`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 73904)
`protect data_block
PRWCrbjUKdE+6ol8Oajw86Dln5L/jlHtT4Iq8tv1O/ggbafVP4Kie1lWpoyG+dbW3++87r4//KpY
1R/fQDCHxtJ/Qz/JiDzFGS/sjNExTYPgIBdHw9C+4/r8TLjxMq8/xX1MPf1BlH9U9Mj5l3eMRGr7
NJuK8s+ubGMaqlSvT+YXvqVmykyr03bTYwJP1KuS1KMJ/M7B0bi6PR56X4QOAQgamsBanhlPBnsa
BZjIlRfBlZRLJCZeJIKPtiN8rN0V9b+ife2YMVxnUcsO1uM0qMVezAT706Ge5em0sMe7zuQKrBLr
72/FXUFAu1yVTuPC9432vciHU1qYarhPDoioaayIUZMkxwOF0FeBGoHvffe1SxdETcWCmrAlBRIG
6JCWG3mnTK1zUQfP6w5iFr6Mn3IGtVcQU1Id+BsMuRrgsXyJS48Rc8uddWOmzt9v/6KlLiXNVOzJ
+0WdyZylPya8XTMotqiWpIFHTH/Kr/6df7axChXaFzJalySs9L3dqY+UgkPGQ3NYVC/jwZ3VqwTY
u6kTFzMW5msjNtRDeF3jiK3DM8srhXzMe+GRuJnJ/R/clrI9PxgN0vWkud9pQH6yxT7djvIk71HR
yhYAoMDoc/Zd7kKJBL/9O8px+Amcmy/YTx8avjt332/2G/8bRPpajucG17SfV1hYS2w7z10cs3su
uECYqiElTORWKJ6BoAceHoHPPqUSEkBeVYI0jcrY5V+c+2EbPsvPhZjT9MsTiP6Y0/gwIFrgxbDj
syCZcPsY77KseOduKJ51dKlaF7PPW4s0Wvevv8GZKeIDm5Pl+UNd80TcVZ8rsKYqD393vudg543S
uhMQ7+AGpSTE1BHEAQAz/sGmo68AA5yDJUARCHrO69OVGvJdScoarJBlMEzKc7nYgi6geU/dt/wq
763D9IgIMfF9h5N8wN1WBUui8pdAoEDNeRsj5DICet6k9rY5YGCOzUvO9s0Q+Phuc2XycSOQXEcZ
JnhVXM8MZF+2HkIoUyIzHmQAgrUSiXQ8rNFoLgtoEkftf3AJ8CLO8caeUGhKcum88pk8elMYED1P
HQf0xh3a0nFpx6odSRT6dG/u2bgBybSntU/1OO9cnEKIIMBPVGkVR/s4C3i5Xb+io1QdaRZP6BAH
ifRhfIf+36WjTRe6klxBk4K9Np/Qq4fzNa83vqRsvuSRV/Clt96Qrd0V62pLV4ZYx+WVH0eMqzzj
e0k7ZgFhvitCRKtlHUDqPhdYo1mo2NBuPp2T+I6yanZAlOTm3Rq1LTrmJydrFnIZG5Mt4XxBbPvR
xPhK49RsywFxWUuk5b6BzJJHYVed9Ss07s6NVkwtPLQldS/PcShTjPYQXTA9pdKCzQvGmwgP30E4
vcH+8vyAyu8jUYmGE3xHZDpNmRW2paBwdxkDWx8bfixFtKIUbNacLGF6ChoiNK1IUMrS0fJ5uWka
VjbAg0LV/ZVzH1uKq6ZUoejycWwWxCPpmLKxC6QR44B81UOHK319xmiujg7OxAlWAf+KWzzLGcEw
rs2tkfHc3srf8Tf+aTOiCbMa0KKzX6FXjO9AaukEhbqE5kHH5ds2OKY8O3ojSgBmfgoY6J+0iTiG
FOkzGcwIEFNqFKIon37/iqbwQuMdLbcYiEfv1FkyhvUAqnp62xHeMhiA68QVSA0xBm6oQg5/ZGGH
KVT35gpWwnKzlNCpjErOq5kQOK0fKxOCegd1l9QYCNopWYMajOWc2Zv2Hy2VunEXGC0SRFffq1px
d/Wn7dgHfNkQtq4sKzUrO1hvzbqqdwrHmZ5L+QtE+QmStR+7/gfrXtAhIA5kHaHUXzKpV8dGxW1Y
/TLjvr3rJzdxh4AtLhZAm/ZrA3+Mtcrcpe9ZiTvqzMvDBZ3pqcMz7JOVdMTDpMgzz+woBJA4rGiy
87PCXLItQS/reDhmhKCkN+LLvPVYZqRVA+8ZgV9yGmuK+0Y3qQjzewltNFoPq8zyWiRt9DqyPlTn
OOmFuS6i0Ui7I9fB0eSm82a0vrgHqWasnRJNYcIUleELCiGtFbb5j1ub+yKJIj3kZs/UoCkQkcDD
U27X1Rkvc39Fagj+3oOKcLCep3ATzZway5OOeu5sQP+VbqX1oPEyAQfOKklGhmN2MvgTH/ew5awn
S+D1xDxCrw+RcZv8pzYoXeRIqIPgOYX2jYXs4SV4Vg3GYKmn12HdV9g90EXzj5AMWRBnIJW36vBL
ESKDR5Q1J2azO9JVMMMeF5lnENr/H7Khqq7s6uD3ibaxn8I30Etmlz1eHC2MBA0aYGE8oiMblBdW
nGcMtcjHI+1f1FOOwmv2EYxfPCAj955BRKEAernSo5xXcDLKIYUGCvC8XcHTiarMeb6Dd7v7pzid
P+eXcM1ZYZZg9tKBSABXNOXmyfZGuQN6zWkKcWngsuUNhxd1aYqmB+Ha2Ww+seuItEbqPfBl7UmH
2dt4bRj8ch1irhBDmE04jEYgquJ+8Y0QebAeMQoPS6z6AecWipJHMT7bkS8SeP1NGWgsx56vb0fV
C8lm7S2qTZDOWH5N+0l7nWf5kO5mujWSMBPNfTWpzdlVyPlc9Jh9BmviiywicEskIN//PNV1sNw1
B40eEjoLWw8cWlKQn/8ESTOCUfKKdr7e9G+J98PoQQW9l+r4RioNut9dwod+ehlH3cPi+rXTMJbT
2igl+4T2S1bjjy2nM7kTu0Cnl8/wrDzXk/5jguDOz95a0AGp70ZHAkXZOpSeo/Q0VRqfuodY+geK
UzPPE0WFQI59iXjWjQ8dnWc3+UMtfx2erYX4lJb1hBBfnTll4CDamerD0RZ+0H53qOSkR1ZGP5f1
CrRKl9Nxia8qqGpdyC5XEp9p9m7BnIeuiBTsFksArFqNU9lH7wfY7LmxUbg9wHTNixm/ysXaIgMj
3v8j4JtwLAb7cwvAS3OGFZ5u0lPmwEcNBfaMY8R9PANIJafgbhNL9g0Hqcqs9lw352SefgIvU5LE
DR00o3N/8SqDS7F/5s34X9MvrGj4As2QCg0u8dnaosY409eFtwyGKrFi9wbzit5v35kxkRuA7JU6
okDn7wA8Df/AkrxUIUoGR0JDU1AJ8kHiF6DVkhZdM1gg2uOdrANVSSmd8Ud1Bz6N5v/0uGkdLlYm
HbTseIr7dxKP6GE/IfY3X6t6p1JUGU4HPt1MVcxqdMG5XM0/lwzkXMkJFvVs8TQY7kO7RLvOxh2y
kxhZTFYMBW5w4VR1Diz+NJNS7tbXMVL0hXJ5LihybU8/lw7nAkq0pUvb5TTvj53chgBx7/fDGOz5
VJa/0vojuW5c0XkTyY+Fj93Aps7gBCnU7Gju4nXmOdtBOUkPa/EFLyjYJBD9tPGMSP6/Ivo18YWi
g7JKTTvm/OnszjT/ksjvaimUfLQjnEQd+CV0rm16J0ZZuO2eiDsn5zOivdNIaNohPhYpnpy3/zn6
aT4ai2z7l4KwkWC9kdvUezL/zeYdrfqli6cz/+5Ry78jTToUigwwKS6OX6eafZVKwep+F2sSGQDH
cJ6XVpsNj6Ua4YR5w45NSSFiLglyRySgnyj17/DATLLKYwA+GbOOZtrSqWjQ1pfi/i3eutacjf2H
QYLG38WMKmsS0lKZUsKYu0ZbyfuD5rL4Sxw/bxI4UPcooEnZj5Rj2ZbwfFJIovA57G1QAW0e0kqZ
x3Oq6d9Dsfzuj6jFCrkltSq3NbiXXzNcJy8xH1/hu4wtNjQbmiCNm0C4lXSB8cb2ILtLKmdeBdYp
4g6nwZHBvBv2rOS5e5HswmoiYOfb29N8YyaibDWNyF6o0xXeE3sixl+B9MSqE7G9LqVPb2HlMzl5
iuKs+YbSsr5yGqCKt6/cjv3iIbLNe5yPdhJvbHFcti+5xdfUFbO91SuApOa4CxehMVDAIBkV/HNN
ts3xPsLGXmNPvZWznQtOqb4csKSx8CNa5UB3YDt48AipJSj9KJeKT+OR4zRUvuG8LQQKqFLhoGup
EHKBuaRcNbNbi4QBq1jgteSy5Ny+JGXdTy9d9TAFwyyez8jCTcynY6BhvcbNdRnoALPfiQ5AYcq9
HBPTB/uoj+O2edbTa6+t852E1tdI/GuRxErPiVAYrfTWHwfJ0kAVAhx/wKxbEQR6xuzKmuldHcrp
qItNxu7vRsEKXVLTJFqTr67DA9q6W7cciwiV2MqipwWdDKLIfh/TI6nps/yIuVvd60R59oxR2tVS
Bc0vFFlodlGJBiMXpLz7WIXyPe2ls6MPa+urMdUJ2W+cx3rvgP2kIKVM8r5TbdxoQHbErXbkJh+L
ShRjAIZtPj8vPedxKv9Q5bY/fEL0+yp3GqXlX1wrx3J3AHa4gmDjBjLTxsNbUI3yr+ZVsZxevVl6
SN+qYWepMSfO+PGu6NCFHPcJnMKOx2tcRQgk3U+/oNO9xVKATNclMM3t3j05EU6rNyXssGhlXKXY
hLWQ7coOS1bbrIjgALpiMgELxeEJG5iwuPIonE6HmjQnw2XPC0diy+h/ydKU/wyLMAfvkYr5MIny
mtOuxumGkROMYsEOznGj7Vp+oiFB+//VaJ7xGhKaFBTkaRSdsmFoqkdYLnScOtrebe4sXD2CdYYl
j2ZfAsx019s2lzliQfcakfMuI0TABzOUodV429sMKRCLLxFo403sXdwSPpkRWuA4vZRnsNH8w7lD
tnGL3mPGyZi1kd8e6vjA5OMirLMM6UN1WrLr2XkdE2NMdJQOL2Tz1fGeAE1gopS1knYmflxQNynE
CfDWpziG8YFRgFv8bSUmr1qAUX18gTo84w5Kf01i6EDZ4XrhprXx9qNML7SRcZ5boROusepp9lSm
U76jqOp2SnhsPzsJe+y78NDKmgYmZHyoG9niCGPW7g8TOnofhtKuvjkKCimrD0JPBrOX+IYKUtg/
gXf5OXJKORVdJQAsfZLWQnzV+dSUCVaohU2R9nb8+joRKPJ16oiy35aOWd0MC9y4My78FSVqg9vf
cyIJ4fmgNM2lsAGnPEaIQA4u31soq51Ji5e4H4rkWunGey+bokmXezF+WbX8bGbfHO0nVfWKEI0G
oEp1O11NiLe61HPC3+7vhCLOlZPKA2BRX5ClU2zI/4+eIuc3FB8J6tZhMxRp5waJ631DJeIYkt30
p+7V2kecUmGk9bXNN+LVMAKEPygMJWiEtOrnGYwMzWXQFzkwDvhfyL/4wMfVnWE6uJ17hwp9Vsdq
koP7ZPBvGsQ1zRujFnNhuHPIAhrUipnkHbwDcpGk3SSLVBS9Yk9+Iq7iWktLOgnRwJQfqtQZPHX8
y5zNJu1Lc4Bx6OPCIi9+ByMQqMSSL/EU2RfFxoCKsUsG8s+5YicvWqKXLeTU3aDu4SizScwOpwia
KbWTh/jjRPr4IIb50rtLYH9PEAMRxVB5/uVkdWB5iGI7FxHQm3X+QERx8amKAvz4SJdUsgmTNHOi
0haPhQK7XTyom6rBqq8c+GZzVrUGf9TR1pba3MYaaYcDd4Rxc7Dszw3hEeAG39rM/BZu1I/u4vH/
WQ7JeugHYKn4KH1ofESQj90ZkEd1VQJr05buzFHbDYmfZV/jSYlDR0XAYpfpaNQz3Sn8zK2Tl5sR
zcBsMGAQQe1k+3E6WDeK/PoCidwjhPSnD2pqeMwWHuLV5tFOlVYfpvVLZLZHMqOFRAaOXlFsF1SL
g4oa+C769QwqsaN7LiNXjclqpsZdsZR4VSo2ekAYo8tnszF2PnswXRxiP+fHgKbXP7Q2g67KxqFy
oAhiXGmM7F4iKgQXPRLNQg39OsoSJIXm5e1RJ6neTJQXdMOrsIcB+15LMMcbnE47b3Iku3T8Of/Y
Jh0Y279D5z/x44iEJF5Zp010J6av9ScjNSEkOxOffQYoANZ9ZI1MqeWxxQtVSW0vyqtzykpUCP5Z
5LvstjTsj6Y0a2EVa5rC+0OOGtEu1UBvyKJ9BqqLxpURYHIWpdKstmPbZHsNa2Hgub3xzoi9IIBC
9SiIxE1VxwHo+WeGqEbAU28fu/jPoglw1HaL2aXhioGXsVCpABnImQ0SAFjaE64BPwkM3N4lc9un
rRcokn16UyQ4/ULJsIKPPq90/zMwsyo3ComF3VdafCaWvbUc2KSYNShMi6kvZgUgviQXjhHarCdj
DHQt4U/d2/AQ+V2eQbUWY9xHvTsJjHY64nADOKmOP+x/rRO+3RaTuZfiWN+jn2TRjWjz0gybWTvV
+DnN/AZ5GjnT1ST1Xr6bFHO9UZajcYr0MugL5aAt4fKsn1nIEJCyKxz6yZbZEqE8l4zvnpcXPFH8
7xVSAJ3KQv7Iu6CZCO8+ePwSjQ3M4LyPb6QWRVqlwx3D4JKPQYaUWrZSIOlER9EQ6/9y1ImRaT96
QjwvIZGkvI/9lNYpQEp2pj0KS6Jz7ttiwBoBn4Mu/3C7GfEqe1KkWPLLbn75mpSSR7rf93bPPE0e
cl2/NHXR3OJ0JNBplgkssYSJvNzkdhyjHcLtcr/7+wDX61nm8ZKBBbKD+qn6Lnd6qEHpzHgeyjf8
YIyBKotIl9h9EGRikbvWaF00RfPKjsZTUNLMdgPtNAZ6ERW8N00MTJLfgvFtKfi/mlOP8pkwskEY
LxmykM7BESu/KOakHGrl2DBnJH1vyYI5+YZML7fhnchkrHNTovRhj2fihO7QV0Rfo2X57UIBpyUy
oskto1hAZXa2ioOcbGc6ZE+OglCckQZeZzXsZOUiZmKKlqMgXPCkB5fg/1dfS7SlTgQlnTdZJ1NQ
m3FYFSVv5Mthh/JB8X2YvaaqyR/zO7NQcAfOYEdgLkO8XmQCRFI2rAFCBc3lefXM+al4iZ4UZE/S
bXA4ssV3U/vK1VvSNFjEYRWDN++crF/B8WczIJs8JtoM9W5jSrmdR64F3n4oneURcd+VDc2+oOfJ
m19hSoHYC6pP6RGfsjAUsAAkeG84bNtFqhkFRC0FitDae8PsZJtS5Pr70/OAlgMtlDVq50kv+L2+
CoYYBCaEDM1wEtvWSV/i868CA8/+1ffshDuLH4XL8pslgjokxb/VILMNyTE/XkP2IWzcXKd6GEOf
D/cSHZRMfBU6OsTPvIHdKo+cx5/1F/eTJ5+66PCUt0qLY8oDaguUytXCWU2Z8RTrD48dJSyUa0B3
YCD2CAJc51m9h8y5LY18cJM/29z9lW4Dz8T4mOR703MzPAGz9tA5Bp4l/u/FEiE8OSQmSKTWT1Mb
exwA8Wqq5PfNeaXZzkdlHOlYJ1/yo6cgndQEIbZpklwc1vXCYn5kvK5HDzTCZ20vczUxK0dS6Fw+
562v6UjYb6eB3L/J2IpbGadmcucOJ+6+gsA6PPL0hIJJbYskeXw6l40Nyb2qiG96aO6FLw0bxJhT
qTSfg7rV8O/LWDzo945SmdR/q1T9tqGupKWkImh/wMtc8rIXg9e5GUo6SR1O6HPBzpjqYs5UVhIT
cjsCjwWBELkNTAxKnH2Km+ij7YLSaL5bGNiNSorgBS3zn9NVlgi3H8UCKr0b3tO/AxO/7UqfdsqG
sZwgrLpPoysnop11+VHsLDJzVa+ZgvEUaL3fKPAgWuQ0MBqsaow+qfAbistNabwW3LfGOpBQgzg1
c0YHXr5QORH/MIbvie7VY3wgS79BafjY1dJAbGxBHaIlhRpYjKoyoNHqE6sJcD+BYTK1148DmhH2
8bNEfOztiyCFySWAXMXBUIEHiRQ2Vguv0UCGi5Bm3a8CWfp+Wb6TbEKIFHrDXqUDlylnNniWaxTV
O0DSkv9A6QmHCorg5vvcS23Tv4RnYggx0pSIT+RcoWCDzTg5RhehdKQQ1fvyqZOcNss2JCXnsMnS
9F40naGJ6lfebr4jdlLkh7JCDu1N/bIqPNqc2v27BYIlKRJZ3YbEnsUBEhDRrYx43hSrY4JXXNHf
wgiop25v6on/UB6+B7NrkZ1o9Is3tU4+zGkMPXUEzfgtmyPGW+2l94YfOKTkP7ak4xv1y4Q81bro
aNYL5SY9CUGCx7xORxUpj1IEUqyui1aAjwnKA4DWOMwRegfulaLIus231tN2ghqTbWPBAtNm2lUS
3RcfbM6y0ctJ/YfWHsTjXuPhwgyBajGnyyp5Vvoy4EeS636r1GkBlFHoHiyOD5oPyJmTJeeAVqYW
H6vZXDx7qc+s4D3lLmvXTknocQFw1RpVbTFyMoCU4kbQdHH8hjVf8r2MrjHeRUHv7Yz7qmhZ6HdB
orXDEqgQcdyaasQUGmXNclJlPHzp5xCuMcOeIQ4pousAqCRUW9xNEO84Uzg8qJeBTvdqpNXPlA4C
JjCNFqLdsxPI6h3wJVTD3ejzs/iAkuL+IT4SwYEgGRsUNgoipShaX9+vIKpXgB5jPcU/60ZKmbCl
Z1u+1C16aug43TkAyXSAdyDQa4F4k1JusWw/uLLbxFVDa0prZoADTOdrFsMxxAPzbz03HpE5TKto
8dn1WB5KQcqxroxGxCnHHyIUAnCJp/AhDctMuhQ8xc+D8DbqyuR5q7U3IzYzQm6qRnjojtbmH09z
vb38J6kHKoTadrdXu7YaruYr+oUxLQZj9A9V6BZ3Wkq/2wD/NsxLDaXsAAKnGHtjLvD3Afp2dJPe
iPz5R98wlTU0C+xaQAdFpqWszmRnktffEHNPCPt8XGBWbTlVw1yQnGP3lnqcIU+IrDuzGty4ab+q
7i434OtaIPa9QUTlmwoIX5CZYcl3iBvYwPtLTljmacVUt0VqKWCyEY1KgylDK+FgU8QW6TXNG4S2
VZxSXz9F/OzjL+kKSHGq3cZNoYBUpdgm25umCm8B+Q+8kz7zbpB9c9lh19RguNjGnkNnOS01X2/5
d2JkVTF9mGT8bVFggTaKLK5fb51fYPf3o1tfCkw3vZ56P4TIOqtAHKiLHAwYuOLwnigCuVTVKPG2
RVUIKWo8pTxF8onkP7KxyKMSLNaaHOoe8QDpzsoemXAYWcDbII01xm9ZgLXV3LGKZdXGVJ1ouu++
eJ7h1m7F1zM8XLMYAIyCntIKAGgISFJilYlwdMUb4XBj6+qEeWZ7lUJPIMjlWpFtOV8rJPw/jyw3
ZDl9Lq7JM9VKyVRk6v5Asd0Z4wUnOCHVmZ7OatJWXhVeBQbksdLbMgzIHGG/AIr1sd7/SSzHotfC
ZJ1KElr7TXJqlnKZGzRJLDoPKP7Z+oFgecTACUEoWAN7I+97c5EacaHG3+eHhH6Qkh/X1GOe2S4p
i+lSGjDCbT48dxf+fulbRA1Zgang7p8DvRF5X2roKo6ZHivN1D+HU2u3/DyANsvQREiFUA+4KIl9
udEh0aUw6SFiji2uc5E3rKJMX2LR/YxvkUbqtkAuO4WaAtoE0/ptS8tXRGqUW9RPv6a7s4rAuPAl
rFr0H6tiAcERKnvvAr0jCjHDtfj+YJjkXHZk+FNe0WCoUGg5zWCtkRWq4WgnRMN3OTayZqFJlfEG
Fk/b4f808O4QwB5uKE8NZygzqjdF8aefowEJ3zTqapKc/27zL1TLDeVy+T3+v8czK4+Dffmqcr7K
Hlp17tnMApXGRawdT9w4oFm8qx9S7EOjUAxa0Ran/MGxUaySodYQIQrafVAA56BYlZi9db77AriH
UYfRXEUGIlRmBRfGsVO89/lrRQb1R55myFFef4De02ARC9veDjzR+QGuheSkJpCD+JhB6J9CHVyq
Tc2cECu7pPFnnS2LzIk/WcsR0go5+pQZV+6BBVgJOnqToEFESDt4BE9mutCxJXnpdXjTZJwRT+eL
FnFe1p7yqhaaBMn8qel237Sml29FTv4SiEQRYL105L9AU+BW1RMGor5XpiglU2L1dAftGIkcteCp
tlGPXNDu2Nn6GOTVJ9A5kQg2gQqYzBa/e7j1pu9+L2yxW3SheqcQGC3Tot2Cn0/E7f5XPgLfaV8X
7s/q9ATAd4l0ITydvEiLep/FbIE7ZQsb6GXq78FAbqBT71ybhNCM/2k+LitcS3AqQo+kADlVLDwU
35c3OMsmiEf/AlNyT8wHI4buJH59pY6ABjJayXZlglUi2OahYgRPALYuaSF+T47f8nJvWa67xbSD
bz1feBpVUw7Nh8y7PCRAbFORsWBvayVslLqqjWs0iZrXXRiftb4U9Yb7HPDgYlFz4fLXKpgGvKQd
Z2MjxTxSXLfaKQwLVchhIcvF0TkLbUBcnjj+FlglTN1Cx/5gdlVBSbZu4hosLumlUtV06/UhIaVv
Q0eS5lX3zvGNclv9Y2A606S5C1q8yCJx+uKGuvVzpatNUE1QkGz+Tc1Xh/pFd62cy+sQWnMtQMOJ
ypzQui8hHSkxpAi6JgHHOIyZCvd941mX+EdvdCVLTs8c/NVjxXxZARW2Fuxu7CH6sfw0rOV3eFx4
vRI0JG6nKdVNC/+DnOx+OI6Z+tQPd0c5tZYmSXzNaDG2bKIMD3gAtBc8ewjhQYDwcJdQIzZMxgOt
2s+jW/xUD/DoMUqN2O9xX77VDtp4kIfmAj/q9WNfmE4rFiUrbSKLs17JZGWrQmlFeAwX6vG7IduJ
kCpCNpC8hYp2jHDzNSm075qHlwUvtrl9TB1pXDLUF4wa2Ceduc/mF5kshohsOglfDER+MejFZYoU
blma6A2H2yTOC1MjWAbl6tsohlangyymk8kCCA+BPw8oQcW8E63J7WKOp7s50sZ7oz2UvqDHiRsi
oDr2ghXGMCJsLkBwePHACYbWGL6iFsLZKKe7vA7sLTDUzIp3M+JrfORWjQcWAjyeheTnUhNo+Xq6
nr5stjmYIY9xsRp4eb7On46b4dbz/DmrzYZ/zfzBBaKxmOSQp69A/gIclYUiUEP3mwssDC/LEgPo
zc5LIRcRPSNsobr17BasgykLDJX7tRBknEtNTDTf+qZkJPrxa2o4UwYBJo0AoN2VfJC+Xk1aLyIi
sdKf/p/Lp2ixr73+lU3SXckZ2A+27pHqzCsXbHxgvGgLVgAANSxghSIbN91An5L/U4QwHB6BquT5
juGJvu/FxLrI8amBz7M2EAjGb6eJeIVXQ8TCkR/2EiclNiGERDQzbtelNvbGvhWx5QBk+iiYqlx6
bNwOu/f9um5yEhMd5HxIBbtOeO/9HxfK5aWaAAHMfn+WFz8wGkOFkwlt801MKEJl2WxEgZCJHPDB
/m3aHGs84ZiHaFVueaoIXPm58UuZHg0ApRoNhwKbjKU1uMoH2x0/qpQeg4NWrNBepxK4U4nH6cpD
jpRMIrEpPfVJOsufZiv1EQiNeFk97jGddbbD2VeksGbRTdPuzZZzOGrU+x6+WIj3obgXkBO4M+il
JuNbk3zsDrCc75Ud30qd1Vn9VDrP2qDxHuDFdyHpPVb03wt0x11NQ9ae1Qv6QVJ8jvGt8Maukiza
6/hx5enu8XQIQLJSgIiJCe9FDRrB9g5eHSOQ7DA+jHPND+O6JgQq8prKasEDeH8v2sgfgp3UXoIn
Vi7udMGL0Ur2ddGGRoPkBt6DhDJGAVsvVT+oyU8+C/m21saWW5UiqWXbc0+E7UaKFrshJlUhUBUV
mvKEfytvjaclTKXJi79YU8pvZreYpvgdrcrvCLkbSq5OJz/yswU7jOIlftzp8+hTx0KNlhlZYTwW
WE4hQ6+/ZffMZpCX8Elc3NjTyHP9fhsA9P28sFRnp1yZOZjtO2OJ/EoCBWXZZOv7jJVYDXUEVhSn
N6OX8u0V39VQSiTUxpWEJzvJ7QTGRRaGp307WpsqbutU+nhoaVKBHVytbMYUaZEMgPsIzhHZsRti
oAVfS1FrI8nL1iKijTDxAaY47E80X0Wx6JWML2i3ep63ZHZOMCPMyaNbejkOLu65Z1lw7TzxHrQ/
zehujbWsGZUP5KLUzwIJB8x7cV5FrGDrnCaqEH4YoCObOXMW44sAWLWUkNJb2WwQd5tWHQUU7i2o
2qBkSe6pttpOsrg6QdY9UOh2JyQoP29fK9JgPlGLEaglWAhH+854cSCTAzzMPiUcE04cIkpWQ9gJ
mo3JmZ5v+gn3yvem/KVG1fixy25nIKP3gDq6vvLHeuIIWS+lHpb1Lq7YvG+NYd8+pIxojlq/aU0n
R3NXRauMIvz9U/1hHOx+s/mWE4ub73I/kgf13btnhbLpMcdUQ4iwE+nhbaIxMmprQAI/wm2dhiLP
pLvktr2TS4KzKgvolIQ1RN0JVCgsb+mZzkXFcVT7S35AmyfpyeSVCFTIPRHQHPl2hXd8KHTifG1f
4WKGW7r1gkKPTYiDfVIVScFc+8WISKg1bbefm+OvIOuzJpt1KSddK0wh0kN8V8nFIhQ23dZpD4Fr
XUlHDbdvTD+qCRVY6USAO3zYNJPEYTVig7hXXC+otlR3c1X3tNXHP0Qv+i5YASFwsmEAmAvjqLN0
63EXxBPIExQEmTBEAp0W+Hdi2iemZOg8csq09ILD8DdDOzEWCMK6e/kkgLht4AdoBaGqenGhP6Ir
pp670pP+fRsvjG0o7TEdI4lj9MXQ24jI0i+VdtPhE3ED5Bvlm4eARyZLeGBjkNMvefSRixUh/d3N
dxv1cIunfQz23KfmmsX0BSI60JqNMwbVmOr8tDmF1PNXoiIDXHHyFsr9eBYD1WjuSHScZ8ORu9XL
/Wv4++Lob3WowYaRwcJWCsYZTCOaJzU9LJhJLqG9/hojgs37b2o/C9Ip53oSdu/foB2AJmDj/V4B
k+mdeRm3nlq1mLks6mzj3CXkNau5jQzys9SV2YahZN7Ay4Mj2JtCgSarYz46v+MxWqYB6B1LAepx
X7Lb9K0jsO6ZXSSxGYPTEdusbe1DQGVoiuyWhrjtk35V+ivMLk+IYABYic4zcs15N1OZ3RRX1QLW
CjxT/aHTC/bAAelg4uR8ybpMixHyzGR560gCq766OK6oc64pxGaMKBz69OanOPeXOLwMXWpXNm/W
Uhc8NAXB4ozx5o450FqSuALodyoyP0U6vrV8b4IIf+hw5CIOcZL7ourIU6Vf963+YIR7xhbm7ZeW
3fNOCTpwoe0tF1hIcqFaW70trzVycZWFkqHpUQMIRWISkkBpmkkKi3h+xWAcDw6T2yDmTp0wIQrX
6QaKZ84wXZQ9PWauoagRt2HvJZk7nPOOv7dG7qb5TGl8TwS4V+ypjw/Td3S8/PUZ6AdUfOECDPkd
rS/t05N67HxuCsNjZQnOHk8TbiExqWHzl3SO6kG3DZtbWPlsSfvzePCCE2I0YPnmbzt03lh5qJvE
mzxursRXRzigye3YFzEy6ZHCf7xDbW3GqNQ5HxCf3kytMc6K8Gb1zP3yX+eXf0braQIPAnb18v4R
iQkd1Qi1No6IZKsOOGV6xuWfqyzm4LSIMopx8qqKWlgM3LjhW10FLlAkY0pXF6GqopSUK7BssEzG
7Dkm+n8i04r6jlrkjybLaq3EPhkYoE6z4NxaBJ/UchPwWyFwaSYr6O2umtIvv3OZiKYO58lPPPm8
Et8fox9W8aXNhp176RelYtEybHM1u45cLAmfliibel1lOWEMpakApsDGVy38qnBcg3AFvgjyOZvR
7p+JnBkam/Y+uOZkgAcQ3Reqy9GTeHVsOGX5hfrIzrEUJT4rrB5rjXsgERkII4eiXyfIbQZObMHS
z54QdBwRp8SAFf3L3VV94STl3wXTMoAfuxR55iNeNzPyeLrwHYgPgPAbpcDGuawLmMN6dLVPqRBC
2kFj5Zi7vAI9wKfcxV1e+GjkDoMs2qNqrMHU9wztuKBm+CEhCXzwD8gEmsHK/2AgPqcR/5W6hR5X
VoMKbBMarFwUN4L3QmrSPvM9F13bqZXoO95Tdt5XjaYb8B8BeXL82iRTg2zJwYuuY0AwHUA4Egq3
MZBkdWSsGHiItjh06KvOjMHLyKTPAbWJDF8YuNtsLQQoKgfRuNKvWno83/GP/MbfI06vjofCjPsV
2T4J5MTsVJ0PE+ogXwvkmDXWW97xmvz+DN68G11WButB5lPayxShfJFxdBkQvPSzoOTqP7ZipOXJ
a1LRvABOCnLTiXn/TGwnNivfV6yMl2LeWKR53xpiv+Vcv6nMsVgQE/llt/ptTWF10jM+2KCL0efb
r5BhQLNLyVJunLbTBdJZThjjyv4nnPA80h6fDcikYY62gYzspIBqWigTCHKFi4/tojxJalllwcte
wNxgI4N1pLlzElH7fo/SwHDHpJWiEkJFxImjlb869n16vWPpve61qIPBlf5VMCNT2iRqaHuqMsTO
A3JR9ZU2V9AS/P58zOw2PgUNKsU8KDV5hS49qHBsYRQYmHE2fUWt/rjzoNvynBSyPxORs7T2sY82
bnsrXdQO5os/6P9jZO3yZzr8X7mL3QSxZvFaxgPEOno8038PM10dMAC7D0f6xWB4r7FeCbo88i6K
exH8tojA0+MQS6RzxKxXJ8wtDGNXak/yOE/QBEZerMZKFoPry969B0UjV8aH3u+yqL4fQIpOZA/c
0JU+yOnoImKUT6nntdvRFxty279HGSxS9e1dAI/+DqexdTUiKxnLmO3gnrFmEKo+dUdqNX5p5Hj4
kWjO5xgGIAjJGwhtRrPS4Bn76AhkNbChdxR6u/MgcH1gd6WQgQxiTIQ1EnI4q3l8rCc1QP3wJU+Z
hZ0imSRhyRbruIGVrymWnIhFhSqBZemb71sqVXFdyWId0YKcCMXTzryrQ14RpCqD//5Us06KWVFO
nOTtgY6jIHqlmTfYk1VgFgBqvR+2AzLh7a4AptnnpVNXikJGN5xu1KTmXExIurM2Dy2BzfRps9t6
OOhk+p3EzQb9zQCA1r16zgP3jCbnyCbrx0QITjLPJ8pmo3fFBLMvZ1WRyoVlOaWX8g+CI85HxnpQ
4MfaPCK6f0DHF1C7+yyzm8BDU3Vso4G5zx+hvKl+t2XtTK10NAw219qf82vZU9hHpJuaCI33rb64
L9tvAfFqdHKq4xJ2994TLDDm6LQC1WWB+n1haYCOSFm+gr31bA6FUQgfPqOzRIr1iC7lA/g6/ASU
r8XmQ/TvoOnW4Fgfkvmv/Xcp9g0rQGWjuePKz5PsrIVLNJFgdnxR8X7Few/VW8xtlOmB7m/Fr0Gk
O6bOc78AcTmPrdmZZ5Iwx84l1Sc016hdoDT6S3KlyY5Tm2YbVoXcuZvUhBHbXKb7moAI4Br6CMx6
QIklQ7TJ7LBQJdgeno4z/LhnXiJqKIqkJS5TUgvgfjOd99Wf/loQTR1z/vp+zA4AX6l3/EI4lyhH
HDS+dd/i0I+zhXXrdKiuGnnP+z5OTDbHBQoMrtAwQDICTW9LBtQMeV376JVTScdilI+WwGnZYhLN
FU3vitQukN7spEqiQ29A8ZYvfZzxHYOYF/hD/H/Wrb1c+iTmiuEfW9Da5gWNqhmRbD//IR0Aewgs
tUN2XxNH30bgtqHDb5+gxBztrz+prbV/nDJtMRXP6F1IvvDl13kYR8hbeTXTbX9dqfKUBdzwovi0
6u9OFPKOcxbd41JEyCJDeWwSMGm/1MVflGNkCDjHLWCWdutRK5uo9cMqyJ45An1eCWJq1RrxtVic
vkw8B6xZvdB/pNSb7r+BeX/CzMPOTmhJW9zl3K2U95dHwmybMPAO+aTDsytr04MuzUs01sjyvUvw
OXt2GrNZicwNw9+tVacs6DpZ7/MYTyhCLclknzUTsGDvzZfOOhKs510Soq7Kqj0B3tTiuZfQMPa/
+kXBfMyeYMVz73Wjf/3JveeZloXC0DejSc5iN38L1DbMryYrxm736YmdU70+MP+UqAbyol/6CsK6
jPmHrXdAAEV0TX/h5bfxjPfp6Ai/+KkoAXXAI2Gtw3b38ZCUaZCHmBHW94qUB8bRcu/57HSiLmMg
San2gfAJ+oC04aLwKnzUfqqkjGnezJQPkjV94S2dKykjH0uqT3wWAl+jp4XQvhjR2gyfz5dsbtv7
n8t7HZdQJ6dXHRO0nGeaP/6XZXCcnMrOwoTrWQvUHsBdAetCJVK6Ey2sWXeyOt6If6kk8ohe6Gml
8z0g5apDczUgeDCwMWX0lFujX+MoGIINOHBwgQPssoQ91eXBqnD15agQ+dHRtqJ4b2Tpw3Z0EqL3
JgKtRRv5jaTY+wuDRoyi6AxxN9DfiGFXwTTUMSTyEsu3Vhlj+JFFFxGZAEvZh0sCpK046E9TxqXW
kx0Bdw+Fw0vyyEj8VbNGyXqlaqbuq7i/OGcx+tgP1Pdptudd+Jyr4dyjqpF+QIHzoeAuD0N8FsLf
ZBVcIOnFH+uyKOUNLTDP/Gxwrk/lRMc+BiMOLq2riHTUE5uu4vwypyCWCjA1V53boikeqRZVQzAS
Wvfbx1sQrAE44o0K67lsuPba6CiUxgUU8JoOXFcaWgCQkc5HdEVCgZzwR+VUL4+VwXUY0tUWh33j
OKf0pryz+LqQoPFXxsFv4L9saBYOHmyDlUOgssfNm4TjjECABaYPtYvo1Jw5DtSSeSpD5Z8T8CcB
wwVNOukofYMnVnXAH8o59j1e3EIAtfjG9H1iDFmgIaZGHFtkUWo68ZkyWeNLkiwk+laGUajmQXuR
+ZfV+JPalU88xezpanttI1cjGphZ6JGLaOcVgUMuOf0yd57Po+w5UvX1+7g1qheeLQdY/fRpnUvh
zzT8YgdzXjEgqLAvoqoMglDlNJBj9hTNmHwq1fSzhRhKEUOJGz7Zkqctgayl5iBO+nztB3xwCEA2
MbxKJp5/FJKacX6uoXzqV23ZincZXFNMR9d1Axm/lgU8/k9BDd3Ul/qJiaJUjWll9O46aPlk3dFj
cJfdPZwkvtNrpFwhABWVILer98K7yn1yG19WNlBmzOai6l4xwwgJSsMmz+GWlyRDb456XPz2As+S
i0tnU/E3Y8zCYMrbRwmXjot/w09IMfEr4kdeI8TGkIf0Q7aSqQzOKVvV2uCkaoGkUezW6r3QYT1J
HAT6heDFweHUmLDnZWYyGZteOimWJarR7NELrD9exrLyK0+DMNRB81KkRfuMR0w675UhT8dENZZ7
yvDhpKohRozGS/yUirg4NCALzYlVVTfcdwh5r3a83ObFz/l/Gbqn6TwuH6b/xCrHwhHyAuSY9Wzr
JKqBdLBdYVAUk/aYkd4ugj3GKxeT6gJgL/P5WCmyQiU/0xINgimK/CuYTklshT7cuBIJf7mFMg/2
uiy0LieFNrOKwdoSD8K8til5ZHClPNCg+juv/5a9tp2D28LjdTtbgdr4dVXJeFL6zy3ACVHfq/U4
q6Wyqxts1WeWe0vUFiNt1MI2nwe7UpbC/WBPQGkYx1n2zHh2jASELek9Fjez5gKNt5ioyM6N1NVU
ELjOhfL80QqhjBSC8JGpRBzRYsuhhutUqrh/ZdSwSy4CF0Jte+zfJ9pJg8OI0a79Gcjb4Z1DZbHa
h7bJfOv6QuaALcLjtZVeePXrfI1LCP2hy2Z08u4JxYm7SRoLxqdyyxrPjqGa/4ezNYZU7GX+ZxJk
Lgu7KFplsUdWs3ViNBgGWFwtCc0Sp2YAYmtSdd4h7tiOgonn18ucjixQlhOehCv/3/l8cpiYF1te
+uEGMd0Pw3/uB3a8qTB3R/EFKUFToNmKv17JtiZspUQjoT4+g+k0eniDOdj/IKIpYqlvv0QUJkZX
U3QomR6JHLKpMDKpokEqGw2Rf5ZaZ8wv4EXjUN/Y85r/yjjBNcl6Sx3i8AwRGyjaNksfPgFSQ59Z
gijb+kj1kIDNM34Fe7GOlh+uAQTdRjLKnsp1T8oYDwKiZe9FBDPv0YagluS+iAThhTJj4XgiFZ1r
nWZVvlXe5bpH/EurGUYx80/2o4hSXOYFXdfGMQ2k+WtLRmKtiMpViYHqpHlm/7xHJPMV9Aj5rcYR
DyKEdiP9Wk1ENErTeNE9IKLWOa5ydsx9BPiOUpoUJoHvQQH58nWv12nJDg+zBuNQmpdrEulgApN0
to+2XFuTYs38bL2x9G43zaxRH0PZmndfTiR1tw+k1nLe4acszCNJ9zftUrQ9ptMHxgjcz5x1YBs5
6Q4nZExmexKhq6VVV9rXv1ndifZFk3v6IHH93AqbGWF/9IAdEvP6/g2uzKtprn/5yDitczi8lV/S
kozobVazktL06il+2p0zrlPQJ95pJ4ezCwKQY/hXoMCra9hF9BPBCbkGeielOwawKeDRfJmOuJtZ
W0n02wlqzkA8ITZG1Gt7+1gSrqEcOnhNN03nR5i82vIR5z/M4r83psvjVzYlLLFOx5tH9jMh4kfq
xq3iB5/XZx09aaTHpS3IqxSEVVJea3Z6hcaX6HMPRKdpttCZfeWc02INqckbhoQaWERi5JJpvGEI
jSwO6VsTbAI2is2oIrSEv4D4wOMi6BWQRU5cCcYdHcLZ6v+aK2L+VGOfPrO2bW5KLW4ke7tHULsV
4j+J3jQiVMdhGExzlLrByRhRkDsTMkdOXYSH4AgHX+6tQb52ve8+GZdQtMBhia0nQlZioS+FYy9V
jOUNUJG9PrlpFeXDQqlQTkMY38/jg2SLQ3jQYlgczqT+sDgmcYFaL2iEUZr7vAWh/04dU+xSv0Np
Bw+a2FerFpK+2tuftL7POFl9UMynwdcgQ6+zhmbpzpEwEpr6rE3GZkVXMf6cI6/rHKsm0riTTR81
E9ObEiHpNqEbcEMIG11mYyc+4KuSX1aHmqvXGBmYSHwiAsmo3OenVAsyR9Fb7h9QpvJOBec3AGBJ
N9FeyBNQGdhTD+4+gSqs4IE9/QHEucMaNWpHp7mimWExb7kd/lA/6TGqA7bSlLtnPwMhaaxXC0TK
LeUzuSEA/ZiT2T99XGVJ7uiLzG0mnXO/XVrGJkhktLhvgew9EcF4EWsyXnhgAV5XubHV7qVxzlnX
xyDScSUdAdDoqqSGvm5NzuvgKujcZyqpjJ+qeYqAFQHwAK8NJDDFkxauhp77n5sDSTc3BW73+I1q
QLrPfthY9bDdWl+jRTJ7bTzsoFin6dJN50ts0fEI96NsiAe0prTJlHn23qVK0KcmvkuyEWNjAbq5
g3SWkmI4ywXDm7vIDntxfNIezopaFueWFY6PAYAvWbKvNPlLF2shaYNHUvTwlKIOa/8TM3SLvV5w
CX+528fpZAAvkhamMtBooKJj6X/y0RQSO9m+sIqTUQYOWtiUrE1TNQStQcAJdzskrmaaIjAZAdW0
fPqGvAVgxKsrUy/lpfa0MCeHoKxuEMbW/YY6Y1OowV2koBm1zRJQ/CqHrej+H8FmSAPEO/FfcY8k
J+EV3duG5y7EGIHDLJnMQfs/DdFn/zarjJG1sGJaZtlRygoGQjOvzHXIMHzl7ayxhaXvKAdWvN7C
Vsjnz3/3+2FZKNEIqhJaHBlJl6golK56ghwY9TxrTfNRfPlLwe4aiFAY1YUbro2gz9LAikyMQXUX
e+Ne85YTbcfyMVfiJqUNWm16HD4C0QIMEbxLBSSPelr9VQBMDVkl0tELYavwuLyp5mqJRwiGmjJM
neWspOiXLbF0wkPbhwsXndHZAnr5xRWeiaU/9+QJ/CCstJIDhUrkF9N88abgletBHFHWLWC+Ezwd
jAB8IUuHPhtVq9YLwzbPYzLVLbokPMyTksF2yHwhRJpl9UZQRipMxsRwjJtT7BHI5JhMkwp/40N0
k1P05/lH0eWvTxsa6rfPqKtdKWmU6XVMrj5Txiz+o1A07rEGAfhC8v7HjdQqtVljVyBZS0BzjPxV
YG33iRkXlyaqbIwJKh3IRAVcYxMG9EQ3or/fvyjvzQwQi6cZaMWSa0YDSeGeu2dZ3xBUfxYf9UEs
SO75qPRKSNg/x498M+g9loi6j8LYbA9+BeCvibELoObLLZn2J4kTe8lrkoRV9l27Jz1V/gcUhlDj
V3Kv1GCKOeq/iKje38CsG1gJArBS3mGPnLjIZxLiCivtbYiZ+JVTB+Fwk2nKy62Du3ZjJCglLFuS
mKRqXUoC/jhVRzMvp6iIMwiUt5k13Exw8RbZZVxatdhzyJGTe8m74gHL02wt55IqZUbdCeDZbv7q
VyE139mfcBZyycPO7B4m8BMrbBzR9LWrPhTo+nsgtdPhzq+NsO6B4QcV9zmdrZlXbvFrUYO7+B38
0rLO8O0/c/vqa9QLpar0Hiz/bhiVZJqdxTTplQT1O/ScPHzBYKcllBMGwy81EAiml2MPRbzDGMEV
kcqNsF7Y4ZA1RpGoEWYg3WCgPoatXxKyFTrR2D8BszGBMGsSeRENv8jy7qIegJQkztZ2uB1cC81T
MNnNw/tuLx1D1G2RGa2ZN707CrAh9WeH30qWBs/U1sEkCbsaQivkewF8SEQcyB1Zw7cC6CP+q9Ni
jkns1SBOZ+U/YzYKV8M6v0j/nDmQVbQErx53ZN0Qdaon8KhmsiCE+P4+vd4AHAcsVkjORWpoIcmB
u56cvtQ2HZ7wAeDZrrwjl/oqp2r0YPrBreD8CrKtfXCFJKi8Aj2eFWwtq5M09IZt16c3p99HDI+F
QhqQ0jMmADD1slIUNWv9HFYs9RUAU4RaJ0f5XFigI9TLl4NC5EMziWtcqTvFjvHw24w4GmPSuQUV
qxVxthdMHjheZtCitFThbspuYDbTsqEHHfURhoYq8O6ui69qTLpXlnZv6eBt+9qHEYjpyLQIJ+vr
RxD4q7mPGeKMspDYbQvjPvNmyhruVlG4RpSuV/7HGqP0H5BGvBc0P2vLo5Ty7bTYe3I2wQqdoEpX
FteC033nHAtcNBCaDGqljuLqn8iXb7p9Tt+Hv0GJFsN95S6NPSlxm1W8Mp5e+XhV9aGuwJgYT9xb
FLSjr5cMDxlSGk18BGHspu5dlSvfFS11k9j4F5KrzfAeHF6bwrlWB4HA8z6/aPrjrnasrpcqYsfQ
ilvlsPK7eJdTKxxzgES7dFSEwIsb+CzMk9fwrbI5DRxOaTmYYPjTfLFbnyHqDgdAz0hpidPs6hhI
XrILjsf/BOiJdkvx/pb3U86dJVQkd6c+N/WB5WLAgb7hzyf+4l8s0I7Qdu6OjPUjfYdWXV8UChK8
gbpIieh54i6DUzHLOrgDGc5wzCaHb1VAbfN3OVVtvOgr8o21UvI1rsqO62HCGcthOctBNkuo1pew
T2NvDMfBUydlLIEm+mY95DLv+kqV/kA6KENF9cr7MbJ0xr7g7r3LyMzJ73p49tAs2oPLrSnutIgm
NSXy63UopYhdE6OmxENo5LHdyux9TScg5KHkMDs8XnHZGRYAAq6kHkFQ52/qtkIekBOAPtsw2hm7
O/9x/nI53aDrs1ghLaP7brqx5fH1qiAVtKmd0ZI0kxlY5p+ELKlmxaFOgxlw4hMRYpHZ5GqTS9/g
z8lsFKt/WVZTbZJS4Blq1anIYR4xMgTmnQTgmrjapzfrJr9ww3IweKOZK/LKJDcME+76sC1czQuk
2lSW0w3ek650S0FSkJXA9/Un67cnfRMgdP2j/cZDOwS7Eh3Fe4llQN4wIp1ZmJaHYjM0CJkhkmul
RG2+YPl4IIZLS5AeVw5atvaOq5ITIPwP65BK7WxQIxDgOkIXnerHn+IaxDuv9498eNDNtWOqEuam
baGHdMDKyenfAAn2w4Jwtc2qCgNRRO3ACp6myXVduqPBosdyJosFxxxEabi23RU/4I5NvJCeJJzR
syfHBALl7D6MrimiuDVPJH68JLiwW2j0DL20xje9MhdUtOcmKgS0R40scy5AeZx5dZ8MEt9HrMAd
SIYHB9k61qXHlukAI+icUl8IoqnIY9r+2rEDHvMm1W10EkmNN1c81X8Qcut7H581SFyujNzA0yeN
3FgcFkfEL/kQiVgK/53yNgKdrnBTwjE0yweAzVjzzS2plq7RqcQhfG/dqgu99Lzh5FIT4Rbg0muf
14EFJ3Yh/3WEyRl4DpFVOc8qL2GntDcd/WfHBr0/zqv37VFsfuZQUea1EPwHSbjsadkJ30GdPndm
iCMjN9dfrAQ1INcvLZQpB6/9rKHZkGOuKF9ROtX2HDydZ9SlyRht9o/XlGsju0fMKqVSjb1+VhWi
DiEfYiiiL05YV9t2HM9L3WTZKN2vCcY1J2oNOJuFycuq6yckehRq398R6fVzZs9CrJQ9QBfqunXY
zEOcDxwiei1p5GU/1c/Uxy2hASrKQB4x1rFX2fUtNvp6VnPgi2xzeM3lUDw6uPsq4ONeho87xqnv
LH2ljU8OyCiyr0DldIT+J+Z4EDy77LCt0M2826tAnEeMSjetU0IkGxARRI+xdFAdXVbHeIy30WtZ
gDzTuF1ossLJJFkV13R3ugCO1M3IwNIbDdHDhEg1K1KJeJV9rH866V2PfjaUnvGs+uzibsPgH8cc
2c1rx4uk/Rs7CBqCzgeICZAjgZOeU1841bo8IMAdvLY5uwzWmH5AVIVmliVa5zo7Pz8/gatu2e8h
7ZAWsUYKyMNhXJSMhxkjbOezhx6/+Un0scLyCYAxsMXxIDM/SqdYGAzRBTEs7GOvqS1GhtYygnJT
txDfaJCVOPAMSrFTTMVVPNCInsNUwPBYNaDZtgS+NehfeKxbnFx7srKLXgQNaFC9SdIdCDrwBqfq
Vszx2FkCf+IyyEVvyYibqdupBHqaH7ysZnJhr2Kh9vn5y9S1B0hvZ7udXaogJVpBjw7szw+BRvAe
rP+BYmV7sL/3I95zC4YMUrJxJ/gAMxglAherz/uco5QybAtnAvAjbxIEGVaoH9ihbHYfezqOSX4l
AWtLyMCD3W+lmUwSSA+n+5YHee8W9kduQyrA4cQr7skm9nltxg2TuEQLWSX7po+u/wR0LvBlJ19L
H192dEbCeKhP42/8Aqo2pr8Abd5vTFKwpHIiexxH+C+wtOonn7MUm7nao2LpCyy1B6NUYEiBceyr
/kB63DFKrFPHQD8OSJQFAJcNh7xNURCaNVRPlsTVd10AUmiPHL3whr0150D2LtHh0mWWRyQeA5Rr
MkzadQvuzbR5Mu8EGHE2F8apnrD/gE47l00iCbw1xCvqlOFKE17R4yRJXCDJE/IfHxa79raimLRI
x5tM+ZdVmMuxyUsM/K9dB1VNrJV717xjYLooTrhVg0h619X+o1f8jr7XdBAt4lRYsidIsJjyVUYu
r6aBSc9OOKREKO2/EH6VE2P77WYHqSc/T3/g9OFwNk5cxKb4Elsh2HIMJ+FauNv14VkmpVpc2dr4
tHk292+eZlRj9TZgW1iujGYyCM1oOvyW3klA3BFLEhlxfdS4LPaMAJ2xcQUIMfWzKiHnie0WxUaN
NHGsBXFFDsfCkBBueh8Qy0J8nPkqEedj/6dNXHFVP4vAxN/xT4jto+bmqIPj1vYQe18JVtIw+tGM
4s4/bC08AuzbEW2cIAdDPqYmz2C17KKnHHWMBmc5Wl9O7Lw3kFu0I9st0emFtHHExcICl+0palp2
r76lAX3I2b1CqyW+GrDldH03szFM8FwJZAs34fjHdIypVkp+Yw8xyuivLL0f7EfwyzPKo8MCpEGS
n7QHj8Tx/zixt+J/EmObyfBCloParzGM41v6WAs8vrqyZqGWjx4wA9eYSHiW4iecUSTVQ4/xw33d
SvyyGn9pVolhAglGT3iG3YCh1Bbai+2akS6DeJCmzzm1GJgKl7zvyW0N4RdQ//jIzPpGTkZNylh3
DRMLkx5904Z0TlRDd3D33Vn9Bmnn/f9YBqPq+O+2OEC52N6xwlbRhCdqkseNDzsMbh026j/+7+NN
VG1mjCT3I08zCrRDjc3i476m9lCJeyKpLlTs5tNZPSUVLEA16iIANUD+1tbZZZ7xZPmSVblHbfmq
kEUHDAG7ZDWOBfvTSE9PmZFJevZfXdPkrmsAMhYIcgrkXvdGfGulqs+ECyG9aA+U10JEnQqdU8JW
9RtYKpoYY6x3OpCGoJ+yYk8T8zLt4vUmEbMNnL/pIy0MgZF9i21yCS0+tYPSHfq6d9RqreQeZl7G
9czC9qGQudyFruI5Soh10OhtquReu6cg41bNS5TPePTw6D/MMbBFKxYWSyCQ1kjFROScsPPRfS5P
XQksOo12kfxMKHsMbSFYSmEPFY6Fnv8csNfW4zP2m4+UVP6ZF3xF7VyVb3Rnb4NeQbUL2IBMFxcM
z/ATmN6ORgp1+hiG9rKIlJHJaJjIC6xqNcqflk8sd8WPyVeIEbcijLbcvvLjZPaOW+huKscc0bQf
KxKZ2gKmUFRvwqyf3QME2qOpCQnZTdfZEsgrhjSiobuQfVS87uRLa26XS5btCdkGA+OozAHRYEZW
9Ty0ZuUjLU+aPTwDs6gp0L8CBYlVauU8D6RMhQRow3r4JlUHLznNv7sXgCa7yscFMVq/zboj789J
3ZJgz1o7xx1JDaaUkQjm1YQi/UeSZBjz0rZLtlllSYELBMnmjfnilo1MQidqVJfBVZHRXY4PNG5y
NLbSsz6RursyDBtN22FIQpOyExBdXT4yJYtV+VGKAAQ3M8gx7DoxRTDCuWeMsvCOoKfnyKGImlaK
wJpY2CzIaGWeLGSayhn/OF/wJEAMyUj3EVNWAPl+jj6aABJ5KkQ3j1DtVev/Ee7SM2DlemmuLxY1
JHNg71A3I5Jld5ksSbnPAGbGACv9acS6X/47fi1yG6bCGrrBZnvVFTJ8JbIyvApUzt0vt1VpyZt0
1tPtKs+U3GMAiZgDyKNijF5SnYQ0uOgPeq25cWj8dzRoCeGrDguRWgSQasLWtibIyvKP5KT0P9KH
czc52eKgASlm11cwqN6vgCklDmuJ0vRl3NMilc6pjihu/WpXJdmbWkE5nAI0bcZA30G3kGROdpNC
L9kc+CYP2Nuz1y5DO8fnbM17+d1zO2yQVjBbe9iD6bfNF3WcMji3vXRoFnlPlv+hs0e+ak8uk2SM
EqUHhtqDNF1Ia+VXNy8Nurv9KQ3pSEVqVd0PKqVd7Ojh7wv1hKUNBYSLqEKZAN9XSRqUKHpgu2L3
StaDaOpV8En/8pFdmAj6ZzZ1gths3z0OfZRBz+gIVLUDIPksgL4PUHSKQPpJ9qcidA+hFGsGaogU
atTjuySUfpZw9XL0Vp6lAhZodVbMNzXuVL2V4mqsdF25Wi4ORwNLEWJ6nz4TTtrEsYUPA+5i4ba9
kaR5GSxAxDfxs5o6i/7lh9ujsr9taGqlrDrAOfJAZV6qU3Vxadtl1zVIEc3c5xj0rGwkNKrNLh53
2K7hbBZk0yCqCDpSxainDu5xYRtAQfexOnQg5bIV4zvbtsQE835QVORYNqfLoul3TJkrOFN/6edG
aXmxI1G3tLVGU9l6mBUAIYSB/arJHjfgHlnqKcfJg4269R4wFqEN3Ys8QWk4myGjoUuN7/xAYK2s
jD2ikKr7vJ0vZKPFKcRn+2bL0vNDQiN9iL+q2DIglconRzGO5nRE9FGiK9SPOCmfOhVhPNZ80KB8
sVhcn1I3nyZSGCXUgSauDBpWvNF/E0Aumm7+AQXfa5pmaJSsT+p1TAfpRWgka5S2heGGb17PNUcP
Cm8Qew8ke3Eux21iUjJgwIybYJg3xdsOtJKbWijctLbmK9MNFDF/o4SpNZdlfYB3fcf+icxgV2FA
FsKhSQKrE/K30wvU+2va2TnWVQC3z9ag39Fd8NsZu8IkZe1zJsfMf6I0JgjBWoa6a8uhVO61Y1Wk
7LdlC9wjrxsbrVCe2lZi6qfyustqs+WyXUW9V8+uA3X4OhY5FNQD0RpbvuSqGSvfod/AOT6wFJjY
mqGzsQiwP/6Bwa8ReFTfSl8D4j9nr3wYt5GBeT9mFPH8wSRiKC5BIONuV4F2dQTDyantNNwsqYr3
tKAccuAHAy5LAYM5AZvS19VFLQVtSjUtbKtzvI+agk5eHQ8ILxPw4yLUm8iTDoK3ap0/wLKBp7hB
FCMtSZ8Kknaj5GnwzoXJZ0SraRjktK3KIe1yRdoQJ4VAJchutsHkWWlKJOmawp8RxYCrp8Urz1rd
jf5KMZnLyXDQCfxJhJJtsnUFbvfPX6I7Wycz6AdhnTTy3SL/I2K7DVbB0wl82+43KH2ucFxA0qu4
dXTwWQekXyAyKJ+9QZ0wUMFWJ/iHUe1wsgVZ7liurjb/xy++T0YwUaJz25V3u+WAmqRWPpEFR0Ql
8BJToME34XA3/dVCO0lXQ8qI0IrELrJ71gltUVaOdEZMaH3i5DFKd+a8pPDE0gmOclvQaXARxl36
4NulCKXtz1i/YsdtSTn5cB8CGN9XgIIACax+ePfFTLR26ygSJvk+11n9j4VFhzdcpdf4ujnvhJIE
mLSctxCNzLCpakWqKEjJTPJN2pWWYiTxksxd3SRvShBcLRhjnplQB3HyEz0wsvTicLAKr9Gx1Wp3
nnX3W3cKyx/6ULgajY+d7ChFxlrupaitTW79HNq9wuHcjsZm1AiCzH8bUmW8AenAiQKNGaJnTkat
IRC1MF0gaOO09VIMJaFqxMDG2118mGnRKt0mSKxh80uT2w65o1CEqZFRdksUnAXwReabb5UfEoMh
xRKzpBL8NJmRbI08nxb85rZcVmZeX0+u2XfBtHKMAWL73xcHiIUWqkK+okwXQGL80l5cqkiBfqdY
T17CZ1N3StAKdmz/cAz0kadTtpN27yO10iW0Wb3lOlcgOGlSGU1VYIroF7sEOB90ZhU3Rne5eexL
SR+qLgzuUVgydqudrjgvW+GpTB9egPnU8v4cPZzpqnOwmohHZuRaELHbKwYPaWgJB9ksoKMvHbbI
FHpEAP/i3v2WeuJz8tcIo330SiVI7B6etx9oHEL+LP92hiiUvx3hcFlnPd2hw6UCuoeRgFsmc9Tw
HNKTw4qvPod8ngNJrY8zfN89bqBJy/VeEaMUk1zYHAOwdcrvfTPa2kO0hSJubhnvxZKva+qPKxOk
N1NnVZ1gYuDtNkcqZOhVgNb1e7w1rMC0z2G1s2g273VgI+pD+A6lEMnq50+oIs0oJD2G0tjVHgLU
pOmohXahk1jqljsP0L63EBy2Eawe/wh6BPdDoEqLH9tiVex5kCxRCHjc1LdiFOemsisTMygrU+Mm
gZ2iPj+5ykPf0OxtzdrJ7mY/NdOzw+oHrWegJA7I7FKrxBcXu3GI6w5xRYF2DSqQDTVv6E0xqzt+
xuRmpT0dgxQOfyQueK99/wxmbF2QU1x6/HXQnv67bT4G34QGD1qFPV0ghDu8PxS/n0PxQUVrHhra
kwbv7DozmOC9nGqoMuCzq5qCHQII5auprUkWYl/p8sANuzVDrDFA206IiB99xfLz5oXY05JNs4rX
ykUow6LNqxFKzPkTpApdOFi0dp/DX2HAiZ3HtUiFS18JSSaVqNHTfPFj0J0WZzndU6XJzuUl+Wq8
1MQNlhSNkGTMJIWBwJzCzS/qqfRsGvkbhmGxb01CZoeCGhBJjjQ7DmVku0ip5zgOxaVbYAVFBp/E
JXYy73yy3Wd7xDAv3m/XWlaciCgp2kWqVnay5kmuuNptErQ6gGL25d0KTI0QVrVh1XyCR2laEli3
eGzXcAgZeD4TEYrYF6+0OHByZMOqTxS09EH851jdH0/81awwZMUb02q9sgZ8+4viVXaq59Pl32ti
HuaJ39doTiA2CLhSdmBhdVhSyL+vNzW9YwYz9dgg0105kRBbgEDX1o6GFkwKqUeYRjOj72fnbWwk
Heqnko7MudKQmJ4cLzXg5DdVjyoWaLkrTZPIvq0yvzBMgg7MgFdtWdpptLx2koWEOjFTadQava/a
1pa7DSh6okcXfs9v2oD4YInjRe8UDfunHZaUtzKUYamK9QEwF7cMqhsGXHad5pS5HOWNHyuIHo63
t4SyJJlpEA92PIzhmR0WAmEe/09GsaGhqqMYaejmxYCX/x9mLsi30eVzzr44J8tlMmKGKXoWVkBz
Dju8+vCRYmjuhfuA5N2J/SxF/zRcewwgAU7P3hl7eUM2LQnB3uDxsP6U/hW2K+X6hm2aJOY4yfzk
XUxOboNmuA/nG8EiB9Q396UICs2v38pWMoqaGptUltUlMgMeFBTCO5pnPyUOdolp4guCkIRV8IKM
VW+EKRhHqgF4OQcPquSEWLl38hRsBvRremYBr9vpvqWB2Bqa1cLgfyySb8xBsOdQjFUlrWCgHRn9
QEbyt+/NqPZl84Xxl27qeRTtAblAFlkcFrBSGrapn9G6zxmdPQV3kuBIwKWkmC4ged0FD97mQ3Hz
yiK1Qge5wBRhkP4C0LwbzwCl7N2v4Svki0QIla1jvUIKLQ20LneTA3rvR2vWDih+hEQ3ppyVGHF0
ehYOrz6KI+HuywWSUNeQsNtMRlBgD6+x+vlN7uBJjBqgZ3hQI6E12QGCN06ybrYsj+R9hag1sxOK
1BMspkFpzAMYP8k6gOZuVF5XMqxPC8BGTJckFzZ/U2zrBkYYBd3TD2C4hHxiQpXwnmn+a1Vpjx61
bqoGVdmlRczatUOmfzeDV8VgKppcbMRfg1Q0q0odxLPO/TtutA+j4JpADMG38J5jNKHAMDNEfNkX
8/c5ip3/frzVTjj3GPXRKGAag1AZo7E4spEl6pQlQMjo82ze0Ltz2OqfURLPf5s3BcN92OMIc3W1
ZyOTWODyl0BstvmxLbF1JBsyne3oUQlbJ3oVjIb2sb9ep/n7gF0JrwFNbc4AVqGOfRg7GKd5tSjE
D4fXzp+TszDP3uf5YvaJc0/V3LdIJ52Vg72P5TL0eYRxvlYgfM5VfzNcRhP1SZjKw6kTSIdbEglm
z5GkdNlEb3S/G7lQC9QaEqE/bgeqbr+EounKBeBSNPNHvXqm9epHYQ6e3DwqNE4ORs9Wf0bs1qNY
MNCbpw2qk9GidyZY3GqyrQgxWIQVcK/59byi1bg68uFqZKrw3SDOvAEzDSw8I9seQZLv+uwHVETR
bijutW4SgMPoxds6FOQQTgHEbkN19GjNzrBPqtOL0qRG0J2I3vbcwVGBTedJ0JxYjxjwAccHVa1D
I/9FvYxAMrZVtxCKlAgjlZByU20RrMU5RNiYIlcxZOkQlx3HBmXmNWbSbX6TyvxUZQjv2m0em8Y9
AILWCNCWVjX/ckePXfmkznx8318AoCF6OAIwCEHRU32L2KHs6SpQO4rvzHlRSd+DClkJQw3yMKbT
yRLZCDTcDhY9b5InTJGKn4F5fNlk2JI3jFPrHuC/IebGNnOKRjSp2VRcfguI+Co5vQ3rOpeya9ho
iLYim40qBCuDrBFtN8WYl/bKWCXc/0HbmhmdMlI0K1KuQtIIEbBVRPr2Rnq0Nr9ZrwuFNCIJiIxi
d5a4qmp6eL8WosCBMuCUImRc0hwYXDUJ0a8zbS+gQim/l2HQ9LHP0ERPnXNrYfaJFvFG3ZuhJNiT
znyIVteTmP+tGQvciXeho3+SrRKzInB1QMwDs6eSjRz5L7hVCBCZj3jTX/FcTJFPcRlkwN21jQG4
viCB3GM3tvZQKFaj7CCrOFW+XPdLP+aMptHhs2NWI0AnOguVV2djnhcR/uv3T4OHKfZL6BvI4F6f
GoOD4ZNepFaMSifTrUaWW64f2JxzSuMYdyQqDik9TljGQf5VG4La0XhXG0ZMvvL9ejPbBWkO2NkQ
RDjG9qzC1ImDQv+z5cD4FCNwX3Lhnr0sD3xbb2j7PkuHHV24piN5QKQ0Ne9+RrceUURHpnJU/n5h
t9N/7GFZrdTiw2E2htlQWj0h5aw3IRT+U9+YJaAu+f8xq6D03PBSiCBgtm3pGbSg01o8FORM5XB6
OpW61QKBBHyL3Ec0DYWIV977WUP1gCP4yL7RXi8awXduOUcsw27ysozu5y4E3Af0bT5Rk6UscF69
T2YnsIwdlXSTrPqGJ8pfSw5phcEib5ErPNe0cjn1M9iRxVV5zk3SybZrfXDIFopdYstrT/Zvx59M
K0KbfpumSUPRGMOAhjGMfmCm5SAK5C4ZbHClCgmJajO+Pa40Co1HopmRUCbTWzez42j0Wn+aM53R
uzG2aWVJ2RQ7wGQwC3RTTn/CLXC/0w38yS5uG/IqrNomY+msyQpepHKxB6D2sUyGMXrAjOruL0MY
+lzXvvvehB+bISFFwsopwATzklt7zxDqhTMXrvyhS8Kp5Foiqa8aedrcXtNr8OGoVRYB592bUelY
t9vk4VGPcmQyDN4gMqK1wdHNMIJmhJgNnyjk1KWXPt0ug7gY3JND+A7H08nrpV4V6vbUxSGK2aDH
xv0ez1XPJokB8cj2lq1UIZ4IFFIztdurbDpmPTAC6iDFiMlMtJ1C/EzpyAGacDbE+uf2AU2N6Xj1
6fUNCBxLxMYNurAn3ME79m1i53up31ZTFzZJKJN9IXCSmsUTLtc7I5p6Z9JU2u/UJnS1FIrjKC0r
Q1MmfGSFQlVhtdp0N9VJNDlju+bQXn4dYRsvfiazilfpUTc5Ng+ZVyCExenfkxnjyCXqPNyR1skX
GtXWQ7Zq+4Zu+5LldLliLSGnnNbYRF3bXmCxXNH569GIG9rEyq66Zp3oI9p6YViVturTY107eibK
joMDmlXMEwW9grm7qD8w0GMD/XajX/57U3QLfk96ickbBnbyPp7ife7W+gt9wVzfceCkRE1L1j5q
D7oOPGK32Kq6tKlX0DXPF/oc2+gXqbc6HYrzwFcdzIXj9Oq6TWthu/KMC1Yc1QUtWdsyMiK2AAlP
HHmK+60KIQo/phGABtFAl6g8BfVpMugSsY6YYjAtif1FjRVkiiMB5PiRVSkHUeoCIyK2XQxTw8ZJ
54WEXtsUU1qerPzV0FCMIcxDFJ12J64qA91XVmBVhvqMoupPuEtm2Aih7yWwW6Jq/mL++EIsF5bC
Tn9WT1Dzq80fqizsc/mLyW2VZ8fctGV0Z6QcpMDhsPMMR1Sj+BTE40p10rVR9uSLHjE0d40zx8gA
novcqrJtnB+cg/ExJW0vMJEs8PsFPfNV/imsz+u5qBqjutZbQ2y0qLJzk+FJ9Ngh8l/tec36pq6T
GI0xkRRtYZHFHKfn0INlEA1tFV6IahZ8csCYU8tVdpB4zGfr6/0OcOSl68mroN6tYbD+LMrFD7VU
SNNAjxxv9P7Ryqvfhk6ZDYFoZh/ocbKwL1OZVyQ1ZHpfBJtPUWj1jD/lRab7HEUXdDP3K8SLFH6T
vlT5wY6YR8hK7dXIgeuYTKc8TFp1Q9803uZltY55NcOXPcU26NRUzIQ52Fb53TJPyduhqCvtyR5A
HZ31Js417gcqXy76CebgPqk8VWbNb5A5JtZGyLqxRJDs2YqyGnwPujAJJUL2szjELTSXxucqfj4a
0RT55lbI6TKLtuPBK1+4LnCxnO5LYsemXxBm5MduvYo6kUCG1qpSLzIEXEPx8akB8WEiea37JkMl
O0Q6VPgAoa6MtT1tFvRFhf/R52yYJPJEBc5ZKSft7g5Ihjm3qLHZblgFFARoP0ZwdO9xP+/PpJ3x
JFftQLMWUCK2X/DiUbsq3Lnj535qSZVyHV2XNFisTtCq9J5PNRtxQZIyOmCKqAXMPWSBMCLlbd6p
C8Kjxare1GtpMxxCh3GDQ/Rj+os4rPwJxhJHr02mW3goNt2FoXH1t8+wDPJKqpR8uxefY0gSDUMr
KPuUI9hYSsm/XNLloLkdxjXaXDnzwS7gejIFmmZ3DHI25y4B9JOnzGZZmoU8PBhb7kZ34O5slK14
JjiLWpPPfvQ+Nx1NpX4dnwkzEnISbBeMqwAE3rR5iNo15jC5DBUd9kN2BnTAddgzSNYwvRmunMjm
RQ320uR+BP3rUSVhMbNbFe4FdNb1MeBHYDsVe2z7kEWQL3gm5NaDe5vDajszo2D/RLcGK8HO2Vsp
XQ+TMdIXPGWdeYHYOEizPGA8U/t1QFXOgZJWG3zBSC5tD9agcthfij67Wse3wP+cIm0INbJby0LE
vTaCPkgg92Ik5ggrgzFCOXjbbhlquQROHOvvsklZKj5jON8iJUWuoolO2ihxKR9lZgeTa7ySC/df
GdLF+vTS/ALSQoxkI68UA6/IMVEnGoM9wSlrqqqR0r6KE6jqynS3nPUcSS065PpKQdj01LpYViGI
LqX2xc8Zy3iU8QBKsXYyYemuiZzkjQe+GwrMKQ7HWABDfkWSj348iVTTsKsz6ycLifsiJ1nz/0Kd
3s8LqH8YjkBpUeGdb1awYhFZbnBPiuwD63byXSUt3X2TPD9eGCNesmSssKDD9e7LV4IRnnLkKshF
jzKdfBXLxuZxwQZhx37O16ZCvsttn8H1KWvCWGxBD3ap3vGu66t0fgYM6h9301aTd54rV971PKRe
jkJSNAQOpIoM3yZ3X6HLvR0ihJM97JoShB8RDwp3ngqRgFl6tpU3ar/WQLZAeug2/ZBDf101aTn3
1v+XQyVlLylTBACpgEb/yRE4m2qufpRFpyHbl3soFOgnaKfAsvVOuGAZX0SnQXLQJHoBk92lobsy
ezDYkEzP69uSNd12MkZQGl6w8ZzqWEM+d954HQdWd3NlhTa3j+2lZ1orOupeTPsF1htddOl+zREV
vMaCx41e2VEC7LtkAADX8to3sgVfCFcJSLRwJTIdMS6NFRaZWOzY8bh2bElxNVxwG06G/5m0tyC/
9A2+s9waMm5JnBZztTQbejM91XM0izrwozT3vcg55EALNsxvqf7n/SCKclQ2xRbeaDCcwkNqanjZ
oCEP8Al0TVAfbgqlUlyZvNRYz4cuND4aMld/qFOiMqq0lZ0NtJRUdkswb0TDTcEcAcXRToioSg/k
hD4HT6O1ZCtLJLu02ZMD8k9S7EWxqeKWveKTE35rQIQWCfqn74uMH1SOLJ0+nDMsUKoOCoPFGXxP
Q4hYwWqF5nfIgy2NFN/mv94tPCJZF7pKYm/AIF14ZwVoBZ3jNPgaKDwWSWHP91xjtFjvDc3E2FZF
PREcpoEcASw1tsjBeEj6aaL53ibseDPWaGH4cKSc+XUn8VDmeFMG7r9M1puwF4v5CJ+00pohufL5
NJZLFyZp3RmbdC+8LTCgkLRxjOOprekwdSHTfN1fh+JhoLT6KkStzaWAjkkXYrQE+Zi1x6+TuuCu
0EIY2F5PBP9OsBuOfG/R1AbZ1i/nK2ZCyJWTUrHjKjDkL9qgl2rVPdrUNmVZ6QrcttRNT/k8eP1M
7PEdsZWZEBw3ZHs6zX9Gzs0l+VmZGXRPa6sI8kr16bfizt1awYRf5H7RPnVLltbjxNEsBQ3L+ucb
yODCvmkxAUjjOfhEI+d3pTbq41TYRF8vHECfo1zuSuxFzv6UnGj0xVr059SljEwuXg3BArFJaCrG
RSioPlBXXO+RFOaE2XIiUcjGV8KGAoyx5t1SUn6HqjofmcyEfCElNVitgY1A42SMzOekKbUuQJPy
87nlYfyY143B56wkTUmAHA1bGnYxCsCbrRKmjBwJbCtEBYT3v+2XD9yuZY9sMXCZFK41EzJREhZ/
6UjIDKbe+9wpX4gc3GUoc8A0UrejfXEjFyj50UA1xm1FR9o6q/90EChrAYN2CEQI8wulQmrJURRY
UvOKHhjtUBIvBeLmCTq0580U4yWNg69FzzKfdOGP+p0d4TSEJ2DEhYWQgFOfgARZdtKppe8JWYOU
M72oCgZQsZq5xzPJ1ANwyynfceCJ2lX+Qp9Mqa5yOmMkEr61JhUklPm33T6FC7BsiNfKg2jz9rnX
DKTnLqs/hMuzrOxO4XfN/3LdxL63bPqwQ/BX70+XZG7hH46/atODr4LifnLZlkC2Uej1BMo+KsIl
UOfOP01PFtjiqQ0cBiKAq15n5yWZlZxEG4l9Qo40C0rjpRiq2uGeKtMGnp27e7FhQcr/NAgIvaR1
uETBnmA0cPKvxxuXLJQ73D24hrTc2x9BI6dTd3VPNXF48rDzkj5QuMaVYhRdyMxmhlwXqqjP4YaF
UA8QGlSHjAWFoONdzs/0Zi8J/qPa/NL8SZGfaYoH9AMtSnxSqjQcNzjGTkI9boDpYOv1TTZwbPsh
sWM6dTjTkdUkXcOqJCkyp+n8yFSwZItg0p/Ofr2/B/shfuq2Te2uLI9u/1ulGjsUMOyrkLa/6V9G
4vrU6chX13bHAWtvzT0EXWyH7xQfGX2ggkyWXZTI72eBstFcjrBJlKYtXrFgpMqJkP56ZXAU1zbn
bkbIJXBFZBwutAunv9FwN+IVlB4LZV9ZHwP2yrNm/lmUHmSNs4yIklxFeDyKGp5qSvN511jLfbPN
BbYX4ehKxIT+U6Rc6kE6KyOrTP4uIKs/JPAKyUW/01QUuACFEvxl74gRGy8sFTEAAfsENzke9qKg
/SBlp8PI3fkw3MclquNkeFj/AEZhqAzup3YFd+yW3IZT1w/i/h4pF0+Bzxi48PPa5LaDVU6GL1xx
+oikoJLhsEwiSZfQe4Yl6DrCCeAxqB1MkEKaO7Attkmo9X0NEeKHjj3sA5V/HyI56pQ+T1Gl4MXw
/W9BSFs5Q94K2N7ngBUJtXwJSb0XquEj8i1ILND+jcvXpSZXNBYsDRHiZaS9hXKMz0yHy3w7w8mI
QbDEc6ugG6RpNGB+Jmoh4TpgNw4U+ysBwu8nAx0rg2DXnS+IuF/D3p3PbtYph9FjFmGc2ndo4oqB
6cDPpSkEnW3Ak6EIpkB/OMOaPl0mEec7ZPbG4sKkmbsy0+KJ70eA5KP29eSIYcTphs62NlZtlpgO
L3+oOEPKmFOCGiRIxV3JWLdsdXFlnu+nMNC0vLKWAo00aB5CGFubv5PmZEgHQhI0UQxBUvmIZKTg
WOTYiMGLu6raaLTFBiDzmeUXuYe+4MkJlH8IizLdFmCWy2ig4DAnQHsLg1YBNRd892iRxXDEJY/R
m3VCqblO/xyULN6AlQtb1uVde2aSHe3UdC87lZBlsUFlab9cRpBDFZYK6Iaf5KEe6DftM/vW6T8q
vLOGpEg/56vfZxf0GnP6oJVUzs4MexAPl5kOJdNPhd5xOV3Xz1eSJbnJhlVBXOZv+LEk5V51Hshf
gdGn7SVPrb6M5aymMwVY3beUzc/8o+wlBigvasFbuj6jX1wtBywMRFb5/ZnE3x0/okZr4Iu4aD4+
Rotbz0vxAJf4KaNxJuCXOf4iySc9XoBjWlgCG2Tw0lKmEuI7YEULFP5zqvqaAvn0MKhJs5H3DMeL
tpmG2aVgnhEQLSUNAR3cD4h5bk7nzyogCE/EzC/6b9E7PjqgA8TOZm1K/fssxvfi9upC7KSlBJEB
R/KlVbu0oViQYTizZ/rsWSuTzMwadtDtvuFR9mqcnY1pq6J/Z2sj/9wFzMbk4u7ALMeOYO4lwfyD
NfduAchx731JSlAB8HyV/G7YoGpGBdn/wJja2FUkb8/chuusIMHjHOx2yKZQx8SGun0VKB7nRYIO
chO+63FBrKqisryEfmMBk/05vtWGAHiMpCORLFhNXpMm5SlswpSSBtltrOU4EheIqwjVFWwoZr8d
/mmyN2lU+tMDCc6zUxSuBrwiQYnQ6v/iILihG4U4bRxZJa8xaET+clVauICdc8hdBdh65iA8C41W
S6RTDge9qwQgSAfCifjMkbOAFxhfdzUHwXq6sD24S7AguUMAw9k78niUcrieJVCYmmJZoySv4kW/
2pqwy0RPStf4JCsXV5vKWuxdLMGk1K82zg5U0091TrimRlVaTGR9FxyJxVX9tSc4pPAN1rNJn/3s
vISpIpKVfIPYCUjKgU20QuYSzir1GnYua5tweTXYZQjpdwj/0Z7MhL/jdVlnD+OvxKS/QNJhkeEm
7s9Ko9Kp8Z00v6/41HeXL871dawtdhAKeAf3EKGi+HxnPdJuDRjYF8Kk3L8FYHGNb9PqdpLisBX/
uzWedn8SWf989EGss9WFqZaG18E7eHiH9tVQnhr3A22auFxKqXZ3xMFUCCp59KZ9WG7j4nkBCWJR
UkQFGAW3sSOUtI6tZOQO50LnJOC+5D5xBfZF6n4ThWZzTSFX4B4PEx6nW6EeSjzADqis8WRhoH3S
OHymvgENpeGu1R58MNWg0R9YTLUGA6czH8iffhpb6wKTfuHn7MSZxBoZZQI4HVBVzQbJlSCHRAHM
24kWz0p2mWQ4kHY/v31JhEUtXhx2qqIHOUOdB9EbJ3nxBZBxWPBEd6OcU2vBJ9WQbUQWhkJ5eBG/
Uyo+5nwrGiBxGJLX+A5QjtQ3nidIl7XTuQwhTCTpAM2KVV1CokG32v9xPpjNut+aqxxVJYgFCoAR
Ix9vnvG4x0qAWMdlbS8BWXri4FOaW+kc3jjnq6ltNPvqAaxhvmXQ0eAtsn8C7pifOVW7lZFMkP+C
lLbx7Glm7TomJFV06f4oIyFW3xAj3fuHxJ8CnCXFQtijn7MsGF6VyQe9BN5taH2YoPHh7pFUVZ09
Az0H+A6I2HfuW1PQDL3acKpIf0aFgRpprB1a43HW4jFFy9FRvA9PjCvgmeZj2+9xPOa00pgJc8iQ
yWiZ351uMY3MIEwUImIHfn9vzSjCLNum/hr8WgL3htBgc/a9cQwoW/ZVjr0kXJrtYQQCcs/zwMVd
buM/RIj03RRZ6CDhU7S/U8rvnNyjHMTsOXuk0UPTzxZEbYuvW0yFOIodIrvSmyGgtJ74cb93BJja
DiQvfogZOhrh5miKV/zvCE7bNCZ6iKMN+K38a9m0986AZOzcNvSNne66Y14DQ5BkkBkiqfw8PJqr
mSiTPR2WGXXjHFIgEyHtuTonXpYrFo/N7or3HYvbgbdU9ZtpfbOfa69TqmzdFPYJHzjYqXG3MkUm
hFwZhdbzkDbVEaYR/xDkJg5hmPD+EoMRATg1DoYgAe43YBuajPPItXFcwS6Xq2XbrqcXYrGFOHXz
NAX+ygwCqQnHKqN6YeW82/3VbYK4e8KKwAdXKgxPuVhybau9PexGTDgKPrJgjHE1mqpRgLu+d+lv
OjaSIgf32fxtGi6pcWHX1qZjK9yCFUOs3lHKUL5fXWOJB3UEC64to+4E2SC3vkRR+NfHqOtaGV6s
+YEmkZOTPBz2uLUvZlo9rrsOWj/c2wN1AGjWME7kqrujIJtgDhXsCXo7sRkO4cO7I1nyVNXyHTy/
B9tf4f3yo5prW42uLIeTpjaoVbW78+4eXXYqjvrqJV6DWv1qm62MeBQ72OQNvsLlRCrv7CdI6gYN
7lS5ygkmxrKZXea8bqziy6b3XV11K06G8e7TVeNuJ4zcshSeFDHQCvZ+boa0peNtBuTQxuWBAcAY
iW1s43V7IXi31ljdpiFLKLEZRFWHUc8XJY3W8AjJn6Z3x2BX0W3LSP29R8quLFd1LKtfrEedB3H2
tP6LsTncTOVeIOMPpkEgP3itg+WPpz7vvXp+dmFCg+wHHrQaQB6oTf/wyzxSIMap/97QqkR1Xzwk
L0fHLLOL4Uw5w5/rf9nRn+aBrD8Rtpssycj/BdJqBK6PahvVvdyL75GUl5140MJfSLOK+eoZg56m
plkEl2cuoHWNxBIuK0BCjvP73X/2z9iEWgmubIxwmheFATLLo5Kp7Ku3krWAE5Zn7IeC4jFwlthD
S+2FWd3OJZbUPgcKRUtwCzpzKODHCcbUN1uyE9OBZ5w4ulyFcuFAKst8VZ9pppFfq0KsVxoKsfmK
MGIIWLWz86IOJKtJuDpVT04F9QYme0vRBGZkbRxHDr41GAVHdTS3FaWS/6sUc2ikY1W5b88e0Z0C
1iAZN1dGwQCN3D3zIh3NxvAvwb1AdLBElW854lCftCj7qftcgDdfvSeogNjRc9ExyPgNLyl4kj3C
Oni7ce7RHhzRqueRYSdeeL5wqvt633rwysJ6VS0gHNz0JPvSku9qjNgmXKyQql5+V2842GUmya0P
JtHVDCHxus54r4pUxujz0ae6lB/tXFODY4upJGWNpJA7B8t20YLf0RteAVJKJdWSxCBcOM9kdP+4
86u09nUbAdSLRmspjr+bChEP2SfHG/iXI1h75NddZR/c5otCuIhJWwK+uNXk0FFyTd48YMzeqUbp
mejjalveOv5tkbX1Oqcx+WkHE7ZYZwUG6gaOmu8OVHiULIv1Ihk3x4rb3uYvR3EYgsaV53sf9q2e
ueAS8TiL0pGVhgNTG0E26uYOU43eNXLvY3kWQ9z/x90k7ppYLtjVkw5SzzUHi8qcuHOAFgyZbU6P
J0ubdJiUlseDa+BBmRrkfze4S8QIhGW8C7l7/ITBUZTLvJgbD/zF83YxasN2ceBA5/dbmu3kjoJW
iyKqmmyeq7fslvsyFyNL9kpkt/R5E0gESX0N774T7wK2awm3wSMM5I4lK960s/JxehJVtFmh1NkH
nZMjZjUh/q/ozsrbNStXMAt5hEwR8VnBzVPv3Sz3Xma8ar6oJy8LBgY8N3oQHOtNPQLsTXXHP7Cc
cUunzSFWi++2K6uCaI9VXyT82qIwwTuIBAF1cWIDZsxHCkkntYmZk/TH5YMO/dD0z13BZCTWjjg0
jIi3Ag1vyengfrcZucu9Zr1BmClpVUYKhr0E1sb8YRehLz5tlv5E/FN+VvI3Af/CoE3dXY5n5QSD
b/Eg6vR3+MZD/l+a6WP9fJhk60NG9QiFgeAqZoTblOkUWzceGE3Oy5Hz0zUjOjiM4Uz6F2utvVc3
UBzo6hYZT+PmfgHETbnRRA0ifpgfBu+aLX2wFkswL2/5XzW7Upzuw2QzZnW8Hu59ByQp4nupIy+E
czUGtKcSg8DiaBVBIH6LYzdbCwg/WOSB1JoLHLsXwydA8cTFi5+f47HMH68Wpe3FnAWv0jFtQZyN
ijyt5G0aGMc+LI7tkqn2l1Sfr90407pCQFE6moDrneMIw+M7xdEtLyfzEFm95gth96uWjIMWp0Eh
lz1XDM4kydBPBkA2os0KB4iJtHnyt4eqdAxA9RXGvuPLSjQe8zK3GqDwyUu5zlv106ml7912Ug4z
kMXOZIL48M8rrNveqBAyNwYMdYXy/etetxuT+xkExO7aTJ1RpEVfIExPnIfzp+XJ+FXP0nW1sUx1
IfjyzE7PIF5voNepzQhJtzc/mVkw0eZjLOEt5g97X1FPPRmJqdyCiJzlCYEEUOhqkIvy3OTc6MOg
/llRCJwozn6wjcUsc1uToIgfnKpmgf8GeD7o2Us+Npe2QRWTyJsi2aT8Dz/mO7lf5SJztofLEAc/
HdEpo/VXwbRvrTp89f6K764g/J4wt/Jzmiu6JOJlTmpGG/4PmjE+wQaOWOh4Xpw9kUIsmTDJMHJe
eH3CqHzo0kaTzdaR5uYCUE2vbZxFSw51UBVjZDh7DCwM68CxsZYuVam7fxXPWxivSWm2alnPIdi1
mhG0gtxzMO425pX8uYoifCoYJMuWv9fcOYZQzMPScv7dMapwosMXz1aEjpup3mXd8rurAqe5S9mJ
P7foWuxn6yCvNq8/GOaexqN6qPNdEvppaoTQ/MHn0102nNUCi/obuRcqcNfr4ABglcGfpDydKwOs
vnPAmEo9wP1ytSzR7rkBg5O3zmv2alhaVZimKqb7u88YU2Asu/o8hfgZazRTzdjJCu8eQl5FS9SF
/saz1yOTGiQazJb/aQ7CfrOvyqjT6yX4/928y5MDQReTd9ouJ+gIkUyHvvAbymwknEluuc7vfdOP
WVjM/NJJ+W4AMUtt7UOq7sJ+fh1jo8zlpE11+Zr4kEWn+HtNiF0Nwmws/VVyFXo0URCnCOP1NRSH
c+wiohuMvOb28Z8WUE8578IDF+dBeWOaQC/9t2uMfto7NIzBHRIaqj6HX8wi+d0Myp+TGSAWLKBd
3PZ93KKGfXHiORgecERJc1ZDAaqjs0zIPEk6nKh2i4byauCRKrYlrUYdzjO5Kw1kNA0isRl07Xou
+8o6ZgfKJDb86V3mxg2NX5j66FD3DRJlJSBPWzde0V1a86Oir0PxfDoY2lyNbVGcvmIs1pq0BLlA
b//o5r60UV26i5GMnEFBSNugS3ed6UsBh/K+VxPEaO9a0Zgsr0PQ+GTdR7+H+1PdW2iquBRg6+QA
OVBGdKbfmqe08mUHw0kO3vaP+PzUA/Ci5ihLW/YDP/HAbyeMEhxOvcQfYLILeIfRV/HNpDhQsZiU
0JnzIJVzFUeVWmbX4Yu3WGK28XoRJLtmgg9eZ9ala6sBlv5l1W1cA0TWzQ+ttimkGmymA71R57rj
6Z+8H3aC/Hsqd+jcQwVmn9+p+VKl97fn2shX7HLLLmxIzt1drgxD96tqUscuX4B2I674KJpw+Dox
KJhEsNklEWWk0MrI2M6qdv4har/YkrkRirjicL/sOMuPzP2OBLzHXDFU37iuOD0ZxtmfQLFTuGd/
5i94M8OlKp440OlDEzb9CtWE79wBhGeVNDdiHVhaveyLS/SC9yx3Nl9EyZZuEqk1yB1o45ZgA1vS
AphSDkTB240iH1HzF6qRJnQCeqZ5t8sgL5BopsBLt8rB/6AB1+ExfcWOVdpnZUOryVlZessVmZYo
C9JuvsRfzwiB9NbdkEGFzCUaORSrupIrSUDvCQeObXCa53rkxdh5hmd76vlJ134zzEyRBHr1szM0
mBRlRTjj0dpcvc07jigLjkd1f0qWj4LPHmciOKKNlQcT8gyIY2zzVnLLY1TcO/5MsXDVTN3aZ1Wm
Le8F6N2tnUxDR6mcpgSwnh+TgxJ/rd11zVOWYPqKLT0a2qU+163DE7gXO3FWjVT4yk91CGkNED0M
uhaRmYlsXsV0lMb3tRlhXL/7II0lhtwLfapPoTycEK181+zzMw3s8WX6KV8r5j3oLhKGmZu1Y/vH
oXAN9n/an+6MB8S39YS7qe7ubbSnEWJuZ2b/V2jDbwB340tHHepXxlolkzlpQlh/GntYmYmVt22/
sRpwtygvvpK8ikENqidrFQXAWq0RigclfIyG1U+MD1NM6r8KTRU8WcghAkNE13lHfK4f6I1DiroG
jlF6ykVTdJ2mgwHka5skHfGE3iMb4ydYiU+Xej8y8yif8v3/XbMXmOFvCumgRv4Pu+rwSu5jil6q
Y8Qb6/Jj23H8woWQOsT2tmsp5DozmG4vlDs+vTlho6JsDasJUqt3v71qVgj/VAfL/3I2V+43SjTQ
etcDSb2UAe8hM5NGp+AsPUMoOUHQTac8ZnOd+f60dhZ8nok4XEQ+/wmYZHdTZXVm7pqzLI7/jSiP
Ap120Vq7hklOG/aimyqH18l57ycjp1mTLON58AjnA8k+Xq+FKzfSGGYLCSYlWBLqc2V09XD4IYxx
OCGp2XkJAiMg+rgJUy6xwkU7J43EunmzARrDOwpzkEfFgYJ+qcTauRc6u6ZxVI+JOWzUavSuHHfA
z53q1+LADcLLOciYf6SI5STO1P6JY/cYCGae5SPYtYjuDx/MAU09WMMoW28MbwqtbAetOSchZjt2
wUbGA0ETVJfo7h3dyI/JzsaXSm+IemultpUYOYCvOyt3qxzczYxgxteii+R3kQOZ1Vg9pGYnbW/X
DgoymUoGif7CPSYej1AdMr4+OaP2DO9H4Jh761u7JdP1Iqk13+L76Un5snjFej0gzqA2sdbhWJTq
Y/7DvLhtC7wAqk4hCHwUjJY/ci0yVUweYLs4tQOjrrtFRHHLfkH6Ll0WayS3I0yqF4AsAx5ygZBL
dZuhHJCvLKpU8Xi9JCQnmjZkyj/zd+q9Ukc6t+kFhLLelIH7dLC1RRBa5Lo8J8HKjbkjuf1MjclI
5GRF3dfAXtdaJA68Mk1daMcGMklugEwK6WSaGzBHsicJzDtYRsqNCvUCGDexUOJ+0HsF7GQXuG+y
6D2JMc3wTyhmP4OWVz0/ZD97qdDxXYzFUWxo+KervPbpKbhNpXbwYb9aFB57UMI8fQycs0Cd90I9
7wU0RkmaXd++nsQ0DuNWu/7LPjsA7/in3tqE6DhPGlWwCYMXjg2fZSfY8/kAztHlYpX19ph7hlvs
ENpxxVsQLSmf0leuiB0ISJoiqmPOflbsE7U+JktyJwYgxVdBCgtBMk/xwUSjWldZsuCF2mQOh6LR
l4/d37fHD1eLchjX0r0zGP7qVmUcWS0FM6wgTchkfhK64KUadTOCJd5OCK5uB1GsX0s+w8MBqReU
2v/fa4vUBVlsBZP9IgkHNjjyvuCBTE8bASWtJnIkLnA7UTPAp65PqY7j6vSdsFYz4OBkA6BolHiF
uDfgVZ6v+oIcJTwoZZhVLC0k1lfOz26CO4sv0AzbLovCKhDON0Mwz1VkezJzNR6nEPE8UbCZyZCY
g4jUYsU/BsfUfJuEQqKNuLeMp9GC+wJFANz+MWvtxl8mPg13LruxEdCNYGha8aM/SI5QnFZ9OEf7
SH+WGCuqa3/xQsNYaBDDyj0HKpJqeKxJ5BqjHMjt6HapJFCI3LzVoA58wNl8ulQjPEEJcDj5Jq81
3c/g5OVFKPtnswnUcuYLgR8VhIkzosi6EdqnmsOfATCBkKyJLEUB5tnkOm8a3KQ2g8SWRwDwcC7d
jEHR83E5bhq7FFvzOnoOD8LDynOOeoeYySvsSeaJS4zqRU4JA+SfOR68YgzdwPjyG9Txtn2hEayb
P76q04RtK6rQNcLzf72GPkNxQC5DuclgVHmiC8rYKA52zKXyayWNvVqv4MZaFZRsb756vT5iYL8c
P8GLpUX3i/dJvQ5J7dGzOvGdwxTHF9QlPm10FlkUJbpo2gKbu1S8YAk86asYqnKDdZ47JlIF57vK
RDbG9a4ruB5OBGk1j8rDycvhR6PfvVQJi2QqYGMHthangLoUHsKVM9NZwy0zxm8wprOCP4j36cdl
iudU/QONabQk6DQE7ckhFJSne6+l9vV9vgE2OrzBAdI3JYp/mOFca+kod7eAPxNVf1kykyk+QfsF
B4nqZXsT95on4Y653UAdPjw08iHeR34B4O0unI+ruO/7ee3UlJPjcFBqXIZyJ3RL0GLYDgd4OXH3
2aHIEOlfCmcgCUxl3D1+7eqrmOhMuiS9UHwebzCjmn2+3IyA5R0Mp8v45DaKhbL6UFzXZzgydgAD
0HwOCwWwaPXIRIeYEVApOWGLQk5LSLorxBRoRh69zAtQeVRszjec1HuXaNtCuLWUjWk0pfJ1134F
jVYmUgOavQ3gwr1CmmX1Uuw288bt4O6qun+WNQNey3sKvwDl8VM1eTHnXlQ4ESXOtDXca3COASAB
+951JHcv0Rbe82Hh8iFDu2rynl4lSUp09yKJZ9X/w3ojQ9Wyuzw8FSFluvhsRrH/PAYNyurfIOZ5
M7plE8y8x6c9jjl3f7RZBA1TeGUdg1WH1y5AgOnZyHkILgFjybNp57Dkcy1sP3b7Rwfl4zzjl9p1
Mg5069e4mDRkAXp0Ta7Gti4znYNZH9PiVugsSViCuhkgBjXcUhkl5SBz3S34z563GVTNO9NIgfpx
ci6xXnd0lA72IwwNbGdrhm1WYZnPayKkeURJOVt7RWKXwNW2sFaGXVovx4921eBfgE/6qNZ7xfdZ
uXnt+sYaZHzwOOoLjykwqD7rWb+aKYj5RVsfONzVJyZ62ChXmuECh/BFlQZksnzs+fJtXKISsy+m
NuqlyyBQ0oqjzi5fLpU2ZIGvyfq7IEzohWpAfzYLre7hz8ps+nLsbcUpVaNp/woraDKPaxHj52ZI
ZPSRjQvQVBFvOjAtSyyWGW9ZgNHajlNzelf+sprQpEzW0HAlOwREvsomyj88/GbkVgo9F0OlpI6X
Fv8TA/QThmR8Y+A85yu4nyvs9LQFnasNLun3trTFxOP5d+CCQiOC/DfqjWeuWBMB83PpEtgrRx82
WhFd/MwQxPvadsHw/OkdlinBgdvjVKEoyf3afdz/EHnRR8bVwI1FNk4VpYk0aVYj0RNRwuB09nNn
dxK2Y9n3UCGqfJtVj18t/yc1zUgfBZvs6BVvOBZZUcRX0tMJdyn/MbcN1InjtgMFC6vLhwVDWzpN
Z5yJ0vzmJQ+u2lG95xxD2qg9cdUjj5bkpjmbiOriNiuV6azKm63GopHSnF45VqZxDumu2JG3Bq8X
SktX5Wm35GbHQN3+zFUyaGQvAUtSnzZZ91RIQICiLJyNnlLNu8a+ZUiAXq2b/XLemKmuv2tXRvvq
T/VFbHZberyuWxPDfBmnf/afpeokAuraY6jDQxxd+grK/R00LGocXxEqTxegH57fYPSxuKMvzh2O
M6U0qyalkEQEmvkt3daou6joLOR4Ob8PJdOPHspVFjGALsQ7B1aNu7Eev/vMKpUpT8P53vJRRdZ3
c82SRl/FlFaqjphVjSFVWNcx3S5lkxlKZYFpL85pNsdQv9YW1USaCJhP1w1escklgdRGV4rdlaLt
erBECVtK7138BwZiTzPIYBDooxx6JPiTTNQG+B1Uj4zOPhbkL75v37DEt+fKq8uSbVr4b3GuOvAF
XuRyPSbq33YzyQQXaigmh9zVEQ5XRLBti1YZCQzV37gEeR3tVCsZAUkzbdkWP8syzMYqCpVYDY5N
iWmoNXtNxq6aMJMkrMGhBADkmE+0a+opSQ2u49qkJFvYzbJBbsJIwSxI0MaX8MR+hFX2R20GatrY
QWuN8ms+Usi6UZkmqQHdGcgR9YNmn3dI1GUgvAsxh3snqHT5VvgTq0D299k3oLnnvFR9nMImOiEY
QgbTY90natSgMwCjVDZVo/qrdwTOGB/0CiueQ0+ANa72YwqHFuum6EdUfqdRgjNzMA8n8lNWdbSr
YHVBJGpRFcbDuWGrEo1dC/t9sdO0HZmkLHFAcxOr0tI13lkTvj+23h02Ex74tzF5Ht98y6MrouXW
Q0v0544xjy/k3ntsa81WtXdGNZfzBwjdq83SRPUxY+/g+tD4gzR3WEGgVulXpC7qaWBKhwbE1trP
zqjC8jALI/BA5VCTJYF/PsfsAjIKndiaLSvyrNdBbZjbRzl+ZIplBYMyiId6nFK4+SquP/PjmPCN
CbAd4PDPpUp+BiHiwHlJnIQGnFzBqwhCiDgFLCGst+IAqsqMQVv1MSCcmLsHtOmIpj/eleI7ZAvl
zuSptyuMe8Ee+Pn24E6p5Jp33MBj5AfnrJE4yJD40kGLGnmoch3nFx5KGkOIEbH8ZFkfj25leLZP
HOtFuX6K/EyqcyH5P3eS69YbtTASiG6wY6vckx0j/NV1uAuu9SJu4Ei+kQDBm+0SNbqxtVfpqcsx
K1UfxCKnt2B7B4H5Hhn+s+cjryDgC2YIrc2/n4nE7i5ZaeFexe3/dgh9GuNyRfdvxM8V0kG19hS2
c6i1LaQDOrG6DhuM+B9WYpDIQmKFZjyGge3cH3MNZC7og7oue4ikpZGvpMlOumjeLglZKbUnmL4r
wujuMLIqtyUXgu0DoM8bsdZwpIvXeQ4Pjugc6DeFyROi+V8WqQajCSUnFpyvMfAcCvuoeWo+zNS4
yglPWhny946B/nhrOOFYejE8XvQlgMmQfHX6OITJUCv25ySgH2ePssK5bfMN+DjSZnjO7SG1AYwf
+oAPE/IJXfF3u4T9PIXrtr+F4WehvNa4oe4JRvv0kTjG5kxS/bGs5MKbI8ktz6DqFaM2452MlBqB
SI9XRhJW5VC3lLUQTgt5CqPs+FogxjXcjP8gO/H54fKYpqdALnA8ffv3SE6myYGqlrvPlKXn1R41
sAWeitC+dSv1EDj0QmmO4Msoe2VG6nTnlwnzr7+y+70l6F8KIcQVU4+om3QAdsfC4dj8auOy/xLn
Qyfx50umCIgMh1TgljP5s6BHHOYv7P6oZrHG+OFKZipgCA320MYe/edFPd2qwHTjFhUrZ9J7Smok
uccqRPAwjJpk/igiuHKRWvLs1u/ZxLUE0jsBkih3UX5KNNQYllQYHW84+BuaF4RdLqmcis2JjK8c
C2PLuZzdiRB5LNqgNtl8T90+lCbyYKwxwWCeiHMMZlCW1ANrPzrpAbSukqJriaym52WyhD5Sa+Tj
Ha06Q0Chk0q81LnkfWfi4m8Z6xXds5yarfXFfo24zzMPXggnfYmLskjrhlGzxPDQM1oy/8fs27Pz
sbLCWPpmYPhmeYoyL+vazUPt+OpIYD3KVuwhdS+0eBQlYESC3HBQyrGOnY1fxmcXSWw/usVBJMH+
7OzK6MrVm45jH5MOsV9YXoZtJGY3VtBdueAyWRLNMfE6bNgmaXCKgN2FwkwvbD2FVOOhnCr03s2h
S6Cm3poJZ5W9PaZRUNrzJ9SI2LcG4NigrGOHVtdLXo8Sv99FP7UQ1FLXhnZd4ZRiwWKDtVWaY4Bh
NRDHNYCHhY2WzjA/n22WqN077AMrJtM0djs8RKqAZRx79KOsv2b/G1TYcPi+XWWmam8RVqGziWXF
4UyYSETVuivJ+6F8zxu7xhvDvgWZaNSLMFbdumTUfEsNznaJiHLFdMVUKVByk6BXcaTvGb3jJA9Z
Sl9BGX55nSSSlBX2GBotqNG4Rh/e1ZswC24XjkTGgFLQv3kd0VyXD3g+37gYlgd3VG6TydRf5t79
iPKHvTbVhR1kFx4lUQIvzmivENU9e7PQeLqi2OfNweLmLEi4lfuXCW94pozihF1v36d2X2rIS+sp
fSG9VXTTIzsYVepnsRD+AreLrZPvt0xmWYQPeXjn+jwTzv09VgpdpE7TFt3vpRMwowEeRwMW2xcq
ffT5lDd7YRXSLwiIubhjDt5p8rizAQUwX7lukvOGoOYFfj1FyQCLv5nGWSNksQEeoVlykDNsW1Zo
FTIh2cyP47ikOeYeyzVXiMp3OSTyWrlfoC7Mg1V2vYayDLDzgMXcRCXW2mWElsW/gWz1l6wgic8y
oOA00Y0dQhpTbDFG7ILVvqcuJsKOmaM0h9ue7MPYfZ5iIaj+nWNeS8ZLBNk/LKzhJeLLBLS01wT+
Z17SsakBZhsZtJmRW1bC9SckKJ8UGqSbWk4knZjIOhcxSGSxzw0D5bEGzWdBhEGDqrHT1b0r6Uaa
ZmoVJxX/Y4cZifDKP4fotLLN1UBkH+yt0E/EJbuE6Eyn2o6uMtNjGvXyqldytAHBUTJLVSvz9JYh
CO1Q3AHHU2BFa01KWw+8QkneO2dcJ6BrJZk+Ayaf7AqP8QP7oSCotSD6vC4feAaOY65/WEKz6uX6
/8t5/kRUEGpprYqAIaMbqhlZumg/2rAoLF/JFFe+zL9xMgGx56seJL/B8N0VLNHGkhd/GvjB8kAt
9uGr6VvXH3pEeZlYurlTnEakXvVVP9QuyDnaJE4ryD5sawctUYZZAI13F8cgjWUiNGRjSzxrz0dc
cUgCWbG49QOYeAdq4FTltoib1MDkXnB/RayGqHinTSjBiB2aUW4CkNEqsjAlM75qVeCZV7F01Fkc
TwUvsTin3qAGO+kGXJ8IaztX8gDXJmsodlFqbQPOXAZrFYIU3aus7TqwrxLsYUxqkvpa2g4X3cKS
POrPIhuc/4Z5/tNgLfOKJGO91BrJWCTbc4wFgXDAXlRzkd2FmAnzhQDOttk0QlkNiNVyRQ3gVtyr
ynjKIKiHGa61JAk/z5YG70xlm8PDimWOKh8dg/iHS+akMPvjYvzJWd+Ql/Boaae4WNuznh+skwY5
/+kcLMPiLsC3gpMnF65DhnxygzFH0lWEv6SwJFsRoaWleFuOe40CbrUhSuZC15u1r3GhvRIJ16qQ
5K5j8+nd6Q5GqVSbRcr5mB2sAS9s91YTYc2PHtRN8FWkwF8PuJqnt9zL0YKvjcs5V3bQHktfvLYk
KvGbaWMWsfqdqa3fsXlWSTZb6S31E+iO5D0NZeH0KgzBFzer4MMIpDAtflv+dEmh7rarHHzCTft0
ycMHdYPjXyL9DzUQmEnmWux4NfR040uD0Uzx1n8N5V7NBd+3KZx35+wcpDN+f9y73Kcyeg7Rn4nG
pcWylLI49+qc6NgwDIqyGry0fVISaUaDBalPm0cHn8AQ/BuhbiRJoMUo8q5mtLXm6aXIfT2hbc7z
Luh/zQ+By9QN+TYTmxbjMzLQO3S7Yp5SbfuVcISkX/ujiBk+f71S7y3/Xx3ZCJQysqDkUTt7ngHu
/QdZamEJ5HDmAypkTSuWvRJXiBaDa3vGhwa9jMu+hv9cLKrwydfiPPtqFg44WovIZVyMQ9D8b9un
6tZ4BF+mCQ8h51njjRBYBAM4DyHh9rUQIu3W5KqjcVB3acg70aZ3nL2swfsIqRiQDeK24W8okBlk
y3XgFXC9dC3n67vMrUCCeup/9kYbt7YIhOqVfV9KoyWHcT7vSVFNdEPpIThn9imI/IhVzUYCTkwX
OeGz26zI5TRcV+OV7oIwUBAoYTKGkEBUYya+GNpD9Qf5AJgYHzaCux6KT8eK12yw1Z+xRQ3hSC3Y
G1jXwCrWpdz+AfOjp7/egf5Xayg+IR2tohjcyZh9ppHLeoPJyWiBvROleS5GOO5UxBKThj4RPkSZ
8boTgPpZ7XhX8bHDwA4dLida0tRGQ7rcoLrV9ClpTkG1g2bffbAJaTnGxhLA9T69CIiaXFuVjzLJ
d3URinbl+RXGY5u2/TSxXcp5BKZiNZo5udCEcBtZr3STKbDouu2e78q2aBojpW/zDrdnny+uzBSz
aOwFBcG2yY/nD3UMTguV0W/g5nEGiil2CHUXmwPAplHc1x82G8na+FAyckbl4H9RPlr9M957nj6F
QvdPz428SyUwKYs6MtY5KO458txWpzynOgny3KgBniqNU0/vGoHuXARfrdOqjtE8SnFp6vCu8u3f
hV4Xg/N+p3byg/qfhsWWn4JzbF8CwsqoYsdLTpPH315qlVDXMq9GF4s+O8OnHG2xucTIOaxlzKoz
RLsWYrDymgjLil0YvHFQcy8uLw8/wnNGpqxAOHQNra9VERilg+9mIpKhItyzezivoKVa/Z6w1ET3
AmJiCCUt1Htn9Rvpumkhrzqww2d8mPmfIZT0ZbDZtSRS7sOkishWTwR+2BLzD+xDEJK4CXN9qSx0
zg7vXB6Tw6Ck+UhPTBwliFckhUPd0Mk0KifFVRdnl+ApL/CerGKh0RLF+cTwA+6A9jl7TWspR8IF
Ylw24DVZSP35C1bBfdVzJJHG7qGn8hXNhBNpMalVzvDvXpGCMk3FEdbC9jn8O1Dgjcdq9pkQ2icP
FN1N3EZXMaJjamgLdAP7ii+PWbJiwjJgQ0GJ8gys5qxwCrVXf0iJBAleQhywTq73KjpLzI4Qu8ke
WhZAHeM1IQIHv7faeG95/qLNjV+wjnSsic4n/Cfeuaw3w/SIwkwALpXcA3cy0OLDMAUmuj/swQ8L
bqL4ai6jRihf8btn1QqKDQsYr7HuMluCUZN4/z63SpXchtEuEoXVThVmgimgVM4bfLxRka1HyFYU
xMNcSJLkKBQJJAtftjRFGgR2th8LJ3GOwlhpnvZrwlROhHIPnL2nSnXZ95btL1Q6l46y1jbLok3n
s73JI6wiyf9EDlyDjas+Tz6jbPeuYcRVFQ27LX5JkfPLWJ77oCRm0ySalzd0eLxGGULTTlLCowA5
dY62h3BOlwJnOqHips71d2cttlQ5/ar96D3sFE6lcpdNAG8gocpKkUfIhzNhPQvoCSTKbVm28K4T
xuS2SzDpFrzEcPDXC0fHE8QYz7FJg+Ysvg8XOLDnv1WoxEBOT8OQAPwJL0vzcZsz0bcIfmxO2ty9
yxleRG7y0hp/c0kDcKVArsY4DYy3AjXSo9KNaGw82jjg/aNB86TR0ys8dYURH4zvGxA6WTou0LmN
pCmtHOZm1pd5EdehTKnMQ2ZmL1GbGuKWqUFPtSEm68r3wd/9UzAOrFaILxwDwmQAl/mGvgvymRkF
05OSrI9H8vP7Ja7GuoyHvLkL0+7VwLQ+PjyN21T35LKZl3FiYfKJDTY2MreHEth+QQTsImRqsJ0e
svxEfX7tZS0sNA1nt72bQ3NWto8ss740tLR/PuO5I2vAQkOGKQ6PbniikbucMB1ox3Y+S67/Ryya
H43U9STJXXh9FD4Flm2Onj6YtfNdeaO3++Vb6vR3QYJlSjtTR+E+9OaMl2ipokX/h/B6VvYokh8H
FAWN7Evx9fR4aD45kI8hmJ7n5PXw5XlhzB17aPDin0cKLQLOASyr2lT5+flDOv/FSnLfea3QtsOG
nUrh+hcU4LnjOqm6rlByDtDXfkOlmLaD8dmvzSX3f0kYxXuJ7hvR5jeqNvdHnyO97x4hWrqziNnh
GxIjS6Z5zdYTcbc5kmDIialhOoHx5oHI6kJm3L6UL8seuZevqcLfsIOoJ1MxleX+hgExejNkJrGB
iR4kdzW9plc+dN7OEqgIHV6yxEOEi9oxlb6iqRCePy+IOXo3dKzIApwuKktIz9n/HGoWcNk1Rv60
zWPNHwXr8HgbkpW81mTwktJyUeKpHMurKCWh4WH4YjY1vEUnInlXmQLYH4vwadl8C2PaTNiMBVB1
2j1MxkNkr3+cPcuF5lVZ3yNA621FENebgia/lHR8YeTOuTrfMxg/s3xWmV8sIf+tGz2M9KgZIWx7
dRae9p/HwyindnwWvE+wxxH8cdVwzwixyuBqjYEnC0Z2G4c9ahs5TwQmjivsspyDeDhAdsMHtSWE
KMDjtNZ/F63Sw+ivGz6YcJBFfICpgYQTlapLUiYOXFsUHpel6okmod+DugWtiR9H9VkVqAoWG9tV
dXaV+tTgtZTeKABTNTzCfRLG/Gd0zzY8tGristU0Qb/cr7sZ9kQLx+J7To7cbdF3QAvT7RmItCz3
OsVPQnZx7rZyoVxfAVJUQOOf/lHEyOg/jwWGYK6VamzAE4E4b6hzYRbEJRRbkhu6buS+GKEzAFqR
b1OTleP+0sP9pNVRH9akFQBwuVydDeCk+xlkkexDDzop3kygGBU+LuVaXLjyIbTina3qG89TlgW8
V+85NJjd2S3dREKfGReQLDOwSZHelZRwcPntB8n+hP8cAJaF+ocpsHibKoCsO/ESkAm6ghydDV/Y
p3g5QTDGzbifqYnaAcHdMKprzAwzlQ9b+gp1OvaR8EWyGXAWxsFMbqW+GR6C50N9mt/UrW3bk4Mh
7HW+vVRKyG23Jqowf7v+MvX5ysFtTiIZghNQ90bgZ8yOs3X24bCfx+yFVenvChBsF9ptcN7kODck
tcqp1pbfPgt9KH7OfS5OpOUQfCx9zgAFYnxPebLqu7u3Qlq6/3Wg06ysMBdCtnk/VdT8IBVIWSFQ
JxKULmG4QuXjgS+E3+1juJKuv4hmJBuawvRIhTXbPswdgQjJeD9fTwT1zy+Q1qFV7kz8bQwO9E+i
mY8nunq1VpDlRtztoJuKMuFyd2R9LVbeF2HYeHKtGSaC9PWNhGNrtuXDndjBbIIBfOYZHEAIz830
ET283NPtluYxGQRZtRv2hIEqf3zWxz3bAlPUXfeG7JfGsozh5i6Vq1zdqosXJpvWG2S8t2geAox8
8SYlXsVc4kfPsuGtGKQpiMUaMN+CXqEcApmelPBpPu7ygTP6aBHyZToTzb4ICcEd2b0Wh7ZhK/Nu
ZwiVcTpjcN0xA8F89PsDQbwZX1s0vJTWtXoC4U2PStbph139Tddz6YoX3qU3s8sdUkQCe3eqKR2U
Nt/Txq164p7C3r+oI6dazly1dzItGMK9WO0jjvZVFaIamKzpDr7XIHuumXP9zBijmC9oWk07Lu+d
zhyR/nxf3d5Mva7IhJjSz3Xy5SmmaDiuQk8JnAmc2EU2ifYgMmZ/dUc5yu7ENXH5RYOR2kvwoAMA
viPikUZkFKMlfd1Ie/j6OHHcDvkJ0iT3j05QX4kkUoQk60JUiUr/E2yZqlWt0whHm9eM/QR0P2my
zi/R5CNkaWoWzU4JRqIGF2cbdSd/uDJpchSuko7LnAwFgZc3/ocFXCLsXmX1cB/wCIA/zHKIy/bf
aCrtdm3iL96gxIrbPhouNKi5ibEEuyaWQMyrNwYdwHlY2DD+wd9WlJlLP5z01I+4twb8vDQZC7Ya
tcXAY12QKOkaFjCEIm4t3aZQyV3v8rVjC2Hx9Bbw5h8hVt1q1YpVvXw8jotqKLezshkMBZcuZ0fb
nhhgVCCQsTPQUahdhgrH3KAM2Y7fB9a8AEtzXwPOsXCR1/RjVkK7lU06B5Lut/ZIrO9hJR6wyBng
Bz4wKuWGt7xuflKFHja5B1DlGJLXJdVtd1L4ieDx1ArwX423ed3BrNLf5j+FJ/VasZqu1EZ3nxE+
iBi5r7M6bTE4+3kAnhIfHQNxPjKF43hgKPIdTNwBt4ZxluWfm050Zz15YrGpMs091iDWzPz+Fye9
3PpPlMlGUOGsYiwhpkwGZsPavYLngznU8FKHgqnGgvHKN3Xcdnm9WDl+XRT6npr7qyQz0jRSaPBn
ec8SJ6Kt7GCfKAI7QHKlWbF3Crx4JN54tK9l2Rou6Av3xtk9tZW1B7B4sfg7b9kgCB4P/8cNbm3F
Qf+X5MGyPcTk4qaN5KByU8Jeorionpr6B7nbREfQYipt+CuKqUmKeLIhN/BXagyZr5qtXR9kMc2l
sihNxAUZh7JrvQsNFnJpg2gcYyhbJq0m51JXvFwGl5t7EU157PE+oTrZvb/6H0cgZCUx8hLPa7D1
bAu6WdTsOuy4bugqjfoK2SIUXHhHKa65RcnFlEvlByfj39nVWtLr2BAPIjdCz66wIfPFt+Fy5f71
yVnxc8GMeZ9OS4xwdiEPTxJ56k9k/rj2mrjse8nIKQEJM6jzx638vZSo9Dj7/SBlelGKxLqGhAei
EI+JpcV3UGw8uN57N/rmvQzn7YYpfAo4/w0CsZcX1xUVjM67G33JDMqRjlZmi1dO3B1IYgLjKSbi
CbSM8HMbjGFalos374JAKqiT+5vQoeJNmvHuCFzKU8ObepFzXq0ttCRHEku9mrKJL5xoGG2l12sj
L06eAdFXXJ0k5JcCj+BCe9ZAH7V0RR6+29IjVg7RGm8RtETDclO0NnzcWfsO6pS90TdSWCiAEiPR
mAj4bxU0DaBKdVqSEWVgWYhGUzOowAuyRxaML56bx5MQIVIBUE7jEnqfy1/pGZgnPL/X8AnnSomY
KF+dkUHJbv5jLv4wFbb3zCEplrNITjZ4LXZPhtjCVYxbA2sls9NUC2OthQtlFankrRcXKMEDLTYg
1BZav4SdQ5/Ry64+OpYUe0mRFN33jCOTw3Q/PpFXyl+apOteqSGKt8ZsUHJwiRg42Lhx9mSTEbTd
EY41ChnzifnciPqFnjEnzCzoR+3B7F5FqaSUGtgBt0eiCenFCCofWZBQ6p7RSSo9cp/KsxoEktP7
GMM9u4o40zZydcqXF0yTz/rgsKlkPAREiRXV5Hjsqw3KkMm75ePtSyb8Dm3V27+3NotpK65k76v2
iOYsSwwUk9FqRVDJV4Ruc/gJAhlAJuuf50+L0s6jX1XaVyghwgqMJwPj2OLWqFf5Wa1BkFemdsEu
ucifYPKnRfaQ+6kdZ0Qke7b9JVvHkrwIko6qOgMBYsrrJ6UocCDwIP3hL60OdLunJX7hcVFFUywB
QukPO9rSaeMb50y9ugq0U65FetIPWdIlYtUmVcT8PWY4xzr/M5dpiaDD0MflkgwaPLYKEIo/86Bt
mng+sBLTFGMPhg91OqVq++a2ExvVM/+R0gjj2M/In9IGIbvCgig2ZyK8l84dTHASGBFwfZYIGx0q
OuCilZsYQmrvxAPx7QOQ781ByKDElw9Mx6Cf2d4MD6rYp3gTpj59zQ6XwTJwYb6ZsQZXMLS4NGpo
mX+gJ+PlpseTuIBYbFhLiqiEXijH+c86NNXc7lQYp3OGBTkYBBOR9h1XfCwQOsbdpDvaggLsSIXi
ONAhcR1MBBkBlQGr7SXOuhBFkdbSYiC+vOvSd2DhYpKI1fLdtrszGzi4cQWFrl/FkKReCk2ab2XO
B8Bhk4eRp03d/5NYeKFLNMWutSBPuTAGzD5X/8Qmp+AZS9WL6A6Y0oux/idmTu44kBZSwzNI076Y
Lq/1tXQ93L03jfmldo7x5E0c6qLdMZSaK4IepoTJqKkSrQ0/Jy4iCOSg8/IloejbSY6DOZTWPkEk
dznbgF1U9ELgU/6M6P3HJLZVS+0eDu8pGd7iiZXR3+6LEfBwN9u4SPyDE8zyWecTijXj1EqaX9LI
S6CDLPXFCBGWO6z0UwI+SIqR2szIJhkM4hGB61Y3ixifS/fldO6TLZgkeIErdXI4xnkG8TVowvEr
AYs3/P0h044NWYYcJz2rY8uhJMEId+r7YiuZxY6NLToCtfaQ2+2PLQ3nloPu0izvpIneTQ7/YOJe
0hUY7Cm29Fc0eHAQV+fupQ6AtavuhNE7gnvAWB6e2LXL5Oi31mA0JPtJUhY5V1cZotlJxksKZ8Yo
MI6+XA1whkbHRrYCBLZkp8RXUWqhTy/12Ag7w3NB5YFWhu7s+1+cqEuZ3j3bwr2PIuD+pj2ywzLq
o5HbSQVT8S837BPiGbFiX7y6qsd/Cuq8v4VrvFnSObBPkaRrqmIrRI8EtfzMBtgX8mR2JSkGmyyx
Z3dxTckfX+vQ3c35txjNvAlMFxlxLRw2urN9DHzCla+Luzn88cxnjiJT9l6+54HRFiXLlrlOIMNT
1mDvAHAjQp1+vDIZlELu5rFNy7sk4Ja4IJiivs5fqo/MaKpZJN4BUidCOvcH3QX/U4IqcpaJ4Dbu
ab2Gh8ok2bOb39NohNkjQY00CsUb0y3e24Ngd6mW3OHa3tP4lo06QHnb+z3x3VVpwaLY2TiCUjkz
WJY6O/OVXF94z2933/U4ufepLLxnOcwvDGcyEdHroxDpUgCAWIbuH/2pyMs7uCN7vme7qnDjlJBk
lywVUvvzxctb6bdVp42KB/4SkMhG5TxYErTSYXVJlxfUD3Zbmk/4CxDsqkrE0b90wsluhy1mcYio
72L2emLW1gCmIN1UVztKl70cpjrpO2tGsSap335LZtwdRn4KdbCsrk217R0UUoULtrIdyWFGXjVR
NkbYVLuUihxpG/Rm9rrLs3/RRQyq2AXTYYUPe74RJxiJpROliyDslm/iV90PuaC96OPEYxvEVKYT
ciiFbkKCBuLXnzdZeNhtcPD8QFBpuYd0Lvfxw+Ub3tKOTvE0pKYRe6yRqgdIkcQBwgmifPTW6f7/
o1vAPOIuds+EsiuUxf8v8/08N71uXYAZSezazhaOqgfk53qDMWXKkG8OFVlLR6ZpEPhyjf5r2eUE
j/9Z3zt3d9GZ1ioMPAzonys4TT/zScjV/XEdy9bKNizUpaewW3dtO6znIEo5TX41Ro9+i4KVT49l
c5CLgN9P4/hTPbtYT7QPzy9/GGNfZ+nCeJabta6hz+44WgjWeUsac1Xo2tZXDbrphEbN1tfhr965
rY9Dh3Ba/eJWJuUoJLs/Q313FWNCygtxBm+q+0t3b7LzwipeLDrAiA9sVeHh5wo8bkEntxqRWTjd
88226I5HbomPUqSeT7+pBQzZv7q5X9S1yWVbF4qT+bAkGh7VBSyNwduc+0CtPOqnHi1WDevXYED0
KrizNWgNnek7yPLFq868t2FpOzp85b3C6R4VRBuGgOMo3Oa1gA6N93fCHKzM7dgAvXpCGVFxC+zF
3KgWqmsiDemIG7+Ci/qsHQmAlrM5dLfzTQQFjGelmiu6PGwBM2Kyqx4UI4nu8u+PnXXfjlz+rHRG
5Qs9riM+sQA7CAf7YDYKes/dgB/YgZRO+kglhyA1HXHljipy5+39HeD2ai3+7yeUd4X1VLT9//3Y
iuWoWYlTbOYojLDmRMON+I6e8iMsrbKJY4vdi+7xG+j7zXQKSGih7UcvTyxeeY7svmIFsRmp7rhi
VaThPemDx6S/f0GPuDuLlSoVQcPb9r2E3k+lCNFabxUcHhmtSrLLeKVXD6zgnqAKs6cMdKadQIja
G/qyPHeVRJZw/InBjSfpHxG0BhGzjRf50B+MVrgCXuJWzQFSURYd8EtJZTn/WEd/RpgqxJBezpyP
2QHeKIAEPojv/VpbWMz4M3emCSocBSprHqXo/ub1hVlf31vgTiNPj8/KLAGJ1m9xrBTPLBRmPVHk
1OsUjSX8zIINmPA3me9HSuJ3qjnXh0zjeklvVtex1j/1yXCIAubKp4qgk2jSt6bRZL+Ww1KL2JHD
RmofZFj8hfPkuH+cfmpoLTp4DB74bCFnbeWVqThv9mrYa/tsVsQkF4i5A+XW2gDUEZ3y+NytJgHP
V7Dt7kABH4q7kNNBowZKdEmKcovQYvi0t9lthKTA/V1U41IGWc5TowY22Nf4pyl+GZ0ZAhGMCxf8
vTUrKeTsCnM48cQUki5DEL3oHxaDBK1ABnSLzE3NZ046Y4Xp25CQ+zgHhDVT7SI2y7yfmBUpIcJe
O5YYelniCAnmFkw0Yb0abb//4PBOEfHPXZMuceHyg5KxOJCiLBVs/+JaEGlDDKvvS/4PPPugTFQL
LvnEgdDe36FKc3CPKEW8MsOzbRgEteKEZ25p2cpfKG8aPCChMEXf95x7P0GFvxnYWOzW66aPiLfp
r4sd3NIOTAtQRNWCqRq2S7tQGtUfl3oBBs5p0qubezbY1zqZ18l6O8IDuvf/z5UapAP9FDCLbFZ5
tCLxjLbI73mzfNxhfL89EMLZGp9ePl34Akug9vX94TGHKz+0tQ07+lFdHzU+kMhfDxMPU19rBxTj
tdlBucZs+3HQgLv4DWVLe3JUTbhRb7fzvKoZMtdf7cz3KcRRRm7ACTOMCXbB6J3Spvl54/a4BouF
glkYEd/K44uZz1J825IcxnSDYxICraqDtYqpuMZYmCjSkcUa38+K0zcI2KhxOEuZxAwQS7fbD+5W
/yLj3mUma9uKauLHaWeq0otDZ31lAkGCYELWJBa2mvZCfvyc19f01wsF6vYaPmITkMGHLrGZFYcJ
0KPydmzyHIcUOsgIY623q5Az4AyAoNT0iA8200nXGBinRsZmrRuf9j9z4D6Vqd8Ov2SBvwk8G55c
HM5dbhxmoLrH5O2kBnnYGIHnToTFyVAqUERNOxYhkmRh6435+28jF8c6JoodxDcjqDDF752FHNmb
F/SOuhCqJjuDO7/bUu3SCAGa3IgoIQdKndNQpJ2ZXIRERIrmH41jcZVCDCqHkTqcyYJLGhqaTK0X
tfVx4bS86Nr7cbCf6BcgpSVYSk/pgodvBaTvNO/B/wEDmrE1KZdbmEWZWCFwqNpPJGWHJac3b419
XIxJzR4jvgZwLzhRHvVt+e0sxlXxiLSNHjl/9WlrSpYnz6smVZheWPYGzbBId/JMpcITpjOrH3gz
gw2nqiRRhm+3MRsowjuCqB7tnhAuWVuh9RbkI58Q4ws3uFKT7NaMZceV7cOPh6R4TtCJDoCWH33S
Y4Fxl5zx1wAyAtTHXwZ5fUDpwwKYLEepgZFKTnvOXaP2eApMxODKJftHlMOTopn3BZxoVHLUbzpd
Ilj9HFE1xMw1rQ8y6qtVb3ABYARkVrMNtf0ytw4bwXML9oIaM7NCcMlDJU7MpCihB8ZQxG4qFz1K
5NSS7ZLgLqiL3z/ZTiTYNgDSXoJgfkpRWyVYq8o91U/Hi0kptlOIi4CsfRLLyOWnYjXGEQChdWpk
FJwzIXL851dXUP6yBdZRRKthXNZXnYz1hXGUEAfJS1g/lFsioa90WXCmA89W9RRMXNkIIEKPN53i
JkCy2lDb1RAzkpMIROmVTnqG96yt53NQCwN4XJJs6JJdITE9Tsth7sC6NWOSdDA3Xxjiqt1JtedM
/VOhQW1+BEXZRrJWs1RpKCqHGhSQhd3RSQD3Mj4ZCxCBflCi/hbWtAtgpYYZtMHNJR+BlYIesHuB
cS5SoVHC9UaE/KbVlh/FiTyawEXvWmXYJHTWXzXkvk0CpGw7NFhUQgRdwUKojnOh++y69nQX4/xJ
X+xNKU2v6LQcW5w9T6LzNRgae59t+CU+A60pU0h9y/LP9pQWXgqvjv4NWvAyK9+O4hPYAQRMuRBa
pM7Z6Doa43ojoxFdZYhrvqyMtPB737j0Ksi3GnnflE1uFeZQ3RzqRGO3f6p3xKpCq6Se6MMEBX9X
/Tn2GK4znlbbBO6omp+zZH0HmU+3k1DdaAs9uTrGgjKm2LGE4yvZuRJwEI/9pFG4R/xi9SgxuASZ
T+NHkXAFebKIoMyO1duFVF0+fuah4fePIf580yjNgHCjxrtlE1DP+xJP1VaoXP51TriwUGEgekta
KmMJsR8Cxn7Fv/aOK0OomQBnVYl8WQNWq/Z/Z7z4mcwSsxSls/CY3uXuA2OY6wSqPCY8WvUPcAWT
6SE9iIZkhr/I/9MnSMB7Fp5rOUHJsiAnzWLP1rMaXhNQeTNyqdH2/cAxLTuLPzxCd4Bu7zXs0FlE
LgB30QBpN4AGvKbyYhyXEhd/bK6MtCWkAAVTs0s3vg3IB/NtzJoqS4+Z4eX3poIn+pGOXG2OahOx
FPBO127EsnQVUyNEgQVI/YVT9Nx+FP/EzRyFi4fWZZPU/sKOFLVJ1xstyyq8bqIDW9kz6YkkcJMi
6AYaEwuav4iAS/2d5W8LBNxPeU7R2b0l6yDh/VZlW2IP6lt8kInfc8DD9Np5QZ7KKCxT2IdeHdBA
ZjnWvq93ICnwTULsd9A26xLD/XxL3wd0aAXWK8FNAXZzAKs2TPA8w0Bwjg1SI9HK+hEpIxJQ+MQ0
CelWnhM7t4iTKzTGd5boUK+OkLkk3qx2+fbBvUBoW5laQ2LnZNAPBB4YJYGpsJ5ZdCepv3MJhSt6
S0w1fQjmvQWWMkIuawtycEPDSb46HxlfzVxAweBTu1TVZMiX10IIPWmnSs1aqVnOJDYPrg61SVTD
noHH4t2bqpVboywcbXQlPH7PDTRjC8vsN7RMvRoBtnnKoipMrOk35AeLAWByLouWLdhqldqOIAsv
rODsbsopKfh0N/wXwRccTizOW0xIMpwlgDAPqa9NRK+JNjOQDyCSEgSJjM+U2K03PaEjTRaKZ5FR
acxO1HDL8Bt1o8vBdrFajKcQZBI2TfeTm0HVTl594Uu0pXQoDuY1Qaob1lAZIQYsG67KZ2qAZIEO
jCOYU0WHaA592r9obKrry3/JWAIU63Mx9R7Bm6GhfMbfQ4Yy06GLAUb9JzIX3F8EFXhc5qft1Lq8
zZwaFS3zXm4zG3vtjsY8CG0XNldzD0A0p21SLmSvM3ZYHQqelKYfYc9z35XKE66glUYpFmb86WVx
/YXTYeKr7Fqmnhhj/VWnTyJ6CfG1KeGAd3/n4APSeQAbRVedRzWVRaCQay+akjZZpQW0nuEcWMf6
wzRRtoY9IwzT+GagxHAWAWEgUuULe8ROMvJm52KnDS9xt0atFalDKYtIMRk2AYwmOgfCsxnFVluN
eFImgxSDkROOcKieJyhboWWwM12OjV8C7ts8Eq6IMwxo6RZntUJI54ExyUlCUN654PzB9D2ncXqZ
z1uYCDiQXHSOVzmrI+1hWyWBr69e3zNUd+yfWXtPxI0L48h9DCeUQ7oBfCA+ON0XynGMe7fnku1N
aUI4mhfn6NxCUfCC4cRb+i1pyBDW84izwEblUoQTq7YVQsoWo+Mj4LhcQygpVynOIDYN4dDU4pNc
38DiTyoO6B1Wq+4ezSpSpK01xmYwtMPqBbyiq09wvJln/8YpLi4044g0SP7DWqoLkJ3Ce0OAKF71
aKYfsU559oeWahslZlfkZpHfYVuRo7pSWo7N6fx3sZ3Mc1JW++VsqzdAO4B66BWjFl0RZMsYRMxw
ymfjHYfkEJrwATU2IYCjOhBFVukgT7HSn457SCSKoZDNlQb67iyBYMI6NSJ/wh5GV1qqU68Y36kJ
l3ITWrY7IS+AbFZFiloWUQufZzRPy6iV9UIrIu8Y4nxRKQgSA8nk7XITMUIFGxNaMs+c/7oPCadm
BgC7eTE9kwg98jQkPgNazYenev9p+Y1On+hqB/HyVY9q4qNmwAh6phkdd19zaU5RsVLq/1ICaOV7
vl1est1MhOQiF8gW4FMyZArTyv8GpNDV3IeLCqFvAGLLtEFzpV1kxzz6egDSxzxJYNyyhRVSOnjA
r9cdrEGdfEQDc48KMBrdJqtsTpJOZsP44nRt7faa0KNn+njpEjZ/iTngWOqLuKpTbH190P4YRQ4g
mmMsJDvBeLfW0MTRmmJq93x/RlTNl+XeY5ew8Cnh/gdB8kmahPMZFCRzCafWqyL8D0qQGRaduNhV
odlkAE+wtgJ4YmKUWLq6qVOgg0TmzAkuVMbGMQBB1kuuMTyJ+Wat3lmopoGAeaGadq8XUK5smqKv
fdPbXUYK81nqU5t0xDjzPBknvGyj8RTaJM1yor3e5ONIwRkxys2UiGwd4lwOmO6BWnC/lyu4SC6a
bV4YqtlBsmguvRN7SZ7uf8jMDxDIqG9ALgm19jTybMTMF3Pl+4CfjF0vU//bGntCHYwVdxT35aCP
jGulC1POE3EQaMk9MxrEtjZpRjK/1VOAI8DlatplqIBDO3kupIiom+P2CaJQEZ3o4MWEhrIZqs6I
I4a3CGBiEtwAwPRJwpqCA4L+Qbu40wUulQact9gPXrOWuPqFcrI+UnM92jCnDu6zJILGW4T2ZZtG
kuF7VNxDyOpi1LpUrxIHHMf+pp4FEQbaIYNspHc576oWkmb2yngSbTFqdV3jU26bKYfdmR/GGmzO
eSJu7BoTY+dnErJzh9UeO/CjwV55J4pmSCLpmn1vI6pw4fJeqZ2nme52snmAUhNpF5n3ftq8r/R5
Gg21pTUdQ1DQaaNB29zOcdzxdB6Ze0vjbDbpe1lGW+FrlEh3AGD/cmtwFGnUNSCrtufGttXpxRWD
UCJnTS55gXNUBIqiU3lhOr5D/petevO/R3uPYD/nL8EiM9a5EETmNT8z3ELzAeSwoAfeZxTmejS5
ecHzjA/3Zv8UAQwoqh3ywz0NHR+evPtj6Yll1WDYKkXz0kjznO29QPddbiAs4XAUjlaQYZ6e6LRU
4deSe2dsAoYYQzli8lVfR65Ff1BnLK66YLZSlNXHHNF5PRaY2XUxWq1/aBcGtD8siqnCCOk6mNb4
2SOTukwSooZiRuEjDRHN8wOMZ0PqwViARC1+g7m5ID1U3razZe0WEeFpKXoIK7/TAEn9hXPg9ik/
boAIhx+bP573VON//rMRyUjXkD7E6zjRD2DP2d9b+KEy9F6p2pUptmBEWdJwvwFXAdqkOmWoOEaq
bSOBn89k4pm6g7qUfavvtlWzqjKvW1HmHtrNPXoICb/9T7oxTBdgFill+d6I0xjFHpmLmfYD+/1r
RMI//KeoJ6MIuSEyKNnZ77pjJ/lYTAQWin52CgiIXJbeC1b9vVbtAt7Knk73OhIgBbX2FdgybPHq
ZaISnMDgjTHm6Jfrz1No8m5ff+yFqBSF6lS0QH5vmrOBjvExx/UJQP/v88zgpK+jOIy/npPI2nHi
xI03qc30/gRFBNFixhQlvn54JqdSpK7L+Gs0ZLRWMR0Z8tGr1Ng1Ekg2bbOzZ5IhTfNpBMpmMxng
R2onSqZZnLcWhZMKL5FLJYQU9kx5bkzb1nkfduHeT5RfDj9ngFCUExW3zus4fqZUfXTbjiVeBhpo
A3EyvjKaDkuBIjJLufCJy3Vmrws3QibS3Fo2xxFwk+cLJxpeLY5Mq5MJHUqp7FXp1wMDOsCLeaXO
i73VL4JfVevOWcEmsDs0vz4as69+wdSFNuRury0Ire2SH2TmGa7X1JrzzPc0O2VGMitknjtRdKoa
AdWbXaMdazdHc7w+x2PW6aFs7YZE77u0m7R9KmyElo80tAVgsY84bWJUTukPD+Lxm4ot3/H7weMS
hfYxzEYiXI2zcViweYRJgv+iRffLPpjb8PsNZGpj85sw+ZTbGDPsH/YjiQaCW42Lqw40NbSJ0RIc
xytSS5IbpENbpZbiq+v0eBmQGD6x0sem9fkmoo8n2PFM60flgNXmmS3elLzAHi7NhkWhTHrqQywz
g5t2F6cvWo7rVxOCwDUrPJW81r4U9Dt4WUMs3ggi1vkMDuVfqU6dJhyQ22dZdf/JfYyW7h6oUoYI
mNKPWtD0rJzpllb8kqAouXtWvAfT0+A+nqsPlnad90KWIqbRPh+mqcwLqE3AfEKuzzcZ8GTan7zV
SCrtapTyFzVi5XNCG1pRhr7uGI+zDpglAHp6WxyTq+sdYp2D/YZ3ai5nyIqEKbAfwjsktD0f37W2
csqs4Bs/LsQHqnjGePSZvwSmVFQmDyP8xiiGrQodd7Sa6+XH6FgbgpOhVkuwr60w7r15z+esrKBU
WY8cmvgBNn7SdBnk5a/Dc33uOwidMpadhn5iadoVvToEflY9IQ3KQK5ddfPeH5Yq0ChTSnu3QFpc
aK45LlYfXf97jDnYKUCL/iCyG6paXYv0FdDnP0fqFRvajxB63BFuMUXG6fscfQ66U7of7TrgrPLy
8YiPHMMKLxNRQa7TIS2FxWskrVd/72rsmCjDhe2AaqCVI6JPqmcaBCzZ1B+13nq0yTT2nphtbaln
VEsvQlbcDVcs2GyKOxhj7F9Azinn168kq9Txp2ZKD5srEAy76X4WgvZ9oWNVAQNyJsiJO0hF5unt
J97CaKmoTCD83kA0wDjK4WAuUgRqv2KCoaPN6bRgjnnBldDAzRIA39DyOqLl7OqSIrI8eSxzTNhv
RqO35H7gmVWuEe4p0CnmC/RJ1CLhxX0a4x8+kiA7l+NuKe6/VZRw7sF3KWIL9PGSdCG1s4bsEYcf
xMqZPkyi4d8gh+2RSZTEy2pqFb6we1RCDLZ9XiwM0usjfRWTqzPfcbpaD1nCvQd9GncUbpBiC/qZ
4lk04wvn3uK054rPQDCv2wNKCWrXPMb+AkGe2KL0ATpEGnY3GYg3WPncyVVm/clu17BaxypiXUYd
EQ9iPdBN4R5AbmXns7wY/zU9svnMKzltzyUlIoX7R3FD9kHYqrJcRQmiR7FPBdBg6rPOFPOAsmyk
4HwVWUvrLrLahKUnud1HwQGY1xRNAAXs5uVEROz6C7QDrv28lXKjLHPZLkffydyuanysFWympuwC
sGXecbiFqOPDZ44FbzrVWhNTFvcymWVbaPtjqpVByPanr9hM/Uen96qLkydyM71LL0iYDDo6Dz7w
TzyfTR6T/gkD30mAWa9rOXkqx4pSjF+CcxmTcI16HCFszug4fle/7n985pGEr9H4T/TNOcgGhnIo
/mc7SntTtIGSPR1BFH7v3/L4G94u1JyYxIhsisAk6KwG2Q9vhYKNckAYhBGfFL9Jy3BIsjDBthTC
sUSwNXWZsxhBe9e9LslW824uJzrdcqAIEfYkaWnnNhC6LTebs2rXjtpmHqWcw1L9o39HIEgSBV4f
6mnv1KlalstMH1EitlV36lk0vep+t6sAQhYpp/CFxTi8qfkzpcBtJPCQuY4WV3kRSpwCIZB34FWT
cz8fQaYTHG7NHpKt6s16pD5r46xAK4bpDI97PoTKbkauOD55x+nSg4pGKZHDbjLXKo/wGEuz0r30
BG8hTe4sVJlvMrNblHxjPxy/Qrhyn+q08eaagADbwzkW9Y0nGsyZibMN/Xat/hYLYW2kFS18JHqN
uRrBI7W1YFwbI9msI60MS0rHdjhVQRqQQSijIUj00pMQDw9pgmcskGlqqdDJqQvehzE7At/rvTQQ
JVR24BNvsem0lc8DmNDw+09MAR9o1VItUQbGll4OhoiCPDI0LHnCf8QLC6Kqzex0AwPD+c/1YpdQ
dR+9GNtSQzEbfMO0euxUCZXd0qKNTdVsyDTib5NkVqgngGZptvc87nFHqcFCUCJN8WHouVXR1hnU
nZEUQ0gYiXLI/8cC8sHdTizSCzJchaPXCfsrru33201uIMUY5bTd6r6+7Ocq2fVdLE6Im+2c5ts+
a3QSlh4myt5eyNtaESDP6o2uY+teSjYWJAS37wqltAUeIXmERMKnNAcS/dzDMkZttdzX+I2LJpJG
qSTopoMDtljyvZk0UD+hgRXOxA6wKnktzqfBb5JN6j6pS9usy5EN7IDwUoq+8a6uBA6qciDSVa52
4TWKnhpBYnRc1VUl7OyGiRmvxBLFM59WM/ONSpJsuiQ+bA7jRQZ1vzz+Kzbz9WMLOOlh7H35KhqC
Wher16qTSqiqTiCWY5FmLkuCfVoTxlMr7otMT8M4RRH+e/PFDecg8JoniFiGmbb3IM4a8YnvlCx7
NgZnE9S2CodyuJm3FQ6pLSUAgRAI/jHsKyYhNOLQ/+l8tUjCCi5C8JVut8NO7EVNDlzpJ5PTkcSH
xbN4i+ZNC+RWq5MZx+IA8ZYCS+xqBjXFpV7F8FpxYTcC1xrUqfZiGYl0gx5ePtdLhwCW5anJTc39
Z3JHN+avCXXFUoYL4FB7k7RSztWDfrup0LdZy2UQef2kf3bC1CQBc4cK57oqJTFDU/wnY51Ht1ts
tyKVtkaDnCIVK85DBQeJ2xFdNlfmr1MGAa+qwwRrKJkx+qwaz5NnruW0INcxceH8SGinyZLqaXe0
F+RSeN3o9exXIP7pMdL2MBfKN3vcne5CZJ24pzUHXBO/E07tHj22kTDcmzfpISBLDblZCDbXqAEZ
vXBVzMrPj8WwYl158zyUu87O/W7rhUk1UPwA9zFtiAX+UsvFFaNl+EsKVA6VIN1VSAA/yvEddnVQ
B+osFK+Y0h0v9oOpjHtMWpQmt80K+XNFT4FexYKjARR/dKAiePctrQTHVSs3OYNh1I32N84PFNiK
TgPtHNgLBkwXha5AZBqc6GLKF9n53Hh+g1HhNwW13UGUq2bL8/2YslfSEdCq2vD/P4GW7zp/27FO
vXIUVvo5wOdfCKPZNwV+rAQjh5AWewF3eVtqTq2XIbDdXXaJDwQUsvECdlHYgVjxk2n3ZNdAU+2s
edYrrHNNJb0UmtpoY6rKfimq+dBvGCQjJqb8njSjXAkusEIXXuuUsYbqvpVxRsR/IXPUnHYG2krj
AimA0qKW7zBq5ibOXT0qO4hqz0KqORySOLMH50xAnTKVRc3xanHm4f1klD1ftdF5lCHZ6gPSTj96
85Opf+hxESpYiWQfJtyBV8LwCEfJAb9tsxyB8mcAe/9tIKiyGhNb3eYu4ESxu54bOa9IiSqwZPsh
z5uCrrHL13EeK9X8tQD9lereiToKz3WOnySfWC2hvIzX1gRxLgNl3FMQ1v/A4gUGBFCjMvPZ+a04
+KFoHAoM+ld7qSR8SoKkPZsif7iUHdibi627U8aHAkE4LCEpCi5y2dJ++g9c3TeDB+8iTba0SDjt
F4dKnGrp4PCAQhIetz+tVNN9KxH7K+TC9h5Xncf6c7PzMOk5/a9mqcn6yBJ3UlpVHLz0yVG1k2lg
f2cWHrTovkr4pFlb4XHnBF/iA+h/Z5tH1nh5sNsfrEbdEtQbfMpAxk3fY3plIijwN1MZ8ZiK25Zz
4UgtRz1ei3GU7w19/BPY+GuDLyTXuTWyPBZkCKp1pyQT8aSU3Cjekq9JzTMJfkGJirq+rpHPcexT
AZeTf15p8g+M0Kb+LDPLyhffOEDCdJmw8gagRbNbtErqvwDoBfkuCG7g32DbPxCLIHrmddEBTgBH
aTFNk+w3JkRgWqaDc29ZltDwoLWmGtQ/eZXYp8hUJgxM6h6SesbgarPww4Mea+s7zeJ1THUqSTmU
VV60sZ2GUr4O26Aw4arGSTJhObFXQIS29Uk+7dZnBbviW0gCdO5d/Z2C74NMfzE5dU+MFP0e6iIT
wLnkqtiTkwKHJwq13kykcMI2p34TTZLv5bmBq+Q+jUwgOaytjSyAU3YJdTpAGxk8rG0VMhuT01+y
bPhpop0jflI+aD1JdJJShrs2P/+dLKxzJTN85DbqdS7cANT+24ROSrllWMy6KxjsjblNs9I9ZvFa
wqDXjLww5dxeLMGvwYKTVw33vEAohdiMGv+kuC56uq8GOc2JLrMIxV+QaEgGQQ8yuroHwGsHhtY6
/Px8ocn886ksUR4z7X8C91wk0GePwufSrbUSiDuouG9sforNjWPb8K0XOH6SDqmQZSA9qeest182
eB59q2I8zumklRU0Xw8wdnMq/SvqM5Rj1gcAzAJ7DwLXwo0jUQAiO0Rc+qXC+bjEAcE9Wcy7MjKp
RzvglzwKwVDqSFaGzvGPqr9TjG3bG9QbC/mJyUOait/VziIhNmGTpBa/Mt3riyAYlAf4trlWE8ok
kQvm2z/q4SDf1GtDEWZaAe926mYuNzr8Nchb90AhMz+EpZ+vAiVUJpho5zAE+x/CfKzp3rJLcddC
abOzC5rnb0HxUnXMVq86DsTy3M3vQT5X2p0k/T2Ol5m0Dv/GEyEymwcGMPwr33UcppW9kiN0tL3m
AeQqtv+40cpVRFK+JXg7r6foJ5uzP9iAeHhLvPTKEEhNLDNTYGFnaRPs4dGGEWJDA47jo6De4Dhi
NVidWJ/PiIA2YkdgIgHcN80u9gFcxGUFWBumw0UWWFIkr+73YwVT0GwXAFJ+lxRJaofXiALMSYBS
wpuQBbY80/vUQ1Plx+VdbnG//4gUONkkK75bucLaJZIEqrvOATUSpWw+jUt8i11dAXW3A9oT8anc
6kN4UMf89gLMlMYcBpGbgzF0xT69BeAIwuodSWTDXAOiXLc+dgGIEK1T4YvSqm6lXeL64t5wIazZ
gfBH8IOfZm9OUNViqiRVl7HLdBKU7WQ9CsCofClMAfXxIwlHwWuUGRFTIat4JS7kP3pfKmBtx1ij
RGvpQYLWjI7z8bu9QoF9vr34dQWhjmR/svYEjBTRFjg6ANJJ8wENPTfKh1i5i1xxTrHqXS4H7tX6
82dpbfS7tSoy809mFUjw8DTW7oy9i6NIMyYEY9W6LFN8G6sONq2TpQiqnKRdembtZe7p4qcLY+Is
CP+qT/TbBoEQFgywkVZBGOkbHif29M7+RenimSQoYxt5IOH/ssrdauvrffin/Ku7rK2eYLow1G4h
I9BmlZv6e0/s5FvTDijFg5FPtgaepB9SynTvcEjexiVWnRm2F8MONRGXeVsh7RBu093iYP6wAdqp
/TxFqYy7OUIshVZZ6h/2u5pMwulp2zBjF49zuBSbBgOmU7N+8RohAnX0LttwxK743YvoxrF/tuyq
+Y80Egy8x+QuE/yPX26c0Vf5Z44pcQ7EDU/P+u9m8Qq6Jvl+nNAFI3EGAv3DNZxQ0iwihCBFWL1F
Qp97B06FU1YcjvQ2KjHeq3K8sDefjoV1RfdjBtGGHs7jib1ddUrVGKl20wYorXs06y00khX/Vee1
mUvaQDcyiVXalru0xzLz3S9AY6E/idxeKFPT+esNKbrqjwnG5nd1CzC266zgtbpVtR0leNpsQpPk
abRd/EtrkcnOvt4mjq6dMkWfKkrfO/4zTRr1QR7eesmK4xXx2L6Voua3x5XcjSJQLyTsnIH5yZAz
5oJuKOKRgB/IKau5nsPJJ7b1Vl7vmU6WoGHyJ6KEceo0AmWWk1jxOYgUeYPzVMMjO7vxEkjqysQM
I/YznfNudhyvMPk+ik0xllcqsKbdVKqcFZzypelUNh1+2yquB5TiCH+4bn1SUXPjk8LGwDpRMGiO
c4k91pIAPJ9SdctOOl8lfm327o7WncCk1tIAWMNw7u7vt36TDUJJVsQRZY7mOYGvTMRt6gRQvfL1
VaBZd9lgK4s8frT/xeRFLgn/+65vJaRiGsN3pEJ7sqyfS3oMy4rf5mZd3U48dIR9ggqIH9/qeH8h
vR6eLNx+k7fw6oeFBzQlBiFS8rxSslMg/yHM6mPwLMvU3858Q+xENfAZi7nwoRMcTF0jBA5gZQgD
3I9clngQS3Lq7AcqCdG+443wgL7zBesjYKArIVqy4vLFzEfRK5FOogjexShd8w9hGZ9xiwRwgIom
cFmOyNXckyE8w8eTux3TMvpcpgOoiTxk5cVj68iUy2qnugV5TALbGod2v7fAuWBnhjIMjpUoQQfG
vay0xvKzSJwvZdD9b6NaftCnm4qeZ/WD6WymAT5Qp15L7ReEOsdv9KMgMqmiDHT5fjzIk82Cnwjy
lDSneplMXyvFoI1vgn1V/Zu54APhIaBigdSCzCaahFQNfSxXTFbCX/L/ibLs1b7G19x/IW5ZFBZX
ls+AVACvY1hlyGsYJyrNNPJy7bYu09QJR1CT0ZAerQzOkGON7LXMvRQ7vUicZbF2mCajUKmTH4Do
H7Ik/QwJauPppXqucOAzlRmdTQVbZHpUKgDZGfswtKh9eH1Va0VsUTOI+Ic4lp6QDgTUTiZFLGUD
lFwgW+zYEnh9443RgP2Kqg9xs4SmoF04m34/sXTzsTEcR5k6O2YBTJznbiMtALXCbQGt3XS2L+eB
qnNjbrXuUWqKL/TLyv2w+UTxySs7hPH0C86nNbIyP3FbvhtjAHPT9th7OIDYXkzTDE70y1tWvsTy
91oGM9gDdub0CGaex+rp7PJvm28RhHWUAbyoobqHfAQeDBUy1JKGct5NXx94UjTML8srKcQETkRY
7y9JlGhAJ0MQ0T0jmb2fc5By0eSyJC9YwigvhPtuv6b8yf4YwvLneN56moV5P4GrQkft0Va3ndkW
FpUaRJ8sQOjAXVlshMJwBL8Nw+jAmQjn4CCqyfIQp8aYX6mkgdBs+Jv5zdidmOX4ETIXVZjTWIn6
+HEMYTh047drdlu5wO6HseQt8/GA6DTvnN+4BbvOkZ95ZIcfj1BZuLw+03e0GyvZLQliRyLyz5Ek
Ig4ghP9rCMXTgJvpUCDHcOUYZvORRechwyqSRw5/uFPlbeCBdySE/CLPmdQoh6zIrBGZ9+WfQQEY
N0GCfGHcnxG/s3TPSVSKntBLZOZDTfoNrVT1tovvRWGrhfzmb/baHPXruGiPrcZdqNjySPRof7OH
ue/qAXIevR3whjmf/sTytULyRqnGn02wVHpt0YzUzdGc0J07EyFKdq8lFI5GTaeGAbZGxloC/oin
R2C1Rbd+uCZWg9JPk5h3qIigCKKL3novjE77/WKzvC3rmk0Ym9mCrO6g2xP29yIU36bfBnJQud/s
CBPDP7+Lr7Z+vvKmNt/pYdzSdfv3ZIzmrE8tO6pOM+LV46IC0HAoTz4D8impEJcXdiT81KXW5Dmc
xapHN2zjJ3mwJLfPc4thIkhJTJJ9utK3B6NTY1YMUSr2nX6H4Q1XhBCBwIfEK9ACGJ0gTyC+qIGZ
g52DmohNP9FRCd+DUQWFacFdM8WDm1Ip1qZ4EvKtNCwuGVrRIYSYoCKVlkgdLloKuzzk6Ve6FNQu
lyV+E2TrDZAJJfHk0ZVwlt6Lq/xH2vX+wcX8NIUKPIT7zfipeVmP6/h3nUv5EJbk71WwQG//+zdy
g4TiCUQrCfjPG/9N1kOH8rkeWWiS7o0RUtFmR1rOd7d4/R+U7XpupUu5KKvFXxGoJRu++cv5PeTz
aUy62KRxB6+lv8r+YbNQbSw9L2CYW6+SyXkCjDQJ0Gg7+TSPyZOhj2bDhR2B9Yi9FjZJ0CdDC77t
FxvHOE3CNgoJAnwunhhkLMFEUX7tE9X9dZ8HwJTDBHIH9hlCr+uYwFdNUwndMTlRasHk60tVWB+u
sSQHuU0b4OI1u2VxJ//Tbz2+rhtgmAzYM1L1a1t0+WGTlm/k9ylfGplyjfThjHITwXqjhGtw8uxk
i3u9GO3xvH/A8dgTAKyIzoniUMCTu/pNRlezNgH24AGrYgHtVXdes3UHuGVzcfsZT0Qoq7CnYu6o
Z/Og6YgRIfqvMS6HtYd8pCLGcwu6RXjZjD1fIZsJ23/zirmi1R1Xdu79Pj+B6m7pwyds7gD5aSfF
/AkUtf3aIP4N8dprNouYPk878hB3R9wHMJGLnX8c2l7+7NYF0ICRmN7KJWTDHh4lYnsglZLpq5zy
t9oEIGwBt1ga9og8KY6MpAug9hvb38xQ2jFXgpGHKhmlI1y7HNNvlXhh50hXee6hk0JwXUSW66Ns
02wzzMvuVhLZXV5bnZoj05s5fa9z4EALP+b418u0tDQZ5bz+lcsKBD2o0hnfwSmtMsuj7NJqOdoi
bj/T09wmP2vUj3CYK9j5bTRgrXymkW2FsZNO7p077moIXU5hpHhsDwXdsKdCov4BpFBwIanvl0oo
LmZNSeihEdXcK9ek/YMONUhacynhtS/mRKJanMCmWKi2MPOaq8tmkDbzvJ6XAkB9cSpCyGyVMrza
Nknz5mw7txjro7X1cfA3EvOql4onGEHtpVgF76ruiGbbO5uSKKbH676bb2I5XP/4q2JMx3X/hzx+
+0gdDdFFGR2KtzIhZ9jGzdVyiHbLf2kAKCfWDfKXlLZkZpHY59vhB5YB4T8+relVMN8O/dgOW1Nr
w69WDXX7wqU012ULOVhFhIq/kZCiCamnekB0HU3HnsQ4vMa11B//PVT7z0KbOnm648RQdoN9Km5n
olMXdJq2Jr9lPPRAqPRoYqGHjsEiaSw+OxoOnmUCWSjPHvTILbEkO2wTsW4ieT5QtzxFKzSzKmZ8
QGOXvZIqhqpExJIyjGVWXt1XA8HjDUeHHIJaVTFiDg0LS2k5of9Db6D37eq0MD6nPf6Qh99gSM/o
asSzDqrwaalIQlF9FKi6H7yDRlroCXnnFu9CT9dk9zLEfHsWkj8NnH67mm4gOpT7OjhHRrLaKWZN
KR2SFwF4u65xmNEZtE2/S0TCPvwMMoeulV3FYMeTsf0MxhPBkgkvceJr9Fb7Y/94lrbtk1smPPGW
odDPCmZSlrQ664pZdAvg5tdpum6TblXWwW8jFiSQ8wvHVAYXFrPwc5OiJxvb3hZ3qEQSwxTBxFJb
mlttevwIRz83w55RFmalWYFoAyjoUm/pJjcUjUlOdkn7z3NDsCUbT+mUFb0p0gMf9UzV1vamILq0
7DqsSRev3UrKiQWkxhNnLwJeJeTDe835yaGRBfN9B+021au7XrBeRmkASFpYrK73weGDJV3eG1by
5FEdx6g5qbHpC9fymQYK2c87arMeZR7Egu0PXJm4suZlCkXQgZiKdK2CYETWXOkWBt6xcKkr41XI
mU3zDFz/ni4NIBUS5mX5h3/ddw67r2pagVelI9zLPAc2j6oZx0UZvHKhF4TdVYE1CN3n/Ph5wZve
SHKIE8gDo3DkEyDv4dzBKH0EBK1sIrYEGG8CO9ZuTPfvfqs7jgJABqkH+t39Omr14Sx8l/8UDUg/
EG1NQ0qE749o90Y8cjszL8j+22AZjS3eolcytSd3WnaLXonE/aRfC6qY7Th96ct15CPn8A58VySL
hz+L/y4pbAnCMShGmtPxJb3sIjP0wgddFB6rVOPe4OBU6PZG7yzmbNt7M70+E9mMDLlqHzmNCJVd
klAkwStyEBbPwxNGlZZ8m8MZXgZ2PznPESDpwPrOkHObzTU252fzdy5ayx9gSE32VnRV59tk6edw
Sd3pGXcj/Aub/pZAzMkcnNLfwEaVREKcgPBUNj3YBvkj/tztVSVBnzZbdsmbxWZUhGpX2dWu+lL7
hwx41QRc4AOY9v/VxBOuFKAk2r5cSBEzW8lt4RwjEbyNKTlww9mK3zPSuhUq75Mxb6WQ2pH8Ik4m
9emFmZWfDBC0kYs5Dt09ZDUfipY9jmqOwkNK7PxCp7iUnkPGWUUnnBl/qIxbUkjB78ey/KYlViXm
oqFjik/c+FtyU/JahsMEPZ50lTyTBTICVjQ06NKHXnsz/nGg5ji9sirkYtSB+iAe++k6EvElnTwx
VefJRf3omHQ11WRDVtnytaFfvuZeNWoAR+5pZH8M1B2MxA7jptiJVyqnXIYQqEAHf9du3ztBCQe4
wPeIRNWH0L0UohdLfZQn1YyugZK2xX+biYaGKZLW6sLdrdjHi4h69A+TC3zW2Nd0rlY51E8Y+ofJ
/PdBGGM4f0Oju76wfKZJDmbRM1d2Wx5xZTdIndzVBPpSLUFkpASd+qQJhL8fAQjfolp9MtsiFbWu
aYge7TUbD3RV31+YRmeTp0xS0c/RE+GP0jdEAR7ZxlQ3LH2NjATvSji6YqeGPSFtnAyx9bAxxn32
IGdR0EUsKeYkCJXQlQXl8VA1kzFGqJcYY5kADA0mIdm/HrC+CugBShE3kCxcXYHYpHz0UriFjc9E
kichZxHh0e9zT7OPELUjEx6+/1+WFjIKob3IhNafzkXqIzN5bPgm1kWc9mWJGOr+Ox48tV+FeH9t
qViZtiFTJIPdedA3ZkLdWkLblChsFHzyf9sjl5XnNgVZdCObTFlsv/xYAJ9r6e62ZGF7FQCBH+WY
TOrb968Aud1rQlzJ4cYkGUWs6oZajUq7oYGpEwDwTV39phnjh9HlGe1hxraHAOKAnp8sODci+MIR
/U/A8a80bvR3WKb1t+YJliqpg9oY4eJEtNU1tGpaNcg94sLwf9rtzrM7VGdO2lCb8spjZJslRT14
xkS1T0SOGvevpNv2tiYGnp1JESYf8rd9sZA7eRQmWEyRb9642/UWdPjuqHi700mBlQyoeUy/WPkC
yuXYXEy0YW7xAlr7i6ookiuMQRUBmM/hN6K2CBiYSENLo3+hVWFsEcoIiU5fdHWExSvZfmchiUWi
VPAqSCm+cTUuI5mWMbNHr/LM+A5AeTb7wgWelqKtQ9QFPM+hU66gJmHJZiu7s4bBa/N8A7J4HG/9
dg807wDA0KeQ+mt7VPBjp5g5QtD05zAvgoricrxh4cIWK6a9wh0QztMqh6HY6/GiTpLiOVfEWDod
Kq27tWaGII9M9EkBedW1DS2LIgd1dtb6rl5Zh26/ovfyMNiNx++jpkwWZ2wzL0em8xSSwGXRzK7f
k01QietjOx1mWDyrC2ROyopAZUpN4xh2KXXgbfws4auVJuaHCkyr+3KcZY9oZZw7vjP7Pawd9CAZ
S81z/IREum6vAfcWtkL0nk4LYIHh7gFbmDpZ8cHvO7QVZrQ1U/Ku6yGaDnEdUv8YjcQZ94BWmSze
7zpsTAYJIFqLwit/mGVpI5vbrFKj6G/KkRG1eetwJIhWkSq31tpfLCdUaBAQIfixH5hTeQYFEEXb
j5fjYCGOgZGWlDd5sRu+Y8Qp2oBhjpYN033ch7pjpKYt7q6GPpPBMON3G5kxxza2PSKQtzDel51W
JzesXdjzQnNH7ytCtbk9czAdH8/hi7jJ2amTdV3zijBMAt/Or8oooqWCy7Fv4a6Wuv4nK1l2Recq
EdUIt3O3fzob1NowTZHeQQQTYRpoFbGKSw7ZU103nvUvvJFxiIEPw0tmUTJ1UdLSsm/SgyLfShLU
Aok8S/8iwS/wRLVsafWuBSEFErVKwP2URjxe28i+sXP/EJ2n0KXhHrsUZ3XWzcMPisQknI3x/+6D
hVb6WTAyIbXO4YO3nW2OZd4vuu1S0lJ1Y9w9aDkEtDFMHpeHU6f2lv9eXViCtk2LqBljyQdi0fqf
8LCoqy+JWO/5oJZ+Da8WmlXP38GTCZ8jhQuSsxSFh5fPIVEL2CRENGy6auhf1s4w6QYqtnFFzUvE
Tvlc6Wo+LzYjMOTLYER7Fc4p8qEI4GXNZTQ3vCZPeyti/ClQGPUTj4dv2yHRtXU7dltpBDt5CUgy
rDQNxgQFIum/iUQUMjZdWPVIcf4M+SnI1SFh3owfkkbg1CX/MYOl7TlhKX1TLuQOPvNW86eIEghu
Kg2SZ9aWhUqGHPPpvFighIMBh4aXZQOcjE3hJLVUsHb2VEmIrssyGA+fYJixP3FRex/lq4OCnX1Q
1am2Ygj6l11oaf8vFNxmI43n6c4aGXdqOMcUH4AHIOxVcyHRUvZ1kA8TRq91t2LNySLg4xxNY4x/
6PZa28UIBKu0i4Djbv8cb4+tS0PKPx6tsp8kYWIC5xZ9Te/2vImGqWz66VnROpwZDSCm2VdoWQ7K
CLyKB8kSxC4MYRb52kaSfdQwTD933EtHcwvbWBz9AqqjSHY7ypS8sFxr/o+/NCzCgC0bJzrS3/34
wXvFeUK7RIlvGk3GE5tQpsAjKaWmON8kmI6hXzwWTaPPkBEp4NrwYpA4r3qdrC+b2QYXf6zCadci
H3iflVe8G6ww1ImTyIFuKPjmCM2WzDsnY+SakqAFlJWe3nTXFCdBbZWbLafHCHJad8zXiIDJvBHR
2nAvOrRmcUiKtBQlCEGn5+XXDYuLUxQqOvD7lsgfDc2agsZ4fUuVO7E1elr369tWD/Y0yyKHgW7f
FffVXvw+WA6nKHJvAOFd6m2duBAaoV6tVALiX3qSR9rNyVk9SfAGAyPudjoAWCPcV1PThaPChgB5
jylEpNdBqjhCrjFtqr95CSLDVzVpuEa5cvtUX2PGwuse2VhGzSvqUzWZGc8MrC00fVuk+uUpwHWi
oGcKPwS16Cly1FChE7/3UYyipC5qH0EAxjKbj2KybRg2BRil5yyCZwXJiBNGzmTwfOIu1LpH2H1y
Wo4VT29IsDSOB4EnGTtOYe5NEbajab/WhtqSY/2fVtP4KOq+wkHQu1KjXwDAvNu4r/qn+61858vF
V5PscW1HzpXUYVtdTeguX4BsVU3I+WWmsbbjNEzIxytlnl41zUWDjb5NkMk9Vup8fC7Caqr5Chsr
JpHxHB9vBfhdZgVOyUhNv1db9eaHbKWiG4ZVh3EpFuQoOpnPduZf0HFnrNUV9Xrg1KnZOylb1HOP
g09O+bFq7+xEKtyxOtjQEVz72iVSYUYC+6Ii87n9Gmb8hfrgotElK+kwodXfe4RRl3exE/3EpHDa
6AP1HAToaLqYpmgQjXap9Z/6OGq7+JsziQUdlpdhzWNz5DRkulIoPtymO0lK1NUNnKUzLfLU+cdq
bRmhV9iS7cpbWAtePqNdfH68OBSJ1h8HgupoJcythdTBfYsePZIfCq5WpQrG2EmrTFn66GLCl48g
mKlMpGM2K8xs0BOGPgQeiWoeyjLkautDRbpFFJ885itZprdxrcSfhSk2la6qnAPlEAw3kLZ+4wm6
TJjQElxSWJOHjuAkHLHzu3KqLxRtoqP46EktzQ4/6sfTVYebJBCegHandf5t6vb9Ex80FAVuhXUr
wxxgNbIX7dAINK+2Vlh9f0GQdHZAHUwgIVB4ZU7apMg1p3Y/BH2qB9bRaCTQ6cMPW+24EmI5uXUZ
vKmJKfj8Umz4FRVIUYjKuTYUtuxDK/mThKyY/J6b7jPq00dFk0is6skMq3II2y+T8JbLE8TN1jcN
0cFyUV5TutnqYTWM8FwI5nY/hd3XcKT2pDcF8mX9uOIe7mfX8MVnLxJhv1PD660PJAgfpsi5Cifv
ydzhqteZCUtcsMIJuFuqK45uLiJNFcDCFuP82e7jMJbGk+m5maN7YANzWFeJwtb83bDD/lZBO/+Y
jX6bpTDwGl8QFR+XICRK5jLgI1oHXUwTZzUylhXEO8u/Z6+KwQNtVjtgZLTzs4KceRZDZ3pOTQjJ
q3iGhAeJRRkp9h/nJicPzd4GCtEGH+peMZ2SfyoSf6drXa32CNmi18mbnjDSEw4HQ7KhXuXvAfs+
DeM5S8vpnBAHa9IRRUwqy9Bz0DASfDSpUuZ+95UIa2MsdjBTc1BzAJoOylrCzk/OlI3TZN5+5HJV
tqHSCJoklkv/Hh9BVy9/XiiLUrOIFpLTeBybkTc/VotJIsLoP9bJVGiJzLkTI0edkD4lr8y+IQ4p
BxK3/xCZbqo3crLxkuLn8Mrt2OHRBADdiFg6i9uBx/mPNowaremUBijMJxKyCzK7cbWWnJdKrktx
QZzzMt47BMvE8BP8ZbcEBhk3zdg0n/nDaMVoACuDcb+VEPmRN32zsvWoTJ0dfrQifTMKnQuScdW5
EYQOpAh4a1RPRu4hPjOAfQxVtlJYo759z77nNC/4IIzMRBcLdjI+kl41U8mNYIQVXni0alQmGKpA
aBTNp3r8UpFigvXXjHfMe9w7uNRBG2L8RP6b9mUajMuerVKJRWWnymsude0VfTkegp1b1XIQA0JP
3EP65cBdoSQ183J6lLjqig3hsCKHD0oyAlG+Qy7vk92hawzJD5/65QaQAqVktcKMr6mK5Se2HeUc
ICMkoDKusoN5aF9/g4Hx8QvOgdYHFYXyiyS3GiHZZ6bH3rmYw9oUK4GzTIZ3P14rJ/HFzsZLHB6X
2TTlZTzjSuEBYWkAALnn7weG6Ii6uZllBDiQK6zXn31tPtjbKK1TKA9mpqeobR7B2R8NXtLqJh2z
h0+V49mce+pu5DeFiDXWQcYV82jHLoIHG+LtWB/1YCG1dCdXL7MuwrYLAV1ChJGQGltYibPxidEo
fLmw16uuHzozbZqMxLo+X4ZYKezaFwma99HlvaEMqid413fMZ5Lk0oGAMPSt7yEy4jS785UT5Mb7
MUxXgMQfDhiSH0z5q/3ziUB+Ed+OdlYLa8FAt4vV8nqD3cTB9kJEjdPwfNWmwf53lrzaBNUQo3q4
ouTzVjC14u7/BLEssyh8ORK3IHlhAT1SGtW2GlTfXjDpLjG7u+NzuWfpznmZZS9vONdPcT9TLWey
a8OvEb3aBrsZZsgCDqW/M3MKDujIrwvSkaZ2a8AuDMLUkAzopmQxPuAT84xxAbYOc7PbcYhKTw2x
/348T/HYZgVnzJBcDVUeQfmD0otJf3iLm6oBeijpC7frtd/L5wUAIZ1PvIV/EnRJfYqAfLACnZ2U
92Tv8hOFyyzWPgZ3Vd6opyPs1yPAYq6ln8ZpxykMtj2I9+h2sGB8Kw5kPDg0rEYq8tEPFVYWgQEE
1I1Wx3DzXn2L3GzOR7Jl4Nruskn0yrRKmCOVpZrFmBsAjB1Qp2Y+07RDpVtU5DMFECNAepgwD1b5
wOljAC33SYSvp+KCAnLwt5vdjRCofGCL65Ogi3JHlzRGAKG91YwOoQa4o11EUB8AWvTMIFpMNJkY
XxGhesiMZKaiFui0kDCCOuV6GxtITY5b7TCAp89tx7r4Mcm3Cy8iwXsr1ecvW2xD6xwaMShE5sGg
KI7B8Xh712Xc1gR4/4xMV3HA3NpEas2jpTFnQ/850k8YgpYnEK5SENZ4Wvpqv3+V/H002KkEsZlp
pzzHN91AXov6VPsykkNGo5sGLXw0fwMGzWy/SK59Kz+xkCnsXDDyCj1yW6vdZRi1Lviur0dohUwA
kT8flpupw6qcp+aNiqO5rsxplMcML8J2QgCGJEDL0oHIcSfXEAlgCRppI1BpJl20C5+Fl1g9Vvyq
bObrsxRggBd+0o5bN1GH7cYKJVcuxM2YuE4FmdYCo4O2brJzHe3/H6fl+QcDe/aNV+mJdQyPLhn7
gtCMSu4r8436RvpwOVkRq8fH3kCDVZD16cNkxOo4qVjNsmN+XBxHvFx6p9dG92N/c2jtnuO7E1T7
KifvdJO+e1Y3XLSmJdE/LCdCbbmb+h+mDj5zpIQe4c8R31iTQN4RpYeCbRX4VO/5ISvl3GRT0kaF
FxrRqtAZj2ThuwPfPEa07AB1DGGSMj20fBhJJEjRFp3jOC7mbEQY2RG+IuVU1SSlUNdmLGtOGli6
NugCVuGz4JSeTS8FFPGxN6gdYDd7zHBTXpfcPz55GiHrG31MjjfFrI0QBzQ+ndEboW0qtAwmvJ3K
URzX2FRThe2XDfC+dqyuDij4j07xzu5GNcFJ4GfH/KJ7Phk4B+YH9wh36XirFqXBlrjzS5K0lsy9
IgMa1kRkgp9IoD8rfnPMT2efKvM5HXE+x0zWCpnKD3TPRYUgIBbYtbdnh4qm7zazMf3eJo3vYnQq
6n2yKMOuSQYYJiyo4efIyoTmMxpXZH//9HSOAiKN4NyI3m17lmcHn42Ee9tcbeabaJEwnJzjI9kV
tNCtxl783RcRSSVkEOoVAB7+rRvbNgfYgiJFvbWBQQ8/NJ8K5UCHEpCA+ywcguLeNkLjOqiUEvLD
fCCW8xixH/UFO6uqrLiKfmisgjVM6dgDPIOCVqlhBmOQAZYL+PkiA89/f8snn7lcAjaCKK9wICGf
mQg9ZGIqBqrYDS+AtsoveYfQvVtOMJXkUSFLejZ6iBP7gMhi1AK+rlZNfmBtoaEldC625eCWmbQT
KJcPpy/FUDtU8UBosE2f58E18TrECIll6a/3q0GI83H7kHiFn4RxwxJL0BnHOGnsQQvCpPnTfV5b
nx0ikknL3GawceIDxZj8NBlP36K/L01z6ouTmholg6cJACfvIWmiwTpTix3nBzPtQgouOGiBOMnM
hG8S0pW6GnpNPEazWDyziJ964/6ozJZAjPF4DS3JK3n4GQt2hm8qwbEcwIuGv0f/I+KcRtlzWjAL
a+0JgnNSpMA7AQzUKmURaFZMVdANizw7zjS/BJETDpHavThjyQIE6GMPm5+pLRyplzuO6VAGllFg
2T5LxHhNRRbOih2He02T/zZZPaWmQ5SSOfrPGlp1EKQvH+ILe/9mITfeF7jtPSD/OwxadvSost3r
bs9QdVELJ0RAXs/nPZSlSU9eWMpwebtnWjRTTH7vfdUacdbkcreOpnkZNqyMoRIKQtpxMV8fJhfQ
2iSxHtnr5seJg8PQGItw907X05O5iLJJRhmfNL9/NBtQXnWVR604XHP8Fk4Mc7owi07y7K88/XqJ
pvTtxBFoAe3CDny4uqDntBywZpVq+OmO+qicUEoQ8bhMODucxUKuFetQWeZaKY623hiZUvTAJj3t
YhkusMltQvdSJGPOV/xKmUSzyjTF3gfy3ireDTrx9xaA0P+qhEcC1eWOzxg0LClmnBXolqZSiRgh
D/8j+n8dLgkCiyEqWuKFWDDAQj5g/U/3e1VCa+CqCTJ/J+xUwLauC50tsCX9VYw1Fz14EgbHqvTz
57nFPsv5wgGmuEBYIVcS2RCKIMdmQNmBbU96mcAAtxy46Kqugu5zijmeIQslprkXvEo+jj9jwX04
vuiYjEa3HJ1mdHy+vQB8milZ3bRIGNf+/CwfS0w49fn8STo4BMCDfGHLzOS7GEAg9Ara2TQ6Oi0f
FzurugOqIkJds5TXTsPJJP8GCuIdeODk1fAHJqn9n/mtOSAEZU//P6w2w8m/1YgN7ymlgmXaCndL
HRqTT9iqsajFXY5A2e+chupAo+ZpE4fi9W5dnnkZp5eOpLihcWTkSWGaMb4Ed8Kcmr7Zz5i+BpFl
1wqcuDgBOfshQPYog1HciJBpoEL2mTyCcGV2mOf2ZcPAnxNNkSq/IXzdLu5N1y5Vg58Aki4Ld5zz
duh0Ku6+aPI0RH2Qbh9K647OZuBS4YigoVcNMxS6BAOgJtK2BvMc/NXpYsL1u5Jr8ZWlILARED+P
iHdPpJ963X5yhzbRdAMJS6czGkIamZOyl2KPEv6I8+Z4AYTNuT/DVWeF7EA1KBK+Pi8EgQTRi76G
i4RWcHLig+hJh7LUT2kDQECsqx/J/drgK3hd3JuL6S3rbUIFSECucFqm3hsBOe2LhPtNfHpzRfjZ
tSS2zwEmBQayCDLdGevtymloEc4YsS4CXTFA18Y4GW6LrX1vReBHVG2mErQs/6SkHO5GuPl1WRmH
b+IOsx/w295URKbONTacGf8iuWC/gSFRtWo7lv0y8fAHHg91tuPSpw+cOENNPcC72+48unzqPRDc
Ly6CjEc0WnO5Zp1+UP9hnIDiOg3qiCgFGW03l5Aeo8/6GyTeO0CLuEVzYOAMN+jiZy4iPMwQu1oH
dKdw6AFycY9FB65AXIsgl9v9IEnzytCR6TdDlv2AK+nXlPvTwuLSmqXRrX4fss1eukAyj/DWchqe
pgX9yWcs6JIiG/EDOaC/jhhbiDpMqdQ2Z9wVgwtXZh4wRrO9pKT3gaJx9Po+8tokkkd0Dk8dDJ4A
x3rdx8JkEgXKNLzDH68xt/PlX3lY+Ju3JXDKLgU89/lOpz2KfhlG3xrO0P0R8Wqt3f4+wk64x5DE
mK5hYnxTgDj73wgEcVv5VnwCTZuWyGx+5HyuDoS9hioWkxhBMc+98mEQ00lU7oaTxL7C/ucXZhd6
tEY/V6zaLVzCt6a7LosQUNqxGGj0au1aH6UL7M5yvjuqm1NbXaHvAU2rgRnDrxnLfxX0wNr5AADu
XwlLmLNuKb3ppRUSg5fMD5I9kQW04Mvhmq+cDiLBd8v9HnTruazzgd4W5OoHLgLN5o+CyPENe8cB
CaLnwPcv0K+YWZCoZr+dadJLWNBUXqVRlRJKIjauzXZvj9EVCcSSYmhCLcEh05u6NDvgKWnYebvC
BuVqavz/5TE6UFL7T0hel8CYRCHyagIO7gQQRjo/MnB/7eOyleQ70uGmj/uDqPXGkUiIdFbG5Pwl
gsFC2gA+h1tvcpT0RqGP2qHlrp4aJ7FLdA6mWqPyyfFPHhrb7s5LAY3IwgYNQ3k7RHD7Rky3oRjO
kUq/3mWcl3zxw6f22bBLVYTBy//NGdkVI62UPWQ0OQbcYiCkoRd8UU9hDWkFmPpjeDNdroS/OPxX
knSboarj9ZGFxNb+SOs5z71GVpq6CkeTxfD8lUcQfrMtaTFeDLIBjV3dDbattRqyoUbuQU5PvSJ8
S4O03AzTxrtjGpmkNcUBEUEncOhA1G564buYDao4cSuTciJIQm6fh1fGF3LHrmFYvUTPZs8FhARL
FPkxMQuGIOSDxHi8inEA6hMByE2qcpgpdoZgITlrO/483ChRFgs6Bx2KC/ghJ+4XnQPmu59tD5e/
GHH79M1fJX2MhTVXgHEKDcfWyXdm0RIV3Jz0ubLjBdcbgSHQ6hYGs2Lp9L/dAveDGCEqsYeDnOJ4
YyYmmzBsOH/jfrQW26v3H0Fx5/kC05jfpPhoGNxaZ8V3WHpd3wLbQNXJtK1YqLb4jgScrjjPikat
5siFMxkILat/M32onhuv2mQN4iu+6PaDpZfV41AgxdzaXqDdEPV1USD6ZI4g9fkbHxyhxctdhE+Z
Dv0NWZtyUf5lB0s612OKzFIbXRaI+aN+zamzf1EdDFkANNBsIOpYpQ1BnSDnygfY6r5YB1z1Z8hY
VLi2dfoTJUjzf8k5whphLQ6gzh9CxJkW5TsUZFxUZKv+JlkXH74tJHnXyWJEL5aTd91KliBoP8MX
F6/KSgWatNgT+Bv8o3EAuL+o/rr5Y6kodvnQEubVEwa3WN3/WX9dkbnXmRQ1UgTV2iOIVJw6qTxQ
pPsuY5C4tmgL2Pa7ClvA8Xm0XVXtiXHpB3B8lQJ0o9jVjuqa8Sr/omYv5jfiepLd+hvLLRK2cjMl
84zLB75fX+DytAjg+MlN5YcGw3b2TaNoCm0MExcnNj8NGp0UzOE6oiwcOA8e8PN9YtUUEU6gFluD
6ewZMUlspg5jz/c4T9YHMfjs0kfdHk9eFY/AP4u1oWL0bseVCtR9nAXefAbf7rH4+FldcITTDM9h
9zZ1xZIu1qmk5Olbs30Bs2xeIH66olv2dviLnYdzenZdqRdz/QayCG9MnzzoDb7igxRL+Hlx4mPj
UbMoOZcMIat+JkWqfguA/kEsx9JA6C5G+xs2PWIjeQW4U7wFQ+2mbChrDkF2eGCTvO638HekxCtS
byCsNJRUQ685tLfblrcpmsRP5vaRhYlF7VQYiv8jz4FjHLlGa/YzufV5j1ghblTGlsFc8K3Ultzt
+Vt+jkBLHN8zSrQn/d3NAdx/36vbxtHsx8+UaLx7STu/ASBJi/rYL7oIJCaFLGAd7ZAd74yNJJ1u
8ntM0Uh0Atb6ZrVJxBs9hApINkOcaUfDVghdSMjprYAKItxmzW1ek/5YM9Z6D90ZITThE5jzvwNA
rpQU+ES3UzDAy2Xxs8fhWA6avgfb7MoNo3Xklr+37X82R0a1HdgKRrMmhgZ+0XIsDUSajmu/v5WP
t5g/aQML+pnHhK6i7AYBzMKGP1JRUjVSTj1mI00Szy2gl9BcY9EQ//hQ1V9tfTtIIX1RQnGofLT8
pAJMkJnvSNDMXXer+id9Vwj6uNainnjhKF8eFAeHkLvw83URLiSLrRXbFHAWW6+do5UbFeR485m5
NpOvLaVtQPLJKwSYcIV5l2gwUxSD2IlxOHSlmSDgeJd1KDsRSYiIP33NAql4BuHH/u4G0M83IOul
NCIK6gfRW1T131WQSTT4zGSr5wuaT6t8b4WudrrkBMHFHNdCEBYXoWR0aCRQSeQR3feavhX7onKO
ireeubuD8VVBk0xrur3b4iPrv2qPYIyb2ACaDe3iXCL85AuXuTV94R3ZacDQ7E7X+epMqymSllLv
/ZrGRtgXlia52H0sBfzLCVPCOi6ie/+n7ZZL87BggL8stebMwtzRHh2Rv/CXq5lpAHOmuaCXoUi0
RatnSbrFbz0WH/rPxe+rodS9ssJOGoW+PLmO0b2gk+4PqSJ/jIyB3S22SvKCfbj09b7T26CMSGru
6qzs4frLcUla/h3BevY4Ovy4OkSUXUAvedSSW2qQhu0s7hPvChCOUvPiHGdiFEUbU2ShTsL1hJqX
Lb/f1DefNqWNBIXglQUFsFxH/L8osLr8Oqgy3/QGxRmOUOqnX/7YQxpZTcHFRTk3iZaEwZNbrx99
EQnX8phC6AuLndkjvv6zCtojz8Yyb6TYsMYUEKv/ET9M0wkGlbaFwjv4tj4pmwAvtFHSsPlsFXMA
X6xipsrqww7nvPgOeAXckUU1/S8dH4pys/tUGcwumCoAOiFxKemIBuSHgyEdvf3/B7ekWNhfc5w0
HvtiRSEVt1GdvTIDmXthgNRfXbaXJ75XektuihTzvdwAZ0WOJ6EIHrRWZWTOOADfZL+pY3mxlqa6
MktgwY2bxL0wMzmYb/AgvT15H2YOFoR4yc2Qz6ZtzdWXXYtU4YZRTOMHkrMVqfRPaW2X5mXPb+Gr
h2MQtdG3J4nyQXPvsIEB23swfUMEQqpnAp0xBQ9kp19deWHARM7uNYhKh3A8J42ouODsX3kRV36W
3Lkuf0U0K0tuTAKNe4guae+nwT2yjNmN9HVs51O2KLR8Jxb7cz5InaKS0a0GDnEBdWk/uCX14uay
vsNQr0eLKtRYjgoQJ14hxBxxn67kYZQPaswUtqnGeT2xpSI16zF0dsfGyag6yBFPcWWlvBq24Zf2
s/x8QIc1Vzo/kZ/STk1N/AHDFEiJWmY6VBLeyv3csr1bFNic9oYGGCEGRyCsUh/smLpvD57+JnS9
MHsSi3T67wYZQW1NmDcO2TcS4hJSlNAGlDEREZbFd2GKScw9SuuKv5HpRKsKR3eMSLKunA2MMywY
bxyoxpzJyQwCV+I8hgUs4t30NJQUB3Z1LykxbdR0HJ8ihzQEz3UIKiR16LDujCD3OlQm1kmlhz/f
cBLtLzGg1JnowKzA85sE7SZGPHGsR6/7Tqy6sGzICRs+4j2k7lC12+tdXmjRZBFOs0pM8WmdpiaK
VQfkJNf429KIyN4CPY3oKux2JLQWFmQ1ne2vjgA1DkkCwg/e+GuTSXAYvdJjgDEKVHpgflDDvclG
587EahTRuSmclBPJqFdFTRCVPpmNbBPGvb/kiOogN5tNS5qadyAr4yyNjMOe+03bzw2kdL46IUw4
N8S+k9DdrhiwncIHoXlPlgVv5LxZLL1LuuKFe9NCekdFJUCl0tXlbGiyUWe6zeHCU8ZMt1POjbG4
1UDLi2qHP/fqRHhRECoXBimcDWKCbbMtniFPCtyVI3O2VpoJ67qcN8dYt15U3SsFgaOSCgN4tzTc
VszSOIU7kZRegsd4vJxMhQYGzvPzPHnXI0HdK/EWo2yainbT0HiFas195mJEroiFoW+1Ir3x+Q1Y
HmSE6zlS8RUHOJ1rTQD7uXM2ICC5f1u2r+tsJRaqZXLPjbmPwIAptVp31FFbqHhhYkr05mHuXifV
GsT7OhBKdP4StwdjDAkNUpzTaTZsQe14Sse5imFyuwblklj+6S97djFTh84O2YRTNCZjh07SN18j
eKfrVEvvR22KBmGC7YFbOpzwUPI6JOGjFYYco0AZvW3+0smXmmADhJVXblob0fk5wclRwC2B1nbS
CnZrrOvDPlWhVsDUGqUf6S8v+sn3Ih5cR5CvRfyeLeyw4X6w8SdUuQWFy2uny6RLU3Y/OT4yVuC0
9gLgPGQEecumyw0XdxXorOAGQ4wVagyDwDtlhqs6W6yvO1A5ghHzmtdIkaP4yieZP75npLYtUGY9
z6EAX559yhXsFmS4aK1PVucQ94UPdWoIfs9Bv9sEPwNiPhfhMyF+frzsNI5B3535gOf4aaE4Mgob
CGf7qCBHXEu7PxlifgNLiGqT0bacN6LA+leQ5da6Xm7Afn87O/bxMx4PT4sIe49TGfx7rbTgt8Po
vUEhIwZMl7UM923VOC04fINOuGutW89z9o5+lx4eDnktqAREN920EpNy5VyqoVPqelQT6p/TERmT
kRt3wLG2g99tog8VvUE30I54V4/fcKkNEWSAPn4OEzksAO80MM7dWpRu6n3twRTLV3GzjvVcB86I
/X/X54I0I65aWy9HIQyOgTZWEhx6EmRcR7ZTlTLy1hfDVRdWtCtugjXY5yMVwo5Fqx1dP04IG1iI
XmnBj+vD92f2QtAEAnhSlX5glIERIeGBJQ41dhcwgV/ZJ0GwZEQQk4kR/62r8AbBmDxZdECtYP97
Jy5OTGF9VlcpJgpRrbrM1u0MlNWnrZCfAptqMtHvJ640xnJC8SfO3Xy7LclkRakw91D6i8dzqRbG
K9pc/G7QiziYTPhl0CjFzYZEs90DAuk6HPZRbvcryJPbjRi7duXRLrSnLwBYrkqd04OZr6jQbhv2
tLr9HIDLcH4ukruqbqywwRLFaUOrQdNHyki8gJISVoMEmmXyNphnRuBH6VJotaw0PAR9NJ9mG76k
SePSPhWVFbGDe8blQzYGhKoXNGD2/8Y/faDZu6Z0adH+9HQxqxY4Ptaa45rPEQ87O3XPz/iKPEuZ
kAr6uBUUgykStmfMFjbfOQEC5q26IXU2OPJBPxMXFot4fqhniNp1pOIhhsghHeONZYOqCbbzXw6Y
wQwJAN/BGSlxxN1NLQmsaqMYw4VI44c9OWaDV8wtOzxAuWL5pMjOLDTW+gdTyvWQEtzHdGySns3V
fmEeEit+BGdxduIyWYj27RfjcAKfZd4FnaMSHeN7QJvIBq/eWOukvpgNOwIr4aHO+7a3KrPGk44m
YqUZeU0rmMrCc+8vesZfNJq2gqNwRmdu0GZvPVYGNh+ig+aMD8d++sMAdq9OcSTg0DT0imAokK/w
q5mZvO+2boxlsvIdJAXV/0Qxd8wJuatIBRWJ8TjHWOaFsZEQcubLxxjJ0gCjce6N5m3bUBE1GFVX
yXIRbeI/WsS2DeiJj712Y6utnn6cDYUfIvrz9hCfTt0IB8CDPfT3dWQY2cQqoOM/bq8cf4xIgIfH
fIOV/kWflMaOv4tguIJ5DbjYOnd+2wCe3xX+qzvolDqmxuZ6JlLcScAwMtA7A2tWgL+pCFkZyfHQ
Wxese5OWmMmq32qBr1/CRSTckN25icHjAp8rj5hBqL1o5L4tW0apayuHR21vRi9+Bmw77edH6wVF
8GLdwE33pBCScwicLw0tehIRggkvcRcbn5CD+PFiPb8zy+jVbmM/wS3aLy2IBKs7HqpEt9Ch2Eql
dT4TFu1s8gzMWvbB8nFZ+QbWJkkF+qWKtJzYDlBIILd90yCMEZ26L0lkK56oxr4dA6oLOfh69U8Y
Tm+nPVl6Qe2oETrpHklqvYNxTFGqO7z1kMGzs4ttBIGRY3VW9mhJZBOuOjJ0dTY/GVWyro4qnNR6
U4m325n8rYYfINq3yYe4G9z0gBfCgQ0P0XSRRQi6GKlxjzHJysc5MsyuNbUi5Hsruq44InBym6le
bY0v5GIshsfPLoDpKgOO2cLaZz7BENn+tE/pf3o7UDMkYcQYmPfTTyqCWTq9kh08I3LEy83dYMcK
Lg85Z4ZO2FnLEFZ1NemmqV+1QKnyeJcuh8cj9ErD9canWCglpctXRXGuxxHd6M1bFhJ5E3jLOAw0
cQzSNGGg6Ke3jhGOGcd9l2k+/HEmdbeajRYaGlD6dcPFF9ocqHQaoP4wVSPp5+jZ0jWgCB+exufp
r1C/RvsKniTJrtsW6DWJv4ynrY9QvTNgGQPQvIP2NTYKu+0/oeg7zmdWwwsbtrDKy5eed0cl5uCA
zQNjpkvr00Dfp6+kepq4N0X9LrdiUvRsPIW37ATKaTSfeGv4jtDvfFK9HW5IyNvQTA3UbvWmLpco
cooRb3tqNRHgfWBt6L/ZcVRTb2b/Lg3VSVazJgCEpQ2stvuKGTYn0XzN6GL+WVb8tRlXBebP/5Jp
bTxd6gQ/Cfk++P5ngN2KZGFcAIkMoBzfVBWZhGybgofMleMAhZ6UJ6gOGNNMP+kpZ5XGDdBbB/xY
k02H4l+MD0XGunIXRLFxrT4iZc+yMEWPItUufRa/wk/gYodZm8xWJ4HPcCeBqjd17TORnQvBwqLk
5CtitLnPpKqwJEbDm0iUv5EWtOcU4xs/BC0qrNUpMN4aJjqdW5g0q75SijFwHhB/PeVCwoiDsR2n
VbOQ9YbzU3X2Xn8sNtP8y75EF3VCQYdG5c9mvtZf2gtfdRncPBTTGZw9ZAec4PTckjJvsjsx76+V
0X4RWsLyv1bV/SYbdt/Q9NCocarKxu38yORfH1HlbnNkYlgM7dAG2FtOpTgb6D+QtmiYA3d7ivzX
vWJtvK1F7GBp+0alPMWLfB9hzRuM9G/TCsRMwAJuoXmxK1C7eCrpjctSvHczxwv7On24vVAn1sss
QJf3BLUPLVqg23MHk9y7zNvM2Io8DaMhS0LntcSXtU4fuT0jEYMnCWVsZ/Wrt0vmqxLD21ikWJmc
s4eI+obZIDA5YPk/BpF6zKKdbE9BaI1bRCsb6VfxXg1CYXKU5u063BgKOPJUakHPW2WXOkHHiRna
Wt+DL8b/1wJAuk9QMTmPddIapYxkCccmHl6UvaE+rnDpR4d4AHsXQLWmAfzGl4JayPq//W3AnWUb
9X4jARZRqhvRb9hcniMQSab5uIo/zzRp3iamcGLxAMZEHdtDpBSUFLmldv+Z7Hkd2nBnXj0BSv4v
wriT52rvjAEMGfwGytBrivHm8zgmlUBcnOQjVgNGm51v2/3U0wEBG4VyJbNWAYlZdMu1/hQG9GS0
qBuCAySLq3JsF/ahl+a/DGpQWEJm1yGP4wuBqTPe0geNWS2ym9wHYr1M3D7M0UutOAG59zetDK1E
FjzgPk89p80Rsd9cO9UQU8Px5rXNUlgP3zD9R8Q76tWoNFY7JtFm1bMHItPZCUwVuPWm+oeD7UvL
4FxkNQKkCKiJVlbIFE9BVN1/YCXII/D4nwC89coewGYxJgxM9+FfEdQM+zYzezH2TZOwTMeQVM+I
reQ5neeb+AvfvWtNmlxnIR7hZdwdf7xKcP5BJpgDTZjb1X8zPoWROJk41A4vNXIlH6v7ETGmQmme
nJO73JCyMLQygJjGcfkzglKblGr+sp8hb+CAZwEBUy/pC1uQqpnYxPOG55Y8KUmbhCfxVI8dZr+Z
o5hRR8YAzMGRWbGyhDv3FwSIvfrDCDBgGr4e4II/yjglFXm6HEXAek3CIPtwsFEvtrvwJsPa0CkA
cHdZ84k0mOyUgnXzD+sfwAgFRCVMgFsWJssMHk9Bu+y/JA/S4hwm8q3I+KbhktpIHHyLTew7r08Q
NrDe1GVUAdSJRpRVLDHF37kqJrrZJxfef6vcIuwhPvwNU7CEF6tI7p7HwTH8x/BRduVXTTHs6W4C
HZ3+aupHfgb+OimtXaZAaxvti6in7dw2GWLHh2Uqco0VZncKpWcXHz2hUoM7A34WDpb3e8dhMwcU
LaR0wB1ucubbS3fRxHn4ShZkeaf3md3aflyuvkHF45BdmU+ZUQHW7XbM/ApTJEJVFpjUDIM/7KEQ
NYweLMaZcdLPkrjqIwRQJ7ZEIGVI9O/f3/VriaC6LsRla83V6zPJDPAuwB74seLmTqPea8A2KvNo
11SGSUa4C3XMH/9S2z4m/BEBG9GFsB3tc5FhNfbjZNMOH1qbfML13s+0oy1KpqfgYa3F7pfe5BY3
Yyw9m5gQbk6kbpquudLwEgUgvj9y4EoLUiivVxiwCw/bQ+Nu5X/ow4RFG4C6JdsoHuIsUcc0tBmI
FQVGMmGckKiFzPCalp2iQio2KFgB/W49ylDwAer+5aNaNVL/doLSXTLQZJrwuJeY3tAnZc9sAxAi
pD9KmVc61/sM1SSyzp+CXoJJ+JISO1U0zG1d5D/mPlGXjI+TtUA1Mf4+GLc3R5uxiGfe3/xACsT4
9e2pnzQ8IPRmyy6ikAGY081IX4epQMk/yCxak6gZpXKHdcCVhivqjSKbSlOfESNDLjlzkPYZdiSr
WkX9t/Y8B7aixiTj2hwMU41hl+Gc8OKHpSkpSR728eXjl5PGEvsN0byZSZzSWm6Fyx6FNWhQBkNl
BCyUx5we00DkLJ+hO/7Oy1QQawHdJHDg7iizKtzAFcqyO9JGPzcF0AS1tA/4nOr83aJxTdaHtzF1
y49TviAkeJKOyG1XtmaGOeZE2Sd/zrMQ8Kja3uPJVlUV6pbPxQk7+FdezLYJh1d+bVtbSqO6EDOd
KytV7FWDV47zeWNKMn22WiKzFLE7LyNCl0TqjeD8y/gMqnKrg3zRI8/KAt6+D3YQg8U3PR8c4mOF
wja4ZtIcZCK+gewRZwiUXmcPJUR9/xTuBSY5Pkohadkx5I/68Tl2R83vqxuVoj2XVHjyIEBRRMzn
4nzLVkmwHY2WPcg5DtulWlDXtxLSQbqtQtNXWo9BxYQgHsDIndN1K/ePcxSZMqv66ITi0oOUQrZH
IzlSewnConpEGBX3fuwpY4G0B7yrfvtVPnVzqLiqIhRGD31i4Ao1nGRDYStzsLOAFEXeS2F+lq+G
3teyfJQHnV4RLtymrbGV9TbRbjsVPrDSZxBcGe6DSLqp7HzpsylS3nvGKVcKNlCCpIa1sqCYs5IH
Zp7GZKg5AS5Cg6KLYhcWixor3Jbt5YkhXXAp8o1WwYCohfMUZ9y6tXQD6NYa8S0RqOfqnHSagxZE
oCXYRdfHJpSUQ23ngTnd/YDD2zOFC/RqOmXso5PI+vvqFXmIc94Vu1j5DyL4lEhdzgJz+EfLpc1L
aoQ2Y9pQY7C8tjvZVsSeYbp+emtKi1/XT1VCRcrAKox+ol94asG5fwQLpwVTyGuNnU2cc36u3nVq
JGdHk11uKsBxtUYFhIqwEo6bbzdFlE8l1LpPNLMBORTBnk4GRRPeOaGvDHbfRxdRr+ayKt7pm9Qf
zf8cdB0IWGA9VZ/6e/VQHK4defEVkOUeEvFB87dg9SJb3nBjEbJj0lfSfD74VbC33tBeXRR5Ufnd
wr/keUv5fjRcbNds0AqdHWNo9OWglMsoS2wR51tI9dnI6gzhRIi2JpUMdAIO+EXHj7xe/Yfa302O
uWWWo2K+s5z/Grep/th3N5+BaCL9u5smze+d4bQ8J+8qC3dfiK1kcX6UFRxxlMnOqsQE+rbBGAOS
BpTZu8wpNaSJGS9Iy8SIhcZcwdHe6rE6/Zlk5DuI416l/T6JldPuvAz7BOTffVok2RVgbdL/fGGA
Fufn5Oxs3Tv2yUO+8x17RHU5DalbCGr0c0kNso+js6hJnhVocRYA9p3ip3IUi/rfuAfjtzncrmZ/
zkSFbddKmmWW/SQ044AFipxSTeEfFyO1hD5JtJ3QRKhVY0Sz2s+AGqHiVwSbomk4F8YeLNNnADq8
zN9TVbGFLFljz3bntPsYipDvDzY4Of7fScGcek50+F0xYseMrjMGBwMLA13MQc5cbZ4HoKnnJa9L
O+0SWLY5rZODjJiZHRKkJy9ZlQP3Fq1yiemqvenk8XHaalozY4iylzt+A3H8X88awi2y474EKisY
WBGxeSTJa83CrCFLC2jjMzYWdhD/RZVA7TnswTluxjvvBxnFm9wuKT+JCJgnT5ErhUFlR5+8evZj
W/dAodHOsi4rieT5/EyK4ppurmnOzaGXYUpfnpQ9UQa8esbkf9ch4dUChyvLB8Vr9IpR9zj/h8GK
d8YfEnJ0z71oZBtKHyW5uvgyzqH4CVAJdGisH+AJqhV6neV7iKrl3kSfUbpF1G55wM+C42ChAtCm
w/pdkTW1kcULW2ZGTbfCyIFz6waTG5EWAMuwzAIm7Vj6z6RVw7MHGRiIFdWzaPhVagsbjaUdJcZ4
FePYJvXuvwewKMwOyPDXsITzepEIh0e+CvWKiA112GVCIRRWORVfk+FgzxkyiizjV6aIImrz/eWW
fsg27asvlyTumM4cbyuoQNsMHccoydlrK+MxW5yZbGYSAtcR1Gu+sUnF7GkAWaZCIRxraOPwgvnE
Ko60PJsYnP35hng76j4zxOySurrzhM5AgA0cPJFOYmg6OmZIGzjXWd2h+BwzVI2lCnUGq+NUSzFH
t7XoS4Cd53oNB53hrO+DI3AT2ucZikmE+A/IYZ5av5lL4zjnIzHEZBwIS2BAXDfSRlfKVtm7ueUR
/GSNQFakqkmX6ElpHjh7hwMUBY85nKkTwy7tTPzs4rbcgnfRO+KE2Rup/WnO+3+ntElwVcvqwZR8
9m+rPuY0BtORh86B/MBuZbLdvzQfC4kTsYAWbTR8nZzFdxBWfV9m0KDhu/vZVGVzdd++Y+zymtF0
oqn7k6rS/TEtEe3+FOWEjdA8aIwSsX/PKrYg9C7ENiePGZ3Sk+w9opxjrBt3FVzB7m/eNYtJWekm
Mqe/+O70L3r3UpnlEJt1wOAjnh/S+EsM0gnABsnDmIA8dE9kP1nGMOsOS5mT12H0Xv+GmdrmaaJQ
C2t3Q9v/d9v3NayR53fSNucUWPOuCS9H1ouFetIZ3YmYZZNLFdqtUup2gNzULa13l4zpEQfFXlFx
4s7puHjuSnrlFjx/oUbU3p/h1vP+E9ZgCKBzSGMCG1buQ58Oq/xyKMx4QIoZjcQIjwtdZbVpW/A+
G9+7KpDSdtPiPnnALXqD0dsYCm9dVPHYR+hyjnr/XoaY2r3hsxAnJ9dK1fOA1ND0k5K2xPPzYOKK
nCR8OkjM//3dQQSXRYYkmJ63ug8vATgI90jgt4XwXOG3oUgEA/9vi0kMP4nzC2TKu03wqVmyq2lY
eocWa3Ji4YBouPPzjgwKnyWFqgHYY5u9s3hRoFPfZqffptWxOpQaTfd0/O1iIfbWeRdwzPjx9Wz0
Ww2AubtPadGO6KQnyKnrNNCeCl8ZX9mbSgwn58MRckGh+BcBxWllNMADDSEU0EvTcBcYQXmx4k7i
J7uBb5axhlmhXUHmog4Qto3yn0ltXDaYB0BdYgjUUFWVk3GWXGOKYNbQzNs1MpPXH6ljZ4J7GZtM
ar+bZTeBWS7eBNOl/f3Co3qBf89WLrBVXjWDKG/S1ey5tJOwqnxa/gYcZDkv6svxjbmpIVnitsnh
VJ8QpVYcAo99XF2y84Ipw4AFecR+iPaDCQgemrksXnLHWESqFznszcWnNACPhbOtwlsXMqVAMo+H
WAMqR+brzJ8wAfb9V3sfW4DsJWdGONEYwt7OGQcyAYyVtryo9yvN4I+iycpHztxAMCM6uANqem8S
V11prRV+H5976lDlmvW5P8W8Gd5cr7ajOzmXXzOXdvlIMjacSjvptn0gVZsKc94oeTgKApTp5axv
sP0FnBpNy1pcK0zcpUZnKZWTdozGTiZ6wcF2SIBpaT88CD5WS5EzVHUtQwW3+kRywDFnJEH/F2um
+KmEEFsfSXOU27KMyToyvw0QLaYKJm5TONyYQsEGyuuv/g9ZWFWbspjnMecNaSh1cmJ2kVr5rGzR
xkl1QccgF6qNEQkF35JN6nt1p5Eg1zKht9qr/N36y+arGVF2NMKOd8q4oXz2xzJwhTR1Iu3uMz7H
EfpgcCLiDKrlYeBPhpWQnJt6yLhgIFC77pJfeAC0HeJWLfGVaLqJPPd+jPd65RRHSVnPtOgU4MRl
8MBgUxK7YtOdAVVfWT1r2QfYPPzbfoUOiCUQ5FGxw2e0t7Zkn6M0Hz7zIyjiT5saOUDggMm7EDE4
pjy/FvrgKH6kJWzcyvl0btPU/RiGpR7zBQi+wDgMf9p6v15+eQ5VjNlVfF8sXYyYiURpm2K22aV9
zubVaPJUFo+GJ2+Xw5CVNxNvm2+jXd0/IsTKIWc4A6ljDlnvMwdE4AX2RmGGSWCPn3i5WPm4XiWu
IlJltCRRFEKC0RPxOUTzd+wzt0MIVC54GbqY+IuT4QkeK5sb56MyD4o5toP0Pq7X0Qs85t0nJ8af
YF6yJ4a8oBERjduX0Tm/xkTJv3oVBur8ow697xZEE8yzKhB6lKmVUluth6cCN/jYAlSiBmHuwIOo
zYGiqj467HJomBJ72/Ntqh3zy0LoDFRkfhjv3RghZZZYrcM9eOuF3FfBs1UX3tF+dgto3Iv5aqA5
42ZWc35nhPheAbfZsEe10mAzZ+Gf/UrvoV/wmqmGg0FF0sTmaQn3ncFdZkBlxAPHoPETzOmXFzmp
A6gXS111vZ3UoGm6+WhRR7I1Ft2EzFWZ05H4Im1X8LfMREHgYJN6ufTRk/Y9c9LO7/hMR6HVIUSX
gnV+ubdfaVV/rFl3duyskFhVw3ZsC918oghOK66zLWN5cKBXsgwRhpJfgwdhmUqt4RhBR60wbXJU
1ULoMouweGqEJjJB6ZpKmNIz4zqIHUESFULux5D3ZlypTwUrkJ3w4dmmPZQxN2n5BDY7+QQTyZeH
FPKrMxzsgQXBwOnrnW0/RHxnicYZaTsq6Pzo3BIca/wU5RFqRpBd46yYUkltISzM6NTC0rJ2/Vai
QuViX81OwIc+Wyvtn7tR0xQB5NGABZnoKs5btpmTffryPwai2MH3yZDcuoTO7L7XkThcbWeNW6vS
h3m3/RapYMAMdrqS+lN+JzUyUdJfbQlof209ANQyyHS4kWEAmFKMgMPMbGtCVLADsSSfR093CHzs
prSUtLuJBMGanj+HWafOKMfsKgPxW8RkFwy/9gULBx17XJ0AtuYpGQ/g93dVh3C42/Btg+PvUTKD
mjmrmg2EjoIAmL9E1eYYoiMGgSQtizk1CztnjhVITKGWI+lNwW7XBpLvoePvlaIF0GDjTFn33YGp
FKfpvlKOa0RcwRA/2lgavgx75QsIAzjw1LHqmIfm3oCH21VE8Ty2bLZtbWkABxvUK7M55/r0adOC
jSPWkzF/GxF4wMmvpjdbIKdsXsl/3/zrivg5E1VhbcajlGgxESQebrcW3kyVEi7yT+T3+B4Ekcib
AKg+Kbicj+d0s9yMfAHBZkRB908NJXewytGDcqbTGGaFrvIFnu9Ch1N6LlU1SyRS8vFsLgIILEqT
quSHkTTMxyll7gpFwWbTBFL3ceLiKzM97hoXGShnlMtisOmU0XguG7ZUBp2Dv7qJmik8EZTdN3Z9
fv5yFd8cJMoP9VifZwEWZCA/qAZeorzw5YDUI/3DKMxhoLkdPxRbGMG563I8LZ49lQvojUKsYfpZ
GRU8+4CX6/WCj9oj/ROJjTkjozDCpVK4PsN7XtqV1hE8myMLCqpWBs+WJ3OwASoo95tITMLUhQDL
a6pgodQXllvKZ8rCfSDyml45xdT40jxfFsT40CaMtM+EI5p97dzhk8n8Bh18Em8hiTa2ZrcPY6qE
nS0/poRkQ21tzu5XIYqZsbuNYqHcPDg7Oig+cs3R341OQlc23igNLD5TWDV4mLdUn/ogJFlk73km
KE19W6GWudi3BDGpLRU2Zk8qXvD3lrRqyTsEwY6/sf8nx0Z0iDRKzLuf/qPFKM8d7ZuGiMynuYOn
7n4Qvblukt8Fa4H/Y5rJJT96jzjeIB6Qo4UpO8JarEgRJEyefDgJkB9zxShMhwJ0U28lWjrli8pp
a/Ys2zgza01tkkkbf33pvDp0Cys0yi+YyGo+mdTmO9kNg+pWSOyqZGgnehWZht5b9OMj9JUnRpzQ
utm8hqI/HjckwGmzzNu3TNIjaRn3cUtiXDX7JLxP34/C+aAy9FW1AUKvRznXGdryiUqqgcmX73C6
Lkgl6LVv1+J+wvQ6n+7iX22UB9/NmiBQu1lkZDwK1EaYgZY5MIRmP7G+LXLGGVrRRd9+fb/s668m
+9mMR199Vutyj2DzFeMbKxb3ri8QsFeXjp3+46yf+HatjHui3cPuB1OyTP0NRR7mnnx/TZHGDT2r
W1IlNJd+d/PtjVq2Xi62vsBX0bNRgVcHpdCTc2L1OZw3+tpE5Hdt8yT6iG9RTFpfnsnNpA9rBYqM
01JtLpGBdqe/RyVsSX6B+l0ouNM71CzGZcEHt1jfWLiBxkFNtLc4x4if64moKtBCOVS6zaHP0Tcj
02J2LAB1/KVMF7gfLkAq8W19RGmgCAuA84H9s4S9xdKeJhVMe4AzumVASfd38h06c9XQrhaJlJ3e
jFeHIlm9lXuBALAnzxVS/wZ2rPZhb3S3gs7CxwF/EjE0imfw5O7wsM4CDT36P4YmE+CerpqHcw0M
Br33yePDprO8fmTk542yhuejKIYvRXPn1LG2wNYxBBFW6ShMaLdMIoxG/axpxuu2ely10XQWrBKG
s2HLWjhdmKxLlsT1UqIQrRpLli70MTe6Vy/oqaeaN83sRgMnf5AQCU/+ffwIHXuhEmbLpmn4tmBs
7bfR1o/exhL5XdzJ3+zv+GPq6ySExtGolMEdAdHrAmyQk4odPgcrmueprNHkp/4FyUDEuGmC1Dza
Gt8mcVS50KMCvm5qaMWNNxWFl0vKDE2cJoalibB+YUE8cGSj1Oe/+U09htx8ywJE036VHr1d7TN5
A7ROSQ5Ld0Xqe8hHWrgJnHkyLDtD9KVNU2+ElV52YW5b2eNUQky5jLXWSRoFX9vIhkLhWkqoS9EB
OVBpGjRiR11ul59e0+4hVCi8BxcHE9JQhw1M6b8TOKgpeyrFx7UgV4nc2scKFz58gQj6abFg3its
J6MnZqovi6abe2sP16VhLJ/nN2rgYnmnzTsNCMr7njjfvi+sBosW77QQ/MyGfJwQpYS1miVLHUpF
x+/qZFpN9X/LVDWFSjONG8FykCkF2f9jyYjnAIEJdEvNfXFlzl3zO1xSXyNp73sRcHaDJUNfC/Rm
t82zGI7pTYSMk3oO9CUKTF2B6lq5e5HNCND6/s7Zgfugv5B03Df2IAnF6Lu6XLSO7Ooxh4qgAtd5
Y5g8efafRXWTaGo0qIbm2xXh3XVX3a6jk5aABX4b+s0QFKY4XxzHZVEDP+oJCqL5jcrUZICBOD5e
ZenPwh4NrtYLdGpmtUXJQGUyXCBy6BHYkb/SBMKSB021zmmNktUbKp6ASM/vYN1kt+ZFJNmFt5eE
hlOy5slcPeNTb1VjXWsltKzKG4F4MLy37h/+qZkTL9Sf1kr8lpH8rhlL6akLt05GScU3xKYO1hBn
0FbVhRPwOHqdXDGS9p18MyStWh7BWa/YGpjyAya+RvY7TrUcbNQUXkyHxYCfFO+xD3pzeNi4LF2o
cF/wEd9T4GHGG+LrN9PrL2izGR9MC3CHGRyMPlFVZPT+ZBFzKXiJ/Wckmy1uLJtVNaRIk4VfkOD4
WGpZxLjJ8Lv6pHW49RfHWoJrWLeFtSN62LlXrFnRnijEq1I4donUgIoN1HyUoCahidxVXPqxsYgV
EJ3mjZrW381mJr3JGiuROIHyedDWcxFS0W27EBiF/U3zERUEpGMBI/PW7+89NvVLqhDen0i16Y06
wOMIkXd0a7DmLvrPoTaj5BX/LLX6a2Iy7ZpBc+m11tVXqQDkSQb9nvlf3Y2kenfSp+T7YIELw/hy
N6yy0X8SD5prGhABMjwboj9kjDL8VJv8AAV3c+MvfPGtUSgVah8x9pur6mnprtsOfL6GsvqcrV6t
Ugb4+G+Bhh48bfS65GqMqn8+4pC1UDHMCFYYthO94+RBBsoPyAdXbvcx2I9Ve6ec6zjve6LmIF+S
5MYiBkIzTN3W5R3lXydi+4bo8xEpYd2hinSZ3NA10RF0gfWOQwZbTRzBfxBKjgqgy8wk58H3BF3C
d1+KlVZcahAPpgAHBHken3n4eKSUg3ex4NAl5WFk4Sj9hh/PtbmBE5M69mi0/K2PLEITQjcV2TlL
7ETvc+jsmNNPZtk+EVkipmAs4kYqxdJ5XPy48YHbVoXvhHSjJGbNt0VPKHwRozHwaXX4T+eqRmUU
/pNpnh6VdiFk+f9ZZcGXYEVRQ3PCrobMGUuK9+BRen4L9JvpwpaxewIS+KdtbQP3KPuhrpPsSTyb
mdBzJdY295yJFT7JoimmCRN+NtYYPkkd09/sHmwU0awnlU1QPq2CRJ5FbqEnRQIp+guDe7ovagjG
uCZpiiI/hbfZXabD7CaGLJE2k3sY34UdMt3+fxWaY6u1WgCMXwXhPxmISlvWqqRaCWSpjProBxoC
J+yMG42Hqh4nytybInyOP86e72vYxHwHyjOCXu8z06ZyjU9XMulDJbZIPtzVKWLc42zCua1bp0+a
Kzuy0scb6lrYkGh53FKSB/9Pj59Ry2Y6HLP/T+k0bGwriiaz9Aie24e7pUSM8UKSyNpDJEkYA/fR
tj8yKjOeVn8NADcX2SfRC1JPUJZX3sHnESVbnPukfdUJsuqk6nsIZXfgit+r40at6Q+4bC5wcF6V
/oeGME/Bcw/7DKOmCGx2bKs2MzyAXK2HF/iAltTiOLnc0TsLW1r3adISfr8MLXyabTQfHCkLInY1
WyXgcnIXhDuj6iiVPuvFIdvfYotApbiE4Hs2CkmE5CP0SBsPlEYcQC7owQSzQ5n6gO04asGQMxJh
PWSBeCeVyNMyWX496zkug5ikYNU4rrkq6vZenCfzKw+JYdCkOZoAE7A1/qGmqJEI2/iFq6EdcsgT
zfsrorrwcCzrzWtlOj/f0GVDI+1Z8p47ymNMBNtkZ/fBAniMjRBo8qEUhnY849NcUAz5SLVu+UAx
LF0aDcmdnyobqLsFvjyUKvF/16SlTYOP1AJkgPgzRUuy9lLbPRQwvLIUCqMR7CenzJwW6fbcz0K5
6Ywm5B9/gLBbNQeXNNIpUZ8uFrYgGaUEFKnXo0kxT+xib3bc8Z2rMcISrh8tOOTWGDsablhquq9d
WH0PqWgNrzGpIzRKSQoK1jXV0n2y++PAZe53NqrljlJdJW1mkGKOPXrfl3EYuxH81I/jouMjw6CP
heLx3BiLsH8FJ+UIP1GMShlB8den6ygPmfoz8XxpWCUVHTw7KbcUuW4myr0trA0ewM//YmdbToyT
4NACEM817LVzfDVm9CnQjXqCd9u6TGL+4+IzpEhe8G7gqpb/SDwFRA+s1oxEs6/IqFR4t9U2JL7Y
ksIwpv2JAddyQuPM+pLoAUWjZKSH4JNqccr1IGJ++VcZVuikBRwgNe5jG5geMmvjNd6o4hSF43hK
BBn3UapEZz2+Cq70k/iyiqhipO8hJ1Hix6t3hFxbfCm/G6/RwKrXIoPwrnWlUXsR7c9gRs1kMZqG
tTDqsZDx/01HEe/cwy/7zFowQapeW/4NFIbCRfqPMOKsG57U9D/SN7P2n278Jm6chXrFI9Cjv1Ox
8TenExGe3+uH+sNXl6xYvtgjeoP1HAgkcHS3rMAkrbhFGPP91ltUM3vK8/WylneIBqnDSECntyvH
E/isYISbSp4mJNSVcqeaDjHCdAYMQLKLwDfE+rsKAT7OXkji3sRk08eYoiq+DK+elEsj58+1Zyer
Gu4IRZVqmKkIEEHL22ZA15ftapDg4Mh3fzo0A+NyA69zNg0H+FIyK/M0eb9doMXWw/Hfg36VYUil
1pIrfTrSSOacLHP+mY/LfZPJE/IeEOo93w2XEptnQsLjdEZwiUgYl5yP6VM0OMuzxKmtls5LJQN+
5klRJRhpx9ie5cbJ1BocpoQtjo4sZ1kcP0hKYZXGkSzDMZhsVv+8sGBYR/J7dEKQmGvxg3/uLLBZ
F1M36naTw43ZfjlWa8C8sVo32m3nFx8PGDJl0muhKq4R5WzuPqm8mHFr2e/MvrNdbeiJ7ixfZw0+
o0l34A+kcBNvfK1sWW8NZ5zPerH9+bkCyr5jxuvWlM5y09K0Vvw/IZswEkIlnuwnYEFeGR4gs4gZ
OW84I73cYanqjCZT/JRaUtHjSU8Ix4gUsvGwXrXT8zAtnRyQi8GA1m2DheMr1wKgszHDDE4P/PQ4
4Ohjq73PsiTwkD9LvrgWDB3ZmlgpvSQBpP5xCJNMItrYnrEMQAq2b377lh66UYWfl3zFz6Lmeg9x
KZaMXLD7VG0PpwOjIu457KlbORl8drHfB27GgKj03VfwZSI44HzSrKpj/zTpG6uAQIRPOZ2DuKQ7
YCncoOM1Jy+N64yK1GMQqO0XdC9mMOnsei59AAVF+iS+ob+gV+KKDZMX5NxD0n0x6N862yeiXNiq
8XfbyzSfTB4yH43L62S0gCgIUWnV5ueMc6fSifQ2OhXxUGVJFWJSG2iOmjQN5E6wdnkxkzV+7boO
mF3GYBryUpoCjoqGiV8tYPMvVgxlb9z+p9Cqpe9Lc6QSV05uxhhLEOWsvscN6dPYEYME/o3dTnwH
rb9+/hpX2Nu0D7cHsl+97+XzU1L8NYmyS1opTJXZrYUuc15J+96AT6Mbg32YVsxjLI975PgJTwga
8lNz/hNkBZ0kZ8sCaSLuJ5CRIAZ/Mwu47NFr1gtb23UlMerdO8y0KuB6kd6IhMflFYKCgcO2EJ6b
fSz2aUclIoITkvCw7bJfpJebPZPZfd0jh7BMFbm/ATrUrrBacYzzoROlMMsG4cjVovMuV1WmkXbV
/u8M7ao4ydNCKUj6yGdmsgWBXOyM2PmHzWyWaSlrIUFBFL9r5pF6YG8rdXIWKuXrXWt7G+BMm14z
GKiYEflIhYA3vO+M2dY+mPN/yyXUOJ7hdZW8y4ONeiRvNdXV0du8ukz1LBfp23os0G4J2zDK+LGx
4+LaGtLKjQhBGbKhzVcIKM79f3bjQFahXqiDnNReeNidv/tEOrM6RBSfN2Mx6YbUVzOrqWKC28h+
Y4L9aDwuRQ1w1T5/dHI5l8cooi6HS9x7nLn6Pmv7XUZS3zFXkx2sMc2UNyRtnxxAL0BCw4yDnBnC
8CqCu9kHaEK710HjANK4pJmaRQ6crEBNZx63Ft/i5Wkq0aM+E26tkQthwxq+lFlt67TitA1fhTuD
rhjsDdTXufbsxoHLm+v8Oe0WpmafrfgGzTmKNaLfVoXBhmgRhtM2ksSJzybeN6ujQdNRYYnl2LCR
GxSjJ9Z6zArKh7Wcr9r/wF6ScmYvAbajwpQ3Ws0anyh05rUGWPMTt20pvH1vFqMDfuOSHjYq013d
NhtQJHSnMRsOP7Azg5+XnREyKfs7Js0GFx5vUjtdq8txCgKowMpb31aQCnl20kAMAl95IjPEl301
O50NMHb3dhY2FZfRYJ41tqjNE9/Ed3CNxCTYxRWiHQHEY+/GiQDUEwZMyXz7RLh3auE58G2P85QA
5/3hfMZS/ZXvCBDDEB3WkJvIhuZxAr0f5//lgjFeks9w4lvmfdyKGtbEyrq6aIPJi3+SfjGOIBuK
P62tu9EfRBdccLOOT0n31POMnHOoL504+ORttC69VvXBWdhyZCYYRSO/YmFV/FDHnrfOVLH4RSxe
+kLoxL90tnzFE81C810w+/vPg8N/Ls7pY5YWgLaNIA9vT0Qn5RyrzlSrD/1CSW+qeyKk3+ehVgO9
gkq6qgTghEi0qAMqX6yVHp1oWS1XnaqDso/GrAohDX/m1HGbR8NN+FJWlVrEPW1wPsJGA3JR60LR
MKCmNEBNwMSAH1oGVqDeHzL7k9UFppCfN+fW4f+ae0U=
`protect end_protected
