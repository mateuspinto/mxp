XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��m��{^�k6�� F W��3}	����m��s͂��Iǟ7��f�]8��w�*i >��Oݗ�y�4L}u�zrrp��|����X9���6�1Y�� �����l��ā�0#Q�:�d�U�9�l����/F�,ݙs �h�*kָ�����(j�c�:,�W�Į		���י��Ed&�`T���0�x�x���!Dٱ���+�����ʃ�y�?��
���и]��ߕ�!�'�W:w�`o(�3p�7�~���Y�
:�4��Z.��]믗[˜�K�nӁ � ���=�p��{�>.��S���
���'ZP��$��@��P�hS���AT����t|�Ue�,0�VnD3c�{.�+�a�?�ȀU��~�jT`Z�H"0���k�1,l��e��k���Tv܎)RNM��#"��L��Q̭%�<�H��OM��؃�Ǣ@��@��A�D��f*�>a�!|+f�0�˼�J�M�,J�4�q�v:J�є6<a�{��(�k���d��2���4qo��߸b�'%�x�?L2g`�*�%[�e��a��b��
�*I6~ų�sk�h�˱�=�|�T��cJ��9�!ʽ�3f�Za���*c{Eq�ߎH5;��G׍�(�����:��.ph#���>"�( �pr���te�Ph�>z�ROj�	qv���{[�"��Ң��#��\�� #D��?��x�2�kVԐ~�Yc�m7�W��WO����{�7�E�>��%�i~XlxVHYEB     400     190�/��"K�����@��%�$H���؂��M��d�Il�,F� �h��2�|ې���;~NQ�U8�8�t�&_��C�h~vu���FlS�%�X$e2�I\G �7�ހ�"���:n���<��ؤ���w��=�2�ŗ��`�Ճ��/s��ɷ�s��+h�S�B����oIAB�fZT�e�>Q��M ����/�X4N�4�p|D{~)�=��x��L��$=�������N�)��{�O~��v׭+3Iڨoƾ��[{�7~i��B���١<��ڈ���N\ԕ��3}�!qhCp��6�7�ƃ��r$8ߜ�I�<���Y�J�ԏ?6F�iLd���������4�U#��e������V"��|)�N���o{���Zfr�XlxVHYEB     400     1504��J�V���R����Iua�' ��GKIk|��x
8��rO���U�r�.8����O��k?;6]=A��zp�@�T]E��؈��y��� �ɟ!�Y'�c���g��nV�"�{T�⋿6��m	t`� ���E���\Lę(��q����Nd��99�1.cQ���T��P~P��\߭�%p���Q��'=�Ӌ�dsw� �>ޕg�x3e�*���*�O��L�P\��t؃4>�\dW�秱�"��֍he�;7{�9�+��gD9el�B���F�~�m�v��tD�-?�q3$w��/�W���y��`5����tr����XlxVHYEB     400     140�$߀���K7� S���/17����M�����2q��W�Zf ��G	?e�Q&b�0��m�����%�������|��]\�+H�en�Gd�#�҂�gj(��G� �X��.^(�hE���p�OP_��-��*��̔�9C��r�\�����9
ʡt�	)1Ѫ�f� {L���~-fQw��5�W���rlD�L���Z`p���QX�o��x�Qg�<p[ZN��
�zݡ�^�/�.��ͅ�o�K'ą]�;j[�y�SD� T7��/ �~��/�� x�*�ݣ�Fn�� �]+v����bp�u��4XlxVHYEB     400     180fN�!��R��޹L"z�6�>lna;W�&3ܑ�_40���V)�rTA��s\�N��Qq��3�L"��eYy�ɜ�|�)��^)��&j����I*�ddN�ޭ����.%)�o�w�ܵ��jL��X>��F���}���r���#J�o�UQ^����F�L�&���Na|8\wE�ed����w��,@r���	�T��2���Q� �eĤ��B-Fq�b���9o9bχ��>�o�����1�)�Ł��ɨ����<��/`��������!��w��$���_�6�2�$�P�fz���jO?=�1�P��B�������j5<����H�_�Si���4��ѢU�����uDߥEy��X4����L��e|�XlxVHYEB     400      f0G��NS�S�H��a��}@�ng��2�-���eg!�ٌ�yI}c�h�zN�0�쩆
w�?���P?�bx��.���5[T�!�GZl[�KD�OՙU�Q���eGi�WK�ș	�^��]ح�{"������}3Y��@�XlT2e)��H���L)_�n���h4���cW04ؒ�Z�P����ŞoZ�`��]Ƨx�����:�"a����A׸\z���oWW�ǵ�����/�v]�wXlxVHYEB     400     150l�n_m����p�B��#�@X�7HR�~W�ځ��F{�+n��qz �>�׭ k��64��J��O�g�_�z�&�-��Vh/���=c0ʠC�?W�%a�K����t3��9l@����[ܷ�?zk�L���z&ꮌ��uVL@b�$�T'�w#����!�Dw:۵�%p-��v����C�߳}�A�۸L�A����ઍ�F2����Vʛs�/t.��fS���/��^���b�lD #*�&f��m��7fm�#pߏ6I�b,;6�t�/1���3������i��!V9�˭���1{y�J�����@9�*i����l[T��qSL	����nXlxVHYEB     400     150�j;�,'�c%�3�Ħ��Ҷ�?��{I������(��k㧊�)8RK�EW����JS2�EцE����~�mNU�xz 8ڹ;��+PM$z�O�M tr&��������Q�#�T~U�ԓ[��6�B/��������ZP��E�9u��'ʔP~<�q̜�~�sp� �4�]�F2{ЪK��U�d�?��(؝�(���cF�ُß)�F���*׀����<ub�n���͟j��x���dM%�z�W����lc�ͻ������$؞�;7��f���M��
g^J\�!Y��wW֩,���0���%����h4⹸�,ZXlxVHYEB     400      e0ug�K�Ǚ=��������B���D��I��^) %�	w'0Ȯ�[����}8�Wfz���4�*�6K�6kC��F�1%�g�kR/���4c��]ӡ�vF1�б[�"�{�����F}>b�PN 1+AJ�g���=ˣ�1͒����++sژ|�x��T�]뚌����1�j>�љ��OP�V�>���Z�Y�F���Ǉ��=V��)戍��$�zXlxVHYEB     400     180Z8G����V���>ǚ	���J�c�)��!�gA\�F�L���CBta,���SP���;���٬�J|�N/4�I�뼝�s�L`�t�Q�aL�`
�	F��EPg_}�s�e��V�]�ǽg��A+�a`�25��O*J5c�>>-[�!�u��h���������,�H8��d�T)��x(��L�M�ƾ���'m/��9C��T�+��.�\��5�4��$��L��J�'3�	�B��ڮ�R���im3@�U%�-[�e�D�\�G�+���v!��A�vv4D��)#��/�ӥ��cZ��|�8�?�{���@�V#t����9�ߣo�%�4���[��W�h�!���S$�W��Yi7_�LwrcUd�.�C���᳀v�XlxVHYEB     2f4     100ư���4Ā�fr�pm�#0�OG\��-J;�Bl�k���/�'.�A����(O���0h˱3ڔD��8;h{H�!���.���p͊b��Que���J�s`�*o�`7�h�O�&sʠ#���w���K��j�����8��e�T��=�7��sO��R����w���������#d�ذ&}$����/�!y<�;X�u���ECܟ=h�b��w�xk�XևO�}�<�����m�0�,��1_ߔ�S^I:�̕q<#�