XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���E�Ό��u�т	3J�F�!��5<�yv�zTBj��C ��A��2U5��4yp��n'�q�o2ϐU�݄0.�nV�H�1�u�+I�I����[g��X+�6W���j:W�9�� �J ����׽� �n\0I2n2�^���z�YM�>t#���S�f��B)j��}�,1"���b%�W����-~��=�(6m)�E�t�~l,�%WZ'C-�.��t规����TNVX������5H���!tg���O����e�[����I�7n/��+g`��E��ϥmK�t�Q���t�\�}�S�� #�b)@K���Lѿ	��o��[u�w<�
�7Z�?�����#C����H@�멫�L�	�lQ�55t/�^�RY�h�\���:�B��~�@����d	�uL�9#��E{�Pi���S0�Z�IA��C-�<xA�J��&��&iޢWvj%��H�y�J*\-�{R��-�38��̸�/S�vE��d����K�{D�S@G���
�|���6in�4�[�7VҘ�h��uNx�
ѯJBk� ��:�UH�w���]��y���b��o�DB���#G��OQ�ץ��Ih\9���*4HQ�k���@9m|����+��?Y�#���X�+����`�o��-Rr0�5�Ł��G'(��չ��i��҃�)�0�w$�rٕ��NQ�	�Ⱥ����/%�X�a'||��#�o�qD�F�FJk��Ag��+3�Per�z�s{��_q�m˭y��ٸ��SH�С���XlxVHYEB     400     1d0�&�{�??���U���'�:!��R1Xٱ�iڎ��h]-���r��h���8rW��!�{�f6������gb�p�ՆbQ�<�;��O�e�o�������O�Yh��Z�NK�V��_e��v����(��AP�"]2�ĝ�¹t��ٸ��o)�����MS!P�W9/�Fr��������y���D�Y�@���-�g�X�^uh	�G���\d��fc}�:BL����v���Y!
��p�z��"\eM^_m��`�aH�	?��l����_������bQ5�vIΆ_�c����h����K������ה '�'�N�:������Rp���o��RI�����x��k�.u[��NhM-�<r:��@�����3�+�k��.�]�A
!/��6��|M*E��D������~jG��%�����$ȳ4�����픾 j�&D�4XlxVHYEB     400     140/�%9W{��th���']���4�
63�nIB(�}?�����L2��2��ʃ˶�����I���3/?z�j�K��AM���=��@����Ք�Ksn)��><�6zp�7>C��C&��uP�i~ٌ�_D�Wg��v��F�'(b�&�'����JruΊ��%gk���*U����=�V��'�D�ڰ�<��"����m'*{�)���J#�
j�:�vO+�|D��a%1����X��Ê@�l���W0/�0��lt�g��4�
Т��A9�F:�A��p�q<���+n��`�oL.��[�N�V�jǣ�J\Ԗ��XlxVHYEB     400     170ws� c���T�*�X#G���2M�o�/�lY�5y�N��$-FƝ4��\�2�����B�=2^�gS���}��\xn���VG�@�uť��
Im��#^�oX ӸG�6�#'-_?`N�W�ݦs������M �ճ*!=��+�����T�����)J;�d��z���3��l:W����3]0^\�QDl��Y�B씴��;I.R� 2�(�}��Oܤ}x%������� D[����j�M�0LY�&7LU����H����*sym�w�ր1�Jat�L�p�'0���0�!�t6�8�;���
;����y�L�J�f�蔉�}|N�����4���N�:��5F��늢�_����XlxVHYEB     400     140	p��=n�)1��HLC�y���,����I�)�t�-�J��2L������Bu"�=�R�Q
�X�Nȃ
{��e��U0�3B(y��S?ts�<�j2�J0]�C�K�E���!�?�w0��z���k�OX��X٬�V:���1�n��oPf��Y�����n��IV���u�j00�4��uH�}��� b`qj�1	��
#[�#%���4 {�#�� ��,�'������/o�].�J��:���W���}���-��lm�S��`�ݰz"�	4Zε0��=
 K�A B:��}�4�Eo����'��k��poXlxVHYEB     400     110t�q�ְ��B���_p�j��'׀;���L~倽q1-�㢹~/�6{ɠ2z��I�@p������X�6�<�=�F�sR�;\!`��]'���@�C�`9��u|T\M�\��K?��jG�<�r&{�����P�Q�tDS����To"/Qp)UNw0LuZ�h��݅��.�К�j!�k>���!�~�	�-tU!��~vm�wŬ�@Os|8A@�"A'Є��y�(y\�0'kaGW=uY�
Ѵ���W����;�cA�[�L�+͞�0Ʀ�5�=��6DXlxVHYEB     400     120�*��q+�,5�#0������i�-��������d�,���B��������ޅS�0U��IQ���}�n��k����:j�I�#�����ItG�y�	���A���X�j�1g�A�$��>�]�聰����
�6�AR:W5�y++�����H�HY��*�'�z Fxrj�ق��zEr}��As���cĉu�97W����In�IRZZ�KN*����gv��>A�֖$ғ5:T_���"PP��BS��s��@"}��B��uX�$��fu��M;x�L 1��g;XlxVHYEB     400     140���F���gb�G�n�����1&��J�p������OP�1���3��I��� iFr��V�e���uĔ�r���'����c�riJ�J	��Y��E�°�i,� ��EKX~k�8�x�1Fo���7�ͼ�����2!��]�)��AFB�4ތ5��@��������"\%�ۿj�aRz��hIUX�K���Jڐ~@}�&-1�X(���������?w�:��;�W�Z�6t�,F��^�����)�Mn�r��*��G�>������jMY`�*g���.�� �<��	a�������Ry�i'0���F���XlxVHYEB     400     150��`�;f�L��7���: d{s�c��a���
�X
jS"e�sk��i��t�O�)�8֐ �~U(6�J�D�mϔ����@������?�����?�w��}�q�� {Te���u~��!�R?��$���N�����5=���I���;W�x��rL�a��0���r�.r�/����)�c�Bgƛؓ���f��XT���H���:�E?�����F��ȇn�&e��F"�kۻ�pۀ謆=���RA#*�ގĢsEVr��ࣇ������Ge�{�סּi�>��lg+
D�9�^T����Z�A�XlxVHYEB     400     140���b{G�D�?�>�eNd������{�Z�&9=;��^?�\b�ʥ������t<\~N$ �.g��]��|{�[���zD�U�PSr���^-At���!�+q_CRCg��q����Y'fXE}~�H�V9�C$���ȵ���,Y������0���9��\r�R�Ķ�]DU`,ߦ�-wX~3����א�g��o=��EB����uʍ�$+0����|��X*IB
��������-�ܪ.��>��J��kx���jd�gR�>!Hڹ-�Lۇ�.�NzU�Q��:�m�EW�}l?����rI)XlxVHYEB     400     100�-��\�ᰱ�?�^yA��:V�Q]��%��R��D�;�YVs�A�1����*jL�D>���k�װ"�N���z����P�t,��_��M��T;3Ze1r��eX��:h��L���?�zC�����ř��~|c���t!A,�P��WG��������H�E����K�H&��E�Rm׼:�j�^*\�,>�^�����?�_�q���-+ њ~���x��@�A�?��=�A�ex�XlxVHYEB     400      e0�6�D�O��9����I_�B�`�zz>W^�/ѕ���^}0]���F�!Z��ͭ��O�g�C�?�i+�F�A���MM���𶰣0y�wD
�p�,l�m����A���һ�7lr�%ѹĒ�r�Qc��$*�+�����D��`��B�C��$�"����Q'F���Y�/� �rc�;�f�Q���7Hܭ������ 2����?�՗i
�E@�����5��z��PGXlxVHYEB     400      e0:���H<Q�:�[L����D��O{zsN�_�Gid�@�p�^�0��Q�n'lG��H�5�{��G� �3xΆ*�IFO�G����H
�s���_o�-��=�F��yˍ��" .�C����V�x���';���.1U�M���dA=B� l�5�3��_Y��� �˞ĨpB�2��>g��~K]d1*�U8K�r��%AQw2���j���ϲ���K�XlxVHYEB     400      e03����ZW��3ˀ2z˛������[�V]�rz߳i�x5ķ�v��ʥ-�9!M\�.���k=8�*H|�Q{zbb��� :{M_dk�:O��Vo?���B���d1S���B�8A���/������|��<�?7G5IK�V4�I �*A����:�z�`�,�rŴ�JW�Nd)t����n�V�|�e�G<�r0�F�$�g��2�S�, �К�3�P��XlxVHYEB     400      e0��yl�a��$E�Y#��=��q���s�5eݐ���(�Pv*�p/�]��d���C"���i;hi�&�
7���-� �����~�/��gS�G�c�qk�4ҰP����͋$�?e���
���d��[���xT@�j��b��eN�0/��Wq�yM��+J鍉����j������]��,��~N PYS�=1��"��;T�Fu��~��(�4|��<�T�XlxVHYEB     400      e0�"����Ln3i�x�˰2�P���X�d"�g��u��8T��d����Q�S<�M�XGe7���1��u����������
��*s�O��-��(�H&F��[Xlj)V2`�">	�1l��0RҨ���A@w�5�vQ�9�^ئ/�Xg5����P_ʵR�gdp`xV>KP�Wm���O{��um�Ǩ��r��do��Ֆ��Lh��[�*3�f�T,��+��XlxVHYEB     400      e0Ab���5)4O��/�Q�I�ȼ��u���y�Mb���M]�&(;I����(�v�]l�%��,�!yҪ��gr��t��5��O��'o������A]x���[?��|�ww5����0e<З*}hT��F���j�IO/�LJO8����լ���L���;��T?�V7�Z����ߢ�ZE>�Y* l\H��JZz[.���k:3�co&�H�F�-���XlxVHYEB     400     1c0��	/���K��N���F�.�|E�9��$��;_:��}A
��!9-��2�3�V��㣫U���D�k/:_q�ȃF���DpM+y1�3��n��/?�}��k�srj�5 ��L�j��"�fKѯt�zƠ�:��Fa���P������m��˨O�m���-f�N��QC!ڗ`�>EC�h�43)��DG�rP2j��n�����G!6�	>&�F͞n�^tA���T�,Z�p�.o螲$���̴�j zܩ�����??
ԟ�[_~�ߵ!|�%��:)]�r���al���n��N�,� k� Q��y��p  Ҍ�$�[R��z?�%*[~yW�њ�B�SG���|�葡O��FG��3l���� J���i����F��l�Z��j���P$em�IAF����:.V�ל�!=�4D�XlxVHYEB     400     130�Vv���N��I�I�\��>.)� ��C�a�R]6��;`�f̗�u�:��ᳮ,���gD�{v^B�qcwU�h���E�Mo�K���2vƱd`717N���W���t/�C�u��j�.n�=�2��e�"Y��8�O�l�y� ��� �C-)���>iN@q��;�5
���Y�ԯnN�-ZQ�gL= �9ȱ�(�q~JDO�~�E�Č̨=�H��FTWĎ̉(����
C$�="�lb9�o��V-�){y�i1�̥d%�Fu�ԋ^8͘��Sl�=0K��XZ��g0<�	�	�8XlxVHYEB     400     100
���ޜ�t=� n�(	��a�`;�z�H���^���ENJ
Y2�
�3i�2��}����r�:T��ou��HZ�#�g���#b�?��MЖ��"�d�X)�����|�!�)K��$�B׏�./�æ-�vJ���YX�_MsM����m�C�e��³Evn ���b����,��E	2��+*��ޗ�Zf�e��n%�30_�`��b���ȋ�V��ǩ�Z��u��]<�i�u�̕`�XlxVHYEB     400      f0��F̰Td�Y<�Rz��Ӑ"{4<@�#�X��)"d�tCx?(�����b�9k�P����P����@H�(�}[!+x�v�q%�>N��γp�E�k[���+�I��]Q	�G�����O=r!�\�r �h�����3�=��MŊm���!l�N��%��ZM8���qC^Z��;�~���I0�������6�\�[�&k�ʯ�P�A����tg�8i��1�������XlxVHYEB     400     1508�~-��e����|]�Ǖ�O?U�A���0k�;�{s B�:����Z}P��q5/�},��4�;�g�OO���|B�C���x�ǜba[�]ژ9��=���&�̺��	�Bݳ�,�Th����A�j�g��@a$��)굈A� ,Y#5�Dlv6�|v}'�1{}�A5��Dq*6րq�-��b�ƃ����k��34	���*h�L��`C-=�����	�����.O�r��lz~�<�Ӷ�۞�K�D���7�@���yP61G)�q�c�����T�R�﫚*���K;2�q̩�����]#)��n�$@7y�xo��I������Q�̾XlxVHYEB     400     160��Q��;6|_JH���7@������r=��FOY�<`����Hc�E��Uo�Nss99��k����{"}�]w5T.jFg��������%��k_�# `3��_�������%�^E�.GL<X�ĸ��y7qܙ��ឝ9Ǐ���q�z�o�� �ZP�@x}����������y�.��kH!?�;�6<�W�N@�e��y�e�W3�K���B(���s8�d)��$k��n9��*|�׊6c'<������:��Ȏ��`��ZO���t u��N�k�_�b�o����L�b��3�Ё���0S��%IG$I���p�����"P�!����h�(��ukc��v��ھ$W��?��Y�XlxVHYEB     400     140�ctB8=�h�� �k�zOџ�HhOҘ�3f� �@N���ږ�����J�G ��Ψ�RE�ő`}3�U����"5@��v���<����Ť�R����|{������} Gl�z�_���������4��er(��4`pʱ^aw
:�l�>+&0ǚd��y9����ޖg<p�����m�C�M��!���+0����1)�]P��V���33�R���ehYi�o4*������w��2-��ss�#�3�k���<���O��=
3��:^�a��,��~���K��6ɠ8�j��w��7*��0җ�^�XlxVHYEB     400     150u�v�eI��Ҁ7D��5]Ȼ�)���ߓ���{���,����{��vt�&�M	6�`.s���-͢I0�YY7�-&����Y���F˨,d$�ה�&k3���\�ts������E(��Dn�������@�ӓ/���͚&��[�ьH.iPh]a�:R�؏���蝄z�Z	1qD����6G�!Z��S����J���߹�-�
,�i0D���V�ZL� ȓ�� �N��-�9�h(��4�+U���^�����'�����go��Y����ZG���P��0ݟ�����*N*�[
5��G��֏��{��>���℅�b�[�XlxVHYEB     400     190���?L �a|:de�}a�@@rr,Ӕ��:6mA^r�� ��������┓ۦ`���0J�0�#'X~'o��t��F�G�%?@�tc�z���ְ�q�F��&�M���#�~�
�n=;H%��L����$���c�_])�}��J=�����~�-85荪a2W��c��I� �0�_��n�&M9=�%�K�s����Q����E�دF��\�g��4��#����fy����aK��!a��A����x*�� �j3$kD��y%�+�Q�5-ۼ����v���(�6��/�i�oK�A��}���<&p��ZrhJ(|��f}y\FM���@�셄b�B�o7�5y/�N��+z��(\��#Km��A�cޟ�l�.�o2υ�?7���*XlxVHYEB     400     120C�;y�"�����q^�+���1Gr+�
[��-��������G�[x뇷�Z@���؍Ӹ���j/}��q�,��O�U対?�no�"�1`Y�c��Z�{��0F�ۗ�5}���^��,G�$Q�Z�_�H���Cd��D^��w�p�H�T��aH؅!c!b(����;��@�t�,5 �y�;Ԃ��nW�v�{�2��t>C�s�;%�h|clpu�F�X~1����~ ʽ-�I�~|�)9���L����I2�
V��p��Si�+ n�N6g�������j�MXlxVHYEB     400     150��r��޾�#$)p+�f�iS�?���h�<9�mFH�tYD4���25�;hD"���E��0�2���O�Us�Q�����'���}�BNk�(;��S���ETȒ5$�~K��G��������+OgQ{���YF ��K^Fu0���p����J�_:T�_�\ DjGؔwх�?�v߶�A"��V�{�i�|"ڨ8|0��詓~Y`�r��V 5�$~���C�Fw+}���I;�)�O��p_�0�".2{�T����0���-Xu`�t@�)�cȔ�*��`�mu�W@���)j�ݖ��;y�HˬN���ا�%_Z��3?}�P��XlxVHYEB     400     160�_4"� 3|6L̩�DU2#UP��hV�kj|# �}�N�$��k�� ��o�ͱ��g3��A�����!��c���1�����ӊ@����E�ďT"��1�,JO����3<�x�?�)�eTo���7a���:u�#9�&�/K�z��t"Նh�|�F2ȭ�OQ�FJ�k��D���Ti0�ŎVr��n�w�s��?��C���H$q��j���Z�����T>�O�葱}��P	��}z��H�A�*��΁:�{ ��gKx�v�.��7Q��0�4�=�m�a�4еLb���AX�(fί%�A=8+�P��B�%���%a�2�P��}y��Y�݆)�+XlxVHYEB     400     140���C2��u��2������2ʡ[DnLLe�N9�IɁ"��lNX1ؠ�c���絰;v�=hM���u�+>��ˌ�����
��;��|�j(͗#c�|%eS�y\3�=Ĩ5@0�~ ���((��t�a!���v����V!� a�)O���I�C�C]�1��#�Ī����2��0��8j��1��B�j�D�g�<(�5i�{�ݛQ�(9@�����7�������R��n7Ô���9��/[�'5�JB��)�<����MZ�KO�_Z��2|�eyPr�5�MƔC�I�gw�)|ș���*O�;��d��XlxVHYEB     400     180�,���8���*/�]�M��؇��6�&���Ѣ��C�������/�;�)��a���Ӝ�z�kk!L���@��O�6����_�L"�a���P��?�s!km4��Uf��i���(�=�������b���[�_����d]igVav��8�o8���lƹ�E.z;0�I�n�C[*W@��:A�W�E'��.t���(�.C�μP?��j�V����� jkϿm�ֿɥ����ߢ����J��D����W�ol��6�&A�M������h�.0H�ȇF�7v�!>�'�:��z/,�9h��ʗ�{&ו(~;�J��l�ۚo:����^�ؔ�e������a���	�����2e��z�{XlxVHYEB     400     130}s��ӀY~ �`�vGcfC�@�X�H�y��X���
Ϛ@���?�E�V6�q�x���Y|��:2�hҁU|���.2r����ώ(9��~��<���s���ats����0f��{&ɽ����B+�Z�5L�6&�Z����.]U!	� �w$䑁�o=���P�_hcd�D\���F�s�ab���Ƿ��/κ乊R�8Ƭ�Ǘ���ʂ�������'�^�X�X)��;�k�=fu�I5pՏ���&�����%6���X�y�qxb-�I%'a�i&<�օ�3���m�.�!�XlxVHYEB     400     100�)z�:�}�^���GK�	@X
�ÔV��UB_s�%Ù��b����2#�U�bޛĺc(���'?|�K0�嘢ٲd��8���x"ǯ0�ﻢF�cZ�~�hO�M3Ͱ��z�>�7���	˾^)����W�8Sps)�l�	B$Ti��Q��,D}{�Z��n���K�r��U����9�d�8��N���]����CB��P$����1x���v��N\�ÑK�ܿ��Q�'�g*;<R#���2(��"ZXlxVHYEB     400     120�&� �ï�! �z��ڠ�	�M0��ܡ&r.���s;�oc��
0	k*�'S������5C)
�j�r4e�nY��df��<h��'�ڒ����<��{YёzY��sw���wF��P��[w���q���A^j2'�Ò)Ó����"�������<�X諙��\��{�t��H���o�Ţw���\��ޱ�4hn��6��S���eDBڨN�OpbM�M�����W1�lN��ȷ?�ة92�~+AI<n�W!;��η
��XlxVHYEB     400     170W��mw����7�b�u\Sq��[���8X��hݣ�����;�h9���� �� 奟+p'�����c���5k2�[a�5�����6E��%�uwT*O��2Ez�Ae������ƘH@8�.���������ˤ;��"�Mv��(˛�0���R۵���F��ֽǈ��m0��g!ۆ��IΆdf>3���	�f���T��r�T.��*G���8/G�U "�i߇�Z������6��,�x�eMQ?���Gs/M�����	!v����s�-�A+bg�]a�-N�����.�IZ8�+ ��(OT�K0ǢP��>�eq��L�J�l�P3`�ĝ�;G�sث���e�
D��!Y�9SyOZ����XlxVHYEB     400     170C|Q$tn���Z�[��#C����>3�o�qmH�����j
��?�LF�L�_3���u�9~�;�x�~n;��'��a��WP��
i��pH3l���|G^�4�9����d[�<��X\3��Q�[�f��u��p����ۙjC�*��Me�5�!���_oi�5��GC$w�u�1^b_�>%/�m�9���4Ib�N�YS��Ps�_�$�x�vڲ�F��-�L��s�E+F�ޣ��^�Y�3q�1������Ek�I8��"�'�E؞0_0g~8GPȢ���-k�����ŗ�H0�w�Բ��P3y���j��$F�M��k�5����pj۬�.�3LE�RS�MJ�i��� �����{�XlxVHYEB     400     190~0�O[;d?�-��m�j#��Ó��
�N��`��w�y���ޓ61Q\����	��XD80�B� L�i�B�B�������X��P�N��J��(����x�y���Y��P��,t���
�bs�.���;V�zK�v$ �:�nn���";�؂��Kz���kR�.���!g��a��?�(U�l��*G�c;&ؽ�+��亦N��_S����1U�-j �!��M�5��y�-�{03ls^��Yi���:2&��7����}c&FO��|w�-����p�ӟ��1�ô��!�TK[�3�a��	-�)	n�$Ԍ�i�&p� �@>�3ǯO���9ْ�
��D�_�?t��	g�US���>�E�Ω��wS�d��{2��O�ۆ���XlxVHYEB     400     170zL��*�6T��'���������#Rr����z�Յ�1cǵ7�=]7/2X�� �	��V��q#�*Z6D�R�Q?䷴i{�v5�	7߉�aX���(o�0������w9i+L�7�Sw����[��!
Y�>� *ZKg�E��\|�[�p(w��|�n1�vq}��s�m晴@Y��g���|�0I�	}{�����h��7B�81@k�����1Lˍ�/�6?��W/��7*T�;xXã��)�����Y��];�`V��e����\��>t�"�K�8&�����u���m����i&����_°�%�x�n*	EG��a~|$��"'�|�u��(���$=l��>����}�5rXlxVHYEB     400     150ߦ�c��Fv�N�>}�n�N�i��ٜN]u;��FPn�*
��In�oI��.����SC�i�m��5��s�!ۛ�����O��eɵ`��W����Ճ�$�HtB�G�!2U�g����xU�`f�Bi9-�Q?	I��8����+���D�ըݩ�t �_��N��p6������cg��~�Y~m?���lA[�^�+u��2W��wulâ	K0�٪�S�/��w6�~������_��t�_�Kr�:c����Sw�O���!�����KiH�&HF������7���,v80�0Ց��D���5&:�a�3��tm��}ѼXĬr��N�~�XlxVHYEB     400     170��7O_DdEX�a�������&=�#� T�)�h����۔�X]�\�)�^�e�m� ��#)ȏG�oj֦ʪ�D��[l]f>e��$��;m�`l�T��n��1a���5�~_��C�_Oڠ�I��M���3	���PH�a\ՙ~%������(���[�g�����p����K��=��|�Y"EeҔＲ�s�)�7yh4'S�rT%�@U%F_1���&�.�E
;{�W�l��>o�2
"%re�����ճԸtQގ_~����5�Dy�U��8�fD��3���[ef!���0�n�������ж�t�1���8����g���`]1T����uS���K�U��7���d�0LXlxVHYEB     400     130�<����6t��sN'��c���4�n���y4��W(�B,��o<�d+���O7m�sw�������\G�Vݍ;c��5l0��i
E(Bo�������Qj�
eh�N�ݥ\���p�:�p�����_y9��h��o
YCWX��+�qy�\��\�`�<�]����7�tK1�讉oE9|'q.��
���!����1��#]���K��Yy.<�l�2�;10�͏1��la�`�}�G ^�5�^v��G#S!P�N����T8�Ƅ���Y]%w�O�����y�"�9#�~o���Ƌi�XlxVHYEB     400     180��R��!NI{CeO;h��s��1`yni��)��F�h��?4� ���9��^b������!�K)$��k0�B��XX�ν#���zdS��lUT���/�ՠ��&�ٮ�^�I�Eb��D��u��7�c�w���;��-#R��G�ٯ�y~~ĵQ��PCc[��!��Χ�}Sby/����V=2���	_�;J{�iN�M�\d{�F"^�PO5K[n��r҆"���|Ԉ�C4o���P½�է!�Ċ"�;h�����U1��'���7���b�?IU�3/�����0�&J��P���wa��t��O��$��f�1��}PnHp0h��������[c��L��LG���N+���ć?�݈F$���b�V�y�YĈp�f�.SXlxVHYEB     400     120��J�Y�lDָ�<������T��?	�Y�L���.�S���S�jl����Um��7�7r�+��M���x́��{+4�Zu��<��<�h>ٙk�~1W�{|��]�Y����9W"0�|��1�A��_�I�.�x[?��B�V�I!�@<z�������}X���!F�*i��D;sLٚW�u��9�xOPj$���$��a�`:I�0gl�mؐr��d_*<�+!��e���2�[L����s��$�6lp�=�ٿr�xQ��#�`�5m���q?c�y�X)�XlxVHYEB     400     140"���Dk4%�7L����[O����}�._3��I���V8PXϨ�<��o������&���8�H���'����}'
ӕ:oR��_��uV�E7�Yڗ��b�X!.9a���6ˎV�|B��q�̜�$G�\���M:B7+�d�����C��z�`q���G�Dw}B�JEu��=�#WFc2�8�	����f����/��5?q��R�3�m�� O@b�ٿo7�;=c�o �	n<J�����}bz1��x�=���EOJ~��+0F���"�=o��� �ؠ56ݼ��u����P!XlxVHYEB     400     140��w9�dk�~dm��2� p@}R�{5x�U���Ɯg�(�C3����8�?�_}��R5ԭ?_�!�8C�$Հ�,%ŗ���wM�t,Xk8�g��}���eM�z�'���hJ����9�IM��}E��&X�J<&�9�sڝ����=��W)G�n��oE�'�[#��!sut�֌���xq[��*A����?m���`���ϼ�Яb�v��Qr/��Rx�J����~��_z��2���Uc���|�������П�1#w��SF�;g�"~ňD�CbD2��`D���	!�NpO#��Ʌ�k��ox��vi��4XlxVHYEB     400     180�K8�u+� N���;~��K(:��)����ǩj�h����+��C`E;Y���4���ubi���ZI��LV|��~��֓p�_a�ɩ>3Fq�BLS'�"�"eﯓz�4kL�V
�6ƦQ+�KB8+�hK�ӽ�p��u�a����"��eZ2f"�P�O 8��	aH�k��<[ݯ��ޣ��j�*jGp�D�@ex���1�I]<�I�������&ga߷<�䏖�$�$X��wS�o�屿����C��DBBR��#:��}�.q�=e�[���Uő��Xvx�C��ޑꞋg�L.6��ޏU���?����O �^./;$έ��x�$�Ⱥ��;��b��;�dOi�x
x�%bvtH)�]�XlxVHYEB     400     150e�L&PTR�9F#�z���?锯�iU�5�"�K2�Y�>ˇO�7�0ID�N�P�:S�"�~�q�N�!"�_��6�'�m���`���uzR�R��ێ��[����_���]ٽ�T�H �0e3A��|�R���L �|�܇Q"!��~fC0�4,2sJ��ع�L(�Ot9�`�P�j��Q��~D��mi#�����
)�ui�_P�ъ��8�9�-ݕ�"- �\�7�6�\�Q�z<��I:�"������Z�)�Ey�]���p�%gmo����۶������?K�$I;;V��X�H���l�A̺���"̞bj`P�����6��XlxVHYEB     400     120f��Q��KH���C	��
#]�0�<���'G,�-l��2�r}��2���w�Ҁ]Q�t��.���S�]��^�9��H䱽l��kB	�ɚ	�g?�t��['�Ƅ/ͬT�s�����>9�P�e�x�mRc_&s�� ���˴�	�Mh��p����ݒ'�N}ת$�>�Kq�1�#B@�I�HV�t�^V1�?�N(k˟S��T;�x�y�>����9`Wψ�6mT�7`��)3Eh�plsѣo`�/Ǒ�oN����j�K�(q�0���Ŏ��/�}�XlxVHYEB     400     180)Z���)��&j��t$%���o@t���>9�d����;���ΐS����B[�M��$
��ee�>\7�Q���?b�f�s����r��mX���k��a��M�X���ڄ��&S-��H)�x����@<����*sN��Q�e0dN�~I�;�1��i���<f�����L���t�<�[#���@SQ���6l�AJ��DHY�����c�>`7�����>����>5	�M�5�?��<��ߞ�Չ���ƚ��-�Px)���FֵDS?� &�� �4;��5a�1��s�f�ֳ/�.�3��xLŁڥ9�n��K�/�������}~U2�)�{��L	g�y)J��9�qP�$�XlxVHYEB     400     150��6���=�D�G=T=y�u=e@����n��:w�n��ѩ5��&�w̂6�5M����d-��M&+�h��)O.�͡�!s����輭�8��>�	$|��Ok����kVl�#T���g@�U��2�XXO� �Ӛ-�ۂ�-��hm�����*���)9�[��,_z9��,�L�3�	&��m����l�6�?z��2d.Z��>H���8|� E��^a��h����\|����ςC�o#��qr�J���^���8䒋���qH˶7d�OQ���~�+?�%K�/3�]�ڕ�ׇW��{ot���G[���2� gӳ[�XlxVHYEB     2c3     120��%�ߟ�F�mg����}�V��C�%�U�4r�G���X���g>����R��.��Ρ:%4VI��5�.���(�,�"#��r8���XbjQ�}1�ӪQ�G=���F��o��. =��7��I7�gV� ���m�~����߇}�Yb�U���6�P���b��\[���m�{�/?<+����L�}I�ygč?�u�<���P;��sY9�s���Uo���C���A����u�,�W7g��X�Jih��͞+4}�"W)w˃�l���X�p��òPp��C4