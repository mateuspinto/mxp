XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��
(w���)+��Gs�7f�*58@(X�q��>��Њb?��`scl��A2>H��^D���اYh2�8����Ǐ�	_,����i��槏[�ú�~z��_"}�VL/�>������_" ���[Җ��,r������"D�ͣ0�v���i�zM�i/J��E�ԉC�"��R/�c3��*\�t2�v��1ɴ杇���V����p��k�%�~���?c�� �?M鳾C��c�ݙ�/�������� 	��<3:�s뼛�P��2~`�# ��tܙܜ��{�=M�C��S����u���\(������:��k9{t4Y�}�r��P\�c�����}�#o�rcT�m�i��t!����v�ހ��H�]����;�0=��Ez�{}W��J���{T�H$Q��ϥ����PO�R��L�Y^�7�-"��`����af��wN���|ak�k�m[m�@b��r����SH�#�$���
���|���x8b��iD�dV ���}�ŭ�^��/N�frR�)*�tf�N������]���l���ͱ��ooPk�p�Q�l&�?����9��NsS�ZH��0��{ �(V��<�`	Q^�r>7����=����+�U�C�=iļ`�j�j6�\��#��s�F��9ś�;S�G�t��SH���j�9�{��,��?Ɋ3"�p��k�y9ݨM�;bi�2W�?�)&�S郀ċ�d^�I���O9����H�S��"��	|.M�XlxVHYEB     389     180�y�Ҡ���>�c�bhF]��S��y�7!����O�h�-*�H:(-��]��؜�R�[�������� y��
�nHi�Y�AT��-�-���p;�i�4�q�?�Mk3�Q�da��)�˵�'�vT|��T�ݹ9y�+Ӧ�(@_�
K�g�] O~��XM{EG��5�V#��p��b%Ѩ]j�4��&"�伯���9�r�P����py	 ċ��� �E�"1����.〮{쩝�����<Y��x��#�U/)�g�9lRV��tW^�����(Q>Y��H_2�<�D��~����O,
�wBV��f�=$���B>��\�<q�	�-S�-�������қ���+ٞM��#���o�Q�O5-�