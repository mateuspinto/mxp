��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���̞:C���k�K�-M�7&�fϵ����O-x_�0�*��hr��Pe����\W3���Nļ�վ���2�G�f^�5ז��:���g%�|�2�hj��8x��oe�aX���z�&���߮�����#�Y˞�(gx.&ֻ�U�$��; �����Y����M��[�v�1,��{�ypƛ��� ҅8�Y�/�W|��׉i��'��l�wO�d�A�/�(��T�6��jO���� 7N��d9���J�Z8mCs�������ҡ?�Z�D�k����sBD�rR��F�_���1���{���b���6���	�	���7nZ���[Ƣ�p���3�>�ǣS����>uP�Z|w��g��}�p �1�G #��7_k/�o�����Z�{���]@͏�Og�6��Z�5b��~�kN�(<�j.���{
c�~�&1���w�
��=hFxr�r*.7�"�(����Q͸I{U#t�V�@�gš?e�hV�'�	��@�_/%� |�O�{ ��y �gIn������Pį�67Cx��-�2\�_�Z6�������ȅ4�3۴C3f<!	PAq��4������,N[U.&�>�}W���kc5{�7!�H�*�V�Z'������������4`��4G��_�Fkc�ddNg���\<���yʮO0J�W��/R#�J(���W#���9��Ԣ�Y�d��k����y$�Fgr����*����g�D ��'���;j_���ՄF{5#,"�Mn�݆�5���/��A�y�j2=}Ls�J�.��E�F����nk=�>��7u��R6R��`�ү�Uq�b�I��[!��j/%�7P����˪7{%�|t�}�.����3/hE��@$�RA�?��h+�6�̣C��W�D�@[n&ҝ���� ZP%T��6��r�d=��E/6W�*2�!ĭĂ$U��녳��>9�4G���Z�݃
���>+���!>��	g�_��@!{��S��l�⊆�f:6nsc�� ��^%KM�QµmU%04e4tb�ΗΤ�rI��b>!��ݧ��뵲��X���H9SH��Y������i]�P�8�B���HTA�xd���t$Ys�`-;�v�/�N�I�޶ �^�U���?�J���gA>C-�����t��2���`�����"��;���F��#^+9��+%�1n��$�۞��/�Ա�}�V$Sn��V~����� �UQv�b�v�kR
�R}(���k-~���U��2mP�B�F����!JFڣ��_���ھn�k�&Krh�,<�zg�c�ՙ��X��)T�fd�A蔮���$*��,&�c*�f6n��f�*܍�<�F!O��8���*�.2C�F�)�3uʆ'�x\��|)�x���=��r���@>����C�WE���;O���m���[2%í�?E���B�X�����Kd��z��.�e���s��̮��^����0�J�"�7� �
Ԙ��Ѻ�뻓�W�S�ڟ�6�,�l�w�&�l�1P|�_������]��aX����j&���v�L��Ew^����Y��d��}֥�_�e�.�ZN�(�+��/|��_��_�=2#Oh?��c��Ӭ�qj����9*��&��Bl=�s!�eA�A����ͨ+�������vh���?V�X�ǌ�+���s�}��tF>���1I�@�׵*�s�-uܵ�Ѹ÷�##Y���2�0A��	�������a}����+���'^N�-��̂u&�^�k]B�����i���0�7��U� p���s�@�y^�y��w땇�#�3+= {���D�Y^��Q����,�+V�����6:��Xz��h�1(�L����9��`�Z��f�\٦�2��t��/%�\���ܵ�b9�%��ő�z6 �@��"N�Ѹ?(��� �`���swcw��AZO�_.�`7j��!�����jˠ+�:_�����I��z�� �����;u��EQ�H�Q�v���a$�����P`�v*�;]���*�{��EI�6�y�l%��M�������U�ѽ\�;3�*�0��]%��E���4��~SY�"I���iP�?����r���F�� ��D���~@�e��L��ۮ�(����V�������SYy\�'%4��p#��A	�I�E��k��f}i��F�3&�x�d�(�z���(�ʴ|?Q�%��S�^̮7O(g҅'���RF��K�����~���_�@%mH�|�1O�K$�I�2�t֙��J}�������z�vL#Q�܊̚�ގ�:P]��p���馻ŀe㷻;gӺ�U�7oC�����%h;�k�a:�2��Z�L�R?�~��zP*-���I�Iڏ���<�����/���@�����w���(4u�j������Cw�������>Z\�BL�Q羅F*;Yj��&a߬iC��j+`�W�	�\��Q�n�򻚜�5��0I\�눳�Zf���e������F�z$�盛:	�ƍdB:��A�.1�<)�}'�'k�+�����k�Ō�����w��Ǆy���Y˔��(j�X�Cז.�_��P1'kQ~#O��g i޵0��2Ս�Pś��\�~O��v�IڻC��߇}���w�v��׸8"��Kg�3�ճD�P4��������O�P��(F��o���t�L������<%�[(�9���a�=�4�yJ��Z'�.�ٞ&��
�����W<�[�K�]�=�5�Ze��d�?��Z�d~�"����aA��s'd{����g���[02����&�T���F�{�����+�P[��cyAZKÃ5ݏ)w8!0&Q6�N��sT���%\G��!0�ͣJ�|�0��P�����@��ɍ"Ԫ��|!G�$�֥�o���
k��lGbp�sa��9�]g����'��)��>�\z�L��_�i���[���ٝ�Aü6����.����˔-͝0��aV� �����[� UY�-H����Xś[��Kb|, �m!�>�\�]�z�6�����a�j��#�S�Z�a�7�[���;�.��%q鶝�M�d�l�ʗO�6�ح�-�կ?e(�m�dV�D��`[)3��^¬��P�k��-�Ԯj����,�FW��}�Sp�]��I��K!�������-4SP|~�}�����ďw�=EkϹK,w��k��<����-��^�>�>z?�	gM�A{�t��}Ճ#m=���Gܥ�M#X��%\�:�z�3�k���~�8��!X��_��%����6^T������o�k���0+XB�i��+bmB��9��eQ��\3�t����O�F?� tVBk��M����?"��pcwq	둩�r3ޮ���l��ړ�X������|�������6�٢�fR_�O~�VIr��n	���~9����o�Gd��+.���|sy*ɢ�(�0L�L���i1�M�"h_Aऒ���V	�[[U���t���g&����;�Z2=�ѵ��'���򯭟�-��i���]"���&���o<�-y��6���<ϔL�D��1:Я{Z&Zx��э��2�e?pi8Ag���zb�aȱ�V�R#���pȨ7�E�WUu�� yX��q"�r�4�6�v������Ͷ7 ���9l!u�j� �˲����a~� ����a��:��� �R�(�G���q���h&a���=�|E�.��B$yM�V-ŷWq�Vt�>J���~$���+��M��zE|YR�5F���$'�6e��N_��->R��|YuE�%�&׶n�mD�1��Z:�g{�a&��#�B4~o�B����%�6�=��޴���ؼ�E`O�m�y��� K�Cյ��c�˲�֭s҃3ߛTP�A/1�������M�Af:��(S�K�л@����PJv'�t;�J�T
+����r������ZBĖɑ�<O$|�j����P�lc��˲k{��#�u�Gk!x˘�����9�mg͉$��]��f7r�e�T	j�w�P#��.X�>$Н.����o����&��;]Y<� �[Yk����KUm�j��P�.�a�W���F/�e�y�o	�(�66�7�h١�W��} ��Ǘ��w>�9(����PM Q:)����J�ˑ�����	䀽�vU�A��@���#��+Dn������	���O._;v:U�AA�� �	{,�?��@au��U������H�1�X(�d-�/8@
����L/:�R\�y>�����L�Q�kwP�M̡�)�b�R�0M�����S�6���֨qJ$������@�<�S��J�Ȅ{xx���K����'�JpC���=�nt���"V^�!z��q��8pX���.e�-gh2D6��!��22����\RNh{v��5�3�_��%��ǅt��c��L�v)N�(�8L�����Ȭc�Ɛ�r�y%�1���
� (��pB�k�;��i����^�bngo1x�O����v焊�?��K�v�	���h6�V/@G�ON@�!8�Z��r
�[Mj��1?�S֍"�
QlI�����6��Q(a A��8K&���Be���}$�\&�%�i/�M\���4�`��I�1���
�n'�M>�4i�r�o��V�b|���>J�d!$��u�#���d�g�1�\�D�c��!:�����?=��,Y�DXĎ�S�1
ͬ�ʷ����a�}ﱟ?#5�ȣ�"E�x-�?B�3���R��>8�!0�<����{݂�%Ax<��X��&T��]��z���Qq��pQC���⑒n�t7_����)�I��0S|3�����j�MT�yM��`D���@�u��Y�^Q�����.b���J�8����{���������ke�r�=\Cm�(�\W@�3�y��:���6�D��:�8B��*_��8w��=�"��0�а�ii(���#5�0Tu�XQwYY���YS���҂������q:n�-��i���0�i_�k�:�de��6/q��vö�+(���+���l�U��m���	^��I��e8��_~ �ѽ��/��u�
�,k���&n�=H��I��&��b�)\H�l���2�SS��߽��>����J�k�=��
>q߉��-�k*ފ�U��q�Z{��i����^�n�\0F�刊��C+A`�w3�'��P=R�^�Ə�_����c��๻��U�;��4a�Jh��Q�d}�`ax&�
���I��Ҿ0�cz�k�;���\|����VUD�L�1�񚥟�.&�KĀ;�}�Y��ÉÚ��ߵ�³�1��`+5ߚ�5h���4�=����;x�ZM�r�M۰��j�^±}
zX"r=z����l-P����oN�D8���#UW���y��=ĩ�6���k=	uՃ�w��np��c0&^s�E�C+��l���C]��e�esz�BS�N�o�[���r<x]Z���_R���B����7�;��n�%���{���Z ]��#v	6iP�f;\h@o@С�]��v��T�YDf���q�����l�#%Ӛ%�2����@��m��9
�p�O0�������p���2�1p�`Z'�R�;��qn��D|c�G���]�������lڀ���g�7/R3�}���Hc����5��S̓aђ�g��g=�D���J[w'���x��%�}"�ܺ�[��(5Q��$V������W��ߖo�#���1�_�)<Bz��%j�v-�����������fM�v0���:1^��&w=0�����jim���b�d;5�6N!y���+�@� ��mC�x�[��?�G[2a��;����ox�B��YBA����=���/���C�v7��{�bX�l�LaK�B�l�X$�!G���#u�U�
��"���䔰	���O!�<o��t�0����
�U���o�F�ɀ�e�}��^FNnM�55��1<�Lk�F>3�nr���f�q�e�&m|fD�������+�5HG_�Խ�;[�;������5 -�o�8@���п+�>��p*�4 ��>dp�ňm��n�Q`�.��0'e8L�C41�d��UW�1V��s��h�l9Q^Z�������@H��}|.�$��o����&#���9��X���J�uS�L����Uc�A*��F�+	\��-mv�k�}z�D{����6ۃ�ڦ��M1��E�$�H�dx�����QӐ�6���kP���j&c����AN�:	)Ψ�Վ�5�������4k�٦0�͒��	*�	!}�n�[_��4��<۷ׯ9��nX�*��y�Ύ�R�`��}ߺ�[�趓�G�T�H��J�����*]/?����'�U�fS#d92�e�x�!K�٘1Td�?i%(��U���d筅"�?l`�A���{7��)h�%�zZ��zy��{3���ց��Z�7���$e��}�dªK�u��v�>�ʨ������-�%4��v��'dO=��݂�ў<n��\�beұ_[�jr���|��D��*���V�6�V?�G)¯�e�??f6(쎰>>���u�5囆����!�Z0��d���1>��%�5����&�������H'���������/�/��Ϫ��~ gGI�ޚU
���"I����;��=��d�G�=A3���[R�x�2;����;��v��x"�<߭�,�<rۗ���yM� /%:�z���r/�s��sk�0��ȸB��@�C�V��z����F�][5F�KO�pL��ΐ)A�h�F�����`M+�.;���]����Ĕ)�jU�9�d�>q�(D����(�HR{k^��ELE%`EM���.%4芭8kT��oE]���|F<w���?>��y��(A4T����vOD׉&�V����.N���^a��t���K �}_ð����C�����^
��F&ss�`�|iu��T���7���3��/vy¹=���'"���	A4��Px�A�ȕxfr|�݉�[��b�6Rt*���E�gg������rI�`�{�Q����Q2AZ��V���l�	ⵉ���hZ�8>T?��<nS�s2#8�� �1�K��0�1�s�sa��j,��B�u9���p՗�d �%v�p�xMV��Ncd���l����(2�xW�]�'�a7KW��ז�4Y _c��לd6��n0�I�q(q�Z�y����ѡP-!�*Fh�=Q���6 �.o;�.��	\br�6�=�p��/RfW�?��m�@�~�N�r��!.l��g��`���1��y� m����#�^��h�iMjU2T�ZW��BY@�J{7- �����05�L_��υ�}���ya7p���������E]f��|���V0����R�7�O+��3x�w���D���hs�[�='�7��t'3���c�4м-��_��^�F�J9,iw8�	����U��a6�|�'.I�}��.'�n��햐�L6l5����z�.�U��*7W���vR��Z�:'�é����H�Bٺ4R��k�5,��%}R����f��O͵M5_��d(i1�ԄE5S��n83?�.�>Æի�����f��_�>�76�?�@�/��=� ����h�ή�T�I̞B � Tr"��_���$B���ڇ�&��VȬxƖXF��*׏3��͘�/!��O~y��ˌ��1�l��>� 3��!����������]s������W�G���J2��Q�J a���#��c=�C�h��}��$����DLߠ�ȌK��h.�"����Q��H�a� �4N��(/���G�a�s�c#ȇjpuԦsa����q�j����(>�c�z�m�Kwu�R�x4�����G#�wǂ�<VB�<h?y� `oˊETE���P�^�W�ׂ�ԋ&F#���\+v�bs���Ł��??���=�|����?G(��
`:�^��ZL:�J�3yI�=D@g�RY�r	-�vtv?d��*m�i0(Ŋ2�g1YN�P����h��1�����]�W�8 �D�hB�9i�%�n�\�Jb�����q\�W�� ���f��h��?`�u�ِ��K|�u�;z+gr��ӈ|���7��Fv����*vÖY�L��܂[h
Z����:�	�D��͎4�<�'���� ��W��KfM����ur��0�_rYE1���N���L*�� ����Bjo�×ˊd�[䒕�`�拨���q�I/��z��+ݠc�䝁XPqw�%,��C��r�N'�r�?0'�ΒN�\��ʅ�-��E��]J@
q� >��~�����;�!� w ����6���e�";o��/�iy+5���D�I��+�q2�o��234���<��{���՚!\��.40��?>Pg"e�)a,�!����9��TmDi��f����Y�z�j7�?v(�{�O\�+C�:�~��ɍ�9˨���kp��X�u�D�U��n{,�@��ǫ�̳$Z�{�T�}��ɛ�c`c틠��֤������,��t#�#��X��Qc��!����!����b��[����#祔�_2I6cs�e��j`�\���G�_@��,2����\�&��	F��'��iW��*�~��� �Շ$bpذ����^�J���[��j��xi� �O|�k6��i\�s�	��n_��oմl��1��A�Jt3�eq.X�OSF��`4w�����P�w{A#����J]���8�MH��j�$j���W@��Î�W�fT�a,�o�N2٭s�[Ωp��T�1"�U�aɼ��]
=�g�D �b_l����j�B�O�����E�`KUr'뺏�����H��ؘ��6s(��O����+���*�ڰ����X���by���/��A�4���Z��� d��hj
E���a ��"pˎ���;����aFu�c�r�b{j��Ι��ܿ�qY��T�
��*��r�0[
����u����lO��l@0�rݒ��x�N>�L����
�eM�����,`ñ1j��N�7ܱ���v.��"N\!5��g ?��_	ם�d*Y��!�'�(���L�.Z����p����#��٭uvDp喴�C�';�z�ľe�k�
m���oͱX߉���!b��zb�0ʤ�"�pu�F�Y�ܧ���\���ƾ����o����LU5OxB`�DSNCg&O����*�����U��g�
A<��OX��.���%���R��	$����Iʲ�B�KUc�]�N�N�e�Ĳ��ѠA+s�.ɃS��D0�l	�8�#ѝ��i%�
�Ԁ8{��8�Fg�����?��F�m,3��a����	4xLhK���]1_A�v�ɻ>U�&��JVka����Y��oR�~�%���wk�`���u{��'^dNҒ�B.	�����f�׬ݢ�����Y���W�<H?������W���w�|)�U���/�{�f���v� ch����G;��nR@А�B�p�{��m�A������9�~�p*�:I��,P�4��jtv��H�D�R�0��i��5���<���䘮B%��!8%�����g�"�Һ��Ԛ_k�������~�Hw�4`�L�j�ҿ�&���2�t:WL��'���Tta1Ue��A(P����C�;l�̌,7�@}��v
0黮�B[�rΘ���w�}�=w=}�A��u��뚑�M>a��'��!^7�W��m\�cj�va��APڶ���^d^�O�Gs�/!u�q쮧��_:�|�Ǌ��y���H��-LA��5���Q:�4vNA���3�0��H�p!�B?�eUk8�����ه��h�fǢ�bjK��4G��H���D���`xy�`������)�{v�#Fb1��Ԙ�lkyOD��<k�*�]������v�<M�q�@��$�<��/��0o�a�Eqe���X��G����E�|��� F&��]I��e�@b4
=N�ۉ�ÍAO�GK��$�g��^�ZV���
�iTqk՞��f*�3�$�����{ܳ��BC�0�/"G>Ew����mJ�RB��+�k�k�.�u�m;!xW˳�F�o�]���1���O%ͩ�Q}mM��^�G
�c y7�c�fv�`i|��6�3T��1�	W����2M/A
M󆝰t�L{�ץ�5��_ �T�?�Ϯ0�� }ڕ�O�)�c��b%HΘ���&u�a9��v	(0E������F-H��N>ylW:EE�rb��MP�5��X$w#��$t掹�&	�̯pp�!����F��Mc�]��F(�%����l�x���R�N����U��zJ3 �ک(<����/�	�,4wd2��/��L�x ��=={�RV�r�q���^%'"4v�+���	H�2�֋2���] �W���-~?�';���R�����W�u��ѹM�����%�a�ؚ���*ǵ�(lb��a.H�v�(��s�h�c��-Z���C�� ø��]��x�ٮ�+��P�Q�+@ȘӗQ�ħ����@�A��+��+N�|b�>� ܂b��T콬�w����0�6#l�ȸ�N*���[����\��T\�$E�̞i_,T_m|�KKa��� �Wv޾�(7���pGbz�[N�ÿ�?)+U^��|�sq��oO��3+�����"g�G��m�bNpCW�i���������$�+$�Q�q�>�����U�+.�#�[�� ��B�BkO��!ގZ����T�}�GƧ<���pZ�����ș3�%�٦;�3i����q������C�a_;�l#����j�~S̹�
�pG_Q���S�(H�؍��f��I�>_Nb���% o�$�eV.����\6\|�xXRJĮw�42��,��w���d�s�>O�]YV]�:h�ے�N�7�E�>�X�;�)�Ņ�a;%h�LN-Kb~Jj�w,!DȒ�Y�s�6��R�B��۠G}��Ҧ�ͻ��X��0��Ȧ�c����u�L�z�)'kK.U�2��ԯ�}?�?�͐8��ەh����M�|�����9���8�
�V�l/�h­�	�:��E!���UT������l�@��L�,҂�53?�ٴ��rCTY��@g����h+��̕�/�!�5wnS��y�Yd��J���t����fHk&�`C��4��M8Wˡ�ly��N�q&�ف�q����cG�1��cXR�ӧ������s�ʿ|��e�
���t!�c��\6�w96$l�_�$��F��<е���O�s� [��'2�J�ߞ�y���9W�F����Y�e���Ec��[�_Y4�Z�@ov��s�����~�e�!�1KF&��3'��X�H��m����������4:Z���\E����g�$j���Q�p�.X	��_�d����%��n�e�q��ij$��v��L��5Ⴠ�
ee�Z�e�7Ml:�}w9v��L`ܙ\I����2u�g��|����->�BW"y��v���6��m�k�ԕ�=�
���jz9�O҅��N[�mvQަu7��(�l%��"fK����l��(��_DdbumH0)���v�썧l>x�a��_gQ��OH��#��O�n)���Y�i7��� l���=N�X~Ѥ�U�mקJ�k�ӆs,
1��cu��WK�RUS�����-�����%�{I�tB�u@�	L�p��i6���؂�����?h�� ->Ԟ5���:��/�c��Jy�X��I�*?s�E�W
p�ݳ��b	`����ƚ�|��P���ӓ�g�nt,D�K�ϫ�Kij���J0��5oJ��pRk44��q#�/�F��+aU
�$�	�0jr�E��\����O�2'eEb�߂��3�=3V"���;�/��k�-�����@�����7YX�b�X�LK](�zfyv�9narH�F*K���f�o�K1����)T��p� �-
U��-��	�4m��c։�"VBH�5��z����p˝׍�{m�$r��Ȟ`6=�5o�5y��KopN��O,��]�=x�`7a�+
Q�r~@�bv�x��@
�új�3����q���D��-JP�zq��,Wղ%���6M�v�x`0̊d�����U���=���igO�yF* �V��7$x��������'Q��$tG�qB������D�r��y����a"��V�k���O~�2�t�tam3ކ�xa��������ͨ�ފ9�&�I���a�}�۫t|��'�"A��2�,S�E�S���!G7�C���1 �ߐb��ϔ��?k˔c��fg�c5gd������G���Y@3�U��f^#躑�o{�cnx�c�na�!���j( �������W�k��0� ��W�$�:�׿�W�8���BRKf�d"ܹ"���
:}0G*^�`A����Z���L&:���J�`{���`(d�JEÆ���Ǽ_�_qp�U�@X~�0*:�y�ΩE�L��M؝y��[��J.O[$W4�8���w��8��� Y[M4
�J�3w."2����+� n`���7����٬(�������e���V�95��|DJ����4�Q���؊�Qa��VJ�2fDծ����/�HU���L�KXO���в�(0ۉ�S�2���
����^��F�]u���o�Z�f��Q cx�شS����z"�8(���#�mK5��$���U1k��O�
kw�'nX�W�8OW�Nz{�xK���ot���a4�F��BLl(^��H�#�òg{���*��ѓH�B���Z����~��S��*1�Y��e�R[N�e���d�Ҟ*�s� ��jù,�m�c%�&���A����®M.�E���#�-�'V�د�����ͩ�d΂@{;O���CmA&9��S�����V�3����5gR�C�7��PN(W٥�[��yO4�KX�f;�#'�7���y�f�n`[[�`I4�Z��+I�ZM��R��<��^"����׭�T��n[f���m�y�=B䋋l�]VȞ>>�OE�ն/Ƕ�ĉ�ʄ;��6�?@讝�L�f��7��룰��6i�y�^��g���$�Un2��D�&�gD�,vR����iL~�C�?�i�-�^�@��;���0=I���s�]��u�j�	�(I�Q�C+��1�ؒ�R������"U���E%��[��/*�f|�d��Z�!���iw4�^,DW0����W)����m�T���l�#���a�&%�$��}2'���ϝ��xk�����T�����d��V������#�� E ��@�~i����n砹9 �l�ۨj����h�����3$�9�4)��������O��BE:���N�U.�)|]GѪV1�!	[�G!\�����jl~8��Ts��a�˹,k`�i�C�e�C��`ߩ��x��}�2b���G&���-P�;9u4k�#�`u/�(�����"�S��t>V;�w6�%�-�x�?��Hw'*���_�G�T�ۢ����zY��'w���w]k�2�O#4��}r��b'�l���9������t���$g��a�p�W?��@���;ł�SA�#L���I�?�fT���*��8��pb�����/���4qƮhʪJ����2�4�7>u�,ߐi,)���B�C!����f$����Q�C�;u#o+o�T<�%�Px�l��k�p�Ա�t�������d1̛xK�:��M�!ۮh�
aXm&i,��r�����$�᪵��\�촖�I�s�n�B����w�uo�g��)�*��M�/�W@�.��_�R�]���>�~������kC8�et%3^�\ؾ�]���1�YR�������?�F���fa��圉^˝��p���;E�e����E�/�N�:��H�ph���yG�M+��8od�e�Ϥv�P9��j���X<�>'�{f��g����A�a�!��}�מ�pp�w@����5�u�I�f4���y��$ъ���VṆqW�=������y�c����f]ƃB3}'�pfL�X��$:�p��񁴍Ӣ���6�QQ%4{h�ͷy�0��}����a�>�;l�,��b	�5��{f����tnU�g,��5�wWhQ�$�\��l)��2��(��F��ȷ�.~��i�V�g� �ߞ�SN���c��?/�38�.�Rv
��(Fj)�ݶ��Ş)�_ީc��J��������e���ƨ�8���
!����Q�,�X�з���&H߂V9*���{�����םY�7*d���fE�"8vC�X��n~��6���Lϊ��%!*�߯d��0��V���.����$Pay_Z���p�y�/W�48�B�6>L	���a</f�3�eVŵ��
X� x��y~.��Roܘ�͜���)V�D��� �Bz�S�NZ\�U�+�	q�+9E���p6>1�Ug�>yK�w�.�W�iKb�;�uͯXx���l���#�῾�P
�΂�/���p�q�>�P9s!�0�D�	A� (� �J8�T�ه;tBeS�rB)��~ w�0Wh,�h��Ar��?`��=����S�M�8�Z�QgHV�'�:�4�̠��L�
�_�xJ	Ŭ��U#����~6�Q��MM�S�r�N��������SG�1k�?�v���?�%�T�ɆJ���uX�2[=�eO�d��vET^�ň�=X�<���>���N�������N��IE������D1��_�m��!�TO�}3x;K�v5R(��Q�Rl�2����*�
��P��q`��K�%  ��6/3v�)�Pq���GD-=2_V)��["��8o��b�)Һ�Ό!1��3:'���eK*�6��{V�`����|� ��`���q�/�	�_V�Bd=�_�kap�M���`��_��f�$�7	�g�(w3İ͈(�b�1V�ݑ5w���NYF���ov�4�� ��8�ߧ�#�����r��	%W<".U���d�>e�|ƃF�wƓ?�A��T�6�Wzso�k��)Lϒꄖ̉g�8wX��yP��X���1 �Be5%�����H�se�D̕��������1}�T7C�L�����,���3�W��ļ*Өb����*�5v|�v*m��k�5=5uۊp���gu_.���xY��Μ{�븘�q�G�x�H��وF�rD�tG�;��[N��Zeo���x�3�~_p����2�@+ٵ��z�P�#L��r �D��P�MM
��買�uھI��z���1�y�9v�v�\���,�@��D/���}BA�?�]�L��kć������DKJ^�s�d��X4C�8�	�l�e.-�{��T6� �����Y��"
t�M_`j8��p��&���k�V?r�P
0�@W}1ڴz_�����u�!oV�Yw��{ݥ���,L�K���c����G)e��� <��2s�n,<�q�J?��)�&ѯA��"ngC��8���|A���Y��B5����c�[2#Lp�ۏs ꖟ�4�mE��>����?�> "=����\��7>�6��b��M�!��	����Ϥ�"��OM�,������=��r(�$ŵ��qz9�j��p��o�z/���?�P�#	Qf�Z��Ӛ��aܲ$�t.�Z��A'���B�ӱ����^��`]�q���k5A1��h�DFN�D+���p��j��[�v� �(�����0_�!�ߥ����e�����d*�M(ǵ��˵C�>����#ؗ)����#���_!��xi��Xh��!�u��nz�����/�}�)Y�N�K�[�GVFhB!��2�4�J5�_Q��"37{Ԯ��	t�R�5�:���Z�K�yMy��b��|�����o�yp*3*`o0K�p�v!�z^pi�2t�6�+��-��.��A�j��4��r�����u����,Fq�#��*G��)�T�v�.�F��.�Q��d��
֤���<u�/Y<���y�S��	�`Өҭ�	܎:(N�hIq*ϧߙۯV�2�V5�AfC��������p"��9d�ŁI@j^�M;C���?O���Ks��.�;}	A_(��s	�ɻ��~$�
w�VRQĥ !�κ!�x�ד��#\�u�`nx��ڢ�Ib�qy�#>|$D��2ti3�k�����YvÊ���w�G� ��dȂ5N���������yF`J�c��s�9����\�����J�����O���Sh���^�}�)-{��;u����!��J�d���U ����H .P��&_4�T�����:e��	�(bT<N	~ÿ�d�sO�(�q�4�isX�L爩� ̭t鏋��;7w��xNz��7�*J+1�jJ��#���V��]��d��ڶ��H�5F�f�v��R�X�Z3x��������x�Z��R��_���˶�9hnl*n�XӚ-n��v���]U���e��67�aX�MQ�ɞ{�i�H�u-�1�Î�AA+�a�W�	��F�B�]�/^��1~��(�����Q�GF��� ����i0;�0�T8��>{��댄o�"�f%Z����|2s���.���m���1�8�x�Yyzt)2���w����X��ܥ["{�����	�n@��dU5�,.��/6�����v<��o�K�P~J��l/A5��I+X��p�1J���*$�:ئ��TB�t-��aZd�P�K:a	Ք'��p���k-�[�Tɧ�Ce���I�����m�����C���dWtT�{�j��E�0j'�_2�e;����-����I�����Lw�������A��D��M�~�j��"����`���>�m�[�)��>����ۋ��/�?����][N,hmK�ԩ�m%U6z�i��,'M�
�;��H����#�x��.�A�HZ�B�1`�5sH -��k�-�R�Bn�ȰT�[�])���V�$0�QŔ�~�P�4Kl���u9,B��l��|0z���0�5����=��H(��c��R�0{=���R�������i�Y�3��o�R����W덆�,�^�x:ż[6zG'�O�	ɮ�A/��c���	��$39��S����yqą*�;�3��HKY��}6u{����E���6��D��X��@�ATC�h�� P�G0xz�b�X����?��:d�׫W�� m-q�.'T�@�Ox�MÛ�z+������x�n�n.n���>[����h�Z�O��������,� ζ�w���{Db��mEP�'6��7�n�}P5~�e��0�?h�5�WЮq��3?b�QߤM.�K1�����$C�ȍrnw⩑Ld�{�c�5��߸�N��{���g�N|R΄�y��,&Q��."�j�nK�7O8b��A�(W��?���b����b��y
�eԙ8�߱@5m�OO���}�yM�Nڰ�A[8La|�J��q���o-d��������l1�%�B����� �5�[t6��JR�{۞?��2گ$/���ݑGI*A[>:1�nC���8,�ߒ,���'?�#����4��l>�CvH󒪼U�����Bq;͂�8��=���9�̲������o�B��;�
����$:�a"ڣ�)�@�˙�ޔ��I�� ��rA6a��U�Ua��B���ZB���G1z�c��z�ȕ�D�C���r%�։�����Qu�Ҁ�5