XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������V���Z�U��]H�K*��R��&�M;S7.z$�Ǒ�t@I�y��\�ǰ�Z�����d��diZ���fnGb]���t �3�̣!�Q��3��O����=BS#Ν��_��D�[|Z��
��U�K�W�ֱ�"]Eȶ��J��1�o���T@���<I�a�ԋV�����:��Lc����.	3%1����\�?ƁJqG��Y�$��!`}0LE���{��gE�Q��Jw�S�C���]��g���qo�Qr {dAq��
w�U��Zb���.�4��:/?D��gD�Ѝ�7��)��4r��'�s���8 M�hD`��M��Ji�`�($��TO�g��,�
.�h!�}�����&�5�F�M\�[$�� �p`�a���?i7�>�((�L t$�(�r�/	�Z
p�8�/Z�[��*B?���'?��A�R���%ak�Y�qhb�(Oag	K~����['':cot�AU��=�T��2��#A����IX�?���d*�*���#tBJ�x5m��g�m��N��Y�"����p�J�N�A���ky���ƏU����ԨS=\D�-��!\c�m��&>Z_�^�f�^�E�q/�j���q#c��e�퍩�@;XA -��?��(M	��y�}O�%?�碨�Ȓ�?�~��IP�UC��;�h.X)q��e�T��������Z^��r�[�����(:6�#�hB�MPx�l�%�o�E�%���p�J)ld��D'����b��z�B2XlxVHYEB     400     1a0n�i?��J��YG�.j�,8�s�/AUIR]�����<r�^�m��?����e��J��rr��o&�oJ��P�B�,؞/c)z�~�'y/&�kϤ�&�ފ	�N�s`u�迭��aJ軍�Z��Yr�}N0�'��E��%�;0�\�U�� �k*3��M�32hn�f?[9�t�N�/�l�A��&�<e>%��Ȝf��$�1:hm�|���v��d�O���`B#C#����m|�K����^���,c0�P�=��fwϽ�~IC�(r�%��Q�����R���sO�X	Y5З�-�'��(n���0���r$ ���_h�*Ȯ��8�*�d���I���1�*1�2M��o��U��S�$L=�W�j�ZsP��~�B�# �/i��_+������P(wB��L�\⾭;5�#�@4XlxVHYEB     400      f0�	Z�;,S�u�2[��8s-��.�`"���Ž�&�A�,�x��7�cLw1<9�	��C>n~�E�Vx/僌�����
��ט�էٸ�x�9-��J��s_o��`�Pw|���r���^yX9v�wu�*���������OD#�.
� Y�S5����+Q�E���z�����S�~_�?����IHF���E?�m��)"���ȥ]G-j�K���
"E��^��XlxVHYEB     400     1805)�\7~�M��I�v���(o���'��3l%o�Ʌ'��LR�V�/פKK��S=�~L�,�.�L-^_|���f�`:�m@��E~Gr��D$|�__����r�3��������e��.I$��%k�uc@������	X��|C�Rn��jb�����n��xf��aet���B��Z�{��O���ڃ���'����O�1�.Z;�����V�=I
#~��x���JB�x��#(Aq�	���ԉ�t�x̆]e�㔴C�ȟ�D��/��
H���5�YC�d��*c�T��	ֿ����Ψ'���G�3�u:�����6j��?Az������KNXx>
���D�;�h�o�c���E|��{x�	����H��+> �Ie�*F5'w���RXlxVHYEB     400     230�qPڥ�r]˯t{k�$[l%��7�����S�e�U63��f���e��\ȸ�8�ޑ TP�)�6x?x���i���bB����QC�8�F�o���"#��y+����ܐ�����ֆR1��R4%�������c��:Y#�S�B�3&mP�����Hլ�����*Tyk&EZ~0 ֐�ԕJ'GT�9@�Ą5�2xCg�`�KD����KU9��p�č�ʍ�~��G�!�e�����+Y�K�K7M�����B%@�	8_�pU�2�$�-{ j�3�^Y?��W������2���aW��� n��Laj"Y�9mbH�̕E
���:�-�ٚy�q�?��r����ªk�����Dxqg�a_�|4�R�)���Ǌ���;;;N���<��&�6׳F�F �4P�QF9篲�< $:�O��E�)]1�X�)h�1$*�D�HΉb��$��CJ9�
3�,�ї���Z��ݴ�;R��␙�@�&�[֨j��ބ��Y��d�jH�]��Uώ|�5s���6Tפ����â�c?P�r'����~�Gl�̀��'�XlxVHYEB     400     1c0p����g|���Ɇ���o��sy�r���l�5RHz+�ԓq����	
�F��k)	���G��&��Y4�0�?瓡ʞ����=�s�5²��ZJ�ET�w�GNN��Bǁ~�W����Ϙ���)�wO�L�,@���P��	:=�u	�
Ꮼo��wy�i�魆�dL)W�8Uz2�c8��#����E�3I���foIr�K�1��mS9�� �՜�Y_!�ds-ZT0��*+Y�[N�Єq��|�����{X�2V$JE��r�Ap�?jA���[������6���G��Gy ��g�z�n�j��l�%k�;B����RP ��,N���Z��l����~���	 ��b.��YjVk�5�ն=����ߏ�]S��r�a��)\��5��0�n{���,َu�`��=|xr�PuHD�iT�dȪ�//uG}'U��j^�XlxVHYEB     400     1a08��RN�N���K�d3�e8"���lwk�m��~�������G��uv73Mv��Z�{�I�u4���2mGL��[���`Ϧ2V� ��KS��!�4���a����]�_f;54��AR�כ@�p���Z�ֹ�x�Q[���K�����x�`9	;��^��vQ����m����v86h�p�m�Z���M���$�k�qq>�1�D�y�݀�!�v���Qk���IX��F��c�ۢ�]�P�!0!a�y��b���X��$_� ��jvV�#[�`,E����݅.���f����W|mm�a-ڢ�aI�����k+h�����7�Z�y�f��u`	hwm���4��8�?=cH[]��;h?�\�fi2��4a͐� Z��Tn�a"]�4�3�d��,���3 �-�S����$XlxVHYEB     400     1a0Mru���	�"{Z��Mb���C5�˰�0���`J`q�z�b8�CQ5�˿&E�T�G�f��Q��"�T�[��jh7��i����b��A�%�Jy��T.Ƭ��R7���e�~�Ċ�o�3@�S�[a(NI������K�`�P���5w�^���a��<4�7R�[׾�7b�b�!G��$�Vn�����"8���s�f�ٍ� %�S�X����d��>����C����!��mf0�\���XwC��U�;@�m�=�7#^	]�����9M=��dB���
�Lr�qY_*gv{��s~o�ޅ,dO��2u�3�٤���7���@G�Ϟ���y.1Jv�[�����{S[1i@G��������= �?e�H�9��Ws =�b�h-X���x��3�}���j�*��h���:�XlxVHYEB     400     1b0�{��SJ�_�DB����*C��RR���!��^v���U�I'U�+Ш#�k�VZ�����ԅ�,%�}�#�Z+�Ny�[z�_�n�?j��/L&)�D!1u9�yc1q��s<@wk��``a�7�����k����^�����qe!��q��]��o��O��E�r��Տ,��Y+� *9�̴��8U9�s���u���U�<���F��a?[:��'��?I�3ъ��C�Qw��*�=\�(� h��n-F����yc��,S��Ǎ|#��v�tL|�KHB0�p���(n���A������O�RBg�2 V6ٓ�H������֑�Ѵ�u�+��|ڒ�����⳧Y�;�~��䗜V��OH�}i�f���$^����n� �Ӧ�>�����R%��3Jۜ���k��HO������˴|�	G=�XlxVHYEB     400     1e0���=�W�ڑ�b�����@4x���*M9ĻWGL@g ڞy��@��i�LAo�����ζw����(�<��B��h-����q��#V��S�V�i!7/H�D[4�R�6��>ωY�I��CFv
�����5�AuR$�o�{3��P��%��n'f@��$3�X٧�@!�kh������	իe<�j�7[sȌ�@s@���۱;�A��4���(^�5����zPQ�uH��eJ��D�LyI��\�^��P⋒�N鬋�昱�IA�N�Ƈ�(���i���+f�h�%�����O.f��È�->��5��e�ܟ!2~_~[��WS�t��<!�����6�,d���0�K�	�kKk���Ӎ�)�Kx�{��N�d���z����ٽ�J�$��&���˦���-�h��	ʖ��"*@l7x�8s�f�^;T[�*ZƋ�ö�i�'�a]�M�o�K�sVOXlxVHYEB     400     170n���T��`w�"
�M�]f�u�Y�d�wq�w ɿ7�o����̲	P��64)=^��uܒ�R�<o�yتL��O���S��;�<��B���9��)gBS��[�L>.��w$��m�M�����r� �<(�_6��a��{�mG��t4i���Nhh˞k]��ؑA�D�@�vf =���h`�1�mm	J5�0j�~�'�p���AG���Bt�4�ˤ�C�t:�Q�|��ěv"�H8��4Uj����7�o��g����vS*���#�Y]1��+�`=9z(���f�鑼p馇M#�Y�����5�'��2�ÿ�Aq`��e�)܆[����k[��2�'����T���ko��a#��XI�տB����־(XlxVHYEB     400     140����z;�Ґ���V
��9k�y}Ɍt�x��6��������"��-<7��=�`�^���p�a�3B�4��?c��%����=w�+U�	뢔Yw�Zo��c7���_�]�*��|aE���߶��Z�Y�JNT�~�gtóJ,����������I6��J3����Ljnr֖����2Ju�Yt��w�#|`�^����N��Bw�z"C�j`��^������Vм�Š@O���)eճ�Do��$��wS7퀶��/+�$Dp���_��^���z�i�e����%>8,#����^��Q�Ø���,���2��XlxVHYEB     400     140��OD ����h��p�e����̊�m|gR����o�/�~d'����r`�T���ٴ�^j@i�f���ndF}��w�G�`힢B�K��MZz�F	Pfx`CX3����<J̔�ʏzr�$��8�9�ȑP����589�u�"fXK3|�k{��T1�b0sE���)դ��>Snm���W�A����͘��Y��L�{l�t��G.�����#��NZ���� ��E��R�}�#��QL��8�[�Б���8�_�,<�MHit��s��O�tDH]��4������mp93��+EK<���+�:,�˳S@=XlxVHYEB     400     180$��������(�ݼ� ���$Q���x}�#�w 
����	W�iu6$=g"G6E��W5��O2��7����#���*LS�kX�K�ݰ�����O�!ծݪ7��T����4R��ɕ4�����E2�Tv��į&�?�2�i���:WH𰑤5�m��a䅘��3t�\�·�}��ӟ�p��t�BV����uG�Oh%,ȵ��߷5U��,Z��� �b�������
��<��L����,��i�����;Np�w�;�%�Sس��4���ޔ���hWc$���I�Dz%�4�b��-�"���a�姲ȟ2	oFb�TAi:r�)фN���-��(_�;��(��IbG��gd�ݑT�{��qs��-$YͫʾXlxVHYEB     400     180���o����<s�ޢ��w�R�-�%��n�|�/�� ur���g�2ߠ"�O�ȩ��74��2�=u�>�H}�A��g�qY)���4ګO�2`h�e�3P[����	߫�FF,`V
g�������7��<�0���01��*uzm��ے�pʋ��+�Xx{�%%h$r�~���ȉ�y�q�
!x�� �aQ�u���~ڒ�%
qHЈ�a���	kF�d�z4��k���c�m��p���g<,����ܵd!Dx����ol����iofӵЍ�i�5{B�0�w�=�4L�M�x)�D��6Ͽ�\޸�˨n��i���%�q�f�:�6_��_��ʆ��5DH�,��G��,���A�}%��qp���XlxVHYEB     400     180e&��tZE���E�.T�<�U^�l^?4]�e���1�,eS���ԝY�X����- ���_C#J�r%C7aB���P���@=�������ˊE�#��J�g��m_D�C ��X�(\�+��m=�=��L�)�
�/*,�Q��W��	���t0.ޫO�(F����ʙ��Z`�a*"��0g����}�)��>',Lp+ ��<G{'a��� ��$�R�?竎 7�<�X� ϺFk���K�Z8h�R��Z�=��B��q�:�R��]#�؍�K&�\ �-El��?OW�N�#@,����&W,t	�N��w=��G�[��$&��x*3�v@�䨑m�y�����iO�0^�����>b�> �գK7�QbXlxVHYEB     400     1a0#���Բ�u�4�N�g��4M���ר����!�B��JC���)=��^S�v�W';z5�p�r��muO��W��),uk��ڷ	�N�z�Ԁ�����B5�S���>4�R}`�A��#�"� � �����H����(#_21H�a�'}$�ؤ1"���6J�7���}�uc�����^V�ݓ��T�Uu0B���s��� TN�nA����S����޽à� h�d��9��c�>RX�]���J�Q���K��!��<[�b�|7���+��'ߩ`z�n:>��X������[�ͭ�mN��c=�q����ϛ���9O�-)�kӴŅ&]��M"�'��>5����*y9	^l8��:Ҿo�\�7*��8�Tf�a����.�AJ�ZU��n�pB��![�K0�nb�XlxVHYEB     400     1a0���80� /�QDǑ����~{���t�I�/;��#&��2].Z�0�ׁf��M��^ۇ�H׾�N�L�v���������Jf_�ģ��0Ե6�L�Y���d[ԯ���ղ���*w�m���=�`�94󢜥kZl�u�;|�ZvbՈ:Wg3�ȭ�CFqJty��5�y�����I���]��c��JH����-N�:�%��V�,� G)���&�N�m���uP,��/���b�Ui
%�̨k;Q���V���׎��	��K�Bu3;YQ;n:�`ZR-�^�����c��O����#���Ϫ-���a]����wQ�g�V��[ϖ���}�8�,y�*�ܬ.�Te�/�_:�$A��
T��u���S��Ey�0:�hOg��צ�y�;2"�߁q�b<�m�Zf{W���VXlxVHYEB     22d     110R�ɶp��x��
�+x�G�����q��9��|�N�r�y�c��ޤ_=�]�7����8-�"R}�G�Q�^8���컬�I���Y!��~���.����[����cp���(�0�ҠBt�1�G%���Ľ�a�!��7�;�+&1-��@�]�5�f��T�B�
�t��a����� ��Z@��=l�VR�����ݝ���V�v���&Ǯ
���J�$�{N�kqG�ȕ�e��v��Α����M���M,е��k�j