XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���k���H��;���L�~{�JC���q!����u�O��O��a������촂N�__���π�h���������uR���?0b\U��R��GQ�w�ӏ�����-S�cd����n��� ��%u��3����`x��`-���v)S���������0�<����n	#�?�D�;K܆ K��A�cd<�[j�z �p�yI�����.�\:>�񨉙�m�����\C~���:��{���C�c��E-FB{Xs���V �ț���X����;��Phv�	
�꫌_�s�7K�b���r�YY0�e&o�*/�X|�`<S:a�~��z�,�2,��*��l����ѫ&I����F�N�?A�.���17�K��c��������J���	�UH�n��S04�QS�Y4V�{��{�D�Kt�*Ґ�����xz���%繆�7���	>p��z�z/e�ﭿ��W#yޞ]}{_�� �#@������(80 �f+�;��6�vu�[h�,��"VC��7���=EW��J�&Řv��Q�tM���7��E��7L՟-�{��`Є�����˙d�%��NPF�+��y��X���ì��N��&�*N�߲w�`�X��v"����Q&,x���"&��f��EP�M
\���<���x�`�Ħ�Ա�
t,J:���և�+K#߳#��~&�_Wga�J�*�v�4�Y���w'�%���M:C��i�E�SUD��PSLI&�����\-�,��^��� XlxVHYEB     400     190_+Z�\1�W�-l���Ψ����:���:�Ny�Nw��M�8��¤���1�rs/��;	>���/�m9^��I���S�Gr��[��������Ò�
l��2;�d�oI�E��ه��ӓ��z!;���~�K��V:f@(�ђ�/�sN��I�#�E�ƷGQ'[�A�	������K�R��H]�����&-�>-[b�s _��d��jÓA�p~���>��_�Ϳh]+G��7:��Hz�p�63��>���:U7t�g�4���4	'���ET��|�A���	Pf���Q�O��~}���I �a�W�<��W�쮡�tD�9Z�/��Kl�/F�?kq��t�b�w�O1���P/:�x��w�A�GB�R4��2�E� D�T��� ^�XlxVHYEB     400     140�H5Yc��!ݻ��J�ܙ֐(H9וgs�OK�{��;f19EUט[��>\�(�d,z�����9E���t%Ǆ�*)r=��c�F>���Ɛb���M�����L��ev�4��.�b� p����"���:ʹ#�p�5���h3�_{�FP�R�qA�#Ai�Ӂ1�k$z�3�.8�������c]���5����ZwǤ���=��و �l���6>�c]�:sj>��>�hV[]`����K6J'��B)�f����I�)�rĥ��RxpM���,kT�G��Fvّ��WP��G�;���X�z1�0�����2�XlxVHYEB     400     170$�Ɲ*�Qp�o0e��6$"�MV��{�a�=bJ�Ɨ,��fAN>�� O�c��Y-9H\�2�6,4V�<�uD7E�$fw.��#���Z����㻖N��"����C�ub�Vm�-c� ])m�jb����W���?�����`��!퀰��|={;�ɫG��C #>|?��e�C�T�
Ƅ;]mT[(g��;���י�m,�����#��LZ0�u
�0]y�
��![���P	P�+[<����Qͥ9P����/(��zJ�=.��� ��QP�lbIHg�vl���������T���͋�.�h�[�<��l�ӭ�����(����5`Q���Q�Se+�<W}�S����\XlxVHYEB     400     130�%�k��{���Og����� �p(���7�{lc�#���-\����b
]��AP~��W�C�o���j} �o��9���O�J�bR�8(\�db:�5�m�"��M������x��;	a�w�? ��YQ���+�A�bũ_�d�Pǝ�F����z{�@Ȃ�^\��m`gM=/ZO���D*F �
���> �_Kx)�\��������	��$�Q�w���B48���ul#����k=����X��m�1�>ѐh�Y��7B9�����Ʉ��>ȁg`��&�XlxVHYEB     400      d0���� �\��UR���8"jq�����.�t�)�wpćB�
�l=����@9�aĆ�������d�0�aJ-�5�1;�k�eZ������� �+���[@�An��|z�`&�����3���4	b��b��1)���5�69� b\�7e��3 ��$Uv8��V��[�3�h9د�T��C�vX@���9�����f�`TVs����e�J�XlxVHYEB     400     130�l�(���W��%�J��U�.G6>�����8gRƦ%���˺*^��E-�0K1���J��(7���_&��!¯y���`����� ��p@=�f�	/9x��g&��Yt�!�|���Q�ec��h�L;��ixO��	��*(�)��w	�\�5��@���ɚ����&�ŉ?95>��/sH7�cC,�5wj�\�9�`�=Q�g�Nﶀjl���/�wEy��#��̽����C��l�ӿW:��"]���e�g)�A�b��H`�mVq�M5��\O��Sx�������E;��)�XlxVHYEB     400      e0��|R'�_,B�k/{����'sU<��P���=nt�]�%�h�T��!�����1��9�N����Ϻ�,Q��E��)/h/bP�؀���i�|�w�sw�9�����$��E9��0�޳4<؀�����d	Gm�}ܫ�M�_$=������5]�(�ZV��)��a����k�ߧ'P�zd�U��O��0�����G/�ȧ˱�Ŀ	��"�=pà|F�?��0B:�XlxVHYEB     400     140��RIvY%g20#E�W�ʛY���k ,)�/R����ٺGշF�qv?:i�|q��,����-�8觴K/sh���Y��,��fLF^`�oY�
$�]��' H�Bpk��b��3{�������6!��k�ZYy�N>|��U�q�ð�5�q���5C��e�?���OZ��d���Wo�����DZg����N�f�w����E�P� ^�=�B�ųz�QnQ����;g��!�(3Fʆ���2ީU˄<�V�����`��`�F������B�α��=�LXo��� �p���ꀔ�Ns	��n�PVC�Q�)K�p�g%NXlxVHYEB     400     180�k�{)�BJ`�ߧmӖ�C����R�?l�����\[5��+��,Y�Y.3c�g��Wz�Or?i' ��3w��~3�:�;��\x�H����
�y���}^�BpƛDH��m���4c�pIa�ɪ�$�����ҭZ�L�)ԅ�����|��`�H�'����U��������%��TA<�=��Y�l�jP��~�z�447jH���Л����a!����R����<��ݿ�5T��_A��s���Q¥.&��N��̟�����`��v���;�2@d-���Hg�JN�nHU?MfX��Bދ��i�FNh��c�uѝWA�i���G�;�c��TYj���W���̘���;�k�*��w��9�(MS�XlxVHYEB     400     150���|\10��KW����r��m��@.*�o؎$����E�R�w�ȹ�~�������
��@���&M;�jva�M;�����~��.��'�aQ[���3����F�q6����ώP�=�J�FX!�Uג
O_�E��:Bb態l�$i^���x���Vl��IF4c�T�@���F�x�=D�+��ij\\�Bͤi��z�wN�γ.ɨ��Z�)an�羏$+e8bѷ�z��T�V�Ǭ�R,a�=��Ю[�J��nb�Þ[6��2f�C�aSI/�U䆄�Vu�d���: }��a�#����.�c6��_��*ֲS��Y���[�Ne��XlxVHYEB     400     160����U���XA���b2!��C%hY�/~C��Y*���+Ԁ�$C	ф$�y���~\�B�
\����Dp��:�kv�/U[>V���`�o�y]s���A��؎��Q�d�]��&fv��2m��H����4+�ϔ �c,�� �b�}
'X&<�����4 7�]""�(.\U�9@�*(��_����#P1���������6_���M�u�M��<.�ڻ�S�hRFZ\�G�I�98���/�*��E���u�������z�����
�5t,�NmB�#�]7��P���'c�$d�g�_�i��(�S�hN�2�5/����/7�=7acZac0�nx,��^�K�=���(	�XlxVHYEB     400     130c�7�t�'O]�a��AsP���K�{h�+Z&I�W%�HC0J�T
	�{f4�w������U�4^[�� ��"~r/<.�gɫ��p��%"YX,J�xl@�ZuFs��N%ZF��E`N_�'^����jݘ��'p��'q�;��kϥ|6S������H5a�>o[�k�i9��Cti�J�E#���:��;}n��]Í@�,s#q�~U�7ڭ��#� A�Ѓ��T��tI�Ut�G�n�� ��9�|bJU�4��hv�mY� 	�_���b�o/Q����\��������]��3\XlxVHYEB     400     140!�q�9c3�+���l'��(��� XtB�e'�`�?�Q�:���cV�Z��&Xݛ,�K0��o�V��ZjUga��YT	Z�S���z�q�����|�;07��\T�.ct^
_�{�vvH&�L],�ްL�_��=J-t��6���lr�[I�.�/5��������'&�uH�Q�"~��If�*�t����-�{�q� ���������V?Q>4
^a�,�L��yI�\��![�� u��.x��v|gƧ�����+� �i�##ݿB`��^C�J����f�������O�[ـ�GH�!��I:NՉ��3'�XlxVHYEB     400     1a0��n�ҥ�Hh�c�H��d��y3�:���~�Z~��.Zl��}�rg�Q��&�V�ȉ��B�?�I�W��VNd����F�YVBM���F���3?����-�1��a���s��,!7��z��9pr��	��O��w*3x��]Xⴞ�󇍋*l!�S�`�J�K;��hC\�����Gf��D���>Af�����)I�﫜���`[�%��[�q�/g_�&^b/lP�?s�j��&�tk���ȱ�3:�;+��q՜Z����!�$Q2��b�J����g��b9'�ZK�^�t��o �PǮk`_�(T4-��Vx��8�>_��8����o?��D�y
M%�.@s;���} ��F^`�협AT��*����g��$��R�E�;[;�BS��̬_�˥��L�EXlxVHYEB     400     120�է�;�L�BK٪����7���T�=�Jn�SlZ�&�������,S�^�F-,{����yF�]+���K]��}2��2�)(��s�P�@#�]�œ�.q�H܂T{�`�D�t����/�ᮞ������?�OR�w����sA��IN �~.F'<����:�B�jI�FI�7��5؃D�!GR����̙�/�_Ftdx~�h��Q�f��ʇ�dO�8�oF��H����N���fy���(����UJ�Y�7f��@�{a��c� ����E��o���XlxVHYEB     400     180�dbTH���P�X���3+����Fy1���F���Лڵbl������GC�cVqxX�$kO��Ԋ�^)L;	��i0a䣋2�� 9�1o��*t����*�W��`���'Tf���Dp�d�<���|�;_=���1_S>é]Iԣ���RӾqR�<��K�DZ.B|��z�^�K݅,��6`�>���t,ͤ)�`t��D����uS���T�����Q���4fi@d9Z�أ�C	�6R2H[�;������$��RJYad�������#�=$2�Fk�����DC3S-I�=���S!���Z�A��`�v��������x�tlz�}U��a�
fd���t�����e�dG�f�9�b)��tTF��1�XlxVHYEB     400     160��	�G�|"�=u�Y�Cd"����3f�<7N�)���o4�I'���ߪ�j��Ȅ���n�֚.:�k�6߼7#%>eO�f7���&�]#_Ҏ��D�)dL�����ʂ����ek�'��{ s"�ռ�Q���x�Ec�`�G�dga�U���Te���2��nua�1���G�I��`G	�>ː*E$��]���A��t9�h�m��*�ZZ�ݟ�#�+|�B�oV��Y��f�͗F���Ӊ��ԯTL��A�k7�!�-Cf�]�����M;8�2`�]�w.J ��Ⱞ.-CV��͔�2����R�!I>NUD!�8?-�PЖ��\��.�F^k���^���D�6XlxVHYEB     400     1b0���;���	�AG�|˨Wjnh��v+n5���%���U��6���01�c�a�	�NJ[Q�)zϿ�C�0�/��bq�+<�=%�o(V��Z��W�^��\�Uie:v���6W�!�b�Qd�m�D3�L���gJ���3|�����1E0�O��C�nU�,L:�$����+��!x0H�>u$�4#eku��D��ly����h���j�F��2�̒1B�:����ؤ�wo8?�)���R�8�Pߚs�5"rvQFQh���/g���b���M<�q$;ŉw p��5́3A�|�o�f�9�J���M���:����D�QbBA�Z�������ؓ$[�:�O. =q��V6i^��������e¿Ғ%�~���1��E�Boz�,�G�e
���UڷHio�#W@���w	��XlxVHYEB     400     160{�u�a���$a!HQ&���=R~�0�����Eꠙ�;�/l�"k%̨ѡ,�,s��ڕ��k-,f)�~��CF ����҅Y�D���	�y�g��F�=�#��#���H;Eo�@���Qdxְe���>G�\�p����ě��Z�`^��3 4������°�&%�]������ř���JWdi:Y�p���wa7�SM=\M�jM;ܚY`!����_�X��V0 �H��>��C����LY9\C^�]���M���͔bTe��!���:Ҋ��_~����^�o�܍�j�j�j��8�f����r0���t��M��ڰ%t��������ک��XlxVHYEB     400     130|sro�K��ь�ی�T��e�	S�\�b�z��Cn��|k?{c��'�`-A��3�ax~��g}Q_'G����þE�+[{d]��yp�-��U��ALI����#dK7���	Å�1c:���z�U�5�Tl�Qz�T��A<阯R)P�4(�R��3�����z�\����m�BL���^2������dV�dHM����NK�_i'��C��=�&�H�`ε{����,3m15�oe�7mk�XI	�Cj��@_����ŀ��Ƿ���}�P<��h�[-Z�W=�PZ��LS+W��*F��XlxVHYEB     400     140���]@���L�f�3�6S�di����?�Ҏ�?>~�͞)�?v��S�e?X��MHLv?"���?��l�*���GGol@3r��.�*�Q��a4����� ����#�۠������cv�=��FQ����1�7��	��kA��=X�:Sp�gV6r<Ħ�O���i�6�^���0�h�R��p�9�/lMbCͣNk�A-���e�Ym���-M�r��א]�o������007윭�@	�/���k�d��m�lp��%�kG��yD�&2��:�O���c)t	�w��e�2�=����:�����ɜ�AB *��XlxVHYEB     400     130�8*eo�O}��!B�MR ���˙c�JYu�՝�K�ҋpU�A*���+Q�.���F�������tO�x�_C`=s?��5�U�'`�IM�I�l���oè`��m�
M��g�`�vr�ӳ�C	9"-�'�����ϞP���3�����D#�~��������G1����Op�+�\cYM�� �ȟ(3�f=�1������f8��ڗf;�U'��0����p<]_�m�`4K7����I��]	���@-[8gXK��2�L�d0u�w09�Jʝ�D���?r ����XlxVHYEB     400     140KS�O>��p�͹>�Gx��/Q@8
�&E����n��:���^�@\dO�o0$s����Ȕ~_w��.|q��?d���̶c�����n'�g7���	^J�91��s�<�N�D�SМ+�ذ]?Sm��mٌ,���D�U�B�?����-GC��bEl�/�ː�%&h��
g�'����+��1�(Y��&�7��3ek��O�<�D��^�������3Ƶ�h�X�;t��x[��/N5'(Qy�"�k���f�fG��[b\	XXр{[<����J{C{�9��8��+�;biԌ�Z��a�dE[DzM�:��AHLk������XlxVHYEB     400      d0���dfIX�_��v��d��B����L�;�����A3��c�mwuW1��u�˶�/[X��H
����b�آ���q=b�|�E�P?��-h�+����\	�4m;z�;_�]t�;��Ptļg��kR��8O���&�N���Fg[,�<Q.��9���S[M�x�r�WѠL?���@`K���,�ȪZbs�CQ�{�95�XlxVHYEB     247      b0?Y1�
��zr������[��%G���O=��
��q����8 $
P) �@��M���%,&�������`Ra����CO�m8��J��H��
���y��_�E�GXK�$�j��&����:�lT�_çN���j�K��Lz#T@Wm�
�DU$�1�NY��Bp�C