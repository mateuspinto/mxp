`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10640)
`protect data_block
vMdcSlQIV3QcrmoyijFha26B5TOsRWX6/W2OMlq8CUyKqfhh9fn+QufI5HItVrCHDPehgZSVOlyG
LIP1TDGKqtK1BQbgP1e/Dnu9K68Op4aWc9lsr46JBkE+63mjuL5Sx1/fL+92LALKRVdBeLTEmBbR
L4x3OGOuxn0aDyzvGoiea7eUddXtfJXkarjhrlRKc4Dr8oX8pEP6S6Qhhv9cuAOk82Yr2ccA+kB4
+j4cUr5sy/yOioLVx3/1xMXzf15+twEWFUgWbVBk9akQ0KBuZQvdO7mofh31PZz+Fvtvu/rfIrDM
6UBCxvOSxY2BNm2fD+l6mImpK67MUjEP52OvzzKcwJItGNVrUZ6KMjRhQqqji9xcHEm3vu0ECZy9
vBQDUFGlK0nkuG32RiP4OsoHSGtR/12FdwttTc3hUk0x/ms7+DIPLAyk8F3G61oO4u8jReizcvHJ
cYJmoAMYqsl0MGoBt5oeRE+E2ANeV3HAc6e4Xh08JQD6MWqQLfZi70k0DdxrLv/xXFiACBxYLkuI
d15tGtTvLDWeTKj77yXjvr4sGi6JQC8ovJmgRxT7Qt5d6e3uNFTuB9rykzzC6QS97S6b4XiNQNkJ
5QqbX5qoELpWAmvIxJhmKQ3N/e/w1iEx53Tjfwy3d/wMhg4BygEFaZZ3iZb5R+F8vLBaFcV3Z8rY
GyVBkrOqncbLUGwZ+HkrldXV1u+RxbMOjNXICVirI87vf5Xbj07sc3L84u1p6bQ3tXR75GgY94+y
fPhA6r1phN/xgtezhCU/I9hjzqemDPgZXT7ARXIo75WM7CXfPVsL2yifYNqMK9aRHO8OysZ+4DJz
nQHbvDLwUealISsVRF5bbjhlEmR9mz5aQSnShyhVghzA3FtBLJrXjdlSykWT2ldVVkDwTelR0QEP
iuhl7i9mf1U9NYOKNyhRQBvHVvyIHBi2EvFv5BQP08fPgf7FKXpy9hfEpZQP0LLD0kPZV4T5eQwr
q03oP3kAb2wxYguguQWb/yCKpBkPQqIlj11lc3OCtesYjMV+AI5q8To/DMJPaUVKfhvLqXGr5vEN
9hxwmTWAyXS+p0SDrpJdjBumpQlYqb1memeSc76P1s3w+pWA/ogRSQw3dbSWOgB4vYkCwNLi8f66
ZdP3i994T3Dc/HBlXj5zhF6E2dZNwQtUxNfFL5uvF6VZp7PEZK7FWtSm7wUhQu3VDkhj5aph0mh9
c2bldJRxdVKPkQse3/s9YI5BFR+K2aOK2cwk9T20HFeqsfuqvhypYgXOQua0PJYuYnDlefXRN2C8
aB9qgH5E1RF5TPiHKH4SUfOV7mYHX3vFvLir5afRf+t3FuazLZF6qd8GQJFE+0yD435XF2OADF0I
5blnEST8sRxWkfbNhqemc7c3NdlMAHP3vWJ2ylZtGQBuidOeNzfLbwvgMX/GgrVt+lfdBknoPhkb
9RL0Y1lvjbK3cuiiZy9SnZBqI+WTdi/eTEFlmz8wzgm3Sgh+P4702p5Wik4AYBrdXwmmbX62zNj2
7MPZ4sQx6+BD/BedbRPjJyYuenJIxFaipE39ROxIJpvMjVJkc1jGbRf819KwIMOuYWPScJvjyZTA
nRLWgvcgEudmaqRX70KA75E5J/Uvzbf/bPsSiOc4oblW2Kr22cv8bhl5E2lLQlR3q3ObyX5nWkjy
oANnkKmi9kBHmtxeC18BLQ4+caBmQJkgcqBQBoXpGJmooUdhqCgvgF8dcM73N8kzLf2R7OjrTR8J
1j3+mwxXPu84qYo7n8Tn8z7ypD+7r0a6CfYrNrAQgzhjPt3wYWDHoP2PjCMyOTJ3EuEQrfnirO2c
zgqB0bbsQOtuAq8rUZKBvC9ak7WrR8oBaSvlUnlKw3ovoUI/Ax18wVGYvXXZ6iNwBfYqeJ/TMwr5
ncTAMZXK9gjk4OHA5hcef3+qXl8AEf8ot0OQ413V7Uc/MY0jdLFmc3RZF1TbKpWW83/QI3DhUSR/
2BS7/C6mS4Lmy73wqk+fM+p1LNktSWluYeeYUmNuhiXsGZ/+mRfwN00iL19nv6bZ3NuuZT1OIPC4
u9qRTx3IkcHUELhuHy+bQCpQwwCrow47LcYKmsWbfgH9LuLV4QUtj9GhgM08pLAQ4CNN1bMma7FU
h/KM7VdAPQV24lNq0qF4z3vYmhCk69xR1QJAhfqMKwFzkgXfyVfDJDyeuaCbOLhbWIfBfblzkMOM
zYXws7d2C342qjsABwZkVOhzcfolwXdkWCE30Myl5LEyT5RAfccM6J8Lm+0ZWTxE0WrNdMbxxzgp
ziDJHihH5OCMVyCr23TIl+NpNBHzcodbQPc5aykPyCfmhKLhQth938EI1VkPXiMbRhcvvNvCsyOy
9Xvogfq36LOyu5Oz9bguhZUwPx1dPEI6UwAyJXxAreqHB0fzkou2Eu+ejeKp6nt3Hz29FlarnIho
ayDai6kNf0E33D9M7/LgPXKCK2S1EMNmGSOordzEw97GQAR0+x9v9yt9O0UJGfbzyIoSkqeVz4Yn
pfW9ire60BaUWaUTwG2G58jDSRTVP3OTNfK8g6ENr7OFlqOW5d9EHqYOQrY2BhbnNVX5Zui8xuat
jOm8nmGeLLpuEpdH6VFN+sEUTnVENaM2B8zmGgDstyPZEQQqIKIFQTuPOkSNWqrmy4TWYxH1Iz0U
H+FTZdcUtPc4BziYrjLuhomp5+gUknLGguygmwazm9aHWna/4NFM7QkusNGY2NIAFwD628zvGRNd
wh/KV3GtBvIKG7kuF26BtatzI7g/yo5R+deDMdefIS+eXeNf77jpgTg14gWKm93dT7XT9Fqk1nLX
96N/JvVauP9VH1mfTMcu+YuUN3b63BJt8z6OTYB3AZsKqhrQVGdSHLTB+DsJzn16ezhQz4B0HoBd
z1rFXeOlTrYzTn2QN7puwRzf01YN78EkT9XbcjKKrkhlv5DATh7X4KhiYZq9dreWx9KlxPjFG8qO
XUDKGeKF49LjNtfN4SOFM3smrW61iFqIkCoPuArWBZkJxlp99JigXA8dzog/Yh9hobmjnZNt/ASv
b+LmHsCs+WziAPYGbfLXFXU49TPQqDKgEoUA6WTpQaVdM3hNj/O1gx2tgAy3t2QfuJNKuzL/wFZ5
EFh+iiZwpHAVmqCXE5z1JBrI/BquR3JyPnLQvsQXbx6Yh+j29YnuKE3Db3X9VMaZTeZhcIBoFHcp
/MLW1I/+VC/WDK2fvHQPkiRw9Z3Qd8l7HgLCkowQp+OfrmTVkKxoC+wzbNaEgVKD+FD3IIzSaqy0
PGqfcDe9WcWr4CG3xSXm01SpLaX5gRyjA10DsRNuMnZ8y0/hMcV76Qa+SovMiqNON4xR9O5UgrMh
aeghyHZxwy9v1Tlub1ZMZ9sbb14BTyDCd26CE8+tDn+xI/mUG5TQ0Cz5q+ZJqg+zTIguRA8IZZX+
Uv1QRJWssAWRKA7OTmNUDApWPZsLDMP8zmmud/9TDPTypekdhSApvriQ/+HZW6oZ0aixAYcq/JI9
Ipz+Hw5LMxhEbFmIhcUgCDSe6he/mK8i+8EryssmZpOpFoeNkqAtaTutLkRMDTpwuQZ2/UVMSurw
FJ3Ep4jrpLIDZxydrRMWkp6frcDFnrpBP7V2LEYKHXC4LIBsmGsc8MY0YmTmJFHBRsmr+KeRhSKG
vUqhO0gk1QB6JhXdT4K9bxX69fDVgkhOysqvrHpeIrPm8SP5AAa0rMbSCXU+BjvL8M5X9dA/VHrF
Pk/vj111bzkGtfo4jt+kcc0Vn5Xu/XF/wbbxEMqYaxGYp0uVC3LtWhRdEqVF3OiejVV/idXAA7H1
NZ7cr1ugYfZfGO2wE2y/HoNjbcNM2zgHc8M6Rl2zW+BbFoB0BrozziwlzX4HmGDddpvbQELdJ5z4
zpz2mw0ZFkuVGv+NW8gW21SxPmEkwfqfPvXo0qOfZDe/FYBkKtTH34mlvhMMKVXhCiVqToqLCy+j
pMG0h3eyQXh1Ov1xbQL65hGliZzEIH4dhAWDucfFpbOawD6s5dDD42vaJS4pYGgr/hjSHSO3/6Tq
9JiW5AuXryuprPTJDCOqQLFmkRF+WEBRKsWJChvNXwjFsMzwja//3IHQTaDQCXqyRj7hzN0pcv5x
amB5j3jYnXZ+A2gE0kRy3gWw2Gre26xReLI/LaIsWeS60bhH7L113WFEmHRV9XbxbP45Dt7tfB3J
VGET8Bnvm3oiftnwl0IHcTbiHU+Q6I+84cVdQAJxJcaraAsrhKgKCteWwa95QwF3pUXID728RolH
SMDT4sz7eljsjXPGpiEDhbwBSVTGQUO/hPGLbfs5YxlNThT9f67QE4VsI3wkJ7ohDaI2NjoJpzQo
JPi58WOEyfsC9Az68esnFnhpmCWPEiw8hTyOLBJFLsb/b0ibe/fE4u5/vGrqi9R81hZywH0HR7Aq
bY39ypcaN+YZD5m+An0TuSLtJYk0MuGZe7Dh+SdFJVAfGHM5M5u32Rei+1FnfiOdn80u7DLfXNIM
EZbvpfdC1q3TIHvfxJx69CoqqI26+g9mS9rYQQgUGJrKJDVUwk1GVS9gf7ICi2q86pW5UMQarQoi
KZbsdtG6jnmfgxcLf36BQvrHBaYmDCX7lHY0gGUh5WCy3dr7tzdUa1dqLaW8ZswzU8bBY8gFBJ37
wFipH9Opli/lZRhaZquXWa+pFts84CQW40h3sgSR/Mmf1PVvZ+PLt/ZUYqSaGUroevNBcZ79gMMP
hbebo3Z5S1lXcsZawVfsVgaMm2c02EJkeYnzn4b2C0nRbBNFphVOQKEWsSsRHc70WbpT/L0AHNxX
trKAHuH++GuOcoJ4Tu+F7RZUfZ76CI5RYPqZiqfebgqpr/q4UX1DtUobglLQEQh8OWa7gajmiaBL
62cWO7c9nwed9PKBnIzMMZ0B92X6F766seNBXixQtQT6LFc+BLUzrNee8gQ7dguJFKThJoci2EqZ
CJJBeHIOpyXABsxltPWiwsXnS+JjMPlou+I7iF9KjzbuRU/8S+hqpZ6Q07opbI1IPiIDo2BOFfBb
1OiR3RloecMv4MQRlny7JrsLJVETY/DQOFn/OaaYxMHhzaNZXn101/MIi6oHgsHhZFlVllPTeZFB
T9+YWGnb6M/Z6QPrNfpSXIJDaf8M333TEf+VxE4jnaLlsaqSiz4q1SQFaC/osc0cLWi/xztAtyIh
SFb6wuDaFMSBgJ/Zrwri/T0GuOVGuamH0OG8ioOYn/uM+L1D25YbZfXustFFHnzFAW/yLvuX+GJa
KOMshQWaZRum5nm8kGymmr+AEydfD42tMWXRHX3LYPumxciXHfQRw9fPIEMWYkW8jCPFsSxzYrSH
wMtX5jhresX0A6I4959J0AelbJv6oeCfhGMNx+A7rKgNTGE0uokLFHHqyFwAEC5mR9NeAbFP336O
J+G/9QvwJwVjouE4zQsUCwVSPV1bA+5gah4zZYIlNxk69ixGQZKqQWH9QIoduwvu4ka2kCrZg648
zyxsNLLAk+hgLOh+nyk56KcOV2iaonL0rE0gAYKnkFest/3/8m3UbL/CM9/w0JWp5UCgH7oCD44s
4xe2iVZEe3IhsBrcFSHW2Yt2/54eGIVEaZJWNecYMGzAHpUdLfEqtKcUADO9qTX4tmFe7UzLI653
VhusF6UqnD40GwTImJY0bxMNjwhnZJsyR8GRb3uBTIjoPRM1ieTXOk1KY5n2G+A8o44ofLsNvIXh
FCKGaVkd6UQ9IINSpqW+jB18DKy1QqyEbBgFTxdDl1OVG+mhSuMgE1l04WfFZeIr8Td54EWowmzh
SYLu0dRaF7eSBnbEEliFnGj16gyePPE5dtjcfD5dkCxh1F9Fi+L33Ls6OZRAt4/moWkkc1DSqSvp
C1aI1rG8RTu3aRrkhbnjF9UoS+lLxO+a03/frQ8xr2kJrvjyBu2fXcdvze/bx991F0oJbJnNFg8D
TovQHRCO26//U0EP1KjFn5BTDX6jid+Hc5M+rwItrBNyqKkPZCAnR1ORmNdI7vMRFAdVnwxQ83rg
LKl/cIN/x7NJ0qp8O9IDrRot7if3RrDR1rKd7YYeWhs+dNyWms0Mjt1kO3TN2y4ubf6LRT0058aR
YtWa9iKhnBBLl6LJzWCAPjDV5RyRrjt3BjvsZnY31Gqo8SVJhaVyT0ghKRIMq6HVBpKE+Odhf3xG
Z83nURqoSE4gQgOberhmkaZ9YoEijs6qgQC0rmVrCCnf2mZ//nWRXk6ILygzoq3O0Yv4GlyeDYvB
WRzZ6u32jZtC+z5OCVGizd2xWQFhWnNJtb0hTk3gpehg1IOT1xCgtf9+yWDxgkv40gCXx72ISELA
RDE9n43EgGcpRmbjjTDtmCdubWO+5NGhJ1JAFAl9LHi1yPYOatbsanPcPGgfUbPLhpvGBm7yEjso
nnY6fj3CYRq0u17sqoxZct0BKeCXNIye2GlMI01q6sks24lvvSe7DnWIhASzhuNPCpiAg7pfaEb1
2rh7dL46fUDNoX5En9FxpbY/kcoDJAu/AlYL2ghLTolhOvQLqX7n4hR4w9qiv8sWtoBdHUxoRMHm
HOmWZC75ffHHC96MQd0tVz1ATb+8MuMLHmwf7lWt3UOlrWsNPYChPh7uDzhPohSm3f3cRHhrNJB8
bhWnWLCbqjk7cW8Uk9A1F/j2+6ZVx8G7tOlwwuaw0C9f62XSNOZJaPz0oBjCfoysMZfy0aHHSB8s
bk9tmfttPoUXqjCz+hhqeBSGQHB24q47u3dPlAi6I+KVx9cQU97GuKWZSFmtKIufApKdyQ4Hm8oU
/eGuQGiXfyaplc1muTOzL+s7G165Xu62hE1JPhG9WpHnoPbGhVVCILT5lnFshLtVjxKlvWALjPPC
ltHQEZjW9C/apFAfls4irW48nYO2rDTNZ2IyWz0J6GsH68OQCrzteXwE8Dtb4jfG7AqwnOLJolR5
+RTCYwKTyLxy4lPKzbk9/vFKDujDNNcNIXOVzqHD2X3xuJ4FaTvgaKvDd+Lh8Bys4T8znjpDvGRT
JVcUZRV06hcT+FYhubkDh3Nf50Dxql+q++u8dwsmpk/bRP/MvB5zJBGnrtxOGIY2w25wrFJcfoyC
KnP9IUQpaW/Yo7MItujKY/k7TJJ6kh/JO2KD1mt4Ck9/CutkwGlxwJ1kQH0Z/R6gnGB5TsykcePR
CzENQ0wn8LpNm6Upk5YBepfyRvIX7S89JbO/p7kSxlaDYNWAy9O/c3lRhuf7Gf/l0nhk1UmJllrz
MUJby5zUalEpCcRmpFCWzeFUAbFA/I5fHajgBJEDSw0o89hwXnGfSdbKJleaaIS1lOdJZpRKHIBm
ORGbv1xJhsVep+XjXZNGH01noUs6no5GIooQYn0lgbqOELAmNLajNi97lBW9ZbNL+aJ9DISVp5rk
YLoNamzrZ2fW/5abyP7lfKWNIKi9NspbCsCrUe4deA8c8y74ResBsEb158jinhV1LLYecm5qZNQf
8Nj0XByVA+pSP6mm4q5/kKMeCq+4NatTCRJkngCEZ3FAWyZsI0IFNA1Patiy/nP/p5JrrJ5Gy9Ur
MlMqYQDFCFZKPNmNXoS4suttf5zmLAZ/UWok4AD3pWHtF2SzSuurAyXiElk3dFFHLl6c6LbqtYyC
1rQzdzJHoPdYtJkut3U46IkrplIUMmUqlBsraoMZpRrbzQwtm1DoU3FsHFlrh2Oz7cpBrpzDqeHz
Z+hmZs8cEvxnWVZIBftEVMYtSmMyDMIu2NMxaLriIjqY1T71ngvUvLEWkWwGvqQHNSjvoK6RjF/x
W1oFutgJ7gHTp1ADiQm5uajUVjiBV3Yo9/W1gkHAFTjydvX3hn2d3HnjTp3nTkyeq3HTLy9tCPd3
jFJZ2yV0msXEPU86bJREs+ti8gTgDb/F7CMLYHE2boSsE+g1lBJJ4sjNLQ2TeD5DVQMgM1gyiQ2a
CDZB6TUvNfIkQk3cs61gODHXJD0429DOxevglIhc/0jrbuBVQG/KIOsFlCX8N1Yzm/T8qiiXTeXv
/IcpZ0zIQKQfSgTxZqM6UpEpVpAhHL9RWs6iw3Yvek0jRSDKFi64BjP9yilVSyOFAtNgY67rQqrC
/537mVLu76F+8BDjhFfyJUToIxnlT47Mv9q0nYXF+wx1D3D1qzynm5WA48FHQQ2K6Xji1Nc0uXpT
H+sqYO8nsPvyX76Mo8LhSeBjALXyY02Zc2TTbaGGmgBbynI8s4IgsSQ1NJohGM7j2cCfr+1clsP6
gqCUd7jNv6h0wEEPz9EjQkk98f9zA/qelmRla5tHQTIORO2dh0zn8fTiRL0xKOImLWcbC3GPpBgU
jq96TUveYtBEXfYy9r3nu4O0YiNFz75M7e7e+SUjjy6pKbY/gym+m8SYtitNydhn+a15gkq5OkEs
tiWu+7wEvw84ujgfOoewY0J2Pqq4412BSJFlxTA1DLtyTGAzt8LBtj20w6y9v7yy0Ndj0nnb6KS6
dbY5WARabteU8T6zgfNsAeCurekQueIzurzai9NKlSZEr9F9OirDXgfDtAn8YTssHy5sm+19cqgR
Z8nIvhp6H88PiCqESSBJB2iUCSETspfh13T9LErU2GwCUeVhn2cGdm9mSATHf5jThbOM+vsoLb9j
hOQVXzv/E34/rVLr5RLTSLrSklzjcvcb+4VYJK4/DePreG4SFSomcEE5FtNzTHQdQVTaTQdwugT3
bX2YwI6pH2/cNKkst7VFQ6xckvKNCMqXyJalYr6mnRBHx8XTX0oZ9RjPbFRl4s3gmLikQPtbRYZO
cCP0DL7pEgHjZK4hBn461C98bICmdpCGPs5A2fKcxuPzCzIdiN6StW1WQmxRJ9YN1uYDSUigCg1f
9ewoJslC0Pgxu7K2Se+oDSH50cyyv3WYPM4MjQWGdolZOUG+cQlXvNYIcnN6xKYJmAZy05zZjwNv
lHGJtMZLb03326yMVvGlW7pBq6t9FF/ifW9TZSf+jqrns0nb5dh0Hfz+4MouVJnfZUsDfkx9apkG
eDkZH/pm6g5/vUF63w3+8QVxBHI4Ip91hN5d+wunCEL0eP7i6FAQYsWQ5aZXbWUwuXp2hah+074Z
C9p+TnNTr7MUZarsovDddI7DlM6+P2kOU0APXJk7vLU2gztyyhVc2sUOAlutzf5hyULY/9fD1Sot
WMjnOHbhw1VGZfia5eO/TXJL0BFuiloyROKgW+fvfwaIiQi9ix0PbtHP2PuXzGxy3FUj6zJJrwo7
MMko9dQKZOR7gH0+sGhmmnmzJBOGFC9/mh2wb8fcNZ04GWdgYlkAjKl8doW4erqrHeu0oUUevbrP
KdJ/RIOumVF8bTNNBtkDTu8cdon/m455WjtyfJ7staMw0DWWtmBNOhsCajnht8MJjMhr3yakQMtx
4Z9yTEQQq8RC6Qxu8tYwq7oCxbV9ImIXpvpacvbXITeBbUxI/XitXgsau9gDXJ7x2E5zAwW5FEM0
yvGyy1Tb0rsvbYETpKuK13N2jTghLL0RXwSww21//aBBEbiomcCstA0SCJ0TXaUrJK21ckSzHN4X
OMw03N194SIQQrAcDlixZk8Ml9fruXjIevne8KvF03lYj5rJSG2E9xnR3ygp2yu+zF/oobTXwToC
SNqWHhyYRQZDAYTphcSzh3/sla/C5W2S7Ml8rpxHkT8fEp802kRClydbbMFWdNVKcBF4NUHuD9Cm
GlwYduJQQqmF2ASf24mDrbGML5wGtjVqpxBSRjV2O9j8cvJ4GZcSU1QrJHOn5RMfCcdTwX7bpQKZ
xcB2QfI3ogEYa/xbwyG2B0AkyPR7YEVzgfGgybjOAiVnQeu6I5o380ICGk5zMcUE81Fg7YcGNFjT
OhDFbw8/NR3NSL1r4XgtFlQTVnlknnM6rrxybxXpmiTuqdFqaMjX+bzSbJxdMtXEQmiRM90kGMZn
+xruYIZ7Heh1kYYAwqktzTLQvAMG/ch5p6/olQL1Agh5mwuCgupivGjQpDis7AmoXi1Q/IdiJL8d
4eIbnfpi38clM30fbSl+eeZXRXAtSK3lObN4JuPBra4MhmLM4C8Kof88j84VCQbNDVf2f9V5LnKq
eMedmuDpK559HDQ6rinkG8L0yac6DHxd0SRWo0yqTuc/e9XKkTm2cN3JWq+2EH6HY0e3/MhiXVJy
k8kbULEX60i8trghgbAJu/JfwcJyWFqA/HRH243UuVFhUzXodcu8Qb2rIYFO56kI2YYSbhhUwxnB
CWxHzns1cWW8pY/k02WF7WAhFM7hwt8flM4F0Gmmc6TwNtMGYFh7UrSZx2DaRCOuSvmLXe17Lur3
El7R4HJJaG53rU0Ba9JdxTEiUKAZIWMy/pEeNbItufcIVpUxLNmCJYJTBKwI4vgxHYRdzzdhEm5/
6a3sw4vlxlMn7Zm0P9lNzxNisPkhw8gadnVRRcRcFSsDjOzAG3kY6QeYuiyln1R+epeCzvJJudBp
TRqSKREpVO5jrpX3B3U8+i6wCVD24raZ7uBcncSPKzwEAU10u5FibHksdixM/z/ZKqLFXhxkDIvo
q7mclg9ZV2+QEQxOdOMd5YCJ1WvlCdG+MqBpR3vdNDPjQACLXpc8K8Wp/IhKNd0gniMACdGi6xPS
hf6Y9vIL1WMwqM8WjHN5t5B1DsPr0Hg55QxCAbwbCLpq3RKj5WxbAYr7K8vV1Q5sBCB3qHor9Vue
VR6DmfogX+hGs3Y1XySIbc7Pev6cLQW9zfrXPK+q724InsUtfotknWLTq1Ji2uPQ457KenL5OLGB
m/F3f/GcWTJ6oehPeqLjWobhcJWkiwbYM+TGN8Kr1WNUV5HWJS4kwTMga+ijnWcstOo5xqmyOFM7
NMkcayqg6deVNQp/bkeVq4bFNwEkkdy5NrlRBr9p7YfQQbP2nokbu4SJhInoXbV7kvEXf7klvSMK
Cr8uVD1GkWEc7jZNyREdz7pzK7bWFhygOjWsGJQwHfTrVyet20jZgQe04woBUN3nJnR3psgBeF9A
DflfvOCQRtzFadh4r7nGfFPmA7cMm89shhgFLVL67voGXLoQCztuWt0g7pbP/v/kardggxN7pUri
jP/AnZcqSrpAyHzx7MBSTUcskbdumMaV+ToGNCvYrTmIPpu9WbbNmmM9HebYxIuOe+ZQJnCkW98W
lsdRGht8S5ZaQ5SDi69dEVHdQNwTqNnVhfw1kzjeYWKbZba2SterKoM290NZeuKwfmAn+7mdEDh0
KngoH2h86xc63WcPhGy5Muzk9sX1W8jmLJF91EyKizeSi/kKNZYV5X26X+2DhGaeopQ2e6/dMoL6
iIOqa4MgmstelyjYIbUGyvF5AqeCkNMWExH8NTP+PrtdpMaqsR55p+RtIVeSsbJ8tEZEBJgExw7X
Ve1iqcOdyYG4FOm/fhi/SLepxvYG1cWHim5oShv7NB1hm8vYAMX9tyt6qjk/eRtNhHlbrpmXQW5o
dfkMpgMtbKW0RAfKx4XE2rRzuspZ/ekXuW12Z0G4IJ4iEx15d2DzURqmye9n+DGWAKqinwRJxiRw
526nnX/SS3R5aNydD7U9TFzsTFbTBsjQJgVIyLROCvRd0wN5egivhgmNSBjT969v3WqC6jFPPX4+
x1+/u0VAYn3XO3RMljGHMa5F/ijuc6NqWyeljJJy908nUyFN5gizhDAU+b5PnBWqau5WjjmZtcfw
x0ZLMTNEB4C4bD9eHCWlYxAyuXbLCdRFEmOJLRXefAnges9V9DKKi9m19i9Ra842Xj7ybluJy7a3
CU6kNnLvUxayuozFW7ci9m8HP/b24EDPWWQjX69Kkzacd8ajTBvFCzGZYzOpqYlkGcgliCQkHHOQ
uAmelenedq+hlj6vaQXQYtauNAJs9ALnfqZA7FI2n9IrW7CcaTmc5FA3rx4jsbIbasofQDU5/hl1
oLRdWvsaPsl/Z1MGSQiOp4/iDoV6f0s1gIMJLWncSswlhNDb3j7Q6lgzHfIDE9ai1V7mhFTyVlUR
FXEdIjqgDlMgWhDAt+l1bou4KFunyHl75RzSRAyhrdXGZrSulwyNgQysZ878GnzX9/MIGSboGHCf
Z9gFGuhS+n+XxdxXOdFcNtAJ8mnpnsunPY2vWQWiDFsv7nwLiW3bGragbUJGV5+4esqNHmxyYmoy
QFIFpIgua3m7r0ATgo628+Mx5NYt7t7X8UQmPitZ04TDxwh+CzP1nqfGykT2018qtejOZxsA9Rzn
woYPMaZmQTxQJtFfLG5YBhoCI0TMUMQ25Hu4gMEPkmPdLBZkzFiLFt+Kp14UDssXE0HBnv3iOaaS
FQubQJdjcuw0JHSKQ4a408WdydkJGKnHs4/m9BNztV0gh37iW77+YzRP93GmF99teOP8rAshTkZy
R5TrHOxMphm5SZDew+/Im/a782S3DgcgjnLMSuJeIRuhmEBqARk9dWE2gL/pGl1eR2/SZGh/Td/W
do8kgbOkFUv7VU01HIdkNh6e6UgAeEg2NeWYP9crrDMcBPPukYisxZ7tEvNrUKe782BTDpM2csYU
e+prg9zaw53RIaiec/gGQ3ozucMG/Qwp+2wDhCOGHcQTbnunjcd+1nnimzbI0j1Uba6voB2HEyT7
n5lom8EZHLnltApidMhiZfAgSMVrjWCqicy4OmdIPaiMQP3vw3GvUP/mUeiUxorRwz7Pteft8EJS
+rsOvsmrnKjyrSV8tglQeksk4W004VixkEZ2kmTmPhcLZgHlQchiKSpwgBBGlDug6kW27sf5pI+a
y0u4APVrFL/T7WVqOtj+kUu1LDZ0V6vmca4eQIvfzd3i/uDO82GOupa+q+6rwXDL19zAdxZrKkCG
Ao9kZIw8OS98clsmSmWxdtONGApZDvFRjcR1kMV9OB2sFrS6gh9Crspm+4Dvy3tvugLc8GL+MOVl
29xKmgCqfakGwiUZ45F7Pp8AHG9l1D87XUPs0THKp6tWx2T6XFqNmlqx3DE8GhPEkPPUMPrX+DAq
7doB/36DeFfBq+8o2dq98l/g/pAXN4KIu0T005gU0WH5bBumTFqkdGdufofogLU60cTAMhkdIPCn
RVK8TfdFokKvEVK5ijot3eTE9BiX3DOFxT8uPUVqu8Jiz+XEDJIgglpQ0IjrNgkoX5Se6mLVwhs/
tMTASyLBNHTCCtDirI3AVkUUYxVDjX4UK8g5YkPo1F9G3y4mTY7/vL5u6hhCG0DDD/jqTVa5PGds
hqKwELvfUNosj18qSODlXF3eJY97iSXtkdJCAZ7U/E33HpIulSzzXePa2rz7xQFbNir3UpRWcv0H
/tcAyMlrhjs9o66gupZDNTf2w58KiJWfqTgnprHfx1HQwlMM5EEGl1U0EWOy+NuDyxQOuEzHnGM7
BW7aUFdo+OeD2oSL3KRu0OlVA2ymCGMT6A6YmbvlROkNx+9bZ9HAyKOKYnjvS+sjRbuKoFnDZx84
dfeYjqiO34MwhtMc/9ToEq8ZZqwXTPPTf3DYlwMcAfvohc/zJKpZMGhYMzaNx2U0K9S5Wnh9+t5U
+dG6JpHam5mrnCHQg+Q6GaYJCz14t0bBghU0VYE4nIsnvrB3f/bDEPSt6SbBc1Uwj7mT+Zw3aBs9
4lEggJ5kaEiemwg3fPuWT2LK4DOHglD3D/hdKPwFohBJqhPlnmwLOGAGUDmqMA1WgPsU/vexXVlb
UqaHH45Ol/VvLr3q+glKuGYtcs8hyLGpuwq8CUqtIdsVwp1/80J5IW2r3Be0B7CpDkQHxuIKowCk
+ktokz5oywqZIlMxdIo227F7A25aucDVz9SP7dR1OfjSsilEcJQQE97OI0dH2xkq0XXhc4LefeIS
vUw0Hx5Tiui+HnVC9hHIzfo4YHizANt2DBrYA67NtfD+j/yIypdvN5WPCfGgLHXKFs63CpG0wayi
X2I7TyUb60EprBjmtxhyyylCNyc3HoDDzwO9p1eh5bgKuVBo9z2boHZX9aTfaRs2dpaK3UpFaXJT
I3YAflOfURYDmZgdkAOgEwGBE1v33lqhe/cQqP+5LIlSHlySbiocCf3pveqB+Y6ikfhZeE1RARfW
2NVdBql6Bu/N59lR0QY4oEEJ13dsf8sdVwzjEb9T6g4LiDrLzhl/tsJHmB1HNmzYKd/R6qy7yDM1
l04zSwOnjLwIWTEv6x5ECcyJPNTYcFuNHjHfZZ5F3jnA+RgMeZUPwHPhmlZ8jMdSPhOdXngqodvx
wzQQXGvq7QcfPVN0jPhv2PPpZpFx1/Xa1SUGHtsuXHxvIQd4jmI=
`protect end_protected
