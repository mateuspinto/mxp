`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
DIeldUrFouTooqGufzut7xRv1m9gxFd70XBmwyfCCU+1TU1eeSZiKrE81/1Whjnux+jH+lyW+8TN
+JMKQSq1GPMNM5HqYkOC6l5NLrgeLVQWKRdKLyAaBIsYqdtStZF3W5INrrlbQRJKalwhRT4o/Lhp
H19FRQHeEOHcC9hMhxwLNGa12I1qRfJuP49aTW0SCO+a1UJJsf2y9FI6pfULcw50bEh6j3hPaBG0
Dy4FbmmOsax85ipOpoSm0/V364hsH6yeOcKjX3JVbqMRANoAA1gTubNbmer7HuO2quCGAutC/xpX
FhzX5O+Hbjch9N3TQkREW/4PY6FD51RJc4zmPg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="Sb+z1SXNmK0+XcItil0IZkHQKoyXGW1l/jXlHjWm3W4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2160)
`protect data_block
5i0EkaCVUcP+OmMAzUOjW+MO2zKwJ5bGwnVrypatPKYhtkeKfAsLysQNhK3gXPxSMwR76A219xyw
6Nj8aUunhrUck4mYDraUW6azLmuUDy0+1mhi4o4aaB3GlHFPM7PQMk7Age6h4L2i6Cxljr4zqj4F
FAd7YeNcnDc8PvwTfLtnmCVlF8O4dWE6zJUG+qHvo2pNAsYPsz/TuTXcG34mfXKdTX49CrknjfKP
XwF5iZ6OQ9uIrZBEaE3qybhToOrzlqIu4JK8OL9tRRUvffvX64CmozBpvvu7y9fnkBxDMc8XeH0m
kct0tkbPxJfSA/Gkj2ojwqn8ww403o11qa+8ykpiC6ixgE0Z9Xvy25+Ne0+TOuqkGa2msJ2WFs9p
lXzhMcE4ePW5zdc5qE/iQf3nMUQqeFS5NsPjaO8Eq5d7TpavNo/IfPuiz5dSJWQtie11V1iuPncy
DlyPWIpGCxbX6fm2Ka5pdtLVFk9n6HNA8w0OGpF76JYYTHgrRqPESWiK/Qa07d1QYGoAtfNe/BxM
c/rzTv5NoUFfpIrtWu+9FiKolN8HjxwD6/x45FhuqMedhzhpbn5DgZbqYPISJe+QQRvFSTcbP4ca
fTuPQU0C8oSYqB4UuvxSKufHHvJiMtSamhFycN8Net9JIYzlP/S7dZ0TKBT1bOlH6GystHHpUd+/
o3h3gI+hLGBX2oeGAIeh5O8JVkumXOgZsY6t3D/GK6RyhKaeVgx9jw3pmUXpH5OuEmL0ZZga3deN
ArAmXWpopvU+egU7mYP7+8v4QKpZqa6gShnHAC9NZ3G0oQOpdXc1PqHTmpxcjTx68xxvjjlS5V3i
UjZJY07GPyL9FvdZxFRJCN05828W0pTV+v7klHs8uEQkjmbbJS0+cyh2uM5lQQ7o6574oCg40D7M
0XoQVbpg5A5xIT/9V9wjtGtfTJjjI0h4XD1ZNacIpVXn2Yi6Ly548uaX4hZHN5dkPL6JhMD3UBWo
dq9d2OnJAo5IPCvoL0MTtC/cSGTzSHBYGBSuVI7nAgbD7iZFZVV+3uPN4HhUo1ClAC1c3MNQy4Av
nyOe0OMpsGxT/0K7tYBx2a/jsxhhW9Qzs/2/SgRRUgsftZIuL2eaF71AtYBVfaL4ATqOe8kNToIa
6ORBqHIpnkhLpZvOKVHgVZH8wlLFANxc0rSXt0ZzAi2emWZKmBrRriHH6/DOm5wHYQiDImrlkibH
UTOw4zN8AqqMQojWtAVIuTZWffcFeB8c5TwCDqOceDbSWw77ncLv5Q4wWShjwxdi/wRDqqbmnKWU
K0VuIjoZEgpFXUSFJ0ip7Vh7UTsUjpEWI9H1DeyHNfmpK1cyu3Llvf2Af5mMC4rhji1LRCVJoxY6
E3s7hBsBln5I9i5sDKzaryADIQtOHUm8tOUQD8d0y/IJ39xEoBu/Fc/yCR72cJTZdYpGXYO2RmXj
G4ENnRjLwt9iDlbHnfo1jELGSu6wAmwbFKvEUegtgXQAOfj431HAZaMHSUrTCEsyKD4O2xN2Dkvu
ovnKBp59+/gpFP9O1cy+r2md0KNihgyGC693hogg59bNJ7R4JdxXoOh3AoBVDglXqxhWAZ8LkJfm
tUd3NjidG6h24aT5fMImF5+ZLEK9OTySz3ouE8B7X3JK45naTf5wnArcm5LBV6k9RI6PEb/gjBB4
hhtLIVJdT1rHx0rm8mebRBXCRXOQ8199WouYwM8Ak340h2i5PQtGLJqqThcVfu5z1O/aCpy0uE4v
3g8h5Fq1KEi7Yv92g2AaGXgLRgTCgURkeSxceMAJUWam63tRjSgTBEI6CVqeyZGUAgD3dF5bXOdd
L3JD3+Tjyol4rN293cn6v2asGPlw75ZfV1JTui8mHehd/hnoFPICyaYwFEsMTKDw/yYPJcaOUMj9
eh6Fwe/NK06yy5UZqhBOD9731EXwPaQlPnHY1E/XfCxz2dBpp8M3e8kch2Be7+XsQYEdhMRwiRzz
SdvmqIISSatlmGb1ylcVEoGrqzm4hsf16dRVfELcYAaV5AT1sVckWs2+F1W6PXvIEH8+INm0tBY+
P3H3/ydx3gVxKxlyfxifNOfXkeJAvmYxmvo0TphKYeVMRoCI6EFfUuZG4pxOYidWIpJsYnoA0ywY
6wBwT/YVpsVAzU9cvN4cSz+38EnKP+OG4V1giuj94xF25NV5pc67GQgF1Cjpo7na+NejL9iNjALD
PxvnbMnuA8hE441INCpN9RvrnRkRsGGvlXYixIOmeUeBz2T80G56OjCUh2mAPIpJZQ/FCkhaMSl0
QV83fdKQ6GoVkCnwJJdnVL38WrDeZOcRVgxdYFgtJSzM4eRN5s7kekgiily2+7x8NXHLVEj2y72r
5qQUgnrJFSIAWCEj5Ha0ZDDk2kSuVL5QzeEyWtU7A+yHHisRTME9RdWnjivjcJh8ZU4BLadBj3Ja
MxzstItXEN5eMll8xKjZ2oUdSUM9G/aasjG1oJg4xRjKngDJhE+h1IzU3zxKCeAihrnMaEwtK3gN
l+wDeubCts/JqDfMnWVT5f0cdBEZQ4VWKRWMhiKBor7jDC/EvBPs3O9js9G6zN5HnW/7xQyvAlEe
/8EZhfaj+tVOPkxw0zF1ESzILXOlw3cu0esgvZne1HIBgeQRiX7zowUllfJiiL0JkWCgMOd2FBAp
Ygj3MravTeQYP/05ePl76c/vlBr4POtZjYrfDM8HP9GVRfF70aD3EbVMQfOHbQeAtL8D9eE3WJZc
Fnv1AN2e1SYearwiv3MzotkmPntLyHwAOuLy+DnlaE9PRJZoEhzoxsBNE+6rGVoeg9bVsNtzZ6L6
GehPygCcIkPgC2Ir8Plu25Svxlo+CgID+1UDi0nq0PaS23tdlimFkzuuRxKif+eFFhFf
`protect end_protected
