XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��'���w�r��Л �p���S�:�p�*��L�xf�_�����Km���|��������jT*U�:߻e@ɴ�.Y�k��7���o�&��!n��	��4zy����4
[hj#ʠ�	(2��N��r���:5�sec���+0�EQ�qz�#	WB\s��Ce���y���WKAA�^JK�jȩ<��)��x���iMv�n>j
3�d��h�� W�`��y�v�?5LR�w��d/�S_����um6w?|e�7�^:�S���X����?[��9���m����i$*}�_�^�R�H�4@{� �s��9�	0�Q��FT�'*J=��������[|�DX稡��e7(��c�sZu9}6�HQ��c����^��/	�:;���~.q�6�n����<�|�s�"ic�o���#���J]7�7�$=����g/�e�p;r��6�Avj�_���,��G|��:4��J�
��Z�k<oIF�kض��~�\��sTv�?����t��n�.�Ss����e�G�4�`�P\$OZ��?�,�e��БqX��"Y��º�l�|��"5=�o*CO�����]&?i� ��18�g�^�sٚn��>R�L��|��̝����NS>��u00`�so�N�Ƽ�V��-�%�5VM�y�W�7 Ǡ�=����$c����S�/����z7^DATOc{��ea�)|��W��8����qŒ,�c�c�(1+Jd�z���8��霠��[��r���}�XlxVHYEB     400     1d0���`/�`���ϖ��cpM�I��>wk��Ro*�8H2%��DP©�DΤ$<��ïf}�	uZ�3(m?@���v�:ku�@�Ӑ,!�A� b�lᅵ��NV�T��- ��>i�!�u�P���B��c<���Uw��N̰�������k16ċ���+�gsQG�xG��( �ȕ�Db<cb�M��h/� {Z5A]�7��! >1-�|a�_� W&d]�#堙�����J=:�,�]����y���H��w�� ���F���l�����̋8���$Q�M:����sf�C�I 4/����:����ѿ���ȳdGϑ��^)�Y����ﶀD���hŌs�IG'�X�;5b4��v�o�M����hMHD��tr�ɬ��fkupK؞�ڰ1`�ܸ�Xv��j}N�w��z�C6�a��Re��A�W��ܝ{�*����m��gT��$�L�z T+����XlxVHYEB     400     140<Rc��Sn�����I���-��K@R�N�Q�)#dH��ݖ)�ܗ��l��{,K/�d��C���s����5���To�����0��� �|h�q�l� ]�zMkY��8��ѹ�L�F˓�췵�Nn�J�r��m l����`y#R04�"j��u�� �N��I%i����3��-S%���{��[�{a�,z�l��5�����"VL��◱d��.��K
�z�
]�u�hU��|~�!X��;�|"}.��-N�9�a@�a"+�����NRҩɚf��!�=~�->~�ع6���(�TU�;�T XlxVHYEB     400     170w��}��v�_j򔡘*��y��ݦ9��sJ¢E��ʾ�WN �0�Q�wW�_�tد���?���!cu��<`���s��*b"	C	�y �tq'}/*'eN���B�g�X����%��O��*U�L ��>C�21��,8�v��}��6���I�5��Wҍe�2�%��xDy�`R���7W�4(!l�[Y�9{P�W����v��x�/6,�]�-;�>�F�u{��3��s�=Tc���ҿy��*;��5��!G1pp	�s���P�\ф���)s����Y���׈�6gѡ�}������T�0�4�Sl�*��7ᅍ�G-iF�j6��1	���#oP�uB�>�DK�V�*���?>O������XlxVHYEB     400     140����4�3�|z�� 9�{L�#��x�$�-!�	�gIhr�P����΃3�����Lo#��W
oB���1y�Eq�@�Z!>lw�W�
�R�n�r�z������f%��,K����3CM�H4��cYt`ޫ_�3�zlJ8H�x��S�����*��^������F��BgNӎg��]>�~�	*Dۏ�c���n��e�R+2���Qy�f2*�1"�6����cQ�����#�����M�Z�k�����Hb��7% e+�E�?����3+�W�/(�P��4}MORi,�C�+�8Xד}���K��U�~%m��XlxVHYEB     400     110����'��a�C/��{R�[�0ȶ��Eb~���e����]�v������"��e
�;h�*�^s����� X�i�BE�#k<��vRG�|F�P7�8iE�m}/�::v�cP!9��!��%J�a�%
�n�Y���pΆ�X��~m3Ǫ�<	��|t��87���џ���\O�딻��d1��c�t�1�[���z� ga���G7۲<7�E� ��W��Ѱ�-{_�V�~/x�n{)��?o��|�rZ��cW�݊�8R4��F��&�,�XlxVHYEB     400     120�H��4ز8�1�aΑl��[��jo��]?f�Wb\r0�8Uy =c���;�r���o���]�.\��h��n�U,V5���T��E
�������4F�4��ɏ9vx����n ���#�f��;��_�p-��B�"�[#o4ZbJ��s� ڢ�^���h*�C]Mg�L��R�����,_�n�b>�<F-e9bE1�����EPAf�U2�Sv^HΥ9�/$_�=�� Pe��3q��6�ZAJ]�qdIF�A�\/HN�p*�@d���\%,�x����|Q��XlxVHYEB     400     140vV�ź]��;�f�R׷��}�~�����L5��:����|��bE�Y��yow��>(�9^�LS���gr[]�FtY��h5���7s� ݦi��B��{�xQ�7ֵkq�x�q�T�JÍh�LW-ZPYd���i�|��m���H��6�����ڙ�U��
8���Wa����W�(�K��q�4wZ�K�C�C汹���)T��<���<1���t_|�M5r��8�	Ҫ��K���g7�fk��YT`�u���jw�|�%*����wK�)�����VOt�f�e��0}��^%@�#���O7#b��(��XlxVHYEB     400     150>�,��m�?|�ݱ�ܺ���l�R͟m) ���#E��b��Jj�]��K9�c����M�\aU΀"�v����!b}��Y��e��:<�SHN���Y����;�n�H-����p$ ����{|^�pЩ'�����x�3�e��Ǣܷ���:�ZO,l�2*U�l���o[$�w;+��\8ƿ�Q}3c��G�t�E���,�y\�E�	U������� ��%�����Q��̀}�4)E�F�Ґ=�1�0�q"�ҍB��DUel{)x'& ٔ��C;s�D$�w��-K�~��{��6�j�[�U-����aSc��փ'�F�M���݁�SXlxVHYEB     400     140�3�o��I��nX�!��7�y��$O]mV��jz��ޑ?4'M�~i�g��`*�YO �k0�|K�>��r;����4�y�K�n�9;�
b3s�[�&�>�߽;Fv�֧R_&�eQ�cQ�W��+|��h/#��`�8�H�����|��ߠz��>����I�'�uo�)���!�ўr%�i?�@Ev��ӽ_u+Uj	!c����Ϣ��fV֍�#".��G{K�t��Le'�^U$fq;y�l�ۅ�޶�N%WjD���헾�sɟz�qp����������k7����qHw�� ���P�]	�ܫ�(8�XlxVHYEB     400     100��I�1������x�H^��}�]�F�udi�@�:�^(�O`���S�ǌ�k�;T�Zt�R{y���p��ؔx4T�x�&�=��(��Hʪ�{���~3��#�Z��{m���yrx����
��V��]��U��NPG���)���_�*�鄊qE(W%t�`�a�di� �*�&k�u�U�}�?����"�Z����r$�F'�331Q*��s?�'��KM�@2*D��}�B�ٕgjU���h)�p&၇[���$��XlxVHYEB     400      e0�e�V)џ=5���ɦ��*B?d��><�>Aڵ
u/Έ>s`8^vb'�����#���Ț4�5~Se��ƢiF�x~�5 H�b����� ��<�z��}nx�+�Zo��R�`�;�{>Vn�{c�m��n���U�0�L�uW��W���\]$�"0�~���!0���`G�Q4��9j��|�P56���C`4a�$�)���������ޥA,y4��XlxVHYEB     400      e0M#�[�Qa���Ұ�\��[�|��w�M�}%���@�A煀���%q>S��_�*׸��P�`�֣$�s�o3��cO��'�dx��`��+��^i�;Z���t�����e
/zMn�<�z3�Sٌh���]�H5b.�n��1.z������1dfλ6�s�X�3iA���4E����^���̦�j���D�9
[���U�]'1�4�4)o����y��XlxVHYEB     400      e0�HΕ�ڎ[�a��J�`���Gd��O!��e�� }�Y	-��*W�=�;�ǐ9��^lѿ���_c���]܍�/���������������4"޾qT�pQɞ.�����t5��O~H3�:<+6�/t�H9k�-?�F�I�G���[��UQ����ɮ=wKs�7� �(��_�.f{Ś ��u3��=CE�~o�Գ���z1�KXlxVHYEB     400      e0�]B\څ����;M��î�)e�6~X�I@:a��Y�6��g��1�[�`�a<Ph�,x"��^�(��.���RK-?�2�L+��"�nR[��E�e�E�-��P�$�?H,������n��b�(�^ �gz���Q�Fi�`��7���\n\���R>D�&%M���G�[Y��0x�W<uZR2O~ ݂�cD��\z�/g��s�`��t*������@XlxVHYEB     400      e0U�*�:Va�U��T)�n������v��Y�km�����n���G�]@���+6e�S�ޯ(*nB[�6fO=b��\�(���Tk�H�Ǉc'y�,��x��}LV��F�i5����B�,)4�g4tEu�Ycs��t5��s*%��	 ����:9�$��"���29{|�/�3ՈJ1a��%��Ǳe����i{dt�~�2t*;����ϑY8�����@�XlxVHYEB     400      e0�p[QŢ�tp�^Ҿ|�DL�����L8��-�h뛀m`��^u�>M���[b��"ߛud���?nM�ۋ����!�����9��\]'�O��17zy_Q�%��MV��x�x�h�);_�7j���Sv��[�$bʫ�h~���܃�q|�<h�[�������az�0�?3�r���0�#gOw@KK���?/�v��m�I���}��# ���e�j�IW^XqXlxVHYEB     400     1c0<SUЪ�`Rh�|�$��Is�Ij���⯫�f	ev�)���L��2���0�n_��H�7�ƨ�������^���i��n��V9䣀0?��e��_�D'ь�1e��Z7��|�'���U�$lN���O���6�kV�b�O�q˻EV��d$���6�=p(T�0ꅔ����z|P\PD�8�̜�)l=\gG�N��*<<Ni��܌�j����:\�.�5�ϵ�*�R�[����`ԙ��TO�M�U8�(�3m����+�҄����c3���މ�ϻ�����2[�ʋ�<����a��!���7Ԑ����*|��	���C��a�o��#�E��ǹ�2a��R����L1Ca�ļ��k��Y�6��u�^)����A`���Y0j�N�8��9��J�< �+���Xq������q��"��ê�o%gTh?���:�AO�XlxVHYEB     400     1307��ؓ��1���4�r��p��"2UI����$E���I'+d��?��h����~1� �n�m��I�}9�Ϩ��Ie��G ;y֫�2�V��Y�W}C �����v��<2MEg�q
�E�&�4�/���|��C8�z�����LUkX���z�]�uSB�VH��!9�40O8�~�G��1R�Mm�c@<��ס ��o�����3�
J,�I'��Ad��S�F���i�0fA��
�E4m�I΄E������R����)�B��u�F:Pv��WҠ�XlxVHYEB     400     100�J�x�,�Ռ��^����FD|����3?�"'���[ ��vI��F\��>	�R�g 5���z�{6�X0��L.��`_A�
�����L���,��v6&eZJb����9y�O���N�S;���^�Y"�
�a���~{�/���>������,4�/]=% �!S�xo����2g:?0X�da�6�[mKe��|����#G�&�Z�s���rW���k�2�)�x���?|�l���,u��4��!5���XlxVHYEB     400      f0&5�9
�^�ձ~�АU����Ym�]8����� T2P�V���)��,�fR�n�10�F��VZ%A�~����I^In�B�����U��<���wD]#>|2�A���,���!h�K�5J@���"2M�h8���/�k��)��3��?�)�b����W���|���(��zy�� [����{B�q�NX�-&��Q��gVk�R�SG�F�%g
�k1�p�I�Up鹆XlxVHYEB     400     150|a��R�|����ȝ�e�Zemw�/�v�ж	�߯젴��(U�@>�C�r)�8�22i���(m$�tX����c�6	K:��kL���X��Ⱥz�VB��2�) 6_e#��� "�S��=�rغܖe�e1LI���V�۔�P4H �/�Xm�((�����i�w���r������a�_�B�Ȝ�xE��k��D�e Ɔ4��mkl{��Y;�|�B �,r2p��cNօ0M_��m�W� ��
< PkI��xb��6��	���5���%��[w~:�g��0	'w�ztL��2NG�$�x}=,&��ʷ��&�Y��h���-���F�XlxVHYEB     400     160\�%OŰ�X��~��*W���/�^�9�F(a��,��H)�%���)B��S�M.��Z(!��.��š3 ��UJ����Qy�A�帧/��Q���A�R�5�ŸOө�BE%͡�^�2�\�òz�3�!?������V���z���.�E��!�ᨀH7e���%p�n9��qO���i���=�g7e����p� M<���\��Kᯇm�K��>�iv�2��<��{Z�V''���|\�o�w���ɰ���T.~�&�UA���fAQlsuwp�WK񭦸px�	K{%�wb��&��������(�豷��9Ǘ���k�̥�M,,"�)��~����XlxVHYEB     400     140!~X�"��upg��ب�uR9�ء|�ȨD�jW���9�8�j��@�p�k�ȬА0�(���`!/���k���ó�K����)Q5����4Ȝ*o�TM��t���|�zόa��~�M+#�'HaJ�U��- �B���ݢ�e�n�v�'�F���[�8�_�I*g/|�꫾���*�dE�}n����"z�VطG�� ��&��-Aܟ���YX��~	z�XL݉b�|`� ��2/�:L��$+����'�kO�F[V��쳸����<��7O���jW���eg7[9�kG��k�E����f�d=��ľ�XlxVHYEB     400     150t��ڤ� ?�����?���S��d��#������^>�?�q���l$���ǽ����]8�J�f "QY�
�9���)rJ����5^�����K)�魶lh�)��?kD`"I��n�����g�]�5������^pWL�m�aˢ���޲�0�+��7u���g�OS@�k$�&:+�	d�m�w�]�{���V�u���d�Vj1�m(�اȚ-vq��c �7X����f��i�$�d!���.�1���a�����2�p�'��f٩e�8��o��UF;?��z�� �����3M5A��H�k'��ɝ����<��f��A ��bR��mXlxVHYEB     400     190�}$7'&G�!�$�z���S����*}>��ɰ�d K�.Z�������f��T�P��=M��`��T�Vْ��֪�!j��	���@)��p���6��g�;rR�
�񓈒��v������n"��Ƙ��W���D�e'E�!���vH!i���s"�P|5��2�l�0�ek�K�XafdX���z��g�q��$$��fd��-�Af4���Ҿ��E�i�E(m}���W���Z`Np�;����]NJU�lw4��٭AV��uVE�ϊ��(�bl䄼P��=����/����p�O�L{	�?
o+[;���f,���Thg�,�6���L9����P�"��G��r��y� �
�tm��1r?�»�.�2 W�F��	XlxVHYEB     400     120��o�8�����f1}�W!lyΙ~{9�J�.���K���v<��b�r~Slmb��w݋��o�	�E �yΉ}Y�)y��X�.ر�~�ΟM7v��X�1J�)�&��1!P�c�4ʩ������r^�Ќ=�SW{ܒ�[o�u%��-$b�z|�־PA���b]�5��y�E@����-=����+:��g����BQN�҅Bq��!�J� I�;:Lu���H?�Ѯ����B�����I�2j~v��f��Q��4+�|��CO��Qq���^'���1��Kg�w��|tXlxVHYEB     400     150�4���ROp�,��:�e*?��뿘1ƾk��R%Ig跍��!�0ӷ5��MBN�@�.�|�ݫL:�ɣ�6 5�$����X9S�Q��c`ŉ$D�̅W�FT�g�>A՜��W0��A*Ŏ w&��-�cf�)�',��5#)G{��9M~���!E��&=m����R�"ӦXt�~xP`��{�ʪ߿��c���!���$v'n
b������ٌ���g��3[���6�%us��,��77�91�O��S!���i�9��V���c�	���7B�ۣ��ѐ��I�6���R��YY_�Vr��C�&�KR��E��vҊʉ�B�C�Г�����.drѯ9XlxVHYEB     400     160��ֵ�*H@�W���;'���M/;����D���ŕX~�:d��5pT5H`��(�� ��v�`��tNp�"`�`�|�`���{�Z�a�׸�W��M�I����$����"%�1�v6�'g
r�68"�4S^I���~"����]����	>�4��o�{��b�[:9���m��,>/}��Ig|��}���a�6���@��4P��O�!�-V4�x��@�ez=�=5�s�|�I%��A�oi������v�!8�������i0��ON�|�U�x�5��0Th��ɷ��:�]=���<�ƒ҉{<]ѕ�C�T'4�q���������(�����f���l�!��eaOGXlxVHYEB     400     140����d
9��m�&G��3ġ
3չ�Z-���5�]-cK�Nq=%]B(�8R]���	����2��[1E?{��hHKr[\��/}����˛~롑~L�D��Դ�d(O������*�WV��$�=̩��{���$�����_�����iG�8�D=����7u�Ȣ8���6 a�lۃb{w���A?&�)s�M�n�3v�Qd�i�N���%45h+/5h0A��"��O �PWV�(��7ƫj�:O@AJq'yt�LD\x3����coͭ۩���7�[���~�~���碱�?~5Dj��b�zXlxVHYEB     400     180�oN���۞�4 J.��[y�J,�\�<P������f)4v��h��R�V��D�Y}P~t�̶E_A=�6R����I�^nS P�E�.��)���dL�f��>�F��b�ou��4��x�T"*��w�l��a�QEz�S�W��ٲ]��Wؼ�r*F�3:Μ�rK'�}�B�r�w<ܔ�`�l��Վ?q��yAЃ��"����!��>9���eU�!��:�X5��Kn��V`�J?vD�)�9*��oܰo���̥>��I7_�k wM��ja]��h�5��m�m,�f�B�KU�	4�0zSG����aA�Wڶ{>�|b�H_�	���a]��N��O��(�nf_D|b��@!H��[�e�IqW����3<�`��iXlxVHYEB     400     130d�{54�rB@��@�a�wQw�֔��xyS�@>��vD=Ւ�wv��x)L;d��O��E�/P}����͍đ�,��$ъX=��Ƌ���$b�������,�%�!�O�";ẻ߲9�d��e��<ۺfC���A���Z*��k�Йq��OqKZ��&���c��s���S� i��J�����:9��|��Y�S����	c�u�6�=��g�Dۑ��	��te���a��1�N�0��\�#��dњ`�3���	A��� �>T��P�n5+Vvd�R�qH�(����(����$}XlxVHYEB     400     100򟓳hp_L�ŃO͵���G����d����j�/����9	8�c�D��Ǣ�KwW���eY]�����XCʮ۠&n�����1���۬�����3K��^/
x�H��n@b6S��D�ъ�is��]���p�=u�S	�߻i�;O��"*b����V��38��� 2=���I9�l4�ʴt� >��\t�Nр׮��j�`=�01O���
( DR��p+��s.z�����M��yE�D��_f�V��XlxVHYEB     400     120M
��6�v���렪���/�/��CW%c���ƒ}b �)���z���������>	�������
�;z��ն)��=�j�K�����Z�˧�Foφ�ֳ\���w?Z�ң��z�38��HHź����.�.�i|�o���!:�T�fcg��P���_]x}�9��qX�X��舫�i6X�3��[l㬿�����G��~uȦ���_��J#U2�:$5��,D���|w�M�����2|=����$]��4��Pٙ	�#�E��:��XlxVHYEB     400     170Q�l�p;7���%��F(�4�EH҈5-=�ͭ�\V�����0�Scxv~6S(��H�#����ea4>���X#��������,�x��g�t�$��X��&�g��ܦ�tZr/���&X���ܪ�X�PS�n�����9P��i�2LQ�)����2�� ,�CD*�v������2��-o"�����I�g��W
��{��n8
��jp�O�i�`�iF��fgх����o��2"�%m(�m=rU�4�A9�LW�7-Cq�2�Z�\�|�
iԪF� iva��3:~_X�}�2���?<n5O���6��-���󜊬r�ON�9\& d�$�?�.hw�{«����r��΀1��af�XlxVHYEB     400     170�@�Ő�Y7pS�fӂ�������������`(�p�(��is�X�Wٖ,��Ց�;��w^&��,�_�����­�PqO|k�@�x�5Uy�y�3?ÎSʢ{�W�n��!����R��*������d�- ��y|y.a����S$
��>C
s��'����qP�*-��nu�]k9~$"�"��j�l�Ӑ�#�J����:�γ�s�"����XE�7�Q,�[
�&��JN��ΜC��%M��� t�^��ĤN�>\`u��dxٮ��.݄�����Ö^��9;UtK:�[Pdp���p�U��� vΰ��n�:ve��� YA�H:z܄��'�~E����xT2XlxVHYEB     400     190X���FX��9��k��f�&��#���JlJJF/6h�Rf	l�4��9T'�ųW���q��b{wHi�7YU�� -��	�����.�>��V�8<W�XU�8x�6��z|Dŀ����U(#3P����Jڳ׻��ȍVΑÄe����ŉ�c�<��P[��#O�3����gtw۴I5�����̳[EH����%4���;�QT��f�l�[`Ƅ��u��q�%܅��G-�W:U���Pc ��a�Z����� ������)+��b�!ĥ,/��G�:����kf�J�J�����P�����pė�$�t\(/�:}��� fR�����h�'ْʷ�^�(�-��(N)O#��w�l�]5UF�'���p�R�����XlxVHYEB     400     170ؕ��U��r�9C�m1�R��
��e��!�gH(f���1n&�
P���U��,��M�g�T�3�|	���_lⓊS�s���o�����k+�{�bL�7��Ɔ�6�����z�o��wL8��&�B?_���;ϦP'��C�c�ȜM�JA��#�81ei�M�)�. ~�/�)�Z8�y�b�h� �R��)=�?V��e�L��B�V�8�3h��������񮥽��B�}R6�y-4�?{آ��(q���`i�~)�����F��%�g�a�Q�|L��g�H�J�������Q]Ҭ"��;�>��7
��(5B��Nx���U�'���ք��B7�[bv�[W�����;�h��" �����d�qXlxVHYEB     400     150`Y���;�W�.��&"���pZ�g�aJ����C�g��r�ޱ�H� f���n��dz�Y�D�d�� �����b0��ٕ-����*0"���� �J)�8h�?�.Y��&�o�rE	^W�AN<�R���y�F�r9�jxW�c'}.V�ģ~��&h8���	nqN�[�f��۞6��U��&x�����IF�g�5�<1��ύΈ���YJ�]����#mN;ƻ��w�?OFbt,�3��B�옧�˫\M��6u+���|D�c�䤦���8��w'FA������8w�d��7ۍ	�U��\�￐
Jr�Ǖ�tL�#
�vXlxVHYEB     400     170;��蹴j*����8wPġ��>�[�i�Jz�Rm!��j7x�-r_����%ڏ*X���]K��.e�(r��Srzn���g�'��Y��@�b|H��>8d�a��T1�
:9���j��ۈ�:�ɟf�3�$5K{ �K<���e&9LA~��D�#kn��\Gd�;7�� �������3�bd�F 37�8QAڱ��-���?HNf����[��%���g�����[=|T0%��_�����Y�l𠞤3W<~��>I��8���z�v0.����'�x"8qS�CnN]��m�����#^��H�'���ٟ�W3,3+���������h֜.�ȿ5����M:�k9XlxVHYEB     400     130Qh�NĞ۞��9������s2��%����K��rB�>�='��V��z����{.A�x�������'���j��6�K�����X��(�ˠ	��A��`� ݅HA�x�B{�Y��>������-g2�����)P)�_�}�h��`"�p�}N���V7�Q�yY��[V~���RE�(�(��}��xh��.�w��w��}�T��Oa� ��lV��kTq}ʐgn\�)�������7����J
� �k��{}+�e8�m�R��eE�;@�h�&H�z��֌^^}$8����XlxVHYEB     400     180�q`r�+��1�̡]w!�X�P�y�w��H�̋���������j{�p��J�f #�	N�3�Ta�����5Q������Ҟs����\S����h_y�*#&��')�����u��2���� a�7�`��+��7�H`�����'Ĩ;<�\�ǌ{4�:�W����+��n-y�Qx���S�quэ��$�0��-���S�f����il����s~+�G�3��g�Ƈ��g>���}<�
�L�����9k�����a
T׭^��TkN��?,z3 ���_�����b�l��jk_�hWӢ���C*��T��[A'g$ ��";Q#`��M,y��������'<O!��ˎ�fy'
��E���gk�XlxVHYEB     400     120�Ʊ�B���u�rE�c�}i�r��Rs�\I�M���&��%R^Kmح�@
X2�3ˡ�N����+k�O��'�F���܌?s5|���/J�+�����&?`V�=?�d�e�%b=�#��hB7y-��Z��B)�����.���@�
hB��n��dZq��x4���K/ _O��c�ʑh�Rr�aTA�����^�}8�0�s�SڦO�N���
*�<��}Ii$�^#�{�Z ���rl<)��H�є:�?���H7��º7_"vf��.8�����6׫��GXlxVHYEB     400     140Q�Nc��������mu��'G�2j֐��~�J�py�nHE�B�qZcH��?�&�7��%C��_�{,ݎ�},Z�3C6�?۩��f?�ryV�N  Fx�weoH�k���Z߾3U�;wO�~)0��*��D���as*�T8-ٜ��"�\&6믄�z��؇����I���5|�K>QS�6:Y��$B[V*S�s�B�� �U@��y�[l��{g`���`��\�GRΗ ^B����Q��l����p�=k0&��vZ7�L�n;`��� 9�*Cy$�/s#_=����A��v�nN   g6���~�
���#XlxVHYEB     400     140k��A�I���2�-Ο���-[�q��:l������&�0�W�1-�Z�?��x9~M�TT�������a���������.k�]p�ʹXV�������p�TriṘ�:�NҪچb�?�'�rnI���c��EF7�7m�o�n�JRYv�Y��%����;MQ�d�;�Su7��F^�*�x��tz�r8���Ě�w��a�L���QJ�:���?����_�G �F�-�ښM���5�+�͗�Isfȃ���M�8�"U(�T�<�E��ĕS���;�q6���1�:�F�����V'�.ϸ����;����TG~t�rXlxVHYEB     400     180��^�������G�z�bB����e-�����s#C|NB�BU�x�"sؾ깙Y�dl)z��L���_�~�|�μ#�H�a��Fd-S��Y� ��3�A~@�����+0�x4�y�u�lHP��n�s�vE4,h�>pm�'�'вB����j��,��#�������a������z�C��?����D5��C���WP��������t��y6DеBp�oG��.bn���ư�0�D2niq��G)�:f<!�%�%�I_�� �Q���J'3��8��X�wC\y���z�&�L��Y�ߒ�[�EyR������#Z:��-R��~��&T?�=��G7��{!�;%Ɋe���hXz�C��<>��	&�}@�XlxVHYEB     400     150 �����@�\�t@���`	Fv'�i9(23��>O�r,h�[���Ga^-\�Ř�k4Fb�v��ys�dO�9g�찉.���=�n��k���j��v�W��hN���ȝ����O�gh�����H��P��po?�����	����Ț��W����Hk����Β�kr+�#F'�j!��gW��z!��9��o �F����L���s����\�>˷�m:L�]�.��4*���G�^1M���:�V�:b�boBT�����GF�ES`��8��ό���E��Xs���:�o��:\��;�+c��:{���q�=y;X���F�\��Qw�H��g�R���$XlxVHYEB     400     120V'�;[ٛ#�^hl���B))1)X`���y
8� �Q���G�cs��kZN�e�މ5���}���ۓ]�+�Xh���vEͫN���x������Z�$F(ju�aM���LT�?-��A�ܪ�j��w	E��y���?�p]GǠ�~�Kf�
E~?۰��d�i	:R]G۱�A��m� �i8̲����K�j�b���^š]A2��|�4q+���I�z�{�R	�'C�:�v����;[vg�U0qH�b���|N7�0���<�c%c�` ��S}XlxVHYEB     400     180�Ln]U�j7:}�
��^B���t�<����hW/W��(�{\s�E�P�d��F�^W����1�G�J�a��ڠF�n�J��D�����UUd�zĬ�V�%&�Y�¬4�M�4%�}��ȸ��U�v�r�>���yi��5��#�!��x79{V� o���� = �cq
KK%^��M�<!��L�����[B8�����u`ӆ�.�� � ��0#N�~�K��"��i��0�Z�1"�~��N�N�#O�r�zB%� �&�7Ь�qa-Y��]�WjE�ǙFyZ�	�Js.�K l�H���]*Tzw$���Ɨ��x4��O��9-������}S*�A�|$p����� 1�L�P[y�(N�^�z��}����͵ߝts�%Vo���XlxVHYEB     400     150���@<[��Q2ƚ�t�f{��n|iAF�u���}�����Q�%$�	�b}��f��8�#<~n�Ɏ�G�P���ؚ�S�C�ȅ��l�@�=G�àf+��uSɸuU�[�mԌ�8�[�m�?,X@g��pa2�9%i�V���cO�-p,�N������'EӾ��2���|�.T?�-V��m�+O<:�.��XV+�b�� n�Rd�9'{I��+#���P�ܧW���q(��!l�Ϳ�ħ�)%�b�b_��3�8@� ���3y���噤t�:x����p����5*��@�Z
�'Se͞Y/$�?��nFA�Ţ��Ti����2�%XlxVHYEB     2c3     120��TF�R�o5	�#�G����E��U1�~��ɼX;���$�R��x?��R;����Q"�������v�Z:�EJ�cF!��'���n�P���Q�'����J�8}L���D�P�ͳ�#��G�?e����w	����4�39���BB`���C>S���Rz�Y���a�����k5�w�P�Ɯ��n��1���b����s�!��w�Sy;�I�S�w��j�F��Źİ�4)\�����4g�����'�ϓ�;*M��	</���c���n��*�m