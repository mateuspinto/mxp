XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���+����X؜�XPfr�.)cߚ�g�_�&V�^���T����c)ak@䬑!�ң_�A紽.s[���]�Z�]�2��	tǉ�B,���S!
��R؟�
x׻�Qs�"��}�$�&�b��XB\�V�)��9��?�A�)n%�����j+��~_�g���'���F�B	�����i��۠�U�M&�\}�vg-c6�i���H4T����	(��@�}���NM{.'.�9�I�ȹ��$� ��{�P�S�Y�{��tX��@��޼t	���P
Wك��G�$K_�6���f��ED;��t2ȒS�>]��s������j�G})ȳ+g���h�˶���k6b	a����:A7b(2��j�p��{6��d�N9��;��퐄-�����uV�X�Y:\+ly���+Ã��})����+zM7�׹z�D�U��W�9�F֍2��;�%��'D67�{}E�k~,�#�_���*U��g��+U��_���S�h ����:��k��S��-�A�� w�6t�ۏ
Uw\����&:,�֓����o:�)�D�o�1���?�H_r��&�!�e�h4zG@�a|7jog%M"��s)������
-L���������ϙ8�o<��N?��g�i��~1q�1.�k\g�kʞ�V[�$� �Z�]5�?A��'��*�������{��E�i�Fꇹ7�=�]:�`0�J/ �U?c��X�336ՠ�:� ��J<Y�b�!yz�L�����"XlxVHYEB     400     1d0�HW�*;�MA�W5/�>���E�,X�-�UÊ�7Ü����=���tE��\RM��1�%��$�jc%�L�(��"%��UԜY��B���(Ζ�M-�0Q�x��U�r��rZ*�������߅h��/��6ў#� R�y�c?��J������n7�Y��Ú�s����Oq̌��5d��)�ww	J�w�(�$������%�r��9Ú�w[����c 12��Lǋ�F��F�lM��=��,cV&����iI�=���T����n��0g��[`k�i��dyU�q�\.M�+7η̻�pIf��%��[�r��!��$�T(��%����w���	�R��#��� ν���P^�k>�&<$��Q���fk2(��8~�Z(������=�P��:�Y����Q��e7��{=�7��gk'���;+rF����(��~�/��@[��i�Q�:I�'�#XlxVHYEB     400     180�ݮ���ܾԛh9\Ɋ��_��Ua�7��7�<�r�~mM���_���Y�Øl ��H�O��!#��S�w�vE��������ц���]�Ҡah�^jl��+h��.l`�*�FMA�3RG�c�]��o���
��#����#�-��xcZ�E�ޅ�U/HZ t[g�:��;9��w�E@��b�Ib;�rӅPV�ԛ��U>�*��&1�������2��瀾Ж�l��̗�)��짵n�O��'Qjbz&���o,^�v�;�D�
�� ǌo<��2BA�5	����܌�m����(��!�ؑ��&A�#y˫Ƒ��˲��3lb7y0�;U{1&��j�_��w��>��o|m P����� �bxuTXlxVHYEB     400     140H!�����D�\ۻ��H8�D��v��rΐtva2A�f������F�1<�XY_|��"�Q?�;�Bd�M�&��9����c���J��+��&-�[��#&�����Y�p��H�(Jι�!
�m���� P��:��w�Հ�q��Ԟ)c�L�	cNU�ͦA�;šG����Mp�P�����-��o.���v�Pr��l�^t����/h���eW.�M�1>���-�v�݂[ ���r���-�ais���Im���E��r	n��k#�?炮�DI�ԩm��//�ڄ9��"�#�zRf�S�XlxVHYEB     400     110�bqVa}V���?DWN���!(6�]�3��r����FA�;��L�b�7���_L��*��;1L�ڄS{Y^���UI��|w�.�k���UR������KL��?��Ǡ�X��KjΥZ�a����'$�O�I�!�Qg�3F��c��8�X�c?�e.�D����d��m��L���u���;�#�>��H�V�b=G{օ��c�r��Lя]!Gp����Y,��a���u����;� Ҁfn��g�喇�W�vR��8]�h�b�QXlxVHYEB     400     130~9 K]LP�O�\ b�@�Fu-�	πc����N͓�%�.�ׇC��ڳ�gL~��)(�9���Dot��vk*e<Hn&�y�b�6�m���H�J6��D�Cm �F��~#���8��S�'�������	++~]"�K7��(�;��������U��ֵ��G˸�0���aU�uM
�2��N�sa�E+9@u� _�ߥ%{`TF��/~ZJ�髗p$��#�o�~S�=��^v����(�iGl���.�w�-c�S}��r�Bx�W���ƀ˨��k2~c�º�+�ړ�� y|��t�NkXlxVHYEB     400     150��#H��*T���}m�������4��'�AK���'r�eR����~F�?��۩!{3H���x��óhJ(@����R�9�Ho1,�>����;��\q��6px
�)��"%p����7����$ˬ��3Ak2��x@�x��N�n����`k�[�n
(�	֢z=H���z�b|}*-�"�Ë�3�y�7fU���r� �:����R����}�e]+��{Ks����eT�k��/���_eE���m���Ӓ���b�/V��� w�-�7����K&�L�}��efYs�2sAZ�9e�]�N�GPZu�&W˟y�gy`�vXlxVHYEB     400     100�$#���_?�'7{�2�qCpC:���ߌі��,����D� ׈�>�L�_�;<�H���(�˯\pëBg�NgEY��eUS��6�N�7���ٴ��P�D1���B�V4m�r=�!���8Ep+g�O�u�(H:f��Iߟ�&���[#fY�dL )ߪ�ʈV3��7�[���X��g=��N��}��n{A)�L�?����c"۹�oPR�?"!;/v8�I��7m�əi��^L,��XlxVHYEB     400     1c0Й1�+��H�J�L�wd��^��=�6��Qehq|�0'G���x�TN��T����"le�oV�4t�ew7T��<��`83&��X����ڞ��2�`��>���j�=a���d @���-��j�6����Cr���I��������`b
MO�fTEp>1��T���:X��4B��?DHaopqʭ�N�0ej� pP\����A<�Ϲ��c�V�������2���ɱ��N���yCtG���@�gs���=���1@�:b9��t��V��X�Q8
�k���|5&m&� ��d�֮�wP��}�o9N�2Ɔ����	�^�o0�g��7M�b`\+ڑf�����~��K�B�ѕ����*���������ߢD��SԎ�=�I�U��Q���
7����:	�hr��ǳ�I��;.��ޔv&�� !8 ��OX�XlxVHYEB     400     140w}��+����ǚ���=�|R=Cu�^���YNXl>/abəe'"ʵ��*^�R0q�S�;ؤ6���Q�Z�I\��$h��1U����z:��,�(�����~)��FЂ��8��_���Θ\�����s�v}`.Z_o0H�~���^�YK���8zO}�f������j)׉�{���!���'3��С�Q*2$R༞4����o��6G�{u-`y�(�AY�qI�8~�K�"�x���Яj�e���(���l*՗����f���/er��ۋ���S쬄��|����E#Io,���k���J��XlxVHYEB     400     1a0������|� h�i���ےշ���QwH�N�e�"�������.#@�BΧ4Dx�:���Q%np�+G���䳏&�I�;�R���W|�{�VT/$DH��b��%��6�u��3g�,���;�b������l��!���P�����R�:b�G�k	 Y �LL� M��:G
�T}���q�G��$z5�-���4�7#���#�	��9fB����ґ�P]��Z�I�|��K�o���A�x{f�G����BS��S�͋�R	84����..Pp܃�g���]�`&��;m2�v��Y.�?�<I�Ӹ��zZc��xg�Hנ���?�W���-��x���T��~T�_չ0�����仾���(w�$�ݓ:��Q��EA؀_�n�8@���.���t�qC��%վ���U�PXlxVHYEB     400     190Y�<6�-�Rф��Y�4��4t��WR������%��2���N�a�^�")��P��:Z��+�z��6��e��{���m�$�U�[�Lg�i�S:�%랒E�aD�~D!�?2��ʍ�1J����Ŏ��,�hf	�GDܞ<x��~*^; �>�?�W�G�I)]�eI^o *k��\w�21'��\R=���j�hO�
(�"(@�X3	g�3���rs�u�酑�#&E��6.�d��# ���1�5}|Qi���(|&�良�Q�U � �+R�R��hF�GR�Ζ���9����8��)Z�f�Q���p�MA6jԬy�(�Nl��A���g���K�)���_�#�=u�RZ�pJC-D�5!��D�{��� ����w'�OE��XlxVHYEB     400     1f0œ�|�"Uz��t�If���L�24"-��(-�qIri.7n'xF������Rs�_���x\x9v��:=_`4/���ۅ�/�UX5�8Ђ���z����@A8�a	���֎)�6ȥ���݊�G擹�pϣ-��p���%�ܔ�4u��c�M.�����+��솙�Sj[D�b��њ����37n�hoY����T��p�\}��������WC��oΪz����O����3HO��e������5�Y+��Qx-�ĂL�m6��?Q�y�H���q�z�ʷ$V0�fį��R����,F�`
�࿐�D�
��nX���󲦞5��������B��G��k����c��7��崃7���0�؂6�~j��(��K�`o���~՞^���G�J^��|)I�g��r̤ҙ�>�3@���yq���p]I`��ޭU%��s���Ӧ���cG�q����#u);�<T�����"��a���XlxVHYEB     400     170<Y�N��2X��b�b���ׁ�`�=,'����V��+T�4v��5��������]nS;Z��c�Ό]�o7ˀ��g�#K<��m��5��[{�S9=G�Xj��b�	�RaHf����q��A��(���C�&�T�ݝ��5��`�����ѐ��n>�.�H�����G��z��;`@Ĉ[a�(_o��O\�1�ȵMV�7���z��\<���8|Zo.��r�I�� S���օi�5n�TQ��A6ך�i�f6�\s} �+ �ـ/���e���C���ig��/�Éۀ�ə�G�v ����8�('F�P*^��E���$����� �D�a��WE3�s}Ul���3��q��c�GU�fs\�XlxVHYEB     400     190A+�,�4@!����`R$Ңu�ZH�Q��R蘐�C5[�W��������0����o�'�b����W�����p�}0�|�)�7��e����-#����gE\�;��7mY���(u()�m����vX �Z���'��'O��8>2�o��PQCw�@��^@���^��E��7���Ar�<�H(!Ql
t(�$�L���zH���/$�_֛0cH�Q��unT��b����t�&�$tm{|�^��R��佄%m�V�������9��Q1#������ٚ]z��2�c��=��M]t�6��ʛG%���U�_�X�Z����b`Ηa�')E���\!�)=��?���}42���#�?w��D8k$�����O}����"ڣ�r��XlxVHYEB     1fc      d0�@��p�n������{6-���d<�bt3iA�Z�)	���$2��x�9�rG,�k����-��db�:���L@[�x�!+��#f�S��*���J;ީ��v���� �ߚǢ�RJ�̶kΎ��k�?pj��[���#��lӤ�AUyi]mF>t���i��C4����}qH3@���V ��=J�Q��T�l�������$�ext_n�8{t