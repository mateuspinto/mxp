XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��J_�uzD��緝A9@���?"������'Hߐ����6����B�%�Q�x�Y�s�X����� sU�
M"�=p�_I'�y���Q؞Ӏ��(���u�_��_���ݻ�3{'eę��Ќy1Fz�k��L&�kװP���`z�ry@|��uЄL�(��Q�1�If��v׸�tg�����J����3z�߀�g��{�qJ�M���!����v	���6���-�xt�qN��[�L�����U�K3�g�	(?�jٹ,�p�ӕ�x�,�?���Ըbb%�}��	�ONl3���$G��쥹v�kda�b�_�P�O���qL�B��ӗ�'8�<��49��&�b*(��=�2�K4����@�bL��i썀@��si��w���/~����a��MO�}5�]�Rqt )��Q/�ι�'�p�`Ռێ(��c�����R1���-�<y����O���M�"G��;K�|��^;�K�3��>���R�d&T��|�
���冎l]i�2���!a<��H�4�/qWA���T�6���2_UQ�J���	��ԦM��^@��x���,mLn^���W�X��N��B[XӾ�l���A�0����ɚ���j61{C�XkUq>	5��ʖKt`&��C���jM�+��J���P��4��ң0��P�pj�/�)��Ў��!D�PF�������bܩO?|j�m�E��3m�R׍Ù7F����X��Xd%E2�sf�����Bf��XlxVHYEB     400     190*Y+�G��'0�f5�6�Ҍ�*�[`=��?#/�uKa�۫�R��h�-.-�������Z�K��9+��v�L1	�{4UkV������1	o���%���l'3o�=�m�UZ���~WIXAক�`!�0���7?m�夭��L�T��Ars���E6Ȩ�O5��dL�0J�!U:��xe_�W�`ˤ����Ar�xE���K�"�=�+i�`:	tq�^�w�^�*?A�<v��Q�]G�p�ĺ��X��x@�gR�#��g��n��H��5���'��Ooe�Wۄ�6���i?GiG�����B�~�04�����9x�h�0��翗���wRr�Se��ch;�?#�ю��fl�����?��<�w������W!ԵY�eI���׍��!eAK� ��XlxVHYEB     400     180J7NȦ������5���<d��ȶQ�\�"
ϝ�uD��Q��Y��j���6}Y�u�,������`��A99t�~Il&�K��d'UDB�vN=���Y%��L��}�n8��o��cD����3K�S�c=.! bQ�{����n_� �SǐN�E�;YT�������`��ŗ�'��ɐ�Ns��jb��f�$� ��Wk��E׭�<����;v�y��pRIq\�E��mdt��N��Ց�G�(F�W�3�f0C�a��zQ���A�DY��՟&H�s&[+Z������BbfW��úk(�������h��@@��h���$�L����{r�ib�������cK�g?�� ����]�c�@��?j<۬2ߕ0XlxVHYEB     400      b0Ŕ	�X�hN�A����w��w���A��{�vPb��Dy�g� s	u�moUbo�6{������k&b����d\� ��f
J���?I\� �z��4Ls�Z�@�}j�RVa3?���Z7�a��_�W����ڼFa`�eB5��AO
q 4�q�=�ނ
��j�*���< �~XlxVHYEB     400     170�R��5Xzn�۩�� �8��t�E���8�T~���e8̪sSM~�;�$<G ��s�'��B�P�/�0���$X�ϑa���2.q]��wBc�g�6ؤ�+N�},��4�=��!�J�#����))����k�f�̓
��j�l����0b��S7/�
a�u,�Qu����ڪ�O�h���2�����Q^ˏ=}@���ޙ�C�l1?b�{P�)���^�`��0=+��_�_���
���N��6e�A��I?w{P;���P۟��/����	OY�
���i����SK=�߳<� <�B鑽xtB`N��ϧg��Oo^�����"S(�^����-�~ó�G��&�j�G*"�8�XlxVHYEB     400      90)!�Ks6�'��� �<�p���ZҰ���GNw���~9}��ص�$��.��7��I�~+�!�ͅ@�
K۾�u�s���Cy�6��+A�v��b������N�pȔ�꒟T�)�~�vz�[�B�@�I�r4�H����L��dXlxVHYEB     400      90������t���S�sg�0��j���P��woi�M{��P�� �`'m���г���B��<]��4B�^a�"�d�Y��mY��+����'9�fq�������	�x\^��Iխ�9�ˆ�N��M�$8�9��XlxVHYEB     400      90�r�wR�K�J�p��ꯣx���}�+qU��P�]K&Q��P%u�V{� �@u��������|�v�����v� HMQ0����u��K��W��瓛>�)go�YW�����se�gl�N�ˉ:��U�Z�XlxVHYEB     11d      50hn
��B��v�� N�Lp��{U^w���;Xs��Q/|�o��;6v�gݟ��Y�n���h"3!�A»E��IE+���