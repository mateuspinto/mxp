`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25696)
`protect data_block
Brj6F/wuje0CqPGc7I/VPwwQNQ1gCXVsLZyQilassJVJnBtui9S+BLCtvz8mSe1yOr0dsOrlgRJ+
XULgOn+PJfGIFivF+VFwKI14D4tAcQGhThwE8nG9sAl8v7D16g1t/osi/cwWc3KN32K7/+iR0BvT
om2/8LrcQ3O1dS7FpshX72eoQPk5B5RuEqLxfHER8orNfP03of8NKfahkhPWLv2TfuheSJ/pisG1
xb0rMX9xynHPahAUKC/WRoVm7kgsRi7yKm6p7nNKh5rsOO6iEs5eUsp2WbhOXHnb4ddPA9szhMk5
5Wlplkc+btDBBbrhJQx3YuF0dUm69xQ/T52fSoewZR0/N08KTeLWYoSB8oSOSUBm1vFit9StSpIR
iZ+WRitD/CJiYhExaibzy3R5fkO4O8XMSVvEW+MyAv6E4yAxZDV52j4OaGxgyFkBix/oPlucsbTV
lXsuzKAJCHMS/4dSI3F9jXmGrlDMWT7r3trmqLeQgemYxkDOB9+4BNbNWPFCkV9d9BCJmnjL49x5
2HpfBq0lYu2RDqlDO9VzIrZwO/sFyJ97Kw0Iknd8pVdcKgebldzLilOTuxFmfkmz1X3Dbww1Mt+y
B+rfmlzGfi7CcjzYVBYcYju76sXSD0QZae9jpCswTIaq2UcYVe62faXUUzdNk6tQIW1xiftbWVpM
xjlTSdNPT1tvWJZWxJI8GwucEegDWEz3IMpkuPJMFwx43Tcv8mK098LEK4DUhmp7l50nbF9V+MRu
XBAA8e2obL4l8V+1Npx3HmAb7Y58uZtQmM+v3cYFPFKHzNJftekKql2RmdVnFWC9Lvesjsxpykou
Ra/tbrAuMZOdDKU5UK7CAa2QxprpUwe91uEBXBWm3dDPFYxpYahgsTb9evL/3muoS5/XloOsv4Xi
CllfXA70s9LiFWPa3ItE6yHIK2l6NGEPiwmtqmL8k+FxUrQYqSwq5Xw/C70KC/m94wWTr3sJc5sR
+EjlypCZYt/twgBPOrGLTBQIkklX+3+EsqqEWiM5sY2ouwa9cW3/1MavWyIGYaGWK6AB29ds3cJm
t9Q/jS7QvzVKlLxudGnW0r/o7AXuPLFrStU3CVeZD2+dYLImbzbWHCekeYWesH6g5+SfNjgDuPxD
cCViLYSpkaGtmYTM7qbqsbXzDihV8UZPlsuFCZ098ylM9DJ2IE1SgEbMe6Rz1+e7I1iK9GHVSUyq
W22tcGyGbmQjuDUnYCitWKpOivkZMS9YLToAY1RIfuKuj0P3RGux1qXLGQ+Wk2ei5N99bYfKrIoJ
BxtJS11XoMuyPyKaoMlLtSyL383t/w5jdqvKLWc3MgJWvJKYZLvMete+DcpOZmAzIdvRt46hXbgM
PxCQBhkxwL2tBomzU7BP1I6bGBgV8UYubkHMPpQM/BCtwuPFeXgUDH2jIaK2SjtZbRdcNR20ptwb
zGFi/+sCMSLDZNCRf6cxjL2zw4+ht0UWv/sZlZh6xUZ364QH5gWjiEZJ9+axWjOWFYuPhYvbN+ol
YENhhDbzqCIVAb1tdoOe2wt2hLLhzvLVK0cYvkmOTgBiTM5Jy5e6R19+u/I6k8F9xU1MwcM2xCYX
zP7uN55qGPjd16N+qzYBXrB2Tf1gadihEv3Cfov6B1ulOKDKUpuM8g5r1xfB8euPo49sBhIlriZQ
GZ9tQyCvOmwhnK8XSuCV3WJf6O2WKxSlGjabaheyIn6Zo7UGK8cvmIaVDolI5TM9kU3H4nVpKNfv
Y3L6i+SV1e7K1dw+G+1oPV932Vjn6yFlHm/bXEPdys0lX71pobYGPGpxvZPt+Dm72KbudkL+cYtW
HjNCcB+ZVdHnfB79IYrCPvG2Wh8xZLlRkrEUKehSbfiw3mpAmzAszZUoB3M4I6TX8vMTBUvfSIL/
6NzcmnoHrKkuLSK1GAVu8aCZNXjidhrrL0tO0L9s5iCUMx8tgOqMMs02nIwENomAyF+lp6ZW9TUb
joMBJ4CGE/XNR+Q9AklglxY8cyncX4AFe10C6ILFmR594o5eLn3Ak2kC7RO3oXqHUXmH1SuMSZ7m
HQ711lHpAEU/+RFiVddibO72WwnKWyBt6Cj9rxL4sx5RUQR5Tr7QcBP9ZS8tKNg1QJVFlb8h7lnq
UZaJpgPA6EeOw1uNQ4jk/3x76BVxcD0JrFbXDlQmEnlMcRVg7dFVE0VVCy3rQbSSU7MRMrk+UcPG
2aZMly97H0vQeurq3mpJT0saJrBE+eiqkhEzIhYWJNwg9KtqysDE6xnbBl6ugngVR0RE1VmtvxZm
5YJRHeFTHvnyVcqEYdf+4ZmClsXKAp5xDE2lhIZ5L/nlMhJDuHW+qe3I9P7Ttd6EYubYex4nr8Uo
NTwsx4aDda43fwkJ/FAtDv0nufIFSIE90tdx4H9eHRiRr1BChoTmNeidefyUkwe18Inlpc1jG36i
pvkD8LYvASBK5ZfJrjPu9jZvqkLDAr6hj/M8f0yTdRpMf0j4tS7jx1dBUopnIbTFgvRarKpziOtM
xtCNZtp93WPSJFXl9vi/uy03v6OF+w4rsq7xC+Jh6A4+f9JzIByQi3TkWL5X33sEPg81KiAi1nZW
dpeJ+jkDHph2P76XNFUnq8alS0f+rrZZ9IErN5nhDsg5AE5k9hpJ6dgs2WtVDYfERsSlm2ujSF1I
SkN1p6CaxCqDqwitGTLtbWloh+6mt4xBAAIN2QZ20sdot0cD9jRReVRX2cFHnpZl2/Ad0R2Wn6Hz
zyf8WCoJvdcotfiKbmU8W99yiCVwqCArUa5XxmSA+zul50c2oDHaHtZnviolDmrKV8JiUCnGhjF5
2las6cMB9YfJlE1tGY8iNiCeAaJ4d5DHVwkFWrLMjaIVuF5zWO2/tc5kWC/oBYKQ9HV+JgeYlgKz
TixW27epdo7i/NSbW+Re3nl4IZ0uF4pCuPAJ6L8VqCpzK8nNyWJXi0PJ26UxeUu17JSYOY9Hbc9W
PDKEP0cDeuBxZp3CAisBqCU/te2qABnbvF10W6pDRNyt2uVIZAc2i/OAjWAASjAVPxaXKr1+QPzi
axgZAVzJokJUgqSrSqKSlVWePKayrPJI7g8ovlj3UKTXQOtvdTaHLYKe48hMfBlP4F804qm/z5U5
bjZFzMhRjIfPxKKT4x0xunYbpYNKkaV/KTTybeicbGnKQKwu/Qyu3X279ocEfDooNLAnpIYKEzjN
s0kfgeTCD0e34awSLaDKlKqwcTt7EzqrP2KXefuMaoZoJ7WGZjbgxzTptSxHa5GhQDIxXN7j5jhM
Zaii+bVLN0B/Ki7sodUu7PWCJAbd4EMPBg3DyX5zl18fnwtL3YIERBWlYiVDO0e+Cs4QdJMhqTOP
29ZfGGvBQHbls5TEoJIMGOxBdJHtAF6AILzd5cjWObRxlOo5PT55RmmctCm3FAc1A9LWkyurcW2j
wFpFWNmlY7CbI8gu97iFlzWrpEQZqloMDvE01xn35eXIBm0XtnIDQlrcXAHlJqVnuhnb6py5RovX
L28s8q91sDRD1zcURQp7gh94M2wREAR7nap975bW3zo2Afnum2r6+1yMdpkkvGvwfV9Nz3bsyFVV
XSloVzu1dw5L/5Qgos7qMNOqbfQvZ2ZId0ljArNWpe++Pq5xFFu32ww7/g85G9WOZdefVYgK610A
fs4MoC7+pTsvx7BPoz1Z5+ip4Ov9e8vKF8KSOCf7mpROClhsvk4+VAQVN3CHFGM2R5MF0a8lUqrP
p1Y9zEDwI3edjQfaskcIoECwNc3gOMw45GUz1qZdehqdOiJO6H97n2402KeRJ9uvnneoKa3CY/+J
D+3yZu+b6ucQKfCqQ4Q/MOJAYI8ARzdIeE98IyVx9MMeE7C8UhuR6O37yADE8f88gtBHvPRCnSGA
HZ3AzpGbYKOXyThjLCWq6FXwM4DvFcnydH8IRjwJPYBl4qp/+8S2HgTh/lZytejso4hm+K1dotqn
pkeSjUxRaLLsKECIT1BbFhrshLQDbp12AI6fTKAHLeMbybLr6vZIvNV34clzl1JQIPfWdQRFPWSA
HnVIxhfhcqKAzB4U120VDRLymMNNWft0hM2ciq0r0abRcnT7a+b06XW/Ti3Pj9nbyWqOJs+kbz9M
YYT1Knb8CxZQEmx9uxxL9u0mpVl0n8A/TUSp3ue0ertwaLqOfKD2za8G6c8WmzRj8xXdt5yRrjYe
tNJ0dq1J6ZXbX+9cZ8pnzv8IFaqPAxMZcvUlt+uyuQPmK6r85t5UCP6kRTZZy92hJaE5cksVtJ/K
WXWAVva9gm2CfqzgMTOVueor0cQqF3qTMMRNsCRc3tcH2okFVXhAMpZq5g84Mp7sr9je238kXM0G
rdTc2oZRKd9s+Y1lzaiAkJg4hx9yBRyZmBOvvfBc+gKYIj+kQv5Yg4o0Kb1dHk4KJBi5zcuvY6kq
F+YCrhMv2e2+GaJQHORjDxOdWv5enU+Yn+v+2FtwdDD5NQSLGSxa2++1kCn1bja3G32TbJEXy+W/
p2o4knMdPZjiD6SyEJRbJsF9kOdItHHCdX1VRiHCBMvLM/qnsHFuMzL5lWHwmCrapE3h1bsLKTJi
gLS/eEk1D8jBxrz7JF5NFZIfaPMs7P4/Cbdcq0OJe96BGNA6nU8+ERCKqRYUPmB+U1kDlLHR/Y8I
4Msn+bmk2h1B7BdvUVz0gSR9ynKuMYGuV0aph5eI/bi6+LybXv+fQIDrT2zfJKjZRbdx99hnlNzM
lMvuW5zAjNZsGNSf3juRf0vYB3wXvsTHDTk//L5BBlcnLzlKu82CoCAyfuZbJJiMtnPucDXHQJqy
szpDmM+a5wnl8I9zN5T6Gr7clUY+0DolBd+qXEHYMNg/jLRYAb8RKQGgTV7FLygq3MLmDKvePz5F
glN0LtGWgdOoxxH0mVMi6sUwyewL+MqnQY/J6V7Z89M0OVJw2otQesUhHd0tYrJWjqpBF8txp4i0
lk9ILt4lSPK10m051k159Gaek7w04rcB6GAtsv7orHxAaFRfycCeYzY4PZn72ymIYyBbwZ38h41M
OCb4rfsxidZMmXlBrC/RHyIAdvsXNcCfiDGaktubiSCGNqmnHHjUbA6ThZuzeyPsnHvoqRPV+tpo
h4CbDHPb9FU37edw3AyKUryasyYSTbBbxiq1jd8Lq7KM//IpOtukA/n+eb1vfWsp8M7dE5WwRVEu
URlSiBWkDfNHe8cXaCEZ48Q7reFnmd8MTR7Onh6B3cbxiFI8dv1hsJuhqX+gn6rzsuqPZOY4KLCp
njjaFb5Y9LgT33NTbC+u9mZr510p8aBP6ZMKmN/0qTeauZDwtxVouDbvwwVwtKGelm8nY3o8r6iy
DCkb+kwIVRUhNbnMgDc0L5B8SX/IGP7tgG39+51SthNTiwc68KXRYwU15DizinR3ZPAxNWTRDvxu
y37Z0ACk9iOwEvwv1kBkPeHjSBsLl37wyhFY8oJIY2sW+V2Puc54fMJf6ywnr+cixDC8Zi8OjF/P
H8dFGfLJVwn9rK/MFqgYZ0j4AcyUVCSib1bkOhSkrvwCvvZllT3tYBo78k+4rcFlW+0XpO7HGPY8
1xmdvdejqrgH1G0JzxCyCHPqOodXJx5JJNrvc7jGaUZoZf6AX/EE2pSxQ6+UhgAq70t7shcL1Txm
qdZUWd18k+lvX2OoP2lzNL2Dz0/DCL1YSEfiOxD+GWJx35tnShWwJN4YDGY2lpIOeM9oT3YsfIkJ
UNQ7lrgv64DvF9yy0x3Gsh7j2bvntQBY/4ofyhnjSQ7Fsnz0Zqks9EL0CvKTP3y6Bc8vUcTu83vZ
JfBtMW+Rr7UwskGbkiDxFZbczJD6BTFEV42knHl/fACv6W0ux6bZ4SuHo72juxbMWUzhL+O143gr
TJYGcKl0E5cdYwR00KoAHID3Jzf/5xFs+tGeshjaYvOLgcLTgh3N+AZNQuAhu11QUP+KmCJWbaKz
v6mK457WuWLBm/UFXZzPBWPTlhUnV8UbeEh0jysojw879guBB4zKUXZJX6aKlGGOcUEJYqlHM17p
9X8D9LVSrQlZvYIrYI8A52+yIG1C078koDHKtRHLcjmmJSnUYFymrAkRnWDJ+/j1Vawe2n20N69+
TyWIIqd7M3ut7CFn8lPhi4aH4sWpiiSpd72O6NSYTKEEd/XIIMFkKAj6ZVp8AL5yex2MUqPVYOcj
RVoQ869MY5Uhi2XI1sS98HTpkAjZ8AGhdAqj3Orcq8rKcOKSyRREJ4y0ujjtM4EHjh6uOsUZ6T/N
t43XEaVdqUMnGHWDnmSJRfEeXyDLc1VOiPULqUZIbVJ2KcgSLAeXtHw+wCDtbw0RGNizXmJ02TzQ
+flkn2oIVkMf8XEwT+N0+TfzVvaQddbRMnZVw3C+frs6DOHVmqBpqjl8+0JzlxRqaHsxSBlm+fzD
MpKT+UTg/j0VmoEmcAA97yXXgJtgK2DLwd2vn0+cg4hq/QWfOKlNTKSNUUFc0TjniTOWB2GRAdzY
5ndsua/tQp88Lln8rTF2qJ8MlrLuDbq0ec2/SzO2vNJZz1ovA1gPaP2OgfJMiLyYMxl41Acx9K+b
TnG6iF5eiAcKelGc2O5/VJAWRbx9NThVbXSMEvONjtluuRVCTXu6WgRSIEkOwnqLR7FucaLkDX9n
laRseya70VPUlXOnsUS2YEiwmjONGoNknff/JbBwyeGTYbWXkSL6Aq4WQCeobmJVQlKu0MV6vLgF
s+uouBffQkRzBpTf1R9K3kMKnN/3MgnNI2F3NpieLtApPS87rC0fK++sw+xITeNTF3PPPjSgffKH
lJQ1Zr3/omoSNywvA8PvAlx2AghidYWY8wzIAhrT5xzsuPqevwUeB+7DHwCA0WLstnVAgZU8s6iq
FJuNDYuPp367QhpmUcql3gZjA58GTwqExmijcMMUNwz/GhBanSgH4twY/I0lcY9msH2sH2WJ9IKL
FoH/ksITsneVQva26pjj+6xvmTuGLqQnnWQgyPiCx8PpcIs25BrMIWgUjX5BzhdC74Ig5ViBTsmj
p2h1CjrrlxPY9zPa9dFboX2LKIrPBvKINWem5NjYARWHn4jNRFylLaIw1w2oyE44k/FVcWgWLHaz
afcLaVoXyevlrTC7TznyL9apfSKTVJ9u6tHEdQkQke+PF4MP6Wn73bPDEtKQb4Q1Cs60IL1bGQiu
iNZr/vGAw+qDEG3Z3ifYI0rgSOWgKJKgtYCeraKzes9qSukpdavhdln0Vvtvi8LbVQxi40Bbtg/O
xOy6w3dQUeSj0dQLm9xCvRD8Qsh57BCbUy+3RceW/rnzmJb5wHKCWraP9JqiyNzi9LY/fSVcPoZG
aNk3sNQz+NKwtuy0upKfwRVZ9R2NFw/N0bZVQdIruATbcwiEyAIYXuC9c3hVXeiJH71J+Txt328Z
MMMU3XoY2voYQ8Gzt8J7KWfXZd/KE9cV1I3vmILU7aGEcJilfvCmZuoAK8YaxrXTCCyfN3ETej2l
EvmGTYPJCgrbQIAYFzZsfAM2IyGTjwBIuwO1p5Y+l7U0oQ5mEpvLOtH2R0sibUzq4hmV7eTEGyps
FUEY/3IsAjqnAiy8xu73Kw7/rUgzzj4kUCAVZ9XlQRfmUudb4GfYANEWbgKSRCMTEh1RxZoBgHnL
6Bd5eYCQTtYMtvaFbuyLMl22WkutIT1xy4mDLdaw7Sf5beI2HNeCSVsFIwKcnd/7P3Z6y37aGlqc
157DC84jEBzDjf6jhM5ZRyJZYV3Kfa+VmkGlCK7ZVv5ckQUmjIO7UbtuwpWQTUcMzi+PCNvNOuPi
QbHBv5X3/Z2Qfa9vRHFrDHx8xWzRDkzKKEeegMfVNulys3ddhaHVrGpbqPRrtRU6qMgcMv970x8q
N/ZKXlIwyLo2U1U+f5BLSkVHw1l6hw1tGaSRHa2gAwQ1abnnhikAewQr/TMjSXodwHDFHzxWgqr9
WhuMXDIrR5Qkmwe9OrE0kMBZ3J7HkCh6cjWxPjsQIie5mkwv72DRbK4ytbMRG1grNtB/ux5qX5Yp
cbD5n25D69VFrZGNgzQMYFFrI9yK8AAIajWxD3+2XkaWWxlaJHjn4OtqOdUqDNpG15g8h4RDSr/T
q5olaltR4EB0w7Y09VzKIYtSqg+XfemwvDEhLSPbVCF2GdFbaPxpgkr1XrOqBfgbpagLwigq8/cy
SaiBvvr5G2Ob03LcuvleVjVCuzQ1CW+Pw2pFbq1VZCqRfK3lXRbupYRg3fpThkDUw6aNB8JbtPXl
iphs9HV3EP07jH/gz/1/6RpSRU6D4/YHLBJjHkGv//ReYPhsFGCUchLav7pKv5XUj1iNtXI/sVWn
vr5SpCd/pCXstm5eitgUNgmTFD0HLI46oPo+2QgQSFAs7KbsIE2cdAFt/eWA/U6mscTXpAqjoK/k
IbEEFmncIdShCenarEoAiRgIAyhy/YAXtD9EuCjUtE9QyTueHygA0Z7J85p7tXAmNRM6aEb6uPt2
GYWa/bVKreAzVRH+aLlgC7gkL3Hj78TWmi5eN0EwBQfyiLVJ0GFBuUGFjFMUo8wx+sHPML7TGXaw
m7M2mb+kso9RZSbdVuNhFCpMkGcPLz4niCYZJu+v0nWgGMc/0jXSzC41OTuIt3jMrAzsZ4lycwA0
a+aMBZWOJyQbbdCQoQ/S5SQ7K5LqbGqnuXAAwGtG6zq5Z5Rj+QxibVHaRRQmMhn9Tr1Z753nw8v9
wSLDRfMktyBoVEdSGanZtQg7RHPyQEh1xbWvp3W7gO9noeqHejAtLIizNuEXF304skpN0DhIayI5
LTucP/hz+HyiWoDtMs1aHzZPu8jAgZvHZTNZJb9fhdlI6zOyLp0HYS6lvqh88HgXQN+nCRXWA6U/
ZRPnHzL+sw0x73nN98Havz1746QAF0wY3luUgXQ43KW1zhR+vYF2yg0bJSV1y2aYCh5NU99zE0uR
N6caAqHxKhbG84YMeJO94SOgoRTyacpyiFD8fl+aVYCDbT5hpQilnqwgcTIWdc9XFyrXAKWEldE/
wwIidMK1Wcouvhqd48IMbr+M50Yt+f36mkUdPcw5XPYnghX/+Yli2MQQ77u/ZhAt7xZ4pofdw0C4
grH2y2IhO4EppMPe8u19XdyLQnXMwONebPMW6dIB2Eo4jwGtszDBuG9SYi8MjxtU1464lVOVq7Om
9pajHi7nM24TJBO0d/frC4d85+ljXlW5kejt1lGTV7ffclHmsKNvpsrCKGUQycXQg6kXuAu4x5CK
n7vAJFrgRHymEnZef7pX6DupNF204GXEnste8wLrdQSLFv1xla/xSTTwFKFhDNhsV5zeS9EKaLi/
UJ27VIpY9saQjd83JRETARwyZym1w5BWMDj9SYxB6EV2kqOvIH/7h9cUari3EELSXkUoOPtzKRoE
6h3eKzTUTDnuthiPUeN5yXf5pHxJcZgB6F5d54iIWosSYcua70//gydD1TmeVaGAGvO/qkDMsULd
KRCUVQhEbS025L/TYyD5oLO3KYV5Mm4xvQfS1efPY1prunFz4Qt6d1nVuXEDNFMzH+0X+DG3lfec
OrhKh0JP1oK8D5yo9Lv+DWsrXhIgzuO+WACmnrD0HdgWpE1OCP0g6jsHerioKxhKgIa6/x95aEqi
RnJ04ereUcdF0rpnxhGMOQ2b231vjNBGHYj9oq9VObs8t7DHVldOfDiF+M73iY7xFqzMPcDOI2zz
B5cZWlBMzO0Qbn0gECosNcUpNMpNFwHWZhyESfUlF3Mt901B0U4PPxjW4pwbDHOwgf6+wRSBGTkU
EwBQBLn2C8uIYkPi2bdtLpLisTb5vJ+nXvMZKkohJTKKTs2gEXAKW+WN8zE8oqtbUdKScgRDY9X+
lf5PyVobxp0w86vorMeXtweXuAYcJxExB0CYaMXIC2ZrqctzQdjQ73/jr2RNxm1iAEqYdSc5FZK+
DplrFwIwFSvOWGh12EFy+8CxSZxxwaXGIjz1MES+LvDCE9kztTr/Jqi4YOHPhqTxEeYT6NGGtZeA
Eeb+4OzxVyFWmvhRyVO8/+i0qvVl3kP2cJERceu7lAc62BuSkVP2f+upiPYqAM7DeePeEGuCNAyW
7vGKvy0Lxh+VKXEaXYaAW079rMXb8lHYT4LAl7z5LYdgjHay/IRmUZySA1lt/9NDGpD4WjajLISU
xrFvRBY/D4C4yLRkdlf8SI7PwSgtcCM7yhHMyphhl/Ldh+deo7AYjLrY68B3mojbUgFres9qGSdZ
9kqotQiRa7ZVPN66yK/40gD0no2qm9KyvJ4FWqEA0e5oZxoGKn3pHisDSOqAHOtsPmyRJCgZL1Wq
4rCMtrviiq776wBlSiOk5YxZaCOfUwNMBwhRcLRBgyS2lPI94n3WyKBJAy5rDySHjolTwIXkOX8M
wN6+2nFq4gWZsE4bb0f5uSEngW3uXZhYdS+OfSn1KAT6YfVs2Xry9CY8HeN3jJhWuvW8hJi4eVe3
AudKcssIZ4dQeoNoNtLoT9cZcQ+ZsyIJJ07YsUvaBtk2G+9mUqQZHzq3T4NvnML1WvBUOfwZ0cAI
6lTTGuPipD8Q8zgO9uQzHvchL9oQHY0OqdPP4A6F92qKGYWQpqHDgiChblCkCcuOW1TEOVDJGKyz
VL3RH5XeicjAMQ4yhKoQJ9/u5VBOLWDFW74MFaCvv+YWe4XDVYV8vV0nWi3Lk8tV0M0rvMkkWNRY
jcGqfDyFWrvvGO7AZ+cPjTMuPCnfk31zVNayWABL1ahCeaPbeFABEb4rgUrS6f8anF17Dx9VYQD+
S3b8Sys/DbM+hnKWz2ZZ1K+4xhrGLjwwgvIrg6DfalojLQ4oHOOpC2JBUd4TSIwO2blZpE/Oyu++
Tck2BgvHNrYP/BGruz7Cv+MJVqUJRaC+qDaNfStB6erGaByzEZtSsc+4VOmPKbQXKuEFif8IMErI
sly2Pk+TxQP78hDYw0W+kO+dQOkVY+RriCLmsa02oo1g9aW1FnpOzZtlcA3uarPcy0NpUYIATFJ9
TJMbdYHmxNtcLxld6Hm1D8U6zXfjngnsJqDLrfdBQQ0G0TmFraVZFnV57aG8rD0bErKXE9qRnd8B
h+r1VzOKtNzLK10ypS1U6HOt0zq8xPIow+tvQc0pKL+nL6wZkRozlM6BQ8W+hb9bYTcTlIsIyQ+o
9iopq/MQ/8IahrmezjGvLEebJJ+/QJ6+470GzxkP86NNWWDwMmwmq0ePHeRvx/naucPIDM6LB1Se
RP0VyVB2uUyhIF1tQd3++YM7ZDf2Qj3FuErJWcy7itL5koNSaflp6m6UHwmILR6wmsd9NWfryxee
qgRlcFa4FHInX/S16yspBQmQzm4DdA4Lc/U/mT739/kNy311t0TdvpVDCSlLkW0TQTZNm77QIPWq
j99hPJBkcxqmJ8TkFnseuPkWxymLEyRGcE6UI01I5nVoA0GyybaIYNdD1jCgEeGbCQJCS+BVjGGD
OgKl5FuqqMmpC0KVmUDYBSShY52lbGF4p9GT8YtoXfOThGZheXWfn0KYKDnL5jpEU7SZweieZVYm
Z0q4uxRkj5kVjBQd673FuE3sdL+qLgIQxLb/u5u3n9Bw2Ymh9cGExfOcbOeeqmQ8p1oD3thcQWLT
dDUTeDK1+Pf/QXc9qkLbuufpl7fJOuOGLF3TSC1GVOQEUOc0zyvgQeLIwsE59NOtfTABAQhFXb4W
5w1nOzslXJk1xkWCQ3Vs4GnU9Hv4QtRNopI3VRiZPSVyA4F2717Lung7X2d0jO/Fgl/JjcARJ60J
/fH4qnEP0sCq5Va0awj2iEhu0/YO6hEM3KkRJBdWOEhT6mG7SzXKgNIg+zhQkBfmBsZiZbkVK9cv
d/ZkHWMPmcpQ42sjLo0oPG/hFYvwkS0OsUDINBiP/Js1mMo1dCyGtO4NTS6eVCZasfPgvIHzrWJf
3FFEebbQJbkR/GvT9n3mG0fyU9uZ4ZHGgPS8w5IaVxJp7o+z3vAeEKOETG1EHeGqM5CEzL7FWZ8G
34SjZ6ZGAeBqwoAvX8WD9abmvD/r5++Ceb3ZGg4alCYMPVaqhQzn7s6qgSed0Twrd5oHicmStvso
innbgaUapTf9MP7UWpkgItRQxYY0ALHF/jyEaR3f7Y+HcyG59RM49Xyf2cuBHKUW78sYVr228T5L
+p5QfQI3uQvi7UIZqOaSbeoRtZPvSEoJSyp3Ur0ZOSkCrMAIPpQkfkaOBeDL80rsaxxwAX16KTpD
WIWZBnuVNHzbMYVB5zFvl3JORNmgBIRo3589Roqrc/dhZHPmglp7VdarWGG+DECHJO4xXS0U/ies
Y4A9uZLTZaBMaz4PKhcuf5QT5x5jVhnohS6Trd9FF/P6Pth7xUJBbAymk/wXacGiCfxnzeeCZkCG
XziBAPpowmPcoYkzQ7hr3262ddO8qTG0kS+SzyuFQxo8GJMIFBbttqpgE9ytfaO8h8uL3srzHUQK
u60gv2pMILHZ5X8y3gvEbtv8PDvQ6JmAmlFFkjofK3xP7x9IjRCBeN7k04KpECqylfsImS/MBj1C
QXNBfVAPqPlkFAtSj7ZNm3KSbQekFqhgR5sNPJOSlMbUtN+lWRZ4x8JjwF+IKF/sEt+Tx9VyegmX
wKcah2yP9j5+92QIT13uMz39H4poRKH6Rs7ecPWnzPisR35dRcwvXJPgXzzc8pkyAMQJdSGfHr4e
bR/+gkTDBYhRkjwngAwjpJio0V5RCc0vOXBFay6pCWsvlCi0T2o4oLwNF9NYDAfAwO2b1w9XWzGt
WX2fJZkT+PjHMWDshN+4RIGQSrXM/ZQNqYTkaH9qlospYzShuXDAQwRb0St5nq15FiAEaLvHlNf4
6t1YFGK6Fqh7CbsDgOAb7+Tb4eBzM+EVMNPXgiuOkVmGsvjKJLwQ6L5T6g1lq1Lms9kKzpwtaFec
hHJpciDOAq86OtqjzwKm0eE0W/P5jVE9xlJBoFj4PQRBNL98zUqkB8efvtlqkfbE3QMjIDW7OTtT
iIqnyV3Oqov2R2Xj6eG4FOk7v7rWFaAiAMwmGo9sRFnGQVu9dVCKPcYy1YjegRMbXE3O2T1aAowR
7veOcETPxIF9kgNhBDRI3OHqzqZfi4zAzRH6YRsG2uVBzpTccZG6Bemp3eMqiEXUXnywSdeIfJrl
zHN+HByEU2UI8M3+MPFe74wxSzmjE3t0cBSCEdMJzIdYTnc5Z+Kv9/V2AHnNTKAZ9EaDBKEf74HM
UUjNCgJ7emlm5wMzcWu34aFI8TkbR7F863WMMZwn3VcO+U04346gG5U8S/VFfixcWmMcmCaWad7I
Ma8O6Yl0vJm6sEmaVhEsy/dapVL1xvic0WQoNIZfTT3ELFb2M/tr8i7cisKfD9vTB1rxqbS2hBHP
sZuk94xgOiSq6lJ5SvHcxObQT3hDt9x7e47nZuLs9wsTdIgeFlI6QPeVeVKdmwwPCexC1fcz6RfG
oYOc2YMvaoEp01KX2Z11ABlnXQxLqlBiIj4roYNXeyUjs+rgAtuid+iIsYo3plJoPrjg+RGnSJSX
S9WpXJNPMAJVxPH/7W6AVZbgVuDHb4GY5ZtTAKDoFrD6v0id6CFMUwxRa640Qf2FfGdEyxhEYcSe
m6m0jU4XJ3Mfb0GV7k/fw9F1qnMGNVIxIjsXsNcUa1GT7dOu02NuYrEBNjZgOtyoWzi7guaP69W1
U8xA2x+jFnwiWDH7AwelndnwWfMrSvFa9sYmVMzP5Xkx1K7b6bBXNKRCg/e8C9kqlziG7WwmGmSV
eMM7SvPws3fHwbCPD17hOOYdDDbRCQyih11uvj3G7CKnhhVJuKzj5W0PxthO69Z9gadyKqGkcImu
6eNekG+3CmIEIsoC7w/7w0yy46Na3FzjoklWMRQRXtr+zxc2BkdL5KAHQt6a22JfIn6BNoHEOedO
EX47pQx71uW+s5T/4ucrqS6LBZUywtTAPO9MTP9MO5RXof9irDrRGwetPhg/m2mdYKBwgizt7ZEH
SrwzLhni0imbMRA5z0oBVgBZdAVkjWNw8BoTWCUkJhvgOB4z40rFBFGMcoo8+niRdUm21lJcy85f
E3TdFUFAU+3t7py0S9rIDbaX35g7nD46Peq7w/7cVo6l4A+fuVADMGrwgmGmN4xw7tXbULdO/u+u
h1kKivLZM4bq6hnDERdIj7lR16BNoJHpMDc5Qw5E9y1oWCku0ZW3UxBm+rFaSb21aNHpLon0mQMk
QFeSrnTBVyRXV44CGpmq5tLakiipRtqbWutsVqOyhsuKlXc+vHO5Y7JP3tQ/h1tEcekGHtorKRUa
fAtDkbG0QTGRFbEju9vB+8DCg5UQMGsqNSQUR4fXLyURapmYrSxnEiZrXWKO26sufFj5n5CsjyC0
JGcsqQsvLOLQ9NJgo2Etf4Qk/UIB7D7Ku/tX/YtpSvBiigUNChSKgLk1XP7XxKnAlD7ntejqoL9d
YQVj6xn55HvTKHETm7xeKYtABiQRLUyteqvhXgHWt3gEhxzyvjZMS9BVXKBejXRLYmZ6dZrTdNxk
mC6jhQLXmWPLVLSn+uIKWLCyy8C15Sqr4B3CcPcDHgmFzpEuYelSEFQ7o7mEcCBEGoZoKbmX/Yiz
j7bPFAnX1INtBsHLYdXjPVFWaZJMlVmW/hLLxRn6lidyMv3A7MXGYmLCgVxSUmqVnRFTtA932O93
JckMA2c1EIOv/cCrQk5MQcYUm06u90/0KCt+U7p6Ycq2vkAmLqNsQxR/GH6rutZvWUOEU9vV14Gd
STYk97F5LwqtqjLSBRGCZtQYCu3Ns1wI/HaubqtOZWkMLLm/wPZ1lk77wgrRKT8boDUHtCsLQe05
vid2n+j/IYQ4tiqo5bNssdRfjHtvu/yb+++XfCzi7TSLdigo9B+RznpXQjStkJPxmEpPJuMMNVr8
SuSEnlUIF+jSxoLsyH73sYl6xCFvw6Ik7kCqjWMZim1UA3LWODX6JuwPMocQYaWVWVXIZOpkg8pS
mgTIHmlA4YIZq2I00btwxp8LL/kvK9+tr7n0I/kFsrICtsI2KUDRIpjiPKWFFHb/ImvTx3+6+cG5
Bc9CIfTVu2iW1co0Rh/wwkj1v8iM97/3S6JJ6VVh2IwUadP+OWPXeQGXakoTSSHz/aP5p4e3BlcM
v2YdkqsRceQ6b8QPL8sPK/uBIQLdjj2giV0nAVftOSZQcPosT1Y/h+nckcP2mcueLqbeEZDaYEA2
gYneHpHX4pp0lEhYagwy2CohAttrnu0CMlo0XcXDwHowUIWAFTCj1sbU0+VsbSw90o8aGSeXaDeg
srbNzBJ5GTnWRcH2cn5fETj4NfP+OWIh+wez9yU3goayxi05MXwW+GUZZaat8EKVAEjwQK8cH3a6
wrsD/L4xcpKn6F13v0alrkxAS0uNczsulczpHZC0Rnaw9reXeRpBHsXNwPcQ/8xxbTMyWF7Fbh+G
4T9VIiaeL/EGUzEu/GNGPDTXHKLtyISTlyPbt6HDISy1m7hiOPUHgN6rL0DDxVp/tJaorSBiC/CN
K4R6QcK3JydCtFkUAUDMxO7IUiUkByPFFcX90p6CLRi56MbkOEbl7v6surp8rRTCZrnhX9jGsHqf
JYpmM1il21oqRAYQ0iqc4phJ4yN1Hy5AFuIDSGIfg8ClY0tu+EeQaCKS9Jb5MzWbzX7zNpjwP96y
bKNrLMrTiwUAFMPb9QpFh/Ibv2yVTgvL3imdsZ9o5K5VYHzGWJRWhjsiO1o+O9HOxsIAz8H0Qn89
GikU7pUppYL0w3P3i+r2GMx+PasrrvyU7/GNK89dD4qMqpvoOwBjwND+ckUiv9bRnLLtreQgBB22
J49Fh9+CxcAyJ9pF6ctCZv3KJydqn59cYBqrKLaEuVLECKwXc3GhRzgofq7ZMQVG7c2UZ20AA8LJ
6n6RYgO8noZ88iTjQeCIMdJ+n0juiWNfh6Nu32FmnT1xUPJrhEtOjDC3tGUMWqYEAvsJ11otBQEi
Tybip01vOa44MDBWm/X7W+VCRHyxcDKcLVCkyeuNin0xpptmTPfuno8cXHbWSCcIBiuDOs4IyWbj
082yB8qbkl49XAT0g5ej7HgmNNhnZ1ZXPDOas9mvjiZFgRqSTvsutv0PK6WCQ4uY0DQLqDC9gAkD
9Og3XKzITP413mR+gJLDj60hg7xSl8zz6EfReuJnZJ3iFjIK2U+CeyukFTCeHzQQGT+uTqiYvP12
vu+phh2RWAoFLKgYrNF1qgN6QCXU9zL4GA3oNol5GbHvnVLL3UzAcxSfdHZXVcrJ8TQNmC0TiIgM
jfEfMFYzOJPpGy6lzja1A2YR2lbYAkYKDHiI7AgRahhBEn6C5eS+sSU55ZzfyiXlEwq3MeeMH+XU
VjfZXAxspPxooNmGh23ZxrxzDwvPOHJ6jzy3s3NFdR3MEeKBS235Vvn/Mob9/FPtJ5zlK/sjwdyx
DehFfPOx27H4HIPCr9tNrznYIPbJo9/z5yut70dGHs6qAomJpkE+gk4RGqudavr47WQVhXL1euiO
8SPZ5e6V3axvhuWhuWB63kZ1tGGPDaaMZ3DM1Wy5IPtpYEk/PReCR93EatQIn6LvQRis3yR/crbp
LJReE2O5RnT6ByOwhrEQ9hxfNCe0jLZXPNtfIawC4zcrPeuRieLPWPsOBzbooYAq/cQm9ct/+oy1
TcDIjtbMlK5C2QF9bHM9TdOkjaGxolsViKleqvkIYEpOsA8IYxX+TeXaRf9ZzQo3Y4YtO8jIgA+5
wZIxZI0EG6zXik1XpaJLNCpYGuF7mKl/3e8pBde5lDwGSjQZjOseAx/HW/pk3Ze7g3mCr7z2x0Ag
euradmxI4jtTHQD5VjALhSknhkgwhyAx6bX4ttgO3a7/vRVBHkszO0IO8KowgDIC0WDFJ1fL08i7
sPVt9woLSkowDQvAwdjIPjMCcSUujoKJw4L7Ut4U/ux71ZqfE4QxqWjp2/hBqJ4MDQitDmU/FAJB
Q5TBfW3yGSdZUkfpZJUasCtW2De68E5xHIBr+q2N8f2vX0QWDyVWs1HCbNIVVH0mMPR6AcyCp5ZZ
amQlcC1j36noTMU1SKs5RFXtdhflTP/QGvNCrT2bm/WnsYQMgysSZ7oaEykHsX+oieiF8LPS9M4M
jEG2N06xXDZjE4ur63pBqZqTgnjRoTbykBn2HSWwcrnZnhD8Fy45eVpnhY6nC+4OkqE4ha86TP0+
+/0KLFUutSTiW6QRcgv2rkc7c+nk+MSQcpfqf+AOF4NAaEv3UjQstVEQdbYZR4SS3u0bArYQh62B
AqRvfS3HY4+AZ/rxiaTUXHaPA6SgO1FJRYoorRq4hlszQ3csqFUzNq+nVS2Sb4BqWmU5qQinwe76
5XjJHqm6ymYnlVBOkEw9lasxW843RNkPVU6xyp5ec27MvthN3dVCZI5ThXF8KB72BmlQ/OElFxUT
xDs+uRjLvlMTeyGPtLCaAmO38b9AZHAeHxwSnGteBOiYYwFCMTy2SzE8kd2L/sLhNi3VnxV0wApk
/H2dwZGukCZ62Bv5GzAnZXDOrddtsE9015G8cmnPETkwLksExrUxvE3XmvP3uJXY3SG6FNxbcW4v
rMWT6ocKgmWugGQWA4pFMGgmQVODsjWvqMhQ1d+jpnwQr7u6hiLrJwu93cJJBAPG4SflzCaPrbX8
HyC19QVfxjMdvzXztiNXG7Nee5HiaONPQDLHir/EmiXXCKxScwMieu6MprlycBxEEW+mCE4tjG/2
Ivcn0BFMYCgu9rDNVQwBb3b9fV6KiNYLpPXCzvvZiJpXSriFLWVBMo6TqCPGw68IxSxOFO170OJe
AqYBRPL5t29sDdqvt0Op3I+inkN8j+E7dca1jnl8dF3+8tkb1pmuNzP8hT/zCbJMWT6dO1qzWiY5
ind1OvoPR5GAoGb/kX3Hc1nysVV6PmJZzMc0Lu269HHuDZCD969Iy/YGpSbi3OrKNuhPbdTqfhes
22bKJxhBF9KjRY+UHHfI0faACdmq2cYtBHH8WUG0ychjYxQRIeSMJPr0+JR3hOcSeM/c4q8suC6S
5yNFq6J+q+GsYuz4NUoqTwhDc338NFfLi1ofWMfUamOoOfiPekjWq2P06CxaAmsYUi6BPvDAZs9c
T8jz5pC+ipDDJTO3sCPva4YtV7THrHIxU8yEcItXncUzLbrg1xsqR0HDDwtlkJFYO9muS+3xiY3D
KhXNBm5sC/pBNb2kS5o+ezxeHyme8qPLfO7EPiH8h9FmTj1AqNAO25bg2VJkAQz2UgqM/PcdyvNH
zuRIRhBLw3VEm96XmlCGmKWuBj0lRvNqJ4Hy5yDrv/md2bDZpUzoxiCLZcFU0RVBKIKpRepdITFM
py3p4huDyMr5mfxgfqLfk1w4Oc/67sxz0+w15BohDDplTN4nCyKpGPs2VVSNvcqIGlLOyRJpBZff
Ny+2RH1RtFO4X7N+9aUO8PlAGRSr490AXsz18b0IuTFe9Qr7JVaCfADhONE1IxsfQRz8eyCHsvc2
bwEvN712ICrJgnCtAVE6g0ZiqQCGEX2s3WmD19AhRhnPZSYDuInNeFM6Icnty1ZEKiUSV2O+SFCk
9oBZCVjGQu7Y/gWfEUg1OSyyfCuueti40sOO29RBVuWrecFC+k3fLOllNrQbKJ7GeU23sQorlFmt
vjTeuoMZk6ltXzcTUQ+iIrKOeeidEAE1nWvToTdPWz2gWJNFDq3WEwsF9rk7wHAVvzf4C4oVVl2R
F+P5Kd9LWkQlHT3Nt1//i/Ib3o5MYDbQAmNk0hCCfINgm3kmPnX01vze5Usy9cnbWDHHwwPTd7qC
NH6+x/qvJwg4Dha8WPEoIo9hRcXVGNamRp2Nw/GxO/jRraHCEoovh//9ytbxJoC5d570yF48TLz9
ELqgd1MCUVLFucwCbrOXbJIXYQCuI2YmrAckc3S11BDxWKUukQW+w4/rwXHsGEis5Pa0INCirUdO
NpvTNIp8MIX3trmSwBEq1hhBLzDzzalgtqXx2zM6Lo6njeE3EqzXjACI+hMQFwdszqqESgSRaovK
oFhWVwnmtsE99+XWnOqGuMNjYrCLFg9BRVVaFrnslKQVMIXTXhvNKa4A23wigkuTCqXeJtG/Rg//
R1NJSQyos1X0mZVqNcGc+iHKerADIXYhhUwjknUiuAcfNGcCB0l+vYphLP23gArpv5zeg0JihpSo
KmCEOwbk9vGyFn8dQAhpXz6JvJt4jwH8iWxKfGmgRqhb/Og7pmOMGR34fVKo1c5pWeF4F7zIAV5k
McenW6PZdyN9i2jOfMxF+ZfTSK80Mob0o3UPDrS7ednhm2kW19vEQWPjbxLwHc82stLJyEnSB/P5
Gch/nQnNy5kLc8jcGeDgEDZdg3JNr3tcqXF9bP2s6gle+c/iZ0BXW0twcBR6Itr5d0O/WhDL18XJ
JJcB3OdFZs4Cag13KYNA6EBBi0qEnhl3i4EXbri4RoDbnpWrKm54e8KAJC1pHnO0w+DJkliAzz5Z
bqS34obiQuoIYZba49NwInWFlq7L8IRTwr1JlBegyK3Ve9HOL1fa3GV9kikr2yHIPwEKa7GZAWDz
63BV4jQRDC02lDMNKxbNvTQ1d1v9O3IF7BxIsXG4Sq2GcFG3CfKDS5Ozn6Xlqz5NNSieJfM2sZdC
tACo1osZeiONyEllqUZ33FtyqaBR0gt9OutC4NsEIyd1wwuyhBTzWroz9FUoSZuRa5nWC3qSdWZH
YIcz0zBHzw/XaCen00Ap+2CI8BnN96SRfv1bion1kvaO69KJNwDAN2Agq36IjugyVNuDzbk84H34
vOlfpws66cx7hQ59qHoS6muFX8GPi5ZkXKeLk99zDd1H5NZcS3ufnj8hNqhRvrMT/TFIIVdkSn8E
TboFaxsunFsgKZo4oZO050Ri0GgB004IoJb0SfltfJFgvrcttKvWQY7AEzZqNPr4CW3zaes0qlmD
cETl/qJ0uz/kZU/81DAgKKt9APURgw9B/JcOlKmU7yU21nlwC3AXBTPPwZkWlm0vN+kd255AkL5i
ln3WXWb821lQXe5f1ekgW2jqsvH+GHDkBNXIsA3HT5Ph7/yFhprx3uYX75QJHRVBldV5m8YqRiBI
HXmqa4D/RyPDYZfqkRDBpLUY/T7ZcTvkP77rPgR1sC+kmqBEAVuT0OF+M8NnTE3gx+GkEj/iHdno
Up0ohTtdIRKBPBPylh+XwvTBfIEYBYu4YevqMtXsrdZtHquaP0vHG/Gd5teHKznPBzSK8qnDkcN6
lQjjsRY9ii5igr6PrpP4q9k4FHUh6TRhCcb3T8gMyA3feSYT129eacsEge4drxyMKbnnovTaaG3/
Orb4KXdk4LgWwPCY+bO98i9ImeDvX+uOkA3DwuceSJFTiFisb8kNRwlm9jY0Evfs3AWYrLJuijJe
s4u083nF2p55c0zufopuL7LIg8MLBWGm+36NdUhKRcuBpmSWLAZeP8PXzNP+wcp6LrPAfUZme5o1
slKEn/ZjWj2IoHcEJri8Be63hETs4YLselurBN9M7f2QODfcyq2NTHA26HYmN7GOZrw3Rq97r9qu
bv/sAuNVgKsLTgVGCFv6x3bbPM85tG7KGZl2keh67KVrrSZZGnAiDOXbP6rEc0htzbfMCiBNUF6K
ccltTkMvCRYw8BOMqTSSNtKTjbpwE1nCn8nk1gGVY90GJiqAUzGzG/ipzPGi/SjF/WXU0ev3fN1O
V372wkboKT3V3q0O8GVgQH3wI056ST6/1q14U5Z8XEkh4z3vZ4A/jA4mar9gTTcUahShvwS9htUR
pu9wuq+4hidc2uDU3YWLJsRQ4fr/cleuzQ8mB5yKzP1Lz1CBupyTFlKUMZk3ycgMvg784wAFef5A
NoiefEevrGjMJr2/klNYAvy8UIzAyagZjcG70GV8mXhNmzlSxBvZh5eej2VgBCdGM1ZmNk0gUfSW
3yTnRwC3enc5CmRUgoZ8iPz6pW5jgFiS00yp0OLfu+a86/mw0GrHS05XHbSq/Ahq35NYNJ9dLd9M
+EIEdOyp3mB6UDk0T428l4Z2Dnq7Pvkls9ESDzKCEne2s17fptOvQzkCL0Gc8gDIJyDCWy1ufL/4
kkJTYCKjK9JJ3wa5C/HF9ypJTjh9rFoD1G7FehR+3zPmQ2c7YrnuBchT+/qBgzIWpXRAY1rN87dw
w4Sgf/5YnUsbq9+E1OukGPN1ZmcUYer0pZVVso2xmEHGG6UsRQysayDjbSeBtSDf0UjrZfBd3U65
f0GO0pSYDRB2arNgPAmSmvyJUHcTMsVZMomkEnTowyiz//oAKZqLIoAEbjl4aL/W2jculca0MAn6
wiJPYlczomca2qQp//7bPbDKYYpPU6eg6E8+RhKn+x11go89XpXKCdufsSl1pjK4tLZm7ldQtG9I
dysJs/KefYN4CSUjYD1jvjyrCHEgzjmHvGehuLeOiWK4/YN+NUJekaZIzFf27eEYevtXM7bV7RzM
pUjl9w9I2TPjsbhbxpLC278qnRTscki18iKNyYYo7NU8ogKV6fxsCOqvcWCQI3kcHBFy5LSIWBGx
bVnDA0GAhmaav7/rkvL2iwRpOG7DJuvW8r8yoMfrqMTEfp9RBOod7927PR0/cRU/zUovvr7QYOZZ
/bXdudzj0zOAEOph9UGBz5qM36bx++VcvI5FZzzEFRgxwYROvn06hHXxIN7VxiO2cB2MpAiUlxeG
xgeNUdZ3Oayq2EWCFzJ6NgAekYldIJPY5Sw3x5hIYE11C9mL5Pdt+zs6wseUKUOL6wd7Gjuhsx+y
qlCL7VuYJCzEk1XBrXjfmUcDyIfFJ0nNcC3cbLJmpCGYoZ2vqqv0TfQN+fL4dQ9c1GKhzShc39gd
1d3MzMGfvznb/f+pOFAdUUfCYHySu7SSREzmkG9TtdHBn7CpwoBya8aZ8bHKi+k4AuuwLW9aHQIi
yLRV7Ku5GrArPR82NPGmtXUvtjJnY/WvzpkVNB/4ju76dTuRiUysmF0MsTId6fyytOQuFJtoDmAY
aXeaGF2sSmrV/umemYA1TOEySsxZ+W4XJjIeqiV2FmFeUb1Ctc2GoCL3ZzFz408DO+RMANv7sB9o
66F/kpIQgiCkc3KaMpTe5eZnzhZXOKe+KqZOfJHuZlSxU/xwDGdZ5BH6I5HBH7pyzWFW8WflkjO7
a1Io18FOarpA8uNrb+tikNQxBDtuLlnYOqkybeYRH3SlFvdbfn8Dq2W+Ye4S6jYS6mojUVpBoIEr
E4xKizQHiC0lJ4IZGto+EVZ/yZMUyJ0lnQ0IJRLyh7R+Vka09JDKAr6b4RL03ZFK6U7hSQbRJW2y
s111eDjq7al1R+YUzvj+5iycfmKKsDfzDh/h1NlELT4ycoPYRdvH7nZBj1Z/RUqO0Qg7UhBg4JFk
zpofMDPVfykJcpjKXowzKmeHUUDt6r08l2bocJYAqRbndz8X1LacywDsYcrh8AQ3QOIMPxza2s8g
BYEAOztcYzcP93LocC2xXxiKdTjMJjs0VJDMqZoGwtGcqH8EBdZwnh0ot7c/iKz1I4GnV+mUrEJq
ryRZxH5TC5Av+m2QjpbIeG13lJyZ4b/1PSSlHM/AIiLVOYcf3gA13iHj1Q+xyY7Nh0Umkhvb7KUm
FaTkTUTEh8WNxu/YWGn8s4pQL9cN0xem7AiQbcOObVi4U7n7Df6FEgfTiUYA6q6IPuAFS81wAZqG
nDiTg54nCMd8N+x4tpJOhq87XE/5hCv9JrAg+commebJTrgbeRWkymd//Z9Jaft1jP/t5ErMMlKR
XqLJ4OMHG+e0DdAfCIvAje/W0tW+jbKVwO0jwlh1ICHrSHVIxGowvux0xcfeK8D2dhyO22l70r5v
QirQ6wpDxDvrAfSDaoRb7eAbaxBu94qNnPK+JnL9uQD0JWEOgbhlXHn3R1SfU5fEnGyeNk/ij7iy
Ri0Kj9vyUydIsR9nYkxE3MDC19h7sekNAtKaeJhNO1mWGVX1wbvnRaUV05UaObdSpxFQF2zgHtxG
4BeO75n+EL9nvA/M6NaBQrCU977Ow8/c714Q/RnnyUk9VSI+Erni7eO/NHMZnXoS87wzC8+pvhhn
F2X7u3vT34XRvfYUawaScLW3KwpPPDxp6byYlLPxIyq3OxJ7cYUgSAXke/E6w011z20eTDeSW2Pb
mxI5P0gnc5ywlkP1DWx8OCOIKrk6ctQfFcHVKXblYANOCHq0iWqFuT6fH6+7Z08dmlldli81vhaz
fFxs+0/422f78G1NWVU1MqmBNv+/HBF+B9w7/3asqEkB+cgmd5n5lpWgmq5C4ditE2xkfUvMaCmL
BzmUn5+i/v9GhSmlLFojxQOVpu8R0cjfZpjQ3J9SVeRLxRJY/MNvWRfSYE8DWrbb98R7Bfm07i13
UMX257yLhKK/3bdqU/IRYJ9UpPbTn00HbP1UbMO/TSPpH3c+RhwjrSMgKD+AN8ZMPjOYgrsX7MUz
ppdNTd3Ciddi18zzIrbtQ683rso3fuS6C/ozTLSWOtvavpQE12qfC+czX1ede2HavV/uhTyvx0WQ
mCUHdmz8SHrc9CmMyDkJD2ts2D4BGX4U6laMwY/Izm8rpj0fqnyw9eVlW6ADCgSEbUqVnL1jzRST
pxe3Z5qOPZo2OA9zzV6sGXDqeg95PII9GNziL8ZTX2+hngX5zuGI5K8b+x1Rj1gHfm2DOvmQG8eM
Ry8erIiwyaRVmlnilSdHxPmEKJly2jMvdKzCpExLQ+udf+kmZ229POlUNr0BuDOpX4A8pJfzvxwR
6hTqHby30C0g7WV2JwxCm7VuuNpiWVHktv6ezqOrrPtRnLyOrAA8DHosmUcjUVhvOFbV+xKkNPgc
8A4hHmswCm4lO+tYgBVaJRq43pEVgt3HNdB14D5JaNcsFAVmnk5qpRZNc8dyUW7S8gFSQf6mhuOW
PO1xocf3ILsJOOuObSFeRmc0BnFEo2JPBPC/3qYpnWv3FMNmOA6WCEDibXY/Ge9QJp/KADG7I3xK
jMtL/0PSGWa/xit3aoMKfX9F/A8znPgIvUi95c3dUw0ixlpTkvcTYwsJurhK23Ij0dVZk7o5P8x+
+l3EC8lNdQVr9aS7oTgpRmRkcSQULdCSaxPS2Y/lby5dHSC9EPaJphQiEX3Yu8Y2uNKMnY8yVa6s
EmHOJnXYjeGv08IlYNxFF30zkpKTzOVsq2g1nCQfaa5QAMG4jROX+lcL63qUK4HSXARF/RNCqqB+
K8JEusv6RLCVDGj3V+/PfA3qqC/oiL4CjNPCpv4TIGiX/JCOIIOGqy/UZkg5GjEG+Qje2Tjy6BS+
68lC+uZ+AOgjuK8vL0hjQWM4jFWmBscK8OZphvCTtAREnsb3SLftcInrZQS5X5xOmFZpan3G8XWY
HN7b3P4safDSdRPV5xAwcd5R3vm7XtsE/v0bP/l2AiWkSdRTH0zXNlGifvh8tUh96TdlYIKxtyTR
FRdlSSihP7prCBkVT2/XcQkCEhVtTHsoNUw8YpmseqodQee/63t08aLMEaudjLo8SMegxF2Jyoss
oe+EcQeRJekb/jbgBdche2lxMj79yrLwEpmbqD8+KvWGszwhxgMW5PXjU/Jchm4f0TB+BMtMx5R6
cXl9JweY0yP/ZyppD3Xm1HhuC2G23GcF2e52t2P6DyrIS+KRZaDgHJRPVBDddU0alnqAkYIukZ37
Klov++kr2ozFAAABT4BowTAAFFVQwwdLzQz/WGiJafWNOH3w5nEcMoOEGoLi44FLex39iAWwqtkL
2/ffrbp7yam4uCgkR+do6WvHzi/TEiFT6AsOzcDDVX+cn0gnZzM2ZzBWT8b/OLFSXGnaQOWpNrBK
GZPdDbqo3k6jS4YRKmMDTFWVsonLBxHzBemGu9qfhOYsRnEZtDnYzUlEN9cPbviiXWjNoupYslFq
I/CDj54Vt9rJLhtthXfw9awqV0wesVgdS9gMU1/6/iweCwQ8lecEvdCb1+8fsZewbsoBihHPUWt5
EKloBHn5bJAytzEAj02kGZWGRA3R8VrZV5bMCNCVIdiC1Bdh8NTQ6EDaI7TGoH3iXlH5Frb/8+IC
ooYP8k6pPIL6lrnHLVBSLGNuVytIM/Qclk34cUhsD6GpLKxgwjR4bN+r5N/FMmgaKs3F8dOJI2f4
MsYEv0c+UOHnK8bwG4TWkr08s0pXQ8qpsr16q5QpgPRfZ/oAJqkgUkaFvofMxqywevf4V4qmGhjx
3Eih8j6Ib+9utGEGjHOgMc4rJ5LQa6+LnqAbtePYFEeTHWg8VUfeZ8Hj3qoqR06SWQ4xdAOh9CKa
Lp0HygnmaI6VE20w3RtsSXSnaPQYjvFez7qUyvxsl1UcNVd/bvY+mqAItrxVWX3fuxiEl8TYnyOC
5R3V7H2V3Gzq6tOhkrE52CjPmh51tKxDML+Kmrp6xnH6La7DjmPXGjDLwaotmrGOWXScR0AdHZGM
o8eOLgO8oKc0bxPwr7OVwvJnIIrwtwLMfAvX8gZB5HJd09N++nltZLXgTRpQatoqaguFU6MLOtGf
hgxnmK0ksUfyLVuh//EhK1TIhPcGo8QJ3axgYlQah10xpRYHrxXWciU0Jkvgi7k/XtaKuJAKv+JO
d+/UHJdzYL0H/JiJwtOMnlG8eFteI95y9UyeEXlQahdudUX4BVChtrJsDMm09qyiQfVI5SUnxcak
oCU/FQRJ/hsjyFjLIxxSCmjU9SfcZolFN+JXs5D1LDZlw/Z+WGDByU3MgPcHVhZswafmIeE2Zmsv
Y1nwZ7X1avlB9xCuJbTNAxtUilkuOXe+iUxTXOsODUXMcebdEpxej4d59kTcrB+v2bo1eKHGkCwV
AM8jWwJ7CD8fTAbTJPIQVDvtiPVd8wxgwYk96FNsMSrAEjXAzo9CdnUL7VBvOxmtCt8A04acY3PH
oqYE12mB7IgSaQFuli8/rYAoM/iTmYcK/R1Njq2xecW52JsHY29at3qB32WNmBijGuRXk5pVFMB4
/VvE0wH5YwTeDfHLH+JA3twahSt77h54cxSjMNNjtD1200jf4F5YzOAq+aNWPrS9p6LSH3hWKo/C
RCuzoianlPwAOyHuSPvq1Z2sNJh3ySNZHdYOSGjg8a3hkEtF+FRn9Xwx5mTxzFIwOMy5YVl/ITiT
uBENwjlko1wC4sFH59BeBC6UUyMdqCJY7GLsxNI3al0lpi6HPPeJKP1iKW07D4PeBjAGCdbApUwu
JgVggijalNFyMxYdEbPyAaSOcmL0j8UIDLpH9dTQlqKksg5Ms9YZx8MMrw3KdAIrpoafx0a+yM4p
JQBpvovsj4wDFr/KrI1Q0Pe9D589pRfLKdR3wltZcxKn7S4dILS7Q6WwaUNT4ZbmSxaITSlGN6xW
qhtw1xzCVb1lNcRrspwDakIwsKkbBOOs3Xw4BahYiXHAmizZrn2VVhaW2cHCIjaT2qMmO3ciOx2H
Wxg7vfvhLrBiHfX5n+6+xUC5sB4PjHyU/9WoUM7AtQyD9hn44Yf4pdjc0viyWiSyoxkMC6pqaIgY
vYEvFBNzmpF8JKux8+I++sRsqg3bM4Fjh7m2HqAweKcbpUZHrnoD7qHSAMmLV2T0365qIgYYgTbu
zce3Fe9RZ6O1vUJStQVmcQD2jAXsMFRMZHJDE3+Oj5HUSp2g2C6DrnNvQJZiKaW0navBNUt8fLcH
mIx40xT5z7aGjjywKQ/ru18HsHxxL9j+qa7pT7SreQJTMVAQNeelBJRH2uqYU9z+S1lx+jTYTVqm
uO1H/a93afXRg9rapL4v4+ifxEE5J7ZZ4raxpGpD5Rs35Zq0ZBCqfImXTYKjNNMEV+tgXETHog07
QYodi8ztbJsVXcdkllvYaLEQSTfupKoOeyclyxMcL4AhoCMm0SVUV2gEuYhlO3+ixTKBp/+2v3Tz
DCmEba0JkiaYf0Gr7YEfWfbckPjMdSsf+jIAHPXY1drblz6OiwUVcsP/Pb9EQjio2xRqjn1ifRmp
MP8TGl8fjc5mrO7N2p7V5SDfSHfZWGcr8EYQpQZlb2jdSLHrAZoF0DIJoaMoXs72xQdty60IDBP6
CiluhEshqTbAhYhikdzJtp7M9g7A3kL0J6/RMwfav7AIBOWEl1NpNfN0OHAHRXRbgW2wdvgURMM0
VgfjRR+Tr1lSSBFeR4imlBuwlm2bGXjy4k0h6T/+4gdKhXg84aizrN0SbK3itumieYaQJJBb7QY3
HObnNfL/YxawINnFO6/7RSathxj4zfOwG91qpwHPZZYdjzWp1u0kWH0iRQPxqhVXxEai7nJmQ1aF
Vhz0ekqq7FB9DNQteBmZsrSX66JlB4I2316Y3xTHaYTXf64AVdXAAHjU1a4T8afjgL3OumNeP6Ls
sr6qn58k5cKTH77EJhHbtq3UH8Up3BtG1Zy7sPg+2K0fKncrurdp5QVO4NfttpzItx8WPSVR4YvI
L6w3qwc1p7Pshegg/WVgZzfVGqnPlwaYTbgmIKr7OOVn9WTpT0gCTog+BJaenzxGaYfqmDBaarzz
U/pYQss6fP6Yonc7S/ytN1jKme9KABQKnCQMvbYrNdt39uKxKCsXaaYHZHXyfBbSvZF6QPoPzDhI
xLTnUw5dSJcIMtP7K9J3jNs1LPIaoy1IMHid0gjuhL6+5Q0YI7Zyv9S0ahCrONBk+9ChDrrYc1bD
82wOfFwdKVGne0wdYpaeoj3DE/GvV/0yJJ/+RGACaRgn5qTQmMza1Mq7TXfnohc41PH8HwSEVwf4
71ZB7+5DlTLC38TFOszSz5/4eAsBTY55ZcH1181OGaLadqtQTIQTrB20p7zn3GYImGQjuCvW9HeZ
UdPAYW57KYNVdyPJ6CxLDQUf7CJq7ybBKfboxfF59LRgB0SjkkCKN4jrd6rrY3fCbEX9uDtTP6x0
KjD3SPqrAIWStbV68KyMPhXk32p7YWzh3P/MbY9Mz+8yDzZCx2QdeD5gynZFt6jAHRzPuiGA1GKU
4skCQnqCtbNM9hkn1G38Zv9PB595wkQ5TXDAI4LGL48+GTfRoIRpmLJhBxTOfN/2IrD1y/w8wde7
J4vsaPNrDEoroGLRa7UJCVGU2qb0SxOrNeAbvV2tUcpsdmU+mn0DNZC2mkfjtbpMmoUp8StDE51R
YyXDIcSPEO+rRT31S6dUY3f552bRlOE4N1/I/brBYDGT5mo/wvPPs7XjLedm6meAlnKr9tfTqpnY
zknT9hxM9MwEgU4Even5twHVsQPBz3q1RC+xbBenSRhZZgDcqDyBjhsJLblSKdSZkN/MH6Js5pad
ihBLlqh7WM4Iw4mXoobXzrPHhYqEG/oA8ibURFyuq8k5Rrr5oudhL2xUdHrrcrYtDeFsk+DmOaq9
a+RjzvBsdtlGwSC3pYkWC527CFG+PXqliD+v3jDKsiZgVsuBxgYtOGrfEvFYf/MMxAhloZ+Ar8hM
evWPXh0OCdf2B7buigyhTYsfxHeCqtV/kgnSv/XW0cTKrGles0PViPa2Rh5zoUxbCOdhqCxMFrbE
k+qKPPUW8CAByyzBkXqn0vGpu4f4V30CkR1xp0LzMXvUThUD7mAr2WpKdQPGZgFTJfDXOnJh2Fz3
mX/tSMDK9y6/VOxspH/5rqwAk3uax6kTDx385HXqkv6qedtdHMErcyQiSokOqkQfGRVnsDLG4AHm
sqPXoCEKR+VdVSUZo66JSX1PlDI93xbBTQO/QPEmS4I2+7Oz06HyM0jbFfB96jnpyC068Yydkml/
WSFf4EAqVo/RMF9dnFyBkmGBvYynJLO1Tdq1RASc5rILJRFaSSmde+4iM8v8j+nWso5BkuYoOMa3
7G21DrBRB6AMQGXJqRn62e8HmgNhbKITlPXrWNk/UJIcIXwgKYj+0kkO04lsn8RNayc00rlX87Be
x7m/0SO/NBZJzNjVoBH73SLMOytyrg8A9QTrvF7QBdm1EC1nip+3xBILQaEB+G1+h24iR3TpCj27
QVzYGqGm1p5B6X/YFfaNotpjCbvqWJvCHpTgoKmP4nSgeCjHF6Ca2RKIa8JgRXBucPbDQy7r21Yr
U0A4X8PFG1I5vwm1Dyue3hOeFXWD15VsonVD1Nv8YZQdZg1A+49XO0mUdevH68TtqVyg9BFWrA9b
PgfZaH6SUV2QpgoTrFYhYDH9m1flNaVtB/XdWR4YhRy1zmF7yJa9bMnXPCZc/BQFHDxoR7BaJfk9
HOafxd1eNELOH662GMRpZFAVNW3FOmj9/SnKAiCHBukMo//KMyIO4E6KhVjCbIf4ClL7q4HW3X8Z
6HS1N4iiswIgCi2ELq1pzaK5fAUxUu2EDI8peNqkLdUVhzOJKPJsUTTpRj35FBPMTSZXf8mxNFDn
z9+XzQClf3T/g+RkKO/5g/JCQfMzY9/87yICNbVyCnWAz8n4BhhWCiJWBIoKbSEuJWvOBc8AGdEO
t1QtXQcfFnEk9TLUCdgZ+4VC02gq75/4bqC572piuLCQ0v8Qo3/7SATckbRvVjmPhXWqp9SwdGWw
nlyPkBgTSXZWvKBM/MwSnxDUWXPO/8oDzSBvgGGsAVyqBbPYczOTXTl3KLE2niw8G2UxzqOcfoV4
PTQQyngulUKIhnCYSpQ4ll8joWkddYNo5jcA02StFTH0oU8txnQaBVBZCVUtfKlIxH43tuEuoplR
nmpkqBORiuz5Z9alep29ibPpWlt1xbKkIFtJpSW4QA6Hge8gLWlkzI20DRgUOef0aFMkiC0FeT8h
5fXUWWFAaBDSp23YTldd9jSQkrZFMIQ/Kll+4egOwFF0s6yvGt/LGxulnzEokKjBAgc0v/og8aOs
Fxl0kHNJrMA11vxXuup1QPd0infjkow4GIYI5fnY+Lm/Vr3ObQKR0T5al5GEiBqVQhwzRCrbYgK2
hE8XNmvpaXZwSq7f2omz2C2qtmzJJzuJsVoPikrwPjHAms42ZNp8yBGnePO6ZymRxoLyRt09Cpxx
+C3O35cAEg7nqCLm5BsiC9MUGPwivMExLpx3VACQ6ajI07Uj3Mxindj6vZZa/RZVNmhlE6IZRmVm
9krud9ORErQggMvwk5+3UqqAm1f1H2izYuVShMuDYC36kh9a4/NIMcdqoqxvlNLquT8uP5hR6Rmh
Hj13neKoAqprp9Plg+rNWYbtelICmD0KPdhOIPC3kPkvCrZ1+vjanInU2inwKGG7jBkmXpZTSEn7
RRUSLimvJ4e9fzJORwpYttZJo5ab6DlK8x1j0DRJ7pJBjq80KgZZxFsXvu85zGwId4s62ymWshVW
TtpJ0Wup3KLYK5KkGD8/8tAoro3wIQeNewPcUiGaJPqIOwm8/5WnPkCRYKRQClQGDIfAlP9Q9O20
fSOGOcQ2t+wRgV3UC1OGb9arbhZfB2OuKCl55uuZ3CYoxuh7PImXJF195PXpMhYaRxw08ywmIuwU
Pc/ArFFKfOkp1cFRTOhCGJHWbrmUlq0rrTsJRWiA2OIAiPnUz8hQYnERq/jYClophyn/b2gJ8HG2
1BeUBccvQSip8WTClR7yOy7cACJ3RjbmDZU4Tn73HWDGRiDFbDqB9aIjz+07ipF8GX/hiijFlwyP
uezTVP6TvFm9NpKob4Od+m+RGagMXOJ+ZwFNdnY1A8s8Q27jSw5JOQuRtoEwzoX91oTCqCC7szYt
gcK54uuRMx1ov3cXSa3MNiORzz7Mq2U/uRbvIGCjRPhGeOhtqgqC1KLlF6B0gksn253fNFdzRCyY
We/r8GwFHfb3/ZchhoOe96bxhKt+45TPPP3bwqYs/lCKb2STHSrWtxnMrkcf6q1O9/f0VLwmTRxW
MgApwapNwzfK7XoXcbtFqKzDKUrZyyRI41CBSlFHPyID8c87xcAixMg8QJCxiVVq2cByI7cC338r
vSoC2E5A1/Sx9YlqwjiXVEUE3QhXXtMMlWgCP/1EK7R5D8srbCvZKy06vn4X1WsNaKojrWMJ1PoJ
39/jSoymH0WV/2p+Vv/NJavrG2xgwn1HreuOd4h4MVaQj6uWslDHxyc7Q0y+mEtIBlSWZBHZdO1L
QzMNREGTmdXmQftyvIW+oAU76AX4W+TpsZSy5XPPnwgMjamMKbxoyBPo8M/AchgSLSawzPAFRRW2
LPVkxSTmUdJlVQMmqjVUtITHMO3xsswOKy8VFMcCj9Gr1fW6LSvRwX+IO/spLNVkEsxcQUWGuskh
BnWT5SJBkZFMRJjur2K8cYMcu9eLgPQeDRz0cr+MQRMrugyGQT4Lwbx3Ty9xCB4wL7TsEdGod9sD
8CDl/PkTyLrKlVf6OEnsdwMFCsYA9Cd98AzQfdFCgXZ70YrVLa2dGHh0tqezJsr2ps71LfkpTE2k
0t5zIOvHRKvkbkvUOpwKO0nUZWArkJy3FZv8TA4fJBYVbATIk5H+fhLvatcQ8SPQAk9llFMGfG4h
9sVpLzDOur0PyOef8oCoPD7siI0yQf1jTqcKZ4E57LvsNT2V3OK1soOQO0fUYcBsHJ5+PzhP0fBE
PcpKxBuHUzoCu6KnnN0W80iYSxYetUHLw7nqOIZXWj95yZxSd7NFltpYMKBAe3icnPsFFfQtUcUw
Bx9NIN487LdXlOQnHnWmDDv8XjvdNl7lfzselJHlmj8WUeERz9SFLcfNBEFD+2C9QuK4e1+sNuKz
8D3Lz6GmUr2Proa8yvbbUhBTdkusiSzwE5DKVg9AhWhti7utUEgWnMHIe42PapqjWYls2WS/7Bgj
PthGk9OSj2MjRr9gWRMgyLb7G4bfn80OO2b1ZiBkhD6Qj9XoWW2uqOCKDOzM6ybapjljfhZ6ILcK
+cgV+YSR9xSy+ASQxULFYdgMgHJva4AI/9/Tx61AXHCzSWo88mUxv1GueRzJoScnJPeeackhjoo/
hcyQm1jklvsIFgAEjfr+lCgu7sX2zYkVpZ+V3u+jxBbjWNZ93x1idAT88Hh/cqQDiUa6cqnRBia8
MgyR8C1IVS2Qi4dptBAdEoQelhO+9vjvcSht+lkBsAP88EBTOENvahOOPLXxsyeJNnnlAG7HosJP
Ok1iCso3FSrL4dlFS5ueRQKPqe+IZ1/5Hqcc/GD/H1cy0aZDPK9pNng4VUfrox37mcRSxpHku+hU
If1fbQ4WLN5Z+PyQuUAslzTM8yT0Rv8EvuC5M+oMCvstn5tDmzDL9ly1m3NX7V592XKtn9+EQI8I
TFK1emy5G2WDFdQiXidcumZQb39wYY2udcG/9O+okW4HZv+Xyd7vq6T388g/OPKmbw4xKqjSFAfP
b8G88DhEARjpGBg5hX5+ooyUwV5XWh5Z7kEpmDeGsXGxv3aoybWRq1k42ScppqUHQRgRy4Dv1UF3
gWl/rv/tNvckCAOW55antB8vRPEPKJpXfvW+jEJfSsTVBrmHgg7wvSJI4BygiZ9S2EfoKEI2P1XY
oQSZSK7ocYDEu73nRUXMaL/90US+drxVBdMa5lIRcrufLib7B7VU4GcFZuvYqq1dg10eTs+4jsPB
fXxXVcDG7VOSM2UCOw2nIl3UTZ8OVK+J6fneOIuE/8tCfNiHJepucTIjlm3uuZ5t8zcDsBeG3VVI
3e5AG40Fy6tx76mIeDH4qDZ2viRDCGkrhNCWUmUWkGZE5wu+lWo67c+wZAAl0IXZIKU3wHmO6hEb
e3H9IXKuFl8RdV6Z3Tcd2QtSo0ZvvVrvXgBXscutIGnCHkjlHwAx05w0dNMq7ONgzYNNLvto4lrn
Z3lkegO9XZ0DzGyO+LKI4B7CYM9zfPPQMRkzG2NysB16ub2ZXUhDHrVVzYxOp6LvXmzbjm6cbU4D
6Kb/KSYvOu4lxLA4R82MNzw/n5IwUR6iGO1ykKp6cL8X23pMDFpd5MGvN3Gs6ixlw9kK3ItjKN1N
bbFjI2YrJauikJ3OmegLW8+nywA0dTFj7kVRdZChzUcXn+YZ+YMYrNwpHzRmj9uRVjKXhA5bOM82
seGYAjMYTYAZZK9G+4ZdgXCe6VavQdwBYTJTI3Kml2JrvVE2B4i/InQdd7UR63nbI0nD3SUZlj+O
NwMSGbkRcriZK7QITHAH+KUe7BF12TbZU3bbyKLlUUOKFM9JcEfToMplhcjPyGW4upHd4EqXP7zd
6/77JQqcstyIVWJaEBFDL+gPTogiqMz6qelwabEj0TCRruro25gwjVjDHRfC/CuimRvn9a8zprQx
u3A3nO43HPhFOZTbUbpa81gHIJx18zwzFQQE+RelQDV24/JuzkB/itInQfww4NgQOo/PX8DZR7+i
do3DIdCDH1rO7RRVJ5i3BBbS4MmH0ZMT/NrnAJEEZUp/NfvWIS9N4iZKEPUNoG3n8aMUzmWhlrAA
4K+om7220m/mJ0Ef9vlmAoVqCCMoYbIzW31odYLGz3hHxK+z3nHL91xQ0F6bMpQm3pkJCgbyHh7C
rk5m4AGq6y2KKzyDsZSi1+NaQc4pLnzaUvh1j1OkElcD0cJZhpQ1SX86rqry4hVgebluaWorlFXl
WiZV7taK1Vg6G0YlmHrj6EhsuZEDIWl8uziq/j28C5I9i1XgNdGuozL7A1CRcJwnwk6ZJJA76+KB
GMgLw9lYPghbp+clu9JaCDkrNUZd0rwrM0LGt9Cc3eCBPiazd7lFoSViIbdsRWjwLtuhEz72/FUO
LHCLvX45gWVAEpi4++M/k2qhChpNFrlRWAcr84w6z+c/OkOwDivBzQw8Hpih2dek9bWeYGAvQxJC
/9pgmRONKiU62dQ+RWpmKuuYXtQ2vkC0oEW+YD5KBbTLdY0ztezXaRmi5Rl8aUJBcjjAYoivir2G
wAYzR99hi1GED5sVar9sfdcVZbkkGMcHUssElF5qGRvDQXpLwPfZCwBVmGZipbaE8W0Gm1Q2RcDH
Vk6tEq6QrsjCU0msewUQWQk6hXYNLhH/wVyOggNupGj37hImdyx9L5kG4oE5/ILri839lV5qZE/g
7GVJ3H+HiLONRk9hwIMJjQbAn2CRRbH31NbLwR4KnYZidQdp5J3CPXlf/JvloIR8YUJfnLgpX3ks
F7JeX9ZA1WX+l9/0htTPQ3rSHLTh7/OQA0egVOq/muAPWxD0CyhpPScPN0pVpBgp5k1FAdsAf65K
/Pvp0mWRtJjim38sD+Hl+ud+3eBQxUZoPHggCWU+ueI5BVSVsVLF+M6CE/uwO6mKTPl3iJtnENav
Z9nYJkEaluT0Z1FUpRiggn3pt41aFiwNELiy6PTcSF8PsdotOY/FbUxeKhE8XYmqLaiIiOnfLewS
/37RdK+II9MfehAx+j4x4iNVLdeMRqGqaqUaePXDYiseCDvxI3Cf62u6f4sEDc8DJFn29yBYnhlF
HCzlfCjyvOP40lSPOrJTuYc0ZsRdGUyFIBYCRejZ5pHGt/rdO6yPAgidYHYLpuEe61eHNtzU5Pdw
kHRw0dYKmE6O+0VHl/SBEAoVifmzdB3fUvTasKMADyD4xSvOfshIKmR2Gszk5g==
`protect end_protected
