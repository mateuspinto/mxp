`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 928)
`protect data_block
xXhDKvpLu1t3zlcKdTaDcKS3sKfexz2ufwmEcqNjM/ZYrUo5seeOqNJ5JHzUp+MMr6sh0lA7dxpp
gMaswDYPJsAydlv0k2V0qgUfMmH7SOvXh8bnPhqXajy9gXPyF4eBPps6fVfqqkkC+xmCj4Bs7kcE
0bCLZT/43eFD8Vx6GjAaX4xd+wCc+7Pa5r6nNu9y6Mu4shWK3PQOtI2C/brgKtLjuUPPvojiBoqD
zRRfAkBYd119La+/nlZUSy5oBeY6YqModMvOaGiRayfe35LSl6iTi8ccznw/uD1WsJTkg8MDr7Cg
G6/LbpSu9NIJhzNQ+UpYQ1PhtwBOlJofxMVgFcBSsrHabEZHh113ZDCRMyTHpn0rKPCL1g05rKbE
oaXT+mVbyouXTQ0+n7zGZvrPyJxf2DFve0Ue5b59cGFSEtfBNFrh8F8dKKDV3fdzsEgi/b6UOnd6
Luh+yL7bfgDKBUH6WdEvwDg2rkoVhUXq9j7KaRucJ31+IS0TvbDAx4xHRiBexX8d9cRDGQNnWjM1
pEaaENyHGIq69AxG+EzafLQVKbouD8t8dLDp57dFiCC1EvLnOJVdVzadHp3ykPI+xB5bNS3zqwLJ
QfpEAaN+eN7bRKEFeoMgI+t2qSob90cRhF2NX4CHZaqe2FTABNUEifpaZKdJpMpS0S0pdSrMMlci
n62GnGENiJl8yyirvjNiKpAhezu0tTP3LBbZhx6VHihSUBb84B7ybgljDEUtjgl0qqT2CbyZNSB4
E0L85YSpAND0/dfAuWcC1+rp3o5iouCvIg2ANRXGrflm4zT5yvDuKUFdQY8+AyfO7moB6UtD4P+A
PH1kSiva5lZeGxU980RnnhhQcJ38I0rugdzA9FTfxspmuNgIegmPdVUBBBTQGFeiWcQK5w3uqhmE
BpzxDHBp6aP/lvxNkjLgstL1q7biuw7bN/pPsyjM3H9RNpHLtwKzut1rm/asoK/vJGmjrkQuczit
3Jxw1Uz4hQ3eP8CCj1DZt1HrL0W2VVke4VodebR7ZLVKtkOIKBKal3jxAIvYHQt4vyyXbXzirq8j
apNBhQSA/IyOuW6g4OBmU7i/vO3oP1XKgWuu+/eGoY8dlamfQdqskJDmpc8VGTMkYYKLEuOTJjMz
1/DJLC1qsn876JRlhTvZqoEv87/dbY4OHpNhIfL7pkVDTABH+sRpbwiJ2yqz8wVNnEM9mu2NvXmm
Sr/VmzsRzqnuamszXfsyZA==
`protect end_protected
