`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7472)
`protect data_block
0USWSUGxovGsyBJteYpEoXZd/YEhywK5oRdvHV/WUhSlIjzFgiQXDBwfzZkjMUMr4q9y6QoF+BuE
9qkAgvUkUoaG6y4YMFvXXAWpX8E3IoCmyv0+CJcPBppiUHoNJ0H+HhkGWjYjysVBL5hCAUK12Xj9
bM3UURYU7V5dvegwHdNaGtQpH7fR4fYPqISs3oU3/tKMNF3bR29gj5gjVasFLTfFkGMMtKQksxkk
9AYSxv5Q4k9eHMkxXWVHqkngyiW7iki0twSG83VJJ1k1NF5qBUm/2pLCKPK20JEyuxgNkk2g2xOo
CxiD3ZeltHibjD1y+F8l62EdhSeIXtGQxCvJ756eFjIvl5iUjwrBquVdHuIhBMD/vPsrst5CM6v0
nGcROJHQ9p8fnIzUaCQWODRvY2Hv3FzvowToAU3/6fqSv7vpNt5IWJ1A7O97ijkS7ZNIub6jYlh8
xPkRvbG5XMgTaD8Y5J3D+jJx+brM/REnSY+bgbZ/WixtzUsH1kGZ/u7U+ijRFElfvzvSboA0+izc
73Ft8PtojbDN2/vdPLW0dY69KvuHFI0H5xBIKb04/BULPGGfiQsfw9hfsu0D8YuPXb4T1ic9gRyD
b02ZVTJKuSeW9KQ8sZAxcPmv6MJlLzPZYs3Cpui/cC2oMLA3bdq94Qp6HmI/Xdp6tipT/Ji+j9Xa
0C3dJ4Us9N2A3zAMmCKzu7ZdqioVxKO0YQ2sCYzukNCT2PP20ri4HyzeFFA/gR4giQ/c2XmSRgfY
s+LVErAvG7JmA6mdJYaQwK4A/GgucUTlF2MuQVRRqdvboRXW44lZmvIwDRhuHWIepquxWvoDL1r4
tCTPYo1di71fTqH5TmVYMJfdkbrWIZfzGvGecueBq/kzOfrspT2KDKBh8URVi7n1xEqnRXzMkWXZ
4GVHJSBAFGUFctlVak7Ft6O+5SJ1HhPcR+OWinjOTKYjzLqAIs2RZnwlaeR8kRuxwjHC15ztTR6T
PJQi5luskO1aiGASsYLsYpbcYVKzLisEv6PppcRu4t4Vjc1vYuvzhGI26JJBOGKXqeZEhoFc5wKh
lpQ2ZrCrR1AlptcTczZmayx3Ms17fxu333iY5FLH5G7pzhE/MbmJBC8mlUl0hTgmqH4maGfk6FaH
ez9h5f6KNcIVk95SKOiv4fds6C2qfvGRUA5r2NDrxHy5lbQrLv0BcxxxlUvl8lvipCEBWGTOxAIC
/7u55bPQWRtMTNEXxy3Q3dNXA5AzLfYAAW3uJmbDm6TqKtLXtXfsfJVjPtubqxhC4OuCbAW1tGLh
VRP99noBAIr6PxN0QYOIhQ7jSNXyGMVL00AT7PYOyF46VzFiYqL0HL46/CyAhT6+i/92vIZv5MFK
HNRLWs8LeUBGk7ftLi6y8CznDqTxxZ1Nebs8zOVVDFv/iEzRSAbbRXZaATa805av4oMHh4QRLJsx
BTQlFrrbe7+Eak9w4BUkBoM0wskflc5I8F5ErPqPZ2t6O696xmZJZwinl9p/ka2d5SjWeXQmtD36
s9ugaANdbgXTTlsIoq3tfmj0ePvw9a5LSVGjUOlIqERNZXZdRTn9dp3MDrtJYSwnZWcS6qmCRclB
PLYEItsVpzHJAQrA+yp+NGveAQsEKbLosrxs6+XBy/30cXpgg/PD5e+i12ShasfOz2EVi6OpGNaB
1tXO8PErmmXeTGrv2iGlQSULf71e8FL+uNUD3PF58jvF/FS9/7kypuXoQ8eShPVcdkyJLOaBh1uv
7+A41VsqNQiUv7c9WhDDV79FC705bpY7ONYmFDszPJM+yZP3zOyntDBqyscL4XrGAr1TPRC+nLWT
lsR+iRp5a1ty1kST+FOpTD3EOncLM3LL4Q4kDVPiQROfWH6/yML/t+Fvg5MnEb8byYO1Yi2NUOEZ
yKVs4wpwpQd6ycCXRQRSnOMGUR8qYpHoO4V5lK/Sukp4oLE1DSUP8rx0RP5QWPDnnbQ0vY60LMwF
llD3RGHviFA8vtb+/wYXoZ6f8Zhw4lkkSt+Ck8mACaWv1UJI+mXxgNf2dSjzSpMxz9GHqU+j6mx+
UuFOM31HBXnJGLgW7CawzgKhiyNIotC3NWO4j3byWs4gbbnHqob9zTh7Od9X7PWlN8AXd/zOk4+h
GfPyshXGVNjuJzbQxnXgb1o0Sc2cY7Gsu6NqwiCY6YeCgVGWYWJu1IB/quaMmM+qcLYHwDqvCrHz
5sbsHFEQOqQ/KUSoCForyYzp0HPZcg1e2ejSPriw0xVabiIjvyGcS3oUmvz764WN8GA3Mh+47n2I
2MiidSNmFLABtqJNk3NSy6+UKbVhqgNIcykPG1LJppKYWsqQls/LkcHFmrMH1w2bC0WmP0EQGQmc
HHNI2tnW/UbzuH6E3hv6NqYmqLbA2mTClLXuunHHUmYUCXi21IdlpLI2ehu+xLmuL464q7jajHem
sLwL0u3qPCSaUu5o9bU5y1PEdwInixB8FTiEJqY4LE3Hakr4/kaEhePqI1v3vF15429qbCAfjXlG
MfCQVWfzAlONh/InKCndqlmN+OBKRweuhNy/io8NZtttyX9cdUFn3guzpPy45Nzm0vdLk3hwle0c
8kuEV4TnslulGteVqKIyHubvCt5jW+W3eeeYZVqD9hh5TZVySpDOm6it7f6LV4TnBGjcgwrSH7dR
tHPgAMyL2f/Xo73yVHLHznWoQsmZHKCOH/SNvmoxIVUWKYqYcAtq6nZla1ldioBLagOs5bGBHZdc
Kgqu/WWdCskxXiMzlKwFQvovSOI+S95STUVBvr1BdDFK7+bnzScu4ynyhLjATpQFMpqcsDOMgvJh
l3PISC7t4ahNVYJAkkhsE2tHgFxAsWqcAPnjRgWYvBNvlj86JQNQkEaxPgyWgphBurmQwUobQpIg
3F83yK8kAN2QG1CmcP1Nx7nehdnMg4TkTnzoNMj1wLsmBzr+93M66plSQDy/lfLXye/dIikczcI/
IFN+yDTNLYsx9PXmIXJD+hTUXvCegua8QjwBxCFNjrhkZkRMhNu8Pwrgo9ah6o/KLCGtoN0f3xzt
x+etvjH3pdElUCpiscjiDxZYWZnoF6ax73Lt8grfMzQiDUUNVwSXH5zJE7Qkghuu1FUcrxsHmC8f
dfQMdBGX91Kxd2d8SQKZNUaKpTKHuCWJJ6ndvyOxR8HAXDXaNnzY0ytPSNSnuBBDSU9xxeOyDR7k
UUHIFVtCIpppXzzCARtcjWisRVYMd+SY5Pj0U/zfdel8WDTMJc28C62fkoU51MzqHZ0GV/P+PBQ3
6J3NxHCuYu/jcG/5K/K0JYwCCM6xJael9vIojYnXgZIYyXjO/1GSLPRlxw9Hww6by/y5vkHWesUv
fdEYe6BDhZ8XO1R3DI5dKo9IGhBdVW1K9Bvqv+EoW39TDfP3VXWAxjAEug1ZPjNtevu3lYQX79lc
bQSZqWYt0k3Q2eIkvM6ccB98I7/BLSo20sseUsAefz1J/6g5FfwWciTS4kwSsrwCtxp2MJrNWl8u
LaXrXt3R3zJrr8c+uKW/d9DdxQ2SrLLga2OcqZOQO5aESuxxWFavCZq+yhr9V6Rx5/zmjHev05Wx
4rTCOn61dyjqSHkySh1tSejxOtrhFUR9ZiHf1z5nwTBEEb+zO0i3rC9avkYUeNRvHiDkQPAme04a
riRIL2lYRg4NaW3n6UJsh4snfn9M8V0x5/6q3hLka1oR6vXgSwH5zS4h78racQoNU105EACU1iy8
ADYsFkEQe+rYKS6Rj2/mlzCLbUjQLtAgy0079tEU0bT9mkDW6hYcCrAWV90JrX9yWU6+j2ZX8+lt
MjGr0wRBzgpGXo6h1zaU1yLzyi3YC+emRx2UHkNztybE9UnUb+5CzSn+1xq2x1+2UzskdvyQ/RD1
zIbz9AMzG/LiBVH7Uakv/6KOyF1I7PKy1PeZgh6VZYDA46TL9Uy/AZjj2tmV7Zjgu3ERXXQQRJFV
VZRA7qx5lCfUCIiIYGhsrm4zogDV7xnIApGRWoOj4gmFa4axmrstwT9QA5aUIbwPVoMU+zOhreWx
AbrHTt+jSdJOuUCy4ggcHMGQJOsRTVt4jwsNCzg/rrBPj8iQjaaJ1xdPGWgYPrZSVmAasc1vIPFj
982VMv3nqgDkPuuEJS0ZgfOFGw1gQ1xc1bxVWsyXz20VAVRdBYjYz5INslFGNviLlCS7A8P+HOn3
Tvq8XVrntqwIVRrdVljdzTVsrz16G/iNxNZp1hcT4HQ5ZhMXTqZcLD/gwG/ReujxAQlrcgoEurpw
83ZqmyEOunBAIu2HLmAyWs+rpL8A21DcgBclzHSyed48TsCutOHo/IwBqnsC3Yvg/98bdPBr8gx3
em4nYNDumLIsxP9vtjYvC6Ix8QqO67SaXVm3myA4L0TIGgBLWtaAwceEo/sgOxV0rCV0DtdTFU1O
HpfIPwGCwgUH7uxvTk413RHtGIlM2Sfc/KcS694IlAw1l/pVeppNxs+awW4xeG+0yCh4Do3dAOoT
5Lib98/RjLPJQ5tKC9XJGt9drV650ebIN6W91HMcAaULh6hMB0OjIYax5AX12bdQoSeglushokPW
jg+aWTXrRQawTSD9Xs95leLfUHZLm3t8MsRBhNdhuPZUaGJvfB6Xhv7dhMz4q2QJKd4LeiuU4WJu
SUyv0wl09/9ZWtjXWQN1lrg3T5yll6cV9/49cjukLLJMs3xhj54XQ79cWV1G9CKdUiru883xlF9H
ExbyFAfmZgwmvU9hfkh6dzZYVkpJq8I+HpOiT0lRfcOurB8In3NPlag9QM3HyC+75N3pwJrq+ieS
ZC4EPKv/SjWcpf7s3golw4g8lXzgFHSbzCkw+BP0FR537heS9ngN+a4hw9cpMaZg2irO/1CDn52G
ObSuS7Cwn6oN4CyXsNVt/s4cqUvIrVn2vW9PEiBiUDSto2yE52Evee5yga01xTJ3/eQjkZN0msr/
rRDuBaxhUWfT7nsTgSw/o3+aXLC9tF3KU27g0m23MDk3tY8XwisSkjCOBgHJwAF4NGeL7VdyhHAg
GdHy/tzwHP1nULDa9tF7/nYT8YDRMTttppi6orMW5KZq/mh96PhdHaRmDj/AYXHHfOG4n/leKWfb
/90NqZuY8igWO7fR926QspNLJnIiOprjYxMzzSd2EDExPoPg3AkTFhq9OrP/1mPqny+HRbadijYP
ZJXuyfiLojI9lExExliDcN9IGibgzAwWBCCa0zwx74/U3fDuyQ5dJrCXYIRLfPS7PPzhqDCqNEzH
hLluO8jZNQDhIbZuz60aTLgKsBoHj5aMEjUkgKzXuFKFtacYnV8XAwnta9cBDRg/wecYBvUi89/p
wkoxZnx4qbn056B/dt3ooZAJf7V3lvG8VLmcwR1yUC73FiZ4GbCUeNeb4zT5SrrzyLvJN4+LFDf7
ApJp++luD1f4KmKA2SPbxWCFxkMmvKM4c+hWbiuw6EiXxXSmOZtlWOvrCB8y/oxKAHqZ1q9eFdpp
nKEyrDjYIT23xLl/ZNb0Ep9cdB9WaGZme/4Bw+BDoCaIY0vT79Czf0dZhon40N+K24hWjnREUrJU
wBiSov1q43XL8k5WXt7yp9+/m6zmPAedq1ahR56dblCHQq93F/aaW0vGnQRBygt7qQlarFLWUd0T
Wxnz/P6h3udsNN99eeWcETNgSNXIOpfUSux6W9rfDX18FX7+8v8kD29Z4ME3nNqKiJ6juLQG3R60
NGhaGzHQitlf3900PJkfqRPvurApUX3QUGDDVwXjEZ2oKGCrLNSkwM05Ss+IEYqL5IM/ch3KNRq1
Vi6s5Sl9IiHmK9BgKwKRhUSnUvt8glZgjat6Y7/4ri9sWhBFs7Q7dPFoThLdrreXEpvUJIQlgGwR
LKSAJS+s2m7zJayW0Q4YsoeJ9z0Zz1HTV15YWTRIh8HNVBZHVQyabP9Ey3uSwm/xw+9LuFTIXpAQ
e+iKvLOF32F7qGNKyv/Q8pE2c/cOI01y7JgCwQJXjblFZbnl6yj39iMOsUXuT/D3AszvWlj4Y+Ur
OmooF4yR7PlskDGO0NUV5A2/1Z8gpb8BtklQDfE+VpJ+iqNnfr0iFWwaZwaxpNGCiZwDhcDJxpde
Q8dB9ZW4SZczNDp8l7/mv9NCj6/w5tRyQbKg9yUU6dtUHGJ+u2HDVIl0fJeybMe8gEihaVD7OAd+
2MuZqJvHaIR/DVhvuy5blFxdTF4hLmTzAkIU1HzKBnIQcdhwMzHms+QdKyYBP7ocJ/i/a+5HmWJb
xhKe0CLa3KoayHrZ5Kic2NJcdlLx8FXNF6xi5Oiva61uSalup9DBwPtwTij5CXd6oyuW25ASTiSU
xhYxVDJEL2IcZ0UND83HI0mUK0xPMF8YtUz4gPsuXTXTLcXOw6WpETHD+m6C0AvD49042vk3KpU4
Xy/C3Nj8jTUgcY7uaPmFZzlJ00R7yWQ4yhDd7gQMGkRdmZi5o53GE9SZdr7V3m2PkOeEvlgiblsg
oghIZux/Ebq2EeyO6PHjbsSn2fscF3o/nFxbnJ1NMBJYaQV74hRcTe02S9j/Xu/SmRL8bG1rg/iz
8eCgJ8FJ3C51kzpsWF4BiiSuHQusB+Y10rIIN9bXqO3uyvTdroaYDTJZdSy0duI/zWxlM/0mhPdN
A46wrQaFyMt8kVNGfDl87wIA7Uv1zt3EjWzSINkiVRWsOWh/9b8buG6VfDEzfGp4MM0kgyPOqnx9
Ee/JlnJILUCUQsaCsyZmzCZIV0hj2uuAz8Ytk+vJiWLDhWLyqkOtMc5aELAKF3+LJPTxWIogMgS0
DJulOn1A9tuq//ZaEMKNBJ2AOS5WzkTyyRPFlpqw3WuLVULg/WLYBliwzSo3k7tuuKyAirIA7/Ro
YSvt/9bpQWpkcyFKsEjzYPg4/uMmhq4yXjijjiXJ+ID+I6g++vg61mr/6/1gcYsv5LL3FOkF1EcH
wzslB4Nlo9x/RdR5SdY3jNxqtYuVCk5gvU+/4MHfcRy/+s7/89EF3cPho50IT1qzTRB/YANZQUkk
YnsIet8TsNRsD/tWS9D6S6uWX9enR/O1B2d2j54I2yNrvSFb69MKA3HfTaXku9S0xvxLFgBuu5np
/VJbF69UluHIKweGAV26Q6QBkVevEw3LZtwJQ/s3+MXLOo83IMSWTHCwguPpatOvUFXsHzPQOIej
AIj3akBM3lE/zaw7lT5vcCpscrMTz/YmcY5z3MjSmw+j/DyPelJXofl0P+FIm+aVJBLr+VnyiZal
7jy9lVT4yuJOWM/YfgevNL3xRuMEFOcafCbyRkDDlHjDb30MVcQ3Bdxz9RUTN+Ngfxs+UhGz+hFn
e910JCcjXC/mf0b7R0OIPcjLhHiEq9n4tXx9j5Pi9MGFIHYwCAAw1SRc+VgZ1iZ+MMaK7s6CNH/r
7tjWTL0DJUxpkyIZNQZw4SyPlPyaPoCSI/b+PiIzm+NWSRa9fM8fv69IgBalCf39W/mMR9tAA2FP
W3zvnTePGYp6E0u2tMRDsKdxrYUcUonNpae73h2G56KTR3ksQwjdlwgBik806DAAsaHJ9AlcP8/G
/ApI8j6xE0t9XqbQxONNs1Y0Bl+M5T/Yy0pjtUajhFZZd804ElrnmoJIRv1mK8gu9L5WOCBpxpYM
a0FJ+n0HtxTk0WfhwaeZUhmDvMnYsQShaUQVtQH4odGG47ooU3B2JUWdzflE/MEKIo0nEjUj/XCM
Nuy4SOd/RhX41WHeKW4R43uNswnn/Yb2l05YnGiaqrQTH4x3SBd3+NMHFRaBOl/7ErMjElZmiV8V
OOcJG1WWkUJ1gPQxvtclMqYkeggqZvhRSto+fhLJsc/AqhmgbtM2fIErO8v9wLlUDrxH8+U/tMN3
zX00kHTQBMWg0wFLL8FRBAAArju9PXVU9hDnHP40WCeSVLaRkkwycHLj07Qmg/1Ob3rW7vPJJxB3
WURNna9+UQ4WCmZw0RNER8u7GgfVVhNXeyJ72NvzoXYBVB6awkOGLTH93Y9t3axgkBpIuXz/269E
jFjvQQFiks/IGwkSU7xzZABlqk6ALPr23eW4SDhbr+jsGtlkcqMEliULbKLLaHr9CL6HFD5vF7QN
BU7r/Z7/jwPkZFfdOtgRQfn4lQKSsx6EBfm0oVaBwzvD9LHlPedLct/VLtjh3FfYIQQy4pdTUdaV
It2EIrBaFwaP9K7nzgcd27G96KEE8lLKo5cHG2n3NMHmTkIyOZFpiFNFfCBasURhuUV97Q/1uM3Z
ob/10lSPMlcspbJ1tRSMR4Lv3tcCFK+BybIieZsA0TEWVFrsXgxIBHktw7LAsN2tNOxM5+dkPN1k
pl2d33rcLjUoUeteOB+w7/B64Vzifq1pFMHSs4i8DH3EJEaz8QTyL3lFzt7ur3sFscixol1f+cC9
UBXhVuAbNuTBtPSnD3QF7HHersKnXTXfj4t0wINhvw+Pr3EKq5yfgFrwA+DZVtMsLy0MgRONA257
6smX3G7RqkHregIPIdh/w9Lk8SB/cm4+FWMhBKAYopQPUxHLppC5e27NWBAAA+evkjPvUYkbT6bQ
Ncb3vEUZbho3V2ZI8JHTiCpo8JAm0s/v/uF1DSR75hT9LVM9ldaxH/GmYzOiHqCVzopKWdOsTKXs
CmJ/f588TNMGRjGOiB9TKuBYkrg9rUP2W5ezjGtvcfL6TyHXRQ+lih7hVQKwD4rHaRw0XDKzpZSh
3oNM1z5ZvcoMNetn95Y2BAcrFuZ51nFu9nnK6/CDC7KWWpj/f9qRiAZUkfEb2UXKs7fVbwslaj1O
QTJfxA/sErd2sE6J+GVcI4HelNnQXZGIo3mAFhrLgPlznd8aLhPal/sJuuhmwZLGUeufvMMoDBhU
r9DV7qhfeOVNCW0qBKH+wK4vQfnz53+GyFXx54PkxJ1DWXu5fjEGOBcgd/a+V/uP5UiNrdkB25zK
xkBMruh/7vV0nfAhhxv0wVkbAETBqDZNIhrYJwd2AU083uu9+mN6TyEgB+wCSZKXD00vAQ3aex5B
bBDPl7NqRRgv4iZEK7WNn2y/8QLKszn/Xeos9QU3drnyzznjogJG+T4SzgIjUwknrobmaty0rN00
eoQcdIFbyWCIdHuODReNw23Ier2dAovJhxS2NSepmQKBt0V64l42eO0Ra+6OXFgrHgFTyDCjmugK
uLWBBIrNCFJDcZ5JiRYkaXzEPb4LuajWiUl21Pkv3SLamowt6MOCc9Gp/2M+WeHStDf061wQxSDr
8oQbzZFrpJ689ajJ9BfbPRNET6/9WckpA5PNcXpo1/gyGn0vYnv4BrXEGTl9SmUEuqhioWb7F/VG
K52YSe1ekKqC2F7UvMnDpsWoW7dgYfBenzyk97CvZ8sJTyGcM9oCDMw2aObkgG5yKwa7fXrshXH1
REOUuDVvMdx28riT9fuhlHnmASBvKs8E0coXqpa/AGl+RaCFdcsHa/i6A8SvrvviNDwahm0yo2TU
IZHmhBSCDr0davU8eJN49U57QExhXkv/wq13CVpxGMrWC3o6CNtGSRyPiDeuEa4w2omvjVk0ouPQ
PbjyF5REDJ8p9nDn1i13Lm+/KuSYn+I0EcZIZD7U9lI9H78qnkvrgir8dQHBB9NeH9CQ7hAPYbO5
iJOhjog1xjeGrGfGMjj18BqlNxvMB1wQR9P3V721AfXg/zZqMgIUc+0NVaKVj28JWykiTNsIEGio
FeypLBuh105+ZDQH8LJWYu5wrI07mzJBqzCuPlMNG2OoTfzyE9rCDhCRLXPfWL9grvJEFrVwV5x/
jhMjkd5Gj3cGptKfgd72K8DHZWu4C4yfGkbxTaBC9W3ZK52VvhIjmo4Ou99FhdfJUv5qEYdYsYl3
BvYQPmDHmZ2krCdLd0qw0s+Am+n4cjNyv+5GhVdqdnSXkIFDP0gwEH0K0QlfKWQbWRKZe5ltvyzd
KdNEzm9IVNtLXNp6GmjvAgS7NkLDMHIUXKCGi5gqckFEFoDYn2HyWQNxWvxsuBkfuOsz101dqaJv
SlnQzJ0=
`protect end_protected
