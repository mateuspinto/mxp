`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 928)
`protect data_block
Qq0ZJiisYfou76PgQULyN3iGODU74d+pBP5oge3mtGBp/Nw++Z8T/TysNnRoTz/92/OpMO1XASY+
vhRRe4mI7Cm15Ohc1+9ZDdYFa6i/5YkZxGA03CO9tQnKGG6EtCjJksWbH+/eUB/bTJxcJWNh4vBT
jDwBPuFYRfe2tUEg7zsJC1tWmVu0Y86aySXvCHcP+Hs4sVHl/Psk/WioaQEf7oDExni84HoiBfeV
S3gZfKIFIsAJ9t3op0iBg18sDWikuLfl6J5fKWmW/F0dG3bieEyF+iMMf6iTh8AJr1Cynk7fkfkI
dXM2GjrY/OawYMkE0PfeAlm8WxyR7Nh9RxImXF3vAcoRRnOv/v9FuLWMfc1aizDHrqWDdxGiFVLV
r89s4uCz+fQci/ql7WqrH8XFNGUe7qARH45bhhBZ+O4C5kE9Sm/aDvBIR6hQ3hJ67iKPTRdAsMKD
P8YPeM/8ZmEwDLTHZ8APVuoryfLye/HY40K+P7pf+FmeM+VqhvYmH/uMHYM/vQAzXNVL3KPsvU4y
3eGVQyVMrtHegl+Wje+9PHL3tIZCTH8OAZTy8elJAzCJKXIk0iU9rXH61f4noxtmb2Ca93ZfQO84
ls1bsBht/qtF+NEmrEzsk/nyUNVD4/rrrDWZJfES1hIEjaTcRDlwVuCwAQRDgzs+fQYIskoLx4DB
YpXf8kb40aRUTVIL7WP1SPHmhIA0TZk0FtLlmYMlU6BB9dE7wZcpFQjjcLgxMTNt//Fn3CGP4by1
eHbVrxAQ6sOBWYpeYGqdM88ORVLU54kxHn0EokGokYXvYOBEATXpOHzAs/dnMyqR7fO6L65zlxLI
fPfLoXqYGjmVLIwckM9WiI7K7hbNY8f87vFNam1eIrdSsO+5YfbPbCSlAyMCdG0Leo2ZwZu7kHod
5LKLEipD5ti+O3Kwtt+XPRuHnUr6pnQ5JMX6tth7WawPOWfOiOGTKLJ24poJVKJfEhqJHIts3RYq
j7gaPH3yrhuKt3l0ySQEmAp/SoJIc5oqB0slWoCbA2HcOBYs7XGlAtiy2vyef0yydVgqwvAC4EZt
sGZEt5dUMDLEdhjLMxCPdhpgZZTGH+njjeWMQkpekOn8Y0/8gKl4pzZJoFDYmsSuoqugQKWlgpvw
YRFRbtNKOCq5DW6EmX9XgBQoxyvR8q//nBW86HSr+qSkgO50BUrhPULdRTIZOCYEIXfgZKBdq7El
50njQC0C49HO6+hfeC9vlQ==
`protect end_protected
