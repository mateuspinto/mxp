`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2368)
`protect data_block
PbY9osurrkKjnV42BwMObpoa9FJMes/mXZjCRdXmmSP2NQb3TYM7I3A23U73WJN8kOggbXgSlPsI
AAXZ8HwU2EcjPlC07cLK1qWamxkCstuJDBaZhAjdOPY7Q/T9iyKDCBEENceahe3s2+JZDybo9WsS
8w6XckfZ7PGynmuz94lyMDWW/64jDaZQzjcLy+OXiPs96WuMJWSw6eGCF37iDFOrlq6QnFzLA1NK
zpKyHanJHDorIPpq+j/pyDIV0DMRew0FQYxIAkmwD9S0KKq6DXEntIihFiQWnZ20gPxmHHTak+mW
PDnEY1OYQey6QQ4lwIBBjYA2HKz7eesgmUC6fbPgLqBVqzpf+A95d3oimxQz8Vb3SIjk20zR5DV4
yXqCONfsoANTGEVqp4NLmGevkdTqTuUuzbgTGMW6jkzMAGYbQZAEaMfx/P/x2VONaVGNlDbLBg48
hryV3JkWG+wkRYLSwsGW2lUHU7Co/fXfE8wHuewDkuIqu72W8h+sRn+4ut2YysmsIkj/nz4k8mM+
HGqSRfb4SuNhJu9FjnpEEJLsbO7nb75OUCVQbqF91CFSq+BlfPfMogysF6f/BLllFaS+vkz6AxJJ
I+eLEIayz7q7HEqV5W6eqpJl3jJ/pZ0tKsqwuN7qKjQd5PRXCYrBlEKx0J9UYAi+zU2bYSsGHo7N
tDJj1npOr//DnlWowp7YzqPEd7RwRAnuH1UjHgIR2jSYZBqxuH94oGnVmIzNuF5F7M0+u3U6TJ1z
rrxIzxkmzvc0HjFT/eE10tNWT/mg4SflJKta/lyyzRAUpEXug6RFVf9DWZ03A9YKyHhYwND+gUW9
8Ahy/X+GY/J8ANO7RuRKT+sVjkeSzw/7tgHKip9z9zeE2FzpmeR88ez3sa15tN0OsNX4DTTDdr/O
Q2wEcqGIco/otNt8ahujxAdeeRFO9etyXfZ6gPmpjyB9LEGn+71OhkZMUHJip9MA07z/qYSPRBlO
iOPdzXSax/ZqRtr2zzzMSkKp0jq+dCqfZB0ErA8S7ryL5rqVmEvlYOcO6Og54pBUT0aWOJQ+8qg+
LL9UbBFpjUBt5ANoLMNnvIpoTN3KIu5aUaWnVhErUt7ZskNkjK0TPUGWrxehIiIkdo+GnzbYxh24
Pi8jMURFcANe5Nh7lhLNbOjBDwB55wtSBs3DeFkYmpV8IyaTt5u/Owqnx4uOolPl0W3yg0A1ohAh
DHibKxrJ16o1MmegEtnLkrumAGPq/z143F2hET+w8FjnJCnPsF1AmvCwSd/4qJMteqwM2mAMNqkN
VLuEqHoJNSsBdSQ0iNveMnN3tAOyhUTPobIfFl9EW7XGD3+M1Sj/s5AufOxyiCK+iZ5x7BwEZsZB
R4Gvjp6uXzfsiqxbr/m5YdGvpo1CvzAY2ulF/1KgvXAbi2gOuwc+ourZVZbboK4R9St4ZW5cu8NE
4IGnopLMBOpc+jf6lUxwlrJuNAVVzvsV7YUcKg0DO3CHZrMmwfVrJjXz+AkDVbbEmL+1cAmGs9Mb
faQ/klBj0ukJQgxefMw0ZylmPMeblL2Q7jRjxELIcgLnxoeMMUZgYNGjMbZ8qHhHeAEZR/ZxJnmd
vhGLgA8WLvAG0hdfoM4YKOmAG3cCC4luYln+WZNOO5kTkK/n+oteYSd2fyRadBB0Y8ge6NjChUC6
VpS9QMCjXpl60q9TmDWsHduYXY/KkmMGP1kGiJf1G+RWwMCJayWx62kjJVdDz2G3+PeosymiqDtq
nSTC1fZF73Q3VNW1r4X/e/PkyKWnUK2xFsFF2wjfRVNuDUYn5S7YMM/yddJUGzOv5sa0zue8eROC
YyzvoyIdxcI01LnTvpHv97IWJmhGslkdQFq40DD1z09mxPQY0DZytObRdq8+skTvBXH27CAx/HDg
/tqtUy+iZTw0jRVvfc8dYcsRzmwMIoOUcIxjJpS3Zg4HJ6g60UO13Dzhw1iw5mTJD71nvkzar80f
s5hkEwVUo/It4UUBYVG0goeagNxQITHTJy6xa279oCGVunAi1pl6l4C9GlZ7xQ+RgKTQB6O3KnJs
cC7OIJQEy94VRmIWkLiJ2MT2TRnikC58DuNySz6rPK6VLeTVTXAGCCzacNd75WmFmtaO/W/8jou3
hx4xE2nAEGjQ2bW+ynREk9QGPRxhDE/9sa/QcLR3yFtBr8nwpzsCgM4M2Rmh/olNUn76Zf+Qwq7p
9QQw/8k+4NJKnou0hV52jBC0nT3apFkvkQbC4WMh6Ym3NE40dv/GVk1rAsrCbnKTafDif5x41KeI
Z+spKdmnL5Ppgbg0uX9Q7Eequm8lJIvw85KgRVWh/d1VimwQ3utRlflXg1qD8ziGqPpP8j/pouWg
4JcEQT6DSsNgCcZsj/70GF5XVkg/REWCqU3if6u0oI7Je8vGGmqMn6oMmZnjFCUCSfWgDlXXK7ga
WfpC2cOcn2eZqPgPwmwStOmsa4pI5NKpVTqxAXA4Slka0+huIOjnY63kN/PJMMbdqaOvoXIXtWmb
2tJs11Il/+QIbdzCRSOEg9DFglIDu2WxTa/hR2YKE73yEXFGmzhwhX1PN++lP+UlUg6ZvMZGBmye
0S2onydsCpKftNZkrksBA8bnpcnHIlSrPwpp234m0fw8341xMw24Ths8Fqm/ZWKRbzU60dKttAwA
6JWjihJMBGMJBd7GkF4NPAj0AEXBG6VYKz5xr2FRYmRmb/uE00rLXMw8MmMo0BOROZgO8casUcpX
tjZdbKBAAEmcAmrgtXi1LLqP1xfqgHMF6O+KnHr4q1tmuoRYaq2ixh5SzTYmE8dgnmxT1S1yrwyP
q0SJ6RMz+Fayymg0OHKYSP5nAMOSyBNz45MdZjczZ4X8cxTXJ6Fo1QLA4d4ke8mMeLqu+L8F+3NA
OpMgjDmUA1UVlqpB+avatZjJFt2L5OvZg02Be0q/1t/QrVYpFbP2diwYAYFfZ88cEMezCvwYMWPU
161IFcvtWpiKUhkA1SnX61nf0eu0rhNCQiYRFWWUEf9y+X6J3r+o0P/xPDyoshP9gBLYpJfTCT2g
nm1B+7NUPN5P9yXGGDbP+3ibifPtAS/MSWIpC2nv73Nfie85m2utc+phMsKqoBqh9h9sTxIM2h93
VOlkmg0ohusoJdAqyZ3Zt0o0fJ+rbi3L8QEYAI0EgQ==
`protect end_protected
