`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74304)
`protect data_block
0qWIOUAYKnUV1dtnGAba59WgH3uKGjnfoN+yPzoviuBrSENeyBXlgSUoXGZaHhaPRLEdEWuUW8e2
td3U4k66+kB/6xTTiIvXzVf5UvMc8kfWzGswPuiFcgfp7fCAICP4OSQVHeNVK6QqrT1py9RblNnm
vBbH7e4g+nFLOQtnzoUQ2wsJ+LCOapzNsxreFSlbuKVQQqPhaY4DCFJrn6JUvDE/EOsBFFao7Ti8
6u9nPlrMC0eobn3ffAGO3BzeVssIYlLMy+8WsFm3A8J32NbnleJQGE3LAsxxiBG5Y2yK8n9vXAb3
nzUyAj2jsnKhblTjsEfHufFwhsHxWa09Xk2GewG+SuVs9w589Gr1ANP8sEP8YoXo67bGd8JtIcB9
/yaESCU5yOh9O5fq6HcTpimJIlIulF9Q84JoGwTFv378d5ZI6NMpaWz+sDevcD8QVmvMG1pP4Skm
jwE0XM7VKJtyEbY2h7tTCSa6DyOqI6sNmtdzV6wa5hmL1P3PyrVC6DDI+X/2cYrAkeFZPhOFyCof
9tUq0pavKanhqafCEGPaIVYXrODCG00/gfL5EeqRnCMwq9HIp5NQ6gH027+fj8Xpy5nnZx2DVM26
GUNrR1V4/a+WkDID8IhrZCVthTMWNfEeRBpNsBGbiiz0TJkSedBSIx5N2D6UP1CDNjVpKccrzRIN
ogQrkmT9qJKEj+hL7ufrBwRRBbPPEidUL8LhOvpBedakIl0HLa09bCIIjQoC1vDW1W4J3mDEn9oz
lJ/2WERis00PVbwPQvDDdmMKI78ugRlBAL5TMVVnJa/QuXzotUSyBDunNBcWqxII2lr5pFWMcedj
m+YjKiPoZPm9U38wNIoDIGE2/6oPPuS4rOjlwKt6hkZ/0cLhAZ4wnCQRpBL2iHhpEbZ5qk9hDx2k
mkI9vT8j66jyrTP7r4EUzZDwsnR77e9PucM4PXK2MvdaEL62oW/4RzA6b3pChyWt0MVlpLGqyzub
vKvCS5eklBsH7NEGO8shKpEE1ylSxwXKYFyfb8Mlgj7uHN+JwI3FOceEmpMEgc66m+DOF1s0kR4W
bGhoLsRAucmPLsIh6iDfxHovJCEFULs71JWYJYlTMFC1a0xCfC/t+efd/fnmEmmabydZe9Ejg8bL
qvxYy04X4LjggC/YSKCAJQgZGVDDNuPk321Fo1hdTHOCagt7sBvJ3V0/oe+wpUgd9QXrKqBF9Cdb
jvtjO1NnbTsMzWRGsiCz0GvauJSm/O8jLBPUao7DEhHJQepH9RguSBj+n3eBAHpVNLVottT/+MO1
AbmVcHsxR3Ordnw+ZQK940Xrr7I56a/uiNQoAB+uZCkrACE3zB0UNupeLK502z4zqOn24Fqx9X9c
rqTWuhdicZ8fIUazy86DaoKwexxlF/1foABNmCziHtqk2AQ+K/UvkmUpfikySmmNLIbJlFmrrs93
mrZovyW7gjJ2BTS3aeqCtOoJEvqDrTtyyZT4276IFDS6YPXwTqkPyMZO8oZ6A56bycMOuLkaXz3P
bBpzuPON00ml+gnTHYtQEAXLdO6ibW2WyhXiGqFvqo42OetjXvsKfLgXwoNWxsHZh7cFgzo6zx8T
D/NERrAoZIutyyQGO9ug4JES4vkT0/KegOmZttrqJ8twJl9VRe165wAz7bR6G0Cl7hLzV0wP8PBW
IZdhHam4L8enL0iqixIJnCcmgsHD6tT8vXHY6R1P0g5l1BPdcG64m5b3hK0Ze3x2aRj3YrU16SdN
QmH8ZSCohseNWKF5zvdfHg6By635Enkj0mwtQ2C3ve5v1eHU5AnjWA8rRsdtoy6fWk1CN9jdzabd
dnEdrEVxUxryDvoC4mAkwwy46XJjNmI8M3jPhwcspqN3xRpS4+vUCXR+0IrEV6F/LJl6dhuWVl40
zM0r85RHvgUC8DsUaYEXT0b8FXcmCiwL/zNwALmYltFna+ZaY0AnJbE0RtZNQzZD2ZHS1+s7Jq7J
fgRSqIa7Vt8rr8vvhVMYrxFeX3HuufcOQ4oSEbu+hbYheyght7DjI8o5tWol7fTlsFbhSLHNd9vH
t0S38Lg9vSpn7WfH3PAQd0tnEDzjA1pysAKlflmA9MQ80IQpO5gbAcYiqmlwjdvqjj+mA1A0jUXv
h79u1Q0EVY29gJEaHwPVZISY3/+scaEs5qMlKnHTnUcbaROeQN+WQQWHadnQ/rWp0LU3b1HCYvH8
sG2mRAMsuiYM/xszPkG34oos26FHOMnDPUiXvQwDTxaXkkNr93DFu87bR3KGoVmU66s/hWa+XntR
SHpHtPG2PLH1UNu1zsz1/p7TWElH1xAG83kR/FAc60lyu3TsuUivPKCaVwyX76QOUkqwqEYUlwGt
mGWgJD/Bk7Dc/Gs2yQ+I0D1YynkJzX0FcoWgTsKpEPKW76MPwJIJGt92GAJWKDCTcQ51xxVOgId/
m7N5RU0eoSdMrFYHE36oxRlqAK20TnMC0phbJ29y8phxtVd2ypmIjrHdc0O3zFQxN7VjBXQwixWe
c9/V4PFKl8V2yxTe0Jx0FciWqVUA+8E0paIWy1clgpmfwbqPc5qtMi5QA4dA2GaY0/gzVefIvEuJ
vVpWxsJvU0MxN9icGJ0lDWDEF8OlOalP7FdugPetlS5a0Vpj4bvKh6Jscy0OEmrjXDMAWZ6v9qs2
Lr3Jd1UzTtUXM7ZBz3OD3m0dyk1SaJbOrGCkSYDgWgHg+YZ22xNssqIuBUx7Y+Ft58opggXcNcFn
B48bsFFIVylU/sONJqYtxjnx6O2aKFYMjpCuTqdSsVK3f+HKNXsin0r8TLJIIty8G3bsrYlQfrgP
HwV7P62ELbsTeCAVgjcnaYmQLAYxgqARYN7L9yjjZJQ1IUdZ9MQBq+t64f6oojhOVBhATMSPtriS
AdJCeIxAXc3GoRFY24H76xcUwcJK4fRTRLIGjmph0QPledHajR/qixtXu4NcOA4ehWEmOQfDEoXm
3rpRqNWkQaLz+UgrrtrtnufeB65ZuGPB1DQ2ZNr3+zomXYkt3UOY3gyw6n40XdKTBHYM04PLmabw
ksr+vtIKEzXKN0ECeq2ZerSJX817Kuxs40aX8oFdj45gdHF7T7lKj/9VdgmRJFzuwb4b0a+LzNzb
IpQBNKFxGEYxF5uLf6YSvbsJXum40gGmqBNRCEbRHiNPIxBACmCrZQdKsiOzAQCvm+KlDBwCdgMj
8+NNQNg49OosFicnXZKH4PModDStaXFpcK9DMZIi8PAC5AyPFboXGqhK0nspUkZSdS6JK1t6m+tU
bT7FxyUSOVi9R5TbKiXg2X5wJB9AQVvzYt8g8qqWFu7Nu3xfyoMrgjm3CSyY1tv/Yt5kFggj8kAb
DoojBY1hRpvAlA+bPBnOxZGS1ha0wVYR1m4KgEqy9u0pbUJZYt/uq7t3TnnjbOiKu74igqIUtXcK
8F62sSTsXr1kOBInaukAjhCzds8tU2lg+18auOK3S30HtRbHhJPxkfQcaaAMuJpiQOmDvYqBCiUt
ueLcIdBChiTZ/HseogCZsFg+oxu9R6wtJFi0Y8gETy3swgLRuj29Q8OWcHfdL2ncPtIRW3NOnczH
PcO/uQhFzfApb0BvymTqIytBJNVRL5lvowatFCSS2rOhF9XlNmn4X1rwtDWPBnus3vx+xWTNoFVL
dpxDaKkdFmxQd8u19YiFiGjyePTQsK6pzu+lWIKg0Y4krZC8GfWa0CW4bvoLDUZIHMOnFPevuyQZ
YwoR+1kULZGWTVZoUnM8wGtqk4WvSG9pj1BO17aGbaeMIAWk9/OkxayB9wCzipphd5K3TUxgGlVt
NoZkbbXcYHoPRMB/UtGkuz5Jnw0gyVkedFEzB759q22LIPVCZeFBYH39IOwti3sFrBhvEWbtoBra
0sA4pa2zckNklCOwHY04gPUugrIamy0p3TYZFUkRTgPdGpKPqgFSR0uITdKcIqixkh9ezsOXklqV
JhdrrTmJ9r9tuGhg0KgNQw5FOTF1SZPPmYljbFP94kmEmtC+JKv44Yes46GEUJxsOet6NQ97pPVV
9qmL0uFadYp3DiauuqWmew/F3tnt+v1exi5bQr/+8z5IsRVrObolHZP77qHQJkkoCNNeVPwRxG6Y
+fqBy4BNUqX6TIJSDsg9Hro9qehzGCzu3HZqdZWhb2bhgZ1eZYYvNQ+Q0nlsst367RHEgTmnoPLv
G+e0FRptC3iGJY+qKNSvRBesi2zmKYRDnsYqzM2yQygyP2SZzEvSik/yF9p1DyG3hMEVWrauhaSx
VPipRll9KTFdU/DDQc3nZmJVn0Qk/NXIkCpA8a9zOfOaD3GL4yoQsNI4/H0pOTYF1FcfRwoJAzuG
qTujL0H2A4ciHKMDYK08TeWDAH+iLHOuoc8s+SZeJ2dK6iBW5McDEL9zSfI0pNpssEJyGcj07gJ0
vQz+6uSPaYtLOy5QGpuiykF+85tfxDgmozO7YdgfgKFuP6Cx81dFZN5Gg/kG7QGyFKPwxf74TKzh
DDQAS+BWr/j3+pH7JByHpIIZoq0hJxmpzriDa9RRPyPoTyZ3RJLn8lW3kTLKDFhUY1NC/noILoXj
7XJ1V9NAVlK5wIrhH9JWU0mylx4rKAgX73pS9wiZRqgZWxZdQRQNJtD8ZsM3BAtGI3z+9uhX+Zpw
2SG+zHMPQJQ9iEHMk1tl6SWao/OvCVb5d8MISUDFR8bwKtJGrZczZ7/7O8oviUBzQSIt7WwaBwVU
0VnGa4xFG3hSSIe4x3DvteFg5nYbwdBlPTSQa+8QB97FuM0w1bxxIJreCtU2R6w4DX8b/bAvz8mt
VtTwJAoMW484/yjttToh2GKrWobSFaDzVQoZfTMBk/tn46WX34uHgGTP31V9ea+mpRSaaW39DzAl
8WH7yJECVJ4mS3XCJtDleqg+6Co8Bl5PVfU9fEkiTVXA8HdY9df7HQGsjdPEQst21OwSPJ70XHEF
Fg8iPF8E+qcswf2s3dfDNzb2DeCpv2psVAbCGqc3IkWaKk10vJT9bcziMEmEcCu/DBoFQC4mhVYJ
8qZPVwNuU5w4fXHnMtD2EWR1kVohv5vUCQE+1xwLAQ+Ne3bSrHp4ReNKQYKTgJ6Ia9jz/LnoKiUU
yl1AbId/tUklN6yahhU9sPWdOI5idV4pwvCVntY7gPvMWjgFz+/2kBp+5j8AwucBve+BmFNw2adz
ofNADkPNzW3FfH44RyIutiz4nZSaWqobH+ZKJ+Oqq+AfKQKfcnuprZUO7fq9WSJ6ZC2UjWpVWRpn
JHWj4HYdq7RZAM+cbp3zP0GSrhR4eOPKO3CJwpkZbeB21vGHZ6qd7c3d0E2U7EJD+dAPxuAqizli
2Yqy4GT5Rnl2+Iva3FgowqCfH3IgJYyev9Z7TZm0zV5VV1eW3KAXTIybNB0/vF2gIiNu0XPzs5Yv
xKxrRjdxHoXZ80anFVgEAvaB7wIGBzZRzjPj+Bn/uHrBOGox8gJy5P/NfTR6I7i4sS9n+m5WxP5+
HaK/Bw8sL+khB2E8jTGbGyPdagoUN+Cd/Ivo79UfTfM/2ZjutUNR9VYp10ioAabwK6P2WyfXaIGp
cEGeUW/LShW8rdshFu20YfuJ8843Nfjoiq+retH0eMBCJazfNBfd3Eaqh9qqWMQvKv3EbSMxBc3K
ebZk3g3/g6mHu7m5ljXMWdr5Jbr9lPWHbN6wik/kmShgOs8oVjLYTADDjgxm7zJS1qDz3q0VCDSh
biF4mzomGgwXhdFbxh+7sUWIerxhBaRKIpfYNk2zL95ieKccnORut7IjEoa/SbgF1l67Nh1G90bG
FBaU7pdKAPDAONtQJtW7YxJcJk/41DaGeOpLqLAGPIjup8V4BCISoOfUjKqineR0BuxwMHe21ta9
NIRbjGB2XEP2wzuX14KGdYTiHKiQZrtIGFuy9XtEeY8hQNMJh058MCFWE/rGLhjcGeKYHcLN+9F4
qk6IKy7NnfYVjmL0V+raqWYdHin53Q8Rh5sU9t1qJX0V/Pzx/Vkte6M5HuSlGHu/AnBTkYs1kmFc
VRIGOT019RGKd9aKdKcH0Hu74aznmKA4LcTEmHYqOCcXx+JGoHyiFa8scLorVGZGwckba3ylRnus
qEehVBSm1CBC002PntwAMLudF/K07yhlaaNB8L6fw7oCHB1VOy+a1/AbvbEQc3f7DfLgWptoanKS
Cj920pLEbtn2cAyDBo173vbj4y1yLrnrS25bACOV0pq+L+mNRnrJEjJN3UdJixRBslOLCqewUmXZ
q7pp46hxlcpZ8s0iDqaTZEQ7qpWdfWLrpFWf/cIrNgCOozWdgBDQ00WbpG7ixt7dWrBDHDiNHpex
xI/hXhSixML8ChE5n8EdZXbkzVJRkG+gez9jn1iu1HmomFPMWDiPeONv8eDzRLuAwtuYh9AmZLqF
s7aeO9rOvcXKxBiwkJmR9qEdPxoxPXOcJgTZ+zDXCCoSkqabi6AoDpOqv4A+OIaNcMlRJD6lhmYf
8GP8ABlrZBd1c5HnykgRUyD4baSqkYZ2/RFBNkXaEMeslWOHOoK6OzYs0FSFYiYEcOKvMlgM3WqZ
m434D6RH43F6D8WzkFWleuzOYVlG501xGHchhVsNdhdpeHnF3OpLktsMgeFhZ3W5F++784ZfsXp2
ksPtjHmuQJWgHN51nYxR9wMexYdj0Rjau7vUNOmSpoEpaJrn8nQcowPK0oT4OkCQq1JO3TsFmf8q
f2wX2J5ElvW2mxJvKJrR/3PVvQSn5PLybvroAvhjZ66fuq/LHSHSBTV9ZTXgu6L65Qc/MgFQmyUx
QhM5nOahcM2H6gRsSszVKBF06/g9ao6VA26DLdXyBOnvDgiBJ6m7c+7/hQPLQKVLekC//HvJ5+L0
qDnhuS35kxzvZTHx6fy8yzfUdISrPdzJtS3dkYEEYp8mau4XMu2obHdN0Izf+lMO5zf2xrj/IKj0
vJAV41E7dca8sw+iYrGxyf3S4eawUu614ocOz96KJp0lJAJvuIWDi8O4IaupOpZEdIuw6gb4nPYi
DXu5qIqF2gRcYzkq2hWEOwPhckDE7ZNeU052KUMhMu+BFcvDp8QFSdQygh44feaypqzONDPGn18E
do2SDRXzz7Xdc8ueCVQFXcAwh042wNLpUse+6vN6Q0e3WhvjzmdesGO5oo/7DlfjSaycsHvVy9BG
N1pxDA4Ih1ME4AJp4ijBMFzCdGL3r9lTKRWgU0qHqlapjWIx4GVz1sV9TYU7cTJ8o7I3g7uLq/Ou
tWQNVaM5u89d5vpPLRz8VNPpKvvUga5iiMmI8KYhT+/p0T6QWyvY5bVQkGiQzTs8FaGyReUA4187
z0Df6ZPSGtRcOdHRGAVcq8Nvf+ORCqqE7WuDgrZvwsYi/4RJ4YVloN+nEC5b0e9NY2nyLY3E/zXS
YNp9PD2UjfB7DsGROLUoWsCIfYb+XNbRWK9o/u5UhHqusPm10hI+76pQmWbjyKqPdr+NnZj8J2n4
aamdDsMO6ZrHLgGawSeFYM3/+I6gkSMGsHQcfifSRys5Y9ZEqYi3wvVl2pVFCPxCIsM1tme5/Pqi
ZxUdpo/kugmpq7TjwLQsgXAFK05/aguSNqmgZMFOg7r0LXwNrHt5HA4oHG2jobo+jfDZE8PNY/0p
hEVRzo9bYRzfP5EAtpwUjVhrIjexm8VwiHP6aOe1oNY2OruQSP0isQyf1c+t0ER8hroEnfkzx6fr
GgMxSqmMcJJaowjNUJ4Bwopk7Oj8ICs/69nX6OTudc0x9dAMC9hQdaQ5Fw4QZAr4WqVs0Idbb23a
a+VriLiFoo0M9v65Y1WEzhqNCZz2kZhyrTVK3ONAJVVOpaKWkdEG5rYEDjKgImDnp+P5vYLU7l8X
v/tHCd4Sq5cO4PF6GwHSEIsAaLBcAI6rmz9GYcRhYr5+U8eJYmmUJlrVHzAqt0J908Z5pekBQPtu
9AzJjHhcUQdjtE8BeJjboZu+RgiaKtFUJYXjPCLM0v6xp+DIfnqZTI2T458UheCztWGXVu+kwKS7
6r844HpX2CgOrQY9Bq+j7SLUSx4+dHiboZMI9mI3oas0LVuIPtTSSVCafhjv6O8IHT4Vj/a2tSEL
WSgugiAnABhlxRWzBr5rRuvKSG4tnlUN8ILIFIVEpvHVdkywjSommGHLWKSHOZIQ4SISv8eDoG6w
ay9K3eaBOQ2PT8AWDjD+ggiSiFP2XwEgA07+/5ju1WQk75VBQaPoGld/5w8+9K6/75axGCRN+b6n
d+34AxlcZx4IsSuhY1TuclaitqWwztLbf88UVxm+SU4gXi9vYUo/G/n+900S6P0HEVu2bb0r8LU5
UmFaujKJlIgsBEWq8Wg532k63AIbssC6pYQtzUfNplIvPJSfdAhZTLN3xAVqW1yX/j//mRo3DI6n
3f+bj2gZ7wMCzh9vtb2T9UxWNSqP8atreCkr3mOYwioIyuuJ69QDoc/hISCeqmv4OaE8nGmei0BH
votvh6gghvcwuyiL/rbqzzXfCK/WRc4pVNXbj/FSLo7F0S3NpFSF2A4nGff/7KRYnkMKB8YnbAir
SknM5BbhIOtFSLm2vTLRQe/OO/MSCoSicGOKcfXWU3ctFP6BRsLJMe3h/IheMEPvfIrrwEeweHN4
WTwH+LLwPGZ8zpJ7jc6t6lJ5SYgdqbzvykUHybnXMt3y4vZCaPI2K8UPYBlQeE7TzEtsu3rj1MuN
ivg3wgcgWfLY8mEb/ifWe77qoZSue/++GxfMKu5XAb2I/qM2HjEfPmZAnTXJyxcu2d93A9rfCi/5
ZPt9X0c2ElsB4CKlb0XzqM9zWyUre1wJrtG1GXp1SvdqL3WvxVy9PTGCTn1Nb/55KcJUvYCTr0Rm
qA3WT/C/aEUBz6N/XcnRgtu7f8VSrceQWhWrxx5jVlERcHhZWq1FKxGzLCE4A0AEkIouRUZe/unC
UJTEWUML1I3hsv/XeFoJ3ace72nUwup/CsHCh8e58RXUjRrVeOYk6FV6i7EUma1GV1W0zKYsPfHN
IGbx/1SKNMngNe5zQx1GuKng0bVvfTfs8j2cBLUth4i5lV+E0R26t0459n78HQZYH5p2qlCGyHtI
C+VEQAftOaV4uUUCAvdyb1dP1o49m7EyWyd2fhlO40BVc3KyR3jqu7BHZUxSV+hlMI3jezS9HqFe
mhA/lm3BYDkbTN+Ov8y2WRO6xkSmsiHqcDmoCdEjVI8uqxW+BVpXFO2Me0+GSZwHZm5EB0+6x8hs
7FPmvrcjd5hVPFea909C1Kh281ScJSi22SIJBjy/ardQ1dY0Tz6RNCexo4WPJe/V1nKxxJ1lNPMs
IE5GXG8m/96LxzpoFblL29hyGzuANU2wvOAJsych+R6FipwWMBqpp+3wvwkv+d3fUEXhCGQ9QRz6
/k+Bwo3HypL219G6hvostA8ta7JSdetOWg7ndqau72PA4xZJ+VAhCJraVwX3lwkLhPI1cxOYfmz3
rc7p8ajy/kDcUMob1CHgXBO/3bHLp2pOYOFBZVMYuhdt/3sZx0jY7qcKDkOiyQNciXeYj6un82uf
a/YXVQkKrQ/snbMXfwtLb+dTkKsBxxw4fODKMXiITuIc0XBTDq6gk9jxESO5mJJGpv+VydbxHKcI
F+phaFWv/oewno0K9TlyaSD2LytyX7+Ct6j+BVEO5jRKu7PRk1vrQelMd4bB1ohI7Bkib412ALxO
tVEvg4QvQ5PMXzwwVT3kCYSJ8nrR/Dkv85kXFFT1uH6ULKu7NH3mW2r0NEaeA1AVTbGXOUY2too7
PluYc5aMwYJzA+FoUMVbi5kYKiPF6qIyUW2KUhn3/SxONKunG3sJhmKbShPA6hHEH7sic0etS2Fd
/1e0r4SoyTX4MIGk6GrRv9aTk+1EYSag54zsgzUYT8ckCVfKDd2uoout+xE9tL0sVFlWTFJiYUas
QcWewFFwdtNMnxDPtpANng2zAEGvNoObhP8qluVEAIW97NVVA6LGzRlRXXxUeUvYnahGODzQhryL
aHW/m0g9TjzToJRK9m2nD2rToFg1gUjCb5rxlOIZsVle1i5alRnZ7gDUuPx9BvcXDIxvQu+4/WA/
7XKIDMj8nK11yzyAOOJ2XQl262NkdeV+NfpezeJ8KmqplDR7+vBj/1g/ZyaAxSab3yMJ7ki0XG8p
j4RhLVb08fVxg4D1+xF2iRt+Qoiz+gWlcAWfEbO9bTPaMBlTsER1D5HQAasICXK1S8CdFfD4Ewhy
Nc2s09gYJ3mUeEUCunVKpQavDfXaa3f/AZB9WMxyQ/09rd3aSHVZ8bj9pt/2rRogzt6QPjblQJRB
R8TVzZ9ChWNhGXQvh2SfrwFOgx9Qgk33A5/J3S8RIALBH/vk1YF62MdgLShJ8G5XJTI0pPdMXu+0
hfdN1ESqnmZofSHU3E6EYOIKFXmutLbCgCaUlqfRoS4yuWCrHau6LMVhG7DhzFp0cfTDiQLzZWaI
oEdbQ7yz061E4HMbwsR3NS0ibYXkM4v4X99Pg6AR7lrsXLNpci7d/scZD1eOVxAzqHMh7eZHOUNm
b4A7fUBJIrdGPYyTzX3EQNZeZjb8hyCF4LrbKuJA3rBwu0AlmaGxCPrnrJZibThS7FyHWFQnmsyj
MrCNuGPBej0fEbacjJpTlXrM9cKmDShmwKS7gIW300ZApy+TGXxQhsBjBorGLDX/WWN4yR/DayZ1
u2R7zMoMhvATyzg7G3RhRCOR+c6OcQZwL5xKQZWkR6VrANKnCJMU+88OZrn4bw/kirSxIGC5d8R2
pJ5ItJ6ADaoGtbd2mc3XQsurBnKRUtOuUa226Z12+q+iF0q1R6Bcg9rG5nqNqs2m1xfJY42S10pU
m/cx0n+6QGfd0Z10+Zzxd8FTj08GpZ/dxx2iwek48XsMlo4cFhm/oMx3dvtZTea9iSXcgruRTDGJ
msNf4K5b2Jkov/ZpjSDg/cQ/wAig807cC6siRtwq9GHEmkzIMLvP048GJI0h13G6vxpqXiuA2+gC
WFqIEYp4MTO3a8K8BnFTvnL3aP+gAIDXY1eUxULm60Ww7dBEGz5JRtzuBcH3YvfqadrhdyC9W3YR
oLMWy24T/+Qe8mCBkhmJ4k372a8yftG+2HOq1cRivG7F6ZPbot6ZO84jwbQYA1aYOOpzjghTtpDk
S71Jv0NSxKT+F7YpQvJiRpuYnE/5hkuQoXycNtLUpu5+O4lV1elABrnNj86jVdjloubZCPAwTct5
H0ppwZ4iAOeVL/XI7khEfSHku6+5llxq0wI2JdNYGnq2Slyoggb1C4tSbtWpbHH24nDuosJUdjpe
KtUhRLuRSyN4SRo5Iq2IPQ7qzMyXT0n1evTDeuKBsxdtQC0yUud8uRykrRMolUtA9xcqz0QiRKP8
GspQs6CS9u4uVqYs6dq1QeVWVsDc38gTNlYCLvYQMnxoaWNdBRvw7dus0sKhzbhK+GX6RJKC0kLj
QLKvB/QqnRioISi0RqR6zuaiJZKmayvffFfF5sXf2dUKq7D8lk9m8yq4gUtw4T2fg3NhPI4Ofi0Y
zIkXBPXFcR0eJDbhQJz1V6wYFgR2zLL6gGs2TQzLVMfU6Lmil37E1OJKQtujG6HSOJqk9bHdOjcQ
qm/CC2BfSRLV8bVjbPGmYcmJsWhUS4pAWzCIy+uDCPAPbUhUl4Vm2EDx8T2mMbfMI3C1i23UA9vv
zv5hC7rC9bFHa6Yi0xESHmpKp+h06JkdBvhdyXTBfDMrXQUndjtpIZLi2WesLUe34kHZO8pBfb3r
FGq8+RGPaoReesMO5FxLeDOTymTPtVmZmGTHwpdeKXJp6dIAYcmX5bvo3ylO5NUEwqrEI5eVGiGf
41je8r08LaotNCwSnsB1GxLeW1xjLxsaiI2MpvZovhfdvaPBMwegae8JxcwD9QoZ3sciHM3YALz2
7pZ0Rq8Z3s0zqEA0sB5fI/FDBl+vMaWPvOhSFvBUciIRA6wNLPKatlN6A+PFdL8bWjyKUeIHjHby
MES2ZV2LJ+q9v29kjexgsb/ibnxVPabJw9vWJcrv6WliaZyTmW+/gOV9qOgFdcHalRBn7oLep//w
BQXGYy78op3u7TpF5k/znl5r6CCtdashaxWMcKjaRKW/kSbL1uKMDwWSZZIlHZxr59sFpcq2Ci+M
qGaJjK8X/10Q4Q+JALJBW23O1zPByIyaE8CWV/WG80kbzJuwDIFAOP9V+fFYaFjkbxZb8JW8vs00
72laJw+WtiG7YfxmWz09VpK1+C4dSSVHHMAs39B+KmvlMgL6b60Pc05XoThYVoR4cVSTgldTs2ME
5C7czQaN6dBZ6Ndvpdd7hsyFi2Pw6RxXm/U9rN4Ht+MmM/PP7dvOcWc3rL4vATKe3prC5NPXyoNU
Y9+6FT0yyg7WqKi6NRs7icaFsXDSR0xxRXNqV3es4Gt7z7rpusJGs3ehNvQ5ae7s3O0CzWQcOMYO
kAMeScwuKoulT1k0d0/ZhDX8UZowpoLafSpdqJWsLrWD5pHFCd2m6udEAxi0nQsOzm8CoghUl6Ty
g66QhIRBySMNoEUkgPJ1ZYDMJq9Dr08XrMu8TV5xBJxqP1fSqx3MmeE0R2dKddWPROOmCbe33DJl
sz4WkUVdfZUJaMwbDh+xlq3h00+iuFSbn+5twwCzLwlxg9hxY5KLEuDSr5DRvEAOyYjPqX/Dh5Gy
EGQfths5rjZyygwVI23T/0q4M/XdU4kjxFGSHxH5dV+2+slOs1slkcQwUasMBHBlBfC9H5KGtP64
rKSUkmSDOu+A/CMjfbXcWGpFy3eXHjX0JZiQcKivM/WRa5fw60O2pNTEF77e0tF9Qe1c2Z0VQV6x
D/YB5TIm8iEHZKZEY2dAfFTg1L2Z0xS58gfmEU14qfCVi+n1yC694nqW+2582BswBmrNJ7ko/yNc
JM/KW1A1wa9P7Atk/8acK1hYlyzLzhNkD2l4C10QLuGA/eOci1SkOOhiQUgkGPoCv7oQIOeyzmAH
nFRMzejQEbx6IkhGL93dr8Br1uTd9gqk0rAQ1PTWrccLTwTRWY0xzS60pOnzxDImUpIldfP11BeS
QYEr9mOI//OeZnFOvVkdxQQHcMmKVdgm7YxbliyRtB4bhr1e03zcczgFOsenyVbVBiElgVpAxlVE
hkCGTGSTWlcR/yIJ3v7knpz/4UtFOH4UQuu/CDLeP+2uD9OnpDp1Dz2ZeT1kw/AFMxXXaVP0x0vf
ljbJO4TFzfGdk+/tJp5jZ8FMbMRXR8RZUHaj9oCFGSnT/kCrqMm50qcoideryuw9yo616moS45lQ
834s84q/AQObOf3+TOBFTaoVZUDYQ6AJybNfZ1LyPA9beJWriD9IX7hUa8Shx0zZivIwXR7JDzdQ
K5nV+B4W6eMPfzKVQJwF+K2XauoDgEPvNX1qZfQ0fDC4ZYXFLiJJNvGQ3hw7sRfwcxwKHji6Wmg8
GVaafjIqG9pTsJfukq79gPqATsNRhM+/QcPssJQ79oDaomc6FuaM2cvufsy77HrYfLGY2iHRo7nx
HNtalTpfnRhdIARkceovW2yEBCFk+oB2S1CPNvmxY9qPQn8dJYGcU0OW5GExLNi5I0b0MQHk4nm+
e/3JbS8UL1Cy0oZhNZJrTu3YRfgESY0/Nbqa1wXef98sPD+DZ3UcmS5OMTBl/SmlwnXWm+n7Q7vc
yR1T8LdL3a1juL8LKhtUxPMYJiWoX6ZBQHVvQ8RQm9WIFKZNYeiTJ6bRMBi5rI57jrw2jHEggYgy
+mobqcMIZuhgLrmXLBH/JXU8vsbV1bY6DN1K30SWIv6qlNcMdeeJj/u9OKTSfIWDc7Y/DRsUbnkb
o9BDTGOwqoj4HM4wZTLoiweU5QWV/5PjFXNCTrBZhfdF0jS5CBZ4nKRjMATQSg0VRCI1jZJw0sbP
ae7tVKK6ig+oWcEatvrcVlH5g/itrJGGNcQ1VmDXsrtqMLr3FYlysf4pmj4AH2TgAM3CiPJjQTWc
4ktaUQv6upph+ZHoAqKjNvnzVHWQG3BYIlGe6tGUyJ0dOXzTYk10IQ3LhMokhSSwZS8DvyIQkZfU
ci9t8uu1U/yagX+anlaBWZePgojfKAYgKqpkKKpopf0lHUedXxZGoQvc/K8z3JjnXHBeZPEIASl0
V1QpNeqFPUVoMJkbr/30vdqkaFLFca9DbYYvYTmPdwNiom7uLcAApWjQSKWkm5HWMdsyCmdPxUmf
iXkNVt2wvtNBwzhfmDmHlWcvJ41aWt2UorftIae5DNLBYYD8wtkT5LLsBDM4aJYMCVZImFonJeVU
jXi8SGLMMMmx8brboCZ1j/YgevP+BjgxHsTvgAi294fvOkYcEfQ/UM0Mo0eiyNU1ed0Db/Iq7Wtf
r+C8f1JOE8gbUSGYYGo7utsqc9Oc9Wet/glKsdn6o7eiIJ1PKu82N8tozxMm4TLc1JpE1xsFiEhc
iJ0d5hCHJK+jvYC+NNFHeIf9J6e+UUaM3yVpvhkVML3K83hvGN64wf9tSMG/2I285e9ahbnl3POg
+UQ2D87ZfDTpI6tFynj8bXgPKtChdQ7+fpE3ggE9wwkIJhdZO/FL8fEjWJII0xFwExdrQTxlWUVX
OE+wvTlUKECUJyZkUqsy1f8/+02entka6D+SmlOCqDP65zFsGnEcjcdT9sBFRwz6da8nuIG/CCYn
SCiumJ2EhdgmBakaGIXGXg/G+mvDcqmqbIM89Z5ilefAWuZFvKzkxZp0+NWcxu5V61qk3AzZWE+S
x/r0GJKzhBAI2u3PLf4qQlkGvluxDmGsq+JFHKcaOHMBDxWZZdzSRQJJj9bSUE3ajH8KF8xZw8xI
ANeuI4ICHjcHhsSXyzqh1H1kil05uHUO8U6shIHJ2n6uXNgzHtkJZOyAKlHuOdA1fn9U9EUaVr1x
SuVsXgqtoROHXIjaCGKpBvLpaNDN0WAzMgtxTtTpisw9B7giApjtAXBwaZlg7K+klieGmz9FAMow
6VajKyu5c9wjf4EgF7ndqbQXKC4v8RjnjTWfIH1/4uFYz4/5UxnksPtYDv1VYNs53hcnlvXZTcDE
UTpkj8nMX0nniIHvU0FkGrw1THu6yKxIFkuZzi0zSvHfrejMvxcHQctzBHqaRUdq9hMkjI2eq3RX
WBrEgzCNlOwi8lrDcdcG1E2u2GF1YYHFgLR7RP1IKgfTGODXk2rxs1eukSNqQ8VTDmSO6tkn6l+1
ZLS4gpCsmYSmjMnJgi9TqUMAmeOUt3aAQAcNsZjI3N/lHlbggAjDtucFPo7+f6WU+LDEHeA5JpaI
AzVwomw95QKRAmniCaYn17qHapFdQgwQEUTtex5MNbZrIk/7J4dnN8vlhsotPdT2bt90+3TeoFul
9oY2nLR3a9PBtvoCQxUkhS86S7ShPbJqW2tJ8QP3vLN40Z6r3NCOfivLmwraQHHZslOn6e96D31M
YttgVIbhhO0jjXRUaS/DEex2o31Yiv34AT2BMzMEJDmH2q1kknO2h2m4tahpughxrxIFMDbQfx5w
Zf/BGjp+4QFgPz5LBiEA/09TE+gIiQOxArvfblmqzJP9jX1oPT5u/ztBhhttA1oSCjBlG63Hnpio
oKys64wf383B2ufNQiknnbUlEqioCC61jWyF6s6MSmLBC9POssL/5S7iuh9Gngy8ImCQltL0r6aG
pC4Ei5oQHh90pdDonqql7fchKaPMR8wjyiSbf2YwI5V9Au0LF1jrfPkpZvh33kuUI7n7gnw1u/Yn
Nz9301AAmcd0ae6oIq8kdJ45DrTxpigRwo1Lqwld+PIPquzYjZtpmPAEG+UupA2dRVtHsZuU7bYi
8Bpfqkj8tfAIsn46jVFX/FUJZuP4pTwXdXKoo5Z5KRz0lglyOcDdDnyaGSIoCWvboMKL7OABqGib
HgyWEjf0cKC/5KzVl2Ci186pSZisKBGcYYqnbXuWuCVm3lOhyUut19oc53Vo/ALWO5HDaamU5w98
molXqFPE1sGYCnF+tEGTLUcIKr/wI1Jaacgw8PaJQfM8MOIeP+VOeuDg9FuEgEtAbd1GUzko9n3j
akK1x9HDJaZeX63lfQiecTOJSz/UVSIZONdtFhuwUL7gyvfwHsvWT0i+lquik9OL1Av9kBIUYpj5
h9x0CnF3D0G4FKOhUMpfK/eODvFv2GN5mR54BGehaV/keWt1j/8xMvkHTmRump9Wa0D3HnDi11PF
cGdlMUq8VEFjysesAjG+5JqnvRd1Y+ZHKrua4rIEIYQkMhkUf3GO+s5bIqQEAuF+Wa7h1aiuTGjO
50/q9PhErKi8b/eZO1jxEIY1tU+dX8TRPoyYN6JArUkLJpVa0EI5UuAt34uc1B7ahFxaQgZv1tnb
daOR2r6ErytrE2RJOX2YnGOoAXTvYFWrdV2e8aza9F2CSE5c8VKaWXZ4vSG6stk5M58SQ45K3c43
W4KhIkTArtv5HlQebWuUZzReerJ/s59BF3w8SU8Bz9UDoixH/yxt8FQ+1sdX4bdRVhyfx1/3ND42
iC3hPxjSGd9Nmo3jrUpxu9qZIbJ0SEpeQV+Jkh6OOfJBGtepz3lDmqASMJAppoxtf23lqZNyvGQi
lPzexn8Q/m+9nBeCojDqOWQDaxTZOUKQItNoiCLzcV77NvxLQIf/SFE0ExJxkud++SfwMgmQVufx
LW88L/EhkDRhkSD64uTAQWCgeM5wICHYiIHZdGoH50e5wjBVVwVs5ZW2/YKBjj+SjCHUFjj9tn8I
ocDe9l6uHCfVr8ChLCwjW9P5DvW4leqVWI9EH4Cy6fJH2PFvo8UVNLRo4pwYiJz96rZk8knTvp6U
AvpiWWvtXLFVykpLwJPYWpzguNVj+e/nQPyfG/mHrjmxrSPCvyI9SuOOKLHY9PeWQbXF6pyUYQ3p
jYwWZfGsrMyEiV6gFE+r17j79RlmTq04bZL63MuDtpYVPvxPjY4E6vixlQ2wu2576qGb0b5fw38A
lbJWK50JDajeeCnms+F9zPtKo4BKZIiMiBZ9DnjZvfPKIds7g9eHKw5Q3k1AGSf95433EjVQKPRB
SdNVhRF7+TGqyqHp5y5tisCNkjPbiVagl8GfoLXGumY2PSgYKPlET4WotRBhqQKrBXiSSTNZsMYq
1icw4s1MECuFnaGgqZaTRoPM9+Nx7vhSiO27mp1Cfkm0inNoYTDfgAhAlTGAdt8XgZWbel3LIUgV
cv94QKw7TRInW5FnoOOnzRTRU1m6pqLjPWhCl+u0d0Q0ughS8c6TBj7Eexbt/OCdBNmLfgu/rE03
9wJIHrVLGvSmG5hxsToI5U3n42zp4z2xW87iFN7YQt0Hp3WkwxxR0jOs22gU6P5FFeffWHYY0p+F
XT1x3H1oim65+vqpQIQeCCXE6cFVGUZ37/X0czfHpyt6mtu92we8/nSDJATJyyot6Gng7ihaj8Qe
IKc75H95vpmEpiDEH9FR4Y/pYVm4veu1thBbb12yr+qHKOnUdbauv+K+xUsTHVDHmEr9lP4owTfW
op1JSkbfWP7eNDrzKzkGTgNu9UsP/gbSG/Kh/5yzNfKOxRmrRZf+Za8CR8Teqhs7jrRpNy3xs5Vw
fnHqLDAkudjv522ytDy/Ts37umTHz4Qf5+z9PEqK1UvT5uHHaQGFbYlwRAkqRTPffUtzQh1L3uh/
fnSamrWFFz20mmcJdRVMyFbu+M3NU2flhp8OxNgdF7gIl95Ou8WylhRKNf8vuN4axrZqC7MoN16f
KZziGbbJF2/MxIzm1X69/URokEOReltuDcGHp34UTkrb7TY7yobDlCyOuUvrzJEm+7cVvKiZBsU3
QFh/BlxPwWdRtRMlbJjKq6/b/9ge09OnDeipBLYfMdC8h2e5gHID4c+Bs4qCtQV/1+7LveGgSFlU
sSAoJBnjB5NDKOZjDkmRu6/UU+yXYw35A6E2n6Gufc9fHa2Gty/JhRtobM1kbu7qHjZ9BqthMVoK
ewh0KhLf8vJJmZHFo+FlF/74+HIQY3Yg8WWoX4Mx/REZo2iH1SZAtJQRF7brfflo8AJ6xX/egHpT
TQuzm5F7h1+z0bAcvp7Js32hFRYsaZUZ4pVnvWMfpvCPnUBxyGnM2j2khid1WZv4o8ltt+Si1w42
hFPx1q9/nIxf0yEsMBlLAnwToZnI7JtJv2flLNGKzEL3w1CZObbAO/yTuJqCXVtH3O8ogWTAZ/Hh
MyANwZL66dfw9ClWscw4o7jtZwGU/sK2gHGtVjeD2goeZ8/W/vzlhhqPTYtnttd/nInrdcxZsqin
LtIzpXRgcO1bLBnMuncI264oXgepI6V1oklut+xflV/BBUxlgguNjmTy4mL2cfPjQjbeNO7ZxEWF
Yc6foOrhw+oKIWXcshGb+L9JRXa4kgdhHBVDbrEvaBX5RAzVE7iaodokUWOy9LXgWBuFMqzzSD0o
B2GIcFi343XXZFGPqFCGP2OJUhhYSIuBV5PUQeqphiHZT+FDyMjKwLW69HJ0H0UlnsRxpDuqPtKa
hL9xu6iS4+GIKLXR3ML4zjvuTG95l6D5n5pkuLjjAUijOMV+K7uRr6EAlYq3DieHcJDdArEJmFW5
b0lbotnmoXHokA75Jnq7XF4kBSMSH8/R67Ob2oFsjQKjIt/yB/Ltz5xNqcl7K+K+CeFmwFsItTzJ
8EOvMCCEd1l92cF0dnMTmQUT1y89Hq5MJJPzgFkyPgfTlZkRKigABgK0oxeUY9FVw4bJJ76k37A5
5+otjVgLKgSLLtY/2n6Nyfb/8wGcJD0u9l7afdaRZZrgo7lh6fBPj3FWGGV4iUJEBWR052jPH0jr
MEM7vNDNCDTX5a6S/x1gxsB+mHZ1yYYgsthlOYQZ46ClyQ6L1wRz2RDRynjMqC5hee2NIdN0XUEm
2pBkGisiKAH2PZ3m42r8KsHKaawbE+oS7ljtwZP3GYbpZ9/A38blS8x0Tz3WC+P235pBEh3w/QGY
i1KrewEjaGvDIk/cEfXL68f0149ovVejzW99kms32Su/eYDOxFo3QxdB1AtOk0jp4VZPudj81Zoc
ImUWCJjNrjksNBsOJhP6iTbPC8f5xT3KIXWqLtXJAllk7s1kqJ1KSQ7bYaQrmg1a0ZJYQZImgzP1
M3JeuUKSIS8TQvghY7itTxUKCdJXLS4cFo+RcEN7fahLhEatu4htPn5+TzykDHRr34D2XGDYqzrE
UD0QnrmYoNnvFnFrZB7mWuBqsIOLBuSFj3Nax87p78BcBXfiS6d5Ls9sJdbaE8Tg4VQBPn1blycu
tjttqqFT79MPj2mRCr1kDkOwM7aRTOX4Gszhe3VY46jmTrNc0vuXFyogMRyA/rwY/bk4UctU0t4Y
RIDtRWfHaIdzSPmfDPbJpYsFTFluBv3+axLEL478Pi3XTxkpcM9wV4bN1/StJpqnnFjdommMREos
MmC/Oeh+WuQC5qDK/XlzMnYi4szfZgdl5D5u9jTOTMJOmuUlKETirc2JN+y1qojcLdw45FDYsNEK
ZjmSy+Kw60LayU4jPdlFuUPlcLc605T81NIF3XVDKqeMwl/FCmtlWKSVIHB6NTHxXrA4NSf9WLD6
Ei6HihfXs3PcsRVpG0lMvJuU/zXbsBnFwssQ6wkg5tJ+kPGlobdBoGhd289a14KqO1cKNoeaueSh
Mb9Vp3bfQJshvh8ucqCA8q3IH76ZH3Q/Nhmkhxjh6jN71gEphWUubF8IHo/5r8ghsY3v6xOUSCZN
F6XQXln9FBZ4osUx0VtJMhpnKHd4iXCwwzK9CBWWvkhdlIzfS1+xMJDStOxrH2tJXUd6ktqWsIYj
W0ZcX54nP5Pa9xbTVRhowMrjUkbl11CaY1pwtbtrBxYZzA6fEly5hMKBETH9CGGKQQG6h0HydbUR
2q3YeCZ/BOYE5JCz9pTDkvKs6zYjqFB1+p4NMBxWOl/NYmQcFQF2KAWGTiEnxtuSP2NL6DXwGJXk
VjjRbyfzNVkqVNBx9rELQBwHqFvzZADSQBJ0DEkfdXgtiDEDGGNOBjICz39RXK+pTyceqyxPRVue
AhIJq1odW9Rqp5FWlrJmvo1D4S6PP/ED/l58O3BBo0S1pE1f2z9MTWy+7rIe9MUSgQyDdWh5SXwu
IiH73W47cRSyb9xyi2ZpNmZmBWEaqE8+Iq4e8oJTrTy4wYx5buAS4INyXynmCYcAEUe9R3PVGiRx
ee6jxCjGAMrILManCylee/N8nFW5STzjT0oY/cCSiOr2lob1dlyPwRKVmW6m2SH3CuQ4hDeBrBlm
rLWyow1ozGcn8n8EC8UIMJ5dkmheRvf2q5QOCqtnkbVdP28bOTqS0sTd78t6DrOnZHGZK53tpZRG
xj7vy2+MYTRBthNELvCBbJJwWn3a9i6QJVvLx+KOworKEeXKjua7UGVMYB6DOS6g1tQw58AG9CeM
S/U6qL/ebMfaHjf3HDXT0heDyDB+4wyYKxmv488o/Z2XBWtkaIvZeLiVFpYFwpLR/9AoeDP6oIV6
xaYXIz3vWajLZxtygmRVGg7VCrl+5LtZyyOUF7gcumg+aF31p6KdQEaAx3OrKFtIbA+hWF/wRVYT
nEPxJt198+n5FwWo7Th6UVRWvc7jz93pzN8FaEJqvz5BRdooOCqkDyMunp/6vC/BkBAbIV8TxFje
d0ueAwHNQ6jQXhCRlIvXCC60FJSLSUZx7vCBRdqiZ4vSyI9t2IhmyPPieKwMZpqoi0t0ipEKycdZ
c4eTqM0byCVIw6tJfYR7IR912w870ygCM19hL9UIn4T49YgqYuVzhbEjY1b4KBhilzQJCjEQCmkh
ukonLTw+WAj9keEJDFh59j8n/mkkZLGroAFDCCtef3hQ78+nR9oM9sZfrrCoWblbrgnc0G+CSKpO
BStd8R2Mc9qiPeNUXDMN7XWQ8EQlfrS0UwY6ShNHOi+46+1xSPPL9joRrfh7Puj71oNolBZkYvOQ
9Fo0XuqOlcbRyfRFyNS6AI8TAuWgpw7GKyGdN+kfdz9YTW4L4N7Ycc/RGh3yo9sLkRav1f9zhs3K
RTtxbFK4vxl7N6R2UQtAYmd3/V2D4znhsNPU0U/9E0NRhkszHfGjXL9r3lPxbDVY4t4dvnuTkfKi
Pkjqk/zxvta+AbWQ/VMTBBUck6sFdaNgiwxnF6qh1tHZmhR4ISzOVARnMH+9Di3P2gXO4hwkmaZ4
/DNxw4nlTt0pD640UdQGjzxrMwRves2OJUTXVeLeCP3t48NgoSQepMoelfE3v4Mr02kcp/yzjz70
hLVQfNDyP/3QuWzjC/c2ILZ2HPARXuods7D7+H8OkA3MrNXo2KcA3Pe+8RmjE1Nv5x8LN0Opzrzt
udVW20zm76RkT2ctxmrR5e04QsAFpM7o/5ykkf4jTDGvTQofYKpyYgtduQIRtSQu3nQ9j5/A4AOl
KqREVGrmZaWfGuNThMpsGJACNcbpEtbgiSdStjkGrc/qVHpCtWUb8SqZ05BPmRqBB1FD8L6TmsWl
GF2VdDLclD/TdAdtYj6AoE0ZQgiIVOU8rd9i8CU4blqwEqBZ4NPwwiaBNKNg1tZVrRqST+3jdrv5
ssn290yqZCCtJ5c9tTb6U9yzhN6QSoGDJYYTCHtr/aQXqsZptuqYTUxORAVEyijfGpY4ZzCKOf4N
bjf52PYXPWpyFCWgx99yiBjOhXto3ftSefMG2lmJaF8CznwWtF/YYyxU0wcUn7JHgeD/3X98c4/i
SK4BZp6iIIo64tPWmVgCk3xEklZJH6iwunGlMikFuG9SqfSYfP7PKiUtgkraJ/RUZBM8iIH5x9JO
btiMzh8TzMj4owvYa1H2De/s2alAT0CzOCy05zMhOsaYeNu7ADzKBnNzquPFRIRo3KaDzwxPHMSV
o9wYm0QIGQHTIbtCkZp7JWkAJyz4JLXJelSs8c+msJcN9LlcIhBDGYD+TiPFDVIVDF6veXTu49NB
sW4VjXzqQaI7DnCIl8oFoAox/f/OJbKz1N334LSk1pXsmDm1GoW3NHDySh/uy3q80EpwVFQb3gNv
ySMvXmP15uztMUVU7Ua/N5Is1siNUjMM2iDUHuh+383uQsNVcuqJYyvYQ2Y8CCQSktoC30DxkenH
B54YXHNgXUvAgM8c9Oe/7WCeLXfrPxtlecIE1yOMCB121bOcqkeJroB32vkjoZ1Pl8di6ncJMsxk
AHA5plbAWFfWl3rraLxNnd7nwOS2scKeG2Tphbk3FGrG1wn9HlHxwytIrtSa3rDkHoeQ4XvsbdH8
UDOGVlFhvRNXIY/qVeErfyO0fXLTKgU4mQlku6z6hANZwXhklpj/CgHAF2rJf6yHbgWntcvg/Adu
RNTxl6US4UhG4S0X2Wol+BgbNzbwHl+yfO2Bxps21fYVaJ1HnEQt1iyq19pxKf3kbHiIfziY4Jul
9sglTD9EO6w9FNMlfTcCla+PQRpyoobLXNUCzhRVoIraBn23XqGxu0lHw6SPYDE/I0LHnfklo7Ss
fgY5M1D8nhIiNsNYvS/J4UgyAxraH3OVTlhqjUJ7feAIh6gGU1r+ohXk857bgTkVCjhgzcOegQN/
7OnVTnqBZiLXctYzBKQy4gTDIvrjt0b8syhBzh+XIUJAPwscst1TsACpqe+lflQSCCVQjI0c6mMJ
Ms4XrvujknInmRvMBvX/V46SQ6gCqfN1tDEOm4ug59bPYFovuWjUP61sL5qzuw5OY4i/Ks2LGKXF
ubyIP4Ftk1YjM1Pof+YfvOGZ0weMsma3AO4vP+X86zwyS0IJyPDlFZSGNbd6dvCUnB/WMpCQgUE9
2GUP4SAqOAqrGKCB6TFK4NsfOYwjtLaj4kXmbff5WmPozU0i3QjGdjkZIQifEWtxeIG53O4otPw6
04QrJ1aiXJ1BhBXEami5TlVLHa32IdTR2UxX0i6v5LKVuFTEWXcLYT3TWvNY4Hh8RspL28pWecNd
P3j0CHPE7SDXiVAZXFThMUq/QX4KScMuWYCwCJMlXkbF0qBp18QBUV/WMMg7Wds44sY6PpjwfEeT
JHUiGlKWACWp+il0EGlxju0QBHhTuKnrxjkt2PoXcG4lnSBu5L/U1AxEuiZmHRyb4AmwA8D+M06a
LArlvwQdt9XP6yiykpviLULTGyjlLY1EuOq/gl+/+4bh5YdGoJrBTGE5Zi78ZCJXfXlvO4KlDmsk
3+5UN8VC3WzoscT5LoAn6tfICWk9XhdYVInHIZjbt/ZO5kqzqh3eBw5vanJqChriQXcm46KykbA6
qmk3jfBBMEyna5zvytN4NryeuRG7bDCP3WHKIrwJLnkKis0bk83wvDYWtTlym1Uk7g93dWvd6LFJ
Eb1/nVY1jORJ21csyrXHN5jW975wa+dOGw8tm/cAbEuIukCl9dU0TNI6eA8QY7ePTV0oD7m+tgLj
0KpP3jNm+ANiTTt28sgmIYPp9OAxFVzljZKKZMdMq8ELtCONZeFGX4zamPOJDMgn703s50HSYpzN
oSqZBrgzeWwLXo7cKcOboi5FwQjqb5uc3mlFn9xX3P28lNPXAx44kZVhuVtF4GIQ4DiBrz8z3FXD
PJQVzAnS4H8DnWYUZaQyH4247sifb4t8R96vzducDddnsRoeAxsj4ML74uGAGTSAbElFTUvwFsUG
XSp0I2cuhiYsODs9uKSqJxjTldjlD7/rXx6uqIhlM+m2du6+ACgKK56OiCO57J5t3SCHUcQf8BWC
aEzkYA1j8aeeZGIHwD8dmybOQhCj8WP3YVdugQwYXjXVTBiqBIidQWRITCw1BrJRXh+K6uOupEr3
Foq7zyUdJ+0653Mn37cVHkodhPUyx8FY/YLOS9D1a3g3vdXZSg+SxHxYFQYKm+EyZB1cq86/6abf
qP+scaHPrnbRQy+3PNLSoKyOWNvw0Hhbdx9059d6+zuL7+zjaZYI8iZ/P4AjitkNUc9HZIMDcaov
E7LCWOSkfextcDkzmBGTZ1DOFHWm6MLQI3cWHZris+ypvHNMAnYZ15OI0PR94Og7agH2OofliVUo
TgNxRjXJQNxFQvNC5VFZLQII4Px+TRay4MW4E2PbJvEQQ2uZxFGqarxPJAt0Wf7KuLxOTPsGUT8b
mRFj6IWM/R1UFEw3RJfPcjgTHsBvRwomSUvGUZO4sqvKo4YavA8IAYhtXpH1umSC5fqJdZQOiTk9
ctcfgb72Ei7iFCsb8TLW+eMr1CU+MtN55gK8ovLPjdEK/DdKCV1Y2L55lGWtyTcsNMi4LSqFF4ZK
+lNGBX1cvxC/fADsFiX6iusrnaZDzUZENP0h6013xEhI3+1hRtrM7DxuKhrp4z6I3JzKEPtXAGga
Qf7xUVs/Y50K8FSZOZnA4BAqQFIwSqoDy7fDaYjGBOfJ2M0FMf7Ygd5/A78kD/RsYezxKoNW6qqS
9IQ1cgBtaWBxZyKf9StvzJlo5epacgOqM9CuLrC65LseS8Z+NmGw29MvB5bhmAj62FJ6KpWBgdr3
yBGmklkacEckPWIo2h1xbqcpBKkZ/pGhEZhybfW7ejLAnPb6ScmBaIrxejxvfWmxBU8+e6BwrnW6
OPZorQyPgCT57VXbOLKTc79QfW1WRVrzu1+LyOssjPOwjFNgVLgPybEbhunaCplgxSn7PIMmB7qp
slhEI5l4ODJVnKZKpo90jeUsiwz13H8hyCWfcwUIDhvJrl12D4T4Ju08BzS8siEq7CuFHB9dEICK
hFuxTbJtNHzoVKS9344aSpXmZa9mScCwOS6hsk/5fZwD81b/EzZo+Dm+ANCQ3/PavL5tKvtdWSNy
PQ0V4t1/Ic7Vf+Q1KAfUiqADXZ0F6nel4NheGUTthtKMRtoSOKwI1R5tawe4RYVNnhpK+etfYka7
KMQpvffr4Kuz6Cd41DsGKYQPM431nvaRaQK1IOvj6nESpn0xfq7lQ1fYVzw72ptCayZmmiPRPNpf
Qn/E9FSHxwbbI6uGqhCC3z5+DwrRN+sCZHmMXn3FnxgGsXH3RqDkx/tGmHEdOy74nemcNM04w4QW
9td/ZBNbHdJ6kqEz3dDwyAUw6dzdmgQGpd5+JmQzrUfXv36niyVwPpeDu7J1MvAV3H93Tmq6EoP2
zRAABBinAmHEKEXOejJSF6Ge11YwW7MIVwnbhbZEdEncD49LeC01Ks56oVn/A50r8nMn4O8eHdDe
LVoh3oW2AXtyQOIbV1fGWtzw40QIUxRf73Y61OJ53cf/1JFjX685+bH5mnwG5xLMuVVqXZfAqiBq
Yp+jxgI0E8Bz0EyaaT0glbvQTCyDcwkm39feIaOBajR7xG73ajcEOd9pwDsArR02MGZV8skFI5Ik
yxH1kRrLeFWG1vYtLpbv2s/hprr67UI6zmYrmC0yT3xHqCsZYur5UczJ3ISQ1yLYj7RY9wcoJ+3F
aFNVmXM8SF/MY+AHts1m9Lo9UphtlKAVsi3O8g5IGSHLpED+iybxYT+kp01dJ2skYuj0RrWOikav
ndAaPwpBFsY00+JE+s67REYK0353vi4HicJHVR+5NXTBPnIXPzgzPGWNqOnvBbAbdz4TBwY0PVfo
vvQkWeXbYCnfrfA3evSqgb1cvzkHnAUpDbWjaSQnidLARPBNHeNYOLkCRdjZEHXpNjIyn5+11LYg
UCQHm4fT7YWF8DEQVs728ZuySgyQxWh2dbKmjnNBZEX/jEqblFFxoVk+rY/6w1hGoYkpzpY+GIo2
ydZXEl1/F3QW1hNFZ/6rC62T6m+5sQhUs4/s+lalt4onuOdbCc5qyrcqVvMeDtNerM/wmVR1cTuh
MsxSNKejAGT6irk794oiiA5OLDq1YkDM0RY2WOXI4lXA9BIdePq+xuEFwvusQP3cy29hBOwnfIOk
O+5pVCVLRlFv1qv4zLxidlAk3cnCO/jMVOoiodh0r4r6ZzwwSUuJqwgssMvZKpd21rv9qPTIFNg9
tWRwoZkxldPhT64hxLHA5kmMoRzEhsI1rvEBXoieCBWYfwzMXf45d8mygNhgkXYHsIDrZDoqJbZa
d5Ok721RWuRvC+amsPueXeEf69o8VcmxprSGPmVR2yMu6pOAe9yxyDOHaXG7qZEUyDSdC4qQUUZf
4wIKs4fy/6WLGfj50nU/6KjVTC8jy4gjeylyA8qUdp/gQ5ZBiPnloiZzOhZxnDB2IzAWlqSQQtBI
IgaeKipI3WKts5jzzn3nwj0Nv0xZ9JQuHyeD7WRHrugQOgNIph/F8hCJJGR8z0s1anElrPEghbrQ
YtjVh7UFw7nN7ENPSj2mQ4QuWNRIg3KTJUjBy7x8kv+q3PhFX3zv1kmIPJECx1E0QNM8kttFIp0b
A+pAEAB3GUjX/Kqwk1Omj9hBhC4k0Zz11v1FClfkKDkyily0Ur1yKoHOvDozv2hkenv14OxhMgl2
+UeG9JsXDQIqFTOtsg+CFUczcpPLwfCBXWr7FQzpLSfoY3a8qbuhzXpezeGcq7yjbJnuzCuPuPdy
vY9KSS1yskDkhisBTva4Oq2ov0KNW+d4g/jfwm5kpJxDBYAT7EFA4dcfkzSB6pHSHLSkTEPDPT06
V6Mjex9KKWkCiGL3Fjc3DzUJTohJ+v3IzRJQKCbu7ai5Fbe7tOliaUDjdDAZvuGJC5nPf/0HYP3h
M5mtJftBw0/7mACVK6x5rKfPk6sTbMR5cHATgJ9V3IMWfutEFc8FfhdxVg+p3HMNDHFe5QlvMzlx
5fCJgZfDIs8HOFSRzG+naQ6erf1nBDeHwEBZx/oTobZi2xDtZ9Y9OA+eQLldg0ijy13J/e/zVbMC
YyWMk/AguYf7W12PRev72dKxgWR8yJ8Tu/IZrYvuJThPAeQg0zgfX/18rMF4FaOA6pWeDA8mRmmm
CbWhuEyTQWSMWOavWnUBcvcCIc3OXipsVnNlQdg60XZC2a1acQ8YtKUWsf1hyXJFjEkllYNQgg4g
E6peCZHHKfHLPNSjAUY6pqABcl5AesK0bPixKo+mpH7ZnnWedVvCij/lFQQJqrjNTgIOxU8FFpzO
cnPTHQ9zEnB0C4fy7iBDLcPRZE88bVHkfFun/W70XZbIQ4PWob73ww8ZPJjeSMlpL97FHvQ/McAP
6bAqeYNGCb4JXlXJLMq6CQqYVfMFzIDYL83meRwg0BOz390cWJnteesKnViDvE44HeIvjpSSrkBa
xxlasXM7XVyAiE8eG9/XV/Hvum3enSIyh/6wtVyWE+YLMbsqdmks9vnbpy6jjLn2VUS3gQU7pkYU
eQ8fVVRZAbsFPUhdPHkYImpLZYSCg2vFeBcLQQlUsBM9t98fZuPb4TawaKN+gvRzV6ZvCFcsihA6
cZcrX/EhjTXmlXqnxJqWRHI79exYNr+LKZSo+rlOgJsp5rQAzoq4RfEJ5PGRZTcgfQffYR8tCMUA
HQDkZ7EmTUC/WU9P9HxHZ1wou98Z0VdPph0L8XEqoouVQydfK5j/2dwQ9FnufEH4WZoRO+Pof5zW
f63m/upK+L4hQfD/Ad2hmNQ9/78I3iUhZbr4H/Kp3Vx0uAuHrv9i4q1SGYz9sZqnszYmSklds3nu
vuBtqnGT6UgqoCYM5nF9mD3ZXQL0jxfP6jRYpts/ZErLwCGuZQmquTvN47Rci1NJDlub7CQZRYVf
oeMcH4pHC51n6RcCzTUCSJdZRtVx150pKGd68HzFYQUbYzU3Sn2zWWnJrXt8+0j/ORc0lkULlIWT
psvZ7iBPa1LgE6noGhxF2iquVJKK9LMCFwuU7JCI0ZcyPmfFx/piBCYgmFvtQtNa8AnoQukUChV4
AS9kqF8giC2yzmkm+A+m5em4P1nGDLYY88LQNkjKALajcq2j1LXJMffju/pVRp/l1pwEo/RE0xwW
kfzokCkBJBjdR6TAw61MkYgPF41uE6R7Q1Kvs0KChY2a2xomPEb5ybuWpQimAGDEeCfexU/JMm3b
61WTCvxFFIT2cghfRIpWJLhZ9y8VWn6jKvj3cDEs7ImIcWIpwdXpK+bQPwDpGE+/0yaWnAZHeOOS
N2to9QdKAn35VSykyYDi/MFGhJsFbGCY6/M8jT3CYyiz8aFhOo1dC7S8KIVIhhBCjqRSiH8fMcro
mmhvlnqZ6ByWgM5tiAJmzBG9grChuw9eel66V1lIHFw4yJrI11rvAtcxulRrGdsT3XL6MzP1IsGZ
t9LHCkHUklNLDvqS5kNnUGkzgvMlE0PPUDvQJ+haQfNTGcanbqp1FPec6lqmgiE0Rq2Q33EkffqZ
b6pJi29FLPE8fI+jW8MBZuo8KRWZfsGVf+7HI7jlYsoxfZGk92QqAvz5ZJhuMlfJaRK5TeK2Rv7t
DHqnw92m6t+4G8Qd6agNIj2xZe9BmI7cYIMnIjRwnVWsF6bokoloUjKPfqwlT9S94SNUI1ix8a6e
Jxwa3c2z0oWFH8jTO89Sneq8W5845pT8tSYmYD5riZ9OD+xnZnEvFd4VPmavDe1qNkUegE3wAs/q
UAoSovpxUnp8uKOmrAamwsyNUqPEZey7YUwsgDVkAhrYMXefIWmBleRRFydV8hauxbbdWsxnkswL
CpAs2zzo+VcrhU2K9Ds0aQNmxM9fQSrCzzW8kgXaUdZdtEWN9voegblbdPxKCgtmt6328V4oIVSx
bAH7Lqr2e1Pkk9xcOBV3xbqbe2CM+70dT+UjwvfchHN8D9+2NnG9evxbkYntDm7dx7rGBMxAwwyE
ED2mm150+kx+ZIZTe6IpWg5dqG9t/v3gcUsruWmKaF6RLoIWxnwnQGN8JGtspEEp0vXL5GHvbFyw
XkrX0KhoutEe6shsNqE6T4/cz3kjebhmPinIlzZBkbXttmxC45EyhOGX8kL+PcIngs+eeJJuuLX4
HwupRPQx1kRcn/l4iGywj5PoUxBzkN0Z8bNHKWbquEmGe8YLj3P04IqO6gbG45WPXHh+4p+ntf36
hrMn//Xmwge3MAuteW/3mWvMIkwoc+sG9tLtjK1/8/+s5BYJkl7nZD/ZGu4K885U6rZjSypP8IJm
LL1GWNQIif5h6N4SMiY7Fvh3gWVYzYEkwvVysT10m3vZGd1ay712FiwJiHUk+y0eBUhTwhCbcO4R
DbrU9T/m4uQnH1tBcJe8IWwnaqskPGrH8/YV5Yn0oqX66oiemAFuNSLnILshnoja6WvoflbDY9Zk
4mIzqm2doENK9TJjs/6P0NemR2xH5QE1nyNN/E3SN+e8jl5OAQUqrJ2mbxHP4KHuLbunrZ56hzt0
17n4EGVwcdAJ8UTzZsaWfRlrvcE6KGCyI24DcDq7z6HDVxzjslJuOkHuzHI3w70aW/Mu/dKPmL/Z
9SK4aoiGRgbTXkOulk6ED0F1Wo0Fs0RHzjSuaXjE8v2MPzNtM8NGt5qAY+uEJ1JIa6gjUAbJ++t/
21wcDw1UOJcmHyKMJxVOV4cbcLE9NKnBY+Tewkz1a8LZ2YazU0vklbUdxmiJZFOZ+3+aicjal0hz
j3/VIzHzIXPa1vbabTub80WVdevgAWGwy4h2MCMKSKnsMY+jqZC2Ieu7AYE+DFo0aI8UD0FLLbt+
zAinxrOlYiRW4mUyjdYetplQ1Pgujj3kaiWt/qk2OC8ywFXIWUr99z1DP5aYmgyb9RpPUT6O2zJW
Ks8v5+06bgapuskw57m+z/7ApwiFkTQgTZ5x0cqZaQYxvjdsbBnj2Mm6DCB5266m8JXiQnvFG6jz
Oc9dZBfrrSabLx4GzLqFMVtCPtriUh9XPE1j90/Rrt4CV1FnkkrAxh3tOi58eEcfl1Hezr/utMii
gh3StaAM+SOi3n60NXiIy+ZnYxM3WFIfQZjyRvtjP0KlJKtHBDzBF8+Df6/7E4lkFTTxIzDiU8T0
ubPA+omcAglv3J7EYkCbkV8B4vh04fea1eMqM5uPPNFi/zBCc/XKZDfgTpCrAdwhyqcp1r4zK298
n4ViySY67HjDFo8u6V1nQXwBPktT8UcLGfeQu9qAkYp/01+Sub7GdeHdOL8tBh6poVs9/b8Wissk
ZlQMGzPynW5AwekJJ3yR9Fs9EkPwRgKzeCP46kxk+u2bc0uvCIVU0z9QFYoHz9K4zc5uhC49UhpF
3XGil2biMa5HzdSkPAWyh0DHm7u5kIvBsjTYlQpS+WXtxPrcQEh6Vek1gOTk3YraJA3G0WQ9FlAY
bPc7FMLBfOpGziwoIqzAZQK9tB/qUXW1683H1ZnDBin368yhwGjNGm0QENouek2gpAGiAiWfQnU7
nzm6/sy3nnIwHSi+b/zaWzjNkgLurhG4P4F3anXOk0qq5N0ABqJ0PLV3SRkPpGj6EOhJH5UyYXCP
KiA6CGnczNzLv9mi/rO30otK/nr7GL4IY6bvADSQT4kx1KIUEIUWcFJtwqnKYOhHMdsw55NSZipS
PwI0cWY6Se0FESc/oXxgx6TyANFkHLQNucKzEQHcB9DukbuKXrIi8AQMzuqvbJXIFeozcdWTJz1I
OdWgkqILa0re+hYOowC7+tm5O2FAa0e0S8lUN00aduY02oOn1cGeLAOajeLdiTeanxI6jxF8Zgfh
rF9SRZgKqez+MUuOsgqFhpXoDOcH6yVXOo+WE6B755fnwpEgnjhYT0nYM7aVWZij//pFiatZe34H
jXXpywhnu47z1rAOfgQMSVtqT88Y3U+f3YXPJGo/JDrO6ZgqlWkSYF9ppxGv6bBCiwjAaLuXJhT/
9OqOqqJDhouAoEwKjPNdXfdP8lNFPpCmSFKBpdtUp0b3Qcqbt/20lgWZ0X42Ie33puohpLHoG6Ub
HZTgOz1+5OO63l0w0o8DYS27q+Bb73+OqOWGXUDgBUAsIKG6C5jH2vHiumrkBaFQka8g00NOijKP
poMS7TU3659RbP2kjx7lxSkCsLFJnwBWTKamtTALD5tsm5Bz3K6AYMpzt4rtgcOHgOxO9t8SFMCL
fxEfFe4TPzOEijMjEcI+8nR5Sd4lqn36bwJfnFgEPLHeEkhVGpyX+sYvOlyH3VZ8X/oc8jgtXiMw
8Q98hSUvOaZKVxeIjv22ds0BrspNYy9dajNLy67KCXBC5s/txjaczqk8s0au0cfMwoI0k0JeWsN1
M9uktu8v+GRJh0aTn28aoIb22BAhaxH8RbWMHPVxFfucIyfU92qMbX6QxpmElpXOp3P3r6V1BTaw
M2QJeyUwjSMGQrmurk509IUycCcgIJdMMeJZGBG4HCPfZqn/MtoHhCNEX7E4Jcro2JOV7al7zprF
4mnjlugH/lLN/czmwUIFFnnlLNwV5IAzvWaHrcF0Nt8O24Gv52r0xxtaPG4bAgxZ8Ip0BEEf3Bcs
+RaEBAL5xClNdcVe4vG3b21P7P9RZaBID3isEdFjsv6QRTyDFY3suAdErTJBBPg+QYlDb8iJ9+jF
+79G4Oy5sCfpn/dIJL9nt5RTN/iRJvI/veXRhVBzwTqw6vvRtGI75/cDzrNy8nbb4W+Mkx13tC8t
/FPmQ2ChYpEPzupcYQIQeNXtA7EluLTvmadWtuWx2KNUcrjKNr6ISlIXlyu5Z2+a8/jPNlwlqsIe
uzLmqfr4e0452qPhtPsyX8J3zU62Tl6zAW8HivXdsMe79cfYLtl7fVJAdtEDwIWb32PHW2nwNOBX
NNH8NUKwN47n5fb4TJXbJiFAc8gHrGh8OuYv+rlZaezxj4SJoXU/aSrywzg59WMmMFqO8ppoQiMt
fp+UF2jR4+epr/vxX8BmDkc4PICYVWArXS56SerBTWtrgcicANFzOUUQ/Z3HlIX9l+wG71o5mAOe
5AQ0X/ObkRszas/xHOMX1J7p7i1SnSzlN/hhwL4kspgRgnUn8dwMTN21UtQB+ozUY1hB83hGq2hW
UUbkuoRtb9vtz7Bjkm5Ex2GDOYK5JuN0A5AGBNwv3fX2+wMLoWnFdYC/qXuVEnrIQdHjyEg0JX3E
60Dci+jf75JRrPSZr8ZBkWY2Egngb2LzpzcCETWLadoOBaTj8vc/BhU73RdPjhIoaHnyuTff/jdH
4fd1QXLEmp0SE8Pc/A+HeUh9S7K8GwDv7Q2eL/wQR8uwiwexBi9nc4GL0WmON7q5BlCGE5AdH+2u
uXlL1VgaT1hvXr8LZaClwOOcbr9mkzdILho/y80IQZeP8hJGpEusr3r12PvYZnl96tR/ZmHaqmrD
L1WHWOW0wj8TxmG2JmSaLtHwoAXaoiVV6BAVL9tkgQUPP6Ou+hIVFQE79EpdDXOQWVERU9rL4KQw
S+0dhTOuqM+DKHh9CIT8TBbpCfDpPLDmgymIGfR4KfcXOhtoYGDlWiD/YrJ/BMsWGnkPgSIcpxv8
YKHbOlK/Uk0C/1EXYVtM+obf2YFQP35XW0r4U21V7dG2GAte1QXGvSSmGOPbOPwi5JNG+ktX00++
IYox3dSikHMM9dOz4pY0TUD2ywbtVGriM/+GwGJCJRF/5HjUXBCToXcPPYIgRgpFbB4y3WFujisY
uPp0oXH4I5dgBwhPtG8b9BHZvs84w8rlK6Wr+BssgDvsALIK/z+2dMywIh98Z/dVSmP991PGrHdm
yBZcjB3KaOuRc+yQ4l6yiVct64xTTodJr3mf7daj37Mweu06ECJJ7KBSDcyC/A2LmKhCnu5O2/LW
bFEXpPxcgD8fyAr5MXzxdqyigUp7tAOyQR0iZjBRBAIPgFrCQ+7Jv7WPu3QPEEUOCz3t7ZIgfO/G
VSWfkbNC0qs5OsLbBPSC2aWO4llJPBIqJTLGdh/vhhjgCkBU9hzWIuD4hgVClE4V4kkX9KR2gvot
p6MACUQcKcU2/n6mPb2sAk6ibwbWTCaadNpMO07joQyO6tXJ5Q9SZezRZEC2bOZ/9swH6W8eR8Nz
uzpStEKzQR5Lx5m+NVsvNigYfp2Getpv2dFSbvzXDdZB1fGuoJpo5AbBD0d2lMpvX/Yl8Bl8hd1X
z5BPdZyVteoIsPNQ5ZL5D+XD8lPaV1rm4HiwZSpCMMTndbZTSJE/DcQbORi3S/Gv2/Ptve+H98u5
lPvZDJHTifMR7RKEbI1W/HhKf/2TQp7XPWnAaWl5pOJwrzW5t7uc66bpnIBlNOvmh9lAHoxAcCJL
s6NxR5toOZoSyxUWUGjk9XLKX4Qng4k5kIAP0U994rJG3ksjdsM4dE/E/sriVg3jAajyV8fiTfiv
eMlZtsgIM140dNGPgrxTay8foQJvVLS3yE2r+R7WruphD5S2w8AL0s+xZPgrBVAF1SpD1hSVs6iF
FKd2ed4/ih+6vgOcuOXvTw8VW/FkyF+rO29F6h7Tu5ev1uZ3OGrfhGYN4YwhadiYHI2YweyIW5Fr
zp6zYBEywQNlML2vpyRRsHFp744Fy4GjatBtZHTnLxUu1WNwuaS6Mf5Zb/qOk01jpOz8n4eT6IX6
lBYhOeL2GIa21KhD+GkdgVjBMQb0gpUPWa0UN9nhSCQ4Np4HIWwbeOUXuZZ892VWqPhcXpvq/WcA
LXQjOJSmhG2uLRvLJGr1X8fpLots/3zr7nr0EAiRDnkcWi2ZEg/wnH6AEQwJuU3evG8xZgt1ZdFQ
TsZjbpXnwdqwySPTxjgqFFR6kNL+Dy7y9BfoaxYOBtxZB8IfzK3RHbaQWqQIheoeXBoTX+Wq5Z9+
yBZyPHL4K2tiMKkSKpeKwIxt4Qv3aQhsHPR5TUhRyEOHKd3dhGqrIEZB4YwudZYIbcqlNM/7V33d
Fsr3Q+r8wGYvTk7YUOPBDlVFe2DOqrAabKdvvuYSk4spJ6U1pdqzdD9ocQKBgl1wQ9TRlUVRfdBd
ZFxgv8S7VzMoMMPmahHtaLnrgQqB+vwQQdZV+Ohv+LCmM3IfsjzR+Hof2yJe58Gi5HbSEXfbbXfO
y6UGpwhvMatScuAm6fpH3R3QybO338Aiv0sXqksSpSWjn8Hsem2pDWua/m4UT6TP6xjaWhXIjYjq
UmEA9IqieqYQAmZRiqtcNWHRjH6PhZ2iqzv0SB5AnqQi5cVHHqZ0TptfG1faYN6xfj0KKATRJHhy
tmqkjdnBJRzU1WNsE2oShLkswnabajbj0w/W5tw5AaIvQzPLEL2eOfEXsz/CajtfH0T8h45eGuVB
qYLESb9zC4OpHBlaYhso1ODDEmrtXB3cQ+fdLH3raoM7YhbkoRace2LUAuBHVK+qL0GsV7RYHj4e
AYL0Y6G3BrTvMnAs17X/5DYd8WNhTB5rgVs/f4rR7hZiy9brENM60X5uVWdRVuPxUKJ0TuSz6u0A
sAjALJfAU1NN1jbOziipo7+iN+fv0o4/XzjoflRT1qd+RVQk/nkFu1jKFutLrKH9S59BSADIqcEt
NdIhn8/949GlkxGaKR9UBfEXLuatOO5kCnJHLOmS2gEwXGCLZfkzoeL+pOkJ997ib+B20swMccBL
LxehzPKhyTaYaHZcntbBxXo+04m4qc1h+m0ovRbM19PTFZ3khmRaOyltxh+75V9e6i9JIVJCfm4v
jDoxd+3Qn3/yD1vNk8CmkT69FRzE4TgLaNx3RQm1+1Kp9JWM9bRN9tcAi2NsixqJbw7j8t68Hz8k
YPxwqjJbLnX3s9NIuXR1vpx0YVi7Ey7BaSIfpljvAtaav3E3Dg5XDQvSlfcia/HWPIZ4bD/q/7o5
yYj1fsWgeQ6gQSCo4kBVAzBcv34HqgdZl4Lpl/knQm+wFR+m6jDn3xNC7FTuWNpAHeJaW7jjKASQ
riqui/g0IoRZ+2EXvJvx5hUrBR23l9tyqzurbhWEqUF9v06vL36+aNPHMfUYXnsuInpRslJ0w/EP
6UIOFB2W4RaNm7Qz7LZs+C91D4QCJGNZSgLgpc3/HPQE8lluGwTT2Sm/uE2tm0PcFX1kpaYWOzUs
7O20gFbut3DMsyzv/4TbulegfKtGkflWF4vWkA50tVMd4ccj5ocLhYvfdsfzbpgU/Z5E2TwRUVUP
SwLJvfc38SUzKRrPSmUxUQWLSa++zmLnLLCoOAQttlm+lWJ+wYlPJz9lp2l7DYTY/zEsNKugv7O/
MIw837duJ9bWKLjOZPkZgdewnk+3Uj83HmQ1BzlolzGbBBnLF6BxMQQNGWzwbdRw4I6D14oib6+n
Uv83SIWxVo+qTJQDGpzMmbnbQxO5+4cs9RmHH9bcqcmtWCvRvpUPSee9w1XNZ1CmjlpJCdDDxmTr
OumSyy0u98F5R/aGoHrAnxE6Zw/8NKR2EJlgLvuI3iq4zTB7bjMXGzfKB3gg5h1H7BDuAELisEj3
T8pr4D+i8aWhqNx3eUipNICI8c5isdW/BzsVh+aeLXLhqbYQZEe0JbV18EKStBohkUmDEHVl/uSU
SinTuQTC8HKcAYNNFiq78KvaX20MHs969dQnQpeDGzxZ7Q9Jf7e28olK/otAXzgRKZuMc/sA96QE
2+ABrYTT2WAWNyoB1CN8F3LvW/porDCgG02AZpDA9o5TpwoVP5o6YZGrZ9sr7rNc070PMsEjxqPk
N1oPTWVMrCzHuX7Yp25kNDA5WsVAmbi8Z09Q9k+vS8Iqd0QVlD/tAdYWdIRmtOqg9FAd4FktEv7q
Bx/jMQFmmJY/cJIdKmE3o5e8e+PWl8LDp52W+q7kia31jD5D1uUHMRU1y9i8VLbGaiV9+nJxJTtA
a0VjxexSQlNRg7UxPRdPF8EGGDReeWxkxKb1mksRIO1KxNeYjOp+NY2K75sEzLNaLoalZIVcHv9C
KWux0j2lD4WPu5GrbUU2EEmQ7AucCztwdzkGyFWqQImabDLDbrwWs7PWAYrhe5Wfk3gmVplpXS/Y
N0MtHIyZpRWJMQCfqKPRBSXwB1kGhfhPIMrPMn8qrm4mWASWbhpzNNW8wk644KUWc3N7JoCu+7Ww
vx8ZPN5Q5VDDcmF8jAuo+fYDm+xTPqo6cibAqqQvdnl+nd+avfeS611s/h0HN81zgGh2qK3Nz3Ct
yNsABxBfoEeINm5eG1+bN47RlahAdGQXmvrFZJlQbva2zDBJx7AdeZtABPfX4vfeD7pmaWqHTrHG
baWj+ZSOfgRY96ZFSc/qzD93eqfKkTbM6paHm+y1Y2c+w+igClsqIcfoGTNCvRv1VrjuIVif3QpJ
EBxxyc50MK28Yu+bWMfvaFWHiqMAeXlm/PyknlvWu2yIv1KdEESMMZELWEzlLl9diqN2aHbuNsVx
ixWUNoqCVJoatrHL+ThLw12G5d3MMVfEmaircmK+aenIQc5oPsxp8ag67AfSpYG6kdgkJpPUZTWG
Vb+tSfFKuQug3VSlbntAzZiRplTKFCCbO0OQdO8/vN+aDRgPRNk6ROt5CqqnR86NUDpkL+Lwz/vg
vy7EmJ1QTaxLdgacU4V9+T4XjqY5CT13VjLyfaJjqV6tQQe3FWzc5ypqxOgJ6MjruwBCi5L2zMn7
MGnRBJcGp5YXiLgeEOaUmj6PcSPsnka/6kcX+fw7J0pGvWyw1tauzrxCfCT3Ka+5v99rfOLmJwW3
Ln0Zb63yh2467QiXeiJ8f4LvfIWYA/vXrKV/A/hpejBG/quRoXXxwqHh+yB7O2ivP5mHpa9fgZ+c
vs5cU8lyIM2b1MSIXlFZCRFoBBIw1RmKeTszqm6xERT+UJTSHEh5HHgk1P3cubGTztGp1PnBXin/
hitmar+v8r2QoY6+v4zakDpz15Up+3/vCeoo50aX3enr9fipSNj3t64dZiSH7yNj5djBP8VUHq73
FNxuoF+IIvBbz8UAxQtuCRS3A82jluq/9Rd8MOwjeutkAwWVeAcx3mP5iwj17OCbh1fmmsVA4zsa
snwA0yxL4nC0NyDuRMzUS8wCuqcBEhRMlPV03/vuyg5x9FnIZLmzp7UupbslLmO8C2KxGNcwN9Bu
Hoeg1e7aJe3bqgVgewvVJfecy33dssysBercZigQGAFVVeSqRP5uAZObLPLI46LT++m4HSxYeqKb
SFKYfPdUIfiJEyDl+6hyuLo5Ej5zjkbgwztB2QlsTyAaojlEkff3QE2d9s7ZjC6In0+ofVMxu+1A
mmXGT3fEQuIFgNoap16uQASDZHFwIgXDTioFGhcSI+YQF5tSY/wUH5P/q8g2QFeNmSOgNWJQDzBI
5YxEPG0N9jAuewBvJtNGHMFMFSGyfCBd6KAI36FGL9vjHzMHfM1rbyShEmbhcZWv2S4CFSiqCSap
GyA+5xe2s5B/MIdWXtkZtADgPVRpgdbzLOVxeXwcWsY8FrT4ItU0Ybby88+trRGNOGz6MVDPQa6U
2B8vz3o9OZ6szIWCSAHJ6iJCNNoRsi1/lZdPVY9GyTpAGeePouti7aCe8EHS0z6c75VP8+iAXPKR
Hler1WSFQ+tbzQBXHaILG9hjwVSv8ouzsxESxGjIVcoNyIK4PNzpFTFkqVuU39cVIvUicJIOHHLu
ITvlT5LCXBQ6xsFvSVh2lMkd3dRCIuXNogJ0pnbkIsD4XnkMmO8QeiuNc8OMDU7pVE1S2e4MSngg
OTvCp3NjxOrI4yc028KNgD5nQYEbWfaZCQ7mm2uDysrzx+1fKHxEa2qms1kDUcLMzLSHxn0lgMQA
dUdYcPjZAI48x9KwAOz1r7OrYo0ycEymDw2wo38VhWc95jiRuE/6Q/I6P2GHW/jYJx3W6pPco0jk
/cZjta9V1k4SW2E2xIzt0tGebItA346IczAWmheGn3r8tOaeZhecIqb/A5VHHt8MeOWjhVt/wRmC
K4dU+IISMherekXCxT9r/nspX5DJSkP3Zeh1NMiYQajqcuT4dEbwOQ7ZOCGy/BqP4f7x97EsV9ae
/H8rUjjlr3Rkr6j1KXMVJ2x3KCTLFak9gw4FrIJW6NIssrCeXya20LKOFfSb9ozpuKbxbEXvtx3p
kI9A3zt0NNsD5Rnllascl/9FCXhq7s6LoSv1NqIqlmpMklkW4lNs3Cs991HGQT1qt/wgsJu48SS6
IV3qATzKUh0stF3nHxeEZwadHvIBCiRgwwAXKxwgHdfBz39jow4/RO+UhWaWr4lwKOXiI7bcpUCt
oN8prcH2lED39JqFSG1DrU8Ly3/3PlRQZTwvyfnzZXLhfj86UAjcBPjD34VcvH89XcUqqFl0qnpj
YOR/i2pmAuXLnaQAVhlR24dID+tcD9wlHukJY3WIjIVrijMj52xur8M/copvpsgD8WvvIwqEgwdP
m+e9R00ahwUzl3wa/O9xkekjI65AlRTynuIjuurWnLuGoQsN0jNWVTPtq2TMxLi960C82TG7t9KS
1hH7vOw0LX+1/s2NB+flEcU69CTWmgARC84icR9n297ae0TaZxEu2Vl3qraFVVhp0qTsKm4jXren
88qVi1WtSNa9/QPKV7tXb99HaIxXesIrGe8cHVi4S1l5tsbqkM1UV+I89K6BZzZJL+KzKv5YdFMA
GgAfCAdqICxlqFvDhViRzTzvpYVryfRlA+2XKVvOLzLpRjuToGe//P7ochHEMzJsijYvB6FQ5cpg
DPA45lyOYL6LsTPmcBtNiRfQJei3vsSTKpuM6Mkb752R/exqKEucnzVBYw7Wbz9jTsEKWSbN88i3
CAsuHNyy7Uq2YUdRcRHB169jI1nGqtQEiKr1DWHj91l9toUNCG6K6XIbPOs78QTw/uUrogXUZBFG
qkr/vzeHgFHsiSygF+1ngrV0fYQfx249Vmn0gCgtbVvBHZmnSBhfuHlM1/dF5DgyiVE12E8da/Jl
6AEJ7U+8iiiznF7onBQSOuFKWv4iQtQJVPC3zrWBXqeo2u5d5L2mnMs3M77LHAUk9ov9brxX5J5p
6LZPjqFU1OxC7M69BFlQNVsbr/ZQys2gkxRPA+JJUs3XvqVpDDnlmPyD8SY4dod75SMCkF8fBwuz
Uf4WJx95I6EAUEydRkmBhpbqM6nRn8ypPz2bOSVbfjeGDCDNnOMerFTS+k/JeObQbXRWzE1OLJmZ
/tjxcqDvwMPKl0mKvg/tjas9nuG7Z6//XeXfi6ZsqjaVeC0elGX9eRUlCbi5SKdqXr2KXQH57Z5j
nsMRaAEdVFU5alGet7e/6eScgEuIzvqwtXMu47vAuf8+ClZnlCSEesfIGwKFGBJutxK+ry99yauA
t5rNG+N19r8glzr2uCzzV1DHo3fYw5HvkzBdaaNxMT6UhMtsCR148g6W5x9SvFGKgs/oDN4AG18D
xZm2QyHehjLC9uCHR7j8mqJYONxxRhj2zlxRNSXwQN0/ODhDjR7F54mqYYwZkn5ypQI8yiK+RJSp
oM7Uhkq71CgR6ocW9Z0rJ3mvXBiIX3azEBhtoZlMBb808d3nvhQg4AzZ6RaTVs5JAmRgDq9yv+nU
tKiRyrIASWYmP2ZSBVk5YEEjOcslSg54IHDkVGKuzZHnbMaPEiY4zrmOpEBwgrNjUUo/f1UoBP1V
Gx45miC5CAs9xC85pXhKwFI3Zull85odtOJ9G1teT4wYjbZ98rC57pX4i8fZU1F+zx/9fbt/sz9t
dFXOeIkmgP4jN/U0/7xj2IoIYRa/xiRcuGFMpMMy6qwahH1krdNV27UzKTC5RXAjx8mIYWiRyftz
50uNXQq4jHH7VQtPuQWLJ7HH4i9i4K6mr9uSFAndgnZl5UT3Ppygfxh38F+Lqukk0aUJtjPAmzZL
xF4uVag0iPNYfQl41rR2IsfNkuomLPEY2CzITJDkexujam7GbFvTL7cvOSuk+oBKm+N/qDlKUUm3
R34UJGNU1tW3cCCF4B+mW7OZfMFTiZEuc4kgj5Duko6ETeMmmTa34lg5QxEqviQhfF8xYEFSpVxV
VU26eNAcpuVJan4wH8tIV8qNpO0XcSPWebbR5yfTlxGvt8jalVyTaqzid9IfAJt6GznVYUrPhtD3
DUPZsP7eOmpmQDkv31fTE5dE0Kp3LVbTFHnc5G+fJM3FbttLQnn2xEz4nONPX13hegwUVt5BqBvo
mQCHsk2dFaIsl8VR+Sx1sEspY0qkN0L2hooMHW0xVY0ccRLFi0xOV4lTeojvcv3OwuN8S8vKIoX1
24/N/kFtdTgBRaPSNlCuly1+jswwrbmZRVQKUenrxvlTGm/9tdY9bFBbrn9YweR3QqdZRZbpjbDz
2Xvc4X9sJ5MrfeFFKBA12dv0lPrvp3pecA8rF22JeOTcai1SiRifg727Ge6d2gPysyuy2zEltlIX
rWmdsKv+v7sNAbnv6ohDAxzewYFLT+8SsLsnNxbWOsZjjKjlhQiHO+kFgueY9CntO78Mx+nwY9xN
of7mNTmPprKGIyHS3V5d6scW6UVkCs1s+fvxqBoXp6L9c2VbcKua9e16EUsJAiCsACuj9MW/P03h
e7B8oMHhEz69JKjzzdOJl17/4Np0EiSbPUlFeFSdLmaMGIhmlNaC0cstfMTtjP99V6BFN3pjziMj
FtGI4gNUbHB1HmylHh/Qe0F7dYwBjc0pMeFWpN3OCX1salykRZy74Hwel5bCWby3bn4ndRhjppRK
4X13B64VOnxIFhDQ6h8CfhKvghzbB9KvAXFJyIQoOMnc5P11qlAfkn+dlFXqzv5kJXjr5KipMF0x
4rGVwNTHCOTXP4n5gXcXRWX73Du6ojGJ6R/e1gTS0bXKQkoeV7WmjYl1tYxYt4bwfrO2qDtgZLeo
31X1UU9bx6PdWjr+Isc+dEq9GFrzGZbcCHu7CBhLGS+CretWEZWwDqKTSgA6LojIJ6VbCvFp/O+u
/pFNfohDZlcnqr0dObiUirtC4rsQ8kZGqKzro86jTtxRiD8CZQWJwhR1E6IjO+O1kKddQF/KIZm1
5NVdMVZYvEWYmAvZL0iI+ro1MMDkZmzCNdzr0EYJerb8uVDoP9LQRsMD/iuWHPLUGX+LUL6AjCvr
LJ9px0tzWm7IM9M2O8Vj66gMQ+7RCbLYDomVJSWYuaXKwaxRahg2252e9njmRnNjS2NT6TqZlot9
PKZquMnJI0JhypOCtgkDjxz/D4uVhT0Np2r719Tyiad6SM60X+PqAS1S25wyCYqgkImMad/DHvoj
Ne3oqCs5Jpr8t0JCOH8xoplcUI3N7/lIUcH0WGeHjMHOZJf6CjzsHTdA81xJ8JBPnbtaPNvcK4EX
Qb5czYKIEMMIy/2R/GCQeqq9wyeGRQfNmAS9+fjPFEAmvB3y1DmNJeR52r8PBRQIDp7lkxubBoxx
Rnox4cl7+pA/IJDpgsEKuhubwLU1tU5ihoho+VtCB7JdUaKpiMBek+Py4DQ6dA5lwBoG7WELugWA
th60d7PLU0SsP35CajwkFngWLki1SwCtPZaiE/H5y2qZQ0oyyZkI3t1eVO8bzm57e8QL+lE6g/2y
+ZWl79PtqRfvuc0GPwXduLVTidObvWWmPi6wzNIpOswRD9D+FPPe95HT9AgOFW5ouHL/b7EqawRy
2o50pY2O/pfBAUbVmVE4cOoQfdsDyHReLi+dQF1IGpDZZbAaJQWT8Ld6F1aN/E8oDlfH4BbA/Yla
fEcwZRjltmFHLnA9hGQuYoo3sm2WOR9hxoTysMQPPYIH/D55Qfhk6W0VFsiJiqaCgXqfZKmbc2rq
hKj2YKHhPTElyGjiJ382omvFs1ycUiH/1DTiZeuyhSGuCzorFyQ3O0D/TMxe6Nswg+/fVA5+x12F
LN07fdgJ4UWGz0n1C1m4pS3bAzKmJxS//1tqhDQlk1WEGPDBBrurqp4xgbas0k1T3lxRdd/ut4VZ
5s+jU5AYfvyOL5GW43arz8uoJhXg5lukp3Qp+iC/BDg+tVxCQ7QDmlWeY6Mp9BeHoKc3gqId8oZ/
sIjbp2pDTHSPXF36WvHRODD/Fv7ARI0ztsvvAwDOTM03iBSe58gDAJCY7gEzgWiQx9ZyoGXyCfcf
Xr3suWqOFP+Q1Ju74KD7FuBPpcYS4shtAWJzon6y6wggPGIsUvDmJ70wPXyGXtKbIGv0aTbvUIXE
/rBRZ78tJyLAxFYaFBnMPIh9e5WnSMav1nDqSIRVZIMmSUIUvewoaEhK8b/2QyOJci/rC7peR6DG
0qZfXATXqqZqEw0Tg1oqnQpWlanqU/OvD7vN9BNVp6lHPDOS9DESAJEkNUAKK4BOWc8n5Nwg7yz9
sosGIjNa3oyOa2k9cnuNMGob1GEoyPzdqbyCk4ZH8Rgkw6Ypo5QrxHGfTrSECmKRo+lMXGLTOrlb
ruNw3Vw5y7EEqdfEMQelcZOVL0iuI/B15B5X8d4WEYmgSDdFjjqb9YpbGKufVUPm0njuirF6jMeF
MpesVQHUIfKBJCH2F+bHeq8TKS6Qh2PmB5pFPjsKiJtY3XfL0Bs0fv5/NH+W/WJS/IQWPmINkPkp
3F8eRmxVf8+25pA86Tlo8JJ4xX4pV4Kv9sUeUbYfMPopH1KCGgYuADAsQGz6c/UgW5wS2TmyoSlG
33CwaOr7fy+7BrjIY/XZqSSrnfGWwfFcKTMSeRTExVpDhxAfPSyDIlNUg1cE0TSXEwFLD1IfH6De
kcapaklEtQSH6YminC8h/TpcHd1WVFQsCEN/WBQZPiBJggRlzBMElEWThgKBM38alqSqN9NMa4WF
DG/YFVeuSYjAStORtA7qFFLyLK7kwxRCr5VGrJnz2PWchw0hVqh9Mk3RsrB7PKKfDqjPRLvJQW37
6I5F/k0FCkYHgMNveUnEK1J12aqwV2zSGJWy8ymZh11msBZ/GTSiacFQNHNdCKYzhLIt9dsFDLkF
6hPsYth0GGTUot15HMxOcm5RUIa8sfoIp81Ey1tVQV8lc+5Y6O1BrQ1rIyHpKUs9IBBVtGrpRgh8
EqEIM1Ke2xVXKk9HESq5j9X95s9Qh71QzdGD+84oTX78gH5+ScqrEd1iCmXs7iBJJe8ZmuJpFkLO
f/GP/lbKX76SwPLDo7ZCX7vJTqPCE1iDNSPO0x/SPp2cIzqrcNhiJUC8P2kN9Qm+LRjoy5RzF8la
zOK8TAoLZz9ldgHAzvjpzySnLBNTwk4fE6+ox0eZed2shY537y0/0ywuh0O+VktyQFIXe1FFUwK1
Mf/V3I9FxYNjgzUj4Kv2JZUYexpThbYiQOFnu9TTW8k7aQAVEh/Y7p39nP4KVdmCB5jrizeY1W/k
dznfunCcipQXUJ73HlfyDuQxdwWkq+lYf1LlQAQiP9aVc9aztlXa9tJHCcULD98LZQTuoaebrRnG
5yHT5jM0TNjFOfdegChIxfkunUK0vJKQD6dhjDerLu1JHJrXr8tSs/SLO5O4or/E4MeksZrZhL0w
op6AzUJWFE2r34JNcnOGEd5y9bPes22JNIVf2xQQNMm86+S5bvDCtFJswzEpwSQQoqV/EUBHNLuE
OtUO97ionvuzOes4pLvdKcHNBPOfudv1bBqkZVmalOoI+e7LIuSk+hvqPNL3Ri3Ke86+IOg6KZ54
3tbHExIpaSg1iX+22iA9uKCiiCE9OVnV/TvP5B+ZdIcq+wq9ve4bT9MgJthIyg79pu1o0H+C6N6M
t0feH8DHMYIis/xOHbEmVRo71fIEvraqjZEhmmJJLu/dnaTpWyABCnoqXbEM4l0uKUVdNou3da+W
W2xsxsFfj2uN/snZ+Pn3fTP7SY1cnvgJw5nyFGEcVvQlXppyq+KkhVc5WRSGIVkQ1wzL8jnYKCJe
YQ5SyNUvZkogqaSM0mYdBuhx8IpWIhsPpNRfKTEPR19m0X05rlQbMbeeqYw+NPHMHOYLPoglcl3u
QcGWzjC2VW9vSsnxbRZYvKtc4oLLcPLuji9E7v6TbWvuYHdQ/bKcKx3VH9MqwbxO70gCKs339Xra
HXiYxYpLn+8QAFQC05W9E5FJJhPLpEduMAvgGeHJvHWJayvBai731wsrZcZjrxgEHshkOk0fVM4i
9pozC59RWI3bPYRjyDEBe3F4WNV04As2nc3vZoav7deGUV+G+R9KOgA1aJOIafNXoh2D3sFHPXfy
Z/5PeFhYOSeOYgcV1vlArOvKNL5ss3voPIeBQEvfkUAEBr7st623xVz9oGwJnSTyL2rENUhORYnN
vuyH0Gu4kbsK+ODmIqNzvVUJc7DSdp20OHFzlSLCwK8EDErzBPQvCdpTo4wO14rdzc4hIx5yLqy8
QNdkDXvso9AFXa+9CcCnyuNDhkDAsAp07bOu68reh3Sk7BQ9tFisOvtSpv9o5ASfYPg6Uu+49T7i
BXmd2iMt4nfRqLg1RroDeQVztbw13xw/DzWMoZ2s3sbsqSgPAfwVzzX/I7N5CglvNnIm0etoclXp
Z9kqmhkfDgUQBIN3U/bYr5PUdwUA6rDJndtbPsYn43//tG0NCAnOpn+2+SIJVY29vmAZTP+plaEZ
QXRe6IytvrRuF8N21t5WBlbqV53VE+RDmFcDTorGVu8rZm4S55mG8WyBpTvpRPCZ1EFuWmr+jvQ2
jJZmkZiq7wEhOZwiNEJMaDi2xTtBGSahkGwssEq/tpLFy32k0zDhwBKl9+Zl45SZLXEcmp3Sa83P
WQdDBK93fdQQDTeDkPhwSAU2OAfOUXHSzC6Q7cgkZ0/C8UFH82DhTglT/anqmt+AjiKs3d2QzH7A
3+iJDZaiOpFcen5F9M2hmivy4AMB9JdETKtP64W5ZErxbtFAjfmwRUa1EarAgYrc1qyaTER3Uobc
3fwy9rhJUhfjQxRKLQCWrWUrei/0VgcBS2lPdGRZ0+IDg/HN0ZHEyuFBbmQF6cG3VASV7twKQAI0
HPbzt++18EdYCd70E1Vv13uwap2VvCGfkkpz88acTfeEv6Cp1Ym1hr9fo4H7Invk98AJTFWx/+bK
hLjUm+sZANrr2c53Bg7NtZWUAEzsLcY0cbrovfuHRG7L4r/tyuQ4SA5VsvBpGScR+uqUjqFdK4h1
Bwf9LULK1JMfAJN5OnR45OMnViIurAxAAD6PdLdIRl45roDcJl50n9S+7O9B/QRrqtXUg8ROFRB+
NG9gnql0TQI0J2jU2IXtbNlb0qRylglOtB5Rbj85rvuMZTl0jMVR3tCniK/aVEI0332+D4WjuV7u
Uhtk/VvpyLHcrzr0Le9+q9r30btpzGpICezqkJ7PJlKd+76O3tnsuVL0Za0KcQTrYdbGBzdmnscc
o3XQWCCxq/4SeK7l725Y0dqR3sQF7HEzLJjCakJYypX9RNoag7wT7p+iQwyS8yrrQX3M7cgQa8k9
Jeux+e4zwGwxMhsKIqpWYAvHP911xPvhnXLN+b5DSLlH4LUBuRAb+vYzBhjFcvCkOvfJSlsOu/R+
kDKPB7Y8icWCNPoJCS53j3iCOEIGw2Q3k3XLMsKvopn4LhsaGC744IBWlHTvYk+QMLGVBJSILHaW
rLjnk3H43b3jMxeZzHi/i9wVqCjo3XnM2iLrHK2LCzcfwoUSFy72g797gRFAPAi2EHA6SFuOgAIq
DoVFlpEJqafnCIv53VI/MISb5TcEJUE4yK5deHSqJzwsUjEgfJOmss5L2t2tFobtVeY5PPvjOdY7
3/tcG+eejLiAC99sc5/j3mot57hvfx3e7maDKW9oljV4hpq5GP8iup0ZmVkMVQHCxvmkEEWpC8QZ
uyzYtNQZBYrmHuS9oiS9XfozJYP49LiaCnTiO7Xj1V6TiO1ysNyMyWMt0HK1dU+M2Gft5tyqevxC
mM4d/OgOO/VZXsVIiOWQtuijWR3Fj8Y7CAJoOE/QuKtIsnr9/7vbdFyIlr1V/b+iN2ciYcvb/XDj
nS1ec/py1CaVpLZSgJg3kDzRPi8xtFEeaYLNFDxjr7+6zBG3wIbCdBoNr1V4CPrTjXnAOy7yMn7d
PgvQ0KiuolDHzLzAFcuZzpyfcMuEFuUsmcHev0IJeFZPi7Zl5yK5H1PUR0bFdRk7d9slP4g2tZUW
yry1QyTLiTAEUQ9s96Q+Y2m5WqKDlly1uSeazfyPL1oSApOV6L9xoSPzMvqEmW5T328QizEFBUqk
8L44yQ7k2+7Y1RU4ls7DvmMJ2Slom/mUODJw3WDJUT1TbY/6N3P4BNeyscMRQVFE4Z5tNbDNwCJV
SveT4WIvQ4Rdy/Kc6atUTNUNKdNqypvKQbJZ647UU4pbaoAt1cWBafOFbra+yuGhPidoArPrSqnp
p1TPKrwOcQacA0GQerDd4W8p5vwjgscm8gqFQBC2SDTZ9BLz/PngFLpY/qMqlnLvKdt7v5MxIVOw
Yr9KT8s6HFB7XLgNhFBur5NfsW3U78cIrOgNANmwdetw0soh+Bz1D4v1MN+4mjZBJKf0asMjZb6j
tCvSxHngNLqETcVjddYKmvhLi8+WOox1CoV/8ryMpiD0h/JN/n4PcQJV3sB0pz5ig5OceHtwOSZF
kVFyGzp731tRcPrJriZmEKitAYYr39D0cke2jNZ9H+qrs9q6wifswmHaaY1wg4YkwbEfiEO9MnaR
H5XFXap2GsnI5rNxK1p8RX4UXSa/aLTk/qabIHq33bQXJceqaTjHreOI8J6TF6mboJlf89KliXvm
9wnkxfWsWODwOef0WN1gR+1HwZ+MepMc72gMQo7208EGf5vYnkIA/xbH1eR/e3vYE5fFBSRBdFTS
X427iS0c2LdHQNTEC0FsGeLftgBlChvSLWEcBgpQcx4KLu6ebFoEYrir74riPuoDEAhWWQVph2QJ
iv56rruFk3VgjsY2XTKE79DrVxLnGKwsOvmj9QQH7j9xb8a+Aysrbn8U8xCV0JAB+kRVr4mShrYT
ya53tZbHKg0dObPlv+D4RAlJrCdSUoFgYDGYI4kT4xtiMr/AtIWRjNcBOwzACr4j5jpK/ul+hXLY
6mRxq6HikuVZagAfLu+qqxG+M/KDptjeG+s3mXkeiQcuydkw0cP7VOfPj2TZ8Oc2+/pVsRATMDHd
wUCv4+LUR35jLMMbAsXIGreKJMQs9h7rH1Z5AepN6YFNLzI2AdEEj5p8yXe9/Jqp3Unk+R1c7mfe
78DXp2Rgo3jWzHeQncTSqJojXzOMxbblVHWHTn8oF2VSuMXHykch1pehfIh5A/+sEmrZaBbaSXo0
F6RtFR783XFYgltITjSQG85WjyND9Oo4EG7oRsGrhcDSdZyzk8CXjstQpdjcHj3dzrk5Q3sZwe9T
N8XfxzG/7eo32w0ARfHNzphmC53U7R9PL3uhB6qzP84od2aJNCWf2QGVBfENHTUQNI/OoPnwD9Am
D86O4dz6hJmIChSAMEqmmR0pLQB4bdF2Rveb78eFLBnm5ypa8MB/W9rDbg95c4yL/maRPm7DytL8
gCwFjQRRurh6eUIOKaCnOeHObxCNkM/RyQpxwKf/7GQygwqLbZ8drBm0n4t12BWzML0BQca6brdH
ZPoVASXut77Gly5p9NZV7x7NaWoavNioqlJEtf/v1MJGteMw3OugCEBXYCeAJh3/VVsZYRTscOLC
iIn+1cBBTG6b4Wvji/bh5u+iE37BrUSNnEL5bA3qFmdrkKgExzyUQqfgHIDth96H6MQkIxqxhbyM
AYAJG+52ne0aAspSC+8ICut1HjpMZXjN9450Os8pxErCmeERNBkZcfrLZuAX+RwGsdzR53OZ/vBm
6dd8aPGChpwTEfAGV3wqBmv/uz9jJRiLnd9syCKvjaWuJJ+Muwwd595A86SftL9tBfrqh3fMz0Rg
UNGCwWkPAq5i7ffpArr7e9oD0cD9kyt3EHERxPphxw/TM8mrFaLKezZL3V8zCJbGnnMCuRm4dB8t
byCvOduMmld/qzHBCoWgdb11jxNbKJIstpGL8vywWn7EQ+9GscKC12uGSnS+5iQbsnzDQtQAesJW
kPtsi2kj0LpnxS4tQR0RRNBSyG/kfWRKYjcmwLIywvqCrow5PQ/GgGVmvqvTFYFNJLj2+hi+J6bV
hYhp07mo7tFrKbZl+1og36He4VUNxcis5CPTBbCq2nmQF717G4ELV/OEfukJ//RnIP7utx6lDi9I
p1XQKF98ICIDDsyd1NHTGNo7y28yfgVxxGfXXrR2NYdo1BDaH0SdJQSpCAS9d9XvtttxxrrELopx
5GXQjXplBNPHGQ+z0MqkJHSY4CHVWwe4zToFcQAweBdWaqcm0Ex+SSSIxsuMHqKe1zxGuc/y75WH
Sj8vdA94ABqNxxw8btnQPOjHMZhGJXl5LxPnFtjpQumFUoP+BhZYI+7ORrDHJlCxR0BFS7lPbDum
wmfAQd9q8VxySsKmfqtKqVN3qU5neczy6Z+xliB2lZdPL5YHnBVxDbMJ20egws+F7HWPvNcrjML8
NOpyAT6R0YWVL2V34tdfeO6Zlau+nX3hIw1ZrCaQfiCY1F8VIUSq2QOIkbLvJgTqzMpAO4kbPbSE
7tR3C9PSgDej2X7SqtM3m4L4wRIJuYHPsnhtxryMd+3dZYVXZpk4/00KWYRbgwz3WGEeC0dWo+LF
3KUL9fixoAtpsBUGtxbG9F9FMMixMxnZV0Jmw1Z6ZOPz/d0+RvXuxp2qlEAlb4FFV11K7rqPe9Vt
ix+EV6kfW5F1LRoVDSoxK7puqTYcpUUijME0nVIqAz5Sjztyu9MmWCaWcOzrc1Q0Wz/xO/UYOnHL
f4Yh44+w4v3dlDpo/09c/yMRgGa5fkigsg1Tet3oEbNuGwe6hyCwStVSsg4rZ4dqLxmLiLG/ad0I
wBozGbZCtmyOmPmzJLyQkD5kprXAS3owZ54tOVtE0TYUkhf2Odr4oEPfZggRs2FrvHHgTM+gT0yu
ZvGCkSn0YlDgh7xQu3o6S6WKMWRNOhEw/iJtflYZcV8LuJlxBbKfOGQ861PSTP5fVMpBxFx5I+Rj
n5o1A3Ijrg5TAa361gsUVtmQD8a4MOTVqj0HvRMDB61JcLS706K2JT4I9fhlsNU3kEAOGXzMgSV4
wMSLe4zYUg/Qu00jhX4DRyxTdOJSd5mJ4mcc2DATx+9k8PciyYCW7cxLY+v/mKfxHfUgp0hXY92J
KxHDZDD7V69naejxBaCAaOfx6zxsxIj4JCG9FLkiaKynMsR5ovRaCuT3r7LiGdMJoelw3fo3CQXe
V+OCjJDEAMCp7MAc/EJIv6kLYAFUPtGZ9PpuIDQDze1xJfwHupbYVbt36YgtUkGhses+XBtxqxu6
UUrLfal5sIchvSOmjbJoaWPPJTUlfMUdCde8mxa/3WFZgAOwtR5SGojIsDkUHpyX8f1sxCaRpNwK
u1pFrZa6RFmHkAT6SUqAVXXS3Bivu4oZE+1FvIdSQHkEElFF4asOXZXow5km9zgpVk97QCABzxAk
hsu71Adv9UHUt5zZ6Nx9ewz8gYg0YX+Vcau1DtaSubMEM3okSRziwwfU/aiV9McC4tF+LArSSHF0
7IEj0Vn6jpDXEHQ0/4zmQw6MNgXem5lwagsJ2+GsLoblSo/pNPmkkpX5tV8AyZTDKKgegkAMN1Lv
nyXpHrnB9yBJgePbX36hKITNYWCVlxvdErRLzvNRvDfKMejj7nnh5tV/y1WPXvH4c8xihozVuw9M
SHD64yWlfaYpB4N4NAjIjD50HAEfXQPRC6fHH8IRqj+6uSprE8OJoQmYFueOp7Z36oSst9Kr5QUX
khHg82GZgr53gXVVQglagjbZ7N5qHXzvzOaFcI+UCwdz4ddcT8vRlnwdpyB5S/Y3vsIqNipz6TUW
/j3+AFeA0AmEoK7qZZntZidSqV2ZV5yPP5L39+FsK6C25j1L8yfdGnTLfG/6tcTLsbHP0klt3UlA
R5bhPGwKD3+5jOMGqUmmnrkRWvOu8KwaHXEQtbeTKxFZQRjQvNyPJtNDvyeLOAJI6OVCZ0C67j6m
skG6B7PfTSo6an9JVB5kwD3bN0vnJDIdQTj7G86NMU4G3sIUbIoiHCmZRzH0Z4+NObNr7auJjZ4S
tFX+VqNpUgUNwF30amE++dv/NnK2m+yf9cII+UqzjEIwMcQnNTs1Bg73LTtwUHSmvlXhuHyL4qiM
Cs60V06HPSCKaH4zCP7uut8q34d26+DkQ39HNNxt2xo90nf77KcGVpBt30N1Nm2J4IFaf8g4oKTr
6eFfXqLGs6eTgqZzo2j11IfWpd6wIqqNSxKQ6yV/prGhxC/qa2divd40klvgQyktvcuqBfNgU2XR
UQ35I6iSNULWFww6oXeIP//Ian3HmwEl08sJpp/WYyXtsSDtYzSL5RaPsI3SSVY12B0pBofPC0ii
7tKE0NMCGHPrzlKFfYy8ZP3aXDd3GxM0/mTatmFQwv1mUoy8BgDrDutZDZ1smTvfxd6ricq68U11
k3atEXNp+gWE3zBfGgWLFD9m99Yi9qKChzeM5xDM6Zq2HKLfPuxJclv0hKZhFHc6WkonJc1LQwJz
ddT036ZWdHpmc7LcLUIvb16j1krO5L8HKWOmT6XXoxXfbwTOWPHKt91JADpQX0KZA82PDs4k56dc
MIxzqMPLyqh2KXfDXZX127K66odUGGrGUcmvAjoRWGmXcr8guGBVJckEhaeT8x//kHMLxm+UWz/3
Yl/DpOAHyXcgy2yrKArpIzSvf0AEMSmMLXlH7geZW+S0aMuPE0X04doQENco1WJ7+KmQ1CV+jc7V
q1NmHA7I/sJfJDyBmFR8hC4hoNxv5x5027XXkd0u2z4kVaOQewrJ3wiMS8qGqWSnMyT/5cbL02Qs
5cK6vllW4SCgK1Ruwb9Ft0CcnGeWH/vPtiUzxT3LEUSVSuj94VtYGcWfNrLxzXMdtu19wk1KSz5P
y8TL6mE01usQSsGxJ8KxrRlyvBScIJ5Ju6hAN1Gd8hUw4lKccIEAy02HfkRbneaPRZtpXS3yEcpJ
jaLfimkbfBv+jCC5iJZgsLA64ECze/gMgMwMblt1FWmfzEN2JSrlRjfjtkfzOxSibJDwvp3LbtgJ
8/VOJ8jne5ahcz10ZjiOePVzkcuC+jvxqJhCqZp+n3v9TI3kfNv2Ft5p5ESuvM+qZfRHmAMdq8Id
BAdVhokcgZVXErr4s7rppNU2kxBDPxS4bNrcyemZThM3NSJoE24VVrPfcDJvKEEdylGXHTV19vi0
/+5wHEoc4rj25pEmm740/t18rV9iQkzc37/e8fczBjF7lT/iLxGJArqTWwHva7mcHwB2qkRINWNI
WClrcmmnmL7lrf/jSfskxN/Khp4/ARDb5Ct2I+Lq1eW9VVxMceJRvZY2GVTK07XZOPk3W6xUQP0X
6s10ztT98CA1I7C9iahzlcrwjjkFuopQS9IDrMo5llrsW8gPFg/aCtrxqN4bWwlIRU9Red0i/p3E
PRCL6ayTLEauiJhmnYdyknl+gHcfbSPG4unoMykw2yI5lwM9dT5VIH6B5BxfC0ESgP1SNL/+trdH
6PrgjusRt4ib+FrH4j0S+Q2mBnePX46Z68qS350kg8w0WZR2TOOaO0eZ1Qj2iaXfylt70DzcrL/l
OrtvKCjH9Awf4AB/MoyyqTfDY0qsD6veelFRU40gRckb5YG2AGUzk8Atb9RaGyvxVBAiW43Zv4fH
wD4zmvWPrLYEiXoVYClu2/R48Ui/zeLPPlh0+cv7ll9wD/s8Ya4I6CuLFbDMg1kIlNRiSPwQl266
ws5e7SacYwjmfJttMmUX2YXBnhCbcwkrhP8Jboecztf8F/6K+m/rorfax2GZzMEXlPlYFnDyMAQP
X+4xzLcu1kTeiPx5OOkjfxEDss77lkpg01vpjjN1yj6mtjyt13iO5DCNY9KBiDz92cBb397/lHDy
OJVH9paiOc1uUxZRrZiy7dhPj6rS0OtpN7/FTeGXjJV7VAUbjS09E1OC/8KQjh1xg+JdnOprYgHz
FiDMrXosL/8AlcIfimwxcVXWEjp+E8n95KohxhgvNk5KpnxOdKqQX1NHyUlwI2qKTo9eRDhSbqct
yZfo7dtRO63ROT98ZdnzCs/mcLvlAXSO/QySk/SSZaPQlKPcgsyUOvsgG+7MwKDiju1nBb9fQXON
MDwYTdfAVhI67e8Unq+d3K8Kb9iqkiX/LK2kwVio+PcaJ2FCvGGnHQ3FkByqvdtTvTElCvDhtfxr
4shhWqFSzui7wV6vISa2C9fnmx/yBAjw7isPiikD4B9hTbprpAoT7imUu7VqnpBEyBlWAxoDygPU
OodivaLUyVA0UKt24LsyYywtrmWbwTdx1TtC4wwsomNF7L6pGifq3SJnX7Jgz0VMGbEe0dM0OMUF
gXQ5/JYTFsm0h6jR7N7dbVAWjll7NvfLS1TEKfl1m4qsH0AX0MXe+ha4/CQOQNIr4mUwNCK5puyr
lthfGZ4Z+f+3nXaiSArzjuPy/3XLTkBTNysLuTZdLcVnIOebnl6pUbJitZKoxoVzWdprJ/1rWtFD
jDYgM/g4avte6XT0gVguWf9Fl3sacHAh5tXW5HdDB7cpy3IM10+D5VgpJv+cl4yUg9Ayc/YeLGc9
xztAEJaDwygIKuwxIqOPKJuvhT9jiCMvdC51/ncVDAYsADBpCt0PUi4DU+WDdQPlA49mkPZRPeCs
m/hhAR3cQuardjg3bnurWSURJPwjDf6A03VCpiIxcTBpK4L/cOK4mOrDSKTRAQbJ3yDNOQYpX5hD
EOVGAAM14ux6BDdbcIad0HF6TBp56cXu2a+raEPtqEaWpn6mVyizvJQfWC8EV1m6Yk8NyokVE73e
VpJNhnngNWYKvgY2avopR0fa6t/TuoTVnTrtAOm5wgH+N4C8SrE8FWm6cyukA87v7byRIeA1dCAV
sNv+M4hk0HWcG/FV9D6S50Ms8y1d2LTr3cZc+I3R1kWcf71dosdQkMd6IUBTYhRwejYMrIoQe5M/
nHzbPJ8Cmh8j4mxT/KBq4xvNERXqTaDeqzEi1hEHGRlfOONR2Kh0izXeFBcCAZyKaCW9973j0ciE
1eGAeEF2mBYjt9Ki02vjWFdlXQ5kciRWx3VP7ZLAM6OKW6x7kfWKL3oDEi1y0snwvQDtiCf3d0Ps
3oVdb3pN7ARTyh1+CNZ1yurJCEMa8Z5rSS+yycBgO6o92KTYmvmCH/8RIdyoT7B6GDUo0jtyU6Cd
H/9GECVVS3W6ZqD8UIIJdmyUZwhMhL6T6gb+BIVmSjJJfUwtK/UlyAjTZRpQuAVh+njBwCkdEhQ2
CbOAWVA5jFOvNEIA51jBUw3q3VgXQN7oi6YLuKwb0A5It4vwhFUQExmkkyZI0WKfA0pIFTIIOUYK
2n3uRmN+c+4E9kUpt3QuFp2yqKKCYkfvT2feiL+CKdJ70f3G/9IkVM43svdK4ELJTJuFqdS77RqT
iN4gbKACjmR+zpGQmRY59wpzevCjgvCtTehSUkw1nYVCVbiSenROVNygDCwekQEusoWMHBm1RVHh
A/6qOZKJEJMs9MR2Vwn1fSvjfFAlmfWOlQesV+qwAePjX9zoCOU96Exk/v07YQv5hCWkgiEfBV6l
y2NSriSb8zgReVVxZe1hPrUnqD/xcsFtf/uKMc5ea8J5SlfkvMJcWsnALIB91kbsunNqGZCXOpBU
bgLqU7ho5DW8mlh3nlOt5dPErriunKzYWZp8tJt/0pNjYSstdOTOKqZq1yTCTOsbyjFFYKKRfPpK
MHrutffW7gXI+MQ3QDQ8rjp5LPp92gOdRaOklVrpvkLpKF02Q/Rz9XHt0RU9Oi+j8XlNuvggjjo7
NuD8ujnpdYqMcpHsBoH+eOGBnlTXP4NraFpElwbV0qzFq1JxIoXhQJbqV05V35c2oQowwypfQ0zR
/YzoSmCmv/9JQAMix068G7SYYMeHraVZNui82vQtjzboV37lBsLLT88pjrXeFNP0LzNavwBm/nug
z7dh/ugFxX4fg7qtlkV3G3TJJ5uFiOr4navwuPZXaIG9VHOgKCBDE7Cdo5wf4hg0ZP58SZyF4H//
5H3zTzehaFPB55Ke0CaswSWM5qmljDLqJsm98tZj7x51kH76dzq8e6R8wVBr/UKQ79aNKSvf3jbM
tjQ87O9rlsf9coypB/RGHq2Y63oBA159PDOpBIDcBl7Vl0pndmfYbfIr17G8J36lt0q264PuQ1qu
Jcuxwm8Tk56tBrVTcFAWH7qVPG/6pXj4LJsQcVtY4uV45GliUWSZ91aPtvZ8Ud0wF8mAJK8TP4cT
IpIMyceyQV/fcDj+JQAuwhZ7yx7lI3NDCoeKM49tKykiXA4YVPb+T6zpq+yJF5UdMy+CLEf5tWv9
/bZVMXy2B12A9KjrqeGNMWfTwEjh+LyoRv09cQi/ZdfRFWoXMMLgcEs+0mLFVc4XVutimCRLCb7y
fWzufQtb7sEHPf7BZ9KcrpEBPNZPfKYSmJH4LJubNEeTO6ObXbBsClc/LRYyPMn7FKJRx0/vIZTA
AkQxj2gzu2wYlg6nyRqdDeZpAx/tZGGapeSJPzsWVRCy3pDgarCAlL7GMZ/eK7n+ZeVdclu9OLm0
JBuDcpchEdC32Es8PF2BBgtIXBqHnypY9+IbuJWqdgW8Dg6yWyle6W+WdL3RXUu9Xn4TK9D97whH
n7YxiHJA6Ob+ebFQlxzdf5q9k9gLF6YYJEGXbYj/xXq4HW4l8iFyObRH3/4JS16SHTxtbnhPn3MT
62YZGXUnYO+IhkRJlzvMIXuZR/lJYFxpPmyB1iZ6ORoiAPnX4Afm4/4C6Q3SFj2eU1lKQvmb6N3F
Tp1gbBN30cVXeIyQ1pntMZqPktVA0/fdJzEJdKkgyeEm2t6X3WuxaC0JpScBKrNZROUSVa9tMkBp
Qy/VoLpvrA3NTL79Fv0sS4ioPGybSF4VEb88iVxm36OBxtAUj80kRTgsMQGH2Z17s7WApVHYl4qy
t1Cx+rFfuRhBV+wy882I7PwCDRklI5oap9aJfqNcgWxoj0Y9GuZw4Dc+mu1TcJzdME24JyxLzPuv
lXGeYxZ2O2ySuMpAnGglZ588TecMDou5ThvALrTm3Ymn7OfX4y+qcxXS0LED+At7y5FFY0YScmc3
gLvn3RrSwEVHNS6L0pxL/me5Iq5TApNrxY5eT26AsAUf3WkiUTsiPVQPBQUU6OOEpwmALJuLxGlS
R4G75jZvukPH9lTTFX4JqTNvnnV2lkkUQjtY5BHTkzS9CKy6PgDdXKd1sRCIcad4/XZCFIZZfE8j
yjjHIPwji5zY8KJvtyh+5rXCRPuw5+Ma9UrxrX/joh4k0b+BoKg8aOAdVfatPp2vmfMDgoQWjfFh
gHEGXa/4RUpsTGhcYg+2LHWzsv3VtU2SmroS90gbNs2No04ppszDVIoD3j+IyBiM/T3azhF6jMfH
Lue4VX7WzCto5ck7bcqg+S1PlW0stdIYaeRu2qQ4g6nUjyDrYtSjBdE8NcgG+XmtyH9TpL1eUOlG
DBwoyN809tAo9vpMIt/oDNe8nvHJhmHBjyNFz3yLmRfHVBoBQ6ht+u9nZiLdP2rUtCHH6Es1yJkc
Fl6nwPk+kfU1QPhjtwTo0kb9evnPacV35rfi6bC2OqMNCgVb5lkgHdPmCvPXwbECl5ryiToGmd9V
sN8C2MURuWHWZ79hMK5jE6QR2nDq9SIre0nAxDMjchmYRCGQ52eEVkAX9o0cNLOK931GuDNYibJN
E8pDCVAN8QrvMJOWjn+bkaS/0J2te+ldopJCM/FYrdoagLCEOCESMrP+2q3+PAuNcrBzEjTIMQ92
4COSSk7nRPj06nF/EmZZLTxu1PVUwK4ntIeE1shGyXvGGHFAWvnzuBfvF4PCvp6gpRu568qmFQYx
Ub1YGpe+Z8YSmN2pBmaeSa9v8HhT3BdStCorGR0D28tjEfol0SsbkalwfgMI273UjtgslcHYfYa5
EFUP8BXzWK4mAMX3hB8JPfQB3nCBScufgrfdlYeHV2VhT/Sh1QMv9bllX5wLjtbJgQ6kQdUstyjD
5S1e4RYmn2lbNrSX8oR/6SCS9NaNLphOuFXbgLfXXc40IRVFX/gHh5a/9eISMBlxh6J+pRpAFueD
D/8PUrI8WpwM5MPlnDiBpYIXdFG7zP1RMelNuvpceJBSysyMdgfGEng83y00RDAvFfkybaTwniM4
dQrdnGwcaun6hVfMrQNh1iuBu7z05fEOtSQcKUjiDoENCCUU/LMPzIaIgs2BaP8YY9sB4iyYNz1/
/Q0ukO621YXXjdPZsi24lNbcmeWAOpQhpfPjT56Cf4ffPSPR+DTBNVs9NzTWGY+cbi1+D3QSup9N
K6cwhW+De9w75ZdlSlyUbeiUTV0dYZ21/USVFrJ1ijgLcDroALSRteG00zxs9w/Z8JYW94Bk9gBT
sUZoHjsUc5mh74dApNwZCPpw5hML4TpbK2vAqNGvlmxf784xJJFGOi313bmuSLnrKRHXKUIs7LH8
JT7P8YZ4Hz04tc44F18YC/rHz7YWMBrAHUhqq+46uUat8XQgoZYFt1TkDHLo6TGlfmWvTHcf7Ct8
S1dPoFuMKu3/MYS6dWnNfexvus+8n2P4QiluoWRRBj2EsmT/yKCyj1OlmDx2u6cAv7djKbmu1oD1
1GmIAQH4EF5dSCVHnYxhUavJ1YIhRFeMC/uBGrzmaargB6r1qcfVnGGCqgMe/yV38tR1RZWqGbSG
72DFqtBrSmzipWSncRaSpTss4YmERwr89lzhaI1+jqsLcQCaTefcmkvFtwrM2eZ83r9LohgyBpp/
hWN+kiXapfMtPksXGSV+orsK9nRgJwHgYiD72X+2rQas5brjBZnwkjHSk/9UPHoOuQL5QX4TihOY
NVr7BMIQQFrZ2ZLxWdLN6+uTpoC80igoscjBPUdTK0RiqtZQAnCj83VRO4+ftDKTikt5Yw0dFz3i
4y3pD+ArDgVrVwpAYWVxBSx0m4wRNJQSoRRKsDR8LFjqtLSnPX/TVHHsF5VatmQqHNmkNefrNLUt
e3/9fWRkN7OF7V4Eezv9gXC0JZIg/y6xV0UjBENnAmWXH+qo+sVib3mfON9rtl1NaXkeg+jVtEHD
eFsC2H2uymMRUQW/DkRZwIFLCPAftoKVagKNIyjl5R6ukbVl0kOBxTT9ktHW99HAnk/VRbd6hn36
k+EZMBUBBUaF8fzgP92UqtYtLaZwS8Laz4x5ciEbZjhtFb9c/6E+ZFXhT8VxxuIo6wqT4W1NR5kY
10iv21EMz2kzMk+8HlghB3OloDD9zAVI5m09mvP6g2feJA5m5fQXTzgGWYP3sZQXWXbaH/mRT9pX
Ku9z67I6ds465ESpcdyGKeHWJ4XknXVVDNxHELT9+K8WanvZ/LopjiD9nirp51l4wGx7ClKUMDTy
Pe9MFNDVs00bL89VuUIi1Ih+s2B9IJFBP5b95LmkRtPZ4Wz/DnIYo9wkP0ZP850J7utQbeXIcZS5
rml2iWt7eIaco4cEtAMDptH9lzvX8CgkV7j+oI6zgWIHWabhF4lgPC2HIz8muQ162GN/SD24NOmb
aII854SUWNFMB6jRqe02DkmC941CSyEjX3Z6nyGxjwq0B2fzhSpZrdkFF4Mqh8zQb3FMoH0yXwIu
cqOlRk0/6wgxHDkT8Y3Tzc0oYCpZB1ibx5JLEfWLye7zDNPn7ebxZT59JUXvX/jZDH90P/IqhXeM
TEB2HfcOznhc6PCQgZI2aebuk/d6GJ2lRp8s45vvoJ2rdEg+I0h4G/G/nJkxnQJ+nmQNuI650kB+
UUv6kGgQKh8dr/XzAHmpbC2FMqmx1pznBCxZFisM6J+6EOm1c/b8vGgafVEyEnPNj54uMerS7qRC
3/4lEgP9i8FHogg8gZnwoKBCrP0x1OMiGfdxMjY+C0YFq1jHJ98wD/MrrCagBXOrZb5gmgtmHcZl
Fmz7Rw8Bq8POpc2Y+Ifu6UdBhj+wjwcH8WEH0S2rQQPpwOjPz93aP4UuEe5FZBuLPDlLlVLg6wTB
qEbZoS7h41D6mE+x60bEdCB9+GTpdJA/ve9kN2Rbu6gSvxpR1CzNgR1h4quuYsDrGa4ffhw+hK4X
ow70rn59gACXW4UT6pxyskv7gR6mz1dhnLfoDtUw6Ymbmpz/6bx12SN94rpOoQlkyxsjWmXy1t1C
rIF3lknp+9YTqV4vvFLTuuPVXGUrjg6mNr16q0HmBIAjIfVLRPR4dlGIprzjBwToPkZiFE9R/8Xb
OTlz3NOeP6shKpEDZxiLWD12jBx20iBY+iiYg1wbsS/avNuDjHMFGiPPkOtbVPHZiZ8Z29tRZQW9
DCYbh3jglQSogPF/BCYez7TVOEZXuT3MrjSkUCuPvrAucQJQOdKkXOgnO3qV793+UsjIzVBSRWhy
2Be42+heeWDfHwKBR+uA2V5BXLHU8DjTovAYOe/3SB/ukB62ZXmAdCR/uyl3dWtTN06dCNCd44Lv
AA6ZbZLZ5d+gzoIMFnP/yNa9vFXVPA4sq8vuk40tXDG5rxJQn1i5nTTPPTmCz3HQrrWPhQiC/jI0
Y4Xn4lBiFarjmK0cjsHLieW9xihk8jiDLBNahotZsuHBvRpvQCM/GQ985KX2DaFveTwfcSsfy+zz
cved+SkkiyHzM+HceD8VDnt5rkKU6JiV3dS2MgZUvP9znR74d0uDM9XiJk3DU5a7KfKM5JUMjLIT
luWU1Q3j/R0DE1OgCSPPa991pPP55sZzKaRuL5c4fmnAH91ulULhogID/E1jcv+CC26hhYIgnjUU
Vf47krI4Yqv1ZZLNG2vmDuuzXhzngLOEW9qsylUrJT6TnPHVAxsI1m+PwOihSXuDvzJlw2YyhWO/
nnCbOiHLPbJqxdg7NHPS7+hmoOasmVIEkrd80jgNDDGNZz1p5H5ICREZzT1UIunGWTjPYULL7xhz
5Bc2R6MYTWhestqH50Je2iHLvkJ6PDPuTxiFEtQX4WHSdFW6qs+IziIgtyxLQGuqxjXaYpQW1feP
pPE/pu0bokTzmrMTPokqjTdAy3GUGUdo7MLK0CQrNnVOc3c5pTLztu7C3Kn5tcniJVPEI/rJEr4V
urNG7GzWAC8VmQOCaCD0NmsqP1izNJtndk05+RTv34BEa9PMhaBnkeXrbV7gh6HW/vK6/wxXfXzy
mP6ynvvwPd6U/hChYeklLGw6mQkX+7r8B8BGMiCOHnSbA9XxUt67nyBQgHXPSl2pP688hzyF76ZW
5eyHIQJpTzfqvINMW0E/8pdrIKSgIGp+9xW1Am0aiJHDSwXDNc+L5wzoK/V8kXxIDWkxsO9l6bve
AaR/jp6ZxcqOSpigHpeznbJyUY7fFVN5FHk9UslZXz1Kc2d9STZyiqXh4JGXT2cM3edc1V+Msniz
b5KwM70YTks0gW2KRxjxHeKFR9PcjFdkiNHwbRNhkCHIlMdNnAH/A4k4yD0z94WS/gco3MJfWazz
60wTaGrfV73DVQZlsxFflWnIoSRFHBhdo1Aq7RQoyp+Zd8gkDmSU5z3PHGGcoNuSVkWyboWt8wV5
Z41ay/lYWVqTsMfyccHi+Lbksr9zJdUGykhEwP2INsYLGJRgZEPF2xh5VS/soGGeAYacAWDNOzFY
cI6IviuD/ruI2V87bbrSvubKEr0R5sn4E8hZxRmLstRT1zI/aPp9kAIQB0dAef3lS6FDH6f0eow3
TZLIisqVf8Z9ALtf1Oyv2tsHPwgv2+devxeokeT6YTrV4LWo/ZPaFS3YOxcsJ1JrkH9DkhQOlHVt
GWM2ymg8+0TDhCeU1nSYkFry8zvRkytp6RAGAL7SZx+qvjjY+DAzm1e6cxfzPRnZ4zpuEP5ipNqk
06Bs6nwJjbjoq51Vphz6VG5571ywvjMESe3weCiVqYVT1JA8UBWhZNsbD0Vfc7d/IkGblgDY6/Qi
8iBXqNw/lk4RBcsOhZQQItQ+l3mX/w4srzuh6QEe9zk5bCZJuE6jy9k2BRJFBNWRKPZE8cKrZTCm
Zwzf7wB8vfcabqw7rX646RtwVZrA1/oiDrfQrNKxPKbS0Zi18CG0cruedS7obtAd2GR3Lu7Ei0kf
g/TVKVgYoigspmiWMuFv0T6hXfiEUtLmTyXPEXPZcYp6QLyV17zRFFXizCZiZsxFREeVhIXWGnVx
qZBrl0VrUw6BKf9uYuP6y6tOPAFfiZpGx7VTfpAfHj62Xpuv0VzLTV2q0UEOdkpQFvtZV/s6AqJe
vqTwVdrrbaGi3M9SinU5JwBtb126GcS2PrJr1yyjDBDR1MNBLdXmXKHkA9EIEtBOm2/n0OHCmd6K
qCjvVOwAhglcoCFZQTIBtL3qop3qz27EygjNJduL5HX+XzWDTpcpoYD7Pzd9hfuzuVc0bVt+FKqA
80yypvKmTDxnlPKtCMTN5RgwOuSTEKlYFvuCWonzGuB226rn2dfVcr+Lw3zk7vmf9pcIRvpYGCSv
jYILs0kgKK+Kh6ZkizWH7kEG71PoCdosklM6wDaCXAJq21UclVA/z/3JtFL8Kk5i5odQ+L+rjf85
NDbKVtHi4eZiNt2VvffBhIqeg1sYiwvWbBJ2tJYR4fCJSkAcDk+rW0XWAIZZmf+b4aGuW9DE/bVk
Vgm4uUYGRepMRvQy8CYIKAaJkh3tlt8FY749xW74Lodm/kSVfdBk1Kjih7NgR/EXMfW/YBAVr2V8
lhwabQ+3MRmJehLOQo2Iaaw6Nw4AHlaD9VSS/TKvlazgzWL34x+p5FBWCEdO3KosYMdRqg4/kjPb
TpPtgHfyiLf4SUYt2AuiLQGCFhX/TEJHVAie0Y6yCm2iYEOj4nDINQJe0OIx1Qq2m8zbjvl7VER2
rk2+j6K+zXgaPIG0KjQZGmiG6M1ffP6xTgDGRadyxSQJCYBW/MBl4ZpcDAdC+hR0e+dN7M7YSlkG
ISZW2su7G++bADEVsuWmfSvrZDUQtjGIgAiLLKj0SwTF/DKRn+hTW1Lt1RPoJuaDcatBevtaDiUw
S3OwWxOVRpkiLwVqD7GXrt0Tn8pabasEOIH/6/XKRTBub1oxOnRQ4iU2buebF9CocK2IFuhrfbnc
WyRp214q6tcN9esDepNRutkYmI4t5GpUSPZSb4vMnGRDoQN4ZmBBd5ds1mVIIVv14l+yJd0uIWJK
aB+Cu8hngvcCDMGNU3mDM7Hn6+IoxUHzxR3w93333DMxAKFiQrb074l+QQFRjA2fDDCqvVk+hfOu
DGQ9u69wpiS7HiIv4HwrFVkjajP53P1iqFqohoY6RNSPRRy30Rbfmqp25Hd5wZmtFxDFkGIC2eJv
iyM4AfdkAxl3cvxvRqcfsp8WkhxmcsOME0BnZ76FioygMfIrlYjhFnXUQKnOXm7FuCcJythD1UCW
sBRpQLDQt5m2E8wO/upMA2hy7LLm4RYtXraUCd9fzXWiZPrl3jTxrcvuWZejq/HYvQVOEpcLRXus
6Ks4uWJY2Mg/NOfiFGPA2HkjU5XxL+LZzu8FWgD9gvbDFLyCGf83RBNZ2m8xKpRKyB6X7uelY22P
s8zKluhbVPALF7hMUmOhPZ+VDU1etb/m4lVbZ6epuPFBWEfB/edcxz5QxM0yfm19jX8eE8r/q91z
mUqUTuU3rzV/iVKk72MXMJWvj+CR3teq2m7E9Dc30a/tlAYgrZu85kf49qOk4ddRePcfHm2iDcKu
xKHyHbtvyBbgj89D5ECjCy0GQpBpHPO5ZmsXu0Sk07pq0AkNM437vqpXNZclrwfDY2fpalb03LRd
rGSFqwOOZ+U8BjLQXTU8OyjA2AEeDE1zpdcY7cUf5QqJsnziaDNkbZL/kvKY2emCsIE26GNNnDHE
dC6bThZvFk+fYEqaYkaY6Zv38fGyTxceZZ/rpnmoI1jvJ2aul6s4oVz0ems/PJTvAv64KXJ1C5Eu
78o6l6LrJyibDEvSbP/b19Gw9WtzpwkOj5iCbCVIp+iImScrfO3cuqWsmHP2jU9ENBNhvjBR4iKF
6+nPw5YZKqhDJS4kx16Z+rknAjHboMOt1QqdpQ6frxtudnqi3Htw1bhHiCcTBC9a5ox6tpUKM2W/
H1eRbz5f37zmzKgDksCOSuuHywUV7zOV6j2l+Eiqli0PwuW/dYUVn5uiHH7KtcJvyjsfkG4YSUnD
DWLX3nPFBNKTfqe5kWlOeUWPPq10ElFiqzUGBXl8TScJ+5n9X2oDbUzfiFoebHzOSYkcKEUtJ4u1
ZhaRF0Ul2GNLXx/DZ1ndn6ZkxB4CsTh4LskmL/cfyQC+0bFeP9UKHJ2y3/8nzdhIpZZTRLfxFeTB
bB7i972GpUgZsoWsYFdyCE0GVhq6LgolKcjhuzIoIThvbtQylxzzGIarCvgwIWeP5VpmvUvETY9Z
6dVSt2aY7w8DFafkJCSag0RBPQP52yvd8960EN1wQp+IgNTuXZ4uWB9LTBwpPueThEK5CWV2Nv9A
xn27TkXDgr/ZIW4mniTVPfodaSqoc+t90e89+eDzyglcoUcg3x9KjQnVXlUEV3yJsvV/RHgMeyXa
BePAJU6wZ9jZoX9Z/vCxzhxBX0cd+lFf0idsShO0xODo9XpG7sfY2+2R77IrAoaXY4opZy7BQJUl
IeEwNDCuQCIxDnh+t744JCscIYkhk2FOHB7U4blZQ8L0z3lUBFgZQa9CNXV1WHWIxpI2wc4jTc3D
sEbAqtRrL+7gOXsjR1/iXQ7yq3ghjKePQn3J30SfFPlZcAIJIkSNeiRK/rptp92pQuja+hBUJSOJ
X7DemTQX+7GdltQNaHcYi1bA9EgWEmDjHZF2KHrFo28j497BzO2X7Uh4D4bj7Hbr+PB07MSeuoYp
9rTxdd4D46s67WkIxKyuATNg6INVoAzqqV2LdZOQoXD8yQFY9Cn9RtopQpU1waVRMBBcvSPzFfha
q4IJfHBEVuLvayGIcYcR+vC+OkcnVGoUuDluhsxtsATzWqrMYB4hbwzRSk6pLHShRzhLyBYs9e5v
QLOFzpDrQN74mfd+Ic3Zj2dudgb2jiUOFps2kHzYNNfPnxc0IUdVap+UiMtr5ghvA0FEJQj+Cler
XdicnsIPHPqbVcY7kIZhxDqvg3Jtz1upd6CRPqzwpsyoieVTYY7CNJdGSa0lZnZ3nqy9X+F7YWT6
nFBEWDmaRc4Vl7omYoyvZQYm3LeVaQDfkWuAniq85For0sJovAqd9uwih4UhDAlzm8kJnva3a3KG
4AMWo/Zyc1WoVOw93ErsVGCOmPLHUW+GcZqqXVbtkC0tOjR6hYORVr78NKjFLVOIeMsrCYiXQ9/Y
v6dHsvz3n1dP+00JoSCfe00kYIWjQxcJVz4b9ffd1yjXIqTcjsrrLJDv/nqAUpNYXwku2MSg3s5q
ntiVFfC4HsX9m7FLACF7fr3QARuuN6eVcvXL0pzfwQk2fy7+EkXbFVl3O1LydGccQLTRayu/MQS0
yS5BKLwiTdKP9JeTG7olrBt3Y+62t/vEkeRj0IPfSfrxXrP/bXQQfVx1chaKl6JDtQxnpZUYOU9N
D1oq0nNRCTcGqxsRFwulLyKC4/1z2v50PGAQaao2Pxq7fi2RxSqSUAe00VyXptCobTm/nffcwx93
A09nq2+27whQ0H8o57LniCJEJqmYtcUlcaNfTPCOFipV2FQ+VR7z+yiaz3wE6I0aEtGHh+9wBrTO
/fSUxj8kxKD44tzbJmTwQ7U1OYMNe5GTJbWq+HnHTQAVju6vQHPrM5sXax0M+Xyzf6RGO5wiph0D
2XpjMHfsQ8p2lkOBjdsDhN3ZF+EPInPsLGf9XMVHYIhR1R8LxPEI32pCrpClUhB64uLPKIrnZ7LO
/4TmGdzEJCP+Plz3owv/51P+Y4X+WQbWFSSrlz52hQiA4rk5Qr4v4xUsxihHhR0MsajcxWMqi+QM
nWwJEwmPo44F2rD/4ztdHmabIOotB1VjxEbPoZH5Fu8c3uFvWFXTW30I3LX5JM7V4XkHQHMHqOmF
mXl2BVU74cTRk4n8I71jJ+sC9eTFdeqnwmM18x+iW1mOIIUENq0h8HZQfl8LkZsJPvSQUlR3jTbY
Kig8X5AzXRCJQK1jE/MraPwBlz91ZUQA9STOXp24KSyzm+ifAtHGUVL6p8O+z9kPRaFWYWRy4/rl
xGKP5hpe/PaGy1/m9ajc/85sNsKHljFtj4EGSLeN6iuid9USWx+GJJLOZeFBg9sJfooq4jhK/Y1M
T0Hp3wv6lo4udytYIdyDZwBdZlczn6zmPggXPcNmQoomk4UqNnG5KH33wjEKFINwFNg1Xdbyfx/6
gBn/cqZl9MGAT6JXIydyE24RyVoiv34LLKhq79fm/gROBBF20ODNkvZ20EMmoVCrMfdkTFJg3xMq
IokS/Gej5ElwUXSg7tJnEOpJG2vsGeK5AqzaIT5uCQwJrBjYoUFGAMln/dpN7cuywaNLu7QsGaX4
kLWRVdBD+cqzQi8RuhQf6gHtI0gkjb3nRCjtB6Cdkm18TCPonNIVmdfSl4VS7DPt473pwDsgHHK9
+wIERUnE3GEUdS4cj3/liGfvs+TATCBes8RHcZwRuDMO7wW3JIfBsr3MyrI5Lk5GWxqstd8b/sn9
3D2hL1+2CRLyZkiezF0Ltbta5djD4D/HtK7ec8wjzjkKY/an3AQ1Q3Tifhs0Izky1eb3/Go4iutX
AkIlBcEWxDDhYLTdebU3bRafeayNglqxBVHC3s/sJCLKE4lRzPlTA4EdBgTlPv5IZ0FJ+vcFKakT
w4vYJV2ZkiT1rZjBhG+KpEtGqrIUXkV0NedCGV0YunFCzrYpt4DPRNN8wB8hUUimq+27z/rTTvr4
2DoAUqqZ4oQjptIz7Y4GX4W6sLzuBjfPlX0vc+9IH3ZOiE4RFUW3sQLrYf1q7avJdqa6HOadjLjn
XN0CXWXSNmOo9gx8YHqZXuw6eIYULakdqzhaupAmfdMQ62LUa4xXsla6p5/hkrB4hcZjZ4FFjQiX
QEXfDQoQ1R14QrrzwTOB/Y75lYNemzqpDl2iYpZ1S1ew7YppmcOLhBmsU/18lRvypAUBjkbQM6Ar
Op2++w2VlT3GHvrfrv28oaTKRJvCNhFKLOuGXA5wslLJS7lSLPYsA6ebkNiGxVOObqMoOYuRVhPT
JsRQ7yQW+eGMRGkv6XQktA+OAtq5PmFtz7QpL4Tk6k3tNB90E9shffSUfz+osOf8TMDO3pW2D2dg
KEsVXMeAKMgMX53WGORzJvNu7gtn1MKUaDaX4hUFc1ZEemy03QupiGHP2YDH+e6jT8mdBADtu3N8
o+9U1ttDyFeaEVec5a5D/UXXn1pdiIlgUioqAgGlFfLkstGI2ZoRMW55SgLBaiuf4NQYPqk2qn4V
PSVhoWYT5dHbmiB8VSGdAuQX4wrSYOwtdKpppkxhjbx86xVQImvVPmtdft2/hx7rMmXj+vMCN8fe
RXoBqbey2yjKj0cCsfrJfTPEVjLhdbEP4Qsz5JY+c4UAfsQ/nGOpuBS/Hfk/wTT3GDwlDQU60WQe
+Od005V9sZixEcBogN9HSDBHVdYVr6swhY5TcxsJC04rujznMU6rIc3v8mgZvaPrllcAtn7q0wwQ
kikduTwP2kP/zJs2lNXkELpMIwTaiCz357s018fvPK/Ox6NsYGSuvrXeKpFITDT2ieXYAMTJMJMG
xvkl18a9v/ESeiuB6WbLqoKNtdMfedtb5zXkOl1LhqSIf3o3B19Oto2/uyaMceTzjr8gfybOZVTE
qY2M0ztpmVrB8tzaBTUeNl0V9LJUQLcXeaFQ15mWIKGWSfNpu9r9Ayk09IgxjzK6dki3D5eH4Heu
fNKU+eaAAD5IIxb/P+nSCyRDvwgNOevZYUab7ary0Il5sofeokC44og7ngh96eUmjOC4akicBjP/
crVo65sm7ilYEcbVwpZm/M2d9xGGGxwCD00LbTi1O2mWOsF4MBu8PgHuAPY2bjKbFMYUQEISVL6Z
hl5XRzFp4HM8ETwtNSGv26vqvCYJnFtuaYrTx6DfAo5O3LNoBRy0PHGMP5VGnVtF46h8apapARrI
i7M5/aurezfzsZFZJY0jkn1FCTWJrr3O4fFYuLAH/NvWRtLiofVMAqdc06J2xCbgGuTouZrpQDb+
XitboiJYuJ9ggpKnD1Hny5E2GJKYOaFs1h4fN+FC3bUBR2AyHMLT48ZBHGEi/kID8jux4GA09Rjz
GEg5MC4zWgRmqOxDNeIDrfA6Zg3TlzsL9hO97hNROS18decGtr9sZuS8DdPBX6kIc2ATy1112MZv
gZdqgf70tvRykuqZKfdQOLQC0LEWffMepguoU8AkaQD0y9I4Nyh8USBBNdhArB007z8sqxTYqnC0
D09GNrF6o4UEoy/BCiRtYXSJhiRm/MIuTI2ZO8NZN1NytRlUNw1JXROHwYxkwJ3h5RSmqor+oIQm
CSybHFwAih42fwbGBePSZ5oZND5N48Ptl1sAIAHLJQt/3gVG55s8v5KR1JZur6Ae/mICcdhWGZiL
axi2L5rTMUBsJqVTl2es5P6VCNeLY+poBLGQjotKDWRY+m/x80fMD3RHRwRdIwJ1ARUP1ZdjbF26
UveNegOpW7ueWlAWhuEHojTmmZzc1mpxMPXXw3xTEZ0luP+vbSRShRvBD3vKWu8TB7fLZKL5EL74
oxEE1t/zmDD0XjDy5TCeicCixE7Y7YERfTqUwX7cWdZTfajKExgz7UZjv57Y4O0/LkbrYhd8tQXt
MmfLeN3MX31WgWKmZ/aYPyqgTrfk79+eo+O/PQjaJR8hNaZUWDALECj3XtmKbN5XjiiofmK/2vTA
njVjN+PrmIN2YkWFdMotsIhhZT20UATXzYRySNSQl+N+/qCR9W4LbLzbTh0yukfEEcqQWhf9PA15
1NOATBKjYDidwm+VWVWSwJ78CUqke24VAK1QI4hMqIiSY+EJnbNSkFDJ4XZySis+mf59Mc/y0Tfk
qqO4oqd99etzOq9WvzWQGxHjqOJF7iHc9OSKAwlQWjgok03lJs7pw3qkR5h0NdXbfO9VxeLQAiF4
21BiiQqYLQ0ETgr5LWgtiFkWz+900u98bsig3TAnBe23ZO+XkGnaE4HsTKiYspCtOOBCV8irL4nw
0AYvQnWAzSZ/SMIKSHZB6Y2C4Dftq93ySNu1hqWZQA3nxGS/kqyIpF4JDDWXR1he1kL4xDc46dfM
9FxcIzf+yUYk+1bionaMjTRl0h6rToO59y1wYB2aesS5iecwy1ksUBXEPfNaozoQvW836eWyVBDP
X6UXXl/VAU42qyehHt+rMy2h40dUDcY3wcJ8uFgKVI8/+Mfvmtkr8ehWk9fdp2ps5dYejhOW/7YO
+Z2c06tzddsOKkJI/ld6wjYOTnGqvJG1t+mmIPPFTAjZwkpkF6R0hHXIZRYvPvtwl2b6sMHvaeCM
c77AkqjTM9FwpNsItgBZ0E9hNXMITQmetnPB2WjsRXCsqM+Yd8tbwoeMssIlbrdbZGylNOda1X3D
oOORb+zyvhBFGXRfppaUH4wBdntSRKPuCB3+ps5c+O+dB9beWC2lKu6ZpIaY/E360Xue3bkfN0WI
fp+/i6JpTXHhZ4KpAclTKYTE4uVP1tPUc9KNv+tXASu5tlCWeYTsyEb714hXRGeTxvbsYkkaI/w/
bD7qgKaGA0yPNmqNRApPyB3bwKHFtQR7iiq3OfkM/C8dore7Zq8Io3ij1Yq+ATz6T3ejkhNG1Wow
P8gaM3+6d7yk0+QEiId8esr1HKYGMyyzVHJWh6ApfyaCgcIq2tzjaZblNdA7wt8kaHKNG7PyIdB6
N2daE7duuDXXsM9abcLxhePHpvxeN4/8UQC6GEIEIb8w+9MAy+YgBGArLV24YQJnHMO8e98peTcm
KYaxV1kQEIjcRqDcy11CbDZBS0TsgOg1pqaQjZQWDdaTuhov529JTH4Vy9+fMnPl7XhuvQDOsNOV
8RTEO9SqcyHvXKi4kwczd3PFIzVK47UbFZiCldNl+cpt0C5RUheP2MtdxsBY+vJe0i6wxBVmZU05
mTlScS279eoVQIPitcINoA+rGjAJCsi9vJpcCe1LvmbOQfCQrorHXvEKVlKXw+81zcRtoQ8HcpBI
Tiylbfn+UvU9c7n6+bDtyG6XzNNTOzEqwmSFM0xBrmS4uV4AWkfNTZoOtQe7XgcxHv7Pu89FbE+h
WEvXu5GxtgVmFwL3XS1bZ85lUxT3jAQ1O9ic1zwKDdr47RAEj5MIwa6CUxGxX00f+gFOr82aXLb0
mLPqh8lW+iQxIeN+1hkUl/L3Y9040pLymJcgZKk2+/JhISHE4yGQWja1MWi1lMv2rQ+C26+cNNwc
/bKnVaMRWID30D7Yuq0IpmjwiZgSRaiyAUYV/o+EtKo2rp7vw0C/YxtqoIwnBvfgZ0kV9lj+EvH3
BfqaZmUU5KBuyEI/lgi9Jhk/iNgod/UYdzMuNCzS323DQcfgBnkUQ5xe7toPyjlJpAV6cwKySX5e
7MEmrdO43age5RwLxyv8KersUnDIDxHVF/tcPuXTmy4H0QAWruLU0B0XC47qHQwt2WN4H3rnFfqx
Cj3L7WxWqMiL4LlbaKbkKJb3E9Tbijp2Q+e36Az1SqwGV1e84JiAJWQoiUweUvK78okpEFE8xOUB
0yHqZHSQGK6xTYK8mjlv3cVKHTIRdcegC2pftKWWynqXkZQNmB0cO7HB88JLCpiNek8wEqmIKJfK
OsV9e76GJUL2bqtJ8gj4Dbs1NVDWnVVkWCo4JALhTNbLGb4lQah8vb3DYZD2Wq10Uvq/4gyuYM8e
muYL0z4buyYvrDXYmd0BHsjE2C2GgyqQOXGqCdt47BUljvo95wRu6l8MXZ/kS/wWWq7Q5zoFSn8v
CPmyzdd76i+ZV4NVUOmCKoNJFpF92NlUjW6mP5Ym/fe7tJ732Y3xoOUop2isu0Aj7IvJ/ag8JAzu
LQC3nhx/Z4eQ4Is+e/LazrEsalU9xTSGAVArICLTCVJpXJtN+zMYCm2G1pPSgOQwh8375IkgjI9u
a9C6Q21wTjUI8dwFC2xhyyd7mvHH7PBIX7JROaqJ5dO3hyzLEvJu9O3B5pFZyiAM+2GgV2jJ40vB
2vSRQvBjnfRBT8AqoI5fHsNdvZvPQz5uGdZzsd3tKye1kq1MBJFwM9yjep26xH9IX0EpOJLwue4e
q5dZ+MK00wZgs11SP74ZuGSvt47HmijP1oL6zKzTy+P45k/ezuTg2iT6wbpcL81lr4J+YsDfYGxM
5FGvcm907s5c1C1gQyMEIPeDfQ6WlgYGE8tCtZAlV1/g+LyI0Y+zkPZ1Wb7x2Cq0I46grsGXoF/c
PoClcSRUOXvfvs2W7xCeRgTEIeV784soyzgB8AQtpLwpSizFHt0qZ+qF595GI0mvl6MNyBcflTHe
X0c3nj9excii/qAt76oTAIsFfAJjEKtzNi9Rwqc9M8VP6ayOxpvCW3ILWiI5ARDxllVQgyRT0ph4
q8XNtPdhAnWYkG47sENl/zwsvJScB0eyH0w9sa0/xpMMB6DjGI1ZHPMaQPdTKzBODrij+XSvlP4b
XUcN9l6YDWH274UbVWkJt8XnxnijYTuIhFqeLPmheLUCVfAOXYKS8TfrOeD+at69iiUAu+7/KiNI
DilNgS7wLlflDU5C0rSgkJl027zzaBy8PwiZd5X5pWAThbJLKldVKpAzuim0AT26KJSrXtN+g0F4
OvArmvBju1rbYIsdUx8zZ45p/TJNjGLa9jcZDJmANT2XQKExJNBZC9d8xSTcyOxfPTq1zkPO0sQb
E+VLQoGkHg9wZ+3BCuq2G1ij5MZNj7J5Soz8zyfl00vWgQyjlhX0jJiT9a4fjZi77x4H2xW9iJrc
yCacFDt/80SrKCVfUhCnCS1gtOrYq0DmfqHxgQi5zGxBfNEZinwQjxDR/LgJySPFandg9Oru3IZ0
Y9a4G5sHVOc/TqTuMZoNeMYqJie8BiRXyS/ONk+o8aBw0Cmr8zGHZJfNdybwjmvXmdfVNXBtKQjA
HevImHjW8TGdFJWptVGMO1+t4vE+QDRxEG+cEghXxjuq4FDzKihHueyA26cl3PuyPqtkMA5R5FrE
ITcpIkMfufrtyJiADicqaY3EpH1YAPyoEfMTEbaz1w4HDyWjqEWuNVz6eyfpTe7V19eXpiowjQck
mXNQAHPmDpbAo7HLi7nkM2t2BJWXlJU2mrLJIn2TD2nXiU65UegVhh4GBDam4nPBjpcR50AqgI+4
0IaaElSyF+C1RvtKNOkJhcK2qCTXDovv5jk4kigj5F34tiUphrZX+ot/H/Cg0qY6/eXU0/iSBEY+
uZ0nML7p/hbRDAfpV02KKAtJ8eRfJASFnKQb2dh+DQQaSQN5JHcaH4iBcTCtj7lSX0TcvrKXVIiT
yt2MtpBsLCMS3wxWSoPIel8tAhojPXI2WNNbQyEjYzcypqPbyNoPH8VElbENVbc4x8DvecJ+qqoX
xmovJpaWyUrD2B7wZE/Cda2lh6mkA1Daj0JlXIZWfEdt0CawMcN31WZEBqH8SsiRwUAjZHMaIUpl
zU7iLPIJnjlJmA04H09IvuIfzqQsa62dBEIVzK2pw23nu54FMRK2AGFbiMfedysWhLHmDjT+JGx3
46oUm1gp0rG1digNNZLMd3NYNLEpEwiLpMghh5HJfFDVneAdFBz4Skoo6hXoanJ62zXf4CdoIQx6
GGlQRlBIIyT4XK+1cc4TUzPbdQ9W8vfZAdLRa5Ze+BbTX6Zny6j2UgRGAmlJNUZp4e6PrnkpXY0c
Y9yiiDFeAGrC8fXuocd0QA4H8fafW/qvXv/3zJu3Pk6s2VsBgsb1RF/F7Q/LuYtLCmGh6VZRCf8U
7hvoRUTizKBFUiIV/GV9wLnCss1AjKKQDJzhOsd+F4xKBlrlNT/Pj624nJgAbuP4joqnlO0dpLRl
LPzJRf8Yxrt8eiEKnFLy47Ir7cWnyIWG5eLgLOPdC6zcKu2M9BqSqGtdctuD3aiZeClf7HkwOfQE
pMGSfv5HmiMFACgvzMyY5gN9NLelqK8kTTOXk2jzGG9r2T2/TihB3v3j9jPeZHZhuheYbNDKhw9X
27Un69xx9LzxPPPgGWBwCYgO1ZS26sogODmz8l69f3gnjGudI/agD2YTMAx3d5HHO4rlKDiur7WS
5zeOZAFKI7rZrSBLq5/U3Udpvpog0PCe/3LFK5czjUVBfu4ibp2+TUK1xAg8ANK69UI6Ok++q+Sb
IAUOTRX0tFGVNsr55Mv8+WpKpOB/NNXe8ghIye4U1MgusLHkdG2y++u+m3QE6baC2CSn6AQVIzWY
4Paiz3mubD/GNosQvsDPNTqFruOPWaAYSj2zt+FQVz+5vDvWJI776EbmcpeTkciXS8DPuJuZhozY
iE6C4052FHI2NXiIwpeuDtGb0aHYLisZ4+Erj/Hd/DGS2mpj3nBxyQHi+1lBHcV8NO14bBzwL8A+
FftEPuBsm5HUXuzLmb41yLztYZ9KQ5IOUxi5S9cXIlKT/OgfyU476gT+kGuXM1yCMeL/GRtD6PMg
OKAMMoYL/7yTGcK0VXRGEl74nQPcyVNKaM2W4j3N62EjqZLff9mgDPmgHO+BtGIsrRhS4CZ2ShDT
PaimBC16B4e3cqdoBSiDAzlWxwVIZq5kZMksF4PbY2V7OCS/bY0Kz6J6Y9KWqyA7lIFI+DfenbkB
kY47wfeJqsOWOhykTVIwv3QXVCK9psCXQ+FqJWhAyHyvl3Iy9myFNOQNFvkAm68QrMdMocFqTC6y
gABlxkODfBCShZx+s0cUkuxu60DTdYihBClDmrTMNQI5pvGFx+utsWDNHfvewvkQLw+ZqwMxF6sh
/jyH02Xbw83OmVjYC+6RoFx70muTLOlT3PEwp9COeleP03bOZMfbSVTq3kMT9E1OkZrUrBZhnfui
cfiLFktDT0DqbabKKMkOJWAA8Thc5oEDxJpaAbSv1dS2iDOHADx0bulqJjJs8BBAMjLiDBnVWZsI
Si010cV3IxIJL+f+tzN19U460JYCxjRfWybXnJkW+kKaPp2NAvPsNs83oUVsLJYkFu8XJgq1MMkV
3nFRl8YWw/jF2fyF3EObPmy6xDfmraLKchSrJ7Dt1c+6S5KDmHh3vDacIsdWz5unhQ5cu5xW8nFl
NxX/xIVoTbz7HnOkdKYx8DWyUEymI6WlaEwTc6YBk8A39wRbxmvuvs0hJTio41Hb508h5bddYc6K
NsDoKthUjL1PHvDmcFrM9IDYCO6nbmyMHFReXvGTRiM44c1us2pY3S7w8ptkR55Jdy36dK+9zNUt
uD6u1lQj9HFgr4Wzvqux+n1zRcGJNQMWTE7S3Vs575UyOrA28zFPUWD8DwnD/sUFIC8GrFVkvxGC
ZNKPVOu8DuH3cQrG64Cwpt07OfPULn3uKfoAoHe+9KSoJrfrOlF07cb2bPgynC/Oz8D6JlRPA0AG
pc9aZmRLLZEAEoBpEzwFzDY7cyg4Q36EUcofcn5mmKKcqnp+4SiKpN+7mAGPrVK74SxPrPpR5GjR
N/OjVhmGdSvg3Xey3EHekLH1+BhWeZBCX2rGy3CSXLHqUATN+TG6tRPpqGNBze+wx2mP/o4Z4V5Z
8Ni+u7lmgSHHw4E0O1/N+fAEmW3lUaMgD3oiIBpbFTAcWcHKtgSs+VfD/LwuJnMuaqMPs2yUAo30
e1FKW2c0GaRiEQHu6/b54rimUFUcfLd0IcKf5k5pUEvZoqIbRI9td/HenBtp7X9FPerH12XbqFbB
/VxxLw39deR3eSPXdYNVUe0AFqQuEgtQ4afzWJFZkPGy36cqxLsq5O/fLF+ILHeUv5Pzq+b+skOX
Dfvl2Zawc3EC5zHDxeROnajqXYfyF6J7NMSl+YBIumFq/VZfhBKL3lwNWaiXFZdoOxd8HhKMzl2V
gedArq1HwD/rHi1cQMsNKoihIy6AtukIsPAuiKSOwKVQW7fqxApvG2MznLhAvOIP9xVpYESOuYfJ
7IRAD+rpxXduPYN2MTo6qAxWiS5JdN9PlovjjvcAst79vPwW/h9FZWnAKy4kA7z+IZXsxObQ1qAz
jdQ9y1Q2VjmoK9XXAyjGB0//Vs5s0lhn732gXOf4HDij5Q4HwvCKZhtfNUwvXMCx0EalLVxLL+bu
A2ToP+0LTCOX1+DMjkibhQPTxP5fJ8Z0oeEjX8nAfvAFE5ZpXzjQontVmWlhc1Q7hQEOjTmt/WXN
3rf4FSe0UjT9Krr0bCWM7a4eDnp5i3egxkqNJd/jGKDvboO4Jq+PkS9MKiPx7xeFZCJ+zhuuDnO/
+u/V+hzWpxNm0/+XoGY00sB5av/pMUVehyNDTN86z76sjLYrN2+Di1pG+e2fvPkPeupBxqWVJdDu
8mQn7oBeYWtuERTNBqMEoEa13jTrhTkoFuuTdoaq8oUO8jjNoUsUsHUutW+Xgj5sArMR3a1muKFl
JuDADPu19SHAdnMSgto0U0/OBb4Pf8aytJeaRNUGncPzonqYu9edZUyj5yB3rQe0CPC0na2E825q
4ED/Q3H7RCe1iy3XKkKRHCIawwj00gDtNDFDEr3/l+O5ThuUmf81nwV4CzEvUijy7UGlHTLbOWAw
1E57/X8kYrMIH2oUKgE2myB9XU9farib1Ktoc/PRKPIJmK8uj43LKyW++i4J04MGGXKMOGJtGwdI
9ck5PMBquGPAvHzoRGUN27w5o4YwrSBqyYceVfaRJMxOduBHV631moFvwxmwlfX2oou+uG8onDfu
l4sb+Vr49uzhPyjLFtC85hKVD0yB8kuEeTLCQ31va1V5EJVwUlPm0wUxnAk6ZZpmCDaczi1rrXJ6
8R2n3a8msYkHPHwcIJUW4gJUBYRZUZYzc4QkTCLN/cVsqPLXoeZSbAyvZ/Fr5fVEiNiaDG7yMYX5
xGlmIXCjkciODe8UhnJtIaRHiDhnUvusE/MAOZoyt6c/wwfiMVGAG63LhBDawlPOpyQeyzlePugn
2CWHGFjNEI702Aww/4N61Nmvi1XB+G1yF8qNRVB4DQFMWeX6AxC1cZgO8S21k92vOnxcNHqW/2P3
EpaGoAAq4o64XI4qhiDqqwVKeOWv/AGA+ByAraa1H6LajxjsANw3NkUyjkGFJm/WzkBqmvZntcXk
gdmmB4NlUTxeUG2HgIpZbfg8V6VNKpEu96Mylh75KlzfLwt95QuVaEnmL2uOQMD69wVOwOrqp484
L1fRE769TBOOV87s+b04dRtXkKbvnWjo/Z+8G3Pbavxknxpo6kcCzN8uhakanI7hjynuR/TGDme6
2m2D/VjaSmzTJlaI4qD8kSiZInMW4KvnO9H11IXze7jxjyokjANB0sS43OI4bVT93WWTPsPIWpfF
x20Kn3Ggl1hHADPfQaiDPd3CDkzTxH5v5vqG66An4CFbIMTVs7IT0Wvwt9yjStkvOkaKfQL1dket
XCNbiQdUwmDXO1Bmck3LGp5s8ZTZtPJCxgBocGmx87WVlRyz8U6R9pcbiVex+NCoDcIaI58VN8pa
Uqpf2Z97ZmygTf7YlQf+I+SKhdMr3SXu5NHrn+lsSzCaDnwfw8HvlmqeVjmK2ZtcT2fdbk0lw0xQ
T+owTiHSdofwRp3NAiXXt+U4XbM1PV09KdLAb+BCxEa0CF8S6AHL9A2RGhLflJEgQYTY+k+W0jKV
E4RfsLM33yzU0MKfLCgLDxFerWzRVLoPPG1kIDG8CrdWBxPeo1lxGgown7fpc3Ej7xVa7DnP+t5e
uOH0CNKfLHRKrRtLphJBOMR2tASFBA4zYr/Ie8pT87OQvHkArSpN0x1GothTH2SftdoSZRT2bUSJ
4LA/Wfi8FoEaGz8WNDV351Uoezm9qZcHmZKe/Y2F2Kw/bZf7IuFboAihsvRfhp5pWHO2wgNQmAQJ
HvT7E0I/EBlcM4+/WMu22LXmu65ZwSAtzOThDnse3PDi8gEAQwTT9y3RHoyXr4sY048xcMEi2Jqb
B40YnyqNbNSwA7KI6XwRArkij73SikR97DbazBdOQ5Jsikwu0tEWYVpoQ6/MwYXrrBtun8aOsyXT
X3dqU7M7ESI/sbQzp7Zc7MDPoVd5Kn9ctv7hELVNLwCOvSHvUMhavx1/J5kfU6BhVZOcrC7v6Kcy
C4GJlcjvH5E8MsqrjDvAOsJf2LL0wHfJpgUfXW4icfQ0nKRqslSBoCDiFWtImUswUkBQqtqP8iiP
fCqmjSwxnyOn3L1E4HlQEMfHUJchq3TpRwT4vrAUV+1Qtw5a9sQ1KOwnG5r0QYWTxqKZ4OhSoxBA
KF+cLnPE0RB9442KZaySgRAOBCSGJlXATDVXRhjT0i0z9FbyWOiIMCqoXl7kwzK5SfbD1LhUACic
AZXM+QZN0R0wyK1q08jzmC+CSkjxHlr9QjSX31tlkvS7g5JCYkoGJmBR2dnB/E+OfuobCN2VIej5
PlURAQHF1BwAcd39l6teDpfqe+KuD+XdXZRst1uI+e9dl2So5mtUPrw+yA96how77ZbbLxYeBhKE
iiBK3Uja1xJWPXc20Pm1WV21DJRSpfk+SaItMNrIZjFRFzcQr9Nj6CFV285ECUZgJpXkMb58XwsR
R62zhh8NAHeSacVabtLOrtIM9A9Xun0xZQZC38dJv5SbU0BAzQoZBuDTsj9EL9JsQwosrLRxSoQ9
yU3Ofv0BKkiGIMNcHF+sLn4TUBuZz6T8Vyz+p8UlOhTCiH7ah14tw2w9cbMLQKw4MxoJ2m4X4M7d
0pHit7QR3Tubby5oD9tcF0PFQDi3Y4yJRg99R+Ed5mrgtVmjC/tOrf+xxhnsFwbkh4AU+8lQNlbl
BWHDOpCFtZGMm415ayRnRSIyDVBc+4OVpUUJHjXFvlEZ0T4tS9JRlD9OBpJQz0DWDO/mrIZMt9KZ
zbDJEwzChzdxt7p43+kUBkNqx/KAKdQUVOu4YM1fj9986NfBZU/f8YV/IAHZ68JoXaSG/EVmA91Z
Z5gqKFn5fJI1xV6uSqSfLelSOatiPK9TO7opJcRkBtBXtVg531JCyo9KaF2C3q1lPJWWvkNAhGmW
gcHIdZHEc2KLFE6KvvMiiLKFYmbjv0kX81wICDXXHs4lW9/MD5ChESHSrmK4D9KzIaDQMwbSwvzo
YFzcD12ZEJisZ0D1vw+3+hENUyqWm2tdFVDdqB7fmwb5hUNph0+Tn7YjArAGfEcN8kjJHuxz1/4r
9dKcZsgAVHk7LoEhxuJH+Mc49ScI+naE8/DlItEXxmreeoi07931DN+r7GCskdlJLuNxpBmecrel
mGQl1g9jivez/9UgxEz6Nx+Y1WV1oLFGFKSQpVN4sxCsCOAXMwYl/XHNPHFK/y/b88NkUcySN3b5
XURETgbw0kESYG1hrvk49iZU4tC0kyb69zKwt6D0fN4103/d6TPqjP9i6Xu8uK7+B10CNDSP9mAz
9ErH88WQGjKVEmc7f0gc85stnJU77c5BD30kO5W6mSuJ/dVO5JMZDC1kjjS0ebViBYHVYmHmHalJ
l+G9py2IRFAi0huNOY7SWkMpah/KZI5K2S9bl7CkBIg5VUIBzIy0xYkR0vZTzth9/Yjih5YzyMAp
csZasKaqhUoNYlGlA6myQbPui3NJHKfmUBFXN358bM0U0Uwsyr+Vj7qq1keaEWVxGQ3Qbu2UkKSR
agmJV6FygOWooVi+E4t7/tZI7PlQhJamKl5Jv/R13l5280/z5/tObs80wi6TP7Wq2jkDMLzuxqqm
7y3C+qL/LlaCM6DnkEqdf5v02UCv7KGjNIbCwvPf2P81/Mpjp8PwWZJo8bn/bN+JiGpp1cVY+bY6
KKubNw3jCxpjBbWGJavnPTf/YxQYB7IpNOmsw+8AA21BeEhOazMBjldvBGKuyKiZVdvQpwg33li2
HhoEN76AfYjXHBqJmDIjB/BJ6e94pPWRyBbnhNBL4I+q6qsyBeutH5FAlCSOO2S6IxwIhcAa3nfI
FtZmXo16qETPkBuLIzW9THtinjigmefYJmNi6qRZCOoK1ni6ReftgXNf7UTTa6t0+Y3CZ4IhYPtK
tFC1BEMNfLFIPM2Giuu5+MUDb1h3AnlnoIslSc/qhof/qBC9z813WnDFWp2Yhp1vW7GLE5Ddm//r
010U/QM4VL+V//8LUQH6diBWYqHYcaBGGjwtS5naA8oF/OlSjVyA8xR9YitGpz2JaESYUw3L/FkG
Egwh5lNZ+eFD7i5OW1PwZram5Br2n9J8AUN3xauVvcH7oD+VHCXqAbtQ6ho+o4onwx8V4r6AEBoz
5eLiPUJk25e9X6lpmdXejONvfsNFQJqOtIMCiyGMUrsvI57gNz0TnKRKnsOLIAbnwcN4Cm030E00
GckALyOtqlhEVphrPHDQQ4YNvtZMN1SdYNri+RFx1gY41eGDVHt1+d9cULiVpgAisskYzISMgD7g
XekxaOwiF8rlUkinRHE5PZc+WVsg7efcbiaUbh6vqHZWh4xIUpOGiPuc2pbhBzgemQGQz+nJaGsQ
5o/skiRcQdGfH7HLW1cnSMFAC2AveUI9LGYixg5M7OeaAXuLysnoYVa4gxjfNSJc6j8FSYGipvTm
JnvRrJhVYyC+iCr9aHK0a06A27DD6+1s6UZKNSc9ouo93WzenkV3OMHue9l/L2pkpvgYMULsYE13
kPBQbOE+OYhTSojaUh6AgdEmY5QPZTTDFowF8Zbmwu2DF+0lytn9ZsvTQ2Yl0GGPv9lcba3ZMjxU
xO7ma/xeV0k+/FaB3FOyUX/WWjz2rqccuhpVphroEZVHBb9ePhQKXLwdB23kvv9W8i8pmqW3bgag
pCr6qTfCFkrL85khMReumLf1TJwaJJRXsxrF+x5NDwtYCrNDQYVcPVXn+GMLojpnKnWJtTOB/O8J
HYn20Ko/mBSrOREG4cI14OAqVyXbMKWiYCFSLTFUozBj47Yq3mO7j+D75lo4ZKmdqWwM0MuBPcuL
ujlsNkHqDJwyNjPCQRLKNuzMdywkLovxvIKhLFNis6w38+53RdBJMkpaZWq9ouxac5EZ0RvDM8Ty
iTFGnJWn5z8DajEaCjGICV5XvfdY2oPjZxY55cLFZgCu+LAjzNHt1Nw+8C3ddA7P4PwvfbSoaveV
OTtpBHYNzRB7j4g+LERKCCZUW+qaiC9fWOfymvTww0CbTvM/n8TFySc+Zj/XdPVC9VAZpARbiO2C
MmFtGqP/5J5jWmlmKo5VER7AtUXNQaebYjwYHBMlbaVUx6z+n5qGFu0XSLkfOdcTN58TpQt1Ev5l
KWZeg58p/vg8Xx8mp/xdQmoGdE2u8LkV61LdbUo17uBsirVGtmX92VvADNXMw0qqCC3olhblsqVD
ItYjd9k4AgxqE/dUTzvrGLNKUXEURYjVqJtXKdP6elBRecrU4hikqCTddPMOfMr84OmZfFj+1RAM
07njWU1u4y+IZuWwLQzc0xkKgAuVkoAYEU3OgzhACC+PkkiBhEeFplZR8o4u6UHm4wk5KWYHTf0+
kl78OHS5D4gGQAzQbSkIGGb0lQqvpZYVGa/8t3uKpJ/vzLRdexiGkqZW8KipAUFEHiK6NMtAkSBO
JTU8TbMFeDlznp1XdnL4xwmCLAU5TVOLyRgqslICFhwrsP722nog23nkCR9FN+IvRirUQ35sUwul
TxqYfG0Wxo+G+hbM0yVALAXKRcqtaSpQZcXdvudfb/4idMTChMhgmYQQTD79Gn0JFiO0ne6Xih6n
fRBIHwQAC4KE9F3Hd/voYpITEHGXuiC/JDKMjnNiJDu2QezbMeZJz0/DdqP0OmeibIQ4zPIX/HhP
0m84jrckADtUb3xMuHuNnV/xKBqPCzoqlt0SFUu7iYA/mie8S4e7YuUPhQA8zRPZ8nYspIyPZtzU
PcaKJChkTmJ5C09M3f3V5CSDnzIfQHyhMEQMyxaOPJpXfqs626URIR3SabJdWIFqpxb+IgDs3sr1
J+99b7RwVFsNXCqq+TYcerqOsRJR2tDF+mnChOZbyJ4xEoMkhlY1sEJw5jJdGn+oVBizb7q84Gnc
zfjR83amFVagdcpc3bywQnMQ25r5KmYLcX4tcCtaNRU05RkFZQC7r2tobwfR86DBQF2e7bgCsN5k
/N2YU2xEWhH9lXq6c32e4p+DonxZaUf8uCbWCpGEqfnNcho+eJY3dl06cOGMxnGualYHp5MsFMzP
dprzW1MDzvTLUtOM58qyKo0wm8qRXP8j9dI2cRzCI3sR8U6SYrIxVShkFqMEOhOuWwhDPaRaW2m1
BFTlyf+3uJf2wt9tAWGzN1x+8YxTXiT5GUxPPp6nfAnNh4SRDOTy9VqVTo6K/2h/bTGdkgZd+gMf
lQfxqnixliZNX5FQdQECnKHZvoYMlojoGf/wmkJCx8/5ZALdX9eX2LzGlzlvbsInSQPMVjhhbYag
AUwjKyF8hVQzMzmAFRFzD5gKs5he60gn2qxPfXi9ekl/PeAn0XY9t1xUxMc5ZBmoP2gmedxhVbVB
8I+ehntRQwfhaiUeXcnj9nwqS7hErxA4IByDYuy8bPAIDoD2I+tW0BMSgr+O25tXdlZZ4BH5EFZY
ODYc/Hk487Ya+q61/5aheyykoVdi5x0Om/AnCJmu271XkSaXb9ZeVKOPIEB5birWx2L6CNIYZ8vw
0LRMv7i6AjJz61qdsuc3530+M5hIIvWe3KzvzeKfYhI4GwmOx+ZKCwu+9rbyTq+ulPjKGrs2WAHw
iui5xi1z3EFBrMKTQ4QuLRLy9GBEL3aEZhE4Gu3bX8dHPmB5AJ6z4yTupe7eNn8VuywqvJkfbu0C
osCtFaf7vKJhLI76uYw+jVIEiXjnivD9DSYZkv+MHq/GW86hdowesvNuVf91EhjlLSAocfzyFL31
N4/vlZWLHCf3j97X8MU0KsYrkbptrCsTHP2G4IHsEuZUV7LO4Q3Tus4ozODukHJOsEpTMqN3qHX7
de8gsbrwEPqGZ6T+BO6LFZA3K1pJeNrqvYPb09Zzv/dWnusYMjUeP2q57xqhnD4dv1S8AeZgfp9Y
vnnc/voRBDRpiVhxZ/O7PGdViB6dfl3Hux0QgDuJN9rLjsyDGvJ4XysdewAc9ZkacYLAM+8Zuwb0
mBexRheR4ErPN3yJxWDtf1/uCNNS2PNUSabdi9YTiBFyRte+m6TrNsrw1upbu4VRxIX8xbSy6SD6
oSdxOMBvcWDyMw4CS7wlipP4Dg0NJHjhVfx5dZacWpQwQnZ2cj+uZROg1M69Qdc+2AtNBG8j1Jtc
Jzgf74ocg+eou3tytlpyH/eQkhPC7wJcN8A7LShOfEACzuGOgrcCJQXvKPjwRsYJ9IIYW8whW+4r
T+ttGfP5uSlMceFLOjbrJxtuz8RV6Bk1fotlcLL6YgktQst0x5Ex/R6glsaM5m/jvS+10YehHQCc
YMzB5kEowrey9IN1Y4gG0qntSqxGAnJicz0UQDzYG6syTc0FRxTD20FkNm500NqFJ2qvXT2Y4uo1
gD4zdNR8Vggpa6Two9LwHWdAw6uFl3sfarE6pBABSREIGFnOnN6/OZvS/b86NVqLi4rcqo6HM9r7
wRV4i7MF+LJobLmHUGKIIi2oMlcfLfZqoU028GITFpjwqlePFPgpCPD3RAM3mj/vLlddnDseoiGu
6FEVdrc5CCQ9aDEkgxhfIx/kUtKJEt/6nGG3/mGQXxfLEPdH3093WsXHoJf47he7Hl8U7uvnWQmS
qxm6thJUfNJpNPdhf4aBsoO2isvIOivexx7pOtEoA7reoSg5Av36Aq7yNAUkazbwiVsRs/dMZv48
I+NvZRAR0pMCdbFJRaFBmyv9A3BW3plaRUOgK6P4JYxASoa5axXXVmiOFhkBTCJVTQNlDHPSxxvX
pRlf8wb/cOmwWMLEu8Awq2QchmaYaq6gseXlxI5+/T1jBmFZVNR3JubXNnNBFA6AM0w7NvZcc+d9
CTEq11e8xUYtlOdyrxdII34Y15yQxchftApzymJtC3moNhmPUkMtSlXbzGl9DCh99QCb0uSwkJzr
NG9zMHawKtnrbgwZNjHxyfqN174SI+sRTYLbLAt4nC+G/1r6KZDm2xNrAH0dZp6zryXH2tcWpHkY
4itwKOnpmFnj4KIxhU6jvQUOLd4uncjFziam2OH5NNP5WMQXeAIujrE4A5uuSJ7td+OE+Cn0M7tJ
5R2jMIVsPoxLhtSGULH3YhWFHP+j9Cjvb8zQmt4M8wIWLJe/dTAGs9W1TjxtW3TClFX3R0mjvNeG
ns99d88IPjG9oorDga80P6F/wnK3mYjOTktrTVaDX3rZWsjteH4+/XHuQjRzzpIY0Ad6zX10HD96
8Cn8aS1syIH7FXRDY0pVeGuez+sBTKtdYFObzVYPWGNJQqqVf56USm+jq9hGDVwcLfQdJhbPPWjR
dPBblieXe52em2s1i/8jkpGjqZaw39c0XTCX640ibSYGCdSAKMm6OteV0+IWWfAXYowsMD8fZCPS
GfcmTAeahpL97txenVkrYFjIFRJa3jsVSc5RTn6LEU7FX+qE8XvkU8Th8LqWVtLjrqwb6KlWhpSe
kFV6thLn3zsc9EuemFRD5mO2fnVNAnEQFgQfzcAYpugJMQCBFSp8OKlSBneWmWOutjyoiJm1j0P3
pAZKYlw9e9IdUbIxDJR753ixLeVJbq7rgP4OnJ/z0YggXjEMrF6Xxgl5RSiaPoYyJ32elZTrmvQ1
McL4sTBtBJW2FbKzItleKjgaR9WSQslxJn774CmvPMKljF7TE21u7Ff102u0d6ur2Nymf/UWzphZ
UmB1mdP07bNB2GWtJUSNBSU5GQVb1V3Ewz11vissm/apWExuTJrVdN6LJeOdOBmjvIX61gKJeDaE
yvRJjtob5+ctpQ7HcPTzP8qwsGtGYxDcIhbrmx6mUE5RmJjZDyJlDqjsPCVnEd7z6kc/XrGDq0GG
4YAcc11K/sbKsocZL5xgJvuL0i6bf/fMY+z4qBuBCsDKy3rN39q6HMuMJMxX8AcgkhD6yVL9UTAn
VKqZrI8zqye/FyR/3Oe5icNVHTZ/BtJhAL5IPlJ1bKBFpEroZmLeL4D+/PEv4+ucH1Kf6pdoTHtP
hBMghv2ZWNuP7pQcNFS0al9BCAm3ohZxG1BkRiJaXHfNggZKjnQH1JW50SjdFxAWpBp5MfldZK12
OFheVJJCgVpfbI09shRAs/FJZ4C2/I83+oJGzZ9d9Kj9KD4oLd2Nw3kvLYv2IZvK2TKz/+oZjrte
0yVVRqwcL5lGxCPY1qSBQalQnxw5zV5U2HPXXEnHHb81pDk/VsCzq/cgewllUHvCvmFY0LgmWUbr
Ol4gpUQYoTY+deEGG2CptRlQuJBhwx8pVpu5J4KSjfP45TkASX6aYlwez1l/zp1b/CZ2Dti0Tko2
lNxtHMGirZpzNeXq+dq3ctRVsV8tWazCL5mclh0z7UxbvUc/yrAJcqvIsT684heAKx29ldHLBobA
kKjCC4Ki5LIGBRpnZDh9oYVjaIKrbrdZaMWpKNvgrLpSP23QMcxKOkTXtbUMKYWFV0hq4Bc+xLE+
514ZUE/sZbk7QosQApjQzhNQ6sy/NpawgQ2e8/OEk6QSR9bUIWVlMX2heZ88zUcoen2aDgWcWflN
M0tKndRv+nO0rdzFO8PQdlmBClNjVVZ7k2Q3VgnnQs+S1jDHNfWHlh4wvdrlv2zKY/q4cK9xPt9A
ORfZNFYsecAir01gDeigiFTPX4e5ktntyzWzxJ3jDE19AwO+9N3YOFexWfnIfF2eEqvQIgf+72wd
GvGszlQRnYDIo7iIE7FYjZLbD2H9bFl3gic4lH0naHQtddq5zavg1YjMMPUMOKMpkdMolOX6gD17
COSD4CeG1Iyw8EolLaj2Lqnb7WfEOPmLFlp6U2NBMUj5Ucri2KnKgXTk41zyDqVt8V4VBWJPfYfr
5MkSs5dwIqDpOIeiRyy5/ABl0qtCpjqJAJ7/kZ3sq4VEP6twFLRrxncFSJwzhYXDMTcINSSVCiMU
9SPoqjLtWB2ZqtqYzUnSl88cZswIboVpfmlzEjc9ol8vfIaJMS9jnQo1AlFdnQPeAZ5RYWCSZCgk
IZtaDOAu53M2w4EVe8fXQP1Mqw7szZut+vl/mIxc9dJWMNfgjjng+dU6lwhhecm0pVHwP1DS1+rU
0YGGlBOdaprmCmu52aSwsh0gUeLTkm5/8pE7VyOPnQ4r5glilnoXxXFUIuIBh/MNHjhb0L8jvqVE
7RAhs5Oj0Yq7MalVr1Zyx15PBt1czinS90rDA8kjmshjA+hrYpLL10LbgBq/9c6usCke+DnLtZUh
7aSDFL7fuUI5lq51DjC8AYcutmGZWJEvfQO4J4Xdgquve9HT7OHievNwODtpzjaz6Os0Wla1Jicn
qxtAZ6Nx93FjedXIkT4v56VLZzRTDQy3x4Bhf1BuzLCTNIo1jlzNcC4G8fCvMbM6BrbXGJZtjx3o
quS2jjzpqOw6CArmCaazcruCG2VR5p5vzRPjbOgo1ObRjQ4fsj06aA7AFsLXZTuv8AeUUdLZthNQ
06y1JAEOigkWt5AtYT1S9H7C74xMIX7n/brbGwOVfYPZ7pZWZ43oH9WZVhQHY1XnU7gDDdEEmfhH
fesb4wOdJqGlVIaqHOkuH/g5sR8J4eYQA6C3dN5pkJ++iMJ9GQWTc4SpuvVfoDr1gDXLdZWVa0qI
ViNgnaNsvSZ4uqrYEds51qOTiEP2rgri5GZ0YGvhCFrQvX5+/zt8W+ap0Ii4812p/ogAllj+6uoQ
bnVuSgg87rON2BuCPCcGCe1kVycfoVlbP16bhEwQPQYvYngpsuWzI5HTOcXIdjdp2DJMpGdItc8Q
MyRggGbsXdbeXDlhuP/6nM3HXJgkWMCRebErdXf2GNuKZw0gifQtkzrDSDnMg6NElalPPZZym1AB
7FoCVFgMSTndn0FRJPQAVOF37Wik5Wz6HUVErX0G6vGhR0GIJdq2GKplg+zac0EZermfTE4epp4T
pXSoAwJltOxLQ+Y/iIZuadt3b0GqhajO7wPAbaWub0/4Iv5+RlACzDLgssfX5bkJdBng6TQ5lQ8v
Ks87DsYQ0IpNuB9Mu3T95Fa5XZ55lOIf/IsTYCnEdKnimaUoVYFh4Is+bKR1Q9nWDBa+mEsPeq/P
xyErLSaaTxjdejjcof74JO7gxk/OLijdeCLMsf/oNJNPp4fHaNsktBylrhAj0NR5XHh7kRkn9Bkc
eL1y7CAsEPVviVZvuNiF2DPDkqPEIkYcB2nx3XVV8uHhsXVRJxUmVcIiBBED/QItHC7is26UEEor
EZeVEjtvcnO8q7Cj/b5upR2Qc04tjjJhDo9s+A16pKmYWNky+1hAt0g2H/wx7t8dPPGLohtqaOgn
71e8Hffkz1WRuOkB354JgrB+plCIq8trFy/IDYjjjfw6YW3QiTrWnqhbBifo2jS7NUy7xI3Msq00
j7eCxWgB2KfJkvwnEQunD//SCz7+Fv8zcaspiI4L4SGJCPIuBO/8xhbzdTrrWPXgbIfzTi9jej5o
2QQBfJ5LrxthsKemxndpbf6DxMnYYHy1Y+mgP/eYg5w0avCLoAmIr/kVov0hfRKoxm69y79mjLYG
d2KjGA3jzIzllWiIc8rj0p1i9friWgr8Thi5wNnmXCCyYCozHWg4Ku22RCID49/dEYbPmoPi5frS
qV5UuPUeRRKhjYjX+BLMIazrw/Vr10ECyAS/dxgVytObfw/jCHp5GIqFJg1YtCP6753Qdg/2DpSV
CnKhGXQ3y15WyiBeH4X/OMOxQklv8WpcJEYT+XZkpuE+px7RAplZ2lkS0stwONwuUAqx3VI4ZMru
UKx/rkdhjLvd9E6NXJuiyTNczQtW1n34DvMNV9S3NQOA+P+Ht0YezOyWw5fy0gi4tzkg1tM9E3Fa
Vd2NUc2jVABXuyWYLfR5mT8c7oim9kdG/RjghCtB7LWrTCH7dOlEh5onbOHZUVFhFjSwxLWD8oTE
/3yENmzDnSJ9Zn9E41GJUZ0uUpryuxgfi798h2eFxDdQAiIL4w7pptukzFn7QyMyYLtisOD9c5Nt
INE3f7LuQYgavbKid8sDA0p+FEUsFfAa/Y8o0bQqi8QhydJjOBASVdU5hRiYgE0M70L2ObDCwqdx
sDbRfx9eKbKk961hB5zFcDT/JlnkLT0equRrVl4Dd70x7EtIJc8DquWafiwgm7K32a3XSNLP6GN4
CD41ZWjVQBQcTP5DoBQOa8zb4nvXGNrD+DECBoLnUHzK2Agf/itywz53xG8glh4HBp2Xoj7+Zgb2
aYK5UHcDLGVu05OoidtsfK3LI9Z3JNp2quwOQa5OE02yHXvHhsE6y9Qyjx7YRQleV5l+PhcKqupX
CrT1VNNhqg9mzzlkyQcpIbChNV1Av3Fm18Pl37YUFF7rbMxv/skG9qdD0C381NOKRm9BwwUS0u/z
l4HuzMq0CxEZavx6UbgDcrH6oTBMSITAxcwMDglxQDMRszbyawAgT9cwSToYKd7uHESY0hYdlvTC
CUpFA9QrSTXeS7uUnYIFTKWUu2L/0tdvIVR9EU3LCVI7LabdePSTKTh+uj9pYCus6gd8VIU68Qd0
s/iFst9XdAtSLDQclXlYZRfRG2XSZ6y7eb7QWav6rVssBSWpMF7lZnmvsY5+2yMmOonf7ANKYS3V
UmrL9NAkWc7uLPr+4TuhLEp6yr21JQH/Dd1S3G8XjUxyXiFPgCOdNls/JQdrmkhicQfeLxrwhHph
F/eeLvMuNDYJ9nz/WRKVa25hCfPm+PP/TGH+VshVSvRoY/Rj9YQSpkxOQzLfhW27q5Maq+zYhhhE
feFoEDSbOaI8Lc+xT+/96l7oVzhRfijil+7+MSB5cuQc/0bLEO+LjLyET6JByeyn6VHEvDE/4+Om
/ofJuLQR5yZBHbHIUeEQkkfYbcO58IA9hX5aYJr4jOxJGWzKxfeIa6TAps5g/bZh74cXjNzd8JPM
G1I03hkEfGl/ybHXwmKaxgQ7Xzgy1QPHL1WxMhZlV/RE4DZjtDHbO8uj7CTDuCP2TgRYyLXMDCK2
63F1M3LSYargYyHpyxU6bVPSR2O+RXBlAXZEjNOBFR4mVUblp2GeSo6gc/zw2gW07SGrm3MqKHkP
E2R0ixrFKX8+gedvIPyW8KMBJAW4QnkC7kVbXg5oK1ea9vemipN2Z83MTNKbDtNgoR49kzVl5qme
Y6uSr+Nkeek8thhCYdcvva0Kqlktb8OnV6Xbt4csE4hAn2WsBJIEkX+GFTiwq8hwlfIhNUh7K9fK
7NPK6c8oCOPfU+cSAtEdNm/S791wB2U5RQic0hooX7CDpfdx3U3pUbuKZw5VyLOqpIrjpG9Pu97i
skuEMYssVh1i9hTWUx3p3Y72hlni5FxHMo3qlQYzT4G5kxHL8fdjBWKG/crMoO9ZDvKHjt4otrVy
DM5+m7PPsrHlwxtuHbmzRs+KCLmPpCkL4iPr0plhwXx9BwvNv+pZrTa3qNZ4MyDEsg9kzRl2M6Mj
NEwbap7A/R9oIze732B+NPTCbw05xhEZio0Ne3Lls8DKMU5y7ajGHepMtYqkILAcS/0HOiSYQXHT
CUSXaZc2zNFlm5hIRvVPs1MJdBH2v9XsZilJpsM7UU1UVtDRUguIhvYdcYy6RYEpMO3UQqdGv6FH
MPfVTlaKWOdeOuP0RI4GKahegrzadr3cb6eIBExqzUHgNZQ2bD+R24qZekdV9WyyO9Mrl6B3O9WE
JJmuqmiIj1VJ80xLjc94m5IdRFEvJ1LtP0v3wX+7huC69drXTdWLPJSHMXj8IKzScvto/z7cS/u0
eYSpE6I7ImudZruq8TkMEqQORpUv2cB9tgiZSWTjCwcA48V7XNVVikrRSBecLe+UtRxeTRxknOSV
kYc9wCgmfGhk0GO1p9yWCLoPxfG1mfz9IfV3Co4ZTvfMih7wdOmqKZQF90tFvceVi/ExVjPW4ndL
cv7PsNkffrSSjpces9Um/kiwpsP+VwzSMjFvZr7L73pW4/41plTJ1H0vihF27b8xQdG2p+n8ff0N
bkHOEULJbZHXLus0JcYzH8cfJXHMzrUjE8bTSaZ6EDLAHCwLSn5s9V/a6/86KMH9AdZpVNWzBdhU
LY+J+Tbi7kmAQGETC9o0OSMWaIAD4/wmELopb7ZdQHtN4i30M29VBOwnriypw4i8lZ7KVuDzQrCj
HWkA5KiYGYo81mYHq4yOZH3ove8+BzP5kY/348AlJzm93YKC9VArZBjph+2CQii03DufImJiqpIq
wxIc8sNoc5NfT3k7vRwK2xEdrr+kX6WT8Fveqvz1Z2ejvuwaSWl/liUIOwhx/mCvTrUosLJOVjcp
mo0tn6Wgzd/bZPzrQhnPMZztzi5fJOk8IWiUEN2ZhUpZFz1HRFDxfHETeqMXIAxCxsh34d404joQ
iFK45aXoBEXPfYt/P7felfXM4rDpa0MSYlYGSGrhz5iNLuq8CJRWCO7ZBhuassKFWeRzij3sLJ/Y
pw67xGOEF15vb16jBaMa2TBNxM7gERXbXNgHWTbe9KIJnf9+xWG8uO2EocJL/5ThnYwHecGZ6Trq
xb3riFJZ6ZPzGJB4uu5/i1iAaZE58zxz2keKe5NLIg6XYfm/DsQD54+z+nG6zgspCqYpl0nNCeBh
9wDhs4ofBePwpVI7A2+eGZbuapvoo0rMtskqJeIkEoreXTbmVm0FJbEeXCueDR/1IOErkxVVjPVe
MjG2JU3jRN5scQ87J+qSx1jG9z3qsYZseznp/L4Y2Dkm9QNKVkoMN0Is/y7vT0AqeWqJ8b1lHz5s
s1/HZf+RMC0WJ/fn9mS3Qm7Lba11Gze9cVWOrFvEpHtF60Z1bvdY/apSkqs4acu17bjEilmt8HN6
+prQC4DjvtgWEWQ5I8FTTjrGjYVCcIPpkRYtYu3Ik2uv293RgbUNB8PzoqFesMHLwnS30vVUlL2o
R+HyEmeSNzH3xKotpYmBKvDMGSmQqiar5TEfOEiIHCcquD4wJSgwbgTYGh+ejWK8yG1CT1kRqisY
Bepusb1Gi2uqBAtDqMrA58ANCzbFOKvT7jlU5WxXUyWqqhHigpi6d0hD8VfY+U7sveevafgcyLTJ
yUd+cAHMOI0Mv2D/P20iHt3C1oxAyOlbQWpHRhMVJcB88avyvFghddCr/z0psyEdCHK7/wKr/Nkx
VK/K/vcMR/K8kRQcbwFCrUsixIjU2BwmfujR2BVRRCsC9vjXTcYsmt1MQrBYQYV5vasjJiwNpFpH
Zcjnu0COyVIQfeUQ8mMqSvwp3h8lvnqEDcs4sfGgdcPSZqJ+BJOoSr00pIRXhRiSYqVzqZ6YcZ3M
hQ2lGNL3zBpo8xCdguYVykPAda7SvlL8SAFES66bdcdtZJ6ZypPZw0F64C349yTGgjggm9M/2WNQ
I5yZWFIXDdjvu00MjdKrcJ2b6FsGGi7m0tA8/mLRpHq6h75OBYwJ0iACXCAo6vslszSrgKLoN87F
eU6Cvx+6dfYYVKAvtn5FUOovuDUzAZg7cKfl8kMyV0q0UNECtWZTvPhdDsmycVfhSKeLwLEN5slf
/G9DCBciH8gREFc38rpEOpALmJtlBf4f/EEjW+PWugPy9/39Rj7DKHedsNUQHT/y2AoO7hozIjE8
9k4/IRJmNwDFgqai6eJ38cUQoM1MbvsZzgCVO6eBcQeNqllTH9MhoN5Y7yivHYmitCWkgTU4fIw/
joH6CAQub1tU0/0IO1dgCY/vGmJC8OmjtWlN94vbv0JPsn42pYeQAyWBwR6bqQRtAEg+2IiDjJg4
w8bTTkWv+Np4GZtcqrtv1aRD3tePNJtVcqfKvoZg68WHcUx0VGL2y2Ky2kdBUhPHdtdYBziyDWhi
gAbuAgTnsVlFQqASHNVjeFT7S6KNnKrKZgaAoxDBFzlg+cBTWUYBF5TYE7EkZrs//IYiVyC5VrB1
hYaC9kDmGa1LzLq4L6nBbqssz0NMVA3XQKO3n01IO0/DOD18DfvkbFFPm0KwyClPcZEle2kmp2PT
HmukIdLqY3qcg6S1cJFCHgD5RzdHy4Hc2gy/gmd2sHQ2w4bSH99KQWfDQrUdsKTD5WarI0UrjO9L
VayNELlPMA9NBLXgrT9d7sAj+3utWvF5vkBpnu4qsSb+3b9mM5Vw1yOAcHHppuslonri44428ekL
XLEFS36UOixWGo5RK79BmLaxCB9YsL2TaRNB4mtIcLcUyDU4KUy8y0vgYBNLlncV4HykEBjrqJe0
J/L2TTDOUeRYSypDV0tVeMt6CgBSZXRaGdBPNi8npNFYTtNxirHoXNz01dt13lpYLtrfMykt7AZT
mAMdXsO21Yg0Ir6B8fslVeNa6VW6MJpZjB88qMjsH3yW4/poA+RZySiGCbgtQis/Oc2uavPjJuQH
VC4W3PMilYjyp/YszNn0a7dXZbcWAU4zxZAJgjGr8RG3P6Ux8gifu3yYMNiygjZCfrfcdHmV6dVa
o6+tzVUfzksSb5UBe+5n4OmIzvqFvYfz0MZw0Z+FkEGFcy0byLGZVya9VSJBhTee6kf2YJ87sRaI
FEl1L9V12Ny7z5bvvg4yh1OTNwVuGwLkkFJI1cuOF8dPW1uk2sDvMpjzeW3caM5Irllpi6o27WUM
6MkiR70cQ3aaf8o4hDoNcwjI2nfy0sT/H/BoMesmvZoTvP8mtNMvNfF3XjFXbbcSK8QWncTapx6R
E0qjPHZbLm+O1cwC4eG+7khBBmOQ9MX2JxxEtsApiUOlz4hIzTXEazO6iWT0lqfWOUDPNGfOsBol
t4m6bc8PE62YWEOCzpHFGiQMnNraZWaW1eoiGoo0rStAjesvaNSHrufrQ7BnegYZiKURSTFu364X
WQjZSWQ3vD+4qmGlZzb0C8QyeL35N/+DFZaPnURFdxbp3H/QEsbyUW4YR68xsFCsXZOu0NumIPNp
4EBZfpbODyqTFUkS0W1xON6qXGuxlJf5or8GOFi1WFxMc0DmN8oo/llcqp3qFxo9QKC8K97lPaI6
E4p4xGVoEkaB6J0+Ii+OMVNI5+48Tq2M8D/zA/Wqn06aCFcT6ASl7GUsP7v3t8XLzIoNUPLdfG9s
QEba4nUWX5u0FEtsJInKR2fOWX9zf6zK0b5Z37mlW6ORVecrmrzeqSdqTFzSBJoSEXh/i2umXDkX
GRiDLV6Yil7K5IiM6fzR3itD9N6YAm93Sa9lneQ+6lbAO9I0+XCuzJYmuC544O05PYK+0IVTScD4
K8tIalxmkLg7BVTe1626WzaOTiolpjQkdg7bRNvh0tu0JkKHzPzZQzT0LYoX2C9J7w9xYnUQyYw1
wfSkSwNoRkYr2b/lkfvepdUGenfM1WTltzOja5W4RkFN0k3XTSDpLMPsW2+GE0IjQibv5TTu5NTY
jMMmHsEsgm2RqiHDieZXOwQUSx8pYDDsSmrDA61bF56LMRMzLLDRactn5eJFXYGwiGQt3hVDdCUz
Za2QwKK7jp9N3Nf0eiCj/nYHbmXUQbJa0H5zfKBCAl5q3jUYfctSx4mRm76z6aa7rDgPZiLiEsW4
Ty8FAcTnb1qnb6EzrfjZECXw1oBw60Pdyiwl1uAf/c0ImqoFdB/9LwIM6umn8lD9mjtfGING+rLM
0BgE2J6Q1tZeJw5i6OXtcsAhAoDH4abqVQtJ0a+Mky6zuWVlQsvn/xXTL8IGQiIVFNx3hi8PrkzR
9Qh0pOjXxk9c+mlwpBwHCA2fewtANenvBQXlrkh4ZziS40rWLy3+nkuQL0f2hhC7aE4hfMualKnD
42iXTKUcclXE82rB513GDVYaxvtUribk+n8QYPMSvLGMocNm8dpvlAJ/FHoyAj8jGuNbqTCECvpt
BDDBm+6KyVeSdVE4R1LmraWa4qMHVtpaaSRS2M1KGzS1S53dBj4MT80RFun9DB3EJIN6Lxmaevtn
fyYbxs0oiFk98ytwfSEc1VPm8pGplpZp4OmRqR3077yTwq2ZEhoqzDzMSQK32G76vZIMJjmV4Fg6
BTAm8vH73GUvFx+b0c9ff6ZJngwFzLMkOH5/fB4Q/hDu5UoQQ7txJ/EDgBQs5s1AGZ3jtDyNbBRF
sDZ/Y5tCnPmEiSFFDdeOwhrQ6jUgJzmsYzWauIlZaaLlvxFVK9k1NgHOF2I0oYDytLXA5FAAge99
GfClYy92lV7XyBvIF/24+OLZwkH7vsAmFVAN818uC28oxxMOAdUFCA/4C3Goja7ZmACTxoC+eRLm
CgTS3bjPcj21SrISDLgNVdMY55ffxUud1cKwrMu1BSfLB8LT+zvNq1DoeetDSKEuhrCBfBnr7Ih5
jgYGEv/Hwr8L39Taln6KZrfz96ho7wssWOo19f48oeUYjdGTmO9rm43rb68OYW8U9CN1nKWBGEr4
1Rra0Fiq87mngquJACIuW5EwN7D4qW/Cc5RO7rcQi3OABhYWYQ6GjXyAufc3IqwrS1n3aTSLah96
ZwBXjtdeBLp3h7ML/3ZpowLH6Q5MPIozLPkpezFTRs4/T90td7Fz2s82rnEpSFyB3DlSz7QLCTgE
379ac2SoCBgIcaiGzWbTVj9Ak3CRliKqUGaTdkDZQBpHHUdK5oRDYlRFGtKA7shDfV9UTiw1hCaI
rx1Hz6ADkUJRlu1A5jqB6zh10kuQOVgZVymvJwgPzvwDmz9PV7WkYPbwIWXbG3FZx1t4ugYElsNG
wtaUb50rnQVonHLxxN56dHEls4sY61g/k+D1bo5gBxVm1onXd/Jq/VUgbwQnm9X1JFtAQW7Jss2W
R/Q/acqtvRyFuOp4ETMn1ZaCSjOh2gHQ4qgruQKXNTSBW6RPuQql7gk/VoCvrEESs5IvdW1QYfTs
opb+Le+kXs1BlmtHoZqe8P04/kfNaBQfLDisLr1oDJxP+pz1kZhT459Ur1uX3SJOBp4iU6tfq77Q
EdowKrayyGwPaR+EiIH8Vx1rG5GxETcaVCWnMu8au+F+K47f7rJ8H8ajVUNu7bpGQJ0LGAxuzjk+
pTi8BdBWx7ToJWHnkGZe3dH4t51x0zeLeIy/ur0aM4E6B+y4iaJ0mjT3Fi4c1R9v3MO78um5vavl
pTfw++vwxz7Zrc92oHebnbAmEkjI0S43iMm5lwN/i16djpqy+vqewxb2Oh0CCY/lHpnilKPUEsPX
l2LLsMgZUp7yy/BoSmAqsqtDhRpUCXGpbIOrnHrkospSgzeF7SHNUfShguOekiEOep1fbrwpqoRy
7taK8ftaz38ZlNkYP9adt3PY1sNVujqlAuZWSiMajWY5FB/yt+6AmPADWiX17b4RSAOKgsjanQiY
fcpzTweS5zdDCRn4lWXNobPXvFdfsVYZV5yS+JeOvMdSLJIe3bsaE5kqBF1iFlxUYvr20ZLpGMHz
Y8/oUfTUQMp3aB1hPLUZS0wh/rVrESw/OEL76A5D8/ojY1x7a64V+qGMKpbW4gqOy3zWto0LL4/4
vyPeHSeM81Qn1V0/bari05gqTYrXl+hrfUHUX5gmZjgSfC8zvFdQWTMVUkkSMibB01/IL2NkWUgO
i7bWt1q0AHGjnIGP00XeyYco9b7ar9ZCAd6/U2jJ8bPsXEkEHufum/cMCsXgDuzPJs++M44XlCVK
1bq4O42sKrTBrAAEtItuV4KXS0V8mx4u3AJfPYVJk7lK1oXpMPDXxHzTA0WohlcYmw5dPAJMc6er
dPFQ8DWmISL2LPIqPPs0LPQFhodEAPLhgracEeqtLovxwyEAWVeE269I133D78u21BomED6Y5DEP
gxumLlgi4JnxkcC96DIRRF34ZP8MUYfeZ64EqFDn4aVkWoim7qJlh5QhauOHv3SNzLprNhuWx1QS
sSDRg0v89g1u4OSZdPugC9PBvvRqRD8URuu5bKFsaRDk23gmOW4jkmNhuwzfZbgOMKsCTje0akdd
BFAys5yN/KTceswq0jhO/LpYrEdSobjqNGOI9xds7nshoC+zGEiiWARIUIXOHKuC7C73DoPX3gXO
+V71KjTxwdiY7irBSdE4Jcc7RA06qEZlOc/utdT+1fQEIL/wTAVn+2RSbnZuzUUqX4mLmIOQ+kQU
KIGRKvjuPc8lEeMP+auGIF9dkycGRYyn5oARgOKs/8xGtM0L2OIr1OLkc4MPXX0fUhdW/xUq7sqW
g8VYpSHLRgc2GVWf/ArcmeTbyp95zbfya4EfnXACiEjuixKire8EjtESjahwsOI0QraJzTU2jvUj
Gzoad1yaq05dG5yC3HNC0O9twSVzYGMtN7OBzSfwRnirm0zo8dFexLfLW5PD966eUiSmMEvj9Nae
w3iWeVUWVncel1fDBvt+k5cFzgIape8qt53D//4bRH3iBlXXi25tJWEN+BtmAZ0kHSMfUgvU/I4q
2xh4xW/LWPH1OAD5zX8z/mc94WJOOaywZmSx6ON0efH9JUh4XRai0M6gmkD2pG5Z3SgIgN0Bnj7H
gwNh+FantRL8VRUTptJAEo/H3ncI+aawG3Oco4blT4YrGBiX7xsE/nLn5fA7gUC85loGzB+5rMS4
JCw+TZ6kGh55pzjXMIoKFmPy0nA/bqBh+ewQJQSoCyNDZrPhtfh4TSNS3FqoSpzF0tbEsY8qlwV+
zY24Kf2wz+Tz9Q/x+Dq4NpzGMpqZH7Cb8kcHn41Ba5xskI04bXwsW8BFMH434vbnsV7NCeCDP9FC
8AMWI2wqQp7v3ey4nK1kQ1I0/+DkWBvwrVk/RApKqwDoH4wWBVHNSmym4bgbO8RZsyMOU51IZA3S
WHWVmW8G0XWzUgJcrU5KnXXDwcqiAtsP4KCCqeDhF97MdwlmzddOkAWVIdnxLdBA0A0/1APqd7mL
lP3C/pkIYWfzRO+kgB5+vIK+kPpSaNHfQacY5y4MEgYFKmv90R9EJAEvdyrc7iTbHx9IS4PRlRRz
phAvOGJYHfJAqK41XmVYwPBWF97mr1gvd67w0Q2IYvMCI8Km/ZoTjo6bArUTps/vBuXfUuydgxB8
WsffoqDe4gAPj7C/ALYegUUEOM8nbAvFqune8U4zIuODhLP3qRibmkHd5azF7Rp2MfAQnqDnDQQJ
tP9P9baIo+NNAn1PkR//PZEToM1ZTfljzEKxNppaE/AKLiwZtfpq5H8OkzYmsTkf70i9w9Xf4Skp
OIAFRq6gajG4IR6uH7HgJudVxCaf8scsmfZBo33SaHhhzwrL0R5ejqKX4v1KPT72ASJB/zKwwQAG
7qZr/Xex/bJIAtmXJWWlsR4rcX8u+DrS3ZtSu78XkfyDnYiwIT7LLaoaf8YBvLHtKsgb+bD6H/PK
VQHDtMaRZZ8CSddnzxuc2rZD4mqzlWvX0pJrq90dDHLevKRMLAxZtIV3kqXoTvaAmj9ee42t7t+5
E/6BQRkbgydGM3rjFcYd/q+zDOni1OIhfraAm+3GMr+QNj4s4EnAmJNXQ1Qu5MeXmoHnigo5co5K
274GD2rQLTrgdDz3thskNHayv/ld7dsSWpJfhqZs7KUZyxkItKT+b6JLonw2PAGSaIsdJHZV78Sw
iQKU32PMZhMIyrZgUs+Ov8Sj+wg3I+zXGn6ZHJxCqwvCXgKTOtQ6EadnQsnoI9Rz1dMiD3f9wQeG
9iZFjQxvUdIspUIbC/v5Kw+fxJg25tPyJfOYftyOvEt2M90a25p/a5M5ww2vgosDpEPxzIED+XSE
76N61hg3REkd3gfBsW3+MQdb7l0loO7le+qC9GRjJRhGNb2MO7llPWfjhOY0qIyIM+IjgW+3Mcrv
CV46VgnTTn9Cej2OqdppZmL/uPq6oAbvgvQ7OR1fWpTAu6GffMlrcWW8xZ0joGjXNXtF5D8CG9Jc
5KHD0fjtjN1BBld2eV3OVMZtX6KL7XMmn94FzumbxhMEKZHRsmDvukx5u7Y8ONlDdtH0E0Z2HB+6
ZkJxCgujUTWko50A+J8cmJ0dCD5xQpgZXjqNp8vx6Nh74Mv90GdGbzTZhGrENw7rL0G4MG4+iOVK
zQAaGi8AnpYY0IZCTY1eLjC7yG6TH1I7nbJIew8cFnyJLP6U853BliWtMZpf/XJPyOH0BeLIFt09
QtTrk8AnfRVblZc6XXjr3HJ5yOX0t4AMhJbbsTDK/8FYDs3dskXb76qXxa0O4c72NhJJOuJyVpoC
Ul6H/a7jCxDkIZksl7YOCdwsZjkLsXv9EG1dq9Ad3FVYI1v6Ol1heC8BCNS7IKvFAKqIkb8NABhJ
4kmMEdVML4XIMEFf/Eadmr1jP1rVJWNGEFkioec+TM7YZGZiQwJyYaUy022M5GTUX4uIC1+RDkni
uyg+DXI6NJZECY2ZdzFJmRu0Rmw0k+8adgSgMhYcC4HcAh6iABD4Keh6Ufi2NMmr/hx3xoPGzzrj
+l04PwvSVvN6kRGFMp+zUh2VyVS8pOoz99dupbvu7Mj8s4Xj9gQ5vkO0/VSFeHOHw1sYktF8eZq0
NB7npUvgxUQyTYiGJFGM8mFBW4RAkqPyn8EjF9X2gYYUGHQsbBKXGGywfPslnuxWhKSKdvy3pq9B
COJbtRODaAgmRfaqAMGHUX0hPbaZH5iiTlroAZiK7f6dINBlq1R8QUp/+GRdcDTkYj0gRbx/a3/K
n67XN88EEoyPgffTdDT+zzVbB9ZB79q8p5+q+/E7d7lxh0cFjjQocmYhl7n8LOkmmPAmGmKhjmUC
pfENTUN4ngSu7A195S4lOi6WjSnEJsS3hcGM4VG+DXngtMM8k8oRfYExbo9l5mzzY1dhsFjhl4Kr
5tklbdAMNiQ0ug7sPw0OjkMxX2bQBAV5xroZv5qv7On4dsZC9fAelWoFC/zNxu962G2f7wi3M3Vj
ioqfnKPaOkfy0FVGqa6QTphu56wfmSBTdA7aaNiNwqYtcN3U2Vtg/3nzxoJNRyPaDmzS3B33KZ9a
4dPE5j+WQA2HEyjbLXCFQsEyeUdeVEN7Xz39+1PoHX4W/MjmpIU3Wufh86Sx5k3JjX4f+7MYEf/S
S/fA7bwsL4VGVpUUcZnk+FducfSnRm2cON9CYicY1ZBoW5vghUl5alCg6cxXKpxvDoU78gS0AO6U
GQP4Y0OMVYIGyBWPhj1eKbolyQadqe3SFNs6HxKrDeHEeG8icOlPJXywfuplP1ks8vvmnqv3AEAk
e2Ckt7z0flGf0GSz6cWJ0CQFGaiEB9U0X9MkVRIC6DzoMSMsGdjoas3S/nHVTcn/db7p+Ds1dDxK
4bAAm9vGmV0m/T6oJHdSre0Rnou5PBb7tfMqSvfWNTMjhKlPCeQZPjUYm9xswKvUiwyHksTqG8lZ
+gxz8qcO/k4jhwItcKVi4R4GCu7PoCO4C5iMZ/xh5NHB7E1T3Apc0EBqwUvb3czxrFBgswSwg6dv
Bw6qoDytktXsXp20hBJFt8mwXsey82X2HLHpWowu14u3d1Z0w53C+aM6DokK49ScoHJIrqBt8Cov
XDunuX0VVQAwD9GoPXIVqepNp9VD8j2OU6dD6XO/lN19c/m4GiSPnS0RLkM7xhXUQdhok1qHfe7D
UFuGGJZpvV+JPS0hN4mFCt6sKMoCLnlP+tNtMOOSTlq1OyFxyHGd7v+yBdGPgzaJDs7vPi7fEqKX
7DgcIcxmdRnQc//xEk3pnaafSfye3aR6FVgcEKdpLglkcO+lKAdNt2TXRtdpupRR+a36ZlsvBbsK
5faksb8uOEMoA88/kXxnHDobP6BLc/ypxHPLQ5Ha0+6fUmVvBZvcVo33S7qt+FIEKvvV6G5quYWt
vrKuND4hhK4WDvVJEmZV0mDXS9XgvYpCZGDwoui+RA9VF9XiOsIgbPSZFS6Ak2f8r/wfIdC4jeNk
i+qVdUL2Qh64A5GAZadeMkE/KQlbbiJaZQomwabxlj2uBqxhlYiP8TLyYj7rHmyPQLvihU9BMvWk
IiNvS7nQZPI6UStEMR/VLablBdPPpZMYPtcBq1Q5d5D1DDhDBgyhGvetE1/Y6p2w4jhtvoNtxhPb
37hPYVKGy6prw3SsotrSbuyqDjWJCYlTS5ojo9tJnfw/N/Au/Uw6soJRMB3BaquEWPNaMajXYoEN
lESUju0sD+rDrI6vz7oqnFjzNBYP+g9zhHhZuv3SxFEl6ucybQe9zb4nc//XXqpLmRLouklD99TR
M2YgqBClE5Gc4qUIAZUFXVop+d91z2WeZqx/ZTBBxiWSp/NjIdHC9ej1rEQchEzkCtNDmxeaUQAR
iYSrNespgW5C9/NeykU74tGpjCVsNRbt5KlVH7hyehjI7DnL1wpTXX3/fAU8gMB2trWTNX/P/pB5
EslzluNiuIyLbstDyePuH//4ZDHypuq2jFIV7e2B9quODS5nwyNAlcqpnuFOMziXZqG13l7YNyp9
oBDU3c4unVVaiLrMi2DyLPq1eUrqJcMDTL/VNmTvd59+ixXxtOGY5SERZJo+x1y65WySfPxP2wSf
JX3ruuvVJl86uPFELwPeuC41Q4jJ3WN2jjA7xrgGY86nwpSH8bHiHVlqlom4UiE5BPN0NDZuqmjz
rO4xh0pT8pc7ELvywcjikRv5VbTyNLD8PSh/76b3xerL92B8u/cYTeYJS5CHu9shsWFIDVAPpkMf
lIa6YGb8C4DiT56xJQ6IFdWXmq7nMQSkSCn186TSGzIgpCBUgA4KKGK8IBdzHDgpLNU1ur7GLV4o
ZdXhJx1jeEccPaYiUtzOkuhCwuIqbVax8naHQV2BidXPd/VPnSLEmPqnJ4BWJ4KKXSznY2NoamEr
LhtoDsvg9Z+/g2s09s7Dwe0o+OEYGoVZ/zqSBojPq3wusSsevJ/1wrkZBh988R5LqSGeZq6Oxzt8
xGvAccwCVlxFyg4xsEiz/Y6ueikMNUwLqhbsWMCM+j7RrlyYSuumAoIWaUT97WkwPErJS1vbY7JX
GGspRu65sBMvXBlqpThK6jy81yRZTCXI5cv8PMEbTY2ipW9WqB6dSGHR5QjPEBzxrQHSdPgydqzs
AMt008zn5m0XOoIuTrOrDPAZd8eZlSfuMY8MSpiBYHfYmA2BtuOJIzkaIMIk4Pkkt4tE4zdRfoB5
4cgzHD6sTMhnoAXvjAsdVuucH+sIKBFvVsFpAMMHp9ROBd3NJW8AXgH0V1/q3Ij4KqBNLoQKA1iE
FaTdOTeGYJPsS46xS1pbJ9UE04d/Qp3C4GqI6kySdY2njS76B75IOwfmdBVs0BCtK0VpvaVPbN5t
DbXtkCr9/H2++ryvQlXk2aPFx6r3pL/CThLRbY5AAqf1+S8mB3YASvLtdMn+GdHI57H8lHjE9kD1
HOHfospXQZLjXcvZ4LnjYPCqkCiic0pv96fpXhIGFiQ9e2M/Ldg6vrBIyyMEWA6EhaQ2D1D160Ci
gvfpAdTgl4NYdxnxQKKKfNrfEcZGURKAXKQtZyduaCXFAJJK82LqJIIpc4zI+JAeGtEK+a5Hz+pH
ulZMl+tNR+jOo00hVveyvTkG30r3uyZtVfzr64dTidu6bWRKpQvbRmFBxYOCrEJcLpv1/o+BYJeu
ZNsw5KiQmM2vZz5+Gju3D7iNjwj2G4RvH4b7ySXLd2IKGGOkaotxQRM29kHuWavlC6npWVilO3+d
AA8IlvRJHsGxRbpDfuDDicqe06DuE6LfQMNgeV2Kha4gcCKrk4k66T8aubB2uCGR9PCnpWZ4KM7O
on8rVfcWLpgdEl7G1D0hb3KEIjVzUVbP5iYfGUU/upbTYxiEDzmWsN8mZ3JWopWhPDfeSslKUo9L
/6/Nc2e88UY+Q6htKKRaiMUPl5b9hg9AkY0zQZSX0II2XNB29HODGTOOi4/W913DO7Jeggm57USO
clJdxrqGjmELoKURB9+nbHYBxBw24VAHmyjlRLIN2Ws49SfBl1MysmlcBdW4o0PiKgONnuMy6kbk
vy01yzBdCtbUqcZWlq/Fnh08uhSb7VKUBTPcVHM/PeV7xhNoHh8gdD4mSAVoTcnprwUcFeeVa7qR
1tlfpp+m1KFIuwiKKUp4xNdd6ksZvVM1WoaVgQrKKWSSaHsQWK2DAXqEuSusqNjbpw/IfUeUXjcx
u5PeLdaXtSFbcXyWXbGv3mQLH31a+0XKZXKkbxCNhDoiYIjyIUsn9YwDTawxw/R/JtRrtYYBL/GW
s3elTNWuDPR/7swNI/aQMspsBv3hrwucI7vY7EgT7S1Ktj10f3wXrvA3T4YwMm3YvTAC54l2DZGP
rYlX44jCORjbilguFabK2JHnAcpeF+rh3U3gyJUQ02N8AKPkkOmQqSDx189TR5ru1Dk2XY7StH7P
Je2I5XLkji5QpdZ+y/PDSGPFY2PLghrySzd2mXY+02VEIAbe12ZFA6/mcTkbC6hEJqS+LayKpoHo
NSaq5IYPRFB5keF38WVyAO8Zwo2uYylwVVjUKDHp39KP4eBPQUrJTqKBGFEkK9n7kt0u7ODCgmBI
2LbwgGe0mRsxioKEHIAn68hZtgXbJrSyjM1NJCAn/hfiSfgRs5QD0VgPwyF92DkLjLGN33MxagiJ
Mxz9A6rwu+LWBvwK+byCF0+wvlFTbf3XULABKdCjim8t98VvMxQF2iizvv6gPTKZSHSrfugOzuJF
kMXhIHiWXjjDQl6w7pXyerk8zF90gkLA+cNv9bj/zBcffr/3krdQdOpF6cbdTlzxkkFK3QpfyLqA
K5gKD0mb6X9E/LI+uKyHwfdfyCP6dWnhtbElBZyOZYw/G0WxsVQPPVbiR+iIgvEGAtVs1I/rmHqA
0eAYZQ9t9FNx4Sf1lOYB6SCBsa2xZl1EZPpB1iInAs1xIXOgpHFfH3LRobT73ONuuIvqTGlij5CK
lfj62jVW2bMERXMl44iddsvMWd19+Xw/bEZpyP/BFnZaTizkRmvPoIUYwa7qdOKm4HzneEUJaRvg
iQkf4sixnRE9JDW2naZkqC2QuVNyfhvep60T/hNTWnW0jS8XOvunP5K0WGvCEqTJh635cBdY7HA+
xIPomTDofTHmTFtiO0o0hoNCWj1IaxYSW4SQTSLOuwYM
`protect end_protected
