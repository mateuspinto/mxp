��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��Ь��-p�l9qe�p}����y��L�Xݳ�,du~{�/�mt't��UUe
�"WJ�>��.���as��^�o�r�?�>��{�z0�2|K:��lL��+�4gejCx3V�+*��$���$>n�e�*t��I����5y���/���ͤ0�&_�[�ڀ%'=E�JZ���^��Y#״i��\Ce��噤�7�&Я%�
�r��ESƿI	��!�"�XN*���8��X?�(�������=�z��Hl1NE|���qכX�ʦ5�C6��7������.��ۥv��6É?�%� �.ۯ��<�b��r��`�x�����Q>�T]E��������1�S�J;h�nR���D>1�B��`��K�$����8��b9�zWG��9p\����$5�����L���kO��}|��:pڿ�wt���f�,�2���x��
�{R��&3F�CQ$6�#˦Bξ�T����{4>�Ё1�(�%���9I�E�bV�b�F�j�m2���;r|o=AYG���jzYI�D��o9�?tXg�?�lO�vef����uX`�GaF��G[�����M(�ФK��6j��U�������D`�oBS/�@C�Ӷ��wd��'zT*ʣ�,��>�ۭ���^Ok���_����Sa�3��1&x[r��t?m�������X^i�b���~1%""���ĎRج�;�����b�#Mo��+8"Y�2P�M�q�3O��	��%��$o#���s�q�������|R
:�	�*�I���{���v����Qnk���REI���p�8 �j"K�)�7�@�Bh�lD��2�u��0�
R��R�dJ�r�/��8�k�e�o�m���xR��7���^�|��p��s�ZC�_��gW,��|��@��H��ɾ��1�-�<ݣ^�!����inCne<�2��A��4�� A��DЍ�xPw2a�Ќ4L����I����Dl��tNѡ1�����;�����y�%�賃�G�
X-���(͞����#��J!o����#X�_@�\1�!GY����%�*S}�bl������$�!�He�~�cIJm1Y-�4W�y Tq��֝�m_�=�h�ev��\�=�F�v�ه|�8�'et�����$�t���J�:x+��/�
�����g_
Fꌳ�Z��bC�I?h��ޠ���-͏�ta}T�"ռ����Ɏ �<#*�-t��.��Mi�E��P��×�	���SB?:R��dV��t��ρ�ɨ��e�6&���>~��h��8
b��;M�RYME��4=���x*E)���l�o��D��>��Q�>G�c)��,i����F���/߇ۤBH�J�P��&;�NJ����"2��z�����M�D����!8I8�� �$��f�����4B��@��j�4��U=�*N��fډ�Y�<Z���(|��uO`�H�t�u���Iά�������m��% 5(��!���eX���{��S�`%��RDw�,���*Z��M���<m�?��J_V,�/ɮ��<^I���=�?r��h���8>a�'�23���\R��[�/ȳ���=uAH`a+F����B!��fU�?ί�tA%��?�)���9��P`	�:]���F�Z�xkL�0�(�p�j�	|�5#kn%�e�u�_;�k���Д���"���֗��%I&rp���:���-���$��4��^Ga���7	���!Jh�E
��D,Z�nJ�uR%�ɩ�gf9�E��1
��4M!���B*�5&V�%0��2�u�R��l�gR��X�p�NUc�� w��
.�#�&1@��;���	�D��|l��(>�Oj���Ј�]�L�BQdLȟ�n(I8�[xU0z�}���N�C�gQa�X�y����p�Q�`O���2�tu�'6�R��*���g����kx~�hl8ϗ�ʗ³"��7.n��l��&�u��%�t�����%���G_ظw���mm�
���8ᯭګ�pe�U&6H���AҌֲD� p%h��������*B�x�IgxB��ݡ-6(�N;��l~��
�b�(��ҵ+�kM�q���)`$f-t�?�ڍ`,$� Z����&�z2J��m&D�m:�=n����n����Nq�������#9�Ea\�\�o���<(#��%�Xp-3�!V�$="İ� ���q�m	WB�Jb���B� T>!܌p��OϪ�ڱ��F+�IU��9{�N���z�q��6���z�'h� �$#��按d|�"��-x�P��8Pe}	7��ڮ�Qlx"����\��3�i���$��#�	�*��i�U�9T�Q�4�?���f����U;A̀���Y8��e�]��H�1&��lpt���
쌑��H������3�`�^���� ��a��B�����;�I����l3�d:���5(�Gk˯!� ��Y;�WLP�U��T~����q�2���II��wD_�SB�&�Ô<|VV�5��
�i������pW�L 6�ؐ�R���y:(a1a�7J�&#,Z���q�"t�L��N�]�2�T�ﶘ��x��{	ŧS�u<uc�)-L����72f┹&G��8���݊[�w�i�	���>�l6\2�+�J�6�ଣ�iH�I!Br͋\�����y������ED�a�����Ҋ�R;%�_ӽ�ڇ�}_C������d���5��^:�k�X<l�N�-E�����X��
���STȑ�n�2}�{���hסg=����Iϭ=?�2�m
�C������T"�F���C"���VE�sQ2r��'�^��]m�&��]��*��Ɂ\{�+��r����I��+�7�8������F��
���q���np��b.=��w*_�NYuW�S�&��fB$V����y�yJ����f�Δ?w^pBM����`�:2��D��J����TN'l��Ң�J����F��,�g��09(���S�<c9�������*�������E�?"���B���s,]~D)8�8���;� 0�6�Թ�\�`�qhH�Nr��4�S^aT���_$��~��o���f���QL��j� �4�@[�T?�	��v�I��_m��T-%�+G�pq�F�(���4#����)~�8�F_�y�dR+���k�qU8#�Yl�3��l�*��ʘV�4��b2q�0!SP�t�E��ڮv�m�L����0��,�8���i挊z�=)M�_�FL�����$4��+���!��Ҍ�M�Q�5�(�uh��u�dI���\���½]R�d	:ց)s}Ťb����Kd8T&g��'���T��+��X,A�ٱ�|:��fm^���K���[�b9�m=y��œ���_��G�G7Ā��v� Tk��ݗ����vX�eZ#�}ܞ�zr���‥y`4�ub��2`���2y��G*���3I�(
i�\��j�B�%? �.�H��iF��w˳�)����>�Ӿz�z~e�i;k�fO�z�|�;����A�b�b��`��[~����ꖭ�@q��pxaC%��YjUipD�������rD��'>��S�' �f�&ڹt�Q��3�����.|�L�IaM���N	�E���ǯ�	�NsP���}�
�9#����@<�� �?���WS̟1�s��I�H�t���cݿ�KWlır'	�s��Qb�p܉�)�w��(��
�R`�/8�+���yăp4j<���H \0c�G��OEm8	.�v�v��-B�<��;����B�1�.�`c�����q&�ʳ�!�J8���K���}��ʮ�����;eҵ �"+6�Q���ȏ�	����͕���cY�
���g��O�St�����$X�	'i�(�R��[_}:�����sC�SY%
��ϊO��U���6ko�6�wrJ�-T`�9�D��6^,f5���{ ��I���;�������/���1�o��\	�E_4<�0�8��J*�}�v;�Vu���$";�+	T73dm3/���1~���H@Иio�%�ra��2�8EW
���y,�خ�Wa2���V&(@��|%Z�t�vM��}h�1��H�Le:U���;iЧ჎b��-:����=��_B��Y/��넚[~>��0�g#�b���w��<�������P���n+�aiN���a�����9C*4���ip;�|I�����,\�MT��"��&�e�a@�����G���o��[��տ �� ,fe0��I�d�)�� ��3'!f���D�W��q��8Jw#-�瑜m{Μ]X��$�����R�8���Bai��d�L^p�u���0�_]99\�}�Kb������$I�����o�)'z���R���8D+H�Qh�ꅊ!�mt��v������}[Y��]8]I�`�!PpN\�ZZ��V����&��ġܪ�H{&4��e��!ɄO��`P!: r��2Šj��5�|ŉ~|�e��.��h����ɖP�h�B��d�.�l���t'h��!�P4��!�p��Ɣ�	�g�]4�Bua._��t֎��@���omL!>o������j{_�YorsD��9+�:����X?m,a0��t`ͭ�i@t��@�Q�?��c�Ϝ��a�A�M��X��y��-���_�lK�zhИ����RY�"f��Gz�Jx�M�� d�r3^bs�3ѽV�
�� ��a�nQ��aq-ҦQ3�ie��(?�1�UX��	�,�i���6�*�U�Z�b�l��5�H�N��0�YuJ���,�`�����	�51��a� :��b�Q�1��zp�Y���c��p�Ч՝D���)ˆS�ǋ�l6��d�ě�%�#0`,=����s��+*h�)�����EG4A/o\[-�7������xsC�R3Ui�9/�C&8W��!��&�2w=x]���ڃT�!��~���N�O��+��A�J5�4l�~��'1�=CT����������zSV�6Q�*�Χs[V+��#���x�Ժ�m�#ŮW�h0����%��9��O-�k"����N�>d�)��**MCq�0��l2UhЄd'�E�����6�ӗ5��6�S�b�xt9S��0S��n�d]E�=
G���uF�a��vy�/�K�5���[��[�)�����»�J��Cg��x����A�a6W�\[�h��Ƃ�'�z�Dΰ/w�$�d"���eW0�n/��x�^��i)�[��U7�|�[U��I{n��<�T��@�gUh_�&�I)�V�z��[��r\L"�_5�9J���gA�*#��X�B״+�]m)� �oHXg�۩ Q��^���l��S�sV�h7���T� ��)ڌ"��ش17���d�~��C�=riP����<�%���ʬ�FK���Ł�:�0��<=�J/ϯ7?p.�p3���ʻO�R��I���́Un5�P�ư�<ن�U�������<�J���Xп��ϛM�S�t�Uc4x���H��Jy<�kYKL��J.*�#�Ҕe�%�U��+�,��H2�?hQ���9���왝I���X�� �4�X��%�v��[�@��Ӽw�'�L��:���]��5u�F�Cd/j4x���Z�0��M�ݮ�h:$P��e9��3Uk�k��h�������^��tsۉ�����`,��t��I/f��O�D�=�|�}���ǩqq���7���xV�9T[�]��/��nd��Ē�;�|�nX�e�83�R�"��KT���c�:T�����=�=P"!%O�U��tw_?ǈ��K�&�DQ�ju+�J�<��ق=A��5�m]�T��$�r�SY$3볠UK�?����"�i��J�!x���1�y��ɰ��A$��Z���A��_�Ik�&�@�ێ�!'�B-S�����(�e��\��+[��X�R����.p��IE������5#/��l��2�K[Qd������z�>,w��Bq�w\?���t�R����M�8B����lD�6���TqE���:�*���]�[`�@��u�E^A�i���8é���6^X
z�䣜l� ���O��2�M�*.��2Ό���:۰˔�!�@d�	!_ �-+}��#AX���~���>�"s�Sˊ��@i�tÑ��c9�R�I붑��l����RA�28��N��C���a���~�\����2We�1����{/��bh�M*���)}�Iɋ[ �}E�o�%M��*��͕�?ܼ��4C�����
t��H�w`�����F��q�'�S�� �Sr�n���wW��5�q���"4��iYo�	���u��j�W������#t����%A!�Ω[����)��C!��!s�e|N�����'��{Wp�0"ڢz�N��^��p���G���U���� �}QT�GQ�.�(*NA�C^!�?�^Bf��>�ƶ]����&����qOi������UO�Q���|T�*s��	���B���k�2>�s��x���u�4s!&V�Rtc{lz�_�Z�^H%�u�3a�b#�k���'�	(|SB��E>KA�^�bӡbf�m�A^��0W޼&�R����z ���
/�S�}���q>�t�Ʃ������'W/�ݝ7�Z
�QpV��:���y8��L��>�_��Ÿ��
d�R)*uwn��3�y��e�{���m+%��xX�i_|�E}�N�M5z�~��ɽ�yd�Au����,�w5��%���hO��0�D���E��X�)Wx��IM#��Z}��U��e`N��ᕿ�^�r�۾6ġtJ��*Û����"\���n�?+��,��ϔ]7�'�.�̚��<Z�B���9�I���zYĊr�%]��7[}JA�	���=C*�}���������_���c����U���!]����FK�'T~�ʑz���;C�v	�V 6BI����b5+�d��_k��f���x�]���9#�٤�wD��-6�6~�Va�3G���O�V�'���}=�0%a�fOHVjb�,9u1YfQS����	X0N/����>�Qʻ���Eh(@�/+����џ��)e���m�b�]�Ɏ�5GPΝ���	��+g%�y��l���{_�ex���*vG�W��D��ß��b�r-��sT�t��N�P>�w���6�Of�^~�1���i��]��,¼_D�3f����9��We��zw�Br�]R�T󶑢]g�䚃��"�ϝ\��7]:��B��I�x�TL��8��\X�%��sr���6��s@���|^cv9j�FHJ��Nŏ����gYJ�����^j㢚a{������L�]�ݖB:(W�G�T���O��)� �8���>K����y>o��X{G�81�w�k)M4?�������2{�D�j,:&Z��!C $h��5lt(���ruf�N��_Ew��O�¾�4TP]�*���,Mn�����<��op�bכ_�F��V,}��:���H��$WW�h8������bQ�na͋^��z�!��O�T��E j)�,��A��ޟ��J�ٶ���]W����@�I�>�72���D��'_�	���u�|.48�ߥWOt[��B-�*oEvg�,�)�1�r�I���+Ɖ'��Ek�W��a,����(��fG��,)n�Sg��I�e��TY���(�۷UzEv�sV �ka	���zO�^F��wH�f}"kB���:�L���]�#�t���3��`QK���r~#ܻ��
��:�Lf;�q����Τ�l�mG1���M��r8�g�ռ���׳������+�@P��C!�����1KKM,���bf�������yCbѩv�B ��M��]bU����-5מ\J���v�u���!�x�ĕ�����`%9?��9`��(g���cmxb�c��֣:SY��e��j�v��A(���.*	���q���U�������N7W5Z֮+=�8F���N�GJ����3���(�I~�l��2E���}��{jG䌰��쓶m�l�?)Ѽ:2\ �<�] r�tK�ϗ�N1iA�Q��7��b�T��2�.C���'�uF��V�@��3��wU����\��x���2z���W�.&�x+�0BW�<'L��D��l.��+�!�����:0}�;!�,��*,)�wL+wU9�8�l��� ����J1,2IJGx� JcM����������@��<�v�M*�U��\'�i[�N�k,�54�E���v��Ψ�}�v�9��m=F/�t�d��ȅ��􄍿�ϖ�JQ���cn��YPE�+n�/�6^��?��Q%��7�	kh���E92D�(�õVy1�\i>6�YF�Y�'Փ�t�Z18���>C��Ft�H
�=����erc%ٲ��؝d�n��q3�n���=�ߺ�v���#����P�F4u�1�<�E�a��W����}*��~�8���b�l�j�����/�8jV��bT��8��U1�� g�s0qO�ko��6��W ��Qx���lۚ����E1���;�acВ�z֪\�?zI�����l/���d�T�9K�4��#Q��v�Y��,�j���-]
��������|j7�~��#K�"E~G3&ǻWDo�er[h���9HЌ��ϛH]:kV���1�lC$�q۷�����c�穎9��)DB�ջl)Z�Fd���o�/gwZ��H�����d����M�V\�MH�T��A�\�V�T�y��I���u �k�}&ժ͂���)�����M��o��P���XI�aYnl�loN�����t�1��P�q�3��҃d˵��w�(���X�E|���>Փ��e�C�(����Zbu
0{�������+���J�oӅ}1\�j�!�\ٓ�=-,�|PU��u
�6;�~z^����O��-��:���t�܈�kJ�r�Vi�7�s D/�X��ˁx8ٟ�(�����C�F�X����H%E2�&�D$��MSD�
Zނ����,>6J;�~3E!�|�������Ň	ȃN��C�,�y�ѓO�e�������Z�%ZSmD�uH�l��3Z��#�]����{I����wu����Φ�0OO�b;�;���j�'�[/�5�6|uB^\�gtm��	��=�d9f�ƺ钂�k�&H(�:���>����E!��Q�� 28§$��) f� �C�Vɓ2���r����.�%�K����Z���v5N��ý�2��f���F�74��v��.s�G]�ݍ(����uQ]�UbaFj���NN�l�u�������K<�(��B�Z�5�YM�o#��>��Ĭs~��oXv����tm���yD�S��<s�>���#F�!vn4P:���+^�[�Z�P��&�Pۯ�X	͇G����z�.�ׯgD%�U?�x�	���wd��K�m%Op~�^)���\Ɋ'���j�M%��c����taKj�1�J6�L�c^������6%��c�H=ה��\t���tK&�+^#p�I��k����M�J-E��D�#�Ү��W���y�idh�n֝~ߵX�*����m勅ɼU���&����111iY�WE�R�P!�����ʠ�gȢ�s��8����C�	�?4��wZ(!�
=N�6x>�?�1z��`�O�CO�����V͝d����LH@�R8��4�^:���w�H6�&4�i�OW��B���q��H�м�L�C���}��� >���k�vD�k�US�4OэG��5V�< !u�o�4��V6�GZ�	�!��:���K�p��3�_(���_z��0��w��k���ݒ�"���`�'r�h���y�-�8iMІ�<%MAQ#��k'�ݬ��h\��8儴����rBp����_�i'�	�o�:�m�����	\W����PO�lvct��F)u�2Ȍ����Q�rW�6��^�_����vJ)C�u}Hԙ�#R�Nt�
�1�4�NY_H�8v�\y�T[I���4@���>[34IUH�L��6q>��r�tt�����;����w�W�'�k���` �� &#�Qk�?���L�!Ѻ&���I���K��:���;֝�x�.s_ђ����"Yh���֊�d���������Cr�2���v�l���҆^��q1�PT�\��a�%9pJ���`�S�fX���eh�A���_���L=
�%�h���,#�A���ɳLx�%���`�Y��ͧ
�e ���ˢ��b��儮`�`:c<�)�9�?shk�L@M"q��Mz�3x��)g��ޭ���%���Ȑ�b�EYoj��jӴ�&fyQ�-�{q�!�}��ڪ��c�{�2��z���^~��Q��L�r����v&2�2�3y�k�j������1s�n���AF}�:��
�x��9�^>���Iyu��G�8f���ەӤ� 3
0��9���q)��#�k�ׯ����T Jf�� 军\�jT��! �>lgV�E3r�?�����u_�������م�Y��r�<,�	������R�Y�܋g�$ѷllC\(�ys�{��w�E��Ga�2FR#��"�X7}��A3c�"�V���%w�p��Y`+��(�OX�/��B����R��n^:�W+�������qsu��H{���EB����9�%�>�~����6Γ��X��M�ƪ'�\����\V՟�n�~&�,��N�Z�'��'�£kR���s��e���)��mz/-;_�ʾ�x�*O�ڿ���tXH|�Je8Y���-����hmO����rވ���B���%���$�8�
�ՙ:ڜ	�/_��CL\����}d�#�L"z	ty�c�	d�=�۝Q�O�1:�sm���Z6����� �ў����X�Ї��J��t%Kb��'� "����\KĢ��s��uR,h�(��k-a�y�^�>szǑ��V���Z㾗q0�"].��������j)�b�p����u�MX��H��Z_G��_꫊�������?�I�b]� �.?�i��q��`lW�}`Sm5ȏ'�F��-섚����Kc�E�F$0w����I�	���*�Q�N�W��¼���
�,J�J�{�B���5��n=t	V3ST���� ���#��r�iOim�����)�Rz�m�N��GBi��6!����ҁ��﭂LlQ͸4W���N���>"�^g��H��F2��7��2 ����U�1�����(]T������*���.�b�u9`iGX��28�v��O����������M^Pɔ�%��i@�=�q&N[L�C@�"�]ܸ�`G����6L�uf��i�c���fp�6xU wi{r|C�����x]�e�2�́�<=ؿ_Qܕ%��p�p�����Z���������U:r-a���,nf&5��ח��k$:~SBRഭ,Q���h]~)����&�;U:p��~����+i,��_SC�]�e�$M=G�r�W�i	�y$��ƾ�"ɽ��Mܒ(���l�'w�*(��G=�����y��&�`QM3^YS�md��̫X�b�b64����4;�Zb�4Ң����߃�Hf�zkJ��'79#
��r�k�}ޙQ�&L�S�K����E�Ӎ����)���W�/�p$M��q �����s�mC�X1��>x5(:V����]~��4����״o����L� -�o֖N�2�g<�sm�������Ѡ���:i}s��_)��B~����ϐy*���7��cHI�r��ka����ut8;��r���5谆?�Iԋ&P�1�m�b��]\:L���F�B�Y��.�6�QK�,CUW�6�@D2`u�Ў���ј�>�m�#�#ʙ�iqݢS�	�ߔJ浕,ڳb�H�T:�_�!Y��/���L�͞�d����`
�^GN?|�uް�+�o�L��@�d�F���N��[����dK2`�D�9C�`�J��#�<���omJp���*,�mFQ��M�c�:VO����f������D�%�tU�(oB6��~Jq���<�Ƴσd���?Dz��G%ƽw���d�b�2k	�'����H�"��v�.�
-]n;L�(���K��N��=��t�Nx��z;ٶ���YU|����e�
Iq���kn�u>�����A�8���N f|��^
uU^g�r&V���w��)ZF��6_�{� �-��s��%�U~�Z��i8L*�� x�0c�X�a�sC�p��.�e!H�(t��nI`-j�شm�)5\���W+ٴø���S
t��Xk�[��׍} ���������Ak=H�mcf,1aE%�Sc�}K����8�h؟q���#χN50w�&�p����j���5�M�fQ�^s�.��ߍ�3O˩�4�=o�
��(\�=Wv=4��4��4ү֨$�$}z����l�N�߫j[@3�Z��ׇi��Ă�ϐ�������f��N�0{a�:���G���Ğ��GK�y�0G�eLy����>��6�~��E�� 0|��T�2�,%xo���pNÅr�oY��8�ۈ�^хTw%/�c�B_#�y���cҟ��o�骎j�tw�s0=�c��*��^��~n�P�(�AkAmi���/�g�d��G^�읤t���)#cSޒ)�c�(���͹Ă_�Am��q �M�I�.p�0�_�䰒�_˱����qm�(��{1�%���(�\�xՋ��W|r*#p+Y�5]��x7S��Oz.i�p[^(��'*΄����X�Cr������">��02�2��0���{^�	ݟ�ʅ-���0���9?U�]K���V%�-�q`]]ԋ�5r��hH������I(�:�=NE�<��_@��8�up�|T�:���&u'������t�����J����+��q�N�i��|�<kq����'���h���3P�����)��T��iߪ9�ԏ��ve��ƂZ��̰S2�'5�ϼm��$���pk`K�����~c�D�������=Y�~l �_w�`�g�WD�3�R�Q`�c�DDjT�S33ˠ�FW3J�
���0'`VnzDW�Qme8�����S�����qy��E��o�O�>�d��D��ƹ�],���ͫK���C��6I����+�*0(:W[�FK*��K���΂�w֮��!��w<��ݾ�j�K5�#֔R�ͪ�h��5{���+J�`٠i���!���e���W�p���,V� ����z��k,S�c��lE5�ҏ������e���~B�2���0)�n�X�YѢ��������GݟV��Pi�w����⫯��L)�Y��2$ �bؐ�q�o��	'�yQ��*�d�8H��pP�M`�sU�{�u�oZ6���8�)=�@��G,����D��=~��zZح����~7˴Z�����rZ.���,4���j�ߧ��L��-��j�R�P��A������-|/���.�e\�@˥�Z�qf�����	e��ա�_'jU�Ta}��9{^'�P�=E�}�=Ӧq�F mi�M�%���=O>������jǁRH��OL1A}��6A.X:��l�C�Q �
>/����M����m��0�vujB�&�QJ�Xy�
d *��9�
l^&�����,�0 s�P�I`���T ��$���͡у�؁)�&��9}>���[�ڹa�;|��.�����7okc"��ez�)��Gn��'<؎����[Y˿Z�WFK5-�1�_}�'��2��v�I��7ClO�+�����Bp}oЀ5�^̚��문�JŒ gdY�վ��z�n3L�5�񑖣E!N����ohbb�V����h��y�7�U�HMkBzkA��$��e�9E�XRI�z���ݰT^a
-aBJ_��B.7��W����[-��{:.�	`_�ҕ#�O"~)IA�b� K�%Z��>��׳�4r5� ���J{!n�ێ	'��!���
�'�K�'l,cCYfT9�b��<���[��ex�)xg����@b|�3�k���ԇ^6e��C�������(LM�u�ǟ"3J.1�f�Oq�?�� �:
8�ìuY|��&�����d�@['��|]l#u��< 5��܄���B\�����6P�R�n��HrB	�dbF�]'($͇��d򤂢=�T�R>��#��ra�Tr��4);�4;!Y紫s.6#��m���9����TX���ʡ��L�r�T��_i�8霋��t��n�I�kU�ͬrF��S�m���v�:aGC<A�����э�1>1I��!�dҳ�s���`Җ��~��C��iPW�C吝w4HA8���i����ۜ}�*56������c��B�6(�?.�$Ӭ���C�3��T���c���x's��:E���*
0���2g˳��}�֚;���M[�֬��h�۝T{.���Ԫ(�J=D@�FICp��ǹ�t3��3�t[Sf�x;0����3B@��,+0�k���%�6��k��������_b�0�xmQ���>iߕ	�M����_��ܑ�ߎ��la�C�S��(FJu ���)�Bq~D�����(e�gr�r�蜾-v�w@�Qe[MW�A��1[y%e6@3e�T�?�����D�cYP�g��y���s2�5�F�|�����1��}Q����̡Uj�zi<��c0��-S�4Ɲ����Muۇ���ȥ����AŔ�ף�Ȃ��c}YZ$lY�JUVVJg�7:�]k���*}�(w��"l��IAj�P�o9��uP=��`�v��/�/w{��bcjv���S�O�NML ���L�8�9������}.��֩����'��1��#|��5u�o�z�1`�6%�z�Ժ��P�+��M�!�ō�x_g�:�,�2iL�y�;���F�14�ݒB-�������n�E "�:���Y�V��@ƠimȆz�%�@j�j�j���MR�C�ܫt�G��d:q:�D%�w{�V�P;C$PP�Ͽ�#d�2¨V�Z��ޔ��5���l����O+�^�)��[�ߵ�FĪ��&1���ۃ�&�$�I�Hm�F<�����Z}X�#w!�����+l*DF��z����C]������Flg��.�aS��a��Avx���a�G+��#
����g��[��/B�°E�c�YM�ayQ3���=|̒�b��j��sr�<7��Ih�t���I(��
�j��෯������Ɖ��([0��������R��ҵ͑4�k�,SA�mFj}��2�e��n���q?��j�/��w7�ۄ�|�G=^8�\|o���2�� ������qLs����\x�^N������L[<���l'���i�\�b��/ Z��	�iEa�G=ۺ����5�����C��x��3��ڦ����6��1�L����L������F��h���6�������l�,솰P��l:T��PJ���%k�h�����������\�s�`�cwf��m�� 
��u|l�[[�I����E{X��(��1�u�6%�,����KPҠ�^cJ���r���p?�v2��q��A�[
c�iԴ���1+.?������z�:���{ps�σR�@�>0'槾xN�ի��τQ�I-[�^9��x�#CFl��{�$*�?F��|`Հ����"���T�,��D��oA�q&���F�e���0D�3FS����>Q��bU�t��փV��TVq7/��F�� �4��T����x�Ə�O��f��e���Bc�].��dY����SP��$���܅B���@deң?(��3u���:v��ZZi�B�~�����P�_�^}��i�P�m�p�j��p��g�/h��S��Z�Q]s%��cC���
��,�y���Q9��+2%5p�b�͈����Yިy[׫Ԧ��Bq:�	��5����_�߭zS36�v��ӥE�V���m�t.�/"�}&��Yju�G����8V��ta�p���l��V��Z���b�r~�}���g��1Dv~S��a��0����׎��*`ܯ���s.�of���ׁ���u�c7�c�<k��W�D+�(=d�S��JC3/1be���H����q<g0����,u��^)}���/���3�ұR��V��ɉ��b���n@��=�v�Ʈڨ�Ŝk�:���UPb鷄�_�]:�Y𷗿"���-f`�:+9L!	�s~�4C���/7�m_o�6��0ܣ����xw}|�GS��t�1��쵬ꌭ,�e�����E�GC��F�j��9�sJ&{	���jH;�&G����?C�,A4��V�x��}�v�_4�amQ6@��y�hvx���z�41"lߴ�����V�&�Kb1�O�S����"�pK�qL����@��t6d��U@!�*�`⿙y>2��mU8��4�����[0�TT����}|�y���ŗdg���Ql���bV�h�?�Uc���j8[�9�0����[�gz�d�X�sf�b4`�e���FjO�1 ��<Ҵ�&W�9�V�#��Y	��0�SI�9���lp`8L1�q5l�o%��Sɟ(6^���f�z�y��|k9��`ڪ��һ�O�����m� ����E IX�F����c@�
���G�.�gA�վ�`�� 2�d٬��ͱ?��������㡲
݋um�fE�F�n��1�X�F�g��7%&˚�k�N<����[C�4NZ�V{ ���iHB��Jn!�� �6,�E=(�X���� .i΄5��O�?�m��^;L�į�@���g�|KT��c�"��r&y���j��
^���n;�g�͚U��?�s��yuZ*}7+�&'gh��Eo�O�b�,�I��qG���#V~x�{xec�b���N�Y��N���.G4v }-6}dô�EJ��/�6�si��3��Ϻ�\�kz����;j N�Ysh!��������ݵ�����àDYb�����5�R�WQΛ7�{m�V���=���xe��n.��≰�I��W`Zb������>�ue�0����t����T�1LU"5���؞M�B���#9��E=�v�K��"�d���Ɋ>�rӐA�����aR�&�<��u���m7�&$i�(h!��QK�c�*�ML�q��Ʈit��A�*?;WhV�:8�y�9�A�n�E�0B+� ���2��I+e���Ʈ�%MT�g�	0-ǜ����O���E�me�_�D��68�8+3�lS�Ϣ�)CI�H	NAB�S���v� $Z�!�Xeq_�hAӥ!�*\����F����������0��i���795/h���i]n�n$�w�|QY�!��S%�K���)�XLdn���
���/>�-����ȏs�2��Ⱥ�Ґ�ջ���m/�~R���Y��_\�=�*�NWeIJh��4�������A�$�b8���c�+��+b
��K���g҆=0*�v��o�O�r�[E��S�~�$���b)dD�����C(���=�Aoh���{���뗵4J?��\5L�_��?DŶ��u���9�ܖk4��x3��X��r~+����;!M'1����vB�V��m�~������_��tK�����_��/���s	$��ɗ�Ϗ�W��d�
#D�'C֚���J�z��'Z+		\:�j���q4>#�[��=Y��^��_Z�,&k@�u�$w=�����g���ZL�o�nc�$&��>��DA�cd�绋�.�$T_Nhh�R�E��¯b�3J=�gؓ�q���{����SVk����="��)oа�px�_��.���*�`5��m�?OW��"�^��xu��>}����d=�4(�����+�˽������v�D]R��_�nc9C�{+�n��aH��܉�>q�J���F��/����nFWGS��Zihl"���:#-�I"�,��{�ΤU�:'KT��n�2z3� ��o*�$;m�z��Rwx]�*>�Q)���A����(']A=}8}\ٹ�:��)�J=�m��4�y���\:u.dˬш�e��/����f�.&�u`,V�1��r�`k�U��D��t��5y��\@_���oqn}�w/yi���N��2M��V���d�w�)^R޶�]��Y�a�-��=U!?������
���B�u�F�&�C��1�PʺjU��
6��
�Z�H|���P,����?y��3�����,��8���%��j��މ�=9��g�4�\�5��J����Љ���쥤�2 ����5�<Of��Uh�Iw�.�Y��^~���	8��ߔ�||�v�׼ K��I��Q�e} ��B����8q@+!�*v�_5;��2�!��#k�"Κ�� �eJ�ܹ#-�~�(ۼNE���#�d%�R(�b��� ��(b���V����������:C���}��[�7�ħ����7=ez�on
�<*�(o�g��#E�i�V]N�:���T6�x�ꞇ-� ���-��\�`��*���2^0�sB�4e�
�QTW�^�i5�	9.�b�����t��f`b5Ope�
�!�d��4l��$�� �^���X�l[C�6��%���[3g�gⰖB�,��өµ�ELE}�/p��E2	������v;Qk��\���<~�&AD�����Ώ121�+��4?��\�s-]r'(���a ������TR�8D����P�F:����[���"O=��15��:A���A�ߝ;�ۘ��Y}9�ۣ�̶w�;���x�ϰ*ѨS,(W@c�K�`�����/4J�[G���	�7�	��}���M���6��IVF΢����Q�wf��u��0Ō���[��y�/��5�>�gj�&�t�Ѥ�^h�3SQ&�,֣vs�*%�2�$$U�|0�;�Z=	���hR���4���͇F	�T&^kW���r����/���'�V)/�><�����ڰ�-^���4D"�*o�9#/��yE�
2L�Rb�����DÄ��!��&��C���6�=�|_��x����|�%)X'�5[���c�͈�=�C���B��+sE�O֋7>b��f��p.ڽ��f�4�}=�W;A1l���mCBZ/xԈ�ҍ�h�����9�.�~�)�魠���|�PJ	b4Sk����Y�]/>k������K�(05[�oQY��u���B�5�@t�=h��*Ě[e�*�[_>�����j�w��b�$�<�E��
-}�z�ѽ辡���e����h�#����?�B۟E��]��*h�)ڤ�t����w>14}��f_ȺJ>,(�Me�f��L�V���+�O\��y^,�v޾d\�; �͉�����k�I��l@lFAZO4�ߴ�������ڨ�l�_Z�w���'���r�A�5MX�6#e�ش��B�n|���cR��� �pɲ�ħ+8�Ȉ��E��B��1m�o��f��Ƭ �cj�s�x�z�"�~���&���i���b��jN;LjJ~�3�u*�fp西o�C�1��m�Jo����WGeRk�T���ie>$hD���_"҉��s=��������TM鼰2�WwZ����)��2�*��V���v�&�]��a���ߧ���b<����7L�ͬ�K���U��ϴ@�^�ƒh6N%�k`���@�r��1f��*�I�Gg�6���t���}|�<d��t/�R�y͞�U���y��P2t}� u���|������غ�Ӊ����L�$�����Ȫ�='jn
���D�@Ӛ���-&��8PU+�OS�>X�Z�"��������:jE���Å\�s����^�En(����M@ NO#��	�Eb�\|�c9S��M�跏�s&�:��K���<���\Erđ=���^yh�2H����wx��E�������@ev���U��9J��RY��ď߶�P�i��zP�B���ԣ6�Ujh���p������g�{nW�'=�Cj]���Niۤ�db���	��c]�_�N��=~�Z�_C��7�����~�Qlu=z��'����ǰ[B�ud�c���"�X/6�+R�]��m�S̝�m��L��"��7���X��H����w�msN�tD?g[�9e_�J/�bW�Y�*��A��8�x���!'���g"�Y��8�@Ե��_�S���rRFIo�A3�k��k+�Дح��KdMOi��n����c�P�V��L��;�p~�q�G�m^T���|�b��I7���ȴ\�߃qlX�)k�kʪz�X��L-{�{�����;/p�<�$�@	��:� <�l�v:�B��?_���z��o�A`�X�$���>Z;·�)�B�bw
�n��^��e?��JF�.Uʟ	���Á�WߣH�".ިe��=��B��)}R#�Ѫ]x)�K%/�*�f�D�jP��jgW�G�-��
�,�	s��Q齝�n/sM�^a��T#`lJ�����f������B��F���w�l6� dL�v=aS�������\�p@�=Q�Q��_���~t�(L��SE�����ǰ�w4�<ųK�w�`�l[�G��$�f�������f뛴���KgR����gd :�;��&f��n��p��C��b6O(-�����<m�0��T�>��Pb����jRO�����#G��´�2�[X��\��.��賂{۔����S;�]zXPn�� t�s�������O+�I�˂9L��7��B<0{�)^��Jë/�Q�:�4��ܴ�܇{���I�p�*�2�l:�=�,��bu-`eVw�+�kT�:�I���������`�c���8^S��B�����'��ۓ" H�G
�"t4��];HM�+�8�������l�pn��N��Q������J��t�"�x�;QŖG�;����h�XN�Pm��NGS���Z�tȮ!���o6��N++ ',2f������\ى�"T,Ƌ��+���V��-�v.��AJ�;>���7K1=,�w~
�^!_�m���W�����93�	蓥K�����k͟��e.�Y���i�띁�4r�4B�o�R�m��}�9�i�G!h�������Ψ�Յи�B��#;�)�$EZ#�+��L�i�i\B�Cj��pXS�q.j�t&y㒀u ���l���H(G��zl%�Hp~j�oe�� q�2z�AB�L��Uw�\��lcKھ~H0�
������w޶�ok�6$��O�S��&�O7�����Fl�z��4LǷADX��P��Y�.�)�΂�u����&�!릩���d�� ���G�ݍ���a�R��\���Tu���L��e�ez��:��J�]{������[�2��������Sj$qu�zu�J���Z��k�%CP4��Z��F�f"��FE5�]�y`�q#^%������K���,O��O&���{�p�fP�u�ux)��tG�K�MO��=$�5��8�"}�3��������:�ʙ-�#�L��I_J��̧:�U�$\f�H�|V>�S_�~G����4̳;��7�(�!˸�lI����e���Hg�����O@kE7r���м#l�/���X�l����e1pen[J-`� .3S6"Ȏ��9LI!"]ar�G #���R���pI�t>�{*!B#k��Χ�5Ҿ��x�1UD�}��e�a�%�����8��Ɲ$蘆��JD�y���S��M�n�I�o'ʙyK�i�@-l�u�Dh��1���
���h	jq��ģ�J�V������ϻ����b�k���]�¬P�.��ȅ�_"*�L��쨘ІO%�K��ثi�q?C�:����pl5/�<�I��^hJQ�7��UZ�����g��֐��h-�K�b���Ɍ�
6</_�'��G� ���s�VQ4�#'0^���@[��{�<t�%y̢mq�4+Gs?��%%$���\��g�QAjJ�8x�jb1�M��j�B&�{s@8���������A��S��o-:����_����{������#'28V������B'1 s8.R�H:��1�7�P�u�^�5C56[3���u�3:L޲��a�e�S��7�JZ#�W��e��'Yi�a�D9��{i��=��]mN)#�."�f�ni�Cp �O�
�Hj�-�=)98=����7�`��Kh��34��|��>{Ғ5D_۹�,�Dp��^e�g|~����w��-/a� KwrIC�i��Z� �0��C�S�[��n(_ꜛ<|��S�)*��b*o��hϞjP��}�a�X&1Zy���Ttl�|�KJ��id^:���QnK ��=Bs����>'E	��������IZFIS���v��I� �� �= D�ॣ`�ÙX��]�@ ��ϭ�c��<�2��c�M>5Q�năg/��(O񋂘f_���{���roUt��V�2O��O�^>\�3�^]Z+�{�I��%K�+5�Ix{���k�^��C�����F�e6q�UF��G�\B1�x���)��P��|p��7أ?��bH疧N�r����Y�@ȵf������&�t5����7m�r}>� �f$�c��I���_�J�b���2�� �6qS��GqB�e��J�r�	&���ǐ7�_��e!&z�ɉ����Y�Nߛ3��@�h�5�z���UŁ�Y����Mh�k��y�
OzP��T��0Lv����<��*<s�D�����o��2b�Nvj(b�Q����W��o�߸��1�\V�� �8U�P��F�����n�Kq;F��H�x:��krX�.aQu&��fZٽ@*R�%	�]X���N��-(��K�pP?��rгΥ���ֿ�ǚ>�yl�vW��{��(�)���t��}�y�a}u����Z����X�l������m�1��J`�����a�����0Wb�L��������2��{g �I92�B����:}s�Vu���O ��8�D&wi�*F]�����)y����R��.O�4Fn�9s�Z�Y����H~n��ؖٜ1�ުbs&H�,8���ڦ9B] ��^" ܐ����F<��\"�VGZ_�NA�7�˷+��ψ$r����kBڵ�/�D��^�gh��&#R-˜w����k��?"S�VQp�F����U�uPQ����B?ohA���\���RI�d�7r_����$bZ���u�rC�j���6�wD��O;V"�I8q�������g�E~;\ɳv ;�
����@ +���k\j���%����Bߎ��M�p�P�soɻ_/b��U�U�"�|����S�z#eI���p��hў�N��:�wd�f�
��x�S�T��0汫;�{�ӹ(g�'���lӅ�5K��?��OST��T��0L��Y-���IeP�ʮ
�+�]9�tj,�ub��0��!h�����:0��^R9�Q��o�� �b3��؝Ï�6&6���l���]�rg���o�0ty�?(��5�M5[���9(˵h�g:��B����v��Cy���3��G�YRY.Mwe#�y�RJ��߷�̄p�4-�-�+�G-B�aC�X�V�f-�H�ȨPi
:������QR��Z�d�V�	�+�?�v�������U4��~�N�M���Т��v���q���T�]�����.U�F���oA��l-�1�S��~r���(_����)0�\�'��b��?�!c��	��&!���]�s3�pQ\	!`�U]�%�z���\*�dԟ���i���t��Fu��;L�2�/z�)2B�(K�֕&�9�H���e&W&�%D3Ew�P��\^%S��Kg�;��,*\��ħU<]B�.�?�B�|"f�
i=+��oի0�'2}��\�i@��l�j@zn1�?%��\T�P*X�W"7��C���y�q��t�xqY�Vnf8<U	�4��$������|�rS��μ$>}&���19�A�iê��Mɖ�_em�z$�8�p­_tLםg��[�:ɧ���������YQ�>�W%P�`W�@*�w����M-J�j���V���(@��e�y�e*6��d��d�9��������Q9�ϕU��A��X��T��%�3���;*�!$���~�ς^2�K��Q��0�2�եד>������A�Uňr����2�T{ێ+���L7�H"7y��j�#/��I��1S�w��@�s��j�L��R�>��A����D,lQ��R���������t�~����`ڭ��;�]��@<���Db�i����;tݟ(֝��=~*@�o���h��ߞӿKY"�P��uJKZ��Ҳ�}J�\V�S"\=���o��Zxg�!���C�n�Y� ���:���v�C��(~��q�:����1=qxN�"hV�,MU�/���XR)�lg�:֭sI$�aی�'?��
��nG\#��
���@,���;�j��:��·��$4�_w	�MlG�Tn����QG�9��J��������X  |�w�wRN>��1�Q`1o��.�9�|�l����)P��5z�9ha��Y;��%�nť��-3!A֠�ޱ?����)En�����?k@�1�l���/A�C�s��_�u,�bQ}i⋷�3���E-�w�K�˖�h
/����F�Z r��"�1AqLJFg�%�B}��h�|�M�z$t8lE���`����i
�P6T#�	���'�?k�v	�
T��XY�'�_A'E��پ�����?^�X�ç�*:����tr���u�07i�sR�K�xܓ{
�ڂ����S���U���]H�[<ii�������@� P{�hZ!'�1�EW.�p�j=59��8�4=h!�S���]^Y-,hSh�S|�XL��	�*�6?s�e��.�Ѷ��M�U�!�(��ߑM�NI�'��T��璦�&�Aw��,w3S�'�oJa�P@q�8ɼ��L��?G���im�xd`|�kFV�DLs�\�p����7OLoU�����`�6�M�΂T��2�";e*��k�b�tBMg$x� ����)�1͉�@���y	��6ߢw�8dѹ@�pk��k�W$���״��(�G�6��->�+?K�R�K�4�a�y bF���K�+��L%���*����n�{
���(�~<s�p��4�J�7�է{DF|�xo���I5�҂G���x��A�|��~F�:rD�36�dJg��A�^�o�#��Idsc�T�&Oa�@��u�ٰ{��,:AR����������=�̫���)�;�D<2�B�g G�-�v�S�Mh���`����Nx��r��K`J���-N/��� ,"d�����%���!r�4��<��x8xWE@͜��&O����TAF��ЕL'�~�Ul������E����
�|wwJ��kz�X�٩b<����L8�-�[;Z����_�w����Ė�$���ÒP)��
�7m�A�Y��B@X�:Ww�DI],
�h{ry>wCA�e\nb6/L:�Q���p3-@W�{cx9���^)1$7��s�n��8�����y�G؎�[ƞ�}!�D�l��^����Z;��ya��GlܔО�H��փ����{�0�u��l��_W����S� �8����=!�⛈|�j�j8�do[����-��G�ڳCW�_O�a2���a;�br���