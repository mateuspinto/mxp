`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3664)
`protect data_block
0USWSUGxovGsyBJteYpEoVP8Rz4ZyQkaY2NB9Glv9ZMbuBy2chIpek8TrEfZ5nq7kcCL4rG9hRUG
Ax+FsQ2l5lHLPNvvR/g4jS7Osed5Xz3XVR1HS6jglA4dNKNFB5QO5J00bjrBYO2pr/mkKSqFcvgG
cMihIGE0H5eHcd1hh9jW8mZYngzKWL3N1JslrpzysCQMeAa5C369p/Rg+LnKhQgL7cJJC/DulAb5
9cKH0oMENBCeld6C8Gl/oUTAafXZyf7nTAHPVnU3x/4vg6ggthJjQ1jDuCwh0vqgt5ZFPrw0KeCE
VNKaKOr5POg0biTckENI+RZCA4yxZvwBRXtXaKMzh3fYrD7W5PwdGMVvkbA64Gp25puKajE2o/PV
7tGNbGAkSb+sPLL0ywF6ZBNvw5lGeIYroxhjkw1G4YWXU0FYgO200Ln2SyBSCsxKkOrz5afcEQWY
3CZZD1m1LpXaPeWYM5Q1MFT1XNr+XcbAbWxk519Q4C9AoFshBBZdjS91i+Benax6S+biguCIWOpw
mJ5KGNam3saG6TSW0r+BN0P0fdjh8xVreavgGtWG9I/O4ghFE/fTChKfiP6hPlIc5u4kW2FtVmaE
upsIZdc9l7tR1AViMMrX77Z4Wd1UT7ePvOdG3ImvSE5+/Qh5u+sSgu4s7hM5AzvBbE9oFvoOEGSZ
dYtrtyYNTOvTatRLMVIkorgvUB+o/RWGVYkIokGVfrKaMB5Be9eP7glVpv2pIIa8mW4YiN1oRrXE
XI2MnXZxQJmkxQZvTVOXX1XA2PVTeGF3aS6oXwuUTYP7IsrOysv2+cj3gLAADIjcdNP8K20mG1mK
G1q7M9jG0jHlY4PJQ0kYtYrJDv2JAnumyVewp1grpPdgIh6CMXC6kvQ/0bhGI6+zMtss93/AMvLI
iZSML8/wH+/gMjB3AqR6MeoObsWMa5L0XrhfnZM0uMGpbSSgznoq3dzKrhVISwh00BtBb1FAJI4Y
M001T/NKzYyXCR98Ig0bKK60psIwXmkK/2ClJLcE7eCJFp0GM/GEJ1e3qeFF2wfsKjxfn4r5LU6w
eie38a/9ucByUMx4mEQM0mII+cFl8meMhaxrOaqIyowlmd7B6M96G6J3VfF1ubLPM4jG/ADrlvph
6zRZDOeYO0Lme1Wehp2r4+m516S/tWCwUc9tIHOXJa1sJp+a7xq1UygipE9jPqGx+JX1OnoDwVlf
HA9VvHE3malAJ6ZWTdE9hLo1CIKmEDeonD6ZP2YR7EzAVC0u2JBRBp9BW7odKQh4M/+1dJHqlUtP
tL1vG9YtGnPKSWI/wS+a2euvZM5JWwOVKr967orCyOFpY/YobVDIkrUnBJI5jLCaa0K4Z/qWqeSn
4uL6bfh6PwOwPzAs+LtN1GSJcenZG7nGivR+TT2CXjIginOQPDpPuU/5CIZCprsIVFov6e0PjA37
AFbl211zmgOJE9MX2V3nvG3qE4cwwl7lEhP/SwsGIGiYtev2lYh+QzbE4GuHFaix9XfkmVuB73HY
BSWHVaK/TtEM6tCUwQanzG+HkENVlRoU3JMIuYHoB7ITvHJemPgDqWIsPtWpZM9fL76lqMS+7Jnw
mJQ/i9aHUG2MAHc7tci9aS8EX/ymAkGlDmo+G5CW76zeqB+mcKG80Bq+TGA/lMxo1ZxX+NPm9LmG
cpfreqcwMwhlVrFtItpIH6GAUxlkWCjgTFtTdO2KuGI7yEXwd/WTqvywg/bJoeQTyOQrP3UICIk/
RIRNuoRs0bD21vrmLnmVdSk2PhLCTdhPCrgzDMsDdIzcJ3XoB3F9FRMqTyZkLy3Ob9G/VE4C7KSO
bDTNbMTmjMJEXLJAlSfuVmsAr2E1I5YdDFQyT86ronQfTcfpGhuXzwE3Ok0Tw13S7jOzL7NR6FzN
n3Qq1BCNVpSJOBpPpF+j2wkrP/iRNMz8/d9LD/9MKgTT/EJjKYyqUphV/hmC9yfhzDEQNc+aQeVI
yu/uO69vzgRyMI900/xZ4Hnp6yZgB8+fBNVtQea7qQnqcHRPJ1fWsJ8RE/ICHCeeK6TAnqQY2DOO
GsGg4WylmwcLlwaRm1vv/u/vYasJSUvgs3Uu8+r8Jqug80EkQCvBuFhBU0KEwIPoUoHej6x8AvAQ
sIyxjoZxekfog/Gb/h7oZ/N+BXwr5rfWlGVteR8SAGJ3Kma2wKx9jMADJbKPhdeQmLLrubiKOIT7
UGTdF9UP8JHCmxVGx40xoSm8AzR8r2fxJpa4ZVUM7UD2+Zlt9dYxrDHf4dh/FEzqD3KE+GFZBxxO
uaFLKz4shBZ25qsMVir4mcXAUgLYhoalrlr3B70q8f3D+pqnLhbdPZ1lwmXoVFC8UmB3lqysri0J
9HzzMk389JPMIeSxoLclgEW9/luw8CHw7WiNEMAlftN4BzEmOi7JGv7ZR0xtEc2QE4StedBZOd/x
Mk+zyB2vH1ntGXdM0a7XxYVibavh8z2vj3vRP4DxqUfXqb4RLFpoz0tyDiaJYAJ389S6R0FaUNhU
HLGdmE/s3CQUc8jGiudNI3ebu+/uB/LizYdvIx0BHKKIvJ9Hv0cGnskEYLBZXXvBbV1JsDtUXHc2
GrURluZIGux5e6btxp53ZTlVrjxu9fnr+yVyU67ilz9jEwq1RnjqR5sD4wjEoLQVqf4UZBWsFchI
vmcKT9VKbmFYhQyNF64C6TtLyehwEEAThQy448RxqVJog0d0nR7racL2hBU9wfKjg+rN1MHhvtRO
f3u5qF2Tn8xnYfDPQsfDOzgwZBwXUUNOYUGQetaH4WJNELZmdKxrDY3XWVhSh+GVA/OXOdCYXCBD
dYsgVpt+qnIg/D1QcLKSG1hbB+bIS1ef6DQX097qrSFgB6SiQcaMUYMkS1VqD1utjq9OfP1gEywG
zONcUN2M1H4DTBinrTWGY3JsZ5pYy7MdF7Y+X91tO2XDCmOEnobYuOkfHHBVRshz19WWKpKxpr+u
aicQwL6rkgPTd39UIavUzlCvZJWqwbk6FkpSFg7jA3QmaqY5+dPAynUa8/0s8a+pxE9v/1Kz8fNI
dSV6lq4b5PUDJcGM5qzvg6MnoZS6EeZ6TRz+R08WTRBrcmPjgmyO68ntCofkw0M8C9LbaI2pSylI
3RTxauT2pb2BsuHDKwbPsQBpwYTcs2kElLjRb+WtB3eVobBcJCBl5ucePEIJP1eQlsYi9MjEyUZA
jpR/7mJ9GpdxratsraTlr8SGKjHm6ax+VsjZuuN1qpeKEQ9qwaVvTj7Ps3MLyvIPmi8qmjawH6pi
VTYXRlMrWRSxN/wAAu7VhW7Zmno9y7/Umilz8+fHQ0c8BWxvmucuCPIOjKM03dCsvUiWSVqQKTnQ
a5GpMCCLVK+PvLJCLSxZeU+LrHMIDqZ3FXjMSW/zm2EV/LHCV148oJxT+rm3yL50sTt1JE7Khfiy
dWt8F9SFfjeS/2ojSpk3d5YEYi79WZ4MYuHiHHr14+oa1MXSpxyL0ycKKRmmNogrc0MZ29kONif/
MIUpsIWnzjD10/8vVVRUkgKESVU7EqBVr5Oac+KlF20q8F5Yy1Cw5t6BQ9TZ9cvl08kdCa4I/02p
x1Ud4KIoN6vm1tTpucQ0+FwD5HIjNPjpShdZGvZtJSy0AhZPWAjU7WLYnt0ZpFupRF6BUxCion9X
HK8TBijz+2Wk4xX/97DcCTXrCPWRB1TWLB0Xz1552p+aBw06kwiVm+4at6qIY8ULl6MolazX7pWw
wksmn9kwyEv0qEvc8tS3A8Q16z2ADCrdT22jf4J/t0s1YS90hEWZKRZjajFBRrzy6RKuR5galqmm
txUac/7IhlreA1egF0JF6d3cMcPDPvYzl2xkJZIknvoxqT4oXBB9+1vhMTNCJgMl6J60yGhaoKCY
0uOkFoOj8BQz4lr9TadObRNXnOdxvroFikYwVbbbghgF/E0APswB4VQmCOGHmBEN1tGRcfj5V4WZ
WS+645obIyEf1zAKVqWIcubP/HadNu3YG7xHgW9fnGLcwRoQ2vfIjyXpRBfmulB0dXAxMUHGHd/1
eBGeE0acbmvcZOk0PNwxdHxY6QIwylq8QoHCQd141YGnTcIFonegCCdx41oIhmn0FpxXAxZsUOgX
7qmKUnVx+VOFjNC1JW62v8ncG/GAmPVRvzjKolEMV4KjcLdaQFBPW2GR4YJOAL3WIHWPQYjHQonw
NEW+Kx7/S/9UcEAzYeq8nDfrFg/YqehPnpndb0ovqhu/1IX9+DVnfj8axI7dZLclD/GFhgu6jzXU
Rv14eNVhpKNZoP4TnYWLn2U1bB84ooGLlj8emFZq2GutJuX8bNPGz7Vl05XyjfJHvM+7+Ty/s/dR
LEOqNAkpkNY+GR7r+LxUQ3d7YoLfrwSa9No3+byNG9uCZ3XUYmpPWwmLAX65pBP3lbNytgWsOmXS
MgyXE3iy7HaUft49Mwihk+yfb7hNIXGVPvGulXcz4JVnWKmKQrxwTprKNfiqPpbvdhSS93PKo0ji
GdBJIZF/941ojEgMyvKkdCq6tPBgZmJiZwAlwIV2xNiDtwwCLc2Ki8bAvm/YAeY3Jv80aBC1KQX2
nbvaD9Lwt/e5P9VAs8bEv9ffwxUsDR4LFZEHmST1EmgUo7zKSk2S3ddh+XFQHe+tKjZNRLD8maqi
joNFPM4WPSegrt4aSvUb20e4Bc82NknoWq3HkN0JNJix+05P8TOldftLEtjnZvAFOuBdPfBgMSXk
hAojp/T/zkwjbnPSVxqVZ7IeniDAzlJ7JK1V33ABF3NBva005QvOvg8oP7/DPDJVi1Jc1m5632UO
W8oNYx8Itc9qHpapFShdbJGLxBEahOXPCN4nH4YP0i5jyTc4keWnUhkytx+lfmhdw810obxVk6fm
BoaXCaaFKeEY5xi0vXGcEg==
`protect end_protected
