XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���g�FN���o�g�����"j������f0��r78\�>e���9d�[$�����T+�
F99ފ�Ve�w��4xPв�-D�)Ģg-\���������L]�<p�b�?t�7�Z�����0�k��u����8%f���?iJ�^+v�e}����k�[���(f.:^=���t-	��'��D���\����kt�w��!} �v`I=��]�R�~�u"܀���������'՜Uh7%�ʳe�Ow',,QM�XJ�@��A����-%: !&��A\\
���&�&�����'����%�*���[D�]��;t�!>,n-I�[@���$���i�]˻��d?E^��ڡ����V�7q����̰O,�R���0�/t�$c�������1���vU�*�����#"(�0�b��v"$^C�a���H��������Ʃp��m�0G��/.G�l\�NHq|
\��B)�V�:ðz.�I�ՇN�F�&t�^7�n�e�,�v҆$U�Đ�-�qt��|�#���YD��N�����u�v�f��6J���1"LK��ES��숭M������7�+��Ei�ud%�M..���q�X��v&~�w6�?d�Q��L؊��m��ڧ`��k���JUaӚW��P�kn2����rϬX�D��n�vw�K��@�c�ˡ%"���Co��\g������!gnSp���M:�䅓H ;�  ����BdhJX�W$m��،Y<�8^��޽e$�W:<�JmXlxVHYEB     400     1e0c �,�@:�;�.��H�Y�w5����>� ��0*/���x�u27��5)�*U�� R�f����u�x�n�JSl2 _� ��k�d0^m���B��|Xϙ�H�̹z�%Iz�K���w��-����J����!�}j�`Ä��4�r�:���Z^[�%>��f�G��|j^�|�����Q�x
8�7�&�=�gg
.LP`����j��ww8_�m�2T�hѩc�A�'��I2]�P�r�SMp�7�����t1P1}v���'C\6E��TѺ	��0:g:��li�"�yn:[]��Jv]�#bb��+Q��$^}���`��Y*'���Opt9����8d�X_�ϫ%��1H]��Ѫ���K�A�r8 e�>v������8��f�\ ۤl��-ۛ��~�@s[��\���A/��d�;�"\��#A7d�a2���X�!a�	<�C��ޣq�}������/��Y�wpj�6�d?���XlxVHYEB     400     130�Rsk�}�{֥j\��K�@~��Xv�&�r#�zv������N�����^k��Є�Ltq�� ���IW �k����/��|���]�;�s�����CJɤ�R�A}�M���R �5�q�.����gq	X��LU�I�K����ҩE+�8(C��=��ji9�A�hp�����MŃ���������$������t��C����;Q�tЍs���>��	�(��v����列�J�w��q��A7.�k�۴�ec��iэ9����?�$�{�1JO5�QB�%��`�׊��R��#ihXlxVHYEB     400      e0�� .�0l�t��e׺]v�'�!,��dZ��N �|�&�%d�¦���Nd�3�]~��O$4]0��)v>�!����ޚ��H)�<�J�!��P� �&؇f0�(�:��$�աp�_�X���Q�I&�8"ρG}���z�塚��/'�&C�軸��q�S�Q�Ic�q^R�[��h��!Xʒ��-o�G�� !F�S�K������B,춐@�FG+XlxVHYEB     400      e0�l^��v��J�%1\��$OG	:h6�>.��@hqI
5��R�������z2��K��^�?�:�P��=��+Cǲ����h�|f��W�,=퍯�f���x���G�EL���^5u��#/�q�4����'(�d��_QVz	����F����X
��K���PLWԳ�k��P�ݣ�&d%*n!�䌄��$<#O�bt���,	�z9S?�U�4��?�Ѥ�@��ދ~��o]XlxVHYEB     400      e0�F�@�'J�4�d��w������Lҵp���_Cl��V��#�[/��~��	o��T�����+�{�X�g?���ċ�e$��V�5oh�4nG,�b���e��mX���âb���e�ui���Ww�]Ne�5��-~��닝��O�����D���
t�Y��x�ԧ&�U6�yIh�0���I w���⾾,�!�y�v~���[�
C�E���XlxVHYEB     400      e0	)�bʼQ�ny�x�? s�BQ���	l��<�(��5��$�t4��sZ�rه?%'׋�D'�U������7"akY����t��� 8a�K $,�����j<St��8�d�`�`�!"_�#�8|{����^h\�!�Z�qm�~}�@��:��� }�Ţ�=�H�o��w\:�!���M��$e��Wu�Lٖ���������ύ�E���(vE�Q�XlxVHYEB     400      e0aQ1K���0&�ұ �>-�9do�{���1�ȿ�nL*�}��׬�t�i ���![�D�aT�=�����n*��M���D��2p=J���O}�)ֻ��<q�݇iKR �k k9�?�f���Bɱ�b[Et�:�$4�5�rr�l>nm&f�<��,���ky�>Y�W\��«�{߫|>ˮj�K�H�6����7��eL�����q�} n��ҧ���XlxVHYEB     400      e0�"�����������l��~�������	�)�(�A"�*\�D(���T,\�np�7�I�^# ��c�./��c+c��Z!�@b����-�n4��������m�k�x)56Y��Bd�C�#�B>�L����\R���b�<>$yN�����Fm&"C{��0#{�E�n�������X�>����";�+�����<A&�/[yq�p�K�S���4k�]�8��XlxVHYEB     400     1a0Z�/��u�,V�d\�����	��,��M�:����g��Ն�.���O�^�25dc27hF5�Oő8j�j�$?~�2��ĥ��v�һK�������ہ�}��Ȑ��]�X�9�'�u���z��EI�ݡý����w嗵i?�}:_��X�Ҙ�~��Qನ u��n�E�H�*ݬ6��I3i�k���#��Ľน&;���o�����dE�=�V�t�Pd4x�f�Ȗ�We�;Z!LR�_q+��;��VŁD���<���DuP�̷wϟK�Ys��p��ddJ���>hK�?"|���)	Y�8gΦpec���70l�1�Q`�(�ĖS�����ni�{?�ؙdi;�v8DK��~�ݨ�w�h� ]��$e��Ĕ`��!iNr��g�XlxVHYEB     400     110��	�L1��E�I��7g�R��gts:m�Շ�1��yԭ���y'�
Ϫ�z��̅iG�r�no3H]���%.e6L�U����� 1��������ޣ�]1�J�ے�
uU�`���p�ϸHo�'Af���)[$?X��5U�FFftf�(/FE�+��-���΋|K���ex��KJ�h�J��{�6I��-�R�[;ug�e���z���qL�feL��#����fVI ��Ȓ������#�;�$e��ɬ,[��!�J����0�XlxVHYEB     400     180ov��:{��1wX�a�ܯ.>�-�k�-���<��s�Q$t��W{,����^�b;ߘ���}u����J�����.�"mC�w�\��<;gA�Bֻ��
��q���8��c��wX7L��E��Z���&w7���ik�Zr[n��կA��(u�F�#j���8,��?��E��EJAԸl�?�K��f�RN�9��ګT���	���)3}��g�5-1��ޭ|�+N��4�U7��K/�m\����}�. )��m��x'�޽^�x��K]��ゆ�_��ǲ�s���S�Uu�Ҷ9��lp�c�@=#�������vT�$Td;S�}�h�}�c��?�loNv>�/�Eo�|n�u�p's��D+�b��_sY���XlxVHYEB     400     120�f<;|�{�#$�э�yef��uRUt�)�� �9'�n�ߎ��׺�Mr�> l��ͳ|��(Y|�8�J�q�Xy+�˽g6du�_���NN��b��������Ut��G��+�[��C�ܜ��l�/\��ox�N��(��~t�R���BD��w�F�\F0��l�|��y��1�<�~F�}�^
��̑���`
ƞѫAܼ����Ƞ����rJS!���S$���Sԇ}��Af7R�:�RvZW�Ԛ]���A����W�]@t��ǰ���J��eXlxVHYEB     400     130f��?ҥk�Y���g+��_W��փ�!�6^E,8@>�@a��S� ���>H�|�)?H�@evV���j�KEz�i�
{�>��r�c���e�cÝo+&��l��h���L��t�V�$��eݨ��abr��-���xLR	qGJ�h��}��@�7
��H,X��B� �� ��W��f��ӱyM#P���(#H�2�d�	j�<�����
�J�7���w��=	�kLc�VF5ق�����q���<�2���Q�N��_��`q�d�Y+����[���e�c9iӕxXlxVHYEB     400     120�0>�=��/��f7L�:;��7	Ӳ���&G���濎/p%}P���uׅY5ZC�bYe����9*�<�g�j:vE8�G�*_�`I� u �9#LGh�޵��]I_*A})p��)�h �4�gV��z)͑�OaөL���^��p�s��+��k����
~���m�	������}㮸-��uE`7��� ����F΢�:��-r�lk���5=9��oF"=��C��$�4�l�f��X5вj�%t�?�M6'��4�[e��r*{M/�XlxVHYEB     400     140�۠:������z�=�@2n��䢥C��B�)���p?{h�6UT4�K})�Jlm�삿?��A
��H�hk��H�{�V���A�O��g9�+�,�{�"Ʊ���G�N<W�6)��6`��Ա7f*j��5�=Q���Ȳ�/h��}޲H�䳃_��VE�<��0-�L 6�'�Gb߇B��:��#\�|>�����&D�>z4@c~��E�>�^)�#�)�pZ��Hh�1�Yǥ��`��Le�\Ŷ��3V�~s��6����	W3ε1b��[C�W��d
���?�2��x��<X�׸�O|��8\XlxVHYEB     400     140#�pԒU�͕8k�xv������m�9e�?�T� D���	�`a�����=ʡ���t'��K�?��\��]����V��FV*J艣�O��e�@�1��K_�!�&�L<�=Fql[\���+T�[t`#�!\�N�7E
4�x;�g�h)�|	�u�X�f���v群�E~��pM�l�2:/���6_:��$S0�J�,�ڹ��̵�i��J�Z�Ip�S«PT$���U�z5��ρ�E��;Ӷp�Bh�c���d*R[����;�0��)�=w����\�p�@�Y�mj��@���]�
qr�?�'�A����&Z�^�XlxVHYEB     400     120B���fIc E�$dcB�ґ VX����_:�ݓS�g��)h4ڣ�lNE ���}3[N|�y�|pa�kT�a����[�Ji�l�K���H���y�*���������
D����4�Ǥk��4HoMָ�
�&�y����=�AC�3e�_��eu�ݦ,Hqˍ�>���B�4C(d�m��u;�9s��=���M�}H�ܨ�D��#c���P93R_R�k��7 �֔VV���3�Nh,�(`f9����������2���E@��6���=�;�6;�,h�w��XlxVHYEB     400     140�@*b�Mh�[�,���9-��\
/C6Am؜�d��[� ���0)�������L��1g���ふ(������R�ؼ���0T�e�� C:���������+5`��Q�G��h�qhM��~�Bvʔ2��H{_p�dZ�]T{�Q��#�Uh٧HB��˅��2���s�O76��J� �[ �#��zC�nfQ<�n8�,0�=W�E#Q�'�l�O�l����2�y��G<u����Dc,s��y'�!�E���$]v�E-��Q<�/u�)�W�ט����p�?M5�#��?xE��v�bgT����� �i�XlxVHYEB     400     120�� ,t3v�;�|���P�鞸"�F��~#LH����M��A���?�13P�I�8��vL���� 1h{����������	�Mq�L�qP��'gv֤\���8��ٮ�o40�ÌD�_��F� �ot��7���]��g	�{��]d�3��
�{2^�y��4�Jrڄhy2��A9u�;��g:���z�(kO��鹱!-x�w�Zs­(D�d0���y�mV�!LD*���q�R�>o��UKqH]	ۄ"�,���p���R�n���/��Ơa(��V�XlxVHYEB     400     130�攓x�)�i�Bc�ߎ&z۱#��?��`'���4����@��FuMv� ;,�zQo #w�:QN+j��,~MWǩ�4�}�z�ͯ��ʻѩj�����J��@�������cN�T��{��K��e0̧���0�ۨx�D�Y�a�C�$Z��U�j,d��j�#S�������I�ٯ(��6kq򤶣A| O��χSzG]NLyã{#�a��d�`��'����.��Z��Hn�c+��}`�N�w�a��	�X&J��ͯ�I�*S�\5ӯG�6�F3RvQ�R$�0�Ɓk��!f�(J�eS:�XlxVHYEB     400     120��5����D�ݟ)�M�u�+��[űr����Uz_�8G��B�4�\CXw�wG�/Xw���
���i�H��8�>�����|���Ʀ9�(̮�#��������U�����E���g��+�l�!C�����/p�q�GlS��]��lJ��P�Fk�x=���w4����>�D�7����R�Y0�KM\�0��)��u��)��Y����F��蒮�,�X�v��������M,F���LJ% 9��*��;�R6���!�ʨ��'���ox�4�=}��v	����>֓1�XlxVHYEB     400     140,�����qM���T��@17����,f�Z���������Z�M|��6�U@�4�KN��v�XF��3M��$@׷S��S�v�����<��3{�zK�p���a��k�§�bb71ac���a�Cˮ� ,ݥ��H��$���`vX����3�ҍ˨[V�`@��X�	-&�_!�1��Z"�B���ݸY�Z(��7�M����'Εy�_��G�q�vw>Eܮ��+�n\䇠M�iѽ�/�E����X��@@%��N���S������Ԃ�[�w;֗�$��u��d��O�n�!_����s�6�HXlxVHYEB     400     140#�pԒU�͕8k�x���{�g�Iu+��� �8>�]O�@��C��"}?�˵̺R�0��������1�E�Za���Ȗ�;U��������=�&�D+߁��{Uf����UNl� .�aɷYu���������B�0�`�*yǃ� :Y|L���D�L �Ƴ��n�^����*n��r���E���L�x)K��� ���ܿ�Q�g���(�_��v��E$]�׾Y�t�e��l�t"������[��5�i��J�!�(ŦU���P�+Q2%N����hC�3�EeS�c���Pʆ�kܙO��3Ǘw9�XlxVHYEB     400     120wm�#�$���r��� 0z;�z�opH��m�b�ܟ��(�T�?s�>Cnh#����C��[UN�H��3����$ji+��� b�
�58��'B@�RC��/W����MW�cRr\Ҳh�����}��/�P{F.�r�O�J��q�LX��V ������]�U~C���T�,k�6@_��o{iau<��t-k���)fTYL
���OJ�L8z���	�7Xv�~�_��s-�Q�ծZ�K.�◉�4T\�a[l�l�e�}!��"�̖����g��F�G�݅XlxVHYEB     400     140U�<%�T�5�~�ev!eZ���O����mK� �����և���uӘ�̂������ȁ	W�+ÂA�Z�P��������"���8��C�aC�J�������%SEq��So����~p��,o�)��cyiv����P�j!XN5Lqz=��9���Y+�#�sI�z�o�Ӹ��~d_����!(:=��r?�
0/�0�p�Κ
wZ m��i�(�\z�֒o���&���˱��_�ԉ��?>�̺ޝ�����@:��*�q�'ue�
Wb�&��f2�_5��K-|��
t��$x�l,���,*ZH��Ԧ5E��XlxVHYEB     400     120�� ,t3v�;�|�H[ω�3�6��7i �����Z��vXZu�������?E�;�\83�W�Ɠ��H4�r\��_A�d�m�}Q��hcyq��fS�h�Ԧz�Zu	���c�BCu�Z$�"���9ܼ�ǰ���u�� �V�oet���Bվ��ӱ�&V9�{�\<DrP�)�rb̧�,�:4�(�����y1T�?%F}���1P�I� <��%E�ht��2:U����?WФ�!��&䲑�V����mm,3�!�=��[��=s���.o	�o��XlxVHYEB     400     130��f�p�Ϋ0A� �����E�P"��~ED�=�Tn񎰋��Y�iˀt=$Ƈ-A� ��~��k��̯� ����T�����m��V��
ǵ]Y�@q�j;k]Q�=�O�mR�S����`ʣ����У\��ܨa�2�7�w4��
]�}}�@�M�@���l4x_"m�i�B̞wSԃ��p.Ο�fM�T&��h#��lXƋ�"�$*x;�c۲
ϖ�7�6��	�6q��b�� �M��H�Q�c6��0#E4ކm
����<�B^����|q�O:���e�
L�o�=w
�!0��XlxVHYEB     400     130	��~�fgH ܦ3�}-���6>�74P�P��׹8��ӫ��Ƌ��.��mBʫ?�_�;j�A^��}���6���Dȳ�̀x#"�QvZR޾88U�ܠ+"�+��o�y����ҝ��O�s=x�+���A.^Ku�����٭}������������o[�
*��s�<95�@�<�%.��e��Uu�����~�>��6gX�lHU����C���oGu�Wbـ鸚��W��C��!�ɭ3�'	��|��d~�-� ����K�o�'�MDT�@l$��D#�0/��а(So�)m̚�Ҋ^��0�XlxVHYEB     400     140���PɶQFA�pE�R��A��P�f����>+!�oUEWNg�I�ѣGL��[�<0�-	�Vxs|���� ������6���a͓��X͏��һ0U�` ���{Z���E[�;{	���s̬�n3L��H��V|y��CZ���]����bޞ;�j�T
�Ԯ�_��H 8ʾ�����H�c��~�M�9�������
�� �����'^$��^X�hm�U��X��������`"�iZ_8�Tz�����S_b������A���v�W�ՎZ	��I	+-�ӡ������6�gN'āu�c���ڲKWM�����r�O�XlxVHYEB     400     150#�pԒU�͕8k�x}-|��jg�1Xܸ�t�9����O� c���]��k �S4�E	Ԩj��n���1���k5$���R����t��qX��9#�;�*��^�@n��j��{W�K�v�Êk�I˽�e'��X�=���s�E�������b9�4���z7-��%���v�R��ţ�N�je.�SΑ��Y���7����������l�ź�a�<����sI4�B�`�ݯ�$H�hc&v�@����Q}��ꖒ^@����^r�l0��a;�6ux.��N��k�R����t�s5����C�tI��,Gc����?����R�XlxVHYEB     400     120�H��hy��R�-�)�/S�d����sC��·
�l틁�����!�0����P�򙺠Xncw���"�a&ոʹ�����A�z)[SH�h1�3���;���v�*tUW��ÿj�z��=Tn��/���5Ĩ[�,��e8/�2�L;�_��?_݀V�7�`�?�B�^C��a��wtY�?��,O^i$���N�u�3�ͻ�[-{^QQ��i����#xYi�����̊o��v��b�Aθ/2���F
��쿊�T{��F�)H+XSY�0�����V�&9i��ZcXlxVHYEB     400     140��G*R@R�����"�SҔ	7=I篼�O.��'����#�|�￾��q��v=3<U.�%I,�� ���o���e�$Iz�w=`���)Ƅ�l��emY�&qY �ۋ�%�<Wo06��Հh�$��[�8�Zu���J���Y�3)���+ei��D�覨nԔ�X��DC05�H��k5���h�jϢP� �f{9F���Wq�D�ׇ������7aG�jFbv�)�ǩ����Vc%�>�e�M��8�8��Ʃw3��6����|��(@.`�MƯ������F$j��K�yi�]Dn��?�5���޲XlxVHYEB     400     120��V�E`n���K5]���B;��V@>r{���C	�9�'�$���<Sq%Գ�~\L�P��l��t�%
�0,6�;�+d����U^��*&8��&t@u C�{�Gs�8%�sk��KH�e��J�O�i	��Q)WO΢;`M���X\�B͵vj2���B�ٕ��ʩ%I:��@�E8�;�O�������EHB��FG�\��;���c+Fk|f0�M)�,��@��N(=�_�z��鼆��`S~�
L+u��/���b���4̇߭$X�cچE��#�|3͗gaN2S~XlxVHYEB     400     130�攓x�)�i�Bc���b+�d�ć� �/a;�4y��J1�R���s�J>��-�y'�~���q����2��������O)���*0�{v9��&@��{���(��͙�!Ht��b�
��!w$Y�oX֭�ݑ�jr���u��E$�e�ڼ�u�w(���E����F�-h7�P}+iB٭1>	�+?��V��h���Jao�=�ё��n+^��]L*�i%>�K^���8���-}��O݄1-��*�#�M��K������l���4{��#�y����c}#�t-jw�$I�6{��үWe���%XlxVHYEB     400     130	��~�fgH ܦ3�}O�ҞrO�6���QK����e������(H����#_/}��Mm���8��+��ZϰG��U�l+� x2m�H���જ�D%��yU~����Q�h��+�c�G�Kwk�\��&�
� �	�~ Ԗ����H*~����Oe�˞͗��ģ����M��Ԯ:-�4�c?����y�xi�YVO#�Bl~��P%Oc��ͨ�h�l ��`K]��U�:v�����Nr\�!��'NEi���}�{��c�6qr�6�69"L�x�>�=�׹���muYqXlxVHYEB     400     140��w�J3�"�ذϤaP����X���"f���u��#(?�� ��P�r7��h�����&�L]c$!�홸�{��5�y������w�ȊSg�������4+�5��k��$Ӫ ���9}F�]�W��^�&ҟº�$3�(�
��=
wxS�{��IP�*��:��yO�9���h!��^����K��cѓj8P�#���.3"���,$��]���$�ㆃ4�3l����$'v+�����gF-l�(���,�!@��@�����	mKዘ��P�qSB.��)G�����'q����ΐo�y�X?��h�f+C�*2XlxVHYEB     400     150#�pԒU�͕8k�xKg�8�5]��J���VY�1�@���Y����"�FL�9��V��u�驈vsL�����W^��}t��{��[c��22w*j�ɞP��N�"]�ȋ�>]̮�����ks]����z�|z��aif{C�2.iiɟ���5�<w/k�l���U�<�&yGucθ_���<*�\lՖQ����艎{�ܯ"�{c�������9�1�ވ�R�@�Y$&(һ�W��`�% �)	%�SI�[ߴ�"710���z�1�I�0�'#0S�ҫ~�1Ҿ�~���g��{�ZJGM(]? �ұ#�����C�&�04 XlxVHYEB     400     110��<lXˑ��y)E�v���0�����5:-�= Q��&�yx�U^�~c��^ױ'|(_͓�?Ե`�-�e!����u��(��n_���ʲ� �&�A�����,���Fc|�����U�f�w9��U�7�j�'�B�gr��%I���O��Ӥ����?O,�rIM
<��=}�e�h˜��^�9L����
S���![��.�S`��	&C��l�YU3�?b��ts��뮏����{*�~ym��D6z�yW��7^���XlxVHYEB     400     140��΀�r�CB��XS��@	S�ESR�F���\�U�m�����PM|㯫^�J{du����xp��q��m����:�h���v��$8on��k-�������wӯ��I� ��þ�������zD�����ZZ�#�L����͡Gꖸ����������p�[�ɑ��3�{|��+�/j5۳aZGR���R��k����w���o���ȷ����CS2�k�0K��8	�fu]v;��"�؇��H�"��+q�c��~��t�[�k�Mӳ'q��9��թ��>��L3�=��'9�U孥��8�,�^΄�BXlxVHYEB     400     120�� ,t3v�;�|�Y��E��Z&\לl�"�%��'$�	9��~������^?m�K��+\�A��㫷%�'�C3|��y\Q�A��ꇡ���`>�@�c7����~������ �}� &�L~����Z�"�G8��/?Yu�m�\����� ?�ڀ����/�ϚLk~��R�����{͗K�����
r�@�{j�ݢAq�_��T�;��A t.ϣ��@>���V�x.t�;p(Q c+rzE�Z��d��d��U嵇��%�S
 �"����XlxVHYEB     400     130�@�'��_�Jy�2�kq���ǐ�fi~������`RݑYƝ=��r��?���I�	]kAP��垿��3)x)��šl�'cB� ��>�q8�ye�V��|��<��A{\x�%L�A��ߖΨ�����beu�V��ωA�,��U(\�� �+l4{�Ǆ�i\�}jC����� L�Kj��7�<FV�Ձ(�*�@**���7��~��k (�##�~�2���A�x��`�b�1˺��d�b��[�%�l�� �2St�N1��d\���\Qb�tn�BJ~���I
W35�&y�`�Y=�bXlxVHYEB     400     1305�k�����vQ~Y=!����5���4��
�<�_�{5p�A���x�k;��Ww�b)���.>���Q�8PI�f���O/��UuOڮ����Z�n�$����y����l��/�)�B��*p����QV����6�'6�p��z���&�owyp1�4���}U���Ѓ���.���H��jF�%ے����Ď�fj��yZ�ii��:� E��`�W�8h�R���TU@��K5��>�e]���@�������P��x5��6�J�j+�G(R�S<Jg�xP�*>�>���C�㡮���XlxVHYEB     400     140[�a���=�L��Ϫ|B��̩/\��yE��ϛ�i��p7�ݰ�P��.�}�W!�WG2<ɗ� Ho��Y��=����w�Qס@멲�("��8Y�����)��&
{��r��V�E�6|%�C,�$ �m�2M�.	���ˠ�F����,߱��VuB�-2�t笯����%��Mw;H�l�V!���Oa�E���z����l*_�ҍ�uA��Ϛ��h#�õ#tp��h��z���n��AF�!ߛ����\��q��Ŭ�<%{�b�#!�jh�5#=��{x+���@2�$9>���Ji���N���=���7|�XlxVHYEB     400     160iϥ��\	-��D�*�1��d�%��uqe�e��(���'w^�q��^E�J�@ԛ2�O���o����ߣI�ڗ@��f��a�����Q
a]�B��O�f�[Mbu� �^Wnh��Vu�\_ReJ]l�5�ۢ6tb���haDF�SXU��p���󋖆�碵��S�$��6��/�"j�\h"��k��ק�P�#$�!+��|;�p���LQ��[�ݭ�=V�[��*�mU����a/��i%�T� e}�����D�^�Ps�a�*ex4�����x��̂���0wу�' $J�TG�������f&���=X��we����m�kF�2/��$IiXlxVHYEB     400     100M�]�4�p�CB��p�����EiѤ��ߘ��^���{�ާ��)H�Yq��s��9�@�7%�g�}a�;�����(�KRS��[�ɫ�ӿx�|���$g��e�Q�%)y�?lI����i�%w�Ὄ�s?JGA#�Y�T�HN�>�¨�v
�ى�U
sU0���*Y�k�\�a��Q�u>��'@i(�>q�6WS���cQwY�7��ӝ`�[�'� >���r���R�2���L���!�#{5��jXlxVHYEB     400     150P��dH��lE�Ӿ��>ao�RKY�y^��W���P9;������~8*����)������oq= ���|��d�Ɣ�6uJ�>Y�be͜���}�P��װ�\W������_Y��3�Twa��(|�(������6�؍�܃$��z:pу@U���f�r�_u<��x}��6Wv?x�L�v��fv�>ץ��L����~��jiQ���(r*I�T8��X��* ��	wA�3Ի��$ mok�e=�5���6��T�c�//x;1,�F������_�
_�u��2H������!��ú���Ⅿ;�UU��?E(�1�6�[���v�*�_W�XlxVHYEB     400     1201}��LD�K�;�����V�>͂t���y����U{�<�"�&����/5c(�\`��P�A���#q��!���~>!��'��d��7!�^B�� ��i��dD�����<�K����� ����� ����	A����(�Jfzif�F����k$����kI;�#��E-H "�6���xI$)�8J���q�y�oH�Q��|����&�ۄļ�V�dB��
�� ex|��r�$�Vu,tW�
���ڔ�g��BNK1D�UD��q�,-0T��N�.�?�K�gus^lXlxVHYEB     400     130�T��� Y;�����������@�vz���4���=v4�3��w-"���M������~@���&�R�������˂]e3�s���<m�����e \�^m{4{�]�3�����]�Z��L�&o�	z����*s��$�:Q���j��o��0H�4߾z ���Y�"5 U%��a*Sڜy*��SΖu�=_����BQu���W��f�2g����s��;���hs҂��8�f���Ã�@��Tz��60\�I�%_*�ɡztQ�%'ިC.h�,��9��m�n	�'P�XlxVHYEB     400     120d��d���R�U�!����I���zm�C1��:��UR�+d�5MA������_:����BMg]�hc���o�K�����HZ6���s�iZ��wؾ%���%�H���N���$0��̌Iپ�d�c_=gw��v"�	(�T�e���K�a���Q�tAsZ�C�2�>D7�,{����)��(&ieS5��Q������~F���Lλ�������-ENdS�}=��# g�Z���>f/���I4��X��z>bGB���ŋ�_�ŕP���Q�DJ�_8�\�7cXlxVHYEB     400     140{�pqT��){���{1��^:�ŸQ�s�&uz���V��Gh�v�����*0��c�i�}���OsN4/�s#�R{>����Rq^A异P+�Jj�5 Kg���V4>D�F[u&h7q/��*u�={Y�����s�1,4z{Q�{Ps�~�[��]��L��JW���4Z���VԸ�I[�<n��_�d��x����� �x�eܯ �����Yd�
��ł��D�#:GO�%�{I@�� �c����_�����!-�-�8�V��A#X:WW{Hw�P�Ui��-ö�7�z�;�[o<ө(���
� GXlxVHYEB     400     140��-���X�%�+ ���K���e�UrNr���cbȨ�*Y΅��!X�������\��F���w��0��Ѯ������x%1OB�7�)�lx�mYR�N�Z|�X�L�h�-�5���&r�qi��>�H�R�1�����z��˖|{��������7�G
*/������U�b^�~ǽ���o2DH��`��#�!r���(��+˙6bĥ�P�z�[���ע��d0�u���֋�nnw�Ե�>QG����%���9Ȳ�L<J�Lߦu{��4�ֵ������bVفX��"��m�*V��������P�
XlxVHYEB     400     120cN����)�O3��pgUU���7�J�^�kgT!���` W:��U�9n�țJ+��iʶs��85�ҖK�=f���m�j��7EZ��ow�c�g̵z�Hb=Nh���Y�0���馹����IǛ���"�ӱ���D��8�g)�X5�ѭ��4Ϙܜ��,]�m�>}*Z�"m�5d_f��u����y����8���'3y�t�a�Ε�2�=p��P/W~5�-�T��b_R��F-S��M�h+�<rI�u�+I8O�����
�C!�R��X���xB	� s42XlxVHYEB     400     140�v��{�M]a�$ِ���#�^�Q2��7+Od4J�F�i�.�C�m�r�r��?�3[Mm[]a23�g�(dL p�r>�X�}m� Re�r�J��h�hs��.A��&����v�� h�����4'?�fq��\�&��.C����<�J�{�"[I���m!�#q�ɺ
�?�e� t���-�8E�
O-�Yu������pq����������2\~p�u���,�$�a��i�Ƌ�\_��}y�Q4�3B�o��+�q��apt:^�eO��񯳈Oфmd��dky�dY�ɕ�K�����Qj���G��x�{PD3���ZXlxVHYEB     400     130ÿf���kw�v��w�����*��n!�]/�s��f�aӺ��������5��/�o,.�}w�R۠�-�T�LK ���ZP�0�w����ߑo���hu�0)���X��TEQ/Apg+;�5�Xp�8XQuh������9�@������؋	�oE��k����ِյI�e	��%�A�G���c��o9��&�g�$c&B|sI�|�z��;����g�IYӑnVv�i$wgCN�� �F��b��Gc~��ֵ���r�I-�b�/�Bg�{��3� !����*�I��<��?��eZ�Z&�Rd RXlxVHYEB     400     1604`_E����!��	hU K�T;�b��Em�T1��6�J�2�1a#R�Hy��&�7x�s��5�����z���I�j��]y;����˜#����S���N)��$��Y�V`�H%3�T�zy�����2���ru,���k$Q`yh�f�"��q�;0���%.g1T�*��7��~���ֲ/��������W�Y��5S�=���zζ��<4Ǎ=��´Z��>O�eZ�ls1_���Ę�`����t��DI�^t�1U���к��K$�
�*��1Ό��r�Q�c.M����$<TM��K���1�hN�U�bW��)�����������m���ÂXlxVHYEB     400      e0�&Qk�_��[9�ޕ�*?�n�X�"g�����nwh��N��~�2�Ÿs
��226,Xۥ��W���7܆s]�i�����ꊶ�g�w�cVP� KGH+%]P�<n�A����b��ZC.{�M)e<�F͢�9̼$g�Q>�������ZÜ�y�i�m�c_���g�#cr��旭����VK7�`� �A.��C���-C5/=>3ぢ��l��XlxVHYEB     400     150)�z'G,Os�vN�&�ڍ+�0��'^�r��F:�<�T�
�A�3��n�)⽽3Q^Ic��ߝON�� )��|k�~Ĥ'@n[⩻�Zl��B=�蜡zV��'U���4s[7��*����pS�8���P�����G�n�(�滲��F�\�d2n8��Q^�:�AQ𫏍�i�[t�I�3ɇ������<�A����9[�̩�cyz�Ue�J��?�<0�m�3c��*/u��v-	�5U�8�YJiy�Z�`�� �0��ǘ�����+io�܄�Hn�����u��<4��c�!#m���>��$ɋK{�p�D$��4����ɍLXlxVHYEB     400     160��?Wr��
$
rϻ�,�=������՞(by��+-�XI�j��؞#��`)�7�DX�p����ht������eR
*���X���|;�l;��%ر6~�-G����!��M;��ZT��g�'���������Sz������T"|3K�N�&���j�B�fzh���i��X�gAH��}�5��#��=}��\���~��iR$x|��(��_B�VoVK\QQ�nwM�[����8Bf�o��+���c�.�|ӭ7��ꛫ�Ma��Hz�����!��I���7ѹ�C��!״�t�,���R�ow/���|��@���Ѽ3���B�x��lH?�z��_�?�W����e�2R�XlxVHYEB     400     120cN����)�O3��p��/)��[i�|N�r�g"kCW�#���:v�^e�? �ժ0�>�뷁{)ǔ��y���-�+^�S�";T��PF�<o ��3��C\��Z��<�uw��]nQ�[y!��0���)�8P�t�o6�H0��<��	=�ՊS�9�nK���%�I��m����N�5�_���R>E�zw�>�
V�}��h`�����|��K��_G<�[r����"^"�Iw�HL\jA�*y�ff6�08]l���BC�'�`y���o�L�d��pXlxVHYEB     400     130�8�hw��2� E8�{�b�y��G��ƫ`��1���5��B_��쳭����ܙ�f ��x��'�� �B����\@N[����Cb��﹇�#C-'�����e�oU/sS�_�� �Q���߶����L�:�ٰ����t����!���M�	�!���]�U�Z-�m��Bն
C]����\M8��~L�W���+ȶ*g�A��j�� o��\��A9ͱ���f��/c������]��E\��[���c���6�M��|��	���m����3�������̜�� j���m����m}XlxVHYEB     400     140�0�I��?�z�@�I�kB?��E��)ļjJ+˥$]����7��JV�N�4{���(�ӿ��/9�p&���s�����ĵ�9����;���;�._Z��*�T��.<L�(��(0�=�B�i���x���Bh��T��;�?�ԎD��_�H=L�OAY��N@5gs$Y����|�(;~
u̝��Mػu$����a�(6$��\&Dt�=��s"�P����y�\��S��;$fYg-b�D�҉u_�V����H�'�s*n��}��W�z:�O��&c�2�N��qn$R�Cc��i�ϒ�v���xy�%%�XlxVHYEB     400     160%Ί��wh��Q�u��ܟ����R����^��ʛ�U�?C?;�٬V+n[a-���� �o����xȻ-���ą����C�_gW=��Ÿ�ȁ��:(7�ݣj���uH��;�0�дlu�.y$l�EEe�>b�ڠL�v�;�W>9���2��H�~[5VE���%W*9��r����4�F�_X%"o2�O��4������*�y�H�̮����Ws?B���c�ʰA�����Le:����Ň֘��hTѕHS�i�=P4J��V֢�˂F�a0v�M?.s��zfH �U�K  ���F�²�`� ����9������]m]m_C4��e/��@џXlxVHYEB     400      e0"�p��o�%�h��.�2���B�G{]�<��2)��ۉ�&2�,9��N�&�[�����,+3��«9t%�[q=RdG������rj�k<��F'h�����g�/r���"?��d4j$�|��7�?V/oQ�ބ̊/AQM�#j�h�z�������+�^�C� ZΌ �@.�PG1Q����2܌�$���z���]aa4 E�Ԡ�9��uT�[��o*�`XlxVHYEB     400     170�ٺN�ۘ�t��P�0^!�]4�LH5��{���V�T%�S\`K)�v9�
O7�/��toS��f��9�Ϭ,�}z�dq�%&ZP��]��c�'�_r#�;�8�����$i����G!y�lSRgo�l첔WQ�,�otu�?�^�%���h��
o�ڏ��a�``Bיu��7��C�Q��)�Zm��C#��ġ��?�P�@���[2_I��YÁDa����芡>������9ee�C��mm�֛��0n�fI�>K)�^z���(��kW'Z�|Q�A�֖9O��L�m7
�m�,������ݩ�3l� G����⢻mZo̧��G�+ǳWu�� �&�Z��eE��P("m[[#[��XlxVHYEB     400     150���1������M3�I�Z��Σu��~;H��z��޳��9�~(J�2#�r�i딟D8OӜTn��@G^��mmIV����u��d2{9�9��Y�#�m���y�����l���Pr[�eI[ ���-�]�<�zG�?a�>0�a��_�6z���i�F=��t�Q��"��|�/!y��~�?`�{��x�]r��ű'�՞,;c���u
VT�ԕ;6�}���C?�Sɧ3�o�
�D�p�V�6q�c͏s��hI�~�@������(�0��!o�9,O�a>cn�VV\�!�t���ƽ�������1�O�bu;f섿n�\�a�0�}ǅKXlxVHYEB     400     130U�Aɯ��ZmXyl�4Ʊr��$������QNjJ��n�C|��)��shï��:�a�S4?���M���<��>R_IV�>,k*�T$o��X�L"���m��Me>��� z ?s3���U3j0y�4P�'κ$L��G��۠�.BԘ.Yt�95TʽaKKx�0�!S��C=��+�p[�v�V���[��.I��Ұ^W1B��)ɷ~P���vg�(�@��iI"�i�Լ=���u9<����^�NAHG0�ǭ��t�.hۅ}+�5n*��~��i��&�Ɛ���w'F}|�nA��dXlxVHYEB     400     130��총�}�aY/�ůN�H�G�^ �n���N�(ε?n�	��j/�9��`�db�Hj�5�F��{o�����4?{����y�������Z��	��oZ�[��]npg�6�Pְz;����
l��A������I7��.�ȢH��1���0�Ɣ]�:NW;���e��y�j�ǡR�f
����J��z��l�I �'���a�t�z���/D�T���(����
�5�!��+��\����C��f��!��!�k��W��^�ql�X��=�];���T�u �U���bƙ�WZH��XlxVHYEB     1b3      e0��/�����i3�4N.����d�$R"�Ar��e�;�Qd���~���	�Ƹ��EM�H��n%r��T�W�WP�5�b������ڠ�nw�4I����J�⽵hA}1DI�$w���L��Ŝ�^����B�Wf�8���( xs`l��R��������pۓn(�ԵO�:�����;u� :�5�3TJ74T�?�P9�D�ˁ��B�JV����