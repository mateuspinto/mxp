`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
o44old+CTal5kXyCySEvcOJwoV0ksn2yZGRF9NjW1WDTWjbNbbt83qGfXNz+82SBSR/eMiTBsF8N
3ESLNBDDGDzPfpBoFaihi6jwDOPjo3i9oOLRpYB2hlLuDXXz6Tn+lwe+Y7E8+ZoFMlvcOe7Ysc2K
zc1dM4LJ9/pDfhGkL12a4ATvRezJdxCqUuU2mnVZbOvhUXl7O/T5ov1SKvo6NW4LujI9cmUX5zl5
fDMoW88yGGA6DctVUoIhAA+twWa4HA9lcJqq76xQaabC1FSJQdxXR7mr7cT92pWCUisIWMGayBL9
IYFbTvem9Y0wHbJxWrUfV+jWMsIdAz/ivKm9VA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="Vlu1pH96XUgOaJQokROm4cYIItxfPbbvVmQzZssVgsE="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16464)
`protect data_block
REySVAgwmZOnKOIn+H1ucNUu69iu3TL4L3h6nOjMY9uikQtmu4rJeRv4QSVD3cXIrFuYoqLEa7pn
ygCxlgD89emDyEintk1Z6tb477PCjyQVFMxgArg3SwVt7KZDwRm7N+bZXApZDfU16YoIB2YCuGbV
KbBFmqyA8ce5EY/Z/9vJdFOLAsjsJkBC7+GGuTgHt7lnS8s+XlrrM/+2z53UtDgAWTIRS1O8B2yH
vBjP095T6bXMRIokb1dBx5M2s7lY2FbSE0BBGnaZMaJFBTS3BTDcG+QWCqWrvE9p1Q6epBLJ7/eh
rwQkc1fJPCZVZEGsoNwLidfH2PI4VtIQkZuBtXTu9rzRTq7KR7EGhVbXgweLyiXU+qcVB5sx5qJ4
lYvKl++404IbeC8t1Mmmlfvy0jU872P+kL3/mi7PfmFgwZknkIBO1VdKSu04bX+cuwikT9zRkgvT
t0ST3cwa0s3at9/DKBsNvBk2b+HK2StAUvKBlzZJblw8j+BwaCIJO4ZTFyyjMdquBrwLZpnNb7Ac
fzd6fsvczSQNPEIn3wT4WHpjeS+qW4opKSEF9E5KWrgsdG5HkrkSM0jz/SEWNw9sTg4NNgqZZtNj
CTHbqTKBz1ngpHKISbX+DEt7P/4+g6RqIOSV2C4492ZD/Hpq4o+wldjOaLa6Vu/3ItHu2s/QlgVI
xXt7dAzUjwagLE7NEvva1DqaNm+UQ3otrhXi5x/aa+MCWK5TFAN3GMfcXDnvWxLeivSWKPp2Mad2
lEZd4IPdlYNIqfdQeCYhT4oplwTh+ZpNWs0VtsKC4WaiurSSUhYaKgD9rqA2S4qr9iHMv34KlCjN
arbE4/nKUoS2dXiFm850nhmbufjwZU6PvFkIIEgHET4YZucWI341jI3XCi8ThqeqAgs7FP3gKK8x
6IdHu1xs4m+hfdtwZJV//Yw804jnMNGv79ZGWZg7lAQr9tM/LIjtYZ+S3B7gK4DKEQmvsy6vGyjb
lyH0fXGI3T1krs1HJ3DL0XKIuNpTROHLUcj4qQE7HReH82QpBJTrhaLT2Bdks1OC2e0HKta6aQfx
/dTH3eHmnLZzGsndt7Cnvm72phYrRIsBaXCcLe3BkeJ7YlpMneJhRxEK9n3LsFTmvQFGlmgzgdcJ
QQ61KCxfnCcXkVvpBBWUbyRvjm19IbgK+zNorcDMpLxfCp3RlVD+bpnGIJeXOiTDUut9QXZqlZcs
8l/tgN8tOTo4GJMhrtpS8cDYRFn4TfWI/hQxEj5lom/FeINfehLrPvehMGpYrlUaXm/W/2/uj0Z0
E+EtkEC+C/iCUITNYu48ASaO9xfPRiEGqvfjm0PEEIR19g18Fz3HYV40F1bBTxc4aU2BaRF/kG1/
F89OK+vrDDPWsySzYL/SG191COvvV3wN8u8VPDj+o0kOS51KFyx+rWlsAAqXkDeJTfMCU5/saiNu
Wk7RMAaZ3eQTBXrNuEw+AD38HcMzBRlNw/pCyQL/XSHw9fooN7Tzl5V6A4rvkP231U9wEiGTrOs/
GHewI9lkU5bB2hkgU15CjZF9C8qSmkMgQUuSJAbVH5/jT0wu1zVEJcKZaiAITxogUJSmQ0HWmuUb
UFh1Bdv9roSGqgs5I1CHQaEgKxORTlziKCeAZCTJ5LIBK8VHbyely5+kMDKx++QzCO/OH8TfIZL6
togiaGJjrhExI3hQ92s3chPaPhTlcXW24ZwJWy34USJDxsPBDxml5AdP3jSKQK3Q+fpLwYJt3Wrf
/H52SZZpLB4x6xL6d1guvCA3JpjxxOG8opLGZwSQwawy3C3S5so6stcNGqUw3IsQ3OFP368n39Kw
E7NxFoWR8s6yDHEfZU37lGxkcyIusy9y6cZZYtM3qg+6LE4nsU/CADUE9VwV71oVQHIWuARCmWVZ
YTPCF2XbMRcpjnoDleKrCozR3JYtVOHJoodF8mtJvsZQ/eM9uIq0UPlABZZy90gqlOZkcwxNQonO
loLIsaoB72O+7yye0/8QBo+OWAXSKi3Fi5jTS8U2BY9FE1YxkHSMth4wbKRri4P31Ec8+qsxRRWo
OJ5ydPazFHV2/ZnHHd9gGhm34Bh8UBd5VU6n109CXODlZqr1x8KxnfsIXFSmRo1O7/DtcQQOyWFc
H3+Q5x4HqdtB99PFq+zFegkXAjHxwwOOo3WGWdOufEyYN/uUpsHBN18iqWIWG4suc2XiarLHM1I7
139ePtEpyyYxwGnuc8ZEmZiU984GVTzpIVXJHq78ciIRGerFrMqnP09f38fy48TjT0xeeprWZhF0
HRlMYVKx271WCFazWNlfAt1B2QocZno5Ue9tPnOjg8JYO+ukmDCDSa2LLMr+gOaICn53CPiIELF5
7BwYEGk9RzXSYiUIQOFVHp4GOuIsMEHymEHrn0psTsTjfc/mSVkBWFpRicXk13ERivXXD1p53piy
K+5uXdcAN/FyxZdPimYRGBMgTXqMclD9uYJuJnouJz+EWrfh29NBmqnQZMAFZR1y6SUiVNYvSszJ
ddr1JfHPoga54K49hJJxnfS6/+xJU+T+a0S8/XLEDZxioCJdd5aR6YORCVgNN+iV4dziXP2hNYpw
kd6VEaQplzIRdWUPQ5Ss992ezXaD5KMOacCHkvKTQFaplgK+62qPFDeOt+lQ3QOHTQ2IsaKSnKJ0
iSi+jL/fEzcH/ngfTXD5T0+YcGWAQ+g7wf+lTJiJJhV79N8zLPsKpnACxizztk9q6pURfF+nn3mp
vQtJKCNe1avbopSGR6ms37rUKZx1GeUKRno/xJCtjCU8L6UDaxCbqhkMG3I6YIwUBtmcvXkplg/2
npjc7bnzdeJzDUDxhXAdgYbudnyj9zaJ1YxkJVdg6iDWEgUehfdM5gkf9T96bpj/RgebxW7n81yp
lruLtxXmFkfuj39mSbyp+Cbth3D6NV24GCiuTSlK8rJHbblAC9DBn5bx9sKlmWKzLVooZCEUgW37
UuHV1YbA/UsYGjGC5/eMQEvxR9loX85jITg62pnoOVvR/Hd6XGbCtkm9Xm2k1KliFthXkrsvFxXY
+KSE8lPEQh6tKVNCdPSoGt7VJWaXOgCRPbooszBExniNrPJszQcvVFVjomd59CgmrxSwzAi7NAIW
PfxXFhQ2sgK8UFrmYhYUPSy1WcMYmF0TqbzQTgE9v4ZTGWBox9zZY3yrTDDJNFNcHgcv3/hOew8O
HihR6WJF3bEHpdeL0QlGgdPOF1noJ4+a+t+fRiw0IYLZ3XaQfonooRcF89UUnLQNgXJuVxbKfcmh
iV51KGje4Ebq2YhUgZBAapP74iGYCMoJkDZ5ixrxBFrOdKgVE2QTug1/O9wMa8Byn3RINzFLCtOR
1QjTf5IxUl/plYXcFj0SgvQBobovmQwdAgV+YP74PSQ7sQGAaRNHJg9dqy8R1AUq2CjUarAJmQEw
wsKGeaSRydpgxufdPuumSSzcdm6xNeO02pfh5jmobo6eYpbW1t/YdrD93xjq7u8a0Zgj2kK3tBWB
I14xtyF3FwYLnem8rB3tKTFvZIbybSjK1Q9Buj8BF+HIKirYkkm90bGKKFwLumlKFc7UDbgvK03d
zet1edFRWX4bem0aelZgts0gzuotrIkqFT9vpilJJqj1C6XA8v9ocrOgDNDzhS51InXUgM6lcCTJ
Jq+DlQ9IkjCQcFJ6R3ywuVPTYoKtj+SVqPj0sc0+Y/wsTPxJF4OaVQUbqV6z6Jqp5yWWPX5JAMSf
FjsE/IPNlmTtvBq2vtX/gPxenLThRg1BGSlmbqc+NlrC+/x/Q/1ELkmFolVnHA1ee9FAbZwZi+7P
371ix59Flq0uyar8iD8omZQWJ3dVxRMk01TG2wh57FVH+xsoYipH9n2i7y3nuUpTrpweEGlGszjr
7eyDCWJqnhfnHIhRv6h6JU50GXVy9e/zFXUqFl+AzUaFjWnSCHZOVtLM51MK8QSqGMifHLALq6Fg
7t+9A+S/n7cIUo3dRwZtX+Sxtze+9i4XNhqTH7ijsqLtd3/xwU9lVO27S1T4hbLR503s1dgBDXlo
dlmSZWuihPM8i6Mr+UOdSkkFOpMsyjnb9Jl7dOotOfRm+iSRNHYrWuohR34MXBigAMxLpuQFamtb
vtSlhElsRxZk730p80UdBr6Y15hhLRLq+3wpgrAg27nDYTGN5nXA3Jn4DbjcjdQxwMqU9JxpsZjG
4vc06Om/JqwWK+XWJGczRyWkUx0YKkDj7nW0or0TBK5XkcMoeMHG4UebgH+2DGBxFC7cyEZMnz4v
6dbiHKAXYNQRTfB0WSF/2MhiMYlk5jHeChPG39IxgoTSa31KK5NQsyk9YeawKF0nhIEXXPspSCJA
yS+nOacdgHUr8M/b7tcY6oC5P3bxitn9iCq2CGFNNLCtkIHKUi6SaI6mu9nLkWdIGu+h4+ktZKC/
ZbKUs+mCd0rtAD+32bF5LDdZuHT3LtJCkM+7MHHcN7yJNRzt5jCeiqsku8e/9FOxlkPld0H5CjOe
CXuz4I1wSGRNGr64CRW6WiXVD3zDxAEtTlPAZVpo0yvfurrNhAmatW1ezOQlenOfVvE8Ub4LFeZF
9twl782WM3b7cQF+kiMeMbYXqpAqKyNhRi3ph8euPgIH4AMXVp3OsyJ2YLxvW+91efaxwQYtPCev
7gnU0PZUeFYR/iCwUbr7Ds9VSyuhsFwU75aYU68zxqAyn2ZN2c4bE65xRZnSb4ldfozgmQG6Itu5
Ai7N76bQw1VHC1GlO5ZC/0ygwhAFa/E/zPnk7bM/se1IzHCidGYhhqV2o+JoKwZp5znZAdU7tQou
+dJ+9TVJtTi+ONROx73bzhZvJFZwZB7KncMKVNDSxGd/zpsIp0/V1kM4tM/eGiV9zx3kQ//a57GM
7NUFmkwq7QzDi0jukyxBbXEx2AcGUCEcAsg9Eq+K9YsDml/u5494iEDKerYTAbtLseX4/bwUM4FH
5X9CnTkM999nrDENKHlebICLJbk5Rv8m/gvH+ZQgefqHqAJqkRM+zbnY71Us88gad0TImeF1WTsn
U8rZBdlOkwdxIVxIzm35Ptzsqt3Nak6cc0uZksdaTgOS2gJilucicnoJbZiU8VQ7rbbiZf900Gp8
MAwoFiwLfBit+vxa6d8De1ObBoqINmg+d4wpKbAXjQvjqwOKArwaasy+6jGS/HJN6VhokLK4WUok
Whdr+YEtQEP6mt1FMyGzk01EM7EMzlxVvg/+F7BUCmoa14GpHhAt1I+riqzstSWpywnZsLHF/k+A
HBnG/T9PBybe6btoHwnuEae2vExlyTx51KhKxQ3SJIsupxX3f+JHQyRM7C9BXhVByE8ZYUIR836j
vHYONsQUVm6t8PDEgJUCtRUyD3M1op/GpAqC/JOItbQe+3GkTyUa+JcGDrjhaitf5LVe8rKN2N+P
EyNyGqarsz0KRloxYx/qbTbFtr9GlVj31Vni8AD8+vDyH/8Up7S+LyyI2FzqQ6BL5w+Hoz+6IDry
f0/XYkP+lbThjflH6Z0rhFM10nto/TFpMY3W+cQFyAf6AOYQ3LmAmLkm5iVSdg5SykzQ7mVcjp12
cmjZ4+GJdgI9OC7nJfB0Imqtncw5Ez/T8h812YYPYo5E2yldGInQm3uDC4/nAHjkFJLR3hrsMbHu
843tTHRg0GfiBfxqDvzLExpHQ4hsSB7e7Q2122LM7dadIsaMqBb5hEvlLPoy3A8PWfcxZVsF60pF
+ddDfkc0k9Jo9UJ2qtT0URzcP+brJZaHf4nD3KzBhEo/zHbv6CmBd3gGL8FS3S/sBBtSITJrZM40
IbvS5/TjCGdpve7c2/z4TT4QKci9DztKaXQT+XUwOllErE9/+LthDyqVHvv/tjvfTmfqOhvWcmRr
PASUxqOxXN3R03AhutzCPKCiyJIU93abgnOPvozOjApXWgvOdO8NAQxDeXaZOeWRj8cL3c3DJADG
51V5mpLQ1MtO5tzTRGilr2G7gfd1ski1RSNqv+hPeoQPNSklPlrDDRzcrQEQn+ieVSudGmVnmYGD
rZSqPtHKHOMRQ3FyIr/LaTkDYCvBLHtLBWwT/NliOXZ92JYLY8MFbRCByQKal3NYrFcBvCkqcpil
RSYMuQdJ1d7FXiuzv2BAl48xtENOL+KEiSa9QicBaS5LtnNwmoCE6i7Aamaq38i1sFyKbVrBsR5D
Ky+vVvXz5fvJXV+c5Ns81S3+NFoEEbeN1yu/vORNswnu7e/XkhmYgEsM201LCrKeog4HtBGsX4tU
UbnPV+Dr68LbKBXckHBG69U9+ClgKv1vO+mxi1T2VdCii8XmXxx5clcsKW7wxyrlWutjaEbcMOIi
1AbGDXKhaiuO3i4KJuPwfIlEvph1WU2DWxwgnLng5EMLKaTWI5BpRnGuw+4pbAs/zeM/dlzdEBlw
+JfoKhpS43HthsiUaSi/mEMFf+5kWBuQorctoMJfSE4Mimbn6XGebWNcvLbX+MsHtVvR6IXEx8My
eb1ZLkMzkFSbVWuOyewMjfAXWnLNENoOC6jU7iDQfEk8LBGpBoQdNEwHDbne4KAdgtZMTCwcW4lN
KP6EDWt2y2qyETBpVZiQLddwxBSKJIIZS0vwtTgLI7YREeQLuM2CT3eAPvf53+Cy7fZ3pnvp4heZ
shqmJea/B+obIAQKsagRkrEBgtTjjSC0Or0DFJE9IvtzbeHi+0zNT1mD2SsmAoMLYgYdK6vDVlCh
EIMEIqLrpkHTuSX4gQpwOPxaD/8psl30baqgPtKx+/Dg+o8auD31IxiQRaFi6Xf/X0Ie09xMBfp9
tufYcn8mzeGgJp3tAa+yJNMzdPaIb1dUUh/Lx2B8v2tCRpkIVAG+SCcNYI3DI2kH1gVD6noZz6wj
r1jvKFltpb/zbn8Jq4nUfejG/PoWlVkY4oL5QqiVmnac9lrPBqbjRhQqud6ZnL3REfWEoTR0vlM3
ogZopdigoR5wvsnAowAA0latPc/HsZyTsxAKlbaB0u3bVSsfTyn8YnjPfRr90f17WSryjIn62Htj
TXV9UoW703qKheVt3fVOxsyJ/57tHTiNwxAoBYfI3Ortd7DWLLDLiuoUzPC0yb3Fa6T3c9WiNGA9
SSdiicOU2/A+ZZBVy8+g2IYGW4wAIeuAZWa27f/MncarnBiddvig3vkF7WKxqWHD2y05F5+wgbwa
+F/ctRBTPbg7KeHOUjL3KXejOBK1OkjkO+D5VAb2GM1S16oRa82KgyOcU+pu3Qdlw587tYHEJubG
8PAeY5bbp0nhKDjqbsBHQxZ4HMwF6U/otsrkP+Taf078Z4NrmlSV2QrWIuzKuKF4B/PsOtKZDaI/
s1mHLQXKLaHjCn6+IelrwYx23zK4+1fdkG1k5fzIIi5w6gCiagR4rO96I3MNPw364In9BnLe5CJA
GWISNtb+9zX7ONM5nqhIQ7RARWbErBXlDpteC/9WhiCrX/XuMdL9yhW+Qke5jkerfbhHH6ez2LVf
AzNwNyfjRXzhmRi89SJ7PikqcdsZmOy+21InFJzKtTWgvhpRji6W94qVxT1b+Cf9jb5Od2NSPiKC
Xu9C/hhKHW3+PKVGHLPMTSinHaTYcCZTHmrlNtkOdSl6H4dKj7TBCunLjgI4L+vSIlsHl9mt6VPI
EKZgfGwzF7VddDBdSn9UwUtlPRynXyGmTY+8kg3oX9eog5KRXsIaN9vpbvThSQAflvA5rOpySk+8
g6OnUnUtWLgHZgg7Xt9lYywJlpf2auxe/KaEaTIJUPLyd1jJdM/n3krpX8vqGTtxwhyBPJi2/I42
gET8NT/zpSD97kM83s+J8KSf8S2HOGl05wq8SnleojknfsOa9VtvjgRM+MkwRkG9ETPYVFFM0xN5
Rcz7vDNPsZ9Okv48ncHmDd/CXafjA85CX4jcS9YAgHHHyHAd7r/LOMtbwIKXidcCxuSyYW85AcpP
8ct+eyFN/Uf027CXj75wYnpOVdJHfQB8DBqvUYlsWffYa8OTTAmLAmCt9XJoSb059dcCPG5j3z5r
k1hZAglysMH5wEnCKJE9nD2C6WJL2flgkQmxNV4uURNyWGESYIcvxQw+vCyqCoAp6tzPk3q4op3/
KdiYAJifxjwNCAhoFD/FB6xsBvJN35gJpL9qchhfAL1VyOZjPNc4Equj8p+qfqUDFcI7HUDfIVnN
80rdzqkOwhxUTtnVLX5tXrRBp0hx06vKPZxioFXKVsJwPzyLS4VcC41LGILiSl9whTbQtNUbAl7U
FDOdVscluqZXudCaKQZuZg4YXntKG3CRbMyo8F+q38SKO/NczSDJs1wpIJLlksbSPVxj2l9qOKDt
ARw4zzg+rMIDtZWJg0mTAYI5CIt6p91UfHzgRMhgUEIlfNgpeGx5rxSFtb+YmcDin7VDk6fOn4yQ
59RXEuBEjm87ElrUIIBpaA4jJ6dM2XXqifWRTSIOBOhabHNC8VSyXIKs3AxB72/+UgPmNYCda2Gh
MP01x9R/EClKunot+p2cZ4zI5+L1HMxMjMPsqLQ6dremXSW3pi+O9JAzeqlBVm0vpn2xOAOm95sZ
ImIAo7XUssOQ3NodTmr2gSkAfdv9OMahhW5CsySNMkqNYh9XP1+3u1FgYfMF4oPqptFk9MS+nqS8
9qqKJsblTAJQ8VLKPfTf/HsEM5G83v8JdbSoO0IkqW92X9eHudzbL5RewUSQZHaQIr/GRNY+Cwrd
EL3zGiILEVByUixEazAUyJccvGZao7IkDd4c4bmaOMc4rVDZLU3FqxVd0KTOjJN69A+tGMrg/Elh
nWKn7jDYHJ4iG3UqIoBZ2zecZQoylvUP0ILIDARTBa4ohT4MYNf3K1BNbzJaoIgp8coaGYJaabQR
i2KfDFizZOVfopn4dF7a19jog16J3NuydY0ZntC/e77yKbnbQZyL6OFgv163lL6r8jAEht0ymR5q
fLl6hCO4DOx58KhmKKgSTLHqxXSvMcS39kbKSKAyzwg4r48cJ4JrjbHM/YXVqDKRH3BJIKGkDhYY
UJjnhrsXv0XH5iztg+DC6tqVcnEyE9acpNOsdbl8Q1PI06MzhXfNKFhlg5xBllEZDjTYyNqKUddq
eaXzPJkQRwdwHS6BiKf26DbclpnyFJKOBLm/MqriYVRHhiagA29UOcDlbIdB+v2f3NJCPSUL6xul
O5gx3GNuSDqrwJ7Bl7TZtGoY0Wtx/CybKyi12RAIxWfz4wTGKQzcDKfxsNnBY5XpmWuszHxMqYX4
ZmLU0q+kLg8jI+jcWpWRpIv8blY0ZfAv4qiKIW9TU00hu896Q9HvrPGSXWRnINkBBuBXSAB1JCq0
qbKKtB5YS0jxRH2+yZDId6xii/MjpGixwJSJdgMVcQ9T8Drq8PkQJksjGlqkeBqxqZiyer2qBLIt
6PCLj+QIZ8b9KjkB7OElv6cz11nAeLcs1ggHHxzyY50+xqgmqtqUgrD2Ur2HIHYxsRgzohKtwPVo
7FNgNz6byw7FuyHdUE7Zu8/aQPZ7r4dlHXRSM/hH+gvwz8IvRemrEjJJNc9cnIDarYGXVr3PD95i
Ar0xx+9NB4KLYqbeI73bmYfwah4qIywpXSeGGh4b+VDRI21ZW/+8xcEtIf54W0WdzB1Ue1q+fMJL
H+wkqdm9slhD/jtdYsBKa286sYH5W2EPub897pWdeS1CUVkh/LhLjtdXrAg+L1gHYpr7PoVXmSWB
dHehcRpKrFtnGPaBgNRTuNox6RiHYdPvjs18Yt81/pn8X1eQYHVycG2gWBh3SAjtH58ozZ2WdHYC
Zti1ejYk1895/N9tOpsX5iOfGkxCutfql/iJA1jjPK/mWh7GL5DJ9zQabZc/VbEGNP+44JOtqIKb
IjEXC+t8LPGD8He0i+aiapV3AFiT+ywl521AiDS0fiiirTWNJG4kbsQEescasfzDBjFMSsBdl7h6
E83asujff+1fttq6fBxTAqNrO+AsxnAerRJXhm3ssVMJlzVZM9DYFglDGEk7c750+ds+KeNTHF11
ptKnglRiQ01OYOsseoZ7paB7k0LCejxTWMjCIENRGzRDY0AW7duT30U9Lk6TEOjayPaXpXNR3kQv
ZoqG1jnxf9iocmHKbRG3ZoqDyZR5lIo1UvebjZSZgYeTR5SC1tDR6dJPMMgBSy7UxnOCgSMsCR9F
LfbOiaI2u3U0Xk/tv1hDR2u3iW2InJiLVLv6ZcfzzbOabpTEfUNDWrsEV2S++Ee5wIJitkNsAGhz
FayTE/xZG8Unrw9zOLLl5zviJJ+cq7NhZgMfti9rK5PrNj2pM/fnQMLxhCCwF7sPJRwwQCS3v6g+
PzLwmJrnL+owI3uGUy0eT5DFk8IvGvBdCVkoXCNd05ExZFzVqcotTTS6ENqZmYv9pBI1hDZ709wA
+3CUH2xUdaxKaSFz5/9KAA2qQcOIfGPPAzKtBBRin1DkaUDygadQETtRjkd9yTbT/ivVDEVALpqL
CTcJX5NupKnM8Pk72rTQXLN35RXUE0WYW88xlKzxEFw/GzPU8k/5rp9R8ekKn58FKTlPk7f+KLRU
cf6vpE68lKTFCWmZN4d5It+Kt5jp/ZacLvkkp8DBG5MoRV2onXCEIl9AEwzO6NqSzDhyOiqG46K1
UQeQdD+qJJI1v1rsrUxT7zDJcWqF2Cwlh4uMTih4XeG67Xw1KwCnyTWdT9XdlmaYjSXdV+Ilt1uE
fQk5g/ttFK/jfifg8FcHNxMo99sCNu4MnaFv3l45yzXn6+hdign176Brt4fk3U7yVeCQ7n49JNn4
w0F0/EECI97JkeOi9lKk4jBaiDlv8VdaznMT7eotcFybtoILFWO5D8G38wxTBq1AjHNO6Mj+WZoP
QMOWn/Sz+O5c+xw8w6ucxdQBWsO5C76e8uM1Aie4LstELDgAIhAgyf8fOvN73MyZqXFnPMmP4GTb
n80dwoB12Mr2WoUJtfIfzP60YoXX8+E9x2JvVJD1tlwl/WRdou5zaikk9VGBl5Te2IjT3A01bttz
irV4z5ePHxvlDNYkf7NM4XzyDeGgeYfQaDWcDIaG/TBdTJrAIJJQp0JGbxkjvMkU882DhqkifXty
TXM6plW292wfzYRAOSif6yuN9AudgtV0zvzJy8zTa3Q1EZNFqwMzzLaM9wZF1PW1r7VQOwDBuBEY
x83ICV0v0y2PQsmqZClLHA7XKzi8QpRlPmi+DX5BImR1Op8PhGSDjqLHPbCNyJ03n0MVdwXH5i7h
Iu5GUaddEc46YgFU4SIaOTSGFCaX5r6+MDdTtc7dS3LPLW+LcC1uiemnQl+IoslNSRJUxGXsKUiL
U6g6AXnv+M68JUTF7X5Ju5cuMXBPnrrC52gtZ7hUqV46/LnNKEg3cPu9QJFQAR2wh/euzJYgj2w8
sswjc7Leqze1CLXv7h8LAZ7RteYAs8FkXCjvOc8n6RYvrBdtu4A5j1ybrWhAOpUBlBOb5NoDTc9S
/fa6OJu0ncuxsL+qlML1TFrzQ20ZqJ6uPYvYOnAuk+Wmp+XG14F54QfFl4Ujlg1ixnxbtuV4i1Ru
2otT75r7zi6twLyb7+Iqr5ZMbxr3xT1wQnVjw72lk3MBglwX9RLKBLfbcVYdoLAvlJhhCF7V3IfZ
OoURm5I0x5gIaL4lixVAE8bTz2hGSRoO9pQBITo9CJ56pXd/+Se36JQXYIyF8KIOBxV2ft2MNXjn
BoKbqfaXWHezY1ZZKS2RK3w7ICwoc7R09+7C0GndLZbwjADiDvwErhDKVWZmTBKAFWqropWsjQuQ
ul9ewGuECiZKsXZ2BL5/KVJuRY8LMZE3EL+Fu13Ki19U5mEpesSQ8sdicjyP5sxkmss+DzB/wF/3
QxNm76vVgvvLmgTPw4Cn4LFe3QbdCreVAipWNOwIMSHblmhcPvQxZnLhbemxIVfLkpglaTD3TSgQ
XCvwngWkAwXzMTgovItPIAZYTYcJO9BIWnit0vwlw4qoRjK0PQRHzxg+7/F33/YwjCoUeaI9XfA5
HigYlKbqpfjREyJ1DGOS5GflPTarrcQgDgckoCDaIhYdTPAmoHYmO5gvNB24ozIRMZDw64s6d4/9
P6F9i36xF6P24geeBXnNyrxIO0glMoED2tOeC5YyAuE5vIZAQBVsjMNb+Tmvd448BrlhyN+B6zzK
uNbRWFQpqa76nYH87kG6TpzWBg1eVHaRZSU6QVHW+X/v1xc5hZh+eY3O6vTl8oj0mr09r0IHcwOy
TO9rH8c3AyAGR3KmKmhPB026Ysw4/aAVhg0ujuo60L+rc0Iy/Vw+ux6613ntF2ZtEQxXIkt3xEBd
qmDh+i8bJVXsWhSq7vtLDBEOvPcmDW2siCN64rkoqrSBRWF15eN/xX0NPkP7cJg5oEP6vdmSCg/Z
2Yj0EhnIkNdxrFoIBZ/JSKPIMfAsLxvCwRH7HfsjnPjvVTW4HH1VFH/Q9LcdbxBIcqfuYsw7w4ne
VTPpYtDBzvRHjNlwNvFZBRkcfOn8KYQYEEO3v0mTSl/3OI4t+JK/NH/1OHjobg50mK6DAn7z3qCa
vdeCaLL16kcB4q/Zst/oFRJiVcI3/ourJBprRal8hpFqh1yLTZY5JIuo/SC5MpnL1THtjXVWUyQp
UgC+pgSj3YxdtSBBdaNRyM3BcwhEj2JEDJ1N/XsluRcFq6oP6Ti08icoZ8XdYj6gPcvess3CHZHP
1HPOmh6f65I7Jq/VJlEJzjyYi4A0AnIY2wN1MCRwne43vhbVFlsbXIlTnhmfzrwk4UQ4a5IO1dYC
fFG/WXYgVQ19ASaAbM5ogjNxE5on3X+gxJng2ysoC/Yidx3IRnjINkZVNzlDnKBvUzQI8HfMTGbj
cBGWUxVGT7vmsVjIiscUI4QkCjr8c5ytHUwuVppzybWmvHpiBcfE5VOz6JVQeO+zmViJ1tR1+0o/
pv+GLxPBzl+FJt9RKXsjGySuzjUx/VfVgytj0yYwLevt0s0Xiq70oZjqf/uqsNpvUEfnkXE+f36Q
0Aa9eZx2L+Yx6ahIbPwu5KHMGrXjP17mR5qJHp5p1QXSL7iVNCbmeVlULSqBCGEdRN0R6GRjz+Od
WfaBmEROhkBjtglqidW2z/mUw3Pz/7c47FmEFzRSUkixRiDLfnmg0BCIDRcOtGAWSA+TtoG5R2to
w2jd6v0wV59/BmofWjgLJN2X7lZolY5FSyK6t0pCv8de1ueuvh80nCUln92KC+CYYlPDmHRHCctp
9tTjGbuf8B9xS4tejb/wnFw4tMJtlJEzY7jeZl9bQS+rDnDsHWZrLH4T6aCdg2ZSgZGRNh4xdkVd
XaN8+jlkwFw62Q9XxXanuFJ5ehlHWh4k9BshiWfY/E3I89cedFqzVPDGtJRa6EaZe+g3IRXoCS/A
jyo1WA1GxHr4Yzigke+O0BL6mNMyW/jRR0JnsvbdxJUiLq9OvLqK1E4iZbrq4eG9vx8r//Q9SJaB
QmKLnYCBBHq6R+xQk0bPrJ2DnwCaKGecCY/O5L6+zSEjF4K4qTmld/VXi+ZxXsEmqE/FRGJdxbDq
AYlt62F0r9P+fNfOY24yde+iwxhwv2RuUx7TfntM5YTy4rTM0AA+lsyEWDpIB+5uy3QxHMTuN7+R
kXwc2O/HJ7/DwZuyfKE6x+y3bsc4bxOGdZSSHsi8BImzj1XelT0a5fKl3J0L7bQG5TJzgm5rKXpu
po68NkUIo0Ze87CXZX/c4bfLCGjwakoPJQK9xpjokI4oNlpE8tmVxAHxflc+zpYkt0aqbEreiB3c
Xs6tdlTYdbcyWEDDQ5jNNW7U6lEAJvV97x/Whrem1tv6JFRfVN+bABXTxuI87AnhXIzcgVNwES7g
bzKXycKiVEGLJR4ZB/UpzeEAoqw/In4M7/RG2/gwYn5GKamYzEvrTMzU8h0fjGyc66PfAXgRDi/2
eJ3mz/D0/JproSPsO6FC6RbFLLIRy82QET4arvC/N/lJMLMsT6UNk0XpeWx3+L/bB6Y6uHLAiZIw
3EkwioQqLrIAiN5Huwe6EAgN3ZB3ElaEIjC/an4fSJIsvb6djWH/f9EhR3j5jKIXwrFqQrLsX3di
TdWHx4TZGCBwDdYTlc4cLs7yiEXxirKuY1h+8EbZ/IibOxKOl2ri3L8UhtKaiTv9ZFycfpJb8TZA
f80PzyygZNIk/AaZZFbn43Gdv0CbKEB6ei1YJF+GHIGZzI6HZIGvkL+bMsh4zWb7nTZdLEQpsd68
w2a6KinW15kA97I7oHiOcu2xWeQoQ7gIpf1lYayZMgpOndLAIe7nMEezHgpi+Ihuojim9bYbPmxw
WuHGV4oQoRRYnbjgA+ngOwBM2K5aHVyUvDkUxwDzrirDkQyI/PLeFRVGsUK6CK51RkeS9qAmCJSL
ftZVZr4JA6b/dZxCk9F4biZsymq7guiwv3aQ64ZDl4/CA+tGMt2XqHWJJZi1giQaBCuYk5knpJbi
0pF2u6o0UsmZTBu4fV2yL3MWcy8IvlkccNCM590TlB2GXUtHxJChztsLtyp/++rRvWRD5LBj6kuq
5NTGsJIaidD3QIzS+Kzp86V3qnC/HmaDhw6ItwuqNi5Nnx1aPopE56OnXIxfgQJ+Slz1eleJgyjP
AJtNuTQ9qIMvVTgyZA/p+jLAgG4LoNr/L1Nxl5tiZv84IcSNQTO880Aak2pXcsHdKsZJ8DarCpC8
EiSMlpMvqBf+48H2f7Lig9z+f5X/mJ9awa8tx/nnuLu6yagVGGHEOLvezWR7Q17setE7BAbkp0xO
7B2xhmykAcGTQ9eLVXcdV7bWs4C3EFH7kSabs6r6NxzMR1liEmqJ3RlSNfwYFV6myxYZMxXgdk4k
1l9MzsjDSJV2f+m3F+uNt7tMaU5ZUNF6lhxp84jNGIPqzNeaivEMqGtvlrredSVpKRrkY6mI24fN
1Z3sW679V3hdivaykqRoCPYO3pSmskH0VfXqwrCOhWPvNXPeOT4R4Z8CCC94gvSsbJvRq4WeraLl
GChL1UHMrJfz2A6HA+kMxsx2wDlKMno8dCNxSvHUca/JN0UfpZVQ7kruw1tSHKtoJXkTlaQFAT0w
6J09lxoo6Gci/543yBi8F213H7FQgi96j1tlgTJYWTsTM8intlsBNX+lwOXi9nj/KJWHPdYyJW8a
cjmvVLFna1rGuHjJdd6oi6inGc1+En+62pwj6BUt24mJ4I8M9cjR5rVuxjYUKbVv3L49peMGwu27
LHEK5nIr4COWvLwfaxeeV125IFqvov8G3Fp3yQ4p1/TF2RqEA8GGtwlo9UDKMLteGSnVQRPbWWrf
LWwxQ7KjKfs54WyjMHViPDQg9xh/rbWUkftJXPZF1PqWxYYYsInpAxJvXAlpuCYroVxPGrSE08JO
PvifT1wjoiAXCj2Z3cNYhxy7tlWmJ0tf0RTofaqlVbYFRsWjrId40q/jU2YRMFe5+9D7bBZij77M
eFjGo3U1AUqtS+feezMOJwroOD5gZk+RVDlnHAr62rY5p4n00DA/dsKYh0zuK2Eep6a/avdmqGm1
IVu/tPNnnldUwwk/ve4fHC+3b4kMrrJMepPmjQD7a5dtAIYcbqbhE1K+d8ufGaDtuaphsub5r1f3
jwTJduBY1LK1MWdLbaklGDOJQIXPELA74wo5+/WTa0mdTJZv2P6S5ATozhWFvU8yW2OE0NWK8/vb
01TNDr459ALYJX1K/l6q8htICFK5TAvcwYpoBpZ5OLGbHFA68DTnn0tmyAjPaEFw2H6w/hSFL43/
Zm1n1UAjqj2APghinHuqcgcyjIaurT3vJs+EC0Qv7NLUOBZlKTo9ItnQSBh9UWYp4iOKS60bIVFC
+csRSPVFHIw0oK4JlzSe1ILM+AWogLTRYepNtnLUpMGmCWqRl3MsWkplHOCkuvq7e8iOJTJzGOWL
fRhqa4B0uPVU5Yk4eLGD4jFwHbSYSSc9ClPqM7vccYUaXoB7RnH2VsB3BuLc5aJjt5wpdAzNrH1X
wGgMGJiBKitsYQNhxDaXWh+4RbXIq/Wcdrqww82jRdxJ9lNWSMXJWEgVnn/nqnH3o0W3bkQCMztq
D8tV81/1TduG5/5v9Ga04Qjvy7U5VIZDhk4s4WK6S0hLbfllAHcwG5iXtoEnlX35q3iQkLa9S8/+
nb6QpVxnLpV+/kpu5WT0Mb31SJm76pjhECObtNdwzkwg/eFFIGzoL7SKR7JKM1+1ZtqkunNXa9hO
YqHtWF1SRAMIfRtXKwUczeN6Oy29b3OLRKc8KZFA7DCEXGZUMjerwL+AciL9tvWPc58Qi7XEsUxY
Ly6hjufkCA5eASfBei0maklQIgXT1jSc0WXpluDPFzZMQjryF/1bcAA5XiylekpAcojYYbaFX9Uc
1pmSDkngYVjCTPEeAmqwg0rx3VsQs9OI/H8poHvTxnHzhxhDlVu9LO7ByZX7jAVXUHE+P/Zzvs7B
4L72hVT0Oqs/PkWjWvWIeo4r3IX9n86jRD5nAc1WrQAB/nz5dwOmsFDZPyIq6/Kdk0LbUJ6qVhp4
2SJOuCI+7VIXCehANfhZNUbm5bJNgI7/tmUHeBbPXyzmFtsShQ6F36ARTpxQn/OW55EYE+hY8DLD
dkcgXF/DG4K/rKEsZri8THF7s8+Q007t/SclQUEDQG+vEly48gWQFgii/7OOYZMa4on79QBjSvgb
y8EjsOGS6IP/Nij5xijBlClId7etKvynXSEktpWGwiGZAUvMgtxnJ7ebAP/VBcbAgEClmooBY1lp
enEcrBoYvsWh/zBz2sBdbUlWrTguJscCwtc+SP8/Jv6Mqt7Uwl4QAubifeu6wP8eb/f39q5VtC30
7wvIwja5YnsB1A6aG/SmQQpD1cg1bCn2ZV5WyO+9YYFK6uXPSm6/xHspUlmguA+znp3wgfrrvEnB
ikY/k7SVVulkZEdbEPjFBCnWIyo+INb79VZE4DRMpC/bL6T89iIJXQseKloSii92G2wTGdya1Ttj
VRZtKt9Xzw/87sZYPEIkZyjhuhowzK+KPsXVA1LESGrz4shP6XbNIASVXRaRfVbyRT7dkBna9weQ
IADIvSNPlkViwLIW3o7HacQMeEDGf0T00BwDG0xBQqCEkvkWLWMlEWDde9u8Pza1jhU5sN8Aj5UE
cQ2zmFLytmMF0E6Sl/2R+WrbDQpwfo5Rad/3KJQzrAZe92y4ijQCUTaQ7KaUhTNf5iH3uvqG9fA3
NN1X9J7oxct/pI1RftIZ/tSqoMbHcF36QSXdo9jMtcg1puMclUtRlUFYuk+/XEQ0BDY+IMw7C3aH
0KLjR+8GyD2THuv0WWz+3sNefZzqPbT16J68pV1Klg1teNhn7lNNlEzZc8dDKFKFDOMnDBhA/98b
2+0XVojFJoX+8h2KV8Gq3YjED3hgM6A7fyujc1IAV4k4Gy+QpW/yfytAg0mtFTLwCvZ7IUVTPFE8
e+A1ErntoSIvKO/DFR3dF9b86jXP6SYnfMFVHacY2VnTpCUA+PZ487TUwBJKfuFrbdRo9s4eX7zH
dpLdit1tPvmkgdnHeouvTFlY7FxWDlWXU8PDlK1ygqmAXM6gNvhsy7QkFjIw/scCv17SEzeJyUA9
BtCYajvhx/f3kZnHFBy9lYxXLmn8GEAq01GE6lciJnft76ZBf+c75PnhX4o+Rs1LoTgZJYihF8Jx
eqE49sFakO7M77rBgReGexZTEZ/dnonDX4Eaul1inwePOP1iz1AUF9x7xCuWgl0LV6z3nikbB5lE
D/rQbzGS0GC+HLqdXdcAcV8GU8k4eWh45Dl8/NXqu5aSgoF4VGVfEWgtXvoI2vqDTsodal4cay3b
ugc1WpGOiMtvKoJlVcXNIakMvctR7FyO8hC29GIUKuHoF2zNxpqFrMFBygdFVJExxb6jOCggfezT
QdxaIFrJzXAVVU6C0pMvrg3k3IdesOJ/z3UQ8oVsszTrrhcYYokD8pND0Xh0ACbGW+kE6p8Hj/3e
CekNegY2BX8yIDCwcLx7ou9BQlLnzZTAklRm7cODkTYs6ENb/tIzDkbosXnNhxjTGLNhB8LZo558
MCRGjrFvu1vad2qz6Nuf2c2ytnaVJ4mihWd4EpBzcGjkt/y2KdyJ/w/LTPJX+UUWsuEkDomAHkoh
pBX3h3tewbpz+buHDneZINALLuyZlY0eAPE6vSQnHEdLMhEH39IBWbC0R2TBPXITz4mrFQ6hYes3
Ef2/eaAI+yLuiGvDKtVHRMjC820Ux5056AloQFkgET/DtXUrTaRWtYjVWmyJixermIeYbkyKwCJX
EGjIwd8YJi2wnnRiV8wse6ULd9clWFRYROUnTPQFc6922KBL79spTmFQs7O0rNDwva+j/sd6GsGE
Wts8Gyqyz1IzbL3q1GIAGyLLtH2nmf5OWsmrGNuYJ5BCcdQmDxm7C1DA4MelmS3t7z3PF6NTQgUC
Cr7v/4iVwAki2mt0g2hWi2AsVDtEf6RpcixUtg9zFTHfYfWowYIKN52gNsF6KLk/DIRfzgUGv7bW
0BQej41BKLEQC+YW28u3XGvnw5/13Dtet1iI6yUHqC3gha3uybjwIoMRDki6vBsPys440xPdomtB
aFSdJbwz3lWOvIsNzns0X5bG8QOGoJq7oNmfqLwxKpGZCvusZKth263pmtWZxJdotDZU9PfX2Jh4
yJECQJVQ+xNUch5U1PiCnUcb//T5aa1G2vjNZiiUi8x+yPgu730BcTPlnbUTzGhlphRk1vqaxbTF
zUCnrU8sbRWpfjA3fi0ShpKesAlzT5n9Pn9NjycJTYHinMy7F8y9eCLKdlnlC16OZlaNkGgyoHBu
bMzGMPoORt7BOyJ0oa+cTZiIniXHiE3rknJLy3JdF6Z4VWp0tcoJQQ5ix+mXFh9m57o2TRFMnd6i
uQTnfkpRgcWDm+hXsh+AgEB30CDhlNkTmRrDYTMrGNKb0zSSE6w4gk1lfC5Q4SbT3WLmtqR1P1qs
gvAAxP7uKZ4lna+K7XCzkp7NAz+7iA7bjsVZmMkO3PVCOS04lkU8tnmM6QQLZ9y2qipydDLe9KyS
2t7e7R7K6VY8WPdKmRYaIKejD9U8NAcVRo77vQH1jQ+FVptcu3S38RZBemkTk8IUKnwSBFvgijZL
9mNGajKO/qQ480GLaltH4FJ1MeL6dfg9mJriVTe1XlE7HaGuhuGSrIpxjrcfbimT4FL3DpMWsp1k
VirBeQBj9GXhX9DtC7v5JD94u/9Wl3/WSByr0i8Sfe5IdPCNu1dO27OtFaBunzmr1c3TNiYHOPY/
BitDvxZM9w5CHkGYc++RdH8bgpA4pY7TChlWSYKv1UsDP/bb6znvwxaNM5PxEdFL3lDzwM8Sa2rf
1aMNurKXDPn4S2rjqld4Pr8zCXjcnLePxNCJYOhJgbbWDozOz5aNUK64AUcXY0wMUtHnVQOtO59l
8BYxOJtDog56Rtaa9rMPehV1kgCH9+LoaOemiC8Ksjo9/j/4e/ycryahEFwwYjaFD7cK8FXgmZ07
FyLVDgfc1wPu1+1ydwaz47C8Eo7Tf+C+iwHyLO1efw538J+Q3IxRpHOLZJFMZwRfpDG0bgKChIbd
H1SREQXrl7ehufioU/+AUds88ueS/ng7SAYjtJVJ+rNhCrVd4QcUA+2YkYrwnJfuq2WzLoh/9a91
2UVDWhTz/K1QEtoaxg2Dj9RidCgmbW20LQSVcZNqFqShvTXQUHjhGv0Spiaw9cDosXwrCfn62K79
Ikx9txC6xPnNcfhNbofTwRgh+rQVG6YsN3QY0cREhHzS5xOvqn38pAE7Xhvrhy2Jk6xhOh9jnwpI
zLgvaHnK7IK+Tyc9Gzs9XLIu825vE/rqYClbIZYANtn0Sst+883POJtfqjt9M/HzcNeEw/JeVJqV
oqcJ/N0Io2O0cD+RuNlr/lmSVBWTloOsOddVpOmDH3P1CAS3sFA4sHrO1/6DZY05ZirGshvyxIup
7pePP//unwF7tTISxGzu1kECY2ZczIpJdrStfcoTA6rfOTph1JTXI8rxQdWcsZQP/qCu9QXGR0tI
/oqUfnyLW6dyAnnSDoOKUnBPtfLc7GsxdPKRxdEJPdnA0IheJbwLwg6rqUI9egOSL72Q51TfwkIZ
7SurvVFwq47fMSNgRCUw5ojoydHtOVuoRQDDTeF9Vj9+6wqkTYd1h+71/uBsbi5behI5m3ePgY6m
ErqTyfnyzIGA8XavYm/0716tab28NxJAPCISXfil5IBs9xixdwQMfmrgPcXGzlojgY3KptDg/tnJ
ehV5GdQhU8Tg0ojuiNjiS4maIubajJIol16nCvhGUEHZeAlot0RpnzqjamSaIJRcOyXydlh6JH3f
Wc5g6dpYRq4w25XHGgY9TPz0S7uj71GiPrTA1JHeu5j75p/L52WheIAW9lBcWuSTcmLri+Am4YBc
wiUD3jKemq/uVswcH5exRnx4R7F5jDhIo6DcpomEAe7v9360gfBKJlUYwD16W7MGhKZ8VsF0E5Qs
rykusmr/cEylO12T/ZTJYNABhM/u8XLlCRK7cIIjALChE6s7O3X5oKmOFpLNpAN2DLfbcZaNDV+X
qPQBx+FFBy91NPoU9oq+0EsefuGrh8HccUOwTaAZdvjzBRd/gA1J89wgGKbLAOJB1N5od8RoWoUB
smz2zstEADJiNkDURDlG0fFtBMY6pu+eMhqSZOrUvhg5IWHdZDfFRF33LVtVUO+pzJG9tHQmfHT2
VYxxMrtk7/mz255h/Gn283bXjPNNZjfYuRbSoiYlOsbSxh2tZ9xpkNxdjAUHE4Z+l5fhw7RfPfHv
1HOUXtHxBdVXC9DtmXQqs1uiYVzncN+T3FCbtEVDJG35bJhfVlqh+l4kI5qtm4JsrvBmsP4Oaw+A
+Q+bT7sh53uxG2RX13qucuQt+G5bTCINW6eNuMtWn/1At0t5BPnVfIufWeciko4KxP8j7z6CWKGr
cS3PO3Y9oWOqy4VSHXEAtsrh/SSk5mlSJ5bDzUtF8oUjmxQQU31qqxWve3DaJnH6Syxy/DWLh5rD
A0jcdakDsb4y/EZGUaU1A3O1DKbfuhacLpyCGRjGPB+7nFnPrCX45TMAvcrjshsPPMDf83c2l8+X
6mkO6F2A7GE+p0eZdhUkIg6+m460Ol74+XgW1GHsAyz+FX3x3emxzYqovzpTvwJWclPH7deBHwHZ
AORMzeNm2arrTWzNSiAQZT7rMrp3shKZyq6gI3GTK7g+Ag+NiRvcuh4VuXih4FOGtp+WEh0W7gUN
c34PSBvLxcImOcOJ9wnMgHi993NyxJh0IVzqhXXr5V1bHf4envITqfCI8R3rBrndRAt3WIPNzm1B
IhOpsZRbiReuasonDbT4LrwdvaUM+YVj8fMrCI0by99Ix7z0sI9XZHROeF4RWtrxiogI3fXP2Bia
j9Gkw1XlI+zdQkcOxM7nlCBtxSM8pKRBPk82mmtmEiQEKCL63+CoL4YdcCzV9KaLCelWKY80F8iJ
IAeuRhjl61FXEiHCgby4WzO3wGdmWi593f1sBqsi0aKapWcMtKasjAfxYpn6Zxzu8EA+wH6LTJsM
f9A40jHCc3NPg5XtG70UrJMfTw1lQVfABz4qS8EU9a1QJQer81SqiM0qCkkdX9SxW/L1oLmI060p
SylDZ3RwRGUSltbMz/tLlwbIUVHCRmX7oGBJ7Qviak26fWimLr2Ve9ZXyNlCYuxe+M4ifdg+EwUB
+zmBqnbXw1yH5/9Jm9lKIK3KbvivfRg/jlvOQuwYLwXIVXwGTMNTBBFUv8Rk5t62OvzCP+o5j1Dl
UIWKirDtcJuEOUbFt1Wjqa9rZWIcyHuLZvJjq2Pgea1B2TMZHoWKEhDj9Mi/3TJQ3OeYFQ4//MSC
VnXDqU4BtIIFqJy2qiXSrrP2AfuNVlvY3oa6khIzQvIkupbdsMLJdG9z4q0wKJKbJDGao3x9EmpZ
fw0idRHcrNClgtt/TJJsG1KF6LEWU7pk70Bbh9Hv1qTCPHTaPy2yb6SPmLzBRPeZeTgAOAe2+4EC
HXX2roTYyrLG+Sac+b9G831ewsGyoEOfWdViYO0NHvfp/LG84xC/x6PWh81AZkQ/
`protect end_protected
