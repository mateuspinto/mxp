��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���� vU����U�a
��0�j%�+1�X�aJ�t���W
���{�+���&��o�P������ԡo	r�.m��^z�w1q�K2NS�/uVz��.j�7��S"74,:�+��G�nc����O��9����?�����o��\[ۚS;.�4�L��q��%��g��z�v攌��8�F��L�Mx}�㴭.���h��qH��sl���k�-�f���?S~ؐ��SP�L�/hՇ���*�/ЦdY��4R�i�/ImY�ھX�0��˼�o�HD|��#H�=���� �;S-�3� ێ�ȏZO���}��j��;&��t�w#�e��_���țh]��1E���f��Ss������	:斶[fhM�	 �.O���de^����Ƌ�8"�`n�K,�(H�ʨ�ғUZ}��`��!��]�i"�U֦��=,5�'S��-�Kd�N�mV�������_��&(���� �L��eVYom��U0ɺZ!�(�m0ŗ���}�1�)�#����96�vg>[�ܻr�%BE.�kFE	5�^�b���q�?^�		j?n*\'�dP�4�|4:Ì��B+T&��jv�W�I��l&��|�d���L���c⼘��F�=�C$�'���Z7���C����lp̊/�8�G9�F�Iݨs���x�X�sm�2�TӍ�p:tb�yZB:�	��A��ܒ����2IZԷ,i����Z�$��]ow=�C������/� L����K�� ��R���� :�E@u�����7B�&?��OwB�u;�(�09�T��{L�q�}���3R���G��h.��j������Q�v�����LN�P�����T\<��w�XΘ�Nc���c�愧��OQ��C!�ͦ`������ր"�w��5���Ӧ�y����NDQf��rdB[�%��<I�o���׬0��+��ar��xx�ms����.��/U���������R��-��x6T�SR12Ob����¼'���<@����	\l���Mh�:Ceo���r����M�`�Ш5��ݰ:�c����FyU\���{�@7b^{���Vm�H��%\�z���E*�R�x�b��F/��g#7N��?e�i:`;�$��:������O�f\�K��Pz�cf!���@�s��\��h
6�����Y�ӿ;M`��O8�z{:l_Lxx Al��M5�����V�h�k4�oXX�����z�/�;�i5����7���V�w㌄YS���pN��O����30���6�e~�	��k��X��g�~uw��������ɿ1���֖�)�  ��|T�	����ߦ&�~:8�1�n
e+��ۨ��UMZ��aa�>��#�Ȳ>>{֙c���^��Y])���N�Yfh����k�0K���_��3���h�A%a	��+�'0Ta@�a�$?'����n�A�	;[�}�ȹ' �� ��@Y")ݖ7����v�����r��#�fCu� �?�ՈFՆ2��x���_@~��1͸D��&��6�����i�u����psN[BR&�d��ԆU�
�^BG�<;�b�5�����K[�
�k��z�r����?kh�/5�������N=���L�ߒ���H tp�ȷ6&2C�c�ˌ��;KVމ�U���Њ�ُ�����ډ�����Շ3��X���E�Z �YOV��+>(Į�
�=��Q���2�ƞ�{I�@'���VA(�Y�!D�T2�J����b���>��u&=�-����ڏ`���ݣ�@b/嚘�!�r��t���)�r-�ʪ}k�*%~������C���т�ۻ�~j��h�֕0�ݶ�ڲ�_���B�kw�Lܹq:���y��GR�A.���b��N��d�̘���	*;����0���a�u������y��^�`��Ʌ�� )�W�6=�]Ği�����m^���_�%M}�o�N��{x-5�lrh�>M�|aq��r�|�:�v��N����ч��c;c n=��� ��Kܤ#J��!��>!D=Xu*����ۮH�q�����i0ρ��br��4a��3JW�˦��B�����]�QIG�R|�A���N�4��z�����B��F����,�[E��X`J2�I�����aS�;vG�%*�T;�S�SA�W ʑF�U)+ڊ����)F���<qN��-�}�K���ӄ���B��&�G�G��c��Ӛ�v�G �Ў�A���i��ڡN��{�o�YU&s�	�NQ�����`���*Dv実aYz����U���� 5T�u��_岗L��p�>��ٍu�bc������T���K���#Tvu$Gx�1h1��WVq�"R-����v,]#e�)�S����;3�Ϋǯ�F��э��Tz���i����b���&	h��k ~<��%�0(n$v�׊	q%�����k%�{����]�ھ����̬��;F/"X%����ås;;��S�W��^��I���4SsCr
D�u@\?�M��u#p�	 �W�ڬ� �a~��ۅ��!)g  V��l�Q�zFG��I@������M¦.r����jWL�^"`��5�m	�ulY�~�e�縨Z.�Z���t)�^����ڌTv�և������
ʔߗx�������䴑�|�J��8��P�	��C5%?%�~̖�<�ܪ�҅گ�lV��b���ھi��B菁*�a\��̿x� �^�����H�~o
��`<ݰ>z\~KË���������4�
��`�B+������ \���7{�O�B�r��JG���1حnɯC+}�����w���=<y�-��V>��u�=�Ɉ]Z�<�Z�c(rF�5�^��8�v��;�����G\=�$��E �G6����;19a�K�B/����>K�P)jT�(f5ˤ��16�����$�<�ɡ���/��� ����(�����$�!����x�f%�\,�M8qLj���b[�{�(�	��G��y�\����ԦBN>��(�x���y��\��b�3./�fg����. ��t�-�4���HX��qnF���Fi��-�T��k�f0m���ְH�=��_d
'���5Jl$� w�׷�m�@U���,{}��ϑB���Ad2�Wd��q���NF��ą/����BnD�a��{���O����
�*p�!��O��}|����*<�%d[���0ӝ1;J(�Sx����Nc��{��/���!�?8��ϠL�س2�о�8�2��g x�g��d�,��{�O2zfR#/ىM��9[��;���+�z�ȧ��M.�����ɕ�I�f�2A���f���ko�YB;������k��-��?+5t5���E�@cֱ㫏�"��K��
�,�>�S���Y}�5!ض�w���g� z�e�Q�������=^��bz�5ט��J`��(�|�Pe�눺x]#S_3M5���	���c�S<�Ј?�Q*�
ߋޅ)�G6.F��x#���3�hn�o�.�g/��[d�Ùq5�k��`�B�Їa�z�(�܅�% ,�M�5�R�z�#�q;y��r�}����GƍF�ϱ��HE�G���q����Z~��Ԃ�g t�Y4-�UKA׌1��`eG�U�%"��V��6g�����'�m��)=v�ң�����>_�k���u���� Ց��-� Yҩ�Cl3$F;Y5��0À�<�}j��)�E_�۬cY�Eb�������y	�d$d那Uͥ��'k�`9������ȸ��1Ѽ*�m!M�&��7��#��TF���Q���D�~S6gn󯜛���#���I�;^�w@g}ϝ� �l 
�� R�|<�ԟ� T��kZ�57n�<|x-�����@4{��C�u��?:yl��^E����Y�G�p5�|�gM1j�-�wnq���V�U�;��?�U4#E}���Z�`w���yS�J�׻����M���~�x#`k*lq����?��.b9����i����'~4��W>9��*AФ?Ae4X2Qu,�pA�D�O'^fY�iت��lP�і�Q�5�1�h%6���@��c&�CFr�b�.U.�K�����.���-uy��*5�f�����D�����9�(y�C�SY��z[�~��M��abb�.���3K�n@���N�0�����|-�">������Y�dV�
��ޣZ|�h"�	g�.%���JG0��|g�o}�/��+c`�ޡs!?�A�|�@�K����g���A�٩�(�fؾ������uCGn��@����Pg�H8>���Q�t;v/��b.�X�����ȸ����¨1R6��{Z�S�#�$� 9���zT��_��|��Z���G�V��#�3��&����OD0O>׳����ƽ�R�*���:�I�Xa���Ic�x	l`�Ub]�Lwa*iido�Ai����i�-���lQVȪ�+��F� b��*�Q�/�Q��� �}g��5k�{�35���n�v�qs�r�+-�|W2�)��1�x&����hQ��
д�Ӂ�Cv���L�=" �VH�xU(�L�1�#c����g�c�L��P�e���uu���Ni1� �U�n3j�W��S����jX`��Y��z��ƹD�Kq��#e͍$�wYS�4~3+�3��{��Ix�R�j����6��&bHHM�8Le0-��[|djZ�a��G�9E�ϑ����X2'��Ik��y����5燵��w�^�&���"��5�NGs!���C�3�"��7���޿�-�gW��`Yhwa	_D'z���vJ�ߎ���]� �zO����]F�3��x��U�b�7R�Z~���g���#R�p����hUڭ}���WG�D��)uZ�$ʈ]����OY�bC#r�����|*���[.�>5���f��X�1	d�;'��<$��U>���.>dʒ�w�>��7�U�U���Gc��Ȇ�~DF>r5.��fؖ� ��5y�~�A����G=�&��8��ge��v���P�ڥw�6�k�������	��%��8�!M��3	ɕ����Q��6�P��B'��5��W2����|2���n,�c����M�\��;"c��*_�'N'f�nt��<^.vƀe���@���#����!����R$y�l�j2D�t"���49��w��_@+9|�;�u�7(P3�M���E�7-����K�1�VSJO�2��N���é��_y���gdVf7��?�BP%o�����aQ�?3�E�e����9cW�4�fc���wCr�4y~� a�T��i�9�m�ÇN�*Ry4~���f�
Q	ޠ�Нɗ}␎����o���Yfx]4���a�%���Rэ3Wb��Sw^:VC5��u�u R��m�����+јق�����ⷖ��Y��k����/z^P{�r���}_�b���q�OPv�W]^
�l�����ZC���Jj��ʭ��kx]��st��;
�lX���F���w�TJ�ȓV�RwF{G��)bu�|`��M��վ"�_6�����X	�5@�6`!��!ѻ!apk�za	�Z���.��m�=0;�<�-4U��,4)�����>�ag�;Ŕ�F�ٙ~�lt��b�aʬr�@;>�M��PO$?�L�9B8Z@���ݻ��s�;U^�H��6@v���> >c�O�B�&�֣���N���i��|��?��FY6�����JO�~R2+��U��	bSԸNqhA?��u��ޝ-�`tmIP��&w6��H��@M�H����H��u�A�1N��p�4�d�������N �a;1;o�ͮ�|K��b�'�P�����<�u��mB*>��l��\���
����[e�uA�����rp�v0�HA���,�{�A�`���/j�%�.S,Qs���)j*�ʲ��C�G3'�5�c#id�H�ueZ�
�^|)�F�����R�¯�Կy�țsܹ ��c�u5�P8&� }7��+8ސ�t�(`l	��+!L(�7��Pn�mhV�~��&(�螨�kF�,ON+ȅ�'T���K�f�f��c6�͠1����5���>�ݻ�H=�+u�G��mע1�vas>)�B)��_���������5��^�	���t�m�f�iN��ׯ�Zu@2�>ӍX�O����J�@b>�� �RcC�.<��n�I�Kͅ�~�˛�<ro?��\ PЛ��3c~3�*���*�1S��Lx��!�:��aJ��#[�����&��h�G�͒_E�*���!� ��hL&�rj�B3E^
X
��� Y���	�� �@�V)Ds�\5�޳ioK�<�s�0V�����W��v�U�k'�t���d�
Q��þsM�� �{M��o�����.�i��6����C[����p��X���Z���q:�!���>��ġu�Q�1��Q �m)9z��3&�0�0��ueU�l���J��_��W+�Ml�V���Y���-c]����d��_�A,��<*����&X�Z�\�̳W>v m��W�Ê�d�:{���a"�&*�y�$ �]��j�q�Npi�����S?���q�
�&����!�L�H&~d���Bɕ�q�|[�5�-����q(p��,К$ WVa/S�q:���ݝ�%���[^�O�֪�0\v��]fM�6�v_ZZG\��;iB��u���=��7q���l�ٿ��j ׿{��?1��2���RS��|�������EFӅ���_ڝ��V�c����S����'�;~˖�W���P���7r]�~�$�k鸊�_$h�L����R�)��_�3�l�jG���<��I3�	�G�T�c������:������� y����{��LT%��!����i���	���- 7�|cMW%R7:�">�υ,e9�+'�e���#�d���X!�z������q��C��%�РY�x:�� S����VQf��?*���x�L��i�_�aw�;������@��P\t����J|6���L���vI5���4�A����4�yӣN2��f 0%�j�Uw��������zuƐqJ{s^���ӯ$�"��V캚uy,mҸ;�;��)S�!�e��Jߌ��u�3�E�l�ԻB����֮Wjb��]ɕ퐝�<����&@̯��s^L����	�}�k9��~%��y(I槦���'G$'\�S�.�"�Ӛ�m���Y2��|��C���GytA�5��4Ú q���A`����%���d���MSS�����a!��5i�6H	|mI�5x���CQYj%4^��}]��'3M����=xKLm�,�V̆Iǟ�(�(�,�O�ݤr�.���{j�+�t�	f�yʹ�p�k�.���pmR��Bh�8��-ZxnZ������3p�)-чv!T-��]!s9�R�ˮW�+�g¾�Խ�t0��((mg���/�ih�/�*�lf?[,�jyv�)C0gy;�O���l����B6�{b�w����3ò�:�5��������qD`��T;h���{ۇ1B�?����#����������5/�0�A|��m^��lh��܊���.�U�fܭ�a"��^N��8[ Lu"�y:�j��!T ᗨVQ7'����f��^��V����5^�6gI�O{&��sm|6�@/�7�0�ba�2 N�4ΐY2��M��
��=	8��қ�V�~n�f6�cy������8�c�1L�C��z��ɺnO�q�ɱ~`ˁ*Jwk��GXg�i|��������9�J���+y�����[;}��Ћ�����O�ǌ�2\
?��b)�Y���=C���t�W�zxm'����=ؘ'�sӎ�Ŝ�����tk���-��ȁ>�Ǉ5�<�"���ˠt��!6

�d,<�Y��m����|)��J����˰g/ވ=�ʉ��b�?@w\���$�_��)?�\/G,B^5
�@�������.�-���L��	�i�������Qg��7tqR+�W�D[l�(3~5�RSZ❎�h�������t� 7-p����Ʃ�����I0O
��*�l��EϐP]\̢;���.�wD,_�B��'�1/�d���P�Y��p?�ϋX�������Θ���������H���$�EK����j��;e:<60s��TbF��������� v��S^�}(�h�6��݂�t��?߂x�C?��%�٩��J����~���l����9���+?˛�,i�D�R���[���e5'���Ы�����?[p�}���DXE�S@��QD����/p	��"k:vO���@��~�O��J��b���w�D�8���M�=�1k*s�8F�K+W]ء�72t�nO�����\rg���^���@lp���n�2 O_ ����|�OA�E�j�B�?���q�)r4�l�=�f����*^o��.[�&X�đ'\9�92+���7kvW{�I�fVQΑ������3����}!0L]c�5����R�ɽđ���xP\�뇫�t�c-w�D������0�wh�?��Q�'�u�J��h\ר��V>C:Pq�m*y,����V��=qx��R�D"���(�� d>U%
�v�I[���|��:��,ɧ���=7����C����H��սp����S�X�I��>�ȁȕ2X���M�}^YG��rA��xC��HX�����V(�ӷD�D�E��r�C�K����MTv��e���	{��n�C�V[{��m �F����-���,��Җ�0H��֢�B�2�vi�9֣��R��?��,CO�4E���>U�u9;>�9+�v�.���5P�W�!�射��Z8��]�w�ώm���w}���w�M�A�8EJ_�����h�b��x�1�-�Y9�gc3�$ov��w�&l��	ݔ��q&b��F�U��'2��F���W��_�'N%RF�>C��� �.݆���\dұa(:V��c=vᓩl[5�Z+�$h���X�ŀ%��`���؁�Ɵ���������/V�׉����
�u b��ۉ����{!c�!����F3�L�qM����#��p���^�	���&��[2�T+-:Q�s٥/����y�;�a�N2"��,6BJ���DC�&���M:HM��88��Îe:�O�؃�Y�$P��;^�H�����~eL�
�Q޸4@��bV̒�-l��G�FM<sHx�E�Mʩ�e���(K��2�pf�Tvɱ?�9.�x����Nݿ-_-L=�燹�#�tSK��(��k`R�&�H��KJK�2zp��7��3��Ay�9��Cm�_����P�����=�pt���џ��N��4�{�,�N��t/G��;ܙ>y�#B�_�Sal>��@�7�վgv�x,kZ���D���D�T�E.���(�����#A;�w�0dX�`�rV1Ti�JX�MtƪE�	խ���5rF�T�ˤ6�kc˟9z�<C�L���� >�[KbR�^�-�]v�D���7�Z�{�o[%l���>�MZL���%�ዽ"Q���Hhz��:�!\� ��hŝ�u�)c,w>]�	{^��Z���:��I�������i�X�ⷾy��q���D�?L���h|D�tF����)����v�K]����n�'�pOuP,�r�Ls���ϪwF�n������3R�pz�Du3�O5��ݵ��~�"s����i�v�Pt�C4�t��+M�:�b�`�D�WH��(0)��L���lw�ũ̻]�O�J�_���	�!��X˧�8��b!�XF���)��ï�f�����}4Ń�W��/^-w���#��2$�}UuY�@!�7Ϩz�L�_�˝��g�c����:�M&�1�
��v�DRS��$&�_,?�����6���5��=�!�h�ƌ�X�Ge<���@?���OΤ�l�}ȃ�#��}L꽶�$R�m"�Ï���p��zcI����?�	c���b�N=�ET�(��8���6���k��\q����>���Y�)��`�@ -ǂb��Y�p:���ĕ�HIE��²?C�4�Nbǹ��#	j��	���|N�p�͕�(��5�ڒX�fxz\%���(^*����ݧ�R�č�͉����	ρ ���$��}FJ ��&�e���Z��oz���9L�Xo�j�d�<��.B��N\���,�&L����o���'$Ͻz$:�����4��ք� ���p�)W#Z���P}����=d��I����@��]ɇ�T9�+BJ�0��KoI[�|I`^)p�1��{p���\˕B�����J�>�N��\i!��ʥ��33��(W8�Y|����k8׊�O@�!~ 	#H�{t��X��0ŉI�i��tl�kC�$0���o<���~Q�h6Dr�Uoe�p��k�;��_���Dd|��l�`?�.mp���J��b� ���E�bĘZY&�)��W���(5�8F�ʍ�U�}j��G7mmI���rbN���������F�R�!����uSvs�u�W:3ȏ,z�/(b$�"��0- Bp�^8���3I�����5��7����=gA�eHYܒ�*&���c,[���0Ӯ����+�i3�xv�'o�R�%~K���D�<F�It�w@E�0�Pgk����GW㢉k����%�_�OȐ�.�#��d�n�����=M ^s{����Q;�,BU!u�Z�6�6��B�)Tc���Y�;����L��+�$b�7k�	��3�'�����@b�9��:Ъ����?�9��:�{���ʏթ��V,���9Ek�㐔'aQEP�~�kT�,�"j���,����#ю���}��)�zR��F��spN�z:�Qc��x�PeqH_[��A&w#�9-{LNR��^L��p�8e�-Zf=>�v���oQ��VN$x���eY\
�������@�h�g��� �"�k%f� q��vR�Ӑq�vT� ���s�JF��yK�z!��vȊ�\�V��$���}2 0/�j"p��؞]u��L��bo)r�<4p��Z�׋�gb�Q�6����j�p����fM��5��Q��1�ẘٟ7�Mp�Cs,�k�%���Fklf z��Yl���h�X�OW򳳺�|(��n������2�ɊW��W*��RI�#!�v|ozo�Q����5\T�N4`��ޮ�'�0��~�}=rp�s����qv*��4p�i���3�#�cPԳ�u�hxEARct-�@���; ,>au⟴ےM�t=_�p\�O ������B������z5 ��L�.3��������r�*�=�M�#��^���2�Y!����2��Z[
����o9t[�'�[;n0���v��S�W;$�B�j���d3H�d¶�v��͊�=2=��o3�k$N�"T�7��H�H1�x��|�\��ed�ڨZ�7!�x
U�0�h<>��`k�q8v����KdQ4X��+�JV�Բ�����y!�f��}_��?��RBK��Q���Ԧ9yŬ��R$�	a�r�@��|"!��ȋ�eo:�XNR!%�f[�"�ӊ`Z�N����R��"Ȩ1�]G�
�U7LYd��rKp�0��G,3���r:����Xګn��v2�����/�\���A6���g�۴K� �O��R<������.£��1�C2�@x&�Я��1�M�]a�XT	]��Q74`�������N)�_ P�1�O||��(���0sH���FW���e��)�S(�b؋�/OZ���Ϛ~���R�Q��0��q�����&ضuQe�®���j)�Z�
��k��l'�>iɭt�q,��Op(}�4L�C���D�Y�66H��hj�6a�ܧ�������}✉\٠�#�+� �����l����CnaWyq��?[o4%C��?-���`�?z�W���T	����t,'���x��q<%�y�r�8҅��@i�����Ȫ���vɧ�py�g4=��h
"R�������3vSR/����P��@X7�m�Rd���5�/�PqoW_�2�* �((���kո�A�̽�I��PaJ��6A�ܤ�5�h.1�{!���������=1I�VJ� �ٽ�赹-�R�_���)q㤨G�7�RZ/�7�.��0Hcn����P�e�>�/���p��ɤ�q��)���;|�1$�]=���K,� �OJ/8���G��e�?�\蝇FPz���R4����(�$D�%���fD�m|�y@8EҩA�y=�!ic��$X<ڐq<8�@c6N��9��X\R�a��
�o&y8�w�v�>��C^����o���vs�x�ǔ9O	G����bk�OMH����l�G�	8d{�"�o
�w��'b�͹����A���z����v�J4Y�Jcd�4�9҃���'�s�s�<oq����}�J�ޝl�����-VZo��U�}xVp�	#Kf��
��|�����B�e�F=�h"��F�]������_:=��m�kS�(x�5cH��K�?<h|/Z@�[���B�Y���kc�����0a��8ZFXW�egܮFC��C#J��멼
L'�Ya��Ͽ0�R½��C�@OPyB*�ωq3~�a�Y����	UCobX7wU0�蚦�@���=,�3{"�%}24��.��i��+{��c.՘��Ȟ�j�ay|}���C+ ������	{B�Jjw�(x�0臎6�&E�>�W�3��O������z�ҏb<������~ O ?��0��(�y��l��,��G�u��z�7�*���Я��y�����5���6{�?1|��"���=S��r�Y�-Ę)!(r��J��ERf_��W�Y�o[hQރ�
��(�����piBPN��O���j!���;�uȢ,>��c~ӣߺ�"
�� oibJ�A�Ph�QsYo!�S�w��%�q*��?as�����vX��C$1@��kU�Ȏ<�V�F�\�T2���&��}j0�4�	���襻=�	O��&�7��������l�x�����.\�ȣ<�!T�Bo��=�}��$����j��nS[Ãf�1�ԣ�}�u�������>���  ��E,H�V�3W[�	������L<��^�,��[���� ��[L�������,�`9����_�������N�V H�x�};}�F���Ò�D��\g�\����F��
���ĻU���G��e�1I�I�q3D������+@o�O���?{υ��sN~gg�m���>����w�q8�R�/2x<����羚c�E;Ώ�6T��¦p9��W�ZbMƆ�8tkB��`ܧ�G���`~LJ#k���9������R�}��;��!'L>���	b�x�������6�҂*����Z҄������ݳ�x�#q\SJX���җ�_q���om�j��T���<�]��J��T�\�F�:fǿ�2����6ھ)�M1�O��e:]pSL�ޘ����J�mџf�\����Mը����}�[:@ F�p+����$<O���E��B06щ���}�_4��HU��m��i>�~�_�P)���9J��R���9�1�߬�����/��o�|��*p����N��0c��Zľ���:���2�"W�"j��L��ڕ��ryp������!ԗ|fM2	�2����"8V���Cv�eԽ>��O�]�*��ϢVk)��q�1A��oP0��!EhT��ݨ�1E�hG��'Q0�*W�5	�<ʻ�?�'�y�`90o�8��d�W��Y5i����NtK�G<$v��$$B������u ��U����a�bɓs���k�W���fY;2�3�G���v���_�t����G��MɄ����̙j�e2���L�۵82M�į�	�mjm��-�{1��pgZZ-Z���B��-� O�jsk10�Ed�[����{�og)��#�G%��8�*el��de~�-���p"7v�N~H�	���ҟz� ����`�J+Z�u$)��T͢ja���d_L�DToa,�_�� �r�(ߍZ�7�~F��.
z�ݙ���Q���0��Մ������&0�*�U�߉�x��D82�.��ڂ&y[8�k*c�ˋ����J��_)�i'�]	i�a��F�4�`q�ͽ?W�_��s�Yx��Y�S�8W(�	&_B���LI�WZ͉W�e�<�їR8�X��`U���c9l��~�\^|� Ѣ�& c����e�>lq|r���isq���Ke� !�&����~���c��y"l�o��mZaJl���,"�`ң��F�[���EJ���)�`��M��O�v�!���b�����K�d�x���v