`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`protect data_block
DH70PQxgeeL8JVJAn2qLw8QAz4kZ9uG9/NGhcOP37+zU59Ir3Mdq+u8u9DTWeYUEKAKu/my7L2w6
GyTZZtSidjixqRvNuSOL/zxL5teUE65ma0p0dyl+78HaIAh9j+MnNXHD7PGWwCVia644YUH+vkT+
KnbuZ0q2vD7TkCAJnowZ9RIe7Cdqe/Lyi/q44gx1ejsVHaEX4C3n4/LZGVfHx/u+k4H9tN6q+Nwh
BL1Z53cepXDpkQfOxGX+UZkGxGeRzrx0LyqRkHD/Lk2fOvLjs/dzwC/piAIcT5dS2ppAQsMmR5Hm
t2NNEBISNb+EkL+8uQhyGrH3c0DewRkVPETBZJ+LDwNjZ7o2hEmScOHLP/TJVkgH8Ln39540g3SV
1iq/fJCzHzB3qZAjFQFxGNFqDL6qjKBkhIQh2q35PVz4ZOy1niyr4Jp/B9uxNtvrgjArV91dsFDi
9IOAeS+T52ExCnXUiD1pZB4U0qMPfQkOyIeXYhWzTMsyyQXIjpcUuV5SScymh8UNQ0dy2x7sg5jA
Z32ygqSWSlGqWZr7hct5ozeExIFC8K0Jpo2KFuwo1xS7hNvQ9tQr7sUR7w1UngdQ4z0eFI4vqy0Q
TRAWoTsGgJLelg9k0+WYD/b1cVjQ0KkYwShG0iZxrgo7/1TCRchLvI3LEJ2C+S8aPREZ/kTEA4CY
H0WKvhLq6dlWt3HJ2p1ejowEMq9LNm4RVxgoLumurIHJbyU7aI70IbYnAYd7ItsfkANecChWrFKL
Rpu12GFU16JVqCqctQhEtsSAjpuuuKxahaKvpHEFfDWEW9Dd2T4QLhsXeaSeplHMHhrpKNtVRDZU
Dmexgk5D4An0ANq1NKdjXtb7697ZtD8//4Wkvm8DKX9CpviniZ5SeEb3fEVAGX4sKmyiIps5DHST
to/SE2OeiLIea0zaCvARI1nn5+wOhuxT+u1jl0LugEX+JObtRpYqQ99sEi1FbXkwz6v18kjF3kM7
oqsNmiITrdHms2KvrqdxaMKN36KuHAo1aJDzNQk4cGWzL+N4aJ2H77/Bt6l3rN/37RQhs+dQjxoK
YSz2iz1T7PD/r42FLx/pz8kBPkwmocBUCG9fFcyZ2z+mnGyrN8CTP+bsrjluygCG+yBmgBqc4/KH
9H0R1BD/vh44z2S0/QIhtbGJqKsCaUjF8jXuC3Mx105mVjm7BmyngKuhgEIn2MDk9nMOH1UZ7mOo
hb0+BhUoXApUuLlFqIab9fGYylDPei3x3q5syMEJF9eOA2tuPqRhFR5qE3Lc85gkyPTiRyKtj4De
gap4Q7PmBX/QUXjB6CKUxw/w//QVt/jHmcwgFO587C7foYG5dpGm3RtgpxLx699lTCKxXwDWsQCU
f6t7Wl1IoVsC8qSKhtUM8ltdTam0I2VER/c1mziXeuF6H17atQKwYdUqgr3kk0fW9LrsTBCl8BOI
bf5ZUgOZSAch++y0EqItAx8zbUyAt40Y0JG9Li3FT1y7Dn3NzQLYwnUYCbNE/LlC8tQc1RwYeZ2u
8X7eKx38GYG9M204KptQZFBQDrg0UYrn3Cc8fMJ1oOVqWbMEzE1U+CglHayRIrhUCAjDPZXw+EUO
HEbO+9k1w5ODj57wn7fEkw0M2/L/bqJHN6okwY0C3iuvV4Pu/Cpx7HO2BIsDZKbXycw4kbysIxYW
ZeNcRkXJXfR6Wi+ULNaqpMB4bOTbqd1PSildqu22SqH159lui/DZlPSD6t+KdmpKtQNRvMqYoT6J
FtgwfSTPENhkpAKB1IfeiW2DfBdr9jHbw+QQo9QaoulRdUlYEg+Fmue5+MyvuxUjvNRW7VBQCODQ
bZM2Wr89MfLTGLOVDDJTydJzUKeb2kPjxIeJMAk7DOjGHbWiUdFZbR+aF666YPXB2g0QyJ4ezae+
cqLcZZDodfWQNu/Y0J4XMUVlleHzPqkcWG+blwTb/nN72Kad+i+HvvjD/wXSS7LZ6d0reLPqXoSp
JkZ6PxzB8C20RKTOmPameG8YIPyNy6oRL1VBZ/nvhlYIvL+jPkdWSOqnzImPkDYKzvRVuQICWQX7
jlvRN/1qVAkXA1qjyeaiwXcSn1xjgi1CY6rfvIDQ/c7PIcQrQHz5aip12I+Rlr2DT/hrVfxyPMv/
9KAcOAHRpucw4KZmkyhFj7psfYA7rxXRlKzTxo4hHdNmH1PIMOw4VX5kIGr5DP+xSwWf1CdBTyFv
000hnlfd04jMNqMOvNf4ETNg2GbaUo8qb2Ok3QjZhTDDhy5ithf4D1kDFI9Ar2MPoV4hT/QiCh1D
sJOx7JoN1n+0cCmzoPhKnK8THZl2NWmAnO/Fh0wj30PXfXESgw2eYBV4rtWerOjZm7860wo1RWY5
saUhU8JbuXuhJqV5jrZZI6aQleS0t11Tpshs3oyJXYNgledGLhllpKuDIpFBAntxRB/HXcVr1zO5
AxwcmIAWOU6zldNB5zq8a58XTQV2cLzbAi65v0iIahLvHpB8XuI5w6qXazmyktAXsjQNsmnKZ2Ux
RAuwxnCEI4afqM4cdPfiFWW5kEbxyMS3a8o88sQDn8Pje42MtlDIPyYqroJByDBB484UVxE556Tj
OZsNtMGIZtLqmZ309d4V3vlLn4ghT2ObQF068oX5eoemmCcA7EWKaplznx0qslpm4X7SGTGwRwj9
Mj31qWMt0qrzO9w6Kyq1eOpDdfLbt/LHWF608DLMqS3wmQx0S0sZfNtiUOH7hyMUaPEdtmDpeQJq
QAPyVTQM6cr3PjCD6J11mPlCRXCzONpHwIN5EWoZE8A61kPygfZkPJ6/dtrV22xfu+2zyVSVwXqB
CPaWFDLsMMsHAzjaJMUhkdlhRp3GuW3bIl7SAzfpftc1Odq8/w0Z2yQiiUUd0xzdvei1f7sTRs0A
zNWSfnN34pi0VHHvCQOd3zLU0fkf0EkeWArgjHeoFVyu46Pj0V5mReGylzAW6Rcorgjm/n9UQYM3
Z9xHbGsGCfqGzp8TSrXOsd9drVFXxLRcYBO06rApBGS6EfKyFSOVcpfhrp5CXcU6HrPhXVs4yddw
TRXmBKeI2P7hjTfNwHUvpmQ/NzybIoZRl50enOpmksOvIuqHTX5hWVMcMVd/i3SYHxKte/0kuR4E
HCshzXFxr5X1ddeYa3gYNnxwwNBRhC6Xg6NMVE7CmDXd4eyS461BBUpEEMb/3NpwsSISDfQeFzSN
TqqIKReTD/0qa6IqERC512yXcXVRQtM9JxfIvCYTFmQfYNK+FbT0S1f7hHGYhYEG5+vtNjYT9dlz
0Gy92cjCnsrZaPIcyQBRYbib1HIcffnV4IgFNmUNodh3fSRX7XSS9tTUkvi7a4FhNmmman9mOYI4
JoLmJaF8Dh0bi7IvFX3YohTnQodT5YacquBHC5KNk5RLLtvH8S8K00eIMv7D5O6c7oQB8thsRPLh
1rE1B7qNnC4ymKfPHwp5jj1nUbX20Rw1RsNt/mbCCKehGkqmNKYG2k2g21cWgDun6gVdXh2TGwG9
GvBw35v8V8BbXMW8vZWFrC5RFLDUjhyO1xmNMtvuow7C7qq4vfrit8ikYcWHNapzYQf3BTl1Y0to
dYJkkk9wMa2Z3V1RTOvce7vZo4MK4GZYkpGgXKpuJJF/mwxj7pCMdqxaq3Gk7KfzZ47RhdmUqlYL
ecbBIorjPVhCPiBfY/nP02XFzbuynuK3dilU7tWOCWz9eSpufg2ljWF9n9a6IW1jMbpRZke6mFre
hX1lz4zP8yToZaKsbTAotddnG8YycU/HbCoGnUCvjCMEM7mTOzUUMVzpnE2UV9QM1lPvR6ygntap
7NWGa38pf2xVgo2+yGlCqqkhTsFXBGfAYU9X7ZfCXPGegsILmMb8hOx1fEMPxbIRqTKNrJpEbUcU
DqScVTHVfwtz1JGsXqptJzVn/AzEKoxyYqgkfhZYH2+lB/s2Ve75dgDMv+LvDQoVc8/fSSt3OOf6
lXCUt8W398/O8SG4wY0fddGk2bsAV9dpfVFxJyFrJrxDCovisH4Xt8+blCcteaMBdIpNgd7G1DOu
KQ2hguTaXmacOQ2IHNiZz/rEpTUBugjPyOX/YF13mbu3irTbIPOguWFLyix/VH+d3UF4tJwKySNB
/9ehZgu3kMt7QgLUVR7g/7N7s5wULjS11Ujl9xj56DSggq49vP2+a6aMybkdbvZ5oZoHCYrC5Gc7
MGEuGhMlsD8ZarsNMTjNg1ot+qcm/hneOgreWVtP4kFUEmx+9jcLED+PLDZpKcdGpbERNLXaC7GN
sfInnD4c1O78WRsUkJEV8oCymaHxxijH9HnXf6DLujujvUB8N0UoKF6I378eImI+ECP/pTayCQN1
PNuAHp7Hs+EcklGdsVz/yCSEXEX+MB1Vx15SgXMy1p8PrOqLrrDkHUBVXnY3Z/viWzXvI3VaCMJk
AjaVpVcZdDpkF799UG2+fcz/X61S8KlfVQpkyHphUVq9u65bF9TV9WLeNyTPbyqviqDm1YlySTqZ
dAWEn8qP/aIF0Q4qzuo/jEaD8S1MnsqnRRiJ5T9ZqfbyNbOjaQdVIeJwNQIezbscnAHzMbwze+nP
+YXx98SVgtuR+XVkDbK7KyqtZo0ZHUv3Z5+ipMApq2eMqNiUs2XlZP5FrmA85m1qY4MHtN4PmJoR
e01FaiIy4IbllGgwGb2z2A/l07+0OLZ1+3pq
`protect end_protected
