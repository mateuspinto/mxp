`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
D0AZ2SqmzjYGgqmOgQF1WbB+V/8UhI5a4UB0a5aRYXJsSeSW2edaGzoKITWlPnVJKq/5VKVI62aa
VeIWKObxcjMtW+/tsM0ZoQu9O/eEmGG1syWoH8ep0xO+ntZHsGhSXOhmMsCU8Q8fhj5pViKz18i5
PHEnitMLn42CMdM3U52Q5eYDSKY3lPpAhLK9hkLBpJacEgUw3576uJp6CE7QxkYT6vJOAH5cnuzI
TR49UL0hfhUGBi1H4ZzM6xveQA0qE7k1VHIUmjM2vLYBHtJl7bk27w7R4twUkjQle+Dw4E8GJN5e
k56nLvhTt74PJ/mgpjxt2DpMzAXvv4woMN+Hkw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="+cHx6wfkA0S0qM1JVzVhQ/OcYD97c4z3MT1ynZfwJsw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2464)
`protect data_block
N32i+ZkmsEus6uDguHLQhqVQvbv/BuRqFXUSOHtboHZAMiLoP2qdKVdDHarNv0QgtNrgtSV8OBPY
l5VYA5+10X2E7VfRJFnRAF09KWREjQDah1ePBEW3w9RaIv01YpPjLEmb6q0qfWzD4kCUuKsV9BuQ
agweRWEOegYVD4peGHQk9NxJYkl7JXHBbYoJFjL/1tM+Y707DCAEE1Xg46pSiifWxpZtmK7OuQ68
EObGMvokCsOoBwJszlqzqy38khCbLPWyV7GiTxLmsnqp1jAs5Cn9G0cQ22fJMXrI0qTBflcVB/Dg
vogT7sfc1zJfbHEVsIBfykcDB+0esDLZFkwNviyz+uyAzegtPTrDo12c9cfExYnmyCuQ+9rf37zr
y/5tXUeHvIug3FLV0ERppay9g5EpRE4Q6eslJftIHQcc6G3sIT7g2BpMb8zT+Ym8d+89cI9Rtc3Z
sc3C04ZRWXrArB96LW8u4hmCqMg/3+CeDO3mBQPwSZbR819XlvmTtdr0jXLTMMoOf8P6UG8vPJvq
yND0TFEiad+h6qNePc+yKGyGGLZysGVk5iRjeL29r+1wv8ShNyvLYtUs4Q2Zw1t9qbO+J8VBGLwK
eMqZbjH7YOGz4vdyZ3p4G0+3oNxMHBIoeiGmIDeDRnKqVbPDWFC8OtImA9a5/pIQl8F5LTjT54nO
rYI1l/R4ija5mPec9rkx/cWvVPj64Zd3GUYgVrJ/yyflBey/ruXh7DMXQHlZhvU8bfHfWY4LOBuZ
+LcBddD/sqNMcivbu0Dy+jDNCCz+dlKp6o59hGyHuO0xXBLTkxYGQwdJxRJVTk/OsC3MkCyFH9UA
nxtUQC1b5GGQ3MYA7dJiti/0JuM/6QFXwr5oths4WfDFtCLAyfAzNa16O2ABcKRB1KDcPBPTIeLZ
J8xYPOG3WGVQnELVq6oddHv7TbfnDr0vdcclSKg/EE3pJpbcRazMxXIqwh1pEu3swes4G16fr+fc
nlA1bc6RZFAVzGlkg1YIgayGlnD+A7e7zdsEAYhgvw6QBXGDEa6M9qkeUdN3LTvozGLFOEL/QpfR
76umCxEHEnwt0GJgembrybDzDwyTFwNg5SzMFD2lIhRepOHkboZuHbKnvaQ6gu2kKaA3lTDLxKy1
4hsiBwWf/Qo34n3sM6kOI+26ciPLrytw8SBqrS/avHpiNqlOKWtPgYsUJOvu9bJnGle+L9xM2GCc
BJKb1Ua+StaLs2uMb3T9oYCfWfi/C5mc03ZSEF92vbMC9sMI1+W7mXwbaa96JVp6lemb/RpprKh1
4hzc0HOCl/wqDoN1GPmpUPyZVN/mhzRlStetKiSXk9ihdm37LH/reycLd+tH4j+U3FGs5j98vojk
DJ9Hb3ai9bl4mxXmtsWzoVSkq9cWwlUj36FU+i9Fn7vLIeH7u/Ami50Tt88YRx+MMiF6H6mPdI8i
UdfkQDUDgFDNCndLGGaIhqfr39voEDvhv+b73VKRqFoZaI0jOk0U0GSih3y883QVJw95XUVbYMrF
ypiMUNxp7NQ8FRJgDjmyT6v+WJxIBOORm9kLAk06pXcmLpNDW4CMp7tr63d5tSD5T/3dPnrwGWvg
OrRn5RD3cpHxv12ewWNBO5habW2FJi/hUoZxFyzoxhD2BSPI/X4qokzdI1WNRx8OiT2eKX+LOW3r
ze/eFyS5eeOXqOL2FwSTtRLvqck43lf8r9QfwQE8q4Xas19Fv21nZ2R19u9F7Vbu/HZAkvlzZ83K
3zi4nXkHJok9SjWIrzY2NUXM0j1JzJGmxtq0h03A9gPPuSYLHBS20mivrJBah2fi8ks2ikCBc2+A
G8rnbcawUw7pA9vPEp87ikULpKCm2chRYxLi8+n6YinJqTv0KkHDdJhoxzxVNrfKCj8xD5E3hgwJ
oipAR607mA1LFMsLNQxs+bij/qS6rdRoYQDCnWEN1S9AHADELwfNZmZiR+yRhkpXld7ETI5zxnlr
qBvmbqKlQmPG+Hr56iODjEBAAmJwW8jjuH5EV9RUeHoFsiETam79nIAKrKW/XzJyCF0jFIrqkJoY
gfzUXyNcBHeinZHI2sXMbX0/NRV88zvHgJuexQOYJflvXrJfE98AMtUueGQv/TRuMDnjDwEDv0rq
HEe15HLXiobS03r+71/tCY7niyFYgNcXEjl6ITf7/yHNsRQMWMxa7rxM9gpwivDFFpFVeH8OzG7d
m4IQMt/Iq2keGY/mlaeVclOUGcng0Yh9N+y4KJBOwOr/bNdMymDkMCyK59FVb6L08FLsJ8VGg0un
lCJUNm6x9sbiwflT+R0vUXl6a6M7rRbLCBFeyBmEL2C/u2brRChEAX14CVgAMlTkdlU8mND4EAQD
NsMGDuQwm98NvYEwfEmr05zmcRZ7aDFGISD6BN6Sxcg0NeKjFejxttJLIK7YhwtwLSnQhTEeQaqg
dD1xx7CFM5A0mdq2DghhZFf5vkzv9P/7TLMdD9n1SpznzZ1Fsc1hcJp4UNHufitUF5p9vp8x8Z76
KNS6r9yuD+63/xedVaKBeq3ZSPjYYmjZoXgF4erpfGA+seSkB8pOGM7fYVoFf1F+wHye5V4FNUDl
RDH9P1IjIiMyGleYNjCx9ywz7O6GUmPGud5y22pteYXHMXc+xLRAPylbyZO5NwzQ4vfy2r9702/D
O5xCn9eEMNyGP2POHEwlJi3cthH7TNDj7YE3SIx52bAv0gnA9aIUrnP/fJgx4tYD9Jxe+gSHdQ8q
Ez52I0Juzbwe1Ucn1EE5vQkVpaZX5SMGpmsu2SMwdHjOXyfwTbE6XP4AAFUvp4Jxh3F3LpRzhuY8
GIFLz0yCM0iWcrUQo4yGzj2ozMayTK8+8rSOZpgMZ15RFsWCaulIc8YwXaWdYzgEFu7zgNmxWcIs
dp21lHL9REHSN1QS4Fz6ua4gbFZyqObsC3NVvLhWU5raeunfUiogcPFMno0cgQSAIbfslxnsOfDB
Y4vc1Gkqm9P5bKI3ayHhVoVwmo6a2omw2bonP0e999I7assO4p5hptJpqqKGm+e2iHfgsPdfUiaQ
hU1M5oLCIe2Gzvi/A4eLUZanxCstRa7dCuv21qQh4iUg8rGY6FkFIgyahgbmNEF1moZAkPbsqD3Q
UKF/Yg2wmcuj3JD+4fTlqvdRUA1fdjC7pZzwJS+KQQRpsMW/p+SuuOMYlQlIr65H7G94U1Z8nNtg
ok9lETTPqVg6Zan0+ZkJ/Jk7rLugdbXFs+KHRNAPb3EI098DiCrwKdoiGYKhStio6tCzfLsAHcsw
hzpxUGXN/YIAHatj3w==
`protect end_protected
