`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
U9J3BF1OzBqcoI4K/GwfPKtJQdrDBM/TBZN2A+qoS4tOJbR8zqWh4Q7T4VdP5WNBlQTjd82vTBw4
nK55nCKb+qDMRtkztNieJTIGpPyPIKfGhrE7GcgbtValUhStfwbDvZwjy0s6CPNU2K237J80W5wR
ZolwaNHqIxDbgJ87YcWVJP7WLXjMirafN7s2vn662iyzH5APzEFnUETr4V669aUJRX/0VMpxet3K
xYUiZdcQf9EzK4AuO2rXz6Yz2/vCmuPbozrnOxh9rq9E0aqTphStozsTMAO5ehz/Hnm67Cv8ofRR
+uzHzmxTb/w2vEdiKnC2HcAIKLITTLcCdHambQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="2E9+5/jXKm0sk36WSKyoHpvuyZK5oh1GdQRQ4St7Y/k="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3648)
`protect data_block
qNn1Alj76UibWE6KVnetQLXfdTDxhPyfhR8l81kDXB7lTHi3Ne2C6dPlSCZ+zqjGhMeOEc3huWQO
bUPT+5P6YHh1oeFP37LVu/sgK8f0dixK/v0bzBLSWyiE9oz3Gl0W1M1DKEKMISfwvDqxJdPhcAM9
CXMphTo5hVlqIarCfi2DipONUEUxVXuspTd+0CgubE2he77qd4sOug3b6MUI4VVvTsJ5KJWkFj4u
N8ew/vC05xOdcM041XNY1wwwwpe9gVmhCVrvUE5i9LNI9+/d533HBiJUJQu82LicjxwP/dB8zg/S
kzlx/yRxEJ67mt39jfCx9fINBvp96zVW8vm5PvEAPMhrFIWCMwVeDX061y/I1RNHCQfRGo3SmuKZ
Xah3U6USRppODGhh8iofGwWkUcWEQA6VHJmSRvviyEboeNsmJupBe3MCHHa/DiyIRsPTm3Cm2IfW
typ062cCO+hTbxgZ07JPTLe7uzBB+MKP36ZLXhxixH9kZj3R6UQIH6pkKxkURw+E2CK1gewyZTbB
KFU9DA7p4rUmmNI13UZZvE9vgB0i1ZuPHP8Eqm5vUe6pWcQVnR1LMxCA14n9lFVyFL8D55ru1N3N
vIZBRR7i3faTxqYxHMQHXs9kTqCJoISZ8OKjBA6Z1NYfVwnSmGAL8xxKypuMii3C/pMCqKU/JR9J
346RmnZby+NfUPP78IKekW73wPXn/++fKAljcZVMoelCSW9WomN9Ff+QF0IQookBIKTacnRBRcqb
0e4XOV1bqiqBoSQwYZL8ZF13eeVVBWuzODpqIHK+7LkZYg6xWxu8Kxc7oNnB9Do+Qph012ZqV3lR
Ky9y0eL+fa8rG907mGFeM8qhIcwwlIxf8u4ryK/W5HDDS1vnY8FPRvEVewmaAPfWZsmed1UWyNs0
Nxn3ENzQ6WjbsHRRBH6rTXZRVyUaeId5GSHMsTq7haMer+bLxbDwnstrFgaDqd9V7uJj/URVLJv2
6eXgEFiMSSQoUvbKdj6ExMXjM/KimwwjlwDWacpe2D2VsmEeewP/fVa1WaMtRxOY9eM7dYQnl0oN
62z+2vG6fKXHdv/tzTprkeq1krpNzM5BB/9r0VHGssLwZ0tn+YKWrGEwnIbvpEue0ClXBqLwxDR7
TIZtxmFtGymf3m/KdsEay76FTbQQq0VVrg18uslloKTiBB0mflXHZ5KHU7ta/CF9oom/iMt9NCRS
KRLEyINPsU5i4gWTSBoOR/53SXfg7Dk0FgXpp9v2wx3Mqd5qDT5Zi6DKW6H8Fp3DUBzr2Iy1LNFZ
fgUUMgvVavsBxE5RKDjjUJ1OSQylFJxkO0CddZyyFTmVmvwnTpUmNtYEAhPIclbAAI/ohW7AOzTz
34gq9CwOARpVpUYfHTq7NumlgRYlElGjzlSGuXa/htgIT6g8IsH/wUU+l7E/eZ7n0zM/VlEoxzJg
nE3knF235DiTMmSxv8fw0ImZj/rLiP6l0NzDVPVeRVC6WeqBWbTVTL7IY07HhKdTTnKb1dns9u+m
BBxcdMwJeXmGFyEHw0sC7cZUrRkJZwOxmxSZVlyeT2GpW4TAFjaGdd+orfZtnIynhtQoLWJHYyKC
v0E3dLDDwKqfhgHpouKWgbtgVsA2xkDyqzdgZnYWq5YuxuWCf8JvPLsidM9n+1zMNlaohz9jIr36
MmHOk9UF7xzN+lWvdyaUQjdta3xXDsM6Kgf8+GlJ0NJdx6BidAGgKi/bCP15KUdDKL5ZqsYYVq7s
dGKxL2EtFz79WE3tu0ijA1LOUSkXOdDIYoBABnDx0mh02kODofMi4uE5v7f+noWBCXJ6EwhP87i5
UtkX8/LVRxHoEzeqzKlygF+AT6r3VvxqIfIqfz9YoVhUeWySzC23A3MI6O/epsbouut408irs+J9
vdEleIeg02t59SHo+Lju00BhgDMaFIySYITGk0e+PPNLmHzGlEmlAEz6SVrifBWXQfQLVSg/S8Tk
wkWdfk2PsusFtdADRNiQPH6YRJKqeMAsVMbC7LCx9N8fyfhe2IeuR6AYZp20tuTk4AlYIu0Dccvl
S7AivfKss4ATJEXY2QWp/bZNE0wTKwLdAoQoHCTN+fTcaB3NBmLTLxmt5umD1hn7ikHDSx9Tt/jy
0W1Bqca5cPVVq3dmeZtfUceJpoHJf6hR21JX34dTAR/sgA41JmlRIdttao4SJB2j1G8wyGwhB4fD
kQ1+5uTD9QUWOuccDrjqEKbjs4+lU2DBlW2hTcYWuFyJP5vMR3bfiWXD53uc5awy+ixrzdDzqSIF
b7FCKpYo9wvH3rjvWI1MnrHsHxiycgmS3rqhgzuYlKEME5WkG5IwPcZpw+FMvfI4C2lkmWo9/s6x
Rk2fRDdXU22K7ZTucZYlpCY1jBfGZIk0PqTtqZyGNYoqVHOjvHn/kj7k/dxzq350UylG3WRlzh16
SKJDSzIlSM6jOh5qB8xT9OZQFjXaqozpYluRDczBsBdiNLmcTRWtOlkMIMevwdyZPQ1TUeeUB5ul
5dvUKMEyjjEWpcC9sgmYTpVEs3HtJGTors2rYyqsMDjPU/lLwKTeZEAIACALTvgnstLml5esuNn7
HH+8HX+sIJg8LxGRjLunc2yOKk9bPXaabxlXUOyUrjRbhF57orNpH1rtq9XMnk9jUleTUgndAQCs
CfySc3FTNJDMh4wp1eaEjL4TzyeHdKZFOrke5tpRhKJGbuoURJFzDctq+CSKryHkKyxLwzCZRKD9
P2gFVLahtijm0Qs43wsBntMX+VKaOIHu9bIkkzI0RlgazjeAkPxzkGJZjKyaj/di6poSAhkdmV9E
64g0sPxExGoRmQbCKntA9f7iIV5LRxJNDjqFGg14fb4GiuAJvWCsz2GbGz/lDessvA+jMe1rheVL
qtiUetj2TZXQTsI4fjNjuJfVA13psickAQAntuLAtGeRIamiijLZ3DZNXcwjvL/6MUC6IYKLCD8a
qbzY4nwYICr692liy+55W3AuKsncED48NTBtZogUCiPO8qbUX3XbLFKk8OZir6K06RQuxRotCKYw
TXVByf3uXwUZonetCSlHZ+paVAmgxQ1t69AckChRd3RvKejuwZxkwUu4CUajJEhScLrG8JOcSYPq
1gAz0kGWFy7YbJ8yrVD8sI51usp6V1QsbMJjhyvKXHCKSRQy/Nu8WAe0JLBba/GaQyC72ja/aeVv
O+biR1nn/xmI87l+3i80Au4actbPuzOWSPNynfe0xtKIyvifEGE6s9/ROS5vkW87m61uLzPbFSW/
dFeWrbZ0fXnfDyz4SrkouK/ea92vwsdWGo+jGUb+bD2EylIt8a9tf4oTLSyLJFHEQZ+DXxQuQSXo
WSMw5HsgwSdyg2Zf/LEzBzgCstfszPXygUTHwgFx1aVwV0Nc5k0E7LfVW21GCrZL6egw6Xor4/Co
90gncK9ILwsppeNYQGJ+IdAiG6HTsb7P5DiAahXLQMDP6NV2mIDDqRpxT+sUqHZQxqe4I8vnzzKj
hNz/M4Fw8Vh8A2LvirvefWg/PhsuqRAYcOYgWUssf8dypKJ2EYm1NdAboxX2GQMIdkcVOL0EnoQS
Wi/wA4EFGaYCTTLfzLV4WfcVVV3/tLqr+wLK1lWThhXSnsERXzHlIDNSrR0MXZOAevp+oq5D5L59
9mQYj8vWtw8H94ELZ8DwDpAjYfcePsKu2yfu5ZD6qVYQmvjV/8Z1IHjcmKya8hbxEx5LXiZu2/nv
eRQ7Gq7Hid7I4Mn3KJVo+4uJfsgqjmBu2jhvmqda2KMHZFxbunitBcmGMGOBGkIYUq6W236S5AFX
MPoAgCWf3iVmTnyeUnfgvfi+Sr+9i1lQP/mZuAQMZW1cHROOnAc/14FUv5EygcmIPej1D+6Pp8s+
8x2AsVK94DZ87bcPkNk2r4TFzUycJy40zuA0ejf5gDUun5hEV1eu+KIN4c4zsjnvT1aM0KLxgDa/
sobkc8lyXQCQt2AvWmkM40b2nzgIQ7qZrBw+Oxa5J0dky9bfyczTA+giBkxjIU5hDtExtJv1TpxR
Zz7SbyJnddp0bc9FPUb4dkR0VoXt4URwUrD1RW87Mc3wh2Bo8tzt2+FaGCE6pOlZvFqsmIqX3PVD
E+4Eh2obJtNC6r26eB16TT7bCPbEvFMM6e1mmnP1V2FR+aRAaCnLQ3Y5cIjOnfFy2mH+LfcdSzIt
vDlvr0olqXkcNXB9JaPdfQ/FlH+3Fi8AdhSkFupQOICqaepoz+ZHfM5/Wfxz8l6rOJyoXmwqChiM
m2PJ3wB16hC/k5i8l5MdfrS8P5owxow8IUTn9AWFv5WcPvuu4QBNQs7Wi9oG8j4/fvnxABBCEisJ
caVCXzygEfXbE9OpL+JLRF69dTSQSP6J0n58GHmE9R/eDXpB87IrZ1mPIPyqfhUsAJ0IYg/8yXcs
9N1shcStMi/R4LeiHR37cGWi8LsQ95Cc8qPrxc+31GyAr3Z0mvkjy13ZDj2I9LZKCCr24Bxw929/
qDSBkzPUdxVzD6/+BbC7tT9c+hqIQD46S93mI/HrPd3n39tpPaP0cZVJElPa8IKfnlUkbS5xI2ch
tUJcfUvfZZ96CMqYmI7HXBmeFXmeMemP53aht9EMhojbbJw1Mrl16i4R8KJpED+f875Ce5IJ8e6/
ahTzpUiQC7iIl38ev7FNFI7vQ1dibW0d8uqe0fnVNKj9QzsFM5vHlN+QCDHuoCEWNuYqu8bK89Lv
Igw6stzw85OsIcsS/nwBn5tUyWfM3pE0W38oFGykJFbD5TskUWbN+UgxgOQ3ELJ0gzcqnnv7JQpJ
lnZkN0Ob5pl0wCX4UeYScUW0c5BBhggS//zyaMuGSyHfpaFdq6THvIGuTMZ7gl/31KPnHcRgoyhB
`protect end_protected
