`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 73904)
`protect data_block
O9EwfxGSkaOYId+eIL/QCLUoKHuXGsUNpamEveEtsWr5tLRcDO6jcV6UyhMmV/Cm+7hpdKHdfant
Nko47fPJ107R/VfIxExoLUZspjWz3e5MvvhRYLs5EFs583cHNa30cpwi5twD1TR0MqHU7euFQa2P
/4v0EZz08ngGDAVHqZ/JLicSw6+TG64db5Tk8+lcQGOQF2uqyIr7qGXVM4cDAzIXmBsxthA1/+U6
NJxGQp77Z5XEn78WhXgfS2dNZQS2enEiacW0zz3uA0WydJ8VMWBkJQGxGs5TAodVM/ECXKFhjakH
8nCAcRe031W7br11DObLIZjKNPYxZUEFqQHmGgjtHP6wG80CIraXLAUiyX/EfDzZKpSQiEPC2jbQ
FTaaO4ERGokFpqIBldGLyMZ3VK466LTtlW6aEJeefvzx+U/XR8KHdALqm77jfoQXzkETkeFa9JRi
pAB0GGLYv7C8kGphtRI9NjUZqavTobbkC18icORvH1tBjgngNwJRALr5pgoK0A8YwEo1BdjmDcYS
VQYmp4orP4fooWq3eazct0hLRWcEXetEv03crYvMfmpddXLFf4juboOTsTmxdvEXMAcBr8zBlA54
Ivhv2GieaspYvsN5Wr5VUKnXTtUlJsdN4qLt3kYAHLVoKI1ftFQIiT9/PO+hph6b6rjWhWfYRk3L
6ausAaVO7Pgwa0hub/ZcdDeMV+243A7iXNgdBxeLakuACUHtx4H6btomymojhNirYCYSF5C770hZ
fTXo88+kwzVKNYyacnrlRI1LUMvJKXT/CuV83xIkZ3ajw0A5yqsW5KpFOyfL+yOWNN89PKDVckj5
2qwcKnmCDlbpvLGjUattvEw/H4/zDnAX0HgeyiiZI1/uUvfbr76EuMMo7jfsaJhRk1K3f7gYnL3k
6pp9oX5ioh8bMFa65mTOjDz7RS+iraGqpVedkI2LR3sZFVEEynEre1burf13ssgJoiCzmwmYf5iE
f37+rMe3aebL1doM0KvK93UNknID5jLBmsBbbGtaoph7NiP/ed+thC/Ey4qRMjcRhld4+/Zg5Muj
/1oiWeE099QhKqrjrtmct8/vnFmaGZuSFAWdXesETbfyPoUrHU+QiECe+/lY0zvkKv0JjidyHP2p
A4rGqS2TLGyRXgWbkJ+emzIGSI98NQHm9FPl8TS2bmxyJ35ZYlNpM9NDu4y8H81nRYOB1x/JVEG2
mbFHBebDMCwEzV8j8nfB90J8Zw61Yx6ek9H63/IV/25Sbxn/MgTHcrFF9Z4lPoYdTAs5TaKKQyPy
rYQyhYazsQZFej91aG3GwhcR/8ogKSjCn3+FXDcaVpM8QUAGQPuhOlmDmonQs/BKmc/tbDZpe0Im
H44wrAaaVccnk+Khc2ZTTZ3Bjp0KieK1zqh23dOEhAZwnBGK9jmghkVFkQnbIj9sXQFPZ+w8P6O1
2gqtJy97F8JkoopIJnDzPFvlDXcMeTb1ivMvpT7D6gTCS+QiGkW0r5lqw6H3OkOCVR4H2sGPHdVE
GmUt0iTRyTqGEwnBFIWu/+fQvPn81f4N5XTx1OoHWklHWgAo9h+L4L9qTAkUe7wljRwviMR2GNtj
2hVyWftejJDnLdCyFM8YFj/qJoNbfvAgvfijN/LcUyJxk0IWKEE5gVzJGzuMdwwhlBjycWS9H+b6
L9S2xHpX3tVCvsDezW/dgtVG1BcPSjxB2JlRXBuL8z9axi7MTCGs0/XASL8MKVc0C1ds8LsDgPr7
11tGLl3/XwvwXEwMnvcp+1+P20ddmBiGJPZUlFXwROctzQdjw25pTdFvXhIkwJDTTLqkipE7f+Bd
Hi9Ij47w67nSobg9uxbCWMQk0ZhohdEALXWFM2PZsAElW4D87OlfeihD0yCeb27SBG9ui7YytaPo
g72+a8xMqpFGoI7Ga57XeceLEx8P6JlrB3Gdhv+ICjN9RBfoZK1M+71OFkx0M/vBF3mCxcz3Mj+J
ofjhe9LLRMbAE9AeJVKOJ3wMBl8p3HtrUYyyc1C/gRITw3czrHgcX8p4a6tbMxtFdvcxmKYzwbnh
UVfa96KL7WoCZuIpzaYUnAisWPBXLfm49OMfZv+1he+OQbVlskS/+z6zU5OqU6xUgQeIKq/QtFPz
fTziAlanxIv6rtSbK6itGGXaCUO51wEHWMEHVZbYgwTLqfuLewbLGXz2VM+Nq8TlQA9ppzaoO8Uh
3Wg/4VsYbmuTYOGGxhpXeZRDFYNTRpw/cKVJgj9RVeyJ6A6+laHDMgazXndQ+TEZyyZbeIKzTQDQ
AdtLmFilHso6DTtLvUFZWnhv48GYxW0SVZLonlxLOfCa/mflq+xDsECXgMK3OD3YyKH/IUN/BWlT
b9iZ2rryOHHkrmB+Wl0+tjFQUamJXqckT09nFEweMQQNirvvOReC7kfWYCUULPI3Vo7oYyo20Tqd
NIkfzeoxZhpNUptK7yWyVml2Kbt/ai5LmnnqXJda5MtEDpj99FWw7a0ee7EIwzRrzdL2vGlcAP+n
kkckIc2VSQM8fGpVzh129mPP3Rthg89UUZDO/sg/DGajHyUokzrNGFCLbkuwOBDVRPRPaODSqEpi
HDFQfvEwgeQlsGzw0lklzS28DyxG/4/ieg6vSwRnk9p5Ca139UCgdXVL1olnKZ4kp032RxCBYJne
nYEDIWedTSThY29ftX8re0Xf04KEGOQeJnytbRbNYzgZ+HOKKq6JNBkoX4kOAAF2GfXBDnto4Hxt
2uxf94eNq/lf/o2/Ke5L9yEbf6g9IRZgH5n5AehqeCdu7bKLbvum/rw8XBLSoBTRI1fgY2uExqfc
nycoF+G8HLHPe6uv859yK4C1HufdejN87QUfuwd4OiWH4QKmllD9k3u0NfpzyyjT/4Wid0TwJrIs
3un+ltoRB50Dt5v0WbVXt16RLP1ppuP5O2PlyF7a/jYb3r3fQ2J2ZvWPI3G0bNzxvQYigddeL2QX
F2nvwOHPJBWwzp4NhDGdpvv1+hrN92ykIColvokX2vZMJnwCTP6sKML6GU9JB53FOKTxUjsk1+TA
KxZEcllympZJIPlkKspx1xDdt+HseaiNzv2spuhp1Q8+oLXdIwtCQ/IEEpoX2FzrlmPl1g5Bjk3M
JyjcQRd+Kq/ee/FhZVTd8XRQAx8kQXgxOX+2wCXZBfHlBoCXHAB+OpKspMow4mUdLCKc9pcCV7qQ
31d8Rl0xZW93ly9pfo6DgYWpNCN+2i+qjAOZI69eGlC69BNwyPD6zxWeNyTTjwv4hwKA2eRNuPAb
8I6VOm0+KiJaUHLGrfLpKDXPPMf7OK43PeIdOT8iP7ZX5GCZHL0r676HoCgNU1MsbmlefcSeuiOp
2tnI1IjOWgMhVlvyHeeLP+TWK5rlmmtbSpGhEY5pPUvYfS6NmC/TZ0CfyKIZsq6MEH0FexW1eCH+
7MiafMA6A6CmV1NkVxlkesfeYQbkA2SVfX0svgSnnCpMh2SdEDn/+Xc6XMqanCCmwKo7vvEcSFvE
YrNuKhZCQLxvV5Nc2AMhY+kEsYsq4qyWUXzKBfftGIKMnbJ8MZ79rbPEx9mO5ZIXbkJ72+8xJjHA
i35aoFiEhGR2I75vNjl8NAIx/B5F6hSYtdb6tlogFG+flYb/WfLGqguaSPQZhP558d54OsTD1w/P
kFup0xTj/AKpG84BCZL0e5KnJlSzyebOV8ldQBdEcijXCB1s2wWgznfeKFI9TTQXWcc9sDEA7nMz
pNJlwaLZXN8/SrrBlkq4AjI0C5PdKHeertNBI0OBKjHmSpwzElVNdUiJQVOLQsesBHDr2FI3T0+k
MD99ym8j+5K+SBXxyb75b+2e+FG/2tISHDY6CWw3boP1k0gpfw55ipq6fTU2gJQBBWZXu8fyMrIQ
StRvSck1nyysGgjEQJRn6ao0lTBNf2pg1xKWKXR9OwRlDL1EMSW4aF5U2ZFWdOhTO1NTBMrgcEaO
o/pavtyf/GadhoaHksWpG1UGg2urM7kkMMkUiKuBRgbC2YjIbKJWxipG7rYHKY5aRlutbG6cAtCL
oOdlHT10T8p+TZo3o77jd0o+6kMeFbYEdvOPepba3abHbmJA7x2dyfR5iTyTnfn6SOI+pE6GbQzH
j2EogXpXFjnNh+t+/aHjQn3TViaau0ND9DphedmOKlhF6BdO2c1B1ZgeO/jQxqnbwD/HhMiZ+tMI
lW0o+Q1Zraz7OJEf0gtnRCyz8g7cd3IKcANx5GdRRTcCGdV3egn2kFU+61R9Oy0wzn7SF9aXaazR
Zl0TVcXE/+rb50o0heA68YZ93FUlEd5PA4vLzCEWb59oqPutrFl3eNp2oU8ekmvOhE19H1TAz3YY
9ZjjDbWBQ8mfA6Y530ABQ0fD801LpPkvWgjJ6F1oB8aJjIa4K75vdaEe9KTPkASvvfLT9L/SbdGY
/Qe315dn/tNUi0AtGpLUvQghqGFQMKIHebBYSPWozmthil2JWJUtz3vyjK2cxHqjQhlImfgi3d3C
aTrJcGtvhit1zNZEvz1nw4aFGUZ70sqMZpN7BHgDKm+bhEVmeUmnKrGvrclhhZzC0tf5lUklFioO
wJNf0FkqffKUieoEi6UtjAEcWY40f2oKhsKZWbZ1u5KmZTxlWdZAIcTh2gHXosW0V1qgEYiurc8u
PXOvCHmEuGwJpkttECYDVvRdqCKvMTdpitGzBiix8UIQ18SiEXskHH1lvESKiJRt6GJzZQl1qPbc
a4Hk+fmvSfR0dTxg9KGNH8K/dtCQsVVlpJUzPvc9kZ00Fkvr2yPbwVQIF/Mhc5EW6RvJhOgfsjqN
BRRKF1ysR0rfAs/2YVM0bv2Ves371IoSxCZre68hdZuJuTUPFx4RbE2VG6URRzF8P3fciAd2s842
y3tiVA35Q/tXMlAaPvFYLiIq0BRt2MNfmaEFbRVlUr7DRXjbcMv0/AESdcrGU130drxrq4aOpvD5
arJaCdP10wflmLyHkbkEBYGnDtqSCWbTAr0zoF68MnIRq63pLWKASqHUaO3xWqsJ49rIsCvxeSX6
6x5BL1ygOdgZNXKn9MH/d23n0FknTYU5nm1RVQxcU3AsXCJqwNEDZMdWxlY4btKVJJGbqgOjiUUw
sQUXADTivNjDDNWd0RImQBnbCl0MW7OIJchGqERsJ7Q73hzGrZlp4bu3aws/rDVx9UiI2PoA6zqH
tg5SfsD2JQi7dbEKKroYBWIKcbBLRnWpUhC/cnZ/hDtAVrRmUCPXx17+TVulmKxaF3EKbP2MJsqW
H50epct3hvsI/Gnd/8xyNZ3XIs3ph0ZmCAMnzWF+XT9dE/znzh7TcbmR0KjbsDYfLj+0s8E2EG6u
M3k1dAqDSnxX1HKEpMPeapdt+h/14dmTnwoDtnI803YBbptJLLy35Qo/X/QRC/B+PS+jEnVnOzUl
653PkGcaGP862wHJINbbsDfRZWkYsO5LZd1RdhlSags08t//Rsaf3Do3ZR2UOPzFu7ZfjrOGHjlG
BT/Dbe+MV9Mct/Wn0YfPRaxx2aASC1xk5exjT8JQ2LmsjyoudWuZTUjCRKh0Awf0YREsZ02r7Hzw
AJBh5uMz3Ko5n7tvSqXOM5H/u/X0G7w+3jel5t99qgn+1pVK0rRLcRYqZBbqoCh50DZQpiBW0amh
iQCkMa+Ixk1Ski/DDOZZ6ehqJRox8xucju2I4tMKcY0LIqbxUy9zdBH+MQLZLwK0v/RYE3czb10p
teKG8ukCbD/rmwzwXbWGcPKoLNOE4FBBXuiNnLXCBnqwxxq6Y7/bNPgUZPSAhD1pY7JPO4JA6hic
tQDdkZsbHfgQ+ccLx/i+kFq943HPDApie5KRkwLaR4qvPga9tN8o7nRXrtIHjBf3LNj1DfCerWFP
CPYAonIxu95fvujnD/b1/u6jYnUynyUuBE8jOHWDhIuYW7SjMolqloYXADtco3Ebf5QoKwf6quUj
ZUo8/T0/mTDA2etQ1hxTaRENi5p4IWjb8amS53qCQiDLZQB+FX5kHw22yN4hGPyL0ZHXuP/CoYbE
FU0jRUsWXXRro3/dhY2wCyL24RyO7GFm7d7cg6q+xLeQ5BNqQBAIIgkBnUICI63Lg+8nXcbuWYg7
LrElrhNf4jMSlHpvnOpOM1WTs73GXgWPo3aaTKEpOpOwcXl77tCLYXt84LbnU/bExxKDuumtafB1
ok/eBynENroHtBYaGTiIWQDEDcorXfI84f2CRWuKtb34ok0BYMhDzdLhMoqrM4Uitku6J4uZ3JsZ
MUvQWNVU7hBwfSoAxTO4ft8sIb2MNoxW544dEZOpx8T1HZDz2lSwDE9ftRHDfvlMdggL2fQJ671N
1MK+p1EOG1hDKxlskyU8riVzb/ZIs1f4HHC75rtn9OnmLZTLL9nm9zXzw1nJr2xyaH3nxCgYgCSb
7tgAVkm1vunIauxJ2QYb8vMNtqV6KsGthbhuypdgLlcDsZQOLlqv9zBijI2w+wbp4wFdbEFhmd7P
vWjLgDpR+ztvHtvfMULcAygjjZbaWlL8DdkpcNRPDwfcfLPD0k4tQ9xL94QbYfKaZOpkiix1inc+
e3H3wyhoDU9Q0iB8pSbftRIa8TrFFrYwRRtGlgd+aJNssh8+sPcs2VSyBgWfoT0/eN6yMhAfpQxK
ecP5bWu5eQvRXT6zGASPf4rXzhKyQFBkQinXdKMpkdl1yDbdcKWd16D2HBfDF1om2pM23R762h3U
wcr6XePcNlPhQE6AHbIg2JvZiIjiGTMuTcwvAQxdbnZymhZZqyAxps/3CkwH+SabJx/9SlemQ8ti
ZqAtJT05vrsHmgYUzjikW9Oi2LCq3+szyKcYAUK9Sttg/V+p+GG6YHA81x+W7Wm5U09JUo6TsXwo
r7mI+jzM+mL99Xqhj3bac8oQONXVLPF9/U3SgkwP4aQFIZogXEby6Orx3oWf8XjhBNlevxsL71tk
QPW6zHyG+3snv0d15bKW3jp+CRNn2L4vVPA1d3kgOzdsmxsd6kl+KEl/V+8/X5YXh+HcEhYoaxFD
GYk2siIe1z7OxiAb1NIhOZUF2SGt7SMzJloi3FYyANWTDt6A9oQCjuo3zrRoGC48GDkRjxNiVT7Y
3EuODhyVFJuOqHDFxHe1i9XKWi0b20sGj9DbvUy6z581fLwzQ14if/D1xsZtzRTLmuwkrnCjd9fi
B/jFz+TUrsllRTFx6TrGvwvym3gh8yAfib5po3DmxtCCiBVlW0rXjT+IEX1kHqRtvX9KHaH8/GH5
NLiFrt/nFy/gCVQga7WeOFldcso2UfonCJEbJi+dl/0Tu7VTapFedtRy6jqqV0QNizVfg4ue4Bv7
seXIeoBHsS8MfVFwwGp2hlJwPLvLK+5QSZsygMaZt8Nn9AloBnoROy+DP0KsGDYLGy1UVtydXhWx
WDzpvw2wqr8b83iVXAtbh8gm8xhVDSvyrVK8MqM/v3AZdjJO89fGlch8Qt6mlEgTYv1g/YvsAuaN
w0ssAiIjVpdHhqNCdw44K2T1czr1GD7UG9+6LvyKTvpeSieaRVIe9AeZEgRgSyUZ5ziZJZ3CB+Qv
HW2tSbLvIk4GLSzqR4+w/yZSEzuAcy//6RZflmlshh4/pFwycXNpfxVQPHPGNAwRx/XgF/XCI+pR
XuLHdtzojoJiQwpIWfdH+fY5mTEReqhSeo7LVg6pqe1QJRf57j4wuYiDz75Rx3MfzGu/3i+dp3pT
Hz6ZGJT7Ko7q5PfsS9wxGXY5fMplkaU5ni8sl9+bSANGYlu/0xrY2IEOYix1TMWIW4oYCSDqljaL
uXBSjb2GIQhx2uZiz5rAfwMDF7Mmc8XgmNtG3wA225mXtjqtcCijzo8nstpwRLfMNL16eo1jUnjR
lONumKc6DjTH+K/DRwkzxapb0qPO6uRbWPTWfTgG9sx7iyq0hnVUzqHstvTCYMgvvikSs7LqnyGs
oMTCV+H/iVlesEF4ZLFWklxG6AH9gmh/syCen+DcXDvfMBGgsumKwzdOTudtzzNwP4wd4dkV5rB0
sDtK7UB7m+iCBrkqxmymTYEhVdg/zvMlicI7aE8Ro+C4lBicaMj+xdZBECqXB1afPUI8zVXkRphS
Kf9VZWMKpSNng2jhRbNEytJWp/AdqAC6UtXGiudZpNUETrh08oReHfzrLDuGbqoK5iVfRR4PJCgJ
AYrw5hH2ibhDS3F3l2z3WArLxNXKNjtg/AN+SOJ+EcYAFQ8IboJt3rHp3MqfjQfgtYUvzeGrqvKD
M5FH8r+0MzvGlmKWDOKC7cKzEgGBQU0CL6D44qqt5uuKC3ak538J/8x8cbQaRLqg6nwwWdKYaLw2
SyMvV0rEEcQVFhqlbLBkFNKpUA+8G5RiTtci8iopFBRaaouY7zwRfE4hYVJsDUxx2L6vA9rq9idN
3/8VQKPE+/sDHBd3DenZGSj0iH2R30XB6nFraODRCg32cjb+YI6iFyZnnr3BwyNz/zDDylCJipRr
B0cKLPhTex8tQL6140TyN5n7IDukDuena0SG81bE8lXykCqYGrvJHM70Cu9d1BK5JMt4CHNQohTD
aM6qyK6WrnllsDOMx0KnSjlwWiJgfAoAvHtaPsED7RNFc7umYdiRKQjI32O+uipJdBkBgxbakQJ9
SV8m3LiPh+VeGfR7HDXTRYAWVjql2vbye2wBIG3bllxAQhfca6HaRUsKPj8CrP+at2P7kSlZGvKb
x82f41s60fzgU8Z4ueaGR9wlGJtXq/KMZ09VH5X0BqO7o7QlAm0PGgaSH4jP3Dy9Nu7x4Mjj5b+V
ZKyQ2a5jbf6h2OWgDs6iXf33YUuH9NhlTf07NG5ycokYMAyVo0IqtI6iSz9gzALMeUfr5nKmGTRq
sqnQ4O+eR9+V+FgeA8C21rsbrjAaMq7M2I+CXOU5mnk87qasTEfh6sAnLLbsCh+lxZlLYjywB8Wv
bngnhHSpd+pEImJkkiDxllQ+T1q/NOp+cY6pRTsakrQPez7mo/oevtHuoSXEfpEqBO5xUKYM8uup
uCl6ZigCs+tTasSok3enuQIe8iweB3uIUVO1ufJEpRbJXUakjzRGwJAn3gnzIlwvD/tDSzyZ9eXc
Ysbe4t/WW1qYUMlLcS3uLkQuspethQa/2VAT1VqbLcIv6SboUyMilgAA5PAKVC+bs3SHwVsbrRYw
AIaWW2XCqxf+Tq9gzLJtC3pAWos2bbbNIMLngrxXIhqGq9b4aWXdlhZDaGKD+oyYFb0L3hWj1S5H
M0E/XyKOUYlODNXUetmRyLwBs1Qa0Yx0Nh68PH7vNFBxjkEcrlk3G/2mKvOO/kPMvafUKzXUFSF0
NZJjE+vxH8guQpiLS3jTIoIsZVsP7ai6wBwr3714SyMOmnzs5DfUOW3aVx6FOG6eL1RtCO7+mF7Q
kOkUnP83BTTG0cdKHY4ssnSHfvUxp6+/0k+RrUyDirhXiu24TxZEh1BAcm/GeK4mRLMBmJH+cIwC
etlGVoNpc2poPOxS9pfd+AcWW7S+mR3vpCRsy02SA8rs+gJIjQVs4vV5LHSKUItY7lyI8klxKQIY
OO3xieDOnZayPWreEwmH1L3CB/sX+zfKZrnORh5i2dTk6ncGA7q17eI7BEQc2piZjVQZ8sNebTKB
pusbcU2BuhjFIzeXKXj++6W3hdXuO9ZD0GEYmNGaSMQt4rzGPQyF4/pC4uPi0TaFqZ5+vhNppOgK
jvC7jXbHlk6HzTcjZTVRoBqh6cAQvAu9wCkpn6GG3ObeWB7v/PDp2yPD5jTTmqzeNojfOHQCoULq
qQAJ4QrkBw76waVdlGDPe155DPXjTjgi6LyLLE8oaqKzocC3YxaHAn0Ll5BuzsWrItlUOgvUb8Er
DHxsC3iYHptcHfFZORQkEthaocSZUeR1gH4uLjMzaKHxXQY7WCbwhxwi2GwOFekGWwG9nNnu1gn1
3JHkUniasaLWbYwHWq00yLL94qFZ85V1kf4quox3+OXi5hzpAYZK2f58awoRraiHg6oLb9J5ozcx
/zdfoHoOKtb398NDgfVGJu395za5vPdPnq8Ha0PvsbFBgeRcUkVLZrkD2RPe+bE1mBU5lqJuzGr5
G45s+dx2RszFDbaJ466/+E+YNYA2kso8KFP9BZ7IsZbhJoYXjN+OeAA/6OvUMDLC1RDLtXeIDs2e
emqNKpWDcMzICaWpLVqR52x8aPWaZaApYyuYPeZp98PxeyDSafLi3zMWcGKwda7o0WKEZm0moWCE
93DGOjVCZjLIwz86V0F0R0/MKptgnkDdr7VlPfSrCVrD5h1MvmrlgEXI/Qjcs2hjI2gOgeXvmPSC
GbWbqmhXNqBHzMWgjeysReSiUTJBB/cP2DpWV/RaXY5gmAlpmwBfds92pmmc8UUVrd8bmC8Z7LT5
58CfdL7iNjsReKGWZXzjNM6vZIBZwMPJu2LsbDaXq9EhwKVAg+vvkrCYpRjRdYiFl3vlRA0vsFhU
sTHX4Au5TbsNrfgX0iT7f7Kpox0oCJG4JtFXx1te1zOTMMLsCO7PypAAe6mF0vJ8R6OVYETlTmRD
bIaSJTYN92ZZfnQLX96fma2IbUnPSxBpCYuMARDOE7yT6/XPqXyQ+1o394FkDY8tgc7CKIuR4aVR
7Fal7BErPayjXuDDUxm+0PZIyKjBIOhOqSpPx6b3vRhx+ctnfpyBS7XeLVFHNfHzXOWXszodExx+
hLScvFa8+c761E47dJbBFcVn2L2tZS6cj/5OpNW0j7MnS4uTJH9zfpZa6zUMCb1qRzCqEWK517FP
B2ZmTW+RSozrCihxRZHunk5OAZsP7scBvcu64N9sW4vU1pAdcHCIcb/49bZdadrFuJYvVT7JxSTQ
nf4Njt4bbTUg4YY27jXM2jvgCPZ+7B4WJ8om3ynE4hZF9EUaGadzA3/ai19hn9E03r+IwJIwPvjc
JwEq+28X0xS6fv1L7qwTnZFKPGRsokKOHhBMIFyYL2cfheJC9/X3ons6E4ACQM7wfqwGTxp9ekoC
xB5k4SjWRTn3+r00rID5srGUZoUo+98TysUUeAc1kQaZHpK36mh4Tx3K+jDMb+sEDo+PJCy/CMmo
XjwazE9GQsQ9EczaM7zJ/z9ff8S/6QRtbU5AOPiScGty7ZAZsVCd3BmWsen6OyfGbizQhqQwD3Vg
z79Fv52zQN4LP4/+cH+xkHlfwLDH6nrNoBbAi4NWtDu4rsV6WNyD6P4y9yJn0T104/7C1g5BYP3p
iBzVpcnlIXjFYTCKdj+E4PRTjQMwywe6y8GDBpBMW1JXYcZBn/yjhdDsSI5AZrnsafM/io4l+/f1
O0IeUvdAY1DAPBm+AH2gGOT2gUx/SazMlmTOl2rD6xd+xGYSiuHT1QviEQmAqD54NNGdwaycYVg7
I0UTGU0XdXzJvwB1CXHvloYXaFjzu0TK5FDIHDvcWKD/fpb3573DBSETZWTNeRnwnkF9662yQbAy
ljjtVXwIAMLq6dOy0eAclz/NaCNMS3cuMFBC/r5er3PNyT1QDE/IO5vQA7jaYtA9/yp6yr7H+7iv
+tbNfG7/6EQ3sVNZ0lTmuBQggSOLyXWJTactqL2i6U7Ko9fqE82pEfAeniVm8d8BroCwU43O0HIh
nxNNn+npCM75UTgWVfDvIB8GHk5KtxnzWgKdhNO2mQfr+lY5qh76BEN++mEqGGX+5NhYoA0MZMOR
HAxzE7Mp3nKc2PscYemcLxq/slgO0ykB/0q30J5VilcC29rN9VkTsHXrTMEb9Rs36Zsb34AapU/N
C6Ix2tgpCqFT8Y2JF1+tmpkVn/HmZUIDXmCwEPksoS2Q1CzEwdos2wsAR+O5LnD3GTXQVuem/YBx
yHWEMNvWjDnsimx5x1gIbqQ3d//zbnXXbGbtSrhr3u623uFIt1/zguXbQP7TgLs1zhV/h3OVFuND
aiZvdJOwgr537FYnSEwq9c314bjNqVVM6f0lO/bf0aGQl/U7n8s/BCgOlZqMg4DPFhG8TYd0iHAZ
92rEj4/khijVv+YL7Ed1uyRCNVT3oM3tMhenM3VckQgKVQi6/cesiuV41isTEaKwS2DyoXEg0eTz
LuVBcXhdEE128ZhNNl40lQ3yu6FMrI6S0n7HLuGpP59yyC8Wrkwgb/xTDAMbhv9AQ6MNr9TtqAIV
nM7AMMRia8lW7kh/gPT2lSme+Dn3lq9b+PPaWLv4zWUAgvltXyZIToiKGXmOlvf9gR33/fjYWifR
NQmgu8JIXn8hXVkLd7AjZSvhwYt0G+NzNhXZFqOIoJFZsjSGM234myUOG+8Ddy73ZOulNc5RoozR
nsNXILRS40N0dOXchi22bkCM7y9bECLaLQ3DSH/cFPi3scGaSCSFI1Aq9VYZsiZIj4Wp/kStI1Ay
JQ2+dAjmTADyftqC9SA5mY5W2a5ciRuDtCZou3Nj+HGhjV5k0CDHjyKcX5PR9htbt9n3KMYeM2vU
eEaGTPY4JZgvro0fBM3FgQBcKyASlzjwrHm1SHVGhPl+UQmgpQ6fB4gSqmQJcgdTdXRW7R8pq5Jv
vYZGfemPtnssxa+KnbejdR5RyN5J7CF/FN4uiOCBdFjsKBC6pAC5Pcj4H7AD0DsYlnM49vD8Ey2a
nARHHWNIECAyfqtg6t+gxf6KMxneEVHn/0OrxCh9lo90qZRboPDwuDLRolkhkPsbvnIpwVHRuu+w
gqihQqa6k/9/P2hWXbSpUdsZrbGlR5Fl4klfjekePrNTxNpIZ1Pj71Bh/wdidhcUVo5DnvBj4ayW
19maMt0mu02lGLiXoG88TG+tTA2U+aamiRAIMvKEHEee9sJWorsSf0VXYmpPNTI3hJk2gONFnvm3
RRTvdg73gQTtRdeeNk6EHZ9ZJGOoe2DSerH8KPPm6Tz4Rw7xcFolzCdWerVVng+lA6azcoWg7ckt
XHk8PfoG5zBo5j7YjVY67lN0I7W8whVLzrITxMnKhr+F1VmMf9kNcqo52RqtwLoCw+3ow6MdLvHw
CP2XS45/E2hjmZIJVU/1jwXViylApfnEXuUeWryMcJdVvFXAknQHyEJkKueYhb2ENZfy8SV5mu+3
imMJmw6QebXA+h2PPTVcpSK6HR+eEy+Oc8XL0E0LD+npl8exOJLIyHZHBJDBJLpQlzvapLhuWZY/
AVi4mUR5/M7J7sG3tHoGcX7dEFXC8bRVxrA5DX0p3J2qsVfGtqn1tcwjZ7lGhsnlIBMccq8/OWdu
Zws5Hjb71jifaY5YO/GGA0t5pF8rBDVwSGurI/xo8FRKBr+wArXoWEJp3RP9orOFov3iZAxyATcL
3Ql3ojiCA986UKIobNFPotXKQ66D5xM6YJwMuaTqJOSpHEq0JDuTEpPmG0LSdK0YFZUmavbeFhV0
1PCZGeJa3+jIoKYtT8dHZfFJ+1okWL4U7voSCeUj3ZwsWm/v/WwZTA/iOH/1pzbkNKgQXHqPQd72
3ndwzoX3Ldash+RWj38qvT+d1YOUPHZfC5oL7oFq4N55F9PKlGPybELJSJGhgPdF+T8Q7h4vbclo
gdTRog4EqWJZT5r5S0O56lM2XVqOxMXBuSkICzs3RneY7PxUboAvBvcxzxRabLKGRJxdNfr2UsGG
917LWz974WTGZu7Ulp/1LGzqW/uZrz5+efOtvFGEH/ygwiXxd2OknAmZagjoOQYAU1jFosaYsXML
nWMUXpiiKNTHKY6pji8qtXM+O854k2dYMlAFObpGioY7xNBUXyw/4T7MCoUh6Xv3mnbMzOtQ3nrn
6mWxP7taaJy4nFFHgqqSNBhmHLpczhmhxSm2dME9Qs5vNI7lj5WskIWydcPu82qcE3IziRSRm/4I
nUiKmz9JB61DgpGoCK+K9Xdq3o42OsloaqWy70EUKPWsevo7yjUJGDUA4iuUQOmrTKAAjzYna1vo
F+Pw8StUE1unGo4u0TOBshW6Gjz9Qkjo7uxZ8ngJnU4G2Fyw7a8oymX7m6+WJ3Aw70YLFKGkRkim
8rzptJjxF65Rr4oKb4mxKe3J0kflmDrsF5BxGLGEPQ5Ws+Blzg3mdaZLzbaXvN0ZKXfnLhnncPBo
4EE/x4db7oPqNgX/ofN2b4TE6hYJOdujrpBQE5UUcZCvYoViE/tUKBpbHPA5Os2FfVr/JzGulhpe
h6r/m8ovQn1EUtcyoM7osh0F7dC/H3Q0K1xmAhrxgDpPOXcklej6h8SfHccbTUi4Bf7v+1hE1V38
2ZFmonrZ6948gXhzl9dQHo+mQTGsRY54lrEE6L7P/jBXp/0KuEcFwQfwct5qmtIxWMvWTFhyKkJQ
l5S5C5boBfk1XTzNAJNs2qg3qOHcZngjDxz5Prn7gueMzIeoqVfS7Spbqt5bTVW+lWk9uy0JB7xW
w0/VLNpoE/g74OIiCZeeRTYpZ2Z87n3WlKNZGvDpf6TL5Hkr7B21hrkMMnWBr8AVdJXM+Ma27RHL
GIA/glhJp6vXhW/13amiC3X/KB4BjE05JS8iEsfN/bmuh7Y4I5O5U715doMDyh0zQEbtyuH2Pcpt
39blv0Laua6Yk50ljAYDkeCNTHgkoM859XFaqM/0P2B5snhPccTuh0I/7fpmm6gBibZ8MKGEwhzp
zsirpKlQtzdfoYJlJ4p5rnRlKY3x7rDs5A8Vh+Gs5KINT/Hz0gSuv5Yv0/WMRTuxjQ/rPZ5Tdk88
/LWe+GIpMFNiIlG5oigyJKv1lJ2T9yJrIiilmYS4i+LukKvWix9tPqSn8eeGd1OG919GzGNW4PjC
6zsV96IY0PQZpio6qU/a0dsKJUsBRVq4XLdMIHvuaP8dsZFmdMId7lHy4VN9gjXOz6pXuFfsEIxf
nl8SbKRQyNWkjqrZ0Qbwx5w8RuUwU6pQnlHqbAgHw+tEjw28gIfyC4PQ7L0kUBRZRhvwgxWB9s4i
pjJ2xmA8mS/UicWf6+cHKLscrNvTGxUEiuhSDbVWXJgMCrhnW/9EUKhxJxa7/zXJYQhme9Ubeq0O
MdI2Z6jjNhri1Bz/i1M11ojnWBFJm7KRZiJOhgmIHGhrbj5qSBQq8NyLPRkXp8/aVEpLj/sSn+Kt
oihrJU0DZBEJNtTIJHESZT2bkA6wnSB9x4V2zwSIBN471Vh+e9gtZg43clrzcpuDhFWs/AsmFcaL
WatldrfYQoBIAp5j6gy7uU219eElT/mWmXnxNKt8JIApv9avNE6tC7tCcis5MaPVQ5KwNw7e1KnB
ozYCecpqF8QMMXBWXHRTK9oQRxgCab6pJ3y2r0w++ZRbrF3wwymNhyyp8dM/1dMM462IwphWbOBb
AMGY2Vf7erxdDGG5TEx5TX7hCwKAKq2bQGXZPmDaMYeApghhq8nZfkF9OfIGsptSLW7JSMn2EhZd
R7kdYL3T2V+E5w8nHNd4lB3QwvsZtAxiXgqqqTj7b9n6LKWznyI6LroZgTEM5IKHNHVl4Mn4DE2B
+CynTjKZ5kCY34WY6uJivzgACO5krvPUf2jEdZAOXaW/nbF0fnytghr3BFVAUT2wq5S3pHI96Anb
FCwm6CxSDzMnV3Rd9SCqERuxz8APB0GkuuaHoa9zWniVDMML6KeRZLWgGTFUnJOrUi5+gUPvauQu
CyX3LAtKveUavdZbC4uIWkZQ1Rc0j6fSW6b3LblZKj7+oEjgkyj/TBR2Phd5XlQUaPnFeNIEdiEZ
PMyejHiHcqitqaEe9FHyIV/QyeM9o1C7wiJypoTvXXlI44WNFG/ZZs2TJ2QFUDBMUhV2NQPU8SoH
VTEEA7CZg4nSCRGO7+jjDbjSz+4w3PyZOgw9IoDQcm6uRYMBOsw69NFkp0xhz4csupZThMnSx+SW
EMNnTlZ0iw1wXcZM5HW79yDtAsl/r8OPhi2JDBhIaVqtFrAIvpCB79WEf0Mgmp/cjG6YxTw6sTg1
o3UDbDblHutqAmfPg4osSJg8Vm770jZwtIqUxoiyzqneG0gLz9wXD7lyo2S4TMWbhEkVCl/gdz9n
J4ruDlcOCJabJQ/kpuXbp1pzeGyQPNtfg2XYlCFzRFOJbX8OWWjUwevprHlrwgOZ07Mmg0ZHHnAd
ZV8/2+5j7ShAJ5iZjcTIl4xROy/jIuNG9Hl6T2x3N8Tyx2vjagm6RcmapNQJH3OyE2XZaFqzIrSp
P/T5x6ThEMgSs2wN1+xxi59owaZOSX7it0FeB9sREWbBI8/K3KBINhCwtoKmRdZg21To6qTYINLl
zIYhHigQMo6a/9FzEnFlKHUGZJkbtDksaKYmZOFgDGa4/GfIPCin3ctszVajTgrXClTz3eef5kBJ
NOZG1tgwGOKnWvd74NrK9ac+SGv/PKxNgMoQA5NaNWSIbzj4rhCe29psOD2wKF81qJ7En0JywOXP
+5N0OwpPXHq9YSAAIpnNDezZEzCVM373H+QcMkBpIBWgF5/MRee1Kx6v6IAOjxzYJr4shnzGU38J
9y1Cb+Ss6H6xF72s9pm6Q7Ie5q7dx5cLMR0MxK5/zxosJ0ovfjlUV0K69I0W0j6QvgP/ff3Bd8xz
mt+SBxay2n49pS0VV/VeSiQ4gTBWLA+KRnqxd1Xj5FEi5Ojv/IM7BnnymPHhtEtv6h7n1V8P9y7j
+A258SOrMMUTG/2URtnkgUwgwhttQw3Qjp9nxgnNqvi/gUjroA8pKI2E37J2mHAVFiTT6S/rhhzn
DgF3viufeQXIs+8SvYtyuLSaVzOYLJbTwX2wu4EvnVe1KU9L3/HxbWMSswmTuehUfsredKAnM9c7
xrDMiK5aOpw5lB0v1VwpfSzJgMq8ozE9xmzyQAxuQ8H8CgkaJ5Tva+xFSbsM7FQvzpl9quOY1r1e
+EbtBrL+gfTvHcXm50SNDn7CFGIh04Pgeci5LAl+k1nWjnwy5p3zDjSm8WVZ8lkUyJJtQUtK2z+s
xOdEumrQJqHL9ODAdhvV8E0LG3knztsSwgjHKlwVnYi4/dgkE1Xj+GFeHOmtrgFOuEv1+oIUfj8X
6/3l0khk5xzQj0OJk/KDMtDoSKXxiCBYvY0aRS2Ok5cii66CbqzS72kFznfVO2Zm6KOWMHz/FIVh
5bcERyEXxuLly1RX7E9R4oT+EGIF2igF17qiHRsSSKzf6DPNmXIW7DI6ObVp+bMYeb6HqxMBq51M
E74I2nkoDZv9TxJ/KhIaA7EySqUrOtcWS3SjarpayoHB8AFIc8kOOGgShukAZtpzdUJ/CIG79TDX
cKSaDuLRNvfIVTz2ELJZ1uz982jl6H8B+FE4N3E0j4dop/pDTYcyzlWNpHOjhJ/V/glVmtf8QAGT
N3GOr65DKIMxs9TK6G+b5omkztoYUHyPVvorcYWG0ilsfO1SdOcAfUljJKEZw8PuviyauufPTNQc
7AVLDxJX04tTneCzgyr1QvGR8+ga0/KGhdUkiYlwmFVq421KS+0YWQ9KjYlndYgE2IkAJL3p9uJ6
UrCXLEoqrT5dSlournvdxtTrdbGYI65Jdcdn/R+W58qTOkHKJJD9QeU4ph12zIGaKc/P88JreNEn
dgcwyw+0pPjssvLpSddBMwPAqsqV8R56BcGpWfxiDECwPgZQslaOzwT1XwAyC0uc++i4WLMhU9yd
6WTyeqTbTpcpwiYOLcgHwIo+XWPIUXKlCQGUxqr271u8tgEKaT+AGZ/z5R6h4tPDywR/9flt6H8I
S0lsYQmJJZoMnKEQVwryZMuQYpkgFWrEG5JfiB8StJCqvYgNQvuUYQwqxcnJrDabN0GfwestRyAN
Sxhy/vpIaJXgwNS7qrb9Oh9FX13+AavRWQcnh+6X3GO5YeDT+mqvR5VYYH2BBay54G1Y6ANWF6cS
15mHbWuv+lZK9DIHPPQu6EIL5mS9lNLqAyPZi3YwuXJAZVzGGIMhbbmpjbVsyn79WWyw+4n/Wm1y
KlhI3pnJ8RA17OTcOrI1wke0rLYZK7r2WJentlvJzguK4clPNI97owgXgG9dDH9R1vyqUc1igxsV
PjBVTS4ZDORIyxjFDYGXhATju7CvrcVVZvDP1Awi9IhX24jSo4jYiyOrfnC4uh63jWXrL5wcnns0
8bbWuJFtN0p0mMpc/YkHhmB3qGyB/6gQ6C3zuOrp3UzmShmNxgJyGgr25vg/zWlq8B7kTgA5tmDr
Qp1r8wNGN7f0KkwR9zXX6gNhTrDY47ARg7p3lIJ/eiL35A1mSoz68ekicffEvaoavbHN08P6VaUo
8Ob/yKVp1Crh6eb+kXSUYnrqzKGsUhDHwo/xw81tJweTrxIlRZpNSBc7HaUlUzlVzcvzijZH4nsH
aGKV9BbSxSOn6s2IVWaxOrMB+ItEHHDDrFOhfXjATlM4JVYW9WujczZUIai6qUYtofeBjOuVzxow
W9EslK3xLdKkHi8quwa+U0/H+366IqObGm9qQzeoxsjYmRqzZRvMBPbp9muOXSe/aI9CMt7lR5GM
X/klqRI2mDtRPVPFeid1NmpDHr7OoG/VT9JncRaobbPdDtU4tf9lTQoYxG6xO2KAfba7WYpvQm0c
N9r9T8+O40bDY85riR7LwByiseG1RJdheK4Nh/N7AxHwErX7TgBx0RRPoSlN9mHA/rYxHO8s728J
vskMzoCGQe+fyua0Pot3HytoPTNrcvFIcgkMuUEJ4fFUa/Y7jcuL0116RXP2qxHEUBJbf4hHKMfJ
Pgo5TbGQKZypoesm7vJ5Z8Ms7wQ1TmLIE7O7ydnCXaFXAtYJJX4/nfbfxJ9+6b08aN6tkc0qrMQK
jXWA2nx0wI0TpVhsJ8KnxHfpHG7bjGOI5EVec7tnAzHb4gqi46yO1RKLxU8CW00nX/JzA85ILF0n
mtRoowE6+CAsURcuZ+nYWWTjgVCIkYS8yCY03J5ugxgrH6oMVv89q+ECLtO+18fMiMnfP26x+axX
DNIoU3A05Ude+KGo/q7tIlRGrssTSfEErfAindCpM2eCr8R1ITNPISEuktfkvqe/chgDChn79YXC
g0smYt5/XQchPVu88PkJs/e3JA83HcMtEyJd9mS5zxe67wSIE9pr8sWmXePVYux/7IXqLqm/Xc7Z
LL0AX178zvEbLtfMD6KrEDDbk0KnfvyDgZZ8PEPFF7NFZBE0r+owlnJ5fktjPcWLxKHUGwVnTLU9
FtNzZ2hJhaAA5ojK6arwpRnLnWwS60DLb9o9bySHoedQ1jTWbDJ+nnY6Yavv+s6BE5Q5SnfXq+Yo
xRtew1ob3OrK7OtL7nh5XPKI5sIX7qQgw7J7Qit5nM274CzCXHfx0WcxZUYUfmhWE3lPN4uCnoth
byUqY+bCuvE03PD93Z1ZfaWpFSGDGDrq+D1pHKi23cZGJP5igAdIVQzNBqlWXySpuT7O4haa1T55
uhRzVbp7SV/CjWufcujnR9qn1CMjMfHBFVrisFi1Evx2iDmDWSBIY9GzK9kdbsQPBpi/vJPX8B2C
qOQ5yvv4klaC/IB4dRr4hKZhCtMXkakbcvwZiiuWwZxgYqqpPoeZonjV54XfaPojdEZuQ+ZoHGbw
glZj8hyBBpF2lk0Kk4pz2q/2Jk3OprHzlNL1JpUiL67jUPy9qkCqjDfzO1iJWg29avWV8A0EeRar
GTIntcZzaWvMviBgaAHguMnCK+D0yg2lVnTeyjMuZyMYkJGZyJGLu6yhesnWBG3JSORXubL7mvSa
mDFS+TjLPmhqPZawjXWl7kchyxdakYm7baL7Mr/epmbdt4B9E1R2lOL95lIZKWZHhFaslPK5ftWd
extWwY6oQEL423wVwE4VcqHT7DRisjn+wuIqnVV9k9U+fa+h9jXjUMBcydl/OVrhHjF1pEA9YNqH
WrbsHCsDtvnYCdS3b1pQKrlSeVBBjSSCctDZhwerb4azbreQRy84WpX3tgQC82A9zhBz/f6anLP9
84Lg87RRc9vPi5KaNRFrHcsk/0+gmYk+hzv0M11lzkQPtRL4IvwKgfjXl5N6GBl/SEK9KfZXf03T
8wuKBmPFKYF6BeOyXgA9mH9WYrcF3HunSpWJGAoBjvVzvplUk2Sww6LBQmUm+X2tdUrhDIBTYxRq
l2pR87YYE5pQsvif5DMuX6ayv5OcCs3JAWJ7vfLlR/MIOrN+m3A/5B/mYDNoMcWTFaHpmhIfhY+E
kclaz3tbvwF0Sejjx0uKgyDSTf56+HE4AuP/jg5v96F78kxs0P66UIqoRvbCznx7HdsOKfkKB4YE
NDMpCLxJ3DFpHj+cZFVOz/RTvI1/AYDqh1ixHIBgFcMshUIUqxux6Q0TNmBqFWgtBBArRA/BVYF9
tDkIQ3iGkcGbZ54nMPOABrrlEDXpiyzJmV+wZ9zoyvR15GoFgKndKP0ZsUgIh+spGDYXplFHr1Vo
xZ9IZcTqPHSuaa4+5GAmdmEdbUIa5mbpUThojkERXVDjtyD9GqNkP6y8sLArgKX/eKew/xMEZJRo
5i2kVFrUn45rZRdAGt79Fld6lwl9Sl3NcMr4CC/yh6cb72YVyfpFTXRxnjAH0A0dYANNFiV/w1w9
EwkDHnByG2NO8QLoJBoSNBHEcdOPbpS1/wXhOjBl9pdBVtzsPKgdhWX8hlG0Uazyr+jXb2YFBGwB
5ugS5P2OS1pG+SSyax62kufE6NFQbGyLgoOFn18rR42GmepmGoaJQdymxXUqvlvac3OC7yTtO0AN
Os2itWtI7qrVmoTXVM5ccD0I0o63a46u8NO6Sr7by0+NFpgO6k1Y4GqYw5zXOuKi2FiPijzYFNS9
0VHC2/ocnmudy4JFTbheuFvRvN/2yJnLcEGPruJSFQTzmg7H5B7lLtd9JgDZxaWK4nEc+dgX52Me
Zd5Y/Q5AIAZLuZZsN5rCc2D1Ma3Buzylj1EP4cdOGt8eVPKu5x1CWGuLWvbt3ik1hvKjuVVqvz07
9RQc7jJsZneKUk5TfQtS5yWvK6MaqDYcTHqNLTC1zRNSvcMdlqziV7CpdJdqTRtPiqp2UkzN6URg
LPJ1EDq75VEauumnp/EicxDj2JymacpQ41kyUdXeq/DHUdSgKamNP5ISWpmR9ajfGW3lg0HtN4Tl
x1EVTejYSGesjaJ6kRklp6RFno6IZrfowaSWRqkinx8RK1A/RIaEzqpXK6+uzln3R926p1D57T7S
P9vI97d5pbXoS+DOHyyDARNqF7qkSGlzl011K2h3ZudxH5RPFjzTqbpM6hkrhJlRVE+UCpS5xmwT
rdgO4SvMZ4vWiGbxL+ggIrnqYT7Qxd5tmxh2tImOM5wCskmPUil66rbI4Vyhuc6JtcVmptt6o4mM
liVZMeqoL4LdsJN2jtSKcYIQezryrNRcedeeLQvlkLeCjxAKzbTUcbV8rHUgRwqxe3h5/96JpzPK
+h6k+SEzKVV5EiWyz9dMNFz9oQMrG5og5QPPAqc9ck86e/wSgxs7tz4koOEfYw7wX307ZWhABgsx
cwhPBxE6B4uVxCQLySeCXEjHV/DyxanwHG0M4VvsOoPgF3ZgsDZA0FLOIXa4QAVmeVdxeyV8kvr7
q6PcVOWyQ5taDsBBVk3ifHG3wefw9vtigSRAU4Q2Cuc9vDQLDXkqHgUY93wqLdGkF3uCqva07/kp
F6s98YH5neFvursyY+e58l5e27x4yWzdIFYvEqDbDsnvRZUeHzEPn4yCLfoxotPU46yFbtkZdGch
QbZkdqSHQUxQnN7hv6jTbvM/1HYsThrXdenOPk0k80s0mcq+lpE4uJS9b/IywEECBYwJ2MUAUwsn
v/G0hY6HEitUIh3QThsNd+p4Hz7CENPNUqdHCo7njH2JuEc6qxxbN7Vkq19yGEMP7ZEStJSrl/CS
wBOTcutXjc+0RKwZ4pgXiFTwsOpCt52oLkHgkkY0MiKUwgzdtEbSXkbdLQwgkhmUTkywFVc1zmfU
lzetMM7v04DjqhRKqxbcEXAKOhO59IVuGa4IvzlDj2yPFg0Z2FnjMv+nb8CUR3T+7n1io6wCtQAu
N/xurSbYMbl1DoVupaboWtEGPYZvJWstnJ1h5jJ59aYE8qqjiDdjg0qHxWzlYodR4mcij1THkau8
fZ0Zl+SqYgzksLs9rxL4pALuyJME2wiYWoWzt59iy5JmR+i4DSW7Ei4pl+kRct2/MHby+3chK1x2
b/BGuX7YeUycIZL3B9mr+lOUyt6IyoLtafVTgTevotXh7SsrpE6wdGsbq1KpjwrImPaZETUYnyw6
LgH0eCXfc0IPquF6pImiERudYXALN10KQKW+if5Q8L9t+dMn+oIQk4hBkYyapZ/+ua4JXyjeFzgd
YJYM6Qhn5I9bNsUZETNbQoc6S36s62Yi1asswMWl13yNcM31UJ598Epi3mYEhGRdY/icb9nhCa/A
MPDYwAQFokNoyyrzaXR7qRiujjKKk0rMjb5Lv0HqFfsLngTg1Fx2zKK6MhOcWZf5XBB05mtdVj2R
qt2pAxSXw7dmwxee/eHCbHEYg1uqjoBQmQAYVt5gAgoR+36bK9SF2q2sAW8CvzAxmnsXKdqGt/zo
RzvC9sQ6SzTR3VqcMTkSTpfXhcHCzZ7UW9lsDEmbgOvAZRv548Hb6XsdfI8+LGWCSiP2gKxYU1A5
0SH33S0PGT/0hZ5EDsYc782gX5CBVXciAtUMNHV0XKlbQtVd+WbMHUMrvKduV/a+6STtnyW0N+nT
+3u/lilSFCTnSK+qTWhSHZLJ7fEB3vJKUuMps552zmoCr6s6a+LnqcZjWJ7rwyfNNUwtSVEPu+EX
/OACxqn7Y/k+yQQZ+BW7SoImlGuF69jG3nY6JjNy2jzVau39pWxGhgL2gslny5QpfLrvFxYzVquC
fESCRuKELUT9P5AdARC9PCKVg1eSIXgJjoqb7B9K2fxWcBfK84ytOdzAR3V48ayiMeF34kfX0Yw+
VaP28Xk32z6h0I2rblhU7o67Jb7EhLEtHk7xiiT5d6NIUML9ET43GPzpDRg12195UXd12vqqtsKo
cT2duarMIrFeQbLmIAH8hJhcb5cYcVMB9ucK1dawSgk0ErKtbAtqUsSy5tC3eHpQmG2+bghuYoVp
pxRxdoOznH2raId1TA+KD6H8Gntkagf7hmgWcZNG3t1yxG5ZIPixyUJCS70KDLMC1zM6Oro0FG6I
3UKtS8iwPZL34/Y/2PmDmJlACIwK7PllH4hvCMDKpQHpJ81t4ChzK58mOu1ZelPDVi6Pi/ijuABk
bSDYA3vpD3+fpdfPfdJmxL+NLHBFNF+2bbqruB/Q4xGovDXVdYrNhL5Ut/CDoVL/YqFziJLo8ZJD
fjtdYZwtuPdwmCBcwlXqS08x2Za5JrKF+CsH/sr3gJ3GO6jk72VX4oZZKo0Spf0WDzN10/Xt8TDH
/LIltW0B99E9l5PMWz5+JOQLiJrcCBoen1NEH52iLbg1FILgQaXtyuKsTGdf5txqGn8GlAVAH7Uo
8B6eig/Qxvmj7wtexkI10/KLWRhpskHl0NKG29ZnMOAFBw8FyieWXd1pakf3VFEKkNva7GF77dkv
b/DV7hGzKQZe30AwnU5W+pU/b27Sunp2eq3F34OUo43Ya8Tpkmk8b8Rx2ccFJZXCpwxkay4PeoLB
/YZW96UZrp6nLjjwSrAhR60bVr75EwU8QCTlYLFqMKp8oCbWOMZty7jsbddFsJtUEnbYL2TswAlM
LOACJycBNU2s7MN1cpek2EV4BhZZog2WpSq8vHj3dVUdSQK1hkZ+KtJcx8otxsuwWRtIJrTEzpJL
mhyfaGdqV3E0mB+5/ea7bPnjxZ4qV6/zJdngADKq+3A9lGbU9VK+hLrgwHaTwIQtcWgYYr9tqB2a
3Veuoxa0rx0TRMQ5Xl8pa9yA5BzJilkwKNWIvq8F+RCSHSJszqtP/TmhUb2xnwFTVSTD7EU7d0go
O057sU9TQ4LTmVQzIybXLn2elqJAX5hyJnNwbHUj6++p7sL8C6egstnBPTSa3+M2U9sh/Bk/ozcs
MheXPeyTt1iEtLZkyUF8fIkNFNkC9JcpcQI9I86v5kGnXx/ftZtiyDlCza+ODVqNrwL4V39jp/lB
i8rxTJmo+BlI9+2q5v/Dk5L84r8lJlxgPUCWMOz/MFxIGTAiJWzPMosHdh4EhDgA0+4WVJprx6O+
Uuomwal7WoIV5Fc0cL1gXZ2FXt/aYQGt+VbG3orq9PaUl6lKc7bKzZPc3+F7hL4Omcc6tFGUn57H
Ou1aFpGg9BWJeHfc+wZThFxDqOAfIyUY1bzdWzDN1+oKAG00ru44PT0T/fdda2bauNYE7C6f/p2G
YkVMpY5ymE62sCEpUuBcscxY5bHNVeNgjPh8wr8FtR68I0ZN0rwg7km358iUlGRFJh3Bk6a02SjZ
jANCKWgyxwgUcF9PZxCoSuHo6juQkhB+/h0d7fEE6+jCXD78ZhqIO7nZTHOEWKFT2XPNXpfr1W4X
UOfQieZVaitj/9MgCRoTonDSElYh2LCjj4U3snzxc0XDlglU52NGNRFzSXa2zNOQLh+oAMU+XOj1
0CJQmkKJ8sJNDsZXY/K7SZLOs5xVtnPM4RR2kn5L27KbZo6L6pWNvGmx+PAPQwJocNKP3FQdgkwk
ieissHwQPyVn6aF/vq/jc2XnWTqzTfa/V6iaf0/J9/8JE7lcxqtAdIjxXOoHndpoHMpZOVT2bCHs
8+CNo5xL44WGhEJgflh9PrOm08ygC9rbxe7100U1JtIv00MCKT5bSUzyEWlsR/Yk/8cecdIlTCGj
KAincfKyBrEMZAfubXxJ9b50BUD4/m/0Ycyb9SEsIxWaHZPxX0nuxcHLy50bdQc2+rxW9UVePyCt
SYsPqmG5sk/eQvB1t/9PN/aySYK3a0okKxKx9A0cxG1vGKZfWnyAs47rGQFTe9rq+cp9xL4HrdyB
BrLiCEhtEdZ8UJpMJuuJwvzKtoQH29+9+U6dCf7UuYVIG9ydVaCm7cOgMRFjdlr/VbE8AjG596FH
jMznMjIhCMUWLEHagDyM7X8JjB/FIBSpTeHPi1WHbC3Pv1Oh8UqkxlkQ2r3ZgMhqcHAmPKTqNmVX
S+kHUoEMRK0bIDGLv1DN0kJRslILR3Nddxs6myZQ3Dp6sTbXSnl4b4mCtbNWJJuek29jQLq43/27
OG75wER7k9Kga1v799wKS6XNPuGUqGgmiOh/U/0VEZiFR8t3Fx0NN2ms610bRghIW+CPO9pfm5Mi
4Fsq+ert0l0n8IiCXx2Sh2KRMJerGGbVXvCPr8ngxTAHHZQr5tVwCUTgHEgCPBtFNjBmccBzMDfa
6RIA9QcxTRx6dRPBcM6rAUnPyXMl7Ef4nOXH+1B0BUhZnvKOv0rJ6mnM2/9AdDHoDraCRfuPh5Be
FvIZ89nOtE6sXW2iKi49IvtzKa9fv/l8XRGb386dKrSerr7xBpSzkFw6YN2xWq9r8wrptCMZNSCe
sa7DVQXTtrZprwbXJ3BuIGM1MgNls2/jyF9/++XQfEHyslM+RywBBv6FBp8PO63XsKpaCQ/AEUzo
5l3NZJJb4OqZv8mAvrKACUKRM8cjTTHenULf0M/gz9AgsMXPiN/Ki+L7j1Xvao9gYUUI5CYih517
0WASSg87T6lE4scylvTXBe226oN+Vo1rwwMXu+s8w+STW9ZKuY33rsrNjZ+rheZ/k9LqO/mvmY3u
vXgoDX/T7Lq/ZJr8ue2P54Mu3/8DeUcmgbLAx8WVc8E0kxh1SnQ5Fh6Tj8QA9ngF0R8RrfIyvI6s
2A9qLIRzil9pKzQcSLYy4auz7CFgNCnIkwBiK0DuuaPVFPTS5BwXyj8R5l9m4u8uuiDz8LpicQ9D
+NzqZTdkWUV+zM5nMr1hjOcs6/jzXlfiQtnCtWI6yao02heuILoNLgnar1l+8W/XsTuFbCVL4xbk
5ih1ama6JFukExpYlgz2pKbEE+chObIU/HGSWOYh9iVdvwncUIc6Rg5ohMCWavmfi0SPEsJkCwN1
mQFtuZS5cjHf2MuvaoPcviz4FZ4SgLGZvz8JmEcvOSRDn85t9n+W4S1J6TC2/SRsHjHa48uxc8IH
teDWzBj71Ox3bi97xFMAxdudCxVLv23yUKRgzwR0+fjCSy68EzObI50nT0BvZmXpBPls1QKvAsVJ
PPDowd5R4cgPj7e5GMvPS/iZdw/gNov2YcFqOT41yiZoZzRA5X66UcPEzdvCaiYT6Wc5gSTrWk/t
ZW17JaWz/Dc1XeTUGUpjfCT8f8VxFpRFoDxBVOc3ineoaE8ixQJfYApUMfpppQHUYhUATpsRLp8k
L5Jk79aO39xkxfK6YiTf/VMsoNOZFi3ikoSxrGw4Pw3gBl0Ue6bqXMQ72AO5VNplzg+kv5BgKyHA
rQhhbPtoT63ZVHf3pVlOAwyEZwkHCsoDzJDvRxVzJwfQq/kcZVP54/tRNoTWdsf74VoR4tUlUtFz
pLZNNtkvl1QG2gkT9hfvrRMYY/nCZMi/YOQO9bRKHRzFq13QtfSXCh5YNUpKoAGiEqmHG0kDljcb
ti+pMSWjBQeDC/DrAas1HBHvyGogL+3vW8X/c7Zz7I3wy3i2747GYuX3PqRx8oXo0XTP5uewmIsO
s584Av3O+HbmEYJlpg81lCHuR5tXaNx/af6VpxO6eeYnKvmqGuCgulI6g0PprTAfWUvbzW4K8bTH
5Kq9XFPI9+G2N9VTl1A1RHkKlDvBIS06cEGLbL6QOYeBe4fBj9zcqqAeha3K0SpmJVq7phmWQxYn
vutS8BWeOjRQmMtD/6cJLQ9J4ilyy1jyjvSEvswmifNY5b3Xe6ZPp/xKb0Nr+0qOQNhvIZK8Wq+F
fOLVeyO9QId/OiLpwjsx+kQYWVOezCXqpOKnhzRPgeHmEsL4lrpjBirVKZwL9EvbxxZq1PkyYcNA
ijxnw7zNdUzqOZl9Mrgy7XxorLc35qxY2o9JP7obkee5V1ZA0OA2ORT1C2pwCfRKUjCi6XmoTAA7
LdHTIT84qzqMiHIBrieCCG/3XEPopNbqq5Xu0sG2932IXIYjC5r6nJN56vOum6nsYv1SOG/it5sY
Ff7LOSc3H7ATAYDDS1CoOwV6vmPode1LfWzP151f7jkf+I/8DzLjgiHaH/F1z1vr8Sb0LDwNgoQj
yQOBY2EgVUerUsrSGqteaxtYkPZ9DUKCrgfcXL0fydKBeftOym2ZLRpbjSHiqYQWWbET2jBG78ip
A45jeWvUuR9pKxpyA0hJyjxqDJjseNrCACKlEFh8Tbgmj05w1g2zyZHJjHphhQ7ctvC0BNR7oOZR
DTS5NP6cjZ+aXqjiynhCGLLMlf7fOij8UkoXcqGcM8RVHrILQrjlN/tc+nukflJ9ji/KXtA5PhAV
M/VZCFXD3rtPni902XrzK5erqMPmKZoccYZfeL7P/h0lI4pIMWUuUc3KJlHX+nT1MZNqVRtqieET
9uh24QAmaU/bmttcrW6vCnjBcCDmZxO75YtkiBK7/HhltA8z3dQiNRyEbDd68E3D8zR0U8cL5gCD
Yw1NOk6o5pIE1CuZzw2y9OfL9ZMansx3mO/w9DdH6Kzdnf3QWn3nukUcwJDZiziom8mk4LPChhd0
nUdkwYfGMVCfkfk7zRDnFcmh1fhGx/yuoltFNToSXJQaQRYiujCCPyFSt1MuyqP7ndCodjyamjF3
XK4VKMdWjB3sDrdkKayN/otMPihVKfDEMU1HNEIMS0/Bw65rHhbST42czX+bLYp3u7qo0SGEQ0dz
VEZ3+gjSzQVl+GdqNo1Omy0CxAvyhN+E3MRk2899NXTbKcbN4p2YmExw/Ofaq3M7hLlQGoiENIvx
q1JfQTTd4Q/abRWpfMRyczQk/dmK8tgr9ZvXdcGTTuAzG8L2A8lCdFQCkaic3CN/SHJapcA/QDny
uf5XVIz1SmzTJ37atwLTkgJsdu0ggbk94FvvbJsieJV/Zq8dS+2nzt2d9LCpv+oNsMhhoMFVHvuz
8Sj4J5Rhy45Pif/MkcQW+45c3Fna5Gq0Y7ONlcpuPOuEUG0bQlvt3QfIOOvKrmevb//pPrVF9BjM
WqZK+ydTzf7cMLfhiJKWWUVaa/cQ1XE3bX7MFlKNiWaCHR2o7GSJPV71O2M/vMGDQb/uP3ZuVUav
VnSMuVtrgn3yhLx5K8WUte46C3B2ObaH0ydQMn0XYxisSa2fiRCNWtU7+xAUPioqkfdPMVTY287H
tSwxb3PJsbCfRn01S6djPVGLaqSdqz+qKPQ0PzXPj20MKc0j5bnewuJ4qH05unTfvjyyWyW+Gp+r
DnBWijpS/kcK78ssQQOvKaFbebppxLJUHUdPp66OWgg45OJYEdoICZVSnUbT1H/+CRUgjdTZYOD5
An1/6ifYYtHF3I+A+OP5JRnlig57lTkVYQVenBDlTu6gf4W4QaZvvGYHi9tDwJQUNq/qUQB8dxre
Rsfz9oDiA3OyTL9U9rw14NDpvDSVo+YKfBu94+TcsT+vbvh7ez3fb7CcocKzC3/6DD2vR3H2znnY
g1rd5ESOGXiusqW+5SXqwgc6iXRDqoMQe+9Gor+A6NyBVtB0zvKf+nNrw8ve/oxWps7mZm8UCbg9
hGIm3u4MDwfXdpp70pibM5bTqULZdkOEQ35LaY1gXtAdSzKHC4V+DGLS6BxiNvaWetQu4jU+SfPF
o1D8NqbMB6cnwLTkWhwtXQae/gwlVNL6wudNo4CpLNlcBwpV2NFvM7Uim0ekaQALNlqBWuy2OJJU
juTc1cL/dWXqRIAMbuYSBXCtkz4cDMoySZZUiJ6hHNrSaRPqWoiIMSmzJ5rQXJwynE25li+ovIjb
UBnIbPfSi/OsTX7BRPRJe9aJwhS8X64tlV82P70twuxYlGhepbPx/OLgxbSY8uWbzZM7Rh/p6rXV
FxZKRke/sl1pRsmdeU6IlSi/hwk33DapB/mQHDV7IZKkFoXlrw3Jvnsx93Y0fbhXUN6zWtzIIpc/
rGjy/GzJvAq4CHOf2GYxUE3Vby3DwGU/5R+x6T098/pmHUmFpmkPYbfxwD0Df5VKFQa6XjlLomSv
O8jDoQz/O7HNsjNhcxIm/1xCwLo3QbnWAti8J50YmGp8mnsBFBBWGJAGkWF2VWp2lMwPLJSEufNG
/gs6pg2yP0iZF+Pi6CPACacc1Uo8y3beC1Nd9+C/jkLkV6yrXp+Qx7bOU/NZGvangfEDXTXfy8c2
UaESz3dZGQh9OY/slKVmdjk7dnAzrx6+9UOKBAydEq/q1iIo9aFlQmd+1nBQFEiAA0RiwuxkfEP2
HReR/dYEAlaEaQTID9alrLKGQJeOVpRAoDsRQA4ayPz9AycG8BONUt27b9eLpHe8xJbZRz9jwdNT
r+0sYgShVfY/65fjYna86CcalDaLrAVBVYsOA6JdRKV2cN260m4qaCEu5srXrbFk9zY7DFxILqFC
YthquSwnqtPlFzlI/V1GgPlOKLQbLvC1lahb6SeQjHWCO67DSRSiCjMSm3H+WB+w7OqeFB3cq7zS
LktiMQMAGGYdePArn1jYnas9Hh4K0zreuHnsK8zSKMATinccldESSupe6SR/YuuvDHOMVyMcHHDy
l6dnm9Xkv4NH/mndoKV0JPITsDwcFhW31z0lfR2sbG4rKls/Zvg4mCWoZ3YROO1eOqrjj+TEb0Kf
gmRGWf30HpLDVfZibKL3YZLi/DTtORUU+QyC6jUL8V02ehrmZ2cgkjEJ575YW+KJdvD5wFXhuF6e
2EdGx+pwzKZjB1Y0LNyY70zOjrMa4M4PqALovY/+Re2KA+w4O08XNMUnEz5BfoFDKtPKW/IYq4Dv
gMyccVwblpaK72MNFD9QCAFBZKbHNgyu8+Uz8h6IezqsRiFLLVsvlL/Hr7G7rEK0cGbgtvIwEWdq
cAed7qbRIK746iYze0Iqww9xCejI96XElWL9Ju0jBAP3/ooobpPrkvuL57Q2pnYvRI/cy1Sbwnnm
OuTVAy8Nkn10t/NkZvKXHspIOsR+GWJLOExHLYis4QrnHw5ZNUz6cgLZPBSkouqWebACRygkhVnQ
Z8YFH37/u9omtt4go0VssGzIFHnYfOEOlRlbhZS625S98rUVgUbFZhmiCPn1W/3YxgVwlaDo4+hf
bL6Vv3ugmZVzF9+AMApuWQqRVDOByBIZ/mlVk43NcOwZ6UguTMl+m16z2xsbiKbLXpTmcD3LyYJR
w3EM7xzPYyMLPzawVi1rU1GyO2OGyzecIyrl5gt30YyUdlKGkrj0hGuyJYJPwtdTWqnWAKdnk5OH
VVpEChLm4UWv97l9cN6L6qHQcdcfn+vqgsZFj14gx3X383dtAS8mZg++0urdNIlfT/eIVNgWx1Is
xOocpvgG2dYSTRaGPBWUrG12KXByaka+JWfB8C937mH9OKHlR+UXFmmu/xIOITp/S2O1TinuenVn
5B11RiKWKIy2/V7h0J3Cntetq/nqoCnXQdUhJOnQUesEsrSKqvgKW6fDO8aXI1NokEutMNBpQ10y
0+uF9nkHJeSeI+MyMjvud4pp9m9FlT4LC3sFd6Zx+YtmFxA7Iz1dyUmLOn2BDblBUX8uWFFhHMwC
JzeBqfEq/cU6LfWtMfcg/UhQAMGjk7bOMj/b5z+UVIw0T070Bjg7BmWWSx6LsbUQPAhBeLh898N1
tq8Xk+ZBWaXWZNL1grg4LyGNRFrbUEoConzjx2Zy4TqJjOuReLk3KagDFX7ScRQxD/uyoO//izre
TY0cU6/i0BmqvF4UItmdFasTj/D3Z2g1OUSRjQU0zzUWphhSsJpKl0/PqiB9QMTl7bzyWgSCzZni
JIDOdBHVOkbHjMPoYmW5ceuhtOQfSRLt8AQRSzsREf84p7EuURwGqCcX/V97ytZspLvXn9yP5IGT
RqGikTdVijreMpplYXiyuee9lfvvXYfIJgHKjXgBw0OpzuBKnet6IzPfRA5GTphXwVJt5Af4ilZh
IGo1l+wCzoFuYyIoUuMeF/qgpByZOWuDrLSucC8uT/PRscDYAqBJhGaIYN4AdqoI92yrdHMRQTmd
z4uFjuPY2L/9vhb6i5S3Dr07mhS+r2ASEX76SObXkEldKICrgo41KYMDmBgewqXuSs27kaA6JM7+
QaEa39XXKZ8IRv14zofXDqDt74TeiiD7wuQcRPYFQkIMzQa5karBveOcARn9/G8fwtGLsz0CajGS
kP5q2SxesPZIW8aolyC9c6WjHjDuHAJnM32BxsOL2/lbjqqiF0T/ngbnctcejVF2c+OFRsKlwy8F
nc3Ttq+n1+ePc8tvyAPjHFy3P037RiLpQgjrxyyj5RUFv0BgtlAAtsmsx8o4ro7OnpBtxO98ZjED
jILCAfro5UeOPjcZ8plqffHq1dt1B3Y3h/YL1uqnIbKXpUTSQ8j8mVH2kTwp1cL60zG36azV4Aoo
8CvaK+JJm/UkZ7T4p2m8OaOWGn0b72UAby0d5X0wXLeEIuGvUcLGaBAFQxFMwTc4mI6uuVd39S/d
2zcdxrUU5TAxcZFSF9SPSsAjcFmICNnfqV4fAwRpxd9CpNPven/DmrkhJQz+EDIgeP7tTgAhcQjy
oIZ7S1CWOTaAzE4U4/Jjefr54T5EXAmJF/HiS94cb0TdpwjJXU7zpCbE7YDebTbLjWzURZIqdSF2
TSL/4q687djA6mHhPVWE/e5foinOHL/NKEWQ7ghshDB7RHsrHhRXDMO8iSjO/iTl17WATsoxhR6W
liWjExI6ClZndeBl2MiCUKy63Onlr+Qej/bebktQzxsTUILAKjO0CkShbpjix2OCfmA0uAHxFn35
TJsJCXw1Ru0XHRSUIoYdg5NNNX9aS5d5zL07DrrRNHmfQouonTxjqcgli6w95jYqAAK0XplSypdq
CrIs4STf7FDDyQAwZ2SgJkUrESHeQ6a23P6hnccfAgZThf2IH4s2ydKkhIh6sCFKTjTSJDMvz1wS
ZPubRfYPtXrSUBB9epoEANcCbTSyKNp/qk9F1ulIaDlYYoak+N5ACmOTAlJR6jdaT5+7pWtEwhhs
E4/VZCIBJlTUfeFGI3o+Y54kToCk7d9U3jUZSyFvGYA4PrKTxYcygl8kqhKWaFNHG4VB1DoNb2WF
B7Vn0jItQCpMiO8BwrZwqGpTWZYdC91JYW46O4uqMRmkjMqJqzwPC15g+QVagGJkD34rylXgttGF
OaW3KEYMB1q3+9iJMrRpgGFg+ksWZ+l0Zh4Z89uHQfw6yQX1fV3WTvMGdhhRnGAk7xsxmm2uWo5I
AHDFSS58BnjYg4WJ+p7kMW9VKZ3rILKfqS2zlOFkvdcgJD6GcfcgnLF+p1g9l6gzm3Vd7IBQarIG
Uw9cXk2d9XNT69A5/jHd2oXMTKsqnowwdL3ZFB5CdL5XPE3qgRmyGWqv6At2zCgCw6lbxLTF76zj
du+bq7E3WkhGDrgBVXyT/UUDlH3fL2ushU59QzW2ap6tTvdoWB9NgIAYkiNyf7Nd8V2TYEKIviem
0XyaihdhESifuLc/7GxTWCtzC+LzoKTyZfeQs2Mu1Q+TTxfSS0bxHav2E3Bk+rYLR+uLAIsjpC+0
n+golaz2BPbJ1vDO8LNwrylCWdWGqtZLKYC/Wdxi1vYuhHpNiSzTafNKHlNTpNR36nDh/AyiXuPq
wZlOCMSjE22qKmCqQEj70usac207S6QjvAX4NZkInTAECPQDDrPTZBE7tjlSe3IaonInS04/u6w3
2lDzv6hRjKwutEfYiPxtPYQkzwYulVNWRJalqa17IrzMcvwMwBeb78NlEE2dKhyG/M+oxKr9VMW/
eOrvv2hhrncwCJZ8WsXGlJ3hcFRMmbZyVMAZlNPqVYXqDV2PGS1uVSD2iT7ggyYe2k86bq8nVh7k
uiWRmCrJazcaOqhUX9FfsiQ0OK2tApY9z5S9u8hwGz+0bLARAuRFJwTnyN0Jl4HMGvi8Ycco/DOr
yIVKD/agvTUOzaJfiig0xcZMIBjNt6UtnSzlG+SrMVmSZDqYZux56ucMjzB6GYUYmZz+OZUqEqeU
tsxCAe6y3AjRxJTwwnQjY5uQ2c/Udvet8Y1IrZDQL967NZe9PCKizTofFfk/vC62r5bLN+vKODPz
2Sk20J2KZYgeWMh/lJSdkhkpHwcfGBlEsRmv71IDZ5vXF3NUlJLnzwg6n3QLwmDPl4eZYogi+JAn
0KlB57eV5w1KF0AEa+NN6QtT9U8y6D+M0j/UAhQU/s4A8ol1fQ/6layFfcAzPwrLsEU8dec0fe01
eXjVVnD/FQzVX+Q/O7vpG6JwXyOJxZZa5/1AmMqFQ3I6wGnbStXpNhsKwWZSMVbEaDkgqDBYx3/9
SH3wxePgkc2p950kWV4NLHrH4dE7tgndqAmxkyQUvuHezTCXt1HzxwfBR2OA9EbrMQkfnnF7bMJO
HNFOVQDKvoNqLVHAPAnh2FhKM1mvhFwEZwJEY7+GnR5ryxItP5eQxxeEghBXZOFeEC4Zr6XUN64O
VNjPYHJq8efEt6NSJd5cfRKrVMvFJkQeG2aJ9DKzHE2KwNJSZ6+kxtFnJnBLKYJIX+v/LhQ4Bp+m
vSFs3P2hDSvrhhHNGdjtufFLlIH4QWw2YZQRnXs0Yv7IRaqN7yNsi89VOI5uqIWEUvhiiCQLGLGY
RtT+BKbuO6WsT0Ov7e9CWlroVvCx2zPNv+xlm6Ei1NdDOh8PJi/EbjWimg25il/4k/bumc4z6NM5
NDJVx8DNA4b3nJ1Dp0OjmK05bps1uO8H4tpNfOX8Dzybz7j1YLpF4eSrdWuN4rlYxVD454bmTTek
K1d6wqqyukWg0qWP0ssjerbyNu+jLQNNGas7AfeNwOT4JyWkJikmSGnVAec79yCnJuBN4SB32vDX
zVbrZTkr8S1UQjAzZjvs+q53Ll9m7jp2oF3HQccF46glRPskYGJ33bewr5Jp6E2rCojXTE3dihLH
vVKFTTPyYAhUYHfCWZ+ObEs7FO19DMIVSgzbt0jT0i/Ox9DYKUVxbwcbH33dSqT/hg0pdZgaKJH9
lxGlPJbopXiSEsVEXw7O6F4K4FSu7QDs2SwIB5fKjoHnvfYFhh5EIJHlikFXPZwt/heCwRf9pArp
vwfGPlSjQbypumDI2elbJ+lxVabLBh9ZA2xVo0B7MHGhzv66EIYxdvy7hLFA3jpsLH5WK4ubu3ZS
bxFlbd11EgjyMahUHsByHUJ1bX8ij1c7Dy1XWv/2KJykh9fMZaCO9KlOJBAH6N+x5S2VBqRHGxFI
t7ySTePfFAc48aU4NsJKrrin2n1Zc0PXd+p/f+2jtJuFJeZjbBJwU/znCWdM6y2PjDZcOl9RZPaK
kdNyCEWIPrMzvoi1fyfIZEDRQfYn99XOC2msyM0hSFrRufMhc5Lux/+aRLMoa4/8W58i2Si0yzYT
E7iAfa3qHPfzRhha4zdXRyc/whDaXFEdEQPI710XtxSwddfrGLJpG6WNJlY8y4sIXVPsJpY4sKv0
sG3Ga+ypvhDkqclKCOxa2egyf0iG2FRQoeNbd5pG/Rr9jmf3wNGq/iTHU29HnTW/44WSvrbDbyeW
fT0grWJNxSDHLqFMZV6JJ6wBwesPmmNl/uENSmAv1T0knXcb8QsghhWHcSX7NK45+NEbqtu6G9vr
DYOD79p879s8b8+XlAS0vSeo6q6LxRXjrQ198fCJ8Y4IfY71ybj185C0Qzbnc4H8w5QKmEYz0Lxp
JEvLPU70qpEXm1htH40Dm9o+eJFT7wq2dOlKGCuUAVJvU9ZFNVmZbHMm7CzDPGTEFEjiq8uPsPv7
9BFMpP7u4tJxbdhx+uj+DMNnF+vffY/XQMYihFLeHah5PL855Uiy/2WC9rGHYBF8soFZIBX1JtMx
FbmAKj6FMbvBHZr/j7os5jB02Rn72muE/xwOsq3QGAMC+Mwp8wnXe+4vEhXIdnvEUgiddy2pp6Kn
lNuMMrPxMUzb2w1kLVglSHx0QN49hrxc4rpnXk+7HuZ+DLZ8xtoelmsTS3RrwOdfH4Ei/sCnFt88
Z+aGUEJUK+7foI9eH9hLd4T4aX4Jc8p6GqfXO5SGuTxo0hQG4Ty2nytPhFTmUZ4Vt0+EYsVQIIRk
B6BxysPHqko9XlWvS2ItLg3M+U+ljGjY/AiW8dDMijakQoGReHg5/71693r7qk+9lgRtlfL+mLBP
8A2xscrBzaKygqqr3nXxn/zhd94pjWSEZfHbyx/24FTkfMqLhZRx1xRJacrTUF/fFFeTo30OPob3
ymbgWz11BE5jjRMjxWLwQdt+Ruv3UHrrek5b9J5fvvIYrU49v2o2n8FSzLtcMqHAUICiApoiRscz
+e3aoCJhjFedY5v6a5m0xO7In1ts89mUoBHaINXwIZB85nhDLdho5+esr8zc7xu+wshuwbMypRMD
QAP55r8x4NHVXxvOtjzIxxlnbebgpoplrSxQ2zzeR1uKAN3q5vimo/XlsUkKBNHqv5UoxaucB3TO
8iGf52qbkygedqmTj+I3ddvf180OCE1yrRk3IvRoQ6usENVetP9W0hX1K1nclVG/Te9z6wd2EAyn
/bNzuCyWSNBAv5AGESyt+cXG6p4Yx7ewsB9dvRnZhGqkfkDDJuB4UbzvCzhGPeiDeo9pzGST5At4
5Akk887msKtCrZK8BjGyTBXcl1dmEJjgEGFPgdUa3k0skOLSdmxg/uzbG2Eagyxi/l5U81G6dyTm
VGN0ePho9GTDDIejTDXLwK2FjgS5z5MnsCpdxwTR9Oy6jyCfA67bPEZKS+2ugUoYf2A1/WLrcvne
PBaoKG4Xh32PlZYxsvE2N38ZGbysZzIy3ijnCRO/J9CZPKlvVOqYiD/3omFo6KmbHKxTsVqWXNEN
+m5PgpaprhGQw2Lpj2LzmsK/znmUOoY2gtmOF7Q0fXYq8cwtEY7hep/Z3woHVzkFgH8AkFE7Y9x3
uwMouxt67Ya65n1Ay+QkQbHS3yHtVNqE0edBonTiWA4hF4pbjV4TouLGd48PyDmZlvxKIeWnVhuT
fhZ/Kvk2DfLsq22/o3WZMy3X/9DvtOLAi0UgmN+/fdIRB+yI+zrdB31we4kRNZXL8EP9yuFdNxid
F0ZtafM+XoTDT1KcClDhbTQIgDHFCjfGJI0DHoXQgRs0DwJzA9NuoCKPL0Ya0oukb+h5pB7ZqRT1
sDN/eRVNC9J84iI2C54HU/z1S/uEg1lIzmZq9n2rA4GPrCjzLzbD1BVZq+kF5fypJYG7sXo832qr
dRf4r/4eefkyFqKNZA9oYlGdSZGqQYW0LyZJ5VAEdNweyt2NM0rm5BHeml9Flc4JZEHbPjmAhxeq
b+Oz8zTwscOizuL2qFxPzmplcpXKazu3f9uGE06rK0FYfCfMLYBTPpCmW989re7yJsvVB9mwZrk2
Mdj/XTuxCQmKU9v3VC+vN55cNCYL0FWK/aFWZ/wwnXstHYoGBoz7A20al+5PeLVryameKrjtQTCX
kukE6DiTw9DGbKgpLYW2GT1AbQHTa82gbkUfVbC19XzlrLL/doiii8DqilT7Ol7OLTUA248+BZxl
+oIpb1BZlwyUtL4HvEnahVKLUwEBPFOt7+WPikXoPTOnpNOT0rfajtF8tyvJSwiLiImOe97bGGyx
K+lHWKK1Wt616kvTXWyPwi02dcwZ6YHOIgCclRh64LYrF9YhI+J7g3IHpHWGpWmjUl/HcQYGUqWN
IazOf6PVLB1TvtXD6FbYVCZ3HE1m3v5tMOwa1reeybPpNZZ6G/SoJj0RCxLCJBXyEG7RzqrfvAqV
n2ugS1VogIDBFlZivPvXDwqFTGkndrm7lTQ3Y+pDT2tu5IY+jZQu9s47HqImU/gel9p/naRMiU6E
U5aoSM9Py8j2tKMc734MydIO4j7YHUAInaThwGpQh64c9huRoWU0tNwerYNlonjmP6ZBgCmvR4v5
MTsvoiKvXews8FctoZ8efRlpsTkSuy23QJxQRlNjRJKvkhCe02wpr5uLjpCsDKloy7Iq1URAEtAV
Rar0RIRohbnWtuW8+hVEDct4BT8st8me5eEhRkSiUgKh8AcO8fxPiOMB6b/ixZ/7NBta1w2xZunY
YN6o797ys7xPNNJ6iIWqIWvl5crYilSK/rcHcRinioFFTMvQ6IOl69oBtPcGsLW7v0AhC1JaMTn7
PWMAx9ak3rHzzLVXlI4Bh9Gc3oLk4xc7mt/T9/OFsLVUjefSfijvKN2iNc5LhNyE3oTVOgDLhxdf
SuA5O7AirJQmwvZdE/D1gQigK8xaPIZWvTbVydfMz7KdSArJh24cTCNI5GBAr55UGNhFQUpwIqNq
1TubAsz8mBxNOA81S22zr2lKtSWRoo9onswGXI9Yq/8wXKamZpdZqoAa/NZzZtRxYMK09cXZ6UFb
cvFKw4tlI7W8jMbmqJIH0Kpur0P2nYEQ6zKCrdGGirQz1JutqSn7dbZk63B+SY3LOsj4S+nlVYoZ
m4nqoEwNzmgyiyo2MpxFqzSxanQAMiDlF+308IpjB9M6lhiqpgXOkZLpAwRv6aqyOZU2Z2muOB2s
jYCGOoIVIQA0dpbZnal5CJhfEiCQ/MMhHG+/zoMoO8X9f8+R/pMjJIMzVe1RSrfMZwjzjjvgb6kt
e2+zrOVlD81TWOVpdlrqx1eUfYlA9y+XbVCB6DK4v1XhOgEM+A4vm055prTBrqMUr1OymqPE4TQz
2YlJTMaO7HC0AnsLvkVSgQdxbbf4Ll6oAavlPE2y3nLHdQQsVTb4NbICOKtGI5DLSCRmTgyUop1d
UHEEh9D+WzQ9GO/0hcB7u2SJZ1/glvYWd/YPbZ2yHg0PSAy+MWLMzLVJh73LQIPWMJ2P0vqSj3zS
2iAAnPQje2pjkx+OInQrr2447OapaY93sDFT2MmElgNPfBIwT2OmQccAL766B00NLGEgBUeRdZ1m
UL+6XOGzbX4YVAEVjaEbTQ1LkpMoLfPCu+7vwTPqT0NRnX/x1qP/gwQ6/Re58mciDd7o/nmTcnUT
1kdP7o9vorQ1WPgUdp8AqhwrE4EwTz0AZug5AC7wZmKnPizrA+jDWidfSoFSe7Wazzlb9X/SdhOv
xw/RxA27a45I1UJPVdxRR+kvLBz/y2LvQZjVE8WrFeeEIl+vSG2e2G84cdG+raQfh2ID6dWE9MI9
1ckwP4DKR8SjHlOJByweqWbqLkpiGxgQO84/cC9edqBsnybQf7g0KhZfCnS6/dmpUIppafEO+b5T
XiluVk2B3yaExw+2bgPhKKqShZVFj+E83XWFQlRj5jHDNiKKFhpuAnPSeh6tV8Lt5eQ5rimTvpOL
fbS1Kr4wR4dCtAfoPYG6Oubv7SZdQx6lLG6Vtk1A50Npqnmd9cF6I+j6AedTiQUBMAm3RI3lk537
Nz4IIdlVWi9wanNR3SqcGhnQLruEonf6xLqLW4oKYjl1woCVWWcVyhdE7dMTJM47SUGJwe0wImPo
hZuS90dlAjLbVaCwX5aRBXLHGmzoxJw/eCUYI5OSeX2HU24N0ymzusbWdf+kdivbZy+bDM/y1bIX
DOtlQK9jfwYALLQHOEaRAo3B/3M3qqIW2SJ9uVKDugHZm8gxYTwLjiGMGOEDJR1hlrXzrFvtwGvI
WCGwG57CqOFqLrLOIYIwSjrT4bz6lKU1xf4NJhy5zpE1L3XAPAaknet5trIdVw1TkryD8txQDyFk
tmfb1/y9QjvUTqmEEvjrb/GsX/qs9dfMFNYQzFX9UWSk/Gn/rbiBAMqacXsxyqj6irW1zKWF27nL
0zBhWB0ymAfFVBc1lBvmg6jiJsShMgTzoh/Slf9EDvm0QP6l2yDXVBTYjaNNjt4MeoVA7MLsqZI0
EYYjwFjjXgJVO6f04szNLvP2SkCI6nr6N5eBwve7n1SugR0/Hx5g6JDiQE/tNOmUbD3Aul2zrHtN
u2TDkozo0U/zeFW8qdg1rrVYEo5nT79xwkkdBXPY0Of2HVCUoVjFOVl7IdianHLR0umw0SYtdzZJ
QGIDrcl0nz5YH07un4NiFp/+bEG3JyqxeAtN7yCzchnkFjVDw3jXIPxDZ0TL8y30tCi4F3qFsx9K
nSuZDxd5otyO5tgafJuLVq+CBPbAgKrgZv+saIRP7woOxMixmgyAWSohAZGo1tZgvth5MT1UXFvW
gRThkC50JlaPjuU4a91k+Tlbw4lgfnx1f8eMgNvVYVWRodyqHcxN5aXRVjvIKW6P8r3l4V8BkvEN
3i6mF/ZJ7WmFI2fBO2qV5WF8pq1rRLo3KvpPNUhuyA6/GJZTEndSMakvlCpmdkZXTAkAGToVDeLO
3wtpThwfkIg8vLmMBPipXKCVUMcDX968jkWMJwMU+Bo195RmrloiOmBjsTq0SjrFyKGM3/AECzmg
xsYVUmKUwGpQMV8HoHssT+gYgL7zh6rVmD2X4IC1NVjWEEbzbPGcDJCOiOJ4AWp1TE7Nix9c93sA
4HUAFlX0kgP8+b1P3s7n2+mWeqtExCUlwGV5gSoYRjRyaIFznpeMRu5kHr5j9ygSky6UUCniQb+l
iovy0AxYELm6jCUGCwuyWKtwqqxDeU4wpu48huqwN2TVfjzHRrzTwUw7++YLHEBVKACNs13pUBHK
hzz+E6K7hkVs93AcE7kwqZ0L5KxOmz9dpEWvysK+X2rM21JigRy2Xo6GfSKU4DDZew2jyp7R0OA4
oZBYzXHWk2OHX/2J+GJWGm0AknVHZvSHXH3YGv2ly/cF9q1cUQGiqwnjDB5iQAmLslG8PzS7GfVf
/Tw8SX5bymqma2wyrCGCygU0Fc5DxGRk4dwJveZU3niRYGKfL8bT654ckIcyHZ4vjR8iZ0Jr3s9t
6OikpPMk0eGcH8/22ZAOmBvExAqeWbHDmfm5n7nppVEjsgvW5EXlbBd++ZOM1m6fDMGpb4nYkIwa
uJ54MvRkAincUW/rQPZ32JseT/kHdX5dIx07FYcon5fHcQ7VggeLMFSfxIuvqTMyBl7od85fCLiV
RgpVdIoJj969phX6lSzeMNqd9NO2yH62TXmSI19FMBsU1dGRxQqtkif/NBPLGTfxcXHtnDWgnrqb
uuSeqtwoj/NMASJdwQI3ItQslGc4hRyJ7EB0mx2u0ld5jtutawEwY8wrHFKkHtxqY8r1cJf+I3CC
JIyKX8sP/SFRaeLp/kSP3RJsYD2Ql8/+ENPP8ivSu77M0ccRz+ciqvh+ioiJ10Zs2ulvp1wADvhq
dudD73gh74Umv+TJKHSpznh4BjyqV5Y/UNBsaUC3n/t8012P1j9xDfAW6x0dr8W8wY20VuVXup8h
Bju5Rl741IoEntm7pGhXTuQxGlVeF4c11AYeDrz1OtpjZI4u3kuP8GB498AAVIoaxQi/Fg9u3jYf
G6pHeJgJxuVHW3MXRNF/1WV/NEDjgOmti0L/S6mUn3gCGEswN8joFnuvuIPFyjNydj04c6VequM2
EoKncWXAAc0edRqPOKVhvYh1yi7y75WOTGjEQhcHzREJfP2H7FITkytt8S/lO8jAVumlaaTuKBsw
3dt68IhaYd6lxPeTMTNEDPfNZVhAN/urfGlTZSWXHnAfmAvJG3NKBzeVvwgU2jL4pxgsPYATIEsV
tsaNWdLKV0GfCP6GuC0RP1ak3COU3uwLovoVs8O6UqpbDgAyd4b+KIsUqLTHfRGsvFh8rQ3KBNz5
8/wezIxSvIkvmMFWwMY+6jBfUPV+8A9Tm8gZe8OlmlyVmUBgF/izdhMgnwUjAA1H4KywVncmT/PY
o5K0Q0f33WCrDzBaPeI+sXfmAuXQgspvmCxOxZHT7tp82Qrg9uxH80hb0nGBQQco8kLws1c7Jaqi
cJradMP1DfiGtF8B7437eNCb2K7Rm7BfhvLQN2vaLl3gunBx6bkPo8oGzwfw3AZqWuQ64InIgQEa
t3qB7k4h5FTfhRWv4oFcym8XvEfrvmiZqdaplt4b/Vc5xYlkOBj240rahjsiIFj6oBqg+Nz07NMp
XV+M+uzaFsYkLxS16tV7HKhr8HyxmVuQ31rix/tZckkSeGrjbOy5dYvdF+E4sE5gF3ygLhqKbDdW
YOVCKXVFyi+c5EQDgv3NJ0tiX/YmwQAUP+KDFcFoQay8IiM4ar/wAfrVX/x7TKXsN/njQ8l8Y2rT
gBLNuQT6t25d20grrwN8ItdJnm3OMgYcxzutLd/nVMkviDqmHQOi7qcbco/ZOLOBFe5v/uRBbX9n
8cov92MWO17GpOvPTuxULU8it6GxTYfY2yEh9aYnJVg5tBLxzWd1apuF0T0TUpJaCMbOhxviGI6g
CzrgtpoVFCPWNdebNarzuBfj/0jpldNRi+zTp5Uj3mVFgBmizjWmf0beVBquN675ablC2r7ZHvr0
lYBIFx7OjWUgP5hD8UPYMfjlb1r7vUbdqJWhBhF8aAzbEYt6RBqcHswyxQZICEC/Yi+cYg5ACHAn
nuzKRbhWaHjus6ok633seRHaPfQQodBUOy3BGSlWFVNfpp/1c+kcknlcb38eBTFUwiYDipykrRlx
6Kn1NQg2FDe4bkMt9nzHvmj0fgeWUZDjiZt5XTaHy+3YUxfT+zcHDgOFVdlMDDv+NajMaVFd1uK5
B2sUeYLd2k/+xsRfMlUXK70ZtFZFhwHn9VaVK5As2x9tq5YuZD8rqyJ4blKv3Tk9RWpQJlgeyQoc
rIZZx/M0aEJ9Hx0Z4j483VoDNQkOQF8ZteWMLZC3Dxdut8y1E9yZlUgerupgUqewb7XgRrYMiuvZ
xbqsU+g0XhFkavTQH8RINoP4Wjp9K5RBCUKgFqPXPAO4J9JGXQ3h3Ava4POzJcJ1+iy1KFqsnoZr
8v3ypocOMtpJjN38nuX/NCwpUrhz4191RjjSWXDGZSM4jfvxWofPBWAkSROO8V9gomdwyVDyQy3g
QTVBJus9gqUQLbVZC3vQutohSo6Il0NBaeB1QgDAyAtgCdTmExgZRlyt++J1Q9oe/CPh77+OYf3h
eB7qc3LVHQwChLAjWtf9Iw9tWFBKxTrWcIB4tqiZifii1aMDQCf8OsdQOj34dgLNVtClUHdiakv8
f2HtvHYySZQrR5aHVmNIfcX7XBA0AvXQFhUBsU7IQkI8VALAHodBCrAAU0yVUixfO4s666jbDeTY
4qGg+2ByaqYboBbXYpMjmC81qe8KsZWQe5+5bNIgchhknly8gF4dMbxjXBROTwuY6bmmqWY/fQef
a9bgwcA/3S1UrKwOUI78Wpqk6lp3pWi7NCneMaorNkUwDweK6B7eNOlnIEWuwGdeY9IzQwky4bLY
NoDe4xa5XTbNd/hER3sF+l6RQ18pqEeb26f2RqOcpXAENe3PEYcD/K1mQbvGYOWKC77Y5hextwsQ
0ES1XypEuBNPcaTJ4Wzlw4byGBUi0yMHoN1AcknDCRePMZtIpWV+LbQAcp+C2XamKrh1qzM0xwp2
zKiFk3Cp22CfDza3KKQtAyrLSbLZmKKBtQaK2wQLAQoYem9yUoz1q5Bau/NBYKQ5+8hpYLDH3BFQ
HktVxYioQmqPMfgaJSkpf921yu+6mPwHOQ0Dmv2CQdAqvON1UYuCR1Okx/7yi6DD8qslfV4lHF05
YQoHTUk9BwLjy8GBYffJdOm/sTkCmEkMRRfkHMvKhXKs/QIO4IBruGp9vLSrvwreNv8AlqNcbz0s
cmS83xe9DDL1vL5DUoDqCO3bT7IjGRDZ1YiKVyFhB/W28mjQHssivol0xUyw/cUW7E2cNJ1K/8zT
5G4kHmYxYzMDjs22dkW/eggjR8429/OgUbhv3zb5D2RX1RM61h2HHiUtijm+y2c4DUjbiZkxatFq
pqp7HOnsn/HFcXrgMGp63Em1jE7HeBrGn3hxxCnCLeW7RYcJRfuhM6ynMI3dKWedH/g1sJqK6+ik
5DMUh13sj2agNgEXGpWvgrvwcMgdh4EIv079LjUUL8Gn4nOKfphFRRpxGkOJ9QfnLF95itbz3gMM
vZaNvaIb/3CgP/TdwInV9L9dVvRVo2/G9D9Yz5+PDuGrHCrSOEtedO47MbfP2br5I4/uA9vPwjpf
0hO34LIRQB+Np2W5wyKMxUQdP8HT2Lh1OanRxXHqdjL+zsbJ0OEHyhrwG7mrBPA3WB2+2QMDvtW4
P0eHYwlN7vvVPa123Z3BNn4wk+KNKm8fJwoKM3163VCd7I7m3z+fqXLbKSjl1dayp9M6n4dVkC+T
ETT8oRUfu7b/Z6kfJYBDGX+A/mrReLMf558oQEcjqQCikjJ2YGujYgl3v3qR3rqrWFns1vIgWYVI
UCQZlrbm8MpYOYXaU+pQCt2dVdKh7QQImuBrO6aSf3OBbWWV10ucbKW5oup3A8yE3k/xdKtKCYgh
xjSWmMau4qwFKDZciZjBA3UrxagA0s4SAOFFbpAp+RkCFbckVLBfN2GW9FSegF3hMLVC9lWYkgt5
drRLC/AeoHyyC8fRaxCQRG6kLvoj7khOgubePqsg2bJCOgu/WH18xWMNPauwHULCE52mOyzT/TDy
R27gogUDDqU4jv/liqpejnLpQz28El7CvHfUhMbbEsJDP/vGhccoiJUJLfKhXsg16PQeQZfF3CNf
pjI28DxxBDPCllCjsPIsjAapDe0WtjxKtDTQpr3Xj43FBabAHZYdkj7mRw9eCO8XQndH5PDlEeKf
Stzh3bWtTC3u9k7OV4HVU5wHt3nBmSJ/Hbdm8CD1CYheqvNoDTJDMDvmju/6RDusxfYqBSACsQsL
xoRyvkuFXbrQK6shWWvj8o5ktKDfEh9c/hRB6Hc0xC/k+ywWOduAtI3BlBb9WUqdPfAIUlUhLeIk
X1nHcgwlis2Ud2q0ESTuTWm4XyvXEcY8r/k7tyvlrzwYxxBpUfBfqS4aQyXQ/E98NIsHMiA8MBir
L1eu9BivDLSg9wmxyD6J9dw6lgD+C0MIyVXKYfZCyl665Kfp4VeIvGUz4o+zleR7NGRUd+PTL/Gr
bAqx/SJC93xNIBiwsms0mBcb5gbOgOfyotVNHFUuZ5cR0rGYobqPOqaFI53N5gWnm7+9SsRHNZqm
lTmvoRRviQiYTyrWhKBmlMlrRh1b0inoqm8w42cLdbch3+T6obuhf+5E50poQ7FNViAR+YfFxbQQ
Daz9goIoPqFknuqdA1yUd/C3og8Ego971IJLk++3zdVh7kVFDrEzx0ryNgwOZRXdAPQ5IoaLbyGm
+nvYoOa6UuckqQxyK4mKjGpVAzW7W3dHf2qJYni8RpYicq4YaN90l3AQ28xZSeY7tgEAbaMQ2xnr
BRyiyaPg/p8nojASs4qwvYdIBfRM4NVKo5g9Z6UoP/aScSPWsoW0Eu2RMUcBISTJVXaq40kr2WP0
hVbgh5mlJxbdVIpoztpxmzzKfZCKPwK2h98WmimpQ2wORS1WWLVvKl2I6cKYWMWPbopGnF4pZ+GR
mE8G6Wc5YzPXiZ5zMrdiB/67xHVlQaQPoRulxoRWapx+m9N0Jo6PJBxyKWAS+Pdm83jdX44TMFUP
irVadeICW842qhepV3i7qB+yv+SqxEHo1YdircyBRpIqE2wdbhPi/SpImIIcEugyCYZwmQ8iAu+P
cqDNuR/k20dYtj/uaoG5WUnV5X4wW1kvFocVyu30xqXnW/zjmppfU+ehQIz5CQnrmmpBDhl9H2b8
nuW4JeHysVXHXMeWJ1Sd2XC4Sr3yfutwxkdiyNCQ03zC4+rbPVphIqfx1RjFJZ5czKGLG8uDjp8F
/CsNSHETTyVAYxoTSsSGi1O2sqx6gcmtAYFb2iEL8lil5voWmcWHr+na+Av9hcdOhI9xEh1Kq+JT
obAA8ggA7hDeRClPAFkrT1nAb01xV/LPPDdaleOXzlwAmfgM3V6v6n93mQHatjK2K9eG8ZI9GOxD
ocsZvCAxneTqQAT4gL8pZ6HtW5wH6aX1MqwPzN36KC/gNVIL43IUFsRRjBfEwFdgYPVxsnxwXctK
jX4M57m2QiwQuAx5YrntK5mcNtNyeSCp7tZzJPIxOvqVQ4smxLWjH9yyN8WrO59MT689gqfFC1Gs
Ny8u2sL74GyBvWwTTtjkxSaxLQX+k5dASI8+Mp4z6JS2sIHtBzpIRxl9TWffgGj/4RdM99SDv0UR
ayRZexkikj0kgxknEe249avQEzBTJ9p3u7XjTuMN5ZG+jb+uJoK1dGNmMu1vsKgJZFduagu70qAu
o/rx7haxhlHgKKBu4KODAcczFmCfsRaxAtLbqcunrNpzAQU0QAdhYMKdYe9i/bm693tK943gw+h5
Sl43dq/AkJYRp3AXdtSFtybsX4sUtWSivvZKG7aKDi0oNo9PrhcSXJqIJ0m2WVD7ai2VYtYxb/GV
FTwQsfraTsU+x3uRLoN70e+zCKCrmtL0eXSm9OwXjUUQds4QKSs1/876oEQzaUNshNXf3k9ZuUQy
2K2Nug1+jztZWCVtDojFWNPaOHyNZA4F98CqjKOA4xLQUcrJe6rI/JsQTt/7jZjHtiovQxR91YDz
PHPuowcDIPzuo8AVU9g8oQBn+dhfvJ/L0QMzvU5TcaRl8r1mmp3SrafSOJK5wDaf51MZ8Qg7YtSh
y4/OiVLJqzLWQ/U7XFM5wXJ0uAv+IWut/S4hkIQiTbwnb2Df3aPCkdoIhbnDu8GHI2wkAkVISzOP
kShzmKV3Mb4xcAk2OV6ao2c0+qtfMMd3/1i26RrMDQNnhHethx1lIEJlwvNtQ0PRBXtYp026J9L4
Y+fQrZpyk4AI9WJbB3wZhh9R4YZgPShH8b6G7+Oyh7RaH0J4V5e5HshNXVR3ck6+KbsB9o/1Loke
2YjOto4LztND+7KTAjU7ZOqYB9nPeSt8fg6610u8j2g2cxlDCV/LWq+qbv8htqoLikHjkZ+eAlPh
umtQ5hG/zvtCGWSDbODVrSH4Tq1XVOxkOeA9LhUiVLjI6kWNqyzh7JlI+5K4dBm4s0j7SCL90J3J
SGwcTZPtTTmocvuEdi12/Y2XDrf1ATDNk3k8PUuWmoSXr7/f9rewoJ/znAuwoZls+RMVboAN+xnU
9t3eDmFVt1S2PTGF2qkuVaYK+b3GR7DBgqAfn5YGC3E+sL9Q9MA0Scls6JaKqGfQbrT1W39Okk5A
jXKJAEK48DbsZBDr2JeScvhgxef84dXfeQRd5n1fxNs0iJox0W9mymE8RprWIYn4NYuQVViKNyhR
K8avUIfLqELrqzqlqNVeAAEVNvqfyJbwne1K8xI6j1wZxfKCsKJObUkkF/UT6R/RiLzjr1+FO8XX
vy8FB8yAs02mr3eJqHC5kRiSmyQLqh+jqRHDv6FJeDTPQSXsaySkHVFcy43hessr7sF2MncAa37/
dsoaj1GMyKm7fF7IUSXL6j4AOXwdNRALlBvY3EX4U6O7Dkp/7+EHywDP1P95T5OCGscorze330aa
tppnt3LgZ0vCTuVeSGW5xWf8ntpuG/gjRXUMoh/cOA429z6eO5WnEyEtW2jQtvh61ANTetORrppE
4JCkeIhkcoMEvNT0CEmpS50Toi+mLg6JT/81xZlAmEVHW6RRBxG/6vaChACrXI7ed3nlmIcEdJ2b
KYjrUPgC7oQZ/9Aqkb8nY5oxR/FfJDChaWpJzfv0om1oNePEtXOO+/9xhqnM8e/tU1pxCnVvNvzc
2imZEleMIHWb8qkiXv5tn8P5zIv9bCrbXQSUKsj5HF1yhEA9KfWHthSzIrRkJV8wlx50w+60iY3E
0wIkXbki5DnbT+xXOKNMfHXqLLYYZ6hr4drfCQKudChGBF4Z8b9Ctqw25M5/AsUJ8nnbuNwzwzWq
fc7OzpAdpcFWFcs12e7jyt9S425BhgNQZBSQneTydGu2owSOma9ZZizisuLU4LrwIDPehsDpOpC/
8rSzz4z55UW0lH7NdShlxkfjL256WifIIJmO/CLxl/KeizsOOs5CkRUKR17XMEpo++zuoUAIFIFj
q2cveE51lgjuVLbcVYGUhCYZALXLcqFhOUMD0iJPQ/fOmKruWOjVSFxTgr+s2yfBHv8gOCR5WwPw
dlyUvKJjyI+7pjnaVa6RR1TtKcMPewjGGfKzsfGZartu+iLqleX0AzRZe6J7kZkEGDLPc6eip04B
lN/X+aXb0sUWtHiDkF/ZciXDBXLq+QnFxiYws2NoyW+3FTqzXThEcwV/2/4GrCdHiGQlIA9k5gHa
/mpYVn2w2fE7voHjbsmgZzqpl8EjjvbVy44BFkQGAokBRNR/xsW6zsgtqQw2HgikN7Hm2KQEsCDV
uqq4d/GDgvPi76Zs6eEWG6ozxFtJpzus41X2NYfxkoL/uDclABA8GaWCZZ0AWjRKhpVu4yZM9eXh
jSGGUJRt+H7pfTEx1VjzEF3mATPQcH5wNlU8hRBh2UyOtH8sk2ZW3WYgorpZd3hdbuY+jczJAccj
P+oGEgyY1zOKUfsh0n+vqhLoAD4iDq1dFoSGLhUtkq7o65Q6ax58g9JjYQNrZyUHvJ/Uq3Zu7/Lv
L25mcjPKkqQJNMycKKsVHJuFjJojYjnID656VAkiZ72fCKKvNEAXXay//nbKtAx8jbPgqjuvSjR6
p82/TCST3rrezChZgLJFmYuQz/rTzDjZMr/YCMmlQ7aMa/Emz7lGHeDpBGZO4CazEF5+wWXDGKyS
p0CGI952W7vxrmPnbsoubc0fG/JVDxBziFRhyvFaY3vB9C6TsZaiB2y7702xQ+30UzLj/TFghNMN
WszgxR15GuGwb4iI7+KM+AM9xPNVEM64EHpwijcbD1QF8Y/jXS6dthnryiGgD7W3ugjYx8j1f7L4
bFUclaXf73+YdTajhTXaa5kA5Ki6k2KFdnpSQ9EkRTZ/xi6KQTZRBvH0O3kfKRW3+QQwJR0ab4Cr
RbRoXoBavRedDvOK9MazR/A+CvJkmJcnnoJJRxCouDEetY1795oy2VTsNH2FqvMMZUtekmCtlIsB
Cp37LexfZJ4aRvPQGYkXDRlnxWn3ZrAWnMmlIpsoTFl9bIl0YqcyUGd0pCumeA7uChtC34hHJXh/
jZ/ZxTeOzfHfz7eKpovGYFJFBYY1BYHlEUQmSr4WcAga1xPmMSunqlas5/XRk2JSo1ZvMZxXwmpT
5tuMjDJeXxc2VF6SbYhccWLSbMgQcP+GWGJIVzqSsBfm8Mma8E8p+id0JKXQ3leG57ESzvJVs/un
ulcMZb1Bkpmiru9xo6EJdn5KoL+PL3rpGOLVsx5SztrYApqE3Hp3/j9brV9BUdaiDhvzEMk/cTEb
w5vs3OLkfnIUGaZBllsjI3dTXvNs5EZGNwIGoqt8eC+dd0vO2ByUpfuuoOC3IEHHPxt6T6PaDnQK
eOk7EX9UG6P6GVypGeHr6gNyEvYarrZovp2JxrqnfhreYsKbZcNl8OAmyNJxuxzmQy3HqyVx8441
ngdIIiHF7Uw0KFZgsDZ6k9VUa9TSthNku87Sl1ERm4cH5MX0y9dvm8FMcvAIdn/aI9AgsSIliBHj
GUfpbbCNruicTVIoaEb1+hhEqwhViXAnaVie654RNqaFN5eCS5VoCl9kJVhe0IdcbjE1QO0cU8nT
27QMO4IAB3PQXmZK8isOexyxbCluj2DFqpfGnMh9w2AHVX/Mkan9pX8nSmkCOpWTIC93EW+jxNZj
C50VS6i3xh6p3v09sUweEn+ro7DxxRRZDRM4OUVOu/m9U8gulLS8XCCxIRTL+IouwpKDTZ9cW8mm
KtjGSBTr0RdSWw7gEH6xVi63vJBHe43sxSPRxAAcx5io7xODcFhiiC59aL/z/G+p9nZ0N8/I/xZ4
8fl/Bg5ZZf0prEGj7lD1LROO2hh5WzdbQoH0B1emJU18HB1enW3pjV5xXDQwc+P9O61Jg7zIuq7H
SGk9at4s+wT40jxCclxMKymnEUhHu7OJ0evP8s8bqTjhJWkJeGZnSqXB9c4kr+Md1T81dMsBRrdY
oTNpQTTp5kpIAmanT8x/kmIqIuEAUrE/mMMOlmyAXsgJb882OZvFpwGWPNrFrqBLSq9s3Kpt3kPN
hBp1UhNrVtBCyqUO7r5adig2URZBgL8XrOYD9OrhKWrImo0C/IV3ksoJFSjqNrdiB7K6yVosBpn1
xxr39T0/vc5ZShHXlN/kgTroqYa56fZP40fZ2/sxyXJehlrJvu6pO1/sBo9n9/zYrvGOeMYNDgpo
5lpzwPcAup5UKu3B8YjGahTr4Eg3k3gmeh9AooBTKo7cljLN4XeYcf+ga4jmm2Bdo+aLZYkm8RtP
klGdQEvrkaRUNsUQKSdEMfS7+MV3mIoGk1vkTTtchwqIa3EpiINbZbY1r1jrc+NQ5+ZpZad6iseB
6feJV0BtOU2Bd0C92I7DNvjN5TKsQypVw3HDjTLpZfwm1EnvSNfenXLoj2MomKAqPv4lYSUG8ZX8
PnxT+027nxBQVpvtlXruhluOEskJSUffIG7HZbjaXAuOkuM8TvbeZWYpDNgbIgpkmazUqJuzma/5
PhRYxvuCi1/0UWD5Gk7NS+XlVnrwLeDjqGlQodxO9eRSVBXsAgrl7yk7bdoPKZyyXTQezx73vle8
FHx5GGLIssyY2xws8QXqf9tt/je3VyTwVD/ze1gFXQ54G5GSyw/sKEtNs+9zNgh8SU+q/1Ba2uG2
zTXIImndUoc+YxXkc9OZgAGI5yuRIKoR58HCwSK/lKJ1oN+PtoHJudXYvkv4aiZi9fLv8wKMQSqi
pQadtWY5A8BSRVB6IgO6NWhX1cP9VBYXLhImHq6QlcLvrXntqLc5m5MviUFu0BZTPoacegEZoq6e
kqFqB7bqs4wBrb9OvRnXoRp2YexnjE1aRM/DaJDAIBsSuQoDq2aO8q1jImMWozCyqeFe3g/baV1A
5kIhsCWdGqYvMz54Saa9BE6SkJCCtC4LpY80RCjFWNnEAJYMTLVaeHo3Zusl79s6W9PlO9na/33o
nfDQVlYOWSqwFEvjuaMCp/u4A2q0JOyTGjOHWKE98jzsitokPtyymn2nFQ9Ts6r/PgvV94Dolz3F
xPliMg8sgAeNiEFhyPC4Sg42315acgho0Hauxb063fUwtSDqyVS5oDn2U8TXluUNULoJs5XK7Wry
yoIE3AhmEkrBuPBlcBb47Nu0TfEuuYYXIZ58oKGZuVL7aNRYbZ3HVC4aAdbzMRdPDktJXbejJhz9
FgaBSs9QfGfys2/kv5cFhW0z7dp41bf4fsgM1rW4Ryct103CaNIZB/dQVVETFK9Mldz3qmNBLKaE
9hRpWs216utKVciRFxUoXS82ue+1mfQhwoUCA+Lppw255eQmJGPR2n1Z6LAwqVdpVTVEfJowtkCr
yU1i3ZoS3nm5Vglu9v1CZsCHkneOxogJYPyLXN8qQOunQMxhmew+KVPqaAoUXiXeBNEHQyOPDyXk
P4zH57mZCHSpVnLw985jBxvvBfd49HGH+dL7pa3jnZvTOEbydkTdtJ8jtN5vB/bA54LAU1Rh+bQi
8wIogGeNCHjT5OWXGRa6cqD1M/NvdoQKj/ug1zqGEWBDP4l1P2JBnyf/Plks99iOS9mVGfAAlyiE
vbJYAi/EQ22eULw3u9fYkRiysYjP7JB3n1WkqPUGHdr5S1m8+nSAl1YTMisUVz0vhUhwefMpz4QN
onGvYz2UaJU8lUEqjfFPv1q3FuU+aLyDOLh60ckKbxC8pvh31shh7STRl/7DhDayPwnrfxaQxjQ3
FVcS+vN3ODNqkD95yZqNp0KcnC1p0EkqVaniypE8avoS5jPDFnwxmZ0Qit1Png8lYtegi1tHwBg5
+x8+d2YizxbktTl06ECIio2m3VWoDdTYT/K6Kq8PrFwypOONIDWg6erIiXm9OtpR276cpHD3L/T5
dxJQfAUmr5JflqAPTzXiaTR7E6XSnU9cdO7kHptA+SYHJ3cWdKkecrBbpRWtXBf4wgHHb+U5Fybq
RsWMK/dF/TBCFpTe2NQCGcKRZGcrL4oOKmeP1B1YIhHkHTzWoI4Ns0lqf8CGEx7yB/ae6JZLvvKP
CRPAP48ez+aX0EbUKw7jXZ069XxB9UkAJHtkOdF98Bq5XuXYRCp5RwxkjD6c+TmIBIyEABKAPMgc
6xPhAInFR2RPSZ368ETE+nFWfOUu2Ycp8IOsYpPMSSl5nEjdRj7VOX0pwmUsWjBUvYw82vJwS0Il
28pJxEMIpH+uNOGPOsu2VdWXkAgzjsaXBrazzrsB00kQUf/LjiXmkJl8XWz8HCbwgPK+WpRfNe7m
JLmqUpwkwLAe9v3cv8iNZxYCv7jQPoAKXHQfPpJTNlfbG/QYVfpGpvt3muTDdUB3suK0ciQiXgfU
mZJycPfw1YmwTW/BhQh+n9gg7PYNyMrE3SxvQPClTJDQp0r2S858kcEBNTX4YB8/qBbW5QvNByrs
oMWFxve3cR7athmnXJZzJ9lyzple0+hAFwWTJ8c8vmmZDxYwu5qBn8EE9l77ves/7inoGDbzQq3H
WzSdMld2JHtUSsjFWtXiTNDcPYd//QHfS4pwg/vtR3Uknx7e4sB02PW/pkRD3dmANE3QMdDeCsCm
q32d50h0zS2YYt2RX0EtchlFhC8oezf2qnloh/U4QvK+JZ5PkoKxB0utWLDcZBb3HeYo1AlKpLQi
gXp8cH7GPVmWaC4JvwWxWx+BtF+jHV8J/KHu3U+gWTCJoe62pPhu2pCGbEouHmJdbhYulwVlSP9x
SJzRrLVDD+EcfJYFvvaoa47TpcHdwBFwGIpjnwOykuqkSNZII3Jj4shn7g1SLhgf5kM6NyQ2S6kb
ICWTpYXKqOgplNcT7ohd5Mvp+0iB+jJWud+sYtKPvjUECq8vwM+e9ppMES/hFmMOQzRg8hY0NGhl
+mBMmbG0kkp/oU1glzM0OiDecRT/5XrLnak14u22S6TdvAnRVYg0bmLOvkTQegXsNFZgH2Osiz1p
QvGOLquzO00mUNjdhhHd3PMBrDA0jdFae4UAdOFbfqMGDSwM/EiDlbn6n/HADahpSyxtl8mYxl8X
TBCAHHklBKJfIz8XLnjjn9Qd+tjPNhA/tYRJzhrjS6tdKiBk8rARjLqiarmX1MxnEdTKxWaPWQFH
loavBlVQkT6kNh0Tbtqn6mUmxFUqdhS+fPF/jvQJjAQ29CdRicSUsNvZdXCGfpvMQYTda04KY3fV
vk+K+vVeX9dFjg7gozcxBc7XtHP9Z36xImpG2AF1Lh0lNoyh8xUVIPtSzVZB5XLCzuA7XoNCD7gq
pPx8e9Uzg68tOI1bS4bwvh+6NV/hNlyBEnIu9eEzpCtbEWl82iCmqMQqUymEvS+zYfbRKfSiPPT6
yuUwHfzn6t7zvEy5muUlrtaAgtFOoHRdEJUJh7md9Y1ILpXoI3JI9nXYU6hnF4g6d0T+NsNCSAy8
5P4zXh+n5CtgyngTBrWLY1EiVFR0pmXsgRqwEdrOcsPY9L2MbS0wxoT48iqC7iu71K1sv+4DY61/
KJ9gL/ZOkEcQRldz0X2zlL5CxN3MhGzIaB9Ho44fw2vVysYi0wl+YvJzgHkbh3PX/GfgzAVJ9i3z
NQerdzDiOPQlwI56SjzyTBhPv+3eD4m8uIZqsN/oj0RlRwSDN1FvNB8WuZ3m8D6h0Vj5D3Mk78+6
yL+jTUUCYy0/lSzE28qK3yM+apgw3AWymR9AIARq/TZzWZ5JSCMC8MO9+XgnWpk10BCu1M7kAD2Z
nlkt9Ah0srWt5C/BbWQVfui2rCoG2lq8ylg8Rvdpg0MxfxWvh/aqjpx5Ts3ri5vbDcs/PlA2xRld
lZxxa4XNpOtIZJMWO88eo2Tgk6R3FDEZEGjla2+AO/FlrNorMbeMQzRpo9D4p+nLy2M1FtzuXu+7
BxleLbNGInXeZz1f8zPsvq/stNENiUwVuUa+TvsO9oWxm+x09xwt14pU8gswr3jiblIBqsdhiSZV
yU+F+dOtm5Hkum40sGrHtg8N9U13RIdM8uba9l/c3LW/xzI9AudIrmcp9Bw8xUc9tUFaeHPyNCPj
XE2xpxg8pkrWKRM1RCcJxPfMlecNFnaBsiWqDmgUcplpUGt5hfhV+908D+uN2wdphyVblphadHbr
L5cDw6lX6w/jTmc9QvMyHFAB7AEvA4iAzo6d8yD+3lAMRVsDA52j1VqyYjzQAWYsLDoyqF6qxzVo
csiFYizn1x6y+td4NcRlDcuQT3BH4JTT9p7zNw5RprtAtGdF+jw6kcBrFM8Q+mrmjl23hAL836+s
2WvI/f1XhyBoPjJmqnSVXDvx0O2/OKCBEja1U71v9Ex/UP7sJOLSKFqLvMRLDFsfP7KiTfE7A27s
GSe9VXEUwQ+L0kSAV+kxH58AVpfWrNyzdj3MvLey5cqHVnfPvFt1DH73UtqYhyE3MXs5T4C1DHkW
iCwDtDnEuwnDKaigvMlVVfII7hxE1i19NcPfLQ3jg5DG3waqlXXbIyIytEctiw0vbWy+VsP5e0cr
pSQVYxsUssA8Xzh6TcYoy3TzbCmUpnoResg7Ci7jG3KE2XbVZ3blYUeib1ZqTpPmwF4CU1jcVd1s
nY4xMNfqmBIHkOPCXTw8Q1Dturu7jNaDcQ5Ql+HaMNtR2KBAgHHhZAXQH6fkyxI1qjIy1O+C0mrz
8R6kq2BjyiJ8IWANrUaln3TP2SVqgoC0M8+oOOMAJzfHTj6B/9fbeDH5syfs5PQP97IjvB09TyDJ
KRJrCyP0OiWb6XQjpXJIhk3ptfHCytErm9Hb3i0medlsjhz8w0ZPDa/AN27cNb1oGPIOAUUIghLK
OyVIBRMr+MbhXVgAcTWpvcwUZls/wo12uAHT0hj3reoP6fGYifzzIQNOzdlutqi6pNBYB0biQ2vD
47atrOdDP+VGbVzkMQWeCne7VHgwfqCLQw5WouasDH3qKtaHQ9NJIG2RFJMOGB6ZY6LNlZA12z2X
q96vEO4Q/ptdAUIMpQHN67e1M2tUuqlcqLZeSaxjY2YDFXoggPHMZugwdXSsQpZbj+X4hdfx0ImW
xNk0sg9vThg5NwhaytMN3jxfAQ8Do5SFcROH+t5hKrCj6t1OisnGa1u0MvQoAkwbWbGDKpswwMRC
akEhEARDh1AwI8r5A55H9K0vByv2HdWZZaEBuJs8jXsKK/lhxtiLGeNLPERSwHX+VRZJDSPc4it1
XcmzzG78meJewablke2GnW0Ga3VJMVu8+St9B79ayIlhMK6krmKhcdT3ZwjFZGpwV113zBIib3Vj
4PLYngQcvOEheWnqrX4iKfO/lYSprU25MKJ4iK6DlEmBWmpjjyimbkdw0FSLNnMswYkWVAE36LAb
Y7MDt+2eR/dkUF3Gyq6atp9hf0laN7hcq6V2M0DfbPyEHSl649DZ7i9DH9Cy2ZnY8+tylszBxKYx
Oii8zOW9LyPWMknQolnh6nDsAZzgT4gSaQ3IlCotsXq8VDsiTa280ZR7rGTPwG+m+I7h771LDT//
TVnXdkVVTXM8//7RDewznvjr/6ONoDDnFO5n6FCi2WQTprTNUaKZqtJbTryyhg1y8kmwwh/nfZyF
QzzjI4Wut5uwsVUDkI0TCLe1gMoYEz1PuaRl4Jx0D8JoXQjE+UcP8dZ7dj4Dp6wbP5QuvqNtK2Fl
W7bHhRo2ZduVtoxE1vDHwCoaQ228eQOPoUH3ba1bZFKJ4Wsb4U2bIV2RmfNtTX2PeDblqKuIr9rr
UgKJiLpI58QNN1sk+sW8ZV2cLlMXHR3lhk9UvYHjM0tJH2N+Z1fW8WhDrEEILYMN4Mxz6UciWfku
xnt9fCdP0YYaBqeIY3e6/AWSvkRwlAC/+og48x748aD6/b5NFIRX9ZTS4TI/9APSUsH7nztUv8pW
YGUhhPHjSxWJ5ci+5i6foGT4JC4ykT7Ap5HqvTSXQz52q4k4BYERBe+btJg88Qbq4oAzKQ99/Bde
iXCXmE0+mJSOPS9pgZbwv7t8oEm2cwjDjuHotnOod8H8pxBSZzF4qCPDEKXP2LtxvewUi00QTe1/
RmLr//XuMII6G07+7zpxK44r1R4vwhDUDN5BApwpoWorlx4reKHIYKT8pCJpXU+whkn1fV4H6ohh
hRK5omI/nq1h2yQ71j1VH0n1jm8QVm8M4RX+Exzdy3FGuWa2fE/t9ZIlruc4l2yp1tpFrxC5BO2a
1WTeqiboo5WI0HrsPTpGB9i0XRYemOkq/JsXUEB1W8rLh5PUOOhLT7+DQI73XAXNszSAWXsE65Xc
RGXIXewW8dexSiIgHKI+C8ruXPtL1OWSYUz6AksROqPfQew4HpJphVWS838q1T4HCTZPtFZnQob1
yOmsDtloMsAhO8kn3kDPw4p/a/SlaT8gyPgrpUhHRpaBUQK78lRRyYYq1St3lgTxthtcTfhMdKZo
Z6tDZ9BCM8KWvm4rbFRslBGSb4kR0ZJmE0T3ei9N/NvZCqLpFLMVZSpTP3NU9jn3Ih/+9vABbBIu
mN/pTJ/8aPK2ii1jpKpUcdiklEK1hZE+f9fTsbYiT+KQghoZJ4u7tXw000eusyyVXD++EA8mwRY5
t+lzx15KTBOdsWi+zNzuoBBw5aVpSPK2EFyPvY5E4uEJyc7BLxsfkDGCB1icbfd+4ItyYXd2b6G/
omrldhTYTDp2Q8a+tHTmoMI5rpeal14h46eOtjsuF82LSYohq7uzcgYwCCfnIeEsxyTm3MiJd8tA
ig5NTgYQnXtRiDyjsp6Du6ctsev/gFCVHOf4Lh0XvdOTpvdns+rLFxVkdaYJ+sbNTarIFnlzWDOV
iwPzpNA6m5VMF/FTBEK93J5VFIiN/QX29YbqqYLT/RQy2esvWLqVW1EXfBhoWQ6iwqN+6GDAyPIO
OvVO5nV3e7ZrS8ni7uviUSOXcoM2Sbbnx4o4c6kdhufMxJXwuzbtQ4SaOCGM8Ad3d7ZtX4jTTkuV
8rSciSfUrGMDnSzc8ZD9+5NU58dkwTvgG+HQCLG21MPnaLkQ83balyw68jodfeTOxRoZXecMZ4/w
aox4chXU0SLLbhK0z24lX/Q+2PLlXwjgTL1fTOksDa6q2ITWNk1S0YsMBJmr0bzRrDYneVAs1my/
cFXYtALs5/fbnOpgPvhGsykxd6999yz+dfwDZ2IHvpsnghuSTgSh1lTeVVAomCgOGEq9jV+CkRor
X0EQxr2DP95ZPxryf9fQG+yIKKG1ptlXPZFuzh5R4mD+0acr+m7+v+jk5/y0G1KQj6pZVnHckcx9
6r7QJknLE7w/Aqd3z8737U5cpmg9xjDKhmm8tcvVUG0hCOaoAeG4deWRQXJ/g7IBNm8igrh3kYds
UCyW8etANuoRBL7X53P0Q2uS1GFqJsAEltikvj6K6KDMvvlYE23ZnORzxbj/LxLasTJDSRl3ds5X
cfyEpgecAQ8FNwBdRfLMGB7xgE8i5FcFNo4S18JIwd+wjtGAimuWdT4Yws4LwE7wU8p8AwGuqz98
0ZGiGlM6NGPio9goZnBRdzuV3vX97FidgOtCjjaIk5mOgxb/CRMxeVHzP9CaxAahk4SznspanIUf
W5NxNFz5rb6NqJe9HBH/hLGeHb3Y1jbSjgdJaKhjRb6zLIrq/EE2/TSZfLvGS4x9OS+ATZzjXaWg
ebifspp+lP36m163wmsNCAdUzsnh2BzjUYqW8Q383ZTUQ2edfzP8S41hCDg0Mp0kagFZ6FmUI+Lr
sSI2WukNig/IuNjP95YZXT3EeJ9VsBkrPXOq5dvdYUJUt+Y5jx7Hj3C/dfj6nZs1NhiYp/kzuh/S
RkNWfZSY506hzAiTjgzGIyLGct4gpBe9dDqPVOmiAxqtKNE54a9w4ICsSiQRkbo/C9QykqFfQHIv
Vk2GH4TMoBmEkw7Ygq1HU440fsePnHuXmD2bQwWNz3e2Atll+RLDr6lh7gzcHcgMjFVWqXrQ2tT8
0js9TMS+Hc1KUlcVPTkkOWfDQxO+P54oik1cLzFTOPXuHTbxdeZB9mHuj+xnG7Uu0n60qpJ6uT1W
k7WDkcN9+bkda5uki9FBMTiXk8WDzTu57/qCrUr3k292fHOpe6LvavUUWpNWy2nZvNU/Axm/CJxG
LXgtBegu3hcQsb2BEPA7V8Lhk4XzuOE3/PNUH121uxhGECOVf33vDWrkkE5DzS9KfXW4r5e0vXk4
tPeenBbNYZTgPaIbHg6kK7onSRSA1gYJjOqpd0uFlUUeGsxrX4IpWfjXb1F7HPA0LlLvW1ET/bKr
olzIjNIiwENjtUjiJkk6uMV3ApDXDzQ9UhOX1YUM8hN93F5Us5Vav9uqeyEV/TGiilOCEiGqolqB
3cDC+IT2QjXjSuIOCGu9xsrFIs93uxISykyq3mFfGIyWTxA1yGICfIGlHkFB4lmWKTmeCy2w3lPv
JqDi3WDITRsumUqCd5qNJLYO5B8Tx2SaT26fP5LWm1oajsteZ7K1/nxCRDIxOpNdJ3Z/Zdi34tFS
QxLwhGPAmcPDuOvT5569iIE0jcD91ufN9M9MH5JGvbOznm/VJ+4FSAsbzT9iqrAvq3a9OIh0jeKB
aGDnpOtuKx2Fq3MZTmO5LiyRjMJ5IN3Oi9FyJBBsaSNeyUr29h4I9jBSwcVuGlH9hNlgtzrZHg0J
MTXlaME0HAOG++LZNuwEh01P7K73FanumNWXIofeur5YD1JIBDYfSg6ZFQ14rVKUHf8h2vgmU7LC
BgIfZKagUoNWo7/VhWOdm6rRfZc4uRpbapACWpAvb1vzvx/gIxM91vsAAGhnWVaLEHPaup/8WbrC
7lhcUtSgMKKfPA5ScY1NpFwauC0z1GqjfE+bniujY0W0lifbwxLhssSBQikvoMrc0qV9Jc64Nmjw
xqN8P9Fcp6VvFPPfz0rtiEvEtqxGM3HlmzE+wtx5xlI2VJhmqvflbI50dUDvSiDO44G4CLLiSU3f
E2O5SE7PRXIvJlDeOUt7kw8IpLI/EmgdMLtrhoFdGa4h02I6Hn238wV4th7ecbT4oy9GlLE09KMF
TKrMm2k0kLoBmahWUPBec3v7sc060XBDI0r2rhOIcNw+IlRH3FR3+eff4SnW277qQkBob7ZQydCc
fh/ILX3PxifYDFVHm+IUdsiRw11BRtTDxfbEaapynI84eaH5Imp+OF/GGk1nbP5AXTTAS3SwOxTj
NVQJQYvDBpEMSgPdimNJXSVxK8TLzDFqUvP3yejF4gJEAp3JXpvFFGkMY8qKaH+LqNhWums2JjgW
QW8Bjxf1hakIwshVlaHvOeM2wAKB7S5eJaRd3ufac/6duonYAr72jcGcTgK4tk2of5lrl74HASvM
hnA1mEs2klhuBZjNrCfSDcQjnnL1ST1E9SdjlLIOjTtJNsAjApuutUSX7rG32hWFndGpZ5jAltuo
VGjudraRtmrATlmAlkj2KgAU0iAamva8qy5xZieDsX9oc2lAk8HyGlPIOvr326KPpuBbJRkToC7c
9vFSFoUyYj+FcpnSHHuyo1F7TaD3iaRZj+pCTSRYr4Rwf0f9QlVx27l+irWZdy1QXyYCMaqtot3R
gunmeIIBY3t6cGMtatnpQu+LycuQwVRY5UKVbr+7eNsfSzKS2/T//qwK3GtCVrXjWoxVoWhkkxvh
/y12rLMBfQ94J/6Q+MtrYFTRrfQIx7Q3p8M+XDHoRadzvyqeeFsLCl8qhDCLVAZglwO68WUKUM8j
FgxBRC9pjB+Qgat+7r/tUCkq854dqd8wsHi6RFvI1N/vD1bzMCQxAeaaM99Ox48unALLRiVgpYJ9
BXUkgyfN3jdk0QZtOVGEusMjXUW6oexJOnXbRBFithw8d+YylZYEGBtBgQR6z7r5r7VMOi89Pa3D
f/N/jcntiAkX4F+Ph8XUtVEXVNgs3BLc2v3hb6tAE4yyVe1P+kxuQYFf/o+r4RaWzLyF58DpSgR0
a+2o6k7CbE0zOx4pP8asLe5WD565ptPNzLgJ/Q9qWZBBLfz7T3EUI6CXMVTZvuLSIEgpjtWWc6Xa
Icyw8MYYrV4aoAIJx9RnguT1waPonN/Vqe478FOBLCOUusd897p1iJ26Z9/3G8Yxe7p3z6i/FHip
ciXN/xh7QuExwGuuppCBAjtii5mRkele2eOGKbwJXt5H6XzXz4dvcjRh2VzEf9Twu8pxDt/ftPBg
6FR2BbD16RKc441CYPjbIkHsJtv5p2ukhYX9+Vya/LcugiPdFnqvYPdadr0zkRuiRJ4H73ct1CWH
umjP6TVi73aRG7LAQ2jHmzRmmGb2Zh+oBlmBwczyXU3BQ0qd++NRn/zozQGoRE0h2DhUatAkk56o
X9OWQ0AG/0nWYSw/8Hdh/g+r9vsP9Q60xb99+C0IN2Tc5fceI0+on4GWZr3Of1dJi8itgErMW4/H
AcyyPefgx1Rr+bo4a3mteOBFwyN9vUKod7n+KBa177QTvjO7mOs43SccQz+nZArWxVyIu8LoR9zs
WyDOJ/vkZ6Txl2c+UsJuwdkyxK4pbqhC+AG38H1sjGhDghk2mZ0ST3Mn4K1Z/gm9Rx0llLD3xiwt
i9Q2vCqdmVmDHWpWr0ufwI7zOhL4vuzbbYVwpP2foBc5FTLkMEa7pAo+qQnLw7u07xRjGqf3B4JG
pRKBrP9IHl4oOdFbRlrxAbnworu7aHlPOEmiL2VLCmUPd5SW0P/cUn2Rl0+kiO5koVp0hLSKf+H8
336Y6YaQzJIGYz8FCCTRM3yhpBlM54sFNQEpdQcCOUX8Jf2YM2pgig0yeI6AaxxRHqyDp7pX+rnQ
k8qk7F/jyRXhdXzFOs4TmGf/P1nmSw5FycJdGuuVyeXsZ1F5zMTqw4Or1UGXmb/U+wvsWTbN+/yt
eSGaQm0N8hB2MZs1rB0QvRCdalQFBYIk64XPPUr8TxpKUQztIFFLCa1kstdTj+dkK9KHbnXA0ngG
O26jen31AfuOuSyg5ZEm30T/hjAwDdtedwBqzlzyQjTpDgQ6VQ+izo1oKAmVH1I8g+0Oa5jfrqhs
ANeuKDBHfWbDY17bKhXgvYLZnXsQVwdruj3J8uSIFUcM92CXb8AiVOCL+3zMH7v1PPvU8j9rMnfU
TDME4T+bmYJqdRpS1qIWQRLsf5jiFMbLy15iD0IjWm1nffo/7cgouMbR8V95+yiuYF3iC6tbG3en
xS4lyujZ/IL07bOqKfL0IefkvwWBlVmzQ0IDffn3iLemGH6wMTI8HCD5X3iqBgwWjG12HizYSYuu
0BgJfKE1GTt8W+MXNLjGt+D8qFfLyaOwjJivsMzDjAt60oZ00k/EpgcdW/b11cDGMcK1/IKy3dM9
UgNebdjfSm52EEiQ9ErWdZZGFusS5BYEYMdXRdwykh5eoGloTaGy5aJvkFN+5eJZl03Mt6nhmaH4
rz7eSZt6op4+CsYGGnkBI474XhwsYxiCk8CYIWG425bXSdLmq7XgBa6aMK7k9JpQ30gIYF/JBBtV
vq7Z80UuZ5tpqCRkk+VsWtQ3a31nTpJRhDzU5LRzoqy8KsB9ppjyCXnWpFSpe0OP1yWzZVsv0WSy
XjdSa5M9tapIDWfF/EAC35TBImEzDK/itRgbltb3SQcFfB03sAuOpWebfZ9Z/b1yCOm3duQdiOV2
6zp6yCGZJchUdVmS57YD3wc9PFTafY0z0A7HtS9vgrXkviTegYy7tj2Vju5YITV/P9sRFu5EJV9H
zOMCLxEiIQBbp6eroqkqdPO5S2iEHNQ/Fb6qxNeaznc/9fLcSY4e4bqKtLeIkMUrt3i+gf1TaVgD
gieqQN7+sDRHr58gz3osNxviX2o65ZIfagaRQiF/g29jz6474uFBrlpjIsP30tCfzqBUOFnKfOr1
J7E5P1tgOZ7t7CPbCjVcRQBmmCyD2h7xbhsDJhy91cCrneF3D66+ki7w3ri2zkOXCzsZrE434jiL
9aW18CdZ5RiYpx1e//lBtccNRPShg+BEBFA6R5BqYmaK+6hlzurWOT0O+GNbr8dS9RYjzgV8fOvx
cS1zWgR7d0NfmBVE6+KKU/ulXbZ/r7ZOjVpQwWZFw9a8TxzgldKRad8Fso6i+WMDdyTGuLeqE8CX
NjwohxgoRO0h2zRXI0eK3zK2dHCFRforoemBQnLeg+dqYWi5XcXEr9daImQpFmXQWMaGUHzW1Ms6
ssmoJj5lUFwZ/m0Qu3niTOOdQwREtuj2oEyB2u5yTSNEGJ3I4Pd46m3JufCztB3rwxXf3AII5hda
yvkVXyf0dgib5EcwPDW/l1DoAfEQvpVZr0pb4sB4ItwhOkfqWd+c24l4ZHvLsd6+MqPuktn+YTci
VCj6n47rvvbfFDfM4o35NfXSsotay3tRTfrAU4QO7D/OmgCIdDlD0tCwQEeqRqSLjOOEU0vUQ8iR
ydWhPIAzsXc7/TuXcr5GVhXOCrLu3S0X+IU+fLBR1VQGTBzc/q4PEgR7iojws/PzCLO1pneKUhi3
SEn8jbiqmBWjVgZ2nAZUYHa6uVssCGvf2sSSVm5AVUUkcZ27Vl+r0sCTNuqs4Ijrltlvyb90kOJx
8/Jk86uWpN7XZnH08+cpvgSpN+ETcayfaYujfeu2NOyPwiyZBIZ2OozkeJ6OPSpdzXcsijN3aV3o
bA2Avm9CUNGlhr1DdA9wCM5OdYm5Eta7LT7uqA25k/in5jmmudJVwQzKC2Sd+bhihGZNb4qRyAru
Ywu8hXBV1oBGOFEj5vbhwv6g9btL8K/TviZEZH7TkprIjeYRKdy++6XQkrnF/EMbZ/Z4pd07KJRO
1d4gsU+lN3lemP/znZKYc5dPiFDhk9aIKgEMFgBcwnefpM3aG4E7MzIDUtmyBHBZhUkCkjzwCH3h
jJEXM08Ir8l8jdF3TgT+GMUNp1VgVbfYhsS64k3Nu/wgegikASgYiC8iS1u2lRUHt5520uFfSPUy
W2myLNM+d9xr/yn9fOmU0FZe4JZnnQdxwiTP3J30HMXMxm4OA5NjvojusC8NjV0sHgmVzrBy7Qnk
gQxXGdq7Aul03S9cSAdsWYJMgf2Uucxwxvoy59+Jx72rhU5vWBKDpuazqktmDYsm/Y8L8hBLIWWY
uec373hyidhs21+5LyelVqIrGETTGbUkTiYmWYZ1ZL5B4Zs5TOHhr7PRfsJBPC7JrLywb1KPWQ02
tUK4gBK/fpL1vrQYKNOVqsBsQyRGDcKJ+h1++ZBVORsRFlkES3xlNPYOEH8VJwEjI1tCDNNnv8b+
zdU3pcD8+Kw3alFToo3FgRNwVSpSdxZrnXXU5ahUSBoQtqM093oiKgQDF6O37z9v5PxdgN3jBF/h
2A28Mxy42pzQ4bshkM1ZtQcM7snF4KZP1de+AVkll14/T7a0wBijMysXe6Avg3jvWbnadOhRXh38
7NtGo2BwRfadUcSRhlCrR6g66eg+7Hf0RsmFaf3p3TT/NTtMvMrNrnyNK1QYRokldufv2FfnLrqw
R21kP+KGL2hYGPcvAQErsozn8q3T3ErppJskO5iaVTBtIvw+tY/Ag3fEDgksXDWRyu1T8kRQcRYd
nX54FZXOJxnqiMBuQTjn4CzMxzR+1bzbRK3oLSDRDMO4tKXJj7lFEjm7gFpDjiggGmciAmKOMl1Q
DHPP/NzLel2hkOO/g2iSjNRtO0uOH+nn0ZfJiDP05MpGxLja4KSx740Cucv6EyZl57zplVZRMkrc
0rpEiTfoSKDE3rISDq6LBDKjb4xrRLkVpJwIUMS83RmHWNaF8avwPFQpY4DnmKfmi32NYQ+g/Dkd
JaFGq759nquldObCKK0s++rzkG0pj9hydf8UKZkY0mKs1u9LPgkBgMzsLBBZHf49iHX61CqTkJUG
9Vd7XxEkA0BLKVs22Q3yS5ZMvmvhJ2bOKZdHLggONsE44JMeXicDgKRdLUABdq+7sohkC+/rLZJK
9OXJGEf1tSkThrsQYRbf9yyXJXXFn+RgKuvpwnxzdvG5plfsZvtNaQG9GUWfJ3XvozOo7Gy337cx
vY1V0bbBbt+GW87RiWa7ESkr7FiPnQgCdw054IBlE0Hhfir/+MyHHkj/W3/PKhmZYL4YTPvP/uLX
/CiY1HlleHg7ehR5DtE00eQPa2uwZLj2cEPpW0Ke/cFBeqz9gDEq7h3YpBXbLViKSacm+1Yh3qX2
MRHcv/KUCadDksMEwSs5dMEFQHKo6E0Pu30eo7Erm9Sw4JBFFRnT1yeDY3KHv2dsVIOMuoRVTwed
EIM2+0C/sa3ZqwMWtAGoP4wfiHXe7zQCN6Qkn2j36/6Ie+Mj/qbAGBOWYXtI5ZXINNcnLdbVklIT
4OdMgEbfejA+3Vw94Yx5GtQKl++uJgV1+oHvxBJqhx8XaoZrmohuF+y8sH3ThNxyM4oTrMhpXQr3
SpONlVG6UDobaCZamovStLLVBJd77izq8R+VIyN5N7YG/J9laF76L+Jxgvp4ijJqdBSOG74JazRf
9OFcfszPsmhLl6nF1H0dsD6EhA8SI9E7EvNvn4msBFuaeHB5uaqiOZ8xejSp0VhOMRgGPkGspXC7
DaAWd5njBVpcsVBjK8GIT5WHOFpUVaicz1ii/SgZAeYnyCNpbhXW358ODMZ7pb2BZrb2jR0b0Jl0
bUmGCNwPCBYb9xyihdRxR+vGRYCGQqmoUlzJ7SqhdY2Io1HuNMqu9AEa6hXh2/4X0BoWzKJwBF63
IGI5y2akKsh2/vn9caqYhv3LyBEDAXk8YTlCHVEFX9jUt2NR2gYkO8ba9wcg5ejtE3t4lgUOA6RC
l6MhKmzvS4IoKZQ8LSdBrsLrxPOKwbORShATrhEdjvCuG2uUwQCsQMj3NDUtQ0Ht9fDO8HiVyQYB
j6DVdvTuOH+NzbXXrmkJOSB8HEF/EVlSAREnwdYsq9tTO2Cob/XPpl/3INdogmluriZmOV9/ia0O
25YanabORqM+zTCKkfr3/kdF9nC5GYVYOS69PR90iVrHuNUbMM7vbIV2rNuLjLk4GDEHeIR6ZAx5
k7Y4OBGstUNz+4Mj6BfRizHl6poTJfjVOcXzQtNRHvfNe8TivpuPW9Wwdd9ntLlvZnlTTsfF+EVg
+gArkcQDoRVv570cyWJvhU1ySxNXeFKDZtKnmE1fnsAUthbTdNeWm3ncKe0JLRcZIEqR/cEwAHzM
2Qcpy14cww6iSok+3Iox1h3aokH3Krv8ZXgTU9YiSy7XJeTDJGsiOkdrc744MnSfmr46wW+lsyEO
DqHL8E/oDBZZMP3P6cIrdZ5UamhI7v8Hhu2YYBcMB/j93zYcmdYr+hxuQ3UsnFKJKqxnIzwNMIpP
ZEg9nl84WuAoTwme40G3K7TJgHNvXp97UfWY+0Pd+PuSAkxeadgyoiwTa8KiFzgAHC5gSYe0A6LD
XsE8mTc8073GCxTZPgofheKw6OPby0RMyCw9G01l00LPVqZQzrtvwgvMQ+vQi9XdqjstAloyckzL
FgUdGBWOm/5U/Wb9bvMaDruV3qcRCR0JAfUWZF1hGv1JUrrTxzPT+FgNMf571vsbxZqbvQB9PEK8
itvQzn4OIoeWbGoTXU2ov2T7gVpXsNbPGk31c4imYGUCFeEbd0cFmW0ajwDXBom0y1/IGbeZJP2g
yWuPN/gmc1lHk/PvnAeTjiD7jLLI56rHVDRMQ5jYtZDi2yk891phl+XWtLV5cy2ZrhMgbNQuvtHX
qKZhaIvBDIqNkcLLG2s+A9g1Y72nUEqInusxhnCM/YQGdmOD+VSq2jEZ2m/FT5Y/ntMm+YQZxnMg
jGL4+8JuyjoOZplnF0tE2KmVcWPHlY0j2DTaNVTKTO6NFiqsmRcyCK//EjUsxWiP9ZLTlTbXsotg
y/IntRxKM0Mbp9DQ0e/lxxA0Li8RgIIoCj01HtgbmRmavPm5FE8wLv2ZrgLbhyjvI2dAuwF7cUKP
H4Q+NrjZwlkfmof6XeL9igpIAynZQpCZjRupCtBW4qBP7t/3sglqJKXv+ulEwk9cwk9v6CG7pWBn
/9BaiN7nOZjWxUUBfFnwAUIjGFjgiLUa988M0m8ACaCXfshy0vbwfA0ZaH4GDXAjwuAurZ6cC3qq
Hua9aLjxHDDbLwhfxXL/m7Nm4OSFXYWgMiAH4w+B1+qy4u7EqHPR336MSKXlezukY+ukODZgyMX9
AMKaRyd6RuDKeipyYDEep08SlOF2l4i0OQKec7A3Qxy16wR6Xf5AuP22HVPOOBBsF5U0x0eSrvWN
eNPKFzpwBAIo2RNbJE8LsL1ZzNjjB3p5vVOe4KQSvEbApT24hCyfA3PmTQToF8zgszP3tmbLAUJV
fUfU5gijhO0kGAHCctkIX9DFpZFbrM7fRxlpY88+UXGmqb6UrbVtWvbs2ES5csR9EA3vR5ioL7cD
yRWmgHPsuzCN2wFN/Pbryhku+sxE0oMmshTyk6Oa2AAxPqHeaLQH6lWP8yoBWpmnBUZPYUVT75mr
Uye871B1bYu0CkglD0HX9CQYJTrnDM7nATJSQDs4855iBC6myVeJVvgbZ1JKYXopSwXXt5nsuzkx
HAStk9SNTJeJ1akRFwAP5lx7l3hGXm0gHf+/UlpbOGCa+OL/cARPdI5VbzrPeHJqtsYPbLZBbrKD
43p2YEcjVF+E23gaOjuwe3RSfwrRM+buHW8288RwGmrsSVp/A8sZYKiXvHmGq+0MTcPTz73wMM0W
rYiB131IgfXkNvx1at54Jp42vUEeutYTk4u6PvbJGVojuA2JmwesKsV5e0OBESRqYlpFeE8UL+qN
3GETFRpjWCK6J+v57af3cptzx8FjdI7pbTKfnWsGTlQ3mPIma0CCLT0Oj+k6g/tCi6+PRI+wsUJq
F4ApO59uGElBYZFIBaT7Yponz59tinn/KlXBllLFm7mS0qY/P9SDIDgfi2lAU8wP/45bja/GF2fX
2/7hQydIr3zbrSvag0jyRSKKR5NWsl5eoF0kUq8ltCnXR5FGB9xqDluRKYB6cSH/y0Lpgil82kyX
3zQ7ftbVg4vLhgPQq8B9fbYSpQRee189qXO3++IiQ68Um7kGqFdhf2pmm7gN01B6rGyzSLyBANTm
+dTpgPcHJUdtwN7RV2Vv1T4dwNZDwZaBASzPgTdG7QtOoAHFM/gn4C7jW97AIIkDUVcLJYz03XJL
veJ4Mypu4mq4qvo7iTaJxlXK7lgYXm19tYZM6ly1KcYLUKzMsru1kf4RATnBdkMLIaC1UnxihI49
NmPvkSfVytnDQA8I34d5hD42bPi5TfAsIanO0H7q/a6NksTnbG2CHEIhXNydm9XkkYmspnuCIJa3
9zz8m802B14tZo2q9SSNn21QcqMaheOgAMlZWGszIW8K0SGYW0znrxxXf2nqJd7E/IR/kBZ9auV5
wu9xtVlY51H1IR7NzykLccQS5k1aJIFZL74+CiG/uv6LL4J5+GA5+QEPHTzquu+WCGGfMntwKMLL
qc/huW8X21ZgGOB0iIuG0GTxrGvTwqMAdg7cNNPKTlVjwvfShnP0LNxJPTSlzNahiY2yObNKkApE
eSA3jHYLB98fzidPqPiIRfdAfs0z/0VaX5U2eiIHQZXDvCDHcw8Th6QcvMdY+0qqGhxQhwwzYp8B
npvQh/jUq9PAYzp0GDd1JZmumbIDQNQIBsDBe8W6T/w16He6+2lZI1Q4kUwYseTZhtMLDI76tzlp
DGKM9tEUC4Br2RMMVysaUkWWPz8H2yGWV/011LQuaIGC2rOU4/1sHpXxfhG5klI+np1Sqd0Xydgs
Qwwi2YrDL+sIf5tZlwLZP326UjOvreAhCiRgSuKn/908nbEF+GHTAt866nLD2j6AXBEVJ3YcxBbj
TXd3rTc4Ea+uqTku+1gVDWyyKfbFR7GFewbXe3jMFRipeh6Ti6CRBMx2ZRaBs/xnVrrVm0DAk/g9
mjC4lqEFNUHDEG7zvLRNA4fMMEyiIFPOF5NZMzkFjkU59Po/Bt1M/fSQFRzPLh0aw4rPc7XC/pxK
XxP27kgWgTCbZfF15H+UuJEss+ygRE9nMuZ3y8f9i+yvHJInFmjmpfbywX42S/mmajw1SPwb7e+6
JL97sBwsXquzrkRbPbGHIwk74bawdC5ORFDyqJEBU1T69oQgrX0SlZBZYcSHWq+plIav2tWv7dHs
W97xl/gzX753Fliq7OBhNScRoRV6CdrwCn012ughbXknO1XHEcnKeupruqB1lRhO/YehtaKKw2ju
cFEfealDHKlhIJlMKqTRdNNmcXM1HcpXoYctlUTwBvq7kPGDbVe4qsUYKiCf2t6uiygDv+Q3FCiZ
eZdJYUusx7ukDVnXl5gslJDWJp/E3TP2a4BjjdlJwFU5av29l4ymfL73iem3203m/6WTdNnlEN9n
hXjpsCS9KYvzEkSYODClCQ6nRuqHA1xXS2OWuhnQjYCPVDcNbe7h2kssvoYkF1e2Xxr1v0zMHWxV
8JqBHEdaAQ3XRW9iC3OsODeprTH2PYFXK+e7DFg3f5EvYLbtP6xUTJprF8Wb+bS4lMrSX0UWf6a/
vh/nO5yPUY3cmo5+3HXXTUyPYLenNoewQPlXaM4Cre+0ep+KMUkbgT81nUlazpjYYkhR+dqrsPeC
gdSXeqxed8/JdAgaA8HIDOpmtLJf6pZKTiFpeiLdSJ6E+OkfQDNAR0+9AdKcGEqJd8Ii6IBIow6y
2Cfl6LG+hZbkCXkUdND8bbpK4tsFzggPzUVVaROMNU/H7TB8BuiKldAZTrspuimcJ1b+qsfCuc7w
kq7jsMS0hHgeCmYwmhmh7sUKusD/gz0iSR13jVAqiG/1utL0Bqxu386q6pyiG34VvnDN6RYxlMXp
0iZtl7hXOAtU0lK1FF3zkdZ28C4zrEzYgN5c2cmqlqfNT5f7q0F6u1wsjMrCW+hTqrCsqlqd/dj0
Ad1LfvL6hIERT7eIjG+mTVv0iTKG2wndAHUkg67OMsN6rdDQJQVTvhw8VewQYMnbBfNVUNF/5WOJ
ptPb0HunbCs3xyGMya7/bZpXkhl9dKJJJvdTmhC7jOd0I+iTDHJOuje1G9b7MVHKq6caaWOTjxQO
4kwfyUdGTUMfBGS0i3DOvwfBkx+58EJgoistcOkZcUF/KfQw7kpzb2H/aPYtdp9GyK83qhrc5Spl
1Wo1uDZYdlMkKHHUb2W1s3sksmrCXa/aOzDM+FCRNsy6BqcFU/nb4hOvyewFHKuRq2gBEjqVVyXo
kbHNVahq1VlfkAAhgGJIveQLuqwM/PYWiracFneOgsGsyOFFrKLXK06DRsVUrjIguQej7ZHb+om9
++ojKy2w490sgFEkckB/NasD/U8rSKZUNeP11E906EuPYWXgLYCh8BE9jNkFGpY8qgXATfkNz3Uu
pXWn9CoJ9fvpuAs5nNLuJXFpk4KcJ/8lWg/VzpzGnVQYdestE9EoEyRlQnDZeJCBo6xOFowNQbZz
5v0Afur2ZNjky/EYYC3EPKwiYdqYk2PDyDLW8gK4GbTCqBerXCrBJ+EBlIlEkl5NdNbaUb5Y49LI
hegqgutCgMXyF97mtV/YF1WT/hvvi/Zmb8z04ydNGApabSZdS2rLJ8QRr01dZDgXTpVg2j5NQEN2
wUTlDVNcjoU4FPJb30oI33+YGvDOG+7x9fwDCPSrvto4cx1rEsAQM4e1uiVDqFqk+5Ts3oppUKAf
cdmwnGkVz9pWKB8+HtMADfYU8PqRzZtAejUMJOwXd+r07UE4vnAj2Exc3dALFw6oLuuWPhc0O+FB
6VPSuhhBFjHnEBWIUFi7mq4NNq2knPhHq6L2mRm622Mzfq0AbVb61rvcbkAEwnRq4hIpIX9mADvJ
6F6vbF/p8x3yFP73c32OZYJ3nvoy4gf16PPHWwu+umEV2bbZHI7GPtTc54xGLTvG4DnRwfqRg83l
xxv4aijHIYRfG77Gza0UykUY7zBr8e37F5ChNrd8WBR/XV1pDs8m7mIgeZIZfYF9sfWNpCdTVmir
i5zE72igy3n10dQ3sGxcZtl3GTurdGW9bD5flmB5Z4p7jPh2+DYbF/SSYwdVlbBwewBO7Qc1T3+m
398dfFvWyyc/TM7l22g7hBVdBGXbmDdsUI6jiDDi4nCmB1sPTKZbt6K3YzL1bb76mKXZVfG9K6rC
lkbots9b0VHkBu7iMzX9f4Ux2DK5rh9CzsJIpbwJf2jqJYK6qM5WaA1TJ9sWnpO8A6hhGV4Lgq7V
6lzDCpiDudVSJYXfiaOLJlPUgYvIgCHh5Ac4WVmnu41ecAivk4r9nU6NYG+pnXl0hiJvLtuBA7pT
MG31L1tg4+2UvdBWc+GrYtOc7Kr4Cpgzc1VhgNNhiyyFhB7ofaYI9DCmOlD5p6u6POL2wxgUqNaI
+HkGP2mPvz5aN0HELUVRoD9DUw8rRPLxNpan8JJe/SBxavxAL37ciJUiFLsmZW/ymJIy9Pu2nSw2
RCeKIkFhZ2T7dmxZ+TwDj8LugIYr/jB4fz6U3B9ZrM40Ebg+PigNVx3Fyvp/h4mIu6oJ9XMEX/yG
/GCuDPf/KrUZddypj3G3ywC6NAIGaLWLhigwYFVEtnI9yxxPeBXOTKmKdoN4M+GRAxJICy2vpISw
0w7X3vbTJDtjYaz7bDgwn5hrR7iNHyAiaKAGsgK9Tq66wYFTxiEEJ3f+1vCv6QemXW7GcBDzBkdK
gXAtPd57w0nfK9Qt6wE4n1CS8XIZAv6tViqTMpoKalX3QXXv3mLeO493oqXQ3a4dCKYup3QB9zBV
OdW3+xer9UnCAI2vkcGSj5urZF3LObibid1eacb7KYtm6KsPtvZmh2f1FKsWiBGecMCzOfoE3cnY
/J5xX6hbnTCAIBaVqfUiLh6tmf6nPDjyHbDKfnKacyzzLQ+Mq7oasj2C0WLp7zw2d7Xr3DlxrCWw
EzGIgo5hCztkj/6i/lqQTluzmE0UbWlHqWZDkQW5BM9AERXnz57exml+msOCDzcLtJMA1oS29R4+
C9TAsi8zgd2iScfTrj1xc0LqIEsCRuhkl4TN08XVx97wKeM2+dhYBwz4Ljg+ICgU8PeS5c5Yvkc1
O6HrKOI/6Ks4LSPqJnV7mawYc0r1ynCiCzp5zHRFFRED39wsLqPUXqw8Qefdmxa3wgfgMYaommMa
1uI8M39OBEYJEUW0GcbdQHfDJqBUx3ha+6rGicUU15a99DYNSFA0Y2XmLRLeTvns6Lct+H5kgUa+
5jYfent9ydosliUuNqz8QnwBSp5D90MBE7lma029Qt2Q6cEIE+NO3VHE+WIWgsasJUnCgZ4AdiNO
lmmP46wJYqFZQ7btE8SAjuGvGRRxelwADv3QmQBO7fRVyjbfFzH2bGV50Ob2+Ze5hZjv7ybURFHW
m9hhPS84RYBCzpJS5bKDVHQYBylqp2r1R4Tj8+THr3JzATjSezCo1XKHL5GplJav0c1EUEAB9RCD
Ys0g33cC5z7hGGKNujJ5Rbekx0TLxITSHDTDQ+w9p9+NMjYADPD+5WZ6vjmKUPyA0VJdmuk10eR0
sHGXRO/OnQ/VUclWwooSnUM9K69Vx5hN1Bp1rpQIjZHe999wsXN9Ek3C9NvjBGzY1wmqYv7/9KQM
TGxVqr5c2P7UchV7NOSOXkFqjsZngwGSka51d/slHKwlvK7941hs82e8tMOCRdU0IDVls3VPNhUT
bhDeJrniEtth+pMr4rtHZWYPz3fNQD5wgaCMZtlrCVpMG/zL8BY3bm/RSG8lL5FRL+l2QlNNksa/
9yVVXWKA9h7VwHNI3Nxy2Oj9pATM6QswpManbX7yczKffxflteH5wdFp8vCMiVm15uFt+x4W/P44
Vr1oQgMZmyFEfuk0XsqrUXLIYezLw//0IEsw4wmsGBzMY+ZXD6qFG53RoV5EGGTkqhM7njrI4rFA
FnqPC0Hv9S1PeZTabm7uDXrCKtqpL+4flA1wSgTQLCYcslrV7PsEcBY4IwEny/Qd7p2siQq40QH1
mPJqB21sueN4bi62v/aHoHo5cGcCE6230bXJ4Z5U/qHipXFs8+ybhU5F3qYzx5koGAg791/2s2tA
EgQx6QZIADY7WJDYmFR/B/eMR47AoXCgLkYQ0d67NgpCAdDmPVVg03QIBwXX396HBa5eMcsW49AL
qalVaeYuUOhgBEAI4DZAOJobQToyBoHP0RtxLpqpiimZMtm6pk2lIDYwL+/TvVgwzXnxi67c3kY0
VCsNIF3y593FY6NacbTami0J4TjVIqcwjgosLkDfxy3MvYGi0jbVwv5LKkRfNeCFARFhdsAcV6xX
6zdQa+2R0/Y1cv7/gU7UxAPOjLH+MmarIgunsFCVrHuzcEVu/Qm/QYOLSqAmK02fxZ9nBaiUAr52
MnpelaIflIhueuhu6gfDdwgxaya0zsGer5ECcKrWwb3HlNNBtC4K6Xmrx7AhYpzTTz12Vyl28q7f
LPvIgUbgeqhQKrV+6moP6AhzxmATSrnrCZEJxl3xNHRP521uHzQf9r7tku/rszzkYv9WfuPTF4rv
yGsWJc42mavKvv5Z2LE9CEht9z5bff20PkFUYRO6pyuJ71Un8NNfeBgLSqYv81PiFJqEfTkIiSZu
NGPOs+YSt1ZMvrLdajK0TPvzxqP5slzm8Je/XMtYyt1eJL8/KUIgRXavR9m2N+oc9a0+IXlqzeOd
hI6y+mIX+AFZMtWeg5JZrZG3beUKoaLxpC8SBrBasoZJg99LPEZFY0myDqLb17MZOk0Z1CeH72cs
L24uVewe5nC/H2am7LCZ0V/4Wb8bVm2hh9u3mvuqVfjZuMYREZoSfxMD68VPu0Kld6KzAN4FYoXs
53/CQmO7rQJg131YrE1fkn8jaySDdoCIgLPWXdBLyiOYVZTisJ6u8ToYvqKfCTd79eC2dPyCXfl2
WuflwJMSS/lpD5tVwmD3xeB9SZKt6lZj4o1AekXIrfxI8yuezbJsJQnr82klqD5mCWGHGBzCs0ky
Ib/5qtbWZkdn8s7vxvg9JBSzmRDzFV68O8FzgdlwhNwNzj65AGDOzBCFtTDk+t1QtwKKoVnJksuj
6vexFbk94o2fm8ODBM5h2KVgFuBXvNsN/y1JPZD0KVkvbCunBUSeINCJLm5ONx1fQSWWr4LzdYar
TZ0+SRX+pm0uwcWqDOKum8pqHJ1gly65cOmYDNOtDwgfQWGbdJGJYgeYMOtSBhf4gAgebPiWvFlo
HwoaA1EmBnUtcIilqAlLLelJ73ldSkNuPsb/7WTDYwg72sZvwnWNLecvkBiHiBFjRuwZB12pUPwE
uBwGtM1ETdnZN5oYui/imGyaxlNx4A26OI1e7TA1d/SeQ9Kgqdrf7KLJjEEr0tZY3aHdrbE4kYb1
g0sxEiSetf2jFF8AZPBE+8/wWQyNs7JjGlQJsgcLlCQQDaQF/Otc3ir+84j5lpJyYO6Wwlm/64F0
us6okTS6T/y1CNiLCFFliR7jFu2mjQ9B+udiAiQodWRq9mJStsJ77JO9xROfaB/sZLlAFctRS4Jq
RJUuDS1VRygUAidfymZVKJkN8UxtLD3TjqcRTX69sS+JcbedpqhuxnePN7f1iwa+YIvKbqV/2nfQ
TiLzU/Arkof4+pNg1yjUX3mMQWGBqgXfpFTeGGF2Ah7imH1Lp6E+lm/25xztp9X/wjRUDHLj/NJv
+jkAh/jKJwGXtLH/vYWOD3ZlYd5EULHgV0JgXkdkBtPa6JE3lD2TLEZJUKIO/FkljQVUj/tsKpcT
Um88+weZTgriM5rogR9iygjz0JM82yHd0wEGGK3xDl9FmUgI6m1c3CPLyNTFJgBA8G799+5WPDK7
rhzDD9VS5Ov6O2K6YaGjXmVeh3kumuzchK/ARDeIfPQ4fb3uaOE3vmj1KEAiBSFH4YSBKfAQZCVu
h4Ek74ejBJlyiFkhLD4A+nijtfkSHN8592k0I+kd03effEbj47jFil3CLQCv3HOaP8wNPMvlFXYl
FeUjB7YD1s8bShSDJ3KYlFx4Q6BPDyVeO5JBxXswDe2A5l18wdBBVPhbyF43rGoisIL4S7GTB1VC
pcPjp6lkD75ty90Pwt/Rb2TKbp3t2xur+xK3qi7YXCFqNDxw7aY+Z+IcsQq/WY4q5BsUFj70rsb1
w4LJWLVhorCM6ulaL3xpWcnIggCRtea+IivkjFG9hyWpKaH0qQu/p6ENfxwTG4MOZmiIhlQlSCy7
sAwQb2iRyEg1EJMRTIZnAN4r1ASY0jU/aJcmwJNRoWadjluuKYbMtSzFaXQcEwF5dBcLNoY+UbK/
7wfC04A9b/+T6MFGrMcMg2Ht7tCD8zBU+8+6tE06pJBBhxW/KZE5bHvy7PRf8ae/QSVb7vUx9OlP
yYM1UQzczrEHTV00udjj5hjaQambc5okMzqV5L9frc5YnNw27wPaP4BH9ndhjTUPQS3Znrrpt9Jr
JOsqrecvznVoJcjDJMLKkt8uSnxh5Z58DTs+HVyGRkj91+8/txJi5yb606A6nr92he42Cf1YTxgt
sRq/ceb86VNr+UwZbMjhoKhXwpaMd5tN8r0WsW0kPxALtzoLDl3iIDHdYZ6KBnKT6yJvHpbt1Jpl
9DjWrasXMumwGaAeSRTOmW7lSexagpFK5aYZQTvUu0Aabfwygr0kx7pbfCpGqi6kJfnEmIjajYyR
XH13WpLAgzDKhLP0vVkAM+6w/d/oeehADQnIWo3JxP2pFlGjxpYQOWT2MBwvrmulrAG4jz6iWKT2
RMASUUdrA4O7CbO4H2krV8RF+URAko8wdNaXps5AGs1W35tx3L4alBlkLFzZJiLMGuYmHC4yufSB
N6ZBx/kHyCcVjEgw7XozqNtqVVc1qrXHZYW4OE7uwJKY/t23HwLN8EFuKQiCt3A2rnOrSYxBygcg
cw+DrOsLRob/Ri0FnpDvqI6Z7XhkGt3O5/ssmXETmrrVZ1S5qvMIge56eYTI3G2/CZ7/hUY9ajfK
3sIurAd3mrqN5cpW0BhZX2EL63Vp1qUpKNH0/K7PViTKEi2E0GuooaYxYfnzwsLN3BwrVp67k+1X
wLK44nFZtZ/s2bCtBGpVD4tO7wxsrANmfzGB57YKrYlBHUsy35/nlp6th/Kz891t6qukmwlTD7oz
JFBxBqS0xLMR15QTZl04Q7hnKLIxrH2UgScdAFC360THUS3ImBXlsYhaKKdwaCtZ2TzW0s6jNGbo
lNSjRzDeX9eY+I6Q2RJlQc/b8mGRE9g5HubfOcTkdzfI02ryje7BpDShnSYsf/4qTBDHQIxYnPFJ
yLJ3qDLM0p8WYHOF+p80zqqeooXbhhKT1HDoCLw/t0hyYzbAR4GBnqQYJlTuKKemqM4iR0K6Me3Y
jVtMkf8EzRxZQbtKFDNbhIzWkts8ndwFi6NrBzpn+8IceHmN1NbLGko+dfxtU8fHcTV7WtjE7qs/
IOWRlMSNM9cndKLNBsagwGprNs9tub65euU5Aili03J+IbH6e3vlsYNZi3sVxlGAYNq7Rp0NgljT
qXiA9BXHyqqZE5AC2pYqpkQsi3yv4j8h/u09YSa8R1IVDl0Ys0ZBwdOJNUY+lbWGxek77mKvaBkl
uCbLiqiwJN4jFmdiaY3x0q0IMHzCXokZvM/nzyatBx5TQKR5gSFnsk6hfst9q5DvHMvcqSQnVxaq
kuVhe4AJHIIvK6ILEK6RU0tzrszuy8BdIJlKcvs2/VdGFEaARLxxb91JrYMZncUIr/oxJj94UKmr
OajZOO3J5cPG1OGqd0L8I5ti7gMyGGAmSb2H5P66Nz011pTtXIyRkFgRRHNHWdX8ELYT9hgOnYJd
kb6kRWrU+810LvodhLj37DqKWuEGBSKIJGcBq7bbe/orD6zQYQlNeb/R4Z46EaRVdyyoV22rkH4P
9JbZDN9kQGCIBD3tGc3+kA8sPpTR3TE/5dffKEJTpcW9UPDz7TUuzjEDdTVg7E3ujnKtdbkiNyZe
JNl/xxgV1a5Lq/DLja0JZYqZ8k3m05x4FIsNGp31apTrefBLL28bQ3scPBbJqDU4m+/Mht+Rz66b
DrUSkd8uiMNCUe2u4ThDjGlskTYI5/51JVvnj2Dne+GlhsM5VA3sBlp0rij0HEVrGAjjXmWZBd2P
WL+Jmt7RZebLJAGlkt6jTnY5YxhNWEuEB9TPHMEwFWwgl9Z1UIwH8siX38ZYxpkIM5GWMrb1nd9n
VtXRmtDgOA/L4kIO17cdt7qZGSbRVYgTMUX4rZFfyfNYyK93jsLvH+eYMoTfY6uCJRRumGRnfU6Y
QF9zJBKFPzThPncAfkB6G5ZS9uHsfajQm7Av20+dPeuF5jd4b7+xXbOTEn9NIG8HfAn2Ya7ixoYn
1EW3wOtbfC4c7yUJBGmgEj4w9vXBwKisgJfr7Ix/onmM6kN4FysI8tU4qqK3/Ta05HNb/ucKw4pg
7S9EjTNjMedYR//vJqraYhwpGDGNmjj0v7FXuL1+ZEeohgPVra2tcm6nY2/hXcVOw28Xqodt4HLj
oiGYMOcG8j3XnjUDcORgdZM2dglSer+sqU+xZDU10TFOGU1G/E1w1gMs6lSk2Sc0iFBz1TbRnegN
CIlkthcOBaiOwcHDwkOCex+/j/27tfMZJfV6YG0FEnaN2MfB1B3VU5Q8E60VC11NPUKnQmu1DYyJ
AcXGLQARnFuelkS7uuMUzc5G5MNPiCR0lo49oEM6/J1hAtLkwoGcJYif9AqtuCMWJgmN5CFFvaJm
nQ9ooRg+GJxzUnGWr2+nr6KoG1LjaWTrHWIDCrus8ATNz7uA0jsy8Q2Aa1LEgCTg7qc3kjkVSkZJ
08yvH2RXYRkpZi/6TWf1I09yoS17xwMPWNEAetCD4hat0bQwZGQ+ix0meO7+jOp7v1WhQ/Ovxtl/
mbXHvUGFRa9Om98eej3gB2KMs1FpmMKMY0vni0mI4Y8fXTZH2VNJE8ntjnM4l7u2Sm+80sZAUU5S
TyB5MosupRKYLYEgLcELSKa21/FEEcuYrvcgonoPljUwdPHn3ZOay4mYhLBq2NV6sdzqziwnnrVm
xnPP5euKhr4RKGAvzAaHKBYfdGSJ/7ahomxeng3qt9a5dbny9RcCOSILGb+qbMf4JKUcwFUmeQqp
/Jd/rYS+cLfj4L0D3uLgSpIkLjuKJJK0wUvQaQV7UOD05ZGlbRA4Y+pxzGi8mULCjoHmPg9Lp1Hz
+Boi9XQZ6Cf+Ynzg+bNV9ek5qg0ZtA6Qkb31N2vmm5kSlYUFqHXcSuXBT4ZZFaAYRYYqzmLV5B2J
DJ2bTTbQni+p/btLUQgwgLBULWXWTyKxCjjuoBj/O0v2C/BJ9+vtQHi5lhlcmLI2Ol6d54nmobzp
d4LdZNb5NzNd3mApj9BPCSqYW4nf4YWV9os+AyhO1KndpK7rYAlu/8HqawZDd4Wcallg+ytcRLYt
emNk8kqBy8CBa/A6mqZc96VEVefq2WMw+1F1+zh853U/jf2KhhVQOl+jqHADYM0cdvjlExZAjkiB
PJ6NXY+GTR83Sru3nnXV18lod9tMY1WepFmxy3Md+rUjPbXdnyVEJ4TkgODdmNwmEOKJx41Q0f7e
ANMiTphY1UjH8DPqNKOqv5Yntq2IPl1eYzLhbSFGV/XY+SvTV3QBD60HpoXSZOjlR6rewuOOnmGC
Wm/MPdyjmnGxNwcWZxilGNUoTRfbMT84LZ1lBNYfslz1zYeIi2mJQ4rLuQgEYQaZo/xp3HigKU4g
JtO+NQvtoxCGZTxbS2Xt/diehmgLZTChsmQZiv9WI9XtMBgEIQ8nJmjaSdYIm3lcLYni6Y1nh3ae
eXNWPtgkJVfBHeBZDLWkCy4IaLhptyfY01kbzKJGGATVf/JPe/ANDAqjYt4hNLEvXPJ1Y+O0+cd5
/HsnBQ5kX8HiSmNcdkS7MGuqBrrSo/8pTEyslOaMcVz9BUUeI1atR8vPRZo2qZiJQCrFVwT3MVrl
zC1KRC/cplQzJeE13XeU+ZG85XHksV1KSZ+gTTh9KITO4twNCjDzdrCs3BUwlXkLTt/Ffb58F9Xx
Nz6ZKYyG3LSBWdC1AU3xiDVK4lsAs/TfdJeYiGA4FZWzOs5rRmumH2m1856hyB3dMKQQeFCYCYvD
/haqYeTjQAGiu31e8PrnZIFqN/TPoAyNjeDJmPtUzl+4aiXCqo7Qbcmc/t4S+muzJcTrxxbo33vK
OwRqcNS4jg8p6vSh6H5pLSwUvwaceZ4SvB+JTXJ25/f3UUb7PhL58B5CDm3O820v3HHn02w6Ehcf
PCCFGbdwn54FYgJt4qtxUrFdMLBjVdA8ZdN+A3FSP2YgTI+RfqpEkvVeRqFeVKMXgLWoN7DH0ohI
Bl6CJ0S/mI+mLaOKbF1v78lvnVEOI6jA6vMECSa0mH8/UZfZ4u/1EllIUiBzgUllgbRGq5TLeBb2
tSl9GuJ+wiyCnmXlxTpD8Wo8/PDfrXlFGxh4yu8zN05PXyZBuqRFZEfonlquUIa5ktdklrqvtFcI
w1lFoxJh//di73b/Icjq6frLsGr9mx5d8TAxxgg/NC+l+RicswcFnRXbmWhgrTinAKJCfTekzC2G
Ax27QxpUW98RAgau5xXCmVH2KEU2cyJlkzXbJ3waripweiJNiNmup87zgyRGsr+tWz8IErwP99tH
B3lJH8iFM1CJDuBs6VajQTCRLbIXCl78e0NJNk+foF31NZ9gnwnPdEIYZPeo2xBMrzwP89LP2Pmq
8N0nfWjpswzuHg8ecqCWz4GJEwhuLULCYSO2kPfJ8ywcRJWpnHHWce9zKa+ceFd3EoNc78UEIqNv
ohUscRoKgSQaQLF9m/5jy2nXvjViTH2vSZE/36wW/9NN3YF4RNrDGDw2l7tdazUYLxxGV8QD09SS
5QT2B4tmGD4Ut3+HT8lquMcGcVWsoD0z0XYVUJj5+i7TY778jaf4hVMB+Vlm9cRiC+GH59ZVPXkN
M9moTr6dNF77joevZBsSMBc6neeG8M2UizLysZlZGEiX1IKezjEO82RjPnAnwX+rgj3b9ITDXpvU
S3GX4vSUX7EILJnV5P745Dh7FCa3S17qo1ZOifoHyNCfxMDWAQV9hW+8hiL7YD88KqyNprbi3Oly
EeQVJvlVBrCbz57mHku6oFaUvU5PR8HtHMjDHSpO0/UfiB/Ot42jUDn4MyeulK48pD/NdeUvpQuq
5AxMn6DAvHZQTP+1z+0n/PqOA+4zyGv2KyvepYQzvPmUhT2M0BlDpipvZJyW9qVrBNh39u7oAo16
O5XgHWC099UFPivv8SLTAtjOqvUDSmijQjAYVuwfgVwLhcsaFRyXJhDdd2ZdcHiHSVuNKxPaG54T
hZFVy67p4GoIVkJ2Y+UF8IZLzccQ4Pj98pMw43yC3cMVYev3T3m78ycNyHJGfIs2bvOoa8Dc6VfZ
6eGSut69xaIM4AGil9vTpzRiPNvnDvMG1fuY6eqSGdlmfJykfxVG2gWyTnzwVOEV7lR8V/LxGRZb
Jp01XT22gAn/Ms7SAhapJr75QPpdismYLgcCtyRKg7363ia333Ejq065RSVdB6qHGT7yW3l3A8N/
f68ou1CL2ADn8NimoQdDipL7GdfwAm4E4MNpApJUQUzHQ+3qZ9zg89wfqfhzpAEhU1QFDnfKEUyL
SzLC0NYbqjmdDb+h4XMOTQ/N9x643x2V065yYwcHXtEsCLvVoVdW/UiDIsvFhCW1ApPvOBb07zy/
HqR2TmTT9wtWrBmlHcJJyPO6Ney0JPMWPIs/z1AmZg1gkMn0mP5OK3Z79mb6aaKo6sIdSviBBYna
SubTKbxqhU9slZhfKYalK+1vBOMmTONlk43vKsbkZgvmApkmb1jHYQvYHCA6vo3ZgDjRyYJN87cL
hWwOlDuV0KmQPI9C5JCPYYnl1hyiyyxGgZy+fgVWGmQhaph4K5tvi9m4BrSC5Ijt89G2L6rTSl3S
ayRraZAPWHCfj9XoQTci3bu0rIlnLNJsmX51gnCtiU5maSgM5TiRK5fuc7uSz1WT9xhaQohrzc1u
WcI1atm7EPa0D5Z3eFQZB/GwyfAdHN4uywDM8/JS543ykHVDKktFFbiPozKLl233Rwlio0n/EOiL
mMeLfR85UW36b7R4jRRQRSynnjxDcHG+nSSZoFbnSjvFyw08XiU4H/mt+Z2OD103kLomEbglyMjB
BA3XcCClbTshUAnWCqVwD/H1hU4uCf1EEgewkWXUEPpY3PFlWFDIU/Qm4u6gMQ+FIeQq62wNg5yx
8pTzcHclqjCTBRz+RGNX0O0Mrps7yFtjaHe4tVjJq7Bv10p/3Y6yRotqNMTwFI86RfehcC1+S2gJ
YUzAUGv8vdf95mee7uFIsirBVrrVWMzNV2FqUtOTwDkw9AUG/R1uDWKjBRGDxsFVn3Vk8/2ekolG
GREncBh48Nz14ml/4dggsJLT+8ZPO6JOF8D7X+vnrDA2GNGA1OnUVhiPtQNXmZoAGnIbqG5sYGxA
yI5R7Brc5Uu0kvwOz5hBRtv4kG0FM1u4pVnI/zP4oEqKCOmelzniNcqaoJG1tGG+1ESLyZwSCJOz
1ExaWA3tQ2GDzKCc5ZAUNch3rJmp1mbmXblBFJjYpNpFbjIgqLw1PFWD4MU+l5bTxfW8rFOpbYRm
l/9qg91hJmsfoZ1/UXhfWjrYPKSQRyS9drl7j0pSjhXw6I72jxogZzTcuvVko/ezTVekDO0zbJin
cCeADlnhCV+AWQue06LSMHsoBy8BxHdrB6CiPAzs9O+A8aYEaaxmWWCZxp9q37Y/GI7muJKyJSGx
hFJuEg5Im1xisu8yjOWqv2l//9NBV1KwO2qZLriPpWZNTU1MtQN3rFEdy93azy34nTEuwhJrehc7
X+E17WIl0twPRHS+7goBNozeCL0Ta9KSTiLnTYygwqhKjqmi3OLbmLNIZppKFM2emENothcsqo6M
pnFpeSZ+4whxf9oq/xIDv+D5KVcir0pY+UajXPKUjDgjT5dTs3gB9WJIbecvFwYKLkc5nVd+7tRs
hG05xq/d/6DjKMK+7zHj+SVK223R001IHt6UHW8BLKRc7JtVSCabxqm7QUE74MmsOeULo1m+az0G
5X3Ja0lK1134m3Cer7dUDTBxrRhz3hwkNSQQpmO18SQQ/ejbLXfJsdATUkAXrVKgU0VtzOfFP7+J
8zhEpAKNWKubsv9navqPOMZat82cJR0ldWeNsdX3IO2oqqJtDVFrzBrxs4rc4w3i5z0LaEgdpP9y
/vn7hn0GcxTFa9uZPEqayxvs6vAyeRcYs3Ow1Tqr5ikIYtiSC1d734MFVVtkdtdvl7LhJIyICLW9
SZIIHOkb6udzgHLpzpNqBhqcE+AGqOFLdiArhcxy9lCxLCh8YlhrtFGFJFPbCorZ8ktN8q/QlDdX
SeiMhVImpE8i9d+phlj002O9B6vFkV1qfrM0YaL5i+RtneA0GIEIFq4tpV9pUgII1VZ/24aJsMZS
QtmqyNUBaNojcB0ZHWYJ8CBMiB0pmGrEOSLNc3sM3ROthfBZlNNuaXL46p1JcY/KAKH0AL0H5f0y
iZWdllPPYCIBOoCiTwa9EusKVnjB7OoJ5DXbDnjVE5w0e3X/2LHLrPqHUGbAkWai67s2LSZL9OYi
d8p2CVs7ClVl8mIMrcabCRs3ct/ZYfcT5YogkC+se2LdkVbVdc6kMLzSrFv2yxm2KWGRE7nVdSAf
mOJALYwyoyOBtJmXY5fjCqmax/XD4gIv+hfErwfpmTKgoRh/cCSZobNUCdeGyAx8A/n96jYzGvsf
41coiY8G5Aeg8DGcK5/doq+4Ph3PrtsvZ0eRmY9T62zhyGc8I/rsolCF9SGu4Yf5MxGDz9h+ICAz
nZpkFoFhdGFr+eO0v5Nd2HVovUyoOUWKKcaoK1plvBmSw6ZLnpjQR7UP2+SEBPonUAEZrdCwfC1f
1YVK+UTmLcnjJoKD09BHYjbH6a13ldpI33DC0puGxOvNagpg8jUBF+MV0QOgIrUlRy3cvbWj1iC8
/Jb7eTB9AxcPvgwrw3oiMTHbjFH4qTcnJS9y5jpEg5wAMj0P6JnxlVr9CjXKdnykWygce9+vNWVQ
wfwAlLS8MvfgzZIujWZv0QBWNKS0QoeXSA5rH6oOyXXVK7GJ9/odOcrJjEcpgQnoYRFFgvRVE3KZ
6scLMI2o0VEvovWUvVOKopGS5xQX92QAJq4cYdlhcDqcmN8pFaWG2ue1md4qtB8KhMCBi6wMbdjz
k1W0R7y2KRFM5p6v5JVPe2KaXFRWrnhiSR9d5paowEz2fEHCg01CK8awSBkwY5UYb/j7/hD6Ejt4
0UtmhMk/dIioePgnq+a9wXaxBQUw05lqS3AH0qCcW5Pb+DXtpY5gsOottAW5JzFyb+pps39SRfn4
mFvhhXxFBRzSPMLlU2lQApOkuIlKDN8Irc6yEBqev5kwFQQPYq9nz6aEBSVa/5rvsJZdYTnaSJLM
tdQlytW+TPaV6WwJimWy86C+V38ZiW7Pr2G+TB96UbZ2raTnpNNRKcwOjrVzXfkp/xCUff4hoVtD
x/wv2MD8Xj3ThGT1V4hHkbh7zrZBHjL59lsCqv92ouU+idztgecpSfVJnuU2KD0bVhjoc9+5ocsp
JSer1mdF12qsPoEH5CZVMP7IrD8wddi/m4S7/av37M/C9ja3ALTiMl1NnVUBqNbuDQ9FK36tWuF2
i9y5XU7bhWwWPiOjApqPJn+jPR2pbQ4gFoMC31Audc4gq7WAVETXmGzXKYAH3kFMQlV/yhFVqgte
KcUa9xiMwNiswtbeQarA6Yz/V7XARbaIB4bEDAEoGsHEwHsBRHxCz1zI5rrFmIj1PtFH/rOYoRS1
Kv4A51LheFxjk1HnRz4YnAbqm95zkI4YnP9KenAlk27zVpQMf969lzFVbibAHamcHEkhSzDbzZs0
qxByUXKrvaCHJ+VJDcgGmdyndESvPqrfzyjaPFlpvxFDEbrlvyFoKgxPp5+rSzdbTdJWzFSyrLJ+
qf1u58dAAPQeXCSf6Hh5YGKrObLE7183jmzobKBvc9OoyDv1po8JudZmN1syb/A9TCUUvqLKTti8
BaReyW2GIqAtFMIy0ZWNgLgVpEbEzFr+d3A7mIp7G/8jkMwg6nn4C711Y0iybOjD1RuKVBtTcr+p
GQqQjg0YU1qYkynaMWcwfIln5VRmU8K59BaGvnzczYSeKLrahCFg8AfFMDlUcD0t0EqnOPvv1V4E
BYvN0V2qqt0aaggOdMiEnEE7jteX8VMTDHlM3Jwr6UwkKU/jZBsQTyawUppJYMhCAL9vXhWeqK+P
zKHREh+B52gDl92Ji2vondIyNUxRqMLdI5/oYVhRC7HM5rNPMx5E28xg+Ao40PJV+DnoOBhgNQcZ
TeFx27yDj+/FlRjopqttAUh39WRo8piUPVjXI16wba98Sn0ze7XFlGOhH2FE8FgqEGuoiuhsTCPs
OzR1D8LyqRuNsexgIwgXQrzMpFlZxEWF5100YSPzvkbHvtGzrFKvWsxAcpo4SClu1qVGn9E9ql/j
5fXd04jlfzpB97Ps9dmPmqybG51F0Hfnx5mpYLNLmX2Onp+/CcamlTXOk10qd6QbGW7N6iNjOAU/
NXqGEBWXszR84sYruVAEE45Wmah7ifBsxJY8xPpsTlFRgaGbqMcn/f+Ms+RQSm92ng7506gD0BZ2
tBCYxRDtuVyBRZmm4d7u4CyRkF8qefI8B0iapYsZn6zpstzdrqF7WRsBtUlvTOjX4YtzX7opSxOd
G8s9vSvwFJTKcd69aMkBFc74ZK85iuhQSHEd87dDQoAf8BzmDAgkDugA2zPH6G2t8OY1FhLQKA5C
RoM9VI4BDvRq3Gp2kaC2RymOtxMP96NCe9O0PfX7sq10P2outg9phyREiTG6rXMqsWdU/N1EmhDG
sgYgMYzGoSX6LfXpLHCtgUK9SD67qeZYe0T9NbXjzbMlFwGXUpvfFOi5mB8QolONvESXmLLJcEgW
DzwW3ASvw3qHtljwRyLx1VOWnhr+7nwxPBG+j7XEcW8nOPzzu6c7qFLT2lkctb3P4BwTcZ8yXiEB
+WDWkRTPc9XQo5o9Mu0Tyt7wzBETZWU/jhjxovCPU5rf8yF6TZqWr/ybDxX32hitxlhfe79LemcZ
OYuzmQBolQiokDGjoarg8OVihbkXI+aPwtvRvg5cNrLJVoTvd1QXx7TFBbvBnQzjEFnDWzoPTWsQ
sJBUxZ5JFqdKkuHo6hbb65iQrJiGqcriWwn36g/WAqPG2HQpTDDMtorg4inuS09KcBl1n4iWivIo
8ZwXNfujKMNR+Q0P7xyJLLNvXRon2dA9TZey8f9xM0LfcmuwY41/uyu1uoy7/SP5bH0HNQvL130X
87oY/6akYJYSF1Ih+wYl9YHPxO2nAdkC5rcZyV0OSlo5XS3tBMNcNiHZC8RXcga9QRpw9gfCRqPz
jIMI820Q4kefYNKkaqrTNv5Sd2TMZ4LTSvyVplkxaHvWlWO+4QbSIGPjRmwJln1tvJUz9/RCJsXs
XHCbGlwzzImmYMLxqa4Co6awTwupl8oX/4EaMljzc7OpZ3RRVEcvAisDaQjr5jFfZjzs4tridJdW
BSW+P905fZGW0j+/MbzWLAAdhCPDq/UUxq4mcTt7caEpljr4xzjPqmMxWb9QxfZf4+fr985SPLTU
P0Z8ZMtxunCHV/sG48aoSHtUhljyyW1PI5FxRodbJZMW96lYqFKChXhqejJZ4oFrlYG6l+/dIm8u
fZQLF3ak3/XGufgXwHr1D99Ygpy+Za3wdj7cvLr7ST5ZFNoJa7fZ868ry5e2tH3/fVlUByBYrYbF
pJfdB9hzyWuZxbbaG+MTkhpKrS7f1TWM6/+Lr0eC3pOUYJpVBhfJVfSOcUnk+1iqbbJVK5Nfeivi
vqV+nrZBTdr1od6Ma9ot2UFMDafPFyOgESY5yYciN9yefa/ZPhzIRYWDg2EF1iAbuv1YdkE97/5R
wqex2FYTiw9qvDeAksTv13wLHBIiaSDbaeCcw+oluFCN98YnFsFcLwadIkJ4IAhbasIWJCNslytI
VBALxu2aLGyTRAoFxLTngdtUe4C7bJjGgeA7W3MyMCTKDg65owJOe85TPF5/Qrzo6/XlElprKqlZ
H0qK+7Hr2ULHUg9Im+aJ6RE7dvMay2g8+ddXUELj0XxAffq0MyDo5B1X3ThT3X+Ihjxy8FXIbQ2n
WqPYs6ciqw9kz6S4pZwhN56+5Tso9gwxtVMUCOhWLa2l02awzIh741noxeyD2L86Ljd+edLwP2VF
L1aGAPpXuNO115GwuXbiZBRKX6IuaUyvd4Tq9+lj+a1y2NXQXVg3AFuUKRzJNKFmXTiKSdTtfHTF
dhrMAcEynTUtURFbpRy/X510QP0kDXXHisPcniLbP4hh+vJ0bvcORRRe5C328BtomIfmp1S0IqWS
ktoCr/9X0f06L9/NouSM2jVC56n16taKNp+N//1lVfoAy71MfrDkKZK4tG/67J4qOX+lpWkhM3Lu
VuxFycjt29TGhF9ikghNtu+3zDVE1/6KgGLuuYkL7oH8BaZ1eO3E8hWKaQ8EhLOI4XCRgYyyJCgb
DGGO80HqLK9J7kogHBsqEkGcz/xpCHP6ZdmeHMzMqLk6LFqTiaOt5wvgAX65Nk93zYRpWEK0lB6k
sOKHgS/wdzODo7NjMBINjJvd3Dzgd96seZMwpF5URMoaAMfPYO43FJ9rnTblLcoBVr0dHDAa8JcP
fCopdkFnrdh6fVEKJZ2LMk0Eq9L/sMEti2QqilDPsgBp1elF66F8kF75cg2ieGD0rHnkBnlq7hPD
wWQ3ikLc2fEMtlaieUenMovxjL+k/eRW2fwEEFYXHS34VqtIPqNJUBVMB4MmV9W7W91DmMQSgeO8
8J7ryVj6oJjHUNwlbQIemQoNS3jXhcKYZlRWOqpEwyrwc4CKgeMThmYkz6RVGjalZ6xJQeoFO2hd
Nok60MeSKbz68/neXNM+2C/e250T94IOJKqtzKr2mQd20R1G+TdGYgPE8qIECsnx/5aENk1v4y0x
RydEeLDkNq9+OykTAIAwVh1yxrlqtG2quPTDx+T0O4Oxc1ROXutu3+IAUT4QDUadKxgInmpv3bp9
Zaa+dyt1ldxNuWfMwcilTryC/RKRZTEIbzJzALOZtxSrw67BfHK8OATJvoX7xZkTY/f59q7aPXPc
rnWIuZyixXaDgdJYLFRWOTog4JsFzlQgjR1rFMiRkBBnNoHanHFLozcLTMCFWlEGgSZ7LUOmWypz
wlfs/56ZQxHF9ol6BwKIzKTf8FFqKqc6CGHPFmRoRLR3QMp+WIH0v2NvSqDxa9BNVo5aZYplttl8
JaD9Px9eITw2Y6kMdcWBAcr28frXxx7gyND5iDwMWKShvhhkDQ8bX7+MDWmZOKdSATm4EUwhIm7b
FYQeq3nW0FzedoaHxADfmupXmLJmksY5E9xuxDNYEwSOoEMqTHj6QxMaYzbBJZiY4jfBNCARkhnn
mVQzWM9qP1/ol3meahkI9kMWozwMz3+gqzE7hSzKGhRZu60g0rTKyoj9kesgtYHR419+HtvYC4y0
QjrXzg6LL2xcG+iBhDYcd7Jlq8RRbY1kIgMexEzPqourqQHKEisT/Ad1ANBJmHkg9mtCwIEQsDev
6p07BUCKrUCq4cbUkVzeR73iRb7ahNOPTZLsevWS41EhFw2dfs/+gv7gcsAa1OzkuvKjg57NkFSE
eiz0dn+lJ1smmX2lSXPSF0Oj3VCKcyPZTy/t3aQT0wrqqcwTUcFe4MQTqgeI94iiKEJ+u5EWTyJj
Jo2A0t6Nyvib9OwmWgcvGNwaEQ/lK3T5rAlvnQ4X9iUPJ8Ex9wX2VpPNWc18AkaHEWPWVPP+/YPb
mys1VcpNwKQLKnumuhy9iV07fuC8fpJw1iVuWejwFjZWqe1FzwAJ2XGR1evmuLkKcvCgLv2vxJO0
yAlSmu3l6lEcXJ0T7g7jca2eOZoMSGw87oPfpfWHskwUB5B8ZqgTe3eGl38H1I2TWqyUfB0CeL2W
P1GIDtBL4XglBvv9EVrJlzMoGKNQUqzM3biwy/bUTkYqkcTb/aykPFsRAYseuOd+uz04T8M9zV+A
tGQF9ZfHP+Z77zwhdeop5J791OtD/sPNiJVnV3+Owv9gYgTAl1A+wCHkhkuUNKwN2d5mRTT9roeb
ok0s36CukidpDcXgnLTXA0CLAgqcp2KwQNVV/cqczGNdcpyNJy3hcKz5x1qxaSwA2Bd6DHRCgJVS
n73N+94eJ4ELgQ4lvHyFmv5kw1w0+dBa7dDA22IkFcPDmldL+HBSVmxNpgLCvb2fgpr7U2SMpq+3
yw8cWBdP1YlbFFEMu3TTNlQyzMkDo8gT4KCzsTHHjZb5GBpZgsBLBLKNl1ysu7W6pL6UhYoxNdS7
Q3f8MFTwy7fEyjCEoOQiLTdagxf7HhWygUosn3HFd923EUl0UFD6knWKThSNV6KX07auVxDqLjIZ
K0WwldAzADrGL7DTOVee+46YDcc807kHGFDGgoXcOHd4/IgGX6WSQ2eTMHl/tN11pV/FOvZU123+
JuQbn1cCQYfJ4XeFQ9DkZhbErI2yVtG43XT2PSf4SwGHTfX0E22bVPs/8zd2ofvzr3EDpT78dm4t
dzRDEGvlFMFWnymKQozTET8XMSoe2Hy4Q3/AN/gAWk4OjwfG9CidjvEjpm7IE5ckvfpdCUQEqfn2
SR/3lAv5qNSYhCmJcZmRCCwbrOJfp9UG1ArWk88uEwkluAqgfNaBZ0GjrlbxfMRut43/s3oxF6mN
iqDjNBqBbkbSq8Z+jmvSQ18XnPzxDlpdEI3ACljqS++rUJGvMOPGrSszT3iwBQ4+bf3NvBI44D8l
JEDMkmzxfeuOtjUSITQX2j6VXr8QnLh9SIKBI6p6Jq4TKESYU5LkxuiHTiWqPsT+aXJAGVWLQ3PG
71HNbtyelX78n878ytnAbJIsKgCf7TQRWcoYGkz+Xs7SAJFviSnzypkPms2SObfrnAr4CFZzE1Tl
qaGBlwRBclyHd18ymT63G/yKR5Ht/n8dA3+FnMEWjBWimpz/WoOyMog4vG6J3PiRaaEOy7KjbbTF
edGAx4f7GV88UeTaIyy1zG8Pppk5V4pMXESvx6v10ZkFNI6PVHlkHbqJ0+8Z04wa3+FD430+GtPT
tS+6LS7qKW/ZNkuIZeifyaE3CPSs8+CfZtMoRhDDcw2BmJk830tSIfJX76CsD40hfZsXmhwQzMoK
+K6u89Jr2iUMKc4MfSH8/PgLHEbW7JdIGmYO9uRtyrPz3zObLF8/QpYzArYsuBXVJDVQPfRHr3lB
+PllB1dAn1kAJW/beicaEgVd/CjLfsRersptL4BzWe9OLQnmL8y+BKKi+2oAns8TI9Qbb5hok0V1
fDDZX1wApg1sUQnuRP4Z0GHQiDlLxjFaAgo5pG5IVxwdF464TpnkKa6qEzp0wNmcoxwoB3wZT3oT
H7o8+FfnWBY01s/rQzCVhWpjLtnjOKMKvx6n6x9avsA9UV8Cbbx/XuivK1XfcchvUx0mbDbAybg7
t27n5yVmCDKD7qtWuqfmTZiv3ovayh9vg1e0b7fDEYvOuMavJ+TyVXXLwiC7CbH1mSjjK8mweo80
d+u4sm2gFJ3/Govv4jMm1EShy0FWAIRaRCHbDC713jguTe5HZQ2sbIk9IYQFIEZQ2ETPv18q0ypd
5NIc1z1gDqrlqsGA/0cNKSuigJVkHD9Gb0kzbL7cLlYvwVWrf19rKMfZ08GHg9iO42yqdlebPmIl
PSEY2VHDdIVTN+mCilps014gGIkwJB1BiQtnDgPuz/dQC8nbOz+eMbT7umWSuzK/DlSD6UvwJ2Ds
uuk0tKtMiDCLoobpfz8uguuvqQ8b6xG80URrJQnvuDgAz3G3xjAdm2va7SMrD/QP/msTqL4T++xT
Ts3cy+zMFjE7II/x4IKlLRdm6VG8aokH+bD43momuAb9L195C1Gm1Xa+4rwcKShKTG7+TlMnP0/N
leOR8yAdiLf7lWOmOZvCTDQQfWAdwzA78pw1x40P2cYXAOjxvHt9VOXdReWffOk1WFmvorg1xQVY
xlOd9tnFfzKQK+6Z0H7vvibr175RshbNJNQ9fGliA6Hi/mxlQi4DDpeZG//pp7DsBxWdLOZc+mg2
t6YcT+PATQh5Kj4bLcHMSsadPdZpajIkrDjyp9RWQFmHLfhk1vZYv/+FJajssd8DLoByNc+V7gch
RQjqS/e75vWienJYdsVsZT0e+9DQA1jBUsu+RUpRXAeoorHHBxV89accYG8An6ALlMMGr/GobT4K
kqrNh2bZHJQLD9vtjBMYtBVnRSCGkMQz/ekSw9n66h55F0+gwfUcl/tbR/dYFM/oVk87DXjJMVWl
zOIJrasKClxopbTpJzbjz9q5ehe/tjuL1IMUR4JihyNXP9yTOUPHoilvhk4oRVLMJLZxu1k5Dqtj
N0CYf2BIt6+7mZQW3UTq/5Iwu9yPZgbXtCydXkQUFkJGhSuC96d5nVy9KtTXOtNnijlPVHgNP05L
Fm5H6CywtsggFPsbeNxxRmypIp9k8CrurolWbNJHhoC7tf34BkJkvKs60+rL6lKDYtuzdaJIN5VY
5Yo0aS04Tw7mRK5iRe4jbZqdYf2XfwWOYwyE0afI81gLOu0NUJKy32OZ8YqYTArPsNtzr7AIWGyJ
gL+sQtp07iTiSMxmxV4rZHzuPYRqlKmNfgVHEvauXKsAUfCw6zHLa+e6nigJ/EbSlUHv2GUoPAnI
Vi76amUMgCFvX4fiTCo9JN2bsavyGtmEj02PNPPUGuX84H8KbWfb/Z8i9mlcjwatHk//2hlms07x
TXNtBnHs2NoAMvw3P6wCKWqpgzZ0bO69h5VYwiG86bqHiKHQZWirqNC0Kv0z3+WW20wQUr/QsxQi
WtPjWv2uMiW3793TuIfKrJTGsQmQ4I9N1H3T3V8cSNFJvXhXoQdGLHy22ZpSHpCUwSV4j49RDsMG
1437jExQizUC53pBJMkDdCjTDKsvuC7S0qJgm2dhZPstzmm9RK4KEW9d62YoycxkLijA5QbdvuBL
eR/fE/E5rvSG8ANXbtRrzDdjM9Ni0lfOTVvhNs4e9ze+ABS6/5QfJQ6PTWOJnqCB7a4Hh+FnPmh+
B3THZK3PnrcpuDwPEN6oZHu8BjiQAnx7e5BMoung9xPtB+ZlYxB4wjGPVfIgXmAAlA0wAS1MGWLh
TQRUgwX/jrh3yZV3EcklLosrYlSFyidTarCaNIBRQ0czivgvtW0NqWl6Fs1hcMG54LuzM1jz9DNP
z1bHXXwGrYve9wG46d9YGQiKGRIzcWU1YHCxW5zc7Yuw4BnglPyrCvLgJ4i+nNQ5tvwqKuJ7dTWQ
reH8LuVEcpHq1dpsM1nAgtIHtBtrN3QYSn+98+6ggFcPKBzH75LY4giruds+T1278i71WEyecSxj
wlIIA8s/JKuAR8sNpKwpNoSdrYNj07XVu2htW07WIDbPjqB4DM++100db7i6xsJPo6mF7/HMhD4S
QE/bn2sUKJUsRlHrcj/61z/mowYXHsWybOyVSjMzmLupBlO5ocYvezo6Ks2djYl0/3ho4ytMSj4C
WXL+l3LCr83BD4RA8wB7tHTTsc3T1hK3tbeWJlBRcpDQzqUdRygb5b+edeS3sdvms/KQbm8yo9Fd
069h7QyYVLp7EepBJFyWA6ZBCvDx07zdDj0YLtraVTQEi6zGQL6713svsBQ/V0L/NZIOBDOB7EB1
Rt90xFFOr5ZFd7uambGtIzGWMaS51BMQYmDHqUNFVAztys/1Nx0MkVkM0HMoe97geBkddL8hgyrV
mrf9BK5kFvJFDHvqQSpsxabNEHMppCtky217hPHRVmN7wG9cD1tKhivUQg02pPMZGJ+lJ8hXYko/
jMNwwU7NYBnW+FiiZgh+8Z6fmsBkf7VlCnkKirNfvqLM89sC1BVMZiAGLY8xLR7tHXMxEDxjkQL4
ZZrVus5xAOpN+vR0BmS4y0mqrw8yvtixbQDkUO42wR9DWQhRAB3tmDgqBXLWW1twJLDkSxcAgdtV
bdH+IJsspODKcMSXuKfi+fQx3tcb1kn/pDT0nMx9pMBJHQRY2rlj3/dZP5NCQq6GdQS+z3cOogcW
87WiSdbNKAXA6VT2+z0+gJYhG/vGKO4oQUM1e2Iu8tWLT4WFLZGljsGFT/+BaBRFg5WyVLSyItqQ
cwj5zhW+pepkxdRp2I1qUrFp/w77vvJSj8uMjSGFM2hpI4PyG4Kl2C3k/9So1E0HevHlZTnu/XQL
/VZMpoZUZTPBQ4lZUxHL/t6/nnge97QGm/Bo1/qBYZweOX/Bs+w5SBqsmk4ZE9C3o/OEoh+EX/x+
wCwHoKaBO5gxSgoSIo+SU73aO4ZmxQ/b3ZRqLhDPLus1K8NnxGYoD73CcGSzhCywXtmDywEhGtix
/9ARwBSZCEG+IypRmN1/3KbzSHxnzGaC1HExWyFrEu9iEzFx72OoqUrfUb7hvh887/nGjXgiHFKW
NFEFFSPRM+RsapTkeofiy6tD46Czuh4ibfPFTofob485YlUpaxiXP5xCRXJgEMGTeUdLWIapbZXd
u+k0WDGc00XqYd02/j+6qVWUShsLo5nF5ypOzmMhCA7wdEQ74B94l/R+t4mOzCPgS9ewKOV41kLJ
CsGM9oNq9iu/z0M0XhFqNiMT4mCFH+2HcXl2I506i3AyD0Pep2z81chABt2J2LUSY79Ttms+ehGc
wx0ucp+PJm0M4UKrxBMT0jVzXpnGJYicD7rAA9ui3fC54LDE5KwejWtRCLw3wH7gD0s5uqG8dYWr
hDIeKGxsOMwZVNrHMSIYo9lx/fqwZXVBL2xs3fu9J2rAmbVq/q/mXzq6EWYMe89R7q/cWMmUYu2r
++NPjz92aNwzxJW8BfwUNmTnTpisdEMJMRtHPcYjacd9sReQ5VzmkiYR5f0BKqF1ylOlKQ6D/NBs
JAZVJ+O+jNv2kex8luT1rRFOHxcm8CTv1UcYVDC3+l9XkDSrjSp3yYTyTjbHqH2PWFm2YL2YUAfZ
VuacTTwm65YppGrzqf+uFfti6crGwiZjx9giVaIhmCTKlxu26TLdnV0Uqz+SAKqNmVFQn+dGhvbG
sMQLGlLirhXvbhjbE6BsVAp9JS6NXYxZH65mbLW7NnAD/mBq47ifRY0S3yxbQXMWv36NwJwHIjCS
wF80jpuAvVjw8g+Ebr4PAiS9JvnsM8ly6iLb9lJf75XPFm0a5fw4K1Un3sDXoCHlaLCZeoLBPHqv
2b2ElXrf0VSB2naOZK8Azg9pPNTolDDHYLgLQes2YSKzxy8TCC+XIz6OGXsXUcAmVWxrF7gXb2MV
pjGbwNlx/OaR5YY5uO/t69ERo7tclOFK6Rh1L4jzdUR1X7YQ7Kmb2bmEhgKyY7cyO2iX0dz8vaf5
+n6W/5kBmTNQVE9FOzc5SLYiJMsGmH1lms79P7EAh70Golj9ba7yQtTBh8h0IRikLeqLv10DGxGz
M+fUbZKiPtN9IQj6RYZW5vw4xLsX/zyhN8UEIAaCqaLAJWe4tOohIV5fXhwgM65QIyThNdpKnpGm
2HdIhXLqwvTQ65PvGSvi/uTTMHrtoQU8DY6YaaidHIB/kAbS+yflvPT3Y1impzdLLYA0F2+3RKqC
q2xoRUoi4ACy4L/Pn+B9fvuiGbNOXjJQCeU+DnOGavCv38Pw7dzjPeU6Amg6Eoghp7TKEwuJ7IXS
rraYzImFyMM/KjHBcmWiLvk+J8G8/fMUiV89z0ySsSQdb5uIK3vWlzrkePFzyaFpxipm1LrFoOax
BJcOTXBcTgjmxU2BwZIYrftw8EIg+kqmq33hVRo2VIuxollw5sZAbOv0QNjaUfEaMs+yKQ3eqYi5
PiVblBdBL7JyQA4FO20XqYYxfo6z1/I09sUcrd+51SrXgj2zpMg8QlZ6E2BZwHCLBYbUp5J4wvqQ
u/BY6iuZk4IDZwUq7DW7gShEWAmXgrBgy/ROTSBsu7dazai/xhhjmhRVthMnUXfKhIxvlWNerIOI
ZVUEjJUUni2XeS2w8HCvJZHt97qnorWypNa6nbpPxPANAc6rirvTKgPcEszRK4BJRa8gCv9c2HNT
WO6ZsBwjmC+W9fDxGGLTegEQ72ZeQZk4RBpFhC/0rKZwlPDt/+QOCLYKXaHe+qlUu3ulGIAClWDt
9G/HWjY8Xlrtxl1fzhOHzBDfljvhTAJ8EuMAe6E+KziyYYcSU/PJXeYj7azoHuzYtQPX28c2Zez2
eHpd+Xd7y8VSp+p1iAC22/dj81yTboXvCx87SZID7KTA49eQUuMy1Y1ajI+JgPiwqdzuxpd6MlB+
q8O8IHMS/+0UsUvqwMXbfp/Ux6RiAgoqG3h/Bsw5czZYMn9PfNJTxg/e+Vn++Qvp/0HDGg9GQNvg
99018aZrzijBQQ9bw3GKDqOkzfdt1dRUmfiOMwmKDZwzNFybuxFW4DdQdobO1H2IJZA7qMkwQSmo
jsYLG/umKE2+4jAxm/g7tErAOkT18LD1qAvWFZcVKt0XKyJAnkKzw9eddosPdc/Ir/yHoVIE6Dl3
SZi6L7jxJwcgu1GICADtqI7uHiwquyu222+jHLR1J32B6kElfq8v3SzELU6Be87ai12vqZKlD1ov
tM0xgHkNEiu2BcYH2Atw1dvWbMedvm/6wfMPjseioF6USU87MmSgaizT+5HgbikwB4HK2Aui5yr/
BO9b34yZv8iKBLw10cTRZHHFUtKlVExQk8xUZigDapI6r9FzAnRExwewoZmEgvq8Y/w63kUsE2Kz
7kHcbjUfxbyCHzEVJOvGlg6X5Vs/lyezJx+K9ZZW8i8iOSNBeZUsL1+dKrXujF+w0tALyhfXgAX6
w0oJuOJmVipQs1dO4X1P2sRuvs9QrdfJm3MYfBaw+o23ClR1McKWWNkaNINFQ4WEU9rro2/2PzJs
UffndSiXxtxfTwQTKA2hSH9I34gzzZ7kbnbfPd9VnfOAZWMDp2P0ehecAbku6g5+9SXYJHHOWZxq
aHmf/GHqy2dx5uZu0MxEHq/55RrHf6ZPj1vWBST9Si0v5e5040fkwek27lHfG21aHdA7Y4A7YcFb
huwg6M+tBWPBPjj2Q/O/6wgTL41xYqmwDxx7waCnP0KEiCRIRL9Jx3gm6lXpqRyZzBwnrOQrLBXS
6ySfppFQUyVdVcQG9y9zqJrl1c3iL72vmjiOSWAZjKnT5VWzYt4QUNhu0XSbsOxJYMgj4Ih+WiRi
KMFqsnpw3IaRDfZTox8DnzW9A7TOAk/I3ZEO5RXlFp+DbNhn7wuSODHfwk5Rh6WBoQa2O12PiYjU
enB4yLCRitr1IL2qPFdMedf2B+aZ8kW4F8PRlO+rUPkf/JIktzdn2pMy7w1lqY7nADKzL83ArcX2
l6WXEdx+K9+ugoVbzry7UT2nkr8Bo0r/uxqm/2UzGcZNQBVycY4RPJGH7Ft8xQz52Pq2UHuw0Ji0
5K250NyBTk6Eeq8HAtmPXEe89J1dsGh1kvmIX2a5lj5xnaW6Z/n52mQLW1RoiPYwWe9WfODnbmbi
DfYXbRgg7NwEM8bflZ6wBtoxi5ovxKVTLD5SL2TOqwy6BH4jMTPbTarMykxOeRHQlVgpqSw4QEmp
gczmbwcrxwOYEJdMqJGvEfVLm4J7ZfSaJRv03qusYbznbMD+mFKnkgIMWCQdhy/mVNwwNs2UF7mQ
SALtEPrDBr4+LDWGl1fnz9M9mXjgmRhr4VpwovH6sZOjlhjCdMPI/nSuYXGZ8l6+ddVVacTvPzFH
JE8zLkZ7Mv8Gden5IGmIDS6zvocGKJ51McKf+PbzCXnLGvpsWPmICTo/OCHVLTh35DtfapyAj8Wv
RrigQIDNJWFZED9EbfT14BJlNRa57F273gY5t1SlA3olBQbMOR52T5HDU4GDIfdZjfUSsMl3XMue
+D+RWPKEaUFnlbY4tX6cTvsyo9+tRHodSrXkEOBI+LuElEGmLJIhoIxFTg2c+SToY2ok2HzEY4vl
PK0y+bE6vz0fhcPkrvw1vSybUWFrtpSMh87PfBR/onR39vTkuvvD9x76N+ktPLvAurAV/z60+kFC
/4fQm2luwctSkM3uq5LgfOEPPclBwxNNgOFR3+PMW4zxI7s09KlhikHHFxyye+G+soKLMvNbOxOh
RBp0eIOvoccGXAYZNiEts6XtR824f4oUzu5tTaLUzanHD+uCEyNlZtd8DYIb5sQRPGyqQDoCs7bX
4TfAYODOS7HUQhvDLgfONqGEzrxPjkW9U2uG3CEWnP6tdEn31MzkktDquGpzIzSd+oKf+E/jOlQ9
mLjup5trGlhi/uUf1GRTexgqU830ebRAaE+2Q3uqyQMkhbgnO+uBN8bsKviXzfn/h/RRob38fbfn
nQa+0Sb6Y/JGcngAHW3mRBG1z+YkRpHUAfbGRSCZDwTmVa/xd72RyeXVUjsQ5B6UOXZid+o7Jjsx
8kcZzKuY9x74tMCFzb3NJKyy/QEJWI+BVHX+vQeTgbKlfsYtno5wIUHUL25+jTtKwA9+rOsOKlBA
Y7l3XaMIqPuDia8jXmzKUsTUc/rcdXWgucDYL/W4Hg6LAhglN7p+gS3P9DYR8BZgx08DiEQaPWqL
GC7IgQM1juwrM51TxzJkK2i3PqsqnxMjrhJm8kB2JGuDJgdRoAvDxnqAw+so0NrKzMlI2nY5/uI0
1sbAHrvQPVG0lZJ7KaDHFmL6yHZKjhCu43sTiBzrbzMkpvq1WPlW4pkCZSudeV/QXzk/no+TbGFR
bZyemOZWWlS+2kpSTOxx52uyeL2l54m5EKHBq/fErdXAG9AL4LerTmBT4miFhqy+t1qRCv2JAD0p
D6rfjU4OpSTKWLNyrD+cUtLRUPKkU6h2Qgfi2t0sQIVnLM9Mib5fCdW5ViaBLEg+xHzSjk/o+QCZ
xlBUzaR4RKfv4HRgk5zypDZ9ISC/vQ30n71Mi7lhnvIrBCw55Y5oGZRV7y6pISS0S5PxeieSIHgv
YHv1COnvQFW/KxdRthzVuKB0Wogi6fitsf9U2m3kQdHBhHwfIQb4orlzDtrb5VVgXObEZldyviUH
V5HWmJRG7JcPRpv0GRVzOMYYohDLcGX8s32Ju7kzNsRbL8I+rCCjcmftVB7ntoMB4bIs1v+Mtw5Y
NvVaL4kmbha+MJQ/vWWLqNGVpVasWMFkBuuX8Xa+oZaivmeT2cbPyX6ROw4dU4tRGj4RmMEHzqPa
nMZrAeNb/lDsZPepEhe6va/4p1mJcyJRJ/ETf9NRMYdgcAkJ9cwOzStzvglzZxYh+8lNaNX6KLS1
GQAh23rtY/DlgdVTtg12kvQXiIg2dVkND+7MKNImyQSSuVJjf8YCfoaM43mfNe2XlbHODQsUYstT
tGVJ0sCUkRVuldNZP8zZiZVrrvE2g4srn87RUsEiIlbm05CDKYNxg0WFjfvfzxpXUTl6LKDHQ8qp
hEFgCOyhegjG8t13UJwK+BkbpY8OKXDJ8BplY2OtaSb0X9hJ3lVs2GcVeQlhh0349K/wYKPPN42G
aLxm0+mRwDURV4QCd74tk1ESyfg1I/SG+SouLAXQdjMedEdBL+1EmXY+Miv7MR8j0d/8LxrsyXBS
fAM2aNWQlHWuFETXqQEvZVaf3N+6lH2qPKR6B5cbGcUp0EAe8RC72JOHjrpSXV77K4EXeMqv7y1Z
9j95lp2EWVwanbiCZZmgmSAhpDIgZ+lMvUO4cPyZaQm33Owhqm9hxwanW6VUZTcaoU9zdJOcQQBZ
/9U8zolaLj0UpN9xftX3wJFtQhM6y32DEgoKbkZLJD8MDwOKzhFMgm3D4yOgdjYGJo0YFTh2FqQX
Q3gSQqifRYsuxYqz7UCv4Wvyi2X2kBCAVM6unWQpcacsmDvE5XBOyaWrFvf86MpSN9UiPpvcVIsL
rgmCatqHsqFO3ILzcup8uJ6l+RwFmPtWxp59/JrO1n0MPAqP4qjiCsMgwZcGQRzicqAnZs+us9VH
LBWIwCLvD8s7olP8hPj4umeY2nU/3IMVuCCKOG2faHHpMLkWRIH1/CyRP5Fx4n0bctk4dSTU3Int
JkBi9VzqYpGtblf4C6nQlwMQIIjz77yItX0aojw6EZENzkBFi48XHXQiLyrsvG1SQoGnChsJ0IYG
KYgOWxNJaC87fVljsvaZbsIi0VnmBBXC0jXmpttKQFve6tdRCJu5VpfFiSC/XRwBnZsjSoFodH8j
pVPydP4JScj9VNkqVvh0VquIGw2sqqcuuq/9wVCpDe62ArYeqkf4r7sIIXkemZlBPKAX1WqRtMvx
kZzOGX1uv40KPDEP0dk8X287Y0CGSzSUO74dJciwaP8OXuuFCUiscHWGHdzGjCpCNK1LSgFIEfmm
dWEPibnLfwKUeOlGNcmhQIsjkmgLnD1uzhahDsHztQbd/XlsVSMh5XPd8Kba/+SxmwHztOEoP4h8
lB/xpqIV5vvYPmRCsdKde9zXnhgPCdbC/rOapGaiwkxRzSxsrJDPW6A07xeWSm8qschJU4oIm4VC
K6aKROud4RAqYtzf/xJZm1CX7Tvni2rbfKoqKRG4E/M+cN5yAPyqLGYWCiELISBp2WEG5ukPvp6Q
Fyp6X/a8D16kgLrV+0FgPVELYpulaz0VvqFymORyty7GObNb/v3gU0WwChJeB/0M2TTD6ohgx6xB
n9BBqish4Hx5/EqeahvMwdnmjFtOOHpyHvzThJz4jbq5qgbajrUCAiOi5Wpjex8qmOJyCks92uG4
le9KF7fTdBzgccUJ9xyN0a6369ce7kwxhjl7MuYOCBBCRNUSOgmn4chMjKHc9Jt7ReejNJLL/4j/
fCXnJ1/lWDpCdXtNlDB7j744ap+SVTsUx/cGvQeRzSFwNDnzr+x/f8vMQcr8TCXhKBnXIK1gMdpS
hRxknmLL89FUKSRX9ENerbh3RtVc+G2DTpgDLZW7nSa6uqEYoYs3jUcO+57gcsfbTBrknc4PIwDB
Ko7Fam57Ctq4R9CDOr5SxfCUKCp9ZCkS/AZVgNI9nuL1ZL2AUtA/RciWgD6SYUHmiI3PgiCl+h/M
GRw0S+g2KdYSsCVF27yDnG3zQrryq4npPSUUUREuYdJWfXqoc94TdtKgD6gzakJP73z7vIFr7r//
4W5Qv/QPz66y6lyMiZWwhmGBBzQYkb6wgzuvpE2IboMXnDcDUx2+ete9sM8MPyPL5OH8/0fGyLGV
Age/Bg0n4uECZ61QtGz2uvmw4c9+TbBMOMZkt3L1L+QiHBzulbNtqmv4Br0fuPhcrAoXrYVnj/Si
/nqRNnBMa1K9DSv1KkSth1WFdVc8awRI4k0UmBdOuZgKidMwc7iAZ6WxkjLbkw4zjhw5L2PgZIC0
tJ/KFDX1NbmfL4x8q5RsqGreoDJ/Jy5y1zfMPv2bfBkSeMEUcUOzCGn1xpJFKqm6xXudlr+YaVBc
+uLrW3cd8UTHZkqDspRFb75WHUSeHo3QfzzjWnnm/7VF6CnYLmK2NRGLcjkqkA0nYAMYk7lO2zPV
BIrYaJgyp2IjCXtzWwNHIUcDFBofnVPDFDVpVP53GbyWF8Rau5Tn3ly1GKzB8DN8nCWn/255a7Zf
53c6oFlMJ+SMKWY9u8B5qDejoHwgccUdsyQKzsCr621WLsZqeJHl9bS4q0T6A0YhnSx5cG/4/t6F
SgGu7nWhVEAYrbrqScRMxLHMMcPClbWcOhUejJ5olyrCTVZUI7P3FRn9NGfUaUxOMnrUV7UwwinJ
XDypIeznnwqEY4hiGOlFjqKNPvopvXWUvNOqD6dWoBIhHlORW2DYL1G5dWlgb8tnBlyJLZuZ3wH4
SmLrSAhVRnkgxXhjHVJ+0S/KT5zoVatxT7iG+K5tMOHStSdbtajNWh60Daufw3EsPMXnNIL4oYfx
nqbp+Hh4fOimkp9ZbQjk7FToxRDwTYHxzma3EYY4S90qWlPpMPmX1vvNvt8VavT/6aJXfPAUsUab
n39o4ajGhWMai5cYe8sAcoR173hkCcpGl6yU4X/IzT/eN/BD3RjPiYPTxd4nuTiuwjZB18dh4/Q7
6yChGn9dIwLc8qrychBRTHllUv5pHUj1qZhcrWMLFYO5Ot6og5wtRC7P32II/dMJrfS8OJaNumVr
QCRwTlrem2u76QhIO5gY7cwg4kPQHax+PJw4wvfcJJLo8xUZM6/tOeEGAx4KsFsDDXlV+6kpTtKX
5eOrgCefc8U3AkKMETGWYfpkQKfNv9fUiVPlmK0l3ZYfd/FLQBchQZiIKvTqLKM8YVZefs1G7aEX
bVbUp1r5x+S9dhzaonx4n6z0Edyg0V4Axmsp5zSH26enXifQR+sdE4oNwTMC8nxOA36pb0DWvbJ1
2+b80bgkoocwI/aOC0de2gIxIZ2B7FSf9Sx2UuRXr0gYUDa0S/moi3/VWYYrEVudvPN6vB/uHEgX
ZagTCplO3goqATPw+IPEhclshPgVWUYqTmupVjadx5yLtqL41B4z+xK7WaLDYBp7AO86K6mQcRuW
3K2F2KVQCMPU4ZsUAAHB4498jqLzHXTAwvgvEGXq06W0l6LQghKThpmNUBj/aLt6UURUwBZ2c/50
PjXS8/ftjPsAbpcB+Lfhqlwrf+lJng6yLA/tkNVXuOJRVQA3epUn8OJdL7l3Stg0r/RLRXII0NqA
dDV8/jHZEXLtKld333sj/ORIWvxIBNkK9DAqMhRDqsOD/Con4eqkBsHjbkSSWnhQGKMrw5XfUZ4H
Y1/IH/dtYFYt97cnWWm7tB7LxWf3vTp28CpS4MOqJjavGrxZLm5NDAUyGAVoJYGUHcHUlRDXrcIY
Cci2GqBS6Lyolw093vHaqPOflCfo1izb0IM2obvVGY9qrFaMERJqXQ21EYxutiQvYBwtz0xrQO15
BUe1GKnYB/uizoCVyI3E7dCKprLgs3wO8Lpgzm3dIF74g7xFUpkwl/d4ELusbjG4XwWK91sPzHIE
0TOgo1xJszsH54sFzFm6eqqv06HD/IZR1CgZI6/pJcyD5w5XS6YMvPazB4S7I0Qxn1hcDWIPay7o
FGkhXLmGm7djoTtLGAc3rWkOpyjKgm3t10eo2Eqb4E/0sS09S63sx7j8Dt3Ty2cIdsiJDXXUVCVh
/NNqKIlhKGmetVSV6iI+Cy07cRy/NyUs850dNaPPo6PI1gmMwjnMS3Y6sMya/ZYMXDNseLq/XH7i
MyWLWhyOHFSxNPJlSPK6ZH5Jz288hANNbiYNvABXSnA=
`protect end_protected
