`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4176)
`protect data_block
FF+5gqd0b4iwvpqy0wpQEassZUjwDIF8QuidTzWAGpEgFDWO36seShBig/327JYCDYOPn1gDXpb4
7bQQUxto9EYX9KaEivq0YsDbn3jLucAHKOC/bV1Z23n4lDZE7qgVxUIXqUtuHatYkrWB4wan3CmR
JsuV/Ff7ETUdI7W2zog+AT7RqGbwjfO06Ebu/F+nude6ZWbi/JV6enxjkmYJ3I+KBeKCHxvBgv4S
3PejFKkn3LLj8Sr+kp9ne7K32I2PpV483SHUtHHkPvRhA/c9/i7U9SJig463i/7ZaIfWkpc1CLwo
mSdradDy+Wh28UE4wvAFetqzraBnnpGI24YafjnbKWyg9Wh16s6vSVYUiny/kLCL/sicrS1KxbTn
AVrxwreewbDA2kJ8eiwErWJWdmx9cd7u3PHnUf+4CLmE/tYB3DBtrSrRogqOcI54cgfO3+iS6lxX
abY4/R0txlnkzQVWoD7d6/kh6KcQ9O8M0AYjH0Wq5YcspaU4JqkOb7q1KNq1rLX8DY7AXH/Lmtii
shywAyiMGZEpJkFVngyb7JomHWN4/ukcrngeDQ0TFLkhGjvwFuxSxQmPU/n/EQ3YFb3iucdo80No
a6vfEufRNp8QcxFIS5y2UcLeN5SFCZMdZaCEc2JUxQlYpkO/u0+t1c4/vA+sq5teI+erx4VW3YVw
cIQw+HjouxH4DUbxrJ4pNdnnF+GTWzVBokiiwpxsVYklTY09jw44Hv2cRL/HslXJwgEVnqFWQAGs
EM7jvIjJFAzM7dm/cgH5kpsUSq5gZEdg8+NZ8UyfJDeKfZYhPASGxvr29cxQbkAfDKjRxa1juFjG
3OqhvOecW5j+3g44lRXRVmYi5lcfhlPHEBViAka10ePRS7H14uoeBwcyrWGqExJ/oU3VgCX7CgEt
DDaNUrA3oKAVCBOE5hsK76XQIEuiuBvSbUrBsIsyQDkkhl/VgaAnb5MCtBlwcnCIVi6hh0cLlzXO
pYNtlgl/RQ3uLBkiL5cr6HIilw6EYvas7M1teSUYYYUTIiY3SI2MXWQBdA3a72saShL75DuMRwAE
3D35+PzcUQFuxV/WzznXj815OJzzFR+aejGac+5AKLhNozSQNZtL0hVrVMGt66ycn6LubHElpDkf
1oCb5FrK1+26uYrF+1PLFy/6zU23WDcBH8jCFdWLzOubx8jz+NwIcKOZGIEIt4odRummMle5/QVZ
8VZdj05SzsnNoltbZm1D8OkrEN0AY0NlcKSREHtUiRfjSoF8Vd5OtjHSTTxptiIYooyVgjuH0uwK
2XwroFzHb/51ni8X/FVFyV3u5wy3EOlfL7aFAWavA3/Kxm+8y67MkSn8aJt9y7YF3YzLVQ6jQpNQ
5/bhHVg3hxzV53JJXxG2ze7i7rjs9bq8a8YeQXxlNZ11fEZ5+HYVvdDJutHnsW9ls6wO5DHDMFDg
8MOp6CGPx0QbNWYQ6TLxs+KpZDpXL6OBHpEy44hkHg7excIi6z+W6tzj1b2HzMkDgYYmwadZjwWq
w9EyKFfTjtL99h0huvog6k5O02gWp+7LwOfcqY08poWOnkDpARUyYjg3fcIdP203NQHo2TVfG1aZ
/9+zC2lmcdlvGESuz936t2Zi0DPhiMfm3/M2O2jborySWLgwHiimyIVru+JqjMMbwRvyVU/KhgDc
X3hAojJiX70vqLrXv8H87t2/J4PvqJHngdGrDLZfL5ArvbxN9tU3ivCJCXhVgvToER5jNtXBjS62
3InPJDtJJSMcx3hZa1grE57UtEW/GgWG+FVHZHZpp9nU4bAm9FhZdkdCKv/h+cD43pSFr0BMk63a
dqrK11FM3xtuKupxDN1WmvyT+LgyQBdP3ar5IheY+Y7IbFYoi/AZC9mtZLfidiS7BA5fxFhlSMXM
6C6w7Kt8U1rSdbkGTDN8fhj/MMECoUEOVwAZVYNFXKgJ2JpJ2LqdRgt+SN2i38P4mDqAby2ceTy/
wDL1cJTCUeEGymE1nS5KQhUAzYKAmm2BJArF/cDVbzHYpsSpUOzL4DxMuL5TQpuSs7c4kLMRe0uM
ZHQMj0AUWRpYRfx37iu1NGSsROzZfY0fgz9CFMtgMEcfwhawCvbfL9/wSWyPLXhRVOyR6Z8+KrTW
+awgXkq8NUcLEqh1G8mNWxj8KDzOkAUfULLW43sS9UoNP8oivuAyNioy2uli0TNzPde0+EDdKgaz
O5KE7XR4cpo/vRcSiZ/oMxQC4Pm36xu12mXbhem5/RLHlTCrdEhKOKeXg7AZSzmsS81hnTLL+ebj
JnU/99yq9JVBKBeX3+1EJ0xaRaIioAzB1ZXobt1gdVTs002vqnH5cjdYSR+jsNtzyWXKkhNKUx72
Tcx6Jdh1qm350ks3aCm8hkDoVzzNiyDe4nZDiNxH/yfac0rySOWGjnWBP5VT/V6Ma2J7eRakZRpq
2lXOV4wnunFZnzZR/zBcWowCOYXtBHlaKvOdHFrZimDMf6D2jfrB4iuBmOVBdlSsSrn1/UrmP+mt
QmPYgmj8ZpfT8q0j4ibn2Jv/SRyKH13xINfqhF1dJfugtCCCLRohlBMvXWLntxjF61mpK5Kym9lm
V0MxYFnOGf+2a0Ud5U3NQ7A1Xx8GKkJ5Bc7fZwko674XHUE7Uh0xwhLYzQj9XSNdp/NvqcP3Xh5N
eI8SPBgGj+nDIwqtW5HyImoSHIgpI8DWpFdZQpgAwp5vK3fetElXuC2mOy2KmW3vm259PaEkkd4l
IM0vTvRwUbcwGqGVda4OcsHA6gkBTHnKZYLCdrgzKiEpcou/JEyXTUG189Vsqi4X8RjiqG5+DdXD
2jdhbsnUMt83yUB7jq3mOhE2CkvO5qTAJtTFphRL4mgj5EXuMP1Cyuhb6/TMZxkj+qpczrH6RqWe
SLLqPgRWbhjMqZXVqezdajkcSjmDNcBrS53DTIZ1JRuVWSQ/5KxOuuX0k4k8YgIh3kDJ5Tr2YhjE
17Hb0CFkOjFDKtthgIB7KYJPqw2QAVUMJ6cIgqtMzcxMoQD26SqK1A5q3vEN5BbREYqCN0qHhvEt
yLuFgBa/W+RL3YWEa+ouBC0L+Dpc31yeygDE0mFVIakI09VsF7BZnky6Ge4jey4VEpZhB5sCvL5t
T/XzuKjQWWuTNN5X/9rX66rWCgJ93TigCdfBAIIMgZp+T9VzUoVhiN2n0NHpaVYtzdEDIKH4puHu
v/zrprGmnog3hDcuvmwJsuCsKmS70EJZrBTfhnnS8MyRbpq5UgyIr8NwcqHSsPnRkTGsAHivvGu1
9K6wUOI3emDr6aapHWWjk1dgSqYcY2C0ZTxAg8bij6L15nk3cXKRJMgWL6+7eKaGjuIYBwwKPQVa
0iJNoflTITIc1TYlIdtnQH+mMZ0nyE2Uz8WPcoFfKhiovvkBJe1LoDfoLwvIvQsShEQnR1aPH+jM
fQN9wzOvOSmUNQGYLYw+JJRfojRHhRchLVRWWapmmy0vTKwXmIwry6xOGLWGEUoE17DnzcLI/+uP
Pa8cZhAVDIcwnQv8eDqRIK/YXdyUsW4TG5kDD+h5Mb6jpAExgoA5SkS172JoztVsjc+aKcwZxRlS
T6Zhg8TtsYACn2UjFC+RYohNBfHoRa7TYjc73S39rDGd903gyyF/FNwRg3JnbMEWckc8SObYAD1o
J8cGXcVaiKwlUg+D/aN5fbS+4Q6vlyinXcKGKqAoumCS+dAU6HznyqRaClMd4U7dT5PZBCy6OGTX
S7ZZ4/t7iGMVD9Oe7V3TbOj9DcGHgFgsA/xH01PxBUmKn5t7pevEscEtOEHanu8zCanHQq1OwZfX
CTtNJ1vjJo4P/YJs+qPQVbtctyPzoRFzBuL53dzGJ4P+YsgOgCuZELWytNsQWPmbr19YCmVZ9F2u
foC9P84P+w0xb7WMVIqNwmgCaWsz/GIiE6PlXRI3g1rVT4jlKGCTJG7IHLStgJGH36vpvpU0CGqS
EbQ/9n1NWZ9zjibRXbCAGmk0YTuOpSSCqUsA1EIAEOyAUt4RVWOcQZzcQAOKopzoh8eeqNAI62Bt
r1ZB+G0v7TH15f95C7vrM2A4n+ABgacyLTpoqNcMQwmcWF0ewRJo0jQW6vGb2l6Jl71ccNmEnJAk
CYr8Fb7wvsubJE48cTCGptlHfsqbVzxbSzFS+Aqgv5fEUBFLpNnEacqRR4bCNEAZbWlxFPZvJDqf
HWizv1HgpAsilDWcjykgf+V/NwmJmkJuc8+IfUqSIEw3zm3kmf+pWwGJfSvT/rFxacNhmhQAn2wf
tAuS//UPB0nV3uUt8rEl1hn7E8ltuDqwGMHhw6k3QVZ0ChqnUJgjoNqA1gzM9j7IFlGtBDJlFtZ5
PcsS3tveCGGYt0/PDijGcJUIPValWRwPFvbJ0zqfYW4mEj9+BkaHJx6wWdlr1wjNgdsFH0xoT4/U
hxrB0cyPXW5KNJQFN8KaWndJ9PZnXKN9vLs2OZ2l2XOyetqZS2sem4Cpzs8W/cURZ5VxezEzHTJL
LZ4gv6lQ/uqWz2gnQ5xGQm3TtJ+m9nFti3LzTFuIERRBLShQas7ckoaDJt5dUbHSBjhOz5E3UR8E
LTU8F2TvzWIHtUIwcAtocy03jkJ1+g0tQM0eAa5pObvEqS31YobUHlst/uJlPfPzZgEQML7k+A5d
azmxuiyNZnmhLbTJEqh50vm4AnbsPJFwrLKkl0UcljqPwhkiz5fQmgTtGJGhj3eInzbNW+f1wQnI
ngIXnpHi4wNMTpS7XLfgaB1XC2Cps74w1FIfFbWP30oAv89zCEYxO3UGkv+0lojfgVgq9FzhdqKI
cDeoz3UC3XyFGUcnr2Ee4byr3Qneh2vonASuHjAjbfaJ2pVwW6cCXSsSbkO2XNEefpsD4gk4ATIt
KbGkwdu7jmpfHmxoShmrRhuDaWppoJVM1OpVDEeJGxFIzEKN9zJWq0TVSSVbrw6BznZ59AYoAeSJ
sORuGDb5mjfxHhJyAq/96PRp69rKkqxZm2BbqQqiU5ipjztom7+FPj7DC8hp0WrHnz33U/qOdMuJ
rXGOydOJL0/3kShznYu79TGq4CQ7qDAryrSR7vvW50qVnWaJUXUSM1/JNMKLUx+CNjF+D1Mp3f0S
x+I2Q9dufbEs+cXr05SSf/vd9U9fyTDOOh7oGReaIC+kkD8AZ8ZBrFiIQ5nLGfkp9qU4sgOq+Yjw
gMVkEEIKXIBM1HDGvRazN0Nb2MgzUnT990rMqQ4vcuPIkgOUKrGHP39plsUJCuEu3+CllQdRE40H
w8fRAvJVTs+Jv6srS2u7YxH+UgM/c4xae6zDDmwVs590qIZHMdudlHj01vRaSJmobvmLCZrVM3QU
Tp/PzLeQSlf7W74nvSS2d0KdLe/gsnfuKfTWvvD+Zu1+Tjlo7GPu2OPl8nvCQTl3iX9SI3HeI+DX
JAKI35euAExXZslAPSuno33XKwU/uenqJIkPubGX+xTctKgUowtoIDwFnXOE0Ne9kkqpF+BFgawS
fO1cd4or8Br9Os5u/kVERu1pI6wnwf/zavvgvMOASVMiRbqB+iJ9ck1aC2ufvwsO8QhY1WpfTuwS
+fQu1tSc9ABYlPZg2YHy
`protect end_protected
