XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��2�u��,NID5�y�p���SlcpY���Z��`���@h�D�g��a��<�j#�[��>�""�*�H��*�򵙎h���Q:9�/��߀�i��Ι�K���H��X���S�e�DÉ�ro]�D.W��+'�N6q�ո�X�M����0�fb3�D����*r:9k���p/`A��\Kܠ}���Z�u�A��#7��9��y8���F��óW��o��ʩy���ϔwc|���V�U�D�& :�/[L\���ZVOP��f��Г�$�W����#���0��(��t]���ϐ7�-$��*7�u�&~��붅�[�Q�M�ò��\����K�(E'�C�B&k\�������2N���^
�����H�t
��}�3F�O���z�&�����+�&�p��O��ͤ�����j�e7��r��*zmT�RGc=[T��"V���3Q��H�X�KN<���j�"�Z���y���:�N�n��JJN�2�^�,�C,b�/��JJKؚ�i6�����'(��8���P�B�fEm�T#e�f���"k�o:H�4-�cr˫ʲ~�����߬�V�qQr���\G�� ^N.��jK���~9k��<�����9l���K�$X�b]��+J���~>oO��.��SJ�i߂&^16�H���O�=�=��h�IK��	�Ci���UJu���^�2~@kz���ȗ%c��R܄�
~Fݖ�}8�J����B�}�uq34�A���7Ɲ�(F���[o
i"XlxVHYEB     400     1e0��,�<�D�.��)w<�ѡ���?WJ5]-,:�@ �Ngk@�Ϩ��oh�UU��Y�w�<�M/���D�֮}6oiBv�J��w�r]#1d�6�qj邊��̶�N5�_���5 ���q6{*�B9���q�&<D�Ss%6�I��i�ů3.�z��u��]/�{(�����y���߿�
j2U���/ ��tg�z]���:��T&�2��p���c�,g����i��rw06Ⱦ��TݱW�J@MhO�Y�Y��F>���)<zM��l�I�Ţ׮t=�����a����xD ܞ�)T�T��T��.O�YPTU�Y�l�2���D��U]�n���f�)��YE���e��&��n9�4�����;�3@��	�|��ϲ����켾�%mS	̶+����n)�Jm�m����HWm[)\d��K���2�#ahMҞA=�$hFo��"�=��2�i`�����InXlxVHYEB     400     1f0�_+`9�}�
=�6�']�G���i6�#�r>7���N�����}�T�u��{xմ�;ܥ����d�x6`R�Y����cmR�ECI��+�]��u�+l��x�@�t�$��b��Q�~���S���:�����eW�yh�M�?X�H�e�Tۜ����xD�[u�
�y��1T���<�'�J�~�5���J�?y����i�i��%s�h�8#Li���)���!Ğ��Rmy�*Z�\ � ��!N3���rz�ـ���
d��K�5�7\Ǜ���_U�*E	6��X��h~��E��������D" %��(s��(U�z{���T1?��zl�g�x�D�aS�F�L;,h�C��-�@orC�"����VmJ��Sӻ�k��N�:H�5݁^U��W4жA���_�"��LRf����}�K ����Ul�h��S}�rp�,I]����� p�z���(M��B��v�Bz|�1��K�����oC��]XlxVHYEB     400     1c0Y����U��X�g�E�]4�'��v2c��.��[�[�|{��ǝ��D�^�;_\Un�+��KH�q�v��p��w}(��Y]^�A��{��Q+����H~�/αI��ڌ�B��V�	&�8�*@c�3�R1/+�_([)��r��A�[�Y��=8�7���m��Cر%�5H��CNNKw���	LY5��RVW�n�>�Q*g#s�O1������c=9%���'o��/3=�]_�i�;���[0Ӿ�VFVF����3�y�������u��>i��[/��Y�AL�I�zȢ��v�ҧ�	������G��f�}��~!*_��j�B�.���˷5�������)&+����$mꅳ��|�䍹q2���(�Lw��D	��`��Ӵ0Ԝ+����GOW.iK6��`: �qxm�s��ݓ��AzFn}E�����=_0�pr\XlxVHYEB     400     1d0�Hoyl�ϰI���4\^�w�=+#\���H�?����U�CJ�_-YƵ�:��C\d^�/oF7A�=m��_��"J�ro�S��Fe�J;�,���s� �Z/B�G#����\�PjwҶb�W㔞����C�5k�F�Z14%����V�S���#���MQYb	2�N$�6c�6 ����N��<�Z�������7z��-j�5f:����}�X�_Φ�x��2����A�;A���Mn((�|��͙Þ-�v�z ?��<K/K�P��Pֽ�JmV��>�|X��&5K[�r~���#1�	ܪ
�c���WZ(�Ǭ��E2W0?F�����~W���OUd�ޱqa���G	#��q�E�R�Qθ��K��D�kV�x� � ����+nYB���񱲱�!a> CT#EBW��a��G��g;�5Ah-�UZ_*��0�����{�� ~�XlxVHYEB     400     2009��e�6~�E+�ݕ������$�������㣉�y�{1QXZ����
��d���z�*VvT����j�jt�l���մ\���ܭ�`��n��b@�����a�r#��	T}�B=gD��8���%+�?�-L#�MW��HR����wa�V��3��������I�d��J`�%���!�Qݜ�	��c�e�i�����ҪJ��V���cL��)���LC��oI���Gτ�"��o;�z��v��uju��R�f���d"��	��)�S��ܖ0��o����7�Uc���O�����0��W�K��_]Ebx�R6Kv��S�{����9ZI���I����)co/ܮ��a���E�����#���n"�)������q���T��M�5�3��l!V6"�,��O?�@�Z4p��be�,������4`��=Ib�f��lWz��_�5��;|�p�4�9�`^��a)A=L%D�V]��pP����5N*��=o ��%��oXlxVHYEB     400     150�FQ=�h������p�@� �)u�y�=1�s��
�����~���7G�"�κ���>�!(����9:Ω���U����c�������O)�m|�x>%+�A����S����#�,��=yG*����+U���ϑX�_������ZM'f���8�R]6������|�݊�aFB�#���D2Rfa��h7X~�$h�h�����UG�?���A��c|%� �:I���Z4��Uo�?2��P_�	�y�u(x�I�3���u��a��y��S��u�ɝ��D�|�է:�EmY�i��e%��M:�@B�y�wu��_�����)�8�i׬9XlxVHYEB     400     170%�{�}a�աaE�xC��Wg,g�����_�D���h:P��{�`#_gY�0�58b������p$�\ �b�Oy�����k�4'$i�%��^���h+���J"���5b3/�W{��<.��-we�rƧ4%0�M�f�ڮv_�G^2I��>��p����j��>�PP8h00�S:�L
L��#�&���	�Ꙅu��[r3}l6�p����AM�]Lnd);������K����(�T�/me��f9 �W�Cw6c��!C�� ,��ϡ�8��CRb��U ���Qp<b����c#���|=���-�5����@��9�� �o=��4�+��{�(s���mx�d��{]>=I5�XlxVHYEB     400     1d0�����	Gm��~~��w+�f��[�=j	t{fsr�G����$��\�_�T�Z�����Q���Qi� ��n#�̶�ўF���Kf"s��T����e����,��J?��_<���Y��PmX�@�ݶ��V^���Q�A�����r�Mn>o�.�GQ	W��S���ؠoѕ5i��0���%4x�VBn�pRp��		�!z%CEc���w<U�Kׂ�{��7�A>���`���wV۩���x���dY�B��E*����Jy���I����L�;S�0ɰ��\�Hի�=4S~L����>��e<Wi��y�!h\h���P�}|��-NQ)`E6���U�&3V.�Ȃ��+��������^����,���ş9)xD+��f>gi�i�1��4I=>e���ީ�s�'�%׶@"N)1�IW�ۑ��и���X:�mw�!��7��^g-�a܅���`)�XlxVHYEB     400     190<��L����=���s���l�j/#��$�M����*��y��s�A.�����C�ЮQ:���s��h�%fV8o�ǔ�va��)����y%%����R  V��C�ubi
4�U��Q���WZ�F�z7��)��g�}Z�ۛ&>�[�͞2��{'ǹR/����F�c|�d�L_���8�xK��Dުb����r���4+��-�s�����뜏���M�3OG_����@����q�R���ʟg�˶m{�`d1qt�]��\J8mEI;1zo�m&{��*z�V��T�W�w<��ܞXQ�; >ì���|�s�pO&�k�0#zUb��U�O�����9b�-^�h��� f�b*�}ĳ4���UXr����:y]1���\,�@-fY�yM��t YXlxVHYEB     400     190�[�I��M~=x�u�(N5lr�>�p�m{ ok��b���Z�9�N�<�X&�m�72��H	�#��5�u%Hvg�f�C�Y����ľY�ם>��_=jʵ$�fƷR�J�_�S�c\����E\|�Y%FR��N�3p��A��vb���T�."�w"��6
tK/�/w8�)؉b��B��_�ˁ�e�x�S����Y�yaO����r�h��N Y�h�;���t�hPZ�����|����y^�j[}F#s�_hra�s�6g"�I���j�k��QUC)�\�!��"�]�b#u D�^�0���m�ʤ���*8q0��C>*?��苡�#����&>���j)A�$r�;_��݅�q�#"�$��[��C�v��Mu�:�D��];��G6(2���XlxVHYEB     400     150�`F�|RU��sO"�,�Y����U�˰�}ܝj���Rp�^��P���0ɮ�tXz�>����҉�4m�=,�lI�3_�ZL0�H�U�Am�Ն�����Z#��a�7�v|sə�yj��îW
X/��OXW����X���-�J����J�v-�7G��0+ꏹNo2&�؜��Ji3�M�^ ����D��O5#Y�ƈ����Ug�4|�Y��X�E�m���jG�\�M��/�cYQ��|��n�P0h�26�x|��/p����dEy퇴��ȕSWξeh�{y8M� ��S��(��9Dԡ���ՙ�^�;���Ϟ=�WFXlxVHYEB     400     150���+8Pm轺�?� �}��}��چ��ˎv��+�l����E�^�����w-��P����)7u]����X����9����W�	a�*�,���Sep�W}{��яa���i�M�F�+�4R��.m���}��߯���ٶe�\8�*���Ѷ��g���.y�E�/�y�ݿa����ȿn�0Y(��Ǿ�E۳p��C�rO��(�t�t	� ��U��R)�$a�@8�����  
{���0���
��pv(��k=�G�f��� q�jU�z��g���;C��I�T��_�Q��OY��.�F��{~Bw���`D]XlxVHYEB     400     1c0�q[ܛ[�}�`����pw!�q�:�6'�����Q��Dbo��mH���hsP2�I!
7��s�1p��D5�A���kg�;�#Z���Nu��ȩ�.x�H������}s3���g����1翙��@��-��PJ���!�ˣ�b/�z�~�R(@MI���Hs�Ŋ��bA�?RPy%VMm�<�D��ޗ�J��s����y�sc���m�Lϖ=f����^�z[b����M>i��r>Ì�࣫#�I�/��M At�ə�
�q�]�B]��T&���難��֊�o����oH?p"5��M�@�V7�����Hh�ߒi�?p�5JDӴ�d"n[�l��d�I��Q����A��V_���/��V��ہO���V�Ɠ$�:�0>�l����, ���VU�PF�`��.��1B_������P�US�`_��XlxVHYEB     400     1c0=(>Z��I3����C���9�P��7���y�!�秷�R�k��!YU�ii������֏���v�Ad�x�U�2A�{B==й�W�ӗmJ�J��.���Z�$=��љΞs)K1B�QS��3O�$h�a��}ȝ��
��Sz��Ӝ�����v�pB
I�8�Q��z�q|~��oKg�k�l���=�kn[l���3�2+��	�i���`�N�=ش$��Va�2C]�����pPn�b5v��E�� =���Ka1jC�uF���L��!DD¸>)|��w��R���MV҂��h%:x��x\���ᅦH���c�ZJ�Pj1t��)���gB��Z?����n��W<���� ���^��k���n��)-{�m����wF���؁�d��y�f���F��7�dˀ�ZZMX�W�US�����Bs>+�	h���iI�]ձ	[.Gn.b���XlxVHYEB     400     170��-$���*�}B� 3j��=�����	'av�a�0�(�2Z�X�g�=/E�i޾�F������JBQ����2���25�K��[�+����v9D�[BH)\t�}�I;�3��r�������i���PM�s�g�|�8����v��x����t����y���������%ܗ	yz:���dG�MM4�"a�r�ɧ�F�c'��
�� jA0������J�9D�����R@TX-�h?V
����i�q/���R6C�]2�t��������7
��P>��v�@^�v�<s���5����i=�C���oG]&(� �?���Yfy�l�8�ڇ���������K�|��M���I��_���O�:�;�5XlxVHYEB     400     200���*���<yB=�+�3`��Z%���k�u����ʈ�%����Y�	g4t0R�%(�)�	o���&�V|z7i��wɎ� mVC�_����ښ��X`��W�_�G��Nlm8Jv�+/��p�G2
p���V��Tgl�O����O���EQÊ��|I�2,�j�g��V�-��o���(����N�/����b�R/M7Ra����Enz����.C��aŖ>5���QuB�t>�~~���`�8Ŗ
�����Z�gYcǚjT�K�����D����p�i�a����z��o�S�����]uT�_|A:�͆�~���:kiB�e��hcA�>���]3z��d�Q$|�"-+��㜽�h_x(���~>B���7*�1�]۬�����6c릅9^�̏\>��=�ím]�z�\_\=l:U�4��)^?O\���5gv��f�sQ �G�l���އ�7X�c�7�{�u�ef��ȣM����e6$���/)h�FXlxVHYEB     400     210�`��Oހ������i��+Z2֜?!uFrۉ��U�&7��y�1�lM�:�}<Q�C���?�LD�dQ�%�~S/�ߘ�7�3<�/� ��p���%��a���C�BH���5	�Q�@��L��"Н�BH���lLG�(��kI�_�dc�e�D���Ss�q���'����p�� ���l{�WƌӮ�Y?`T 2�K�;
�!����龜"�(�eN�F�`�K:=?�U��n|�˔�,�����WVO�iM~g�*2�3�I���m]���uY޹��7�"�/�V������k�6\���ץp��*q��:qa	�ƭ���� e^�.&5�/<���,�Q9���zZ�<R|V��<Hv�0<<yk����RE��>Z�O%�b^��C�KY��*h�$Ia��Vlb��޲3�uw��by�Fd�_Fn���^�XC`�b��wXDQ>�p���C����;�$�r\�뾺�Q,�oܙZl�3!�sD?�K��׀:��� �r(��W����Cub���<$H��Nfc�XlxVHYEB     400     1c0f�Z�4��������w��o�_W�+(�A�y����%�}��4���)md�mZ�6�WB�@|$��-̍���z�Zw61�pmP��Pw{p�Y��
��Q��'7��tMB��.�x}��M�o��Ҥ�.�A�����W��:C��g��B%�F.6_�� �{����^q�[ {�BAcTD�D!��=��w��t�VJ�&-*o¯���o�µ��^%�0��$��]�}|��.����Г�[�Ԋ�u=���ߊ<Ě��^ʽA��:ẚ�[ݮw�OC�J��g+�VWe9_�ݺ\B6$�:Y��_��p�Ccʂ��P9be�W�PB.Ѹ�e�L��#���Ǣ�d�IE�!�Y/��h+���6y�)����8&+�Lt�H[$��0��E^%���w����,Pެ-��ub�����k;�ȐXlxVHYEB     400     160��:����j�|+?UmҥO��%��`H�
������*�/f��Y��g.(0J�\>W�(~�;+�w���hR8��0ô��k���� �	&�]�g�|�ֆ�A5,V�?�6�ߛt��p��@���̈�#�eo�̭���6j�F$R���!�; ��m46M�BЙOӊ�=qfd���B�c���H]_n���28,�	�s\I�G��,�����+��y�D��BD�C�aMok�0���D�H7�y�Q�a�6��G�p	f�k1�ͳ>77��JT]���*��d���J�uG7��4HY��vg*��Ѥ����Dɗ���O Q�ѮT����.j�k��5�����+tЇ�!XlxVHYEB     400     120���^��-����j�������.S���m;Գ��Ne7��ܰ���ke�U%Z�\!�_��~WJ�$oo~p�1��&��w�tJq㸔�끲�y�ֆ|K<i�7��,M�o	���9������)3u#�Y�����o��P�*��㌭d�F�VC9�1���)4j��ü0&>�b��V� +����%��B��
H��t�MَK�����Z,�_w|�~�e$WVݴ��,��ҠQCi��%���[�f<!�pĐ^��T(��+R�g6����%XlxVHYEB     400     160R�Q�o|﫛���i-�ZD�e�H��"f7�w!�gB�6���=�r�Kܹ�]��3Zb+�o�2ƃ��c��H�R������F={6�!�xE���i��mq���=5���HC�m��[��|M�;p��I��PՊ��-�X��p����N� rFrE����W�^|;��>���K�!�C�z��UA�M��Le���F�?�m|�6�g�L������>���7�X�EG��4�}�!����͞��b�Т&*dԂ,���<�l��8L�
5mG�?8��Y�7�b&�1�{�|��[-��#��B��t}x�,
}�Us�8䑿X��r�*.C�u	޻+��*Z�"�+��Z�XlxVHYEB     400     160��Q91e�*v��Z�ۭC�=}R�4J7|�`H��q[�/����w��nar|��-���d��|*��ɻ܋Mpf�>ۡ�y$�2�����f�e����x�#y�M��/`,]W��1�� ��bY[7�p�m0T�D)� I�ȾҞ�3��V��S�m9��5G`�=���寰��UM�}�U`�W֮��T��/��<�0l�%��D"�$�<9js�c%J���F^�w"V����_�3�D8rs}����|f"r��7 ��̷��h	v*U����:��ɩ���D��B��{|�^�ɱmA_���3�^�1x\��!��*�%'j_Z�2� =hkW,��%�0��'�ߙ�XlxVHYEB     400     200&��j ��R�qXvlj���'e��n�RD�	��g� ��R���E'֭+��__�3���>gUϯ��>C�~x�D�N�ܘ�m�Ko/��\o�_�^4�����4UR�.�F��&K�>��/�C��cO�"���-7=������w�MA�����2M�O��x��q�9�{9-��?��r?���4l���
*������\��.��9f��ݪ���^�ظ��BK���!�O�rf���&��S���ҟ�%e�FN�e����6u�xtXr�I�4��<Q~��_��V�������Z�.�e�a&l���^�u�<���[�֑E����do�ػ��Or�i>A�<��3_ʜ<|L��2�����ݾ1�؆G$�BDt�xה��~����˟`�_��"r',�1�FϩS����H�n��p�۝�%�� ��5h0׆��O�{�'�2`v�(�sD��X�hL�[�~کm��G73���h�|��ޜ����"�)���.c��XlxVHYEB     400     1d0���$
}�{�D��B�>n�����tl(�p�4��,���������������%�����5# {��'��� �8wY7��N���8��Z��Yy<p�G�ݷH��Y@P�@����ʨ���h���K���潑�d��g�}F��9�'@�"&����*\Xm>�ar�+[Ĕ����mX��� d���m1�N���h˂WOǴ
��?gT>����\u�j���=Īv[(�Ԣ޺��I�6N�ʸ�Cҙ�J�Y���To(��J'|���$��4����jN؍&��%�a��I�LB�6���-��Q��ف���}ߦK��5����dB����iDc����|�pX��]�?�ͺt��V��c���WS�G����u����Vl���8����	{CNN��1�P�0�rgT�D}߷�`�:;�DI�f����]�#���;J2�XlxVHYEB     400     1c0W'	��Q*<�8\��x^��>��	!8z!�#L��h�t�V�v������"� �17�75����x�}��W��@ӷ��Y�b/v�|<��ҳ�$z�h���.J�A�K��g7�.j��_�I��Ԅ��E��yuU8�ߛQ-�����7deǟBk�veA��%���`�X�7N�b8�5��`4� w���=ɕ�k&����
Y��v�/e,� �e'~Ss�R磂<K�R��щ1�������!�L�LE�\ZN:��D�,�����呗��!�DݒkU*e�; 0
�"B��������f�����[J�<З6�X�<�L����6�(��oiЃ�Vý������q�����!���TB,�����-��wm2)D�%��OЅ΄L���YV1����U���Ԏ+�</�k?���	�VL�IuZ��\	���B�͑�XlxVHYEB      42      50m:����F�r5����-�|&l�`�=M0���'R�f:����ה熥hG��w�W�|���P� yN@b��AA�