`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2368)
`protect data_block
2etu6N0x4D/A11nv0oWE56pXmc1koTGgwq1vGE2uP0Oqftgy7SEpHLxZtDXtOlNZ2yzHMdyxzQvh
hZJlK165HmlZwLythGUnvwPHkmVSW6a8OjxZX8A1ml/MKi9k2qxamW9vEdzA7potE4u8hrhyZ15y
UMkReQU0Ckxa9cJ0N7ywuZBDA8dUxYVCEZBDrUNYoBqdKWh+Fwojra28ncP4bnGqKl17Rriu/RmK
eLdHu3hzATc7IfgSbO4x9i0+pOdteTHY4b1SjHjXvV3iIhANGZ9Oo508FUInMkW5BDB11p1GjKmi
C7cXFBBJLFvXvBYWmUHC7l24UNSgJuyeKPo5v6yPwkYLX8QFgdSZ24euw2Zs5qigLPU5batvGKcs
Yj4BVyfUUeZEEWcWgj3qhQ5sTO/9TQPInbR0jR9+eHb8PG34JkuxVpFmCuCCL5KSvjL4mcNIIA41
pTUtYuJvv9PSKb5X8FcgQ7/4SVzPqoODl6VkubNvepZansdJJF7nldQj4rOrMeKt7FQUiOeEzEJE
swZuai9Ke+okv0wz0kHWL2MopsvLnFve4XR3ZIJNn+4j2Vhno1OIrwWkpoisuo0WVqsZcRY830ga
AgZfOoGN15G/MF5d4elMw+UxXUKXD4esXRy3VjeSHXFLTTOEqpGT5vHRwLcBhKVEZYrjQI8y3EJy
oOQ2S3oAZ6GnGs/yGLn5EoEX6upNJyjtA97lekagizb7IA4kmTGMumrtB2Vr1XwWDTetJsWTbNQC
z5l5NM1ocf5qJg71L6OnM/fe2tI1h13+fsxV+7aKlluMquA24BiOyUoWD5FXUBXWY3EGXYZlQCD5
ZSjH3VtgcALatwU8qFtX7sAE6p/YkxXZoc7JsoPKamg6tsLhosIc7HL3B+bJRwf06tjD8IUDiH8Y
PX7xIr5zCimd5wBEoufxpNk19UGXcrbxpCVaTnj9FKbit06kbmG84wPSuTMjZNu0fxAYRaQ7MUEB
IVjvVwd/odV+gAIXRLx/GsWTY6BdId+P4ZBz7kVOYq+lRKv1gEGHK9MtljNUxfpbQcTPd6srV0JV
6WrVK60FzCM4U8Poe0LOwR8eYNY4p129vTIaZiX2Y2lDJ/Ez3e8Ur5PltLAKHhXUDc0uIWQ+grzI
9zG8ACUDlDUHwwoit/mVaj4Ty/qDVAr3/2H7KAuuUAAef1PqtHtKU2aFImRXW8Mf826/4JbROGo0
dL+KqV/XLZRdngQql0S5+vnwFAJbIXyEpb8Nwog9f7tFGxP4F8ETZ+fzPS1/4oDZjt7dkeacNyRu
wUu14CsFYLZ+9QPwh0B6hr2LRMmhO7WQkkN8ut2iPaEolJcZnYHnUYRR/MY4L/OwDYsTj7cA7jd9
zMTY5mW/VvJC8HiJTLIKVcOF02lHUdJ3fZ7luxga5jWWYDEOPcOoCJQ0iQlkOYzJi/B5CYvG5U95
0bstigCypl0aNRJDYeN6yyeB2n4j5eT+0okMFfEWZs4lk1YTzktYmcF8w9dpNTZ/N1t4hQih/LNn
ouFcQU6RoYu1ciL4uiAQU1RBGSPSbooYAojCElx2zxYHym+sOGbmDF7DI51o0oxkoDyyWL5lPGCb
jnqc25bMNzGIwSUm9kQI4hj75toFwG7jkF46XRaxzGaq7r1y949ghpLbCuAfcXT/HiU2V4zb2l3K
IsWJSN5UOwXzOuje3wMSiLAwmmKQqg/KPDCRQwF+FX2GzHuC8aJbH2207WvBHmjIhwBeLuUs9YUF
YmQJZnQOXdyYQeGkN8semkJKqK1yW5PdzdMHw69N8oinMdVnGn2c/ycpmGBsZMTwsBEGWETHMulv
CgphW7yNYCFKsCd37WuYYdhD3tGF6HIhJYSXSoYf4TxR7J1AB/FuIaWXsfByEAHh8xQpLsMHmy4l
2OenIZYT1o03UNCzi3akdEWCykPpM2eWqz+nGw8ZsextbdyALgxo5mhNX6KkItV1GA68Zm/nd9ZU
Qs4X+PV5sDrD1TXIEEBifCXcByJaK/0TjkBxWgJdl4Flds1Yi6zBaq2GhtRjtSjs4HYd78YdrBX7
jP80oUEfHl5NqHYR6gV/gM2b3DO2rqogcnaPAPnuvuhpukllcnwC+BfWOJBU1wkXzxgI9ZAKxM3v
/yBlrBlGC6z06dGI/+EGiGKjvtaiguPcnvVF9pBoEAfPwIDlqudRKgLDsjh5QcD4fs8DmXoLChei
LhedHqoCWpWm6xJXIKv/x3+uQ1YxiHX5pC+Da1SC5wMe+hNxiO4SHyekRjSrTIo6SxmxSEAUoxZ8
/eKymxajeZVXRRKo4OxAlDyG0CLw7GT4j/IWMpvu4OQaytrjCF8PN80/IGF37dbrjDhYbB07RkBn
f94F95ijKzXHNmsrI87w1x3RO7qAcP18spP3llPLyMQf1z2ldw4zQnzhNclFtUE5q4bQq2u44wqA
zsjT45mLWHl66bgZ09JN6cr5qStNY9x3W3z/23tOq4qCq2RMcoHAESTi3zuRm2ude+6N0Z5pSGxr
VsOUcFxEe7EdZ1r6mATkZrFbCbCJrGBCq4d5u6unPE4AJpsWi8Y2VEqms+cbvzemhDZW0BwF8d/f
C783FgRL0tjOHXY64FLelEvG2vJWm4rHaxQKXenzpg4MPLINDiwG1Ve3QKD6ZuBKhBtEV+QQHrMB
cYg23f14QUgREC2jtHN0AqKgm6Hc6AGFfuJ74WOIIYyRotQxuRWQxNJ8fSnjXS9ibb/XowY4JdrL
ILHygY+vTk8WgGkC0gwGGzxHRbhTh4wUc6x86aR2/MlfOW/tvblcZQLRB/+xNqeH+gmIw3nxMI4P
+gnzgr5KFV5IC7puvqiHJ0a9BbGXJz+bN9Nr4FBzdefsYOLzAHuW7OY+tIla5lwrSwOdtRs0WwGM
7U/fx8NnCTyqs7SFojhQ1f+owcXzINSPXBbYZDB3uZc/YdFAkBmLSiLHoyCnWi4IsPMoLEQ3xtlS
tO0f5AKocVNGm1Jh+xx7F3zGPdp6dfM3FOLUxbtO/PBdFqWJO+ih1vfcSB3oa4vxvVxdXZ8SVwDV
sF2ER1NcjboSlnN9Z3QgbIFOFZ6UTYucqD+guzoE+svGtjya+gn3BYqYIRTdjTVwmEzCOHGTvrZv
0/YGt23mGD3mZ7oM3939B21IgUOcNJfWbJ7SGKsU9g==
`protect end_protected
