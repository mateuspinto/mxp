XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���2�v�3�Pֿ��������ϻ���ۓ�Yj] ��E��m�@�d��m3)��|��#b�h�]������r?��±`�G�`�r(�,9n����8�1�MTC���P���<tТRl�RYo�UL�L|�E*M�ӋƖǾba�qe�&�|Z6��ln�Mv��$H=}�~F��n��Vg������d�=7a#h�)��4��.�j�ve����3و���И���ߥ8�v��z������$��0�iA?t�N�IX
(ؼ9��{ȻOY{�yb3�Ա���#�[^E�Eh��؀9��4��ź�ω\�S�	x2W.^uf����5�8A�Mf�ĪOU�2�)��Oϊ�i��r��c�Z�ЀQFJ���6K
	����ɂܲ>_X��J1�1�5g�|TH�ĸd�\`NJ���G�#~n�R�v4���w�y[1� ���h�H��G��0;��Kݠ��~G���!: ���^O d�9�7k�6J��r�\m�M��������q/���O������v��sc�+�W��=�̎En>�ݯ|T@5�����<8�x�3!=�2�RY�h��Iz�@�D�$zr�#�O�H귲�<O!?��q��_L+����>�4���8�������O�J�S6k%X/�t�s���J2���^P��o:k��a��s�ڛ-li,h�05K����>�L�7��I�`H���F���-E��͵ �K#UF�:ǘ���~���b��R�T��"XlxVHYEB     400     1d0zC��c-�Kްť�ȓ�!-�I��A:���5�w�*�(2ȇ;��9��3�&h J�3gw��lepa?qB�R���`C�O`2�F���D��w�-*Yb��R�O��ڃ�ZQ���^�-2�!70�;�S�FuZk����[��#z꾦37���c"��z�R Ŕ�".��K�� '4��w�Z[�_��
��|a	�j{�^�y�����U�3jL�]7oz5����[�aɸr�[N�N����=�>����Ea������MQ�tܡ�W	���N�4a�ZA��3P����o2�J����5�R�3�E	f� ���>
��9��=R���	AkZ��p�L����|�S'֥���.*�ܰn(�ae�.���9�!`?y�l��2�SB���h(Q�.�i0㓹�av;�
@K����vb
^u�&�7y���l���v/s''t�f�����.Jʆ XlxVHYEB     400     140��?��?�_���)@�n����[wnDs�5>86��R�d���Ȏ��6����z�52�ZoJ�-�I��[���U��Z��h.�3���lV��Sc@/�c��[|�0���x��Y�y4�e�h�����7��StJ��ɘު�4�)�	��H�a�K��D���S�Đ�G���$�ɠߐ��x����$p��!7�I8&]��&��9K�~:��	L�d�:�A-�b ��B��,G�*�:�#���`�h��\�\��6�i	-�i^�EI&Y��_�����K(���ag�u�l.����Mgw�<��3ؙo�XlxVHYEB     400     170�y��r�QEkec�,c`��{V��U����q��jڪ�N�s]�R_!l}R�NO�;�ա��i�F��t��#�*�ֳ�5�r�dx���ٟ�9��:ѕ�eh0Qx.����^�G���Ĳ�%`����m���H�~��`���2d/��rɼ��\B�$����Dz���|Y��m�I"=&���6�l�V�kjQ(b5�Yn'�ݧ.$�w��7l���iI�z�$��Ͻ��d����=�7�5q�5&ݶ.�.��49|�r�H� �ۊѶ�["\w?H�v;�@J��N\�}"�S{؀��eLp�$�rHt�l��ѺS��4���-���9��Vm��Ѥ����L[�$  �I�XlxVHYEB     400     140��o��p�VU"������%Yu��ѨWu)m������A� �F�����ݠt�c�ji$�0H�_�x�$q���rП񭬝g�@ׄ�o����f�G��λe�cEu�P��~v��3v� �g���: �q./����?�s}��lu��Fy��ƥl)Ltӧ�Q�Ͽ�
�9�J�b����X�g�����ir�,&���~���ϧg4{܆[�M  �ϙ<v����&�0KSR�P�Gԛ��f�"t�4P�߄��$�?H��o��]j��Z�^�[DKV�l��?��Ƽ|�q�nMPխ��L���=7���XlxVHYEB     400     110���5d�,p{�uZ�@��5��WK}]��kVz�h
F��E��M�����8�2�>٨�Tk�9b]�]bٙK�y_W�=
v�$�G�d�p��h���ޗ�$��3�~���l)��p����/�:Ik�PW{H����!(�Ѿ_�YH��:D{V���s���"*2�wQ@8"�/�ެ����~�z˫�����e���Td'�c`=>�W�]y7!�aج%��q�lP��M����9J4C�K^﷚��4�{u^XC�A�;��.8%XlxVHYEB     400     120�����ӝ4d�\�]yj�3D�ɫ�D�a�r�lgB�ܑ]a�Xt�2уy�2DF��J� �},�"1`��5�F���q-i��'�A�B4Gz�$�*8�&\�K
'�����$�k;t�QV�&_*m��6�]�.��}I�5�ý>�Y��g �ߧ��ͻ43�D:�v�IZ�鼾�Jf�S�@�!-�;�ؽ�k��7�>��\�d�9$����s��/T���(��t	n�+�"@[��T)�VL�N/p��ł�qiP�`}C��G��)�N�+8wdX%�>XlxVHYEB     400     140~J�����	X�zo��[�) �R�2���k��noV*��T�D3����߿T��)Bw��N8e����*E-�g&����M9 �(X�"�O��o��=�J�[�2k�G#A|7'�|�:`���H��Kj���JW&c�AD1�,Oƍ.���7�������m*�yZ�PL��@$�<%��ܛnsJe<+�y�Ve��!�+^��Ӛ�)��&��gѻ�{vA��p���Az
����{�Ǵ��I޸����c�f ��Bs�xEl��N͑�.x��b/Ǳ��,����b��-}��6߆�i�П)��E��?XlxVHYEB     400     150��� �$a��3mQ�C��:uЕ�o��f�	�ԙ��S���]Xި������P]�S`ěr��:D����E����LOıD�Oѭ��3~ۜbHu�g�tB�Ȏvrj�_����a�ρ h>�۹d�����p��ժP�[��-FF�e��J���Z�(�Vef����C���X���8i6C����<o67�����6:ȳP�e��K���g`����]e?"�3��O����p�c�����7�;�}�S�ڔ%�Hj�J�ң���l���x2x��]Mr�G+�#�Q�M5m���}��I��"�]�k��\��I�D�k�Hԗ2ׁ����~�XlxVHYEB     400     140;�$]�p���T����M�����)2��Q��� �$��6��\��ֹ%u¨���+4�H���0��}Ȝ�j�q`�+�pl]M����l[��x~�� {E�f�������>��ǧ�n;u�S���F:�'-jZL7Q2O���gY�!y嫼o4z�($F� X%yE�|�븷��;o��v�]*C�F�=�	�� $�i�Pݔ��B�=`#(@�,>^t���yWX�%C��C�[�oo���q�,5|�:���/ok��I?|L2�z�-#)�=��Βu�T ���޻�[A81Q �2��d$��N+vXlxVHYEB     400     100k��Pd��V�I/L��*�'��A^H�D������$�s�Ю��$�v�s5�� �ut�u�?�Sh5�aI|���NM�u��/=١C{��i�O8�"<��#>�cn5�����RwzlW���Z��-h�I"�ب�:V�������Ω�x��w����d���-D�?ş�:ϙ��O���N��_�~�3h�F�����}�+y�����P	�/����M<G�����M�}��b�'����|@��R�-G!�T9�XlxVHYEB     400      e0n�����I�ќ oq0D�b�$@�Cy0�`�����ǐ[Хu$JH���{}U5o*Hʩ!4��g�k���v_�+m</]���=�k�n����B�f�j�JE���&�����`�b������J�[�'�j����W�gL��w=�WH��@�la^XI�	��
J/���S_;�����(��Sޡ���?)��V����k� ud�5
>w�&Y7@35XlxVHYEB     400      e0+��ۺǃ�X���]Ԓ��gS۩��^�y��j)�G�
�2iD���/Y�wg0^��(�G@��d�${�`�@/�k��Wg��#1I����Օ��e_,��4��<j�i:Q��H�xo���G#��G�ܡŝ(�K���3W���Ը����D���&�#�_��-��`)�p
��S���k���Έ�B�G�F��
E��.n��}���#Q��9c�v�&
]�XlxVHYEB     400      e0ʶ�*ی���4��Ҵ�k��;R��H�ތ���ZNy��àB
���^���_0�P�%	�:��o��F/aC�TP���c���P���\�ߡ����i��*"&ޘ#����ߠ��E�7����_X$��i��#��15�طs
�>5�8��n1����+���&v��=��r�A��A��`�T�����ѐ1�h:���*��UE��#�"ʸ�7P>�&�:�CXlxVHYEB     400      e0�>c�h|6���� ,"SKmQ���4~�줄�g�	� 7 �]�Oh ]�S,�	�>�nPv�#P��ˣ=|���Ʃ��q�p;]+�ͼ�
F&4L���@Y���Ƞ��W�v����.��r�E$?��Kx��oS��t��*�Z"�Lԇ3q������e>16;���؈n��L� ��� s�JgcXsܱ������$�S��1VpJ/c��EXlxVHYEB     400      e0¥k�O���+
>(�����8? G*���0�UWE���;q��*B\�i|�Jv>�=S��T�B+^g�*���4��؈��{-���F��a�m���CL3_�׻����������ɿN�n�Z����7�b��D߽Y�eZH�z&�����Q�?6 �m��K��;�3�����Cd���U1�R�Q��h���Sh�DT�{�-�3��Z���y�.���0��YXlxVHYEB     400      e0cl�=�5�{�D�/a��ʕ��ۙdL��MIV�A��	��b�� h�D8eX~ݬ%���qj��������.�i�L(��U}���+����j�tm�r����%\�s��TPo�`��`Drݛ��U�
kj�״5���bs>�0� ����@4�G�\�S�(� b���?kdG�֭,�[*M�7�'bO�ƼEBI(�=��#|k�P�م�=&�<�1�kCXlxVHYEB     400     1c0�oɾSz���	{�0����WC��>�m�[�`��v��]a�WK.���gZ]ݑV�E�"0֋s�bDFؚ�m��*�ܜ��_�7qRÎ��fW�l-��|w�ޘ�,��y�M�{4Inb�4��B��~�#ʑ�r��v)<��<�'t�<�����mK",ƨF?�\���e���L�z�Yd�j�]�L����!~9UM	o����4��?�]�|'gĥ!-̈�"���H:��8�b.i/#���zš}1�[����r0�m���ij�fS3ږʚ(�XF^��� �@�ͥdG,���0�Kqh������yP��#�g��Cz�tC�6,���}0͍��o0������A7�n�����lmR�{�y�pg	vp���E5�U,5׆�0Ԯ��e$�Z�Ů4�����vֈ���Hy��M��Is��}� �W��XlxVHYEB     400     130�*��Ȇ����Ԓ嬽���
�r}@�Gܙ�z�W~�!��b�:���Wc s�C�u&9��@�֑V<}!\�$7A��(mg`|�9�2^SS�T_�������v�?a�����*���#����M�~db+©A!a��
E��1���7��-��ܐ	 �Q%��z��%3�k��!W�ֵ��A��W��[qFꙟ��eX�R��?��_]�Z��h��Ī'��J��K8����n<����Li �&g<>���d���"�jC�=�*�Zk�͇�e:�u�U+Ʃ��=XlxVHYEB     400     100{�Gk�Y���g�5�{ %;�*�&��k��j55x�b�[k�O�=
�}�2��X������v��hty����@|��m"Y䐹L�c5C+:�/�� ���n��xPw,�z*����:.�z��(�tF�W�H0w���_dV���ҋ�	�>LJp�P���wy��#�(*�vK�Ih�#�6�/X���:�}��]7�+B�e��+D8bڱ��2��y���3h�[�� �,1ő���ZA�1��ٟ�XlxVHYEB     400      f0:x��A;5�7%9�V�0�LdKq�9=���k�m7'��7Fwm|Y3{����l@�1�)�9��%�\��YR��-Xj3�ڽ}H�G,>�0Mw��	�_�=ߢf�k�ia�$��w�eC^$Z*�"h�N��������Bɻ</O�ܰ�I��-���ѪE��,?H0M���k���zq��O�>��I^��C���[�a��3~޾6�ŝ��xfw��v�����i`�+�wynA��XlxVHYEB     400     140p��.ݮ�}��Ӫ���X����p'g�>/CS���,��p6��aцBw>sL�A�Ѹ�C?W=�	F����V7ƞ"��""��v���n󖀖���&����H�G޲��`�5t��	O��Aھ;��4[���)'"��?�^�=�.����w؛�ŷz�n�6���+�7]�4�}$2�fT�n�E스���R� +Ы�����-໥�R��)�	�WZ|a���o>T�&S�k]��5�8?wz��%�l�

Lrҷ2�^K
���y��̷w����" O��R��<��;�K���B�E�Y���6�+�J��XlxVHYEB     400     150�ۋ�R��`�h���`\~~��	�_�V������Z���i�nL'ɪ��'[ޕ�d4W���]��h��M�3;�Ќ����1�=��uɣ�
���=���u�������
��E�\'���謾�{���)��ՊEv�-�Q�gG��~��(��a����i�P���[2��R�_{����:��)��8>ݙ�Q���kX���#��Ƭ@|���~�]�|���@3��(�U�7����'r�jCUg=��$��>q���P=�+v�.���"QL0���'����b�?�	^"��Ų? ܃�>�������Ӌ�Ck%�\�}B:6�%	�_kv��]XlxVHYEB     400     170S�)?E��4T'vH^�~L)�J�sڋ[�A.�`L���Ϊ�� ��Gl�����m���q�&�9A��|Ʉa�L\�gOש���R7�;s?�u��v?�xB�,�/t�7��u����qMM�@�C�?�ٴ����8�ޙ~`�݆J9�5�!��WHY��9y��
��G�Ԭ1�f�˧<>�p�y^�G�2�����<�*Y��Y�Gw�#�5n�����a��{� ���iŀ�p�̹Ջ�I��.]R8ro��=��&r�ɊϷT��+�ǫk�}�[�m����+���c��]�#-�E���^ٞ�G~ŒB�.��k,��և+�����A�	}�ӻ��5n�jTOr���D�-�XlxVHYEB     400     16008��0�������%��&��@�,k٩�Ӄ��ϳ{_����Ƣ�����������u���2�]�\m x�5���om%A�M�<���>�ӡ����[@a�����7����Bd����Ű�_�G��#���Vu�e���M��j�,I:I�w����w����c4���k�<�����R-J�Q�O����לߪh݈e���Xh�x�F�|���o��Z� ֦'���?:�z%�l��"�2��b�ge	�0�@j��-�+�$���t��0a���r��A���	�F���X�J��4���ASѶѾ�5g��i�F.��R�UbK�Q4�XlxVHYEB     400     180�S�ٰ���Q�y�����Y.�u�Z)sgh*���6�<�"Wl��V9��y_�!@�U����ϩ#���$��a(c�S9����M���~����ETZH�����z��c?Z��a���;�nI�/mMf^���	�o�\V�S`��LV�y�Q�0�BA��ZA�f�	ӚI�E0S%�Ca�w
�>|�{�x�7a�Gћ-U�Yy����s_)��i��0ꊈ�� 7����?��$�-
�
g�5ܟ�	/��ԉ��t�H����?�,Fνͩ~�U��i�>�T�ڪ��%<md��P�/Ƣ���kӀ�	@���L�b1|�5�����Ǥ<Fi��'�V��N��E��{�2lJ�0�n;6=u�쪜;�f�x8��XlxVHYEB     400     100�\:�{1u�:�ܘ#U�<����d�Tgd��#jZ9�*�^\D4$�1W��f�*3?���s.?x���>x�vu�sK~���l���������!BDD��SL������k���f*��A�w�n/����������XF�y���U�j�n�GXV�A��'�>n�q�jq�k&�P'x�f��h�آ[LQG;���܃Zav��밽W?��e����U!k���lhg�Y�+���M�4��U�s4�臠�J��E{XlxVHYEB     400     160���ٻ����>p���>DNEi6L{w�?�(�b_�=�3]��5T���AIoË���F5�HI0@{0Ht�Q�Hh��a���]-�,���xT���,}I�}E'fOOM`�)�b�u��JV��3���9�?F����O�>F<��_-�	#F�/|5�|��d5��b�aPX�q<{z�\"��z,��!~�x�/L:m��#��G�:�-9�=�E�^��f�|��F�x�,�K���!���pN���(B�Q�K8A��@аT��b���
��W]��O�J.2�q^n��O�BCV���$?�}X���4^ߴ*��Rn��M:���:�Q��<SP�B�&�&���XlxVHYEB     400     160#�՞�:F�6l�-�i����}�l��X_3��NB��sk#�E�PG�~�jq
�l]F<B����g�s8����d�s����RD����p� Ņ�����ж!o�	,l����CD��	1�7���~���܀�6X�IvÑ$�tĽD%��a�{c*�7==r���1�(m����@ҹ& ����~�:m����wcy-f� Y�=d2R��y�&�KS�@���oek�;¡G�Zn�>�1����\�i�H�nb_�K@���NR��sc�C4���	H�ThX-~������Tɔ�y2�1,Q��Q�h�����V�/�T�r^�����)k�p�3L|���k��d�Ty��]��XlxVHYEB     400     140E��� Z������	4n�Qi����6̟��8 ;��o�9��+�G�o�9й=��u3wQ��:��IFL�|���(4��w��gAў�����W�H�hg��E���-S奜�����P[�[�E.ߩE�/��g�;�u�gjXJdt�S�jZ:��'.�vy��W�!��
�I��e��r�_�������Ȏ��X�,畤3�X�О�v�B�p$�)�.��)�x[�A��?��svܕ�r$߇�?�.l�d�3��R΁|���c6�����&l�x�~�˛ή��.1�
Y�8�u����s�KI[�%���}mXlxVHYEB     400     180�͎`0���S�q�M��0����VzD�ʠ��b�a��+=ƛ��;���e��Y.j`��˫�2{�jo'z.�8��~,�̚s�r�3�ђ	M����7�������P�� @��i�Dp	��lw���}�-��i�6�s�N��a'9��\��^¤��t�J'�q'�����+բ�M07�z��yt��E�G�D��ǅ������A��?N}CN�/�"��������;�$�4N/L`��t}-��+��/���}�3'�m�oW���H��dZl/���]����C5�ʾ�2&q�����v(].����������c"6H�QR�.FB�9����DjW��`�2�s�;4*��k'y;A��1=���XlxVHYEB     400     140�l{�N�PF��}9b����ЃͿ[o6ۥ�����*q��_��k��s'�x�g��Z7?I�E��ܙ�v2���9�G���X�y���(�ٓ���Ę:��e��u��q�>W�*悰I�ʧᬹ�|8�.��`F�Q�"���h�����R�Cf�Ԓ�WJ�(��k���V|�Re���`��D`�K�!�-sþ��� T�N,�^�`Gf�������"L�φ�x�I�pi��s��"�	����NoV�r��9�ܐ���t�;ԏ�t�o��Ys��X���2�>/y��i�=0�Q��K�%#�XlxVHYEB     400     140��ࡦy�m� Ed,��&h́�?W��c���,�c0@��l�����~��5��_U�P������	F����2@��=����t�Nn��g�N$����ai��7�Gǎ�;_.�˞R�v���sTF�*�T2�m�EQߎlx.j�la�z��D#V��.�	�B@�	��@>���RZET~�"�
"q-_�=z�������I�ts+��t{[��ԋ�J��W\���1T�I��f��5�\� A���`'���	O�7���z]�O&C����h�����o�b6�������u�\�lI(�Ɨ�.�|M�W^XlxVHYEB     400     130:��O�G�+�}�H�5���u���L`����=�gf��F�c�Ĩ��| �Ƹ0P��ZQѩ���;���9ŷ�m��K�͇��r����u|��h�u�.F�]k�	�g_�.O���J�D�Lv��$���D� ��՛�8��- ib�C��Z�\�>"����M�U\��&��l �6X��1(C��u�?�� �g��[*��nӸ{�:4L�b*����iQ���^Z��Y���E�*�ǴФ��u�T��QW�����Nk��W�:V���ϘI]��juj'H�i?�^b&R2XlxVHYEB     400     170���'q�¦3�S�����ɺir�*���Q.d޾'9�ƽ��T�����HL�����kqWvP]�i2բԬ�JNȬ�eX��1���[�S@Ņn���<8yK����|�Q����8J�t������Ƶ�"G�ſ[R 
/u�΢����Mi�h��.^׋�!i���K,59æc�u�	���OD�(�(����o���=�7ͼeˈ�"� �/�F���&�
�2��B,�^V�� ��3>�g������E3���
��s4���䄰wj1.��:%P�|��	�Ŭ������˺�}:�0�Q*h�6���&������e":��}�sfh�Ѣв�B3�\i�|�V@�rXlxVHYEB     400     1703[=N�h؜�7<�W*$�}g��!z�f@bW䜜��<�V���ܧo�c]�=.(�C�^�H˵��M1"���y�ZB�B]kK
d7R�(����?�AN��U� at�g�B�Oh�n�b�h�8sz����f�p9'貌TP`�c����zr�Ő�����0l�:D�!8��w���^�H��MA�Ze~w�xjL'�2�7�p`��~�Y��ꃐ�ߎ�R�-L�SO��ga����~�,`+ќ;�P�K��O?JO*�>VNu�eA��h/8h�׈.xa�HP��ʈd����"k�!|K��"�ۦ��:�34��U	���L��E ��dvLΞ�ˠ���&����!�)9l�&�`��XlxVHYEB     400     190n*^�	��ۄ��SzNܪ���B<&�.�<62��6e̤X
��O��8?���'	��ӿ_ö�͵�so ��`�:��Tr[N��=x
�Uԡ�i\AK���J����NC��H��V� Q�n�n-�Kzs���@s��=���l���WN[ӛ�崾�5-�L-e{�z���FCF�ƴ>��e��]���6jC��K] d��e,�����ŷOC$�P`b)-"e��t��!���+_�n�?eO,m�������$���~p�3)�S���pCZtw
 ��~�E�$�&�S8d����*z0,���r����H��V����1K����҆D��%��sg��&ǂF~#�()i9:Nx>���c�@�3D�>XlxVHYEB     400     150�<�@"���3���4&F�-)�D��(_Z(������Q�X���g*�Ɍ���.%�+/w!��a84� }�b\��m��ī`q�x���*rô���#�F.IM��G]Lbx����D�ub���L��BpD�iaMZ�^�2��@������ƪ܏�P</du�΢�fS�)���@Ǡ��6kjX÷+�j��!W/Z��Yyui���.`X�����5�;u�iԽ���:w?
��G>�4��(�^^��6�9���GTwwv���m䋒H��[�̊�}� ��Q��#�B6�
���!R#�/��W��f�����ȉ�P�i,�:����寲�>C��XlxVHYEB     400     150\+C���#�Z~م��ς(a�V�w����|����Lj[��Q��~�tӝ��T׫v���������N�d4��Y�(E���"�{eĨZ&E�]�8>��0�OM��,'A�&��7 ��P����|�'-��c��ؒ�>|�3t�@��S��H}z_�0йv=HvŅ48b-���*�+�㐟�	�Ɣ�IL��d����u������:`�@.�������]R����x��OW�"�]��V�b��L0�*��=����U��]�w�8�;��+��TV���6��nH�����z��D�
��JS�I�j�q՞�C��m5#�wXlxVHYEB     400     160�YK��M��W(20�0c������Xo��PR�&Xy)JT�$1L�E<K�D����e�U�$�6/I�G�;����wP�Ĵ�r�\d���N�X�a��Ů�[$��	�|���Z�g�w2���RZ<��H���&������� a�>N&̾��e�2;���s����s� E��3���(o����V���O�Ɇ�s0K
%��>��j���,��V�	� k�2Ⱥ'	<B�<�Pp���2�9!Bi&�%��DK�MU�Ctt� ��c�kU�5�[�-������f�]v`;5����¢$op�	=�[����Ь�b�z��z�kV_�m���=�XlxVHYEB     400     140U�TУJ�*	Q��v76�m���.����3ݤ�2�z�J��$�b�N���yV���>��̉nKn-�(�|s�..�^�I-�����k�mejt)c��'���r���&,<�O)�abYy�Q}w���= Ps�����.H�_b����O���}]p�y11+�K�6��őu[�C��ju�3߳��'8	���c�&|�&�P�H����&dyz�+��v�s��s�z$���#��%�>�H��>E8	�s+]�s�J�&Z�v�J6 ���4,{u�X��t���	w���O#�2N��	R��{�?* �[��Uc��ƦXlxVHYEB     400     170�Db��_��NsyIبWVc�H�6 %�v��(�ݫ�����U��Q����G-}{֎:��\��O--�l��0�f���rĩ��i�ȹ���~�*�̘uh<�p��5"�	p��������X]U�J��Q:���`i�|z�i_ߗ���LĪ�
��`:AUUR'T�@(�>��l��B��.Si��}AC���\�x�Y�i�hކ���z�}*W�(F?��)��K�r��]��Ѻ-��X.L�B��*�^U�C��Os�P�M��A ���z�ၪ�����	&�0���T����~�;��M�}�����ֻ����=�r^;���D*�)��i_��GRF�H��XlxVHYEB     400     150{"�#UIb>���E��g.��8����Ep[�\��:��Қ>��9��!�V%��n���	(i��e�4⽥�ђ/�]Lm�7ԛ�n���ߦ���?a�󬇇ϋwcba�#޳���)��8�T���z��(Ϫ�E}`���G{�mE������_��f..6KP��*R%�[�#�7��1K<-�3�{QX\�WA�`GB�@����5�BH��^Q^���:R�=�o�T+�$���L��+x�ϐw0����������9�9���ؕ�96T���]�,efs�Z������SU�P��`��O���+�N���%t��q��M�b��3M����t_XlxVHYEB     400     110>x�t�*2�rq>�����j@kZ}��B� en�$,�#����je�r���[P�-��[�u��qD2��bB0�	B볻#�����o��
��������zoF���1ia^T0A����t*]�d�m8E�����!=������Zc�e~@[XϲkĎ�Y#�C͕��r���t���ҭ��rBKSv0F�g���m1g5��/��?��5`�I}�nS�b:��1-����3C�Ft�J�톟���������-�XlxVHYEB     400     1507&�9��L8��$�q�i+k���^�_M�`/&�T;-�z���~����t�/�t�Y"��YFl�B?�g���7��"���:��g����t��&�*ѷ7��4$@�]^�`�t c�����Q����iY���T��:�������Y�En��t�?&	�|��V����� �}퐏�l@H��b�ܜ��>��lH̋{Q7aJ ��t\�%������Sd�׬�?c���f&������������%��V,{ �q���J��5n���^���P`B� K�O�8ڤ�0�B�:�ƶ��M������<�e�J�a��|�-Z��^.��XlxVHYEB     400     1a0QOD��uG��"���WGT�]s+����j��Q2�=#���� .�Ό9t-"�:6n����*�y72pM8<t��|;nXV(*���j��(��w=ߝ��݌)[�p�^a���G���6��{���M09-C
E�S�;�*����i;��(��9t[��<ݐ�q2!�΢� 3=�KqT�ꭸ2��
Q�*���{�>G���U��ߺֶ��v�ݭ�0r���ɵ�s�lV+ˤ�E|�X1�-8:�:���с�O��2��w�����/M�B#z
�[O��'�Nf)�zY-�I��h�b�sB���	��㇙ŝ��Y���߭�ڋ&� �\J��"@��~�>���ʉ�=й�J��ՋK�R��]�G��#�T�'�߽t\t��us�G���pQY�:�m;��|�XlxVHYEB     400     130�*O;����%��@uYdH��#N�\��J�!M������ԬT��0̳�#~��,m΅3ۑ��=E;�|O��ј\;�	��p��L�=��wlK~?��!�?L�uM�u����̄���G�"�nd�trM�Fy��h���W�:[B��Q;uұ�ٿ���[@ۀ����d���r=���r�/u��lu��I稍����I8z�X?zq[	wlh�szU`��X+_�`f�<p�=Bہ9`��5?Y�o�-`��_H�^Z�i�nÅ �Ǝ��5�������Y{ݝ1���g�Ew�|9͐kP~��IXlxVHYEB     400     120���gL�'SU����'% �x(a��c̻3_l�?���y�
V�F��Z��\���9��͛B�Ħ��.Č��>ޣ_Ł�+��oWfG�q��x�X�[!n�y9�����{�[���z�@��`�D�	E5Ms�5��6�S�br��#b���] �["U�M���H�EJ��	Ǥi�+��� �8l��3�Ba^(=^��[�!��o��qE�ǐ�{�k�c'�����d;��ɰ��{��+�:-4F\=�[�R������db� ��vL;}�dr�~�b��)XlxVHYEB     400     170�v����(���^�H��Z��*ߌ͡[���|o6�30#
U�`������Z���0}���B��U&���,9Em��%O���hϕ}j��z`������J�����t����G�k]��+��������Z\���-V��E�������w��9���j��&�i|^p0CQ����������4��Ԕ_	�74[���	�W�An�(��%SP���x�A[p)6o��1ey5¾!(�08��ICt�]��'E�[�\�wN:��B;AL2��V6Z�m3k�1�pH�	��2�/#�&)�0�m�����9.�8mG���׷c T�v�Z���w?5�N�X���!,SdV1śJMؚ���XlxVHYEB     400     160Cf�]+�8�	A�:��W\��m�[��p�K�gd��C+�0�����v�$#�~�ئ-3���fV��{����Ê�7����`1{E�4*RmD@D���W����F�ʭv��b�P9�ɺ�I4��������t(�Kk���{=�_bVͩ �j¶�^�5���"�B�=Sp[�.�܌�H���� ��P�\�J0~{@8�I��N��얀1k.����Q#���+����5ŗ�1�᯸�)��=Z�:����`O�-~t�ܑ>?p��.3�g�E�BŌ���ᆆU�	!��p�K'Z�M�l�8��[����?>#ߣŪ.EEҗ��e�Px�7�{ʦ�]XlxVHYEB     206      e0�~`�{����S�1bD��F͛y�r����XG�`�Ki�z�kz�hڶsdD�S�7ꄶ��U�Ec�6yD�0#n�^�y�7�p�
���&Vp_�.pg��x;BX�%�<`����y���e�c��{R�$_���$�aż��V<;��kV�ys޾!��װ������R��l�Ǔ!��rqc���=F�֭�*�v��cn풵ʑj����&y�u��