`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
VGRs/jcDtqg9wFsJmISV2bf1/NI+ayYmMm+6JxYTZdKtC2kC7nRf0oZNdphOslTfYrNKNd8vGM/D
911hhVbRRDF36GGcB4LhxejpuE3tlgBqgyYz3xy1iF/m1Q3OdZTjk3Tcco2UfzjuO7P+PBMxKtgM
6hf2kb7roxP1Z5DrtOQLP+YmaBH/nWbQRhmabqnG+9AtslPm3dGzqaQM1rToovhvTqYkJry8lY9R
z9HxgYGrx9A2PB9ftyzBUvDYcK1k4MeVWSV/FbXdG7mZTwqeRgofJD8RfN+QGC+0+4Mfw4eac1kp
d8GNarjPAB6IZ4U8D7OF2TexTe78IkWnT3owCg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="I7UghOUnofLqjKpE5QqrriKkCz8XdJ7pnoiTvr8HiCA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17984)
`protect data_block
13L9+9pkZ4ldzqWlsvyi+8VdsDVbcNiXKnctBIQtItF35gbbIWFBxrZBT+yGzu0ARRLLov93dJ2v
D1BCKGQajQVXb+ItYEsZWSaRYGqEbOrCSE9qxrUgfbaJBwnOEIiY4j2P0QZ3FvImGeWzBtNriEa3
m3OJOo2+qBEP19Nq5mxJ0dLgH8kh55Goe8Qc5hwOF0I2mfEF6KCuSlT7RUjg9KvHu4frfWmk+jKw
EZuccTdNxOk4yuopmihxXNHO67byv5Xoetp8TuEUPt+X2ZWwkHJiEVrRxV0se7PEqk5RkXUm42qa
xhx3sg7KRFfh/8DeBctR35oM+QrCBxwKbE1hdD5d2GVkEXUaYAUX7h4XOfSB73cWF5TNw+rxqshr
2PKhTLDGx1vGelDil3C+vf12ecwxEDUV/DYpAj9wURr+RTX0y58Tt3+Zq58nnFGV9lrPl2qCium1
IzSLt814rRdKS1Mdd5EnLG2vJ9X21vdGHl5jHxiRqYNVdvL4sSWQrUwyTaPviqF5Pf3p6mEZkaxb
OYV/Q9XD0iu4Xq27aR99gIU+M8RAjCGWwlG8Fo9/0VxIUPfuLHNj48rdwAWyrOr+mlq3IXjA8piG
/y2WnhGTRgahMdudfnZkyWyjHggTFkUGQRyDyveCDR3fCbY/qBJ2jotsJ0NbP/ARbzqej8oUKtTn
WX7WGRhBh8iEEWkb27+OA6z6UtVEeutx2CKdZfaWR976SnFqelryanpI0hDE1IX2Ln+y6e1SiK2X
8gILaYo+GvS6/h5mopMhQ1QWUfOvCBWQrHWhLcMCRK2lYVgfUq3xPT0fF/bFPMl0hOu0b/LkmkJk
ct4FjfrzmxB/p6PxHpQO8I3IOKmriFBmB3RvtFU0HSfev/HUVpZiK2aZWDY2fwIlfoVStZrA/E0p
LtT1aaMTtj1xAQuA7UxGPGr6wUG8SHpDnZvC4WUqlkKIRooLpOs0SgfJO7FvQRvH5lA9UdKLL2rA
3P7VhxIuqOgLNEf1+hdnD+4uhtIxcq7yREm3Drct0toTmzH/w7uOmx6/rbP7d4zQbGqjGYuFBP9B
vUQUwnPnSsaVyBnk/FF3mA1QUVumYcj2vwgMgmS3Ob/dnREcLedd/FWs1sU1Lyuk1F0Bn+8IsfhB
+v4BIpheiD5szNJqIvh2X80Ul2Dks1tB37gESLo+MuRdwbr7FYvjidF5/BreYuZ+A88+B2AilMVp
b6xhZ82XE5RIeqQ4okDWUStqnHPENWDPVB9nphl+TTkcEHzofmBejysew+lrgApFJxJX/ZCXAadi
Wk2tYXZ13A36mpQMVgxrQeIvPyhu0urcgvZzAyUp5zwvooNAwtWQm+vCqZHfrWqnxxT01Ylevd01
kam1A//rhYtqYH3UoSJfCorw/DB67d58MiR9dtXanryIYkMgVpp489EJECuPgrGL45xD1asyr/mu
WSlfFqLLE0KrdHa88OvOXSufTfXQzI5QpylN05u2CADGfN3Wv+9mZe6IYKWmmgx4H/O1B6GYNHtl
2AeGy5uUi+VYC7xSWhB1oGxQ9NG80W+LMB0qm8K183ENYCxsms/O8wOYZfeK18rcyKwS7fpAqH8j
5rh/D5xHU71f7ZJYbP5w/l4ycbiv9iNmwMu9PY7GC/e7iJhxGUx97ww09JPVaKhPMiBJAbnZLewQ
8xd+fOGJAIfcwcO02v4VaxjQbcDZwY8ZgTb3Bxv472BmUjBmaOc12mRS60dOLn2Qmr58ky3vrley
BwnTqE2GY/B4olvqT5c0CMBNFUaktkHQ2CLu65c4lmINyxBbU1XVrFj1ZgzKHqK2dpHA5XINaPbH
5iDI9S80A08P50joi3ZAZsxBCplrpVu37owNWsscvoPpqY+VUEcOSbZJBL5S6IsECdgiZ4H+zkOZ
5lb7vifLl+VL4HMKX/XAcsOMglmbuYVu9LgbR9qIa+d+zdxQIj08J04zcPy5iGHZNXHmaqzX+krp
16+qBvynb/L3UDgkKXyKEiSYqe14Ivi9qEcV/tlHkKvS7YXDSQUZGfo7mjG8TsUffQFp32PuF/ZS
PVKqV/sPBYX8biFneXhvuPdqliFuOLK0av8CmWuXf9KW9vFZ92sxj0jcB5hNgmiD4gKE9kvp8SOH
jjy+A/dVzn/LUgmDI5i3hdlAy2IRc87nhkfEZkSnT0NEpA3HAmenDtzkqeiImGDhdUN3ppLsNONU
wzur0P+klYnSogaWsswXWqWy38Hy8nBtu+h6Jr2JGcOb9OFChZZz7voyeIVNakadTVQbgAMe4KCP
5FV/hHY5VUXB/+PXI8O+FJxMS/6dksluoAm/JgK4ZQ2GZEKile18MkFGgqRD4PZcvOXFlB1+3cb3
ojsx9DKk6mzIxM5Ma0WX44Y3yDQ1atE8mGualqkTw5nF2A7DK3JKL4jxrd7iTSPDuliVtja9OaRB
HIB6DxTfELVDHL+zz56yx8GI7uQKlKzaZ1q9SWPV8AKfSyTB4sAEdqnqHQWVlgtbZWsdWZdH7ohv
66iDMXdlFUg5v1MIxJfbrlaYYgGsM3CcbkqvpfKBsVOr/ByBeJbeIKGvPwLTft4aES7h9jxD1aXX
v/smdT74Tm7zxxzB71ZwkMHvu/ao+QZ42NUCj++r+KrryQmeZzdSGn85YocuZ6+tC/NlZloJFarE
zCGhkL7VnVkT0ngQHD3b0O6KN9X31oGQairvydxAW944TkhKKmd5TyhrubfeZzQ9TUVkEAnzXD+p
Xy41MYu5XKHnmH9BxeQn79eJdMVLniuO0/7VzhKklxHw/TVK3cXrz4lmIYodwIKNYaq2N/nWu/r6
ZF8nZNlh8lVNsJ1ChaiHhU7uGC2oJr3975q5ZXKcvk7tMoWVU0wxvwd8cc/F6pfUcXv328FUJ9YI
pFtrQ/zdMnlnQaejaj+4opyGWNqv7ZfIkKMW+LD3+wx4nW7lUQCZbfeVu3/NHmc+klx01kLC7Twa
A5QCNeLvbgzr4Tx57HBhvqf2BRPJ73aHxssW3HZBvkAHRyb+Yji0sPwOVHuJ3MWUcDlMONyELprG
0hLpdBiA17TQnWHxuqnKuIVAKAPUaDg6K7ahPR44adsDewiYplIRCk63fbMCWXDMFZPHe92QTvhi
nme/eNXR1GNr5RD8Q0wUxEal03juurx/k9ROzED5Iv6tuglJQbmpuSydIdHfFW3yLDc33HXqWFIR
JPNz6oQ8Ha50gRIDS4EXuD+ruCR9+BS8x3I0+RTBe1r9PU2k0bA5zm0nu/5Q8JX9Eoh/TuYk9l2l
eMxkdzfCKy+tOql60KQkpRHCIO4aoi/OqeFDxjV95uExk8tCj8v68QZahQqAwJsILNtCy34epuNX
u0CrK7jBx2GAr8eks56OaTmqlQ0HNYUjdZcwCB0b/F4tP3sHriwnxKEjSIYQF+atZE/Hattz6QR1
Hv+xTLYxm4VJ8lRFPFJ9+XRoO4fQdkF9aZnd7EsK5851zcZT/At+gRxQ+dzVhnFa5ZOr7guCcmjQ
OYmRMyhhX4KAEjsVKcymtdK0LerCHEQAkthOtG7p2ANTnRr6ikOkmq19Inps16oH+gSokCrgq1PA
mdtdMeS3VloMi2zVo7BwqlOeQIjNCOeZWvx34IT4cIuT7WAI4XCxijRjrcniNHZMrujZVZWhW9fy
fwFqdeTy6FxFQcHIAjer+ph1ELmCBR8FD2IlUuMVrovShsbqyfcvzqx1TpVSHtHmZNmrgH04IThS
fbHgJkEIOv10rYMgI2Mze1ERg0X7pOpu/hdEQbyfRg4zHL4LP+gsr0UnpTFwEtnbMjG9zRA8Mn6L
2haebutu/BZr7m4/ZzHC4h2dAia2m78ixiILLnN2s4LOY33D23vL8k12RzL74CfqGMrL4iVoFQZo
YPovMyNJijVzCpT3RTF7ixDubskvMQZLq4CSyiEbY0zNfje8TncD1szWcIZQxLnHAoOL8FikAIrh
Dn+FZcN66zjwFMOdEs3xTzBsrLEdJb8NxCghgsaKwiOLXlyT81m3cyesTmCyRFDE7UhwkrMNqkES
9PtvW1xDR03ag1wxHQ2Pknz+Bf5ZcgH0mWYNf9N08NqpdbCoVt+Oox8nzphvl0owOv9BiiPlRALE
zbOh4LRdiw4ne9f7BJ2R/KuMe4d7lHoYrb0NIYfPsP3KBEf0Wt6Uw87JZB0v62B/Rny2QpThmDfH
yMf4jGmvlSYSYL+PoqLiROZ0gDLdORjcLQ02g4wVx6IdVMd2E/ybLL7wDHQ+Q1rDg7Y8/I42MP2V
kzG6/4j4zsnq2qlffGhK234H7etZR49yf/lf7GYbZ6djVP4IgaqfPOOxZsZzEzM7liSzY9JjFeYu
yl8SJipZzcHu5BkvmubE0NL8FbJgzhRssOjt5UfRMWZOP4glouhTHrObDP7uiIJGzkDgfk7dGt9L
AvSK6Su/pSsVRdhJQNdY7QzIAA8Wmg7DhKo8AIQ0sLnjI8mbgg5Asj+/v5GgwuR3T9t6tbQyARYh
fL7EKYJM8M61yWjkz7ajaO0iJlC7X8uns/vt8Et2sPQZr8EuVUf1yRTdwkt5fZH0gleq6AHbyoiz
zqXkxajfzzhvmHhf4pXv5Cos9efogmwrenGsXxMhLbJtz3vgpI1rjPsdL8tXOFef+sUvM5b7qvw6
u/nXRCeFXEv2vEK5JOEZKzu43iI0vIOzsdC9ODOktpO10sZlqDTFz3I24mOo7nBbJ8Fid3t/qKf2
hwBGG6Vcz/ogNYCecnlHv3xacOINOZevpCPJJoif8wfBK/djSaDyPV8VHGjLcf+F1hvPMdbtC70v
0wpda/bVlublOP9JSLRZENptlU6xnOGBYxTYBIL8h7vbc5P1XbFI5T+RwTGSTsPPkXX6oZMBMkk2
B6ReFolqoA99vkWBit4KPB9P9lE7GEKCHSjJQ6cO7y/YA1cPfpW07UFpChOrl3McjfxrjA7KOMXz
1sTvJKSs4woz96SZ48DbyewG7sbIdxCK8zmJzPiZodhzn3Z/krZxclsW2JaiIfkLgl/TYMOvLyFn
SS8MaNcEaOqZQWkJNXhkN5UIxnmWEYP9+mJBwap/d/miwdEr5o8VHOfT9OrX4fEkmQsrotqXy+mn
zpUkRmG/JKS6p6PvdOtQDIkWiOoSSbK6AOOFt4ZGQj8drC3yhhsANAq2aSofPxe5jJxTqYcDkn61
lBNZprClBcf6aczrdRFobOgAMTeQz02u0ApusmxPYa/XO4gIQ19VeKD6aJER64Zawf8E1YNch2aj
8wySeQhoeQ25jBzBJfTgMvf430IfmK94dLmTDKE+7Fic6Ro0Ifi5dxiZXjY4ptQzLHLRdepIV5ZW
lKlqDAQGR8kb/Z+tQZatolw+RXNb7pjpZRM9Nxju5nedX1S3miZaGfOdFFN9Sv7RJZ+Dn89k34p8
3+XMrwoXkOOnj5kaXBbY38EOiX5Samjai8SHKqjXYZ7wJIxSTwHQU6HQwfBCcfTqjk46yaCLZr6j
6asz7IQ0QgvkfiTJn6K/nBeZ4pbLv0zdwaokv/QJvy872MA1ENJTtTisxFQSTf8e33lCIHFI3xSC
GSrDjNW7+aoiIKleDOnyY8mY/8bbimjuXpmrdyxw/lFZ2e0yrXKLFXKxGMpiSzpqcCuNHhdhKnBj
chTVvAdnMbQChXtE/0yjKmw+y86hu3fmaU8JRSiduH1Kw4lJPbaq9n8ieJsWJBGTxLkOF4lXtit5
Gh7PIHD/rHYxZp2S1QTh9aM6e6Ye62aQO4eKX3it/0whkZw4AW09q4/1EkfAHL030sgFs4aQ2sIK
LxeLnIQnx8OKbKKBP2Vtm3NF1By//my+BGfrmNrgGG6FjZui7FyZ6zXLZQ/qWizElqsA4b8RhgyA
rEJcfbkYYrvodZkdwPer+PPFlWth4g0Ipx5R1Xq76OYcoaBJccEt+qwvGv+eFQ6lI0bk5iubASTu
K/KMJ5zVxCEHfIa1s4Mrf5JF5Be+0Hx0X6a0hN3b2MLxM+GUT0SnnmJj7Z6LV+b5xVfDedvfTi/e
td4AcilYWOlAfl20o3m9Vq1JaqeH4cFOI++AwyX2HtQmjxZrEADo6gr4VTULNNvhaBrKDgp0744Q
+Ho4426Z8fZHjvVLo2fWvOGXt6M6LfVLn5quoElRworFcZVN2KkfQtGc1mOLVvpgT5oYfiT+eM9v
31c7vl+j4h3lxZJo/SXLe5T7X2bhljxdPkm8xMj4ITFScXHWWhrXZwxsRgGJmCSQwBJ7E2nvOEuz
9EIBYv6OJsFP75sbvUrGJwIbeAGwRyUvtUdeZoJvI5YKxW/JmdsXaN8SJMSyBPTYoZi9AvibtJUi
TA04+THx16CF3GG7N2krHG0UHtQjcDhg9yVdanEV1l5x+KMxcB2kUGrygJwKLnw4LPGDVgcFqE57
71eUpRb7zvnKqsXAhm5BT9arqLxn134QAzj1WnqHkPTS3sEMGxzEFOZMDGo0lKwBw5/GWiG7/Twk
HRAcALwXWSJsE8bNR9eSRsuZ9eItcUQe3/46tVVhdi7szNtrAU+DNJNqkZN4cNyfwu5hKvGlj2Jl
eA+kvz0kuslW5VVycMnj0Bl4sJaUH6DhJmtfVTBE9sI21x6AkYDE4nO6zIk9tTvwipFWuvnnSB5/
hCCiIxt20h/O9jf6vkWKyl1k9OFyE9doAQohMkZSJ34PfUMhmecWDN2JComvWmgxpy6doDcWEFZf
PYk9Q9itAlk4eOBu6gXRr/fNzBdDFRgnonWYvdr5fBgRx/uVD9GHAsDWXeyW4CohAnyeRCeR3DIt
FyjgIWd9KIwT+C1METTCis6OHNILdAAXWK+sBiSf4YF6joxFTj0AbpAxbMWIyA3mzsQb0Vwlc7pF
VB+8jn+Y/dyg2fuPCyyW0yatvJQq2FwMMuiUEkSayXt0B6Im+nQVYvglGh7F9T7ysYEathpgh0Wa
ecdtC3vc+mHuP9cTZPJeqK+6Xa9Eq0pH/OtnspqqMG8loZ/F5aWBEtyBfSZvJQegGCw8ciHOinmI
caFgx4zlOJK1vSukiAs+BlzB5ue0loutPTrPYqdHeQRM9dWJIZUmrCVBsNxiO+bd61K3BXJbXeHL
96+KrwKbAW/cXq+s2tTvYpnRxBQ+KZ/sjZS/DprAWcR5kU/QUjCozeS+LgND24UwUe8f3Vbb/ozt
noLGYfHp955EcEOVFcip/hJsHmxgCdGG+mJUJeS84F5WX8OETv6JfLthKfKqjlPJ5Nvd+lgRoADR
jjNaQ5tKDQVRbQDPlKeQxymJIm2RTuSRHUjrC5uKItE56vMoRecDWIJBet4xSaQpK2UT7O8Hvbel
peD//Vh3f9jOVvjdssrE4WuWb0ZRVm9vJ9PJSuAcUi06QMMw59tiTBBYMRiy8dHwmXadnOt4zu0M
58udeMKOYsNhwH1VOGQjhXeB47qlFx3ZQNr55mfgEhEMbAZkC9JjrN3fsApbhXjG/85cHwdtcDWS
Dk9+cgvK31xoUsIdMOi457LOfeWU81hIx8qhG7arEeqXpEV8qmfdn2LsWPYuYd2JHnGGURCXBtV2
DORBccYdWenlAOFmL6d98MYQp84tsfQxOyy7+0jbveRnb+ivc38VizLmksFZ56rNKX6yFBihGzcK
dV3LkvOxsLs/fWCVL+uPujq27OrsD35z/Prlz59OdM5WRxQfkwIwFDMlpcSNeY0SfuoJ6ihD4jSh
Rt+nS8Yc/DXdtKZUtvs9TvU7QoTmMgnNF8m7JgDG3m6od0eiqxq2/3/CIu4oHQynw0K9XFEBfSAc
n8ZbI9VgJFCUQB/KIu1k2Dkukow/ME+1GtPR9f1p+1pLrgAM54a+rBHmzMUB7h/gVsAEzdNkY0+h
gLzzqhQNYPVWulGBShfi+fJl7X5BFFf3C4eIxFxeooCs2rbiI+IKb9sbO0d5OuGseBBw570qN8X6
QyvQFIZDVFnAh/yfqhe6FpT6XRkTMzSCE83LfCsMkkqMwfsI49x/xejH9opjrpwc27nnJvqj9GaG
Ald9rjMcbxB72+MX/Auvdq3+8mU/q1SWRNxyVHg1yEf0K+NlorhdUq0JP+jj0mwN5cwmjTVR9uch
82ynl2EW+WPZ/kUDYTQ4qF6A82yiYpfXp3he1nGu5bOLHgwAUj1/HIRtf5GBWIov5mXjW9dCdehx
GBa5yl9ogDV/xW3GcmfA58kxA+3BikxivoY/ZOjpGWPf/3dKqgK+qQsMOlZGm4Ink5aDlVmlraww
d0PD24XracxpW5WCUXD6cBM8aWtlepJ27QSdBD7avvMSaJ4ge/jqkhw/kDt8jc50AFjMfiLS+HXG
465Dxm/ReoSGBE+qdDlNEryvsuT2tVbNJwPBtiPzTHQF0Pb+Wm7hqcl9ai9PEj2e3EH23bMPyRad
cJTzJQ/z3UVRLC5O9kqeOsY7s05t4DacSSBzeCsHR/J9rMVg6d9F3kq1smAzMVO/fWz3QhI/PiIJ
JrPEii4afbpLc9brvacptBX03QLs7tJzGyrMzSIAZ/05NLNwuZoRB5UgjU5pT0u5ilxHpEERJXVQ
hhxxT8JvG+iJCOJEgpx2X4AzM2Io+hHrjrWk/7xSwrBQx6fT9YaKVBY/Lq3bthnEl+7+Ndj65giM
iITw8lOmp9f+qRJSykzwB4E2mlYgundkLnGG7Zu8NxGOURSLAaOO1f8wcIiwfBHxhMvaFuiaOule
aOQv7woMbsviu6cADvwAQ9vj/I9XzxvvD6XMfLxq/9MQYHWTZL39Y5hAcnscyDqoXbGqVbBx/F7b
FdqhkaCBpHHhJZqEv7pCYlL8qcwKNjIVw6Rv4xtUUMn+uPqWfEYjZhTsE89teDhpVqzW2/ejpHhu
/PxKOzeS1GlFFx7qLE9cSPFZiOwWWn1MkQRh9Nmjr5f8lAkRaLyoXRs+mgJhFS0a6KW7+HEsxX2S
SeuI32+vZ8HatquN/z7C7cGVVIkkOm6s+ryCeZPsebaOzjv1s5BGcF05aNab8z+uU5FQs3Ye2XC4
5mEff6SQbvAHnt336jG4GN8fkwbm2x3OtGltikwNGBz3Ptw8nV+MT4CDEj8t5QNHZum19kRo4fOE
j4UyfJJPpSZakLF5oQKfXuj4ne03/5N6b1x2iXjuQy8W1a4UMOBLQU3+dv5IGq591VKSMJVHbxyN
zqFUY7ArIaOOFviayBD5fmHNWOxJi+689cdxfKpULkQyfsZ3RQRydb//2SBBXk34bpiaGoHA2Sf8
OQTDhmp4j4rihdMOPzaJAgCz+2iqy1LY9I6jP9Lk1N8k7f1bJw/0we2dxMyJcWiexlTr6hE0oFh0
iWYKMDgAzHgMHfbFDNFgqMBtNp8yyGP6wmRgCVNH08ADrJVeJfefEGNIqDH/YnyoxLYmRO34iAAb
Vd7NKb6yMFQReJE/OAHeZbZNTwxKYpxj++TBsCYXRiEvLxpWd46XeiZ98ejk7zKYnrj3WUqFEdPs
gnGMM+L9Drcy6GWi1WX1xbeCsZMeK0sUAjjF+uoa7NXcOXbb3+KDFZ/MM8XLb+CHuYhY7J2MXg7b
kFJSRmKWkPwmwgXEnXtyCzoGA0TfdFP0PUgoggsilV4Fw7kA4s5MdzyUVy0Cn+sJaiSGQCBOPh5B
32BDjn9ajA31qf5vSm/PoomFL9WtlegylK/XRFOKrz/5oNBQZeHpVCDfypHNMYYbyc7LWzao7z8C
AMZxmVBBQJKMCwEE/Oxve32By85JYvuI99Iwg8TRd328AGZnLRZwodvdE0MOCNhKToEGS3FBjlPR
5xsoNSCQlLn6VSAwikKagaUp3O6pWfrF5QHQew2cHc0nGExUQgixs/EKk1tnqic1DnBj3MGBQQIy
c989LmOA9AL9qRxSQ997QZWAtGbbM1tvmgRPdwvycMyJC+MxtALxBuRx/G71UYyrCZctVFyOgweD
ZdlStlojrY1al3//ALc1ChjP/DSRtiaEtvw8TNYmRe4EaxXS819lftE65ktIjwC2P5HzY+i6eDU0
9wAItsE/nvGTkFpNQxfec5NznF9Sp/bgbR/xdpNcYXummD3l+P9aei/gFIhqVOH2+W44Wyta9t0Z
/ARy5NoZD32nqIN+AeIFhV6MnbSiQjpoBhvtQPaSxJ++43Xu349lcxrPHVBulW+WaCaadULQXcJK
oe6jXgeVSDWKj23fdlotPpyHr5RCvguHStvkWT/3IR/SBmsiEqaeOBqiOoRm0vgmHJyOvg6Rm9E/
Hl+wDXpl3Mn+WAJWVlztlArOicPktzjxF9RFrgLwH+XSIGAJWLLZSAjLlpOW4vgPUSwGWnxtwpF3
c6mXCKmZ9eVgWcbnBDY+9VIAmYrZQgT6Xghl2iDxjUGfQ98Scl6WJtkfpSu2Ng8gmCENmoKt7h+7
nv4P/J60+vlrMADXweqzxSvBfYeoyyLb6WWEXwCDzO9q5PGsmxyzoIjuIAAYV+NsvHe/npmlk7hi
IS6c7p+kQHqnnoGNFMXdHjwAvN5VU3dowxgJIuCsfcbvIDHH57dgBkNiJlYXcwZ1aI/CW29gkgmJ
qhYS/zidFi0jzR7RgZoJHU13qhEZHW3RKHhZTDt5XraC0iG4kMhmfuNMAtNvaEWpTA5qiATl3NVs
ap3KLlX3NzJJAWIlP+z8QYQ0q3/sI8ITp9rRjSFEf2vcCApOnH3QpU749qOp7ObTUKvkdYE+6HYM
oDEcRUEXxpbG4ODlumRkUtcna2mEJSgTVeZFBD4oc0yRM6m6xwzXdujoSaFhusaTwi2MH0blYGoi
OqTaumtQ8cOppm9++VLVmIt47BvmK3lXFo80PylR9+wQ4WKW0LE1R2QNX+RmzSOiWQ+Q+UfF2oHl
5KKGjJFCOy/uXnvry/uyEYZzLXgXAWQvXFDuKN+CO8uBWo5M+mbXnvKsDMxG3/6bn/jQzn4qs18W
ssMplzC0w9sOQkskPdvGJweHqatP6H6KGXx1a6UNieaUkPlhlA5PDMgDPYbCi7ar6ifuXzwlIWBg
EP5uJK80VzzUvVO4FlrMxnTAM86+3rJ930bAJt2KEEMTAPXL4GbehJ2FFEfWVA3Bsm4BwypBBf/R
uwl+R9DZ/9eXFn4e5xz4ICnj2NpItUdKWo1eSetPB+QxZ/jqccs8c8qyNdaLHQxSoiOmUfgoasWj
b6HCTKYzDYJv85+LCR+h5nkHUkyBeltTk5lz+ztnz+PF5FclZxMNW50byVOegc/bJjbEbV63zXgf
lWBLamuEVz7yjOwSfMcPpO3h29QNgD124pdCbY2oGQMikG6yCgtzjRX7EaMVqRDnFHcro9T/xkqc
5+ReFjj0OfkYpZWl7qqctGs7Dvr9+7GOeZZOCTSr3vtzcP3Fus5tjwHgBtwdxHaJLRO1Nsv7Cx97
fyOdNsu/2xxhXpEgtlU+FXTm4hetwLBwknXiDP4w8qm4YP8jxGZateCVRk291xhkVAAy5MYcfCE0
Kj9RBNF1y6nUtP0V62yjxX+Ovwf8TNdzKwxyhHncBQOKaoCWpgYwPQS7eAGsi71cxinqFE1UTNBA
dwg0f6v9UcnSO6jS3DnJIOlrI/kkOWOoEnzVV8ZivKLGPrIB0TKODGDrV3VCs8c78nNLmCCaSNS2
lbSy/UsWX6ZdWlBNfBvffcXaeobBJ2ULcZrd5YoMDuhshyZIOdUObJV9OiGnJwoVXGggMxOP/hIs
nFWfzWlq5dhvLgdVM3t6qNzr9oqge+Pq9Bd0JHwKHmfZvT63MRu8YahK4OhB9D8gaCGRTpmfzeGB
wNp64kDiJFJtcI4m/np/7p+2VWM1UwGBi2Bpvd2W8HHXTfyJWDM+bT2lYC4w5X91pqUl5QyVuL9M
spmrV1honm9CUzQDANxM5eKspK9vMNJs/gxB+Urf3JhkOKaTEviFUBYa1A/pLYrhPfeerKddZ+ry
1rVtct7hQFQJ3aBaGdnULxBLmL3XuC3tU1RXCoyFdSVDpSaFSjKW9oV2seN3qbncApmFxlI11bk8
kwhvy2AjjoNsYCWNrV5jee/clj6HuuF0d5fAA/4heMzDNrikmzNAxpwcurbZa1K3VVDrnQo1LtRe
o+OEn9ocmjBftNchmGUvxlUrGN36d6m8jdfxdBf5VUYL+dLTFRovtw1ABOa5lSekzaJFxIBnK4Oz
iGTfHgROu1tFyY2GV+ZRDWBTH3y5LY6yZmQOEfQYNIXyC4MeWaJTSAUEBo3WljYtdq/Qg2DTzT2s
nfBf8fpqVy0UnquGdWW/00gVzpxRG9ZFUFbGclZTcXykwqHEbPAkRTWX0PtxHbOlUNJnVagOZ93O
p3kSIEY4qvwnlxUjcKHZbw126DeoTTorRqCJsGWEjrMuGnIY5GWbEG8ddx/PdPGe6401z3sJ/nEB
jQZ919Y5r0PN6TDiZdjqcDrScuStWA1QFMpPJzTpWhhSweKx/j6ikPG+Z8bMODHbvqnuUcih5MjY
Z0yVM124dok/Z6UF/sClBf11oXcBP3MxVBS1G5AWNJ/lYFPO2J6C6PuaoVmsqZ5fjY2PV1VOd5Rp
F1dbgDr/S8ysE2pTkDNY+E36yzkgPr7hcxa9jUyIxsixLpxohAhLuw1OoeVuJy3OI403Jwgn1MZJ
h+wRUlr1gFi/c3HTgPlkxov349SpUcd2elCtlWq1PlPvv5X5nLOeWxdGmhqL7oTG2JC2c92jJaOB
MyX9NTh9h/kblZkAA5pk1q5uWX5kgjCw3YM+diCpfHYGdYCuOOSI5QcTomozLhgSHp/qOyyko0UX
p0ovTprRtOjKGnPgt+67iJ3WcOQm24ar811AN1jdh8WiHqlJDbMB7ynQLIJ6J2gmUFlLGveY0l7o
vhhj0aiUM4vPYEQK5CwKK93LdYTMfnRiwXsL5Fd8MiYzNrxMbFfSwiRfqgdyGbJ1dQNmdg6MbxJJ
a8FiHE8P76afmrU5/brMAQPpyuNMvWHWFqnYxR4URXW2VL9WmjmZn/NEpnqFF8DGXgqPyGk3qY/E
CiA2SOXesFOWe/T1VyMi+5Sa3t9GKnWCHRQE6578ce4ACtYm90pW3lNJXBJ8HBp8ShkGJXTAQtez
Q202BnfUTqTVYwQMx9zQj7xJxAYCrnJWVHx0txMHFDUbG2M1y/DesxtJO80k0cWpPOOWCzbbo6Wt
av3QYyicUQ0mpQcPQqVzucuUFv46Q/KO2s1IjO2/M3L+qmnAPBkb+9UXFAUnG6yIb5Zoc7KQO79t
ozuexO+YJ0RYDY+6K2M+Ed6j1EvoetlV4Vnz4l9I8XLGNZWcHxPpdfyMegpvxoZ+F+zy2gp2t2D4
gTt6z3M6hTImvGpUMeyqwFz3QF+d2MYZbvIscuxekJrqddtYiy+I5j+U1owC+cAAcqpnvqqtkHw3
QS9++jIT84cBkJB76vh9CllDaoI8bIdplCNpgWqQwlqfk4STKaxKbmWFv/FWt3taUPiL6PXb+XVZ
m0UWkwQ2+tpOt6CZAl4aS8AyNzRmgYqxS71I4Kb/XexV7CLSPmR6tVBVIi8RLvxO3nQfAsQZfLeD
TlcLr0qK4VaxoNPPZkjAKr6asSN7jDxyaNVUKwRwhOsETJlaAavjQJSaoxGwHo6WMJL2UGYE1ONo
5C9Hj7dqa6LDFb0w0T/6ZzFz5/6KLqacQ2Ue8fHmQxZzi5IY5ahfcd4DpS7jdLoQ75V2J7KCEku0
MkcUVU2VIcLJo1kwTNrf1RrHG3gE6G2FEDtsnNIOxpcOI+2hEFCL+b6VoCnLpp2S5XB6ViiZSANk
r9l6GKG1gI/pAlXg3RcTU35atu2miRasQPQDDlQKKKmlux074hlR6u3MWpGtmQHvo4/RSZW58rpq
ohQKcL3BgSfYX/Gxa3A8zMLJONFpW4wkvXTbvBDLtRNsyBtGuvoXHeUGTXp6isAo5iuFNpWFw01E
R+d05uIqgslI0OaIyuHFWSF1PpbhhuFzP5Vd0Dgr16qx2JCucTSFNBg/2zMRPTjRb99skmTSMrXl
a/gkQS0KOQ83G/f26Na+zpbjEkefo3VvnEKQQkTS3Yc7QsSsyRbRq+XM2bmzKd6otwSO6LYGvsck
qnhVMa/ohyEwUtSHmv+M0a66uovcDL7M9fHUeIL1ainqpi5Pi9O0RShs4xE/wAqD9F1x615BX6Kk
AbpOo50/4j6uUn2kYyTfs7UpoVa/tMC8AnrJ2/T5KaAs8Tcio3xr8BE52nlvl96xp07QruTu95ST
4OCsu7P3f2B5DpGno/qVodOcuTHFaZQnSEFlvW4K2zQnDtOXkXsP5OQiVtzeG1vassWHHZtjQDZC
ZMFE+E2Bca2BhHEn16VvllQMbicC9bYGc2QnXCIlvdbXLn9I/rW31OKJ/rM3Z/OsI/SvclHiZ8//
koWZonaEy4NytQA6aogFcZf7uLZ5yA49VAnpiIqEhs0pdNKpcK8L+/PFnIaoMbg1U1AKw/Q5P7Si
IceJvPEPvYp0TCYolW1+O3XTSJMAM2968DYM325O4F/YN0T2rYRGlDBiHB/ItwlnORHYMR6H6Xcc
0p80doe2eukCajA5SdgzMvV5uMd9HVJeAbyOtuc6upm/SlMEGjHPPHrL1D/CMJDP/SLhWoqkpPOZ
VF+nX09eyxoUfCsP5ipfdC2aKIOTm1ku1445AIST86cueWUskBt8I2eJvZ5aPTGV/YxnO93S/g6y
OTkaRbC9jX3jQ/PzDxUCxCuxxN7A53EOW+Gf8m1F+oCdRB7cmE0vUCvKjLiacZZ2lzy793RWg9Le
ey+s4TTDlPQpfKZpvI0WsqtU92/1c2rXE2rEJgBCgWv8YIxvhmpC8Ov1KkW07UiJP3AXFD1tVUGs
3zFSuGBgKI1T0aLgzWDaQWys1NWXA6gIPtQYz0GYs0pHpP+DTx50QT9vDRdyW9eKbngyfGs8bni2
Ab9xP76MNZpiuBUrsV5nIDskWaRgjLA9O8ZckqaXrHc8GWhU/q/GQ4aT5WqBu9KuygP/PFx9v/Bg
vyjxoqwvB+5jhwtsdlLt6BLuhoMoE/n9B4QCkq+NZ0N6c0XntdoDqiriPnpzwQHQx2chjlDZjSvo
qBMaq75KnxnKkkk/4ZaydSpeHTdpl+Sxxa+hTLcqsDJrYO1j/+SUCKXqNdzu8lKGvz8kR9lV7Y7P
O7KBhp51KQBVB86+/F8/9X0LVjOaktY9N64ekrgo9ksnsfY0HlRN3Ph/lju1ihIKjyobX+wLstcC
sxiZJAHUtt7o4lvd16yhAsy7YD0E766JByRW5WC5A/BwPsW1OakCsnyv8YmDqeS3/ZKmGmQP7pq6
jaKa5aWxSJ8RLn4lPzxtu8e6L8oW/jtkFm5mqeuPkvj7TW6OR/WERJLEO1aK7oFxkmtOpPrtZ4wv
QZV2H1lgz+xOF6ISL6568Hq6yvr2R5FIFhNaLrMQe5i4xlUK99vJctXV3HXc1fHTyDBESE80WMMU
fB+CkSzddctURqGHbwJ933U6EeVz9Rlc49mpg/0tM8YeoYsz8PgDz5KpfmU5Q/OOZVpipFxbX6iM
P0It2wj0XG3Chi+kHRMIBNFrlCTeaMnsDx3yqQqlteAjWIwpaGh7mBlyqFSndHKODRQ59uvobERF
MdSqAa6V6gg2BkfkNB3ixIIfM0GSulkNoa8VBcXUggFquCaK74+Pvsq0l9toKBiMspwKW2E/wab5
QtutFRSPq8UNomYqgcQvjleJ9QU1sD/TjKoZH32JDQnEYm1uMeZHOs9z8+G5gOB+fzQgeKIpfWNY
GheGxte2fwWWn9HzUDDlYg0U59Anr9hM/A1LPubnTYRE5DHvJNvoa/iE+z2EhP+F7yv/dl6YNJnp
C8nTdiHK3W5BA8AxgcDKfsij7eTdRsSGekdh75Dpr0jR3gA8SOKxtaaLtlEPx6lDSOEu3vv2A+dj
fbjT/5Zq+SjyP4P9iHeeB2P1I4hNnpuk6ZJYqJDk0Zm0wYIkjRBvSHo8ZNWq6rSx++ioOwH/1bTu
hE9YnuuCJVJsVcPEx02TfuTw2B8AswXh/zpPKvbTgt99YLIZEnggNlWGvvgvEXoMiNeFoaxBwJzY
MTmi/16j+lkwvWSZHamtPcPlrpBscS12EHyXlgOpJ1+hmGiePBED34FOgJga0uQpVGlRp5blWqu0
FsPrflvJTV1+X5hok9Tl3Py5OtviWE78RYFYCDnmrYPqwOqbDIP6qFr+R4NBoHpqJq4/IFGdmGHj
11d+uti5EeDAh9SWF1vUpzNxZPFI9drqtx0q89yCdJNMGO8RxJywPRi9ReeInHUnhxrKQn3htOsl
KPg5BZtT5wGZVEwt3G2oAJ4fQNoQ3u2ONSZEZcF81tG3Ff/Lip73VHWasJdXUd3oc3jwMVn7Ruw+
hieSIKgIJ5AtbpkrK6J+P4Bph2upP04b0RwZMdiTcuHVEXX/6R7OV1vUsGHb3QbqhlLDVFspmANU
s+W9U1PYZgi7d1gTko1wc7K8pWQ2Oe7jAc8HeDOHSKsqv8aryvxM3/N8bx7PoE1r3vJMcCVWI7Td
QpU/DlRxl56lfZYaHSarRWqeoFX1hROXpHMaQl6RUV+L7mz0/Hfbb1uWccvS/KlcutSnk4sw1Edg
AxESYXUi1wnpllz65zc1/bpv/a9/qtMlDnroONRsAMk59JmrheHGA5yx7ptSadCCRswrUwIU8BmM
u2QDzPNfIlOkECrjs7WJMGVknBzo68KMg1hnfAAnfU59kJR3711GORztdaqOqA0jjYI8AiTGCaV7
8l2HaaByIc1cXPkYavvjNeIOi0LIxd4oZQFCSEn5H6wd+PvyFM0Tv9f5A06SK9CmTpidCwO253YR
wgXehQbjlLYOsVb8e3GnHeJO7pHXdBxvDu8OMsfOM1C1xONC0K8AIDux9LW/BTDxi1a+ENqkPQF6
AtQvJu4fCvEikowMBGQNP+gveM9VGp2eBguOTtcwn6qYFbv0HmXVYTDBaVrG8b463nGpWUSwxL4e
hdfkezwVfvdoW+U5IYcmIgH0/tBtxCztXB0MtEDNWmTk1gPFOescbQlTtpPJIWMphgEv1wxgiDSp
V2+IfiUXODTjGyueCqBmPbCH+Iq0EjqawOFvPSRgPEuNlRniDS0fAvfe3VPBM8U2Mzu4hCAHN8JH
INoAP/h6+fuBMzjC1ZdA9+arkqg95PcaTT/T0d506hrelYTGn3hPb3E9jAexvX895G+CO0PIrfgX
M0KiXFduvsA1RdW5MwTnZG0F24T2rOXDizEnucWsUc3r9lj34xfDKvZhgk8HXUN4l+zzoqXyUYMs
mfTt8BEpVtHBs9Rmcnzem39nt9coPqigDABJFZOTmzeqiAsdVgZUq0Guc7VB+/zWXQ6EPFemPj5z
tIsjsh1Mb+r9tpAhFrlZBs4ndpfQclgAtTav8VbLI7MdN0dqArLRImf5ao7GTlVxkk7QliItHKoe
jlKrGNI2d52jGAr7Cs84vVEe5l5VyaC5Bz8Z/csEgYbuomYq6TvMmBxMoHIZ+f86sFvtAVpDEN/K
VJlEg537Cl5ebfDvcUZL3CHAPtLvdvpfnSV1yJHyu5T3cd0zg2HcGHohJl16U9AL2j7NamhI5C5y
A8jo4Bm5qRy+5jlLvZP8WV5Dr1lovQN/HEiNozWPfReVTOoF6UUGNiMBEzMH7BgcWC6pQS1bfB8x
2B81zXSKCvjLWJt7Roio4niH7QSAP8q7ZEVlwVKqEVer85Kjia+luE9y7rzdRZy+1jT0vHpdQjCn
NDowGAjybwuphvBvvILSEGVLR5cGk8/Xw4aylnYZ4OZnPDDZlRax392o1QxWzX/cwvbIzRc7UudU
1hAdnpxf1j/veNN4zdnAzo8A9ZtZY65sV7Js0/ezPEQpA3YcG029MfQc/zoFv7JNcxzKAL0fX6Pp
guPgIbjRNHpE6rAZ11iHfaxa1sxs6HcA/7qm53i82woT6OteAZiw8SGCJ4TXarg44lnjB2LMbCRa
KJQqJAvMcW2Q2S5W7kybCnbMBawDLCKDSfBGhIaJom8bMmVfsI0GWs8LwpL20/gBoZ/+87YY6shg
yHDWZjeXUszWFAtgt1fNKOEaQigUTuAkbk9tpEY1f0valUX/PJC8skH/y+vOw891Ny2I1SGwYODc
l3BZi317xNfySZxOehYy4GZUI1W0+ZSCoAA2Kr5oLx88XV8AsCngabqMu7dK1JSPVlMnD+QcVu+W
UR+m/P3FRhwPUrVQfRI/9LSL0TMEkTYZ9wuMBTVSkuNHQCru/eIgY/gAXA+xnmgTIoPMGcbaZgxp
/YHwbde1vH3A8i/WC9Cnij+VLu2WxA0ccRP0wCfDAJCN8XAUhNauF5YFm05UsFsoV6oKWW+Tn+1f
1Fk0nSegZ0HPDDgHIak45BxolXWWMnZaO1DpRqlXvgVfeR3jz7fyUMARW1KM3OSPjQwPqsi1KYgE
D6UYXpvGYJ6ku26vfFhs17EQlVSYObmmqZQS52cXIiT+X9bQcG+yBxh0kYJ6cl7lCmyFiuj6Q6cN
0ZaccojMcuUAdTsrx2WMYDE1zesEKxkKyH6JGUTzmD5pufhFYJK18il8heuPZBSBdjacvvj3jjEk
Un4D+S4DD8MqcZAaceC/3JkTS8MOUjxBkuGT1CeWL2lnnBnplgdu/mFJpyERDS/nl/uyMpKPbme1
L+uewuqX7C9YSmG9EuZRiU4XywrhIr+DfMdKislfMl2T5THGV1PZZV1EdZzgR5Q2pfwnMKS7yd2/
CJdl0egWIYcEusy+47Egqck1nGsbccrBW4ki5Ci1acqSvnBA9oG7dB9f+dFtqjZkHMRpMmt4a1qn
XYeWUpX8CxQPJM1l5MwfD7TuzibxULXAWB4LriRbSdYF2va3sHlT+q0gxxfXsH/M8hoE1kp+FQ5c
uNa2Rg7zaA/eMSxkf8oRwzT2iLVDdXgU2N15ghWjwUyyrhbI63Kg1qj3IjQzpxpnzvT+roj3lT2t
DxgxAn3Bg4OGYNnDT3sOQB0GH7LxKxDMKUxebWjW3ZkaiLX672mum+rIFSyaHhjNaTW/k8zl1iR8
mDuP4Zh3w73TI6gwm5GqU1bCv1AmL8BMYfKBtCQbyf3P9073TSHPZGS/R9XCwlfEWhm2rZUiRcJR
UvcegF4S/amnnLPaK8//wTb2Wg9K6NyRLrXsNONDS3FIlFZ+ELpK/yNWR79G5a6g/S++EANGIQu+
6PtG42ajJt6MWYqEpJu7itZMgOz1bydtmAZyWCHXhCCbXi5sYDt6tRyEHPPU9LR4lTz4NOA5nwZP
R1JXCQtR7Y5YQa4EUn5Wc0GfPryOThjZZapGe046Z07Ator7a3a0YNdaNBnXUV+sz1rofkKILOiw
M/N1TvlPpmOtgi4TBWwLf1/UvTYhGkSLYlBCTYAUzm9k+BUdNt2XECgjH8g0mlKZKdHUnjjsxRhP
rp24EwQDRA1LEKt/bb9h7K4ExL0Xz6X04I5mvGcNiwIpb7AmbnPZzcQ1tdaXgytqlkTBMRS+6g4W
7QPbEdtwthzVxEUK8LE4VUqhyA1X8zNnBE0ShzKP+klx0pU9md3s0t0pO9PXTT/hCa6XwpFh23II
3lTKWChW/sDTqNFuUuCzxtwrax5eU7XD+NJtuPGQXlT31nEHiSQEx/R+qdmy5+dy7MtEvYPRJRIe
dHVO7G8GtimeuPnK5A4SpGr4HpCEcMrbsrGSYEMIpmYp2ykLYg/FRJEsYuvKAL0lblEpo3Jvv2xm
ltpI4AvDhIxHwTGHyAjYBE5Vi6l4iXHD3vItC+Dxxh1CQno5T1BghdEsbBw6o0079q+1NJ/iWZvT
SgrQFCgYUYBvI5S3K4xnVXzdxDDfuwtYmOgNs1yRMA8xhM5sIk2lkiQmT60JvIWY0RvzXpa8qqFT
/01VnBY1fVfEdUoUoAnm51y03HW49ra2kwJZfBrgn7auMuebxG95heTsqD6+3HHHo0A9C7sAomHx
EAVKnsAFjG10Uw8cQqDltHrqkz7tutDA0h2IoQ1+lv9jL44b7w2l0Th9qFQIekzLZq8frM6CES6X
sHdBvSYcUtR1u/kVWNxDdp3UKzlnnZcyqJPUWNZTHg8Am4QDYUcIPvFCiLfmDMHygL/vy19TURDu
ryQOjpk35BHDH+PtXyXYHUmCcPN308657zjBJmCZJlyJZ39khC/e7tAMiTh4w9IOYqYnG/rZhiPD
1WcfNKxIIs8jzgi9UHTyAicf32r3YmBbGyyNPBQNmAOMUovf/d3WNJrkcHX6sDVlDEZfP/v/U4rn
bmxtATrHsaBhux2uVb0SbfF0vEUQ6+MD1VM5pKYdKTMpYmA4ZN0rsri2yKcyNcMXWYuyi9OE2rEb
8q0dnnNuRtmrNxARET+SqpFO1h2vKGNkvDNbzKL/BJUExADkBpkbovaL8w+CWaTTvdOOCX967BK6
CXa2xF+PWZK5Ejp8JkQuQ5SaNigMcDtBBU3FvoAiqBvVyfBfpUr3CXET0wHHlYJq8m3BcAC7HP91
tgjYZ3QACpQeU3RmD4RIPP0Oq6CrdIPXwAJ1w3XcX+4CyvTruWJWQLZJLEig1ra71nRdAfo8azrw
YNWJG1Q98KjNhQmJYy4ZoLrR+3w3XzWkym743yAMyvyGgoAPCoUFu7n5PDD1806oENtUofd6tpj1
DblO1FSZI0LjqQfoDktZ8BEXc77p7nl8nSPpqbeOQ0b/upqmarnKmlM7UF3QXotd5TIlwrsdcnw4
L33pp+HvL5ueyw+IJezixc91TErll33hoYKYjOFa2Jt2eHdHyCFXlOJfHD8vCKqxCQtWagP22iZE
WzpV62olSoUlOSurACpCnh8aGoafw3ugJARu06vMbSkUdt5Phtdc6I1wId4/WQVvUJ26SMdsPffK
qQtc2hTwjdUt9z5A9LgeuMoFcZdyhU/RvxLhtV2qiQf0D0hFSElzVo8cJar//bmUBMWRhwOzNicT
pl8GpQfowi3Ljx7GR+bEVy//n8kylhu+XyUXwkrPI7DMS1MRESemWt5ndjfrICLqUXythGiihF84
29MEdMZvcnFPtv/uLzIQdzBtvG8I8NzgYx5xQGVvr9ijTr5jvj9/RC19/nOLtb2bSTYzSLokKHso
/7DG+IuLVJWSSvDTF//vfFVxK0r6Umf+c0giCU+Q+COcMxU36mamNJS4+6yfRCkQTKppnEiYsE4S
MIqtYsP3ovIpwSwnSWaSlBymbubxlYF6d75U/IGxoKeXzsYwYDu3IvKDwHyVhU9fzAX0WTSPCPUr
m8vCkzD6gDWNAmSH1C2PnB16TnXrAlJlI+Ouzk14QZfBSUwD4G2ZjbmIUBiYtresPApZrdurKCYM
lVcHU9XJamT0vw+H7BLlb8L4qY5HVfa7z/Xbvcdb0sjLmZaOCCh8bO0GIXOE+jnOpGd1F5+bcko8
XBIYBG3z1FWVc1Q4L7mElHnpVIv16BqXq9oufVs4O8lGFBO73LZe+v9wt31blSas3YUQVP4JZJ6A
KgrPsDtTprKUvgVEK372h4++EqVS7OLe1GGA1rb+kpG0w04rdFB75FHoS6qKXWy/ADTPOOugG3jk
c4q4W7gaRgY+aVQsRDI71s0kbG/gK2EaXpKC8tOx9x57TkpRu6ZMsiQ/7wJ6Dm66EEO4mzR7DPqS
Xe/x/nkRxWuxLO9lW/PAqdIFsq371jfCEGdW3sAtllr4RYd2pSPyXHgT0KPx8vwsYykTFapklQ5F
dIZuAPKh6WQG0Q3jpT+btJerW6sPMVGbQDf2FvlNB6Aq1RWewUAig1T2bULE+9PB0uPYgQMzpy7v
hX9Xjt2Yu3kHr8AO2bRYELZEW9uQA3T0l3vHpATjKrw+BGx6dTPCQErqo6wn5JRFpjKbRLv6OpfO
xREepZQjXUbu37Qp/acZpzk+O4mVyzidAPYRuyI/Fe20RJmvgKFeu8Czru7Jjg81bmXepQj35S+H
D0UzlRXfOlkzhxNpSwTnNaX6jzx/hMIA8Pf0RvXIFZtvkAZtDKWDRTIwKJw1rex03bVRG8TbCjKH
QIFq0VbSHzQTmMmAWjSaVaOlD/XfYoW2IMi+IX6lqDcsJUDfeFov4GqBvi5kRHSKmS8rYlUhQqbv
GrSf1RGo1OqeybdDh9OHkkIG8SO8IK7bYFa1hW4xeaGoc3lDQNUMb6vgMtePuOoy4PTAxqvSVgNZ
Lx1vOMlSQdYB8AdDfKf7zs15RfKe6UQNEBJs0Fu6SZijrkE+9d1Gfg5ZMvZ3/Pz103Jt4o8NI49X
uVTDDfA3Em5tyEHr2Am6TXorRvtCc9d2kcHmudEkB+UiBH4NUMpqd9q9/OBsa7OfGQF+tyaZFhde
DdWE8iPB2T48Rl2Mnaj9UYDlP9OnzxtkPVAR0YnWUHC1rOhpoKnJh9HVnSoTDXwWQddW8VqHFUHk
lksUOzv58n683FGByFX/ZR1OxSxRQhzremNMZMfDVSETExqkhoNA3936LAtfpZ+EZvM/NOFLuJqx
ah9E5Zc9b/juSZPndiEiXHywK+sgJKWgCn3EWAASc2xyKRTF8GmbgIcNOvXc888Wux2ds/ST2mfR
+79jW6ZpaOAjKoCocJNbiaBiK1JPGD1JBwEx0K6kyfGQlrP7wzQa7xc1lHYvRE6FcIUVMXxMyFm0
ll88qg2Ib/P1pYhX8y+h33YVOBxaM6zMj2RDwtPcuJFmcfTQCYW38JW5X7FjuV7ofWowxqKGp8mX
i9967FylrnhztabD/pvYehDQ2y86GxnBYgFqVp9uyUEAvr/7BxvOnVRykEnwqgjUgC8YfoKhhFwu
IuzFV60gValeKnPTb0e23Msdd+bh0bP+h7X6Wty+rwVXvt6oVcVS3myxcvqkOVptHmzDUuNKXRsQ
ZGAmCltQ1EB9SYnZ42gCJeLVytdmYny5gjZfQ6UMjoTzsZU1UTPP0qpdPSJDwUnFAjn3cTaCg0WH
4K4DrxIWJzkT+mbWWGzXxGL9UCk8vJ8U6WiliahxV0AXxeFI3QsXKoo5bBVGOM7kNI11vLW0en9r
frXaBcTUpKeR9ZLIKlcVX3em1zvC4lkYHzMVqFLlKUbsqH5gP918RMHj4mmqycgkkjgkY547j1Wb
BsaBFphgou0PU9z7ghTTzmy9b/Z8A4fwn8RlAMpjqABM1HN6dKCmRVpvjkxGYeuqXgGYgxNVDP79
t9+ykxX6z1GlsR1oN6m27V/i1RECcr3OiAhZ+PrBdFRJvOw/GESkPnYYJYd8l7t2PbpHN1g7x1Ht
SspKBvD5aQehuhszKdJ7ll2kYJXdvwKLgswtrcQXP3i02xT/kD/lU3whaU0cGGpiwl0IZwcCtqCb
ubASHdEqp9q1AwiCtBbSd3KkaTcysgcynupKGGWosq/kbh5THjP8qsLi4/uEyuZJYC6UpQ2ciGqO
2NHe2u/1zvNyNKbgfNCSBp+fNQ5eEyb8zTc+/Nt1Pa0lHvLruGSKrDWC4nZ2HGEikd29GXTAEHVc
aFvLBPIx6cDGXvVbs0qvzPFmUyC/WBn9tMM1JMulV68bsiFfpRdgDLoF1bR9jEH1Sy9A4mQ/Yk3I
+j8UFkPpwXgNYEChXqOjUSzE8w/guY54h09Y9AvmEvzhte+rAjM8cpE8SKlD0w5rHz4xx2qy8cJa
75+ucNbVjcQVHI67kqZvwKDOvPHTdYmvU5eeX6nrIIPuX0REqu4iHJ7kMVUTAnKkY3MNIBBL1mRq
y+gcsyqfoS2GrVloU3zlRdcbOa1Wbh674n+342ScX2ZF6R8NZMN8geQ3s1cfcD320vryvlqHsw45
Apssm5FKbMOKHEehI5WsfWXfPoq/2M5WE2S3Wu3+GC/3SSuMbUkFWqJXjIvnwp9npmPlOxxvUiji
eGtvsULqeFPGwo5DLFd8/OmvERrF8pmv9w0NSxMQNOFVLpk9XoKgFF/AD75mjMHD9tQo6NX1OkQL
Pg6cD8xLZhLxGikczPd9i36Ls40Atp+/b3dSKLBFcgdauHmK6skQPJZAxQlSgOTbmVhg/yvvqGou
ki76NxV76NQF0URi1Ts1ISE0mg3pWJOdei66KYUVHQ04Na/OfJHnfHHx8vEebCVJr7uNEc61UX9k
rvb1hFW+a5M6LO8U6m3yUFMLEBXT6o2MC/GccuQ=
`protect end_protected
