`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 928)
`protect data_block
0USWSUGxovGsyBJteYpEoQMYe57U7EVv4KgCh0gNmqIMNeyn0NylMhbEz7Q9aPPbVwnh19A+zPnJ
GV6MX29zfY0sRtJMTgHCLe7xS5v+rr91hEwovxoqyL/IS0irnoDaJSE7SgtFSp8WdDmswgukHZC8
YW9IJaInHng/d+a1Bw6flqUyZV0BPQWUQ7EcT4B2SWJZHGarVRHN9ci1ZvBHH1kpDFsUr9Dhb1DW
TKyzCH7qCVZM+ipfkdmYhV3c75LNAaFU92jKyYuY7QhlG1QRz98If5Y4oraPSB501OLiQbjmZb9N
23ut17hitcQN2NO7wmta+fuWWCV0xodeVXOFH+wIYSOnxmqtzWAEv2vW4GK6U5nB1lojg3aeEzZh
ewWpj1Cr5on3YqO5SEE9oWXQhNDbOQ0l38MkXu+5k8PcK4H6Yjshd0CNwIb0KQISz+XzTWtkRzV0
gCKJkRs2DZW4y0QrOd9miwYSE1XWL1ymr6NAEs/uHkD6q4l7NnEIfEfVmJ1mKGevpqgk1bN3mUfC
zSUIgSvB3LFnuPbXXHzWLpNwEgxu8SQPB1VZfk5XuHvGTGjagZqtPgiXFUzldvoFut2GicCwTUQ4
cRBuWCvf9p5tSvNiE7HrtY+gmew14VBa+XdPk5nqIG0TTTHYvXnAQVvJmU4p9d0FrESWA9wKYwY7
TLkmA7/uG6EeaMLBkU2mm8yST4gfA6QyuKXbk6N8ZWGI2fvRk8w5Nik5DFjr++U91XuvJj3Mi89K
fH2hvLlDdqbpdnTQe8IFW8Rpqp7RBwYXj7jOYPs8y72irpIi/gHzR8jZhRXIymdp+4xI5rtbjMNZ
9J03B5+giFI966He8VwI+qTTIA6uk6qHzacINQPf50CklOVqCvJf7QpAsuuIcTcd+oL0JX1+4wYQ
ksI8hnHRZPbO6a8fMC+wNVXKgOI6rZI5rjL2Uf28/buMUWqS9NqGHex0V9AcvAV4EE9PdJhiSfzA
UXxftKuux/tmDL34TkznchcrpXkF5KX51OYyNc+wqBRYR123wEB6C3+M6JXffiGV/MZBXIrs9zeT
FopNf0MO0qbOh9k80Vf2xiUrZWZovXJcZtI3ESLQ+Tne7qIkYZFHybmT3EnT3evZi1laro7J9KHu
3aifGgVfiK8PbkxHYG1jG1LTlSYF561NtiPzRi5eyZffh93jbkmH93Im6KBEhLGKJRBHrvMk+lA8
anftgL4Ahnny/AbLE+JQDw==
`protect end_protected
