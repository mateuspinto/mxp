��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���UIn� ��V.��T�B0\�|��K��Sv:���g	�yw�ЪQH@��������o�gL�c���|��c�Rȹ�S�B.��
Ў�5��wv<��|[��(��<y����(wt{~vq�H"bs�	N>�rL�y?�rS͈x�v���,�؛�p�#f��߫�$�� #�'�\���8�M)s���M�-;!�8��������V�e	�����]0��n*E�(�+_��#��П��\A;�@?��ھ�7�Sg~�:M^���6�G5�9�ǡ�}ԥ:@�`:2S��� ������"�iz�~F���U
s��&EOMo��O&�i�?��k�O�� R�S�������`�;E�}���.���N|U����=��6����~�Ht��u#|�|N_:2����3��g�$�wd�
�l�!��.w�$\U�GT;y,�7a�L�1C�֧�������^f0k�A���� fc�<3�c��W�";�urCy��w-�#�+j�߼�e�&��nϘz,#���͜�b*Kj݆wX��n�V�"6o���P��R{X# �-�߇R��땊������JoՀ��6��yY_:5�ƀ� 1#�֯c-5^���x�	�yBZ- NpE�k	z� ۜ�̌��]S�k�b�}��J���f�m	��7J�N�qޫ7�B�`��������xv�;i��H>�K6�+#S~�]��K��*]� �e�e�}��J[;>�-��PS��Ђ�5N����+&��iL�]7�lΠ���}~�����*�&�J�iR
XZ�9A04�j���% V����ᅱ���1��Exא��#�Ӯɧ,@���*������ꅁV�w��M����趾��R[����n>�[S�@	�af�"�n��AE�kJ<nVlzx�)����#��j�<��i��6<Y5�5G���j�ғg��#���N�)�rO�s��v��ޠ���)@I�?���ؠ|���#��t���XF�H�43���O�?���ǒ���pP]-kM���i���3��%�p�ԛ
�����R#�7�̡���&��|�2�P��7�'�v6T@:�Έ~ݢ�����o�`f�qOWB��)Wɝ���g!}%4,ќe�x�F�؍]+I;��tR��|.�fӅO4��"J�S|}��*,:/g�vU�t2b}j�d��=V�o�N)�Q�Qw��B:u��cv���3N�E��>"��2g��A����M�R<���ރfK7Zw�,,��;Z����e��l*��ʛ>�.�^j�����;��`��h�ȵO|u����(=�17�-hP�>��6ݓ� �)M�jL�IT+��Ώ�ɁJR5<�C
gR ���ǻ��-t��{,����א>N1s�s��2���$0��a�f�S��B��S\��xM?�H����͆�����n�ê� b�k��,�	V[�/ �8?�0���R"u�5�����<��Fc4�_� j�^y���L�(�쬤�j�Z��d�͉zC�]<3���*V�K�_���G���fs)�����"A�&�U�7�=حN��RJ�c�f�T�0��fY;6����� E�\_kn?@���j�]3 U�,0���Nr�o9&B�`����v�m�)����q}��6�C>� �	Sp� ����@�&KV`vэ�����nb��b	�!z�b]�GX�oV���y������P�G�z�&$�K�/ډ���*�dNhzM��7���zh�(�ų��aE�Ca w̖���5֊�)BJ:T�<=ϐ�`F��w_0�W�DE�%P`��z�U�'�b�c���L�v���5�tٛr����8��!�{����s�cv
���ȼehgDaN�y����?W	�ލ�(����Q��Tؖ���I����X���--H����O�Ѫ7)��X�"Ѣ�kh_qt�U�Η�"��a,6E��,}!�E�R���fΘ����fC�Ѫ#�-���?=�iʛ�2;*,�����`x0-613���(w��ԛ�*���[0����� t�p��x�ao��S�r���0@�X����� [£��=�i���s�`=��9��Ǡ�Kɝ���'��H��m�������|�
��xl"B�7g69O�n�x��6�zX���q<oU�tq�zɘ/됴�Е`�d@��H�.��&��;*6e(K�ˣ���ڦ��ń`z��r�ɰ /X�E�e�;���B��Z�F����"�Y�eΖ']���%�� L+h��`sA�7J�]��m>�N;d��<���1r�jGd\	@~�j/��X�D�C>���M��'�^\�p�IX��l�;`�:M��ß��0���B{wEd�橅�������Q-�ay���{ĸ[�driou�����?�H�T��JRq�S�3�9=��]��F*�ѡ�A�AY��U��w�	8��*��������<K�f�
m�S;��ߓ���P�����Ԡ�]'N�n�Og���M1T�i$���o�$/&itH0�!Rj#�Єh��՚�יh~gW�M�2ْ�7��nR w�!b��(�rM�ބE�ꈡxdr6 �x��I-��R'ඐ@��v�W˔���l��lv֔�- g?�hU�7���Y|w�	g����r�4?��@�x�a����cgqz���a�%�O�y ��(K�[��#�d)x{La4��Li�8��3V`�������z9�V{"w�rQ�`o��hYQ��g�͖X8���W<�l���MMɹ*����K3��O�0ӄY�q!5J}����#�ω��=��c� �g��OI�n�D����sli��/V��<����=����~���{���^��Ͽ�z���fq:��t`.x��ԙm��PY���oc
��o$��j�(#� ���r(�E%	�y�8���R�g�;g� 6�ḍN%�_{��Ĵ��8cm��~>Q��-S���������{J�!g���(E������Ñ<z�M}��D�}��hD��O�=��C@,��*d��(v���k!4�Q=ܷ������Gsr.����'&�/�G�d:�)r�E���'rR_����,�����g4Fǿɝ����1K�_�
�F��kiyd�7l����ص��x,����d^��'�u���3��M�>uTzQ�5~��h����s�ݏ�r�m^�!��IB���5�Ɩ����A��vg�<~VT?�7���pKB��_�[�!´N�>6/��Hw-��~��Z����0�15�L/�Bs�V�]�0�I������m�����6�*���^��d�ñ�m�.PO}�_��٠Ͼ�AR��%z�G�M3�R�#�<�&��;�n�%���VW��%L$9FenEG8�i3�)���a��6��m|�"�ow%��<\�1u3���S��U�7����x0E
#O~/��-AN�iK��-ӳѩ�K�`Jp�k{���}��汥����F��	;�~�uQ��p��:5	���5��(ɍ()���7�O�0j���s��]�d8�qC^.��ɯ�����Kf3Q�����-�1��O<t����*+y�C\���h$���7�d�c�P���f���zP�$IN�8/����
�k�i�q���a^�b�����k�%^���*e��G4�I�j��v&�W��/õ�pTr��y� ���j8�_�;�H����;���kѢ����������]f��
�n;�����7z(��ϕ������2谵����͙�5���P�Hے����hH�]qV�q{,���$O����Ӻ�s�r�J���S�d����˼y�~�����2�1Rs@�0��0�(K�0�+z:*���Μ��g�0{#�NV�b(�Ua&BD�����5~�ve����C�I��)��Ǚ�|s\ʺ���4j쁡�e�u�k����6g�He'����Q�αE����[ɇ �ؕ�!=�X�>>�-у�lҚ����ʀ�@X%��_�s�m�~�s���ᲇ�	�?Tgh�CH�r���E@�L����c$�-�<�;Պ.eq1_���f��-�r��RN)��C#��H���(D9u� X�v��_���*�Ϩp����㛧\e&��=�2D�����{�M�L�E�V�V�υ��[����&9|7Ъ�݁��tµ�Z���_����OD���p,�3h%�w�8�{ʉM���%��R�G8���t�T�wX?Nv:V�|)p��*�zrjj�NhJ}oÉ�������K�@]��p4��$Y�3�7�q��W���@yC`}5 dn���3���B{J�(�b	:S�
�˸�X�ig4�.�e���>0yV��d���V�fK�<����?��p ���K��$1aHf�h��H9s_�q+���P)�Bq���D��V;׽�d�?���Yfv5A�Nu�����Q&���gs4Y��[X1 �sfLL�K�$�4R�����3>U,Ȅ���IzYC��A�O�</��KQ8�!kO	��k�BO�ux,]�k�{Mn�}Q���`C@O��9��� S*b�b{i\-��Z�B��x��ryc�I�-:*��G��ǐ�GU�?>|��_�i CĂ6��w�U�!J����%4eiR��@�$�v���eb�Bn�VP���#�GP�ϕ�R�/�	9��U�)�7��o���N�p�{36�A�� ��g��ZȊgt�];_��Vw�$ƅ�#��w��s�^*�/r'�^��$��btYR���8~�$���r9��u�y#Ө�΂��4S�8~�7D��$BL��I|�M�peB+����Xڌ�k���8���x����,�����P���v�����m	Z( ��c_i�jcjD���g�V#P?8)v�\���T��@в�� �����Y��z/�nق�u��M1�4�w�zi�O�
h�Q�Mu���;6�s�Q�_R'e&��T#�8_z?Ɣ��"G+�s�
���g�w���0=w��$��4j�Th����N�����d^ag~����j�1'��7�(���/��(���.���
��*��I}ɯN$B�t�qP/�E(9H�F��H��	O�Y���������e.6��m���p�l����cs�ky�*��8�pd ߉�R��h�o2�N�<���e�!�M�7	��ݼ|���Z���S�ε��m�ٷr����%�����t�� 7��ۜj��u����Z�(�m�J<�jB5	xH�ڵ�h�"��s~�.�8U<�5YX������kDLW��x(�S"�E��s�b�B��b��A�]�\o:����S��F>i��S��/�+�a���� ��ق��3�],������wu��V������?ðX�p����t��[���Z��4�)in��������g�N�@g�P�P�r>m��h�t��rJ���F�����=���(��5ZQ�wy�����ݡ�G�M���J�+?��H�-�0ť��F��J ��N�,���CA�9V�To�|�jVo#9�o"��9��rvP	�G��pYQzv&M�����R�)�R�������t�9���0M�Y����k���h#>ۨ̓���ݴ�sl�B�*O�b�U���6|�<=l�t��	��N�?��,� �!����w4�C���t��C�E!z�AC��Y*�¨ŖU�V����WwФ��Q����Q�\��!����ߌi(�������Q��,Aj�Y�t�'龯�����4���LQ�T<�H�<:[=w@�*���t��I���1�NGun{�u+6�����jq��ŷ�ـ���2��	]i-瘕D�L����a�Y�����RC�����8�w2�V�fI�3���k���:�wH���Ok�6[_�̴g9�u�w��@^c���d�f�������d��G�����,E�ᴁ=�ͧ��,�'L4���kM|u.�N�0=<��$�}W:�`���_��\��AF��'��~5�N�s^�P�����C��%�N��	éC�*j�J\>C�~��΋��K>�N!"��?:�G�x|ٰn���A���J_i�%���I�/�s�x�.l��$��~#�΁R�սt�Y=�M�fX솃I��H��
��8��݇j'�7 ���b��<���Z���s� ��aS��&��z�=�(�8�Z'��&�>������"3�PG+�h�1�:��|�P�(ʼ�,g���6���a�Q�MQB����T�3ٷ'"E�7Bx+�����5�~��'D6�7�	9�ޟ�Ig6�P��˷�+�������>�Rj��QB�)���o��P>Q(t{=ۑ)����e�̞�T�BYc�j�K���}>عRzS����b)Y������}�~fg�@�_y�&���)o�q,J�筤���Ӝ�CN;rX�8p��9LؘK 2����J}��~���TԼ���}s�IG�l{� f���J�C��`v�
=M��^I
�>E���ꢑ �Ю����Mw�\�|�8���{�oJ#���|뜗� �;��e �b�_��N'I��h��0��V�z��}M��l�����sSf~�˖I���{S�c�F!s��RfH��)^��q�b�������<�I�J
����g3ӈ��&>�n=��Y�>��3��C���_�k�j,�]8`j�����i'��H;�� ���R���ܜ6�hE�T�� #>��;
�2I\/pj�K��8N)3l�0�Yƴ���
���T슌�p!����%>�L�T!��A���A�4f_1��ʉ��r�J�%=sz�Y)���_��&.3C� >s��($Pj��c�~�0��WSb��������,���8w7�����M�ޡ?m��(�G r�9��:�i�((�Q��=74�O ɗ�Z;M�� R�e-�'͐��
����M�A��E��Y��
bM��A�z��0��f2Ҹ�(�6�L���v+л;��avQ�)�mme�}�A�w�6 hθ�����f�戶��¡\B� _7���WdU���ybQ��G
 ��{=�ÀVJIp��삋�TO �#R<�{N�ĐSn(%l�TE��	;��i��x�azɎ}C{���S!e�'�ӎK�sQ��-|�~���Y��`��RT`Vtk*E��'� K������x�CXHD�`B��\�*��+& u_'���09)~�c��H��I��V��T �����k����섛���M賶����h�R���U+4r<:� m��e�]���7�fS胡y�%�F 8x��ѽ��֌Β�S���&xh��'@�u��*DN7�?J+a��j�i��ю<��Z��FȬ3��׿���;�?%�&^���bW��� fZ^ヮ�<a�",�*]L�xg���3��0�2�2�Y
����
���*Qm�󪈏p)�lt�X߫6˯Q��g'����������i,�^����+������.GNU���K�!�'�K�y�>�C8��⑤�d���aG���QRQ%��*�jt������.�ƿ�bNm�џZ�H�������2�J�ĝ�;���?��Y��|h3�:��XF��v�����l{�J2�'����u����S\2�@�[�P�7�Ϫ�>��$4P��z:���\4��q��H��'A�4B��i#bx��w�]D��P�t����b�5*��W���ò��8xI�k����M1EV��F1S<���I�
Y&����L��U��ﭓ�d��1�m4O���˜�:{���L���:�bM�O��ͳ��L��b��(�O����@Y�Ŝ�-���7e �Rh)b5��	�[�,�/h�+�C��V�m�3:`gY�L��Vi��^О�L�������D��o��q(9�v�ճ��zz�A(Ȉ�ې�5s��!�� �Z�^����!��w���a��3؆�1�M]P�s�H���n����D�\�XI!B��yᖙ��_K�����G�+U�:�2{�TK�4�6��d�<�͊E�����ĭ�����.�Ӂ�R=p���)i�����G ��P�"�NWs%���p?/=8�Fs�|�aKŇM�$�[����J����t����4�˸PG�L|3j)�׭:9ͣR�������W������4D�)�CZ�~߇�t�%��Y�wk��]LP�ǉ���c ���?�Bu�H��|7�f��ͪ��m#N���8�</%�E�f�&��3�����|�h	gT�=�&C��Fk��;XH�O��$�O�5�T��	�зbkr�).������R!c���I�V�|wC��e�:�����L(4�};���q������H����-S��leZ�mA���5� ދ��.' ^��	�2��g]�W.��铒%�eB�▘���~���q�#L��n���4�f�K���ž�����A<F��b=��Mg�ڝ�T��ud�^��G�V�W�N���>�~�_&�_c�n�a�(��7ndx�rux����LZ�O�Xx�(�t�q׬9@�>����-rXl��k��x�S�ʹ�DdK%��蛙x/@�`��}���h�$���,J�}�NbJis8�U���J��%��b��J���]�es��ˇ8gw������;Ǝ���G�n��&Sv]�k��ycՆ�q�Q��-�n|���&U���*� O�س�Ќ�w���c=�u�Y���1W���ZBk�c-����6�j(2�5�/��63���D�={0>MT�B�|cu��5��P�vUk�91&�cԂMS4�L�{U�3^��(0W1���f�p����)�߁�~�v� t'��+hlp�ܢYd�G�M6����v�L�x�;���Y���-y���G��#���z�!ߚ�?���ˡ��KCz���<DP"�r��6���������,�]"nDf�}�TY͞M	{)r���c��3��rE���nB���{WI̻�{CS�A,����kV�E<JB!%�9�g�Q���{t#w��6#��w S�'�Zt�ߠ�e��Eb��~��U��[dB�t��̹Pu�֝�Գ8��/�>�Ni��
y��.G�ZP&-���g���U��?�s�|^h�<Qs�c�d�m���z;�x�?��h��0( ��E�� t����?4�(o�W�m���M��IN��+��v�|����D�Y-=�Cڠ���i��g.�
ҟ��^
��_A�)M�X���LB�����ߜ���g��J��$�O���a��j�Z�m��3O|Ic�vŕ�`q	{��T�O�B�:m�OJ�`����2ؽf�C�AŨ����[�[�ڂ�s�>
�ؔeK���/(���n@~�LD3.B��6w!��O35L�dU}�B[bg��i#�9NĆj�0=A���ĭ��W'�L}������? ���x)�g4<iz��&����}���˿���d0E����xm��Y�c����ПqXph��m�*Z%��p��s~����B[�Mh~D�b������N�Vb�Y�B�I�X@��%�T'��u6?w�K�Ymp��#��ڠM�ӯ���D��Uv�ٙ���q�ėU�cIa���&P�Țiz�~�U�|�|�I���!5���f���`�2fM�B��/��b�l��D�6�3}���Y�W��x�t�d�cs5$yDo�FB;����ӆ7�-��e��K��)���nd���{��v�/y�pt��cmf�,�r�Ԏ��M`<� �Spfd=Zz���u��{�Z=�,��K�nm_(@AGI��&?Fx��Tg��B�:�����e��k���3���{'W�
���$��RUڲ��Ǡ�	f��D�v��Q�r-��#b�Uv�yyŚ�R�D'��&�H-!����s��%��YJ��4_#Ŋ�b�x�C��J@���6�z:6����)xb����"�y�kQ��2�����œ�w�;
C֎�1�&�V�!�|< w�YOx�I��)G R2=�����m��8}Ji�x����xN�1��f}Yώ*��`��K"<�"�ͬ���Hk-���̷�j淸��Ө�bk�;�K�l�������+n7���WG��<T*e��'�H��_���>C�~��%�s�TX�t�E 4���j���eqbv�I�-�I�p���G���_y�.���%�/�������`�Ge=B3ͽ�9V��'
[�HQrkq�
��OE��!�*�챥w̘U.�LE��͕��7�D[M��r{����f�/1�$p�mA�ޙ�N�6����>qD� dU%�{�5�Ҟ�eG��/T.	i�fH���i�څ%u�!�;�XPՉ
n�uł'b�.KC�G_�[A�Ӳz���^�|A��F������Q��Xp5�d�/�r9�aG!�T��!7�ǰ��_'�8���*IZ
קġ'��\I�LI�6 :w���9,��B�| �&3�MO&��~�i0�D��J��e�h?<��w=��ls����`i7���|?�bg6��Z��g��8^=g��>V��(�<�'���/c�,�7!�`b������xy�)x��kې�@���
����I�����5I_�t�2�)���h;m���?�S�!լP�u'o�9a��D���!�t�)���o��d�{+BC�~����-��gH��S�g5eD��>	�3��{�T �q)�ЁɃ�O*�DV���I�,�ݞ�u�04�9:�uO���g[,��4���y�D.����z'.2�1}�AAV\�alk��
�������I����=n=Di��ֶ}���nٲ�(ϣ�E�;�=���^�W�{��폗����x��S���EF��Vc�w�`�w��m]��?gp���$|����1�C�5�>�!�����f� �^��� �e�ⲧ�+��6����P�t��J,U�1�<�~̞���Q� U����a	����+\�e;{9\��^�gI0,��]��0]y�,d�d�sZ�����j*��pƽ2��L.���]��kf�7'�}���ʵ=�8s8M��2+��8��÷�09��t�-5�Z�@��:�ź$c� �r2�z��6/�v��'�9����%94J��g4좫�:/��?��V�Ya�9X�]h�m�7I� ZA��lqG}x����Px[�\�W��yb8�����:�+(�߀�T��{9b��'�S�[IL;_sg`$w���d����6ٻ��B�����:�Y[O�}�I>Ϭ>M��{��N���yM��)wE��E���>���eȷu�Q͹+B����E������G2�L�﯉V��f��/�hv9��*�t�w�f�^��[|j�Z"�N���x4�����1��$���.��E�s\"	�l�:�9�l��Ik��bW��=�e�0��ә0mHBe_�@�}�\K��3Z�=>�oz�~8p��~N�|N���0��B ��{�J"b�`�h��gY�}�����(�S�\�ːpW�7�j��:4"@(���X�G��Nt�MB�6>H7�-�<�Qô�negϼt��	�����ߩ*��7Y���;ȑ*?Q�ǲ��:��0ƞY�����/!+o&����+�ی�}�]1�k��c~��Rj*���:����fj}��C��S�=�7V���y��]�@?��B����P}���.����'Af^�wy33�����@E�w'<��'�Uuy�Atz�����s����h6?�)&e`�w�ڱ��/��ZMM�{���׸]��ۖ�M�E��x��1�~�d4}^��X��NǏ������XÒ��0��y�'���C�Pu/�Wg��(�<��f�+���H���&QץN����q9�4�-�� qq�b`W��7�d=��SznrNۓ?��4�]ɽF��Pu��g/�H����@�=�#�����t��S����C��
��bP:҉��sȜ^����,u���NA�?Z�<`qX�kq������W!~P��lwͭ�s��V�1�C}��:���Ю�S�歪�4z�rEb�~�e%��D�]����Az�vO��D�HX����a�E���
u�(�9i�ޤ�!:�oc�Qv�6�(�M��g��=a�����z���	zW����|Mם,	1˷ay����i�h�M�7!�Km�#�Ҭ.a�
��;�u�F��Q�@�\� ��;p��U�ˈOKt�r���,a8�%��7l�<��Y9u'�'�٘�/�3�+���גs�v�p�;����� �tD+�H�V�F�ﭦ���Ϛ
ջz�~�:ҁ���R���_1�3�	��M�=T����oQ�-�"=�C�Pe�#��Sl�z���nhVE!����&�YFYXZ����= J�_qb�#+��+N���^�Rf�2�jb�	@�\�Yo�F�GX2��R�5����Ά�$�M�3d�4?�i��:Av��b9��/$���z+U��J��
�&�_�%j�a٦�KЁ��;�Fj�tNm.�
��VRqyc63�nB�>箱@Y��!hEh�qz���$_�ӧ�cUQ�:��ZM�T�)o_�N����eNδC���U��d���>�5�-�'�ũwTj��ni{��m���٢�b�u��@��p�B~C�g�9+@��#��A�(	�0 �鄽��{�[j'Z�qR�Ƨ�Bpmx�tc︡U��`%���G�mSAuB�$�C���*1�G[y������a��6@�ƍ�^��. �*Z�<5��FW��MX7��6��E�ͩ4��#��"/w�I��e-L��U@���8/Y�;�	u��� ���|%k:i�
�Ȧ�d�nqg�Bn]��K��.{��'���xEKo����g{�},�z��WZ	w�!�Tq���k��#�]�����_��O.;j
�̌�t��z^pzd$J�_���UV��^������cL�b�9:��?' ��>A��
Ye�_s�T\�t�q����o��� �ŰM���' N�jF��V��ci�z�r�A�����x��Mm�:�¾�fц#�����bf��,v����=���$�pkek��,��Q�zow�o�L �wL�A���%�`1E�+y:Zk�Y	��=�z5*jk�
0����������1Px#�s�_ �����龌��B��T��G���7 ��r��ǰ���9U"�V9��F3�u�z����~��D�s��PS6N�s����O;Գ��sj,Y�3��Ĉ8���a�6�Ώ��b6'n��5��H��S��	��T��t`g%RL3_�^1��&_ɡ�">�jm*���ζ<.�OB*���K��.�>б��OY�R�)�U����Q|��T��l���|Q��u����X�:� h����-4�@�"��(ފ �'㠶QR��@���&0w��;%�d�}ow��ʯ��m!(�o�:E~b��-*B4l��{�ڡ;l���L0�#V�=� �%�k�޶.��%���z�i����@i�y�t��[3��3�-��>��G{�,茀Fx-�]Pn
��F��}�O�YhKu,KQ�j@:�3�@��1������x��3��[ࢍ�C�	������g��rv.t(u��3l�(tp�w���K�g��w<]�%?�#����ie��{ey�Z��ߵ�0��Pz���釴eE��j �z��];b���E�ZG��/��9��?\�'К�~�R���T�+A_+ZgZEn��S����S&�f�km ��ǥX��Ъ�rB�u䙽�I�>e��HZ�_��Z޻��Ђ�t�X���!_^��{(r��8����Zg���[� 9��+�ۘ���������ܵ�=��{����h!sx�Ϩ&�n�NA�b�̋�F~Q���o=����>���˄%�jGs�q6.�����f�>�Tö��Wy��D�U��Gy;@XO#���8�qw�7��oQ�pngb1H�'��2�g����zd�A,I��J� jW���7D��3�5��{O+�X8�|�H��Hsp���j���ʁ�6B���;|����ae0���&�m�E�>��^�d�Hr���s��W�2w�}���\]\�����p��ER�s��t��)K�1D�_6�����ճ���q:�	Q��_.�����M6�D/Ȭ�/iDV�o#o8� rG��Nm�Nl����{W��_t��m�˒��[U'��w��_PS��5�?�`�r�_;�|GL �e;\~�(��ǳ�����'��׍)�g�LYt9�i�@���a�`H�?�)#��э���#��d����;oj�lܱ&�P#�K�za̍{8��2�P�˂�8�͈q�����C ���S�Y	.Z5�Bl ��D�:<ĺ"�Pڹ rm�4u���q.71�o���o`1U���5���<�,�2�� ���� �Tu(�tw�5Q��C�����Jӓ �=~Ϛ"���7������)�+�#�)�����=)l��v��iv�df @�t\���0�uv�W>hծZf���P;�>����h�o��yU-�R��_Bŗ�6i�!Ͻ��-��N'�:���sP�
� �t�d�tB{�Q$c{G�Te� ��|�
�K]��+h~;��r	;}��!%w3��	x�1R��En�t�=��ZD��d��t���(<4�y��dŨ"��C��t(#��_�A��8��i^%͡ЍUx�9��YEe�X�&�G_����+�4vv�=%����Y�������:�O�7�B��e��U���/h(K�fnqhR8�Q��qy��P8�@��STS��={��c=��2흒h���E��b��*���(�� @�m��u88���Px���u0�VHG$%��L��Ш�mlU��Y����:�����N �<`�)c��5g�R:��/$u��{�Y��Q�ݠ�q��*%�mC����o:Nd1�e�P�����H#��G�&"�S�a�e�Dw��sl)�N��M���j�b�c��\ne_�E�` ~u�zk���c�n%6"�.��(��G̞�Be���P"�3�!ǜ��?�tȥ���W"LJo}�al#��ӆ*d����U��8�S���ڷEm�_�I�������6p��Ľ=J0H�����ƗC��(�E1�Z<������`G��j��l'��H�=8��o��g�D�0�>�μ�����z
������m�e�-�����}�?2��YW�S��@�d�-�Խ�՜[	������'�4��~&'5�Y��ժA���u]{ ����¦�j�a��ZD�y[@���+>"|�VA�יi��&��:]�aN�\8B�vd7���L��p� Tm5n)��5�o��>��K�PDW 4v�]�.�=��̒R ���Ѿ]8�H`I!�}��0�>h.� o�1��Y$CU�
��s�����X�RE��$^hrF.=ztT��vݪA�]�
��i����)�1,��j}�=�p��{�$-h��c=���T�o8} ?dM���-K���ǀ	�+�{"#�UX���I�����#��h�G_�y��/���+�Q��Ҙ�=�[�����C��6�
����࿹{����Y���D�M9�wM[O���o�N����qID������?�󐿾w�<T�%��qg*&��mѳ=�����&-�N�������O��(�D�K%|Bd�(�����ڻ���YLyA�`�s�9)������މ�k,���/g��%�.`'Q���6��sW�;�_�^{�=|�/b�,���+0�ͅ+�{�YW[W�h�����FAa�_�`������
IϿ��x���1A�V*�!�z���uAP�����I�6
W�1��'���FɱTQ5Ӿ;t��X�"��e%���/�:�*�;���Z��Lһ�Ӷ����f���)b�C�YZk�Ʈs"��_<��&j86���,cLg�Nt������^>��E�%]�"���P�I�p��֠��37\6�bD��1�U]���z0╱�;{d����L_�6_�o�8Ch� _����
8�� ��`o[����{��єv����b��V�!�`B�z�ډ���KC�����;��`c�Ww��KԦ��u��|Z%�i�	�\�
�D[ͺ,-�UL��̆���� ?��B(L��C5�l74г�S�wc����\^1W�̜-�e�/�X `��i!f��1^JY�?��O�!���Z�Ze�FV�_�pƁ�]L�"�/��ES�HW�A+f��a�q���0�*�;Q��rP�B��b�ET�hIj;_CK/�"��=��4qA�d�L�ܺ�s��>�YF���o��	˰���ă�&�Ԓ^nN�2�zr�+yH��t��j-�hrٳ�21%P͔�b�f���9�z��7F���4��r�eQ�n?'�G-@�Vb�Ϻ
"Q��)$���� -�/h��U^���)�_���h��qד�Fq���J�s��Q���\kr��t�]`E�W� ������I��=znh,%0,6P�|A���Z��	��6kiCM���/�W��Ɯ���4�݊]��\�tM���o�:�aP�g�bKC�LrS�,��&��_RJo]��GT�x=&��w���Z�qb��v�����p�������~J��$�.�����xu�ɇ����:�<�[1�]��S�M\�L-MD��^�"gN��D��b����a곴��w��|1m�rKx���jk,��xх�s<�as��q�Hi����>8&�����Ҽ�7QJv�7D�J�4L��N�|��"��<:߻��Z��C/���0�SƗ��ɴ���
>�\@ө��%�a��ژy%�N��P\X�]{H��(�K՜d�$�r
ں$���	Ԇ�>fٴ�a��~������e�Ŵ�`�Ҟ��ͻ�����i{�u�`�n�ì����c��|ܛ����?,+��K�
6�ӡ�oTdt���z�m�Z�	�����H��n% \&��l��<hd�<�^�S�d9�chj�_r�˓߱9[rf�j�U������J ]=M���Zmpc�
+�F�V>���^�8�8'[,�BU)�G��E��.SlL�#rQA�\��E��wO#�M�] �ŭ�o�e�Sg��U<�(�K�����eC�1W��]POe��*��Xy�4y�,�|�`ȶ�7|(C�z�:���z�a�
;��< 
%m�9i��f���{��4��_gr]�(���z��h�_�h�Q���Ym�n_��y�s�^���7j%�y{L���mH��w��A�����I��ߴ��RU�W�ur�b�o|��Rl"7^N�+�Jm'u�{j��gT5�K�-[lC��U�=>��O�dǨyQ����v��l�׸�:ب0���e�D�6�+٧�����s	��=#��}�P��=����j--g��S��,�A�{R����l
U 1Fl��C�F�ͱ���� �G�p��G��{�p )2��lÍ�y�ř�uPr����D����Mlt*��E0�wN;>�T���k�=�_zD�n�e���eyxich���-��r�6���WP�
a0� %��6��?"�t�3F,F�{:���ԶG!J\ ɘ̺� m$'��ԯ�OQVe�n^s��j[��(�2g}���:����C{�`/�G��+zL���!�ț.H�/���1z��-RC���4��4�Ģ���%z��{Ɲu�r�.+�8o=ɿ���.�4-�D)�A�u����̬1b��7EĜ�nt���-��?�7P�8XlM��N��U���w�S�@2^��w����H�����+���;���)�����Ck
��6�,~��14�*JVށ3쐯Hŀ!zF8l��Xu�͇*����,gZ9��L�q��c��IUr>��9&��n���mM�7��z���)I�U��&sT� ����Q9�� �H�(i&_��o�R'g+1���>��п�.-����V�K:��V�����i��V��*��=ytH�=��K4�~&I��x4�w͓��	@����А#�lGj�@�eEPS�{ǀꁱ��2�G/�����qf�(����jy3��< �}Ҡr��:�!���
�����GN�}\��`6w�c����ۈ �N�T�]:�$.0k܊L�$��!��-�S�̽,,5��r_�9���xvʨ���W�5[ZB�� ����S�(�/�u��d�X�>J��d�Χ)�tE�&����E�f�!H�:�5����w )���1�d悴���O�;5�����jg;��+�̞��*i����A3�)�aN��>Ց��&6]���.�D�IBA����߻*�ڬNJ �<^�<y/�r}&@��w�����0��M}�w�$b�zl�0]������Ծ۽�ף�!4]^�g ��zߝQ�w6������*�?���ta�H�}�tw�A_.<��9'����H�cW�xx�g+F�h�6w�ی�>�m�Q��h��JA����kD���1��>�WC]�_W��`S�Q���L�:�9���� nB���Xp%�eڤE�I�ԭ|$o%7�`���|��]׬��Ґ�"q�A��G�p�q��PwDh���l�B ~8V�'����Ԏ�g}Ye��ꇚ�i¢,i7�b�),����df8U�=�p�J��r��_������ΔJ���-�=��:���z�tm�G��瞬�'�e��s��R�����|<F�b��NeA��KK�G��iL��>�{�}u�Yd�K��M�[)��a�Z�^^.Y��a����J�zU���ˈ�@S���@r77P�@�M��0IJ���.|4��o�~���!�L��p}->E g5��R�³�����$~^'���̤wG����˒&�t��O��@�F��}�A��^?rE��?Y�C�G�?f̏�Т0by��E��������r���&��$��3M�j��l?ϙ��=��QՁ�ޏ%u�	n����gS;���s��V*pɆ�C�O�&eʷ��4O$�;uh�r39�G6�|W���Gb�ܼ�Y�/��ŵ��L�H>r�U\��q�\���6���:�	[z�6�p�_�D��U���*L�sl�z��dT�j�(���z�u9m����#v�9ˢ�V�QJ�����MC���

<Z�N��͘�2XK�Hr_	 %(&��ܦ�F �E�Cc;����rA�s��$M��u��2F��[T�o��:f���/�����})�˗���z��#�|��]�I��4 ��}X]�j���:�T���T.o�>�D�*��\�K��QX�Vl�V:�������pd������z�e��[��޲�����n�Km,�CilDto��a��K#y|�[;���Wp�غ��`]W%�m)Wh�9�����D��<�aӊ��?3��3T���"��h|S-،fsxi'=PB�;�t�B�| +-l\�D��guS:oc�V�RCe�
�Iq����+R�e��a�$��R�N�(4�Y�#?}�-�=�b�������M ���VQ�$�L��^�[��t\Jn���/Ϟ���8�I7��۩o�Q��욌[2f�<�'-�;�e�15�R��$K�U`Q����$����Q��/���_�.`�Y˾�q(;y�I��>[�ڶ���L��Hk�_�
77�:<��;��ѻl���1���	U�ݡ��՝�ّ�4Xa�.ꝲD֜
4wm+g�|) ���i�V�]��e<��Mr�R?6@^�~��R�*�_[W�E'���{7v�;҇�|NV,�M�e�.�&W�Yc�Ƣ�^_��iE�&~�l���Ĥ��m��߃���oHp Dd�(O*�]B^/�=��������'ܠB��'2�>=,�����g���a�h�������1_�Z��
���	4{p�?D\�>����5_���P���	�OV܋r����s,p�S�d����3�Νi��~�n�C�g���po-�,��-<�r�)�F����	�I<��ԟa2d�qu8�~,�>�f����\��J����p�1�.�2l��� ������e�ڀ�~���/a�a�pKꁌ&~��W�+5����M �1��/gƽ�y��	bfC�F<��Bc���+.�O=�6�w�T�P��v/�b����U-ܛ�ˈ� �:��+�CB�������H�7��f)�F�c/�ܴ��+8���y�Y�?��cB�VA$�C�&<ݍZJ��!8	Ni�0?Z�E�;l���1ԕO���"�G���؉�q���M�������S�K��$c�Qg&ϑ�D�&j���KԞ'%���7I�"�g��G+��	v�j���xqLK ������j�V���y��j�u/� 0��ʈ�yZ[ò׶��
<5�W���WP��n.j�2+��:��/�JU�C�*%����@2�7vT��h3iQfh��I� ������
�e�����'�2�b�)���9_�F���D�º��5�LAt�8^�)��2zR��y� , ��$��:Q�*K�%��#�^���{��<?(�K�s�\!]�L+�����;��h�7�:&j����/��Geeҳ~s^�kP+���ըW=rp��f"k�b�3#�J�?#��<�R�6��ȷ�%����Lx�j�h���X	я͐���R�T�|�a��#Q�y#up��Ȋ&�3nK.���l���7d%٤o�/dh:�^6�t��ȼ���:�~9)c�o�W#u*��GFC����*Z�<�ƁP��$Yl{�$���q�g��ײӭ0W9G5�1�o���R��	�RcPJ	�]!Krv-��Dݚ��6׳gpZ�-�rʚ�	�y0�S;������6i�{�lx��8ۘ	���	ER�j�Q�X>���14��I�i��DQ<W~�Ԏ�<���,�T�q��60Hkk���}�"����.)��m��������>>2-lT�D>P��������C\�:�*�˧3_b^�r���D#fW)�u�����x�u�\�<>c��%Y�Y�Y�;+@�vU�����f��R��F��k�,�(�4M���4�M9/�ٙw\,ԍP4 ���oOj�<���!��9�4x0�"V�N1t�?Z�4�g[d��n`�U�&�4ǅ0��K�Ǒa�Y@w�,���9��(e���k����� zU�BF��u��
�骞Ծ���1uh���ޣ���PAhN`���*�т��q���2>���e�p�x��N|��(���L���|U�*���-�G����B��`~���G�%~9(�A������
�~���~Mc�*�N��N:6����//�ʎ�y<g#����3�Ǯ�]Wv��Yex���0�d5ę�.��K�X1D9r	�s�*���LC��lO8��&�vε���z�^Df٥2�m��t^|z���\����ŋ��a�m��ABe���]I^�+@�ڱv�u��3�Rv��+�r4�%�X��N���<.��s��z{��n�M��kd}�-]�辽P�e`�;LCR�~��-D}���@�k�]�ZH�&(n=#}�K��(}�:���[�f�M���ց��	��F��BZ�]Ӷ�N�i<L�=�؂�\��o��Հ�]�I5I!��p`ح��os]�i�q��($�u\ݯ�kX��~7R�V��	���,#����� j~�!!Ox�#А6��\Șt�q.)�����4��LxQ��3�O���e��dtK�SO(��.�b�Z�������_�Ei�8��3�@=���,�=�&�$8C{����a�MF�hL�}Q���7�i~�V�j+�[Vm��yj�,G��N�
���Nz�iAM;�8�g^�%����-]5B��G��d�������!'��\���ŔZ҇/���Ml@��~���g�dST�~l���F�5)6���^��X��:�a�	o�3x`����-��?�6r����Ӽ �P�;�[l�-`�5Oj�dL�P,�h?��`�uCMVWP�taY��[Go�D��/:�q��O�z/&��]��(��H�%�BDu�Q�'.VD-����b�ܒ[y#�$N��+DX�خ��͑�i�a�J�7�G���hǍ�+ �i̦�x�V�%��e�Դ3h��/G�K���B���f��C@D�hCM�V2oӢ��e����+̆(�F��X���ݼq�\��[B��\�W��<�=����|$5�	̃�b"�u(���"�Kcb߸��J���0w�z
?M\[�g��p�:-Og��!nt��I��J�<7���BE�Sר��$\i�D9��F��Ts���]�˘�4���w�E�ܢG�����NM���E)/;�<G�Ju��7��?k�����(����[��?��s:d"*Xf���É��m�ء@�7����OI�
��*��s <�x�p���
��I0&��D�u��
������Nث/��M�Q�%߷e{)�*v��KR�44����C�����\����qR}l}�@(�U��a5&Ak2���>2Y�Z�t��R��R����^��c+�)`Y󛌏���$!E�
Y�g8i�J0�O����ԃ�j~t�=�ҽPh�8�3�؇��l�+��#���6U`S��@�ī{wG:��߬򧏘6���+�o��R�/w�.Ԡ2s�S�yx>�ܖ,r�|�R�D q�g�{ վ�nN�vP�J�(�< �E��,s����|�!y+s^����,�����-��P+��$���}P�ga��
,͌�$��Q��G�t+n|b�|CC�Li71IK��|��p���և$��';�/���=+��8Dl�f�������B�ces/������%AY�*W�.��5��}HM�!w/o��irk���%�Bz�(�VO̸�8��5DJN��J����*�FNؘTd�j���h0��#}&[x�Lp���b��}�v>L�!)B�0 d{��������:�+*�b��A��x�ѻ�����JU��VxӚ�w�����8^d�ؾ����mk�9��1�xI
�~4ڔ�̑L�9�{ņM�滤�FQ��V���"��w$��&ʒ��Qc��{k�\��8����m�%����̏�W�nn�o��7V*#|���� I�T]����|=�A�P�u�V�#�)0(�%ݶ�Nu�=�ONUz�3u�RuG1����ק�MH���������g�㽐M�D+#2���/��Ry@_8ン��� �8��ã�����:*�xq�l}<@�ٴ����#��X��Q��U�h�,��v*��3�(!�a[�� ��q*�t��44���6 ��|���Q`�$"���&ot��xݺ��\1�2���-M����y�tvO֞Qƴ�z�15R�V	�iS��$5���=IM矈w/�Z}�hJ<F�<�!� ^p=�J���+-�}�� WRe ӹGU^� S�(e���a�����yV��(�
�4o���ܹ0�m���9�\2��n���#JMެ��.l����B�yN�k��p��+���_�����P�_|l�e�>�K+:�cR�2�nLW����Fp���/�C令P:���_�v�2�'�vp8�� ˄O�eh:H�2�*�8�/������~�&������I��t�M�W�ds���� ����.&��(9.*�>5V�fm����M�J�N*�{��o�RG�y�������aT9�r�/��ׯ�V�z}"1����R��?k��3�+2ݷXF�fRb,�{��"3 ��f� ��hFQj�y�/!�:@��:���[�^���se~�nu�"qק���M�"!�JC�cY4��`��L�&K�xH�M����zHy�qvI\d��G&W�M��(��M�K�(u�
�>G�ǒ��l5w[���0���u7�(5ãS�3��@�^��#H�ĳ�݋�2ÜE�螌�7���+pn&�ʻ*��� ��S�`����Z��Dq�ɤF!��E�t��q��]^!�FB�S�х����jC},�3�h"��VlP��J�bH��J�1���)}��㫤�������yRչw'-�?���}1.9UȠ?_u�zS�O�ja������_=���4�m�y�,����^��N�"��+��Ͻ��Փ3�<Eh�t���rCΫ��lͬ�VC�!���nК����jF�����B�$P�W^��>K�tO�ͱ�>M�����3����a\-@�*u_'ޑ]-V��I���B�
��-��;x���yP��I���R!Y�"S� kL�s����J;ĭ�*��j�	�<�D�c
'K{i�۝ 9p�🀰k�n-�_kIܷ��z[�3�n�>�<n���L�9�e];C�4LhR��ʉe��l���:.��j5_!��^�x�f���JO�?��i��y@�Z���2�����p�/��J<)A��
��pm�x��k�xS�{�K��d����C�x�j}���EϿ2��c5���V��������0�v雀�p��t��iD?�Q�j*��%�,AͰ��)�D�pydEn+�ݯ�"��-|xm�%�����A6.V�xHT�ПP	���*Yu�!����fvB�-2(�Ʒ!�x
A_�5�?� V�
�P��2c1��Տ��:�x&�|�~N�Ua�^�l��\���C�Y�:�2�Yvݎ�8�[����M,�L)<g��Y+��z��Y�W#��H
d��#uHb����.e��h��U��s�l��D�i��\ԒT��{��^�iT?�6@j�Bݢ	�8!��ARV��L��b�)�\�V��:�f������Bnw�h�-
 Գ�L���!ʑ�]!�����iE�~� �-��j9Tfɘu�}kH.�xνF��j{�Vy�*��a�G]S�ڷ"q���Q�ld�f\�%Rڮ=��L� ?m�Q�?�c"N�V(�>�!j�����آA�x�9�c�� �I�x�/�B�b���9G���+�(�����^�h�٨6�$~1��$/ws��<N�SI��RNJ)˻ms�DET�5A�C��\4�TH�����b(��_ъ2����-���>s|�F}���
��/�6/$s7|�'��O�<���p�gl2���Z��~�Fl��(��j?��B���������@6����n��j��uM��q�E�[�����8��+�ڥʍ`[��̡W\��Ą!�نdĭ��od���s���f�"sQ�e]�R�V"�Vf��y���tV?]�J�
E��V�(E@���q�J�k�qTR����Z�Az<�ږ4�������4�N3�*m�#g2)0������%�5�%
�	����e���hZ��e�^˃�������!�L�'�g�<Jة8B�l�±�m3��t^���H
��Ȁ3��@�*�B��H{�7��3�,I5&^���T�s��������|US�P��x�����}�F,��gc�V��X~��?ơ�Ӡ岾
�9��THI��z�o�@��������G:��a�'���� X���_�q��z�OX�L���(♶���(�3M�|:�g^@h�EWl�)ʅY^-����Y���U<0�Eƣ$������#�c��˶�֞�h81i��/��;H�ɦw� ���yl��Н�\!�	��{���o��-Rsg��)�`�*,rgyV.�6ڍ٩���6X�o;�su�T,���B�C��Z��/aR���g�1K������������唔���Xf^�*�"8��yU*W�V��D>f���I���+ꘊ�e�.�,�s�z��y��/B=�S�@��Q��p�9HG4�:�q�o���έc�{�x��Z��(��`��N��ƺ�f��c�z��V�Y�yy�Bn�[c��"�ɲ
txT?�V�>Ŕ u�r�e���mIsE�)��NK�J�n]��y��X���X��M��Z�� %��߹��E[2�G��mxA>��G�l4/�����������r��,#�Jf𜪻=�������.�(��IV�Y��G���m���F���Αh1f��r�U���g�Zb[ ]�� &�U���H�,�hpcX���b����{��`�;:����G����<�TARW�^Y&��<�ѺwO�t(�H�%R\!۫b��d1O߆��Bҳe���s(���	��>�j�I�S��r����+Ts���� ���9�ޕZ`#�!3,*/��#e��Cn)�3:�:»6<6#��f���{���� �xƦ���|�d���n\�Џ��Ah���K����\���S=�q�xL�.3���=��1�L���vd�w�'���q��	��G��s<��&�c�i�G�ʌjT��'<����í)�(c\ݎ��̇V�����|'vE���Ј/��j��a��kK����[k�k���6�L� )I�an�Q-|������f䪱$Ǆ~����T�s�d7�Uzj]~�%<��e��GZ�r�!�/����F�m��.�b����ӡ}�l.�P0�@'(��S�`xfxh����K�����i�wݭ�)�W$(Y}{���l#_�EpVɈ��[,�n�ƐJuᛁZ�K>!(�u��V����d\�Y)���T���>vڴӔ�����	:�Uk��CW�Q8����%�ca��t? 9vO��m4v�N���G���bx���9�Z� {{%e8�[3���V�]El�\��G�D���x){%��$��W�qW���4z{��A<�gV�������2�q1��=�(�`� �ܣZ�
�W}�E�V܈�6�^<[�� �ƞ܂'2B�R��܉�^���^؞��G�b�12����474�=fx�h�k�WN�(dz�3uI= �>2��>��
r�h>QYC�������ԉ����#�� 1�h�`�d����!����W��Q(@?�f;�[�l�|0����mp�d#;�x��`\䭿U
|����x22�EJ��E:������'��Ph�s��Ho�[�@+I�q���P���7z6���/�Et�9We�+Q�H?`��h��Fk �UB��O@�q�z�����J,��k�}ū�`���� l��+Gk_Hz��^?���g�y̙��}�/�Իsj���c�#����q�1�j���Ik������\K��hh
*�NS�.\L�!/��gejW�Us�ʝU�c{:D'��c�:}�����X[�;��t�{A �;�&���qwq�\����'��e�w�p�'�s\H�_��ދn�P�v�Ҿ��m.��GQj�� �R�}i�������s0��i�7%�z�T�A(�q��H��+"}�=5�@� _��(���!ed��#w�Q�] ��O��v?*��Ⴒ��K��Q�zQ���i[��K��3ɵBz��iP�4(�Ź��>���C`f���~!J����E[�[��UhH��q�ݶ@NTu�i�/R�C69�-l;������<n�<sF�fh��m��'��rr�x����M2K�&������>���F=#���!S�2$9�z		���kL^�9��~�.`G)ͥY�)�¤ہ���&y>&�?�Ʃ^�< ��sM��Fb�O/}�#|f�v\D8���D[��>�e�UV�7�5�O�P�~�x��N#e�e��;��ն�>G�󇆕l��Y�(�����YhY8z�,�F�v��'�qx�%�=㡁�3`����`��a�_�H���������kX#\�N�i��3��nh~d���pw�lL���XO,&���(��E��j6�,g�����A�뼚:�(L�tj��1tW�::��᧍�5�@�ގ��@)O����n�	�8:�<[c���s���x�]>Ү�|i{���`�v���U��c?�B��S�%'m������!��ơ>��n��|H-�V���NW~"@���S݈���y�ް�L��X��@�chA'�`�C�x:���"$�U3�z��ř9:��U����}��+�Ѿy��Ґud����8x�S��_Q&���$��Rv4`�������U���ei0|(d�H+�d5�T��pΊ�G)����='7���T�Z�~&��pŭ4G�y��3���f�S��0O� " Q���{���\"˛w����L@\��2�Q@����$>b�(v�4�U��#���Es�a����Z�*M��ভF��mX+���y��H$�����9Ȧ�
�W�\"�ʀU-7��o�j�G��iz��L�o��# ~1�i�l�K�=:�qy �R��Ay�1�w,���C�ҿ�"4�Z[.��xXY����Л��D9�F�sWw5t#֊|����A�NU�5��{7�c֥�<1�R���P�a87- �6叧O��mԖ�8�J�.�?Kp�dt?_�`�)�?��Gq����)������,1�J��%H�Ǣ�͒�0��Ŀ�C�����}w�|�˄�#o��Qa�8T<���@�ݞ�	z�§���@`�Dr�\�0A�|Jc��$>7l��*G�nF�X���Qߖv^����O�lH�f��p"˛04�Ju�&�����S�X3�I�����(Z@ez��ҟ�خ���6u����fօ��N��`���%���s Q�OʕB��?���[�b�#������*fc����)����h�"ΪQY�F��)g�ږ4~2�<�:S6���n��쯵���^8vr�e������I�'	���]�r�����zFP2�:}��]����[Ϯp�o ����3����_����;|67������/@[��k8�w8���#<C�n�m�6�*��� �UF�Ez��Ń�H�Pg�ii��>BY��W�~�t�k�b���Yd��k��A��X�Ǌ+�3��5`E���37{+� edUW�8�r��Sd�A�|S����>�� ��Cu=66�/j�S�;�MN�Y��ږ����%�ʣ\�p���Q=cё�[{��76�A�U�5�|Ex��:0����K���pwl	�Ah�s��d��x�!I7�~��g�� ;���'����m�>.r����*���떏�Ľ����b`�N���$n �@f����M�b�&b*�q��r']����t<.�v�r1�p�Nk��m�h�#S\
S6x�>� ��T�<�`{�^UJzܻE�����<Ğ���֛V퉸�)L�hC��̼��BL�}�Rۧ<R��@��-�_�)(�(��aB�Q��Q����Z��wU
k3o�C�L^�㌤��̔7��hXȩ��f��Mp�3��1����Y̩�Rde*_�(n"���*
'c��Ϳ��o�rV�|,[hEv��ql�@)Ѿ)2���<o��8�]����1���o�3ԇ��p���!3Y�H6�V[�-%��Z��[�5*ݿ�w� ��o����i��!�����
R�y�'"�g�����|�`�~_⺬���	���[Gz��C�-�YOK3�Gsy���w*�M<��
�T���/���$U�}�� .���J�^�{�ƃ>áx�ݕ�;N��\�[=�����=`�ń�����lo�#N,h�ɠ��D�~���;FAs�a<E�6�#��DgSK�r
�ԎѴEfZ7
%�e���_b�
����x�H.8��
'.��ATG�| �)��x ��1��g*3��dlt��<r��/��1Z�h�5�ZeS.$�(q}#E���m����������1E�;$�RH��au�v��x�
pJ01UyԒe�*�RP���	���(� �=0B ��a�+���?�jx����,x�k[�ѴB���F��� )�)�W���ۮľФ�c2�&(?e�Do��7�oQ�S����.�Od����_rk������s�f%���8�nr�l\���-D&Y����=[ʋ;ʷy�[^���������b�3`j��J�����v &B� �S����90�m��5Bg�::NZe�<g�HFQ��b8*.�� �����1_���.�����)�*�`�lDϪ�Y��XP�%�}l�txM:×�Z9�2\����n@����\6�(Z���vz��I_���������9�#��r�d4E�� /��m�X�Y	����3��x!��\�Ќ�_LӼ����l�B̖+NB'���<�]1�s�ܵ/ ��!�@`��w�60�د1wV�2�׌'y৊Oa�0��*^��GKC��"l
L���bW`y�:8f_�b�n�!�Z�	4y�a}ek��x��RXA�����&?���*�O�"z�D��E��B(Ò0�Gz3hV2�v�=;��n�)t3��z~��IթU3 ���8�H�]�+��N4-��[vR���S���������`�y��ܕ��~Q�>h~�M��^��;�z�^���y�J0_�R�|��l<�*��J���3ʴ��ۭi'%�Xb���jmb��*��k�O�N�HsH��z�4�����ěS�A2L��Q7�-��;���Я�Y�4�QLϣ��>9(�.S��KB�S��<'����.b��b������6Hq�o�X0��#K���h�m;O�<����I�����ˍ�l�V�د|S��a �;��֩��A1u+X��j�1�_����#�ە#��°E��������|0�{�ҹ��1d��򔱉|�s���La
�4j�<y�� 4�C�.LMΌz5cY~XS������S��^h�m�
]krDb1�6���K��g��)mH9j�T��؈�t����QlȬk��7���q���58=�������?�0��q��Bk��ݨۚs3�ݕ$=�_�܏gw��b�x�V����i�����@�r�#x��v�	k�$c�7�ɼ؀����c����Q�W)y~&��n8���L�*~�:(v3VH��,��ԂT6��y*��?��ه��_��j�;Є'�4tr`Nؔ�R���h���2u#B8�0�_g�\6Hr����f��ȕ���W�L��v�I!� D���ӎ`��44�����$Z����aZ�xд�Hy�i�ǯ-�3D��>i��st�#4RIC?����;�9��8˗��Ǵ?���H�t�)�9�l��.�K��{��2d%OԵ�~[�tH|�a���:��@r���z����z��"�ЅXG��<)���9��L��v��28�ʜ�!{7�q��k�{>�_F����E�L9S�|������=�K����f��PJ�ӈ	�=�\<������1sS����b�!8��{�p+xt�I�e\�J���K�#���d����`JS���Pm�'�ʆ'T����7���)@��"��M	���m�X���C�?P��8j��u��ԧ8�݆Mºg��Ĳ�	q�5����DgrG��ϱ/��!��?Tp�X|��#���iG��I�K�������t�l���_����rXgS�{���>�S=�U �Q�8`-�A�>� ���3�8���1��{ǵ�Vֹ�jȘh}�*63��W'�7HN5|Z�/9�H�{BfJO߱�gh%�������f�k�*�Fa��G�b���To(���m�%V�U�u��}Z��!�Jȳ��V�V�U ���܃9j6�O��7	w��Z�p��wĩWB� Ӣ����?NP���pgLt�xQ��>�#��˅|���J1�}�[~���ۥ�o϶JK@'�z�H��2���Һ�ǪM����2aꑊ��o���fF[�'՚���D��zD3�x�bG	���<�"�9�r���"����N�"@ZV�r��m1�N�1k�F�#I�A�����*<�X��6�S"ڼl�Mk���O��#t~��m�6�7�U;=*��M���ԄՋ�ޱiҘpQuYۂp�0��mjK���.p��_@���#8��e���MM�̛�5��jk��ǖ�*���#X�ۈ- D|�dda�է�xޖ�PJ��u�#��7��I��:$�:�K��>�&�����F�2m�kꊆ��O�<��9��|OJ@���ʓCiJ/ۜ#���Ip�&�y���i�Ԩ4vq�8!V8@K9w��xb5��H*u���Y�p����`�����h�ܩ�L �"�?`
�Ft��A`�ܫes�!���}���p.�y�6m�vq<]��t/t�ՙ��-�^�qFDl�l� �"48��΂E�j�B�B��I�D�gl�v��+��V!6H��y�g�GA����9�󮙁=�<\��T��s�5"�݈Q��i�nZ���˿�\��A'�,;��[b���V��0ǚ�oE�m�d�
���?VH/���f�Ɖ�2(+��ua*�b��|D�{Y�u�z���X�\��eϕ��\��� �xm-���S0{�r����!����A:W�9bciS2�a{��ߊ��9���4j�f�W��XkZ4�?ޮy!Q���14�CQ3c�c!��H1=���,�kv��1���0�A�2;fJ�wy��l���ȧ����Ȇ_���E���z���{�ÔH����r�NE�&�U���ŏTL��`��-u3��N�ngW����xT�*j��Ym ��������d�j6���Kly	����z3�[�H�IX���Y���&d�u1����jm��T���w�Xp����I0��C7���C?�f���z.��s��YW��.&���.�����i�׬z�	���!��%xM�S
_f���4~�i�o�ᰥ����8@��o���s����>1��/,�<3�R�C�e����l
,�TAWV�)	���QH͂���(?�]�N���� �B�8��+��>b�/M=9���>��l���,j�PO$����-
8��|(S�=:�#2n��IY�E�/'�0s��"�x0rB�G?��^(�#{D@�^^,#��Dd����D��W�^�&/��͉����R����
e����6I2^��W�QD�g��%��� >Jyb�Dt�n�s��W�̷'��O��;�Ƒ��6u��Š��Q�B�\�Wm{r��75&��a�{�PF�@�k"Ov�iC�a%/���KG��r������H��1+ɊD�lZP�F�lA�9y����:��2*�ύ�ʜu�Ǐ��
�6fq���l�H�L�2���:�iX�9f��wn���x���h�\j�����1`�2�FAQ�8잔��ue&}�q�v_!s~6��ݒ'��&����`��������8���k���F@��4�+wg ���>\��<� �ƃ)0��cΐ����t�"N��O�TӼP8hm}S���ߕ@�4�v��mqN���F#CB&Z��s�k`<�`M$^)wb�e�j��,�e���� 	�>�;�ց���*�g�wL�2�5����CT^���� Ƹ[��|0P��J���9A�s��L]@o�Ԑ��x���j��������ꫣݪP�|]DK��g�n�����^��.�Â.��} �s���l��u�:?�O zt�f@�!{+)�
v �Ӗb���]wX�	���C���G<���㲊)c�<��y���}=�}^�C���2�j:'(^g�w��:*Ҵ��\
�!���UƝ|Z�(�jGG�@�1'n����iq��x�-��b�3e������C�_��|lR�d��q}_�_�s��9�Ú�z�����2��U�x���X�c=n�ֳ��}e��4��YJ���vff�/��f,WJ�I��Ov͋�Ur�l���τ�z�?b�[~2@�e=�������zM-� #:ĜE��zǃJgA�W�@�$�7t�������ֳ��=��9��W��ϱ�`)u|_��͖YsE�.�S4��\�N��q*�\�Z�ْ�{9���C�AKۑ`����8Sf]�(��ܖ[���e�`#�pJ�D���9���]'��Mz?�0PF��'4!�G�*����ʼ�!�A��JA�gD%m���� ��Fx�}8L���n�c��Ə�6�^�aX�_��Ǳ��F��f���4��ݟ���6| �L�T���q V#lBB�=���ƀC�'l��K���K�Y}�+��@0>�%fƘ�'�h4.��D{�o���Q'9�kG�US��J��px��忩��V�P�*��.|.e��~���f��2[#q�v] %�kZ��Xp���j�ekd
��p\"��4����������kٔ2'�Bڭ���[��Az9�d��::5D�K�Ix0+��Hc�oKo�w�&���挸+w39��w�t���<�R���d�6�:���d��\ �Ahv�qZR}ra�MOp&`�%2s*�DY{��h��L!��jC���Q//��xS�V(s�{$�[���e��8�zΖ�^ud��X�_��i$�\�ض\��H &
xq���d ���j��s|���׋����{ky۽�5��R����K�[q�N�n�&�N5�}��԰�丹,�����aN���3K��d�)�tK�9��@�g%Jy�=_g���q�/���DDwT�`}�����^��d�UOzZ��S����|&w���OQ]ǘ6�D38��2����ҿ_��6��l��"b�Bɂ4��a�q�k�:�����Ǿ7���K�����B�������gV�@J�^�ꪛ��co���
����qP<w_j���F�����ZZ�8yu��:�Y�r�#n�x���Y���c���eǥ��1|�(�f��ѕ�����r�/����%�jPDRfp��7H�},["c[/ؗ7�bᦄ<K�1��z�UB�ҷnX�JsR/G��E�ƗlO�KlNq[�|��q���<IoL���S{ Gٲ�<�����l$9a�����T��4�H��1h�m�`�����~Ҕ�����n!5=R�S���rM��t?���(A�D������H<�
�0�L갌��/r�ӚS�hK�W��%E�l�������EB���04c�ꁊ�+4{N93��Gs�X�1}��B�V��o��w\��	b�+���g�v�
����D���F@���?7S�nE�^�00�[Z��D ���
�p��aV�E��� ^���I�!Ȕ)x+&!F݆	��,<��:�̚�t��|XT�&���ԛOZ�mߎ�)*&�«�m ����+�[�4�10�<�+�RQ�6�H9u2
^��Ԭ#�*  M�K�d���f�8�so�l!5S��?��.�u�O{�Ʉ�)b��ɾ6�c%��ȇz��<ɹ���*�EC�b�/h���~^y������\5�5Q߆�p6_�t�%" T����Q#��p��9w�����u�\��U�oSV�[�qr�c�6�rFObǲm2�Q#�/�OAn.k	*���3�F$�0����H�1v>��m�棫OQY<E>�Gz���G$2_�z�D����to�1��-+:�]Y�X��U��~h�U�I?	���m;��$�簖�1Dk(Y]��	ݥ%[��.�2tm|91�[Vw�8�E�C�݌K��QiD��Tt*����Տ�T��n��ne�"�^�B]��� ������*�T0@.���P$�&U0Z��U0x���9̬Gjn�`D� ��q����n\>\�`M���Ԯĩ��È�4��G�����2"u��dP���"Ň�CP>^W�<��	k��fp3���{r��(�a��t�繆N��M�A�N��0Jr�^��s��ӱ�� � �p*4����'i
��:�;��lW�L=��$R�wq�a�Tz G��&��E� �"�7}k��^���Lb<6��VL�UY�����6u�ri:o��V�s�����V�I�E��M}�
�w=@���<{�A��~ ļj���l����jY�y
� =b=q��x�(�g1�*U��VS�;�F�`4u�o#i����<E�r���3+O�� D��i��	O�!��i�YZ;�����w&*p�s��*VƏͯ���N�N� �E�GX鯤n�쩫����Oc���%��A�1T�!U�!��B�������ѱ�i����D��}��.z���>!��^�E�G
���#�@�	�bI�{7VEp����h j���B2��`.2�D���3&}:�=h�*�I�%�/���1gJ7�Gגv"5�F���~����Y͡Y�*^�ݼ:	�0<�����/J��|�z�B�$���|��pß���Я��Υ�=�׳E?[+(1�#��{�3ʹ�n�a�;�,�w���B�5�E�t��6��%��AA�cWAiRn�U�؍���G�gJ����������G�Ab&�d���2�2�)�b��71c��~p��0w����M�z���ٻ:�E���p���Y�	�&a���xF3h���Z:5/`ji��R���q�'gB���ў�}^�ǳA����2!P[��Ǒ��2�]荜��b��(1ޞ�).�͆�m(�/.�3��:!(��G��G����Nv ���͐��Y���(u�/��c�IMq���,
����'�@+��cx����;���T��̋\H,�5����!�5�nMy���*@t�7�mj.$2u��S����W5��aN�:��{YlɌ�#t���W���3�����7N;���8D��R���ȁZ}������A�Nտ&��/�U����nG���V�qD`�W<ϚT� ��J���F��P�&�9�#��c��ıD	��ߛ妫����w�Z�N5�&.��0�ø�VE��ym$Z���Ex{^}�凗L�s�)Q���QS�p@�J>��670�e��%�v@��%c�BB�ƽ��ɫ�/(�u�5� ���^L�,:l��h�EbF%�(<"��'9�:F@i��B���xa�y��������Xt�s}���K3oS��V����s�H�����>���m ~ ��ٻ��;�TzQ� yѬ�k�'� ��C��*��2XS���[�z��`���?��^���^~���S�Q����	Ɠ���W%��7��w���bOx�zj�f^�N��8	�܏�ޗH��pn���0Ƥ��S������k����wS
�ǐT6׎97�Û�a[��=F"(*T7Œ��t�>�f�G�j����Y�j����<-���ÉD��6O�u���l��I.��݃����&��Z퐒�U�O��ۆ�o*팼5֭kf�>{��΄�q��u%2���iY�SDr+y�='�3˛��������3Ep:*J@!��œ7�=A�0m�M_$����2��C'0ܺ��1�_9�e``u}OB<6s���.�V�0R�H�S>���/����UӠܔ��p�[^,�ǥxq:��G���{ZY��|��J�ݙ�Dv�{Q���ml�c-垘q����}xA�\>�oDx�Q	�e���_���&S�1�F���O�8��m�/���6gE����75f�ư�D6�y���-��~?������$вg0J~Ѥ�6s��Lu}��� ؼ�˶ۓw�S���4�eYL4Э͐��*avw��(�*d?s���f�]�x�\�=�򇏯n �>i+� ��U@P���w��ϔ.����Ae����+�Fs휇��Lei�q�F!9�KS ��L�C((d�j�jl#�|=.FT�i��+��YUDm  `o�X����e�&�|:{�T�g<�s6t����������7�Q�v~��Kpfc���Ԯ�?ŞR$Qs���w�(�� �"��#󊒵MƈMD�߱=C;LBf�f5�i�\�r.f�p6�]�߼��������%��̰O��K��@5n��,ͩ�~|�9]2��4�}%H/o�O,��i�Xt��zDI9�LMd1�D"]�g���yC��q�����I�g��9x=�Al�'aON�
4���P���o�=�_�z|���x�����d�����cL��6N(ݐf|v�I�邦��7������O�I�vx��ہv�%O���}ϸ���?��Y,E$1��00� ���dr��dexO��G�ϕCtf�?V�f���|�+�j���ʑK�_V{����J�4������t1RСŁ�H+���`�@n���KIzph��P��e!�^`����P<��+J�,���TwX�C�_�|�el!\�.��m�<�F���۫*�Qp��1���&�����2<���«Ř>�g��3nKLO��4VP�B��?i���<�È3{��.�Y���P�Oݺ=��u�I���h>�Af��-��o�c��i�a��u�건ش�掙\ً�a��q�$=W�$�X~�m��»��#oV�b��\\�}�O���JUĆ��׹}o8"�Za�y�Eԓu��u����z̐�n���A��8����9#hI6�9k$�W0^n�G�R��U�%�7(�q��^1�r�@4���x�����J���-��28��>�n>ji�6D\�B��:�th �e���2�1�ǣ���Z_T���V��� ~��:���*� ��"��$̳��!i�8�苉�+C�/����	�ܻ���ۤQ-(��qx�soy���#qgnM���ӈ�t��%Vs�tm2�԰Aɳ���e��2�6B�D5/u%�>$j�~�lNc�E���T����3s�'[?�e��ti���5�_��EHhP��*�O���_�M0b�5s��"g���a�JM8CG�ʁpl��^m���kS<�r�A�s�Z=�O�y*/�f
�:��|��5������U���w�Hܺߒ��`1"��Mh�&���s�.m�O[��Pݻ"=�S��"|�k���}6�kTO��Ȩ���-����e/�`��p���D5+.Ql�m����B(p�*,%�{�c!���AfUb{�>d6KvQ�ކv���\��vu|��Ȣ8�&��A�³�gP{):��h��)���ݑ#��v�X����4Y�?٪.���"���������e��)`���{f�q����<X�V�Qt�����d_8��b��FP�=������^�ef	93����l:��O˕�����~5t�ul����Nwµ3 ,fY߱?�8NeyýG~^ç|TB�2�{M>���mp8(��8��F��[Vtk����)�[�@�g%��ڻ:#�<�p#�뒻�l�P��Nl�M��R�[�9� y�����<�����PU�r�+*:�D*��a%]�ə���:Vq��s��Š�ҁU�����Ʉ��K3�y$�:ԗ����ɽՉ?\�f])�ۖ~�H�NnYV%���˷
�-��4�(&g�+�0�)�
P��>I��g߾w�ƙ*Ri�20��_l�9u-��K�כ/�6%�i/7��|������-y���nu��z����D���]J��坔�
�����Kdd��y��O��xS�l`��yV+�DI�����Ĳ�A�2`��	�Op��<�{I�V֕JB���{�c�c0=�Öa�nɯb���3Ô�F���J��)��`�2�* Z��V_\�����d$����Ψ���n^��}������iQ�T����������a\�,99/)�&�Pc�C�,M-����JwA�	�{J��]uq`]�n�C�6��<�h�c��$�0������$�����#Ō��2�z�8&8(�����<�dZ;Լ��S?]�1�uk���5��R�`Lۀ��R9l�d�DP��8��dZe���7V�p��<�!ozR��)�Vü>��;�Ɇ|�a�S��нr�����G��^���p �ݣ�a�?T� �$;�[�l��e���5}�œ�>0eb����
��T�|i�i�M!�5��a��a������:�bo����s���8��mH������X���;��"8�b[���'ѡ��~��Ո7��!>~QĠ̒�#�K5y��@���f�_��z��j��LR$Z�X�NY��$��@���������H�}����oCjq�:�������y���a`�!�	�9L@/��GM�L�{����khM�d��8��y�@�WW��j+��s0��aR����O��D�퍼��\x�����:�qN[o���߆O6
lCc/��{��3�f��]�C��D��h�-���̢��Ƞ��u�K�ƻ�z���l�&�w���M�χzy�*���`y�Sm������"a��o����=�?@���$3$��'�H�O9�zr�p��0H��s�YG��'�?�v1o��fs�_HL��nW�Y��}UHBPɜ�ֿA�����bG	�ҽe�>�&T7���g��z��JZ&Q�4_������#)L��t�<#<y	$����`�iJ��;�3��"�T�k�m`,PU?F�Þ�J��"�ۚ�l��$�i��WǾ�MQ�0��.m�:�[�넨����+<w�&2�<{�"��[���t|����R�r;��n̍�d�Zv��ւae���pw��F��J�Y�����v��
!������1�#��~�WU-u�w��F�y����	rBv{+i^�9F�hc���ְ�I������z�fE޳]]>3+g�@�8������	J]d
'������5g :�E鞵��L�Gz'���|�92�A�S����V-���#����8#i=�ޔ;
u��e��L:��m��⺤����U���zqnN�����`qg�A�AP}%�&��1��B�I�b���g_^&%�5�a������_���L��ɟ"$z��,��O�Qp���]�U��IGFIn�
jW@֧th�H�vW�5C�lԳ��6ɒX�3��cf�Rnje)�xoJ8�4[�E��ZʔX���0b�HAD��TK���\i����g�w?�����n�<.��1g�����:o���6�c�1�������)#\~�����F����2�H:��.Z�~4�%�v&P`;;m�Ɏ��2���ʩdY{8��x��}-�lD�/\t��
ڲ14�S�;���!	��ث4������kk��[)<���VQX�^������Zr��7V�:�I%�C0*pQDA>z�?�}	4����"'���G�p7O.���_�8�t��x:�i@���Kgᭆ<�KD�J�����2T��>S�[�t㳞��w~[���0�=�H^�Qȿ�&�����Td_@�]�,���1ލ	ߓ�UQeKZIT��V^�ü}k��)	,MM�{+u��Iش�C��]��B���/m	�c��؂��B��d`��M��������na��iI��b3XXt\W�g��t4]��}���.�~ь)����>��^�I�Z�h�+�x�=�B��H-|�.��'��s૖)W�l|��o�D��k�8SW*قO��X$��nK's�	�V��H�	m���	.k�%wد5�(��0�XS��Ȥ	S�Ͻ&��&�g�:�����֯�PU�ž5���^��ӝ���A�����q!����f/��1��1� ���`�:!�PQ����p�o���<=r�j?��	�l�$<x�"�*t�4���k����~v)|���؝�F�!��<s	۶��ߜ�
JK��b�_�Yh�J��!��[G@pN���3P��=H���N:�_uoz��MMU'��)��S
ep�dG��=�y�/���dC�nd���ta�k�{���5�0��[ӥ��0�3�3�ס��gcF�i��"3� Ns��Ǎ��va����"Y�/���b4��N�\����	��D�/�i+X���u�!���o��q��Đk����)dM�3���A> �x��=�8����ia[�ր>����ɠ�I���P�/9a�/�dB�!H�9w4��D�Q�k�j`�����+3���9rx��۲i���o^H�laq��*k6
�G'	U�r�ы�$���$Pz��`;XPGT�"�/�iD�ev�0��ȱ���B�{S�Ϳ[B��6U1��|��v�L��ZU, Y�%�I���������U���`��t���/�2�,_xiЀ�=*MF?��l>���$�[�����1��:QL;|��I3N0�!�t}3L���Vnd& ��O�d1���w����7�&	|�v��^�m��P��G闞h,�]�:'��JX��Mv;�ٻ&�P��Tb�-�j���n	���=[@8O鞪I�?�Y7}�q{��7(�U!����U����u-���k�p��9Fw�+��i���:9Қ*+�{!����.��jW��}�ju�l�(/�o�j+�*G�\(���*�����q����E�	���>Ɓ�Hd���<��9�ˏD}�B��+5�b 1�j�?�J���W����2��D�\W�½�i���I�G��ˏ�=�-	2�@2�;���Db�uE;�J4��H�yB����& g�r�!�Û%$sU�PgZ�7HF���s���i� �>�������1�v&����PD����b��s�a�ӎ��Wc@��zd]�7TN��~ ���B\9ಥLG���`�Q� �����8")@T��}\�Y�_.f�{ɆyUR��/5����/4�f�[텿.��HV�AN*�Z��1�^��ǀP���2��~�q�'�E��ַ�f	$9���r� T���?��5���c&#�����b�aM��F$�u_ 70����|A�[$`�G�D��ܲ7�7��2{k�lNYCt�&����~���sy|z��PI{�� r�A]��k9���<?�>�C�S}��ʪ�U�=�M�X;�õ$�o��QȄ�r�Ϩ����]V�0fn�2��T��O�	�����(�����	�O�@�<1H�h[\�CQ^Z��FL��%�w�Bd=[�$�eb���
zf���hp	ζrBj{)��H�C����Q�\<����$o�'�ߨ��,Y�2�Zm��<���ڿ�`��0��n����Z��E*�;c�#���kb��s�Z�h���ǏS���I�̰��%�īf#�-{l�]}�6䙨���Y�'�Ok��؝�덃�6�T������c����`�K�z^1Uڛ��œ����DG�g�r�²�������o|�Z�<ȭO�`�3�2l�2W�@:�H�i����m��=���f�E|��`���f� b��j��>��K I0U��=���Rl��h���Mq?�?���J�`�q�ie9p�5�U��|�f����R�V�>�[����'օo������-�.(����l������+��Haە�"P�$`�?8u��;Ǽ�Be�tC�2[�S����-�j!O<8p��L3,'׻��<�G�I��ɱ"���"#g-��BҼ�I&ړ/����
�\��˜G�n�'b�tp5,K3��_a��B@M&Q=WmOJ<|h	�oؿX��kK�c��������Wx�HY�`��d�TӮ���,s%1/���� �`i#�w�t>��*��iBؤ�������Ɓ1A�1�^@sK��v:�B��f&O1#	l04�g<�K7�(�ީYq�kÕ�r}���Rx����/QՌ[�Yr��8{��������Ǟ�Z�r�Oc,z���)����P�Ek������8gs����W~@C��=�A(E�	�Ÿ8|싔'͘�&G�4R0��� 3���6�И�@�q�)��M�Eh�A��2�r�W	{2d��t�F-+�Z֖�����/3�x����e�ϔ[ivY��^�s6�R���I���UPc��dCzv�+�cӎy�g� �����/�b�5��ܕ�1�c�0 ��\�M��kخлEF�1Y"ό֏�0�"D�upہ���c[�����`��IO���5>�s;E���G'$y��v@�w�J^N�z�W&����ޥ�
�np��M5{,�ۗQ��QBӨ��� w$���?�����T�������.�^�����,ֈJq]:9l���P2 h��j�w�-U@�j���2MR�G5t�2����G���b>�|T�\��4QREr���2b�{ �j9*;U��V�{��+)�ɝ�m.d0�X1����� ��Ю_i��.8:�%|s�t1V�o�͋�Y8>��z��|�ڞS��{�%�8�Nٜd�茣s�'��I�J�S��<��0�x����U/���b+��'�3�'��X�6���d������eVN��a��79n������;����i�iҒ�T���xb�U��sX��P��
2D�7?̠�d��W{t%\E*�8�柚7��K�.x\����;��?�pc+�%5+�@Ōj��;��t�!���GL
剹���<�N��$)e;De�Ʒ��L �������v�v� ��9�켼Om2=ڠ
څ����ǐ�x�ֹ#橸����j$RZ q���H/���䌒�>
�	b+�¢++����n(�^��i���t�F��r6��Ͽ(��%%�p��U���A!�Ny�4�d���rYEb�gG�.t�Š�cv%���0�;�^�xVJ�O����
�>�hs�ΞLglR��ѵL��n�ke�͂.B���oC�ZN��{���x�#h+}}tp���*��e������&ֈuk�V����~��UU���%T�ԟN�zY�t�8s�j�%�%\��OO��-��l}C ;A������\$�I>��=�0��=��:�����h��і�>���aUcV��JAa=����3��S	�� v;���kM�(2�l��/B�ޓa/�	`� =E ���lɪ|zG�Hr�л���hgն�O~�;i�M`���a�y�*��w�S
2祮t��ܵoҨV
;Ji��|������0�Lf��&�'�&h��¢,� �c��ؼ�?����X$h��]�b��fsF��9�rW&���/!d��iw��OP���#�e�/�ۺ�^�M�a������VI@���mOu�N{�AI �ZWf6��*1ʞtc�;5���֣$5�t���9�ʦF0�%�����]��#cU��Z�Py
�7.�Uݡ��Z<�`�q7E���[�%J���k��o�}#��0�?'��:��@�4r,��0b���j�?�Ô�"|ս�X 	�z����~���k&J��(�)K[�(�6��K41r�ܻ�2��&���T��fwy{M���ȳ�����#�� &?�f$|����_F��^�����Ʈ!B,����������[��d=�ݭL)/*,�#��G>�W�N�J-�N�I�F�΂iy��L�����m�z����+��9@�w�]A`�$ W$�lv����� �0'���>�8���A�0rs��z(:\ty���[��+Tf�^����Z��X��b�_��$������b�\����}�1��TYj�I����z�>��mBAŨ�mX$l5���F����ľ)�b2_�
0���No���H/���"0�8�����Hmgn�$.-'�g@7s^�t9	�ׄ��x�p����\��i�O�o��-\�n�m<e¿P��}A���v�)Y���8�d���LRh@��0�X���8�Yd}�͐P8Po\ #���3�� >j�6Im���#��]	E��ݻ���t!y�l(.�U2��+�� ɑ�f���s��A��P#�/#���]!�!c��IBF����ύ�y꧓��&`�%��a�ޏy���D�Nd����
���CY���w�>�����N(�#MY�q���D�{�l�W�N=>���4�Y='��0��0��7��'XIsxJ�L���.����J��5�M)�A@2d��9 '�?T�/�q$dØ;�kk��N��!c�QC�������j�U�+������9oJQƧ�4
"\�Ln".���*�<���6?X]hy��yn�Q��Z����P0�}Z��i-�Y]�E�[��5�)��4�-q���"��uĔ�w������0��^�uyXF� ����4�9&7��������lY�Q��G�ٍ��&��I�	�ށ��_T9m��WӖ��q���)
�p1�3E'��}�+���`(6A*ǟ��T��#S��EE�#r�xɹ9��ŌW�Ԕ�U���zΟ[����M�񍺻cʲ`�&�~��	��Y����=��C@�,Ez$\���Lkbկ�X��Fз�Q�(�[A��ԃ���̦��iz��@F?��*�7�R��r��;�J�'�Cv�f���7�)Z+�4,��rK?#񅟗㊇P
�q=�-�#�m������^wN~�z�ąs���W�h��c(53�(^�����T}�\�2�� �����B��*���ɼ�?��=��;t�x�I�/�d� �H5�WrS��oL-T'eYQ۩�,�8��菔My8�u��R���m��r�T��1�bR��%"��;�%x	������ �!���v5d�j�}�:C���i�7V�&�=t����q�� �9V2�h
|��[>�[�x�/�v�[(JL��!i�&�?����e��hO��l�U�U��^+�%�^�� d�Z_�2t���!��m�o݄j�-�sW���{�-`�g':26�BK�z������Jɮ�L����y-���)d�a�-'���D�O�V@j��Ț4��fR޴�2&Х��G��]kp��gy�-~��i�
�kz��s�^)j��EI�
n�
ݣ�#~�� �� eUɴ]�*��伊�J��k8.�~Q�f��#ې�����U�&N�Ọ�4�l^{yd���U[���R*F�z�E�Д�����S6�/W��"k�L?Fur�^��;�p�Gn��%v��M�%��q�3�>��{�V��{I�x�=��\o�|p#�N�&Z����dU�6(�P��⚀���j�FW(3Xt��9?�̩0i��� �隆i��M�qZz��L2Zj��9������i�+�nIX���~A�| q�� �iH�{��S�gD�:�p�{�U��������n
=�1���H��,��R�JU ��ʰm�gw��7^jlo� q*��c(Ӄ��_r��-b���H�	{�I��ZѻZb�Öv�g۝M�dG�/H7.�W|��O�\$���/��#����]�A?���3qlnPip9e^��;i��C�`?`����7EN3��t��&���+��m���\T�0�ƺ�E6׾�"�_~�� #�H%)	��3��d冠b�Ӷ�Y������^�"4e�R
�-�]��\�!x�v��G	+V^:&���c�H~1����i���T��C@�e6B�����Eql�}?0��s>�<'1@Bt���
AІR�9�����_2��ɸv������$��j�M�o��d��3v|IiFR���`����zXt����?A�9�g�<.�0*�5��7�oV����;eM�.Dg��rOC��Uv�Q۪8�7W`�⩸��~�i�'ϲ�bd>-e�Wh�A�L�����e�C�;���@����@q�ް�d�+&���ʪ�W�|s���%����e�V<ƿ�]�>Wc����11��'L4�!�i�F.M��dm����XWK���&����;ni c�O��?��l�MԹR�ϣ�V]�x�+yf���fa5O���}�.�٥1JZ\�I�k5<�Q�2�����0A����a�x��P�����ѣ"����L�6?W�z8Ґ>JH��k��BExW���l���hJ)�k��i1�g)��#�t)Tm�:�eH��o���)}=�"$G���A�~�L'�����w%�F�@�y�	��C7�����|���BQI�QW��g���4>Ck�&�z�ϰ�N>oE�ל�����F;��e/�d07O�N`(�S�>�6Y,^*C�b�^|� w��m4���I`�5V�e�#�8���K�>`f�G4ġ&kf��n�(�����66ԋ��D��������'f�:�+�LF�_�'�Vζ!:	Ulp?�w��8��eބ!
E/$�c#eeWw���n����ЌѼ�����o�xّ�v�7D��M�cs
�`9m	jx߿Ce��P��q�nV?��)�OT�շ�)B1�����K�RBs�m�U��2�����!a��+�~�����h��ݲݦڋ��4�)z�j���o�:6�����F���U����տÄ]uQ'���Չk�S�y@,��۷(�n<|,:�DO�R}��XA6��;j���K1�ha���iȔxl�0��AL$�0�B=n��ԁ�&���~�x�h��Q��D��������$\}H24 �!v��mQ���{[��pu�ab�� I�hk�b�?θ��1���ƕxu��l���hI:;��������o�C�1���֋��ޤ:�B���׌���P�܈����pY�v�_��:��6ª?��-,fqL 6�2Ϲ#4#��D��f��BR�Ѡ��I����
�8+B��ڷ]���xo�}r��'c8MT睴�u�0#An?H�WY6�:f�ؽ ��cic;��0��=BX���+R擲Q�q��I@z�*�섵�9�����)��$����fg�IS�>a�:��Y�ĸ,�:�b�ϰ�V�jC��ʨ���.�w��އ�����ݙ����<ԍ
`����0��m�%�|�n�n/��s��((l�ь'�����4�<�*���	��,���"JG����p�a�y�c��km��H��X�O�g�.㹅Fc��(�75�=e�c��:�]�k�Ӌ�Qa��T�*:j�����@�Ѻ���G��_:װ@c�Me���K�S��ކtI3QK���c�;P��s���%s5�Hc�v4���T>�\f���*G�$ �I��lT��ͧ
t������<׸K���;��sq��P#�W�w~�-�W�ʼ��4{�UCG��G``����5 F�អſ�i���H�/㊯�ڬ����L�n�(�`(��׸t�"Co�X[3�MP|���K�
H!�*�����҈�0�.���gY�}�{P��������[l{���å�3���GQd|]
@ ���k�M��V�eb�&���R����1o���C'�n�)'��F����oA5����H��(F�)4p��w@QCȀ!��dh�9�+�x������j4���t|?I��-��K|Q��@����Nf��L@v���*�WS�#w���ȡ�C\�$��nhC�>CgKk��%�q/�֖��O��&wKp5��#���V�>UR-q�;�;!֓@U�4�6[�2^8�g�����]�\��kLoG�,-F�Y�rA
2���]*.	�	��_L�;��JZE�>ҩڞ�����I�K}��1�q�c�&�T�9t|�t��?I�N�[��(��z.�y�i��"��S��lM�'%5m�7��k���sk ��F`�,���/W&�����Ǟ�]a�����9��
�%ުv��(Цؽ%�*��A��r6�k��QOBv�������RR{~�:���RS�Wc/vɬ���]��f��l6X��3bF�i�
f��!�x�~��E���*�zg����
�Zc�E?)))p��b�vmM�:�W� ޶=�
@�X���܄�Z����B�9�:��6.�K0Ǎ1iQ��q*�zB�p�����$���=m���<P�mr�ie)"��{3?N	�6�<�sCW��<�m>ȝG�H\r��������j2��*O��/gq��x��|i ڼ&q��q1��G�8����5كg[m�6��>2��a��n��Рl8�b@�W��m=4�� �71$x�xj��̡���zՆ�����T�E|�F����Q�ky�&�˚����
&��h��D����:KRÏ'h�B�fqKK�����Ja!V�>O����B����15ܼ �m@�Scm�}s��* ;g���,�Pe�o}��1����l�t��F��)�:�V�Up��X�clTU5��������1?�O�9m��](�#�Ә�xS��	��C���������>��C�E�J� f	�8{|�2۝��	c�B��Ӵ>��r��_�b��~�M�M���[�/ �M�U�'�J�o�7��n�>�>6�B�D;�E�np���g��( g��r��X���(�0&�?.�5��e �$ǳ���5	j����e{�į���[���䅙T��@љ#��\&S����V.�Z��#.�E1�D'����n�.��l]�f���-����@��U�7��vb�п�տ���/�:i�ݫ-i͜i�,L�/�/!��T2Ԕ�~�0��+����j�0�@	]�I���i&��M)yV���������X��\~ZA�إ��O/���M�� �rcǼ ����:�tGi���@M�3�:t�o� �jx����Oя��=>ҽ���e�����k?�|MK ���c�E�,���sf�#��$��,3᥯����q	�w�l�~j��SЁ�İ�s��k%DUWX�8H6O��#�;�ނ�V���/���֠�m�=��3�s�G�bK����<���#)�lS���1/q>O�΢w��^�.F{�(&y�(8
�;ل.�'�S=�'ɻ�����_�Փ��Y��{~��D�Od�#{��A�'�h�`�r品x:�e�TYN�-��W�9�b��~u���`�sG�7��ԙ���!b�~&rC���V�n2s�l�[	22~��s���m����h�b�����������c�'��m����6�J�0�#m��{������:��c1�ۅq���$1����V��%`�0@��g6�d��J��Gm3LȟzʮX���lTH�ԢcU�[��sI����(O���@�Ҧ$EV^b{�}�Z��|������,�d7�#u�#D���7�������pj��5�L$�����M��׹G��θI�^�KJ�����ħұ@W��>u��^���w8�0]ؖ����}�����f`�k����Y?%���|�Z�|�p��02��
�X���CH���()7ǋbL�W�zi���i7z/؞!���X��WtNs�A��%�C�ſQe쭣���ϑ�E�7!��`��$�;*<Jz��"�ɏ&3&�]k][:�;;a�i�Ouҭ�=yQ&#m�'V��F��E[=���nP�B��>�c��8���JG ��
TEOͿ�~7���F_®X-�H;ؔ�R/Q.w	���k����֝=�����h<��Kd�tL/�Dڻ4���>�O�;�9>��߄��6� ���\ms+��%�Q�Q��M�B�tvQ
��?�A�y�w��I�O
�q�Y�a����nJ3�z�2��Ƅ�I�R�{�C�[9�-GK7USg�}{�����n�@F(���CTǒ�?�9�+�1�Y�����P��y{)��$�Yu�i@R����Az@���YE���!�F��_��_a0����r��GA:�TN/�${$p-�d�ǚ�镐X���%T��%ϴ�n�n���0�vϰ��=��'H�;����'�������S��8��6�����"��}K��GعaS9���Ȏy�Z�y �H1+Va�˧�d��|n�T*��-R `he|����88���q���x2�7�l+�/YjK�S8z,��� Ǿ�E��?�xB�����ޝeg�@I�gr�h�s�`Y��)-uYGm�v�'<���6Wh�!����	:S,l<��N����-���o�YH.��Nl�^G_lE����K��]$fՏ@����G�9�������:f����������������.1��O�[��Ϣࡳ7�%���g�-鿂��O^��������Cg��ȥW[��#*i ���%�4�\gXcy����W��)�h��j'Z�����FvE�'�2���"\RkA����]��f��U���2�GN�{��F5��n�-�y
[��\J��:�!�؛���ʌD ���Bq��n<�1�����Mbb@i��Ti�<��ʆ)��xa����Kk醰��p�22�۳Ytx�J�9om�k�����xr3v)��9�V`b��&=�Ͻ��rS�����ho�O`�d��$�ŕP!SBB5g��M�\�;�oJ���B%ަyOB�N��j�9��Ι�l���zz�q��ᱯ����]�f���M�,\��(����[\�� �ߊ6���I��8�!��v@�C����f{�Z٩�jS^:�p�(�M��lD��%�T'"���i�.W���ŧ�a�$5��FN��a�<Z��AQ7����W�U6��y�P�{g�J��S�<I%�.�L�	��m[��� Y�t8+v��zjx�ODK&�9�R�%W8Zy��(��V�@�Zr���c.�xܻ��iMa�6Z������S����"1&�5���� Xt|A8��j^1R��Nv8��A'����y>�4�_�\��Ο�$���vR�p����$�G=�2���ي��L���Ӑ�U��F-O@��KRZ:�3��ZD�]Tc������[���}���H7�
Ygt�1i���#��U,�6�o(#A\)l@P>���=��y���,3�@Oʨ*8!'2$6-ȣ3+/n��y�G1�+5��G�b}-�s ���8%	����(�����kH-��� ���{=5/�y��E�4�f�Z�n��t_Ҝ��LdD'�`hl�Ƃ+b-j����1IH�Zrc8�$�� ���D��h��:=�t5ޕ3��ܿ��*���{�[�U�:�3���p�|�e�!���b��qfZ8��[l����p[h^�՞Z���OL8c�(�A٫b3��KT�(����<^Oh)rD�!�IU�N�50�GK}��!ǕA#0�#�*�ܣ�Y�qj�B��b�J#���J�����̺?cn���\2U�ܽ$t(��dXu�J\gD�U�b��^۸:J6{���@�V}�!�����\Z�&$�i�8��r�E���'!<5B��"G!��L�Jj���DQY��mp�[\ީ���)~���=C^����I��(?&����[�s�-���+X�`Ƞ��
�V��=�V]:�dk�0ߩ���ܢ�f�n�T8:��ϟ�(��DQCp0n]�˧�s�?�2J`l��� Wd%� S0�k����:��-���Q�K�L�ƾz�:�Z��y^�h����6���.��>5X����F�QȔ6���K���E)Ցd��	5{��Da#I�.����Wj��ݼ�gTm3 ���67b�ec�牌���C#�wT�$LkZ���m�t�{�oW}���_�]R��m���5[&
�UT��h�D>�=��;�1��R�jC]+�XHEрG�c��_�Z~�����<��mɰ����9M̑SԌ��e�=(�+�W -��"b��EUZ|p�JB��4�#G��#��{
���5����p9t�A�#���F[�͝fR�
[f�eY�Q�����2 �,�ϸv��u��K��~V�H�����}��`GQ���	~��nɴ��|O�_\�9=��Џ
)9�ԭn@E��U�v#��r�&x#9����-e3�3V�:�s��̍�j�+�pp�n����w�1�e��")�-&�����-=z �q�q�[6]?t��y �;P4�����QK����a�р@��A����b�wҕAK�M���Xp�ů�:DH�[��˛5d�m��|Oh_9{���F��tBͶ=ߐ����Y��o֝���QL���*����$�v��x���&ݷ�d���}rչ�h��u��Kg�@����=Q�f0 F%u�Nٽ�����*�\A 	����\�k�<GhL���CF��\�cb�M�DH��0�5�jT3��n�����N��l�����"b�"'��'~��EҩQA�~�7�s�ξl�,���/��۩O����N�"�Rk�ͼ��>MC<�*7(X���'v��F}:S��'����F;
��{�J{�Z�P@�m�<�-�dĺ/�����ѩ�v��yH	�3�^�E.�Q�iT���N`q�{?�_�~�x��c��)9���ր�!3M���g�|!����B���UU�h�ȏ$�>�d�����@�x�+Hx��ک�5?:^�t�7����B1B���l.(㑸��l�ՇҀ����>��F4�(jb��{
�V�����G�R5[�k`D�am�TOa�UD_��.8�{���_�NS�U�A�y�]������/d�$V�R���(��v����F�M
P�T��8H�l�\)�b����;��K�ؔ�o�K�1H�*)^@y����+�1۞������}#mq��6�彣��Nj|���|��5^�ݹ�,Gq1�3u���|���9=򿽴��6k�2�D��r��]�a]��ܗ�w����fʢ��q����u=<oC����"(0g&Fd�]`��
J��w�P� ,��g<w�X�3��+L0�Us9{�w�ФD�B�-�}ů����}��L^zP����C���KZ�~C=v�[]X����o(����	��c��<�B4��R�ūd3^=�ft�mn����[�t�s2T�Wm�$�z~C�p�f鑹B��55��j��+�SJ�9>��ow3ek}>�H*��ה��0�������ߐ/�vI��Gv�N�/��x�	6}	�,r�C���k��zE
F�䷵,�W�a<��޽@|o���ph���/A�~1h;8�7�k[��,��ғ�d��?�4E@�%6%��*��
��l�r��Ch�8bG|�P|� �s֨�Р!�F �{�J�e�;�_�_���4:i��)�I	�U����Y����XN�?9D��,SO�d[�����(��w�	4X2~�G+�pen�Љ�1Q�E�R���jk��o�8��v'ċ�o��,x������l���ޢ�{^���']j\��Q�p�;"��g鯁��}A�����h�)��K;[%-�FU�(hm��ne��2DS���;P���c,�Z�%�r��T�d�h�8.� ��D�K�{Zy��3����2�b�0Z�D���DVMC�8�%�$L�\�L�h���kWrJ^�6����_�S���LZcTJ\��^�H�G	���?���t������DX8B��?D�1̥n���c�\�C���_���WmqiW�C҃�&�C��e}���ěHYf�h���H�p���-'`�Ȍ(Ql��h;��M�����*�`��	�8��|=ͻ����Yk�~��,p�M���!>-�GlIVY�����A_��L����R8����"1��6��R�y�P҉��l!!���Qć�^��d�ܲ��3�:2KdzU��X�ת�Jf_�X�����P�f�Uz|�
Y����H�o7g�Z�NŊ\�`n���Q#˯�ϡ���P�`Q�cxՠ��賀�ๆuo
[nT+T��ˠl;k|F��Il�Sb%�'�"tP�v�ZY7,
�T��!�H�k��bioL�*PPC�#���{����_'�9�&Z�P�� �L�;�M����v
�T��� rC:�X�����ۉ�&��I�6jq�3�Z�Խēb�����je����|��K\�^���T+�F;�B�r��������.>�E�8T����h��b|p_"��e׬<Y#0����&a�p���=�13�a��},���iHb��-��?͎�n�{���� .]ZK�қP�{��TG��Y�g	�0UJK�?h��Qy��d�l# �儺�o�)@Kbw�5�71N�mK��ˡ< �J�g�����V�soFE_}tM���^�~ͬ��KT��nh�Ƿޚʁ���8+� ۃrh�5Qa[�@��)�fr�����t[�v=7>�aVB���]�?��f�ng|B��#�9?z��OFF�Tį��4,��ѣ�(F��d���Ϲ�?����S� |�Z�~Xq�1m\�B U7S(��B'S�?A$���u����O�jJƣvl�S�<=����Iv��~8�p�.y�*F�a,V��CKkU��;
>���^VN=�Dƃ�Z�<�{J^Q\�"4�K�t+gCad8���0̙xn�oG�J����'��ff����ϔ�ӸQ��������qCtE�v�w"og(�y��t@�Dw�@�*y��p�g�-����m,�Dm��:]2w-�D��s��E�^I����q�8�|��M%��7^���'�$b"L�
F�H��%>���܄p�b�!���[n0�F��hqsOZ�oN�Wu�ּ����#z���u�@f��8�d�v�E%����r��$c䮕~:��&�w�a�:OY���u�|��e�"��r��F���,��[h�mP�&-A�Xjvȕj���}U���ɍ}[�{���4�ҟ�8:Y!�e%��A?U��T6$Q�9	wx���PV�)S�V�a������(�\�����������j��������.���Ҋ�W��fs=�:ݒd�d�k�+�G��YN���R��z!{�m��$�����{] Z��Χ�������`�.��,����W�wc�T��R�E o�m�M���ndXr��(�6��|�I��O�Jk9���:(�ђ�V��P�H�`�CѠ4��Ɠ�I��<�<��-�x5�]�/G�5�F	��,�j�d����:g�	�ﺤ��D��	ݳl���0�w
��Mr�����ت0�LKO�L�nU�b@�g��Y�H��@-���i�-C�����i9={���{��9៤s�D~�MY�����:�x3�����詯�#�����̞㇢�x�Z�aƵI��`�z����MK[���{�t��t9Ę�+P��N�W�
H*�*��b�Ɨ�I�/t����S�Q|�����϶�^] ��[cV�˨m��U�U��PRf�?�ґb��f�c����`�狮��kF�Y����*����~���U��R�XJ${��γ7�2_�h��oAi������u���O��`�c�4��a��{���o����f
i������ݫ����a�!����f���d�r��<��5uj���v�(DD�Vח;�d�y�gM�����<����;�hQ�:Tm�.L����%�s7�����$��[7�Pc�~������?�`^��2%�����o��եJ�	]��N0�I�N��"�D3��0���eo"�b1���R� R���+��=b�}{���x���.y�]h���5�b5,#�*l�aO$�`�l�������(>�w��KJڬXr�j\s{Im�w����r߅0��?t����V�!u��-���?+ģ��@jE��Vw�S�Y�� 5U����Z���o����[*0h� �
���Yܺŀ�\����##��O;,a��l�p.dY�
9��Q�F˞�I\u�%�������v���Q�]�W��F'Wӵ-�վ���X�8Vh�J�B� gJ������S�o���i\��!P�MgF�W��<a���v	���
�sԾ�]"lx%+8̛�(���F9���جW	�"��rWuC~s�$Z��+~9VF�(�BB��J��J�(t�A�˳<U�sYkq#z�D����-a�\�s��d�wZ=�
�iؙ4=�����9�6SH��K!Mʺ��gT��ȊC��������`-�T�w� Z��1�s�o��	�	F�ƞ"�W%�~������yV���	���m��
���̛=bky�����=��2���A�c��*dF;�t����%1uYi,	uX�QSI��ͱ�M�Z�����MA�|�o������9+�@o�Y��Rr�����*C�pWf���*�#�����vEA���ITs-Y�K\�>I��}#��u�e��'��D�tZ*���8_l*�y�g�mي�SL����F1\�w{�f>���a��ީY�Ճ'ŭF47=m�{w��4Z��Q+-��-�qC1����`/��aH;���r/�a�	*��0��R�j>�pĵ�( ����.#�w�{`h���I�XIH��1�c��D<�_v���h��C㶕z\F/k*��"��_�z!�g���������!r`�>����!�U#�&|���Ne�Z%�{�e; ���yP&�X�����s]�=�$����e���}�e�ݰ���{l͇f4�Ȓ��f�/�Wir��t`�H���]�	�k{�Y�u����/��G�2����&���M���m�VS6�Y��.��{���T0ޱiƻ����#5Ͽ��:+(����0V��XA�O��,�S�槐R��Rw���!�_���*�Ö��jk��,"&�HǏ��~M�Q�8��/X�W �I|�o�ΔM��1ͧ'΄��_� ��rg�߀��=��j���+�8���<qE��i�JZ�7
�X���Ĥ0���<�`���w�F ����M@�p�:�UC/bj){��[Dԭw�������&��5G�����F����k�8v�SM���3lp\Denl�r�[H)tn�5L���o|��1��}�	�p+U��8��(�BDq���ܠp$�����o��ePpڲ�	�NZQ$k����b�vD�N�Y{j_l4zYI�1��L�5���d��Kw m2��_�K㪂��kF�WE-���M��T7t�i�mb�Gٟ�/��(&J�;���|>�����|�Kjw�(���{�����6=3Q�!@��-���&��QM�����)9ѩ�1�E�u�8�äpJhC��zl3 �g$��0� ��6YC�$'+��w~��d���2�n7�^l����nz-$U:c�ę.q�/���}��_���*� $��]�F��h��#�MW>��88��e�x�a|�h���㚊{������������HL.���Y�4���0K�Έ��:�d ȘJ=N!EL���nA��@֯�I�ЖR �b��V|�0ˠ�d��1��2nf$%�͚׽4���C�og�T:#j�k�tA��~�Vѣ�~�R@=��M}Xn,X��w�^�n�=�Я�2(�|Z.N!t1�<0�%���ۇ(1=/�K.8�G(����Zl�T���l�T�7yr��Ȕ�=�T�s�-�P?MVk+ajﱸv�j�����+	Ũ���ᣄEɓɃ(��e����Ge׶��՞�+�䑈Sj_E)�?����&�U�~�+J�E	B!��*iK>����.],�Õ�9�~qk<�%�F>�ٽU�;4����\w��0P,���������a���>w���U5į�b%��L_YE�ݟ�*���%[ƔǛ�)Kc�Sհl�r���/?<�)T��B�^�3\�(�U�C]%�d݌��7%�/hQ$����yՔ��q��nT��[ ~���?oO�~#%�t��{���=�!U��:'����p�H��oM��e���@O�!g	��ݳM�L����<��m[O� ��F� G���2��2����[4!O[r�>hP�o?o�3�.���%�\��ݔTY��T���e���E�(�./r�7%�E ������|@2����)-dW+��)�R��\�쾃W�G��ts��4���	�޾�o��%�e��o�k��1�La5/��׆� EPd����Ԩ�y��@Q��E7�X��~Yfo!���kgz�E���&�č�&7��^O����Hj[M���{qn�o/GG
W1 1� ���q�/�	X�����֫/��U��礲�.�/F0�]�WښM9�A���@�,��O��Yi��`g�)�|0�j\���FD�_��v�(?"��f)>cD�1�]��M#�%�J���T~v��-�����:��zUy��-��Apՠ����-�@�
���f��
a�c����"ϿqZ�<�7�^�6>��\��-��N�M*�I(Eӹ��I��UIَ^Ѩ�7��<�
��M����6_�L���6�)|��8�V�:0� ��ZL��>t�!%��0�Ӯ(F��ǚ3i��u30#<��8%�m�#Yt��"l?�|DeV;�	�&8��:BFy�����c7�p����$À����P<	����0t���~L�b�a��o`�����K�b�t��-�%
���}o�L���t �*>m��'U��S~�"����Kh-�$�P��tȬ(Mh����]�jj����:����Z`��ʻD���7
��fh^4&v[F�.W�S�=��¯l^xY�^�uQABX[�$�^�%���Co��X�*��Ʒ�N�]���#���8��'z�X�c�����%|6��0�l��e��gzP/W�
iP6�k�r�{0�-f��DI�L�RP����g���^����j�cG�מ6R�C1WHRy��}�r3b5�Wv_�������asff�<��a��d*��/j�L����A^�(�9���We��N{˚@&c�ɝ6I��R�:y;�nC�J�*���U��� ��lԂ>ː�V�?��	-frc��w�13m�%x�v�M����a��y�����n�~��`�����X����ƍ�+v��k���/���3Ѕ��-����7�Z��P��<A���]��ˀ,�'���i�ӫ.��b�Rev�0����R��C��N헭�~�ż�7"X� -�#�KE���a�����R�6D��3�?�!�ІHv��Ĳo^
�h \�:Ŗ���+���NT�w������*b�k�$�a��_Ց��]�n���{��`�K����H���휴m�\�50���ǝ�1F�`_&�`2(So�,<������I��kd5e��N1ӈJ�9���3.4�Zn�Ԏ"�M��P X p��"���Kbu��(&�ν�a�α-V� o�]��$�朁�����&5s��t��~�u�[��,ۖ���
�l��ȊʾD��� ��Dr�?�*"2�3p�@ɒ��{#��+�氵P����倿�6�6J���T|�[%�#�c�
���%�
 1q��I�́X�Ė��2�T�H�͌6�aʅe�=��@�A�]&�RILf]O��{����Q�8�Wݠ��T/�ۆW���p�|%ŇC�5�5q�k�������<�P�O��6���~�a�M��~�V���X	����)��֭m�<�dȬ	γW�P��,��o�����Ԯ+���1��	�.7�^\O�k�r�n^_OH'_{�s�G ���cR�
'[�g ����dN_ʧ^�1���,��2f�|��������+�|c��#i`�q�u�!���4���1�Q5�A#(w�xq�|����Z��^�*�>����ڬ��AP=}aCAo�!&�׮�<*-��/9�Q���|��Ñ��-=�r�qs�U|.��'�ú���!�*�ӽ8L^Ja4-n�LkWy�e��g9���Ϸ�4�F�[\.��9��Fo[W+��Xw��fҩqG��AJ	X~��,�B�YoF �Y%�ڢ�L�����oIb/ܡTK�u^�?K�<����Y�Aj�VV��Ȣm���Y��H��Jz���3��]aN����e�P�Z�v�d'J_z���j�۠��W�~"� �o(h�:W�˚I�����%\�~�����?Qk��;�m:8]f+�!�^|�����J�Ҁ�8�6������|�%�����Vm�&�/�l�|�,��������޺+2����J����ۂ-�,�k���;���^��Z}�q�t�2�J�6�1�kaj�/}��M}�*�����[e�E�����Y���W��9��A���F��df�!��*˱��|9���f��~�7�ɭq|���)�v������*T)
w�W-d� �&\GU��dj{��F�!Pĝt�{[U�J$��lVۛr|�z{
Ba�\���?y�bgk��һU>"��2Ӟ�a�Ќz�'!bk��*w#p?XÐ�'n�j�]6�b���0XA����:2�3h�#�qN"�cA�O���-����*�_��M�1�5�q�ُV��h;ȃ%���;7Ku�Y2�U� ������b�˴I˰��]��/�h巺�\(W`��i� ��XkQ��u�rKb��"ծ�4����h]U*	����Hֆ�d6VVaf&�=�b}�9��e7�-�#b;l���k�<������U#��^�ze(z���C��r����@N�)��%��J.G0|�=hF�CQ��ju'���Xۍ���%��)�ƌ���ۜ����17w��	4XAL�:<��V�C�����*����Z+xָ���>�2���܁���j�˂x��|T�}Ϋ��o6��6�(쉮���܊;�'���G����O��RuP�j6C��Z���5u��}7Bt� /)��KU&\�bX�'#�9�OtK"���9��%S��Yen-����+h�E�L^����=���0X�2��'Z&��%$x�.�gj��M8rjah_�:~��OX9�7���5��] oȢ�H��źg<��m��s  f�>���.V�V�l$��:m(��$�W��Bdت�~I�r��La�d�؋� y����b�o2����($����QS����{�P�(B�p2r�@��c��0���<"O,/�d��Z�;"1�7��}C@9'͐�.���&;6�'��r���zF�����0O��*�bBsy���x+�ʖmG,�8%��Bs{��U�j�y ��gm����7��,^�G�7����Ji����O���
�$�I��W�����qn��-Y���A�d��$q~��C�������O+���eE�[�a$t��Q?�m"��`峆Y%�v�B�`�T�K��Wh{�w�}!���ֳ.��c�63W
r#�5���@iH��-��Z�胋:u�4�6��H-W��N3�2ؠ�K��8�Q�#��\8?�<����h������=BԜ�?����B#z{����$+l �?���_�H�6b-̪���w.�����P�Yg	��XbXW�g�)���wU�;@���wU���G�	p�?;��h%]��|m��!�.Q�H�Ō*^�0�;}k�"��׿�s{D�4%��c0��l�c.2������"������	�Z#�ɪ�|l�F����+��ts$�����/�A;��B���h�#� ��pD�>�vA]]�ád|E��o��V�Q^��od�ץJ (L��)|���j:B����*4F���*�|.]l�h�3��Gg��3t�
g���d?(�Y�CX|�ž��k�V�hd���
���:{r��
����6$w��ʀ�+&F�dE�>W�B���j�*.g~`��|��sW�7|e�r��h�0EE�ޏyy�F�i	�퓊k��)����C� ��a��v|$���9q	�<{J=����fj�]Xv7��-y>ЏR�PR�{I��jH��R��tb��~V��.��~���]Ya=��*S����Ϩ�o�%q�78�[��V�� ����8�z�
��n�ow�)�ٟ�>��Eq�`�W2+�5�V��}�)�'3ČuT!Q����i�o�h+����ʒ�������-.&9�j�������a���4��t	c�F���r��7�]�{�Ӷ����޹	�U��C85\Z�dv0m��<xm�;����\�-�ܭ>��� ^�l��,��@�/�UT3p���\�.��UѮݐ-��׀�1F3|��"�?}��̾ځ�����"ǝ���
t�B�!^�6e
ZP�!��x+"������#{,�����l���p�N�[q�um:��(�~s�no�較���/a�R�>�2GdD�b�.e�!���`���7�ֽKT\�~/b${ψKw����>�}	b�θ4�x:"?�^^�*r��堜���v�uXy�o?4�n� +��=�m���x�dlR�}�CM�����2��"'����IQ��(TO7X�]lz_��C�	�C�r��%������e%�&���a���I�j���CYB�?�����-ָ����a�� .��om,w0l�r�����uzb%X�3��/�W�I�@��5o�|��a�Z�E.+R>1"�P�$'��+~΅6�w�#��˔�v,x!�S:,��$��U����*eW��y�H�(�ĸ���N��v����Ľ?�I>V�.����#:�F�D�Qng�f`�9W�ټp��ݵ��0*������ލ��iSq����(%�Z=��-�
�D��T�]��~D�)*~q��պ�d.I*1�M����7�夑�0���r3h�B:B^ �G9��iBbM}b®˿����aU����Q�>�gHx~v���m9���Ύ��ʾ�87�5Go����"2�|�DGG&0�G����W�Ӹ�]�L�f~lImЩPs =Ӡ�	�i����(x�P_D�53�z���b`�*�9 ǥ�gxhjω1�C�ohv�O��m��栯�6U]��Y ~T(��M�(E��q%���F��י}���
�E�'[�;Aϩ���j�uЅ�W�)��_E&��=,�æ�cI�	���y�?��ַ�l��<mS����Q`6!�Υ���Ǻ~hu�QO����I�=ժid{0c�QV11�81>�r� -���!�He�8&��eb���D�5��9��b��Ŗbĺ���^�KJX-T�P�x7�k#n��(�Rh��b��N�&%Ȅ����\��!m���*��L/�Ů�$P��SJ���Yo�=��~*�fY�j��T��D�����߷�����Gz�:Ҙ�%�`�\��1}����|K)���8�|�A&PځI��@Ӳy+%E������9�o�w���V�SFg�%���W�.�̨�������޿�6�����C��B�J�-C�7�#e�AV��JT��h]?��_ ,��xN��6���������σx����>�@:�ڃ�0�{��@<��Q<��p�.$� )A�r��"��̑�L7�S@=q�2��J�8zM*aߦ�qn6� ��W�?�:V:�g���ABJ}�@m�O��?y�:�V��2�Xu�''X5X|Q�J� �b_�l��8��E7�Hf��-W�(��hE>?Q-1��#��v��w7��Zď�q2�޿ M�5��v�u�w(�\��G��\�1�r���cFS�
ے��/O4�اZ�WK�¯�@��C�M��]��q1j!��b�҃�DT'�k�� }��?�ɺ�+ 0o�o]Yo�f�� �]�MP�:E��z~�O��kS�H�Eݙ�'����0a�]d"�-Ŭ8~��w�?̭yRg C�ur}_���>}e��K�;n��T�D��)q���[�_�B�[��Z�qGu9CK��v�D�ql4�	�l���� u��K ���Šr���Κ��d�%qJ��Jj�?�zm:K~�H�kГD7$���k��1�2g0�T�n-e.��`���S3�J���p�q:���!V���3'�)W3��CF���<�"��a���wQ���>K��|��������I�����������lS�!<��e�;hQ�[�dߌ��ϺLϿP��SOMK����R�R���>��o1RcS���-��גH�t)h�1	�wӋ������i�r� �h��p4�Dg*U])X��e�[Կ~��f�N�(An����};drui����b�=�"~��_��N4ٕ'�:����=lBˈ�\6�����4b��Ϸ���=�cx����YŨ������Ȝ���1w���=�� �Bɦ~��n��Չ.�.�!�+��XДx�S�X�(�>��SSv_��l��C��>��v\r���>�궳��D
��q7��������p�V�K��H�n+z���o0�J`_}�t�\����b#�2\u$l����Cƀ�o)`t6�u�* W�r��P��=Ԁ�a92�]r̝e?�ӏV��d&�j/��ψ�z���,��?�\~#NDq�hi�S�,Y�������*!'����H@�5����Y��mGPR>u9�r8%�s�Ⱦ��B,�rQw��a{��	��oui��}H�=�0Ȝ;�\�N��k��cV�������m�Z��o"A4�����/��	Я@i�b��U�!Oފ�끪�iڢNL�jӺ9��b�\|��
T��p�kr_���
����J=�=a������d=�{l�t��ק�);�lG!�=�X��s2�(�U�W��!^ѰwZ2�{U8���d�2׼`Wk_t�d%������δ��o�>o.J- �TO�s�((�c�7� ��⢭��y|��@�y�2�|.e�P}C�X	]�@��ڜ�F
<j�G}xD�u�|mP�)��H_o�,l�������w�fj����s��m߫�����?�t�A���������h�K�}G���4F4p��j�7(�Z�������B|ثz�]��	Ÿ*�>��;��25����S�nU�]���/�6��w5i�>���_����'�C䦇Zpl՗��1���y܈n�r���sA���KqD�1�kesٵP��A	����*8ϊ�T�kk��{�8�a��~y�R�����S~�d�8��
�o_��s�Y���m2�a�9�8Pn�����F�Q�k|N�OL�Q�0
����ӅKݾ��d�;:a�|{�;0K r3	c��]�H�`r-1�`��k�	�CG>H�%H0�}^(�ɜ�u��g,
�x�,g��7ԴL��d�؊�N]*��c!��h��_��p۰�MM3{��o�ID�Ĉ6^�dεu��0�E���(���N��	yb��1�39&(P
6Y��������MN fC�Ʒ���܀��$��0�9�K
Yb��i@�����g�]���㙷nKzn�ixN��j�"�c�[ll"���V���P�f�r�?^��D�\�7S�ME�n�_e��i���$����jY�R����m��Ӄ}y(���3��(�] ~(�_��^���M�yv4e�; {�N�~�ӕq��%�-�;�y���3��`�?
a)�ʓ7�K�����8`}����*�����2����c���������95�=(�r È���'$OA�# ��N��O'�^Y
[_>���i�H���%,H����"Q���O���dO�x���z���p!	��Z�D�m�I�էμ�/�7�����!Ŏ��b5h�v��,��tb����'����/_�FvdY��O��h���K(	4%�9A�P��}��$��vfKi3	-��3�!x:[�#_���IB��Nod%R�~���g�vWt$��X�7I�ا�.Wv�� �ULihz�
YA��=��>����=�Dσ���7窾q�l���h]��R����Ϭ�-���(��B�)�ٮ���ԣ_��Y����)M�6��z�C	ۣ���A���!9�Ւ��΢O��Puc��%��f�����_V�z�졊�wn��e�����C�L@����(I��~��&f^����3�՗��rV��i=@yg�l��s_`v��fxL�"I $8�	��FH�{%e�VĲD|���*�����4y�����=柎�ԱE#E#ypq;�������R�)]	i�D��������"|�lZ�x׺���4pTTY�ݑ��Z�.��8~�ە�v�M�2��.E�@�ӵ
���3��C�~~m���E:=V�fǎ�qO0VE��X=|��=K�����9Ё6��m�WK�"�:R�b��t0�v�
���$�R� ���Ӡ�/�a�g WwuČ��;��g�G�ď�Dl��z�f	k�pEm[:7�_Vy���a��)Z���:p��&�����
g��*����bk������u�=�{`�`�@��+�nW�������-M��DZ����hKZ 7��� 7$�7�<�.ߓu��&Q�-��e�/�a������VD�y�AD�������z�8���6�2K�#��o�������(5,f-S�0N/�c
�f@��l�dG�{r��%����y������~uݤ��f3���l�_Ψ��1\]�c�P��R���̀|#���B��_"t�H �����*@���a����o�h�(��\$ހ�ܔi]����lC�-Dm�rn+���GN�n-��*�9"
Y�.]�G�˹,��.�<�먒Q#䀌�"agE��S�6pE���u�7iJ��mC�n����� mI���:<����՗����OCX��w�����8��V_��wCz�7
�����wD2�p�H06�]$ڹ�����`2<n�#z����Z�h?�K�5�#ɩޜ��<�X|3�E�#���3��Y�[5/3\鸐�������H��-Gj����اZ[�5v��g�:AE.����x�2MW"���� s���	�� �?�\hdғ=�;�~�������y�)v(��A0��ϩT\9 3�̓.k����[�p��O���qy�i�]���4s��X1�l�E� '˔�
� �$��L-I�� i��t��ڏ�R	�=9��#~�}'}�U;;B����k�i��2�E_Z��n�dD�L|)w�l�%�<���{���z�B��#j��m�낗�c��g��s��`l�Ӭ�$R�T��Q�3qG�z���\�ܼ�FD{X@�R���<|��{zCj��?fkiÇ��h�!�G�^�ϻ���4ڷ�\���zağvO�-	�c���#Qć�*Z̧_Iut�"��J%3���!Oۆîѧ�=PڈH��A$��