`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
gYDYuPO2G/aEJ1cNsG+xVzWQTAe+ryXDfqdtwPbzSKHHLwS+Uz390VgHomsTesEs/zREQTOHU0Rq
O7x74OTHYGg7I8XKSW5bDUsK9v34lbdv4CnN9yS5ywYqQE8l+n3hcxQNXGyenYaqnNH1Ubrbz9Wh
y+bA9+pds+UlOb+xaNdcS6WQcrXpmJ3PBFQOGwSBQyKOuTNLe5qgpoNJkuibb3LLfUS7JU+0ir8o
Q8bYZaNlI/rV10tj8aw24HJEGDSMB7VqkbP09cjzHTQChEt9F9kxQl4QTg4kTxNlvy6XixcJbT5J
6cNXHEUBcIEET+t4sIHaW/cM2FF8RFiyyBdB5w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="PGOM+O0o0t4ZWOOva/QU9Yn3LmFTVbvnZ17oaHoRIm0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13856)
`protect data_block
piSg5O3zMxPRFqxUOVt/7FXHIJ8/Kuyg0IZukb1DMENnkPq2M0Hl5SWjytiars4527VM3EjXZPi0
233KLZ4JiA0TpxHTD/cWW66zdWCPCNmCISocvYp0W/ejtxV2RiPyRHPpNreWLKkBffm5/gVo4c7x
I8zfjRiFUaommo6iAcIxbdM7SvvOjEuDocUnYYJoj6/ejuLgDmiBI8L71F4RSWzoZbru5gvzZFLj
WSq1Rv/J839dILutAlu30M3TcTjBIhmev0PfnRhaUWly2aZ7QpVwtG2Wkm42VyhiOYatQoyeQGZ/
o3jtPuUjf+1vWZQw1mPcsZtwcX25ktOcSf4retkGTPS0aDrFsioXCRMEQs5IZ/2PMIF6I+nBYeOI
s7/+6Saifaw4sTvLgOjtGToo7mjuy4lbamEcPD0xwYtccQ3tUnsFoPalpuYRxstoFIYZdB0NCwFY
99P3o8OXJ1v1TToHb76UVUApOjvfbgTY6sQyHeypzc4s8wa8n6O1Afy/UDPC5+d5EwAEz6Y4jslm
4hEx44Y1rfcAIw9AXPQy1pGk7eiI5S4s9gGxNdCHr7YcZHdomoK0wAMYvbna3rh32g0+dio+CtI+
ItEqICPaMn4QlzvrV5bNNQlUGkwc6ZrACMCugLLSx0KpObkl0Cpi4b34I+TjUzVRgyO137Kk+a98
laffo77wYj7IYjZrAixT90yD04nCS5UCZI6B49UVjn2/sdn9cho8CaXwZxjRIZVDBmjLXROfVOGK
hKQFycbOMc8cNwZLDK1uem5TNUa7lPsL0dDsmlGn3G9gInJmA/j3+1h2GgMjN33qifu+Rd/wIt6z
q4jOM1Ast4r3bE0unskz6IwXlUZqVBZbSRaFEhVdxa7viFLnZY0V+o4xvIl3Uuh9rTWm8WYCBNc2
Q1YWeimuTQyp0TCOvDmY7yz1CVHNuvR17yFu3pvefxZ6jE/cc+1Rq430wh/a7TfM3+yVZkBuqmfY
HnFzpq7XlfrrOq+uesQiQPLM0vHGmyG3VnN70E+baqQ8lJD15wNmeWCAEn6VTg/hrMXtUIoJqIx9
H+uZN5YQqKoVrBkg+vYTvtnTZvYTLyZ9C/MpNOaTf2VXLuuRO2pNKv+Z2achTuasWZOFwoy7d28e
0CTUvZtptnMMcS3vAQq975+ISp7nf8a/KQUd3TEftTEuvIhJZcF3g2ZyCuP8xtDoxFAe3UkVFQyf
buvTdn8z/OEPN/zC8vxlBR9ZgrNWqZm8mgpwwXii3QJhBxVEcgO0/X++K9L/eaAnYr8ei9+auI0l
fYsNVqi/4+m4XFmVNJGNfBgEUeGSfBrljOYi6Q/ncakdWEeWAPRuK1Ts+j7yZzFcI/NE0p1slN+w
pNJkh5bz9if4wuKn+xmD2SofwEqBIAju4lDCZ0dQfhOEDdfBtWM2v9B9NTgyy3QjMzE2Zv1Hhdno
2zZSu6bP6mgvliVJoeDkAnsSYoRJbXzt7HCJmGShgAMaTGaSSPp55OeIRGgf+PQNlTW+2b+M/4da
M0QD0p7jYwepvz70526m1FQtqIBUtf+ZTnHldRDeyVyfwWjv1U+uJ/ysTsGCiRER5kbCHpiSQlwR
cCBmDL4QbIopbWzpbd6h+LF9uqc3SRvkc45wzhbOJqsWGpOz6ewshcZfNP0/+990nZx80nAGLnu6
Xs/VRNRauzRDb9qArr16VFbj1Atn5JPTIsy0RAfjIxd0iHgFPl2xdHyF6CSi0Z0FXEcdgVDx8DtJ
YX/u+IvgaxLPQxRtKH8xAegbTsbBuXXsTotLqEdprn95VYgJDn5BI2EQK8DjbRvxflKakceh/i3Q
JBxmLjgBi42l8VatIxvx8jikDyqtcOXyAwrbz2sLIMwRoxWV2gRQBdv1NeKZTq2mTj0BlJY/0Upp
hBalodwSz1muoIM28Zh9gYfi2kHbWT/s8YMECJKsCA5TBHtKeiIplxi/PvEBHSmrT2Y+UySkVqiX
+A2pcL0HBkU1ewB8lmNFfe7HYb/eAMcTqqKnLRUCs+W/kH9gAihOQhEtJnMKPTOY6INfCkbGng+Q
C9UJvRuhDUz6fJJ0TOpKVRjgVPQoPVjXbTrgcziOyJcQ4eD+KiaPMEcGx62bHgjxZv62HFzYfq6m
b2GzyFBfFrzFelKJi+QrgdwpnPCi5CcrQp+SpDWuFNxStMkGwmDHU5K/owie3U6Vp+xMK5s3qziG
U1hj8nUuSNT1TMXR7RB9I3PzIfe5jMKSgtMF85udoXJoa7JMdgQR+t75zQNjMSaPd0MhRbM5oCrn
c70jmteIkjy32+JpOy1i+m4feUPXUEFarc6xhbwPYNsfTVYXhS7U7+BoFsiBN4zRwwWmJrrCuUhP
E3eZguoHG/sog76ga+h4VJYsutlJUmkctIWxwKcPqR+eY545Dzt1oq23qf2V94qii5mxV1YAo3dp
dwwz3RAVcps/FCbuTXQP8tmKQf66QUfmW/fajp3xC055OI1BzPBE7KX322GT1HIX/Y9qggxASU4E
SBfmiE5alBEmXVLuNCqiVzS5DHZyBgPSZfzlrxdQuhVAnlJSaGhyXXhNXm6yoflcv2IGA/SxelVZ
NTg9AryBL3qcQEKl8qwcye758bImCAp2rCljTQXg+2Iual05k4ZNH0DGFD0RTmIqBibIhDan8M/2
DHTsSfd4OObK67nYwjwu71sp0XtXI+Pjjin0mZFBCKBgs8LQUAXGDkLfN9Ba8Ziy/B7XzmIW/Uru
F9fwvyfvA4nfsB/z7l/B1FI5Tg4ec/jwocopQO4bbYcEK3D13Vv8PTiZLGnbWGJbUSw0jqV2lNen
a/nmCxM0tFSR+edghKE+6eqqA/nRXO7KX0mKuQ3S/AxDcZkAIAXSYWmvsp03CHfGi6iASz5PW93C
FdQM4h1jM7S//uGixdMWe7ya/z2tCB0juY4SiNCPKhqusyzaP5Ko7djujxLCyCevDgJhjMZWrqzm
wQtGC4KMzTedGTkimdzpxHT4tMbTFsLFOm1zWdIC5sSzjTCOYd/llxG04PcckDT68ru5zVwcswGO
ECrsqU+pExZPuMl0vzwKVKlx91RIS7WfzAgmp9otbdmJGKEa0heIDjQkJ2TMF5Flz8sdBl7zLd7Y
jl7yzUCT5Nt25IZ80DLrC/jhFCwb0WZRqYU5lJmliLeFX4tQJNE1USLLMSC9v2Joevu9/al2nsDs
ukWO6sn+5cgR8ZKkG8Kb7GxJiNeaK9vymIxJcbingWDmJElBCVjSmPnrehl3C2zhUNZFmGSrnY8P
SRsUzxlHaFeopUUhakNVpNVbGiuLwM5kecXC5PX0U+UJgH1VHeHFZV6gsoFWX8Y10VLGqUogmQce
MgZip7ALUIcp+nSRVxaVkatkc6H5LJgmPZgCA1FRHbNXZSPr6tQLpImVWO8xio2Kb1WcoB7xOtXJ
6gNQvSBrisnMTQHCf6GZ4apQeTPZmp5MzeS8/l51TLd4G5O7e7wIT5zBCLuigB7zrAets7vvt8PD
lP45lcxdSSQBur0dH7T59obJ55Y+oQfUhJpTEk9JjqvUqxsXctYn1OjGu9qLvA5W4y0fg20l5z+E
OFWcPwGoqFQbyQhrpMRbfaolfRRIBHXEfe72yUslMVKRrCMR5O5wvWxHfiVGJlOeUqyurbFCPk7E
ZXwmcwR8JP0uNNxD9Ymk6NNmaH7jaIkPZXGOAjKjcgZ5Ocrf9/yp8PZYXqFN9FUpHTXFJg6tTtyb
nGVyWxPZX+FfX+P0QwcWoKrXyBwRRKKd3HskDCBr8QaBvOBytCK12sf7x3Hc20bA9IlUteoYQFcz
Tl9h9QefET2R9+UcDszknSp37rYWcrp5SpBZdiA0zUH2nRgHiVDju+wqKkm1iAJx+j1bpCoo5dMS
gLzE6Yx9E6xT68UuzCkz1UoPHk+Uz/md82lY8foZO7ZbB7gDOQrXMLDbmtKqcb6G7V8VYHVn0Nz/
h9ThT9NMHP2dQMpJ1Fq/8g9UoFwuarpWdEmx8Tj2/DTC16+vtlw7HmMZgz3Sij4W7OcCvJf0N8Fi
uDYYFyg8YR8ePPVC5Pdo0VoyvgusA4X0jF5P93SZDoDjjM3thhHi+XHDVGD64NhVc9opUT2yRcLs
5DeRWu60QIUhR8LbwmkegWLcplzrgVjY9sGVaMqtfIZM37e7ygfZE5ikrNJBL7XwBXDLsp4WtBhS
/tF/CCS45vVOuoaqYAIPJzdSTG4/5M8BKu4pMFtrWz4wYVpoPdOriTC3TdBchy7qs4rIdDKJqe77
dSD6BqhMycD+kUl5s1EWGgxo01TmKOzMJhk8x4TO+iqXgma71yO6L5ZSY6GC7PNmq+odjdEZYu7G
EOtSBEcWb83IWo7oYGD6NhvrBOqzGXRiuM/IRchshNRXw7h/47X/ls55FbIWMf8clXh3U3I8+9p2
xnFaP+prEXwjGReOUk/21z1kpEw1kpAozilQwNf0OFwr5mkdSLbX++8eCDx9VUgcgs6YClodoT5b
USh2ZMKic06X9z9Pnv2utE4lg1/wN3OGCp8+kx0erB4lRSQlp8iywRMyVqY5hrBYvLYoDS+MjaVZ
UYj2jjVzbWiXbnEMDiTh5G7rqZyIr4vhWTioRfCtjDdIg8Taw7NMdSkQXsfYBvlu/qQzNy3te9oh
JVHQDhZDBmzhCc/Gmi7jxnoudtdnRFIW2FZC1LqdTtNla+s0EtmrwefzS+4dWzR8xSyZGvaDngFk
VVbqKfPc0hS87kgYcMxfdbY5BiqRpSrqjU10xPX+mdN9D/rDcVeTb+pPKtZBiK2L16j8tDTbRGku
8SdF5CLx0VPE5RyhtG+EC4PBATfF9BRjz8eyfi3eqIj9D5r5tCaxafnNuDdmW04w+1bh6W4HXmZP
NcaNvK5aVVwdtdhmLGcKgwYe1kkuzeomitTomgokcyorRRHcGSukp1aUvCltKhjShO2khaAupxio
YV1A3EJ1QAg7yqFV2ZfR6GVZxZ5YGRm0xUz/MOVTQdrsgar0WriYlkZXnHbA0bK3bDIW3xJkvZZI
l0/4O2ShEWVF4JK7yNQUmgT2zSvpsqi465ETBgJPIbugDXukeZ+SlrAQotCykHDF9H1b7AwTJOnc
dWXr6MOvyZckWUJ/YFikAbAAqiIP7yDJrnOvxyC0m+qtfBrBJtc7ZJ7krX8uliEaLAkwIJ3f3x7x
F2BuMIo4TC1PjLG7TWcpy5Df7rFuJMGdIDs0Nzvm8Q8aJvzlKOblN5gTH6RLZRMInFFvm7zhDvlI
DITKKqKL3V5GPSlOEesrxVOvwViQfjdypLSyXG1e1f20Ehz/GxhH+dDWuRp0Lo2a174z6YVwaYRt
CZpjigQPIvAIjM/Mm77cyqgJFmqnffcS0Zs3/Drm/lcHjhb/AkPW8EVXuKylTvZLtcyJcLKSx71I
f3aRlf9ZVUN7CNeDCxppAQWmHbwLx0iXSxqHe318niEVdU8Es5CPtkasAkwrxRawbO1ADyYEOvBf
vw9OCiAlb5vMONxHzxCS+4vXePZiEi8CUYvR0LVATzaLQt0+WgZ/rLuNw3ttNYN8bQx0N/pPFKqK
9UVBmIVFJ/AHKR0v0T05jQVUCD2RJuemo8vJrtwYlxq4HZJ2QvMy1pTafZfJ7EpJzYCaq4XsMdFz
bIo5aXQ9e87jcxLsWjhv+9gH0yAs/zAHEZe+mn61zq+cPqj+oX/18ijNW/AiseMSsCgAWctd5rdE
uvnORbYTirR3gNUfOXWGWit3iNdYZ4AGJ/Mbexq03Y4gg1n98Tl6BErFi7143kL8e+DNg4vc+y8d
xoMP9AB2KMZrVdeXTkwls5OsZcozRAkL3VLdvmC27QB3v0L+AA7zU5ALYkm7M87Tj4+GMnk7k9GO
G8mF9ehSc1ZQ8irKU7yYArIXPPNknKJcYfSZZ1w2HU0YIeClgnDkCvVo6YZYDLdGuD7xoa2/3po3
6mPquMpu6j4Veg41mS+4BEEJm+LIikl5P+M6jg1DMYzJbQDKGjDDiPqeAc8szWIGEAQwckEB3dhA
YU4NChKntmzhKXm1Wff83sAnaFTTmvjguq9quR5lxrEgVwmcRMj3cDrkYYEcEP4KjejpiCEMMjVR
Ym/9sxoDnUj6G5iyMgrTmZ7ytDNXw9svCxjyBURbUcYHZF8ze8tLx7IwGtjShWaVyusp1zx2APSA
+Q5Y/C1dXN2VHkOmOgbgkBxlchT3edkrs/PWjSNQ9I6rX6xtUPHS3jP5D+1dzsiwBLxGhxhH6XNY
OkD8lMkOhYaKIhdDrAm1E/PePNsAIJ1dO7PhvjAy2kNrKhoxhKs/MX3fAbM8jHIS+QT2zJ9rdAMn
r3Yk9qW/DD7DAqsq4Og4hXUG99hFNcjyG/Gn7a8t/4dAaJWC2t2uVFoijMFHLw6YAi7OAeNNqbya
jABW4c3o7gX/ynDMlJmwG3qmkm9ErYjJHEik5tvUex5eLAiV0Nh+a1fLzlso5jz3Ulpq8BuKY0h8
fIvdhdn9pJo+ihvlo4XO/LRY9yCoxnlVgWsUh90Y2SwElYx16QHq2lzuprmFCQUi4IpinjRmoOMd
Z/pOLFYdMKdVz2iNqHSI/HRjAVhlgf6JMkD2x/bes9jzfSa3WOi323wXidb81gjy+LNLqmzHXIi/
fzNRE+H4NeMvsDLedF7JfxImlM6qTRrsbU/q4wT6b36PBpRGHPio2q3lmpBHZiKoQVFlDAr4eyI/
0unHizeGZkOCbNwSTO4ubtM3GWKsb3qvzXGl/bZ1tSOjYsp0P4rpMr1dh9Q3YeHRxo9FRPORp3Oc
nIDc0EogrmpwxBzpbJVINWQLWDcGkrzMQOJ6bBgKeTXn2f/f1OXki8dHssn9zXPpXNSvvhWf7D3s
rPjJ1LvoXMqRYMQRQIbOHy/piT2jQh5Jzxbj+lGRuzhv83TPmS7T+NJmm+xWAs9Pr+HcqwFp1EIg
5LUNcbVq0FlxiJLnmCbDVGTND+fNZ3/hr8x7dy1Q/Nm8yjWu9mMDZ5ks3EZMbLlGdkSQGfedPc/w
S2xdlTgBX7ukQHAf5g1/ffXvYApBfoWW1d/u0MlzFJ8iBzf22w8RFNgz9WL5uMwZfxiaclyCVSYz
QKYJprJCl2INmYa6RCoZcojgVfnqvPpqtPdJFs3g75R9FSkzLQfhpuzFrFW5XkD3uWOokTaUCevs
Cp09beyMHYn/bq5vl5NlwbjqJ9MvKoVlnWLAngPxxgTCQHuONWSpXfAEdw/H+Z1DbyKMhUhImF4J
3sjsbIb0QR6aN6/7oxaDKhEiPfixzpcjigG8p9OCnTdKyXZE6rSQreyA132HWP03dANZVbWi/q1a
z2F2zC6VDWfV7K9wmVAyVvFQQey4s9P95vFuIXixwq1SZOgHN4hKFPTzN2uAdazEnc1jMlco2RGC
+WwobOgezdh+/9D/ath/HbRQWFMYgm3pEKR9vZn9epmZSYP0/+VZcuncA/zyy3+A4JovbriNzPdk
uLYgGJqhqAiJ/8+dDz9PyYTMNHWVOhc3aMbTSxAWsIYyczcmrSpWm3rYW7WoewGj+bvpstMz/TFk
PpPj03xY8gHG/HpQDBoYHsJ7UlHeFTfhSqGIijmCiiBeDgBt7A/VH0R9rFxIoJ/0BfhLyB7jc9GI
8U1VCyYktQheBoq3nXZ5kd3UMGqe29RTAOl2btIEiy00RVDi7TAkkJ9WVRLQbPYeL/pd5m7OG2nP
wgoLnwWj9nr4Qn5fWrj6S9lg5w8R8ACW2i9jrf3uYVz+ecpLSU9w/rE3fYizTKU4zvKdOUBGcJi8
Vy3yjQL6M257feFCfnlDARAmgYE8z+9bM4AYiLpzEXofVFVoEQMULATp0bRid31msw7cD9nDnkKn
daB+Mux8wGQ2+ixqkBRBZ4erV/Fj60Dfg9P7Is5D88MvHV/UdDuS03rGwdGHaDZbIzR78YjBJuLl
OqL7qZikrcKLby64HVAqbF6MhDHP/vLfkCnA4MHKmJl+SsHUbl28xMlh3SPzqpetUggZ23FJLDlq
vYk0AMibMT44KbWWQTKZL4y6ydpxm+Rrp0NWHVqInnGVgiNZuDV88FGcU9sv5lGX4wqA64/5IG1R
AWYAYNPxaxsJ2M6hX5l9DbypQoGzFDn7xo5Bnr+LPA+NxfsifstvZDnwPvVHy5V22KQxenYrmWyR
IzAgmsAMiPJqwkaU9Ceiy97ZbyEF76uPU9nHCf3m6PkJ7sPpcO6zcnW8wd4Su3W+zISEl9MDvp2V
s2EViRbL/iCP8cnlc9OCsjXv02TIaWv6VVuAJHq91Y05xNbypJuzbUyW2qeVivS6Xs8WhfiJ194U
7q7smjZokLr52Ro/4nqvDOq168FRsLICwXvUnl/hIatj9AthzHDSCvS/oRCsMBJfloVmIYyRh8O/
iHUhrq/tOByJbI8Yuyqm7WexVrMutVY+Rtr9bZ6Y4vdTACSXE2KSEj1jfCetx/jWkT3GEzQIfWSV
dIdcr259sGE4OCh3SnnS7aXg67TsiYrVaFQRNVp9WU2JOLY0FF2bDJV53RZRBNa6WBLWrSyU1hll
5mWfiryOB5LHI6K6wFEZogQB8exFWi79XAcFifX2Wv1xhcJhoPS/KodxtvatwBBjE934V1bDTQh0
YLXM1bOX965Nf25bKHHuxURqaCtUltYd3RIHXNM9LLQ2pEsXiONLlUSbZHOBk0gYq2kRsAlTt59D
mB1LTAki7DYnUZg2BsQqHWy1JhR5Yl/XZ3aX+Cc+IY7T0UP8iRcj54KcpTX6tav0vxbAmWlqBdSL
RmbStzfTMOnyVjY+wOP4LGG13hqY4tcj9gt3Ou1jjnK7EQ7+0HlApATHB7meeIBDIuOVdO8Le5CK
SicaZrjSHvOULrd1KFwUtp24GH4Fbhq9mtw5Lj4NiWRG7uWYnXzR45c1CNY6Q+6/D/UMjopCzr53
L6rxSKoANJI0EtFsUtWozepwQsHF04GhigfCeR0+TnWFtA/4UnLLsTkJtOuw/a/O5hIlskb/VDQ8
RWaeJIHQHMv6kMcXZOJF0s2ACvHEJElFmr2UscZOpf7SH9wfojw4dxrNDxyn+zg/dqYfP1KAZENH
6xE+ioJHFJkTq011DbkKMDW/qkdje4jJhWbhzKD6xTxOGpGeP0dJdYCMIrA6L6erh/1So5wt6OTL
5FHG3VTaFDVP2yZ4CZVptBV87I7Nl/HtF1TGtg9UEdyi9X5FprpkpD8Gi3xkx8SgxZn7b1AM4ZRE
KgsadomOpdTzglKyhtcDvuiARFAUbIGnChpv4Gr8crL3Tm6U64LlpXOAKXcVrhzZkuxAXYqvu1Wr
vihqRFAf2RIFuxIjAUNykIiTw93kGX2dae7+UAmx4/EnnUIUTtkFm0zqZl7bcDq00Z4sVVsjExGJ
efdMD0o97kzAkp1Ag5c8AuE0e3uzPufWgSp8U+lrPAjUrcEfLPgZiifMvn1nINEDDzy4jhisJxqk
KDiXFsNvVRXbpKVsybw6577yRHo6ApImuAxxaGX0DtmUBqyQprU6/3TjojY6xYzM4IO78mAEbyZq
raFU+4CMcDZPk8MzWGUUCEx2GyXvotlttwjYg9MEJMwF6sykQflG/M5m4pYc/fz58kEqHnOv36mT
4at/cN19p7qi9X3FsNPVhss+aOk+T6SV2zSFKU222V0Mjqsoc4olFZwBdw482aIQjz88pjuSSU+M
rCLeDWONZJm9CPuykXLFIvRKMh7ze6f2I4pOFaZbPDPVQ1R9abx1zmBhNUMA6iTim+TBpEZ5qBgg
SDxxt65GNuEcm6yxsS3MMjOaMHnm675RU3tNRqfE+vT6RXqup5Pfo3KsnYvDinXnTxdnG5wHc2jS
6In4FBQuB+wf+XlcsZ+EppSgYU8V/kj8c3je2RKa1i2HtPysAUNeo3HTlLR17fmapEeiCUXI61GJ
bYL3w4NhavdgJ4HqCbCoAE3QG6UGBPQuUDu/k3BhEcprtgAZRORyO+7PoPcktUHkZwVrrsRsczWH
Z7rDVKZ/DUAYtl6uCZhc+Ec4YVRvjCgVTot6rVrQ2yiX4uegykdKx76YMOcPyAGa6ZiThIL6P+qT
DkeExVvFwzET/rbNYFQkiub2k6t4Lcst1HkHdD+XGtIwTeyf8CFGXxGZudbu3IRtLt8oL1vMJ+Ox
Vi3194goc7iV/WeALyZIE3ywhWbw1y7XFSsP2lCMRVnJj2Mxb+O0fzApE+1dckBYO/ekwju+4fVl
Xo7X89X7GzNLEF3apiIigKf/6DgJgXMbaCkw5bWdM0g/zPUpbRDvtdHNpzmJ9CGnlV3dAD4BJFaO
Bjou3iRVfNIMgU1esuMO7SNRFvTr/y3nmVM5OYheBb7SaP+fSZo8lyqQq1pDxYzviG0wZlfDaG/l
jfuEPZBieG06wmL1EinV91nxCNxJAu2l+f9S3xvr0cf4LBmWkciJvJIFX7POOiRTMyrnHH8oCq8p
5XuVN8qD8cuJxy7OgWv7lAo5qytilz2/uFfenbsYxHj6VFThBYV0u6Lrj+EjFR2hTIi5oepAMTo3
NBXgocPd6Yd3iLVGNW25HbNA26em4aqfzkGSR10+mvsbQxSJKhp03f3sZgjegrgU02MCmh3eT2Ba
cZa95asqNo/WJGpQwsZnF6J8zK6jcJYbdk0pyPkbGDT38cjGWn6qV26Pk7268Dho+fVr2wlK4ulK
Tgk2z5pp1HWL11OtswEkUjDtT6lcnMaSa3faXckrJejGtGDZd0+B4hNcqYpJMGMKhfPTqqFPuon6
kO+eY2h7y/SREwPyLV4tDkFaaorR5M+Ic+aIBC2AmgjfTbT1m2oQVYF1BcE4eiLZLVbZBeIC40ez
bitTMlvOa/jt/A/zYJrIYVKdDlueZ+I7h8FqnrVfjjC9TDPahgsn92wpNLfFQI7AJecEDga+iJK9
nlp1vF6D7sAYzzCr7E7XSlxAw5vThKy6+7extV8B/RY610TZR269VxlWdLMtoSlYWB7klj+Hth3h
No9+9RzIesQP6IZVz3XFNEWfigVdJ/s0NGSxpHZ+JATBhW3r+07satzNGe9RUXmt1yrAGXEN8n9d
RNdjvsFGOfmhT345THKmGb+Rx6mgbHmT6eeskFpnIRs0IE6QwjN/pWVQsDOCmAeEy6atTApaRjwt
ubXobeTQs2OvPH+GwuFYqAWGGj0vZB6z+PW23jYvU5MOb6ChZ28QUffzI5oZEeawBoKLGhUi4hVV
aGhAE4WSZOtXOz75YYVJitf7GHwTra90l0On/REPi7088WcOiVMswVWP1ZAFaIxQSQzU1xzhnOEU
79aaIVuuzpmgmtWDmQ4P+kFg/1fgu0WtY3tGAx2uHDrUMlqMwr/bENCCVAnCFF3KPB56p1JezxwE
f699bOec40gCvVqjtNpwlx+S0yNYYYuzcd1gB26KROXmsT2yDUz9HN2PY5NcnSNSZZmuQfhOraQY
8gsB3VYFjFAvsfHvZg8XEgrwxExsccYrwcXxnQWJ4P7HQLQpIeNbI+Wg0zDb6XdnUf7RzRZ5mNXq
1UKovgolhwuWr61JS7CfT6oTIVWV4o/9WgWcOK6yj1VZU8v5R6hHb0A5ksWymvhjYE+qJXX9tU6b
HJjZirJvYmKHl6zA3/4epFYpg2gg2NoJXbEQP/ADkoFXdq7sc54X2QQ49SFHjFHW73kN8/qd4Xp2
N7PM0RbQqozu0fJeXP/SGfOB6usifJ19fkCiBdJ7DmPybONfpnZBFvePUWdpQPMtv435rhEODsBs
AYAWQNSQpIXxEODi0KglUdOJCttoxh1IKz73QPAP5bPKvjNZpeXYvyllfZy3/lfrEPYRbJLbOazS
o7oKLDBuMQ/UvZAP0se1MdF8ZytS5HVNDOZamGCZC3Mp8stxcyJRTcGMmszf+xIXgZYZqb6Mmj3y
MPSdSss+iaeR1bRBUb/FoAXEtO+X2HsHP8flRVUNjMitEGsfkbhBQiLDThhWp0McRHu1NTZ3H2zW
73JWNJPruadeIrbAhicxbsNu6Kr9nTBTswbzW+yMrbQEsiLcRb+hRxswEbqQtL2g+ttSzb9jOZ4P
Kz5z5XS5GtuzZZSgCiAOWMqdhGNPc8Vi3ZLv1giDQt+KF0KNqCg9scujR7vxPjKhYxVa6e4akQCm
napYWD1gXHjBtmneEkV1RHRjPmAa2EYxRTHia1gWQTBksIE66QxT4tHW2/qRzMxAiSlh2D60sTge
VCDrO883Q4QnFPul70n0fir8XD+9m7Rgqsz76QrINy7k3orzonPTxz3M7ExpSfDREgvUR9yT9nIg
H5KW00grXLHA2QlQIHSEiObZDq7u6u+SAirr6lxiJEjVBdd4eIZJUX2MC3ZvTs26nu2h2vShokmF
7XFKHOZyqa0FWbYUlkFcZMzpZi+mQyqPccDP0pssmc2TAchxaPYzsZFs+l8gGkgewIQjEvVOmRjo
ogdgCE9EvLF4hoKPt1lURjzT1RrPE0eo8Uq6vJTVrv1A6znLTlM0XfGSUF2RhaXR+d3X5K5CIM3C
Fvzl2OzVCgTE6j5jOOV62bYheWt21eoMKvefp/w5pQx6NpY/cJI5Zc98nmy4cZx9kjN6lAk6uxf+
dJQ061UdQU1LBrPW4TY++Z3fWLU0erWp8rO9K3gwRwuSTDdvm5sAv4BHlqEVRnu2cHVo9PdSt2Pt
GZ8UZFLQW2+0vC+2btMxyWNMhi//zjWx80V2wZltYoMXn7FEzmdtWXpyF0t/fui1vXisSIRMOYzZ
84/wJ2ZqB6hpakUWvlLDnjxSCdxd1i3VcJwu/cC2xfFdwnkRPUcAJhWX7AxwzRKuXM13bHkRd4q8
nDK8IWxPOXASEr09xHT430qNDIV7C06ugRuvwrB7KuFzjZiU8nAtoi7W38yOeW1+mZcGY4ttrb8o
IsX2G6Xp7o4cKFnKObBOuu/wqbNPGU2g1f1HJgwJ1TJSjOc6xNKdQ6UI2pwq2W/+F5ZlnoK7lKdC
DbPzp0crhHADtJxxNJQKKueK4+imQlizFFpdRehFmIfObRRfTJ2yUobUu9pMv18lcljKxigJCsIu
UCZzDrDsGyZyimo4e1omso6zKxQbGcRVOIXlGLqJ2KlJfCfX7U6OZi2RPmhkQfNrOm/aW4i7EG43
9peNPUEsMHIrRm2KzLKrxwYnKniFo/hoGXwvVtpOJylA4Nz0Q02InSEf5GdMlvAOlQP0MGNX8U9J
qcVoncQLE/U8mImWwdyG9p85FDmmcJxdqv8mdJ8UsG4lYtkp5kOAKl2fPV1w4tEUKbwCl1SqsulT
7UDgQxmL3JqyIIzfbglvPFuFL+GZIKkqzaky65X1Ilgr4WD+X7dMozUS410LjfRS/RuDNuhRMzs6
xpocr2q52gsX1Ba7cJd8CdabQCYO/DzLz/Bzhk5VImOgLbnvoPYxxDTvi5ByobJW1tWJeYIsPoEm
A9/JifHWQ+2pqmmMnnkMDjA5+YgPT1eCffJjW+7DHSbPvv0GW4KNkTMHYLY5e9LAjvhNFS3F18T0
z047wSk68kUCl/lh8+kdfPXTU0jLQfjw5FDVgoxaFqu2wxJu/gwRXE7Et9n56K04w+tGYPxSD56u
AuBa7Be3B7Z+vCugQHibXvWhN9WqiaZLE+iGuzoCwa6yEj3+1FGujfxUtilRhGTT53uYRavaij00
Ai4k9dBpiH74MEd9dvNMbuSVvB+LFA48lLGNR6G6NDlFj1lwCcLnx/GIVSVLKPxtJ5YvNhHx/56m
aXGqL4/eW5fNVCCCusQVU2KzRNNw5teJecnXvbCFEpWvCqRgD/YwuWapZFNKsZV8PU/KlDWZo3VN
xATDQjkPrb6BBtx7/tYVPmnVz/euM82e1M6AFZLYgo8Po0GWq7X2LyGVgB1bpVzpkF1WKnlwe2DH
Bp7K2831nb7lE1s73LqZC095XGGw2CQdAH2RsdMz0T2LISMdEzExjmS75wluhjGUDM2LHixs7vXk
RjYb4sgKBWxhz7huu98SbyqhB4LRTyUw/vfYeTtjDngMCDK/ucWWsjtkWek54ywVgnrpBfIMqv3k
OHDGGewgl1pCk5OMJskqKdXrSAXuGIO1KO0S0Tchla17MxBkZcmaczlc4DQI9WoN8X/6866xUTaZ
zfPAvYz40m/TPXaxyr+nMy4DgWYmsa/GaCrWQfc03HfDbg+ujVu9lh+KE1m99Ymn8pJxpdOoNb3R
QQ1FuCK9XqRYLEeshoneCbJ4i9T7DsBEgTwWpd7mNArZy3z7pKPVqsXJ7ShuRddu2NlhewHPQ3dd
lpXKFmsrVhRLIcIOnz57IiwB1+nwhCSkWuBk5vKQYOjkhRO4O49Sx4lVZ4TsfA+YivS5knyI+dad
CGB31ViXVtKYAxANTYyJEi/kdYv5CWVlVAWAvS+/RQcL+DIQ955uR8/dFIKVViCQsijzqBK/jyGT
t6qt27PcC442/iLYpXMtvnNTtupNId44wIMhqtbSwQwMq9xfbX7FwRXfsj4V012EA5lrJMFG1C0o
89TOnCsPWcFDgmEPwlZQkPVTZRW8BFuQ5zHS6UePzaGXnonD8KMViem5iQFLZUsf3gQvIRL5TW0A
ugh+vpmimpMPLtfcO1X67PSKaoOdrDmY1TSclfDxLh45h7k3hH9T1VsW6Vr/5NXkSAWfdPgViyYg
YiEm87D5uyTUOutMARj73dAifz2PIwFFwW/6VOYv5JE6NehBHz2ziSx8TSIs7bEo89wynVUjTwz0
Ye0iB0EqO9WyhVI8ZvghJS9UcFSXoieiSizumyUcheJ4hQibPhX85qqAbJtN6PR/ckQnofHN1tmf
0Dr4UtEG0n1Mu/7qfmPSmbL9aH3PfLOAkD2d+fgydYMFfQNlsOWH5kzVnpA0E7Nqog4xDc59tZY/
L4hj5e+GnGPEfGVGIXZmxUi37AHSFwP01dScEGS7GF/pNi8QwJUqKLlSPaWsly0PT5qftRYoeZyA
k9zgMCokazZlJcAQmHLOvgQp1cWgQivd4CKJrB43/c7mhlIw1OOsPAzFBvuRBDnOioRoshkb8LtN
79E/8k3UfJlS8Xsw8+CnJGYR/WccA8g/6UWgLpUZwMzdvarlZvIfdZHuqomqJo9yvjq2iJs8FJ2m
/oGq8DpG0neJhKaDgxXRGMnyI+SZ+SUTYxjwz+9L6wwgSnBG1lEBH2zH5TMrPrLQyF91WyyW4Bm/
0yKnyfFW+YGHCd4dK/ub+7PAoPxWAStVUqGi8eZFf/hw7QtLp9CxIANeiaLugGdxGwu87TUGFTtR
S9q2xXY8flNPw+zq+qUVD92EHuMTLvH1ksYuHjlhT72699OEUkDCmwxHvsLMitEmB5zYSmRB9w+S
RdH7oD3k1pGwBjjeDiodrd7SD18/kwknveaL7KFWQoAq0r81BdDyh9catT+YhnfCQ+2qaZ5TThc6
9bMt0VWGYE3eGDu8DX19e5oOn1uT5K6blWsnE/EWJWcdaJK+t2Rzq6i5qRIZ3wRpjQ7lQh84WlB0
V3Qa4c4I4Vq+lhWW+OSW7m60SXYWPU7XAbTGRrfWXWQax5mV/aKHOH4Wtn8WCuzbHiEOTJdX795N
gYfVuiZgkCL696KnHAPvXA+Pn29vb9MnofhLc8xohXBnXNnfpck8dPz8eGgDaTvlsxWsWM+CE5I7
dtazKLl0PMw/tWTx/BFfy+DpxLZR8JJLmLrVGAfHVRfrHoPv8QCOpuV83RfpiJ0XHKR8Du1IHJ4x
nmM5RFlta3ELPhrRaevEWfGWAzvG9OL3QbQC5PS+377ea1e2D0/qu50DeJcZ7AeRQpI7j6Y7g7Rp
5GjIIjuulzgeZpc3XMdpjuG3prag1lLNQuC44LpD0REbMnKhLAHZEmKFIj1EkziVOVNz88ys3FoG
XMgZ610bgJ4XQ2130q9MHnM7ZOtyHWzbOj8+27t28fNwglKNvO+gYQk7tN0c2eE5+AD4YnSV0n0i
1SL9ECq7MIx8QNwKT1rVIU90waNLX1iLscwS5b5/1SWU8PFT6rD279yZV5uJdX/Y6uP5NrQI8QA7
IQ5SII4AWVlWmzWk00oqc2hp+ddaR3V5j0s/zuCgXIxSR2B3qcZW41oMgjEdCIPsQo+rK+8KH9Gj
XM7krFiMJAl/+KhYCyGG2uwdsC6vvE3DqD+3V7K0wx3a8orGZWdHmlJG73tLK5qdRYmja1CdkrzD
vT2VMXjmNlWnfGLktenAIlyiAwtHQ37AINScZ6GRpY7iDXZxw/Ro1Y66iMBWthUR64JhqDejgUgJ
SB8E9oKw6+Y7/Xf/z/rkTwEIBOR8bwHs0skkftGXuatAQneZI/LCHXCM0VUbqP+v0uBtndPWN8VD
Tq+SfS6sHcAIM3Kc+KP9Vn2jAH2ZgDx/+Zn8cV71BwvkHLbNF+U2HlAE9sw+bZ1VhsGZbAyBnH9/
fZPZyuzs/5Wq3CyxAfUXfikNMjWOe2za/Jk7FP86Sh7AFjQ3JY68SFIaH9z8qwtHegFE9yvVfPBP
PLtwKzq0RB5Od8q0ozYZnxmImMeaZlwl3G559zThAUo/2uA8i6absCx4ISSiRh5lJTqmMB29iUD6
9UDbZGljF1c+PKaBZYzeaHB+UfN0J297FDjEWTIGs05QMNCQA2xv+4/wcd51TVq2xc3sfbR7/T8D
UCIbbiv/QlA4O8O0wk72UQpbaJKgQm+6KTZjgf9C7ZDmaphOR4OLlZWicVC86Y9f/Jy54U/wFqPy
OrEkXBlcTIktHtMVdkGpWPbcgpAcITb7rKokGVocsLLZTmkxxPXwPSzfttCVVshmfkjD5kq5xxnj
cQK7jYWAIkeFhdRyhaEH0jxZP803+G46enNaSZvRkwjKgAbukQBafQ//lAwWAVaQOQX08AobXYy1
Bl8TJYBukHzBysqMx6wH2jr84myHyZywuxfMtTJRH26zq6XqZX3VZhirof1cT/RF/A5jkG5CLyVk
mCO6pLSqMLe2Y5fZo0r7dMUA5VhZ49dpj9KPlT65yqNbFrGtKG4RAg+a6hadvNSeLAdAZz0H0gRd
ojAYWXaPno2hvIXwCZzu6zd8lkxoz2keGQ98KHnofSbP8gs6SlcdLKD7wB5ygZeJUIQwG4ao+3Si
1YPIbwp+S+XIVUg6wRMHHoBqKYBSo5QMErskj4eGrpayNPAi4MrcwoPbbQNXwLDQ/OGMZtISSYFm
gjvRryt+e5tcTLMeOQ5i3uXO9qGLDpD/8ZBx85NQicuKdjJkjk2le1z4xhZ4VODnwCGvAxMPbnKm
855/CUKnHlR3ALgU4rWyVpEeaQMULVEk2rUyiPfxN2pbOQFx/K4U1N+njUUMObTHnl1mkPxyqEb1
JFaudAyXqSWZ5vJJfbmIOXJ6eqaFcYJjW//b3G2dbaMOFkpo/4NFrlGWsVTWrT6FCkFtP/g9tlhD
NtpHMwi4Lz6oQWucl9UZvSMYdIxMXEy+Z2ejkFt8XY/UzYaD7LIsOtbnsleQbvgClFWrDdlo/b5S
Y8mQCxTt7SnNHiMa6jMdsF7F0+kQL9YztdR1igpIohiIUovragjUWNtFaaiDiMLmXkocWLbLXyOI
Cc9JLRTDuWeobgg+/S0jU8VHL7xKYfoCAA1TzZ6HkK2T0EwwDOehGEI6FDQ7wlpUW4xaUSBPYUTR
J9ziYT1hnS6iySA52rXEnOlVtrjseeZumkGWAtjeOBJg+LizD0ewLQ4D2uCMUE7y/8UrgZ92OjJE
x8PTCVJxrmKfoJ5cib7NOqhZ3JsWtFSts01BWHXj2wTWU9w9X6AH02F4T5YA29xvjYVo7RzQbe5q
b6KU/nYynrGLMhRe1kJFbA18noEOqRNd7bmCoNVGIXn44mwblVnshuW3hETUTLi7zgtSpVBLu2QR
FxAkGIgRrjGx5VAUqsyTKA4JvgW/UWCyA5k9ypU1CfUK11H4j+FWa+xMKUW+VWNEn0xN74SW58Ox
mH9qfV8yZ4xWwSqruWiPaPD3MaU23huQ9ZtZ9aqGsOm75OJ9q73x3TcM4bx2I2xFTCVrUOUAZjyp
hDALAL81sombo+hBYGYa75Hg+aCQ1XrYH9i3qMk6h0QmyO7z6K866m0uQafDIRsXFn+SpDhkjVRu
m+f8kFqui9PzqWAXNjXRJORkzfDOtiLRO1IQ3jGTS6II7AitdMD+M7hoU1NEAv/0xYuHQsNqu+b4
JGX0DBtVBzaHx3UDWCaJs1OwNvJyTRPt9zOz4M0CDPdp7o3QQXvvV2pEe9qwy1NZCdsy6EY7Zb1C
nllL5A7YT5yHuNiatQ9Y6Uwa7JNQycN7WtyjRUcRii9gGM5NOOBTFnYopz7n3NAIJVVactpMUmt4
Dcx6aHOJOrs80uhSzktpfyjuI2UbCyvL2xQLEvwzGJi+npVmVc4vbu2urZ/Y3qmoLsGj7kDLN8T3
/E9NnSro2uJdvyIBJa8eqA0fASd7Hu3nN/+5ZkOTXApXtZygSVlTvMjJDsQ9G55dc41g/dhkDY9+
e+N01pp9YbhJRA+k2Z5bHqm/L/4Xsw+/AfyQWvifJrFQfH6xipRwx0/c76LEQh7Trz1uuIRxxDfh
GG+yFa4=
`protect end_protected
