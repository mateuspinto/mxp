`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
CCcpSY8TAnE+QQhnjDRP9i8l3hQvFOkE2mBRcW8yPLSZlche/7K5uhYF7KIHCyr4/k5umLXdyx+F
pQImQtPUfqSKOBfBB0qpnr35o5VoPfTN/aKcxo8MG4FI5DFCo9uLGWCctHvrt+CDnzY8lUVWMDdk
DMRokFO4CnzGx/ZHhJCNrJeWCdWB8CaNv/xJP7gHKg1LPercTuK9dgU2vHK6jV5WtL6Uo28Xm+n5
xTbwt/Wzz7tqz/6cZ4EFZktctoCzhyL+kHOt8zXShNlYW7r2UNmTPTo8OGtaa64bmHBA8kYfUyNF
NL0hw2sO6MIAtCblG+3GP/7WuToZbXAm9CejEw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="4K5PRGgwIpkkO5qoQhjvuO0/NvGeVDBdue85ilNIuR4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11712)
`protect data_block
w/cKq4WiLYcmEMM2cxBlaA/W+TVkO5gB9KStHjzbgY+ApWawqPDQYI1GlRdK8EZQDwDH1X+SjwtD
X3DJKCxSwyLg3A2Tp71Ho+DTuHPgNQ+BcyJ67BvxjF+aRVtv+aczMw6wZKtuV3kFiySYuSBMVj5m
v4pR3VDYMKh5EFTmTIcXCcWAbMDX8UsyKqhw/59+CxMA443RsLMxV/4OFO6XBudDgI2fzpzquiWz
PKWQy/QaHMROcBlqO4krCIy3LNnnL4mDYM34jVjvvVB+PxZqmGGL+FLG7LlKahgPAQaLtnuvOUOS
Yr9RrmziqaT1/dKjI0XpdRxOvg35/JVwp5Y6BHPZ3vlRZ93/V5nI45Iq3ziGZJfCAPkc4RzuBoeO
xDsypGiP3AUQJnhVzezJUydDdHGXgLlZdT/S23LFfCUGCy5/uJ4D4JaI7SoHMlbMxxd4WhKoWHmN
n3rXp+I/G1LTdeHZ/IpIYawt+1yeHSfpenfvgcQcC9hZuPrAfU0hb8GLfSo+1Yd7rffihZDAokEI
VZqyyOAlgUMZhxZwPoOMdFi/t3w4VkuXA7sgYgPPlh3QvIBBiCewFnZeUUwTe4eoLGXymOx5Hk79
a28ve4T6gmAjhjLCdDirfhUgg9j7x+yJ20dtp9Jk8Ds+XReT0hdaehcM1Eiahj1ZjNDcT0gHu9Yd
T3GKUyq+xGqiH4rE8jTFrBv7ljP2ONofZuFm3z08aZRFzCETR4j+M7b/bJFaZ9wlGKTFtL1h8BLF
KzDab7of5c+J6yb99cuzsEkgSYzoKZ63mWnmiFUYX7WMR2Ag9LFq/WFSjKQqRWNQGvAqjw3pS+Hf
bF4o/QtlLZ5TKQ9+X1/aiwySzgcfng1Mnfk4REu5OdVWpr90lYTxh+zUma+yX1AAY+qA+USw/Uv2
bSBgJB9+LEcnmOsd+wxp2Icz4MI/Vqe8dX6GtS2zFyF5HGRqI+V1LWn6fxProxlvJOydgjaEbq1E
TnzXYv2anRbwCKTx3HF9+bta5q3CRzHs0XQieyEKOtArHf8Zw9xgYxiiLS5QWaujKliw+jQ4ieoz
mHxDEA+bZt2QI24H8DxGv+nvcPsD0YxigVJ2m74pD7KxJZgaiijJ/HkdtwQMnNpqZqYZ92YtC0w1
/clc/I5af5kknnNMxC/u8K6xlanzDybj2r9Lt9FOJ2DYl8jZ5ZheIG34yviYKJ/Ja4bc8efJ7vsP
cQsCwpRkeXBlRQA1xQrwMi2oTOYq6vKNhJZRvxJ5LU+7MAAXicg6i2u6c18k4E1Kdi4qvxAVTbZe
a9r4lc4rvsT/tiBvKeK3r2j7JC4MTEUEi3YCIq7UoLD3HZtUYT/A9Vwj28Rq1SF5lwwMe4mnELMb
6knd/0j1ibJKd/qYqtsnheu5kdUj90fnunPNzXJR+KfFQDH85bMunUyQACnX4jKuXbfhSDxRCagh
Q8F9+xXrGdKKPq5UzBrMymJpmyltN6O8i6iYkWXNeY7whZ5WevW3aZMJcVOTxWDQtf+b2wnZL3F0
rD2EAUrf+TMGd24qvaaJTX41jRBuHORYqYAgGTmjgz6kuQOyJteQ8Oy4cLJrFPNZ2cr8yR7OLmyh
4kR6PgCwa4jOJu819Z3I2vBYHUKBg1ks1BNKJU1uNrnJxCUc0Cf8X0wGow5jeA0qcjXRZ5hRmrGW
l600nQa0rcl5zZ+FsfSMvXAeLtHRlcpPviBGOjl4ze8d14Sn6x+cqbQOLuDqJJ01dQVJJuv5fDKT
BM31Sa1kNjdpRqfIXplV0+F1QUNKSuat9+775kzRMs8tEFXTomAsv2GOHYVgmclbuqlaxq3ccVXg
EKSGi4kAkY+aoGdu+xj35XNz9J60ktyzmgsmM/63Z6fzMmYDhzp1llAs/hTqNpa2XAUK/kbQB01m
fBiPEdBjGdUOzdGiZ2E6k5AhBp7pLjRwgbR/mR3BBVjf8eGB/7CnKObZDjryvGMC9O88vwaJNJCS
GRHAyac8nmPpgAXQ5t6TglXnON+t0xGs3C+c2e4iC7cNJoedkdAClTPzyJfTcPV/FMgSdioAfZz3
lESqKO1zzJ2vL7B/LMmpomqc3AF/kDK3L/V1rA75uSZ7LUuYex+8M8aAQOb5/HRcXrAW67nlGN2C
tFy7Xlu0WNs3Cz+jjCqOKHDgV3ffs5hpg01HLyMBmvHidNcXz9xo1ZXzFYPTchyMw9pJRJZUGHGS
kV/uAYMm4wXQxL9X68Nwypx5QO4Vzf5FGLciVhcBC3piCmJXxInaSY024uV2dwmvPPWI/gBCEX2x
A21cTd98MJkr7KfNoOq2z0JH4prpRq+PHJBPU4gk/5UYw4FE3HCMs8GbtLDfyZwQ9fz+dbbH2sK1
t/5T8vnPlz8wlhrPkfgvOFS9d3Vw0k8wk+RC+nXPjzrXIESkvhyRkNqyXZsf+ZxIpavy5nkvD4cl
PGasTyMexjoJEbF+prenQtQTt+owGuND/AgHaC+KI7bQxDmSfEwEsLrTygP/YqnpU6IsllxZ+LVk
yGA/q0lL0N2URLlZvnjjIMx5quQmGkJNgmIYTfA/QaksHdGYDSOpGfBZnWXK5GH9zGZniUnaTBRt
/a9oqAdupjH708O9V+HpTK3QzPQAlc6azv2s9OgEX5ae1d7C9WtcKJey5brx7kDFezG4uThgvZBs
g0TFPloNqQM0GpGLgw/JFkNqwCV/X8mGN6a39lqxe+++Z6Wnx8BKtyk95AimD3lq6B3mR4ghbqpI
KOnknGAKzQsYbhkKZy4heTSJ7e5HR5Y43us6qdR2E/4A3qMyV1Vo0ieBaZOPgYPmyY9QTNQw5XHm
pBt5F4hCfK6KcmCoZSCieAlyw7wraMeIK7wDfD+rEzSzsQh4ox2lqX2A/kUUe+fGunaDjTxqba9L
EjHd0a9QPBs9JmBuuHAOF4zfR0yeexYIfhN1TJf6zwpz+yp+j+FmjE3fvK+VZIk/OErey8qytySv
X21A1qvjfoAyvAj0m3w4lDC6VO7W+M1MJokNSWmwvpgi1uchY/AB81RZLv2wLCLsJ+WOevjHnaCL
J0NJfRjPr9TS07GsLSvJUgfC4CBggWxTcjl4gvOxUshIJDHHGI0xGwDgP3fMOML/6GWa1N9LPrys
aFQogZQT9/9rGN4iPxTqFSwFgh0EDViQP64oCb+3pW1BpcvwkE0mtiFusczpV8zz/Eb6Gaxh6cqI
vFNqfRzHXL00/5OjE7Y/NqbRX4s9fIrNlOeti080khJa+3pJX/9MNtJcSfPiqAItW6eNaeJKjHE7
av2BhIKHEIlPiadouVnQmATEvYUwN4F6UBoLKnpvzA0uFJW5Ty6nfdMgGAonwcT8Kyc1BORqP+Mw
94cQ+HPmTagPZZsMKa4gkL9LIzl9jtn2x9Rd5Txn2LujBQe+Kzzeg7szi+RAI/5cgVrasp15jkVV
GFVz4H0EdECL7T3MfH3/263hVv6/2CWGF0d2pnxoZWU7SK6OwmtbcPdxW78mjVZNXTYTRV5lzvUz
78wNHnGUO/Z6sVHG3VYWbNsv6+REDHIa1Ty8KjSsmI7zqv+oqOM9RqpUbTBuOB4r0dEOiPIs08BY
Wwk6mUPBWt//9OrUT3ocNqPeRjIoNlbv+AgjpXbw30Ahd4a/nDI8K4ZD0lfCtlNrYuygc4N5UdlB
4pqqKPEKwTCd6KK6bwk2ZSlhkLR6mTw1bQdUtWgBUVib3kXtWr9KTHt/Bz9ic4ztg0gVLYq8nRMD
NmUUEKloca2f3+KzDVdD7pFxNVRaETDR+rN9cMfDvYFxaRqp3F6um4g69mpZkPHBe+vFv8CDmQTP
9LNqhCwmlqaW2KznrU03fHwFqAQnz7dzyDYA9zQsUFk1EWWSumW41/CbHOw9FX2f63BqAJLoxTmo
a70khusMkNFmc6VldeDK1kaN50pG6GbQqsNmiQOEsj8wo0T4RtEq+wcIIjryU6qxhEXWrkSVpcUO
LxArpitNKPGz6o7+BEOG4rQsnhilwsaR05UIRtIcTyelE0vZV1hwgQwgrL+xdNKToo/VghXp9EFT
w/kvj1MqqR1+iJhsxoA16X2DpLTdd4k7vvvsFH9k/lS6pkx8irbO+kwKivsRQq1b2Pqk/ZE+zPlw
5HEE7578XBx0j725Z8qOboU/9hajJzkU8w6J2V8EFuzD0c0URq+ekTpALlCEPRXAP1UTivVbPQcT
gKhDihcDn53yjdbWdA/XMyfc3uczmRYLHKjTMrW464far/G3brsm4WXwlVVz+KhWJ6vxC9GsMZdY
l2VzSMsBZl9N6Fet82fc8uZq7KXrVXlBqJ4HQKL4XGIIVe2+H5sa+KuEyCt0iB5yiyR07qiBLKjc
Kan9whqMHjwID+N2CM5M4DA1o5SbYA5QHxvPcx023fhL8mjDA0xz77i1xCNfAsFPEkZg2CJsvO3U
CAWZwrD6cPCI6hSIRHN7La2B0ZlSyRTDaKc7Zz9liP2l+KB7d37bXxJL91lMvyvdtssAoUFM8buY
JTJZHJxiQJKjVZV6TZSkOX24oKFcC8coBRNL9pn/A+cgWWlZ7kEBYqtkbxvIcTUVN2g1SA53Kpc4
1ZhVR0pQeDHNGkYThpEFcr9clVABJIeBh21p4sEH3MT/Kx5wv46nE3trmv5o8al8O+hf95oFFjWK
pqE61uMG8Ny6xXpwGvv+i69nRlQLYbDGx7ojZivH1YQTpivXWSl5PQQlqyuMEhpBGDhiCxd/xfmX
oJquCl3R/wQiIEXPdjvW7c4zlCdxw+yGqqQj9AMKEd8NggTomec1j2WebG0XDUC4RcnmaV9kMbMn
twgGxZqX8PKcuotwxqmonmNL5swhKaUo+te+3lFeKKNeRVw5Aa/bhhh63TdgB8rrsI/sValkPTZb
J275XuHeuccaDm6Q0Lox2KzN3424uiKwh/xjad4l8tPFA5GgxwXHdH7zwfy3vulzd/9Nq4qFP2r8
Y7H2u7GO14Dt8tavZHOIs2V6TNlHoVUcG6bhlN6Zn05njTrwMS490iWLZ+kqMh4t3pq0sMnrriJy
OBskz9+EWvzTCNCIK5yMZH9BI6kyDO3PCcMlrfp+QHD1suHstEKcPitP+XFLcY3ve7rzxHdHK+x9
AgdCtBavIX92yB0A3yP5CI/m9Vi2dywBHrPfBt7eWKmBxWLN7sFATioSvjYDdd3ABwF0QGIM+/Ph
6K9j2QZYitIqdT67L/T6nWu2e4SRzfvUKFHE+YmxfpVRDNy8xRZx1sfpx9hT3GDhVAVO/oEnfpbW
BU+dNR8Bi+Uw3tx3kdYVts9tRjJWR721ujP5eNLGzHfR7iLQCfk3mt49a/zdMYckLFzEUhDn9A58
oLIbFhVOdg01W70IXlf1b/+FcVm0y9qEzFCLBxAjL1YSQetSslKBZspk9WvKc6sOAIRtnHTFi3SG
BwShkvuoXYFydERmxIEaJclY89RAxoI9B6eRX3A4IiOT77iJIPkRn/ctwDwkDFX3CL7pq/Lg7bYn
c6q1bZp4B5fBwzyo+vAE3a8pX5woTLIPTKud86LzDEGXLvHpj+dLKIAwQ6teFNyVPTIquE3zbauD
Atb6m0UbKuA8kecwSGtslYEVnIpnGwxBlVM06eZ0fiTWz6Ahfq1LOk+WYA/3pn+YR0+utpqc7zCe
DAIrzxfrNLSs+spc3tuAyNZdDBpeouS0z2iOiOIMJNPJMGg2Kz9iZOCMCnx5WJ8PqE/+SdtokEKG
FqzBZSOzUh53b8ioe7HuHiHzGKYmQg3HuPc7YhTEh6a97AadHfFVzmnqgZZJVz4jiFnUEBoBgWNc
J6p0eIzOcYpy2BEzOgd5DYAVyxUvaMG/14ZtZMSRBRTpAk5VSj/hjptVwlBSXNA99ej83IGk4XsU
sN6r9tOIdQLWN8CLa/veR0NiV1CcqgaGZsAojJKgiYcW1ZioTl+2MLP6imFTDgwCe53i5/S1TK0S
xnW7kLwMjhxgKIrkDOCSKeyZngqpqskP1Pyt/QPVncCT4EP+ebyOJk5JvjbscgciCXlxc7ANY7GK
/FLZWbJWPw00dEkEY5M6ETcSCrHfbHkrN2NGvyvcdZHMpHT+DzCUb2hqyq7JL5bvXxs2Yukcy6YP
QwHBUmqM88mZMg7KAaVf5ARLkxzlyV9V8zBcPU9Uj9XLSkL+ZTJB9fbwFA4B/oIIGfvl3Q093ow1
REV2rcHCyUl9MqK1HUMZA1xBGNHJYCry2zte1+sidioaddceuDbyE1lTHZ8xr2H4xPhpnCZJL9vu
ilW2nFG2smMCgCscQp80wK9BreszcYcMjAjLm2GRpBB2/i+SnrX6jfmOGQroAxpU0H1mO1UbNXVX
E9OWm6WFVevK1F3YQjSOyoH7Z2koTNFqLChWmkDHu0Ql4JHYVb52FFJXIT4tADLcYGSYrwd8c/bu
QC8EWzMTFdDU99LMcze8iM7sCdpeaVUZMuR87rx9OC64DElojQXvDNFjv/roT9JNyG2PEh4FFqZk
+j753uZHKNfyFh6NbBmJMc1IYfZz/4+x0sni5XjTPSw2eM/h5+QfdQtDREca9CU2cBGBQRrAyZsv
dbTm4nIMV0dkhQuDwsWkWxh0E15BE0v22WYuOSxNI40h9ihrNVR589tWiuQoTNTnJi7rhQ7IC369
X8L+NUUAl2DWbSCPr7lyOozQJqpNuXWTvwD6ZzoSBws8Jsm+HcpcrWwJKLvxS9aCOFyD1akjQEUj
ERyZOI16cGHxumMwY7ygnoPYSprIuRwnOXaBfEC6vjxA/DTTTsH6UxUl52GVN2e+bJ3YgeVeTuWq
Pq+MvnfrCN0/JLWpWPTUX8WNyVhRYSh09OSYvaKt8BtdMwQngg49cZ0pELqsUstkgJRGohfGnUNx
uMvxpbxE1PHB5a/0h0TgzhRYPOLV5iNr8wVVxb7ushxp5UE6M/PCzMTo211R467pWDKqOOan4xb7
zVpwvntAVlKNIP+vPDiImmC8TPjB8HmPz/+s94qvjjzjCAYsKR1OhDM15APJHUCLd4mlMrxYjc1e
/HJrZTIdk1Mgu4peZLvqOGJMXgBXU4j5lPSt9M8oztc/62sN960hCc38OB1TvSsZEjGDIzGK5+lx
b6LRmhSoAVa1inNBmDjC8dQXvsS3DZRBKjx8ay+FIjD7PvRqYbxlDVEnvyfnJ2k9BYVwRdRyXTOn
A2mjuk+w1XCoHxDV6PjTqX+ZBgo4AdXYrtFoOnQn67Dfp+cXzM0CsnxCBbttlelGpUIrFrOVMtxg
KI3gRqZjOMulalHdCaxSh7hlqaJGBpNoE1XSerqAoxjqxl48kXwHpnbVaqv22LcXJcOu6J/zjd0k
9TNUw/nMUTc/fdtHLbDLQx0xjT2Rr6DUze/qwYTOyB+PXqxDGlQjrs8tm8CDdIgf6n57RjHrRJNK
rUYaw7YbTBcsNzlqzCboIensjRrPSlZxsAqIUqnicEHIvR046G27PPlsf8IHB90v2nl4IBoo2KVL
mRoXz8bdeOxhu4dvs2s9aOJ89RMpZqlrPaRbYjhmIY3Zf8ywcxLrrA9r3DRkVhQLeQ/dTbkNAMuA
LpCdLYVxbF1oDsVqEWve+aev6fIFXdD0q3C3UswsclEzB4uYXwXbbgpNJJQBoUsqGu3bjMGqD3xd
k50p3t/Txtov5LL+ih00GJtn4r7jeLrGvRq87FJm5WRhpEOxk/CyJIYRd23XSGN/QRWAfOXAmlY3
0wlXr6qNUib5i8ClUZxvH1uTMX60JyaH5ioEWXEhFIgF62/cRc21WXuANH9WKa+tYGFe9DBDS2x9
StXAR37EESw1LT0ask1OJCDuxzBNc6NMmUhH5G3fERCtQx88q70xw8PCoC0XppsptzupCMLYsDAv
4lQzOwAFd70lZAa41cjipb7to2fHNHDiQl4aT1z2G2RCHBtfeNPBFSETeAPdPcv9wLNWg7tYwJ2s
IpNCb9Ia3wCVaSC4Hfq3wXPtfBaveFZylPbz/9cKoh9Gc8E43vc7gzEquFOGKLoeZZbCtT/HlX1P
Pa0PVPKr0Rt3zmy/xWvLavArwlVEV5R++sxatfvKJADdR7/sokOsPHu7dDKh2O3kGLAcXaUUK6ea
XIAfOQ6bd6N2xakUOOaBQjAESSgnerZKnvNQPgJSxPxQ/Au4S4JGk1m5w6ttVSpvHGVKwfE8tkSq
UIGzB6yTF7F4xtq7EX4pEdw6udbbQu2uyw5ZSVnpZ+8S7obgt8jUMimry2TBx5d9rkxpvRh9+Ji0
ZwbLN/w0vIGyvzIR77MTDAT2mFyP7MWmyvj/vQMiByn2YEd0ZiknXHJ2zFfwpgyt0AuCiuDjxoR7
YqsWaWrQqdaQNzpJbpykGRGIKZGAvM8arGF5/ZQG+rlO/R6Y5RYbN877sQAGdpuZZw0r1b/T+Wnf
u2ZWIp78RuRDPyZzOZX3cHKRHKMvBcHGn25X7H8BwpbuNxyLO7V8AcYH6zwUNzL3FBwVBZ1XZF33
wfeFd6hiBwSc9S2qXu4ncZC9kiBJlFQLu4Rlo7r8DGJ72xq1UmUgzqdi1WuM8PjJGK6ssntZMfM4
Fc4Oilpc4Sf53Y0QrDW1BVrRRCr5phoxKPxAGI9Yt6YdYIl2Y53MM0T6qPE5ApN/Z8r4sDEuEeqG
9USgTJZLZGSpCKYaQL0T8e3itQJEjiw2hcGZ51tCGJhw3yP9FK3imJg69rYa1Eycwo1Ps047UXTn
B/bHp71kRjieg7OLC4aFR6h5L4mwSk0y7VWO6sCnCjaH4iLpyzGNIAU1B4jK03TU4+c3YVrp3IzN
FURr5tzl59TFueTbPSLgBNPDafTuCX+iuTvbkfHZDhsCf3Cj0m95A6MhSKOQHAAZgzx726h3DYDP
0oMw3BUFHgT6dILp0QZW8fKnci3+jqpIOs05GCLeW0yYYf85iiIbkCj+4z1w1O2khHTVA6n3kvne
P0ofmueD8xX2yqi7awW6k+BYEpFABEiS6YmlXSm1QxSo9kbgh07HGYpkn9GQh7x8bcTSSaqOOxb0
DOgl8LRHadIIX7UsIJXRi7nrQkqYypHNPmpF/iVADgxEMBF1x7m1YSYw2I7FNvcGcHovi/kTNuXs
Sd83ncpIsyEFtBdI5crOtkwa9vAUXc2GIfG2swB9N4Nzj1MTZ2swYj42LQN1xJ1sOm2heFMQXnuI
MtVw/s3Lr79D8X3j8gacXr+KBHPRU520eQ9Pbkk8vojEFZtneK3BfSvXtUoFMcYJ4nQnA3YhfUwU
xX5mXQWQ3APYoSJmXkzcrwLhvSzhFz0S7y2mPPDVmaB5MJ/YzSnVwyVsbuJr3qECC0uH5CmFlZ7Z
bhvApGIgNhCRg9d1mLXJGWKzoXEtgW3KnhgitOWPhJmMvn44if/h66zOvVNphRFEa9tlbm5GRBLQ
P6St7kuZMWG+9bEsHGjSITe/JD/2B6ygIbobqrgqJtrqF2uObsvBkhOBdA540TvQc8/EBUMXbziP
ydjIaXttUH7bLXtNGX+WA/rRUJz1H4gMv/bljv4xs2Zh1lmfSLCUpnD9NA58+TcOg0t1YCMGBTpA
WsW1W1/bH9dDI13/k2yF9WkQdXXy3Yvwy/zBG6LF/utyPUwU4QTw4GMZY95ROF/xBdYvSazLsgeC
eeXcIA4r4Rb5QCChemjX9yHs1vAavX/qN+LVQaJUOxEfCjdAaKt6pEg/j/3zdqyI2QR+YB/MAxkw
ZGjxjNL6GmKN7WY9P70V+wx+Gg96IUvi19KsLbJyEH0T05L22MgQjNsM6HDLEdh7LSTFOojXLIqz
yQOp2GHLoaJwBpW82c2VZbYjs+A8u0fosNcEUBcwJ/P9LPZWk4RnD2AsPsUonnu59/WukIJ0B2YX
NgJcPo0H1biS9oB50kHVXEPSYIAbH3SATwuwUica4ep1NFMUcVMWQQ0Fmp97w4LAR3cRZgFCQUnX
BkBk3C/iWJFjjwrEKTd3a+dCdq4/jlnGVVb8j0UbFs05uvx/eHlRo5+XjNkbVqpTsnvI6C50ZLkf
8Yt9ZqJNj7EcdZdPYqAkA2lJvVGTQGgpp+4Fy+PPolEqaJQdL/QOlJK3lXeCy96v4e7/W/TjEm0e
/dCiMdJWSh5zIUSgZtS8biXTg12jNUfCl+8kf1OvFof4LSLITaOIny/lBakbzJ9F3jqpsLFFf07U
6sUgh7TdDPbgrklxLLUSv/5F2D56R7Rpzj8x3UMV4Lv5YvEJ8we0vz5IPA1G/Qx6S+6Z40ZBPc98
h4KoDCVmM9oiiuC+spbeO6Dm28hBABwf7UOXYn6HHOD/DHHZDPX7iybQJN1iVwbgGgSeyjqlf08l
Zjy+x1JuSFHdUKFOi/VjjKJy6LwT2MrVpPALq7vCR8PVUWYhoJhBChE0l8RmTjegZOIuqxShN8TC
QoG/NJLltMtcPtl0GX/unHSnqhHUyCDXRO/GMb3y/7tYj4zl/v0Quy1NQ6d6yBAz+LGNkWcSDDIi
xCfX9IVglPkKwgsvs8+l4m0YUWd2p9aw3KPegcdLWdevDYMSqAAWIw+tfIYeeaiwPnmZpr9NyQQu
sBmDn3BbgyZAc/W0ZSp2zBSvpjFf/hqsk9BNHpGkMVeB4OvPVfhTVYerTpvJuCaCESFW8+0Wvkaf
f1DOBFcSL/gOLyHudaZB3Y9kRYnDHKi/oiKHpDiPYwOvNEQH1loVs4NWle5HdnhpxLrE1rRtZ0Io
xBpohD6LrnWLUQBecTXtOl/MfhalZB3Nae7wVC5C5XdWMVIOeCVDypAu6mdd/1Z8e2s2hbz8aUbN
EmmjHbmZEbmkm1KFbY3Fr3sKiKVUR7HaUkShsI96HiK6v3Jd7b1dPH/ZVsOLg/uW1Ja7GEI+kNnD
ZgZSUL8Mw2TFYSB8/r8SjsjFeU/mM+pkCkzKVTyVRpilrPebfAMEfaunfUYLaSUN3OkOrV5V5mYm
iEAsPKFxmvGpuz4WFPtlWme1x2Z5q1FrJNgYEp13rOhCsI7hc5wTUB52MOf+1pQQE4j497Tjmwcl
njkO68TtzMfwQ7iZ6ZAETPP+A7+bNhaWlyh7rJum25Q7s49vmttyUVGT6cAP5aO9Z8R0ju+fXT7i
lZRkK5JzvCohaditCXriJbXERkzvAWAoi7vRDZbGRSBokr9x0T8eLlugjRpqCFNQvnzyWnuW2yuW
J4PnSnyhhFvbTOczwrqyhRLI50SPuzfL+wb0ZErJxjXq13+2WNtfa0IlnVi4YGi6z1WzmlGlaGjs
0jRYNtuVGCeYagAJeGR6FK4Tk04U6Fm2yM+Rk8WryUOtzkfhoa88SJ2va4P2GiQi2XcLN0sFSwht
BbFwePI1be/3ccwAdyGzYKCNRhSYiC+iE1T3sxD4jBNM9h/ML93zPmJ+bU/PHZs1nerOLXmV9C95
fU+QexphL6st6oegQNZE2LpgpLVkJt4CHW8CsXY54GG8CPjcSxNQhl8UdgR0RoAEPpl4nVGQK6SU
AoD0acZHh6vcZaExjfYu6W+hP+Ab44pTqkVnFvwyt3zxE8eRu/BD8Cu9bmTwGa/2eCfQeIsaSCei
KnVPp8NBPiRy+AO133lYJ5tgUNVpJfhtgbJ/gpEgE74gGBmda2GpUf0SyJl76HTBljhNh4ZcLx9e
JfDFIlVQoK8nC+gDMdWHycTFGPJwn2azcsiss+9fbpMDHTm3BLKRCf3kR3SukkW6ec3E2C1zi4I2
1ilkbPj2IUcIx3VLs3JGh47kOGkbPr8kKCZPU5Yocu1mVjL1tZfQTu4eSDQw7J7l3+tfvAlcjvoR
ptvJOCrWemp2xZXaTQlF5fDNlmy8ErGKeBWDEAuKpBKHmjz3hbpqAObAusK+KNqOa7Sa38RMkDvd
Ksq+eiE3RDVYnoSePX91Jcw0nAkpKSBtMa7EJUmx3nGG9VMCKc0KrxO/Oxfn0EOSqVDWINiByvUd
HfzKbpuoDhoM0CRWU1z9I5RC+9Nk1MS2GQh2K5OvavbCylhmLdWB9PPXi4QzGSC6Zn51pQmtw5F3
FQ3mAdB/DSb7CRZ17rtSf2PdDM7bt/RNyI/FR+EX7exp+Pl7Zaq3adNYTgtEtcDCdw4hhNsjma5B
pMZkbAqp8a758+IvYsntMezC4ie+8HWW4UbQ97dPY3uPMPdLl+Or46+vgoBihjLymsOuq0mQQCj8
+AxhmvRr8NFqfHKzuHKYvdUT1LcUJkFTAEINew2ZwQYAT5FXiUDI2xGawEhvZfLoouFOvYGhN92+
0Yks9ySNiWyilU/S54zOiBbikImvxy351aCqgxR3ixGhjR00O/sLtsU9S8Yb7LvilYYnOL+a7j11
Vn/T5YiA6HhiZaJQZaMIqzv9OLNfbuyvq3v+M8FdaoxZHr8O8Hp/nKEFt81PDSjwoAldaMDKKXNQ
+IzAmG35VNoVmWYrMkq3V1KdZjYb2D+MPtakWb6YHwX1Ha772/ip6J0OoqNyOFmo+m4OjdIhVw2p
OR1aGezxtpAmvTKUWFfvFI45ZehUGGkfu3n7GGA0Kl4UyhM66L/YHXdME0G6eKSFoeD6dLorBv8z
CiZu/OfCYAqtY6dK3jRuDRgcvnXdwEq9u6h/1rziX5W51hzn+PJ0bsAdbhdpBl5+X4J4YZ8lsiiT
gvMjah0vABMOFdng8/qI+QyP3PhDGgNWM1TZ0Apj1c5JIqzn0tB0txmf1RFL+fHCzMYideyDeMY2
pckcHGvqi0mRH0L/w4cUpqJZoj9wz69YDpHu4bCi4xvwXjtOQz8zwX81XRxqY5Gk04PyiejEs3OA
1sUBhLfNsyr+8TEJlpLyy0AcBX7v+HQ2/jk+tejzZANRgcYn2d0nd1/+jtlQ0htiPdjYJR8xl/14
4Dfd7mrOXlZovZOUsluhgu7TESqciv8IfFCuWePzdc2Ru28ZcODoabFLFrYEjhqoZO2KWmOBqI9x
9ICAKPbsDGvEVsBe6CHxi0++AEsj6UW7jAGBSWzH3alyAplog/lQUDYx6+T95la2EWHlKs05jaCd
pC+W8nqCla/kxqvwEWMB0tChaEzIYVd+1AcvLeCsbV980RzQEhDw8DctwH4N6TXTkPBWLhrbpbnl
mnlb4xRaM/OVtVyBAU/NujrMpHTFyQ2kFyZWSPb4SYemeEx6oH+XoTG97afH4DaR6bowjhDElNF2
FwdFzBqnQH4Hbw4ZUuVzBk7TV5ukDqYt6IdCQsElhhTVugUANiBsYC15ca+tXVzn20bPm7Ymu0kQ
43kWVhM6+uf1eIoawSpprZqAnmnKHo0znMLHoEXzXq5imz1mKuATgFENqdYkR6CBYGvD78HBjkd8
gg1opI+HJMOnJ2/UhyLc9GCnFojTC5LYQYiv9xN4reGu/G4AHfeDimjBK+vXB8UCTYiymKCAILDl
hH2K+cxie63WxaKc6hoz5DRAeb9lSwb/0xJQkhiUWs4TE59BCL8enuwMBo2IWcNHeTq6j9JHD/PQ
Et9nzbyuSNLBwHGeyaiOyq2oGQecCCcC6tmGti8Jvzd2/Jbx1PjQAffq9uxBJl0ZyTEuqjZ+ag0o
Pd6hYLBTOiAZzuJKXTEBsq9ekamej6kFKT0V3YlvocdfIZhayIs3xOIZtCUzoS+lhI2Ss4cOd1e4
N7muDOfCQ0V9rIDaF/NdYTzu+5hBNACVRihefSKif5UKB/f75cL46Opx1PnoAVb9cBq97O7pFZoq
AYCx/jrHzz/1AMb/CIXplpjiHQ1/LCIVrsxH0Ju6n3fLnXl7Lx992ecMUUEpMXAjDd94hcLokfJw
RU/Z1qFUqDb9AGfuhx5sCFtVfBQ15kTAZqlgGPVMpgZDlzZ3mBukUzrZbqzy1NNdNmhdaLlWE+u/
PWDflae/Ny8ifpviehdmBy+D+dF+qTf2O7YcbVJwd+lltrQmEOBblhqStk6CjPoyqC+yaLhQ5KKa
ywziNr6J4HxQfb65LD25c0WJMIDnqx29yTUtmD9WKSuEhWS5LfrmPvtK/OkG1tBZqLHiEONEOP2b
q79gXGlezGv/bEFWZi9OrcPUUuLBZCOg4SuDWw7rsCqHUG/MbOFWa26a/9XrnI+T97aVC70omQjC
JM5XMf9Jpxmwz87bT55KtKAjfPpCbHqVWcP+yQUiYbyp80iZyPs7/Aod2LJiG2NIUihF9MGoR9ka
gQIWYWnlgHzmr9cnrvTCgsXA47tz6BX6dKc51Em9jqrL1pGIEn76ZKVynaiHgSNG/y3ZpGRG0bFg
xGVceYffZsTv3zscmWqD9AO5KhysQh7mucV3yuCt2PlYmP8LAQysDUUMUITo1YgVYDj18voXcuPl
4Y8bjH5g0GyYEBpb9O8aTCxYhavHXBEF5eQb7YIYirbJz947Z7mId8QO02Ilv+ZuDPsWuI3MiO/w
vHyMWElLsC1lN5goPMCIxfUg1CvyzGYgpT1yTTQSRo/y1v4oMkDZEi+/9PpGqqLmH4X7UuUo1ji3
ZzvZRN6C4nASxp2d6HDhQgiYy79WJVfGlpWwSSf74xgin0mnn7u4vcRUlRVZzRB3SaTHSizKWJEd
Ckv80G4tIFzXdUbmF6HHATHSSFkxAaitp64eDv+PpeCcgQF1YyeokIrBIvnJUYXB8sFdtvA1E+EU
p5FqFTBIOPIf4rq6GSVW2NDaz8o+ef92wS1IcMUdyDfSmGQEjE71o/tO+NisFiNTZ+vGuzEXy6z0
cczSXZLsPRBmQGHu2RhRde8r3mLiw0I41ZflpHeB1XVH8fCrw+6TgvPAAuYf8K105gXUGJCD98Uj
0bRkAYN/peYU0qHhfhVjTM2LvM5Skow7Pn87kFQjyPSIEZtXj30XEhAPTY1Tu28H/H5mAib6gF04
xY989ok/fAF54sy3rkTI6pXjy5vpoWPfbte9DJlRH/omDLXzaYUfmSsBAKyWKvcjeS7tKXnV5KyS
WM14bB4Xq0eHGTQuUQRHaHYF1gDiluPwUpE7D/V4Af3szMtyU6gwiF21lIv9AesTDDaYOSxLJNCk
/rZn8gAIR6Fn69tFq7GvEocBBfElVzRcPJfIpOKPNUZBQ+PoWSOpKbXjinIW53/LCwVDTyVuPxdP
TOWXoEDOk/QjZ9me4yJ1CW0xAfJkMjJgpCtu3Y95E8CQr1+7RZnhzh7PEKAnORgMyx/cRnxIZ7lk
OfOnLOnJUTgJufEpvA2Tl6vLTWsPOdTb+fEtqiXdQIb4MkSIAEGJFIULWDmHyEZ3kZQ4RQ1LW78C
TRIgE5EjbKoDTAmqm8vm5DKXs7WjHuBK/s1Qda8kFSBjvMQKNTUkZDPTnFYpk/RWUXy+oon6JMp4
mIT4et48lvCbc4uQ8u3lRN0GV4Q3G5P2lLJJE1iqL+HfCoSs9o66GcqTtqAmO9XmnSpKMx7JvVzN
EdTMlhBqg+acguSz2r5FGiESiSs35BuO1reiN4g0nX/eiY38NuKGDSb9OD4p8ZuvAgeWKrDxS3IO
Wupkebbye6eJKRz9AbDodzlXXC3i/cXnQnIYzGVErQZsqr6/yqI1KC0E5gIhujlM7mCp64izuARM
0mAcGAVbUC+CF8fpqihjvVkMtZ6wVRLn2ztqvxMvd20l4RfBOzRkYwSPyA5hvlguszW2uhrM5QMm
zcbgwM189l2hieJGjNUGnd6PQzwGWXMFtrp03FiJv+iIrAJpJtxiIUsGhfuzUL5C9mApyQROZ6T6
r0oZAdKEy5PGf2/bgBcGYb6RuBlJ9jkErmIT
`protect end_protected
