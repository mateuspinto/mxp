`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
bZTSX1eTeLRclfNmAUAR3R3AaRgVsWLHNvvLKrwF69WQoctc3sC0r8IYpo+ScjqIC8CImjaGvdNt
r1xGG0wcn1CTvck2e+HYaGVwGzwEkCUzXYdFLKkvULERBG1Dz3dvHsMltZ4QgKof5BbQrdN9E2FG
7xaJwfkwbj0Pen0rA+I1ndH+GAFJ3HmmasthmUp2uP9388bmGkn5XG7axdHqC4CnHOnm1bS5lb9b
DYSgtWmjVVcOTz6fsBB08rZEptHIe8wSp2y5jM/CkQQEVv72Ma2gnL2SKqzcDlrZeajIsdA8LHXe
n933kemEirf2B8ppLId3UQwk954vD+iM+/FGD4pOlKtRHPrGy2SPzLqv0m44qIshv1BfvYAm3Jfg
CvNhCiUqQ0jK+1haPfQ8zHRkxODpO7U5WkNGs4XhmCFqmUw2E6le9pNUlVjt1LfRlrV5+kJegi6m
DpV605JPPUYx8gmSE28Rs9zMUh8ClPJ5jTY8upCf0EuRKkbdOfZd/l2rehx1/ToQzzdIvt0IapCB
UMGM1zBqrxwosuWBI7sbP1JRSw8msNI0tsPKmnubXAA136tGe8O/tcd4UBn4gQQbFXxcQyPnru1b
iZHseTF5CeDL1ppPsZOdaPLGuSV08FOCEshhhFjKIidx3UTpcGuiswalFJIh6idNy3l9GWklamHw
Kpn4Fm4mQ6Ypmh+RN8VndVjFyRS6w2v6GeLTTrFeZ8dqyijgsck6DKOGMfHCedY351/vHdHXtXHu
E77KaGpl2/vDH9bILT0PvSFa9b0cH88MVkOaUTNIqP5KQKmoszkNoln0r7wIXSlxDw4y8CWGuRLv
mieDt6vh4ZdeAN5SM88IbGQRTaVon+AehAEcQy8X4nKo55dO/LxxaoHGijKxvMwT+gC97p/ia5YM
MYA28fdlqg8reHk1GofgpNQThU1snYlpwSPj4hhcejtfp5QGKW1gLbl38C1jDrKtqmmWiyEIXPET
tKZc9LqqKlQB3CbrGDUuHd/671QlQZS7RV3Ek0YVP9CupK3NQaLVjt5GjdJt++zB0gXKRpYr1AmE
8y4x45fnMQ/ngUtX4w+3QBRZmN8j6RUXFp49JBpwbxrD+rZUZPhwUCtab3sas6KTyopyXrN5CKX6
VteG3RafQFfYJn2nJXRd+YWYMC71oYaBLFcByJZCkn7Yuj/+FtbOCv+KJSjS8HFtqGwAeLoesilK
A5tB/EQY/3cwO6aKgpNkdlEABW+tMBcHHj36m2HP9zsLsbrM6uIZF9clQLGIjNxDcJ44H+bRdMFS
j9SBuVa+cDqRr8cmay7FfIuYz++zhwVHDG1V0BTAuLvBe3BVPw+YIfHqOX/pDuU9gk878oPWS1oh
4CwBeX8TceKkoB1aQA+BXAf9LnKUztHVP/WiMphhdWfbFiAYcxiAfyQOQVq8o2CC5XAGe2RzSVSB
kZsmZv1A+b/smlu3xjcxx6OAyRsrJOv77qmkznHb/2gyBlr7eH8ayyp0RGuTMvVc00ctqH7qeCq0
O/nKDhIfHPQZnxDJyvRB1cCaT+ghf58OUuuMVR1LQqVpNQivkoGkU1JvrUeHIOre1jKTrRXIrdyk
92A8QtDQinAQyJb3zOePprMao8AQWF57IFXw8nLylM51G8/pHRGBT/FUasDq+yJH+0nqFmwYfQv3
PkjZu87QH8H3GzA1NzL04BQu3FDwdwWwF74FmXbSccSdlEmCwYA4lMDX7vpEYedpOCpzKEzlA/Tr
mdQnthYfTYqeAOWEaqpd1nqIi2y8OW3xYXMZgZ3Up/xfxr6FdCQWsqBuTt0XJ05WnhXY5VbwRJfG
qNhBBR0Hne9NuIBLO+dEfNLuuW6tyw/plHbUaxayvMz56az4QfKEexmfW391zVSBmB2r3u5g52K+
gecgVAT5uK9Es1WXR/aYiQqtYEdqXYNwDvIvvbMHQDEWhWPZdl2AZiDpqJhR4fstMLqY0+Wbxii2
pGA2H7naD1zP/pywsJgAY5aa6e/XPGyOEoh3eR23k1ylCs4Y+AfHe74wfBICQoZRL6XPzbYTrLta
QrNspaQkUYf2PLQyyA2hvMnh+J4tzTEc9xy/KOigGRAO9CIy9kyobepEQ31Wkr6t/g1k2FVOyXl1
mheBxDZr01+Clyc89k6MqFnvl7cdHc+bwDXTdIdiw3/1YH7nQ01CLWj3sViy4VYYUSyFXHhFcP2H
In6ZpRzuWeZHMHzeClq2TaI3nAa1qo8NfKN5itpbapC8QzSIQkaoswCJG+iMJzREFw7o0pGyrvXn
FZnIlmu+an0DTFEC/eI+Rs8qp/vp0a0rqGPlbxYAyk1RN75BINBatYkiGcmEQxw343/nJjJ9TNpp
Y7+UYG3RZXLUIcVzdticmEXybEb4YqjBHa/SE+usR+1Emqb24QgCYhOaKIXWBYgw6/VHnN+NEXPb
HlUVlidUmYvHQoaD4SKkrZluqpz+wbvmjC6F44SfTDS0RoITDkuDI9YxcC2n3hMmyIshPhRo1bLG
OFYMC+hG/stDsH6PMU0jAM5pFxv3/5d0FaMEO4Tu8EcLZBBPXG73svW0PDBsTeT2XpN8mUMEii4f
n2PjIi4rh8SynEjBKe1DUvfvqg/X/ygoT9AeAYEfzlmu0osd5G4lI+7i+HJmMZo4iWezGQXwEoIh
xJR9zFz5FZMzYwMfWzLHBRIUiRX/QJ8bXNkSD7V6bJ/501sWRPBCRzQgRrMHG301RRIi9z6KPBir
IvM1NsBCQmnjJxOE7308YujttxeEAkrk3cVPsLmBJeHO7d1AR0TSdzPfKrRxa5Qq8nbGj6CMNNZU
JZcH0OOqnuoxnI+/qHS0OignYWfyfJ73gcZxDBJtqja41x8T+N4qTwBRyNKkfSGyCWMT26qUbpxo
8vxqO8hzrGkS2r42THa7SHk1Qetn41PKm/sB+2bxwunPy8RMU91tHg/WaGsuwX7TGgSQ48MzvERl
obH+kzYLNHSPZY2MIKuOxhSEXzXpi8sOsHDnxVXqUF4LAOQ58UgUhWQgJTZ9kIgbWYmRoa1NAK/J
Y5T9fTkPsS0OCpqpnQuH38fjvBhE2TMLQtPX4PlIrDdVtLqqUYF1tDF23H/HjBqMfC/ZKZCZZGTq
OA/9XCXOx5m9nHtFk86Gm+PhI6De+t1MBACOl/XQv5WhjTcFIsDyG+b9hLP29b4CPw/xOwGRNRey
UVfjlNG6hNex02GoWTx5K7EgJeKb3wymZoEniiEpa/3KZQ4lI1yfbbVwIWqj9ukyIPtfNkCckNAO
b45X9Z0kTR10Tm62EbR5TxAJ7ui4Aq85e/Y9mtoSCksahjW/wZ650i4vpV/2FN7C1KFREyWvFWXG
TEjPHMPbGYhMKw6G2we/mbXVuh4rkwOMf82HCRCY1JhBVoAH4XLOlN+v54tguWRAIc+eLADt06id
zpCP961edLKNWS1AQUzaLrX6OeV6pJ3ZgTmwFXe1UceoEV8ma25Lonkzhy/m6eslyzHEm0bBCUSV
6uwfAK6mxw94ioAbvDtQN1eZS9cVw+DmwEZXslXo6r0Q1CMruoOA7rweIoc8GYxZRqv9TJC1iBuo
CBG7qJE0r1Mo9FYV5H+G0KRAfET1u+r4QinWtDT6E/2t90mbE3A24woTlREI+vGoYpNJBflVRm7G
ucx/ZlNfuXezInHQmjT/NDGfy8r/nm8VxbBDiPq1FmcwaS47cQS2xjLcyWJxkN9G0wjv92UlQqNY
tmv/1e+EqnkAF2DuF4IDwS2lY96d1IkLyyUQtjzPsJWZE+G1xTuEW9p3I7PYGYRwpcw/YvOO8LDl
XgbvSOR9TPLuTXYJNKNyeMFzzkvvMSk2eEljRgYevRwUr4dFRg3TRs06T+APXMLcaF6mshU4ravF
+YqNFYp1iBk8lO537g144Kv0BlICrOPmHNXBjDiVm11xhGpqLl1h0M1OMLfNe0tJy6L1AyVSMdJs
GSSTICfBplldyBBzfxgC7iJjAovYXMv9epZsalGcm2YEPw8j/Y4RY/JwC7R8gIGV9dp1UV7D2FaK
hDLLOhGIXeTtDH5bPEBKXt3ZqVz7svuRdlvuAQtyJBSdI4VCsboUr73ov+8O/iq5cD2wlZBJDNAk
/tdWIW0gu7b0pOq3g2JdKnILAUrpdgNSiOp9Ae43EQLKi4ejlGexgGApl40BRWFtkw4U5b2++v4W
VKOsEyTVmJpNqAEiEv4L0BaQC66/+5QeLv188zwPl4RMYuQvlz3VfttKivjEkS+9mtWW1DDmACnw
Bbv+7NE1dVYGrvNFIa83S0RGacPuRxsYn9eOikfQgMOe7nLSJKKVNMbned9qEOtnbvVi+Ax1WIb/
ou6jEHkd2oxHl3zaKxkWSaarOyDnlrtGbz+t/XskleBtzFrVO9pFRnZdvYSaUbOUFbI2WW2bnXzq
1X3E1arpD3JU5XyvRMpMecEKwR6nMReCCeqpzj5u/kaMYtlplY+NY84h/B9qQQTHhpLLJnyAwuqO
Q9DIOk+tMBsyd/hRbU93rW/SjC9tRfxjCbxV9wsWhKtTSF4eZhuW+SohrSHPaqWTFtG/6U5JbfSj
3Sr4wYxhOuW6F8gm5MiYgYAheCGrYusovNv0ZmdvoYkpM3IhgzLk4wr2QD+oOjPuvAheAucegEbo
Hacz8cubm6SO2IVAaudhW1+SRHPTchCtkzmceN2FjclkqZEfpBKUsqbDGfBmONOhMPzClLPhmhtk
+7h5c4i+uQno8n1du3+uo3Rq52dgwqR2R6W+a8TvWWWngrWjT5zrOTEyQaVQWp6C0MNs9FzrDQmT
Ct0FlJTsQmF1I+lcmKjshmDL8SRjGbl9/IBGdxAybUOibKEh1/X/+SzgCP3cl1gohXWXaNce2INO
AMV+D7XCjcI49+L+dbhXIFiE0TOjittH4lNMxaPdBNrh3PYy0OHRs71xp6guNC746irndMXGQOkz
jkJ09th+uMma3KxwIftNaMfujEGQfJKKiw48/OxtMLR99P5MiqLtbTvoLjBDl5j58wmoGoAjh4hk
Zx9dIMS5tcLijws/PtVMddRujQ00Y5TD1TIyHaQo8HxpeFBLD4l1YIlgFxtsLpOMawOWxnfMhUj9
V2ebMpxvT0YPEoVY7vyBpwUhe4ybqhTcchN+iRJQqYgZ/Mms/G5O5ymSfYDXvRYZLHdiO35BwWSY
tELs+OKbk9UdlLvyY9dUXg2msJQ8hAEgysZdGVQMf2+0AXsIuhgCs5bsUcXlQKZCKAfUmasxoH5b
JQTHgN1GUxvYPZ4UYv9+ADtEs2fIFmwcDpfcvdABv0F5rQ/6d7BJKp7vCsIHsfnqxRQ1z/1z1YNE
52BTtlqATeTk0fmqZQRir2b6pGaggEhj7QPgH43GmGu3G8ZgMocH3d2GCSXA0VnGlrx04DLImnEg
IvKyE49ZLqBLf5atGbpDPT4NP1FMeNjhBsPYmy567ho7LmvWji9OcQ+Oe3LrwiJ3h1vmP/yAcusb
2fIl4wpNMsfRizUbsgoyl4jNUpmyaYoA6niZnsIA/f1VeQbyu9PymluQvug00lqwcgyXPoVIaxdy
3tDQmDNi52comPFWSyVwSeam7CswTuuRJoCFvhG9ByUb3XpOYlRjdBAQx2fu3xIowKF4a7mqWjqY
5+6T83vn1cI/wIun/JTfOD1hSCxSOvUNzbUl+lA7sRENxwhxXQuWEs8XH731UErmUR8inMxp0Ox+
mf3ZcmfTbqRMXJ+1igEhrg+d5Sa6cEs8hlPaZOqyV93iB8o9khIQP/XxikiWinz+oWguDckgECMq
BO7HE5Oi4zpuYmgcQIoIipYxSKUNda4B2SGLPXfxijuNOEM9e22Sl4zZBu1syhGT6OZb5Dfutmq/
ZVCnqkVG6rpCSwn0yvC842XkY4Py7F5juoyLMAWURpUzluQWCLGWOinwRfeQQcH10hXuyl4+M47n
UDkBA+lsLNvO4iug15/mmvZC4ovdv4vOBiCj+lUGUdupQdxt3hcPEok2e4OQ0xXG2KIdw9tCa4xf
rfNPoFGi40s1a80y7umqqiqUr/NpU3Se5NsJ6KDfBTuQUR6Qqa0ka1YL7qL6IvJHXemsrSaT7HCu
c6cms5LsExWixDFr4saj6uXrFnUJfTqEPhkCgXRCl521KuIpzUbPH5z3nRVmdfStwPC7MM3beV/n
CzVf/KH8hq5LlKd+NK3JlMfdf+jlGEtdu7gd22etnp8iTkXg3HOojih4okQe2SEpJvLtiKBvP4Ff
HBWqn96xwREVWDzEBNSpSh5pjECLwg449PtwzI4kuerVwAtyMv5O5sr/50XktVau+d2AGpOY9HyN
xjtefWyYhu26eAsdaIwqw/S98rQY0vX657IBS7Ka3tqVowe4YcdklhAjg1mc0hyiF5lSucCef1tK
7ux/wfw/vjQelRO4PHV0J5MBIan4RVuXAcAiPVzIcvkDGRMlMLAQyB6+Mng3eKrboCY2zZtlmd10
E6ZE1mww0QnuGGW7Uwj967FWk4gaGwvje27zpZl0Kysqw4PGtOXEpIdM9+So8tY8CsFLOZ8GX1pK
5lxYa7K77W6x3iH4FvR9f24dIIKVI5yTgyctshaiFqYHslUlpxEA/m8OXVip0HFVZC4qlLtbPbz9
E5bRh8iQ6iNDHWybkgLu7O/q9+pPfPGyuPjWVq7iRGHDi8WubQo7dT5ySNIBfRh+k2afMC+y58ka
aBV6KYVTZLItAb3xyUgcvGuwACuirUuo8eFKCNEUOullgiL+f8Lp6xM98lAauJJRhZMWItzGPZaQ
rTytlW1CRboj6Ux0GfKtzU4bVPhaM/Vdq8YrVu+kyoFasHDqJKTq2Rcx7Hjk5xx1EZTRyw50ohWx
SThyiIxTlMRPkv3H/nQu+f/7HCJltx8g9fFXOEutMtji82AG1Qcoi3k2Uq5xYkGg/uou4eVjjzrg
Hr/NQWxdqOlZItM2hdReXFfKpdfmbgUL6LcKxXVvnMM+CleH1KaEVJQe74/y1bJ6t9T0PVwDh7mw
ZLZVTcNnLN/sYsHMJqianohrGM24+w2zOiUp+w/HwRcmYvdB0oTQUkXLr4Ej0hmRqKZBjWvBjHSN
r94nGQWYIYRus7fVpIRYH/sLBzcZxvBOd7l95ICnrF+QmBYYC+KfqivpNEq5ma+xmuvrMNRGWMBq
3Tb+l1ZCG++rshv6P3sO+PclFRCNAxJFHGW3I5fTfZBHVFtI1fX293BQx+vxWr0NxiyEBCHYDbNr
YEW0fzTYaUu9X5p9kqCzbEP9VV0kp6BJBIULy0Aux5KjBCvCdlVitQyoVdxdn3+mC2rVwkToiGhw
Eei9xeCNgrVUDjmccGpS/SRfuZprkGVKoyxn2kLouRDslcrJKID68jcRQlVUZXWGtEDH5Am9ZBbb
7j2M5CtwNc8gh1iY/1chMAzAukLKzN9a3tMq5h6PhZ7Ll9MzNFSGbHKF3uPy4tus4983YcKW/857
3KI23qkvRFVw7SFbMwiYFDdsCEPH1bw1PkgB8sX14waq+BpQL66tB2przzcd2dG/ASm7Rq7siyWi
S/fth3X4UYvzJMUiiZPOGP6Sk6z+2xwn+tpH6qbHU3L6s+Q77jLxnR1cDb8Fe+XCKqWYX0PqDc1l
6UqCaG6gtm7gUyD9va7mrO1s3LKzhC+PnFu15Cz+qIrdHViulfdomVxnyeMMfUCh9PyqOJEzI7N/
8jWG4Y7q8HeH7ec0i93LKLB4oB3A2mlbn4XAT7CkIl1GT4VoMW6aOlwpiTK/k3bx1PEiu/tmeW1a
3Bmtj4pVNVJ7N79uHjBC1NroWdc5iDJ0XzdQJfiSj6JPwcTkjSRBaHBEILxObtr5eg9DNucxEcPg
UKZL7A8mHfpXDB7ZJIC/IYQcOZLSwcsrLmyrIKfDvOacWEA427sJ2OzdxZW6OYynHHlakqYgyjmj
55QPJB7qNfd/wANhVyfsALnEYGKAS+AX/BdxEpZVS0R768HJo8qwSr1gnWALHypts+ulEIWWbyfS
lWT668CUJBcNjUSRg6zEXDob2ZYFENTqaFRmi1gkyWKb7g3Wb170FPm3Y4SPzMY+X+om2BTeiQO2
J6Bo5EtVoCzCxEWEA7Y8JfYZHJchGStgPfjLP7cLcfCeQBeevYSCPlA7tEEX2Bjzq2D0Bw808W8F
60+HdwNgnbtfManWGs/WXpeHzja/EptkYKJRtr9+i7EdMvsCUP3DynfEo9ZlIIwvhvVY0s/7Gmid
O2tlwktsfpb4Pqf2u+dnvKXXNn7zY98gRCwfXH3eKvbbw/Kr+fmU9Nm8XwHzyT/Su/98esjrbOIb
4m4C+w8tY6nnMMMcyooLLIwQuAv1yhP/FGLCbDoh2O9jvRf64M1BQOIxOalHxklOBl61DK/SVMM1
XICsZ2AduZi8CMEOyt0jIOpSG2DtU0k3Uma2SZ26bhHGG5wbcM5nD1NGJyxRoknhq5B95EE0EFXx
a5Qc/uGg+7Cm+TzwCjkG44+L/lPejglvN1Gb306Vm08yacRT5K+FkTS8giTdJl3uwbwUfiwqgVLb
z76ibI7ncKhnGCRyxoITmw==
`protect end_protected
