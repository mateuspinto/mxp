XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��	F���"���ۢn�89CH��1��)�#�݄��ݕ�
j�` �!�u���5��I�������q`Cy+*�Qo"pee�d��fM��|��s�,���U���b��O$-H[Z���6
"8�P�A=���0�f�\��29s>b@�`�E� 1��Cbȹ�*`�$�R�Y�/G� r��4����6U���~r�Xg�|�F�W�&�X}$Q�Q���Y0�.���I�9}1��9�$9؀t��5��z��RK3����h��\��=��!���2AuEt��>����9@�8V� ���u�
j����%Z��\]|Dts
g�Q㞟�[�����Y��$��mE�������v������fT�F4����q��S�ΓE��2����!rYH`���8�=*���x�����\�KK\\*�k�4:u#>��%]"��keV�?+�l�ta��خ��� �X�+�(�?�����)S��d�m������j1��G���"՛{��ɘ��@����h�*E1o�S����k¥������ס�sRi�������� OAȩܭ�]�oB��4N��8���$ö��KN#u�O�L��2LC��k�
��5��{SAZ��VlV7]������o_��"AT	l����z������_z*VN���J�0���=uz���N
i&m]���8�����{p�Vr�'�OY��,�m[xꝞ�eqͿ��>䧷Bw�LrdN����\"����рXlxVHYEB     400     190J������if��y�^��6�x�;Sw�݂\�U�����U|JW�%��18�N�@}@�
�p��v�� �qqr�V�)ic�!��g<�L,���~*������`k�U�&О)ܜH'��.'��ME�Vܰ�V5���J��#��?��Ax���Y M�@K�sxpx��$�"�I���
i2۫,V�9�,H�a�0ͣ�*-��A"Q����/-��w�:�`�׹	�jV��5�B�'�c6)A:fB�$.�� �w{@�$�{�h��q->W��s��}o���c�I8#�rol�W���Rd��]�I��/��M������hGP��<��;���]1d�Ǖ���=G2��h�jS��8����d/+_!�pJݺ���^�����M��XlxVHYEB     400     180@/�bJ�1��������,㮣Ǚl׏`l+pIb��m��i�����-8�絈f���;��< ���ia�/`R�ӋeG	�K�v2n�h�E����{	���e$�1��咚W��P�y�[�iu.��@�*Xȱv�IIs9)��)}ݭ�8ai�{�����*_�d�>E�	%��[!�G�>���a$373b��0��4�2H[���g�g�X7u�;*�w+���&KK{d��A��cP��X,u%�v��X��`���? E���n��f #wR�%�*Je��Com,2�?�R��]�^����J��jM���i�wµ��H+O*�k�R��H�������D�d���j�8rC���=��XlxVHYEB     400      b0�`9*5�t�XM���V�xH��uiٿ<���_���
��������N�QR'A
/�b�[�^��>�҈i �v����e�^:B�J�uv�kD���EMX��D����l�=R��/���廛B[]�籧S}԰'}��/�!/#I�q<��S ?W,'IV�{�n53~=��50�TXc��XlxVHYEB     400     170�^%��9�.��&=%~��4b�:\6"���4}�VM`GD�q=�!�x�Q�,p���fc�'0�J2�T��_����*��/�[���i磓Q��Rޝ�!�؝�@a)'�^|������j�;�	e��51?�{��a�RX�	�[Ѓ�V�\��)!��q[1�'��ê�rv�P{#����q}^�3�U�ό'�
��A���gEH��"���Z�G׵Ϋ�ϴ\�"a�0�A���D�p����	�L])�&��C��(�t5mDR��C�HV|c�����7����5 �~ix�:y\�Q;G�N�Ū���1U�����5\����
1<����~M �$�>�ѿ���˞�����XlxVHYEB     400      90�@m"�)
��N2�q|�y7'سQ
�6&��PZ���=����;�����1O�@�҄r�� c���MZBA��>��6���$�3�N���4�NE���ŜLi�? Y����Z[4�m"����L{-{�Ĺ��XlxVHYEB     400      90ǀ[�H��;oJ[�����S�����!�ӟ�3��K�OUV����`xX�7�b4�ҁRO�r�>��*~]�Ty����v^t4Zɢ 6�	>1� ���<d��W�p]]�{"��13oG��Ty�Ҝʛ
J#�~Bo�������,XlxVHYEB     400      90؞-�M�62���z+��$�F=!&q�g:�W"j�t�Z�슣V�㥊TV��F,�,ku�~�mU8��y�J�S���hMwP�Lb{����>BI^���J0��q-s�.��q�Q��aDy�vV����=�X���XlxVHYEB     11d      50�X
������ǧM��Մ�?
d~A��+�i���6҈�1��᯺�a�F�t@
�F��6JS�L�`�؉�,�l֨�