XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ʍ�@m�Y�`BPS��a*6���Λ�)�Gy-9�� �4��E��*��w��Sc�'������o<��T02�t�����]ĭH����If���t�_g�c:����E��ͦ�S*��g�[�h)��"����o�CD��e��j�)��7�`������v��Ƅ��e	��F&+�!��$�x}FC�����: ��K�
6۔k���>)V,��\@o5�m?�z�J�����0��ı��E�xJl��u��ŬT����dft���턨g����-��>��`��X��u�ۨ�56�>:��=�N�U;�x�+�ɠ�[��7�T:�T~��+��D�K\dg�<Y��6DQ����m�慁��������!���$=����6�y�

YS%	��Eόw�?IDiӨ��I�ls�p��ce��<-���������X�`��)ܴSy8�-�va��"HM��v\/��K�Q��J\�Jgy]1x/{C�(O���E�ڊ��W.m��#�9`vP���p�A-��Z�g�wxk��_l���ƸT!�>�ƶ}=�=�xgW|��U/��u��6��[�,WLc�z���{BC(�߯�%�G::,K}��D8J�`X��:�܄V�Q�ڦ�]�χ�DXO��ٌh�����צ¥�#�����g�3ai�_�I�<ǼImkq�wI���5[�aw����Ҵ�Q�T^4;�/Ey�#�4<��y�Z�Y��N���b�	�V�����%�������D�XlxVHYEB     400     1e07%I���Ȩ��g.b+�B
�'z�0�̾oi,���4�T�W�r��b�;�z{6��-dӿ]f#F���!�o�S\G{-�O����ݚ�h{@��j��U���=�jPr(�K���^͢�E�}d_`/�tc����������F3ٿE㪀�CH[�]�?&��^j�[ �+��
\���l}��83��//�yW����*�&Lp��.\��VW4<�J��oCRG5[��|�&����A�"��n�7��_,3���w��Fw�ć�N���,���4�"g�uc�#�%oM��N�k��=�2�lꭏ'E�Z!t��rG~�ҞT��weY�X������.|��.Gp�>=� R��Mx��Y�i*���tReZ��X[�gG�)w��|#x���3y����)�9uN/a36�s,Q8���y��A��ݴ����8���ð��*M4�l�י1���L��ߵ��g��I��fO,�qXlxVHYEB     400     140���Q�<vRs�)Ha�5��7��" bo��K�/c��`_M��E3�:
��l,�>��9���T�y��r��&�kܱ\�����Gyu}�t ZZ醦�0��̊���9���o�V�!Ɗ�cs�I@UanE2�ʶ�#�5���,?�d��M���� ʆ��;-y�v�s�a�gr�0l�$oc�QH�����l
��>���~c'�.l�]Pyӿ��m8E~���i|ӇMq��:h�)��D�Y
����>�k��j��G��.���d���A�U*�{á���5�9��z�E�Xs2ɷ���{Wn`\XlxVHYEB     400     140���|�X���K��N���6!�� Ɍ��	���F�~q��d/����qB���X�����l������x���ܻ#l���]�,�&�	9�oU3���I>��I�Y���/\�-OT���b���d���*W�`������ ��`<n��-ɀIY48_��A��C�չ!g�4��Ȟ��t*?=#_���.e!\����9}|#����6hɰwҸ�ԃ���O�&����^:6y�U+(BvJr[�>����0�`���q*���lF�i�!AHJ��{��H�#�.�wgO4��� �N�\�Hv��x��XlxVHYEB     400     1a0ٞ7Cdm^᧰C%�
�6Y���{�/kra�����ל9U�������:�b��S���@bo5eD�;�'.C)8�&��9�j�Q�^f��j��}��}�������i�T�s�V�tW�B�?;����V~Y5	�M�;�9��V�s�w|��˜
����ά��3���a�oK:ڊg��W.@ko4}��%
e`
a -��a���<X���^8y�B�p!���-��0)�ހO��@Y�-�w�ߋ	ϡͦ�AM����k�@ݧ���v �q�يPu�-|?�V�������A���(:�?�F��k��qd㹜-�\�v��M��p�x>]��3K��=���g8鸩F��6�fc>����d�J9v��u���	ym2+`C`E���tUI�{r����q�XlxVHYEB     400     130��L��.�N�	D��Փ4_���fĴz��D��t;c��*��N��wjT)�%F��	��*T��wb�\�J�qc��)R�D4N��Q4�Y�U����F^x��&)'��j=N3���L�@�y#��pyG���Y�ǰ-}�K(GBi��FL��1�4O_Z�	j&"&�	�-���E�#r}-f}�,�g�:p���q������W���k����Z5��s�pAm�AhG1�����\X���>e�+��ƫ���u0
8jA:��󩔁4b�`��=^�����e�Z�3���i6XlxVHYEB     400     190"��G�w\� $t �tR�Ι~��o�@՚0"{zg%=�`�|%����A���3�b�)v�?�~��SZ��m��b�,��\��h���O�N�g�ͧ�����:u�0CnAEa�Lԏ[1sH�q��)�@��s���"�7 ��:@oۑ�����L�x��8��2ߊ���n���lx,g�GX�N���z�����D؂���;��2�l���p�X��s�8�xo4���0k�D~��Y`��?t<�x�Td�B��fr�]~;�?-
g�^�*�vЍ_���LG�9'�%�ьK� �E��j���(�h���)�*?����p������
=b͗�,�c��zt���������HA|٦���%>/��z�UA��}r���@�XlxVHYEB     400     160?��Q�����F��_���=�������UU�b� ��U��}'V�4�H��z���X/��b@=t�+c/X?�G*#�P���j����k� IP��\BjM�RԜ$���,���	<� 3��{�-�9�C�'������T��|�4�&�
����&�D�\����M�b�<��'d�@J#�Y�8A{��ĳVUȳg,�zV�Ǣļo8LND��7�7�HK���+f�@ JMIV������08b^��Ttg�(e*go�!T����t��Ex#�4�"�-����L�~���#�շ���^\���ua��-b�1�QSb�������~4�0Ӆ�X���XlxVHYEB     400     150��,�"#���N�	���:��AS=x�� ���pI�N"FN�U�q?��9�e�޿�zz}(�gua(����I�/��͢��g{VP3Ȃĵ@��I�a��k�c�>G�B+1�G2J6ѡی`���P66M�����߲����(�7���l�)�D�i���H��Ωϔ���3�*-K*��#x��p�9��X��<���YN3!�/��1Es����	Ĕn��-��A��2���rB^*����t��X$�>�����f���)�o,^M� v�����ta�ͣbF8�8�*��AN����^�m�{!�d��%I�r�)+]z�gu����\BJ�XlxVHYEB     400     1b0���>H�>�۾�:J���7[hN11"��5���f�t�z*5���m>� ���j`i�\A;���ʟ���B����\�a(}b�i�OO��&A�##��7A���W�<��Ԫ��kTz��W{�AW��3������)�%,%�%��ś�W:WL�,e���Ǜ��s�
s6c�Iᾔ<*]�r��/�}}RC�/u#�v1߶P�*���Hn-�?�3U��,']��W���j�N��c����~�Z�2
>���AXj[P@�&(H����1�C}ڙ|���&�1rE��Z"O��W�0�q'��A	EV�[Q���[x�5
W(^L�-6BZW�H`�%XX2�f�����*6��(�m��뮓�v�D�`]�]9�4���i}�iN#���ci���tzHU�gU����+�ETXlxVHYEB     400     1d0�8$2��9i��}(����Br��}+��r�� �N;�}�e�"!]���]����8��H\o�S͘��m:-�˂w�*�w�&]s�"
�aSJ�"lX�:�`Wuq���q����V��7Er'TIj�! c=,6�<<ѸMi�N�����լ�;�nښ`�R3T���Z�����x	Q.6�,d�D�����_$;S<�,��+�J��熓��ܑ���2�]z�	(��FLD����L7i.IIffS��m�f���X�s����0�������m9�و��S�y2�����gvk�WϨ��R��Ԏ��t'N<�P޲���DбE�{�ﮌ��7L�"_�����A�:󮇘�4<.�c99�ż��;� �((��V�,銳�V d�4�y���,�s�����&� HS�۞���%VMHJ��?�?�����fG�tj�[=l�XlxVHYEB     400     160N�huU*Y��mޗj�	+Z��M�aD��ot�z�&��r����r�V׍�F�Z��j�j���r�x���������{t�ݹ�"�>-�"^ʠNP�}�2,}��;O���3�/������a��Rx��؁�dՁC��3��L��^���8L�K�Wh���K�N�-ߎdp����|�Г� %�6=��|T�Q�B����9���d۹ ,=�SAƜ �1���]�ѝ�$�[a^����$�l+�>`��� ��+j����O�{&�����|K-(ܟ�غ*!��;��Q�-�֝obG�3&^F<J���S
�Ѷ���{U�U;�+�&�u΀#������;�XlxVHYEB     400     130��o�̽Z(#�T&��^A&�����[�7�)����~�ُ�=�ɽ���@9iH�Z\=,Z�����L!>�vtt�ui��X�J�8�+*r�@-E�ŝ$'�%�#0m1��"����Du9*�-:�]�:?�}65�ˋ�y�{ۨn|�B
����c���M���3
,��F���Ad���6yGj�R�g��.���S/a��髣=I(A-ǅ���+�۠��2KձtuW�9�{ 0��}G��n"J�uIo�������R�z$�<+\D0�v(����r��S��j	��<�9�2�eJ����N�XlxVHYEB     400     180���o~�W]��?�fM=��'���H�/����J��z�~�4���y�DT�D)K���w�q�Z!�����3��؊�נj�2u�"�k�u��˞�ۓQ��p�K}�y��]کG�E�9�W�p���	Z�K��.��w/`rm!-�5H�E+}�*��?���]1!�u����[Sr=�#;�X�Ww��B�m��	�;��X���z�DJ�!��x��1pʦu�{� ss����ӱ�Br�E\Oޗ�
��R�������A�J�W�f<��Z/Ӂ6P�d��S�yD����E�q�o���}����_�3���v� ��6�/����B�P88�e�y�����#���J|�/�K�����a���ż1{}�,�XlxVHYEB     400     150r=���b���n���䃛��"w��G����Hsz&��b9YU��L����!���O�3�h������U�^hx���g����*O�Aْ��~L�:jE/�&��X��M��S?/3����Á�����)��6F�i��� �EQ
^�]��Y���J� ��lيLE�?6&ܘ��h�\�3LVwjު�U}�I�w;-������F�/W8���:T	���s�^~G��hkAQH4�N��b�-�t�>���k)D�"W�z��G��d<��Y�9PM����6
����5�l�![D|��o��G��=�q�&��7��to�6q��F��{�_>XlxVHYEB     400     120q��k`Λ0�&�T�۱�"����@�]s�C�H�Xj�Ձ�C��� ,Y$y�Tށ�k�o���7.�k���E���O}��������lmhQC�塖��X/Rfʴ"��R�#P���&�<�ɨ��~E��o�qT�I�x�����D��ʢ*DoS�ٟ���������)c�j3�u~�_��j
��m�=m��p�d�D���5�=�����
[�ܦ�a�/�C���ybW3��b���7�}'�q�ƨպ)�[��M�@T��!	������2sc��F�XlxVHYEB     400     100@,Z��(t=�q�:*_d(���U&8B�,�-VSw!-��i�}#��b�oq;8��$ϓ�����jP�>�0���wh�}���451ΡB�!F�D^D���^w��FC���\�rQ��m�чٜ|�W�L�J�e/���h}O����k+-�	eǮ���%s�}I���qs%uc���%��ƹ��]�Ӻ���FP)�L`T�x�<���㜔��v�����i0�l�`���{���u�fC����XlxVHYEB     400     1a0�X��;�1�W{®�sͺ�.(�M���2��"���Ie���Uk��+�g�|�w�D��zbտd�5���x4����
���g߹�@�B=�Q4L���h��a�;��ܼ�N�w(��F�U�A��p�,n��!(���1�~0���)S-����q\pb.oR�G��Ur@��~����H��4%���%�Y��+�LM�m�	z�x�&�*�h'��&Ը}_OCr����P��g�I��gٗ�m}�ď?,ۍ�x���(m�#p1G�������؛ض��R��[��p'%IGV�bC�A�����ds�?	�2'�9��������J�ݜ���4�7�� �zir>�B0l����z�&��!����QiB�F��6�]�|}�߸՝�XJ,��,�s�,� q.XlxVHYEB      27      30).�[U3ΖcR���;�{l䞲���"b: `K��u���F