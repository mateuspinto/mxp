`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11824)
`protect data_block
6ZNkSEgpxdq4blrdOIM4+oZDtyCxiO+/2qytLWxGgyNchr1SyYRB06j5NRkxVl6AAuZkNNCWhKPM
ywO+eImMrdrS8l2JyC0obKK6rV6BwlaG2TSWpalfStnb0R9ltfodoa0K6Jk8Xe09U8rFtRnU+CIy
d8ymDrv/62BRXX3BQCSN30kG6mvNZql8DycpvRk6ubAMPKtbvZnF1Uq67fa4gCsIv2uWEiGF7+OQ
iZXigtLnGaHJJq+3Q/9HmR24D5QEhkC1udehC3TlBoIPOZuqX/e2A1BesP+ih2H0r710CIx3LVqu
z5VNzpSL96l0dJUrvk9GmJsTa1ow3qA/JgDLAZCfpVV/O8goL1cAJ4/6dK3JfDsTkMDOVKDbM1oZ
VM/SdnN7PsyzAh+AgmafFqe08t3Kx44/EJq7ewn6/RI2N618oTlOckt5K06bCo7ONBJt5w0Xx1Qx
l+Rlgd9fuS0SAeFoTYxv3ALGPn4mzIJ8sgx8RZ5vt9rGJl/yVGj9M+tkNndMrCh4BbymRj6ExLV3
c+6n1I9XLxcGngymLvS0p5Pq4Tm2EgiKiHuYjRURBnbl3CfskkhGWu18zWA552FccUN/d9jOwFZZ
KMx/iNgHAM0CGtqxna2cVJmkyBSUYa3WxetYxk95kVevJJYOaxsLcxJoX0oZro8BCY4GbWhhLWZY
zfcHu7TSe9WGxxDZfZxvYuF4UuGfK2GHEqUUJombFp0/mwvnS7p3hczXBhXtLtKZFH58kfCfDJok
DOffN72AUjPdsNXZfNDKaFmIsMsEEbG2UtNOzWnArycCmDFypKx9yniNAhQly5fst/q3sg/j6o/V
D9LDmo9B0Z5kE41KCOnIft9vJyn657KTi50DVDgII0WUUYQFYv9pCixJZGlb9RHGW4sB7+2I2qwk
9Vc/UIUX1RK9CFI6MPTWdVrhM/0a1fXs9qimH2+4s+hxPRV8fl/q3tQ2Z2eQQcEg2MeIOHoU/p/v
6fTXezMT6YFTo2OI33wcTrgGugFyOgXfYdQ+aTykqT+F2b+ChixTfqZ08IS1Z+6bMBd95A55k/m1
NOF4k5dQgbcoEDXB0Dj2h5j/9WvyokwqSVdaBqT+/M6auGxlmP8ZiacIIutW3p1hzD5ROb2HHg+Z
97gaV1QSeKB7o/bAqSkT9ujeOYTY+eMzEbho/DIwDKnpb9fST+vceTDXYbZYoboG+LX4zGqqM3s4
8mpqOLhsa82D+ObtsaDXc9b6gKgt94qpzRMaMSNCwTeuYO4q5jtiCCHd8TgqQmFC0jQyJHUqBMqT
eL8yP3P7qsJ+lHsR9hEvz9BGgYgzKaNv9OH0PEd4sMxNsMZhfZoEEHTu1fsoDhp9iBC/r3GQrTs+
h+Yis2A2EvtgoZDVjB5iAvLNvvmI77wYvIpwa+psj1fegI34d+0DkjkestWNLXKeaheMNqynuAf7
QdPA/B8yW/HK4w2Qq0EDzPvTTe8Ic9LGCrenkCZWbcdNJyf95Peoxwn4P8QdT+VBe7/TovrWUuGM
M/HmWHZGCwmbn/IkrreCjA0vrvardcyXc6gwXgzwwNjvian77i8xAWvQ6O4dgmbc2fYGw3qdQ/fN
98bvI2iEk0wUQ7dO2eLUZHegdGg3dd+YuyCZ5G4NZ+eBHrd7N1YXPzecByEAZFs0fxNSCYSQsb1y
uQ3hmLQaC3YAx+jBC2fx+AEEaEaBo24GsIbQg/qoqTCiZ42AYapqTWVtOVtYlW5DTXmm0LsEXh6n
ysHWEfcZjK8uY4M7rr+qFwa7ub3WRGuKlOA2+NJgcXT4iQ6NOn4KLUZiw6hGzc9a0G3zjPrGtgC8
5JWrwfz3PJiPi4YQauMfOwPjNyfztbPC5J31qnINlbcQgM3FV4GV7gr5dR8nIg9Ptu5dECU/yLii
omoPeswRryBQfvmo0jTbg0QIoAgQbqScVTQy1Bij7PSGKqvnORkEqu+BjWCUtdUHkRWj87sY8QgT
0LQ7uIqjKXovzcDVGB5zihsrg5XS0Pa744/so8MKhm2UADqVPuVgbniQrMimcNKpGtisKqSs6t8h
wiGNN9tzZEQqX0b8MKh5dp4sD6elDtfg07GbI0PGEJpcrvKbaKDd5u3b2t59GZaxEood4/h+qJtv
yMeWcfGrWlsA3LojnIBaRlfVCphv3giYTFv1GKijnpxsgSz/LvcXM6M6CoFZfIB2uQkMrqGmqzfx
MJIaLYuyQ26v/aC+oZGtZvuu3S50G2vDdRJUErkDMUJQxVLSQunLT+iOkdl6aJM1FOvinIY5Wl6f
pb5xlR790FEKPYG2ELAjM6ADurxV3Bpbp+86i2NKlaEgqbQMzSlDABZaMM/IztVjG1BXfGU76wFl
lyMxuBWM/4gI8MgRfZitQIX5G1cw7GO66D+zev9wY147k2+u2+ju/7hVH3D8W28csR6K7DP9MJCk
H5VDJyPY/tcWyK4Y/t9ijKcztYw8acZosldBTxzL8CzGhzsEe4JS/03Gc2zNMjypPpLip5NiuFNz
2v5OKo5jt7FqvVYBwIQHlukIbUaDB6mtdVJWjdBgYhO5Hj5dMwAa+20UYyk+UGfqxpC9sDm/lWoJ
19kcvtAIiahVMAyqT6Do0dIDs5T+kwhQQbYHX1+e/KrX9U1dTqe1LZlcQHpoHco7fHOGagd1BZY6
qvh1owy3i0ClKbo96jrbEcL9yFew6PKhMhumHE1LZzoUi8az1zy0KPQFeyiGj4ukFf/53YnXvcjN
AX9bUcbyySqCjyR3TbuLOrtNuCaok88lpjfVqxDQ65Bpyz4tAxOqz0tv+thZI7bc5WdcNSyVnmBB
9c7smKn+qEnaq3+t7+LJ/QwXjF7g6H8RHH+X1eRalvF6cpmOpebAc1gqlqZn0kU+5tnqdApHcM4E
AbiU4+uEm6VaofRcysbHA5415w/UNdn4F0PsnoKlpmFM4qq0uj5upGeLhcLCiSPh9fhiJh2Xo71L
3Oc2cXKZ05Ybmh4mu9zy0vhDk/cHTdj9wEodTiW4853v2Ht0hhGjMiL8d5hbvkkxQxfSQPB4+4Rc
neLWxDnmggYbUcB88RUG346rB7HeR+A9arhaBb3Bervfotul/On2ey0dxltCsraMvLeeAObMM29k
IZz6X9J5G40ISklz+qjeHh2JFI1Qv5Rx4JYXIA7DXbShaXontzjfAHMTCF1h1r2fUJvhEFPwsHrz
JBtZ/KW7PoPsqibUYrrfIf948y2n1mlwTFsGdEd2aAiSzfs8zSSL5/dF1CwFZwA0gI0q0SB5niYG
43Ei7Iu2ThYVJLjI8FyM/Gyf7dVAlQY7EuR8s4VJxXfx5qutu3xR7n2x3VaL1bHYzTIi7Y9cf/+n
6oOBYKANNTVpPMLj8tDZTAfJYEI3r2rql+uC3zf2zuKCxF2DFft+dtlTk7FtIAM/ZCMbQTQUtH5h
xNh+VZtALCejx7kGuSnXPOBFRR1Y/QJEfNt8VIrt5NjLdv38MoXaNZ4QN+kOnYBhW3wrh8/TSLss
FzBbr6R7hUikW/ly88E83rcZyG8ComiiCwBmBzXi+3SLo/xlWB9QstOCOe2DWGlq8LhG6vr3np/M
E55VN/Q05Z+81gVv8Vm6ju2Ehy5OOUhR/uz7TgnTqDINMXsZmnvg1PuS/kjc9EG57hz5lbOcsWAA
7Ipf1qNqfrQpoOPcVgENtMxs+2RJtApbut7ugZnrOUkMj/opntjdHeX9a+k5pCcjyItFx5sJOwk9
QtHF6jxIf31cjEQkAsALCd1jEFtN1jmr9QHYYM9yhk0csF45myJL4iFQmI5daTJupof8Fa+hCjJJ
0WLmA8Rs79JPOUIjS//i9/iweoOWK/sypJOi9XoOLwFsifOIBmEZr84hlNvDVNSteTW2v80yQtqg
sEWctmmopTwJY+5pJ68DADx5VknP4PKB/EySuQraAjqFp2ufBMIWVPmGl7+/ubdpKIl5MqQrKwmZ
eWm357BXlWBhboAAZ5kSZH1CMR0rm8h3bvaisb+DZMw4DOi/Kd0adKsHg9p0ohoiRXwMbkLETdbH
cenA/QWx4x2ehc74C2y2gIt0TWfpNS3pDAPl1SpHtPTgsyj+YxIoDgp2c8QErc01F1/C4S6jP5ob
Bg/zO8JCV4ADp/PPhn2lmieaEeJWm8niZDDcG1+NoRdp02GZPT11rBF2TUNkXdyHCuRRIxjBrLoX
MsxWHmOIGe3MW9/ldh5bK8pIqcRhULUs/oPipdgHLiIxVo62NVk83QV9bP2yi7ry0ywfHSPdmW3I
eT7rwwdB64m7nCuqardNBxdi0lswvQCNc/PJjT2nYnxFinBKRIcuWYUq5eibjhhZY8TGfi4Xm0YA
A2Km408y/yV1w/Z4BpDxSd69CydOzLpYsoodD2PkvpAgJxVRXTJEOX28R/AtGmsLsJzAi2vqm8et
Emgekmogrb+/pqWtenFShgo0kcSHItOPbQVTd7yYZ/Hl81PyaZL5jxbDpgFjM9KO47jymjXWJLmV
gzWhBCxh/00Fa8zT8YwfQcM5B3onneOfwZ2fdAaJdcqSjUzQJbV/zKohxcuDgt66WJzL+M4ibYwG
68E3Xzci3JaKBXqjDfG3DsWm8vR6atn+UCTcKv9oOvKgMGj4iNCbYC2JycREM+7kDB2YXE3E9Nwy
UemUYcmscd5QmC9DSv05jtcg3H4qdkSjDyScsmSlDOvGc3g7nNNt0xkxfTC8QFFNaIJJyBkQxn1Q
3o2iENEW38eZi4doC6CwpD0H+jGGcnbnrzzK6sj3D7pe3yRaVyy2rmzQVTcCGbuvvt2UAqIXQHG9
Vp/SSnrwP3DtWT1pKvHwgdV+RmUdgtY5qk4+eaChr6XnajcxW85Gc4n4GE7+r8N2Oh3NaBjhaWc+
/pTNg8TdxhJ3BZgTbEzfOLcwWOGWj6oZfDcXiUqMs+RISVxYlo8Ow5ONtzKhm3HK1jEwgEuAHozD
X42gbD6+hAXNtDuSslFwAi/HkKo3qUmyi7y3kbzR/FzjKGODENxfFaSWstwRCqlpJ8Q8cjjbVxuV
WIXKnCP8s+luXQR4jDeXKwnH0K3nDoVu7dON7ARE1FjqOXoujlmK4R2Op7h28P8b3fdt3qsMBqyr
MSNDtPnUNZ1y5E/MXlgKnQEPuUmDYbpl9u8GfHrRyoP+wXbF7mxV+U8l5W1mXnY+c1LGGhfhl6/J
WTcUHHmqYH3EFQ0N20NgzMkA8/zW1nJ7KndRkTpxCa9uVnLyFrJIgj+WPlrdq/cxT+fb1u3OiF5M
vno7ozU5Uts64kyF1aUmDc1EFk7/ZSz96nflG/oJj3YJLy9DOllM3kKqf2Lq9RwQKJ/cyZ7ifw3d
w7QSe86YLxnWGZGSlnjrUBfaHlOjFgbD1fQ3652HaAItQzzYV5iVhuTB/hQygc1O4/1+s0wZvB5+
RObE/S75XuAARglDF45qWE1tTWoGA1OI/8kdZHW5lTdPbhnHbtxAk6IOI5pjsKKEgrDfakXEKaEO
oiXvVELcMX466GZS+KyovlC0WssQOEebtCeULmmuVnlUkye0X2FxAm9kr1aQbK0Cj+NguQHXNM6v
7mLCAe2kjXh9/yuVqa1OhWDcegjW/W4OEhB67Ml+LdA74NKbCwcZups4RraCCfI8XA/gOuZLXhHC
lIVp1RO9lroCX3IEw2rIoevRcNuzIKKdnBxkvR9p3KIGD5JuymdpfgWtQK3JC3Gd+LxislSPzaTb
KzuYGPCSaOTUxo7z2lp9mz93Vh5x8VOToSt5BqFs+0OmL3X9yMIIbTS8aUu2rlmKZWxkpbn9RmKr
SIC3OV7chPYc+jNapdH+kKdNBDvMYuQ5p6Uau+AGoM4RTPmyRd2ZfFB98BSbXUMFaAcOV2qwHpEk
rKU/scdHCUWDt5qD55GxTSkjIC4yEhPiZab5wlXwPN430t1OQgQ+7103+DRKugTtvedr8itjcyhr
mpFluQACEKr9XHVZEMGVwDBv696QcCpiR4I/1DYQA7pfLXqAH8jqqZOqeTLom1SPYljLdzY6H1RY
eD0aQo7PRhC4WrtVxxOaN6MByImDOTl1OG+KOUpqbHQFCfGSG22Wn/3fJVzgWY0D7EtH9soX8Ny+
FARUgHHIwDRAxiIzxnUPa9WnxTwvUESX/X/d3Nctjq0a+gjJHbedMHTQR3v2OQf9qO358+P16khD
shqvnCkpU1M+TUza+QtR+Yf7IDQbU8YRcuJcZzmRF2RdR+phil4PYipmEyMYgvZvPRP3YUgCzYx7
D0iVcR1V5qLswPYUy+Z+s0iV2HYk+zKynqQIegy1zq2WlctGubp18o+wGh1X0StuodQfc7GivELB
G59kgdRNs/QGRkYNQbFHiAYlFpXwwAse6S96LAES0qEpCZ9Rnq0hx/BZfhskW2+AcX0c2dOnC5Hk
1OPXWukkXkMVMJf+KHRmOwpg7K4zXo+NaBU7BB0IOtZeiCOkEi+q41jd3IgbE/rsfsqaw4cTWcr5
nzzpSM9pE95k6I8keANW1kmvcYdQ54pXfhWsb9jpeEv9TFdD6PFTcW9OWK5qPgM9be9jo9gFuDkb
fVOy8MH445jt6gRimRS9V0y9zrEcOVnYjSv/ETNISMpHXbXL8UcMVW+vrcfPJk2luhKiHtNvj/+a
ZEM5Mf0imyV9PfFgxa/h3/FAR4OGvGkNbJ+xiSYNSM8Eyw6BPFlrjNswoGJytojnjaDi8oygr4BM
OEbLMfYDZn26xUQ79+IKD/TGWICQ+zA31h3EwvBrGI/ZmfwJygBbxPCBVCqv9d4tsg0/d7STHX//
Nfz5S7i3Vg0Awz1+mZXJq0P0+4Be1OLVkna9Z3eyckzG7X02JGlb1HywdGYix0TnRQebJL7Un8BR
7CknVvfzV8DTmHUUyAwphn2QDXaCHeiTfbCFR59lSgvZZFsbxldllFQFAWSWq+HiB7aRsE3x3Awv
gUQtjeq23PtGK97OEI5sg/Fx6m6k1xIgpclx4Qp2ZbwFSCE03RXaIHALYtpbQE7+/BCQp7S0/Mwa
/4bOCIx+s5x1FhaVfx7tI5hoqBp3Zq7tuH2+WxIbgwgEzgE2v+IZPJflTWbnUfaZkkMQlVLDJRTb
Z7lMXeNv2T2O6nJwYUAGYpWyVhCH7EL0L+I/1WlZsHI0pywB1j7Nzs2RBj8/v4AgcvcxU2YIacqY
/XYAU0JX7OzCvthP4dmulWKYfh5Lzc6qY+n+JknUw6WX95RKPpEBW/KyN/Gz/kCkrbH/5k0s26VM
nM5l0wlAnBSmGWUSnUigpH9xDvONKsc7MxCE7ywwWgyQyTgf/D3vGi1kra6OB2LYoJfPYOKIdwoX
pmtcx1u87Qp2D5jYRwBFvE0j9Y2OlheT5NCd3PDSWtWtDJIa0AHK2iHa7KltCVTtD+kExI3b8D/s
Co8UcwWb7m0y/4SGmcLg5LNDpPT9wjnK3SwBgt1ppurX10zpaum9aldrG9uz7AFAvpsGmTHNP9VK
I4nvvWJj0ao4Ho4CA5gmINbi8OU2XpJrxd9mfIfFYmUoLJLXJm+HmxO4qY+OdWmLRDhpP/7lJwUg
ik3SkoLRPXkK2WKDaXZ/23YXCl7QLMML5aocfy/natyWnJchDb/A5itvTv4YQASsyIk99Ukqllqh
2TfVdFJvWoAh1FfWHdWmA5rUBKl3dqBqMd9pzzyG0GbFCcg8DxEUpYIOOgucRVz7wX0JNW6UtkpW
9X4c4ieuH4D7vl1pL2sOdIvr7wwCDohVDOKEuvtY40psZWVUo4qLkN+J/dXniw5JDHR5llHeG6Dh
Yeol3RzUvahEDgDyK1TzqfISRWFQR0ip5c8iQ1kqNYwqsNM/4AHusCQUK4Mdqx6ensUFyRCsuHSD
GUAFmSCd/iF7z1MEe+eiWsWs9yxqxKB8BS3a/np3TPug0/MPslLTX+3DIDV11QArkbr2fT2lER/g
A+YTtAoGHi1fy60Z/YBWXDxy0lc2nPau6qphEfoZrDgUGrA8HVAIOa5JsYkYH5kzk5MCAAPEYMaw
tQ9J5Kpxha+HsIO36MPHPhO6ygoRD2yRZQAiCGl7qNLpk/YnjhJ0yfNqQ3RaB7j7avlDmQR5pQQx
InYwtKA17cw0d/bZbApvILmKtc5M1v+JJblKXHsnx0jhJFdQmr6x6JBxAvjiUaQybODF6EOEdwIl
4e2484QGVPFJtlOg018KI1VzwQ8b9pm6PfrvlN/gCpgAZ/7wSrQaT5KJ7Q21OQVo/0jB0hCtZjQo
NDTFYs+223PaiO1req/5pw/i+9SRT23ETJGh5qdU0UAfwGB58VayOQZq2tlkMv0xLWqQYhTIY3zs
MM5vMgFO0ilcJwTcr5llZXLQ9vOb51ZZI3IwKh1wnYhIdcrXpAOQeec3kjBsFpP/yHnPYNJntvNQ
LXi+oJObOLX3Ejgt8dfOUF5c45ThsvfPfHICISg9wIbhcoEpB3PLzPwaRN7qw0kdLq7eDubXJdkL
Vi1aUFIwvwZge5QLV498Q6Ambz2vyHiUDlijHBeL5tRKFy11ldps3PGWITp1oDn+GIT6RluPoEQb
JMlv7UQz2bPrGG3gWoUnSqJrix4PMWBrNlsUPHenSTetjOR1Wf5g8SBynpVpDopwFKTNiqw/SHD2
/fp8fHEdgqT6Z+MBszv7GlGyDBwL42W3sAM92Tqw+mVk7g7SoDfogO1rwTwDVfgWWHFKAWThtEt/
5LpvEdWOlGbyEhdeJwumE6YiRN4gNS5c8j2cVXhqPGgx417I57mVt4dWrcWl0cW5j/TTj//LCrqX
eLEMlHIk9VARYW98IW4w7Yuse1wVDexi2B9OkZt1Y1GsVg/j72oQ8cuuO+Rb8Ou/tEaunbegJNGs
qtIimTa2cMO+QFQ5sDnP4AG19gc+sLjcR3Y9gTo6Hs2jK6E20sOiBTbAfz1S4jN+FbnO0t+j0BJn
Vej2y4RZMA4yAeevAELbGYlyA+xarhd4BYQF60LfIVp5UiOJS0R7omGLYiPtXHD0MHY1KyfH3Dp6
2afOuDLZFFJ/R+l0hGoX6UAwvNu6josC/3nYtpZhxIPve2o5/Ypgh1bepCBb5FZC9cZU7MLzqzqs
8/OvHjAdqd9HoStIZRGPIQlC+8UOQOy8cm3zgI5WWO1AFxSVC4NbRefXuSINNrPD2oGPDykG6DA2
hWPO1qFJLP4+CfJEHMK8xQmRR3KNE1F62HaeJBAgK/d3ffE21xGOdAC3uYv2YXwBqk4KAnXYAp93
fh93TZoSbmAYqHsSAlT9dO8yGnbBzWdBCV33yk3+LYhERDh0+8nIKRvHMISAPMiptbglAa44aZli
KnkFXIH0TOwBF4xbNLDzsw9YhhJxkp0TnV5mu8zLH2qCuE0i2ptSAjgbM1jdRQyy5XgUQNNS8qb6
OnXCKSghouhRGUJ/k36sC7zA2O815FLlFX3hqyiw2U2i8ZpfEXxm2LsXIe/YAeO/aeczWLUSm5wo
x23TDrku1hobSKI/vw9nPj5ufIqVq7P404ggVTmpF0nL4UcgKWGmMoqrwcytrVHShtcAcS/YjaXS
1TwUDdeACZLZj9oUhAB1aPBMEVd68g/Ygp1nkw1SeAvdUB979uIst+GFPY3vxSqZJ3ec1QlBaF+9
BuY2SRB271B4r3P8WcKR5WUESj6HIg5sFHhFSuRYHquhKK9RXF0eX9Vlou9Pg3Npz5I/nlAYDzLW
usqKa6/33kcjswUu5/gi9nFVZL2XnAPflfUPBwPuLz9kNCMU504XnHe+8dDEI+r0AANLQ7b7FOSH
UY4wZwnpCxy9C9ukdVWwbGZhRKI65fdjdy7hI55aJd0Oj8c7x0b/NWzGMQ2gKk9rSUV8yB/u2r68
oRAcBIj8iKiXoB7ksJ5ESYGNwvzlRIZFKArUxC0hJRub5kFChgt4sh3bNYobvl9hjoVxXOFrbEJv
C+W8IidO4J7LeOvKGsQAZFLg0zH208/plHRbXtOC/nWulaMMFPPjzLdKSaoBE0d8R4LuA+av2siW
8oTpXTqxMPmJDvC4VO4ovUjAZbEFwL7f+9gX8e4S0v+t+ULTouT02jZv1TzLmaWuiy/oD5WOAA4x
9j0BUN5HoL9A26dTs+VXE13V2sL2z+v+zjTM2pRV9EIQ37vjxzZAO8/716Yyf/+I2Uvtcjy43sRF
mQbq8ZxuNobPJ56CNyPwDlpAVe8Qg/ZueBKJPvopRg//MTjY2u01ozEGaeETUy8A7K7nLvqM/RYv
ao102C1VxaeARyhERoSrSGbUVHRNh8dBk99SkggHGnG8JrD7mLehf+A5UPzFsx0m02jQwsp7Qn7w
e6mmyRocqR1PFBu2sSEP942h2ccr10SEzOsYEmwHSeOJS1Cp+YKbqtBx6ZRREYa/nL6TFlL5tmER
qR/IzEIO+WGNFdPxthZ/yNGxH5PsSIpHJ+6YDi3Rh1lEMKu9r9EH/GOmw2K7WMKnYlhlDksAbBlX
kJHXB0qWu8svpSW5GwMCLg1wT3cyBIHPpVraWaBKhVPSdbl/BguVKCLrL4o5Vq4jtLJfN0cOsGll
Ih9K8mMA2iTJqXrN45oEh+9iVOCpkBVNXCM1Uf5Jh5mPd1QQNWQl2jwI3wIqM/22S/abV5XQX2fI
WFsm3Q5dmbUDrnBBvRN9u12CyR/+SMqF07AXbwdmL2ReAP3BnFWFPzDT5u/wiV7+kr5BnD1ZFj06
VIXaCCao2Sj7D0uF7Z6saW2DVl3AI/YZmFKNiVC4Xng2lJhXlQURw+r7TyeKySDQZlJbT6gFGa8A
8PhWZmd32mrAOsUKZP0LxVAg579Xynl4hYSxalq+xJQI2/Ue3bwj4IBpuArE/sclYQhMJZs5/TJD
tsvdVRjuTLms2iegrIBjMeze5S23bYx2+H08Ohg1ynJFkxQI/1iW+Y+ILuvAfKcZWIIckbUQaHx8
2djR6ArqU+fSv1aCLMG1mLVOuhz40yMHgbW5c2amxpO7NwMYsCtGSNAckRNBx9JgRMdjilw96u3M
lddboF1VMqhzoO7VbGkq7fqFbz+V5N5OnGMJDFl9xntyQfK9fxDzbFiFPv8pduLQI2emaV+OXROr
xGCxK6xpZpR4dQ+IrY/++5BkPWvcXIfIRzFVP+66d+O7c3Io57BdkeV51pwVIAY+MrYRJlzD2N9Z
/KO8EbYeNfq+JAe2EeQUPII7ChOBVIIAqcAGin2OhHYvjs0PxaBw/EEpkF5hLXrNlqrUSCdlg/hc
XMLQKlMUEC18H4vpvqtorZOyJnAflLjWBwATUymbBd1v9bcauTDnkDfoYKonfYsW2Z3ar7RjW3Y4
ETznmWtiyTHqgRn0FcVKWP75Uss3hJZROk/ifooB/YcZyaQv91xiexfH/FLEaHTdN+s+wZGIXJQV
bBq0CB5nohR25DP7bCxhEAQvvLPQcBzAjz/W2pAn26UEhA2FaTuGFub2juHlp7TLz7DdqKkAzjLh
MmGdqYJOcuD7tCT8VfzQTu1JfNWvxpMuE2Bz3Qe3bZpuFwhLSw+4eG4Z5t+MhaxaiQaHSbbIPEyr
VScBNoybaanzzEbCayBqOUVf5sI52tziIMQafOTkZbxRk2nCjRy3JKlbVxbVabINTca1JXZlgt18
6ePP82miBLOlXIuxebRusmW+hwMCsGERBL5m4LfZDOTaSu97/YROsSLosSaghIg35Ls06VU+X22P
h21Q71t5mFggTaqkZP3JhNH3pOx9hab7CKXGTgH00r5qUG011gActYQ1+CNl9TFPnFvu1O5+biIG
x1IibyrskPf28aIgK9EXbdchIShKC7giOyMT38RiGEz1lpi6T63k+G6iqx/3fHRDbl1W0OucZaTz
sm16TrIr5vBHkOSvFiHg6j1YYz1idFlwT+rQOuxQvgDmSg+7sfVajAOtb8v1jG4At0nrGtt562do
dMnbF6jc13+hO2Ai7sil/NFktO2uXDFTwB2mB1vPINRpypVgBLu1BqQadnryZ4ckkMSIco2Bd3h5
RNyCwDFfbqHD6ssAH+z27CZ/SzAZPU4QYNzvlo4qBhr64kzd10dBEHYYIfLOgYHxGAk0Ujp6vV/K
+8EsoUN+XfpUvEtT5sK2WtHI9eyDQi7tNgbD3i2+i4pgNnAovlK+DBa5+ZQjl+wJ557KbYLnrjz9
s019q2OXlyUF2qQ97kfvHERka2aN1GIOb/r6Faz6ZZOAPjppA9eM0GaZOkinLHl7OyNozIv1JfEH
2Z9WapMJttjnqtTnLYddqMtEE/+Xp7cVkMnzNnTJLIQsrU6SEE1TrmvPk6Vqaaok0qi23VMfCva6
jX7GRkM8ocZ+91DpGKu7TxaCj4PcsSuyUlyTEb96j8RvpZtzBj8lRm+GaO7P20tnWbTuhKl7Dc3e
BuJkJ2TQcBfNfNdNWVQawvp0V8iRsMSwMG/2cMzBpnov6yss6Gx4fTFSF0uhTF/dkagFFdeDE0+3
DCmfZOUK7E9aaJwHfmdecYJEiR7DHtwX1PJlu+R9+6Hd5f35zCk90P/q6Qj3xEgJ9Ggs/+I0FoW9
RyyK8uAUoSmM5MpE015g9jRJY5GztAMwiOAQhHK3QXgpv2eWHFpOJh+5JYsSRXuMCSL6VitOxCvW
byQHO3Jw2xv6YrcZwPOaI/sDRzgkpggmsnyo3Rj9Lf7eHwewyPmEvaENMZgkddBMcQGQwp7HWmUa
AstmiU2xWy6A6J1CRRiL6TZDX9WCDvIakUuclS4+/m0yVbfrA9JIHi3gk9dMDbTmh3sY1WzazkZk
dA6CbO1mca69X6yyvGawtjG43gaS2WwN1p6pxnhWKQtEMSsKzEOLgQIscDuDFsL56nsrK6VxYfoH
fzp6VZ7BEuYmqBV0RotbvYknUbK2B8MhUzuE1jGW7JdKY7UFUYCDZ6gFqdZ5Vm8j5lnZh2rTnHvU
CoHDl4xySvnvg9kz7drAEQq5Cl2YgbQma+BxJh2LalKpeUBfVjC0TMCoIKBfs0+/mp9CC86RVILP
E+D/Spgcsw3GMgsQuiOaIL4rROClSfwaVO4zrfm2I/C5GUS3esM0W0MYB1gYO3Heaovm6906YRS0
YASqEei52COkw0JwPH7+hzDOHnXLz9KhXQkbyBfT3sVzhOSMvGON53XHGyMt5M2ehQJiOc11ERWM
ANiWve4WaMoeYEvWvReZheKIH9ckh+cwV2Lh76X2xhUlkEmTjh19caM8yC36cIrtPO4gUj5lWa3s
nr+NMOntu3uNsl5vyFmcdxZ0Cv5IYolPZSdgFlNwudqt70WA1lpsDLmbzeRCMAbgGg+WTwjznPnn
4zxZUtU7yxM9DLTDdxeZBhDg1le4/HZ91ESku0M2rH42EYVeCcYZ/z9Gl3W/P4AUQexOMRnoWv7O
knf12tbKtWzr66+RpCJFa4cObC1IwHfnRSoix1VEms9Ex4XC59rY0fFodACWUPkV85Tq3tVmVbvy
HCVmGkPNfJNC+TwbE0EEmKNZLAT0bij7yfM3o9uPWxLdbhTMK3mmrTKTukNcIjc3VGKSc/bE3CzB
BnBqBM9tUVWKffCiTG1aHbyI4dI38bwdUeN0TCvG/Avs2i1Bj6HFX2c/rq/CzX2JJsk/3lcSQVSE
TuIxIOOGS4eqilt6639TYlP6XDYwTUWhhH+F3N6tprwPr7wmJlNrQKOW/vIp4gRXV788aHpMufxZ
CMWnbdaBOHkWhQ9AyC7AlbXS0vdLLy4HIHsotMmsJQt3pHbDnBgFtzDBKdCIm9wNTOdlA46K/oW2
MQQx8PNe0tl7sudPNnr9t8wzyKHoPwLXM2QQcEcKKgxfrtUAZRRbB2UeyvmPTjb0fjNQyZos0/Y3
iDS+vlLjy0eQB/n9iFJwOda3vY7LuW7yvgReVeK2XwJo+4nR4stQTTeLvUf2noaLEDxYvrL15qNw
cveGbnPP2yehYr5pXAYaBXvE/4iG2M/j/g9ks7u6rcfxdvDpQmjtzmJZXNgTWmt6+KwOrAGYNTIY
BJU5BAeGsg94yI27H4XwIfLIABMVodwxAX/Q/w9+wb7kZMwCR5Nly+YdXG3besZjCMX+52MDTbxR
ErUfhappyxhfrJpcMWN4zS5WDq2ZFYe4JT4UBVXrcbHvFn41NrjJSQtrb1LVbigtygp0L0ptJ2ZQ
xlmZcCtsOHA2nDsCboW/mgTSmKSI2gjSaFpqtwjwvOdFmZ5u1og98zXQJ8o8PuuNo6iAbxCIRJvf
QhOIDsC/OB63Efuiwvuz0DK9p+yYerOz+O6OCrtGLHxe34KEzMijfLuqcf86PxVWNjmVfibJs2dU
RVGkJH2XYmE0N5LHaFQzW528uCzG8wijcWuNSoVskyAeRz/1fY41aPp19K8FSfuNMv1uVGzQ/MyS
zOsoW7dGTACO70RakwwMQNWuYEvGCLKlV/num+bfyKdeIAWxkwMJtarhy6+UHF32yJe/dXUysV3l
qxokAa8ubFne7uZRjpoXvRZZI3OP7kRZhcdMYCwWPEg21fCrsUGxkP5jVtk38qmrEumg/6T/imb0
tGANZcERJF8WjKJOLPSz6e9rl7uwCsFiz1ZoMVyhDEqQrk7rmfUanYGoQJ2t/N/cH1Ri8cQ8qd0/
E6zsZciLTP6crV6shknvgwEX5zr5sDXeMw9YHjDbxSQoVB///tZ24LER4Le6WbK+7crjEQrdXI2/
HczTMCXt6h44niF2DB8568WtB57BrmkRk8AhKfz7wMvIU4Y9PzpMD/VOH65oEHhCQJcrmuHATb8I
4+mrOayEEGVGlGugxr0tRWyHDVHCdhqDw8cpHDIpop8brLy01PDP8AofoRdIg0u5qS/WcLmZn4aD
g2TqsMJi/hFNfscPoBDhvwIM3nfT0gFRk3DUqoYVw7oqLj5Z7Sy6IdWAJbOQsRapl/TQB/vyWnoT
yFdQ8Ff2Yha9mq6Am/e0pkOFSCSn26beKQjMoIx7XinIopKnsTw2OkVG3YftAuP5M3wyzGfm+yrN
bq5a40TNzpCuxf7GMU3eGO2cTsf4cua8PaYKgnIyO7rIJuNUraPhCLQ7G1nMnwkucAdakcfARkC6
k5ukNNiFoXQkJ6E2eS28x/t6ZpBrZcrn8uFaT+aw7Cvj7ABNSdkIrUkZmBvlBiydLTU4aPSnfJVR
RLmewuM1muIPLOi9mk/KNXXJ/MBtQzRFex5z7qwPPvcHXXB+xoG0iCsOgeThpKRyTI3SytS295Rh
nSfBFV20k69OsQ2yM04Oe1XUVZ1p4LD2jotCjpp0bn3e8FEfu1Er2rhE86XltN0ATjUeImaBpqf4
ul48pUB/stRXsLCESmhvip60z3WZpoxB9a1WzVvdIWtuHYvdO5NJoyc7cU84GGUjz/ZaxHa5jdSQ
SdE4ZV616Y/eCoG/Pult1lu6HHgDHZc4d4V5Q9UrK0GqfGttrAJenzIdGMiHPZJIVIc0FWMBb6sb
HZEGVPsUq4w8vcCx5r0hG4FI42bO0DyfOlDjfrGA+6kAg1A1PXQaa/KrjaAKZgCzWV7mvEj9lzwE
ONqM3vqMcBbelWv/L8SpAAa688V6VQIDzVJ+3SVctBQUjM4WdEWvEFi+lYn2sZN14SpX3eV+M5De
XxSipo55Ekh1trdVw0J4AuwzyBW7JIJQ70X7nACMxdT52j8ew1s8E8emFiyzGDVu/f3UdLh/L+8k
cpBB/+uWfgII8drhcGuIqQw4X1LcZATjh1cC2MuF2xgClas80qBC9J+l24W2BzF2mAuOdQU5PEAQ
MsYUmUkON8WM9x1Ev0uAdUKbfO+Zm/vye4Aq/+GpGM10YchxtN/ZXQjgMwrraZT+CGFprX86/c6H
wFiMuM3awuDBeD091Ne5B7zurIIFEYnN4Q==
`protect end_protected
