`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
AkykdZkCOt1h5up0rqhhjuup4OkVCtLn/awd2MHkRff2XfTxozcnoz/9GWCUVjD7gN+YSwVX983F
rtz08heFIuoeqSd94agMYfrBJcRkRY+EvRfx/n2itSAkuGTu5OHbY1ZQ63XBoxoC7AiBUBqsWGWG
oB1x83GZ5+oyWCvNpKTyzJqqpn93+MRZ3oQJJ4rMGm3LftZTV+wr1yc0omJAR5erqLeId8RHCybs
vymtUFFR4GA6IpvjexYPcf332YJh4e4dml4maIuTYLrT2V5ie+8NyXSkmOqBTGvAMcv0hc4AHWZE
x1C6GgMTRG7VAU7vZZ/I9NKphLwmsMo1snZMeg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="ZQOBkSZMroN9VJUiDemvwHSq8MnUdPTPJ6P689y0R9c="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3520)
`protect data_block
h+wk3FsBYUHAKU8QDJDWzru9stw5y9z+oP3QscLTnW/4rlxSj2M01yLBWvSy1ZZLteUkAPLjOg3j
wg4uLUN6feGAUJFCfEJujaa/DA/Kd/7iPiyqeAQi1GmSE0SlL5ligzCy9bV0hsvandkmUPRi4NNW
ntFaoHrKh+iwtIkq8ATPK5TfC+T89K3t2xDgZpKs3mx2w49LwLzpOnqQufqmLcczlUsi+lORYUUG
conKw2xYqgIO1Lme0aPM17BFuYSbsuDdkXBk3Kh9gXroPSN0is3AUS0/3AqmQHoiMH1kVKc2Lnuk
g9rZ5Zwbniyd9bE/UQkLl8ta2f4TKbspBOe+jKU1YRvvGY6cNSZrioHPXAgzWmwnMtP+GPJr4Tve
x2PL/B4qf1JVFeOyz/QIHxEda10ujXNU+vsVJtyvAaMssvyoJXgrllm10xyIdMWbmD/7WAYEuEgK
B+V6DQvPcqdr9cysaShgoScaXS6dL7/f0jbHCA+DZ6/p3HXZnQv9Gpos3DMeqm5G4pW9eiNqV5Ae
DNAWG5p/eV3zhl+QfHQZXNx53Sl7OxbbGeMu6RZNXD0kyFiu63Pa1lANKE3SY5dnp21LZaALvwDQ
dTkxT05YqHldIcca8TCKSH4BwPpEipuqT8m2noWvQBqoi9I8B63eCnhCzoq2ss/MPqoWNfCTopzd
+rd2BB5N5Ib/vei1hAUiXkP3O/PdnmnRDCj6uf2wYnlCtpbLWTBBZLEK+G9iQnfRRlWxcPSqwlSk
TiS1Qo4zgT8md9tu0Aw+QXDXaXr0qBhI5SovGSTqWWTx/AN0HBqpnoXU5QT4Nk1HMwPmhx9swN2m
SHkWbYoZ/CLdRnvVe43MM3rqhF7GDsNyScrjtvzuO0GAiU6/lZ2uIASwt3FpQxXYvZEyholovpbw
8642T4oj85Y04BPtPsZDwrlo5DTMm6Sy2iflvWWe4Y0l/iUVD5fEKU1IFhSHjuIR1Vh4OWzZLF2Y
l4Ur+H71QuwAWNkn/P/3nQRlYYlLcRcps8tNf3twBJIcgNT2HhSda7GmsWONSa8sc6bgYp4D4CIf
Aofz1LTYHl69GSNhtAty5aOesXeD3o3maR8zhdxqg695qhabTp6/rXwuD7Ww1k9wFSaheBf0NnAx
ojjev+Ef8iPbw106nw1ZZ4EqXaqyccFamrCkcHY6h177XqUe2+oUJUO0F3j0/QifEMpNZNlOgDWN
jeXisGtxFWbtieVpjc0GqnnarsALrj0JvqkByWZ1jrpjh3MX/BGVfZmmsj5rlwGvJqADYS2F/heL
wKf6NTLE1LaDWZ7JiszoG33hhSAAlvVFIN4i90L7Mz6c6GNA5t+RSh9kDO9diB6vTYxWdCgb/fMi
UZFCwGL5VW5qjCo4O03o5crERsoVTa97VhclyccroLE7k3R3YlGnDVPRs6QFAY0U/zfQIwEh+83l
sfp8Qo7/orfZ9NNjrybe8sOxuaBIGsi9W7K6653MJk9QCf6E7lLuFeYseHWLoGlXX8LfakIwzVN9
rKBfcjaPppZLJFzNHKpIYHgCTp+P7J/Vp0zcoAAKfPwUu3EA4X/MTpnEgFYQ/IGtliWA+UPRl2Zm
9AmN4m1rufvpfkh4t1aTT+QjKt8xANMFGDiw6Ft42lkQkhGOiRYB/gYJ21jpW+T4FJvM73/zVdK0
E8noqeWrzI5NeDsgRVvCQ8ZBCh5Jm4cnaHvH//5KGoxuvmmjqjlm4AC4dHulz4+spe+HJfZVbuLI
te4DvoP0YYeOibF+MYCBwIGQYo2x+lBAFAUZI7YFyCw2QxoNce6/KR24Q8iJ/ufhWszy0y+3X7u5
of7tU0me0UeDMKBtNfOm8KRX3+5uqX9oR/7aCf1+phomI6qNEKorEZM88hjnpQJMYVsXAsP2jSkJ
/q18nZWBNrjUVnibVp09qC6gM4vv1e1vmLO0ABbu4ISQ3tgh1pbNHeQil0v7nlVFsaQScVpAYong
K9hcQhJgmk3bQCQS8supsE9FMXbYKE2glbhQPoNeztPD45bfT/uHXSi0dGjPaZWhMEdjdJSXhRdx
xWLRdylYwnR2UZ0huJp1T5ELG0TVXVl2i3V6Udv1zKz96wIMUJZGUoyys1rz4wQrzF7IWo/zPLMO
azlPw+rutJej+pG6/Yte/T7bwBwA/4WK3qUQ6TX37xD58j4hlw3y8g22gSilLBqpg/dtilO+a/Uv
rxPy2EtMd7hZTkPWarE6ZaI1iw2U7/9ROetKwaXP9QSdjwSAX/NZ/iT836wI3qLEFNSAQMeTTK+X
ikbzj4FVoGAr6+is1la5Z9AvvdcZGOgQ4gocZzQFUIIF4dY5ZsKAyvDluMWI8CTJBYZdoSPF5BgJ
xV5mYGgUC0Evs1v59ccATCVqk/fea6fpP3Vw61cblsx2CoYkjE4woS0AVrQM1o56Zt2k02DDVKC8
RXb/MEVGg5m11oIm8fdNwT3dNIgrjoorLWN8fMI0Tv1jBe+1WIxgPyQ+90zOb17jBknw6yRScAkB
nSSZm4qnB9iLHyNlgjz0wT3N0iVm9X0RI6KpRxbVCzC4IQD7Z/3SnQh9y+BR62pqvq0eIOl1tJGC
3QEmRkHnj+fCk78fsdeEM6BTPh0mqCNzvYoS7ntz/C0VpR97jDXH3lPl6kCjn6KGmzDRTxC6j2gf
GkSIXvVJKnVt6wmSwappUD7urS8S9MAR2AiyktLKIcdzYXrJIqZUNmd8jYcuYIWk9ZphJ5etjcdS
e9EyreuRjHl8r5A3NmT1i1AIsmHBKk63it4RQSvf4a3TkyUzzSLV57/plmoflN+7+pzBu0hYH9XV
lcE4y+Fw3kGFc5/N9+mhhvSXdX7zmFhSREIMICEvaCxJn+61N9W4Db8D4CL1+H2PoRzAGg10xDyk
jbR8AIIcG11vPIpWBNRV4j2pD5zo0RPuMPXD62J9oVB23rBRLKWx+JwAMmLCF0k2Fdcf+Ex9pT6A
jM/ZHuqzAzVjufsVUxZpMm7yDS8LHZGsVWRjt0xgLLgo8iRfFSmtF3kDInxLNEvC2kgj76q/nnwY
XOhlV4eBtKyegv62nHgdZFFGhnZwreVL79ha0mrsvH3SscesUjablh7EV4ZMH+KwRjAvCj2LOg2s
jaWROpVZ3JYxNmsxgmiam28/bN2c+uyURaO/E0fM5383M5WL4DJ+z6PNofulNOCqodR6V+BdEFRk
Iedbe6D161oVjLjbOSCoA/m6afBoAiiCz5kqiYQLIVzDvm46YahAOLgXRNPgnxWrFa4Pfq4rzcW6
uVQnhDbW+jw6HCUeuBwHRtG1GLLpmP/+TGSyzHrMm38Q8xCkdzRaNBvP8bLvySOqvL2M5e89cyky
hb6uhjNGFRulsZADHIPegEmhnLcsg/IcmhHOyFyMD9mOtgau8rcZCgM9KOsJIKmQ/uHllKDHdjcw
J5zAT4mgL58H3YNpp5vivkkioMq9YjBzwsAYEwWAl+6Ykpj7c62lyoeR0xY7RtM6/gF3FuZ5o6Ik
w1IbPSxVxlVfaHCJIX4aszOzu6jaGSr9CZ308ONVQAKobTXp8OCKu9HCYVg8oNXM5hidN1B5lu5d
s29HM5XUTkhNjCbSxS4/AW0dWhmnn7UENNLtGo4+4YaeObDBfKT+361fgKMdSMBN1+HW6bvBdf/B
67KAn8CQ+rWGrAiTsLoIiiWHbbGaobSwYF1PGjJmPiYW7VNXDPyLTRpD2Ur1YWoOw8R03q0bMi0Z
AuWiabKYyUf0f2Hyb3y5d+A86pZXsBqzlCLPF7AVfESYn3OjTGRopP9GyES2OxWDSJCIQSwLOLH1
hFsUqtTkboCmpUcHJctuTPy8/ih1lGmxyAxpsEDUzXqb11O8jCs6UainLp8QuqVqMMEG8SkVyeYb
2aBPML4YN9iujvI2NUZBnRbsWulS0nO6fnnph8dH2V9vvO4ZBX2HW1ob+OR4qHrP66wF0LvZO3TH
vesjn4aGlrDz8S87RyLN5i73SO0odUcBvXgF5ymBZ5vEb8TE7n+Un8GVV7wDINlWpkR+5E9Uwl/j
zDYxQFtPVmDK6evs8KRZ0FmwxO9LoDSUn7m531i4soh6fveicCnT1/YVUhUukmevehsDccxJhMiH
CxKuoLAwzUXMzZwjE6JRcls1LlO/CQsaZzlSJHHi70vWjlqjR/TRxEwC8HtU5qVDoYl/1rHyVJuS
a3Rh5ECqHKLlfERFl8d+i0dnxvxh6VK8S5PSTiD+IfJZWnAVM+pQr/RcjhmlCwFrRE5FEeKwMt6p
mehno8W2rmvxXh2iJ/iz8OUyXcc7AeceQzaFcj7BIAss7yKhDbZRWD9LB+L5gMoVyG7yfYp3dUrf
NLmZ5t3Rsq3bc4SW8dY6wqOoKeaENsp1Aj3zUA303EBoB45qSN5R4/UUnFrysLWl2SsBt29/+Iyw
QjF62Q5ZXERo8y88/rtYtCItXTfIPNZYU9qftp4x69CegA1hk7En8qgkXDt8VSOUyeWLmuxMRUTi
YasDF/8YVMRSPursN0wPxgeZr/GosgVaCLqGhTl+N/Iwarm3Qgm0LUGqc+P4/WZ9jnsF1PkxsYW+
8bow1rjTVwpWGndE2zEjN/KY1ByZDa8JHwOzThvb6Qdz3QFx0mb4AOdyIdQRWpMTv9AQC7t+ZiGu
8gbhuan9l6JYWn+5LtuD/5xZ1AGN24UAiYtjYjP28D4Ip59oGy88ncSesg==
`protect end_protected
