��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���kn*�PƐD�K��휊1���Pe�0�0C��Z�[QD��ۨe����W$�6$��SA�Y����A^��w,}O�`���/@TP��EK��?�s�$���N�����G�n�t�b��X�h�~��H��������:�z����n~�����/!��NwB��u�i����!5ĉI2���;N.%�k��V?>��aR3���1������1/~yx.�yAX]�����I�j؛����� �y���e�?B�a�¼�:��Y�V]΍�Xq����4�U�9	C4�*��q�Z������%y�aAF[�P<9�X/��u ��rJf�;8�VƔ�����!M��)��'�:@?���;$p�����s���v/ͅ@k.̷M722v��
*�GD��@�\������u[A0�b��>� �~�KR"D�y-�,)j��"o�4eQ��:Fٺ-`~1�Ii�XU$�IC�( ]vr�$N����D����
�i�e^��ML32�|��ھ�2�ݞ��pE,˄�J*����I�c��؟�᰺%�ӿvR:�k+��q�AY�����W�~P;i�ki^{\�W%dN2�M&
s��^m,�WB?�X�CMpn�� ɩH̴���V@��{^�ʀ�ʕ��F����W��iO��x�����cԀn���槈��u�8J	�M��4�4����C�����$���C��^~���~�2o�m�ы�5���$)&�3�8!g%��fa��`���#7Qdf:<rBW�q�懲$�|��}I�$;��*�!b�a#�cE9���J)���<� %����)��&B�3cn��=�wnC�e�>@Ƀ%_��p6�qm3�S:\샱4[@�
�SuU�>|�e�`��1�X��I ��uʭx��U0��U�\AI��M��s%���
����}��k�ݸ4��;[���}1�o����S4���k
@�C�� @X��< 85=�H��x���Uf�n$�Gl�r�����M�bט��;d��#IA�.��c1��l�0�
���g��0q��2^ht�lH/p��|��<z��k��xO��)�����(��>m�a��.����!�z�l{0�΍;�݁�ʺ�#
�y/��u_�F��'������Dz�Ɣ�ä%B�l�lK�`4�B"�m���N��a��i����,D��0v�v����*_.��u���'�+�i#����rx��lWUS�w���Hїb���P55L9�h��s/_�";�8,�Kj,ܻ5���dM��
�{=	������Fz^��uK�| �U,���F<qwoYTk�!�o͋��A(KT>�M,�YL�9���#���W�����M��9.�d�,_�#x��7�̾���H����v7��b�N8'���gI0R�Y�K��J�tח��]��4����O����Wآ�i7h�@s���!g~�l&��[㡬 2�!�o��qਂ��l:q����,Ɣ���/�,):��e��Iu����~0���42XYhg��C����}�?�?��S��rvaNn�r���d/���!�ؔ��H�[���z����m~ xCk�m�j9W��nVi!�������j�RE#Q�۬ך!��r�50r3��k3�)^��̞�
�&m�Ϫ��쥨Ϳz�dPBu����ϐ(�ʜH��g��_���ϰ��BDm��,�� �<*%OO�7�=�h]����`��3<�~����*J�X�A�a,��0i�E��6�-���Ѓ󷪘�mr*��X�Q��T��)����x�h$�
AEQ금��wm �E{2�7�@�cA7`	O"	����>�M�y��ߚN!*@���N����d�iq��Yf����G�v-�.E�y=m��;�̷��������U�d�������X+�q��G���r~����I��f�\��q>*du�`9O���3�_��\F��f�7�O}q�ؘ+s猫�p[`�z���!�