XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��S����v�(�kQ�ؓ��:�h�~�)٨.@]��1����J�൧:z��Yy!�?����Tǀh%�FZ~х���3_�Z� �j�U��yw��^^%}� B���S������ltf6��<Vr�4b�H+֯l�����|V]�Э���(^=��}��4�m�����s�N8]��	K�5����K	������1iC&���Tf�$��1�G�D,xR�Z�/j��+���}c��4a6P|N��a�� ~��Ł/ӡW���Մdg��|�O���˔Q(��Ӛg�fà��z�T�T��q��Pk��使6�	��1� ��!����h㙿zQ�p^Ⱦ�\�SI�(���J�F�3v��b.���>��)�����Vr$�����PQ'�v/�O�Ra��`�L9 �ɑX�����2#v�D����q4��4�k����#�3�43�]	�[MKgo;g{M�<2�5�p���f|�>+�N��j�gQNӵ�tC3�J�i#�*@��UR�tJll�n����ċ�y�j�m^�J[���3$�x�NjBɽ:B��E���l���j���m��nj@H�E�Ǵlob���g(x��6�tz-х#md�1�M+l �E�p��y��:,+���b�yF���U$Ѧ�\Y�袕�n�	�~��
լ�����mNt��w��O�L|�I�W380x��W�`9<�ƭB(n�Y�%2�d.�.d�,	L����VNa���{�:<��쉐�S	�'�;ְa#Y��!��XlxVHYEB     400     1a0���ԓ\ݘ6��Q�~LoIUB>�������z��hb��;0б�1���1J�%	��5y�J=g�>Ekr���B��((9	����}GkĈgB�U9G�c�^�#t%��F��8P�I����eaBo����v��Ϗd})iZF���"Ҝ-Q��#�l��*ز�$o
�˻�s���ÛTO������<sG���M5:�3ށ��J����+q�Ky^pI��Vjb��T�q���M`�&P!�q�?��9�[�tkc�0,��s�/'�;3��I������ߩ�A ���V�p�b����X�s{���| �����9�÷ky��eQ��>^`������ɢ�f-*��v	"�4��Q�X�)�
�x��n`��o�Ў����V]5�� N�XlxVHYEB     400     1b0����+���qe(:�kQC�**i9�Y#\Y�v���JF��BXũ(mO���BȢ��Y0e#���e�f�Ξ��W��%U1R5P��ʕ�<�q�#�R�P������y�ҧ���k<�8~z�}4uֵ�j���!�v��~h}��a�
��aV����R�Y�Y�����W�P,� �%�I1P_�����|��� <Oa�s��U�nK�>�J���u��⸻"}'8����Ġ�ozr���y`����Y�;��Ml~����[!�u�i-�ɿ/xM%��rO  �!��Ա>≥#:���K��Lt�o�I��As9.+��H�PG��(+�������*j���e�+���������Ѡ��p�����Q]?k��ƼNIb�~
��_N���Z�8ڷ�&=94�8���|9�!l��F��p��XlxVHYEB     3f5     130�U3��A�O�Gj�����io������[�񛘒�?��N㳏��1�U������dP^�0��M�\k�o:b�+^7{�/x��t��։�b�Pkm��V��B�M �f��ؼ���7?lH}Ԗh�x�ۚm5!X�[�؍(vӵlK��A��4ٽӏ�o�I���^�������IGQP�����z��++��=F�*��\7�<�ɡ�t�R{�J��k"�����Sп3�{�B�Ǚ�zc�v�$�ћ�<ّE �cT��ey�J^��-��ð��*���� *z�\�@����i