��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���rKj�U�_�cZbA.OU�H��0PE����r�C��}m(j�N5��=����-oU���:�└�����&����e~�W��{��H���-vQur��ֶ4'G}�2�"lp���G`��{�M�'L�i7ְt����J�vc�~��q���֡?�2�r#�L��*�`�F:�I���8�	��T�e	�q%L�e�Ms�))��.|L�6�0o\�^�¬"���c�W����K��y�f�=�+�g>���d������q&��������t p���n�ʑ�Ȯ���%u�x	^O�K�L�|m$���S�ƭ<��D_J�㱿�۴��y�g/<vZ/'�V4y�ƏV�����6M���k��%Q��H�.Q�:�S�X;��Y�²�����ɓ����*B(��,�f!)��M ����
 �N	�z��{�:�+.]�4������锅v2	"���ph% ��t�ps�L1�k�F��Ž�[3��JÈ�a�@w��Q��W~�͚�;!�{��/����/v���������􎳘�&�dC4�Ō��7H��Q��t�O�̊l)��sM²j
D:2ҁ ���ib�Dj��3�_��Fӛ֋Wo/֑5�Z2o�:��.x�i�W�d�I�l��0t�d���\��-���Yfۆ�6X�"�-� 8���'8���X�%(ey7a��¿��V�UOZ�|�9���������{֕��CO���WSE�D%#��`Ey��w�i�h��PL8�Q_���&u�l���i,�H�mW�j?�#���p5G<�\������ʊ�\��𪑚�8�_���2��~��xp�j}�o�Zn'��o)�>�+��_��m,�����\I���:�Y���
�p��.5ua����`I5[��F�>8�b��cv/BQ�B��}���߹*�1G��T+�������v�Tu�v>�9������  �<� �$�:�K���t!lz��v�.]GS��%�zw�;�߈�s�Vk�~�
^�L����Ǩ�9��0\R�#C*�H���k�D�h�Xü�YZ��zI���6(�?�'4Y�s	�f"�|s��!I3��-�n%�2ǐX1��B��P����ڳ�o|���o�y��I�b�g%����`X����-�]J�劬$�F����q�	���ܡ`FD����U`�k5�Ύ�k$����Ue͘�X�ؕOϛ������& ��%G��ճ3#HF
/\�Ne�K\�S�j�����pf�+��1:�M$"�&��c�Q�r5�!�����66p��m ��t�th�qn��u[�	�d{a3k01��7J:-]D�c�N`�Ǆ�E3P�������q�)"�k�� ����[θ�@)���t�]X���HL�ғ
DSmz�-��?�Z��KC�|�r��YY*�/�iC �H�"����)b���d�Y-1�����A�]��'���.�3���R�(jW��H��ӑ]�̓<���6S��5�^r�d�l�͚��6%��F���ڿe��IM;�Q�a���̐)ܩ/*��{q03Dv��^�����!��,E{h�mj{���ݐ�9��n���?$�kP]�@ߐ�Lz���l�~�a���ϾK�H����I��J��Q����4TYJ���P�e12\w��D��DG\Q^b?r�`���s6)N�����|�+\�ٮ�b��R��|eIJXC�ƕc�п͖=�ˑ�v��L�C[<�'����[�b�v��.�/�5��k� +��#J�ɔ�|��k�_��E��`��eh3��,���z�G�)k`�䉂X��nz�xHB^)y�L  }��
����ߐ4��[Ą;y�"��i.��@_����<�*��M0U#���I����rأ9O�@��ĭ��M�O�'��5�q��l���� |Twf�fN�Q���K����sĠ�\ί���K*G���D�0����(V}�>G�4�׈F�Y�Zm.�$�䡜ȹ�Q����އy�&bP&Q]��W�, j,:�#��#4�1@d>��b�Jxs�����������JK"	D�$�v�Ѕ#�E�5e�!T\=��0��ط�׎kb��Q_{R@�e-&�rc��d��E���4H��V3��8���̜���KW�H�I\-J�z�ѣط��[��ad���~���1�m	OHݾ(�;Z�V����9���oZ�%Z�L/�|r�����ԫ�M�'Stl���&߳���x+�*�O���)���4�;]���r�j�V�Q��oi[(yY��-�߼��m�������Պ�%�g~/"���v���0^X<+�f��U|�i̱�)s�G��t��
_a|O��!6Ҟj֎�Vd����'��zÎ�<�o�N� ��ȓ�h�?m��.RQSl