XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����j�t���gncη��u����������@M���K8!z;B2I��#ZPk�L�CX���3�g���(Z����p[�qb?�D��!�M|5>���o|JK��0�4��jNpWX�b�Y�XVo�#���/�����(#��Q��Z̾|ja�MA+��*��c�����O<�ϴ�3I`i�����;�Ӂ18�ݒ%<��*χ�F>�B���_��mA-v<�M��NyC�$B˸�%h�| 8����?������Q-Q��r5&��i��Q)9��5B_E{�?4�SFWM�A��n�@��~%�d��V�q*��(T�t��ԬzQ�k@j5�*��%`�I���������������d�:ږ�$/��s��L��p�q�B_��ԑ���� d���9�È(��/^�F�Rq��ƹY!�����|�tR�}^yn��|��*�Oi/���x2�0I�^kAuy~dj ��-wbL�8C�I�W^A�cO�	�z����s���c2U���9ϥX[)̡�수jh�ދ���w��h���Zá��;� s��ux��i���.~�i�$��X_�%A��:i�a�Z�ȫJ�a/��������	aM`�R<��z��8n�$@��L��t���f���ݥ��'��5�,�����>c��y��7���8hB��
��
����~�3�R�S��Fjp\i܁��}+�`V��xab�r��a$O��&��3��y �{��M���U����;;�q5P�4XlxVHYEB     400     1d00�P6�®6���]����h���HU&Q�Ep�
v<��:w(	��q갯��<O��� ���w˸���̓�����k��kZl�w��NO��g�����������K��~�����Γ����_��2e�T�2W*G_��Z5��jq������:�)ٚH��3�p������Z�{j��-��q�3&!8�+��z��6���{q�њ)Jv��m��z�"�l1ۖ������Y�4� $�����W@!��(i�P�LZ�� Đ���<!�,��;�J72�6�~�KfQ������E�QT?������Lr�D�w�ס_T���^ig~����qn�تOB� з��e��܇��n��^�/�;�8m'D�&��TQ��6a���y�]fҿ_�(�U�:�H����e@9���p����v�������p�31�=,MXlxVHYEB     400     170/ɭ��A���l�í>��oq��̓�9��/�<f@]���a峑�4����ף����%��JS.?�2h�"2^U	��i�N(��g�W����� .�歼N_��%����^6�˺ ^a�04x�y¸�������]�v�3v���3UG�|bBp��uN���뵮EWh�2��-r3<�-�k'�BJ�>l&j}L 2Ѭ�)�?ަ�2�U� ]r��;Ȫ�@�0\}�}�w�-P�h��U?��/c��뢘��	�������Dː��	��+�\��o���-9��]rM��:h̈S�q�iN���|ˁ��)&���.��U�d��?�{���Cp�~}pN�	�n�I$a��Y��Y$>f�T�XlxVHYEB     400     130�����Ŀ~��^����d���S1I����������-�|��B���Ԧ"L'NKR���a��S�ͺG������78o����3�΁t�\�M��ay?��=�=�^�t�`�Q+�Q��ݍ�OM�߄����r&p�u�9p16�гPνe�a33� ��rό�!)�k���W)Q����i:l�%���"OR�,�������� ���)���̰ʬzm�?�T
&0�vw�`q[�wN��e�x{⊟o�S��͜��XG�;m������Z>��j��1�Ơ�Q8��ĕ��ɶ|?XlxVHYEB     400     150%���}���P:T2U&N��@^��A:D�:w��UH�|�
�ݿ�U�U��:�BQ2��h8����d,���.�;Ep���!���"�BQ�_љO��� ��~���J]<U�-#��|	�s���� ����ezV��H�yH|2�	˴�=B�
�!���U	�ufb��ƽ�(s�ˆH=+ٮ�a�ݡI��'e��»��<|���]��x�l��^��_�M��`-�{$y�5=�!�����]�p������W�����-��
�!'j��!�%��������)����u�cJ<���Z|C�iE�9����R�{��~#S��+XlxVHYEB     400     190ժmHKL�6���3���}1���S���0����l���)J�pl'XSw���$�kwk�T1ʿ�@�r����c��2����Hת�֜�oy�#2���<a��꾎f��6">��TsAt?,�5��O�-Q4#��P�챣x�H僸����XAg����-3�]#9�v S��镑���ۢ05EE�����Tz�]<�@��A�h������eVi�,$��7σw~���9e�n%�'F�ŗ"�)bLaD�B�2��tp�ܼg:Epy@І�D{�u���HGK�R 6<� wP�8���V���ҹ�5� �S�:m��vx�_`(��$ˈ53��A���>��a���D���H�CoDp]3��zR�j�cib��ov=�� -5�XlxVHYEB     400     150ݫ`�]��UQ)��	�������OnS��^"���Q�z'�5 ������~@ݺW�9<9�����S��̯�2(y�Z�X0 ����+H+U,�W"��#�D�ї�b�Y���)5���;�@"����]��A�:���ջ���7��?�w���Ԛ�ʔ �]�@c�O_L\0d���U�f%]4�A���Y/vj��N<o�c7��b�C�
��W4���=n���B�������ӏ�J�5���7�vC2>�W�ſ8DCJ��Rqw��ȃr[�"Ʀa��x7�c}]p��O���	ۼv$����}獋�i�
�__n{R�[XlxVHYEB     400     100bt~P���EM��}2,�C;AC8�E�Z��O8��诠7�H4��ρN�z+��u�J��
�^��U���8��zs�62�go���ⱽ��՚�\���GB c��mN7D�e׳��c�ޠbk�!	x���0�l������=���\�d�rX����E�sAJ����5E]Qa(��I�1A�S%G#]��c�gs�+=�1aH>t�{}! �G�.��ʋ�1��z�ͦu�I���P���9�pXlxVHYEB     400     160˄��F�g��'�'��>��8x�0i4+?�[Y���ʣ�3z>��'��C�2]ŀ.���Q���ZEZ$��g���)�t?HjY�O���a�c�=F�y�I��m"�Q�a��;~��Ǯ��l�Kg��)T\V5�i��~�D&�'�.>�8���a!%0�8�;ܲh��ՠ�NS���`\�B��zV}#H��;L���P�:�#,���+�-;�!!��y��u#���h���V���ý��T��R����O��f\�,��e�%���v��s����3"�Ё�|����g����e7Cɮ�)䭘a�M���"�Jn���@E
��ߴlc���܌��C`"d��<TBXlxVHYEB     400     1b0���`�#�$�/�N��M*���w�-_D�������{��s!l*�����M���B�zoL��Ũ�C�L5���^��tk�fr�ҷ�U�a�D�D
T'�b����ԢvWH�����e��	�j~k���+3P� ��"�9�O���'��=����q��Ź�Q9|?b	?�,m�F蓌�F��k}/R��⢹`���Z}���^#��e�����rݑ613�����)��[�@W��#�D����J:k���m�iGf�-UZ�zZ�#�U���2���6�q���Ld��ݮ0��-�S����צ�I��	�y�Q�
��j����n�� ��Oi��Fg�X`��7>2G#ͱC�=;��
;�FaG��a����W�*�l�l���C�z�g%�Ї��0����:�]�Tot�cI0��XlxVHYEB     400     170��PX=�H����p��7%��B�6��WȬ� ��XO�w:@#"$m�"��,�gh��]�+I�M�q���w��vg��*Oǿ\����pXY�S�54ϋ�U����bP�<�5%�0wȿ�Yp�'J���yz�fP��,V]��!����'h�z��\"g9(ȭ��jy#r�d!#� +J�g'���)��͚/by������F.�q��b���E쎋��ؘ�M��3*�Z(�f{��Pv� �g�=	LwXsS�'�W�Cˉ�	+W&|�,x%X0�4J�@�,��&q�o���+'�k���S�
�.x�ȵ����i���� `v����k3��k 6	?�8]�2@~X��5��/��N_��kn�oXlxVHYEB     400     1b0%�x
����>�H�;;��^�L�d}-���M��5~x|Is��"���k�$r�e����u|��X�Lh�$p��̀	>^�������f!}�0qU��h9R)L��8����c�+�?).w�A�yY�^0�t)R��$���<����?�-���JI
�|l}ٜ�*2m���X�0���ʄG�j��٢��F�g�K;�ΪsuF@/x�J�"��(� tC�̸�S�i�����,T?Z?����i����D���TJ�#o�glX3\��a�躤
X��r���Ci�J��W��DE_�=��/���dWȂ�W���X��b��
O�$a޳cZ����[+��������R1�/�-aJ�km��/�R��A�hh	N�����r�wF]���fƖ�Oد���1��'�I����XlxVHYEB     400     170��U�N���{>GËr(�y#G�Zv���� H�g�@�ÆA?�9�:L[�M�O�7��od��ގ�,&���5�{< ����.
z���pX�Z��TIڱ��; ��t!M�o��FW�
Ρ����KGz��-�0�O�k�Y�9�G�6>�7B%a���'��Wם-C�`,{�����F7q�Y��}W�f�~�?��L1��[!���lVM��s�K2T�@"|y��'�bZՋ	�1=�cA�Q`rn��y��q��0ix�3H'+p��z�c-qo���Ю\���P/}�vV�3���
�C�C�%�Gc��*�����n����v)^bP�X��o�y/�ߚ�mjʳ��^Q톝��iQ��]�L�j��#��XlxVHYEB     400     170�d�����tp�4��Vt�/��F(��W�-@�\��8����]�qg.���\,�:=����۽�a�ی<風�Hp�G�7UK��w�7�!�A����{����ͦ��:���:�$��Ƶ$څBgf�
=y��+��ЙZ�2�l��������C"�'� �G=�<n3��i�A��DVf>�$X�Ɂ�rH�cd��Ԃ�}N%�|������WZ�~l�`�=ۢ�g`ǺD�w�^�@5��?�X�9f��̉�����K9�����z"0�d�N�Ÿa���Zb�m�$V��$�l�	��(�pB�_|�#r6Y��Eup�`�(�<�=�1�f�?",���@�Դ�o!ƌn>��u0�M/��Ș��XlxVHYEB     400     190�B��l����gy��9��|���w�U��Қ�~�Tj0��EԬl�s!�?�G/�)d�G�����lH��
?�
U�����"OE��ߊB��c60��P'KIZ��W&Ի�cn�����
n�m�Z����w���.�{6.1�*A1�%�"8&��r*d�+2�r(�{���i)������Y̮�َըe~���>���U��t�X����&�f�}��L����ir��}Z�mT�eO�+��|C^�ds�Qܭ�v	�*�0�3�X��y?*7<+{:�shi?�Dl�0Z�0cw�wf�$�%�P�O
�9Me��);����
f`����]��[Tz���fb=��/�U�]ѱ����@#]5`�!�]s���o���Z�� ����0g���G���T�aYzn,�XlxVHYEB     400     130D�WC|k��Z��+��m�C+��`�������_à�['�[*��E��������NpIuV
�aV���x*%���������~��9�02h�U�i�����X]��	Y�Z-{��aO �x��c�c𯅘}(P�w77/�ZG��䙚n�*���{'�;�%����L�8� {-XμʧYu����7-G>V4���1�(�B���r��>'��u {:V��l6!�� �Ǽ�oM?�{���\m�<��b�w���72�����o�_c��
����*u�g��A�3+�lL禟�XlxVHYEB     400     160|����e���d؞�Cd��ԑH����}X�,��0ր���3C��P��a[E�%����>��&8Keؾ�/T��˟��G$}�����*H�]kѷ]iVNM�Y���H��B�Q��V%���Er�T+���;:�\��ӄd� �x��M�ġ~�	��B�[֔��+��XnzS�����fm�d�/��ö�EH�(��~(>�v�(��x����Jp�&=k����u��&�\���E"z�:�1�Z���˹7�(�� S	�̌��L��M��m���;�F�_��ޫD{�:k~���+$C_7��S�a�m�jvkS���t�#��!'�[)	r;&��(��,^�`g�XlxVHYEB     383     150�IC��IέQ��>)GD�p:N�_QJGĺ\.���2/��5�?��jlm;`��7�]o�,������u�rn����t(qz�n�7 ��n�"�(f:����-+k��e`�.3ԔR��,xc��yP��W��}��x���?�奏�& �jI�﷧�{kԛ�]�)a��>�|�o�i���g�u�/&�HD��u���/OaXF#�U�g�\��j���ߊ��u�Z��a���PMs��9)sXa����o��@���Maf�N�i�Y=��-�eߞ���#��ai��$��dޒ��<�lg(��|���[>X�
$�M�e���Я���Ri���