`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
X0NMbWDksFJ6iTSTLu2vn0hRWhMIRkH6NW2XJheWXkFw2XuO7DtPhbHyupWQif5j5cgLo7XShF/W
JT5djY1LmeAZdmmoI2o/9ea25XL+TKBAqbpSvWHCdge0gip7BMYELTW46sFm0QFGwU0WjLZHqSQY
EdiWpN6JOj+pPsQd7099PmsdyXCYWvV4vs9d7FBMNFiuH1WqAN9LLIC5qh0Aoxv/yNC7+jEvI6LS
o+vdPf+RhVl1XGmQeRxemH4esRuxXwvHGwbMGczybvYRo6b99EdqMww021wnhSYM4On6zQfBRAvu
2Cs8H39hDYryNpXmHDcPBUlCzOypoDG6DuIpDQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="5IvZgbSSOujFRIZ67RNXUOrYLNDsChcOePd5L2i0aFY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12736)
`protect data_block
m4KNafBjG/FjoYkApogbzIYXjBg1sLFfGWUEdJ7DHlNqMVAMlCJJmfwL7wWCcICIaalclEVe12g6
pQNsI7kEfPJNXMDDt5DhLVpjduyFOedq/0hcA7k+jZY++OCppAmEplIUTLZ8WIkWnlAAHVGNY0kj
vS63dcbvHtRlQ/uOb3KZVtgWeiY4qXeGCh4Aa9IAhd/VBBeNi70dEMc/4qURLWQ8MZpttR8gs+Et
KMVRJHGS/8AsFULkD6PHux1Ni1LJPwK1Vn3MN3NVp2CCSQVTYgApGVT5ZIWJG93fhgdK4X9QqN/4
UafkDV5hCmzA6U3ZVkfRBGf8ROSuAsjQI2sjFzhcX6Z8OYwDU4c1mVOEjxs6OzOVBb2Zlw+pZ/RC
tm+7f+SJrdStXPFX+lR8RU+ovH/bHu9YetwBlmnM6XQKUFHimDanG52ZWiwcGChNBxZPAX6OqHuX
WdJoIL21nE83B/TN0OrkyZHFogW4Rd4mw++oH8rQP+CavTO6T1IZMdbvSKj7odEFOp2MlPsnMdrk
d1eTLL5ffaDT2muP7BypFQLatZWU4OpRZcWwq5F6SNq3HmsoT3Undw6KiWgXgpni/32fHJaoECYz
/7HgaftvcOqM9V+9Al8k/fkkOEZ0PY6SfSqsmkMuGUNVotUyLZK2DSekzLcN9GUcObHCTECvPbN3
aN2fzQZR4McvdXOqqIr1/4X9LkVCJe73zDFN7VVnfcjRW8TCTBjGonJN/CRQsKGsif4FkDWBBpSb
0cqUTlyWBkch7rYRIVzWLXa34nEkez7TBFPWuDqeL/dAcdfKSkcwnluG2LBiE0SBRvJ1Rhaywbhv
4U52BzKMTeKQ+NK7+DKdG9STOgkY6H7LVF3GW0I7I2vgSG6UY3Cg6GN5iJ/Kns2x7/im/fv3EGYR
OIPn/7AQKVXkagFeXeWluy/bI9Auuz3UAv1mO1GjeXNCKCLhoN+CtKdg/254zLY1R4EvoWFDyyD1
VLIWmyuGweHHMl1sD64p3LW+Udf8CqSIBOB11CCwEBGRgjwslnXZ4TPA6Hwg220wz6K0nwwYl3tl
6axPKXOhR40NEnmge3KDDr8jy0pUvncwaaTV9m0WKJyt+WBFa8pisAa/S6Ld+BnVCkMImtj67DyE
kjby41SPO/mJ/e3GziL0yLZPn9uqYy5Gx9Al3AlB74zOHHeTnhFS+hYzmAROlg8sj7QaUEWVlB0b
Byr1dTHDeBbI1hkQnQNFfJEIO/95T1+KHeWjp2fJc2QHs+3qYslWAJBWsFuvf4PRVJZTgRucYung
fkDs1T85qAnw5RIGjELfbl5TvUVDTInAlgEy9LlK0yWEqToGQU/YKq529p6EPmNt+8xWoygbMCqM
rGvsOha+PWgUGLSwlWyhmDz8E3XuoyqRoFdk5WHT9qdGT556JlAlt04lcHwUBBrMFn2ngZ/ybOvV
DU9gYB1H+0vWuCfdRBcb9NiM8riy5EdVcpVce8dS3QGksVew/9mj4N+ql/MDn+Rw50/k+Wcame6u
sZju8CSA0Twe8Cc/7K/EIHX2bzsYXps9K3+FFu4w+Ef89VSKfoGf/zfc4SsU/WgbPVRZN4mxEli1
25FtQ8LYSBSLYGRxW9O7dWvLU81xHhHLivTfwaki19mHxVFSNDiuywosJbYB1CjeeCaPOqM+kWen
LPito6PFb/1dJwf8ZbIAfYr8xrM0pMYkcVhu0erCM7sBUyu6gsd33VSpDPky8chshODmOTqooDzZ
XARy+m4yNYATI9drYMiAZR9SeDGYxiWt/D1Rx0xSVdumMy2mf5ba6q3F87BJEVFgw/hVQnoh/Nmp
FGn5Jg/H2J+qzaKcdxLPN2qMxyYKUe3G6TjaEcOg/NgI6NhU1vyLWHUqD3Htzcc/7rOHdrlbms+A
3OBzoM/0ZTql9FLWLaCoDjQNIG277F9GBB3xQqzKX20ni/7qBM+OwvjznZKlQuw7ORVBNx+9IlQU
SE4q31w4RuGrT6F+poUSR6Tegi4E03qYhQ79I8IBeyrdjcnWeewcx83tW2+yOc0L3dBShZcFyQLz
oIqjinsP7ooZKclR5IkY69FM2iLD1LHqw1IbOGs3aAeaNWTo/Hex5hkzhrdFTdZ70PSbyAwqjo5B
h6ga+Gmi55bhTwxroIHWw0Nw7FeKNFsImvmDQGCWE/sD2nBk7dnddtnfWWIYjqrJP61Y5qdp26pG
W3SmyKq81QK125r3Wg2JAe/Xx4Q73u/TwaiJ3yy/A/SogemYrrSX0x9BUYiUTuyQ4Cfp6GA+eDfa
j1U6LjOiOqoVUXR4a++MV/rgQos/5xA1LAdULe/PXc3UJFJxZ/pGhR/KEMKxR1OkYp2/KSyvDvOS
9wxtEssJBl79WL3B6tcVXfnMKzyNcUqrX1QaprXbypy79ZR57aG52epnDF6XRna+4EaR+zszT91H
/NcpcPDGZasDmPNVRWKu0B+TB38N5bA7fcy6mG+vj1DQ+H5KuyElX64fQcYqeTc1HMVnMltlIhjJ
2I3+WLeN/WuytFt/BSXbAoUxNoYlAtL0JCT2B2f3TlADJZBL/xi5/ETibLoRm0otqmgszFDfZAU5
Gm6hqTU8YgGkWmDtTDbhe/o7mbZ6+DK/xdadqdzkDnLHWds+CvusR2XIJBVnN4yrhLI8DgJtmpkN
eNNYSSbBOJ+6vyWVITWUSw9S4qwrVnXAgrsWONbl9GPPek8FyN5AFqSS3XumMHjdwLu4d+EevbdX
Lk4LJswsjLk89jR+tgXW3DDJNWrwzNUuR5TWFY6uQEwwQaz6uWpdFGxj9K7X6eaSKHE1aZOhDTXj
dViVS0JXaPYlb1XaNWdgKQRRHenn6qFXPE8ydxklNdZ3cMgSIK/Up/OrL4IG0HeCWaCOnLBTSqfK
6v1dZEZhJBCKNnaNueormA0Peb3L0kGi8ZJZdBuFe2w5h+Y66J6/GafN9ZlEuCjT9lfg2EwdeRYa
18dKPfR3Ubpbq8PtXmAVb9PVYK7tGXJ/d9NqO6VfVw608x1JcXTtP7QH20wf38sRBbipFnPbY8fA
uytHSLlO9G5Pup7faJF3/GtMziXqJLR16KtXwBihU29Zp0Hc+ZDqYgg5fFAempCG9y1LdGSHNLiv
AlrnBrhM0lE2aXb2EblqN2FEDcAz9KwusINBaM1FojO5G5eKNuW4KpirBaf08fyJOxf2PZTBGLp5
X/UyIvb0NpBIG7/wnqXkezsYZK/YKiPGHP/eCujNVkBal6ZYkkAwkbRXFunjnPAbap3cB3Row+o1
jC1cdE+uI/ouEf6pPGFv84qPuA4zTTOE+U7aXDloBkAdZ4v7YbzXobIebgB8ZD2wsoTSN7vUz8ux
dXCTDx/Z9Zq+FKdS6hkXmoAAN+R6nHZUa0wbLR+tJ1C7lvvx6zrhWQGXBs34hQJ7mfhSEtZUT2T9
0Awc5Ooaq0dbM3rE2m1NEBa0RIE6WTW+AS7yRgwFpV64z9QSVeRYlGkfomIQDBld+1r/FvQmhNUf
crR0M/qZldjiveCC6E1Edn6M5nbK8rzGWcvt42pxWBSm2H8mJY5xbRycfoGJ84Sz1ehYzkjesP8/
+1dLHjsYItiyy0PBoZd0pSD12QhabEOEHtM615iJzyBNJMBFjdP+1mt/tacICNCNlW1GQffAlzAU
aG3rXg2Nix2xmVybs+Y+OX6MsIfB9ObSlrKwv/ZLzz5rwcRkVL4aaKfCkkp0Mqk5M+JZZWGWtqNP
KRp3OEMAAOcERb/1pZs+rMdjtp1eVsb6foyByJ5RfORQjGEG/zD9YpUBnRPifsn/+I+G9R6JKa7V
YL6HNg+c7olOkIiwK0gCeeVVRrzrwRZJv8CFRTpD2N5+ddHy8LzxnG3Sq0/ZgNGWnRpvvbNwFWbt
TsU0XW53avlYQMctuE5DFC0ywvhCDAp4zOVblL0HC/dbv70VZjflCqU11amiYFgE/viebBgZzsBB
8Pf4Z6Shw/mlfpnI9fUNPVOu0ZV29ry2vsd6JUoFLuPAGDa/5W2YbZz/DbbqMk7DoFOAPloEtULj
y8VIiUw1BqxudwhZuwI45jNOCMDVyhm247xD0KaEXFo9RKpA15BWEfJDvabUYn7oO3g2+8QYbYds
yAWjclUIsU4iOJ8y446o/Dad88LLRBLY5oFgfJHTA3kai2YksuPPLuVeGFlwz/ZcFvLj3RfKdk0F
5Do6wvfd72H0uIz2XZGdPeQWueHvgzbpmdFqz2M40ztmTDkJJ8U378jVWZ34rgRNWjLbw7xokwpe
N+H2tIbB30ac0PDHwleBS+9WH/+3yWHLvPZoj3zjgKRkBhDAwhjfTa8XYGix956bmC6ftAZQDLCP
JvtwpN0QSNc4W9/9vrSr8XSqBZYgnYw7Tr/suaOqwyiEezelnn+wtfHZV0lC33vQH+Eb2uYdHK8g
jaNO9yyr9U021MOf8lk7mc6/RjS4CIu4+aJZSBz7KaCuRTOSa7Y4FT5ziv20TrN2YH8p9/9398up
XoLA3N1g49fnYq1Rqi9bS5ETuJSDNhovAIlwzGavyZiF+WUVR1lOtnnhvOmabJER5RsaEu2r6vdC
0r14rmrGVy3+BV8+iVjXCb7Ars4sfOEFk4F3vncg9Gnx2HvzzYmp/2oNlLW84hY0xdPX+01Yw+M7
EeGn+lbkRHA95JYwSYTLQHle0tEgFro7u3vqP85EqPDqY1lwMienp7E27bUZcLxi4llBgeXfNZ2L
dfqT0UbU5HKR4c6VT/gYr2V2aOfjgllIXm+0hO6YjJADEGKWIDxejteHI72dlpnlT9HtkIt+Gxxx
408JJhqKGi5bqLEBMtwKkcxAarbTHT6NhG7ZUnAYYMYvw7GhukgcxDZCqZAR1s+o7j2gWVF7d9V3
qfCM0FXOHzGWNU2kM0fireGOHDEftbTaG9MRQ2J0J1o/DfDSaqCPQrPdzDanxctIQR8gN6zzI+8w
DeeL51lsy413tZw+UAXc3iPqr80J3yZUndtmgj2MPWORQHqCtdx4Y7ZhHSDIEiDPWGLmAyBwD4G2
heeMjLCOo7BzIxgpdjmfq1gD7xS60OBhqk9FdV+/xZ4G2OeEbBOEHXrTOwSNq+HqxwH77aJzdOWa
CHRpn37e7wL3tLHvlZkzUjd753iTGqAY0UgG+Yu889JKijakzK9bDU4c6AUmRHFVDMOWe8RRSh28
KzVnnpVFsvUf7pLYIe2SOEt3JqZNOg1g+pY8VGkwbXzlPG3o2DdgTIPneZTGe2UAfpAq8ZSJ/Vhu
9/TzpCpgSG2dy4sPaI5y9VIdsCiB+teVx+U03k8AdjWbk5qsvUJlEB8QulzkUxBr9vkTI6JA/MbE
pxuS9E4ZDdnqxOENYmkV8qd6PfQpw2TnD6wyc0wRzQ7BjW728ISNUWIoNrOT13m/fMzdcFjUpAG2
H1MMISzNemk1Yx6rX2BJZiz6eOryWwYCqAeJ7Csu7ZlZ3ouAS0xOwk1Kcs+aBxGgKwPUzoLc9/oZ
iCehtkXRflzQkNVQDgKZLSEEvszphDlH/kKdIdDW8dFNNtPPINhs2o33w5N7r+Q6MqSTmFmly+UT
S62uVtDxq0A7lcHjorwHNN7S+maAi97aIV3iMoODC3tpfHfXyDvTRVVi/o7rpNPk+6lJEy42Odug
2EPrS63qHtCr7l4ynXqBnTVlgexARig1T0S0HH1PLw4b3kx9bbueYqjw5LBHnPoYe6EC94kg4j2o
Hqc1DFrPnWGkaGff31e6SakiqmFH6k2gBiZBi1Vx9SEz21gPIJ7IlbGFs62tIeqtSC3fAc3t+qAp
SAV/k5UfatO/YlaPhDZSgeGGgxFLAqrgi8Klq/e7lBSQH6m86ZnFlqiDkiZW2CW4cr5UecqbccSV
euKw3cz4KqbpWKMQfeCHO0wOoA045oPKhUH9OQbW+togFXBr2EkQmykDHagIiY1XqQxkrI4HNWaZ
ky8fnBywfE9l2UVAh3XWE2T9O9iHD8I6MhWO1W8xELrKHwySNuYPs3byhbRs9koysDiuwjGxgytn
j2G6Qw14b5HaLJTdOeORHQVWXBJjLFOsRlwEkX/Ghp96ZHY1s5XhaCA8b0hvEO6CkyaL03AiE7qC
Lz9pPMNfhYy9uR3y8bnHfUUyJVprx5Jnm1pfMa6qYntnpETI2sMoBXDZzBmaVdJ5gxZPmlYMwsCz
JNj2SxsN+i8o4tcqvUfFDN4shyUKoqCHwefkKWthElbzd/2ZRLjwDojWxpbqIYo/JhUtqpr4Jmd2
+4t2x1lOskvn3bzP5PZVAq+p+AVRlxnt8fC985XzdCqCfDj5+3EiD6V+Rm0ZJREwEjlumUnD+z1R
nqOkhq8bv91GF+zArepuC9ndIg/bQ+zoIUO/mdOgI3HaKIpMxByNAOCbgi1hyD3eB8OadUb7vmq3
thU3/VH+B9GjySXBkSSpgpOA1EKxlkKFxS5emm2RgCckfHjVj64axWnv7z36mnfHpvAPX0ROs8mu
Y6Plnohns3awV1zfoMZtYZhkH15zvVzVXNnSgGhN8Gi+jin0V1ZwY45tvEpD9OBC86og3NFz/Rb5
D8EsYXPYKqMmXsERZBPhVGMNJVtqJg4gCEYYXjJa3UgKJjyBRWvQF6ljCgd6fWl2gfy/o52h/thI
QWG7IIVVP/iHc/F0Zttcjx58N0FIvH5rXkNgrlCmdmnB4qD+anp85Io15tUPEPHeHGVwhnREFrzJ
uko8RhzaymHq6EMg2VFAYZadHbs4KxFLf0N+D9bGc/zOlWM78B0izYK1hJ7dtCa01/rMTRw1YKFG
voKM2wkMcWoX71kLtyPM3UiBFfsBjF/fDOdwnqj2vkCbBSKK7h8UU6sfLqc9rhtjylpQoESnZiIg
xC/9FbjrgzGBfEx0Gw8WECf6EymUbZOSrmzYCrBbfQP0vJqBS34/7EJTYmWzuEG4p7QtWrWJG2Km
pidnOnvmsm6njtrM8AOGaIvp83CLgcMSJdTfvzUxvnqEk70yoCJja1Zg03gtw+feZZTB8Mp6o5iu
40KgZGi6bZCvlITBXwwUIJwdXOLzGsIU1f0NETrgjEBRkHXTXOL8De+Egn6lcmtCmf82d/JSq5v1
hDB3O9XeZyDUoAZGHBWe31TNgC9/OZReEcbhn0VxydxVMPRNSVVuhg9cM3nh9sBGkr5xtGENrSIL
zInjFQGagGRuQLwjTNst7eWKlrKE/PfynBGseNEoueZDoBJL+ksxZRmlkasbPzb4xLRj2NBrG/R0
Z2WxnhjrUQ1yYAtOkXmHTmFTNxe5Xvj9cHAwr0mMR9EVD5BCkoDi/mWaNNcSj6SKdOgxQ05NzwH5
E63yo7wq/KElPojiqPYKjjVYyGmVLKuXyD3bx3tXCN4D8/WbSlQxGvXiMuG8ztQWZPq5JDQOfuHo
U4ZguuRUMzO8DFhJqCkt21kFy8ApeleoCmIalweWArgnhio/vmMgoBMiAtQ+lWRBLO9OBPtY6EFc
zjV+kapABF/yHhVE/ozjJ+T+pn0W+r85csLFLwljvV11hEh0JyryNcwy9XL/ceCSTRJ78kkWg494
BeXbZIEVBHkAhpG0oOaL8Ty1uGual3nAevW60DuvDRALocueoH97lJD9GbqaKTEFQ9dGx/k8p58V
SB3Ur1cf/KuuTDP82m5Lb2WogG0CJz+AAgC79eiqTrn4Qc1VymhT885fOKiOFx1veZZVMGfVvelk
fXXMbym8RkDnqxpWtzkSXLbjrQtdIZcgHh+cuk8dzrTY0glkfgTGT2ChvWv46JiRrQe5bUVtAtWK
y3Zc4yNNWfSZcoECqa+digLHV+2/mtmOCBgThuR28ecG6Jn2whoRaJJ7H7IdS/A7RZae29itZD5P
zQC8b1WagPDTU3c+KkiLyYCMNOhUitsIsfoqfu6aAgdGa/bI4Adba1lcyvcNg10Jn0PjDTzMtXUF
YWeialT9yrx6As/TotQdC8j2MPrsKE4Q9A554WnuH3UWw5Ec+5LrMwZYe9FwxxYXAhNU+qX1UfQv
ndlKOStoWwfawmOujLPRZACksEtnpSScbDJf7cFszE1xRZRbLJMT8lV+0QMuHzfy7zrRj2m0PM6w
4y+2KPh4poihCCWrJJPAFqDO5Kr/4Qj/9mly4cnmXBrxzO0PCqKQpk/bqlO+E2Euk/r3UKD92HQp
6gbKz+YlRT9SaqXk9+vj3/cl+H1WXWehDSfAmGSv8lIqkwZSzLhlrSVr9V0q1ZGTYspYbQyPrHFR
9LYKcg5qKlnc8VxBwFf4XHnDS18seAlavnlRZlUR41TgYVT9LTUc79Zlxxy/KqgosNlKTVEQTYRN
syOQfNprGPmdk7egtR1PzDOd7Hnt31aZtsi2IhmzKfcLN9fyFhpfI+MS4crvQg4RRplZaUc6IyS6
+vKxUu6EU14i9PcRYB/lNGkRp2tpFPO1I3AH6cm8GQIfj08g2ZswOliTUBSx7fcZZtyuerZGnGJq
50BCHO8xQm20bYEduyouhxFG0FjzrUIcPy5lVJVfqH2PDFewSWQfPIaVdoxo++bW1MN4Oqp8WLJg
YpR11zEvjxhomFgNf0VJ8iBJAmYQjXBfgnGYY+aHMI8dGCES9l2HjarGj/LDqnsMzm8iJo9/H8/8
afkDNtdUbCYBe+4qCpoYeB+WbN34hwNNfHoX/Ocb+buOpjoStZo6cL6u7/ymHf/+HmJAbn3VywC5
NFQtDGqSqM9Ym6Ge7pNcI6t5JNTTiAb5YoytHD/ehHRPiuGHkFqR7g+Ak1E6/KD7PTD4a/uaIWPG
cXqdQHVqLXicTCCtiZ7+3mvYTDcCLtwUX6n+NXHT6jhM8n4v1zCwosnr+xuuzBN/nYgpuHj2vaX0
4Ji9fZYGVQ80jWvtrzB9/o5RiUQAFnR/tJXnrcD9o/CG9RcVzxC3QeWtW+oY/vuaowaxtdZD+h4Q
q4fNA7WW0XTWx/y0oz6DPJkP7pQ9GJ0QGzLPKB6N6D17pE/UFzk3+S1tg98sA2F/O8S1N7xXEDIH
29FUoW8Ft01R4Vm9FOtjQroOdr2XFpMy7G4nHSf0qFNiNlc5jttfX4CoSNwp5RA22okmogsXxMMd
Ua2CmBAJRD94ocWjE/llwClyMshFXWsVHZa26feoHnemcG1VCpCQSlGWwk5HEmo2FnTmpGoQORzP
4pnPfJCmTfCOPtc4VILeXTRn0ExlKKq5FPC+ld2EN1tnIN1bGuiHnrAV0YNI7Sjf/8nGpWJGm8yZ
KKhIiLCERy2zH9KzmSak09+wFdnryyGg6cOuFxWvHiZYHiKAijYP/mfh4+quwWICBUJIw3qMiUb6
dJ9P6qLe6ylygknCeTVpLDKvkt2dnwr7i+Z1TN2tE9C0AW8tzV1zPUUU7NU/iLutH4QVPrj4DOHW
SGZcas61MDIpSfuPaiL5+cK4sbgcWHCd0pZ3lH99wtK8YarloENYxm1Pcw9e2/XZcBFPRtseZElC
9M2LExlGfSwVeozJH/q9Jk8f6BicTmhWt8Iu5HoN8mSUXe2I7M5H339EHzymn0Prn94FZqZ0lU4P
T/KY67VV3STjyeVTOa4bfiQfeduTIVi8Ev95sJL/P4IiAlRBmKpp/Sbupe9vbj4TC/YlOq3zxg1n
PgrTvaZOo5m+Qz/5+NyCxoz7gZj2JGdjCplHZwV4/f7cu+PXRgdqJCh1YXwjr1f47S9kx0EkVmAq
ptkUWCEZTaSAgCrZae7VclFriAmQTKgdPlsqh0PcQdkOaYvVlHlYyvJydoJge6lx5nfPTbdolNdT
D8nnNGiEAbHksGcau90KeA35GGmW/N5M45aDUfNQ+BQWqWAsdVdENxq8RUdclauYLRWe5v5tXCJe
4Ffi6GdBzpqVL6fbI0R03NxVgM0Iyr1/n+/VYF//M11CGGZj1id1LNS7VjvvVHCuuMlCU2kgl7J4
2t1Q0B1FeCBhOWpiC+Q072FHrFZCiIKiAqz0EEL3IeM13S9hzGLgWGDouwsSBvWpKgwV8x/7Lbfb
AMe6KI6R5Rk5qBEm1VOCRArF7iAdoYtBzuXgrtliEL/VAnA/plSBbDU5jCgCKvJXlm1zapl+iocG
cxFwWcMNhGw6EmfAkTPvvxpsF7ZSxejNQZVK7fcig2mdzCxmtpcXE6ZUBOVTeBp9KVGI6aL8l5f4
TGBDWeCI71sj+lIIblEpru+mMcFrd3WkGfYdKcQJ1hIuQd3WQ6+qgbA4K9aDiJcqqNEs7kefRuAV
0w2oL3Ti2NIgz8IUX9anFgtGsvJvAymA2VAfQdfmVRvaN0ZTWhM34Jk6igQ6O1ZsR7YKXmRBMKEr
7gnJLqyAK4KV5wa/1V+8c/FW/z8epzPBzPS7l+IBRCWxw+Lhhqi7HcIrFMw6YzuSF4tF4GS3hDvh
qB7XNmmgiYf/wRaHUZUoUBweN1Gd8lHnlhTagBQvvOdW5DcrHixA8hiJhP1JhKYLL/WNJig4EV+P
Yjxu/+pMlQCBC06JJ0eNZ6uWauQChhkgkWfXV6hUUQPzFMWvrUN89DY7mpMtxUAF9WTvhFVbhXZV
QDoas2Ir2HckGmJd6OLaSsGW/72nDwIXK9eIObpZV3zoiqIfLCAiJfHLzNooVGZ2yv3Mik/1bODH
bneCTu6XkaE2i0DGgrWo4ESffrLoWL+9P3iy0aU9BLUx7D34N2N78GIKJc8BukIaJ5Y0DvhDPb1V
elPV5ILxGHlnaICKzTBUPXaX0xos9PNics6dXGYSlArkAxwF2iTgIu86Bv2iBuoz0cic2ncvGYNv
P+qySqk2EOz262WgaK6/EcboJ/AuWvPIogT0vT2wp0VN38DT5YYp5kVDlBQAN/pDkTrW4aLVwx51
gDkY2NuIFS8cXoJwpGEDagGVyfNGwfS9BFNOlgBJFdEqVzi1ugdqHJipil00k/R8oybyl1tK9szv
u+oWvxIuEXqy7/HJalFzg+Heph1IrI6kHZpmutqy886LhaS1VILA0kC2RQO+E69NtAXDPIwJOomP
E1FIzib6yjtTlFO7C6R6RWlx6QhDMsDSdTTCyNygZpBEgWK+YOeK2vllBnNnkE19PPVqkroBUtfl
IjWgL35t8feHcFU/k9NysvyWAyQkKb4P9Rp1mQRbV5dP9cemEHTTwck28pc+q56nK79SgU4yoDbO
W6mG6hYPq6KLQ+kYu3PWwAMM3gzoP+mgcnItKtHqG+g2933mU5sQXJR040asmMlFhPYZeLvw1UX9
oS5iiPsJnXwTabBqmUZzoqy72UERMcl+j54HWuMwOCF1xWRivPpXUHg+6ga2j3xS8mtwZRX4ZMhJ
aTj7swPMQxM5xvIwHSqPi8nkIx3YQZK2jWz1HdffP1z/RyIwFwUt1+bZhlAvX2re0VSU1Tcs+jZZ
kzwE1Ht1CEe/9DWfks+JE/uvnMvlnGrzMXuvBq3AxKemIN0Es4xAIQ+uECWf6f7vHn+VnjQ4uf0w
pQM8O9IKIaOOv74llg+7Q72eu6kdoL80bWtgxtfd/vQL8JOXe2KwSEuKaRS4rXcaw6DwUMPN3YSa
RcdbiG+fo3U/TSSkqJuCK3aEO57czluqLLyTy6AEZTHkcpQsmEEsM2Jxx1accItsabry34rz8uNt
hw9J6KpCWBbMHi3v/9w8iZNeWLo+BYhI6BwckXrgwTrMFPe7ew0JVciwuqZRPBqWrJ23qbZnMsLl
fIdPc6YSL3jy6s7OHmo37Vr3/IusJWquWIbQeQLr/5ogAPLKyPVyCIWdkjhFS9lMDrQd4Qlw1in3
yTSHDBKpNxXSG5uCMuUiR8GZ4hlDLQKyMiukEmcqxVLSGax5lMBZ5o7AkKA/BpRTiFJ4hDgTIS97
ILkYBqdhUsfdFPVQR5/t9YI8qpXgIUtXgjtL9hnxcIokNg6QlnIhIB62RGWZ606iYYApnMaHP2PT
xH7R/Kr2EMQCO/Pu+o51Ld05CIMaOvWH+BDSpcv3R4uQrB3fgHygUYSDiV4J/2GSEKspaDXoFkhg
10h8ghRpF0yXc2sFxkA78nfPXOpww7ofJY7/1lw4YgFxl6kKOL+zaXKmIwnxcqNoVTD7nZ5Ttt4p
c1Hsd5Yc0XgvW/8qLCEhaNJZek4JGM8cgypUcn9336+MHiPsScvhFvutMh/HAgd3EWnD8i2ZUB6o
xA7+FChqctqJCuOIsJtPcxrnW5wK6AF68flzevxvfQ/u2naHv1VbB7Kcu52V18SaFGG3gZvSqZmv
SGDLsHsCCVxsPc2qWXwLwyMXcFPeIYxVpcwH1pMQpiLQ2cub6fKLhszOPgTXp/kZv4X/VTCWkkKR
bnzLFwMJjCthkbKxElv+fu8CkLuTqL7UWlq0LIEN2iVV2yij3KKxxkq4owxjG+fMdx4o3P1pY8Oq
7NX2ey7p9nqDYzOIJUsUnfxD65jTViMSPuVTiivGvnLgiqOx96VIAVIrllZWbYlAib2vGZyfjeKO
GEUVEtm769pIPpZBIgvbxQeXvY1SHvhZYfqV/3w0ZN2ZrJK5IITfFDxpFEAgkkD6qgfDqzdn3jnQ
WtY/qG/HhPNCuswcweFY26B0u6HxKOE9LMfYoMhgkkw7Y6fnFUboQQ+corg/oqIyJ7C1dlKEE0pL
9UwYnBbBcsiP+P0Q7QZbor/XIF6OfZpGGjoj3X+X7h3aVPD07ip9NA1EN8eKSNbnWxVGWryZ42Il
w7DYNY0eoolmGjLN60aHuz70gaKi5j+jzYehv+q3ceYoNmFeNJSyvjaEAw/sINNFjIzJc7WxWuPr
Iz9klhY97B3RM9xgMK1jDFppPFrvMqw6eV849Msk9BHXdUl3Kfw/A6YoIUyv1/soMEjvuRuynqt1
a83orvK3rtMYpds77n49IKnmDVmJ5lLdh84L2P4cFyFBLvnoQNsDOw3dloH+QLOu/xDsPdct1WzS
38ZgaaSed3SCuRV9u4ws/oadRKzNf4iZl3AO/kQsqh7lsiecQDW/Nj0/6walFQB4M7o93K/caGOb
iESzvaoTopD0hA0VzrPXaRvOpx1ZGdOvDqa7r6yl0uPFUBG/Ar8oqXIDvWp4PMWJkHSTiqdBfWLB
pRXlwl0BgM/MT/jutOQYT/u1MO8PnHpIdWEMxLwKP9MilL5wf96dpIUZ1/e8Ms0b82U28Oblmg6D
xa38Ftrk7EB5d/Cfme0CnZEgbZ7MQrtGjEICEhKXLnTCUSx2UdC3gYIds6V/2mLoe3GtmXPYtXOv
lc8L52uP1dpRjU7c5s0pSBdxFh+p/uQ65S5hZUU04Jd2scRXK8gCuyRl75UN1s/ksCHSpQd69M2d
ltbmhLI3BTiIauthHQ2czptv9543bdqVCL84XUYwLbt7iPmCu53aEpzECOzD8p6xrbXzmXFWKcJJ
ku1yOEYHbaepy2qftiMP5xcwcIyi/19uiELEyID2SMcq4KO0Nzulsxj5MLWRNAOxoLJkdDzuRAad
tpmtMiYiVVtkfxS4VGvDYOl8H3BnsexoabThSJ3sq2DcUayTtEgaD3KCf0pzjVUQsUrR1CM+ROQB
6s/9LHrueUkKrWO2Hbv6nXh0Rq4gNHMD0aV+Vkdoo146u5qrfu/dXj1zZIEDaQJZ61SDMrOqtaIi
DqmG3wiHIIiy2lI5yvrm0qNp7+QWBPDDDOfw846Jq5MjFv8pIAfEIjjXs2MnewZ5pKd6OBtv8X36
l6d8NHprs18yIwUs3DfCz5ItUOJ+z9MM5PERtMrvj6eqq8v/bM4dU03dpMLmvyCW+6kOKf3Sgvdc
Fm6jRh5G7cZpV9I2YmDF2CpxS25BJh9eNeyz3RYB5O4WdvIzQ+Vn+BmSSdDucYZHDcAYymivwCHh
kVfABx+sZ+ijMPPJ0tFuvCebeeAsimIo5jiDvpuSe9SFPEvfZ3mpKx2364NRa7aDjcPRldh/HEMG
85QGIZXdSJT4e4/Ro7z5gPQ37NAQI1rVAvTVsYMmmu+ml2l+IpUnF1JUCTS/OB/E/h9Djbw5ZfMW
Whxlc5hLzF/oKIhVayfCTpT9Tt8j9uTeUQTBO0FcSTbuTI4FmogIL38+5spaEwnjFFq3AR1VqXN2
oyAAcTttgssKXzggfxsAj9VRx49V8AqRhoOTNKzWmPbck4/PCRExwqPkwy/+Y/C6Juz809KWK2+G
KKAed0bDlnBi2uYRPZcJxovaPIfBjf333PkK1jaBfKNg1BFriowmuvhUPeftMZHt5J49BvLEVD95
z8QqsWw7cdAhb+Lmp4TyCq1VVLsAN+HiQa/kUHW70Ol+OpKPvVCEvolJ29ob1OrPf316CC1CJLC5
aVUjlfz5DXq4+CAQXj71fBTbjZ7dovp/483nWFkfwTLkltkkyvTUqw2hNQYZ9HcpV3hlsQ4vBNy/
jwn9p4/nzX0YOfRDVleutrlIZ1yWACNiaheWjbMbSnhu/gB/vJcinCR4SOR/+r3rvh+10PAtFMUJ
q1tokJF4bL+EHnnBv1vAdQPyOU4m09CcE0WJAcJNMGSB/xgD3qc/HWsfPkd6Dk/e7BUwHKOH7pdE
XVUyNggBC3UT6bUQILumxCXU81cDhQmJLKLBJXk9224vmvNQk35oKylDR1g4RzunboIlL522h6UC
0Q0PFxfwZPSJnMlP++hNxmtmJJFFIGhz4+rIFvZOsc9AjQIg7vTfjVz61GIvGnnjzxluxZ4/9Z52
XjFqAu6mCatSmJJuhTcwfIWuJQPXiMDAGWjed3VN7JN5bgmRfGlI8y3tquobl7Fao/jCQW6mk9i7
VAua1SAPbfEifCH3Nz/p1SazRG3Ga5S5zUT3SylHK/V05JzkFgY9g8Zhfa5BT2RcQJ7On1rWZok4
pPCvbzWM03qa8i2QXKMGW6C5jVUeJeSht/WS2j3vI1UsYcqvN8LNgap9TLLS1dsPXfdNo9ZTRfIa
hFht3ouzwMheSZMeIXURahtwUzzv7CDj7FboldQa3VHPuPp2i28uM7vDRwL9mrr1JBfLSTWjthrH
KHyH0S273mxJ6mMF9QsXMJ9OplM5Y2mzX+d/FBISqukyByC1gRZU9yeyHwgLBSnnqJckSWpmKSB/
E5fdX2utJUkERz/DnIqqKonl/EW9RH9HEldpN6jOwf05z0PnpftAh9f3Mh3LqpWxPtezLItzHikS
YfUOCxza6MeLH4L0mBQxvPfVFTKoBCqhqXs5JXZlDtkLyLfYxai6BBYaQZj371fIcUvINDsrSUd+
lqqfsFRzojii9GpWM+pEeKHB8ieqPQk7AS5+Bt3+XwElAFmqXngw/ThLZqZOix/WfLNjtftR1jKg
l1jMiqmvyY0KLm/aG9bwgY8W8eAg20RYn0edDn0hTrmY2VHRCdzJzt3CGGwHF8kU2oCsg20UICz8
ngG2HCC+XCb4hwpdNzpOt4eNm7oscHm0TXGWbkhRcsyCw6zmb55PfPLNyIrwOqZ7gah8S1X2G5WM
SXvOe5+Xa1dCirPqT6G+Rpr1SH1S5BMVj/3zou4wqKCG8FXJjnTrq3v4dpsftroRl51gyoSxD1C4
3/MTblF3hLRfz3bhzvcZpTtM3RWDxeR6F1cVqh9Hp0oLVp4DGNP20doii2Iu6W+TiCEAKZnyb05Q
sIWh7lDkVdnBxyRYvQkeQCmZCUztDC0sItu10IAQYu416MVBmgECcZVMWjy+uHf+PUFW8+zA2oM1
9nQKTudtumnlEwH/IsmphywI2jcItFoGyG+XJFFpCc+PwZmL4KGh9U4MMsYi/HdJOOgr56ykMm7S
EytMsww6rwVKPgnEeioDflgOu9Fmig+sDSpTPeyPaJzCsvgvUWwEJIhcy4a/aCzG4h8QNzCUV5nv
Decq8arF5+j5kqho7Y2Pv7U0e1jaudv49YfPzCKO0740MnPD2i+9Pz1AMcAUB3t/xbA642zbL7IP
ZMaVbG7X8Gal6V9nELCSYMeP6P1i9U3q432uBk8269Gvzobdc4YoSIrT9+fQGUFLGsSPTTgqR0v5
k7rZTEOvTxR4gvUKVNPw7CiRqHQLCs+oEN9fYJem7f8/vazS/y3eAxhw41054KKQ2Vr+ZDF5anh3
phO5tmaSHW9TcBYdsQ9QDr8Z5no1RHG3mtYlF4e0Bf2ZaSnqnqEbCu8SUS3+6kZoXWM6dZvcRTPL
ngQm7pcTv3d+KpYaI1XPzvJwHOOxvDDYkurC4lwz5fR9OAd1fIpBetdZ8hEf96BJtg8QsITf5ZZ9
GfWtJ1tYchu4Z8bh1+F6s8+tc7ik8lBh8vH3sFfunbOYdAFvisDxugs8SGLovoc1+w6qqjSgzeHZ
Y4xTPVnqXLwcTBm30RWJiFl5vnfuE1z1LHARcXiT5ziteWbfddGEiJLulwTYTPEQOijH1kME6T3T
NW8ELxEjSPeJD4Wy8TJS+Qy4t4KU+HtF+r0SK6RkTqOTLsNE2hZaetdSoVPxc1dIuk9xLHUK4wyO
EkhzeSzcULsJ2kiJIOJkdKc7L1erZ9otslFpZr5YWOIGD5NkAJo0JCkdYd2jPEMT2x3OfjJLqFR9
TA9XQYPqpQ/CgQYEApnjVIk0ldVqyfYT5bJiuZQj3LyZOPOI6ERAOl59nb4FA3MzJaFeG98Nq6fR
EUUaqVQKZJC6IyKtBW5Emcb8aL7Zc9VTB/alkLCETw0B8h+VobzIi1Fq/AmFjCZ2LUahQBCeDNB6
pcUSER9IUYN4DY6Gvvq2U/KxCe9nRjmWoa4yON/1UpnA3SRYSp1hnpNRg58ElhZFiG1HffqIWmuw
a+H43N/dhUiFI583jsqyUkcn7XFQmkYpZcdQ0wqmg+VGwnyXLQILu7bVoYLHvq2y480IYvJSrPC8
4kvd8fCBTRXp7riHu7f67bjatEzm/ymrHTbyg2DRocf9l/64TdcT2ziGHFTPD/y27nvNoVKQzJEf
L6a5tRUwhCkjaNzUZYk/pleyx+ERY6nYWINYmTN/g4RIDQvSJX9h4pBnGoXHTMEJ7u8/cy9FdeIm
9Uu2Y8X37BpfL9BuVRHaN6H6JFF+Yl4TsMhzBx0IkEy6bJPkJS+WcGh58AsXKGogBPwVb43hiKzj
mRUu64dKeiQ2vla+gcucfN42MOyGl3PFeg==
`protect end_protected
