`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
NhlszBO37Lx31XDtnW37Wk/PBn+mECvFhJpg0tugiAesVYCSW2Esm9mpXlpyU9WF/YwF6sdp3XRl
0WHLQDk2TZ9K/Q6tZVflSBqBldz5rbq/NKulRandHhOj9kJJksMMIzjNu+Yh6ejgS2mp4FPVjGjY
voP6xN4dF/GvHaIf3QUDolkALAMKgrDNmVEXEKAyLM3J6B5Lp9cN4f/uAy7AhhXQgAthYG10WuIv
IEPpa25Xw4Uvsfaa8WUZpG+8fFM0+WtrdwawzA66jOcqFKd3gtqMxdeYbC2VVealLJR82ajqsXgH
jqjYwZ619Dg4gKKd4E7muR0pY0uh55EW5KkBpw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="tYa5qn0viUzLWVbU6QdInF+t85yc4twbUYqpuZJGzb4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6512)
`protect data_block
kiv9PFI+O8O3H0GKZpytUrpXqZOFnLnb1wL5i+9+dM+mQAsX1QufktIs36wRs0h1prG6Xt9ujB5F
g91e6nInH0Cg95aj+DfrQG99Jq6TX6apA9Q72t9rgUnEUs+1ew2qrT9BqXhc+u14uwQjNhG5IJ7/
jMuA67qRomPT8lGJn5cYpASADM5fxtzI4dVKm403gO+Rqxv9adq0ijcLaDFP3m+0MrpgbMeWVhB8
X6VR1W2N17H/R2Mj2W4LI5lBRaegUK3iPGseskEQRT+pS+BdyQYs4QwKPfZF3GkEvNWN1gFj/bfP
GqUSKg2vIAswYzt/HPrKhGLgoktgb5treMm++fG67UDlnEsNCGKL49ueUsNfq+bvyQNz8MHZGnY2
FCYrgTGBCiiuA6lG+yZhDrYT0LYyy/l1dC23WILR5Q2L3fIxlclossXWfiiB8XDOCpTjmAT56zkQ
INDUMFU7qKOX9ryAsVAPqeKEZsmpvdsk+E/cRslhNJCpyYV/D1sKzcT1CDGp3ajCKV+nrDUXnedC
Fy0n1Ymv//mnB9ycNaeGpJXGlT8I8lh87W2U8R0nJYX4JcKQhgejDG0bDoEjhD7WOLDdo1YyFoFx
2/dQlb32smh5s+dIzAyejY68zi8RNqWrP51PbA8ZbKVOJgxNNd9EboZOZi/kHiO/xPz8KPAEb4Ji
flAOKwKF8OdVzWmCMxIkvJJX0up76CvTltaRCDVkhDo4Q+rPAUYPE4jCDM7D97S2AsL7gyC8FKyJ
QhZ7gz2XwCQa1f5oChANmaAyKCBvx7J319RVtQX2PxntZ/Q6K3/Q56C7g8Q3QKMD2KU6PRX24/xA
XlQRg7I+j264lCsYz6lKgOBU8NSeN+byn/3aZ8sJNCmvqjMp9Xkgq3h+79/QdJWThBtlZFUASIIs
0kzAhSxsI+Efy/VzsFeeczbuGGYDcftzl/PPKWmyh8lNZfd7/ZNccM4+arJ56FEk92DBM+zAGZf9
xMQ78Sc8nLg5CF7P0THdnMj4ynAMZzQQxYyKpDcmCIzS4mXLuomjX+U0q7kkWSxYYG8ICE16gECp
+aY1vAW7spM0Fpn7Aipll3CSBJdikeaVL5cuCNhgEkJy1+sPK3/U059qlcTXI5yAg7HF1hHw8AZn
JcsFhbNUYmVhWPTtsG24MnvBUT8kF3QnLQJanRwY0szZdL+afE9vVM1ZqgByk+TpYd2ipzeiGCsz
li0RuoE3PBLgLq9LFAkg5aC4SW+XBVeGLV6pkDm40BsSY+YaqojmlvS2BB+LAJZJ/0Jo3ZgRhPWn
mzqcdbu1std6VKk82bKyVJZyLJ9FvAZ1FnyFIYIfE4/ZHovNe9r2LewGasFukQzExrnUOIEKcW9F
bNXY6MIHr6+is5VUxtt6B/7PDLge6TlENKtYfAlLMRY+4k3Mymy8X93ORmRIqQwojraEjGs3oas7
r1yv42KoUkVqdEI/FnDtoqSZdJDJj0if8FYwYXEoGElAb4u1GcIZPpUOESdBgcCX1w0BzGSJ9qCB
M+nD/lfPebVawWAcCNAx2VUQSUQWGBGUeNviC6U9SSmE1uAbUaP3Dn5WGFw/DmGU61SISEr1sWay
fNWmxuYsJdgJP5UKegUJfhZFfNh9iB66bZMTZIbdNo45lyGXi0wHtg8u4P7eHIvAsDDvoBfSQrsl
F3Ujt3gjIgoy56fMkeXoUW7AVT5Enz8QYzGc+ZD1zz9orVZPJXHD01OyHu1yGkm+qDB2KusLJkNw
YjUprxJCASDePm8RPtRj6/TvXZQWaabPoTaX1OmAtgRTpiBTbdMi0NkVu/3JJ58X1KT/1OEPsd6x
3eZCJs2SJ99wfDMBLlpHkARGHqEiPBdgBykx5pQseZr+hmbmr5zrExcUZ0doe6o9DKmF2Ojxiid/
AIZGEZCkFFH1JzKsls2PTlixDDn4WC+RRg0xciYS8P90iyq4baJJVf2OH8FxzPS+9LxdUQH1mwOZ
pfjEujolRNjFJNVg5gJtN/sAMgKsBgdJvH3nr8178ek+eMMOk+zkgVDeRgNPSy8hATmQNktINw3q
NkXeifYWiL2HShx8HF2HvwpyxI+IC8c7HRy/BK/6nMy2JdA/LC2KQP3dhgWGI2Ci6geSOehMZ/xz
bsQv53Jg89oLzpnU55QsIJVkKNMIsCiEd8zl1ILldRLcJqdzCpBJqQmfs0JjUaxyPTKayXzHBLcz
jbfrZPpRHH996jyMIBgqPriJcBO3krCglZHZcf4xqQR8TMLCkdqQRdAZTB4hp5RiC+08TAXPI8jm
5nTbM0Ojq7qVTSL2W+8tq8RzOMYE0oWVIXktbQKAev3GnqVG4+54kbXwHrNL7Cl/Z5EtmxjjteJN
aoCZ0DgF07RDXEH7HZxq9iHakxXmrK7dwh2DIdxXMqMXKkCqfAoMkdJLb9J2jtLasCrOsVGavy3J
LyJQOECuHzEw7hfc7QTanGcCehsHBLY3G56xeRuYf/DV/ebNten/fs8QVVWpPNn0EKxQvfTF2kmb
3PXWOh7JNbOBXjrpD71EHjmRy3N4MIK2g1Ilx8dE3uWETPgtZrGMuSdMtsYJf77MfR0Pdpixdq9R
j6EkCykqw1Rs7UXyjfVBPX3djZTEu7rOO4C3WKXipFtCV1dnYgYVVuKeEDmWiyASrQreiAY8CB4J
GuTfBNUGtL+g+gxNOBPx6BYTwp5bZQrYvh/Ul5DevG3tAMhP23mJV3qgztblxiclhm86ssUwEfTX
yIP3WWuPCukPBGUiNnQSgoFQFej+WK7bfKN+0sCNrUDqLuO5fLJs2YmYQUnqtdxkgGJFxim/oiP9
vNyCvterXQ2vZ9F4Xi0+FnFKcZzaoREAmhzYeFCNRY1wYOhji8ZBt0I5p031PTjcGCHO38hLNeA3
UhgKwyNMrxHEMx4ZzKIJ6t6asv/+oKtlrkbEfWUi/SNTZG1gIcbWEXuu76oIndCrCPb/8CrsDGav
PNKEc13uAu+v9GeDBbmGIZTK82k3EvS4NNTCvGMzvpZy5elorCR4FbVt2SXdSQUZ4nW/K4VVbhaa
RkDm85wVL5Ysp2p0T4u3DTrxy+NvjHFH3ajvrOjX7kJgsF+EVX/TB0tj4aPGyoCAzmt8M1dqTgl0
P0Vi3M8PSOD/CcYdA4kzkTWGlaRExPaZSm9sCLknvDgJl5ETYzZnFUq5IpCpYeJKVQ65afSXvssN
T9D2k7Q6Nwx/1kmUAcV9d3gmt6lo8j4MTpE37//T3go3CW1JFmHVxuCgYMOWtyQ9WIelakmLmWoA
J5UVKBX6+Xi0R56ZyyyPHV+Eks/C9kGY5NGbZzyGM/EZ8L6FQBHymB0R9TbCL9XONQ/AGIH8UQg+
ScIb1/02SrGkP12r8VPkVnwToiyG0H9jOs7VQru5Hb7BJaO7N1oB5p0Lk3EmAd8Ge2FqANLcTkzQ
7g9vsviJE7ndiEJW5D4nbpinLXPs92/ZzGP/vLClxpb997Bi8yqJ1l7ASuuRkCH1vDg5OiXXrulE
Y0kVkekBBJu9d77f81IzJPIxtBSlRrapDh2kdlYfqqKrdWtxULGRx4E2rtezo3HOtuCd5a6LRtwH
uWpRP/JcFmUhDqvFXL0lEeqCSwK7haRFNR0NQFtzfIatxlOKRs85icU/gobt02B/T3NII+vdI83c
x09g0zbRjY72crZT4dhTZTHp2c4uZHcCUcFDi2xHFgIKlBK4+ubIOCOkSLbjOov8/BGRa/n+WpeQ
pUvVA1OKEzIlkY2n9XlO4oHOGD1Wvidza4oMGQN/MdO06dJfqhErmoOSZo2X/TckbB3AOdsYy3oT
hByHsB+t4Fa38hDbg8POnXydmu2rAgNzTxxGCF/k8oL33SZf0lMx0/R+HbAeUeBW6h4uXfrdBwsQ
sjgXuUJ3Vb2J7znhK2NbjfkySFiq4/NIvgRzbYQr3KKfvAtDgGZ7wW4ChVyDaCOITVZdlN+mYItA
AEOHvVJuiNAC8BTOJmYa0wFIwdIDeuQJFIjP4RyyDKia6qLvvF1w2rMSXoDMiRM9Rba3bMAMeE4M
MZ9VE73bsbKTMePRiu95KqEqxdG5AH5UyBCJ+CDikQy8jGxDHALcjmh+7966HgKRtaI1rdsVG4dJ
opHYNceU1JakNNiDyrOX7iUBk39sG+uYkgpfQXvs12bQ/Z3+RinEz7ZN2BBJEUq2/onyQw6gpZ6U
RA9a4YF8zkFekx4d55/H7g7gaqX8ZyQMjgZC9Up24rcYcF/pIUr5HJCaLIQn5Jo5MZjVcaWfEfkx
W1l/Gpz8Yk6aDxUXEgbJgUA63DiQ8D0RuEZTrRoyAX7WuSLLqZ4I1XbEsrhycLMJVneLIMuuQel8
Nw7tdNJRpka0Kd6LPxxDmJWHj/QWwYQeGMLnM3NmqYGAPeVMc9bfIMZDJ2onYQKEJbQfQZNY49k2
toYVJJaN7Fegpo5ssE0hPAbdev9cUs3bmgMHgMStZZhOG3yEQP7YIjnuTKwnBXYUI9Gf7CZ4M0GR
BJedh2kP2lSAqJ2TGWYPexD3Iv3xkw6BmgoLAYCU7DRijZo+TA723KwYAh4lG9RPcTwctwLRtdzb
Jgk2T6a99nFbcv2OAShKZoNFn3FpK+bm99WbBlBdAqOu6MbTlP5DDroegzoLfWFm5hTrpWNK2UMP
BpnXMgyT3zNJ50ZdUa6kzjiETF8Ge18nJ/gChWW1GpDK/xvOs2+Zm7yxuC5KKn3iE48Ic1CYkchs
a7BZRQ/oY3H4VwQKCax/eb2GRuM8QQw8phvsGUN0hIfDQQAScP13jOiJoY09SdTY4BE7gWoURt5N
YXiUiN9hYuhFMVL+Z+YtoU4jE2LkbexWLBtdzJGRbcBRJ1mD+ebw2usWHnC00qw+bN4F1+JqrMZU
QUZJn28EwUgBLYx25R/c42fxhDwzgmiiO9ZBn7uLJDZPEEZmngnAIlpC+nrVJSnOMtY8tm4mqjix
DhXrSRnEMbbfTcY1I1JBk7s+688Gq6ti6cTX9MP0GoAOEi84OxirSJ0yPwcXY5Nh6neQpEbiDphu
Snj40gjn7TUxIojwO0bISQlMVmC9ej5M74q7Op1Z+z43oHr0hedNHVufyPK3JMwDKfzqEUOz34o/
4XEBV2BjSulYLcgMmd9JH3/QpcrPK6n4AMqKFRM+r5YTI0LLhFtETpgjuca+RWWZ9Fa10NsDaUZ+
jZsZwHwy3op7uD0I/C+xZiFxG6rDfxpfn62EHOOuJcv/GOymMBlM7AJq4yrl+Ko43xtkjpgvoqAT
Qm5SYXivXqugJVenwVScQK0t/e4OY7OaXTxQn5w0UuHzGeGo3390XOWWe7I/0B0Gw9lt0rpXaz3C
m/XeW4TDmMukf6thCr2/22ZYMQFKroIoZxXV/EPKWlJsoQ8+9sh2Qg7RWx15n1ljAh9BjPmYjAsO
0YyuPYX0FLJ8tk41SfM4RpBL4Q4moeux/J+HbsEgPbz4A4sROPR5tQ+6E10TkblRbN400kwomDQn
4R/HToxOo2XE7fMaWz7RIdOn6s3IH8jX6RE2mz4nnGWpyG/xqqTKhcUpWqs5o2J/f5w3VwhU+Xps
FA/eXCcrUhkgchaNwkZKW4L36Q8CAAmZSxzrtk/r0i5HdsQ2bjjoddZnMTt2+KQeGGahri01spr2
kEQo8OO7YREMn45MzP29XKceh3ERDUHAFH9/DnXGxFg01mWrk5AGP0X4NV/mJEI5BRfD8QBRk/2h
96VZdmlhUOUxk3FEI07OScbzNmZ2Ziniu2ZnOlZJGUV15g2WsdtPil9d5VyiAaf26CG7KUoOiJJv
Ii2SZDpfigb3CJFdx7dLUkd4msxHbUKirXyfWQzbEJqh+vMms+TaXi8y8dpvhwJLTTDOeikL7tuN
6P+hmOcvtHm8h89E3EjoWUK59aAqjnpW96sBJdYGOPIjzaABVqlwRiIobLmrTvJC4TKwxdoamoOk
+EFs14GQJ+5FKbmPs4gBXEZrdD0iLNdQF97gg9Cil6OxWfIHW+YrJTkooYr4KtoPODNYQYjaVMYm
FHXOylQA8pdwF2AzdDLA2YFz2uF+OxEZzlbP4nNdS3pExVC0Q1DdCFxI8OBU8TRQ9igmyOCkjXYu
moSvpsrTjTWMkZyBvf5WaPvOzW1e06CcrHrRkBWwrT0+Ds+6AT7WKV15+IM7Vppf8CgxZZhJxizj
fo30hWhFXtXnLQARcOAVlsZfTNSUNZG99SJiGf96Nu3kVbyDh3zfA2ZN9MOeUewsQU0q4tu7dMEc
QmRK0v8CpG6DXODbspnDs2P2ZQV/8twN3W5BvPVzjXzvEFda3etYhIAE2AHkLpV5LqEZ8hDtU0gZ
4f1aSZJ9B20/vTuc1yEmRTSahYQSDxT14pvjq/nRBJsiIxV2IBtrEj2kzv0xiFSJgud12Q2d/V5M
ZO03E7pcCLhszWphVhwkmwV/rlIH4DIW98JU/CSo7AyfpzGsyyJwNjwfWC6MfGTcOLf0IyTWFuAJ
QyXqCf1DhSgrM5GFSE/GoP1zqi+q3KPfaSYUfA8RNBRfTcSkB/XjR8I1ZcrKaZpS1NO0aLHreyrE
cecxG5O8b/QwlapXH8ZxZQQeg2W01DJLtSdt4WEjIxnTgrmNSHam5LD9uZ+8TJjvHMFtzb6xePKI
dT06vjNQiqhhF4gJof69jHAOMGGIHFQ19ly5iimnWBEHeSLwHc7Wum+B8OlID47gqukBT/0Sae4e
Qc89+c9LuBMXHJTHmab63TJhIIr4qmzf/Cw6WWXmtI+z4w78gHR0HcNwclHhr3Ap3VlQdTxeNLot
kWw+EenEhio0N1uX5BY+Im1D15Mp2XRreF0PetQSfIhJjbBUTM2dQTT7mb8nz3wgZsIYRNZkS2b4
82n63d7EBk2MnlrIGTbLQaTDgoYhFPCb80JQNfMSOoxq+K24AAPXOpYxdX6XFanq/pRvS8cAPlL2
6zv9vkYj22yIxc4WwDEPlvSLMzND1I1399yf+8KCqZ1VVZ6sgNz3X9VazwEFdxQB9aa3GaG/roR3
RTO6BVwv35LymcEeK1BRH7/Ux7lfjmh7t49GR/za8YL2nyn0kaEEeyhy6xq+ASnPRNGxo9YNERUd
uh3e/3hBbOOXI9nUvgTeeBTL5GhnsE2rnwuUb3bLzwBAa72Uof1sUIOyKL0ZbKOwjZM/1k8oXyyh
fCZNHLvF0xVMWAcLaFx1oKsyhx43DpQDBcUt1tSO2wsKBu6ZeztlS/78ArIX0wLYaobQkihNmVXG
5mtRapwDpJaZWMgOOrHAoNDWSRJcTM3wUFSnh4+Rakmjq6PSaLoP3cjiFCyB7o1l3YRAn5twSM9z
REHanFiTEUwKdnDHFrJ0DenTRNObAyyYrJF1zVJqofw4UEVBr1hEV0N+y00W5k8/U0tNlnSQz0bf
3/a124TwWwJwK2Q6+cFNGKVCkI1Px3BI28c8nNY2jEAOyQyKt3cixBQx3E7H21WkaMQAjMTOBkUx
h9zmWN1orho0GE3NE/yAwBH8AHQGRotOCo/VhHxOd2cyImPrh4LlrOJ0JW+7DB14p/xqlMFdRAyU
vBLmTOu/wkWuhRYHYihbbDx/t4FAajp1lds9/aRWPvD7sT4yyXmRhX4j1QNiabsYuVfGtWTPIz2/
txM8D2HMNYXs3zt8hu0LH+SW8U40raaxszbkUHsjuWLHx7HI5/dDq6+sM8zgfya4TvCpo/vNCLj/
kNtWTDheXtghlmjcAeBGh9YjuRoBMdKXy9UOwmED3Hk2eiPY9TZffmpQLU/AYw0llGObrz1lTcP8
z2K99LEseL8f8WgPSlR71KIk/R9rQn5dlF44C2gPdexJ0Baz7P96qQbNQlgLGKEWq46Y96nVsB9a
F3UaUAfJyIgDwyW3J5q0jtVawq9YibQQp5F2Y+jhPavd+GfGXPfU9pgORKKtrEyF2ny4fJUpyuG3
+oI2J0YuUjjnc0r+2k+uiazF4/Qu63+XQQF55bHAedO2AlmFF5WgSP179nBrwhkoq/BU3liIeCFp
54ZAH/29SS2mTqrij9QTZtThqE8olBPSa6hVM6iyEbMnqj2SNkEgcfiFkpHHlnNUAFR3rachpsLN
RMHlDEfRgoswL/dIb6HmiUiBBEUp5J7t2Cp0f/HCrWYW7Ducq2old5j+TrcL628iyHtUFfaMxZ0z
6UYLfY/iwCOYg9/qcGHwRb0+em5hiL3NKcdnbTw/Sa8tYIkeO25oE2UAtAI/dx1GAvsna5H7pU/0
6vYDATxICzYEoFELpA4Kzxigq/5G42A7s7+MH/IaAyypBPRBNIr2Igdo/3fn9ku7BP5svlBi14C2
z2SrIsdsV0tBhPjOEn4UfnUiMa8dsC1CmiyjfiihDfp2vEf07GEcRqM3sluhU81vm6lrKVw1jJJ8
ywEQ4uIYjVYoLXti/U6jhkl3jGaLsjApY7SpWDHj+8wgDfF7oPWXkjMOCvH3yZS44mUgjtgjmc47
GSBrFPGY178JkZ9xExD1Fqq3glDPcypCBjm8jYkY+gguvSMTomnlg/J3sW8Kl0UxSnzipXh5eyFu
sZiEl3ev3pnmELsV6U6fO2Vtji9J9+xi0O+yVeiCpuP+el/gyUqsBGxJ/RwvUeFvwbwAdRR6+5nM
1sjwlQ4ImaleSB7SSQi4cLodoMDBOXWMpsx1JXhXAW3RdiPZac8MifkqCBAFUFQ+H9PMq047NVri
uDKt+i6snwEBTvG9QC0=
`protect end_protected
