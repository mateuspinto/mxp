`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
G2zerGrq2lk5nkKYVaHT+CW2mYbQym1e6DELve3LLiO6CjHRbPTs1g3LCdv9uyKHP2g50ntUpkCZ
sFEE4dgRQy1BmGJl4jTsQreAWvw2tvUmKgLGhCFJUrwXq3TpVI9+JWZIMa3ooLA+VTd14rmO1AZx
uzQk3OYFr3zdqrOHqkYmogb/VfdXGb1HszYbkC/2+CzjaA67Mkwvg08niXyXBhQvRsokArhBMpqx
mFwfg4Ghv2Xgnsh6mGszbVuDEkIFtzpsyzoZCCQssP3OYMEKMGANnqGmEIHOMcEKoLSithm/nWo3
U4i/f+Xe5wzd9HKNSWGW/Bzt+6h/kAkMBKMJ5A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="1pDv70dnhTE/srBFJHsYLg9GLtY9p1WW7VqWRGXy1pI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5488)
`protect data_block
gfqlwo4MShV4MZQ7q+iG5QyU5rFy6ZvK9Eau0zUxO8OKFGcB653h7IOkgbmX6793uza+AbxJDiop
q/HWZpb/aF/u8ZISz01ugRL2qV9q+y9kRAQHT8t21FzT5XWpONskUQjeaS2dQKKOroTHD3GCanUf
bNRfmwyqqy/B8jICGyRDiUqzUd1gNHPNllnW38XZVEdBg+spjoR2CVeKnNY7Ge0U0QzMIixRs6+F
p8c3mIh+dygOphwP6HqzkeNbihmnoWGhYXOhrXTXgerHa13i6Obv7tIhPfdIH70huWPsO9OrPCXF
fXR9wD9UOnH7YtMYWFPkKAOQX71rvvw+Pk+QSFlLMThVH1iIF98wnbKsm0Hx15ef5u79a1/Vw5Mi
GYoqJPpDUVQr0/RHCXOVrHuXYpVEpZMdhTTVPRvqyq9NkDuoKTS5COKJoaVRgTCdyNTFWfCZ5mxR
RRmllH/mEG9WS5ComAFPt7X6xQRAXKI6/InDzl5/+m6fjLWQG//AVS3DbLrorPkXr6VeimQVipme
fUwSixnIWbFTPbsrsy/2IbnA/7EmJp9cdNDBCyx5Gynpf+eRRrBqN4QEPopiGaU4lSZTbZtwhKpC
dyBeWUW9aBUnEUzWTPkeKXuoPqzE3MQlzC5ytOzTj3CNV/XfG9mBGQI37GSr8t7MZkRmenY8gSDQ
zSkMTLb/6WfN3oIWN2zE86pWFU9QfUNNb2ki3O4Xk+MDyLmC10+sjHGEB178p0kO3JE63gMBgTB+
FOrHEJkj4ie8f6fKQy3+rAnq6JGJ6bCP9WTtalVa6FqqTmI6Z59pJzcoxKwiriSqWjnybUd57to2
LyCpDNad/JxXBHPJF61l359GnXhfz7ipvxnOg+ZHZViA2lDnBeX1ERK0emqUBU9i+u532zlk18Wf
HJcxE4hBrMpt5IG40QltG5ffNICWD0tDAFTzMiKbgNlbVBCNeXgfRUIvkjV681uwJlzO+Gy1fyLS
ADu50yN/hgJU42+3lm196zfBUpUQKD2B5ApytEMG+N2aBGxGX9ZAdP030UbT8DQfbZxcPlC6ZeBm
2UkJ/BVQlFUQ2uGUEVuDDoEg7Q5JFObzOMFFH1K6PwXenz3Wr1oOVeGFUhfoixwCFM7K9ytpnU6T
rT6R3FESHEV0UYF1IvBYl5glWoTguZXGj5DU2PF5osry2eaV6ciEmvl/E0K847MYQzLmjmD4Hlvp
flX+zwS1NcfOfFEa0BlLWCxN+IUCIYb+q7gcAuYO5Nty8hkUpYhUrj0nkBobcVwXJcIpoWqPr9Bi
ZlnG+OCld5oErTftmPbYTFbetAla53FTx9btdsTkAImlhu3xAisMinpTb2OxuxO3jpgEmM822QoM
MH1k2c82YHj5ei8vFhyxznDWkkEURWhfpbNbsmmD/vGnAWYHHbJjiyIp039z6ykSYbplQRGd+iYF
CUwVq09U7NluQb10TGaSWzJdL4Qb+B8aIbfvnlOL3t3D7NQsv1Nf9XqgTlgNoAehf1uzGUly9ew7
GLOXMMAUpLW6o/axWPW5TQ6dx93M+9ZhQKSVCHkQl2YP/zWevkOAN2KoCAPq5PCVb7VO+hpUVd0k
/3rgdh2LHWbP1PvMMjfNX54+TRPBk7dpbTG+aNR6pI7osfze+cCXTfvJvUxnwjgZaORGz5XKmsFL
Djrujq9nR2ssNNThDowyS3QJAYG+VhOELJh2GxnlcK9EZXlI0XxdXyIYL1mhiVbh3LOdsG+gvhd7
EbSoDx+xoHcFgG+G7Tpynr0gbw2proFZRs6A7LeuU/uz/4rLMYdNFsC/ZRw6Jy6JgQDYZ7gGbF8n
T7I1Gix/UXyqTFVA0iWTxMRWesgv/cuBQlIhAbmpWNH51TUF4a1D8zc2ykUit5NbYS5UUAGo5gF8
lt9p0qN11IeQsGjY0NNB/2TH87dbMsktIbKZVRVbzxB/K4RKMJc25poFva9DW0IrLGJ2XSCiZ772
vWMvNaqIlw1vtBHXunkNu/NDBCXAqnqHEQk01TmKY9IF+wmzsUrDeGmQULsIgZ6X+pOl57yKlJl8
gJKQawxUeVpGam815p/0z1dmBPcUqWJV/GyeTQW325dmFujDHyGoirLk3C4+p+Rp/E7v9eiQ7v3a
K9FSKO15bpyDEuGmfyday7m5SorigPkwBpGf6L5ueQHnxiBdgsxuiO9GzHasvD0gU7qLbB6thr/n
WDS0URvlQd6/+XLGjH5nbZ2/M0QGfGFXSc2pArh4D71FNYBDP/HaDrkdyZG5rQjr0xjp7ArsFHuv
krQ9SJiP61Mt7kxsRAIiSiyOX8zf4+JukwarNrzUP3ms6Uk5fGp5RBPRaBaTCIYDhzDdI/Mf7fbL
k9kHYSUUB09VEDLKFl/gNmyG/U78lbd6i3JBK+hSdlUPgcLNgleSG5djWPiD6VlSqhWZdaRr0Eo+
89dEPbC7TCtym0MuSgJyE/cPpYvVTFbkSYeWbAf2djNIo4+t9jUG6zmh2vXL9Q9SkqHGSp2+H6Kg
PmGSiE+7g1aKLo8z7LoMogTnkIQDGTIaSD7GCUHCP/+4hSVJDkEMZinvQNkq4ito4bpIKbKSlkWf
KLFgp/1eOQ6YfLwsEHsCLhkXynj33a68gf2CY7c+6Mq3RBAjQbkahJyD98/9kt6cfuCSkxngJLwH
guvf4crnK7uOYomzNaOqTzeL8VyzZeQw8VPAaAUh5g8ujWr4R+BqsFTqVbVStqZmRgzTbq1QRoVi
OZD9rXfgmwXH7U48F7fCLobB+VRhYnOf7duEqtuV30n4Ti1+SetHsiNVosD1Bx+v5Be/hSoGk4mN
oCxJNlHsbUIAM7O/o/Sd0dMQtECETEUaLOv+4YJsVTQWOZgxD3bczCegeTkqC9I9ojan1xexHKS7
03TwlpTEKytDXT+IqNlMt7AC0bLkcYP69NfpwxRrWkm0vhDK7tdD7IGYUMnMepumMOmbTzr34wLL
Thj8Zimygo8VK9FLnQBNOO51z0fjYjuMD/UDqDXeTqwapk6BIOdDFmjG6E8YZ7Fb7w0xwEMTjtxE
suy81kYP2Kp0isFim+ZvEH0HK6xe/51UfViF56g7STG/zRq6acLIZFgA4WwDVvJSJQ01XpAZ5N0v
gYRmUE1oBEyphP6C1RazrpF3VeQD3fpc4O5oVaskOsg3T5k61RpBERILY02xSIjb/0SWRc6OSnqd
Xgx5x5nM3Gqh8DFuf47LqW71sKRZzKYWvMDNVU1GyZQfF1+vvOb4xnMgoFIp1oOyokqa7EQFtDeD
IRohWEQeDuJaUHgibBs+zZjbml/tMvHYwfGz48vfm5BbESKC9wre5jkKtIzhO/q+NdF7sgH5woI8
OMDAe6XwquyCSTlg7YErUabOY3Fv6aZ81qDQtG2KBwBrBUT+CHmPHcrVqqz0oP1IKcYDnDkxafcL
qcZf7A/Wp2R2oZDobc68WGFmuN2eZ6vWunbb064c5xEkIc51YsfsI0xN8JTOTdRgEaP9HPifEaKN
OJ568V7t4UY+XTE8oG09ftkwDemVrkII+FSoiJojomwsZrTYUSlFSzCfLhQPEVyyWVzW07sQmA/R
7jatWW3HefKXzPuaS8uTe/aQvdh0cIZlQTTKGHNFK6mqv4oOTjWd5y8rvaMMREVNDQG8ko3K/tb7
WuyxJQ5gjVM/yeSV4WqnWdavFcSdIbexunDoDUBdlDmB85J/BPdMnXyWtY0in8n71XDg05Cb7FNb
C1NEaKCDfW80e+BhAC5dVaEn1QnHYyi8RtpRQE6XfDwLMZIHiMc/9yugNykZFknFRPnRb1SVo/P1
U979NUcSLKVG8PuprBbst426uLRl8JefEe8kFZaNUQ/yusAWJ0zsSEbNoYMZo4T5b+dvXlBUejfO
C7a+GGpWnNcybrNRC08KHr6zyQTC6GJk7pxt/0FwUY4QR1I2rlGSDySupyekoyDU2oHfxnbNYJsa
fUM50t+MQ9WitiRA13cgmOM5vYXjjZt0rhoY7LA/Xin/IBCOOwGOm5M6sBxJyKVfw1rFUZ1OV/Mb
2mKBxHBD8Rf9d5Hnm2DywJmyK+qUlPNgw/yF69W5lVNzDdo2NxDuO3Mtn8Z9JBSKl+7Z23okg90H
7HHrieah1dAG0YqxmB1Al0qTopm22jEbJ7lM3hJW2DJaKzY05ra3S7BySF5hooXRtuG/ewM6c0+c
5Chd6/GeB3bSoLPGFZE6rq/MQLxiJG4IOm7GKIweX+2AUEiCf02q9mnA2dl/EwGRzd1nmdwY9Nve
FW5ndPBwd+SQ4pGvkSqqmevux+HjbCT0ooH3maX7osi/EBA7PlE4/9IMMna5ajCEv+SSt3QeUuqo
N6sqjUx3Cet4SA+CbdL0rz2ZQyLZmfKUC3wsf0gH2uOPE1XiBFaGNTQA/2nk+pcbGa47pR86PqIt
rwp57nabOMn1MZXcYbb8VBCfg4Frn7kTZwM9QYXZgI/SUjyFKetZ4XKspSgcpA1BZQAdFfMz5SED
6JTlFzHU6mQlIIuHzzFTXbTWyt/wY2Aly+zd44K7X618pT3UnkdDzeYk6BV6ct9emMqLm1h/0/sh
/LUbt0XDqqciBOvRveWDp5qVuGZaS+4P+GuDLrXsG3g2tg5wHrHlR0kccW9nqBHbtOcsgTnUsAI/
NonAa6shHfVUyJyJWd6xeqbpR1/+ZgIVy0UCjfkdVCX37f9ZKnKbbKCHDcvpjUFAFW4EC3Con06q
tSqUbUk05DacZdZA3py3e87lhWdWG6ItVdtLOcgzmWLmvWf1jYuyXYh22ag0WYWrToSatSR3MlLS
hz4mjoBslmOpxe0J4R6hhot/VOtq7eApGBZqfDlA7ja1Gj7AKER9sFCJIbQwzDem2AeaZYC2DpJV
Anecp07Ak1l3uv3e7mMPYdwIn2h3fgUk7r9XN0xV+OB+yREPIR5Y8jv4G+3yi3mu/zUtfd0cSt9F
mMgwH84EuwCJvlBN/qvlbHK78lAgfNtfDWyOEMax21vTTN0dSakyyZ/dJRCa7QbhjJECQLsxpxgK
bwKlEQs+nDp0bhoXAfO3Cd9RwwnpY3lUzCIiZWfLGfIkEQqQ13DKo9gdLvAEGHBtpGN21AVMrf0w
X4mDTSIC1JOnn2EO0k/HS2dqzmpN9rr1tNvJwt1M2FXU/y/qWeQNDMM3nRiLWrgMhK8uKWMIZfh8
bR8PWwQZwfbNJU80N/R87AC5hQBXc2Vd0gx2YqZnFJ+n+b83fjk8Om+yDsFAJUOhDeEwuRaVhCJF
SpOl+/QKaKBfXFjM2djWSEKpZwUDACF+685MtJxaI0eHA0IGXqzE6MAZY3L0drT/Xml6g1BnUrta
XRU30gZP0/m4R7lSfIvDkxA6FsVz408+XzFSDf5cxo4tQ4UIANVIeGbNnUXLIpDS3pYS4I2s4IXS
zz2ZkjH9YpcRgMDnhwrwhCSHY1zhpRVqDYI+AGAtgRwpAabxJvcUHSSnmSPRjFDvKImdLRbIKS8S
TpSFU4c1DNEcU7iid5dQc6DY17nYwPrc4Vtj5coCo37YwDVKCMCmjmP6Vl9tckU8mUtkWAAIeqw3
PCxWHp61EP8+P7XlfkZcw0TweAwMyq2+GERNgDFoW+srsMqRgecA7md94/Cmcf/bIZXJQS1rUpux
Se++BTOVSeoI9MifxD8LnK9QUleUkTqhBnIgoWH82ZtaEpcyR6l3eGM9rFkqY/xTvSNPs63A89jK
nPx/32vJFr0tzncvgGUuwmXcxAIWhR06B4waCp1SLV7AvpGM9c2RO2RvitV/qo47rvkrqFT5LbyH
+d3l0CKNEUnGTTi4VtuMd5nb+FUamsjvTUk1C1ksrdO8hl/9Vd9hcd6MV2+fchQ65zoXLq4ECTIv
HvY65GOZfu2tdACplYoAYoDPcvJ2JGjSbQhTw1xADS4MDDl+2SxHwTqeuWMB0x8zQWciR0w+3/re
zBv8WeblwjsmsH+1IOJoc+wxzGAdl3qRA3E1529XRuJkgfAJgnbC/v0ZjlRIupc9N4lSEMxXI7/Z
mARH1YALUaqkGrlRqVMcsB1/2gu1c2gEyt1uT9ZSwmPd/OIPxu4xx3mRKJMJmqbVRtT98jpLqzKx
i2txW4fns8qBvdKKA36wZxi+Ty77Tzs5wQ6gIkqHheDBXHZA7y9p7jBIxyY7C07yTf0OWh7Htoqa
USwq6DX1FNHYo64XugipnqKBSUrLw/8xccAW6OqJMq2x67id1PnpmrFDU9X5741EP+3OcvCyRS2R
wPxiYUYB7MnK0FJAIeFCqAStpLBhmZyPaReZ2RKiEuv8HjPqLyrJ5zkyRrrmkd/bofwcklc309NN
BYugSoLtnP99js1DTYMsLG3P/F/5g7/GLASYkdAmHJJlaa1KDIRskHMCSDzlMMlUFknxKUsxdd3R
G/ZjMzpIIF9lq7OWmamhBi2AMcrJA6NUe3guVqhPdXCKcAdB1VArHbJOhW7ZiFb+qHBDsuZna9bZ
TdTVGHXoGwvuB7X0EXURbJNQcl9bQSpuAImqLS1SnL/mHm/sykPcYnZ/0seg/hhQ/39LfjF2g9Fe
jlqjoCLFoSeAjR8ticadebvv1ylcByXHx36F0FtVF9OpTphSc68T6jjmOtbsWwBJDH3vOSp+d1u7
zEgO3e+HBAgoxzINVTv0mHOLixCkAolQXOYrFCpToYjYPdiiVVh7XvtrtcXDDLyKnRSs7QAiUnqb
G9m3GiH2O2mYS3PCmYHZqYkip+ji/bCXgVgI/y2pE8hY0SYTZBbTLuBboCfcZyudWeG5lG+SHSyj
+VwIlwvqAyXc+R3O7zy+eqcKv/DQHBukGPm4yaxdLBeFjRP7zLBYWC6kdG6d/mv4KfnnJR9UVlzw
ZrX0au9TA7hBhJkUyYtr7m8VwwjSqb0g2enFzRzqWmB45TR7nsCQ0r3Zd5eFtyQKwnO+xDEXVK1l
5qZTZJZB65IxSrVDy5KgsAY+ncTx1lpznlZAcJXTT+2t6S+ry9gWO0Q2gd6iAZCQDbKA/RmcqyUj
hrM8v8SrTb12BfgWxJTrEBVy7gbtIiySTch7WY0aNTHRwL048gKLEzBSfbV0nVidnSzRB3xWUiol
9HxeZHIpVJgi7R5AG3NLC1OxQcI0K5+LMDkqcN/QXfk2Cp6vcIC6/CRhsRLWGKxeeGNOof4cBIwn
4zNQE5ZqRuCbJU1H5ro6i+WJF28tYhGTd5cjA9xMGTOlcmeEP8zKcnSdGx7y1TvBCx1atgALZk68
E2TvbAUkoV8Gt4Lrt1crr60k/WMhCnq3Ccbn1/3ir60njfPZOOYgjWbtZjWUzpk4ZtUTmx3TGzFg
qquZclOe+aiuJqkVIYoGmw==
`protect end_protected
