`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
D0bCefI+r4ZbOYquVx2BMxedpyn9LR+6dGrXyvqbdE/RkB5VvQH6cCnIdwOUgPakiRHwpfdmEcd5
KYEBagFiW7pcGMNcPSKFILP3YgSsRpFf9zQgvPZYHcQdvj+gMuGap/eQx0X96ViE+F3TgC8zORt0
ckV3347bMyMn47X9z3t2GYNeFIhA50XqC8e45qHGYx+KdK7c98mwRDfx8APyqQ7p3d3njgXYFubr
oGCiOpUcyPv0SHda1qxpniVcdWgsMdGqQLP3hlLszHMIpYyotJMiUhPU+s8xeofMKABVP+oQfuTO
ubvCiPFOeST2P5+G2X3BffxLpuevqLYwUSeKXg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="Srs3eAZN8U/+MXXJya/Uh1wiM+csPgI4BC/j+3xRjuc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 68736)
`protect data_block
lJ74Q2Guey+P8F85VXRTMfaEXkfzXzUYIT7nhHuyqImhnBIno6AgNUuGgbN2t6G6A+nLQgSK4SZ+
pVdaLelOmJ+YUIcwlQ78dQqgnUKcCpZfZIdkfb4XUYjvCiPxYgcqsEW10c5iFaLz+hGn2FZPlM7N
96kvfGNAj9Hds56A3eeSsuRrbchKzTezEyivfB4jASVnXsPZ4AXMLNPlqqzaYD6VceOiK1cl8SA6
ltH1V0Wq5aGUVIFaZlB6kFbYyCk3Ns6rmQxve4nqa5M9fw3J5tpv9OvVj05k+trSBnMEyW8eM1bc
0Mu1ktx4Tjf9L+Lhjy0Ezo3VYC43ANQypzMy4nERS6raW5RFZlZwS6IPzyFtJ+jIbWCu5Qku3aFg
cgOYNtn4WPzb1txBs3kLdhuHJvLj1u12Xa356pUiF2Mw5td+q4JMCmit5nNnkV7kbyEfuZHvrVt7
AKuO+tx8CVEuvXddqWPM4KvSn7NISXj/AcNTHLVNob0b3bydohJ8rUu548L0bE10mxZB5PahYBEL
yylDQAjy+QR9w6lXm4KUaGbEWqaceyFtusrM3nvclTXpEE0lXD8QXIKytdXW484ho2iSB49rjL4K
8PnG4fbrZy1uhSKCW19ASqWyykbO2l8YHhxNxqzLfLqxUI5Flxn/o/sBhC/kAp3n0DlmqVsFW2kv
qYmB3jLGUPxXfewE0jrpdBv1Zc9AU5Di13GpYczo9YkrE733Ub+KkaVFykhQ5widYFm/4JTOloUU
RxCgbAfzPer+mZIxC+kls9XhnjnIMb/osIx9meIzySJCT12cW2+z0F8NoKlkz0b/XBbnTi9k8MnQ
qif52KpJWsjGuC7yVI6B+EJJ64jZwU+GpKxv9l4TDrs3ZpE7oxqdgmrz5OtR/Wz4pyTa0QIZEv8U
7EPffVpOBYLmL9GEXwdtCVNZn10mRHdFswSAGIHBpe63/0bCFF7UpRgHi7X1AAszCxj2fY6d3CzI
NqMRgk80R33ZCjEIbrfburAaEQ0T0ZP7OYSHbfqds7EWMf7zDXfZVZwGvOBgnORe9T7GOQYS7ovx
D3BRBlg7L8xKSaTT3hoyi/XkSe5/QnzFY3pdbWcz/3HUUvX9l08Ihcrz4jwgQl9KQz1wWVlTsGlr
RXCIqoeVF5vvX+fDfVCo96ymlUW8gfBhSzI1mPv5N7OA2lzkBo18kPPI9yPFwDCVRtfj01ljdQfs
zlEyjGKUBRHpxP7CGMgb/awH0iY2ktb9gFSJc4RrnBVD72j9xoHzKOthyJNJWRhB3kpJN2iJMalA
actEqdCd4CcFsMymlvHhx121XM486gDCNkpaVut6/y9v2Re1wg5XuGrmVr/lLY1NU1HWLJhPxDj2
6zRDRpEKTbAjWQTXuwgjmYr0z2OSuVxke+U0ThDcH6mzNic96nWLWxCdkkqyWIk1G7Yi/KQeOELU
0e71C/WAjQJaF+3TNAeyZ1JXOKT8KyPksMgSrIMscRcGzoJnesaNDfYMchcyZFOWxYj50O51TNb/
uVfFI0WZbO9Jfqw4YnIKeKkrmUdLg6auPneWaROJgm+jQXSsQjD6yvFsjVVkj3APL8uykxrwe2b7
cMVvl+jEMSpRUSbY+mbZKjfV4eYE6yWf/2ZvWbvq2Ime6/XGvnpSaFSjHcNF/AeaRgJ1/tidkIPa
3uZhknrpvl/oguHJbFr8l1a+uFm1XYLwH3JJFnoa8BRBAr2ZkSO74XF0zT7tMny278Bgu7x9vpDb
qI2G36KezM4T7qSVA1wZY0Lpjmb2Nht1MQMQhdaOvT+jYFCUHVb7djzJagub0+s/w46alqSgHqsF
xiWgNCwfZUh+nKc/C2D3nYGwRMbncm/nHAiVWj3IibX6JQlFkajlByBWnEKj6aR4wRLE4wXZ+WPY
XJYEs2r9IoN+lAyZOQog1ZSXviEYAgHC8CP/h0nR5+H85WTIxVq5dsHfO+OeNQkU8zUDhXizNDJb
c3Py0KxZ1QE4BlRJjyPRgadEsa5YsESGHarUbuoayTTv3SOiocUSYgw2H+f/uwwHxvPDgU3DAea4
7YY04lD1gNrzYygaFgKRayy2b6ZqiP9QA/9oansloLyEBX8PL+G2UGZu4Oq/7c3XHt5WcReeyJgc
PfHu0eliLFfDriZmkpk/qrXCijrJ9Vyrwlq8GUO9jUgQjCoZqbvBU6ZbQPC/j24hmDsBpngWvUz6
NqZuXyXWRk16ml4yTYUtBxMR28Ru2iN+s3F5/SMR0T3TzG7ONScnIJY22G+UHZlH5+Vqocdc5dxG
omEYfA9sTRX6AYGyv+QcP4sxQqjxS1IBKzIW2LzUxEcW8q6UCRVWIY2VMZrIekDZODcUYtVZ9Hlp
HOJ6JXNd6QwCAfvhK32a2DUfBdorbpNgEKJrcmb6dfL8E5I57qdqFdQVrWzyOWREi9ksvMyrKrIN
AY3lKLLTSkoKpOJv1aJDJH8lQOTLU/iynU3qNyF/dn3PIAtpbJrwBwsQZFctNQU/T5zXy8bdmP7U
EsVT+AJqcEGh2L6xbMCy+HIMVi348kFgqmUj6sE2c8Y4dm/vlHv0eg0QbhXtbG1FJsk5d7ksGNWb
VMSOAIweCRyXqcn6G8q3og3lhpmGXnd9xG/P5NPQ41TVSUnCM64EaPvUh6RkwtDH9b+W/QG70Zr9
rSTln8CvAJzeHewWzGYVz1ZooEGLDDkiM0o13HFb3j4r9Q/ryKikj2h+WFENs4Jn+4JTqTTmiNbM
Nt3D+v3pyRXAA7uuLzG32YJfqbL6wPpaFcmjqIxks+oa+H2leCJbat5soA/mZBaUTO9nbOBCDxWX
iCIygjIBwcGk/4l0Pav0MeusIKijt93l9gzXL4Zk1+4iU1ZV5kvrR/LPoUTkgzYcCWOsKZnW5jce
M2t9PxvsKt/RzQIAeNzJae/7giw4veD4UFjzuehwuyvY6LoLrpx+L0c+Wtv3yCTYnRqkqFu8TnEc
0K4V9SjEdNQcIECqL+ih+iTIaiHdTKH1vLMj0SZSfXkrlAa36pu5mLZaI0BgZvB4yki44wvk2+bO
HEz9xiUnUQWwfUHjqoiXwAimhyJJFuXXrZrUJ4VGTzd7ML69qQTe5u/FMLa5Pgk9mVgfZvQ8cbeD
V30Cqmq/gEly693xEFLABlQl+4IMLzm6q3xX+XltKFqpOgL6VBjTew6NB3EarDJlA19/Owlojwyo
RckOX9j6L5La99b46AfWNs50lhfyzQeW/NvWC3GnrRCnViiKsE2vncRw4YJDePm53TkAXZ1cDWfN
NVy0TQjQ+DcTae1ny7IG3OF6i65YvAqHaIRFYzThFkmvEnVhfPq4wiTXsg7fTsFo2iGs2osOQrla
pUsVq9KoB9luuSRmTigqFt1EJJm0AP4KkvlLgbULfVcwhpBpsxXr5q6IvajCuBwKbV+HbftODTSx
zMno/JitBsFeSZJwjiBg61tGPnvEUOCFnoJ9Ydd91p7I+sSOcPDnV9JY5cGIV7Slvs04lxt4Fi2m
k1J3IL1Bs1EKhuFLyeHA0ZZRwUz+4uWO1VAuZbBBTNA2imyTVHyP/iGACgE4NejThPT7QrdJ1Ww+
Swg0aDJxWcdKTiB+sj8+cEZdUi8b6maoBqPPY+3NKbPDeeBq9X5HSlnFwA39RA003Edpf9o8Ot+v
y/omhVEdL4gUEZzvxFhmR//qU/ap/LjGmN6OlpkiZI7Pbu30bWo8NFauImN3LZxzDrDEwwcPDgQx
uRA0b1t9vDWYyV8A1gxuLbqP6zUyRvx/AeEx6QhXiCNUV4lgI72i1BgtzAr7BAM99rN1z4RqFD3H
TC5wtCWTcZwOXIT1Hm7Ysai/CBaatPfpDA+Fs1nX5qZAzFv0PEsFee7ki4bXKPFBCrZirfOl3yNm
iNHk72KEnW0DQ2LQnS8mM7EKaQbtJqhoCteCBsspV/AtFVPM5KwA04Ie+zF7KrHZLPbt9/xWBqdK
3ZwrraWeHHrzyvImQlwO4HlX9KNeVqk1CI3QYTnIXA3Kwrz71La9Lhu4Oc5ziWc+/sLzhlEVFTL5
t9UkZLIYyJDGf6hue8ZWqttxEWqKExY8B+EzfV6CoGR6/D46bee9zeRy8ce6Hn5b9/CAO013L2zn
QbqvcQySCPU2jvJzbJJIgPc7SPXiEI/uUljd3/5WmkArrGND2Xc3fjm55G2lQcNBBgJFwoXxo9G2
ylsoGxXMmayCcRQIWiXsC/6TpBc4QcBXpQPiSnA03YQcP0ULO3WRxcwn04GB7Xmqc0qrAA/iRcvp
3UH1qHhNB22uNI3StKbdNNWtfC5aww9+GTfzUH2QQnYnmNlAM0F3QyjfLTsl50TqDmqf2yI1Z3fu
NPyupNwRPt5pWWpFVSjF69KTWG+6vhMUGgZ1G6JRvg9jVrvrNksNh83Wzwveru28uSHMgXna9ZDG
PI6ukC9kEr/2Q1uWT81qn0pZZpsJhEu6giC7zmyj7Mw4fXzPU4eIIl+jMLnOKnUh9CLpntNwkEaB
ulhIAQhNW/rExOOWKATWdViMChidU9huhENDVlag84FsuVUflxde1LGDfUhigEqW6rAq6LYO2zld
20hW7m2XGPGoWky/S+h6m7zA9mnVT14nAeXchflY+l8Hz+q4pToOezfN8x/8/iSz+ckpAegWcRB/
VX5GzLbxASsYz5IZK6JInDYlt71H2q/K5rT16G9nvt4Rfl44Cr5AOVlyAb1B2VDWsTVe8u8vlJdG
xl5iMZbJYd/hyQvCSNA7xW4AWyO2INxU82Q4ZBdNklZFfN7/R+YZLjtzzIevXYs9zT6z5kdx0Q0S
uj2h5s7iJ6VhjRp02gvuw4+AyqL56ubcBO362ME3ktR43CUTrCkUBmmC39jtUzz8/mIvv/CTB/ZJ
LuSfeUIHE74XMgoYoLQX25ddBjS2vDYh0R/gphtY4efAKMSLB8x8WX7Mv8p9j2uaWwRi345vi7Fc
pfRf6PSjrdlv2s6NqlsDGXQxQUXyhyBCOg2ELBKrBihU2zmIO42HxdOYw/b/TwYdipGotBB6n26A
NWyPjxYUtOfJMRkB8BbXOV8uXA4y4bNd1/FbO/IThtFzgzI4iNYMBcX/sS604T3dMI6jQZad7k0S
IZ+5/fK5hpkKghWsYffoxe7g3p268oFhyjH6l5dROofzgkHqTkp4x4KKdSXVVa7lelX7q4cZ6oGJ
DMrP87CrnMO7oNy2G1S7AFdBfLkvpp83X+HIEtJE+oj+7U+6O02GKQJYYrsSagptTIwF6X6u4mag
EAxOVSbD22Ek1bIA6tZWdD87ZTVnrXin6EK+hlyYQUa4dAjC/SsBFnV1sZtgycsdwG4JkeSZ1iwy
4C0LSShAygOaTaoinEiTDRxF6qX+dM6UQTVp/uF+w81dfWNxGgZPaIQALl17Db7Sy3pDJkwRYA1A
PndAiaTZn2j1gSgZMjfXxuGaB/0Jrt5WfS9AsDCJ0Z7sPH9wb8DJQfyqHaHJBX3PApibsWzZefdt
EWQ5nussgcGkTytGkv9irepGGFvFdlTpheEzAi2RWjMA8pWmq6SNVUs0Vv2iW1eIfb80ii6WGzLb
GI7WONhPMN8/+jYQEi6+Kc/r+K1QShOsMi7VSy7h4y8h82xnRk9wi1uPE/mEW7SCHE4HQQNQ+kZ3
42/TYtfez+XtzeY0dFEjdcvckvDKFRhRvi88UH5LA3FOdzLqFtUWQBy9kUm9xoVXQ7lpixKYyhOI
TdJzVAXTEsqqG1AtD1XIr/WRB+voR1VaHCi6o3fYXOfIfGn/5hl4hW2zfw6rTS/m+FBcHjQkaF5F
KhpaO99YOzUFS4vErskwp5ZBvw7rkKDkB4K6zlRVR3jzxeOXzpj+h08MKSQQfr5QBFed18/ykwzv
AnjI2YRytjmQxmBiSqeYXjOUsfq8wFS7mf9rm6/ExfaSoCyat5bdCssboicIgjCRHvFjqG3hGwv7
cZcaoAt98qv566ElMGDM+g9eaoN53hoo/dqKNEeQhrY4CUjC7BOutbqRTPdlDW+WavCkMFjNKfur
imCWpMdlYnzRXcWSEsz4FQdMhqJEbaJM4eHe+wazghH6kazCzNbyi9u7IxNwfClxreBy/y10Jpri
k7adM17Y59KvmgMjDhEfmUPg3WWdMcpskX13RjyK8IKSt30H4uJ8F7pdz2ax3YOpur8fyY/iTr8x
lkY4NvhTdU3oh+sT9xi73EMvCYUKZfWa5pRjs2K8G/2QxuOdAs35dKYoa6A/M4vV3haSQCpXyJd6
SMNhXUUclQNR6vxmLO2aEIoThmTWYmGzoBcQXsabBCwG/NZ8w7TVsaWC97kUwxaPt3kQpHXnLcSX
sk/0MYs4UQhUOKyPi4GaoJ1qHJaFa0/jyoywMCh/VFBM0WULDWvLtIjVBiOovkyRfcgsDq3IqBOG
gNr/6FFx12sm/eFoX1A3NJBO0CzEgQ9DWCVHaA2MSZ2IS+WzEiOxIOLCgdDlo1lLvP1XmzrgYohe
oiQyZ89cll88mOjby03dmafdEJ5PYhqmPnz6OWBy9+XD0An7ohUnlc8QaaMRWIl7975FPeVdRSbL
pmxx0k81bIcOF/cejXBpYT/YjiJKfZn1whADWKh6SjW8WLnDCBO/dnj1yT3a7rYx6DT9GPAJh6vP
NkKIOTX7WqGcoKPSWzG9q8NrkAy12v/uqOY85miVqly+dgVozLZ7p8dh0Vq287k7CaOgLaFACjRt
gmfJgoLnbXzyyzoz0WUC+miK9VcYPQXsw1+kzyIu8sONC6Rgd3YGy4Ybb0ncfgz9RPaMjAIl1u0w
GnZ9hajrqXtHhZgjJJe1ForNVbnIOiyr2T05i9dMFD1Ub+uC6CCpWslSabAQAVzsHtOMUEvUcJul
rn8BKfXgzKOnUB86QoJBpOJ4UkHVb1eGtmzzPvzMLm2ozEiOqSqYMdtqyiLavt7xuNBBeUdbSaz4
1Wdu4Y7LrW9RzXiz3kdF2zES2vinCJsmirreSw50NpGkpVq7FqN8R3uux0QE6i+e6hsRmrd+MQbx
ff8YPoZI8DAQSf/SR4McsVmYRuBwOIKiZlP9UoLJOYNDMVi1Hc9jW4s/HvFwbNb0HIphKTGkyhv1
0l//5cH/sjPlPLxVBGuky/PuyNUtNv91EAK26nQQ2MrwQqJB3JO0LOnHPKZR2bSVsZREobKFuwk3
S7D6iNhz1loMDREbLJtSQ79Y38pJEtkCmwBpZAMjHU/6DOzeHOylT9PyNzlUO2sugc1MBMO7SNFU
eVO/c0wB2Q0ZLrmdNoCGjY97nyXAKiPp+wG5Z+y+BYU9laUuCk90PBDcqFKI8/RpqhqKrSYBe717
ffB05g3qTwO7J4bV7SnR1LtufWGAuEBu7woFNEFmjldQt+7jVc/AHq2R3UxcBGBt0kZozWby110h
y2nS3H56NVsQE5XC8DcektwQDKMZzUvhGQSPB+qSmdqHelnPV/mWymCUc/D6uqPan1JButllkdug
p7TvhcnC1weLz7jg1KcZr1kIC0lzveigTKzf0tE5NKzjnelc2ONdaLwgy3Q2wOXGTwBK+z5bJ9Ss
jWxZvdwqxEcZqxUZAKmxnikoGy4i5suTCgWEP3iXflw10PzXtyUkBD/hxC7DyQ4HblZagg3y7G2o
oKq9wHtwhhmyjUOoFmC6E/QT0y6+fu42JF8QsM38jEe0JuiAen8BGwQF+d++EvhgC/8bGy+GndYl
3w1xx5EFENsucJndyiOpE+pKps7yIcauYUz6+RebSmFOSZ/zWL1dHhHXkidfA1xey1Ng8ZggVDVu
Jwt9psofi5JZTRJxWVkCJJj+MOEMEBs2IyLlMf7TJznVSwhrgSsp4+Rj0fQB/fCM3I6moWOaGt0X
1WDnPR3UiUXzL4jph6WLTDzI0pMA5F5rd2ZNz3X/zqRoNgtm9UlhWYXZ02erKS54Tll83NzDR7x+
v0v6yqcQkgGY8BcrU8tj69WW9/rJfUTSOJBattztW/OgLwor2Ei2RBJeb7TizbIcjUpLY5JzLViY
auBtEh5rVziDRP8Okioy9RCupwSuIy8O1gbwPOxXqfFAHPs6u7TqIh30oZ3y0Zfo8FC6FgmK1/qy
IS+9pXGlgkMHmhxNmkCyPXG0/s+ZcXGO8zl0Y+kYoXdYaQeLIHd2TLxTg6eemzKRjAa3CERWiErz
qnp5yAgXE1FIdoCuVDoPEaMdm+rHMx7RA58Gu3h/kzcs+I2vL2GYo4TUS21PJQaM1WyMOKSSYo1V
qPeOUeYBeaJRBasnT2BTAzZSgOpa1pYcDshGSEGE06txhZscpsKziMWAt5ePhogtwROdF6iqay5L
3kQhovAh4CSTrTrwYlDUMIUWRRgEODWLdGf/KJNkotwb6e0NHGu+2y0UL2z6o2sHK6sokrEyBg51
1U98MTDVgE8sHMntxxRznbvgOaZ/JOsQV/aKLf3V2EqXeqTO+1dTCw+ckCUcVDJItRFauta3qRHZ
Nod4Fm8aj2Xa+/ZUOPb3ci3qBE+sqykokIlsMLW/QdSY90aktlg8Ah9Adf1bjzFOLKXQScrTb9W1
2sDbmm7k6+BL85//4B7IwNonU65B2e0MkI3ZIDJ62+5m/7SlvMbibgv9mElakg6r/zmZ7XPFIZQB
ahmt+ZSlaYUl50Rfe29cD+hNGGKJH8m2KcTlC9zqqEGvoZsp6OEckN8kWO4+MwyH6dv2+DqR4AK7
PjHxYXpX4Ego5SZ2jm4iYVHY1T+8rcxH4oq2jmtYAhS+bn/Z4iMsOAO+MCWzFYkYHrxYfyutNTDi
kxT6nSUWThWD77w+x+aIkTxapKMfTnBr4p6OSoveK2l/B18ibcyTP2Y/qhoGWPhDcoNw7SkXfZml
sgYUxm8sjlWyGcW1uCN+ErIhZhhdvF1BcU+fZcnM3MS0AugqsLYjNu0LrnsZEfVnEqMejaI1F0BS
ZzVVnEQO+1VLlkKcFNk4i5XINLkgY9dyyU+zlSUUJv5pa1CVrEfkEYjYyt9Zv/Zyh5PNjPVREk4e
5iiWWWjYr73bb7UfBKnWma4GbRHClrQR70DbD5T9LEdxHn5uY/CJAIgC5VnPQFXT1qp9vlhOIflf
sD9C5JJlhtEv1QkFfFEQVHQLZV2ZPxgt7UMz+kg5Iayvw+LOeBmlZTogUIiQmijR/NGiqnDm378b
o4McliArQ73VmgeErCNQNHcbbR8yJvCRN/vxAj4HksTf+YsRpbR9ZiEQtT0XaeLv4vRD8s+h/8PV
U3eML2P3raZ0KXtRQyfZk3J17rn2eUm7aIyPj0MzuTyZ+hO6Z4ph/9elam6pU1qqy9nsGI+w20Ve
1imPpHwuX5G0ISlJlNtFemR+y39bggxVprCOiW+2eGR7YNnSSbtj0vQwFc6nfRDPIN3pRxv/e0ml
KCpG7sksLT3CpPhrVVu1tRS3uoBVMvObmFK83gSzORpSaWjt0uElBbFc3apEzSzqOvT0OKvlccD8
p5aphTshsaDpuBalCfC/8y6BvgU+dhc4rIAwrwvt3cKs8fKhYuDtGQOKDfTq24JsEatCbDnrGB6p
3EGR6H17BaGEOmzKQpqdhb3h9LVyR9w+geK1YeeclpSvd0d2SKQ3H5aD3ETGuDr04WC6MDQcptez
eL32v1M89WLqamRiyvxxg/wBcR3YFz2S3DZzUqzfLkoiUf6uO5TICz+DYnPF13SMfLPz+tgFy/Bp
ehu8Hapi6t048gMr+CAoitiTTtvFvuRa43nejJKDYukw94m8oxgNueZkNGp+cknpJ13VXMpA/MRd
bYCZpMLbGTqlxxrOEHAAZ6hhXRaYFUy1q8fcZxJRrVRvwaFbrYo1+JTbMrX+HMzE74AmiUlhohnJ
jE7UsXrzOhBE91fP+4S9fkKq0y5soMGdrehG+jk/o1seUYyVnaXCSyEoiYVDL/RmwgXZYT015GLl
dK94OSfO9KxQKCJT8erf4O5YVr4YeCuuIL3+szunLXR5XEQhy+J87QiA1dIhpBSa7XKIVIOawssY
rtwltFftt7cEjhE12L+LREZTyEZYXsaZNpobTOC8gI+7kmB7g5QTHS9Si83SBuD77VuYMhZW0RvB
uapAym2IDlDbU1ZqTP6JU1fpbTgoJL7T+3m+IJrmBLW2HMHMjFntUKXH00yMKyM9jw1X6ILVnCNl
aqOcbWe3SkC25GIys13XnxZXIJPbCDjHeIH2viKMBjMJ2HIg0/63gbTbU1dS+JHVqnhcrboiPzH4
lWFRKekRwd6vPg6Jn3wTCiyqQzGf61lzL1D8Ug8Tckc1gvRowXGbGosv62D4b5Jg+cyHeEXSwdIt
yT3t4I0G3VMSP6dIXGixWy/Ne7vNoDl7yPOEmo5hgcqZdJytYXNxgIcImpRywXpR6LdPQ76r3sAb
LejDiphZa5AQDQVKI42vYZm4nqq95TSzsZ0zLtJ6wBBDtVBCQ6PjWCj7z+gvdwVDXd+0BqcUrjNd
rNiYe3rIJaNBqUERcrL4xlbhAtSNTFYhJmkwiBXvj3wHsSNP23Sl90Kx6kgHQYFkbNpZrGOEvJOn
XDGyfdSMyWKFL7dTT2rjQLdgcQhcoa129JRJmMlodyTpwvhIfNr1ffxL24YUhDeYUzyK5M75cokx
2Qd4DhyMVRvYlXhJ7l7Vv+kEWswix81ArPCTzxbnpdo++YzvpcEbesiN7cSyARLsDJppMMZkNRfx
6Ew8bs35A7CUyoH/lxfqmPIc1ABGqwVR6ip4gXC5VVvVZ282ctTu0Edks0XBcaTiPlbBXhetcPq1
Fl6af6Bpj+31IATrlablP5HwLJ1uVr//dad949agviT3aUnJ/rVZrcYEf0o/N2/mZIpMFG/MjqYO
FfVobUNLNXH7vCLNpUKxdd8W03MpEYVbhDbbvFp7DTWarB3ukYiYNH9OLObP/YYN0mTk8iadNDy2
j3qqCS2F8wA7gRNxvAa/eS/rN41iMG812XrmlJBa33npon46lj+NCEOWjZZ0VT5Pm43FJw+ygk4L
3lhr0tLeSbOBZtV0hA+qxB9HnNAvMVKMOAfs3vaNBAod3cHCbcSqxreBWjwoxRp8MAPV/IPeZxoN
27jJxdmdt1UNvt7jdfKxT1f2PrLKnTeBVoKP4lE5/TZ4q7fbxLvpcR7KMfbf1I9g30X4CmGms9kl
yot9xpGBqW5Bq7zLcZIMqmV3NyQv8Po4Nha34I+SSrrOVhRgx0orwQo7QJnMqXBqHzayJI7iYrOT
tdi85r0Iu+lt8xTnUYmQTD+D+Ivy1zsixODhYRGNF+YNUDx3E2fQa3KLhFfq9QDWsf574Wxdkmda
t1M5XLRMJWSfUmCxMMHBihFmsDFWUmBD+60+kwuOQeGTvuu1N/f8bbvkzFbR0S4XzSZva5ese0+W
xoeNCHYgMokPzsu4KtV+suu3pU154S6pAjvXFc6Z5NeMvJ0CXN84NDqzVd72uEBv5hbYWBXTfH4f
6LK5Wtrsvhg+ufq7tRYSdxQtvjPudU5wUlJuTXDMdgMNrRQXadT7qweX8CjS6jiU/UYXMly/fyio
8x/D0Xp9YmUnWvKpuCMAxmDNtVNHNdYx7SRotPFb9Ni2Ubk8plgpImBaCuRp2zUeRS3gVGKETXaT
AmZhlouO/2cGIgfOnr5v2I0sTKR75NXgbPVFpTSh29+QIZqPu8mTByxh2bzMaofFekAB961EXvOa
e1I6cBDKBEKjfc6GRxCr//wTBaGAXF9zxOvgnngAcagyPc6SZaquqkigyy4DRSJN6kxazZQmU77g
P0QDKgQv57JH/OIpm5vRPpAqQp357lWkL+duy/yRBo3KgjrZq4R6ulLHEmhKpr6jUJvBKFcKpjjF
h1F7ItwhEBoWiJpeGNEH5m4KURXI0DaUDY+2nGsl/IG21tphXnPg1o+k0NCb333JIIpdRGYUHo31
WwbImXuWE+w9Q4d+p/tidi9x3BFix8Yuo++2a6Osw7n+QorkAqg4Fm/hJf8GTENf7vyZXE1Pf0Rw
r7vqqt6L/FNUpJLng1NMlU1fQNMDVY6/3O8S1UC8hw/GpGVbFqbAkQo/0GQ//AnT5X0ulzOToZIo
xGvgCYP8IlhopHB6bJ23l0KGE574OLy2mNpOd+OBFtQlVzJrQAFSbHNilz40CzxAmIPaSJqKTGIu
FJBWBR9ZRNK7xnS0zy6OQ38hLuHQjqg4afQk8gkOvPuHY7kfQNiRpp5a+8CXD8qFrnKcKX3trdiA
tV37oggS3iBhq5S2CRmbkD8bxVepRZ2o1prYXGGAKUow9sCO9sZu8BbGKsENJWyuaM60yFrayI3G
kHGVj+sS1BKn/eSjP6on3S1fs4WJ1Lm1mGaBNsd3uInm5wux0luQswbh0GZT+ei90JT+0z53Lm57
E8xSqFafU9AFrq+8ZCW7phpAHwXJaYb/Qky6AA6GnGtMfRWrafNk1DVoOZiqbTsr4/FHnfDXNMdo
hinKwcc/FCdfovT0kMMZsEPjgteXmY7CF+xlUEpkq/n97JOFfRdNLxo3DnfRSekmIZo+lL0Lri8z
Z2X00eBkL//613zzziVUA3bhage8iGtd11FrcWx3LjHm3x2MamEzK5/2rq6F+obyvTl/6h2UnOwP
/giFSPCB3ZBNeQjAmSFOIbQ+q+T1JDG9L5vQzUFr8lYbuwGxXNaBIblLjRi3LuCpcmTsV6teI71D
mOuwgygMm4DqBGYvW/wzkpOUYYm3Gn5BF+gkDJDsdmdv+ZeKxs1oAIl6OEr9wGQpoAoz2ieoIPJb
NZIv6d/rOBFBpvubFEBhLKQrpKUSDDalCZK/oUgODICc/ORj6WopFlC6CfbEQDpgxpaiRP9CXLY/
7BVQYjvIhJ69EMtIrMajUB9ZMVILmhkLECe5uCIwj3F1tJ1EzXDa/k5xRoe3zPc1y42m0jTcpRlv
IUPQ3RVK4owGArU8UAFqVrzoGxcI33ng+YIdEH+dBpRzmE94iVOlMPvQ5sa2T1K13rjnXvtMTvmA
AKAprvQltbIAC7i4hCxudm7W3tF/RvFIq5lynd/CVmh/0f3gpZjMmJsgr9aBIolKiy9mgLR79+Kx
3X4VJBNU4vodfG+XtwqI0+DLqkweIPNsEk9uQT7P9em6J+gXnSZYTzXo/0R50NPAV1XuO1a50dKN
WRda2NczOnHG5wqGn+J1MWlYvy0Ejx4VhhUCRbsFyesDlJjgiNZrI30H46hMPAtfyQJXC4ltbsRy
4uvf/1+VfnMhsH9f5RE5/AgxOKIbKmERhGevHyM5RspwHn+HTG4kSpsWuoiRXc3pTpJ0vz7zXmju
KpxBQHMvp603shVU5XcwxYne61U+lzkGdT5HcIER7vI0+DTXYzqMPmjU/uH0HVUw1RGtSxmEQJ5S
6lr9DB+qdJzgJJfWy/tF++DYMMypgbgBgUT0L0geWqtbIuBpWOj/g+E7HE9iE3T45bbFD/D2T7Rl
gsa2SoE9cTnKM6J33ecuj9TgrKqVLnfdyvxf9jlx4dbC/WrGdyHHi4UEZ4CSmsZnofW/W64egmPL
CmNVmYxpfJdxiAsBgDHUCqDF23qVlmT3bgsC6IiJmKvONyfgPUAYOdQbM2zdyfZSxxdnhtF4VmbO
1dYssL1r7QW76njwQkJJSVwFE+iT3LYUeIcZGuPXE2NJ4qo+XhPIiD4m+8XldL2scgw8jHZMpsvh
XM7Heij+BRPcCVXGgvnZKuoLw7t/oXtzdhRvog/okrbK4IZgH1lETxK6EE8/9i1ZFvp5bQdLrO+j
dOyh9PumO0Du2+azDpmuMv9mUaY9GpdKdLRqR4BWujPlskNKZ5JXmgyz8Djp1zMIJAP3n0GoqFI8
NJeDlPc5TuXA6IVheCPnXg3psoBCPDdN1ugmJb6lF9tlGtr2qfIhlsNRMd628XkMZwZ2rlwb0tBI
WeqSz1Kr2SjnpiEPvwLwCHjOtiF9RisyrkX/umB7qyW9Zr2gO+VPqlI7Ju+QK7hUNVugaaIBeBCC
ySPKbHQRNgkLq7dZULYJp0GOTqGgib+8RDdEuA2z3YNPzVC/YgDyxW5cImf7u7d3vg9UkpJQUZFr
c8f8H6Sjet7aqBcCNqgxj8CrHg/NOyk+hJFLAmnORrU343xXfDCOz5hsP96g+AfrVhc5618o6o0s
G00KT20fkrJZp+kzC0LqF/5lWSBWq5kgmyPqk19X0MWNLkfeP3LvDkwGTm6oWxJDGq+GD9izKpIU
nnGzvCUdyQM7v2pResTTRPGXy4GbU7/hAMT8IRDLi8hupXBC+FCBcefLpVEYGCIDukR1OI3+3PBE
zVPgypkTkT9y7GqnsseGuiHB2wXLvD5fBYyzAHdxz/797bsReU9NHE10dPec2RyT4UlrAd78aGzQ
FPlzfaIhbdxqCkD8fMzjktf1QQoTYhKXmMQsqQuovwkc8ZVpTAgw6qFn4sWpQv3Pv8kUryIGqCm3
BQgFpamEYpkFcBF1XOkLHhsgdCx+I75xOX/HEM79rx5OtHudma2tsh2frEYG2yT4cu7FcmDToLYy
+mfCPQXkHD3x9T7EquBnhmVAGZ4PuPPPbpbBkr2NHuaIl/iIp12F3qvn7yRHnGcCkYGJx99T0VF0
9ESO/vB4ClEZVsOsMMIiMlJcmPiK1Q+ekA5CQPiscZ6dNAvjr7udpbJw7S0nhxFAA2uT+M8t/oxZ
+EeQdCH1mHmM95wn0mqodadCc8PYxx1Orf85CfEsVwTIXZRSp8FKKKtIWVqtykUO4RoqOPGkoSxZ
JtRKARmyyUTh64oyLMqSAP8R0/Bzu6UvlXm/1dLjUNAbEtJg00nwx/u3W5jA2FS2NKoywQp9ULNK
f6Zl2+6qMz37QyQYHjLasdnrMu82shC/tk0WZuN1JR6RrXU9i1LgHPGirYt+kgZ6o25r7AsgAV2e
yiAFVwSr/rUn19km85xWrEGq7h9K/ylHZRyfLbNtO+iaOnIgY3FTle2Hnb2U6dDGKsWpAfw1L5q1
cHqk6n0MR6pLac3mmpubxEAXWvm7Gad6z+rozubo7sPTDasY1hSMwURYRiNCEYrwKkci5vS2i3nA
Jxk19aONASi71ug9m0Ic+1Sqef65li0crsijKI9r/IzG2fOsgbV3xGlGb/R5/n8UeR7eEM2zPPaz
fQpggoRGfeZdtuYCMLh9T2y6OobQqvZtPgASuTU0l4wre1WjaxZh42THEFnD9AYHqYDHFpAE4UXr
jV+KNTUxQhPQrBpcWyecqkyXqSJz2J9jsIzfmRvPoINRraZvoxsigDAm3Srq8Umq+dKulMydxGl3
8/Qrb5K4jZ5vHOi9bpp1we4yD6HkLvFknEk+k+nVZQnAthsQWetQXpmCAfVLd/9RGvt7WA5fpJoK
gSMGPDxqGaI7sA9neu+7LAXIOeE14h2qPjKDXzKsMGhATyBPDz7LNEAxoHoWjHYmipK8WtyLVy+1
DkvZa1pkr/stbWNJfSra+oSwkiB6o+gizAMUB3mxNgEyVLfa64oqE9CRtqFtPmkTk0Fk5xZBNyGj
Zn79/qHfjAktW4f7JcgEHHK0+2FPyQNbvvXvKMfKTmhGmNn2Sq6L/Ys7pOB0/KTP9YYS3CRBklY/
Sd7xpVxbGzxXiWxqJSzIRnAe6whAa/TVn30r1VZ2a7y9N96OutG7Nn/X/qvxfHB/ZGPRR8oIvPBY
fwH6O+aWdTl+RLomHLZ/ApqngJLRzDA6W1WgbqClHnPOrX9Y2vjM71D8EDgBnaQ598RbibjmJZzu
a35fUflZQSMRgzmMm/jb9zzZ0kSEZQpSw+XdwAsx59zfd+mat2524fJhnq4J1AjnbzBReUPED9Hl
cYk37uWmPHgCDtxu8tB5rGsExg6FxOYem0RRJYLgjkXd77mUnH6hkdyNE2iGGuJPUgdGtqTY5AN6
GNIYuDSvJYGS/GhspY65EpS+f6c68Svki+lXB1lY1xfCmZTDPT0TXPZrtVII4zRs8nKKsp2zoLSq
2pSlfXsWVZ9wnx/geiLRHKICe6O/xDaTs12gxppNZqRJUuqZQVjxxu7rAciVTUrSl6l8XjruOigI
o3WrOdYAjpijiAquqoUmHMUkMz8ugjsObd43WtnBw166dT4ktTlJiMKm5I7kzOqbjNalXsJjy2XV
GbSPxAlZ8Ro3YHksibLw6loOY5zmiUW0P56X4CKX6ch43Gftn3FuJttBUqGCdeAn/NlCCgqv9InM
wKjLgZiikumwv2GFmuAa9rLEsIx2WvNFyFAWu6bggzOaHaj4Ccn7Iq0FCyeujSkTM7E3ml2wG1Tj
ctJLePemfFu0X05vIHIKeb40OINh8UnT6hC/2u+iZHW+0p/6dUC+spqyiS+RndLz6tiLDEVl+Yyi
9BH85J+kH1kuUgKJUazdghgvMi7rqkz8Xv7SMhOivbv5VjtE/PW0jcQJR9eUEvvRtzzIFGdlfDc2
6iPI2VVPhsuY9LUu34TBSNVHYePM6Om6lXFRqNZ1KC6AtSH+mtuCfE4zvEZaK6lL8mvkQs9YAwPG
HqI1SIz+8TOE8LWZvai72ozzIIBhy6Gz+sYgOzdDux1wurKuY6G4Hxsy5/lShMWlubavdx0TJd8F
AFzjViOul6f3Aj7AhPDZf21O4ayffmyLn+Iu4Ae6ukaVs+B34CwiDokxwiMFKu043urfMY1h3nqo
BJJpLDfYmpFspqtrEYrYqjRESZ3SxK3mbROorUFSL2aS1GP74tiGwV6lTPBQ1XSJejzgf1WM70oq
tD2qZMdy7aJkTlI/aOdVnph4HbM8RWIwqaeO9KB5WvYcXYaMISkums+dQyQqFBqH8k7jMYYjn0Px
KNlVPQm1j0IvPMKFwEZtaHrQRD3xCAOtza6OMCWxNOLIjVxGBssZUTaF+YXwhtjaISqLG57NoIfI
BUp1zTIpXaI6mEQ+SG86xd6Zam7uNCkISrZPI2HVIY0Wfjx+/LsYv6aO0+BuBWman/xDc7WynITs
S7GnIBkPkkq+gwFQAPDOwvfnDGG2BVVSPuu38Lfx1liBg+pizY7yREBLGBItRRrf6CZMkQQMLXD+
Ir4i4eYJKcYfgTueTMTs5+0WHbxZ0FHkc383ddjLeuKOIy7tBpSCqrg+dAle6SboDIpAPZRoBoi5
ekbbDf8gfb0t1zOTlKAoaywLpf8ST0BuHzghRyhEKk9DzMzPCy/YkqfVLVESxzc2icn+9d277Drn
PohsebZCSAkZ+rxSrhzw1wt1SWDVc/iv5sekDN4rOoKDwCIchFD+fzx8b/VI9i95BH9C//SUEz7n
ecTcSEmgodsJsT2j6zP+I1ZNHUpD8mbjKyZCtFFNsClUdoqb1ZUsg6M3+ie7JKbgSDF1yVv6QV2c
4OgnM8AHzJqwcZlhftW4YYY/65l71UmJPvmLOAEJZILZeEyGQgFEOFCMK4Yddx3fOsk4zTK91OsD
BMfhmXAWxiFJlf7cQBbYaJWaAT46f4AzDnQ1jiie2H0CmpV6hD2yfUdTkuAYBdVtJBdwQMzFW8Kp
ERH5rbyAdiilksPezIrNneyARdK4WuYucpz73H+/X63o+dJaS1PPPWFir5hFyTVhfnzJ1aiGif2c
1Gj7eOVxqzlW6fXgWBF3NUjVtDmIOyQAs5ZfO+NOiT9PSxULtAgJilYGniqkjMmZBdZ6RxHUU1ck
flB5ixT92rlcVVE9F38IcLvNTSEYem7hXihA4ZKOm5bpl1k//TcreJFRPWcdorNlinxuMsKIU5dr
Zy4dCOEUIv+LRvKSKR12wsx02fl/U6eGQkX/DXl1iA8z4mIkeOAI9oZvu3G5WEFIdvCv8J60B7v5
y7fA8yoRikKoY6puGEUiqSFBHSR3stRymn65zyUSDoy8pIPGRYjIGTF65ATN1IMPybRjAT2NgUBk
+PtI60CzV2o9aUBHa0VzQvyrgF9QXc3vVLFy4DT9/814etguCrNj7qpFwHUDGYCetjjfSL+wmtJy
EuX1Dt5nzxvmFlmJCpKFWdYKE6hSMA8Kx/MJYIlkf5ydvvP70GAog3YB1hrawEO6sWZw0BI5cKv9
ScdA8QE91LdCOKrXi/WzulZonNlXe3vIYS/UnNqn0tN6qGQD7pCySSeG4POYgVomSKf0PWBOydV6
QU43/zCkPKvBh2uqmSkvjz/4LD94bNXY62ZGo19l55QplT+3fhKZ2iy9INb2DS6UGyzgoxEuJrKi
w0MNul/nR/KtHi+Uwy7NRtoSyeElbFMOmSIBRxR7WLTJ04xeY/eZ+sfnNyk66sVy6r6hV0iZihwR
KlznqIz6/ALHl56meaymeQd3S6HpckQrEE1yxFR7sT4gJDrhr/6sB/vzQaUPFJ8plccYNucJYTSu
UR6KXFmqCPmS5vOy/PpNK6HT8YiqV71MRd2GU9wsnRxlqY15mpVyVVfskEtNz2TeCdXehvbIY9KN
1TzUXMOrcsqHusWf3eFlSvBwZ4eSetoyvbrXG/+ghd4vMO330FmZ515NmD+zbwnlGRFter6XYmwm
cs25b/nAC5q/fIn4C8oqxMM6zADTJOLGzPb29u7/pUyFeKF4V1lZMUBsQCxfa4mFzL5Uw/J9LKxe
/wnqpdN6f0EK1RYTQ1RA/X2fvVnbDnPywJRxqMYoHj0TKyIHMljO8dgpBxa7GpWJwR1mWmlbD0YL
Vr+CDI6DGRneLzD+08h6fU2OEXvTaG+djKHV9My5v1bUFDnMYe6Xn10glq4h/pCO170SyQdPoplL
8sBAFJa7NJYu1zHV7tzDUZO4+JuO12rCDoBxSOZOpqd+XhS98tJlBs+/8Pflgj+Gjo/Ql8brmw/I
9J1L4LC0IYVQz2zNExpkIUON4V9z23mZ0j3B2mlU5lLGqqHXwF85dslVSa86PoThnXCopF56XIc7
GxVOWf62W/bI0kDToR2dGs+MT3uaOgguCfjuxLxLIEoLOfHWExQzF7Z1syFsla5ryJUYxZJJ9//4
tju6ZkCrySAUoV277GTHOMCz8HuB/W9hCfB7cIn7VZ1ETCM+DLlRa65LGlVGRU1XTHt/f1XFSPoL
z3ZJAnKJg7VWZuNz2fE+4R8SyFv2OlUWeo1i/DQYy8ZxBMlpyiWudYy1NPC//oiozRxiD7rzWZVm
wtW4AQm86wskGUkZW8h83gRh1RFPyy+HxZyr7aon40E7U/x1SL8q0DJvTMQqQCCEBjOm+pdZa4W/
cDv3MLTyl7hBHAESaY0N8vMSymv9ku9y+/kyc+IeV0Nq3+RGH4aK2S1WfeJzaJLi7Ub/QiHwcNJ9
jhLI+fOfLE0qlL5xAtrJUa5gQK5kNiJUCgEdpOvw2l5dKWp8cvKvs8OlrAbFOm2cAdAlrRj6I/In
hO0DwuCvGVN40zmckd1qU3OmNnVW+55F1Ambll++aVWdt/ZvVlXaIvZ6YNxKof4/1U3zG8epRK+J
laovTKpyNCXmYJw+2qBc58HykswxpS6NWYmGi5j4me3/whqhod9/Sei8GgB10YxNWf96a4OENKVg
brWKl0JOFUiz/4U/hc2rwijJsVSYDKP9oPmowqRr4OAd/aTivEmLCBi9XnABeg+nxInFmk7aJ/+y
N+drY8iEuedt1UtCs9FKvC5fw9/Snc/w7ch2u5wXjsnq41CaBthzhFPIcucQ3BrOF0WJUyOzFmSv
nKV0eqBk4be81mcF3LicA/85D1rSv0CCB3UOEoZe6cSElSqvzVIhTDy3yBVte7QCMEWENoNBzLz2
CPUA6HYrLPQAk92ooHZ0fvkd4rJTlew2mxdcmsVZFjHCpxWTvMUybhD8dfaaT/fxHmsVZYTmZWtq
7JExz0rls1u8Iw4f1Z8RsplS3bAC/kMmFXLEHDBCCBoOBWOgZ6jLibAmgdrVsIlb2Fhv3t1SeIqQ
MI7nV6RzgQkLnojWxQjKNQXGYnV+VPxeCP1Ta8LF5qORnKOUgxZ0pb+7qHDtFAnqIl9LOML3ejr4
ZObB9urQE0WBuDvtBjPV5TUDt6qO+guXszZNrDNb19Q/j2i0hWV0HKoa9keyGnIB4KTOYYO9vm1/
4k26UNXtoPLUQ+fsT1V5I2tQ0ubQbSskRsKe15fWKvgXoVKuBUDpfPVknY4KPLTPMae5z9yWnnuV
ZdM/pkj7OQ1zwKOCh77Ey5QMs0hvdS+5eukL91lzQoL15g+HSmzXtldkcCibOdx9b2+A4hmAQAgd
g0HJJOYJPEF2UNj7esyuBHHxs8eDdASC2I/sj87tHk+ub8PqZP9Deo4mNxJtOn0uoE7G49v+ji9N
gWRFkOCXJ6BL3y85kgH6mJNIlADZMgANo7OcUpae0Dx1LphQvzghH59edy5Yug57+KNaATZgYPdY
trBOer+8FvfKu7bJYPrRA6/Mxe3Ujlc+6/OCHRgi6MSE9SKNNcgPqz9sDp2UYIbRdkhCFNdOGIZs
Zh3LHzMw077v0qfWTNYm/kjLuwmboE+XXpsaGaNS+eYv+cFSFup3CPmWG6LCyLG//6QSRfR94XDJ
3VwTSurIpGAePA2V276GKO/WKMec57a+yRzr0JnEnhGbVpmXKEi5Bx/3Z4MSLfQLeyYxFkEeUOSh
Y+83sDSQN3MGAeuGLpicC+6MFpQ7J/Boy+UQOFtp0SkwFm/f6cWKG4IR764z1pEXghZv+qh9FfcI
fxd3YhAKawNVICpIFALA52dPw9m18I1lWR0H/c/MqvVeMoKmBzQyU/hZtD1ugQcATtTOVlLBrR02
tP5BDeTnO6BX6zXnsJuxFztuEacTdvt53kpJh0OqsyxjjCdj2fPGAo6BF+PpHuJGjZs6NSP8ai/d
KFp2Zk7JwofnrOqaVXQhFQdLlNhcesJyOya02rlJuICNdjHmlbsK/zB5dzL+wMNnBoxgvwBVmXQO
Qgwlt4dqUrOuBbloycfSuc/dM26urxnwDfYIeN13WPdT5YKKO43RIkmKZ4VGnHn7lzWwbtemoLSV
QmqYP52nYSkxQg6o9UwJ2fmchUAb30gTHM7ddQ9XkLOC16WQUHHJDODdZETWea+5mbZvdfrrfoQt
yaplHQED4neOEWDiO2LhXVK0F/8HT60Gi0L010e1IievIfQNyNKXw+PEG69wJC0CSzfqrWEHO45R
WuIg81cu2cUz3kPWvn5eVtZXzqXuVqRdRKmL6x7HrtLe55wDSm0OMsmYHOledE61z3SzIuHoJAEV
OxJKp7OKgfXRMH8bo4deOWRwW41wYWRRpswASgbSC8co9+KrLpUrOM/yr/bjuUZKkHpnt19IeGG4
bQCVM9VfDW6YRXdZswkzig+uKd+euBP+89+09ONwuHMQz4L0WaypY6SaaCp922ondsJnjYDibMC0
ONPycs0f1GNcY/BFV6Cjndza9DKeHKXbqejmRgub3Atjj3Saop8HawM1PH8KweqZjD0l8oIUGqbU
ImQ7Nw9H5GZhiVA1Sycq65TL82yDJbntV7k4WLb1UEc7qbNuJDxwzYC+a2JTYlm219Hn4t2v6V9+
myf5kjvtlpwqPhbMZgPgc0e966UEhvjm3iy9LBeQykMzGLwwPmlXNj7VupOeZuekS0NV64Kdz/el
Ams5ieYI4+hrQDFw86Bp+d1V+ikd0gdAlFpzhuVwq72gZHim66r11x7LQVeaNemUSmoBvhdKF/B7
Fm+Ywh3FmMMXb9gwSZYXMtI3MGfmCdqPUjFjKPtNPIjS9h0Mm5kqLbFxMJiUuZhep9CS8HDSxVud
9QGhSDQA+si4+76AK7xR/kjcnpnO0QW0anvAeGR27I8CN6zWDwA8dx3+Ytbc11uHaFTw+LnFsHAR
XwVHiYcl9u2CMmlgVfENC8cllUQIXcIn/k0O4YZSiYCn2ujdr+iUtv/b/Bvi6Rhs4livVt9Z9E+i
7V6UbZYOGa8kdvswR4YPgnjESivNnjBx2VWFF6C3eUSfbt3G2nRHfqMRwDCsdw6cOeeeMWQ0fV0F
m4Q4Sv5Gj5zhkgr1afEoAN5pTTzz6bsQ7abP9Nmvx1eDXm9VGUuqB7xzMP2cezM03GXUcwNpB8tm
J0MnzrMNkrQ6+bVme2fmgnC6SVzwyhnpb+iiTPKbX6PINIHqzyHkUSMl0PLP3Ck+WUo79c438nNh
xU7tO+EJuF651k5cRIbfIO8rNRZ/qZGec8yye/UpTEpzTxbDgrrOPtokCHD0AEccY1f8Cv0yfh91
0YPKExEgWrtUnQdz74/VG7MNYIehNspIeYmj4DZctAJtKQ+dIBSiSXeVfviK96HtVlHlSyc52BWF
5fvVKSxq/bbLgcSzIQu8uX2w5x7u5ZJhMbxR2ngj3ntMsY8LpGgXmKExnPcucruEmaJ+i4s4OArc
6bXfN7O18ai81noKhUciLhWYKw1CzgIQ9JuC6oALui/3PMT9qZPfM4smUEaVvYakBQ9ELqSIbSC7
+qw8BdyzkCCKi//nmm7BY52WV+9j7Ytw2eMey+FC9J6/PTXYrXEaDcH+53nZcBfGo7J18xSbMK6G
4FDYhg2bLh3oDw2Rn/emkLfIYelaJYGvGUmqH2SKffgNZwgtvPL9o3ZddKET4f6XSyZASDYyqrBl
qYe37Ahywcuh5zJIV2m5VBFrF0nKlq4SfLKDAy7WkyJfrnZmeWns/DW8EZzfF4R9A6ggZlgmYqJP
s+G5Fkb6M7VdBSY8ND7SZRjrxspnV/N6NV2b+8OVzbfL2HYMK/z+pGsH9p2Zok4mcwLxSmN+pAV2
oYtBj6dwPhtLnzAzpBV5SAJ7fbLyXwfxh/InXmafKJDzzhASEwxQXs6iTyOMNT3Iu0hsUEsmkqC/
xxT7hm1zzmsBfTqifgP6x2M5vwDU2QjB9j4dquDkFItUp9IuVqRaxp0LI/yVDmu2TmDGCLOzVxZQ
sDzVIKF2ywz3m2/7wsA7e3pwHqZBmY6RfOIBdt1gukqsIkP+6DDqTko3JT3RqUcfenwjzx+7Nspw
YwcXcL9Rg8XQukv/n1Sm7i5nJzo4JZEP9Cu57qlLcJkuVV9YMyxdoEQ1EIJB2fnyuMl4rogxnk4h
ySDlbveCQhAZj3sy7U3pkmKGsnDKWMUxCzuEnRn9eVkdwafUivqjrWyVC2VieY01oARCm8GPRF3m
Pn+0rUiZwph0OaDxW/1IO5yyIS2fvsxngqB+yjeRALc+V/s6bwOnXUOz9kOWbaVJOLYl5jxDRvWU
AeT+hwG/7QCJsYc6/2Ln0J7+9yWTx1XoXljDGbqCPUR0QOCPGuFH+fSHntuzZeLNHnE0ppNx/Qq+
AfIik85w94I0b6I23UaWEPzTRzqow5lmwQIo6L/Z95ar7y6fzkyu4SaUNVXKjmTn61AJghZOVHNX
sTe7GoF9mg+hAynTA+QvBA82LYJ+Q07ps4tdueUl/X//MWIUTOAuKyclYYpiL3jSONH4/ex0cPoJ
eaioMT8zKoqdZmzMbrilSIYQUerGU0E2Q/ZVAhnL4amPzP5zLQ8b0Lsd3uqGiNpUo4mqE0n0uGZl
l3G9MrAAVDVordaDONP2xAyk0xcuqworpQfQ/S/TF1iNaWR5COCGkk5URYZYsBK9HnB/u+V5fhUj
/3h5vLn9rkUghCnhzqgfE/IGKg0EZPYPqYaF8NOEPLE3KWauouQYklL0xffexWCLY2hwDgGIuUwF
/Jy92++4fSzpBdOfMDGLXexaZZb4UeS0TiP4BzMap64uzQQi0ymK99xPHRM9xLsFqaG1aJNHOP8y
h/BU5cffHfYi1GEVui15RTBXFaMaV2kdv5Jkb4vz/2XO3R5w4kOgqTHTk9WsnenUV1g81+beeXU8
prmbnrlX3g8TNZx9E//aNNUAfv0np737WBNa7p9wqYQKdVKVe4/cMeMD54N0i9UXsKZElTOkMb9N
8Aro/0GGxTApFKeLUxkX1ApD2/OJof2LA+tiOW5fMUHvZLUSIsMK8c6J79UFF0nr5cex5tOL/E9Y
t58SbdBMg5rguv+GTT12SN02qvXlYVurezoZvYxLkaPq8OvSM0hKVfplVbN8ErBhPpMb7fOSJZjR
zKbWDN/eH4aDlm2F0zCnuk3Nv55QTXHYn6quYavqpKRpjEM/P8wR6JeMOTI2plrEJTy+ySuyguvH
M3wtSvFMmD0y6pJ2AnHwAlK+gFji4zUCJqQhbwjT6jxtqoTRfbN0JaoBMDfcz0FO+7VJh3OaO89L
0qftz1gHQcQUd4BkKhxTgFX9/C1Uf6+6pVWzfjn6T9W/fFkvk9X801jJkI2TvbA3/FtKW3ethapC
BRyMqjRgLgyGIK3TlqCC1EpSgdzRWaRXmwLEey/Q7oK2f+Uujdp4D6RHuNPiMFsd36nagNvsrFNm
z1RKpB1H5MhFx0HUb413Dix1JkYmv7B/BCPJBQ1zPZ+K09ukire5Ly86NYjuoy8+zcslqD8fuGj7
4wNdRuY3NCFKMhrP1qItdSw93bQ/GRErzWJpCmr1dX+mpriojBNKSEmKhKtMVR0sStCN6q3MmpE8
Khe4ZvPoId8R273WaFVFzGCYs7Dx4Wc4dZA+g1J7wkmjaT3goC6DJxr328lALmmigy+rud+Io6xF
6vs6d6bL3s7cThxv7sOSuZjx5bL+nsD7+Z5+/76k2ILJoxdDAmyPpuOcP31bHdi+gDWDPA7w31Qi
eoTsh8lcbDnoEdy9/faxPik7KBCsMlN/Uj0nl/U1VrwCiqQWWbtZY+Guk1dbVIO6oBDXbT6qvTHU
6pjNx9qh7dnOyhcVeWHRrpNvazXx54+Htwt+TNE8kwT5oMzBVwOhJsO+dZyOKVpGMIzDQXbkVpLu
sle6RfoGWvYngRHI6oKS6Y5PbvFSxbQ52P4qOdKgxKuvbPJHhNkQfmI8NqLcJp3iDclhNXevHmW4
ZjeUdi5BtEjM3FmSc39T9ySqhnF2lsMvVGPfl5o6PtSrHlYFF35XFW9mSc49s3TTl8JGcU0YMRsr
GRQWzItjZ1YHHphBwl4v78a2Nmjgz8qXf+97a61FeNq9QK9ETrstVEvOdfEpeVi7HuH+Bs5kYAeU
L+fRIXlanZtTiXlsxtvXaoNr3jSNaEvfpiEp7QpYDsSLwSYUzFHgrUZeIx2I4Mw0Xh/iXWInecoG
mIHxFekImnXCm3Wu1t8md9GRFMSHTrgUCXFImi1ixX04u+lSHipOC7maQdmxfFG+r7jP1BG1fOZr
TsDljbBHH9G/vjWrjcJPU3GgzgAL28hAM0og7A2wq8mXkG1NC4UUtG7HWa/cDQYOAatt/LpkXUM8
SAK3hAaE+tI/YTROOaeewDH8lXlLGkxyxQmZoL4ga4Ff5hFbiWsAx03n1AScDvY8tOJqheDGkFIe
ZrCyG4MOatIVE0ePSHqElDeAKOv0cUorqYZ+akg2ToFmuDH0RlRTohz88C52BBlr5nzgFTvUY87Y
sKlfq5jdJ10Atds1o7zruubqgcFn656kCoL95o9ZgTEm0m7ZhX9C2XjysYPwBo8x+yDi6ofom9AO
/UZd1Sd41T2f+NRGG9yIK5BTr3GTaB5VjmU6AQuwhfQpWbWePxFuH7ezy9IVjdRKp1xcx2VFwbkL
s8c5xYhwGM5lDcoOXZCE1IBvVk0kvzbs7iDWMDqQGk8fcRCXPWNblfO7qJRpRUC2mEf+PtBSCDAa
schNWNFdtfAhEtMhkVzNympS7Aws168JoV6s5vueeSQP1njRwvGPRZA5U/nU0RfBXoYn0mYyNxiQ
Mqmz7eZ8DpLJzelCs2M80km09uMwpBx/JzSRGOptKUx4STiW7Dxq2AKjksUr12OHmbykqRuJpMZi
rud7/0Qtwysjjbw5e1by396H+7Jzy+SJFqqZsqsbZ3LmbIcQr8g2Qzj82h2B60fYMs81N7KgYFe6
MjtGimlqVTSF+gIV82OOoGS6f7Bu5ia7PwwD95XTEj1DWr8g7dB4dZzbCsRrulqOnscipHJWP1vp
ioc9LD9wV0gnnkigsGZjfWP2NDP9xja7JldLp75NbgMvlFwvfKyGkL2SWRTa6O5oaXYJgDLPltZq
4vkLrCYahVTb0xmn7a8LONCMSvfow12rIs4Hlc9VH4r6H9VL3lUzmnW7H7lD9bS0Zzd02cdNjPsX
uHHBG5w9qvzlbbtnZ3uaOBKT5NL3IoYNcKgdm+9vywTOmwfosdktutUIGQnqeaa19alfOppQ8qBL
vPwTm56ujb15s9PaEahjCoVQ8jJ7PS8MeGrh2vq4j7V8Q9hkaC4QQjCRJ3YmG0AABVPmt2VnqT5Y
i/+bN81m5Kwntm8fmWx0LH3MbtV8+HJDrH6b9YCfgfwqobalZiymw/JnHjRf72vpCdg57oCRqpJK
hXSBqldwTMII8hyVsXOVDH33qR/1avlcmvMf0gxGLU6y0k0gXJ9YNkn8353zwnKgpHUOXz852h6j
LkCnSTVk8TDlspodlX9zoBRgwj0aMhP2+JOZvfb3Ai5hsz5nQNFYTO37V3ID/g541+8TQ4eCm9TS
GjXbnLsENKx8rnd2GEapvHZMYwYUSNQfGNfxW0ey5Y6lBSzwIkKRKPJkI3PxFip9jsJ+j4fUovNq
MwR1xujP3CQv8jN1BTkQzaTuxVaArtSQjpBj+FaUFlWn86JAN2ujdV+kwEeCHX+yYY6d9pQB/QOJ
Rz974MZUpdnMj3Qna50cTOfxGmowqmJfW/KBVG/hp7WbQmfgyOtT7w8iR7kRmIvGMZ/3bfLkRiW5
1UO8IluyE5ctVDatdll03G0JIvPkFXX0F9QxbJgHob44IpRApe9i/0zVwUUHKsZrUSYcmXPdSKr3
5LnsdEWPHgNxJQ1GQW9WOFVRuOTgghQBcxbTMwLFYdtdUVxBQl/DFsX3wSbPcf4lF5pUTbJddtzS
rj+w7ZpXX5TgNmIh00rXGzFA6QX1f9lxutsrV5WJe9ICaBFKp1/DsLe2HFAG6GJZ6oEzGx+RNFEb
o3IIyhOiGDSosstKxKCQo61Q98QP4hnlZJzk5IxygzMmHfTFqAT0uzh5J21FukWMWc5yJluw3sRW
HtJSHizAbQTuPtvmpjiLdWh37Gl6eekmScZfD5ovsRVIhyE/OLEw1lu5waWbu5K/iHy4k5+X4cSv
cmlhspW1Jush1D9bjwe8ARaSBwsXQywmVZUD13MKt6ID86tZAWZlqwEIyl/OwHSbQqIXUDKiO6b0
iGcJ8CohWWjVArxAeA75OVuvtkBccV6kextL6WM6Rn/ICQtajgs1dG1soqhIYDVF8SieRNP+JYgj
In2CcLrTh+Zj+oNEaQi84Vc4HLbHWJUpG6nAPVmRYeXi5l4R0iPRlBJasysb3CbgG2boLkuikK2r
bLZGG9koDfMxqSTF9MyUGKJSc5fjwgILnJP2bOVZuToaS25pL6p9tQO8d4G/3BM7yeINyF5r+yWI
koir1H1ZAU1HhwKwLVjM/Zj/ijE9JcOM4eq6ZPocWqT5Iop8xXFLRIkG4PR3V2rVzwdHRPzxxkR2
6hVO/3QZMLgcAdXoDLKRF+nN5mB+DeE09N+cJxE2X59uPgby/C1Yj1U4UbgCBMI4NpHBT+eEk36F
E7roGyP2hvOot17uv91lRkysWLTqBbfufvHkyz3FWPLuQkFtoamdRnEUjCkGJr5VEPKMdDeoGZ9e
7bH3M9+y5dNpa7p4ELK8Od0oHlgySrgRQqLJ30z4RV40yI5jvZFuyJOtmZ2yiIOS0Dg/wqYE6BjB
6oOBtI6fsDmcJ7KIyFWXRHyYnC0EgYzXRjWMPnb7djArIPcfB/xwSEK5fNbHISwPM/J74gdY9way
tJ4IsW7sC/IWXNUEJj/uJlv31c6Bs6FnavJw6FVpYIQ+WuZfIg9ZQPDB4ulRYLf6kTUHgrxtB0Sc
phOY6n7GBUkF5rP08mwMufEi9IJ4tvTBDPP7BqEdOp/CcNP4niYonJc48Nmjx5gMfLGv7tL9fWhx
DBQN5M1AgS9uygcO27Fkgaa66v63QJUcebtHQifn6+G5wUEdKB2RG5xlgRtUg0LUFI2FvpLxFLcF
J3l6KSSZ08UKS4sCKwJAmLA9eZl8q9zZ3wi/bUy5JLXdoayUedYFfxQXG4ovuci4Xrpupg70vq8Z
l3Nq+QdbEr5YhWGsi6+eG5sfi4iG44EsQA13JUvRpR/9hFNv/BYTJ36vnoPxvqtI7WV/j1hBrMNJ
EEqozsfONKCF1s7sojiJ8571/fDpYZGGOTdh3/QQrdBo6JxvGrx4bVk1EyDLOj+QkyT1lumXrpL2
Xog06bJGR3l5ni1jcMRUui8Ssb0nJEO+6vjo7HiOvcC+iaO4o+1fHu1MNLcFWeN4EhkPs9LtmVjr
cOjnnHehJpKuDUFPNgjY650CkThxqVwAOk3wVgVXmAnVMBNc/TzRTKJ1EhBR9IXLCaoZ/bp+8b6p
FJr+1R79gPWllxybGTSGdN8O7dosqi+UsAy30WeNaFUfis/fPHQuHWEIw0ifGQsi3cM2v10dCAXS
FAQxxOpC+uHnkzuiB2N+DIdWhx7HOUWwtVo8EsJRELvmSdIm1CU3KeZVIUaTYFy5unphHe1+sjKw
N23eoKaQJfgYDMTKGav+ctVSCtj9J2eTxMoAtnr+yySmUrvuLGeCnLMHUQk77IM+CED3dyPCE/ad
ap8NufxPzbkdIXbOOOIFZ2uOud3ZgUtDlcsteygN0ekRWfMf433TNbi9bwc+1N/tv4UuJGn0fTDT
lJteIyMIFXa7BGPtgcS+OBaDcDCcSdKRiHhj3TsneDHxhw1fq8bYLr1DlCQ42r8Y1Msr/AXLtu8T
Wd4/VV+YKhWY4lxBQSKDIEJFTU4niMSNV+pfT/lh/AxKqHrXzy+aQXxk4IZ4HcMtslCn3Zf05Uqm
sYmp7kKtnJddj+dDyKyBnV6MGcLM9dabfToHO6WgXAb5rg+zfet3aiwVqGWYbw+Kk+vv4HUXe+X1
lkTRRYumZ96bmRZIb9NzT99Kzq35nf7kpPXZz1+LP/ahAqj0och7LwnlVl8OivDT0i5NxPtaMNwQ
btSemyjMw2G5jOxRH8b6y0IuTBUkfRUb8erb6x1mYZzbYftxmfg58r0sLkI9dHVavqr1MROB+B2H
F7tRligNodOSQLtA/55vYPykUAwPDvTm/3oiyw7SnE1rouhAJ/OKa0VjdYX/ITu6GFbICLJBrw+l
0Ype5Uf9Gw/u3O1+BQ9Boq9+rst62HP+7dserv5EssVd288A77rKhjCg7ELHARi7f3ZmTU8/fP97
WRMuoCZhxZNTAMi9Yjq0FT3pKgRY6tClnbJF3eQbxWNRt81R6kGHmLgLGQgwH4LibM1KFhmChXHR
5HXUUmsKaY/qt4MxS6i3lOWYh+R0rVhcGgL9AM9Zc9abklSUTYgjM43v9yYQHhUMtjEL+5X66Nl9
NQW2x/uNUz3CnrmOkjoG7OO6F0mDrwranmx4pBMM2bffu1SRQHqTWtpZqnC84SY/2WP39pgVKna7
5Cyw0g5UJ8M+1CTTJ7gtyBPIDAlyFLVCwODQtsS723NM81XinKObm9CNy8goLJBD074zwCCKfNZH
fj9NnppkddGPj7NbnRlEsapHH8sD1RytkMEx5vK/d1VeAsOSiBSMpDENKMLVZfNJdYp1TqKCLJ7o
XDtCUqVZm2LheHHhNpGGbpTNcGfIaM61DvIxprtTq6L1NznG3NDfEPwzwwp81YyQDIXTsqTdhmey
sXstU62vTL+0Cz7OD4lmCWZdSb/9A3M0DkdABekAM5ISDcc1dyTz8Houc1U/9Jv5+NVETFFbMgOa
ywHCEV2ORy0ctvD9JH0hs2e+1mT3Em716DrrvXeQreMB0YcFLKihf5fcTu4QCxvDRuXXq7f4iIVB
1et7uO+hwhsSdk6AbyxamGx/m+gRshsh5a4isyG3u5SNJ8OQM9Q3jNJPBhB8mBB3hwgkEtRcm7h5
uXEE2Vg+czwsJQGWaKB5z1HFWozgqLdcdXcwMKTnQXdzucqWyhioKOnxawC3TJQs+YcHIm8W2LAg
P1rc04mW8yRMlqtpVidPBqvK+JLoW5U5wqeuIMb/UzhAhpSayGc/DhYTleHrAuza1uY9XHEca8Ij
YJUEZx1pQFtWQEkXvIQc6hUZLLD1PYQEdz43KRMGhaRkTVmRINLo66l3lSLEfQgD7G0d0mChEhWw
7N+Kcoo/s+WVYAQZQzue7zRXLKYW97N76OiKz/0GV6tFEY1HgrJFdgYWPwRDTJeBRswdpAx4BpuH
KPlwPo9nPslwvJhrgmnErcFpoWgTBReseAU/EwME3VW0VL4+tdXrBXqMa7fG/NXCVI2wR0gVj172
4881KC+dtS4edPSl/wmhDzizE1IpTxpHwZCzZJa2km0hXFA+1yeXrQRn2VIdsAPF48gUjxq6nY/2
sMUEZiWXMG92eJgRfR8GXxN+yNaGAEtatJJZ/JTuKu47PGye7T2d5VvpF/XthpkPykCDGxfz4Aed
UjB3V3ZQH5hgdtvHJhMAAH/scSaE3FtvqgOoy3Seok6QH7OtPqZYUvLo31JwVwAohPQKnF0EZYp6
cm5zaxKuATSwffRlwnaIONU/tOPD9g5BQeLvZg9mIcNESEM8tA5pw2JJvHa2DoabPwmPJvYii0Bx
HEukVAljjSxaY2cIWgj9jc8kPTv8zhWwzyKUR/sQqs2A7HWrLAtN+wfMjpxiidVG1mMHvmFRltRd
IKDvYnIpFQ277xruaKlbr+EwIl20bOBTDTFYeBP+XvdSBnhsC2TCvG/bEQzuGeVzttONeAH/dAF1
LjeT+1ob6VAxP2J+VY3tuU1e/9oE7G+pmkiabl6pdc312y0flTnczQsSBVsB3F0gDR/tZH/g7+pf
+ylPWXQwy2bymop2pGx/xk6t73yNmzYihI9UaXRkW25bQwDFUSoPKEaBJ4K4GA8qzmG1mrnrm+us
yt5yowN5C95JD9x5uJ7ZnurulMjpIhmrqmOCM5Xi0FGniG/0m6FwW4SfK6iz0Dopl22UhEuK9Kq+
D9/ACu5Z5ukW3REF/KQ+N8e9V8yc2twNPAqpdMCO0FpWbl2biIui5dyW7JqByQ+aEH1nD4j7JAHX
/LX//B45/2kPUXupNJIYr8xjvdEML3IuummAsTTp0w4dmv/Bpgqf4Rt3hJuyo2BP9J921C9j/p2p
ML8QZIwvGd0tNGiD1R/bkYX7vD0iN8T6gblA9zDARxcfVLZvexHR37iBWj2C5p8P/tMrh8jMii3m
A9B26XZCoaXk44gZh1SNvU+BHqXZa+mhaFuyaGEZWm8gjbU48gK7RNILDkxJMOKORq+Ot8t8z5Hx
0js9675WpvwYh06SH6xoMRV2TGH8C1QuRk4i3rdBLC0zf9nXnl/nAes4bNqmeDOvdBx5SNuoFGiM
JWjAwklA+p43cl4lhlsJDL8+OWoi5U94FBlSYa/kyPoHPS977o9hr+VWMHQ7c2Hp4+uEOs9tZ4EX
7i/AdctAvQ0F/wA2I9uCRiKkzPktqNoPFNaxNdeT6T8HvhinCMOU5NvXuXPMozZ7/41TbP8waFsT
35FvRlz5zq1vEF3PWMLJcwC4Fvzu9s1xHOcx5mhJhNvEi9GI+qOnLD0Ej3Pt7EaQ5b0dESVvCs4v
VvtxYxbDvpozXnvBp/EXqqX8UfDu3PnirWKIxM2iYe2lXclcElbKCAwmTSmk6czZ0pP6X0oecwUi
aD9wc1Zht+HK+f0AwiJ/Kcp1R21EBxKIgpczmpnli7ozM5h9U9xg1O8iYAvx2YUCMR7Cb8bd+zRh
KpPT3K2yPxvEoxFM9/mVPN3ckGNBTQrMZ5SVSnRx5kIlYHO8pqARWI9A5Zj183k3MlQHQvpeHj+8
NStDgxPxhkq990eXVskUgBzkm0ax4NVhb3nleaPeG1qfRqvWxRXQFJjzTVjA+1myYCKWIor5z2rq
GPXB2/HxjmgpW0qUUX4cGppi5rYUCNu97K4tULBSYX3KizyZNrzMU8JW3CPyw/flRF5T39VNA6lM
U6MZkTcH4x40jGj5x62toXPBqj97a3orW7qpn2IuG9cnKgFlUmpAe8I17QV2OpMygoj3eHWeaBYM
fF5cwEJMh5y83RB+Nh0drbZegbfPUSCLzFdKeqR4M+bwib2ifXR85+QgjW9eJSp8iZ/Dcw3bbPzF
cpmaZHzNHLGsncA9KgIdolrpIQ6h+6OYprfY5pl0Wvczgv+lDIsf8ebGY0akiqN/Y2IwzYEMeKSB
ReKm+Ji0edo72RgdTf0Ra/QlxNyvXRuSdE+JnqWbJ7tPgCY6Ulf55TSAZ2qhocgVzv+6w2NwEM+G
VAnbGYDIhW3Wt8jICGObyESElpPOESVNtCzXz65a3ODgW/Gr3XzVmTZeMroyRKx7A7qR056VodnZ
WaEnvWFjqp/KUO8I2dH4TxZVCP7RUPi7Nc2+igFVKYf5oqda5ScrPTK97s1fMTZciLMAnB1aytP/
dTK3pcH8wWsdWssjU28UPTDtFZbZEmKpsWUNg/h5eahoYLGrEB6JwOVOO4ReOyjLBbeWMHBG7Tph
PdbD429ozhRT7gYq2HvCBNofxFxYK6YxrOdMv8JLUDlHkN2KuZeluJy2hrWficDunVbH4hmk2nUT
MyyAqqgmciA+RRxqSgpzNtYknj7XuULN5offwabA3tkPIfLDLBjUhdhiwqS0p2IiOLCI7AvRVPii
GpsIcY2mhhbEKf3RgUWBAQIyY9U0qiYX45bejMACMqQ+DZrgRmPRluGPcTm/bHPhLutazzu5QTgW
LDVXWR8TfsE4wfGlXrr2p3Tdo+KP4Awz9g/u8z9tOB8eFbnkSIzDLMqTqEJCeyHWWMcam1/9+oAR
/Z40QmW7LsYqs0vRI1Yhnyx9tqY4SNyzI9pxtx2is5XuzXB/PnUMbJW+i7+Qmj4BMBACcFku7tfo
f0nvDmVPYVq7dc2KT5IenJ55qg1/XD3Fmp7tkkovPinlvlIUA0Xo6YAUO4EfgS2FK864H8eF+EUK
j0CMeNP1kwCm2WT3fGjXu7ONjsc48W5n4B9hnFGW0lEiDu7IlphwuDR+nukd1BQmHA6il3g7oD+r
QTIEQcuc/T8FqsN0MPRiHc/jT6RxDf0ygxAr3aomhRHttf7GWs7ZhYMPwpiXLZaZx1NgPc7i9JCy
5dAMWbKBDMxsaSRtaPImgaDKrUPYy4/CKmbfSlrS2Gkjt4hPi3h9oickBk4pMrYbmCup5wMguDiu
1DdQr8zLjta8bIxfDF5WBUt/HHBEeJVshTYr+B/CGKM693sKrll9mbvV1ZzlW+yi8a4EDkvO4nkE
kz0P0jNn7FqUZcg0k1+/V6zGrJ63ws5GnWNRWn6G/mqPPvLd/0TmI4RVG7uYR8OM8Q5zH/EGLb5K
M0r4xKIawQhTn8sw9zxeo+KOWxKrkM77HsS4c9lco2dTN2Hz52Pd55PEVmMvSEqTRgLhe15SiH6n
527idFsIu0dAhaPnUS5Hw8LUkNLiaEr7YAzwE65Bm3mZsgHQnPbpSJy1NA89qBsik8bOIU82/8Fh
QGOwaw8tVsRUbDzLqoF+uCQemFX4u5oamDOl5pXyOxdfXlFg1keaInON7V3qqYe2usMeXzvIsrgB
EkiDa9+G4J8RsfUkG8xvuHC5KxqEQrY0OI11XYxBo2IGK9l9cghdpG+bWvafIrhc5LuwQjPcuqiV
cfpgMwMesZs+4UJVNBhEqAemfYr74TDFdlvnxDPMX3fX6N/4T/EQIQuYdraiSCQJU2icjNoMmDDu
4vmp298cjY2vcX46aZvu5gPkGqWXBJIA4VHBnysQKb0nvnvz9fFPfh2jH+71Gc6RRoAolYIXFpGP
1fzZHvT8Nhz9lPZIVH8Ap0juD+x/Qxq9koLddsov2vHN4O8toSWKcbHMzaZtcadICbjsf0ZULbhi
d11RbivRuWlOStjJx7y7/pi7jxPN7NarkVPOxtCMCOuYuLy7Y58z1EJNiAEKulImA/Gplap1GKeq
AOZ1qiRb7ZdA877BSm1QRRyi0SkEKlo9sAJptGhpLHw4piyZUWzt0E2SMzXuDXIl60h0Z8qFF7ag
wIVkPnoJBzYZqH29Fg68ElBZNGVAaU2swLHrgC0ymxvUSEnUrw4FLhU/sNFiw3sn9EBIH93ZgFZ3
HyXkXrxtovy1FORLZANDrck1f98mLZsjto7o0//vQ5ufuYJDKgGeAdlQh4OIjEfd+/ZB5vk8pooR
/3Fgr0403xlz0ocO8It+OUDsF3WfAgPgX3643SmAFV/3IvkexDXf2NC/FM9NzNS/licW/BGEbnn7
u/waJ6cZOvBycPMEFg30Kn+LxF2wBSET370PHPNJC98aZ8khoyHKR1tew/HO6mMf9vJkggEC/xXT
UhEyFvgUZ7Sdz6vJ9na0ZaQ6YbhmtyqS6hPbnRS3H46We2Ih9szzGwXo7adhTKZG7vJG9yvn8Hm3
docT7w7neI7Ng5ik8WBpVDfjIR6sV0mkHsdPW5jXJ5UU3DnT8nGDKNrWGcGrGRLeRkujV7gHEO0A
K2ByUmSac/YsrbUZ8euJBp6LQg//Nf1UI8qhGXsvyWP2DpGpL2wd2vBLjtPi4LcGKRD8rWNZ2dUO
nSskbvpF0Q+51Cia6jDlEN6605FVi65MqLXP3ywuZMVfMNg4WThi/3tqwL/W8EjIX1+j2KOiXJTE
YuKpPsuKNeUpyHZJJMig7JzKYQSNcldVng/oJRKnToWGkcVkrpTW1m8xXTPIlLA8adxrH2Jbv9Nz
XvsMCOYMWj4XCph8kF+BeIKZV7oSk374nt1kGxWfasJkYRdvPEZLkiUqiSUc5+a3YGE81gwtWTQU
LgEWK7NVWtzwhXX5vh1ZKYyvPXUceODCOf6lDopJYAVy2PnbcKVqUCSaCxAuw7yE7xXNVxRdjsBp
ewzPrv5eYFvsERlM9IjyU4znVDMDhGCp/H3Ki9qKmFnrsu2agN5eW1P4Z4+NHNpX5H3keZ70/+VV
peFF1tcwqgwO9RYG8bcXNebG6qzIdkmOhQ6yF+Mj56xdZZMm9c8BN+dcmPsO3eGUXQw67V7Nv1dw
4gjNaKf+jsTqnZSAVgleG1//DXR9Q4SflZyieR8b0TFMQuCurujm9h7fGvqNGC0YTZEHsphA8zk8
rxKx5NylP1N6m26Dkt/ubSqwapBQNsSesnS1Mnieec9arfJOnsrivTWhL8wwYNydaByWRFmzDZXs
V0qmerIqpp3PLKU8DDdpV/mLfHoFeOzgYjSAwiBkYHfTQEl2Ntq5A27LzY7zsw7BnxWU7f5KVed4
qT8wfXfYtCjDjGLnEpsbI57Ua3SotHD+vGofszpsf7Ddhv5/MGd9XeNR0i+cm5YM5n4vKfCIHwAl
F4SRBfUfXtToSejHfo0nP3cpXE+BadZEe4dxe3T0kWHVDIE8sRUarpVaMwflxhQ0PV/ZHVfQZr2Y
v6+TcK7LzwuFftdwqtsBZaJymZ31uLCaq4nOwuwVoyck9pH8nBrXb4eFIkIs4UFW+DZoMMN5Vui4
YCwILXD7BHXLZOx23jCewVtxrB2yp2Min600UJF1UQxEKVCrjfZSBlsxVSUXIBUFN7HqC0t7yxUK
782z9gFrkQgcqirOxTiyodHFmCH4QRapyImvGeV6eXEIFexgIvymsXjkorKNonqJbhqZMYHaHtCB
W47X1ucTv8ZGzfL+YSvOmttEGah1ApaeeTbYV1SjXG46/uomJ04TzGTksXbPfGtXKkb9bchfVCs9
vgai11EzKKKGjoiSkIquxC3d5TUFnAfq5D6pLcLd2iHOTrHNTplwy7YnM85gkRBohdu8D3Zd0KCx
qe4W66MMvqbIeCwr0MUJyZLpjvPOm+5N+YcEOq+wqwG/PwICBfXRyLk/Y1Bp1CPz63uWhcKih4BZ
RnAG/YoHwL9SrbaXVnimeGgmzK2T22q5GlnwU6HfQByKEyWMLTfRpe2QTIOKh+/NYO9u5NYc9+5M
RHfEMsJJQsZ8h9qz5ZtotgtTiUi/cH6LXVCzHYedevcDX7vpxgZ6vCBZQE1gE0g9/yMlT125wiqZ
QVgPUzt830m4a2b/xIqk0go8OI3VDdwcpQ7V1S/E/zeAXReJvP2rH6+NFXlvAPmvkwDvCQyU8WUw
rH4uCNvHSIF/Xdcc0NPmk62hSXuMYxnSoLwsp6pGvLnn92oMghYhV8zpDsX9YajQfZfQQAgxnCfy
tRXBZ5CXTgzWIl5kyp7bxqo1UG3foxIANQr+FcM9lkHoSJsY+HFffVaa/8mtdj/346aXxnNe8taq
uLMLWx731cS6qZC79iPylFwKXM//vjhCW9f64Po+9io8rCR30q9k+ZOKq3Yf27NsyxY5Wa+7EeEf
iMv3bC+jTYTjGBEvy6rFgt01d3qsJqLyDcL76ISbfXXSWWLgW13CIiPmOa3tF1HY7anv0a3wKLC7
kKzvwItkZDdYjtV2iXV7GwsqiZa52GikWJdTdUe2nQHn7eCjUmguAsgcHhxSvGzA+gF1EbWjDnOW
EB6xCj96ApG1Ff7e/yCCnSUVonLUjo1TZhd7bXgGWzIQVRhyCG7/sjfgKiZxIosYTcikncxPKjuZ
d5bIDAgVvghRPsE32KDXPvTJb8FS0UbBDZwq+4D33Md99AkCIhOee/k498qPfjLpsUt6aBIh5uBD
W0PlHS5vLxcLmmB6QEhJxi24UNembaWD0PxMTuDg3bPXq6tgibJBr2VKF14Smaffe+fH5+x/+oEO
0mHWvGl/iFBqox4nXSK3GqFsbFUnfqn8ye37DCwWxgFlwhP9sVNTvFv41PnVcLjy7Rxmon7XG05P
mfNHKiu9RSWvXfzc/JZh+9CIc3vUvSwrk5XmDz0qC2CYOiSGAUVRjm7xDpDiiyTsgMGY1RroeZPa
crwjFLc2JKznRzcjE1Y+QPuit5LTDloYLghhKlnvz6Vl+pHnhp0PAF0oWXHJ3/L9ZkJSOZrdzPUo
dzO+jcjvswCum/ZNnq5wey6kvtLhO2mZI/X5hnBMNFtDy2tjEOntOLgfBbqTx17mscQuIEX5orFl
UNSYGi4fX0qdylw0xpAhbTkStCCgCi+jkdHLu1jSzXh5eUrXXCGJi3rwmsiLgo70aHyQQfShZVej
nUhJR5Yig3vOPnhIJMsnY4ruUjTpg5eDkhvfEWcv2QaOsUNCTMBp30ta+ULgTbLe2hud+I0XJ6L7
fxBYWkGv+/3eSKB1o1S+4kE9dSqsO4fr24uebnUgkYOq9ruW6rE+g5wDaayzy4E8Nc/3ZeZQj3Li
ZaFAd0E9zl+iRbcWLj3/Mi9D5+4+SNuUBjE4Q9Z+bAloFoOZtz0JlDv6IneuPwYnFv1NrZQBUtrn
GBf5oJPsaqplp0TqC4IFRV8q+vpZ7fwTI6AR1mdsWHTEHPKUg5MEMTFZYcU3fyB2HfMAYhf8P59m
jUpSTctCy1S9MGMdqOHmwjiTdVBIYZED9b0bZCHffoI5ooQPAy0RUbk/DuATmwz8hmbEDSxYPi97
s84axKS3BjtKiHoRMocPJrqx0hbMQf66VbsOczjRLJeK4C07hMP3wOOLlNftBetP9YxDgOR/JDaU
dJkNVbO1Byn90zo678JkHPa5eajwTZy1O6bqS1MwkgtHAxHAKyhbYtmO2tza0aL3WDtAx5h+p8R4
OUHlrg1V5FOj4bmYr8jlV56ApY5sv9rATkqycoPePr1o0nAl9Fd9qOAfrF6VahjuNitVvv1bbVAL
uoiRqTgM78PJqOmFkilsLkK3hthj45wczoOOqMGOWVcvEMmFCJREAOD+u5eORc743+Xj2jfYBTNt
xUM+RbPWcnpyY7M9/aGDWSeHGLFl0UV7l/1X4+OnARYiNuIy9QEeGjuQToqHJIFgukD7wfoxCldJ
+6+wHWj8Yt0PKZg9zPgAn8ATdAxV9rlOMuPvuiHraXlxkvOJfHKjw9xl9iMYkxN5Z1sQ9rWcUQ9W
7lTSqPYtaX/cfx83CSncAk6wS6DvPqhzgRBKUENSYTsbFUqacH6ipSZ2xaYezmf17PcnL95bYlp7
2vxQLdR0JUDurqd9Jf6FicLqWlBxJZZibW3XOLWYnkKMBVNOTz/+Ym0j8stOSANwnrCJIug7I2NR
3Gz58cWChFovo5l0DSacykOyNITReJRa7EVo3rgrMnyglkVmrbgXk46CFoNzgvZextfMuM8X2mjI
Q1ERKYfHrdk6G2ktHK8wA/f7ETtVLXPascTEND3gOpLhI9TVaGGp50307Roh+RQO7t0+Ia8udCw9
DE1Q6qqkslAtyM6FHQmd25CeRtPgSvpRhLNS/jkotAQbGGJosjZCo9w/PhcUYJjrHqnc9PejjhfI
HkxgKMSnkYVrr+zgRZrGCeNALTPC3iD6vMxHTSFOzE0SiaAy7jVhNrIB07B2GmRcpHIpXPchKHuI
8+lUFv2ooDvrrGd2DQfeg6nfqnSsgjHNXUD/0hgPd9zAw8LeoG+TozsrWxc/PC5RtNPUJmUu+Zta
UviLHNktv10YWTetshyhqnZCItA1Tkt3u1vX3M2WQp86BPTN/3x8If84T+tV0+MJgQteuiWfn/63
zydT3fWHAbopuZvnGJZa6Icm185tarSFQp17y4d7Eu0hl/jAJYHCk52FaRFkJucl6PtKJPIhDIdi
lAQDUrEQI9tEWQN0W3JW6xuDDsiAoiJh8XKa6y0AZlXkppwP417iAQwfX4jWrWYF0dwmEdezCEnR
BDKg/RB9LB1BUiuRzH932Y38JrpaubbicO6GTDSFg9wLKuajeRDD1Y/IuFsVU7doj/ZlAgOhC/i7
dotwrwgVUlPDnVyOtivED9wvctlGCWROCS4jxQkj3jJfXXZuSzJBLM9F298vG+DAKb1/dNRqpOro
ScWSp6DtDZSuJL0M12vIH7vpj5YzZZgmVuBlBN2isumEjBLFPOrp/SMq0ymwRANV1nzeS/+1y/fE
JSef/Sx5htej93Gf9EDopT3Hicp46Crp6REa5MEvJA44HyKKCFSD9SnabkzhurpLIjujV2R+y9sx
4iqDYHnmMo8KYnGd51PY7Crj1XjKaBy2ikVppKQdAiAATFpJ8hr6azYRMccR1nq26OzMQYuZeVn1
zkn4prQWrGk8AvvxDzi6RlFOpKY9KSpWMejvEaJDKjVPxYlz2jD/HsXou3zY2RGT2WmUZxLB74KE
gJqBMB0RmsCLKhGfwrLb7yh9L5YT5uFJtLC8hMTxN4UbltN/PmoEoWQq57bSvk1afHHHZTR6oihJ
o/dtgTQJ9Y5gIdxTdV6NdeudRffEmO5+TiY6sKqciz/fYWJK+sVw8htYSjBLQutvGfAhCHC50zhO
nCDDwSHpKFCkslGc0OkBPGoIhbDO6Ws+Wer+700A8Lmo0ptWenI5TDEOOQOO4uMsk43IhiqpwaRU
Q/akNITkht7eSRY3iKMf3jtBqhN1pTOA4eqOe54b3pm8VaSPSlfs49rvR+aDuqC/U2tEnVtgzzp4
H6vl1Mj9GlsT1GAsE5bWaK9NuND6Gc8ECf6U0jSQuEAiyvKN9uytUOPOKWksP7dNiIoru4DN+8bu
yMEuPyJ7vdw/x022xJ+tSzF4F3swiebrJgCWGjphP/JySe+9Q1j4E0CXGWifoiEp0iPO/7u5MCHQ
vFruwjcvUupNkM33MYS2EssWvef7XnDBr4BjOn7+kpfLlRaNn6Xs8ipiZYPRskYALaEp4ikLbd4l
a8OwsFqaKdHMBd1etmYz5j1W2xF+MxvYlCS5jsAA4DvbFD+IEb3JwN/heRguTnZV+xmVAUTXKpys
NbHa7i+xXIrRZjqMiOJziJOXdTQvdUCLKxAPXLJtjA2rUbC4cUSIYjkBKeN0mkllHDvxfxJmkEFm
t5kLJTVFXFiKJeVzcJqDr5UIBJSfqUMx5VGnzKJi/KAi1zPD0HIS3qX27dHfmE/H2FedFKzMyF5S
6K/3lO75uoMiDMzmzaw26f3ga/j2V5g6vakHLohMw3yx0t6TkdVsG6kXmbYJFYsRTolTWR/K9x+v
phOBdeMLMT0gRcrRELsj08QcdU6rJqcZyvZswHCqzfOCwAaaZ222AChYP/cyIGyCqygy0nj0f72n
5IpsfNJeuoI9uYXS9gYve2uyRRemEdyPMVwxPXVNQBh7bQKPIgplsszJsSqAnjqAfhIjiEBL2Zl3
CKvvUM0JQxZhb/aTbmxiPtGIY/NLUquvoca4ado24TkVbF9LFSf6MiLq/1ZKvcMs1efnpI1pLteb
QulTjve6EI5b5NzFkfdlusyLcZu0joJxPpnqKeG8m8vC9q69mRiEdFh7hdr1YZP9Jw+p7Tov9nc7
uavoe6jrqw4ckB79B732V0OwzWOGBxk5FmCOPD6/mAmPv7g4/CFd04yUF3DRBecV9v28N6oIdSsF
eloln6ymX3j0ET2FLfjLyHaadSbPbJsqpNE2IL7sZDSOnU3G4OtCoFfDEjJeOUdMHgfE+TmZIr0j
QBzhJRMFKsqY7Gwyi+0Voep+BWmtLMWnPiu5fMw6ISAlnMapSRCaE4l8lupqe3ulGiS7BnTMiqIC
kge7Aslxm93lS7J13GmuSmFXaAdeiDP1clQvg0NJXy47JC/WUxtSpOKI+Fz2Z1N20L/WuckO9IM2
gC4brURUXcDzlKCcONO1/BAwJ7VYkqyhNiQKkAvQ8JVooMvrAYV73CWSbotxhcIEyMjLHT9i/CKU
Xx+65ahoaXosDvJR48qvs4MKe2z7iMdxnPXWLLVyX+0z3XY7qSRdxmY8yA1oCWXEOtsBSlYNrxaX
G8vK8mOHIUZ5S5OhdQ1oZ4ttB/XZd8c7bZLZxrNwLFMj6IpIptQIMBFhl62WpcXoMiDy0aJ6HqNc
2eLA+4INLJ8njq37gELK1RZPSRYwMNPPm+7Z1pv/SgZTpOXsyiCrMwLojCzxSu8JmJy+q7dqBoCc
1pwJN9dFm9cQZWuRlHUyPWKKp5d5Q8qiVBzP2DDF8qwDhX/ONLXnOfws9nJ3afR75jzl1hfYoGYX
SXY2paeqTxewg/sROSRe0s4n93KQ/Mvg4p2An97wESRLaDWEsY58cVzxveOliSToovrAN4FPtvVR
fU1s7L+MekdjUpTSAN/loYQdblX8EZyq4/b+WaLkA/SduR9QdFAodaYgWx2PbHwPAfkTVIVcTtOY
KDgU0wmvrnN3dLIyMQ5Wi0lurWoL6UdmKsLQMH/y2q+HB7QHximxMMaGR1JLZPhiS9jur1e7UVKi
+H01MUI8spzb5url+M2QAvOcCrrssiRQuXWNK7EitEFhQ6m5RKe6dA3tXBhLBhL9FtZt95doI3Ek
5p646yDkGFDbvblLnx7mUCe2gvDkAtg5imSLzIurx0aVCEtGlm7FV5we/3PhVqeOZQmgVYcK3IEg
O6KE+XuIAqBJYZHRtF+Lj0shECrU9joTE3OD+eOzUjbWJZxW+yFRnllz6Ko0fSw6mWmq+shfq+gR
riw6DXGtMnhvk4o2ClsHRzwf90jLDzmDhd60XHA1LIgf9IMAwK+gJCgTSR8TxkPKAGAiqRSnCdwB
3z/vTIgr/v2ZVh6xUFSoZibwywpYTrRhc9t/iFwniyKuTyoL6lqmBb7rTzebi4QyThTLT8vf09Wk
jL0IACWHehM4WBhygeF87rG6g5G/VNQDr+LGA9wLRvGYikhKEkzvm+EdYCc9NcUND7XdsHJWANk/
bqGXlu2k2mmMKPADoSRm+cyTXUs2LJYL7d+G3NhBkTNK5GmaAftIhAN4T66lM6rgLhDurhA0P5QW
Vh4D8Us9fRYFnHihaS2Mg75eWImvZPeCdJnN3fpNh/vZIBbN3daXsBju6Xm0p2o/oKd2mYPi4VmH
FQ9C5ggqFJanwMYRejKIlDji00RmglNN/8iUHRazCrQQZ7r9RjnfIeD9AtU+RmYhJRZ6G0GHNiUB
EWgS4iFDFMTBQp2wiZL+/zklOPIkvEqiLCobrInMoarnagJPyzq8NS8t37ixDzJ6/YqSYtJOtK2S
CoQuGr9FE5n3WhYiPDczTMp0iC8ZSGR7oAawitgYAhN6iYIJe/SKFvObrDbgWKEyAeaN2vNeYDow
9T/vB7ZbsNHVw0VAgtx4ZSOMPAdOMkhMaYQJQ97quCKI5MH4Bmx5c3YA4qarAMALr4PAdOB1tRkh
9F+s1RoVRTQamtDZkP8WXfKcNZ08FiMeFN2e67b7JpX0TMrADQOzAfsBRIAgDKvWyAR/92jk3SAN
g9V7PoJ+sjF6dHHTn1JuyV7NJQrM7I42nC7Nd10gVlXI29Q4edQqEvmT/WCHDvwA2ZTban9ZzVM6
3VH+W5KLqlMhbo1BHQF8CavwqkFm/aPJqwUuKAS1sUQsDEl6JgExXcKfnkzjZAQfxGETzJOoQb29
cwoxnVWBHfDq+yQwitFUO2UazYGyfONRk/raGwXsRFjz6EOETQkoQaEypP9NKcIRzDEIfO8Gu+8z
blkyQXc6cpTPTKWST4J0IWdrKdMEtyK/Dadc8PYTCHhv1zonCpEtdoYQf384qGoVqMnH/sALuX30
qyS0MBw/TkjYNHnrPNSeW5CaWWhWmC1d1OMq5S75y8JUqGU8h84I355OykcL0yNxMSaK8kHghCn7
8LRPqFfyj2eo8G5QJsLUTefxCOPkJHLABN2OM275GmqKWyFJGQZUryFWEPvZv4obXFvINZiifiIx
GxTfiqWhJtarufM13Q73F20ATcT+z1bpnXCgDMZMAxMd+2FmCJDur4P7rIhd8n5omQ4WAy5eSgi1
5nPn9qq6raP08pzNixIYv44U9A5YjZM1/80UYaf402EUMgyg+XlpfyGh5BKHIxLys3iI6U2buwgD
a1RgkPbGsPzjmvJyLTZDsDCLYBAp14wuATA8wQ4kHYJw1l0cUsdm3u/VPejgf495qJtGUwTo0L/N
fg5V3/kNWDNR4MEFI/QnvNInZSoe5oR7wh/ELQ0tcidHsRDGRz1713GABxsfSbReRa8Qxwm7czTs
Gohs4gxD0vCLbTHg973aN3yYP5EfDalLDhCk+T9LX3mUMgEZUmvvMwOelx2ahUze6c0WJ2KmMlvJ
wFxk+KW7jsIPw9L0yOXi48CPkBQP6Hzz19TtgUWSVRT26t3MQgnTbgDwXiDKkWqGVNqoMg59duGN
7p0Jb1KmQS+BqLpGSZPOa7zDJvwxmHb0Eq+WRuMwPf1s1qQAKKwSODuGukPAU6kQrM3i4yJ6Uj4R
Q5qmuwMVs9HlcAgHMi4ZQWi0sSuCkv6u9i1Gw/J0PSBj3dFe03TMn+w9ee+V0OSRFbHYsOfdlDP7
Hg+OVmyxcKx1yi3ELFPBe3jRbWi/Hex8uqkhAIdxsi9KgIy1LakJGNG7zUFziwKFHNOPLaUlahB9
B+DQo3l4VAM6LgoxHLN4hRa8r3/5PBX8UfTR95NfMv8LV4g7x1cax2aC+a6D7vBQcqpuAooXrMZ/
11j8R8jFCUOW14vKq+8oqPStxHGxQeHtR/+cTb/MBQKPRG9bjKpC918Ct+vkrcTQfqo5yNHzengh
npGdwYf5MQtG2g3kO2iQ90rtf3ECIzK40teYmwjnx7fQ9vCApS6j1qConUb7IN+5sd/pD7+rvtsS
TIpqA7aH/ySveSXbShQY5rrZqUCoLb4zSyj6xyyfELAYrA5yrQS3IAn2s6STkVMCd/ilS4dbBnQK
uJqsKN+wdXk3RoBnWuJvlL4Jb5qw8W464E1Z98VtcwZU4XhykgQnL0YBTNyRau+oCDglD+IkR+nS
A7BcDuuT/bta5fw8P0jUYfBJ6PM16qYq2SfVOppYW8uo8db+qLQBf5/54V/VB/BGqKd/PKOovIiU
+IjAJdg4DdhhflfOw0AQNB4fgJzfBNKbhnTYA04xYDUuWqd1mIsPilYJhy+bn5XhmdclLC7NLXKO
DSs3l1wcGNzR2jvdmBj5OWiRWmtIp+kOcm6AVX9aUqFEd4fGu9o0LTILDajntExxRnzHu9QZ/ASS
gvgUBWyyoLJp0+Be8MOR6V7QkSHDDw3i7fXfjdu+I0UlOSmC3NKcDshYex5JnCk+1rT2BJspzbVf
x9IYX1fFzfmqO0T9HBhASl4fCPe6agDPjhG5e7nMVWzN3yVEm0rF8p3NaMLm368ozAB6Y0c5tSzD
J56U5HPuIyPtiB1Z0BJpmzlrESKGebuDKuRMuP0ddCwWeL127MRai4iKM53SR3++ZOE3PUlo9fRs
w9/Bg5JVnedCPjsurvujdYQvQhC+oFwdec2S0Gq0H9jWfmhb/K1o2ly8sl6SZ86sDNsiMqf9Aw72
Y2hMo8W1JWtnI4sfSTtxnqPonWrFR4b+pM/EGOuPTW4qRj0aPDkwEt5P+kF71rBJ/id1m7hXN9cP
zjU5jq3/vI4Xq55Vfh85kS3uZsMjkx6FnT2AN0nxUlmeG/51JcIJTZDcAd0aCyHQt1P8P3Z4IiG+
1uDs5vOFgbUjslKrhGhe6ELmahfS1r6BRNlHAP87BAK7xA5ZtZWRxl54pudtLPJTKCFRqGbYyJ8w
aQz0zIbRXtw8z1eopdAMJ9ZmXjnMjb/3ZKU+LsixxJEqPytHfWb7y95nGFrgAgPDsreKwg0eF1XR
JcutwhggOlNBrnvnklFtmpjpxM4MSBPODBEwfP9jUvRHfm6rhEadp0dNGD4OUOYXgQ3HJlFRxzkL
TvHUi7GWZDd3qV6ia+w4LmLL/KBFsxYZcqbK/VeW1TK5Qss93oGtrDspARi5g6KsVakk7neO0aXJ
ri3Z7HBht0qhBaqnADaPw7m0EYO7SnDXS9suQleDD6Bfmj7GsT0R4S/Y/ZMCpjZuo72jMsg4ZCsd
P9MneTcsP92pwKPNJZep2DWUXhGWVU8bchCmsGmVwfFAPIdOJNNaOJH3BejLyfRJfFr0FyySxIk7
ymMNqHQoJd1E6+eVRxBy6UhVKz1aYhbPrjWyBCG7W9AcRGwXvza0bd8LYxprlWDGzp0L1C+aCyTZ
gsEXOQACE1yGR6rqAG4lQmPrUjvuVkFfol2WYl/UU851ZyDvuegz9CBaYEUl66OmbxAdjJqme1f+
aWi/ZTBEpmktNShZxvqVvJWAvKmO9yNG4ZSOmtGxjEN6zkkWrxVPtFH+zpdB3NH8NUosI+a4wUdW
efMPLH4CmP/Vle++s8hv9fOedzzVM93KZXgIqWIPDxJMhGqQ7ZfUa2YI0HbCCSi3GRd6hlUj+MKL
YRZ26Wr07HmfFZ9PB9MMee/KmYomXLv/4Iot2uNGw6uOuF/H+IVQafeunkbE2JEMGlxA9S/jN3XO
qH7HpblcJLCxaMzpu/86aicq+ZhZamn79wHmVw9KZvSmeRXr8+4x9AGANTUKD31B6qw0Oi5/L1GC
Hbg+zfYIh8x/BNAbP36kyhPadJIOafdkydNmwTI2mARgtOR8B2eXzed+ophvAOHYJ8GtQgvVW1BV
rD6JfLYCMcxPyJ04aKGMrNzBU0a8XPjnseHcUOCPEE1IXnM5t03j/uIEAcg0gc7Z2wrcY6dfcNua
Gaxz1zlsAqW1ihtuZbIYPDrCpEtrilvwyUCpE8OWH6jgQZkM4KS+tuTp4D65DdO1j7c17Bu01Qq9
8SK5/c3pnOQ96Wb4+NTI5Vdj7n+4+H79K1az3OC4fsNQMULAPoj4fE3CMHIAqfcLvQHv+w9uXPv0
pTOog6YcWPN13tI4PSsZclgXPUZ4K9uHEZCHaLRTOa0TQHrt3uKl6rQh1Tz5CcCfxkGniYduRsaF
Gr4/AUU5nxj3vAKQEzYHNz5ZuF1icIoMld5iTBeoySETjKBB1LkQtlNrZG7nuNuBK9nTIL+fufTi
xIXmv/3PHCPi1aOgLY4FvRjz084zbTHKFFOanJMBjcpDebG5O/4WcoUO1FdNf65oqwEygNA5LPPx
S0dVB2teDSBj6PG0WmO6OH9rwBYmFO98fqGE+rpk5Yt/LvUUfbN/rntvcR1o3IvUFI7glGKvZDZY
4SnE0UkipX+D0zu75JI/vEnqEtkv/BkTZbkDwl4qwSelzi95FxlEaBMvxtx32glCT7bToyVgK0eR
3PRTsJBGAFfK0/awtIRCC4HmkSa8EU25aSgqcIpwRCkLQvA7x1Wmqa922EwKdvD2T55OY5aySFfz
sIa/7eOEySR+M7gnzNrNAMZGAmB0OOyMLNNcLwlmif9m2GKglVdOYWR+sNbYf2zKotlx8lMBMQoy
AyD/d1QuVUf3rK/IwLWOfgxPx5d78cJjS6D+FYMQdWCL8Y9X6cMBEyfC+YRBTaBBFUHvtmEu6G4j
zCZQ9Gi4Q1E6pQB3VAfL/3kHWiGOiC2udJKfaG49vIHXuoeQDo1AGWA7pn+kfGkwROQgJeRtYS3K
+EB4NlUBavM9Z7uEC9KEvkxHrtBzCpqS/K/NZSq1C96euF48sb3tKldV/F6grT+Nx1m5ViMsVNOu
SCr6KlUeTIUNoFW/EyKRT7gCFw820niN1MA8m7RFh9qkWt9SZmaHNGbItlk8l8g/F6THzS5RkymI
XJuKmFKYIQSxIKXzgk9Jqjn3EL2qJlBT9X6gAit7iBctKbN3Yn2o0cTVvLnu7D4qhydkzcvkcx3e
2NGkgLe88eMhTlShjj/884PEHuTICnnetuk3YC5o1uK9WsfiILwQ+Kj939NwTyyzxoT9sQ9jxl76
BJuKAVa56j6et8c3PZFPFlEnBB/4iiYabIceRZq/1NHG3KqX4e0vYfNBjmoL2xFNgVMj+YlbCzmE
oFUcnTXX/xVOgEj/zXwCKxfQNKzqufi1PgbRAZVRngxFXMlNxTBLLycJ95203aLkIbhLG8tBpqLz
WUPCiBdNFfY71PLuzQPdfCu8dQ9BRwJlMnd4sFcrUBJJY2/oR1EGaSiXk8WivWGe4JTTXhhHKe+M
6c+TpbCZucZSuiBGA5KUNNPfQw1/UQdEB4BLrG+Zm13KqPzaY14+g7kovgMP0u+HDkTwFYlLnCt3
20I0KzaS3U0AmZBuXmpWl4ghKNoGjIS7qEBUhIJyPas8/oDC+DxBwY/O4kREASic5lB3J/YoavhV
/Lpy0vKDDgrvmZ10oE/hmgKPSux57FwpIGyRg81qyXCF7uh/2vxWOiwC9wM4aK+0rQABMXdtSywN
Bo70XbvrMfipiKoZFppKY0q7fi4ICLrDor/cQuVYTjLGBmcKUnDQPHpDaE0yEU5K2bw3Y2b9X+9Z
eTzL/69P1lQDeikzqtsFFEnrilkr2i0SA53GGEP9Gxg2/uWvNWfQM6YK1wRFQdR0Zp8m6E/MKlcV
oNP/1oLmhk3I633qCnHO3bD43jrhfUxx873wICXwTXDaDCX06xN4SHI7Jszd58wxygqDf/k+kjN1
RlMyyG6DTeQM3JLOjJeuLFiSDRytPnchGgI9cIJZeExpc8J9VlhNZSQeHoUw0kZEW6ld40ugAH48
LOFGv4O6oGR+pBxl5KRkfUvJp5XTKcAd9GbFzFaz/Fds6ovw358A/GVmId581dHs/UY5sBgmP435
eZj/QpjJjUI3ebBMdHnznfTbQJhFHzqvQ8kojg0S5FyMrefnyz4BKbto7clo9eUPozV3n6h+50yS
mpw2OqblPrK40ek7atxkg+wfg5yCfInmxTSbCgAq7N/glR3lPnCSlSfgUxLiCO+i3Ah6JO96WHIU
DMuPd9nDCXK7TUCLpw5vdD/uHGSXgc7tRqoxFTfp8PNSAfkwLusc/Cd58f/iwPNUP4CTeLrfK5BP
o86gEsKVe36S0sR0+sKIJHRHzk96fr9tOoZIjhNR5+KZ+JeIun6AkbfWTgb4sPd2Iij8UJKTGK2f
3wSJNPsQazWgI3OKpTskRaRq/WZJE9AnHko/ERFv+u7IgbGqCL73QPEia0WALdvASAAuuDkdYrJq
N4r9XAykRPdJRRcXbYGO7zLzGH/JuFxthK+fLB+46G7Htm7munWGZG+BUCFYC4p8tmsZf1alHfzS
HbllxmzBx4h7585157ucjPW/TqWd/uRQsPZToCJqhVD+9Q+AqPgiDmSxNkTFFmngvYSDHKAeOh3E
F89Mw5v/C03BnOrZ0YI8tScrBsy1eF/EokL+d6UBRPyChsSfxin9AElEoPsSmeY1+ZhSIVnD94un
GkZXk2DjxHy1lUt/QujzeUGU0iWKj1lPdyuOVmLQAL1k7qc12m7n2qQtdLaTqjXOn25+Lk91uBR1
rovqOoQ/tqxQQAK32ZpFKG44Zgw+47xuV/lzwMe1/ME4HQ4omclU6e2JFjw0S55d0lAOmQbBf4a5
Q7dVcskYkJO0z95DkCw7HCX1y32OiXbJvhlk3wt+CSJCo7kzgUA7GJyJmjTPpHUPgLdUOBraL13k
qN3GCjFPWnESB5WTgweaeXIylzIGXGdO5t+RqQoHEN5Pp0i1Re+0o6ohFrQFq3lqD6FTPcv8lprD
qj9meqHAaPqjM9yFSBdaz+Ia3HQEGkKe1i1aTbfSrLpcEDJ/V912IRiv3FctNz3EqOSKnNO2y/X+
l85km2iWNzQyLazGoYx6kwKENVZmns39+HSKLzTlqsT45xE6cMZB3kTehvIC+CDkLB83IYypKnxi
r/fa0L5s9lSWFVWzP32WeU5aIAXPHPmR7xxAFoKdDM9dAuee2mhGLi+H5yJTel5AvfVZiN6TsCg7
NIuTVb2KpH7ymLxPkjQ2xdAP6EppV8ONXWZdiEfn1mpCtRe0i8orBOY4YBWsL6ZE2a4TKbhoDw47
nMoSN29Nr5PFOi1dC61k5eng8Zet72vtKSeCv5TXEpTHNLiSH/bbBhWYl3gS444e3y/k2F55mGIW
6rcOnRWD2jS0P+EnrOx5wwPTgLVKgDhq1f9pC706nz2aDS42WdBMcbNQqqrmeLUD2FHPlY1HHXNZ
yjJxIIosaOKS6iOqRvnvsXrwCZM4iN51MJAqrtAg0Ch3xQRDuCOlgpmPRotD7CUKaxO6kdMyXWgs
ZaOb6/HvHN0bI+mWEUUTHhoCYMyNS9QLwxeV4KLVprbwG00w7S+ttJ5QvINVDa+E0SBKspdof1W8
pOKlRcqxqnzo7DhF81JcDcUU1OqKecysE6jTX9v4N8ev2ze7705dd0eeYMroaZfMc+gLNqdcN0Oh
22Yki8EIOa5mBhgXtLz8fveBCRadbtycoiuyOHF9kc0if6t3I/qHxdw6/kzs4YNQfGWH+OIshCMh
4fSGYdbWgETkCru//M0U9cvbh721VgRvJWGeSylDt9u7FicTzt28yrkFiYH4v4weuNCzO+EXlo/c
yR6Rgy4KJJWD2JRr4Rbtto8remA2RzzGHq2zBhY9EsZf5wWEfcviKmYpjFdpYJNFKjHQRRsREzVf
YqmZios9TFjGSBYVMIfzAHDeSui70YXcV7Kg7ICY90XIy7om7B5zcImQ2mKV5ngIY/zEKLthEsqT
hW5hSDrCv4/dVv9+YL5RYHz8mkOL2mIb3Sit2GWoxLGRofazfH2eFdHBirEm8TdFa4oucjCzQS8L
69qDftS7vVlmxpLEgKX6uF8x3i6zuG8Lu4UTmoE7FgK7fSr+eXKhJihgXrB5IWDj+R1LU7Eawpch
40UUmC75tzhdbpkaH7NH5KhU9a/K26yafAA1p2YaiTsGiD5DPenFurBb0FgW4p6TvYIFMDsKPmdq
SDlLbS933RjykdbDScxmSdyF/XG5reNBqGVBBbzUgoTpNhx55pXOItZfAnqs/amXv581dE7oKV6n
z3+UWSUrq7ZrSuTga8/Yi59XQpvjZ1YK6p3D+Z7an5ISalEJYmLf9EX6TFOJ5E4c+YaR1mXo8EmS
JudM61w5vdsNcSCvSs8GseYG3O+lcicwwwCDDIbYSXDLDRGc2170/rLqFTNAm+SAW/9bBrR0027O
FBRQwY/+ii1ojJIGGb4dO+1bH8BJqYyilcK+7pnzMoEE3Z/YX/OP0bfpS4AFBkvXjvSIwJ+xrHDZ
ojiYuRUxpRCCjVDlkja+Xvz2PkX+mjbQzPC8lhxPzA7W1g52a/Q5ms1VRiS9BRJKj+EAKMHBgUbS
ZN0kE/xeCoqv+cRioKRkluptFThgJb5QlboAfqksYtw9QS47OEV9yzeEWwNjJ15Fx+uvr5jVJTtL
0P3xjdMY4mOZIgQi9ouiDQuqfICEOQXbBYqy4BumrT52mDMte/h0ORlO6sCU643QzIW2T3lBBG9T
FPmQuV6Grzt7o4Z3YLUmeIUukAdzoloxMAEMjvfMJbakpNK7PbtwJfPoYucmKdvGJkuWTwXQHrT3
A+fvgre7MtWmh4Ne8/7hdjtVIHItXkYJhtVQkUYEiKpdr/CqXM+pZUOsm10kBTGpbUjLARUAueDC
MfZTeLFTXLzumjWAF33J3IB2sLvrWta1uTvBIRLkOoTusjmi/6ifQPnROvbfZWx/Siw42RWyMOhw
4pMUX52ZN2HIuNHaLGg4iVuif0/g6Mk+y2ztuUKa5YOY4AlB36+y6WXa6d3HFUYbDs1GlHDjgqhb
6KOO1GS+g9e2z1Taa2z5t4a7sn5GqBece+HYhyp+C2VAyuT5NurZE2Nbr5fKRR0Pkoj789cF2kc7
DpCzUBEcgRjENFN60rDfBjyL0WVofihspEByp8UmDL5vZyRUBXY0fVLuGh+pawfI6Vg/scjaAhjk
zD0XCNFX2OLubCz/AsmMgHiLxqV7S94VEmNJ80HSvtvOF8GgUbCmz73CKxjvpkdxRwMQjtFQGxSI
dFBxiGviJ9EaoYqLVsETQz7xiMdEjgAr7w4tmeOCh0SUL4VS41LfzcNSfnEgD6oIPzeO8ji7/lPc
PbMWSW7caz/bp8qJeTnLJyQoLBUuhGLx9P2jZvhLe5rSPRYhzXAzyj9i0fejIEi0XyaBEYLkWOyE
6pg/B6Vmt8JNT+B3eIrPFOHrx7M7sEWophkhlNFk92uqevB8DVpxtLxR5fzSnO4rwsejNsPLbOsE
wSZ9TgX+RH9L6aLJ/FCgufNQa6+b/ZpgjelTkbGrDtLM6M73VI+3LTK4nsApwj9ezg3/64KdQiZ0
s3kko+FfvcB4ypD1FOEP8YFol7mUZJ4pKAem44lYLpoPVCtm8Qy5lSKaZxb69pkd8tBxcEgesygg
5NdeLmFaaSwbM0Ns/SHt3Bbng5LRmGUHS4GNL8i84f99FCazOofVrLocBfptHKdtjd4crp7SGZEW
Uo5oWHLaVn+g4U/H8jjeEdCMn0bJW8Zg12WtC56IlyoTslvMEGOY79J4fXK4sPj7yrizU72xPazC
7fRoIhWCrceVI01a2sPuN68fBsokdlP7ZfHTaPpjh+zqHog/P2DryiEnt0nLKrQoA8990KBggOqe
vNzzh7rgGVSm/h65IN+n2gxf0lMM7f+yBJRTLhhfI3LCHG4BRJRoWej3bVevj/5zfGm/VtT7osgK
TFTekI9hC2uq6CdFL+M4VqiouQ2DLJKHlpaEfCWWjpgdPjW/1UqMLE889+IdKpHCygsXc1bRuHga
/kNEMN5pmNol1hA8YzFwvTVnHOr4HlGBh9Ag6m0sP8/9yAklEOYK6+kLsw61k+yhg1nlhQfTzHw6
xQHtUOeGhXaFqjz0B8uIRW/g3UvDz2MjL9NJ5lW30fow3SNmcRVvK+90G0zhE7XqJMUNla8RpvCb
F5cAcLY8MstTdwWLJ3ipDyrRmsyzmhX9Ii10x8CwvnMCRdwuXrY9LSd7KVrSj6lODLonL+8unbpM
8WV29vKsEho64HGCurZBNfWTD4r5SbIbKYl4D4PzxPAO4WwbwGppM2XqniNkm7XUEmLvd6NVdNNF
o/00HZf2ck8ppYcNchhGqGiB8L7lW7DhNDbV7woy4zX5Ul+FmV8VLtzM00KhRX9RwLOSaZvSM0Wv
n/eBIqE5XgtoM2zyDcy/0pbtOmkGLZ1UhR3OShZUtrAwVXvPWZ4AT8NnLRsNmLMsYO2QYkHG/VeB
N0a4i4bNL5U1MpjyqmdEgj/hLlZ3hgTXq7qm/G28DjB5DVhvNYasElD1DuXWU8eeuSAd8blwnYCn
QK+D9lU9sOZOY8ySFSa+6QkkKqVcThEDRAEKGDOkZAr//Igb9BEk+lCeyxaaR1lpHM8zAFTaH71Z
DIshGD9H+OPZa6+lbFCGiTwVYO7luj0+tYBZZwme/ygqxVFUqeLoOZDOB0RohCYPcpU895mWjoXO
YYLomxsx6UFrXbdv07KNBdj9qEjILYB4XDlC5PPEyapvKVvVzT1tzD76NGOOzpsR/LNeGP7i6TKi
of7CBkl67TQMsFfPyX0V7a+aztzhqb3/vE6xoUAgxZJcwJPvTFfKwj0hPVH8GUA2SDWszOCyA1Dk
BNwP1QJSeWN3UouyUNm1KiumvB9/aColiGl9PKOzdiDzECQ+0DD+vbl5C/nxSEDJGebjKlFig4W2
QsZkmcTiSXCzh1QoYU0ilAIoRVqDlWefWVbzsIz6PQmIuMaUDgbSwhTUXBere+QvfmRfJwS3c97V
inLOoXD5k/cWERFd8Po1bVrq28ZZS+pV1RoQ3USe8sWyIJny3nMmrFxmeqKreVdfzmDyy8cSlzcA
7wIqlZsNDdJQX/2kn7IWn9gNmGI3/4LkbacWJNJOKVBoNFWsrthEpSBC7azYZIVPXpL0ilCdafoW
ZzoAkTyy+GtauXMJRroKlpAfx+Y/wnUMGYei72hqSBFogogrqZRRRPL6cXIJUJYCqRgZEV4Gi2qE
e65xQTCeE/97pTN0ktru5ostQkd5KnN5MWZq3JmsIuJYDiX27/a6qou2dmhTg5Otq405ByqpVzmL
BXOT9GszNzplJ+XhxAjzoZe2F9DQNLfxAcXHAgTeO8jDBt0bsErbYNLi3GrxW+9CvKKzLp2RGx71
9q4/ljyQwCgxJeoU4dyzRiqGDply5MRTZJY4AtmBgWpwtZnvbejJaibS8/6kReqW2p1BzlFxcbSu
fHH4Mq97qiDWSlxI6HxoynZkP+1tvhwsObe3ilQDSY2nzYHCrMYgktiRuISt46psf1HFXrUtOaed
kn3oiRBl+TXG7lTPy0Q3hRQcAfvbuNu8zPUa0qDwvawfCM2P8dQLlDQ/BwyRnYl/uwDOix5j78pj
2aOCTXOHt0SvDN6w7IyFIIjw8gR0d7aosV+eWs/+/U1/4Xx8l4DVkNHrJ+9AMoozaSFxU1ms8dY0
jQJElbFSBPcC/xSu+2vSqmELlbelk0zsMlmuNV3xfTvxUpbu17kVEOwvJoW2HslRCwNH8l9vNs5S
Ao2gf9TKRydsmjDtN/PxR3lV+O+0/vNs20LZhhSDE323ZtuVj1k1QF9vnvRsu+AUUvtrfkEwjkmY
5iGocNB3tQVO2joctKZNQiz/WCicwWfyD+vTORA4DapZe5PyDP2Ay88GAq7Kyd7DRReJ4VpaCaua
9SA6x0pGDrvPYUYUCfNfzp/+ZaChulbh1Atm8yiwVz0+RKqgFCUbvwtP5lYjdz5RZer820NjfUqX
tUdWtMrxVp0UzwLdswrHoPQacND7sEpr1r7u0zMyESrbHFONYMqEyYr6daC3hIbNhlwJ/QopQOEJ
OjGFeA5eP3MBxjsX3OaS63P54CbaSNaT5FrPnGIH2F2h7SN9KFsy9KB+OXDRSIG+SAf+Gqe2WmxZ
4H8F8dXvDE4AetmJQeybk0h1slbQosVpuUhW7Cnq61MBrOCsApl2iXaiN7pCzwnQZgDAg5hn3Mrb
nvs7djCk8Y+4Pr64mG8ei04LKwHVSi21rX9J4EfwzgFceaQEn2+ZuMJVQ0DYw2TQBuD8EPpnq2uZ
lVRtLXEZDCkWHNVnxlieQES2uIYQpM8+oM/5orqPgQ/D6XHvGHUzfHvl75ln53IMfWKm2bdPDM6x
1jgKBlBh+FdcF9lTsj0/KXRw4dObL68Lhtx8hwGYmhz4Q+Go3IAOkQkaFaze2ejePtl9TTbGxBEf
BkIfhbf+WK/+9vJt1YaCqokdb6RakuXXNRpcvosppNnvtpYsW9YHvFX2YIZ4oqkku4ahLPM/iUcr
hpSpyLhA4VbB1klJHke/MTC1L7G6H3Cf2Wqz56v8s4fxhXcHk9PIUsE8wLQc12sOpwGgpp+0qNco
2UQZKtnbcWsK3siIA8crlbawq8MwcGEvmnhbVHK+zg5DEuRcuqrOp5Og2w6xRet+3rvrxTc0bSe9
3EUQtPb7uI3HAAasiwV2Lbh6j8T9qQznxBHnCL/vKU9U/Xtnfu8hV9KuKyWBUE+1Zm3VU5/8+CHU
AintJkK+n4IbA2nr4dxX0MzSxj3cSkjrphAHsYWmWQwCnK5MUg2YOFm92uaPlnMT7YcI5OHU0cEU
/dzLVTgXR9hurXhNQVelkho/pPdl3P+1bVfRh5AycS8YnXKz4QEI7dbcQAvKnNa4f8Da9WXkX9bi
fkT6rAXxKy2B1Eno3Ggab7Nj6UeV2lhEIfkjLf5MZaiRg6n3CZWvnsagbP/JdGniOpAPDAtMrz4Q
tid3FHXJTRQUuvY5aTbWTzNhf7NwZCaDLAaunIBVAxbM9w6czRqgP/MGIenx3nlul0bqd8xBzgeW
BNwoaiGotSdJqMrrUufkhks7xEYbEDAviTJ1ux6Os1+UgvZ1FtdiLzNprh2JSYOml//fxXIqspun
dZUXvcEbLoxHai23riyqhRlbFZq/JRTuRNfNZg84evEI8jRyU1QK7Cm7u18xFb4cQeeuVpI8vMwO
IXq56ljTfJsIg4ElOIjks6uB1SJtpp1xUulLexZFKHzeX7vrbRtYx0emXU6woaCly6k6rNXpdoI0
4CAe1zbCvKoptzGcFquP0LXmrIkqWhRCP/PgiL0aMBEMlS0psQ3iVSDF+CaizzqPQs5FLvFbTvYx
y2X70EqYjLebx4HqHq2S3aAPU5WCteBJGx+qLE5P81bt1K63nejy7GX3wxStYBGmOkAW+XF5Wz4T
EQGADTUIHX6wkpXzowk8drhHH16XaBTRLEnI7xCxcT1vlcs+wZxwa+n9u0MBQMsttjTNMyVfD6zp
F2Z/qjJG0zpLDmj0XJ83qT4dmT6BoKmOuocBeVDs9fGQvG5V80lRgkQZScJkvKevmBs9TPdjuUDZ
704RZ1F5grUX2bhrN/iQPwbMEGY7S9tMUzittlD46xuuMa7rfuUQ/XKmYnNZsUVTirmNLQBQsUPK
4rp30C5NT13sCrl0yiBcXyBjqe4ZBQcBkvQcTFSFmXat/+155Slj78PAR/WFrhd+z/WlWCguVkDJ
mtxn6Fh8l3IzzIM1fn7D07HX8MFNVmviY1LZlQvFyvkeOzWfgmilF/74N/iXLP00BBo8v0rQQs21
vfutHwHqM2ozXSpF4QLlXG2X2HYVUHlAIbLYR78gGsqc/jtqY8vrGvS4hqGvKNKt3KdwhGnqlID+
kAWjCJyeb3UHCLu/4WBvhHWCUVRXxE4PfrxoTpppYoqStJikAwqKV4rFKTGYxvL5B2oQXnp7QiF5
OMMTkXRavnmrZONjiPsKje2VJkWCa55h4MAin6feF06r0ThSsFy1nEDaoBcxc8uipGkk8Kl1AIqk
ebYyNJgA/lACh3mg8CI5EiE1Tr9hzNT6HUMdXp/LpMpnzUk/BW/eqTdC3am/n3ItY59iHY2zk22i
SPo1lRR8IAdmuHLVvV5phNvAPXIvPj2gew6HuUwx81CdsYqtZr3l/KTXmnOpZTLZw1suHy1wT+Eu
9AdQVVzOW2WvT9BZvOrSUSnun4+onStkJZaVTtNOQ0B/fQVU8WnlWeeapQE3WlW//ovsuCsnWJAV
Id+OfajHOFAKwO5zPJZOz9SUHsKVFEO8MaN1vtNFxJ96Yiy9Lyky+esFds9FJ1NSbd3NRWOg9nch
0vLpf6Q9UMdL8U4HnGMG7FsRlokiitPUgk3tiBtu9C/0GuZ3bHlELuPaIDHvum1jLOmUzfcs9r/J
5owN7j4WfbZSP3kQNnUc2og4Q1m7qZ/ggwwBjRfNOxP6gHMhgMMk9RiSkPexWgbqBS7A6lk9Oz5f
8Eu8rQ0hh0Woew0tnYFsAd3YbhTm++wibjOACzmotYPaLOJA5ot5Xr3RNA4oqy8P0yqUnn6WoFck
0HVhkwW1+imWSMmow3C01vfR2tSxzl9EqU1wmw6wqlibCwFdm4MJ40ULRIuHd2CfA0SliccMGzL1
fGvBpgnWyJW0+kIgaDn7McE9IkKjyhmu2IUS6IoW9LB4DZNJtIm8wcms1Ws3mOzpGbC3xeuMEtkx
qATplsBOiJ8ocaANK5cRiwtA0tW89D56HXSYtTu2R3FA3KkosMQiPYIB1wYXhOJyI277Zf8Saoi0
dbX1i6q8a73CAmMYRd16WjHTE1rUxY3c7rLnlVY9F+v1JKyrw9XEz1IsHcZSkQkazlAQNo8vvDGR
z1bkrl/q6hAbRESHSSp31989lBFTQdLk27IeNlOuAkLLBkuWv7FX0Js/CSsdfS6g09KWdTtTBLWw
JYJpAppzQPqKKyGZMHlm2fqZFMSYKnbZ8wsoZ0hAk650y/7Qnt4kukr8Y12cDM6PrrnHf35RDncW
L1VelzNzLMAqIXGN0ybV2amkWblCqrNeE5sDZECjxc9RmeAqez62JLnuKGnOOGmEk2UvRdt6I8uT
v9wXcx32GQMI/3csXaf9zI7Oq8PERaWpF8D4YnJ3iWUFLziNz9URZR6uTkq3LKFjZJyJpvWJ97r7
uMMi+p3OQrsWqIE6/IsZ+sCiFFEJY421fwI5d9Z6ZZ9N4SFG2SH+jg9i4xDIgPQFSEDDUTXxOR4H
yLU27+seMgrE12o8TvM56sxcL95kr97YVOMY3MHrbY5QkgjxFI3bcJUZNzd1+SpcklNRNnqEFCJ/
FxUbb/dJndslEcMdDYervhZCT4QWsy7Ap7n9rkrBA5bYHa/ABd7RBfcHaVw5c/YY+hOvU1T6CWRy
FitAMLeQ+f48z1sLKwDAm7xGz83ROuWyP+94L4dkuV/m/G4t2ErWlAPopewlXHB2Gq6edMs/2kRN
LFYkBLm/qQZnlJ5SPb11nakIe7ZGviDESonARf1ujrSpmyd8XndGaloQnFTzuaZLgyLpGyDHEYE8
W6KC31Vq0wE0ZQAHNAEjDEwuDV9Df0QMyg0NICdpPGniPYRUv3GHBb0EhIKkvXmliTWSqD9xWpjU
ejRwy450Mw68dP9cRiTCjz86t4UjeGk+wpks7Jy19KUi9MrpbXCXioLp/7R2sL+3/Pv4SIMhaCX7
WV3jRE3m6OajvxKtBZixgNwnDAF1DGTZMjZIEjg/NaCUseusKtt3WBxMz8Xe7HDvJNySdkZv2l1I
af0pWl9pRPn2is9C2ZWYwtKrkt2nv9mK9+LSgOFgsyIki/XneMlMGPEpn8x17MmTO+R252iQ0pCn
9zGD6xy6K6QZezBewTFsIwtlkO23xhsirZ9lU9eK8LhrH3wf6O67gnVb9cnNs17olSAdw1hezels
tu7Ag0m/RFhsGJmJTTyNylKati4tmuWWWJf/RDRcayx1bGIlFMfjotdNrtLy/9UnXjS1DVItBitO
xLy6xRglrNBZv+DGOoyHfk2A+aN+bVNQ/kBXp9lGaxX4p/JdALWts8CJD2uzn61skANsyAi6lrkW
u/PxHbp2bfza8ut2+YBVsItV76hUJTkInZK2p5g78wJyvP6hVZ7mBDGBwtgE3KRUUwdkQ0uUvsg1
5I2h9D+pSnd3rn033ado+6Bbg+ajZVrrn9xjYNzfPzsj6pAqalP9swnqIEff12Mcapx7oOL9TP+t
51FeCd/1AMowtvM8wEZVEPNH1EHTs7M3ZsdpM9rrsrs5RbC8wbcSNrFusRwe84mMEfCEaFksalBu
4xG4/rcvPxvxMBpyffLMJGvrTaqrXAjyWNs5LjXzs1EpVBc9dOqjrH5YY/BOTLvXCH+7FZt9rZTm
z5ufcPiwcMjFiGgAAxNh+nDz74empUGSVZ121F2Sdg51yLf3jLTwgYnOTA3l78q72gWLyjCJDSn0
doFVc2iBHrORhpgd2SrqpU4NSbxTOqp7ak+R7bpQO8VY5WA7d5N6NQlUZZocxY4kAx0Zp9hi52po
CvSSZjwUfgC5V8j82M0yNnqgrcAxOWNzeS/tnF+aZuDwaE6YXfO1OI5p1HWe3scsRbySYr4hUs9l
105qfpsiLm0BBmYqHxv8SfPmbmL7+TQ7xLufB7b/IAu1ccEupcpJz0ROrpsan5RRRe5R+RrId+GW
nV4pJm/a1NnkzCC2ggqfWffk5NZ/TOK7geGDk5gBhDdeEm2l5Hj83QJTWwjbiw71gzRegV0GbGtN
DtVJpxZ76VDkWmAkBxgqndRUvwGp6hBWDx7gHam/ILAePUvrJ8uje9w1hsi8uHySKEWiQh7bhMch
up062CraF0wwallF4aLRKO3e4ZVzQ2seFSDzFZrD4SJ24xwQ5mrcwv7DzK09DP+f9lLrAzPYXbJp
+yuZ7ESPkU8h8p8itS0kK2pKyLAEJYtWUdM9lsKHXaFTZ3fBG6QIn6s9MV36khloSp8Bo3Uq3ct3
W4oullssTTPZ7JcMPLG+geR3jlj0sJqaes5IrXp1z/K2x8P7YlO+h4ntVpulQJYgQUfcdzVTY3it
+vB9pLlZG8EyV7b/xUqHsDPWO1nZoK2jNxUMgRlP4iiWLfbIt3udBgiU6heLReXO/iUEUOHwsAfv
YVTHRaTB/qgcwWxSiP2EYPLaqlqlmpUrsap8ChQ5k/54LkHSOC5JVQDd+nbPT7dPhlvn3AGlQbSX
07i3xLwWAKrEmQIynm8Glm0gLkWoS0P0rfZcwWXWUN5LfySNgrBeIeSKIiG8st20P0owIDuN0koA
W61hUs7fuTxdl1p7cvFsCe3OaXjqffzMohtvnQyfnUpkJKXi7CjnRyDtmtOWXZqckj/RtUJVa94n
LkV1B0asuQ5BiC385z+gsfcRGIfhH2UsUPk4WYna1p69RsTPI2/vh1COCXqu6UZcYqNo6OEDRcbo
Y2EjYIq5eYTlSkEF1L66t087Je8MGPU+vZSNcLwSvIbOI57IpsaCT/IGa2cCl0hXdDrvGy2SAujj
B3s5XSjozn03dnCDgiNrFKQa7akaAj1dlHBO4rz2vTUrBZEcBNl4c5BeSfkfNPrjbo4HGeaXVrHl
LMGFt7GvlHB05ok1bi4KpteeZrsUe/nCiBVeG16h4TQiMp+IXhjTd0GSmzqU6ODJvmE8u6pd20nw
oJC/3BzmqCRSSQs/g+PANSWNSMmAm5jHy1YxskUkZDaK0SxGWDXGemO6GppoUarelOTAjj6tJXw/
wyRSlvf3N9sfgBxBLadJCYQKFRkpmEQQoLcIRJYwSS27PTZMo8T4666ebgVKivHtff4vBTDuAA68
oUhLObvZ2c/hxMmOgDOyrmPU+brWYAxIoN6h+wWnIQ7+rg9r2jROhVYPlz/hn/YR75frMquIlnXM
b7DrRtHZYQeh5EqOUf9iYfs7b8PZYv8F5DlNyimvahviiMJqwPSagS8uQxq5VHTdWYQgdqQ0gRaJ
5xQF5TCfut316oARvc0bwixq51CzSft/13x+rW5sUKubYfLHVYFg6VwIluODeghvgAqsAp9PUqqJ
gL5pfwqz6UWbKaQWSq5RhYHSZ8zBhgtuE5gFBiDVWYyFXN04GxTtUOtnkGh/si6zdl1dp7m1CJO9
b+av/XGZliI8jM8hl8jQdJGlikD9aM5GI6qRH3BQhtIFLrzMaxmoO4GmHAwREcT1BqNceEbsW99L
WAk2eFZCoHe4MB4w6Im3MxOZTmXmjI0YES6iHj3DFkDYg0de1vNmA5umjtGZpPYYFwq9YLxpK0BL
fS/5D/XtQSKl1enupK6Ghk2X0YpV6MDUYawq5PME8lHHsEXJp+h8jGJ8deLez2Tnaprsux5I7VkY
15Jo5xbqGNOdUVNG8HXSjDt15PyjViTvoATm0UmYIvD/9ELSqsLQHXbgRI/zIHtrDjU2kY3hXGr4
meHP7CwWa1e+sZ8Ds8ZSG9Gam4LQqUlPUXV5RNZwx8jhLLE6V55dAwuiMPaIpoVjlES8UXYncHJR
s5soQ0hZjFtEYctsWha0LjLr3eTwZ92gPzuoL/GllnJtbsI2Rmu53F0u4gdcAtwCM3hJ9mS20F/N
t9oJQg4uyEze5VLVm0pe2GFe2AtsI0O5WXpoYT0xgIpo4gE1PfEes8K4rB/ZGs1gFG3MH7hmmwWL
3BuT6JWQ9rMSpt5VVmTxDVrTlrm3PaZz7yTddfEPL+p3R6yP19+sjpIzalqJh/FtiSrpLvwJ4ZR0
BYzD7QwGQfS08RFDxscXTPZSAFKaWXiRqeb2f11Wjf109x/Uk7WzA8++qOInJlaYyff3YUeN3lNI
J51bpRzM1/tFIwYzRMvM37VegfuJ81s34RUVi4NUX2nCctPZMBkR3mamlYab97B/MbC+s1oolJuW
ANwkPu5+T7uI8V8cg5zAE640tJElpJ9BrNeervR1vGBuiwkWw6GOpS8cwXJom/bzh8cfJM0pA+kq
4rHfhB4bWq+8/PQ9jdtq5rao3KQ0fVDbgZfniiH3Df9ZPxdylbdvkBBjdNKFMeyFrrDeT+5zghI/
oiwsdkHy1zRCaRAMAh7OsMv6gb7JcgcqAT/ShMYCOqC10uCZkKJO/75uQcccMwyQonmheB353ML8
qPsVr9/yDHUu1KDzdp8J4aPv6uWDj39xMtgLRofOILM/+QJ5ZPhijFIL4EG4NFjVhKFREdrVT+XM
7VQqJcEPTu7Nhcg/b1UFasdgH8KZ+qL2iQXT/U4/LE97OyD+v4zYxCJrGQSfDSHM9e8t5sW9SodS
Bqa2zo0459qxRCrRyV1WrIX96UDu4N5L3q4/tOy7sl/FCrwnx+eANpK3slEVKqy+Czm4lk+NXWbi
124GtceeB1koQZRoqa2V43YH7HUHrtBmRgJygOkjeRqkezyZzw6QJ9WDOjDMgPqWAi90aFR86V4x
NAG8hxxwa9v5ti5xxol8hDOL3SKI4M75vj4pX1kOIkdbQLaPoDtdrJDdeXiECuPIDHuoYqPZk3aA
1fw1Vj3EGKKb0AYVTzARAljiBcBQpICLid3OCrI9CF5q0HcTuhp1j6a+/yGqEw4jCqNBopK2XC5h
a9D2mabgLcHynO4t5mQJeTKKJl3Y+/MhlcIL5uto5UJSLPiDKl3uKIph6a1C1W5GgpD5ZvlrBgfP
b2o3EB7I8v489+JWf1ESlbAyOkvHgF86MlgukxsCeSYZiV5UUqwZCOvmefrkBuChr60c+joimfU5
YbHOsUzU4ykhqFQua56eQlQarhBtLuWtexLFM6L0hyAIO5/421HMTCi8+c7/7W2085uIqiByYQ6k
bw8SIuGuQPdOUhHqOppBPS/wlX4m1DhjdEnKQib3iM4BzA+p76I3b5x/+rySAfaqbQAzvQ4caVPJ
egTTh2Etg4ODHhUWtHhhapbZnzwVp29a8WzfQpTWKdV/CKUb2e5dtSKgH8yIt/NVp5LZ2WarG5Ag
hVaSgGMUAk3b2LBnQ8f/Jj3VjSI2zaSqvJfy0vVvLNjUAJ/4z/Rnt+JUFsthdwulkhqRVYbGl4sE
V1KLb/c24//ayBvSX8HRMov93rjaObRO5szv7LjczQ3+mcqEXe+qdClMdscyPzH3N3c0RQXkvKhX
xvL+xEFBCpmz3mkY9rw0TCatLttSVCnGozAytOla1O+pkCSpGTA0xEDkCEZLe0SOCo2f0twtJITn
U6Rai9Qt9PQAvPTPg9R8erfWePU8mmIeild6K9n76UowrozQdvVjX9uZtoPb9eqxCmmZr/+GRo9n
EKXk1j3DRYAKDUJjoR2admYsWV53jS3Wg8D2yF7B1u6ogUb3RLzHVhQqEVkg7WePu/VqZIAT/zQG
Nx0wfpYSixLILlODwBXHGiWi7q3bUej2YPzHplig/CacHmX0w1gU+AIk6xh5cZrLqxoZIEaLecXY
7b7s84lLmDPda05p6iXcAolC2ZMfQD65JNZAOD0bBj06x0DCwnQe8FYmQ3r8If+uAKFVmriRPGn5
tbSvGI3eX88zc7+fYH+Al0pNLWXyGD0Wd3z5TTspyNTQ9txvKiRDVR+758ic6AtTnHBbkYj2t2yP
+G2/RmsuITgv91GI8HZ7s0pB+FXnEDdEIUocIcsbiM86Ypilvy+dJOUoYtmijsD4/si4eo2ZfjYZ
OB1Yv9d9tSd9ddYevcbB8VfS6stDhLiLSlLh/RjzGmxoG/q3zxyQvFFfTyE1Ld8ovI+H2yZ9mhlG
1mXJMgLLU5SMoTatVWCiuyTH9G+ykbzJkBYQz/n6nUCcIt+dQ5opafpvwZUCLryMD6DQOfdMGeAa
Imd6WQJauKa5S/r0Q09/U3F26hv+2YMXRVxaWLp5AFJmeM35h7jzhxEE3eEdO7gNmeGBXz5+BEhY
qD97U8MjcWg9A+0s7O1Q0fCKNmdKt++jRbq6B/44WYzOUNBY8tsoN7CsiURadjXFwxaIwhtQK7vz
W7q+AE+wTg2Di9WZMgAu4KXqJxDPCh60qAFSAJt+JB+16j+im4CQnWjncLpRGWHz7/Qv/2YX66Wc
jYxydcOk8TO9gX0GdRtX48g9+RavGo9ruSPFSmEWce1Pnuc7KhQ0wph+Pnt/61tDh/UmREvtfaKj
l4yEc8SICh4RTc1sOXbYe4fpYjBOZYJF2J7VA+2Yi03LHjuSt4yg5vKjr/TLGQH6f+Mh/2pwiMDb
30YSkv1Y9ytmUN5COFpxk05v7Mds0rBF0Y4E1PbBeSuPxRn0Fic3e7XGL9EZG5Fo2UpC7U14F3DX
0qCz0uLe0KTIZRL6EQUON4/IZ3v4HXmmo9xiPw/8vFHmMKZq0LJFLdwQMKFUfOpBAS6d3WdkruPc
ajABIE6fAcVgGuUoFb9h4clXDDZmeqZ1s6yGIqyPF04V5Dg6jJXoPgwtONc8NL2ptZ0AJd1Q40ZS
/VNFLQVUVCvaNrXOglUz1wYHkpyJnibScdtKhVPUtkUbC9CnzkHlPMtTYYark8wIuDxsDkvbGIhf
wH6RKsECQVCf8gvRM7wUqTXGQthUvBbj43a6kh/4y9anj8gcHw4opZVZ0SRtK0/oDIQMAhKlJHqB
rAtNIw2/ogglJa0cls3sbxjCJiuqpKvJaG4zYFIy3idoVFboWpSN2lk3bTOq8WPJ16m1L+Uv/FTs
3KA6QCY7ah3Xhn4H1fPztR0x72z/SfOuNPGZGICRm2yGAVKRLGKA+2rkM0BiDKbvKFm6QvZbIw8k
rMfCOLEoNB21u5VY1cWkpaTT4bKxo8vS1LRI53cKsQ7fK6WikW1TKCiXjst+QVIY02g2vJJC5XyP
u069q2qbq09YtdSNo0paU0nvO6AHV+5C/YRwIFZFHan807yVD4NdWV2DtNffExDqzvcaiow8ZeBw
SFeFfzNFfCRil6sA8iaLyLj0w68rlQya8JWX7RAuLvA8Z1NYtXe+mWg8FPwfs9VrRE2rwPUQ6uEO
P+4Y4OU8TMpDip065xMSZUpxONksfULz7JYvPa5CyV0tVvp63RAJET2lyKtTyGPVy68VVVvp1Odh
LW6/Cvfo+8u/NphV7fEnsVU61RBUHaTGZrIC0GYJ6cjTMTQdFKN5eOOMgkHORV6l18PCnpRxxseg
KA2Bh8ADslkCrKkXQdGyAZQsv0UAURUogRsAEOQgSFN9/yXLouRvWyqJjYjwR0emXryPgEH88Btg
G+GV+UPPSwFz+UtUD3Z6vEXLHCJEGNga7fMpd8z3AZ618KCmkcPcu3modwW5AyTQKG1OMSNcO8ue
Td2E2BoAUAyUalOCEESmlotZO0NgH9WUu5OxLP6w0YwWXk4i5NFp0XLuCOKJJrVokIDmjtRklbT7
nkAeeDu5Nuewk+A8Iq8/Lt9uiTMidp8ml1nPhWaoEuLuqCt7/bqQKtgyo+btJiEY8hwF/yfC7PZC
DB7z8spxKijBv3QU/6dbmZVwVjOw43tQ/gZeQSRhLPgdy4XKUWulFZDJlELigKV1s4ONo+JGaXGr
zZTVkRD+KGTmZqdrevdp/+GYlUQHb47j5ob+iHWc0Z21UsuUgYLHgoEpS7rJHgx8wA6sojRchnTQ
7NsiCGwlLMv2AR51rGLxE+ZIaF4XG9fU4r67ksNoETY1LURGezX/C7MLRxhZJIkyr5eflEGm7GMT
oLO8rhB00T86D3hAg6AB4uCHKbHs7N+kAGK/ntrWdf9pIMXQR2wasMhLybLKcuLCFqx4II0BRk1P
FWeE+BnC7/mn82W5IFzTxDKZxIF0q08Xjvgeppp31JaG46uB/ppcRBw9l1arAzbgXc6L8W44DfMK
LVKNNVQ9WTS9Kir5xlLFq1guFgErOonc0WdKmiClV5YtZVeIzfKzGCuTbEXHe09oYC0OtufBGLof
dRnytBdQ/kr1aGe/c73oh1NcptwfaVG1r4iYRENb4X1ju5ZH28DKMscDJHCd7tReMByQAsYKoXwg
uEUD2oYvHV1e1kT4TqV+awqRT+GYgwlVbgYO4thiigXKgdqugZ9C/O63Jr8mZJi0Asp2lwOfenu5
NCombEckSeEt6lNrHDswCerx8tWgEWbAXcBb9EqWUU/Tk/Ugr1pEbH+9UBT/jw5KHIYl9IabrFcE
/njm0SKgf4kK36/+fVtDUoqp866NeJjjSnMISLJM4AiU7IFPrw8nKZ7Ukhtssvxq/R3qb/GGvloI
dO7DaBTpEZh8pE97vkYwZD9/xsnO9IQoRckLSj1C9KbYEmlqwppcPb4BCGl+zYfqY37/n3dsPyQA
NGEtuLhPToSGGj5/ANmfumBGnlBJW2HjZD0/mWWMzjwOyppeAuDnVqxQev0DOD3QhoyJpXTSI0Sz
FHq4wjmUKQjUrC2EyFJUjhh75SSEnvyXEVDcE9K+2iL57g6X60l4/4yav9Msg0EzBd7+Jdx57v6i
SoRfQI7nZ5tshkMoKaMwDAS+ZJMlVzCtYu6AGEfQBuQOjFNKZaMxClOkvce14h0Ta5zU1YafriGX
yUXe5FS7c7zhcryHu4Sb0i8l2FURLnCLnFCSAqplbbESyc8nDUEfpBiWEv/oKMOhBYAMthnhsvrx
sgkIIR+stJ/0jN3AqlpCKtzpN4LW46oUSw/XXkoydcVCb9ybOxFFcNjMiigfL6Ed+6e9aqL/IsOj
ooTJTxJ3D6vzk7bYfA/2NrHms2QChm22TIl+gnRvFGkOb0TYeOZjOWFRexG+XeRlg8xCOT2Rm1JE
Awql6qUyQLaa4q3Dl8GDlgL3jZ+1Jcea61Ilo9bmovUXS5eqF/bytwMfp4nrt7XJNyNDBPbuvS2O
OkbsdXMRfoZtp/spl9MBelFmA9+T+RuWPsEJTfnr9SWbVfsHNsknK4KpckD8Ok5/SeTlu5XwEyYz
Fg50Fdk9wn0gxafS8gndmmVPtNnONjNJBj5RHiUkzVH7oUPRbwaPDslBxA503y1hOub2ojIhj6mP
PRvuZXofmaqfAivJQssfyzrUNs/vBdkiJx3mf0yF0wbrRqj7L0pD6xVz3DvUhCRw3+pk9tXjbX7f
/8CzoGi/Kf+5NoEKy8813USNEXNOUrvCKSwbhwRf9opNyEJsDOzDlIxaMfbTXH65Ips064UIvcp3
fkk0idCz2fdpSCqjLcttbqEr/ibmPnnn5Wfv0y5OXyF4YRY8PWVA6KPw1+WA013fNgmDMsYPBiRw
Zd8EcxDHPPtoVyOebj3njxc4Wy822YN+V1+hoFL3QXqzqrAEs9hDc5z49DnslWJyzpt0+tNJXdEq
b61E1pzL5h3s3EnC56jlPhc50O8SdnzEm9TMGntybRYcuIeTEUCxR1oD0djKvsIJNGpxMVFNqyI7
j9Izn3umsTyBFW6gvzpA3FEzVeeECak0mQiCspa6RGQA+/y3iRQSk2S2HwBMWK8vi18HsZlzrY+Z
SGszjJbSbwHobpWy9Z2EBsEdHyRQrG71RLsu/TtA3NArXOFiOYVeoHluA4hQLaPpot7B51ui2vs+
hreRX0Jxl7+m/tCD38UGTXnvJt2RxlTbd6rwniHkXjlTjeuUgfQbOU8Ss447kBs68ylIfAMP0eF/
+7Pe7J+p2L8kZBabhO5DqXekzuIKD4p079jb9oMNpTO051LCp1sWQEiyOzBdEAdm9620mnttSl4F
Z5CNHOalqOwHB5Ed+WKpEWMvrPtninWUX2zNHn0aNwFqmzzPxlW4nOMw2Ynr2MVn+RdJiMp2qAc7
X84uddL0T2ck5+7UWFTbv+3BjfdnvEYkq62fcMsaW77LQRa+gAO3aHZpVPByjKajADnR7TVqY7yX
6zmsEFQllMy/GsTMQB56FosjovoP0Mhy30vxGaIbF1IgD+busTuOjVy7fKtA/0u/LkkK3xmMtgja
xXMBFihBPNpUDo9S/Q7yXKag2CQqV2jMgklz9HwK5QQAWOAAgvXaF/gpPGbqe/rPYPTYEv4bB69F
WQm37+HD14CXkpkGBN6qAZVILwk6bGkDBw3rGQITuLMYEZytuBIJS5LQWP5p0W2RJRnvUT77QvnU
Fk46Q8GudatkTUhfeWuYd2Y+Y6kz1rfBOx4eNzkT/qe9GG4YtmD/ukoutNhvVRxhVZ2RaqhXN+WC
nsiZkXRmIKZOYZ+nq9CTUypqDcZeInyW+akC5d064txQa7rRYLY70ra1eh5bXT//Eem9UjC98NQ/
N/+1ruAzLPeyygKUnak3ybS7DKMYIEYGlqVDm9uM3MVR2a/JebMutbQOaJrFetzOLEzFYLpL3Ukp
4gb9l/xzV7bH214wxQ7BkuXohaifnJMeWfB0i/c8FyTbh8Qid6zDdMlczD8oae9O0RheqseOw5c9
0Hlm9z4vz8TNngZ5UA2RAQnJQBOSEtWDFn8qzEZEl24HTj2x3mq1VUU2Te5IHGumXFkLaOn91cyB
iLQnbH09ZjhaTJmT2IHY8pZdvlg/vytXYxELTeWoN00ffVAyu9J4qpFG4mb/KGG0F2QCw8IohLTK
T7yCrOt7fdz+4kT2BkYg6/foEs6t9jdIS2YKIQTSrl7TejJHLb5isI0mHmxxJPJTA9kDYfRlv16b
aa/J3eJhBl+VJX66tBZQ7KBuYsNk1LGuB9AxqWrBbryVKN2Hg9KYa4KOx8m2aNsFFvuGkSWJBjNI
DAR6az2aTRI6KUvW5yK8MVpYayQzkornWXgayIRHcElZ7K75VG+TaNCXINgxg1DLpAOTS15wNjcE
qQriDgmV104hGOH3pThb38e3VvgzzV4IAI9JiicFNFVO78NN1wTDXF7g/sxQj5wcC7Z0ua4P/1eB
zFtxAh679jp71KgO2VV2W5yGylOVPFrHBBzflcV2XHK6KDEJ3X4wYsLkMES6/5axf5tJF4Rlo6wJ
gsV5s2KCnUEuCkryPHShA3Kurk/eCE+hcpMdvG5fzSNkr5sa0bfwTDwG4jCdWsgG50/qAi3gc6/W
MFbIfmHaxjWxrqZRpVCHHkdNUgIlEcvbawiRWi98/gbQ6ZtXnV3F6oAiM80EBO+tjvDkBSvq3ZGb
TGNgCBbJuRwN398qcgW75ZR6uCrZBqFzOOvCCSwb3QPu1EQ8gSkvsqMPKVSxBWpHTaN0rGr3OQ1i
1k6cWq2tvbzy6BAmncea9FFhX9H03H7qCuCUVeY0PNd/4ANtZKDDMKvgJ8kzLMOPqsjTH4GIx1AP
nOCATRHPYAH2QVlF7J1Nrt0XVd9SuKvIca21JbAuqGsb/YUZYePCxcczCx1hZQaK4RAd9TL274iM
eSw+yRuR/6xJeNokgCdR+4NOzP27DkC3k+iZBTSNewVCaVGeDyplCxVhLmc83gREmXwcFEk/8vqV
Eqb5T8chhUtpRl1+ENFKOc1rmoOjfC+SiFy0C8iWU2UKQ/0PZ/VJFjicYSBCeQudxwa4uJCa+wmW
EClvFniNBoHRW7+UpsJAgRyVS2AXbuLHQAUzVHKS0H3QkKZsxyRTJcFKldfPbCHtxQNkXBUB8Yk0
IrKEvmOMfKL6STDcmfv9NutnPEjru9IUF/O2EFITSIagDon97BULhg1yNmRuDEjYYXGLNgCe+DHx
yJHrIZmRDn1z8XCxncHcfycnEMaJCDgdUhUh2l4TVFSf73eeo14nARoLxZgQ0W1XxcnSlCy5sevN
+1i46wiUpyfYVdisB1HVQqELQO7yXKrVswLGrjCVV5kPaLB2o1wdwdQWxjJo/fStkm/0/rflE/A4
l7B2wg+yZf/eg1ARNnHIycECErYKenCjSJmGUHR2s5/xPecPc+m2qAVqT/DJng6EEoqihXTbCVtB
jd5xkmRg5Rf8AvGSppeumG4VNEYhOm6jqksjAkHq1RZlK9VU9kSvN99834KozSO3tzfSKsEtA4TK
98C5c5nXuRNViP3y2AuAuYespc1o9a792+tvjmBZos7F8P9mbOd1RlTyLZbvr48Wb2uydjfw7lsd
FtFBsseXHAUIi5DICE9IUBjMpSQk6vJLonw8Qx2yYAvVhU8LQHNC/82pKipVdjT3GH5dU1PfFk4N
pLz8n0FQmLoMX00uVYpwLVGRw42yZ7hh5MEBJwXtrASM8xIFzZU97ZrkekfdwesCl76mz6FOt6bN
Bj2LnSOb2ih/dJc6mrBX5bSc5OD8Q/1e5R+tHLjpviN69b84IAzVxRgZiQEzPsq3wZ8dFM6Iea+7
NJIjWn2VAGekNRVnppDSGSK3PZ90FBCqEe3zhS1d9SdvCNSuOuEfuSl28Aqj0D7MZefrbRpvucfB
3oifzw2n1W0ih+8EMKfs4Gcmjy9clyMMQ8ZWOnUBTlyLJlBSXkyP1NhCFMw8atn9vlw6R8T6Q/ap
NQPyDDaDjmU34yWigO3c6MHljKZtYGCBtqZVXDFUCUk/robV6emDM2DvUASYP9KTyOnlvlOb2/K3
4FZDGxl6Xb5vyWgOGb0nrcrLqnKXXs+k0pI416Pzh5Jid7z9x/Hv44w9Y8CgzDhRGJi6oo+0ZLp6
8U45554LXsDc//qDIEnmUsmaIPXryGRYQpv/+rOp/G7n4YXs4XBYDzfvxrfb/oVBjuk5oSHLlMUN
Doix0KQFwUp6TGONDrZTXEHm4qmHIE9BHT7ZtUZR9Y6tfyDmsQVFIvDCWUFVT3OgkVSoBXMhunI1
IZSuJhhLNblm19BBmsZ5TswLDPVsLiGttLEpNcxoamAkW82UlpJ2zeEM9dfYXUUo0KIbigwM2iWH
92PhYFoa6Jdd+BEkQ9GGkWDmU3N7PON5HSZQHrosWDlQVVy2CPaDmHqlvPDgDtwnhM3DHJffcOqn
VQ8ADJYATLleuhcYvAr4UflfqMfNTj8iJHaCuZ5Awa2TN3Y4J/xi5DcToXjDUfgDukJL8Mtn6bDh
UhSctsxlNDeOE4Az5NFP47tu2vFYzzwer0aUywC66sbLxhoaNgSfADr4RLavo6qSbzwE87vlZM1x
t6vGJhdsRUvPJKAGADlu7hqBfbMacphuHx2CfoTgabxVD4E1+AdBYqyA4EezKK+ZFpm7GULIbZ1B
4r8t+ShRehpynyVIGJhbpoRxYckus8bAGbI3lpC3KOZj6Z4si9whEGbpo9T3bdIG2k3rqzn7nyIs
pFdYUB5tmEKo/wvrQlkCyb2FJhSXy6xlJCwOssxZlnNeUPulAF6e7ym6UmrFju6z4aiex18rabi/
v6IjrTmii5+4CJ2onDQOqdnkS19dV2O/8MtTReXdE/QCKnUFy9fXkM4LbRZL4s6Wt8GdMpVeu2Ht
LzrbcbVCABTc33oYrCAyM8NeemdIWCaGDc8QaU4lzThMCS/JDzbJ3t7775GcLk56/O9cJA1l9WWC
1xzUltnnGJF/JSURk1peXw7oYIpg4OcV9t8EEY4kJW0nURpGj8AhWApOf5roGwPnWnYeMHuMSMuj
5TPdX2goDqWkMX3I3rdp0u8VLs6IlioImXnVXz/UABEar14vE2PO4eDYMIG1dzwKBsgzkcSVDnnJ
yHz0694p9dfhiAqfqH9WmvRo67JuwgDPIpZAkOfjI0Vwn28pR+nUlXRsBK5Iq07E3/DMNhpvb6mS
Nx1QwK62qVf2wShMZvTYo+Pn+zktEelmw28xKPw8/2mUCbo/tITWUVUIs8Rut7R0i3q2HVn1+Nhg
Trbc0tdT7LZYzCGdHquLIkXgb04sDQdOQ1pX1puJ8unRhMsuM/6a2435a2NBrnQ1kzB+ESfKmW+J
buEblHNPdiWgTZvCXvnk5v4osHr+srXd0lcALs1ufy3jSO0XHM/81QlSn24RoIxRQMRN9sVq9OW7
CydYcwlYt1f0w2XNKfmidYDWyXXrVcGV8MFQVYNH/Ed380AWdgf6kLWpKkrKITG6rxOVxDkthLo/
cSL9YlklsThDydSK4c/+/b+tKZdMKNbWBCz955hSyiN+Kqezu8HYRXehGNn4FBM1BOkeNDowtBag
uhmq30oKwtdUsYE5oQ4XJxyYGX4aPmdo/9mUGULdLIr50bSOiPbleiDd7QRoXhJ01Twu5F3PpclU
IfYRQcGQHvtWbQLukqRApgY7fuSUoHR3bsyfjMV0e1LExrzjQrjTM89YVvyM+Fg1Zpby1rmp4AbE
SiAULuxRt2fWUYOrkp164LECm5ehkv89lgLuY+CoqqUTaJyH0Pd/HOP3HxVsWRLuSVWOrEmcx4lM
hMFdDdBUhz8FlNxHvamaJARTNUhLUHYSdmBmMXe8I13OlSV0jRRwy2l9+AP+sAXW8RytT/6K7XpD
5AMlIp8sIk2oZgSXdFYqD3NUo5CU0SSPPVUzk6mTWj4oZR+bQnYpYk45yQqx32TL5MIez14lOeBD
/oz6k7UEruN++/yYPtIcpkqDAz1RFklO4yRQYuEcFK9eN1kMyuVYxcVuMkO13DQsWYilPXbIRyEt
zvHgqvjQapsXG0ZEKiFB+pngXM4HGyku9az8PaZwFQTdRJBbHZ/Uwt/kETzIs326ol4r5YB+1D3Q
FeOQi2tih2uSEBvBfd39NDSx1/FJsD0AG0mEwb4R/dx4lkh9IaMGzsOwli4rfayUfvIVFUn5QIDm
w0Ss9yqKTB2B/d1Ywa01Zz8+i1UErgT1A9tPUI0FaPrkzK0n2+B/0CkTRZDa0nzoLnwYGcNJeF3l
o5wIEv9Lk44M+PuspBxrNqy7UlI16BWspJzyzFcNl4m5urSTSih21SO7DXpDAq6UogMXjfNBOJ9W
0woFzRfUG7v8+Pv39ZIXDZK7mhoCeT8YwF8pKZn9voq1mi4y/IKizn7DJoKCv6J8GnkRf0i6x4up
0bV0zJQACBcq/bZzqMTHzTwli4PGJRaoAHjuaR0A3B0Ft7pTiYcl37FdOXRnUdPjWNypmliReG8c
aavwK/3JTiPp483gGs+0udduOIn1/2UtwDJcIu+FAWMRcW2QaQc3IlLjKZ/bicUWbPpT3Vdsynwy
qoZdh2GXdYo8h9A4pX7+qRCqZH77xdtddk6atKFeYSIJmH/0KYi5McTcQcNWdoiWWZJNt3vCSC1Y
76Z69IDQ03ir5b8bLalynydw7NN15UBv7LPbltxNbMvMNE1D4+nhPrYfhETA6w7K+u0NaQVFbfq5
vLeUBwDtPainfQjkuAZAb0N7NDFdncBmYBTgfClCuVW1CP1nvmuE1TyQrRZ5Ene+qzfd22F5aq+c
X6NEPviupSpu+u+Hjq0OE15BmbktUL8nGBvtApC/AeXOyasYjzmBG/PZQ/tQ1DH2Yg8gBQjlIzW/
wTQ+v8g9FHgfLnQT+zvIV+Wsa/M7RjfjVoI045JKVBO67guBedVWa7A2LbECDruix0rOVNiSROgZ
s3H+KDIfT1BDTpucgJXaDjWlfYpT8QZFrYbMup/KfVraWd1MLKn5ArHkjp2c/TWFYwb9vS2fbuPh
JQ0+BGC8zvB/Ka9ane5Wsv3/Fd8AuEdrdOFk/Vl9tLeT5XNRYYXqrTZhW9iznIN5dtqCP2YRN/px
kFN6zhWVFgJCmEC7lqyKK1lsifBJdQGv+yIKWNfWl3JCcyST2LpJhjLOQ/ED6HQXn2KzeodAbCO5
jtRK/SdfVeLrlvsTKN37WvKqBl0GG8bq1ziWTQ1M4Puo96SAQIkMs0B+ZfXCCqnJ9NqTOTqhjz1w
1D5pmL/nx/GAQtXoh8eYJhM2NvL9SKd8Pgkj35EueCvpgJdLQVn6uNwZpG4o6XAGvTgzoqmRR4D9
jQee+C4x9UMfv13MTlapz34/flOsPCmCgh2f+ger/1McPwF2xcq78vMLxptSQ0nf8gq0YB4TX4q7
TlTNOEtf+2dTjOWrN9Q67QlP9efu9s7PGLpgTFEG7ULisMfl1pKL7lw4E8pgeFUgbnEWpUCxhPst
8YerK6yapQBGlB2mlbXnUEP0yCGs9IeW19/JhC+WxBHamel45Nzn2Jrkwkx1vMTOasGyx/pLqGEi
Xsly3qxDAvm+xjge732QeXLyusLNw8RVIEHXh6fAEsLix6wobmiewsEjpsC3IilTo2jc7z3Az2HV
szhg86q5pTredjti2d/J6lbV9IzlyN+Qw0e2EzKAqL06XYexvjSuh/rB88LQjPRmzD16+AR2JMS7
kck7Tc6G/2GMeTA6lPdAdMhmSEcm/feYWtKnRj0rlkx8oDYaojAa3YMCJebEoP2ndI/G8whIaydp
t+9KBZ6dhBJZ4Coc5v8R8rOg9OST7AIufbVXvXjCSqGJJInpBV/TWVSdV6l/1uUlVWfwpjyVu9l3
WqG8Lm1gEDaFyMPP0uEVrVVf5UY1BYrBT+eo+Ycku8qz/8aH+/QRVQILOTSR1PZlK/8/obVk7s0E
Q6CgwcYql4+GaF/oM4HvJ11yrXcCqbxIcVw3YdXYm+j+oHGyKsUI9m67lnLqdomcqPqF4pBsTVW5
sOwcSlaFUDPUfSaGfOjDvUPKbW7AMPGWEJ+9DR05wtKGR0GCNXNKl6H7lwT5HrVW1xARzGxjo2bq
H7dVghEmNTRDMyac6oqB1o1AW7RgBTMfXc6nogVYC7WUnkLmPLLnOIzA6FdC44SX3Qf8gb96Vngi
TVH1Ilg2swqAIhFxFfXsYn3OycwKCgTpf4S5RJ1cxL4brBB6NW1todT1ULBsWBw6Ji7mSfyQStjI
YGBYMaXA9G8INeJw9Aqcqsy/2E6W4vADVrzuzgiIJSZE0nWZ59vqH73f8laoSqYWpwmfOWRYjgcl
HUMNWfRMYCsBsxEBuCOhCp0vUUBngRUYGABFZA6WHq2xVKGG4aN0ZL+WGNZY0EWvus5gOA3xtC2D
Y5ZGOXRoCIAJ+/vQgCsZ5OfOOwZRFAsb+9bz/u6+l+YrUelcMPnUcVd6+KEPeXylAmMP66po46nb
jgNVJFrRNheiQXUCQIv2ANawtL7/yvClIhia91r46mda1IwOvrCPGimXJkoZMiRppdP0bQVZYMWj
HRCuG+1shFD7z9/0ndsnULzBkttv7oLcdoBF50aLTNq1g44h0XGgxfAg6ujo3WM4GgwJaG1Eyc78
BRP+AMsUocOSMaHsPNOghmKkzhn4mIj1Wlxc6bZ4uxU0jVc9cB08oMvhT75DDe8EiFk8Z03Frvxn
0DQAnKtQCRu2GqHY1uWW7jnMWx2MekSn8gUydPMrzWQERs8TAgsgZD3i51GM7qc6KtV9LHl2ZQDu
8I2LmECeEpCRMryxPpLGzd/BU39VEuKAHgU7M420ETFvb/U1NVwFMQgLV3URjDwZIjUBkHjzvG8Q
cOJ/bKTwBXzWU7IUy8W6oJZ8XhJdqti8LWV9RIx29mLcn8H9+Rf3oYJCR0WUHSxoLkQ50UwK8YF2
19R9ElCvrCFkxa9sncqE1O0L2duEo9qHviHP7vTYXCu/5QxaQcdbmK66TGNl/UesF0rRBO3gCKgl
54so97RVX8c+tTWE72Z0Xv0NpomgrwY33oVfw0uGVk4IPnIcEu462rSnXeh+pbqOtHoO5IxDlH3W
4u+u5MuSSRqKpY6bLTW+mD+sbFlSEqakVkzq66dt9fiLgMm9NYAuqMENGO1Pkk1KUYm6wNhhV3Fb
p6Z6lQ6eNzNWu4OWV6cIU6dqgVLexf3ql6vJwD9NX/GWikJd6rO7UEgp1UNS8p2tCiuNvyoVcufn
gX9WinB366Bke3kdjy6FFMEXR6lOeHUTQsmXI34Xt/q+G1qi2Jgl8/EKZLhRMpnQIKb5ICtt6Y9P
bAUK2qwI+ORmToqnIgsan0INf9E2Bs/xp5pzgb6MhDIpWa+JvkQyTPiTM8ibWSSresYT5SwP5quR
huN5AjJ02nbHoctD4t9Cj3H+4VfdZAQFquqHn56+9D/mToCbdBzf93r05X0DvfFBhv82YI/WAt12
U9hUQSxJ5070G2BleXVU1Hf3jNaZrekD302w2Pw+d1U8R/FesY4TwS5rK7wGX1QXgyZ8bnVewHp4
ng/tfCksGOYksVbgiYYXpqScu7FC7rOiU+CqU1cCWs1hRlCGlTZqAOcyYnw6L0Yf9RfMWOv9sLu0
I7HOBX40KnKi7GSROt/Gt4F2OyP77dSi9SKx6QmQHVRaG5mUm0QkEui/2cDRRx12Ip6Q3Um8gcvb
ahjvfJ73kaKUBXVUt1znar54otNrXYsDsOD4zmEJJOiTBY6mRV/KFrWvmIUPxnb+vIHEBWhpCa56
cx/2cTETrmmY+j8tmtYXdHbUzY7Emtk39URbfWANJ+WfAPJxH3Zcb1S/Z1IguTbgNz3GyFLc6aug
HyVXfzrrWc7Z9lWD8ovoPvnGk9iijqAcKLr2/B63/6tlqNMP3hIuWMfuxNZRGoPqfMYOYYqOK/bV
vHJhREHs2V/Wn5Qo3UVANPIibmZzOgD3AyB3Tp/Vn8mpN+Qz7JBdJ3pfvdD7ozVZmifHjo9Tnywx
tPqeseO0GgeJka65nAToprm4GlwWfuz1oJXhCmqbkbGXRxfY2pTYYHGcbRc3gN++l+8RyUIBXGyJ
DZf/mvZ1rgQzboSk4ep+PdDdlwURnV1r1K8aADD0eHb6uK3DN87KDzj37ECH9tXDz0yoAr39kZTu
ur9gCf+MOIPIGiyKt2Sqx+cB36NMNlN/CUW+ISLACiUqFmRiBTnEj9a+fBRfK9qDLx1hVAT6Betp
nG8/g3PmHKJMi6zANFgPi6WSzRkUdzi1pIH20jqQUVjkIscykWtsYOPkMLRnhdmH6ZYRb50wfKYz
d9/8A5JZxXMYDTCYLX0oLPmcZvBAxV0YrJ8P/4spTJv9Z/nL62QMGPbgxOfYVK2IQHj+dr6KzXHs
Bv96+ppQu6D87oCjeZnApJXfw/OSm1rrfY4wUqkvKDPOrtBqO3UvPl/Is6MUtm+NA+pzUE8nawfG
iDlApKD2YY9fbqYjpDv8P/4dSsmxdiGkSsBU7n2uvYujJDwNLaobCxDjswIN1p68k2cyItc2/HyH
OhHqFPCCOsRzemLZy6jXrIrGOuzMfSJyVqjHvB7rQzZn9nptFAojNF1oiSgKP4hchMoRGNI2Zp1i
Ad9E3QZgdM5OGPOoLEyapW6kf5e78wNZ2rsLH+TGanWQiAsDQMD4dCa3/9lD3swnQFwinCNrzRLZ
LhygfVrPkm0ECuwu7lBwFZiFOTTmNQrTmOmhWJ/JWr8o34QlQhzK86DgYYKPuEeg6s5TMdbnB7b2
DLwzJezfaLIkp+Swx2w59M6F1eemryDvGL2VIBYgCQn8qrOwNG2IdbNe0UiV3GqV/xwBKBmRaLEp
b8JjftgrjVBT9phEQM7UX+0Up+dBVhDWOCEIEU+Gj1JVgzQBZEg3TvSaSpoYxXcJQBwSRoL/jhJB
+JUr4zkCYeFWzuzcZ4NTaBzssNbi1i3QzYc3XOeh1Xs5819hvmB5mhbjls8pd1tRDfjcaasDFi9G
tjL/usUJHKVkmh2V5GXYKTO7Ad5QGbjM4EPHjBNU1JQcXw/yLb6V9ukJC4HzLmLgQ+Cs6hEHGoXP
eV0+43DuCvPtm1PUbqMmR6d+eSZT0QLInqQBGvp2SB63QYy88V3/tnEMWQHW1EcMynti9EqvuE8p
eelsrSZEIEYU9YDJlBCqZLtgmJ/d/iWZM1JjwN8i4gyg80XSXk7GmCIvGhIobLSnC1LH1lJbk1rA
/AK1qQopuFKUNVp30lD1JajvdHXK9pPv4FfrvjgvBh+sAQNpe/spcPMYi+0xmodT0OEv5UM/JDe7
NiylNJjAc8k2S7wIFj8zxK/kzHYgXCX9dRs4ZA65zvETH8IqHUKEGrSF3Lko/CIejQFqz58EkQmN
F/3dlXu4z7EK7oCMrD+y3n58eww6zJzhl4FD7NCZDNsskvLpx84oVHix2Ut6eVQf27hbGSLswSCF
z4v6OsdnaToeYsNF0VStBdn5ELXTxpdcMBq3diQfXUAjGldrcnPi2UkeL8uJ/Qe7byROS9voRHce
ylHp0VFaX2Ip0A7gXu2cO+7FBEYXlLJ9ufcb3laPbZMBxYF9asztugIKDEZgkwkTQZ5wAZwlqZZZ
uhH/J/zGIyR8HvWP9u1Qd05Q6rb6x6Y0HSee+LrxQTdaSwPcMvrGBBS97Qn5/us1GAFrpJTx0kSs
BglLhDH7P+vMfEBytLKIGt548XOE/g3+C6TO2DDm2yY0+q29F6coWsMM/FUFAZiUpf5mxl1rkvN4
yisNbKdZCfydL2bAjiqQTW/7S3oaPcJ0vbxy11fHAJrFrQd6wtGsS45krZ5J7ZcUcZ1vsOD/niE8
Nu6oWhyTtbPiwmK/8myD5VvrnXd4ZdC/fzMX0039cpaYc3xo4ukAPn+HAY6lFHWW4Koe/1MuCOJZ
JOjo4CJn/gfmiLaWCHCtsl6w518bTkPP2y68Q2Y1AqVoTCbE8k8BbQzx199gsVdUtUUVtaCvF5HP
kVqRMPONLQ1pndm2cM8ulqsU8wE3L3WU1zSdYE66JiM14Z07wDUgcPKkeSd91mmuw1xfz8RHPQ2X
LM4XSLSI1pcErr08YnA0YV49C3uDdPyY8qrGOSTDK5uVIjkIO3Dz25pFB5xeVTQegT2fZ8rge2CU
xnc1YenEEb9WZwKrXA5v9F3MpDFt0bt2sSOy8sfZSvZ2o1ou4RXVEIk0JgCsL+rsiQtb/eLFp3bg
qplK4VZGSdzJIeFt6fqGLqm23Yib4+1D/kvN2XztfEujTs4B1Ltj2ih40O9T0JpocvZTVPaMvTPE
n+7sBTmJPnPY1za6G+hzp0wMXg6B14m1k9ssYZ6pNJ8nD64fWP6aJvEtllEV62LzkzulLGHpLJPm
HJymmRPPJyCyrqKfU8Ri78VyLXz4qBoEDcZuLYegXLie/6zI8deZCy2TVbb3sq0cHLpL6zOrRX0Q
UyDgUTaaWEifoSLdNBwgx2igFHCtM05+AyE6i5BwfOZC9qF42KgWHzptQTPtAtjOHr/lVuxxQ89E
y2aYNxVaefArFGfKB3QiS8J+Qh8tLfYucRw8f3nm7moKlF40H57KI72R6Xov0Y+T8XfeJqO1SN5T
r/ZLHnGPMigv+zU3EKghWP4+ouUkdyeZcqui//OCuwQodgbvUW2DjGnqCDyj106Tx3zENcSIdY+U
WN281fbPWjMKUd35F1cTJLN4kHMzWvc6z6d23ZDJRDtLjS/GphY6ZYMbnGIMMhs8lzeZUNNHK1hj
KTslTOCWv+liv//LPJovddcmaMPfvBzwfBrI/REj4nTeIyDJw+yAgGv0jIzvX3JgJcLOUo/UQC8z
55MPraHsKYq76fRQrCJB19UFuWMP2kRLixc1hBRttLLxVu7xIE3Sx5CXeK+XzwD/WGmzv6+KROGm
3SQiNMCqilC5AKPsTTXeLItN7mWoAPH5hPFXHln9vumcmhGlcpjM7ytROamJiwjIcHruSpuQkTi7
4rCQ8U3vzlH0DDsp/mJq8HvNFpUgACEk9wIMOV6y7bbfwUINqMu5XYd2MQWGR0F/E2et58F7hztO
yMC/aV7vZoeLEUfa1Q/os2uD+FMxHYfQqHcC2zZdGpRZp0t85qk73ZJImmOd0fbu07na6uul1fLF
dLzsZas1KcKmvEDqL3rsAr5e/pv/kAkaseDrTx+rTwxH6+Z6wcXVdWsEcsCYqrY+13PcKuuCcg9c
GPb8i1fnfEqszefBU+Ks12vs3vLArvE+BiNv2G9gqpXAxJlfczEsdk/UxNG8Vdd1ebE3A8Tyy1wD
UmwilVF+keExR5d8ZVATbnCha67uyKU9WhDzyolVw4ZcueY/BdZ5l6FiBJ1CcWhGZlOMkHuhrvPY
mbCQhzLl/CyGMsU8/JARMeukjaBSV4s7+g3WYetSpaXNvqWNd5FbjWuDp3jGNm/HaLJJewVW0f1H
hGE0mmIblpXAUaY4kv+Kc5EpLVL5xRQXPHbb0mjEO0X5LXSKbYGzPpoL63A1WVXi7zq1x6pPrfkU
GejbPjjz/ChkgJp1Yo/zSulXOiCb2p2tnC6dzsIYBFxOi4qVtY+RuELCclzjrM/fmf9ZcevoUapj
vgx3btcIkjCuNVVJyIH4KGqgSQ4OosAR5kR2QgWBm1qHB3iKgTdjXCiw6BhYSALreZ3qaci2iMNJ
Y3dBE6lt2sakI+4SljxO68q2quHpmrSkozIlbwTH6IHFoqI7RX7AxXuSG4bHUnQftmUA+OCKiD2j
ffeI1L085nGXliKI1yIff5f9L7SY3qtkWF1V0OldCzFqMlfueZX+3mXTYcKifsADMv7XAoey6xwy
yBMukDggglRVnsc3p5TcDgHPg7urcmGGvEuEKXTFBL9nYulOzBM7LFuKSIQBhwSEhimZ8BfxlAO6
vajmFIN61tBN5jYO9VnAJqthvZ1pGBlzSXImwe4xlBR4+inixCvcW70kOZbgVky19oHd+N/FGEKb
5bSwxsuBdipaRIwpvBgXIIn4FVOFIfKDM9nsYH/OLhs+J6KA9Awwd83gLHWgr6/nUEa37PzJ1Afa
0h0ENeQGY+VMHGWGLNLgNkEjghdLusQ/n3DSXby8Swgfmsn/qaDQsBNuSFlhBflburvMd/ccNTlm
3DQwkO+UYYXJwJNbvSuMQR5gK2LUWgAIXQaogdrT5iTmQBDERUg+8bMDcpbPRU+JuoBUi2aI9M2o
q5HnNB9tu/5AlOlzbzdgfF1z/XlXmABFpY9hWyP/0yYRiO9XfuKcDredp/XMjcMeeW7liOUPffSI
aFDT6FapErqsxRCEL54e0e9gbZwxPlJyPjGlsTktkyl8O8OqcFRdNpfZygrsI6z4WqLGYTA3LTy5
bTaSjoHmHvOpIKd8Lao5iDWN4uEX6h7RsD0ZWF0JLfIPS3xj95C1osF4fEkJvJXx8QTJktF+0fyj
g4fz/L4R00TqVAIDg07TtBQFqPX0z57D8XKOQdazAOYMLtIfPHIoGhKzzUhlj4aZSfSElpRR2pTn
Tbgyr+DIhzH2WSwhJHcsCmNrCzLdnvWaIVVmaFiETT3kH+c0KAfvqm89zY+0GYRjiqSqa8g/X5Vi
7ZHE1ARk3XZsyA6Of41usSOGtpTl11TAej+3X2xdiL9BS99g1oku7k3b18jMu7eqTGThDtEvmUhc
LBCSHnrfrzaRkluQAHAfgUiMDQ1P1ct1SWJYliuINqxJumdbHw0kjSeSjDSNPCmJMGfwOC6UIBaR
wznsCtzNuwOpepvNMPo+Ou8W1ByGZl4ZowGHxbsuhsfOg1xIHT0vEt30JAclu3XLh2mdCdBQoFao
xDXZHQLtwbt6pBVhmlsvRXaujp3N3hTA40/+Gk1oMfxOHUGJgGbDdz7qjmMwreO0VxJDpLDZ/9BN
ZSVAp20Cmyt//Nngs9Yg6GywUAF3nYq4DSif+hq8IfNxQ7gRi9kTVTr4DOM58mbo+emcjxDPhZkl
F8LZYqVAJThxv6T3TphfDc6lJQ0ccKMWEryZwiJN66iLMVwkoaWkByMsHAOGGMTxrKdTNafiBops
5IxQr1kXU7ojBFs5mrBrhfwYBHZICPY4tRbmwqM5czg4Sk6xwG4e/0HOjp66i/e+rxUACLJfn9rm
K3UmrjVvg74Zw8CqKPJm9hg4OkrHiXzbLse8BOIbk2yd1G60kCXzewktjQ6aTehf/f2QFexaUOHk
E57lZroEWXbQ44GaQiJDgjdQe7Mmzt1JbhimCcIvQMdHvGCHi6VHsw3angyguJpArbtOEjBXzY/+
h99muQ0LmtqGK2rm5oYX7KcCgHn9sP8Vlase4grSXXXnX0zta7iDjZT74LFDsoXQpfxsDvPkc47N
Spt4elZ+apJ2b7x1708Y5Oi4zTdcKYXTE3noFEArVSd9gsnl1g9mkUsB1So2Z/ewxk3NLH4iV6Lx
Oh/Fd98X8bA9nZXnV915MHOupartQ4C3wmkAcgZfpPLjnPL67l+OZ5pYXMrRqsDh9oSB1UXWZ7Hq
RiugjSU7vEjp/4A8iy1nTZL7hcsqP4pYekub+UvqsPFJHB0uigXc/iLL7amuFe/1f1nzRAAUN7N8
R7LaJfrzhkBomhxzJKemYulRuBdO75R1bMT02DoZmCl5fMQ5I6jDaQAeTJo/Fb2VcJN999/kD1Pl
HLNVZyr7RfEHmAiC4rmIBv5qa+InY2/7VAZDGNRLW6CLAQjnM6wiP6yrGsQoemm/6LM8gHmbQ8LO
/teZlx++7s78RfnObwkw+xHvDDBs5KGdqWDQpdgfocNl6s3CjVDP6oVqNcEimJnvXLW8XsuYZfjV
Q6dsMSTAAvQyEzhDNr7xnmQ9C3cGY1q2tFajDUkj4ltyR5CSFOfuCAdZCq+56k62mPdsq4xDLIWh
5tsU0q24PDH6uYif3ToqK49oDfJf8ylr8N3mkrkUZ0RE8jC1k01p2aSI/jGdQK5Bsk41Q3dK1FVi
GUjtq0SDkmk50UOBEnQ4N8j1hjyo1GKpmHkfaj9QRxY0Slps8NA2GYrIFin7JtvEgnvDIx6ygYUM
0oxsNWG+ciHKSn3WJLGDDhZteA6YDfG+AiQngWaDwGUsB2TIyLvg9M+UpDBsEtbuVJ2mUczVWZxO
/7a5J+7bD1g+OYDisAZI9TiiMxSNRnVYlhBuER5Z6I3zHlfxoNsiCfLeAR+oyzhOoU8Gcbc3DQS0
mA+Jh42kHB7RKEP6yNITP/JAjn9qQkBV7OoASxAbCyVw+3szU6srdGQ1SyOClHyIxD1evH7vD4a/
OqDBQcu/OC49z2xKhfrXGleyBKjzBK910vAFTrGEFggsem0ODw8f82bVUOF1z9vVsxdsMrY7EMKx
m98wZlpyIJi4SvYbE9gPQJ40L0RpYIbb1Nwfdb2hZkmS8gQO2I5H3KJFMr57qYTTuZFx5pAEqP8T
k4vrtZnphaDV63PYVKGWZ6D+rQ0SMrOdG77D29rZwLUmZlssG+6cWLMwwzIEdCvSiO4jKQ9Zl3IO
v7QcEbqJFYOEbGvo3GSIp5jBnYsX3ZJAmM7IlXP9bpRukESq+eNSfTou/qNX2XEcrrk2JYYL42JF
lOxl46zC3jFgIXSREDNWQ5IdA0Mcb//v2Fyca/gURxIB0/5sBkasjxXfWrv8HLMy5YYaNAjFUFov
sy78W+1moCo9sQNpuCJZoCJuNyYMSqtkUE+OTJkxSXtN7MnQRn0nXvAAE3yqWOzhEVzV/8xnY4AO
qwF9m36PfM0g3DqbWsCzfm79HCDnYgroaEvXA3VnB8TDuDFMCDeeTz3m/5n4vyFXH5+ngVWD9mbS
i6mmvJsbGJA/kIdPLGFb/h49gKAXDE9kOP0PKQtVHDVP5oiRcX2aBo6Z+BD6nXMQmNSuz+o5/Qz1
i1HH7L9I5vsY6JnNxOiKSVWhq4GYLzuRYZC2xGPeeVhnhm0bu5PTuAtYSL7sYnN5ZH0SF1oAV8oQ
ZFb3RPkb61fM8cFU5zHc/way2XtvZCMZZ/fP9mSGLm2VTtQfQzWybBrKCLISbgt03OOJXxA6fasm
BOzxIGclVSXIEeivbGnBw5oBk8/z+Tz+Y2b19YIeFgXN+fBt+xF5eqbC69NApJzISCYAivZyqsVP
ihxOeyO4ZHsdIXCwm501QnskL4psjDwh+9eNP1+WPboUm/8TJ9ZzhRlmYwMHF/+R385FKvATXry0
zVxyOLXR2BT3j9PBnSq91uihbPgQJbHCpqpgemhEB5z3PWCFKEoTjGoaCET2SpkAnQOOnUOYqhJw
lnicES0e+g0KcrdUIInumq68ibwHvDRrlhekODsf15j7rPqmVlHFEH3JT2IJfW5zFjIE+Irq6RTl
bRWsVxsQk2HHiakuIVjQVJXjvNCzJjyMxxRyeV9i16CNk81iPUTdNPsJRRpXWUEDIbI2Tz4QJViH
MIRNMEDNpO59iaQn/30IUfH24t4M3C+6hs9BQM3yScqVlbt7XUQSyhnt0l3JuHr+icZYNC32kynB
28vJ20VmGAJ6iXTTb1biU1R5k1Agret+2JoaMCMtz00jX6uXME+h2aNuowhp8MdfkVjF3bFUb+CF
JhhNWJz0HQ9vUsCcl3ZlvW1RfS5L+mVuRitUaId7pTYVWplZSAD1kpldCuAyx1A1YTH6rx7OSDUU
zaAHWw6dkKp1SK4hZgDetBOmdLtpQDA3BDrUA+OdHEC0oH+ldIlOgzxGjMN1dkhYSCg7nccffSAD
rm29BZV1Bhq/HKVhL18KrvweTvMcNdC8st8SnHUS9xKlaw5I1+uG68bjrM4H0Ic3AT+OlZt/ngiV
GtnZA165s6k6kNYcIlqHrEbUiguj7R9qDls2CfT/rEtTyIy19rzHTytHhoLbuu8P+ylbUlDBlJ8p
H88sAeKmriS/q07CXftvEhi71cLs+DKuaQmn0Nd21AUvb7HHAW45BZT/x8tj431eloutqLR7P0P2
HoH1D++T53o7pGC/VvjAxNbo6W7PyI5No92qAulQQstM8TY8ae1MuYecBqJJIohrzjUxx6+m2aaW
00yMqA0o3nov5x1zeZAUC0ymqpMLb+x+ArxxndSbfVH3FfxWcW3geFdPpQSTfbrMQIRFk6H33pnx
IuQYdmB/Mp6r7ImWziNkn5Z8d1hz+14zIWlQIqtH+IjHoVf5cJsUez3qVk8TDyfAAZR3V20PNTKM
bxoov3RYtwp+Kq0Kw+IWLeUS6n5cHHY7FONTI6esqQ+KyJpt+dENE4RRBsSL94GKbFFKb9zlS/2o
OXes77shOhGoLL3v/U0llpGUzTEjS49BPBKAV1KsxkUFSaZRJ4cH00gwDk0CJdDkTGUBYZYJHTpv
edvSBZ5rR8+lCA9aKQe8yCxkkQ+7IzOm2eeGX9MEZ/t7+JIH1gUqxiJcNG79ZsyiJL0tyQu6THkQ
smnHKGiMO8M6o+TutCQF1M5Dzv3PDCDb276C7xobBapYjEPITc+PbLqdfqyTRsYJJGhUB+cfFLRQ
d2LWoPBuYTFchohFVnS2WsEyEWLJipp32njAG3UAn6Ujjn9r+ZMRMV6TVDbJ9TXsjwGMlbbtlWeM
EvGDqKdjBUjxrKgHeauIWnbzxVjBFlBp5YnQ7syFoYRURddLnktmCTNo4z8b9QlnUa8CP7UoNjny
NjYYApDJzEipp3NAWoyeduGGVQ5dHdSQUzVMPvxd4EsHMXzkntTV3y/GVdsFlGcOjRtVc3VZy0Iw
4pA6W0x96ADdfhqGH82FDF/xZ68nM3EjDRwAxm7hNdzqy0LwN6D8lqSM7sV6Jv8iEb5WzbzGa3o3
TelrBScDLhx7A7CA0c8Bjgg0KyAj4SD7yyk7INVLi1AzuN9cRoSKL7Csma+sopTjmZmNVAg88ygQ
lBNjOgVL8UX3SVXhAepAz5X0Yhn1m0GkZVksHW1dMDUZojO92/l4JUBQNY6CQkdX7/2Ns7vRZ4Bg
hVpt6dd7YtMbUrXEaSi+ZntKHZA7qFAmGud4hy3GrAAx/zwfBL9DuPoxs7Bh0lB5Wpr49+fYW2WO
1Q4Xp6jQ+IQGFKgk7z+PXcQT6862bqgdqWb1WgXQz8MVIvCzuNmFJo6hANxVhjIohWN3zRrbTegS
RZ3EkeoqMBTg/4uSulwpvkv4sol8tpBjPOKx8FM4Aa0lZ8diCPHYlQ91paNE3JoK4Xlyd7QwpbFb
CawVXDtvf/WQQQZ1uA5a8AfdFM39GPCGT3b9LqoxnY+Y4CDI3EnHGjMJYNgizhqHt7MVrb0VE32d
pxhk77JYnePYdVlE9LOVos+0BeeQvQVp+HK3syjmneMw7KKKalPDkL6Z7I30SGLhjXYYqrm2oXeT
xz5UDIp80nT94GRo+yZnKDOwdn5Zr8FvQ0vJNZPBmE5hcSluxFNUljM+2lZrVqpGEO6K55yhqt2R
PRLm2SbTC6gE20mPv8imnRpVJf/mb46qw7L5IbTn8C9Gh5O1LclAq2Cx7SA+zkr4HGnQhtwzumJo
p01rsOr85mV1f2QZJr/eTysab5+8WtIIjEc+LGuUEDNKTa3+A/tixey3AK6v0yala/9Lz1+4zxvV
mv8XysVWWDZMhm+bZOwB/bEQVgvujmhylZIk1cnRd+EcedEx+HYsHjNS+NxGjyImeT/GgoVvhGU4
55RnuvCzL+EDVC39iUpE2dSFkDNwTqgoIPS0EQx8yw89eemVIPJ1KNil8KjtE0kF/FKRk/LfKqdK
gqpn5VDE77/il4o6lVnGc9ORJx0o1aLgOXBwMpsH1p9oVso1FilpVGog4qjgvPpJ3l8wT8hSbUkH
H6I8MHr9eaG4dZHsCrJtxXyECD+NI0PDjFVnQX3eaE71E2JysFVNMvqOmj8uOKY4KcQ5Sfei0XEU
+a5tZeWNyet8Sj7s4qo3APU9gp4oMX07q3JQUDj8V0O3MNUpthpSFP/vjfTNe0wUUdlfpr6ON05o
oyBN95e9SYmRz4g0G8yXJ8RVTpFwLH4S9wUHJEcWbBi/mL0hzhGVpUkFvX+UYC9Hzkk1FyOvEKLY
jN6s+ypFoZ3jZ88m6mGUsAgMtp1w8ixa1DyJhq9uRkxJE2wh02/Yue4tmGl4TdZQRzUiVHjVsDiX
GVJPkiKf31ofMpaobI06ee6HcwLdhUQufbsqePMBPhB+GiEa4NpV5YAmLZp/UEN5mYP2ZfrtPyJY
6gjk0il1OiBm5Znwkr7vhvBGit6MYONncNbx9z4ay39ra8/zJAD/e+eB7AfUZGRXe0ZA51FioCC3
95Zi8S/X4vjb0X7GjgrFwxgV5KzwdzO3RGgaUYhQOrBOpqcQyvmp0GA/yg5AQsh2Gl3/gavLOqAD
EbfOGQ3PDufQ/uakXnsOvYFOqXIrFt8IkQN1FS5ME0Y7/a2HX0kdO0P7jq6mQ1lge8v+XZmSecTP
KdQEx15ZUU/pyjDxeKfw5c9nI9K/WAVNkjJSZEws9z+Le3G56pyhzmCINHnjPhzUEiXCDV4GKQr6
I76uNV5wYFDCD8slpyeBbkNw/8puHSzND1nTKPS1d7/xe3RSC/yGJvQDribNMxJWzgOMvbbzGpyT
zFBNauFT7tpB+wJSshsSpwnPziLGFci/ILclVa4nigRPjp1vsEgXZpMPxoSlNnspIxhyRH563r7U
qcJE1r0T+I98y3+kAzXdztjElOrJTY7Iy9lpi01zsmty68R0Lo3vH/GbcyfMvyEkuX4G6KMrxgXQ
0eL9A2lbaeJTEeolgLg50SHFWL1DuQVDZQVjgZBbKLq/gmQ6z1nr8ruTtkf3SkbgPBXKKEw/nHRJ
zjCggwEfGkrJ9uloVqk4rOmtBQpiPArB4SY88OyZI6ZAUmjBksYSmiLt0GSfF0ekPdizwBTC8bES
SVYzJhY8hrQrW+ToCQzpO5tn0WjzOzzmiX+mIe7DB/a5qTxzQpbRma9zCGwK0RcpFIMCq/CMqCQ2
xb8NkUfwian9fIQ6jP4QL/gpzn2XO97hvORIDorQ/2qQ1mwUp+BmEWb7Lm4oKTE4mbZwTqaD3Jcs
0nXA23w0Mb82HjFy3QAyR3DzrHvF8WPtScpNHCyKwwmdDXorO9/hMomThmLZVtW+r+RiHCpwTHpH
tclDFjU3vstEEzfzPBsjllflrgv30Qd1m0niF4Ts3w3PRX3rUWUZ/R2qfjq3cKOEJ5UCpfEJFGv0
vhuo9c36haS9dZh+IAyYtmMWrvrxOGlEsvvfC369aCu1bvFRu9roXTCypbyKhJ0L3Ly3Lgyg4zjw
y442/wEAHsiKTPUVNmWZBKZwuMpPm/6d9QEs/xMB6sci0GP7FSiueoQMRGvHTjvITMIuhaai2PKV
i2Orbh0mTotBVOR4dKHgxaBJH2OCdcXY5lcb9UbX53SW5er9rsE0rrKhp+R+eIACYkdxeuYvnbez
fonbe0hMzczYKh/hSeaLhIIEK5MJjU52wznW7wHvsQlBLaTVWVimGUGj380fjk4fOKBHNu2+9CS1
CXGHij3Zzlr3KA+QuQQ/11KKQ0V8Z1VMrf2iIoFxEayNsxkd3Eww86EJnuMol7ORgtHqDGO/nvY7
danvg7eOBr5Ok8dIyFOruVnMiT0l2nDQp4a2bDiZTe3fIWj69FL6X+PUcXiHnIncEnsdaC1xgDyO
WuBnOTLcYjerx/U+4t3lSA5g2db2FZ1bmiKV54wLZE//meUhfbViF8qczh2fsgrUf6K4FMMhKG1V
fM/j3zSnxdQxVvUwWz9jB6s640zgPuSuzZS9yHn8SKATayHDOxpqXuGA9isILykcWWZj+ZLMSHrg
hNrqoJ1yjHWnD44Sa2R+20RFuJvt0ZnL5ujPRMww1cXI0f5Ylmdcm09NwbOlIwlE1qw4Yp5BP1xo
Dw0+jtywyjI16ljDBmbeKF0eiNQu7NTdWrNpNdQb407JDab8ffyuTd7BHhDTECWp6iqDg9Zs1HDW
2344YOBbVRy4rJpPPb4ttswo40a18R/dYKTrMqYz3JogEbfHa9sq8YbHVc1RdmDjfrv0ixslAZtG
zUui2viQ6JAgD9476i86yLjOf0DvgfXRLtmtV6TGRY/iIrom1NcJW1UMbB1pNchmtii/Jgtzd4QM
ZtRDx8vJ7eZL2ipSFunI6nfXb986tRpzQxxgbFdS2Bvbkg12f77cJ8JcbbSIJ7xk2CgZOWCCLpd3
ghXluaSv4rL0cJezmTs4DV3QXZSZ8FKHqZWFa+0nuLK2pftf0hMacgdUsVYHr4WNdgRI2KWbaZpS
2SK53QCPYS8R2mSxujFUxw7NvkLwBAkXCG+nJP+tA0gUNsllPtWroU49scAsy9gbuZ2W8gwzJaGm
qHGiPRPilgbKrLPa37I0i7oN+1wDWU3+Kvc0G19OuVTMJpHpxUiD27f7PSzccu++0nynjtBskzpl
GHsE0LGiU681K5sHENM13+5ZDYUUd7yrCvNaT9JIwR1fs4zvNW1HEazGXYD8R8eA7vfSuieewgPl
B/Av6+JaVHNB4BqTVdhrZUJWtxO5fsVi2ra7fz4Qf0aD5zk9cTfaAnUtdX+2/lF67piUQbjWv3DP
TEwB7fC6lrBTBGxFedh7Z7y953Ewt3/YVScJXVAPqBpLX9YjJCj+4SWZme8l8Y/QPozTt1LKZuFv
VtMqcR7739sy5EpXurgHDOKagXB3niXm6G/eg5nCYiHYS1SDy3m8jo9dMDz16j2mNVqUNlkOiHDa
1KHhMI2GZuKnR+hA+A3qM37iSsnGEE2MDK8zv4Dr+OrdkC03R54WcDH2AS01LyfjA9NLJeGyVVhl
UZUXX2rqly9MofNOBK+vZLzcGpPjLHL0zD8Jf9aQBFyMuvwlWexjDN+BAT8YLGHQ9xgIH9rkD+Ll
27teS1GrThxHAglZJEN4B9zAC1ASck+YGy1AOHqp9IOY/r11i0giP3sEIUWQO6Mel76GcgeDz4UN
RsBsws7zkr2LWQOc0mVBwp+L7FeDznlbohQO0eyn4jeFO8a155qdHTdXTShFCF3WEyO//3vbxhbo
2jYt2kNdPQcwyr2ulpRO7C3MLMuF2TfxpsyG0qqKhhZ1+ZZymKE+O5iQ32OhYmrEKL4ruIvDuLhg
yksuYIWNg8xDgrnOdGeyTToQKXzgXRVbMGzQ/NMWJd18fa6MVvEhf8FiAgVb3RTZXD1sArJUlyKT
lpS1qLEhKQm+gMxlUhohWlBXOa25dn+tpKpKwzVX7+lq/H+gVTab59VEYfDqxh5Pxe+gPhKtiGWt
Ayy79+5dKxC5O+3ODeRKJRfccy2jEqZsOW1aJ6/7AaKln8bchSASp7DOpn/vfh2Q6LfRxZDKwQQF
WY6r5PfK262T2pjEcU2H3yBb0yOsmmqui3KZcxZ+wljvCDNZO5pFPl5zE5IQ8pdypuNmt+AoCagZ
ZzdExqzswo9cLcw1SU7nzvNavCIF6doexfz0ZDsm8flzdI8BHXZRsoqQ85BSfXILbTrcRyJzxdB8
ezSgeK/nXIBjn68ODcO2io92BV6Jxexb8cMmkq/fgBa4UYX3noCfvvWtLFZ1tBOjkq+C6tOu7cJh
7lfORYjPIJbE1Hs/GOx3jkURdBBhyILpE40wHTLl9u8zrZ46BSE0DZloQgof668nJ0cIrE6bT6Lz
fIZzvAgvTFz0XOi0I83cVRsSemKBYiTrULgh/vqCOBSspqkTyOzV5k9YP2sP6HOEVl5qrrWqrNun
c8ppG+loDdlFndOL2qqaABO7yVY1TO5aEMQSB26TLI6tHZZ9W7yNsf7rOo+b/ebFGoOQFu864OgQ
iRN8T8d0et/nMkDiu2Enwdnjka9u2YmrW/Am9lvPQBVOvpiBVrbqBPREMZS7EbznDL31DSfN2n3X
ueWmK1VHwmECzIW4EL+szADms/q3p4ejjz+NuWcLQp4Rg+FhcGvbspVEp2j03rXKauageExQ8Qw7
RQlbecT7Zn20xM2G1O7iTXhcLg19mWHWzPNvGyF8bCGbF2YW9NtBILgYsIqfFQQ1b/CeiqL7FQSA
VSavFlnQq1Xe+2fZ7OYyohxD1erLIHmDxRZeGGSLlyJYbyOw+agLLk7+tUi5aS/xEaPf4TiX0/Uj
LUf2j8h/44GQEXgok8+jhtEKKNb+x8MRx2CH5TSqmihf8Ig/vDipyYdCzePj6HJH1ACBKX4Sj4Pt
DpihlnFT6ukffTLgqG4HzgDsbBNDSawbWJfjWkYLys2yJF+RuRc9QIPnoRpky2Snpxjt8Yf1Ow1L
SPu7zkmnzm/4/nJWNAwJ7gwHN9rb9GD4G4YN1gPnt6uBrwZRcZ/6rTKmkIS4Xc1codZA/Qi2r2ah
Z05wt3fBaUgYJ0u2pkr1uFj0y136IHBCoepzv29FSvVNWrEcFvAI5GC9w3u78JiDBiG5EkL8e0sz
QYM2+vZmGCqZsgLpeEAt8u+C9VpJi15jzCzTobO3e/U2FfrdWp5IyclCSm0PmhCmfpoXNmN7ofhb
YqakbfCy6zWbvgh064FOw+PeS+G3IgC10ikPjOVXAyZyMDdzC6zRv5fHpWIOA8YwFW0d+4b1AoFx
N5Y0DFTWPAqZmm6jqdmwzy8HvjT6+sYSTY21u/TmaxPfDVRCW65Rqf6TZnvg5DEy+au2EF5jLfAs
V9NqhIiJUTSraI6K7Aeo0omavo7C9V4SYlJpbZ92IBEaIyw6uPilsNMoaQ7PijQlvYfXxQoAavYW
MqA/5w3h79E5Cvs3toiiqO6l5/GolFh2DKmgEdvluPEww3jvWwfmrT2rEUjmyXhUTdLaXTonmJV/
Ct6rVaCYxZAshN70dxMvb64svnH4MbXaNiO3CE7Ux2a/x0VOTU5sNGaoh2LYvY6n4UXzHxCdQMk/
ttXmFCqQmiBppmhp1GlCjbLbkBC6zQmUMUsF6qdSz01hEvlcvQAKgIaKcPYNFhAOIDNY49M8YLl0
xpqKoIOlSFlbh3K4TuoT4jBHOLlWCdEaVexidy86yIZ9mtF2Odn/1A1iSv4yjWH050rt0pRSgWYk
xowvV+BITM+DEca8CJkqy0v2iIrzwRROyQxjzxICi5yrZugCNn5fiTGZZSFlpkphGXu83xrImdD2
I+/L8w0RmjxXC0t1oT25KbWIYT+yKa8uSYfgaCjxcZsLcxhU8dmOznh2uDU6eZCwUtyRGb98DJXu
QSdWbXJgflSX/k101IZ8LqNf9mleAq8sR+BsvO6GiUlV4ALRcEFBvjLfNWGPo4XdenZsDwlxbPwL
3PjGeVX+CQyI+Zqn+gU3+YkJTp6TpF8jrjVLxvoh7TBlscUd3D0jtHrNsB9aKNbIfsd8dz2DskFW
ofbs9unKuNYCeddV9bdAnOvzWZxv0pwra9VyheEIBILSnQXnW1tTDVJOvzliTZG0f03i0Ig8gME2
Egm1Voh/et2t85nDD0hfpK8sMK03qskBdPec0E4hZ931zlpmfIVJYLW6rhS5XZRmo7acNCQtDlwH
cDZprIapOKyMrmbfJo+Tm7lMlGeuBMM0hxA+tadjvXF0HOmstfvwWZzzzBAyHGVllwp5L5SA5dg6
Y73xD8twApchfndP1NlBTexyunRa9QpOyKBUZ6CQ/pbb3qOEhmJV/38ZokKIOS+Kfe3KbZ5hC+W+
ZvUeoSOWF2fszmTxiSehKuew3XWbdPwkczpeYqOz1THZNZtsJ9OD4Ulv6yKdvae8KoNIh06EQW6y
aVF2TzFAty4vK6jyYJAx+R5WxpfLh45wGn7ArpZ0vS2Y9po7c5HQ2MA6RmS7uwaa73EaLq5vvRUa
OdOXNFolrHQv3zDY6cFqN6U03jwWFdeNoK7GSnY2xuHw8Ipk9yFSoES8JCHhmrRG04vNri/22ee9
bc3hb8bVwhp7kWwBQSnx6ORWJKIucap9UUNjplFVMgMOscOBuFgbijHP9z+CHXxYfrYO8rngewlf
pprbo3TMqHn7ZlMzQzHWkpFp24WeJ4PWrCQcagtWHgQneymrqur9tyscBONALogRUksbtA+YxX5O
i2S3dcNWcHLAQcurtPTbiv3y2m6goi166x1UzgnHYSIQZfWcL4vL4HYe4EF8rq211DcjgOmLTSmV
q+FUwbjMzsUDTHIRsfsgP1l9SsW4tosG7IKBhrXFmQhmMMQwMytaNAeyO9qefrTTMfJwSQ42fyjK
fWiMdrrDhrkH+VcvakTa2GTewwD3NeqYZpkVnivJY4i3LxUoRhsTQtwVxGu/bHNtwdzSJnX1eVWg
0Q2AOUvWGhv5O5Sg/Nc0SuC1oiXb5ZvWxSda6yWIjO6874oCxK+ALJbwyCV6nI0dy6tHhopHR0yj
m+PoyegAay9263OF5F0p2EIpSDUwcEd/Ijy349SL/BatU7hHF3yCY/mldpapPueNjbS78sMFduMC
XvnG9WuG1+w6f0cTVnhOg7hdHqV9I2hmWWwfApp7tkoDpPRtx1Gxilqbzm8LNyx+fcnetc2ImC0W
BoKvRcOm+qjwcGI1m56F4tVEGMl/dl4E+kThHapkhMH/oPSyGsz/OURfB1uLHBGsi+8ylqNahejF
MTIurRhvmiJUFHkBtcT+UhK4EChOSo/KO/PPma7zor9zgJluLaKme/YA7okF2ngZ0msh6F6e9RzX
Mo95AKwN0MdRMYq0rXHNlKEETjPVfEGP45OWCiiiqQ+tNDHjDAZmUpFmQg2+E/QhArCAtkrUYyBM
6Tz5IaWgVLwfrz61Uaz81SUu0IqLOZEL3v6r5+jcdJ8DvsprIK16JIrysXZ+Z96baQ6y4HeoXo0C
jeUFGZcRtAyVeOhhWU+MBHJ6JVJjBV3Gxcw1QaohxYqTSJGTK4Ep0TZcRcM1nxR1Cw8oOBvRUze2
XFD8+573r0WnFXtyzUNwoxExowsyFU65V5UY1QafVrL9pjv4UT09IOuiMlF+G3K17hMhlkzL77GU
Lt+aPTw2BVB/7EQO/VGPKAbBRPlxNrsGsw9uuCJhMEUSfJzokLCBlsV0VCLVjoT0v3T5gSDV3lti
vaMc5uZPAQLwxywHHI/D8CJQTCHKe6QPyJ4LIMlbXB3RDZ9ElWlFBtS/FMUnQVDB+L/oFsnpfoHz
A0MU2Z1lPwPWymbhthJu8a8i/4vD7U+PDgVkHBNH+8AidZoKHKWbnPhzKQ7UxonjGATMpOvaH4Ac
PfskSl4tkfvoGrOtc12TuunGmKCCEtg/ExTCsKwTyuODNRE0J6hfRe78rOFmQ8FJ9Lilz4F86CyV
jVwygDXCWeBVGpIipy6xlDnBtN0eQfOmSJIvohFjfyFgvHZPppAvWHWjqEab5WXMknNd3z+NCLI1
bCf9M00pK3k1Q9PufJUDqQOH9AW2SZfn/tdxT8u3t2gg2mfWn/WGPW8WifrLJwxFTXYK
`protect end_protected
