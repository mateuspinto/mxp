XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���	�,��~�H����r:��q�,��|鴯c��(7NB�A0�Ɣ�����$�A	k�h�H��%�^�b���>� �҈�^=��b�h�ZX��#R�+1<�?5�rL����ZxPܹ����A���ub�g1�M��� bc��KZ?̵��Mc����5�+^�\�b�n�e��[��$�W�����	��fǥ���y4�Uٍ�Q2!��0cn�"<���Z+a/������N'F��;�r������m�{����fm���6<��>� ��C�7��F߂d_��� ��;�������9A��a�!c޴O�·���m�አ�Dp����YP���B��Rٽ��+���W��@$E�^�o0�;�<M�����oX�s:�պc,�"���
f|+?��\Tz���=��LE�#X߉�x��
�E�ұG����%�b�*�80�Jg��l�w��LQ�׷�6S;2.Jg�L?�W{����� ��s��W'��Ĩ ���@�-1(�;u�ƶٳ}uRݜ;9�nѶ!��-���w�G�}�KT;�/Hٙa�Z�8����I/h�u��4H���"��p#��Z������c�oE ]�t9,��m�Ō}?*j�2T��<SlI���Xy�TQ�w*�G�L��Z�Qx���o��vT�vo��[f\!�}Vզ���R	bf�Z>���������vO�s�?P9�{v�hiZ<��_t*��И�Ƕu�p�p�������/E�2E��2�XlxVHYEB     400     1d0~dJ����,E+_W�N!��b��ފ�t�ӄY)��A�.�0�*��3E�L�z/o#��)l�x��ϭ�L�� ����x��b�_#�������K��v�E}����G�
�(y!Ns�yZʌ�������e�g6�`����:dl§e�J�9�� >�9c�����	�<��x}Tb����;|-�S���V����C�����$�M�d�E���:�ɇ�u���U��cGG�f�$���{a�b_$���G�1����r���̉#�Fp�5��~`���������yr&�.t��S��_��/D�e�;̡�ܽ����r�]츼�j�mO"oe)� j\���7����t�c������3s����.�Ѡ��/��f�aH{�~� 0����[��fs���u��V�p�\o��.t�cY$'/܌3��sJ����t�r,���^DdlLb���?XlxVHYEB     400     110�+�[oM7�I�\��5=�\%:	�Q��
I]qu�"\S��wc@񺶀�Ϲ��t������&d
�C���̦&-��ѥ�[���'�vh�(c��x��uC�����E�t}��"������:)�*��]��j./T�b�͢f���k��Y�� ������B��(xՊ�8f&�����WP.�>>W?��JL�]�~�E���j��jfI���xkǖA��iy���>��:������I�C-��@���̩O��p7�x����XlxVHYEB     400      f0D2�|X0�����F�S�� _���B?X�D�zs0��75I�y��_���eF��`׳ ��;�2<�sr�M?�
s�����)kq6�L��;eM��a^�XF7��K4(�'谦���|��{�DuWm�ݖ+��1��2H�&h�=�hz�J�R��8S�0�\.�`�]�sۤ6G(��L����H��v�9T�ץ#���<m��"Ev��J�\k:�zR��r�u��ݬ����XlxVHYEB     400      b0#�ADe���p���T�����4�(�$q�he�{�jD�z��ASB��_o��� j�V����h%<7����xI{�$I������]'���#ͼXv��#kK  $��?広���*��E�(WQ�9;`�6ng����u 5o�B6�P}ZwA�$�̄%%�{���&K�qH�D;�XlxVHYEB     400      d0O�
5d8?��i��s�9J���;F^/	�f�̞���(��^v�p��ER�%�y
։Yg_�<��ڔ6�c��,���۹iP�O
:�_#l& G�&���P���Db��ͤ$�X�T#��$8�!�<c�JTۄ�������O��R��# Ys��<FL\��Ԅ�FI'�E�~���4��S�Ϳm�i�ah��-���|iLfpXlxVHYEB     400      d0^0�Ͳ7�*>��t{�5�k�f�c�l!>Oly��q}�(%S�R7���庭��׆K�����0�C���\չt�4f�#a�SڄP42	)�J�C�����K�v�Jkn��2��9�����آ[�D�` AY������)��v.���Q��1���^< Ew+�85ݘ���'7l�����u���b���@8�s(�e�w�ʶ����3OcXlxVHYEB     400     120��� �I{����Z1-�|��:7�e=e�S�ۇ��� ����hV��G P��\g�'w^���ӹ��I�a��a����>�>o<���q3"��G��,P��G�X<z�}���\�M5��qQ,>x��o9�O�sD&��s��s[m�4l�3�Yz�a�"�;1��4\Q�`J�N����r!�`|��~L�o����~�	u_ᵱy����2)�
�>�!I��W��."��f������H�ߛ�� �A�X��A $t���Ӌ4�Du��I��>�"dXlxVHYEB     400      b0x�s�s_L��C�[��#�-(WO���|l��y�4۫t�a�߰�|�!�o���ƳōF͚O��,\�r���އ�&�x�C����ӹZ�C��:]�:ݳ�S����b�s1*��kP��/�E6�Q�Ve���Kh��@ӈi,�#�5�Cg�o��)<x��D��2��XlxVHYEB     400      a0�e�9{D����a��ʂO|�Wrd*�i�Q� �N�-�\X��v�8׼�}L�)����S=�6���Mm���]h�w�v7&��W����ㇿ����}8ѱ�y�Nz}�(kxHQ��,�z4�eZ!Z��Kf`J��9>2p�aL7�=6�eǋR�d�BXlxVHYEB     400      d0�l���HC�%H�)�΂�*�U��en��)x�J!b�m>��3��b���o?��{���墨b-ߙX'�h��IV�(���GA��<��� �`�M�����Άd��}G�Ĭh$�8�ܮ���U^��(IP�\�a��B055߀�R��B9��L�?!M��q�2���\�4�T5���0�9�\_ដ��*��Fi�(t��"�u��	XlxVHYEB     400     1809�;��0*��G��C�`�+%��",p�L�ma�n�Gcl5V)����S<eɩ�0]V�n��{�v�
cA?�ܓ��z҆쵻���i�a��p{��{)ԁs#�+[D�s!6\�T� ���b�s�I'~{U�wc�8�ln���ϳ�Z��C�ú���PqL��fB)�j�}�fF�s�����G��A,0tha�|��5^H����/���(��X����LSC��Ԡg$�]����|�+��A��W�^�]�.*��{������WcE�1�X�%�J�C\B��j2���c>�vAR��"b�0a�l��|U]������FPs��#���Ho��)���KL���{�is��UIp�g�߮R�)v���̙��u2���� m�XlxVHYEB     400     130f�S7�P��)%K?�cBb��Q��������}��bv�}�N�H$���p�ڋ0\��;yU��ᶢ%��^/�Е|��pm�9#kѵ��uN����~#�h�d`��?���R�B%�W��E�N)��r)�.Ji���c���K��.Z�͗eJ���x�U�v��b�:7w��V#*�(�\0��%N�~���M͐s��-�J&����bq�[��v(@#Ǝ���7���]��ZA��zʎ�o�'�|u`�a����K	Dz�7ʭ&��Iɺ���F��Q���\WM�@�XlxVHYEB     400     110$ڤm)u��R�r�8���Rn�a[��G�1�x��L�ºu�v��_��Ч�~ՙ������#[ӊ��i�'�Z��1qC�ʽ�`�Z���o�6B�K�[�@S�<�A�� zHfk��'^����;�\�i��*���*�.��s��V�����c�l	^SSa{����=�7K��&i�^�KS��TG7?�8�x��'���X�d�J-��U�,�r�
9[M�/1�:�P0�N��{�s��\��	��)�#�;Ggّ#��U��ПXlxVHYEB     400     190����sZ�lZG�D���ՈQQ��
�L9�iB�%�w�V��]10c�k[�o5/���2�gd"N��7��*�"�6��Ii���.S��a�s'r&�P�/`�C\/&Nw3Z�=ĉ:ry�лΖ��K�Jjr�5�N��N�Ԗ }�<�A��ۦ�IS|@����{�7�^�1|AK�Ȇ�R���UB7� H������)����ʆ�w3�N{��{ό�������&B��� ���Rd��L���-Wq�᪍.��- ��z�١8����/��q��e��*���"]�ޣ�č�a5ʂ����t����,���A�^ڇ�2ݩvI��4/KCa�H+��xc���k�řc=a5K/�؋����R�'
&Pw�]��A�2XlxVHYEB     400     110\b�l�$�{y�ݛ������uϲH'hO����Y �id2J�mD���8�x�~�4�j.��^|�9�� m#����fJ�r��'r�E�S���W(��b�i�$��$�p�`k�q�� �����uO:;[�-�"
����`����υP�������`{��FUln����F����&AEC���aWk�bh�P(���JݯQ�[)G�w�&�ii�E H��@=_D��B\G��r8�#�Wr�C��Q���=A�$�C�XlxVHYEB     400     110I}�@�-��=!�)MpY�3zJ�א��Z$���#8&����ad󨷵E½5�Y���|z�Ҍ.�L!�x�
����&�M�2,0�����L�M���k;P��<1���">�����YM����TԺpw-!;U�
��|�.3�S����z?�~;`c!��F(��Xbm	�p������}s3�ߑh"���"�^ErڛDd�)\���%��Ew�s	Pj�*�K@�t�a45��b���?��+
G�8��	�K?����XlxVHYEB     400     110���A�1D�@���ⵜ����/����|�*��yc8���w�(�G��;)��R(v3JP�F�8mׄ���/��Z��p�!�*�ru�P�Q<F?�`T�\&�>��I�k���ua���YQ!�NTh#b�-:3�dD�h*(�MX1O�?�F~��TT��I�2M��Ĭ�bq���+ �Q���qM��\
�9���5�8_8,��p
G��<B�%�����|�n��Q����_���;���E�b����
�氀���G�XlxVHYEB     400     100֭A�J� ���A4�gC}چl��5
��[z;[ߎ�.cɲ������H�Տ�LG��B��!vF�������F�p6�^�si�M�K�����<��ӿ����lܕ,Á P(r\Q��(迧=g��s��/׉xw�Nu�c�#k�'� �."9�O�o��cKƗMڤ�q�ѾΛ8����״͐U���Fײ�-E�����|����JExM	�wU�\<6�'�$�[����5
4��}f�XlxVHYEB     400      d0�P��`0N�yQCu�C��:����0�"T������Ƅ�g�E������э�&�.�L���%�t�NOc�܃��X�/v�HN��Ȏ�6��D����-��T��;γ�R��;� �d�F�K�^�@ob�_���HH�L��-�>�6�.�����)ݹ�7ڋ��z-���ۊ���T�ʒt��m +��8#
ǹ ��R�g�؟XlxVHYEB     400      d0o��=M\>%}<E��ƌb�t�Ơ�_�YmF���W���Ք-C�ZH6}8��W,��=�?�sm�����^f��N"��o��8IG�N:�L��1��ج�@���m�	J�6����ux�RU���U���Y$�H|y<��H½('� թ8�u�6>:��C��)�VMnK����\���E�$��c��R��h!��XlxVHYEB     400      f0���iU�!-���l�V�p'Y�)iR�Zy/�.����Gx�oOB$r�P�t��[���&њ3���$�N*����E�Vi]��Y���9ZlG���.�0�rG����SZ�9�d���]�T/� �;�$P�{�.�B�q)M�f� c0�{�-�X]%%SX*k�$ŗ0���j9�]%� ���D&@���[=��(��yH_��6�M�ӄ
>.��������%@	�F�'�,�E$LXlxVHYEB     400     160�*�?�h�VZ6�e�##��=H��ٷD�H{�(�C�2�4eb�k|oCj�]�u�mp�[�A
@��Mz�n�Y��1��H��
7g2r,4�!�����a+;��Kg����J��������I�DH�)�]5��[���{��b/��-�-���+�F����Ι	��<^��HH�E����ឆ� ���%o��J�zҼS͆f/�&��W��[�i{�$�E�ȵԼ�5�y�~c��U�+�wZ��`5\�pH�B�	 �����MV̲s8��C_Č|���w�;���3P�EF^h��3���! ��piWz��n�%be�0��h�'�!�A�u���~����XlxVHYEB     400     150���E���b��KV�Ҝ����
)E��Ogj��1r��L�T�J���Ѿ,^G�����|���rf�WW"���.O��K����E�����9�Eb��id�����~����g5���4����9p��@�%C:��(Y.e����YnT���W_��ȓ8���;LH9�q;��}�����W�T��: �2De�L�0��q�7*��Y��R����N�|cbe�f��,!�3�>�%���Qo��T�(4�=�E�\�C�R�H^��ȝ�z��[P��\�3�}��-�e���y�}��v1f�}y3��I���!�!۶Gʎe�S��)�+UXlxVHYEB     400     100S%>�F�k�\�Ag�.�*�+g�i�P�Id�ؽ�$q��rM�2��0���R2aAgE@�y�Ɍ}IS1l����.�����!�Ͼ���u	c���21
�1�)�?��e��8P8�	�����xXϾ���ySB��4�ڙ��T=�CK�(��@��E�ڋ3	[֧P�*V��`Ӓ��B�=q��U�S㊼��#�ꋩ���i�EG 5�~ljj�������q��z�VT0 ��Q�O9"�$�>�XlxVHYEB     400     140k�̇7���MfvU[��S4��A!n�H�B�>!��9��K�����zq�I�#�Y_��)3wІ����aPh�
}�ԚG�K�j];��e+�$uNM5j\p(�+6��m�zM��wM�_b��pU��m�wYkԹ˖�Cq�)]��"�����1�#2膰7m�����zC��,"#�fT5�7��.�^�6"�l�]��p���u��e0\R�s�"C��8@��F�[����bW��}ؽ��TKcziKP����d���0.&#=2h\m����/:�=%И�J��D��i\��.5Y��V*�S��!���XlxVHYEB     400     140�&��}�8�ë�>��y7�'�e��R�ދ+Z�3$�� �B���F;��Zlg.�y��R�ؗ��T�M,���Y���|�)A�XF�B`w�/!��ć�.oj��K�3=�T�r��d�9#�b�?�F�
P����ӓ7l.�_��	�������y��<SЕ����|#uq�̲���O��ĿcA��^���@��	|��X�̀����g�'��%u�X�' n�'�}�T�G ��<}���W�.q�Ԑaa��� �Z?�	z�0GU�@*A�ȶL��M�;H�j��������`�Eg  �[���XlxVHYEB     400     130�%�{^xs�t~FF�� 9"�S�KN�D�hm'�o�ȃ{�/@� ��Q�N_m g���]��#��HS���,��+�˿0=r���4�_q�㵚C�ϯe���%C�] ^jܪ}�U�I��b���'�����1�ݿW�s ��j� -Z�l��2tp���2���(��_IuL�0F�����h/�2������p��g��S/�����E��-�������7P����}�XĐp�b[h�����,PC.B-K�b��͛�?3¸(��*�!�T-���f;"4
��<��s�iـcVXlxVHYEB     400     120�b͍���֋����5c9�pe�c/�����e(��64$��b;��Q�o__=4@��lbM�� k.�+��=��j�.M5�Y�sc����8	�����%�B҆_�}A�w��i���2��v�8q���9��*<'�mr7��4[������C�$@������ă�H�r��$t:֢�{�Q�����X,ǽU/F��O ��-���.m��G"p�t=��zꑤ.�@�z�!ŗ����-.)�ɍ�/e��v�����YO1'A���ӂo	=Z^�����ǵ���̉�u��XlxVHYEB     400      c0��]�U��8J�:)�L�}/݈^�T��X��7=>����}-�����k;Ӹ��l���b�TDV����<t�o�L�/�f�TY�h��Z1M����5��q�M�� 8�,�7�g(�����[���$���4f��+\������Ϝ���|�կ#��b�(=I������k ���� dʏ�u_6H廷	XlxVHYEB     400     120�����޼ �B�6��b��s�&u�6���w��Z�9�=�����Ҝi ��$��S}w����ǽ�!���*BoΕ�U;���"�
�|,:�
���v��"=���e��
�<�.�e��mgM�"�Je�����ZE���k�g�)T��;�`-�7t�^��5 £�=u��<Ƭ���[�)T[T�yD�}�R�p�z�|W{g�y?�*�<^k��T�����W�_��������u�>�>�n+0�v�a�km�;!WX����,Q#� �n	��9z��XlxVHYEB     400     120�C�և��ͫ������;�#C�w"O)x�D$K����N����膍+󉥲u�5P�Q��ei����m�c����~-띨��UHm�����1�-w�!gV�&X��u��Ay�h���Θ��"�~6�]DGic� ����#�MA� ��GkT.�����LE��T�y��0uY	�5UP0����B}���;�>2�hvtp��˟�H����A���KBL��,��D���>���vCZ̥��=;3��:=LX �K�M&��Ti�3J����J�����vXlxVHYEB     400      c0fw�۟��;w>�����=�Ct�׼z��9�6$%��s�Z����CJՁ5���;��ّ᷒ �؎9�1Zy����l]��W]��6��ґ������R>��N��̛K������쀂�Kn%�U���j����s��� ��'�J<Q���r���嘹py�?��w�Z�[~�~��k�3��%�6�GJ�C XlxVHYEB     400     120��E�(d?��e���}��7�v��Ϊ�~J9�ϴ���A ���c�$a܋�jI�Oq��,I�B�l!�GO͓�Vof����$��˚�mɏ�'Ğk4��O�����7�Z�j"��F�$��h�
���{/b>'p1�dOr�qO�.�(qUj4����:��\���2�jkFpPe�>�"$C���Z�����5c���ai�2:>f3��z����yf
7�OQ��1���Vlg)^df�ʯ���Nh��N����yE:���SJ.�[�hn�U�g���'�XlxVHYEB     400      f0{����.}V��4��P	��va��)�g��DFz�+`�O ��IK���% U�����k��KJ`v ��q��=X�G���Gb�t"SL[�>Ei�y�l���O������}�50�� D���=�q/�Z�REF��<�6tSg����J��b��Q,OAr�37�^�t��zD,��T�e�qu��zC�>�5��c�pΌ��Ou6�,^������zq�V7���E ����y�Y�|�XlxVHYEB     400     110�ȑր�A@٬lqٴa7�#Lbb��N<��ӯmS�׋z�ܼb[�U�#����<��z�n%�����T�$�ї(�8��v�W�JV&K�x��m
݁��3��0i�tj�݂Iև�e�͠�y�Lb~ـ~^���^�J�D>p��7��� V�i���V���C->�3���96�r*��K)�p�0sL*�|U�]���KQ�e���"���T��}%v��ƕ�M�H�_V܈����ʍ����$�jyCH�b�<��ɶ)#tXlxVHYEB     400     120cnV�v�K��&����*�z�E�Sc#�_�[Lٮ>�|��t��S�'�t0L���aALyՀ쳎��<����?$�]�j�tC�?���/�0�qW3�0�����7h�]cp팪6R�M"�
ݦ�WD���.e\�/��a��,âcS�k����Z@���q�#����C�|�>P�� �{�n?������P��쓰ݳ��y�J���C*Y�J���� �:U���Q���=aw�����4��D�
*t˶d�Bz+��Yi�_�LvXlxVHYEB     400     1205��� 1���k:����fXV�T-J9s�Ն��{��yv}�}�.�]�Ov�Z��v��t�w���
é,���)� �}+L�2�w��/mb6b�&/K|�[Ϡ�A9txw�Y�}�A�U�;EI�	��X�ٲ����v���yB-��I���KDD��:$���J�ę[R#���RP�?���ߔ�/]vy*Q@R�rK�:������w���Y����l�u�%32�mh��/�V�vO�N�4K���Q����ư	��	*xی�{ο^r-c��t�0�XlxVHYEB     400      f0�$��X��[�٧et�M[n�Į2*�`�bp�K�Q����\�y#�#�NΎu��_�z�QV�F����ʴ-�}$�%���DC����%��M�Gz�x�0��(�5o�[!�E�?@�#X5�)k�.!�ϰ��sv�.N�%�Cx��]����ej@��8�l��HvI��O��{���l�9��J��Q���V��B��!8G�%F�����0���K�.���i�/QG�0>���]V�V��#XlxVHYEB     400     130�/L�@h��8�t ���_�GR�خ��|��a[���ik����w`��e)<$����`���]/��;��-n)��+$l(�z�91X3s����<�}t�n�Ã�\��G��,'ٳ��d�Q�� ǗC�~X� ����%S�Ij��&@�ܬ�i��wVh����\�`�E�ʩS�����O�bv�d�ת�K�q�q��v�׊O�� ��<��QI^:��2E�l�p.��fuj��ѯ�sb��������^��;�4g�����?h���ˤ��3B�Z��x˛}��rB"��9O�4XlxVHYEB     400      f0؟� ��L@HGGO�5���MF�xI[�G5&m�`J=��V�S�Uy���|�3E�iZ|�9d4���g'��� 'cU�g�iZ�m6��S��9�V������X�EД��t�x�3�oOp���o����moiM@�t̜��=��+��|��c�X��i�K
?���c��2F݀�zi	�Lhf��M; Y{�#�����i���)νĒʼǫ��n�y�P���T#n�XlxVHYEB     400     150f��<.?��<Z�/U\��`e��S� 0{��~���v0��"��s��_�H�'��!D�>��!���D�']c~�3
���%�h\����n0��n���o����
�rd��ޢ+�ј�����Z��|��ޟ�@������Y�]X�G�#c[���������Ez���~"�+�i��-�\��S	O��]ǟ�t�Ff#Ch��H\l����� Z�`.���ی��앺J��
o��3��Jj��YK��
j�GW�IM@;Kґ��i2�rAZ�/���[�p��ʰ���c�"f���CU�	,i����V��]���-�"���5H��XlxVHYEB     400      c0;V��|�t�!���ԣ@�z�ǌƛ^A?|�R廒�|@�.��+mO�zXIl# �(qUȎ*6tC ��s���ȵ5�>v� ��*�B-����\�}����A��*���[���c��u:	���V]�E$�5�^"e��ri��X���$��ǎ/�	�x�9(^ [��lO��F���7"b���3�X�-�;�3XlxVHYEB     400     150������Eѧ�����z��f@�sC� �6��!�F�cq׻C���=�2�ߕ�Kpf#$#n�;�{ޘ�c�=<��������<$�� ���-�����=��
'�D;��T�>��U�!��b�s&H��6��
�\L�3:MX�ԯz���BNâ�I���Ĭ��[�e~0�� �ݍ��M3V��T����T��Ak\���w�L���ywZ�ȻX���;6�0^�joG$�Lk#�z��P�]~���|bO�ofz�<�!��"t�Is�$����=e�̎�!�7:7ΡD�1# JsJ�L�پґejMh/��?<LrZ�)����=����l���?4$+�XlxVHYEB     400     140~�ٞU6
S��r�2����^k�J*�q�������u�5�H����9�ҿ��7A\�߬���2�|�4Vi�@+����5�BS�N��T�ש�M�m�z�� |���c�x��i!���ĥ��2q�P��q����Z�4� �LѢsc�̔*q#�䯋�朷�z,�Y� V��˾�$��� J�������6$DS%kO��Wx�,>���"*~����C��!� ��&����\�6�L�h=.lA�v
�Ԧ�H���Gs_�P&đT`Bej�8:m���͎Ԏ:k��W�J�F Z�'I��L���XlxVHYEB     400     100�1�����rs��&��S��|����@&�%�ۯɽ��^�(ш>)��vN��RC����/\�E>{x�"h�}	�(���+��:�m$�;�G��ɿ�B�Sg�佝@ھ�ҏfxLj*;R'����k�h���C�&z������H	��)>Y<̴�إ���@ryo'�*`�q�j�Sv2"���s2��#�ً�H�a�$,�9��"�^�M�6�r�J9�x��Y�r)Ħ���i�B"��YV*����5XlxVHYEB     400      c0a�Y�mPq~7�H�S#g��+?;�r���P�.��TFIft	X��f���<oS��M�}Z*\h8AiE����>.l����e���4.T��K�_�eK|�K�j���wJB��q��q<��g�L��xڔ_�[Ke_��?7���7��T?Z=��*��@��I�=�5���B�Y(~��K�c��lL�M���H��~�XlxVHYEB     400     100�p����;c N~Q�n�h)������PX��5���x0N@�A��_�s\�3��͵�4q�-G��s���;�4!z��GK�j]�C-x�B �L6�(���>�߹��4�+���c�ūv+���(v˰�5fJ�,�_yJ]z�G������������V��A��;o��g`"�E%0�b}���¿��&�a�#��b���Ϥ��<@� u�△�P5w���ӫ<V�U�Pz�
@�L"�Oc7�m��~��1�XlxVHYEB     400     110%~�b��o݀BB2�w!��zpM�3�S��!ʽ4+2S&U���f�(��(���wT#u�w҃]4|u��&qU8�ՆN$sWv����%5ǯ�c�	�&h����@nc��r{����ӷ�g��<������c.�B��8a[)�X����S&�y� �vBƐ<I�O:���|E
b��4>�}�r��I�_��J��;F�+M�-m|��[�]z*�A�����V�_l�<�;�+���0��'M2���d�dσ�c�ߌa?5��VE��XlxVHYEB     400      a0#&�7j�#������d��u�?�{�&+
��-Ym��90T<�_�V�Ϸ[n�顇곛�ߍ浤��ǭ���ľ�����kن��/�fN�����8���R��/������p��{)��V�$ʒ�jqT�>�?w�gY
/�5�mk��¶u0�v�}�Ѡ�XlxVHYEB     400      e0�w6`J�����ۊZ�R.�@�ΥԐ@��ٱ�6��p�CX�Y���x��:�4,URR���G�A��0b]j�y����d��H�l\�a/ŶJl�'�k��\({��š���0m)G,l�C
9�	?��c|�%Y ���6v'��M� N"��1����(/6K| ��mj�R�6�QAu��G6 H(	2׃���vM���)b��ݵ�*��a���!��XlxVHYEB     400     1a0�k�P��k���+SNΡ��;5���4�b�ZI0LS*��v%�����Ӊ��������=��Vw������D�+(=K�Ѓ)u'A�=�~V���Mkf�]'�2���h!���Y��S��H2;SaOġ*J�(QOWk�rF���P�p;��5gU*��%�歈P�X�����
�0��5�*$��;o��a�ÑQ��3���ʋ��foʯKro��U�՟@Ή6��_e���3��Jx�'�-�$�-�$���� 
N��	;�> g�7��J��E@E��  |��_{ؚ��|A��@j�)�s|��|����"�t�#�2%���Zua��aq�CE6����)4�Y`��A�&
UA
H�����>;�?О�x#�x���jB��̃�t�"1�jL�k��	��ª��(Nh�XlxVHYEB     400     150{�&��=vЃ%�p��x�f�X� ���l�̳Go��kR�&�'�ӣ����HD� W:��y���:��Hٙ��/9�jV����>\�*g�G ݁�Ĩx��7���'��ᕝ�����V��8�W},5��nn��:P�)��Ҩ�;�����âED�.�6|b{��w��e�\�S��~$��n2{���.��p�f%Xte�H+>rG�H;˩&�m�vwϰ��O�~&W��}�
$}&��:Q�ʾ��w"�[�
9��������X��k������?�>�#2��8�,��Ư�&��������֛��2N=����_��1T�@=BvXlxVHYEB     400     120Rߍ��}�� 6�s��6�v9N~H�B�X���y�<�Z)e��s�?*ͭ��VHF��X��M�)���� zt�uȖ�os����fõ�d1��_�vW�f�p��<�t.b�����KB���]�͠c*�ţ�2z��\�dRW(}������<�r�o�1�����eܕR�g��r��Rtʎ��5ZX�9��	3�F}B�n��/ǚ���a��y
������e ��¹��>��͉��c��*���O/��
�7�7[��Dπd�= �f�����b<(s�XlxVHYEB     400     1d0�
�I�<����Ĝ�������8��o-ʿ�4g�b�qt��lqܳ�o/a�X�G5L�p��g�h�8'�e����q�X������R�zUci�ރ��KX���Ձ"�����n�����5�.!���<8z<)��(�A���l��ӥD"e2�r���>�3fvnW^Iw�O��,K���|Uc��BU�+�&�b��\���E�hI��]҄xb�u�m�D<��2&�~��.��J�)�����fm4$�j����n�|F�h�ܘ�臱V��(��/�m}����������iz%�kY*L*Oȕ}��0Ъ�l=ǳ-�8�R�GjTJ�%�0A"V��γtM��v�w��U��o [�J�d?ЦY$l���Ǭ�qT�Q=y<��O
�W�\#�f+��	ut�}��Ί�_��i�=]q̈��6{c��Y�-�s9j����l�U�a5 b�TXlxVHYEB     400     120����nǰ�~�F��jB3�J�@�׭�����d�\"�(�e�W�ڸ]����)8&2j�֖��?+�̳a͐g}����� N���.�3�@k?#��� b>g �K���s�-�3�T�(�nՒ*�sf4/0c�J�caM.�K��*P�ՠ�tʖA���\ڄfƬ�u;�?�����
SX$��p�o��?�X���?��J%���v��잮@�v����]�p*-k@^�k�����O���@���:�(��Nvv�XK(���x:�˱�!}ӵ���}��K��g�*{XlxVHYEB     400     100��Z.�
�#4J�<���[�?ַ�9��&����{􋸃H��Z�T�]��-4˟ٽ��)c�g��^1yl؊[���tv#>cįsr/Z��f?o�O��8�?���V43lj��碦OK�����h�`�Gܬ�:��5�� d=�c�U �l.�Vz��2�rTې�+e���[d+��:hC��×�bB��Оy�ϛBǩ�g{�"萚�=!z�by��	��[�2�qt; 0PM�2a��~�F;ܖ�\�XlxVHYEB     400     110A5+�(&I�Q>,)���ծ��_St�^UdJ��	�ڜ
��Re��tub���S����[a�t�+>����>��V���mM>�7%�̦�r6yl��H9�w-���*�[�f�Xp��̮p��Q��ِH\K|[R�b�:�h��g�Q*r�O	�ę��'�L�ђ�I�C4�@��]Q:R�J`�,<k6��f�8f�����W�(F�4���d|Ր��z�*��&C�H���N@HJ��z$c�h�Ts��2�?�WTһ��%SXlxVHYEB     400      d0=�ӥ�A��ҝ��h�e�/��Aw�a��������7��y��+��_��1i��x��&�ϭ�6vt��!=����i��/�Z�Ha��ޓ�GH烃ݨ�ē�]@L�/XO�����������{���f6�f�.��Hk�Χ��ns�%�� �&��/���Ǆ�S�����oeV0$�vv<&�*ߌ��D4|0i�XlxVHYEB     400     100SQ�ov��#[K�P�H0���sJ����q�q)�/孯���y�&/n�$�2]J���,M��qfi	s�6�����	�T�F�pp>�Aju5&�Gs�D%Fq���[eW�pJ�fLE\�S�-6�鐑��Q����eN� gC�]Zn�P?��ྒྷO�l��
�$굯�'k���s~IP�B�}J4�h��V���0�H�4��g�_�c����0XF?,���j8{Vc�isxkF	��L�2�s��h�L�"���.XlxVHYEB     400     130l:H$i�j�e�/�p\.CrdT��u$�B�\�jU0�Fi �kCN��t���Оy8;+���U6��()�2L��SO�&J�0*������#��*���8����%� �K�B�A�RO�2����x7��0%$RlS�)��ֲ��׬�K�P�������7������;���z�\o�\�[l�D���q?�!��@�4��!��7��Q�mO{�6Zɥ*���#p	QG�U4��{z5|r�+���Q��	Q�l����o�ծ�\�{}7����A:l��q��襘�]��L o��و�ЬeXlxVHYEB     400     120Dk!��n5��m�x
�h*���m� m/�u��������rY����3��!Ry.��Q� ����G�(Ƥ������
n�QӅV��&����;���}�}j����@d��;�N<�m=�c�8T{��
]�����B�jf !�yf|����Y��E��o�0z�z������1�����L��*
Ol�J�4!?�$g���m�b��%F�h:�E �ag0;s_s��#� �»qO�j�X}�RzpXU�_�u���G&���J�m�A�W'l��4-�8��_XlxVHYEB     400     150%�]}�������cV��{���E��_��gN�!�6�bS���&.��L(ׄ;�Bn�ELWq�s.� j
��A9�(x1+������V�)h�]-B}�#@'�:¼�:A�~� (��u��uM_#F���xjFLمQ��q�u�!��O��w�妡�A@�k	XK�-8J�L`j[ڗQ���/7���ؙv��w?s�{��������7��*��<��lL[�]�j��8�WF�a�O�}��v�ps.qu N�Ej�T�H����
.�\TdT6�1z`����Ηbf0�Uɗ��V�"���Ĉ,�m�&�=W��6�SIS��f�z�n�#M���XlxVHYEB     400     110
0F�������0OU���[�E���v."��䜹-��6�<���NO߼.h:�t�$m�T��~[M)��듞�Ҵ/�d�X+5|vt���r�ĭi��ô�3QX5��xv�,Z���؞[׺ә�/�a�z����a�_�4���WB����J�:�T5�C03�=.�*���jۺq,�'�#��0!x���?C,�-�'��&_|�<H��國(/)'#�s�� L��^�yhT�^���o�`�I"	�@��mF�|׹�~ u5���qx���XlxVHYEB     400     110ϩ���8�`'Fհ�g��#NX��8�+ ��Q�g�ڙ�(��u��ȳ�D3�k��̛鯈}W�#4)��d%sp29����!�Ֆ�רvY��?���5�R�k��t���g��>�I�ؼX����R��ex��+�%���^������#ܠ�J�;�֘�>�m�/8JO�[�ȧ{B̟p���F10�-�_�,�b-�47���,rz6/������ǅ�*B�'mv��w���_�h56d&6�]x�BAʉ�)XlxVHYEB     400     120�^dqlΗ�J/���t]Pp�r�$��F(�i���~GMʰz���t���ms�����{���^�b7��-��0�ݵ�KN[��_���ߢ�r׺<�����FUpXg�4�Lv)��6��l����'R��6��"�Ey8L������u.,B���W�47���y���[(�A3��;��	q\��W��۳
,�mkOP�F<�r<T�(��M�6n���2@o@XT�<h�N!Ӯ��o��-Ѷ�' �@� "v�(���?Q�j��(���b`���'
C�XlxVHYEB     400     100&>��~P��-@���D�]��Ɂ����ev�
Olܞ�P�6��E]����5�{͕���~֌�u�;��&x��B�����s-Jإ.a�ޮ��)����q#
QT�ɇl�Yӱ��'�Y6"�.�Q��ơd���XNN.��E�5p��4���d}�mFK�_l��rP�VՉ-aEFAK����u6�Y�5�7!f<Q6LS�
�#`��5�C?S c	�R;�DFL�j��J����!N��=9qV����P'�bJWXlxVHYEB     400      f0�/Z��e{�?5��cJw;��"�0}6����bw��ŠQj#�Ǌ�Q��)&�O�(r� ��Ќc
�{�)�u;/1�_4�ZH�ʶ���5Zg���dvVA�:�+Ҵ&vE9v�ه)�S�� ��7G[U�8�վI���h������S��~���Cl�Um��a7<MlI�@��O�?\1Z�r��Pt��o�RЏڤX����{l'���9��HGϰ:����e�V5���ʼ�XlxVHYEB     400     120�lp������	<�O^�����t�(��ر*��Ѵ�x<ޗ�`x���0ޕЇs;9�蛱�)�/���U��h���KC�X�bO���e���	Jn�8�1K�i��pa���R�� �%��:`tbqR;�}��]��?�#��e\�mǨ�M�3:���ʵg!��M���C�X�.��2V���"%��/�ֹ	ᣮ�0�����k�u�'A�Ѹ�*|z�u�����fiVDpv���
�!�����rͨ~*^���t����N�B��I(8�?�od�mX*����j�XlxVHYEB     400     1104�_�UB찢wL���	�Nq'fZ(d��߾�m�wFn8#�[,;�|��+��=��G�s����Ts�]��5t�9}JR��+Q׭��LW;IM���(���� t@NR��[�������V!O�BL���'����6�+]�b���2>ɦs�K�P���FO��G��\�4m;?J�N�Sʢ��Q,ڀ��>�J��5�z�Ƥnqe��^�<4�����i�6��o]�"�QyA8O�y /�s�Մ��5�ԭ������"u�,��z��kXlxVHYEB     400     120p|YqӴt dv98 uG�{@�í��Y��,��2�]��,w�J͖	��0#b��<V����1��o��CPp5r[��&��Ə-4-U�c�Ơx�����|�:�޹[.�d�_ο�|��Al���s���WXX���o������_*������kz���b� ���FU|t�c�4�tj�VnK�_F�FJ����,bG�R?-֥��/�̕l����g�v�����?��fᜒ��޷��;g N5ףui�<[V��H�F�WO�΄h�*��٣W���XlxVHYEB     400     140�h��őu�*���`��7��:m��-��=�1��s_�^9�I�(t`��5�����L�]���0?;Pf�7���slfTs�i�.���9�9a�5c��a��>�)��yw��-ڛjHi�KM�\{()�53�����Wd$s�'6?�~t��Sy�|���Ӵ��
mn�8%���T�o�g)��	HoI�{�����-��
0��K�-��)Nv%\���c����r�'����h-��}v����To�3�<0�x6��4��`x!c�.��d������{.J[բl#�4ن���� xIB@��\�y|�i:XlxVHYEB     400     140�b�k��V����ž���v�X��C�w}��`��{�Z�A�!�Ĵ�X]�>�T�e��h�J��=��@��v���87�g�@�x�G�Z{�<��Ln>����Zb3��*$�}"ݎC��%;��:�*���Ӧ�By�c��-�uXC�f+��sҙ5Ok+��r̐U�Ȋ�]��k����
��_�����#�l��itX,����K,�wv��4��ApFo �T�=�B�
yU�0��K,C}buAy�tf *=�9R�h2y��g�1�X����Gغ�j>>�Y3��YV����O( �&U���:�Q�ԝ��>��x��%OXlxVHYEB     400      e0�AD��V��tJ(\��������d>4V��L�&��K��õk5�f#&t���Yi�:�u�e!ix.���%�|&�fɺ����r<�Y���dO�������No����Ŕz~���~��i�L����u��ءOO��W�H#Ԩ����F�C\e#W���>�W���o�}��hn���7,~��)3}�����̧��5y/�$��r���oV�S�[�1yXlxVHYEB     400     140/��=��n�) ����M����/�b)��H��lxV"��o�LIe��)�QV=Tظ'I(�e=��H�m?e��JaHW�&�i�Y >��خ��Y�0�L҂�IHڔ�H ��^�#T����v��J���a��K�<E-����)�/�p�rfɣ��אvg�D�Q:�[��ozࣩ��b#�-|���O���4����7��l7�ܾM�Ƿ"�V��?y������3��0����ߖ�S �Θ_��A���p�k.EPs�Ⱦ\����X���1G�6N]���2��?��(Ð��Ǵ^�y��`V�uĆ^�!m.xXlxVHYEB     400      e0��I�vv̌��.!y�1*N=ޚ}�Kg9�Ir�+�B5u@N���
Q��aX;~r!���]�-[��eg�2�p֌!�Ї��Ag���n��u$} 'V�`�e������}�L����ϧ)TX��/U�VW��T�l��0[E��L�R\T�R�V�e��T.�^[��?���oQ�(;A�DA��z�HE�3��C^*�G�N���.!���2k�������T�"�XlxVHYEB     400     190�e0'B�t�׶*�Yu,�e��b��Pa��@�R>ӂL�ٺ?��E?�gX$��sձ�^P}˓��T%1�m�������g��*05��P5����Fɋ�"���ޟY�l�9���3��<�
��'>�9D�M���-˅U���HN���l�9�$Ëa�.XFG�>Z���k�{<�>�PG��,�7yP�f��A�a�Y�at+�dd�$0�0T.V��y�<[� �O��`�	MM�4��$�B����M�3�̥#�zu�l,7�m�0w���mhWO�J�����L.�ӓLc8�^�h�$)C���^�n�����T%��� �;5	Ke7��̇l;���!d�:���%��H��g�T�!��ӑ�y�Ii���O��cG� �1�SwXlxVHYEB     400      f0�f�M'A�� ����S���xi�D�YC�9��3<�B>O���ǽi�h��Xom%��I߾��*¢ÔN���2� ÀcO�StA$f�=hOyٙ	{����>�g(v>��:6ȩN�ђ�T?�֭��u9p�����͒fN\Ius)V���P�}�X�F���#)2 E�:,�9��'�Ņ�����
2I�WE�~_泇�p�#�mi߬�0LU~���C�@A���5y��3�m�=,���m#XlxVHYEB     400     120Z}�DU�ܙ�6���nD�P7f��-Ჾ0r�T��rR�'B�.�،iy�n�̓��H����j�9r��K��5�L?�%qD`�|�~�z�97���Z(C8g���sC;��g��+=�zp5)�_Q���_�ԟʥ����m�^-����q��@E�q�1_�'j02�f��a�u|^!�Z�� ��V�S��H@���-wM�o+�{�'���p�`!J�u���Zx���K�(�sx��F'FW���\�\o]xܒ��GPA�O�51d9ig�XlxVHYEB     400      d0i��.�8Ӫ��$�j��-�P��S��J�	�@`��Y�����^����䵑�ۑ�]s��t���4�̛:��q�Y2
LH76�<W�@|T�o�,���]�l��Ms��"�e`���}�=��� ��΁�6	�5�l�$�7b��JK�V��������c7Zñ<*��=K*��P���-'����ȑ���M�_bp�y�0��������XlxVHYEB     400     150����bR��id˃x�Cn�;������H� ��w'�ԯ�Za e`r?�^_"���5�Cc�1�d)���m/�眧z�x6N��r֘��d�l�b3Bݖz�pg���^��D�KT`�]�D�u�����7����O���@4�붨�|3���ګH�q���n��q�I���x�q����"�V��� ����E��"�Ӊf�gqT�{#���v�/Y���:E2`)ʈ	���c F61'����$\��S��2�t6����x��A�*��tZ�L��3���:�B�<�2O���K��Vl��"����Sa�y��ޖ��%K��Q�]�iQނ�6�hV]�XlxVHYEB     400     180�z�JeЈ@�m�_O��`����#�_x`q�'�a���iaj���~�N�"�E�t ;�=��w���ԥ"e��G@�p�	/.#6#��mWTX�<b_�� z[N��Q?8l�J����d{���,c��+�J��Bm��g-9�"�E�U�k�Y�n�w�h������@	�)��k�X����$a=-.J��/�Z���O���� 100��l,�U��LX�0��tu�3��!l��"ڲP �u�m�
l���>�O���/�:G�QH�>�P"�9)5�I+�nsZ+�����Q\Ϳ�JP\ ^�6ig+K��ė+�\Լ �ﭻԗ�+^G��z�R����^��Zg�:v2&�l��d�f����F�k�XlxVHYEB     400     120W��4�iMT�e�q�Z�| 6��(����e�	���֡� 6�$/�插,U��g��po��f�݆��������E��	sr B)2�2�*�~n�2<��%���!լ���ǎzؕ�V���n$�->��W�j�L�� YY(0ꂓ�_)Z����R�v,��0�!͈۝�U���.F��gd|�9��c��}���l�"����q�w�hA�;��#7Q��Q�x�D��c ��4��[���)H�Oy8�vg���٤����5x�XlxVHYEB     400     180�n�Cw3��b�_i���_Է�`�D���˵A�T��#�SN�Xt��Dt����?��!�&�X���BEZZ����~	�O�y"ށWt���_��l�)\������<b�ֶE��鱞-g�1�^�j�0����"p�G���W��5-��y�fZ��L,O�<p�`�X&�}z��d�q�	к�R���V��U���ۚ�{�04�&ff�-|��8���&T���s{H_������6\F��~!�
,�Oq`�|"��T��]�)3	���,��[�/ӡh��c��ψ�����B���H\�Ʊ�t`ߕ�js��ٖ��UB~���pՏ�E%���n�(N�˻�OU8�py��%��Rz�)���i��yYXlxVHYEB     400     120|��ҵ[e�}k(�	4��"�������B��Kԙ �p���?sW��v�i������9����9�|�7��5�v�>Q6�ٜ�o��zs�!�EP �t>&N�@K��P�l� >��8�$�4]�ŪWBZ�|D�����j���d:��*J�M�i�	�R2>�kCb��n_ZG�p�@A����0W�3>yqh��Y�Js�f-�Yҿp"�L��~�@Jc����/m��#y@{��Y��Vn/A#\���A'ȆH2�9.t6��7h]3Z/�,奜*ʥ�$�XlxVHYEB     400      f0���� r]��������aN��"EO�HW.���<�+�d@��B�z��Z�c�_.���4 �����e���,�5�{��G$+�S����we��(
w���'�^�A���P�=)_�p�`�yB*$Pddi�����c�5�3o��K���Z6�^��t'�{Z	�����7{�C0�����<�(�pH3��P*��6��pN�4u�P��&$���O��o랡of�C֕�t�ݫ`׼�|�XlxVHYEB     400     130���}	kQA��v��nO�V�3*<ֳ�6D5�a�b�ߛ�"L��l�;*�1}�O�$�̧Q�Ӟ=o�ϕ��뭽7�տht"�MK���֣=�	h���������nm���V���U��{ˆ^~��n�g@���a4ȍ�W!��X7�f3-��?�v���/�|-�士k�J����o�?f���T�g����^ ��F^W�v����h������KA>H�����|�Yd�����ג��X$"6�*Q멮l�?�O�^�uJA�x3,�K����c�\�_�o��]���`���)D� 1S��XlxVHYEB     400     140���Ɏ��H��S_vj�t��g�N���m���e�X^�{o^{�Y��)p�Ňi�&�r�����&�D�b�OL��L�X���� ��N
��6��aVe����y��U'���qmaۦ�
y�F)��l��.�d�}��j~#L���1�� ��ш>q�|���X�J�F�dr��C�;�2�{s�L��3��ܬ!ʺ��(�����|_a\br����	����|E��?��f$�~� {���ؿ��uK�vqV��`�-�T����5��Q5��[����Rkp��'�[�*j	�������3Uq2>�sk=8XlxVHYEB     400     140��aw���c.]�D�<|]F���b3�{���Y�����xp���\�J����,w�IӃz�-�l�G��B�e>#4�����z�:Ѓ�A�8�}���f.RmAc��7A�A��NI۲�۳��-!IV黨��%��|������!�aQ>r�i���zhYW������6�Y�����)r�8*qN�
���Nը��ػ��_A��,"�l�E~˸@D��a�ͷ[rrI�Z�s�q:u�K��	�v_=x���7������x�ES20j$�& k�:w��r<�&M��-b~)��JdnO_;�!.��sf�XlxVHYEB     400      f0�ݛ7�@B}S|4�l>ƕ���/��2�X(k��D�G��yn���CMcL�ß���3��q,H�K��d�e��?�Bü��Ӂ�Q_��V�����.ϯ��&E�����{eQJC���F�8�-�NRO7�
�9�R��4�yKL �0b���b,cUu-��s�n$&r���/cd�"S�6��&Y�wH,��Z9����:���T+v�W����i��&\Bɹt.���pS֝⣚_dXlxVHYEB     400     140�J%�4�!3 O��*@�'��F�Qp�G8�����������i�9Oo�U�~�g��ѹH��sg���yz�������[)4ti�^�{,��������aS��Ѿ`��?��hX~	4Ⱥ'���#�ӫ������8��^Y�M���g&�,zچ���g�D���$�-q�����{òr1Ӓo��ل�M���3�wgXF�q݌r&������K*R�|�6��g�$���6�	���!���Ĵ��E�okF�x���3n4ے���u��Z����I#7�!��~��X�	�������uKL�}���Ad�b�?vq�XlxVHYEB     400     120A�q��"�WHY�ѓ�-��������30I��s�ax�Cl�o��7Y�8�3���}�F���;��d}������D�b�fW����Z��2 T57x��y�6�����p��X~N-�ￗ�ե;�Ř����|k����^"c������B�v���a&%ݕ�3��E�E�H���:˹��
Pj ��m?�RO9�D�GMm�I�Χ�溾��Y�W���݉u� #	XmdAGa���}��nZ9]�?�m��H�!� QYL��3p3�\S����ҹ3� a�sZ��OXlxVHYEB     400     120}|�ɘ��#D��tϷ����i�̬E��,��x�?�x�Z��>lC�Á��[k8HI�X���V�l�G�~��gQ�}�WM��U����r@8��.t�����I_�8��us�T�Z�D�U��~׫�;xy���P�\P<m^��K;7A�� }�VaSn�_�k���BD����lc ^�SL���{�p(�1�oO��@# lo��$%]0-�nl��]mf��w
[@B����q	�l�t˵(Q�L��LV�pL�눦OfU㒻Ek.��I遫ǫW�s3XlxVHYEB     400     1109!���]�&�k��%�^�g[??�s��J�*�	��(�p�`e�(�P�	�����muy<�1���ٕO��\YJ��455\CɭnPtZo�E�q�bft!C��*�����§	|X�I��ꦪ�W��r�~��M2�q�.mf�/m����}�r3�B&?�����ҙb/�e�8��I�I�'#yƖ��^~�q����2=J����
���4��)�9��w4���vhAݹ����4��W �|������g,���`j�Fg��E��jXlxVHYEB     400     160�5���ۏ���/@Z�a�ȴ�(��^;���P�5�4�Qj���N~�j��I�eX�?Q����fG����
RN������O�DszES�]��'��Hָ:�b%�����ۈ������Q:��ᵿ�#|�r�Yhٲ���w�i�43[
���%�S�!��I�K@��ݸ ,��O�|�O�u]��ꐚ���H]���:����v�֔�,>�5�Ouk���\���l��R� w���f���P�!5��iQ]m8��cv�Ȋ�:���]��Ɔ.��p0�jK8�����u{ڗ{ ��C=�m��� �	BFV���N?M�
kK�c���0���t�f�)	/vQ��%��eXlxVHYEB     400     130;�$�T_� c@$����̤Ѫ��F�������R$���>1L�����ͪ�f`�&ƫ&Ֆ��΄z�b�J��#S�
5����j�l?mS�;��E��҃��.����a(B~\��� z|U���NGc �Qm��D�M�-�%e�8�ѽ�L��b�7�C�X�[I$*�W��շ��S�k�"��L7bY�R���ǀ БbY�H����^�[���{�ND1�N{U\���XC^��m�aH'�.\����\�� �H����*��K��[ˬ!������me$���8/vXlxVHYEB     400      c0ۅ �ĂMx�V~��m���@!���tp�u�/$�RU�����G�r>V�
xF�2Q�{��M��1�k����Ε���b@�	����<�?*z$l�!J�=�MF�p�!�E�77]�A��5��0��ٖ\����^�`�y�G}�<-�t�^�'�gS|o�&?P��|Z���ß]�5~5�j.m쉙��<XlxVHYEB     400     140x'�G"7PޞR-��xڞ�o��=[��=��{:�-�Wu�l����-ӠK�)�<���Oi.����p:��X�	й8�h���%��<K;�H~ }�et ��򲼩ɪ**�3B�5�������A��D��6�77����]�$�W��ɧ�B�#  ��sӯ�V�_�yշz��=�+�W�ɝ\�%O�_Xy��Bc>Q��
�_���A�e�!�@~�XK�KQ U16�uP�M���7~������$�~Xȭ���V���@�Y`�OV/;���z3�d0;io[�Bz>N�Ðy�ĉ�݆>�ޑtg�Q�/NB�!0XlxVHYEB     338     100�r
�u]����b���(�����=�2ͤ��3��� �8����Bcq�5������ݤ���^�7���=Yо�۷Ϭix�_�-�f���M�A;��e(Y��[Օ͛�ܲ+�*0토8r��w�	��vO2Ľ�)�����.�x1��,T�:K�I���B�4�c�o�il��g�g�Ob}~P�x�\�1[g��c%%o�����R�u�?P��ҨX.cW��6 8�a�P����������H&�� 