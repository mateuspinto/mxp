XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��y��?��]��#��BN��Ngl�9���t�JՉ|�}5߿�
c�yN�8�v_��l��\�L�C�g�}��&�f���~h�!��֏�gfN;ݨ�Zx��	@2�ZH�dLϷE�"xK��yB��wܼ?�Y;\�Og)�X_d�h�4S���e��ާk�l3���s� �������QP	�e#����=�'�"������J��ƣ!#��ll#:��w�/ߴaYU�	�,tk���&�vKSQ^�E�� S?|u�x�?2���)L� �V�>A��`��;��կ�EA(�,�f��3u�<���F
�--��8Z�p°8Y\
�@o]PQ �|@���QTȐ<�/r��{`T�:n$�c�k���>�;v�@�������k�̀,����@�U��u>�٭�i�cJ���^z��iUc����>�������2g?zNc���	����-/����>��9?���c�����nM$H���2���&�/ ��!L�X��'�����`����}��V{�Vf~Ԛ~��y������G�&��T�)��@S'u�?=�>���0B,}��i�G�ћ龰�|/}ϸ����N���!!������Ux�J�3���g�Ҍ�cT�V}Q��]Vr���.����'�ߋ�����R"�� �%a�D3���4�`�ï#(��讼����59cx�� �]���"�Yϻ��y��f"?DH8 �`�%��~�!�����T�L��i���u�Ѽo/��fXlxVHYEB     400     190���\�.�J�gy����u��]4C����.hjWR��FAI�g����9!�5���Q��x#	���'�%�KDX�BX��8�T�F,�jḊ���q�����Dg���1�n�a$gt)3���jI������������v���
y�Hf̈�7�7%�"qʛʼQ؊�c���ؓ�`���E�v��#�.G>ޒ���t)'�$a5���Xz�������A�'���w�”�h�b� ��,�o1��|
J*}?�xTmss�,�}���7Ԡ�ŝ��Z�f����M����[��Ǔ��x�T�-�_7J�P#SM�TY�(�ʅ
��d�1�jlr}j��
$��Q�=벏@��so�{�Rb~Ee?��)��*�B�����e�%�Sp7��՗�!N_5~�B�+XlxVHYEB     400     150�������7KJ�����G��L+�J���~��4d����Нo��RǖDB�'J��iI8i��D
�v2$���W&�c<cS�j�=��^~υ�Ƕ�Ӛ���cr���tH����HW6�bE�
�Qߩ�p+hH��
�n�7�2bB͸�4�������zMͲ��Xگ���u��:,-4�����N�#=_���Ƕ�1c4�uZ�c*��3J|�a��,=W��nE�F�J ���-��
�ݍh!���>�S\B�b�:��0�u�-.qe�����\va�n��Do���HuT������:L�B���Yl�z�b�XlxVHYEB     400     140��֯8JKX����	�N#D��g�ݷ�ۓy�z�&\��x�ݡ� �D�3��o�5��W� ���CV�����V��k���Hc^�A���F.2O'0(OHS�n����ꛑ�m�[����������)�4ܵ4&�:m`1&���������Ya��Sr![�(�P&e$��2xH��Q!.h�ңZ1
��]Z�����JB�c��|����4=��99���`y�� ��E;#KˮL�/�oJ��|� רA��P2�T;�4��z������ST�Ōڬ�HW�8<E�X (���	S��1Rb(:r/�[��o�XlxVHYEB     400     180��
�u\�H�������zM@<���s�gxEP�
.' 7j� j��1L"�M�g��-�����,�~]v�a���TN#��;�<Q�t�����R�j"1�Z��3 ������ͨz'�֍:O�ф�4E:Q�����wC�[�6s��J���"�i���i �#������R֤�f�b��4B�o�^��y7".I��?��W�6[e�y�b�3z'ﶛR�Eur�!_��ҋ�~���*��D�e�#�/G�} ��;��d��Lu_��n���B��qMȝI��'�Y�%�\�$CQf�[�q��gnUd�}�ը�u�� f����G��8���1.��2�F(�M;�������� �����Ĕ��8dm̽�Y�+��u�)`XlxVHYEB     400      f0(�S�c"ϷGk���t`_�Ѹ�F��t1�h' 8�W$��|�zSyF�<��}.xe- 	�ϗ��Mg`H��K��<����w|�d{z�J*l�Pl=s*��:��;]
Y
hL
���2��}�֢	��<G{U��I��C1�V�>�P��:6���^�f�şR�>�@�V��,t�c��)N�9�<(z��/�΀�PU�ݯ��ĕՄ��ebg�wv���(�R����Q��.��XlxVHYEB     400     150�Srcl#m���_g��L�-}��?����D-5l��W�"�m_�-N5��ic�z���F��fN����.L���>]r�W���tI�9��s���#�Y�.p%�ޝ	X�Z|�'v�h}�7"�c��$ѵ;���$n�G������+����q����Dg����+�ΒP7�[Ɍ!��0�kK�Lb���ØZ{X�1$蒱a�$�`�����̰½��i�N��:8��"�n�7����i��0'��zؓ�ɿ֊z��@5�\HXC���-VT1nڭY]��-j]>���u���\����埁D�s����&0���N�]�XlxVHYEB     400     150�v
j��,�A>���w��U6sA񵢸�ߞWLΙSG&��t]�_9�g��S\M��	B����n��_*�$]�g�?x��	w�i�HRup�I{�8V�RX��d�B��9b���*��P�/J�\��p����<�щ�,N+�n�u�!!�㉆�*GqJL]�Â�N6[k�r����+B�ӱJ�����PC������XPV�Y)j��^�{x��{�n����d���Z7;O���57�����iRv�R0�Ao�Q�^��������ɶ=8&��Y��{ް/���8�Q�B�h�F�t~[�<���$�ջF���)Ӝ�}"�c�Hu�Y�L�1p=��
'}XlxVHYEB     400      e0�|b���zp��ǉ�dz,��xr��G�E�HO�zxP9�q�|Y�vs	n��	�#�]h���kZR��� ��vƁ�e4� ����p�q����+�.L���G�"�&���"��t��PCȻyr%H8_����.�EBn۞h�� ��VI\�o�c�4��<�0�X�q��l���&��3:������\R�h��/򼱒� �R���� ��XlxVHYEB     400     180=�v�C�u(,Q	��d�S�N9�:�KL�C��p`y0�l������o�j1vN�4��͢�i��EO� |��f�<�2�2~�5u�!��$�B3{�D ��+��
�����v��B𻝀�R)�`���َ�Wg�ưԁ'4��sLy*Xc�����H��a�iKB?����=��7�~nlJ���D��>��:Z�u���2c��(�^��#���[�yz}}7^��ߠ�j�����!��l� �:{|���p�P��z%P�q�{F�&���:���M�	���;;�zpת����������v��ָֳ%���m/��������	h�7���,�D}��� f?*�����֚��JLd쭫�-���GXlxVHYEB     2f4     100eAZd���xS��I?�$Z��C��UE�?��h���PZn�|�������9x�R���u� x�T���y��o�(�)�7gu����b-w��J�P�"b�ޯ���8;����'��@�^�|�w�f�W�%�uM�ů>���D������r�iB_��`��� ����>Y��J�e.S2W(Z�	��kz� >�TZOx���\i8R^�N���S�|�l!Tw|Cx���4�]��Jea��,�kG�����v�|��W�