XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���� �O	�CM��������\F�k��J�p3[,�sL�T�i}!����۷�;��7�G��>���ϲ���^��bmlb*��j C슥K3�t[/퉶3>�q�/��3(��ș��W��0bF�K�dа�g	
�O�C6*@��ⶶ��XI��ᆆ�<X�db#���c2G\.�}��J9�����$
0	�ҥ�����@��aV�+�	�L�a�p{hcF�m���RR~�Ǫ�n1:qoL�ِ�a[��	:��{-oO�ڤ̧a�#�W�=�i������!��"��MZ�i��t)�:�t.�y�\�2H�b�����������_bu��#�Nە8ך�|�}���֒u��Hc�lӞiZ&V�ۯ�����:M��N�A�a��]�����8; �q���4��&��K;�
��VNJ �:��C
�H��E��_MvBt�{P��m�RG�e��Hp�"��BhMI�q��CͿI
����0U�j ͯ.#vC	�WZ�i��L�y!����_C���N9⁡.�8�혝]���֦�*��Tl����j>d����.��V!�!�!�J]A��DE��y���ڱ)��`8�-x��r�-+���!���K������ϰtH4:��ԷW�;�ik�t}r�O�{l�&�Yi6�ߕ!�] S�����+�q�d�\�選��	:6sN��(��Թ��	d��X�]�����Q�L|ќ�:+�`�x ���EXlxVHYEB     400     180f [[5��R0X7Z���-���L;�z�[	LQ�d�>L}yZ��ƒ�1�W��y�6qCH��v%�%�xR�W��w�H�5��E����K�����|:VP�C�^�׭ &�Mk��M�(!�C�[��b���Q-A�,���k1JS��5�+mO�$�����`:�('|r�ZI���*kN�)B��9�B]�P�m���Xpئdi\�Ř�Z��!���n;UV�=u٥�Y�f>Z/ys�D�lU�������}C�2�h���� F��؅\�y��@�T0���>��ل'�&�ZB��:���s���)xU
�&.���׫QE�h���k���C���x��' ���K�*9�Cv����^Ab�qe8�J�XXlxVHYEB     400     180�C4n���i2� ܀&\
��������uG7lw)~���2!e<Դ���T����\��]j~�-{�n,9CQ��D"-��)+md,��T�:uNɧ�#�nl.|-A��ZhFҩn~�=C��zߋg�x=�H�q���:�����`�P��m�2�l)�lj>�����7����53��o],.�t]���(��9�-V?�����,��܍�x;�"�[�2��唢���o��ֽ�D*gNp!{EȖJgzqj`&F�S���GPT�}>h�a��w/|�t�����K\r�m�55Ž��:61i$@b�!16�d�$���YˏO�F/_ltr��y�]o\Pn�]6��˘��-���ԉ�?��]���N�n��t�'��gXlxVHYEB     400     170s�l\�?iA7I2I��SH��YTG�S�f�_���׀�rpW'���ʩ�K\_Q�bj�"�7.4آ���5�D9�|�X�����92�����6�ΰ� ��T>��g��a�����o��NHnSP2�ɧ��dΏ+D����)����h�㢼������z���t�|��{��XyT{��s�f�;Ȇ�O��bJw�{��ՁR}$�������,�\4��I�=��t�3�}��þn`�V/�0B��+��L���f��L��z=�yکEז��d[�e#$	b\��p�*����*@�@P�j�����l�h�� <9D1%����PF��Р��
FȐT�W���dx-�|E$�.��XlxVHYEB     2e8     120��rv"����#�=�ۤk��/�}�xy�`�@�=~曼����m�$���F,�B_���{^�<2���!����:���^���m��	ue�3u��>��4�������~h�OƾF�u�L�0��a
7N�K�p� ������ن�7������1���YR�����ƒyCqjTX��;v2�K}��#�j���� :Y.z]���k��d�f�I�\HxK�iH�H:;ͻx��"2�Je�3��݋�L��"L��/������"��ӷ��ހ$�