`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
tB6Y8Ow7j6SxJehPu3U7ZZgxxsNs2df20g4VJq92r4eh7kTR5BzDWwz6mSwmQF0lj6MBy/xxtxBd
SKexyUH1Ac9CC3qqfJvzXX7+zhbdFac8yq+PftH068/bMGAng+Z8EwHga73QWdzy6FBY6dVA6+rU
CwAqjUCMPEcf0oIr+fZpk1/j6O2xFRhlTBM6yvojeHjIEiPrJQLgR5C2Jd4V21qRninb94TW1CEP
IAy4VUcCDYfj3a8VDElrt9MSeEXh3MI6zp5sGEEhL9CZDuKDxq6QhVzGB3BQRvJEAvtooE1fnurf
jTKh6/j3fyt3sIfSYygg4loiCvD5Mf79KTefMg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="Z9gx6ohUifjaLaSO7PyHHqFo3l+n9AQCvPytmZezK6U="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2368)
`protect data_block
fDqSBvlL4B/gr/1ddRIsxXDMytOfFQQGDmrDjJGhjS6hcq0kSKXDm7wDxaw8qM+0jT1vzzffuVsB
Cg0ShHBtC031rGmNNibgAAzkEmMNhru1d33ulEuXogdtcU5G95Z06XpixnoDIA0Do7ezg6afD+Gc
eMOttgn3Oe0mYsgMyqOjwS7D8UHAsnOrpO46Zeo6aYo4Nd3Zurow87gGBBYPf7nrbrzyXhtgX6Kp
LJxbDD7HCQbeV2qp6ngQHIKE0p5K+kOQcYw/vuzPNQ7/JMPswoeSsRoF5QwzxciBu1zP+YgCOVjh
bqjtY+2ndiR6EluN9swQfaUAnjyapo1AoarFnuyXZX8xGWNDXkdXVK2qCZk8oDxwGOIEhFeF+HWF
ZzAmytDedAkWttRjehNrCTLDaqE9pPU78BXkkWkOVWadtOkpWc8V1QDnea1oluPy2++0kYRcytsl
RWkUDAtAfe0GxCrUyKTLLA+5vAkd1sAQ8+I8xgeeBz6vt6jaxrxhBwSYa4kU1ulp9acE+Hsnb5he
DdQCWmg4TV9VjWorVg7951lvSks5lXaspfah9L0GNL91ijbajg0GR0rOhQNz9PrON5CtlPA1fheB
jMKALbHLxePVOFe/8FTx7A7+6ezloOGxLVTvEEn5N3THD9opqjM/NuI2t4BYji77uoopLCOwMDtr
B4aZcRLqwRY19KhDavmm/Smk4N/ZnFdmfreXSSaFUaH192ojXhLOClvLb+t7icYWDX14C73R+wJn
mTMOejg8T1NIrcPuoERBsrXvjwPlGSC4BGAJ1XyMsWtPAHxY/wfckG6JEpeqSFJie1cu5kTlCecN
uDywcvaK0RVG0O2Kpq60yApF/WkkFo69adPBmxz3ALleV7mcpl/ucB59i6LSaE6WkluxAPqzojM8
0iUAz+VazPJKeRguw009D9A6EtQxNTDdK4+n0Lb6nTrQViCYr55m7V5e27fdNSOuia/6fG3cboZZ
0gIYn1iZY0nLvpcDsiPwtGhzYedKZIowapBf3P3lEX4Y4Gq+vhZgcn3CgsPEixwS0eagUgfo/kL/
xyPbK6RlmpQDIZqN7HeVlnlEIVbfPHPzo2WADrV9HxqoZgc/I8mUf/T/FF1tPxdo+J26lK8UwbgS
oSjcH1ZhjOEEebT0uyLPjXmVy/axNN3fmn/5gAlzOBNdQiPHjpNk3L6Tshea9u01kqWq5Kchfcib
/6M9rrMINCwER8pbm90eMQzS6gh+jXxdGLMcs7/vNm9TV3ktnrNNOF1i7pcm5fM8KK6yx9Qe7Cne
7hD/55oi27dJMs9ZekJRtvVXAbQdID2VTlw0WY5ImbQxhHfq3Jlb79CtmuV2yIquRKbn8m0oaLhp
5RnIPF2Azglt3+4RRz8Cp8RJFOlGfOfM/K2Di5IjVJeGS6OFM5kURsuIeym3G5s9bSWK1glNbnbJ
JccK5nmmc/RmQw9G5PEq1BjPhYhwTcQhrIIudVfZzUYomBYaQVOIN+WDO8D2w6/aemaJn8u2lzK1
9XdXIq9akiFMF3dozuSwcrOmz3JRKB+XbJwjxm3Wz/DyZInQ91NUPouuMq6tID5bhX+GXWvVi1GG
jI1JYPRPRtgl2JHDs9GD9DGm9CMFK7uonDggnZpL8bG2nRht0HJ7ynZ9gqU5/bE4I38zOQlft88t
eB+sWQR105KhLf1yOfm2al/wUZzBMfDD8A5YqiAYDScUN95PUUvmUGN/qLEt5nGiM9hudmbwHoEd
bked5Mcwu2l4L2htUR6VaCnqPyh8ij1E5T1MV7WhcVys74PZh+df5l0nH/mPmmkrqq5q2Ziy7LxJ
LUCTuJtezxKOFsCw0xBoDlEBlT2h+B1/QoBDR4THJsw2u4xceJDy0GuLrVPZ8Ei8aQGEPw0Szce3
/ltXi0A1Sl9KXQHzjzhmA1qhXi2TzaYFANTborAe5kcUxkbAmL9IHoC97d7DXTdyd5w7uqZVDvoT
YA/qP/fRTXXTihiyxNWCESZh0q57ueBn9JqvHsENJr1J/6SQ28plGCCw1U2WBJY/FLLL4Wy+80KT
9X5/jM1zy5n1EnLSmyf6N6MCRHcPILiW1IqQ9Tb7dFh1CK7vjoFrzwZtUNmjnL2Ps2HJuPVwpdhf
uyx21HeQ4tXSMuHdEhvAdjCYjkl8cAPRqBQDqjCzeJjRLtwIWzuAUP+4OwO+z30qoxVL9SuN00OO
0v+R/orkvO2lMVHdaQQZn1/A6bT4Z6cjdNlLZ30W/rgRfw/N5Vdp1Lpg9Yn/JN6LJBxh9wqy3LeI
CiuyEFb3N+1B5OxCtSgq7xOiXNMYLceVTHin578xDakfSfUsz338EGH3fDUZI788R3NaAOsjHjeH
NDkhtQMWTWYMAa8KMt28YWKLk3J6VS/TmrupTjn9wYI/F+bNP8jAwpQ6JuvAAEAuXayyl+qC8eP8
+MGhTJi+IUDwUxOIcFCEJd3cWG1aKNSomOo/+2GyHCx6ZAE8OQR0ifxep/r4C5TUF8vmVVsHX9t4
+DGUxXzdedc4/XHzddkapgMqtMPfyLJuCj+lq5uIKVz3Zi+cNEeuHQAuVLO576JWtt/LiepesBxZ
ZcY0M/oZvA3IPyp8/MIuQNOUGe+Dir5aefUiHQANhwj6fJzrsDgBiUjrzITePZu9rfGFaQ0elBj0
Wn94iquYawY8pNRH8YMDFFIe9MaF5v0oPJULjvEfHhsccwl2vixmPcstaSuBqJ7twLOHHerieXrW
yxFCM6EGBKciX0Vrn6dY1DD/oVKSpX0zaQrtkYakIgJlHpD6L8mKKrUhzW/r9X257KjBSyarlKD/
CxUMV6anJM0Z6hIj8AXoK6Bp7+73PdYD4PuPNwOaour39Ds1ycm0ScGwCUOYYiotO7pWTJSPpsz8
vSF+FMSjXxTTgjwf4KRXCVC0UvnL7T2dLY/CyeYVSTT3W/9VtaVECCPpiCH80618hb7EvruNFCpA
3rpx4ppDiXDFsd5iIwdmn+YkJ0pDi1VDcRAJ7VTq0fryYYRUZy7bEoDQ7EW+gcsmwqPhyErGjVDk
Pax4YjSEOHd4pfQrk+lJBoS8BtAOPRwFY2c7EWf1I2SNjG8/98afkOM04v1qG9TM8eo8VNNkkH2v
kgjyWwFdlrCLjmAzHw1PSQofC9xRxiH4JJYG7kPSEg==
`protect end_protected
