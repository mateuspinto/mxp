`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
W2Cj1i0tF63ghwRGVuVyvkAM++EeobQDVpwfGOb/V3mkHVSWytrgj5qttgUjsDqDx3uSeVzkEBnr
frRzYlaY7L7dMjB0oxaIt22/XelP4pQURlQmdjle32Fg3u03ph7rptnW64kFHTM/KPk0lMSyli0F
wUBfrhISfuzrhhZGl5o8NiTQwmCNZpPYdVKo6DSORxBGEM6ynAtOA2FTTFanVkTzoGIqKMH/Vq/f
PndF0/fcb3a5gK3SPBnLy0W0gRnAw/rxrJri+lbtE+sQiYwc14pqoLIQBCBfh/lLFZN3yoHwS97S
w5P/EUPiSXb2ymTELast+oZIKCEX7jrpRO706g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="NokSfV06WvgEL/PwNsuBIISnpz8gnX8UPMOlf1Wl+q4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3056)
`protect data_block
a7bDFUzM6YFY4DsBwVr83nzUxiEFBYz4U9F+tFjQhQJa9tzjkv/gA3g1xbrg9nX23VVlGwCsUieh
G+BbbhWkQ8GoaboXDcz3IXP8XxmUljXtO1Rq4yopGSBpNPsGQT3+P+yPs4uZBXPLq5T2gcJ2r+1M
fF6z69iCwQRYRjq6L7RPcK7bhPArhJPPBS5/uzIWOtBnacuEseewNp1orZS0rlSeFvdbPGEXHuHn
xnApOhJda1JrrlsqVrG3JZyRUqh6Fi7p/EWVtQhhYh5h5uZA6aW0cQgYqf4RW+fV0E5Hwsym0ZgG
wh33CN2gMs0tNEcTuPPL+oJF9pKk3UZZz87gq8zlXtE1d3SJFBXUG+rYVYWFtzv57Dsvay+avuDF
GUAiTzbOQDy87NmI0YmAN04/Jf2OoTs3iPSa2jaVdcdFsD7n+k+uV8fgEdV3+KDVJ9wJA70J7ONF
0KmUK1xFDiQ9fQkCdaaVkqwaJ+JINXq0zfe2qdQNWxhnsJBFhS4xhaS7xlc9Yo+H3sGIEjS2vQ6J
pgXmeC1wzZ4St7iSpcpZOEZmfdrTzzJMaM01EGJPEjly7Bx8Q7jNGCLjfwy3KT5dNToZvDDRkgqD
/wI6McuT11s3kDBa0v6Tul9Umm/w27VMtoyoWzSKFv3nRfKbMzJJK13MJaV4Io7dtzJr8xpE3x7v
TMbu8lqJliHepgfIO8DhAPHixIhkxQGmGLuIz39KxeS3VT8+bNeFg1RvOfHct4XlrOqxFEVH5C8q
/P3GDil2Ux7sdUuH8kcpX/I0q9aJCp0H9S75ZHnQVr8bASkg/lXon6d8a/7QI+ZpkGeYzlo2dKDW
QdVN2FCQTqFdLLj3HMWbAhn/xlOykccVyp7kE6tECH8asKUwPJu5FHMQPL926p4Eue+SCQbkWeHh
KaOFzQwdDB226o0BWL4vq97C6UVRxyGNIAWLzorf8/mC85nzpkUVZBch7xEg/q6W7WCtniImLgWX
5YVygV4TSDeX5DrZK8ZLGliurqsXU8xsoECmgb4V7F/aqy0VECV5Azxd2h2FegYqpNeTqiAjz58o
RR46a901kTfjtd5qBSw2M7KqpmGjfMG4GvQ6t24JsJqK+4GQy1di0cL5qaaP3f7qnQEQvem3Akft
ccxbLqOLdWJ2B1faoW46Cr8c7mPMzkR6mEG7Gt2Q+a0qTJdDhZ8zSTVZl/9fIgRBrtWdU0Qgf/AL
tIXO/R4cj2MO3EcTcJHjRH810jVlAIwJ7BgfOUMiqDruPczxVL4Aox7uajEZCJhYpR6KCvblOlSD
5rwuM6T+f33NUnh6EQgCbn5B6uMwWOUc7LG6g4R6PQykG79m7arlLkQpNBUUGD9uev0Q5+/H2VlG
zoXuq+DksD1xU83PbuBPIUkuS1uyyMLsAXQoGzFaP+JDSVEkvwtnxwQMfvbJ/qzqtPGEJ8GT1gys
I8EuXfEBpaSl/jQXDuYjN3XtkJH24xPx7yQt101KRHxWd5mQCcXB60ivD19JMtkku2a2JI/Td2lA
lLTcAxALnPeN5Culp1jccfxry1aEIeJTerb43ixE+HPjZEtbZFrm/fr/mqHKaBSoIuL+8vDHq8yC
ZTsO60xe3AsCJDPmhZG9jVyxqap9fzUo6rXWw6CVEny+DchO+F3Ejyn9GDmd1MTBu/f9Ig+z62j1
RUncuWc7n5yRFCm9UeY1ppQ6uJmaSoZ28hJR7iOdi2EhRHKFRVA2ppuA8lLA0Ba0yL8zSRwaMqvJ
1DLdlgXL0CU0OMLyVLs5SZa7VdTrktXVtYi5vOxIQ5o/up2kUCzawhdk/T66AsX9TTbW2OkTsMZ3
+VskcRer60+Kchm4HgRyqjj2PVSGa8hG+butzDVIzhShvFhjTZFMBXbm8UJ/3zg3Dd77GKDMaJWF
ycCl26nhTCG7rUZ5tuVPpPQ+VmoBn8ckPYIuy5GhqiNx6laLMFq2PbNiTbjFvT7o33QGMdFnvgy5
UvhEqPEsIxBKRuIfYit7qoClcnX10WpxX6sM2anf3oPd1+kUYvqpES59jgXGqjHX2V9FLkony2uw
f6Uy26NqX2TQotMAT+NoI/vtjP3V+76ABQ5E3QAHq92or5BDUXTKN+BWuzjbf9Vv0/fqcojBRibR
znu4SCI7gJWUJyJL9z/9J5Q8W56so52qxx01iU24Cxt1IagB9HsrwKey/eUNBp6mIjpm+3E3qvrs
lbAFCRxvQlahyaiF21gxtBCHaqh76lTIATMpbQNspQJCEGdaqmYP0jWMgxPEvg4n2NIKjxQ9rNsA
X+jV1ninjx2pAiZ381m4l+L8CkWJt8ieYwplQaLLLh2MD5QXtnOrH2sAWGDDrwdYv5C0COd2f38i
bmY6b9Ijft2jKXGISppGBJGvhe+Y8DWfD87M76mjg1AYzaEVfEXL6l0kbdLNCJZzFldEnPeYu5wT
p6NpoQcDjHKUxuhcfTMzhUHvUkZMgqegGj2FIeiL7u03AVoTL2jD9awMqw/zeEGU2cnwt8lC2wv4
J6JwduHZcRP8YCWn7bpGKIYOnQ4u7FLEzG+d4f7wYPPsHc0TTVt9RpAy7tpQcMQ3QUcRWb8TBbdp
d+EtZ7QCrTs8xq/UhdSLY6LS0xblkx93W9xLI4zK9H0xrhI7JEm78vnw3k+ycZNk6jrqJ4ZdV39W
36TDlt7q0YvAvyQG9dTc9Gg5FpsnjMerbFU/1l1re3D9Hrd3JX+CflRGGxGvPv4+7vN9Seo+WMcI
Y8O2Vbs3loN7ng5f9SO0Zo5ffB/d6WZFuWruJL/ATAWkLEYi7cc8gvrTlG2SVuxlewiqU54v+IxW
fR8+UDdTK7qtrfsOGiB6PguN60dxxFJSJDkYIroivhl2QFEhhH+VidudjeASci0x5LOuiwfHxNZn
bxlPRwBK61DyjkrSWKm2nbN79mNo94th87LYgOFcjJ4qo0JO2xmHNEK9/EfvKEjxriZBQlDkVr5T
aZe8D3gna+4YtkClGnpVTkbCW/DSAmqdQ+/v8EhphCHJDd5/NUQiO+5LvZuCnyWuHD83igYNMA7a
3g8HH2llU/aWb2/QQkpxhttMB00BjYpn/DE7AIecSD8gNnazsgnNQiDgGUz88BknYYdBTwnGr93B
M86qhwAq4U2oukD+rw8uo5znBFGZWXar6e3wgpKvTrnctlB0FDe8ulq39A9AqyrOK8cW1pxluGaT
CqRocP3naTX+oYMfMFxNaJ2DgVv3tPBX1KqS7B5eoHAyYO0+sQSxmR6ggqgH22yQoo7rUxt4Ssr7
UXs7uqVHwWXmYiatITxZJwyBnzyRvRcnEIHPsTC7JEvhBKePyLwXnAJRi8KIIu1hKN3fV2xOIvTK
NhtR+L4kDkMVj1PwLM/kiIrjeQ2J/AGF2tAX5SoLaBELCNPDlbfNNfpFXx77KtWyuaOWFDlooDF9
Rda/ms1qxyH32kMeCPH49bworW12YvhYIdy+7JYI/OHud5FbO+ueBqGxJHUZNUmFI6SnwuzhWPmL
E34jgbyrGt5IIvJz3dtCIgD6E3OuFELt8jPP7IRJ5W1El8VyCXC0saeurZl85Do0qE3Z3DH9183Q
q7HqyfqhjEj/EGG2J+HMCLlGZURNEwsJcVXMKblFQcNq7rTxc55UhprQRw/pI5Mptwc8aUxoSKdk
gTbFKS+++p+2alXlerpeshzd6+XIF/xrQ8YCv9UmfE6b0+dygazLzTLBkYmwJxImHn4tYpfW6kmz
LyGkoM+jWckIofsX55f5FAfPYKaXDflEhqUc1IB+pNXqGXzFNGnT23lvmIRGxUGrOhgqiHbjMdv4
tbQhKilaNLW+IJMTLO0TVdsp+x09oyVPuVMTfwYNbhxj3k80vi8jwk+XFonS1FAlk8SZ7gFM4VY3
15006PYIzECdK9EqQkc7WTGNlrGxXcaUZVIy6Qq5ESnCVjHY20HO4K1dLFmjGLI+ZAOLoBAUQvhz
+hVmXySC5NWw4vm2sZeWjPiWadkKV0G4oQcJM2iTCddt09oOfmhbGJvuGfn80zu1vHGD6uh+aCQx
I0OokrVdrVESZqgZ1jl4Nlrp3KYk1WexwC0nFMmWiv46aCM=
`protect end_protected
