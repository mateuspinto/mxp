`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12016)
`protect data_block
pHsHF9S9akWP7dqTZMI+wZSBt/nN01ZQV+h+Mu+eCOy9USVpmb3W7DP5oK2sAFiR18h0JUqgpOEE
g6wHxVaXlgXLr/n4X0yvfxMFkXtuaX0G5ecudrQxcDNaPNAfGiIQ0IWAqwyXlVzOSRwXT9xcZCRP
WyukXJlkQKbRzv6SCH+y1+ZuSFeiYaeTW63HIOQRzSSPyOEbGAwVQK0wgbblFP1Mge3+6l9rf9mL
3Smfd8x9Wa0ra0aPK2Ios1vPFNyPtETPC25PwQOPJPA32ufo8YTuWyZFHyjqPyLZbFKNozTNHR8a
Lvb9jgRyfoPqMA0LUI6pma+qAqnK7g643vGRqJOccdkUitI1T6G3b3b+/h6gvNCu7Px7AhuhUeQf
z4rOE5jYYzfaJOuuBeJMrwIcU/JFt8DMUX76LABthWBgr///xEHpUCFRUQ+ZWv09cOSXgtMKzW0g
hrM9TpFm7XLlb/MiJD3vgMxEU9tAUGX+Tyka16RPHxJYGwCOSJAo9lKo/nun3YXbVC688W+yWQec
CGNnvep+siLSKaY1RgkzV5TW8zz+z5tEpuSg1pMFrm+hYjj4xJb03sZQtAX+3q8Bvo0+IcgHPpuN
joMYMyn7FqdnjRze+9ipDcYw++BTVZ29vow8enW043rYjB/1zqEVfPlZxSefak88DbdfBq7Yeb+v
Cq9aG+ZekOFzeWdZ2dx3/a/b1qfHp/xAO2NoMzFJ8Ddsdt/yaIgdlaNXW7COCp8imCADZRRyehu6
qP+vuzb5+2MQ+1qmXw4EMbOlbMYNeFdqNDizCUJqYbk6FRdrR23Uq1rtv/T6hvZaeXxtCl9OxKU/
9odlhF4hvJd73SldRGDZ52PZ1p67L+QnyaIEOgDJCiRCFX8G0rgdAcJCyCJXfpM3Wz8+kJuCK0Ii
E7hFMhy/PBvwWakaT2xhwWyWUsdxdLIQA403UxZGAilFlpOHNom6gqnz5OXApW1Mektyv/SHc+6W
ydF0nV1DiHSwjbotA0EGg/d+YQg4Drm4VToAS1UAQLupc+ee7R/Ri9g59x+9+JoM5309uVa22nig
ZrwWQdirYzHGgfNqL6ncS6lYWwOB/4DrDHdjK6Qr5idFvwipEsIlraHdURGMloiCkWbMHejnedFg
P7hJ7ht6eIe1yUM1RG+jcZweqHhZdj65yuN+Hr3zf8gcDfxnDSY/meXMNUaXnZGzBis9Dc2gt57s
sOkL4UmU+7+ZxuotwHsc1z3IPRDCRkBK7176FFWuRSGQKCUqWsb7x9hMs1/vUdIEmHJ5QcQBW8Hl
9P0oclffex6Kg+JuZH6KrMJjmJpYSR0uomapFtDsk8Ant1hn8daSNz6thxfd9njFoUpL+ai9vBIb
OGsh07U+L6zMjp6mLCHPvtYGmq1LKph/hZfFfFxii7C++KUmrrlg8spSML6Q+CDclRxXgXJ0x4EH
82FO6qsM0T1H4NlBeuFjKf6VIMs0K0Td5FiK21ry8lF1JmL7VHV3fs7szCOYt7uMt3K/pk6e18hx
3E3dW9GvpwR7Tlw2JCswqYspSjKWY2qvxqU1LyiwOj3BRAXKXLM30F7f48pNz8N7XmGaYAzUkQ1g
Dv8wdkRBtmt1x8ce2BwjlZTV3FlJS2JaJSIEEug6aivbhEiT5xHmRLZkAtsFl9u+/01vfB0OwPQp
tS6p100fMH+DKUI0oP4LLeMEEaEycLvpU9j4P2q27E2Q/m96XTRrY0wE9ME9IZqzznpP11/gxYWh
x3W/XRaIy2Z0SVZtX46hOKDiKBImRHKbgdtqQUI7PXqzC/ct9oVNmoO9k5PgaWnIJNrGOtZs0Uz/
ecoS2A5Fc4zWb5m3Ynuo2NZ+qaciGcCS5BUOmWJ9X0XEgkeCGTF2zfVLQGLSenC+JGlc5sadoAdd
S0zFlJXbmtWWjbJtrIBc8zNAucndpViIfGyV+MW2W59IE3RtzXA0ZILLRHwr210WtjH+USP7Hn1x
1NLsOHx67/1Kvrnww3+t3hCgC2P8FVL77TBxr567PvWPjUAghDuXe0SUDdfyD7r76Wi4JX5XqHvU
q2CdYzaymQTotjzrEZrDp5PPFwUzFeQc5sesdcTjE6Ec2a7P0GFZhLdCcFOxxscfk+pxpkSoHaWx
5WYTlc3dpMX/f/hPeBUWEmt5JQ9QVx9mPNPUTtClxeVDBI6qkD3u06KPgpsBHbeP+jAz6tVC8MsE
mptketCLlJJtSX6nX5ROjmBwNoUrQHvSL/c+3aXSJV+itsqFVn0GC1r8uLosPlL1Xq0wu9olL4Bk
HasdGZN2OBWook594dIMR3cMOzBHBqx8tEbbPFOwXrZjbJFa3C6Vdglf/tmAvjcmnZfYOgyhWI9y
F9wvbLscI58p6/owDsll1XrOeJT7aGFCdS0HW0+SU6aaKKT4xG28R2KH93Nd9GcBFRKmeDoMTbpV
E3wYhrwc3JFpUSwTb0Qlj8tH1vvEd6C0YcGus7zcl9m/tAh51ex5zT8jTGC5MWXcsSTR+OBTT/Zb
ca8JWTB6yBNtNzNGW4nYNMNbKS7Gqfj8NFjgqvUIWNQ6li4A2Q3l9+lnzTPTEvbx8WvzSZpEJnXw
+uvJ74TDBbOwsmnTYOvJpr850OwK6NyzJ9aUcexhW8mJEzGnXOomc9rSqRW7PkaGcFY1kdJUeIU4
1Aiw6h/32tKMlTnif7O2Ki50Gw+KJczDxulCwH8pamXiBPUKQGJpLXa5kw1PDEZ1EFhTZV5IuyCY
w7fEMn3kBMIJGQl00+vAWGTI3uZ6pGx3F12jIXGvrCizqU6qqehDto6vJTJyEmk4HUAxgrwg2prh
dECQr8J0TLr4sJzxLN+/SvL+UgnopvWEeej3Gi0L+ZKYYnFTqt5swZdw5LY8EP/mNJutBLGZKGwU
IfGiXtyyy45MwH+xQJSelss0Ob/e2JRQSxU+Rjap9JqLgmjXago2LPEzUHaliajBjU1+rmwnV9mg
g6mWXWMvMuCH2+zEs5G1Xiz/oiT001elsn1FAa41S8jcilacMjeuFTjMNoXLqFE4cR1HJ0//VGTP
x5Rg8mbh3BDVz48NGmiWISEwtE1LYbqEcvQmeUYC2y4y3Jv2CyNgqHhrWSEl94ZFRztQZvf36ylT
SlFQPYs7fmgnYBMO0IXgsr9eQQUBZQGo/CNqCrPOAgbFsPCnGDN1w+TXUy0vMPwKtsUDO0+xW7YR
wrMzQsFl7/Gy+9O8xj+KWTLvrvNkkn4jKtHUSumZI/R3+yA15lylX2VAz4bcuJTlWGtJlbq8Su33
s+vlYQFe36JMNC1uj6yHrXJmGH3m0x4ZcP40FVy2z6TAv0eD5FoTBbhKnbZ2eCkXuiRqdYaHygMK
jB0KQpcbRJAulHK3vxIWzHxQ7nRn11nJQzVNDaQY/NFM2SFzcajP+yQaOZ+UDCGizyEJHeFVWjnj
ptyt3eWK57PHn0Tya2CMCUc6g00IG9Z6FbKZtOtND8b2WXOycOuRWitw+mpMVVydryxTe4s2K2BY
3fX7gRHCO9xwKkMvws2n8P+PZhGh1pk/tz7zu+mm978+QHHBJDqyuiTx47u/nCLCRsLVshv0yRhf
2dW/irQ61lWbFlFzy75j7V3Z90wf0bir1dQj4OZCADQepu7FWRErag0IRG9zlf6JBRHYA36DY9pq
gjpU1unWPdRQIAV5QAKB3xaB+5AZiywK2nzGNM2ls9qa6mMUS76NVUeHWGOVv3Vwz3z0RoJ+rfC0
MGNSLHOPcmEOvI3swWUePEN9qvwy/34JXmFe8Ky/FlAIiNVAAoGseyUJ+TSFiYMpRPD2ESe0oGZu
OrnYanUn/Un9B4PRmC5rykuiP1xPomkJ4ZstpCwHGFYziIPRzMeE/hy8qrr0RlvG3fy03Qb5C0fF
MJopYbneqaj14JTJYWEMsaw1CQnXVQLMfdZGYaF4Dlk104oC6Ac7RxuEilngA68hkqxcjiuHhhcW
LgP8+2tSZWRb2UXzC+yNe3unpM+sVehYjw+clUIqMqWnzbIyk5ARQMSlSoMLrbT/3myKP5Zrp5eW
bEWM1hcdakg1ZikDqoZBn7szfHYJkhbeYnrudoQ1KltoknpgiU9e6wkFAGOQQ5v2iExxmSt4Dibk
VNquJt0YwAElhpi9RKWv0EEo9y5J8LuGgzA5PkqhHEN7ICzG0eM7YkBV8TMkLUGHS2jh1n8W56T7
6IxuhwaZcK6sQNXsq/7I4Ky5npJ3ii3Ums38ohBlC3IRivwAFBjgEOLxZn8q2wvdz1v00w7M6vZB
k4DA7OtNP0WWMRNHyUouTAkG7jCipQ05vGP0+YXNytrJlK9h4FS64ChbY2r1RDc1AmIJ3GGi7o0D
Ed3vrTlwpY3g7VNUjWKWwPak6RmkwzK/IgkBOXeQoLCvZxJd8M6i6i97hFrF0EUds0O9/8Ks+UUZ
rdTPBq4bxa71tnWlR/O71N6r2iOuGNz+VYGct8fVQNwL6H2iqy4bI+Mbt0okjzeVzQ7CYMFvpnBd
UY28xHuSgRBsa5n1MbDObtcPOvFbefwoTC/bZenNjl2Dsx50w3nQZaYg2uThTF011aMnOuzZbY7P
qA/D6Exfeoyfra+Gx8XBeWsfvHnDSciWi+zfxhxL12a+g5OfO/WcJWmsC9m2d/eBqOHkLEVEShV1
z5LVaifinxChaqTrvmX2RGJHUnWXpP766CRfjpChKLca+Yt/w4zO15moggyHQzT9h19AzeTyX6Y5
cPJ7Hd9vLysyX6U1ecIB8ulFjeGIJMbOsD2zOi3n3ZYxIpepYDga1EOUR0tdUKvZWWLHsY8H4KmK
B7rM1XOOeHnjUjKGfqEsplCEeB7cV4vS2y7hWnjtk+Yy15VgSCeYCQbbGgSKsQYUflzxxabEluVl
M4f2Gv7DJWscQjXrL4bAT33qIyZZdoMXZ15C8Y7WNxdcZsTchw0GMm3agLSk8AbAsV9J0H/Jqzt7
/bUj13h+Bx2tuW1eRH8wKLoF3uImVZ6bCmo5cc8hZVUWGURYjrSdTcfejmRo+xS1EohbeJQrtgdq
KlHi//Tq2OkwRW2lZGX51Rg0Ul3kN/W7x3MD3+MHLy021tISAaRiSbgVQMBtZ0Bc13/t9SldwV1b
ChA1BHnXdGngvyaQYUp4YSrmQj7tHxbVehyZUVDbpbZebAGkwuC33epXMtqUghj3IhRGWssndL0r
3uqC8dNs9pD+QAkgDk732N7KYm6NPovKuoOsOdWIxcG9dU6PGmSehjr/owjKzik5wgD6f+U3E+mv
eaTCAGXnBy0uGYuYm3tONUTaizYgTWLxlHG/0s4KnkkaET09p9nWmGhnkqIpTFmGrQ/v3MUCba35
LDFr+hPMqLDH9goMIkFibZ0pEYMq+pYRPZDChNMsL4bzh3us8BzGFmAbeNJvZ7o2cN/SLvr5COQZ
O6Pwk+d7yvsmihrihrIK8OZIoeIPZkkzwUdRN/XEO5Y8Bs+8urMwrF9R9z8JPQ14JNO6UXwitXcP
yiXeWXV6EvUELe/7QPq4Tp9Q1hr48q7SSKT6K4A8NAUdu7fWhDBYrgIDGjulp17LYlqDXpkkjPTC
tKSec8Fp7i8d0l6bNmtyZGXgrTnUR1zD8nMo5XQNIVuApIUo0R2fVPkZVi7l7X7HqxEx0QvCw5b+
XCrbqCJa9LNiUSJzjxN7SyaLKaYOZMvkJB6ZbCOaOCjEuv1ymVBLClkmAplqp6k4A0aZW1MUeNVR
xSZLIVS3WDDzvx/38IkchTTl23FbPh0jic984vyJzTvUIBIpMP4fdPJUfpVJbhS4Uuh8HE700rvy
9CECHYFk7NpptXrqCuCyhYEJzf5JEPPKunfxbdOdynK773x/fOTXnRRTc0HyduTrphUS/vH80QNe
FFZaUtBe95YH4Zm5n+LE0tmx/8KrUEkgN3+C0h1GaKlQm3XVxxKg8B6pGjDeaJhERmF1pRoH3mA7
V4pq1/J6sUif1Pr+DpHe1Bp0+OL1EMPwyIy5gwd5bSDpmHJqmb7rfZ81EEs7X5jnvV27HoRApf0I
rLYG1LUcHoR11vbDji0j8XwLapYBo+h+Qt+fflD5Ko28XnBjLtyZPcWNxbE2ENKZBSjSEgIapihE
vdspULN1DmKbsWlUEbOYI2nRt0zI09EmjEhPQZrdOqO4Dw+91RxoCNOmCm74hfwn3LkH8tcxfWy9
j8+PAugcNZ0YwIucIQANOuUB/G3MpVq7cfOl0ZdV/Rr7t8WUxrTwrAHIBDOLM/DURORdvymLggrr
3mVhwqbVO8pcTC2jC5sA3iNa0MESx65ZwfAM89ffqOngtiKSUetE3NJw70I3Z4rzvjUWDBNPUPqr
z2r8F6dKO6omOaP0m4bmMQhBqL0qbawgmDxpTCAGGMOlCJ7l+DiZtNcw/lXciiShrJJzC4mnzeQp
wylwbwKoBkgCQ0ddXbfL+AAD/vFApg70Psxs848qsBAKEfP3DNF+u0sVGDtkCE7O1W/4b2EdezP/
8aFx+5kLH9D3PGwtncEB/eOnVWiJOFTP3Y+EVeg+1b7Aa4cyYJtM30Z9ZW3R1wBy1HnvZHahrMUb
t8g9xEPmwbgYEA9HIJ4AK5dW/Lf40nf2KfuUcS8EMXUROnGYAnwCnZEQ5ERd3Isicq4X8gx1xtQc
+vt2zstd4CcV9xFbyJfKV/tzsMCJiLSUyVb5UO3/YpJvpdiYsVmEqVLplzjiwxT5s/uJ50zSPzZH
Eg+se9+U0aBU0XSPHl1NhxVncZsuob1NAS0T3qJzYLYQP0O636EdHj3LsdDWZzv/AUXY1BoN8igz
Em48qmT6AqlwFpfiNoTkoL6g3pUJlVlAfegCXN1uNhTgP3sHYCGdaXzmi0tMTcoJ/DJWWKBaq4HN
IPbOtdBhbepHgKeJu2S03jwqWFeyrBkBVfZgk8UrA5AdCI1LiA7jS+kcb/cS9Sn0mtRb0vH+hPqo
KDEb4WyLszE7raPhkJmuMY+f5VsDGHkVqtm8aqMqe8c7HQ9riFByeIkhgzB6ZA28gtliqlj9NCLW
+rOHyIjDpGAGSjQWMlKpF5zcVv315rDmuRjKT6cqCPjboJbFarI8C+7wXA5hCjtgPbnQ99HzHeOD
beiQJyVdHnklWAlPdYYJgNG0lIKGH25r8Oyv9z5Ds0kt5q51xZRp0LyCSNmRuFYcxgA0nhmlzNrG
acMmnxD+cVJgIK5y103nd0SAONGZch9tBo/CAsVrtKzoHsNERhW+69An9I858pKqhWG6zDKyO96y
Qx5Iqz/UyKicMW3en2X9jZycvWajhQwVtYm1/csPgrB+2hUWwmcfP/8b9sXoPiC7h872BzNc6gw/
eB9e1zgYF/bIlAMZxRl/XyDvXQtxAGS2X5JW7gAgL2g9NlpECm/cQCe0/jDUF0lcC6SqQL2riMLq
YExaOO/P3uBd0URvOBTi0BWo9nTTry0mUQuBDyKwqhvbk41vUut1ERQARmDJa2QpSQHGpCMJEkHr
EIBzOhSWzg/b+ZxMSK0EVYR6ugXCcrO/HWK3Ee1v0iKugrVNDRwWfC0vN8cT2d6F3KTP8tmXgK3l
zqZCr/HHI9An5dMg8bPwJ6+4AxOiCzXYgEORP6bkU5l/86KtdBmDfabuOwxquE2cL6MOlj4+8Els
TdDIfw6j1zzyEMTn8ZffOFvt+lEBADSG0a4CnZkGbMD1qSkQXDMdH+ORZgO2LTcrhcOhWj5ZYQNe
f+2F6aYWcQROmJOtrASGBTp0yiH2r5MDwID9oa2Eyo8it0QcUozXaTMT/ivmi4Rm79l7KGS6Ndyw
/Wsza5X1su02CfeqRpl9lDWric1qMrkBZYpEZwmJ+NO0fNNCCOVAD+J+tzrYlsX8LjEKbHs1S1Yq
SMsd8O7OIi/V4mZP7ngbV1gFgmWcAqhzjmBoQgY5Kc3N1TY7SpYabgJvQzv3n0Jx9XAwh6qBLwGQ
quiEW5mPTk4xf8wL1UFPt/cEhTZyX1U5MrOv3xwlWBZtYeJ0peD8MrKaJp6FyDEhNd5ajw1250MG
bJ+kUN97hcRfcCSfYhmt8PIC0xVwW1KxhwoqEBoo8Ib4UigdtvYMS5BmbvLxgNJg1iHgUEzAKE+B
VCSsoaIHMYi1/+V5uKb9J15vGNQB/pBi+OMgXQYjTlFaKJjY7e+HLVoFnplo7nFJA2E4FQnRF1pq
CtohE7BVuvRt7KdCrMQkPhvZxfUbEA+Yx2q5HEVWIsnvDmX1xPrU5oEDfhLUXPFXgPu3+qasDSr7
e3/eHWpJnAKJZTcMnwHwbZtx0FHWzEn8i5pH8WMaOvmdWUG49GnvN7njCv22XKpGUnIYfuxbuKl3
Kt9CbZ0sFjOHO9AMwne7pWMI0XSgKl9y9qf5z+7XbsUFzTQFXuK134zkuqYsAkgB8c1MsL0g84Cf
LFqSlzMhJZkbMMt5wwXjURmWes41+GzwgOX/EhTcZANJp6kv1gPhAeYfBfAHRjnv3a3xrTfv5whf
yJrN1BfuyFKv9sWVyN+v7m2B0AFyb5Ierg4ozI47DtbvHtCTsra7D/CSJdvodrFAqlIkOF1CEsHM
Vn2lkNyu180oti6N8xMotMEMEtIrtvYW/ptDV1HT8KCWy0S8qeDsUMham086en+sQY6wp/x/bQt3
V1YjvU3UiANQam1bBvci2yJT11HDXFztKosZGZy5mOv+DB+yJ0bWPU4ym7lzFSqtcFQHaFAiBGcs
kSBSUD8w9gHxVwRGOfrVGz1IE3NJ05UUgZmIrEEPb3qWwOQOAhIx6aonMdbcUV6FXzn5aokJxe4J
AN2JbP41Frv0hhyo53C7Y+Tl63Q2oG6F1n5FBrB7m5IbCLQdDm9yvBC+0/38U1vry33RwQHtORMk
hRJYFTAfllOr9F7tJ9HwSqNAHUkD9jwt7md1bOpn7+CFisyOXu1NGzIxT/ra9JHUpWX50S1ml7Bu
rbyA3IzxWFL0QOM+EwhzTt0YG5xI2m9jOPc3cOkYRRSQNBo1tLs4OkBnWNcnom2buw5V6NWA39bp
4O7+VplH/W2tEsNQi9a/AzvYMfKa3mxkIkOGoIxa1kq6QM6vyCb8fa3XcBbXpLKY9dK/S2uYVd9Q
nLyBjlIleT9XJ9dPZ8KIezLce++J+g6k33XUoKh5g2tvn6DYeCygein4dIEky8iVDhsE+en94tuu
Ijjx/QhPsRQz0bBPvXkMCIqV4o/SCy7cE1S7fmcy3aiWrxMzYNBnnLRzWvEyrV7CAWUhGalgiYCp
Xbj2WKKAvmDxDKgaom931I6zU9doJwi083jdM+7aCqKFcIsRx3xdu5CBoUiAeGM6nZGzBjHmsQMU
1Ez5MNlNHJL63LXhIqst0057yyewA+hmudtlBR+RLC+pWyTxCLyWwLb8EwSV/0Dpy66GHzsZB7Bo
wBckS/DIfICYn8i+MHFbAPJDwRiup0SheDIBrCs5te96E9UC5ND3yj6CKYeDKjUsRJK+/HkNYyUI
W7dWqcJXDT59fj7RYwdapgRliuC3ePEHabJwDPz+a2fhI7/2dIzJk1OECJge23G7Rgl4VdGxJAZT
4jWLhjW5H+wVsYsgNHiMr5oV3Ai1zUSvgYZlc2bGcxvxF/bevOSzuf5rObTM2gXrtNUYhQpA8/Gu
m90NwA7qGQuxe6wL9aV/YKJa3CdKzzpeojiEqLDil4bbIyVksoSguKqF1xIhN7UVP0dbKGxbNruF
jRQuo/MuRo81WwNLzBRFh0ONgX/G+8HlK+kf0TdpYw9nzFTYZ4JtP0h9WxEIaOa/Z8te2LJwUB17
1ERNWoXMyvHQjuD1o4pLZgoIZO36jdNpfxNPvwLtS6+3pziMlV1MyHjt8mQhLP8Eb7vtG54S4u0c
Gbtj4Xz5GHbSUaImtqmZ3UY5Fqyp5oNilIXh6eRNUXZRnXmJM2J4gptwbLT99qo+gsx32DGGm5iS
JRuE6Wp2IXEfEIWBTPZwYbj8XbpNe1BciOB7fHmA1wnTB4n/HwZ3w1NNFQG0DksDzdBF6NHzZm15
BsNd0wtML5a4cPoyAe2mnLCPYN1zkF74JzYA9l8dyV7GEp7DKZUdE363jHNMg0qbxPTHs7GXO4UU
HELcjjJxdBIXbYSp/Q4iYJg0O1mqQ1ayf0WVqYh6ywSJcA39hnaRydOUHpyfqPfdCrNa/74UENnM
WqrE8ZbTiWTRbxW67kaOhV5K+aOiF2PMbzrMDCCwTTUbLzVYiSUUAFtgGvHFOV/mE4K1NgQQe864
NX6fi62s0/vAFPlBtu3BgFMA1mWIjT8UhfXVzJJ5xcsyOWl6Ksil+8i+WCxpc7larKnz4IXQAniO
VgTFcLXi8QNW/D7VtWPwYbeEFw7dv9HRPumZm+QPHxYR6jXFAj6GMfzgWaNH5oCEHW9gWMGzJmSo
56IGX9uBjuCYV9rLA23/hVG/Vny6q6OhfbH/qLksBq/wI6ur4JsIi8bu0VSHvV95hcF5gM50T/gb
z7qHIGiPSpwmZH8UgSlB2MUfKZKFbWbJADbnwvTHBJyW/fYA9XaSFQTBtFGYvbYwJMGi0Vbs7hAs
aOyK4fjrBYG6mek5Ou5TR4TBl2Fb0qb/VA0FmtzOfMIIhhCsBFEfzmTjVDhVjBFA2G3iDUCFqnBd
t3l8yrkMWE9X5/Ie5X+Bj7WRy94U8mhucEnYKUY8eicRvFh48fbKpQj5hjMDYLcAV51E+ouCQci3
LKcBvUGneFtbxLYdG0i6ucmHUwtxxOxYdW1HADvQy0FRihFki6XMC5qKQl+Epa7ychkAv2UqVXqD
SN7oZV3ucU2PzOUU20LSdxOshW1AGNtZaj9zCnzkvHAYEdEyxaCZiCQ/9jYPbukUwFmktZOdoK/A
HamWmMT2cWg28U8Kfbl+g/SYKP/vhsJ5LITU5kr3E2BOFujKajcmewkWH2TnxXyc7XKdxwtjTb/G
pzLNVLaLp5gJnfGfUqW+tBnDmdIkHRXSCDC+mHk19oFYgrfPYIRu9m/eNJoFsns6+X28wQcEGvMS
QG/5QiDkgdXwJF36Ftx+HAr87rV4mWxXOEl/x0KlF7y7lc1CXjePR4lf6BoTNpmvtHt7M+adtCD/
s4JnypQTqNVPlXKJI3A10Vwj63L708FZ+XgakF6/ZkQk31inGKmsbtNe/l1E9DeXQzciJnMcNt+Z
qneIVuXqIW8W/B6+69M8bjX7MCi5topjGeU/TDfjNCYlbKOyOs+0ohHxlMlGhlnyN9qFeeTvT2Cm
GgHS6eofHoz3oAilzC9ifAZ503Uwu17Sk2h0P9Vft80bfI+x4kEV0k7FtyQ0BuUgZVF4nN4c6eVu
5rzURwP7V90ftKq3TsX07g9JJB9YLtWepQlL4X7T+qyTWXNdrA3RKAAiHh1Zvv/sm8Uhcf7XFjxj
y0dVQ4v0e9nf6ptRfO2kId+DsSqMfYb8vEkbx/HZB6Z+5rxXwwRNbjglLkfDFrV0XE1QdDVWN2Ol
UyqfMnqZ285RUgJ9mKz8uu/s9MAczdnoao45yzpwT2vGYdBjw6/lh5r5wcKXqJB3cqXQl5qYKID7
05K1nkN/Q94g2FA1H75VjjPdM0qvgcShUdZpwHn2leaj1+5aHQTACkblTAs7/Ftux97JgDIQs9yL
8ZuqKBCFvfGCvTdT30R6HUEftWsytGMnE2OFIXBPc+9uLZoJzssXTitqYdnBlEY6+1GbrTTNvaKn
h7mYnpzGIgZVyLgES61S38rPLX4cxEYiRYEF2DQhOQ+OdPkD8gppx3lPQZuUuh+bgeoZ+wwR32Cl
y0gOx9/u4Pzc6cOdSscRuDAw1Y2W/veJlqKfog2Oycqti9mOCMkiO3/D2EV9yvbhlg0UAJl9h7DQ
8qAZCQ4043ZP4aKHK2cecdLyMKcWeo6zNwEnS+t5++Duy0BMzuUlWP5RRa6ryFEGLlgoYL5JVoNm
6I/JRMYG7rPO0wL0P9dYz3qzva7D0SC8Eol3aqpr1GnxnePlk6/sniAy7AlPZuy8WjQ/vSNyBEvZ
zvVTd9KvqGI7ClGhYgwd83euKwHmrE/X7LU4hsQ7eQHn7ijm2UXMBsCqC3eCeTAMbJECyqWO8DnG
7f2Dxw0mQAe7EmOb0+09I0XGGdzaWE4VU8ab/ruodKPCbNtukeucp+eD5yIoPuv8fhUfZuWiU0xK
AfzZbovulD78kx7e03NTyle+J53V29GGCuXwi9xtNYTBnJTuHSk6wXO0xtQnYbDDAoJaolaswNtV
hbPJ/OIH0zUMPPx4wQZ4IaIsUOB/SzGeGWISEhPoCSfu3gFLgY42MeyQLfbMvk8jvurvzSLClwa2
XLdmGA04SKYZnXpYjsSsSosrkh38ZhEcrzBCBgPerDM/iWrXLBtKJ9qbB+1TWz823lVTf79DY6ae
/ayyoDPoqUzHjUq6HW+46AIikyos3hQuGLbRcDtEyE08xBDGZMnDJkCFWdUQ5iYAkEdn1pTBFDJz
TPhoxebio7ZzWHQVTXW5y9yMnxy0Jl532ImRzaifa9AlOMvsDqYFVxRDbguUHjnTpyNPKif7Cwj+
tmnfxSQmpP3CirbgkaEzW+HW+ayQbTJ17O8Sye9bLYxUgBjj67elyFwjfv21T82ca8J8HgaFrbZs
qo2ucsp94souQs0LTr+laQSIZtONxhQyj7Ps/Wi4UN8eIhwYn8zPeqh+8BYxOYtXiFK4b4jAqO/p
Qk37Twf2TIyAdVzFPeD69hFvKq4wltxJC8s3bE+5zRV69qX7OrGyw881jzMnd6E0FyiRWXT41/DL
fuY/usD/CG1lpp8g8/XcVtJjiEMwdMqYUDiSt3nM2NFnBAupE4ySlkt40/6Fic0j8RcrsGA0UvcC
+EvT3swMR4ucNscqIS7etcCftZY0au3Z7vYfSYT7zx2KZ/sdfUgm2gCYVNjv8OpcaQ37qOyFrpfR
b6vq9VSOCoQLhYPRRuELaCtU5KKaldFcyRyDowCnK7k+lLXKQNimZwKTb0tzXVVZx+nzwPUIv3Z0
yah2ZJ1tHDNIPEhCfmns9s+slhoZ2Gs57EPEQehKTx/pU80MuRUcNxNFFlu4Yx/qoZHX8YiG/R/g
V1Gwp6bp5PNtsAqH6Te4KciwcEESWNNQ6Xh7GIaO9cyCempoxnDX5HqyNzEq8nspirxWQWfl2BZF
9md8dg0xRdhkWpEQpWRv4F3OdPmKsV1v5VfLzv9BN5WVyLUfFwt0xCg8CJ/Sfwn5Eqw6lyXAF8md
0PJ3V+LyDDTqT/5tkCEfSQiqGEynxFQ5FgleWw5B6dKMgfAmKyovVyPEtk6jO9lZQ5AuHZ5Uz3mg
uBzcffxsagx6EChF/JhYKSQg9DvJ6EvXvIMQHPxGzx4ddj4vcpmbEKVhbSGT0GGp0L5uV6hGxHFR
3l0nd/UZQcIs5IQUFpQVPW8idhoN6O76qVnywo8OZ7+gr6nhSAtcWakIDgd48zKxnnW3unsPbaRQ
NPyxYNrI8pWJWB/1iKIQZkOXdt+Jz4kiyoDoCERkNlSSpawGpsBw04jHvSX6sm92WL/2KML+4Bqe
apGB9ObU3S7pnLnpg5p2168wquXCwt2Wer7ksCfh8B8TqmbuIkqxHJ4wruL6uZAoyspyyDHAJscj
I/YSS/62c/S7KrTNdX1zDmIMzpmPlC1boBYQD78yfMyvMf6Ezmw+d2cSMgOxxU+8JZhoPQ6uXU22
Nz5W2U3Z3OXuVi+iEH65odaiofrQepRJsIEGjmzeCrVR8ksSuRavRI2r7sbFC2CYkIeMHDAYSGMf
w8nkOoEyTkEY0CMSAbaiUBjro4eSqwIjcYy0bi3WsaDxBPVwyZGLT6sfoRQiyiDU9nma0+/M3fZP
mPEbw0fYwc47KuM8aT0lQ7q2hD1a8fz15NuWfDhtfGEkYdlJi1aCcVCIZEDBAnDcm82VLeHuDhRE
kfR+4HhyS2i7g1LAxiJk1lB8Px4zS19KpR59/CYBd6UfmpuxIUbSkouUotr8vHuZb/kdlHLe+1gl
XH/dWBwzzjHOnT1RqReuTeZMrg1D7whiUrqMkwqhAoxHE36SADvzyKciLPVYLmoXmaf1ii6WCvaV
YdGxBCTM0+UcKModHv3RGJN8F1ASIJkk9WrTAglPuCo0Rv3hjhHmS1Ida+cRUs+KSoOdzWCa57vD
MixymVkDAGm9SBhuM/os7WhLu7VQUXpfNjGRA/YlQRMDJmRb4MfGpeFcmcFSJrcHe5N1OEVQrF4T
DR2qkT2xEFQXo5P2f1ZbdWw+xrtWS4D12vFM97EZQq70Nfx3/QdysC6oMUlSf5C7AO+GXZHyxq+7
ISPJUnH89+6Jr+NGBrUiWTpVokTawvhwq+QFkHT35Oxh5QaOwDufTyEsLF1nkx7SWlhPVltvOPW4
M65NvoZSflCjocVlxBsOHMUSq4FIlAI7tuQl/30psl7DHdOzGFg0HMMtXCyQeZv94NakSFgDWQYJ
xxwgZucK03UAWxYnla/auJ0Y/8sspwofdO3WprdL21DTI/REQUUNhv1halQmjgcCdR/WpIeEqz0H
nKxgJ5xRwgWf3TgNP2+uy7cuu3b3Vh7ODMCqlFVf0gc7vE9x9tLP5rrGOoYk/7XK8FRfQs0WY3VU
AYJHkvLmqpZKO3809kRZ9G+rUf6nL8BaMIczEhJ5MT3CPyakKF8Y535iAgqEv0oQYUxHwdU4qzmu
d561CFWS7nClhmEOpZxzpyZFYrCpPMCibkBXpiiC6AeqEPUiOpH9m656Lm9qRlks25e63gykm4eP
FMaE6a/lG1SFGRXw53aVUskK+tMo08ESnQcTndXb7LJDWQaAupsk3QnupmsCW2YQpHLQKGk3qKJ6
f4Q8lVfOj971VExJ1jcJBJw5nv0iGLVWlG0LKjniMBEbWCWS0wTaYpapKmGuHrUavKOXzoHriN2R
pX6wFR10ul8GwPt7IrkQb2tNVuHneH6cT42rWWa2nnL7+moTVOSzuAfe8EydVL3vQM/Jc5CYorFj
BAJkpDaqZ0nPIKQYl2vLq2cwrb46kNsRdMvtI8aTJ2otpy5i0LG14Uq8eVx/9tTpQQTAK0gRYOeB
3LmIIwi23FJ6fjdWg9+7TEGplagu73El8bR58uEeoNWhKg32Mp6Hgw49Zq7hAXgBZyP2WeP4VWCR
ub41I/mp+pE/edfx8yQDwJpcEaP8O3qoVASVeBiINukcFwvwLZFysErC1FKK9GoJWhAGo8C5zQlq
Z34BsSt5Ayk2fPQ3i9wAlDiGLNUiK8QZKcaH8auzN16CUN9nxtFcISmUoXqDtDh/zd2OBT/uRSOo
cFu9b2WnpN/3WTvjM7vb4njRaoRwMAGIVggq85MpSNEitBtyScbf7CPvChr3NhgwlP7/7+Mzdu2y
NjHK2GKaf9x37XGX6Q51c+euxKwSkHTdjzaLUwSjkmxZqUkFV05q4Kx5SwRK0S+n86oa+TKQBado
0p7ATFt2fVGyzpovpuaBIMXAccp2JgIaIhqv2WysnDZhzE6z9Vgo2fbC9ly0qEV/9rhqD8vwE2tN
mpW7or7lJH1K+b5HoJh0MV7SGMwXj241CqNdBMDbKfHzamdsfjDhRNF1+cRhHveZcUDHKGVY6vTD
0rwnsPkD/q13/Bohenzyed9ehIQXsWcV/2uuBXAkHkfhfyAYfNd5tBMxGcd3JHuuluc12oYvS2qf
11p7PoICkiTIp06bRQKqFGfUCoTqZSwEdVIpKFWMxeyXobh57Uq+BWD8hCqBV1xAcu0YWL3dkE3z
PBUj6v2vH04Uk/uABuQJTL7vyiT228g9QhmCMxktGXJtmRSD9S+VGF2Jlpsir4dpH5WiyEUUDHby
R8SCo/dV749epXgApsX36bIuJ5edwdDMQWgJf8+YumXj77bpNWry7HFyXFEZfeOGl2J1C4lbS8ej
/ND7ld1+FfHuytlMrD3ABuG8vz6yCMsxEWzzaWttpf1ncShifLrV/jhVNjTsG2ruyh/K6kbHzi9A
u+6L0IVeJlg/CpZkVZfH7LK7wCmkUpb86l1Zf2sSikaVi1ik4Pjnfe2xluQpSBtfHywMAP3eXkM+
IN/rzwkrPaR0TCKTY8TAH61UEc6niURh1jJn0zMscnVAumutvPhzhOURKV2DMg==
`protect end_protected
