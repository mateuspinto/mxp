`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`protect data_block
58Fw9jn7zDyTA9jSpR5E1y1ZMlSHtRbwMueEPKkYNKdcOVbGAHTnoykgD7eangymV3m3wBHDD1tE
AqCDmzS49l5TIq/ZamANlBZDSNkoXpeWw4VwXAFduOQpgCTTU52WAWHfPmey5OBYjXsnSTIzVGls
uinU6ZQR2el/uYTKrYNTEYamvDtJ4vyBcCSTr6UvUsVLUPfnz1+EUEeontIIttZmXSkRmAjIGUnH
7rQLEEwjTnYfSh1lxzfL/4ndgKfH48vAcCSysWwT4UkfV6arZdAJbEsI91neLZihXXbVMTHpoEKA
UrIBYtwKtTnn8tWCsEmdR9AAVoAM5JjSoOUoH7cu04PlqrBAYbbBElfxTJOlxJYXCRCb1WSNmIr1
i8TcGji9hRUFCPlpJtx56jji1DpAY3dPyMJiV8IxLyFu3Ui7v+/8sXre/1KCkZKhPsYGlKI3OJ4M
yN64oPQUwBWA0blbEvZC7QbxC5OK6Dm+BKKmUabcrBsz9T9zJIr+YzUv+j1UD5UIx6cpQz8lUoII
FIQ04h36BJ5PP5WFbIzmoJ/QjW5AMrtAbN5KlE8FdnWct7T17dktcF+cmdE4S/XhQO8iIZ2+OKXS
aBAre15bgIYdYORE+WuGzJsWgJtoxFUmiFaZ1nJ4djJqtL78SjytShCwnlmdCSy06QR8f1YEkPPZ
AXcqrrgClnRMmweMZbgo3QCzSj2s8Q6u8P0l6SIut8mjs7Kcg/NnfoqPBWlbsYD0IyD4Pq33s6nx
OAbV7nZvXk5MTv5juvW1bGEUI+PUojAVBd+Ln+iVMMhHw5iLDb1P1WHpAZEAEI+A/wIbLe1mtOvT
9m7aqxD4DZW8mmdxoOgBl3fmi954x8V0xsv8NTWPHDtGV0MnSLti87ORW737R8sUpOFwxhR5BG9L
p7l6D6+aSe9zhrsBYRU51LEAqX2GhV6vc21/HC7p5Mvd5zUxUW2yMRSse+8vXLbiYnqIl6TCRM/B
3eGQ3ecoJ6vzzbXOSU7NsV5s8iZHF2R+yp9QWPGoA9exTDoMpxOhTsXWpyigupkIrWnwTCh14VDl
IJU0DguaRhLev6qnIE8tQ1bY/MEw6Ig2/QCnipoq97gQmLq1sGgPmOKdXpKI/2lDSoZHRkYj2ydp
A1lAuoR/aRU+Du8A2syRVo2tdvTszzfG7CW3V2RvbCew7RDDD0kIuAUwPu7e8yyoPVmMHFqMAsZd
hK3qpxJ5FbZV5nVwJ5v2pog4f8kADQUsmaWxPRBbxJ7WMDa/nVa7/A4ZtY8f06T+NrVXcb0meP7Q
VKGOpkn6HmMaw6KD3lzOsNCJNPmw9TegkymAFpwW7VsMqHvvFWdMdBWT66/UMjFs4Ac3qFdImoiG
ARgU9t/bEVD8T0Uhz2e6NHwt6aJ/saXd2A7RYy4wb7RgS4H9JwFuowr7ZwFqphtWVxTipVcDPHw3
HuUPPOSLoh0HA8hdOdHc0DnFf/10QVmdRwcCZQiakU0PqHnQW6xplo1GMOgCrszDNm8whQXlVlfS
Ej/m9oT5EDLBn9tFlgfNUPp0VLeBhnFSXAapJCot+CJPVZ2Ec+bJd4YTrLoIQmGvRohyjO5NORxf
rWsM8TZGqxJEWByxodxCrIcwCSs1icL7tG17uUmlYbTAf1S/HAaCRwwWUwQq2ZHRhTGy82QLsWYW
t0ew5Ej9n5EW39byWavEV/WlD6lw6Qt5QCGvmVZjll6DqpQtm7LHjO8qAdCwB3C28osoz5XdsUAL
VaXWgfG0UrL4EK68SBHUqFsU349JTFqcIkzbLZtTjwVO6qmcKKGpjABoR4Efqpm4WFlTYQ5R46C1
SI6XpGJdNMj3zdJlFwpgcllDPXstGtWnxZkS5+g3OV0mbda153Jooa8le1cOV1bv8agegd6+IHI3
9ZJUd+i5IRCbmPxmz4VY4yQW9QDIdfcrGPB8VhzeSv0uwZocob8yukuHcOrab3ckwEwy5fpxbNMF
ZyPE8UH/Redt3mXuyTH6xRo1PH3BfRQjXUP0dWgHzBVf7XqjiYg30UrFj1f7+KgmMtQ23gVTWL2m
9Eml2tT0Vmx8PcENKtsqlbllH+FKgXh1JhZ6z6JPlCRPSVLOFhaIOB1TLs5FnMVX+2Q+mWTlrq8o
C5nm7hUfL2YYKvIuVecgImJ/Ur6Dl51WdE2qZ7O24gY1AIfQDL+2fNwISFkaZpuNHcfRGXtKb1YA
tFCI+B3cNJYSY7PTC7+kUFajWyCvwutKJ68KEa8J6esGrEg3MuwV9qgMF6KHfr2XLii8WyVps/PT
zswgAeVY/BIULjfh6dRghkVty+21xP8/3lUzTPd7+NuLPXNwP13upTmJmVhz8HGz4AImFqaC6M+S
kmmPQaBLXD5WFNs+yw6unCZDg963FekX3HJtSBp6jeceHBKFsJxHQOwdfWI8l1T74pWGkuHo/tnq
RJJKasupIjzRkZIh9dbFepSuPl5nhIipakaBWp/hwVUp7mmDXvFa8/1Vl4H4RJf/X7pyQXyCf0IA
MRguSaK75nyGx9ubktNmRNYA7pp4kDujDJHhaefprLLm1lWgFi5Br3Sgwkh6s2RoFBUEdqSQsg3W
FcwRDTnoc41icTHbkFL88LYJuRN4l39e3SRingvNzwGw/eQT8+u2w45T8MuGZIM/OdrsOw5GKdLc
FcLktZfxNGDTICTCJ0XRSgYDayaCc+e/ZxpUee9vWJaCKIVXbDQRd2WRuPyski0M3jlOCz0fuHj6
p0cznEpfHZkqGpGoXLYQVoqYH5oLBIXt1IY8HTduvckX42xXtMoNyVhsAUg6L8p4CxS3kPAOqMzQ
f+N/3wgHTCzJFrFLI9fWSusZYhr+cuSWqMuWrSx38VpoGRpPIypq1krEXW8IyWnLhYN3zhXTOJ6F
ZBdIKMPW5Jz0m+cjwrrIDSiiOXKAsm2JPYGwIOSKXOmKgGFaguwnrHXIanoUPDEAqA0cxmFbLYu7
H0YO1uUtFugpzHI1zgDFP9YXzuiTEaitvQe6InxMAEe3kM/xIW+qtzD73g0CQcyujuIFKcQ+KVYj
CeYQX4sOcmNxQ9YBqddfKqefihsQ1rP8zGBc+/9gVJkU4Tubq5Z1zMTcB+BIdtlpmul+IUc/4oCd
KrDIKeZ/gJTcwoiz8Xw1tCF/uf30neK3pScy/9cuiYkNCL3TiuU0MzbFwEO0jv376uctEwL3VsG7
41XlMB/fGZXH8Qn8yIwnN0eLC53NNUknVppkctqCWNd0tpNKjKfDwea4jYFrrQxd0OH57EBxvNgZ
aYeQ482hqwPV/Qr3SkGUa6zwAXbKwxsTaWADnslUCCmIi+5InmjN7uKHxnbSDfFf84OWMCjf2rSR
gdOhE3QgyePvhH4KkZMI8xC8Br5jEgytXpRthkmRZsDI7hxK0FaqJDSRAUmAufDK7Kd/xqyEZ1j9
cizCtIifHqh6UHl7QBuoVlo2ADsAZwp9zJqPUvK1NluT//pigveE/KJ2v8jDYwoV4sk4YQK9CSIp
tmmhOV4/+yWS0jMSXn7d3Rq2QSxDhh5EoNO8UOwnE+wsXxuCVxcP9Z2HqqJFyTK64/wctHp/UCDG
OVggxLpy0g+p7glav83PIMiM8VsGh7XN3xggksHWTZ4mSQ/IDsuaSrCl3jc7dzP42TsAqiTqd/nd
1+gfUGFWIFDMB1uxQ0hDhiJjp6oVVRee8wVgW37OdLCG9cM08T67GeVvBke1M1zqs+Upf6Rt6gG/
YuEhvseXlMCt2FvX8QpIo1PgklqlGAKIM5s4Kf4ouXOjtpdMqU/UQmUaYanBcaOthRYEiDgO4wTS
/22B2s9Hh6GWHHQS5bLfSOV9jzqeVOImZV1WvKNt3Cb0plAfUdMn1kH5fBKqtknJ0nsKeTXRIjrE
/7xnN47YDghnbUQDFGEBW0ads2Be+t3n+1tKNJoFGJjGVdvO4xWFxiwUpLlA9uY2OYzoNPRdHgd3
giDNAtvc/JMds1X4wQrci1uaxMo8qZkHhi2ZaEyC8WlkgDCHTC78AxtH2pORGgEGYLzw8eF5cQl0
DuDNd6VmNSJwNlK67y7dOKqCDnAK+uS28ukTAeIAsnl/CAFnUBPnqa/tSAjxbMQgwIz1IEpjKNfW
ASfppPUyZvYHJ+9ZbU2GuVCPmagi/D75e60+pqHAyN7IM6KUgKzTo9ElQG8dHOnj9M1bgsoLVtrR
6wmQ3BqmYNtvbmCwmRw2hZjtkSsl5zdckcibIfm8gTPrUX2wUoQu+OV8kBXXemJYS2r/la0T7IU7
iRL7TPVAYuWh910nNQj/WfD+G4ZnV9Vw80WZ2Khq5Q2Pa/zSPzvRRPnyGETscYKrZJvzy9GFgkTs
t+wv6D8KkmwQ8Y1i/3ieNH1X3YMwyL2oF6NdT2YSEAGz4LvwuHScTG+OhXfiv5aceb+pAtVGmbU1
322nSTTkoehmxeY0ES549eTSoY6AKNseoq48GJ9jaIvZaiMOD9dBATuWGhKu2zX+hMDGwD/9yqWA
FD41UI5YAszgUQkpPSS4Emyf3yCAEducadFgxSs0An8WPlpVbODS0iELCQwi3Ng74STmTF187mmN
tK79BkFa9OQ3n/XIPtIn7KJNcJ3MNpfTqjHlWCgOBAghAQ4QfcOEeFc738TpjIFI1Gg+QvygtFZN
cKuMwNfaCTevM9BMR6KBHoQHSwSydABwG+Zs
`protect end_protected
