��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���@�ct�: �t`��k�r�i��ʳݴHEL�
i�ޗ�d��'��p�bF�P_������Edڙs?L�u5��[�_7�o��߯jĺf�m_e�	]z��'��3�y��:�6�.����x��b+�큔f�ǻ	dR-�F���kU�1Ѯ�Ķ�����~h�� ��@Į�/��nB#|9.gA>&`6,ܕ[S���2*!��K6�>L�Қc��B�(�!�GH\l8sY��n��ʛ�<�����σtU�V��og����$�o[�7%+{���D��Tz��+��=��<�˓k%�6]P���Co�x�X9+��.�5O�/؄� �SQX���}�|����G������愊��&��-�%3���ר��6���=v��R�=�îR��ĵTFp��ȷ�&A�؀���?�^S��-IBE��)W��_�h���}?�� N��/ �Ұ��n:jǘpVeF��jG�e��z�Xa�z+���ks|��-�he¸�Oo�4�]��8 �|9�=2��`cHeE*n����K��q���p�z��\�ZU&���9pV���X��J����ѷ%Q[Ψۢ�����N�k��ng�a����M��=5�t.��U󁯀^|��ȗS�_^��`�#�O�j��:�N�7`&W{ ��B6����	CU�ھǣ���i� �"�5D��'V%�탼e�]t�w��z�܍�}��x�5T�m���w�Fn�G�!�/�^+>gբ�X�Ȃ*�|�
��V�dt�ыK�$�D�_�8K�gF��'4S�=�;��`��߯�;qC����L�4RUR65�պ�ꇛ*��q�����Y~���ɻ�ەQh���C���@��@�6� ����ԃ�'ml�n13^S�U,*�l�o����7�9�}�e�գ�� �������1P�()7���p�+<A����q�[����J�$i!ʤ��ے�
�כ�j�q�O|,�����@e#j��j����-Q�{'��:�>B���JH�ehY�R��J5a}5
��/��P��Du�Y	aH�*ŏ8��k��g#�P߻2�-�J��# �7�O�wC߄�M9�o&%�q�����E�!�׼z>���zy�b'�%z��S�0�$@O_�X�P�Q��R0���nu�R}�-&�S�Pfth�ŋ��z��V�s�24y�:�a�؞��|Y����w����5�G_@0*���b����ζ���JE1F��4� ��w�G����~��e<�a������j�sB�ۑ.�6m�n�le�F�M�=�nL�b
/����8������[��.g����:�����d�1Y.�|�kpՊ��p�@�1��җ�<�7���f^SlQ�5�G����.m���W����	�n|����X��3ԷX�ơB@xD��0֔[�d�Zc��Xu���fu�Z⠿� �O���"�?�;2�����&�;M'��
�j0q]ݛ��si�Sa��� �&�9��jb��2E���Lw�d�;�C��5�r����Id�D`��LF�<(��-X�FՑX�'|���J�X��������P�D�Y�o��;�'��Q�'F�ē��D�2�]�.}G�m^��S�WA��O��ы[�&����b�݀!��ބ�����7�4�Z`�cs�f�D5��xukVsp�{D�P�~�M�B�ȅ�o1X�Õ��$�y=d�Oy�[���h}��TS\v
@ͧ�u��h!v�\x�-Z��]2*NsJ�Ŷ��[K"R1Z>����ل����琅 �	zG#@N�v|�g�)|ޫJt���4�h�jiMCN�e��d���Vi��.�i���c�u�	9���5ڇ��+�X�.�8,��5�J�5U�Y5f��yɝϤ"N�w�ơ`�m~���`@�p��mÄ��Z�/��7��h�͇b�Ae���:7*������3���3��V���dM��T�i���ww,�񢹱C �� ��Yd�A�}ГC����9�̋�����ߛCә�� �A���x~���0]�[�D���_KQ6���&�̊e��j��ɧ��/�[32T���B�ag<7�(�����	6�S��G!ZR�Z�u�����־�u�����B��c%�{*E��)/�[~$�oG�*1R>D��ǈ���E��6/1��,/��5��Q���%�*�Q����F�n�}t�>WY�VB��_�\_H���ϻ�ȭjyV	z�:�,L���*�Y���!V�u'�;�B
�p&`�?�H�#�4rɹ�����-���Ԩ/��Ā��t$�Çx%P����5.|�H/��������� (�c�"zy������C�N݌�p�xx�(�z�n�� Bf2�^��:���d�=.���z(��y��B0�J&��V�8����sgh�s~�	�]h�,�c]�����Jk����խ����/Pؽ%�\�گ��7��/{{��`gOY/S�"���,�dU�>��9�a�h<o�=��fRb�����'�֞�{�Y����j3)�b�X���XGڿ�Lײ�g��CB$�g�>5�G��@�'V&�f�l{����C��H�&U�<m?�#��V	~�Ζf�T��ö�d%�{<a�t���`<��CҨ�n;���tڂhL�
���|Ň��ɓ��ˮ��6S�G�Ae��(e��!�i���Y���ǥ��t�7P��UX���-"��L}h��L���ʔ����
���U��_����yV��+fF�p�wN�58~3��a ��w�$��;�!��&�@�P�~:m"ih&�S��:���[���u�4���u�0���:��^q��5_B�!A�8�H��U�i.FgN<n}D<F��������o��Q���h~�qR�\�*ۼ�>�^��عc6��졛+ԨLH�����dYCg���s03l�^������;�K�@[4�2+I��ʖ��o�O��a��2�Υ�*XR8G/�<>@`�շ��V��!0����֢��ץ�\d�2w7�<�4'B����{��_H�ͱ�P�[Y p�f������ăB(}Ą�P���{�X�y&ce���4��jhu�-I��A��!���.KZ��[q��8�ͩj�(�ɺM�1Fq�j��⟕eN���p���3l�j�Ul�{,��GB��>FlA 	� �EAéA@Khmߣ�Fns��r�o�ErKz�8H��a�`$�׺óΘ�1��������*;B�T&Me�$d�~ט3LG�^���l \X�g6�a��|�=�L`�E�Uc����4I\���O{��Zp[�|�ȓ}:f̍�K����"�����6z�W�n��>'y�<��7���X����_v��A�-�K_!e?b#\��q��,��Sb�9iH�@v����_$�?V��M��Yx�����H��?5D@����hMacy�o�g%2���q�|@�D�V��+�^�y�y�ɐ��ߣ�`L@�?%h4��Ѭi�}���@�;�&z��㠷M�_r�vBa2U���W���9cU5Eʗ?��>@���Q)Q�|�(�'h�	�ƪ�8��tBJj%��Hafwx�����9��y����-�����s#�9�+��݈� 쐰�.��cA�ܐ��(�s��w?�^�ȷ�|�	�>�F1N�sk�3�<x��HCLy��;L)+��!aKX�V�g�hJ|_�X؀��'�L����_�
[�ڧ�4 Y���C}3��a*�ܵ��8��ϛ��J2�� �X�
q�qh�!��3�c*Z]==]�Q��1�ψ��|#��AuAo�d��i�%;K+v�?x��`3VM^)b��0�{��*�w�5�y� ��EC��u���/��䃚��"�����|�;m���EX'i_��wA��z��S�`�@���m���sD��%Ȩr�h��$��!��	���)���q]DQ�Q����7\���}��D��#(�;FK�������k�FvҸ i��(�0��甞#K߻?�&��:���h��_k�e�A~7�ü9�T�v�o�ݥ� ֋N�2������E|;���DIlJ��.0�>?&���´cz���m�_�xGTo�K �f&!�2�+� NsЮ��Zu��M�!�ǳ��d1Zj��ND�u�$/�&�o~��\A���ػ;�ߑ g�߆��rm�H��G$F6Q���]:9���8y�/��f�@�$k{�1 �NF��_���[uY�emɰ߳EC���%�*��~�&��u���6���~����$s�M+h,��>�.���l-���N�{�7������»%��$�/Ua� .)�8ٹ�@����C��zsK&�7�Ws{M�	�i��^��s���K��[��=�
���-�!H_���L�HxӘq��&�ڍ[(U�z���ǅu���k��v�{� �?rQQb�(���S���������!ML	3]{!F���h����w�Q=���I�?�u?6rx���0k79��F�>���pz�|c6]䤶Ր��ӈIف˿��*�p>��E��w<��>�����C��`�B����77#p�!gd�tb"v�3��ݛ����"�9fa�b��o,�W���ހ�`MM��Gtrר�MŠ��_��b����k���J�m@t���T�3�t��>�ǖA���'c�:Gӆ���+δg�U�������3]Q�{�z�Asq�a.�n.~|3ݏ7���Q@��<�#W+2 ����@}��Mrw�9�e��&�F�*|0|��Ή���4L�b�Q���\op�"� �v�\n1����	-�bM���r�s��'����KvT�qN76�a:Sr!^���	�cFr�j�R��N������E�
���h���~#.�F=�!��T����w�>`��f5x�)U}��"o�~z��/+/)5���x0��S0>M�y,��,����� �f3AEF�p�c�d!�㈊�)%]x|\x��w�T��v���'��h����Fdc�)�\�4�][����j����g��f��s�+� ���ѹ�e��UBRL6����o�����ܛ���E,���WZ�L���6RU��"��g:{F�2���'��e���-��v�Bv��1�`�9¹�X�9�W��{Z����S{*�,Dꗍ��r�����~�;�]hyd�L�*����D':��1F�����"���)�3���r�'���8�ٜ�ar�1qf�,�M�I�>d'����I9�ߚ0�$�R<����#DZ�B�*tH��Fڒ��SS;10��Q$/����gE�t�~%�r1�r�،�,�*�&�^ y���J��L̔޶���޴��o�a��˫o,X�G����'_ʼ�gm}|7�1	����I��'kW M$��ۗ�����jb��=	2 ���n�1�D">F�hB��E��[��*1��m��J^j�i���2�~�R}��m=�P��W�e�^4u\���#\Ny�#��d���v�W{�#B���?�E���V*O��Su�Y��3ڨ��6��|?rZ�L3|�[Z��=̅��H��7᳕g�Y/V���P1�K�ͥ԰�.׀��@����u���D1�B�ԊI�^cB��0��tFt�{����.[�X"�;�`.�[!|��4��F��u��ԁC�i@��&@�[����kk��D$CPc��y��:��] ��I�q����.��^˷��9��"Вg.�Y��Îyx�do"��O�2�,� 4z\j皀	)'}�.U]K? {vaC47t|�<
�i��y��Zcљ�F����K��n���(��R�����?T�1GZ�ԑ���&�g��*׿AY��������KTW������JZJW�W���MЉ)����Z�7�d V���@�eI��'��/�z� ��@, Sgu{r��5W>�ވѮ�9Y��I�����f�4�ਅ�,I��AѠ���G�`�j��P��Wծ{-߀�vl�D20aE����m�Vح~պY��1�u���D��y�(?��w%��"��X7z�Վqo���w����`[*��2�¸�hU��rB�#Fݬ�_�k�b��L4!L��0�<E�ӹ�Ϩ��P���g��
5K�"�[�c�->�C���7�7aFTĈ��*A�(<�X���z>��$���:�U;ol����{ܑK���i�����B{*���N<�Ɲ>��9�u] ��9��9H���/;~���#gn���ݢ�]�)d(Ѷ( �ʠ�oo�nA���lR�Z�a���ǑIg��#�H�Μu7-^��|7WL����{���-���/83x��ME�fZ�H�Y���E{Zrq}���2�5.����0&t]9�X�dH��i9�;��j��.����u����"5�5�ݧ;	��ɽ�f�{�_e)�
��D����nx��(�����qk]zS���1��y;�<��5��`N	�3ߗd�ĸT��A
b9��(af�$!7	�ۨ�����ey�t�͙���X�0�|�"^|x�D�!�\��߆�E7���nƎ��4�s�3Iųul#Q�{j�i�ME�Zf�c�qI\�8("�<È����Ș
Z���	�O����V��:�u��W�wnh�>�Ë�8g-E&���Vқ7PW��AO�	xʉ:���m}F�	|�'xS:ߞ�d;5cơ�~����%�T�d�{��Wt?p|�Q���G�B�|����Y,Я�+���VT�|c�k��0K����B��y	s�{V�(��R5��R��ew���D�ɞ7��=�Y�-������L�jj��5^�Y�;�2�HOxģ(������7���ZMux��������P�&����ن,uԃ�֢��$m���)�f����u�Y9��������/\�X`m� ��
Dr�+-�d�\�A 5՗�E����.;.w��c�ӊ�u�@̩?�F'�����k�lQ72@p��`�e�8���Ch$��^�k�d����ڑT�}�ͻ��ңu"�F�M4R4�ûw�U\,��v2F};�E8��o!��@oX^3u`���S,�}:�} >9oz�t��=����g�ǋ9O�=�(�
H��o�S�4��U���Z��U��\��y7��"����^�H��O�:��.ӑ�;��8^��)�u v���������[�>��4�����$��G�>�Z�N5S��n��u}K=}DuBpk��K3%�Q�T��r"މ\Y����?b���Z�f��v����?\�xی��2Waz����W%a����xw��)`��e�/O�z`|�q[5R<��@,r� >=S@��J��ko�'��ܰ�s��VM��B�nm^<��=�×�C�Z�z��ߥ[;ܬ��~�d�t����ڃan��9�TnW��}�a��i5)���z�a��XM�֒�/����X*ۖK�G̚�@(�((���	������i��*���ۑ{�ty��D�M�Ne���\�|}��tJ2$��8���d��޶�k'�I�h�p<�� ����P�]P"�x�/��M�k��QM5�fLd�㟲�9��n�8��E��?��EGZ���w�U���~(��e�.A0p@�!`U��<��K���9��s����].0!'����7�v���c�t��7�d�-|�9a�K�1$.��@���4�&а�O���g��o�)d䓉DB��Is`2z���U�H}]��Ӯ�CP ҆:V��q���#��7��ŗ�Pv��[�s�cQ�֣K�gE9��CSa3-̏8��o��o�ل���fQ3j��U5̵^��PQ�Y(J���m�����VB�G��1�Ŧ=(��a`e��r�>��;b���H��.�㞴�R$޴
�yP���@�SP�b�zQ�^�q�v.���Ȅ,X�&qIJ�J4	e��rJ<D6����&�Z�e���5'��`Ϙ�+�&Iv�!`�z�P(@�3)��4:}�Y��$������J�s!���UJ�|%�Y� ����up^[dz^����nX�_h2L3�����tL���F("����,����&-��i�dx���;�]�T�YJ?@��c�$U�i!-�;�l��)�|�cQ��i�$ΜD`�[���+��	ȇÿ�ap�n$_(�T����<�\���X"ei�Ͷ�h�k�{%u����V�����׺�um�At*��'�V��pN���@{X��̸cLLvXrb쨦�KY�Q{�+`��D�Zk�[�[/��@�AY����,:z�\��Ů}�'s$���� Qx��̬঳��۸���b6�Oq���>?E��MN[������:��,%H�>$��o�L��d~;fJ��N�s���즥mmE��^��x���D��Ξ��~�8F���%�͒����6r>�P�`��o��4��qn��fvca&����}���UKe��u�O���B��`�h�P^��u���q���zBa��C�D�r�J��@af�s��RQuc���TS��=�
��O��1Mm�e��p��F���@��B�Ɏ/\x:��>4L�YBܒ�t;(���D�k��	�qX~%�>bz�8gO��	�E Y&��%q۞����\�@���+����=���8AZ?�ޝ8w�M(�8RB;�_g�3-M�=4pJ�%ᏭC�ը!/�+��)����A�6�������
��A���*æ��320�k�0�.��3�W��jn�s,ˏm�L�%e��I�M7�g���¸�]ޟ`�470�T3���+S�\x��(� �/+7��ƕ��<�����]���B�:M������C����X�jo���
}�Z������k�$n%MF�9�T�P��B{$<�$~_������VA��?gdI�i��gO�[���R^��S40����e�߼�/C&S���O@INTڽU�Q�E��Z��(��j-ǃ� b
؟���pۭ>'1�e1-7|��dZTީ/���v�`��oޠ�,�4�,(N�� �@@�zO �����ZEa�r�{�{B�js�5��0�j���'�i��4�ΎU��@�+}���Mq�.y2ǈ��#f�^�R\Bf�%����z�V�i�G��I�Q�YNskT(��Q���a��00�B��-�if�Ԋ��X�-��Е�Z��JQz�����+����׍Zo!)WC�����~Q�h�bﳼ���b���(�F��hJ���q`j�̗2$�H�q���2\@L��˲�R�3R�Z@t(��,?��N��w��<���x��B+[2kt�4k��k��Je��Vm

B)��匹���q�\�C�[��=�H�w���u~�
z�+���榶
���7��J�پ'R��O�5~�|ZJ������}tF�������l�����G�������ł��; ���^��_$$��/��I׻� �#0�H�=����t��]����4�jL &���z=;���n��l�Hb�d����� �r�!v�g{$��A��UI���:!�/l��fq&4d��M�����J�vD���5�՛'� Nk#��25�"�2����"7����i�m��Z!6�8/��Q��s��?���>�w��g���Z�*�I��\��
Qb̬T��J����a� zH�m���4B��ΐ��Ib쥅u�&N��:��EK"/8F��H��r@��a��~%c�Yv����s��b����l���m]����K,�7i�j� �N��D�*����L�h�3���Dr���fF���a��b�k�wL�XN���s3�g����=k[���Vc�"1k�u�#��ǔ|Zߡ�W�]2�n� ��������>D��!�� ���6כ����bC�W7hQ_/��;����wC��O�~y���O�^11XZf$A=X=C��L�ˡX�չ��n�/��i[B	�v�K	Ն��&�3�Z�Δ�w�;�hI�c�RKe�⭻�rek��M�W�7=6R�i$C��ܻ�^Řʙ+Ut �.#$�v�P����ٜ_�8���ʖrIAI4���-�Uq$��3i�[z[��{�%Ej�S���r��u&���p�YI��E�[Ud	V%@ްڃ�۫A!R�2�	���?g��\�	�A0(�Z��Wʑ1s.���hH:���e	f@C�sMH�1��ʹysݽ�}��; �s�ɦ]e������h��xF�e��D2��[�o�w�ǟ[�98��w��)R�4ah�P�	�?��p�i-��~@���z)�SF}'~bNь�W�X�6�#��Q�+��`�<_�(l�m�x��OF6u4,u-&�	槑qe#)x]���Y#E�Z'z�VTu��(S�͉ :~��0���BB��VB"�f���I�P��|z [�����ƛ[�{p�)����a[��3mnM{�7 dB��S>��	��yR����mB<Bד��h�Ӧ�9����C��A����.����7���-���Z�闊M�G�"��e5����	F�6t;�W[�F���̵��v�~���Cp����`����(��B�i�Ny%�~�ȏ_�qY�b~�]f]U^A�8a
'<�+�ܰ�u�ܧ��9�!J�\������[����+D�V ɩ{�]"bĈ+;y���^�W$Q�m�f�.G�����c������(�?�7�G��`��ύ`����#��<���-/��}���X�9�ǌ�S��Z�t_��I������8��s�ZF���PVB$6��Z��֚?�,ؑȳn�kky�#����;
Hrr���t�q���g@��(��X���q�a+eX�);1��0ߵz��"r>|�U�F��FR���i��T ѳJl�<X?�e�x0c� � �ߍ]�$6 ���'T�N(���Ɋ�X�^�s�j����	UP��8�ctg�������s�0�)�%�E�8��4W0
�а��AYK�=Ϟ$�l�_r��vh�&'F\�������m݁ �'�M���I.��z�6�ݮ��+�\��.}�	(�LU�+t�~{���W��S�M�M*F.���:e�5\U�6��a��Ȏ;gdo��#O��|C��`f�@5k��\�0n	i�.7Pw/���><|��>:��Ϗ�H�?+�=��-� �0Up�n̹N�բLH�6{�h�>��@^I��s�h�x���;����O�(��Ǚ���umv�^�����׋*lj�>�i]���_�kv�ޜ(Vc�������fv�y��'�Y�ll�fb�I*�1�?+\� ��[��ل���[�U�����@|�I���$���M�:1�(\ӷib(q7��74S��/Cݷ1�^tV/���-8�� �&���C2�������c �8��Z��_�5?k[>DVvM�-�lŞvou�t}�d��[��}s:�ϑ{W�Q�3mƕ��㼑-��_�&s6��"��6�4�-���Wv�$���M����=U�0���.����u'��ʑB���c�Y��}jkw~���5+�
���l��̻Z�1�� ��0?���J) ���`�'�N3��P
�wa���d��ٸ��?{�FF����+��Bk��ũ��ړ�Cd�<�:��9nT�h\���X6.IaԪ
�X�D;İ\���Z-���Ux����u����UR�����g0A]�^|���M��	�k�����.�ubg\O<dR��|d55CMS�$����ƙm����*�n�������V�AQz c��Zl��Y�4�?8�����6Q�r�˘�C3B�_;�;���K�,���(\VT���9]
�~���Y�0�	w�RљiU���|$���]�M�I~c\݈�
�p���$e�U�n j��(���� �򽌎2%	���`�u���'��1����,h���Z��Y��X�&�@Ӧ:�����Wu���:�0�Z]���}���/�P�1��Jc|_1�&9o~�V`(�K��Q�̐���J~K$Y�Mh�Z����"J�����co�=:=���}��*��o:�|���+?�R ?*��ȋ�I&K��˷�WAU(}Ė���5�\�0P�)�W�#k���y�����Y��c�_�"�0�~�����ei)b\ ��g���"����֑��`�l�5�Q&�L����{����|F�F���F}y���=��rSg��k�ʹ%[���\����ӿ Y�gr׀9�R�L�a?�ɴ}C�Z�l	�"������q%��;���pj�e�/�	'�:;x꠳�k����g}Q�o�5��L�6x))���hQyd����R��X���p�X����.d�,��x(7��GV��"�P#��3���k=�1Q������[�k�z����!�l� ���D߃�����]�f-B��n�*��yYU��$�5WC��<�3����?0�~"��4Е�y�(!�yF���_�L��Ufػ��&jy/�L�q�9LVK����jL�߻�u_��C��ĶE�e�as7!�G�x�@�%���
�d�E,٬uKh���.�sϲ��i�{�X��zվ�'�I	��i���Iw����g���n}�Ç^x��
������&M*�BX�!�5z�>��(A�`NϪc���Ťy2�C�.S���� a�z�;B4�Շֈ�{t#t4-��%����g���D�ZĊx�ULc�!(�Ey���} | ���%��.W��_&�Ϗ��=�����&)v�r[�ɝ�7�yQ��$����
>[ݬ�*�ț�쉅���;â�1��/���I��riV�X^_�����7�<}��~mH�[��N^3���P��sٰ��J�4��b֜$�9tO���C����0�����~��N+������C��2�_JW�@� -�1=� �K�9���D�	5WhxuJ
#�y���A�����f�aM�$y����Y����47�/y��t��?U�a+e�͡��I�U���2(m;�hlD�$��Z�0H��9Y�5͝�%�%�ߤ%Տ��m��u���������^`y!��V/�\�~DP�W�,n\�ϴ�f��fb4���'ڕmk4q��,��֗�g`,�Wh��ϰf�C����47c��6S.￵�yq�A�,xkb�ĕ��1��BB�����V~[jP�d�W���}�B)׹Po��+�l,�ReI�R��nð�,@.j_�Z^��Έ�ƚ�����픅0G2��ݦ��oE�iw&H����
s����ӣ�/�)����SB����1����#
��f���]Y��nf�3X�W5�8�8��n�T�-%�w�s�mC~ym]=�<�j˼��k:.v�l���f��(&S'H�+���j�)�<���V���Ε;�7�[��t�e���zr5Y*�<�� h��-����>���:5S��#��SZlu�-�S����ܗ:V!�p��_0��ìrW{�:�� ��,~$��XV����YI¨|�v�E��P��煲�L]ll#���� >i9�u��rQ�����5?�ˑ�Q�n0Y�{:��4��T��m�m�t2�X�5�Q6���,3��M�DU�:)�Ҵ�G�=1&�5�b��:�	_yصg��q���~�Z�� C���{�
x~������$r�ď��N�K��!y�~a���Q��M f�2������r6�qP�U=# �8�ԍӂ��8���|����u�`k4��	�m*��5��,��)iL����$8��Na�l�:�����X���������.����qH��*��+<�>p��B����d�}H��Ɖf��U���u��C�h�� 1�u��!jT��ƶ�߯�G��������0!n7�Ӧ�V�~0H��g�u�a��}4;���R�W�h�P� ���,~��u6Ĭ7��#j����w���(��C�Li���u��b�+���4�-��O�m��ltܯ�c'�"��o#���2e�-�@����t�9������� KS�[�w-��4���O�0#�ਜ਼,9�U��i2S\a-g�$j;2�s�%CY�m�(K�
Q�=L���� I�Q$��86J�nų�	���G�+� a���tbr*���W���*��.!4:�{\�*����h��5�����]���P}�xwښ�_�ci��{�,����\���BaK&?�!�=frl���C�Uu��xv:�9�
���Y�� �0�o���B�K]�[�R�>c�����]dTO�'��Ց�"�3���\�ގ��O,dn�^��YB;��|�O�I�w�6'9�A(ZY9��t��6�T�j��/����s�����i%�����|\cuG)_R��ʇ���`7��gS`�D���N����Ѱk"1�2�`i��L>y�x�J�qp:3��q��� c]H�VL8/��&��s{�]�f�3�_��$�V%��[�ڕR��=>_=�+[ �C��Nm	]E'���J�"��5Yi^j=5E	��&�!��C.��f��D������^�=&��<�����i1�]n�l��Ws��n4�
��Ź��/�l���K�Bj0;G��|�r��̠�T����qc1��?��u�JpeX/v� Gz�H�lkH�<���]K�p�����N�3m/�bl0ȯ�_ҕ/i��{-��[{28V������2��?�os�b7y�c��Zh>���l�}�G���3�������gZ"����xo.2�������9�3`n���m��R��m|�y���'绞�v��!�;*=�F�?��k��!�8[�;� N����0W�;Pt��<9;�
��9`�1�{�e;,�S�EE&b������'��~�+�u��:�̵B[m%"�c�S��0������1�����ْG,�h�YQ���U�M���<�ퟏ܁T��Qp�����Z�&���}Hy�)*MH�4�����I��%̦"�k�����X	���ސ_vD9+�� ��}����CixF�Q�HH_*��c�1�&XI�q\I���^,W_pY�R�)~�s��cD�]|��p�3dl�S��CG�y7���u�|�͞*C���W|��k�=lv�
���Ѧm�a,� �{��&q,��j����>���Ճ�4m �1b�q��F����a/�Ef��T`��L�/zD\�����G�|R��d���|�}+����H{�Br[��˲S,]�+	U���̏��}$�)�>7o���6z<4�A'D��a��uA��vG�qF��K2,��v���?�I?U�.���G�ֽ�ȃ8��
ړ�(�|���$A]״�X0��:�:��7!2'6d��.���A��Uj�k3��o�uʆ�F�@i�8�Cŭ@�=�_𛓘�j��\j��n�y�<��3�P�v��#�����#m8-~!�6���MfC���Ú��&޵ ���z� S|��u�g�������r����J���"L���b카86����]Y��)�X���w/͸�9�Q�2�p�E+�P��_�
�c��
�dț�����|*y�6	?�gn%S�dP�ݣ$�<�6疑��\��g�J6`��B��V�Er�J�~����#Z��˲��Yn����$�gRPtj˪d��{�N�/9c�VW�oד| N�5�*r����N?�qX
��x^�1T���Үɦ�v� Rۣ]���6P�8��:/{�a�wn��	���W����ύ�, \nh��Yj�F>ʸ�yc0ds��M�N�(��oqhWa������qiKrZ�G�&q����-��B�k+q���۬��Xf�{�ۏ�O�G�]VF;��U����A��]b�g��]����iY[R8N�� ��:"��e&�dd�C��4�Y1A[�U0�����)�_#��,��g�E���E���X��a^��o4��:��-d4�
\BKk)�����~X��_2CI�����G>�:� ����&T�z5y��C�l>e�����Z�<f��ՕH��-�֨74�`��]�[�2wM:�P���z#/?~M8�� ��0¡���O�>�P ����F�L�SpV5/T��tF�о���D,��B=�F��ܟ�B�����~�����4G��r�K���N^����T/��H8���v�NƓ�q`5 ��c�ʞ���}���W���%;D���+.z})��JjhQ�Pn����I��n��`�c�z�i���.�-�"$d �ɟe*��Y����錱���y#��e~�
�ߞHO#�&;l"@���|?х��+:�;%k���M"P+�f(Ӆ�� ǥ���K�0��}t�㓷p~5�c�Bɡ��;a���-�+5{����\�й�`�.�J��I��gA3��{� %�����]Y���RQ$>m��q8�x���A@�����Y����rT��Έl���.T��� n�a�_nE�.��J���{��KVC��xRI���E�p�fd���%����EhEQ.s4K	Y��st^E���,�y��Ԝ��N�Lܫ�F�&J�(�#pR�ܗb�O�@�f����4���*^B�k����v�W�C�[)��G�MS��ɀ��K\^d��H���Bd@�Z�/�=��}��5+�~'΀Al���1��<ׂJ`�o��3*��J���!��a�E�>�z ��K�a.%��:�W�h{>����!u���m�����!�Y���Y�|3;�]�$�pjbz�c�'LX�#�"=.��j�R�~��ެ3�NܥX�6��?����"Oe��������#�Z�*���?���`� ���x��i=?�ܳP�4��B9k�l��$�����R �H�[e"�ǁۡ��Zs���<��|h�*���Ŀ\"���#�����&�Oڽ�~����#C��z(���?g]HO3H-��֗�iB��c��7	���墒7X�ȿ.`�$l�j��70��fɃ��� Q�ѿ!���[��<�M���b�p|��#
A�V3Q
BM� 9�t�8S�(�i/�-.m�#/�!QnYV`v
Jd�A��:2r-�2��>�|;�\N�?�Q9�3�&�N����`�KQP��Wc ���b� ��z�l?a�����W��p�1��nɞ�#n������oG���a��/���X?���5����f��Y���2o�esZ�+y��(�%�}�1����4s�i�@.?���P�)
l�~�
+=9���@Qn.I��N�e<K�C�=�c����o�n����Gל�G��v�^����]��Q�^�%�b�O:�O���[�	fΞc����L���^�L�j�_h�:�������6]��PG�"�8
 c?4v�2|,�+C0��C���u�l�T�d"��).�̞V��U�Y^�Ub�^8��`�1���LL���~Ј����^��CQ�m>��=�Z"��h&J�Yh&0�çv��3�v%d��f��:]�&cF|���+�fa!Xp��
9?�z�O9��&
Qdͪ�}��?>�愈$�y��'o��\M�?�|%�Mh��M��S�@�z����y��BK9�CE+3P��kj94a,N/ו&'2�/h�%�I��om��j{ł�Z!^�A�̺���a� /�C0L+��p����֯������7O�-�*LA��'W�9��o�:�YF����w��K{�|Q��3����"�+�"�Ծ��3<*�?�F��)H�ҿk��0����t2�C�?�����&.N1~���e�|Α���gL=P/����M=���v�:7:<$�Yb���