��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���^���IѼ�E{g{�^�����w*��0�%«�W�sXw�
sg,)o>�u���z6ۉ_���y̌�G�UD�R��:P�3]mx��.�:�=�$�x1y�Q��m��S�"�5Ղ�L�J.��@��� ����|�Q@������k��kk�=*�o"�?���=����I�����N��+�R �hD ̠���1�0�������g��֖�)�HM���B����و��_�m�+C���t�Ҟ=�T�p�nhr��Ħf�;��F<�F0*g�c�h�N���df��eۅ�l�SYy!A�E�d0�;�:��W����� V�i)���:P�\�=PHOF�R|�<�}I��2�?@�m`����f�82����|�,��7Q��oS�uݦ�1��>��9_(w����t�_���Ԙr��/�Y{>�kݺ�@�g3����Ʉ��Y��A�ێ	r�:e��2�����{��^��iWb;~�'�E������r%��̑t'XW�|��L�x�q�O!2���%~��[�bh�Ja����BkaN�G.L;w���/��J	57�l�h��r���y��-KW�<�p�n(a�!���[�4����#Ն-S�NÂ��u�m@�*�5Ke���`�����5����x�Z� K��s	��J�����p�Ӵ����
���;�aS��y�J�����C/N�XN�$����3*���>P����M@X��I��&�����e췰��,=�M�u� ��6�I�N���N�ԝ~���2�L<wY������?��ᄇ�����rH��<�7��h�Z��ƙ16�H�\Z��M�0���f��-�<Ffٷ��F�[����[αM��,���(�����;`��`=��YQ�/�ۃ)�)�]l�����M����V&!#D͸!l���L6��K[�q����2��;�z�$�f1P>ٕ6���9�IR���o5�HW�� ���E{Ǝ4��<�S�f��&.���������Κ��TM��?O� wwC(Ê�s�fW�����Fi�~@�U�o�)_L.e����;�S���;��O����~���ca���t���f_�и��-��f�60�Do����u��?��^�Ա_d��v(�0j}��B�����B��??��|i4CU�i3|p������Q��-@K�/9���϶��e~0 �����avP����5���M�p[}���&�b���ԡN�cM�Zs������Y�`���G �`��@�cw�����������ݔ�.�$��@�v�T,q�/�%%���3�0!ߝ0ԁdUG/P�IHU���V�8��9-���~��*և���O��y/Zw #�wI߹W���g���\L�z3~��pa�Z/�Z�O�TM�w,��j$�#��Y�[���I?�LuP�ںيа^�6�񌐚2����ե�Ⱥ5ؿ=� ��L۲\��,�C��0��h�&t%�y�����L4��R9��9���MZA���y՞�Y�P$�t����&V����3��k�ľ�Vd���L��V���AR7��,pA�K�qRt+���y�mg����^�$<�=N�8�ݹ��[G�fMpwpռ�J���2����G�rgάv��5Ub��ほ���߭�n��ťӁ�ݺg��i�`���N��o!���J+c� �6Kd�s�!&�*9�UD�%-�ή�/'J�3�b��0cZXuXp;�{�˰� PM�� ��7⽿�S�C�hi��elo�tl8����W�U�2�6�\̊+B��I��L�F�Y8s~T���ټ@��W��g�^��?���D���8 ����Eʮ��t��K�v�FLt&�@�W�i��8�Ӧ�5j�5�2�,��[����@3*Q�m\ڡ���M�k�l�=Y������ǲ�|��X�UQ�y�V=��՝2�%���� 4fBs	9�s�'0i�݆LG-��p��q��ن���6��P�-��b:�BN����24Q��eW �OyIH�V6���&1������#[	�$Ԗ���S$fp6~ˍ�T�B3�W�k>��d�^k���R"^˘(��7D������i�Dq�V(2�����j�:�~��@�g�2�V"cWp��5>���_��q��͊�BJ^���Y�+�e�ڧ�3�mr�M�^bj��o����~ ��� ��0��2B�@��[���[E�<���čt�Sy�ha����q@�k��;����l��8�_��O?X��{�����9t��� �ީ��Շ�R(.�hE��}�S�R�~���4��,璏�R��s���5U �]ׂ�=�[0a-(1\���͹�N��?!�.[��}bg6��؟*��W��� e���|�n<�+r�M�x��(n<�7�Ĩ,�3�$|.S3� 2��>+���A�H�_#v�[�g�hE|�n�����<5����	mG�"TeJA���=n�Q)��ѿl(�
 ����]^b9��l-�
F�����ح���RJ��G�t���У.�\�z�{����ƯC�UfJ	]��c�[V�I�����n$�S*Q*��Cka�Τ�����v\�W�������j�0)g��MVF;�Ϳ���V�7��B�NAuT��q1��H�'}�\����:��*ҹӵpWfճ���E���lh���L�xFU7a�y�0r)�E��=x� E f��d�`���\
*�.���,��-�A*�;i��Z�(S�Ɔ�ǉRD�J��OX��A
Β |vX���u�B���z���G���-J7�6h;�����D�S��n���I���\T�¦�+�\�S����1\��_����54?�h����r9|�<-L������ޚܫ�^�7|)�f �-�I
�QX��6A�<;�i�>^��E�u��҄&w��
@o�������@�U�ul��4FFIh�tY�����u_�1"-��%B�/�_��-6�R@�_����&,��ʙdg}74�#�"k�a��,�
�3R�"wO-��n���Ã�аQ��~,��ū�xi }�p�� w�!���8�H�(������!TP?�!� ֛��w|eμ��CO"�&v�O�6��K���0,�X����p�S-�d��y[���}�q'|�o�4�o)ϙ�D:]q�#ӻaln���6?�C������Yk��	>�7~�����E}W�k��n��=7Ɓg#$�;)�|�Ȭ�$ޭ�b�۴l�p��b����d�?j�n�.��kw�I�cf%���܋6��nh��Yj�(���E�pc�}k�] ��6��[g�3Y.�ўʖ~��I��߻>�;sy�%�C�]C��W߸k�^����V�;�ÑN�ֱ�9���f:�T���!�~O2���5f'�SN��7@�>i�b҂��]N!���MK?��"���c�������������
���f�T,R����ɒ+K�V���J%�PWRm�R�s�͈3H@睎�jH�[���8�£k�@� ����ğ���W�JV ��Фtd��d'v	�E��Ur�=ųƾp�=�mW��I�[~�C��/�l�ƥ�$�R�s���^BI�yi�M+;ݴ�b��F؊�czB}���rt�p��mZ�'�'��{n���#�@~}�(ۀP��hZn� ucz�~=E��0UP�?�$�� ��Ʒ'��	!hu��ܠ���@��&�Qf@�D�����G��A?���K(T�� $H�EY]o@³�[?���s��G�h��S�D����Y,��6���:��/�(h�1�B3=.�-i���n -�z�?.�F�b=��T����b.�gv9���f��cu�M�]ڤ����̻YMTam���B�GtI��RW�U�,�j��B���g��{���j��)��G��j��%O��H:CY���W�  �Z~�4�������`�m��+ȑ 2C�#%�1d�1�%�A�ʌ�%�
�r@�Y"��Ê�#�UW�G��x���erS��#��bf��f{�w���_u8���pV���#�n��H�� � ���Y�kM^��|�=���g�P,�C"�^��\se�Q�#JѪ`,"��{�~��ŶX]��PP/��dt>2tK��ہ`���^x�/�6��e'�T��3\�]{.�3��UJE����[���p����}�|2.�*����'��q{���ߛr9�0�W���l�����Py.A��<�p�Ԡ]� 4PS�=����jݚ��7���/{+��>^�P��Б[ҜE��*��+����$��M5�#e �@!��7�?tg�kA�r{��gvQ�*c�� ���"D�����%@�]6��YV���[-��)��u<���_G�So�]R�#V�pn���=�[�p��=��; ����p���-�0�!�ѡ�K���ϩ��p��s���w�k�6�L�I��������m$B���,�l�H�s�lǹ��h�4�Q
���Wg�����{A��0�'kg�ޜ�]��f@Ǧ)�����!�ãaa������% th��rǤ8!�}N��������"9j���^`�-eކ��P�RG��1eܩ�o�m�H�ѐ���pf� ~�*������v���LU��X�L/܁��߇:��o9�������Z�d�͇p���#
4c��:ﶖ��:��2ͦT;�	���M�v��+�9�^�0Z�ܳ�䓎e�	�5C\�S"��	�]a����/���9N�o�<����0T$$1��s�g��IvJ���d-�"3}�w�Ě^�E7B[��3t�='
�q`-R�R�S�����'��ɽ"�ϊ��뚔�Cƕ6r�{�duh�4�CBf(',����o�����-H�X�1�]���Ba]���w��(������������7t�+�ϼR���[k8}l�w�"�rDލ.Z�۲J��)��!(�\��T�wIh��7�<��TJN=z�����:�L��t���{j�5��.7��C�Qm��#��5�>��G�2t�٣�2ǇŠ� �����՝�4M�#��q��Kdo�b��z� �*]�Pl~�����r�@F�b�ڋ"�͡���6w(��Z�-���}pӄ&Z�Y���yimZ����'K��f�b��2�U�.���s�4��a@�ȸm�`ȈB����h�elDI��y7��I}O�e��0V��R����{`E�r��C#��.w[�� !�9��t��_^���ᰡ��m����5f���җ�����ZwL)��C1qC��uyf<���몍wj��BⲻOB4���R�ӌNHY�����8dQ�_nxZ^�/4�R�s��G��MC�!!ӌVh����C����#5��f����9=��Q�p9b�W~퍥�/?*=�����#��
�D�o��ݿQc��i�w��f�~�ۆ�	a�Q���QX��!8[�[��\�X� @�^{�j,A1�([�6�zd�.�o�՚I�%ld̎�!�!�.<������?ʸ��,��'.>as���Ǣ������-D~��.nv p$�����U���Z��*Gmq����!�W �U9����X���$Vt�5^�`�F+���(����>�
�>	@ܱ�&��t$�:T�]R�3'�-V8�Z�P��%��J��-�QtF�I1MV�{Q�����ΰk1	�nƄCo߯V曹�QV�f�3;�������Z\NgC�+���P�U�zG��*%�2=��'�2����&��	���ʟYl"�0j<K�Kxp�h�<�A� C�����H��OOk$����~���2�<�!�`�ͪ�ܭ��`.�V�`]��\�+�)���>i;V,��"��#�N�Q/@K�^�6����$�޻������٤[���
��c�6�h�<�]�9�ǁ� J����d �(kv�՚��t�Zo��7��T��N�����|֥�* �'�!IW�TX3���-^-"�;������6�	��hF��bN���X�R�v��<�;�zL�U2�bܩ9k�)mۺ=~
%�(�dD��Ƀ��<1H�������K��R"�_o�p_����F��A���K�c���*�I������L��O8�`	lJJ���u�H�lb;� ���7o�~r��T+��Ѿ.����x����z5�"̐Dч��V�+03�ɏ�i�@��m��3�kM��;?8�t�Ȕ�I�:'T!�&�<�-��ԝ��`��g�͇֯!+W�����Yv'���c\27)H�� )���J�6�G����۽��}L�ƴ26:����{�8ּ�-؆��9� 4�����4�m#q��'��'� tPqOY��K�+�OۚZ��w�%2e���[��@�ވ�h�e'�v�����x�H�0��.N/c}e����_�Q�L�D�%'QZd����&�6�{p��h;��	��B�$�����5�YO����=�g�݅�*�d'�ՆN>���f)J[�w��/[�T�u3�O�]���AŸm*�@�V[C�b
�l�4���$��b�A2*3G�a�7
�Z���U����K��B��Mh��^�'&���,[D[�T�'��<ΩEc��h����pR��=s?�1�N=o��`�HVSd��5L�����˵Ǥ����"�H']�O`_/Y� �VƠ%���i��*0Qt��HڀY4���=��-m���,�(�rCi͜o�� ������P'�3��m��T1�C���u� ;�$}��_n6o�tRzxi�.I)�D�?��+�w�<�y��:2�S��|D�i1���� �o��u��[�0%]���7��z�i%^V �'��X��?�X/i�ˑt/��g�%��Ҋ�C�I	�n���}G������Q-�Q?׏��������y�~@X�;Κ+� e���ϩ���=:�5���W�Iq�Os�E��g�k�iSۨ@O���o�=��|�w#���C3>gr~�~�I�[���B����N�8�&�;%��s�/6�*'~���L���Ѱw Qhpr^_�F�	�t���o�$��mE��BC�>���q���1sb��Eo����b����0��_M�I���FYNa�����G�j��D�i������KwDU�lc�:%��B�����	��
:݌C~�r�o��/�T�(a���:�}s�:]NR~�dN�Jq�hl)i�5"��1J�{Nb	�w�&�̪����N�c'_�'f��ii[��i�Q�d��<l���+�cT+��c���s	j���6�q��12~�*�� c_u�G��*#��a9o�"���X�Ht�kq�W���;�v���ŅxF�'�$��@�~�Wd����=2�hq�3<����1��{�sJ��Ka�JE��ibi�}�-��7A��6��R���������n��\�? ��Øj{T1X;²�8�z�E%`�zo����9�����'��ڕ�i(�`���U'ձ��F*�����EK1����\�-
�a_�����5AL��6�b�q�� g�k���>�8w+?��y�9Bs~^R�Y���'$�`��idq�-h!.���d��0��ӂF=W�ͽ3�tG;Z�3=Vr"!d�����Oڏ��ʓJ�i�?7&Hr��o�4�o����}3R��[E�i
	c�^G�[�n1��s&4��AN�2���ܺ�8���E�i_����y�"�]���j'�̎W��2��ٸ�����
�'f҇�\��^AO�9��V��G���q�3i�g!��ʢYU����/�$�i��'v7���G��_"�8����)�ϡ�(�&�'�r �A��-�R�q���N�4U�K#x���y���@씒ru��Z����t}Zz
�&7��}�����y�^Z4I9#���T	����J}�Y^h��d�Z�~�[G��T1Ж���y���� ̌�!�/�����,���%~��[��ZH�L��#�N�}�O_�s瞬&��f��-�u_��H�97]�)&Z���òd'�ObT5�EcȄ7;��7�c�D[��j�|��N5���_���z2&�����{n�Q���ĞB�lT�kqݬM��/�ti+�c�$���nC���u�Gȹ鲞��a2�:�����Vm�4\����2��v�?]����.�����~�m-ʲf�Ӵ�����&t���?���@`�O�p3Wq��Fl�Kh� ?�S�2:���̴�������u7|��<����!�	�UxY�8OA䄘q����+^�Pr4��e8�$H�'��}"I,B�s8��C���d�Lg5�d��D�hλD!�D��^�K���|�uH=M�ANbQ��k{�XT���zGC
Z�]�.�����7��5�y�"��)�Ke�L66�l#Uo�������,$��~*�ģN������K=�?���=PO&_��,�t���b�x�БC�����Pd;e��׷<�ݍi��q~�Mo̡��p$%]���L7C�[��+9u`��.DCWyT.[���30i]z<�݆g��Ox��:~�巃3ɣ��p6���f9���5�M���@�
"Ħ~'ߘ�Y8+0[�tI�%�Z�N��Hޢ��.B2ڕfY�m2����~PM�َ{z��k ����l���_�L4�*bg��]21�EkK�K\���D9ue�T��3��a��҄}8&��6L��z��'���C�]M��ꨰ?u�R^����V�������ҽ5T��&؜��B�C��1ݷی}���=\�=2K��Q>�-��Cc��$,�Q�X����W=&������9�� N�Tק�O%@n&`ȰM��t�PG�dI��_�'=)�R,[����Qt?�V�'��f��� /T�L�Dk �B�]���~梊�:t��OI�0��|C�u�n�0u;��Z���T�By�^1��Gzsy-�r!��l؆#��Z�8��C.����db�VS3׻N" չ$&ސ@|K�x/�aM��:�)�|B�\s����������~�*�R�T��z�j1r���x���˸�4�s�,�@� �Ls�F�~�M>Í2���s!�=���W��?��S�"nR��
b��D�;��J"�$W�a���dy?U3��Q�k|a�lxb<;�8�l��<�3`Q���l(FC�E�Nu���1\t�P�@,�*uJ�jL��K��'u���rg�RފF2.��U������'�C��]s�I�������<���!�p���P���-l3�	Q�^_L���1��?"c�5i����~�:BA|�J(uC�D��Ȅ��k����i���
7��M�ÕJ}k#����L��7O��'�#ah5����Py|�fJ�⭎a�O��[�}�vR��/?a��Ҵ��{D�?[X=C�O�~�5.>l�e�D�b��Wo>�y��*�Z/�%����'D\�>Q<�;�3W�g��s��
)�c_zY�Z�-5�7�����rU��{Z/1+4*�Z����,)��\��t�*�v�Id���=�¥��ڶػtG1s��ݭD�J��BG@xZ6B6\8$s�{����ʞ��-[dU�8��	��"ۄ3�K���o���|S[�6~���U�xP��NkAjy���?���b��H�1�U��os�c;H�PU�.^�Z�bҁl%b��P��}�Z��m���Y�rW���� ��z>.�q��'HIϚ[��m��:���d���·B�U%�9�����G>���h�^!��/X�_C�OŷI�:#^��� ��1K�\�%��������6Jq�ʯ��n�%`$�i�qM~����&��f�Gm�,����4�abNQ�p͚#��c)��4�B(f�8��m�Ssh��ǚ�8Z��KüQ���Jцn��Pc���קeX�|`W��!�7�6��W��׮!"����v�W�FP��^��Q�6��<��\��ǀ,��}m-ygX!D3�� ����5+����L�7*��7���M<}\Tv���sQѥ�Zq��R�2��?Cy%�kyk�@=�Q�\�����Yu%�����O�Ӭ2��s�˸	�F�L߼����5g4tb����q;�Y�Ѷ�1߯�H�������|��~�pS亃�TL� a}��Z!;�E�Ч/�^R�����!�"��tS��k����5��)?���%V8жe��/���>P���*�O������Oh�'b�T�[���4�ѱ��)O�C<�O\>���)����b�|��k'l���|���K:��񲻻Ǧ�:H�=�$e<4@5�i�+^���v�:��.: ����w1������M&�5�(�}i�"���Ϛ
��������k,T�	W�%J������)�9v�;:mz�:��2����8?��6Ӽbҥ�����l9c�� �X ��y��}����9�w�=��σ� ����g���`�n 
�!����* Ĳ����>.��o�����W*{M;F9����z���=�D��� S�.'�����~�-��Fq�Д�f�)+�GktKN�9���&?p)�R;�>�X6P�ɭP߭��2e7���hf*�Ԥ��d��-��l7��������H�M���c7U`#��Q���Tp�yU�G.�8�\���Q�n�p��+%ǯ&��N�ڑϻ:*�;���X��"uvb]�t�>%0�������?@���Y�N���X�i�ޥ6`s'�<�8�����[f8����̉8�����@�PN����)�|�?��?1J�fw)T��J��ˆ�ɘOX�*��l h��ц3���h�"�b�J����	���<�w%�|A�O�";� N-ZA�����Mq�/�x�d�O��^+$�|u�g\2-h�ګp�7��D��eLT��6ST�a�"��Y�f�;�"ow���k�t1W����<E�*�y��$���oO��Nsr4t�`5�t],�vߐ�^�Z�b�	�d���6@~F� 6Z!�z�`�� /e��,��8KPH0�wۘ�!�m.�z�G�8z���gƻ�B������%6R̨V�r'4�g�Ȗ���ʏ��>�P�B�L���M�e t�~y��{N�[_���(�Y;����?��d��n����U��%&�z���eӭ�v38i(V��"`�L��a'���)�h۫�ݘ���d��q��hN�R0.ĩ�5�H�,�����7����r��b�_��\�ӣ!�!���L����� s�u�$&^-�z�bh�4�G���e��GT����ǿ��gq�����s�%�T��}Ŷ)y͸	,�x��M���j�K[��)��(�6}��&�Z_m��W�߫�Jk�4��*=b�Er�n+r(ڙW@qt������39<\@�;�*����I�Y�j�:ە�]qo?i��-8�g����0	�Dy���S��Wtl�G%�����Jw���C;�%<�~2'fC�a�C�WϮZ�jꈛR�W�����O�^��h@�eEL N������؄Ne7V�I�D&�	����[���M֨�m��q�����B���.�#�[�q��P�wN��yZ#�"����x43edN��q}Ad!k�ic����_�ҍ����/<��6$���e)�U�O�L�/g���C��dZ4z�)��r}�X���'��t f�d���wmvUn&�<�ܯT�r�s�{`hDe��J�d܎S�c[��w�N�>�h�E���`� Ca	E*Nw28R�J�Q�2��������� H�EcQ�2w.��\����2��_�f2���ɀ���Y����w"��#(��F����S��Tuz�L���"jW�؉��=���/(���T���3�x��� d��g���㩀<�f_;�$N�Y��-�Um�`(zG�y�!Id�����\f���Q�R�̬�t�(bxd������@MK���EAbHQ�Z�q���צ�b��O�P���G�l�H�����Ժ	͘���rB����pk���ם/�#&_��F���:�U���c-���j[���),�ͫ�Q�A.D���C-]����L�ޠ���_�@���t29VNA��&ꉾ�o�)N�e3���ڮ�)�뱟��Ý��W�sTbtМɺ�"�RAf�'?�H��*��5H�]Tj�|d��C|L%��M��|�1 �Z@	�IE'��0xͨ$�1ߞ�5u��l��U��r��[+�!�5���k]���Ո��F*/BL��v6�zB�?�'�-�6�jI)3�V6.OI����G�x�I����$6�<I�͡�F�N^~Y��S&$��ne���.q�Mi�"��`n���(c��3���NF�Gts�r�����Z'��9_��f`N�hG��c�L���6G�^��q"���M@v�c���]+����2H4�ֻ!�L����R�_JL�S���c�h��+�� >��4x��2��zB��b�:ޔd���������u#�:����F�H�u�I��3�֐��e�O��$i�6���&�����r��0}n<�$���kt��Fp�q5�RL.v����4�G%s�2:����U���S�]����hNL���^�����EN�rt3��[�Y�\2�N%*=^_��s�j�5O�!�����A6)����K�%L��#����D��աW�`��"W��7K���;$ĆBv������޿��;)8Y�џL<�Nz~.�O�x�*G�{�˾�J�`�{�i�U��1U��i(J��g�<pa��rB�(�Η6+�S�]
�?���i���P�AnC�tg��7B�м�T��q��4�,���MZN?NT�i���#�p~�����⊬�
#��3*L���Ί��o����H�B��yl(�+��J����J,�8��}MH(�Hy���	Y�N��R.�����B�x�E〘s�`-�u���>z�
D���|E�g����nz������!裵�k�3�E��G���p����g��b��W��C	��M&Ry�o����إ�4s�Jy��1�P s�!J;��T��7�Ĳ��D���|5`� �,��',q��G�����r<�A�ț&]�����b^���٥�����0�=Y+�G��o�FDzR$���{��<k�J��'�Ξe�xHz]>$��k���#�kb]������+��/����Q��;da�Ro�hk�n.�����ovGQg��%c�R0�zq����-��3<8dj�`w�6����R����B�D��K����~KC2@�-+�'=��Y��"4h���;Hz��66��$	 +��^��A�2�R$ٸ�By���������22�M_����i��+JVL@./ɭ��$��(O�D�Mb����Z�.��FÃ(<,