��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��Ѓ3E#"�7�Ӣ����{������R������i���N-���0'�a��JE�X�^�l׻�*(T��.ݎ�O�e�Ф�N�$��ռ�.�w%���h�s�`q�3�w��@�h�HiB7�D�Ya�?y4�+�}1Wv ������n�Z��T�^��B��xж�2ʜs� w��1��[$paل��'���p�y����M�	b���Uu�ϲr��X�0���S�|CD�(�휁0�s	�����<Q�O�KNR�L�1
�M;����DA�uf?fo	+c�����"C�͵�u1�i��^��6�YRd���yW����%UK�Py[�]=в��aqv\� o�Y�1�Zf-<'��
�_rt���L� ���|NDƟ���5���{9�"�&4��tJ���[1�C��݈�T�b5j�8��y��X*��~�"��a�/�Q���ܔ0R����}m��Ȅ(�/�ĵ4M~tel���X�'V�v�Kr���a�tW?hJv��z�KXO��1>�E�Y{��L)V_*/TJ>� 8
���M��t�ʂ"��v	j�<~J��1����79ǰ�?�*&��p[�Ŗ�Q�%��s�3B��<Z�uS�(fA9ɫJ$��y�����\2{�[ ���c *��K]ôm��������5�i,�HA�]K3QIG�KN�<�%�d��f�>�#� �zJ��$�0����c#-�(7K�@���*�KsyKjw�5?B1�ەHy#��lF�#�8���w��dX�-�Q�k��(i(Q��ሂU��m���:K�T�cG���O��q`H��TU �4#{N�JI��_�+��9ʌ�g��^�N*�THG�2���W&�7L�����#��I�P%�1齾i~O
��ߎ��L4��P�+�5�;���p��`N���8�n3nl�e7�Z�L�ӏ�`<׵�KT]ܑ�`���@'ڑ[�(\#�|l������TL�Q͵,��k$JF<��!���R�mt	���������z��$�NҖ��[����v�Ƹ`�\�)��l}	Ҟ> �0����� E�Lఙ�1��UAKFV��A�'�O��Mm�4��=��F��W9MԚ#|.�=��1�u����x���.�u����0ģ��Y�Q�k��vs�Š^|����3S2´������P��-�1�� ��ci��},��^�h�b�El���W���卿ΥN�o���6�r��(�H�T7��і^���z����:���x�;��Ǣǁ#6$�r��iAL�·`��p%��s�R(�g-�zr��f�ԵS���6!��4���Z�.<�U�dؠ���}�m�)T~�"��9ٍha|fl�}�̷�Ϻ�,T��r�R7t>��lh��7�=V��K�K��HZO#?�M*PF�z��e�x��fj9��
�5k�Ī�Me����Dg��ᭉ���eɒ�-G�=�qVN���e]"7D�l��o��_�!�[����@ �>�������V�b�{�ee��R�2��*i..ӑ����c|���Jmp����<����%���� �'q7��*�4^�Y��<e#��j�$�ڔv-�Vƈs+�Tza]޳rU���K���f��U䍰5��Mf��S�/����	3�[�EĚ�_u}�M����A�"ۭ��+0�5��O��&�v�F�!��6w3�>��{����<����x�}���iRl��|��e}{<7��\)4CS҄9�H/��#`e�B#��V¤�e6�E��N����h�(T8��t�M}�P�x���l)z�Pr�I�LA����}���C����}ߤ4�ڌI~������{�0��׺xYՔ�'2��y���2�u�&��<�>7٫Q�J��/�ge^M-Ucf���[ �T��藘�^�`3H/.�U7����,���~���R��^f#�Aׂ�BC��ߴ�	*���v�p����F�������5�AdE��(�� `.�@�GR�h�����&\9gV��s���]�z�
d��1s��1���>�f̋n��#:������E?6	=	#���b�G63������2�US�$�����knձB�o_�
i�h�]bT|�9ueOp��Z�(M�*���Kx�>hdt�b� t��-�ܵG���z��*਽��g� 3�y����UZ>�!�e2��%/�>1���F��_�R��x�S�6����z�^4�T�]e0~��C�9	��"Y����WVj

�\�z�����u_��0�}'�|�͜�F=�w�)�ӎw�����j��y9/��S�d	�rl]7����S!=�����Jܸz�Y2k)�&��Z��t �v��r����Ԭ��"�$Zµ���'��<'�F�J�4x�͜��6W�c�e���*`S�#��id������76��@��kƏ+��6��W����?�Q������c*�"4y\eCάƷ�8%����RjEk	pz��`YR8���0�#�(K�U��+~�-�2v���6JÉO�2���-Y�}�V{��	�ʨF1����T6n�~'iW�{ƊH�c�P�ee����'���Q��%�>�N@���*H;Uqz���T6�G�u�k ����:1+�.,������zϱBӖ,+�[X�`%�����M$Y�PCWˉn����Y����C��:�~�̖�͒\7hmi�_6v����V0Y�pC%��� <B;ށ ��g�(Ba�}}JV�bʹDF-�*�CJ.;�hS�~_ôqE�d���kx�xáE(�,���M|��rX�����MI[s�fH��#
B�g��L�j�#]��6 �䝳EV �@[�_���/&�x�a'��8��n+���h̐C�N�%�-K<��$�ͬκ�����p��h�N�,��	Z���~,���~�(͟=	vj��"L�)�'�j��s�*(�sݤ���F�d��*8� � S�/�qK�1��y����o�h����B�+��~k:��Q�u!�_p
������hD�5�%k��U
�c Nan�����G�?�G_����{[��)�C��_���n�
u�_���yg4�7�P�7���:6n�Jؼ�M��7�{�D�]{(J��y�������kW���lQP���j
�V���h^!մ��-&ĸ�
)�x됆 �L?�����D�;�Wĸ�4Ls2H�u�[�#�%K| �C������A\�����R�W��_W�6�T��;��0��*�if�Q�p5Y��6��N�nf�Nf��U�'�"N��Sf��氲������\e�8,^�u��$�����F����u2���di��JB��W��xs>���yfFd̎���2v=;�tD�)��qwy�ی�7�A��>%��To���H�V�j���Ž�æ���������4lwe��V!w���T;z�e����.�w�z�EF�kW��f�hd��r�i~wQo&��4-�OS��cQcg*9_��b�rn-䜛�蛉8��bE}C([�Br���ꔻ|/\�	� ��+d���[a�ഇ�Y�aշ*#s� �@��d�G��s��Ј��
��\5b\���۰s�I��1��g�a�m�&z˄���6}����ϓB��cu>šjc_ �Wi"0l��ϖg������WFD't\P@������N�"׏��r���1_���>�:��y���=J._��SC:�ݠ�����������P�:�z�N���볤R��m�+x�4�K��\�)ȳ�Ҝ�|�`N����ŦJ����J��$}>pM4�Kϣ��w9Dc쫜׭�)����k4��}x��w��/�#��{A����Ĕ��@W!�մ0��Au�r�n��p��NHQL]i�3�ѿ��H�=-�1bad���)�y
$iq)G���mϵf������#��ɑ�q$���k_�h���!�9���8G���&>+�5��ն�$��dnm淊c�K(O䚆<+b>����+��0F��֎��B8�*:��!mEQ�{�C 6�b���."�����8�볻��N�-9�)0
�LT^���8��w����o�B��G�b�T�m��o�à�-"�dI�\h���N�p����+�Qb.&u��a�4��T7#���}jbHu�]�0/����u����r��8��F15e�Ζ�y�cEx)�!8U�R=��%�M�~�w"�<^iu��m�n�,�@t$W���&Q�2\�-�=8R�2ShT#AV5�r�~Y'�#�^v�i(�b�tgu��>�<��_E/x$7
�Gɉ��p�-�`��<`e±¸4�������<�<c^� r�9������A�:5h�G߿�k^�C��I+]c� �S6��B�5J�_������G��M��6��n��XIFQ�o���G�1:��rOl��pqV���dfWX2�i��ӳ�i��?�QPh7�{�:Y�ڂ�I��w? �O
6�*�����w�C�\o������Z%H�P؍�s��ˤ��������4ޭ6�39���v�(_�=g��0�	%b�����ӊ+غ�{���Jn���Eu��}k!J��T$��)?�0��$$,7��$������������:���2o��=�����2���6^�y�#E�NgO�y5�hw�A��\E�E�CA�eF�Nm00�PZ8ʡ�m�4E�`gt�?�Ŗ��3��VhlPl��<KS���b% �Ի^=#׽�5�Y(h�_�����t��s4~U��-c.j;�r<C/������X���nWt��h�<��Hb=`�2j&�Y��o�lQ}ZBh���nS#}�o���/���\B�k�&�?�j���G���7UF�xA�a�4��VF��A�k��Pc �d�%]"�9����鼘T�����':�mIu��d��Ԫ�n}VY�m�*yY�Am�F�b	~�w�~H�D߹��^�$6���|_-sS�'���N%?�?b}:F�+_7UQF�~k�Δe�[8&"YNy��wt��i��1�|��� :���񩼘_vT�MDA�$hq�n�|��:�����*����/�P���Zh�7[���{~�G^)���!ɮ�+x�*5ܾy����yKՐAh���ե�)����	#�f�O�O^Eb{��y]�,�� ��hݽߝ}�2:�����#�|t��r��]s�r_Q�vS�{���8�Od�rQF�c^+�ޮ��r�A��T���5�)2MKϒb�&��7��6S=��l��6���\�j��˧�/Z������sI4;a5�_���d�4mؗ��F|��	y�U�^4^�3ա�0������Sܘ��P���,p���ʍվ;: ��}��tΡ�(M˖������;�-'v��u�pě�r[tIGR3�|麪U[l�>���ֱ��}���Q	�&Ą����\¬��(���Ǎ-��!<�L� �V��0,�=�� L�n8�Tn[��'�	e��_?O���ŸI��l��1m&W�QmFfh5�s�^g@b��'Ն�$�G�D�e�xn���;0E�P�RR{Z?��p`_i�$��4.6=��RZ�~KY+�3��4�ZJ->���5�R0�b��m�@%�D/���X���g�	��'T�C)��B_��6�G�d�w��q"�cϲt��+����ǶS���Y�g eB	���t=�3
(�ē�tnJ�թ�-0�-YV7�GO����c
�J��Y��*�أ0�I�a��:�����-��(5�!����h�E�~�E�K�	�_bD������r��x��g	2*�����ŮoT�Gw���+�_4SuYş���uO��4�n8:I����x$�&��Gb!H������.N#�T�F
T�zyu���	)�ɷ�>����K��&|���H��#?��T�T�?Z'�c[c��<��˼}P=c���m�
m[�_8���e�2.Z���0��ڦ8������)
j>�l��b�ր�SV�q��"φ\[�<NO��ûifñ�2�[J�~ށb�;���1Q��5��	�q���wT�����#�#*��Z$p�����E�Z�VM��>�Ei�W$_5���s��g�Qu����0���Ç���A��T��˗�/޼���� �Z�q�
޳��]�]d�H��u�C���e}��o��2��b4����F�����L?n@�W�����5�]W@��cq�-L���g����ܶ�M'���?�P4����]=�L.�S���

-��k�'t�R&u��W=j�2�D�'���Fo��9��=�!�ԅ�F'�`���8��Ga���������; m��X9cAU�p�'�mtK�s�b�M&��<0r�{Y���P�.���[>a��T!�Am�ft�iK�ؗ��t{�^�a���8 q���כ�Xh/�6���� 0&!���\",W��'��qL�����S�����O��ǡ�/�f�5��<7�'�����H����I�HS���}l�}f��+6�������� �.�T���c������j�V"\sDnRR"�d�T���d6$H���յ /i�Zc��������Q����{�F�?�]�/8�V�?��jOu��l�2MrY<�$Auf��{�zJ�����su�+.���z��v��=�T߲�hƨe�`���<U\�z��ܭ�b�w)�&pz�|M���(a7�<�G4<_:�i�8-�EZ�T!Og��Z4���*��-��Ҍ��S�`�2�t��I�HY{��wכQ떌�.5�\w�!��3�L�a�c`Ga�IgCG�/ ��uw2)�H�����aW{���!�Rj쬕:.v�s���!L���yI!�'�yS.�=�ê/�=�Y(=IP�߫:��J��A�?�7��9aj���A�T�I|(�f�E�J�6r�����"�^£�b�.Q����z�'R��ylJ�����<�M�d����cĻ2Qh�����z�������}���G�$���<��[��Mc�[�FSõ~�����U�:����}1�߸�v������"C��W�hm��/w���qր]���ܵxga���!��N w�<��}?K���ojX-��` 9a>R��3��Λ�T�I^fy�/ܢ�m3��~�"�k~&6i:Z�V��=�K���ady�s�b��&�E�w�y3aAN�<��tQ�1�R>'	�g{��_�`�ӕ���K���9m�<6�eV�j{��3�4}�%���.��/V�d��=�e\��s�$�mPV+!�������v��P��� m�-��֨���5v��nU�I����5�qH����bmi3�#~�OKN�+îЃ��u��+���w��SQ�E�t�B3b*�E�s�x����V�+u�)T����6�@Iϙ2�ج{�;؈�������:����Fa� ���L-�3t������G����Y��� q]�i��*ټ�V�!���Lh�#��f�߄(��ߚԍ�ࢌaM��j6�`�<Y%E!���M���h6"d��Y[ˏ���.~��8�J��5��!�#5q���=搕04�@Tv�l��ْ���s��{y�'�����TS�	`2/=2b^���nك��l{ҿR���ޗ��G�N��qz�b�D������ �l%wB�4OCHh"��n�(Qw��S�X���uj�����]�� p��4x��:�ߘ{�6�t�B�����Xi6�Q�
��Q��h��:;�Bà�_�����&�����@[�h�zO�R����Ri�O��4��z0�Z`�{��k沞9"P��6��|6����j��,Q���x��n��[&�[��n:�~s����aK~�0��ڷhu�F�3/z���}���=�l9��Ե��b�� ��-*
1Y�e1ir���B�@�ߎS�$=��%���i�7+9B~����媑���BKt�(|�ҫ�=EF��}�qKUH=�Y���jt���"bz4���V�� ������ZP�~�L����{� �*ml>���'$����`#-�?W4̓�Щ�y8�\R�-J�r&GJ���^��ݺ~*��R%Ƚ���,�2'S��~��z�6�Zi�n�3�OtkL] ��P���z�E�.��J���q��v=ZS�ɗ�K�D5���y-�j������=�$d���.�:K���l����� ��腝Z:���8]�a�&gF�ݨ����AW���j?z/!{z*��6f�!���{]���fa#M��kӃ�@�O��t C���p��O(mv����c��R��3<�x�7��ی�Czlן�.4-#�w2\ha0�x����$�x�(�-s��u�K����B�4�.�+���%��r^1��=�]`X2f|E����>%�ˊP*ٱ��nX�-��TQ�$+�%������ۊ������{�n�C�*���߯;8r'B3�N[������G]�qI�N�Ѡ�~w�5J�f(^6xx��aUd�<�,f���"����<����I�db
��s�"8��M�����OJށ�z�T��d���,n�Gn����o��xx��ͩ6��h��*�a�]R�����ս³�7���E�ZfS�+�osҩSRZ�g,���*W�Y?TO"�,zN��,G��Z���NO1�ɤ��= T�FG
�u\�5!���0�y���L���W�XN���um�x������2Rk���E�$++�N9�2	ӂ���ip(����������MR<iU�W#me;�g�A�-^Hv�yxH�{8<�pv��2d��Y��w���i�6�t��r6⛥2#���H��ag���
nj7����ɳ"7gMc|����y�<� �' Q+Bi�	tX~��m��	��Ǵ����nv�u��8�
 b`��#)����Ձ\��-T��F��(J��F�XN@NX��0b4�薖�X�@�*�V+R��W�i��Ʌ�q%�V����D�e�q����m��^���g<q�U�M�qm��/�s��4�����Ϗ�|��+;y2?ha���7����]?��3��>���zI�!��j�4e�����K+�ƜR�U�X�����p�y�u[c�?�(
���-�V%�h]��F���i�(JF(+kߢ�5�:���ƿ
ޣ��`�7��߫<V�1�iJ�籸�Eg��N�����Y�x$�T֓�OS�$��koe2�ոw_e�uQ�~��k���̍s�x�U��Rt9/MS
�C����VQ���&��$�V��#�Re	j7����~8}6(�(���Btc��v����[�"ܝ���b� 79`\�F��؍ߣM��5�'�!5�7hLl�����ڻB�0��L ���rl#��s��WE+�۱gu(qS1��a�뽚��Djt�����f.A��3k&��3�ٵ���z�%�YM˽|��os�Ŭ�;&�DyΜ�y�S�������3�g��ਿ�����Y�)�3�s�Np���鼙G0!�x��LX-:V��+`BM���t���G�6���e����t���:.�V�b+�z2����U�ǜ���g��g}�H�zXE< �����
��'(�k)���d���#J��#߫uF�TpP��(�k��c��R�|tv˟4��/I�SFTp䆶Y(�[M�� R(p������bDtB�w��/�x�u	����`���Ē�.����,^ ė�2����i�V&W	V��I��������H����� �� cxl��J^�����@%=�e�(U�X�b5�Kaa��q���͊�(�w��/����x��Y���yp�Ո^�]���hSX�t��"ed"�D[���Ac��t� &����O�1����4I�V@��twN_X�f:�s��#}R�����C�������#��_�p��?�5�(�|�2]�h�q�|GM.�=�@�$�k�=���蝋�8�d�u�",{g����.ȫ �tF��sGzv�����y��1HD�g�z3`�������#%�#���a�c1�:U���w��E��\�^��3�m��J@N���=f�HT�u��J�d:�V�͂��%���lٟ�	�ai�`��˒�/�-^x@k��`��E�"OEy�yߤ��Ǎ�����砠x��x�VH���k��dl���e_zY=����v"��K�w%>s�X(�pů����F�vO��ŋ���������Y���B��D����p�+��Y�J{��dE��7��e)|/0<�C���{�}NյVϰk���>;�|	��
�F���� (� ����A�0Z�B�����֕w�}d#�tU�8����:���jR`Q��h����	�9�����?����Y��\��Ɉm��-�P�k1o��� o��dV���_+���A��qV���N{� �]+N�K)�ݔ��?���P�*�H����~��ռ�P0p��=�Bᚪ����ß�%�v���v#�4uӰ�� ��Q�q��F���F�ýU���p�����ߺ�/�Rb��}�n.Ø�Ø��f��SíSq>���Ʃ����-�\j�.J�`X�"�����9�������mx 	�M����ƚe5�׺�H#;����(�뉀D��xLύY~-ss1?]��Z��S�Y<GaD�k�
�+��EK쮻�,(?x��N�(js�z�M:�=RY�u�P�ۃ[��x��k�Hۣ�'�"��f瘥����pZ�$M�NN���C�J��>����O]�R&Ѿ�ʝ���9N$��Ѕ�T2a�}��g�9�f���LP.�� �b�@���,ik�D�U���}����)_gz�B�t��G��|�ٶb� ]����y<,��}$��*�OO����C�)����	
!��P��?�?R�@,ǜ���)E��ہ���j�T�,)o�ݳ�P�΄��{2���B��J�ߠch}�~4a�7h��=���Xr|����t����q��~��)�/�q�����q���*C�������]�� H��pA��������S�o��W�Ɖ3��V��n��D���q��%����U�"UB�Y�Z�t�i#�����>��n�iL˭R�
`�ے%��T,�$[h���Aj�Q4vr"W\�.��u�[ $[z^��>��|
���o#����l)9��ë�� ��֪W�%�A�J�`-�2���R��E��fB?��r�\��3��`���"_n7��9�j5Cd(���̳����e���r���GY��sQ�4�+n���q�[���X�A4]�����#�,���V�)|fTo��ϊ��hHVgC� z��9��6���c�td�Xú�cg����	���{��p��b����Y瑅p9�u��lK���;��k�:���y:oΌtOP��uqBq|1J�i֏P�;��Y6���CU@�"J̺}}�k��7���S�u���n(�T:�r��