XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��a�3x}�l�z��[M�Xz��:.��%���#��u�G`���l��vQp�������G��t���� �$�&����턁9��2�ڸ�1�q�W��҈y\'g��KC��.ɬ�vA�nz����f��N4�M<�+�7��VI�k�K:�����d�����Gٹ2A�D�s-��ǩc��°�͘�Q���[s���C#ڡ��s��7)����2��V�O݌�RN���b;S9��7�Z��� P��<7X��Z9x�e�LS�'/���P©��Qܱ��.A*Q�*��u�,\w��O���*�*����L9�L�ݸv�4�6��_��x��谨t�o��~�wF�|�k�5����8��<:�S��no��FYs:Yv���~����AwGD�3��X�#M#A���t�u�JPg����|z��S�w��P�qW1�S���^wyJ����u[0}a���G�I2��o��y��2cvZ �;Ր(�MꂦB�W����D>�ւ�^q�'�

���'�s��w�0I"eP��.�Q%��0o�7u��T�&W�T�X�]�ԥW�n�n���kLl�To����!춖���;�m�6��yօM�u=d��[+һ�<�~}g&7?82ן�L�.]�X�/1��c�F�w�/��mB�DnA[[Z�D6�ae�Nܯ0)g�Ȩ2��$綱�I)�Z�h�� �"X��Ì���o|�v��x���+1=�����ݴ���'��FAr�a7�,q7E�ط!��XlxVHYEB     400     1a0�`/���>
3�A��HC���y��iY���߽��!��(�-'��u�
Xl/���"�:��/n���"��F�OS������C�"仟
n�y�tQ0;\���h{�r��^��Ta�m�D��~��k$��o�[0�]�7�qJ�ʟ23���?A¹}8fӭ�ɞ}H�!�l���4�l���-����M�O��-�d�|���4D�T?�!~j��:9s÷7���YsO�3�ՆgX�&Dm`כv�Ě;��i��S�\�L;=�봻��_���uۧ���h�9Q�;z��e����S訁��Jm0s3�'ή�f]���k"U�*]����-�GJ�{WdDlڴs��}���ߴ�Ռi�`2D `�� �7�٣�S3�����w���6�3:���V~�RXlxVHYEB     400     1b0}x��l'�dyo�,���o�0%��1Ae�5���V�����Zit�r�:���R�B-E����e��he��,C�'0E���?�˼(��h��1��FPĕ6�	�[ �1�j��8>9*}���"NAW�:���:'��W�T��x��Avf�A��@^�)�� ���3����S5��=g�}J
�� �T�be�f�J�<��fm�T����?{p!1��O����8K��x�љ� VR���'ٽ'����%\b\N��
�-�<.{E ����M�4��D�i�(CR��c6�4���b��|�J����<�d�E~D��Ҽ���6ޚ2�v��A���7V5?�N�h�.J�0��R�s�����L������{F�b�.Gt��zև z7� *QF��yxj��?h�:�����>�y�:�i��"��A�XlxVHYEB     3f5     130����D�܃�.h�7�~���<�H�:��3�y,r��bwY�R��B�Ɏ���r�Z:f��a)Qߘ��8���+�Fq*jh���  �ٮ�u\>ޤn�~b���]���])�?�z���	|e�u���wV�o��YI伊�U�2�2&�w9�����f�PZ�#����P �,� �\DH4IVU�Ы�� o���4�R�~�C���	�]�&�+!݉o��҇�\�I�?E���𺱒/)ʻLȧp��^�\LM�4�%u�PSs��nH���n�4� �/r�p��������ńq@