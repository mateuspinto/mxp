XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��c/�R�!r�����c����dd���42�V2���R��X��a�ۇ]\�v��`+�F(m.?�l�����G�F;"O�2	���i˾�Ф�Ф�CQd����Ag�G[���3Ƀ,���!��x�3P8��Ę���<����W��v|Y=�.���#�y2�>�c��/Y#T�˲��(�W���,�0Hx�R��8�??��l)�(0���<�0���).DJh@�݄��v��;�qu�ɉ|�����P��$*��B(5|��l�^�lw,�Xȧ�(�T!ʷ�9��#�a��H*�i}����O�ia�?�S������=\p@�7�RH�6����6f��r�Rͫ�#Gʧ.rw������y?�WTa��ۇ���w�@���S�#W�W=�䖀�(���R�[MH�tj�;#+�,s4z,��	לx>�_)����;�ɼuW�P����t���G{nG����!Kb��$*���Џ i����_}{N�`�))�w���D��'�#�aؔ���Zuy�4���������,�t�ק��H����Q!}�a��H��E�O���>9_�T_!t��?:��d2D�=��}`�A]�ΌV���҇�:������1TBW���+��K!�YRI��	QW�=I)��U��p�˘�*e���X�Ősy�'T]�ê�4o���}�َa���j�!� 6#]Z�F$��GS�Z�}B6АĖ�N�AU��b�6
d�@�m�?q2TD�8H�l�,�m骖�CJ�?���H%XlxVHYEB     400     1d0����ޡ7p�T�?!�!��'ŹX�,^ƷF	$\A��I�A��fcٻM�&�#`��������k�fP�`ă����2�'�)�-����6�ZD����3 ޢ���(T�:�k�.{��k\	�c��kJ��c�����_��u�-Ӻ;��i�ilY\>��<�/}9����uz�,;},n��1��ZJr��x�EN�I<`�C� ��A���c݆�A4f$	�M�sE�M�I�p��RFW����]��0�j�%̜Y�Dd1��N�e�-����,����§�G��>�< ��D	�p�X�3�ń��fK퍴�Љ�B6�� �?v!!�V�� J��*��M
ݷ�9��q�ΰ�(U��)@�*�s^.-�!��;���Q;t���i�fR~��	'����������_���k�F4;�I����2�ւɅ�70(m�tD�H��p�;��\_�u�wXlxVHYEB     400     110��Ш{�����`�n��;^�N�5]0�l�(y9�2b6�i3�.-C�Q�Kgj�=�P�a�i� i۞����"�i�+.�Q/@
��`jo /(�������'��`� Z�x��se�5�c�RM)]Ѹ�L��#�F�m��G������� ��<V�V��^@I���B�7
8��![V���̏W|��W���CΣ5���S�A��'�s��&�=9ɓ�h}�_L��V�e����[�䫇��u�7�Ƽg�B�R�����q>��XlxVHYEB     400      f0������?H����v�?Ӯr���K�8HgF� 5c���G����dq��������'�}�������ǜ�J�GY�.݊����*b��D�7�M��9�.�!�w��@��gO۟*��ۼZ�%����m+Y�uz}�H�	w�Zo��5����ON�����G�6.'eM ѤO�5碰у �6�3)�y����mp a�$�Ƒ�U��+D	H��O�@�=~� ��簦�j�+XlxVHYEB     400      b02F�j҉Y�U� (a԰&�eCkk�]w�o�-ˠ�3�ȱ���I^�cS�t�>Ѕ��·c���)�A�
_
�-b������7���*�B�?�qf��we�'&��l8R�����&�+��b�(uõ�񻗬�C9>jF_�ݣO,X;zZ�M/�p~|��F��+Gx�3�/�me-�XlxVHYEB     400      d0S|�g�j���Nϔ�M�dZ��	����nm�T������/OD��Թ¢�,�I@h���l�4j�1��E����
k�܆��A��H�s.)�]�a�h�!�SX���9?��5�"�Eg�Dt<�llϲ��F;�4:Z��y��I�J�޻o��^��qњ�+R� �S]�
�/�CW��˃҈�w%��I;�.��"��`��3�P����a��R�`XlxVHYEB     400      d0��8*�/쳆IE�i)$g/�>���/R���q�ݺ��[�e�WS�kG;͖�����bͬj���/}���Fѱ�-��f���s*#<C2�vK��7�KhuAR�j�g�A��rg��M��{1��|��w.y�:+��t��.X[�єn� !+5�x��ź��(�� =d��,�/z��f񌠚��Tu���a�u�]XlxVHYEB     400     120�CY��x���r�$2���	�ӥ ҉�u�$,�՗/�	�c�mqu>T�������"���0�Q�XR#�T��;�,F�fN>%�I�1���(�J�𰓶�#�&ԗ�	l��RP�������xܤ,��5���o�	��f_�C�����p�3C$�/�D�D�kdh�����P�u;F���=����p�x�S%��٘O��!<O?��QF�m�F�� Z�����=���n� ������c����@}���@Ǯ{ẻ8b�վ�?]��&�et�٭S�Տ�XlxVHYEB     400      b0�0�.+�yNN� Fop�s��n''eb�l�W1
I�5����x���q5�L,`�QbR����}�3�o?Ns{�߮���o,}@�{P�Ԉ/!1��g�F���q�$� Oj(�{F����%�R��n��D�̟5O^�"����{j`�����ʊ�������:9Ŧ؟zt�XlxVHYEB     400      a0�'މ\ۗI�4���V�$|H=1Ɋ��>7ND��ءF�O��(�x݂5yiM�6�A�l@��i��Qy�ϝҚ!�������8��?n!6$cc�H˕9kHO�f~�}�~�SZ?�#6V�x �?���πo��E��ے�X�;��
XlxVHYEB     400      d0`T#SA j����0�E�*���ϤE�����BQ���/���[�q*�_�+	��y�mN�����SB�:;���ף�Xݲjr��}+{��x+��Ő$ ��T"�,��������qdvR!+��v�J�; 5�e��i�
#Rsy��ۉ���j�clz(�� ION+���!�dQ�[�uߠ��ڃx7�W�?^R�K�WM�`*>��lQXlxVHYEB     400     180.e&���3�^��UL�j3��p;�����AYM�X���:FHf�1��UJ��:�ڌ��r�5z��CUb��~K���Ь��]��\��z��
�h$���X# &����^M��$���˛B��g}3�"�$o��?E꤁�a6��pW7?�D��8��nN~Y��L�ŪX��)3�Q�̊0�-M͕M���,vӉ� �:�6�'2�E��?~��Q��EmHe	�hJW�����G%�w�&��_���qtL��D���!ȿ�M~�W��	1uH�q�$�Ȭ0��C��LZ��0�Ox�kn��t�7�y�I.�� ���2a
f_H�ɷ_5���ժ9^̇1��&$U�~�����m��K�z����^�>g?w�ks�XlxVHYEB     400     130��u�-V�hg�4K�Q���)& U�#��N��9�Y֏���7��G���s y�؝�7�ڎϿf�W�z~�Ϲ���g>�*Bb�}�0�_�	z�xOV'�ב����5�6������C�!��<���O���5��;�y�03&�X��M_u~�J�����A&� �!�A��[�8!hE`�ޱi�>�W.�}�ǷR���n�;�`�q�#�xk�)�쨰��<O(  �zT5mzA���������a�V_����SԒ@���G2�?v�`�m����#�R�>��}MVio�XlxVHYEB     400     110/#��!�g�,:q2\�xH�/��p�k�����+p�{�؟�K~]���ެd���s���-ļ	'������NN?I*5��#|�<RJI��5�(��[e~xE�Ɣ�]̒�k�5�ǌ�f���X�	gv���>gC����hˡ���3.����nG���H�����
�}m���h��:��������h42��:[�v��$p�����`v�F��N�.N�3��M,�U���(����Vz3�E���e�|��.\A�?���XlxVHYEB     400     190�fO��o 蘀[X�%��7B��4Lf�����vMh��z�:�,$�˘�{_�_P�g$��S��A�D�~U;��d�͍�S�G�A��H��%�٣�=�ʍx��w#�˒�2��u�����	U����S�z
PO��
���&Ƚ�m�����m�j#:�����~l�P�h�B��=16�o)R7\�cxEJf%�JX�˗+�gEee�XWT6-�KLM�������iz�#�}Z-�uv<����5�7 ���0�ֶ���ZUG���9A���Zj9+�;e�T�3La�R;�mQ��]+�k�/"�:5��
�K�7q����7'��l��=U�w�}�Q�����b�T�;�	;'��g3�Q-����&ћ��q�"_s3rw����XlxVHYEB     400     1102Uցc��	ʏ	�{J&B��!�ܑՈ��ױ2�ʵ�����9%���'�	�t6������<�g�ɨ���]��&�U�O�s�>fU�g�B��l9vS���mqxn�R�J���R"��_e��1�Ї� �&����<�Xe%���'��P�J�Y�u��}׀�xr�^�KN��E�L@��U�@����QX5��kի�U�;+`�{G�Tܢ�=��J*>��x�С�Q����D�;|�m�`���� )|L�^����CXlxVHYEB     400     110o�ёd�5.Z��-��F3�`�+_�l��A���(6(#7{؎+8��s��,j��Ês�|��p��S���c��w-	d4n+�`Z%�]��%�;�Ꝍl�S����y���V��e@-L���B<'oM#��c趶P��%%�.���j/�<љwc&+:c+Ea�P���5��@$� Q�!wA�C��U��ƽQ87 �*q2�¿��HZ�C�����|0!~�����ps�|XV�����9�0r�ߓA�l7�ek�ϒ�Qt �koHx��	-��TGFXlxVHYEB     400     110�ߑ0�
��X��%ܭ�<� ��Z{}��1�v����su�:�F��,�G�o�ش�klE�G�q4h� 	bY�XK�N3�&�I�T�D�?B�XM�?Ǌ�2�L�����,�Tο�;�-"������$����T�M-[�r���-x�O��6�MDQZC��*0�h����񜉰SK���Gk�#H!�8E���<�lԉ��P!��UB�$��ڳxz��쾉g! �o��B�:y��A�	�.����m1=s��F��ɰxQ3�( Y��YXlxVHYEB     400     100e�m��H��ޫ-UΑ�w��!;IG�����x�/lf������ �^������i�f{]���Ө�°rn�W�nZ��I�=�w��W�q�k�l?��OG�1C�1!���kZ,ѵ^�s#��@PՐ��?�H򄌺DL��PEX�"}�aN���*�*��V?����FM��3�#��An�5ԩ�A����Nlj<z5+��X����|�(���{ ��~3nd��l���x7�!H�J-��XlxVHYEB     400      d0>�K�����bp.@Y<%��cm�7d&�Y�4�tE����"��+<"��Z�!��9� ��P��Jϸ�����?l7˘Qr� �@��r��5�����}���8���F��7~��J����k%!cw�Dwc&�Jx7P��nz"��ܥ�ߛ��n�n��:�y>OUN�5���p2�/Ԏ��Q���JV0:�e�'�HRe6�D2�8N�XlxVHYEB     400      d0�^E����
�P%�E3{3׳�W�^	��-�R�g��W��T �ur�v`��;�8e�k� ����5m������rkE����M:����'f����7�����OƑf�]d�Jnf<�̅�"DI�Ĵz�f�u��d�i�۫L���W8����N�Sv�I��|V��!3r��ކt8�/�9� .�>�wZ%@���O/��XlxVHYEB     400      f0�r�N��O��y�jE�LX�âӠ�C<��M!:����B�+�Ȥ<��j���Jm�$�b�Q���
P_��'L|LE� �h�E|~��?��m��RT���8(��ڍZ�l��nL��1���]X�����E�n��{����Wu��3��,�Ѳ�h�`;��"�~p�V���F oS��,� �m�?�x4��n5��h�N��h�O�G�HD�*� �d���qHA	�N��o����.F��XlxVHYEB     400     160L��~E��*ho�܈{p��y�E�Ĳ�����BKٹ�vf��h��'cAM��LTxA��ˠW�y�/B��h���e�@6Id�B �i;�P`����w�$p�4�L��P>���l�C#�E�~$߽�g�5�Y�/�䗗z1u�'��ե����� ��$oQ �z��8R8�wв�P�8N،::�>��v����'(�ձ��L�@�'����UV��Y��hЗz��ȳ�o��O�s��B0η��s>H|�����`�r�[e$򄛞�7%��!;*�!��`S�8�I��D_�&t�q�!��G]'��yiW+�gc�"#?�)��v��ʤ������_̂���,XlxVHYEB     400     150���f�T�Cs��I�)�G�!`=�Q�äW�?tI-2�.&:RR�a6�`4�^�+�u�~L�*|�y�b��|�E�iz$��P�*��{���˫jd������[q]�;�]9|��g�(��A<e8X�;5����I���Z轅��PL���䲬{�iX�Zȡp��'z�r5{����m����۠j����~���"m���xx;�s�j����$u20��Q:�w��.O�sO.71O�i3�e�%#�PLx�����F���H��>���#Ɋ�2��zu�e.?�ҧuɝ��hG�.JZ);�2��M�*f�(<ng��s�����7�H�X���XlxVHYEB     400     1004�w�j�_?s)��!��	ƭ��
�$|�[P�i1?�,]�?�9�����^+t�ռA��qȚ��X�*Աp�z�l�.!w��b��
�
��_aH�ĶY8���Z�����}̎ 3]P�7zM�b�x{�l&��r�h���hC��9��-S���i۹s�*��XB��Bte��H�����M��H�"��Ӹ�r�"�&����^9T��D�L� �ʹ�f�or`���#f�D������MGDטR�t5�p;i��XlxVHYEB     400     140BJxj �4j�0Ȇ��%��#vE��Y�SA�/x8����������ԭ�+8��E�lR�::G�`hU�h��u�]
�!Yc%��Y�?x���Ϣ�։�.D�j�� i+ލ8x"��U���H�V�g�Z1 �
+Z0�e�T�ݒ�Tˏ�d=�����*���t.��ƕ9��Z���J�;ޞr����<ȏx%�Tx�M&S+}�7�9ک� �tk>���e$^��֭Y�<W����}�FMqB�������7/���H��=7���*�"�'|$N�I�.�&��Nf#Qb98�����xΛTȚ�Vr��=XlxVHYEB     400     140�/��lMw�/C��Ĥ�I#EF{�
����`�'V�u9$�\��Q=��*
��Dv6��2����)w���	U�LeA���Uy�y|�Ns�Ŗ㰊Z?,����pHh]��p�Orj��υ�ۍ�������� 
��g�JS8�GQ�͡�� ����L��c�,�>�m��ӯ��)Ih�/�<�i���ۯ�Gaf�C��_r�Vܜ�?>����`fƵ����+�L�W�A�R"�� d+!�����u*��=�t�$>�5�tV�>s���M�=HUV��\c��f�� �#��	d���lCW��SQ^wW˅��R�.XlxVHYEB     400     13061��(�]כ�ٗ�-F�_3��{�.�%��ږX�Fn���l{��2t������S�M��� -�!SÁj���U�<���(-H� HMP����T�+���9��44~-J
�m�kv�T�f�ɑ�� T��]�%�rXʻu�]�K�y<�y�����Z���$Q��/Q�+R�!^�F�g�^bO�����2�'ʷd�	ъ�tw+�U���3�=�E0��U�#٤��FM��5�۔(�X���H����&�RTVSC�|��`�*�0�h(ކ*(>�5>��w�k���v��%@����� kKݪLXlxVHYEB     400     120#��?�teCz8l�p�N�{�y`v2���SS�P2���imK ԇ5,:��V:O��: ��K��ψ�T�H^C�'�����?yI���{zQ~K�z��rG0S����'�2��\�L����9w�Dɯa�j���C�\[(�%�e��1�)I���bO����W�C�A��$'�.v��lO�Cg�Ր��w��-�.Y����R9�Z�̢�=��R�0U�eR=����O<�-)d��oq�{��j����e1|aʸ�l���F$�(���.Pp��<x�XlxVHYEB     400      c0��@��^E����J��'�-1r��&��vf���h��~&K G���܎�K�uҮ�[���r���K\���K�]��E� Sέ�u�D�dɒ���z�P��>ī����T�hH.����0Zb�_��0�%�������=fߥńL?��Z��~�"=K�^Y�V��Ȣ���y�,�k��M�	�%��XlxVHYEB     400     120�`-�������6�~��8Ih�E�Zl�yh��^f�%8Q��IZ�B4���|r��DUz��r�a`�j-Yq���>�EF1I�o]E��`�������_ic�N���p^��kK�5�ҧ R',OI��*�֍�[�w�hz���~���LCfZ[��,[����U"i�v ������U����Q�EF���1]�K�RU��٘�\�C��b�����\��C�#s�t�{U�c��P���-�\��3��")���M��Ga�<S�{�� �q+M��&���ʋɬeXlxVHYEB     400     120�:�=����n�#��&|��NM8���'�K�ES���r��
V��f5r�J?;d�Āb�S1<>MS�bl`�T-w�HͰrf�t�W���h�w=[�Ƹl�9Rƍ�����U�
+׉�����=�����rex�S���E��^����ܗ�#'U0J�q���	R �s:S�9���}�^hH����ג�uD<��̥����h�)5T���NX^�Ӧ�a�F�h�8��>��v��Ŏ�������v\(˂`�9�-�d�ycᮻ�����b���cX�~Us	�8�-3XlxVHYEB     400      c0v�CGQ)���^��u�7̗�n�[=Ef.Q��D=��z�%��%<�0\����w��IX� V. �|Q(*Y���u]<��6����m�q�s��!-[��D`I�m��y��0=3專w������ ���M��߈������lu�GW�n����&�a3�I�)�c�<L��ӟ"1+R�xBJ!:�� 	�s�cXlxVHYEB     400     120�;S|��qZ �x�ݣ�3��ↁ��c}��|��3��a��x/ζ�Ί��Dp��}����yE˖���Z�"'��q�]�\KȐ@� ��z��=ж|~@����v�G���ViӾX��\I�>I�'p�x�!|4�c�����M�[5|+��t�Jg�4���L�ʬˇ��o���󩲤:e[۔>�惠T�O�W���r�b	��$!ʨ;|��
�Z ��,�3�ox�j#�sm)��W(���D���w����Ff�h��}�Ok��0S�µ���\��9XlxVHYEB     400      f0���f�4d� B�Һ߁�����Q�ɮE��Gh�`�JUx�������Yf?�RJӾR%p2�;��ZN�ʮa�@����! UMp�V�cB�鯎�n.>�^���d�0����OvZ/<�
Qq���4M
H�g5��U<������2�a����]0�����F�f���d�dU��%d1a�;EAx�d���"�ob�V��g�J���ξ6���Â��7<[�XlxVHYEB     400     1108��\1]o��ғC�r���F���.��o>��@=��ha=0CG~x,D� �(��nթ�i��B�e��W�7�3��qv Y��S8ɨ�ۗ)=8��W9m���W_٥��W&S13Z:I�_�_)H�oZ�ӑݨgfx0ڨdcZΌh ���-��^`Ίdn���N/�H�g�ll}�9������nnIhv�M�<�= ���� H����f���tP���D�v���Z�Tq|�X.��}ˋ��n�Tk�Sћ�&�p�XlxVHYEB     400     120GHK��r��"\�F)�A�����e�A8_7���7Z^)8(��]���y��A<g���6���1�ÄkO7�n��F�dn���2�aކD�g�2��RR�%���t����Vl����%&7ה��ʂ�e�	��׾� N*O[L�c��d������q�UK����M�n��cO gip�L�oR��˟�������+�$ӹ�)i��n �o�f�o_ڈ�����13��B�8��_ؑAL�cs4�~[4��h����������A;5]XlxVHYEB     400     120�Bd�H�)��+4�u���� �4�53FK�~�G��-�4Z��j�l5���;�e����z��y����r�1lp����r�z�<4�;b�yw��>f�>5,�B��aM��H�_V0��ZA����<�z���D�`�}j�w�]FHr���t��8�[�L�_G���8��,Q]�S�U��G	���Y�e���� �&�hy��S8^����p(����C<���7��-�L��s�����r�8U)(����dP��k~C��aĺ��%��^>1��/��XlxVHYEB     400      f0\=�� !w����v��9ٺvE�uR��r����B��ԥ
�0`_������r��}�n��<�Su!=��KLc��/���K��`����|ޛ2�FP]���h�=��y��<��(+���V���&��L�U��O�� 6v��?���@"T؉[���2ht\��@v㑓�s���&����|�2uy������.~&Jޢ	|B��Mg�
�J�4.�x}$T�fe��>f�P���LXlxVHYEB     400     130�R�?[�J�m�'��(�Ol�	�v8�0��Wj,���UX�m�a����lѧl⻲���h8p>7B*K���'���J��M��Vw>D0�\/ZoeS�f���j�ԍ��@��|F��xh��5>aP�~R��{G����oK���T�!ћ�r�k��s=���!�-�����HI�;V��o�Ɛ�J��@eE�>qf��)Y�k1a2ߩ���ޛ�|�i��|��W{F0����܇#��/��FaoMR�� �(P<%�W������E>L&%-~��T�r`���(m^%Y�~�1�A��W�qBJXlxVHYEB     400      f0W�sa���LR�!�4�w0�/W��!v��͂�<����X�H�v�"�O��#�����ˈ�J���'F�Z�� ��M��E4�n{��UjfԔ�i�C�ή�1���\5{v��<��C
 �b�n;09���R�B�~G�m�#�F^��������h�'��&�yI-��Ve�� P�k���8���Z{���U"���B����yYrAХ�/��=��O���pD��[+K^��XlxVHYEB     400     150�Ů�����w2#��@+�]�iz�2WI2��:�u5��vsg��%'��K[Nx�&#4h�9!�U��!ƥZ�"��Q߲���'m��%D�x�o���9X��wb�A�~q��H�(��CК�Å#m����n$þ�3�'H#�0�H7��Q��<
�{����=����\�3C��h#4�'*��\�̺/?3�!5�O���|��D	�hq�g��f���@Q�#�����/y�����&�@����E�����g�f�$J'ή�F�"8M�WЈ}̻��2���I<���̷	�i�7�< �i�k(�|3S6���a���XlxVHYEB     400      c0=�Bi��Ù:�Ѯ�FR��D"���+����06���u�O�m�㬽�+����$��s4� ׌6ϑ��&ٖ�i̵ڕ�Yӛ���(Ao�3���n�.J��g�?��K��i\r� �9�ma�3�k���e�'��z9�cy|%>y�Ò�e|)/8	���Ev%����XKeR
9E��� XlxVHYEB     400     150ä�kn�go��
l�	��4�U�kx#�LrȰ`GǮ�ʼ8�\�V=8����>�ܪUJKь89��x��3����=����� ��h���;��W:���o_����T+��ڙ�S�}�%Y�1�	�P<�I	h�p�����X�!��p�>��R���n�(�o�>�G4��H<Y���Ш:&<>H�=���&{E�)|Z��Yǃm��/�5���Qj6�YL�� ��ﻚ��[+�#��� L�T,A�M�\��z�y
S�B�*�:�K��tGz�֡]\�AuD��x^\M:>�Xp�ń_g�x�h���u�HK�e�{ڞ�=5�^�gy�XlxVHYEB     400     140AF�.��YXL	ű�hn������Ҿ� #��K�#y��X��A��k��}HWFr����\�����3��Aŋ�t+�}���������=��*��l���8�P!�9z�N���TH�)����#�"S}Uɂ$>ؔYv��#�5�؛@��.j�����Z�BG�|���p�贯Ru��$y����ح�V	�_[�%B�>���D�#�([�cI`u9�X��[���5ǺJ����D�l�L�-1}ڜ�Ĩv�
��lv��k{��x���Y��"h�z߭�7�Jn�p-j�ir�n����8��5;��$�L��XlxVHYEB     400     100���9�u���mKZ*T��U���c:�����W�R��'9�$9��a�5���$ʞ{��OÑ��-��av���n�p�y���&m��m�\)��)~e��uy/{_Bnk���%[��9����%�7?�� NjVu6d�t���W���U�$�EW�p
�;G�F�J�e�G,h�7�7�]	�#�\�{�.���֭Y��
/�������}tt���Ղ��~��g�A��I��;��^g�W�q�}��M���XlxVHYEB     400      c09�,���谕�^��7�P|�e�"�K1��f��ԏ�� �-ã���^"e�ۻ����bA-~�5t����ݼ��9U��N.?�ur�뎚!]�>�PFNiYD�G2EŶ 6O.�Xc��h�����ܮ�o� �xԚc8��`e��׃��uD�G��i̇�dv7���W�D*^7cDn%;�����w�XlxVHYEB     400     100��l�˰P�TU��/I��S&qJ��(Q��S(��f�β?�(�ҡ�f���=�=\č"��GN��������uS�qw�뇋�m�yB�eT!s����`'�'��y2��VA�n�n�F֐���9��7�t���t���Ht�r�U�RL��dJ>���F7�����y�&�m��>p0fxqEG�D���T���\l��~I��d�Ԑ��<�����J�[ ��n?������KW�֋�^�3�?XlxVHYEB     400     110�;(iNבl:�A���
Pj3t?{Ws����L�$O����H��v3�gUO�zb�V����(s���zZ
��;4�i��ňJ����H׌?�g.*��Z0JG�����A��nE������+��.�|q�.�0����_�"�����ۋ�C*�L�������~��{N ���[5Ƥ4f�B��Yi�[�	VpRʗ�A�@�����_�y�!����E���)�����|y����̂�mv?~v;Ȕ�2���n1��qc'Ә�W�C ,XlxVHYEB     400      a0�l�W��M	]¨\��?gȖ�ԨoQ������[��nb��C�`��pa������b����̂�vZ^�QL�K |��U8���J��h��@vFc�ۙ�ɫ�[��6m�ohl���c�ё�����$�8�Л���ȼ<򾁉oL�>
Q'���XlxVHYEB     400      e0�����7���L���/�| W���o�+���!����8ff��rkl k��%���fd�}��j����.�t����Tf�����!j0n2�k��F#tl�o�3�e�N�(��5�����.�Φ �ւ6T�I�esJ+z8�z�#�l��	�q�<o������X�ǗG�I��Iq��ό*MT��wՎ&�������M����5��b�v��y�>m[�XlxVHYEB     400     1a0Dc��k�d�`��>�+?���r{wG�/��{gx�,�U��)E����>��N<RF#�?���~���7/�&b��wv��i����N�ar��wp��\�Wa��Q�L��B�@����ʙ�1��$���&�h�s+ƿ
���dm(C)�:Y�Z�󹑼}�Q��SH3 �t_`�F����ϑI�-���B����l�c���b��*�(p�1��KC�;���"�`�f�l�Z}=lx�2T��� �i;��{q�t���b�2FgE���j'y[QMG(�'Y��D�������ǰ��2���rlDk��;z�I��΋J_Gǣ�:�۬L�݋������Z�^B]�!��2��a,,�i���7��b����q9tX��t�SB?X�el2�Ā�읯_��XlxVHYEB     400     150?�(YzаPQ�T*`ѣ��wL�lo�M�EG^m2���&෽�G�)� >�(
w�8L	����,؈� dK�֘����<���f�C�y�=3u��H,�S_�²G��2ه�!���"�����S�t���Q��x�)�_D�J\ީ�\E��4'���� W����������z�@�A��U�Y��o�O�(��CJ���?���R�Pe��3c��Mc��l��ۡ�;�"^!�'h ��'8-jV3���x����ͩǔ!/��{d�;�yТ���S��5��;z'�dMq8}I���M��tm�(�Ԕ1a�iw�NP�{���=��XlxVHYEB     400     120�c!�6�M����7]u@܆�|f,�"�z����#O2U����W"�䄐���X��d��!簝(���Kl�J~A�7V��|Gy�@�?�>\�#��9����=ë�Y�"R�d9�K�k1>�P-�S9)���/�ub�g-�}��I^��٪����M<�~S�Mޫ{催�t`D	�YF�KօE^p��N�=O�Ri��ζ�,�B�{�],�9�/96a����-*��;ű�&6:?yPs�Z��L8w���u%X&��ԀP�;�;#��D����[�K몚(�RXlxVHYEB     400     1d0�|�p�GN7��iw=��z�ƕ��h������6�"L͎X�a��ոd�%��;�C�G�RM����	؏���;k��wg7hC�Y����ON|�Ɵ\#��|��������$~F=DClx�X��5��{�~�}qM=����e8�A�6��9hD����	L<�3TD�p��;�u�aL0� �-��u{O���WW�C4<���������� �^k�:z܂D!������;�2�B �T�>,wWU�j�۾��>�'��,aT����%�����h[4 41�SƵ^_��" �����y<7��J't=��Z<�Ia��ˢ�УC��|\T�X�#�A-G ��>.-�w���k���0������"Y���H�UŶ���O�M��5�w���`�˘��(0�o��>n���Np�6ZǠ,+n�Вv��e���Wk���(���N1�|!���4�.XlxVHYEB     400     120:	��w��8��M3���-ڣ�����u��z��(Q���٢�B|�B��@{4��
�M�
	UA����-�ͻA�`��^	g�5}cԬL������\&��]�����=�����5�q^܋�o��0���@��O�:כ
����P��4T�: �$s�{�����7M5�^ `; ����q���}U�Ke�� C��emc���Ge/�ZFi� ��`QT4�7O?���aML��|�h6-�^�L�`���Y�{	z-�l�ͬ�^˔��=Q���XlxVHYEB     400     100�l�H�3��2�=����.�@|�:�6��u�c������t'���~�N8;�Ev�]�L�n5h'���bR�����%Z"R��_�^a��`m9#]�lsq��:�lIm��8��3D�S#F��/�~B���)e���q�%���X*���Q��j)׬�}g�|+A4;�yG1ӽZ0u�
�#r��#{�o���3V˜2-�Ӣ'��zX��������B�z0K<�9�,�kD'߷�W-����k��\wE#DXlxVHYEB     400     110+3�TB$��ɵ���zk�U3�o�-S%X�3E5���7�&GM��G 'yvWE�B�ޡ�+d:/vm�p�٥���Ty7g5�nA�6���!)�<��9n <�y��!���&�����3TZ�2[��Yĸ�b{�����u�K��_�V�4Uŏ��+�EO��X���$�]�-�zɘ�P5�(�F��������4%U�ǭ��Q�Ѓ��ݽ�̟�E��Ra����NR`~��Ɂ�eq"s(�o|_q��;�=�>�#��A�XlxVHYEB     400      d08>'��Q��.qN/1ל�rͼ��`�������8������)��-"|�W�9��	؍���LHN���Tc�m�W	����g���WvO�Sd���d��&��./ۄ+��M���v��Ƅ����0��~ Q���m��_�޶���_�V]��0z|14��b�/?����X}p���]2����e���P?���XlxVHYEB     400     100'm�`@xѲ7!�߉�pIU;G��~U�eP�~��ۜ�G�
�s��7��G���s��cn�],�k-w +�\I��U�ЦU�G�h Iա^�Ǹ2�.���
����<�%���;���(��L��Qi�x���*~������r�_0t������܄)/-��Kd�����N<w�}b�+�(2�+p�t0���9TZ���)#��w��`L=GB�,��G��]te4�Y���%��GXP`�j�;XlxVHYEB     400     130��VW]��A�6Y9a�=��3⛆]@7ΰ�Z�=9o�}�x��]�3{��I�����B�8����e��:���J.0*�`��[���v�}�]�|�ڂ����y�A8Tz�q����s�C���)9�5u2"�u�9�}�������1iz�t��z4�4��j��7�yQu{�~`�R���pN_����틞Z�c��KM;6�TG��"�����I�0�����?�Y6�ⶺ M��@o�~��i��!q�>��~�RV�k7�ĺD�^�Y�Ľx�&)��N�	��Ř ��2�XlxVHYEB     400     120Rv�#k|�6� �~����D@������B��12#��	�I�T�I�t�������#�,*b���O=�-�d䘜VՔ���s���� A�mJ��$"�z�a�h�����0oR�$��z�,�;��O����96Edf#�O�O�2�L��	ܫ����s�B��L�D�B�9�v�;�������Kt������*aǄ�S�������B�
���j7� �	�бV--�͊ä^�l��>v�����4�jOn�����VV2�W����N �a�p�XlxVHYEB     400     150D�HCN�_%���(4�+���-AO�k�+;�%E��� ���G�Q���e�X]F���"yТG�W�LP,+<��C?����)/y]�Ǥ��G��b�t(G8��l��~��l�P��rB>�Ra�k��T��Ԙ������������Omau��r��୎3���5�p�,H�`k����I�o;������m���'@(Ëj	�-���[R��%Y����DY��i�`Q�cA�>����.)����ߖ�W0d�k� ����P��Z����p�3��d�
�ζ[my2�>�8n�Z
���ޕZ>\�Rx���;��%R�kJ�P��@�XlxVHYEB     400     110�^>�d&Ad�Z ዽ������v��a<Ϸ�X8@�r	&��F�.$B�0+t`�y�d�_�`'����)���hh��AѢ��l��N(濊�������[;�@����~GnE���i*OR�k�7}�?"����l�v��˥�*d���?�s<�˔����M�I�oݥ`��蒪������".5ks�f�)��e}2h]ή���Ͳ�PF��z��As����5/�0Ɲ��ۨxߪy�A{1��$�݉��"��	��qXlxVHYEB     400     110��c�I�,^������s95��2�}�A���!ݶ7)���s!M�m��:�o�0�uE-=	{ <�Q�q�g0��$/=�Z�xa�j,[FʼP�
waW�__��?���%��)ba�J��MR0:N(��(��R�Ȍ�KK���}lQ��R:��x�[9L�<>�������[vr��7O�5�,�#l5_	A8DeW���.W�Y��B��́�M��C��7sD�K�]����
-�q>�A�&�I=���	���6[CXlxVHYEB     400     120�'�}��|�o���Y� �T��Zr���*=�R))��Õ#�]��̅��d<�	 0�^���OE+�	5ܮۙ�ߗ�BY�+ƻH���>q�i�5��qT�^TG���>蝬8˷��6ƙW�2�#ʸqk�T
֑���gE����ٽ��0Y��惑�;��"�D�ϥ���-u)�Ұ&5[4�8^�ɿn���s֟��k������r)��o���YQ��@v�`�I��4J=�Dw�Jc�P�ml\��^O��z33G�?&�{{X��l�xXn4�ȇ��ٯ�XlxVHYEB     400     100+!o׾w���Ux�Ù՜�H��)�w�5w�m�KN˃�&' ����دW�P8����/�W���Wh�m��Vp�ێ��P���va1��Ո�a��xd����/G�Cy���0ʣm�'�n�#a�!�&�j��NJ|�k*�@>S����E�t0�H��P��dUq�)8|
P� ��t�`��-ZkR���]�=�kc��*H���k���_����xd?fy�q�X<O��r��8���m�s�YϾ�!�XlxVHYEB     400      f0� �s\��z�����y�|�`�G:D̃C�b��GV����,G+\46����e%6��e��]�-F�n��h`�7�!I�z�����Ec�j$��~JLopf�Q{�<��t������<{DpQZ���W�0�6D��}�?*��5�OI�|���L~CW�E�S5��d�F(���J�!d%���c&f�V�Y���Z����/gr����_��"�&�p(�59wKbVM7�����XlxVHYEB     400     120i<i�DC;;1�$��s<����d(%I��W8W�|���.6y�P&"_U���c�,bʹ����YAQ��싳�e�\f��c�2��-1U�����p	��q��.�!8 h�+�qC�3%�k�X~}����gO��ҍ^n����1b���xT�Ӭ 9�,4)dͨ-��2(�$	�(�D��\st��4ɓj���՗^E�#H��έ��x�(r�[Ŏ�U<h�Λ안B*-~2�żj�vm�)��I���k�����d]��0H=��vs���V��	�Z2�v�$XlxVHYEB     400     110'�0�5��Z�<������u3�������z����=�M�3O&��H���4��8�_�QKx�E�)�0���lfB���LL"&h,���R1'�����UK	����WM�8��~}Ds�p^fʍ����}���a�,8�=}F�߀����wW*��&���¡�u�4��箔����i)�sx�&��\�x�I �$V��N8O�"=����B
�95�f�@m��ũ=���8Ǽ}J�1�:b��w�jNX�uZ��G>rV$��z��XlxVHYEB     400     120���'j�4D���P�G�]������s���Hw�b9R���� BjΓT�)�2J���w"��(��|^L�O�!�ea�ib�e�����S�Sᢀ쩆�v�KÍ;xE�:�i�CJ$y�3�i�6l��o�|k+�Y8x4�t�4M�nQ4.�aC$L$9ݠ��I�!��${sz��خǟ8�
�Z�l�dS ��Y[��&U����Wf`�1�z��1�{h�❎��e�����y�r�r#q׎�N:��(.cQ�s�u7ٮ��bP�q�1�Y�"��XlxVHYEB     400     140�i���k�(�˝<n�׽k�2p=@u��?���2;Qe%L���0L�dGNы��ʉ$Z���@A��d��59q�D�H�1���T5���6: �mأ8���s;�J
�IW) ħ�����S���5�P\Dޗ6���p���o)"�ojz~��-�V��Ɯ��--�J7�9�`���4Zu�� ��ӓ?������;/V�9�md�^�{28���Տ�C�J�:����Ε>�@�C��K�ｸ�A'�;�����1t�ꌤ��5V&;!d�%rj~a�݊����l^���u[��U��bF���'�v�xE��$�V�XlxVHYEB     400     140�t��R>��H3�w���kN7�D�o/f�ցY?C8���j@�� �,�� �4�l5(���>|�Ig�pd�ǝ�W_����@��㶮�q��X�h�X����
�Z'�@�Y��Q~9+�{������ ���!g3/q`��D��j�:e�2y� -�^SD�6��Z�D�^��&)</$o��[�"��� �&����-�W����Lk��)lׂ��k�`ж1-}#vi҆+���)qb�iV-KY�#G�7�'���1�㱣[�AĹ.Cɯ��_�0^D��!m|�����x�q@#=/8�A��3��� 2��T8*�����XlxVHYEB     400      e0}L���ָn��%C@�"�U�Qm�W�h��s�����͎�eEX�#C�t� .+���Y#&H��'V�2FN^t֭�g���=ц��ۃ�����̾G}E�������}yiȺKK����~��s� ��/�Ǽ�R�`sF��.�=�;rb�	Ė�~iW=����<�9�p@n�)y%�����V�i�Iz��?
 ��W�Ї��� ��0d������i���K|XlxVHYEB     400     140$]R������ �����**�ٸ�_�����'Χ{�\�2Kk����~'�+�2�]��7&�ؼ Z�J���*��呞d��`Ԙ�?�RP��ܭ�t�&n�(US��Vp�g��4ճ|���Q`����U��7w��^�P�Y,�v�jTt,e��Z��uWj'�a=�*�m^S�Su�!�F�Heq��d�����<b��=.S[�峀rT��?��+�E��vݨ��G�ZY�e��ka0ET�d�����BI�U5�i-�Q�N=P�{Dʝ���L	�����Иtmp}���sSq����*�Rvⲟ �����J▉XlxVHYEB     400      e0C8y����L�rX��tE����^�g��ױ\,hأ�M�z�U~ �|��b�H��o.����T�F�}�ԐWn�����z#>5�μ��PY���������d��$��t�?�i�c
Ϡ	��>�l����[[�/��GlHs|H���'��֘�b��6�c��oK���:Dy���U�;	�B
�@�ͺ��!
�;I�Xf�t��9����=&gК���+�XlxVHYEB     400     190��VdI{�ϭ��o
�\���o��G�fG]}�oW��e�Ɣ�ڞ���<:��"S|-�RƶH�&/�qiԅ�p��7\83H��p��Oz�"(r�!��7��;-�m�˳�c#f���B����ˁ���DEv��ITUn⃜�&"j ͉�[�/�����$�{��$4`94�r=�{ײ��]��"��bܻ��
��^����m��-�_�X=�ކ[:�wy%|��KP��=�䦠���E��l�A��%��ŵ�\$i����eb�Hzh������^E�)��ԒJ	��W� �\�!�� R_Wd�~���Z�c���e��Q��`"�Gv��ky1/�`e0��PZH�1�V���x��Üfw�Vt��p��v�n[��n��εXlxVHYEB     400      f0��2)F���,����/��j�6�E_İoO�3����	�&?h���>6KY�[�U����
����.��T
"���C����������~�����7qC�x�Pg.X1�g��4��	�(r ���f�u3���P�0�<H�	>��i� �`�F���@�x̂W�&�c1��ˏ�u�kFlH�)ӥ	�0��U�[۪��v��&�n+VA����U��ī�Q���j�_�����6�XlxVHYEB     400     120U���$7K+"�ȼ�� ``��d%����!�
m�z��Db-�&T���_CM=�uim}a\v�:e�Vq� ��( 
�Lk�Z��LZ�ng>y�#��a�7��Aa�N��o����`�*�a%�pJ����R���v{�����wLGd�pHi<Gs�gL?�yƂZ�R;�f�U=���FZ3�t0a���15�"{�)!`�������|ܼ�0�x����$��BbF�R��o����_0]�js���]���V��O�8��	b5J�O�t��4ҏHG���J�]]X}�{��&j�MXlxVHYEB     400      d0C�&�		�r��od��EE�-;p�y!�6q��DH�A�_�.�-0���gkTYw3�t�G��i����΅Rl�͙b��}��,I�6��<�~8��.h�g��i���r��z"��}���4��h傧Q�[��s�>�����t���E�Ӵ��qT�b#���G��[1`��$��
6�>yV�P�Y��V4��-2,�A��XlxVHYEB     400     150G�{�����W�J�d��["���Ԗ��CͲ\J��Y�M;���_���$�h�H��C�rь�����v�*5�K�VJ
J�ֶC����dC�2$.y�'^�B�Yn��t#Z	�0����(hnߪF�	�����~w;C	�t�F�� �ޘ�Cya@�s+4����f붵U��wHH%z�L��Иw8��J'����d;�]$������P�Nỷ������6Jw�'�Ѵ_}潫g��[�c"�%�O5�h�gh�1,ߙ���Z��L�4���=G�^� ��Հ�x�Y�0���h�}K:+]���|�ZY=�e�3uޱ�G�eܯ�Y�o�"x�>Ħ�XlxVHYEB     400     180�-�b. �d�����i�C������G�:��HW�_���2F*��ilP�Й+�`��j��g���D�>�s����:]�ᡑ!��#垟|&+��76�<����=.ЃP�mY�8�U�K��� cÕ�j��g��zG����s	GՏl�鰻�!�TwJ�C���c�@�H3]�3�{ˣ���`w����et�����J��!;�^t��/ �=���iC���Ar|x�`m���ްHa�3�I����<�pQ��i������o�pC��w�Y�Mj�^'�?.��u��gUf�U�/�{����eO}��l�.r�F��:$cU�^�����ެ-7���S�?g}�?:kn���L�}]��BېŢ%e�p�1�m��X�_V�XlxVHYEB     400     120���{ ���O}�QֶIz��2l�#M����]+��-�b!��9:�����_Gk1ΫA;�LB��~���R�r��K�#y��`xeB��yc�%5�u�f��}��i�1�.��R
Ed�y�mihB �k�5���tʬ�f5��
G��*�"�n��j��!D�k��*��&�2Y�+�h�=�x�o 4���W���ŷ��OY��T�,P̝����[D���[���Y���cZ^Veڧ�-�[b��7"���Re�r�X�_��g��(~ͮ|8���vL�}����EŘ`��@�XlxVHYEB     400     180?Y
�����b���}�����n��a�����D��B6��2бd`�oV�X�}�TY ��K�����ۮUa����/�J�x�����c��>�q��9=�a���BKۦ��Q��a�Mg���2�G$@�EU9�m(ԱG�J�^�P��[���`0H����M$��H�������P|~j�?􍥴 � #��GfzX���%/87�b=$������L�9'��dQYMϥ5L�B��,P��z_3 ע㒝03ڏ-��q�5��g �ٺ���Gn������끐�u�j�U���yBGnL�7Vcj� V���� ��u�+�c�GE'�7_�⫷֕��,n��ܣ�����,��ze�ժ��:�0���W^XlxVHYEB     400     120��ވ�$�@Ю?�M�>[ϖS���������s�*�5����K�
{D�H��(B�:�WUA,����ӷ}nʏӪm.?�,�����F�����k
z�UF�o-W=��[�Q���,I�>s�3M�>����� ����w.C��MQ0����'�Z��R�1N�l�����lƻ� 0�ӵ�Kф��c	�����˅\{,
VÙ��O퓹h���z�~< :�rM�t]C'��|�t�\�&SO�El��Q���ޙo�Ҕ�����M+�������>�r�t�?�ZXlxVHYEB     400      f0E�"z����`���ݟm�gÅ"87{��Q��r}�yJQI��g`�6��z��#Xx��^
��9������=nh�#��;�[��ʮ�NX�����n�bI�~?�>�OgK�Sƫm͚N7��!ude�ꋳ���c[���:�X�3ݶ�J8iSM�|��пY��k*�L��lH�}X�ЪB�
}1�7�o��,�as=��In�Nnmj���/�݌A9mg�M?�p���{�1��XlxVHYEB     400     130�,��_)�d���%М��=BN��XJqM^�>���Z���݈�?�E�����s�J�-�����EJib�P�{⽵6�OKT���m��'�a�z9��5)n���J�0�U*�D}�_L�	~�a �޲@1": ���y�3�����ܓ�v��ޫ��ϐ��o�\�����-��[�bQ�$pBz�	ee�VŨ��nq��ӿg���&�d���Ub�'������� ����"��^��Y���8��)������1��4WG�T�l��0��:��?nd)���_���W�ﮨ��eXlxVHYEB     400     140�zq��A�쿔�bMH�M%�ֶ^��X�k��V*��T[}#���v���R*�SMʹ4&�tSƯk�ݧ���$��v���>�-�öƶ��H2�f��ӴϦ��W��Cm�Q�S@X�'�Q���v c˄@V䄀���&M��}�1�I��YE0����&�9��yY!�5�G���Y��IN�������cz�A�����5g�B�R4��	u��w�G�C~���P�*Z�#]���r���Uy7�.�-B�����P\��EXf�!���`)_�c7"󎡅s(XF�r
֞)���2B�XlxVHYEB     400     140�<V���� ��a�l 848�"��xOs'/.	C��i {�������׊MLz���5^o���ǩׇ�8Bڿ�mj����5�|�d�O�#�;RE��J#1�R�Y���s	���4����|���nВ����dB�u����Y�¾�w��'׸�mμ EUB�/�I�w���y��N��=�{���e3���?��i�T��9�E�W�F�b�$-{�[6x�F��"KxC����V(��,ٱ���C�.���C5gj��;.S,��[B��I���$M6�I��LW�#�0X?`z�Q�i�����eoXlxVHYEB     400      f0����(����G�T�ñ�'A`��ɓYb[w��B�B��&���;M�u�AyK5�~��]h8��h��x:5���~ӔDnմA�@����V6����k�X	H��uy�ə��G	�G�\}����]C/C��낑��I^�B��e��P�H�O�E
����s���3����ٕ�A�]]?H$wq�T����C�i�M�腒)8�e��!���, �%�܊dYf
�b��E^��w��XlxVHYEB     400     140?4�?�h\��c����.X�G�P5#�����	I��W��S�-ؤ�N���-����?Έ
7؃,g]�����T"ܓ}�;;.]4�Z���,�c9�p1A��	�o����L��ҲG]3S1��m����JՁ�����56�:��e��kr��w�WحnQ� 0g@isdÿ*[T������G�^�����I����N5	sHF��Vi�YL߀��Rوd�^����`��\�U�.;�k`�="Wz��;1�U�~uN�Ƴ��M����/-�%�B�5��M��P�վ���.���Ε�p����kP`����.�_)XlxVHYEB     400     120Ϫ��qS��I@�W�dÝ���I�$3�޿iV��"��J��<̎����4�r<xBIl��#]�~#J\&I��ס��r�}آ�?D>���<Z{Z>C���/�~�Σ��K�F���3y0c�`�J��${�V�� ~B�)b�B��Y��Q�ܦ�qp�&�]���E��v,�����c37j=`I[�"�ú��=\��q1>��`��t���l�� �a�@�t�sS~��R��ۈ?��LO�G��BJ4G�	��+T����L�^�%�y�*{��-�UZ��Ga��f"XlxVHYEB     400     120?�N�Z�T��.��I��+��n��ҒQq��o½�!q�|9_�C�>���I���(#�搈&5-�G�G�W^�S��͊9�,�&U_�_ߊ�޹=�5v�v�u��2[<�ܩ[n�C�DC�lE���&r*�"��k;� �q������t��!�i~��&����j�6r�,=q(1�L�Z�����j0�+!����k[fXKW����E���f�(d� ���݅b������p����u7z��a#�>@�w�m�zՊ_�x�Î���l$�XlxVHYEB     400     110�1/�T�˧P~�5�9��w�J���k���Uu|�5����/�G�Igߌ7�y~��I&���t�@i#	 ��ێ�����L8ס�"�X3E<0����6hH5������p�l���-�WY�-t�4oG�1�_�}�d=�V,�����g�
(�|�?�	����\�!�noVC�����Q�^�!g�#�­�vQ�Σ�cې�%Lo忝/�)M,4$���W��p+ߑ����x�\�(ȭ��*��*�J��zMXlxVHYEB     400     160[��`"Ȧ�ywy������Y�`�^@q�u>���h!����&{D�d�qx0��&�Z+i��|�EE7L��i�0j�h���Ad��y��,�,7R����m�#���)�o�R�7�ҬY����
w�����
:�f,�F�#��zl��b�� �����	PX��G��r2���u�EFD3��i(&���'Ϟr:E�I�F��5q��=�iZ��������aT8���^u�&����E��/�Ϋ�^6ׯǡ�+�v*C�ə�����X����G�A�9�VC�q/��~o�r.i�{�c�֊˧�X�@��WG���fN׏Z9��M�+B23,�1SXlxVHYEB     400     130��
¤��~�|�_����l�ś�Q����Yɒ}(�i.�wh�w�����c&E�n����>2�[L-ͣ2ţ�y����8:t�����`��R.�\�W�����\��g��p�H���r��Q�\#�*R6/#=��?U���DҦ�%G5��w�E�S�<?�b��	�H�y��mʑ��6�0�W��-sW�"qHq�D����o�n:��3(�FD���f�6��������qG�����u��	�Ǘ:7�?疹�Mkd��2{)/�\��K�n(�B4�ʁK�Q�H���~e04j���XlxVHYEB     400      c0�M0�[�����%&���2RB���}�=I�&���GB�@�Oԣ�|&�s%̤����z��C�-?i��?��^�hEfLm�ۛ�ti�Ez�]K��1qBZ]�#��/}F�!bp�ΊwWj�D4 �o�?%�KR�e���������T��f��h ����	����/^\ '��y���/���!1XlxVHYEB     400     1405�Q �g!���(���>�䓉�\���M8���D��u�1)��O�X ���V��D�%���ę�Wݹ�iT�J�Xh%�B�O�,B���v����i2.�v�չ.G��d^�V���m+�
�̄-+|�Q�S3LZF�ߒ�^�č�X��@���N�{�[��z��գ�	f1�k-�3$!����k;N���T��z�H79~��&&���M�^m����F�g��1���$3ɧ"���P��_��U�ynt��Խ��.�b��V����1d���%b[�I�� �gq���e`�B�ͻ��ji��hꖵYXlxVHYEB     338     100)^��᪓��Vq�`in�
�0_޿�Y}W�X�dQ�i�W�||`����NǿX��fk���%��FPh�7�B���1�������I<x�m%�I��B�=��$2 �{؆4��ͮ�~��#��ԧE�X�Z��A��flݵٔ�W��??֣8M���py��X�qI��@�wrl�&�%��]�����������M!(��:@4���n���4o?�e���|Sz5<1��m*��D�k	|V�~��%-�5�(�