XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����oU���`���^���m߉ﱍtޱ�
��e���f�{��hA (�u>��߳���AA'v�@���V��C��������Rȟ��پ�.������g�������M�;+;��P}����Z���z\���^'�n- ������P�C�����z��CE�������<���'��)��s�����F)݇��z�;7��X-��g�E�n�uu���܄q�Fq�W��1���[\,8� ���s������yy#�]RM�F���+�k`�-;^q�@���c#-��Suy,x�VA�fa�C3ͷs�{�4�+H.Ŀ�K��%��;�HC ,�v�O�K)��~c����?.F�M�� �h��#��7
J��ZE�yo�>���Or���?���B����C�ABR%�c%�{-�Tm5"��'Ώ��Z��B�dn}�d�Ԅ��R�'b��0��K3 ��	_^��9����u�;����\�z����D�� K��O�tϫJ���G�)��q�fQl����,����a/jG�(����n2N�V���!6�}��
(1|M�'Z��B���
��������;k��:̮�#Ȥ*�Ӥ���"ĥ�/��t�-����ز>�Cd^x��,L�}�^׃U�w��7��$�Bbƛ6OI(͓[�q.�O�@���7*3W���|%Wy��
W
B�9\.�3�R�*�����#a�uJ��߉o���N<R�TΘ���/�ֺ��yϩ��S4	N|&��XlxVHYEB     400     220��נ�,LU-�	E��^��[�vSŶ_񕁘��jb�_�D.AQ̷��I��38�u�Ote�ɴ͵�d�(�$5�#�ɳXQ�a^̥�,ϐ�6��H1�Ŭ��R�IS�`rҼ��3���A������Z��#�Ս�{���#t]��6���]�[��nY�}�~�o�B%��s�� \���
�Ra�����y�n�&�����	'��l��)�C�⊉,��#�(�I9��4��{8�X+�L �1g���@���(���w��?�g��Y�?�(h ������Xo�*�$�D�.��e	���"+۠\��[S��o�vs���f͔��w,'�A1��bkq*)d�5X�3�����,� .pIjw�db&?�E����y�3N�
E�6�\��|�(fi�����i� :~�JToe�|���U�v���'��-,�>�ð�i��_����+Ou�J&���s'!��=~��or`��6.A^u�&6m�2!_]�V���e1����G�)Q�[�7�P3��Vh�XlxVHYEB     400      d0�:��oMp�<lf������c%{n��-D�&�l��A�lR�8��}��3���m�Xw����-�7f�]�Mi��Ph<����u���V4u�M7ڊ�$��(*r�W3�5D#���7��Ӊ�8í��>�2l�?Ys�� �Ts��'�8���QG�֑I|B�c�k�<��d�A�2+!�+�uģ���N�_��y�oz��2���Vj�נ�~(XlxVHYEB     400      c0���:ck���?ry���c���>�܉�PVy?��+��&��q=?�V0B@��^P�P��K�
�|�l;�H_�7X�"�`B#�̠V���R�"6�``	����U��<v(��?0�񳓓%&]��e����7n7���T-��s��G\�?��� �H����m	�4����YĻE�a��W�ߟ:+��&RXlxVHYEB     400      c0H��R�l4No����Nr���6�yFĎyu�3����)WA���Rnԋ6�@u��y-Ts�O<�n:����㵛R[&�����M@�a�]���5K��R�mnRna^X�M��=ɵ���@0��>x����#(:�+}�Π=�F
��Oyv��q<X��s�)�/?V��x���Y7�;��(�r�1����XlxVHYEB     400      d0�-O�]�YJ�/N)��d�.�B>	w�ލEԂɘ�7���"+2�\[�n�JK�ki̹/�y����m�?��5�e/OKx��c1
�sb�h�D�H�d��^|�M��i���Z(*�&,K���~�h����f߯T�+V7��/vɏUv��O��gj�ֳ�����=��#��
~���U2�z�tRb���lj+Ӟu�XlxVHYEB     400      d0g(�8՝�x7�4��TOa<f�>�ÌkwɠD3�X ~x޵۷8�m�-2rm��/-Љ�x��bV/; ��� ��t�e���oB���>�s�
Mk6H���<a�G��.:0/���;��6�Aw�;�m�l1���0�i�h��>�\ר���=�fx�n�Xr����5@�h�;f;�������7;�6�Mk=���A��XlxVHYEB     400      d0�*}��/u�|�f�����j�X����=4ֹ��v��\'�lW������I�@�7Z��9�,-Q>ԑ�}֨���z�����շ(^�I���l{(���!���E]��z� ���I9g�fG7ϬP��jw�/˺5�;��!�U2;����E!`'n���qɘ;v>����*�����6�$	���+�G���D�}���5XlxVHYEB     400     170�U� �foV��-�-K�{���jƱ�~߷�^���

C6�̊Y.O_Mubw�9���L�ok���~�
�����y7�	Q'��u��RpC�R��g���rZ�ƚ�*��2�]Cb�誨8������1�Hr��B�����m�Wo���D�	彦�y��곈��?�<@ݝ(@NwAK�Gl�&�C�/���'���$~º�9�_�������L�i����r��gm��P�oD���[�}��1��UU��H��sJ|fݻ1軾w��@kᗣ,����U��*�	/���%�"y���ه ��֙��VM�ǑH�@}���S֥R߭�-Ʈ�6pX�� 0D��D���������XlxVHYEB     400     140��֟�#+	f�_�>�K�%�9�㋛9�Q�tAo1J�ThW[x��>:I͡��5s�N��+��_��we��-#\��#KG[��S��Q������
���&\
�Ɯ�,SUU���f𯸇	�8�c�߉*M�0�HC�%I��}c�z3�E*�ɑyw�S�'���͕�/X�R��s�{�E�/�kq�$�u@N(�z�	�u}'Mb����.�>n>�k�TE��=�$��!S�p�� x���{�A�����x���b�W����Q�>ݭk�ߌ[xz�(@������Ny�g1�_fs�[u�Ə�~dP�l@��%�S�:LR
˓XlxVHYEB     400      f0�����^���o{�d�D�8|�.z��x	�sK"��`�ᕐ=�H�ې�ʣ�_14����cu(��U0�wp���0W$J],�]Ԁ����2��)/�ɑX�C���Ji��HN" �=<o�5��H�yk��/KmBf�
9�M����H�=S�iv��c���beoR���@�J�CXO5�֠W�f�P�0 Ț4߄Q8�x�r��ר�ǘ+t{���	Vm�~cJ��������,=�o�Q��pn�XlxVHYEB     400     100�����`r��o���}"_��j�ͬ�P�/��!�^
�>%&�L$F���Ӛ���W�ň�U�t�_��-<�3BP~�4;�1nǡs�x=�M��X�S��p�	�&Lk�i��]��y�yw����O�6NH�C.�YO�C3/S�5��ȶ�Wd/���Dvu-f�J�p)���<��&ed�Ѕ�Ḅ����21���*��w7���0X�DFpmڙ���@]��ը(��O,L����_)��6�<��XlxVHYEB     400     110���`���P��a�V҄��˓�Q׾_�IME��QU��fw�DM��|����
��V$�1� D-Jy9ϧ:��xB��w��&n�L%������:�ץw����.i���2�2~ΩRp�O[�)Lg$������M��7*UmY|	r��:�ί02@m���LU���QFZ�	�擹�B�����(�m3�J�~��$���lZ��i]�惘�h!2L� ��|�����OדY�uc��A?��Yz˔���##��}v�L��^9ǳ��&1��\�w�XlxVHYEB     400     110䌆�I�i~�ዑ[��V���ԑ���P-����&�z��qD�^��9 «�iBh�ǰy����K�����oVq^����-���Em�5g
8�~���?O(����X!���	�\��e�x���ӵJm�]"�����x���!z(��-�gF���6?����f�+/+A�����R��X�9��/�(��"�;� �=,�=j�/��6^ɕ�E��D��!Δ]�_������K� ��t��@�ha��02~��XlxVHYEB     400     130��"���rJ�����0��9�)�[�7#8rN�G����i!����#��;�\~���o�ÿ%�i�W�
�;��K��>����?�7����2T����ц���,U�Ћ��k��ֆ�u)A��S����G��^!m[$��1b��R-<�������)����|��<4��?a�iJ^g�b_����]�t�d�N�,jKp���7 F�U祙/mƝ|���L��; A)����+f_P�ow�[��Ȇ�q`Z͏�/Ο�X���zo&���}M�eHq�)7�bo �]�\߿�V�!�Oƪ��XlxVHYEB     400     100С�!v�T������U�X���1'����aJ���=v/�q�1h���z}���N}�%�R�������d�K�1�7I�wjKA���O��Tà!���!�U�� 5�Nk���ft�Lx�f{��h1�S=�I�!@hh]��.���Kf��z�O,�����e
!�\����!����n�����������(Ƶ`Hm�(�����b���g�Si�!����ָ���k�-�Ï^�8:�QO���P��I��5ӤXlxVHYEB     400     100���՝7
&��' �����~��Fk��ρ�O�7�鈯)i�eYc������(4���i��z�?�,�@�XK1�p�rKu0폄�x(g�FxP~X�YF�"�F8���5 ������2�j�b��в�qQz�*����aؽrkK%��]x�����VK����y����L����2b���bQR �}?;$��$�+�����0�0��H�Z��c�ϟj��u��1���THZ��"B�XlxVHYEB     400     100�)�vghK��#Iq.�k��`�����V �7��{�2�g�P�/�	�ލ!���Z�y�G"y�U##D��(.3E�z'��T2��
�
m%�9br��"k͹=�o�*@�p���}�p�%	����?}`���y�8I6^���?�t��W� ��I�À�
��f[&ݒ~?j��fm��m,��҈�z�I��+D<X��Q%@Y������8� @b�B(���o���~��M�R��/.�^�I�2yC����S��/���XlxVHYEB     400     100/'.�b%�5�h�	�����n��k��I�*�co 6[Tѻ�El
+TV������^˳'�:cv�q��wkG�X���վ�uZNs"?߁�>�F�&��B�͈��'���y5�a�BOߓ+�<�Y���);X��8�+d��6I#�t��id48�����}�P�gQ"iLu&���I�zߖ�0Jܬ+>0�� "Y��)K�1;���h�|�l���b�ߘj/܄-W�D�ʨ>�fg�,腥 _�M�J-h���XlxVHYEB     400     100��RJma�M���N�������!qGU�����)�O������$�	2�Ke9�vnۣKxt�#o
�d!��BܺE����iX��)NS3�PMb��,W�y�m�m-������w��AA�_j�L�S��+����" ��T�Z��=�p�`��ܮщ*@8�;T�Ӿrq	�q4�R�(��}{*�m��Uúk��͟
 �<�^��t�M�������NT;d��5���0KEP�,�XlxVHYEB     400     100�Q�/
g�k�{�Q~��Of�O �\K�(����b��Gk�������j���}���s�s1?�g�]^�&��J�h�	��ӻ�>�6qd�����Ԝ`m���R�L�7�ey[K�G�;�g�W8�ƶ��
h�	7^:{"P�_�̛{�t2Z>����Fz^t!3Q�o"��B��q85@��� �����pA:�q%�T�!���P(Dێ9�:�"�C�Y`�*��`��Y�Ԩ�h�&��ԣ$��XlxVHYEB     400     100���zχ��1�FtWLb �W��M�[��C<eL���1��!�uI��_Xp���_��G�(��O,|U�-��(�c]w(�!�:-�>?wE������U��/��1�R�|{��Z������ˊE�`=�F���n�z"��*%��\eu�a�k_
g�Oo'�	B���ퟯE�0{T��6CD⡟��-5��ÿ���;��z�OZ�m��-J��!��S��b�ߨے�N%l:R� ����l���lXlxVHYEB     400     100��Q� ������N����"��G��%���M"ފҭ*���/�>���z�M�0���`i��i2g�P~�>�OQۮu�7�qPW�Z]e�_�+�i��i��EI��92�~���t��26�
��i���~�`��
|}�$��@��I�Dߧ����2��dRᠯ�6�0�_�u��n�A���|5�p��B�>�g�#j��h\����.U�[k+�}��z��`G0�\G7�G����p��:N^�G[D���\XlxVHYEB     400     100^a����i�s���H`,�_���nb8��6�5���r��)�:2�m�
�RC�Rd	J���@��0�Tp���{�Pp���������(|�����(�lV�MV��X�����P\�`��?��}$x�:�'���ZS�9�sqv��m?K�ك0��p��v9AƾgB�����yg�L�@p����8ViHf���麁N�j�>��l��;ܙ0B�9��^��t �	��h+��rҎ�eh�.���u����IJOHXlxVHYEB     400     100�z�Ѝ��vn���2,{��Vo�Ȳ��C���
��fu�a�˄���Ն��d� WF5���U�?�|���s�%�<j���'E�pR�|�,��߈��_�@2mm���LDY]V�4�� �o��]sb(�W~/Gx:�>3@���Ļk�ծ,�H;S+g͗�O���
/ཱུY��o�0{�&�xhh9���/�I���
4k4���Pjb00�Ù;E%������5d��[��*��K F,��KUXlxVHYEB     400     100v[/;������Z�����ra�m��I��A?$���\Q0��5@IO��\�����VtTR-��e�1Y]��*�����PJ��ִM��vZbLxG~���:h�v2R3�:�B��F�0I�^�쀣��;)�3���hB,4r�4��� O�ZF��&�h��i�j�.S �`}��b�[&�Ǯ��{�^Tp�ʁ���׶��i��c%��G�E WH�&`�t) �|��Ѓ|k�D�##��o9Wj��EXlxVHYEB     400     100'ҫud�����\/�5yE^c����[�4�R���4#�r��_m������O�6g��e��?V�+`�H�12q$��d�M��	l@0z}�������	 z�mN]{]�0��gc��U$�+JM"�ڀ�'4C{���5�&�D��9�V��4Nh�[��$�����ޠ��+�vo���4m�$��H��NS~JK�'��ݗp����N����ۄ�IN�Lb2���}[�0:�r}#� Y�FY����dq��WXlxVHYEB     400     100q<U,IyQ&S~ʱ�����\>��G���Mx_����j��S��B.4PD�<�&����`��Ѐ`�����+{_�����z�$�*��bT��������6�r�ڡ���CM-�_��W��_]��)�
Q�8�W>ek\��A���R���;��L08x]����͛w��d+��$�?ݧ��ڕ���/0�B�"2P��}��n8��-=����=-��`[P�먢�����-���(�z��b��XlxVHYEB     400     100��$G�H�lCi��/���s�/$�5훹]���Y����_wh��%��~�b�i�b:f6x�e��}��h~Jf��T��5	v��*���vX��r��*�}���*Ÿ-!�Lqe��Z��[�|�H[�B2�W4��r�h~�ʾ!�RǱn>�p��F;7�^ �vU��I�z�	� �&�ן��$���9v��wӏb��W�>Ƴ������0t�-���"����>����yB�
uKUH_x ����Q�XlxVHYEB     400     100�&]��Zv�!�PVT�wW��F�&���;E��h2�g�fq��5k��K�
ɓ�,R��ĩlk�9�oai7�~(�v(�`�A��Ҽ����.�s?_�z8΅\yqa����4`6Q%J=�;TqX�&�Մ�>�6��h�H�&�t�Vb2,ny�]\�û� �|�
>
sW�IKy��E��'�� o5J��������kY}I�6�.S!6Z|Y���ٛ���7 D�Я 7C`�Kf}�^�ޥ���'P&XlxVHYEB     400     170�%�����OJvHB�8��˄aP�_�$�*R<�*�ͥ'��\�-`�k$k��T���%5�Ne��G�}f)��sb�A�u6}�d�9B�^�d��vP5����y�*��~� V�N���<��� _��
_r~G���9fHЧ*�\(�?.\��l�v�s�k�<>���ӻIPl��S�*(ͣ�).���]A�ۥ���eSA���巟L�v;|0]_�`Q����EÓ-2f�Uj���Sƶ E�6up.��C��w��-�N�}��\��.�vhYt<%v��%���D`\� ����Mp�h74EdP|��4���˥}ȔTN6�j㍩����X��2�Z؇��>bS�Ӹ���d
�'XlxVHYEB     400     100)0����-��SURs~�*��7�:0��p��k�#{�q|6�J������y���vD3��P֑�B�n�U���s�����>��`<��R��Щ��	��5�&���U[t뻹mO�N��,��K�9���NUbI�2���һ�Jt)�`=D�8�Z�{���'�m��G;!����da��B��y��N���;�}|�"�/RB����q��rYkjmIu�_W@���Ey��A���G�����򿈐�L�XlxVHYEB     400      c0��Oc=::1��ӹ�/gXkc\�KUR�)�V���9QO��Gh��YF��!s��#��甓��x~� �&!���H���W�W�'�[H�59�&�8����4gy�a��1V�<�>��zP����m%52$������P5A��m9,��r�m��!����a�;Z�8>��*-l�����X�<{�/��Z�-
_�hTyXlxVHYEB     400      b0��E&��r��p��e��ς�Fԭ�R����@�A���]iz��H-������S����C�n�J���$��`�X1Љ!f�c9g�d�^�`/���ӏn�J���jV���z��f���q�[�-��sM��p�u�'a�Kv�8Xc_�s�^]1�B��4��$.>1�;0�XlxVHYEB     400      90 �6�>��E�o�,m�Ҟ��C��s ��:1|W)8�[�K*��8 @%��f�����b9<?ń��AfAI��aj�2��{ŰdC���=�9��o�p��]*��
ר{dnl�
�i�:��2�!�l�v0��p˻z����M����XlxVHYEB     400      90�Skpl�����P�Lv��⿷wYm:?�-È�!4�,�{���&��j�m�,˕�_���'|�z�l�{.�y���hȼ�Oya�IB6�9�q�����WN�s$??Fo��I�RZ�*m?����;w��@yN�8XlxVHYEB     400      90��8gA� 3��ȑ�t���n�����t�*�0�x��Z�ʎ�0���u���, F��Q
��h���
/,(����w��R��F�HW?�
[�Z���=6-@l�R�',�پ��r�p�mJr�Y�L������-:��7haCXlxVHYEB     400      90�.GS���հ�*�	Y�Zc2�~��T���,<�����Q����%� WJӖ!<��6�]\#v��WF�LR�r�6lT�*�]��>n�e���
Q<�2���hA*�G��x@��RW֚$	r<�=��Y�S�W�)�EXlxVHYEB     400      90 C��?#E��ݠ�E���,{c���H��[���X.��-��	�/��|)�)�m�Fڤ���l���hEr�Q���$ii�5�<Q���UmL x�i�V�
�	�S�z�P�'�F�;��W�^�=�\�4�XlxVHYEB     400      d0�9�\P�W��͸����X�-V%���	CĒF_�xh�<lw�G�K�y��i���P�D���p����(�X�a��L�sPo.�׹�����B�lnnz���G�A&��8D_��OՒ:���U���'��/%���B�d(T��r�n��/���S���{[]V��tK��ٷ�{��`�D�S|�07<V��D�h����t����ύz��+`aXlxVHYEB     400      e0 �#�1|2��ѧ,�^�D��t�=�2P�h�h3�RP�n�tc���K�ъ�ejޡϹ�%��G��Gg"4LE���ow)�c�L�U���c��e=�N��M~��.�9��r�*��yQrt&hD�^��%��:� �������G�1���Ң�Z��*��y�����+�����J�R�L 8y�x����G{��-~�y�儒����İ3�V�sܾ�'�XlxVHYEB     400     100��(�>�r�wR���vs�vaz�eџ#���2�eO� 6H�wߕe/���x���FH|ϠJ0�g�]��H�}�f ~��P�-���\�O�k0㨅FOFv�	P(�D�YRZ�?��&����.�Bq��?U
0��"�����6^|A����n�j�N�����|Jv�#F`0!��{8P9 Wj�O�8fAPͭ���Gl����x���%q�$?��a8F����*I)R�a���L����hb�.�ٝ�o L����XlxVHYEB     400     160\�&8�=xX��Y���P�M�W��o�3䮲ڨ�2� ����^#�iCy51�T$�����*{򯿖O{��#P"&7�k����B/<��.f�J ��ՏK�g�W9CY[Z�?Za龰:�\��x{I�฻�����2C����2���y�AGT0�^���Se�a��4f�V9v/�+q,����r�Q���T����p���1��I��ӛ���FŶǙ�`)��Zx���gݤ��!�h7-�-�Q̽	��� ��x�H���|mL���;�wCB	�K4�	%8��a</���~"��Q,�bg/�\C2FJ�l/��I����d��=��ռ���XlxVHYEB     400     160�2�j�1����v��6�ɝ� _����M�T���eK�59��&"�����=�U4vs��ޮ!�y�N��i��Ƽ}�7�!�t� �C8+7IBz9&LhК֤�J��!�j��P�琢5�>�:ik�M�`%D��:�~�e�u�"u��'sˁ���X������g�Di�P�%n�^MZ_/ R�Ȼ�Ŗ�gA�{մ�,wQ[���ԘsN+K�L��P�o������B!>������7.T�F�g.����WQ$5���s2��`��2L)P�VD������������r����cS}(�Ӣ�_q�2�@�n��h��^Â/�)�w�Z!��K�&�=�D�%H�XlxVHYEB     400     140)Mm�kb��������s�0�ndԆr0]��zc�1U�8�)Ӛ3da���џ�$__�bf��C�od�D�� ��A"m�ه���*��`O�Y?��)��:�s�;�t���m]C���H�������'���#�QH�v�l�{�J��CED��.�EQb5���O��S�&aIY�+M�h&j�j��>A�j��{����6�L {'�{���.�����̀B� N�3=���n�JB_�!�0��h��$g,w�ׇ[��B�$y +fk^��ۑ�r� |��7��v��J̤��(R��cjLqJ���)�FrR�\XlxVHYEB     400     170I�d�⼟�-�'_�/vϲЇ5�iD�}1��7?�)�f�{I?�s�6��WD<�I*W�����'�O���Bg����N�P{�>�lk�Xa�Zh�Ap��I���Lnx�j��'�Rx��g��i�2ȶ-�1̎G��, '��Y���V��c������e����h��Jo��aĉPy} g��Eg��O%��7xm��f�2m��mZ�"�N�_w���q�@u�^�2�l�?��}����6N�춖���(Jqm8h�jJ3�T�����W	�ws����/0��kMm����pӬȷ<Ѧ��;��0�⫸�T����i\8��}��L�b�-~��ʨ�6�MBށ��%��Zl�L��XlxVHYEB     400     150ۋ�[]���ۭ\I�����O�7u;�$d�h/�d�o�\kV�\��4��9N}v]՗ˌ�v�zI�K֦�﹜���H��X�:v���Ga�=V�~x#�}E�A
�C�"k�ݓ=�'RE�p2���
i��g�F@O�B
���2E�@�*�2�S&�����Ek$E�ɕ/��o���_�7����s��h��5k*L�b�J��j�À�bd�!�vr ��(�vµ�f�X:�>=kRKR�q
.���sG"�	��_�p�o����a.dED��ƒ�~p*w�;
+����[؂E�_�V�Բg�bt��o����XlxVHYEB     400     190DP�0��^*�3��3���iǙƍq��ݵe��wF_K!̦]ٿ鏍"7s��(AG�bV�s���6G]�i��i|l�;E��T,[,����(���F�yOI�2ْ��O�����p1�}��C,{�	� �TI���C�Pq^�`"D�,a������N\O��J��H� =z�qKܕ����������yс�/�s��]�s�E�s�������9w����h�h�eM�T+ ��I�i���0u� �u�x�*� �8)�O+O�1��R �ᠼ�K���jz�)��~�>��e
�[����ӸUMlt3*���Y
��;�+�6#�@s��;hI�6�ǃ�k�R�?St�蝮a��}�* �1�7U���<#�|���1��"��| �XlxVHYEB     400     150���5:�o:@��ׄTj�
`�n|����Ġ��q��wQ�zjUK��<����E�م(L�o&���2�
o/7�e�,�g���gϛ�#�<+ʲ����r�����/���g���u�T�E�cD�C$�&���1J�p�9f�g����Npݎm=R�x�#/�;L��,Fs��_���C�����w7�Nf�x������Yz��/5 ��l��NI>�=�w���x/b+���t附�8@��e�<fD��4U�2T��*��| P�%�b�l���Cdu��k:\�>+5��K(pn��&22_ �q�������ի6�r+V1�zm���~�"XlxVHYEB     400     100�5����Fu��P�T��ƃC�ȋ{
�=a�	G�僦V^�]�����Ҟ�k��d�<b'U��#%f��b�$�֫k���N���O��Pə�v��嵻���$�7'�5�}��e�T�������Nn�z5/�3���M-_,y�r1Wct-�l.IaZ4������~��S�x}�ޱy��Hd*�)ړ+�]��|��VӋ�f����U�X�G��������1X�_@��W� g~OC���Ae�8��/XlxVHYEB     400     190�U���y}�}�9��͘��c3~׷i�>�^[��/Q\/:UntS����^�Kj��dP�;!�*3�� �jg'�p��\a-$��	�=P6��z�b����yG�Ŏ�rJs����3"� �fW�J��ԗ�@��u���㺹@�!��NI�]m�D�%,&�c��s�� �����U;R��z R��fN�}�&�vX(�RN�������cTqc]��}:U�^��o/��o�f4u�0g{6J����V�=��"�un��,d�H�*d1��g�V�H��䁀D�N;R��	�ĕZ��z����m;	�ß�
{�X�E�b�_f*Y)� �V� +��,# ���xN�Q(�T���CS�S4C�F����Z��W�GF6��>�	֤לM���oJ���[XlxVHYEB     400     140���4�
���U3bQel�i]�|OH�aG�(9G���hC@�b�Z+�#p�V\]�
_�%E�򷇯-�&H���'+�� �pF�����AH�WE� �EA��US~!��2�>:yeH��ϛ�Ԑ����n�2y<��F&N\�Ҽ
FΙ4�Tݤs�٥��'���)8�on%{�� �����˂V6�0��"d{Y�]����˴e@U�.'���@�b�%[33b�W1wV����=<`Ah�Xk Z ;I�����������B¤O��p���ܓ;��}�
M΍"�3<��X�tXjD��7�XlxVHYEB     400     150���
�@Qq����53�?�w6��_6�B4�}^�6-mPS��k��_ <���ԋ"T��%*rV��x��(���E�+����hq�������^v�L�Ju��Χ�&/$�&t:��~їn��<ڏ�:�ۚ�(V�*�9wo�s9��9<'�8_}��(w�;��DJ�(���M���(� ��ֹ�W,_���
X��� d�N���Ml����8s?�rE�k8�c��w^ڭ��d��� ��j�#��a]�m�~�H�4��͈�y;�g�)a!��?���u,tK�9.�x�q�$�a���	������#d�x���y���XlxVHYEB     400     110)�_�zZ�/͑�����1��� �h��4⤊ܻO�ʝ��ק̿��n��[��䈂1Z����m6� ;�#�C ��E�����bs`�r{�U����M��PyRJ[d�ױa��%�jU�������[�:I�S�h�_�&���a8����a� [�5��ޟ�`�LsV����Jqm*Ay�  ���+p��0z��yl֫ �ˣ�m��O��a ��#$�x�88��ZZl��J�IY�X���T4���d8c$�	\d@�{�5*5�� t�Gsmy�XlxVHYEB     400     160�̂߈�bM^��"8��Px�,�U7o�j�6[�eI�.�}�杫�hdy�͎�BT� L��gB��|Ց��M�v挙������v��H����˱��ٶ�2�� �WЏ����?�E���r
�?$Q0���_�2�k��g�7�qbP4�Pۿ��%k^'�D�BT4����gX:��\�;Q���ƣ�>%�p� �d����	h�F���-}L�����fD��-��[<���`{#�p�*)�טoz9v�:�� D�
҃Uzo5EcBV�����I�{����f�͈u���E����l���ֳ����=�#�g�rV����v�C�m&��qaȈ��SBp{`r��,L�XlxVHYEB     400     160��� ;n{"E�|��Tu3��h����Q�'��e颩�=��b3w�Y	"�2�m�%�(k9�9�7�~���~�Q����� �b<)�A2�����~�:��t+�ٌ�Y��8�Ϟ2��ѹ���:.�A7d�rrU6`�G76����u��m�[�OU��E�I֞��)�-@V�@��<��C=5n=��QE�n�'�A����Rq��\��J��~K�o0�95�{���K!�G��惪���=��s#�~�_�7�{�)c��K�Os{F�7v?���G�^�RB�1�{I���ϳ�ݵ ��,���(pf~����H�EQ�Q�l5�Q\)w�6/�f�Fv���<͠��,�G�Q��>͎R-XlxVHYEB     400     150�j2 ':��P�Hx��2�K��A��3��\V���+1�6.:AEN�j���r� ��K�4�p�V�nB� z�^N�f��/�iAi��SΕ.A5��4��q ;ޓ�pH�:�X�$��X�,�A\��x)Y����*`h~0Ƀ5�E4�lHL}�o6�1�O��[7����'�H��M� ��3C�J��z3�\}��M��%8���9x;����C���A���s+�^��6�����a��%�l���n���w���&�#�*�)�[����	�F�M1s;�;I	TH�lj������qZY
8,0���A�h�46�.��,XlxVHYEB     400     150���V�t��j������z8b�p�B�����p�[�żpQ�n���S�%6,�{�WnD�%bYj�/nfC#�u�����V!p1!��7��O]r8��s��Y�<p����4�;q���^=\=I�n�-$����71`�C1祳���J*va�6��L��圐�;l�#0������PB�G��&��c}�J'��/�_�s�P�?����mB�b3�G`��@?��2��B�Uj�h�d�������>���#(
��O�7�S1� �aV���r0H��W��л�w#/��)�5z��+�P��q��:���E"�̩�������2��9 < ��XlxVHYEB     400      d0|�&�]�ÿ����Dp�O��Vf��*@)7�D�	0#U�gy��@c��$��>�t���,Con5J?����$��e2+�\`��c-�_��&�p,��T��/��7�m�>��}F2 u4 1����g17��·e�#����`�G(��,�-�!t�9��1�����0���3��؍�lO�&E�+�wR��,/~���>�`:0XlxVHYEB     400      c0E�4R�@RLxK;4U4�/rm����70-��V���D�9Ƚ֠I�2��Qm��?>G��Xйr~,�"vI�(c���,�t���pҼ����K��)�� ۭ�����<��,��L^� �U�C�z��q)6v��,dK��3S�Xq��D� 6FX��f�����,����{�<9� ,�vxkg6����eEAD'�XlxVHYEB     400      c0K0o�� �@��NP�7g�g��r2�T�V����`"�ēep��Q{ю�D1�f�˞��*���� �4��q�=�a*ۼ����*�\H�5� ��(j���i���f��CC���%��L5�Ϧb�F��+Ŏz��8U�,c���J�߸\��5�L�}��LJ���+�m�������I�N9�7�'B��K\XlxVHYEB     400      c0��Nj�Jb��8L���i}�L�[E5�%��1	��P�/��'��cIGC}o��SE���]��څސ��P�%�/F��L0>
{�s��L����#{��S#>��p@�P$8X����&{��4E�S�8y��*#U�FB]�
�!�������>�0r<�D�뚶�����3��걓eΓ;"ҧ�XlxVHYEB     400     100'��>b�9���HߎԴ-��yW��(y�*b��vQ�T�]Ū�*��/Vw��q���O���Dv�_Im�ꓜ�|�b�D�S*�A�
�?�ϭ��X���/�(\|�8R�C]tr�e-f^��o(l�B�Eï�Z�Y2�&n���4��*�[10a�O�,�F��{Ҥ�c�t��,��s����ѧ^�(lS��[ ���'.��Xa�a�;4*T-?�������O(��H��B�p	��˖0�H��o��C3����$XlxVHYEB     400      f0L���w?�W|��kd�.�V�o �ű�=�b�3[��RT۾��7�A�c��:���������`)�f������48�]��&_����l��}VF������'1��J1ǣprA��YY�R��ڦ��i�N�c��X�X�C\t��e���X�C����LC��
��ū�)���0�i{�8~�R:J+M�m�g%>ķ��]��Z�Ձ`�=�H&MVn+'���ZvnXlxVHYEB     400      f0�da�Z�����bX�5)�;��W,�nk�����j��)Ʊ���~�l�I�\On]��"�ʫ��G��ǾZ�i�+	�6-ǃ������^D���̆�3��ٞc�~���z�uF'��+!'h~�@ ^�<�5�DgX��j���#D0��Ϡ��rU^���YgMY�!+�0R>�L�I�ulv�v��>r�����c����	������V>!޷i�@Q�Pl�1�Y`����景dV�c�þx�}�XlxVHYEB     400      f0R�R���ȹY�#�A�g6t�%��Kē�Ү�>���Q������1�o��fl�o2�_ШG|�t��`1�F�.�M%�����?�{�<d�1�0�H�|x�?�O����N7��M�d�1��jd)�o��&��C�2��m@+Y���� ���]��-�����+��W�
�� �I|�v��!�u� ��+�M}��Ђ�,�(�c�[*�D�5�v�o˫�r9�I����XlxVHYEB     400      f0��|6�2����M���J�O���^G�����[�C#���ݥ Gt݅��x�!����^`#��=NC|0Z�C�u��?�{*��HŞ��'g����Fɦe�T=�O٣�����;�����L뙟�M�%0�!�(�6ͫIyhق:��8�5���F�F����p�	��E=5Ӱ�#T������Ҏ����"X�& �'^�!���+�O�i����y{_S�tsXlxVHYEB     400      f0-���GDx<�mk��j�ZT��o±zb��-�k�Q��Y�'d�9Fŧ���Y�����*��iö��5��5k������� cn�Yl���L�o���ix�a��ݿa�ϝ��Ͼ����@�{�!_���{�%w��'Fl���1G>��H�خ�L�nA����D\av�:��F�N�l����7{rM�՜/9��2O�Ai$�:���뾜i�))��Ӛ���Z�����1,L��C���XlxVHYEB     400      e0LTXf�� i1Е��S��f���1 �X㞪���]M��(�������pޕ�C؂$��'���r�a���"sc���}E
2��<��������忁"[?�6�%H?�~m��,�ci�����"hB��~��ˍ�gU.�>�ie�r��F��nY�)�*t��! ��H�թ�6���8�!3�:S�P�0�d4�����D�䐘I����v:2�(�IT�_�f�XlxVHYEB     400      f0e�g_/(ͥ�� {t�M���X2����0�̗}�I�S�Kp����+F�1���A�C������fM���k@A�:{:u�V|����{�\��-E�P����J��	n玥�v2$�]��.����%R��2k7BjK�I'W8vz} �� �>���ݒi9q�]�v{�a���&G�K�~�UI4�3�1�䫋aG�}l�����gYc�#���c��B���C�.ԭ)�&��sXlxVHYEB     400     150�|���ȉ���eBLT��Zp�+�NŶ�K��0�mA��.Sk�
�R��+X`:E��V�<��ɪn4> #%�k(k��{.V�a[�^�������Tg ��/�w˯R�^f�a��m�� �6�6	Rjd��^o��,2X�w&����2`){�a��ԑ�'��;�GG~߄Q ��7�VL�6z���`!��[B���XY�s��j��A��kH�G��+kG[���f+�('莶���^����y�r�?�E����",s?�I��Sh*f�͠E�f���� ���F�	��x�1g5��);��Z��D��K��}W7XlxVHYEB     400     1a0H��$=6	���kИQ�;�1�Ө�q��C�*t��Ư�\4z'��o"��YI��op*����&�9�S~Q7�^#b�L`VmƓ��@?E���'��6�V�� V�4[�J˓#�d����6g� ]@��j<Z-�`5�Pu���L��t#1M4���V�Z<�Y6��'��_�S'cF2~V���y������]7��;���HԶ2�o;�kA"�\�?_9{k����Fط�������TP�Qס�/"}����d0CRX�31�1� �e@;ϯ�����~2��Ĳ�mN�8)L�'H=gKD�<H��^)�=����b��9-�x���9�� B:!QG�J�����5Tl'u�A�٘���[IZ%U4�6������+�L�9�ٻ���&��̇� O춻��b0R1v}�XlxVHYEB     400     150��pQ���˛0��������9�&_�zH{��}'b�&^�r�^�$s2'>�`��:��9��qΏ��$	�5�B���s�.�.#�m>�mxD]I��4�ȶ�4���̘pG��A	�4�����X[[�[�j<d�r�Zf�N��b5\�y��Z"<��t�op��r|U�-y(��@�Y�+��q�x�ҶƮ�հ������u`�"S�&`$�DD�S]�>�oQ��i0���� ������+V�L�4�Q��-k�꽏ר/�ޒ���r�����l�G0?�ۗ�Bw�S&�� '��Ĉx�qUSh���܏)^ޣ�{�,XlxVHYEB     227      f0���}[�@md����Oq1���~~��K_Wv��`�S�P�2*T��c�.~�&������he���Aq�Z���:N�D�DϕFLg�ԫ��bB�׸ۧQ��q�˽��u)�_��߼���i�\���{��Nه�+O�A`'�x�z��0a��8�r\\��>:�.�3��?�x#1f��Wz���y8+}�6�#/*�;���n�ң��h~,��{��*alMy���>>�