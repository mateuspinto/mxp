��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l�����BO��j���'u��6�NA�%��+�,�
��f��$ё�����|�6��3��0�����!���Ht�����a�A���ϧzdũ�8O��������������Y�8�l{�{�l�Y���U��M�+��-\>����We�� ����_k�h:?��<M��?��Zc4�C�}���3l՚�13TLD�HT.�˨��+��)� �����L�~��� ��[^�3~�4��H��y"K;u��ýN�@w@�[!�q�dD�4DַX��E��ˋ�g_Ot�?2[�4���q`/�n�^���5�%��}�J�Ȍ�\�>,�?m̪�lԱy@�D�@z$�U�9��^/�\��Yj��:�b\h�)hwe�g�����{���{MO�W���݋oUR����sf�����S&��T�W#�gRR���;��/�;�f���@�fg.�O?۳�^#��ڳ;���k2LЕ�����%!�Uf��C�J�ݞC�	�����;M�&���̵��xo�
fq�mQ��x׼oI��G�f"�{1��1�s�����ҡv:kf�"�3`y=t �]��T�n)��S��fE�*�w��v3���O��,����I�o(y� c!��G\���M�c,�i�'��vj��X�X�B>(����g|EdE��j�:�5V=�^O=w�W���+���O%���s�]+���?�}�����4q/Us�]ds��	W�L؊ߋ���*+W���i[¤JתZ��G����a6�c�@�W,�#&V�4�qD�YX�)�l⳺C�/_+Ve5}�p�������K���э6��#�7�M�db� QE����1���e�?���-�����F�D�N�&:��Y_ ��稔XUsצS�;�ř���`>���Pp$PaEe�6��I�.��E�pH`���#�e%����!9Mza�7�8)Cؔ�h�;F�+8û�F�f������8*#7��3Ǽ/��C�NL�g�`G�S��n�Y^wa�i?Tf~���n{q�7���eU���S��7;v��;�>�=�I�Jȯ�!l� �����F`�SL��'sTBm��E#�g/U���XW���f�,{�S����EA��Ym��o��G`�HP������N��;p�R�tTÚ������i�f%c��2���#�.s�H�ڕ�}_����������{�'F��}Y~$(yZ���Sv�q3)X"��	Uʓ2LU!�,��9*�e��R�һۇw���:=���:�sI�����2e�5��JL[��E~%���7�� ��.Aa�AC0\�(nY_����J��=.�k� �E�R�	�q0�}V7ؼ�)l
�K :�rc4c�X�S��Z��5�_�U�_�vHiS��THN4���n����D�E�Y�?Y�r$գ5�;��|(UX�wd��Z!^��_7���M�
�'Zh�?W���
�_e�G���%z�I��v�j���/NJ'ON�����I�n �1t���-1Uj^Q?�(��z̤�7��A�<+���
YϺ�h|��d���%k �f�G�R~��M�n�J3lmh ��X�Y[�r�kA	����S�+�{��\��P����=E>Ћ�9�#b�K��l@.�&C(���kv��� zH�3V��X��^IP�����Lt��YfyZJ堕�q���m�?N4��j�ڔ��|���|%?IЛŰY7X��؀<?ӯ���5��p`�H�8��V����6�PK!�;a�!�ͷ� ���n�j�ۀS��W��Mܡ�������(!��S��_�����mm�f���ce�;W`"&�K/$�Fu��4���A�=��Ν�8t@�����	H-��#�.G#��������h�ְ�k	�+�MD�D����#ʒ�*x&�f��������? ���]6DH�!D��QñҌtiUB��%��a~"�L��� �O	����~)r�Y$zJ�����ߎ���͜���M�C2���rvd��a*�"[��C=�Lݞ�=[�K���O�9H���W(�_�efn b?5s�$yQD�3��z� �7��jWrd^��d�$#��E�R��Mj�%�a��Ͼ��P<|�<�	��y���6E��n��j�L���M,V"[�"�-���Pu��Z欴�S���:6��?��i�2!6�"���ڻg��ZS�D.Q7�X˻���$l���J��]�CdeΘrv4d%�G%]�*W:�������~�Th�� �lklN/�V
�o-���[�;��;����<��S�Q*j����jo܌�%�F�V�W�3�YKn����D��������+S�F��b0�Ν���>Lڢ�;3C�3M�i�?9��E;��⓾(s��J)�`�R�z�!�]��K�N]��ל  �I����ZA�b!e������Fh��R}vVȥ�e�n�b����
N�?�)����B�p�l�dӕ����A��ʺ��܎/�'�������A��,���t�q���>���\c3����lBN��'DS�
���YU���y�cS��ȳ�mCj��3�,�49��5�\J�R���'���FC�����H7m����t$&�D�J�9�Ձ�7T<Gߙ����_��������=���>Ḫ;J>�ufD���$M���V
���wr$��U%G%��8QB֩9�ǿ>I	;"�%t�Q�4�3tLwv"e$��kD�œ]Cq/�_Pq�-Z�;�e��&_�0Gma��25�a��̎%�'�>�Yۖ߷�~�`��ܘ��m0�Q���K�P+MlF����R���
n��L��%]G8�1,��]� 3êO9���w��(x2�Q��nipT���[Ď)0�%ʇ�R0H#ݶD �ce�|��l�j=o�@�{I<�wE�2�@<Fzh�abV��z�t����g����$Ć��H��6,,�ג�L�a�+;���B/<�B���^�s&i��w?H�e�c�b��~7���iEH���>ϩ%�T8#� ᔙ���O�V(K���Ia�o1��̓�x�&�W"1#�7~�����h��c|䯶����.� n�� k�J9�.�lqS�W �&t2��9^[nz�cU�oޣj���8?� n; ��+�כ�o���;ǬV�G�"�Ϸ�K;A6�}Zh��9!z�>��lN�� ��&�_qn+g<o�t�E��8�6�`�v�q�K���M��GFɴ݂]B�o��\�5���F��"�ɐ��묺��rRG��Y_��(/�F�Ƹc��Ƴ$XoͬӒ�-!�8a�{���A�v�Z1/Bk� T�$?/ͤ��Ԋ�q�/��L7��r���lo�I/?�sݐ6�J��eF�,؉�5_�O�	w[�����55�Jh
�N�~�Z)2��=� hw��)[G�El�U��J��X�ʰ���ZBuK���ZǪ�I�`�;*���:o���Ь�B�Ҝ��`4(g�h�2:��Ov�	�����o�Ҥ�{G5e����y�R��}w�l�2Zk�����K�:(xǮ��������9����)���j��.�i�Aݖ�wXb���'Ma�Z����	$F/�Z.�8~��˪��A����t���}������d9����e�\���[��Ѓ,�������G0O���Y��Xt�M�h-`z�f�ni�W:�^�O�?�"'�8��>�dܝpx�8zpw�����\Y�0G����Ɗ߁n��a�	`k��_�**Ef���i��\���?h��R$jl\"W�-qNK�)*B���l�g���<���l(��;�L��(`��J&�yL�{ccCs+8�m�=��1_4
9�����1��(��U��x��/��-
���3�˴Ge�GcM|��d 2&�1�-��	[jeK��9�YW�QƋ�嵤4E�D���?�o
�z���65�,7k�+"��78��g�)��gȘU1�"B7i����z>��|`�����uȑ�����Zb+ޝ���J�1�x�%̗/�܋��d���u����6R�/��� l��l,K�E��;U|�CFP^��cRy�K�5����<@�3��f�LgO�k����Pk�|�����p1oP�Q6�S��jJꑷ�3�W����}=qZy���_���|+�\�GV�bjLU�3ȴ�#%�mV����"�aƾ�p9���@k�:�^1�in�p�,��h}"�~���	�'8�Rz���Ma�gn`�p��z�J�R��>���J�0W<X������k�`�N�eL