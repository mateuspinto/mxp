��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���Z(���H��{�6�b����%{��@@�3����!UPk��r����
M�C�5�(�~�C��*����i6$��fF�e�H�/?F�d�>a��S��n2q�S��A���\8�U{��UOuR#h➣A��\Y<A-L�p�R�d9�xtx�|���oa�r���t�!��S�b�
@����LD�٤���t�M6+H�5�7۷5�X�ͣ�0Q�Q@�J4��Ds�Y$ӽ�$bbY�Nΐ��T�����eM�9ph�4l����%oK�z�۽�Gg���K4�U]���	F?�X��#����`�J}�%Ed3�XR�aQDǮ�<Bt��L{�����~�-���0]�V��p-�����Ly�1�ZR]��؇��fw?�#}7-��[S�H���#�;�|*:����:�ޠ+��"�v�W��5���RH~��)��Ab���:�Q%�����u�hSGI}u�o��/Q�.�ͩHV���d�y'�)-�3xf��h�d�(�k�?���

͞謃bǯ�D�]�l�c�������/�̰�=�cΞB��l��)_9�*T�(��)0�H���! A+[Ť>#@�5��kt~����,��0�h��En7C��㸻�>B�q.�Hjwi)m���/�0�P��Z%��t 7�h�,W��G�|io�q���YU��6ޖz64�M��g��͐/?C�s�ߪ��k(�I��=���IZ>z�����/����z7*�[�ar+rr��|ue��7�)�cT
���3�8��Rfc J�L�za��0_0�墸:[oՀ�Q� rcSG�d?[1��'�%dz�s�j��J��E���?o�{{+��z���a���
N�6*I��E�J�A}�[�����˯!��V$�Dڜ�D#�?�����ɡ��̖�jol�W��!%k�Ux�h+T��G���Mw7���oyl����j����i��4�r5�P~���m�����[�
}�E2	9ܱ��3�g�!�V��M�2��o�A(۫�����y�/�8�(���K;���%���3s�@%NS�s��;�m6
��
:_����Ц�~�PAøE/U*�D;�q���׳��
G�6a[u�����`��wIw�p�!��QE���@m_����k`m��@3���x@�d����E,�@�i�p��~�C�=�����}*����FNLSj�2��h���=Yw˟7��u$���nC)�� �Ff��:�M��ͩt���]�B�gV�NtaP��A�
�ۉ�5�����^�g%K��ǐF5h;c6�f�^�OwK�	g:���J1IHǜ ���4Q�}�/��%$ǒ����,y:G,%9����~eAg~���E Q=���o����MK��B^EjLK���Qr:2U���z�R[s�YS���-6�f��m]�1s�@M�\+Qo��Ccߥ������;������@	U9�>©�Q7kbQ�M͓;Q_^�}���YcX�~چe|R�l�Q���ӠP̩#K��6`cj~��DpP1u����M��
S�Ż"4,�-���@i\(s��g�`���x�e���
:��BG�$~ �ΰ���ƙ�dͨ-u>�C-��ve� ��;~�(�!ɺ�>e�E`�DG|�ozp�I�ԉ����כ� �s��^Ӵ�d�ʜ��x���=���o�)��&��>��g�?����<�'=S^��
�sr#����ۣ+é��?<��a���ѽ�Eڜ#UA:B���J�{��Y�Lɹ����6*� $H�I�&���f���Aw�mʋ�������ō3X���{�ZH����>��Z�=���4���z�Ȃ��� ��Ne��9p%ϒ0����B吙���jZFP�uOSH��HY���0����L��Uu?8H�a_9:�t����3����:�!ց�!A�(��}D�6N��/3U)Phn�BL�c����Ьu�H�t��c��
� �A�������k���]j�S_��r����"�	6L�ʠ�T�?9���ү��U�	��;�D���2/Y#��CX���$���my�o
�B��Iāv��{|���þ�M	��R�s��9�9+2 D+)'=��h���2 �/\�+����2F���E�.�Lj=�&u�C����t�4�򾉁�ex���Z��S5Y���p�U/j��.��������-���~"A��B���j�3 ��b�Rm�9e�����-11���,�av�tC33ة`�Z��{:K7�2 /cVұ(�ՙK3���"��!&l��f��nK�2mDFvR:yCU.T��-���P��ܒwqE��}�\�u^;V��h1�@���s�f�SP/a��#�<�جm26����(��&o,vj�.�k&t}� �ji�tρ�
)T�i!�� ���)����W$�@G�Re�,� �,�k.��8ԃ�*������ٛ>kb�/��ݹ"uF�4\�	�+���
-f+��i�j,�KSdm��+��΅�n���\�ı #�7x|x┾�0�cQ�����@���OX� �͈R�-o���d���`0Lxn��:�T���1��3Z�a������W�D����ta���lt�J�?��KsR����"��snl3M�D�/�þ.�L��8yU7C��
ss��4݃�X���e�p�_f�쒆޻�Q����!Vgu�w���ۄ~��`m��%�{N��s'P�^Z2Y1�^V�Q��Xz�\C��
���ò�w�VsasU���.0(��7j�)Z�gW�.��f�^���
d5FċM��G�;����ƥYf"��eD݋��.X�El�5лEl$�N�O�ɼ������D�P'�����4Ҙy�%�a]�4*�����K��^�guy�R��b�帆�b�<x���*�z� ��h��~��2����[ʵ�v�kZ��m�힧�c�2��#�C��U��DY�G}q\�]F]�T� J2m�q,J$�8�_���j[ou̅m�$?r쉖xΊ%	���<�$C�PW�"L�\��#��V��GV����Ȭ-��Ѣwo:#dH��@�B��8�)��<OE{,7��	���ꮐ���;��"��z����ɰ���t8�CpC1]-4�#�X��}��
���t���4i�v���6='��oA\��*9kL�����NO'����Q�@-�]#OfF0�-ʍ��2�
�ђ7�Ia���1�Ojȶ|N�6!�\CM�p64��;O����~t@ű�=7M������[���rw�������'%�-_B�,�P��8:��M���y�'�s#W�_�8�94��?�k��p���6 ���;U�ZƊ�ŴU����ɶ�.ȫ��W-g�0�s�R l P�1]X|D�I�hQB���78y�%����;$Lǫp۸�8.(�
g�*��N�Y�y�o��G���n--[|����;bh���UWW��������:S�Yqwt��k��Bpa$�Y�&
����g�:֓�3��gļ�r6��U#"�4��8T@��(,��$ E8�x\�G��M�F�5+G����٩�H�R��_>j8DR)����k���=�O���*����b>х��U��y�
�aN��A.��%��خB7ti��z����,�F�
?�6H�/���G�U$�]jKg��D�ݨ��m�#�OD�DǬ"�`Q,^G��=f'������p,��7��~�j��_t-T�aT(@�pF���2����G��܊�<�x1$�vYA�V��C���@�%p5��{��qI����B����q�W�nY�h�:�+>l�r`����i�ۊX�	��D��R��'���@˚'�A-ۄ�5��Dڣe
��@濥(F� ��.�)��S@��F�&�d�yJ�I�G�����*�>6菫a��JA^k����0��������g�`�*#0�U'K̡��Y2}������¨����]� 0��a�m$���r�t��z����&[����V�XF�.���H�I��l�l���;�r�G�������r�Td�L�vn}y8�Σf=�p4e4i�Wwzl��T�*�A�}aٗ Um��^[����qN����U#ŏ�}0�ݥ��qvښ�s=���^˕��?�Ԟpf�4JB�>3>�w��~�Ŕ!E�7\����E�9�k�t �Pxhal>�	x ~�
�zN�ƊJIz)Z˚6�æed��hf  W�j����������3^Z�?����/ny�o��{�
 �1�O�{��U���w7�4�_-�8��}����WSO���"ƥ�GϾ֊xR�� 1vQ2VY��Θ��Iq.�c�R�2Xs�ǮBmSLBR�@?bk?�hf��]�-�f�T�T΁]L�z�§�ٰ~!�y~솮8�c꫈w�'P&�`���na��l�D��ǧ=�I�G�r���?�m[����v��^�����JL�*��Ԥ�[�H���"�[G��Pά�`JM1c@^]��M{`��WYC�����m�K�_��ݟn9��u=��ۼL&�5�!�E�n[�x�RŤ|u�V�!S�~)��%F)6�2�����3�� 	d�&�����n��'f|G;��b�ͮHގ^ܗp��C[}ݠ*�S�VǬt:v�O<��(@-
����mq���&!ٲ�����0'����N�0S]FXVξ.�i�L`�=�I�^�z��8\�
^�����_y(��ޕ�B0���K���A�wD������X@M$������X�h�~�\���P���Eq�4�b��k��2���u��~wط�|9�^Dk�i�m�J��6����̮���t��(��8��0���9����ے�R��7�,��'��)��+����f�_�)[˛Eu�旅o(�@�Ï��J]��rqˇ͠yAd���	Eu@��u���qۣ;�kr�-b	l���-�f?��Oh�;��8j�o>ħf����=c�_|iʏ^�����䥨��!��9%��<�F��2�kI��(��
��z5hf&b���r=+����t�5� è�2<�z��@7��f"$�v2�f*"H>�êw�����x��
�B4�\.�;y��RϪ��q&3�n�|��.�o�3�d��,�oA�3N��%��J�KR���4&j�r�D����~��2�9{�� ,�.BB%�2�dN*G���#��3�������;�Z��ـ����l���L�Z���W� �$ʦ�Kܦ#rƣ]��gM�)�K�w4Z�l�" �y�2��6�,��9��.����0��˘�H��6��V��M��Y9А��;�P=�gf����D4#b̟)R��X� w$�ek죶fLW�#0[#Lt�y8j��r�|�5�e�A��$/��E�u���v�`pRO�aQ3_��h�,qd�kUNYE�2��rЌ�{h�$�4�)M�O�gu��m�IHl�������<��\��������u�K�o��@Y&ГvR �����1U�쿹ALJT�.�H�?���߯C�Vc6n\������:o���]I1.(�_��p������y
�M�9��!y0߽-�� Z͊Օ��e��?� ���PP$ϫ�T�	�~1gg�?R`�#��g��F�X�Ƣ���l�l�c*�'u\�H	��R�{;�y�/��Ki��T�6,�Ld�K�
E_og�jkS짙�cݺ�=�� P������v���$(��2�Z���ZQ�m\b;!8�[5�L������Z�""B/3i:H	{��?���w8��7W�1
vq�7\��F���8:NT�:�R˸�%� �i$ZU��"�3dJM�_dx�Aq�a��^{@|&gY�2�@2b�yҨ��l��|�W�$Xd���x����s,��uq���4G����H:S���&�ʝc�VDT���8'x�^?�Y� fv�#�����>��*D(u�����D�%��?�,?ɶ�%7�J�����`���K�L_���6Uֺ&W��?4^2������x/�$�K�+v@�p��PS��fl��mf��@P�NO}q��U��`4�T~z�����z�Mg)6��(2�����v���HS�+�uO����U_�aI�MCذ�a�E�-tW��<��YΡ��D>�7�f�0	^�AƆϡs`w2x���0s[6GV*�G��Ä�@!k�o�K�G�R���� c�+2�}�k�M}�NX.$��vn��D*)�Hl��d�yK�o"%��ˎ1���P�	a�bRsH��*
�C����7Bg���y}�'V�dG��B��@��OQƟ;?��T��\pT�I�8�D�Qy�[{����u�G�7y�[�>���T╭벼��1��Iݴ��`������g�f��L��_S
��o��c�2A*�����:��]��%�F�7`V�PӤS�t���%�9�7�h�\��t8�H��x����Y���)lQ>�j�]� �Դ	��2���Џ�D#���Sl.����SFْ��}�&��ܵ�H���7o+	�3f-�S�2!�YA���N7zZ�y@�Z�V���������Ӕt�)��5ͥ�캖WԤ���P��i�r�A�Mr*;n��Ԋs�WF��W/�N���~�H�0�������]�|�bzpIi����@�Q��DaNA\�kP{��A9˵H�=�Q�[�CA�a=�o������E�O�,9/�Gv�ԑ �РQ��؋~���ikU��1`���]�ۛ�g#r��̕�7ƛ'I����r%Cf]d�|,�G	��*U2��8=��%�
�I�
�#�Iem�jG,wF�(�V&}42��x�(3Mud�����9�H�{�����A�-}"��o���E�������ڏ-�����A�۩$��#Z.HW�3�"�4�H�5yn�ee�<�H�6�h�/��I.�m� u1`��V��U�5'�o����@�*�~o+1����&���5V�j�䢺�ʃ������)� \�Q�_7a�&�u5�UL/I�@:�d�9ׄ��-��2��8u7�c!L��$�}&����bU`@?#��`�F=�5�k�k9+���X�A..��F��<[�N;HN$61�3N"E�e�Z�����i���y۱�w�ީ��IܭQfO�(5�n�or1�����>�P�QBV�sߓ����A���1NY����#�;z3��h<���|�(��7�:'ՋNi�9H�O1Az�䤏��tDC"���FҢ�#�k�E����%�m4o><%t��2�>l�J�=�;U��<%�ï� �~$w˽3��06,U��!}��'E�x)�ln����k��
����s�N��m�'*e!�5�pW�ۢ�yhZ�ۘ.���S)Ӗ�%Y�2���������"��I)�ӣ�c��pBI��Q�cΉ��S֝��b��&j�:�>�t(5�����H�B�R�Rz�1���'G�5�n?�V�]��!ʖ��p���z�C���&�MM�>%�>�K,m�aqO=�s�nw�k��4S�s֐a�u�7��1g����M���W�7G��ȩvN��6w�5�ʓ����F�k���l-5R�鲅 4?�K�D��_Mp�آ���3[I�2Y�w��ཱུ��F�Ԣ����WHwS��sY"�8��4�Hɲ�a�[J)aUq���Ky��HW�����y���f�\3��@����L��0���ݾ>�e�9u�e<�D~����(+�Sbv�N����7�6�N&aƀ9e��;|6tg9i?,�:iH��q,�Y\�)�5�'ߡ����L!/E�"7q�鑁�}cN�~ol���r��h�)f�9�N�G��qx��I���	΁�S��B�,
>��؀���hy7�*�D�_��K9�-���I@B�׀X���Ex�kfK�sTƒ9��Ȥ}������b1,K]f�͛����`2����
��Q�o��bH~y�/��/���x V2s�+0  �n��]2�4�P��7�k�g�y_F��O�&A.�27~��˺����:��}Qn�Ȁn�s
h��7w	���㦴�b[��vd�*�� �
[�3�māa�AB�WmU����?n����T�ю�~����+��j�]i�U6��w���R����}(���qsf�D��L�hM�^��9{)8Ia�"����A�m���SU�\�F�;�w8Ӻ��Z*J{փ�191��D,� ƌ�-C$�xE\��qr�[�)]bӥzD�w�l��Nf����=<ٱ �ei�F,���qg=��&m�G�GXl�T�H�<���)�Z\�&W�����,@VXkt��[�^�Q��XIezm�w=�*�]aN��S�ȄM��e�����;�?�	���;�kZA�)ߑ��gxZv�|�j��5DA�/!��́;����g�g;B6�u�7-��H��c�o���e�Ȝ��f��p�"ȧ���d�2"��YcR����
�x^dV6t��,U���o��13��X�}���ij��:�s[�mX��|�1$���H�<`65Í�B�8ae}����7��X#jQ��PTC��Ӟ/ .`a{�c�3�Z���p��-�oL�Zkk�E��i���!�ɂg}���a���tޗC�,��J�L�t��0_�j��:�s�Hl�M<	4=�=�Dh�!�s-A���c�9���� j�<Wr^q�7�6w����JPNO�(Bk�|g�/���ל��z�td�A�O��n�f���~�a���Z�EdQ������%ik��ڜo2`m��@
��z���|0��"�6�Qy�TQ�7�{0�)�R�WY��K���H9$Y��E���-�L�w/lg%�r�pZhd���&��j�m��.b��+�o���[�ca�ҍ�ߙ/���i�y���:Q��X�ң�����[�*�4T֤*$�|��'��v���?�B7���_�WW&g���^ �5��*��P�5ܐܽ�fl�cL�]�j����w�T1[�͛���S�;�0?'��i���u�[���|�������F/X��N��9�� ��_�Ч�5�YE�
e�jn�Եr�;���2Ƈ�k�%�53�-9'`�  ym�&�_>�����BiǺ�(������<P������D�:p�S�<E�yۺ�E�
t�� ��}�� V�k��&���:+������M�lQ��˵������{��������:��1�]ݜJA^����̱?�Ztϰ��>�|;0���\u�p�_�-h}2�OGF�S[�M; �O>g
��攢���@�����`�֋��٫��(E�#������G�-�82��R���	Mhd��#k��3.�Ρ������n���?#q��"ޛ�쟑�����Tj�h
^Z��+^��*���-B.�[����v��T��	�_g�KC�C8���3^
�{�����lQA���A�e��@5_�������+7$�b���%�S����~K����z�� ך�z��?�e���Z~��Ut
W�N�}�7P�8k��DK+y�Y� �[bUN�ΡW.�uOS��}^���o΅lh9�Z���X��*^^>2�<�>}s�)=�@ +��T~��Q����$J�AW�b��n���mIE_�o�󲙬��UV�G?T(�#OV��[
«�j������dA5��S?]ޟC����j߽�I�W��Z&�!WKĪ��ݎ���?=)�kz�O�֩��}o��w�mbb����\�t�6#�ѫ��,g��W�9����Y��[k���AC���#������SR��{���+}��C�p��6H�E 	�)3I�¯Xw��[P�u���O�z��A�*�c� +�F�61G����X`^�	��eː���԰�e!_��G��&�qmf\��� ���>��2��*&5���������R���(�x�_0�e�1���N��˽����j���0ҿB#�,�]�F�E�����e�v�T�����s΀���3����-׽��l�5o� ��PT�-|���R''9������/�	�cI-LoT�vKX�����v��!�]0&�F7���x�´�C������J�D�u3?������[�Ս͒l�Z۶�� M[�y�7N���;�ON.O����꬜J�`��^��hV��Ǧ�E[�ڿ�^Keo^�O�k��V��2<<��Z����.�\�/魂�G��b!��:��AR�-e�_ޤ��ۈY��y{�8�"�ܷ���8f~�L�Q@Wꔂ����T�r�wa��%�[������T�����\�|�Z�tѮ-� �.�0a����P���|i��gvei;��≧�V���==���"!Q� .��΀��C��/��߳ӊK��4�qض�}k�R�{7X�1�ƍc�Ը��_^����2M��W�]�˚ �I5w���C~�oC4���+0��aJℾ� %l��D@m�/�O���+2#O�POU���E<HUt%��!*E�O�[UI\ѫL ehU�7�M^��T���N��\kjW��T<ؕ,|Xz�9G�������_�k!E
��X��x@L.q�|뼿�0W�/����fbl8�0I����TiL�}ݷ�`�L��4�4��n;wڝ��4�#��pYn2*bFE8�-���*��6?���ߍOW�X0C������SF�#�7%Ϋ?=nډ��u�f� J��5-.�]e��QJ��4RgNH���Ƈz_���u��)�����<N��@4?~��Ă2TUZ��Y�����o�Y�w����絁�&�w1���| ���NJ�`�Ɋ 	����,[�+�w\�}1=x�k&F��2�\A;C�C�� N�9/��$�z��x��4�4�{ǝ��Ze�m����AȑH��9�$�"��U�H�[�B����H����eנWi�H��e�� �*�.�z���L�_��ռ�j�� ��IK�vq�'�u�eQO�S��1�X>pB^�3����0�1�����������$�j����Q��$#޾p�2�k�?]���@��
�TYbj�_�	u��-ܯ��B��D�`�^႖bt4��똺@qA蓧��{��h	�ڣ$ް�M����/��^����� ��dKj�cc<ع e�0)��[s;�X�Yb�����/:'6�k���AF��,m7�Yy���'�H��7����Y��u�
Vh�Y{/���{Ղ�v`'D�t�s.��v\��i��'\��0<?I+���s�����<������I�3��xF=������Ղ.�bJc�犙w��G2fAu5�pl񱛲�,��-� ���iA�|5D.�#�D[g:�|��3���4eS/L�K��R��Ĕ�����L҂▣!�_(ĩK+Tx-���֨��}	���CL��a�
�Bu���!�vɭ�}d����M�[���Ľ1⣷��'��R��-� ��N�[`���/Z2S��_l9�\�^zd��P�}ڊN�s�ˇ�<�][	I�PțՉL��)F�֖U�+0�9��&pL.p�ɜ�7?�1so,�l!�XxN&b&[�CA��ؗ�Tg>��W��f�>0Jܔ�b7�VIL6Ӫ3Fp9�h��e�ދj@��4QO�@��k�B����*�9�H9;�ف�b��OH�k���I�p����Y�u��``���m,,�K:���K��p�"P���Y�K��<����z�,Ku9X}Z����O��6&p� / ]����ׇ��T7U�C�GKO%r�Z.z^��K�v�U7�Q��7�>�!�3j�QG������'da��d1�B�D6��k���á���bl�NInV����L�,�1�o�����Z	���7�.�9X1��S'&���h�)Y���G@^/���6��~^Q����T�ǜ΀[��|��d5R�b�����P)��  ��X#���+�@��� �w������}Mb�/R�AK�-gaim�*��jF׼�d�ɾ%��+�h�s=@�r���:>���p{�/�W��u��2c-&h�������;:6����qm��[��ܴ,�����:�u�ΐ�-%)OA�#��m�W�F����ʙ�L �y�������u,i"\U�C`��/�����o��b��c���i����Z�vNo����c|�~jokb�Y��[)�� (��e�+�����E��*)ASQ#-`��+#�V8.��B~q���"���NܻD�+�Jֹ|�6�1JQ
�/�e)Ub�Y�U��F:ZUX5���u��?�T9<������HދT8�>|^<S��]y�u���[��|o��p��b�y1�o���»	�����ygdˠGཉ�;�Z�<���a�RF����@`ϽL>�gj�,f����fɄ5g^B�ׄ��;���^�Q��o��WM���
������Ԉ�U|&bN� ���æ���x��e�@�%љ3��/�tE��xN��?����Xb,@���}�hZ���7����@:�	$Kٰ�	��t����R)�c�4��3ke��#M�A���12eg�E��:W�@��x�bn�V�z�����Vިio��%L��3	fV�\�C��F��T���W��Ê��lȴ&�	&c���0U@�B�0,�h��hn��c����%��Y0�v[�R�Zs�����Q�)��.�T�l�3�=�!xA�n%A���E��!�_�J���W�-z��MȦ䦧���J��5"U���T��睛��©}��+�0-n�X&_X�sؽ��]O�ig�^ui�G������I��[b�� .QG	�`�d!�p��h+xg�.�Q��t�Tg���3�+s_�����`E��r�����̕��m�#`Ϋvb2�R�MȻ�*}b�y���"���q��^e�����C��O6��n��lL�yȨs���x��$OfП�����$9���Լ2<���7�xIm4��;X�ZQ(�IP�T��ݬ?=��p0�`��P�I�U��]�X�x ����/=�-��E�\�I�w����nZ�R�w��	6#>�e��=2���Zϒ8�/c��8u���s��p�g)U���߆`��˽�j�H���BC�����՗�~��,�ԫ?l��a0�'G%7;��b1����[f�mwSZ,�48V~	C��u�@B�l���N"���P򟌙N���{͈yw3;�zn�~;��}N����'M�֟��/�G6=\�A��x�������f�{�#���)_�b��L���C#���{�r�h�k���4�wuFp2�(��-{_^�H�44h��r���4��^��YQ�x�a�Z@�K&_�H�Ԃ��2}�GT@���WaXMhh����/B��gli�D5u[�.˷�ʌ�v�Gq�LL�%�-��SwTpe���d��e�s�d�&�P�����ϐMW���+�N�9p~���:@���TU�	ڕռ:��8�^J��2��`��R���_�e�ؘt�e~_����!h����i(�,�����K)6�p�@&6�x�l�t�"�:�a�]�p(%������o������5>�uy4���D~f�TuL}��lP1��Pb��� =�L���4۴.|�����ѦM5���Ī��Ra���,@��D7�ef{����)��1kW�^�ۭK`��8.�[�=��~]}���?�=�̮6FD���	�ǆY!�0�BK�J.�*�k|��0�����gY�me�W�˹<����8{U���
�	o����"Ej�#U�X�ti������'f�ʯko�[F|�;�Q����N��k��'G�����P~IP\ �O�γD��[d�$Ⱦݨ��R{�m&�� �$G��������=}��TM6�1S3����Sf3]#���%������J︮Y��0T"��� ��e�7��m;!@�6 ֏B�W(�l|j��$�T��j���=´ܾa}�E�p�a�4Ba��:��"�l1���m+<�r5�U��P'!po�(�ٜv�$�42~����[Y�7���4��ڞ���0]���@����W#�=��.��g�5��x3�����o��܏�z%~/����
� ��xlϒ<���R5�KE:P�T|�6v��@+]A+��L�4Kt����l�'@75(p�z%Ž�r0ba8n)����z�aF1�k ��ռ����3��h��A�<�`��3�EM��AM�ҕ2�Y8!j��B�.��k��d�Bq�j`Z~�|} 4�1�m��#e(7瓠͵|�!e<���d�v;�������=�G{~��,��˦D���H��-9]2M��"'��9�s�W4ʍp{���>v図
P��A�a����^FIг�+�k���GQ��K�>�_31�)�6�q$=�`����O�O4E^���3�O�(�:un��pg�l$:#p��(��\v�@����y�/��:�R��w�g���D�ρ\k��|Nw�O՚�1�>ǝ�Azq�E���׍cO�H�)�g��~L�������!A��ۦ�Ěڶ��g�.���	tl|*f,,\.��%]!�Z &�_Ɇ��գ3�l���<O��,�������cؖ&TuH%?����j�b����i�L&�)kn������M��O��,����Pp�'��6V/-G[�ɝ`*\[�ң��}���,���[���^���$Q�ۆʧ����m�m�zo�ng���}cp�@B�gsc��V/��ͥF����t��~��+ɔt����G;�ѧ��g"�b���t��zˢ�b�p��g[j�.��KJ�ǥ������⥈�l	��C�8���A�3��Z^tp�r�إ!ح����e�K��#��x-�jN"�.��.M�de�.g �����.)�y|b?@p"�r�d���Ծ����3��ckP��bM�(��-��9EJfI/�7X<$L��w=/��B�C�`ķ�,��T�c��G�(���|Jb�Co�+�M��3�U����x?k���Z	>z"'>pS% �4߹@�� f<?R"�[l�ٳ�5om ��i��ޛ�Qԡ=��!P������]R@C�zkA�Ƽ��a��V�S��e�@!�5��KA�X\h`[q	�K��s�*e�oE΋��]�%��|m�1��|�6�"3TA�u�{�1�	3�3F���>��pJ������u��F5'Q�����Bg_����y\(����Qd�2:���I�U^�����J̆b�����[M��`�P9���#�Gڙ;��(D�exi7��@e�Ȟ26͂<Xf"�[��m�-:��%HE�E�1��=�����I���AK��W�лR��R�$3�+���{xv���*u��|vtޜz<}Mޅ�����pg�x�fǿ_>Jt�����M7��[�s �+�F�韔�Y��t[N�X0n�qA�8��@����7*���Mc�(��?W����E�ü���v���$e9sl:.�_�6
ih�r�!Ue�kFK�i ��$+EH5-��w7I���i��.�9�'4���iUd�+�^��y���%��H*��\r�v� ˓���Jg��Ŧ����6�B�a�xM�f�x�m��~s̬	�1es��=�3G!2`sw���o,�>��c3�.�F����Ne�Ww����e��\�M�a�<���-��)��+��=ͥ"�iQL?�L%��(@�4i�B;I�G6��Ŵ��S[zx$��I]���n:8��޲�A��L�a�I�]��	��׎v%�`&y�g6h�Z�C
�f���J�g�:��_{L�<���ǵ�6M��~�qq�
���h����䂷B��;���U��|��5{�s��4���o�$�i��+݄x&����wٲ�2������T��Ȏn�ӱsS-�My�xՓǘ�Y(�5hro�ɠ���g�K��{�z�!̗x���u9�� ���l�����{�L�Y���	�͏��#�e�~�_H*�Y�,�R�g	���9��t��RЌ�`ǣ�������+�����������$p$����q�)J���?�a_�)y՟(��3�	�~��n�HM�{�(<�h.'��T�I�6;hs/�YE�#J�}. hj3-��0=;~"*��*���:j�:?T(X5�h\��x�F�i�@m��6_��[@u�U���P���P�'�U}=�'��|]�(_��4��� N����wd�{��M!��j{ C�a��}�6��S,ud�
��D������<���ȑ0�B�l#���#�@Xvǟ��
ٖI���)�e����!
>��4`a�����&���T�yD��W<'��Nc\��z���4����5$-X���wxdT)�5���k�b�� �n�_�����s��^ߘ��A���w�v��6���gPu��w6�h)��E�w��J�z+�?w.3e�?fPL7�ơ�~����߆�ɯ��E� �%E�Ə]�oT�A��Gs�-9��n���m�v�����6P��v�6���9�7y,�w�����"-�YZ(ϪBg�yċ��4A�!u��ڸ0TF6�K���]���{� �W�e��ӊ��Ň�W`���~Ha,���m��� W��z˶mS_;��Q�N� A�_��_���|�u�xp��P�SBCP�#%�!x�4ж�5���*;�T~����D`e��+�*��t
��$)�MH��T�`�<1 1�«H��NġP�����L��ۻ�'O�ȓ z�NW��z������ȇ8�@��n�7�1Ș �!-R�$Z�}!u2Mŷ"Ļ�;�+Qñ�&m��{�fj(�g�uۦ޳�'�
=B�R�h_Y�:*��8���1�>�$��/F$e8�G�F�z�N?L:6�,�[z����ʘ44���O�Ԓ����Q������*'2ob3�]_��O�re X�΅�-Ў�O��	��$�\S�Sژ�c����AM	H�M���)�΀QC�f��G���J�l���$�^�EY�}Bx~o,�vF��g�����LxVI{v���̦�2{t����~�@�v�\�kr�S-:���E��Y����=�\�L�VeK���S�k�43:��M�p�t����i�%G��G��b;��.�7HO�a|MiL2��G="��B;���˯�����/��{����YG�������_���|�$�1����g�eZha'��I{%mX��c��\4AsTε:k�+�zn�w:�8w;�ּZ�!E�-U<�0���rҮ�}��]�:oe���<�<sh����,�#ɚvG�m		�����Ts��`iE߂;������k���mL^QBrB����qK
�[��U��HRa�R����Jcq��F߱e\����� �JԲp���Q3����XK&�3#��(���U��M��#���BV��ޤi�g�i;�b�	>�9yj;�:|3hA������_+E�Y+1��X�IkF8wJ*�m�]�Qf�]�`sɄ�$U��u�01V���y���]w签��EO��d��Hch�5�56
����mo���o�z\����\��m�%�I�)մe�J�x�Z �<>]I����igC��w�X4)�ыT_1^�UJ4��?�v�եW�������q��0WUI�T)ZA�'m����$����l"�/l�.!� 
e�P�fͰP�|����i�]�Z�K���O�4�W\��(��¢���'{���,,��D���Ҏ����M)�z���:���Z55?Ț��O_�GMG5�y�j2dO%��j����Wa��\�Ӟ��*#:�H���1O�3�������Hr^ċ2��'��;���<�5���߬�m�D�/��_c��g��?����'���gt�ɢ��Kb�+�h;Ԩ��!�]�D�ǪJ�
���(.]�[�;!z��j%W��IH���?���O�	i��o��*���$:l�[�'����ώ�T����׾�IN�9�tB����tv�^��(d�ĵ�j�m�\�z���[��X�m� D1Z譭���~�"���gǹ^_)Pdkx G1�E��֎e���J{7�AI����v�U6㷘%q����	�m�X�2����Ϙ�&�W �6��'�^�&�ϫ��L�P�Ч'Y�� ������\��5�*>�ց��
��k�-P��,������?��h�5����"�?�G��P��0H5���z�NL�iy՗�\Z/�����4�v��Sx核F�#6��j��������mp�KMԤV�/�^�r�%�~}?F��v~` n���#��Y`{�G�������W0=*���:���l�F$	%����i
BRQP�|��z���n�/���G��ơv����BsݪzI�
��֦�]x�'��U�#B�I�z�4$�O��9��-����#lb.%����X�y��t!'�n鋽�"$��>#*��ڹ�D�Bh��E=t�*�ȹ�2^f��:�ݽ�٩1�U	��U�Z:D+��$7d�峋U��v���!��"�j 9)[��?	]&Jcqe�m�+�V��?�&T�	�N����ݸ�?od<��d�z:���n�k�˚P%_�W���o�f��b�ɕY�J��]���KT{G:�E�U(̾"E���I�ֳ��C�^���?��ک	0VFGX��C��P�qX(�-{s4�f��[�C^�䲅![��ዃv�ʡ�:���=8��\��B��
��T���I�w��9>���#7}A��\�mobY`�Α9��cn��
͜�[��fC]V	ҡ�O!�׻Ŋ�즡���F��3F"'�ǿf.�Н��A� �����]]�GO_��M��n�,�~�{��ⳁ�{f�;�d'��-'f3��>,3�HUOD8V���;J�����xZjN��p�G1{x}%�?h��,aVf �ej己�'�Q+��Ox�c�Xn���q��^�o���	���xۋ~D�;
�7b��B�Q3�L�V4�2�:nj�7e��1�@�����9�zK�3ôd��*c����hh|�dD�s���=�@�ˤ�@O\�"�ߨ�C���3�[@uG�DT{6K\�����s�c�XY�+|	���В8��Uǹo�~o�E����6�Q�
�+��Ɇ�	[��7a��m���4E�V��8�m1�VX&���	�(���[�A�-�O�gjp��},��Lo��#��v��'��=�Q�I�����hHءff,��6���.cHo��졥�1}<�ܽ�
��ƹ�����S!B3#d�[qYd��̬1%�˻\���	O�����{= �Oz��?�9�K�̹���ߊh���������^� ��*Mm�Nި;�aw�Ζ��×��}����خ�.*)S5p<����[O[����|��j}%>�Z�*,Iz^���aJeޫ�W��v����M���1R�2�'�N��R�(���M_yǨ�P.U�7�a�V6a �k�R��̤A]�@+��Ո��Z)��}{[��I�P� |�"�Τ��]���2�I��mA)���buʂ�*b����9;�������;P�)Y��~�1���w���)�����O|��`iȆ��I��2*��R�\��KEc�.p���N�Ȳ[>\%&a�~���dM�����Y���]��FPi�!.F�B��r
�l�]���CP�A���*b2)�����w-�,?����9\CX�u�m�W3@����[���� *�<x���d���3e
��~�7��j�U����S��ޑ4z�+
�T��SH���4�t2d�:y܋�~�_y�)���G�KG�_�qo��y7OYg�A�f}/���<4M�pfa03e���KuU���gjD�����s��k%�#.��˶�5e\����n���(�G����%�6%�q�����ucrEX���f� d3���C�&4� ژs���@��GP���G��$�HlL;�k9[��oe�������胐?ÄS���K·�1<�Ύ��� �卓��dI�@>����,?8��40�������"4U�b�Ţ��K8ªJ]{C�Ը�O�fA���A�pN�w�w���ԋ��!�*λG&�]e�.�^}[�\��5I�.�HHa���X�B��tnM�]�aŪd��M��|�3&�C�@��#�Na��%������7�0q�v;����K؞ȃHN�7IL�Q=C���<�!�nnX��Kh�+Օ������m֎��4u�����Ɏ��xte�$Ql<�(�����~&��32�� Tt^Ѧi#�.C�t�|��y���A�����Z�Ě������g�|x��)ʫ�l��mMQx�ki��ٟ-"�����CR�^R��\�J�
Zg�ǎ/[��bNXJ��w e]�1���Uf3��y���X醺)��]�WUE�J�}��T�CN�Tcq�@��Vh�%�JZ�'�$O���nc�C�:J��VZ��Ո���J,�M�~v����sA2��"4��6Gn�@�?7���C<J}Q|����Lo"���S$uY�ed��h�YF�T�n��ĸ��:��J�e7K���ƨl�����"E�G-�Uc��
�WW_�q�$�OT��(�S�7W�`��:�A��?�;�c��˽�U�������SǺ��/m���ތ�����gQ�T�f������U#��w&Sj�r"�:W�%���}qd���b����S0V�����t����9�y����03�Jt�O���~f"��0�$ O=�1���%|q�� ƨI`����ԩ���C����V���GI]���غP��. W<�}o�-�����h�
�X�fem0?{d``~��c�\��\�A����˥��9L��	xg���YX����d�M�� |_ȷzw���%-�wH�_�xN�O����Mb�d�d�xw3P��,$�4�._pq�GW��I��2�i���%s-��je���F:��Jk!��-?�z��Œ:WU�܌�ƈ	�*��OF�L�M��f�혚���ή���x�=����S+
З�F��d$d�+��|�h�FK2���� �5f\�#�-F��IE?��+�\�W��k{:����ˊ��z��Ѿ�4�˝��x]�A�T2��͕܀{e��w�H��P[pU�P�Vl��s�s��a�'�r�,:}��"q�v-;�U:�[�l<�"x�_W���!IaP�z%��:�V�[#����r$X|��.V����*�_�i�MY���be�1QoeR.�Շ�rp$(/�����#E�C):�������(�s�*$Zfӿ3 �j�R�"_(�I�Jn	��5�yټ�>���-^q�"d���z�tpw4��
���O�Ż|)�g$��0.�!1��ڈ�K��~.���7��w�/=�V�Tl����FO��|E^�X��D�~�}?�"1|��m��?)��?D�E�e���X�:�5��t����ibkg8�����5*V��I`nu���/Z�8�%;�a݃0��w�hY��|�{��-+C��Q㹴"Qz�q��7+r�D� �`���y;�r ��IWy@�rE��%��(�hA��9d'g�Kl#�$��D|��Px��9�b�	�+@Az��C��N�xB��ulL|���l%���_K�N��hQx4�4�3�Έ�jBM�����Aw���)۲�)���:���&�֮v�i�����ƕ6eTB�ݽ�o���4>���ub�<�:l�3ߨ�3{�۠1s�0��q ��B�S˳�܆܏��`U@�2�� �(K[��ϣ��T�2�������Q/讴�zל�E�U�޳W]Ӳ_4�],���⡅6Q�2V���B^y&t�Є�s��;W8��=ZW
�ͤ?ɕ���\Oc�Կ��3$��4��u��OUh�^ޛ���s��:��|�a���g�^��π��s����/P[�����T�:!0����EQ�ږ���̓xz��`q�`��ϋv.ovҐb8�n,�=���CS���uָ��������M��oq�z�7�#�䞐ܘ6r��N!,�=��d"�D�xS"�O1"��ϩu����V�qP���7��2�1�� u�FZ�0�FF�b=�pz� ���E�d9��j�B��2�Xe���� �6-\�k�Y  ��u|�J!���Fy��[��^ �Q�@���'�Wj��y�@T*[�[9�&C��l=�a1/����q!ˀ�g��7aчyɈo�>�˒�� �D���|!����oK%��K�KљROc`U�1��X��BV�v�m
/S飈�Mk�z��VT��i��t{��{5G�o��a�
��ܳu`�p��鍗\�fÒ�q�/0J�+����GGT��^_J���S��onQ��1o��Y=��v�g�B�j�;�d��9F��[r�!*�E�t�d�}o�n=�������X�uΔU�.c�
]KĖ7W��ӷ�����%C���&ӠJ)�%����{~*L
g��-F���J�����w� ���.^K�)~r�ĩ��"��t�=���^�;��*y���!�8[�O�#"e������6*d�z��?ړ���EoZn���k�����-��[n�d3��h%��:�5�T>�+`��<7�+�^f2�2��m'%�B���ڎX�S�/�Y�A?Z�ﱮF�3�:̽B��#hS��]��5#�X�B�p0��v�%X�c���BD����!���.�����`��5ښf���h�U����&��`t%����~wy���:�9��5����Ϩ��ߌ�>�4�~�z2cA��O� 1,��*Rr��ͺ%j�׌̲������Mr�phbX�s�ܦ_����r�o:�+e�ף-`k���R�pׅۤ�VP�j�C9sW�PR���~� {C��pK�P�9������:`C/���Lp>����tM��Aa@`��b��V	P���-x2r�d���}�ߛ����#���o�ԓV�禈�T�ށ� �8qR4\�g�"KKmR��S��Ϝ�L��*Y����C�#=ꀫTiV^��L����um�+M�g}��5�b�84�(#*&w���cz'�����Bk��H1�X��R��s�F��h��a�~��n[{�P���VM�#e[���b�|�em(���-B5QW�L��}]�Y����δ���
|�� ��2>:�˝��N��@�$
����چ��Dᓒ:�%��6qTn)���3�i�;|U�΂>C���^�fWY7�� ��Yp%���xP?����u'(I����@G����r�iy��E|#t�D�0V��}�Z�`#�P1�"���������<�����T�<��R�v��qh$����lm������5ɧ�VR소��J@�ɝJ���F��tv�n�P�K�uSαS�O��f0�db��Jj����?/Mq�H�1����`Ø�~�M���Z� q�L�`Z���1�k����J8*�&��5J������Q��]H#�Ś�w�yFOn�W�L㣏5Ao}h�Z�苗�:�E��Z0�<g?c�X���"�� 	��KEL@��C��^�X��q���P*��B/��r��N��f���O�@��pH ��E5�Rxv�.��Ĥ�@^�c!}�\�7&h��w}G !�=��)���ccRfL<;G��tDA2>#�%W�{��ru�DBz�1�=�.���\_m,ū9i/3�'Է�:�>��/���� ��E���߬����~B.7/�B��˚�q$P��s����vQ��T7fZ�?�׸�M" ��1�f���mt�D�Q�qx7������N:1�tؠ�y�f%~����BP�� �����}����%�x��X��T&Zhٴ��ڊh+F �+r֐�{6�kV��ݜ��O%k���ܚ�tVVYX�����/��W�Ұ�YNK�Q�X�d?�a�'�l�}�\j��`�B%=��)�M4���v7��XWC�I�tW}7Z�M��8
��� ôH�ѸL�N{���"+j�]�;��(�tY�t�E^�_��4:����<�������i/xq6�w�C�k�|bb!���^�'����+z�/�L�k!�p�>9I�[t[i����i����m�!�wl�-y�*}�la9�O����o�}s����%O"6iB/k� "�"��m[ҽX=u;� ��9��5n���``�!L���$ �/���#��jI�^,�_8G�#3��_ϝ�h�Ukؠ�>/V� W:[P��x�;8�)�Pܯ+�@c��C�{,8 ��j>6�lx�e�BD8�㞚�my�@7��Bo�lNB�c̈́y����ˈ$�s*N:��qņ�Xk������B�x\�e���N���( �}������	}_?6n?�E�!���6��$ތ$�R#�H.��qd��58V����n�|>b^����0���b�/f����t��}��3�$�#̭��9t��Rh~E�y#D�K?���c��
��3�P� A���/���-D��^��=DO���3ӌS�0��	�q<�M��[0�.s>�ڥU��d�)F�Q��8�Ee�0��|%�9c4m��j�"�����{\!���JN�38"ڍ�^"���h\�u�?��B���+��`cL�d%����W�+������Q��Vܻ
�#n����d�Ly�h��(v�Wi��� ��?r&��b������!�(��.���We�+ݚr�����~�m_(^:��-�z���B[����YS{&�-�������Ր�y��E���:�֜�_��	O7���*IcP���\zRr����j��,������tfr�$�so8Q�l4�\k�┞¶Y$�ϵ:?��m� �,�%�f�O��Hu�F��쒪���awj��`�C.�m��Q�&@� ���	�X6
�&��>Gl����ר�h�TR��Hf�aC����:D`h��Q�zPr�n�z�Թ�0A\ݸ���kx��P�Ԋ+�N�s�GC�WʏV&w)&\��G[�FF1ݦyÙf���������,�mZ��!�eLH��([#5�_��B9f�&-!�W1��o�:"hn_�o�2ޖ%:��!}iyc�:E;_�t��$���ZU�V���!������x:��!x����f�܃��~��h�u�{�t�O��8,����7��4�j �ҩ0�8?��	X��=���Ui@�'��pasM������"�����N >3�$i�[��{�ndf�]�1�l�(,��EF+®� �m!.|8�A��~0E�����nPzњ*^�J-GD�x���hA�X�X_�""�P�,�$LC<
���j�7V����I��&���W`�[�#����c���W���@#L� U�}Ұ.F9?1�&�ѳѝ(���)�u��hW�`�@�T@6'�L�q�y_lt#��{/�Y���u�����ϐD`q�Ϫ�ᷨ>��l/6���@~�#n��5/j���������&JȀ�*��f�]��_��<DL�I!�R@MJ���Me�/9���Њx��k3!��qǻ��8��,���]���J�{����������9��#H��?{�\�r�)�����9�Yх�V��%Ǳ%;��y3yE[e�u#|P"ž[𞓇�~Ղ/PkHr�'�d��SXye΂�#��!�j-ϳ��ں��w	������F�tc^k��|�*�)8����Q0�hNf�er�)�6��FX�t��J^�[#����
ZM�v�%�������2�9���01M�u������ctݎl�1���*�:"����5V/���
P=�.ԏ����0�'(�C�7숔��pl8�`DK�dCu�0�g�	DV�ä�0+���|_ޥ�I�����>ɴ��X��M#�wY����.o.i�8�xL�ΌO2r�H^�M9	�5�ڠ�Mt�.�0u`T�3�5�S��L�P��$kL�B0��ҿ�X�D��$�<s.��p�������rw�Ш
�h_)�J=TWK���K��\�o#�e]m'>wC7�#Y��ԟ����<�ݰCw��l�z:�M5$!����g�O6�omY�S�teL{r�ȴ-Jt���߉�Z*�>�Vk&��|��yhH�?��u& �d�ܚ�,:�SS��K��b�Uh�e�Q�i�P ~�����Y^p4H�$S(�2{OPJ
�U4�\� %vU���	vZ�O��S�JB\�������v�$%�E!8��ν�!D,Z��I�"�������+������C�+�Qڳ�4�K��Th9���
��,մщ&;t�5ڥA[�
�^cn�`�z����1�@�ɹ|Y�ԝ����0��^��=�r�����?l��-* ��n�	%�S4���%DX���5Kf�#!`Ԑژ��얌P[�㱟�dk�2��Tt��3�Rc�[e����"�I�w5���^��|������@A���,��>S����h���'�k-d@��R���.��9�q��B�g�[P���ް4�zybw�u�ni�{�q��>XV&Y*)��l���9���\�}����+O6�u��m���㔉�|����('���Z���jbym�, l}�Kd����@I�!�5tt"�:7�Q50\�?��@̭a�~��ШeV��l�f��g⛩�ie�P���̑�{��5һ妇/ν��I-��_� 
F��k�?�s/�͋O�6my���2K������f܇3�ҹ�Wi<��B;K�ǅ����Tkt9'!sY|�N���7��}��.}o�L�-��蚣-���m"�Y�M�2e����"�<���ZRr9B�����	Ɲ1�h�K�Xm��L��pDƹ�X��tε���˅sVDr���C��9�E>Ɛ+(�a�B(�����`P�3:�Q����5�vW�1?@��qf��j�$��{�R�U��:�~�P>R��B�:�Vi:����O��L�Ϥ+#;m����R{�D�������'-H�3�Ht-���'j��s�����}����%���}EW��8�""����峅8�8_�I�٩��]�����6�&���l�Θwhe�%��Y�(�E73b�f���$]�jv���޼ű}���P|@@�E��SL#���9�f���֡�;�]�z�p�Ԁ^�*C�����k7t��4%N��䃑��Ή��5��>Xim�a̍o��D���M�rvӵ���GWw�U!Va�
����5 U�Hg�	Z$�d�(���&�r��PI0�RoH������LC�y���M9�.=c������,�`�x������3k��	�C��B�q����Ĉ�"Uy��
�f�� ��Gd[e����v�<�'�2�*�%�<|�����w�5=�L.�p�,���*���9;A���9╏Y4�E�,���.t/ 6G~c��[\{M2�RN��[�@�+V/�AK�:���q�?��Wz���/D]��
Ds�� ��4�}���tV=�z�e׳ ƶu_dr�^�����j����Ŏ��P���r�F���X����@����uV�-Fr�)�0M�-Z�5�<�-m�e4*�BA	��o�_���e����|�w1]�㨜�Ng��� ����F���iQn<��Փfe�B:�N"B� 1Ϭ�NƐ'p�Fj��cD��c�vUe��Y��)|�������[g�n���o��p�B'_>���עu3��Nq9?/�㾞!�![�"��.�>�\ڔ1���A��\u��p^�ȺT�s�V>����3����}�h�M�+�����ak�Qj���B�S��^\6ξZ��f��V�&-�L��s�H��+d���U�]��s@�-.��D�y�X�vh��F���E��#���-/�l�����F��-C�U���Ϝe9-��@܁�7Oy1�����'�J�?6:����� D�i�HO�Z�
1vr&�47����{�`����}4��[��u\�Ζfi� ��'�s�8룖	���RjË�'p�����K���\�)=�f0�ry��0��ZR��u��,�*û������JLL�E�NXX�1q �Q.r��"G��$�V�8������.u[����q��
�Mys�[�DN���p�Љ��I}��`���V`��Љ$9I��C�%��ȍ�k�O��+��@ӷ�SD��'�|,����
�����|�`F$=K��傈5�x�����4p���ǹr�i�R�$		��Q6���r��l��ߜ�0N�UQu睋�$�����p��1s�������_rؗ�#��^�K��9���R���G Hgzs�L���V<�L�ix�QXi8�GO��Z���偆%.��v[uz=0�&�Y�*�hf�\��$��HUJ
�?� �(�h[O��)w���U�U�<��zs閰�\b�K�;�h��� 6�[�u��3k����0C�b52���w��W��@R=k=9Ga�u͓���	�b����7�bn��j��B��	7�~W
]ie��H3G˸?�	ofAV
h�=8�L�|��:�A����Y�<��Uw�y�a)�;a�#�@ZT�9�kU�^��Xv�@�B�ie���k���9G���0J^��C���p�>ݗBx��X�[7abJ!��?�u�WVH�ԇ�h%�~��.�'�Ơ�(���@A�$Ěy�	��,�Y+)��f��41hj��{K*��\ x5X�����LE�=��r�g0���h�x�>Kf�KR�n��!웋���m�ٮ3!�cg��Y���4L�i�]$�Q�.�z%3O5�7� �(�T�\F$��eNϕ�v:>����t���2�dy���u�+�������2y��;�� PV)�� x�:+��^Be �{*v��f�i�_ݛ��c����m�rpz�f�<�C�)]�GM%�^΄u����#��B�����' ���E������r�>����~~K�f~E��a_��e�^,���G����OY� mp��~���'S0=�����N�p_�dč��~Y�� KR��<��d��Oe��ЇX�D^�����G �)�6�
��֦:���f��c�9���#��7c�n6�����Hq���#1���-�Nʖ�xZ�,��S�3 ���p�Y�Z�nt<���/+���/���SPt��Y��nήH��Y!�a�����>�./H�x�3s�����Ty��ζ�­����ߧ(��e)h�B�U�a�-�N���q	ӗ�JW�o���u}V����:\�D���;g���[¥a�[��|����ҏ�*y���1�����}���:�?|JX�5�_��W�K��1K�4�$���#���u�*�������Xٳ�?�����)��Б�a2^ <]M�K�|AѲ�v�si*Gk�[��s6�7x�9U���_\^+<�P26#��m�1 ��
�p8E�Q��0����U*� !�z^�8STt�T7���wa�q�E��@���u2��ݞP������Z$;����i�_miH1�s�~mf�h��R�'@��ݤ��)�^k�	a刀��b(�^�	���T(!9/%�./�ؽ&��������l$1r���)9��)!�������2#_�����WRo���@��s����OQ���Y9��F�dJ�������������{4޹�0�쵆xB���_��Ы��GK�J�qj�Z��\��r2�~m_��&9[�b��3q��{��b�9��㪎��~?�Wt�( �8c���VZ�n���*�V�����IT+P"��Բ���s��p�1K�lA%�γDg�=����l������"�)(�b�<V��*������p�cJ;x:�'�K���\�։���!@�n�=#���>�R��
�3���#h������ZS��~��/��.lU�څF�yL�:�a��F�f�'S���͵	Ȱ9�y�X8���釥��j�X��ϯ��"���(�ڇ�o��^O���Ds�����G�wZ��on��@�: ?��2A ����^Q"�0� �2��ik�.F)�Q���'c��N��|�	���[�]�uJ�B)��ӅT��
r��ܬ��2,�GC<		7��@qs�e�BA��$��I�Y'��D<�'�U�a��o�7�]��j;^��(�AD1�a�	��.J�q +����#T� ��SS��������)z=���d�Hd���{��V�:C:]�E�����dY��筯G��,�����Z�*��6��~	���/����l��*�L��Í�m��)�
r�T�N
�����m;4�3�ь���z6Pc{£�Gy�����"F�����]���W����L��^�?"�L!�H����CMN��c�8��(w����|3����i�Q�q��a�v�� �W�wjF&������Tg�G�c��Qs�0�}�3'�=�MB��uC���B/�[�����\F�* -��/%#J�%�lk	��b�'���'d���O�9[5\���-@D����G��W����s!@��XjקSN�Rm��?�A?��_02tؑ���t!��	h>?EǶ�Ȟ�;�s�#��jю}!����Ug~�D+�J���v6J���1�1�ߕ�XEI��#�L�p
 ��"��d�2��+;5�g�Xٕ�8EKCA�M��=�mo�a"�-OEz:���#�۔t��y�A@�&��������aWuX-fm��Iآo�?���� '�q';/F�%OlE
�l׌C�0v���<�#TyC����U�~���+�0���n��0W�c凹���2���h����/�0!�#}xU_�}�Ye�[G�S:<ҧ�?g�<�+� MسW��5g�ת��Y �V>ATX�3��D\�j*"��[n�b��K�j��o��$j�R�����=]��o����{�6��z��E�����ə(p���j��g��xEw]l7�%>"v3:_��Ф)k�Ϙj��Y��b�ΒJAveW�����ɫ��}`,H(��\CeF�R��!��H4�j3��l�5���n�&,j�)��su�T��������1$m���k�ȿ���� l��~1���V���@�az*I��)S��` M�F�}�b�*��d��&"�J��=�>�{F�Rgk}a��E�A�s93DQ�$��b��	(eNh��41���,Pg�F��CS'���w|�z��tN=���벯q0�X4�R�C���� ��bDz ���Kȳ8��/&۴���$�i������ONV��RKR����g!K̂g3��S����Ǩ.DW���4�fԵ<�r4=�Z�ֱl@�%f'���'�U��gi7�jpgD��O�
Y���E��/Us��1g�}:}2�;~n)V{iWQ��Ѯ�<t�2����H�V�#��`���]��ke�2�����2pB����]���*���`X�^�F�*=��	�Kg��}��i�P�O?��_"
Ѝy�^5G) �6\ܓ:�ׁ4sk��ԚL�����;�R���w¦�JB� _P�KPB��H�e��Z.[��M�J�`62z#���C+�����R��c��W��|$��txC,g�pnm6��)$�V�m�k*6a���+�2�n�sз�x�ʶ�O6�)_nVf-;��Knr�|PQt�hU4�����&ܽ�XTH#*/I�ʄ��Wұ�������'���|�)��J�H�����t>����C����l'�vhcZ������)�u��b��F�}�.\���D����hmTm#�������Y@���W����~&�yA٬���r���5�6���o,5� �J������:���ڌ�%�����۶w+<໎n�0@��j��}����'R�bj�+N쿇���3(�� �b�r>��Ƣ�5�!W���G����(����*\n��c4�{�������R��F��0��s�X�cO��bQ�Y�^�U��F!_R�zc��V̕lڪ���i|,�#��Q;�r��V#��7 ��N;��~?��Y�����)�Yj}�`�=VS�c!�⼆EI�w��E�8Hx�F6�������uP,��`���� �;�K�%��v�D�z�9�x���6�Z����?w$�8��a�_�m�r� J���1��I��)�x��90�&f���ViUIE�ٝ#bm�L-�H���Z0�������&,�0&�meD�lo�@|�IR,�0�	g�
��%P�]���"'�i{��pX��rW�O@���@0��D$�h�a�^X��la`��!�1��/B�z*�"8#�O��B)g�{qC�[���4��ꪣ���Ԃ�8�5?hB>t_�ū�Aݰi�@�;
�#!�$2��I�x����9�u���o�'���)�%�E�ڗE^�T=\����$�`�=5bs�R� (��Ҥ⦠b<�t2e�����9j�/��1V��<�<���{4@Pm��n��gY�Y�'����]]p�(8a�;� ��tn��i;mΌ	���Gw���/1Ӧ�`��(�b��u��㦸c�M!����.��f[��Ç
�o7"��hV:j=G�:���9r�0֊[+n^#<��36ϓ���b���x ��B�$`@����ld$�[���A�ۨ��\�C�r���W�p�Ћt���O�k�߸¥n��L��̼u�wJ(�l_��]�|���S�^x�9���*a�Y�˿�J�����r��39d����oA ���,�),	�+�btȥ�=�IK��v��N��Lg�{cۄ�����i��w�[�b^>��=�x��'���d8�cGe�[��2�";��u��V\'��;���N�q0�I.���g`)�Ǿ�)��T���DM����S�߱��+$&�֒]hgС:yl�d+�'MR�S�,�O����$���n]�E����?�w$y�DP��CK~x\�T��x�R�Urq��oΫ1�I�����8.B�o�"��\YY�,|�l�6��ņ���H�@��)]�D�>��|���T�kd��+ֿxIq���A}C�`wȽV�J��6��� �hF[��؃f_񴰜iGo=}�-�\ƕB��f��Dvֶ�2�}q@�[↼���_��"����^��:����6��}]���3�UĘ	���2T;ĺ3���`�7�^[Q�]&�mUo��G$�2F�a(ƭv�s����G�t�J�m����>�QH��&����i=�o�1Z�'������&7�'��!�tdr�v ���s�C��F6#B�����F�N�.���h��g! �0s�U>k9Jc��W ��(�nGf	/�$^����h��!ozl�1u����OB��X��xH){�LTAC��6�`��Y
��=�'J�S�8���kGq���ν�Kd9�duLM���fu��lZW���0B�:����b����X�U�f4OpN� eY ��u��h�.�4��X����P�p��U�`N�٨?\�%���~OE��f�3�E���|�:ǉ�3�B����1�#�N�3X��CC��2�����6���0��?W�gz���p�����z��j��No���n��I�ىt�ïZV���wFa����7w����ns�6Ҧ<r�����nݤǫ�$ %� ��-&�b���Z9��>����P��Vп����2�_��G�H��Mr���neF���[���_:w��')��ӳ@�S�Sӧy���1E�q�����Ѵ#b���@|���1[��U�1 �˖�3n��8LCX��
}}���Y��Ms~�7j�5nE�����ޖj;8ط���N�K�G��pyP���馔8q��� �$uG|DУՏ.�Vt��ݬGs��"i9�����t:��0*�O� WT�s�!�y��,g/��w�&�d�����p��>��/ܒ}�~Tk�?8�9t�"��5��������[)��{�,Уz:®s��;\%A ˩
�E�Ar?�DH{�|�H����?�ᮁ�5�_��B�w\k_H�����1I<|�n�L�lj��ٲ�n�-S���7�d����� �Aˀ���c����<�2��\R窅�1WW�^�&��Ed��� �s=`�3����٣'XMao��6�q�_�Z4ee�Z`?�o��V>����J΁RES�沨�`pM�\����Ԥ<��d��Z�rCІ��,du;qfo��V��%GF���
�ŠEe��+	�d��T�i2�c땓��	���vlKU��B ,I85�����Т����گ�,������n�a�������բ������ �+x�ۄ��ּ5Rt����R:��=��Y=�iqg�4De��sͣ�Jx���4�+�G��<L��PB9v{��oCC���Z�e���^�@��$O?�7W����,����d�Կ�qa�֒�����ŭ�h�����#Do�gKC�j��]�)�EEE
�E������� �V�dL�̾$��b�q�n�fŀ�&����z!Q|�H_q��C�У>�iQ|�.r7[ct�hI�R�qiO^^(�c�T��I86�P3u��I�u���v��+���to��g���gЗ�:�Ƣ�������a���o
���9�حb5�gbJ�|�=۠�7��g���a�w��+�d��6�S�_�ʣ���a������K���Yν�^q������o��!��\j��o��q��CU7��b��#�k
�N��c"ԇ�Y>h\p�xnAF^�AG�Gp�Io�6ZC��K5�d���oe\�����q��Zd�`��Ծ�z������M*���?&nLG���Bmzy�N�Q������'���"r�R ���S�Ջ� �e��7Yr	!�CK�K~A�w�h$mm�$�������ol�ލ<Ug1�C:�4�Xŏ���m��า�^gGHe���%�� a�飺%d2�X��3���~{Ǟ��I|�H�ه�e��i榕^�}��h%�;b��4���J0��5�\��ŭ�+��4Q�Xw�׎}Je������Y^���s^�ax��-��-H���,�����[�Į���C�i_s��D(�/����ܠ�>�w��	?@h,��;j�8�7.�9h��ր����"�l��X�Q��݉mfU�H�G�3N�_'��̗$t�&`��M0���7a�����5B,Vh�>���&T�C��w��g��?Rk�.�Gh�S�*}�e&F@�@�x�b��ue�3�Z$%;ٰ�8c:�
��2om`Wp�a.I��͜U��n��/�T4�XH�ߗ����?���i;��Q�ൽL`"��(f)�<Z����"��Xc�I��h
{$��E፫lH}��|���K����?�U7����o�à�.����чC�#n�i��q�BS�fY�+�!��!P�&Ǳ��j��-iT�9Jz9\Vf�}�$�g�W̾�N�Y��m �0�&�)����	��:����Ѐ��wt�)�C�*-M�IOM`4օ�L�:�%�{��g��&P���?��ޯN �$��L�����]-��JC�d����PB���1g�--|�2��T���p��=Z�r�6���j��z\%�#r��}1̀!ķ�j��}G�-�1&����ٌ�=��6�nv�G�����=KdJ�p�jp��T\k��Ѣ%9Ǐ�l�4A�*[��wc�nv��"m,}G�Z1����S��lR���+��NZ�?�j�D��O pH�I�eef-c����!����ǣ1����>xk�->�"�!A��d�g��H�zac��1'����z���H�09�Tk�� >���W���i�:�~4\5�����Qv��c|� �oҥ�5+:%d�:z�_pF3~^!���[�����R�B4�B��LX���,)�#��>��C9����R�3.dIi.�'��e��F2M����-X��,҂�+�O�*���0̗��$P�����$v[%�Į���-%-��4�.�����9NŞ�مH,�rzRr�	dy)�%!~����C'ۄ�.���Yc;1m3�hog3s��UΒ��+��m{u�v��,x�%��<q��Y�9$a{4�!�d#��hJ���]����[1ĕ�'RlB�����Z��%H�-KwD�G����Ӹ�.ly��t��b�l��Κ"��bW	!�R��ӗ %�ت$�kz�H��Ζ7V�mE�L�;�P��3z�#@/v�>�8.��~�?CW"����x�!�(��zQx6+~�@�PlZ1|^mD��.�����)��*{����G��"f!����<�D�XN}1��ખ{8��b����lZ�' �J��8� '���xPVR-i�
� ��چ�38�7���P窲J'T�=У��l��:���A�vG���26j�ʰ6K��A�"��^<�o�����uAD�����>������3��*A���@^�w�_�#P��>��\�Av�(��%�d~%g�7){�� �<��S[͘��6�$���	XjD!F����X��w4$��G;+�T:���>DE���c��<�
4���f�n:HzVY������_�C^u�5	4�`�&&"�)?D���6mo^Њl7�����T�p��ʀ�á�*z��1w#۶��#���s@3���$�
J+�O 	���33|�&�Q/Td�C�V�� m(�'w��?-�	`�Cm�$_J< ߎC� W�qD,���9���;�� ��ZC���sA,sk�S��	�gf�&��-����Ü.�K����fv�#^Hmߡ��$t-�����|Pr	� .�߃�ь�k�D���vwE9�qL�Uc��V_�x��6�a��SpWT�d;��IŞk>2J�<���`�:2yO��S�)L���aYj�+]��9D�i��K�K{�h���x��z���j]|�_!1�ռ�MAM��G��N�kUR��'�݉��i�@����r���Y�n/��p(��6�Z}�[�K�%�ы%�{�Գ4�:Y�J��e�o�4��k�:�
�U�*@7S"�`���������	�by���e=�|c�$=� �)H�i��ə�@�sA�����?4E��f��.J���ι�ExDcN\�&�\�c �P/Q(�����a�����fԟ,jȥ�*��JA+�?������<IH=�#��0���3ݳ��4͉&�[Akm0�K;� �<��ϠW��Eh�ՍT��>��#T:���˺�S`\Cs=��J�;��å�Rv�Z�;z\��%��@�u\��J�~��L�fs�$Ff��6��x�y���巶����f�x���j���	���[��8�}�6��yG!�������P��Í=ȡ�;�t?�W6���4-��:S�|xwgL��XohŠw�^��Gdda����HZ4߯Ɇ��g���;a��%���6�����]G/���DvLx���0w]No�����z�Cd��z*��I�؉2Ճ ֬�2��������j�㝘��,9��>�*�c�M����/G]־SZo>��1®iV�ٴ2�l����yV�#��Qr|ˀq��/��٦�l��'�&��1(IP��3+��o��A���P¿�i' kK��'M�N�	����D����s�Z8<�%\�:Q,�rO�)�o���q�!��3$ ���6��-�!�W�\���ʫ�a���s(;�f7�	^�Wd�^�2��N��JL�Ͼ\�~�B�qn�����g�N���ߝgK�b�w?�ܥ��-�[	����;���Y�������,}���CPB����I���� �G��%��M-�x&�D�v�a��ܰAn|��S:R}��~�<��##��c��ď�8]�-��qN^�~�o��(l��]#Ip�J�#���?�?��y��Q�Յ����~p�"t��9lt�*-�[�~��I�̦pl���T,��8�?�h��S��zl]JLP��SV_�F$�/O@����k���C�f��
�V�űD�55�U��@q�_,Q|�D������]����pI1����	>=C�uw"#Ix�X=�����0<��o���,�~�eOE	P�j䑀��~�4v��^�]/s�o�G.?(��P24�\�7�f�u����U/�
E<"%-����y����mY��x�)߱���c;pL��]I3xRHA��R�fC�r�(�"��3�S���,��������P�wp0Y"OViy�#���	�� (53!M�k}ݩ�/����m8^Wz��0�f�k̹yX�F����u���9� Sez��K��}c~�  �ؘfK��$iK���i�9Þ��)���ML�y�kʐ��`Q��oJ�=.���_�G�uA��^����U���n� IКU���Pra�GW2�L'��0�+d�$^A�5�)���-2 �^^OĹ��h@�mƺ2��D�Ջy2/2�6�	�h��p���ߋ�0��Q�͟&%��̡������f��9݃���}��q�Á}Z=�"�G�D4:CoA�}���3ny�oB1ed�f�s�w[�{���H���+���V��%
?Ӱ+�A=�L�:\vq�a,��Ed�N�H��/��e���������XO���yZ��=�X*2��N�β%�����7|E�3�o���3?�۫�? h�2r'�Vu�Z��n$X��Qf��;E�3@����h����uo�>�;�9B��Y��ͯ>���W3�D�b"�G�qW{{�>/�奷�k��Hʧ��/�[n�q� �s�)~�·�HF�d'H6_C�8c�ۭ�\����ݦ��94Vྡ�'�*u�w���f]�d��뇑,X2�9a�@3~�{6�o(8ct`�Y���ŵ�?o�Y��Q����y���2��X���c�1�<�Mr��]����[���{�[K1������k��� ��L�����!�`�-^[��'NڀW&���4!b"5CA��x���(tj6x��g�
�@�F�o8�'�����)���/K����2�^�Si��fa/��MC��79Ë�p��qq62���=��r��n�L]�8�n�g��<{][�V	��)�6(���լ����JdCR[l���AT@�`$�.P3n��?o�<�ԱT6DĒ)�A��=�	�p�'s��i��y�lyA(�'�+��[��Pu�Ytz(�c����{�t��ȧ0�������&�� ;ɞ�w�p�g��a�	Z�&
�8�tk��m��B����UC��"��[),m��l�z���2�ea20���Ө�M��bp�ڽ�F/hiL
�}���!x�	�wX���a���~�Z};B䴧����B� ��f�C���tՙ�)�&2��8MM,W��ӊ�!eވ�ִܽK# +V���xb-��d��mQްȜ=����$F�<u�$�`��Z�����Q�P.M<�S؝��J��^1�����wDQ��vq��dH14%�5��
�&L/�T�DM��Փ�hs���	��s����|!��3 �u����
w����'o�T��̪�@F��U�sE�=��R{)��7�33kCM�q
M�ڄ��F�-��� �vM�d���1Fp�q��̽�~}�(��+�q𐫆�~����&8T=2G��7K�]b*���P�`W�YX���K�>J%>���<�z�!p"
�7o�%�˾Zr=��6f·P�X�� �m�Q^���f�6�K4Q��e�b�\��Į��P���ǰhB�UŢ��:��t|X��=�w�j���l���S5Y'�䏻KC�LY��Z>y��[[b
}z�9���������$C��=���\���]h�pQ>hu�s�L:`Ï#l�yK]�j\�z����<�-��'$C�6��hM���3�$�m�@l#y� {�l#��%� @�w#U�J<`\FP�|�W��3��T<Y�y{�7�.U)p]���b#��V�13=<Bc��Q^��0S�hyC�nz7*�,I
H����pJ7�~Fa0���"���cj���>'܇0���ln���mC��8�Y�%;��l�C��٣8Jg�Αԇ���K� 8�>�馱���rdt�7��j�i��ިɜJ0��dՃ06�
];G3S;c�#�4����k���%q}�)_ZT�E��jqf��
��K�L�ߦ!�-��߸����<�&�q���"8u�g����tzvϴ��Bg���ƪ-^�w��j��P��ٺq �EVOj���T�r>���F�|E�k��k�QI`�+�la��#pÇ�(՟\dH2cE�~],��(�����}�w'%BV�V���"]q�u�;-}
VFT�!�ӷ���|�~QA�abq�u��5Q�O���L����|@�F(%pz�FmF�-!� �D�0m�	�ͫ0�sG��T��?U�*��!��DZ$����.̼���H��@K�ɵ�ԟ�u��Ƃw��2~ZX1�u�W���)y��[f5v��4�w&�.��UcZ1垮�|ThbB�>jv�ŭ����vI>R�h��U/0��x�@҃>5X��ײ9R�={W��St�C����Ť;��j����#���1+����'��~ 'Bd�4v'�k7R�}�7uO������|���P�YQ�d�-��#��Y�cE�����1�Z$��Igݜ�� ����m|`�S>��?]ҡ:����ϋ\�Xl��jf�4WT��1��K=U����$��6�8�w�X��馼Kÿ�@Q5H��ƍ���d�6ۖM�7���)2sg��-�,J\�ɳ裏־"�*~��W�ʻH��|�9��!*�
Gǀ�m����#�j��[�]��4�@^��J��k��S (�ځw����+H����^M��yc�ϙ.���f^�<��i�[H%(��ˉ��pV u4�v���G@��TĻƳ&��"):7�4��|�>��6��5NY��7����5�4L<�mt���*1�l5�����N&���{�@%��.���Ֆi���r�/��z/�� T���ӀN��aI͓��m{�m���vD^�,�s�Br�l�g�X6��(�����nB:�)][S�܏�
\T|����R� �7�6Я����Bf&��Y�/J`p�3S�p�r��!�KO�O�/(�<21q�]�����We��df�)�W��jR�G�M��J/�\&jc��
���7a!b�X��x9rY򇚧n��B�2�[�$�J��c=�(Nھf
�.׍2ʄ��Fؙ{{%��f9(�i�2<���x������R~���H�m���=�?��a�/^%��/��*je���M{������a��7���b$7 �"�卯Ԣy,_y��~x1� ��a^U8���ў��(l?��<��@q�.�l��RSIx���P�'r5��MtL.���x"��7&��>��!;��!���JV\�����pΣO ���C��m|"u�Y�I_�����9�0�8�1�oי�^Y)Ԏ��J��H������V�������L�m'�[~<c�H�� <�7�8�����_��p�2�)���m��go!$�x#J��^�gw:D������$��Zm�63�3�v��b�]kO�C�q�[0�!��'�t�N5�sc*x�>���M��U����$�`�Ψ�D`���S�p�9
u0�`���1L~{�2�u�������v,� p�E�"2!��mn���aU1����lBY�F��|p��V�DR��o�Us��6��ZiUd�P9:���M��,&�(���N��m{�D���׷�,���BB�-��t_��vc>i�� �{�?v?F�ZP/�2����J����l�������A/*^g��K��4m�\������[�!�	YM���~�3m��K0U2��P��I���t����LfC��`w�\bf-����d��r�>�CѳFlǩ�f4Գ�%m���>vi񺼿	B�~��fu%H]U#|���8��;�Fw(Lmץ�<�R'*�;R��ZS�v�Bx������OaȤ]?v����ۊ�FC�����85���b��ʣ_��{�1ȵ�����뇰��3{�)�Pb\f�gL��<�,붓�LY�40R�������H=&�]�$�u�,b�!6���c�an��N�k�8ٝ8��d�z��%t����9����C�3���B����ӎ����E����^��cD�w �q
�G�K�h5�������tV��
W�`��=���� ����}ò�p�Z����>�X=I�'�,#(�@Jy_o̟���29#��E�Fn�杇_�v��T��f~S���Բ.{W��/ߓ"���F�2|����ޣ����@�Vc;����O�?����as���S���Դ��p�|
�l��-�Yl��jE�HVt�0;0�͑�sv�Ov��S�n�q����֍3�-t���t�\?;�g_ҕ����g��^D;�a�h�u�|+\|kze �9S��]KR�36���O=Q�o7�1� l��~hJ�R�ި`�xV�(�uu�acRQy�+�%����Rq���N!�E�E�8�4~l6��l�	��r���|�EP�6�\��e��j���D��l��v�j�gT����[�����v$8�G��ϼ�g��=���]����*x)1�X�Ѷ��i	����}�u�c��`��j�V"l̜c�v����v�6l���b"����R�[
Q�o�CO���K�|7�Զ�}���h�T_�?��K�dE�w�2����Dp������A̉�ֲ�������>ի�S۞�#����zI>�KC��c������>U�ɧ�w��7��'�\K@���8�g]bj �Q:4_��q����[���Oɑ��%�J��n���k�$U&?��X��o�ϴ��}��<����N�ه�n�'��Du������ (?o��f��\���DD�U�rUKA�-�&����-Z �Ϻ.3P���ب~6�mgiu�"�����@^pz	Dl®2��,�?���H(|9��3v��:��o�]�95�v��΃4���cW�w!�ҋLi�I����]��o|q�'��=L��ƚ�
+�/ �D�v�#m5'���	�6���,����g��ޏintBj���J�*�G?� k�30UߑF>�N�T�����X�J_�t�|Y"ˮ�
����\߸��*R�3�����|e�}��餏pt^��n�%AB~\�Mݫ�1�!�領�#VM��Z$�+��� ?s��ti=�&Ҁ;q	�+v�_�|�%y*wn�����F�ؠ�3Zc�����}P���?�!�ӿ�=����w��l�{SI��Qd����ϰ�i����p��|VF�÷|�溭�6#����)��nϺוK�I�a)=d�?<,�q�G)wl�~�ha�:�ftT�\�U?�p���o�$��P�s��Q��o5�P��������s�N���>�/Cۅ Z]A�9*�r5�~�Å���ε~�c�T����P�Ù��]���9�ƱHW�@+(��~�XG5Wc�T���	��A�=E����pQ=��紵-�4\ݭI��&�KjV��������њ����8�+�-H�Q�y]��~w,��'m�]6n��vr�;^s��Uw�`q�&֟ǌ֓���ݷo�@�o�0b�/钱�]_4g}�*K؟����j�����d�:�f�`o&��RZ}����s{�r;,� 0����l�]ģ(�	�Be�y԰qG�����&��3��������#���!r�z�S��`Ԡ�q�AbRvn��>�I�`Q#��ݺ�3�-�9��a��Ô_(�� �/o������C��q��V�8a�[,��
ώsf����)UM���ֵ6ޯ��� s8n3mz���i���
��֢m`�[8ȥW�-�����~��j����M�m��m�.W��f1�t��
F|Q�o�,�������yV��&�������^<��j�
�yD�t���[��-S�*�$���;�j�cV)��&p^ղ�M[�i�����+�K�v?�8�n�m�k�L'W/��̓320�mLM�ab@�y���A0�` ����6.�r!���L��躟�:N�>��R�~i�|���t>3� ��z���` ��e>��q~��_��a�����~2vb,�C#	&���ӯ�m��^b9ZZM��H���56-�C�pm�tp3|���@�Я��?!&��^9G���wW���Fr�
g��fX�����AOGN�nۑ�Wa)�@�a���hv��?َ������V�H��VQ��+����0*?=�]�;:W�")[�,y�NcBi��U.l.�.-��:	�>3����ɉ�e	gD"��Օؗ\�Ғ�ZD:MQj�v������$ź,6�X������爩�^L�
ƍ�Y�j����ҁ���������L\��{Bz�j����,ƿ�t�y5��H]��¦zY�߯�t[f¯�NA�IC�6%׶�r^��V��ј�.@�jFJ�,`�~3W��K�(zc�=BW��U�0�n��X�q&C?�F���X?�;IiG�D�ag��S)صZea�IH[�O�Z-rc��q���\㉄"����L����`�9 y=��	3�`�٫��iޓb�]��2B1nF5�w��BZ"BO��ɀ�����Ć�6���S��i{)�2{�%϶���p�����]�3mف-?0�KHb�B{f�a�8����j��S(H�)h��H��]�$N��Ib0KT�x���n�s���M�-5�)�A���Y�����&?���z�7e�%],[�i�	6��_�UU1w̱SÃ�WYd�B�4]{�`�y�2�G	�����I*�,W� 9,V�kS��x���	r����(9�[J�b1n$��Ly탗�Nro��Z�?�8�
�>��'�؛�'�@��Cm���镋�'��s�T%�n,�$9uL�?ʭ��7�(&ǭ.pDT�#��U3y��^�8�"[M��Q��6e)hn�u��/D�G�T& �~
Uyq��˥E� p(��b�L�L��(C�VP+��v;�r�ٿ_�,�>Xz�UxB7YͿJc"F��h�_rj$n����6)���K�Um+:��t�(�0^����+[Lՙ<����<9: �{o�v<�� �v4r�r���	���<l��V����