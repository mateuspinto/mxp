`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8400)
`protect data_block
GgHqHSGa5L8zPC6p5UaT529RR2ZSLO0LYA4LffUAq5W3vpQsP2nUbHhWJ4eLTm9O2REBgsFJ6oi6
aQs3WR84Urrs0ns87i80XAILK/wzYk497r1DaNn/kYRl6I24e5NpjgfhEmLIntMTOZN9K71BK9HM
H5YbXyc1A/ULxen+Q8se5SomkH4e2e7Hd9r/eiBmnQP9ygR0wBrUk7Dr08BkPYmOxoDPBeJnCtz3
FJ4k+mt5Xn0QWzd2BijHKeb1Pp6/3Ze+8r+WBwPl50tR7SfMi+1wt3Yg2aC5ESZKZ8x7fxu392pg
raa8Y4Pjudzsi4M3KwE3kuVyilgaq1Tqx4A5Ffx9oDmB7W+HROYvRonrxI/WST1jbI7VPIsI6p/K
wZXQo39pDaOjfb7eRt/xp8/GntCXMZRJrh4yKFyutl3foW3CxKWL2WuMPpi7R8Du1cF8EkPs/+KR
mcusklfsx2qnK4uYIZDQimOtFT3UiR3r3u/DBTQsXQLH/RZhV1noDxutEY4TkyEfUG2zCX3kvt/3
rlSeIoRYRgQhLcYriV2n7ODbG5bvlDI3uUhsSOw80wjUx29F5toUDUJuu0Szci/f8vClEVqLddzF
6tRif30tkI+9tS9s8DyYi28fR1z3VAZA5YBfVjDe/0Ac93S7Rqa02QiOG0WDxRd+T2ie2etnUDPx
egFziiCm3JTCQkxigFp2LrOFrNUb1wWLiEM3J3/jl4S591yLCmipR6lpfQzEXL4qHezBNfT7nCm9
K6SBlnpLmWV5BgJYOK0xBVpbVCYfuGRm+UkmnRkXPgJtmYhXf9IOVgnZ3bkpB76gsK8b0T1eVvN8
D5hhHFuzWR//mK/BFH0LFxSE3dvP1la2i8SZl1MK6kCx/EA79s/re/9ulNmQvwI7ulEWKGQRv0Er
OvUqVbf/CW9dhP5VdWWwrmW6J9LYbqPhVv4MyaPLs2rV0RegSOWweZkKooMlHAcAUpVQ4Jq0tua/
4+FpxRdaVEb/2+jLO6X0YI/hsmjFzKys3ygKcs19sI+BoXOPsQIv7FqKi7ksjPY8rALj63cyMoQL
gEDWJWZg32TxcmZbQrKlH292CY04DV24G9D0oWBWNx/TA6VFJOa/XC9x2KO76omhvv26ILKdbJGv
SiIlnZ1a7nogEqooCOCovz5p6n4XE0ypw83T6w6XbF4oXMhRSVtp25yO5iJhvm/uMrC8dB9e4RFA
B74K1nI5I5XHoYIICE2zVNSLZYaN14lRx2gt0LtbemEG+UdRtquV85WOyu+0RXTzJ42ycF6CGlde
FFx2rSS/fJ+L+hiKCs63nkpf9jZG212zEOiID2brPogmsHTZlV4YvZMFkqiLCB/a4qFtMHoDYAPE
ZWIbGh2ErKtDmusE3ACmQS3UMKl6yJkSFXE9OaZIJAPQz77GLOBh5Td9e/+Cm9PjVk7JY1Q9V4au
OYbjYsgMFngYtN0pHOqyxe6onysG5jYPr6PLAXbcDu4fZRcMvsofARIdEVS0rghtwkmZ7ylOiNTi
F4rNCXQ6t8B4YHlKioEnW4iWPm6bcZS4TP82OGu6EYWGdv38RS9q24LicCmTD/EXIbyKZVoOU/O5
RSdj/xnluI9ExNSnbElDNx/DsB8TSyp73+iI/kY2uEuKpeqTL5Z3JQw6Eh8r05Y5My0TzJby5FAS
W8IdfpCbeD5jCeIvywirlrNIs2IMAI5+CjSr3+P4cOjd5P7xa9Yvg1zsXtjxBh2SotwkctDG/Dfh
1Q6nzjX7DmZ2SsQwuWaTbPKgQMj4tSd4BJ6wCGGj47hc1KXnOS0Dw8EBpKWaZgtaEPIFOUlTCQVG
GuUYO4k23L1PSBjCUM5X4HCvGh0OK1LQSWwSa7zvy9Cqy5T7mdadSIYB7i++lBqQrdzlWAqaSrLG
WpytAxK46hNenovlf2l2qNbNe3mqWJhCAzWDbomkYhCe5GbpEgqCsbQQfZ7LJ/m34ckywtHULTbG
8uNj/IebXwl2/Y4wDtbTOLJcqgea8TN8jty4NDfYZgblYhyk6xMV7wcKv72W2+B0dAFZs6TCrA9z
UtTuqm7UE2p0VVbACVCYfBTkol6pwBF8Wv7RhRiBM/T0dYSajSD40XTr/u+gTha3NGEoJK5FuXZY
psSU2m/bDI/7wUG1YjIhRZ7hQcWYfbI8hhFeb5WVSDLEYmU/AkeWMLV4fgdz5zfToqke3BDCm+AB
GZeATi9pnI14oR/RrJipbFAtTIN7aNJphP/1hDvSmKHprwbOEYNI+YhxrPGxPsPzM8z+v6OFMpbQ
VA2FLn1KmWZ+PNozqjgFl6Pkxqj6L2fsAO3jYQFCL+HShFP5kgbKjgLEvahjefURuEYMrMdQJujH
+5iAhUDISEF93nJx1ECmRdgCd6qP4xnSWMyYxBXwadip65ZCvX8kphUe5AkqLpgJuXnnrpaKHjzX
QUAcV/7RNoCAa0uPcx/xOKppTk001fgr0UQSrgePaEqWXDMBA5wFlmtKPy/8Mn9BS3hd4s7Ob8VF
Iw+hBOAFhF63jExIJFTv/elWEbi5fdUTvvkwZcHBwztqe8gB2mNkgLy3zLcsNjICPxicBb9tiAsA
NPT7UWh0EcG2pB2eG6iNQ9MMo3U3zOs8U0rJ9TlzcOdtWJi/snp9w+qnwgCy/wDsUrzoAp05omgm
iduWwX/Wwou+xoYQnjldNibB4LkhuOov81hrCkkUoH+RpAFV+NYjpLaWEwZ/ZuhxR90UF2JaJK3Q
QEMEz29ioVYKvsmDdnNJ02zdrIj+6LOo2fwsxhMIeEiVRCgiNWFjE2BGyQtkWpeYzpIzoogZAdVJ
tcAEKfCSRiC8xBklW8H+0GVA09Yf/Sn1Kmb+pnJzTe1pUjn56EriLl4HFZLoXKpcvnlkEDbqL3mc
MtekJdXivy+oR8u4p15+ZpZDs0nA3NDShxfNO7c2Yfc7QsRMJpYgezQWFssXQ2GH62c/Ezhi1z33
F06ZF4yt8/Z+lpRF/oRZrZvsnggn6LmwjoU16gQPArvPwjn9vNKjoSWBClJLjTiH8M4hIwss0RKu
FkPuIzhXIseQdWRJgLz9ib2S326CjhRxurpTGvC0pqjPtj0sy3mcXZr+Kt5qC022C3ilefCGJYVP
Lucj8IVj95ya3ES3gY0D2TPw6mkj9DoDUNGXXL/n/74jY3YgRYFqobAgETL2PPa8IfaWgIzeAV7L
DmcLbnVxW+c7sZ2LVFggrbKuKBWzkak1U8O8KLusHB5i9ZFpDD8cq5vOsoOOCsldqjrTcQmgH943
uhMnREiqoEQkMu++Bfr+N5qYyRDyIxWNLMU+qPMGnVx9I6ESiO1LI4v840iXqYKHqwS8o1Jri+AJ
VtjQWglW0yW592WdDOd3pfZLeV1oKbVC4uYaWTCdAP0zSssBagZ3DGkH4JXb6UiCxVsO+savT6JP
gmEzaPnfcOExyjr0ezdJcNasz4qoC2XPmEXgbszyLJmvokebuFeul0xozx2InD1prCy6dW/pDASz
ebU+kRY4VsXptWAZPXiogPiRGYuJXw3qwMnrMtcsSKr7xhONQQWmkNFlvhl1FG2P9yehuBPWlv8H
ItjIUrXF1AjsEbSI823M5m0PZtjgpLzqV7cEaL2SlrgOqGc0A6EUbMkUnm3lfUxP/tC1HHWJGcjV
ade/WZyHPwOmXcmmg5bdClQf+bLju5elMjtnjPnr4bzCxKmS8NiuJs6wJAy+FBAia2PZ0lhf5t0d
3HLqBPNCWnQdj3sf86b5IbQLyXT8w0Vv9Baz+Pap1lhKmQpPkcTM8LKZ8y0aHKrtZjmjmqI+S/6T
7BKgcqKb4a1W2ohJi6H4BDmJ1GRVhtiONF3vp8Xfescd8YfWOIuqWrfU7E6Z9Gjg7j0kCRqjbjRl
hr8fkynmZxgfcJXfmzuwrflCHTRVrWPL6/0IYLt2TFszWVeel0FdSSx4JMGv7wQSWM2GJ5BMw55l
V5D8s9YNQXTGsSd8F+83vN9UypVQjqtBgebAGR90BJc+8XDYlGYn+aQesiX4v28C9KzOngGav/d8
J2XfHVH52GIna+DsWZvn3TWiQd3Xa1DVA3NAtR3LmTud/qQVewPr2cwFlLOZpnNXdQdx1ttcnAV1
QUD/dHb02JMQNoR0w5TJFggf2ToiVNyC7KKUbEpk9S/E4aQtnGHuHSgo+Fac3xJAm4GuZgqP67Zj
nROEL1/1dlVamOhu9vxIpRNfQpUr03E4I395a769bDGyPrPzMGahLLi/G8ANzvXwp92Ao/eyYbaS
Y95OCmwYYFe6OkZhNemSR8dlOYDoiVMesXOsETAuEJPSp624+UTyYDO8Tg0DRGTSWOpKJT2FQtUF
XsFVNsqptoF8MVzucG1k9NPhsmB+WEvC9mCUiaD2JJvHrIC2sDmOrUccD0lAhlb6I4H0lEWzN18t
SDAZ1g2r6r7giuw2zjJzh9zF4fUtmPi1WmTCgtRkDozGjJM61SD9FTC19jrGAS5TQCF81MfSgPqw
ZrV0GwhvC95RT4Nnv5PLQhgWeS8BbCqgfXyUroeEXkwGBteDBmZubW1l6Jk90p0kpgUOb9NxolEU
zmSrPEZniVgZ24g++kJSANcB8ZQnwz5IYgCqDAmXdGWsgKa9416zrUof8i0RrH8/afyDlzVDeIJh
8bO3RNd/r1FIf6Kb2aADl/97WSUdetQ2XA0qhRPJhxQAS/01Y6869ttlI0AhcHE+26M0HvGH2/gD
MIx96zIJRJJfxQQ6HNNzPvIzOG8V3YbODWwOVzg0BjttNI70WGj51BrJMckbevNaYCaxovUwmXdF
9hPO6/mNPTGLlDvVESuj+XT6MLkveFdy7vYId8AmbS2qUt6dE8UDi9I9DXYc8+4CIGDCJdJ/Fzoj
RbEgdwHZx4ltM24VZDvLmQRqteZAbE2QI7ab2VUG9iCjb83xOdsjE2p5PVyAkpjpednEZeI3osMG
PYoZ0B6v1FZdlk9WlVgUFs1AnQLTbaKbL4PPHAFRz387VJZCGB6r5ZDuAhS4e1dOlnBiWJDt4QAz
LEMb4AsajHJYv0BJ/YPQu1fPkAIE2OtJtmi7EjnhFEsg+hezhQfenfxEbyBuk7w4ECWXhKsWFuYZ
DpukJUiUtUZPP+L92H+MU6pYGluJME297Tf8gLqr3Ds6ZQKiU2Ue4HHZn/X+mvNes9JqCjwxYROr
iKgtdwDx89hvjNsHFNZ+7TL6RSrXl1kMZvUaygKi8TaPsWmvpwiwxat2V2GEORsNKty09dqay+0n
YMG4hPJdv8Zyu9URzRJJ+paBzVc+nCYMyABbuyjHA/G9ca0Gq/hzV2t6zbVdoY0Qt6QtQysqU6xw
d/3U0hYJ5M8OSWySxSXDz7zr94UDpFd5C+lDhDMFxRItPJy108r2EuvuyY8I1R9yLDCacuXDIZYd
6a28DoFdkvpPRbthn3y7qQg0vcXatqzEl0FR2kyRBpGIbQ1kxu9j6yMzIjXvZ9VzvRiF34kMgtrz
02Jy4dKr/v317R9N3xxuY8auGmRJOLNFJmYWiUPyXQa0MtI+lRnjQmlTXDo6feUp+xYGJ4aPGL6K
uGt19gpZFU0LUtNhOxl3K1dPmYCMAsWb8QjoqIYss9gKepVdbpnUmVVHPCWyIsZpdxS+Vmu/7P6q
w5JDUOmhesPLmFu+pebVHQkuDH071m5AN90gUEKyaLD8JmLTqja5XKiEJunZ9rZilUKrAI0zYNJ7
7g/ieB6BdKqGVS+jC/iUWM2lTJ1NatexvJv2LxJnVWS07dkk2OIZKAqTWBD+V7bYOJMIRpvT5d5D
Dh+kwJg7zVHWKVD5tT2r0hISzpVrEWgQt7Pci/zt1mAxszlWZB1/uUD+XGk3ZVHCMwIJqJwVsxmp
N+Epx6FOWuWzts4zClz08/1YRsv6z1uutZm7dyvsRnp0LMsyiXqVUIcNRNGKKBinCroZvSsZOAws
d8Nqx7fsEVmfVbTuSQtJjoi/Il4A6/22r6n7HyNAD1eGRKdwP8HCxA600X9hejBSAlLsPmvSpB1h
MD28zlXEQsUshmUdA48BVfcLQM6m0Q0L2ZygR6y4coiKpr4UeHFhXf9a7bFBLqprZ4ItCQzEhPbI
g0I2ky2Y2zCCqt10sEfEJs6tHQ05JwrwUhRzBxSoNkfMvX4zfZyC20sKTRR4edT+JE65YBQ/4uKV
EnXPUYKrOYnOOieR1sdn4u7KhUQnT2mH6Yx+xCwNGJ+W/NkC663M46uJhlOEVTtOUcv8AVVsPZoC
gqbNuHQXC6tqXHv4Jy2cd/ibuHlyJEuYFYOjyMtyXan1dxf2cdHzymZEln2GXS7K/nNB5Wc2Ca0o
byTT30+wR1yg6Q2yFw0zrznSlu4zDQvliflKkd+Chj7Y1Yuc6w39GKNlqMXaaK0GCv34J5zMcG/4
AdCKKk751hM5gEKmnLwgqjr7oRqnrQptu33oObN6N6SZzgWgg61PGz2gb+aQxMiYaq1w26jS094a
s6fUQSwVMLaQygJC6Osfin/GTVuZ1ujfSx/A0P/gGgk9x2+v636xXaT2PcOTw0a/vkddEmWZpGIa
oGVivjuk4y6ipa/y2jTQVxLxDKn9a62mx/J50reWzE895IlxUtSkgqIzmujQPqgvVNJnTeSeA3fZ
zxbfM9Y0InQ3RojNViLKmhD+BDHYG5Iy4qltGBXPKp3xP7XDEn12cspnbo+Gugtrg64uPmtNHicT
vFWJIt7Hcvd0snOuD5KMBbml9zW3Qzv7s99UBw1HW7sLRL6FWjm4kk4O7OVFajsOTY1nwxhnwyoD
lxuXu25SQfRtwCLQyg/5doKU4uCzjI/c5mQGSYIQfUbwtVQHkR8ML+ZRpfjD4ZQ21cmanoj2Bqod
bRmhJFYGu4cpR79zg46al6nCQjb/BVShkUAkW+cfjQxzorZUi46Yy103MRdLWQu5M0vOEFwaDt1L
uocldoBJ2cNUscS+I6YG3+Qym7Sqakr7+7qx6rBlFGMywrM+u3o1QEr77Nt+SLndlky1emHLa+wG
YHg23ck75xTMl+sQk2LzDmAi0HTwc/2QxnxtrVH7o1WmwxPoUAIwLe4RzK98c58DrPRY7NBWkCAq
mMgWE5BHdYdEr1ITGfzFFlGw7pY7/H6xW2NqJnRSm+nmKxh5LzZzDsI3McA2uWJFmTCj63hDb0x7
sqO33if2L29/ZQ1TPyCa1TeNjeVPdRpS1EHAhmkD1ov8/wmaxG14FnpqU8+vXvWCNZocDYQaKrkA
5baC0NH6ESw0K/iSs4Aj5Z5GyjL4/2FuE6UssSAtik8AtLNuubDE8b2K0W/xjstTAs80RDCmN0AK
r0LD2QQ/C9Juvamv7JgdIPLpgCUPuaSZQTQ9PYWiXy0kTe4yp7Sep0jJ9d27sFpFmvaPb7/2Yg1S
W9K+VWlmd0rbTQHfBQnvZBwdrXNNAsk4QzYmH8vAonhcWjxnStiJHjyyWH7DvLZpfEU5KY+TCEmi
SmUGMpPGbxojF67KOUeIkTTZD2R3gidssCWgyQFx2DlZjUkgM2ELigfnGdQWoEoMefwYFMAFueSh
s8aTGPc7jdtxkNXzlKU0SjMl9Cj1+4HACuQNHztvJlNtm3eSM0qSFXxdOn9qysYZHIXc0ykZsbJn
AdTEvR9CrCHm08GLlsCJbtqxyS5ZDgCF16zXH6GWoFX4pLlcEX/DWK8EH+M4a7wkysO67d0CjMXf
/LAWYK+I8SvbFLt9spZgvCfDyjvGbOzA+58eVn0Iblgz0g0m4zg39Cq5My3adgQrUhIsctmEz7mf
uzAhXlqfz4c7+vsTjh8R3dX3ufzRsVz9erxT88leNL+WjUwUv5MSQWPeHru0yUqSFkOptD8REP6O
TK1zki7ynww4ISiheat0NUHnbzxDgharyUDR24gCuj/ieOtAYxJpS0vDbDFTChxjBYfuWzKQeW9Z
pUCGlFyodrciS31HpFvCBWuVZnTCydnzgskCFXFg5O1rFrFGinqY3Ed+C/MxF/E+2aEhsdfJQnlD
tM6SK/tNaOS/BfgOEG9cVH71oOIDWwEelbyNO8CVagpFZxGuy8vNCcQ6jrk+sVwvnrVwQf9hTccq
4SG6qgNua9ih6AXTKMwWKpSd3tuzIxRwuxgZRHHj4PIpNlIk9mD70TpmZvda/POx04l3lss/a34X
i1Oi1KnXDbXkBuiOpGGBT1cmxb+tg2ceWA1LOxOOIWkd3DcFBxuCQdveKyWnrNDZ0//4/AIiNc/i
crTb4ceD6flAb3dOAmiVTZw7jUuQYoem/qfYjiRMaCzQqnq3ZC4HwXJ1/F5CHNBh3AAXmLbr/uyX
HB+9Pp6icg02ZWnjLXqzFXH+dTogHnCtr2g2IhxH1HWTim9xcwVD/rmwbxSryKgF4riA+o5cSHOj
DKiHkSKw1OXsbZ7xBHuNhjAe8qro0Trxl2aVUza5obxpuynwHo+9MrvV5Y/HTsG94ZkXjKwP1jht
ROjh7m2zzidHeSRKr90K5D/78/D9XKyAJhk65zLSO73xEGAtjgmH33f10RFC7brZLNOgOFO/p0ys
NIisYh1W+sCA4DTUOPjjAYvBleGMMslbV/byEV5P4L7SWH65WamkyG2ReiMXlYVI8cS6iNgXLHgN
Wy+WLLVl+MGf0rgmzcpj4MgG1Q6Jag3uGv5MjLLfl8rFZ5urUPjoC+xJMfLRNzSYU+Ip0liE9H+u
MoJCrU4Odu+oyZjGLTderj2rxOfKhd7pWNbH6isewGS5io46ooYsSf1KJ3dqGftRtWEnzgMEVWpo
d2wqgNK/DxO2stl7HQD8QLP+l2QwdqaLj8waH1ABt6PiWehrwt6+XqQII5it+xWgayq9kMf0hZZh
jx3Wz1FnX1ewljIX+oEeuy9iZ+uASmwm0QJX5Z+XBEl4VeyQyfsnFg6GtBbkntMhrZwr6fF74UOH
Hf2KRCq3HT4MLn2lQ+fzwp7AztaDsyxqkXAn//oda96gYNUVXt+5o/azWPMcyn63MVNG3z9T3l6e
ctK4uDfk09e0o425w9ySZ3gbnqfkNXdjsb/b8xHmSKnLE0NJ4v7SzivhWA1fTPpv8mRd87vY1XQ1
nC8AYvY8n+Dc6xNtsm2jf5PLcZCiFFenfVqNk+iA6s9gzQfFu7s/DmHYB5jZ9M82uxvKwzkcFHbN
wZph0Q8hb3yHgWAmTdO/33ymCMu4oaccg1smICFuGrCqYnZrHMjcbKjiRwow5kZbsElo5Rg/gFk4
bNtQ50Xq64G9tCS6DiF6H0bG+tVDIq9AaoDwSVzlICWHOUmAHe4MtgD9H25mTy21RvY80PhizkIR
yR8Ix5SqC0J+Lw/7qAIXrXgaC4MVc3gLW2cimyJ3w1nOApPHVlx4gxSSLI0njJIFoujrJKj1D1la
hdOTzmV6kjd4apG3nu7qhTIrb/TSk/GKKQXATAVx6nMUDmWhWfUrDzEGcjmpn452bHkRLlbknsHX
AbkhZMoqhmvpX1qi3QCMYe8AEyzHloPX2xi5xZ8/mUCN1ZzFBqxyKKG5wiTnZGtZv60ZwOmQVEg/
mxJrzxNSCom4uCC/eyDySomhQaULmogbROM+aYmM0Wr6/po1Jv3dbK5cOe2uvBdaLsWIyxaILb3a
3RurWP4oiTdp5Wlh0h7wbafgRkkt6GpVGgodXMVot6dL3YI1M+SqBy0EwKTu0KTHrxBkgnjWgwwB
qJ3e50oHaR99BybcXLBysPrs7uAZXJrY4Kfrc0bxAsztJp1yLWAn0dWV6ESeD9uvtkk0GEBS7j41
KV8GFIBTLd9FygCyADjFCWVTPdtWWGk5ef8wh7L77ey3BRn7vkWpK0Fuf0TeACPndmifbIxP5qZ1
jDmc1gLe6WJZPNUJYTNSzJ1KQ67/T5GNCVQ/98vRRLRmtRfe6uv1JxhPmtMzJbV8VdqNa7aLO5ra
EYikxm281GOkTG/uEqwvqNZJRoTVDAR4PLA8sH9upkDgw+cWB9ul5L9/EQkUlMF+vfUSjm/uhYBg
Nnx9eK+/R8VBvBe0W7olew3t2z1ETfyebkx734wU4gWEWmKU28ZkLKOsIl133vQFe843kO3W5VyH
JHSiqBuWArJpnhj9ZG0vbeADZCSYV41T8QBwkAsfI4vWV4xf/UxxhCEmhT4mjX9nmWyp9+c77YjP
Ksu/wR/o4qCyMMcuYhH+0v7CYcILrR66+nVEMsG4GZBeqBiqf2JHKi2dWcMmM3e6k1EHOUDXcXs9
KEZkTr7m/34Tf75n+6wAxtGpTEbZ4TF8EaMml1wjEZQrP2Id3szIUoJoxSgMF4Em6M8s4o7gPDPf
BkOfakSm1pxcXjqLTMfNswCAONfXzyLDOYY17Cn/pG0ohSPNnWRrFZtz5I/8cJktyczrNgEugslF
aHHibYMioV0T96hmv0z2NJ7vM49UXfgR76QLaT1QIePNMs+HubaJrQePLiMr2D3k29py8aLIxkNu
OHfZNbUZF/3eC6KSr2hg571bm8lpkv4JbIyAP1XvazVmfbQlmWe+l+5tFrzt87eGOcJLr6eY/g1y
HFf+b3f0sF84rcTbEgVepBIp0H8LdnO3wWf3dBIPI3hvdcFwADcAHoxbUjrVs3WnR5HBXsvN5Ij+
VejKXK0i+VTSYJ3JFiCeQ/aBQZUbXdD3vUqlxp05jByjCTVuKid//ceTRqqeaGhwfwORO9yekPls
bPURP067bYRz9c4oj3GPYIYf6LIoDe8DfHBxWqzp6mhTHmoLqLC8hEGY9vpoWR+OTHSncw9vCfWS
E+SvmYBVGVxsbVQwP6tEd9VCd9IkUp6S6giwhn7lbabokit1gf2/J9e+WjjMAKt4r33C9iFd5ho7
9hAPlJFtrGApFt+tpGzbLI5zc/XO/RoVyJaRH+iR4NOg1kixAkWt6ECl85RJxmlVLZnIVunz4JN/
r/ksfKSRa1o7jJtwsORhc9/LtiGm8mlDAC9qOM2RjJloQ6B0is9DunglTZ9RW6aqXE6ypszBbzal
XFb3iZEtJa6/YuaW9W6FbzWYn8SoO7XWMODXH5dzMLcmaqTx+W1aXdxhkd2zjIXzioKYymw5RGxl
28kN7fBHFn3h7WJVXWCTaci6vsHQ+TKXDPGTewihPP1v24OZIvxgDB74+bv+QB01ly9KvdArFo4O
5oEs9fRI6txzZEMnebDgj36HWTEvrH7r6i8qQ5s4dwOJ45ZGM2F/msqZMjXx/KE1TVwV7GKp4xpk
JfJeOzHbpwzyyBlufs7v2WUZ1eiY
`protect end_protected
