`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
YR1vF5dYUOh8JcukEIx3gvXKFfs3Y5OKmZ7hs+mqxzHFnAlfoREDzo1rvs5LL/g9GXBv4bfX8y1G
YL3aW7XAusa2VpVQ6U7hY8/KqF89AcHFnsxTSGarnXaIEMYKoq7zLzd9lmiks/eLkq9yWD9QGp/8
ciGThlqKBhj7rEdxeHdYVzqS+gmBLfKDemqizsdZHbH0u/abbuIkqbx68jn+qXYtJSMjMTAFQkvE
Kqws8jAT5tDukFGBJF6FG6fztfQzxHVDrX2qtT/chjsrOCZethR6LZFUEAUvbLdA4iNwVEQfWiM6
ER8xJH85P8w/6FBP8N9Il2Wt2ID5X2jaQ68hNA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="lr+z+RVbUqzMJZikBzp5kr24vrxjlIK4KCOiD0JCHHg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 77968)
`protect data_block
kYOIV6nrxd6SK1eRom0JB6e8vIv4ZOKaLUvXQES8G46oqzEFwsTarirp9wksNFVs4nPW7RnwpEGQ
tAyiqZbN+Pr3i8gLT8wD0EKPqX9ba1nePTvmovZHPLd2PJu+Y1w6UrE8f7c6WbnbiL2YcN3MlQGX
nK+8ZwJPNEAyiYUxV0WOZxpL+1c6xtHp6FFq8q63vgKK9zggqOopQ0yctXLWn7/F5ZA6tzUin/vV
v3ytsT3LA2CRPN0CNXhAQ3f6IulOeKzvZ1XWzYnI2Cyz3nyXTlNGv39ogTd+1FwISEZbLYCYhS12
QeFYtu8OB9cCDjZMNzC1nH/vb2ue9+PDA8q048FYgk1UIWscRDVFI/FmEPdqjDs2W35dPAC83oq0
sjh78LEIvCYD/vsZ0ol83WO9NwJlC8fC60dnPNU7sWZ94k7ym19ccBpsF52hwViAIElsGvdB2plD
tBEDfwKYwC10q17XvkRXGKkjJA1RAVmpqYLgbX5V+SiAKk/DPU6pKPygjvpbjiCYhHSf0lhuKfkV
D5+ZB7Rt3OHThggjZmPYofIss/1ssYUTneQCyiznHYcd64bDVVImTYWDeXbLyEhqdS5teU1loDMp
WQBf5xYm4GRz30ysUhslEStVqGzmCjvzalBIM9Pgbr7GcG0UCzndnUk9I61P+77d9Vj99YJXrqob
iFcWy4Ib4wMii9yEaNFONusXmL0+RtYvR0FeL9Bfiqe3FLmV+Td/JKmRR050+F0qPujhb8xr0K2b
v3TsCstuvngUV8YDJHvQCZ8oyQsEdDMOvkd4iOF/EJ3HiRIQXlPxvBmIEqhu6FQnVjOc1d4VA7Wm
LukcivBhLMcGGsKRxdQh1mp77fihGkJJAkrOqzFb3PMK2vJmN1QRvRLI2kkgmurPxXh5KL0oaH8E
Fg1LrHn87nNWh30kFRumA/CI+/NOJrrd4ng1IV9eR16eITPy/ujSSZViku9pynJaS/L2wzn/JZtM
hJjqpmWnFP2+nGlDHBbmRGTNSRtfOy7kYhIqsnPtenCFv/1Jpf6OrGi4WOeG/s4zvu8XrGy+64Fl
GRY/niiVRWwuCgWjRlkZ/3NDhRlYMUTZNYyLA7+vydxk5KfqVM1GwDU0xXnfC4A0Nx2Y36UDX+dO
xpbGsHthUO0RB6sRoPIJ+Q00XP5HHcDt0lpcJ7Y8+g+pOntdU91FEeBBHCrvO5WOHbWGe7Bjx6hx
CxVeS9AmXCSMBuzJzLROSgUqNpq9mp/3c5FP0kc1SSAF1qrXJGXKUcV0UUKxcBlVvROZaMNh+xCb
WeirVpZQ+sAsY1ZknWEV6heoDPj7jYpsPQDym1cIM++D5jNVKRXOEPzmSjzMAec5nz9XFt1+Rqgg
ZE9DcjqTPMsJ+T/0/b/Acs1/dG15WIkw59iueN9iamp/QqIoc3Esi0e5cpvNT6i5uDWwc3SgWeQH
62hq3sQIldV0HoNGzBb1zOe82UkF5PXbBMcAAjuDsU9RFdAVIJosOzP1+a7w9pbuY8wPg7efovvz
uyREbEd9x4LJZ6SlV0V4spOHoZoxE1UfEfO9GHiOgKG9Lq5EfzExH6i3IOyDFZcXItoVwL6mtvBM
z9/2Gm02YNbQQAtuep/xcGc36sNc3VVmeXZ5yAUA8g5MTtxQFi33LU8jNYWx5yEGHM0RXzrhoz+r
3UB0KMbc63fOjnvVuI+3wPgeKBUHpWkXfLa03yIY+4noo79Uy0Gd3gaoIBhTo3iMZlpBzSE66wLc
LKpbMgIwrogzF9dUbPI402hw0iVc3lzxhPWQ8NcdQ5js/gsO3VEnpl4PzIPHT62RD0u+kxGn1Ld/
vje3HhErlw2YQrlWF5H/flMbjtcPSZ6Al2Mz3fTqvazUe+Qb4iuYC8E/eYAVPWIQhU9P9mg6OJGE
2n+SQJE685jPwmtO5A+/EwOFJaanVdPMhvQsHj/UciP3ciTK8id8BRlVmx2Et6DfrldlhVvykl6B
tK+B2ZhVWKOgm9JHSPEHDxBqBwxuFmxCcwQJFVEG1tNXRKwtsKhi28lDy+9h0wzpQva28ewja41Y
5jHkMnOgEs7n8dUpm+fze3i9V+KujB3bTlBBa6yvMXt9Jscl58NIuw2RLl/3EFY3U06/LnNAkvIy
E1tVcg/poLpSZuuFNeJsszpbYUFBRvONOd/GERGmQbho2awMYHepNXZyjCHbNKdq8bEjsTqn1zsR
wX3PN8yT8VE8XB50CdlpeH+Njy8vrNtOrVE0/slfUOir+0Hr3VRuca0DacKvcfvEf2iV9reS/Dof
/Fw9YtQ1SiMWC2AdVCVTS5D+Ms/qykgMFik77ooKua5RwDg9Q1GilSWP+O3sSUkBDLzZtPVh6+YH
djMlUBnkdvCi+YTPZDsDoIqeSsIVxnPQDwq3FKjpwrpO61ym4RWHg+hDU9RxFLBwovpK2m5zxZSt
qOGHBNcaQUfL/gEHRMDsmwoxTteU07D2O7v8iooW0gHRPaFqtcVnIM4LnGCBC23FsVud3rEu7G/4
rggzlFTqKGYFO4TA6G8T3sf5RXy1whV4J/NyoMBMOlbKVyGmVL7oE8v2k4ef5nf7OjLFWvZvRvQ5
SAjHwtuLn/HfFotGTUGPSsC7ffXCQwHKP72c5fXZrg565IIe6ya/HK8cPqrR1OUPXXhz3tnFzsw4
1vfwB9xdW+gNHE/K01oCluxTq0dMiaLS194T9ddW9RIApFKHr3E/PaZVIpOriy5N789+SxWIqYJ0
W9GUcl27+aMMO+hgRfC78Oyxd6+MZkwPk+J7iXGZ8vJoKI5UyQyy7ASRRHOH/+R40MC9J2t74JtL
eIILCZlpF1lIAUQaIDc3H/EJ5bfokC8wyV2FfArB/LeJQlR63FPHgTZ30HFhLpxvVBbGjtgozwx9
pZbSyT2HGnMvRjcnmDy2pZwoCuA9D9cnm4b146YxJ2OYdwdWeBeqaIYiGaf2PAhBGmqHtSNdTH1C
hbF4jG7jCciHfhqN0zMxoyyaq6r5OWWybEYqLK/jL90+cueIZL5+bQOEM2kA9+7BgPgN481e+l6E
ZhH2iKQZ01PLkI25DeQYD0QEE/tHLaxKXJfaxxwrpLHErfk2jAJVjghw42GJervqzm1TDO5d6InE
1HWvroZxFB/RbGVF3uB8Q60r75qwfQ7RyqQXvPfR37/By15gW4rxFf8ePLdrIKHhckcwC2IFmkqn
Zp2reHOKoG0vAVRwyJPqZk5l6Ax2TU6gbtRhnw1mwuOc+tyf6uKzeYogW8PLKl1slViQGt7IIpLw
03SoWsosL7v1+2PVHUJVerORu372LcV3YRGA1cGAhvyhJ0ELnUYO0p3HaSe0TUOwKVtlld4bCfGE
GABogOfM8tEOqT/rFPmS4BEF7jiYX546leAzOURd10qQihHVyTBJ7FRVQgCMU62RhUuahRqGjj31
LaG+xCpssjV6gADnjQS+IQFeIax9z866+GFuRG50JlU2s0pKzWyYEQMNyBPfayi1aRSMd1BVpd8J
ZIX6ABwUi6xrVql3XE7dDpOaxYcN6SuCMBZiVlJIGKa+uDxPx43Aw8IPsxy5bR6UbZwCHBj9/XCv
cyhwG8HQfDHSDTsm24Za/JJp5KD4LxSQ+qrT/hU/Wr3+JmjlG0Ugvn9tbWYqdBHuUZIXUMQ6Ru2X
7xDpn0LGqLSNODLdvVdtA4XkANvhbnrHyf+C6kYxrhvKtD6HjaV5+u7tRbR85EQpZ4i+5QKC8/g4
1cPHiRbrePuY1eDjQAJL3DaierCPt8Ua3RRNL1EvssilFDfoD1wi67Haql66gIZrThRDQOQ01sHK
wQW4CbcfeMwOAjKRRYGmAiKZrQgkDTMrizVPlHGyq27pFvbWDpmO8bJgHtCPFTdJaE1zZOg3yrri
9Zu/85yxu86fvYuyqhBEAqN7aeaq0YTtncI99OjMq0NpGOSEuGde3FNRFRJATzsAdgY0ARo7vi+6
onPXWb41w8NXMLS/mDdKJv0Qe9z0vuArbycDA/9BlJ/Lqs1cUGT2lrZDw5BDQlrxTC8RuOriI8vZ
p+HkNLvhZKiHgIsCFRboq+XzEvxpqfRo9VT3dUyXBi6xNWPKNgHWXPNMnh9bdfV8cBbeCYJszLER
ND1IKbjy4YcaRdkTyGbRE92cCHTs78t94ZL3r6UxGMA09eyFlqNaeEf+Tk6/4n1/lWLaxvIG906e
x2MgnGmGYCftkOi+kOWtvYlQRgi56YmBwszvM61wl03gJUfyAYINYu358QDQApvXNEFV6o8NsFjz
+xCbZ5IjC6z6zOHINRsJivmd+Ui5OPUPI86puotNGzY17biix9vK/OdO2MVhU1LNsIVtAz9Op9OC
K5NkBhUmTcr//m8abTsldbV/ly5BqPFWzb7EPwW4v02GT5CpnYzocQHwHyyjXht/9RmqrUBmcGpu
9hj/ZMT0smEufDI6umo+uGOWZKSfvWmL8ZkkdmNQfeYdHyXUp3B7/xpN4fvgIoQd0S9Bc3l6Av2/
R4HI/583Cc8kIaVUzgcay/CiTtRPKfcQQSRYyca0ZfkRrq3OvJcHI0q7E2GVA1WSsrAUNoh8xCkk
kZ/QTA91vlzM+w5uTUbCtCF8Jpdg8OtmFKLMd8gPwaPg6v2ZeaVp+b4Py6ynXRMziWlluWu1xPuU
hZr5uqzm2Hf69BlMkT7YsVFTUAxP8vj4MsprbI0BXYQEtCtiIPKMmSo7iswOhJgC9n9VeH3kYjsT
RocuKLvuxOfB0t90H4lIuM0X7SdZDzR7KxAi+xrwTHZcQrC2EuCkKncyg+MpORyhfblCgTvFk6Du
mAatyNRXNGkZZn7NUAr+ScK76lHypsRNHS8pAVNLFgj656XQRcWWKkRsi0UkneP38rgg6WzkN0PZ
tEaMfFEYC0xi7N5ZfycZsDur0uDe2LlyxFgINmK14SQwhnQFy7WFF3B2Bt0L99+xIen7o7LrlWcz
MiF8x1IPP+nlz40Wg1t6MF08AElI21nwmk/2zNwBI2lkW4O2ElRHM/1yHhEXkRRzfyAq0sxP0uJi
PYwN5xDFEDdNnjjot+9fq0NDTnfXwb4j0HqR8RGoCEiMz3ZCqUq9/H7nRBp9p7XQqyyjKcOFsw/S
KtnlefhnO8A+UtrXq5A3QTVM2EXeilPwhyBLCF3a/mYAKdX01R3bg9rQuq8tT4ZV8y49EUh7wHPm
GrIOH4vLOvDW4sYleehH69nlmqg7xFdjgOKQ8X46G+8eFuQFyf9Cnpf30hW1U3c0RexHf9Rzq/ii
H8bAY4IyC2GEzyK3xHiDi+aNZq/tl26HGyV+S5PsqfLApfbD0szMEkryKvl28qX7Kx1m8QMEYS5l
QBOw7j+yBf2MMQv0eAjVL0gcFkDp60y53ZFS3GOEM7i8/xCp5pnGb/xY4kGIMcZ3yXvd/L+H5KER
JwjHE0wHe3FNdi4+i/qcZ5umFsyLUORAyVvk/07PnoC1jEb5ytXeZt68Si3uL8yW30oou6GY6Dzs
Z3Drn+UjD2QmNFySjgcSQyH8eZiPrOkm2pmRCaHuRq3RjObC3kTmUFPgk7G3Ou+DtbTKp9megjL2
r1sSm+B7KUd9+40Kg/8CRvl9Y5Vxb0vgBZA8uoBp3X6PcL6Wu4EA5ek1JLgt/c6V6ycmMYF/RbUx
tkg+hyGepr4KzOdY6U5VkgGMtzzZ5555z+JuEz/Ic1QAdCXD8ZtjJt01zJRRNsmr4FGNrlmMSwZw
/iOnOm4EvyiwYSZ65ajgb0gaBzSpTGQzXxXvSdHsoSKKZCqfHr34Y3FZOlYUXKE0jqoTOQNpbv8b
VnffWGRO0lr5/eu2O/QDMxCUgAhZMbsYA0UE9/It9Q1Zcchz/MdwOvVJlVJBo/7e4KCh7a+CcAaL
a5m+Yjmn67dNIVuBAOdL+yGe2mHowElbUWdrKvZ4gy/u7xq6AZ2JIBgl87tDR8jgotxHnndrM67P
6u41Htos1boJT/qPBVU3vSv7eCZA4/8JkwX6ylFRvCu3zj1KD2mbKQGtuQNWEsUYqedgIJg0Uxmw
MY8n6Um8L9nLNfnlMjoNHRfKEZjmbLeBuFdR2u8KMCyVVK65L3WblqH6QQh6v1/cDal7qhXyg9Md
rglat8PCMxCrFthNjy9I+hfBenUhBPR/Rz1HRYtjM/bABJ6dUAwIuAnHj0z1QUH3d5T/kTJpoTZA
B3BPf68RwyHp6fx/ms14RxF/8L2gYFly15SojBOqOfqyz4AFpglH7flEqMkVK4h75bQNwXA5Ry3A
AREvgqixeXB5kOIzu1/0Rm6CWhE6J4cpLhg+40J1IcnuyzlybPZjvGJD5EEUhEUWv9tnobtIScwO
tRbf+9BTuijrnvzyXJp+ewXrFlCYtxsp0a2KdonNUyqusSAiskKdiT/m6V2E0k0ZamphGGLvlblH
CuT6gO+d8dYKRSQ6zeWx4kmltqpDqZli7qPlA7qtUdYMHUCar2UAYKuw8+kkTJwAwYhJjLMF30th
57v819g+HOhHwvU/s9bfnAU8l/XHoTLW5/6UNvoslXk7BqAyBGsbOlQo5GoO/F9LjndtQvBzM23h
39Iny9nD2AkJ9vXOT3um01VmmVJ5lICN/gvEvaAaxjo1sRoz93otRmt/VqWYGc5Od2mKAx423gDs
ODp/N2WuOGH+k8puXvKhyriRS91Qxn5Pec6/xL+miIh43HD+K9dfF5VMaOdRAA8qYtf/TDeqp5qY
qbxFaWJR6LTteIiICtO3Ng94oUatonY4Kk/H2YHSqRDpTDzMSa5q1oVSADWxAXuGJyBDROrYAB2W
3soJXi5Sv6yPf+beORpjBgx5BCO7UlNCtPyYB1OW2s6dmSFZyPP/aomSu6Kp9h7McCR4iKev9LOB
nUZYDaGnPpjWz6RJkL9FF3XlzjK3POo/qYXiL8xRvE3J/Xhvu1pCZ7DlagKy6Rgy86QZsN0T+h0F
3jWQMxw2zaJks0D1d2hL6teaoel65jemkR3k5lsAekJhWh2wWTm97MCjbDFNw6wfZFaXaMb3mJQX
ad0GfCEgtg5yubUeINnZBRDvWdE/ubXOsXx93lLM1r+rQ92j26z/uRzQxv7mOwqHuzhWEXzTmcCL
GGEmlWog6NL70y8OszF2Eah06Fp89EGnWbYryS3WxUCqdwiv2NsU9BlmtEzbzJ5S4pIhqwMAaQmW
JnpthjIO133zsepmt6EjvCdn6RrHfDxtYP6mCKwIzpnCN+8WEsyXy2fU9lcEfCg8HvyZuQ9hC1hi
L7A0eJTHhkjurnfuuJA6cjqmFQI0YB0JEf2dsVpyOh40SATKoA/NQaeTUsC//xNQTzuV/qtUrRy6
IrUHFXFlzwRBkwpdS4PyUkgw8MyoCX2xM4kzsSnlb+2lhv9ZDaS4FPsBM6uYTiZhYYcqIbwSyjs2
0r8sNUa+AvnOd8hz0hn9TI8dCgaBTPaPwc9e2yY3OMDI9cwZXe/ihH24riGg2cTqEk9Ojs40cgFU
SiZEpL/WSNd/2Ewhgh4adLhL1MmA5BaWtptghqdELpFzc5soxk+LoiirMdNiLaTAcCo6eMIbZgZ8
Tuogho9rL3wDuv+nNUBEI/cjsJHC6WOWGcGXs6a9OCN8IOYklRcRCLqt+SNMJqgR65U//OG/ZgVg
Wtwb3mm20WV00r1OijTp5KeCwWuockdpuXmdwJgGhgfsJK/4/LnlDe5pzEz1JBkZa1ErdPSTRYoQ
kWtrISsefKQ/j3PA/ds1EBr7ZIL0qEh6XsYgEPD7/eVEufH355Jkrj6Po33WHd99pLJp1Xf9MTi8
6VAQLNWKPQZG0hVysWmJepxe2v6wxROe9H/SDTtxr16uWFwMyDnsrzNv5el+cYN5dzOADB88pFGT
PqBC3R8IEfMN3OA7Qv+5o9Ye/dBtFv0j/RI6lnkwxyYPuGqajUfEOPYgIrQKe1mjijZywxX5lx0X
//KN7+lqHlzwjWm/h1d6A/XaDzmH6rNO6eImCQYWDiiZOtbDuD1RY4plqrb1M6AueLnOVVi0myQ8
RT8+Uk5rSTPHw19vWaH4ZDNut4ckLi3sz5jQoPIGRl/KYHEaL3pSuaknD2+xTfFHPifzjVFLxILK
185HemXrkbIwxlRgqlCbHc9Fx+6amexT3KouJcMr7zsD/3bS4TsuNcOjC9bP5A8bT90A29TV3E6T
783k3ppk+sRDFzHhqJxRo+ekQCxctQ/t/VbksMyBuNDksLCicwHa7fml1swKTo+WH2SzRzzZoCo5
8J3KFK+7ntQMaIAu2VofEOBBct9usZdp2Dou7mb0vPktAynaum/ATEbAG+mmPWyNQo4XQKs13eA7
EdcKlLb3OtzfdqOH4CAdEMVNmxHhpyQXCX/Z9faEEU06zqkLyqVkLhZZ0cSjB/pcrpDMJ8hdXZX/
eKqVvEMrnNk3QzVTJkaiq8eiaec1IiFdRhKdTPzPogq7+dprmiItpJIEfxqUrFs7RCcYplDXXmO0
Kg6XuujS1mhvnIzQPbPwzwqdNQEnMciIDjQCwekKAdrK4+o3IzyU5f/DjbpCsCtCkMMFtDcKH2Up
kgHIw6ISfgcGQ3wH7nbeG8IyFSu2esGXnB24JFCCU1LT+pihKvADt2Ahic79x0fB5wm2IFcR6Spu
ugtzr/Np5iUuaCwwm943812UdKvNxeD/yYba6hbamSr3oRzSlwhtTOptCoeI5C9gO7rD4HxlFHSv
ciXowlqFi0f0eMskAj+f+9VTF4zzh5nUVlGbio1ZrReFt0p8EJSmf/s0tyNduE9LODoL4AwBgnvZ
wkvwvz2gd1Ow02oO/AtGOxzAyg4Ln8mDIHsE2U27opP3kyfufD9PkCPzlrXXLPKr+A+Y7oq/rgZU
Tnj0glWGNArdd2cIuQidDuInNhDRINCqXP2k161kIyVwGzK0/hYJ6CtOKqr9d7AsDfZ5MsyVxtkp
9AV8NgEyIvzJckVDbaK28YhSr/OJXdZdheBkl793DSGjCqPnSCvl98y09EAm/rv4EKHujZzwYR0/
m0hmVQciSpnoUz8Dh7vOqrCegr+nA2zCS0zknT2wWNUVsXqbZPMQdv8C163ZHl833QfYKObFalzY
rHSZ2cAZyNoWPgpMUQLmT5sgkuccDvI/qg6R4Jc30HWYEnJZBRwQNRyaYUakspmn8P7RyQkv37ec
Lh8CoGkBEojyiWMpSsAVeThb2zZs5rkymMIKBx3/YJELovE6NLrwpp113hF0fmOea5dR+xZRLdSA
pliCc9gIbyE2QrUxunDqPO1Dr4zMrnvQRe7iJ/LIxYtsH0xZzOObEQbI0r89MrLk5xmzk7fRZxQm
m8zaopDm51EwxExSy5Sv0afsj+OeCJvq3j/0ckqyfdkr9+PRsvO9EiCsqse2+pjJbz+4+occHuVP
6/2ArcyCsQBgq6nNThx4S2WIDpriQiqlLh7mxOzTYWrxod4s4oIBgC3c0p57gehaUB1Zm9VKlJns
35Ymd87U4TQssX1b6GBfXOzIoxGfzLQVOCWB/2gG/2bT8ahXctf6yhp+MMdIrZQ2F2Em1tECPvZ9
bK+LsRDRTs8r5KpHoOL+uPoLYuxFWXJZdKNwgSjc38fNetHAQenJWGcNtjDRiTUzi7fiDo9AEf3y
npDj1QxZmlIPpuACMUJhZjTL81UwbYkFAkcU9B+76qBAvvO/xgVfsLfnCSU3vG38Av7ApOli0qp0
n+QNBaqLOMLU12Wwe3fmzGcE75G1Hl+jqQ7a0fTKO7Ii6l/jzmdFqg7aeIR93eA3H6x+QZ4+NKDT
v7Uxg3eqMR/wwtFmHcunGDswA4bc8uLes2QC8zdmr69nu/dZZT5mxW7u/KVMA2pofqw+H10psBXi
0XVjp8h04vOcPreX8tvCLFmFGGsX/uA9s58t8tYeW6XAhhDWTogJbPASc6xVOsp/yk9VzFei9eBp
Af9ZI+ysFNHp/BKkAgXCK5fnefSIe+WHBiLu7XuaMizwxopUktDcAK4otZK+iRXHuTXEE0Lfz36l
3vZgLMcSVQWbsQL1ebBwAwsVr6uryJmVXJW518ihq1Fyk/MS6TJep2tlPIew9/lruXFqJr0oBS+T
MkY5CfYXEdEKDLvtk0zrCTgGMHouE6darxTkFMp9brC9ERUW84tlCmwhZIPHikicf+f4fAWnPaD6
d7yrQk0SwXwsWi5u0ya6+OpPRAP8P8PAP8ISUJ3VF7TJK1Zbv/9l//9RxHfOr+xsCjwPLCnl8yUA
i12QtPE+XPa/tw2tDXp+y6W3hMv2/lLJNizFAmbOwb8SCKfaB11eklsiNhEiyrl88JkYpkCEqGxu
oIPykYMYrhLdoM9wYoB1YCUl2MREIJPwomhoGqQsH6x/Yr8UQOs3Am8gmdXSVyD3SPNAK9kmZh1B
TJjs2jbnubOR0ylrLsNlYdGBLYkyR/DmVcPAR7ZOHYWSmUDqANZHKiCnaWJeqHr6hgf0W5mMVEe6
Tmc3NZBabtD7QUmVsqjLWpCal0ypZiQB18mg5Er3Nbg7Rz9t5kHo3uy9dE4f6YV7OaRKE5fs+HZj
QTyUCcanP1CI8GtBe5hz1A5FE2vOSC6ycl+DgwpYBdinEWlRVazqfCpB/RCRdbw+I5fzrlKWdxUF
qg4YmW3MD1G940BfzwjYZo24IHvgn3hZxxDAsC8dM9c5oAdUdA+mRoRXQ0bj9h+HwdstADPoO+rO
DeYHn7bitGWXYCpD5ETA9WYmBm6VqbWZCl6C1JckvJMULtnAGqrcELU43JugX4UxeXOpo9SG9AOJ
vAht+p9V7wcq2+kZwAafyi1QCfNGAAie2ioooZpEpScIGMuEZKGOFp5X1a+eGDhva+i2cM65E1ty
I8ihna5lDCXxhy2THeegHneQQ2ebma6xOgPlIs8xRCqFfrYyfCkoo7RG6MpUw1bPsUEWT/vcFuns
j6G6U5uD5T6Z3gze/LQtg3Vxs+VIdhm4lsGVeFMTloJ4q3+kK9xar+4OxZczyNK2L0N95Q0rhROx
Mm7NJGrfJt2BVu1CNvFZBQDWKsjvJ5CyWnsqIaW8S0fBZ7wYGwIItNFy8yKXtOYa2NBYw9LdZSou
NID3FZQ1YVt0ra7ou2AYwC3lHSmZAXKfXE4u57ckf0GQN7rkzndSWGwfGJ82VAtNddU8w3DqfySM
xboE5hN4MvyNJn3lqxFmEQafU5JLUuOrpwuIuPRkq7V8iIq28wtda/0mEuHxyQDO4OWgjuYqLixP
uHI4ZEfwhuzcS/8HBDszv8tZDhLAwrovs0sAhLqp5WeIDAIC39nxyVp8hwYp12H2YI/pzXzoN7We
rciTV1RzuPIKAsPGGyPYsFhy2TkmJJHdpg2lJ1m17Vs1zZoWkezhdItWsU9qe0/1sYOC+hAWoSA+
y55CuAK0+HQoY5ZWImhW7q6JgsdHXI6U9x5sYnMSYh7KFKvvWoBm7ucglbCidWzh43W0NZVrF6tf
ZWK8KYhbQ34Xsa31QRTbpNlV1rJqO27HSGk2PzGoXUxBqgwKcWPz9H/rvmTLc9uAtD8NbkqnFMRA
DBpEZrGC3EblNgHAXSspjwz5M0Wr+uvU1+wsraaEiORoW8n4RxhYsJrrRHeu6c0sluaLvFvzyD1W
2nuPHxc0mXfvRe5hx49Ivo62aHKXoMnCeUhMLrNpx4FN7e1kZpXv5GFzTV4PflHkDHyXUT7sUe5q
KDNFkK0QMGCCMxfdQuKcp80p+Vd5Da6TPZ0VE6IpKRyihoDLGeac1e5e1g67jkb4LeRyBxmbZ0J8
V4q027ifARszIC7Z9kJfLHpeoDoGVXTUeeMbh+B2PEDbRR9zlsTtpa/qLEBvfxJj5h3y42fuEa1A
Pi5JWAtBNcnXxbvxEo/WZ9ZITzuK0UHrodMRlZuNuGsUqdZPeN+6p/bIk0bzA0BDJ1/az4/uUXVV
bsg7Iptxh0Cog2EB22BGtfUuOdH6GYq1RAFlaJHQ9JaKra0ypw6sTwB5GTUXiBy3N/sUfNuYZ0D2
xHsGIHRdv8x2gCiyP4b36KNpb2a3CXGlnuR0XQ2j6AIu/3y6lcb/EvZT6HwFvIB92EtfKFgYN/Hg
L21ErfDt4BLL31mzYJZSNjXpfB7mJuE54PopbzH/5hTgMTd0SBrodWGXkKbq2EpkyPmG2Q6SWzMs
6m9kRtGkVEdBpx4oZlVUlrZ4/Auob8qd+qoZZmSNkNAibB1R8aUkQtzSNZPIm7sXABnD8ovQdD4+
Nhf5S2UeQW6uSgij1DZgoIvAxEwavADNmV3COYQomEixQY7Lkz4Cyy/jzg8OY6L+GovNvyG9vewD
vkx0y36jxbTBHn2zdUQ/7o7Nr/vSGeDZHjTsrNltcU6uJCn+GPlA3AWVqD5M99v3m4+b18PMSMt5
aI2Ms8lerUWf0FXzBxx+KGcQW+94l7OQv6NoukidRKR/MH03uoJgWkpXkeTc2FwAFptD0WgMK1fa
d15rqmG21kSvxQAPk7q60SSX9jv48DQpwnyAajePfICH2SqgZ9GBiSyfyD8IxBbbWNt2g9CZ68ho
x5ZNLL0hzRU26IL4XyMudupHzqGWBna/Kln2L5JXAWCZoPd3FJolKV4e9tlIoc+jcTO4Qd+Mam8y
cAa0Cp1fUu3cQfDWNgyC3FRdiC1XNgHEBj1WjT/ydaSeLkxzlvr4XdaUo+F0BKluSJ/D13mqmLb1
uVjQOzDmdS1U69e8mjdxxz4TWMGF3RJJ63gGUi4CIs+Wm/oP4EAPzks4imVQFVDHZU8nWYRXi9hH
VdLn91F2qAeVXkhVwpMyXjyaEcS6Wb4qCuQZcTUII6+7OmBe9co4VVQ61dId3M/SCjz8fArOeWXT
Cz9y2ZjfHAND/lipnInhFGpwW2o3uxtObzh4TnV3AmSCyVIOYPk6fe7MJPKk+Ft6FkrQq1fe9aHW
nL7A0rwp3ug5iOubFpqqMD7peLDpa11wDaFX8mU26u1ThFt0G6hSFm3nRddMnCx/gIrNsP8Y9XZh
9F909AmULANeBI5GvvvlzW26dYeEFDXD5qwcD5BFxiAe/cCEuJBgM/2+Stydyb9zOJJL2oxWERI4
JFJf2PPzL81L5MBrO0VCU0AvrMmovd0GMs/5PsMhr+4nTbKqiIqQQHbY0KTTZfIe2tDeYEpxOa0a
MJ3dFueNYqEtH1zRovhorwStbKIBVdO3kIKW/1gpFfkt92hF0VxP14ZwLIQtIoWRZGm++V7vGAVT
SK6XiqpI0owUZfALQvLSXBwc/Cw4lPR46PUT3Gc+iL0ensD+vsQ69E2eDACtpG04XTY0mTgnpGAZ
xMpgsnZUETxRFJ/jGoMZaFsWm0qN95tstL77nI3A2dGDy2ioziJmxNFpU+L03bbHBPpragKDE/HD
fBgrH87DNg5sQSqYfYeAe9G4Xnpttcqg9P3OSf6iDf8vDxP0s47izLMcFVezhBjYBA2adlzxxgOb
/eaMfWF3xDjSIK+4ubgKZRfI+BYL3KkWhO5bbaFrcVXXXFVTlm1Qko1zCGf5z/zrDCq0huR8w/If
J7xHaCnVJy5gmyVgX2v1B7gUTgIs8sNuMSKhBmCkuipb5pFkcyUbZCW1Hisi5MyI+Pm5nDISaRcx
/Rj8u57TianioybIY/TFBz6pENiDEPrD5gHCfDCeuJfQ+MIC3N6adQOIggNju+/7UQRAC2gg2ynb
AKE4siLayFFeCsvcE7DgtnC2weou1h5fnNtI5bYnFujzbMa3x7NTNiKIVSKg4ZyoKcCOiCuKKSM9
C68fe3aGwcGPHbN1vocGGhsJR4/F4uypDuyJbN29itEuPzyCb9lZgKwBadz22mzVt3xxmV5Z3znd
vrPovS01ecx3ObJo/YEIa2i85rjs7CxdM8LK8+JCdOqRLC+yHhHsaVkZcX1U7pKxJpiIk+Kv8EVa
kqy1+rxG6TOeWQwKy8+CpDEZwwylUEXvptSQhH3WvQA9BCIPlUAtUF/6z5EffcDFRVQQkDDPJk5T
97HBVkEVCW4ExC/9V1W53QV0QGFuwSaXwHQAdVXZqtqQeH4uJEShEISUcwPxizYdvItKQR6x6j8j
NbVMBZqaaiKCCHtByWOSmG6xwFPnarlJ4isSmyLUHss3Uc+VwKaP7nnFcibakID9oLioExNkXDRk
/L+OCGI85h8r3WTBFBf3bQzRyWxcwELAcAAtFURHihPgKaN1fwZ87705RqdLjtfo+7Qg00dS6qoe
NGZX4H4wZxoGAyeLZ3AJZLoDng9GOA8k4LVfNUCIYUkNA9BqCFOCHJCVmkRrCIrPGTN2XLimp5pk
O4OzuM0Dv3IUb+jqzjW6GjadW9mvNSQ8esYo9tHCaVHO8WsfKbNIHFl3jv5kA40uRwwvCIiNa0D6
YOk7VmxTPsHXniiGECo2KXs1TttaD3KJSd+Ta3b9TP4jh6gQS7eJ8jrCzQtLvXY3Xp4Pf9K+I4IC
3tr3Gv+pqng+c+39Sg/5Wwb6HiqNdGeq0tb2C2y5/n24PrHJXtGQxYp/qBLgb60nJcaS5ffnklW6
6SEFbBgeLJOrNDRt5+w1XJ/NrSoctbOLdshbqDDUthP//7E9eeJ3w2nYD6aLsVzUixOkYsejyeDi
NxB0aJlAUdkJO2EwXUygA8jJDA9SS96UdKTHtnPVde4wP2kCGrp1XohEiMW2B9Ezqbgw/Ud/VnM8
j1RbdAzjyx8b5VHlX8z+2ZiuIVvBqnEiq+/7BItkibtpOo4cnvSuMbvtvGIo+Tl/6/8X8NRECWlM
3/HkwfPsC+KH548Azm8JSdi9ZaJzcc7B+3YV6/Zo+wMk/mfx6YfIbZ8AF7ZFg7lHGcBVx9Icnny4
MAr5fjGYrGIki7LQZxezgweivUlklY2p4tRbUz0QlDlGRweiJbP8GEwl4w69ABZoYldzpLhNnZdG
1pJQwXbquqq5LJ91+wlFmAjXMEqeudsDyz3fjKW7EJjDhSRag83wDYF6KUR2pJp8LzCFxss/SFTc
sbjfxOyR2SAdzXSdRr53lF6MzyzrEzXaVADm3eiMjPyvtDG2Z2lrDj0TpmyLkzCwWwg1saggk4wh
VdhQ3m9/OsC5JQvE+KeZRzNsCq89aMiw0VkJ94eRDl/ShyyQ/lAi9wfdzvkYZKBTvjfYCJgw3bFz
ao1rOF5IpMlYZGxQtXRECBrDklXFsUi6Mnb4zKOEXeGq13Nc2KcdxInoSGTe6yaRCmu5P5rDXtVr
jIHDXSv2/BTxYM11OkyZvnJ1PQGM/yAH7r7RjpyXnLxTNVUa+plJ6EWSGi963Po7fYnoDMIjLtFw
pYaXnroCMPsCmmVQsWuYDxxNqDhVOT012SsrPoiQUdgiGUVz8f0PX+r4ftobHJ4prIF8jq6iMVZO
zOBtSe09ZyTCukSDXoQwbmcENlxtCYPC5tgAWG39R8C26DysWXWCtBKBEqYTf0qveVcpdwR10KRa
F8c9b3JzT2Ccf9pa6TO3NGGpJRhHJxHzZEQpbJ3ZfWb14TyuuV3sKoRkzrOcXiacNgSUprQTxHoa
BBvwIAyTjWIh1kcjdxcDmwKr82ZWTd2amrNUeytvaYDOJZHIG6N8Hzha+z/85BmSSlE0eG83fh4m
NIgz1kthQXfnIYDBhBQPu0iy2b9zv+m6Ya0JNx5zn/LcjehJ9LtWf1sgUhTYFzWLLWZFD/Uf/8VU
gol8hh1kR9ozpst9HbCely22arF1TBess9nRvPC+bFJNtneVWVzRwJ0tW5dqsJFLMpfqszXNNJa1
Hid7Ap2rooyjnKNikR4wqZeRN5q3NfU+IvItQzf6/xqZs8B/WBB97nrmo0qR9ylH1UNROXQ2Bu7l
iXKFc4nhXgeFHGKk+fX7xH5DHtd5Vo4BI/1gilhefadrYcGh18Ew4GaqLok6ccrE8xa8KtqRpkJm
rhErcE0mL4fbfgiCyx7+cvQZHkqqJMi3Ti2Kt5UcBaxwyxknSEDiNsr8YQVRlomI3ijQU7K+muZh
q7x926XALfrExzugWnMtVXwjoaMBFT/frY3XIaigg7pWi+dWBAVl9dC4bAsXT7ZyEhiCh/ev+Zrm
W48tRld4zQczA4E6urgVbNBvJlfRTMv0VKsnuIUSa+LvYe4ei/fKIdZOQTghc8GFCbB9zPNb0goi
ZRe+POrmAHu1k4s+g2MCgh/FzYdovWUpe8+Tkb6Vvoz/SevFY5qCCbG7M5h/rKlBirdCQAQsI+Cf
Jp6sbNMP3X5kUrEnVEtuDC1tukM7wTkfYea+WplL2ZuH6zNuhL7GlTPeJsCs3PRCFFqc8el6oQg5
hA7gnvx7YiU7q8T9dUZ3R9i2gN0QAUfNe8JQqm0k+9niBJTORPPu4Zf++4gxVSRkW5yRRJM+K/PP
01eSeShJVdXl7StXOVcyNs7wr0lMFqy5DKRSR4vl3U5GUl2OYDX7J5pMjqoNvrBZ1Ah2mgWaLnuv
0PuAQ52Ygpaz9o1tV03xLZSk5bktgMXtEr3HUhH23GRJoJSEL9V/1J0grs7mI0WrAkzWyzd/9Q1L
QDG7e0arRmK82+jInI/O+JI/EHoFLBH6aqVX2DO7u2kk+APhJLy7qCLItV+fhoN2g6QIe+wwxlgi
CiYJ1XcBmGMPh5K2i4M1cYC3eR9woZPtf7p9rIepmLgCKgErtNQZd8ifSrfNl/4iphFCcWpnrwkU
z6oTai6uZyikMhw6gdTIF/0qR3nik/taxX90Bk1nwlr4CaQyyFD/h53GNwOqIJROMwhbzCXePYZM
Ihs94fAMRLSalOka/C0L/9W8lCZJxBCAJxBgC7/ledJ6fP5tXDI3/CkS3WBlgJZekHnukzgBNhyH
7G6NxSvpfdSAqZcC4AuzNoKD9qL5IavvjAtRj1gEGNhmjd7lRLiUfRY6p6EWwHeZkrESTBUyM/kd
0hay0ypcqjx3LXR0Dvwp/rHSShqSmxeFa1hwA9q9TEG2iSfDOxuQJNYsb3Ui5a9q3WZNk0BdHE7h
AIzimWhzgOkSi3sOne8niyLFwcYGoe20jmyY72o5mkZemERlP/JPcKfOTNbPXrWIAeGmV+lZ40zR
sv54sLLArhDU/TQ4hvmFpt4afiDITcOZBGfwPdpdndGtWfIeVT4TBH1n8S6bWM3hH52a9oa7wkBK
+SMVLMINi5Yx6vCugIE0CUu3Q4GHmnGHL035NZ5MD8vVBnvBw5MeTDKXriDZVfx8O6zvMnXhcuNu
VpDf+2KCrCMfp92wkazItLDsI0h6JHwNKE44dgm0vPRJAJD58XaEVDIbgyEenHYxOrxVP3TMAiBi
yebwMRj2O235QJVjc7/v/y3HZJGlB514O2W3bUPDkBSSlxbP0q9AblFqybVSUEPZH4HIZB2IZR1r
0EtiuozhTceKMXoWHPJIUL4ADCKjN7kcbZ1tvbxrDIgjwSyt6PGw63XipT8spvn8w/d8GCNEXUdL
BnmG8Qpu6PuPzKBBfjaAzDSwNZK2pv6/oqehIve1JJ1hblAFFRy8hrD5uFoMKfuXKoBj1zptgl+A
R3EiqTuRAnSP5lPkeBJ+IwMVIAAt2JFgo+B8gp0NTcEhMvxL2cHlixatcc4cY6WI66Zc4VT08vvV
NmG0bSLQaMFUb64gGvGdiRWzOvkt13vz9Ch6y7OUm1yednuh4dT2c99QQCRvVVO2MzWq3R7DB29u
yzE3b/yQPMhzcCB6Tp7bPyl48c/1E2u4VnGp471osoaP7iPDzZ7odl/WAvaAgVmab83vpc2T3bGI
+O+J90tyAB1JB0AiEZL0wHeIDckg5KHrnl2p1TlCMvn6pgLOc29sYQS3KTIJOd2a/9HtbwbNrmOL
YPVEH8wz9zMXOD5yNaWFxISQLNWrwOtUmww+zfH4dxICzCv5ykgE+PcsbdFA7RS6NVR6EbhYwBpb
ORRvIHNDgzt/8anSVX7lj69R3SzXjYJvsoYGPGy7+oNGLYHl2Jqbx347H1GPKKoxm2wbEdZ2chfB
udgDxY7sZ4N6T3+QZ805xtLsir6DDKvPLkjp+orJYCYgO6i47nXk6MC424uhdNjAgDIDiT8qXGMM
0uxgsgzKoy6QiOjyORBo5NuxVWiF7dnZ6sh9K+DAou5JcuDzxgVIqT4gCq+LJaTNq6giWvq1Wd8V
0V5E9xObBByR6o3kmIpo7iLS4o7e/DitburQ2nf+eftEHh9DwVD4EKNcGPt9G7KJ3CyvdAG+EQ/W
L/Orej2Cd0scSWvV0hn4Fdzeeew+kgnyfpakmBGBMs6Zjo0Qcfj1V47tFAdiUHCRlDLUoJT6u7+/
9+a5tHHYX++TxkKatSadrYIO7F7epwLkWvHTVHAsLQ8AMixotLuDX5pHsQcxrTY6qZjzAcuLzk3k
+qxBIv0GXjBBZayGXdckIjRCmIm7CnIb2ikiZTeYlmmGT/rByuTUj6c9JKy1iGG8aDG/u3IuwzCX
DzXrH26yTBzrsoeeqTb4b8DrHDeqg7PYyIWvFpG/pFSw7zyk+A4hIkfeuGT/zBN1bZpaudV8AnmG
nhCqGTW9QN779q5BSPT9eTmJIw2AvFjgjpAxt+OOy/3j8RVfjbbn60ANgFTEyAwTVkHWCDX+8mnA
hMwH1Nd921QNKPpq6vahzeo0ghvtvYQcYJbMGGc95UaT53ts0PPtK9BPqgE/fWUYHOHi1EButMgl
DjgsTMmLX6n1xVmc+aa1jSO5swln5H+Qm3TfNPm4wwNlPr7ZmTX+X+vXDKfhZJBqxyUDuji2kRG0
6OL4O8G4Hc6xz9lxYcM7+dp67K6rv6SpeuJwa1MSZ16cAXLH8pSZfDHqmYMMDDs1QevCVOYq0zDz
EwlrHz1j3Nz7fsV6fNTuh9s2hJZ8B2zkdUnTpMWbXrZw54ZSIdHTNM/cdZf8TS0fTXlLosNmekIv
p0fQNsfH5R2/aHWZUfZWwFynCfLs1bW+5VFJ/eLDFm9yidBXK6/PJUSc4IO0wOWSON9mBn8uYJyv
SwMBvI3wo4wcoh/SDk+GycTsONbSpmy9h0jiEeBT1VwEyAKTuKnk0Zg21eivoDaiXqpoU2ANxC6B
XjiNnSN1K3BXtgq+Lvuwdq933PranqLfQa4DSx3KdMdpuS65O7WkzRgZuxsw3rUriwbhuuhesse5
2L+CE3SWznSlBNjhsoddgdOXrts4Cp8uxqcqNkD9VSmRbCwZQRKGjXX5s8GE2XK2vG3kjzl4FPe0
VZnesuTY/fr+yY3kbhIYLTfBkaBT425SxVl+ONu9Kll7zZkHNPtOfQuGxan1bYDXkzDsJIw0MM6s
bPYMwlhkiqgRpNc+DLIORcuhrrLjCh/C/r+Rsprbq4Yj5F3cpDsNrvLjIfplpvH4/e+XOw83kh5y
dL9kZ6IL1oMT2VOyhgxVXLXsLYQk34pYknZtgZolvyvDiWnBpC6hzhUqN0/eEQXNlQvR47//q19L
ya+hUgN0bbiV3jA3wuiDgnMykPPGT4pmrbJ3PmlfbEsR0xA7mQB4mscbz3m+hk/w/nwu0wYGzkbV
ypgMdZA3AVpUnjpZ9LPkExV5gWpEthnK8JBRbk8j6LqRawbZn6CbI1HJ4tqqrkKVuY76oqndima8
uauYFlz5N5sR+I9/B7QcFppTq+38KBttSCtWOQYm0w8fvwOVf2RyCr4pOXG/DeTVDPcpLpq/viE9
UNtJwKrHM341jZ38FE7vlHr9gfGxPdZLNxijLTBCd2lMGOFpcBTgZg088Od29oGTaVnz5uLLc86m
fuoqxyETteDlzZt++g7hGGPPGOT/inSdS5o1nKGjrO6OJxyH4Et024q2+PvksWOlFLmadMnhmWxY
lz8xzTjpcEiesXLXNuP510xIXn+oWnwkhlNyk4szB2ohswylmE60VnMQ1AbOMhn7U/ewNBKQkssd
xWan7Pnk4Z7ysXXpsl2Z9LLkqOI5KXcMyrh5yS7Fh2RPAQfCMhRpHNX6xvr1cG9KgJg5af4TPNfk
Fx1Majbhr0cXD/CSaQrx/x/Rf7hyZkLUSh+e9j3VMEcH7nIG0wzL5cQEFXVcP+CS43GWvDyKXNWX
p3DJi6ILFHkOHN9LmDUd7VM76hSeBZvIryf2WRagBMgwSPewI2uAzMTlgUIF3VeUAnOiI15JH5i/
XJzamKGdIRLyts5z4PYhy+QQ8m/Iv9DbeOWD+2F/TftlLojG5CQU44im548zhMwsM/A9dgY6xtnH
2XBh9xGY8u7lewhTCx4MHpX7WzlHudxYRON83BRYj9Ld5+KlbbSZuoURloRrm2FTCUSW+yKYNZzc
JVi9VLy1X/lHGje3GhaanmKZnuPMbNhrLpu54nPJiufs5edqVkS+vL5iQxU1tl1Et/mD8BudEbMi
tgw1va52ubB9x0NFDPp0ZBbAG1f8jM9Ve3/DFgTpGWDSCPiQKQwq8J9pbZwi3BaXQEfShkcigV9K
5v8ockjV9QbjJuNDEN65zG9ivkkTNVs2FVed62DHJiZblfg/HImVszdIUlDGc+sZVHz4fTt5Usjm
dibQOM9ZvmSOvbJjEgcNEPocDPqLPibC5CacTwyGqW8d2oQ7/iI5JOSuFnFPOkC5Bkcb6sc9PuHS
0IvReTYekA3ZaZXkLV5wujHwJCUohKI47WfhkqvjSz0x8r8JqEP6Md1DC2ofGmkchA65gNZ24ElK
AWEGfi9ZV9DknDdHqZBczRlaAOniFn9eqaD1Ctw++jnk96CZd6zamHprITtsYm9QUmK7CFQykdfC
B5DqPQ2iBhGH8jDqiPS7zNESDkWSQ7i7vLHl85gocS8VqrpUaDWtSQVqbI1jssENy9pdEF0Otlrp
lMZLpxlFUwsuYWb1JJC0nmAMQA39kx/lSNzUgRj5CV3ZjsrEWxblOdSjyUeHJXweViF0HZL5HeTO
4SkI3tkJFtkTfxk1dz36jUdNJwi1L17HbQZfirQTfAjp782eWTlD5hG5sDmHSfnKB43Fvz7U/YQy
F9TmorA9SYR284duvVNdR2lNaMIQT1rFoerH/yAsViSQAynn282+mAEcKPOLuCti0sBv+Y3VOl07
IMl1+lXpzl3CyNYo7P0tvIya+m7Mek6HVjqlUNw4HZhKEnzB7SRNHHVS3e1xEbkXivyU8yltZdn7
22YOVITPgZhZzncTFbCGNP4jM3LQr+ZSbk750+IWmbQVmdBhSL29PIpwLdnsHp0vuXnA/CeJ/KG1
0r85R7yoDUY9dtFdJg67wvzBnmBG3d1wnbJOkPEOGiDYY/mUEmJM8lEfA7RUUrYUoQbCESLuicUe
idQtT7FTbt9kqk63evkxLQrih7EjTnBp6Lau+PjihzS08ZfuD0h/iRZ2MKctu0W4cr56hLYfEUho
YUrhz/935jeV4aUlsBJRAalxWm/yvdd/gSAIwfQ65+FhauqFUZ4dyiczQdFe8WPpIglsNggMzxeS
bXfkrJjbTfdzWXl2Dl9E1GiiA6LadUcIPzqCL45BINDnHaVavYgVV5tsUCQhzuV/YLbrV7pwgUvb
6v7GNOiwlUWpfdUQqjG2G75aAbNS9RMPreKxfxcgf3aRadxemKN8/AYXkGmO/mgvASG7u4YEX6bx
Chz61B2qoN9vxvoeZplR98lVSz9pQAkO11n3e9UqiRLiK7g9ioieL5e50q5ntJK8ieM0JeEZmjQO
U8edwKBMltBik+UL+xm8U3c3nYTgzzKW5puenvFNLNXOsqIWu1dyimP/mz2KOEpR5x5FbDxYRJ41
iDHODvyVjPfFSSKGZAjOJp12DJMkngdUkTBbsYqCpi1mfV9IWeKNMHQ6DOZCwYM5zmPQbrFvyxsr
aN6/J8xVUM199/8Oq2R8Nm3eEXusRKguAsOEIY/rdC7d8cCN97hxpsIyhswS8p9qaQZHzEVUCcUK
dHKa2YNS831m5s53tSoerHfvjBWnW27pnAaMjNhvz6/LfP2oMJT1wAM1WubIvNKo6QTAXQtAq9ns
ra7DCKIgsVoadDApN/xsJdodYA338zYJEasZ7HYBDipk7qcomAN2WTHHb6iiWnEMspJtGODNPWHQ
r1BpU0ORuu71em47sIDF1nj6VcnkRsDJ+YXF+XD3nMK3blBx9hlXW4TmQayK8APf3ht3xycZKPSq
kuufZ4CkhAKOUKlydl/GJhl7uBrTKs22aNGwf9RxZaxsJXnJTKA0e/IHNYfZRMWkO06sEIol8dtl
LOqdgThy6qmaX20FWnPJY5BXsi6/oAwbtgJeEohz99lbxxilvEcK08pkbUv578ubNV7CAnneDoTa
a7k3xj5jt2LI1px/nJ51cfPPqzkz6FtFrH3CxcB4dkzF5pVhsZy2vYmsNjPghlujJ6HMkWyJDWdX
DIYLKt4A9KrCRXkX9dXdmMjeqJL25xYTyAe1e5uJvrhhItXbuUhcH5DI0Tl+q6B9NZZZuGRudMTw
urcfp25xDYPqeITBsUlGmYIrSsS3MhjuxMBOaLr5A4LZbT0GeL7DVMPEhADc0eQYbp+2LtvC6sKN
uQC/13V4BwcEys58GWlXBlTDhFEfTxOcFuSmpMhyZ0MOh1iOhEyNOXwxE1JoWHds1PjWE3Jyz9iJ
7/lmRfYELOBMD46+g1y65FT8s3D+OrxNSZU7FBD1N7n1dELiBtMR50GK03CIptZbQSeqAJ7dGyU4
HdANzGQlUdsEoKZSdbUgvhmbbqtH7OsVK1P/Iz4XM9AzGbb22NgGMtPHx+rzKY1khBJeR5EYLPN2
rxxPGa6ifVTjS8z53hnegYd+bww+ZJu6feQSu3BjTOjt8OnhdkwSSy7RKZKnFlEBgHxRfnT8qvq9
EM+ahGcB3NoHMjCSeJ2RxPhEZ5Z/C6b36mkuGmtEKEAutHZgJ/k8TpWBuHk3KFJJg6dHarkxwa/f
D4YnrVSdOkyKWFIqUvHFFZMHLTgEXe8e0xIcewAyusKfRvE5u7mLL24HGh51KF5JHbsbVG3ynA3j
BLMKICDSJJBmIW23Q0OBH4+VcONFu+WMG4RABYBMih/xlpAyD2ecNlRu+S8CpF9FLgAbgefZ0ULo
fK0qIF318vgo45QPXfokXaeemIavV0HlQ+RMTcJyfR2pLYDX5Fti00qFXQnfBTm08zkUpNHLRk1v
/V4m+I1mdmBtDPC2YaO8oTyWB1w/XFr1Etg6cCR4GkN5MRFczb+cXAu7EKQkHoh/xxFSz02DvogM
n6Ym/opNNEa7zNRLfmKd0M/V4lFr/ovgaDZPHmMOBfIRj1gJThGXd7qG50f9JfhDddL391OnR7nn
QYIiCpjpnGLz37UZJrCajchzsxF2kLn1KxcEe4ocr/3VAWEZX2fCFvP8InnELWPohSjryNKJ2M4k
A0d04ECwX9WGrToH7/T6tqwWQfoZSZ+yVEwXRj7V9lcKN5WVdhqFD5AamHOXgWmebdpWmG3qvbSS
P9mpVat7ipAcfRbqKHKmWDrU8PUgiwjbCLtXt/c8ZcA0/PfKjaVYKYl5p8DzgH+NpFTRb+I/tpSZ
SWfGizrG76T05VzlRKCPGTRdiaKtVS3oGDqwR7hvPcFWmo3UNYYHXma9rc5ueeUpIMqD+FPEyYg2
sv6yAeEUDPpGR5GexsA5EelvcP8C4flgTnKjtMWxTLjPQX1jF/7lqkhxWYl2l0BfVwul8oCAclX7
9d1d+GbWGWAFud0sRpaBA14Yk7dyHoncNYjKd+NWcp2PdAsSkYT0lD/CkXuU31EfQgzKul8hJF6X
f+Y5Gw9Xpj+x8/C8Vmml5dWd8BRQGIZTY3tHZ0iXe5ULPziYgUEhH6v/chmeC3Og6ii2PXcv35Mj
+RR46x58ng3i4+VyzzztNn6Dc8EJBssErrl1JJhj39ezoKCycxMk80Xrbk47JX6IqPji8QhUkD6N
E6HCKgbsggo7YdvR4LxV/kCzASC8zyGFI7r1HmGpzsWy45TGBwpiNKMpQN3tZRE3S6tiqBBCQv8S
ndj65nGW/6BVwBRUuyaCO6pov3+3IbMZJMYKKhyEFPEu8n87nJw9imgzpv9rSk8LFoDCMxpI+9EP
VQyrjWnJXFgtt4nei3kpqTWtZc2WKNbJdJBKhdxtOrn1GkTCn27URBSg9myDp4BauAVvDCFfM/FK
CXtkK/wIenqoReJdfOknV6ZAXYkXcCqaZBkEHKNGSey+Cclq5grd6FBoEVLMMfhLe1Vu+y/YZZxj
0+qR4tnX0BAzcXKuFt3z0zGbZS6E7VdTHAF1CfC8wWXAUJj8HeJPhH4HAH2DiNt3N8pOebQM2hX6
3l7Mzs9pYGkc1l/pKJSjJo8EJjRr+tq2cXIIUgLuzb+TOZ5WLMh+sf95iKkH7zuCbE1/08d5jbUD
4T3Hu+me03fX6IAupk7HJL/IKPD4egHzjTsE7/UJsGP2SC4lsX8u8Vmgh/a4DRWkYZVwBUbuAKcT
s0q8BpZqYqzuIMZB5S6Xs6npKh+56ejiUwBpTaKg4jkC7XGlgOjQEuQ/kwy+xmYP33m3/6YAiplf
s7tkAH9UK/bBTYSu4I4xVOEmEcU761GAH0HJzXsa8vYThZgfJUKrJcsES0St7Rp9h5PeVRy2yKi8
DmbBan4fg1+Zs6irI+bbLf0EQV6ZGZIfaHsQg9b4WFybauIvdDrpKxQpaibYIOTUYmP4grI4RsJp
YKEiLoQiMRpwMqZ5UAJZPhrjJaxFt3RFYkHPLjI4LamrMUEwTo9RepQ9uHX11DOQojGvbt5PKIg2
nx+BkACDo6tFWQ3MYLy7l39wsHRDoCTzQGp8HkDe25XDefLbwjR6cI6ouITJFfVoWRsE2gOW2jaB
zaDJ0shB6DdDItKSfLtIoeCOZK7k8exjoeisu4fhi6rW53isIvnlTVAog/DWENNQEVEiw+PwZL3N
hz+lQ5yJcDrHeTFP7y+ydCbHgZV1Ox9bu7W8XrRAUvMvsYhL8Lj4F9JXbAAVTYw0oxInZpULrk8n
aiyM75LSKy1BoQphs0rlzIV2Qz3f0svyfu7C4TGENQ86HQdjCoMlsgLvD5t6IA4bUWVOCm31WMeR
C0RDasBF2S2syOWd3b57kXJ18qZndbmXjIbOlm1F2F+28NzfhibgsrTBRS8JLKIrgt7H+19XaQ4x
GadO2GB/C/eQu91uGt6nt6isa3/smlOUiOqxCBjNxZjc2eKQNZMfGct25HF1PxskjYvJti1RAlV9
1lSb4FYt7GT3aU/LqT+izl+rc6ic358CW67h3waj3oUu7JrJKgwAL5fDf5vv/bY6TRON/8y5ae44
hMJJAe/2WAMrP5yXAdZH+M1UQMvSAhrz2OQb9Cq7ELmrUeJQPreTpqP3ilvJOmvjImz1V6ZBAYv+
rSouLaX0rLt3Ico9FAkzCAsme+zTLOq0/FvFTO2gqNgNOISUsN99OhR5ffQBbdNHP+vEc44HUeWE
MrWgyn/Sqz3Hx/cdIRNGxKU+561Eh79clCTy1k/UGVmjXi6OiBn/YXQ9K29S39zsndctE52DlVN9
7A8s1CLgXdXSuWpjBjhBjvEK+OFfLdZf1/9u5Z5VH0C7X/YRqExBAXZG/fOoaS1d4+W9u/BJr5ky
avDwiWiP7OaQ7EBQBrdJlwQEiaLP6KJx1cKxkZo+Htzx6Ws6l65jcp+pbkxJ1SIsV+zB9U+x5beS
9OFtPjlTTArP58o/HhmMYSOJkpN+HXRRFrdWDpy3pQMX4Ex9CRr88MTEHv7V3yKNL4+iiRZnGUZY
VeysZNpNpdBRClKCMY/wXoYwAsi00FpZr4y4Aw6assQ7JmF7dyj/LaAK2dbZ2MQd3H6rG2ORI3Nv
a5WiBGdTL/Ym4TItYDwBoiQPfuRz/gcTIEHohtkKYmCijL9+w29fQyz561Ns7OA8xKHpzeJbigY4
/z3WWRSmVmewp7hP5ykOdRpkdU8OMZVkSMU0/escxJFYyqE/9az2P/7vR9XYS002e+U1o9DfrpKn
s8a4Zrm/t/QTlovHUmNtT6wQdsxQFC/+iav2912tu8qqqjAPz9jsWtK+Ywy6VNrx3Zdk9Fhz3ppd
24Pcd7LbdSQCP0CYfHNG1ND2Yhqf1/ByBTX8fg0itRgmtibj/Vw1IouOCZzaX15HzEmqMVHMCaCQ
WDAF9T9Pe87fWnzA4eK1MyLw//Lr/EQaQKHkn8UvAWkl3Lil/mqDxs0j+u9lZAm9tV4UoERx7+1S
VRuWMR5oNQK2J3uPy+S0a5ZunCfzm2cwopTL+ZfWA7CLmRerdMG+IoFS26I8nHQg/UZ6d7tVjkKB
xaq6OblbI6qko3O4M2MbkXL1nWW9WUrbeF7CV8f4lX68mO6bWzyFRXMHrOFokTycYjK+O3lt/2fd
BZruPVXPVUeks8MEOuwMXIWJfXI1fa5F1zFfdT8DU/UnklSEFVGoQILylbXyytDa3hedfLX5qmQo
jrUIHx4X/T8LgKAd0g3l4bBxR2ZMIleJ88phhAeAUB14oXXGlPcw7GW+TjFkB802JwnqGxRgyYgT
8mY3cU1vjsGuGBPYtY2QF5Syx3M3yYkbpC6dZkBicMuxfRMW87++bSsOcY/qF+YpiDLmpQDVHvL2
W493AUO0eM9xiWezA3APtqDHSzlnhww4jhifDdoA3bTucoraLE/yOqq19cE+dPjsdlAxn4Xxs1kX
eu5DsJDn3nzzbmG703rsC0PYsjX6JLlFiyOoCV/XVmMmyh1QVK3JQJb8ZPOlC4M8nAQZFIlCBuLY
ndRY3UaM+vopB3LZABXCxoUPafXzr0cEyR/tk7U4gS0NM3z8hT9DJFSau03ncDkMh+ciQSiv1Mly
87YGN6UhYQssMiVTY2Vtxzs1D8Z6ZcFR5uQM4gP+fUU0f03I9mJW/vB+j6p4Mio3ykN2lbRStFpz
HncTF2cxaSC3vBZ3aVZYrF/73GmZh1w60XhITm06qCm8eLlxuOYsvGlgLFqDZ9ubDwIjsO0TArNF
scwnckCbOBoyvkx6yQ9hnwM+213IIHbWsdre4jalUZt8iPJ0bAf0toGrf5rmcphdNj1rRRCI957m
EVYKF87m8PVlHK4ArFn13ue+nxVyy3VOqgk+pSyT0lyF65GDaf4jG5VKTsQ71N4WPCTdEUuk/1cL
Fv7jEa+Eqw2Q7E8zWahwVOUd3kXRTTFxiyOi7rnhl+p3kd8zaTsEiqJQ4aRS/GMs4iBlL9T1SFSZ
iKXJBWKsMfs2LY4uFf65O7DjdKkfA2nJD5EjtXov2kpAkZaU/wGvPRLjevsCt/XYmSUL4IanoD8E
2F6yuXioHn3H5SHiTMp4+BFGFQ7Pj2jmdPvaBfOjltyEaY+JovZkA+34aZpDqBAYB1EKkBPULCdv
0BGnt327cFJty0DawqxBvziLDiqTgcvOvl4Tu3jUiB+7jJ15I8nrra1wYxjDB61UfLhJT1ty2g03
yl2M2iRFKB78Sl0KQ+qGSF0gMhfsr/vi5tl0fbebkL0KtH9TpY2jd9kYjqWRYsIzHSVfdAg1trX6
JhRuxl+IlKj9G+jAmyjB3nA7FM4KyWEldctnl/NBhD1ku/G56ux9hGiuaApeimTr9UuhR6gZvxHd
14VMixfL0hQcK4rZs/Gm9Yixdl87wiM03iol/346a2dJ1rOt56NSiG20L8+fjLqepMFAw2a/e6yF
8c9VM5RN6YkW9NpaB3etZq6QgIiPZoZqTM0gVyG3S64e1HNRzD8AtK0RaFJWeK8jAnrCkOCXlV28
O9LkODeZeFTJh74RA7YhM5JYgptxi0fyvKs7hmDFulIMdx5jQwaPxVbsBA0VR2qZOvEeZwC79iBa
epHHEfnz4yBd4YkxMJHgPSLpn09GgaybduE1WhugAvS07AQy26G36HwudDCzuIN8mz1F9AltNWKj
S1a5PL3y9+vJOqu8ucmMiyXFmvLr7Y/a+tEXE2nAmUVs7YKD0dPTMtudRcTeN1wfZC0QgB5GFSOr
smd7nr9pnL4sbgiiXCGx+8i5sxpyZVe9bksmSj52S2+DHrP6rvX7NDlGsAcMgAis2MqkaNMSBrsd
cQ9wMLjLKR0nVJewbqeccWNyKUQrCQAwlDBs5/GM9lstLR6n6j5g/hQkj3HZJYgaDwEqWyxq8mmS
0xOAsiwJRZs2xXyzhKjmTxWPuGCR3dpktWvARgE+VHZ+Qu+eyQGCJo3LxBLB4lyJMo2+pfq5Xb7R
pWIQy+dlIinZIa6jYmsdjYWZFR7GdFOF8QCFSt9ARAZO+StYnn5aGIa9Mmus6TFXlu/tD00gu80R
/itLHDvp8Sm4BdJ+o9SnUDVU0Z5LFkLMIq0WzJ59X4dX7MYGexsXSTfsPbw5w6BIRG2AbvZA1VZ4
yPQgSEe/NcdW7DlubwDp/+VV1fK/8nZ3GLaJ6UYf6JvD274z9hZJtRb3U/KZgG2y6a4fEfUOgJA0
55DinHaulgKc0KukwQPj+xY1XpYAzy6whD65LAOJM/gwAcKqehqVX46pVbmylsi/rJCEysxNn0MO
r7IiEu+gTbEEj0UPdkSiCWcbclud9bMe7LsbUUSN1cel45ahRVEn5jUoY/vX4BiIHsy9Rb9qawJ4
Dls5n11p+jssXittJMovDu2scqj9S7ffOEfE0ujnjkWdNTwF4HJ26fQVuWito0l5Fc+Qf5AFMwpo
T7p3PHxnskyDdtQq5AzWG9nwDJYUxchCHtxYQSgKuwWCFVCN7LIZGxVR+jM2jW7z+S3sQi/31GHy
LvYGSbcevvGy6oQYTgEMWVje56wJcDHu09W54wHRPTdEMQiEj58i4nT4pOhPVPQPFLM9mMbX4p1F
aFM6WO4jRHql2rxD3HRFMg8l1Kl7Uyks2vgoHi8HWWMQWUDcEoKwisgvIltM1LzA1r5PtFNdZsWw
v+j4W7d+nvvk+ZDzDUwU3qcq9C5rv9uuHygDJsAgijFg8AS5WHJbk1m4e6eBVLgN0Auw6UefBP5h
HAlikcix5htf5opU3NTMqckUVosK5e1h4SVEYWorg8nqHepXus4hdneXzdJX6lu3Cuu+SyG3OTfo
JBFRHOCZ+OgqEiD2dXeZkSSZ//J2RojIn+QkufC16VtXPUFa/X7TMI2yIhTut6tUlWD31bgVsehJ
6Jxt/aSDaq/l52wlqBJPI9i6siMcD6EkY8RGBecLhPGziv4m9J2XSy8LYRJP3WDxvQUMNreu58fo
GBIPiUkwnG3IM+S6pQxNvn4KVGrIxQvaa62V8I8y7N0FmxQBMEFZ9BaxOw22pB71A3MQGEZJwF3y
iteByTvzlXITsg6QuQcW31A3uqiSvaPP+1GY4ZVgeyLrVrTGjmBOMYh3wRbDHP+JvL+SA4CVtQUd
KDirBH1SUZWs9HIsSVEkAPVFuQulwoEC/GD2JK1kbnw2p3ZCglJA12R14dkzKGtEXZKwtdaKgzm5
UTfjuysK9mipl8iKKmRT7fSHmFLUD/JpGDf3A7Noz1/hAVZSucJYern+UNdk/qLVZfbEj6c04g85
LIcqoBPJhXyo9ZZy1J0KBpJwAgPMe8eLXw+etsA+sArivhRJT+TEuXjFVigPggYNUP9dn+4Mx8bf
HeEcMud8TkiIei1XPbmuNvc21Hm9QcHoW7h6vRGrTag3JTac3tAM7xX1kkQAKhpL4s5clPcjX93z
vYk6kzD9y4QEBPj5GXb5j7JJ05F0Og91xPxoAoHo9j4Dx3pUZGX1RNpO+dxwTJtfp6U/upwc6KNI
ltKjmljMuWZGNSDVpPkjvxk83eC57oAw04JiXl0UG1DkmoqwWZgulI/AoOQ6JAl34mcihmrNMxh3
pHQT5CAkxDWNt7YzGZLkzJpqRViEOg1YQBy5BYH43x8s+JI0qvXVNkCeHiE09A/iPvVAbgyV+fTa
HkBCQu7kuzYsKdNAnOqW4psbnWgM8WbtJWyjNOsmwJ6uNGMkRBpi5+rVNyexxroE2vMfvFJF4spp
mBqJCMxUVBUasW10YL1zHA+MphIarW0G3mO2XyfMpsOXAaLcYmDcqy+3VGPWxAz1yZUfPRgAJFUO
FvNCBAANJJIU491H96QActEA5NN2avBBKr6UyeJGl39OrOHEFCs6M2TQWQT1Js+GAzSFijlENGnU
agaqHmq3/W0qCLr/42LPjtFYr9zRHhirr0e1lxOZ2jOmFJLrKv2u2dh7pwsdpeG5Fn35kenI2PS9
pxivSg04zDGF7anNW19z/HcbFp07T0sDSeHy8KzKA3BKKouvOWE1r4ElD/4SIcwQPGiW3x6rp+KB
hMi24fafBFWhIWxFCzsY4gUPsaHVS+WNB8zBFRUoR+E3vaaXJyrE5QVVZI+Zyd6uQ/yW5/MPlE6D
xLW7WMD3Lx1S4+mJ5LUsEmtYOCvUJTldGieo6JicMBfotW7R6CRzKGa1QGyaSvp/gfW9SnP7J7Zz
34VJBAa3hydYIKgeMmo+jgAoZDaGg0U0f+iw4mGCljBcx4hW6eRyG3RCNuOBJYjeg7Wd6yPE/whR
DSb/XzR2AqyDYBKNDmvIUrbwZ5DbWlyp7EPm9r/mQQblJhWjWF2NrdMtoWeNzxte8rT6Hx/n+E3q
icnmfOHkCuCDWL+pWXrbrmh4pb/dZQoidngo2hSxke0L77TtCupsR9jvibcVw6v3nENjLTymaC83
2vvRftTOk0YTmIJo8BaiDC6I1vZyboiSFfokWBzgKQDRJSDtizf0d3Dqb+N4zrQiwRGb/Ixp/Vt+
wpGuCWg/0s069C311SGZ8ZvwGDVEDM2ekHZqg7XUDcRXXJCHqRULaKKCAd3odtAhFOodjR2bRdrx
Y0nYS8w+Q9BEeYPZiXCnOAcIWO7eNqpzqc+QjSgljyljru/p6Qi20YdcRmAgwvrQucw+59Bgg3Xh
5fla8gzd8dTZ7WFA9IWAXNo1mnuuELSdzH1L7may8eJ/p9almILrC+uqEgc6h7u7njCmxTOhqGeT
bjm3pQvgznpS+1KThteDXEUxu0CKhHvHd8iKL7+KgumTN4iyoRlHRjwrSE2mv3dd8DQE9ShgMJyb
cyVzIqydVP/pzXxLQQOs1anbkKuP/pl3b8kbF1Q7ZHCQFC5qc8S1S4HXN5LR0Y2BUiXUFfqB60lS
CqETkuiCwgpWkLc7zbZ1kVIq2+pTiKMgJKOeV9a1vfTc1TruogdR0Q7esFfVnZhkjpWVZGIJsCMb
7jjpguBPsdq3syfn6r9K+bOZbyagg2rJqWH/pOQY6oD707P+9ab1HwPCQ/d9Oh6grTleHWyUyFl5
WoiUbRSMHMhxyeUAP5Wu+liWWzW7WL7A0xxqRbEfCxZ6nyJYIhD/kpU9Cyv50ZhjBBAdOvGoFr79
zE2CWkcAWQh6LJn979vmXRgIkYVexQBPzXsa6klaXIW71UpvywobWoU2an4PFMi96FIIkVjPJj3O
K0iUHr/aZySco0Kk8tnBKmP15RhJA9zpqTaXA9lI1uv12v8nkep2tNVy1t23Wfzc4SML577cuT72
WzKu2QnPqh3VuPzhIWTgZOevpzXESNeVMgMrYF9lJrvVyRof3+iC939jX8tU2Xka7f0KeJv9WNYD
zIaUjijMhGq/g0vw3JQSqOId7rb4YjhYTZ6u9nvtiRBsVLNIozXCshX5iGWlivz0OF+jpjTglnYH
yEZN3aiXPYor9HmTucAyVlikd8i+aWfpYHSstSU7K0LWJ4phpYonm2KDgxY9OS/8L6Zvzy2eLUQ0
hyh3Z3uAlpaMzTolaZ7yog6I4Ljq9QDTbWXVHgelVzaCw7GXawYDwr6BX/IDL2xbtUq04UEaItaq
1LzI8GW86iY7zB8LFJpzyJtUHF+PWmxR9I9yvZvemU93Vzl4KC+H73t0njekN1Q1Vjj9aG/AVQfl
nd76/9JsJyB9NX5/1J+25aNKabe8Wkeuo2oGj6ePA05n7MuhfNAA8MvTyZey+a2AbRlv12yDNzzl
f8uhCBC6FHoqUziOmPXBm3DewdQc6vb0xpHuf8EAPy44U5Y/WOZfMxQ1X+HDyJxjPqrGnYN4elnx
pXPoCrJrQqdwDRri/x9b5KDc8IzuiaX8T5sWApc3QCCbx89pXEP3ZOXNXb+ipkK8/XQmlsQF8IiS
VzUTbrV8YyEDe0yhQmNdBsnbk4REkgC5gKb9Isj/aP7NnrvQBcNTtrWKHPr4/ig0YrNcuGkLoO8O
liaoCfZkOjOhkEVk5rf2PcVc5nhXBq0fkk5TRdeJGuL2IfieVPwdpC8f3VeLYNPnacx2NVjsOdkJ
jsyQhmkPje/lBPPnjAY06VQlzaiMQALr/LVWpExuG5fm3PYYIFwT3+d27dMBYIqo/eYYTunoPjNj
eVxnfmNikSWwzE434I7eX5OaGY2SxOBCOfQVb4GH87qHhCDyAHQrhsbtSTFNMd0KAIO2hA0IbKGL
iGtS6MphvDtD5TxQR8gw6rO9A74MesXzQQDtxkWkNg1cmsY/cO1ZFQb+uKhSFYvpK0ap3IR+blJn
UvhNOUm9BilUX8/KOXqzMkg/EaLz31q+YtHS8Tr+n2DNgEEd6OZzgFBMUEpgKUr1vWVAl+sZRbMC
SQXZSWk/pZQADUi/xQc/ypUKnTIqXpJNmlsst1DfP203CmFB22HEVkmk2ByrgTHyiiODCy+uSDWX
vYoImPjR4MqLZ6E1s2jK4L73iQtVBn3C5jFpaLTQPuTRr02ZLqM3Jznu7i4zBDQTtWzc3srGntgF
11XbKM1C4l5eht4brvY849D+J4VvanqXWlJ0VZJtBxUS4UNVfm5Sys82LQKU4iVzWbdjLHGTRdjV
ILumLqdg+nsM2f9pRcs+DG0H/NqkI7eA1mvLaTK+LFqywCITSoO4dl1La+yvC3i934jskPDMFu3L
r3W1m0tCh6goRRtRvQCytRg+MAxkW7m21e4d0xdFG7+8BSY2FOiJyoCIRP23/qmj2E1SwvFbMBzZ
7L/YfbLwBrhhtey5dCms8rKQV6WjPfdETSCKxLJEZVWfnatu5NDtQ4oBa6lnCcahkRVGHIP0i09K
sQbuPz3XLemIOk8PgvMywhaHVyM9pSibCgvJ9bNPQLa7JjYJX1XNxhg+Gv+Rz5FLKwrb8/BnaoQK
k23o/4kAYx/9qA835IXlx8dSmW1+blDGCnThxA2ZSYGYxI4pIQAZrwtupauIcRtCzvnfR5qG/SrE
XCpc5WEw3H6iXFIWjk9WrcQFTMUXMkpNPHwtDvqkc8EPuTjB4sJ35YFYuH2pqS4krGy9YBZYsz9n
Bk7o9kiIfvAUz9HESM0/aCYqw29dcvFOjPH0FCC+XE5QUK09AoC7FHctTIPo8dSdynb2TIthniZd
I1dziSs6JwMTnXShPGQq7DIOqLhXPLE4wmoZ4NwA+FUVc5GvdpjguP6GRjtdLWgIAd3v+sBLhtGI
d6vi0xrxUto6+E6ihEsZG6awNeG0m4eB+JrSOlvsVRwfjZ+ZaRLGkHpggNU6dYKnY6Zv2wJ54Ntq
0QE17w2J5CfxO6fgbROphBAdQ1bx4yk4sD2FBgRL3S5fvhhHMPJoGeumycjdVpHqAeuFbRpTz2Ph
0N6L/UmxBkCPG7UETDnAjUnr/JO3wre46CJL8TecQei4u1HzCjm6pdanOvnpzyjTF9tzlZ7YB39q
QeW17SRIZRmmak/dMfJL27r7ZzBc7jT62gAWnkK53AAQHxnucmASznbM1yLLjWsUQtvdX8YXyJlZ
y6k5veV4kIziLWhWvhkByc4eC5VzcXc/SISpeaiEoZdK2MxF318Z26Tykx1E5ObpSYYgwbB2INUT
NkbTPLkRhjtIPVJ/PtreoIYuTcBkMleiBkDXGPYxgSsoL+U6WPuYbVMIlmFBTy1o5tC5cSJ+iwC6
h9E9DGp3Vz+GsBBAU7jgMtW2VyY8arLVElZYGdb4Kz7bqRdOVUMVEarPeGBVap+eMtPOtvyNCC/G
WnXFINQaZodlmsFL70yc2d4Q7bn/ai+gkcpL3IiFEWb+YTsMImMn9K2EZTG4MnV40YNuaRxIhmBn
1dHNgJ3EeipPxS6qjHUGAxXl+ZYwp6AgC61IOTrAgOX3KyAeoLrqoJQa2rkse7yjs1Szqb0RHEM2
Kw4mVhNemcdVk1OaY4ehx7mBue6DK/o9OvSo7B4eix8PEPGg+XrV5LH1hPPSBg7AU883UMcyJI0T
c5leL8KH4rpEfv7Rd5B4GJfs7j23b2in4T+GVGpKzlKr9Q0+RgPaXC1A76X+K/wkYF6q9J/8USv0
wAgJ+bG6GV/4HLZuuDS6ipHY8w9CGFRFipJzisIDfBAa9oNlEF7TYtoUEM2Oh8aAjlboqEA0tzUv
hbGuGJkmZgOU37vEH3RzNSPeLsTe+YFKEolLWPFs/+8uvHJzyKx9iN8AIJ1e8opXddyTFk0bjYmP
nG+or0tznmQjyjYHNkyi6XzqSMSM32SspDuAJDzMLEPsWjk+iSKiWU/H7eTIdOWCeUp7SwzN3Yaq
YO9RBDvOHRl151+9SMgYiJkiA186EyM4I27pFWzQuhJHZfndkQ5VP9cS4legutWFTcaM69IRG31a
+2bwNmZ1lQOgPLv0TI95InD/2cJtuhKQvPPTHstKlYdN/MgdIFMD4ZrHR/Ok1wbpCtGk8JO/VMx5
MfhXCp1ozP3ZxdBwZBSQ7WPHK1DPfi4YdQi3vsiPSeQoywMN1Nxozqnt2WIyvOqmmxns+I3RJTe4
+FDoUVtQ7OUAqW8luqC/wPkwjoHUL3R7EzLTFYmTbU6JlRA7geYOJKYm07ltIjbvn1sZPYxbFIhc
HpW+8unwxKAw3WbN7TDwN8rSIRILMNds5yoTUqpS/vRlZU0xdupQVu6wema2uqlkufjo8zUitxGB
iJtyEkGeH7/zdp2Qo+b8dp15qw3MCelgOx2V+t5wFZHbVd+T1MxLXCgFg+3JgoB8uUIeJzjteip/
FfHDM1D/ck4zToRXZf8T8qx5RRF6EjqvXp2SYaDFn9EaK2sBgaYdBPkjOrbI634kHNR6M6bocJL9
90h2astvgC6YyQ5cYwPUaBH1M4oSIyAAEvJrpattdOU3mML0s5RIx5t8zrXS7DyUQhBAkD6bodHM
/Z93QAfl+gSeLH/C4zxazwDy3GKUt4D/WPTiwsCTKbgqKSopujfmutbQd73oMGFuywehSEglATDX
0jPd9XtXqGC1l3I26UA2OXLHPUeCLCyh9CJW2ohzkUQt8+nPSvRJ2NPMw/ZH+gNZ1YpvFfqL/80p
OqmP+3PdfdtJFgcrGfSC5HuIo6NQ1OoXoRbbGufm2YGevn5V+CFWrv5TOrF4o1fRMvcHP/5vTkPO
VYNe///6seGD3XXqyfmY/L4U9P4rPG0UYGP0G5wFSrrVkwkPyqHasH7AP2yZeBSG0PDemoNElreC
+FnTuRVjwhYeWlFnitRuD1KM1pdIG4VRPN3RLiZx2++yOw2ZdKGFU6oPsFVbrC8BS3h0Du5wAWeK
k4FSEgK0PN/yx6Rw1SjdABCGoWmLIDAdCaxP+ZbV/3eUcr5fAF1y3moyfKGKdxQu4dz+cV3AoyyF
GIoeJcIkheESLoe5t3C9z5EZ1QCSXKbabTQM7sSz+ia44fFTae/a8bWQ4WtfBu3smbEjadKVZm0D
vvoV+rnRoHstqAN48oPma6Tx8DbNCsJDh7HBILj+J7BOV+s2l4iYNnW+lXKNYNgx3Td2HBZSRwL+
9mVsI+Z0KBHnz9cqdDk30fvPDbR/n8dkKrLu+rhnWfK5jn/otxFH2LPJszypi921+bpfDiu+cTYZ
q3ixkrGCAiQtaVhknQm0cdxixhEEKe4RwfohB6PuyHogegDL3+TrgXpO89ajMB3GtKw6diR37EbD
JO/TIpmIm9iS8Z1v2hQDIGt0Dkq5dG7+6+eVY5w43YM9gHfpm3KEIpgOCSVQqJuzNAkxOCmDKFh5
SMQYSHGuaLfsayIad5PMtmpokPkzBuv1iBsZZ5+mlmEJ5pEnruPYq0lvFTCsn0m/3zmlDMP0cYAh
rdx+b5lfqkOxZmdAyHPMEXaPzfhi3wlhfNsCvLvJcUA9WLNFF7eR0Xq+xQo2mbq/VNKFwEDUEeuI
u75Uac+o9Xe1/ggyWz0dM3vPhgt/29QPwbqwRGMyhOMhYeJ51QjNGftY4hgMNIgo4lgVLdpja5/1
GBqHjWqYFOoZ1MneKoAs+d4Tq0Zo0o01bRpH18C2qpUT8N+JvQo2LC43m9Kz0mh7wPDccovZfHWe
71yscx1f6FOaoxUHPLN82tFvq0ZmBJCT+wif17NgvsJE4WfWtq80DTq7PxK/VeVkmC1fTQyYtq4v
OmoJd0jczCUbWOfhLVVQMFaGJ56UB4pNSaMjTb3WpZllTYBJMpNiax228j0TDKBTjJTPMqAlkbfb
yIoQ+u60NemLjHjzGtb/fpF+isiJwqp6uI/0wQQf9jgGitiD0QIICWXMd23Y/ynvrJMyS90tJlx7
h04nm+YJFJJCPfgU5KcdviACT4vprdsYT5k3oIZZY1iNhamUFKrlcG9QNUfQncwiToAPA/Hj5Lyg
v0cg5MNjYbBpajCLatN6eVCOwHuZDXOOdGCwMmj89X/wQ6gRId7jeGdR3QbCPdaYbhuxYJPnRjsh
hb7yWT3kD0Ks7FxA2S2Ec5Krwloc35S7mPR/8a3G1LN0VWpOMR2d+g/9Ijoa95MJ7VXTcOBPbbLc
aRVQqqns1SIMeVHRUiSbbWVsMMLRH37I46ylPmJ3Z7c7x82/RmdgNe4IUuUVVlFPkTENbLwg7uTI
8UcQDUwomKeqU1ConBYdmXwuRG9vuGucQJYGGcYQWMewVl8xUx9eatCk2ZRlU2R9kpwCOu9LXoBQ
kpKF/c6ZKfgFBHeWmBJm74cFdRMHyogEpG5goLcEar6q/bQVuO0bWxYiHGYcze7S3kaTvJb7J9qG
ZbZvKIkPjIaoWoKXiIdbKtLLkCFaTBLNdPn3F9A2P40l2hs0qMb+OZ8n/MWlNCzYcTYhpRJR68qZ
zWbUBGCqztcW1oFuPJhMm7r+CILZjLv7W4FlTGsa0ECqQurAN7HW6chNrXTIK6MZvwfxZjZVMeOW
7M4FMhWRvyyJ/YQRo9W1QY2fEiggaNYLhQ//Tt1xAmn0RXSHzYnfRZZa9CSMo3Tn4A9lSO3a83h/
BmVxP188AgLjOBeObpvVIOwuVgyWhBl7m7BdeleeQSVKr5XuE4QePH8uK1dGRkJO9GIPg5bs6eHB
uMgi6TqaNgEfDl6teLtPugxJnLCUZKYWhEALjxfQBqx+mMYDCoxfXkCZVoKKlMphwT8gD4hQpaAY
DOP9z4eCkBbr7ivpYbSTDFyjchIQJ7UDxHqtOoJQe58Vw1VrhcNvqkoxQn2YiDkqJCW5bIRQduhX
yKpPYRWCfP1tuU6s8QfipiZ0/C1DRK98u0cTUIkaKIrAmESkihLU2PImW/ut3w7rePgszBz7++Di
wR7WsbkvI3+fC7Lz107Srmefh8iroDLFm9/w3veitkbaG6aIP5kWDKxbaLmYNCAobxaFDTb81yRF
E/3qeX75CWs/J1rq1d1efCFuCdg6oYZFGYlxODb0ik6RK0vwRQDb93zg8UKR1VFC6qCZRn4XFkx6
n1yVSv3AMurnfOXu+0BY0MnTmB4WMXimHa55V93Ugpd0Ka99vV7GcHoJUdEst7qW6OLtT5bmyQDu
xRiA5mqQ8EYsYaWIk8bUlSV/5CMgCBPHPILfM3OpHDFkOMBZJHowAGYay7q/YNj3Q6rVcXJ6dFlE
tT+XyyYNyZ+N2atkkFWOiSlamGlAPpcRJE5oNm4YfrkwIEjHXi4D9D4jWaHjjJvPX+7i7xPBbxTA
JJUJ1FITYbiV8p3bqk38CKZIbQreyYyxTOGG5pgMt0e5yE8po2jD1Y9T5VKuBhhmOptd45IvIvGV
m2UJCsJzAHiSQRuzIafE9u0YZELagxE1esvp3V0C8M6UVda6zlm3C0zHcgPccpwxB2Pvq8DZBXEN
ndxjxc7XfboE/ndgfa4C6D83qH8gPL0QoVxan0kMkT/OSmBQt7gu4mGQHxpXMxR+5ZVr5UeGeH9/
c+GawsewGxVCOrbmlQe+hGYFIqYfwxG7dNopNpGr7XWq+3Dsdeih2k+Zeu1bTRgzc3xKmVhtLf+m
RTooqynYNnUyBmYXBVP16AAGSitTusXOsnvI3FW2UvRI7b/RDoKD9aC5k6B+B1yCWAdmruWSftQ0
8WEG3Qun2Dns4e3yzkcScXc6djt4wNE6HvVcQuUr2Ph5CGep9Tjlxv5TbkAZOknVFpQEJNQohY/0
IUC2sxddkTA05uzl976db3HSGCCz1VCxYVhNrXRpkMQymiOERJJ/8k1ge1oV+AGHsGBCr+/uChXe
dMdSym26hx3XYNME1E+/Gm/TvOTtqVYpV8bL7xRVXQGyO8JRvt8GRydQlvqm2aY1Qj0Ox8lG78ee
S+La9ZmgW4xqn0LsIjd4j8a0BswiaddsUMAsI/wyKk44J6UsmgKgcWnMIJRWq4RC154jaGoVG4cM
noksh2rYevB/8+zBdRaokp2+s6s8CPs7g5aUCc+8LkDNrByV5JD9fcsNLhX0A18J9oMOo5gqB94f
RVPCzV5TW4stiY4kcCV6vc82wi/r5GQACAxrktji+w0D62gDyU5hx7IEhADPFqrNAmt1tgHUcUbh
146HgavV4fywu37a8ot5yKVSw3FB0R96iZrRbOQiKXE1z9XAJFxzNdydR8jFNLZi4HIkKkRZBR6E
q7y8IoAUbvb3HizaPXguVCgoqofmRXs9QCsdQbkfnLXFfLNdSbuyYwQik+2NIp0sYzLX3y8WLi2j
Gsd3+4MXEBVNGjsUpBzFlseixX+S1PK0ACjXesSMeCdZePidmZhbg44yIkY+VQi/Cn9nxLUJoUjn
YAOLxTcpKGjOLZb+moBosYM82M3ZiZ6ZC3ZGYN+lpEBv1N5Ux0cf9N67q+gIaW4JyO54ya27S4Nd
VObqIM8pc1aYh7iZLvUWJ1kRQQxj09RjcvyoEVfhQMTWyBlRQdCpuCbUSCyCLV/hCXDaHXFUtOES
SMgxtoe639v+z7+Hr6bRlHcdtCh8IZEHznk1rOjYX1q1iR0l39hrokgngaDnLkF39meiliVe084t
/LvIsRp2dZl/g4KVT+ZK3CG7+Y33Rr00YKa4m0J/FYDOT9QY9VRQLQv0cfSzYAcbeR8hzElyCG9+
RQT+cIxts+i/y678cvRHqmLha+s+7okq3ICXbRB0IHg4beNaC41STxHhpxq7mMVAuYlT7CfkDZsI
zowmouVLKngrIE/sPoheerOgPILTA24cDOw7F3nuE99KZ56z8cqB+r0mAOPCKrwqhSv7SJo9YOZL
KvFhzSxhl6FB/6KCZW6redfDM43e/mJLC6e6TkUyeoD0R9ePQR0ZVM3cliZEfrVDbuYqgR3zBoQw
Dy6pzTMI+KTYFBrrnui1Q2z4vtWhwyxzeKc10M47S6bosTO1uQc8AutuTcsJ8IAQfkbUS0Vy6OED
NCdQLAJMLyTtmPVHLEOHCC3x7S5Gqy1LAldwTmqspRQ0QgFijP3Q5fwverRXFqrWftlFA/PyRWgq
9hGyq78HsLA47kouTuzUiKsoBaMcURWFdTQ0cKkovd7JhNOXxXqda84FSf3L9alML2tjwVVXFq8D
Q8EYZJtohkHdqoo/AUsBf6s5OPAxtg0qQG1REJIjV1T+O4hdJxzcAZT3Q5nlCubbrtcXdJQiTCMS
25hSwHkRw6dK6STzIeSV/36KINiXh0iDUvR1uTkvtuH6ZNsF2tNEX/xG312G3OVa3r88SyFLKUcO
PKymr8aISoBgHsQ8KK4d0Cw0htA/npkVeNgWfzh9d0CH+SJjVn6mmd5885iyzFdPKL+QVJoJQ7QQ
mzyIJ8EYOqm3159nGZQl1WoXfV33nmEUqHU6D7HECHcFoMJdt6dyb2FJ+b4rZ1uuO+X3A9MtooBQ
KD71AzEW1Zfcx1vI98GEOR1FJshOux35e9+Boixjpvr9DNm6s5sphDxMnuEPPC9kgOV8GSr05wm/
SssPj40b+uPi7FQ9OESch5PbKe37L3y8903LOSu3wzKYbF+FwJ7brPkN5IYMUuaBR9WVFbQbhFdZ
FHbIjVt2E5UVoR7YzHwFNjF7YSzS3fwT6mjP0HbnStuvkbNVAWIN3o7JSc76CJSkcdu9deFwRCa6
imjxpEjTUoP/PKbr19zjvTYOggTiQOAZcAoG9Eo80jwDJcgjbEsktFvhow/39ekcbx+lxk5OAftJ
HOxPXynkAJ0WkOL1VyBdrNJ9PGYjdbhf9OO5dlcS6/g09kVeThMchz9GVonDlQFd4yGkg2e5qrov
bhUGBbkbzpITuqTrIJSrSURgRdSz1/Mu2atDotD4n188Pcyw43pRPZultJLNqrna7+szHJPmgBI7
Bg2gR7C3GtSMvbJpCUDISjk39u2mWrBlgyifBtJvnuAp0e8mdbfVKg/bz1pmnzq/X/7UbXAjrPEI
J73i8CoeQTRqJuhF2IiD1kGwsg+GgsEB+EFuTqMpJeXfh0V6i9c8K0XR53+tpzM2vRJ1qI2c6Q9r
ix71blCcW/WUP0PjoGhMoWIN37sNS7L5b/E3AjK0YD2jCBnyWqREV/1oUln87hm0CQn8sWwpvoGk
cdCNKTWbQ55xOIFRXKoR+1YHMwFCOOVmGsdyGgHxfLJJi8Mj30K8ilE6OuWMFQ3prE16AZT6A5Rd
bESsIHTh9LTCvgvHF0QcE9mKRCpnAuZH9Do/+t1d6iLVssBEnKuc7BQOABYUHTrW4wS5x6u6QMxM
eY156rVoTG7cZzU/bE8hyVWcV4uDZffP0fWpCFzxCDOGOGtRsSpCaN+ngjX50NV4FAX8l+5QWxeA
PzHF4HnMj8aVf6o8Txs3wPsUxLeSRnqHnqeidSi0GrV6UTz/VLMoSLozOmD7LcdfXa1mEaH9HuUc
WFZnfWTz3L7JToyIq/YxuEIZqZCGu+tZdKdMfNELej0y8Q/T08qqhOOROgUQApQN3+gW5pTLXihz
IuEGtc6hl0dFBRfnxv3IvQs7dELfDDm28KvSXSMKBNindgV0vb+/cQ9PB0YlTbddNztaAx0k4j5c
wjYs16udxNTlfM1hgN151fBV91s066Q5VRkBOpTmZEhzeCnh8Qce7FLmM1xABNU/lsYA/z21rX9i
UAaharwVux+z8zejlMyPUM0lou4xcbZ1zX6MJ1+pK7Jz6goE2jHFmMeS3IhUIG8JIeaBOY9oRKuV
RKEFHVqoUhT7rxZZNmXoBIXgPpHxwfOco4VCgyZIkAmPM3HMfBbp6smSTuXCNmd9VDLU3/n8yHKE
IuyWdHJKu7QErs4RLzuNIsl+n6a/JqHfuce1m7TKZupvEmStC3OKw5mIIiY6txStfImDP0ablfYp
xYCi3MV8/QaaOVaR46GbsdpK7XuDqWlW/08qElNPdTWtCNXGjBhdbciph8FMCfrjkDBSDVkOz+XY
8epdh/XCIKSCBmYnQaqeA7UkdeJOYNIGXA7Q7pkL70fqp3Ypjo97ZpGUNvxiNYfvdrvPXVhkBZuV
HlVDcA8dmvFDTyC+Kh0l2B9pQZb2mo7n9OU2HNbr97KF+ayd7sRoUTUWbo79TX2OZtz9eZVSlsHk
T4Ho90634dUYWkHN18fg0DjSoEOYydBiu7G8muv66GAlZbygkAsGyeU+LzYkQr4lFv60tY7T5VO6
f88NMYcSpNmSzD9i03NyU9uFZcV4eljvwvsVseX61i+mU98vDoM/xWBG2OXCH4oRsP0fTDnKzwMB
wWw48Gt6Pjp5SbE8TeGL9iacY8+hGjPC7DSnF/wu7ez3cVXLWbgeMcyLWanBH2dTaDeVTtOchRf/
IbTmVrg0uxLuHWl//6teZ7xN5oHblY1ZjqG7sS9PaXBe2L4zPR2vLPzxa2BOBfULlkYZHsC3QTas
v/YQxON4QNQ6tvakT+kE1bKpGZL/S+QbxXSoflNXX1A7FOFl0fNlDy+5bzZh4x4UGwkXTcs0QpzJ
20lXMMoST64HlixbUToyvml7wtBTfXbVEBK+W1NX8BzGWcHYmapufoiZ7HMZOkAi1BP2+0hlvSgx
sP2sYCpcBVCWiOpRUe6K9USVzq9TM9tzXV9TXYn8CUdpBtVQvXVsIr8S49IhcmqNU5DdWz+PZM7Q
4cY1pL8i74bjL6gSpzAA6CivsGrye8y3E3TO3KI+UdJ6SbmM1npejVSX2pA4FnEMoJXekYfx7pay
xgSooc/Hu9b3pGi8Dvos8fyTQ2dGjU2laDCibtJANQqT358xPnJ9+BK9wNhL9dyfz9/f1qY8xCYo
mVyBDBwgYc7t/iBlVTlN3k6WRpQjQcEtOLIX2ytv5F2R7jLpB8g9yogu0Jb0t4xp/5rKlfzxewLM
nEHUU3FMsWAg8aGzDXcFKOpsona6xUI/tkhQmFYAZZdhz6zxjwgJw/k7A9jkjnf43Vf6OM7fAHZS
J9Nr0o7oj8pl75jHQ850qqVEd8Chn2KNZuv9ZDw8wvzlqc5OHxGbnyIaHGHdm2EFJOTK3quxkk4y
Y2+oDY4SlfNrL2cxa+myl9FWuhZIYbTnuEi8ThkK5+ko6KlcY3k8VPxJ7vJJUNW2p9IkN61jqKpz
uytRrV44pEvfcbUFBwBxblg7Idk+2EU2rS8Eupty/i2CJ5iHgT9JY5OX+LzMFwVSI0wCKNWY/jLb
7sBpQQPg1fUj8Dq+jeju45fYV1PYXhROfw1gfkKWVvNDTcHrxr8qD1E81Syc1Nokhle2sztdOMrT
UFc88qiDaTqZvaHMAqnUu7tZ23roroiODZyy0HPRe9234LR+8ImjJDigmNlcHFAkG1Q0X05rgaRC
7yA/pZEuuY+lJdJlNqzGnmXiMp52QIPxoo/aoec3RaBm7VcsYntT09dqwI4n0CE65LgiNMIYhLng
fXpLWU1A2JWOBRjXLoNsWKOagSdZ/KMGCqowkMBbdp2FWZ2Lp4u09LPkCquQFvbOMiObc/V5zw9c
XxwnPtY6Qjwh6l0Ys6vnu7/dqr4/PB8FZITpu5cKBUfhIMUzlwyzJ3kJMHXHrPO8FJs+HM4Ik+8x
5qKjTjOQk2bTJGSjMgFP/73LOMWlSsh2B5U/GWdUsR0bI2imvCT1JDyRpDxxhWKb1LbdVdXn6P1p
p0W1+nrJGqFJi0tRDtA9uslWzbCUn01ZuwEZ5wVNpdyVtECiQJo7GEIOlgV9y5F7uzIGfSUj1SF3
zn7p0b71X9g811ecrPhmLKKMCQmTkg8DROJ+1TEHMzwBklrqW92jqyvok/bqjBRK6Qt4NShB4o44
6g7So7nCSdc3+S9MbLPytWLruYInV+0vopXxBqwhOhBTFGMdpuoS2cpJqkXM+wMj4ShcMHJOEWnd
FVCwbi26i5zyGZQcML201VX7LxbiCgLIS3U+ED3n2yVhV1MWDWfbFewng7SzLYJ20GhpG1YRE9LB
b6SRsv2Tz0pm4A2ywT9L7tPSilnsIOiuQr6RRuf8bSuBFk5erGdnYj1d7jp7SJBIIFrydInT3x0h
gb19pZB9kozA7xU1MP8MAYBhHGmLyUs4pVHJpt+75KJbdHiNyZNUM33nMHHY7SMPCTulYZ6AYIaJ
xowIZAbNDCbKwCAeWMyS3/F/pMDNg2+fVXabAYwHjamf2ejaySESZrKOWe37uRAXij+1tfGlE0E4
mXyFWhtGuAbU6d/mwpq5Kcab7v2M/rKXZD/cTDHdGHz2Y+ypNkijOzGldJUcDMoRYHJL7D+TfU3D
RVYEd6Wrpy/tIEkXMQMAL+/0hTjaeSs9hueYSUBuNdXQRAAKGjC2j6e3NY9pr7qWNZpAEBWZ3sjC
T06mEarj5GC0kCMIs9yQVfX7G10E0r2NF/lzERyOY+Hyp6dQxUYqTbFi0oYgR/yk2fEw3/b7NOI1
0+yrBNF7ps/tCgsvGSaJPCqVHaIMdPqZwkUjFaYBQIhx84irehMZshEdGop3YzvjbNarl9Vj6eGD
SyoobHMX4Lb7Qfhvha00vFhBP3UEdCn5JFc+E7Y9kD67EmkhMvIb6N0RCUem1I1eQeSM0B9pOq7p
fN06TrVVGoHKBktfQxAZsWwonGz3dwBBpPntcwliJ7uQWKKJTkgHsm6cbQi6RiPRr2V05byGGFfP
/35rbrECziluLTVHfUgMEEkOJmxOjkJILTyke0Oiq0f9LX7Te+UfzJ02YYveSw1qK6+cW+FpM2nz
Pbglf5yIpaitepOxXT815TeadM/9/y6/AkBtClaJBgL0JiA5fqQW619PXnK4jdJr1JRxCG29YDln
OUpl1TAb79g9x1BOn3DJUoeuoEsAfzprUdU6cY1JkIwDigacciEfTgvgg/aVvQzXqFrXXA/xLhoa
ZQahlFMBJ7TvhoJUEdgFy3KHwleO26gXPofIX5997ucpGnXgPnvSanDjNIACxSFoq1pfae8mytYA
k2QyfIRD5gdfGvE8KmuPbCO7tcqEra6AgIM7a+ma14QD+zIhKfco6ynXNgkKPgEmxuv6f9FWNpjm
iKagvAuBrEyqJ6gMEOjjmJICEFtK5txquS0n7h7QXQGkYzUsnT2f7X4FqTkEXd6VUoou9Nx76zQj
Kl+D96AdqMZZ4iXyAeDK4VBoZ/W268KAjrVxzajgj/ISlV8kErBOJtnxHW4kHfuauK774flpOuS5
c58m/xqeSW1kXzw8abRIYm7T9Y2ZEeZOCNCJlprvVVqO/zfNUlXCVm20RABDXNl6alNLv53TqPOw
gJA3Fj77GQk7mGax4Hc8TAaoNO61XlQPyW68tTc7RO18nFe5sHM+oXOjzpxvQBNxiu5ZEzD/dRbd
gpWIdArkisXE3qMUpFF8ZgOBPS1PIF5ksDfk8rwxd9krI2gs8WKTxrPmoBornAG6poi1JRXn+vIw
Q78v1E2ih5NM79SuZiY61yxw9xRG0k/01FZVFUQAbOPVoDGEL7iaD+DqhI89Cb23eJduhSZjc4fn
pwbIpxjSrK73dQKJuVN/nPMTWPhFh4NuwmoQxrYkRKrFkbEQyiUPvC6rUdWtNA9WH9cjLNvG+tUi
Y2YlG3fcng43NLOe2k2LtlIZRFIyhp1qmOsoShnivctI2qkQVbCQ8KEF3iqm+8LpTqFxbFek5HzQ
g2ZEcMOabfzUTeCOW54ba/t9ZCr+qn29HDZJPJNW9Rf/QfRDzwysjW+pwu4FnX8cFz8IDKeBqGo/
euVKVOWFLYmG/Ln7bPhlSAyeyZMlRopN08wgFpESedVXWpLAz1ScGD+2XDXKvlVToWdTFNulfem3
Zi1XWfklqwT3JWOmNWM6HgNVOZPvWDSyL9o0LvgM658YxVjHtXR/6XfSU2YewqO6FCYm+W7Bc4jf
jkDh+t0N9J0wVQl+Ce6V7gkMYosczN69IEAKV+n4duKqQWDkWQhgUAtwKVbCC/or00MGHv3pHfAq
kcxWQkIMoI/ufsPl5rPeLWCLb394vFrD7s2a5UoJm1CxCuIKwifTcXyyHHy8e8MpxV7KuhhYw7Ls
5OSob60tIMVQUI9rOeewD0WV6nPkj65It3iP5uVjh7VRoZw05SMo2Lvo+Bh65ROXNT+Ry3ftN/kJ
v0HxbVlAfzE6z4ljP/4h63bzR6lDGCB33S6RONRUJPgdqJ1v7pCRiYzYmRuk4wDXUeoXENzF3lXt
G3d+DCIVAiS+w1jcbhML142v1E+0KaP53SuKzYsKuRlJxHqO3GHsnTP2rzIRm9x6gKfdPDAz7SNc
qc88S5SDD/2rnDpowc0BQ0cyif8p4lbEQl9nHvhgM/BqEviKlG4MvSEVmkXvpiY16KcrtwLyQ3jC
zbHIfa2CjctDONAmSzUHnEK2lKLN4YZLXzeS3fMhH451iFzOMcWm4v3kT/YgNgZdHqGkLFfIZ5X8
J051vCp+keyN4o7VvsY2OxPt2m2DyU943bGhS6tfwP3QB1zaUwrC/74AIB0/7Gb36gQEo7MgMv62
nsnhKIM7ATlnHJLJAdYpqWrHwrU4ngUZrP1MiNgPyOJOGr75UCdTvXNzRERLcWFVfrRA5GFFZHbc
1R/iSfLbgmfWbxF7b4au82SkTAb9zLWfeH27NhKp8qWo86/AdXzeUCMHt/QZJB7kcSZoBgBt1d/y
vmWj6dQnIucIJ0aspbZU6DWVLQ7M8ylU+H+Pn3AuBxJmUqexpF8EttPbGmI9+Z95zJRUxJMxmlPZ
abg5K0z6hAe78qY6uCEO7ShtGLydhfTWmuEm/PsoD7M0mXftuFgOe1tOTBxRG30hQd7NbBLqPbZP
/TaleyyL7+HixUhzsHMt5Gk+Co/CaeQ6LVYK9WGWJwOJ0byjWZgnm6Zhoq0gUhqktWdJ0KpIg9ly
ZPxf4TiXiO7c6tNnsWVtJf0F2aBRv1FN6UfcWduIG2SxDTx0KJt6NI6p9H6NXg8OfCdfozCAg8UP
IVI+ILeoxAgUT9H4pkcxy6bqHwG3iZn1Ogc2B2qjLj4RcIo/BWYFMjenJTq2wGaUPEzto1eYRnex
QLPqXoLVfua3YomAYw8Jvq8JRNLPSD1hZLjbcrwkJ0ZTL/Fexbj8mIQeXiYCSaUdJxVGbz9SsBnt
IZnl5CZzE9q/AK6Oaqvj3N2KxsH4TQ5eBdR9fJhv7tCND4c8FyY/IpHehW5bPZ7MM6Rp0X/tkKtA
XOVbWkmaJMpNz0yqspiIN33kLlAigE0yYsUriMvbri7I9jZV0cLhwLEUPQFHkyt1x4FMYSaZY1fz
mcHllzaoykXhW9n5Rarf5QGgfyGxERMdZjV6GIz7eRO6vqYiJ5uyA7qpWQUoHKWUDuhN//ffrSV8
mjKU3FA9CFSbKYod/+prhPXPu4c8HpmUrxLNGROleQaCtNM5sKGwE4tUiOrOw2S1t6URJmd01v3X
+hUsxLxjE8rhTV0uBjcBY0Jau3cvZqESomJm9STcKAMDNI/uXaRCmztvq40Roz5r1iK0w2y07O9G
jLDWA78npcaK8tcKkXUqJzx0QFPxQrtYJh/0/X3Ck/oEwQt9GIgwpVrSjgQysBYikQvRBOW8J/S+
morJjogke2kO2BHDXVKxy4+05Y1GoI1qX+Z8uthjluxce5SQ3Kf1/zRwKxrCIWmpnW0KC0I/jyR+
Hykhr6tSqitHRS9s04sbYB2g92dtQnQ5w1JrAD2M2k4xluPlRA4z5DBeBS4cUY18hIxdfSS7TQ0V
BQ/HLY0PEvkRt8MAmjelS2lwNrzDHFW6OZxvJqNpwE7MhGi64TIzjcf3+nUDL2aLx0HKxk/bHUzw
J0Vy36SYEgeRxUAuYoLJLyFh6eWyDFlGndv+MtZZHGcHY8Y0h+ZaLASs1qdLTl7M4JFOZpqnzTZ1
89/jYOFdrRy2TvwX0dnHV84QAE0trL1RwSH2tR89LyWJ73pXXenGhcx0rQRj2NMzGoed5YDZnZq5
xQ+TpnH6vvr5ty5uuJFtwtjADwsJip9v5KJLEknqiczHIgm9LM6/pqU9q15l+kPmTA2ZCjY1e5y2
j5lEUlRyMszL4Cs46iyw/7p4tcqwAbd+ZDkfAzOhWGGKeK5IhpeT95zhXbfgJ81KE55fdldg/pzt
A1WcumBHqpIknDqn9R0WMpmkX4mDjSxYYK5EdRnHUB/D2oASeCmzZ6c1lIsUQD2avmOIL3f66hea
uGPBY2TGyGzczoopX7gPpxR6E/dCGdzeqMz7nERa2CY+rVQgeLCdLbBkcWCxdfqjauFG/jrbw8UG
q0zDbtXSCvXWBHEWJpAGB82j8P8OTiAuBqsbrFLTCcHS3R9KowZad6Rbu8iFmEA+JDXLDe24kjjv
S70ixBKaQ8q9N5sxacGGc8pZLTRZd0NEVJ9iGfhqto928FwnA0RBHZzNLLJR5tw91aj1xLq9AGMz
1Yc6S816dxPOK5n0ziH7ARmxs+pR/v6u2H7mZBCvDdLpcbLXVIv1ywL2VHJOxosBaJAfZYCHfqA1
qzawRYfnaoyG6hACKW7ciAtJx82RdcQxQ2VOb4EPXzSK9l1QNgubShTqEb61toD0Y3QLacUzaug9
KhJRMEkbLSzKUjJKgCD/wMJGaUGdu4hYwZMVDmALdJL9aXKJEOiVwdMVar+blVrH1cOv9++rksTZ
Dg9uDztd4aAchDAg0ldacWlnHzhLfUl/TO3ylg5UXlUtCwBfjrpc2wvBVwwYKZ+e7rGKQtiseBNv
58FSvw0Oj/xK2hE7uMLw0d/TCAF7uluXBG4tLznVlDERfwkMfHpk1r4oWtdhYj77m5GLv4lzwYhq
Av7pOewbmhQyiFKsPPD1wMwWGZxo+yHF4i6ghMQ1T1yFFGE+Vr2+BWA3Uhq4Y/QOMatzOTx85nvk
GPSp6rXFhtY1n/xTfeJQmWQz3Vh3b69HRpFOcPTRMEVO14CLh7DyZX3LiFYKTqVvB3Pjl2Ne/ou+
wm+KRJovBshtIf3h7VsiH6h/vX4xxu2DeSepPPl3fKAkghDNL1jv5cSqcu1+BttEzQTZ5Fcd9Hze
dIspGzg+LLlTYlw5NBnHCjUeHEhc1Abj4OsV/yLpXcxnT1LftPWX5tXY2qMlQCjXiiRhBFgSWmIL
uwIgWivBL/cN/oFRPNWHj3dRWdYuUYfO8bSsobGTsLdQmIRZkcdFyZcHaziF3mhEnDi6oSOGm9En
qtozh+XckDR9vCxFA0YPdXokqJCe+dNqc6JrV3HnsLsJ7Gu4JBnIDBC36UB8NU62B1K61WXSWLTW
IqpLJkOoHPBMdOtH/u9lyGqV0RgnNG34yDvmMrYvXd1RgZDoEwH4YcD1nHTHiz7fXL1PlounIb31
ef0kd8fQ/yVQWOwaugHERaNyJ3nZlo69Oj5CmT83hoTHkYvHlydGN+J6MMEMQKdkly0DtZ3zGy6B
rMbpzFB3KV1Lyo1EnNhgk6glxWoj6MgTLR+o/Z8msu2vxKaJCGiBavXgCtlChN7Fb5tIlKxhLDnk
oWhacEI9nH6z2Q8/TjUIJXj2r7yRknatOzNRz6CX1mZ+Y/pULUTEvvt9D3FPWgDkXZHf31VuF2ar
gTfhL5m1OLsEfu5bni8Izv2OZbX0ouz8zN10XHSEQOR8mLaDeSP1MkeUT9h4n7iiuOG/40Oy7+1B
UUnWPpYGtSyarxzpRDuHEn53wUoFo7HMicY//uRijf44eg67vDae0OkCHgwDVHUTZT9Xhw1chPKj
QPMq/HcaG4+DD2PXKxKPuaiGh0osXDf8GoxapbhHpngel70erZed9ezHEPaVYlHQTa+dOFD6+zuW
ouVgB5W9mDy+y4ulpuW/imAzJo34g/i9j/cDheOZy6NbWT+p2thO/ZXMo/tnGvfs9ZGwSkpBXMCz
U2PtbCjcCQDEXOWC/uhuriTIOlh/mKrwKVEvrl8c+et2Y5I9vAtRU5Ga5WrDCmwcR76oHPArbMcW
fkhoiKUIZK1sCSzanPwr7NuvFYznBQdQEFehRYbzB23+e8qT80t7n+W5gPd9XZHT5aOAzE/78p+N
XQhTNV0BO4by4a/F707pZQyWUWQAVQnoaPgQAJyTckxBO0vqSmLfZ2sS3C4v4x7DzBRmpIvs8Cb7
VDhhNZRrSTNykPBY+qg20L3RKVqD+oMiFX2uZQr96u9UuC9t+2u6goYRZg+rbWln3ZOyCqPmKhAm
J1i6NNpCPULTbvyWZJz2HeXFL87qxmPQSxBBe4VDxrVHuEbHBcH/B8MLjDrfmc6xrLGpUTF8dP4l
0AvadgRFamKItdOrCcgFwNHWL867Cu+X9DQ1MD0DG0EzS7dgNnVaLUxDOvfc5Jpfebm6Ahld3jq0
gL7Ax/WtvPDwad9IKSpSCvPI6xlo2d3Vbfr+TOCaO6h9EL9ZXSj3zwDI94W1tCVzUUelvKU1EAAG
63K9s7loUwDA7m+uUn0u/0bnuCCXq5lFgucUf1UEc/db3v2uOb36gsmpHGH8IkDVIr42CYDYoP3Y
ODBaCP9M4Zor+0X3xNjxSlKDNO+djHM6CfxtIkpWuFDrvm36RDEwSCnspbVNLOIoXNiyAQrZu1Fc
75iSnTAm/Awskn9ko0QrgQWNWJ1QTzVTvzJjlLOIV2FNsaewVww7eh4suQoVcQVDsi1Of1fMUfJs
nWEahOeM9/WaqTTTwdxnksIcja+ESed+be7vKaBOK6/3iHIbIFgUG+FU4ZTIoilvqw7w1SPlOdqg
UKLXudhIGcYU5k3eXuwCXYFo7evrmxIqSw63TdpLdeKKozWsnzc7+oRNB7Sbb7AIN7R2hNoLEVbU
mXFcn9W6nogiqSX5xfPn7NDFdnmO+8570PtADjPUHnykX2FLYWkBUNlVPbRg/lOAdSGV+cab87JN
pqHKGJ+55QiRE9E7SOYDBW9mIBC52loHjB7VzS3J4wOOdQuOAa+e1pCp7bLZWeKoN6Bmt8GmoCXf
vfpogDmWXYMv6ho0BeT3wNi4Wss3jjoPMxt7zqnnctuc/ZcaXiJslObK3+0ASMehKWyzSSOS2wEk
q7ckhhPVGJ94WUwKA6An1ZKECRBkGlvrUVdqdjYPazxEx6k2RSifbibvgRuhASOKDXbpFonzYoCC
/3q+/bTdNeoyu2fAaIBeM7qJkUJkjpTJo0u2nTVK5ckkfXMFIkM1gnpzM0LoOy8rNa9/pW9aXSk6
uCIU7tC+63aX4hRQdUkLo3iQYQRzfd3I6qaro5dJxdjnOrOfRCnFyLeOVpYFSMV8sekqIrK0s2cO
Hs9zeGpQJ7E7YYbG6B2NhlSdYWQ2mpsWooYT+luKhRI7MZP3cMZaHNi9MxdxwXl7OxcAZ4B6n1yT
2OsoGwCdKiuCwZeqbalRk5nWf0tr7YtOY1KsSz1Xej/nj/IVbS+sV4SV9X1tuCAwGvgzndlVZ+FG
yNriMbHb8OsrV/VN04JfG3eSxOdaZ6+0DQ1Vi0I9RpWyHPeBO14Cye7e4R4mo0rzomIJ9EXxRSPs
fsWRo6cIpkqcjvhCc+I8oW1aKH6YsrsHS/7K4fHAtNi1c7UhT8znkHrQps0sRo9abB3hoLbgJ0C8
ILhzWze8oeqC+s+kbu/AyIKe7zo7JjbpvtTAv+6RMbOeXsCFje2Bo6Rn/9vMUKcdaIusYCMezw76
jAvfIdZFaQ6WUKJK+E9uyHjTWicmykfHeg1GNIhupnBWCVuOirVZb/J1buBDPWqPuMV0MxlU+3Y+
uBtD4TgNDkjniHWz6E30FhBg3GgwlzpJYCXC1qewV5a2ogiqoZB8AQEE8qkxhLKE5+SxcKgC7bYj
WpgX5BrMtaaekPdEat/aesK3ux+i6LIbyYbZF7gtO1MWOpeMhL2t7qXxEckdjhP0nr54HDe9sP2z
zy1IVSBKdvaSwhwJ08gmNYOsCQdTWKlorgdiA41jeepYZ6r6tkh02/3c4yB3K0j/F6w/+l3f6RYF
ZgCK6c8cKvLT1g9pVGSBAJC8W4GR5ATmjEbIwyKJacRenXDZhxayW1GeiVRFE8sC3bayo13NIcLu
taOGZZysBAZyaFLEsSCv1EklRgETupGRHq1LKLszkTmh/J2yqk8WsSX4HwftPsDdvZBULjeasJ47
FpbZCNvVOuOH7H9YEkQJuZDsbtBFgZkuQe5Yf+gnqMNhupkTmslWrVqov78kZo3RMq5eIX0Zw+Sz
87/GaLvrHaOqeVyVvXLwECJOPuxPo0fUyU7FuA5fwRnwsUushweAvkzksweyb+GO81P+V/9a4z9a
Os8byJNHVC5S4Q7Ej8RpEKKApUpqCcO9PaiAoDHHe3sU8Y8C0RNzWreChcUb7wNaWGkDSR+gNMMK
gVpolnTyM1tPfU/ra2snQ92sEHzGKY217uwc8BGz8ZRgTC11aXSLtX2gvBF+W/cj1aO6GiVReztT
zsVC0wZdQsEkzqEuLHJoyeuGr+SM4PmohLR1n0boIe3dLDK6Luaz8uQyaILsNHGWIeRLzcC7uf6B
f3C0NiG5YqELqU3vvg7rzw2KOo4XmDmHfilasGOBTYw9cp0Z3xPD9KlRu2Pn7oWh2tLXyaScLeYx
95r8DyfHoZns7JLq8M+kCl1MBPC4zuwXr8QvfpAeFH1Fb5ph9K6Rtju5ESLEFW+uE8b9ZIJmIUcR
KIL4GkcAOC4byU/nOZdS6Ra9vHbAXVyYrKiBN5r46xkDloNlIPXpOhkL6PRn8bdf9MCz0rW5rX3v
Y3Fx60EL9U8Ihi7HLNpQbTAU89hSOrO4XzaaphXSJln8SN0A6LyU971Lev/mNg6/Lz2KmpdtgW9r
F4YTwaUT4NFarIHUwRVgQYkr7cfqr7zm1ZhBJDuBsHqc9eYYl8SULHGEZUHzPgjKwLru6ztpaaRx
gE+0Wn5CglRZnR8FrvALfEUTaWBwelD1OWy27LjOsbj3S317K+w5pKuE3lbl69OkkPwaQT0bgYex
rE0uWl7UzEDx17wg0K8KqeYkGMKpIFAjtV+2NrkNE5GqBx7IAVLgaqVDsapB4jl//qN+yZwN7TQf
xXlKFFBkg9kZoz5Ta5q/HrinwPbiv7Tr6Bf7cwmLUlz7XXO9DFAiKUDtEQsqsu50PGWrMDjgfy5W
F0kFMPkSTTyZ41vXRqVvoEiX/Bw/EbLaRfjrr/ny0sANH4UfbUTkwLLeSr1vL57hspN+keOzvV6a
KIHTAHqCwal0/S8u2hXStQFbQbJkZtDYTYwxdww1TguF9X9cWc11Ji80WqXl9MWjwkM+Msk7lTo3
ZyKrZ16soFRLa/I99p9Xov03Qw6hGEHX6IfGbiHIOITSEmtRSOWt1zp3s6we79R4aYB7Rf3EfSzB
fe9DBeTyXGKR2frswW/7yg1kdTcTBWxCvLDmGjyHDczPjeCDoJf1AJosrIe6X7iLVNzPt7oYyraP
ZjEqI9ap9pbbmyrujkGfSIzJakrDVA1vGArpZ46oEd3vOYQ0fyTcsF2tDPHm03Faa8BraWLTLVbx
KFq3d56J+cegusV6R4aOsEbkmxrsJozfFxc64vCZyDc6XG4PG3MgTOYpDhLJqYHtvGJSYJm0PSZJ
pZXx5evT+/RZoZNDX+IuzpiOXF0gzUEBxGN4jWPrLBpWhH9kLQQDsr4lFnZi1WM+prcHhsjyQYZZ
moKs3vpBDTkxuPveSINEUtFB05u8YldKkvjZ0lkeHBHYd5nhVxOuUQsEju9w+r2FMhv4By2loXPG
XEVshySavdU+8br6rpKN3mJw0cepgiy4B/5dyEnGLnEH7v86Tzn440ptNvgGn/S12mPMaatkrxnR
QhZYBB3grPBwI///CSbCQ/CWos9k+5GmxixW1NJepUovABgWjCY/sO6M4FhGInEcVgTGUv6o81PQ
hFwR9OOB47wkCTgyfp2ZAlyS6g9mVGvm4Vty3kI8EYPFqUaL3OTzFWmETHLiCBiHN0LieSIEtk+f
ji3Ew7p9kO+NG81FTaZMpWS9GOSKeSgTbDTYE4pfruE63U5OzfaViXHRWatnwbdIAsN1EW9LYKNW
tfmr+KNwQ2ZRju+LfhmnHNdJSALj98QzOfKHYFMQDacQNJPOWj+1LPhMe2iFe4ekyor0AmU0TLje
UybshRFBx5J6+IE0ZfxBX/5f14l4FzuDk8xyP/35UyniC1atF5uzzeAPfiv4W4gpISkuwE0iWFgU
6U+zVlnOu9D8ZImrTRBWPa4QWHjY3PYuPS+/jMrMGpkz8KtYnKDtr+Qh95SufsdicD3xgPrlQtiX
Q4zuJuHNO0AsDk4Fj6Zz6s80HjmiAMhn5tO9n9J74WZpEJ+3QNSC5rjUogWgAXzahhdk4/IILzqK
eUpN81fLVKCCGYfo8cb6nK2cP1L/nOXLhAhgwDfH+5w97UQZ86gqZzUOJTIPqEQ8ofzcOHvOOzMa
h/yVDDVeThAPi8+WjW4aR1HqQVU7/bSfiSA4ETE/8++hejiTGxNmL9IBhdflMAdnt2KoHZGOgew4
TmNni3q1kEqt/u+KzZ2Ywbyler0gu1p8Odw86GEkGH6J6txkAEXRfXWdplyLolDeQb5T8FtL6pj0
KD2XaaiJ/md+7mj5w6EPw5qskwXd6Wwvb3rnIq0oQgy3oCyxU51QzlDYL/6chtzCuwBQ09rdCTLq
2APu0sfYI0ujZ6TxDe0JkkDs7Ml9GJ5mWQd5XM0z2NlLqwc5ZwPhbPKkpZ+OXXVouctCt4JVeluM
3/Be+3qFcuyAwBxv7xcPqrRK/uxBjzCHE6x6lfFsiOHSxw/gQrTFGjfEFkRWO3oi2bng1CmCQzgT
Cd62hkW7Ilf98Gwc+jHxqNZU60OqxRDkhrtdeNidixeBl4eAy3D2xoS/wuUWRO3DUIcJ6cQfOGVf
Klj7iC+Kj2UH5w5MGSnFwMzlO5wX6RSBwNceUAlCVrRhmiYRyM+nbjIkC6oOUOdvnenldFfS98La
vul876zG1dYa6OYB97z56OQGsQPLE0YrO9RLxAJF/n6q3nSpxFqbZIqSoCN/ukYJxWAkjMymvHq9
8bk7bBZaAGOEobGmYhWwt8mNDHhMvmAtFEgESnYMyz+ru7nDk4ZnELuNXIRF75ahpGI6JkSGgf2Z
lHSwOWwnYH6VU0zpspV2bSUriRCIt7ZrMoeOaIBZVqrrCCRFcbENAZBetXa4/kucrmVu8UqKrUuu
rPf19Tx+nk3NzR/qRPxaNCMPWYf/i07XcW++ZUejgGwYupPfyBntP4N6owY0yw646aRGVc7igsph
mPS/n92ruldJKpmq+WKcdqHDBfOeHcjLUJBn354pDv3h2inT6FRbmJ1GRrVqDpy1IHszN8RJZRLU
3+pIufqsstGFkJfG7nyAEsA2b9NY6rhGXJuMnSrkjEYTVV5fpZQ/TLvGY0bgyGns/8Bqg6Hme1To
pw22ZiWtsg9YMnx9nowuf2CBBSVI6vwGNmiNEkykQ6M1tmUHV9vqDoZ2RpP8q3BX9vTK8BoR33t1
o4Jga2HjSgQJMVRVsaJLRv8QphKiag/K3qe/VLHDNTgl+w+rTKHD0/jzoaacI6AD+/98kQM5xO5c
r60zgT+u8p7H/dhbtVafe/Pnapk9GkLZKfMdsxiHGFz8JMiSEEbj4+GuKGHmS3oHDf6UXivmiLcG
ta+fbvb4m169kodPiQEqTH/C6b2iAbvfEBUmRWdCp05sxVIQsEPa8ncs5XHU5eO7mWsS2PJHzrUV
MDlQ07CuuS9ZPbwhWI0Sp45v2Efr9UKRVvQyb2H7VdUpORYERXb7+pKiOfXs0VYASoyVU3PnBAE/
M/fYT3OSFGA8nPUBqfB5tdNsBIY42qlsbzoiXgUsN/fdbhndYN6STL1j5RKKLNzLHlo18XkjPDc4
NC0Oxq187wphX4Ro9GsFlHAQ0FUnSLVTrmX2rYYP65Hkk609LYqYdtmbfR6XF502NOh3Cko7AyF4
mKaRIFpaf31t9iM2gghNgOqNOQgHl4bheqCDjqzkrAgLM4apgUKUNB5SNqTtsadkX31W9HQWvlrx
6aUdG/P38M4p6NrzulrhX1gekpqxu+GXwHN5GCtT1FilWYIySskclHhd5xofa3xEx2COOA3FATUM
DwQrX+XhWNb2WV3iMXU9QNJb8c2IJuND0KrXjOEFwMJKny5l8q2yWUwjIANd+0wkZJY6IV/exWrl
gBRDjzwIqhKUEKiQzhrTnrYpiZ4sbJB+qzHmkw/7F/jsEY/e1ool6kFhVpJca8P/wbvSkGbPwmP+
fwxPm5GPxxjtwqWKUYAr/xAVFf/3d7oVBUZTxtr0EAks6xmRnPHgHNLDr5keV3AgDadj+XEXlqCh
z00OLTPnvxgakrmT5R+vXUJsygpDXOK9nNsSGBsu18q+I+0qYva8iwBKefCRvfZYQdpb3W5Xw5ec
KfmHvWqDWpexcvbBVh9VqNmKNyI9OBxkxN4Mc275F5Qdm3ZciPiN7ua7KIp5NRuTS7YNTw4Vyiho
AOJsB+Zbx0pZmKYLQJdrxUDulLnlzvvLYaD0uX4aGt+WrnAfpoErI6pvZ15iOe0EA02SuM2WJ8bH
QUF1DoQ5ZszxL3zvkWaPOYy1tWXzQpxFbpWtqc4+a1nDGv9ueSoSsdlVghY59Iejtn6c1RtAX+t2
FC6ZES0JCV5LTWTUWn+50AF66aL8Q8/wJGMqeQnOzroJEd3ZsZt+sLfQnctNUgmbuy/+hp4QOmOB
zaMIBW5LrcsQnjLM5auv8TICZsjjngb/BfTTTNww1jdLGiOok3bPE7I+f1qQynGUyOLzmtyM5uBn
90oovddJx2YHAk82INUn6BaLwFBuyfJ3sjJtQqNxNDlg+5JHZsd9u3wLpXP2EPsZEadY5oF7Lve0
Jf+jtpbYPW8/gF4Aom2C8klInhLoMapZ/xnkgDpxMK3b+QgeQuwDTJk94X+e/q42L+1jr4ibxdLZ
YRq4muVkusq0WhNGclR5C68y2QxAxSOdUO1lvahGQ7MeQDkS3RUFAtZ7FeW1sKvAxBb0KCq1bbp4
KzNnS3sUfnRbXkianFXO3bGAtA55riZyifGLFVaNUpC2EqTF3r0kguGMqFmNIYFVUVhNI1rNYjN+
5LbQY/3V1zga8dD+ZaOTmkTHiJkyl9dhQCjc94ZalfZSu+oi1JxQisyYEFccVXYNB5pz8c/O2ucJ
TIvTAqmsEX6x9t0xAebFw2cOLLIQsZmul7GVhUmv3BPyLkRqwR1s+62EvmOa8/HPCeZ7emeVzfYC
dDFBwfV2yLqGrPPcihepS9q6fJMnJweGp7hshl2/vu1sQpO8OSOcgZkuJugmaRVKCPKVQ7PfNykC
cHWisLXbGQAUcxB/oFnOAojWz5rsRaWbsxFhH3s2rc/Wh/wB2LHqjLU6uvln6046KhBQ9RB6SkiE
4bMgd4hrwHSl3qJnUaMB4LsYK3yhabfxZ+8EOBnLKOq4Y7zBklXzxS/VnFXP1A1fn0RenKsMCeae
r/n1h/ceInnKl0qWDQWQRWYLGilHPKkysCU17j4ytLq0e4o0zZ0gbcQe+wuCNk/yImCSfyDNJvxz
gVeEuLPmE6L4TwsEYEWIhK6f2y0FUBE97iAT0jMYRurRuc1wgDn6sb3UfEYRv/3c0Ok1wa7C6Do5
/nLXcnWlnKZjq7lZldi2aWV/qrKma9LbnOGUxvrSwbvYVs2phVoHeN99ql3T/USSKrf05rSSt/UO
ZHCNB3M8gmI9eKWVh9AdjhP5EPnrb4J3y0RUlo5DnplCX1hc4uig0wCW08O65O5jEUQKaUP8KbC4
20I7jrLsIuTN73mWon1pYkj9fTNhuDxCfZpFjTMAQeb73UlgADVoei49Mk4zflMf85Y4PTXmyzcj
luYfoOgbgfLNjAszLImzqC9Tpy/UmSanKSes8dVn3pt3Np9AYRfyl1q5cc0SmwW2rlr5vBGa0kHF
KpyTZK1kX8GS84T4npFWLdypyltfjjGKx0qIZb/DHEgBIMBjpfxNI3ZcrM+axpDYbW2YAdtYBsOJ
M3TfKtp7zlutc140NO1jKAU9WMQQeTFG/UKsKGOXqUrmCWOzzeVgKA1SIN+4ouNegUsLllKO0QCp
oBNe5rwiasWvSXc7+dC7i/sAl3gp/Pj1cnoETDNudeNbDKcJphdlE/8/e6Bww5L4b2cPELaI7jPy
LpddUg+bGf2xTjL43HmO4UgGtm5vm0OtClyi37VchFRTHqkKYwf0ubheWv4zOO75fCKknmITGlwG
mc3Iz8f8wPkedI8pAp/gYvT6R75dpQ76JQE69J96mzBSRz/939qEcABCq0xCYas0Ymd5jWsKY8WW
r5vtfQQDIOZqnlY+38W/Lsv70fa5lyKptlpnKkyzI21xXuiMBEgo4P6tPJe0GLvBOBwoekq8+n3l
K29+/8kjoVPzCCWWQiQNNUAawmIL8rUhWwN0PSei+ufetcl13qviC1h9FCFnRVM+8mT2Q38Z6Ccr
rCovXiepwkfHsZs59CqKN9cB/mpnG5PeG4S9kOUrg9g95VAxLOFFBjbchajDRJEAJM0S2S87Mu/9
/O1YHA93pL/XUiYB75/3/Kqd8Bgxrc5CoPDrgjugPH6W8ELnQZtBFBMI3+JJfODwK5Hb1dqLu0lI
KeQSwBbJRA/b0fCx9jlO1Vzi/EOV9X8PqvFjQhfC54+CCEemnMQIltrJYE8menOpUaGOzml3p8xk
VUpnaBUsZx6PQXsJUsY9ssdr0puuOUC45W7B1FSWzF80UMJUUKR2nigL/dlZ3eZ1Qjc3hnsre2Dh
sZNoMWqDY+FPVyclEMoibGjA2L9ygVtJ740JRirr3dDwf3PLeuhMskI44GBi6iNXsxYozxQYKagH
LjX7agerta2sVUMM7JRNazoErc3VKjN+PLEKl7MrBz2laFPs4zA37oSFFTZU4eTaz14XBDHQcSWO
jEBMCAb7VXdYTdyjVtvYWX0zwTy2/9nAlQuP0SUR2fBQ93mgFFSll17vGrNjDQFHywTulcEV3s95
Ign/DX1p9iBh5XqBXo8X+Q6drhahdLag1sVgNTC1Be1xAE+j+VX5h843EhMNBhUK6qk0pkX0BAkr
RBfnwJoUuqj+MbC0WdancOIJ5Ihs+MxXrMD6pVqyppcph/KihZgM2dEaiTPJQBFQcjdpWIIwMIoc
RidWD8e9jLIpJ3Mz7l3zSzNPYx3oEmJKCYpc9/OU6+YzKrY1EmFKKr/X1EHquW5T7gK5CZOHB3pQ
BxqgZeAe4Bac4d59sdtdWwzcR2KFrnBx6EejFjIgwY28XnseLpjtJ25PM9DVjkLVR/yphdKdumS5
XsbS9cgREHiTO1rhYBcf2dVtizk8v4U6ffiKNLG4j17rlPvQQRGTPcm7u3WC3byBxPY+9c3UHJqf
HKEJP1FfPQuYfRyB65O+CECY5zZdkzzbInNC5J94jPR1PtwiAOQyq/52k1YpAF5EndgZWxkfuHHN
7clspMbERkdQG7vnZulgkjQP8zFBiaEodEx0mmamOQhP3xV1s+nY0Cxcqtt+Uml/lNhF7RgmH4ev
B+qxJ+mn9i+rS38rObxOt+hBELtXn4KRsH1Q7xcGSthOBPvyjO+40v2tCK36I7ZSPvlVgKi5kETt
b79G8nFiUOagXAUUoMrFIuCkD69im+1sQWnMCw808S/jhz3+6abDwqRY4SQpMmfK0imjc1n6sEYN
zsDC4gy4uw8xWLQJB79NJAA2TfUGCBt0ovu3zde46SyzLHS5x2rJeyxFRJq0eEaesfXbT2ugv6Kj
+X3aaBtcpDSroH/rEMwb0+uXY3LTzpD0jID3ADpM7D3B7quKaQJNdQF/vVSimu0MVPdF47GBVDBB
2O10tQFatuHXgTq2zGZkxUnHCH4w1fcGWUlynrKyCLFmDxoTT8ttsVx4U3gJ00AJI24dJoTHzLC1
oK8LNDwArxFxYm97klHsE2v2Cx6jNoauN3Uk0o4prdP24tSMLsENs6A5dlOvBRje/AWF69LHbIiV
A3E/Zji2R/+Q9Ab1sx3YPsz3lNpTVFQkznI4VXFzLd9bwc3zOQaH90QBorstrhfwjcUAYa4pTLLA
KVUJDCLbbk6XCWYkprNJWHxf07UqTMlZS1UElBnT3u1WE70/E4YhEFw8qxkDWdEAzDJa13Mq4hDZ
9UJdCtZ6i/vrPeXYct4j9oI3milWWqWVbFnnjMK2LX6EnfOCegm9VU6ynAXuhFNtmnetgyR5Hq1b
sYeQQVo7B6xpERgj3o0GUVz+KojNb2MxCt5KEjZLdLu2PHeM30CDsP6TBN3EFd4M51aP4E8OCrEN
ZA+LzqkkgHy0mFqMBROo4ba/3fP0dOT+AUDAbRmwhDAHPLbMxD2LvcBhmUOHUIn8T1dnMJCWLxnW
ntGXncctjTp/Vwvbfy7qy2Mxovpq9EDPAC6BluQhAJ/rMWyqPE5O98PWl5IT9IbXbeT9fpfTwwWz
0g8mk56oQyiGKzYiUQVuweX5v/nQw59a2s+gwr/Uh1wTXcIvfAjtFK/7Bq1Hncthx0U2p9P6GLnN
uFJ1I6dwjo21zlKj2oUd92AUklcjI1U98waZ1QxUf4lUQZ0bIi/mdFQoiF1I21H67WEEIVhITqnM
iANxMRFhvaiUzkj6MJgOPQAhLaCwFYbuTsPp/xKLpTCkBuU5bTb1MFuPfHQARqJ7xtHyj5yS9tBD
tKdOYp4pLBm1ifRu8B7OKOMuaszf/R3+jOYN9ffRqPpEiAeH0CUHtD9RRjoUcRnlxk6yH+IK2Bw9
2IzVrzH3a7X1z1LFDEDjmcLe2m8zjk+JQdDJZ/sX71FlgLM09upZRA/JsB9d5+btJEL9KEcr63xJ
pP/rO1/0DnVbcSAGd9QzpAApy71XOIqxB4+Mzyu5WXQxPu/Uy9LL2wmHh7yt6K1kLGLH+iXcbZcj
0cSX1lrfSJBZz6qg9jvlvWjAsOtMKC7zuDKEZrLtLBOxGnLfi0el4tAIyeOf+7449lkjiItN3wva
5xlJ7n/NyFnwiUGmubv6gTKQwUMQX0LHXsgfDsV70wMUDnFkqKLyX2M0IXnOXaLPNDFg1isznRw4
bQhR+qW9+cfGrANzNv0UVi4i9wAD3lUEK76RYRbTot9U1kdHXtHcTrChWmAHbOEWj5zQXKJAZZbo
xTl1/4chm6aRHwZiR7tzyr6VgHjd9pavevJyDbfkFL6HcAgtBycKs3XmrtzdD414sQg5dCaZ3SdF
UZJjfK2j60GcNZP/W2i1SYpHSfcLL0SNTXZL/wHEycbCvT5vx464jDizFkMsZRHJjNDpnFWkj1yy
YI5KW1WR+ADwvqoxmpkDrhScCt+XjWwR1UajbrRSzAxOcJsZ/OQPcU23IViSst+COcBN4+bFW+JU
cRRtTtZkwGLHT05JS4D29OJeO4wnA6zTiaFwN6EsFSXbZvrs6TCRgvC55WfCgYxUCrMqmqEG+LLr
JKyr5btTdvifoKQGMBM9nMQCfhL07xdJOXZf46SUvHvcxbzci6NwGiKZ8CBA7f+FY+VQXKI3OSnI
19Zi7U0X8BN6zBBYBRpZ2zvSO8aJok23dIIntyrzfevi9+xaAzEEvNNiPTu2giMLgY/kt0TQoSj2
+YRZEkk+3VgBtZ9Xj0QSOnR/tTMDv4M7Bm0rRfol1P2xpsNRS5ojsoxpv2jq3wqpT8YzAQm1+xIQ
wG/JS+MBTysiivnc2wC38lKL6fmFcl8kiFpox0fEJrmVHXAiWk9/d00S54Di8feXiJ/l2Wh1zEvK
Vf7H9XYyI1ZVACLqURQeZ5Wz/9gE4iB9/jOIm43mKsRcQ5jjFVt+DLVBPz6yd0NgSuvl/QSjFZfb
FFnCajZVpYb5mLXZSIQShLeXQzFivDpxVFFjTbLmFRV9jznMUMUrc939fyvV+nlTidju1LKEDFk1
yw0EXniFbGwpeRZQYBPefeDEQOHbkJc6JKxcSOv9m5w7TWdiyvHI0q6AzMy6keOShHj7Ur16LJh+
CK5T6x9RZ3fi4BovuJdmWXPjlx9qJGoRchljcilKns6l+UDVY1XB4cFI14PwHo7Jf+RYrhqhYeIh
DFxg57f0Sc+3HcQ4z5NlTFFTtqe4S4cOjMOxU7nwlv8o6g8rDMv35K9uBY7nN/s3AkxBf6FaXu94
T6lbaRxM27+gCZmYfCu12+lDQFjyGhpWINjIjf7DoGHmct8o1ds1zhgBY0KnaG5p7OsSeHinJWSg
YOmBUVSn/BODXuvTO/EaQJKJ0RFiRjtSkasxDvCSaLEZiR0tclBbZR1+8bgjnxhGX224wOloXaJs
2tiVYKmuyqTSv5NyOjr7LAmbSrRD/ktx/L0fVsLYvrX2BiRzIoB5f3l6UfvU9MBSFDPlykv+rdBQ
ucrgeF0pn0W8SCdLmZapvALgTAUN8B6vwmeV8T8a7k7+WRzIOUDdppvS3wqPX1vNf5rNy1Or5tkF
L3X4dDIt//dJSOVLb9SJ4KABaX6K+H4rsdp2GGrECMXSvvXw5tamr+Z6fBYqOJVtKgVRQEOAY4sN
chFb6ePyY7MH0frR0emHCB8b3zGYT1wU1bDGMStHg6V245BHKuhkTC2Z26n/QG2RrrTfnCKfSTnN
8NpT/oYe6bzPARj01puJIczNf9lVjkFh8wQGVkXMSqtsDnvDDAVFjxnVMMlia9tj6MEttZKMSDny
CtewjT1iZGnzm7xEjGUF6+6ObSrymkwlHdeZQnm6TXKVpubpaHXORAo5OSvgd2apuZEfEvXLr01N
cU/XHGFllLEGlGqZnKjpG2MynPLaRyaR4GFPTvKwVv621OUkuRI5GNm1uvet6kgFqs12h/6DQjdp
hV5GnsrTefmeLwVL7s/b2EK9tmT6MtO4Vm0vO8p/3CHhUMTMC2KHokmqxB869UcHnLXng0Dh1luy
oZaXFrdYUj7z/DctiQQPAuKnXabSwVasSk89wjTAafFVI59iJwrbWGr/uJxYqoEMDYTdeQD/eNI3
lpL6Bmh1bKsI03vZP39n1+dlsIbqDDFmimo/OvKwMcl3B8FD52aKTcJrleloB5GRwh40sZ0HEL3B
WwZoeKn3akQyP6HAR2vP4O65F6vg+b8vMey+q/2Y506aR5iLSjDliFjOBVaEUn18FapORHGXs+6f
LotOX8t5YKtklzvmiP2GbEq4Ia/OC+AcFAvYLPp3nzSCFgYalvQYb8905t9NeyVzoIMiUTzIjA9H
eMKTLhN4V2dGTV4G/noEbhn8JuGNUYq8YsPpLmna6n44Cgeajkew+fTPfgFH4Gf/NfEUCc9fcgo8
2RaWUcLCjaXIGiEGlIeWwFhbWyct8VPd0X5vGsapD4kNlTgZ5Jm4RUDKYhilkPkWob0uBXqid4Mn
M0NtUhraasP+bUGviTbFfY8xqeIBtgYK22UAoq1gGK7Lc4scCr9NmzijDmrSLO0wTZ0CMFNVdUEd
AV81XuCUDZA3NTvlWH+6YT1pD07ZPmY8DVhpbmCKFDQj42HfMi2iJdb2ay+DMsojbn9ubVNNe/jK
F/QUlzWhJzSppxBzBgjnI/VKfI8tBajNHLt6HomhFJ/MIuP9D8bkjzx+pJ4HyYKOPY3r5TLHdh1s
JDtMIxEJl8uJ6lWaMDS4TAOG7Bin3KYTnpqnFZBHQ7yh2wD0KS1STzfJScKGEhG3j55orjP+ns4O
TOF0W/LbxPzsTlYeQjtu467y2Zh+CzJNkv+hinXQ0s5YnlHKFaMVfPivLHOHAoi7TDFjZfjvD0+f
avZJYLTqbKfBXfOvI9alsOVEkSV3UGVk6eXMcAvtKCQMp6jhhTSFpraCKTFHZV3pRx5fCDQf+03D
jEr5Ukjlu/aYVZmfwxJhhytlxVKRBFkHgV9hRLopbR1f6XnAlJx3Ceec/m5BQwjbsoXRnJRhpzIk
2j/AoIfbxv772yAA/XUT6uC04QSrNy44mkL4bOA57907HJJX/CS2Itb+wdOx/1t13U2VDCOi+OBe
ftQJLzNwS6pVYpVE85qsAg0cP5VG4JVzJdWh2jk9Oq4sZm1s35Q1eWznw5hha9peS8L7tXY+18qc
MAyQqAISvVUgpjx40xhgpSK6ktTNeq56Mmada6Zp9lXpc6Xlq/TWloN0iTSZARsVyWPYsILQOWBw
OV89dpN4yHa388SYmT2YkR/wWV/RGNxmrJPiLkN4R/n0gclkbMj/qPviNu/F7PZiHpO8oOhik9i9
epIXh9H28iiPkaCxhJUqUKx4VMMyiHVLPwqMci1lWHDBMbpuawol2iYXD+Qp8vnJtsYngeCgRoVt
3ARzeswUrMlDqK0io0ubPjzlWJXgc5wLRIyaV3NCAW8412DAyxzInXHUREaaHiMNrXrW3sEMsocx
2apOVOSoPuhB1bIHX/kXnogI39omNcCuqSXi1Ze2KOpdFyxoAgArBtgJOqf8m8sZ2MAJMvN0BQ5b
0KYh9+okDCcBNcroV9fFLgxM3YefX82YeoU8H0LHWLh85UpgWG+KOdm2j63aD8Edm2Jjuu3BL/GO
m3giV/vYKNq4KvuwEOsqnKKPPETiX+nATuAEor351qj9ePu0olt1v+GVYKNey4LhOhUnOW7MOVKo
w+JVU0yUazvz/ny0Weyh/lzHe50A/X8QYNVSgbZrPeYPGOUhzajmsm/Smdp1PK0CLMNd0vayn19K
Eh6Qatjh8gkprbxzRIURR+AeVDiSBWMJZGsr05GJBmRUTUHGmAxCw0tA/lRShT/a5P8+UrP1K6sI
8neI5U6SJ+jCtMWn8uod6QrNQ05wqw2TWvF/i5uZb0qgMkf+FYOayRZk+cZRyhWJPDXKi+f7YzUj
wuhItbdUMIWPMslYjcJcZpyzxHWV3e8+unaAvrQKIJAsHew0ERNA5E1bBA0tkw2PebTNVLdCEpab
2G3nUP2TEBfz3aTkpa4dCKaijsetPg8kALAoiAK7/DyWOajyGbu1tKyqoU1k7fKRXQ8DpjWn0uLd
RUYjMPrASzuvpQbbOC+OXqP1rTwtXXcwozrZSPNjNtHMHxQMIsLwveMk/DBk1lunC5VDBKmVLJ4d
L6cEVq64oGrVqKYsm2DnP4tRYImEcZZfvwztTMuSEv2vI1AmY588wfyY11L6t4SBZQ8KZeRfzW/7
YBiALfiMEjh183705qnnyivmK+ZLkYO5J/44TpVk6YRyB6AZkfNfrPIIQBfKinP14k8++y340t8+
XBqZH1GJjArcFpXs1mt08tcS53SADM/xluzN8MueYKem09vPcNJU2xGA+24JNmFZlqOHyLbt633W
78G8jrlZogUaYiKUH/3hPhH9Ifp2djFe+vugqyFIoAAuVtUtTPrs2zMTjWeB3ZAzXcc9FtUANP3+
vcJoY1h7u/MLsV8pXsI0DKPMWtzd9BcyhqcANvn9SS2LImLsbvckvvZWHlvH0COC3f/17A91lxMh
giv2ZYr02nS3G/zpaZJREwd5vQ3joNK8+8sH3OujgrKyeRLZaXjJNGm63EIOKlmdDuQItBgcpRpE
nebHkx1BGQAe0TLN6KxM9kK/sU4iaEWCaNHqkln7r8gwVpk3S2DnmQq9IGlw9WjZ5IkenCjHFqGS
6pZhrZ4BMfRsk3JhcYgW40iIMxRHDkP6GYKh3MKff9phQgf4A08z/gyOBdJcqNt/VoVdJ7PvfUHa
1Fuc+losNyjABGvThYUwfrSr4ky9y7cbomOd6q3tDyUK1oneeX/h/7vLxPoNpXRJgYilvi0lhEPV
wlp3Nb6emi1BoMX9zDgXWg6m/Nw8aFU1dtLd7i6qiH1kmL7oSg1WlrH5a2f6s5jDMYekPZMNYOM8
ng9ah32Lsh2V23aTZ//eseuUrdvA5sMnzWMOW7/5dT96wAyC458kEHzznZ4NbivDB7Yx5DycnexJ
PyagQNpXb6qRHquL/FZoTpQCNd0xOGqO5exw6VcqOF+4zr6khi3DFdnDryWvODLMRuOat08hoVze
/x3RayTHKqYawANee1SDuMChSbTi5dgj8ft2lOVi/iw8K1uEAbW/PeRFzsVBd8xo/4NnbW1VPnGk
/fSA6iVrdWXbMrTr892bpMPDN1pTsPsRTpyuED6zQ926r22dlhlXC86dZ4mxLMUyHFegH3Jjs0my
rNHjpDBPTdwdioDGmZbUmSm7ET4ZMXoGFm5MrRlSwD8CgHZrmpbVu10Xv+ynkHQ08DMRHbrjTAax
z/4EhOwWriVY/fg1QfQf61bf3FZZnNMP8e9E/XPcY7X70VmGwmdYQURJAT/JXRBn4ATsveOXUSdF
PMAPumYD0MRVmFVejRCrTeq1BRkXzPipN/OLMACTbaWMwTqH27PedZp1eY40LwORXMfMDOaNdesQ
FWWL56h96C0HjVvZ5BkqFXCHUDch2JhTsd4Ycu8raoUXjh09sDANMDfmYhSCGYQo2VGZq5jjad2r
Ke355JKXOjFAULNv6DtAnGQF1MERtqIA9PWWZbxnPDuD4wpkNgyGLbAPimCzJaIWdBUMao0oOCFE
AV0XxnzmWYhhUxc33LyatbmwZFGIGNHFYrMnMXb8/5UEaf2uYWnSI1aO8r0ikyO96YRtY8hCeinS
0H8SsmPCdPURIiGT8XI0jeJlimL/PUmmH+pKy1bZ1UMxW86eEfi6dl+T8aQypNkeNR4XMAC3ipF+
GF2KK4kjKtk71Hwywj0wsmUoF8k9lrX+0eznX9ZhAnPX4vzCfOZNCpsRiqFQYFwvHNshsG6Q96gZ
i48FaW6ZT1GR5HyppAdl1iy8YJNgv8/Dtrg0hNB8Mhd+zhq2IVjsIEnfh/2C5oNmp5DwDYikY/mi
gJXj9x7gaZ/d90TMilUWIZQCdlknJSaWE1U6ItAYJztBOlnIhUcKc+EJxxZOryDeXyLcDTHxI/b0
b6222SvAoDBmDPDEYKbepLL//hUD+tM6mP/TolUX/U3htduKZim48xhomH7jQJKtN9DTeA58TfCh
yHtqW+3gs3KWVwLN9xGy/Lijct9r6x5he3swmoIhxQEa8QOh/ccvr0/qCuXwUQZzGyLHi4ql1kLl
SoU3WErSiQLOREtXgKFttcYN1jo0JcStpvj42qhSaGaRxlkduh7DjMofSZ2dUZGDKYxXr+8ozAWV
MIDGN8CrNtPqB7kHPz+Z+PSM79rsRIqwjp/dFfF4VjOHoIVgxoOH3GCAlyrBS9RF5Si6PST21KiR
3g3dPsWzbMZoghqcSiYKdJWu5aP/z5I8Pm867YEkTmPLlSkllMBOM9mAEqYO6XRqAYk1VPw8hbSW
sINSTF3gn92NxNmAdxeJTSSby3vNmh2Q53vEvuWvFiRuLKOSd1vjZEGo9YfEgPCH4j4hrj5hKnyn
3KmejD2NwkDpYit4WK360tvklV5NXdVMC4LC5zLD0hZJH7c1xfsIKz/5uSAGrFQuv7twfncoH4Av
/D2tu2jlSCvEmjLiL3FApDKL/+2HLnOePR//Ae1swYl7epA7u3xh8UcN7AgYfu60QvTN8LGqt4m1
pvaH4R7yQ/gh1smRmogNdwVAfREB6J9wv4ABzWcjWHOhAKAolV2rKow+oDnfYNiy7XK5D1s8d/ts
FketoZVXFpbZjOP/9+gyHRWjFBqqNsj+QN+0FEhSSPekDMbxqulAR9TVCgvJCFVuXPazg4uzX9Gc
axs74GcfngLN6aY4zwRt3aOTwdqiY9Kh6ulkJ3soj7SZauqlDHCYEQfunKkmGLDxdLGdRk4AuhtE
goYKbuAStBInL5VikKO3BKvH5AHq3hyhHkIPrLsc3AES+kOwV8VX//wfWNdV4/aqZcHC4FOhJRck
GYZ31PdADAcGweW2Y3wVHmAmxzCG+AvKm/E04dCru3UoGg3ZeawMBetQ9DWL64uFHBDIr+quZToF
XYfqaNy1G7sZ+nw7dp370zu7kurweyhhkSL9RX3C6cNktaf9dyHorG0ZkBYEoNyJ7ahdU6QFwtkJ
Q8insbMSkXobtiHf0pAL+3i6ozycU3FCabE+U5YIwSJLEyhMOhakrU1Mz3DAdBiLj73xwqfdjXpu
PDZc6OYLRBnug4KfBFMueAgCYinwMKKuK7eoxUq/5MCPOHpGnpiupRn7ahFPzNclTObOlM14BTdX
I23fPpDtdIyuF+Ovqph34cBNs7EUi6sTwbctn4Wg+vTDL7H/8nlreB19XhYlcUSW/itLq+8mxsYr
s86KUK6qupsk56y4BAR1FEeFdyzDmbBswNwg6yzS/i127wsuwGLg1jOFjYlAUhNPJv5G4eT7JkRD
0gKfdSW5wN77ICrmPhOphde3MbKW0vQk84NRZpZu/BwwxbgoDUglFGxc29jOTlxjSOy3sO5PnWm9
7hkN6AccYg3XD+PZR0ROMU202W8tr7a3/JZybo2smbW8okvVu7XvJDPlCjfKGG5qiUU/PoUglGBU
n9gTbbQmY4b0r3nWqApsKdryUH4vIg12bdhwOjCgGxDmrFSkoHlN0Dy1tEvQjAVc0DZE1FPlA/6q
O3kNuCsA/oICf5caUT6HkL6Ttgt1oqnbRRyHAtaZQ04dF5hgUow3Jsz2z1oNKgCnaJf4yuOGN+jf
DTKOjlVRuKBrMXWXjTIDNXxIJK2z7HS/h7OoeLUjasj2lNrpHJdcHThUEBHazalc5J9alfELk6bK
uxtXnAScqstjw+aseiU3sbsYCg1K+/A1kNzsfA0nq5nrxrrti0sy9x2+TaCaif9R/SuDgZ8e+Hr0
CPgbOU/l4qeoK59DRzsFBL+SwgOAMuhfiRx4SI9rZa2XFjs9yV3S8dZhnfnLMjNNXtJ25JypvWVn
togGLTNOHGCVLVbIziASsOFEXy/sITSPkQuHutrbrFJxorm0CmJ3o+StCMTe2KVzxe7KBb76zIn7
7cFoTB+/GpbcH5jH/Zfaddfk3OmcaBO1oKAjHupc6RbdONAywhjCLScqDdD409JFUSxW+PuDbOhH
cg3ueLzi4lZ1W9cWEhx36Zo6AqY2MuxezR9VijobFIDbvKa6Z/W5+hpA06j1xqgXGZJ34oeHfl1B
+0yp1QGrsL8urxmm/sHLzKSe2Vihyn7Je7o+qjmmsBa/U7bD/M8GTsFbOHXieJ88B9EEH4eLvIQl
SgXmcEUyxAnmoSmpUBvjHkiDL2SG4+MWrhtXopghS36FJK75xuYBuPQOceOkiZV8MBH3qA3IIPJB
OVaP+vFcu38YQOby8ROZgRRrMNbb4PoARq8UKrTWmr91Sow/Q4kBPlBw2dSfzG0xBD/HQ8IFde78
3RPdm/wrEcRJOVaEtLRzUZCorNCuSff+Q0SyZYA5lCSzhxIGjhwD7YXVKet5yT7b3Bbz07yI/JuF
IeKhkswcqJKT81cN4SgxeU8bwScVi40/8Ctq9ohUyYHH7nQaYyLxOK7fkoVi7sGoYxXPGTDXI7o4
n0eWmWBCS+A40hJ/ofmzF+MYKqUDyJOgKBwmkhjW7a+TV/gczW8y1BTWWpzmiwy4QIyhYXtBanJE
1ki4ngT5vW1VrDm4jQQRxpamrefWUUNKVS6JPKCule2XV2wgPadiVIKvU+OVq3URoAQrz2jdwszg
fyd++vKVKp/xZKrU/EFr9szMqo4WFKZuX2FRTbGm5Vk9y1sj2hrhTP8GNCA9YW9WwdWhvV6hgNMe
pSses3xXSKfOulqUXBrBL+hix0JMrx2hnR7ogTFkwFkcaWD0GpH83opRTeKepX8t5ElG+0HIZwKd
0RE9UF3YiqcJZtEvtJh3tAGaHCoH/LRbnLcg1KY6PwpImGo++qP31xLFF4bX+EXiFoEQ34YINx9g
8U56ASK77jDlh0ZOv7JZr3vcBuuGS+3D38moZurfLFaDplvK0xIAQGBJnF7PyYvvDYCkemPeFP+L
YVF/5c2vftjfuSP4V15RytBNifQxPmsZWb1crJs7knA0GxpuPTvL4ktSoJuha1/eWlF9uk4z+nXS
8Ts+JNU8b9/v1qdSdA+B9UqX5dJNWrQP2QVVQvrchLGdFioalNvXavnlljNlny2cZ25Bzb8bZfjp
wg+Ow07LrdvG2FuyPC9UE9YUvG6A/6nD9kPfgn8wK54bSs3ml5vaYqwKP6smgx7R6TVinogxnDcQ
BHOqsmXsV72uJIHEjII+Z+5zMrNronPl6VmeZufIN1BFzdKQukjHAXN4UvDLN0F48EhIY8H9oi8J
LiNXpwzYq0hinITtCUFAkuTGjHKAqtlo0knBdNp860EUvcGf7w849gXLxwU/wKilCcF13HxWAtWD
iP/wyThQaDMvBIh4ZhVIT/iTUdEWybDtr9qrJNBUjgZeo47w17L7xdztEdKNdQRS+v7CmV3s5Jh4
QqvwYONOvqYZ32afp38lkh3FXIdDxjj53PPjgvucZXKHGUq3X+ZM6CvnfNhFZ2Ev/bHe7Jl9FcZ8
Xi3wu+zUP9ss2/TwG0BDcfjth7HKC65pB/03JYR13sXXVX1UQ0Z1aSxwYKJwaIdBIKV4LYf41E2g
a4rKqv5rBC42eNJalteZrGpuo1pVGf6f1q3SILjV2EnxrIGAxj97l40m/Slu1AQPQCJXWA2MytTD
fAm91ckZPZIhLRH4etLhxqdc7FLyZqk5vrUd3/BnrEh4jpOBbBHD8DFABG4xIq7Odn4G6RYLRbU1
XbDylv7hm1H2e9Lk4n4AgpZrZX9YuQtclcnwt9wG5LkoIRfEMU+bA3uIIHZghcW3HivvO2nY5KIT
WMqgLBfoj8PMjU7AT2VX2Sq9oYAHSckfVaaH+rBOAChOyIoVlbOwVDGoyItXwn1KG/gamV8eCwG8
pR+1wdNJ66b8+6jGaRB9UeCY6ewoMuSXICJtnePlL3KehFvYtW9o6kgYAJqY8ZfUEFcnomblEdyD
8krLEVFhC1AGf1mOCxGfMrYB2Ag1S0cUEps+aexOPNu5BZD7bcvl7HwBVfjPJcXIHTwVgmRyx9nd
65m4brz9CT8uSQ93SlM6m2UtQwp6O1vDc9Kn2g13ULPfQXvQKJ3/5Wx8OFhwW4/ay2LHGM/VUoV4
Ft0nri4x9JEW5WnqIByFGCqKZtbicKnyHVbNaxf49SlSEtZTd/XENPHtNfW7YS0UCcAEnZ+cSblA
vgZtm7BUc8kHHCTRGQ3Lgo1UhWhsKarXuVZp5RB5bHS5W9a+SwwXRmGAUiIbEJVtA/q0FUC7kKNP
HdOd2+FJCkjekY/Xv7evv16FQqo5+ORauk98nIaR+DZI13NCRLv8QJA4q98rtunDfwdMzk3iftQU
skmLGjshMh7IrFaqxC6BFtBP6J54H+BVDZt60JDMUaReP5REoW+lQJgl6+GSXGzvzgH8cBX1BI7U
w78WZ2CiauZreBuZeR2SvtnDULmE5Nl3fRHf5Qc4pK4r3use9/Na8iKGadIr7vDZoNakis/yjMFU
zvQkuwKp6NXYpMPB78ON2Ss7YVzt1TrAkUGVSmlARQLAVxyTg89Jnw0d34hejr5e8++c3CsSDjRJ
dr7EX41YvCJEGBsqo2gRf0vaqegjJfM/ACSObDeIovqecWkn5BcuYbRTMQ+1HT0SJyidjR/skBhv
2rV2f5wDpF0zQlm+SXiCcg3b3JtoYdt5NOdZJaiiFmRwZoMRs/Qq4ESQQLU6JW8OuNt463QMQS+k
xQoEajSwSGptbzuz5ci5WlW5iDSj+tqmeBhadcCoDM6r/KbLA/y2mPYaZ4iZVHgQMd+DRvsjA0rx
ZvuuazWMsZ9VOBit+xj0iluOijmDKzUQ79KLtXxj+d9ffXXKDL22fHvMMr0SedFxqPVGhlxGjwxb
ltuhJ1+M6GHUoWbQ7hCDlWFJzp+hbblVPdmZ3aRkVNDIEC/+p1CL5TJAjMcHI5ed4X7mF+YUE/o/
K93oaenqvxh4tpCBa/rXHl2G846g34cphnE8BdtsOorkiKaCTVUbYF4XLJOL+QxOKQlQCjvYoVYB
0Uy9wd8N8etG/Udn9EW7ZSClOutbGF6JaSx9fzLuA9eKkyDhMN1rq87RgKWcIWPffmG92istRykC
rzUC1O6k1xdMPONTTDlp10w7XB7ZAPfkHQNt1tJKjxClK3VRHaiR7w5lEa0YaWuzUaKGEswvrHll
yr3xc+H8rXHiMnLo9hEzTkTr0JCJ14UTuUjx2Pt6y/HmV7TeWxVUHwzJvjgYdp/r17sBF2AQjgT5
IpuSUadUAcbz5HSrixb9wCj6zptWOwq+3e7CzhjlgNuPEM0d8sY+ovc339Uizt73U8qGE9RJWkgy
1+TPWam+elKX2IFLRqvh7dbnLv53YKg7oCSB+N9E5ytk6r3iKV+5vLdkI3BcSqEjFwd4T2wFzkNR
/SPP+9Hc2WXbWyYboraeUf5zcWbsg1ntpjB4pPRRLPtapGepigNoHphSgE6Hkif/EO+4BQdERLr/
MI5jvJFdMFDHWpy/ymUW8KoHv4K6PY4HGQeRy17qUBUW8lCMCnuz+7H1hrWf4OSKqc2Vz89EAiaT
6RF0b1jru6oL0V3Tpi5EBQRJnD1HIhfl5Z/dW0ERS0DQf4o8h/pyGJfT1loa9Rebc/7M5qVvhkNp
bFPiQXMF85XhaAHXuvzKFLOIzdS0zL0aDlJc1KroEO3DC1CS84KtoiBNOGFnRMsz1gq/d/DjztIl
gvStpUiPFYSwJmKfqD6+ftKC1E3AUkrdbcSa2WaYydRSmOrL9MaVIgs8BZVbmH7xWO1FiqPt3+/a
YGOQxk+aWzYcPsccjpdJ0kazl8n033QXzk2dSPBTIkVNpG72j+rcStR755RWS7J+04jyC/sD9DWc
d0AI88AAgybksVgDSWWTYeMCeAz6NimiZWqYsKHVjg2ZWOJ+HvIEWFI5YZUVo8OTfYkGLOsbEyXA
nTbl0ETq5syLQnUlQ4lWtkeRXRtZBaRVHMFj2NFiijt3aPFHfFYo6bVLaY70wCJv9pLGyuK9TwM6
H8kujUsuNgq8rf1XR6BAvP1JSzBhjarJHJecnzNoK578sB5Yp4qKje37Cm64JRdYqzeM+hnB7jrU
NewMf6w49qNNxidWaBIH2PHBjUgc2fVLpGLCfO7YBYvjUJdWzHIH8vJpQfekExxdai4tcykphjkT
y4W2pQcHpqoW1Rl+PoPcKOPI1fIRuAvR4E6XR847ZGE2W58P1p+pAEhyJRnhjUVS1UQhYSZ+KGyX
k1JKKpttqY982YETdGsq85QisP5X0oTBLqeyPP1imef9VHnvW7GG4xYDIGCAMyz8uxeyjPIHgBK2
ASC8UbU5NM+An9o6heYSplb718KLbaBrUnNQIYoWTNeVdEVuOTTEjGZdHldR94Y+vlmNkHaxFOeh
VilEOcZaMeFkG7RcbhvOPL4neeuyh/I2P2EXp8LpA6HLEkeoBAl55HKf3xJup4/14XfUpfvSNnXT
ZAKza6adbJxjjZmfYUBTEkfYZHkKAwwREitgmNvazDc3CiEr1SlANiokf/i0pkW9+2epqhV2UJ/M
P4hQUn/Y+xz4u95Ndr0fuGfpnp/bdvYcEEckVtMRquPS1bdV+WAxt8kaK17z0AiLFRiIBnjrsBL8
eXNX0fQub77wFvtMCzAkqU0Dz545fhmNvsCIEtx6wIe+7d7quBz8lt2mqyDtB+vM3V3+Wx1p/Lqu
vmAf5z009vGDKkFc/g+ygvYmFr122pBR4+gdvBYM7pZemLN4mKP1ycl+grQRHXz1u6AJx6A7q+c/
q/b0Wi0EU/MeBuR/X1DmtZYhb8IPlvZNWc1tIQn4cb2702VQxZDw5jIhtvSmFnJfjsN6OZ18lVjG
/0mSTClJo0G/la1W8AtnEAQGTedRpbb44Cp6IiHSfrHrgWoWO2gd45lDyQ8Q08VLGBb9OaWoXQ4d
6OHijkBK5F8M4okHIsKjNxIVlcOzmRtmhy5bKxdRkkLzvlfAtK9vEAMHP13qq6VQdwRQOqSpI51A
tcjD2V8UqzfWC2YYuk1ItR8rXNQ8RYjYp6sgX1qg44x9kfckrBxkR/+EIdtR6rkecej55/P0eAaa
55euAv8/T5poi88z3PNz9VZIHR2ucjDr1qg+wjKhLq0PPqB8qgJtocD7X1NIL/yJayobL3/Tumz6
R9dp+uVmw2zG/plSXOVjoiBab30yOJWw5HZsa1yiVRrBmt2xqeDKmVRYfR1pYVlCxIm0XKRLMjP4
44GJqv7mgwAzEGCn+K4hyzTgnipYHTI5sZ0tUAYC50LC49MC+yRMP6CLow8x8FspfWqKnDzf1aDa
bivM168fIGsOt6q0sv5v0CwvQ5bLxV9KkrUcMoVrGdmSIQheWfiRp2sCf/fdxboiFG4h3zsFuBwi
Z7SHatl4kYR4S88xYZCGCpj+FGpQsaw+FgYA5Kc7ewrVBjedJOg0mlmRGy9s51eJPj23RQmXHDV1
9o8VCLL5oTQg+wHFoF21DT/atxqcSRfQdvSCuEoOohBhPu31SoRcdvb7TbqLa0y7QS77xZb3jnwL
UrQAZzdVIm5Bt9wTsnq5RAk1CWtQpXSl+2n45b9u7PJ0SfiAzbCYbKrP+Hav3tMOcQFJGPLYId46
THrqxBXnUkPPFYggVuivSPuY1QqWUw3qcdnzIIh91pSIxOp8qpmeBoAovex6xi0lK+8G9VMH3MXi
G5Emlq0T5fSs/3RDv5yT1LnUFUq4smcW1BqcGlwa3hGij/TrOMdEEC3mCxvP2hafaZ/If+RjV93R
84OT5eIcqCmSkLOlyakVr5mYCoWcC1H7czM56tc9b/fScICCu7EV3J2BuoUXkdp4SR1wHKBnPozb
8O8ZwCS/S1/cSnfKhMZ3oDcWKvEOFPPW//9dKHcNk6HSGHTqCu6iDAlzBsk9rK4cBRU/JBmHNStb
oyFAm/p/lENeQlSTt1TwAOCrDkAhS421kiPSAqFSyXC7xnrJ0J+IoGbusVxjZVO8qsUKUyAhYxbd
+UB3q3/EZylLTXOqZTqkbkhhO9DNLYiYJRIpnvOG/KEqVVXOrKJwr9w5Uye4+0qvo81skji6Kyyk
USGj4ActLC63ZL44CrJJmeTqimAr1aNJDbocplq2Mqd/jgp9p+9mxHarwpOrbMa8US7gPvJZsQQy
i2sQnD/ksadWaaFXgPbxhV5FjfRKY7ehvP9dwz61YpdDyWU051+WnBSuko5LiOgw9Y7WMI6akV30
uy8ZNWVOY1i9rgjOmUddfhw3VYxZK2I/3/0wrULfjGsZ7FWgKrXVp3KFFKgwjTXpBoTZRQgsolkK
dRB6CDWEsVjgXen3YMv14vMMjL8GfSszp6tDEJPuaNy7h9tWZC5370e4D8SQLanUnfcXOIBNMY2b
ElYQFX0nOHfwoI2jv0OV2TLK87T1pIr4Gu8Aza5geFZz1BFSrfHDp6kGcAeM9fLIh5b+CW4CkVUO
wh8dsAeraxOPdJwK2fTpNNVxGs7mv8qfYPSShyPjklw/FtYwYUWaN9CysCrpTvEh5WZziQQbFhCc
Rgg4LXauEFiy3NU/Df7LXzrB8UTXHa83/3gTSvkr43tZkW4JSZbML+O9xwT+BmMXq3ZeePQGlIsD
IYo9Uk5n3Ka5MfjeigC2lJxdw1THA4e3hOf12lgyHd9iLFM1ORh4+1u5fHzb3KWUf4W7H0HWuvHH
gHWIhub1kHavaJ9euxoPohAiigFcLV5QrPnafmV8eDc3O+B4vgphMhNH7IbEGRDHkJrUB4mzv5f7
t+fc8WQzJv1PkxkkWoflcpBk1ua2kakgChAegfBKLbwj9EVcwpE2TdQEEISf8kLtH+k9Fi1FhUfU
8fNY8RdVcE2SQtQ0f/ySOBE4PxsU28CjUiwkOp9ixtJQhSeyH+JRNvFjQjd9HLktxrXg/KhY7mpM
sgpVlcMO420Ub1yWoBi0EMF4tiPoZa88Jw0GdAqD8Ebi9+8TojDugOdvXik0gUkSXVU92b8RXBdV
72oy3DI6lQWSfy8LyKCcof9ipzGI/lWD7sJ3tdT/muU4YbfMAaSV7v6rEVWRKHoSCJcGFDzkrZ2f
arFrCU0ZNB1khO9M7Cx3qgpWbqgs5r+eg0vBLnlQsUUwY/aPLBMAr0xqPLOPQTc/Y/yL2TLvT8Is
01YvBIK6F8sF+kyQII60rpOvEYcEd622vE5lBTtgx93/r2N3IdyBEUXyeo8VpE2ADsL1SnTyc6cL
3JCB9x3ys7alGEa2mHdIDmzcOVL/1E42mmqHd11h6AJUBwCbIPqx1/xOHZznvm6DNGVr093uqUGX
xtCbBulT0jVpa/nRUNoOxTzxKeUEt6j+dqZGkXSL3i0NBIKjL9E9WKoU7MMGk7AdJLxu/cutX1gd
dD92zzalSJvwtEnikF2sg4POFYP3pt7yfLzGrAc3bsUtREkEM53nzX2+s4nSSvBStcQXXrgchLm3
e+hDfIODFO+RdmuBMPqAUqbuG7un4yoOBR3IRvsMh3Wb5s7Rp0Vn0CTgr606xpkGF9nkhKBdsCr/
c614CKR8WuX6SZe7uiptm6IVqk2MaIvuOQfZkMH7RZ/nNxovgPEbLcnclmnG6+e0mEYKnmkb9lKw
syk6UUGkquiGqhu07SIS/Ko19dsAETboOhlDD3QftSE8qcVLbkhAmhTQTORuhYlZfHs31ggkO5oo
8G4n8B6uVzglxgDhQHi1vwiV38MIUkH/L0HFqowdI1RdSlE97YiD1nZbXzIWp1Q0lAM0L0hjRseA
RBUJRtt0Hjbp0gWHjGsQJIPNVphN+me2djSGtXlESjjXK62+AbjO1EcwYmFFSMC0QcqTuq2QQU2a
nmZwgunteOw+OPE756aiCG8w5TTvOTKz/T0nGox0+Zp0vMXQ1YPDjBXZeE4qa9NoDa5f3ZK8k/H7
fdhgCNT2NP6NIa8TjK4pNS1iQ8ywE9F+u0K6/VlLfEjUYGWNyqSMioeb8zZl17rDfeG9TfrmHyyN
1/cCxQzP91uxhAz2m9g2A75FmCZDRZq8CBf1uHGJ67ae8MVZohjGtRu9PCHfMBKD3ukZ3C/NYWy/
nzHOdhpOvByX0E4DIGDOB+vmb145ybb3zsz04zCLrsRHiYdhwaY3PX5CAH5HIti4h50/z2xQ41Kt
Ku1kebbIxtv04Pp+EJaZ6liinUn/+zOqf6JtYCpG62uqgu+wh2SfI3hFcHQMJMttGgusjzD01UtK
xr5ZDQKMNvsWdjESxXfp5IuAr6HCQQAp7PFJQLkxoSKdX21nrZteITWe+3s8z9BB0BG3v7TR904o
Rj2F84uEXP3txkVkGItzUT9Rtz0XQXUTnZI/L+q/LhdkGaHi9SaY40LPg708XOVi+tEKN0GZnw5R
uWoeq7rSbJrnDRKju/a4nSiu2MYDypouVQpZuH2bDAZ5PQ62GYwYWUYbGKKx5M9rPVwEaF+qjFu3
DQAyDssUBH/YJBzje6JrR2jntMeQVNx4wZk/YEE+Hq1Da55i/ep7nEPHqhDdEwouRTqpBlnBPIJP
5ik5clwGcLl3Myvw7/7w0uK9+7ng4JmOWhrwrGqNxR7g6W2nvmEJ1WSMl+2x2TISU4cLMzz0RW4Q
GeLnhOYCblE1FRfg7So1YXz8QdfRayOZGkO+MPiyN3bdptyXMeAuLA3IrE26lCLHunrUBBNcLhy8
BUv955HUVZf0F6VVyECYofOXbaOwkoOCAl90h3B6deBdyDWGyPXyTY5p+8oYuSFkQQX9nRgxBTAp
dzrxJzXmkIZJ3BsryMn5xDSZLBbtj5I76c1/6i+aK/fkm49qkL2H8FPxSBqal3I8j+VslRIJhX5k
fWjyWUfnH8biICA32r0BxIIzg+de4HXmCkj0KWH8v2qkG0wZQznmf1h+xcrhmPskL5AZdlfuGsSM
LPoBTFhxQOD95SieSYdEgMatzVidH7YWNi+ztdT4dYIngCaefjMFBNoYA+1ysEN5YoLQtMvyCAcY
y+RU8sDsz+48Wbb4QBj/hGKlbSkGbSgzovGQsGgrLTyn9jAuX61rrFYg/5K2epfVpycls5u5rDGv
3ec7T+OaGRbgFct90jtQpfMs9zNPJEiPasvlu57gd3ejjIvfKKWZ/0KJX0N1aOggNwrPKwfWoA8O
fTOGO57JOmetNPpW293UryFptk3fO7MlV6qffS8y4vKZDk6i72Y1m2aQfMWFq96ECdl8mZ8kU0HL
EI73ACzg5qyAvS1Jld6xNGH7cB7NeeXG5qlI0mpnTW6Y5i8N2zUzDZGFShNSe2plJy57RoBP4RCl
VSVG9zu+LdP+tSGZNQaMf2QR0mHHuGXc6zoCVHDyBt9a9aXgIgS2TUXWfSgsvAytAOThnJy6KCWf
eYX/Kxii2nJp0lpmT2I/0ej7/DD9CL7VoQ0XbPkx0GVIpoSPGRpl69FXaAJn1gvD+ZUDHumywA6X
RMqjmaangWHFMkWK4kuNyzVu3TZ6kHfpKPqYoICwndR4pTQXAjXDFmaKznHPVFa3J63CJkFv7CdZ
MNcsxQlK54lUSbFPEChyha5SYv2fB+kmYVBpxQuxeZS0AB7wEfqhdiLrAfDpeZ7W5jQpmbz9/c45
8H0oyWHgg7dDDT51BQnJs/rU+H4c76lQ5U8ajCDjp7/AbY5yCaq1ISqQSiadfaO6xvegWncmcMaB
i1OrLhyORP7LBNU6QfePEkbq6gkujsAOYvS4pajSs1wi/wJL/njRlQSUg9b2aV89nk6K2O4UU0uZ
Dkm9oltUmg6ZxjvcgL3ZHjP+0EMbXYiIsSnFsnW+iqRMPKiNf0Vf4L6KagvGTmABTCFoV8zEHXa5
UVTUEGcKrK7ucIyYSEABrDcNeCIMLPMu37PVdhbpDMJhJArRGctzKoF1VsNvpDqlSVN3RxnHiERk
AivFixwiFJXy7UOQy5D/KToaS9iMdhBSjtd3ElPNO/jztIKYA1UHLKgXxKSqGZ/qJDYdUgaKZ83V
tCEUa11maoAz6rcXY5hpcNk9lgOIIAe6gRz5nzH4yUIrD4zZfqpkXHj2/we33bj4CyLhGkQsPjZb
Pb7B0020wRBgIZBvJzYR29ycl7ZnhWSFoSRagOJguixwSXR019GGsfwQKYDGYnthMXsuDIViRzmE
3zyl/6V/N4De2dPiJxVlEljRGgkJUnoLbxeec5OKGe5BQi56jTR7cmbWudJWwjnP7QT7ShXxDVyC
g4Vwl9CatZL1yleLlEK7+7BqiKZ3fCSAcxBCTXpDTIHzqrcSRzjgEz2KQ0Bi459bF3vOoD88QtnE
akSi+Xvhy1KrkXCkHhJHqp3JlZlHmscLWSHEU7xbzCwAlo53MIsG+c/Iz7JZRSs8WQtHqtH1OLLd
qbKLU8vxQwiX92DIt/pwym+PLBSIQimlF03kPQMLGB7B5R+3aupUaWHKAFCBf4QZOJx7ZapcDV2Z
pvGzCtiqvbmb8JH4JOp1iUvVli1fbYkskqg4TMgQZkiR1sUyswSn7j6FapjawR2Rx6bxanES+bsj
Ib2AXFp+5dUe+ExR0yhjtQd0X4VnhHASm2HnUTIA1gPXz4OsEXlSMLCrnovUPu7PvWLz4tjFRfNP
BFXlFoqyKcG3pWeKvw4Lq2OMH+IxDnmytGaxhCSTt9ugvtXH6yxqqw5dborE7fHN0x9+/hik5Fqz
RxvP8LciilCbZbkfCzRo5/XJTsdqS+Ds/Yz60AH94bCNa9dO+DBxuLbRcctSBMkJrGny2RX0pTxr
1cfGIB4pKqzqIaIQRohx+Qcodp0qVIGlW30IbT3vmAJrnqjJE8i6UCUJVJdQ8qUBuVIupY0rEJnq
xOSHxxfmGrOFm04YH3DwcH2PN5S09d0YK72mKk04KwLo8MW1FcYk2D6IDaLtIiDEQEMIaYJOGEmf
9vwBvZAAZMJA5PN0bbSqm5N+youd8xqfjg5GjxRGKwQGjD5/XPjvqZ7R54RE2M+/mQXCOUu8e9MD
adXGoBuqGKu5/r5z/BO8+R3Bw6gpQ9c3pqRNXTRQIUhjdlZcpslh+Q3IYrmPcQcVRRUnWE2sKYuX
Ghrr91UrSc49V4Qh2mnjsFpCsXyGoYoEIo8GPPmk9CEOa0rUcB4fJuNRAaM2x2THzcK0vfs+qeBn
yQyJoWpAZVRw+zkimBiuzRC/TzDXjm3t7gLlEnzWWvkJdDFxUIERnG4Z5Nb16+mANHo5V9/kNA3m
NjlO9BC9Crhz+GP0O6i/jm4gVTdXMo8vWuHr/FHC4Aldqb9wHGg9g9tuiGlFJ2cVsIbfVIl1VbLF
xcHgHt5ZNeTrd1xy5HoPZQE5rHdK3uDmk8Sx7PlYJU9vINZ1yKlbrqv/vUZO1QipHLqeaXNk+FFz
5JkPUZy7Y5HPpVEc4RfTFyINQZwf7GFh1XbcMPvBAfzd6CCdcVOAYPqRwmdO/o3vNXLFGmeL3+RN
QzyEN0qY0EsUhPrQAQMJdQjCSvTrXkjcpLH3wJYtc2jHraGZ8RgsYDB94NKIpR5z+UVfDQ00popZ
4mbkA2b7QM4Q7FCdV1Oxri6c3IBqSgPHHhxNPOpbFdYHI6KL0HubqVw37DZvRHZA8rcgWxYhj4dI
AvmhDzq6kSplGoBI3/hJVyhJhT3FLOEHUkP9iV6r7A4ha2cAqLwILODXAmuZJRy2Pul2c8SMMTZP
LtwIy3WwcxoLGePfnfsaNtGdmTIjarTD138OrHmnImO0cRW2wFKQ8dv8I8aJqNp8gCbmImIAIaRg
KwIUkNpyhYV4VtSFcB49DNyag3jZdgy6V95vcgg3/3UgvueC15RjxGei7bVZWAj7wv9pMI67JzHx
Vki6SKlUWMTsLFj6BAuaT9XykkEJZfoH0Kh78mJtte0MfNEubdYDYuuuRQd/X+VGEtI1gjKHJTgw
2rgSiRa30yMFEfLhmZB2HO4Ctt7daW7BxNy13r7TNLbPgZxLKcdxRfNPX9lE+Qtp39CktHXex+9q
XMslj0aBmRXRTai9LkhHFd0T6WRoU6ZRgNpszyW3kvpO4SpKwXiHbup27l5ACISCQhiuG+Awaanv
6UoKHyAmEKUA2lO4gljtJxJSZbJO45539PYn2rWm7b+NPxu7XDIvwzWRfoT11caVLPXFV0RPrxf5
/4l0q/H7vVUtqPaUDapgE7M7ZTEK3Tw3IeRLzh1Y5FUhgxdSAvTdYEWmt5wAQaa2/mp15Bkc7qVP
SJDixz2A7x7xdKWjMjl4KRgqJCT3thJ8DSE0ZzbpSVZBXprAHqu1LdbIiTdFTyH1d8dgB7xi0SuR
jBQEPLSZ6rN2wCbpJsjZexyf+YVUN5stnv7dGMLYu8bea0sMT8kkrxmq97fo4MH+fRoC4KOoau9C
enPj0jx6lhHs6TZG2JeukKH2pO+xsoJePWaExyIJ/IOpm+fgJpmYVqbnV+C9mS0+x5hIV+GeGwVz
WpGcTeyGUdjpMvQ8EIvu7XqsK2oLhtuYGrIqpChzNNy7r0Bwu6E34dLn+B6+oiyGGIgPYvQqZRNr
WeFRwEjxEMlv7Lfphq9FVNcRpwqv4hohxpG1JaNbnweC/Pw7MrlXg9opo4aMKAg3tdpUIo0SmRDc
VKiMhmjqjRMRoAa+volSSm0URtW/XELpxld3oK9nnrOLhmKXjD+vYn3511f/Af7tB5PktiPaKC/7
fYDvBpl89+bUyZkGHG4Mf7AYfkDxow8Ykm4ldA0ww4NNP2+f7NpNhbPpordmI8qjfgyrQ7L31HfR
CjaAaPe6VGrbHxYlk13AG+WT5+rYXjcLTFYxiHXsBvAtKwFV6AYkp5VCk/FbmyNG1RO6716upFBz
Rff7hmXJxHXTtz9R7wRHB8KkPM08/JhXjjSdFizgcW39m2bATLryaRy+uNllntNGqcRpSij6R3a+
mWlx4Chmvyv+drmu87DHvqS/QLSa9qUDCumzPzgEeercMNn4moL6Irp4XXallmkQNA6zAt/9hVuX
qGb/cbfw2vbnCtWCO9i9pvThOJYerO97SLAkgRVAX7LWWbvAzyUYQMLj9IYr22TipA4TKuE+kTgK
uOkCG9F81iltZJ6Sj+umuGpHO97PaUFDJvwmcX3CpzajN5rPXLqpz7YZsrnZkbnFLlPTHdDDfIrQ
qa+KOxgkH6dbJanz6eX3w1bWx367yYJLCtc6BK1yWn7lNuoCxKEVD4t73v2qiRZLnpotSNPv47L0
28XNfKHyzq1Eq48vgQXLo5ZaiZ56vY31/sYmWxL8tMSlXzge1n2J4xQn5qa0G/mhIhLvS5ZI74sZ
KdQe+i2D4iRL9lDGUoqb/ws884s0DMhgnB/C3TUVlrmMixzIJcswI8KIXf87bplCF7HTwPq9J9Dv
HsUpKWfB5dNhSCSpCNGWu6rI/GzU1v4O78rITUC99BWXa4XU0xkgZAaXYxwRQEiveaFq3sdcx8tZ
5X5nv1O1o8Yaprl1wh0BLYzaJ05m2XxXz+LUNQpE7bPK8VVklw9ebknhtN3jvw7lkKL1nRQiF2mj
IN46XqJKdDOW0yxzvwYFLsqORYHwt2Pkli8scUqBiYzpXs9FOw2N2elPi8fG9ZQ+pkhhJsDN33fW
6mMIieD+uMel1CbwZjMPAFBHiBuzwyweZwmZSy00Tw6zsQgoC5fTUIeVOPr/ca/hEwUIp+fy44MO
lTJvs/R+v9hmHBTnYgHArtUaSUrAWOaBghRjs9bnPy7chynBhXf8pOT0iYDQ09DKokj1Q2lgH8sr
W6D76/DN+kInb48Ix8x4QEPRYj3Y5GV/WB1wKRr1ojQg9ZHjXptqd0f1Gn/JqM3UQF8y3fLn401T
0Zqzg7iqrM1gKAcaOmItOtwVob6OBK8BVbt5hIN7cJB5bCt7fIcVL2HSLwY/KXVnE6vsmNQov2zj
XAseZLTmp14lDY0O9oXiNS3vJhaZtsjlcPg6xqPt0D1Nft42gdGotLxF6eNQHKvmhGZUKlT+smzh
YgukpoJgpb7UZeYMg3XMvzY5m553Ejzys+F7cufpDXq6/XW6tucYpmH6LG6jVkz436xljSNvl1kk
TIteh//9ZhhfOFOiLs0CfiF2aAs4CEiawyo7mUO7fQzraZNJyVKD0KfOj2355/Vq95Gvoi5IzrSQ
FoaPpr+hbSKW1+X9qs33waKUCVv+yRAeU417jiQCj0Ynn9TX5cy4GZ58Tkzt2jpmRV81tSTu7Fna
yHJEYh71W4HiijRo8QnyF9BnB3h31a9LANxnt0kELGMoPdkKA/XhNWvJEzP5Go3qRFybSKwMrPkW
thvPermC0aboF6B4v0rR1XwZLTHoWKsXLSxaqnuH0LqZleFxmnU0MdemWtE24I/EbshTvM4uIbAV
cEwOT9WFLnKUOwBYJgwZyTCslC4WizmC3Y7YEEWGbiSD9l+i8w2yEohoIhlW8+1i23YHUjqPOuIC
Udg1LaiAVltAIQfW4jUJluETp0qAtWBwTQTKg4X5EFOuk0cI2uwLKZ8DzFfrdBdju4qle9r7uxxI
EZ9kr4bBbrNMKLctrme8KgxgqT2VrlS68FRPgdmTyGwA0Cxd7RvHZle+6GWYpGGhsmqmfMslXL9W
qiEWQ7s/YX2HVI1jZlP/nJ+SpgZKuN9/+fOL5EAZmj4XZq5w7M80q87HMzFTBOkpNTetlRL2DAl5
mvSgY5vvLS6Nm3EqwAuEyVue1dBNGwHxcmGfOAKcYePP6/hEsz7+H8yBH7A4C6PYGNQq6kOqAUIm
pmR9w0ezfvZbzibfjLS2rz/9cU82N9DB9EjM3Gdm0aeN8roHFhFUzpebfq5Z1Es3adp00jliRs7a
OEc6kazwlW+e5eodGejwLU64/sg7LFYSezP5jJkaOw31kToE3+Bz/VPjKTswHeojH9AArX0hm/QA
eMZbhJGlGBl62RKYtB2dHZjS80RmiH1EPv3IuayfyiPE/xKjFjGJ5tqh3jO2Y1ZEbtp/MkjBGmRP
4OuuI6VlsSTU9TnQiVZn5SFFmlxEWzamXPkoBJ7GKdWUps5UN+UW9dYy9cpy01Gs80t9pg+arsi1
9leCzdkeuUCbXbHBTI6K4mJlJOi/WGeI9rnPaQSMqwPJbebm2Uxiov6/OP0ZNsc12x8ymqgGgYHe
ZWh+vrB9//PpCFiZpKPNRJVQXhf9vXyvdv39LaxB73nEowEvubtNPIfvuG/mM6Gyx8G2OeLLGD97
gXWuxHv4QxNjeu10nO4VKWVxv6d5PfzkjEQkZn94bYSa2LpH8fJUei+Mq2PoXRVxD3EWDvnwRKNe
w3mNsocKPqYO3QT4BgoDb16GI4fg+y44J8hX2OwJZh+2aKNMmdElxqFMB0Bx+kDEM6zdou6R2uUF
+LYQxEAKbx/4Tnkr/San61XPgDFiDddbIzTf2e5PP1fx9U7TgqyGAOBl2O+q1YOVuZALXHttQ3U6
y+WfKC8S/tjYw8FA+WkfbDDxFK9kNmKZUwavYGnx4uWvLz55ByTDdlOvpI2adRLDzMWC+7jAq8BL
tPkve3A/pVgshs4lP1k8LUYn54wtOdwA9d32cCJ/U5BwDsHukYmUN/CNSAlGXvuNqhcAzu6SoXuQ
7JH2f7KHxcJb0SeFiiUYDceRKx8VMEowfC5V3V+DJnzME0W8p/csulxq1mEOtuZzCiyUKz4w2MWA
oLUM5eUveJ8LBe93mI1u7uBI66bVLxCRFeIc7HI63MhECqhTkjsEQCAXMf+ZIrmUPt2ELaZcPVY9
J5sW2YHRY11dzK1yF2T4I8DD2ziz6LYf0jIKkL80G8AWSOXlU5opQGcfd1NZNFCsNxkptQESso/q
D5bo7wdhZKntL5DLCIgynjFe/+wNVFEqaw6C02Tg0k9DqGg9sTDAHFnMAvplvCGxCJenAfiKyjYX
Hec1IjG23R9zSO9bJtaJX6XmGvEJ//YGuojzuMKfjwtGFH44ZaR+LO1RgQBFedJHdzWzRd9+Jy5X
4dJMbbWXPtivWVRRDTOPU9AZJd7HnPvqal+wmD8kjbMWeZondLg3ArpaO2hqaBZiE6sonxfkwP9Z
HIGnmgvI10P4O8FoIUlKeQai7kntHiwmDS+17bF8Bk1XLsxl9nrnhAYXKVK9Wx+2r4GEraoPI4Nu
1/zcCcKEsynVvlWOEfINFENwnl0DtMDHssDpG14CAaO2Ge7wI+pV/1IgM9b8sub1NAON9XHLVUeM
3XIRnD/er2DYqJjEYblmNdwkfbkbawr9L5qMv5DkMyoVYewaU8omZEiuurIGvndD2ipnp4aI1a7I
XqwppH+IGKYrtB1AMl8eRPxOy/f2r1zFJA9C7ZT5j25zfREDsQVah452H6DU+TZZBg/9C9wCOoCe
axeTx/8Vj5tnR78RuMxsxswUgq9JuHJbszOjX7i1AOFqaDLbfNTwHqV4VSUmD8hv1xmsbyIgGIAB
uYMbDx6baTFBcsfRE/zRsR+3NNBlAVfaoShi4gkMXG+Ra+tX28+cTnWsoXT5gH95vHVDFaTSxyiK
6KaeCY5rIc7C8ty1XxZSxCEg3dPfoZryY2l+7heyYwKrpbRm+r3LTrziEgcgQWLiqjfo3b+XFN9c
UpFZtBzyU4tqOYIqIxVwF4wJwOowJ5sV8qiaH95htMGAagKhKSYjk7mtGfJ9VfQTGpeBIL6KD62+
Yg1ABr9bF89mPwwHh5Y7OD33B0kuG+ANJHx+ZCLAU4AqEdpXdmvAoKgwfAmDN0XdM7H7u7L3mKtF
ISfaD95MBwE9CTqBK19RqUI2UCA0TLfXN4gdnDE90oHy3Ix/UswXWpeLEvhRpG27Rx4lkIk0F42i
wcdqyGXrPxmj/2PHmiDu39Zwgf1rosVoHhWwyk5DLBOCjQey6eWy5OwrmFAaGBrqet9NuLFDT9O+
77h9AqHOItDVT/frgn6P//avhHtVpfvFAAp7CbP5rwlJOayzqEc+GRY+80BshwXqbtRJaz96fCL5
tNKfwlrLMs/CipqgXVs1j1FgHHWpNauLeNtz0LPwCR4Ia1nEbz8SuOjmbLv+99Ydvye1Tv/2ZUOK
WuNKvwo7E3AxRb/L2SvEV+6D9KQpN6gIqy6R1YhqypcVW26t+DZ/zzK/EOVDPVWnZP4Q0z3HttHK
8icHSqs91Qebgpp+79Nu1bR7rrVQxGVWKLMbHshDwo0s+N1AjgMmJrYyl3WoSSKa1btrx+u0uwCn
s3UrodwxCoK3jKHHcu34uCONQFp99i6Et4xxSWLdkcXicXeThkZHvrvSPHWG3w1Uewy5C3KHTTgO
xM0GVdMNPoNR01+kOeq17G5f35lD9ZWBQ0kdaJ66WpDyxXMhx2hflXXmUaTFnSZiOiQKm2WwVt0B
vwixcHTTAdh7XKWbd7Ct5c6ewlqh0wwVFOba+f2rVbi7zz5Tz8bMT9/+kDvkqMREl4HsmmcsLjRN
DW/jLhCYFRxGxUYV8ShKYp4eZl9tfRxA3ruQD1D0gAUTJioUKJCZvjI191aggidQ3s5qqF2pIg2l
0ybkSl40p/nwgr+4kDsOlJVtMxG5gO6a+qb1E6dqFh7t0QjCCtIVizh465BgLCg6I8llRnKzXOBu
XY8k8X3DGDPLZhlCgVJzpjEQ1i/cfp2pp5tPq0qEt8RLG7+qXEDSx3hEVTgMyW8CmkqrpnBj23Ii
TOky6qfeGzHckSZ3Mpv6j+FwdJZI/Mn+3KmlhDrCaDG8VD/gxPi7U6l62wd0jQM0LvKlsa6dT3j7
blbclnGJBjz5ja55jT1uYkZpUZXSVBgjocIeBDTzxMHPSUKLzzkjbNFwt0B0n6Sc09XVuea1PTTS
rVHmtY1R7dqewLMeOIDTsKqSW+gkPCGfE8Zm11QNRaq+LGu+xOyfTaox+eCv73V63FHNhwYOROU7
8rLH6KZU/MtqgXUZQ6JJUNTZXgzhM9WL+BiEWriK59+AzLeTwCjMX32Gg00v9+vsB/xK4H9rKIFO
rpOmq4K9XjyFx92wp14UR/rC6MAG6BaIaWiAf4zTmFifTTcdp2mztkf8hogAnhcBYG8DIJ/y2evq
q2Db037cwvKXsdNa7gWdg/dLXs+GzX9ELpSPWiwbY/J9jc2qswiKlG9l5cYKoC+8KyTvBkbqoOHe
h3tEXefYkZ9MQu13cawGUnM4x8Tp9nujUpODHpPv6UWcNHWVkFKzAa9DGP6x2mBu6zE0mVI3qlIK
FZPRp+X/UG2VElwB8tC6lk+pTrskCX9HcmbDvkN9FUb8J77gkeq7cV0nDU/LkmchU44/E55k0aEE
NZ2plBCNRO9h3OHcadxa1DhjUTLjzyPhQGGIuuWIAHeq2dD2C3y5XijMgS90srxce7d5N7K0l8W/
F2jXNND0UKenl/VvAOfYBfN1RkHeZI/esdAkwCTCcW4jM2mwpaKdQk0LrvOsFmFetLRQZ5Jxf7Ch
tDTr+gTfQbaAPBGwC1JgJ+/VyYGCHd8PuUp5wjhhnm+vSjd8PPC2HJPN+mEq4QrBfPrzmJk0g4cK
VNEK64S7f9axbakWx68zNM30iuJ9irrkS6X/Dq9ExlelmMrXfTwhQlBWCpw+gRtb3EL203LIy5oh
WjMDOwHle5WAaE3t4A1sO1hTECeDHBnRtSCUSnCylCE4dLFlV7d7wysWMOAuyaiz+lZL7WFM5piU
3hSRPl3OhDzLqabwPaxfjduud/NUI9TTOHXwWzhAHboFRKNV+UXx/mvSos4iAhjmuVyrcs+NOPOo
pFesZ5S8l+gDApPJ066lDBwmm3BB0Ba2qfjXod51SWNKOeNJlhzFZ/Ua2AOtb2VL5cR5FzSRoPhd
TS22zqCczfazNLLOIWyX0X/6A/HxbadbJCheQSJmP8ambQQELvovg9sLMU1rpoWSKXVL0BoqqMZj
ICrXKE5EdeTtpcmG2VETBi9XUQRZ3jJPCZP3VsN5jNwNXEh/n2NoT6e+umQs8IEyt95gH3i3uo5Z
bpeGYUjXgd94SVMeAUSbjh8Yzq14OE6KTF5cnVoz60J4CDm9TOwcXwtPyKKLzZ6FZxbS0wASV5QV
bULrCoOpbe0TPX0UVhgEfhIdVrW+OZaKs6p8WTcWtcJFBdYjxZGRQfJ75LAeMgvAO6l8iGmb4JT7
NjK09YBO6mYAdrAz9i3FpjW1mklZRt6ceZUI7gLBtIGG36BJV/6wpdsbllSwuV53HXsrAuHoo3k7
BYOXXbc2Q5SbqexMhN4UB91t6t27742UxGMSkcnX1oFI/zNZht10zH9MHrtRcGdV4Iv69xRbv1tZ
r7ENFqWbhaN+jjFLdRsWnBp10DOGZ36+PA/+PV795O2wlJ9XAyvf+Twaz4qaYon82zJ+ALUlYh/s
p8xabPRtVAPB6JxPqWBZD5pk5MtG+gl2p/RYqWMeGm+pMfHbGxdJfG0q8p/FsaT16tVchibmVNmz
S8WLTzQL+0vSeTQLcgqeDlPAeW+eZm77XSi0Byovg08iskigF5RiRHXjZiURfYhuIOleDGcM9iKe
FniP0hyyqUkBBEn0vHCOTzN+n8Mx7fGMP7h1mQrrVcCAOTFVfX/KglxeVTBtISJMuUQgZg5t3R4m
RJT+PzVg0oKNm2GVj6F4dk9U7pPiiuK2jw22jn8NLnNR/F9176epXjXZ7BSP8JzNF+eSDSfeTdvv
qrUwbLQPlsoTZc4WnWjIPuQgFsB8YntigBMZNdnVeic5/IKGRTdHlVMjeNgAkT/IvRZZ+FPqNsQE
H0Wayp9QB4+qZYmcO7sUb1XtI7WtlPFLtv+1FlPgdWNmsB/CTBIJMF+V5miI8QEdVKrfayu3Ql24
w0Zh+QhuTmWCpV8PpzvBvqawkZBQbSTgVwjFvQ5XVKks7Zppot2nOiK+PjjVtTpq51HvCavD/cJb
u+wqUzWNIj3JdJaLvJ41yYSDITfauSjCIqng2Ogz4ij8AsqsEFrw36Jc1crMgmwkl7ByFPq5iDKm
9mhwIDfP9Om27JFm5gr1q7WthlOYhZTeOlogPHmEqz40PK9UurBQQqw4HcG+nVN6eIBflbGXY/qu
sy5lipRHx/Ij3KoXa0Ak9iShBFMOFDKp3tKJ5gcdNuMjnZ2Dm+y+eX2I806Li7eS/kSfqAydqjme
RN7KatDSvWnq2XX7iU4L430auNVGdopcGeLQHOJR2zHTMuQx6pA804tnnuSCmtjerf+TbgsMqK2T
wm0ykLc5PiYO2pV43iy3m6UksK4CHXiqwlWeFzN8qT3LYKmtUc6ptByMw4LtOl0WJ91NlFtbctZE
qIWON6gJlbQKrBgpw9vH8F/jx6CU+l3paAF08nGZSlgWSkoYaTn/feLKnVQ6sR262c30bp5yqiSl
ErmStzCPKwjnpp/gBuw5IZNpnyvi7qYDAwG7rRjwshM5/8kEpsWR0VTXMLc+2mm1eFia3Fi/j2vb
IiF+q35+PMzUd7Jo4X+vxdPn1RAavS9WQMyHL6EnGi0zp/qRdPVKZ56t56SKElWCtMaFQ2WVGrQt
yb1IjpolkMew72Jz3kmftzcqPyqiDOpy0UqwacsI8dtmgGP0hNQXJspCOBShzceoKj4JU2xwQrfq
5tzaiVdOa7KoqJ0wxGXdx8UX4NuUXRVyYSFp8gObsEcx/sx1t1n80wUSCdDEKtR5KVpv8OiJjBeg
t+qdTykdHdv1gNCLFgujfkLon8fW3HUTJBGq4jOwUYZJJx1VDqb5dINPgkh6wkg3kCaALThIlKnS
mO4jeiLFTjSagbiplvi5LMKn6QlsA+zhKtx25CivtK0eZiT3HruyYvDRunOpQavwcbcMYS0J+Vzk
0gT2cv/eHQFB1cf4gM7jVGYdVYhltaB8NZZP8NWJASwiHiQZNGclkUR2pSbxFl1aWRb3KSwrfNhN
6cEgPBUK2DSvFT1aOkl7C6S3LIMazNwlEe2GNqlBYJa5w9WS7X+hgkW3H7flumEnNTh3VNTWVe/u
2x+AJVzegw0N9lYpVPrC8t8CFrpbKUHK06m/aSiZb3fDeHedKeqSX/qxbmXLHS0vbT4X4UKbawSW
1InLCmGGwJxyf959YVx1pRmH7qly2lxdWg7ZvCvTyDJ0nfBy0Lat7Ff0OYMmxQNDGqNJ8iQBMY8Z
bb6+LZXxAmJA3x7YdI8a+hJuW3SdExAcdaTVz794FGxNHSK3eUZQ42wXynpLG9OOGURVWpnZL9es
618ZXHIpJj/3av2LuPbnNlHtoRWDzOvnm5Yb/dd7Yl1eWiQzV0CzmCpEjBQ0Ys88+0m8ZFXsnmRk
BZLPvGAmI8wuBTHy+WJZydOfs12M12mAJYpAeEOu5I91pl0wpMxjhCoGLZOfhM4YDrUdS7AGyCLL
VnGIDlIF7IpED4gbQECBqTx65feU0o3rtFKTx7uroSsup3QonnBkpswGLmX+BZ9Gd3aAxrxRdVfy
e/V56OW0wKJ4sGvDyerkgslcsJ1m3ohlsjgF5MIUzRIcagbkcP9jOhnaznufmEv8Q0tCRdAq8i8C
0fFebXoZ6M/jecFtrvKO+fqWU7JNnZEEvJtH6+izmCE/6knz+3W37hiL3cPipYE3L31idz0BOLjM
eWQufLFmy682UZE4E2zE3O0KsuUOuk0Xivb+VrEthd9l+y65lcGFd9J4ZcwZN2Iv6P7dsPQomhBs
qYkEcke/BY0qHci0BuiTnHIWejFDmnQp6DoKzwOzGT8j95VgwE++0J6rwBvJAtjG5YsNebhBGmh/
uLlrUFVd6SnemIcCWq7VkImWKCmGkOzAaJaeR+fYJy7uHziz506rm3scZarX82DkjV+FVLdCc69i
KYluMeyQJUSZquPdq6A6upq/tiddTpfwciEKfF5IVFDuVIvEd174hWd88ZKduKka4ArujU75N8Jo
nAI1HfEH6Mc0FFx0xNiNqbY96Fwiy+dMQuDJ03YZCSYLcbOHnzX5vOZElM9Q4y7JNSbxxWxWYJkM
MG8YQhz7EPt32Uu3rSZtqmXOTAanozAnx2Pr42Wkyxwpnkor2i1hluU9fr+f4ulHo6jXDhQ4BNTu
4GpzkLPBz2gCvvznAWXn57hW5R5yGYp+PN8ICSlc/8jfGBH6+x6IgrYqr1Up5dIVwaqa3lW4E59y
r/3qX6BeLta+O2AQ0xZVhmhxJfwclcAyrprVIxk5CV4ggggglCHThjg6Fn6nGXwLgTwTZjEHej3Q
zjyhwL7XVC0lqr6puVIYEGp3SZ/yE+byd9uGRWXlC43F5znYkJJEehbcNieTiF4+Rz2XeuGjspRq
KnqpiAf6h0fAghmkwgQ0uJpHMjyGIHPkk2vLv0+xU61RJH0A2Pe+kTHwGTnGvnQYC8piQE7tdK4h
dCJP7AULCnYHdrTLfR5/dI83pywgsROjCbM0cqLz+wIieqT4QSOWn8iCkBZfzKxyw6pdrldi49wt
UGVLGtOd0m1WjQTwcnulsOvXg8Ll28JxVUhxzjNOA8yztvFokvXDrwkt0hWBi81ITw2LxAfv94X+
t2XEmTuGgD9s9NPqUpOW263G+BONm2jB5e/eKdKEr4Q1ggBov0KBtxZF9wuTL5BMUCab2OwVOu+V
V22FqbsCPddqi1TAf4AU23zppLS6P6UTbHeX5dwWqsP87gRIG71uyY3yGAvBSTtqAuXiSlQmxSX8
eOevgZhTPaswWBhgCtvwDYQXJlCOqZ+exvqbqp0skt4/XOyeZhEgb+c/YVbzBbEKTG2AdGGo9hSn
kCJ2dpsphw38xaYRk1RqFGiDPi7khRNzGeiyBMgP6aMz70FZGTKLxAL8pDJLIOmRt27Q+9NklO4i
af7OcSGXh3b4eyTgAVVSAzavvDk/+XuKbl4IYWIN4L+MPI/fDien/yV75DWf0JVHaDBXeanZRUxx
gRiNBgG85edxiRwvelBOSmibtWGK50rifXDL72oizZ/OJvy97p0cwVDoVuzbPtK0NjCw86z42Tul
XCvxBXX7iAkp6/dkyY7/0+yS0HO1rhKrmkOE4cbrTVVUIlBuM2OM+bnST6cWDKFM00L/GcqNXF3N
7FQ1KWxugD2HoqSDokLKciWvwU5kkxmVLLS8sImwxGyNZkHa+ayMAh/KEK68BygcXc7X4j+y2nqY
CunGHkXFf/qm8IVBzzwNQiD1G9q6kUOLxXxGBpAxs5cYHBYJ/No2t1SYd2JPIF5yM9tNNJOu46WP
+fgZzWCkLSo/ijOxJBf9tSKm4LhNdqA8VJcyWJSprA2YxTZL4LWMWge+Ew53PLJB16p2TNSz49ea
2oix6uovNRb3qWzetVWdR8vSp3EztJjHBZC3BN1clbvuqX8x7PVZY5QfXHngAp1izHxbSXx5OiT9
AG4T4zUfPVVnJewhQBAkHLy9JsNNDVt1QIoSfhfSGl/PNwvr2MR2ZzKl04W9k3a97zTwHnxDJItJ
+FvIG1Z1k6wZGIQU1lchKA+LoRrRHbhfPsSY9TeVIQ5arb/FSjlPiUfcEWUCOa44lZEylbosaNb6
UNNV6Nk7CpcCeO9JYG9XTZ1FKOKW5k7NDoUG8UHYtY5vW8G9X4XYV4VdcM9VXY8Q4Q2LBWsssARA
hOYiXsSw+YlFrUBDorCjRZnjkep16F1rpNYZbLe3UJx1vwMoH7zXIG89JinFqQmskbaD3cr7ZSW0
KYgXwaOyeqoV2KPcTAuOSg5cFeFBmQzdmiwsWh9XQBcICX1bS52y6FgF9tftae9czQzApkqprVgP
/xHsYF2bsv33/fR2nN7c9iVKUgEiY/bDnM9xB48TkY7/C54EnaENKvJYf0X2RfshcEwQe+nZtiGE
RAR+BjyFVcj4q3Oz4+/HTKlXrpR4MqqsrfnAEJ6mjFXg/yLEQneCQkCCaWYGyl313BRRbGXIFCB+
bs3It6l7umuJs5TO81YfUyS7F+j6aWth6PYWlt4KnaQvarsP91ljP7PuIjtZqTZijZadLn0b+H+y
Au1dM1QFgZZqSckJB5k8WoIzGZCPU7PsdkvgAtubzj/oothseZxrhGxUJQfBUXRwI8jk1TaVZd38
lxlI5LTNtIIPPynJpS/5/7AhAEyYUA7Fz6pF5AR6zY5yKiDkLjETyWmawZr4aDD/wyuJwgHzjNx/
L2ui6hiMBwINBftdZsewSxNfbhOy4qQd+lxYLe1JSl/tSbX71m845y8nkKFOuGggKvsVtbzbHWw+
ImMnDO+BpwwUsWMfr/jB6q89nX6vKGAtOgKDE7vk1p6YScuYhXA8tolUtqdo5LpZBNG6wNnIaP9N
aGRR3LYXKevFdJ7ilmiE6E3IrhuKJ/xdmFZrUhxMIfuDulsoepSGXqWh6JcC8mHwDm4unvej5w4Q
T8GBIPyn6kotBCyDvv77Nl4Zc7qWVz2uPiwDkB+vl2P7tsxZUDARzH4YWvxbqMhp/f2R5noiCWdp
QDP+iB7RWguzTL6k96OOD6Z34iihIZLP1haO+5v9/Z4GGmcfsl/pUKt5zppTF9rW5X1RhmIGj6NQ
/FN1YnpY95voIaMf4J0KS1mERJywV4SjmxpRd1kqDSUInAFmJv5dfYwRikToFpNWOPMnNFvdTwjW
n7mgrwvcTJ0yOfutpf/QRj7yQSC61fFxtEKlPx+GWcsrPGEGsc+TvDWvWSyZ05qp5SKCBGd43mbg
jbqqTDU/e5B+U38fJoLZno5OvX/xCmO6zWIbbORgbSajgdO9To0txGc29iAnIdeQO1OLoB4+HuqF
kTjzsuXqJaSvfTvEmkjQavks3XJ2AuYc0xGajaUdCs5E9DxRxLQCX7/qdlrVx4/CICsXveBfyZ/5
V5P4jzASJ+cEqBLFV1rqSo+Fs+CiU1Ks68A1mamu3UB/DnfpsFKyxLcCe6bpDa4onu6i3/S8CI2O
S8dXbBCYPdS9UC6I3f5ONVyOaixnPztLAq/eUxp3Vaq5IK/NzpkLm6qmFUZvQoJ9qMSBJudJ/hFR
/9CIrjiM3vBA8OwN75AZooVAx0fLu1Zem45D5JpKK46xrvZMLtVdkwV1bnQshK/q6qPtd8XBkZso
Xdg9Gzazi2zku5QW5JkEH/KY75nzRZ1QbHHMxf4wFryjtXYUmNCJ6wjqBIfrYRKAFchpuxL9Fu8I
b3xFOTXn3ist3XeCIQQK9R/19Zhd/lpsOCkL7EuekqgEu1a7aeWDzWecTx/uNvcepTmxsGOzCXZC
2A5xNcuEN8YN/Hd8C9B/DpVcFJ/0aGPX1HkbLPTHoZWMzyAG86xA5MX4C8MBYzLe3/ncvdRbgrmK
p7+OFq5irSwH9WGySWnwrEmhps7+IXwB7qdSOBfJQnh4goiuYyfOHlQ0BU95v7GADJ0UbaU+unUf
g9jczzj6R5hNk8Xt0hiogifUqBJt2kSnkiz6KsivPID9r2yCyx+fdFAcaZ4Y6a2idNafr8F+VCBR
dr8GX1WGkbBK7ZzX5J0v/f6N6HUJbTn6hIpz1zqO+67eNfrrbh7wq2QlzwBJk3zopc/LLL+PALqA
pn11VUnaST76lz4/KH5tz0PYCPHHmKdzsCpZiIhHvlJL1ujsGMOjOK+XkOwThxjIe1WjOYTmdVmb
7ptn0UzIzEhb03SbJ9wcqHUcpk9lI0srnktPI3Fcp0vUQp30I0/bX09N/cwrbMxztP6BHxP4FpOE
0QVuggmH8PozNM5+yb38kuA+Vf5HceeYDGH7pe3vbKIDzXJVfdM3T+RCdhRm7gAhxng1crB2YMQ6
SIFzWYCVSVjKIf5O6O8bKGPhqKC4pMxQ7VLxeYNBdyI6RDGZbhOOeeY820c2rs4oa8hAbfzmUuXp
K/ZYxoV0dwXQTGu2U5k6htvmZdcq+upfhUjJbQbtb1sgo9y1c8Ss+kENBqbKvGnHCY+tIJDhJX6u
B1/LJJAjD/ExFeQAyt15gp8WT9NVWcIvAGrPAfZOP3hMhQ4d3aghJH6VPYx0U1pYs2abh7d5M1bF
jTiyL9+aOFWNaRBXTSulVw130U+6RQ+AVHWqoM59YfgQoTKkfJdjIV/uDEmdU+X5wrTh+QUVSW1y
a2fDh+jgCPL3m9S8DYB5CeKAEGBw3XnUpTrVkctC93Y+q6E3z5Ixb07rufH84l6RY3mKcKrPuWuR
OfCeyt07NVZqeM4sUiWmvYKG5KvEuU7xG9OxZaLhPd2EMkidOzkQ2Md0uuwpCT0Hq16puHerIGaI
N2W7uoms+tHs4+7Q4f78eiNqFSnNTsYje7qRWzo5vurd5ZT+sXd1g0F8GRX5EyU5jKg+UAJv42ZM
k0yjTZWxyZ6mbgf8DOC+3ngX6gtzdJ//KWrAS/JUJ1anOSYjKgWDncah/Hu8a3s6lM76iV5HLLYx
Wk7YKNsNLbJAYk2CNF10GJWf2BRJuaFY4IPcklchnGpdIeMjgw6u+LOjZfB3A/fMlVg3U+5/7uD3
Yp/yYN0E+UnFrI/9nZ+Z1Lm47TtvM0DFw8ZJlKwJTuPflDEQP79TqWBvCWhNr3T8ngz8rJZZ0zxl
uY0qz5ntsOyUB+6OzF9ANLAcbKfsHmz6wbx9E3s7/kw/B0pO2NqOyyYOYXrSEisT6X2fyA0Nx1Aq
bJgKJznr7d2uhJYO/Rbul6NqftBw5cGCEXapNtD7SSJExY1bq3zbD7ZnyyCDxnfZq7GJF2bavehV
s2a23afl/vWsFplxyGOuStMGnA/ulWPNIpS7LyHQw+aM2pKbvlKZqEGcwuDLqjE1eXroV+qr8Qgi
SAnv8ELzrUVKoanNC5zX1yUw8/tbMnVPxziTNU3F8kX3vqHdJkoObG0Ahf6kkrM0ZRqdQH7YLniO
V91UnW2b3QpN/aolKheqc7Oywc9RypgmWFYhKeFl0glxAYJBQZc+yFN+z5HKZfDyAuRF73b6ZLD8
vydp9KAVjLk7SnE/pF8Ye0/gNI2qmnOVs79uhdUlGVRTUD8WEMAlmOkVYocuVk9/XoFK5x/VXPxG
ii3jhJcxfRhqugNufaC4z71bJJem54MkYTTpZggujphqfpaKbAE7rXcsgETSnQ/rk7XyL5Oktu6f
0xsU4f/3QrTBVvFcS2++S2gk81DiwpD7vjBDh+j8we51FiG4YlPBntgiizLAsI5RmXowul1nuWT4
JIYCbdkuVF0QMgGaa9JdRNr4ImO+1nuuaeGGSUsOzu3RyIh7dlUKF2MMhbTqFjJLQ98gb2AFWX7t
EziKtNsZ7HtRUgnYlaMrddNp+/SF+OGvnTMVbNP2wlqVigZCCicspxANIu5GF3ZV+bu6mjpPKMz/
uO6rLag1E2qID4Hoiat/RI214cAU4AFD2vwgogmG+Zs8LukWV8ZZnzhYZZpGTwwtMXfNDSXA/m1N
aG1Fn0IK5ys5oGsOf12hIdQIx4kWHxfsvZIHLKzDyZ5sp9gfxobz5L7PC+fu0wDBj8WzLQXKF+Il
bwTRwHI4aoL1/QYbRJJNfaQyqzFgM+ADJbDONjzbNV0LxEip98vCqTJIxcO3dkwAf//ypqDeKwn5
jOoXINErshvr/0O+Ln10QuWs+nZLg1jPGXEV51Q6EbGbMd6W9crkdNSJX5cx3bP5PVmphgfkqO9C
rX1JStNZ/DyXegOmHPBGVXVw2PuJ5HBpr5JMLr6a/yuyaPjYomK9SaCKfFVJTNSh0Dy1GqWukmj+
FQ9EvJyhbLZvvlpxAmKG3wL1lGo0A+hQGwkT3VUULSJj6V8rA5+0mw6F33GaiXO+Dnfz9BpCjv4d
F0PhFj6DS1iqkShbSTHke8lJdjHmJx+e+B9+Qm7AKf9uPPbEuAvCRk6h+IgrTXw7ARTG5AmhVW50
Pbo4W899rRqk5mTBrAqwlLol/Vl6sZqx12xaBEmNkI4sz1mIMPRlWWxAG5Y9kV6VMxv1nyww21IK
lWOWnHyxqUMwmnjIQZrbNVRtiEdBfbn3ZHHPyiPOEI4AyX7LSKb8Mwk3TiDXz5a0SF4g1dlPW6tS
ltTE2hnLm5cLlxWBv/aOel+sMlbNc0i5JKdevCUM2qaRnOfmV6RXN7b5zxJqWNxFNpuQ9IGhLLbg
hkwwrSFzdd+s7O9McDN6aIAWdUkRhju02XuvkJYhSbvcNLOxdgJU8oOgLQtjLjfIMyOm15eizIeF
2uC1OZ6yTmDSy+85OOLdMpGCfD0sxJEOfb+jYm9/smB8iKcAxR0fxhv3YFziIHxgZk8kqAQX3pth
3YfpSaqs0ijCblmCrypOXKzT5nFOyxbR1Zw+YRBQ2m4462tYqP8HNVlKw80CAUMFPe8Doy6tG1Np
H+PGL+53QizR3NTBhf2t8NfXUUjfVQyqTtOcsP3oyIP1hOSClnO5UXjVsopnMqfmuUArdxoK8JDb
C7B1CXozUcQOx2k8b+evKWCXS43vUIwe0EYVUf3YujLsspuonziDtmF/n1Pag+Fofh967f+lqsre
zhW+6meGRObzeXLdr0R29Rrb8BtQ7UunCXArdYEEnrV6ajMU3H6HzlbxdCRpnhUYLOxqx2AJ+Lmt
PXcmeGn9UatV4wmgfX+PqwHom4a6KJcmrqxfS2trdE48czToPlpe6Yzn67s3ZuQMhfp4dio7Y568
czdLhGhHQKUNaerFWm4xfaA07qAxUzS+XlT8ukZQcrWZIHSlIxMlIUXpeEK4/MQR4AvA4qpP7WAr
Azac2vTeQYo9J/AntBV1n5chJqQn5817lttYh/59cCFTiQ3KW5hCrH/zqkJCVLdYPPzly2fuuj0n
qmUTruZAciskNG/+GOkhIK6Kbjj7iMm7qT6VVcjJ0W4KJUJn2Y5Q49mnR5BTmjmfHVbD3p86IdKD
ICkteKzle/g4G1hn+DVe/DtyeKbr/n6dLeo+xMdjbXrbY3dELVyCcVYLukoK1eTrrA/H0CO0Xer4
R7xNeQ3w+HcJIWHO6tRkC+WqHXZaIgZJIAsjBaae9pk3BB9aPKEChXGRu39Jze8OZlZ2h8vI7VYA
rO5D1iu4MULaNYgT9yKaDTeNI++JvGP85x3jJ5y5FAyb+5U+p5N1Wob9V8uxWi3fo3cspIQhKtic
1okRhvh/QzJv9Tjf2Unaz5r0nz+3dM3zOx5tG8o0UvxXOjBSu0AhDjKofMQpqNoi1ZXNiWOHQSpH
Kb/kozdpo7r3/rnokKwPt6tlpEOAo35RDI4LroVRxv7CXL5u21bzePGJBv7SKSGtHXf6u2hBAbRW
U0aBEWSO7vZ7o08YgMSOtRRNklYOjnvTUzdNhfnBVAEXL5wviBrv7HcrHGxna36LJJzmJPtYEfwp
jGdwZ1wOdcCzodKoSOV8RdBgdcKwiPrGJx4sOwz/HGOuupsdyH+S+Hz2y+SD+ViDhBAS1E6bD2Xz
zX/OWL13J77Ilw0b3YZxtMFP3QEIuleWiwZriGCocth8JANRqKZMbR+hE0hwVbdX49zWmqRlqz/h
s5nlBslwJbJk5kYcnQoMuDvinTF45mRLDi46GnWVzBcEdfthwd6R0EWOxAR/qDamOQX7/H9C/+mx
rQEaHb3+JhlJq07SgeTMAruig8hOIiU+yWKFyzLzstVlrn4D06PSJaPjRCWiUjc98dAu7qOiGOww
qbwkfyMP+clBleouNQimcCt3y4fXxo+9MpTR5nstoAY7o3k/JDQ6hEYjqSVGNJPHVKBN2BVsLYUy
hu3f1EixyFBEilfTjSQmhYP8/HHcF/DmDc7oPSpOX/0YzNunc1KRhUImbuIobFO32m84i2xQN6jM
f9qfAUEKfye8A7QxLUwdCShfb1H0UmbbSTaV0DYTRsUGrQZzc5GheMH+lMyBtSdYhBCkMYSKkctm
gX99qc9bYUaL/JOeRE4p3I7GnAyWv7LdJWzujidC0GgdPaUobOW0/2WJpq07cmuwO+37nyTidem7
RrA48fxeX3p3+FCDNybT2ucMmBBXyGkgeSKSb/TIFPaN4YjDES+Id9cTsqws89/CoylyiERErI9M
kkmW9Tz+0O94Gb2p3LlRNMi22Sie2pw7q5pds8Av/X5rK8blfJyOo1W8rKAnQcySdovUFhItNbsO
WLQcSGovM+L5+/YIJzgL0M4G4cPTcq8b2nw9Ht183zxadWrvl0mvafEdAoebNDX+4sK4EnLZL6dH
XYFTE/bci/9iuew+Mwt+XZT8NdeLJO6Mlh2gejvlWCzxNdRqm771+NkPWAQZ/SKvmLLdlgmKQ8E1
UiT1LnXOaCcrxNB0oMvbr69H/JzBuP75xK18I9Ayw5rvgDYHDm7KjMRQRlSRXWUgCPg9yNRh9MvX
NQyBB+VSH7TqXLydtKgRzl6UN7585Th09f729Zvt9F+DadRKRHTPRXoODlXJAVAQeHmZmkw1PalX
lIguSfCQ/Y6hHY0drk8txqtBKzdr7YBlt4dMhCodP1yXLFfodFBne/6OtlvhKmg7rd6+av1xf2Mi
B/rUN1eFqhZWb2rC5jRQiAmjz2fuKpcHmNNz0VX2PIczPMKWPkvDRczpiI2NBL1sWXUoJG2oLLa5
yGnAP1n/oE6pH0+ZB8ji0NFng64E0jeWOzs5I9CU6P7wGLH0gvaY14bkRofpDWg0XBjGPo9jROnL
7gM9xNPwnaT9X3zdtElgU+XYOMgFTaWmY9yEze4dTLvNekonbxtq+MLGksRUfdAa/vBTw5244GwN
J48Rj1ovgGiiQ+OsvbnyxMBlyPkAjSyutMQoaBBsf7oCvWpg8eJABWFRPc9FfAROTdc/zw9hEKPh
661U/I83p3uQT4k14RkJiUFfBUlq+/ytWEiiiGF4z2BOH6Yrvhdl8B0oowcsT/wxpi+NqWM1ihav
g0RiB46thipwk5gYww08ORDH+OfLjsshWD/8PHqk+6Ctcb3CLFcgv8RyyHTGSO1Uks9+V0nOPwNK
9K8EZaqqRfsHxCWgcDgFTsZiqe3bJ7VjgcWmlFLUx4UdtcrI3vuq+OEBnFPTPS+mwM+cb8LbHhUh
gpE0mRSANbJd0NAB8/9A3dh+UOOLELa0UoAYHkaeG5fubgb7ngjzDhbpUYMnmkSzKEJ8DGl4iM65
tS8XBVH9f4ZWYPTXapLz2jh45d1miW/IngPkwHR539UTzFJLuG45SlO8NupQF3AD1KPMfhYT3gat
KJq3L8lQiSpYYmrsfJecQcjiPVF6fZ/sPYc+Uyzy3qH39Su/nn+sENaF8p3sxFyg+brwsUV4iM3p
MGR8uPLMmY0dp00ySBWB3DO95hzBf0zi7txqwYAV+mPjaNKffp3LWNFIuACMvF9wvOlb/1wXhvFj
6pRArELHoxrsWTHwDznpESF/3vOruL9vbvD9UfelN5wdeTHjAfSuAAdEORyO4qDoIIRtQ3w1/IoP
PbgziLvVhyICJ92ukI8En/5TlvDJf9+APu6BW8TKwrmmejsYupjZf3qhmBPrhERwNsJTQR0GqiJC
G79WCFtpn3Wbef/BDHoVWwFA4REWvx2Ve+HbicZNRrDu3XI9sOH654cVm6/LjZscFtApcKFGQ3a3
OcNZFpFbPGV+xokKpgx3gGS3nvfogy+XYXmy5SjTtrvmyO9DSq9PpOZmVJTTYyVm30h3ioJkxtPh
7edl56uGKuuXboqJTYVOxfAp7uSODzyQonOtHlKrU/1meqAYHw7rqejH8/3p2J+wg7UiUbsnYg1c
niQeK8jNu6xUeez8EypC1y8vouapG6JEBenaBssjQ6Bs7K0mGAPw4fxXt8dktc5OuDSHAQgj5WLS
/Py2rl2BzbgElMm9MMt3lmjlgohCBrC08NstLyKNLpe4lFdYQWQrbqigU49wuC+g2eBK0UTyJ80O
J0cGxm5EhtoUMBQ6EQAPwkn22O2icnLkMPIcPt87gBIdzWeg1SFCGhFFYb5K+RNy0akx6dupfdF6
9ydMuN4PPw53n5pf7N7o1omjs66sdYzAdm0FgPiAvWDCgjX1fr2Gx6KXQnajbOlFEL/+CNgrcOdI
Ua+qZn7DXOHueHvDaG0+qBE9USsXNJ1Y1Lr5PTBySGndX0Irz5eJP3s1cq3fs8Xws89tTZWsYwn9
8XccrV7YWYHezGFQE0K8LogpS6IxKiEQ+o84nYdEvWCOYJzsJSn6K+Toam+r5sZNOyI7dZeeHnbb
gQFnhks4tFeXiDHLFfZ8RLu1OpmIZAg2bquU50flAmUjQWg8BIrMPMLCpIQb5Q58WBQPhRcuK39a
QzwHbxGbOtVzbwBc7sRgaSTHGhGJCHKOLUCs6ujpkvcxmmorYMV7GUNtDmgPtUKsJp7jHTuh9Fjb
3fVb6xnL6oU7shcA2GJ2iBfplA68dF2N2xIPutlVK4CuVeO6UykWpk+UBAdbHM4eS5q7g4unzlRA
4stPeQLGazHE5VEMWTDGWWLNNQsJ+WZbbxkEbtgpoucVn3WMCKOV2u7o4bRAZicv5F9G9NvLnzqd
FFi/mUY96Xo96LEvnM1fTg3eY0a9y4DTEkNeZ+heEtUaWdu8M0YXcBWEbHPTDxf0xzMA+0s4FZJ/
v0JLtEMs1wc7B5ONmjW7CpqScBqAravmzXduE+BpEZyWE1I8dYea57NxlE8BlhGWBrBxzrQS7UnN
OG56lFGxoXs6Xj93GF4XrHeja6Yzywywsd+pq8KQMNWmMIz88WhXSWyGwSIvXz6x+jRz5IAzyVTs
cez1Pvdjd6WwTqznRgkC873fC/Va5togDxQpF060IZkMIfRtQmf2gX1mUcXJetY1H4IWhp9xRP/F
tFDz3EAc2u+OdtlATsDpY5INU9stnUXuWBVZcxJZ+oLKIfKD3KtUv3E9fjX0pr5yOGtXG1rWi5Vq
XTiV79FUqEWVx9gHSJ+i8YmNdoQ9TvEhtn1xhrXUqV+KkBXi5OWnr5k7S9ERO4in3ABB8U+e3BY0
PQ3E7VgYkTcEhd7affCznRiHpFqdcSEJEC2irw5+LdUv3+1q+3geo/AjzBA/f1rcQRCyrb2KH2Nj
IUpYBEdqWXN/NudYt1GHctGU9ibwmz999DhIruNbQgBtjSU32d5KeC+vtiaMaq5de8oIcgxbIy5q
qsLyVjo7BQQihw5zrWvvuFyzChsxvYJGNu0eEEKS1HmAoAWYkm0WmYHvRpgFFOBDzq+6J4eF6hgA
8Ko7cxVU07A8g9O+RdfWtadSQyEoyIUcxKe1Mn7G1XO4pcWFsVEW9+MPqtAye+ukxLSeXzK/b+O5
bU2r5x6qxS9vpe/fhEmc+PD654mi1j4msw4FLyCDUlHnNvlOapbu0xhgPPb4OixE+YFga1yK2TgB
cYm/BCvlpm263b941ThUmO1BgPgU2o4QbEDdjik7QcwG7iY/vpSD3N/k5pR5wLdv8c/u9tI1IGEV
YaM4zKj1RTThUNCtloWh2zDCLuwe2BkqAcoWq63mCEAX3qjb6domzmLMJbW9xSL1c9k4BfbQJfPi
HFYxbx1+5pRmSUo6Bx9Nr6+OsARuicYhdz45c7WDS+WDlhCOOoNlI/XU5Z3tGf3P2/VJSTS6hErW
gwKAi+QYDr/9u+x+JgRXxcVyHNiKO1CrdEK5WXJwe68SeuEMRVe+OLo4dfP3edzyXzbItlU6nJC/
11nn0px4LoJGo3aRRHd3GG84c3zXAJ2CdmTb/DcBXp+ulubHpS+gC+vT46UEdfiKaD27XcBxqpBE
0ijgE0UWk0TOgRSTWxwnqgzJKhH5gf9V5N96kOfjsmnREaKvCl4kxHcJ3SQUrfq5SS441+sXQEmM
WBJHwseokLv+3KxdMko03pTw82U+gjznuXY1Yj0cYDc4+7/ZW5ycSKRNRjO9k2ncO2ai2yQlmTe1
tJ6wKU/AVN2BnSGO0rxZXKNyOmlHIi3NyHjButwzmvbT+uHG3djrXD01L5E6xaeri5B/tUfymjvb
fREsfBiyVO+R7dJOQAy8aNosURS5aW9o0ZqtqhozRgB0/CHzVsv7uPSwynr+C5QIqbwXCfpfT8Yv
WYcS+CnVU5oK2Z3nDc33tYg00jEPNI/Nqz+5SWg1AbCyXc8zknHEpapGlVU9qjETVWI2ec2QGJ6O
aJxWW5cS3mieTXu+wKPKkG3vY9Gxk9TV1xJOESxouoOR6xoxicCp02qH6zuZ1iJxuOLR4tJMCEgh
P+fciRs0ZAs6hBKXeloyJ6xnVmiAMvW8IX2bpmY4vdq065qJNMYs6rKzUdJCyW8POQgSES7Kx5tg
qR/SRhFDBAi4BmoNpkV3Z+zuSf/gF10HIWK3BNXLqbwXg+i03tecRbjQ7Ztyj+8m7May0TtkRfTA
kNXga2tA70xzwPo2qu/0LxVo7N13vn4Y0Q8BvKJs3BbU9YbW6Yc01OgOyRtwVNBcoNH5cGFh/a0i
G8MRpOaFL8YvBYiP4Ct5gsr9Lkpj46samj/Hry7Kp6BnRIMIBmdslwJFgE3yeu+a0rbdLHJp4jEC
OcsohBc55moGotxzPUKww/qk7vnUWR7nzcKhMf8HHYY8Z9oOku4OBvfDaYyP4OgojMZXM+5/59aJ
9R+rnq55Xj+5SrZIHWIASX+2j2JpBW3YsSzcWNHk+2XP0RtIFOMXf1mOvmbr7gue1InJ2XXKgsfC
dzpFpxGECaGqPls3TkwFH+7MDhIwOTvNBscYbGLQBOG5BvbJ2VRRV4Oey41b3D+ylwutxga0c3GP
lBFGVdoMK2AUcM7LvP5mGuI1WEkywhhTMA7z+aB6FRLdqmvdp/HRmXwDGcE1PBZvEZXUGARORXdu
vyS3E6rxvcyVmb7wIKzRWJlsuFAeBA8UJ/bzd+gV1JmGlht3Z0CgEFdoTzbafzYtyjuyJgIbTefW
3RZHypKL/1WtZlxVrmFOjjmP6TqlYaYf07mG3e1bdswyHsbHG6vF5b9sTwAOjjzED92lFIeeqXYQ
Rs2AYP4IRreIho4Iir6JxcrsnyQM3a+nnWVVyrN/QDq0l5/SZQd5smkBldLnqzz/PxhusBjXd9Yd
Qn2pXRcFt9Thu/r4+M1D3pWM8N0xgeQ4fOmogFxEzXZ0mAiyQ90kA/Er7melctKjKnRNbtBsTvWy
/cVhBBabmpDUWXRL7b6gH9JXnjffkuxzBdZE7TQUJhVTyPmXll0fNZV0/qVo6uM0fRo9vzBOEqDw
gyGGCWwrGHjQqM1P3KoDyXhYe0Ek0bJgl2cuD6AQODVPE4A4BhKd6IivupdrMhVqIxPNkATk0S/7
4aaxE/NP/BqpJSPJn/xPiOCqdAPfBXt3op3hHMm9saWLIm3JJRXDQjiUPNKGX1MyvCd/29+B9o9s
clMATjBLKKw5HhSCI6JAU3fjUtIJ3QVTVF2OQITz1h7y64cQet8Tf29mMN8tAFykie1Ke/V2V7p9
IVH8nZK8etHJ7vPVM2GHsRn4lu97hzdlvmu24kY+sn8WmyV8xq9zRftB6qkcuSmz0yALpFCLBLLF
LK6H9niCwbkwHITNDnZgo0QcLe5k/YmEYbQ62hZiaw/q69kIJ5OculOSd4EMQ4t9V+n3cCpDxfpO
+BqX4mWvX1/WneI3ylUoZ9O1cCxEFKQlPfnFpzAtPw73i3d61VIUAHuSLuZs7Y6m0I31aowWluOp
ma7Mx0Dw/0FO3vWdwsNmp7e6HcUqqENk5kqyFXAD+EocvRhk60kC9L3h4+MfaithZC6lNuN+Yf72
ZK0BYpSgEy5+uWu/iYFStJv0UUfWAQJzPl7qWB7ZpYlibGSukXH6WUy3GEmpoNJH0c6uTXJ1DQhg
xZ+6rtxFDBh1pkmtO43H+B6gE40YacI+j3FJ0VTWJ+QkO4VY4H+XDQNwFWHHW5ZPLPz0TH9O52mF
wN+cCxLt6zRzAhy4ny23NzvbfSvDJZ8c17QNHZzMVicUw2QtAbz94OlbgYe5IpgRUpqtfQx1Kx/g
9TGxcoG8PhHKDWfaKUF1V4JS+bpkBaBTcEaunhD1uW117T4ZDqOua/xfZ+j456ekjStdNzlcXdiQ
MBZtYpoSZHvz7WbwVMqjiXnQWl5I8bMQ5mgO9ir6WWTQb12OD91tF4tld96C/MTF6CcVrrdiYTBj
MiAw3HcpYZ3ljInOl5FDl6/Tl5dqalx32Cg1JiAongh7XmJjmSd+MyT8m9B7qk62Mt8ADb/koLEs
HQPwlw41ZMDhN7wVzEsEr4IORYRb7owWrjmSJipSSuVgqmnZygjysM9nHuxBDJh0tTv93gCu9Byr
hDXI1l2jSQRd4BM4iXSIBNKOTqEwAY816WgJIAlKBmKJwemx2T31hds5zPFCEVVJETqALkSOTDc7
dpIdLM2aevpcCOoFQM/vwnFPiz8nO4/rhWndkJq3PJX5c64n/6XFlWXHe21KsOuQkbdBTYcRGTZZ
qmXxVsiQHg6UB5VQhEXLKUX2+6Yx8LU1chb1bqZqHaoevFwhH47j4JVMO3IELMC5/g==
`protect end_protected
