`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
R4yddp/fbY1YDyWWGOmATrbDC2EUoHwACTskm5ulM0sLWAFG3bddsZVEMoCH4uehNQwdy/3hSprm
7QLbv2aW7rtprkWCLFPPnlo6xW1mNab57kQtkaQbH2GTrHO2adr6dNZmHAaBKMOP+9KF6R+SS1/y
9/0e4obJCj6k1tWbSYuuxNgYTKr+ndI/KH/M6qCGGcwYnu0k36d8GQKw6XEVyEtmnDNconDOhDcf
Sy9VcXR9kh9C7ePfYHzQ3puXUTlK6abttOJ5JAQUbCvNkBrwCWUc2ZDXQINWttgqaCceqg4VcN+I
UdvhQDTwe1mcbwfqawMEhkCStJ6qamRlvzZqjA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="18TfYuNsJURIjFMoFrrGtXQoW/MkJArlFwpOxrnqOm0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
xw6GcRTPKIGj2JLsSyaA6oe0yHcxHwQ8CEHpVU2rbSezrx/5n5LJYeMeTfPd36IiZRXr7ua8FMsk
7NFAOWdfb9AvAOQua2sDhOTXHIJsuNsCcZMrcGuK5JKZIBo0rWY2P8KPbONJ7Pu8M0iqqjdq5dRt
31LLmykOwYjs7nK5uXlj9CaxCucdZs5s89heQP55jrKoFsuB6bqYka18ONyiyoFbJSUrXu7rgDdR
kr203fLq8/ilpGQDZpLz2PBPzTYtY7Mjcy3Fq5G3Wdr6tuokl7/adwiOhG3h8swadwFD1SeV07if
AKIMiL8Hvnzcpq7sRvSrtiq9rycuTyexB+PbusWPRekc1VwXxvO9NNF9xcZ/cKypUewcH1+N4l2J
RjRb1elm8Jm/v19nAiHSUNUDlwsWEwozEdjtvskKIJI3WBT55YTsEv/Ir5jh2rZM3yJomG3J4Fp6
8aK6/QhflDQXNr812nRKYUuRIw9AVYp6coTIFVHkkBtqKciCy+uHAaxL7OmUMyo1rsuK+IHolGQu
LNdFaQ4DYoSr6TI5FzgpyD2yq1uTZc6t/oFp96GYvAJo0bIk0WH1648qQfWo6VXwWbLLTorB/2jq
V7SRdJ2DXHa3QKTqHL2lW1jDJuIXEctqzj4VgYjlEtnxJV5aTzhUxUbPsIzCm3bu7WamkRO3u+6k
3JZ5q96U7HamuWsOK9OV5JH8qZJ/q5MnCM6PLTxmd0efw9M4leljdMRc8nuGFKzKNQkx/9iEWvVo
PrHURTCY0EqRtVlTs33DvXWaP5G0lESNaJwdigxDd8+qH6p+vDrkNsvPlpy1YpMOLopuvWIYUJo/
LOeLNMRcCcxx26neavNuoA5Ljv76QMGoVLEu0zZzXlW8Lbe2+NyJYp+5blUlWw0zaFKBOJxWEIqA
mJ/MhJMdfj0ED+mQ+0s0zVxYHyEFqhZ9DFJZhDkE+hnMMPxGmdnC9vFzvLwFV3ch6VDpizMQpNcK
HZ6JeY461OgmADQdDdJyl8fKYMXcrJcrTn6v2W6J6IjD0a3MdUKmevrVvGdwjvYRwWOjrp2cBZbU
RTF1vGRQ2VWgyzikUsMZbRno6fiKT6gkMyGprT3rZuxU8UJg+ZbVpgt7/3NtooVN6ylYo7fi8mav
cyLVlsyCk2WNvL5QThuJJ+PIw+oKUKw5yOGbIn6FJRVFrIjFjghJlZlxfhfXLAQPPmaB1N3JMSnz
x/iiGVCvr5Sw/b13UbISi+So/hSQ6D57uAeUbwclAYzFFWLQgx2SCk6qBddEjcB3rOo0v5OpqQpC
mIYtTF8WOiSizN41ArOqcuEtqKfVSzrOEoDmMRQImAbPxPKag0K65aZFhf/6jorFAf5FNxHJQAji
w1Ngd1vinRCDLkcJuvpc39wejo8sYioSwV2WerE1J3AJOO57Us9Z44Hir4NeKETTIGtbyzdwd0P3
0kfmC9pRrAWU8oXmYwwweayDkREFAaqFm5LCYT7gCxMSq6w6LvUQLuHJ2+1CbFs6NK5unnBbBlrm
XvwZ+HyBZEHRMLtcYZtqslktkFU0X2rPCzC3CR4vNYrMf1HqRX3mlsXsD1lEBzwlCV4pY0R0K9Xp
ByitP9GoflpSeurCPZE+loQgYHAevQ48CIx0kEVJXQkUpxgMrVXigBR3ZYNqZrz91vzqh/68pfFU
cEt0fzkreTH64fzjdHBgyCW02iyrJFiC1BCAz9h+kiavo9ipJe1or7qhL6BwIRwzaYaEhXMAOB98
GYxH42798k44db7Qy77USpJwCOXG7KAjl4M7SwxgBugmgjz/LNnuMx/T3T3EkFKPVWwEotGQJxl1
ZRe1nlTgle+ylNTMHloEvuiyKrY4FHM7shEyJwZZBvlnXdmNgFuOCrZMoEeR2cFonHudnBH8l108
6DNt6MiqhsoZBjHVYnTuA+vAqNgy20/+1co2lsKeud0iIA4IXZr073gqvJpSJNn/s6XxqhY6LZBP
+kGZHb4gPSYcmyUcG4jeB6Sh91Wkp/YIierLV48z3YOTN+vkZHh2rOfA9DYn6VMMs7ZbqOJr9t+P
1Sc239PRyOp/NI+cLEW2xGTsAQvQYo9q8VGgkpFeHZMiRoGdCbXbNAp//41Y
`protect end_protected
