`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
lc+srumMapb6tEiiD5vH2jOXIvWENt4Ny5Es5I70oBqIWeJUL9Nz3q8aMrBKKaR4dOvr3g2Sfyb6
bSOtZQn6c27M2qpmM3avzl9NYqB0aGb53WKabVYgp+q1J2sPEgSmkLdRfHcxZTSL2X/nx9pACrex
wOR1VXL7GzpS2Vcjh0eD4vRr26hFf12n6IWwTOSXY1RU9Q+dP6BNumksK+Fpd0lAKf0RPoZkqPrN
tBn9Yiad7FrYTOCLIh4GtrEKuLuu8eiD6qwbH8A3KSGxZ0eh1PNIdiiyHgeEovBIaNnZgI9U7hWj
vJl7DdTGdQF91zw6F+8OnuOkJJfQF/HujUCm4w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="sVcH1jhsiUQvAuBOBekBCCHbgyTsrQUN0Ler/gqS+Z4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18224)
`protect data_block
oStef3ox4KYeLi+/s/KHVCwWxIiwYGBuUQeczAV5qMnx0FhQorrSnSPOPeFVeX0m/AlPz9J7lmp+
xgNvlHhdOom5ojqWi2Rb/SWHEupK5YdH44laN+AreU2npBITiGFh+b8hAJEoTD5Y15VwwCWFq+Sr
Sh35rijmBNKfjeODghMkmP9dGRS7yilz3PxtRemdP7NyO2Gsni+tCbAjw4ePCXbeE/hAyAryTckF
r1U3fecsWnW7f4rJ40MAfM8LaIsMJ+3qXuayP1c7F3MpwWUHNsBUs3PEezMdfBUTWKrkg9f47S5x
hz24uo3XWwxV1iB7G4wW9mr8iQ93XgdCfKSDCJTfE7eWru+gd83lwmtkLAybU5Th/6H8k6wsZQj7
oQQBoy5nUJVGUhxHHRtpOcLucQ/Q1VwZx+3DDZu7701zcruoJfSxe9Xj9xw+ifrJPIW9Ty5lhA2d
fd1CZ99Re8/K0qmpKD8K69SPyRpr6EhmQsAsytur2RiEzA3CX9tdQEOIE0w7IUIV9TbTxbXOCz1p
Hk1eDQQkWqGyjilouuwJLoZ0WiLHD1d7jtDB8GqCTsq335mMujfj0RfYXGAmjPskFSXW0Zzgvxh4
o6utQ4cNokvA7c/XFNEEgl9BC9KllnfldVVBPS2gGuUY1zNrfkOdScs7j3KiVIxQpVyKKQ0++oEd
jEpHR5k/MvJ/rZJMWLf/cDoCbgoEMZ4D8OQjvAMiZAGoIpAbEdrwEIyRQ4iEfsyXMLJK8VDeDFlO
eB2ecdCe5TAhfNBFPUQa6yzLKcDljnrEf1EvaqAJTf2345zlX4j6Hjq9XO8E/00D9v0GtgPmcgFQ
bYE3GhqUNBOMbPBKUemsFzMNqPsPBHNWi8oqGykxYaHtmEX/Mr0bPlJ13LRYi5kAJLm+P7IRVyno
HYQjyLsqZIC368JYQ8KiOj4/VSnf4PjkOl3UAdLKA7sUaRxGnEZGY70GuC5SCNVPwj2mHIYnQ5rV
ddstB+4Uap3f5vxy4ikfPgNmuG0tcNn38Dx/S+LswIaTRfjA/8DlJF1MMNNCbXdGxvXXr4LJZTOA
1K9brKkbgZt7dTVG912rXAek8RxGgSs/JZFbaA6SlrbTmKObqx0HtwM9GkhaMCxdf4J20pqlniv8
UjG0VKcT8lRxR7DoZTvI0UDR+SvMMm7rkHCjjWL2CwkX7nDSXwqnQhrEa2+iPsPLMOxGRvkW2mIW
MSancHLTn9u6THaotNw6VkDp/zEID3zQeDH0ntAzgCmwWGpxyfv72iLQUmhqBTL9acfLPJJkAJbq
d08/2adodVPWrx6JBLixMQHZi7IAyrcwBT0ftHZHN48gAj66BL/TxKs4xmAqVFPPEcx6UnzdaQqV
s85vrobrVb9WFvatpJq4vlTIdM28MIDEHc7nVe8xemdOz3ehfKPJiErDXY8GdEI+BBIcXgzm/A00
xR5mWBVM1XFv9GR6rGjCZfabxea2RmH5pvb4XFreCa1GmKfx90pnYgnkvyRuvSxIv9/62pYewc/9
8KgGifS8Z7T80Qymc0Wfvcqy4tvFww7B+N+mGHhAPAzuAuVvR6n78f4h0qj5PjsAEOYPqwzya/em
r099MyJYdMKycQecVhmMQSBaKBpVdRmIbd+Q0ZL1OvJpBu+q6vpLEKFCxCdHND4TzCzUsss6UxJk
NGQcmbeXZEzY07J67uFKTXtc+Y3YqsbpJMfNSFSR1o7JBr6ApQEJ8Qw/5W7KqecwV/dKdYT0u5tn
k0jVNE58vfo+xMHKSqxIdg07RC7gjFJVn61uH4pv4ITNDCwlQcw/iISG/K7WVga3ZcmrcXeSDr9I
urj/AdwVaAJHly3lvBuch7DvwVD5O5zdaToE2cAtqVEqHC3Aid6oZjMpMFhg9eXA/Yskfl64XggN
q1Obs2mi+Bnsms04fJBEAjWu6jB1MBj+2LO7aaiV8FlN51bSkmV7efCTgUTvhaHQ06vewDMaIAjL
0Ykrknj3NPx9h8m3H1GNPftfFxJblQxUbEq6qi9Ua8J4zH0OAdvF/0ssSwomsqVvGAwv8T73a+mO
yLat/KHYP0f1KT8MUhAFAf7Cwjoty2lUE+uBdlnQ33l+X3jgEK3HoQDOFTSD1Kx4lbYEn+h46ARc
Mvm0VUzdgKggqHsgGC3aF5/J3MI951tTJrS0ixBaJJaJvXc7fJc3ixK28rhFJTT/ToXrXQrXTsJ+
dlGSl7p++iBghK6BScu/DqUDYrb601m4L2st+u8sN4bIiMVNzVBy8j6nLme++PILGcCicjVjdP/D
ps/2UXDzcZ9qBUf+/2TPPskYdu6gGcTiI/lugkfZ14UnmPMcourz7bsf77TauenCfDfnKXPvz0TE
WxePGy5+K5aWuq2fMHJH6jX3+M3ewDjkvbz1XU8BgZPA20utIoyjCHKmbNr/HD5mF/cXHVaA16pY
CKQ5qHwb0vI3eKc76EugNYZuSiNE+JI0HPp2iq78glYpJh8BJcjaQ+3BbDV3Xb5Le2vmcK/0WeSa
2Rp82Rg4Fxh8rY2LdiPR0ifr6X0x8F4L4G7tWJ8aVcO/hek68FPxrmSyiEpg5yxbyqg/DfsrBkMc
b7sEC52vYFEZQRDKFJFZel3Snqbb10+JeEIrIp0ZdQy6BP6NxaKRrf5W9DJ+ZFISZLfbg+a50qxC
bJNeR8tVJ51CYeC/zDpPVt1Le5hONiB7aq9KLO50hrSRBIdI5lYiwP9a6/TKBAg2Wf74Ek/KxNkz
uj4zR0KS4sI4BVw3BnNaCScQIUcEr/1sFO4+X2kU2aVHC1/i5AnIbeXlItRFOBRn89QKiNaGyz3E
htbjuhkSIwcDRWmwb+/FsmyqE3V+U4JGwUZgR3mq9MA/U8EFhBMLvQy3O7q6NnDucyt2Aqwf3Uax
yKX5lVdpscm6HO+zzU57kAlBKYwI/BW7LdlxaAoZym6P8BLSUM6AO+X0o7om9L7thsQiA9i3z1Fh
4w/oJRCILg3Umy5jhqRe1f566ekQCc14b98E64asuCfGfW78WpploiGA5uWN9Y8cUcouDFsMomKm
k19Ea+szc5XaMwLmDc2BXMxktXW4mqgn9veN9QgzAjQhmPQfXcp99/BN/NQz1gBbQch6FJz5R8T8
QrFUxxSSo0BqkGV/PE7fXBJZ4Z7TTwzjZF9WrD3p+YcrsrN9opYgyQGIDnEJPWRx1sxCw8HFz2ab
B0M3t+kCwi8BGetZQj0K2kuWe0IPdI6HjlPWZq+yvjHYNp5yADoeAgLB0bg975B/JJ1UEYawfSrY
uEwG9QQN3aw0iO+W4pqHKvVpl5NjvI0JgtM8zFX8lr90GqEHCvMBdwoSO6vqxWP4rl8/CIj2AiKl
Z4IrLUpgClb3vXnysRcXCGflp6DgxhxuT0VkW+yVOY0ebxV1R26C8sSSP1hit1FW+cp5M5IIq4gt
TZnaeHuZzoijS9mZI8tR3lLarInBnUx2vavNMErJAcqTxJkZw+sWTOye/wUQoxDEwXvm59xK/2uX
cf5PtyUrn3J5rXEeqtdHvtaga0h7CmDhDlCo8PTBd104dVft9uE43a4D6GCj6F9Y11hUTC0BGdtv
VHGcXWZl58dpJPMwXcJl6n2LQFVzQf0PtgbYm06/EFx9VST31SfO9F0Sh11qc8tlT6rk7Gnovxni
I/zWMUZHYJwU4FQT/KjZ4Evx3MG23RRA0toVfyhXn4qiP6juyJ7GARB5qlIhfq0PejyLVEdIL3C4
WwJ+BJ5/JCCXCRdvkoRWHU1AtVwBL/En8OACuJ7NBw1BJidoCypHKtasTdzYrink4lsWwHV7uhMM
+FiVNEFKeVXjW4zyX5U7lVxRTEOeKcFohCoUdIFq1Icg0eNdYORdj5wyihNb7efz3y2azmPVogcz
HwfgjREH32lziQ81T68wKAF/OIRhdLH0hRHIkHGJT7CgPeyg2zthHnSInTocQ8VfIhMVEHC7KKPe
e8K7e61RL3R9PgWNxS4yJLrpa51XV6cU9lFFkqstbwiR1XLNYRnHNrtsEWbjPp3aeXpxUCHyyDmP
FNasG9DQzaqn7yX9Hrhn1diV1V4upV/9zrBXoyPwsXxNFrbKH4p9sazzs3KdehOrvXQaLdxazCRC
BR4aqaH9U9QVC4nfW6Qc/rhJHMgLYKCHKbgQ6MYBZTpUyWf9ca40+ZMuI68S8SUDqw9Ws/cc10r/
Ymn3lfoxjnyhusKP2jAn0AeojW197W5sjCLmZTu7nOmN1Yb+A2Ov2il0Q8reVLT4Gke53KKiwpvU
vkvDl/ndDWA8WkICA5ydgrau3MFjUsLHWIkDfRcgB5N/E4KJ1G+VxCrZQa3iwD7gQIO1evHT7q23
x4Nn1la9PjGVNmmLIMn8jTU5UPqmCqUcDMX//i1/pwRwhE5o56OOLtQ7TAqMq0n7CXxUvJ2Np5CN
NyMtYL8/LhRpSadMXTMYADFCiNezGWsuq/EM3Gr8AC2MJrr5XzQ/+jeh0Fy+AYlg+2OdhQhw/h3G
jUj/rJ3D9+mYE9OAW0Arimk6zZhB3oXHVq5lj7VPhbvQksJep5rbQGsVrJMg6/QLf+Og/Xotjfuf
pgNfBEp/c4oNj+dafXvFiZCuAmoaaAOvi6O/8BvjzW8yPuKk1cnXwiI9Y/bk+1vwrdqNwl12tPHF
GT1a9EcXxZB+fN+jeavUglDxWFN+Y2bAeU0fWIIZwDc2Za5/iwwL6N96oHdAWqC2SXBPazlko57+
aDS1oxEDMVg/tFtLmhArE0BzilJreK8poRNqOwNP5YkQc+LJmI4yb59TqJleB4ZmMs2Gcqm1e21T
C1SODjFS1FE/3x8DeQu6dqZBu1qRcT77y6NTLjjF3ghlp4yJoyvvGrZU6hnbyNrdXMqxuJtWJliv
5Oe9VkkW29ZAHMIwXcl0hXpvC4QdZZx44473a+XPzSjrX04SfBOHI+CQfrojK1oTBQ4TTy8CBvUv
8eJd4biREelRUtoa6NCVozOjaquvW1VXVpIWy81UuTBeoIfkgGNIHcvKXMBaJV0+mbWqh29umW+P
IBang4z+GM2kh1ioxlDJRYF2aD/kTtj+bkeZk6KeBcpozMs7vgHO1cLjsFVbzZ3bsqfD2Rb+49I1
+Sl7c/GYEXz1NpKDx+SSIfFl+Xg/92jXqq48J9waHXXthEZdEZfv6TGNFxYJv+T/9Irv3r8KYeWT
UCLrKTMRC42e0CV2+u/1AxaFVOlaxzPCxV7qyePs4UOWzsEuIDmIPLv8u9f/HIhqqhDfnGc8VE9g
JPEhymqd6SrxiedLk8un2cX8ykULN2NN4EuPHIhqescLDWoWpSN11g6iW97rw8vyvF+KiIVodyEH
V1sxmF5QdEQTh8XfFfE8hx+C2YxxCCUVAHQeNbKPTFDR6RzwENN5NzXy9peEq7dA9KTBE2k+CDd7
MArkYyRFloPhcrO5KKrXsoWP6W4iyVrYc9IwUyUPvc4Nf8MIeBXyVpac4KYpYEUDWM1EBBc27RmI
1hEZ9A8DxdahDdhSiRbHdT42ujR+u8QC6V9kOeRAA44pDsgGs7EbmZFbvuYa/3/JV26gIEfO4QpB
0K20o5/Ejps1bTu/ftelI3YujE7YxNKlpBtKXW62LgJ7rfkCdEEwBBaMOAraQzO682651fmgso5n
nvFMaRBZ5KP87ev1DhCfDkl9Qh9HIhD6JCeZb3QsrQyzv/ySJiGMl1qAjegdCinEQS0iXXgGf//g
foZNj8h810ylBYYK2penOrZejv8zGJeaulmUTC8ALy2W6sKli8BR7bU9mW9cNE+Vb4bjRb5PS9E1
DT0GIjCIsK666dWLevVn3uxmdaI4eyJbYcieqbjC7+ROSauvcMdli9n1b2a+GWgyMO6o8aXRLPgZ
gPtswdiSV+lau320FnViPGV+7JeuhcXIO/YLHkxA0oqfTBqTPmkVgmIRWzDKFuW2ib7RJX6CdCdK
b0Lsw1HvnB4gredlkM9SqMkNCOgKcrSt+6qEVAvbm76ONweotfgiDrc+tSWpeWQUojcoNbP1ErWR
vfymMOSLspr7GXQmcDiDFiEE99xK05vPnTs4B5Nq0UHPDD68+Jg7XtZwBPhKIXm5nq+8xATkfjmk
VT/FVSPXxr7rD+6QMHyQ/o46XU87zSlIsaFeoREEE8Kbcxbb9BUzNyZy+hFmyujiWOV4Iz3SLLmF
paSNSmQsBrZ1H1JmLFR2Z70U6wv5op/GEbXin4WD1fOb1rEIM513VxAQ+tJBQM2wSV/ZK7Qm71NU
A6f4UL9m4EKkWI/pOk6vlgZVyXRUvQpB8EVSMxW6tl4sNQ1RmjZov0yjTzeJwOhnB7gvZ9ixcTh3
2C89gvpDHVFpWMTkRn23gfLJUVbyAs55cdudCMyZpvqPx/YlE+3G5s/n7CO8jgBGVmeQ/W7KWU89
6t7hEnxtY98BZyq5mJVUwMwDrqtw1O/8xCGOlubi5olikIllSseV6UPpB6stiBYP9JezBEtn9jg8
V+fgPdpaDPWpJ5tPomiU0pa8Z9fa+eqj7BQAMqlzaABW/LDnXtEdXKiqYkcIbuG3hKPs8bYJGGTC
yq2Wg84xeNh7kJc6+EdMkm3OcA0SZjSVn73xBBZ2rj18yAV64w4Hfuu2GO8N+HRaLhpkwe63HfA/
G+T2/Ezczt6xTdgJT+I9yASkrroqkj68YlybFYRYWZQ1x+fnzClqv5sQq/Oj/cs2l6tkw+LO7hsr
xMwTnFHHZcTYxU+pAfbKdGml6uK7tYiu/QxFqEWWGS77PWdnHipQSxbWqx5qFiHvaPh5JiHhd9Bx
oZibp/WMMt90UfO3de07FG3HN17A6vwmznMH/vQJovn4z5vaZeEZCPScYUSR0z/wpD/eTMzjmtt2
D+o8wBoS40xjrCgXOYkv+DktjFoPJ9JnUQgkAv7V1kP6ZnA9wk7p8A6kPwkZNuURzlsekkMvPpBd
pIzeKWoHJf1BhqkV/68mnpYyBxVkBjqXyiD99tNOeB02dxgMw62herxhAn3taNGI91EvCW2pTtbA
ofugzNNU1Gq54ysK/KFDu2WW4hXvtxSY0ScPZozRY2FpgfFlbPdWlWNbHHYEkW9377QGKw7pf7Qr
oknp20t8qhgWjMTk/KIKSRNXBuMAU47tVgnWKdrb3BomxGt7Ps3uZhImH26NpERRwjT+j6DbJN9n
pKk0qzMyfWNvbMdR9Aox3HJ6KTlMCo8DzDC6NtIEJ5fusR5jV0/70viJVqZLB+eQFAyVjYVm4Etx
1QdyKy4BWMjiQ3ahBlorCmkqHUXE6u5npILyaiN4vu8bSo0k4kLR4zl80FylTEVcOBVrZypfzg/I
Y9yG8dqSXLH7DVGbux8mMuGB2nfL6Nx3g1JROuCA8NPTK4BUa6fT3Yl7Wt5UYzn/jL4lWXi9VQSU
/Uv8a0uk27OpgP7PB36HuXK6neKNhqtqVFL9TagR0krNBWyoee+ogm1rIV1D6V2Q8bHmzAFgvFeL
cK/Jg1119KhyT1hcxMsfZNm36B3dnOmOF9v3lp+fr+rPxNpVCsVNqShKaRqApsxenFRkUs5YFhZd
7mBJ9Pg4wvjbdGbmUhgRkU/mU9fpPgE+MSjmwKAU7QT7tjR3RWNcUILgvZ/NvX/YxnRbspxpmUi6
4/N9knLyzXNpPoDT/+3vsdBlYLwoqbhZXy/zf8W2jVMH9X5ZFeFeW39VEMiQe8rQZi2JtrCG/Wv3
45f3pkcmyHpqIY1mJWaT21ch3FdmLewfuZxO9RDZhBB4bun4JmF06veYT5Q98KkgPP2reQdeSFkS
RwWbRnvydZLccA7cAW7rnnYm/11pqMDUSobE50atyUbTYFRWU2E50ahf12z89JF/Qi50YNRh/Egf
hwCZ67CysjzLlkZUg/eRQ6qliWBx1FChDpPPvnJ45P6wxOr785Rc3yMlIaPSssmeXQ7m8I8/mnGs
crIUos6hrnpMJ9umxWE5FFpNguRwAPW9yQww23YnMCKZtKMEHMo/HMvyMLRzcyS48ugbkpsfnwC3
mJRSPIG2C3JqJ0xWoZ1taNR9SqdjuZAPAx4NZPnie6W5BQzMGTKivITTJJc9IR8tw2Rix/FeuXpN
H7vlEooSWfIP9QUe2PUhtL71cA4hJuAmjELuJMbhEpxaXLKfhi4HXVBLdn63+LoQ0CyWLIPMRR8b
gCGGAfWNoPBHvyisFy8ZL6YXg8HHcjEySN8EWPnEcK3e9PMeZs381kyEvKU/XlxEShcJaz7xhXFn
UFomYh2P8iZfuox4CvMh/KQekpBqBjDdYZKf3+hEWn8/b8Sd9LMrnAhH+wkrkQm3d5wlHyBgEoJn
t8NR5M8mGMQ3P1VYNcXHN9qS9h35d5VksiVlR4LHuKVqQewwyASiE290GHWhRnBds46c0dCVSvtW
DE3+iZmT/m1Zk4CRz4qkqZTpw+Mxfb8Q16qhbuY8O6+J35+kymguwZUVTfbP0JNNQC2C86pTSbva
LMWh30haNZKd84xrQeRX9r3/TVxGwaVpyEdcwnIOEFF5ljEFtGxdZloj7hI9l2KONea0RFZ90dBv
bLRge97hDL6GbPyMsECUieVRc1uPx6/wPVChPNdubRLd/0V76E4MIlLm2Egy+wLykbq1usTXm/Gz
zFy3OUNArPZEMfrvlYNUYals6CqfajmP2uOQGAHh4plaslDevbu1zwmRnD2jDYhRtX1zI5xWVlto
SZfpIJ2Afpnkvk1mKXPotjhWhmnMmK6qDdu5QHYnMfMwvZuss/88LFMr+paDO+/brA+h7eb63ai1
v/kNyWbgjXtj3aTZkb3cuE0nVxnIGuzUSP9uFf14QRc+v/lE8t0n9JiqoUR8l5J9CFgNXBM3bQJ0
qz5YhJZRX+8Ms5ovWcCLswZFTCZcoWkiJIYIhMfzVEPuDqnzCPnpML5vcMkxIibEP4zpE6VQrkIX
a+ZhpHkQ/b7VDcrOsLsy/lw59q7G/vUsWQ4SG3qIXkeUS4dX204t/YaEBDufutMF8Az6rIviLzNN
jmJIs9OULGpZgP1GPd1mGBPGXtDuaVYoVIO1tn7Rx7n2cFT2NK+Chn6GNuMzj363OGS/Cqy1XQl2
YjaxM85UrzZrP03qE7QPe6aQQpdGNPppJmssJNS8kolDmTan1zKY/oAfkaYjLfW+5wOHq9GhnUna
59Rf7D6K6UBwhqBZmd6sDpu7ckEHwqYvFQLiHKAOnM/GuLhk9M1pVue19kZa69a+NukzDtFmRdXA
Y43c8M2VgT4BXw4tJTptGdi18UE4f5E2Gbe+zuNj+RYFpwrjC4P2cJ7EYbjmjvMVMsv3+zLAfbj1
clT4s2f2XGbLdXhKzD0z0/TAe8XETk6TtwTKE0P4bXiQ7P3KL57Lt7apo9jReDdB33dsuSgev/LY
JFINqk0GalxkdKKlhm0JFGCAPx0x0VOVngFKuFvmF/dHMg0CVw+xfndPHqhlVbJmJuqLR6JUIv25
dIzrFn+lUHA3ZZgjR03GKbbrzqo4cbBJViqhTUeYSGNcj0Ojvm7hNY2K3LXHtUPWqnjbS2JIm0S1
YVsBuHFi4aUZo/ze8Prs0Y2hf2Dy2P5Oxby0n2qqi7j7g0vPORFb1lOv5UsNqOhgLutNAswBmC+O
9blo0KIgo01JJ2NaBrX5/46tBP0+4eW9XOacgu6PY9r4METxTo5H+mVfkh/Fpi5UmLk9eRSNDP98
b/PwR5bmT+p9lDWh67lnWuO1p9MDu1PmsYVIo5eduF7PF1on8REc07647spd6zuIJ3s1JnYt/SbA
+8cETx1KGZMJ0I6RdZMGES9YFYbrmjnPir+r+qQC2tKvM36HTBzKCjlOpMoHro0kPvqPDAtk9jcw
R0fFi3uuPpuTYRD8CRsKvDYX2bct5ZUkqNoR2HQcG3A7r20g2M+h9HsHh7ZvHt8EQPticvsbNTQL
mJKhaM+2DHEDOEyLleMCtXI/5w+KXzw94Go2/ZA7jti7f+ydsxJgZGf54l5fExLP144Uqp48KZik
2mFTxPxzrsOs8tsvJZgk5JegkuOd/PgyiKfr4u5kuIAayu/v82HwsWGL3Gnu3/zqWIIjAgDTqZ0N
hRBK8pEX6ulj/YMzh3igMIfrH5PhiuzJaSJdQVgoJGl12uRR0JGDviSlGttCqj3zIjfZxtbEjPIC
eWN5Y4s0pCWuWngFSdFOB8Y0cCyKGvZ9wmnhETsVh9KliuzjD6yd5zLHBlMS/6ldf23Fg6Zi5P7z
RC8iALRkGBYmztD6xHAjkidR3s4DZYA12X72QT9vcnheC5hcCRgnPVAJDLp3qTzVPujO8lOTq2Hk
395bS87fSZCqHGYo42yeB2xxlg1m0T2NabbeUWEeJYPzDJl/uwxT5Cvi+ULb8nBiDDAppwLsQ9Cq
0GRFfwvlNi0Jf+6rB92xkM1zlbf7kNMz9rzcccb/OAs53+Kqnh0y6JhA6Ouiob7efZaA5ve2D5Sl
15Ex4vdGr69hyxCH8DcTn4psxvVJT4mrvjfqZb7xhSHEZF/rFgqOMa28cRcKmuDvgGZfc8ExbXev
v8BOIvMl81YQRVidmfux/9/d7p9gFntHhD43LXyKbF+Yved2mZDtgbWhZsJQT2/XfbaWlUOUOO3y
Xguyk9oP4pH+/lXPWIBjKKf8WYjqmLGiT09mzNP1FR0JpAr4XNNLa15Lh7VTERxJ31QS/258aWUc
RuIZrMgzxQAnrgtqZnTqGyvadMW5LPjRaBRJgVhW9Y7pp4jL+LxJU7+NkhJZ9kINbOo17/lGP2yx
zEBruL/uD6QiYMKJVfvQXBcHQeDlpDtpFG1u0YlpdcO9sNoZNL1QqGG35hARYKZK+UBRTQo4MLGI
Ydp2yTkNh9iaV0MB+Sb9YxtTpAYyReawNzuP4mP0wUhG6r7JOAy7xZBRvHjRGiJPHF7L1002c+W5
wxk1A5II4lAKovsAvc3BP+1keWi7W5GqubeT/qW+z218cC6VJtUDu/fX8vnp0HAzZFOpylY+7m6X
BC3Kuc55pYi1gluq9qbB6BUVS/NjY+o5onDWDwA3Xb4ME5K/Db28epcuqHdyfaJaDo/BmmkyV/0j
dKIbcV8+RvQGjTxa1tf/bp/HtT8ZcC8bZSbucB5dnhggSY6HlRNBq63qnsL7vhbvj0nIOoqbgRZg
3K/ysS/W2r+J5Ycu919M/PyWm7LFw8BdCVwrGNWPWYOigqMScc1nwuxjOBLBp6kK6gtLgdbM+38f
B/7Z8OXsTFd8TlTC5tiSui3qgh4tUKzoVVjUCKjYG1lzTMju1pUhxnEyAhyt/S5gl7vtAGA7l3ng
m+zVbGfBjDWevhIq0l3nN7sBEzxWhpVLfPiHsfTlkKncHUvkMFsSO2ijQdcKA1dC68L4IY3rM8+Y
zLLSkd6c3/o+RDimysZb9g9A89Erk4++SdILPyrAML4SHlr0XF+6ozkazIP+lAH0Aofb8qg2e5st
T2cUKot6mPAXLuvppzXz51yXso/v1YRw97cZhPVHfZNUanIVXHNCqB7MzmOrnnFLBAuBpeDrAAjp
Fx7PceQODvv9ApFXT+JIMj/gqQ+tJbiWurVXrOfsW6gGQqhVsSMNAWIkyyxpSgo99NCenZ6SLeC7
vRPMkAtUbZ0BebVrzLsA8RSfX8x3fuRg5TuA3hTKvLv+Q+BZvftkHcXkwNand8ryBrN40Ih3DSyw
IYviyDZgOEIpm9JC8RasC/gwBd4IP0yllEd99jzgrlXytu7esPg22QKeF1rdFnREurr5CQtvBRA2
TV56EHShj0ftrOe+W87m4BuHAHOmTahr4bTwkyd1QNI86Lcm7YKYi3yfN121+t3zZn5uQ99J7T/2
CvHqf6BzPDtHJZ4Is6nxs+QZ2DXtXOKw9KZ056TvstxLVGWV2uSlZuLWyUxvgNHHYeDP82P91Y+E
ffsJ+clJRldDPMbOZvIkyL3ZC1sj3Okh0HIKG4h91reozyomEgv6tMTBb4/7xemr2ZS8x3rAVqhS
Hs/JUE+lD1kyaCTU1+6pCEX2mA7Fg/+SaRfET/efLQjTqSEYW7MueHi+iPAIq+FjErv6U+zGU7HY
AX6PKcSGIPUixsYISQYKzABmeOTboDbF9AtoHYPYMAbVMS44rwAyRGKA3nXNZD+5enTImPjaR5gE
jJRTeJRlyi5mCOX/p9pQ39QQAOL8Ul9tVAot3YTy2+zvRvNFWFDKYgzSq0JD4GkvlN/XeNOrX7Ki
epA+ARUS00ri6PQY+J4LTteDFSIXrxlvksGEBvkaD5Wiuej/kzHb+nxfpMXw1V8sHHKV0nzRYPLr
/+bkxga5dp7evVcoZyNiRU5uHZ0OgHUbkXjWTkLsW+mMF7gmhrsNcsWjh3koZZJUSWhQ1eiQGFmd
xUm20bsnkeSafcdgVBdos3viELagokfqx0u3BVF58UpRiu3y0LV0IUB/Bg2lOj4RNWnFC9Od6UpA
xepiw2v28tflmVJb0dTUvzQKLkh9fBUUBuD1U/x7EK8Zp6JfGvY3gjRAW6Wh9LW5MwGsTGqE3FHG
MBUqlhpLTRYeywkB7x7FxgNm4INEZkrZIQM/eQfCpFfRaCMnHKwHMTi9rNsJOKBcFyQlhJSnOiN5
HK60h/sjBLRaqU6XMiFw67w3DgHS3AmMqPFXQAImC188EN0T7OBBBJF6yDIG+BK29daj01/q357S
slOSZ89jUgq9QqDdm477pcaFc/QTiEdhVe2WMzOVV7XT206QdoApL3125pWKofQMwXUmZ1aNvHkN
uRwrhq5LJfLb3AMslqiH/nEOA1z6v5SWjlBXjLDfiaKMBnYUpMTWAfeQDNXGKl+R2cHVZ35vDjjk
J7nQ1Vr9vLISrypcfjG4R+cb7ZRHpHyDx7V+oV+UtRPMB+qJRM1EsSf88GK5L2tz31H30iLVy0pu
2j59ZoUOVJOu4z8FeOxIYTvFpKAGhWT/OVzN9Ms9qvN4RTxEvbqggTXTiFakRMfBUkO7Se7xQV4D
BcchWTdZWZUGcECKDQOKSQQa+oJcCp0YtXOahYQw+ZPaYQKcPxUn9opsKy0+At8710aH6iva3NL/
i3I+RpN3fb+5Vj+8QX6CSpKurVDSNfSqn2aQUCuBQOHsHkG61jNsserKLmsvP7hdJdCNrimS4H8N
k4ubsTdVqeVlEXcE9/iinwmWuVHgA6j9ZW6Kk+A/jgPwkWmRKZ9zAmIydcsvtg7ay6jVo2sr/OYh
gFf4k2ZQGAys+Q+Ve/wQn5Cp+klxuWaq7W4Way/GYI02Xj82hXUDPCefkWus1zJk2xfaml1D25bK
lEE21GrptTitLzbKwmOeNfw9QKoo23q7+DvipDPzG+Ml+QNeZvqiWykwU4D9n1mO4F06Pw78+1Wr
OjSFWTpwGrwLevE5zHSl45UjJLp1pd0GHo4L6DLngbjdxBFXhXEHxfeE6HNfPjffEC1HOPJNb220
Gd+FnDHMt3I+ndTGgOlBb2Gvr94xKPQdRtT9xLPE0utDCdKQShYkmGmnIyN+Rj4uJn7dLNdlroC1
hQz2qxnZp+JjFSUWlRO2/JYWuts3wW85bEYhNCYg+q5VOeX38n6FWynuHiHBJT/vOwbyqWr1PHNs
Az0Zt7m7ph5IWokJr0XqcRrZn+s1XK5vBiPaP+Vpg93ZdXi+rPtTtma6Yj4gXnulfCN/eYkxNAmd
2ZS8Gqv6Gj8nrkR0mWvIkMsmAbxw3ppInS5YtJrSpTUGclh1ylwKJsNxx+n/XOkykmU4MdUVoX7w
+fadSFE1XkN43WImL3XC23WlVLZoaON39wAiUQMNc232kkPN4OSAUt1htzGZBHuR6De9zdZEVP5n
hNS0Ss0clmFLxj1dzssxk2GIgR7O0WIR0QFaWo8W0xNCQPg8RdXIDDlGcHJBz1GZ+7UAZJXbNWme
8N3xV3MuhY+oVDjoZg3ApyPs+socVkoQi1q3ytn2XpgsQB5C/3P3Vx8MV3S3fOTfFDCFwD0QY2zj
nLSQp+gWmESnteoj0fybqBmMpD2VPbZpT+0mirve+oAeWkYqtuFspzUJHGCgOl3LAfT4g6y8hzKm
zjeTAhDmTYlv/GKe21/1vaIZxRpDvYLaPNEF1dclwU9R7m6qI5SQxqqMAjc3bSxRg3WCYulCeQcf
7efbEX5209DzfuW/15jESQrQEcHG5rn2lRdgYlWGgV7brjdBfbdRpF1WTJbX2Eo3g0wEuANLGy/5
JCtMtFlArG1ruWIPCMQH5meRmuVNnvs6sM4HkcuvYXnmwUHb8dPFkGALJTp3m+HEiju3em/MPweD
R28+L3ujLsgwtCh/CYQedyjIkRWiWym7sE3HvoI7sXfC4T3V+t0bv3CdpBGb9DVLNJTAEm6I6ouB
BdOWhLGKalyY5s/k1ySW0gmRSgamzXbbrwX3+KzsetWPvS6tE45HN2CSFVuILxeE/bPZsWBoNHy9
scixmvfzzAZu0PA+OLQgmtA03T2w+rWhQHAfI/ZT42YOH4Hh+BVNBfSmRhmXndhHDlRlyiQNL2Cs
VCEwG3BqY0OWwDlgJcLcECDi40x78iawcAN7oJzYN+RlqNE2B0ZvUEUDnLbN0x47IlXV4ZnLVuaY
cGVYyG2s1urza7wFgmd17tktvdHDN02KaS+qWPs8QvZQy8b8jGCKOsAj5rqXbapQE3pGnadAFsaQ
mLUXs9E96maAmpes3EBswzqxiloDUDzxehvRFhVDe7v+fNofe5/Sa7JdfjCWYzQV12FNw1u/jNqd
iMsjP9kBsSQOZ9OskN6C2dp0ZVHIcBiz4eiWEOG6pTnXpxRC7mZrWeGj81dEgYPd8s9ay5hUZHN5
Lhdp/herEX3wniCfUW8YBDww2UlbnIU545Tfdhc9mZvqXnxMYP18PcGtGa/OJNUhSOvKpmlpPnUk
NDT1c3VQkvH2/9KeKrlwOFC88y4z1Qc5TKGC3y6OuR1c9feZ70tdteLpXYyMWyO/erxT2HITYpZ5
T1+aHEoD9n7LRuKJ4jy4DQ31FmgRKIGuULzQhB/RmTj2IvDnXXKfr4kmYyAsOv0UyA4kmcICQwK1
KsvMvf/BTsp5scWshkNib/6RMGo5sXJV3bxS68x6fGJC7JRYp5S0PKAYptu6gPvNSDCuPhoo8D2p
LZAmmRl/UpNss1SntXnotcmA77WCj6k0TPNSwEILxWaheo53m1LJJs3mOGLv7sz66fJEDJMcStal
S5crFMBpumrEljwSkLAVPXdFcOS4/Ulk0aoVhSf9OfoeaRjBA2XYW6N4U3bDsaragauFeGGaPhhX
h4VAqNWflCUmiLitPAz4Vb6+d1/OVuU+urnkp4Ub0cIJPZvc66MlVphI1BbpHZTpMm0frVC8ui7r
vuqTSh6pdMFsaNVRYkqqI8OgYJQfXSQDvLjYBcdmGRDI67oYWxaYL73su7hQIiEtr5F8Fz4XG+F1
QkUtm2uThLvsxPNL30/IePqXirsk5VmRyM14SOkuP/Pcm9+a/HqdFHARGmw+YGigv9sdBDkf1CdK
llFPCbf/TB5vY4XgA6OsDLtFHi+wM3p22vtfe08nBc8ruTSgu9Kzz/XQrY++BvBR0w1zcQsWjwAx
H+7Me25/I5Gm8+56ZpQXt2PWsd5icFXAoYjPXGlLk7yuM4mQebV0fcDTCznFKHhq/22TFtJBczL5
J2Vg2ARNGuC47pF/o8RRiYlkThKIZoKy8wwdqJ6tw5sFy5arW61eQu8ycVDuDucZLIFYrptUVzvU
ymzj8UbGq/MkQEDL16Sdu4BbcyboXmTHTRajOrJKvcHdO3WvTLmhfCvTY40bw8UKrj5dbDmmVxwt
Iw1aUTZhLlv++qZDNhTdZkn7jNg1SMSYbiVx+DOaRphPhflYEQbFjtWRwsgIX6xPIRHgwK5GYCC1
QiLXUJ+KH+InIhrh3qydR2AaoGlXAIv5gzJ1mRcPy0dfKqKslQQwAR3kAiEHl20ZROE/NIyejojq
uYJA7WKGgdY6AmO3XX/PUegknaI78NDYaOAW4Dq0Soc5GAUglbcmdJRJG7WX3TgcgFiihLFv/gkC
23Y4ea3eRUzgv4/2pMHW7W6cY+hkQ+6qEnXFqJjQClkoZndmi9Ycjflbwl161cRhdZ1muXPKNxC7
FCBD3lKjHQi78mRVofKGfIVVj8MBM8aUsgRGnRROKMlvcUOvqbiyEgT+r3wAfY2JnLwldhvECFET
yiI+kyjE04t2kaioT6ozvHi5YMp39/MetD5sGgD4oTUrU7or3MYrZkxLVhuOSV3qH5vE8CDvnyw8
9qfpA4I/YMh/hfHGTvMRExSAGI3E7707gxXp6pASXPpw8RqRGcVdpFVO143vjQRlUi+ew57xEEpX
ViOVjELfWI8At2nsSptuy3HVhxk1kCK5ln4d6IrMV0VlYJRyoC7Jiy7yytSY6BlRdKgW6fUzlE92
eCl7QDAbtIkw4qI0Ly20SUHtbqJWF8WofL2IzBii3hKtK+UDXMeHiE6/Ptq6LakzvEwsSGOnhheu
AWPoJjrwcOLraJzoIi0ArGLqbeqQzVC3kBOSrMu4ILMbFee8WLHEY1L7xGS1Gx0KI6sJL8Nex3R4
NeifHtlGZA4oBQj50z3GMfY+Y9Ol3+U7ZqBCDwc8SrieHXV8JzMu7efzQZ87iRPyUL/WM4yWc533
TTIq91EHn1ST2qmugwdCL6CcFWczzfVgt6P66iSDZSaHRZOGPwP9hIMTcWGFx2ms2gRKYDQQDZUx
oGFfTvMcYHwpi1LxXGmF36mlbHTAciJ/pe8b0OoAZkgkQ+VuTXHtIvFcnz7gqIt1R2l1rReqVJ8l
rX8JYqaj3wMoaj+35BhMC/BGaMJvNNOPGiGQrDWcxQRRyFXEeGWWooRyv58bWVGV7nUTpQruNySm
qVtsRx//9u6EoVj/Evbem8FyiDQ00nhi7zRxTxjDMJP94dw1tnus7dKyzyQx90fQkCLE8NxAz6IB
OpaDQ3raiMoBlEe650fS8oJ8f8BCb7cWnXBxuUmuN7yCJdjYGCW8M74j37tZbNiMvD6tHeWxcM83
DgTOYRY50ZzMuRwtaEZqzYPBlIrZ6NVYrUSdbuZT+ugkAHXcHd9UiF18lp2/IDy6W4Zedjflga9Q
t6nIge8mA5oDaM1mZqnaQQc63Cb0FiwWDj3tGAx4oQyQguZpG1xG8gmnql4j1OXM03424fX74/eJ
XfRT/hmgFEgA3qGEuVLSjJHNss923dx4Mg3VaQjN3XckK10NNQrB2es4eN9zH73FdDM7g7dy9IKa
kiKQEUEWzwYoeqfHlXsBCJLR/E1iZxQQ9r86w1dylAzuV40Vde3NFO220dQAYJ4t/4HtFExDw6v8
xECiAUG23THKLJLlf/5KGaK1YpWgsJYoW/PRogd84oh6MjrvCgaYkomrucAGfOkjs8y+9s9KIG+O
/c9/By6COxy/uuAFmaGvaPE2QGhwhHZv7tQSNurBWbm72Ou14dMcUiHfptVW39xPbgmkMd1KIZ73
y5gkA9vlbs/XWzL5GeFprLg+xZQEyif6Mqbg1M1NA4cs/TcRhtLacQrrySWdprKYSe7ovDHI5akH
tHe4TGC3ZRRTp6MaQODYVkUu5caAkOHCK6Wz7+TP3Cmdr0KkJUfEab+IU9x9YtsaEsmVXS6wQE7R
Sq4vP0NYvycjmCy7kYWhAYgbgACjXzps9nYpzshVElZq2Q1W7iTvYWAtWqBRkNwSI/T1lxaKvi8t
IKCxDYood8+ZENkH2OMYQ/GYzn8+w2PMcr9ER4I16dPUFF6jaUS4Qq5rjmBo/AJnGYlfj5qsEljm
2V2cSgUJH4Xrjo/HF7GtN81MjottjEhQ4t6Y7rnAtWpyQePvJe0apcE4rNi7K8eQ9qvRxVgbN66W
wOQNCFCd9Eys6W06Bb1REWM5NvGvdB/F3qstb8sDgpg6AutIg1BfnXrY5HhL4S8sx2J/nRYvFLzS
pNXny3JkRZByf1FhUJJYj1/7YDDjh2bXuAg2h655p05epMv5jZknq69AfCkSwv6f4umRQmXlQkUd
pAFYfp2P2Si4HvhTSGIVQgiq/vVQqhqSQ+JGPUVNpiJHpFVfZx/l/XC6OAy2IBfGp2pULgkUHtws
X0cLkk27zv64Rfu3uO96UfxJ6+HRfI7Y3dqCVserMmBYgVEBWfMZJXxNI7G17976DJvdk1c1f3ro
LXUPZYPdAuAKjClLKMfjAc1A9CpOfEzlVpPo7QunqxViY8ObRllo2ccMQheFjvgYlYi2lxuoPMMu
XlcQ9I9dCITF/qE7cTA3RfPSsDkEOOZyKIDLVaHVCFTW+kCtDo40+aP8BvUOrebmkUMWIAAPW2a/
avxfQW9gN32rgnRFzZ8DdoEw6RaSOBR/e2CNyN2FjIvGOcIF25uBLACX6v3tENHhTqHL2o5ZqHRU
jvaL2owMl7WIoOANunRUYzP5hf1gWVrvwKVSzl0oGHS6Rdz5hunoT2xFBqPzIhRRXkFHTSa2hDFR
2QZiHKB1OFUx5mKKWXaHawvbIYrGqhLBmdIac59QCBYO02BC0Aphm9oDrPYs0ZpkriNxRQEiFLtG
TFljA30qv3LRf6exsVGLxuf2NpngpanEY92SYY92sH8TKZ3u3BrLSmc9dISF3L0zpxv5mFF/vlQj
IngHC9KKAR7Tj5mkLWOK7MOTcnCu9Y3yvln26CqXXohsFdkEfHkcM48G0shsEMxj2UeR6/9CCp3C
jT+PnLtX/eBaWlPH/y5F3b+6jgd86o6svqF6hGxkB2hgCTcB6mjEiN16q1lt+g/DUQHlsOmk/qA2
YZ1UXwmHzPdVFT0e72RPcrINikutZIuJP1kpKtEIlUng9eWfmAoeZXrG3IcVdoytQRBpP7h2C3IT
AP/W8dGGW9wy575mIMtQ5TK4a4HjNVOd44/bYfEvAOtb4h3OQrYa8oolpxJuSjiX+/w399Oc6cc3
13eUorgQcW6FCoS0n16nb8CyeNY5PNAvVNYqQOzst4M111W5OROp1uEZDGWndA9qpGxO8JhIF711
hgB0DH6iUxoLHS+v+SoFO9iC+Xv38dquUhQpOeg5ZHxsPFBjUpNmZUpwN8Y874he6ehkFg2QomKd
pDI6sQU0XgUcRBOtYnMS/lUQbCSuR4TaQDdx6p1yeBs3IBAYEnaEVVCmaM7p2P7sUyvYhPg5UpY0
5QbMoXqpKw5CASoBpjuTqCtSwQ/EZkOjyFMexabejhA1STpIH+ZbHb7bexoHZO3rGQNyxQj4RW08
bl1heRmHgzHRn1843ljP5Kedlx0fJ0DqnwsCIrhHC5hz/j+ARYNJ6AbIgDtxnsSMSm8fdTyCGKsS
IbuHPMzrkr0cuZtx8MXhqAaNX/o5CbEZDIttDN7EvJoqthvCA/ubGnhm2oM+WENYqKVUlteTYMPi
VVIq0KelBVNuaW4pEPTBOLA+ySOmF0uawce20Fe3J3/FBGDgMFQUjxL4ZgWDzgKThrcSHXKFEN6L
yKiAjSESOKOxzV2+YJuFv6LPrcvsuzXRiKc0QlZ1TwJk8hge+cOvCNp2EF6kRJMzS1ZLNX0SpZcj
7/dwtXSW6qen/0ZCBzhg+R4genVHsRI0sI9s4T3HbwXpOHlbojmUsrRp2DUCi/iotUBr3YuKnuHZ
4drXkcbYZvvKU1fYpiN5TdyAuUUCS2I9HHk1z13Ia3HA4nMseRa5y7v3/VYKdyHYpgLebCK8kQQG
ak0RkFTG3VuFk3jlDI5b93Xjh+R+5zX7hWtORs//rOnbwF1dKFTHNUGRVVYrRiBA/yHgINkFb+Di
ElzEtUbuhXeiKtUZhn7LKIQiubk/gplT4mZ1B5iUdDLXZ2T7YCbLDFbsLgfB5PYtf+HAzsI2HR4D
PVh79K3ixb0lawALTnmhXJ1cwLsfDM6mJPWIUCbbyBse2/mjurBIu3P50GqwZYnjNMOH7FI/iGn5
Q8aHcwzV7pdMNHBnHGzAc++asMsgPNxFBm0MVhkYcdj3MvJXkf6ZdxtKpODGZXqVXKzdiyNKMB+I
ROlpEsKxUFTzk47OyrygqHoug+8NBzhh/y0gfCVIOUv+Nh8NRmrJbaBO9u62Aq98ZWOarj4k8Q3D
xfrvv9udfM5/bIVGHTBkw8Eun9uc51x3P0kiFoPnOrxaSj9KkhHXy9jhy8pRjpWaPf7E0hXYFXos
bQ6SQc0aHpv626dnvqeJd2JCrLjHfXBubVVxMZ24FCpqyKnEXKCOlkv6R9uygJT6xLrFQZPcNo03
8zi+uZ8/Nfdduw6ck3F56akwnpfzR3QHDboMlQlyE2WT+yjk6Pm/YGUGVOY1BThLp5z4eZopLN9y
EvercqGIN+vs7Zw/ihzSS1Z/T/DG6DgD0ohVVdU8mipKVGiogvs//k1hAiuoG326nMTc72nI9Lxi
BTY+LtffsSOUKerR200Kr/9AkW24EcfW28zi7GTDH+jHwx9NQcI5M++l8uIvpL4r883kzeV2nEEX
u+W082G9C95Z0GI99zwuHGTG6We6a9B4jzrz1qE4BtLTv3aSTspeGtZk0twZEEUf9S4TtF9W9j/H
vlMo+QzJr6uDckD7OO8kgULWrt8X0Vg93cV7GP0fqbACeqo4GoGqVS+AFxi+Gi5y/I+/cbR/7R7/
uSF/ZWgSKAqEbpR81BS0LbBqFz8tfeESEgH2yBjJTdntB5rhs4zDdTxkGIvjqS8jAT4Jg4QUAx+P
PG0br+YrbSgMVtmWjG9sC23oXJVK6a/MgnV2gp+aumuq0a6I/ydD9/qB2/OUTt/0g2dHLcdPgAcx
XjVyMSrOfULpS69oo4KVo2gwnh5MVs+PIXhERT4KnAic+b1ltzqb5yDjZq5LCSDU4IH1osaE+B0C
Oglw9uTib1eidL80PTQRU3p1S1ZXb6GT1Ddm6aZHAbgmGHWq4gTQGzqostJeeGA+xrJjQ6oK+4ip
uz9kthalBvrzGv1hqMjA0WET4Rs3b4Wr2iFJmekDyx9/L7ciQJDp31mc+54g6kyyZf3HYPggPM22
yL1xHBit0dWElSBh0RArjAENL/rLzMCJBL6k1/cK3lt3U0gTeE9/57q4nWcMGLh72w0daW7/aJAZ
deoPOx2Jt1UrqWB6NOA/fJbedROxuv7gji0e6cgd/P/mCC4cCPKry+lpIOYpPtPDWteBXaWT+6yf
OKWtQmYOrcK66z+zXYwFTcGTT3k0kQSvWMZVsl2MCBL0wA/c1f49415NPQLLh4z5soE0vUtcJ8kw
bwY/eta7WyDLk6KgvBoXmBrc2sD4SebvqQdz+1kRBFAW78+BnrhEwjSzNH5K8wsKFDw5hL5iTKvL
NiPMF+mQWvEa2DetZ+34947QvhjB0a5MWHPq6IJITywIEGg4eJoCmCAnTd0jBB6U3cvCOC+hi3Xq
8GyiL98vCAkbwh1fYl/KZ37+9jDNunN0uWhQv4EpVIFWu3plLCzz4GdiCDsYp3C9Gh7iKg03Of/D
GXYOyw4US258MDVDww27I5Uk4b2WpkjUe3ClODUi1o+wuV29avkGKZsvibMyAh/0Xs78OjkzGfBT
AitulqYLeL/Xf64zO5x1sUaiTbL+9NmAWY3bpQhUWDUtxOBVWQzB0L+7cGySfiad8oBey/ddn5Oa
7lAdjFox2+zsoQytNqEgwitmZnnO2Zeg/dpI8g2asA48357fri4Hz9xIwSNiX9WIjHqolp+78q14
d3TeDI7uniwqOMpQmlkxrziJ9q2zdGbTokhypfSSOIe3NhRG4DoAVvj4p+HshuCA9XcEBSoxiEdF
MrjtdfD588gR/HfPchR4e1wfN4INLiqkoZz+OdIzPBFtXcdHznbA6MfdstmZB3R4Zj3lFilBkR6G
iJZZ+aAeT2AlUDOIm6+dyjUX0FXhY+L1pUVmcJTJac5+JqHxbPWjCL+Zn97Tk6S9/uao2Sdh7CK5
l0NOjKhL3FwLeVFCdbHhKA1MhYdGQ7qwFyWAp+LoPBweRTQR1X0BrIepjcjIRHL+m/4l3gAI9gtR
GKTMgKsDIIkGblbGREiwMCp8p5sPjQL/zKCq1AAr/W3Envpj48Dgc/ORBiIiSS9q//7eZ4PLb43P
5nN1qOvN720mkWPJDJbY2dKgMVY8x7ZtsTr8HUImSZOLXo5DAdlonMxgNJwES3N49mT1zQmxRtd+
GDWxPsZNtt1zvjQ8R548qDQuFi9OtyWSyTv1gyOj+eNeinza+kiJo9tw9gbck6Bg3g9eYZ3OcbGD
7xbmrLvyIF7/jhIN9ZHTVECF2Th289DOsD1vSFtg75lsEylf9Rbwpc2Fp7dhSC+LD21bcNybQ3Bj
E7+UcFa2RAPiwSsETx/wbW1ht3mga5dQKJ19m3i+imN8yYt0RnjBqm+/Zq43kKOqnoWAeaBN4jmN
d1Gv68WizkOImTaWbqoKQnWMsZutfOBHJqwPSTUi0aCD6o/lWyAUtMUc99JSp5j2naLFpRkJ+Tf/
t7OKhykRw6RyXk3FxIK88Cq3Qe+Y9CUwZkAVz6pXqVbhk4jyEHtOP86chzW66VjEGBab95Os3RCz
/JheHg98afnczFLOHepO/MAxBDac/oFWcih1UBTEtZONTUBRoSEB5EhQ/Ho/pbO8Qk2JS1fWBqxG
W2WweiNsEupKGxW0KE63lEIVZR+rwgkT4WYFfjDWy50xSRs4mCdttvNCzXlN5MoQlS0vZ45iAL6T
e2LtiVVj6zlcTEgisG6WKAsI3j75OVOLAM55M//CehWZCbaFuy0/zgGKpJauCXBLxI5RVv/DhNa/
tcEI5r6ePD0erbD8sXWaY3ME3JI3Zhg6cOeH2BB+0XHuVLQwYBbcQbeBdUrLDY1lh6QhHNsR2GYr
x9aANqV042rtlWnuQz7WOGtz7Aj9o5whX/eCfD7cReweSXq6+GazGTaH+xrgcpaGbraqzbQHhIG2
7AfR0P+BMaU9ZgyuosKgGLnuXVWY2wfNITjuILpPmiGkCUoyeLA2rX6cS+wYh1KyKu3bIVfILFm9
yuN3kg0QYnPfuaIgsMX0ETZfVtQqDDljxL2//GVzGS6NUN88OdGH5VEm8qcDrWE++vFqoF1RB8l0
55Arv12aRJtREBfX6ckElHVgXM1cuhEIMyjI1wCGXmYL8UGujRkQlNwGlEcw8ZEv0HYDjs5SeCQd
XX4xG7YGdwgNggVMc3NkoWEQYdLU0HUbiZd8lPfDnK1naYhcjuTLpjV91aqthcGnsniKO8bwB4vZ
iTw18JS/clnMuJdbdwi+RC2v0h3vjECctTfEBuhsgIwqf6lkaCmAgp6ki9jvrGfF1esE1e/36M//
Yf33t2q8i0+OaPUmhnw/iRzrWXSDf6gEsvhlYxnR1kfDz/+Cl0xuTPrjCvpRPWy9eRcQ1hYE92aC
yXS/sZcrlkiL//iY+CRm4kB3zeoa1k0FZUg+pjc+TuqUzZdCbyqqij927C6+Ip5Nw6Go7ncLUBL7
bTsDg6PDmjkUwbrw6H0+k0+ohnV9g+BymSpzKgXsEyvLd+8a61fyjRL0d+9QdHRmcvOglNXfQSoV
kyIXwlcNkHEwNLcFhzbFfuJvhICjbOP7CZtzg+/5Q9oIo6VjWJOeNscSLx23kOB0/nA1DTaWzh04
Ke/X4JueBpzN5JqiWmA0XDSLDEK3wFTmGkmrfWStQHdfhe3GTVXhi1EKsKruVKHpSNpH+EOZC6PU
OrFjdlujL7v1TEthkne2h7vNzRZC5ocbbCIeRJ6j7JWrmTXOrLYB704g3itWU/CB1xsLLCQqh7wO
pyz/30S10lfYcgiI12FJfbJ07iErJD3sda9Q/GaY1hFDb6wg5316LgApeHZmm6F665l6+Z+hopMM
5BuchGq3y1i/wWnSl0t3/jN0Xx4dDJaQacekGgndcJ1d/bGgrHx9p1qzFyL+NxAA0bwJwL3ZPvBQ
FDj18jno1XjJ+ONjLxq6phK8bBWIQNOSK8+f6JeF6CpFM0hIVq0VwdIQWutu1Cf+3jsugnHbepgQ
0SMIi8U1dY8Mi7R7PtEZU1yW6aiZwTV9OPFzL+eBdKehaeyrZ0BKGziz2yRCGDGwAEFCjiARcWbk
GMGssRp5u5LY26D/G9W7ZBTNxzu9vTZXTVVCaLq/UuGd9nP+hGrvqhTRn6Xgz0FAEd6vMqll4W3U
oc8nk6xiD/1UNSwqKSuaS6KzXRdVc0zOu6oVgvyz6l3TUGnCqlY3UmO9aKbFO6bx21pMXtpc2h1e
UuGvTE/kLrkQPIVejERQOejqtKxrSvagQmREZjqOEVVFl8rRa3VY6EU+1UNcRlXgv+DlvJJexQXz
yRI7QB0Hq9dFpca+gfhKhgI5G3bZDpWgD7ZRbaHGCAe24J7OObQhxVQtaDz3biRTlU0VsGrPaFtR
2kp/6cnLkXfQ9glvcKiDVUoot0RgHK3/6hDoZB4fJphbhs4RG07JvA8=
`protect end_protected
