`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
bDP+bwhoc2zQziwQIbuqbWOZvAWh1Sc8QFH77MKOS2DBwUC/0WcE+Z0328m0Qs4go/4qUF5lxpeq
9z6fMsubqeCFS63wLnjECpwsPSdmSaqHvCPEn09fvlDOfgCLT9SlFNRsFzyIl3oznsRa8oc5QRgO
3CZvvEuJLHk2Lx8xiuAGPl2UWcew6rAmRHRiDoOhsZyaXmjowNEdrp+PHVZAhclRvgvdWWfStSJ8
GyjCWnnk2WO1PEqQvK/LTwISZpKKJw5Sq4B7nTphxbWI6C2nODMTLFa3MQqlKAiofwZZb15mQthk
NtSlInJiwJDfgQJqD2IrCyVflWjmN9NMcNUhXw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="g8mccbz8BICdsG48KNAeJ3UfEEba4Xq4N0U6uBK5N3c="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17568)
`protect data_block
0P8QRSbiEStK5lol5VKqIClorPQI+HYTiZJbl5UBoZx18qTJgios/HqoMLCkmpO5JsJlEQQr/GbN
UbkpFM/1ENvZdMqeFErveYwQ0c7m5seKIm5Z/TWwKOynXWm7vFw2kxTIl7pMhetVBzirUrIE/yd6
BFMw6T47il/v7ZFHDq6E0G057a92MJoWQOZ8T2OxUGvm1SCgMAh+H0VNKlHToZsY3iG7JB4UvDfj
MfbcTOFqv5GwM/dLyjVpEMbYa2+OIrhxkEf2ddrORwCrJ2C+3+yJjp6Tml7BPiABa65dDhX3PkRM
EgcPRe7wejI309VycyFACu3JYsgt5pOROBdqDTGHigE3WMTNqYgq2+2If8IGgId+V7HIQDCpzm/q
eyN6iWxvWc5ajlHQHjfdaNtPzglXXDRtK4nzNbWPtAUOCrF9R3rEHHfYfzkA5ENk3QqIGd5qRGnT
Ed6FcAMSsa57L0r/lJ3X7HpKiDEkkPrILirvCIRe6VQ54QRyEhTlDoaHKnfshlI2PRqjVWA8IRFP
rmYhXFEdPnfqFJQstcLO8bT8oh9xCsBv5ufDT9P4oWkGLYDb0RnR5QWSlqtciv2Ej2zcsYOVzSFS
RFvCxaZjMVsfDGTkJgB3jH5H7x9s8Gcj23RGFrEzSDFUuIB9IubfUVTbdTp0B5wEQ5Ay4r30rpAl
l9xbhBTMZfr2itTwk0LYlnvT06DbxIKO4X529KDn9nmayv27nJfcTFCu5Xb5T50PzARCbk/1zJpi
IwuiKokNClE+KgyuD9VByBIPS3pCo/0nxYwUUU2HpRSc4u4WvcaZdzHDdY34iy4948BE/796aUeL
wCiNXhltSJVAy5ljNlHGaYX710D0qmN1pIQB3XzJB6saQ18IRlB48nE7ib2NOL0yb+6yjlIucZHR
qBsmmOy95AWNghbz1Q8fw7mziZinARUd+svS55DR/6M0/fuej/qstXw+cb39w86fUxaW/D/es9+E
GpBesobLzeAX1jgKbDmN3PBkFZzaJareBoiXKu/cpiQzw9FLGh+SyiJR93zRrVgREDnNz9Xgk32c
HdEWoOi3HF3zYemBTgt2xfLKoiYXyj1CekvFo2e0HN/qrhlzYwTIIonvLWI7GVarm8Mkkt/TAOMt
crgg40Uf8i712DfEylB+uSsr2ZjYM4Ovhk9Sc4EqX/z3tJe9L3mRc64gn0AYSTXuTtXo+/fQk5Xg
JLNwy7TV2dPeJakOkKAerRs67cz/mv9cEQePtbZulO0/NG2jX+TgSmO4zynFOZJnPzE89NnO80pF
xyHpxR5zONVMlfuxmI8l+c4UGsV3ZyZmK+D97o7VjCtLARmnlpJA2UhLFSjG1xJxq3S7mKz9oQkp
vMKWDpHxvfiRoBxfuPVnzpysIm0dsQZKi+M7+BOu4RTHQLNCoswDqAL9VMH+rMaFeKt8qQvxHxH+
yC6RfMLMOhcfcoLwd/wDK0GhVk61PnEv3cXNipgZMj/81xzp88rGW4q/LqrtHBzqmNuEqfnuFIm3
qWg09RovrE7QaBtp67TcpTHOl0A5ElQ5nRTtWHJZaPOz+5J76/IrZgils2nouulqdtXVA3pjv5Jd
NqbhyYVkkOxcm++ZHF+Ek3/wAzhKpcFBn/slvMnVa1By+C7z0+Nc4LDB57RFi9McMJTFXWfwq2Rg
NA70b5ORZTmMs8GjvMkwsklGC4G3SKB+VW+D3DWV/9ANLOdMyud/neAlg5BkMwsWGt+l5yI4mYiT
I83tsChr9weVS/OT3DEtN+0+oru2J09ywRegNi7NH7W2znbFbgff8ggslGholjIw4lVzDh0EcKbr
QJdOOAAXcynw8f+ik+z4EPFg0gjGw0o3yvcICmhBmrG6AQsU0EaKwtcW1hHepKGKMry1fjfxTQ7u
flqHCWZqbDND0fn9zvgt5CD+okaDNYDg9z7xIXPxm8UiDYiA4YONFE7ZBMhZ53+dfQoxHL1zszNM
xs3sgHEDnh2LUqPPuP/Rtl6Xilvl4F1XFjEc+IWP2m3E/gVM8ciSDBqYwMakQ8LEJi83cQicZ4ZV
1N6PiH7eRS5+S13Y1oTjhfx1RZ9167Vgw7sepcX/SNtntNIYM9i9jsByhKcVlU3rVPYc5yTOx/Rr
k5xz+D4gIY8vt25ARstFlAtjqLsm8IDzh+vBLEIRAeHSEGlgmveD2p0OhmzVaw7V7HM2MROOaHDC
x3hA9ZR++iIKX5tbfF/eHgzLMcW09ScIXxVRNM46x+iFGleI7bTOqH/3/LvWXfpau6TDK3+Bty42
UuxOzlwrLt9z0/5XpbSSFL6ZTu5+sri/+7Jo2KJxudjfmvmkaxI+LUNpFhJ5HbIkZthVWsotJMa/
oTxGCatTFSvGFwPofCLwmOdSNcXsPPWcvYBf15PrmTqDbrweA8fTN6R76FODJdXbdAZEpZEpOMMF
gxfjD2GS+fqOW0VthX97QYAWMFswe3pAH92E1Dz+QJpZEYt77R/3aBz8g1gDxd0d1KkzsRNEC+7w
DyU5S5Lko5l/7GrlNyulsBFcrz13y2AIlM+Xq5F6HQHVY5PycZq0HPNvheuN3Gyl45X+F60o809A
qkHL8xdl957Er9Ytwl0/nBrdrgDnYZj1LLoC2qVdPWWNNQ3x4jzOxCsf1tGZIoDXtB/WNxLUiFaT
QEDK6DbF0BfgSwZFf7zf1cReUDDIimJ7c4gzXPagn+3nUTJH9SvZEK/jQ89ys9sNTTaJCMEm2IlX
GDzZaUJMSypBB3ynZL/6//28FZGXSIdFhJSoEKVFUNzV8m+rGyurvGHY7AUNaetRu6SUIoGLlcF4
7XSrpLkSa7mLitfBlgfavbCIOZdC3xqNWddfOngN2TWwXKBOIbrDPoMaPBtD5i2NrW8/kTp+GnL8
jo49rheklDAB7pov5vsFDoGI8kwYyoOebUe3lnx56uwfdNRxVkgNkrjd+8gFPZiWua7FlSxFBGZH
UwXNqvTZPuuRxqk4EEiq1eDME4FT5J2+JTWGYP1beTEFgLS/EXM7wp35cI/Fm63nzdmzWUo5pntm
KgpZvVQ08U8WulnhlrPxfDZ3V+sYrB97VDNhIwPlAouY6Rd3snfH3Dpw8evLd12bfGj9KWiUSarY
LxuMwfhXeM8EDA6tqXBmtX5ooIF1mFcyTu/t2JoggwULYE/7wfmOUn6J6grWReBq59Eg81VbRx3A
6z1ijNoIFvkQmSdJuwn/nlHm2v0r1UQcKyNxeoXlnlF5Mu1L5fb6uZyn+C8HVGFzojL7CjuSh7dQ
O5Af3tZ+0Vwke/uGYPr+1VUa7k6mY2JchwZPhLqHkh6c0Jqd74bvREswkS0xZnaaoLWvA5q3qomg
ZI30YWazLWVwOt7I64eSVW3PYvqtmv+6/GRuDjRzmfZ9pRVFVPX1pwW0M9D410toULK/WQxn2Sj9
UhctTP8d17ZydGCLl8qnjyB6R9IqLWD16de4R/li57pRpL5A8AkKDJK30M2ywWFobvgFj8z524T1
Lptd2kaxPoJpkYYXhYz61oGSF1XXBQhwlkLU1geIXbJxyquuWNKA+gocFrxCRGT3fJRyc61hfEBH
kGZ4QqQioX7fbJjRFDfHgPqiAmmu6gToWqgN/NJww1ubOeAGwbA+93xrfHsgaXjSP4WylzVmwdJr
93hQzBksdu2zK8kL/GV1+fAnz6CMcD4PKmWBymwZ7Sea7IydUjq0WBWxZ24UBfUaAou1jd5kFmOa
xNpejiNEvBhtFeOnH5rYrORmVVJW9ibHteQJR2Xxi+99yhGzdm8coSA2yUrp5/y6f3vO/WUM5LBJ
119fLiUb3sqx0hmfTyXTCHAwBh1l/3zaekFK7dVUuHoN2TxUQLcog/A7wOOHfu5MRMm9b51xsuix
bWYCXtVVqk+vUe1/im2SkUyVHZoda9X7Hd1q3HGk5V0cntQEOfWwXTUJ3APsFAbT93kt9aVAZ3NJ
tmoA05lNwKU3q2bB42oduJIUtaOMFSSM07lWMqcXZFNNX+QMQyiDUGYKRc7SadVvDUzdT/Z+BEZY
Lt8BbGRgfRUa257pn9ARjOl7MI+YJVXd56DlQJR0spQ1oiaoJIELBnebfPnKWwjnK2XKSjZ1VRgB
kOc2bQJusb6PzJNx9DTH683YLYXarkxJDXZCWHPtAxRylSpkHXmAJb58GmT6/oEJg1/R6lES56LK
METCATS50C74NMGlwP6fR4LuIDZ4zMIlKI5Ul+UlVN7gNb4pbq5SVM5a1NbNcY9iZjAKw0GZpRuA
IyD2qvqh3snpx2zuvu3yFTzJy2rCnD2/KRa69PGJbLWdZXmPrQPkXzuxQYJmaglxMJmegimCw+q2
2pCxg8EU/yqQIeqML/C+YKw/YUsbk47SgMLf3y5HyDfhTQET67mj4SZ9z2tHSH5GggDYGXYTSRRY
dKZlLORNzCYxTdK+KdMM1YAB5hg1GBf2eYTAzMkSPws0qcdWIS76kw/y9ALfntd0LzOEY4OFJ/jx
e7t+/YXfiriIkTJZcKLVa6cIR0qGapfCQaPMJ+VAOY4k531vRXBFjK6TB6oH4PHnb8VM9PzV9TYR
f5PQnJi0Mj8uZV0NlI+4/IRIX/7GipiyI6VYA1YMRpuVxSXjjkQ7MXlr2a1dUTW+Nx12kWbxKjHz
g2wuMFEMAjs0CvgMozfcFkKq+CtV6skU1YPgOdO/pdytMCsL+f2l/15cxS0tGVeP274DcKZdzRqO
FfrtaCLwYklB/HRVTlv0o1CoLDs3tLz3UYOA6QvrwYagT+H1t+eMuF70IiL6Yi5kzsSh66Gx2QQF
mg/cWM4RWJPRtOGYsxW2nXYFtQ0lx1qXdrIlh2oeO1NZapKhAHkNUqJqrvXJoK5mrJb8j6sHIg7t
knP2Gpww/JJkF4KPTXM+Tg0pDTMxZ0yuT5KJZK4tbe/35DX29L1wjNupVZ18Jp2bG3VC5o5/K5lT
pThu+4MzZxqT8ZchHUbpcZHciUcLYRTMulnOGkZgtDCZmtL90BWFRVSmZSOr4f96G9r67Mp1bGb7
ES19javK/dEv3vyNXj0yWtzE+QPzQIYhMMsecM9OIKB3QNPsoMFWhAikLg75gikql2ohmEAsGDhZ
OSZj2BJhIU8VJk/4wqDwYsKWearrGnU3hQY9gGxB+luL9xGfdW0ILujv4mLkQl3WqONy52ylvxHZ
QNS1nXcgU1x5qki7iwAaC3oqoRz2NRgRudOM6mOmO+5UzfP/FEFfrpHziXxo/8txNaYhvS3IqAQF
6kcTAEQArg86rn6OnNUZSXdyZY/HSFKO15zL+VytZeWu4xY374waQ9fn+3hXqScA/bBNeUhDRVyw
c/KmWdZF7k2GIIY0soLRaNKNj3QC6fdjaPIomqYVHPPnDWXwPH7l3KI6QuYC5Wkk/z14pHRsslTx
jUSzF5VrDELQoAutZUcLYt/dLRs0MPvpBOHT2CIC1lr7faWKno7GhmrmkwoBFXICoYvHsD6jYqzr
0iFD/+UVf4xUK/gMwk+FwdYPKuT03aCuomWBT4Znph4cMk1Mix7jKrSlPakPvhbTJ6psaajKP2YG
ZmmvI1mnWv463B5y6Jd3L8VYTzRthF3FChFLl/Aztqwd9tQnXcn+9V9kE4r/Za6z2w0wmtLR4mJe
+i22fPDYfHE8a5K3i6I74YriBuo5YVgblU+zP+fXxb44nl3TU6pWJo60sj2VbYdiJemvJsRUnWLz
70zZdwDIlh1Rsi+dcPoxQ8TEmI0XRsxxkA/MGqanxnwHQrTLiPpwsqI4bXKk5Y0y5GM7bTaLtHSL
Fsub6n7B5xe2LCy2RQXQ58QzOC2PVIVKbEb4dd0MEOlN/6K+l7dsHfVmIKSMJZ38eKFLYjGALJbU
LuGrUDypU4nLTFAzvmDU+mf7SA4UU6qBPf5YXp5iR+Jwd94amntm8/MzdNDMCBhdsZNrQzW/krLu
bxCsA1ydpCH6nVqX5en4d9ayKWnY8zZDC7cgMETmTc05Hf9MBGRgqWscAf6UQNQs3I3vCtbAMAB3
6SCfLCD4R+GeSwT1ZF/77bfuIHbev2+uPpTCBc6DdZpf+1P1wBCLZRhJKMk8oQOdMQNd7tlOpbhw
HqrX1D2GgaG/qh0AuAKOVrTGHM6MJAFl4FTO6svvxhR1h8VLPtcSwkfno3/CVQNmtHxQxtfzXgZT
zWkjmzvDvrpLXTwzBKb/vFxSXkOzcqv3L2yz+aJpIhUjo+OXYewbL84urKEFQQ42pIN6o708Xu+0
t4SCrct/bk6GRzVlJLunBfYxQexIekoRQSm4cgEt7b+f3NGD+d4e68f15C9WqGegIc9K02nXrnlD
HImVUjduVW+kwu9Bsj+ttlwrhvK1vnbjuCC5tyficHE7E+Q0isFoYSx5zjFlHlsi3rlhyhr3daLX
RwWRt6LHzh2hgL+/yK5+iHne4DWXPj2lP87dSevqBPbUqdWm2LG0vv0woVVA/B4TnWTUtJquXSax
f2lxLNZEwR+B0oqOYlL4b6AzlhBKU4VyofzeHEYk1FJ5SuInzrFQNJWvIV4KqKTWx1mKUpN4sGNZ
xXx0U3mcELHRRc4UGygSF9EVeAHa/d4gVz6u/v3TuXxiXonieqQi2UdwgQFP3/dy9rJmASJfiuxl
xNlfa6vxLfbs4Ue1lxSz5rWkAX4IHa94UuiqH2sphvLlsbqqtWNQodZMUwPPGgQFanmip/uTTg3m
eFKwxjaWQbtK5KTHkDVyiPAuOtYLhNLvP3W/a8rhdu6ZHzfBi50xfd4a84bkXD2wsn6ZUb6CTRJZ
PBD9m0RhnR+OR3Y7NontXNqufR5Ysqwv67JpX5X3yFeYXmEs3th8qHbCQdnDKGiHlRda79AAVyUC
KuMVKVDlyCaDJ1FvtGOe23Gb6x91Wkl7XJOYRDI8Pp7WMedbCG86LH0L+sjVnkoKwkjx7IKNhZnb
t9P7NEaE/eaXa5/k8LCpPc1Xoa8gJ2jqQY/5SJWGCyCOnT50tDmMv5Na20vdRAqcZXJKFLw2fWq2
bfzGyALAOjludZAnOlLsrne4FdrEIqcg2sH7Uf9YF7LlSMTrFJbQT3Dz5C2sQiFMScaDqkfRZdkg
zAi2rjv5gIrvnfpKTJ3JMVcq2BwOsgm91qWmEMp0fVn18JL6OFUReOK7/aLhdC0+6h0kBjwuqoFT
ijbeBwC5UvoH6tsMt0CWHxQ8wl4CTiVVec6XlBEJziEdSio7nxhw5yFH8Cue3DxU8vQr31meby7T
ti7Hm+Mhmgqxwq1nQmOIOF4+6uNA1RJ1q9YH2aXPwgOaYfXgrjBqdQFqJAguPE53lyTiL7AHTXB9
/lCAVEsy7DS7TVBkzYm032Th7W4cNjx9KbGvDG/ehVQVxIT4xf2rBZxPi9r/l/wg4teGUPqFOhS4
G6BPrxCFGji2ofGVYk/jyGJf+vn48iUJAbL3fwLLPfzJsiRxrl00TfM9iD8CvD86huotkB7J7kli
YEcbefCK3zACWRRpIaHRJUyFv/GY6HyJfuoJOJWsojSVCtkVnXMf/NAUBsiHdI9cH5TEdYazuEYC
VdANY5cYTD1LZX8ZMv+rbTDUx1P0c40Sk3QKEgmpAUi0Gn0v/eASEzmQ9hx390RM2DIt8N9cf/xJ
0qT0e9c4EJ5NLXxGdz1O5JXOgV5ODnENdcjtXX1P1axmiKWCZcFFAl3WnsoTIgwpN0ECWSBwHTe2
OpAiRHKG0gEMQghf5R8CHn6OQWnf++gGm3riBriRXs3NeqYHVy2nIBWcNkqDZysu/lAyzUNkI6/C
sDFnCBJbK0M5r4uvqZIu5yYp9ArF/3u1pRqG3lWgIEmdgtSd22I5Km67QgIDAx5f2xhF8Gw1ir+m
pof/m5r3QRrsIRzoJd+ZRgrNnMKi7cT2lWnLN73peh868lPV23N1jCooFDeFWovHqUpaDSDNkhRU
LJMXlDw7aYiKFlAsr4i+Dcd680vhJWXnEti0Ff1idJADbdLZ8JbCcBFhboGh44tv+Ves3zYmg6Ln
8KX+MNyOQ/UadhBaeLmFT2PZjt50jjuHOfGCLFIiT/rPQPRmoMrpN0rGXuh5utemOKG53VP3ALqv
Qb7o0iFKHVEI3PQqzCz+ctIz01DtJEh2WbZezxXjJrZX8gCN1IsCYZimlOCZPATNPsMg1vlaPOlP
mlrY7QjNo3TNx/3F1KA8x4vytxi93LxCQFkBpCGN4NOZm3SxJ7Q4dmkvs+JEjir/HSAX70HhrhY6
R6HDv0DL40JCUy70qye6wbtdQf8sUTAivLu3focGme2C+BHTMTEcewoNq4qrSZQbFv06okf6E/qz
5yLizebKCqRLUe9cVfAeqzjRgjjGzlX0dbOdc9Hz5UBkq0udB6N9P1yz9UnATjw8DSPVhIwSJAqL
dPv+cFRbOqrV+YzZBAgQTkXQkcgVFPsy5EejXiqMIOFgoR/nqxfAmdl5+RSBHNK4bgaRkNzMz9yX
P9pN/tgkClFckviZSj9PuV+Srsi6nJMaIsqpDy5kJvbBb8XKw85rh6Y929pyigVvJcSLo50CZRwA
wrvFkVyUBZKC1v1EdCBdLSUzQrcm+EMKvidlgbcZ3j/Q4M2PZBGAELTypWTPstJ9IqTRKRWM6A1W
fmxREHvbi6R+Kxi6k/W/gCvH1f/EfnbazDWxiih8jUwX56WDipzj61WzacZ4KDJs+vSz7JkJeUz9
FiHLALjBh8C8yGFQM6tHWVaHi/LMYLlPDhq8mOPxaQm6Ts27ba0NjwZJXWJdPSV7nO8PfRikNg73
P1hmscdSsqYQ8mcYFZFDoRtYoVgbd74yYrc64nuQsGFuxhXu8gGLrH8QSAYU+tsMorruONg84ZDw
LSIgP46hXBqcLhnPHTJanb5WPeTn9MT1WKqJpPjS0ZkV7lwwqOJk4i7E7inUcvCbwBHWjXm/jhWm
e9hrbmkPvG33rlRTxZY+GWHr/PBfJuNWcLalpx4GSiEobRuLSoebrrsRA6KF4nnxcmH7VqW/9EI7
zqmoCpxd92IS6MGakUcElcXGxiXJJHxePNp17SpruUepvo8dKA+DhBkKnFZKSMYLuhrg6afb/OIu
iVPVzuSLxdhq/xaMu//ItAfOsMmow1u9B7ZJy4nE+p9e2QIRxfuWu+2Q9m0wngZ9sqQCrcEV9Msl
kTNFYldKPbG3gNeEQMQCMzjT4vt6atr87VqBMpWriCeCT4My3UmX3Dr6DxBO6TwPMvcRwTyRz3YI
xu37vyHo0VQJ4aZvJTbqGJ7RsJLlkgHkSiU1KhSo0uEmu3h7pphDf5vCy+izvCbcExp3HlY+C1WN
JbT2DFym1A1Xh13P5a3sllQBSVcfxyIoxdBB0raS4bVX4woiuRFkhVXQzIAEzMjHG/d+LUlCQmYP
8c2SIFxMc21/zZMiY7wlT0PHW02dzhVhwblkKacw4kdfwIYbroltDdQsoEnAH7KKmpcYI9U5IKko
Tl+m6iocdsEbxR3IlfNx4rZxEfgvx9zVvwNo+0/Swa+8xSeAvu2ZpYQM5ySNt67IJ6SvgYB4eq6a
NC47KbldSAYX/uTxyi3CIdDHNENfSgOIArTot4PQmemNqLVrCdNYFH3csqOWkLWD1g0pPGVAnTgS
Vegp0yyEs8Vxbfxlkb1ukKcmcFIjFHCXbabvIftYef3Gu/DWVWg/dlZrEoPyrEao0QIBDko/7mut
pgEUcAHIspPaycz8gcd0Hy3E/6/UwG63Q7+R43cxvv32XkefIpU93Pg10zTTMz1qCwfdcii0wtrs
58DQtnBxpZoTI2uL3w9Ng4Pxr7dexdZm8CxxqozSCZH1CiR4M6qn3ODBB0yRwwh/S3RmGJ/ItmEN
qpOp06q8w8JenvSduNKwk10zprELo0cGNYRZ8Xpa/WcHvxPfyh8fGhpmVDGQGvLHYnhjj8guDjov
3ACbazEApj9DuH9ysK01kVhVmKiOtMirbJBRiO6wz3lZxVLJxC6FNIqIuKuPE/dL80///ztImzuG
w9C3qkBPe9IoqryusCYA9Uz547RpVxwB7kJr79R1rKC3H9R2TOeWTs3FGpdRaBuBHc3Zq629exun
WgbHRBKCrEk2ZLm27KPVMMIKYQTuvHXfu2Px5dZrJz59ybY5bvl9SuBZEP1JFn5eWPFMTtpE2CZy
jYEVaodgsNBHflIp/FQxzk+ZbPP6Xm/iHHL99aszr+UgeasrceaPjW9EK4k4EdQed2f8wGWVIByY
wwgblPNGfer7v4xSE2x+6ZYH1FyrxXEuUbr/gMagqA+RnFxz0p14iEfmOKKa3wjXcSIn4+VnN/3t
jKyO+Yv9R/eNLJIXLPFlh4X8CDXSLXneAeMmLez9ZGhqP6DKSq9jBVvhnfFKDyGoXfxjEhtRQwCS
05ZN6agaBnPoDjDmppuBZ33CtHcMAhvaDxJwAhfV9vNbT71fYmmH7fmXSJajpXbC07iMmm8cmcg+
mFgh7YuiVhtmYbRdGBtKZEr6cVOI3ndiCcxn+y5wDotSBhpuYuhZEgYefY3WxbAxuZ8aykXhfORO
Xh6J4+9L+uT5d+iKVACr5VCk+8s5kZpCYCTJRj3cQXG6ZfGPsCfbsjqClMKgKr3vcv3faXFZC+jj
oZzatYA0JL608PNZC7Bnkb+1t8gwqVHkaELEu/O3gO9o+mHdvVNnQhSC967pz3N4pNmIJ5STqw3K
yMEmcZ9bohjMe/qDRAdHe01c1XOT2pUv0kyKcifIoJgQq/bUp2taGjnbzqSqQcvmy5adU1RrcX0d
YQxV4cPjNASouxC3v7w140tx/TdnKd58eKoX5wYz38swdq3YYk7Z5dLAYcaHckhhptuVzxTbDcB8
fMUSy0kX2IdUPN3VXfNag8aaZvAtI+WF0AJaaDDHqAjzFxobdHe4sbAVDGDxeKX9AEfi2MbV7ZGI
OUjkQn0ul5ZfCG0C79zXh7ytkiuAui5tUbHvoGfQnSQW2cE3iQkSVWAHwmbuldKF3Jedy9Em6fFj
wsvcru1n3QC4+NzOzEkqgc38XYOXG7TDD74kvfERNwOX4i1Zvk6UnK8WkV+Vs17zKOvhZ4/tgwPZ
jup+iXSml3dEv6PWE5Wcynf9c8KXGm7M6JXRFNVB6IkQ7cedQ284tMwgI9BTGwTBt8Cgr0YE+DIQ
3FoBonTa0cKHpdNfT/u49DGQ2EEbzez5nTRvt4iwzCZmBGPMBlVnf3tQACnBSA4gqiUyK7XPFvkS
C0ZX1k+ZsCcgwH2kBcXQFH1p9O1SGZRcNAjvPz4Ypi5R7g2FddzpUI23hd2JlXYwQeoL7A76fuT3
RHnPg2K1K/vUUqlxRnEiRQbyGTBPvGueWBCgp5pIjyCuXaSLOlbjc2qSRMPi6dymP68CQRLNih4y
xyIIJ2mxRZb8ApKs+Wh0sBA3ZKDszUrKWcPmNmYo+IpilovrHiEiy5XrKV+S7BL2gik3faiar8LX
txY9j4hGOVa+d3GPFsezajhIOaGogrO93q0Renb9bDY128/0kqF3e8fwEnZZwf7aF1LcgxAslweM
OV2pgXUfx5CkbgVIZ5TjGkKak5y0vdnJttlb5IMe48/Ck7qTzG7TOyL+3bW+cUTDjHAlYQV9b4BP
A1i5n6sCQp4i1+4wj7VnnYzDeYG3ei9v2+55uPs4qz5IQykeUW3w3WGeYd3IgWVsPC53Q4aaxMtg
Ik7GCjynZ+ai32sMYcgp2clT9/hTgRe2scO9rNmi7u5JuTS4Hu2i8WLazqu7shKy6erH1o3zK4nI
nH3wPFibEGEY85KKaSz9Apw56F7ox4oTEEhWnM1lQd4BjuxTHIT0s0GZt84eXj5N44ZPK6p1bck5
3d5UYBrYbI2Yq4pR07gJOvcAtUtF03ThslFfLpUMPNfAgjKSG1JQ5my3LSXfgkiBFeAOq9G2lwc+
6DPYy1deZX3W1QKqHrnx6EgCn9uy6EvMYVC3Ya+dO3nzxEdt5E3VQn20BNjOU2gdPsOxiXZbwMgl
qyoSPLrzgEE1dRpz7aiMGTZrhmrosV7T3A1YUxcPWMDP3/ByVIOmOH0ITASy/Q26NOPVXhMrWcOn
NIH3xofgFTCEHl9gAPIgj+rXOIxxy14fawMhsUOxbroBMzc5eTTu/jfmX7h1p/QimmT7SecU9M2y
q6AQETXZtewxiQTms6tfkapqbRMqKkMP7gaCSPgxHmjxIRxAJwVAx/S2Xayp0Y2KimYfXMkW2Ler
4vBZzIsnhu6U1e92iYnltfL3749AJICYfJkakaT4EB8bMTVDKyp/eus29QBxbtizLqK9iKOSk4Yh
K36JwRvlpmVsSZpU+SRfrwazBIKvp/g4RWIvAj8nybfHCjE2L3ROIP/0NKZofSTni+sXUqAO7HW7
AE3oZ3oH7yp5sFb/KN0pM1epDHD8FhO8v4D0swaR0sAU6qKSr8kn0PUwAvTrFeEhyoEn3aeoyKQI
Vh6Ov6fzmBUNKHfuy7oiC5si3nsyGrDJARIb6C64B0D0+qnoaHJNq+kAHStvGzXrmUnWwTllIn/C
EMqPwHTC6wmfE8Ltu2AlLaxbJdHpiZroGVngIUgAtOwCNmDvhOemy55nHppog+cihnMMKD6BEUFB
QuJBBfFb4+aqJs4uf8AGgKRx4SMPsL1RWFOwgbYSpRjsYvFA5H41IZdQnQiJGJPJXSYnJ5GXEpnV
JbDfAcCpG3KVQJLecUBLbwswDI6Ie+W1lpGimSpetyvZyRd2FsxrM79kfJP1g2UK0kMa7jL0OUqr
ramrJC1LXJ2uq96gBRF3KSGqGKdr5lFlLeRBL4Kx8iR3k7K4Nw0VJbIxzBvUkL0kvgTWVymTRuWi
AWiKcYuKeWY2cwCfcNqiGvPNMyr/GFc7U6+Zagb1gtj4ENLsZaNMZW6n/gDjuD2CiRDoIKbAKatH
6Vv3BhS+8o6wa35H8gVggXbDAtCBtY8MYAxVy5m6rvj1Zglx56MB3tgVkZR1xTmQyVwQw2kemiv3
mf6oKNkIjYi4F3xDOi+ZIiJLKbJkAsjKuxokUz7konktVuVtc3WLzkl4pDxdNoXj/jyNcSw0rwaF
UUm1tAKxahpRjV87x4bfHYLjlhu6tt8UwH2oGFWzeAjC369yKS6fdPOt70ielsUiHbJ9kfHF6YRl
EAZ6j4Zie7Er3ff0DBAcwvaZiK53OUIVvisD4xvSj4JkkG0LmncNrBXBlZa8Cj/WD1Mzas+Zcs9l
9B7cTFJvFxv01r7BGfB6aAp6PPqTpm+z+JT+iPWEVMUDL01MRV2o2Q+7/5VWcH9wSWh6awfA/W7r
MtN6Iyu5G1QJb/sYF/q7Mg+Iklp4T0PIS5MoqzIY1OV9dOd2pykHTMN/M5biSAey/GNnsMHEqS6y
zZfeNW3MsLDiJBbaSk1UDp9f7qoqYeLBzlSi7LLPIkeaWDKV74sKMCmScqPCRd3pvB7nP98bvhy2
hd3q0PBwvfV8UD4PX0PG5EFRd1C4Ka3vjFM29ZLkf/kEiKALIF/TgU4CF2baznVb/TIOEfQw8m3G
ym0xEQAji2q+usreFag05e5ycZGsgdHNYx9Qr/tlfoD9rU0Gfvy+YSu1RDSSxMgMqkgrTQf4LBR4
ILTesyr5sKOGZmM+neO5FJpphd5Wpgj1TFUhu9QqVHfACnqkrnwgsND5IPzSkuLTFYKbudS08VnF
Rhj/edjH9cJ9bIC7U7DKQ9G5ENkfB5KBNoAWYywsEAuLkht2KBdW/kobBMTmH7JY5d93eaWcyuUq
/MRjjIXVTc5q58LoSFPWxH0F63y9buXrZEmBaIJRaeSwaWASLtbkfBM7ACwLEAdjrfLXgegjK0D8
Ip0V4lmygx/veP7Lp6Ns0WAeHpdd6ljMPZXTT9dBn7aJ7VAoafOU3PObIJBn1Y31cjjgJ8TRYspq
WMiFn1XVwwJTnbWHVVqJr7UpI+h4RaAMxxScdj5hgHRFmpoDR+igkwnbSpnEcOxZZozqhkwVOmaj
PFPvIxFIfApqvR9Nf04MijzbefAe01+vHLMTf4TdG/4lHi1cKx6ECcKeaBxG+RIOC2TZifW5xpDr
VDj8NrTcRvktpMIsaDg7n/QrxjboQ8/6METvF/ce74oXhsJe2eBp16xdVuKatIfNVBjdZAZs+/EE
EClELBYToCFo1MIbuUgYawMR5uTzXja3rapqNra7K/+CkGoL3ornjiZVR4KfzXWSSAbZe7pAnhZw
sHfrCpkLW6JsjUs8T12KtFtOGuPrYndSzotTfzofz7VhdM1yHzmm0dViQ0C672ONa1PE3LRKRkyh
ychjVOjpmDZ9pZgt3bSMElL5tcm2Q/QAw1Bo8IeqOuUSzxIus0nPujvoSY3bGJrxlHwGHi2EUwBa
ImED/XfzF1n88vRWUOsTJHlGy0JmK0ACOpD8O4lw3unb73roYvFEKu/T6hXUBGoMJtUdZfT+AhQc
Niq2AKAD+4Bf62cwB7Zpewp0BoIucz36NfhlL/e84u2XP4B2Y2ddjN3WpmpeQhkraHG8u/VS78Mx
oclIn2vndR9YlsVfs5o0RtL5ciqygbmkddLa9RcYsw8545Ve96Rov2DiE31q0T9JU/Zw5pnVi1Bq
E8Gid7nrLX1rM0Leimxq0nioy2Z2Hx/6N3TgutMwuyX01KmWQ7jbxhk4lLo3BzR22fp73uaX1kvm
DZCyVN/+nzFbz+warNdBPhiADVisjPLcklzdAyvMlA+QV+jtxB99Zbh9yP+QPVF0UtApBDgOqFZ1
vhtvtIzp6FVqS92FF3DYfQ1UqFnoJNctz53kkdznVaJ1uI0iqC9+CxnHP4qyZbeNqIhDEgQnBksQ
OjMkLF/65sXoL4WygI7zignEXwrRiIObH5qme1GjEBUUtxnnK8AbNAPLl7TzwzGAnPAsFsACkvun
eb5SqffrGgnbza7Pgon9MNWkm4/tmT8sNpmV2FzkC74g2UvYuuIs7g+6j37avgKvekgUC8+tKAoZ
iu1m3KG2w1aBYHewneZJJKVCu7u+2K9lv1INdXb6+z+RzGSlQxJK6I1DhpPpO/1SOvKgsH+mYp5X
gTbbemENguFLvISMqkbNvvwoL49dj+VkAKl4cSBio63UYwwYC35tHe/FuDgwURk1LoYGqzGzoG1v
Rhm2r1IygUKMFUfvV8+OIAsy4Sb3MZf0FkppmA8gtLo6fk3uf9leBZn/a9WMoyC0vxK7u2ZXAvDF
Kus0M1iaM1bO2WK1mysfVqyWLcSXNILXEiTuMP12o6TThdH1yonkz527MI685cAnDe4ze61hXUH9
4lMZZxCwv5SVxJbtG4xlkhLykEr9//Rat2K3o7zLjcmdw0Czk0kl6rxASwTIVytswXA6pjWrU9lw
MXCrejihChRh12jDj49/1zGrH7mTBwgfb9CEXJYKAnHSavYqZzjsAiJH0rZJtGDMl2AQ43N8DyAx
dt007PfMoxAUNzaQJALDAc48YCrHt5b4pNxLQpM8upTtQAPYFCAHMBbZ7pR93fs4h9pMHJcn7e2+
QwbNmvTZTivjvIjysOTHPWejRleJ2dq/IZfgRwwjetQ0lUZbbaHqvsMtcAxF7s+V4HWb9uDBDYRp
oBmLXEUNfvTJLiZJWn6wFDqkSx4jQE6aOBanGptawQUCrvMWlvPvFQLL/X5Mwzd4FsHZJQUaxLXd
6+MFMUH5BOKLu6FVhdkWQU0UkstcGX4gpPh9A+woWff7l7xsTsI5U1pCkZQiRmnzeGTjtaUhL6wr
y+JzHwyWSoVE16b/eNi31PvKDBFWVnqRMaiB3ylkCPNzPJVJxsBuSGB0DDm5eyR66mnz0FP+7Ncm
bqdBqdEqNGV8J1WygcnxvWwTEqA92nm+Hv2qmC3YZRO92f6t+TpOpN0HKDoou4wKyRU8o1tJtqaz
WzQ3dXMeSrgGhCIkAnCrOxTpeCc1m2E5QX8Th7rQJcltBxBUuohD0wuh4YSQpoNFXFDzNbINroQs
xfWIwoLQtGMQlVMzqlAOpCE3ZMZkkQEnKb10z59UAqkSV1MPnB9wdjyo0S5v+I+8r/ZaqNBR9Rjt
3j2YUjbX1VDmQutAHgx48ySSCyjMrkDz1NY/B9ipjJFZfIDSAofnuMQ+M4exQTJ/IdI0sOEXoFbM
lGkcybcGaCcNE7EEf7Y5CEnlIJ8dG1IeK7LJM8iBM/Ty1R58XsSrEEkf/e297yCa6dAHaf//k36G
B4iUpwgEGcgtlXWF4MrzSbNjEv+3J/YRJrHal+KJF6LS4vbn26ajnElZ4lWtZ58xtaNaFS4Cp9r9
P8PG88mxLMRakhiCokB9VQ8amoTKZYNGABfLG46YmOcXeiEPhJPI3LLyzfOMUMxt39Y3GBt+VDhq
PorIshhXU3p5VHmDhZJcYdWwamvscKP4O1aGTo2wgVV0+vMqHP2BwegHLD2UmBqzy5TUpTMxOy4c
OOJUnNcZNqhthEAIuiMUOWYp6BoAJd671d9Ym0Q0MTwT0qoBbsUvfMqmcn7ln3tPXNwp5vBWBJAg
GOHgOEYS2IQ5AFK78XwA3L2fp2IKZhEFcWrrvLvJ5EBkIc6JyQI7hXH736UyWGXnns/Yx+exIT5d
bdC0GJden//0Q/iCMXsBnfnvWAQ9vziekMXBddbEU5PK6CsVWC2amwLe1SGR2+sUrReVa2yyd0Hq
NecaxM0xoZfrpSUQzg2qtddGzvHOvsLLwDro31g4/xrgjrTkBx8XS1NDH62dYA4wiu18EFo5gtoG
AOQxqhlsTJpuwIppp3JB4AQ/9fISMUg1Y0LLZBoVYs7AnSFIJiedV4oQUK8fdkWaQqHOGLSNlTNi
QFHDVceki1H3fqYtxRzpalNRrhIJ49ROJjNXVnEeqtCle+qwlCcHeS6zoWYwyL2brQ7iA7L6w+AN
eBbPTOB7w3Xbi4zElF1oGmSZira/pl2z+sSJNf7gsxF5LXESJONAKtdqIlxc8QwHY1oSogsnTfUu
iq93V3ZK7uCBWAFaiB/GK+jiONVj11tbcSWMOIJb1tnVrc0Q+RDpsBagoi33/oLZi90QNJAq+nsw
17pdm9OQy9NmAsFxap/R3+jfan8nJsYS6RSaFsKUhQH7hDDSOQVf5qEvR27nDBSVjYB1GQRmoQDC
n901zj+t/aNXJu07jDMllmkbqDeyaIwoCI49b9RCsgBska5gPRdZHj6bkVwEesx5lbM4Zo3HrX8k
Dlvl0xo872KSnGCHDzzLuEeCeM2VntD1MHSmZ45cPh2u1SumJyAd1EDpZ09cC19QlKTX/GTN0twl
t2nk/iwvKNmTq3WmmrSKgOTyDJIa7/v1+4E+sCJrpb8NZLlyUG6UwYSUuLO4cVhfOTIUHbaPbLd6
nhxA01vaRV5QskabtqVALWByNaRJm1WmaoY8XiKop6wdguW4Um7s6qPKeMkB14u04LpXchrU+Ezw
jO/QcukRALTc+4Di1PyNZwZ7EGtRhkHVL7eQmcOiQIxO6wXR+YaCWPHuBK3mu7bns1lgqS+x5EXS
+OHZGe9so6QHyLonryHmIfnq7TSukEU42hTDaZ0MU8IdWa0qxwIkl3mwLS8lpit9LfiOhYH30yIK
sbZbtvPQpgk0htd7jaww1Pw8HX42Ub/yg8GKN7eWYNZhLPb2zxoFwKF1KI/QaKXaaoLnidb1O/+y
bz91bN7LYSLnJr8j4xDahdKxdkNLTwZuTPd+G7g2YmDSCxHgrR2UgltCNoLRW+dcwCTlafoN/+qU
v/h1CXI78Vw5TDTIjeoH6TKNY3dqe7Rwr5cjG75+l3QG8BuW9VceKs2nMvifPWnWAayatMuWnrVq
ZLJh8LZI+koNgDSQ8t44lb31wNDMzh9GpZKk0s04CZlpZXeoTDwDHMuIDsk4Wcj3o1oVMSH1ihaB
WWIyi40WBuWb+B6oi14LpsNo5OyNw1vXnhkuvk0N0xobtsAW0bYCw1z8dEDDnfhvxUq1pOZ7ZMVo
CLJS3jNPLt600kuXvGT8tVnIG5LHjUkRtlQEw6MYoeGMeYPT3VT4YTahNpleXjiX1gZ8hgIZVe0u
9fpsww5CZna5eKfuraaQEMqKzDzSa/qFeBSRWi15j1mj9j+IvjQiNskEDCsi38TYCtgAtRU8Wdwl
SYreD3bjVd6OdJznD3rlD7OO7OGTTI4zzA8UOeZk97cwlD7/tWwZu/sLVj0Foo9TB0n9RTzSr0FK
MFvjeNhNdGHJSkQqOm7gtBswyY2Ts1l0yn6poh9MVm5axxfeg4W5TT8nSJJHDHUGd725/Hhud03r
h7TuCdgBj85VkvobPAtBedvZpZBO8Bkhhb3c2YFY9ZcfJZccjgGgC/bVrppeWJQkiGsJsOFZH62b
z6h/t1SleETWDWOGq04NjgWfo2grlFUSN80xKrnbRm2Tk954ugt6nAM8/fOVZQommvRN3YnhwHjj
wH2vy5IT6+bCbiqZ7fdC8DA3uC5Cmfi21soEjQcOxPU4kZexMnPGg1hqIFAp5v1bbnX5r0ZR7l/o
i6Du51gwqBZOi524gpce6haODDIkghHRnw9M1Z5otWJnnT9ahKsJanX3bCnxuOxLxfeRdrIeTV+w
OKP16HhpSOGqi7mnOUnNzNDXFQ33nqJs4GkIMzl7b/JKl97wFLHkAEd6+tMVvLOz9oKw5jYO3R0f
AvxA7mBo8fC1+fOyYNFMIQgXXCW1IBI+q+G6cpzFwwNzqopuhdBz1zGYZNq2eHvp++zs+7cb7j+X
CZEK8+ZY2Kyothp91/2GsRO4b6MjD8Tyl23ODC7ZImwZo8/nAsv7jGstkqE8K/rXG6ju/6bgKRdq
IrGD8Ywi6a0hl5/60yaoiJ+PS4au543VjomSqpSY2kwW+7QDq9qyzaMr+kbAOKNAF+IHDufKCXAP
RXCUsGHK714HbgeNKoptmEQCY+QYQ8/tWAqZQrppViW0mK39MuSfOTMs8pni04p/QZED2zdic46d
ERRwQFHOtGRX7BQC1phP0ijoBweGYB+taG9CGI2nIyoysMf8wVmdBHrxTyQIWIfGZmNIOkGaU208
sY2C/fSRxerMyoUWhmkcT+Z55mARcbLghMENcxWvEk9Z+NKB27hfXUZ4BnpaxPni4ShIPVfenG9i
3NK43anH58XDK/uJ0JX++HAsOA+QxYz0boxAvAKCGqT2Z5G1WBMSnIKX4GeAZ7XWF5S7Kcw8I6+s
nT0oeBrAcv6/ioxf0AY3bemK9mp8FBLt93wJPpHxC4GMZgPbcXNUc9avD7pMdzVqYtwPJsIoiMSY
jhJoSjuHzhygTLyIO5jVSFS6xyIAabGlqut4qbU3J3ZYKz5NUJyIhUvbfzcpWLzvGWAyHiqkgF6D
wX44IIBQ1ydDrP7v0ht63n/NI7Vc0Lp1c+NMkmApfUVsdYiu5Armid3ClQ+1KPYdv7eV1eroE6LC
Qt6rit8uEXvSK6YlqOU7z+p9Le3JB1LI5Yy0Dp6jP+4yio2Yql1gpbfMnThNqmrmydIpeZAyeRzs
sJEtlXB5FU40DdbWP0uzgnwPTLIZEJcJRMVGRHdV87Btwb59mJY7Fj0l2EYN70RkgD2WoX7+WbDJ
VEcu9fR267s0dNN462GPtpV75HnTcjlRKCAv5ganCr0OEEveHHC5Ntkqc/gWthrKbI+zfOVl2N8e
ixNhzROiGDl/rG+PW7yfz91lt/Wk8W1v/yG/hU2NIG7zTWsZj6GYDopSJtQkuqtBpwq2NY4q9aqI
N4iuxGSayxJm5tavhZv+NbYtumNXX1mxSHPJKM+A2YMZ3ZgpiUHGtOh8vpnwcrVuw1qp4fKQo6cI
gd9UhcyYIyeSx/MIZR4OTRLLhUa8ciU0zjUMVnWls/K7FRIRt0qupfF0IMT0VmFdqC2RLXWrlPq2
SRncZ7NB+uctJZcZestH84a0uKJ2Ql6g8rDkQf9dJBfKHruwh2OtZoBoj4Tw+ltQbmxIF9IA0s85
gYPghgLrNuCKRA857xJMdY/Mqut2hj56b8LX232pNmxVjdFxj7Ua16WvKrgjL1vdkeIGrBaELVky
vLj6uXFQsbm3wksuo0Li3uoUsrl0M0cjykr2D7ZwzoVJeXFm0G+7pTS1zgQMn1Ua7wUu+dwg7BpA
/cc2ehG+WsrmzEtZ5XkCgeSIk1Ydb0HCZ3EsN7JN12mBLdhofLLpU5nuYfsKQqTyb2SjsR2kQleJ
QvYfivpAfLCF318w+XAdBKZUhBGbNi2OblDaqmY+G4OifKECz52sPzAy+9elXyYApWnv0N1TWXof
PYoYDYJWdz4VtUfZoKN5UnjRWkJoDdjchMJYdV/0sEEekcbr7vmtfpOy4dDfYW7upWV3622Aabpa
RuYSWNcn0J/L3dME8Rrd3b6IFh0rEAIqTVPiMmw90zhddVTioYFHCt7Y84dvijNVhTc79se55A2e
s2oe07tzUaXNZ6WqnFYqGhrTvFm4SEy+KopVsmJcV9F+1DHl1YQcTov/kCx4Azx1WyAzci0XGaHf
5R0Q3Am0+TEmQFaxAbIOkFxqG22/gDSF4AnmWoqN51rQ5mmsl1XUhbfjTiXKblw0hw7KuYpBArko
jAmJgVw67lC5mZXoCwbJ5+QR2XjKFvKy0Owm7t04XiJIdaJbbYrJMUeHLXG2UabNC3hvhuY6FFQU
P9dVHlpdYmyEa5bO+WXbgxUCsJI7w6Bczft6tG4Ub+XEyeAbykt6WhO2k4bObL6vYc7+4t771FF2
+8YWPzsWWb/zy5n79iD058l0Cw6AU0RJDk2FyiGGCLP1MK4ojw5QufFHavY8uwben5GeGxYpnVes
OxN0RV+NezPGAgIaz/+tiJy6NSWOVx/Sxp8HtTuY0hZe2Q5PRfZ1qQa59F8jBk04niMrPl4eZBWf
uswxQae/fg2FKZd1kSMuFl8ua2njM4zYS6WHoxQgw6XvpOh65JFBP/ccoxuotagqITazaZ7ZzKBE
VOHimcFoUA52Vy25UAFIUPaejGCr3PeSSom3ri3jJQYdYFkTW7en5KoaSqf7/hSg6OjnMHob3KVh
X8/DZxUwji1HkPPdNRhp8dbWPAnN53N+qPSr/88iKjT20nQA+7PbhBMBzWKx98TdUu0LuMwnjGUj
NCZTHPTXvIbFvxdT6Pu+/EVcn1f/cBnRNYqk59c9GuqZXPq+C6NjoxDalzJY4al4KHbjLlMlrdtQ
aDpb4tOzN7O45RMd2+RtcFEFyafo/xoOr7K6zXAAZn2QUjUmXxSl4guCrsUR9kmCB+g4n3PG7JyD
X5VhBiohZtN9wLHvrzVl41jKoHC0vyEiosKqfI3p+kJWhH9URFj9J2ajQKicHr1+ViAWrZuM2SJq
C42uqJSL+N8R9oVkpEuliHzN3ytapVGoi2a2q5epgQ6yxwSIhvxXsNGYgSyZJPPLD0CmPadp1H+A
9l6VMkVAXUVlLnuLZQjp+ce4bMFK9YSY7puGzmqqqTn+Q/8FEKX93hKwi21dg6QWPhPFS/Ifmn94
kHPHaWs0XKBJlVNalryFJH9x85g7Gj8UQfQBcVDjv5P0oWvPtIo9WU4nFsBZ1czhBENMo0BT+ySA
qGbOZr7wEr/BAUEBeNEfwvzfSrWuJjGvOCukXrVZJBn5doAQ+Yck3Bd7B2qq4QefOXqsApeOMUAV
S2g732lMxlcdTNTlOxWtT21gdivCuruw/jknYWyveSP3Go/m7Sif93mgSe/mzCKHZjFqcpu5gp0p
Hw7R7SIv7X4CRMRdecY6dZy4Fp2WIu9wVvyIsBCCnbGYh5Uk9R3g2CONc6MK4/aEf/R6tu1CeZu5
1C2d3K3F7nKlhXFd4mTbYqMGEPIyEe772WSHooiaJYHwLAF/hOW+VE0nIg3nd3j5anhSrEtruZxI
ShW4PHqWw3CSsDAaHgjlCjzimWzGuvPacHk2Me4XvBmOGByMuHRozwQ8bg+jthBW4vDFoM8z1oZc
GhLYiwfnd/X04OBhnwUlZTXxhoBmNm7e8rj9hVljmzMUTah9nfVrvwT0PFO2K/yZcpYptze9I64v
DhBIRNHxd73SrARAkTTWxd6pQstBn0JuMbEIC0Rur05xRQuWC/Obv5V0NVAcZbE71TyiVtp3R4qA
nWoMJRgyc4Sxtv4cprY3xkT1juZaNT10i1OvX5c3eifOMz1DZJa2A+3nZtYQaxxi7tRSpnQjlmdv
L7STss/kAez45qS9ec4lH0Cb1cYyXoFmnbqS5IdWMloghuUWrmIBveVqB6JB8yL5jVliOvFdDAcP
D9IJJd8EsagUWUBqrqcFgjS5JEB4c8C5GR51+d3z4iRG6T6Pp7OVaxHSkpPqa+NR3tJHHOok5fFj
Ck6CCzvNjbxT5vfGEHIi2pS7b42imqJsaWkdHa5XA1a24mk/uHglSt4j8x3DQxLoQ6iucKrubDlY
JB/E5JzFYA2FPP0hQAINsZTcd9fG80TBJzgMrrj4ZGeBgSufP5cNawrCRj136p5vplzmpEFyOXlH
yjx87nsNAiaavdrd/5GqLVuGV3RJUota/P844W90DBUIOKPPa782gtb2s282zJzPNfOYq5DUi1Gi
9wJ2bty3mgFQh0dpRjMoBjGUE7WA/Nxl7RRmPklMLFIfyyQeLTHpiKGTXPAsriHCGnrUFZ6M/tn9
JDg0JyzwnkQ9o/eT40I9/TB8s2XOjmRXA+//ryqZTEuu/UUfMtWAgyRdrRVynfKGR0aKhEtfzQQp
O3KM/kP4EgoeixWYIzIhWnCBAG30ywepAW6bjCAMWCof0YhUWmdLty+zOJMZ7/ypSmOBi6XfX37e
HK1O9J4IS3EK6C6FCkFsGvwG4LYU2VugC8JyP0NZQdnvtURwnq1F4qphB9drOXUfCeV2/+lzoYdD
+EOCZZqLGcdqAm9R2dPAuhIfKJ/AOEzwHUZd2yhRQnmXNDG2j9izP2Ws+KkwCIBSC4rcqbo4sPQs
KQOOqPdIzuHTfSSFy9uHrEBDROFk7iBxNNM/2THmKpnITS40IXrFaSwAD70C6Ymuaysoj+Jq3nJZ
A1affK1wFWPBZ3aL38YrV5TJ3pdKckmW5Lt6JOBdKeBNeKahgcqWAD7DB7LnNNxu0oAA6KY5tgrj
NVZHMnGwXxLKpg3Q/ZGzJUGvlaWPq/HU6574lM/V2jAVOUsH9qK1SUV79Kzkal6QB5wtZjpbFfsc
OSMIJvyp5b0sXzzGdsfg1AhHH+2/ACMCjjJ38NbffEBBbO7teAVW/9SndX2DMsi6YRfL/8KNMHyM
DCHxJf19aywuBzksoYjKmMc3ZNRqlOSELUi4vDF6g2K6er6m3NpFKGLf1gIeyt/Fh+0VGRapeB31
NGDutPjiVmRrEVCjQ6FFIEVoxokW41e8VM7RSIZRQ3Yla+VR4pyz4DbTxmJR+6jZqtpX2qgJvoym
03jptcYKoioygpiU3DjDICBkgErpLdaHLEuUNVc34A+g4OPAAewSoQEfye88qexWB3Jh0lJOjFTB
Ph0JWh3kwzM+pjGoxK0kffqCuqfEuAY+bxqWfjLxLa1TZLwW3epDGsEwNgK6y7s7FjwSDN4pmFoR
NhjmMvh76htwFh1N
`protect end_protected
