`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
B7AS54ZpMEBvU7DY7LXlmwZnTc31mQhijXcXYu4R9LocI+VzC4owVmtAUtHJFC9jl5qgOwW+YEdu
7zfLeJ6JnlOIrDg1KVJ5jZnkDdzT69wZTkCCDhPYhbZL3V2NDpURVxOPgGvIpkFvNqOCFRrnlqcW
Kirkf2YaIG+NRFUR3JudNrn45zn069L9gAD/xGyD7wdUcgMn1CjAuxjCf9YmiC3GbNhmnrMaBmPH
xvx8bqm7P3dpfMRruvsGkjyG1ZzvnqMPnZzjJiS/nYwtgcPF1ZSoadZUvTSGkArDPZHzN0HszkMx
ztUNVM71lUuG6I0Os53AL8RJd4my2ufbmznBaQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="22WNz460ZFdN6tzC3wHB0W01jKxS7yXDKwQ6NteEZ94="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12192)
`protect data_block
QgbUyCSeE3REkxAX2AamkqHkYkIBXgR2/8pvAgZaMOBjcpsiSKrBN6KxwRzWOXFbre7YhjiKWIbK
0YAw1ifaUtBLStL0qJMkAa+Ui6Fi0+uWNYNC8WeJgTR54rydIhMeGqoKj4iOlWjkYY2N6Okrx5vq
yXCh/FAEpHrdn7GNfMR328NPAxQoKgzdoXtiWCWSPKIjNTQx5+vGgtYNnK9YZ3aO2CiP8T8zm/1Q
0iGKdGUzekgl9XBjVWc0ggcArFlTpCglQ2Ja0Ho+JmkIClR3Zr6om6FSr/vFB3T0amKeVvVRzNRt
0KP6Ff3/EDSdo87tldkLHyBq3Fejym1m3y49gQJK6lk+wTEBnl6bm1sHX9tB2EsoiKzhulFTKbxu
KeAhDJQO5aOD6YV5w30YI94EDPN5WAUwfLP4LX0azoDa0LwIs2CRAWLqBIQCSQ8UOkW/88qNFIp5
ZQFM7N5T3RJJlFlEUuFAeaS5+gO6cEIrdZVhMqfhLqyS5IVJV9yp6/cFgB+cPDxMUasW/DVgRjdL
EUMziF5e0zcpfbAmLaxKaO2TJNK0e8CJueEVO8WRsDXBPpkiFXfPWN3SY0P2qb3ZzMP47FCeyKsg
SZxp4qyBIrCal8UQNIopLtY4Bu7rbO5adM+T9fRP0BY/csnWQqb44RA5O2CBFFbquo+rwcNF9637
9s4/XtUckbyc5M5Y+P5xIIWd10aHQTUEvdGCyIocU0ulLQbDNf37XL0uLcfwYmsXFY6vNPKTvl1/
EKPxo8RzCuETqAaI6m2VAWWshL1MhaZIM9aDaeDdf2HMMweJiGaHSveh6iGOfqV1Hzs/z+fM6498
DMGkDOEt7DCFBL++IhCHv+Z+Zw7vEckD2NSoz2XIo/m9n4i9DuyWHuOesSgWIny0d1tnhWjcTDgM
cdEkdu34SlLppFDn+VczWi0tN0nL06CMOYl9h95+yxoU4yozPPlTRPxWpXUB5S7N0NfsgUJRXw6A
b1r5XWtLXLaI72Yn5s/Obl6oNu+3P2f31IKjJDO6YZaK52GEjcobJdUE/g7jdhpnw6T/38yd9rcZ
q+xBOGsrvDOOPlpUsyvbYA9vY5k2CV6XZzqToReYwOdk8hM5GikYZU/htpFqSu1ujpHzT6/buOSC
xhMSaJtl4erF+GLgMzvmtRwzFZXp3/ecnd68uEwkv7qls17rYRyBU/g1EFtpQU+qE0eTFgrFEqC0
HaI8n8TtRgzVoq6MR1mV1mI3X9QpFETMcIp1ga0wVYEDp3lIhKXqCo/EKtJKxIgrG7uXvyAJioVA
j01JiBxIMgJaBrIlc9PSywUkM35a+SpkWzBRjCXo5XHSwQo2lpHtE6DP/zHvXzQuZgjz7RknaJ6g
+rVuEyt0pA1XAw6o3GcMshIqTWN57pCympTesRF8pFHcDhMVlZ30HGO2dL45Iu2Znekn4blrRIa6
jDgcssX82eIS4QLWs/JLa2DaB6NaNXZ5sTWarXxRfACbwAhBCpLTnmt0mqbwLLeM6hk8d3m4jqoi
GVFIaWUQNJU3aGUBtM6xQhR6rFjXQjTF9UZRd5u3iwS2XvHAyEUTqCtEAA4kbs3gO3brDCK9D4zq
zd0OYNLfy/163qi84+8ZYnLPDTzavgNYzndEQT9FgEwuFGsvI+LvJYzQER6Yor8YdTEYi7yEKWES
YGr1hv8WU9hPq/e64otdN3nNSQBAYunXxo/w8udNdqWN8SzTwGwzFCZVKZI7d/u/05JfcSm46UHI
cVYWmNdEN4D/sa6mvjH0wIpKKDvA283W1F5RfMQ99uhWmB2WpI9HVwcBrAhN8l7evZXI3Kvc59f6
ZP/r7R+ZQMq+zH+cQdz/H1orCMuItyqQU1eyYdVq8gvdKRwRsteFr9BspUnq4bGRvoAXwHzl6FA8
Uf8OXdOK2TjdfD12U9HjTOEWTHK7YT0MFCG7ZxOQCoe2sGrjgpXmXQpFRcXN3Tqw/gLfPbIJb30H
1yNEQsb310Hf4/5o7dFnoCxtjNoOXc3TLC+Zv7t+R+F1dbfGMGjRzFhVZbH8oqakIa3TU+n4BP/c
s/DuStYiQgkRY2xn8QqHTtGyx5ynZsYDVO4MDVJnQSo/bCQ2CGHiWHgihBFe6xEJek4dZpJekZES
GN+MXCsFh3+wTEdDK8JLrSpU4pBmB4t1//pnFfhsaO7txtVmkCD9itRlz4AvoF+Mx/mTZeDcqjzJ
LL2WBLpvcR1+QynQh273mto9LXxhftZ2U93SQAfc6glzQTM4ZbaqMgs3ks341Q2U9Jq6ZNr0W6JU
QenuICtFmIAiSEKm+PZRLA6LAC75XkytW3cG4zlLpAJRUF/sUnalyED1e3Q6ZH8H0hVUs8kxI9B3
gWcRmXplU2LFkRr+wIMiTK6CCKv9FArOBoyqso6LZR2W7J6SC76tMknNAPkg1bSSpbRZIxn41ZWV
quvUo5q1Rb32Swp1yGT2PncpmJX4oVb4F4OPO35PocW1lYKQbuXDt5U8UqtLKvqqe1xp1nQZkSaF
4VoAoyRzTuK6/CsqJIy6QT8eqw6d6/fcS9E1LlyptgJqto/DEQodLhGxR8NDsMhboHGuqPb/JUcn
R3Q0BHcMr3zgOGeRb8KLyEckm3A+kjN5K8mo5MQ1JZ1mMbHN3X20wS67I2yv8YoT3Aao/Pkd6MQl
i1TUsnhbsXxcF/lUFX2OpAMGPbd9aLNTzeXDup9AkbwYInqyLiCKS/CJRPfWDeq7+qbmakkJWxbC
ro+963uoTwNxnI53iOvh6kN5xxm0TTX/kjiPMo53B290SmddZxlIVjm7hX+zFaXagoJfW1O+95IW
xDI5WOEG2vmAHinDPYIn1qVd4qIXw4F1HpH19P8wBPRr8NDRDq+DPnFq9Wcj6yp2ynFKT1MKxZOY
4lqOAkSt6gdt4AyydTeRRx1neKQ8/eRUE/jO6yms5pd0NhhNib0EgXkzyXDSxpZ1WJeVwOXfFepe
HgkZS7/q7+cNpdD4If8Bb5NxssNF6Q/AXD7y2a1X0xBTCQuWT8QjI2U+ge8Pz4dhCx+OaqezHe+4
qjYK313r2zITzMtUe8kUCJsk0TQno9v/B6pHEVg57DSkHbKALDAyi81xPAa4jsAB8meGoGszVe/+
zUuquN14uDVF6btqRpsfnGdSdIp/aDZSa9/5QRKFLIQxrh1aLb2bYJ1+k2/qtHANsKTcfVUMWCD4
dQ/NrJ6VIPu7XEwT9dvOSUUBbrihKG6Zt6zl1MgRKwi4ZW6sSHNBqvf+5eqPwXrtovBaooZTo8TI
pVuScAY71ceDUC9v4Dh0cLbNwUaw8ixjriZV0QATBtQwYbSDCHNlRsiw4oI4S8Y+Bw3QDuIDkFw8
KyrYzQC25DxKQf1O+MXAD6hwDGlLvhkYmETo++3r41SnGSWmTxITQDlBDibNeciUAgW+fpny+6Od
dEacd+aKracvLvH6citswP4i05SKCCkWOWry4mmlz0zhKUqnG3xsfmpprGwPZIN6WjgO+YE95D8K
AAhTKnTHP0B/RFU8lSXqD27K7iHggXB9PwaAa6DU6Pt3JmRRoZQ0ag2lSELZvPHTi41bAD9nZq1x
9b6U0rvCWxXyeQCKxqpEhniortV3lr0X7bA/xLitJK6D5nrjhY/TYnOI2lVprpwJuQweIUAGRaG8
YJLXglMw5NwDKPt+u+BUqMTODLG5+RAhrtfMqZqmR5WS/NZIWKyiaBrtmO+FMaqWIMZG+25i3Pr/
oTyT4Lllu33wYbPqDszGHo8NjePJiN6tzOhRHVk+mmT6rfsPUPXddU0w0pFkZ3k/3QAFS0Hb4ITK
6REO6MkmS/npg3+ugWxGZNfHAqC3R1wCgW8wpfZ8MVXcTmHNH8NCqtbKHgd5WDwmhxhv/XlaFrA7
Lr3NRcADH8dKQNWl3zE6VNX/wF1nKW9Znkr6gjVWo5+T0KlOQfGA4c/pqB9t3MzPeqXKkO2mV8Kc
M/QcY1C9aaxSLu8ZWP4n9vmVgUjwjuBRYXDdWhAd6hxe1x/lHNmNZ835KGVy+G0WyiH9b4Aqof2X
joCo39r65O2m98kisHbBIh/XUVfHnmK/DdzaU5n7VwhXKHKKHjsXkF2Y7UwIF8WVSjtrlEG6n0le
Iw0N/6o92rky+sPSqmzdYyHOxdjkm8Ryj/Z3oV96TylGXNTOh0vgX36kJOkhWJUSBxYmg9tBXZNB
4hGlSjCb87aqk4JSbsqhsGWfRL2c4y4U6UweDS9EbGHOHQozl35LdyWi13Rv7Vfa8JL7T8LLGJDI
mN2j1J+JR51FM+HxhhYFTSLPOGRAypqyJHTJ82DBLq3xae2BXqeNFR/hlmet0t3XoSgiN5vpQ7wd
THn33mUpp7BRvnZtn6e1TTVSovYknzoCYPByaeNNTriPge038CMCaQ1FurE80fOGHbMu4IZSmYmY
U9TiXYiHfXqn+IQa9FW4fCsLds6R5KJUsk03qZVBBGm+8X6OXCFrqPD/5mfXjul61+0mzPog/Qcw
Y9BCKFPxkAMzNQFlMLknCXyTg+ewGn77ag7eQCEaCBfC6hULWboqqGxxnPUj3me9nHBEMDfZ6bzk
mpPFWuJ07ZQM5yvIpvPjBguAokPG/tdfBwbuq7gdr35wH8pQ8vROXzazcQatYL2OjuYrPkPlivko
MWVpZzMJ1j8wVGuC8qcUK5mEsVmebtkyxWMmuT07IgeMWuLBVKpfOSOHzEjJkQnBUMGAbKLYIrsG
inOD51kXmJvLKBjYGomg62OalOBC1SihrTehJhmWfebyR6pyhFFN22zSkGdJEfn8H8rqhrWl1k9d
dzx4dWnSRlquUfYDywBhryvZ02mBGYrPE6l1QFw15k+lQ+b4Cr40qn2UWJUTdfzOAT3d6CiHEzMy
ZQbgu77oY0c25a3hYIl3YDiP4qhSe4ZDZmDarZfp/3p4CyoRYeexTsEE5awF6CfTSQx7ZUTjWtFj
0HN7ocRr9bnLZHoPro2SMCc5oFPgltia94nmmuDMYfEUG7fY/kyjBQOzdVRFj2ckOJ67msNa0DJJ
2ME0inllTrZbD/G8MhhgrCJGvPgZ3p8ezkBrzSkMiPJCy5uUyTgxJTdGcbuvMDOWeJeiy+eSoodw
oII4kyeHH0PkhM6yHpkJgfl/DkEm/seegv9dkAsFJmThVCHbZJb0GkosxjiYJ0DKx6jsEC1MfQAx
W+edG688/54XLi09z4DGf3oO7TQA299BBC/3oZMARtAo1D95xILIz/BeHWQeqHDIqBwQjIaMvqs0
yUR1nsxfeB6wD47fpH947NpnlIOHzHcP5hlcoB/zhxDhq/CefY0AcI9/XIGcodw6aYEcWiyKVXod
NciahAHKLWJL47DZVKJPLDDvpCasCLxFSuVv/cxtqCrK/Q4AKvMr+tnJzWZL/Kc7z6H0wEK5TV6j
6ksNKjGn8SdWqnClP9k+GaiAq3n/fy/W1t1Q1DLr7QYI47OX0l5vycJ+Pr+NADUjDJNsNm9F8Nfl
HfeY9cGyyoBIY7I6RU5lakY/Z0M8zocUE19Ch/PYT2922MZLgPuFjWxDi3xum26c7YuB0L6le0RE
caNlYBZl4/OUj4ZOUX69kImk2fE/1SDEQQEGxgCp5Z/o4Dw/rrbqQEwL+NtShs2w4mlf7T8wougj
N0T9+qOgK3QCmoGIYhTvcYt8OBGT2idi/eZUS1+j/Ieg+Li/g1B6w+n+Evr6SLDjlDnvDr7uf2vn
UsLFpXC60MDS+cgkz5YcsCVQEVJ+m+VCzR+B7oTEt6tqjdqhkyiziMUhMpSYI4GW1CXXXQhkzIT8
kml1UzujYS4qjLFlY16T+N3ZEHTvE6Eg8iMIhdX26O/H1xWQqdvxkQEXX0uOIsUuXItJxuqTc+t3
N3dyQ5K6yacDgPRbGbp9R0zDmb+Zoy3KMbT4qNBDCVEBEdW6Q0fPsbrD4on8gkO67NYdWQuoyBCo
YDYoFmCOQGirKis1WsAeEUXMvmemarsVZFTlm+4Jlom/kx2gmHyumJAtw594x1kLzGe8smq3KyOI
sE/UdnLdjC88KqvnrylcAlSP2pxbbGL9TXyOYHCogjoTFuocYjWFRZU5Wbr07zI0QyEGBe2pRGtZ
WfGwrby1GnsqSuSpZiFi69iwhy5h4b66XWC8miPgvjpS4eGD2nhEuwTMHPYcIGNzib0dMzusO4Cg
A5hapUxUpW7BYcvP52Bf+GxIzOfx07H9Lw81NVTSAa4/bAoI5jIaLVXcWn5lDoRKxDg8RbWlTf7D
walDIOQyzF3R6mR6meha+jcwGNlQB5A/6lgtxe4SQzzaZUpNVQ14ix7U3jlGVcXSqbrH22VP9mQn
Jbu6wOnCRfe09wAN8ee44DWRV+gKsQl7Yp6fjNycpvJ4ZmfdkV1tT6rsapRNLO2D+mu7X14gUtXN
JYZHotwyyZx71NyXeMSVMtovjcHcQThoRUT0ZO5Wehg9ogzVahx3pgUdIol4zGjd5zrNeqJfIb9Y
CfGDWVu2F7tL4GJ+cQyEBLojUaOTTkgS/1Oh90dUJR80wG/AHyVII9GAS9pDoXp1CutC5J9TnOlB
FVqMti5RkcfHTq32K92bAdh7eXJm124H/pOWNx0CTuD2528pU7TZPnf8YpswwuDt2WfRFKAlwLj+
ohO+vGRLRZfLWcYUTIOzI4liXMv6jUNF3PTLqhflqd7LhX7PvMvP8fuaWqp+dypOhQHwnP+zTVnM
7V6g4FR0lKlxiknDuWtxWEIAAhX5kauuuv2t9aNJ754nhQxpmLhyVq41uus8w4hiJXy17UNjtkLV
ksA6/pYOLZky+/I08LJGTmxwHa7m2dl/icU+b5N1HKX2Xk3DaZldXvohriylt8sUO6CnmzRRCiT+
TAA5t+dWg609a7mVomuaQzesL1YhYmEyi6jPZq1eq2SeNWvmjJ9qxvyw4KIzhaiq6Z0ho/fdUqkc
hm+PVdHIZPvKJspEgZrgf8WNHNVxwUL6wFCe78RV0GDiZAfh8ZojAeGhTA+J0ODxUoNOeSF4EKk4
SPJYcobPXod9osXiDGRTRtebCx9ktkV9Uur7Nf/bxN29l9S9vpWgWMTkIWN9Cb1aEzvd3rTYp56/
00D2osXxBZlmw4v9Gz7IZaekISiF+g1Ty4/PVBAg2X59J/hQNVCeWFLVZnMcHvxwdBSbY6bvlVpi
9GtOqcgqDnfv4h1o3fa2VLJKvRoH8HvtXgILAEuk6DGNMjhQNLdEPmJKYM+glzH7SSci2ZlEvReu
qOBZktKf62N/PalNBg4uKaPJUjECIenk4Hculs3jqgmAWPg0ZrepxVrd6v8z7u3GjI7xKdM0Z3/B
uNas4vGDSzWJgfteFYyRnAUQrFl7DHJ5+S54d/O3PSRWCiu5wZFkPnOF8MmTsFx0Vh2mRUYB5r3F
ZTHwBwvnoVQ+O53giZxmJDiwrxd2JbTFpzbSUof5fPpQS6A2YEmoFtcRbsC3ALlVXNOqGTwgWes9
jRpUg3QhYjvkiabebAkoJWZRWpjreUimfbYuPiUH6/3Dmm8CR3LI3LEy8BkjDRmwGCtbq23T7N76
S1Se/kQ4Ot002QRbph9retAVnrGLM0ERdZPjwRG+D0iA7bSrh6m6M9t2WelRBkKqfvM9hvRYadZa
xymaLJsKJru9qek9mJuk3NlAwqhI/L3qTRantnGP668NGtuFD6SqpgF5KZEFJP13e5Av9J+N4Ygz
T39Mc/6/LAS1ciYUk7hNJkQyof/HrC1wS6ZvdjNcPlJFHBuo6mAQfIkOm1ll9SZ8F3YFXEP+5oN6
0Mw/wXYH6gbX1sZsgjH9OhiWgdE+cAWHM+LJbfQjyZ/gn2/mzD8U/3BaY/DrIC0f+K4jW0PfcOLb
I/cxVdWz7XcYRdQaC1WXvMu7DxqvAB/0piJF5AqKE2/TX6AHzAzm+Qa5F1W6uTibeNxaeI2xjby1
9v0xTewU9nUYdecrD9cwvnwBhgoUtTzy1I+6XNq9VaXP56b7fyzMeZ03wUMiBSWP2EkAUTNa8/h0
uE/ZLOzYryHmeGffv0JIiochluZ+H8QdlgqiKDMY2dvwzBXZC3UPd3WeMzbMb2NGb37Yy6HclsDf
qTYK46Y7YfaNVVSyYousIIwsx04m+VvYMfCPTaLM+D8nMcm7ru62urowKpr47dMcHNrD5A+wYSdn
H3lY4yZStvOqrE/li+WdtYHPjroNHp5QMWNkVxMgrppA+Y8l9Tis7n0S4ysp5M/G49EzJAfa+BuF
OMfBLqpNG62IPMyv+RvNRj3G5wDAWFOrCNtS2YZLBEcCreILEYRhss0lr469uDiAnplPy9TJVQR9
yCt8Zfhm5fCQ4B7oiJQCluEnRyMEzsFtH6DIC8QBJAL4tgQ4An+HuNqEYHs9H89+RvcGAbnf9W2h
KXAOmW6E/37IqTdyu8scHEZoJU43+fMMjh6a0zjxyXx0Rxe81HsG0RorZ/qszHZw/oj4orSf3TJx
dmgmy3gAIWRF8nunRFC4l8WFxv9wwtllBDXcu5PKdLy5HPq/Uv+HXICsosFu8naaLcDpjrgdwbUh
M42IubXi9HC5NPtw7ABjnvfyXV/KZYBq/BP02K38NejYNGuJHC4GZDrNKmkaNrPPISjD5YcuzS1d
XyOXU83FB7O0xh8N0OoC48aSUpR2H2g1n0BKxxPsJTqOIijC6S/uepuU3tNf3R1I1s1ibWpPUIs9
j8yqnqAAbnu3XhWr8hFXopUooHzoRgGep4tnSXh2Xgs8vVl0q/Zf+UFfuelvSJojVoNmCT6H8FTu
3y+ykHXomeyZ4Q18i6aXRCeZOVmVoS2DVCwAmg1RMf27ZiXG14WIKBSURiCgDsNTTk2ldzzItOF/
c2Zqs4AWTvRtkKOxZiPpFK3chQU4dgONl7AHmaOWLQ5JbyYHfFBAsnREPQYw21+i9Fh0YQy/2ZH7
rHGw4N5n2cS4dF2X2emhJ0BWwOsOeh61NNdrBenNgsV+t684Mf8/jzw8yaMvLePMx5IP4W73hDVF
sWr5FJlACR8tckOLoKV+Wjq3LebF2L3b64q3jG96HoUk0Mq/bfC47BMcM9G5q1PFWi80xR3uSz5p
V1e3tGnGFY8g0GvYZ569fv7+woEqfABoxHqdEiOjm2RLoKnOQmJ8sLGVMMiNBfMCh3sP+83aai4U
Vf4Lcvw5AWTI53B25fmlR0vPdLESMDqP1wq6eOZmjXPKjHH4ttrTeOsoOM+h+GvJqcpaNKOyXxM5
f3he+plXeaoGBGkTxv7Rp4+TCfFYv/sXkxNntxgwO+znJmrjO683nURCOe/QIzU4lT/qKWf3DzPr
sTC8+uiJ7yxWCReplyGptWeRdUHKNGKbt70njxQl66ilWbcNE7bZl0nkjWGEzM/ADVdr7/ljPztD
ayVs8w+2fEMjHWRnGVZJDtKLU0YoDiOvLqLG5Pe+Lkx+D97XWglyxCUw3KMk14tQUsS7ASU71aDx
Qv1ly3IS4sXWylMyTk+rQHEjzOgah+MwA/LYlpp4uyOhYHeuWW9B7XxxNhJQ3Cj2okzHF4ZPrRwK
ZBzFZZirLflnOMAhVzrcw37s371aeXVr5PKQXalWzxPGrp+TszKFDkfB5UAQ2eAYf6ElZmXbYiTZ
UzOOe/NDoEck7I9jgK7o/bCJonFqckJXYYYx7HBKIbmTTfYo2x8M+Ag11MpEw1rXN6T5J/OxVowv
pMzZDGJV2cHc6QQuBVBtKxGI1M0YMHUSXzAgFJaS9zniESGdyE+EIaViKTJI5Pn80T11baUQIUj4
sut5/QIfXpF+6Tje+fZT1F66vs/nXnFMkKroJ06kQOq0rmGsTwyzLaDUuIndYo78uL2ifSShELbk
EKqRI4VrpdBePKmJeJjkbc6iJZk6cGPEr7vS6PeIKSUhetWh3PHHQs2xbNG8SkcpqmQI4L7nyIN/
LBEmDHsaf5Rv3WJpdrtDZcZXGUW0MdtVLWgMV4DEWyCkuNKHUACJ7aJi9wFWwXmqj+/wr/hG896W
X5ylCe7iuEqxx9Nc5+zLahntCeEyOdUkl0LSbEHjJn/xsKbLdK1NAlCPZt+zNE9ekva23uAAG5ny
RxBeT1PfpIw/wCwCyOMuOIoRQbp0Ju2sNU6qo5E9PQL5RPluIf5PqQMEGa+JnI/MObnWCNKaGN9D
fPaB0JFIgdbyX+W5E8gg06JJMNwf/j8fzE/LgdSlFlLhnl0kJbZlJdO007ASeVMO4/J47VCezSar
yTkTeCoYEyAG2P7V1wbo4alF20EAM7S3yiV9UP4FNE3rMJAOyrCByLnnF2XPAo0n3yWHgbFjDeEd
JI+/cMNPr/Y3artQmodZ5khfIYpb5JZDJI/i8NX0N1UMgi6wLl/D6MNaPpPOJicE///snoV6Qr4i
9Gwg64Vr2XIZwFr508iuEgMufj4s9qzM/bGDgxQo6ZzZVg34g+tiJGVpwz6pKjFyTzTpS9TQNBLZ
WWBqvuHNsLy+PAQ+DMIv+p+f+eImLjMKoUN40bEDEC1qpr/dX10ao6AhySi6U4v6hzlSqoSPovR0
zh3zZM6YELtALAAeROqeKapLRxR0/CL577tTkp9f05ZzlBQ0+ZaN7zZBBmFrJkSDk1rxE4c8YEyr
LsAZ3bRiDqcjyJapLSyuUPwjVdWM1AR67NHnV1igNDh319/VWwefcRapmTeB0OKyXbe2gVwnALVV
XHIcEAyGPMQmzOSWiGEKBIruTjiYstXF9yf66PDAsNJJkoOsVNO0J4j0cpkE8tgvmKIC4rLF7qGf
KOgTiyVStUbrUyIEx/yLgO8uq57ilYSXJm0PtS6umwb25ULgM2WP2AMwAFc8rIqILT+iIpW9lQVN
zFbu8AWragwtv8P3/bT0Jz9qX5Q6f81ASFFZMiQdBy4QkUr3/Weo4T0tHAu3Va1hpCSZ1BtOGtTx
xdOonxd4emQybyMI48IV39bvVq+c31JyXpqCo/1WQ6rAZJHop4ixEtg1v5b1aP765Z9vOSh+E6OD
e3aijL5JfyHMQIWcGNY2fdGF50Gc9oA0YXGjWcdZa1XTb63XNQFY5rWJh1fJNHo6loElhaGNL1mb
hg2qng51ENE3qW6sv1PJ9xdExP3FuN5qMluWeWFwvsoy7evWyQHmPIouI0NtpqjsYCUnvWD6n3i8
5cVCF6KZ03zfMqD/D0dvQVPf6El8lTxc+3aWVydDgmiUIrCaIyQxEtuYmJGHOPnkJNT8gss215Gs
cEYt+BgdvYwmA2mJoXz5b02bL81EvqXUrWqAbJONtR8LazbXlj3fB6z/JlbKle+UkE39+2X+HheB
oA5yN2rvDjfxBHq0oNF70HVbce3KcRUHNnhNGY1v82Tx1MHxE+QlNOLrefurwpPqdFH1+dt9f/4P
MhpO8XQS0TpCsIFkTqyb91G4PBHEXjqW7A1wm/7zXdb4+SGuGOKJhT9HrFXujiK6suQ9viy2UJFT
6mmZ+oonOO50LiwtWXuEc6PCO1hDi0uh+QCjn5oxEZU308PUQAlhubeTrblaZ0OJxpFNFdB/GIr3
JDFhiM1Apm/UpoYhk6gXnSu8IvkM1GUGiJCUihGP7Nd9UE0M9ln523uQYhiI2NAu0uA/mB4R7eu+
7D4/41m0/gViTz6yoDcCvJzl/sO3C7/q7XcW9m5+a5LuhpojrkEhgBizkeJXZAnWIEcprxxLKr+R
eHDNmXywDRG/twubpZ6Y6sh/ja4KMJFJvfXkmTV2wL06GE9VCyb2zSLmweT36J9kC0DuivvYlwKm
z4kq+HQ7gKShJeGSuVn2NQ/pMiM1jIsbfknegixfmTzs2cM2+AstqoATkS0zJaZJK/J72sIrsEKh
6lxYq0r7iPP4sZrCid6x21/Df5qddRL588t134TPUur4APubG+S9Xiz/BXTIzp3UnEPQNYHXB1B1
23l5qOVvnfEodF7gKbQ7tZQNQ0uUJWhIwZUppkGtrl44yYgMfSMPh+73Cc2+R49brr9/mV0+O0tb
DR4Mb32CbGIlmSJNTR/M9sl4SmcssNwr4rrcVc8kFvOYhWCiP9veoxYGCFjwXQCxFd0W8gLoHTMI
RaW//6VnezOhrLiHknpgXoeKCnG45H1jOUOoBESzqL1sQKqd9eilZChpdpP33k/RgfZVsKoEqAuF
++A0NgWN82yDIzlwRgq4Sh0jILed6MxJv6A9hM/1dtZNkO+bz1dDCLHNYB2n/bjX7VX2X56sf2pr
o0CmlujJ5vvlaJzhAAntse+u2OpXdEZqDKS0/F7wnPK6q/lrqhR9mo0MwaLGNiEZE3i1J2VUxK5y
RK2a0XYECsROiWaEZWEw0mJKMVbZbcq26OSjQQdvkzAhASngBpy7cUg7W01WZUgXTvhTYWJmAp3r
FldbbZwOSw/EDj7koKYYH9C6UdplVfCItBxMER8Bc/L/jOUr5Iah9RGJk3oQncv4kd4V7pktwSio
plu0U8xKSM7Gwuk/YJUEIW36Qa9jFAMHFRlrwjc1mCm4+USJiWoxGepkMWxuCKON+8I8wdlF5g7X
h+VypqcAneukFf06frMc8vGL41V14gN1O3MplS1CMTqd5UsdPx9uZAMHME5pN/1vIXRq2npMweOD
bcyqCuco/wTzZk/k1mS+TblhKTrpYpjS1pJZNxwSX6KTjqlWKkZ+oK/fwGX0Qg6yXD+RRdBloEi2
y8layGGANWE0NYQJg2pNiqMaozm81JRE9+u5GNQ1/T6dGE1uMw0GNJcUrS92Zc21YvCXP7f313ze
C7IcPWy8HUFNbj+BlKYczqZrg1CgCtOoIVttMxV+eQD9yd4Pdz0NRIOSawTCt5BU7eqlnFQEwK88
bJmj6U8kaLdcUOO4vfggIK5Pn2UCOi50C68VWGHVJmdm7j9J1NE/y0msvCe8Iut8WzT8jvkQ48iu
ZmeJAOK7Y740oc1/6XGr0V15E+x1sbq9fghBfhP94Fgfe+9SOROZpwKt18cExqapKMzUngXggyzf
XDSwZcuedf9B8ZZ/tIG0x07LhpQHaqyczpMNumKGjYURUp7mfybEJqrckjf+NBpu5C6LNLLG+MuU
/jee7mWNGaEl0XlYpQWB9blcbL1qDwhvWaJ8JgCg3SalnSJr/ccok9Lz2XHsBUryrwExFaIHhztZ
yY8NpGmMUC5Yrd23NQU78oIAzMDXYrM8SyGM6mESF8ZoaxDVrbo7ig7n+/eMHtNnbrIaeRVFpv+B
VoZgkwMDIJ9aEs+aWSjNUvA1IhLVFG0CKX8+ovP02MZjixV3AyFP7Ywz5FoVjP55XBEyw/7Hua83
NR9Ammlin5IivyIUqdfAS2glsgkZjaD0nUjaxW8mNrPlDs8ZZeOFPxklL0rbZF/vyU2UTJ+ScLw1
/n2eKVy15oYWkQeqUhqfN1G9gKEfAVY8aYmJj6gX/TqwfXGfTxsJByFsb2ZWiXbpwktDCmYuAnWo
JhrIXbrr/Fb6+zcecEIss4hTmPT0b3TUBGiYOCiH4yLvaqS19TwShCG018Rpen5+so3U1+FJfH4D
ERUf1jaMd87BJgZYMkTkbHd+iakswqgsYv34nwRGG6gc6dzOodKTZDwWaEDfSmRxRhGD0CDN1N6w
x5xSQ4axMK+PRkMLb2qtYn+mUrDi6k7pAL/1TUCFVLIgj6FIYLWMf+Xb59P7bUhobVd/4CHTKMYW
sZVfkry/DbiArAjEgS/oMIz0DhmNoXmUEArXrSM4xNxneaJwhbuMtd4+obuyiLCsPdPldr7spxUt
tQnkl6wYOwyve05xZu8c0I0piHhZhNUCgBEGaeyctleZqnZm6D6gkBVXVtAj0L7kp1hqHFT8Dfug
+dDs+ggcVzyPXo9aCrG16Q+Afy854s84cQVoVp6YjRueOAbnzqBQAyOkwhNIw4dKwmEt/EhC30yj
F+v7RCizu98tT8bRlOKn2puCxluug+p6M1aPnT6Ny+6wdz7S/jIqf2DGGerlzdVf/R1vW6+KfIou
8Zqso51IdEpBJR27/lOJxmCd7JaZE3oxQO/8c9i0luCg4R3AnHLEcepSXyFlQeW3PBCVxcYydqCH
mFWDX9rGtl1TzWCLxkqKZOgr0Bva9Z6rnAfVyHyocG08Oq1Nt/6eWQg+E53HmIXwT5IteQsQBQc0
70owT7qR4rctV4YUDcTrMlfmiWDlXYj+MQpcb5E3Dn+ibV3snwVyQUJwC2tDRruL9AHJaVCViEFW
v4ajg+gBuwXPqW7iBuLbg1/SDYCLsLE97ToxW2VIo9QKvnsb2PjZQ2/+DjXXpM5HfJBI/FIyakPR
LU3YP1/gCHEp5XMlyHKYV56c15V+qtBR+M0pwg13k7FurADj9O+st3Dh+AHWajSpfV+2MOOJXYhw
1P5QAcrTdcXL5bXGvPmzN03zNsxtky6fZprAZ7i82MeaKnLOTqR7G66TthloP+MCqgERnFbZm/29
/W+KCB6acWmQNeoyTSExAb86CYs3MwMFh0VbYAYXqe16fKfcB11kuN10TGviujmyrNPv0GbjzENu
u9kjoRVkXeDxQLy1UsfCPmuqMRGRaoEiuyJi7DZjW1ISsB3fg4YvMhnieTeYnnH9gaFd1JyCrAjA
HqPAGMF2O05kPluLfIyI9Lf/J8DZH7SogD7f/N4moPWomXNvgxvL5/E4hqdbzQ4skJSA4YrhtzX5
4os+zXnkpBXm83QJCxG436tUQs74Z1wl7BTUNIZWW2SmnRlJ0H1TyGRFEaPOt/4p+5LnA+IFKDNs
rdJY3VdsqXyCw+MY6eUZztphC1ho8VVqLB4cQ/4iWZg1r8aFUYWeI40Tx2PcOMhFQDrbgE2hRFc8
TWbSg3ROLsSU/rd9WXHGWyWtiS1SkbYB8DKKTF+d7MdC5w/Fe8ZHsgt+niCCWlRLnQ3xswuCSOci
3Hy/npwV4TPI+lfUS5Dtbg1yDnK6LU2kSYXiF59kENWEbPYFDgERGGpjAZk/G6UMbz98ZcJfApPO
9AmzFfrT5fzTUw6OCey1iENFxfzkt3BxJgmpoEp/Iu5qSB7GR1bwivSFwNy0YtFsOobCIgJY1pE1
bUtHZqBdgcUEwUIICY4F81SeHqpT/ZYQqOIdt6Q9PifPCtKujUvcULJ4cEA/MIBPEJ608D/kHHGU
EziMlGu7EPpdVy2SGBELecw/HnaxXUjpuVJ/sfJJJ+Ssg4iDH0MQbnNgFEKh06UTL59MSIUYfzgb
h+++fcls9Uav7hbdybxkaSgTr81JMGYqizMD0gKOXFHp3KwDmYgoyfpJbIrcamr+r9zMKDjfzvsJ
dbJE7MnvV5jvjIFJRarw6/BcM7eQp+WMhK34waa6ZDLXYHCgjNTNGCYuC4aZVmZ8HFo5ra1KVyJ5
YG+OD6oVhrYWgsfZIVDmJfGc/1rl3DZPTItt6Wo1arjqqVaozFy7GxSezlBAzOHUOJBwv4a3fjuj
KSgH0fdOWZ3QqdcHCeFw/2DYdZNV/RVfP4MF96XGaDeWMjwZGKQNY3vvRBpu32OpoON4+X0LBcGh
Z29j8pp92gNFtjKx0WyDM5ka/yUebOV/xLeqrgiSQrBLIJo/+1qu95jkDz6BJ4iTMByAXaPw5xYt
y1HMdsHSqiMO90I6W+H8uFMeYsxOKy4SQ7xcIbp9WYKZ+ypI5/5AAc344+ht5UD5fvHDu/Xx92ZY
eph4j7mzYB/J2EkAMLPsEGT/GvWqBSl3ii1bL3D88xd29JZYgH14kQ9ett7Mn0FQkA84MMewgwiR
y0WM+LIsPN49/BBsoLTfLTvh1dhjleQcVTMcpEubOlTkCOmBJqKI17+YJdXX5WpIs1PS57uzG6u3
LwJOqQCw4pwWFRDAUGCs/Gmny08qoOrkWPzqq3e2z0KAXfBgsyP4oX+p8RoyBfy0x2mXj61ntGOb
RayZGi1rJstI/TEUSIah9hhd1eV+y+KOS5bz0J8VpJiBIJYCN/5drNRfU58MjHa2NjBSAtPIMX2+
PFXrqUzuOwVZf9k/IYDDO96Irolmi0lNVQ8YPh5hM0ZiYsLMA3jvQPKBFi/3LlQuLn6Q0YdR3oR5
rJlCez3PCE7FJifC+woO+wrfoKHbI1g/KfBqnYn4g8385XH9WC8NtjmxeYKd2NPL4kqi4ZhTDixn
o5s6Uf6/T0XZKAhwyz/KU2V+0IRviPDZkdlJyjk/eWsW3bb43e8z0mz9Cl3aY8ZZnNUcyIcVpIm8
ROvyOwgSeldAksBDxnm3Zhwd2J3GHL9AmOV2bMbsXSEglcOuuPFScuO4S+QZotSyq2lgFCaCPOBP
JKZbR+o8UHr0ikIZayzrDBZ848T6AuiqIT8NyEtTvAyHfsZXyXQjODd4sVktD8plcjX5
`protect end_protected
