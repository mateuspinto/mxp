��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l����������q򊒆�
�X49>OC)�GM��N;s$ZT~�ȑ �f��t�#�sX?G��v���]G�;N�c��Q���0i@kk���WG�o���8M)�V̓I:o���a�7,̀HZ��o��a%��~"z�L��X�/^>���[;b�bv`Y�3�"��G��aW�������1o�^�9/<����;��^�ܣ
RfS��p/�a��b�&����|���������sq��>��{9RF��m#ҋ� q���*l��6�:u�k6¿����B}5�3�T�ʅ��CQ՗�^���|��p+KiH�ʿ�ap��@�]LF`��b�6KT菬㋂��H�t9 �F�L��	3�xm�9��-7}�3�5���&�t�qZ,��H��п͵�DߛU�.Y#���:�1���@VFv���x
yg��T���o�G�lK��u�Gя�/(��X�:�x��X0|"�FP������`�SH�x�����B������5�M�������]r/�Q�� ���ط���@���z��yg(#ùRV�ӹ��e��p�!I���(OeQt>�Q�,�c�������0[ ÿ���C@�L��Qps���XI�)l�C(͗���λ� ��ǭ%�> ��D������p/���W��xe��g�=�) �x����F���	I�Ԉ+2���QrX�c:�3�u+@�$�N����i�)�z��k�A��i�F���]<4�ZX�t�� )+$s&(q�J����ܰ���������6uP=k8Hl���M� 
+��J,[�P���}tT�Zl�j�u�1,`�yV�В~f@ "���Ή
񈏺F�>C0.�@����sp6_�^|�(���y������a	o��d������#�E�E��@�I�K�Ͻ�3��uZ�Tk��_Z�C1�o��L���1���X�Z~(.� ������,Qh�
5G�گX6��0F��=R=c�N��`�{o8��S�ɡ��?�|r�|8��g�_�S�z	���&�Цx�`��Ȝ�ֵ��Ѣ`V0b��I���:翵3�=�'k��
�M�9���l /��/���=�F`�!_K���U��/�HM��ډv�\���3$�2q����L�=��y��U���{�KE��
��GTR%��[��uc�I�3)�ö���dsmS��q�]�Y?��0�S�	9@��n-�6�n����<��rsj��1�j] ���v�(ŏ�o�l/�]$=�z�8P�ד4qX$괻�,�e��z䭉2��ag����H�^���g�O�L�'��*^u��u�.^&�Bt�~�_ж��3B�*���$h�w*���6���������a;O=/�*�Wl�k�<YW{���R�[0��
tt�V�y���q#��Kt�(�)��Y)lB��ܞRċ�%�VэI[%�SS߹cq0j��*��x�!�d��>#%%��(K��3�\���X	�9JC�_1�E�yp~��C(Ϭ��!U[�f=n��UcV�=���O�H/���`E�b�� ����>�yy_�%�㌌�Pt�z9žlXd�:55M��t�V� i�̭��	l��M�&!��Wl��*C J�V���H-�)h�;B`�^��7Y:n#�U�C}�0�=eH�����SU���!`N���[�h�񛱶����^5�F2����Lv|�h��6�9	�܅�v��B3;�2�[��Wt� S�V8C��S�����)�K
���aD.I�	�NM��<C�{�^�;I�v�i��"ɬ����`(�M���5��X���W�K�c8Q|�\B7�`�>B��Է�1���I���աrL��`��ɹ����E���D�~�Φ!9�k>�+�o+�IN'p�^\������i�D��w����'�������A�ZeKc
G1r<���%��޾P]D�� ��
��Ɨcu�C�oi�d(`�/������!�+�5��+d�D?��>�O��Κ	�bѵ� \�ز}�襥��I�MV�b#4m���� (	#ym��/������Ƞ�B㩎�5$8J�a �ubJ���I����� }���OŖ�[ņ�%-*�+�`f�c��E,�|90
n�~�׈�gڇ�
��:��g�:�J����	}���=�bcA�kn�
]��t��(���C��(YI����:	ػ��+���;^m͜z���b4G�1f7#o���K�6��������]@�6��kO!-�(��L���E=�(��;9߹P��a��:DS¤�0��W���	eSG	x��pO!��mvf���`��:�d���w�d�4	\���� �m
���A���w�����,��Tj��~-�2yǃ8#ރ|��9�n H�#�w'g�)QW�9�RГ;H^B����p���A��n�x���t�Qa�z�e"�>y�T��v��)���$����Eސ�p��e��Ū��jx���M�WH%����FD�f(^#JU��*T���e��Ԅ|Z���&����'� !�Eq�
��*>1A"'X�T�j�V\��ݏP����[�����C�Dd���][�pƿ�|�|����Eܘ�K���!&�����%d���b�;)�t���r>��ɭ0��g�i�R[3E�M��p$Z�5+5�g�jt�% �<�K���Քe��P ���t2�s>%�@��٭Fl�?%1\MW��R�EM*�K�#�B�%�P��}.��B��#z�2����_�e2L� HR ^�QgPeRv�_��c���~��кZ��xCҔ8C���A�p�?V:��Ld�K�.2��,ޠ���c�{����X�#ɸ�)�%|���
��<�\�_&��f]z8�2�[nP�������?�p"�p�D6>�\Q���O?=� @`��M�3��k'~��Es�t]dK��V&<�O��`Pԇǔn[�p��{�Y	G���8g�p/�oBs�
f��[�� tw�mz'�//��6��D�u:i��f�ؒԲ�5岙g	[<*�������^1��M�<B�"T�)&	b>��c��Eю,�Z�Ķ��J�("c=����_:���J��>��R��Z����R%��I�\�x�~��#��Ǽ�����\���x�4~�î�@�q3�>0����H٬߭�s0DWrm�+_�h�p��jP��i2[Z�5�=�3�����wl�P3񋳚�f�:�FE�v�@H�=[%�Y�l\��j�W���d[R������#��{`�;a�S�Ǆd\�.�ܻ(M��vH&n!!��Θ\t���$���D"��?X[�|�l6c��=�$vX�> ^�)[��4�[��ܭ.!,=p��ø�H�9 'k�t�ކJO����.TB-����t~Z{J�0�f?������8R����q
?tEb+���ee�ڨ�ލ4A��.���q��uS�`��RLM?��HN����Ľ�<lS�'��R6B�M %ţ<r�	�����uɦ�<�XmN]�-�Wf��j����p ��s��a�(�(��Q�)
��E�����?ů�o���0\d�yl�Ү��ƶ����H�i,�r���?j��h�;�B��>Ţ��V�?#�pQ@�������V?�Q��Ͽv�s"����
?Cj�u=cw^�e?I ���+�S�8s+�SzNtP*�uC5�)��&X���5t�Q�Q�����I�F_1�9gNɖ�e4
E
�曦��'Q�c���z�[ӄ7��EB�����O����8:���oL��MG���Q������D�� ����H�&`c-}���'��bk�R�IJR��jٿ���m����Xk��QvU�q�
K=��~2Z�#E�G��"Ѕ&��M}؃�*O"m�U`El?:��0���fW-���<�裦P� �&���ݞ��n^4��u����u���LV1x�I�s/��Z��ha'5}��QP��:�Z�383r�mf*�oH�Sڂ7��Qv��Bڪզ�)����P�]����!x*�M��4�-}c���j��j���#T{�cɡ!xB���H���"��p�F�u=��=�f�( u��.��G]3r�^H�"mY�QX�qU��^\F�ډP� B��W����h1V����|�s��c4@Ѩ�A�Y��` '�k�K��iC�86�iDj��f�|F��f����J�&=#Dʧ�CU� �O���	`R�9X�}F4T�)!=�SpIH/�P��Q-�ߩ��bk>�mj�����>Z/�a+�%����ş�v��<B�l�53|[�v�]�<(�(�1��