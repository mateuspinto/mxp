`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8400)
`protect data_block
Jf3FOZ1yRiLxDURFFp53ZLEplNn4CHjFYDHseXgMdgwdcSBsjjCaJJ+xSIsORINOi3YWvbMYGssb
/ugQy4cta1VuOMkpjEd71oFmPEY8IHXKbk9noQDeT63nnjtQBP2LmG0iQyL76yxLAWmTRTw7sH3G
ncYaKC+GHXYh7UtkL76oJnjdZgro5P8CMDlF5zGfQPAwpeUFlTp2vmonog+es1DV/iaAYsipSN7b
SZiMpZ1IymsMLOnnebdfGg1nCkawHL7n/JL0xut9dQHIAt83uHNdoCmF5onWkEuyKzhGJmrW4BI7
gTBuc6bENbLBrmPcE8vem2ZQvuA+fprxYRncABb9EwBcc8PoKM9XwMC1iv8RVMeHg4qXixOiXx7O
6ItuRG/Ch6LPVsPGSQxpqxQw+AsVs80be8TOwl6LAezpVbLuYbkM5EKBfuiA5auBYbqKbu0axXjJ
csq5IzYRajk5jXT5Vt9/LIm1dII/8M/ZeUzTuUhjLNr+dxJ1Lf6mobcyGEva+oMhmwLqUPwX177n
WR4v8uW7I8LlhrNUve4BOBMQg1B6snQnUiHqfA0uqaz9sOERaaWE4Lc14YWY/vpaAqFkacrHjVea
RAtuycheu5YKVes4iJFwErKT5LD9U9/GZtOgu+2O2bDl7OMgb0dqmrOmBNk4872G4e89FSkrkMSZ
yuVTj4kM/Iwd2a1HX29Yzfxmqjw+5dZ8iNdsqMGPufQ/3XokMWKcOvDnWmdaDpOTlqUwhJF9rPKO
2c2O6Bjc+PLyAK1s9Da9LbEeo3Kg3tccFUTt+oINMtmZ6gvNcHmjmG2Y/tPexN3dnqt9oks7GgDb
rKx/8IUXJmkACtKiCA+JjSZUwFv56wyrgG5QkI4pELG8xIZ0rrzPyK5o6wRNQ1XhSR39cxc0zZ3d
EDcuByc0sgqVO6UsSRV/tYHUAA18SM2UqX0Blsq0zeNnP3WEO4y4UoqH6rpS0G/2UbQ83zttrsZH
SyQYXvjEIu8MVoIOCzZ/LzmeW6WjOwWUU6lE+4ZamzBrEpSURuci85tvy/a6FJgum36aw3lBzcIk
oUB7kIvVue+ZUwhZSDsPbYSWQt/AJN18izKANzPPzLivyqXevE6bIivPe75QMvm1uAoHRuD+4T/+
wxTfBhx6t11c6midmcLke7Ilq9zCPa1X+A/7nVN+k1Q6yT+WMb85UBHPrY31k/B+63bIe8W46+y4
oanSTlWcB6r5Yi+Ny76hXk2N8nf3MWWzr9sucLVlGqmjIPN+LXWRFLK/H+re5jGrLG6yib4WZNoL
/Os/cRVyvoiJEighbZ2XTqngolLw9cMuIQ2353Yy+GzbzApdslBj6RUzJ2WGabfTRRiV8GXsiM+D
jZtbUdeyNfal4UjFM6z4zJIrV6lNmqBR39/He5iiqcLGFBuwm5+cHPyu61GvadJy/NIkh66WQS8b
bYUONrBdRFLkNmSDNYxEWYeJH1lgSUUtB+GeSgoevc6UwjtoprLMWnqBsaef/GXTRrlmtoKC1i8g
tiVYBRrP9sHUHHzk15wkXXNt6jTAVszbpNpEQTykd+Gc8yaWn+7wDtnKgEybG8mfi/MGErWPGF9c
IAiJrFfEJi/otEzf/OJvzHr7CBYVze48kSxHDSJomsIYv1rr/jIxKTcG6z3mQ7pMhKRIMVcx6frS
IHsrD3tfEjw5W66GWThYwj/nNftd6BaISeuomwDiF5U050D2EHTJYmI2JjbjV0Mp2ZaxhF3j/BxR
N9Oaut3CuPGjhY35bpuLfzWH5tUSXj39c9ngoqhyGcCxYkUb75xK+ocNZRsYtuLNbcE0iYxyRkbP
KMLFFEGk1oMRdKU6Y1BYAN2J4a1LTgUpe37Ay6znMREmYbGtL/iHNuJqX9nOopPHOoJX5Oqx0t99
UwobpyPC+hTG5S4VFN3kROL0gdvtlCs+gDA3BnV+EKgb6XsoETrgT05rjL8oV/YYqCBJvu4xIKU1
Lr673yQCkoZyAhjfs9SBVDLBYX+OPvRsln48usTjrRFewQshyPBiIt/AZGigcqYzhx8OanRTCE8X
kIOsnbRLBx7xR0cCHspO8Jo2cG+F/F7rYRYHbu6YiXGyFDbbDmgplwQiUifCd3N1fUqjS5jiuPRK
pOozLg0V2bHuZOk8vW8oDOFhyOmlwvg67NikjFn+Tl6wdxXU6WCL+dEgN5Flfuqsjyl+WWXjzTqL
3CQcRqnx4Iahguyt9j0vpxo5J+WGWXQl205xfUdJDO8ozhUQdPyGAZT5/lha7R9ZfbePtUFPaDCE
N3SA4CdD8acYP7nH9ygpzx0SrX5WiOqn8nN9l3s+Qu/gLncfKbB8sMwnzKVk1cna3Dfi/raLmVOr
61s8iTeEgfmlfw3vZNJ4aW72YuTX6az5oHX+1UOr3dnlXtfm9QLf759p2485JEk6REYDGdmpHaLO
nmHeapF7vimG2Z3HBxMbrh0AxGr6SqwG+YUjayvv8clV4gJJGdhc4f6bAGd/6s2+SJpMF6JFqszN
EDn/aRA3OAmYUTy/PUiYOKvxt3OYi7qdP8UpNfTdZKru0DKFSFkHbtfTuiug4MLIJmvbKUuke4JI
xbwGrH+YkbM4gqDP9tgi6vr18VucY/Osm+dq5fYR4ARg9EFyfrCCKL1tRyxij6+FKt1TvjH6m76D
D6oNQNtwDwtIwutVyC0Fq7KzOOaYmR76R5orpf7GZ0G3ivfDwgXomF3sJ63VTBk5C7TUYp8gmWTS
pAveh4GGq56c84xd2OVWERZ1iyge1mmoEii+TsBvpCtrt4fTMAfv5fNdhqIJ0sjnF5lspeS3U0QQ
b93yLmPYR5l1f5bJx0Y2jcVhM8If6p7Eq1Y5GnzHp71pjMpwOLuu2k8izvK2zIIdno2gBRvrPTGS
rEiBauH9b6czqTWtU8gT458UNPxjP4K0S046/d9WghkEok/oFQmHpR11b0XYMLwmiPfVKsKlXfC1
ej5Pai86fjnGAAnrDcBZYLKKhwwlPZtq6Fzod1t+K5hdWvjwOD4lrLBzuD1WKRZf0Ab+5PWT5qd5
pRbq1IjU+Bq4gfC7oJeP82K7uS4vYvws/Cbl84a7yfCMxY/pYoj613sZ6a4IL3gC9Yq+r2p+gP5Y
YJzzF5V47PsuQzTiVQUkarUisNA1fuvt4KizoNJp4hafr8s+GM1bqKnD6qZwV0/0SBz+haDH7qG2
8OeTGeyLtp6GrSXsb6JEdzU1h4lfo9TG/tO3iiHSUnr7yvSuOpBk7OSR5Nbh9QZGWkjVuu1+gIwS
ao+OHzMHOR3cnTJJud0GXujEPwe1/KW57xOd+YfJAtDDY6bYwMBlIf8M54k3MAnhZmflzxB4na8r
B9DQolfQsKneyvi4aDJvX1/bT/ThYQIDYQftbmDNPpKpcTaFXsr+XGyRHRWg57nFfqky8bmHVG+A
1dtamMyIYjQnBcpA7tFU+ttNTRVcfbQ2eBlglx49fjJ83ZvWuP2r911LnOWHB521s8URO5zx/GQy
bmJaWoEFeIybU/9KfpLQP8xeTx8XA0mYJaJEgMgczMhn6drM+SYW2fHsNbuFZH7xnByxXteNp7Fp
tG2yWuPIn0un8t4zVMHJR34LGgUWMhnk6mJQI5OqjOQwbBAXRFU/e/7tn8zA4uoGmbRjLHoq3y2i
7HhJDdXzPMOYXQq0j84fbAgTsjg/1LnGTBXW69r5U40aXyRhX/6cTd9EkZxoDLAgRO7Adjhrk2hi
hNAkp0CMS2uYhO0uOEYEyJTPpBB7rSzDgzMFjhpXNL+eAtwO06qmbh+OkdJPqz6HmzzIWZ6cZQ2W
bPOtvHfoCVtW7DjuI5NPX1wcd9Z/8ww927xpWiVVzrmR6zkZDf+Zo6Py+wIgYqv2WNKL1AHxzs/B
myfJbvQmkiNHRAzM9//r+MKqKkPFZ+fLKqbwhZv4NuIMqFe/NUn3ev9FcVnENzWdadw8Xr89khLd
c5cl5eKXC/4q7bYVReiDN0OL65KoqPzX+0QhPQGZ96ANrQ4Vd3x7svsxURkjrq9CnXJpgiw/YjBO
hOSsV+ogvnA0ZVg/xNwW0zrIk5gj/L4dPx6NpdwmjLrqLNJj4BWyUtcZqh/Qf4jXa1MmfLmFM8Yg
+s3T9C5G1OXFW+lXaiM9nAEScrLaJcZ/sVEGzWojwap3dGvCUfAA1o7e7C3BU1MznCf2wJbOCv5J
F9ykyDXYsKbZUkjHQFyoNpmK7X2/LUkotAlbGUG35eWHeIiOo1lGuFVRyBqV0PsBXSSeSGzl1cne
2ndvVAkfg83Crlu7vFKd46gN4wrbQHoijz3MFt+ZHRbppnKQcMOy/colRg95ou2vrtah3XykbGLN
cMpqFwCMyeHjdGtgbzJrTcUT4lJFRGvkDgicuXA5iOmatCxW5iDS5Hv6gByBVsOIu+uBI/DO/ozb
D9wuKPy1gf7dLE5pj3XjpuvqIfgQyZsW5+fvjkprgXpQ+M7tXAtZ5J8eGg1QyX0CgJMbW4npcSkp
EaHziljMGaDQhg1WXnFvCqxXFtjEHpnbv9N1edZW4AdyElacTSnplMe5iCL6ivkTU1qRbKhl4+EN
MhzDou9179w9bexOqhz6l4ww2REIEm9R3MAuSfomz8lkB2GffpBz8/RNwOGZZ9uGBKIU7Z5TVRGs
d7SMKAoYF4PQAgRMQtYSBxIwXaqfa3p2AHOURcxgNQtPLNbY2ypN0P7+5usfc0rZherlK8iCADye
F1QAqsI9KqjiuKG1Y7pCRQov/yoin5w1ULNBZbGTO46r2Sa1RsCrrd53a4xC1kzzO5KykqARp5I9
YBWVcTOC92VHvMitU3TYU3d+39p3ZEy+qLqbmOLsXYhmzCJ2Bm1Z4dg7XktmMGqGbKL72ZH81EZh
J1hJjnLgZHqZVInvC7yQAachLRoMQTChytiP5qdM8vPoPnZom5cpuNflh29xqi8Ci1lSDpnfbw9+
uA2qdek3ieYdI+kaGnHrKnVms9sxEmdglGoTiGT7n0d348WasSJWhHQFW1LwYAlskLyIk8rjP7r+
Wye904+GwCIGimDseVthQ6wrvaq6PBXFWBtPxWuzVtO/Z7rQdk8cvEHm+5PlMdiPLqjJRyhsRQff
hhWiSh9AdiAlsDeFXpumoOP3hLy9ORlucJZcqsMtsVxd9BAf/0Si2vkrcHWQw5oyFPIRqScugV2a
n951iWsOp1+nReoUFTTNnz/P+8i9s5Ay+7V7LaSTbciTFfRW1URqA1SCNAdrXy/3qKbDgr5ryd8b
qLz2HtM96NOh5AfVbo6Djf7D63bDNTv8JLXIEJKsN0SR+J4rSOgSYYKkXQ0+vo8HKIlMqmkbagHL
plhp0P51Ue0eQCAIUVsLW92YFF7ln8ezdBAde3iBKdMy3pDzGbaJydMA5b8jmnURivfveus4EBRt
FKsaRSuvIADAf3gZFLlUSK6hFZz69A0hXhOjdIrGfKc8aiNL0WAWhiRI5ZMwfp+fz9iVAOJeufGQ
oXmsWRPtJnyq2Yb0ucx+Cz53i2m13TwHOGj9Kp8XvlVk2Cd5Lew3d6x50oM6EfZfkARvh7NZc1d9
kByP6vXdlqpSOg+/rrJwAtkIMuu0nB5Y2smkuoHasHv/uyG/tecPl+K1lWXXrn78njt/SloQF2O1
w9yOQTi2OqUQ5LYXAN6rlQEXNEawfUq/nhJ0yRaayVOjhdSL3GzY0Pv/AIBSdW/wQGaR/6mYNwrC
UoVuUVw43ipUZd93Ewc0F9bsXr8X2fWXgh09nd3/Jyc+sORemzGVFOcypwQL9iQEd8u4AjhneR80
9Hpz4Ejx9o5iUfWiPLZhKJ4i4TnO9i9tEmty3qzha9EwY1374rPay+JP9NrODbqwj04HSrFnhijw
793RFdjIEcZhRyCYphcg92qYosz2FZuCiNPafIKAtIHwWRzJbuEnysgyLuGrZmxS5Y56C2W/iaNf
Dg+3O9nYUzhnEJzcWif52/fW9MrBU2H1dLJvAibk159mxnYD5FJDmoMOgLrByIAZHNIU8acRPnE1
a9XIaImvIxEj/6rm72LZhN5LRe5Fo3mbblvtXGBjzkjL+VnSh81GdjS5TTKJZ1EBXAqoN5DZpMBn
fSCfRnLPf4KfrGn3xlF33vrYJDFwXHjDAtOJZfVOoo9dqGf7/LRTT1vpyxgWUdssg8ezB5H+RNbK
7GUhgX1Fui7kdFKdubH3haPghucwerhpU7nEoysudaXGE73IuLeFFnAJP0iAfE9Kk6eOvBOVE2ak
L6mZZo0tkk0IzDA0Mp37dn9pgRYQhajyksVwaYEc/novEuApXpgS9SdBoXtZjXDRDKOs7DYWDO3E
vL/b4siGkv2EYd6MGY9Bvxjsg9xjCtAkEG6Y4hmEDQ94wq+5TvAhFR6JZfrdH4/QQfrknBOmZ+Fn
QcLtqkB4Rte/z9z8IvesmmNbnYMg1zGIzsqerYWLlNEbvip1ETHo73dAs5lJQJqFdcHJcTMtY9v5
MPy4rJ1EWNgq4kXFrBNGvP5n66ON/toWthC2E91RzQjB6X0bJozMWBbRs7ymaeIEd5HPdfkqbw48
/ztzBqdzlmnMH0+oxhRJywzcw1tlhZvcAx8h5J6rU7/UOryjxS+U1+UDNQIHWxnxHh5Y8gs62SYQ
gNhPe12AgjKkhzSXJCtUCtk3LF+kitmOo7uFSLqG79sdMTWzQyEt2FkIO1DGYZiC3rvHp5TH53xh
bAsE9uI6GAUJ3ox2mo+VP30GN+uXOKnglGWRqpcVpwlSfQeqApPFg+5YIkbAvHGRYSq3PMOQFyak
daCo8uLFQxmI/iQtsxc3DzunyuU7R/bgAt/PbAzC3PA+/WJ7GZUL4I6XSuPkmDmia2v41QFTxw5O
a6dQfzKlxMCbc2nBkTj2rIA5kdHsSyqY1vKBuBu2irYJoUY5EKrvKC0Jrk+Sx/UnkwD4SBTZ7kzg
b2Ia5H0zz+pcLppSANY1Hg2xORxowSuzEJobVwtZzsfVsnZaVmKro0YWcRLAFjXV16D8pCtD3GUO
IbIBYDSugiF2hUTD4d+53awVp225cfrBan5SToB98ydy6fiTMxVMW4zqkJWGC11PtjnQnyUMLizP
+WBtVn4OdZR7H3GTHmxVutLcdwP97v2FNEcbsF4ggcN2xQwIph4kk6picwlE4zskYvACzFp0dsoM
B3wYvF3tVPLQWgih6eO0eMKa3wDWbXZWYvZkChdq5t3yy9D7RvMxTax2Uxz3rSazPne2C7MG1CNB
F4UuLG/hV/lObJIDVfAeCq/XE7puBYsAzjebXpncbtCN8S2beias7h6laCqLInuQY55btVze0TFi
YZu3JWiDTKgvuira36N1lKePE7w/fcoEUU1FXhn04jDw3d6nRBa7+qiTxHiDqnCU2sHgzyZYnY53
gPGtA2HWnyUkCCJLjHSVg2I0YhRlKzIrHBVQ3q923+V1ePu0TG3+zxO/xLVOTjd+qCuDu+9brHhZ
OEEB7qJQaI9qrimyqhhSXuI7IFpM7KYb9n3x6BO8G/qQ5Bq+CrvwPlUxf/Kl6ad7aQdhavHrbRVw
ySDB9UTZ6OXOEFoJRH2u5wdAWzNKHT7+LA2zfUeRp8JbXIgxFfD2cJ8NJvJMCy1qfobM4MujnaSZ
TPY/7B4ifMgSOsdwNFA9fEYP6vrq3Nlg5SP6o1tlCsEtxLwmkAXVtuYS3TNzfw36QhnUS0gDQMIE
yER3zSTWNwE11XVC3p0tojhApdgqYRsxUTZUlu3W51kA2L8j8jzpTgCXDqYbSja/uIoAzQG6Dua9
GEFkEgFln3ajDyZcsDfpfPfZ42FA9TccpDD1DNHNt1FJrY6R4S4u81jCYi26U5fGT+/mjyM86ZSQ
ZNu8jEJmiRTOwZa6AZ8EZJZukbJeGscOJamXA9C50phzVIVlY3Jhx3LFKaR6h5FJmb4WOPMfcXw+
h6dhQzOicsi/1NIMIDjwWyrY0Rp0Qak/W9dZU+C1Gm8Rg3lweCkAHCnPzE0fmZNlWJshAD7a////
e8ev6fSXwxVA2WfThs1tPLasSZVRf69HrvgcyQHUmcgS6zNwci6AYq8iAczzUz1XIO4Y++9FPTOZ
FnkW/TMfRYzC7IYbxjdAGZYM81F20bymMSt+HKMNEVbm2gjx+bNgMm1DT1YDq6w+aV9H5TDFvpqM
Lzg430ubtE/QKgTsxUpOcpNz8CLYgdn1mGHe4/CHqAFNRkhV5CB27u9EiO6J2I6HdObc+AacAkXM
x0cHmEOY6LJhYe6D/EO1FKvB6jvzDf/iBsgJpKJ7UENip9Mf4qdzcWIr4VUZl4Qpzn6FwvbDfvMZ
t5efkl/vSxdNTgRH6286z1ICa6Oan6jDl2Pm0dHPHgZZceKsrPGZh99zAGsyu3Up+CTJiN3J/7WS
YxhPsHgmaQsB4vR7BtraUVLIYsrMU1ZYgqFtV5tOl2XSL5M/8XXiM4UIFZanEWHZDfAgxDgvRyDd
gaqoGc7362hDHxorlGsFfO36Iek7PiwLtbNTuFmpRxYSHz+Obck1meBLfDYZdeYcKBY7TMX86U+S
18yRpJWtIVJmwskOs59cgFkq2QoKO2k4Jo55RW/8Shj4ROjFEbTig6U/Fpr7Hqo2PX/nSPFEFUh/
fqoaBC5nxp5X1ZE1Q6Wi+aHxPuKTqLaSKawRbqBkvPAMsPEoq9mpDUj8ZwVoxEbiEdhkChdn37oN
N5aRv0xK+aV/dNnqHa3rETxYwtGIlJQ2wZP5aHlepVRvMNPlojxPhAWvHfvUZ6KV7zUb28Hw8ZMq
3a7zP+Y/UuSJWYSOPldKtPlutha/PP5TCvuZE1Xy5o5kLyri0YvAOccf+I9IjxzMeUjKyfSLMCE0
cY1fesWTxljS9LH9fVcoy2XnSMfAOAonjVupEJxQPGH/7kN0w+rAZeRn3f7E9Dv15YefD+zJNSm0
H/1RHulV13KEBA5x0SRvmJMB9rDQl1dGJct61mlM9Haile43CSzqKQAQOEMUxGm7+yofgFwLUrx0
diweycn55120j8IVwNqHmB7RO8mm2jTtgz8t73ObtHlkg2fxMWTpFIlZER5QBrGeygMatgp2cVVB
LqerwEYU8sWTBs8GjptJoIIrCq7q5t1nyHlflemLmdGqkcJ0OXRHM4mlase8qRXTsIxJMYZSV4Z7
wUo46JQNB1K1TwCO+xNflGZ8vuAMxjmVifZlnBHmKh+M9AcBGK2OuWTw9206jQ+A+GlVr/vR7dPJ
1qZkiQX7ibzS6GNo5DDYw/wtkQDL8usK3W7NpX4RQXS+JreA9mt0UrcEsAu9Oe54ElcGhIn30TFX
H3oHBt1q2FF0R9poA2nYtigBKPySXDrM0tgJhQdFliySdlNQGrLgOJg1QpTmEDhq4vM4Pz4EN/8G
Wue8IGXKBL1UTX3rUxR2hADCkT9gPIFBsm3iKzFpkVeVQ2m9zuJ8MHvDjHAei55lvN/F1zX4w+3o
rzjsGB9MsmgNsPAWRhkN+Pe8R7QwHLz48lE31+8fhq5wTQsCZ35qE0harizWTvIChQPlBOXQBXpQ
TOSGZy2spb7za4txz6zfckuPO7wvCtmYorAgo9yLV69MAIgEnARKe8pwcfDCUs7dUgOQ/CPFXtDu
94ItB6+44tnYhl9Rf0sLAdBtSiAPIVIaUnQ+/pnlb8F/rw0kwHxm1vcu97LffHlrYOuX528UojhR
huYXwuvoW5yU2vYXETano/CHCXeH9P/AAjVgiFFHOIs/sg08K/5NfOajhUXACL+6+022Oacb+5I+
u3FgfNZWv1sCBa/OM8iIeGJKm8ht/CUV6qJSkJ6EJo5IbGrsSrnS7IDp9Qt6RJY1pl3kn6x3Dmao
Ni8p96+uBxzimYXq3TFvOmyM1veYbJhmh9i+ZiJP4gov9OU/TKGFUQyip9XTeviTHUbsbvz10vTB
2wsXZ1kBDY40UWvdB7x90t2oLWXyJuZhJHdh95Jb28qlRqOb3yuCGSRBW1PJQ1a/hXwgz35S+PJf
iFZXQwQXDY0B5CNmIR8H7HHX4sfw0bSBBQ7NOFRr2y8OpOQK875/l1q8jVQ0EsN2d0uI8wwoIM+5
Kaoe+hJwMTmLLDSYBwhhUCo1LIVoLMQWFPfMdi9poJC/pA5oGZwnj6iESsexuzldSqoi2cIZdYnr
sdT/xSMYUDbu4X3swo9ndinMPxKW6qgVHy1MAQiw9eT0EQ8jwsRNkU2wfiVvg3/ftE+K2cZ0eHNn
kvDUCl5mGneie0yBgc3mEy8AphqNQ1PPegisDqN6gUiMJesqB94lw7KMgdZLdPRGufdJTeFND0CJ
Dkxoah1EKSA/0lOATwCSWW7ErWyjdqgb8yqgFOFOVQe+52RT/FjW1gEkHPECABGiTLReZ0Vt6FNP
L1bzlMeM+4dnfHXGGuHS6QxGYmkOpU1Aoe8V+POEzXyUv/ykVbIet1dYRmeSsxtCkCKbKzNojvbj
K1cyTFRzAabssxN1ig/OQS8xt7VRiO8DYLmjT+0u9VNblNgA+zMRB9bP9h9kMccQFV/19uzjOhvs
fmUGRa4Ksh601ISKK3Wis7TJPR/pmkoKx7O4IU1VQCb2rRN123mgfs96qvdpCeirlk/0eVPwFCmI
3Fh3VgF2wOswuR0thRinVycyi3x6dUqqZh/2QBA9YnklAxz3imyYMZ8jF8jsYNMRepG0Nu/Mv8QH
tx98fFRo/GKtkSuYhvFhVho9u/M4n8lEr4OrNbZzJ9cWLyrJQRAiP1L+FXairufQ2fE0hLxRBm/E
i9PZo1ewNK3OI0iIVUwm+woY8D4gOImg5xi/sZyrqXmpdIcXvErFY0DJgivRThXUIELTYz0LiFKu
uNmf1zKRkpoE5XOZCU/iuPS9y+EuJk06JS+UODlyck9Aj5nUlKxBEPurIiVxu2y3QNBrClw9iN2g
10yZOd1INtKBY0IORJJxU+Lf5D6RYL5FS8gqEeNELWELGaY1LctrnawhX+XKwsuWlnrq4XQNry6t
FMpXkyalA5rfaxy6rYMjR7hk82NVWdR18ryXhVOYHstAfxXhk9Yz/DrmLnpYviR08DSVEU2KIbIn
hiL77cIutL1DH2LIUHDqBxuwSTyb3lfXFYH6y6K4xBOh4ViN5oC8DPMb9B7uDc8kpnlsSRZjBy7/
5AOd7GOuC5P6EoMKoVZUxkTmbHXj9198khOoas55OW9p3K6kxqQta/9uGle1Idn6EQj8tUH5nBKf
fC7th0zxwDvZEXeWJHBJakdAZ5BO
`protect end_protected
