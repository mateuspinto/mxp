��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��� k�X7���A��y�Q&�<L�`��P93,Nb@a�̊H36�q��OW�ZC�����>�o_�}Fp�Wvi��cH0�d�_�8��l��l�ZYcTDC��G��-�C��X�4�l�4�j����[�m����;q_�Ժ<_�/x�_�ʩh�ԧ�K��Hg1K_�B�4��X"m�vN��)���|��̖q)�T�ip�R�}�[��7ܥ��ݚ8M�i=�9Ht��&����
fJ�S������G��,�R�2���!�plw����t=��jlW����Y|���G�.�X��XA:�R�c�+Fw]ś��rL`�1E�o�c8�$5~��hTp��;d�%Y�*M@k�1���n���:)�U�N��T
T;1�2�0^y	c����}z�I}`�%��3a: w�!��7��]��qoW�{=عT��e�R����1p�ޏ�}�T��|W�y��3���ʑ�}tB��R]w�1N�׈��n��耏p�����}�=-��-D�V1��4g��<��#Z�����5��N�<V{�pa����a�#Y�qoQsfA�HΜR�NN����!�G�T�Ǣ����Ȯ�\��O�`V��C�	�d	|u�"d���6��OjAVJ&�?ʼ����S�u��,�ۤ�͙pN��I����V��&6�Y���n��؅'x4^4 ���~Uњ�5�G�R	���>:�R�Yb��u��61+��9j�+= ��=Jb��m;�2�}�%�2vm�]���m~ڀ#�7������T]W!�[��Q�P	K	��)/���_��w�=��������lm=��4������(�i'��Oi�!4�=*�����^�X��aBH�Qb��WI�����Ȱ;������;�S=��ι��VE�(q�?�QBo�]䘝0���;Z4
i��ύX+w�z��}[K>^T`+�x��3+c����PS��O�l�y�;�c�j�$�C���>�G4�S	ŷ��N{��6�>��Q���7�-.\�7l,ͷ �x����[M_>LS��?Iٵ|�IW_�
E)	\�9&��+�e��Įa϶�*Ӎ�d�M�g�~:�Ҍ���_+��OF?����np4�32�#��T�Y�i��"x��\�ыC�0���j����6SvW1H�>�;�>�I��L+|��46xAr88��p�pb$���g,6��ڃ�5WF�k&2,�L���#'k��/;28���i��Ɓ��UDoˠf��}��L�s��P/��\��cl	�Ǫ!WP��|�$TK�:��P�мY�՗H.���Ѻ�g;�׵����I��k4+˓�*p�%��^�&!��9�Mޏ*�����1^�p��>a�؃����� �q��C$�:F���K��R�r�޸y�,�B-{�2���e1T��^3z�QtF�")U�|�LEV;0OB�my��6>���J���9 ���/[�*B�]6��:��=�䴠k�����
1!�!�����u��q���E�uHQ*��Ժ�|M�h`���$�qݱ9�Oa���*�ַ�:�0��W�s���ͭ<�� ����}v(.^�2��