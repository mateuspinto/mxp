XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Opʧ���+�9��zM�K9*߳��A����~Rt���3s��!:���y��PE�us��ʸ��� ���U�������t&��$�h] �	6�`O���/���입�Y�wUmy�!ӹ�y]����^�A�_��2�۫��Hh�k�}R�h3����cw��;��Pی^i�6�C����U��T��sx�\W���se�uM�P_�2��Xl���(�1z8p��Wgi%`�9��y��^KZ-߇9=���Ťi��C���(o4�6w���.�T���Ь)z�꬟��"`,m��>2�O|mJ��B�m�4������yИ�QXy5�?J���f�F)�5���t �������u�n�?�����(C����A���5�w����^,�GПE�/k�7ky*QKqp�K���>������'E��W̥�X=���W�Y�R��s��j/0Jd&�={���(�lJ;��4���q��0�c8�PN2fzF�[l�&"��+��'`L���A��=G����ڴ8F�~�;��GEg� �@�d��}��'7�Y 1�\�g�Եt��>"xrG�2�U�*k�~G �N�N���(�ϧ��|*wmd���7��ka�p��.NV�V�Ya.$W7�"ڛ�����.�no	�Gd�D�-�j}��+G�ט� �z=��]��<A��0��ϼy���e���E��ci�^;����7���d��O$&^��7&2�����ʁ�4�䙯��d5sP��M��^3���nXlxVHYEB     400     1e0�u3�ܓzCW��@����
ʱ M�AtH�j/�~uj�&�&٠t#�O����V(��&�=�*P�%���l�y��a\��$x�C���{X���9�BE�|L-��P�m�_�{�����z'�^���wm+V5`\qyX1���s�Þ���ᯔM'D}�u^J6(rV£�n��y3K�����{�c&vG� ��3���@9
����-|H(�CL��8s��$���gM���F �v�|�L%�Y?�%����so0�c᩠�J�)?T����
�ˡ���I�2�NM�q��XU�L�jU_A{�0���^�/X������S1���%2��'�jd4F�N��k�:%��]�x1�&�VX�'��h�(_@�	��$��`���H��6<��ߘ�7����m��1����i<x?"�~Z<K7�;���ԡ�P6{8JӢgk�}r	��o�����	B�L��'`�aN���6\�XlxVHYEB     400     140k�ù�	�7�o>��Q#⪉=͟�j��~�Zj2��R�y��|$ai�.��2���H(U�M�\1��"��u�)^�� °�������hv�d��
>Z�w�<̽�	X����:��7��(�6�@�& �S���
B�n�>�ߦ�
�e�f"�4�d�8B�V�\��d�.Ԥ��8CS�y����S	�Z wV�-�*!x��sƁ�R�B5���Y����3k`?b�K��f�ۓ���#��	�R݇9��q�.D}o�؍ F��y����]����&t��,X2�1nQ/���½��&�摥��X�M|r�XlxVHYEB     400     140�˘���K�L��T.�bCwV�M[<z�(N�0$U6J��rfº	Vy]C�tcFܦᵤH��l��'�]1��T��[��Wd3'��>*�w�8��Sf��X
�S��׳�* �N��iy���&c�噠Q�q�7��tP����xz��tk�#¬��gEm��2�/���&y����F��䝪�|ބj]�E��pQ���\U?R������w�Z���!�+�_���\8I����у����$yL6T�ED�ɍb��۵i��$�����`YL�]Ե-`f��'��|;?F"N��VS"��T�XlxVHYEB     400     1a0�4r���Z�YzL��3e�	Cu�_X���͎��mH+ ����*�gva�T�.�]ip�ӯi���xDׄ�h�Co�H6F��]�OU!T�EF���2�8�=�_�#^��s���P�p��,��X
d�=f o�4�p!���.��"����yTW������l�Z7Ih�
̍���Qθ�wHB�X�&�)O>q�[��{+�G���PƎ�?��l�5��+yeL�ַ��Z���j�U�,�s���e��@`�l��0�-��-K��4�S��Ъ�E	p�����YL�m�c�U�q(�fE�u��$���&K��0o�i׆�4�e�sq���rآ7����3Q�{[TIof�=owR� Y����tI
��R4=�l�rց*$q���1Of��Ȭ�/�XlxVHYEB     400     130᠎�B��&N*���]��U��N�bAGu/�~�$���+�7u8�n�Sy�HWc������c�'��pL��묋޷tD��~�ꭖ�wE3A�o�����{�#p�F�R~,�/���vv���+�����#ý��,OQ 	]�%�����@�?O�'^�}9��(�ز�'Q̶��^��l��4���+J�Ӂu��^�$A�����y��
��-ϱJ���O|�͗�K�٥[�l�LCLS�#���O޸'<�KH���	K^z�q�}���M�d�j:�`L��	��(��m��XlxVHYEB     400     190��3!��eRB(r�	͌|cv ��$�����L�<Eؓ���S�̎���fT�j��ů��l�y��ǯ�G�����&���fq�zW�8�F�&\sT�dǿ�5�C՛JӪ�"f�j���&���&��}1o���F�
�!uΣ� f�B���/`��5���۾ƾ[W�3�"'Ţ��޴��^��l�N�޹YS?��祠��݊Nv1
�#�h�J�Z2���*��^%�����J����3��S?,wb:\.V���>����p��m�t�E5�J�4��	]Y�n�(�g��rFT�+~����n�,>�<Wi��-���b�2`*6�)�x����bZ��-߂��)�.���>�9Vi���t	�p�:m�����]��XlxVHYEB     400     160�&5����L*x�w0I��cw�2��6�$������4��q���7,��eX��?QP} '�^_��P��u��4�M
��#����J�N䨔�5{�����-Ļ���&U���<���tD�����9�;��"���|������ox���c<Q���+��3nό�l�߿���C#��=��h�����L��%�b��_��(@gڐ��9�i\��o�ɷg⪱�sAa+�OΆ�+��oF���ӒO-�z�[>�!�o��`?l�\UhW�s��L߷0?���M�~j�Yw)X����i�����O����x���<	����,��kn&|�7~,�b<֡�XlxVHYEB     400     150���!�OT�����m9$��ū�O5w{���X�����d1�s_ϑ���E��q�M:N��a?,N���Eg@�/D�gH��/Ks��`��4��+�þT�np4[�I��vm-X�C�# hZ�N%l�ͳ�� �{x!»�݆}���B�cnL������G����ή�s{	�T�vH���i�4.��s�tg�a��<=���V��8�Jb�`@c�6�t�jc�Q��Iu���lQf��	-�J�/���M�!I?߼��M��"�ܩ���͡�Ȁ��(V�`������^�+ӹ�>�W{���rt ��XlxVHYEB     400     1b0Λ���C�����^^���< ����l�OĊ����T/O��9�Rg?S�3�@�<�?�[��}e���׺���
��&��t�fS�����A\���z��d[Y~G{��l!?��ݰ�²�*�9���{/�X�f=��	�d+B3�EI�aܶN��;�v>��
�*�3is���v�uʮ"#I����v"N���`�P8#!W�ؤ������B�����(=�դ]���j5���A���{���%�*�.5�I��Y3bh0�R�Kٌ?� QO����i����K:oRe��N��) �O7�?Nlշ�+/�,܂]���K�����@����۷�����H#:/)��Ԣ
�4���2S^��D��d�FR6�)��;ݚ�*��~TiHAb�[�J%�8H���q�-0@`�i�tT�P�Dd�˓��z@XlxVHYEB     400     1d0�N�|��u�r��Bd������{[�u�o�Zy&2�A��z���#�D	=�e�Z�������j��{5�.W�E�����'7�ݤn7�)BL����D��݌=;��f\t3c���ž5�v��ڻ��w���U��pZ�'Xg�FS�U#���J�p��=W��@o��}7шd�Lb|a�f�.Q�<�|��{�k7�,f�UY�#�ӿ�]F�����x5M$����B�띲m=8�7tG�<IZO��׷����P%���u��W��x��Փ�
a��?�?�H������۴��T�%���a%Ya�3�6����m^����؏�����D!��3�8��ڟ�4d9��qa��Y���l"�#�*�@[?Ue�TE1���̗5a
�$Q�t�i
Ǵ�c�DQ�y��<'�e�'x��tK�ة��[� �T��	���8�j<x��\�� ��>ȫ��Ot��XlxVHYEB     400     160�a������hJ;�]�c���+��e�� ����"ւ�g8J=S��KҘwZq�!��gtp�^X�����0�^V�_o�3pW�~�+����I�u-�(*���ppņ�}�!T&r"��!V��Z�l�)dl����J	$Qp���Z�x���Ia�d(>�mjp���g��F���@�L�{����O34���3)���(b���{WF�wt�T�.�L����ii���$) �R��|�0���;EݮԵ��gs�jC[�&�]�	%Em;��Ǳ=%�e�U.�wV$u�?uWQ@�w�^U�4TT�"������G#;J�֘HŞV�3��$�!@XlxVHYEB     400     130"z�稯��۬-��$�~���E��I(�����#��ޖ��ȯ��e�C��M�0V�ZTZ�U����Ho�xo'	O�����SlB� @z|&�ߎP�]yw�dmb��m~��sH[(��f[ܰ�}��p�����-@���4��*� 4�7ꍏy������H J�EҷVbN���`�U���N�#�� ���˔bN=~r'W���L��
��D���ad]�&{�T�j�B6�X�����I�w��L 蕳��,J�-6��y� ��TW;Qmͩ����R�Dʁ��;f�*'XlxVHYEB     400     180���t� �#!���A�}�f��1�gzn�Bʜ���,���z`?��L��+�?�O�	2��[�� I����y8m���9sg��*XKx(´��őA�5%����@�R��C޷t�ɏ��7��'���kh@��Q����k{��G�������5>-!{��O���+q��\#���k;{�M�6��p�/eOU�CH���(��<���	P-�=�u�������1���T<�8�Q�x�{2͐�}���D#.u��Z�6d��Z��l�מȑ�}��G��T�qr�f���9��Wcb�$���@E�[�[{�9�Q���.J¢E��Y�f�%��i�cg�ft�}�+��{�cL�z��u��8��J�x^y��n%XlxVHYEB     400     150��b��q�_R݄!�_ �~��v/D-�P��x��_5���>ǐ�?E9wp�m�tcSl�v�i#�q�}�z��w?����5�"�0ڛ�R�	i�����>��mҒ��^�]���w�'@�F.kU6�v"���Yȴ7���e��	�h�g1*!}��`|=S�T��4�Y&����C�Q>�A\w��i���d��#�f��"�I�u�2ٙkBq�[���d�W�JI3F��vH� ����v7m�����*�?�x���)�����G���G����O1��"NW�UF���>\��)�9���}��+Ș�͛����'I��XlxVHYEB     400     120��?�H���$B�m��ߤ�`����8$��=�d�W���g��8�dB��?��p�N���=3�w+�9p��E!�30�$���:[o|^/B+�@2 S�@�z�\%��nL�E	��x�)��ֹ��ӊ��c�F.wy��&�&+�n��dry�qY,����Ux�A����r��s]Q�6=����k�5� tr�g�(�����L���]A���$*�m*�	"�'uF��?�Eܸ���
���^k�l2Z���.�6{�Om����d��Kl��1b{��yJM������!XlxVHYEB     400     100#�X�DR��j���%�>��A �q��.��O4��v�x��7��':AR`<8V�~�'����B�����2�{t^�k>b�z���8�(��ɒE>������7P�B���U��Q87 ȷ(yEtW�b9$��<��p9+kU)D�v���8&;{����-�n./NJ>�ZV����m�tf:_FrÄ&f��ΰ{��]v�P�s2%�BB����3c����ۼ-�9~`WA�eYV᭪fLȹQE�XlxVHYEB     400     1a0|b�+Lٔ���K�z�r.������Co�*�\�r�a��~e�7�`����� ~Fo��\��%�י���!|�c@�%p�s͒��.^���am��o�

߁��o��r�.##�1;VQ��u���U`�l�}�DYrV%���U5e�5����ƈ)����m$tc��ǩx@xq!�������a�I'�T� �5�t�8�V�������a������5<,�W���l�kRDU�����ʰҀ����$�FU�Dl:��� �6���6��V6��{�^�֛�Ҩ�#���/�2�崺�u˺�(tN�g0���ܜ��/���ϱC�HÆ�˅;����(Uw�X���4��;�������&ϣ�ME�bymV�#�nN�}�A��9Kb{��o٨�Rp��0>��F)XlxVHYEB      27      30�q��JX�\<2���F�I�:�"���[x1$�.�Q��7�F��vK