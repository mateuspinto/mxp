`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11824)
`protect data_block
hHkJVdISy+0z9nio1Qjm/IKCPXiauzrBCACXtxBEI7PALCHIrmIvPq/NyyZ/1NrQmN0m/WM5H1e6
HCHnoqWs4uvd1dq0apYuNtQYUaG+tVS2stmn2JFyXsYcveplhJW7gVtQuohZAMM8K4N1BjwiD8x3
fReyWDeplsIkcgQh5Zy7DT9YopDmMhjlern+2sLDmZSEBeBSL1cTGra/tveM149Bts962dNpKstv
Xp3DXik7b5HRAoyDv6dXh4oMMZwSCNSmc6P8cyCeuZLJYM1pPu6o+JZC0LYvopPkFrVo+0qSnRK9
LjdCY/+aLFbA4W+HLJpxFWJn87nZnvspMb1XphO7nC7tkaufOBUdRTe+z1T1m0oGz1E/SgvVC7l5
23rKHQLwzDho1zJgCSKYOKFASLCiI2rM/cVDCalIULymlriXPSOaWRyrurNAawjUaojnBybXaRJ+
jwlUU0mz7Ejc/mGPrXyHftdJdgES198am+8mKjs7Jk4eggr64VE7geiVf9ikMw4Xat9Gv4xY3zMz
QKIEl18jekUfxkzTBoSr7ab/MG52seJ3OZ6LnbJnie4vxzRViAYwM4m+nTn+OmcZ6GpuYmzXhg+/
K1epW4uE5nmRuB53SUmLN1q9gW1WmAF4xJEYaq0IxL2W55ivLcnFkAQUksDu0OBpHRynnyMSJxNL
krkPPwqu37uJpdNr7ke0da9K43J3TquKjhTDvnmMpfXCpgAWMjVH5GdwWBHopwPSJK+N+GVvvTWG
mo/7Gj3ghaCfC6t2JsCrxHEKfawjAyu02kZWFnrH+2nvK2Mnn6NU/86F2N1JOkTDNBYpRCV6kcpO
BZRXKhAIITadf7XRYT65p88yuphpBHdJzv81ts/eTxfteS73IKHbQFx+6eDaymjBkmImeZ6tjIn9
60BJFCuxnYompyjkH507pecJhZoJ1bGx6QbDV16W8IcuS0zo8sumGWs3lzS0wby/JApqoO0C5qbC
+lq4wMO+SfiDNDR9JnB7dGR2JK6RNhbMdXDVZ+UHAwapto5E5I6G7f3MS0baGZ3J+1FIZeJG/bjf
9WkG1hvscXNBcdqzjPq8SPcsy97wEt25JNKLlTlm+eCBMigLO6X8q5E0Kuvhnk20WrFi/EoNCIkG
vRYajATpVcEjC+wjdfhLzq9mmNLKvri0Ajhz0gmI6OM/APsa3BdePlhzgSm1Es6PVdf8B9R09dmu
2C4OXYlfrVT2WlqUnfNWQ5ctGaBZwknQ2VWU6APh+O36Yhf9zn4KQgHbnoM3bCNsmh5V5RUZ4Al2
TbfViLO9PUW25XzgFvH5vLWqIIq0hcMvusGmjz97DTbceRVXivLFTZZjBhRSzzqCtQKG5JjpWX3B
itqen+BZN4i5WTxInuRjyVQwuEn1attOnF5YVyEJAxbhrBnSMoJzWCUYuwj0nTGW/9Hxz3UnG1DI
Tv2nnMz7eDfEA3Vv6ePLpYXLwQu91pdpR2+nSu2YERVwmsbT/SV2Dhyf45JmjZY4Ri11DmSC/0SJ
8EAWEptRXYb7djVCCAeOtA6Sm7P9bSKSGf5pFXXOgMikDbcX0rSsulKMWgYchA+MEErVdRN6S4Iq
tHBltkxC2S+aw284Wc5RvCGAgNoZt6Hv/aTi1waxcww5WhidjTzjgZ0vAoPeG/CENNYRIVQjrRv4
6hmorad6JIayNRCr1USoHiFS/eBkELvarmYooMbN15tMExK7bx9ZFHNgu+17+S3JP89VYy3Owl9u
mnA04/1xpdw1yurqgp7Puxez22cu3vnvzt7wJ5nXvMlFjqQFIw4H+A7cBIR072RK2qE7NH7XMcdS
c+Tk1FvdwG1ip68hH99VAycbfVl4Tjfqx3A9TTRKr2/fjmn00+kVVQ3GrEXoLQ6ZzQB+QJYu4xSt
pQm+5gmwTL40UL4mBY7qSX8Ph/fCM8jsjY3hVrYafI0DNM5JcA50WmbPJvvjruRBkS/Xeopi0vb3
quz/X+eUnEBjtlFZIlk6jKB8T85wqkuOpO+2vENF/KyuTExqWwbOLNpW68iGoKMR32mQiokwXb69
d0GG3FKQ0s3nB7huH8lfsVjXNoroJWIiXe0YorjHbEcxcEshFamFhhKpFBZzskpP1pLIKVueafFm
Drxf8OGz7yU7tQv35Hr+eY/8kJQEg3w7hHMigr6OpMqM6lu4sJSBhji8+hL30/DpRruqzOJdgcCe
o7BmfjhEvas8uhjLvEiRzaBvzlifxhYkjJwYVbHuMzDwIFCTgdgWe6ZyqdcsKWkQ7StzZD+c59Wc
xuilXwjcPowAL4RbsYqbW5Y0qnN69FTQ/YtjIqwb2AZNAJiDy+Ut3QEPUSiulFat95/b5k/7XrKX
iqsjtXLRuVg52kE7+KZ8gXquESlOs0qHnGvhSxCUQHbeJ7sAO36KOLwN15LPE8lQV2BDxqeSYyuZ
aA8QQyBnLQdc6j4T4Fs9FTEH8PF0QeFg8Es9Uao9CBpFodgNeCj89rKxqLl0zzR77FhrMxUhc7yn
A+Ow59nxR/Qh5caztbiCedBrisnk5w5heOGXxWrE4iqNfEPW5OX2P8HpaQO5+WvWLzKulhh89SdV
wEzICpPyIaht+DrgLJDWS4rCjHLyj2yzG42zKTvH7opFTs85SgWKN/ODyRMXUlu+J4vny2GUrRIF
7aowzl9NY6KnsecZPXXH5FaAy4jwj9MfT6rSQCPOzpPanzFcRZ3YIF+bokXjqkRImMFgSDWuVszq
Yv+oMlM/mLXp/9lHxH3x1pgKvZ9D1Xb3F44Mq9IFk/v+KSmykgF65LyDHPxJRWsFxc7E63e+VwwF
Z0qXMWBtFYoy+OE9TqBZkc25riAvAN/BizQZpIFD5WjZRhJQ0rYQ4bS6ESNcs+MhnmCk48z1ttdv
8dhuVHMy8nmoramir9YG/2rYM7G1shbWrrdOoZ6J+zL9AgKs80g2hU1YPPKDOMuAMnLctsgmkOGB
FA2w8BI76at54zgBd7XHb9Yfn46GV9dBdZ4YICty4iVIu2HXKCTg53h1vpv6VoC4ip5VaEf7dGVo
xCq4KDNd6w8Iwqv5EbXW2e6+idFG8vVmWwLG2nr+LDgPguh9YjtYaGIY0PABM8xFJ1zyoRFmzTv/
qLHEGw9dR/F9Gy7QWLhvE9TekO1KNzxAGA3aAW505fsfXtwJEAnKgHW6TFvgOYrqDzmPTJxL9ZKH
cWV5ERkHd2xDptEkeBN/rHCVoJ4sd3enMgSLWJgJYPFCDVev3fTa6xCxV6p2ni+kQZYwhs1JHvn2
a7nAq6bfI4PWCqUI+v+/bZ3W9PQ3jKAams+hvDj2+AGH/uM2HfLeU6GUGnC+ykR+2LMfOsitsmrz
TzhmzQ5QYcLPxrM9W46mxrT23F7QY+4r93tMJ5Miy/HiuIDmByoOk5qEXho1bvR3XmSxD6D+Vuca
rjsOqckKbpZt9+toYzXx6GdpHfELo/IjFAYiz/JY38wGXLzPJ2+db/8vIOeGR7lZ/GE4igJcIn35
MfHxvCe6meHh0HisRX9ky5vxUADMcwevtIs25EY4QA2K+4BvoINqdyC18FQzMXgSuottzukWWCDs
5RoacEgOAd1cCp9iMQXZiXYMUvlZkI5dErMtpQ88UxYrXYLXH5L6EJL5TQFZqPpzk7BXprslH8NC
EDriVCNReuHIaO2OQeP3PfL2w2v7uNF45IpwvKcAGkIaUPeM4qVVLbbfu36rCM8nXX4cY7tL4vg8
oV9nT+nTZr8O3Tm5Dm0EAgUG6Par/Qsipr4B6otjoVh5tI1/PO66OCTLa0j44O0UBKU7OeGLSdXC
7dwYLTxreQtsjAO+psjcX1geBfcMADdplLuD1gilpIsikxFyO5zHfq7ET3wL844o5M/yPgkez4Sp
SmeWp5dcEUjaeaYiWsKsVPuKj45nluiPDR12HfwvtVMI7snLDloQfZu1/GEcEx1cj9nqTjxTLyfY
J4z18DJeAID1lAS4XOSumSUwtwNdNi56aHejZgjGT9uTYeykbAYGX0BzhLArZAjsN2H4fLcmTTCP
G3xS/v7hySFmgZIe6OWWfTAQlJgdOuwyD65Rbon16rx2WQtTekQlHzHmKhKbrQFMgr9bIOUhXR1k
1a0abU041ElQIagfJkqJ3xB6i6SD4fjk+dMs5Ox27U+/jBgmtXXyhQR8RHgZ7ourj4R9ZUCtodXD
Ybvw4uczQgPtbT5yNGVzm1y57SH72KXPfhrbNDGSph4ILdeVAKTbNGzfNzJip7mob/t7sk4Et00n
QrLv4cUSwU8pgkfu4QMefKHNG6QsZg+aSCIl7RM0rDzAEa9bx9vGnd11D31pfIo03tjw5cNabYMO
rYZBzvq02a0hnKb4bOADWEsMyntHV8S6yhQvyfGjrB0Ho5VyghxnqkOSODxigyZNKAEqVM78kz/R
S82AZWfJK8s1TzOPGYVZDlaXEpUg/9j7C917XBaLQpD6W4RzfznV8dozZ11PM1AuYw2HsAjhY+zx
RRXIoOd0yBlSbLqomgWpGtoR3ilE18DOJtbUSd1hxwBzW/ZYkhrJdsjJhZtqvcXlReyD/GmZQY7E
Yd7gRX/yIuu45FMpC+WZnFQSqwgT4QuLLnL09FRhueYfdr9dJJWXrO6XW7JS7dcfnxGbKAKVaxT2
pB8aOMZn/IDpzXr16XciMQoN2oYAVPGXEbj0/f8IcDnqD+W7nduJH01BMWPwHFb9ZJPmMWJQ5NRl
kz1Cq8gp/p+gs9apf+BqNbWeMMvbLML/XMb0ZcjVpU7z3UIT3erJfU9VfyEE1qqs0Vzcij+GHnZD
csDZoeaKQuh3CqwI576GhYNKpzFK/zpdaX5Nh0lq5uasm565xmi4QkVlS1WKjEIS5pZGM3tZMG46
J+IUsJdfADvnSzKSZq7feocHE9tfl0s3lFxoFsJMVU5/tH8M6IwAHyCQFkpJED2xqTy6546GBLrW
bItSgnFbk/IWwZ1z7G4QsSfaAuSd5pDOV234TWqfAB+BZGtmXvSe+eSJSWEkD1cg/2iC9JsN+ntA
+T/SmR7DHfqP22vUvIYRTuKQ+FjbwklFUpyrjLzDjCy8ZRCnVmenU5TMr51WBqGbV2+XOlubvG6V
cu8B24DirGJHw1bUdis5Lpk28mxUrZQQDELYEnHFUiDdaAksH7Sg4B0hS4jjGE9sH3br0sLqNabP
WNO2ygKE85mDtKgu+Yl9RvWv1lkyj12O266w+XoveBqPsFBoeyJ3QBKBuKdEI0wNkNRV3KEk6KNz
tOupZGegw7ikE5+l2Ye5+aCZtG6slMTaifz0tmGD4nnDH/7HVCYILzOL6n9zdhBOGREg720qDO0I
TBtFugxIsoNA58yEOKJ/4yW9JH+kvOp2KRrsf30efyPN333kXE81tmSCfyAStDNX/XmlmuEic80e
TkoHGkGzGi8NJQIitJehd5+p11M78M+3dA9uRfo1gsEr7IG6HDFaXdYkQwJ42cHfEhTfly7F3514
Rq8hWRISqcSRFRNUa9syn0LpFhCVjEcDKfV+dcGL9qjjeMTqjv5+6Rmq6bQIJt18/VoIL/ykZrWC
EUp7y9j1/FsAxJVXV5oLZK8io4ktQnDEB2i4O3EH+FC4Oz6OILpXAXmxEXNdZaXu4VOAztKcrt7m
3Nl63WzeBWaFeVVtkL1tvcDZZg/yDQ5xDgo9yDaeQQuHZNs2VU83pd4WVh7A5nik4r5vY9Bh0kCR
0B89WNDfEJy/HQESvqXXA51NOvZemgtsjUOd8IXWvFM/vpQl5dvZ4/SDRu3jneuEJ42Befpx5wlg
smsvMi6Ry4dhiF59mLw8HigYZbb3v8GiaB/V2CImBwnwV+WDIerGba2C3+EwVQZ1R5+Bt2yh6VPR
fJKDZEYUPbmiXEAFEUTiwjM2I16HLgIK/rlgh128uAODVZmHJUF/ePYVYFfBit/gmA7smpiGTsPF
+O2Dh+lvXwrf+EZIETeOaZm0PCqogENi+mdc1zUFvL3yd8VwbNNQ9XPvnEL5TYGh/Kd3hQBt5uOG
bu7oNf2aGfANU43CKgmX8yN5OJ7fEOH6CAQkYD0IXD2bSeAI4RNcSoigHIwqcwccDeYw1zRHA7k/
MpL6MaUe+fsZsEs89bqRun/n6/I0udD/tPlYc1n0FoPbmA2LhiSSK8xoPlRhtJQ62bLcn7Vzxq/f
11jsq/3eDWD1dcUMTpEMKhDFasWfjCfLjUiOKPVWHeru6KaydHzdw22MTKP7IpHAkjUv2uJP/Wzy
7XVEoB4/zp9ASnQu8hKuP/8EAhskvouZo7D+wUa5hz2imJZxfE53ZOv95R3bs6+pPSohwrfrRCkZ
V/ClkmKIy6BsA5ZrmMc3zES90/GSiaPE5uhlF4RXKcivKqdoVjEoCF3g9WbKLA2NysiK5zKdJe0i
IKS+fINA1Lv9niEXezt3wlqRqlf6uVypEI1POnHrB14yXl3fYWicRCzHCmPuFyK+mNdy0waBb/TE
POYSg6/6iWqooQXqBOzPX1qjvfV4SFs1U6HcXZ8sgfnWe/H+ZxtVQSAMJmWdlzMi5RimrLTY9Bts
BKLJspECD1/XlYZrIrsGAvOGNXR+XDpiy+h0QMf9MJCu1ibzwBU6XsxYY8K+pERMgmScmWGR2VoW
fqgfmrzIEiqWLVo6WGQ5Xr3zJNHn5DdnDAX0vBwHz/Q2tPlQWSX37jrZM/XymFPaZuFKiQ0IGuS+
VQCiNG3K9tjlNtmfKBM7wQEPgLqKnBxLUHevz3gNtsGGhP+0apKdkVovTI7IuHM2DcbrQHUXdVio
6a/eJkhaGTEA1o0oCN4GRE0yEksK8iyt80n6q8NUxZSvxeDj2zENx3RkKMnTc+kmoCG6YD963Bpf
Qstdg3QvOLy18zvbYmerZdaSu6qKinc0ijgsBDG2Xqy1dLd5C7h2+8rawyQcL98nwfJQq/cT4K92
qcHgz9PztAEKsEyFU0ulAXd8PgoD/LCvxzVVDnAoUI6cGrgh7wJqgzmk7WVwwsLtSc1f6Y6IWDVh
PFPgLaBXNML9V0lKGIb6ki7pvg5SgL2bYoMFXpGFC1O994i2gzh+aK2J05pCEtGY22Vs1FgUH3oo
41mC+inCL49zyofA2bCdxBv04csOHCg8NpH7432Y/sL0JMgc9IlgtPZAeacDOqNAyxHSuh4pr05l
8BwgtRh/1FE8yNypH+LQFxnvVqWh0FCn1R3o2t5+NVWPSrS/z+HnIMubcmJHNXJZj2Mx6Tnshpfv
ylyVJmYFx/Ubju0W1W3N/ayJF8AvUeeQBqOqLg6WFpX8PbrZECSaFtcNsQSPopPH5jSoHJrSS2S0
1yO6byuIqP8f3Pqdz3XEorjBcgHxxT/JvsJJ7jfjxYMpg+o6977Nzz/MU/n1Z1N1oNFIHSpiqfA6
IaIRB2MamHp6tY1hiJMJDJDNrP28/dJ1qwY65FOvzyk0EU3MyCmYte6bolkCwD/uBkZUWOvQJeDt
N7zJi0NCTfJ1BznIBnRONXdsNH1xf0RYGo77Bky1k32talN+EckAJf8xhElw7dMd2NljZU8ybaE2
GT2h26wfup/XndfsXl1Vz0KhjCX5/ypc1Fl2FntFmxHmLCRXqrIydKizZkku+WcMtRtprUFukisJ
VOVhwxxzSwLIHQKrKLu93zpc5G8gQ/sSEq6wSbWGOW+DBo/6l5vFC/cyHdLs29EYhGzrj7Sbmv/6
wQSl7X15HQhY8jsZ7o78Xhl2ZMD9Vp1ARSsiolWKeZj3M86592iGk9PjRXwmMfH35wPco287OODD
VxUqJ1qfkKbDtKXHwvU/4y2SLQ8v8ieJ3dbsUUdB28gJsVR60VK/agkcMTsaUvgtNsyhuZQAMf3W
NaXUvOyaf7KV8e6jeNVE0ToaSpgfpCNPOdi+dKdJl5RR1Q9UZhz8z7YTG61Q+yWrkE4OjMFxFlrq
WICBdX0biGDTimJK9TEEqIPEpfZBZa+0TTVKiFt6N6eWRX/SoSPQ1iaj1k/fFdljquVt5fJEiCQD
ySui4zO+z1u1leN3tGmS9+NMcAoVSiw4X4bjn70i8r1BI67cbDmWSMe2BwbiRf3OiDBrMFh/caz7
vS+m8j6OF1EqrwEosKCJCVFG17O+a7HgsVSdmWz2DXGlByt3XEs3uiP9+3fo2PCGqd4uYErPf/tP
D2BLmjlOiaYkBdsGVXks7IPS1dyo1LIJ1J/dbxAPrL0apTxpR/Mcx0crNFCTh3Ex1W6pj1UcbIbz
/AWIeU/qB/iJYCHTWUsMg4HqCFcFRixrgB6NijcBFapAp/Cv9Zdbm+7v7TAoxs0QRczChld7ici3
jV3H5kLHq3MSo9gwXR9qv3JG0w6A3LCreZtQoDsrpkdw62Kjg9RWzMV9I6OG9T+sReYHvvYfnVjJ
HzBY326CW3dmoD2pK1vYfEoJySVYTh826gCuR7CQfCZyUc+FirklPI4bDfwndvZbaUqIcXs90L4e
GG6BCabqvCicdo/ONWBk70/mozS2yv1cXMbkMAITBnMJ0gQO9rLUFQjyelfAF64yIrR5sMFHLy1N
rpZRGfoHBNVj1bqMhwllklOf4+CW0Cvwfqm9CSRv3ExI0qPUfJFkdu8heg1TpwQPknbymFq5nwk8
DnQ3cgHoOsMF2xMkUkzuMhFdgColWADVx6X3yBxy13a6MVuVcijFV9PcOcClhOlkp2Vrn54XE7mh
e73Aj8UUYJ8eGeQXfmHSi87WzJ1ACv2lJCGZeQBS028UHWD7vC8nE6hcuYnwYqexMDCNRtMJ7j7q
peYwfX/fIX8OqiDzEIbUflvuBFl6R2Fmn69LWaBCNkMxTHPnsDeR/3m9u1t4URMX1Ss1xFvBYg5L
Qw3/q5hfwJo7HTUL+hlLu219p9rcWqNeeUG+3u5amPlVur3AAj8ZcPUzm2DSQBqy9WEbZYcsRWzO
VSIQk7muAITD3+JGNvf6xVOrSRjMAHnyHiHfbCe1HxcaoLfTt8E6ovSuhRvBw7aQfVJmFKUy6weS
BgAmdf/OwpLXb5T8GOBnfQKxI5RxauJnMqxpCwD5W7zWkqmLer5SqbEqWksa3OycnVZ18EwfQDB3
+9SynWuh/BurH9UzpTfzwiX6OtCgCnEM6KHeh3lDVJEYkDqmuhwMz8/3lY2Myb8ZK6slv/haVFHV
BhtqquVRMpUiUnQ9JDN5UzO5kgP1GLBtMVN70x3DIxfS4vFxs3JhD9bEFJoQEwQFloSFhbUaYURd
WnJDhdyP5Ym+T4ewGwDq/ul4obP/12WfzMKblmKK3utxkyaWUoTGuzfzCinPTFKrhM3QQtzmf4FV
iYo64ii4cQmRbKArIm2WsHSFv4rQEkKn2/TIBe/aKHkDp4TptcqTVWhTpgmVgOHuBB71ghQRZF9v
++7DglPst9IL2BwX8SJSMp4IwtzQK+FUMJdO7xQN88l0l1NlLuHRP0VBLKs8HyPI36EWcjVpeuWX
6RQ+X6IWQUnzPdpye9rV/RnDPopINEPw4uF3NRIykNyfVM+JZQtLFhf4UtBL194m8OTb5Mwx6D1m
jQoJC7BClXT4JpChnXrcotENjpVeyRCpOqKqFW9JE/Of3hS7PrEPfhzUkkHvfCSALtpHtlevLycC
gTt7QaXRVuSQ2y1X9fz15TJR0ESs6hP4RKjbDQ21fMyiYkSS/iO4k7YuecW0HTR1VInw7AYNPG6q
0rvmnAN7kbqMxH890LYrG7Gy71tcgtUWhPV4yiCRTAJdMAG45555A1WIwUVeAQ2TMk6PfOLHU91y
IOCQPJF+9KNENO3L9pz5dhRnU3EW+xr3ZA7JtZGAObctU+j8eyzRgEnF+SweSPoNWwTdwJIBsey8
7GkatgWgwOrARVz6ReHBD8eEGoqmjFAaneY+fnHbh/4O6pVzbIaDSt49tW8ljFuTdlOdc7rMyZeu
3u6qEjHbUQtSuWRpMKykCJAfB3ZD5KKqDXnUhclGHgX2CGGMAYWk0muIdMHuvWVN72pjdnOWmK5e
i2vcJ7m+8XWhKwska66nFRgVfj1VXsoaM3rqG/zaAeVZ7WYyBh63aXsjB0isup0h95nbrBCUleHG
48AQ8vq+VkixeXrH2hOUXfqef23NZz1uxChcDrKo75fVWvaPfmg64V/jN0dEoodPsITrEFH1AeRZ
avm9gAy7Fz9UpLXybAdayasPBpE1BYvsBDKZNLCxkTFsiFvaf3EZQt0EeTfFgr8mxS0dlQKJyvue
//PAzG7MKV5hqrFSwkCcDixE8K0nWsWvl6vcb8OFB7EDt8OgFLUIud9e6iiLIDkFluTvkOLy31KW
q1VwQNiUE7Iv/+K80iAcchXfAXK8u734OY8oS2VMzFGmNPeXHmNpHzfhRVG0fO1baZtDVeJsvOkQ
mE3yLAxLKspGP/OCFILPiKYxf4m6YgRq35A6nR4kmACQzSedWsMBGeSg0ee5AIj6E3PLUn/78opc
DHahJkuNGjev3SwFGRXOK5UtTwMRcEQmbFfO3WZ9F62ApicxZXrZ5DxnS8XfaxDqsxnR+zCnuy5m
DfzY8ABrvrx4MiKtqDJXBeGvLZ/XDp3EzLJIAtEbIQjZeVHUhfmUBCGNTo8aFQy7bknIklZBPAEi
Jd2RwPRPT6H15GTN7q+brnCRY0KuHU09BBwBud9iN/QFqR1YPIxva5QKrh94gPPiiBeJIKLrNhHs
W7ZJUBqLGuuEU+Zy1bnGKDxOv1v1XoObgd5orDkTQa1yp02fXy5VFCJNOgfqdAfI2oLgCEoIa06I
rRQW0nKLeQkLqfGluAtDmmt+hW+J1vS4svdWYvQ7zyQkqlzNBSxsmeO5pPRCnPISpoCR42Avha5E
ERdBnYrWnyu/BNl0U1Kjqb+eyhdqQ0SahqaAJ8wcjmq5zBLkpHZonBUPl+442ws+jm8DbLiou0te
lnMPC71lNk8AFhKLqp0occyHm68hOSAIFa2HMaoV8rVl9Q/lSLb8v6btJ9jHzCc9uMlEWrt6a87O
Ga/ihsWCAYLB/du3MUIc7v7RpdGavDiEeAi16d2vsnHDzD6A/mb96Nqfnu25D7cyHyZalVKwX7wJ
Lw/xy96GC6xHwSIL9a+yxbA/iDavWNrxyxEYyKMyKunzONDuI0a1K6cBLBER2XwD0LLrqo9cdKwo
QJoKA4YaMpmJvxItcEOYsYI0taCADg2ET65s9Eh+hDw7H5daOEdKYLMh7CwGeoM7QX2MFYP/5UHb
sy6q8KXd3NtiSU/ocEgiZYqkdjFqbEVRIHVsiwvpPSSa/X7k5jrUr1bBvFCRm5uZOQOGbdTVz2C5
1D3ouEFYVpYDfLNI/65YnZU8YsGaGfC/zCuRIeb/yozLKZZa6vRunFXyIgFgP/C1CxXG8yHbxUAu
cBjHUXp2RkV/OctK/PvKQ16DbnVurDGyL0l2QyBpcoFihbFP2qDQax/dgtGFmpqrhZd5QrvU5jTX
ChD8K/k96iXvyyx+estGqcYaDaBsqWfbpCqZ+t/1EtWLaSYWdYQORm0qw+LVhYgG0E7HZGnRqiup
G6Qcxlc0I6CnfilTtL/KsYCuGP2CXh348KuiSlaPVKu7pR7iOUiscWgdFynmymiM7J9AJkSFnvN4
p7jRnQMCyMGKoyFZjXbAxYwsPIySH240nBcA7tIWJtWppWUujfs4aWcM4fbYFYHP+W+dSR2Voq31
/tuPQ4SOOmVVXVnsY1U1sBjqBEir5Nt3rPJK4wc1uj5NC/FtOGIw+FHa09Bfijmi7jsHGfk6awlq
u6N/Lz/3d8bpeBSnTPHToIlB8CiKr0KKYes8CbGX2Qjzp0npOxSLc55c9w8WWiI+QnkJZeVTjly9
2GVliRv6leP3bTJFhz1zhGKcd7W4/P1TE6777btu7mpEbMZtNiZ14AIGPW7btQK6RTO+SEokjveD
DY4EzQMDUuUn0rdHEFCCFCMWJRwi+f/RDaCk7pDe9kQiVOT66JJ4ec4dEz+SP9vg74HW6Cx8X5S0
0j4f/dlzToSdldD29SrZpkWJvnUI86TfK0t2qhqVoTN9kLnBKPVfhJ/vHDS/L3bw1Vmzk41FpyQz
QnWjEyWJpib9BDfLYcI+9p5Bv1IrUExhcfNH9UGi3kXOMwNhowBd4LU+UEuBdOAXPMCKAXOohIny
B5b9OxZz21podm8zlsDJwZijWuLUQAEG6ON7zKLjZACbzer+h9Jl7QSli3m7fIsIwWMlNXtUD3z3
NNGqZtmZCXsZurkBHljAn8sC1ynMP7UfHDLzq072NXOGHQdazoxQwcLOCj4hYuZ6XhG1bYdvKS99
tspGIPhOmpImXFxzAKxY8TMG7vPB9eEuO2duCbfxIzezxy+cWXNF7TQ/oB2+/wyTvKYlTIrpQv8I
SEWrsEzZSHsjV9944mBxypnJEQoyJLfcfj1oDRjLuwec1B6OHkcM2o7r2NM03vZll2kYPCtfCk2M
d6g2E8uRYMfQ9MLQtPu3fsexz8cx6p7IvQ8eAnyfv3WHNutOA58agfegH898Iqdnw/mk8JLeQRNh
qTtV2m9uuV440IQkHfQo0IxR7QtBWaudigVZN69XjfKiK6q4KBl+mz/oiuvtRer+VQh81N2qpjIv
ktUmhzHySbU0SEU1ytOk//ng4EVMq6fdQrVWoABeFs4ZtF2bteMGmSYmAHdBxhiTbM/IjKZ83qVG
rql1x37RML9ahE48uDDoXUYsyqCi3x7p9j5I8X7+LtevQMe2X02sgY9BP6vPqQnkyAlm3Wy7z/fg
CEKyre5wUbbKl9k+iaO2XhKX1O5tmJCdCMFvMCxLLMvd3O2j7x0OLBU/UhA+wYbAiN22rnTuKACe
guYDaE/NiKYyUcHCGAGpUiP7pNgVvOJTrugkFRbPhjRAGASyhYbZZIMngqGJp0ocXuSMJtnqEaXT
nAC5KOwamxR1JPsUNeriAdFIJ4a2IIRFr+XO3yVR8PZulWcAjZ9r1Vm0upmDUuVi4ZuiAuXjH6AY
MotJTes82BectpmHDXiLzlL6OXxS2Qg0MVeJttB+V8zGpPInBdNeQylz+x5XChTFyofxo3x0tBFi
oQSV9XPkU1zu4/zDuuSU0Tk1uKix9/FVhBvyebV2SfMOkGv2tlh3Ir0FI9Z2PPLIVcaOSiBP2zmm
XlsfR1PstaF+h0C5eQRrlzlg/IDG/I/1zWaomhyoFrwrxDoNqNs8gEJYl8e/lbVz6589IRHYL/Lu
rLKfKh5vk3aXSa+xe8xkjAmEvqGgTXkmuGfUpxu+yc0YabLys+mGsnFu7dqBKVgB99eXw6mpkjUT
ZRBYIuLml3t5nmL395fsbTRc7EudxrztE/OxaBP4JChhlKWyVR8LnjrDGztwPbGA7in8mqU1duFM
14Uwfg9RSJt7NbI1saOZHT/K0ktbPcF8L3B0E/gM4ALUbHcp4p7z+KheyZSlIb4ZZtc4pIvIwJt5
PJcBdIZ6zB8kjWJwyEhLG7fCdr1Wz0bm8ZmNgB+F+3aH1HEkeXjoL7+SOzulM5laIO9tjDfHcOjy
FcOQK4KTPSroy1kzNlGFjo4eIrgeKEdsJfF9lEfaKaDBWtIRPfs8lndiQpnajJ1Pd0mJ73nFS3ix
Fy0UHFZzvekImYiCm+7Zty2WCkss7ye0GkbqF1TxuSxEg/NgW1SkLtZF+u73qAzz9x3wXs21GLKD
CrsDd4bkoPlIYII6Uqx9hqwjcCLQ4ujxxrAm0NF7wugPpWTVqdplDfjquiplQwh5DQ60DFbJJpxT
V7e9GTeHANW2sDhZS1YUcVV/oUpADGBdp9w3K98C5CJHbbdhzAXzr/n9O8F2Hjqwf64UXxOJnWCv
4gpBvynxEvlyEIhVHZBstmZnwE9Fczn/+/8GC+3PLmiBLZUlCoyBgLAV04p4BMhIgYld8rD0WTkU
TY3t6B7/sTFesJ0QolCulfHj4XkU+GccR48t+uV2lPzKBxv0vvcjXkIm5kbtgUjdbbnb66bdQrg4
7RA7lthGe3F2GwEt9ReaROYf2SCNI63A7gWvJWMwnczvEPacXyxGe+35GdUHoPhdBZ59JKhqMDEu
5SMYh5sNXTtagtxvQDpJv2dxIjr1alBzSoHu/md0MlHxoGU/R/d0/5EZ2pvvjjcC5ShqRdfG2H4f
mtasny7hrXxmAaFbzOMmAtizyGKZuWkYaj9hJ4gzOEjWQ3AW53PJjdUh+AYC/GH0KWiCmNv7+ksF
W0d7CdU49OBV/H9sZ/8sB1kCCCBrC6MhTkhitM5wKH7fudaa1aEoaseYjL1l0zQtqLylYTIxg9cY
o77i66E1srr7S5PNEFI00/fQaBO10aR32dWk1orDSf+V83KYTHKfijsiPALrykRMNCb82+/MEut3
TT3/1Q8rB7V+rUbmte088MPYZAix3ysgBKibqsuhgFrOegLUOjD/40NbfViyjxUYAFK7LlBOHazr
4FxkewcJwkulbJa8b7qeO8J51gNWEKaMJkBCI9c4ffy3DV7NV5fekflPYTXjR2cQp+0r9PBi5K6q
teYQGrIyxe0zcE30Rk2WZXzgMDIR4MQ8q30coNdo6ffH/KbctGSn9W6MFn4cpS7Rc8RzqUHz+mMT
kEgpCSwqms8jKGv55RE0UJxZxGuQ4fuPnxKVFIHHs7rB2V3/rDW1s7pEEaJfIekaGce3cIIgwj35
zmLt/5wiRtWf8IHSp5k7XTE9SAZ9brznJUfU7/2FaB2+bIXJrgukXIvEMDj3Zn2KGknC2sB6Aql5
dyV7Ma8D3lZDI2VeMh1yb3y3hw5fwywPJgKchpAVSEbgSeSTq8iefuJ57tEhvAGsBZ/G8uQDK1KS
D9WAYcJQA6305t+6sSZEuDHFBfNesdSy85toJErfFMLZ1XfabKoLsXDJkEQlFPhYbg6MMso/1uSX
XjUnbbssiUmHXvOFDgTIB9+kp8nRF5YWv/T8VgZQOxXf0Qtt5cb7VjXwvis4n4uQO86YoZCbycNt
yvtya2Ybr1USCkImSdxMl/laWknt7pzBv2tNl9djY35P7rcRc1RPKiTgrIgibUDGDpK+K+tk53HV
sIzFRy2SzYydfIZ02TfUMJTq3iG4F2vrNqSSfiMkTM3ot48ECtcKkkHqRJgJGUkjUIfz5C/4HWE/
aAs0BctCrdSL5PdqdyOqtqjr59RY3YkI5Yn3InmQy81N/7Mx1vfsJJMulpJTZmNADI5mqHQjnDDS
gJn/H7jdoXsvBAwKXeaW1tCGxkPhMZ6SJAcDRBAbzB008uXmmLHadI7jMJWEwZuD9jYBcRLVjX3E
gNSJULycHZmLic3SnCDGyNkp6ZTueVg4NjL+LH4c93CLm/QvWiVvKHyNty6nLlJsE8VfnZzqkRe0
cNbvYAbtIb1lD8yIhMNHuQ3eykVVV0LtrIbTOO+02d4MxBZCZIIzbppF0si6ykAKtrTMX+U9KbQ1
jutaufSvugmHmy0dCkM4B3aL4hr0/vHACHDSVHWxt/UN7N+00R0oDiNP3YCbuu/LSLrIEGHGtj2N
IDkeR1bMgLev2Qc/pUjHI1swC00sKQMPJMQeiU9rIA6zJS7Ocs4L4l0VrKopQ6EhBFMvpfCHQ/M3
hLxshjjd1SdpK0vIc+Ukb09vuRvWAQkVQ1JMEHM2GoV8Tj7JBaKoMgo4KgF3Cbf7A0VBJqrlJcMh
b70tzyJtlHPgEaTeW065WGcU4t/US469FTRGF6r78Mxz8/VTZFiOqVBVEo0UkRhTbbhftBT0T7HF
CG2HaimnAcD4cqfnHLI+6BtdwLZi9K32LFEEqf3Zwkg1VqS6zfRhq/xJcdNQ+jNlD4sZe3+16f5B
ENZ6BM0W1YLbhozdsEa4G8oL10u8AWOwkQ==
`protect end_protected
