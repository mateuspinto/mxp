`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3088)
`protect data_block
1juYLsHmOCxKQQ8+Dtud6q0YOHMNS+MxfjRAKQXXguAxMHahvxmdVz8dmE+yGTYFykxsQWhFkqIe
JljjNb67MKpTGVSIVPiHToimNhIEeL3rmw9RbdvjJuL7wnLRRCR9UZtRcX3ygKr72YvUVn+l2Wdn
/0YWndhwRSgiA4e1uQ0916xPFfqsmrmEe/ZmsmluUHn+aBNmahbXqYuBXLqPsqEkVt2nwLpzCJhX
IwzBv4BF18T/AfyyQJNdLZuIQAtjpoe1ESNB1/mn1OGU02ICY/4iCxGY4CSI8guRCbXUSWsAkVJI
os4RKXb9vVU8DxiW+U3uoscmv3hq7Dry1W80H427EMStuM9SSToc9nZFIfDkgV+msYZdjlN2qmPQ
TDKJ5ho78BHi1rKsPr/SyLljk55xFpx1C2wdh3jdFPAntBdXlKzCkEDKMpw65v327vXYyrYExdRq
pIPlXix780QE46BzQEakYvWAcuZyhLwZysNcdeRZHM7L4thXVfvUL9HwvNzWww5JSXVVP0FPP/1B
4m2fnbtGNnhjyDqLdqnVjuxNp/OcKyh+HfsXZOTgHKW+nZyeW0jzeMwNiElfElYBVhmEhPSh0qNu
p+RY4ku9dGF1ATVfgFd9hEIvGmKkyc4tU0Yn1Hj0LfmfFGCkD9gx9hIMo/7pSPEiw081ZXGMu2x8
BgXrG85B0vHlwQYlAm8rjEEQIqMSsz6u+bkYJFh3DboCQw/N5xmPbiNECgn/EdXllpvfxWM1CYLZ
Sc5wbqBCuje0uK+uayhLmfS6B84uR/HHl7W32r+4+e+oYu9pyTyWIlvqWYTnV+lFLVMmfMTSq5HI
ShftfHNqUTy1m5iRx+w9q3VHKSmoSqGItQKcdTS0f3OztTEYuRFNbEsJ4xPfHvr5vauH/24dAc80
glfzrmijkaSwwJAJKPb+phyCWA9A6Cuj7dKBRmS7fo1O0Zur/EHQSYNydmFKw99oaZdxC7XziB7X
QZ4XFhQ8JUskYJSsHx6rDmajRSs/K0xjZ3VLKf0+V+gOcfHCsl32PvbHX9r1XedUAjdgD72ii5wP
D4nV20v9K0YoWVURLLNhfKT9fDZorwPr9xctHuGeqV7oNBzrflIqMi3T+SnQfPy1RzlsAlOKuooi
iixN4urJFLH47STd7HAToQJ37ZjWiCBfcjQDUq/v5IalbMVecJi56GgHX8z8kSUXx+xWILrIy97a
dvvQhPP+TX575/E7mi2wkbBkp5hSyyfy36wulile/TT3HUTr41ry4namPhMwmx5yjdziR7zWdOZ4
SeC55ACcioEjsZFQ0Tm57jkB6nsYjczGlCAsRYGfL/3wpZnYu3aCNImXQpMGztIDh8lP1WeU5P1Z
JdIlC0OrG5XtGAvgk7plbLa8l6sdHuOahvQTZj/igkufJLPW3q6azU3UiSUskCi+TM5HJivBNJ3q
CPUrLUoyKdaSnj6Gud/jwmWm1qW7zxSR64nI4CNG/sKmCQNL80+b5jBqMd/4B+4VsXDwQxGl75Dv
rjdmar2c9Pv3rSxKPjXleJeXC9E2VWjKQZ8eS4qfeAFEfFKif8FLpGGb3eG1MXw4YS/tFob5oUR9
7QSrzn66lt/zLmQfRHqjAWrx5QYHxy1NXsWMh3ojAXzLpWx/7sGq0awMDGfeCMI/d2zyW+2nOliy
Lahk0TH6u8bPb3fasZ+QNlxMNqilUYZjc3f0Q6jaiaCy0KI//8BWqMHwM/7ilVVSXj7YLv0jBW/j
vWxb+KtvpYh6syCz53y1PLr2NACphe8n/S1m+x/ITVRR0IAc/CU448rnAbJLuK9qXccI4fsEydrH
vzXwcq5Xu43NpBgJMU1vEL+y7sL4dFu0FXis+CkJP5mn0yP5u+fpBGxsQhipPQrnVBgMe8gCf4DA
wYc2kkkfidbwwUcayZbwi/j95j9EGi6sXEZpiAzls24FR7h0oguoVsEr2wyuU3iRSyorGNxcPlFz
iblYLg+y4yhq4dzR+uczc9DS+YMKHDg2TNo82mgTxxr30AC2/pVTz99iXH36WI8bS1lpZQSq5zBQ
bQQiMHsgC2dIJtjeQhpP2zs6FViSl0pBtEKv5+QlQkukFhzi3Q43h2+SgBZxsoZYj0vGl0Dn+TK1
0Sr7DqVT0iOPmZ+7UToJdudpIiApsR8tEMb4MvKaTkDoTo2i7YXPkBJXrMh4lzBVGOVMub8uzPly
F2Tnmhq00nBui9NQBlUEhla4WawR4sG5L1hQi8HRVTaltRzaopBspRQV+rLKycY2TaFPqijw0RI0
WKEXsLJfRbPj8UKR293a4rX5/hNuPJHkMNHA9dANE/lkhOY/T6wM7tnsUcHZg2lU7+kQlC1Tr1iT
X16Pk6vmSpIJRjnLxF787cBk1dwq1iaqL8DwvujiWNe5ahwqzLKqnNHZfCIwvlUpesoOxu+Bskzj
Z7qxJF3m8zXLUfDiDnfzmXoWfJe9BCmckLaEYbSbqdEomYUbjHY+o7npi846KQxQZFwm6xZelp4A
NWNeKpVgipFVcLEHWE5P2+w1Qbsu3HTOjNCZzdagYIy8aZAkhh42qXt/R3vF0Cmt8fKGx8ENEBr/
EVBjZlf3o5We9vb8VupbZvwWxyg61VWg+lktgM3ZJi0Eg/B2Ssx9R1sT6ydf+cnPP5n1XZtNjdnl
i33xHqbhI0XUMDeeI2BLsGopTUNAjAyRpgZ+JABibZTu37ECJz9lGzI+3gs6PGEIGUeM/xlBUGZD
dKTf7M99ChEbwCfaXIJE9oeo2cOj116vK7ryXuDvraZCcHsZyAf11lC05H/8ztVT+ztiNTVX1NH9
CaKUlmtBBW4VTjzcjPbUqif/xfpoEKSNgEude56nwGtHXU4IN1Fwn8jBcgYgHL7gOt4TzfSCvAqI
0WSJ252cNhpnjm5pnCr99p9z4QUwnHpncQWtCTG3ZLvjuTSEM6tGLOiD+0REZ/c6Jhez9Ta1Z+Gr
y3gAyX4i/+lwyeN/qgIaCdkFz3Y3Wpy6Nri1uElCEeHnPcYw4uMZFUnqiKiwUp94JniGxy0ulyA7
ej0cCFG+OqvjklJlQPs/9kbfCILkU6H5TiBPx7EnYsj+L4Vi7zV+ZQq1o2BNhFJe9x46EBr0xB40
n01D48SYNIT5SoKfZVa5jUYSLPLZd9yMUrzdK6RzKUinq7G/fTTEC96HT5aIM1An9YMaAhjxpCnf
JwK7xtNUUw0PauXk727tMBd9+IWDzwVELyUtebm6RtcLABXO42F7NGbW30nuAUoWXgHyc+ZdGu1/
6XN2UTnqWm4mgJxj3Vpe074Ip/H5ECDjFzUAZUg9EGDeQqcAVQfCan3sp3Eb850BCS1jYSQJ0Pel
IKL4WcS/9PHtelmsvWwNekDb2rtDI8FxxrU3q+2YGnfTZhrYS/FtRVDyI7IpvyKgbE1sfxT1bw/a
mzNCqlBL2Kg2D+FzTN9ueBvxTmdmKIZ+y+YHJV0ADujqBY8j7noKzqHeiZy+y6d2+a9CXrYI5GLw
XtWk02tV9Sq6zECyOF10Lhoe+Ku74Z4rZGXKl+WW86qW5qzweJpWCWCL3IsHlsmSuFKhOMY3lg7m
q5AzSbQLlDJHg+GwcBvZ0viuOLN7atoK9cfykYuno9fV1bAvH3M6uRnsw1hXhb5s+TbBB9XxQeZd
jFLmVnJTqAbP9bUf2i2fLr6E4EXiwsDMbHFE865ED4YjkV4xt7yKKqhzHaYwMiHfjOlJVpmaYqWY
VN+tHqLGQg5BX+Ttm1hWYVHjD/of+EsIkbPpxMMM7/RaAanKqIRjgZwOTWlAw5D2dV11iPkvzo5e
shdc2LfaGch6bie5NHMuWejA4FTN1/hzf8woYdHMx04VryrHdM4vi8fdzE2984aDNrnDFLm0FB6e
AdzIixXz7F4Y3sufcccMnv18YjjNWsxkS4mhnWIB40tjBsmBncp+ZiwxL8l2Gyl46FYIkFvMtpjb
cfxPgLUYNqNR/hAc1GNGJsHPTBE/JNmHCv6611oig7NO3EFbJ/URABYYYvlP7v6e5sDn/PxBJYo5
90m2YkxFXtYwGsQ01/t8eU2M/tumZ5hokssMVC1orgCh4lMHkuPb0WdQEK3GGLw7crQKUe3PXORT
aGkHVTKltNBr4A==
`protect end_protected
