`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 100176)
`protect data_block
p0qLiPWW2cGw3BvHFMPWTOegTZRiWVvnf7Q3PbJvECEvfExzdZxZLsoM2AujMfWOeSJF8G3mhZri
JaAfsCseRKmy50iWd8veEV/Q/MeD3SoGQEnpZ5QeYeO4dhkj52APVvAuj5/zkkoYiXNMW/RPvToY
p2qo4qEakfNjoOhtjfKvbt9B9meRresKEd0LIpHS9dQ5o9aYnFXh728k91GzjY2SYmMJLuBdDL9v
rfgwlnAyFRr9Kn+AP4hfmoebnzk5zDsijzQibz3NHsAZ8W5mA0qCry7kK2hTTnxi2WAwGeKex5L7
qGxULY0JSzsCIAht1FJj79VxYMVNCgcCjlmjFIqc+hf5O6IsFIanLT7s32A495Dfzet73w1cEPDE
aUxYqX5GjeeYqSDCDN8jR2ZWZ0W8LgCpepAmwgKcDieyXuZEt4wQuEuP9+EG+2Z1IqQEkqBC0FKg
byYaj5n3vxlJROk+4OmIcEdTSoimoGWkNe9vSG86sdlBIU4p12jN5hUfJOw0GetoJR+nx70lvKy6
HK2BUw2IowQxJQbL8fPpXoiZVB0oS2lyjNeEGoWsEzCSIsGeZEF8J8+S8F5p+fqmtpTsHkll9rnD
siSwl+fmcA4Ht0tRAnKFgTPacZwVB4frP7caYl8AHm3BF29sLd2ZydpuDApe98FKVUN3Uzsudj4A
wbICw/9dDdlNz6L75Fri+D8e8d5FxMff5euG6/NFzWfogMVpIbXhjAHthG80xD4ZHfnC200S2sqN
FcXmGxqMV4F/1Qq1idqxKmXt/AHkDvuskIXnoC8a+0eOWkqVQlgkkJA3ZO/+7txdA2kGbUp4cSjl
c6FJjuXKhGRafMG10G7lc/XIb/6hgfpr2k2722uKM/0zMHSnTzaEcOnz8axFAF1uTcemwbFuQNWO
gQto9/h1KSyiLg/x4z0BEYzGnR7rM1oGYXVZ7YfmrYnfe39hHPCh74QvR4mH7Eghboql2ZdBhBG8
70X5OynF9S4xbZd0mw4NxnP2Q6OTYOitRyZ2JtbUBCRrtSjc1lMReqcUnOWBfRo3vuKMwglnJDCN
UXU/3gGsALNPbGPX3WxSSaxyoPJ3buuZ4sL1HQgOW2rRlRgKHgh3ok8S8s+sWOUcxeL0xRuOTgQ5
6M8BmCfxvUtuvS1zkkybbEKqoIfzjHtmvBopb3f4IccPPsMXys8ET+AXKHz7OEBFjjQpIM/qFfaA
NB5V6QMoVyo0HiJQxOfgsjyl97gcAWaxWs61rVPhrcDHi8271WXT1AhNvhOQgh6xd2nbOuZD3T/E
xDYY6cU+RQRdwTSwEytIhOXWJojDRF5M6psUrNq11NTkj+qpw8hpxaLmlm2dykFv2wkKfoc2e/Wa
t/upfTrEmAXi//PyaIdFhzqb3mndliFmEhDDsDa2V315wwJK0Ojnp6CFagmmsHT2mhFQDl4b81AJ
2kWmuqD4yw0fh1sbq2Upli7r8dvQCC4fqcKecQ1O5VD3wE+GJqOIo5eyLAGXXFGDFtyj7ALNS7fp
q+V3KbtlorCYKK0xF27jU4cjJnXKdx46Ojx4SoPHD1A6azVXIdNsUKcI0GCqI6Y7wkRn1yxXqsLQ
kQiziG/vWu/mi1M9/g3s55kXq41WuQXCBE+5Wl9xax/ZcI8wSWU5xxNIUrXOi+G/EvXX6fG4tgB0
mVRMXVd32rTAdLmpjiNCVgabcORuitUcrt+DVFrt/45932ZJQJWWfL0q772zIW8n9otqx7lpMZku
IyNAnE716LI1BzH+ASIGJ0yK4EKwZJ5zdTAIRCRxEj2sDDw/5av1dogTFssxfV73jGQqPbRiQOBv
XRgH7JELpD814u1A51jWg0wfBkHQbLYNCRMQvg5xJvTaSSGUIBCIt4oRqTqopX6N0ucPAVDAoz8q
R2BvaDXoPArYW04JcFb5Yo0SP6GGOLsBLB4+qVjNH2RklNCaL2ZQSyV2GgFnTTOsHiL/i3GM7HUj
HaWoH5hVW3r+EhnEOnuSIgemFapuHAndr6mgRz+YyaFG64hbGKinTboFsN1fXwMLSVZ+trAhKQyI
nx19Rl/ejT0OvRMQkeBsd1j9UBdHuxsfe0uwwd7R+v6O4TsmfrQsu1LVzjfYEm7JI+PuOPJjtuRJ
JnfgsNS9jEG++RvqlbX/aMCgPvYc+8rjCCt3zsyjV/NiFHP+Jz2FA9qRjJ8SadYB8e4u8A9OMLeS
qdngty4AYOWhnOhlq0Fr/VUBpXUZ7EPGK+jZwFzZIpXiGA10YO4n5f+3nB95Q3NHh7i/R5/TFtMX
l9vKpHSwaE11tvuXQTC3Fyg2CSs+/UZ2GGvt7VHwbXwjngm400j6S3RVqL7gTygR3AeO/LcFZXqU
qsSMMcvSZ6XxSoCOdnIsGhhsxUl6OXLpwGDfvRvbXEbtg5p8Q0EnqI8kosmEeA2GiFYf/OxMRnpr
mif1rknPV54cJQJnKcroDDZ7isoYADd1BgFYxAhA5Bho2aYTnfGz6p13H9PoWrobF4QyQ2aqUCPG
IN9LG/BvUyVSb/haTGpXRkopA4r/mxAO/H/casRZjo64HyWcNCN1YF71Wfz/4oiBfxjrKTZihoo4
aUvtwk3wPNbNPuod9ckeISBesGp9soORsC2h5h2VRlZZAtqKCirY57SSSrM/E7m9ijeDg59UAjbF
/OLsOZ/dTetcPc3OCy3bzcB9c6I6ZQDMJdPbxrT87VaB2GKQtgRrVDLc/n1dNgcI7W71vEJsiSM/
+fitp374CQKufnoRwyOSrK6FqA7CMHRKefNyqnWZkInAnJQkuHVo6d3aUK8J29ov1qnq0X3KhlVC
xmnWG5raBvav2fz2qy2fjQUYwe28X9JyqrGl9kbDkkskqF6GViQmfw8pwidyG3QAPX7+/qoXQgBQ
yOSO+9cuC8fZFA7SZVkqgrCPTP+9XVcud3EPmoIrroRZVrcT9ZdpVifyBewrZ/ZVaVtclaqnocSm
571sA1mK2u+NSvJ81A+CqbkC0/CYD/dV//b71GQk8Syy77YcKM8WVySMLg2q0qBirFCTtc8seCQd
8Tjlf7tGWQj9ic4xLGKKfLV/plqaNh2ns725SypeSXiqfV3Lp5+iJLF+B4YsoLYGbV+sP3uEdRPu
Mo34J3pzLN5lwErXxqGARYBeAsIw5RRJmePNmb3RtDvSrc4mhw1NzKya9fLiIYZShFVglg9LHrlX
EiVaHi8KV0nuTgPCbaepT3mj09BQAdOGlu4IvJz9+oWymCJAP0eLsYlUOruQMyl4CxUIbWkAT4gH
u40oP8Lng8g4fY/Gb1FTSk95SuORitmof+daiYHECMO8YjOdILfFI2mnrlqVQVRWHstAAJfpTMKP
gJnBfkWQBRgqi6UHybNyGmiJMXsqo+7OZZ+gvynD43AGygGQ9CwfJzXR0y0uswLMEZvJz+kpKU+P
snTHKrDrXwCrPL2/wQjY/+krvG51fZ7HU1HqaftBATo5RI9WRapdJFELfWhkt9h+kO08oZVHxA3D
iQ9pDb63ep2cCiicou8EGAwX9u8S5iBr1k03YQxTrf2IvBc3GKBKIma/Wpb+Qaii+rYJanYtEupJ
FVx3RoXfqkciNRqNbtaAtudEHXjSahyn3bQlMlbn0mjZ/OIlw0LUwKR9yUGtVuvGEdwa9xdeD1C0
lKGeFne3rB1yMCo8T2qjwrSzv1O1WayatJZ9td3o7pioSHn26f9DylVBK/8cadNx9DMRo/l20ZE1
/PitdXVPiXlNMqTqZChXKBYoC+YFMALSLAnNlk5/Gl5W8H9PKtPonmLz/6wCPr4wOqDz1kC5pLrE
02QUvwkUeMgHOyf8ilAb8PlE5ez+w+8t82sm2w4zUnqNQniqMz7icb92b3NgYK4JNhO/jHfpqd4W
7EGlWvdEPpPIoIvarRJ5GvrFX2lRaM4LYW3IFv/3CDcG8Mfguw5kTtMXZ00cTn+RgpVmeCBNZPx2
WJgvPt2kyZNKtEOrA5Y+0qahH34aiqVQhrLyEybWxgqyI9at4PJDjaAcv+ODcYhZliyHnuDqu65K
SL7upqj5bPzmREeftSpBpnIs3oKlXYcd0GATcLPaBP0s+CqHTwvCrhFb/y2TL/G3xdhnPaNjr/RP
B+HZSughnElUlgb7HMqdQTWNr3JIttDE93hvd29gNzsBYmiNqdXC1VYdipQOlYl3gLTsGukOMtWs
o5/aGXHpi8xjxAMEuKF++cA3VQkR4fulUHZqGEqhvPHtvGugLiuY5QXthcdI+kChvWcdC0wKnnzl
m5Gir56ZmzKxltArIQB00jfj6zga9s0XCpzJ3Xs68XMezto9Bh3OEpU0pQO6wMJ/Z3pWYoVGZ+CP
5i/agKqMHnCi4sW2MrGo37BQ9bsfTFlG2DcbzpmaqTXctn8e039JjaSahDE0FWJlkQ5505tOQLYg
itxiouTWSLpcdmFRKuZFXqyap+WnB57kyYKXDgbM4Qyr/NLTL91+O2J1D0TktWMw7k6oFmejpCJh
qzmbWs4Iw6Y8IHJovJjqHmWyrrNRCkRjLXajbL/IMeKMp3V8pUdzMt0dP4xK5VvfoGJiUvXIckyQ
9+zr4rzM4qjBXspINC6rBeOix1IC7jaeI/UT2Dax6Je3t3r6jO6XaME4H3R9SXKlEoNfxB0P06sn
x1cxV7Bgb2vFcxh3L+VippThIT9KnQEBNw6TcwAbMKzHgR4fLQ3t1WY6Uq0oDo3nBPixDMBhxwRD
BjWbExhECwIiHk5LlwSWedJYKuiRhfIf8O1YzN/K3Xd3ur6ok9J5LyESDVg45XQ0W0QiVF6Afuef
Ck0H0qfDrBQq1B6iL32cpQjpieCuo+670caPzhJ5vkYzeQszAp7fYW5YZutXG/R81VeU2feC8iov
J359aEs4ePZkrUml8mrNrZUUQbjSh/Ud8IFxYreJGjc0O/P15WmXv/X6qG6KbM2okR/2C9kupQr+
NLUapBdIbtg6RWDmVnJwQbJMYtK9FMmWZgyqAx9AGNQmU4gYcmlm44Hx040M/WTOtu/97idlUvxU
AlstG1cau52ss8SZE5V1yIzfDqYw/edquoMLI8xn+FnIas4h7PjHOi1JT1p7g2jLN2d31dFUMR/R
A55VJQ8uvUCZ0viWnGcQ5gZ83nYEbA9oLRenNP2Uqww51ujQCAPIdKn/h/DEtASJICnTqmhE5sJr
/wsWpS3JgIDz7a+xLOLovFLYJrOa00Vq+64AZdrbyMJO9+USAMBvxrQgLMjwsYArBLNUwF2pgbPF
O367caADY0bcmiG0eH2irAKXj//N3TSLSdbfnBdw8xXJQZOy18TgJ55LW/LYs+ZKLVvlbR7FX77n
BzKrYocrfRF7gkBwYjQh7hHdrBt37GnRCMZxZxV1ldAxFTbsjodwgb8HyNmSpzatTPb/x6xlXCZ0
rrX706LNCQF9ch2YjkkySOrvN5b0w5Eej6N7ghRmFF7hw7ARu41gQ/k41TM3FI8EtdggGt5yEePQ
127Av3pSuMZvqVR66YPW9lA7KL+8rqLeFlkDkWoxUd6/4hJ5+8lsK2bsIfdO/+F41Vs9vD/mx4iS
g5DFCPnSvZkXgSCOH4eLbKY4jiDFQXpvKb8YSoJ10lkp8QLm38f61k/XdSCsS4MH+Ur3PYoFssWS
X5BVGsAdsJIN2OoVS+fV+a3DcfEbvXp8+bhfxx663ZOOKe1T2UwB1VNKWdkJHZlrxRieuMtL431s
rIxcVtCMGjuiOp6ujyLehsGInwGx2jQ+k16P5CevRoxzPw5fjHQLYI0lij8D768gwc+Lh3z1GdtN
B8yfnQgTfEqYUukr2Declplrkq6IRUGF9NPQ678L3Sm4Sq9gMZ5Xog4xFpiU6IBWu/e7w2VxylkP
RICnCZr24IjN9AAm8fwCtyP/KdZe3Ky5HcUJNJTD3z9pXhrZoxcMBoJ6gmOzV/R7kZMPBubQSry3
5T93+eHVL1gApf6AplZVaJDt2O68AH6sPGwUZPaf4LAZLusjQeExwCGJAdlW6yG28dbQ966yh4Yv
49d478dHw4zMuiAZa6SEqUCZUXHafoEh27B2lOdlWQXutBbVslck8ZOY7/TM4EUnUgFO0ZgJoTKm
3/EUvOCCSJ9EshWvUpmnyEM++4U9fbn/tA6kjVLQXqygSzLk1EbO7CF+c1JxW88G+7zSM8QZiRNQ
znwtiaVL0NsWKUCdPf9pk6cFEQx1znGzTCqW4T/jldUxcP5JAdr8NjkorUxypirwmDt2/6jfXA0a
VAdmN4jeJuhOW718TgMmexdG6bUX1WSFlxKkv8MDhCVT3gWpWPB2+qwDlXaEpE66EfpISf+TP7IU
aq1GMoNVA007XGb5FJd/iW9X8Ec4fd2+TKWvqEeh3yEvPUhpEjHHemmTRISpRVBk6IxLFXqCaaad
ENJzwI1pSG/eeZHyH6GY+R2xDj0SKRo4P8kABreA0HIUhqEN1cUuN13KXiVOKFXLdtoD755ZIxZj
qTED/5JlUbOqHkXS+Kpt7Q5OkLl96Xj22yoZN/TtebeOfQlaCv9O6izqdepS83jzpp6PQtKR52Zv
VBpu3UUs8+gb7eByvCsUAKjL0WEnloywNzDMonretCAzjEkGdUoJNyTFtZN8I5ViCzbOOO5wchn0
InBVq2h8VzLI1qFNAkU+KemTu0AbH5zwdAGJS5PuNGV/LLKYbGXp12xyGXHmWOKa67Paq6C1ds0X
/sgIE0r0m7dbeSNDQqzSOppKqzXg2E4y50FhI5A3INmO2BR7S5G7Sltnwxy7KIkFN9dUS6Lunrtx
hTL4P9m+WEQSnPG+9SH5yFxxP9pC5ryIMk86KaCdAa15HoC9ERIL7TIjsyq/3/F6wnjcVrnrq9ud
xDna8Gyy9PynL7h57MAd+od1koRqkg1P50xSVWfnxIex0pLIESZAQzgiaw0b8+CApONtEn7pqUC2
5vYoJKBEUQnNt37UDxgMtJgIoYflomM6drDh++2+wE9m+blkxaOKkO4nPFnrWn7dDj73sKrSZ/By
5ldKY2FfVBgG97pO7t9zyjiHsS4d2t7qCFNegR8I9o/Vb30C0KLp9lFHmYn7ErMxji1rtHBmzBD5
amHmVAoLRr1wpqBdnX73Lb9dvxdyhOWiiviyZ4O14cD2pMITVFl0PP0Wk/HWhLEgy+/Jz7pZKrhF
b9AzPP2IxJvF7cluRa3KqoMfqhetqiKv7ULVM5zirbrYXQIvWUGdpHaV3lwQGpWdGeXDTDhFjuq6
sdifsFN/S5VVju51bXBfSvbIt3TEsw+Xt+QxCx4h5VMHjVXZ+ICB4VQpfZWpI6Z4FurZiV7NMiEy
X0X6HLYpGzlzH7xePa27S5pilk90oo5D8kUK1Tlw28tLMJtqgD4YSsAUDZuZyYKxVRIu6URZMhNT
pGRTE7W52T+6N7X8Fu3JPFyAFOy7CB2GMaPROm0pcPazzwq1q5zndza5wk8tw+5fGFUq2NTcABQZ
UU+LP//LvBRHX5fNdJeNurOnXTThbNaI70qt0CBrRQQZbABM55GjKRThZ14+LPmAzL7k+CkO5fyX
8M2pX01yE3UM3cWDP7vt94BqhIHN9dtbd5J/B6Fml4A5KfzI30q27CpZFjumICFzNFI+MB1iaNah
vVALmlD2P9RpWl2JAznHOsFrDFUsWEg9SZEjL6b6UBTiy+EUKvAFZPnIzqc09KVhBzTMuiRNW89O
m6U+k5Sf75y1OfC8WcEYnhVdUBenmUfAQR9CU/Ne4NkVcR7fKbtlyiIrntFKOClk+uv0ijKmxvIr
frbModhP2dSN2PkiBHu5mkvJAHxO6keT/XrIdV1PBCbo7rS5Uw+EHhuzlTWDu4yQ8ZT1uWOseQq8
brb0v12gtJSKjepHZIVlEU7CZ4Vu7KiwyZtiz2z8Q986iCItaUWUF6QPgra0RnA8HPqXhMRX7DjT
mSVdigRtkBfevQsBYf2zo8wz2T53QmFclWJK1baqkwdUygPmBPTPcI8L44bwcHqCAFL0YbsHE1S4
neQiRsIV88Q0UNBgglZMePrczEurXtvBoEXqMn78rnL1NYOGAByLVcQgt1R8rcJQhH2guYo/nBT1
/lrIiLsV9Rd5ICub4Sdo8Owvf0QELT/7qsLiZpykenghmJk41sTVMw9I+8+uLGrh7YQdzZl2bFvf
yyZaDyzdCXlZlgXiIXPhbxXFP/3ovq9Ioc5Khf0XgbMDqgBx+nS+a+PqgbW9iSpSqd+Xfmv8YlWq
pDpq+IKofNSgDOld+5Wto93E1vI3XfgbKRGlRM5GXZYUQ8OBMSln0Wm7b7gJWKnrAeIgNb4ZiglU
ubGjfNnJJE7QURsGIWrQaqzVjRSTRAF7PfeAe3nvH8w6kMOYOqQMoKx7ufi49S/W1TuDU19nQyMG
vavJFNxF6HndjukmFg/EyosgBoAcg9Z7mLrc0HNVdx8Eyu5tEijYV2XVw0L1vBGeh/qRFds35ew/
WxJkVTLWIfnyht8pwgHKIfYC6zs87Hl1blR+f2dqpJkjxKpEZXJHMOk4mL1L8dyvOALKWHtxRqr5
GBv1MPlWcNoqXo4MutymG0JmYNzehrnfKlWsX4dKBMnbPNp2OZ6VxMTX1VIRjWVtZHXk+Ef3Qz+j
ZnZh2b92BlRIprIWiXQxZg2sjJIy8i7bgPfREiowH/sbqESufUbadjhKB3s75BVmjv6HsjslYOXt
X8RW1W2BllS9w7fSIGigZRKx9XVsiIc0fyk3V8qdrj3iV96P88lKn+52gS4lamutpat0S/q/NciF
MJz6e4zlkBG4UBLRIbs4sBMV++YGE+Dg/n5lvKl/FKtjpvry6FTjv6UAwXRskrb8jAe/xxGMENcJ
PG8iHvwup/5OwCTxgxkXgUWHNvSyWZd55cu5yNv8ckIbcipJ9GP56T/mYSfT7tzAMUFxm8dIx1n0
JotEEghGY/zmZ9k69PyqFVoy7pCcfYEjOKV/Om1e5jhzGH/ce+igSKa2VCq+r1+FXh27fOaDuCll
ai5mXXE9DqWg99beLv2oOY6aQPYwha4t+MOKG3F9ZY49+eMo7DKDr/0fwzdPhMqU/cXFTlcaVPho
+gknLnbXX7386HpmTCvn9PhYxZlvxgkFeIF+dirptswjU1RMHwPeii/49hQbA2S/YWdGxQOnwoPw
3UmFH6DOMAgy27bWvVY/si4L2Aaj3Jaa2T9h0DUJxU6cTc/P5P2zIbr0ni3dYvxpdtQNVBeKv/1q
2qBl76sBV1Epx5AsJRxR0jdgwNcQZPrwmj+JmC6KrLm/hYGx5eH843vGvbgqD49SejNf/5dhEYif
iDvP0oXZvGIggodeb56ZK5fhgTRGTCsmPhZxbHqCkcrra1idCMNB68gUMSTd+1foS2MfOksVIPaB
AQibShgtJ5xswrWkZ26Yh2wJI95mQlNdac7fcj1ZOEnCVsYxvg0Wj2v4B0vxWs5twZjrTBzZ+ZRj
cOIPbJoGNYalakuzYYuOZ3OrtdUIz2q9Oor4vkG5z3fEb6Nr0poiwPm0QGt+A8CA/nERoCVm54P4
0ydTajwJiSzn4Gy1Yx08Y9v8I7qMmzxMXwa1hkMWIJme9AsbFv1pyA0tGMEOfWAnPAAUPyL/s0VQ
hVVNVmdp5vg4ob6T36+CEJRFoyCD+MeH6EMp3hlbmGLwlYxGBqkTMlWgiV1IIOc1LGpVIKNg3cWd
ZD//VItvEmI3hw4lKG3dS995S4mN4XfH6qj/1Hi1r+1DkHqiaTLQTes7+Gg9dGMVCvCg8PPagKkg
rF/TrQqUvCCLhRoIry0GnakIV5lAy7fxVhmPcvZCYRZYE4WOWeP6aFHg8Uy5Aslxhtfd/LmMazIp
fw301Qw75Fi/2VCWFit0F08Ht2y2/IKpc4G9nvykgon9hGkEl+ivwFQOTGvVoNvbGThal3TuYLHO
rmuzlVpStX03tq+l+ghujvG1lIhbVlrd1nkCegz3S7Q8lDvGgba9w5jUXYanHSCum/I4uc9ixFen
KuvXN7azFDZ/6y6aG1jE8sc18NOxF4cS5vPq7H9NAx5zDtxk1PvwojPUnsEqOp0K1x1uNzVir8YP
jgIComl0d67xOh0YET+NqDiNyEbeZaORXL/0JpE4viGzRc2TsV5oYEGH84ZvfCMCXRAMCTxDGTLm
JDk9XvyHa98T12fMkzy33U+lEZ3vEgOmnBRe5Bzybt6JFIGX3SeCU8eZLZpwPTPxMLrU8VwVe8Vq
8+VG7t9z0QG37tLn0Yhrmbf6jwDt+YEPVWWWPGkE7hJt+2F4rglnF/XEcXcRIICgioo8/oUnCXLB
CNFWTSjbwULDfP8ZabRRWMqmrAKIKeL6ryHBBYdHWrGocSRuwMv8FrlBhT8Q9t0Yv9dx6MMzXmL6
KJao4z8aR4O5twuo71W/iM0pzd9kPRETkBdcImXg5rij8AE1WnVDKf32QEXfVjp6kHaRnzQ4AbpK
YxiemL+eSGY7VqN8GrlQWuLsH21Z48GVoriws9DZEHPOGLvM3WWjMTQfio8qN99MyFU5OnTJByaY
OEsMGITltFYTYlEBt8lk4njc3PpLbiEddZvDbfSEzuQJppp/+cIUYFx0/Lq2xflvY52eFLcgsWrC
+g9Jg6y8tkqBUxEfhEmi2rtayEMaDvuMVtcLULjLou+AopaSgPI/BiFIrGXaeJLEDmDfdgCimEf5
MJI06qUP3ijVz9D24VteA8qS6XqSZ7cSzVlPWnCwReGlhGHQ/cn2OzNc2VbT1Lhs27rfD59Z9lQz
3yjxU5bpyxg6Ct2W2ZqN/sy0gG+2yPlw0jDRywOiuTRKk6WGgspc+eMuDoX451005Ki+uUrzWTMP
D/do3akzTzelIe6XRRYwvXShsY+5jmwcDrTLV2S7D/aadHgNokWWak7yZizfA+QisvmjG/e0GyOo
jLnJHRXjbWLwB3xo4tFOnSbbCV6ZmJf7cJ+yHjypTRARijX1cejeQj1IANzdJ8UsagttTEPKnt9L
R9Xcm6yhsOet+lvKxQ0TViwYFMUJNeZCb2HVw8MkQTHQihJWSXzcw0Dygsvz7KR5ZTxlMVCfpwot
dkt8M4H1OwuHoI8lHZ3wtdbVfHHPosOx3dQudHQoTTMA080/v0fgilkj/sRKxLnrx+oXyje5ggim
lEjiTF2JXQhTeF1fV4N1G3XDAQxKvFLSdL4wugz0RK7EcYIiECOl+TkMkyc58wmPNXlba/sBxFlj
jEvUuyxD8E0Eug8qL2HR5hth+VjtHAzm2Btg1D77NyrFR2wtRbNnFuk+k+jb8I/RFSVGlFREJ4/5
VuFisT9cukIJK883EB/XIrhTXvNqZBqASJO1M8eAPs5RfRgNlEXqDuMVtX2vJgqukdrPcmfITSrB
w5On2bGnnsJfqTres9nlnRwkTTGCHXtC/sQcCD8vPCs0Pq2dGx30fcpH2vTg7eeDciEEjC/Ka0d+
/33cAM4qeAeF7z5+Ik4exRJzjbyRlAjStzpclzDimPDFhA/5u/3XWIUhL6sQrq0VvYsdKyeWHn3A
8M9kOB5aliGiDnQjXgGAWU0dYjxgku+1biTnbJdMbnsJxyJdlYF9mvM+6CjoX71FiH8EVC+z58Tj
rorwMRpOi3O0BjRfLXkG3p73OG1tkknPvXPSVp1VmZoqrkek8QlhjhJnyBBzDAIJRj/cFiiHFvwm
4z4rdRRFbOFfae4Usj2sGu8AFay6odaVvxqv66AhKT0c0g8nCB1h6HFJF3jcfqRsCXuBOi+ctT6d
M7URXf1eML3QP6+VcV0ypk9GGQUkpqWuPT7uao/CfJRAudYGazmiYX41ZegTuHjqENJ3axrrBnh0
JF3np5w2ib87DKQHZs9BVRPH3shEb8KXThQz+iDVORjL7BpuyyeKvHTFrspkR4HUGwkql0si8h1S
GnAmzDZZG5TxXLxIm0axno2dnkjZ7ok9H8OG3SnPe8V8l4hX0/taVGnXS4uQ4KE+NH3n12/la6Ot
6Y7VIe1mkJcg4MQTo4J7CvMOX6JmmXUoIPKzo4BNoXF2mH3iZfZ5mRc+pyIJELY/kRMKsevoDxrE
vFzGcBVD8wlFykkh7UO0L0uBvVT4d3lqtyla+g8y4BUuVGVjGmwrdDjgzvVMEg/P+WhGT6DQxJj5
QPCI0Q41JGwJCcr9MSu3z7N5bW0IyyYl71btk0jIywp1cRAsnzImWZhBprX+lbI7hisyni8wa8rv
mwixCU9Cd1irf3yRQYUFSCxd2K74I40ko1qOslvP6Go+3B/+ZIXaqcNa8+J+RMzhjxO/koZ1j92v
SgUclC65wIffKHR1lEets+dicrBSpEaCfDaBoWqwrdocx0yOg07EPEFoL5oamFQoVO0jP42/j6ux
LObUs5oxrdcnl7UonyFhXNb06PczH272Npa7s8sBkf8qSb44G5ujxWx56GEu4n/dV8ygaEf4wnmU
RAyQSeFkvNF/aGaAnJZ1C4yt8Lfx7KIRAeEBb0dMEZYxAFBgC7YvQJXn0frqPUgRXvaNnfvkLAGC
WuouCKgmxde+2nlbRr/m7VPemK8Vy3+FFEQJ/HHnFVQfnNb0aIsIvKTBE/BSDI2yKhXrk5Q+FCMX
fyvsWCFY4wxClFcaV3sneDW5+7a67JE3zZng9NPYLqHERsvsX827kEOja6cdWSyFeudT5czUZApS
my8rG1iPeR/FdcqYAb/VYVvZblgq126ROG8cFU5CWLva1nKuYb3QgWXWuF66O5MfDH6mm5k6lbiM
kCh5fRNeYEL/u1BYcFQcHlJIWiYjPp7mbtyyjegVXVXe0ALFihqIfyVGnbI5o0Bb4Q57WhJXGGUa
UVbhwgobzoxqGOQmRO4XnysIc1tX39QSPq5puwbW/q4LkX4LCn+2NcdKapKtLxbdXu8Edgpyuvez
Izr8daOMkHkKwW/0D1LXmOEUnCdxVKLzaRcs5NNq/eCNTKPvFfmExMes4B3uC9xUHom6W1nqFwep
7KiTuPQ+jIkMiXGDxOJwKpfZ7taFUod9ISB/HqDiC4vfTmOfArD5lOUJX7ikidOyxGgYa3xepaBi
eY62zcJz6XJYLhfl2VexWVCYxkxYr7d0AhbnUKiL8/Qx89gu+BH+U5d3k7ch6x0ZZAR0ElXSx6zW
hf028fZ5SJpwdyx7SRrk5585QtBPqVN/AOTXtfgr3uvdzKjC2K7MDQQN0RPWdYLerQNsoO6c+ha0
Iim0eVe7xHSZ98FwkekPXSRxQ7GNcIl/fRG5NxJChibCt+kYjzreqEFbU6KTTK6eD7jII9Fd5dGk
0aSKWPyggqs2bmZ3nSTC3EeI6obbrKuKzauD/zAB/hkor7wG28rBxhJ5+j8SBNiF4fJcS3KW01KC
fvN61vqOi8thsdCz8cPKTCY8pyR4xojLc23nddIJoxOP0Ivxt07GZ9yhaC/95VqlaslK/c/XV/QC
ZU1FujCayZO9KTjdhz0kGeJA2nE9KPzN5VVLuR0mgo7BH83t0QjAbDLBzZpxqtdrXOr6s07xa/4G
s217Zht3v2d6G+/2gs6pdDR0vHjDxd+kylhaoVVH8y/758f+6dMG/1b357xpfvMu+m3GtfY6Yf+b
+Iwpl8EsAaOl0qEk+fzhHvRg4lrJDdwyqZx1fm/+fowKWlP4Ku+DFTonkMRmjshTMZ+i5HqHsai9
BqtvePoB01s8X8evNGJ8+Ec4d6996v3ZQXQ6ZI/NLiM0wecOdUfGI1pHrAAIDiKy5hQat3mwufGq
B64WOv17vZBm/r6lPZEyA8pIitA6ghrqTWhttqfVP+jkbr2OXr24uGkO6GRQd/aiRWCSOlofcdFO
UaJ8FC3yKkIe5oLdMPxBL93/aO60hJmFlgKxxuOhylmeMkb29nqi2QKsb59c2XON2G6rVqvgY0iW
zoBRFrfSYUyDxSJN7Tn48g81IT0pPKIB67NymQEyC/3swXGkuYELogFCiX4N693DFU1jB6Qc2OSR
t+MOnLFOBoBsE93wesAsrGWOzqvNglMa0ysfcRUY8q97kpr6FL9stDpI1QuS1fBDmPV7tHyKG5NJ
ZFyVsoOqZwEl5Hp2+/Dy/xkXGTU5o0h9ZSr1wihlXwun3Rp28ogZIssskRE410oFj3H7hFtiB3VD
Cp0OzjAtBqt2HnuymReycdRUlrN1de8+hXi4C4fjGwOlAt0dNiJXT4hX3xX8CR+gzx5RVlbYjubu
N3pi9FEyOXMnD84gBLuJz45jGPhRYb7HwZBmEkvcqitvHdZR8TuJjqj0Ut6QyXUawWihQ5Swt4/x
qbVYFRZdWX/vxC1tsxQYyBlgfsYdbbt/PEqP05H+fJeF2EemSc5A1t4Tdem/vzUm9N8Yg2W9UleI
dqFqmEO+tzZ9m2SmMJcDqowxfLNY5ZsbAhVhxqSTWSmgpmRVGWDKh/CLAzXu9i64+vAvAGOU11Ks
ncn5Qm20TVoksSFIZAcL4gBexNAlZrcP8f9vvPmc5x9Z3czNABhIzSkM3Q+k6I7VinbvQ1KXk0sD
cPrUbu49KooZbt6EeAH65mjVVuvCtkBlxKtDpRILqxM0uZNxvM2ZCqJE/m5XwT5D8p8cexoJFjfA
9ZklU3ZS3jf4SGd056nuT0KLFxT1pWUm7FRi5704II5YDPOeOoiXUI6itcKpLJTtoJh5shQvhSE6
pNiCDcusGDQ+E/umARVKIIEbviUaazSjGY3+BXZbiJllEKsawP0oixs43gVvFOafCbVTghgaLZlJ
ixQFm15s4jFlcRwKrigZx/aynAOmTOYjuKC/NrPgmlWLoH2dxD5TwZRHevweur9xKj765UDtOKyk
MNgXq5QjeMnIKukOCaEV2XIN6SWKhHHsEeejEYQU6CggiUkpaigCZM3zNwaAS/Q7jRr9OKBEu2DU
1Y8kmRFWoFvQ4fCfU+tn+chWQx/CPlonRpBOeixhr/1WsI3Afyfkwhurv83FgS6pP/qLQkMBqLXf
NOf6HldGVoKqX9zrLXShj+SbJbd1z9dYBcAMUz3btm5Dnb7NjWdBAxMq2dCc/p21caUVrx7T6Ztc
d4Nd9usQ1bCEUXkI9nZXxeiMSdR3R8AVrm+V2ZgJlXjYsg406RAW9OWH3z0HjC8s1i5W/7Wre6Ux
t+wxfhiHR/Ed20dexvvdwLmVeZRTdHZWvlJN899AaOxK7tSwZgp5jeQcGyDzsYO78h3A3EeVg8rP
+CqvwSJG/NDT3oYbeJVFtuY2KngEWwpvO2lhG8IPDsczbhJ56mkC4fhVnmPOrWx8hm6AnLghTW9b
3O0MBJi1ggIU6NZKTqXOg6QNJ8ZbJzkuLdet6Bd41fV1ueQmGbYRabLxaZcsqLZshgtq90h2MdyW
rA47Byc0w0i//Nwxos/Yvi7FOtZH/6+OfD+Jkh0GouzqxdWDjQhDKg1FrUGlW4ajIcPp7cXbkUrM
uD6raE60QhRikDlFzkBMPezUe1UvSz3IPLPFRDRL4ndg8BsaaMKXKcsK5A/LoTjTWtxPqx5ovHUy
f9mx6Vc5/rO6EAPI4AhFPwlzOLlrM77uFSfpTjCPedGD3MRGqiHOz1zildkQAnanIvPAoehndGbP
dx+bQWM6WYbXUXn5mgSh+jnU4AeYCN/JYyOVxuHCGfHewD5NlvARaC3y81K/0nC1nUkhJ1Z4Sv4K
uHx17ZfoZQF+GMgAyxbB+im4HIybz0PeiUswqi1sMLw1/NId7jrh8kvfR2Y/tnIHsIkddCSfJuL2
aKhHvbRrbxR5dVcL9O1/cvnWn73vszULToI5nuC9tE7/Crbe4KuFIUg10plduvi1O0VCT9XCet4w
VRVSoR/EURn/O1qXkhYuBcEWxHZeqo0xELQUmgCnaKueb/Vu3dInXtMjE7r7a26KFZBEr+h5rvZD
X3OOWtLzMxPtzB8u1HYTon5VdRalMU0AZjZXkWHD1lZaKZ0wOCr60zOOvxVYPZOM+YD25HMxCjeL
xnOx2B0L/Ya5H69AUyuKRU/lsn9LiqA+5hF2f9e/jOIWnzs+nOQaDsbHFa/RtLdHUiU2MUaAE1t8
k8gBFR8VYV/ihCv2Jm+25wHibn7CXMdmxDGuCOx4I/Y6f7PkU+sVHK/Wb+boo1AWQcBo8Fc+CYz7
pqZFN9B3VZVmY1TYY6/8JdM2PJWGzkY28qx2KkZ/r1oE6HXfRB7ZJojvwkWcNcjJyF0RaXo7kZDf
PDx+9sui2WH14fNOLRV8xM7ROngWfhbkOYElZj4jBG9j5FKBE9alfqDhzswnDwrUlZzxkTNDdIjL
WxjkCQXqAjXwuZ9+7P8/T08bDagrwykdiyOY7y/ZQL55jBL+ya8XaPsGgJWZFsCEn4sQclgS2lm3
uuun6S14Bw+mwhcigMv/BleWwyBXr3kuns+JcBFzSA1IZ2NDX93YfJZF023OxFBPJQBYZH5vO3AK
M+NCvoGFB9I8a0CTHCKANQ7a/8ey3reA1eRnvCWx859rA4oFHVLrKvlmvQaADVNYuj8lQBs15t6U
37n8CuTBT/IHnqtuURqMwkg8/ileO2uUGA3yf1BxgH9uT/MwcYklrpwfF+t+kOJNy4bS6i2K5otk
R2wbjNTDnZCUONbTO+NBD9nAW2th43Bpzz/n+LIWK9uUDTLggz4L4PZpL8s50KVeexF424fP8S5o
eoYKt3XNZfdHpxwB4g07AsiYCIM0qvD6xWlgYIRlwJN9zJsXgeID1pr0EcIcwWgGaP4aE+Gx1Xxq
xKZuEWVL8uH8gnX4DneWMKkTPlMbcC3Hb9iu/riKn3UBheYjcudd5u+a7ocj643FGVsE20hbXisr
50dv58NOYymNga8C3HX4oiZVx2EOJyrBb8Y2uKeL5LfzEKHUEUhTFlsz49qR1PBc2iYxzSMz1P4m
hkCQBHtXyJ3o/bzQCKLMPo7Ii8V+YyuJhQnr1X7X//BVWTqypOFTB2SQPrhbUm8asFaecOzUN/CV
PY8gyxWTgpLiZV7KsEaDBJdqPxsp3+Zk2yUK9TvooNSxwXOBN72wZZ91Dr5dEcTxwTpKXOjRjgTt
AbHrGcp/8EbwwaM0UYBAbYH8lEFFNiOL6qNRufIu7qvjYzJXTkvxEYJJB85Ux6dcyIz7LwFlrlam
9xFs+vcKsT3OLgb0XpzmaEa0nznE/7aKVf6Gg/PDNkshzQ9CzPO4EzKxmORpud6+SH/DPERgtRJR
PJ5MlxCD+h3pH/RfV2qdcH+ZL7xEVKbV9xUORl50JM0MEB+9ilWn4eOBLXeKE4/9gNzMd1O/2K/I
QOFFREkQKkjpb59kvgWxLCB+14dlJ1CgnJOMYOJPcp48Skmvr62aaO3HUJmLcGitWZmXO/KGhNyL
1Wdvh98rXpGu1AA6Msup2ZNdVIMzGHXG1OdikPW49rU+FR6SasVbZZd42rIgW+TYjdFBRMKPjRK2
BHgudC3EfZ3xmBXcEchcWHPuDu9MNbRT7SBO0gUTR8dzz32K308r97fvRTUkpw33MMLFai9IWwYI
2kMVKnhZkg/gRR9g5KwOkENxATd6SNRHM54BnG7zRRM9Dp2ED6oyIx8otIiRf8S8xB4/lAW7/avF
dHkzKNhkdu1DiDs/q51ILAnKP+y39XqVNFjpk9XbNKKG+Auv56CFW9lOmyDc5kTILVdY9887XQQO
WNpT9j5EidgT2acNu1HgO15VPiErFOc5wL1uS2lkozIqef/mYdLeDDEcEdNdN6YCKlMiVG+uhpJc
i9wmj2WBZ5VO77YhGYOq8+Hvdhb3eIetZRiC0rMvXq6zgJQdiT4M4ym2xjCeTZlVwkiBk6rMhGYM
Fw9/arC6Vk7ybDyBfuAeliMR1xIh7SwAmMaLPRG+tRnPAqs+Rl1/1xl5iAKqgxOqzvXAJH/hzkid
r+ZJhMqrBGxB5iqRWjnq5HIqYd++kcfWETrPkniQXVeiQIDYMjMXVnp2EUnd8nBUjpmwLcL0fbKC
U4w5S4PzWuUlFLyyIqj7xngHakqVoCKCvUbGFKE7g7xWljMGY9jlsOtUOZ8xt+lqwjDUrxDTeAtV
mx+ovoFoECBhI8f8vBUMW0+m2oWEcERRV0cKYk2ZogqYh5l2t70PXW0zpNca27dexpQKIROygOxL
4oE+/7AhqbyXn13xhSoU+8kgvWFlIWcJgIwBmaPp8tIBK5BdxF2gU7rb3uu2xS8rAaoAy7cYv42H
sVVzFfEXlMGWbgdC6sSlXiqgEUtU/h0Z/xHx1YRHqB0BdgPUFybOtvmC2YPrN5Lg2oFGGztW7rog
rsqceAFH6sNO8DDV5dAm/vdCsDyA+GLTGU4kJfb03Amt7yW9vZPO7dzPrnujjqTZf4pqcFsapaIX
/00MBzFM8yRAwPB0Se2qyWdVUnJ2XRk++oxmIiQ+2xmiqXSIt2pfn6svLE2jQbh1eH0QST7fMrXD
2JDdcljal8ko4vdGM0KhLHLh9n+uT1Rzq13Scfw5DFj7gmtEP+br7RPxJprhM4T5wjpggbozrw/G
eQ4hcJbgyeZkFbhPM0txV3+FDEZyyyfLIq70+uqMdMwvmdfRzleFidYm2/FeBsgqXjVVHPbXzt4h
YRcPVHdzQ9VDnb5Ts3vLoEk37Ve8bK4Y1obSD9+kY3QlQC2cZdRq3BYJhDFyv9ogkA/JRUV5I9nS
+FSuoj+gTiNIQHJPZg3L1L2FwCfercK37C51GNSP1Xma07nInbU13v42ymP9PAj4r5iGlvBxDJ0P
G0pc45vPbTqH4QCR13drv1oCskRJ8TYSVUjGpsoe5f4Gn5OR148QeQqlHAzMtQxO1XDHJSop8ziY
G1ab1Jf98rB3yqYg55H8xaZ5JIpR2J9+jLeFPd7pkqkXW/PVUnxbdQs+6Cr+bQi1fry5MSK6e9Yj
rwPMqudTuie2eohvlzcA4weR4t56UUUxmr/4CuVsAJYP1nVczZibwR7JRcn+lTfWt6eIunkvR/Lx
ckDxXFOMqwRi9vS8w0Mi8hSpdIcih8gG/HTEDTOYtQ4GGxU+ZvOnEQGHGJ6wV/juwhRhrPeIp9yw
1pxj2zBfKpF2xu4YaPdZa7xPUMJIGmhHI3h3bF/78SFh0IMpIo9T+Q72VB09hRCGtLzrqmzS+lpb
l1B6CQRoMGNBi1ZcD2As5jAxv1dzMhxzQNleDbT7BINxQGpidSiMTOVDafIVnp9AuL2DACATrtz6
9HKtePRRMslUy+8Db3vXLYFnWcuCdyQNoeUuzkKly050HZ8BBhSDPz/LnRH6UBjQ/z8rpdp8XNeZ
j13m8wyZ1OWwTEhh/BE9G4wxAIMQ4vszEjBmfs7uYRUOY5h7HJ700+TTJ5j1d0Byx9e1V3rU+Ujh
Q+yA5hGGgOZHPKPjXecm+nUOpQvT55P6d5/rcw/ulDTDVtOlI1Nl9BuLWlDuftfPQb2EnuNNAUnA
2AeTghwEB7MHSDZ6GPVJZr3HNLZ/k2S91V35oQa9Sid+Wf4/auxviA+HXxOKtdItsaP/TKM6/UhS
c7b0QVJbb1QaEkdmkohpPeDgELBEdZm5JbkK2jnlEikzI5u7atdkuRTVee2gVGs/GPXxyVIjnCBb
OqOn1vA10gLjjd2VvJHeSWz6wcbqo624sISQuTesuPvVu/is2E+OxlDg9DpgIKQyW/CiirBe/kCZ
s3Pb22gBV2qlqNzB/fNe81+XtgqRl9hb6Tqze7Mew2GQWKINHpp/ISUs4SnkIRdTZ2vCAxF6pGCG
xlPBWbD/SvPTRYUkMAhYV7wBCAGXws8l/QIKDbGSAWa4W+EC9P4GKl9C3JYRSY4TLzj+Ij2e8uI9
0h7fzbeEJyblhKWe3VdVXjkFlTlXdomdnyNTXYTeG2UHuKvfFoRpkAmwJFVutCY5wA810GYbqhmj
MYHVgeviZqcVisSxZj/tOj2DthSfKyPy86XWtx5U7z3ssi9GJts+jpqdH5uAN4SyPxK7YCIhmlR6
0GqTwqUN5MBxBb7sOMvWdZYUR7K7xqge3GL43DwyPA/23FhxfjG+3DRX8xMzrWybd5W7k6WIeI8O
N+EIc1FsSoggbmjwWD9n3JRpRf8FR5dzHDCGlYb/q4uvcKdR6AdYBkYW0Jrbto3Z2EFrCLasVkVo
cCzAxWMZ5xVHPXQrZQzwLoqa6hwa7WlibnKGGrB3v/7oWPdkcQIqmDHUV434nvV7UcXR+R9Jkx1T
rx8voF3BUHn7QGiW7uNmw0QlbV60+PrbLTls8GZ/3nd/VrP7HABIK7+SCgv/duSqD+6VNH8Ja1r/
8JSt3Fp533cH9fce3+FF8hv1DpgrSzlq2hHiUE1ufwSePnBpG0pp+YPH5lJuOGQdL3Oxr0FoelUF
upYPhGHFpCXs5Dhimo6cW661TgmotG9BVr6OoVX2zWXhVGo182SW5wumlYTPCPt7J892KeaqoW14
Z/ycxJ6nohxFB2MinuVTtptCw2HZ2rF76SkrWIUuUIIwRtH4Jt2mBOiszxxyVhFdkXw2oQW9stBT
bnGAp5Gqg7exIBYK+/CUSX8wUN8V9/B5Hxcx5QJOMLuVeYImsqF/5SbRUwfthTMVRpYwCRpowl++
PaymPxzV3yLU8YlNjl469DZqc2asf9kY5xlKxvOGtdcTypU7yoGQA1ShosZo/WGgxe9EHyPPOM8I
UCvhzQmmUQkv/0VzZZR7kKNpNQ3jwgrVtn7m+8vANFIuJdcqnf7iHZf42mMY1UABrgzbjYc1iCEv
xiJCPbTtuiPFZbTmUHK7Bh6Skqg9tyJmkF+VSF5C6yaEmGyCWI4b1c1qQHiuDoFk4ug60ajCSH/M
JVt/NkwgaIzFaXFL9LFjsNB9ejqUokpEwoaFqYJzbdKqeA16e5s/OevxKPJlzRuPuNbHE0aY2Hrx
cD1hQG/jOoguhhqAZKKRqVXKMPHkqSqwBkTndaSvBKoWzd4vRlwp57xBCdkBz4aMEw2kx3ck5gu1
fYWIdZUmA9ofCn+cGkJPmoaXM4DFinqS3ntpN5HHmyh7mM/68TEmR54if39i4DB7j/8All7Mfw/e
jVkB3NKmWmsmCxZRmtBzLg4QQx9z+/5Bgq2KfKgtee4135D5hSvfgiwEqq+0MCxBtk063RL4upcG
r2X5QWWdoHkQa0anuaE8UUJKEARJi+nclQFHB9/AP1JGt1TXx84NeC+Xo4ZCoT1D4e7KxEyKDD4A
CKkMhmOYISJbh+H4a42TN4qxJB0VDw2e9Cj8SZYGZ2HnTMhZaT36d1lhzJQGsbs1JDdQcOeI5mmh
d3GqZIJjbWWabViOylgXjMxDDaETJHDNlHK4wmbhOPTr/noWcba1L66liV1qmvYUEDxGBDkPPInn
ng7+H1i+JDRn1SX1hTw34bvyN770EKo/A1Wl278zjMsT+/V0xn3cO3I3MR1/Z++ydnu+LUz6SsJo
ykfuAyic38DZt6+ByLqwiHHSdPYT2sF44YjkJZ6CS+/mKTAY5JLMlIJ1aOXKc63uBVB21DkcB/Pl
5tug92aShL/x6BStPwQBwbzptq0P4Lbxe5zUADaGHefpFY/Ftjd3SHyEllknUOUEqUGvv26CtzBR
zJ5N9e5O2bih5DXzn+1TnjuyFH6bq21NjNE0Kqun3KQnkLYfiRlNURYuq9Ok+v48R3fC4P/5PJbe
oY7KhwgD4EBSFZDAUJoOy/hPKthsSmWaGk69xltj9o1TgzGZfAVJ0bmlDyxwC0UswVC2/gNJIZvB
3MhVx3xno/yZKt02hDI0x5nsNDwFI7L4hsRyCKGOqTY8G1aENywni7qa7/izxyhsKHcuCWnqXZto
BUq311NK0B8bKuxpQOxSAgk/bmVMCcZ3qYWWCT6JM5hyIaRQ8Tmn0XN8MhddSXHjxPgkUWFo0Krj
MNBUaVXENrl9Q4P/YztJNp9K13HlShGlCU9d6y0cHlunTpF0IpgiGRV6nxigCpk8bTQMnTsM76Z3
qibDNxBoKrpiJm/nEd816osMAdnSN22PYC1DU4YMdMnYs/LUFtipXvrr3D2/22eVStbitB2W6/7Q
cfYh8TaWZVndxSzxB3cggTmd2I+Ihs4sGEXNm10Re1GLc+CjYPP2Go2iTI4j1Y+tacE3WYXt6z7J
vYIU2ou1qQMW1aA1tdcSMmeKZn/XzEtxHM1TGLgN6b0q2yIhNCzRjvaAAoBAbA9kBJVwb6vdXANG
/ijIbwSHQnNS3UK3CUjTJeG08O9OPYNZSITnU4yh8e9OIGxwkyx9oi//hKewUi2WHSu4C5fmzVGb
91kN/70H7g9AOCC6DpdW0mKkAupfRkIkhBuEmY64vL+0dOcXbNcUw8dX2waGVD6j8AhMq14nD276
2kj63zCFBJMXkv7YbUX++5WukQMmIGicqF1zCOYSli7Udd9+1pFwilVCzQF7JDa6hd8W5kjeoSN3
U8AHyBAms1pEglWgwnwgnHRuaNAstXRSDtHvcwhamf3eXV/DwUYEIRVHJC5eYOa0WVYLMiz2p9cF
bYNnEz12Y9KyslYrBHf0PRu+JAeZhVxZLL0V+EAo6M/tiBPkr/OKPU3Y8sa9rSXClB0mwm4efP0w
yLSlRUSVowpwIrTUqjSq1CIbamQ0cyvSc4Jrbt50GB2UnQdsWJvA5FK5D4Ii3ikJ/7KJFOnAL8Tc
LPrVXBUAT1Muq3j6jNgOC1wti0iiCndhXggQT+f9L3bBwev8PwZri3YcjeGdw/ucS39b8Tn6ly3N
GI7gtuNAL+DK/n5BhDHeC6VksUB1TLmsekn8AD1VE9l8kzr8XAcuWsWI58vJEdMDn3Dmp5WeiryG
bT6zgaoiRpfm5gSXmMxa6Mo7rhipagc8v9WMga781dmJrAKiocIZlDxvlcFNUn1vmjtHpwkhvkzp
deqqdKTKe8l98vlkLCBhe8h464RmzJY8So68oQ5WC4BWdzVXB4eW0u+b8MgrP/a1BhLbzcAfHo3c
Is4U433HVP4m8Jpc5nghUwYgnSBPrnFO5rAHNN80NRHsdqmsfaVWc7Nw5EvNjxqu5Q98C8vba0Jl
T8OSBeDAv7hYRkS6N2uvcvVoBqWDm0OkIJd71YH5zHyP5Pgnc7FBaa9Z0M7icWoninknhnti7Iku
u518bvY7vUo4KOxSIgRLY5VVhAJnCYWtzRiqlY2L2U+NALYN8ElZFxT3jNRqjTm9jMMuvMO6fU6o
08nrsYwE0gvoCfVp72z4n3g/S52Si19iFHk5E5ZsPHggkuX2Y7gGJSh/alrJyaii6VG78hTyKmIx
l+cUImFhQu+jCXUNOjtsmbHI4YvkvK/8AuordDHrIqmcI1XAwU2lvQkaWhLaeHzUW9tul0h0It4a
YTpAItdETcrXbLnjO3VnJ8K53v233Akobaj1spPAKRYlCKYFCGwN2jV0gtJyEGqZydf2bSZB1RKV
Q6tCBvKdsIsVu9qOgfxK601TUHUg8SU+QkVwEo3MT3tdkrhzco6btFHTR/VtX6ZMW7FeQBdzoe3r
GD4mdrX/tOE307Dc0w4S03O1IPAsAF4UCeXv4XNp3vbhZC8drJOEXrvNDNBGgOyYIV0qysiaY6eS
WUSqd5XvgCx028DsrdPLzKWcre00y1tITE3UmUhEkVv+3PF8LA0KjeVbDlO26LxgXbAL2KCXJRLA
GkLdzxWn8OYbX4Iu5xie3eZocXqs7wCp2EEo6Dmd9wqRErzBdI+gZn2Q5DxQK+fedy0PwUHTTQV9
X5dKye9T51AQwLhms1HcKj2UW9TdWPNwFSfEa+DCa3BSWO3mg82InOobJ4AJkfjkTFd/5FzeL7nX
7qN2ngeW4QzarDr0A2z/aroF3V73byAMBe0TCOU0p6a/67qRB7HsjkVVX77Yw45dzTFzERk3W6lC
mF3xCGMudFiCD5hM1x1aqZBuwYjF54dyspF8Y5VaXrAp+fiGewm7z4pBhMqtSTTb2fEjTSTUAXCb
MsrvePcTL1uB8t5UXIwrMzIH9QjwBMQ+OmG5HHjpq/MqlluDpOMuIlcBarZiqkBhzuOh6f6ev4qT
nfUYeqfDQkvMU1b0cYG3ySiiNGf/SOZTfInG3YRegYUG2eTgzXradE1SF3iow+CARZ+y+pYX6MUU
yfdL9gj+ur06zuz1cHu+jwZUeTX25sy3C/5i0LPeGAWBMaVrAp26YiIi6S70awuERbxJKMk5ThjR
9E9vRWvhQsyCHqIwuii4OXfIQp5+jVls3XO4LVlI5ow6oymmZG2lXXBPfxD7WhQgRYKfz6i7/xnz
9lY2LkhyF2rirGIgwgTkweJbxKKYYqsykXyCwPx2CB/rYbACnZ85FQpKmYMqo87ulLB16LCWzhVI
+kRxiqjCXk9C1QLN0cujResOy+iW581kmMMTC1bJKjCobRJSmFTjE+GzJ2ndjIVDoqF12Ozq4itN
rZ+0ySHIQEa6pC8ByiTZuBQMooi5HT9oLddsidJtf/WTA9gxMBBNEvg4Jw8K8p++0w42+hhE/oxf
PptDrM69miS/QI3CXkH8v0yMGudTeIwTYCBm52OpqXLmb8AEigoAP6Tu+eMtzYhO92hqLQBXhksW
HcLvbZtmZZMsro62UynEDzlQQOUnJ9ErWKi7mtUV7NwKTwetSqomLTJbkBk7OX9R6fy8TBqA3oks
E5R5eVuKoSWA5YvnR0CuLX0waAWEMsh9DD84VDPqvBg/u8kAZawn6bJsWsn1/cJhm5Gw6NFjJUkP
wGWWu5IPWH3fUgE9D3lIISoEWDcNhgCpJvPY1DzMrh5rP9JCYpKKNRtE8vf2U0NVK2Kj/a7sVBr3
0pV/UVLZ/MHjtceB7GtpK8PeOv11ggC3nOApiWddOZlpNoESv/qEt+FO9BZpN3fMUssrgM5Kun5A
WHhzSKMsu+2rJEvaOU/LCbqWJK7lI+hqdn7q0YU1S546kRdGVZFNKQ1ugQ75woBfRX7/cLG7DDlr
kYQJPOLPlbDkYqrA1My6q/m6wlp4kNKWEfx2tGIPXUzJ5wystbJih4rEIoDRRWvBoYkiFeo/Pe1Q
PDQIEDoQRUFbiHGt4NNEOz/cGHr73r2NCvsh3bSvUXgXQgn5A72/NOHETmugar7AJcEoteAl768o
5En5KTH9/OPnQdxrFlN8T+RjPnNuCdZk7g9LNnUoEPXGVwZVBd66ccoVC5HZsChiiP7i4sfmwRQe
nXdljY9y/yHEwUSk51OuyKioWDVcgpcN/7twZOZDZqRZvTFar/xfwuodoEH4t7JKWh3bESkb0As4
0Hk+i+zYxz4fa3VYH2+dtfjOxGgfvSlJBJF7DMMxGKOEl8p7CBZ5Lj9VJj04/1l8q4I969p7qZTX
msR3EmHMiIGSaGOgJjWesnJ5eopCyM4WmDF7HFJ9+ARRYwyQGalgQMdVvt0c/Z9TLk6ani6BXKOC
fLNq8YafF/RPpvHaNm87Omn8BXxg5Sfe7cRDczZH5U15vzm4KxuZUyfZejpXD75ZsvacFEtR73yV
TrE/fjJeG3/uz/UMA859R1GgeW3I1QZSIo1Z7g3min/LJircQMwCzzqN+QWuYHeJnA/iCWEDYhiU
dUWEmBGexn6Bqu0vXNETvMl/GovkXdQL/jWEFBuLcyuTyxjP5inee+uWF8G/YnTONmURCOQWF7vF
FRJqKn/Vio/EBO+srNpm3FWFKSqEplULKsYmLHrzVaQ/wHCw6OjSLGrfR+Q+HhZNUrWADnOIgo79
6NgLaTpB8LZFMb4K8HW+nR6AbXFxCHYrQF/wjrmt9u9xDmUPS6jZV66i3pdRicrjaPieEL3dCOxj
jJBqRf/FVzbtifwIUjiX7l5JBBdwK7Vh6/Ld6IyoDHblgQDRIuexh6Mine4FV3EyHdvphnlwpLKF
mhGLn65SFSsAo8XTW+09uEX0BrAoC5aj2bwyFVIVgjXg+95MnJh0qv8QGaOa2rU1jN3plkk215Re
hXEVqN+CB7wxcL6ereaSxVi7PZPPj6E/l6iHZC/7gh386xqbNSdne+U54RSRKd1WBsa7ldqhBQYe
L79o4OtYyqX5votSJ58/UleuyLkaK1fxwmabv+TpRNa0TtUyTt2WutzYgl6ToQ6PGSfIpqw7vIxI
HqVkAHHx23L9/SMFF8RswUpp18IBD5Xaakk0PbaW34QvQ8NxPQEnLnk9/tN+zS6R5rfnD0XB8U8M
8af8t+Tw9UPHAaLn4twWZGOcbMpbw7MM94jWEXNwVHt8sI7q8X/903qrUEm935rB91S5i4zMTLUk
M3xqhLJ60N95brVCtjldwRJeh+LNz8a3uSLRRnsZqpizLaA2NMB4A0c9SpxVHJRmZ1ERZ9fIn2Gb
p97xkDKEn2yGVMDU8kAE9zvButXAKxKSydLEQAEF7lgvRpoc6zMs23TESGUZYsrlpVdbL5dutxvB
G67wA8SrjuU2r/12XW05mmw9e6i8ONshzUX+RlMLAjvNaAuzVgf8st6Bimgf5XAGwxMSddknxOdY
K8ljNFlzss6jgpeUfzZpY3vZFzLKuCa9nyN9NdDO8RqRm6rIyQOhXDgAHiqYkCHCiUXkFnTFzm+d
qFHEPCpqAzisydVnP3duBWsO0JU9qMiaYJmViUCv1GJsTB6rNQLjoZukJqDfYRWjKscPmI8HGC57
7NbyRZWtUxKGcSVkQinUM7NVKDBQehJDZJ5NRlWknTkLGAV/LubcPek+tUkyTWBIfYwPQk8OdPBA
1BXDAjriGTwgS+W/V/Xbww829iVlKxPTRnQ1PvikRKANGDC8gDLtUBwq3UUdSWTG/OJ5Zdge3+7P
1/+Q82pk2Zrs178a+jUqGx2YIc1N/Kx5+jQ3Ww3hQyzCn3exBBJUAKDCz7cquzO/dwZYb7clNtzk
wU8SKLwURF2FhKHSsTyMdv5R5ytnjLcVHPicSsC1vO+cIpRrodh+uh3DiHz3BsSeML+n41R4q5I1
mZ0EEjuX2TGvlcAABumAHb3HibKjD+GjBhFM0BpXw8GOAM0OR076r9eZ5yuCnUqQB3zIYXFGyogx
odv2urHMOlakDVqDNmvri1v9bpkaYI/Yl/ijjhtN70Bh37+J9PBo0pRgkAEBPiuLxyhfwimaTF5S
u6Olc2jS151JcbNf3a41nveVYEZ0QqEeSeClOhRQPaZdHmgzY/k5ZF/7VWIsoaEShStbiJ8X2l8K
OTtCdLWwRAia7wRljONyC6+pKpM36O245NhSLAd3S2H5NWYyOWkTUiz6gcomFVlpa35brVXQeTwC
C3arrsFQfX3J6c06nmNi904wR4IMVFQBdy8DbFiJ9iK7Cj9l3DlSasHS+dMYWVe5EozluYmJ5MTK
ooalwTyllfBQG7RgZXWVO+feLre9PJreAsSxx3okpLoIycUJ11d9H1fiHISHw3BQ2UWvXQdvpE6n
PN+rc0en4YHOnEu5i4UtqttZJ7fghDoWxzCBLpUUWb/Kdo6lQ8CDnuYIqkzR7Q/nSAMi0B+5aPdW
l2e7UZwLirDCTMm1ClPAPy++fvxpGwqbyP7GNaOjm3m62PrxeFCi8nHXmksOiuoS2NN7bb1gz6lc
Uro8WZUJp8VnrjSQNJYzCGMkxRrRyCFwBYJxhuRe4ZUdd2u+zSh4mMPcTma4b2gwDaZGP7GzWZTw
6CUXOAcfgVMPz16N7hfxVDw4m8uoHW+hXvRsIbx1JDAqKZXqc0WHTkeeZf4+RuAGK0sT/eJJdaeg
iDkNdWWST4kkS+PDJ3VRy8HKRRmRVG+2SuZ5R7JKE1amqeeJf2epdqXBa9u/aTz5TAn9ZSqdDiII
V/dQF0eVo02s6JFrjxCkbifcMZSH5ly1lt5nA7WUMBpP6yyh/s9xQE5LYb4MXq1TJD+5J4ekyATO
8a2/tTYTdo2iBq8+3Tlarv/gON0r46qZCpiwVZVGGQuWpeOzd/xINGATRSRgyv/Zithbx0hGLv9K
g1Li7X1RXx0eQdPIW/5BacOtk3nfKxVe7ywj9iJqze7kegLh6LxsDRk+mIugKjb98bPXY1Iw4F5G
Puc+sDWWEfeRQ06fKTKx3Ub2W5liqcIlrSNrgL5suBL1knjdzde5T9t2YhPRIioj8+a75k8SOrUA
WNqOHphnptCA5nHbEodYttFB+VpJK7RFgDiQANd/5SBvpCqDhxo2h4rK19iFT8xY3+AONHlpWMnt
RvYIz9tgc9te/m3oYTxVi5S7SFYZNHMjgDOWA3zuvjEBCG8W2bObGAlvEirP8I6y0wSZiIPTKTRI
Gci7X3XM11iqYbsFDq2qivY/h4J1xCHeIZF3ss9S503BETgRkLA8jNrcb1B6etTX5urCT2n6uM7s
zHj05GbPfVbxe8ufUSkz/cyfPUkjK3THfipG7Z7UkWc4Uvb8D3z0MsfR9+ep56kiszoCmDgGlavo
1nzxOJKpqncmWL7G117QPzNPBnfwLYsqhmDtLrDlOMzRNj1Hk7VBnHAmgt4eyBjMX7deL9+zx3z8
vtu1HpOy2v6IBlzuPwomwxiq8QvtfHHJFmTSn4iH1jxNXOaFzoXAEnTVtnG0BUxWrmTGP1eYgM1R
xcV+YJHivPYewsu20C6zliXRx9ntoVdLZX1zgaGq8Bj0GYzehYuZgOZpM3ZHDZDdcQHpQ2OZBXgS
KZw0FOeccp/eU5ngt3iQJUekt3l3/Z54UiFAL10ZPT7YM+gMkwulEFzMgZSllvEmiMbrJeUMOCgK
mSaS6PHZNIXi1CzG7myv9/YttKwc/DxcjvtRN4v7OI8ebXWF6VTQIpKH/uNa2Y4vhQLFbWffmIaB
C4Jt5n/YuwLl6WR1Zk2Jorj7u7mV5tQSW8V0UjGwXIohOrvwFItdBp+WgYfmusZbiR/nsCKb+Alx
2quz2V3yL1xbhYhlGv7SOaT6WjjsgpjIS/ApvVkPTSAlcp9zotG/A8ZGGfRtCrj4RPp/5xZzEhOt
DCvPYIQwBrfp4XM7KXqae5p7irMKc7+tohYPtK7uwUOONQzUstPPuKyJ5A2UZT1vLynfG2eayGN0
JLzoaZLkiXCtKRjXN7oNzgDq4piStbLoX+jIzppg7PoxpFhMQpP8Qj9bae+KSvwGgN3hmitP/Y8r
X8Xr38CUDibkZr2Ox7zHl13Rgpy6d81Rk3XEv6H92vUHFPQIaWHi+atUJPaRSU7Zy9r7zOxFSWa8
NdJr0Lxw32nmbsJl+x0OWfb94WQbhdnYugjP0cbUqkAitSwCiOBsjsTFCvf0V3Pn3oaIB8ZCA7Up
qQzCUVhop2zk5PAtOGg2/Z0nf1W9tIXG/6mG7rMoNELp4/Sn9c6VB7LHEBQBUQGkMA31varjYvvg
qrJQItN0C0bNdxR14EFAPzBg05DIQSfTT9A70ZzENZFiI51UE2LcYkFTg21XTPqMwun4XZ1CHGrJ
LSn5td6RDJrwMjekq6M0CVYE0N1HMSmIfmfl7b7FC0hrz8HPdHMJ4P7cfQzaS6yLNtRqLGOKwNKF
WyxtPJD7XRt4OaIyJ+ZANi57Lv+Qt4oUwyfVPztskaNH0BNbOPKMek5LPflcemy0POI3dRCD+fE3
wwRiub1x64qc2wN58h1Mq9smMWDVafTeI8E7zSQ+o1+FzORU1G/e3WoJAdaGYcaRd+/2Cz2xrnSp
rPheeB0+PAccKvMv79IWYy02aBlP+EX0du+cyLwOs1UpIoOwfYTbBDl+s8xoCnsDMtRKdlvZ4kl/
m/SmMZmPF4qVJNTYFdlDkEZ6bbGCEVyYoyHv7X6oGC4I9tRKr2EeMgrOjuq9i/sINyDEWXBi8IPG
uIbhMtMUy+6Xw/ZAxYqliZus3VAef+91J1jBe3q+c5jfnLu5zawUmCCrq0SyMVakpT8eTSGcpDA2
fqXBSm35dtAMY4JaJhsGI96qU5osdRTnSW3VNfCZwZ4P1ptPSdfi6/37vFJ9Px8pYIJdX3dUdV3O
U9sZD4EqNheZR3EMXDfeNbz5zjuH5Yzj/KD9h84DgqWQluu2A2k9M2Ww+MS3UQ+Udvi23tLFw1M0
vTRO5GcdxVo8O7uoXWHKOKlNBd+e+Ked+BK9OsDVf2mkPtvC+m47ebJ95zWsw1BVNok7Ll9U7Xh6
+r8PjTi4z4hP+U06cA1IPwqPImnM1L8fNGXtqyl/WbagpkQlqkHflUlGMpSfFfxASXt3JjgYiJHj
p0HnPHgfSBuqweU2WnwvUv0LRE//rTiHgk0ATdRNDrokTVAjaJ+ac8TlPkH3vYRuPi8wlp9nGW/Q
yi67T7iY6+favnQhXygcw+0IPdSejpdt1oXl51OovzsGcP2WGrg1myPWhHxV0+7BluW3j4cgNJkB
HWqSZdCDKpGXA/8zNsoXmiWgpbcsNEnQWZaU/xKWsfwDuqCnuSPFFbSB24qc8YmC5pkggzeh02nX
I7XYQhf/JRIqgpmiwKpatCbH/GxmbhqNgx32p2pGHHujcfZcYrgD05Kn33XYoWZiSEOm10VAo4GY
xa+pOkyZJLnQmf7DzxoViIDgQ80551QlLSGc3fmWzq5nrysW1vycAqqJ1xR3KAopXsKsU2SOE6fh
L02ZVbzz1Ov5tNTG/koQN7srEhdbBWeKW7iUPlHHlZPjyrDz5Cb/TX6X7NCGv00aaDL+wCQcqc3H
AH2xA/k4xxrVR54wZrHva63IBpVWxhUmVCGooeZrdO4aNeOwRgjDWyOgMT6FPzL8siMojlaT7JZg
uemuZx94TbeyxkmAYJ3SIDGoyDU7vCP+TfoGmX6qVRdHv6T/JnwesC2I6LYnhNcpEGMA7Vn/k0Oc
RDr8QaXWxkZUBNKrVnTO71Hcdmp9oSe+1dDxBsv7GWIwCjxwOvC0bna/EbFjayYv9qDWCgu91zt3
t24t0JAVqgs91RQUaN/BUQTsAyCl4ahfwlKU1UJD5wVP5izvRq+WxiVC/nr82sEujuxyqVYeHoRj
vijnDw2HAk48lIX+cuI1xzstms28kiLoceo/6ae5EZPuBF1xiNUE4kHkaa5OfiElETAh93xjli90
mxCR1c4vjf19gniNfAstjm0l5bu4nezCrnZ+V8xek4NgCSrDMvXTf5JfStU6pHvRikVz3D3A3ECN
0MovUXWW5S+vK4Ac/YoRqPaVixbj7SAQK5A7b2V3bvtLcJ3lhA9ow6IAIGxTSk+sUH3w1fRgM7I0
LUzkDS094cdp6vFnoD96eQKsLW8N9Nfdfd0mY6diUC3Mm5KAJHO3J5C9tXxoiI6MviBmspuuIPxP
HFRyeTc2rAY+PaopNWU2aaUN+xg4j96i5vLT2PeI95fREvVLd5nYzXNw3T0w1Xst5BxC+6PO2m8f
zgO+66ZszzlMnUROA7OtRxsbi0ZiqfPvYWq1mFdWYdxTQQmVOos/gJh+EpAgY0ijAdYUwhMZWOQh
pRXAq6MNRhfLZ/Q2xDsPPj4QwbhXs9/Ede5qIa85ULbeerG4zmJbktaUXVtGeqCXeC3ohxcVxytO
kKtR+8N9gMiPr/FRm44RrCc78GDNToIr2lB4haoSsfbi8I2Wtj4q+50O+Py5qg5U5Sc+bNCi0ZQ9
exiomicuQMw/gMmn1tRv7oIuU6d9/Yya1HIqS48zO52nltlpPl4Vw/TRrXsX0GGyk0aZwcfteGGp
8URmrFNUP6AHhffSIGPMZTjWwGAms8l6VZXrimhKD5FY4ecc5kUJMf8jaLPzekMuNeWlEJaOL/GX
xHLjqLr4ou+3Tyfx35QIedA9Ul3nHVyVUeulZxd3YQGplSMYUEmFLN8iTJ5FS0i0bZjRJB8nLhrI
hw16S8Nw5Z+Kd0xinVuk5pxB8o7CcQnpy49v9VlnFfBM4JGgNpZT7D1AeOu/dQSkGAFg5aufvoep
6WSyPBgEFR76Aa1dUVpY1WgsYnUFMO+y8IqGjqZKGYbYIRcPmcnzEKGVwqdNOADYQXv8XBBH9xuC
isTDhp2iKzAGt6yjNHZ78ZKxdeqzgNcr33BJe6tWKE3jrYxSK5vFpaHx//N5XIJboG4FjF50FuAT
Jq3lJEYkj/b/uJW4LfqSRyO6sQ9qsCcMV8AglOH1DOk/D4Ryh/Gsnr80HZmRBzZVJHXScXiFbiDF
s50SCfxKmbbHBx+zVjo/tniGSkdAr/Ok9JAiLypBnYkR67B8W8jt1E3Fn/z5To8s4K0iQzhVm02L
nN6LZWvawX3ZdTN2L8BA+wSpxk4mwYbNdkSxD/EgLsGpgFJTlYL8hf7xS4gC7oj+ZhPQgEVHesj4
hSMOfb3LjyDvzpOcnE1Yz1pxbtOwCxP9gGsB1MbVa5z3HW1/UALJk9bMdP84ivvyZwGyqalPLQBl
c0HJt10WRn7q0657cd8lEb3WqRJMybDyFMPtxndO4Cl59TkiqqCuCTB4synEPW0fXXHLaP4sC+zU
loxEKH4ZM8o/1HShYUTAKMlnDPS/vaL7+XTwRZyCtwsPBGSz/Ck9VzJEQtEh9eqZUqZdef5P0d+0
pA6zF5BoKNr8mccDmp7RWuUhBjorSIMhBGmZ4QYoT0nwVwTYPHWH5fuUmYb/UBHft8nT+oRNthgk
XLUyTkWpfRY7xUAflbe/Jd8pVaubn1gpfTWr8kbjl+k3W4oHlvTrHuzyRWtbJKZqSEZg7Jg8sG+5
ptrPkeKcrpA9FRLq2V6Wq6AvK9r/TdeooWGJfPGG+BaVorJX3ixL25p77p8e7AKhTRIyANODPqQU
b5I5UMVOjfdVV0KObGnA/1cmvBt4sE2Qc04dRPFnai97zU5PQqOpsG/fmSNwe5/z0sUziwEH0k9W
W3ACtRDxCcRa0Am+XmeCDgTw2nF0NSP54Mt5HeJyVqwV3XT2/FKobGKAtx7tITFJN0VAx7CxMrkC
4PcktkTHZl94XTXEFoUUmJhvyaaKkGEpOTWWExhsv+cuje+YsbN+T3JAREHpErK3IjTSZNUp+rWE
6mFzOS9oqwMkb7WLFU0QjrMtHu1tk9KSMHd6YF05yWvCzCIjNpx5kuIqr+buyJqrSIRvQtStxrZT
fb+PnGwmOT1cVTadGKkCi/g/g4zNt/AW6dP4Leci/dd2beODHMOl8amIvDKYwb83eTFMcZ1tJ4Yw
O3T8Z5JwAHR4f6bvAq3w0hMyLcOVRx+YnMGKOSvKruK5X5V3P2rQ9Mv2teSZlYCv+UrdnlrT86TM
4gAaVG01ah/54xyKOj0UEPtR5qbb1UyHuJLWg/CHz2sLQDdVAScbhaqwGOnml92wJf5QfjrC4LhW
j820GpZ1/EaXYvih0fol0u4BMvMj2kN3uGPWqK7lR+wzJMrhCmF4js6ENiP2nWqg3TVPR03LrRm8
nErENCDpheTuEDT+deb2+Tb/tMW/VfATZKPIMRf5H1FFSuiwZCL4yuW0Ifmo8nFzhsZLycw1wKY3
izyzGJht3b9/mCXCw+GUyYfZAi8NqxlzRwvr3BNWYeYqfUYTkUS0+qbdeIBXuTso2EmgTYSqza7w
kHKcOZ2khAZq1QLhsvD8MN7xHWy5DE7+u/MvNqiNsU1KGVTupxz2dSAZXw07bwihZovB94e8l0rR
s4ZONVUrlDW+047RDBPgPrdo7fci/ScpYw4JZJa5hYs4+GKLeA9nDZEYhPJbJ3diYWQbYmwNU4Ly
5CdmReWVUhuHTz3NArDQDEe2Rgr3vwlcRXAK92H6u4gycuvhb9N0TMaPSJJGoQFzP1uWS9zxCo32
zkN6jNbuj/Nzee8uROXoFNGQEcs0yzCsYvQVO7uz5ZA20zGmrdMu9HKsYMr+Pa3HHGmY/SrYvbi5
csZtx6CJ32kx6CVjUJ5H4KHbTKKeYP42eMHfqmZSUZIphKJrTdE3B24f+UUuw3jPJ25mRbu0yif0
U/GxrreW1s94g3Rs3nAFlUcaW4FekxRpFZPgv63YHv2k0G3SUe0aqQqXldEQcECc2mLiAM/xO0Sv
mUlOoI0zqpuORkbNtimNaKYfIC1+rmIFb4GT1fp5JQIQl4NPLklyLM4Uio051dtJJoFzA73KHX2G
KvEWrefUNncV3pvDSIqR5tmKTRky3Uv6hrkdJV7/94Z4lkxLJrxGKB1NHt07gU74zOCX7/FhOTQE
Fy/7urcRh4oN8YuRovI30RJLTOAe6sn443M9goqXpnvMqcLn74GZslmayn9OjsZpoGU3gFOnxh+o
tcilhGN7luPMwjjRzeb7paYqhA5sY2mNXNecMtSlZZZQ03EuohF70PMkbCNqnx7HxIVBMoJqJU0K
ZvBg31o9bzmSfhrhrSNheD6cbFmo2LAxoHi6QgmiXVpJfAXnceK+2eeSWUjreOw53gCOFcOZrHO5
wG8f+i2l8Ur3WWjxC0Kzw5E7nSBcZXBlhRD/tyLhg1LVi1eGP3YOUeKqrGDJkADicaEduJS+jMd/
u7y4K0qBr4gjYHD2ozLynaORt691DoDCn1FPnoXsm2pGeC5Zdj0pOdMLGPAHoWojacn1/ObDWkVy
vYt4lEWT6G9Gu5qCPVtKpmbBpe3/6YjRjmsjocYY1V+4vMik79h0A0qkz411jq6ht6zpLVihnFgf
kCTNET2HtMhU2ZhTE4kF9yyn5S4oCs/2IehLnx87h7AnCaCN9fG8RUXT/v/HdVcFBE7cJNe/nC9g
MYV+Nj+eWk0uD0i310jRehiU24yfQS0F0pEY+Z5rJ5Ed2AXXIPlg/381MGu0ecm0O+bacO+BBAbt
P7Qlj8bx6OEZcMlSEUXzeBfGby39Jx97tJCS008Y1eZQv1RJBFIwndnlhDWeyQ1QL6OntNToJM4G
BTST52ZYJNo7Vi9+lUu6ZEvGEnbMh8ZxVBuCUoxqbnO9r7tkjXL05KEfdM0CHtz5k5YZZ4ZrHkDh
ehRSCt29/i1CNoa1gjtxmIZ+dt9Os6icqZFEsvCJUJTQNgQVpyEXrIUPoVMEg3DEhKIbl3yhWPYe
OeFKVzT/jbQaFKV4EsSvpgLzy+Vh6r/R3pGCY+SUv1I1IGK00yUuSxYaxs0qk+SyK7oNJRp72oIJ
waF3DHajCVqSsC5kHMk2/svWskP2gRTBcXmgxLLBBbv8AWaNQKgxZCWEumwm5Z14tkgWazw/oQ+8
1gw1mbSFOtdX20sHJWuOWpHO5CT2L3V3RMH/tBXFJAC3EikH5E+r+64EkU4JStQfZ/zTBxM5bhXk
pTveVHJmUp8tupE/qo+1a8SSLcFmqsdljgpqEtl2W7kYG/JONz9rvVqHCkO1H3OQvDMyRfJ2KtHD
HZaueMMrKhWA390JcEgRrOqFq3QGusbXtbMUD77N+wqLnohw0plWswQLVge2PG2STd7ANuuy5m3z
F+6B9ZEUMqDjkXsBMhj+V7QB+WCJM0VWZsCckHAEvML1ZcD3TX3Fwr2JLjmdJ0w3NiICeU2eDi6J
wHm+K4C4CY+ZsTq6a5Rtd6SEdlyzZCOS9ph8Q3TFzs9/5uWKeDiLpSGWLAeOfHklg8dAOBG3mtyO
rZUnC/ijYoXuMQbQERIVOtAhJYnCov2O8lPk8fbWxY7rCNoKYKOsSpOUCNo8qXLfeRx4MIJx3XNU
xxrlf04hMB/zdv+1n4XMJu9592pIrJxb2n8FCY3TW15oICdq4paSxxJ2hq/CKJbgWbxTSzv4a4g6
gUYpj9Dcy4onvMc2uMAxMTYLJPMFRDjiTXgmP/WpsB6HEeYEHy5mwWXB2M9vGERR+zSkUlSQbsFe
D6DDJxWiDbxzc6G7UwM26SabwFI5SBZAo1/PsnF9smkj8zhSo0vlHlXldAmhLBMNEJEtM41Ew8vT
14UMp5/Rgc08Qsh3uyn1ORXIaVyc86cxgTWTnS91ckr8jMGJ2frhUZyLgMLRc21x8yVkc/VmVnsx
7g3Nfq4rm12L/Up7Dogf+hxWhWn1PFnGX+yUQ4dgr9bMaRMbbhm5Mq3fW/SeNKXYm9pP5I9WM4Y7
1vC2dwfIw5Y9eO4/6WFsUXMRq0NJUvn+O1JlFXnf24WAoLZlAr8umNmsTEgkbpNyO1zAG1fyc48o
nw5kK0eoN9Rou5BxsuimehHWAV9I32J5NhPDfwFgnfuKDgAHM8vMvy0Ua8g3dhV0SjUoQPdJech+
B+ejiU8QoJDQhrmfhDSJP6lrdtEKuEDKdbc7osZa2K3xKfLmA7prN1h34LidP5izKjW4Nr9jXrAS
r3+SHPRIzaHX1Ofsbl/qmpY+iHtkzYCbY6cSB5LoHFDVCBzE5eN/754WczPIPPGQpp8NVbykb53j
kvEgqyVXqjkgURrNrXWZD0x+Otxj70g6z0kU1GCuiKhvll1KtuxbWoQeSnlSRCwMGdfLql8rt/1x
ELlQSa44At+xZuu47EozSG6GcDrXDCQNbf1VBr93VDLHUwae1NXLDrwbqZ+nbsQ5oUUjAAPeglRi
l9oBFWqhVylrvjH9LnApiVpWKaqF3nRtRxYdFtZsiDNvRJA72fya/2maepxuXfqwge2938DsjBTV
n3Xj5as322cQD2r8njhEuXCpORKe9nhficWFEhSYTl79NvrtJuH7fKJpMiI2sSmPvPsxCBFt5xFQ
KgYwZvJIeyjPOARBw5PEMJBfh8ONSSidHMvh9MkJIVLBbE5hsdZagKWFFrOv0S6yyEjJdlwlnJWP
L803GRbH4/AiRu6MquawQRq0YILvQUa2yVAQLZKqnodsVoF0gAoI65ifRH9FLK+PMrQGGWomCqHi
IqhriWTjBmrcaQPflzEa0BIskSIUzSQCXsDHh6yW0E2TfPLpOdbAUnsHr1sAnnhN3ZUZUxWIGR/a
Mph+6zWwW3BIZdIOo6S7PPAYcmA1MpIhlikgHTyDBGraTAfgVVAWPJP3uAT6z+R9py1HSBNSOtoF
1GJIjvbHw/c8K5bTr92fyCymy96LHym4bkOHmLPu84NTrVfemioVWVEvGRfL4ZAwpZK6CfQvN5IB
IIMHGrXqHZ76jCunahsrlaoelp1o2dGSLY9NF609Yw7JZTljmTh3MpMg4rEF6DQUJCjzU4/wXpen
Fpamp4ffJFYORwpPohcaqcIrUsd+BhVBpXlIfDYANs4yFyxwz6Ahq4k8+ExbqEiFrz2zQihBB5Ll
O4Fqy969WzjHQdvSJfW4hXo4ZXZm76hp6p16gBdpZIXpqxMqGpjjTyuMEKd/4ZO6LMXDDuZ16oyI
q1Uyl+Ly0oRWEOIsgjTq/cT9vEoqVGJi7a2ICk9YjvnQsmkX7MZuNje6gRmmqed9++hcVg3ojdTW
0eJlMlQPgQHAo7hcJNSZehe0djon7oAd9vl68wjkGXGKBOqRfpmoQV106dSlt2qtTbFet3ONYjvH
bhnzQcVRe7h6Lfco/2WkJgxMZjaL9eeRqgTA/6ug6BbDv/VWUxxubs8PNJnWMVDkVSAauyUWkHLG
clh2QQmATsrrzJWP0dbQa86vNH328cWs+uYESbNo8cx/sywUVlVwPJKp1A1qzdqn/4RssQLhOmWF
OwvckDimgzi/SeNUSBF3adoj7i+FSCR/Ceq7Iy6K5jdWjn0YSeUuldbDhSNt7Der1o0er8vn8wru
3bw/05FAOsbGe/1+uKXE6DD4WQb+uY++0NZ/fY8NAh0rzwjaK8O8cfDdE9+r1MuhQVRejBg6JI1g
b5VWhknQNPp7Rtp2NUm3pjlg0exoG7mOiuZP6a+tgr/rwl1xfgQbkyIGFztgztVshYjwiuc1Cp9K
0wfSmVKgSqtTtxvjdcZEXY45Kqm4rFHNcwZFD7Oyn5bz94Y4PMln1/EGm+ZxgY7KIWUfpNg/DXZI
OFWjCHp22VjsAnlU22uTWpjbCKS1U2NRoeZe+hDo6Ye0yc1EOiKA/8eSCjfxxnwgDQX/x3mwZsPW
t9IXynbzYmQAdlO5NprOqnnr/K1wb/luLCrMIRojA9wOL9piReFLAu67VDTpyCDImGfXXsvSb4UQ
V3AktRbj8rmnYxDhHpbzAZAp40V8kXhjOxM+DVZU6/chRiKsPYCVLoaUWdwXMlBdJ8WjzcsSTZ4a
mkPC6pZQr4QQJy0HLiSSyoLi5CIi3XOD/GBaL0kTzLaVlA3y+dNRezTfX65LtRMuKJSxJmUrTc8c
en6QOQgKypIMvd/UzfOKWs1uj3vrqqzL5+RVn29s/la4MICPqstfrxVjOKrHxa9Vm3RrjZ2ceyZC
h2TrRAezIUYELULlGJ1QWxHV6LWNOHKM0kzNt5WQUAGXAob5Ndu94p087X6HFl11B85xuc3u1Cn3
o6BRkHImt67dwt/lcNKBL+MtmUswaklmsy1M4Hm0DqesVAcxlu9XCg6PEaW6aAXcSR491HERMspG
6Siz39bm0MNzxCSMX0UONLeQsi7E0a57+hEwMmKvb/C4jAKIPcHnp+AFgIBgELkK0tTpJBqjHgDI
ufpjRRn9XDLgIABoJJf1iTo04NGLgKYvN/e7YAZoisnCIP/yfK1eMqpLxzmrpM3wNzHp/oViQADT
nb9odzw7jiJ9NfcNEaRszd5t0pbE6dviMDfM28nBgjvoN0kY94tph7XGtb7gH2oXgja2TkWKFEwC
Qi9Wj29xAs90skrwinLiF8pRiVnifknr7zhFVovh1UMIqy0fOzYk01nqRY225FjuzvJWfZWlEFUV
w0AsmBDAy2z46Oom9vGSMBa6VhPsjhV5gEiOhIYoRaTW9SlXlVCUnp5WlQ7tkyFiDJ5vC/BR+OVo
UhV/C9hkBMfRH0nXWr9H65nGiI/BPKAVOQh4xULVQth0Hd4kj6mQ3IZFA4n1ADcaLC+hZxwDPsTC
LMHeOFXRXX+wPb2tIBHraoCTDT8PAx+73rCBwtncAAZifOlZL0bxuyZ/Ea92zkSjybMcylb2xIHt
MzaQZj7JIas/fvH0959odGVa4Uro0gjEOAQo7t+uucMRh097TPpxCxiOMpxGUcD1V9KrojX/4c8U
71QPY4eiwmlUPIcJ6j/PXseiVmGekUOrE4WpUj+0rXPHdIVP3u8aMcxUIN//kd5ATUmvjptc7pXF
1nRk/m25ekRX8hW/lFkhyQ6Rk7MBy7LzpXRSz6WH05G14y6Ig2JLViscYGw6grUlCTRNYFLufDOJ
Ya7HffoSbsBSaH1uesfXzrFtaLjOliWDUiJH8MTiWprCCcwJoE3Gr2rVj0fQjhCvWCdwefTpDjSn
jg0/zaIQy9pt0Br+LzpcoBg5o4GHkhJVcUsL9SChEAXjRcSGi/94ETvBH20DuMYuwBJdDCKiA25a
jbt8IZBykinUz4j5IdZw4BAAKErSsz8zi7CKQ4x6Z/M/8sg1h8rYKziikmdBrV/mc7XmVMO3CfHf
rPs7q/xWDVuYzh06o7lAEJgDG1bprS+ZD86EfrzL4OgMPcrqQAJGVV1n16vWcf97JAgzTQDcgM7k
a4b4A2bbcrESGqyPZaoxuJ94UFQSKU+hyDGseU5SeWfdEvn0WfibChsSY7dbdN49IETv9lVj1vZ7
zvRjwQBo/cP2TWSQuolyJzaX47UCPQJDkDAPYSRKywsd/UyinM4R2n7V9jggkrxZ94aGt5oi9X/9
kO1MWiPUiFjbX3bSSssnFEFgVv7v4jJ/pnZu3w6pzx2CQsciqKAk282JsuE6ffVDiVOKT0wtkXAF
+DviuMJcCfColwt7RtET6qDScY5M7J3tQqmRKH8UIYfsPGQoRoqg2hvJCkRwCBNGE+grhtyIIFbO
fkveldsMWPekal6w7qAnMFm5jNd8e7RP82rrnuFMtSlSVclWdzUDgVBe02JaU+knuZaZXsO/LF/1
+JCenf5OWVayhlx9SxWYm+nVQSoDzlW67OTotpp0+yJ54v5cbjyAksRU/9/PC6FJDcnskt/CUPxN
UTzzr5LUs7O6Y+tWH/w7j27ilx+yvdpYJPAnTOEBMSBX1cMHweqdlYpU5d2g/npgzqq5/WSsl54d
rNBDKKjo9/GqmmVgROuGTW2z1LOyTB0BBGwqNGvv/nZS0E7eGjgRfc+16yWiHMnx4lSHVxUhgZkk
FlVJmbRV3AB/ycAhxA60o6mGFaaqDlbEHH9NRbWhFvZ0+je2oGR8Chx27Kg51Vjn/vheMDmUsL/v
773Dcm/5hZxWZk1sz1cTK46+Tp2n9UdOrVqrqBqQ8F7PHxRpoQIvynRsBJpmCgzlJ3D752PTwHEh
h+8qxMf5No4hv0RKlTMteoAMUcWl/jlw4gBs6PW6QgwkFdsQ2WmK2KwdYTKnVgbKa4k0xBQpom9p
x642Dr93IdvYStTzomD68EaaPhEYs+stvpyjsfHcjUyOQXcj5MPn+MBVSX+gILp5wfglUk4EQ5QA
UoDuxzL9RsAXru3LT6ugg//nln2vP9h+b+/sY9fwCOZZ3dLDPv0sAwL/mb4q3X0vXp27hIrQkmZF
9BmkXs47NyWBZC/6QniPG3csZSVsJ8HXL9QZSoqG+duU8G6qzN02mtXtAemKlnqHXtjl93wrnS2a
iBb2B9tTAYYoZNaaV0mOhgQXWM4d/XKMQWOTDg10YJkvFcUbrgWNNIrxMPiyZ7XG3XVEdPcYi8f7
Vrvrqeuwo18eLZT+O19aEwAKSOYdHJOGg2T5/YLIO2PtWjeNPTsgFGXDyzdZrAFSbinksQ7O2Hn1
aTI90bkpLeLOTmpodKBUaOVwVDOSiJl/rQpj1vB0zDpqc9z0o9VeIx8vFKX+nARQK0wMGmVTpeDY
RMzjufKrNPzD9R8lILUdBmClSB3lmMos1wQlmFFHHNVW4tw8Yccstc7otKErzqDVqh3A4fIEwfxm
acLNpMs2ay84Oadd0OlVQxHiUarEDFj/z5cLS+CLuhvJI/K8Hmps0QWbiddqAfITiX4+/m+R/6Jo
wwag3KS8zyL3wlLgdpcCSMojvTcpOEDKftLecDuGxq6qJKAArYYlp6XVG3bhC8Amo7NEQNMzEjxH
+7BebgKheywgNYvtORi4pRF2YJZPaUkAamMA/A4rRujpRum6z6Jc1I+2oDKrfNq0uRs0cFCuN8i3
Io5LCAmvDECNv6dHhqcWkpKdlkfC+0Qd4Qa4QMw0jcxOu1EkKB/y5i1xmnBdQXTPAgsj8MjvGMre
rNZDMuVPtesJbVG1UHEe88M0snIpy4HpIflizEMv66/h0IaEQYbpsSrA8msAvnbPJQDMZyKYs07F
AAAvp4RJY8GektjOtcAS8DV1KRl2z1xK4YQH+7vSjQiKgUsfqtV0tcm9PVRn/AivsxxHqbM4pJCd
ZmTmAclpb1HC/5jIaPHVi9DxMOl3b5EgtTHW0acMOwraJLf82X8v+c30Ga0UpFsQZCuVtzpFz9B3
nkFyQNa9iM7/WoahK5eqCdrJanNOQ3/P3W8QtK7ktGIaFhlYi2hNMMibYKUNg+iVCHm7aToJhUJC
9unvevhMe2o/COWp49sQsjUBK5UwIp8I3KuOHwd7viw4WkM8FNyMY/0Yj5/NItdBcT57B7sGM9C3
rARj6uoIJ+MdcTyW3kempskDA3giuBS1y+IogqmkeZxKXKCdaH6UI7X/ecgCcoSMJOdVdIUzplSV
Pgxfx5f+ra2GWgod1o/1wYdsVSavC/FVG+7QD65Nd6WRMLscxUfMBsGow+FwpWZlavOV3Ulig+CC
4YpcHs+sJsG+lANUff+CQCVVIdE5LwK6c+E+G9waHHiTxSkcZ2obdMzUxHCZthNcztIVsac/Fng/
jhgaoIzl6OoCzZb6N9G4Ag3ixZx76AfVbnq5EkgqicNZtTo0BsjpRmKqRy+NcAmRf02KOGiLza0w
i1KGwBXqPBfWTa+5ZtgUMsObOSk2GwrhWJUkd4T2tQDXPjMz9qp4QLWRNzrFrWZZxwgOqXah2m5H
7lbEw2v4EgdnlMkB70WlVJ6+PJ+tCKN8SvQ09TYYCDpW8KpJGQInM9hGHeaXsqXdS7PWHGtkYQlw
7hVGGduVinm25M+8d7ku9EX52EvpfC+bg17+dHH5MWkIxUKvrqz2LoOGLUDkjT4pubN1dsjcDQO1
DghKmRX+O3fJ7ZPY0J6LJouh3Cb4E0OxiJtfwTgQmQ22M0suxSZ5gxjg3zqFc0vSESGmcGDB233N
K19U5sfRsn0vcSk3f9/gttUob16mLAPLSxw/PxUypROiNhoTBQMgrJf3razkG6H2TUoFXS0xx6En
W8d7pYC9cyG9MnuH9+7Tuwt7Wh8ESCPTtRgZZb2EKUSnQU6RL1frDWiudW1sntRtDnuCSJRvJPMt
VAxVNCWndVrJWalo9qIXS5Kxsj+Ejo/7zKDeSjMIBmS85HVlQOnjSPUdxK2NI7VIZdM7xt7dWh+K
/p0VXPYMMlMh0ZPE5VUFsvm9M/B7CVFrEtyjKAbNOjTOqaEdXntNUNzATCSfqOL7HuxDh7A/4xEr
5PkJAVPGdCrHBd68h0gxR4BDVT08re8j8wmMUR5o+PAIZDkCZVHGhOG2oYNyvFZwFSv5e462qpNe
I0rJq8/ZjX4znTalD6/Yfy3MOcuYDBsR8cqI3Bru1I4y3BbPVSHLg4KNFrPSm8a3CBZKPCDIoDYF
lsZoiyMwYSC8F7DknlN448PXVbIYPIFpYJpPJt885++Rh1OZjFJoCyZ6WdWMnf5/4VZsH+Se9ICw
uesdwXYdBNYFrdhpc+4wEFya5pAp5YxS/vpS2mqg0NdeDRg4CQxz0Gp4Go52Z2akQ9ZXwRbWBRji
0CoJZv3n10K6CQDP6Xf984JNn39bMuzkv2uW1YBzW0q/zTOHHBtR0mHguNXU/WcntS/0m5KBOjLl
Ba0t3RUnjRMi7jk9daEYXr09S+UcZ+oCxnmWfWu6Td/Iz+dYoxWnHnW4Ep+8B7ac+uqHixbM1eMZ
830bJTEWRMZ2/2FwYfhWIVrYaVZFrDbN1gSaUYtmMiW+WgOqsi2peUp6izdgvSLiOqrkfuTBj1jW
kSc2xNR6V9reRbyLqWHhIpaOr6xvno5zJyeXQgu0IhWUl5O9ZOu53gBCyNgP0vaKhRt22cT/dWZz
Pek9tzepFrgriR8y1XFZsRvU785E1mdXknxFlmQeglJxyOy2aKS4AAHzvqx3lKvxrd2HaFAxS34K
AljJDfNOzswlafXNAyQfwi1Q/pmmMvOCdqGiajwanLvez+H8OZ6ICcnq5/BXPXlOGkVQ/zwGadJS
z/Y3B/CXoYBzzm7taGqadrVgvlQV4CTheISWdsVOIIKqvikqALff6xW7WKE7zUceqTPTfqjpNlyj
f5S7ZLPUa0+P28aukRMIklBdquK6ak1DvMym0bo/gkVW/vfE9wYk1WbOuiEZEuqMeP+IhfVYQOBu
mn1migBCUTPv9nCbVNvOaxN+/zSm4I2hiKB8Q4dIs8gMHLp8SfKmEVE86iVxU13XvmfDjlwRvoPF
zlvBi9UTpn3OXOIpmODLllX9zO3KdjUHiToSg25AnTyzcHcnG+lqMnsCztzlZDafwzOJB+W07ZZB
Spu0MUY1M2ZiIk4K/GW6hS0udB9tPdIbGek+quBKo4563mpfbGHaTB+fH5m02s/DS6HxqpDpqCmX
AJPCLcpnWmugf6UD/H3cOgtLDEtjiuZwRld1+/0Uu6J6Ef2OJsJ8rvWUxL+4yXSyXxnGvDzY1Do5
O+qnNmg04WYx7c+g7TdykBv3fvU0662Q/NaST6qA/Zk9TrzXpJKAlbgCcjQHLdW326O8BV9FT9cF
aQc/Assw+uxyNqGhkP2i2ZoS4yZwJLxW0M8CcgTwCpQSCfp6Ye6sXAz52ih3RUjB1noRtZVZmTjg
JQasbVUobeRG7l2BY2TVc/pXrrCPG/oZVWGB4AyT+YneayZQNphB7UZSNrQUOwfT46URvb7ARo1D
2o9IAn8FaJKvgMTxeukWZEIixBKMrWlqXX4/9R8DcdRZzThbAzP3kDaPPRCEfLbJKCUMiQThPSFX
t3HOJ6B/HjqEKtn1UlyZMUTlWW2Ud/UqPSllIN+EhhvChSVm2ue9A96tSxMRepJg3e2Wq5+YTafG
aqkJGCAUnQSP0VkKLCe67U+IQ/KvtK8MQX4cwhZyQu7N8OOQtpQwaTy6P335atPI200e9BLO8Ycz
OPrivjVOqUr/yooaHxZY65MTTBiPsVx9AuKwrRDltuvJeBYwVxMkK/UjOlMOUbkXh1N1QJvOYe1A
pcxyokfQeEEUWCnbtZTHwKwyiILCgzflCS+hdLAvfbb0tXhCOjOzl5HouncMJScj67iGSh1z4F7N
i9ZkVjZ6lXgOqGW4cn8gvDAIdkZP6S5i5cXXjtH4zrQDDTX60z1gbAQ3oYeUh5dz8TpHIj4YDXDJ
UsjnbiejwZyowMW+EgEu0WDVYpCIaJFb4pjAEqjIF8SnkutiDiNWPYXRijI14MF/BQQjhQNuif1Z
gxxpqs2OGU3f5JormUrN2aQAtErCG7o6XtkTf/KgALxVOLRQ2LQAXCA83+38M5hZlOB9P2n4SsbE
0LdxA3WXf/EVOfBGIVUc0Jmo3oENFuUfb/2l06UFj9MTlSAhIzF+Nd4zubXD8HYPs+pJ06tgyIid
Lmf1sK9iXLMu2P32RWcKP+ybp7MyhR7CgRBiFul9wUoCXLhsWnwBZggsUAsCUkM/9UxnXupVpaNm
7aQmwZOR0Mpj9PDo2ZffDdq3eYdP1FAemweBcYtYMwFEVbB/SvIWkp1lLhP4PcnqJTBU9+bJVRyy
I7QjHRG0OIgXRQwamhrn98+bYY98/jK4oIWQBJFvcTTP6kvMQKAucAP4ge0ZVajoSAcmF823ZCJQ
kGKSJSOTab4lx/VRJNbRXsq1Yp6bg/SR9XFT1mmh26ZBaqA9tmUwJnOehrH7CrJO7qmyg/pKrgIU
CJQfBMtG6bK1qrZ69MRexJddsWjS+rHz2toMvnJ2LjGITWQIRqi/+l8dfHNeQiYzwYkgs05rfuBP
EXv+GfwwuNfQe/XIPY00vitAAkK1+eY2lGMRbEpbinDt2H2fC58w1O0NWDreEzMnTEbqe/7FwUVc
WLosURs3mxiHrpBTFE06c7XbgFvv3LPQjGY6PLs/34lnmBWUOQbnOCTUFKL+gmmX8Xx+m/biVasa
L4julXCq15yFwfFFu1hV0gfGUPKAlyFYDw3IRVwM4SrN6n+cE2c1wM6MTKf/DlfZFCxcixRR61yW
jr+q4AH+UFG1u2vu/MB8avqmsaFOzw8R+6hxOs+fGluew4gdEQ56rhDp1tz99eON3vRB4bjkMMYT
bs3Gv3WkXhIrPjlN8lCg3DRbvD38JwJ5AjUNS83ENXVAwMTSvHS4kUhxlfxd48RI8cDiAXn2asZP
fzz+y5NpIio2nmrHXgT9yuVAz63EiKaKGZ854BoYyA4USR55ElOiaHtCTFtHPj5Hg67GBp0k/F4O
WFXa8depBDkcHWVq/yWG06obw0UAZBJN9FTkHTZ0JuCvvkWBP2dM4IYa4d8zEThq82Lscdh3xFeE
etA+8VH1nMp946LwDuav5mDjnXV/d+3WJpzjvf/Lz/d+c0VcxkXAPKjrKWyE1SkvqgU5AtlXM0CD
xlkjON4ZeWdofeIljJhKloUpbPGJ6T9zqB+eyyRSyEhi9rbcNs3n7Dsw/rMaT66veqeIruDrPF1u
CQwxcSl5qVds9WWYgNYMEqOddGVTSjtz7Tcr4d2FRa0xVSN4Qa1MEIBFHXIDBl2O9CgZpgdg0vjv
TV4o29Fqig1KQyHeS0AzZgHJMyyr0lJoAnM7EnxG58uMaEMC9cI6sfoaQN209XAPFAKU9CCgCJej
tfAerfvKi/4QsP2PX8w/e6ny2kKphr51fPaZFE7si5AULHYanniOKTc18VjrXlNZNhQbGdS2Y6Su
W74yACnJX4q46vxWDIybUws53ZOvGCoaD84au0dcp/LNKMylWgB3uKcm7No1IrZGnIAqWO8PIkcV
tCidzCYyA0lP2mH3ylv/IDtPJ6ca9g03q0noLP99Zsq78y6ApbfQm7W5Fuk9MiafLArVBzK6ycN3
813kNmUEfpKC7cHHaU7viMxgoZ4ZeBzVDfTH4CWPVVzIhIcJyEcgE7zgBe2Izzbvbrsjpb3IC3mj
hOV1lBw5NUOadMpr8pphvq8deaH59poNpYcbKzKhEaY+UMXswg6R6633TD82n5zfRlOBL1x1CGcW
jFioBQzvTAK6fp4jV15N/cW20x0lIgagmF9i9JdApp9A4HJgOcOeVLHVDzBwTx40MwXZlbQTNNOG
bpeK8yz+yOYzTRaWTPXRoU/gLwE6X8xBuNHGaEeaUiYdsSYUAIizM0wPjdH8+K3EZsQWOInWUpJO
EjXsl39rgJhgNMIP/gR4NsUULil3ziKZsiY3x7V3OYKg0JnvHj4PCIWY9njYmABCGTsfzNN+t03+
iTAkeppWaMdAj1/x3hDdydVTz1HH/aLbofQOpCk/rU3zD4M2zcoL9DCJYWAoPK7znClHrYXtz93F
Jdy6EUUbNwpzege5t7onz+BnF++MRmxqe4kn5h6GS5OlK02e2TdhJcJ1pupTTlGkcf2vcbJYHWy+
tHmR3q1jDQdRiwWg0KKhGnkdOy3SMGZDnLYU9uoVipAkLiPwzlllX8vIbsv/puI7h1a/otlCf5Jz
FnkwfLRNSR44DwcKpDgk/0NJloJunLUIM5h+wZGQPnYoyyhEtX8wG7gfVJddZAHv33GpN6wh7saV
vA1bbTi81KVlW5w+5hRMu4F5fJMmL3yeZDydvtJCYBxn4urolq0khwx5tsBqGih4monBhXO2Bkxj
X6N4x/LNMPc48Old6fwTjGIHS56hTP7ideacOy7vcxgmppmSmZt8gyLT0p/d3SznE5H5GQjsNT7k
XZRaN0lXEQsdRsNXvB71KNnGb4ArKCLkzWvGkbUsa+uLqkXreZF5FW0fIfu2Pz3LcF9DoN8VnbsE
2Xx1GlBvMUKl8/OcmaVqdc5NtQzWU5+/CSNEEFHZMqOnIizSD6SMfkTZ5s2xv9S4m34j87zYXz/S
e8si67RhGTlqtGuOTMZudySSPKkW5+SZIXYYYBIKbhL81g0gD41Q0Y1K/cFqiw04WQCdymq8RMfE
5ejr5h/+ieim/7Xl0Go1Y+zHF48HOPkNHnVb0OoggnDkCoOKk/P/0J8kRbkAF4cQC2rPtb53sMTZ
3XwsWyl/mKYKpeM5uxvEkvRUy/CFOJSjPMkN1ihmLUUwTl4GU9FqvBgel/gcIqocO4YU77W1E3LS
NTiSSVIS6vBGb4uF/DURLdcTMQ1wBVvnvHsBccCg0Tcx/lCrNDU6aafEmDkzm6dVCURkWrYwWKnb
l2a5yRPjOFnN0ups0TvH9rIF7CaMlMpkE0jkEgSLtyk+fIvqzw2qxUa9zKUOxovD/Z22YZ9YStWx
w7ehYnk13fLrR9s7sXlg4NPioaxLGXKfjAg1VC66RNo/3TY2tfEv9tHKSzJJvcDvlBvqo0r7VU3j
UFWOG8BXjTkpMg0/DmLo5ijbQtb2qCct/hgM1is2VjPG+fuM0+XMYVfhSUW9p9HTzFHFQZMotwuW
lOReWapCEc+gPwqmXdgXotXRWJPB5mm4hrIODTBBfY3incjiy06VHkpy+v+Q3lOWpfGr2o0OulS1
aQbLhdaWixxeUlnw26f9jAbPBmqhQ8Z6bJBQPIhSHkIC660BhIi5z6tT4GopeJpdwLXVSnr7QUme
zvGlhjsGhYEvDUa93Y1BxOyy1mgldpETRNw4ayYermrRKJB8Imul40XfkWRwEJsBNz9poC9aS97o
ZggjG1ZQwLYom4VmKrncelP+EAtslxH3p3guQoe1gvtt6KQN/4id7RRLH5QPM23EJqc6EQO0xjWA
ezxX0h19pwJAbwpqR4BFbKJT99O+lI77BEJH/NhKmNOA/730obC/EXUc3B3oxuPPXmlCfXec9ijM
4hSA1YPNVijHPPQ5vqYeCh3xzIZeZOK6r4A3sDVDKDTvM1+kYYVeLgvKzAr3rzFyh6eR8ZtRQNSz
FFyFxGdQmJiK1t7SI9NNW2Ibzl+w4KZC0FLtxmrsm0K1cFfM0/5UfKjrTISFK6a6thZ4mQQ9JoaI
RcS4RWBFfb67svHXtq9UVkfwjNcRe9dyYVIJvrhZMoKUnGp9y6vABudFAtmbyfoMRNDFopR1dxIP
GCTwUGC+LACgkfiQ6l1tC2+Slj0u8LOz+f5zaW+IEp7G6A2lDoz1UFg94873sA9ZXCr/L7K6ZvT4
2OvFhewBmBYy1hXIOVqdfY9MZIDbd7Urq9ZyeuOSYVEguxg6AyDFD8mw2zIH8L1fmrtnv5B1+t+i
1B8Sj2yPWbZ0s2z+ErAcPmGeDmoZfd+AqiH6T6E89OttztpbIfbBOUoW5DKKmMeQTs7/qKE0vqHb
jMet24nGHM3xrA09NBoq0+OfBA/rrzaWWCVR0cAuDEG6J7TyuAbdUQulkBXq6dG7Ko4l6XYQPeqI
IGeejH8OZ/VhO5ejZtsMlwAPqHQOEzIK1vDIq+mxmdi+rHimxBXxwB+5+EuOxt50OCMbTck0/8bw
FCx/kID9eLFb6L7Pto8OTrjZ25HA4GN1tmSXisR9Bz8D7Z6POfELm80vrDSn9kEcHmtycg1k97HP
xAW76obZdN9b7Z01JjXDswVtKkXNM3FVjuF5eKpjwloFi86Cos1eQYkNORB9cd5VHikMq/dxUc7Q
s+2aTfgSIU1jsQgTrZU+Mmma4QUzSKZnTN0qL3gKuhcOM6RrgvFMTFSu5UmMEUw3pTRjlu8jwlRz
rUFL1lzvkhokOWU2KAYbDUa2xRN1QLdIfOYf+pkGGSRLvV7b2gOI9O3JOpmOYopFyQkdp1W7PQdb
p3MhYcy2/1jYn6+j5kLW68Kqob1d5roFN3pE1C3yuFXwimA6x6JWmjIMeFNkW9lpcG1DJQPRPYQo
nxK1ctBHPAtJhzrMqlLBjE+ciWO7ScQJDp/2VImzydM33e8FsXG8mOdDzS9k+/H2k7316ddaq7sN
VixQxJjVDN7HtiU3clu27FD/2x6yadyDXs4g49uAUstORaS6j+3PE7OH7DlCo6riJX1oIoJYx7Zi
ZrfGJyr0+YztRljnxTj59AVxaQxfCHPypREeKwTGTSSM71Zu3EbTsHHjIFT/M629H4As7mcD23qA
UmwcRU0NBtyJRc5/CBqDqikhQZoLdA6IsJdqz/zheA2+MzxTRxzpror9LHDETiz2WYFGfNCDc4D5
UnN7Xv+YCGmKpGJWhS6cBfyg2vbnpwKjXG3bJw2d80k5qC0Qr8izZ/RxD22LwsFRLLaxzS4huCQh
Rqy+Ne4kcZjr1wZer3eNmPu2SpzKr5Ka3YAjTBuHiQ3LSRKaJKV6MNG14y0J9bT7YdRa1w6Kx1MR
eqwnGXfz/ZRC7KcQHFez7KG08vHcesb0z5fswpXjCjuAe24XZ9SIvawFmGwoPPgKe9Ee4ulnDiYA
38SLt2qlUW+5HbqnVJyH6fIF6ttHVNmtAf8IMMXYmez8nvYGYrTtxwVJ72GWFYRlJnMOdXR7P93+
wOPfUQrsjev6Ons5KF1LfQae4X0lRLBr9ldks4ywb6EKzXmbQM42J5o3AVrWLr1e9UOBDEHlVH4F
M7ED12Nh1O8EYW3ESk/p5vg7An8WN+zm7mOcEYXeWLR0yZdG7AyWs6fB67BcAgVwkIJQx39j/wtK
nirLtjAd0iAGH05Y8u3NZuHwUSj94A36xdy/s38sS/H7FcKqKETNkujvGAOQ/Fh6Tsd053BZADAz
kIub2wwQHupeUgeuod8//7VbNT3kSDv2xTCperwhkJ8eGuhfJ0SfJv6+8Y12WOLau+KipEDlPR9X
mzKBOOB2uKcQ3qAyYfrycT2nQFOEVh3rrfBaXUUebDBaP3dAeImYTySL0/kqQRJcrgiAlkMT79YJ
W+VuPKemQgWUafsAMzL7oO3VIfw9fdv8lQIl7hUIYtO35dvjZW2v+UOMKRLnWynh4bQdbg06Qedd
ljc58DN+vu5RFpTJA8UlFDs/NTldXu8iFESsTol2Iz2HWkhGH6KK2Qufs4+EJYhJ4oapbrXNQxKO
p1S0R+PQ2hNZtsDMaI7/tMK44OEDjKTzkNyuIm1TApqD3HnXcI8UQ0Xm5dVOINr9SiK53WcII0ot
9HOpkWJuze/kyjYjYeZ7seF8kFt6u+XsjZqDKoB7Ce9TlpOdL7nVfYVK69Yvv8rCpdGuwyqave2E
w3oEuaTtUNpO6tqWGP1irSYwAiBA8AlLQQKauECQ9ST+l35FHjt330yPOwdL3hSfz06ReNFGLfdy
0B9uSvBw7RdUshsl3lrRmvMGQl68F80s7KyaiuIW8L1aNUda5arYau6DLS+flwxz5yX+DsY90Gwr
3IsZzD4PhNQnUjpixpJNJBvZVgs6WmxzRy32/ljjR35JSa9+MTJVTiLpeDFeR5cWknSzqkT25EN6
1Ekg52Zkq9amHuEOJcGvGDiUInqkFdNfqe+Glukfk21BFAShrkGrwWK9A3p9+972hdr0EVnxwW47
5owP/JC0rpfCr0GwuiupQtlSqVlki72CJCFuaMwCxaDQZU5stjCNXwiUvNBuwomIV8oZ33lxQdsA
V9rv24oYKz55/clTokhdsgRDEyQB1one4P+Etr5mriqQgnzlmJln1UQ9lxOlcgz+3OKHPLKLIMSC
VQ5XE+EV+Uwdj1Yu68uyBmLgdPZXaloec5kLJq5UNfFVb2YM0m37Rh2MBWR1CyUOm1G+DW/rQmrp
76aLVNz3mwYNsoqiJmTApQ34IMIarE+gadikCtggU78OJihCQgvRdI1+CO7Hrdy9hXax1a+fJTxo
qNYx8o5dcoOwGYszMl9HC9KJ8rSyKuNf5ALgMaYLiQnHKtx0uflXrPu7m4FHdEU0oNDOi8NDZQn4
5Lgz3Em3TAGiQ25ALEA8YBV36iep/dHhzcBM90vUGmS4rLps3sn0+19+rjy4NOflpQg/FuY/bNiG
j2HIQDQyNIbvHuEmceUoHxIaxM/P+D/WVwFSu/oXYGeRLPiKveoOhPDxYQaigBJuyYyNK7tXUsGq
fxH20DUlNJ5TPTjb5v50mkcv2TG4gK60XEPX8GTGFZ33nxQ/vz2fA5myjw8yNuLKN0cLcugsajG0
kZZdqzgljOVZ93CgOB/kJyon8Ft6rLDlfDCPsq25l0zDwAT+7oq07NMw1nyBDm7kQUwSdWYML0G5
ekzi3qQ79iq09SUKoqTQZazIfPiZKI1gAEoy96Y5R069SRIsjD6ChgBAs5dAcNDX5xx70j2YlnFw
3VVa2mOG9zxXWfZsDD8F73RJZ3RAlVYJkEyqomFrITVYWEQt+UqYQb/uupG48ERPNdRRNqTKgFk9
X43h2UL91DvjxPQVHErwXnkUvVc62klaJtTImYAZqUK5YjrKoYuaf1x3NoIrFxegc41tbxFgO6+q
8KWNIheprS4L5PkDZ81xwhekqFAFNhgAwB06smDr9hQ+NXEs/uISN/a781qNsOwbUF8rRPnjNnH4
iwlqoGIA9uuJ3q7teOll8D87+oweJBjpjeato6iOFTofONE/0k6TezDTLa44aP0E/Zb3amCkZtA2
3amzY6AmTDLwr+Zjr4sXKHmynf0fD0p7n9u4Hku3zoIgekFEA3vNIbIfBYSuxy4v7fiP7Dkg6KZe
ykOzXgUy0KfB1k7bokztc9yIbDOtQ/pxkymK8lsDT3AdhmLZBhGfUX/Fv8E0ZJDAhrMAxGkTJQgf
6rtl7wU2EdmM+P8BTr1DKaWrhdZIj4uqVNRc4JyrSkBnWGBnP/lgwqFQn4luPhG7Znv60sCS+ao/
k4qbXC+J1PhGtcEDH4HFTL3pyXuVUyvM5pG0WBJub4JjiRROxPNctubDGo6yBAb2LjmObhHRltRH
ka+6WwRyQEtOlj6HKrlky5txQ+jVRDgCRhqURkvdYI9vwNLr5douzwHlc1GJ9096CclUZ5hTpiv5
7SsLMNWCMKaO9Q7Fc8/8Q4SRwTR7uJF5L/cDwjxbuq+XYiLgS9pYEXBDbHAWT6gHRUIrMNX3MQA/
zFs0dRMeMFmnpR6ELvuTqQJODX3olctUIwyfhyIbwLBgH6ab94wAQKOsGGLQCvPPd3R7ZurUP8AJ
eUHASl0RExhufZQz+j5Gqv+hs1/IHybt6I58w9Limao/Jrmy55jWjgrR2J0OcN3r4rb0B2fQd7RP
isQitLm1YPxDEGN/xyApfjBxDs1aKf2lBTyGSE7MtqYjnHi2WQCZR157PGe7ShJ/2x8K2IPHAmJ1
Jh23J+VyoY2SKMa3y5QSiPBhXDM3pD1YnPGirdweVCVgEyCzwwwHaeEBnv/1GsnpX7A0hDDeniqi
H9YGb05VKTuAA6rzHO1C5PWU8XJnYPrxV48TLeEgeDOTwUDSREg4lL3fjtMkH3Xr/QjeAZyZS5PD
QuvGKg1kggUS3tCx9PLqQp4NA9Ygc4TUolL+QRvi/uSVcw2eawmayW5Fx4WQ9/M82/tZ2ITowvAt
/MCRa/ZnRSf4l4DvaXR9zHDFVybj7lDuqEcDUfL7gltTGkeJcQybgkekJC+npeb1X7Lq7CAQjXq4
T996il2zIy9l7v/4c1nLfvJd5zp6Ymjs74taSDwaIhoHNhfppoNM7l66qQJV+rmXIMplaMop8xUB
EYfIeb4mG21tVE9C90uUK3Yjeu9kslCk/XKceAyzT5X0F7UoFfZLUVVISvI5TVuirAgjlQYCk87r
L0myIVglxjcRbms1Qq9GP/DIMuuoLNCsyefr/3Y7MX7g87p07+ucTBW04Rmt4CqNaIHYtDmAKQSL
gQqSTM6naomD1eQ1/4Hr+//fdwkL+zyISY/NCoC+IzHsbAJm3doTp4gEWHSUIRai4CXFjwZ4IJQK
Bh3FJdss9e+Yn9VZUpvhs8/6Ow/Y2ok1K/Gvn1JsdZ6Igja/uzTOf+jPCvxCC/7/qTHreMnIgw/5
2UUNuTBgAr0rrv+4NfFu+R8pDOsFM4BLZQmXotVFSdrDxOS9Ycr4W5TblklenIZHG68tZfczlEHn
v3VgiNgYNM+Yc+lHJEXZ6rSd9VQyI4s1h4tc/mtyGJVVvHgCEDA6xIwDrphqfFBWT3ZunEa1nwjx
ECDHBgf/6dJ9g1kBgccfFtoivQzUuBzgY+31As8rbILgX6XZi2WIWRD/NBlBaGKJSAN6hrsYyjEb
yhRgCxTbJ4EyGkTROKINkAYVRVTycAf4LJ4bFbjxfdlN76EHX0iwbaD70VssdKCYBEzQD+V63rIE
ILMmph7ZRt7k0cQZ98n8b0lSjR9vj3rYgUqSQ4W/WspvIB9AQV4wW2CXAU9n8ec4b/x8MRGmyjFx
F97CZm/CGgVazDRMJ7Rl8m3UWPlSrnPoPjBE2/D8RR6p7GXSkGYo+9RbukA866GiRFVuO4ejtN3d
XSIRe5XDsoHuv2PW/XrNieu0MA9wQqL3c17EKUh1zhq7RpYin2RKdHb+t3grdUOUksrfu4PRP8M2
5dhcX9tcRE4fOkEgd2LR/ebRbzSdVggLNkHe16wAMM9skAXXCjN18QuDCM1YnAiyRBy7DOnBEN9I
sw+uXU81DygEnSs5sFsRu8F6NYQBPxPd4hkJl4l+1UN/meGQzmgNXhQbKnGLu/wsGJyWg7avQHQ8
3/tvST0sDw4Lr4c809kay1ooNA2qu/YiuzUfdTATpCXAckZAFJFmXTwrMR8E4MpdIWu2RwEtKZ7U
LxruKGkVhW/X4w6pQZVwYK0G6JfAfj5T5uZlQTalsPDCo94dxFpdkx2eN5OR8Ib04uOAOg1NnAtc
wUx+7te3TvWG6WPiCiD6O8oIUOcxSE+svueJDwTcUg7xS2dhGxeEwhbrpp/Bxu3mtjROvmOepDFc
FzUwV+sZJEiTX/sTzJza5DnCTipdMChGc5Y6NSphU5+GIEYxxZA/egFPbqOUWg/ihTsdRraIowPP
Ffd7Kq3t7vafp56F7rndIZP0UBJsGxLeErmt5K4gG4NnkmuWGJ1totxXSJT0fKeXlzOWLsCE5CSE
jVg5PieSagGKhhy5mFmuK62m2NtVH2ykGQSGe9KlHe0lLMMBCqJpJserRCE32G227bjeykgV1cDU
ua8YqS1ji5u8OUjkR9LeMLZuS+7Z4T1f+soQ9eWZwAy0hHmWBNgoCzAkGIaFx02j1DXTOH8ft6Y+
VIvRJ1tZhusBH3ycmjqxY3BonAxqgdVpIzZVnx4hK56KagYL4kAW0Yf1waEn4i5dSMNQJpzZPG8K
ZRL8Iy9w29rkxxgR8gX7lx3V+eqIbcBz9YfkpbXoK9Bcu3BEFDxY0nVxoh2MreKSTY7H3psmhj+5
6pQDfEE0F9qjpGbtWt+SOgqQPopKT2iyg4XXwV82ewdCAge8DkHr2il1t4qAN3jVOiPXctHl/QQc
Bwgvyzw1eLILdx07NpTi9a2KzUCIi+CA0ld/4Npnq67j33RqnR4ZCG+Q9GsM52uR+Bayqc0BAYCK
c4QgnUDR0Nj/4k4yxPxWSmLuhL0aE7+1GuI8QV9nMWnFrvFSlLpZ9IY4YHEbP5XT0zLss+cR2rfn
e1uIst6at4AkVB3DdIbEs7PQ44qLGt0mAN4nGxBgVD+40xdv7Rx+sVBm8BFZ+exHRVHfw03qwtNI
v3h/eOt8cMtHcAJJ7iNFxCdKzTq+M3W16ikylBNLUxJQ0WOIwVGb6aCSadRUh0G7Qvou/rFHoJpO
uKOreY5em8ZEa4xq+uh8PI6hWtU4X4n6TjyNKZmTeY9J8tIqvQumuG1xWhs4bYU8Qv9POvUm+LJM
n+fNP4wKznJw0fki1pWT2m+hM2C2ImlDkd0ibcPSRfgundB2EAuxz7RIYRL8BvFSYihtyqa4af13
fJ+nKrStWy1b/L+SfXWL37TPZt9HoNCSFVvnTZ7Ai2jQbjhGXO29/hcEwe1BLCSme0Fcu2sFEA6F
OgZ2uqUJM4EH8pk9MpzASojgN4ajmPAp3MZjRITgO1MVcvhvLVhb2ZnPOUkuPibb6RfCRdNp+oPJ
BswsNbJjvyvWGEcMTMFCF9HfNKLd4oyOxf+18tJaS3zGNaqCUphFX7aNrDht1tE6iXzDV/4lYfHW
yf+BB6scuMyjuv87eMcBB7P0IZmhUWnPOAVcAG5g4JjxxxOGvXdk3q1AB8PqnNdOEZ/RNFbayBcO
Sn4rYbOL+n/tEjNL1cmMMqcgENIOoKKBcF+g/EMO6pwsyRVS4KaG2oQMH43I3m57QB4TNlI1cbpi
v47CYFZW6IQf/EZYu7uhp7u2/TjFdtZBvfTc39R/YWiAbhd7ANEpUXt+b2MACRQX35a7/idakwSa
pMpMa43vVNMXKCyK46+IXLYWhJJZiCYSTDXLgUybV+x0hAlQYKh0bl+1p+CS4Wch0VKFGJBqOrir
QjMWwMKVOkBasyXHeE70AHALTioq0AACPg5+PBdTyH9ltkXNNWCC4fQDSkEqrgfiosEJjmc61cYT
UjD490F9T8U61XZHCLZH20kyqtujKFaRZvpKaU+WqoLOzCCqckTeDBJPalVIgGBVeo7/vXOrERNA
uPOGD1kKibLaHwy2zDHEN+qgLF6CF1lySh1kZgATK5pbjIT+f+l23b8ptwT+LyRYhWpBHVvd23L0
QlIoqjgZn9cScQb9YOYTs+Wh+qrW+PzOq7OAohWYd60V2X6BMOudSIRHEpbWoaHDLv+nP+TBMfQc
4JUn5fEmnd71wMGP37FJRS7t80wQ1fpdyhggvvX9Sb49dNzcidGXSIKr5ITzqBgKf1jY0FdiispU
yoWgK87GJZDwlmgCjlK1/PbdOLfXPSqyGNUlNNZWsUH8eB5ZxNjMlAm4xDCDAJZ4WgZAzGOkIfel
kiutBYqjwT9pW04sEdZfBkWU99TjQ8HMGiPZ4sOJVXyPnMX30+VGz54KKCHRyvWJ4tSIIOZEyEFH
mWTbA7zBUMA2CIfTxEKteShrX5nqD08KbrI2aN3y+OkGFS5pCzvPH+RXX2LRSQHoBDNFOnlk15qB
OZIq7Vir+ngTsDgK+pUvIbf+3Xvi5TbtefHIEFUw3HY+mrpoG8vpcB8hpAI4ombRqE+G5Ab/ilzf
6eI+TJumqpGwyy4Qfp3LEtDZc2i8dRo3IHt0p9/hiZxwSi5N4d9KmTuR48vB7hxiSdNNXs9rl4l6
hKK83uuyOB+4g7/QOG3axoR9jCcDLmWyhRHy1B5xXoAfWQ5SBM1Gk8BGwLSNcWvCt+PZPTvv0qi9
lFS8R3OE9hRjxVqufecZ3V56JZJ6uf2zRAVlVAJpmxE/FJn8whT4B8MQEcX4CRSjDEu6sQpmN7eA
kN8RQvirwdd94kfours8Mhd+H1l/lEEs6/hxOqg58pDolzX1/XkRURnvhuuQ1swMBfpsIYxEgJAJ
3IAtaJ5MUpUMQ0nwfBuNLx+1BAvrRgfxpyZDGqf/r8QYh/m4QLHguYMXRGlraohAStRdmqISTLh9
s9WzS68aeud2O/rZHubBTb+fXRKUICA4lhUG7Tgdj0BZ46/AXKt+3RR1dtH2uUNIwEduvZR50kgU
MAWqahfWImSv9nwAgJfN802YytMVzBYr/Mpc74ljZXvM3X+c90RkltCkFz3mKIURaOPUQiIaCXTS
YDd+2LQvzPZYVFhjnWw/YQ5/CKu2DuM95FSoknaxwlklG39rM7zyAU+G6Yxjr8S7RwUH1b07PPFQ
iILA1MCCpDVtBLcbtic3uIwpk6iHsWaXyFhNN662F6RuhVKiY0PqC4ukZ8xHAJejlYiwaumgEvhz
8egiWxdhAxR/XDVUV6AiitXDARMsTgyjcscQ9VkQpqujrB+g9wXvnVliWcCkv2/sG/XlHmAoDtFF
QIZgLK5IIZHncD7nrFd7LsuqZHEPH1IL25sihL2Nq8nzJ2zOw9kjC1ervx5UkWDBDbdlFzKyTKMT
vkC50aS+b30J95WYS3JD5N2w8VDi+6ivH8L7SnbC8OdZIpxYaQVz8x1smBaynJuHJhRqSfnJx4SK
cYSN3ki4iW3Y03bSfz2ltCkcFe95ChU8jKlT7dDzzwqKsZ+0YT7V3i0I6QWr4yXG5ZoxAj6H5jfZ
NLOKOz9/ANzflSJVi0D8Z9S/+uvMS7Reuf6FkAaE07xl6LAIVmwQnusxv0pqOoArEgnCzmmXfzNQ
d3OeHpD9Cbih5O8qE9lUPaO0eO+2MtWUt/uSBSYZhpbRVdzLeG2V/4zT++P+Ts5MOM4ZxIGpFXC1
Ffc3mNWCD5owcLz4b4bZ0SnokZyIzO9KpfiRfIYxnlWPpAXGr8/3Icq40A4tQMGh0nxkVfXcb5Nx
gqZY5xefEC6hkvGIXoPI1hwCWbily8TPoHSDBzOupn+BUP3zlpRW7qJzVbF2Gx19BvX4yBOOBIA0
A2iooh6Y/O9BeAQPRjZ/qnb8fuOEuKmEasNigm/T/frvJTDRhDiFlIJkjn4fLsUkCEulLLUg5IWt
6y4Y5555Tf/W65aF+XSq6mtXMCJ69l49jwcCJ1vOMPBSi55RTmdOD/E/Kfe41QESEvBoa5oXgTaO
8T1A6IKlDXxVGE83tHQTOrANqP807/jaQeaWeG6TnOGzVQg2qG5yyk/NUckyY777CbFmqgDmTPLO
rpGUJy8OZFJM3hbtySZeX4UNbH0Tm7qJJNq6loNJ3qDHcqbayEhiqzvxndGukm54+v7PthC/TPOm
kYErMP60TI37EB6xcxFnKRakBJq2uo0qI6sJIs5cn8kEPWdCBYEHNTntsRBdw+DQR8baqXHQxehI
OuENAmKDFv+z5nKWYGMgGXdu68cRj7fMWyiraS5HBuR6M2nxJr7cnPfaYVXgIfPGx5y2snOLx6Mo
7Zb+ZlVqrlJKqBxbFSUL1mZsMLW5FdcnD9lV9X3ylnhBcMuvZJ4TGNSyd6pRQG0YjJ1pQq5gzbBs
CDbDu4CTn9vC2KkFWuSfV7h5SHQcgXEAXzisvCiRWimyPQCbbtqwHtfRh50Ur12nykEjcfzXj3nS
vtYG76oEN8pMCh8y7e38nZDVfJY+jfrYvfjevs77u/PZyLCwoRuqJd0yY/2mXx0NOTuV0BGfSFsI
M/6cmzUNjpGVUi/alEiC30Y7eWDm8D10+TlTG0g9Y2cdjQyAHPYVq5KbJV2YgsvhuKvKCTgAHKpw
DRc1cN5Qt/XAUP9mZRB86999L0ibP0pX5Qq1oYnGNFND9+M3W+QFv354poj2Ai9d/ffWGQ47s34A
QdGP/iv7/XQJlisWNZPG1Cc/mYp7PuC5rtkQQfxKigfONOJ/1scjEQG4hndisywJbR25qvkubZIj
eUEvQzYS55fWOQlU3HVn2GmbT5kYxS7jBvU7yWPOBEGfuFcwjQ7iXaGoKfhU2hMkJcifmH+LCZe+
wEO/drBxc9zKUJz68oSZKrRinM8+NrnSScsOZgCgOs0eJ2n5kAqTD7efpTl8BModTZ9TMHDyFqeb
tdX3hmmtTb32LXaXbgvJ7mOZH1Wo+FGY4J2xOOAJkB56WIEucN9+1MSM+vvaSbGvIXLWNlAt4v8E
PzaR+BMc/sJObH/4ObzZrtrVcpfXnl7wN7e3mOKHqFw8s8EyIduF1SxISww9yFUvrZ6YJdYcXJ7j
jNhAotf4V0cu7s7AbILty+gTujMCYetkcopKiQrBl/i9lCJpMnUyxAfKi+dGCWhPpDWMVcrpnnEn
/7mbfrOZ00mad7pFm17hAFc2kG0KogyIjYdhr9VjLn9U7S/56Ord7Sb5krBMc/BE0ESjYOeQgrIf
DOexufr19KZNZP6ppOHFTHsK3EwHMXbUkZu0y4NUwvVd2It2tM7vRFBJs2RHR/h/y2aO22mFJhdO
zYXxN0VonzOo3WoR3YB312WeLSnwk7zxnjizu1p5Pg5tRSeGFEmv046Ihj6rzLsaQUfAAAGARG7P
xSeG1SI+23tIzBjZ3B9BDOIRzAi0wldyDaAbwIyvloyu/eaduXS8A7MTsNb8cctAJot7hkTUf54D
TZJCP2R6rHJ5TqlPNIg7dXKhy0MjKH9jbFd3rSepcdModcZ/CBkYQWXmjKfancUlIqHsf0h6iSWh
lT0DdY8CX66MJZXaNysC5OrMMfOu+Sl9O1X41d1omPfvX7ZpVo2wgZ/p+GNdPzZ+LUuWdq+KwlLv
tfVljcZYkuBewpXmScVeQiezCZru7gMPY67iWxZyVfMRDJ17h/nRAZaROUTwfi8lpY6rNEiUqloj
8CAi63o3I/QbErO/or3eAuz39rmry1rqV7csAHgG012u8rUe60tWFO3/A9K1qsB9u5ZqnTMTmBiN
ySGg+hDrJENleW8LiSjOTdoZLwePY91nE1zHt+GGwmXvYQcxHnigF7CRdtNAUCjpnBrL3h+gIB0s
jiwcYSKodsEaH3kPeZIQ8m1Sv0P2b3wEXS8SUu585vDs7o49h5LpDZwCqjL0wdHpLX+0d0ByGh5X
RQKC+zErF9OT4drzB3HQFmG7rg7ZmAknRSo5E60Yf9zCPtR63fRzOwUYSLFBeInl8rviOpk9xoJW
/k5F4ZxJesjxE7LQQR6CLHySUw2XB8kXpEMr+iAWkVH0//ZhuOnRKf/5snAaatrDSHoq+B9qqMoR
dmHpHPuA+OfcNo+agr6QhkR3Ck0rWUyGYRq4PP5Pll+s4cmV5gwrhJMRv5Z0JJMdnMsFV2dxNDrx
HFxvJfFsRVSvHbKqZZ76YcCaWAn8bxR3/PkP09RfrQOeHPJpKSGHHT9+uUvO2TKSJhqXZEp4ibK4
Ci2IgKytBZks7Cb0O4Sd2k5IcyrP9aSFTIGcqirigMeeHAVvQfUMM12coVl4JxEUMUpwUSdpAG5y
WvUwShS6y91ahfuqcbbmsGWugTLSLlE99/Hc6ZZ8sj7atCMtBTi/y940O9fRDJ1v9vYLvcJ98OBr
P9G0lKEtkJYN+lC1oGYeA3bkCy6U2GBqCPf1HGHYsoRG8cIkhoUzK0Z4FO281pV8XX96lT8Nc5qS
ETYyyGgezGAnpAoUhvBfYhpSS5NPLedVeL479AIhNVnHz9MRPwW2OUWmqU/pbnHrF+U+NqJM/F9G
B08e6cvps0TWVaHOdpdF5J/76O6dWVI2pg8YZuv22SznKriWPGKW/4ECKmdYW6JjrmiBIwu40K1E
Fc4l+CoEk+R33FN1Mdoeq83de88mUV3i8HBbvFDa53ZfZ5AwcxbwbbHD9J6ZUBksoF6RVTs3AYuV
QCW5529efRvy8Grosh73STZAA+0lGBXuWlAxkQHjTWwddteAOwtkMWdVWvX54iz+gLhi5lMIExAu
y9KfScMAV1sCYD4ruu07OIY3mxQV6IJVvuIBl1sJrwPyDAgzVDm/0+/WSF6HN/qHD+RYCCUhYDHk
uDZfxjiz/Uh8ZXa/Z3eswWQ6gau48PtZB+nkW7/7yjdXo9B3+ID5fgWosADFOILCLrm/sa8ppTof
AUW6R9KQASMXVZpp2icTPJ6AHVWvHedPpC3ZEBlWX9l0ftNN6/tn+EPmY2KancYW/2Tq2s5KtOHo
kOno2JHix+JhsnXK8g09j0BL0gB6nwe1gvFNy7vrUBZ8+3D16TFouc9BxWiLtm+U4LTeF+Rf21CS
4caTMfkIfD6XqJPD2I9Blwdp3Gt9TtElHNTgUAwvDzmRYmPjmvagKWwPXe0dmT8VAQi0DbGGECBg
L8GFYV+uxLQjk/ufG/aALSjtO8sO51eNf7tslihB39QocvIXE4Un6aH78DFhDQ9vcPblek20u/Cv
LEAeAw1rjIOejfTbuVSXrGObgM+4cUofy7keC+42zlHbVKZSsIZ0R+Kr+zfkM0lVIFyXDGPbEkzi
c/U1owEFfpyw6vHxwpXHeUxmH+RP3b57/sLPyqQG0eMVNIYABIlYTNDMjRUnVRSUVjV9zh+wXGAS
pXrDB4uFc3N3bd67VC9pduhe4PboznTEb539+fs/qUyiZPSLA6f3fS88IUZTlhKPcxF43YRmzwC2
WfU4Bxnmg6sIJLTE/LuDsr7h39/XcfBCw10bbWj4vh7qXX07JEEC8fz5DCOPDsB1l6XrHaSh016w
JdbIV+fOCaAaGkU5isIy4Qv34B+eYR2LM8rhO/slPht1T1xw6Te+G7v6lg1daKLNrFvN10isGpEq
/Bee3BEiLX4EdicTVm/DyDZ7qtTCwkMpKQkBfiMIVwjayoY9AzBiXPNBJ8GqJJaQv0iwrJs0lECf
sGVlLt8nGSYGFjugvo4OpkWPdmO6tA1DVBxj2WtSaEkO9p5pMCVs2TLZz9kUKDvk8Tb16wa+OI/n
8mhZZqF3OLvC+JYLFi0TXkxgXqUANBiP4FrpySmnR4hm4ZysgpIEb3/YhQiZLCA5q5i8fY9+KFCa
ql44xTLRZCy+1ieF5rq19SQ+98ZmTlo2gfsDT8Npbfp4/dpQ8LuVEj3Be7k8jl8punBaGSwgikdt
7SJsv/nagtn+lWstHl+1gnpE3aqDX5TFnt5QzFJoRYErfTcpDm0KzVZMFK4VXrqSh1g0be3CeZdc
JAmDL68uFBsnLNrDLLDsfqK7KlrGMirGFJxrHsaGZA2PMxtDK0KMYIdCK3C6Fd+znbPuGkyescNg
euD7mdzNh943HcyDBgP73brBDR621nSSoI4633Q258Wdv9iSYt8TMpHP/dDpAK/RELFRnWYSFgJd
MtTdgFRhI5VoRPn8P9jU46x9xmfh8U90xgYKwOzbZ2uKdniWxsOgQCf959AzMIzQKFk4a8yq/YvX
JzXWDO+L0PaDw+lR/aXULWLFH/RRDiZLS2tG01dVjjvYbsC3zAh2g8X8jBMZEYrSKLzx2qpCRoNr
PtIskLH4sC1TSQXJg58xZcZ7cSGOB/KgkDET8khEuXzs6OatNmDvUIEpP5gUGn6Sp2RnwZxWZrL5
TxByi66cT20tp+SixfMW8Idisz3Y+1H63mCESKLHlP4nz3gMAjfQdrxQ8MrbELEb9KXnx4MKuSLL
ivhD90p83lYhmVeWk864rHlJFDwL7eB5Th9M7HnlkfMUwlXNKKCgLfR5wZh66r8DQBgWZPhCIAQ8
37Top+/8+X7DCFBi5C0k2NrgZZxRMpITUPDv8GdK3ZCOykpGLmiAOsox3FLrxOZ/AzIUQKvMfyKI
Km1i8Un/CH1EUhFSou7FleuDPh3K8aSj88YeRr8Sn08i6RQ0/rsBo4ZykW4bN1jmYSwwX/5YtK2W
H6vkn433eV+fygQvUpuTII9bhLFpRg18Q20OgEOpJUuQ86N9dwSXsi7fs92xaV0+czNQIo6q4zja
UdSgLD4HETtpdy+UyoEJCTCsaWpi4jv5vKHnZ/Dyp4H2HLsdcDPURQ+ivHpXW2Oynaern8KH4Ua/
bMZ4yx6hj9zXA9bYg6izSJyeFarBygDjRAtKisafKjg9UStQVKxSSseiYS7kxQq0hFVlsSrvIHro
pFfyZQTUF7ZqyQkx5d0kgU2vvg2II0u8DMDTW8/eTFOG0627VWYA1rk/tKPxGLrchR0ixgm2ORQr
Iy11zVmtL0uSDJPPlSiy+Rc2tx1HkgiCNy4pH0S/ZQ5s06PbyTY7u8Z3lSOyj/xwoIhFoPb9fIRD
aB1h7tpp4dCN4gwhss4myaw34AMlvBOazOmecSZaVaWuQRqXQFdF9U7hRRgaT0A1cN3bT+cvFzNJ
BzsInq0K/FxJUHOwujSRk8PF781ks5VgknyKWyg3O2/IA178zo+lbnnQj1BAwP1BeQ/hzJ2C4yfs
UIxEjZoQWgM7nDQmWVfiLW7EqbyQRGZo9+rX7xLDYdKobc8tUUD4TX3E++kCsbZBXEmfia2R3Uxg
kvVZaoftgSLtCj857qeRG53EfOkhCm699+W7QkbWpEZnaiQy8N+LW4/WcjXmCBphwRrKOSl0he9q
IyUWuGvn0jwB/OBcqZ7a3lbBthRlj/9Xhf0kOCRKvoHfvEI9UGuVoUKSte2xBf0/UQJna82Nv2MW
xspxaUHSBQU/TliysmWeu+uCP7+UhrJtv0WiqN+X6Uz2fYCcBf2dLoUNaS+zRYi/EXZIBC00HphH
CK8rjioTYHe0TLuMIPJNXNUA6qetmA9YKd1Ca8pajjQvIa2BRXAfJdiHb7QvDrcuH5PRThkRYrpO
pWSLBGfKuC1MVU4m809cmMRHwb2tjTNr2O4uqUPTi01dh1lKYRh8uooggyDFC7YOqmBn4lU6+us2
zwUnA7z0XxyTyPHgG2eaym+P93fIhV78xyWS1PeoZCJcRpaE/qFfNUpRJwN6cklEe6CYf11/mrM+
NHSFTFsxEx9goN7OfxCnctmVT3eZnyPKJ9xJTnx/z5P9fQtpMOI9h/syd/idwbBOEee0DXJuWLiR
KGJuqMxvCZHHGc/BSZTZenX/X5GBVsDQfBad6bvI9jUOuT91scfytQRTzagqTYuZd2dvY9KJavVT
UyRFLxCmJJDFJBm3YMLlp5u1TMGwrtwSueWLsdym2yC1CQvPNAJAMAleuIbMSR4up/rSN3cSxKRc
eT7Jew/J35jQuFxwTUmlpjJgGccVZNn1OvH3uDcZ3nD/+tytpHyOVOTk44JdMEKoaRF0KMyygaWR
nIv1WjybrJbQO1lSuWb46ceJWPieQrzVfNJsEysPktETAXCtwdtd0FPp8KXkwlVIIj9CtXjYGpSQ
3ldNyGCDHLRtim+y9wi1U2vb8HTfS55lhIYUmC8TeSYSN4LEXtizlTe6hvGmkS88dxzVXIHFyglN
REbp+QHkfKIySNP8KYjBmJEW9ksKlQQWTIwSmE5+7o6nz95n2JrhCu/DuD7+0nrTntpaXfTL6go/
Je2JRqEKZqhEpBBePNDKowrH5+gA8nC0/7DZE7LBiFv6UhTdRgK2AFThLcBc7cCKVEI/EzuX5yiW
ydD4QG3tftWKX0arNYdPgNHhXkN9R4bOAC/JuIAaQZn3twCUB1/4lX9rOd0MD5L4skXyhaeyoLy0
sGOcg3f57F/Eaext/Pd1IJm6LFGxGthIH/3kZTNbT75z2Y1gUzuEKLC3oaOFUPX/dY0jsCf1IH9z
eQQWlZTDzNIx27IRCSRvHtLMW0dNT5kMyjRQ/pb2kt+NxSaLEY3JHFiL6LQxVuZ9oAnLoQZmJwPd
a6SQ9uu5zYgRB2CfCW0IsdL7YYODpVBTuthQCJ7i7LnXXfW3KtvwUWw9Fc0/SKm6x4gkn7Zdzodd
GTKgAMDLHyyYieFNvKSDlLGZ5e8BjpwMFLWXFbOU5FUPlFY60+0O9dIfjL9USbHZlKy778XdgshF
SvGJb+syJKayz4WCMGIY01z9x03KmaImoLg7DUAeKNsymjjjFnyVyD3uBt3/xuxGCWk0UESr2GKk
OrpUpmGrZVljxD/Z/WDj4HVuBlo9fzbqfBEWYDVJNARd1rW4P3SFe5+yENkYLCyMaHIUhxU1xk33
KLW8yl+W3cdOREqz395fFRvJ/x0oQ/VUTHbm/iDGumY8IztXh5RMlK+3B0fyejEDf2dIK08jJHwh
O970UUri5R4EmpwWtCqQGsYrZf+RyfoSkejnDVT+M6rpvSj8RSQFRTAtWIZ4XjtQeM9tsACViy+1
7cDGpCAalhLaPoVc43J9ENlFrM8BrMwX87uPgpinnqhQQHOx7gGwC2M0pn+EU6gIKUddewN+R+lb
6PSBJOhbpX5oGDAJ2c3Xpm2Tk+skNzOAtQwD9k2WECkDTFW2H1GNyn7rgWMsLB6TytHVkVJ5RELH
uvwM3L21CkMqLIWpa3HWdJ9/Gr0FjLtgm78g9/6+oKf7kv8vXgK2BcgtYmnMEAVrnP7lAsyN/HF0
Ijd7q5CQQSEGiQAFfNL8DGXKIpNEzBXjP2rr/4surGdYW7eog1VEwT8DY/vV5zfgWsoaIQ7GvEB8
XoJn90LDrW4WVuNYM2HheeyrPyXMcYfozqEtzJKxcw5nOmzBEkG/Af3EKRI0lY5diOtw4FUQ31Ll
KJ9yv6dDwb/7rgO61k5v6q8AdVPVDEyrH+IGE93WQoiaG/13jpA5EwEaohgA2ityIBwNkGgwT0d2
aewFx4Bc/2iPtyS6ebOa2UQHB/tpKw1dUzzqd9lvid0ysoNQ0DH+I4aTy6H6fA6Xf4MsbWaRbWUl
oLBXgt8xPEeBKEWlAi+7f+f+ygesjzEfLG8fbVqYGG4aTnqC0Z79dmnieegW7e0YtrSRdlGLh/LK
GkZNnryWPVe6RtHYEhrFhwOrrjQIVARE1roKt4jVtYj28Cwir9QAQoh4HJv1TdqAU2vdQpzsPOJB
z4anwDk1VmnpGDsG56s46e7TcxIi4/vmnCl6ORKh52jLWAUGsmu74Cl5UI7Vpeb5YnpIyjhtwXkM
GNy1SwD6CciYzrskO+pmNezLR5QWt2zlgQb7MOPoXVyw3+CzV23kSGaRPVtN0T1AAmqWp0faaqS+
uPK6PJlagZGYlsA9Fz3MEO9Bebl30YASt/Zwp61UcD/I5cRcmX2hK88CNDdOL4c6e3bXyGWQqxfR
hSOxTfy6TL5ib4jqs+lAQUSsloYFfiwHzc+HXjNkKrbU9D2RJuSTcmFkMjMec/Q2zNpCGfhSFy8Z
XNYVnf2Q/9ipBn2GC1kM+Fdp6xFO87Dl/qzeFrFt/QQtwdVdTfyILl35jj/2Gj9P5rfMgxbVWvIG
H+Nyp10C1xTdodmblX/xrAFB+IQMCTHaKTO06ctn2jpGgdp5j7qLiVEnHPyFUT7ZaXfKYPQqZb5I
izah1xO8z2j/U/NuY0oTBIClzDQF1Nb/nngG3FK/YtT6dWO33JKPLQJWn0iE9caOprLYS/L7sdLX
JnI1SCD/m+Ef4GBzJUgmJ+RgbY+6ka5huT/dzOGUcBROnWi0PUADVna6s+S7KoeZxwsk20aZIHFy
S3fZsJNrBlnVWb7w3uvNz+pvOAN6ril3GiGpzK1gRz1toO1mg95ZQhZD86A0+YjU4JSuUdKdmtEV
zIP0Y95pWVIBfql6MvuBxaL5U5jOZsZTkmXMmJJM101y6b2/wmlDOpkbD8d0p5ew+DA7QJRuADOK
c0iyoJQ09zr7FzYE+QKfh4MlshUBk3SgMgcwBqMsfdmZPmH4cGb165vc0ngOVEWZ4v34DXRXzurc
LU+2YX2UaOzc9L4ZDPqFWnT2bBv5qVJcG2sf0j3GkEHadkQ8eLP6KQcJOZBPAQPQ+jM/pcuKHjJf
tsyzYqlz0vCWezD2N5AxFhSP/RPxQmbeMbwkYEiaQLoIP1loLOQHEnjYacHLD10PhRi4kMBvTiuB
hvIqA0rmBW/xskA7mIp/DMoMdSQpFVLvOWqvbsrv6W2nDJeSnkmrHP2+/E5eLhj6YsEdWjA7Rg2h
B7P/fbXFxTw93a807Bn7CtFg+2YZQpVTCLwBl7Vcp7UoHhYdg0wLIoseJzz+Zk+Yu2SuJu7A3RRQ
x+ho8elJnPMwhjL8grtr9qseHQ+0L/QO0MFUi0ND6EWX6musqs4/W3fsGcFXDPl9yRp1ZWDHwPMG
uQRrUzj9Js5FFgGDEZoY4ghyiIZwN8oBLF1I6yV3ugfCLmQ0a2/EwTk8yNpTJKh6V4luorPhiZBS
iV2b1tS8SpaNKAdvcAFWcEL9hlb3ZZqzS9XP40/Iz+6oqSf6e9T5PLCYadz83Q282QqFYf/hE6r7
K9lguue3h7YyoeTl5ir3Hy1RSYueqKzDWurG3LgdZJ2feeKbL+pj1Sk935o6hWvB44p8Es7jTfXz
rGpkP3cnBCS/o3FSTRISp3Zrr+9GfZr9pCo6LpXfJdpKzgGRYlElfeDxH1QrFHGN6D+xDV4geJ8d
N621uhOfnTGWqlE+j9oSucpo3vq4xUE4Ize4VYptyiY3VJtBQWyv8VxDTjbeMW2q1dBlZiF3MxHI
owvr4JpZqSKD3x5k7JraQLCIoDW2Ts/B4d6ny/mouBhAs4it5ERSOizrU21COHtiB2TqKlUGA3gr
g3dNmrg2pm5gTH600ZtksQ30IcoOom2Qfi1Jag7858jdG+pU8RdUC+V2g1EqTUbgFl6OEv5OKQ3o
MpfM9lvty95pI/9Wj3iIilyqNQlOwkX57rl999kUBM1UwTs9wHl1ydrF8U8k33j6CUgQBSTfuAeU
LCQ1emyqVzsUNSD8JUIs/8ItSVW+vk6c8b95hPcNiLXPSmKwZkPwg92K679KZnUSmMIhZDJ19vh+
x6rA8Ak2XsxMa/QyPJdBFwODDBFllHk7WDkN0ky+JfKJB33wWYByOP/vsVtWNsfe2GntDXJ7Tjmr
s6kfxWnke+MKHg4htghpSgKZ1u+tj/TD2yZ2GLR0gC6oDoN87Ylh8ZIV4mBN7xlrK6rfQ6hhOt4g
AlsG7oqJsUY7WFubkSYnCK1b7I7/uAKnaZvvnKn8EsAX0EE4sUZKX1X7Z3V9ZnlNejt9/50sdxqY
FEW5H88du2Gtqt5wAYnkyw4tnRM1YCSc7rzxkfWPWrvfxqujN/5ToCdlTjOztuAkOc+Bwc/pIdB9
W+YPqysq42bCRenMwjwd9YDi0xnSyXFkhJtUgoRQ31fK7vIwxsXerZe7RmN1FPU6b4KZ1Outx/5V
IVjHNe1fdhOyyU/hX/vl8QQ86YIjQVV6rcuhMdJCmVvgDPSZDduFiYbxKHlstD6DEBM4/CRHGlef
fTDFhllQbwHK0yPpyZn36h94y02D51bnj7vCvS2NtgqY/iokX0ZmRoK/9brHcZ5znq7CQmfUIzky
Nv4p+PIBU/h8Sp9CcR6wUCmF0IQCOI+8FTwwFBLV7V8vJ7ml+VWwrSHb6dD25l9uP8xYo7HEyeYu
BQYEPdQVy6yX8DpIkfS5uPlRpLJ5S/fUqCHTo5J25CisXubQlXwWDR83aSW968TfQ6ytSEBdYpGD
6NOh2boB1ZaIIQQzjS1i+KbiLI4jl4230m5sVvEYK3B6p2jpJq6OcKZ6WDZr1AE4r7yPh+VBPWA6
DjdKc4BWnBO59plUbyJ70ubJW0AZAvdV5gvalBxRCkjw8mJB/M3ChDPUu6M+1uxocitrRorNs4gZ
zerpOpkccQXkNF8ul7o22SNe04RrgydOUzpuwY3cIT+zIWHJerZqgVtGDw8Whd07Nw6v6JOAcFLW
H2voGNAbzqbNLfSQw9BZKlDA70ZIx8hk8uCi+hCgh/7Yc34cQIVAIunexktRgoG+Jsxy4veubG1P
NNaJLB89POTbn7Qo7mRoClB9bd3NvzxffFHbKzUSYttFzSq68C413uFiTOYdgeIE7t8W6e0x61hK
iST57ctXlsJtzh2lgaML/zk5IwzpktPgQ16LC5zR5HxT341Rul6mCHxskSCjk1VabWRjd7gsHeQ9
hbyWC0lRnUycLelm5mKzXwr3BRqBMrHMTmZMv7MpqnoSw1txHNcTmjw6rL/B1mOj7W4mYy8ALz/V
bS97eUHiGI7Do13R67livvlqs5E8JsJISuRbYbzR/bqu4fayHCzzEGalc4ueWAnvq0D8erOhB2rE
7VsjZ5iZ2IQovBn1bXbRDOtqmpvkPL4pz+U3pSsUXf4OZ1idxGxeR3GCzcbDOOx0wr7fOWFXd1n9
eEhaDnhYqC/ack+fZfbeR5MBEz/+bnS64o7g9MVxIa5/mxbPRkInyknm6I0Gufsw2K/cwtR1nPCm
lpCmv1cL3FpozUdGPDR8lep46wiDwwdmvnjdildV3cIiPp+C9pfETao6wxtmIvPuXP0S5ZKhq8KB
8m9MDvrrKELlPaI2l0W0A18TJxR0wGS4oxpL22INtYvt81UtcRE12GSSxRWu9+1QA4+Aee5ci4bR
k5qKaus0ZoO204zb8HOVkNLNKDEU3rEfdq7p3dfYAL6SzQVVrfgfwurLDBmR8X2n9QG1nx9mG5em
3kGX5C9tXdGb8gTkoECk82mxkZUrKHIMjfta//dmgaIgCN5WEynYaff31SrRZd/1Fwq5bHKLgIl0
eVAqI6lPQ3CyHGG4eV7xXdPR6QODppVOWqfKBUfQaI+dljqY8c7IkOtqisY9nzq5jsDHQkPv+PJr
EiVE3ykwBeHQevqbKNsTwWyWjS9r0mveX/bW/CmP8v7WWxGlvfxdiSO4CGiSGHaPIcps6uHAQOzR
wSQrGM9Ofvcd6277G3Qncu19XSjzAOAT4cCOZ4mIPo2aasdf+rWw6NB1s6LPto+XfNb9FFT2xHS8
J/5ha0+ifXOQElXKAiRdva0Cic13v5pERlaNnGrkhLEza+9UJlnVDvkM8nUXF8rTms0UmCNSw8AA
vymkmvvfXhmtXPmtsYtla4CV5xz3mnl8b4BaRSOETO5Jvkst+hBx6umWwgVUxnrdjdcad9eV/E/4
tQsK0KUcWWAbwQ5PBEtbVOLd022/59UwCOEZtZ/+ThRSzdVpUU4BI7GuMkmFNtvoz+gR22/l08m7
r1UNVIWINXVPPwgGv1xLnQIi9joQKiYQLkL9WwG84Ge+Cp0tyEv0ptE2VZAAENXHZHImavB0qDqa
d1449Mmx8mM/U4/CfqmlzDQoBYUhXIe+zTPrEXyUl1H0yoGkuIiUmnPFN8dgIWsPheUU1ANJGVeY
6WJLqFdJVa+kggIB2TTi7sImL+Ogn3EjT2h2YzX6CNXxfIdNJK0563ak4CU2hoycXK2DEK4OvlAU
zMglHUU7yhCcc5w5GjrpYmVxGQu0y5SVkRU+De86cUzuQTwvS09G1MyFlMPtMWBM52MvtezGIMLA
pyABpj55eRf7kRy3WXRkCbCgbbPyfHzGzpnOoLSYsztLMKDvg63qZqZsVq95nWZ+3rH2At1AkGIb
PO1d/1eBk4xU203YjZTRWa7mp5F2XmbFXIsH76scfXINUpB8kq/bmhHvOypEOqtD/nbYNZ2QT21j
1Lx6yPhLMkfDEu3XSM9K1sqZdqizJjHImgMS5FmdV286qq9vQSFE7yLF6UA+pQfx9uK0lMLr7aLG
e74PlTPcL+JFKh6/ULG/EMvfSkoxOXlq4yDalz6zIQgyTZWb4IZenHEDzBbTS/akzGz/Of+1HXAS
Mh1n01f6/tifeTqL4OoArvA36UbWA9u4QziI6frJ5JSdkwurEqr8XWWcE2E3+XP7T6HKUhahU1PH
Ld2h3W8dm0G7T1o4nRtwp1T1Oe66hvP5wv2ujukjIF2TPgtSXo2kZUIKBf4H62fCj4Md2eG4xIve
NxbD6PPlQFNX2A86h/F4EyPy73tEfcCz7hrRfLVfyFItk+vkTRY511PQVKiWtil3AjexVtYRUBnx
cuZxGnqHDAjJf8Hzh75Gv5l5ggdWzBdZmpvNbGN3ond/z6oz99tNYPbbEIW+wi2TGm+6Rxjbe/Gs
4D5N5V6sgk+Aal8t9+145B01IWoK45xQIVlJo0BOhbJPvUWWpYKGtdfHYmBfifmO85HY0h9s3fDo
M/qRtUdjLEQRL1xdcY0dcipgFx4mtwhP6mOdgqA9dlVBgWCD3/osOkjUJqV577XBcarqGuyIG1y4
w5VM+ImR3CRfJJ6pHS23wjRPfh24EdLxrBpILbzRUdR51Y13qLaFJXxkSnviqhcEA/86+ts8jZMp
6nbqxNd1GamQWDO9yl147314v+OzQX1iT7g/S/s1JiHvXaQUJ5zzsZ2d0D1g+6yeEf+c08fJ9yCj
iRFy+5W4Z+REUBe2DHHSgxXtJRQYYgchJ7eW94E5b+EuLQnmz8HUdQ2RepXIzYD+fp3Rhp43jCEK
G9ryUHBSsyt1hin1Y7VQunGmR41peWaEA+Zy2yN/q9+jVGDIe4o9FAZot5ug5UeWJIcjMXhvt0CC
4dpdoCOlydO6kRPHU2Dfhn9iV80UdlMF+55s94fCSQdf8Rj6FpCBbVfQcx9yOwX98Z2spKM71se5
WHP1/HoORvM34SysNHZcw0RhJI+qbN0wU3c6pD9dybYKY29RBv43M5sM/H4f8iOTI1PEwOnzKPLR
3vKKw8ExYjJI8Ali7fw3B9kd33bqOS5SYSiLwTa0paPDxUexswS/qWkmdpOfxH4l5sTdCPGWGCZo
aQqq93VismYg/aw220ROS4puwW3AA4nOkAFMjfmLBFr9Il4RKidEewH7GmaFWlrsK20rTlAewZaP
7nclEtSBR15jXTzPGhtkrDUNkKYMAmxlKx6tu5zBFNjsaGvZJIQQDRPu7viP/TW00rX5N7ub7CYr
beJwdhgvwBVCCYzAmwGpcGZ5D4DxSIp2aVrIdkqPWengvzPcuLcZsa5F+YiW0EascoSyDOUIsmk2
QyiZKzEVZU2tYxO4KAc3jUv2V06C/PbK3NRQpnzMYCDtkWVMVxhj+aDlaicL3qKnFk/NqzwpvgE8
KPnfAXPa8mScUZNq7xBPs34OyW3KTUvgro1MHrpsfSG7CNefsnO3usw55ca3i6oHBOeb11+8ohlY
2O+u+RwG5o+4ADTpEJDm2+ESRrJmGSKjmCUm0ny+a0Jlj4jHoiVlabKUdYfsmuvjGFP+QjzPyGV+
893zkP20/e/4z3qzrj3vc/B7HoLbc1NLG8/AdXqQKGtrkVYg3Bs13v9ehLqAsG0esNDWKy7YfO5K
7rAGjn/+wao53gdfCyrdwy0MFZgZHQgAqrlUOc5jUhsdrrHF1tEWE+ADXvHwgLe3hxEGXz3m6aOo
MUDLHqaIO7R0Gr5GGE1NxZ+SCsOLZ4WvhYwJI9cu9zWell3RRChkbMYRn4hx8Ujh6GZ4KCrbw8f2
xKnGN3lkIpoDYycWU2+97zRpl53iiZJU70dYjtgJa1FuSEkzLERNOYWg8qudgrqyoWsxZ9map/SS
8BXJ0J36YDF+CI0qot+9xKWRz6vtVctc1tGaIyfl1/fI/YpWxQPm0y6RWRm5manXbHYag4LjaFzO
KjUb5sAByBq94qkR7e9+lKIenqOL2/jM2S45dJ43CJ127ii+WtAsVM//TnUY+dbG+/Iefv1Qdej1
DlQSeOi3vu8ouDP3Ksydca5l9Of8N0iYcKia7nq0llltOPLUxn1XDDb50wA5kSoXJGwjb+j4qHBT
9fGXFLCLdud74BLnMnl3Y1b6ykMY9RloWlD9E5PNAyeQL9wCB/+NYHX2AlpAwdF0M0ITTWHTNaq+
7dXo2MNqmpRbg9dQ/VVzNheK3D7CZa7DzXU1hei0Mqn2kqcfBR2v5RE3T4RGsgqN90YHJBSvR8ik
QAz/KPI+OYgSH9H6JmcQd4daaQYDUCP+1c4Uo6dBW4v4kudojlaEBHEts3hCaDJ/WIn9z5AeoDQT
KgjWvY6/lglMrZq6xGWTzw1ZYBqeB+91YJLBbzW/hv5IoFFc6fAS6w8TsJuyAAFT5Gq7csLF2JB0
NrNtXp+vwALYoIhJ1Z+MA3Rt0Fgxo5llncR2CxcQKJlVSQ/6xLd4+4AehP0Nbg22DXbHOJnSADSg
tyoH1rDDoW6ibDnnADTZNBsvtA6NY2Ah30MLombh4NXioGBjbUpob4e69DZt5su3xnW53oyNcXEA
rmffa9vg+2C1hPkvOttZDATuFs7svzrChrKfT4zsUR6FDPmfaC+Az6dVmOGMV/ZqXsOZhnW6LopE
Mcy9xdu61drgDJxN3lcSHZhsZ8zFaE66sHO1KDw0mZNG9UTfQE2j9V3EvumtDMOKln1yHRrwVyAR
y59BNa7Pp+4NdBskLeO4lgG/8yjq+BjyYSWQfAiRhes28rEZd2LaekL5c2ETiQfIZgZYVtSrW2Wr
xuAk4m6L7jBZ7PvQVecURpomgrPvPq3NGTt3B6h+Ef4LIJ2mXvXOmyOw8va1f0jUhpYLgTclFVap
xo5JqJNmRYkMM3BpkTK2h9ylicFT1ZET8POtlYgsTuoWfO84yWjk3rzyxavivE4xHLqYvJqSvczO
xzob590hKSQ8MlQ4XhX7Jrd99C1n/RHUV/SIhYt66JrLzk/SZ1+L7mqTJSjrWOryJs8pAzDnkm68
jBI1Z9odm0Ucx1SQtmgPqs0o9Jax81p6SJcJYQMzAvv3EQ4KcDTSuhvdwqcYRNyy00MF3bjJ8c2Z
VetbJqI0SxiBkwXTtg72CmC1mgfagr8PoDbFXwj7xCHVbu03iCqz1e9cvffpmDPtaUXR2yoGPSFm
oqAVUlTCmW0Bu0FAKiqW2c3cIH5+0u48AWfYldRblor93GMCuz0Pq8p05Bd1kjWi8rLqRXnnnVuU
E89mbSyJx76qjfBY3Yftm5r4b9D/2tpRymMsNLidPpx0tqi7b39hzawP+a1U+U+MvYsXdRGAyzZL
t024Jn/0dd1lvpzKMfxhawtYVv8cysLGAMAv2k9Tg4Y95VTluBVg67zY/WQFXeHJMOr6khCJIbCt
vCKdKslDLTC7va85B37gad0BW2nKk2125hE3GGuw0rW+zmpayiSVHl+HU/0k1YH2W7Na5lpXEF2r
HlFZygFLArDdZ5DnVfrEMzYINgnSay81hfdXhGhIjfKmqAqU+0au/ghnLeLXgXU9nQlnsLGmv1aO
IBPe8gZ0lq05IIYOkHmIajha2zTIfs+cQOOdnBt1c7eQKka1KSZql0WN4d3MijPdks5u5eMX1EfY
gsU/DS18W+ZVSu04LJpds38hWXRZgLYx6s0WD9fk4KXpJvW7z8gSA+W/VO28Y5Q45yJziJraUHN4
6pBCWQNRTZormxaBDG12jCH2bwC+mxgZ4TGaNls5JVttnNbQgkhuZSwXAPaUxqzgOfpSvzI81era
ORQm1u0nbzeTSCWf86tsfLye2qvLdn9DPWDWYc++wuHjFMIApSLk4mlJJa462UHk0gNukbH9MgUy
WjELfFq+60pxo89RXbDZ2Ds/MMrQB1WyCmLyAdG7IklQyZBMPdSvmUan50bPWjAdZ+ZTHgC5xC1Q
QcL1k/I2c13aG2M++0WvO0nnnJiHHLaW7PFPcHWUhdCZPXQUKeu+52b/L/QAfDgKHAWhLtPPWjgT
idM7TejUr/eIe4RDW3+iWixjybFMNJj1srAV4yeRJe2Chq3ohX8bd6Sv0vzAcIl58iDbyYgNPLRL
Es4JMxQOSInPBH7Ykbo+SnnjbqEnDLG90+J8nuh60dGZ7YBwqhRkW+1Q2fqx91n9OkFbWmYASxYA
B6PB8OtTKP/5n5qQQZR0gtzy/0doPkqoscP6IThSRKiRA5PGnNVkCahKuU5bRELpwPr9BSsYg74R
iW0wMe47seoqsOCnSKCKZxG9bJ5RLSddFA5jZ/cvSDB1iPwFPKhOfFjIz5F3mgCeJfC/UlLyKxyu
OylHZv9gsvzcK/OIABJ0JQEvHsoyVgWurWlWA0E46lRzOLXlDVKD/2l4m/sA+aF9Td7LCW3JGZY8
Jqm9PKKjeTV6zQU+O/cQACdREzdnet014JSsuV9E7FXLoKn4IDXu1N60kJ0LCSnEFhiQxj6rTrml
Z17cewuVGkW7TwDzNKegpRzr6AEy9MQRj9Aj4ck+iZ27NGt6VCXsE+HDJCcJWdY6XyFJBSi7HEqd
B6UTEyaMij2KVUyMIn18rJMA/6dHcxuC3iyHEFX3Kqfx3T83uAxL+wYNBw+lkZ2A0EjIRjg4TLb7
ORhPgJaN5SC1d7m9GQOaY+ki0oA63mc1kMm+1QGDYRnE8im6z5AW122OwqZ0B04SWbPIqJtYis2a
vjTUqT4NaNv2FxlInuhtpSlmeEpYeEF7ymz6sndwDST6nyvRlTS1gz/yTHjdzoJHWlF3yAhaLrC1
j2qbaqJOkDbYXCNRKmdpyDH33amVxxEO1bZvfwhtwQ+pFHJcyUGQs94iVsXy060T2uOhFyRJ8Fes
O0dn3dj/uvs/8N4l704VKtUVBxQNxYTnCNjAzh5qexb2DRk7+miZTUKfwYteiVgxpWaA5eLtIvh0
p6myuUD44X0FJGox456ZSITlzK8Iz1Jr5PLaOQZfoMDtvZRbNTPEeokhQK763/Gyxvqa+/Fas7iT
P02Px48DmdF70tEOg+L3TP0rS92Pt8Awgak7eTgzW5HPET02TSPnUYhRS+XiG5v1Rcqj+aNmH5I7
Ecf3A/lpy32cjlW2aXkUK5NFI4KmSMyiUveaQWeIgSNfxyBVko6ntZtJvIGBPLmApSNjK/XI/jNl
YtL0Kg4HZnB41uHajN63dV23EnvAw3RzUsb4z2VqiHlQm+AOCYJ8X4gSSLxHxn4rGXRlUFOuntQn
fUIOqKlvNK2xKqZmmlr/FrZqbqd47fn0evS3A1cOEumkBNU3ryY5SoXEzwb5T1D3qJGt1LYhzCuj
MBT6onV5lKMGGnk6pSkvP090tJ2cLGp2p8OjeAdcUuFy+DcrfZDRu4qLKykbWL23eu5ajK8IsYE4
C0AKd9HF/70TYw1iRgBBK2NK6cgO8bxXGq+6j74/pJOCIr8kMdIuI/ArqMDptHyctIIRCrlFW/Vp
KOAi/RvA9vVYblZj/iFyArQUWvmdFBkjS5E/eJN1jeso0IxsHZOeifdl/HeTCLCqqxxgeFI7JWxN
7EMQdLnlOX2K8N4ZvqEwCrm4FYuPeehMrKrhKQNPuQJKer3lYWyq4GNfavYymcEcuJnpe0OB3lNT
3T8GEBHPMBfjAROdOsEbi/X7WUlW3ReDyI4Mxq/M16OsnyXAXOUEHm0OdFSM1NckUJBoaQJQ3C76
f4PyU6olg4XeBfiTztmpyT9DzIgrLeZveeaszUvJr/vWmekW/120U80LJ1Xt7T/gn0fVW9Hm+09x
hZAm6T5SdOwpsbBw9+h5r5E8Dwd1X2fBigEiFG/dwXMI9iqTfvL8LWVp0YVEHkxK4gFeoJmYcbfk
qha7ZcZh3Wqj0DL0/Vw+t61mWJiSOaLXDxrSYV1t76fueYjyRIhXF95wT29ip8xGwtRXiZmOWaqo
wWaWH63K27H3Nke4b+mTM2Hfor7Lla6BhQhl+zn1HUStbNs8CqlI3xRicFOJ6e60Y2W2VJkyIqwZ
vDRGA9S7gWw8eV4gVioA/AZm1a4x/X3tBvClo33Vw8M1m6o5uxu6ArmrUqNARrVivml6TL8F96E8
QWMaXOUO6b6af1Vx18zGnkuzbwmuhx+2vMMRIRdfIieJZRfgMUltU0tKfHqfY5RLBIDNwmjBIl2V
xFF9BKkUdoBjDXQWj4+URB1Y3ehClcyNTAIxjHuSdBELbqapPRYRcV/i2jyxO3YyhXGDsLwie+jv
YGPXeT+tjFCZa/6aHhzvAvYPElTW3V+a888dLOTrarToGj95CptG+o2lydSfLyvVcrU9jMSOwnOw
h88KJZPbMLySOtBo9Asj0Yya3a7aXcRJ70EsweYJYVQLAWuKdKzJOVMvTia2mHg4NI+uQzjsHeku
3LmWoovVgTcJHXiokjmSSgbwdOVCZmOVCcM3O2PIX8o1BViaYP8v6zRL5mRP9QqwgE6svxcp56lW
/I8SYq45d14nzQcxYgmPFgsiC131EOL9LH2CESNORWgw1oFstp/FuFUz2kNcdcV6mBdF4JtzwsqE
0ejavt6Q97pF58mr6Db1rHu6IQrR7f3PwTKNnapHtF96K4BiSm36zr+jjyRFyV++tqN93DvCOJj/
jiFxTdCZHCVviRQxhPm3zgY9uRmyA2LOyladb5oMwubEpu5TC2iBPO45UVTu8ckWp0B+NAxH/vmS
PCVkWQddgXFGy2awWWrPRfZj0UVDeBFsisRkF9bp7Tpqr9GGcMYWlRpk7hV7AZZdfXfsZXcBpf7o
mHrs45fHg+jQEDRFrmOJwxtwM/kHf3snUbRfeIXvvzRA6Z+9VUWTLZL1FQ5M/fcTWllv+gBZLr2R
qe4QG2HC9VbE4sW5jBVP1PrYgjhwtZxht9H4SD+QMsPGW3tasJqPDCY0f6Icbvwc9i6AFwVElx5R
87DE7g2YPmTuacdySz8KwXfZe9SLwNUOgv1S2D2fLs7hhwwyAoc9wroQZzWgxZQ3ekRYykEU4Kki
owUttE/AypKMrDSLbW/fS/upmkXlcVpSIh1xYmiZL3Lpp3EqzVXYI+dvmO9EEV9FEjsAWWBe0Tbh
yX9cCZI9TlGxZefZcHliBfwmYJJUCRiNXHm47UaEiCLQFXCQtuDfFGWKQgbZpMeqVlE5qUaTljP0
fnALN7I3mvGtfDAAdFwnFhmuCjoIN855BDwJg0zJ773XoAOa52dlfTWUtlsQ2X1avivGvAksG/4q
yBCIA+93sgIQYHIXxPZqieMP2QZWLuEOdvJb+YWtjB7YA79Ecj9tNHZ9xPeNOZx5X86TNvWXs6l/
oQ2LW3rzPLRV/5Nc95Nby3iq33x092XUP5QVGwtIKquagJCFYDPlFunwrHvft39NqRvbZ62aQHPX
5LWUnkffsTeNKEsb0/GRo3BxzB2Ps4xlM0+PgdNm0FgSiOCHkMadOK185UfH0v7Rc9ROLWiJPM8I
41yYY4l9Q4G+3qA2MfdZ8BcVZy1J1f3DFNnDJByG3WAcUET/aBTVNPIAdlrQPWzHKjt74ZQ0vWLB
i9N2r6hMOp37e/TnWwFVQ2CXBRzHSZ4/Utfb0IhkBjzWzRCEPjJl2esktPZfFElnT2m2Tp6XizQe
GXxqE61rh2HtYlpOghI3NihVLvJpYvFlDv7OmgpdDCSa6nI73Oq6DaQHArIlvFIUc332kLOiSQVm
XQ0oeuGfla19GC/+XUbwolygNgq5VvuJmHNSPn5Xe+zfpc6j4XUCyZpAaR25Ltp9GGSwByfND6RD
a1VIrAfSbPCZcDPbsv9e81+r5OKOBq7mUfylLwf31vQ2OPFfWw7Vv3PAJ7EgbLtktPzIUKEM7kXH
R1Ry1AsxXFeeJBh2lQvTcqcuLQDKKxYL0HvYzXujWkXir1gR+0fX3sf//Oy1yQcCV565JqbluHBz
IHlGV5Ia7klc8/5/VUleFdEE14RJelBqcQArMMInAaU2sjz6ScDn48xuFiblnNQPjlFGiTFFYPae
Jx+LdmLi5/6jJWzDzewCI5JJyZZ3C8ZmdNMabOMgIVnYP7EaujXIBIwqsZEh74EKJTmhQRJf0jUS
1ah3StWCX1g97tcLrVyhN4HoCPKrLPXyBBtPdlcbgjRoqpskqFFXKezr71/i1kLBgekZ9OvW8p8v
5kEjEhiIKoMgm/Yp+9YAHegxhRIe7pjntpdWJ4O4FQQF4S3WYPSW1LxLckAE2oawVhZKnE4ZG5sH
ZxAJLiOfPoiglYYPI9Rh34/BDf5drt2IxqjWf6Rd/6sr+n4EbBdkzaxxOy9mVEGjUmK6HVfkb/cl
1BJUvIP4gKtJRq7mqC46qFXwM6fYeFvxdQ7RqdzS59RVC0GWGFOCYjLrAGinqCXmMz0Rab9nAZkk
pVlcjmOA1PpFJtTyoSpxEJC+l6+Cchi15jYd/PUlcv1WxwdNhFlR972jS2mpuAagQSXCCCrQWyJw
vzZYTTRp0KiRqAhdESPysnaNIbCCzw7P+61cOni0FX61vGVOXGczPgLjrjzkRMh5mXL9SbQL8iwJ
SSwkIi5PWS40xCcPh4XjwyIQwusVp0ewTTLu7GHHlZemrO4adGlkXGAthyoGg7B1DPg4G7670h+m
NzNRWHS5Mttdx5MwMzjnW0+wOBPgwDrd1aptEtifcBTWOHllLN4Qnb5ew6v6jbbpJy8A0SdkHayD
1qMlggPGB1ZDo/y3dGiy6vaG6PZy3ng07BwDyaXGiDWCzFXWafRIU0w8QiurTUNIyUIRu6+mEhmr
oeJTeQy8Tdb3gBhZF0R7CmTESzxx4WGStjIUyvh9LQtB349G1q/QDnTbYvMD2aOJiN/SYtHexoXB
Da0eu3STzrpnPmCiDMe11tFi8bdsfmiAJg/9SDGIVzozojdegm3yMw6Y9tK6je6sedXP1AI//bef
a/cc2ynHrdzKwqii4zPX45PgD+luERmB5KwgMC07dad/PlM/AtglYwSJWCt4+oGaZlXUgtnS6vEF
3sevyOCdM0pfoBdJeci4PK9xYy5nQpyeHJDt4m7cKFCO2L4xGERd4L5kM50Kc6i2Be7qcxaMHa6b
0VWReqZJrDls08N5sTxGiFbi1YlCJiF3k/3OcIqjiBnryTU7ROaOm54fkKJ0DkpGNUuxfFouOVUb
NNiVU0T5N9azmRf00LtC9d1qjZf5NdN05oziXNDOQOcc7uxiLIhNiy93O3+y+y0nUOFSIXD0Xi84
vagWRGP1DUs0Hh4CeVb+05dmbrbPE7KU2o1eEC2Q6SDDGSfHeD2SsiaMxR+v3yRTWrTwgVMLT7rP
kDuSM6rBNNAfBmojjhiI/jnP5jUXWBBNZAgamdX+qr9sxPxOKwsPc6job8Achb4CgePGqOo54Ipd
/POAY1YDOs4m/tkg9XtJ3vt3+73wukRIkHXcqoFJ0BcS85oH5RUV67e+OXt4Sg1PD7RiNKhDUcSS
JNbSjxCMs3Z8HTIpr+7Kom7iGTnigH6ncyg0SjNLFCesUHb6LJwMRRMiJmlMGcrqj6GJaIC8i5N8
qZ/4EANRPwJLyKYli/xpmkp7DxuiSWphZY32btvx5+F1X7UyxeoJ/Xn0CTSPkDHotzOB2SETg0dm
GiSpTq4hAEGoG7oMHiOmFDJW5IEtGeWypRuJZMH/KiCTwdfZfvGxAzZ8i7EQrVY+y/R08loaJKvF
wi0DlNpxIGZntoWgd3N5keuBdzOVWObfuZDRAPzLZJ8d3CrN/+dnsquWCQCdS70DQMn0SMsrMlnE
ovLPlEYuKAfxxqyDKGGo3R6LqtSdRry6wA71R+8jXwRRkJqEf7cgheWMH+JeuwlW74ZuXSvB6fxN
cFfuauKKwwBeN3Hik69UjEnKgVGw63nDH21+/A7nF4tRek4pfIfuSvuJRWtgs+Kode7OKevQbPU3
T6ZBbVOgFTPe88Kj3hZXUlyMVClYkyomqWBzbAXCc/kZJ0QP+xXmkuCcokHasv+zByI3Qgi7/j0b
Zd5n6IINn/xf7NtLhxLwStL+mFCX4bnmfyoi8Lrp5tvXWn9lyD90aLMRt64q7Ydk+2pVuV+Gulae
LFMIsg9m0tyfVKj0RHVjJ5dOA93RqQDQEvkl2H99/G7ejTinI+K2OmuNUMlqLr+c/0EpwQl/ir9N
uSwOLZnjmw9Aw+USM8HbuqxLxk6YSpubfYZCQU/ZDYFmgJtSLzkhEYkJ6y7RLbAocnEbpOut13Ev
DUFUf/HsovPKoKkGqGkVNi2+2crS8oLahVfXBi7pmFd9XCQKYUNl304j395t/fAS7ovs9kvej3TE
cd82vBDKDVXIvxxGFosDtnDR2QD8tugncsiWf0og09Cl5lPzfli/o2wZPPY6HSGuUelVjGMVHKkV
42snkpnGtJGMCs0GzMCLEcr0H6L3i3ZdL3y3GPxQWsvlq37x8JmZ5D7GgcnQiLHYOVOVTZU0eu4M
cr5edB5sRk2f2Xok48YseXf727V0J9xx8TqaGTCBG0PGZoQw+FpySF0KcrkuH8b1Cpxtol7XwsrN
LMztblOcWxofs50sqpY7hx/H3GsJvL+c4u7Zz8TJbsM4uyjOivefNYf+FdJRvfpVipq66QtIH1kc
M1UvPLpimZKKGjMyttYYVnvajP3lRa6SOfxjFNJdeTsVL66QDpzIxO4JqjyEfq6wP76zJxVkCUOQ
Cocnba0heUhu0ZQ5CkK40XjuuLctsezMq6CcFVky5NDxSm3eO0FI4tE2GjvPVl2eCKcE6wwZA8rv
no5DUyYjEMZnhm8/0iAY4+QQs39q3Hgf5NO62luvmg8dwHtF4QNAMf9UYDe3JP6v0GMFr5nkG398
ZGn0By/EPOwMxDQURR6Utj5FOyq/dGIox6FaRlxEsR1cs/k1YnFGwiRZiCoAD/tg/btiapOb3pXP
UuTqJhYamBmVqeqDTKA0ZWVEm8rDZqc4/xYRu0jwgCVrav0bAaFHVpKqZUldZFs3xmAfpek0dIvo
9TCr8hSHTWYyB6i1Efw64+RXIQCIjyB8FD11JqjBZWyEQhLKcDWBpm18dJFMZLpKP8f/YH1n3tzP
FM863Zl743aMs+EYzXTBFJKjn8nj6TvXvq6DoJX5qntePQ1JVc96/EmibCIKzDXqlJrcQO3X7Ko9
iM0tjHQ7eaBmg2ZEcqi+XtjCUnsWyc6JbfgDKZcDcb7O64Be14GCsku/KnI570Qf7Q40pZBK4spE
B7KMfiBBzB4SuovyCu5uDzp80UuW39n8XqZYd0O5L2NMfA4cRl0H7OWIorH6puwiVdHHvjua+EjJ
cPHgovBQpKcrvMXwAlavpCyMIzAvZviGY6VMGVtCo+B6gNHwIZ4OEQGWouiiNyi+i3u8ZWjxZXpv
BZgml0/rPtMtYBVzPrG98NfX2DnN2h6wyc9S2BJqqZczjOcVlTBC+u+d+J7q1jvcxHdHrnhqDJZN
vj17D2yW1gJ/l+xW0q5vLJc4GgHDSM8yGsMuisKFOAklQXrpfAZ04LsbmPAZuBRnFq/q0ham1yFd
EfjXtWIPp61VLlWd7NhMgty+ldp3u1/EgaHpH6Q4K1I3PGIdzvWxQP6E+gAprJGGsmFL7hXp8wY4
BM2pHHQlVBCh3Dsl6JaOHGQeUg3eTws10Azo8s9z5ZGW7eYV3BNCnEhpDmFkn2iox03XZwu4Gpv+
2I5aFYzOoa5GrPvLkmb+XxECi13SHdKnNVt6oe/LeTz0rHbfemiP4oKh3NrBihqzArn54QU1AMhS
D/Q14xVUZxsObZmnuVIlWLcInbRbiJOxJ6QNdpFEdQjAV1uWa+cIZb/YKW8a55lrV+8QMSXpOGa6
aaTpZF62zj37hloD9Vbd3R6iqtLNUO2yRHEkq98BKIrFq8mHTd/K+HNK7s9BsYL/vRF4Yns85EtP
OyBB50qyM5XILCtSL/0quWHvmoBYC2iCvURbCr5wGrTQVUe13vHBRG++kRCrZMbVMo7j7CLwwzEB
GQAGzYDUM+azLdb5OwtW3Oq8IH5RRer01ADV6kSucQk7tsvwUAGhCZuoKDLQ0qJ//4QUrDmZiWRm
OUi5ojlEepk5YqirMOKGyzEa1ExeCCuC/QbsCnT6lL/1xtBtAOxiSbh0BJueusQ3CQKFDce3V7y6
ImrH6EURkNC2QqdrvXwXzX20BLZ4HGqppkCihE0nIXta4Ivrjo5oNu7WE2habSG2GjED80CKYqZI
vf0fxgyyGqYX4SXkzohRJd8gGn9oceuqew0Mf+vQC8v3EiHMNzc0rPr19Z5zN6ceig9JVus20QFv
UfWYOEMzsyBxAvf+SacLSWY0B6buS1QUHk8XMBEcXUMmMac4IlrJVOCmuH0f48faxn5M2LjEChM9
Jh6pgA/ErrQyh9nc/rWtCbP1JOV0zKLPvpP8QkOFi3zVepPP5gGsx4To6EaMcqpk2yArqCVz6Uhr
QxbzfZU56s++cyF2Nw8t2jMaqyJXx3DwTsUEex/x1APgZFTT9Ad8lm1GCaZa6CRszltd5KDZVhCA
0iPKrEU4+4ouSMCX7MK869d7xs7sD6aTtZ9e/Ty19lEUAi59slCdeOwsdGZusCLEFBBK0EnPZaFp
kV3P06orX9WjJHSYYYCsPMzBkdZgILIUtrl/xY7bG1SP77evC4z19qIwq5Y8kmGq+RgubqHYDtX7
fP8Jx1Gc9VAtNVIBqDECevdZy5UtM/eScFvQpVZbt3UuGKvBYoA6BRmOQ68OXWI2VE2MZgy2Q/xb
MpL5MBa+ZoL6DpRiYJflLVg1h//7xa/BhshqUYyv6sA3YYQmtxyIxrQ0VybaXYxv8mAsO5OKpZ9i
K1M9rYADAQSb/ZhOgiI3gH0WuCZe0vVSUAkQCmzPEx1RmX+34nTOotXxP/2Ll6X4SgSlIVqfXGOh
Ih4x/3gQkk+Zd0h1A3S4oUzzTvoN6M7LtQy7KxmcepJEkM8yN60zjuqYbuOv/xLocop6BDw/9/0J
Dd06/XOBATQjbnFbxNjSjy6WpgH9ZS+qKRMtTp+d2IWQ6jqcRJB4chgh7mY5EhlF76iG7DLQ1JCQ
l9oqCSVjVZHkAfrPzDt14RSL++kFBt/fat4WKeH+ocncCibbrwPwHiT7TB/2rlXkFdwB+VzP2WKV
JuuDm37XyYjhuBIKggdHwWaZNpRfjUnq2NEmm1Cc16D6L7vk8xaLZZ/40lIGh/aJrsPXdiO6iZ+e
sGS/wwijJoTUrbyKSK4Mz5u+MAzoDqsEYfQiMAkaDc/7sMtmXmnp+k99YwqSjTn0H16n89bIKfu0
+JTGtTK6aTNXPIk+f7gKnrUpJXLJDPxhqZCFf+1lqQQl+3w0atxr2MVVljsDuHvQE8wXaKmD/xy0
CJNueCqVjxRi1XvHYvoQPj1BXsLPu+6pwoNPYuSQmcKd8X4VHu8WAOFCwLzordTu4YnsqJRFKeSU
pmM5Y+IRRh9A5HDRtVeIQDCdkfrJQVlX1neol0zba0syUK+j6ub4aozHGxsjI3bYmurfEpTvzWgY
DXuf1Qy6uoYhzcB6UZZA+LmggyOg749QnqxGWUBehkfChnuakp4jCrVoAoCWMAsGeR2YkKWelKfl
QDd1Baxsk3AJkILgAC5PsSHAmjdhFmsXptJFB3mNARE6RkYy/dTsPX6ELGwpjXhbY33x4U2trGT0
1lMu85sc1x6Wan2sCwTv36vUNUEipUyzoStppRfL3KUp9Pl9AMZSBaEiqPzsqlbagGI6Do9V82gO
ISnqBUhejZ8irPlaoLr8nbxDm+UMuRxCHZ0MKdHsIAkM+msLqBlfTW7kLRKDMoG2x4wzCOhAQqq5
rCJ2aRVqjRhAcBlHCt/HynYE4vcoq2bRTGxqVeLUx9TNP+4yUZanwRjqHkjkYz7SJR27JazInU0U
kkmCsPaSCzSlnSBYlhIaMIc7HHXaZL6mREtOjY0ziIKkvqBlTFhhI3fbA0Vo1Cv4xmuMp/ITB2kw
y9bp/T274JsxCs3nPSR/BKQeBQWZFnOso8BAkfjC3nxRFZ0OHoGj7qFpLNKnHqOUMSX76V9Iu29q
iU9VblUKcoeqyEDwjQ3KYMA3molMt6Y0/EFRmEBrhY5EM9n1am7s8CHsn8P6fx/0DMTLQXl4jgnD
KycnyhoI/RHKV1IK4hm+hZ0S3gvcePW0EbD1mj7QT1gBeEPAlHukz+CKlGxgYGdn+u1cq02tb+Ih
0sa84xwr1xKE7jCuVO6gBrnEhBe/p/+eo0JyzlQGdjJiPp8e6Qe3QO3kVc1K+/0RiQfI9bQfPNfi
oK9e0ulftwZihUmTmGtVylb1DefG18OiWVUcTzSRN/tFGGjeHCSxsjWdmOu/0bFJR4P+vvs9AzU2
EhYVsA0hnQFeI3KP8oyCaigosBOGyday7rENlz9Y44lQ6cv4GdvWzWgnBlTrsFrpmQjWqWdEzpkS
83ehl5Qad9jEbR4f4b1nTtOzgVsmoX6CFPM8dNzKk9ZkFzDw5P/zhdnI5ud2iZgvsOkr0ID/UQpS
gg8ar97Fl3mU61NnirAu1qtwOsquRDlT4I6lGbV17SbPlThpfacNGtISH5hmrMWZ4Uoc65OyQ1Pp
TSLQSspStJeCDgRWiVYozhFq1s+g2DV2tBLv0ZswmrGrWVB7L0KcebEVxRrVZTPk81VXQdT5B1KF
//r236jW8RGyHTa2j2NVuSyCereG+Y2/vF9EXSjbRmGFnf2Tzo/5egFORqa44xLYNvkKqWlIZRKv
X2T+BFXfch3jxo3wLWN6QYRZDZHnjUyWzjmgesGYAqwtFtEOJpLH2ttmP4V1QwxGOadm/E5WxVKs
kNwV1CZgNOcOIF8nmTiLPDlG2P7vPs/N57is5501TCSwJga5y9sTWlJHqj8ZsTgzDPwlORZ2rtkA
9fHEzpsGM/T0aSEI+G7VQxdvxOqHy6W82amBm6nDadFL8PGRz1Qkb91U8adnT8RqPGjwQ2sG48YC
F5dLNc3ch6vJVvssnIwFc8HeVj7GObxPBNfb4laF28j8pDyR+7SkGbHuApYv9xlnihaj+64gr0if
wiFwh29F3PyEVBs/rMTuAQmrw1t8OpurFExQ34ut+rigWtRU4jZRgXHFDM59kJ5Sap7qfIzrnjxX
0ed9s/j/y6MLATnQ3d69ZRsflquYNT8rOKZzurquIFhuDncoVTKtMQSXIibnVYNlBDShzmUKqGyZ
/JY0ZPQxrc71VI783CFkmAZukvpkGgI4Baag1iJzBbbPvH4N+Ta5Rc0XnZj6h9l90HT+r1LmbH9X
twiBK4bgAroq1uVArtyOka0/+7zA8zyPe95Hpid1mvADhhPu6r8h9j9cBX7tx8FH57qKOJbvw761
o/JtXEtfZDbH2PC7VIH9rBaVHxg4WKpJy5zKptugKSW9pQsTzc0AlFRjGnyaLqGYptBdog7fFLR8
JCP870m7GwSd6Am2WhTU9BIPrZ9Cv0yND7mJ84j7tlrQF67UvI8Vm3AFCpreYpxiryMIZ31gvEvH
Ui+awpXClz3cJ4/GGB/k1lDpgFIQrJwohhEa+Cj9BiWQccKpLezXLfcACfk+oCuzy8iC94O7fM++
sjoa7NCwjsgAJfXb/orvj2tXzh8xBHbitLyh0HL8qeX06oQG8XLNI+DSHbhv6ZoqP3ay8WKXF7vG
pBaBj2MXHfgHztWjj5a8euipl4BZ3fDPQHpgMDi2SCIkbPq6NL4BQE1WvN7OiL2CZhGT83wcWPzJ
Etizb+E9mk1wKCuJD7ul3p2XSSdl4xX6IsdrGnNElm8FSmQiGA/R8ClHXd1Qa+816IekDhL7RAsF
6RbwfX7D1s+OGJFIM3OIuVr4elVw6s29GlGkLNWRyAQsDfBuSCHvJgJGPfXPovvHs2t1qrHvq5yW
cfuoDKkuWh8Gd/zNdmfhPJg6HwTl17ZEs/9rfvgSfjppGRVC2os0jHw9HbRCxwMSDIUTF1k2l4+V
06J2rOJBMyJmFln98+pgtJHgufT4IocSDKdfEYfdC122lytGpP53siAtJa90lF/m28GH9uRTwpvg
nidqeCakrmOEDqn2PE4ULAj+DncdPyMBQZyTGJhJ/C6tsR99e0+OlfS3Iv1oBAL8DYjsGonG3OgF
lGcgzRGFElaRKUh7bYAgfDeyh8QMfG5eBp9+PrD/S9LgJLWqK5F5sDC7HVez81GIQxBEQPgxr5hx
vAXYhppI0m5Dc+6O8a6RS+OnQzrt+dQPkM5Rl9lvbbBIAUhXkQCCEN5UJS7ifIt/3jWJ66uasrc/
KWbnl5BbiA50yhjOcnG/NxtO9G/Qy44tXS8mWViuAm4bt+8FSvflgks2OkEU9FQ+O6UJ9mycCOGa
NmNddSk3K6LGWB5NhwOxhw94erJV4cDt25fl7KoNgbgFB90nAl1iHMnFV3azC4eBp6dOAFTavOrg
XQR4FWF/XPZXoqeN2Pdf06wNVc5rL9SHOohIaPQTZVINZ6u522901bmLm6sXzgkInuD+d0xOm2d3
5tg1EVNHHr86/yNvYIrVtzF8EtMLd01yRErBlviaaT+K+sTgjCekaXYnP3710wwPkUPftQOotwCe
160Y4mMDyaVe1pfEdIcg9yyIEr1RaR48xxbXUJC+2zt9gzbfQU5+U461qpYQL7bvjsDd6rxSQMUV
5BgSe2OVv6//Gu6ULtFSGxBzFAs4b7MKWim7GbADRH/cQENakCwkSCMY1kGmXx90U5p4JS5B5lG7
S87rLZiOU2L0F+KQAmPlSaZNnu8pG4WA8RDGKyRzSBuPql+p1WagTkFG9A4wHqMLkNjIWy4g0XQM
CPM4LvsXOoVA/7lPN0fVnQ3b6iLmpuXrDFxfdyLMFYopzTvmLbCvHa2jBb0+jQw+EVBlmg8/5yx9
YWnO7K9zIsMi6jOpEJ4cUFkUhgs04xMoC7EoWGWNdjTYouP4WUi0lZ9wWmIeWCO5Yv6kwmrOPqXK
VRRzc3yfAkotJTKefLP8YRYKH7Cur4XOB27AwOvcH6A/2n6mH5q92hLuWKvZ81/3WLFcx14R5zs1
Lo+o0yAkdhpuCWJkZ+C1/z9L3RMZYwHmA7PsHnwOTLCG+josogxFMtF5TerQ0+DUWBagAVtKK5C1
Y3lsmvuxKta+s29wpoUnHlNIymCwXitsFgxGm0ZzM1jEa64kNX46eV+Jx5/KOngZ8KaKGn0Jqhtb
KB5ch65+btm9QAr5vBvxdr3hy3Nefbc/6Bvn94EelF0Vj5dUx3nKeeNT2v3j+dNBznD10n/iFUKB
mryK8TDsdygqugJJ+A5uIHsgDZ2Y/6joJUUVni0i3pEI5Vn8PnRTYImdbrc/5dvE8biYo9mWbQhd
GFnJttApvOu33L8PfYx471HEV0/Bvx7t9wnWf/UlDOV50NPS/BDJNmIOVGWEVhWSz6XnhOWjpPKn
2xcNlGAl9ru9hYbEhe1jfaqo49Fu/UgPf3LZApeaTeeyh83I7yEvmRjwx4YrMeSusUehAlACwWxH
BGAdSaj17RPXWD/SXVsubLNzyhayd1o6keRP/6fmioeBQD2mRl6hg7+EWRgrZq2L/QHoBsVAtZeo
NXIPBAL3qkbnkF+C5r6xY+xdn6Swe+tynaU6PvIervq1MEtEZrUDnqSivYmp0tl6I8BhMpfG6SUA
Tr+b13xr+ZJ4il+Bi43dqleHwLEZ2w2sJCTqjkzZm6O264BPrE8NYnwaIQXG5DD1A0Q9DvrumcBV
73fE4gioSgd6pngkm75IqgXE7/PWQ2v5bELO+ZrPGqZ8eFqrNSp8PbcIHsaTnSIseFGgkdve7CFJ
qYcemWWaW4vUm5+/sR2MSECwxdZpVoCBxaLwkBG1JVp6h8Go5aHVrypI5or4zb5hK6n6/khuaTCd
1bLlbCjZ+vs0lgYw5kr5/XAEzGKmr+tifuWgdMu5k4QgZepgudKGb1zjvAMdwdTAuazi7btqBkAR
b+0Oem7pluFs+HiooQuzjmXOVPERlOsjVbXCpIukQ/0JxUx3/S3vaZqOGdWhB7/ejMv4MlA8mcEk
LtLtlWUNWe0RbXWl4M/cH5I9hz34DDF7ag+AlLTtEO29OJaTT7MwimxICaWqCjAkvdbpxtzCz3Zj
wczWn2FKyxvdmoOjAz+0Owdpxi0LdbmFqGsg0eDzBK3putboCY+1PksKfu5aUH2VYC6xLf0FeL1v
6FwnzISmmZvZRMWx0mRnb40dH5mvzv6//0z226owa8l7LlJWbkpP/48+umnaV+AIb6DJcb1cp8Ur
no7qwAMJoJ+Uxa04nxWENNoBn97FXpZZfnG9YIJeSPkrINich5mZUWS3k2KI52R6WXdGekut3BlR
6Je/VQb6e65FCCRqOsGLoxquB6UIkefB6mouIYi7S7dmjgIPVi0RKvdrBZzxHmhZCJXRw/w/0RYe
Ug8JVMuqthZg1GKrnclQ+P9dRaj0JgWot80YbvHQa3CpzqKFuIGDQ7eeI3ZEBfUVMNAl9P8wwn8R
R181f6glhd3lFllX8Q3z545jwuqDfkG7npCY1MPen7XU5YsT6Vj66SUKQnuW1cNMMATYNf7iMOgI
cDnV+pxhR7VWtChfRa1ujcTxX3H2X3dxbWiKnsm0dRrGHqssfyPc6qiQkak3wL1PSJdY1xTtXoS0
yHbHlRbElg/vDietjD674ZY2w2onVQ6PIvacrZT7imiSuL1ujUtYpiaTWhw6NhD5ftUAVQ0c8shW
ySzi0ppXhghYg+LxjxEZ7kHGkxfukuEtlg6aZwBqDWwxut/5pAviqdylY4NPwLyXkoQhtuqrbny0
VHkSHf7yHaxi9nfLdVtFl4Vk0iOBYD2Jxv4tGCVVOAVQU4Yw5pDf7zIsd3pxpPl9+5c50UYU4Z2U
z6QuQiyFKn135u6cSMNgbi3HZ05NEx79kbZuJdTRsxoJI1lIi+/FrvDgmI3L2xfDbotGzBsGoCVc
HnDpQM9nns33Uku+u4JptkvdkaiADh7cKPDbzBEkKEfUVLL/HUcfvPtHbE+BDVSe+FzGb+cwU6Q5
yZxDyuesvRRBAg1ApPs9ToeSHEuCkKvSe5iE2p9mmv3kHqAMIRqU6bBWLIrggmub+mK8oZgqmceP
rc+EOwHK6XYdSL5TY9MNnx2nFQ2eGFQaqWT8e/+Gt5GiYDUJ3XLvzybuT401PZQAT3zMRcZ45LSU
cj8LDmW3Eo6aEGsKM9zEwGFVvq8mvU1rpKV5k/RP4XrNcVqlrcrl/CALTlLz8vcJN0Qs6KPwoiMq
LoXulYNOMxJWZAmWdBRGQGckMHIKrP7hKqmLR+D0Dk/zDiek1qqBLnw3s8TIoSf4hPnnSxk/FcGn
jwSQIEE2suNlseao43hdDkFPrZ0Oj2I1ZlsLz7j4RBBkPU/W2NMdQU/VnGd/SkDe05LOav5JrhT6
fwSpbii2fkItOB0ux/JwectFsPRnwvHh6fXqGs1fHjnhsDCGZ6RhvfKtciQJdN12F69LqPScG6Gi
kkmoHa61tl/nviY5BDeYJhoBWeb35spy/pFhqinpWT/JhKX2YLXGXDbz2eJUgYMOoRdCSYolBlUW
MAcj3Gm6OIP/EEHwCCkiPwlzFccXk3xcVx3ChjvlxaErcQrcuXWkYSUlGbR/IxIg1w261MoMeZU8
HcWvu0deUfzdUrsuT76JBkKf0TQkuqNc8eEfOmvgPnoxB5U1yOr3/EUvnoHupGUxaEKxOo5b+UEa
RxvRxNFRQYkUiT7tQFx/WJYWZVNlMT5pKW3a1TJPaSdZa+SSJgOnM38fUh7Yvf8VK/JL/JrvFbgw
TvpRp5yly+NIP9ajpp2LU1n/hJr/eCHfvvVnswugfhcq0l6dCLuOae4RtMJx3uYILvCawdqPubz8
Yt2TdmX7xWHeItEGub1Qcp0zYbHhuPOKPfbgyVDRtOLDpUz4tRCOvfd48PXFcbL8i3NUfXqFKPDU
5hl5QtYSs6Lk+s7DTNUBZFu1TBR9ReniHYnXsh+S4VgrrnYB4yin8Rnsu7F34FNTo0qf7woCfqQQ
AgBySaKrAoRaq7htAG5IBLLbcnVOSwE86VQbPDuH9pndzm4zlHw7yN9APJdcVzHgSmYYkKtMZYFC
0Xglm6ysYugZW00gqICAS5idT4eABu9u8XRQTkpmW3nIY3YOiS1b0562UOfPjodhXbY8PkCjzVNy
c609nfEJeSRmb8TzFg0JdVBbpoTKyRwKc0lJ7uttegwFuRUeOR5bsc8olkdHSiAEPrrsANNPxAbt
oZVSsgxK/M0FO0+5yYFWWPoZu7Szf/C9zxfeVJGGNB6Yh+iPerqPsGgOIwiyArrVfE8nkaUwjyJ8
7iIfWSG7phrA3gZqxXwpdGic8dwAZaiCEOHmV6njXImuRvFE4+lwpFOnUedmKfaM9fgPT5gFOhme
xSPCwyn8bRPsfiyHGyhpeDwck54Jd3hcaZ90Ll3l9c3SMchQ4ArwkobeR2erptyHeKiSnrRcg9d/
ixFdufOL2VdANWZF+HllFJxcoJeLVe8X5bypp02+ecgfxJzmWX75vCWbgbkH5C/YC1wVPHYXDeub
QXeIdhtxABkem+O2iJaM1SFtZasOWNfBtowGrXtnVz5TA/MTFRrktWhAM5+/YxMvOhIc9aoGhauE
xZLLfAFsi37XDXLqDpzUUhay6OqqJsnK/oBiJ0oxI+0W7ASjXlcJnBmoa5ZGIA9+O17ZqegBdYSQ
0EX2hPrZPeZUPJ4l/ePy2KPjyOzH6H87iZXY5gdpmwyPeQF+Fm7qjNmXL7hJxQJIKXBsNOk6eX6w
KNdyzPy9piwvqiEUSjjiTv+wMp7mbXlD5tRZk/39RRxsWT2+2t5SQ9xl1w4US5JdQ31IvI3HGJti
n+DmOgYNuZSC49Sl31xuTcDA3ymXjQcHjz+Jh6zsQ324/vkVV3jISEj1w2PV/AFcqgXluSzg91Ww
L0zTQV+87Nq4BqtP9xcsBwHY4pVF1ASZDnR+xp99yODvhSIC5oDRnwRxcZXeGQ5TdtavEpTN0QyK
NFM3z1xFh1oz9WeLAeHYq8k8TEkIkzinKL93qqG0pWFIP1nE/mBshhxVqcakjWNfGbqNwo+yKA3S
iYkBmQ1ekFkMmeSz5Yh1XyDyhF6pEPi0cT+6f5BZpA+iEdhCg3rhfG0sG0X2MZrk/gF6ZRrh2Yn+
QOUpqAed9VLbedt9pFV4rP+vVnfZBDdP9OlCOwbh+wFoQ5+UUPBpGnFJUmImDeMDcVTLEAWe10zp
8e+mgiHrGN+blqxsWBXC2WCCTc4eAFDKOQ3SZgL8pNtYqh7jPZVhVnLKicyvIPkZCIpiHtc+VlOu
YYLing5mG59l9VjT3KKGimw71RFGG635zZef213J7eDnDjzoamZBB/zweqebOpSGsnlfXJtnIv2Y
CNmoOdC6eexeU/UToMPEJi8vjXcLcpd6ldtMf6w25K1H6JXInjY1NBUa5kyNvev7edgG3l4Jc/Wa
Z2fvzKdKLvEK6beEKDLOubcSIQ8Q2SP2b0CHcQYAZWwk4L8NHHo95yGcZ4Pqa1Kvu/p/7LKfOSOf
Q3IZEXUX8PMYQEpFeVxZD25Hfe3hIe8CycMua4eHYYWk0Ua3O1HDrOos84xsFVZASKmF5rwLibfK
3yWlJlkPX7XQSvsZ/LoQsS2pmuflBbiIZDChOhXmlPZ0tLDGgDqlc111e+Kyi4b82GgFVd4a6Owz
xKJYkyOaL7gCL6XoKUuMfoXQB2pxh7BH/1u9mALTxqVzbdgEzu2OfjZsfmqVcYpcFRDEdaPQLaur
vNMDSx+s0hHiILo6V9SFwPghBp1pBVS7RXrVaKjE0I8Vb5usiFRLiAKu4k6Fa4+WZ1kzY7Oei732
R9wy6s5zZ0gFT3a7kMcfr0yQH8JLHf4pivyHt4g6luDGXAiE8GgG7cSX2+7cJKvegPqIZQSa5pOP
1H/vhfr2YQdjLkupEdnu09lXT0ZAm+HrG5VYUdbd++9vA5q+5cCpdaYQv2GhIl/M/+FkHCb0LLWl
g6XuD9K+4OY5Qz658twv8vphOMk1glnVxXbAmbeGyOBlcda/zeRtVp9Lze+8D1cLjT45hWFE495X
39oe+57odn183/7xolAwIfwrerXT5xt5Lp9wYOdN/6UqDWnrufJYggGYAlngoyV9yDVxNUwG7pn1
2kvyD5gc/dfN5gjBerAn+14Jb6nj81X29LYZ6S7ecP4B7EhpTxlKUX3nUUjCNUvd34uM0IjRZa6I
sJfzawgX5ekRSDT/SBTSuSkRVD/Tuhg9fhJR/HSUi7qOWcNWb6dAPm68mQotfjsxE94guH+aY2S7
u8WBNxs9M/rxGQDoYL/tr4K2gIzD1h5RdAz25yWXyHScguKS4zDjMCApYsWghfqASoXk/YNvu4Lc
LWICxZK31IYsDnLXCOMdMfjmAO1dSSoFHp4/wMTkxMJohUssIUlXTNM6BU4IGriOUESRUKDV4sVO
6kAucq85etgRPagCSigcAgP8n5e0UuaWTmuesyuggg7ZkDXvI9gvNLk67P1/6iX/HIGQwnpauH9C
cMGgMrbfBU0gvSjmCUzs6L8QFT6Q793qZIH1+3rAepghfQCV7dKcsSj7Q9Sya7xYjiJee8eCiEO0
ErPKwubvsonPRXUx+Va6yBRdhyDSySaBsZcjagqmEyFna166SdWd9MaT2ILMibPTM+nPO4vzoNcX
wggFOvXwpguglDyXBRwvX/SRZZKPnabbiUeGlnJ+3FpbnX5EeTntN4+SRWe2AMX5v6s7c89TVNch
iIrzGMNuPXLq5ZipLOLPf4nPCXisBgfJfBHChtuHABbT9/+npDcGlmF0PR0ho98QGCpu5m7cR73d
RT9xjg7dHiaFe9J4nEBc5mqPnfa8AhXPSvXC3X1ewnN8nLSSub92cJhsFnRlVPymWoZsuCObX2uw
Xh0aL8A9PQlvbTIuuNRavYOwlJeLJzCf2o65gkTK+hFuOrJ+gBC4VO+/96DQjMn6a2gs7XSLjXVe
AGHxKkSCJY/XIPhvGTe4TsMUHOKPSpOaOa3ejyg2UF7wiLHn1vScy2AmDFaRSQS1liGwfNHgXWmR
4nnExTrDKCiGtVc6/7gemQeo1xgmUR6hnSRqceCb1milago3oxyyy1hqE7Zb+J37UAnNq7nDeIna
B7yZS1bmFxgg3nmQlXzli51aoBoJ3h5nLd+VQIcGAnKa6NbALb0ddbKCnqbBwTkhLLG5kQtTlpRg
24kH20PV2sW87wtKHkvJL3frgamsPgTRZpGea+7P3m0LmxNgB7QdrPle77PCvBlAznqnFbwk+4rr
NMFHhKBFvUmHY/21DLBcRj5dvrEJ9eOloJ6wKmplZ87Kaaa51gm8dbCY6e54U/Yu0h4KF+cADZs5
ZjFSZBJMGgPaAnUd/9pLcgZf8e8LyyJ6FUxezm0r3SHYZimO/w+jBx1gaiV1sxGVIY619jPb5QHl
CuRcqUDHbPjn/MpKIPtZNU3VkzXiUoBSjLwY9It2usGRgCiBK99Tw7KJHNLKqEufKh+Qjax9bVfd
DC0XO9ruSuCrVsiHE/bz/z1vhy54lhnBjNwc9zJO/h33yBC4nQkK1l1X1QRPlwpGwto9MKqaywUu
AibWaYkuc/Y3k8QuJ4brCQEL+BNfdXltB0DyZaP0aNrPf2a3+SMYSmILij2Iw47yThPnq8rT9jnW
Dba4VAaH6Qk4NnZhWZ8A2Thm8fUL9s3/GBf493U+BgBWhI03KgXW7ZBFUIvbW7/hLBRYv1tjtDCz
9oxvxNP6BNOjMRy9+2q9tprNj6WvVjq6DWt/h/yP9yKQ54tH87ixm8FmYCQfL+4m/fNPvC1j7jHg
el6Fe2XkUmEqZGTV409GU5rAw9rz7BtRdTzjwVuvZLkXdnTKP/Ynek69wEcV9yGYxByjGLZ7RaMt
zEwE1bCJO+m3SrfUKz7HsfctfJu0DC27QmApC7STnwJBei7gxqWu7dk207Es2BCX0AM+AwcyOk8K
gMmypDHaODkb7ef7KB4VtUFwdQpZrh5YHmUV3PjovWUnF7zis4wn/55eZgltIAveRJNDZMi4mzYa
wzgWrtyEclcEgwFKVgR3dZprPTYf6O+HGWnm/eV8K7XombSsEDeQvTDJxguCAOQ5Jkb/EsYMbz1J
RP64hcFP/PhRzo252at8vYauMGdUqbxvxcueJwYc+OP7vaKYOpw1a8gL7O1KovY7Vof61VcUE6l2
k3d21yFUybt8HssxrmqdEXPp5//I5D3cH2gl3wMD0jyT2FvQsEr1Z00bJ0MEUmZ6fOF9Jgktu2Zw
BpMHEwvS6iehuGtSMF9JGo+H+usDz4+r9vhuw0k4SQQBZiRs4CZaEgCir41dQL8RR/IddbDh1Bi8
bQI+GsXT3BhuHcZYjm6p8GhOVaY1kQnnsuxs3xGhbxFIiLDThs0jYadTv/kMfL/w2qNyBcP8npFA
Qfg8AnyP3TRFR9CAbfznMKteGNjeyyXYxHRO04TketzoKiAxXTE6vgt0wpyAuezy48Crq8Quksbn
MHI1YutmlAYPsMGmVNdGaq8Xe2HlyprNjfY6Tze7BRUHU0XWEf7tOKSyIujBT8JpHd7goCdDENGU
Pj3LYGzbbcjG0bX8tGYN/yDXLxgdbzPCOs3hnlMRBRO27PT6sboIcQNEr0EDO0tWiyK7OGeCQBjT
fNgs08PUpHVe7HMU4eu7x64SuB15H73EeP7NayI7XmJCI/n6qDVzej70Ayd33ce3k84sJXc7ZEmQ
uuxHvSPsnXNE1kZL65v0b5OHQOxVrzd2puSV2LPiB3S20qFn7T62w933/mmaCYahSt2dj0j+jJZE
cH3ymeICaklb4XToZgncoZL1+2+lqH8BnZgeXSRLAiKWcwk3ibWyrRRMtwaLuzwc/K11ilBko6pq
7DcbaDNla7b4zMOH04KD+JAstyDFESLzphjiuzdf/FdOKLp/60kJkF35SPnNK5D3jkYheH6r5Cd2
2fKHs8xu5MvU82cXiOi95hPqxmrPUDHeyCjFw8TUCijdRKED+WwH/83W9ycr2E5vHnKt8x67py8E
yUdGHkmL881kyReX/nwSd6Y58048mZfo5vDlcO74AJbrjF6FFdanz7gxyrYpgizA9dsSwGPtoxsV
LQz8f8DWRyQn+4VVQt7PdB6j/is7R2eXnSbYSVKRsGyBw4t8a32Iiy01JK2JZ5JAijAPIMRM+xHi
DoPLoZsGVdguhlMeViAcQApaJvbvX/nhLwUk/UXjnNoO/ghRDt2C+ZxE9CKH818+SV5ygjIV4eGx
B79RRYCoJzkaKEaK+zuGKpiiDKC18XldsZuPSJ9Wq79CRqtNVNggjYBmQWk1cc8OWLccQkAs4BNE
OMXCKyBajm2Qzmf+lxW06xDhruZtugfaFgK/XdW+cDrUKpoi0X/pd+s9TYuHwpx9Z9o5kG0BpfzH
qOOyIxetrzCqgSSbp3hZ0rWDoTEoyFPZKDlfFx4ZCGcMA3WQbFYVFFLMUX2hGZ6cu4bZtEuOvTnz
WyhBDtfdewxW+7hf7yaPo3hpRI+AtGTK7yiQb/UkJuyyTPeYXjpsVBkPDDzhiHYPliD6lnZhasIK
j2qY/JK+wh4kOuXjE1l7sDp+l4lFDmqxA7L1+C71yPgjIuATapkJ9pchNt3RdC9u0UeRxNwQIQAY
DjFr2/25aBhX/+G1cBG7dGBAHfOhpwbmJd9SRtYFd2eofWRCtxn1JWszEjL735t0tFWD+o4LzvNC
oV3DZi7Po8o/kOYSFK/y0qpXtCAKiqKUqYoaLal+75Q1b/xySCpdRkwJAzxxuqKFkOx5N8wBfn7D
cOYtoCc1qzfdmye+v4tcaJT0tzDNEqgZ6ccViHN8ZTlh3K4eBkznUI4VGuPIFXj51p8FYqnP28My
Q9hrYhktMHvdvOzPWpmlSXn7jKtk/onFE+OxkyVOb53vnRha7yqdWRgnQWqFSZttR+IqM2wNGfiW
Po994ACKwsPORkUI4wnNPrfYfCSn2XtyyeO23VrNi9b+EmvM1Z79lHHfzz9Rc3LwPK5OiClwGMKW
7KqvGfKkjsCmT4ATdVWXsK532WaEZH6eGpTus1jf1RjyFj6oH9cEZswreL1g8Utxuv1ZyHxrzRby
i5QSrzKVVJJUC0llNJqTDmabjByJT2MqMHMGyrrKL8akjlGn5x2dM3NJozNF17yOMFGYn6/c+W7M
X0gKZ1OFkPy03IK1itPuDS6aLaVERX9MxRNyz0CYHHV+RFqvjE4R25cra9KXL/n/2uiIrrWUxE+4
8OGl3RFCcBwVu6IUAkWJXBDIBWiJNAtpfhT1Irq2Eb4NRg88cr9Q8ULb32bTW5IZph4G77zr+og2
Fy3UvWjpjJqUU7DfayCSxH2v/8y/eLvs4OjhdWBKRDdI8GhvvlxbN0Tm3tUWzU9W7HhLqlFDqA51
oPVrqqHcxcm2S0b/dJ7OwE8qE81Or0tY4OOQzKB4JaBWLo3/BzxyM+euTxTwV3iyvU/DkmzAAq+i
Y3S81MiIGW0WQkyAd/JqVrJFa4/+3NGhRYIntvvS17c70Ynp3rhnDYbNmP4PhznbEtVPMXkbssVD
CicycaTccpK9vq7RmoPiEUbQYCgIzxBe9q8TTdlCHOOFexy6DqxJAnn3E33yWwMPJDHiPyuEvnhH
l026uaSRAEbzy9wdP9X0zadzGnFEcnYU7Eq7zwgcDVaOm0nr2IiWdUPapU8gO4FOvAnQ+XminfoB
Ta/AkDedf8g+K0whGR9FKIY9luneShK6T2ozcNgFgoklRk2zc/WjNd3U+Nn1yhRgBqemUGc+by7n
HEKHRG5pYHUsIEIh+2Ov4LdkeYJWh/Cvmdk6xl9yK6PcGhLkRQ3jK0+ivnsq5LZfIPl1/YeabBpb
gZJlNaXumvVxomFaQLaEYQEcl5pNYCYWiDP0QDrEsVWzqRAyOYz6162r57gzlQtJWr7X1RruQzdN
oPbSMYQrDeN/iRE/yGBZHGlLohtD0CBSDA4I6hT2n3eSU8SAiJmgYvALX9ZN4lOZaBsdyOrF9V2y
FuYpdkTMWOd3OSwWlmUN8WOLt4iOsu/xCen1csjwjzw84NrXplLv0IJ12VuUNYk2nZkkbZdZ2ubg
k0TXNvFiZW9cS3j7LQQgcaBDthLbn3Jc5t3XuY1rBgdrgsa/vJaE8tipCMnB/lfKzlFCZ8bV48SP
COU4Es73Lcp/mcJkH9P4NDb9IOVA94Uo+jssvyzwW2nkG6iDU80WTK3Qdq4InEDocQH27m95WcIf
vetxGHyzuB5AFUoeKSLvQy3pD38GgxDoq8DNqjYmgQfbgnoJ0JRjRZ8n6sCnmdVLoJ8kVFpdTERy
dzRG9Sd1jDcAJ8lzwS948wssVVu7m34yWX8Edjz7jLyNWGQNq3tPmzTHPfLmDzL5y2stCKp0ig50
QIE8PJ+s2F36BSAZC47CaYitfWwNcCpkSumpwuhw80hEfAlJiPuFE2V5BpaYLgDWBDhW36+0008n
ufoDM71mPs5zBwAZrLPMvbZ3uHwXRG9vIaIaOtBJ51Svovo9nCvcepmhMA8AxK4DTKgBhbwNETsb
ewwtIt0bU8p25CnBZEnw+JzR9bz81vIiSagjtYUa0yGBB1HVQx/F7SM3RUPHBFrc2eXFDGxXmPXq
6tQMALnN2OAKHaHcAhAzGxNaZd6m5gWRmMexewxRJVTOUF4fBjLvB9ZjiMX0rBEKqC5NpTQpsu53
fkYUz5W0XPbu/htoD+u6b172amMbpYpsz32cbH/JJzIJ6hJcNabslffHIFaAkjF1RHSsfhhRlwK3
WiSryvGXQM2CV7R9izAc2jZmB0rLQMPdSjerTQ1zniFKVy2haaNiBf1IosLvvgD81cBSofNCwn/e
vqHroyZ6JoiL2jg3RSy24nOL23z0vO0ZahG9OOjSZx8/fi1RdqQWCD/Y6GoPayiKr6bVKipNvhUt
sDXqB7blSNH4ZMJqs36qBOKjLWTWEE9gmtzMR2yd7cYBxgM2NFvuaVLDwc8F+EYWKoElejXqM9Hk
HUdL1NN+Ep9R8in3YGT0fAW42Ny+ODuiU8avhtGO7ktgwOHCEUstx/36YRQp9eOLgVm+ohPbnR3W
oEdaY347Fxn+9TAtCB4DuNY5ekWGx9EZOH2URsjLg8Ua9GesTxfWB/yNdoXEpSVpALBzBO/fcHO+
5+ZF92Kzjg6Citq5iNizSEs35HfWJX9RNasHs1fTfa6TJgOAI7+1LS1tYXJ4QFpcqehiPxkAS6rp
Cu6tozJWlGztLZGkv64OvbiBZ87+HKlGnyeUWBQPY9NJN0U/kUDwHHmar0UA+DyeXI5S+JA32OA4
DJyFRVzJ1VAi5+chMZWKsMvHQUBpiUVWxoEer7qHKCTUWGvpmGvFRgNCS0SXHsXaW+XolW4uxPJM
F8FKiJA/ZYNRzYh4JFu3UHQnKXjtF3bC7KPUtdRFcyV2uB1KJi9FlOuA72GoIPkcnVaeLpQoLltc
wOQBTqHnByXsKvn5bv8TjQU6tHwMFB3QJ2PpKUqNwePjnsv4CCbEfszvoXtO7trGAG+TGluHZoiW
9cJCvYpofhHtJ9Y3Oib3gXlghoYrsBMsJ3vIS1z7CaW3aa8+FD37sqQKtgGOFRQFf5b8j/RALPmW
ct+NCDbvCiK6vohXXPFohLH0gTebw4e5vBHkLzIf2LDDRZ+xNA0meMdDemg2rw9Pq/J/VywDMNMe
wJOI48oypLsQCMKQ3XXUMrqf2m6F64AFf9sxgwnOceaH9BIbVnidkT1rO1NVMiP4677liaZmH11Y
jTD4hT1aah7wMAFa6bNpVNJBGXcxZeTKVeZrU5V+2PsTrSRSpYjFCPcDG+g8eJQ9Hi/5Ty3hpreZ
aB4ZG7/+ovIv+dTl5T8KyKgJqMHIX5BPN+cFWU1/q4f7Z+7dI18YZu9yXUTXRnTz0rJ8A4rqhhk5
akWwKE6sJ/NL01afnGOgHN41ySpP4yqX5wsVnEle1V1N7emyfaWhtB4WuLmoxRKAHYLHzkES6dwj
QBGTsUSF6i2D+TKkkf5354HX7QCgWY+4JU/07uCO7w7UDU6qVJfGr1gwE0vOPiqgGJeg803fmjZi
oBYbcgrZ+mnfZEONn5ubD4TQ72aVOgTGLGrTUbEfyt6vXsC0yUk/QAzi1GqpIMFgAWDzS40k5965
RYRMv0K3HKdTz+y4Y6P2tjhgh4ZheBCw8k4Tne5Ba3R88f2DiCAyNIJ23qRPFnVyuqn/+iRZ+tdn
oVHD5PLzyfr1TpNwTMD/t4lfn/RuVUPqkf0+zYbHuwgADkAAZKx/h+nYEbCpBx4U5vBuN7cj1Kmq
obVjFjrF243z6cSA2n4D6fbEaOULKi5VQbmDRppccS1BxAksT0AJAul/VnFY20u/kpFOljpEVU3Z
S8blDR1Os+xYgMMG0OgO6hZIQtOdIxweKLyT1E6S8M/dYl6uryiL6GtFmJVSUHGq5FAKaYBIuTKW
8HswHRaURAsyd9vtlOzmtI+1tiLKltYF9E3/o4Mpt/XhlfWhBAeNY2vONBJGpHFSU7LyFd1mHtUA
l+TQb+1O5hXiB0bUKARPicYoZmbkGEY64lwza3woAxq1Yge1LzKfbXQm6kzpvbYAB415j008+BdH
qiDrqKIu4fcz1cnpSh4wZYFp3NUpvv5Jk5/DId3IajErxOhgGLIiPT7R5JhVT61PFTluOsvZeZJK
UTB9Xs5gRkEy46+kD/Bj4+FFE+MkkD/pDiO8IqNcGCFc+cga7N63/8EuYrA+KAHcOM5JL71LdlGd
ZBZOOWsJCB8NECcTu7ogfHakg0SO6/JPxd1v69CDs7Ko82w6y2tcrqcS+gC2LCLgWxi6UU4rVUvk
puc/rHqlzGtlTZRMhJorfPKtP2JXjLo+uygW+3EuSISQQ5HqGEuugixMSS8pm6gG7MX9oEfjBio9
3AAGpf9plAI4iV/0/AXfk1OMES0m6NGhi9TFGHf5hOz16AUMEpoSgNJYwX8wDCbtU8TfnEHEkm07
0beZTmNM6xUc7SKFd2FPGHbIzRPWoIy4jzy/FpfSBFX+sc4Idn1lUnDSFrCP8fQNDLIr+K1hXGHh
hOA4zbJD6zuhOPkxLGjf1T4/WPCb9rwpWo9ImPSpcrZqEyugiKIwyOC42hDPeAe1Y6Zx07irkHMp
AnM8fjngDsIB1GPiMGWC+tjjD8ROYz7tmQjiGqj2hg/GpBuNVYMSPA5q9X2HPN8j7YnVqi7NnfUQ
SyfpRMSxvikNCXKjGBLzC9IC4MraHaOhez11IL8Bwqx3O7hdqbpNRijw33Y7HK2tWOknSygUU26Z
p5vv45B/LCtsC83mmgUPvURypFT1W0oQfkzf3RUcwXybLt/yAZB6TwoxgMgcNhw2E+E5ISBgGPOk
OWFGoSr/xMD8ZHpaQTkdWXRW+TO6Y3uCfs9p60O7s6n2z0xh2QQq6meVFCL8SXKYZ2A5cflKBXTO
11noJoO4Bdlhb+ZjFeZAKyObGxmi1F0E4NcIzwwRqHZN6TLydW/ETjBzDuonruM25NxItRUq/A2x
ryun4JMsC1zGYAj1afoFLYunHc1GjcpGs6w/xlwm/tUhULpu8iWhpeZkwT1hcOt4qxfTw75hayqP
dc2tcvZGIVHwsk6YhwYj1b8vDNEhHzIrVK5dOF5mAVX3wHs0ZHIiB3SagQeUbQn4T45DWWyA8Yyp
BCSPB+IELZG+ekLt4oMNmuzb9F8Yk/HqX+Nj7rsWUkjjUUTRp9QMs/eZY2vjJwGC7p38RdGqTjs/
FUF9TWYxABhyaNxMQf0xh06M/w3iw98cv+Xn1iig9gd2AnRmn0p/gci3QJIJBdHxcxgVfCQsxAgD
QMNGNwKAeMiAN0gf3lnfJU4yvOZ4m4aOdpybo9WRVaneQ5Xl4/gDjs1lHCZ1R8cCmEbaIzXRWbgi
CHRZUZd2UwZZvvrat52l3UbX+CfjQXCCpdJv+gBeISUubIXEIbK0vw0qRjLLxhw5XNJH3VZZNUfm
ktFra+a0FR9p2p7n9Hb6tSj99HjZ8bzC1OwP7ZA3floupsL16Kb5TxhhJUMQ2jQVJplLG0MyKroP
MyXKSCDhzLROv5V15Z2tJ5o6OecfeF1wnh70iZ5I0ImzBeB/d50GJh9XXwwg5tZjMDlBqVY8AiVZ
7nJ4Q12G6Ebu4/2JEQvDcntskAwjz2Da5ICAlFF1QSSLMFU/r46zDwWE3SLd4IUaAH73/DAnx6WB
iJzhqgwqTULGeDlmsDrOlm+j4olDTXcrro2b+CwHT2lM9HcndJyG2xVEZosv3tcp8ld0v8yVTFL/
Rz6+EvfYn1bdum3QMV+iENRLsg3EX1ULEbWL73PuxB1DhLk1pL9ukT5PQ+IJXdyAfOdlSSdng7nX
vyGBBhuhWTC71Wd+pTzddBsAlEF+olnru6zNDbf1vSrqCjPpOzkYDtXZyOEU+8fa39ESe+9J+eZP
GiPKIo6iQDsav16KpxQ5TMFpcBcRtjgJ7IISBj/bi4JGDTVTN2BxKaTQNwCEnRKYSOruX+5J70gT
v/5nsRmj+ZyWHdaOFAVdfQBc6G7/XSZHYZUGszp8BqFiEdSboBvF6u+JbNM2cvMqQT/kR6ZxSK+x
4EleyY97U90W5cumdoUAkktwV9/Uf4BbuJZ6deSWB7vEVUQr8iLy9iTK9ONGNbHqBGoHNMAOuS/U
3h9Dyfr0pzMjl0UNOI+55g3igLy+2Kv+MBmY3UvwysX2HpLz4zf6nYGUpCU8rTtVO3WPyNNDQ5KQ
x1oMvr1g3kxVqVT1VVj7EVC7QNZCf9hxlncGIJsXj3/ES1a7VFHnePiuiuxeoIZmDOGp+Tp72WBF
ifXNUT9wwbCnVjUPvjVIS9rNomWLyxLaF9balhzbZgnHHa402Yri7MH1FnP8zSvFX+Kjtu7ppr0q
rnaUirtc/xj64H3RxciLB6isrWwyOANjEfkQXmQQL0g5Uaa8oiah88kZetkd8Xk90OYXs9x5913v
LfmWROXafyTeySj4daSIJRKytMRVrdyMuD4Whjl3nMA0tkRXxGWp8vwiA2PdM5w/HmLoW7IWzp+i
ApofCiWPhwOZejMaayXleNxoR72wGxq5KqdXXL3+9RLmvIJuNSyitlOoylELx2wSMLzkvH0ZV+Bc
BXaA5qPNMkqS04mULiLmH7ggHQl27gCgEyxKbM6svj28GqiWrcWlB089UnzErZNoTK9wnBMwi5MA
VoPY2oZDom0GxnE+W/EXsG+BKiO7oJjIxzNbPV7wdj6w4xPfQf2eTGUoqh6yS8a9ej1aLkfhTrTL
I0ah/vpb97XyKPRGKyxpsMYaaJ4UhXDQFidWBnuoS3iIbFqUE9yA0ZjwSt2HEg8YzjotQ3v8Au+6
Hww7h0w0Thhs35nyb3ljVIO1yLtKlUXO9tKXyeRPMby8yAirkTgb2xJoftf9XNp+8k/LAe1ybQqR
5Rqe9SB+kxM6fZd6RBCF/FOFICLrTKD7sMBdFE7ney94QdvTApsnqcbGwwDn7XaX3U5y0+XvsWCp
4DwSiV5SGnJ6eKFL7QrLWlywFzSr0gOquIaNZwDTLZ+b6vh5tfwNiSINN30m3xJpwapG5Qp09XhZ
oBulsrlkGc/kPGoYgPO1c5rYYrhbXA0+2Hpa5Q4UhuG17m5N0s6lsE/49xQZ7XJStccB8Qz0p1Xh
nt1fhXRYtMWNKpigUj6MmGoq9UTxVThzrKTQTJVDO2/DtuXlC992NlBKO8FyY0EsAl6AcWnI1C92
BusiZLOt4fZK/uY4+g0E/WVqj+iz3Z5MXB3/bS7q+x9eO+DkBZXOY1MeGELsQLSiR8z/Ks8aDHWS
i2Q+nKp4R37dCumjG6CXlpdbES/aYWqEBOlZa0FBGjTqoRZq4Ddai0l4dhiQPOc15/XVh3uaGhq2
eOxKKpHDab9AKks/5UE+x8jpkC9F/2bD/YT3VcPVDHRJXBUcAdho7hYqxBbT9dFFzg4lCD3lLtc2
C0uI9q2/zVSqFuZE1l6IQs7QBTH8LgRuufx506eFL/FadtZLKfNyqhlnKKgFKO03xAlvKUNNe6Et
RaHlyrBFDh7n0tC0dmJGyTzYrsM6G05yVMnDkQ9kq3Cy1hS8tkmScieK3rrNz4gE9EWXkJA6L+7q
VRWrTKLUfYnx3mPbVXrFivdVxuZpW0BPxWG3kgO3qBEdMYm3lYfeSy66hbVoOP1QSA0x7YWu6Lai
h3RnFDUddI36nsi60xytnGb26A9GD17ZzTvFMQy15ApPi0AmW8f180Mu0coKQpky8NIsL+Nio/s0
+r5+KJ1F7aJCQtsRCocySAZ8/EeNj9ugqva537SaVBMv/SmtvWOkXauik6/v6z1OxxnGJ+GZvfAt
5X+ZRo2DjPDeuHUuPfPFYf0Be11pZPNDC1FAeBRb/yGqUa3mZELMbnAwCoO4BU7o+GRT5iX1s5PQ
f1LpLQEzO8qItXKej/Fj7TQkIvlSD0MoHMEOUKnbTYjNyhGTOWkvXvXXpsgEy/hez1KycWweb3OU
qHGJPLtTNsQYZGHBj+pkM5AIUsikr1q/d+VM0m8zsFiKVUi0gHyGVjOWGx98c+3N0UR0FnBf2ifD
bbrYWjdHx7u9+IkR/A5tcbVXS33jv3BGfp+hu+e2D0ZE4aVGQc1q/Ml6k/SDfw4pSbBwDVfCo7Kl
qzD/kxQut8vSNSqTTAX8NUXzhoWv/DFZdMHmCzf4nnQH75+ny7Wf+l25zf7b0oi30oJDF59a2ftj
dKx3uiBrfRLIYXI7wXQY9OrMZwfMqHsZj8Px1wrkqPHvw8LM7s+K5mtYSCBRoS2XmgDaJdKM5yq0
QnPrTcoSSheXWdjwGMPVNLnJBMjD9WyfxUlv5qYJv1EsBHGhsKhCjEJmstBsL/nbK3ldPpuyl/cp
Mlf1N4Cn6923xWWPrlsFowQjxlD3SoDrfimnsCfk1f2J4mYkPI23jjs9lsduEm4hdTIzzyvbdQRH
ZI8g6EccmIDPCWr48w7kLmbyKTzBdGoK5v8mICXqklJ7oZx685ZZmiNLt1SQ/3fkHYX3hPQJAEFI
9Dm4splN8v8xAfFDm/B3W9Cb64BYNTjICuv3H3ohWltedUvJt8RF++h45xiFzvX1ezcqtzqNadCX
cfPOumZ/TdbQa3D3vBvp/abTBQVF557XtRhWjmc4Ri79CbS9BWuninazuQ4XNNXMiADwvaSJRTSl
ekWCjtbX0hsoDeSHw8p2yi7oH919/S2/MPp0GvQ9xNr+nkWhMNLcezrwCCZ2HWZFdpf40RsZLyMJ
4O7cQ4YEOhVRw7tu9n+f+KET5c8vuP389GD5GrlQR+mPJOHSgP8VxZHrnoii5NVo/8RZ+fC1n1gr
0fpQ+QvP6vOKUPtHYsB4t55iSOtefkENaQ7dkJyb+ZCvJsCVvdW0PjkL8YhR8nX7pUiW8Tg6UGy/
dILFOYrJTtcj6tL22FJnLhK7jIh4fPCUbiP5uFvuG/IJL9ieFfQ2hTW6+SYh7QnIWbieOpNvx42T
Nb89P9Kz78CAhZV6t8LKVdHvZpS2sfz167AUI5CorqaErwCkA2zDruu9Ff2F6qlveUbOAwoL9y23
BvR861nK5Aj82YFUqDpjC1UG70ZFJ8JV3wM5F+4cG/mmWGFYIvTj+zF7I49pcmzlVaQbL8UmGTRd
aGZX0Yd5r60jAoDg4TJxlPI0Nb1FuQZ7mnTFMINYdtuC57fqjztn5cGuwSeiWBG7OUNhTXAkHsF2
IiXdb1GBplTjb04uZnrhlVYHkwYWCteNMM6g8mxEbJcHxfBbkafbMMTcfVJR4AWuAZ1lxaMguCld
6sn5oFcnODoNlwGQBPiGLrmdyTYf7zs39WUs5qjulevXccHxryp7pWSbwkLsv0zXEAiS/27x8yFZ
NeY7bdF5YkccFJqCWsHGc69YEKJMJSkK6d1CqTIbuWoNg07SVaUItl7h6SLIYe2/q+x7GidpEY6Z
RRvYT5MhvzqNe9DjLq68Cq3Zr03c/Yofjg4cFbT7kCudNNAGW8JfjIWR3GlNMBgRwaV76fGCSuM1
490pGnjS/GhJt5RyqpP0tWINmq4+mVI5WVSoV8ZV3vmtwlkurVpG+6W8QZJNNm67YZqgd6IKIJMv
QQ6h3rgYm/4Uny2F0cGx4QjeLatu8OJ7KHQg7xqqBiDzTZQzyM0OHsSc/vy6ba9WfXeHqX83Nbgg
Ty1BFbX3f7KoOO9WqH2O566dt1VrCa14cg7d1FWwx+0Mfcp7UDMO0l/EOhhDyxRLVcREp1L9LWkG
J8PZ8Vu+l7wm3W7Rrr57yLEY8o7UPo0KVbhuTTXqQICKqgz6aLICI+hJYXj/A60Scu/TWbmnj/l/
7/mLDjkwidWC37axts3l2qw5PquNqEh4O2ARgaRgtOe2lxc39yyjw0oWCcd6if2e0KhfPEVuSZvk
sJqitIx+ZMOTn3yccWgsmvzq4n7Ql7lAhZUsdQTIJbRsWJkIOoTsIN/wzSDn2FCo3WdYN9ZmFVqA
wWID+SghOBhGqL0xlyP8Pesk4lKKVG2Cve/UXobOwlVOxDyC+RttZmNAUd/OEN2abYdK5drfjUSb
93ABhN2S9k3qeTv/xMFqIyTPl9DoOj70Ogapdh3gu5yOKi6aDhzyAdA7nBiHBswfht6OH7PvUX4v
z/X+9YH1L+OXIoyP0LqlzqQGDGF1Da7EFu83a+vPc5E8Om3KOveYkgNNARXE0FTPgyat/45AZ4o0
1XPTD94BN44smuVrfKd6T7sV3CBbWlgq1NwwdCIWr03cflKDeeH09OlmgA0mIoB722D9uVI4i2QH
5fMvbT/eSyo80qtMlxEmVjhtDqKFU01BaPT5FiE/bTMiTkYMtnN+nLkZ+E+fBLLA6u1eM0mWhGSs
unrcTmp0OzQxs8mwhzo4K8iS5EpVu4ajnLSeCG2qDut6gdKcOJcf9Ff5xuO0+MpI3b2/w6LBySMZ
9ootiLv7pdVNY2nOjLa0wBDkSNuML2e0NJPJm0VXfCTHQCYOd4xvzntEhkV1/J3ot2h84kxenfUP
l+C+tdDLSrA6P5PnjLnGjneOrvgEIf6AX4RRvmCnjGota/dUcSKvFrj6otDuE+YTMxtCYlnD7IeS
0H8k3vytkz0Z8rnu7j+UdbuCwn8mvxIQ6imESq0Z0GIOk3H5DmQ6LWA1dsYMlZQ1Kig9VncmAXb5
tDtqYRaloSLKloW8S8pb29AFa2V9F8Kwe267ryvERnm7FtzTVIBd24uKMxnnEp4EcPP0NTIzH6CL
Y4h0iUQhE2b65FFvPl7IwuQXqhUI9MClihJDOb+UftzNF4xpa3cZmhkBiwa/JbPatA1x5L9M8w43
+Vb8lL6Xi3FLk2T2y0xRNdNff12prIJw6gojIFt0PAnGzq6+mxZh4mNneGtDKGzkOVc2g93DEf4i
FcP6EAtDryFgQN7tpZmR4I4Td5r6BfBIZEb83lY33NJMQwt49JXgaCitiKSwxPMmya7+xk9ibtpB
SdBD9NAQ8k0T/bl9ebzKg+29ndxCUa0FHrI+m7k3md4r+VR3VHKMOJ6sCGjIKcgLW1Mv5hR1zzSc
8PjdwektX5CnGLC2jmjV3CWc69bkvEAHwEtNf96gerfmdlG/Eug1gGfRnlALA29ID7JOttmxsVCh
M4XQuhk6BlBTUFPy8h3ikSl2rvj5UAqd2CXlQIaE3UXkzdYVaT+QRFvy0RdhnQsShPQX2oTsE0Ay
BrC6qpHKhRRpOD/oJOeueSfTnQUYWAGhlUyUqXKbvaG3JAoekaWVU2UJYPiFOrHMsaUER9ACwVqi
xUIgPPfTdQg2pgi068se+yULmurAlTYunoeP8bxXvbDJOHJYsQ8SM03aNyS8O4ACaNumqjq0AHq/
CBNz1V9z/CawDLAMVLTWj98kvNecuF2bZsS2vCIEeP/taX4VGY+1mlWyKHuufSTviBLZWvI1VrP0
rZ8BCD9SsyUSTouBSqwMMHgYkPEwoQhcBQBIgP6YehRywOOQBhBkq3Dl+cT8dwVVg7Pg8Ntkp7jY
dgAc53ekMSh0RnvFDqAvTe0sk9lwcfI7NZEbXt96S3QMRpmYMWy9V/rlydD9bBx8Wqeh4j/yLANv
sDuvVULLtQ+vhS4RxWnHPezrbTZt7Epu2CL53NeWAvE4LJEkJh5ICnoz48HAF7gsv9qgwcOsjI71
9RCgE/maHbF0sTUsPN9lEkajTowdsaD95jb52FsoWc2KHcddkO+A51UZ2Q+A64A+YLo3hhT8MCTa
o1cj+ovLJR+vAN8fcNIL2q48jLmb/bDbDiSUCpwDQb7Gg1Bq+47++tppWZcYitVWQu1NV3FViM1C
zm3dlMXoTeK6sF8d4XNK0dc91FIcczwu1GVb3jMIOGdsOGI9CtKT7y4xco5o3XaT7o0AAxu7GXfx
oclvUPmd+quN1FkWoeQ8GFmLmu0cD9l3A44X9DVgFnmNNBy0Q10cKQAZrmf2FTQt4q69r4+aCw/T
qi/kzLsIFOqQJjN+WDKyGKuW0ktFgu/+fvTo9c+ZUPvqGxMlj03bW0cvlJt3ZF7hOyKRfDvMWX2T
RiwnudF71tpAkYiuc9YRA0uQjVS5E/EDFmGk4wWHMxrVF01iALYSlaN8tXVGp5jwfNQey93pBlDL
c6PXNP+VTADqz6jPOupjsoqAmttaFY5VmQp2fh2/qp21XQLfMeeInXHswGgdSiAZm2qUggCT6+nQ
K22360iCfKyc+XpjNKSvyx9zZ2p0CxTxsnPTliZc/hBs2QG+JCun03Vtu+UF9dxGIgkbVvuMc2oD
Y2TktC9kIfC7Yx+A31EyAZl1SBGhVYn5BZBN8Ox3pNXsNERslwmCXBuKv5jNBz/ViFd9xNNuoJ9K
ZfSMHqcv5OkjqAeMmOt8K2gABSMAA1zb0bduD62CRUrGkofKkFVEJns+YFn/+Y/2HW5iyX8Q6G34
YtgOLlQH2KEg2/9ja/OH81ENN72ptF+4SDvj1H321lqioGlpXzfqh2QU+teNZrqQK3/CmS4V1ygh
u1fEIimJcBxDQVy5h2SaQjkwSyr+iynMOtDTrIARlmhkO0Cm0SOBmGVG5KRcB+xnFefaPyCBI+/T
IkAt9va8OTRQION4O5cIPPFcxA/229R/zMqrtKwhVS9q/WkPCuuVbvhrtlN2HPEJvJjS0MxJtMdP
H/zivOhcd6GYKjfoewS1wWi9QHyIc4NdX3RPzFtaHM9khp703a2wLgcj2Gct0S2Wu7z+y/yq2H2N
Y3U0aE7QHST9giNyn+YTeIiGFWlQ9MpaQTBRw6hXdMpH5eKNZeRXKs3ZSkhfN2r+kTFOvtX6kIO5
D96o8uth1X82gIcZLlGWgG6mBhcdTZc+z1LbYxhyoi1YsWcDQFvHhhmJo6E+5955F7sbRqfPScvK
wm28P7fpsMcx/OtlOItTdDErEpEmedA5NUjnRd3qDmI/u/XTKv8P5ki8lgdpJ4FUXNj3r8RGQ7Pb
zJplAMNqR18d5vuPGONj2uvlyfS+Qww4rvseVMnxGlK4MDKjAxEbwl+XualQUgd8EjqbWM2u0viR
A5KkZiY+Tva7L1tmJjJg8BBLYfGGqAZrhKqujehI07qiK/Jdy2/USQMEvczSYbqUF3p0YZ73fuKa
Uc+U1G9RohEYk+IvlSTpADznmiQsIN5sj7titYHoCX/vHe/ZYGdjvJO0ezGnJCXdenkwqL5wbFov
UsOueaCxvHf2EWLfp78dhULpsLc1Y5MthimUeNRv8xtdieTS/y6M/Cs1ILEB0JF9dh0I016/FBkg
818nDYbTzjOqJ8uOaCeeuiKbL7b/90KdqaJVG9LcQjuwYSSf1lLL2QQJOj8gIMn5g7ZpgRBCzU01
3Y0Lhtqlos1zNXHVXl7f3z58lmUzgkaSAHIrhR01YNsNTF+wMOUBqvf0TfyX1jjW5NNPOZnMyn95
TRg/RpJMOY2nIl/tvHhQRTTw7XzEiirIdnPVyvJyxYG9x3aD5+0TpDegF6Bwqg0qXfFeSIMzOyN0
XDX4FoTdjYX3f30F4UGlIPZ7AkhpqcoN9KLyRttCyhNZvj6ce/yZa2ChEuhptERo9C2I7/aEEuOG
BGyR16Tn1NQSvb/s8g0iZvb+4GAPsSWOnjApWqGmCvOZaD6EPzC/X+lWWQLPl26HwQ+8iFi5k1jY
LKHTIvD7vg4czFJELXreK15w2Mv+OevvDq3lrcf4xo720o7KfdGJiMl1CSBbfUuK4v3eI5ePUy9O
3z95Gcqq2VEEY9LS9MX0YkovWri2iYnuzZtTHEdcvUtXEVqGqNocvOIMW1pT+D+HzuxJcgVNb9rC
msk12weLSC24/S646Xc2t8L8RCnX/oiI4HPPHahs13Vt4M9GCGvaIJwv7YmAXB56hJit/jP/+bOt
C/q3In68qNVfetqxa98thROl5PBQT9cg8oFjKylPOTUDTuDNIDy1bFiLweZUNzJqsXBqn831q3nh
OQAC11FL7Xm2SBikCsnHMFIRPaHztRQAvh/xNGoec9Vrzv/1obtupUgdQBuapnLTG+0mM3szDmGf
MboEXggGLNdbVGMoImRWBQr+dMjY5ZjJzaYZzq0QhlYnzFda1fTFMGY7ER7Hv6h3CLjYVLGQfEy7
watit7pHvOuwSHVesta+jmWca+xrdMOc6NmRDL/z5NEoHapfa5KOu0MuwdTuXFh78osdvnVaKBhW
KQWZSJ2em85L8M4bo0viSkHOQDVhJ4MH9Fyx8JoFUi+c51LQmDVadEpgpD8tGFhah/un01736HtW
Pi7yaXUplaVXtOXI0nDbX8DZmBmDv3f6bX/BMVyRxy00z/C6bkkgWfnUgh7UJXB2CFfkCTnj9MiN
np+oNZqsJxTDJ4L4M489RBvCMHSV389+CiWP6nceTEDjMYGWXO1P1R4lARAVWdwU4GicFsXcfYUS
dMeKGwktpUwBEqdjnTGfpBr0/N1GNd5/Ub8G85TywFoNJO8mZ02Z5sb3l6hUcOgmugQH6yuyEzUi
wiO54F19QJ5i0+VtD7MrgVetrUkeNw0H/cwbmFsiQxl9yRdXDenXlkNtBey+AhTNTc4ON2EzOvtJ
ZRDjOFkMY0sgViWc+2NP3yoffavEHxThpMqyvBcM1iwq4XAJXgROQL3sc7KyB5OKY9qZ5gzJwHsa
pU3XBVpGyKd428eC+YjO7gd7+0VgITjLz5SH+H3EGaNEEYbhCd9KePX0jPFj43AxeEn5cPpC9wwz
3OIjQrwNBZoq0FkoY5iBigP4GVJo/bUE6kuezHWo4v164AU4Mgjy7JcZ7ZAYWa7xg/q0RTHrwvex
0evc/wjvhiIVcflwg3B/Br8DUW7miY6aC51uRO8ulCQbUyrQLTNrZUiCjjS1DbNQjfK+SrtFBitC
gjmvVoPCS2xwUUppq3ThQGXyQ2D2GE20Bxa9zD3fuNc+EdeSSorM1W8j6LLDzGYVVAMtxp0id5Ek
er97z+3RPIWrfrNetvAhZOdWF2J0drvHsvnhQGcdWo2dmwRsBIw/RsHodOA+3iNk/Vrsz8XsYqFz
sPoV3fBw7Rdvgs7qcyJDVLFl7upKnB8VBRwiFIC+VLco4j/bgWPGJ8c+zuhXuWaUbFVP4G6JHgyG
uwyzJOP0/9+y3qknT5vSoljyZ4GSZOVqUsxJ5AHvz/A8IGMfcZ7h+ljyghc/7GMNykMoy1btN2u4
cJODruyOYwsWVi+vtrcnrk2wf7d4Q6kUEyarCNzwgM9pwE/UJUsf+MA3MEdEWdF6vahYrEwiscM0
Mk0rL/WlbqNkb1DkOr6LLLhOpXEH/22PxJACqHP3cGqdb1BAtpagQ+q2KjIMQVoacqHXcEUEc/o3
nc2tXUBPMSz0Qhab58pIHBtAn9t/1u8z6SnMThNZ0a8VGRpedAl91ptkT6eFSe+PtKLc/IG31BKm
Fdx7euU4Xipl+XtE/TY+0v/QNQv5ZupUxyKHtpvBQTR+jIxL+EfrXr+bxbnz7Qmejo3UgC8wG6k8
mUMkUAHAIkUD5sdOoqkMJEvjk4T8eQve+naCAof9wkOGehCPlPwIyj/VAWCMDGdpnvXdhcN5K74Y
jyGn2OJ+qptzYfceCIThGBYT1RKzu8wzAjmFEvbpETSoNUoMOV5+k/Gmaj6GBylhUePLgkq1BBXk
qgsjRUDc5IwuqeD/EqLSTejNjQIE8AOdPZ0LQHgBlZQ2+/dUbpoQjEMEW1DvjLwGdA6/pTZ4GlkG
rqIyS/qPwCy2yy7DJFxT8oLELC6I4rpjABrOGZuK/qtKLfoqiMOfOT5Ko5HarIBzf0UhCgZzIJDZ
Drm1yOz/uz7Q7U8QPmYozS6A0tDjGBbqFKtMwn0ZtV19/alIpIa7misDU25fHpFEgcMWJl335ObZ
aLA7Jw+RvdJc/h0wPZJyd0N1ZBvkMMMLSHFCXR2XeI+CV57mMC2nsBs8O3Oj4D19/ZxfiDwUagOx
FmS0X5pvop0dwNVCld32Z+XMCQDzSKocnvnCJufc889QJdN+G/v2nrW6T/V1ihnNdkZuZ+zgaCkd
2KAU/pyua66D9szxt5k5VWE9A52mPDst40Z+rK5xJLwS+UE9un/rHzlmvsTBjUSd6FkbtIzY58ez
I7rfYGZ2XxWGlwKKPOs2uL2FKPmrAe0YZX7IzE7Lg//ohCPXiu1JZbFogpybIuqv1VBVnzDjxKVL
LBYNu6HqeQuc1N3TAT+dqMk4jZTLBKn+Y6QDDjhDwk/ZgFEOHP8afmZmE79l4QSNXi7mAFUEHCfQ
pDY9fcF209S2OH2/ChdM5o04DLR5oStu5C/k9yXjWSt01EZS5flpzuzBH8N2V5eZMZHnr/Y8UYe5
R4+PwHbYtWUbrpOtb/TaMuW0ZdaQv4vzLyunPcrtJprG2b8i98kXgrXA/vJ3pxlm7o/tf1L/Yh7m
XlftEUuBcw7o3aiUHo9upS71aqQVGFWt+fgq8aKYudel/1azCT+HZeyXpcMBumWcsJUWiCNKlx++
p6yhzUWqs8HJqmDWHUD21j2NcZzza2HiBF5N+tlmiYwyzQ2yk9TcPrjMwDdScUgjTIPwwqxN4Mu+
J1GFsoeGz0f2OE/97SY1/H0VjQ3V5FBKU3cxglBjmUGOG357fa/s0U/6+n96vlSSDd76+8YLtHHB
JzmdQtXTaqPc/CbRKNLtBTWopYU7OBqDAsuNMzcXCuy/A9pyrn9UfpNUkwQMBr2WCKiIgZM1TNjY
xOf/2clO15cFSoh+BEqWs12Er53ynOvLp9JoYHeqJC54+0ACGjJBLZk5V43TfXKnQG1gm1dsLQMf
LneXs+UzgpchfnqWqhFwQExuEZgZwaZ0ETT7X/cAG/Zs8G4SAFKof8rUi6FBa3oNea4kaUCIFJ9u
9FcTcxGs9ZbGCv5AMF52Y0AzRUplhAsvgPTp9b+esCfi2zejfI4jXxtZ4d3K5szdFTX5EYySwQVu
Xka1g3N7a+5uPo/IIj0HC0xPm0vA8+Zf9xoi1UeBjwC68iTCtr50fHFBYIj/KZV7g+bWVJrHj4zw
RWISNU7YNr2fWOV6/ULki0vbMVJnXFnrWop8TrUfaBfoLrfS0xLrcMAbvc5VGRRQLJgwQpO9IY3B
LmvLbzKgn0+KmoH05YnPBuS9578+PyZHhSUL6X47Pbiogjffnr9a4kw7/z5uPqgYR8PMWIoQ1eo6
GC7pieG5JiOs4LYlPn+dQpUGAPPQzoZ4QSXfUytK4FK1K72ABDjRmuEKwb9fSoQ3Gj5DpIcRwGYi
8lsaHvzJH+FsC+7f6PbL9HE6WNWwZlUwSvFwvHTNkeRNypyTEdRB6HfogwzJEzd1aIv7fWMW5hPr
quuwxNPI5ipaEDS8NAv8LH5yh5MFjeCS5Mgzan3+VDfzJQPHd92gx+uZ7Ul7wK9tnlg05gfYQ3WG
Jva5pzjC+AZZg+yQlK3mFLHP/exQSHupy21Sjrfuhi20ZGqxQ9cv8OHQSGvW40DQiuLFcEzS/akY
TEgqBxGsg+5PhY573iY9TVI4YBDLOxBB4OjKbV541MIlFZcWchOr/ebjyPLCxHY8phrkIqTQYyXO
jVIJW7RUh3EUgLo0/XuOBgxBvivaJ4PJgj9fsjm/1U999mcrtn4VMJdeuxeVCSEjoUhUruLEvdg2
AtbYrNxLAvUq70kBAWwKR0VKRPKCZSEGwaHQ8CXWIq/QbPtqSLXgIVkNIeoOe9oB889vQQUnD5cC
1NgsB81st//SDyyyq6O54uz2YG9HoyoNOi/udEQckKq2jJJ0PRuAm+vvX1RKpceP0DNppmCmloOS
/ad4bouojZLoI9OiBW4NtjV7rY0z/J+gX5JhuSdrnGJ2MenP8XJIkqtCsYIWBwbowZOIJSjUUQWu
3TFNvC005o+kD9sT7WM3Mf6a/4A+LUS6KzsI/WzNnY5Of34SSDFRDB2joc9m5/hOElJDpaTOdvLq
Pr1sNBF0zubJatLhrfTZzxVTwSnTT5+EwPIMhUJoP41gnsSAT/Ye/GUIKMGK1XLw7vAdIGprwau2
gRfyo8c2ktr2f/vz0Waci68aI87BADixsJdSTiQdZt2BRAGGMRVUoALelJGKhCIE+fNTC3Z1iTSL
EClAJ4obwbpdb7BR6T4C9qOutx5qxwANR1wZgGDMoHEtYZDMbX6xjmyJxQIhUchHaPkffdmmZlEm
92btDytsK8EjBS4SylbpZN2+9ICITx26BJnW2kbEVfKlPLPpUKr8hBPi1EDPxF8omGm5jneCneAm
YlUB+IG6iP6TvxK7D5d8Iy+WoiLdkk7eu4f5mW+ABnFYMsi82BIm6iCvgXHaGPNvwNn9W5M0nWmd
SeWW8GM7P7uG0rfTmwFdtwXy9vhgsIf1dk7dKKVPUuY3XB2JDdDWS1tsDT3PZ4D/jaDpHw2BAm48
dyaf3bxeXzgWSo5rUrxMFVLY/Vb5Ijp/FkhuER450T3raGytV7xVhqJkKx5Lb467ywaO21+xnkWk
I3soC9qtAmepmJKD9WKt2lrjSHsb5aIU/ZTU+C3sNi+SwiUYLtumQ5rf/6MsNOjiju4L0orCsfzq
NSrbQ2+stAsF0yCBzGkgeUlde8xaAHbc73gtNCsgyeHRGhljR60SXm7xYgZ/ubu0tadjENNqAdd0
NSxs4IijFyxSocKkHcH/nJn6Tt+N6gAe6mhXi+10ConRPljxftBOKrRZi4RZGNK6AeBbuWxuiJOp
plxz9NyZSByBsAKf+/9DJki9Xxw1JzJXUnT6jTsmasIivAZuBCFBtoXk/MpmC/wmZBlKfdIYLM5f
D8xuL7qXyt3SuT6MToE0PpvKmVo4Qo4GoWxQjUQfiIpwrd848a/zC1IgjMK8l17koZAK5SOYYg5p
YehWS6VWIAk8KFzb9AOEdPe9tx6XE8Gisz7RO2FRakYkQ/KS5a0VS7dM13HZaJ6y4ArFYqTloUNL
kjB98GKF2OX+3cMtAHyhBZZo3cS4ob1rjRtBCYUWAA5A8kbupr9/9+EhSvz4OFODak5u3tS0YDUt
HQOXXQmew+EEGxGFYMUct+4edP3wydBhsTRpskkP6+XdwICQNePZ0YaDyGyMBgprKaSdm+P8IwT3
grin5Lo2hdfn8dEntzBM/PcXPm6/DpAEI1KRXh+kkoCDC5MXIB9fJASe3O+wS0LjETpRuHpO0/yZ
09bM5KJIgY1ucW4RNi5tpk4P2tOrJ7sa55mDLI//BjLHcz9IZhpp2qMQQApaCoF8BIc8r3lxb3w4
C+P60BVsM5SrVh//oNfn9Y21gLoOgcLKnpIEWZkDBHPdJ1ljvRRfNuEr/pN5S+cH01Z0trDobruy
66d92XR/3zmCvV9BAIvrZwy3oJTuBUSr+imphYVpuuFepnSDxCozNwQLYee4nZmLSUQGY/KXP+L8
ysJ110IR78hRQigHw0XTJXn0hNFtohkw3OEK55U89DOnd7JM7XN265olHMo+wlOxSY1bokcPBYcf
Tw0pbU+dTzzKdQD3N9hSBWwxJ9x6FYRBVoLQwKknyHnJj2QASamCJ+JMQPBkcJ3O4F2lu+vfDhgJ
FIdFQFbGfvy0nQQeF2BxdNLUV2uApXYyCUKpQkK/R5ROg+6R3cNJEi5y7gyIZiJSwrrC6XNM+nS8
T+/lsdbCVCxln3ZM4eFioTXL+MoOhrSYSoDVbsGFdNShQBuDkHA2v9RrOkKYL8aifviU7Em+Lzlv
tbrGrVV8ID9a4W8MZ2xweZTHuKtjC7q/vWmEwupTNjUIEMJ4L94zRTaQ5fAl8Sbt5Nf6gF0rG5Rb
roSRTcrV7lLDwLmwkF3cSNYR6utV5N7ro3mkvUhfwf4JDccTeNbLiGZndRkXIifX23syU0a4npK5
Oh1li+43KGvsei6nO0GtJ94aTUrtEXsho0+/IaLNEzKUELRQiibjRLKq9/b6nvnRTIyU+iRWeXX6
Cu6gIbO5x6YPEannk3UaDNSkjegqpG33RzwOL45dTfGTbTY7gFiiMk/21YUUHlpff+MGZnpCiNJR
UWC2qNWZqg8BpHqNXmFXEX9UjpcW2vZMCoxizzDAvEmp9W4+8Su8ubxUFJ+XRxBc+uOaKot1SjNu
vJL22OUn/lrvfson5N+OYhwa20t/U7P4LcFj4m4TR6r6NFOTQPok2qt0Wg83tubdmJoN+yf8TE3b
c4PnmH1CEgmjyrIFmWgY9OCrH162CPaGJqpo6PiKFV3o9EHnONaiM2qJZBw+6gFW6d0KGIF2wUe5
M+KgG9oWj8z834mpSsXc2D0IqJmEWRDBZgvXPZjag3eQxIxUfS0c/IKARHo6B0SlZCvsr0PNiJ/T
kCOKC8aQ6EvoMxMfnnUjSV9VIwmTqKzeN2GHmJD63g93r91isTLizJQxR+GR2fPLlmy2iAd9Ckw4
NLF8pxPbM2lHv3zkwrwuwp4FBRlkx4/cUiOmgmZap3zIwlKjvMUOVB5tM9dU/1gt/ecCVKpY/Wyh
jRVRzsQvL7B+C6o6mqnuwkxHGitxM9DbxHO2O+Ah/R2UqGsTjtfP03ObzgyjmfkdTZ3uNLY/5Wbb
23ZwxELKR204aplXel+weIdcWMW8kpkjbZIHYU6kc1ZTp2NokVSc5iAn1aUiSMpVcNmB9vxq2BKt
yIYdWXSm9zzqVcz54LV3zAmT/f9ML2Iyl1QtiBpRJOOBF745frkg98DR/nN9HwprZygbVjl9retz
WgZu0DIK0MNHO2dPcyCcgH43I1n2nuaLu1ZdHAv57lOaVlHyOqcISkDz6WLT37aMCWasGr01KdcJ
MIe1DJrK3Ch6ObQqzLjnlya+2hHbTbZWliPh7YkDzugtE/U6MOBQ8TqennTCEj/3JdmXJKoXA3mw
9AnqMVgCatfn5tTbX/Mh4fpvM81KaxFFRlejWLT62i7EMqRfJrUJNIUODd1HnTeKi32fpwZvQFu2
RXZEQgW8E7R8NWit4lhBg7r32whddwIC5JOlHqurzH1/A1mjUdZAnw9uyHEIgN8+tFXIZc9ZjTTQ
dfovz19b5lH1xz4q+kbeK3bbtR7X9lzQ6T83nJenAK0xKQiEyb8DEszoaJRFew7ZibTeMCJI+1IU
P1tvac42yndvhywb0Z7aiVRI7uod5nfO0dpspzoe+phJM2IN6G3WD3hUlSyJC8ZGk/yOLhC+6uo8
XIPI/zzv2cfunLEc885kWHgkLu0oe3OtHtDt66pUAVwe4x9zGAr3ZA9QR2hHdFwv2cB1WKt7MfV9
SAtPyJPsH7Z1ahQgEXiQG85IruEelxoo/4YkdhqoJKGbR3JuxTLsE9LmUdn1Q/0+59ZKEZliBZsC
QJskeNX1q6Ki2OotI12cETsCmorCb7G2DTKA06GVYioBvDAePD8gPTFM+q9I4ubCbIU1KFVQqTAs
K87/Vux2Or/enFLmTPCoCSJhuthD0wV6iRH7JDp3xeGLmM8yW0vltrUi5/vkrin7WENerFEX6uVE
w5/cnJ4LZb2RafH3SO+GsYrPv0iTOvsV9L8uhlJUuw+3nINVn9DZCdA47QVoASmqB6LDi8wVa9Bq
t/lUuWs2WCDZDZQOsInqRbmi5MylCJxowFO3mR5CfOpFHiV3eP8Jepsjv7951NxAV6jggwrzKjbd
AaxZPw1ZqD2zprhMA31rABer0MpKffP0CseGuvssB9aF3h1XHJRfOQN0BNVweRUVeMhywcIEbD1i
BQs9ry2tyUU7/i9CbyR2UyU0CoknQxQh6+GON+jBSHMP4FdcovVSuK2dLfQTzN1MiK9+GMBXp2D0
lbjmFqzUDaK7fQBmJTn4rqyU46nDEpdcf4nGs+DrNvGXo7LQ7mgQ481pbrxrpxDgpIcHyCC6CuiZ
2c6vixkZ+mAAakWA7/SQ82vGoiDgYk+MpBfaeCq3fUyotoirlNwG25Fr+1fy4iiYxidH6Kw3yPRZ
nKLv6a7imMKzq9g99DjwZUWBy7UydGJblbZ4WrFp0ilXT/Yj451u5/80EFFIaP6eNGDxCAGeG3mB
ghxvQoeSjehp8zBmx1SE4Pis6zNkP3IbvUiB0xKBxZH1/AzuOiLAV8rN0ACGhOCH/eONxWJCwj3P
WBoq0C1lyF9nIZHalIk1gOzVr3/EtAtUDu9SVEJvw7MzX8sE+2DP45F97XMcQwj+MP2Xiu9rVB1O
ROQOwIvyZIbDAj7bjTSpUpRnMGw1wyA5JydjEmQ4aGoJH2jWk6qkI9JyAxbOr2FtgsGFRW/aI2Pt
rMWdW7USpV/yDz1ESDDGzhZVZF89uphBaaQb4ohEMVf7mfVu3sv4oExcjlvqyd93bGn5ukzA0o7H
HRb4skpuNrbS/xx20gXJ2ajyBA2Fi/rXxgYX0PUklqsS1TamAhoXMKpsNAYmPU39mfnwIjn5oWIl
nu5whOhKhmjNGYrzIXJ8R2kmTyX5Ehzea5gq1sbGN7BpFrEL0CP92LdsnE78n2OWKS1+pAgkfF7N
s8RmOSxziMMw9botAdobsw+94yvg1cfKBY8K3hbzbPIT+z9WY3lMgSAKKN8nx52mUExpLRypKVtC
hQZpUP9jk5NtVYkbAlG1ANP+bo0u/xh3oEHFsAtGAkCBs2bQAhBkDcYKao/6drrDWwzVh4fOu76q
AnlhpqJXfWMuCAGm0T2Wan04UkSdJuRh7Md1nYkl7Dd5ct204Z2iom4tdJzh5oFOuiYqRWGJr5Kk
9TsQFL1oD6JbmNqWyxp2znhLqDVlMc2YSTLO7cTf2Jqi8Fh+IqllgsrnuRHzbIRjwtqWLBKS+zLD
VSZOa2unekUyitFO0Dyvh+z1hHP4uaFgXiPllG840GYmo5Z4Xcj43i1e9/O+YCwIZ1W0jLPludoL
dFW+d/mM1z486g4QD9r8lhPq9kadQXl08+nOVyu6sCsgtwzd02zWnQbI7gwEEZNgZxodTKXDSLt7
2urNZAbbJ96MxbZe+C4THUY+wccn+4j8arIKpN4BKHCDcNOhH7adyNjLDuJ6V+SNHtlQO31fSvqX
DFl8stRWCLbFOogukr8n9Kf5AhsyUHxAJGPLio6VP38ImK0siEekmR3MuBCB526pUNG8//qn63aY
svDSLkLnaXxDSrBKmeYG9YxR/SDktUjaMT7ZH+SZbhO3sfu9m1yecxLmdgfMmqPxpDMFEyoS8hNN
4qA799vC7sZu+y5zRwj6JWEB+mCNTEMFLg2BYb06ASzRiSjyYSZGBpStHyzGvLtkZWNnWI82Q4Ys
pL1qCKlE83JCj2pZAWEcCxE4e57WbOO5mmql+IebWftNKygzG51omn6zRfmuSXo2iNGsGVKL6WSK
ExljxEuj7m5crrUjhTyQ8NxHhrTiwqDYp75CUWi/DlCNtHa7WczFDG2jScOZ4TgVruheM3iXETko
xRpOBjv6ulx0agyCWtNw51Kp198MZEz5ErPD3OmCUqkMTMzrMT0a3r9vFUs03P5G/3VuLfKTA0e6
LBcjALsmdKx4ubFdOBRDn4FaT3n2vmmPwPws4DHPXOJJLSyQKbiBEjNdkyLW/vVyYbXuwKjYrYtU
TAAK5XIbq01UflLL5vVCjzFXAagvhv8j4OCxWmvepkTEE8zPMxd+W+a2/dPITnb5INk/YaJiGjo3
+Lk5Liuo1+3XCezCiMeedmjQov092QCjVgDqmF77J5cJNQw27KxNrZgCOzvRuBQXDBmKkPhy95NR
jM3GmAHNnpxtzar0L/Q3/nMSE7CrHvHt3TUCnRsrUxDZnd+mcZYwX5m0AMOI9ulpnWUq+hLg22I9
OXhuWU3QJLCjZjq6bO7cJCVPhJtyarDoTK3TX2dSTfwR/tsNw5g6vFkcH2qQuJry2sQW//roODbC
a56n30dirWwFrIC2Ou/dg0qUORwZQ1rZSpZxptGffAEEGpkwtYPXbrmGJ5kS+455APB/9um8ocCa
oRj/gyvbAgLVDxlgq+5HMQ4WoXMrEc41oTixcGVWlh+bUaFKuD/9F9viMFx5X3Zu0VnQI7aIAoHw
Hmij7hUREL2/hCBwbcMcurN5yoV+FsK8OFKhlViGUmdB0EXoHAjCkFfe2ro1wQ4CL8UIY7boyQTo
toP9rWzRWraOcYYnsQegERNFunma4pz07ZzUtZYSH/KWD7nRb/548jxq0yONZejC+Bw38I0Hb0hA
LlcvcpkCNd08g//T/J8a/3gihE+jf4lXakL5Bh31WzraP9gAj0IDGh4dtFaEAKOY0ZnEwc/9netq
ln12X6Js8F4oEctTEs7ubsJ3LcVNM6fUMv/Mqvq20/9zo5ladQhlHY/eTAebWybNzRNX8nv8v+Ga
CW39R3c82eFgKpMEi0acI98Frq+Dw2VTzc7hnR9s4gDmbgL0BioWbnI2VJGcxCzsEVU9IaoQGpZT
JteLOBgqR1NAcC6dddHle1TFjieM8i3BJRKqTl++V4lbXYLxkNsM/itNxFqn50eMVJu9T/zBja4O
8oeNGK+CuhHBRvr/KPx7NrcNiO/8IZOrQ+kvDKMGmgkiUQVlH1WxkHp8BCM91ZiewvOffwANIPPq
ifRXbiXvymqqsF+tjADjUsMdkHQOBZ5+MU5+0y0YvNCorz9UCGUred18jAaM9vRE7JDTmei4KJyL
cqCNieGVzwVbHFz8DlnF026bRBB/G24krm7BwQU+bMXX3f6uFjE6/su72IdzLilQhnGxTKK2BTM4
++UXhK/x8opFF2b4SMWy6PB/NXnGEGoAedb+PUhoIeZOlwJXfMPvBbaTGqrkj+PCJhNptcqKrHAF
Kn1RAckFIxLpEjLz0qhs4VVvWePy+Oa/iIYbCDW2N3NZ+5nGDi9L5m6DS+0gSF1WCvOS4Z95fUDw
OteSlQSMzuA5eZI40LdvehQiHa87brpfpDfsRbAKOLCifHJLxdPNNOY99Z14BveQPimqD+OU/rot
wHcVDbmyYCLH8kCeOYLBuUIi2oyhgXg5cp3d0IjnWoFMGx6iJfq4gkc9qksmnSbJLO/2SczrwZIs
TK4P8WEjnCn146GkABWhke/TTPlxux02IAauWoAyraswLs/zWcVhvi8X2/giVol1dpioYTXBZF91
chmTykN3I+v48zAxOEpU/NeNlpiJYP1+jc2VOy4Lmyw99yzMVdAznd1eCz5Or20aSmjPj/0pBSFH
GwU13X3O8pUeMhlUB+aXoRZ4VGGJyR3g9ZvNQnzH0RAj4JdgpharQYVZ9fGLfmjw13ZVKOa6vAKI
rR1CHxZ0IvfITIsuedXMfsigqfEySbfxLkZC4rKpTIQTbR5U3uFggpuLuj/rWepVi8LKEcluXDQ5
R7X0Rl2BDZjKi0jyr76WQ/uZnHeSyrNpOcgnbnchpVFqNyIkkdu2J/cOxg53s27Krx3hzGlS8foz
Znis5U/64DbudA+T24Zif4+W0Rcgv+otwwDNv6dQy6HUtKh1AwE2dFo7CGfXBh4/pnK6u6zwx2Kt
jykpoLayM2+WoAti7cUi1Rc6P1AYjnbwSdHMv1CAYgZx9adGBWVOJQv6HOFeDXr5cngsxQjARMiP
nRCEXTttB73ZZ35/W5yrgtW4eGl6dukOXmWkXa5gKARqMtc+7NgVNex0eXHeGMa0fNFkSDZCv199
WK+GQBlw32rrS0+tJzI2O6THG7lFNWmW7NygZ+nGMPGhGHNd/GTeDrQjC2U0T9osAbGdN8yPyprf
e72cj9uus75bb+oq/lkkfS8BnfX7Mljh2VbNBcvkJR8nniOLYMwcacGWGpSvGjhE00NLdtK9RIqr
ZkR3xe8c5KFzz3NYYmlMFlwgxkbHZ5APqx8TrlCKxSS3iJ2A+Hx2wgnIyo4WllImYFFS3VjgFY6h
WDW3MjeAlYbZo58QcnAN7duzQ6JZC3o2W+VqeA4HltWbBywkq+rcW1VqVooXPINhokewifeiljbZ
4yvmUmC5f2HIn+C9YIDXQfdnbjhL9581OmIdBVmRMRnzOpN1ZcDf/LKGwqOkOaYjL/xQIK1Haxa1
DRjAbRihzohUDxRkRHEkFlBhkQL0arKC9fytC4nZoz6yfGUoAMQdfXrTnF0UmaJEhaeYEFx8rqOd
tjFzTFDUvNW/IG6i1GCa5UBlU8OlFaa61fAe155DDkPpr81P0m9X/Mx0tCrqQMEb2Vltf6C1ut+3
+ASBJlyiNOXx53ust9+HFvF3DXzBjnxuDkFNhqBLXeRmk0zEZSQhloDCv1WKEbLBCmGE2MM0VadX
a63crGXWgVcsvSyIFwAOe2JWpldtqCx6ovKJvlZm4+C7jk0U/DJ39GlwUD3u0aekAg6jLM4ZUZRv
thyxIJqxgIqjm9/1Z7VcY0hFRrjI4FaNO3t/LFhPGinv+oD7UNH7aFzpqLHiuMcmsM5A2k1q4lWC
bxfmcyaCln+wtQ+bI6HuGj12cdk39R+wtxG/FAzNlene6MfBYrK+ZPPxHJ/sFvP2nSVYwhkawUMY
6boqq5k62fQwYV+fqv2VEwJDzbGTyMXg6yzOu6Yq98egSzQO03E3VPad5qiOqx7Ss9smtmIeeqNu
72jIfgL4Cqmx3BYU6Ycy9fJN7Vo4Qlumez9v8RStgS2IVPQBXbUxjahIq0ut2F8feOPy3unqTB0A
UNhP8SqsfIaZKEouuHoERAsyIrwKIXt252EiZkMuIVYEMc2COlzGsZQ3S/2tPks0EaOToUeT9Rdg
AJTIcSC4JldhIe6ilawhVkIT18Hs2JtfRAW01H/qiw7gpOTFS9jNigxZh2JsurF3ZT3uJFhykknL
ViAPTI19M1O2gfKrAJldxnaHnxXvOBszWezcfiQZEJ/q0wKPcBppjlTRXZpe8zzuzLDCIfifrqvn
lRNi7clNAT8VMFWD3d6Yt1u1OZbydc/TP/jgWXEiWvBFPnooOWN50gtB6lvcIOepz6BzVSKV8iUg
O5ml8byFY5yvqUekAEtq1MbdiaeJIEqyCo6n0cmv9+BAEBgvKUIw1z+XXais9cjTZbzfgLHJqcpt
u060pSigpAY2SZ8xy1B3EiM+r66kPHs8ryEF50OJ826rGjfNDqRLAXTSt5q4pVFh/2Xp4oZrS2XY
d/fsP+79wWbu0c8StXjr1L5j5DX8HH2DS5+xJf+AMUy3IUlLg+hc4/YN4G4RZ4fF651tY73I3Bdg
EN8rcnkJKSG0EwjmRKJs9kEiRzAkw4btff0t6pBzjKOCoxjsNxTIy0JZW0qQRpNc6caQ241zmJji
IltLnXbqprHwF/fIxEeHZh8i6ZdUcKxOMdzc9I8s2jBo3MqRsHLqZP/6/TX/9QBRIoDPdUEune16
k5uW6FtpYwtHJCwhg9aAxmyYgj8mim41Kvuq5Tt49ffRSul3eR6F4pAwhQ8BaIMSr2+U39sLmBMj
5ZHj9sE0PP+0EuthLNw1ec4t7YsdRyKSxsP7a8+quv3QIzK/78NpDaFDKJ4BgrgaYYdEdsmRpVNL
3oNpVy+CtAj8Wxg1PmkuJ0/TXI625fEc3mBVm9UJ7fJWqm+nWlMO5HgeVhnh90Z4b88nAPMsf/ET
SUBsGe/ICMoZxdeCNRIsmdltVcukWgbbh3zrSvCnkXPAiEuDADirlvf84EsFZdxVVqIWQh/B8qV9
7cqG+dZJglifGsGrvDuXQtyCDSotkpPsEiJy1KZMGWiE8b7T/smOFvUal5AIAbFanDsaUA4HvFU6
2pY9fUeuhGivJRmbzIAVrjMEprX7Dl4zOElRkVROyKPC0biLGvknE5yaYfIVRfG2rdpUEu0LHwaw
NQxmF3/twPrel9DHr1Q9Dr7v/1lRxmBss8moLGLNhHjiJr928TcGLYWl2AqLdPCSdFHNX5fU3IyE
lStUHgWOUDa3GUpXsT7Uw3Nf+otOnexB2b4fvBnYcl7J2l+8tS5raWmcuXShqNOV4kzRnFriNXzr
fd/GeeYoIkzuao37/F4ilOU608XveCJ0bPzITjDto+77+9ivhZcj8PtKPQnykE+PU5hRYCxTUz5I
N1tayRTOQqACfP/HciL5Z3hK0loNkdZpKhQFRwEYR0yMkbTaH1dsaWwd2eSi8i1vhpmFFDadJNMg
0TjJp0/YlXWo/HZ/USQ8MHcpubhInGZRMlxoaFpUcEy6TzgvPtB2FOAae/Eke8A+J6t8XABstxmf
iFwn0tLMzDLKNZ14j5in9xIAY6EgPiMbhAMmB76bMKpfIxLPueYnJ5/+9VFULA2kJutQ1W+8mB/m
TRGbMCKczBA+TlYdrxpMpejLwKlsm8GvsunPyI29YBXv43vb1Z3HQhojlwjMxfxx/ujUh3Rr+lAK
hSs18AJDqM6HNL7WX+hm+ua18P+xuSWXa6eokkEF0juTSaW6/tfdGk7HsySO5YffqN8O01I4fqzF
uzfKHQ9z+WH1O15TnweMo4tVrXaty+jU2Av7ubP3NaGVEJRcGyzGs+9LoxindToDciIRzc0XSytl
AtvTdjZbZr7Mcb6etjzhtyo5oZ2E5Mka2rp3/+2b4801F6R/+e99HnmxNJL0G0oZdmptZoNN2Nu/
sjH1DFN+9T8QicOl/rN8LsYDHscX3DC8+4VZKBB2Q6WshxMWb7jTKUpbXuCVPvC8CmKHsGbxjtid
Q1yzn9zaj/kOxnyQ45n8vFZDACYlNqUdki//3aGgvHOC350NKDVw4Y9yeA6ePh9VdMY/aPfKVddr
j7sIsdSrNXBOELo5P/knFaHKSJ25C5c9BfXDakLwjBNIelRpah5pTZffDEAbnHLTdfNIk+dNq6Tm
cQ5CKf+NwgMIKopcRxGa3A1KFjd/aBAqbBVVaFT689B9u+Z3klIFw7+YzWqX9r+qavjmwM4fKvum
rLXEdF9BFf/oSRIyJKTTa5uaHtNHEmG0KNP8Jeg8Vzv5E3Tjk8SEHqV6NWaUx2xzNnLUAxi8fj4z
Xyhz6HJnE6whVJQ/f8jnzK+No34Wtw0S/xpLKvPmrnAFRcnAFq/GFwvsX35vpIyDczm2m7xtHASL
+Xcmbj3zGu1p43r4LdyBKcc1TdgpOpDLRGGmbx3NELo8KZoMlp6bw6+3bGloARK4+Y4OxAHM8cqX
thQqXEitfsazSXowGJtM5FRKKIJSnQVzDb0KslFWfL5z477pmEYaH/vIAAmj404Oiar40yM9hmAU
hkEFmP13XUyabLhetrQo8divicdvSyXKbJS/lRetuLZu/FXUXflHXDNLnk7NH1suOn4htTkijnPx
A38iXVLW8PL8Rj7YNS6VO2z5zx/yzjlIz4LKZ17fxs2DJYcwnrxyqT3cERB4cGbCXBqA12bi4Syj
Nr4XBcdZQxqGyCRCCaJIQWRVegPv0OzMxgbXwaFTvWr2G8BdECvdEEfY/ND321RgucaT+QQKkkVC
mj/DYCyjw2WEsAuYotPCXBqQ0Re6/Y7aW7gbwOX6R6YnFceY3yzxkWfsX76nl/GUQ75YB5TII+9b
EoxQq3Gfc060m8ECZPRrumeafBNbUpSDvuIXG+uPSX7emvDtl5Oh+8lJ8vsy4qeJst+KuZnhSNIt
ZxBb/4Jby/xz707mrV+yJ5WtXlbLal5zbVwubJPVBTifOSxHkGXpLbNEHy8BUDDSAb8GhBeK101J
wGriCJvjEZ9wpU94tZ0U4UDhD0clVNdx/6g2UAV3g+qOu6DSKHEQyNouVb6OLbCazF9p9nvMXwAL
EOtbepiZxDmSU2rN1AOvtCq1ZpYmohvJINkMqJTETlUB8RUzZjIozvvMTVCZg8SUQCUaUIwRKPiw
a7ygW+8rDW7XTPT5qFBCQD/UIzX42IC2aPrhKRAWveMDwe7XXL3i41d6vtnbk4TQSbh5efSgOcHp
qKq1QyxS9mmAEzRVEa1z8ZUPcs9mrAtaro8eyBTA+jY7mEUQ3euY758Mmd8mql/zzVoYQzke2XaI
XnLUSYr+qVCkIxi6/C/yo8dVEah3UwjG0BtZSQqvx8XTIWhvRFJWzFHrt8bywzUEpdFpzBUZcUVO
NZfdmc3I/vJR4fE8ODy6AAGSN6JbGuUaLwn6ToH2u/014yhQAB9u2w1qQklaA7gQ90pM99brtiLv
+ptTI1GYbLhCU5CXblwp2mBWVyvxMPizNDpen+PqFE7pKKH1Np4o1bXoEVr4wGrhZ4yyssE0qALA
YigLYp3+1KAotGcFm8JHN3dbg8AAalzRZH4GTT0ss+hlZRcFr3cKbx9EmyBHM+6JLsnbOFXbwhgg
5HyyNdlmD2rcaugUc89vGrh4crxAuG3JJpQI+hBCWh8ZnAn6Tg73Y8Zq/UYLWFUSLMquKopZTtK0
FBQabSOvG0U50+m5ey3R6uIGXcsZWLOUWhln3eg+wiHv1CSq5K3RjbSJKlG4BtTnfwTVdD2oTZIg
gl5KOhWsrODFuzUC6dIEqcAKoopPGURf3MfCNYusWI2nZzUJIzdSrf6xYK4dlWTJoRTVQrPzAp1H
juLLcX81cqBCtISFdgOwUt7h1VqwCvRTOFNvGSxBr0W8IeOZICohjkg9VKsb3L14ChwUW5zIVNvw
eUBxMLba3orRlz9cTBG+S+gyU/2eFbL2PejP0tYB9uR/vAxT2E2I1aUbiFJoNUCMSJOTiy+5QSW6
JTN+GbXn75xxTLL/fx8X2msLyPVhB/Ic2DWCXvMDqHgNC/8dKyo4OMx6HPXBMBpfOicVulXohhXf
ozWJeM57ohjDAu1jAzbZ2FnTytAYs4cnctcHdspA8DBLYR9VIHJQYpRtxFgj0C+WT4Y8F5Sw62GK
rm8FW+EXWcC+Rvct8ZdZBA+pXE4po+azYDA5lWcCTxfI7sHYrQAuR3vDRqFt5jIgr/zRK1WoZT9H
dGWWQImPMxAQjVNEQ00GtduVSoVW/LfC9/SPUJnrp2WOqxufQYPS10ZNGEYDXsP9xjcUd1NjnB1k
dfalz7dmMwz1zLbQhFYzB42i/AP/yZHTEMfgOwr2Ql+EOlmKBPF2WiPup5zXaTmsGlJMjMddC+b1
UJmB0EnPVaJV3nDJrrFjwAHfXbL/ROixJGFAs4pSRGIoahTs8PfUnfJIkbM51a+qPKQbe6ogj+oZ
+kOkbuFXJ/AhcCdAwqK/o6WnsdmT9EBA0DS4MGTeFrYIt7PcrM9sbANejkgTRC67jxMF53KTmFSX
gROGJ7DiR+v24Wx5gk2rWz6fn+5mvmdWhpr+l9ckLWrR90XCsVah5hQykmd1vwniksqcQ12BrFER
a28XZ0zHePhJMiX67twk/K8sS7YS/5sluYxsIJwjX4Om/cEQ4syF0+6pwLSuxwm6+r0t8G28RSI+
K/z9W1+miK9RIPhtwTpCKvPZBwOfxmbh1akJjPNMrvO2Ige+88XrnUNDfBzHsJu6VeV304+oDkxE
ucyW51+MboKinLxTrzjQWnLP/fgqS1Xv28IHqZDAaNAwK7oWv1v8BfO0UKRMXTXo5tW7GYKXk8ej
D5NzTYFQKV/Q4vGUjSZV04xd8ZnFItqZ/3sk5sqhHi3PRmBGO0mb7AmOBK3kOe9B26V8bleNwo0d
6jpzCREEC+d3IOAc8YG7UuJuq0FFBQn8aQi82n8GA+mbiNDpEV+ewgKjEfgxiUtGU0UOPtoEC249
3Wf/+KbzdQ7C+HceX7WRinbRQ8T4ivW+kHdWEqGwr+CBgks0rZeRMtlfUAQwhB1QWyaVs0wRQvwR
tsjFaNRuNQ+eVMWDRtSOwam+5LSnf6ihWKoNzBqV5EdzWi1hwkTEnWJrt+fljs5LbC9PBRpJMpmg
aitS+IwWOixzPfm8vHSeHwN2hOvi8CkYNMCy8AeCEqPHl7z1c7FHmDZAfa9hYntCca1tUHyc+ak1
0JL6LXxYeAh47/W9AXhCHoL6DPO4sWmdf5fEq6osHUv2B24y7GB10/w74zJmPsgXVrkXP7M7+W+J
Pjj21OaL01IpibE2Z4f/ed78zlmc3ZggAh0z1YrPYJOvJZOunrqI/rLHlw4UJEMhckxIV2w+Mmr4
OxatU9RsOvFA3wp2prfsCBqfiZQ6pyA0ckhxjoRZMUOZbjZGtdGKsAsotYkbpaxplM3y9phz/zUf
FlvPmlQpLKA94lO6fqOMVQmdDq0ZildMDrWxlYiA5SqQwLRkcUQkdI5y3YykEa64lYLcGxwv+RKc
lxoFgP9+Kt+hQq/s1jScJdqURd/hXjeKOo2D54usF2Wp+/arSKXjfsOUyM968xgpHqdP7k0ut8/c
JbWbs/hnHovd+9JBH9QHti27msk655OeiU55rR782E9oVsajMWy+NCb262bRj4w+QD62b4RZR4N6
1zlbn8Aih3x/F4XPDq3bYdx7XEVcskCs1FAKQo4z9A1mr/Teds8ndEBvPT8Wi53kNsa+juIIAGsx
kSI2CRiY4O5gg3YqEK2ObHMTxssJfxfSjLvDRf1Lo+OUVQ0JUgqdnGhd+SH/XH6DT5EuU3V5nyeD
i5pDssHRKcuogPQQ4O7nWff/v4qhYV7QEe2ldmFj4T+mFClNnV4bEUyu71rx7d1qGL5PuT8slLhf
k99MBL3DL6qnQVFbdsZASwOHD6L2Olg4O8rTIz8iIuWtitTNufegqjl9E2GHVntwvFmPBmQ+/mqF
hFv49bxdq/1bmhaeIRJ3/vaUutc9YdaGxD5PhkxV5cEuSbBuwFgjuYyH0aAKkqGGW6E08PZNu/xm
sc55ROiuLVUTbG5VzditSpbolhvUGC1UIUcyuRMfdCFFbaKnFQ0tqOzCLM2OPVJgnVFFRkHAyVYM
OgCFcIRsHx60WDHjnYPjJAXFlUV5DSrBsaJNCgLClIRO97sun/ZG1cULjJiXU2aWJX7lIikzENao
StO/vt+nbDKzJhtaaP7dm3ufKBOXyeavcdnXGLPLJIttyPq48S6NQHmfqOWD6f1xFkQcVQFJrtKD
7CqODUZnMFb8elvRGekAcvKmvWkJ8JzPR98gELqvQLSy/VlFj+dDiG2adhzpJyvB2GAICdTdBoP9
rqsNuL9NPmrJ8K+ypXVhG5MYfNVIu4cjCZTEDeKKdkw2fOcOdYBIgaL6JKSLhMhu4H7a+JVpYDNs
poSGfz4ezJLcl8DQ7yrVssS1t80DQ/gHD98nCcCb+99j4kG4UNO+P7YStyv+QcOOfAbCDvhQ2DCK
upLcJ0oWIODoVEuo2Wfn4KJh+8DaL/NDF/6AMleFT3jdkmhnW8xJoP2jIjpG4wrSoTRsFPvLBhfO
CGDdxO29MMnkveegs0StM7bKEs9P8/s6bPJbfaJtxxHl2uXtFShIo/PSk4UQ/i9XNEFMRz5Sp8zf
/L95aKnNwk4nbcnmZIns8Me3+1qKfmvaxmA8DX3z7t/sI5nMyojbPR1fflDD9dKjqNvaHdbpDn14
JjfDqoa+VqHUKSD8GlVkHs6gjFKCobHOCq+CLin/11tYxqD3areDCSCSk4Dh7PvO9xKwZxMVrTfE
uD21FhP1Wq74I2BSTxcBfFe0XDKqqJcpuCJuvPsoB1xBTtOCNG6jFXPqAq0Zeim36Er3pwl8lv3x
FjVtvbiBsn4lPhwbRG635mNDVpAByc9uWzb8dr66kzT7nMAArp6430T3ztQBwpTU7Qhhf/1mpmb+
yBCyWiv2s0pzzK3bZUR7JtN60T3UKaSmFqxuFRZ+Q7LuEyToA2TuNHUSrcPpzrvOvTjp56JaSgD8
pbFcIcrdOzMu+0jIDPpWMnmQZfBQIKOU1MKSUBfLa3qmbvzY4BwyxKgT30axLcdpifYTbTIjLRbc
V+gzMRGNAhy/LlOn4NH5OY/kcvORsLj0QQUznod4C10i+MYuwsNhQ6l6V7ieyljvS7EyVjtN8gR1
sadxnbCOPWc2DTMPCWa0VILmxOQ2rXodf8tZVj/hfJ4cz07CEBRe/arLnKspYb1c80ptbw7BPnCU
sjpwQbqAlxgm1P0AjrQZlTE7oXuUxIaWzwFMGw5kCFTyEixPYLlLLn17juiUBUYszKpFLLiem3vf
Pm586TXeJwrbkO7ZFj53MXeuBd77gqK/HbBi3bLL2fuFZOcU/HjMulhDyCbdTN00ZPQHVm8jTlU4
x/wT7T8IWUbjlIvoqEeIVyHeh5PcE+k+Rr0P4LIUOqiJQRL494wDS6xh7EyzNdRBjoyP931BBp5P
oUZzaoVVRkj1QyIbGZA8guSrbTGy5mROdxKJakw5NnyQoqJ/zEG8Ln19cpuEueZqlMMWf3edACFt
fvv6pxBV8/maqxCaoqMENZLAa76xiCNnR+dXbLoqCW2zqihZtUVV8KuZs0X5RAXG3j8WCikUGUpH
3HYAMvqER9dzTx+Wbds06S+swHK6GV3h73UaVd52IswgzJDsUlCP2hRL1Svto6KSdYlZs16RMEU+
ISMOzaPI0R1WRkcMvu7281DhG4pB3xP1NQLwch87E4yysHa6EClkJCvysuL+uT/U9von+N+7Qt3S
9ZZ1ezRYYmaovVw+YpqiP1cUttBsDhbbFIjeOeIcu5lXVEp9eIFIiyNY9hkNbIk11kTQfL2yaVZr
FOPZ/Cvgic4BYa+/Hh2KAhOy2eX4yYLwW+PidGGWg82wold0ahMsIvxsBCv7yGr68W0KeZBwIj1s
BtmNjV8dBj5ezj5HiR0FzRUIKJVjVY3pBYmatPVZR9fBriuxsAxezddtJl/toxFficpnih3QLodf
ZCD3ggb6syXx5UoXcRupMkHCivTl70/JVTNE6wtOqZpsOHDxlUaqeBKylkwu4jBrQTP7zUdHA4n6
SJTEIcpLLk+VJeibtD5bPDLkHGYuMOHXLuiAWVH6sS3ZN7AgfjmcTcxuYZaVxYmzBZa+bhcPBGbE
7BQ4UcPybxfmbeR9XKoyt0EKq9GXtkXDZ8pdq+c++HqcvWvvDZNyLEtcTmrT8QfP60DOEXHMUrbx
+DX6hpGa4ykIYt6ANE5igkOIbKesR1W+swHgxzIjl09LXP6Hgr1aT2it/KdF3cP8uXfbaIC8OOPC
gBJsFXYACnMwUk1LHo6KzE6sepBUao8Q5U7aq/gp6uYwQG4zBKoS0dwoxMsx3XdUwxwqIcIVOJiT
ji2syJXYMKfpN/WqCO+b9R8ST8fp0PDQRZZ08sfGI4efnujGAsjtZaguu2RMTi7LLlAgEmUcWJ9V
LWY7TE/vFTbZGIbjWpbUus1/67ag2F3bS52rbeO/CacIKGGRYvI5LeqKXfyf6cuRenJxRHSwEv0V
veiDJEl+Jd5tkFbiA90I4A0JdOqKwNP3v8Ozq79EHCgwrRkLZRXeUakNxU9ZaOyS9WPA03NBIxCY
yeObXW2zPBx5ubVAdwWJ73obRYuMhHTCqAvqUnuT0icIGJRxEyMgjcb0vhRmVjHXIX+eogrlGE9d
qI1NmefmuY2aJcHbDZKpbwqdWYw3uTGcZTgown6SDb+pRozdIXRgFvCHyqPdjb8SVBl0Vug52dpn
txYTwBuILh9Dy64cMBR6FrTljyp5mnsrkG1rR7lPo4JxOls36YI+SYC2U0wumx3qBpgqZ1RZdadH
g6T1KcYDGBcSw6aaEYP45vLsZv5hCsea4OXFhCVDVRGa0I3Mj1pNCckHdGVRakS+leysWGNQk8E7
d2dHtbhK4Faj6c7Vg+Ag3SrMJ2gQcyMzK4AdazJeNQBWn4kPP6PrN8s3Qm+9Z9gP0/vm1YMcXH4b
wMur8tqWd9/spoRyQsN+2DcCpGJhoftjgdctbS9TOByhd9tWh106p/71k3IYY0TF/Y6HD20de8FD
5A3SbEePmdERjhhippRrV8chK3I3ygy29rTjPpI+f6B8398KnTR7p1/zUzlGwjfoQqOHfSXegROD
nnw160kFw0hD62Zd856642UW8Y7xAtbytllwT6adiLsbdYOLDEElMtaXJCIUWc1yuPnyb3JfS2tH
1n6JnSN8BryiSL1qSEyPUS+VAywZE8m6sh6PP1jdNFpTiQugJXhdGEZb+gWvT44I86p2SYDLeFrQ
Pv6Lifkq1I0vbizk3rWX0WsU48Ly3b2QTs104JhrVg8WidjiSplzEiHcrB1GmCZpTSkEOxDxRSC7
RtQEDfyl9B0U6Y3mT17GxuxntFeCRDYd0HJSLAb9W/NXb4tpDWQI3f2qqGwvfLDg9bGTm6qAfEMS
HwL7mRg7Cb3Qq27bEkncO8GSlJ9+OSK7LMTgDrkOWeriwSYKk3kUxirWqCQ+YJ5Zbo8DmYm2uz9K
sIDs0K/1pcxLg2FzB0qiMwe29m43WcsTzshgKaOdt+nH++L5f0OM+ghLOlZ4iCSVnVJPfXR5QbJt
nYi/v1Y1xbsBI4cn53W1f7NksnQ0RPg0y8iUdKGm3bTx/nGCMlZ5a1IvxuxWt75uULToNPqH6QeO
Pfg1TPDbQHDZItUvc0FevvD315OLrGNLDZSLZBYr5qzNe8gdMObv/nCJ29Ltg8T9tHPLsl/w3tkS
pkl/x8IgBSZnxaFOPtQBesV3ak67hGjod2b5zL7XDjGB0cihHyctJybYiaHitweYvvhUBpCyzoCv
1o5A4fvZQa3K5LTNcsnr69ELiF6UnAmj10gXWZZ+V3sMxGZQ1L9hn2tAwFd9x7Vl6F6C6sLu+bR4
ebQPgIH8+aET79Q5mp48YfCPVo4AU96Uy2KJNic5JXFVO/fbf5kxcQoHfFRyo2/FQ00cdST/zVAf
W9OL9O+3ejOAO1fc08Tp74EY37SQOAQDPN6hMwNkXY4YQ3CC2JTjCjH1v1Xvy8brI9HesT48u2/N
uevgkaGZCa5dIxkkXBlXjvx5QA4TCZV55MYdYbV4pwuJtdQzwuhYG9Gc7Y+lDPOjcm/6eSaP7jKo
OIB33h+tWjTpgVL4ZV2fSe11XEvtChsYpWGY6RLZZ2wm37OFzSJrXZj1gZm6vXcwmJVaqpfM8zxs
8e46VNPzTImxD75P7ucSQ9Bt1G6+XZupYxfZvEEaPE5y/UHtspJ51htaCrgultkpLsypjDw0eS3G
mu+7vzGJHndBvUrGBxVmvNj3vT8+7Qp9xAuxfGJkuKR0cMNjIgBsnzy1uKMmP48waERGT+mGHKUb
0/T+OmdrJsHUqwLHS/MmOTAyL2LfWDzmrEAPG6M9enYcytrdGA7i2OAfWDl9muuHRRXlnnTnN2FM
tYnutfzGkww9oO+SXD5NW1imyeSt17266rQ1JgStHVID84Nw80i8P/xwmnxzEhI9xgiQvkje3ND5
I9QD4dOaSxaIGsEuHEpj5yHjNZmZDiEGO6yMXFBzu5D0dbbuWcfQXI+thtqZKJiShHSTD8vc9HTY
m+lerL1NI+T9/ftT9ozZIu1+diXdakLmNqSD+BJjU+dqTjOsrOmnySxpyh1KTgXS0HFWAoWuFq4J
CveTVgOT5oncbRlPeQeaL/pYm1PIRPtJMFaEVzW7XlMpRpV2gUJZcik/e+opxClPxUXgTVxhAaoz
eT88FW9sHbKge+dVhjcG4EMqWYdRFWIkA5NaTA3nEsyxlCzurkT7fejnrjvO69aXrKcdy72tE65+
43tht5xWcvAR7Ocp2AjknFuqQ3587sTe4tB/wAIy1T8gxyDJanxmPKiDfjgzrPL0gdCoOCFThhKk
nlPRmvhOqPLjSu9LU0U15sBOdATOLbjJfzf8ZaDdRF6j3jOi4tyzVOVwPPeXoQUoDWglmkXRUb4Z
5ooaaEjDsw1f9jVh4eDkjKeGXRNas/lhBgUxxYjUeVzs40rdMdLSyVue6YoExWm/S96YGMqWTKjI
msEV887U6dX74GCSTDmtF2LgX7TFOLKP6lgS+WXC84JyC6TbXG5bl6APts6vVaBz0Ju9ARw1Ciyc
xfRbTktjiDnIz1/Sp8c5XqruwEXgpbR9EyOBq3yFu+y2K36zgdjbns62IuCQGfMq57DnWwAVNJwh
SoiBDCKqvK96/WoTpQ68JJgdptjjSvwAYV4YkP3NSPRWPBNwfrUyT31FZRA/A4K7YKdpYNs8xHbP
Wx2AuPY91WhdWCKoAADJoLBop/CTNbt2CC3h/Aw7bSsFkWXHwtaZPorM4eu0w0PhJAhexGVlDTd1
q6IG/KOjc/au7ft28TrR+kmZV7W3nTynFWNpME/UI5wZz62d/Rn4MRLQ/6bb3i6/lbfdDgmsijrW
e3NME+0TPqRMQ444YNE/2n56koR8NT3zKobhkjPFukAd9zK944vPjC2zmjOaipWQfk5dAfCKOV8s
iOOXeesG6INdSx0iRjVgSQXXBKGPbOuiivNMAzg3HrVd2IwHFbSGEmi+a9Q6kShD157Vfe4Oymw9
oK2Q093TyZZygrc10Ztb963OCu4RzItKZYFolIiu9+XSmipVY5QOUE9vhOgNE/jSrHCPkaYDUIl0
M2Fy3j7c+eZ/Qtz3RmOYE2afcz+YQh37duv24wVXFrxQyvzNUfp7eiDUwkU6O0S8myuQp7nKtirL
V1FbejQbw54v8m5KJEXIsrHoUoF42kLYlLtpOsKFqnSnZJfy+/B52GaXm9lblY3JDHfxE4JUXAJ8
PoYfEZiQUp5bIctL5+o+hv0iwoioPBYzYKHf7VmTKDKYbQPEirYHyuvbw8Ti7txBb0Inxo9EzGry
55e/emTQUd6FfJcmMimSLeieLprWjjO4bufzYfGBmJM2W0tUyhOa7ADm1afnFkmxxsOw48oaJ/Jr
5VS6B6BGTRvqFV2HjQkP2MZE5enUL9NUtjiQt9OyjrZibgivod+JDTwS6NgKf+hQ8ijMwRkKrigU
FaUB35TogrZFJOAfB2OCzt0tal19yEAsHC0FW+e8QfYg22I9tBuvsEF3S9PkOo7deLqK6vA/GgjO
UxUilMUVVSzXvxoD/vVS7WgFgTngS1whg8yII5Gl6dMMB16z9A5zIaxgOLTDCkjgtR+mwmvPTwFm
i28pnoPxgzrfeSd8ANk/49gIM5OPL1VWUsnYVdkJrIEZjfHI02F+Sp8MMhFwRr7z+fzke0PHi55t
UZSoBBgjnJiJnsOZuqxAugzGEjFZ9G7MVH0A7e3MJjs9VrFPzQNfRBGmiWsW6RfWR9EtUleOz1gr
rVXScJTDzo+PgC5V0hlLdKSD1bX09ykpjoAQJgBUMT+hVG1bP/zvHVvMusUt5SJ+uc5MyciMXklT
bxpmJOFfQEfMlcfZUWAsMXJBQkzfUMTtNOv2
`protect end_protected
