`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
vo2QwP5IX+TSD3XsuXZ6evZCOjAojOM3P3cDbl9x/9MWqMiTaqNobcJ57cwPQj/+DuAXszHTwuyR
DMDrOsinXL0/5ltnYZG5XbXZbnAfp5Xh7Vp0Ym54/V9NnPZCNw86e5hMq6oyfVIVA6Ly12wYFcuR
WCzcFWBBLZ6ASkUP+5LlOXzBPcJ/La6t+lK7VqoSbTgTt9JlzlNwsSgcLGGT+AINGYnmGXknqFgE
H1Wyp3e8JKSlPvJH1B4siuR4ijvE5FTwlbRd8SZLlQSKjfJBiMLF3wpuat20E+gl/tnsdiHmxdZb
fVG24/DAxQ5o4999Db08+iPRxQi8QM/YJdhqKQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="broWGfP5sUtZu2OHA5ce+pPKPR25Vke/Us/f/rKv3B8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14880)
`protect data_block
YixsaUDnhFZdy5dJWJWY3Fyzd7CJXtMh2uF7UMLmNH/2eIHua9Vv4rmij+r/ORfiylfayFGv2Hf7
g5kTledW25rOKIKXuM1Acqodnf/SrZ9JbRbCQJPjsIqnCOnupNWrWU/bA/nx1OE1bcJ1ax+csdLA
juxBfFyAGrAohE3VHm0acGVpQ5U/cvrIYJ6IKFJKuYbjAk3a/KtFoFWqB3vA5mfyVzrdgRAybz3t
G7pKaveKNovyMaRjWld3nECBMpbc+hHjRmfIL/EU18LeUyEf+OQB8KTpRWtFPrvO5UW59a0ul6Oj
F1+TNh/89Lrikw3AeeNkoEOqxRMuSNqbSk81r+8SxZ1z5NpqPTTikvNG7UQmgOnuoUe/odtWMhGC
1fX4gDUguzy+BRA+Jt49H338ctY3AkSOHW5WjXWtsyvSdVLHBBJMFsCiUMoaNjMkKE34DWPI//6N
d4KsUazG4PtGAkV6uktlw9gbQ3aFMKstFk/7LvHM7Q1PVfz/bKF9f0NXkobGlsijEI6e0aRk66yz
5TgzGt1f7tApwyifbQyjT0sMykm8DclFsszLqiBJz235OXz687BM+YAtROWW4SRARcZbyQIDsgZx
jPTFivdXTAZFU63fiyuDf6xLGhzlFcNBPWuRyY3bcoJuP0N+4J68QqzOvfpH7s8N/ZdwKQbmJJzV
q03WJtt3GcKaMZRXvEzBOr9EBEjfY/PoGo/uRktvZuf9fWTxPHElGMe7fQgEX9LOZD/WdDkvOtLT
dSs89vQSQ8ppb71SofkNIF8mSDZAxlYbG0kr3MHrGaauch/v7nVKpr+MPZNON4hRK5Hg0qvtrJd2
qrsUY06ER+8aq3AMzWwsPUftGZsfk9SfxrUwTbywESwrcXsTYJB5UzluRzCf4LP7oQ4cOI3JW8MK
PGi7PSrL6cbkZGytCATfQPhh+dgMBfwE7f+gUu5pbVynmeLX9ypg8qfQMjSXvSz7OiF4nza52EIx
vj3sCwscN8BWA5dib6xbbALzndyZ2zFr4pJ2Fho2SFvfCx43df/AJgARiLN9ZHNeFNVYTJhXIccF
sNGreL1Xib+6U16M3l7mUWIJEIXZ+s1Dw5p9ZYpPnsPBn75/pYyiOfFzG9csV2Rn6o8LQnDjk9Ko
yLSCrcaFm7Rbg0QYt/Y/zn/5tVl1DWRv8hpNZC1xmcbjqkql3R4CUAsLUZpyAMNJkSoE45gwIFje
ZgOZfZ5VHNWErjD/2dapSpYxaIeTcWIkegaRmlSliinwZiQ4zgfi2oV+jr2W6cPeOgQK5Se0yq3I
rrk/Nz8UuSQIb9M27JmsqgFYgPzGUCLDTB4Ss9gUHaegqEudHtrZx8b/1g1Rk+dfWerIj3y5k4oK
SER0q23zHfwu5K+9+z/QEbSMrGoNuBNy/QbhNc9LbR2IxNiBW1Idb2eM1t3pnugI/4D1hJsRPS3s
EB51ae9Tiw70cRuHtMc5OeyNtaaqSS/NICKXscFKQm7Zhg/tbqL8x5xqQfYDzzb8kw4aOb81gYDP
THqVAjuKNJJrLj3My/laNecKXWDN5ew6M47LpRL+0frBOObCJkY9NtU0EvYV6On3n/i4onFF5fsy
ElImuGPA0K374YQTUtYGQVSynH57PVtiNt77T50iBI9KrlknvOD9j5Qk6KKSVXaZcvp6+UinW5WF
1x74GG+wUNVp6E/aHHVfYfN2eNPiRSIHQqB6Z1U9BbCrpNkEU5kWrSDs2uHTvOTgVTSuzORHKKRT
9urp2fRIy8e4USGZyLRqUiW5Gl6hjM31vd6je0CwTjb6P0fDvC1NfTt0glnrtbcYB+5L5yHY3Mn3
NfW5GFzMRI4efnxfaxh4tL1NtfehP4YCDOJsw+D9hmqcvwtiClFKTtcprAbhC23lMSOPMB8vhhbY
imsaPJatT7JrhJ2QsBgRHO31A1cIRSxPMRBPuGOyQsbhYDkaapCkw72CUiGtWsFGvWinYmzy75x/
Bw1PBHNePd/25+2wO73vPj9zmg9JVS7tCCAmKSed5ge2USA1SfiTHn5cKCwrpGQVFN+YVIJHqlyr
zYIeYBFH9kjWV1zh+CNLZhFxxt8nNGZaR1EeII0Xuj1tWJL6Tgj32jVSrtdhOPyyNwoQ2mJ2Y6eM
YcLLjflSP1K7mqPizckHZGLux66dPlImUwQBcwWyjAJA0HxpaS5FRk1VVRrD9U79xbQut0UlSW6A
6agHYAwR0TzrYFitEhSry/HosYE1OWd4eBNfBWC0uMYuEeT7jbLx+nlNqcRR7vR0iqf6TIXd64bo
c/6TIVpCoRiUGInyEaoCEi46u5SMxKPq6xWeDCRl4RB2kPOwbRfHkcF9mayzpjfyTyco7YuFKUv6
W4Q9MUauGe8cxFKYDywO1UQFpgFjVl2j/eYqzHf+y4ARtmMNVZMz42LUbU9Cq1X11HzA1elq9SVh
WK0DlGdZVU1xfP5zIQr5tX2zPFu9f/6recW4GUSWbhc3hr9k5aURWqoZOV9JsQs6igPH+a3BplBA
CK8BQYNoUDBwP7ITXutD0xgQXFt6jM3XcqXXtL/JqpbTfiPGXZPxQTI0P9VC0cWWejwcuKW+Xs5n
xU0F3QIpvtzCaRCRdcp6h1xZG0I/9FkujnI7G9cIZ7XypWD+0Snl4z8h12dKCJMAWMjiTkqmbR07
SugSSotMVviSU8X7RELOr6x73vHqQTWMv9uzmWxq2XWzjBgvneKzqhXM59lvvTOc+geqm6Ey7Xw7
Et1ktNJRNWG91gWGK+BBunEc3KyRvIPQlDf4uRghraIZR6lAYQWMAYkQ6Dw1c3Lbi+bzDTRSWa17
7nK4YsVmyL7435H27n6RJprvGluqqkuxwrokES43VuV8y5Oj5l72lCCvExfnugyr4gHaDBuXQn+s
+AeMT1X1Q0giMryIAbm0nIVM80LfkF4MSwCPPDklryN7apRaccNXBYLwYJKBvdYgvTQAhg+YfwIY
BOhX0DSOWyYcrhbXSsPpkc3wwBd/zTH1UpFwqv2rchU6xorlb2wNFKTpabJXevTcSetylMFVPCj9
il+s9kndNuYmQFznjI12nJUVO0XdB9/3JGJW/jE5+JxZbOXWaCj+JFycoNILX1CODjdtaY6CLuzC
B0I1W/suwKFy0dX0zxaAxyFXYd8Pavk6zHUD663bLTipPnvAUhi6TPLbXgd972EBeRNmR+BakP35
EvCPSdYQkrHNiygQTKPi+ivUALACg+w2yrA0IePAourOs6dpIFYBlJuv25P1R3IMCfL6/sUkbOZk
foG+SWR5kqYAwhCl3YWcoycGQVpepz5imMtMeuObhnPJb0z7R/WnGin/7Rl0Mq+zeqpRnpQDIY8U
ZHjrbvVSVxsa6BBc9BgDXv/qMdTzWy2/pPP+RyXBBdtY0AMxmstkZXA6ZXeqGFNmWzHo3evIyJE0
MpKSEXy3/iQbcxjUUSJVpCN6HEhIsKhZUtwruJUw4rEn+Lrod8nY2KM2T88WlzV2DD98UW1U16aE
eBe1ubsakIRXGDRpyVCuNNtW5rBkjnwJGn4yiHoi12aAngMbWclsYbvIMHln7U75F8pbNJ+rf8rR
bi+d8Ty8AARJVO4cWzeHVWpRUE7/lmV/GaeA7cxQAQKWT2lk3ipmW7npDosasFNtwXk6uSlv9OQj
rAD6LUYx/XB/aCoPNs0WOk8jj9yo0e1TjDEaMPJV91+va9q4VJwMnm6l7mIFNJ6JjzJCEq4WFZA5
a6CSxytGpb3TA01H3qCp5CZUKcA/Ub+FbcmoUw9sUmgqNvbA5okYunTxHKfEfcFvfIynD7xKIjPi
rgB9avFacUU7swGMSfOdoTEmAW7jGEk3gqCXr6YS5eZri/hYurhyQR4cyBlWziMzqsbnA/gn5YNu
VtcaODjSRoP+gjxwDzp7cDxuhpQAjCGG51TX+zGqYQY4ZZx5HJwesxfgfjg0E5tRb5JVsA3F6mod
m6WPHS60Rq9QQXCegX0l6OYLcmiXrPfGqvY3wLuZogBKN3HDfxGKJmPAY/eqXyF9BvyFP0BUUr/P
FMw+rnCtyDryG9QnMGa+Za8oKksLV2U9bDGuX5Wld2OWv4+dV7iaWYrq87kpAyUoZ2ZCsb/rRlR6
Tp1xt7xcajC8akumtEa1yG86UvxmMROXAL2a2bSoqR6Tlra2bICDjC7/XA/DuislVixGhGZFajpe
Z5yV+qJIJ3yRwF5bccsvbFkVRoA5nc2epjS9Ik/lnvd8DQS+2AWURk4wXE9FZBCr7THQGd1i5vIF
3ciMWmh8F3x1WqEuZsQ73z1MVW7ipN73vTPHm7ZtDoxNFc3aPUCLEA9NFcod7fUgHXmwDYek9m0v
8p6exAmMsrJFKdGnjAHmrTrZsM4CA3QmMKYtXRzMySnNekm5RL4Iag49O4r0ciY8EqMVpUTMt1Fh
RFu2keBVb9oGfkJLGBTtZ1zVRbN3jwdksJojwaAkVd6krjgTjgZ+qqbjWxveJUx5xyedR8vYPcLB
Jg5Gv5OIEo6Zs2nfX/AQrU1r4tuqVTYTUMBovgrt9BPf9XaxpOzglgyI1B5DI9bqliZ7gjBfiBJW
oa92bX9VOcBzSpXnB2R7MaUt+Ek+28nu186PJYKpfpjSXAWy+RNySL3dP4PA0xRjdzpv3+NnMogP
8o6tLHz5rOQdXRgIM0Q/k6+PWdMfEzjJo23AdW5GUDOk8tpowfzS70suRsRlb1Z401xCS+YWN7d2
x5bwNoZuoTq1SChbYtOsYanSMaLiC/pfkNuGz0CboQLDWkW8o7WxWijSV191AYzgztrinLSANacF
gD/FO3x7b1qBKvobMUes876q6p0b7NyvbUJZTWKjiXqrj3vsh6M7NLDwizPgDaAwxLWpc28QFu/y
D5+90mYS1AiREJ63WoJY7Ovd9Phi7KpGDof2ALU7JSNJW5ZYlKV4+UKLLKu6J56VlM1yPFg4LOdq
zAOAyjq7uq8wTqEMCQsxS3DIUnCd208fptePZhS5Wh1d517rKtUNF+FzSCWg8B+yBEArKqZl7G4F
+IAruvhPG3T6D1eZfStBXfL8llt0eyQQeQvVLKoVCIWL0OA7/jtJ350dFc8xzwzEKeIul7BP9eFU
8JZn+GRLzPdsQYzwRtoR0ntQEA1kogyLLeSGfWLGqc8puw5ObLoz1l/YRe4nMSBLfKbfTuZ6RyPL
gvE88jKUtW7hhHZaZCN9l9weY6ISfyioKAUA7ckyAj9ZyO787aD77ujalW8dyuemhavVkcE2+5cp
9ydDpQfEAG4vW47XSEyNfMlBn+JLjiafcvePFeyVmAASHazoj7kpbz1Al7vL6S/WfR8U3eDk/6GP
Og0OhE1T1J3OKKC0/OgXLCjs40Hm8UQSz+iDiNh37yfovK5KS66lAb8CI9+qk4F6rIHNQFdOyj70
LtPgEpg1oddKGSI7ecRgLjqGgxQhKU8+0SrZfbGGXB7fHkLl6GNMgxASob3QK0fSO/GrEhIKIGia
3MohCYc5iTrGPFORj5odnChN01VTF1XRaVg29JdusiiYcmRcH8Yck+vsPObEMRyzKuyfrhfl5eq4
x9CtJovmwDSK+bFhosaU9KITWnqKrEcMBM1hoRDFtcCbqRU3N4W71ZyXsZDB+H0pdIld/b2GzAcX
3m/RhvMP6+TOL+eIidfYwFwMSuh6vd5x5oajSORYAmlDcWvamgjlnDONnkEC3qrlALztumctv6iN
SQjzAPCymVTHG0+rFkuOXz6F/7Q/GweoAobb2qcPFksTilDmhGhRnDn83j6aNuajSfuBPyRoPD7s
nOCd0S8rfxVxWBbq8FNh2ANU08mr3nVa0jyJxFsrfrzvRA5Aq1c8HI0NBU6w6PmLRf052dzdNCZf
7a7l6tMU31diacCo3YcT3kaAafO97vp78ma7zP78OlIhZMqum+TbtKqk2/T5NSqfANIfAiqPfAjv
DpCKhGVE2xnw1UNe1RzPRsv1E3RZaTaILbWe/TW+pic8OFaSZ2ozs/mh8vaxvaL6h2IFgY28GO1w
YvD5tWtxnU+RfuT8GY4iEad9HlsOofIMUob2HWbTQw5D14PwVJruAwSuOzS50TKhHtEZjpNDb9OH
PJ+fK+8b3E3LaEKOJTEy1eP2jk7YxCtR9CNKWrC98RSwqlBItDfg0ORgAWl+tDWs1kTzHCgku9S8
a0NZPbMix5cO4e08Nh0SCe80ntW5eGYRwWlrL2r7V8RUIrFfP8SIm1RmLDdu43Wa2gOGH4kbuKP2
wKZZXzcEXjNFqxgb/YvdheMhk1cEyxeVWOt4ywHCMfuI/6guIG7gPs6Ft6UZwg9XMbln6ujPgCiX
XBtU86sM8T8U4/tontdS95gNUcAKOsutiKxtRVAfncNDqQRogvBmRK/F3SEnMirbU4VCd2AbZcdM
iQl5V3MTxIFjx1WBo7dQZi78gMo9zm1qFC+Ui/Dt5xehR4SW9kCXx2CYy6gK981hS5i+nuTprlCr
bNjqJZFlqc9hMpCe8BXvbij+WTRui2rLzCM9rm3tBW2f1lVF9uSSsAL23C+aI5z04SpZEMaPOtma
2MOuMr2qmUOCDEZEyWfDmtO51jxncaQimwO7MOQq+gtCoDaSFUjEUvsoe5Cn3dazSXqtDe8tgM2y
c2R7jq+CrzIHH3MKi5ggMHwmOohvRd10D2neiHfYuWfpJhudOn5WP3N1LoZKW/+vZWIlbj5FZh/8
V5FETkQnWsG7gJP8Lipi94J6wOBTMLSJnkB4S4USGo/noBAoXJs+H2RXZRf6DnzjTMo4D4J7B9KV
TqWJf+pNuDPTavwLjFCvNVLcQ4UnYSNa1kJ8t9/LFU9Cq6V0zfHf072jgeNR2AZ8WUNW5Laz5NJ5
7m/G06WrfhITCVff9x35XADgmyCBydSDgQBp842g4gQPbeW+ANp3KHfh57rmxnZ7tfeVhefmQn0H
dFZAF2bP4fqqycfq/VDmFT2tr4w5PTG8PeK5G7OA1c2G7WovugNwu4GWZLN/GQptJrEaZGeGT3tf
5jBQxZtUL2uUFQjdmpVC2TmBvsZ4SNJtTRWG+ZbuukIBxiqHEqy7pZ+ZShqYLcoKlaoIILOpr63R
+KIDqOEoSZZVNnehFEq3MYaJ2uLmQx7njFf6V9brLdimJ6DOI2ZGMBsruM+UDuAmxpNvxUYJtOXd
Qxv4W3/VjcMdXrhlp/UUZtLHIaItXEOZIdNdni9nGHM9JKIbTmIX8/UcDyyiJRQdOpvy9oFf3PBw
jVw/7kYgnvDaS2rppAh0khBLfnakeSkrUA1DyopJ1TYCzFzMxdmRUEoEM2/CmbMlkxiQ6DYdebpd
dRVsIDj9dXjgwUtcZitD96imqjmtV5OsdGa80/M+NKUYS5qah3TaNZwTTPM7lg9dMZToS0QI53ni
sD4I2+jwi6MOXrNT9zp2Lc8bNfQR7RYOqIfAGGyFkrbH9DuORC6ArH1K+uDtjl3TAVcNtf36V4o/
LjTdfjYqu8FI1uqMF8Yjaqdo9Rikl+lZKYaNc/eXjJlnvu/D+LT9KP+mkTzIQ7bNoA29isw4ugcd
l5tTa5fQeHN9lKEPZccBCCME9NqoNa/RvfGwj3i28Eqca55mBz5BBe8JSeYCYzw7SlPR6H+xmCvg
UbvmMUIS2hSEDOXf/vIORINRU7u7k2bIyMDjhUpwBSnGKp60akC/Xsu5oGt23RxF/f1FkIX2Gixd
deoXvUFhULSsH2uvUIuw0I0SYsNmLlhByb4ro46Gic529OG4M9+K5Ahk99bCiAOvWZWlCUPtfbkf
BQuu76rDCOU4sIOVcB8ciQPdbxcdjy42qvsO/m4ndlXgodD6kNZs9i80S81CbM9SPSGl5JXnKplX
19vuDJyZGSb88OOsqWxp8i5N/TQE4dQoJQWriB/NwDyb0OQkrfzQVVzT17FhxzvLG49wE7OKVoZD
f75WC+PcSieCmWMGkcXcluEx9aQ4RaEfpaPaiI7XDmQJswoBuDTvJx5Buifm2+f4p3bTVt28tcqN
68mNVNxBckwpf8cORXK4gFcnI+amLt47c/ohjAiKo8WYHX8wAYQJodo6u4lpc3bZVFQO6OMwHPwT
Aq8nN2a213hr8u8Kyxv67yKGh2H/Iejm2qoTc/nvaMfsh7bx0dVJrjGH7fATmmqFhleRPJD0Tow/
BKRSmXG/WPXHe5EYnsoOgy4TRtoo1xNYpecZFVDgwwSpZbO2zPzgFfwEafHpXiOAzpjJuVLOp775
6bfcEfvkrSC47dC8cSk9i2rQZpBdxU5VAXFEH2R/it9DIpm+tOi28lgcWdCBPmQCbhPQpeuNtmaE
uKj5QtdaBrxhaec9xrUcDcftpkeDRocxa2qo619LcfXh9A7mjA5BnHjoJTgnAT2QJpM5Z9yOhcen
QuC+J7+bZuvQz127DbsohfHQzPnGut1mFlIZ8QA75SNvnNSrdQNXb6OdXUs3ijktDWSQ2v1sy5rO
xyGK11GgpPq7b6BG38cQHlJFBHFxvx9FwiQr41vuQFiNBQoX7qwxALEeMrHoQhGwBsDZVPo1X76A
CF1BAJIYQQ8i3TVCD7ANhNTvWfiEgbvr2ihRtEU69gP8z27xYPYpuT07nYnoANP7njF+lfIeAcDs
5Yo+/2txSlX6FItvq1ZNkym3sQ/Y9LsQ7+pPtGNl1+QNJIxX1IzwWcVuGHHbwdTIQt8DaD7TvVLE
QTmnoI9bYQDB+N+g0KtBsRfCP8NIBdXvy4k36QoFI5yNG+oKdkdPQQU2OPbJTYOKwaxJJLLSGbCr
9I0n27SW/GRcs+VTM8EnBVqMM9NvxdcUMYGM4Gfmv0QrxBAQ1NGVxL4R6ozyL/Qn2OXW2Fy9AetJ
ZcQWxs4eiSaWVeHAYkXhGscCNEKv/5CBjCcayGdepauzS5bRSeeb9Xe/AVvcKv0EzmNx+mzSEEAV
xYG71qvMY/wqWpz1SdSHXQcD1Cl9IXZsfSVv2qjKaW4ix+p7V6mXmWmXiVBfvHpBTt37D88PmFjY
T9nibOHeTfbXh8+W+4xCNGQsOx9B2lH5p4KMxmeWiEH338C8nXIVJTOmE4PRf/Emv9hwsBKHFWK5
6gkPpa9kI5o1vZcJikqS5IummdcPIPvdAW9u9ZXFZQrbxwvp4kJvz5ZUHtiBSUmnjPx5oB319tYS
vV3tAQQmagTz8ouvHZ8Ba8fE+cTEVkhwQGJur5Tca7TGiKT2R3G+GbSECbpADsETTdSlz2RPLYCY
4CtUGoM710B2kllQzzVUFGbUiU98GedR9IMMI60DyJMrLJ/qpIqckaHdyhRLhpUcAgSgbJg1J4my
gYJG+Gq9f9LnbZC34cXvJhQGrl3XSSSD1uEmSbYHKuggcPkY96nNwwDDYmgXWd4Ape2vcRQVMPiG
GILDo0HMgWEQFNFmA2fhwjYTXeR5a6MgYIpAurhk9ZakqbavrMT24mZ/4vN92nWeWICqeSBmYJ+H
/mLSsgK9TTK281y78gu7dfea+yaNdAF99TgJN4cz8Cagfta6IyCkqyGTiixmMaNQErxv3fjU/r5V
h6/FJyrESH8Gd39l9FbfN5ztV7zkC3HyyFxXd2JXNiP4ERdlErB1/H6LIDcZqHlJG/feMnTpmEr+
IiXYtizahn4cC4SSQZbA8a1z3KeNpmcRHdJV3yzSsmvq2pLCU8/00kcKcp0dExEcnc+LG1jCQIHb
r1UqXWudmWtTRHI6oNhEM+tVOMx8CvO3J1p7hFCwhcUr0//vI8ifadOuzcaSFjZlmzIfe141jscN
pb4sG6Aa1q2NbgYn4r4fJjVSViugruoNgbLL8Gx3b+8z6+Ps8ZBdp8u48BqenZLiK/5EfhDV0D5B
S0DRK5n/lMYdbblOiEEeH3baD5SjmCliq0mfms53L7WDg9upekxqj2m+HTIGOlf+UpE4ai1P2csV
xy51OKbcWxeZXSx9Eh23o/nIEQ8h95cFgNqX5u+BILBrSTFUXOB5TTMHxZwvpxTjkIIziNrjqxHU
HfDQEmX9cnk62TeEsn/yRz4ZC74YS1wZByGpjfsLZRCZKvKhWVTa8pMYAz9j63Frn56U+8m9ulMi
nuyCSWq7aLX0J95HWOEAqpOXXlbMjj2B1v6bGSDnAOqevAKOZH2sTxXG9CsjWLRV5dt2wncOfhkw
aKpkgL/6j70WzD+NXwVRtexAgvjxjfH/3YWF7iDmGxVaq80VwWLHegtizRIXaPkFHcFnNr/dL+gM
M11e5j4YkE4OmuDhgQYRmqUlM1gLQtrno1BI92aKfXdJFgv6YZITx0+QUuuX3rP0PhkkGqJGiBvV
+fXuiuCXLGkYImMTowNC39OZvEsiny6FgBSWcNdR3xcAQNFnO+n6g7m5/0t9B1IOzmBsgjKAmIJ9
SpeAqfcLsrUSYKNsXwzKtuvWvNJJk8tT/QyOuJmFxA2Kf9UN1Y6j+K25eFvnWWaxxQdOvh8k5HsR
7dAeuD9P9XToWYa2ll0Zf83WYOuhG1cBZc9G8/FOkraoMthi95qm1ZTcBdoOjgjBrRstXFndLDEn
IfJX6N8a9SibODRmLqhrOJTOX3vtbiXAkWE3NPRcwuyDVbPQXnf0guHpU0+T0cZ0uPj1YGf9GIh9
KvSFBk55gjlejEHFAgAti3T+gkX4DCX0o31WCGGUozF3JuPvW3TkckXu8C+E+QqIlUEAdyTbUNwf
I+XppTm32GQPsYIvjP2SB6AVcoyFNDj9ycUJwlUNs0D4p/YdmAsTvXBexq33aWMxVxUo0gQ2tGtf
0TPLG7fWkurgOaIP0r5veJDjbPXZO6sBeG/g9T/ey41Up194qvP8ui0l40+zEcq19EO50hZ8VyV6
7LCGnCwq8I9Atx55wdFh+un3Ui1O2O+RFc6CN3Zdaz0LJ2HMl6H1JXUce4LfChVwteeW2Z5400Ss
StcrRG4LGz52/P0StyR9AGgkaZvnodKIkaLgiFTxN55YcLv71L9ZYe9yecUO/MxTc6iyVPyUj64V
FnuOrHfIxLpDGAMtnE3IA4Q9ts/krIiXauWOTj1dkXGdgpUD6W8lhhUpIo5yda1HaP4zojtXSggB
GX23/9sEPmulJ7lBiVvf1SGdNTSQIhterm5lIGwzdUS/DNE68jRaRZWvETcb4PRH+mNWAvEkSCRo
pS+A+AayyaMp7Sj3f68GYl+0mLdqlZISlEfoOeC7IveU1q1xpP7N64odYqs+1w08CJ0VbDp1cHTm
USLgCrS057lCZK9SQ8S5M4jpTtMkzyZCsfWfaUzhsgFaihjq4q30jpewAXh4Qo41dOT5vbiz4bvR
i84KzZnnsqa9De+1yaKrzZmoMIgsIcFynHorsM/Ujg81aNDMNm+O/vyPQ0ff9CApo2EnESB1Sriv
91hbo1QU2f+qLWNjnhZ/2RLbFMM++5Th0SwvJrdMdaq0/ylTUZyYt86WQJ1yzfJvIFGe6Wh2bHIP
DdbyhlYl4+qgxx99YMR/stL9ij5Cg3oSVBiRSMMnInmg+Zo3Ps8z8Q+4L2YmKolRBlHWXayEv4Zx
3aVV0hejFgk82QsBilB5L8msIMe/QxkM4Li9XtveDfaFVuEoskRFQVXDcsQLScnQXpcCdX7ypcJi
ZG9YAxZ9xXN6BR5xg7hRUTuRpPvOBUIvbbalYPidT3pdyIbI71WoppQ19Y5ByYN3eu3ZodbdF/cJ
4/fWsTNEifVBP5c9gpjvtejbi5ApB3qH7AFYcd+PCJDrHIP8LkiXCZnYh90MCpJ789DOoIkG2cly
TQWwzQGyUNypiGmDMiGKc70UQMyfu1FaxBFgSbwYCGL2MveJfwDAaka3PVEBbeEQyrdTqjMn30gK
gmss5JcxrlhEQVh9+hInZW7OoJoj40Owe6yFC7qdD1EGKFTf0CHnoebtz8RauAccVE1DUK5pbujL
h+bFA8xdNSq+1MbppXbm13kfGGPpeaB7ul5V7etKOP145syTzyVLnKchfgxpIDY+56IP4VwgjmUz
ETNu16pBoxib/wlBQUIn+Ym3Lkl12d9JGG3MRjEYgLcC0xdMssFka1bo9pmsgLWOcHHltxQ5tyUE
8mmjkOG2WMKxkiJNbQiHoUHSX1ELTkhinSdhfTOXfE015jLihXSki1lHfgTIepU9l3DLaeGgm7Xe
fjsIRjmpLPtDWrekKdqMvZgfrOl7PRFRY0yX1hDWpXhrwpIKz+bbP3uUcAmPxZ6bT85ocYZfZ5t7
/JhYe30Z6pnCvqOB2AWSrOmSmzy2HNK7rmlD5xvlWueBRLP8Gouk5OQ+xPCLly7mXY+DVcwXokoK
gwbG0uSYR9r+mt4SfrIZEyC94tzOBCnhVaWPwUMymAKmxj3BL+sFpoI3eV/rox35ESLO5Gpwu05l
z7lC/y2D/V82yb186hY1dZ6PEv1uz3gUaw6oZanfe1sipLM3rdRMiuLUFIvQX165fMhMtH2MBcCH
+FkKJ/hm8T6RHjVrePSKKPdX62RSRrW7qGqYWvkRGfpiyp8zel+pdbGSyZlQLaTvhbacB5GFWo6v
ggJFkdSGhswCxnElIqW6EedMhxp5PkIkT/A/EFe50+RKCsDZPZQD4piA8SFMpdAboUuQBnOc2Lw0
e/d3nbU3sWFYuE8uVmUCsj/wt9y50mssaxHrV8XNPyTQbCTPnMMscmDpv2j0QayMOLJnuQDEsjBg
9mpFKvAHAaivo2B6QQCm+RunEH28dZUb/au7/GzSsoV7X3tNvu1A0IcgpwjsOgRNK6ZamNig+5O3
UmvGZ0r9lOSZNBSPPyLUlkBIiElYhhBSAS/iX/igTgC9RgX9RMCejurf9DOH7sTKf01vJdLrpR8W
sYI5FCu083BhOouk/Zq831IkfvCNPw4lpZwaH/z3txtkl3O8TXrO0OrmZ10IBZRPSexmKPJ1TRJz
7Z4igQO6NTmAy17RhX6u0HojPB/f/eCbwKVQmQ1OKO3qeRM16I8s7gsclXeCJbxOwGyIwvw46Zmk
m0rnHtZcMjbzVJ+vi+ZiuCKZpB6wr/+uIfjdNA3IaAJ5R7yk34cQ0rOCspOuz4DmwoGp5ixGw867
8vL/TOdP4h+/fumwaglEnAne+gE2Fx/00XUMvoaks/fsj1IypIjleZ46WW4ROfP2EvowYEwq2RNT
H+18rfyJURUhBPxmvUDlOKNTXiVjRjmoSO9UdbSulvmxYeWu6749E5Uc1K4rSA8ox2L4/y4YWRkT
x9qDH45FzdIEue8/JsBTw6xf0C4qvBvmUyuSQ5AzndgLC9c9x7JPytLYWt2qf9wDHUhLJ37sjH3q
pXlVD0TWqJmMfGneNbKHVyJU7aR2xjQ5m0s7WaVsfohg+5InYedTShfbiIxX6HPfXTk/S4uMx9Us
B5aocCVlrksoFVijT0dSwhfijfasRYDPL+DEZ01A5l0UJfNN178jM1VPe4UAG87/AwQ0k9+RtMFN
toqdgHYOE701NF7UOZz56eLYerESe27pQsE8hx+7ov+fs5txPTxmViN8fFZezbYxan+ue8nAdCvZ
wOgTT0Yxub48qxv1UKstGzvd/Nffgs1v2WcGM9ek1QDQWDM0G3gyAv+7B/n/ApPpJtoJvyaSNPlK
uALdBLAMIw0OjlBPbxrhcEO3KEEJ6gxG8H03hQB2L6TvEYoKEAGyeQT3ic+K9E80vJR9jSoB2kuj
MYxSFkVFiYuQaaWK7x0rbhg1bnMo+v/clAipFZcABFeUkLITw50clkub/c+lOOtI0qL6U7mU1dLw
EcsVJeP//uTTz2t9gDtwQVXb+BFheFqRm28abAqlZTQ3j91GLQnXuUbeOSNbKRbwr20v3Brnozfo
Ejp4gtjfTvo9pAUmGlWGSZFpqPa2WAGdFnctlBybWFrHYuhNZQfHeJZIZystVlwq32asUmaMN4dG
BY9Hk7fVTDTBHr65FU2mRr0EmViKKat01F/AkBrDyPpgdFREptkm7sUv+afZ8CaoPqVsOkNg6/in
LJ+VLM6I6QrsbKNlzTWB06nQnWs0RCaltWE3SMX/62DH3GnzZ1wPe69p/jjlHSqe6PGi0ZA04K1f
JKxxMcADb/9dsF9qNDZVfBrx7SkAw1HMFjHBPBipcO2AUXVVVTjgP6TnCafko7FCI0kEtX4hScg6
5qWlOA8CAQj+LrVftZmXaPzHiZrKOnwi/PNyGBiucc6DpXo3TuAxmTYH8MbuPRSgd+38uc83JSSQ
hDxQ567RuWUlu5W3A20BpoM3wSZ94E4azlg15Z9BTovIs3IVCqaqf9hzdD0vBLBAc0YErvUTz9hg
qsR4SlH/2apG6PDkOIkZMUV529ooQ6GXghlwxfEEHxu3omsSAzyweXBVTgFBrH86n6c3xtRU2vyU
RoQ43VZiCun9XUekK5DlIZsRvhNIMKQ4S+aOw82ONuxsFusu1LLpMfnKpT75euk2DtjexvbYquFs
vj4EPdxVs8/W9JvnJT26b3EUKYrkRUftW18mjP4HzwKe9xhVkuhuSgGFs9TBY1LeCnZUgS7QRLfr
gEP8pvTsIDxikkNr0/4eihpWW6mMcNDkabtyG6w1gp9YvN+KTFH9++SzCSGCl5LQlJLiPND4QemI
+ZPRQbdQ//M4FRnjb3tuolDULie8/T+RqUlMGUWjhPkOijCdVouIa3NjEtkply09WsYKsY571uNa
hT5qFTkj3vFnnpxU0FT4fxY7b8xvOpLcs46ItfRE84H50Noh4gm36RF19eQH3z6scZ4M2nGZajFY
qD+nXcbY8Nj9pPDqXfkvPaA4mIbDrr8hUmtpQTVARJDuYQuV7ieioEEyVoCov17bW7e0Yku226WV
5+Gi9jEqgRhYe2QC5V6pP2xlME/ci9Q9GeeaU/o0mBOUqAFrWa32N8jbU4/5/69T0zEUGtLbrkIN
LHPyGsBrXElqt1/aa4xaGqR15DOnNHvHguKmw3gt4M/bqg/GGsQUTLl5eSIPA6Qi72kwGpdRI+LJ
hkUmHqUDmjvhg1CJ5/TZ56TEacYCpMVLb5pOGM3kfEwPl3iDOKPBxktfLNEFzMoF3QZ+ZLRz8mAY
jok65OAo7L74TplcPN0//tEMq///5vYfHivYHglIkcyoSilScKn+/w17/4VFGAy9llmXQ+CeaxxZ
C38K8ll9cuTXZjzdeT9VU90yUBu3BXBCC5BUpsda1PWsXwX7ruasNbIxq9LmVtVxkwkt0kb93JGy
XjuwaVR+iSGDq6GQ6uwKF+4anl8v7cr3lB2hGvb6ozjeLFlYv/MjNNFO+Z7nHu1TkDTURzZ7eLa5
rmMplSbOAVg+hPdk5ePK6f7jbU0+GPymKNSfaafc/mYdbC4FDA8xYFj+cVAYDSr9lW5kCCqHm8sj
WqJyRamll34wPNZZARdxUt9PhBEo79uasVioC6Tr61+PC9p/YtcCMwVAVxzPQbEUCaQdId0WSns9
+w8KkC809y6aKxYH6YwpNwW1PIHT2DFzpTs9sDnoNuBBL/yJkvPhml72m10oPCQ3Hz9bpfwEkm/2
+SwAjY6aARbhdHH1BIASVWdaOFL9M1NKdD6mMHE0L+W3k9ZxZx+yNXxOaayRjrMSu2AlusuTc1PB
b6dRgRaKCHmTqznf7sxek+vhtTLEpfKAF9ZijexlLbquzLmez/axi6KUpkYegp2y6o5B0HysgoLX
8snrTque1IPSCG4aoZ+aDP4j5ptwtzSs8w1rSo7JnVXHeJDF9xQ3OCW/j8T3vyDoU4c+ViJpDsno
iiUM6MyJxJpKpBh6bQvMF4pK7z0rrNgU75d1ug07Vbw17YAeyjxompZsVJ4p5GMsffkxtwScP/t/
I+v0JGUe6y6aAczynijkUxIhn+ftIRLhjhj/lPIVDk769Tcl26sTXXRM/ZOrD6krv2Jj2V4v+13q
CbwUH5NXAjdgyHT4/grEmpF4YVQzRuI6FK3TJhhtWQLmcmj0/SfmaUywEQqvm8GEHIs3GRjKfJvR
UDUF1x2rB7gCByn/3Tdb8IvIEOEKV2VqxsZU6DxhqX72lAZEpijYOGGnpYlBapiZrtXXHx8D4fpV
hOK+HtIXcjZzXa0SGpmcrWirNNKTsOl38bwoD5+LqLvUQtCYGQmAt56BKl1Yp34OI6tDExGtYG2c
wIVkaNRiibPVOivOXVGe6cX+qYxcX7ga6VPKS4g/Pp5N0TPBqoi+x+cneRdT0vcZvWyu+hyz7fl2
xBnty4C8nhdVtxxVMHeuWD6h0D1doFBfsFcOyRslCKrTf1Rw3vG27VY5m5WQEgDJ2Ok0o9WVmCES
d/T5YXtpEUTdaQWMSUE0HSagXt7a9Rz4Gnn57Jq5bl3T2URqZVljd2I/HEuvI3GzIS5nIqZJtkdl
Q2mdoUKMMsU4uy/WrFeHh2HuYGgQB5WwGkzrsRjS3vIdp2eNo0sX2iBTUXqVCi8f7c156uozcLsw
jis/pKcUzTY08IAaNhisliN3f0NZrvSj0F1mWNyEnZJ9B1wBafbXXZ93w2ftNUQb4WwVo6aqQLUh
oXyEGlGzHMZ1IN+/hAD1Vps339MJU5OrD97wzeZ+3/qx1uEq5tSGgx3dhDyfAD3M38DfslCYj6Xs
ykAcI0HiwbDw6fMZkfoJ67/5/5Y3c3t/jl+wOg3Go2japMKCcLiqvSWx2up/QtY4tw5Bz0QN05nP
OdCg6Xh3esw+F/lIkX62iBXZGXvImRO3bBbkBB/6i/P6JgNYR6lz99vNmrb48D5IacOPPP14clLF
cJcjeF/X7BPwMDnQEkFJPwobCgbiYTYSaC/CTyVIUMnpcgKZuke4zqBzjwiFTUh1eB1pAwBBvnly
qpgw6yTINAajdxHXmOVlyhtnJhJNfn4GG6MVGL2mhZtr08A0UMC1Du9Zw38JQp/4p6FUo7fMFgz6
mstnMeia/ipryMlXUEF6SKZrBDhc+VtS5KdDO6XPXCOVcYKddkADjVBIYZ5+PW8OAHTT0sMZxunY
3uxb1Rs6nCYmE8GwhrykuohFKhwjAL8zWwl3ZQvvRZhBtMtvzAbISJ7Exr08QXBpq6ZsfzizRph2
O6W9xLO+BrG5ET4i2CzYxKNJ0035pDsOOodEkQVGBDkTjZgWYnpogmo/dFrgREiKjDKNnXQX9Pkv
Nr1zbfjuIFkbeBxPqEkVPQlgxCSRfNp4hGXTjMpqQY8+xQFmPeNKzNN5rTgHY+vxOq+/BsR8bAt4
Q1Sr+G9AU0g4epI3As82tvJ15JViaGgva+q0EUKMXg4iNCERVXlDQ8HKK2d4KEDEcLYmxsKPBrod
uNCTRkOi9RMf1F51wES5wy6IpG6LsPp6fQJ9Da02G4ecz4A4zO5tqG//z7u5HcEvpPQb9ZpX3/lK
bv1YoDu1kW/Iehgp8RincE+wxUwDQaoccCKUjXAuuz4yTk8RS0Tmi83drSLSBPMQoGww6uxKCdSP
0+jgQWSzBho47PzFHZj2gC9MR/Yd4JoMfvP+N7PIwP9QrppikADZgh/PK4c1BRw/4MWl+jI1pK2p
Hr6ap4O+wymQ2RS3LEI2wd5KURlF8/gzMJJjqSs/XZT0vsO+yJekkJJiTFMUYYjhYZ0N7K2ppG06
sj2cW3I5aJwHEuuM+QEntwnuGV4mESMkm8PTFm+76wVCOK8ZVQPkzAJF95Rfl368j9crU0Kcl4AH
+t7cxCnJGIZCW+0AAy+h7IqvNteAP/4syc63M/BR3mPxAbHkQRtyBoRAHJd4kskz1Z+Zs3iJGEn1
2Z+9jylp+adB60MSvHy6nUjIFb1WLO3IgFHwYb+bWjO5pH3b5DOGY+qRjmE+goY7sDVKvtwJU3VV
+LswLWlCLCYxzD7HuTdgnOTKxuAqwIZR2Jzn5o9qpuGnS93XmKT4KQlfwoFbbFKKszTAGTWrLAZI
orf4fycT5LLk1dVTGuGXV8qC/NOAuorqivo5Vqb6mPFXSN8unk1dQccDZbDMFj2CbZ9KtgsUwCen
IuvbLRAN8I5QqHDQCr2frT9tRRi0XwKPZnc47IbITRieEFSUbqeIaWBCH3sn/YhR1n3t2C4IR7pV
NzTjV7rQKkTW7DFCICHe4sgtSEgqFK3uzI2eJgst6FjkEZFQCK7HeiHyPYL7ib2/qKRXwSzOgXV7
8q/HJxZOdcfBt+I7kAZk3JG3GbriTftg+TAStQCGckUjvBovT5QqsDLL0NS+gAB5/meYJ3zUgu7a
/EQG5pJRuR2UYmrTGQxurpbhEn6XbzmqRQq3Skl2TJ+JSfL4jcHIGrUusn52nqwB++sUceOQN6fY
amxCGm+5ZPEvW6q5Q+d3/TsfJZcg4rFS9HmnCm69fRKdgX5ywjtVKehhOil+qQM2GpNkM3/PYTV2
qBcYrH9EqIGtDnBXaUXtdyvkCsjugSFsABpowIdYtraONYgp8r7/o1q01q2gHCgV5cWoF2LdgtzM
UL3erVxfg7fZYCqLWKvmzV2P0ASZv8yhEIMZk1B1YHWoQXjTqI4X3xfZgZ8gprI0+yXxtN/Wb5mh
zw8Jz04rQTrpe7EnWqEIv6vyvHpdIbAAjFy0CVy5F6MwjFbm4R0EdY9aYXo+nGCyyhzaUE2oPRBQ
9EC9Wc7avkAVPhJFln4RlNpbLgtbAIHXFEEgtPjCjTDi7XhtBdfZ1gRi/VC1X4o+t5PUi+faKxfK
wWOfCDiUHEZF2UOaXvwR02FPaqSlpPYytBQKqzNF9m+/gCFqYq//AJrBhyDcQ6UaVgbzwbm5DzIY
Azubf9O066bZmmKWmByOlv+kqOM/czcv7/+DqnDQIFgbwYTigZnzopMmv6vtdmnFaNkfDNj6PRal
ep9rDlE/Gv7sjp37N8XwGpNA/7AEQEQUBZR2ha/wTKaMvfjhIGPcQzQixAKVhlUcoLuyFXcLh1ke
HEyfeeymPqfV2h3cxdz/IG6wRAhfQqnVFO9QOWI3LnVQKjbdYbj+d7AcM/fsQ22kffLAvlPIjUjG
CcXIEScbHIq378UD6tIen9xtT69LLzYjYIG/8gc6qRhdSQmutsxikWDOw1JDGNWmnXm0Bygnb+xU
inUu3e5mVfPUGITD6D8wBNIgZQgMWSBWj61VlYDvHKvwQIDqO6KfIMEWOmCWlgBdItZl0vDtEjH4
FwzvDn6fYMScjBjnKOfTzJfrlfli+tv0iUaMRtZfy+NUa3wzH245+yn274nxqTKpBPZAT+qG6UIq
dQXERAz1QE2dQwL9hVt6zd8zCWFOXkCVyT5WUdjOC86H5Eu81PWL/ED6I0MpMUaU04QgE/TuUiCr
U7YkivfGCkqWDHGuFvZrs1fnoCW8KhzDIi1OdGD5h5uiFLy6GCipvKvSiUM3bARuFiy0YLjjanR7
PQyC6UMj/xtUHOTUmT2HmxoNYuXNL0DDeOaVzaz51EHxUlHIAZxrZEZIEFJjvj6kPcn6cKXBsYq6
DH2eoPan/4v7R6kN9mIRB1EEcOkG2UL89mVpttwD/FO9AuJpisSxPBsAS9fFIRhZoaJI6wkXOJmX
ImLAp6CKjbFyc/ebMmFLxcRsyJbmbN3impExe+838T51DsbEdmGFYzhsUUCvgzKvi5AXmqvNMJce
PSYGR+kPfe7MGvmB+6NUNd7Rt8INWLCrs/r5u32G6AErGT/vIxYdfRGb1ng8v4j+w2T0QOjKd0uO
RxsDA1Ev7gQb/m63D44jpyMBQMyjet2qEUR6Emt9caYf8F/RHnpcwmfpsHGEpe6+V7Bt76MUDssX
y542REdKBL5auT+cixO8v4PIu/zEIhHoHQ9tm3il9F3TXpssifbmgidFEBML1n6l5hlkQLGghXhK
2C6nfTStAyrnCvvHR8DGRE3QQB5coNTnEu8B97v+6xpWkVcvBKS+dB3ztsmLRXTXI8DTJuoH4Xbv
oMJJ9NRaiGh5YpEvVyahf9XZ9ypqPZPEqemd6IYGmffO8DP60m7SgNzcUULlRh81zyvZ+gP/mr46
DbBx
`protect end_protected
