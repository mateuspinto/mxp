`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
J5Dx6YxJZaGXJY1e25H8YS7m70iYMaV4XVbAFYNagGfiCkCer5agKOfHxfe8Jkm6Evju5x5bDASE
g6W0fvljiGevmoWVM142ME5BJz0RTwp7ODWCMvjYM8pnvsdERio2ZjEeU2eqKZNOVHNK3/QOD/+M
ttjU7JpEB/kjZwdnaAuJLY0Gzwz7dCiQkIW3+x6Gmlax4nNG++eieZG3LJ5b6NqrP8RdTm8v4/ib
cKJqIShk5gGduAo7MABjcLfq4/+EdCx7xwR8cV8XB02PaVKqamMEfBTMMjNM9jS7LGqkBsh+Xu4g
yHkVNRc5ehMeAtaRcRdimcHGkAQtEHx9872IUA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="2kfM743dNqtZ2jTuz6AVgc+DXX+yG3A7RsNDkwABi9w="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7232)
`protect data_block
ieL9GlAU1S1VhFSabKRro5IGurQOklRyWDBKPWugGnX1OWasbxdwVrid1yzmNWsxHak4+viB/zPs
oLpcTAWp0UlZRJFkagOFkWgc1zDfI5TxSffvpJBHXKEENXQmb9BtKw0GndwD03Kfk2FZgImJBj4D
TuwqLBMC87NuQ68/PYCwKX5ZC21D6qxGCC1OaIwB3C3kVliWH5b6zZGE1RnY3l1ajVyvbN6bsMzv
31vPRTKjQ/FrpS39JTnYp/llbcgfWNEoCBGEoboN4Fg9bzchrsKQwu6/KGvnyxOj9r4kOC9it7AA
ys/ovufVdC1iR2AucnAARVIm/BRXHqo0/7gwg4sGkPcLp2Wqn3UJ4GbOvKjfCvlGLrFw2Ui2gWAk
FqBgbclV/koiDYYH+8Do7SZBVpx2fOkaIxwVnZT0zhSabcfe9bLNixFMvmRP42pzskevAkzG+PFy
gA5OjCFY3SiQm+1cfO5/YyJvwvATQauT3Jsmk69OqoO6Q2AaPQTozouVkGElz7rFh6Oa/BtA8xqZ
ggIgjYSLHvWVC+aM8ATjstHNQ2cRrm8QkaGrvptWJwELbsRrKCyn5j7ws4zxcRRjnCLeIBqxS3f2
rnG2WOx7IviEedPSOZ9rn68R0Ne/LMR8WMA0Iy13vgCtWwDCJ9/qAhnQX4orny+3xWet379AcK+b
cpOsn7Q1m0NnvVYKQF/ovzNwH2quCNvfT5aXALqLYSMxCWPO0EVCbHm+34oeBNY/mHK/MqlGh2tq
/7payov2OPeI5gybTrX0bOUF8CLaHAv2JJVmGLClFM2PpCMP/hVcqp0JDiRC3aFpnYTijsC6Jc62
DipfYbak++jE+e30CnBbGXlBnqPB2JuetnQOq+93ueE/zmysHc6CpjiR44gF1hKAobYkjhzQ/WhL
ZsPrtrR9FZef+KUDnpa0pZokEeOuxYoa7zRvnLEVwxbbee1CL/muN/1IkiSM5JYaBhl8edWYZYqG
YFzKoXEbfOlJnglCaw8FuBdULA3rIkcizVNHEOE/lQ8fBixk9XPqNLGwj3eYs1BXrAAsfpk8Uy6w
BFk3pQyw2M1DbyYSX9rRdYlKFlNzcS4ymIx+SJ9HYtP41+L1sVLaKAF/SiGQB5/uq1eIKvGG/Y+Z
orLREcnYVDT22XAK0J/nx3++OLfpd73GPbVut7QIRHIoJnlpZn+Vr//tw0MQjebEExyG+t7pQh0S
lY1VffTOiEqbyXqtsg5lfwgG6cAPO1xC0qdV3Tgj1pap2VHuPoC5BrDI78myNX2OcKq4MF09uliN
0BXhjljXX2oXuQK00Um+QxAmd2xRLPlIJrfSm1bo/1PCRYqEL64871J96jvPUimN7m8lg0XpXUzL
j8SpLQdlpdORiLxGHqSP6iyaejYdO74g0EO+LpLZZrQHQmeDWoH8Rg+hnqW3coqDdFQkduWIlOLf
fuANvMqaCoNpTOp9DbmLIfcNC2FAuOKTXhK4Mj5WftaCq29XACgrnazHwoGu5GDWnAh9O/sijils
YuxTG0jd6CgiZaHwNnBGBeS3UHIGthHgjssGEdOwochxW+LgAarNbHPZws1fOUj2oD+Fxg5y7Kvz
6MQ6VDjG6q7zI2GFrFpV1VgTnbaMR6SgX/0ODdGmzsPEAY/rUjb9NB3CfD+Z9jYN06KGqfyybsTn
lqwIo/Qzdf2BkfQf1nFFWJChyUqPqiX9HbkevPzTh4BofHs/45nnGxoqROaXB2tm1pbSKfSMIiSG
j3iWr5iz8rqFgXGLDkGlMn/JOO2kpjqNTg3sTQg4EuoCJl13mCwmmetkigtUd4XWwxMlHzKHGcDY
GSkgvWtYCFhWlK34CNWAxstXCtmdaYZKMs1WmTcHyoQRz6yx+UbL6J+w8dxKW6uejjL/OvFUbVmA
8BuaDbkJ+y1ANhMiD+PnxJlrQIZ7Dz8Am5BnYNPI+kuLCNgqnP0hL5pIynh2FR2cxXlgsKf/7dc3
dj05YAPfbGpThy+pKF2OvxieKkPpClWxHuV2DNPgRBpzyiiFvwwVkpQQ38gwh3E/kv6dV6hVIMKA
fjqO4x1nc0fxpEHoeER8QeF8u9qUztaU0XsM6fHyHmXxA8eEkWh6/4UCc3wgZL3GQ9pk4JnZec0/
hwMDDVArEuxKdBNzghzbRnjrVty1qbMfsED1Hp2VGUs6rr6Gp0OY/lPCsZln3Cn8o4kZHXsbXRl+
HHp8PhQKihZHwQQDVCQ/He9goaLIz9JdfQ4epEjhAXBJnqH8krJk1Pdl4IM2fV87CTZQmtcNV3H6
tchDvdoq8ZrgMZkjw6CHzOFXfPTC5CTvFr6s0trx96OG8AzOQ+mveg75JCWGmhUjLg6ota9L+eM6
bCPdY4SLtQ60xgAZ/jv0vI9DDWk0+gX4dvnEpazIY+rfbnRR2ejQLYdSUdkI5T6znApToFhRdIrK
LTZblD4zHX8JSXZSOiCnWUeiIFdZO8kdHX/AQgbuCrV6VaKSFYldMIrxWhkKpe2q7AR7jzObubj1
kPm/TfDiIcN/2iAy2Y1lXnuaKz1GAGF0+utfIbt33EzZY0oj3wkcEyth5rJUDTdrVSg8Rmxtza59
znbIcrHN0Iu8HSADia7xhktTwn67n7w6Fb0CTCvjIE6rX0Jz0I8+/iVAv7BTfIP0k7JzklUZM4fK
EDPlH+5iI4W2a58a/QXposyIM5TXOzA6qlmdJKnd/5utUf81U8HQ9oo2R+SRxYIIajrZrJaK/GWJ
QqeaFrv7x7kM0FPtteqot9Xk08kdAgWu+ypDUBdKxbhzm84T5Ph1bTIknrKl2k1h+foAPN0/5EI5
7/AzuObInGsvDV2A4s1IVGB/iwRDzgpRrEKQWQOkTzG3KXUm3m2dJWKJPK6p9e2+HNFvNPxpA4DW
d9xlqNY1+yCDRneHX0ATWucxAPQujvAAsNNjbk0R2VX0bRqCzTOO7p41hpO8SAu+LhXoa7AAvbOO
Px+GuuXxaDm5UyUKW6SfTWSfNwX/NZXp1SJeCer7KYSeNVhQV4GKbQoYtusqwgjaa6RMEALaGAHV
PebkW8iKXqNlbmCPozkguDZGU+Ry9PSOiZPEcW6M9J59pcq6gwxoiJsOXHhhEdcwYh493FpQY4X3
YPtPLgS4kd0aY3enOYMB9mdwtIihgZMlgEQX6ZCRs9fiHN2Vaj6XeGryd1n/JePbJfCbVkXnVuO5
sRHJHjP600aBtGwDtSFaLuZLhyiyx87RRb+3aOh1Uc0gP0tfbrOZX9SiFejr/TJKmR32DHnF1hyk
RvmK85+dGcqH/yND7Pmdajxe44kycLq7cuCxapdDz4Ce3PR0ReFVp3bSwo6ZzozJsRK9J9RxlN2q
ZSBrSV7IktSMTjtDxjPButnfn/5nHgtqZc68Ud/mtNxop/ZQAl3d9vosikNmztPpykLwL4FhIcbr
AcJRVbV9yhOrlLvTOhA1bgks0QVNyTVMRudVzDFrCPPK6cUx38O3VMXOFxZ48IJ5YDOcrpXhvBzE
3eo4I2FWmkE8RCeP2hKJX01ZfWxS0YaOx4YJl5VdRDL8aD/qs2bZKJyhMCX9S3s72rZvKupvcICI
zEOvlEX0ty7c0eyuMtmKQVeVJQHSOzYnn+oDAqYL6H9fY7PXJglR7Mu8LgjghJ2g/fhfxq85C2Bx
pajSwFB1gRQgYzxpkQtTdQqdc1pHj8HcF9AS0yJFAbjhteSvP0MQvsm/e9fk9JVzYeL+ErBrMv+6
dSplGcdeqHJvEtssqeVjEy7LsRE2DN5aF2Ijl2qvSvHn/QliZcJnrFtOnlFjuwT6AsnqSd865VTD
ahoNeBRRjiIldqadY0lN2rf+DymQsSnhOhbkz7UT/FHt52jELaD/4pnHOKHHFtD52GJpvfKPWAnz
wZ3tZS4Pukxfm2861DhEwf8li40V6zEc2FF50d3FXDnmgbyavxlCi4hKVTKN/jWwp/keF4SRFZX7
m1N9wfPsorO5dZo2n3mXs1hM/chOg04roTtRzhydCJ4ie6vqI1s6cdOukvdskGLfWYEXm3PR06sv
x3mr3Gbp9nN0nmgwVBgFX5ofXrqOYpNttHW1n0C93zt1alx/+IgCs9WG52GFAYMUTWXhlkm+id8u
yc7NKAv+cFgOjahik5xBf8JeA3T3SVJke4JjPoi9VtmTMf8m+AfJM1BZDkKcQnKV5lzU41tgyokw
+8yULHnCZv3PlYzw5Is9ng6v/8eRZFQGA4lUz4rM9Hg2tsmCVF2Z5VvB0X062nXduevBZPkVQiDu
pVGDiHj4iQSP11qYEm8VPuF39Tt/VkXINVR+zTm4RxRZnq93cpWkrWEzCxiEM6fRtwFY1mldyLtT
3/5jT0l7U1CZbUOYm4nJZlk4GwAYOAmV1UBncj4q1XJFy/TpfRm1LbqhAUrYWrt4HZTWbwlkrNbE
NKYhBoEO4W5M22Ka2NvJ7yzoRMOHDPUm9r/tTIysmyRaPGCAmUUCqyIMAP3vf+aHGEwzIGYK3BFN
VKnDmUm97h5epJO7dRNvXbfp6mWOMx+yqyRayhOuG10JgS+n+SPliYDZJdJeVBoaMrkrEaiHhr50
olLaWLUAHpMp2kfSwy8VsQnhUHAVAcquvjTf7RMbL5emkOUhLC/yxrCyNQWevZeaad6fM8etZD8D
1788X+pVNVhxZHpV9mi2Hz6Mgp1vRVMEmQgkouxYYSDEa2besDQ63refQSNpuERMbcZVIjxnGiNA
BqB0gAOkddGC5tAD6HsVBlbL2KRvJbTMYjZ+fomQzwu6ObT2arbhOGWf3dJu4EoV2pPaQC0Vr5wp
dtIhXqZ9pLmat1r6l5AV1aRetjeCODtRTN2JowykdyuHY8rJgyVM3o75nq7pq14+V3Xr7Nr22lkM
O+q+V/NxFKLeO49K4zJuP6+Apoy1mcYmBLtwIvWWCML7F/9PFHKpX0NLHbel2/IppReRvBde5ydT
Tfayl2shiYhdSpki0spcVni9/sA7gZCTU3EOeGJa9Aurjjsn5/1JxT/ltcaQkCR9itDfJ1/3nXTK
FziNu4GcjNFnYiP7R04uETX5ZDeyH+TR9qRBA91N44nkeOU0UaiXPDlxF+iObuMheT32L9d/L+An
alzzv7C0DBuU3WistA0nXJFea0ZpefaocyF96GMBzxYkpNc1Mw1pisQzr1eF1sDEEb90GJP0FsJX
/OBcSpyXoy6W+SODQ6wgt6NNsqcBpWZiEFke3rqbwu//0PP2QoFM2rlaWgyr5nMBo0xajyCz/9I0
Uen/sb7nt1ywIW6JYoumUfLNJvpbhoRWXxoYTHmxc2EQP6Q+vfAYm45tHmVaAXOFQKzKiw7b0uI9
kpd9HBuXaQaSdCpga6BbsaGfAHVUX83p8xz5yq+04vftU5WYOdXbtlEk7lIgK21u1R97g0YQKCOy
zDKKCR7LLav/OUAFHVJ4jymnR5qBgGNfy9GwE6YgKtmQGFZfFZIcs8x+gLu3ee/yfUFXo2V2+/y9
gbAQBEnjc4Wux2RABe8TRXHnF52yo17LKkNoDtAxCxzjcQH+eNSB4QvZ8Yrf+JoR+6h6mNBAmFgx
JzfYWDclSHvy02o/+W1IUB+zpkLZDn3TZ1jWuuiZv5XjIwyIPwUTlAA9Gnp5k0pAf+51bswx/1A0
vaHAR35pih1MhKsD2W7KsUF/Ei7i+7m4jg3CDU7uS4k21gZzXLXu6skt09wgaeO2+ZjNU5HU+S6D
ZuWpKGn5gz59WPaGPCy62V3AjCE3SMS5H0vAe9Z05bugCmWoEnv/MOQ31t8CyoVH0GqOC1gv7wWE
1Usguaaz3T+bAaeJeYiDgiSvGrwzKnmDx39iD/TF3avMoEJRVBsvHfevD9IEP6Wdzh2g3dEhYkxX
QZmW54iPtUQ3PNNeSuFam8lBttD3LDbteAkksL9IPtgInAA0RNzjXB2cCl9OjyLHkyo+Cl030V0Q
bus06OeqrAr0A3ZiKrX5YD8avRnTU7WMYaJJ9Ak0dWaNKvuSVwlUvH1aAAjzyQctgN4Y46lla81Q
xQJdngCv0dtIEijhBw4utHy5wkguqBPEOj9CPrKSBJ0B+SoWx2Uiy5cgq0KfsO2BMgL4sVSlhTNg
we1Xs70Q1UEY8b0vT3zgcwfrrm2ivuxVJ/5KRlD0yBONbjoeBqV+18PQnWW3L06OW2CzvKGzUP5d
VjErS84W/SlqEIrsRazYuHp66sJ6HP5Niu+x8PXeTGiMozpcdHV5DSqbxsJMi9/8rUnnewGbwnvz
HQUx8F93RGbobjkWI0TV7O9RrNFhYnvJiw+9e+pHdt3Irq1wKqUnT2/GA4tj2t4bp++DBuIwp3z7
yHwUBcyMFvGejUXCHbkvVVpsEnerGcKML5XHpkQFM3T97nZg/YJdmoixS8PyJoL1lggJ+WApO2Nz
GVsmfck3+mWytyRd7vu97NWdHBt5eQgfyhhojgQGpVdCmOyeHpmhr7jNQni86bWhanwZssc/mVLq
49UKa73ic1vE36qnDRMCcmpItfJqmBBoWeJfHqfMSTCcxs/2ArByfXJ06u/bADWbXPRrI860KAjc
tLZAxQphhWNuN+v9pkGx4yrhhnLzr9+pm/tHSDZx8qSJ9+uC1i/V8kJge9e32d/ANO17Ey5Lgdo6
UTxrLFXkFwEF/pSD6ELvuO3KhnJR9hrhUhoRtIU8VvLHJ2zMEgqP26KIsz9B9NZdON1jVJqwWYkO
dEyIn0pIXUC7jv8zM9ogTpdzKDdBoifG18QU/tWoBbqhdrDxtW9kesmce6sDT7fMSilxQtNJlHhi
BIq69ff/2bMliyV2zLbw1yMlXH5ggE8N7P314F3t+Zc7xmXW36AVkE0XFk5MoP9a1+eDelKhIUQZ
MV0lOMOciXoPhQhuuHRGmqZoBaidKpELTlRF4LOCIpi9KigCUSOHiFBXFm96vnEJk1QZnYe8oe4F
vHne+RxnZQhpGQm81QoAV8XoUZY3BkJ2btiqgbGTHtLSk5tSnqj7YTRbDbBhtU3sHcvvy2WWIe0I
H8itXTb9MLFZmjgCaHl+6VVmUmtSshwF+weacuYCQRav8PjWzlzJH7K5gbzmDDK4glAQTn1QWk1L
gwAnaJGW/AfHewyLYkM/Ub9ORBl25EmxZnwv9/sOQEt3Efc60++ewI/pKbFkBAiC1etEv90jQiGY
sUtWNeeUhRAQy7w9GnW96t1a5VpWfMzWCX6Gx3BG3rSW1p9166mHBfGlHGKkNoWdJQWPpJfUwZi0
HeCqNYmeEHUX5KZAHSpQD7/zU2zgdNGrNtTypfg/g6//ibMqg0QIVb7A//aup8YVh/UWEpixYXBV
tsK6PgBUmEDns6PZSMHMNcRzNQoWlhi8c5oQMbn+U6Gr94P/JZ0LnLHDuJPwrKMQFQ37x+j3SlPT
KapodFIkWHkbWqsQ0nK06C3DavYHIwPLGjK/VI3fyFdtFpweq2vjeWhuJq7r08GQ/99tqunx86xq
s8VTSyahakxL8H5AaHv9ctQdgL7TE+oIxUbrLyvcouacPCfBG2O3neBeo7HNxq1asHzTElHlid/a
3wAlwsWvUvG46lQjBCFiIJX2TR656sQTRaVki70VVvm59y/MTZyf5vf+9gU/oBacEmkMkNUEzycT
o2KDueWeaczIckC+uR1ZBG+clIaJ+cY8vOdq9QryyVPy3Q4HT61WrAliFTNTB1sN9GTkCJr5aMIf
PQ/bSiDsNyXZMDHOyHDgQBw1/GAw6VRCObcdyRpWq9r9OnDBJjKNaAbYkv3o0J7lABesg7jkmqmv
JSXGCHJgnwmfJhtrp/8mgO6z8SzB5ZI+qkXOrtXD58Vs71LM1adgyrnkt37niObSVCsqUA4QBiXs
UPKmTOGVEpOC/w4JnHUYKlHpIhAvKxTsHe3jGjzcbepyh951saj8C2w/o06OG9ayBM+IRl4YRgXm
WdV58a6wpPgp2KwEaCoWjKlPco9lYCv4gaIi6nueTew714+6OFns8mk+ot9rq3Vo6b7wJZ08qiqM
iJ90/GMMqgSVj9K47aJZ73q8FrWm9DYXj9K5Gkns5jGnC/KJIryPztpkuyc2Wz1hr5j8TtO9JGQ+
QEdRG7dqAZufI+wCXvJDZKZTdkB8msbKawK7V45K7KXTVGlL+kitx1F9c4jWM6cRSvrM65CrWbgh
I4dFQb4kX+0NGYxcW0ukDbDzKyICh4P9ecOmttIYPaL6n+uEoAEApZ4Fu2R/9tbJ2h1Sin36MaDZ
nGKF2UzMu5WMJ9/S1l9xC6mo24K9KZyR3tPkoIzaUkDOB81tUqjTq+F+Wf0HxkN8edT67dbplJAG
1TCoHlT3w/gwTXR+dkZngJL3EQ4n/J4+bmMcTK26GCEbW8AFsb6dhVBGahZGqYGYrmqau9tSaJtq
C6N5Q+78iFjGqorlcspRV5QqMVpLJ8mRSa/bYZFRMm64XwzjegAWoPfIxBDHwd88YSiA4w+rmpi1
Ih1hE967GprKbNdRrePnReSwQmH5mNWpVTryMz5R+PPWh2nmQpEmyJ1cxMHhnMXlDVeEOQ1U/YrH
dlvPNFKS4xuR6XIvSZnBN20/2TzZsMSE56HcV1IXetrAsaeRx71m68EqO64DLUdgHBR2jlAC9NSJ
KQafO/P5P5rGbU5Woz9wLH7+xIpuNl6Bf3M7jZDZp46zaKILYsbE8xXtuL/ouUYaL/w8184hSsnE
xBkoF80nuAefForP0jhtGagf/8P8e7+HKQ/7asbEZzC3R/KTysdbTHUoIvqEGRGqARSx9Ai6bT+m
aGVWZbekxkJMbYAiWgMF85BPZe+akNDmMl4tHGcakPJDCeSzogI4tm+RW8cvmWhgiK1Kf3Gj65Fg
8RNquCZBJpGKlkmVXktDYrCOcTGuZBE1eL3nUWVYg6FD0xHqRd8tCHYOA7fTfkmkIaI4z6bzT9Q8
kWS1nMeVKruiC6+tZ8QTG5Q9FfUJNePazBo8GmogvKV3pkAOlWdev7hZcfx54ZVUAgShpa1VnxLr
jbDUl0++e9nrA+MvrCqPx4K8Zrfzb4f6q0un15Kr219Hdz4Uh7KANap3O8Mm5ltWIg+qbj3LE4lk
Ij2gLQ8Ze5WBA1vFp7ymGTm/vZPgZdq8EPdmmoc8m+uShvKRZ2aDTiSj7Ic1SuFvgxuH5dTF2KK/
hX7K9iNkp2RTXshxdvAHWzJQR+I3DE3U4ufIt8EOjgIBLp8gAyK3wZ1Irz4zNWd8zC0N8/gBVUwl
gXt/pKOowAS/6o4OSfyaoWZUpnH0SS8IlmPeC5gsb3ZzaQu3gqZ13OvF9Fio3fZtc3j4Ev5ZN+MR
JU5hnWyDXBku8eH/OJRthDTjvyol1z3K7aDHi9//q71TFXf2hTfrUCnxT4aXYt0xkwdZ/UKX5fyS
3i5IVJRxr9tgSu72Z/32NZTauhZMJ5sITEwCYypfr1ZcPgr2EfuT/s+XgQs/h6TSpiNNXLGn7YhF
dC8H4BrIMfiWum5H5/kxUxHgJEqF5fNrUzuglPCZboRigMpa3mxGsx3F9PpeuPyW6mZJS57Fthyd
4qAhw+ZgSLfiT/s9NCpNsZMc2JLyE0Vbx15wpx0mLvDLW9CP4xv2fBtUWMotwY7+g596XA4vraAW
slHvUDP4sNjU4mWir3pMpyDBri1KyyYtwz19Y8/2E7uTtDnYWghkA5Yf1SoTodi5gd0=
`protect end_protected
