`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12192)
`protect data_block
KmcL56MVCFgXqPv1SixVZL1VSl9frwYYokDPbOB38Q7c9HMEYPDwIy7DFS7zjLFsnGbCy2IJaZ7I
sbTsoSWcaO2hR6+b+TWM3xYWiLjx705UqVwxjaff1iW3xbbyiubllmEgBdRYVHW+vzPtwxO/5NPh
zx/FE8rUIhvmM5vWZQCisYZwfHnS/qKbIAW0dcYmG6p33vEIzkkGEwOGeS2eoAeMF8ZHVmVRT+S6
ajF4Jz5PvGlpFgZyWg15YfAX01kvZ7AQcRXRs5K9cUbR41Fq7STgGaJXOK6uMqmxQIIGTnuwqdSp
r+ye8wZi/W4/g/NMsLpOsb+OXNwA1yJhlkEA4ApgEgcl3L8EiJQTum4hS08RvIg10r8orWBdYf9f
azKI82CB3xbX96rSkyPfOlhXXL/II521nO+/1j1Fh86owBSo3On7bd/ed+HX94qVDfY68Thc75v5
aXFNN9lweRZ7Y7ZVNhUs6zNgrDjJNhfHqnxkiI97SmReKsuZx++CleBW6ehsPO+TbXnUwjpwI06E
vlhuTrfqjwCKzhgZUfBsND9vtzlDkWdNdTCoNDFGWHPsBl9NNCPMnAQ3fujzYTh+7b8OKhCU+KX9
tAsO6TiWyUUqRLyTZInPGRfVNeWaqCNORrZDCIqpWeadFavphyi/avk6VpmQ1CO38prvZ+1+Zuq4
3FqEW34SY1M+lm+fcph3V1D5bht/avhXVs/vfhswSeiYB6bZyAaYdpe7NBTqbltYcsJrBkQdh4Fg
vIc8Q9s/cjnx12QixyG+yDdvwqkcZOZSHhZ7lQgfVYM+k7lYx6ARGeVaUX7TyY9m6WS0E6Uzj1sc
uDzF64W8DS32OUN1MtXxPQYMBtwuv9B+W/N7L0gZL1RcCnFq28ZfgKl0BFahdGkIDMlFByyusCeL
7OFAZxXMoS5HJo7JKkhsZAYEMiF36CaTratjLVg7RhOU9d1KqnnUaEq8PkBo1YsCGQ4Oc6YVbaZt
k6NikFuY/FBj46OmdQirr+20hQBRskF7EhqemmTiGhjrhCDnfRmfBC9l3wQycvvhvOUxbzCtnV0n
b+cPoXv8bDiWUQEnfyf8QHxWRMzeQhIjLSfLpCB/H73ueSkIJlAEtXIfGzN1hCiBLXif6JPa/orc
p18H91RPQUEgGRw9Bpbyvj6jgjua57VMP3/2X2+1VvTKZ9N2jjCwOzL8b8XrNLVl9X7vVJRqOxk8
Lj7jbFT+k2BJgdulWDZcZZMDjSmHBcuFdEO/gAXqxv1Fo7DIwTxnglileUNdXiSU3Tq9MY7Bwtn7
CviqYS1bsAMR6BwYaj3KCIayiKsOKksyZgF/DMWfPSLlIFzrq6PB2BwiaApdwP2WOm2b60rDxQx8
68JFQUSa3GAJVa311GydsXpJ2RdL2XUzE+FW+O+AYl6bAiKcic71Dh2oacL3HxdQtfD/d5GCQD/h
YewY2es0f01Xn9UUPCBdQCDycXgj+EA0xVeiOEFmABqQV7s+RINjs3VzS+wFcq2w4qQiwc1cNmcl
LaOxwt1PbjFjKFIxdJWsPtafuNPPOmH8Ntz3eGv79O8ojFxjC2jE0ms5W5D+tGaNBm9oC6QFDCrn
s9cB9pGplJo8SiYeR9qtyauVJrMPtOAUIEYJZLGui4FlYkh/RRqDsacqUsczmGn8M4QD3TuAOhat
yznfW+b+xugRCM3m3reEaN9VMfOY0fdIwwEFoKLbnweFoh3yOMEBaCd7VqUu8wK9rfO6Q8A4FZKW
NlQ6XV91lL5EXmhtYQ8boP2wo9Pp6RhnPYFVANNzdqUDPjODetSrQ59LEr8YRem7YISgS1eX2hO9
SJPClJGoHdm00Xn+MgYUUQGRZk6toQMrbwZXwHUKbZrDM4h2tLaATMaPfvLnm25iVc6DCjxmA4LI
Rs3OLgOFmF1H4l2qNxESQlr3vRZc1JualISP8FrNQRRz2swmFKiycmpjTMb+nu0d+pK7BWYNLTQ9
oL5d9kbuF3UedY90taQtSH0/JDdbJVgZhnxof4BbD48ewrdTh0mk+Deghts1viVHCEym9odWrTip
NkfdJZfJ3xJp6ZgM57Wp5VFY09MrOsVFQ9YzN5SAZ8kCToZW46b7RUvDDX7+uLs1X+tRNxe8vkOV
9hFPyvHVGen1mf6riEpcUs58y2zZoah9RQXcv5Lzhknw62zPlCH/n0PX157xi/kBLzo6yfVo83EA
hc2i+RfFEqfNCaz/6rouIrAhmxv4f6JL7w5WhaMctLfCbuE3Wmkc1yETPnVio6nCGKChD1r33Y0j
pr/OD8n1IqERwYaMFdFn2q+A9rNDiOJ0m47qLVgLH1HjVc6bgtl2SLaiIwQEs8sn7nLjsOYkaRua
928v9MTokgWx6l41r7k2caObWo4UNX1UOfBjPfu9EwhN4t8KZHX5ZZb1kq9MvhHUTGGR96MKTmj+
R39WNREb8ucHxS/oeYQlckG5SKXi8lAMT/TF/hc5nQ6A8+gx3yyd2XLFPeZQ3h1cf+WTpXgrwet4
iSUVlSdcbJ8cajzQV6xnCkeMIFpVskexb+nMk6j+U0444aIWUJ7Oz+k4TBpYsbIKA8+JMPdmYExR
DNjP1uOICtSBmUMaKZyG7y2ccI9Wobx/QlZ1CB4URu51rxnSCMuuv0qybDjQEvdHrpx+//kFteSB
oIIDCrVbQxEh9MTO10UXq7CI6IacXxhBu3TWLnzlvbbp9czNhtCxm7j7Q30EE1+crGSsHsIZCVKz
7t3bqAa3g0p80A1L6lqS74/744sfr3AOtxexb5TDfROf8wqUsotcZLew3gCYvmnyKg8Gk9lOun6c
DkXI11sEQosoAJypYZBFBG/1Ph0lwXatsYwenHhd3L4MBNX3uvhMW4t55Fkma2h4EOrlDC9x1qew
hGfwHQfNqCEcwEoAwW2NVTcTaQ4IGQyO+ivjezk8VgTtEVP3EdsshNlZMtru+32T0Xynri4YA+zP
LHSjatR5zhQ54b1aEUONpes0IAVXY1AEKCB2KbOE/J9Pmpq3TuFBIO3NBnM3LrfgnvwSiynvyvRn
Kga9Iq3QH22DjYVUc+KVEo0IVnWC7JNNHnNugfY/xzgZSpq+ghFl5D6uhgM8eTSWWZHwT4dKXumd
uYKBpphfbhgWk7G5DkoOkhPg99qoX9ztpGhXnhaISQy0YqldRNMUJDqaxXrM3oUHM20gtydSRqhP
NPgsVKy1OyXlxUmCaTxaKsjD28DbRPvC1ZS20Wc3oa+UVuxVRWr/MO1uR4IZxri51BeNaEng1r2L
ERzqz1KzmEWc3Tneiv9pWu4/RWzyuKVFRZxclr5nG2hGcessPNYYkAc6/eduDFw1gJJcJ+99DllW
13BLxuZIwjCT0C0Tafopus45WoBk2GRkBJqN/tAPF599lj+PJAeNUzpYmtvGJy+2eyFJZ9t93iGZ
weCGFnNXN6Z+qf5JlGhatUaZ+ThJz1KX+4F2XiB3vdHDTwVroP7DLHJKoc/oF7soQ05vLalL6TZp
HDx7KFFZ3DMB6P7N+iZHht+lzdVw30J+0OBw+o9v8opuKkY9QFVcOU1Bd5FLEszxQ3s37uDqZH97
kPWpNIrQOBadHqGZqEqqaz96hYev9i4D50fOhnTV25ViiknQ0Ga0m0IGLB7crSSMbtxG2l+aDMnF
WtmfD8pDG4c855gD/FD3XnS9PcwcwIDf/Zjrnbb9mponNo0aU54Wq7WQMNvN2uqvSWhQ+xgb55aU
f3+su6V301cZ9lyBLiS7zMdT1LplSsR4JJ+6TCiF7fwIOuVK9Fvz8+lRBT5BKJs4lCVU+qO8unec
Ww0zsLSV/LI7aXGyZhfJff73i4MZO/asdrFOs6KZDpSo3fXLJvf5ikgQEW6Gv/rSPqbfy50gHivn
dyANJSqtWJaodtQg5ZQH4zkCsMO+G8Mjn7LHGRrRkdEg8plnuEz8uIhsNM9fiCj0EiLkhGBmeTe9
w8Yzq0VoGm9SRnSRmAhKgpPQRH+4kH4nBWW1QckyljKkDRfTnyg8D5+ppo86PZ4ghWt5B/L/3kuI
XzyzAkdHTQWSI3uSbXTdgsq0xKed2gfffeSqQaq4rJLKOS/uRrUQySfAcyWMulYtxG3R7gd4Ywpn
T/DGr1uIlPdkmXvBW2yLSG1TdsxKr+5f4fVMB3Ijlla9zhlILQ8erT2jFlmSngY4gqDXMdoRUieG
9ctavWi2FzCtDTAVzz+uR79aF209NsUiPNv9I2a189y0LHb/Rp1dM+/d2wydb21nQFn6Bio+2yLA
bq9qXE2UOWj54mklHC4IdWCFuSJw/ZXddkqsL7dR+MfJOzADweKe/81f16SAFKlTsq249ddwXb4i
ILQKJb89yiuAyT/WHRd3Gz2A2r+8AGpcFGPgwReO2HOHygD6hD5DyDL0+ezamKz9kXkXUcQ55kd/
ZgXrYrSKmbdZOZoH/j0E06V02TSsIF+W4i8RutK2G0YAeAUIuO5W9vWwfSr+0Dv217mdScka+2Ym
qcEnjyasWMD84FZlZsIadBaUWvAg4mF9jN17XBL426Cq12iwvXmZFbGXTCWNh3saA3Rc86o75Qfs
lDhY/O0AUF+lZme/ObcgS8cPELkRWlbhsS3qYj7+jJVQPXix6OZl9h6MHn4U4JZnxtd8BeSybKwg
QMz+X2GocgojCty10fMG7o92yzi7LGQ1zcgl0aGgIVJWOge+I0xE9WwK5hvcyq4Cgz6RVn7qZRRS
Fjy3vmEH0VLp+t8vdat/Soqn2GXefOLDTX4t2lJ9gRhtNEqfyP7LaYPjUdfMmC34uLzxtuu1WuX7
jPvjmNMSQxRxUI6S5DlyLeKL3FQNHS1gqQBNGg8FNlx0ez/ARwpVkb3pjjkPif74G3sLt2c3CnbE
B+5ZsgxjqM9zcb8iTqm+slEAmqwPCAxDgUeF1zVRwTGV2E8oRajsQcE8MO6IYm/9eq71VsRdtzvq
9UlCB+2y6xMfJSuvfvnp4CBgLjDxr62h4Yk9Kiv34Cca/Ux1mOT3iBXWx2RkJdIXZ1GOfRW6+O1k
iXjaASvHlxfV2v4fvDZeLwdghX9iQMoDJykos9YP+lCAM2SY2LSOOELWP3x++uP//zQ+EobIVxMg
jPlj3n26WZNvfEp+Ht0VE33L+kfNEJKEH2jjJHRBKxJY9VGgJPInytS4uprNviXRMi6NaEAizyVw
07wKBJUtIdi02dXCHDxg1lKQ+5iiBJbyj568hhbfsXaWYN71puM1lpoDcAoXQi0VQGreaLK22DJe
7hOLM3neUVy7seeXfQvC2nwFlBT7S/9F6OUCDBLhqc9mh2y2qYWGp/dGgKh0rd2CVfKhXPIwFDQ+
Ifui84JMaLtVVUgw5AErp69TwR6PobvLOp7b1fEYuGjJHB5I0gLznFcsXx/ZjVQ1uPUqqdq/hNjn
nuZLHgNv4wEDp9HqHhHEVKdImlGQ5TAJY2UjMEpofN+nO+FKXShL2B29NE+mIb/Q/jTvFk+L0k88
gKLq9oNYok25XgADi2BEtmOLj0hHqxP1Jw2+o2qImJqZxZNPxNnaoypOKD3WOI8Vi3yAANU6ygvf
3FsWbeV94jDCdSeYE8R5FjSKEoywPd/noyz+QdGmbDG123q3ku6AvkYNEW2qCnEEHsWg5IWvVL+z
M1YJAWUyX3HVNF75TjOUG3nTYMyLBvpWie1lfa9YmgXhWW9mR/vfsKW8zGNUUPG4t3jPXPKElusL
9SfKFe8cmQ+SQCihHsnDEgwlFijCgCqLwAQvx7RkFSmL24miIem/aNzNlAwZ/5fyeTdrSjNuIWcA
X93pbDTEOqJXo5pWJ6RwttaFRfe29fzMShX4ATxVSzIyykgo9UCWJ30Fs7ip9rDfv2vP/YmFYvdB
XpOfS3LRHyAf32Pl9T44FjB4VOQ7bRW+0tz/iA57/64z5PyqjkVqfHgM9jdiue04IfFXDXfXnaJ6
oZlQk9htNnuTgZxXo9uqIpOoph622tCNBEAP1K7vOMC17M4wQRAu9ha3RlcmQtooruTwMb1VVj8o
fTTqIwPUjRWXokmDNxOSTPBko9qZJxEf/iE7WHD4kzT6Hft4i9F38e0B52kMEGHgaVYl1MfFDBxc
w6Nhlj9sVxRNu2YhWF7p5Qwz+INhy23ndNftloqY5lY5gmyFFcCqjdV1sZl1/cEkt6IBaKiNFK0G
8ymz64mvKOVxTfvbkbl4Ehuf2GPWaXPY2VWzrQvUHa12JZxpd7qTuo15t/D99ElulybEZQ2Op2hy
WZwCyqHBt84MULp7/AU67ht0PoIYcGwaX8wbOmVC8gYvFZpXVhne27VRpYsp7SaZcFJuKe+ptKjS
cA4rE5M6HCuZnRZbZjo5CyOIyH0fk+2aLdg86kfxX2CUab7DOqrxjU3qouzXGuLoyL9W1O3wjubr
NxeaPAhQILRPMahXnM9n5BV7yc0fU86OvuYcsADIALlb8TdPWW9203R9l1PpFTa9jUJZcq9nCl0T
r3U7MvGh54849uHv4habYYn9b+E+AwGZRig/VVM97Pd6D3rgjwc2wA+Qz8s269lTGYPzJj0rXDvw
dO5FgkI9WfvMLtwkXLH+o/iQh9LvX2Kcmcxj1GUqc6/xgOfH5p3wNZXfTwnH7Y+iSGKvHTc6TDPO
pLzuh4xHD282nnuEiMudwuCytuwTB0Jel/Ab3m3ZuTYmm1AbqQ+YRDKkj0HdNaVEPDNuo5vh6usO
3szEKxg4uS8r++nqSr1lNbw5Kzzx8CozIoeNKknvJ4bUyJS9RD1dOptoB16XI9OYZ7w6vY/JJmqn
8e16gRAkdds29jKtMBX1BhAKhy8D3hUqGzCDZgA8DVS1nQjRYp6sQv9yEjCOUQEOlDvOvpO3hRIL
pc/UEq0EVu9VoFf1v6UW9XazIFRnMd+TZdTFoAWZK/WykK9GQOIt1MolnZL+ZOHV0tDHBbFYqW3R
1v1YOa1yLk/2Fe9FxXAOUmdVnSuf56/nk4iUtVq61+uONtj2RDS8Zg2RXbpSA6z3sLLshQqtSln+
ijT8PmrPIsPBSiRs/YtLp7PCV09/eE3kBqcnZjno4vJNIBPAM3QisBtGUApGYpUpiTLHfWw6aHGF
8005pZNs1aV9L87DJDSnB+q+gXx9M+V4AY1mYXMk5oFn2GVRfrieKchHUs+PRojSMHhxnaudV6CG
J4gJhAwOsD0iXePLAMyN4bEec06QD2xeI9MAwOuggihuYdrk64qxP3+m54+E4Ff3i8vkB4uLlNbA
+A0dbs+TjLjVgPJjG7hUaQxZBCvGasdDW21YMc7rREXAeZ+r/MO/UhkiyqarbwgnwDMJPvhChjn0
PBjFGkbvRbFx22DPdPAslehr1qYUl9+PyDXyZWT//ash3p59FAxkMsawx27xY5arSER4yIsbUp+0
h9cZ1CPksE7TP0GUdYNIS6RPg0SH+IvATgPguwVn9UmoU1iPOnzKcEoGzLOHYNg65lKnKk6plxIH
lRVAU7SQ5mAv22SWBC1uLbeyBfKcXjpX8YD9GgrDCndPULzrt7ijw1UIv94oZAVi+SPV6RPc4d8n
gTznzXMlUaEgiiP/BngZSldhSs3h+4E6wBDz/jH4JzbbTsnWpLRdszAtuvdAYOM/pNG41uiB8Qp4
2b1clHhLfw70J0bdCmncn0jMYS9dOUQWMW/vsRULnHOO6mB94cwIa2M8+j7hcPKsOzaguWSOkUAI
UGAhfStnmVhxQfcfWKpBQ7SOZdHFnj37v5Cd2auQn7xK6uyEtxOHy/QlV0L1xbjKqrmAFi44AGrb
uaf3tkdM6qGF7cCe3xuFDqRaHo9J3YZ4MdfkHvDG4C5OiVcC7qwSDyhdrbawI8QEDqt87GvFazCu
7yCO5Pbu/I2+GumarC0X8tu7alpHpEYYoFIZL2xJVPOLuk/IeRiHRz3oJ8pIMg/ziJLDA4U5+gT5
HEWG+m3VXQtOn7lMBYz9Lap7qWqu65vXjCvQX+NvqeyPY/xts0LB/YLGxbKjpB84TtaLu9KYaMOf
4FqCbV5e+4GDKcHGTrcq8ucbd2QX9VS50Fu9kgfuvA8afMb6ZgzTmxAlP+LWNheg46zW03Z/JU/d
5eDLsvhT+PWYFyxsWcWpI6aS34gotJxkrMbXg7RZ59nqlCEzXQv7oqMYf7wgAncR6OXn3mJvoGIy
KK59Ny47ECgCHwn391T2dzxQL7zupRGeTo2+JJnxCK9DWECQtDFGy8aLgiNkQ6q91BfkwHQo3Hsv
rfizWLmxULoGB6jpGPSGsRlfYMZ2/DPrb9pEcg9bdCsjTnOaPzSS0vr4ClEUFYjR+PT5hvoAPVqt
kaeauqu0lHlwgCFa407sbfM40CUybEwQSZ7HAq9uBaHVmlj0+sEeYh0At6b4wVOUuOcGPbt6xGnV
/69DcJHzaCoq5MU98uyNQF4UkTgUInDzeNd53j/nR3dCTsFCYEmm1WWsVxIinz8ZaSJxi4MPPjby
WUJvxNFjvIcZf6gl71CYKrtLM2+aYfZntUe4ZxJj/ZJLY04oEqMzuNWK4ZGxxYYvpCSB39dX+jL0
NSJLRn85LJXtz52Rrhg9zB6CS1cHWP/bgyWkkyJtAwNKDjoAAzMk7Os8V1LJ+qlhIFbO+2CYLdkK
0VFygn2CjzWwoeI9Oom7XauqqCgeXUQkFfxxhh0Gb1pgbTeL8+4wyXWmc9vAm3rr6DotOoc2YWHB
FNVSZmB7XQtTTxhYvhixSCOEXjAu69U+6no2CBYXl6DQqIwDRa3/DzOKGiOhV+wC9PxkyRKs/F8B
MmJdxgsBH12cAkB5LMHDUhw40JRFU6rJlm7edheknIK3SS4HZhGWSIPrgw1yo56BeEMZ5Z0f7XdX
y6xu1DBWZENUzf9MXqBV15bCa5rP1otgsepffLQSqTd53pQRMOUPidCDVDCLYqISaQNYEJLjgodf
Xk5XeIb/WN9TcXCHTKTQRG4TbKi2u6Y//U4LNjiI/l5fYCMtr/3xsdfoGTFX8PjIcA4Lvp4Mo66M
rnKFHl31+8ApD7erA2NDXgN/UOUENoapUBDrJMqt536YWgMbRPBSMSxinoLD7TIZ2Vu94ZmwfHKp
0klO0+bsfsPVceqNeBmL66qFWOPZPEplwfEkACNFkFGzaeESjurt/5w8jJhxeI/Z+9aYarnx/8/Q
EUXR24qdVZ1DqwcmQdyWHypDhd05RO3iEUxNPl2nQPIFfAcvCWCT0YPL4iGy1TY8WlboMNu6q4xL
hqL3tjA6u4f6ES4QB9V6m50TlxZLfPC9Kdr0RPhW+7OcH30ffPOkBcwi/B8BgMLduHZFxZYDciuz
ri/SynvQxd5kL+PrHY1/IAQwooM10EeOpUKsabrocszr57oBC2nN1i9eOBWNlT/e4fyuYurXUj93
3Uzo0jYCbmjrcmqMkGU+cvb0tksGlHV2xXf0ilwOSLLXehOC4UL0dbuQesknEdWOp21KIN5PBPJ3
p8UK0f/aQ3drqqDK/lDftH9/T/Zen+5dSzcbpm0oPDrAr3V1uhgzQtbEj4jmIauIgo1XMJWvt68V
DRhBC8raIhC6kn05o7hqmV4tDCCSTb1Zd+WhCJDUgBG4seoWrVShft5b+0B4PpBPfNtXFJtQ4n2o
h38PZ3/xBjAQ9kgiBOXv4aAGwIadPC7bHNG/F/gIXS++17uviupFDgd/gWKTJ0aP9s7r8l71rW3/
DtckfyDCbxjyCLWweOS+v1obkIp6QzbBE0xA2QyoLMbKUpF4Cr3+cwMnVKO+BAx/WYL3XXxQ0fKd
AiWBe0v8QWI+OX8w3r51zhioCEtcG0LHVs92PuGe+R41GokvVwKwu+fes44vKTfrvY/+8AiO9LPc
wD5SIDeYHQJtTwMRn0pc20uwoC81LHV+Wk5E2+qNqp90kEZr/g3WMTIhTL0tCqgxgZ4W/okxWe7U
lXZ28C9lM7LCxKcFmI955M8yWNC6dO3Kxb7ThRBSFFXmccG2EzVjP8IuZQye/5hDJqH4+RH4HqFW
6f652mA/XUX37zpGMaigdvme8I79H3XGW74kaYdpvzr7v3a5J9WUUNILU7GFFjYRIpJhNKMpJIY6
c0viUU++jVgQRgNfFTx8O5IGyBhkT7J2Ul25C9NV4jnzLdnZKrmiBQvfaZSbMC7psBjb9HGjaxfu
cJR4Hynu7J+2jc3ZSgDXYY4EGKVXXNlwGKMc+5mj/hu0S4hSKiK/437VvAnZSm45lOTz6/pxIxUq
kGp103MpVyFb2cznXZ0iGSa/c0zDGoKBDGeEXqu+XThW8ksYY+ZHt04VqF/ew+7I+jtZIB+Arm3u
Ia+k1qpui1bjtD2j5F0vnW7KRfq9YwKU1O3xN6zo0nNNZMUAXQneLAihEGiPiSfTN/n5mxJW6G8u
+6jEW+8WkM8O0N/AiVz08FNIzbH7Sly4bJU26Z0sVjQpzuV4WSQeL6aIvKMVUGemzuv1O+Y2Wasx
JRNiKGne57dXZgz49BBzRJmlzLe8EeYNF/wqdhwLKuPI0uAvYy84Y8fwS1sLrdaOu++8YOEQa2XI
jIHtYSpYMHUlxopE5VpyjqsLpCTmEGIrG0U00X+2cHu2s5UsP8Na4lxU5M7ABFSVr6LrL2GikmVY
fWjX3PMhRCc7HauIhwaOFiONp/8/mjCyarQkP5H9hIKqJAffKw5QfdK749QrSZhAWjsfaVvaD44i
wEY4D1irgF+y6RHrBewdd1TvccapeeVJLPU4hE3FSFQtkpc4ZBs6RwKDd8aSdJt6jrYDXUW/tx3l
xXNR3hb4xIX9N13BrQNvJ4uy2K0xfFrdf/fB9/GvwBCvIlbQyEHv++kF3UfOeMkHxRK+ohnBrDlK
nN8GvdAH108LyPa/wMY4QIvgZNgTWD1uUR9D5Cy3dmNaqpLdxSoqgqELcw2eUulruHjPLrFMkMqS
2QBPS4uHnAWzFnFL9aZORf2Bf8WufIqhsQ1sN9WqQZ5S0H0IsCC8OlAHYvEU3CPcueJuUw5zedkv
P8VXoezyvwjON1rnHDwe6F7bbAbxZzigswl4ElI9ZzzVuBrRo9C8cpr36uiFMA4dHmfzw2IiEDFk
IWNxcev8Uc2/D8eJ/UclCk+/W4qOsrHo4g+dLLcxPB7PNAfhOAS+ucFRPOwoD7AU36kXKjrrYgdf
jaexQPPbVP+V49jwU3xhllJNkW/kuIqFXcK4+eOxVARfDXYK5hfUfsSJ0kxkhx7YeKxA1cxeViD4
HveYLzNSk2ohVsWOeqc/rabauCsRRO6rlUEzEbSv5z+HP4rg9HCohsND0eCmqePO9tN4LjqSyfuz
+6CLPlakCHq1LJJ3obLsl2ye3rz5VXRyNU71uKZPnp8694hA4eIIfs8PtXHt8z0oRpBRRbNXZB1V
iJIlxE4l+tamBRcYnH/RlAkZyNEEhEPonYfBYy2B8nZU+hpkQVrGo8cyJJYxgtR/w6BS0a03oKLg
cvt5p7jPDpiMoqPiOkAbYVNu3tFPlY/tLGLiL/VDD1H4kaKc2vUoUfDnB1+kb8Ma0JWmE9BZ2T6X
b3JLIsydjmfvnfdWFhulPyk8SB2Bikc3tpn/I9yahH36CNX6nQVcHo+1RWbRa2i5VV88QIqquPIO
jWHQnMWdbqC5P0jQEWwhmvIRum5tSPKCeBMh3VyjKtZsD0zMrwtayXgIsLxMyzg/+UQFSv1wCvfX
HqflhfMkitkbp+jLM42VWKGdc4/FqTiTDq5pjKM1ZyH19Ajffkprnz8s5okCaazEIwdY7ngQX8e5
jb1dAkwkifXKPLCKmFgYKD+Zypf9+sxrD9CR86sGKqOkkmhV6+HP1ovNeEhji5w5TSHJOq0cDzP/
bS4EdtXYaSiSOxDWCjzCiTROffhFczwc0N8K8bCkqdGraMMITvBpXSBWSnXnuvtdEka2llM+/tDX
Z2GWXDCVyknchQqBBwtnFiOqfHNzOvBZT6Y8nAtl9gHa4bycRXTyKNrSOLy5raS/YccDz0ZORQ0u
87uZYwamhmb2t2wqw8guekWaYEh8PRQMKfRVQDdqbEys+poVnrNQQXBGTcDpYlzZQ3DBqDZ0YlhT
Er/Yl6zXjVrmC37PTcNn1q1mJ10TI0yO0Ghq9Iniqy3YHkboYsdpi+4lnY1i+EmdlqQORKgAyPR8
NLcoFWDwhHhTOo1m61A178+iD5628mwubAeQe1zYKxIdCUv2Zen13ylNr8TOw05nC3DazVUpHVuo
AsNMQQwovUrU/2APAo0zdxPVhl76xxz7Yr6SsNubWUGZYm4FMgJ3omxfQV0nQVq2egCmny6V9MZe
T9lovEEUYgiey6EhQS4GQBqfgN2WZ2aMU3ku50hY8tFZ0Z2CTchuHDUGE/BKCCN+mtutS5m25hke
WLiMY1c3UsP+fkTrLB3pCeEwSDUcoYNU7KDm1gOp7lFVhRPh6iX7NGhMSoHP0UK2g/JhG8rShqAO
lMRQTtr/5dXGsOIGjctiX+maMqYpwOy1Pwsp+Y0GnfMlkZBAkTv6fZu7tkzYYqxFOjlAO7Gaq2bU
1gHdA9zBoDaE9X4gf0HXbmDF4UtGvTbNzIZsrYutpndTlSu1hWCIwumjPiYHs+ckpoxMRWi6jYHw
gr2FydQQOPk34FASaKjSjK/Bv4tw0Mn1HI/t4jQlNTZsD8f2hiH6Z6Wq0wlo8wqmoOJGn6VVoxgc
eL8MrDvWsd0UHck9KFB1j0uHxOX3ZK1636BOfduIutYYdplx5GxJtwutAHEAv1b2it/zv9ci1jZn
JneUQ7PvnEYVS9tJA2CbUzXb4Z/BPiriM3wDgKLgle5/5N0YdcWFGCZR1kpiNTMAxdppcz+DV5+0
cE3VUxznG4wCqcHKviBN4nwtJk/BUYGSZUvrKebF4cdG33i6Ee4Gcd3REIFCs2DOXVwdYz2rQ8rT
CvmMJFvx51GXsAE683/WFhgnfkXLy8Mk/6XHg+vAQOLOPa9EGwHZmuqwet+d0Tp6+ZxbksjQxBjN
/YpWhqQ75DwyCbArDEAH5gEqIDAgmCREiCJ5p373bn7MnNjMt8eZHYRm66J03ERxHxuXMlhD/GoG
/RwTkp5OeH3yXJYMjWLtoV3ED/fuz+Jnm4MvlH13gpnPiujPquiYd7wRdZRHuzI/q1glIn9pfk43
SyGzgF7gSHcgS6iGhO7gtPzvnzPw4qwRJBD75EzMcimrNQ77bvbZvo6T5iz6h0VpVrODGf8RCNZI
KvMoVB98FXOduPvvgZ1qgk1/77y4H88RNmgBUWc0vbh8RrQYCvgmjxes2Hq3zUpWLSXQA0pU9sMn
/qMD3RV4nWsvREDoeWPfeMlHhgDxvLNDOgiHsl8W2XHCj+z8hAWZ/o7+Z0N6ffO4p7nq0vLyImoy
ABVA9kTio/1qz236AkQj8H6qCMMnWoNVXYZ8YiGf67RYLKHVVSZukVc1yihpBKEDr0TCv8Z2H5fK
LP7IBNNUwHWMMB4FfaBEdy+BDGkxKedAPxzio82ZKnF6FspEbvHUJ6lr8BaXsvITmc2QnU47BH2g
2lKYjKHqW3t9ekDCY7XtOi3J84I5mKgyTCuHi/TQZ+Wo/SmVnDn+Trv3ih6qSH0zGnU5sV4Y9tmo
Ed0J0QYN3q4RwtE9asrFk8f9sJ2FqIdcFo9MHzdzER8dWB0pQJOWzVytywQPxBe/jiNEZqEowbK1
jA1qy3DobwJr5fL5bzSSnB861rFdLOErORMeE8arM0MAuODhic0lIWcl587QeeRE54EK8wbZYDrI
TvfOg5JnozXRl2VPdwMMu5u7I3VXThZX2GfqMXknbJ52pcaYVsCWcN/A0kiInU6tcuR+kCu5Pqip
DrBjgIEXVZYCxgTCR2Z/x+0+rNaZ66Py3uPWgY6N4oP2i99rFiCRLp/qwiQab46lbhB16+Apy0g4
c55vb5AfpHzXwbREFpouHZW7lVM2hxu84vstajF/E/Lgl7HatXklaZ3Khm8T8ub3YicQeotFulos
Z1epjgG2M+0P5ehk2/iBer0kN35A1CFVNf6oIghQGKGxYs20Min3j4rho//nx441gyGdmExP2xMc
w4sNhCs8s8jj281QWlwiJBSDlHdQg/mlVaPbRNOnryuiW+VkqqRwQARVKbw8MY0ZPkuFuXdNwJlp
tzis7g94o26CYQ8Ak5sU02smB4ToRW58muNauRLjXIlxPRNmBzmdVC7qewqX8GC/hGtV93PywXNb
MOdrWr9YLZscmgptbj3n04vlzzzutoaUCSFqSb9YcRjMv/W9dHf/co0xL3c1xUZ6PNj53Qy6ASQ7
W7hYvy3JcFbth0cfYBOy1FzvrXJuqBCbHW5esumzHbZ+qMtthcfO9fuQ/5qKnOjlso5fX+pI6PVz
Nq8oTAnjxuNoTpg6Ij5iwVw+Z8MvMi6x83aw07mDncvcObHkHXTT6wkMc8TBp09OeAngNglTMumI
DpOf6LILKn24vV7NyG27BjqdSzxh2pFmvWTcmxYseVtvhu5q6DH3AZqtvbYo/qaUxI6JJ9Ari8Ea
p3U/G5l98twHu1kbCrGPZOqqWaJTupiJKotgnnNAUKT0ctGjDKnUSMBJA2HtrdhyLs8lDU71Z5ed
gEwrZL7egwq9gw7kScrONDHIGlQB04YA2JTlsW5SkRitS3rbBkpeq/cJuPnXip2+glwmxanFv4J5
FQhPfNU3FpmgQ2enL6P+TVBW/Z2EPSqYsFDBQ9M0w6hXMzkewpPQ4V60j0Uno49tpwIO5tGJHKCD
c2OlM2nsll2d2SQsjfM7rHLK5l6MFV+p76qQqYYy/zNne92uCkblqhBoWJY8AFXZ+F9Y0f0tO4Sm
2QQez7YHIMqIYIcVT4HkSKvE8GwdARcGTFbIL8JxR22zmdaQ8iW+J5/jMOI54SshMdzwp/W1tq0W
S/z48ITYhAACP4lDPdTdvm6xHughAtFhMAZ2+REN+8qpogfigcGDCJvUSqTlaW/e6kXKCHOdWkpI
sBkikt674D2ryNP0O4ec+oy21GYhfc4to3Y6SmITx9T2ip2leiDB5YcMV8Xn9TaBsbc3eXAPaONi
D+GrERxU40hbexiGuTW2DY6e7TKkIX96aXBjeyfme6aDnWX0nGrRRTSySPYdwHDcR1jf4f33E/Uj
6WKtxiBh7NuV0w6xUpGqFk3v4nqtam1G+VmTuWLaiUtZ1nx1q9Ea7gbaO6txQtOnY86Ht5ttcXR5
yI8vCkVvkgsPem0ndmHgXA8tWsyMLY5rdUudPdyJlTMpnDkAMeqSFuFNKX3wWyJ/xmGYv1y1arHr
j1auhvOV+FuVgzGjpTpMY9uWAmVwBwjxivUqoPKNfxCwJSSqwDUFITQ+A2dPdoCtj8HhrwUuVjSd
4u7MlWdkHsBrfnAmTw0CAHIpQqgqALR+JSPePjU6kciSiuSrt1GxxM3DTI2y3Dcl9H/13Wjj84j2
MnO0k1tVdBqjk3MsZKdVnfnSNv4/Q5p1SyrNTaZ5O8SNnx3+93twXtaG/i5xUSYC2aFXtNIkF3l3
BM+39dmvN+DmvL0sPkHT/SwjviSR1FBuSxHkDW74u4rlyzdX3Hul9Ij0ERAVEeDGb2BbZFA0Gtt5
mrdAJeA2kAM4y/Ui2bI9PFXjB7+GGMka1bJUYchhIGpKii/q9rFtwd9YLDEiHv46/KWJwvgwGOJ+
Kkuqhva1sTl/bwz61LIZhRapvXdDYAiEjlTK/johGTHfUIkjBTmoB0JkpIzWdkD6dQMKxovzolYx
p03gntM+qESeMyFwwL2fv0EaxXnOfM8t19SWq7UBDpmLIvJkt+N/loO7GCxgWurmlTN44ikkpxC9
XJUiKLifZeAjuAUon0P9+f+W2mC6svfYUHJFPBLeek7uIO4T5RH9HmHbud8+qj2HwJTCaT2Wz0Rd
Ycs5mL2r2mDsHUTKXLq9dEoiQrXW8ofHCwby2QeqzuQ2e7Cb3rU3KYEZlCK5wuuXts8G8fsL4LsS
bmtMqK+EEa0W+fRJd8f8yHdPnRUaJKViQkwSNkyUpsXLZtke0yb1wzEcm2upbY8j5YFSSTNMsuuM
78Z0OoSkEcGVRE/gOmAxQL25hUOAzmqql+eERbo7kPXLTY3+o6SZQpCdvB0H2xjKLyUHRC4l/wzT
veAc27BLT1mV+RNtUpPBSm+eGUDT3rnXUCRfDLxEkabLt6q/DQvXy6Bh/AJRIft7hBuPVPJva5XB
YQUrFcKyIlvSFtHqOfQwQbpp8bkL/k4oQ5FLFP92x+yDKEu9rVDLglGajDoMj8lCKHYdX5i2eYE2
XHG7Tohy3Woj77ZEtRzqed/epiWB/eJiu/ht4yhP8fvOxgjzNpeWIMc8lc5SU0rcog9O
`protect end_protected
