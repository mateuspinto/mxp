`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
QyPjtULsfihPv+J7aIN7zOPlZlCcR65tSMxcWNIyTrZmxQR08fQWuhsv06n26lSOseEUWAvBLc5X
SFd4sATe2Iw8RPW4NXx/8FjtX3slpAkSD1ZWrwJseKTEjdSplz4B362HJCdxUfVrwTobrM0mebsB
upf7ylC4epFPDMVk8mzXaCt/wDk2DvNtqAO+tKKNoaxPb9ou9m7uwC2HqUcwlclwKQFELy80g3Oi
K4XH3V2+Sv+VV8+kUT4DI3lxftmVKAzPuVoYLRPLFcQk2hQVk7Rcce1FGc0dZlvqXVxZP0iz0Sf5
VKtb8kNeFhS2GwQmQNEJUJVNnzFemanj4B3QHA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="Ku6jzowpTUuLedycoRN2GPcTd69UctHaghLiZIAh1ik="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 68736)
`protect data_block
HpHJRCs3EJuPI/YAdmcUtrxKSOb3H+/Om+SmYXiuYDJHFU/UQ6G1WrsU3bANkGXYDbryx5chkNY8
ssPzcccMLtuVXxEkN55E6J6bsU3bW4wIgoDgVSMeK7B9QlM2Umaaz06JwHIaRw7mso/z3r+xxOTk
2+bpJOvNXm1/PWAi66HJ8DMqM3LgD82B9cRtGsuJtoAcwwXQXEM7OzmdCRdZSVoaS/12Fr4dCB3K
QZ9DOteYdZlsu0HexBGvEgizvzHVs7buUvw+ZqVHpT/dxkWKd7Cg+aV80RvFthF4EvtTRJSjvNmG
mrFb0xKI+W/oCOASsUmLou0WhDUByYY9MxurFRvo9AxUZQIwHcuww1oXlatZhshydMHdhGbLf2JJ
4mi2rBvZYIlEhI1vbkiN8oEb0xTpI79geEbwn18IZVGZrIVwlILVvEhEp8u08qBiRkE9awWfA7PS
0LiW1zS8wZkGYCpCmtRor2wV9XrXyIjLXdReTNPEY/u7GJfrI8SlZuu8taLURkmWoJEa1IMpeN8p
+UdQvs3Es3L4ZYOM3fMgVU2SAIHl303yNxeUhsGDCMeycH5dsFHAo9E2lgqBMdar8BFD80vlpUq6
POXGHJqRKBIXlwEM8psh9QmpK7J4Nxbrx/mEdMCKP599YL583iRZdEEfFargDdEYQdiBifNp/S1R
UYMh1muKK0uJGi6k13P1w/ha8IeBqSu/hSMaa4YhZBny8pQWwZASpMlkPXXRwFIj3FVT8GT5IMPw
7Sq2qlCaRBKO/t47EF+GOVlHpZKRycQ3t3oDcOx2ND1nAaIuVYLn49VQn53z35AyNKCQgkYofJrp
WqjQO9Be03CmcmrhJJBn0aCO6g4YTzHZzV9bon8k6YISjroE5pmosqxF9iux+4HEIvcsiwOQkHkN
V2X5aCavknB+75A5NeBaV15YJBBikEzVOKbEFBtKinr2/EvS5abKoyGpGdDfQ4De4Ql2bZj7/PCj
oiP5mz/UGApXS4eOGhcZgOh6t73XMcLjL2CUboOsTKjDlraRbPUapqDNiWOawZUQch+hc+h8RBo4
mjyKKWrDRZ/kguXWhlAevWopVA3YYzkhI/kMIlQtM4fyw4qPaI3VH/ry6qGrMJ0p5sD8+pzTbuNJ
I3Cain05JJWYpYeiYM168EG6mQmc+9cvdyvNFIHyQaSGQVr8I8pwhEHO5WjVauGFH2fC5EMgFZv7
9GuZeyZ1do6Uze7ujlNPt6mZjMkqdAXPX3IzbiFiQ0FC9+p3vrabFd/nFkPDR2UNz4IHSxuligiR
nJkDR3oeMT1mtlCUs8mP2lYZiKPey3WNcHkyOcAyxbGGN7YznRHuz0NB8oCgN/IbM2JMWSnUPu90
GU98BedE5H3kbAFTLmY35oNOyUSZip24t5a+rPtccAcoyg5FqwdsosJvqyp7h7yvxZYhVWPYqj2O
lMXlTjtb36lqwIS7Bdt9pyMe6QWNbeF81qpyoDA11u31raE29LOFUR7WrR7fcbxPL1zSRBQoV9HR
A+gXilhnD77MJ9XzquZHQvq8yIkMaCesbndvpAVHBbgvFiIjYYBAg4PCGnNcv4DxGdMw7UJumdyY
MZHzDTi+WSuH6Z+I4YilFUimBjakCFtgA04xOYfpFmu5F5FfQR4FsQ5aCUYtPJ9EF+62lomQE2p4
lkk8JKapqRaTJlfTrpIyI165QrT/4nvhy7BVwdlIcSoZcjwToaKUwuEkn1noNcXLij/xkVE9jqzt
Fv/d3CaByB8Q7rTW5FyHYuiurCFXGuYDTY5hjeTwOA3QKqYxuZC4KKwv6/KspvXv2LlHRVDApuJf
W330jT2lwcX6rsdBhnyzr2ANPca/UZJmygmwVriI5eaVw8hSqwoCSYFkJrXzGdRMzwEOfdsl0mdX
NHOZAVVmZLJShHIpm/7WBsFFe1Zj8tlQSmBb8BEa7c7C9EHlI/c8shgBH6M1kkoofIq4G4UsJOdv
N4f3YVGjnTJ7ddmb46oi2qnt0J3rsG+Ne3j+mCWWAs45otx976dbwCh9ydgi+DZo6LdY6jLnfYfO
YIpZdatexs2e5SDGqKIRouH5zbLaBNGjdpr5Rs7GhYLw81auFVciuytRICDkUZq3jnuYUbEVyc6s
Zpr18ao0dmxx/doI52VZ3WSoH/MZQfe958ICPuZ4FtVv8A/UwIIWbOjyNCko1fpTMDehLsZfoUfM
pf9yKhZDmqaJ9NJFMaLVyBtvetlivFsoAlY7F/LH0FG/4jGz+Oj+K71FUu2usrn1WQ84IkT/rw2l
3M4VmojUnGTfWC4djJUqUuYavhSK7eERZQdjTApvAWTwflccvFtQx6jCxH9N5TF1NCrr8QqZ2RGU
bfzIuvxky+jGyzvomuUNkjK95+MUnH9d42PjQ5PjcRiWdvZrnAyYpieRr5ZCpW04+J1ilnLrjvd3
4NXOEOZ5lVHqrQIEesgJKR+qBHYy1oi5QJeZUBIB+kWANYaqWutYU3150KKuH1cwCSmp0XCjSy08
ixzrc6zlYWID5nwjR5tvzuQrKFKCxw2+PxwI3b92Nt3hmQ+pro+Alhaxq8+/6XwqAOyPaYoc2VaQ
q2eY4gXbBkbyBT8MMIgTVMnUhJNJ78yZIxLZA1EuGmxOd4NtpYeMX/Ism425EzPYJGEQ4g3EbcRu
94L3UL7GgROjS05TQmhE2pZlXHiihioitxTs5n0xLGY7ZYzPnvu+aPDchpHNqsMeKvt6PCVtwE7K
YRC6SOrMSfcrU5hlBTmV/yURW4MZRai8RVVYjdK5nTZwPcASn3ELYFEmZ3dYQga/v/dMGAF5jFCb
3R7tcgrvpCwXv7UW5Uo+glPJdgxASRkFZkoROHlK6n8D/pESngusCbCZPj7qT870om1ClcivTGUY
GrE0pT2JQan3EdqDZPQ9CsJmnCjK3o10BBgq95y5r9q3Af7K24R9gRFqWwAlCuoOUpoHYOh3KrBr
yeDovu1ZCGyVexgCRu6ELPoDhyZOzv1H1BOOUTw/JojQQICElZniI48sDTlJ43vOni/h7bjTJ3u8
6eldIUdygFdZ+STM8yFUtqEubO9KY1gvQG1f4xYZBS/4qcIkKxJutf2BrrZxH8mPFRE3e1ytHaIx
g8g1DqzAJhrygqBuehIN5ZShZfYu/kQslLOKdsMiJwM1CiAACgU8oqRy1aT53JQZjjP7QH0zdBTP
QggAHPrMVZdV+NWmTgSs28LM1CYFAHiDCGVOZTv/dIWspkJ0p15hLaBl8trrqFbKxyGu9tNsCbvZ
omur8tMvhVnGhQzRESUan/0JP1VwgiZUF1qptLSEmEjI03CY6Xc5fLUUH5jUfAz18E18qnEsYh7K
4ljOCDNoUHhRNRQWks8atDiMAwHUGc/WKKW64cV5s4KIaX0oY0x/ERmXsiI0kiCJfqeRbnhQXsk6
+6GZ68WCDpGm7R1LNh1J2MvxNyaDEpIgCeNx0GZxqdvNaP+G7fTcZAwnhyn2xIjhr7yD9os9xHDe
87WBaqU2bbLr42SkrTdDGJq5S/ptPGK4/9CRA6KROxep/sOB+GdhifRVN7d4kEGfj9G1n8HUBGVh
XpkjEZE4oAFTd+g7gT8Wx50hKCYPjsEwAw2FiJB9wCoFwePUZbuGnagbnFBYb3uSVCe582lzsuYG
PaFBaYILMZYHTIdkHT+JQCboiW3Qu1hRHsTCAN0aWxL5CliMHehiMBA0bJysoAC4hO7J7SuZ67BE
lo4XCDruy6qXXqkL96fGTevxdj7JzzjYkF5lOR8O9YRaOj3hoLMLuZV+DSTQ/obqbGjKzCS2e4jB
61iCbsdycHIVl7zHrolsJyX3vfoESoAED+mp0oalE1y0Gwkx52Y8ResJ62+2fPEZOvxrKT6X2Q2V
S0FP5dY/t2iDI9u2GY5/poPO7s0x5WZGqdvaLG/ow00Hx1hY8KclcJaA7kt7oyp3gQp65XhHqG82
NIhk33YbqVohEEwAbhsfm3DHPKsNIPO0Zs6t6zj/vrKD1C4krPpMNaOD4/UwlRKSFqStURFXIL2z
zwg8FW1qcZ38r/WPV+RtBcG8322DVljA7vSY34KY79NLlTodKDfxMArmPoZFm8JUaDgj/roP8FDA
puyvg4JvDqoQ6mj02P1UzE6ar8UV8llc0OYY5CWn70YeorP+C0uMWZf4ZqzlWrABn41zQb09UU7b
8p2XbnarkIZdyCpWZJx+U7hWpuzEbKaR5msV3Q5Ss8npXN7l5eO4DiUFEbTMXaIGFUvKMKtj/CwM
XumvbPmIBkIERYA7uL5aVRWonalCo5q8mAwvBFso0WrY8R9v306BGb3r51hdsnGBQbd3ZARe15NY
oG1fuXPrikhEvupsvA2vBqIroKh8aR85bvLddbV1nMFXwycdXaFnh2C7ZSn8JIAltjqqDNNU6/W+
tlREbwieMvDvBxaixY+zw3Qos+PKJXmbDx4ErHijx2DIxWIxsdzmxq4wBJegvgXRNOU5wtS9Q1H5
Cnq01+0lQ3COIFSslYRnh7hOJOVUTODFsR5CxRqO5aRRr2BVv6NJgwIkSlwi0J6/kCL+jKPZfu/L
mW/MZ+BU/Eibl6kFZKuDsA9axglf15SNBvjp4eaEd7hh9YuXXOUAkcvJnfg+fxvjsSq8VqwDuHih
WkRHGjXilIvAZ5ICZWToslPbYyDYOBRzj+dhGg/vy2i4cJhqXi6mBux/VJbJ3OxxkSh/Jiw+uElp
F0zsii5hzJtFPhFgZ+EM4KidBNLKem1gpZc29gz6BNnA7MgvgdvM2S6YoCvdIen6OZES6iadp4L7
mrZfLNFpWgfJb7CtFKtIEq56WlRMwViY4Ij5wEu9t67PIpuW/WiUSxjLYaLXz4IrfILUB5vUGC4c
HknRW4uf/jp01yfT+69F1v6Uw123hOMOuFse13coirw5jSPTtQM4vV1kk/rGtGEbuKFOxpeTcfDv
sourIWsP5y7z7cIe0ksiVzCCMszZGh2efIeX7Qvz3dx9lXTfyx3HKINY6umoOHnSt7DuE7X7unaK
ffellqzpFxeBc9s4TsWBCCnTyVa3Ix21HVA0g4rbiSiehwuUQNxGA0GV6f3iHNrPQWkurhm2rP0G
kNHlLlX8gvBTO8mzuxci4vVMv6Vi6UWAmzVlUBqhNUx/0UvIKVzzTMRzGZEQukY3Qcqk0XR96vXm
7e8m3Syw3Ne8nbb5xzt6giZNmE6wo+4dmgK/W//lvTJrJdgE+JNkN6qUVy3ajkgacDePXhBu5tlq
Q4FFHBuJRGUssZlAR43/NHldgxxiexH/G4DI6aYEvNRwwCnjIWLaZo285BQiNboJ0vqpWv8kt+5e
Zx7oS0sQzckwPZFpWLD1JO+HSZKkn6fa9ZTHdXtiLO1LtxaEPjklvO2jEq76yrDfsCwdWa3pCMwL
WQuCUnyDlex2RroWplGKfEQeV74L+IkJGJ9MS2jybnLd4CMnmmLpKNqGm2tkRFzZGYmb4bxxSRRz
5bK/DswDPdkbUu1a5Ls0LZNzuWYbhRnBWZ9Qs1Q9VW4k3x7asX34ZcpBQqRktjFOSR73M55pugmD
qecXJUAR2OrmSgIIHg6Dc6ZhVpC8cX5M3g2//OZInedU7ZrbWbDVf/c0nCiJFG1jBFai36/xOPY1
LwLpbiKlIGsDHH0Ojv6Dm9zUKizb/AXCfZ12MzyJz2awWYZzJspT50JX7kaKcgEUF8wZLQjN6MP1
V1dvYKiOLknUpLOKCMrOn+ebumh7BoRdFC86Wq5Jcf9FYwOOV84z4yM3TovsVq90H9zHg+5827Jj
EOE7LpLafjTZjku4Qxkdp8QIx4duHBFTiJQRANxdpvSikbOWyGJ0mgMX0kQNdjXGIGRC5Zwc9RPJ
D8Cv2ZqGS067NSUcTgA68pVYV3MIT9ivQMsWZ6u9jWN8kdbdc6ND42G3ARKrJsaJbwAa4esLEG1s
FOQIN7xYuNF/sUjLtPsfdwPzFNGjCJqX3LC1HiKgjjBZoJWawszSKx4eXRa5InJ40pRPbo/F1JSE
PTPQpIC2ZquQR2sltn1q7iCnTRb0ua4TeSK/EQtiN2ej3NXbJoUn53yoXmhY1q0y3jKjSq03AXw8
iE5Lce4eAy1EHV0x0LSGP2OZmvC6oB0L/eav88SRX020PKOcE+ZVXzTiVXCqLUNIAxIk2P5pPDNn
z9sT/TCq8ZBTgLed/rIA422fxAIoPGatOEXfcck6TSc4za6eKs3/soQBsHWlp4avduPlE/QsHzEM
VHIICSV6R6j+fyHrhNeRd1sBWGgWQhGd/vXIw4NDJF6q1iBBDcdXQycYKL2hgGsr44T7oN1mWO8a
QV6wk/aYM+NUXt0BymwfeuQolJt45Vfchpc9menLHYqgLhSDRvAof7Ug5aFVy1zC8OL3SGXd9+fo
Z/2xGmtLyBV6vLSl2lg5lSYIlwl7fc6ebzKqrrp0t6bqwD8FJk9RvYNyDGFz+HgfzEXqa/u9hmJC
nR2rBo5SSBstarmDw/cUhwYJxGeBn/xYjdPSj8s49hI/5VtZvWN+sVqOJUt1Nzx4sNYufXKDUeBp
pOwZvLUH4+btPVgYJcVxO2QOzxcYsnO0i+uJNGL5L2rIb4fiko+B7ju3mdzDZxtwQPErmldHNeKT
OSa0YaIq2YAum2sACcEJV7B4AmkPgOw5nqRYnoeSJHQDmr29t1MFq1KDUKqy007irdxQNd3bn8Dk
xFwY3gyCmD4xw3SpGJU+c5fNuFBzL8B/S5DbeK+UYlJBGyjuJ3Xgeyz6fxFlkixZolnvNADecPBz
ab7EDBEk3jy75VAv0UX9e09GElzjkr4jDoEyrPOPdqNtl/sqcC2/VYfcRAMojYWAYxh7TMJruNvl
Wgp5vb5c5CseRmNFNnM3h6sVtPffiuM0YR/WK7CmBqS9VLw35ZYe7Zt4V55LwWv20xsP/0pGPLMm
InHqVB/nCug1DerVMWEFeEm//fPnnxmiB4VT9Tw2rL1yGzPU/fI0RggFZ9YJfk3OOL4UrHRHNUkI
yjE96ZMHzVHuk5MHFZ1r6kh2wZJH1HyBNwWXKxY/34PwfETfZj29Cx846HIdHj5h8qlUA09P5F6q
CiwT5yuwaLlkWZ4OOdU0KrydCTikcAgauwfhJqdd0/99YPjjzcKIdVWox2eu19P/DFGE9vSm2L6i
bb2vGRMRLlm5NmDZdzUSkGNkf8JWAOdUfMg6IsmvvxUPeOAn0EjKfnAyukipp8gLhikBY0HmjRT8
30m5yhQL1SaeZn2l9eFNgVwF0q8r37ZKB0h1ABPhiBvMi5/118j0r0QDyzuen8GwSXyJ8ONW4kEC
Biu6qyiW/nRhvv73AWRYbJqepGqqsuy8ib+mPR5kdbnzoQMCwyJqysy5cHCD5wtV3sxDj0799lpg
+F+spfmHBZnw0EUicnG/QtWNyGOIHhvnZDgh+ltiNgytsaFn2TpOUMq97Hpag9IKxjbAQ6vy5IVP
wfvXTxyTor2N27gRoJC8khqlGeDcgM1Kj/DrinqJQ+rKHoprWfvjynpSnbCyjpkScSvmyUvkip2l
2+XyiXQL9oME+/lwtgtHoszG3lg2l5786rVt92xhd24/nb8KlBPCVd+5xfgaaFmAacCQtFaOOoL+
x1db7EYC92B0TR0/b6nipxU4F8kiINxbkpvbKwnmyHWZa3N7Ek8+aRqAjHoJ6FQ+o6pNVpCcA1Lz
23mX+UjskKFEVijkUSZtkhwj5jKxDsenx3Aqee5SI9YjWPxWjMbaJWKovI67tct1gz3KVaIouusQ
np6fIMYN/KJs1S7orOcXGzx+A3mVPbF2OVl4fcE5/W9ivAgPtRO/NcZMa9aWXi4lDvIHD2sb2sV6
Vmg57U+RzsUKyMKvQ04enaC6oN6So6p01BWq14meOqKux6SLwRKm9BpX2ug+V90XxaXrAdXtpb9i
MzZtZeI4W/rS0ZrxL/p9JdS5q2q1/kbTXWyW4C0XXWfpYWPalG/D0bVFIn/QRr30BXfKyPW9RtBc
NQ+GE85T9OD0yxK7kCjURF/bGW1GAFxuECKjv/4zcxOVnMcg0iYR8qJJ0cynC83P6AqntGPm2RhC
lG9kBewkqx/omK37lL9fT6wKEGQG86jqejThDCT9ku+zUYfO1TU42RnyAKvoxn0Ph2OWxuuNcNOv
AEV9FLG79VNlg4+idEgx2QsDSKce0zPFhq315NHMklOPRi40lMuk/PLGo3RX+yMyTNdznsYAcoJO
g3XfdryHTpuqG3yewEXws6SK7KMA9regYJ+m77EFMORoCvrKAE7wUHmx4xoKbAmElwM0aspWH0a+
FmJvvPajBZRbXOjyWzF9MMHUih75L2jolLQjq6ZUBvOKwUj6Nn8QdwPOZNmzk7+M0CdBAryxMO4k
KNXc0zpSQykMZASwI0Ah7QEEBOdiaup+hD4Gf3+sUEVZL/XTpx9mXqyDbKDU6cuzjBHOwcSOa+TX
o3ksma9RVzFYhNd5ee5thu8G0sYJiv45TJ2ERd9r7ldt4TdCbF7C/snG+axwfuxSFzHyHN4lty7O
1b3epJ0Fh+g7Sjhj+7IzdnCk1knzPGbPC1e23E7VrrHySKN1eG/epTGprGRXmXU6/LLVLD/xXgcY
GnzhC9JIbAvLY0Kw75npM++RGdLBAZMZGSFQayb9YSe7tKF3Pp5szzByzwZ0uUfH30iXsxYmH3Ik
zv4Z1zwZkbRV/Kx0jTqTltXQHHJJ+FA7834H2iFVXUuSxO07IlI7s1NS8aj5PfUlhw/+AORjxaIN
ly34P1SAxT/G0qdMpqNypxERVZE1o/+3MpWt8u+FaeBGEkqfPCIUkR0yACpPBiKOdz0namMG2Roq
UoZ/ahxtJDLO1nScwJFcgqFM8/MNr0sgjJuibHqzB3yOgXBLLOAvCUx187zUD76Rr6ndnJdT2H9E
YT16z44OU+IFRvXF033s0FrJ+WmgkcaYoGzhMdui03asga+Of4bQiZQC/zcVyna+3u+fw7oXVuK3
z0XVkuvidRE7gpSzVoOA9yQ2h1EaxMtkjuibnZNcb6gNPZ48MZP94nUi2x/Z+nzY2ijj0V86HR/b
MhokTD4aTqqTdiXDxiOIudcfRNHCiLxNA/LIb02QnCOxF5xqsl5MmOTv4AWnktHeCszD1bIwJKZE
JXkeqIrMb/wqF/zM5v5zlNzuwQZPVH2bZCgpm1lujfOiSlPdbzRzoVuYeOWmBp96JgwwFd24Sblw
cG1N41tLxmZjN44ZqkD43czw7uL+3TdLhLwI64ZaLU9Kulk8HgK6znf3Nl306yeSOx7+DLkbbU8q
eualEDq2T1KgSXZAOHuUAibK6MLDPOinAK3tgwunq53LAhEu0ixP2dq97ZnvkkhoD7HeqiWgFeJa
N565+EqCJgRIRX2AKMLjz+42Qd4UKWawM23m7KH2CG4+CrylEl7X4WkCdEdj0/0nskpGG580E9Ky
qEITtss0LNWe3PUSTkHHtibcP6qy7/4ZJV1kA0L26R96BM26uxbB78t1EJLPP2ox18KZvfL+UmS3
GEMxLTNP6BH1Kf00tlUH//WzEssUSkXLct6h4rVk39wphKZu49dDG6La3t+oSdZiU6HoBxn5DXDf
Wne+lH7NPRuP6qUcABNpPUBAV5OfucSySOItB71VpZDlz7haQra3aIuX7OQqeWNA11uENbivjyk5
WT8BbGGeFTohe1gs/ddfi0VeZWD9G9b/k+xH7KvZPECrH9zVtuDcMhm3TOXfsVaWVpcYdIcae61R
v0sNmjruI57jyD9E5aps2QJA2jtFvesBBey4QyXkA+a4s8v66z9a/9SwgTdnIwOCKrT3rY3b7UZQ
2y2U3n7gwHihFuJMpMi26DVjclY57fvmmWPMg72G1EJQDSldGLihQT6tKJuN2iBTTUEHkzswmBoB
pOJKEfm5bM53m/Z5T9Ao+jUr8ZFfKxEzhEy1yiJT4K+NxRFVgz7DeN5BH6OOY88C9km6O6QpNcf3
3MAtcPyzX9+3MNl9LRl3Z1u64OFl3RIHDWUApuHO9M5bV69tbXguDusUyPP+8mi53JdYeEJMMRDP
eW2U6znMj0BlWAXU4kSZiGjUr/DWOeBVE9vbduRg6sbSRrueD0N9Q124qeq6zWfbEEq4/vJdt/Vt
zvXOdYUs/Eg3AysUX29dbqeCBC51fOKwsPbCaXVxP88b8Lj9D6aoABQn3BJk6uo8hppTt2PJbOQc
w/rNzfztp0C7MdC9hIgdpKPbtCA+kIPVHq8mQeRDVtxPfqNHiO0z5Ebd2atEFgNEG+PC+p3pO+w9
Ya/S9EvxL8IQNwKtqYqVexc/F9nK+ocuAMVjnulUTwGc8dFdrGjiq40v4hHK6/WAPKY218kv3ZQw
iIoEfQORxJ73dl/WdaJMZhlC34VZQEwNdymhTCJ7IMqzqq8x+nFcb2aGDR9+n3RMRFJ666D3fX7t
5ZObKkiYtbS+6X5d3KzgyOsWlS/8nAc/HUU6ZdKHn60NOELWeaV7Gz6JPuVl7veIrj/Q3W6NCuv5
z/i86FM4f9PimoxH7sMIJD3CVzGEQ6+TRRItw/42HyG084Suu3XviKcz44eVw9EWRCgTEJ+pMqQg
37pc6Qs2cRbyBpTV6O2Xldl9eKQNzWzM/ry7xigQTwvZInp8+c+EIsjbNbNQMDaE5oHw5KirBayt
T0hXYzuzo1a/tpTCpYhdiqR3KQLnjEuoNv8dP6SmM/IdtdOmiDM7d8elz5PNGX59VErucJ4TZOxk
PAo49KrUcJYN5X66GyjkQT7L4UosMMlLFB7T2rQ93Vv57XNVRQVtRXYByVB9MvrPz/r11Iaj2jAY
qKnMVhRD++NbTjIiG1xt6hZgo/xNx03sPXbadoc3wub58koenKlJh+LwL9+ey6+oB31hyJeLh0vQ
+B1NutjdHk69u4Zxc6e2OnX5i+uifCPGaFgAhcYhWqK4o4wg9ZdF30cQuLDFDrkCgPQ6ykh8byq0
GO4GYnM1kmCoOUxqkoorDJoXQgDJePAP0SyesdkozI/soLXKyJBBERurIXokuJYaZbzF4DEzAQda
VAB6nhfN7VE9wl16bf8l8U9nD+Yfi71Qf+YFPpJNbvsR2y4uaM8snITs0UQMdj6O5CwnsZROz+sJ
2GItFyjf9ldpgPZCDr2SO6NkplNDt/f+rg8gwV2AXs8sa3SQ95/3VgP3992B3I/JVZdHJVYmeX05
OtrrKVPaoBUgMV8Jvnt3pBP6hBNMsw4Wf+60hacesUbzwihglvGmD7XEZlnLT+6eJvetm7mNH4GP
8yH0RYBghQiHhuwiDh8WEeqqUu6dBsroyyVoDnv1JSOBTJaoz5+y/lCm11rzP8OuDyBSYCg8O2DB
szUWBfLOBHD35n31LRYI4xAjjnuXmHJM/LfObL2sfJDrSrCq5+ShZV7YC/Uxh1tMo2Zi8ak7F8Cu
BSLJ72u1FPRUXh3b68mYNsHiV5CVELhpppfPf2Xa525TfbPt09o1IuyjwVNxFzBfqgnJx++knLo9
rgINcawcWZgMTVjyTJh3CLqHCuwC3J+FUfXESC6qLPOGd7FbWo0OiZ+MNNvKHlHkHGLhBIAfEDls
6wNIkZfZyySRi4o0kZALso862B0t7/xukSdnmotOiDpi7LYIsYDYXdjZDYO7tfT3OFQgGDWeGy6y
MJUvPrbF7mAP0SfxO7fe+r0i3+EPk7yFlKkxw727D2XXtESC/6xodqrOuXlBi14mojuyNggPpj0V
u0+rUrosVo9HOpR2T2/io5aGopq9ndqZEImoi0QwWuEqHpL6APKYl8F3m+yyDHtZ5zJHzPkmSfPZ
LkEb/WiasiR0Xwj+2iWdpXOiXvqKlHzRPs6Raoq2511heLz8KmmV/r6dYWHpT3nMU8odysNjoY1l
w/7Y8aZ75TpiRSM9Y1JE/ukz7WH+39tHbSTQRdX7JGphS1p23xwfU9xc8IypIvf54RVW4pmD1b50
cYUjEXi3q6Bl+Ydh8+j93ux6z1KUVKOkZX2Z2VNmDVeqNtmWfHT4VtTlzc1KjlwgvP00glYOmCWH
xthYJw/W+rwqL1He1Zw2w7HfQ89xD5430MkocdGVDf4P2uTr1wJFMuAiVtF1r80corpP/nbI/K7+
CYqSxmc932e2IdxSXrDhmuQ/UBlwkSjAqeAfw9Qi5EKbEzG/5BZELXUDjeGTGp3MrnRfDWvVyeQ9
KVMYmmlh6ehKS3e3l2djgynsOa0kTdIHG8q8K4869OE1I+7QL5mZ93I3YfXzkuWJj8xo5UU5gaa0
Xf4Ycg0f0b9U/Q/oIxqkprxlm69uinweTEXazGYeaqGKW+1ySUuembpro6McGUsOWVPmK0RSIHj/
BisNVBW6+gP5Uy+uA4UDmhX7QGOGPEF6VOWis7KPVaMzWd2KLaqXZt46XZV4tGEevc5Mj2FuqnQE
6kiDLgxz81y7tBq0pCJyHvrTmzOEe02+9WcaoNCWcnrobootgWstIGQuDoyaUlOhb7rfoEtMme12
2qy7sgs1po/lZty7gpxlnXTLG0cE7F4PaPtaLUIT0TO9wa8ftY+0/SlCbD8nzqATQ7o/Rb7KRqky
RfwfS2IDlDW69duA0WSIlA8/I0+HGiyqrj2cKzMclJdP7OgZIZ5I+riTGyXRDdAzcJQGPwKOx1pn
0tTIsky9G3XRcJgidSDfeME3ZL46pzmPFKhotXWWkqT37tGRafTMNubzM1oKtFUm+s6L5wTtJ0Rp
E9u0AKQSe5WECmjh1eSCn1jZrK4TS57LY9DRZol3QbXQ5tEWg3IH8ejaGIuiEtlslat59CQFk6iR
SQhVNgQmri8u3JunaeWFnZR2Qd2U0cNuPoJuH0Kzr1fDwtArl16YTo6StaOuZJPAfBKAoFmy6iBF
jvKzU+Gl8H+Zyel6drEi81F0AYq/Ky8l8Viyff7vJ6OEysT2mVXhGTuhJTgg76Vtto+shwlIjdJq
NYb7GKYF3m2tl6aITu6jwgzhciWdArcHaGUtfB6cBT7Bh6VS/BUnmwGyP1NumMeORay8kQ1502KI
9Xu+kXXISIsEiTPISDHC5M1zH1wycYWAYwiiqFUHoBYcFpEM+WUZ8JDMVkUNMCHANZbHtuVoum2U
CAobjV2tSAH6ETVpq88ajC5reRwzhxbZeP2daB8BW2PdUpCGbAURuPj1xBhBGc1ZNNeMR9FHYwWY
tjNxMTaMReoEGrKboGghIP2sAA4sY8JozNm0h8grZqSjmEe3e3j3d8trv614OQTloVBOw5ZVSVNt
zZEMAAF+r9C96AiHtc7dUb0s0ItKXo4CE7lcUhZyebye+43Cnr4PIqDwGlZffIdghT8NFeCzZfKT
xcln6t9w/HKIBTiZsQbPzpVzVbNOmkYsmphegpBGRe1YWfmlTR7QADnDM5XVj40jAcWc/brIPUXo
ZGPRDOCcxEGgQJQWIpbB7wykEGH+FWPcCpSiJGGkLLrHFNLnNWYnz3jADGKXnp52yQa4I+cGqdcz
UcpaK62A4/ZuxDPKeCUOuPZxGkpDGu+ZpCxzXa2vq8Iz8HHaIgF2m1h6YMJnlzsPxAO3gcJi5Hm3
yCc/QsNrsCc8D9D7NaW0tr/O5f2PhOgljoAtLBD0hLWHd9bR5yWHReashcZHcwvihuI0s9NH3QYK
imb4jp1STHVOBJOc8EiObqIJR1jmGay1rvPMK4RB1qIxgEqQqeFYM6hAdl/53SZdGGf0qs0nO+a0
UEMUkNDBKNQlCu3UfEoTRpYq8RY0aZkYZi6/s6IfrbeFFKbA3947ac4gEYzHSt6vNB/r/obuK3Cg
xDxWCV9m8Kna4mHCNz1IbYCA7anGQ7NKGaBhC/REF/v6S7Tw74VwsS9MABKIJjoxIuZjTbfogRO/
EJT6VhAAnWVAeJrFr7ChP16gI9I5/Pkc9g+6I+Cl1bkKaKrRGEJTgfamr7v0FZQQ34DGM1dN4+Bf
E7/dlSFmmr41cS3OUzcJMk2BfCqhV9LilW6OMytyS8JcH7bhgwOcfeF5E/HPYRnsxMdgSi1aYEQg
qXatiq3mUsmSulikerB6V1sdp2uGT9bj/by7M2NlWelosL8k43hjLsb6SMBSRvn7qLtxHstfGmWN
M4//q/A2kNpVIGHH16XpjLqHwQzYldb73FRSdN57ZBmHwdw15tbOAtnPEplpLV4oU8B9eH32IzS4
u5H32aHmayF66IcQZNSuKb9GtdeEjMu4FlcbJ9GkKdt70yPCs1meDiAhp7gmOkSboiLHb6HBWV20
cJlRw94GhhI9B390Iny91jQZtrkX+7CD0h4smrFT6QLIYoTIvXIF0pv+/e/2bEEeLpkjJmMolvUg
PV0+deIbxpSx4SSkTZTIrBycvfbTUI2OcIFoDcXKlvvoruImfLcONEXcoWmGo9Ti2D+fNL9fX5zF
IOueuRbfABuxS8jLf/GYnyb60+CSagsc9WITu4uD4vyvpnsWboqiaHi3Q0ZYY4mWhOdIGdphaReZ
csB3S7nI2eKmMxg5vPuH11gwcaUWh68vwbOxDGXHW5hR3wEDoV4M9qwnpvI/84jOAESluYDfRekF
OOz/MGeMOuqWW1gKYS6wUTGbDlHCJSote+QxCQeHbIFRdHgU97A9TGxVHqWLQW9JwK3jRjeNACpY
ztwK9SSm+F+zxA3UeZQk3jg5m7z2nz3HyfX16jaxJdWDivy0DZ5/47Jsg9o+q26Am1xDRYzmkXT8
PlDBJOwASqm4KR6sEVo87ryN4bjcCIrhwgDrcQt5E9Bj5Jj/CzxpJVXVgkNWTcyGlX4RnG7hvg3F
a2Pwg9fKb9eDmPCS0I+GDezbcRiSqgsZD5XYgMAlAjb+A1w0GgcBosAK8yOf/Pe13NmG/+TZHg3d
I3OtlMHZ/Adsu4B5UEK+khdJDqIrLC4T7FVQA4NRnFVo+fWhWfJudhIEPRTsDFB9zMRN/gipdrLw
+7NfiuppH9m9APREa1xOQ2+bVTIFf1N5+STiXF+Lu7YIKuxzFnEqxwOnu9GEcEcFvLR6XVeYQGeE
YUCf9HMqCisMQwXWT/5HqzcKqEb5BycFHrwNwo/avScWvTff3+RBaMRl/LYudQcxLUfzf8xPwf6h
EbbzFu+RmpAWHpFzhKOJbwZPFhNqVuLREimcJMSzadzA/OAeakafplWgHWDA8extfkPWNFJytK5w
yyb59wGj9yutBOBp7GawnH06eTFRm0pWuPX93iwXZRAmi3osgDm0EX0u3pEhgiKasEufeFayFsgF
Lb1Ya/1gUBaywUmwg0HvTWmh1nQ5J+8VklRcEdfL2sWEuJ1kWcCZiVkjvv7oGgUcsYmFKPIz7MKA
R28Cer44f9Kee6uHcXl03y8OO96277OmweQbCtlAtztD8O1aMGGqbR8XdKql5blOg1HTLLqmGYuZ
6PQ1HpdhPPdLW+R4NloyMZ6wqL4sGP2j7nKs17hBZmxuL9WHCxut/uBX7zhAhbbjnHpuBPUW+Kvg
muw4MpQgn6M1ImGuGaK01ew0xpMUreC9hg3p60dqUDkl3hUTBJoYqPtxHSw3VEQNgfxw3EEbiQnz
9snW3M4fE5zCCGZtKpvUyehLEr+D9nm4mY7A1rFTogF7G6tXlm8yeM4BgOgn9uKr8wGauH7mYaUJ
Ydfzp+i1fjmUURfZkuiUhFmOieZKMwnVbM/j+Q0+YpHj7DOVDQSDW7p1LLBUv78P+aE3W6TjpNRL
FpEx1eOe5gm2Nah+b2Y28pePzntyrX7uB9F5XD+PMap/WmPcdsvMOowEvmHWgrvtVqjDBwsCzOWi
quqr0XWislpslj9peshch6F8jhK+iQ0aqhjYBpNAv9jZdGQD5uWKsFGVataphq5U434x/Xk34YpM
Lta7XMD7TqTDCV/5E9+Zf03epMiaR7Y0eVrPmGIlXGeR0HpEzeEDE74QxX9YQOJ7dUO6HC/8ywY4
sEaR9DLwf/9akyrY7TClV7M7XzFVSS9bI0NM61NbRhZMX90QRp9OahuZcnebwwkgadIEoimYuWIS
9Dd8RA95my1ALeY5hYR//CePLNocxlLYO/f/85n0qfMUhsT4lCzFXMKvWtSrmZ/zXD2D1du/M1Nn
q3EzsEacqSkWhkENyGFjxrFN35AF552aGGdjOCf43c3DrLMs01ODnttkfQy1cFZFFQ03Ir+4WVgu
D96wiik1R3YNVM8EOqlPUrFvvPt8NJcqGl3MHKnEVbVB2kzbJFgv4+g+w+4kflt0LSEuO/b4ukRN
9LH1VMqjRivtk30vvRb4XPHBAPolVLNLMUJIm08ziUHvCk6DhmcJilExSed9FUIf8TDEVHMMUAFK
+UhyaPUxPnS+BWivsLcOIMvwtRC04YZte7aPb8Nn6j/LtF3MRX3TKi6JI7DOa/RPRgxnihe0mmRH
YXe2sedj/Iwm3hfo1Wr/iPfdlRp3rQXJURv2nzDjSdnGKD0U+l8zdI57P0n+9hxPwkjK7FfcEaG0
0b9uGov0jad/Pbx7XKxN2HtQIjk/sQhyCnDhPn+ZmCdXsYQDmgWAkIQZ/r8Q9DZbbXpLoUzftCcJ
MtGK9h6p1evBrBYWRed3lziM/MPA1pYUxj9aV3bBQVfEWYpbq6zBWMEeu88DpGASJ1/PUHq+B9we
apAQgAqfPGk6d1C8qJ8dHTgsnSSftVZFzKpwkzA08B7VYvPKLzBv4kWOqJFSOuhfTPuACA1SKQg5
oEMb2MqlIAg/0o3Bx30D7+F23pQ1mKtc7/MCwNDVy7SlpztZTGvkbMYz0OiV7JTc1u839efryiy9
0hcP1m0LTwyo43jpTc/x8UqgmbZdgpDgysL46g3C2udBhzhaySxfb7b1L8EG68wdUxzr4NcHNU83
NSkvHreGWEMW7xXn0/VdacROQPA4j1I/kGpO7Vd7evzfap/OxfBtdfEHh6UiW7Ss4xjsXHdTRoUk
jEKp09wMTJ3L2uvxDbbdgVK/06fgTSUje1Fv1xxn+9BDWiCCMJcr255f5aWfEg84EYXCt7japSpR
iHX27U6tW1b6rR7b98hctUMJtG1nXYP2ybZIjLais2zijIOZADMRbqCBiXabcDDuIwkG+yLRsbI7
LWBJ5kTwml2e5rZrFSopA5g89FST1wtd39h9BoonUoJmLH2nXFTAIVK+3mdWxljqHvqiOd/b6NSt
HxoYZv1bhc7+sVnOmpeR6bthnp76D+BY6BWRWCGQzzLJBFTuXhR2sf9lvuiS2DQFHG4UY0qH0zYE
Sm3CYtVf6HfXMtjaaSOdDlJdV7tmmza5c6CBIWZ3Q/CpJNH3BlqSkPZ0hp8BAoaf6vMerzHXVvUt
12fEmezzn9elvU+tdSwcZM+Kh3G0uUKDWQf3miXl8+Vk0dBbbxSt3t2gruis+DMH49aVMZyOMfOA
NV2IB50sNBFoEDNqYtvEB5iUnlcVF4H71F5dWz/Je2swAp6buxthz7x8S1ZPPUTteX9C+XmDa+px
R97Mx5p/GT5k8XIq1uRQdY6bEaYQyYGMznQ0v6chAScbTsy0wFPEwHq/Glmr2vyyAjx0Kc3cCkeK
ZTcIxTS0Abxn3aQXFYXaBpksUK9hrQPoFK74LU00pZS1TtDubYurwKNb2hZB5vtVsuhR6B7Rx+co
2zfTNit4Q5fizV+fUJ8V7bOpI/XVSCiiCZkVvW65i6pc7gHOOyLJHOCjHKhdNo1L+1+XD1qC2B5x
/w6zCXVw976uqNvOQIJHPnnx3uytKho6pqoNyNgMaos8CfnLX+W5sG45kwjNCEjOKwZXULtuseAa
6qy6PiPoe7XvWB54IXbkiisWiKcrVZsH3L6MnVaT6cUEJKlHl52DA+Ag5c98iyi+Jh31JXJVl0wK
6IjbBvBeuBQKYFDgwCvEVFGyALv8mSvTVTZtmVDyEMjY0HXBBO92U+8tcIcsUShsBNB4/ES/hP8e
CzHJkhz1JTcu8s2ApbPTFIlAvnaX1q3HEx8xQM+vYak8Wu0R/xFF/TOjO5CTEKChVmkm/AFSPbra
Oe9ujpWRsCotcS98TFJyityLBdYSO3Y5gXDAZXoS/ZE2MwtJW1KQR88gOD4w/080OtYRfpD6EMyi
vQNoJGPoT+Am0ZkZ91wolCfByxc7YZxe+hxPODCtbL1GKEzvNzGp4JCJQOavSIq7pG/XBvzNnHH9
u+kbqYP1zrVSlgPzbD3eotP/zjVKTmiXzfDMOpB4ltIeFm90S8jk2Q2InBrWEfYB0mHUMiYuorU1
ZefifCOpTz3jfDCCCkEfjUvtFjQCtc3qUKczV00RgYBruk4V46bTRJyrw+SMrL3TnZQXmKsCVANT
sm5qs+OxxLtpqLt6Nt7nYcelH47V8qvuUY+bNPh2r2gn39q+g+bFbqjEMkGcjJVMuLg4lYWNhxG4
WfbV87ZrpwYp22S2Nq19aJp013p/loJq5w3yqpQf1Z2zK8sOeol60JFCHTv2dF7snZgwjOAEN4FG
Jq89lIE/HtXFOSgHtHXMHvx/2GgBRBZSFh2099QHvdFDIcXmL2dL81p+uLje5JWxxuM7sVwR9neA
CAUhdpTUiRocfIK/Fjsm60Ic+OgPyCcbSr7icIIW6RZui3oVC3b+/1MnGvr+8h3olOejbKX/d9rb
Z0zlOtR+K3z1Y2HeMVu+aQpQAGJU5qosKTCC5uNIXixVHnSSgdOVjHOqFl94d0cBVy0/E5rwVILR
o/0P5/h0N3nNpOa2/JPt4QL2QfzaZXq+C4AJ7oqYDU7ojZppNK0gSqqeAHlm2OLaBTttfLS8xl4/
992LCu3jiw1DTotylfuOZwHbavaaxvuT8Wxdukb2nsSKJRxznZxc4itZ1EKBLJp+ErYSdfTg4RTR
ulI2dKAOT5ZfrPvjNREYixvl1FxmlUwuT8fUuvLdLPSyso/A6IsUFhSyySVF3osm00oz3O/hkgWd
xqwbiCMMbLt3UGdMeD6WEmydqQeFTdXutmh9/Sv340t3Qbc4eHh9eGWGEeEJOJCjE67sbTgWQRoC
MB8jn+M/+vhXeVY8+NUxeEDsSzYNr6hDN2lKPxn62U8ffrAGAIzv1s2y/G5djQn4UpxR7xLbekij
nyTpWPKD7BKVPqHMt4fGAFcecye1hzkGrHeh6FmEWYuoELtT1vuq4AZdNFvOr9BrlIyADh66mQyA
NSnbP09BshLBy4RBqH9S8wg7Q6bhH/Q0YdKO7JyY5v7wMR9SrR+iibnRkdDY8+rao9eYFoZE8JB+
sgtHuvA79vHWu77JiUiXPtTYKMXL85Hxyc2nyFnERH6n8h/eV0ktWlKI/0IKI+hklnSMd35vwqwd
vD4KLdPr6oiDcFnPuqBcIc+HJwzEqMoZX6aVa+54cFAPqORPp1mTeXvEzofX8feAzjmnz5uKcU0s
CqLbVWP/jVCEOrwM8/X7/qQgA+5ITNWzZEaLkYgMKs/F9TsZGJZCYIJbojt7Y+PxO/LDPTtFd5Mp
ijMtUqduMgkGFGPkEW85yAPKSIjpBrbE8tQ1IHQqTElr8TJQ7z3nxdG0F3ByDvb93AmwTG9FOGVN
IUEN0uA59uFYyjlC27rULCYpNfa26k2V9uz20UH9WFyLMV1jVP2i7s9u3wbdsDwSLoO5y/1/cPke
FQTIH2j/5enSs6AVLAx4nLXF8LFk2f8synynJJ7B098Ce4CwY5eyiddylRPzoHJT/MVvI3niwdLz
oNNe0rblRrot7VMBh2vH3vGpIwSPkLQZGhL4GPkm6ol9/ggtwb9GAX7hM5u2YAFgyyI4cvvO0cvm
itwegVeS90qP6TbilyAun6m3UEqluDVWqXaT85uQeF9qOGWKBvGMiGrm0C6f1mqkw6bSIXkzvmTp
I8eW371DdLk9uO7uT/1nHIW+jFGNEqK3ZEsTa6qzGHKmcMb2mKAq71MxUDklk9NVsLpttKFFUDia
4+B5w6oOqsHr0i7AhPc+bsL3iNOUtODl4mu1C6CznJtr27uMCJ+mZ6uFgsrX34ds4A9278XJelMF
xEjTUdQBa4b7vfxvIrQJgZ0LkhMjbu4Y5ei5gT5MUbQvKP83FholS9odi/VMY44ZeirPSvz4ruuv
X1uE1pTTpJ2nnBTx/waYlxsPOTwdfOOEp8Hx2ME5A2WjyBEz3KamWQpB5fZewz7XfGr1rSBu90Q7
6XntQa2EHXuhJ5OdFMga4cOi68YcHc8x/7BK89ICcpxVsrxjv7JYH+KqB5J5HUEQxtKjLUwuQg6v
dLaL78PvsuYAsq2wFbhqeYAfTI0TAkcpntFEuba1n/qDsAFp1IRRDo3MqCH65XQUPMgdYP8pfvyu
Y8zWRr3EhxDB4nM+p6qC0gXhTWCkWLdnmmnyIUC1ryvxSXi2qwhlxJ7kfy4ycKk830Tv/QJta6x2
qKAgs8dVUoLi/DugBA5K7QXFPuWFq3sI1bTTL7Luoc8QDByfS+4RiTrHo/HRJ7vah8/z1NAzl6R3
s50EUEz8LPZm5NWey5M26gBXTxx434la93t2nGZPkuLPb7BovjHNFSQnl5YPZyLEx6L4AWx2v5mP
Z2WEJG+CN2rv5rC6f0rqduXCMPaWnHDm4uWA1EwST2wmAyESGWRFr6t5/tKvfS4ejFHfnKgb2RtE
Uan/TYrR//MxoF1v+XKmw/ofNUvs4Wros6pM/wFNleoDxPapzDKzcKui/4OfNIgesF7UgFKU2nrU
lTSnpKHukkqBtKucsCx7fLEoz5mHGshTLzpmI1Ab8/4FmMHTaDQoSB4QZTAQNHX67m3n3ZMgTSZk
7ldpU7BVJYhCw/soGLws6jwq16EMHQURQPg/ujGc61jOyNIrAIoVg+RKeHLQHb+8prUsjnZlD2vf
SiiC+BREziZrhTXlhWIqhHAozhniIzYe0+Ty197n5UQpXjJBgbOnmK4LuabZ8FbsFUd62ZC6/jV/
//7bElos7gWeWBmOsiacWYOLzyJpHr3qvHtMvXGieIp9650zy0ZOEcj5HGqCHKqPRbboTGfjcWbk
oEU5S154ugKYWv+dykcoP0807F5Lh9a+euvR+PuDP120KkyTuNob13ywhSiTaYTj+w7uRPT1a+p9
ht7e5NIEz5TwZauEXMR2+xKbLk7SPoxRPyFkLJ0aGD5piul3uNY12U4fTyMMrRT3ti3VVQjjCKOo
crg+5jKiho3uoQzPcJhk5FO5Y41wI5kCga61Ytbe983EDvnbKTMjzmpO1JcFETwRB5GA6mqsNISX
bUofh041GpfSRTf3TcmFls46TEyUw/BSJr89aS5Z+P9YciwaQzU25igO0PoFObIGizktzzOZ7ou/
vzzUSCn95b/XBsUXJ229lCnfwZz47ZF2MIDtOaI4MtwFdIIy8l17gIzCQKVC/wO3CMiRGSlgVy8G
NBz4F2D6q3H4ToqYQrKNJ2slT9sBbsNHHsC1QpKODrIJc+MsRyCC2TJgxreEEcCBhDdQ6Ns6kO7m
85bwx1ulwgsdU+al6/oHyWvxYfPb5ZiS3oJ6NtkYbZU3FmmZ3VOzydvTpcR1Xs+XbTxKxy7y5EpE
fI9XRqvcriXxsTplUcQx8KtQmtaMzqnNv/ygw1KEsnw9t6r1oWvVJXzU35QOWFHEnq+dT4Ke6+6J
cPVD+Eh63/5i8fEW4NKRpauBuDpV/BqFa58OzBpRqPj4vzpBCuGA4/okLcdSNV50YL+ou5i65KWy
L4BgAQDfyQO9VhMX9quHCm7uk71lWsl7/JcqBBkF3KXSvfAqWSI+4RdWX4MA898LOk712/6cOVUy
4YlDRRVwluUBlQXVUeMKV3oe5bov9tk6hXltkOk65RgdM5P3zRAzJC1b4oUONC2UfXG8TnzgQ7fl
QUUdvANcLVIpDbcVltpXXiADg1tPT22ql+0qQ3dRkGHoEHEVoQ5E29UaF+eEjkuIaCyGKgiwFSJn
AoqHCmsrCimESLyGYkW1p1eWlvz5syU0JzAsWy31Py7ElS8tmzqFWg/rDjYH4L+OxLhvyzjg6TSk
0tRg9/+p5qbHNqrQB4EpK4sot4MJtm1eZJKnDvax5aOpJbQ21i1O1Ne8R3F0DKDwu2TFCRxejSNI
A/OqTeiIwud2PlKQOwLCqDd0r5R/6sC5jA1+X7j32q3mAphh2n5LQPRXx9xe/O9q97oy0fsmnKmp
BHf/9fsNeHRIN38AWJoMeC+TPClQ8tnhFO1F42hwA4sS95FovbCikK86iCLyn/J5pU98Rc67zX+i
moSP8nVD/8HXyWH4m+QPZVd34grshLw1W9MK81VPirrYkfEFXZ5KaBTATYCdAXNbOL3UTvvd+T6t
T/E9FH/1IwmkZLutnzSyTdPH7/Z85KR84IUdNz37GlZ0I6cpFBeFGbqjoe6J0cswG4OSau4Yc111
oXFNTziwOzwOYDZNlbwckO9HtryxJU4b6s0EGfp5NEAZrOJXNAyxrYRr3KoDPkdePSI7lp4fW5Uj
iyFf0jQq8dc38uuu24u9yWs3Eckh/2NqUDQL96CaK5iOozZHPLIehl+vQTCK5hHXq203kRUVZtwR
CB+t2Vk3GFk/ZxUb4wEVhGwpVXk3lwgWZ0IrlpxXTvWLDqBoOaAUwshjpkiUi1qkJ2AAWuCm6r+V
ervIwIspe+RormMISIvtdiRLpeGV8EWa1aXNRFleCQvBDDO9Bxw40jW+2sGxCwwjs24wHS5CZKHP
f70wX6Kp5yc3Yhy/oiBzXwD8eH/1CRDmqVqLspXwza9Tdj67rCSEJeLHt356jaNu2s7kc1VrX2WV
yHyP7s24M4cpYlnHueZlPoUnOnYQBCDKmVQgppLwD+n/PlWOwSXYc67lXYv4o3QfAjRPOzE41bOx
/hPrhqj1EiRHxK8POGH3DTadDGCkIDmcQtL+0+l/2uuBL6msaQgUQAGvzX4VMkz0kP4D2IcWYEJK
JYr/SHLQdUqrrxV/lTfXnXXXTpNBMWHv5IbCVRoF3DCMBiJgndIqJ1T1wWccU3VkX23SdcXI/FUG
vxDSDu11It0XSvWFg7AHBg098ZY+2aYfYCPcKPMt4L6eK59CcZycRa3lYVerwLV2ARkEd6xFyzIl
aWKFjj+xRecyyaFh1OJHiQu3pcJavE5lq3t6OWXk+KgoF2yTZtLlGESrd/SPRIaMwILTMG/pcSkR
sGZeX2f3e/gpdAzwHhPS9QuUAy2oKxcEBEgA9IsYzkDL/lQb4HVz857q9Fh2WwVRoQZNAn1/3uE/
g8pjoeI+AagI7/dlzJ7nCriCh1PFwOlIJCpxQ3kI0PASUwtV0XgqgODBDk7AeKaL98llBIquUIOp
qkM4STSE5BIu9Pw3dvG7GCgEIRzBIB8AVMYpI9RWTjjFfF2lWJguI8pcTy7DZyuGLXFI1Ee7NU78
LpX53nVCmxSHS9dmREUjwBJQDfCFvEqRgYrpmQqbZ5NFpbHEA5v1G6P6VxdU47w4t4cXWXQvfaru
cDcpsE8mPiwe+8fxLDVpkBin4fEUzTdzJrPZvZbLd8sHLVR/tdW8VRXy+xuiU/1OAneXkqbdUbIi
CVKBEx4Yy9tP19VzGaB6GXm4iCzrUVSn93/M22IXHLczYLdgSu8rh+p24r2rjCsLQ7AqsLgKxp54
6vmcBoYIlIKhvoKb8zRME7aGjrf9LGX61Rcp4DzMwVb8N32mlEDiZ3Q8+McfWGYcXyZdOK0f3DiB
eZdIKlJMpG1i7qQPofsdv/pCwvUF/uKsvgQ/LFhZ5I/ZsIOohTX/5lnO6tnDWwu1PZ6NrIhUAPhZ
LdqZN0IP9fsp6JjJ+B2URhhD3kHkFhk3U6ioWdP+ewBKg5drKibptIMOpu8X0OkN29uEaaQh288W
J1ekc0uoI9eHd9rq6QhrSvCBo23HDL92F5sLUHQGzALkf4d50DJ5Lav+TwDtfnZyCw0tZ3K9rjXy
oGEYWrP3Sem87gIuYmESXTawJ91ZuKWNl+zfUIA/utQBydncpFcHpVIQOOsMAnIzWBck9NV92UCv
YkgYQuG+jSnNRUhg1msN1qEmCvchpPg9WNqsZJ6lFPVq1caS6girMh9QyGznUOi3lReLRmySeX9w
eX5vWS84If14IFU2PHykLCCYE3UfWXgdMCLvLW5V6meRz1j2bZSla+HIlEYH/SpdV53y/l8u5NJL
VMal2nst5y6j90wFQOoFRmGD7kXKKP8pZxF7fehMhNTNpiFv5v2CE3QOfJUvlDi5iR4JM5jR4cCe
hZrbrpj3uuUMs5oWHBjzMRdu/fmBjUBwjBOczRycOuy3B2zSwNwXAug9UqvXGTnbQ8TR61S55y80
xPmaUkWXw1k8iNXdqDyof0SbP7IJOfBAKgJzxJEsUwMr0oDCWl6LV7G9bAcWljvr0htU1g9gv/Rg
roXJeepP7GCYaZ2hfX/ze0l45Y5ISLJSzEmjsJ9Y/dSTjIGGjnbvu4HStZa+dvk/ODiYDteh47Rt
9PxIUEpPWwmHcRIxSzxHWVuI5wuas2o6mOp9qpZqsFF+y/G4BFQLJG3D5D2MCzcQbkvRqABKmEAX
zRkY7zdFNBETVTdzspNjfONfwAU0PPv73qnChRLJ1q8iuVW6OWgyYnQns+4wRdpVrMlA2Yi8/BjB
iv57B/w/OU8VeTAtOKJVvTP3ZjwRlezSSD3fOOCnqixytQ1YJAyQDFnKbAedH8AJMqlQL5cxELNS
1qQJtaYTFZaEAFunwxU3sJ/0Fojf5QSSh2oH2U7eVllZBUR4jdLvN/xxcivYoOFa4UdyQvyV3h7t
Ze3WH8y13Dh+4iBiT4db9NHByqhDC0mq1uxSzFOS665zMzqIwxtJDUO9V/CnlV/PDWdtQ3MoiPqA
8HfwqrSW1qHCSDQmuGeWG5B3IXTAXlpFOxqTyANUGDO7mazxNhSH4htzGQixs6UDtpqbFflkcrVP
y/DdG1uLNLLPdtOrMmoczLqa/4733u567yur78f4XyIO/evg0H6oz1/tqs53/gp6FCmu8NT9l09P
XR9MHgeTV6kocQWmx2a2RlH38WOuxxdEuAHOpiIMSoUKuSA1ZwPJ0dJv7z+2Cqw0P1m8Xm6OqP7I
YvTLazvdNdTvXH8eEitx1fa2+uwLJ87er3FCKv3slkJ9dwOJfqodmGnB6jnd9XpLs8UPnvziqtDj
XbxpbTKBX9O0zDvgfWJwRWdeKFHGOAhlDfmkfc2zWCPo0PAFH1t3Le1vyd1BLP67U930nujPM6X6
gSEeqKcAV3gZhlGnsbY0SyOJKCf2k49TiazI01gOx88OmEb53LDmU1JEc/yEKiflZ4oMRsIBEpCJ
g1SRBfuPl73AU62euCCAo8pAU7hxJIR7l26kbVJsoHsMjFyg8yuTqDO31lj1uRKITnPgOofAUnyQ
/QkzToocOCNMP4elL+zQ3bhpD2pzjVXLGedfYb4+55WtY1/dTS2I+OLXHB6IOTlLlCOvdITbq58U
0nBcAP5k+L5AVg/DKGH/FEZAxqOcV6dNvflrvAsyO5mcOkwcyAbSXudRTTqb727gLi6ZxcD9b1zd
Ee4wk+CBuIA7Umzw9SDNesCVvPsWiCs/SRY3/R7O5FdWh+UyCcrUa00IqqeA4aHt/ia99vbbowRS
Ea7D+fZGWqUUkaUB9xdkWcTnIA+87ke2owEKa3TEtB3sOjl9Ma/2ypWsEcgQwI2AAAjiERNeWSaK
fZiFuI8SUcKqGecl3gp08nzc/J5UODti3o1AO9I8IBZ203pCLyAslavRvFwIzT/LbmejE293nnrg
hhPVhapjDhUD0HjfkkFayYLvt5Jd2B41K80LZytE8VxilkNlB/hZktiXN2XAX6IU3K+u5lKKGFL7
ncDovKK7dsRTVivbxTAA+FtcTQIfU2v0Zz7WJI4TUxdr5B1CEC0DSUll8rfSVAEauAn16oomg13f
Z5W7tN6sixICdTHqZFGG7X7BlJ1MQBigDZfqBJH7pohdmE8KLx7go5F60EcrQvtBd7EwWzEv1ybK
3SRVE8qCvriZHx/B6DDH7Tw96tLxv5rj0n18JtvIr+wWVIF1lv+SU5HWbAfEQPTplu8d1SV2Oenu
tw9RlUXnrtE0NMHSumERGaspwnNQ/ywQ4DBz8z1NZxZzXOmACDu97I2gB+V5qpIArKkN5EnBIl0z
Fs1tpwlOBgOooEYe9JNJI6VcqEq98ehnT9phJGVLe2dqPXhbmAU74zcG2THM+OppezoGa0OEIHcf
xrZng9ik3tdpLbV2OJTZBUIvm/1ZyrWX8ISQraD2O2vGf3kFBWk13UIOSXlY5gUuhb/psVz1xEMP
zxwO7ZF61yFlIijZf7vpy7CehAcXlJh6KPE9+7japQymaELjugBqUrXQ0lrU94T2p5YQ4hlNe6yp
R+3vq5hy8cOQAwV5nKwM+T8J/KeCz4XFwhTktOgEdw3ViYS7GsxxDCwqm4hZ+jRCqp7woBGcZeK+
7m+tiy1p9x2p/2A4mmsU8Kyya9ofeCdk08xBWF9ckI37a1E4FKtGhgDGOScX1bxuMp3WlofgcFR6
wFqKZ7DEs3Vm9tOCPM/wFzXKI/4uIN/Vm83ui+PD0Kpepcv6YnkCoUoLyy3XKKMr7ywTQ5agL99y
ZGoispKOfMcwwuBBLvCV6Iy9Rda0Hsyo0gWyNKOUQKQcNcSlaX8DK8gUey5jHxavfWZyMWPqlxgn
e5xOnpUPUNwht5XJpqGrOX3ARE3y9e/jYrAIeZgsIsuhSio/FyBEiwfpOAzLQz/aITypFAzMh14+
rltCiO1RCw1OrvwqC3Ij3VIzUopljts9ubUba8YugjhaybVO5L73EIS2o617pkuQOA9sIxei9uZD
EVVl/Y0gXxGSjJQPV1tXxIBmhaGw61tpFBCXIZcDFHSjnjrN2p7CxU6jWzSCyTdpfnbToOKrhRo0
DChUNKRNvZlP2jYXNaqhZaDoBc4MU0OSK8HopPL5Awt2n5HaDAQFBt8YLSNPdQiZZFs3puNJYIUb
z/jY4ETClBz2uMVr0iySZnYvgdgGlFmM7S/yRWwZx+w5BweMWaAHEXS2TIDs2zCdLVIwsD5UagJL
fDuYY4x5xQ9cdJ8646PRUAJYYRUARoNdH/XMwkaLpId0UZaDboQBkERUhr8A55+L38bxs59g2/P+
PL5gvLRb9hU2denxt4/7pFEeTcoAKawwc2/rQWZ6zfXLUSod6hZ/Jgy5/MT72X8xyLiFmouWdjyV
XgtDT5KITsU5p6TeXe5qXKpQDunqHsOhibsRQonXHVNWGAfB6wR4aFMF1e1HGjddeiggaP3AVZwD
xD/Oejat/OpE43E33SPc7wZdHRz4Y5lMQwhjvfJ59ypNG/dAmKJ5/L/fBedFmxLkCRPIPFiPbs/Q
SfvPLsRKe6KoOdhrT1lYPh2OBjv7oRYvsZkYsSOhn+hqXee/F5sAMYjzjwqUKNIrBA3NoQ4CKPSS
mOpp2xEZffGDwQ7lvYX8lMVSWq71eF+3BQLTLSx7vDfy7YDEQgvld4enTch7vLk/fBwhydA3gGNO
TgflGbDWmsDjlpZHzyBsUjiZnnkOocDbB1O+9A1RPI4L5QTatZCAG2L/Ea252jLNJH8K5NiDHXtF
NI0m2IIAE+NTEhyDAvOxBC5nmWSfreV/xcdGLRAOd3h7YejENpbl2wA7mqnch92+8gZjASnm9+0s
BV3ftpYFXAVgau3IyLdGzHHt6hEEZFTVFhm3FhgTTQMXInQrRPS9yWne+8XNYeCKxdWfEBevPeXx
H1MDPC6YLIVINc4/AEDxCV8COzmOC1VhUYxBv3Z6Lx353gIW59uw804V0UbHTSq+BwiqJ9QvPSC5
ZTcg4QxTwp4R6HMhbLAJqDtSCoVjS49DfiuCt/gbIWXdw0bGx0vubpOsfOSo0Q7Z0MSkjFsh/b+Z
KQyIA4cUSl4jsunuMHi+LaQZBOZxM8Gn2LoMVAqZDCw7mj4Utji+4KLLYetdPBaICk3vFAflC539
G1zQXYzCC5wF9XK47Olehi05IjRL6z9bI1CSilykJWnx7b1xIWv3qCYz753jHWX/sZHNPYm7s9hD
KEbTOFZxcZr7tq7Xb40ed8pYf6vwo7516uW9OSGI9RsVU1tvv/Myis+bTeHfk55PtmALbiO9NmaR
aA6xtLvpylfgAewZJrv770RXo2xcEkq2mDlaSp93isnZK4ijrl2xWH6PGADKx+4ZAXLfR3DZ7jDl
wCzbozTHMWWES8sX2xNRIuLQhPi2WCdMPQcfCbChB6WTF1qY25MjAqaS1OXICo/WGVd7fdczaomv
b1ZqJitJ0kxzIlkMPH83vTAM2Tda1CA3s2yyLoJl1Jvi5wRen1DxlIBVU4zvNHkzAJX5Wo6wZF7e
X313ac7JkkrzEwlkwdjzFJ5Ncw2DVLCq59ymvtieCsurylobFqJq5+oP9OXnlK0XYX1zwZ4CAmKh
+3rIFiyG4qtQM9qxVBNJ31MHimODpYMManM1GDsdbVh9seZivY0oOBxsyTqAIuvjSRHXd7rYTPKr
5UcrPYhqtkygt7yxHlYWrxyILcuMCswOVQoB6WU+LQIHyDX5aqAstAYlIgrxTkwCqX5fJaf/4nZH
mCW2U7PGYF9D6avEpmb2nxGmR0niHl4UNOVTqVpm1nh4BY6JFViLTvqH/9YUhIRSkyChHejlyiSF
u6j/sGBhQbnEqU90pGqm/x6Un2GnXNGxqMoBcsdTViQfshhUtwGj2R5kQTht101cV60hUOXLMOHs
mOwz9qUicfZg2PkBiVzCr6tK0CUb3f0LiD92dK+fjsOXYN5S0KDy7T1cTBV7U5eQSlkkZuUHPhei
E/J1SSIQzH3asi0wyQA1wpRKS/rPQjsYzrVRNjlHL7xf7AVwY9B4tLAf8DvY3fGIQjnThgahxcLM
hroNzzaQ3zhjOfmELodF+D7pb1SJLrUH3FSQ1GX/l9ecnz4i75FUZ7UaJEQArx708H2eBA5kCvTl
FmrJ5NprLAQO5Kkenarn1clTbEF+zctVe4WSftOtdL/hlLLG3PFPteYjGFloa1eUN34xQvL/hcrJ
0qXOgh8bLER+SkZfFi9K7RGgqhU5ufl8/fpSX8RujQPqsWmQtANRqMCCYliutpu45GaAd+C5scY3
2sy8mOdl/soPOaIDb94NHdcIqqZQ5G4rq9W2W4df4WnddFomnxbSm6P5e20VaRoQiHUxkWgQNTcB
Ul4bWmNdQcEwxspDmcCtoukXSACmFCEmecZiyv7xDfYxFFeV2hbSt7oDfNkAmM7YbrfufKQIgjGV
CpWnWeIOgO0etraXlqsDfTzQLSpm0vHDiBqmlOojnqj3sULUU5/M7esagqL2ppDGKIgpmj1I8P9K
5ZxcHaK6XtjffDxREy1UodUD3w7F6nM9m1pyhayWbphCmP7iqMlMcQdmGudgAsMzM4lLVfac5tJX
T9q8AUr6C37W2w5f8diOaG4eaIOAaQMLo5B/U3nIORaZ5/bWRpDAvWHtlAvfrwhu1mZ8LMKiZ+eE
+yVubf50N8LwvQCZe/GGD3bAtiogkKlqT5PaKYJlFsThCQ4bPvuNRlasv7UnymD5EWlYqGUn4+7E
PclB9JSsU9I2nvddac1wLhF9DpmXR9X2UlAAvRnZw9A0UOyjYO8zVf4d799t1LaSOOBPN1z1wolG
v+v9b/fiY43Tixdnv7t0lj5LmOO+UIa/nfksEejvmo0Xk3n3nomHWAPLZJlS2xaNnDIHr4Syc5w+
M3yWCcYEZahjOEiDREzjsXf8n9V7ZuEqg1hm71deHsM+8r7qNEg01+sCGKhdVP4HVOOi6WSCmphl
+jHBocTkCaaqR8ck5Td6PpWChLx6zL57o4ih15YPagAqkcOFTi+1Bz3Kqs5fk5/+aBu+3oKoEqwH
7DHA3wqpokeUCps866Xl1IAaaUfiGUb42ou30tZn2MA3UwTN3NQOWRyaHIiPFtOrb92PrCJKZskp
EwGSHgbPBg2LDF9A3JHnW54UULw8Sm+vsBsA45HIyFbl+ET08/iVbWwkLctrKbsWsHTPHf9RqqzL
oapzRBztuS/JPckZK5QOEEjSxuDJQb2UicvXTVCEqKqvGrXHUST+Snt/7nR+hefanAp4LEeL+UJO
CrF1F7MAsL1w0FsPCz6EBQHkJ8tP3hSmAV5rxhVDCFJf38DW7bnjTzm4vabxXoIwG85ljw5KKSeJ
Krn2ZnLeKYa5nSnPR02YWqlG8h48PeSyOQfGOe7LFWlboNi2uytneuBwRLV426l9f2Se+CGhLG8t
tXclS8orV8hF4TSAUGKnh0sGzuCqN9bIbCjJ55XnYHNgbPZ/lXC7kJOEuy8aoWsmVk+EYu8B5a40
xNSnZoDsMz3e4X+R1mnfsYrFKSWMaZPFOQarJLqoW+2RYBAarVl/yxR3Noecpe+32oRI+63MfQvX
mb0wBg6ZXfz1dHAZa40nxEeamSQS3ek9F4kQw8Gywunde0W7Pk1v9txEuKYqghXUcaYUgKmkugos
zVXo+4Yfw7R9hQvgAISmGELx5jZMRyVzAlLivWrhu0y6ok7K4Dh3qCFgbNNdgOUMEcLbXY7oyuSt
6O7tCHa3F0GLXx7/t1EKdGU+7CEE1S7MdCPryE1P5y+jTYxh4+TMfZ0kC3krvKqZhBzF4BJlF92c
1Uno0QZ2al/EXHwVv7kLWehBsqg53q7Tl43bKvasArVQE7Ez6eciIieARqyuxADjGMrqIfQO/+rG
0NxUT3DycfR6moVEU3AM4QEC5/o+8l8nWXYniMsOIMuD+gTI4CRMGxlI3YF/evOdMKF6tMD/Qui9
oRsEp7nMwrgKkAnQrot/EcQK4Zneots0fMB2K5RE8/eeXBwiIJquVEvHFn76tOpBwjbSl+L7un55
D4/ce7FSojxKQqg+f9BWIC85tTypxWn0O4zWGYlyWTuLkTfEXCR1g9daWiTUojt+4PHrPRmjog9p
f0g41VZlLGH0KBgTzCuid0nQ5G7O6dfol+Zrrli923yc5AjWJtxAT26Vjh/Xex6dOaKHzp9gA+Xs
ntg40Zk+rjJ+4lQsHwMOAqb1EKixBlYXsgStOB2TjB5PnUzXHMZMGQmZbtpuf17vPQEF44NNyvix
cJA/NnbgOQtyhml4qck5FQXs9hpiCN+AEqAEEX0w31suTncpoECVg5J6COAbm8lpqqY+D/8yE4Rc
LpqB9c+jucJIoJXNU5wwpZ/R6x67bdsCut3C6gZI6MZ/cjO+r0l7jXwEQ/ea3BM/eyqJe5KgMFcx
XpLLR+/0vgxF7YlrYX+l48TZUqEtQVD4JnxKnfrPUkIgUTYzyTICJTL/3D8be6ecJpnniDUpYMvT
uOVDIbgZ3KFPO7tiN4biq2D/bM4/z1YJtGbnIc22q7/k0+pb8VPfXFmLczy/b8L1T9zBS/PA2MWl
oOeVDTvr8zREeiPeAaE9PBovwf2r2gABOZBWKbGULTvODpOpDiXIfJou4WI8p0icfUonNyYmNNNn
V1KjHZz4DZu5RPX376K7G+es5r7cIR8rBMkGoLzAUxm7GH2PD6Rjmqqc7Ce22TlErNdfVHIMtORE
nbV50x9LbO8Lz4MZx72JSpnu67fxFmlS8NbSF7t5llC6n2d12S1TRkha1egUZA3+UgF/dNx9fGnR
WzUAZlgYbpyjq7lKdya+wxfcnvFgM0iz04SaZiTRdKInCZIeFDzDbgiPvpKRT0O4SoaZA1yBsuoe
nWnuVKpbo2y0mA3DQXCKMuWhO8MEz/254JOqAQw+IpReNy3bkZf4ITPqaTO27cUqhZJ4JeI5tE/D
FRDM6eltkBO5iYi5J+J1eXrBvotVLR2pW+bCBfiabuMplD7wD4XbtBLZe0wr6IdtWWqQO+yJN9Xd
BRIh8SHL81sSkprMUmC9AEUs6Z2G6kE6MICzs4lOAe015K+l9dPxdKOx8RDNANDe6r/Kq8HJRQx7
RWBOcscyq+nQViQJrBNWdbp12P7D406YxROVR7v9amP55vS+QZso1uDImTZnYcv3DJv+LfGUEG9s
h2at2BC1rV29lRilzMLASgt+aXhEY7GEs7SB2qBWYWEGDKoSIyMgzp0mzEE5JQLFTlkNAkrDWKcf
JPY1qNykHug75vgJmNNrWlybGbFn+spyDrk/BIV5j416DbtI4Lsj6FKE7oUv2DtXpAhv8vboOo7X
SOu5UC9W2pxCzezDSj3K3m/cY/aVQ4/BMF4oziyYPPiYJ/OZAVbs0oj4UWHnHHfTkUfNe/mmWxS6
wU6GnnjK+4jce0auCVkzDw6xJL4TfQiXcrNFLkNFc5ijeM4mi266F8syPerIwlqDcf+RzDq7g5Oq
yfk3W3kqXR+oAK650M1cyJcDkzvrLWuW7A95TGavWo9VDzzRj8HyPjyq9eCZhxTwf8PVBoJUFHku
Vu74kc7k1NA3Sd8g9dAeUnHrPYlXkw1wzi3cuDXBayHiceIYaPqvJdm2PKFHv2zLt5Nwfop82pX2
YAcIzV1naGcyIBJalJaMzg5FeJ76b4ehzOM9uAHgeWc15lwy1lMsYQuHaS/3i/tB36wkfttIAaWp
yBcudFNVblcV+AP6NRTx5XrXBGnxQ28OdsU3mVOURIzsKNlQ5ZZTwUKzEPm4A/LTqXpqy/wS2HjP
rj03u70UjVZ3BoA9BCCbo0bEKpAXRUNHVftvzqTFOkZit8VGOIB/mZlT1R7aguRAoxZEsPbADQE2
jx5cqxcJChK0cxWKiic5CJtRd5tFTF2T/zdvPobH+saioBFLwE0gtW7WzJuxPLeUmSlpjBLX3c6m
9haAq2XZhNjxd+KPmoi0LJT1kTXE0Gpdegy57JDdFz1bp+1SjGtAV3yxm8N4z33ePuokhomqd/Te
7cyDEsOvqQfULVzj9HQjRDT1NEEsJOOhnH8FbcyxtpQsKN1evG9QoKczcTAs6cU2qjHtR+TO/M4B
b1O0q24otlSCcAXTn1RrLdrP8d47l5puJoB2xrKkjoMKCraLhPtJiF08P0yXv7wjk6ejnD8Gi+1s
dTjyQY7dfy2hdtuKNqtlsAj45nhYpMd4fMsUoXq2Iii+d0cKm2M9WlMYvLg6OQW4HHmwkARiLoBA
hAxMPvhqI0lIG3o0uKkOO95H5jiEvpZ4Evzmdv+L7pl3TsE5YjM7IzOIKT9cSovbwzO9YQGY7NQh
z2FhWxceXpcidUL4mntdlF4pNMVcNCpTxhMNT2hH7PhmQ5IJiCf/kIBbYJaPLvDgzAGu2KorVNQU
Yc3+li/KMmBpn7W2o0pIxI0Z6IfjcGfovGv6at9XK/41pEHqnXeF4kMgEKWGvATUYHUZwNp7A+0n
PdMpf//Pl8q5YJjgwTeGmoJXrrQgxZ/opY2YZq1RqHM+6R1AKYA1QEyHSeA5N63V+VRFXIS9pd2c
/iSs2etVUKd6ag6HhhjS9IZWiXE4MwuqAlxk9J5M8UDn4F952+5+93tyAF4BK526SJ68FGBRjOn3
CpWjPXqTz0GrwIDQI3rltFZWkfy745TtRjhztVEl3uuxRmHeFHsRJv9VopFcUrBHrIgfwlV/7gvG
ecaxf07E1nXRsfPG/iHJR1olRUDIUN0ZSO0prshWn7zYJb8slBtTu4Sz/15/OyIIBKRozEphK6f2
BL7wS+vmMHcbfUsckxNrYMWk8tAPnB8igZ2wEKGKPvpgw0l9xU+GLjKo/tm2U7pd3mIyyBvl2LGk
YZBwcy5EFQvQt1JdgmK0PfiZCKUnwTY8/67tMZDxJzkIqeN4t9EGx1mKJNaDL9dNuEKBx1WrBYmE
JpmKjWsRYB2b+qYlyAIbZJryVFIPlWQGrTg+eRzxIbMm5+gUIfJ7WUG9Yx2j4N0tDuTM0Do4udTc
WbR7x0/8YNIVyBrDeU8cNXJOXb+cvuZrEWFVHgVFqft/+V9Jzo66cg+zC4WbsYH+qb5P9TUwb9Zj
FGXZ8qip7920Nr+v7Jsi95uev0jAGyYW3yJWqtYl8v15OHER2e6Xjp3c2cc16dcHo+28fGcgasyF
dfXgTyi87GRztIQLDVxNWvbQ4CtAsj4jb5Ep0rkHRgmZqjY8B945vqlyNb/6UPoYO2TetERpFVaK
0QwADz/teTlHGpbff2J6kRv+PaDIiZ7NthXOq2c65VQsG5VeIZwgNbl7AoX+GTOGaXqvVh+F35kQ
fQB+CdqkaOU5pUy7Ky799X85hicsgtTvwrWN63xAxazHC8JT96yne1wb0Sh80i9IjaLst2xLlCk1
dcJ8XQpUoT+VNA2uo2utynkJxNqhTNjqfktg2muBuwDJRLWNQNRIe7Xf5x0fiP+VovDw5sy5R2hN
2hjiQkB1cqJGtlfhmRAYQDfKu6S4r/vu2IURvLE7N4kMe6aBk0+fGEQGzLc3kdTTC+IBzr3Pl8EJ
jHELIqF1v+p2N9vbPo1g+Cj0Cz6FCRTFzO5+swfkOO5iBns32GE9rAr3ZJk+Ns4/Zeqd/KyxfoiY
IVYBW7SQHO4gazdcHyv/y0Ua8zZcfUg07sXCv+0oIaaDLLj94424Z26QSZnUL/wav7hqPoznUhQM
+gUQLIvcIYxvMFYLwk1t5KCOELBKFF9i/BWo2jqqa2bVYEQw96Zj4dxgr0KpK7RjXbUvW6ft+bTz
p0lRy8zK5qDEcfhrm2pvLMPMtzgPYy6Cbp71W7zrCclLDspB9d/1GfjwDIof+eu8dNBVIu7DbfMG
8TawIfzHTE2LVI0WldFU50rTSpcS/3akRxTH8LhF/S2zkcB7mZZvwOH/PEKCOsI5r0NFkaUDdCwL
0YUDNK9I9+XrrJ6Ov/9v2ZElzjXWcgLohc2TN3pwtG9DsheiwBzSSo3OEXAsxG2RJSH9yRRjPVDZ
yvkW+5mLLto0v8iT6Z1VPsfTO2ZszZKxnQmp2vfaJMI5lqfIbJFHm0rSkn1slBNYCqTa9KURXDpX
DHSMY0S1Wm09HA18cnkGTlUA9gAXEm6TDS8ugz1TFC+tXEGvosDkcF9CfsnqnEXGeVb9vYPwG3pd
jv2IzMMUr0LaOhSbEUlctX8KPlRp24skg0p/fvjEJnQlAO98FgAAhowMsvhTTEZeBpqvJDh4oh4s
x6sMQgw77ZysxuNDlhKgCxn6IWq3leFv1JN/Z1u/UVFeoDIzgmk5euIpfStuny4qfrp+ZD3LUtLw
XVl5QcnLKPn1d1qByjcrcMSnEaiUzOBRmZ4Wgowpega7b7YvEFws9dFP9QM9befo1lkupLtBtRCg
nI/VMITYaca0CVfWmSTwHHk3NQT2IpaLoDn/xgtmrNy4fY6MGa7Xm1VW5adzQ4nEkuUQb7ysjfhr
mI06rue0RAuOsS27Z+1lXxxnWfLJPPf0Io0bOuJ5FN1o6xu87YGn5OBoefz5ndrFlqKo+LHNeJx+
IMWIZJoRuNavIL6nZOu+I8m41CNm8cURDH+Y92pK9CnuXUZ6KQAovNNVJl9QBe8z4n6Dsa8gTAnU
jdhpHDp58r0ISogu29CbTgj77v2LCsgyzc2iSy90/fDe91GN9vdXIomyTdxvHMIERM1Yv7WVBzax
FC9Kk8X878wTsjavKIBWv3q9ekOG61RNodcJY2prN6BSnhtC394+IA4Hinf+++ovVZxJyyZ+xfnp
NqEFgvBZY+1ZbEgQp4UKCFWnsDDjhdwPpUgnjRNl4sn7DtoreujqGKaW6tUfstE8jnEe2yqGi4+O
KHpFRof51IqqUu2wkVEdJ0FJtHhOdkVb6CMrL0nl67VbfR3gupbX9tyNLAD2EbI2SuBjjY+Po1uC
ylnU6vsRxp9cUbRY28A28CBXx0LVzEDQJ9MkzQew8A7qSlCcnrzX3X6gXOcUhP2riDMSLNqAizY+
Su5ce25OyEHey3SWY1gONCRV0nfQsJ/3QjysyvKhDdpCj5YcEuM1noKP408hKDttKN7045V8V/jS
BhH1AyC2L6PY5jCQ41BdCLvTmMtsRV0bhhBiLxStijy5XmHTwSKClZOlbS664S4zq1p6g+u/9qE4
lhrIht3MS4BpYfgXLO3ubZTGOPCWbETd8OgSGrjC1nXZnCXs7h+TA4t3/yVFpm8aFOON3C5SOBAK
g5muyb6433GmCW1RIo21sC5Rf53uRdTxVXqPcZwKQ8ZKquSAMxs0WneTaY3oD6onU6ruhJPPpFXK
otz5REPIWzBJtv0U7oi+bWG5mRfUVPl4JVJvJW84DNmSIfxyQnf5QgBJE2OFVg/8rtqwH7yZ22Vu
1lEAGRb2tf7lPTSbdDiXBISuS08fFV7+JDhQa/mQ+OYxCoMeX7Q34hQhVvPsYsivE26hZE6jZXnZ
zPRnKlnEZGdui1rh3etIoAfpRtAtcdTys0YUZa6GDaQ712sm5WXKfWkMvIGpFzIiGUABu6H9GmBK
/A5o+wzZXSgEAvjaGqJiKXEfFSpgyDIpPAgSyX2jCJeyiXErYfezBnK0NWe8MRWc3XvqPdJLySuL
zBbtK7dF5+0D7LXKn1P/J2o8yWI2dZaIKlJjK/clIX2rpNDBdRxoj1CRzfxtDvCyDiKAYwY9impt
LPeyaFSD59iFFtOM4i10aFUIFBLZIulYLXNoh9GorpGi0S8gsvGdWTeuieknP7utJRfzBVbAz0e5
h9wmd6KF79tP8uTbT5gxwfn75LX/cCdAZ4P4jAW+icekw24pu6GQ31BA4dBe8py/Yxk2OFxdicz/
YTVHAbcXs8BWb7XEB/PixmpdyARBl4TzY1bHVt1ONv4o2sWETegCQHhK53gIp5/f+Dv1fW64Vcmu
r02nmIJRwlOFvMMKfORB87Hvnfunhs3PYm8TuLk8M0UkqUDQKVTSvYp2X+NcS74nrZnouTNZfvG2
9HfKFigt6U8XzTMHm2xMDbrWZFXDHtXMutdR6T4FuISFWcmwOjeJ6ke0dcbdDwJCtcjlRU9HA08j
njVLx2Y69GI0uj5eb8oM7uShx7m+yHYBHM8x4tj4DKqah6kcj7FrLQ3cPUbpA4auQf6hFNyC3Q0O
BnCuQoh+84a39bpJvDz3fPSBOAX0s351Tl+qNC3Yeo8dtAy2lP3GLejc3lA1vwi8n5NjUPkSjofx
Df3fePGuAPizr8EXTqfhAkxt984h0kiESCW7Gbme3Ecvcoh2djlpxvEkttlhqRUngiqq9cibueJM
G8wq6yxRh66n6ZSNJvTQnyYRZH+s3I3YFS+jOC54Uqhhp4OJRP7tBMsT2N9Kg9w2siGlMr1WNuOO
ZnerP6jN1B1722NdYCoMRzN54kZ2RWRCYomAOkhgpQ7aKksXM45Mr+lbO+SC1yJkG3WuKGXt+pkm
7tEfEmPGtq7kLgk/bBpACs4A52aGu8GezvtP/NtfCZxE+VBe4ZDVZP9Fc+v4eJ8QbyORR0kYqEx5
vUGYenpFLRsuqupWv3JuV3YQgGfdU4uFZEumJQt2iIZJe44y2axoklCErEqiDYC6EiSq5uRpb6r1
PrBFrj3a/FtpxZzqoTbBzp8IAUxa2r0tB6920uBTsGZpImkS54nolO+iTqSf2gGLeMKQSFfxFFFP
B3pH+DmxzECc+hWHCuhee8F2aRKB38DCuXw0js+ifreu0h3DIBg/+G4gFvHW2SmB0RAhl1s/qbAW
lpPjzJYoeNJuEmoLw3FLqrjNaC5kOD9C8oRsbphkhon8kearm7SexW7oFSZ0tM9y/N6bcDEeEj7S
M6Qx9ZEN/lJqp58ZlChAIz+7I1FEdtyWzpG4l6+kFWM4UsxU+QhCSDcq6XVnPzBTgbmzgGHVmGjW
+OghjVit/0IuS1BUo7n4GKBc5vMbWp4472ehdAqSJY1f9K6oivpTmgHXgrxfa16QVXQixur4oex+
G7VcbLoi+5iteu8GG8lvAc2K15OiuA02mDrc2eMuwjC71bXa8ZY77gjSKAl/L6spucaxIjB0PT/a
QmV5L/hBZH0gNqoaqmFjoAoY66llch0IxU8w9clcmgJKbrNUqfcZ9a9p8SLVMT2AC/dS6+0H20aC
h2kzSzctKzNt2suxztGMKUJgk4LFVQuz2tuWvwOMYA9ZM6h8JLy8vhym/0wqp1FycDAHWEy14gZY
qDDOBu/ct/WC+EKMPOllkzEwOYXzep6reFzJlH+n9b9tBSd27MebgMCrC5MA5PFlWAZNDcjAcWJR
PktDHLRiyPYJxHoXHJkJHNINsqrrDju1ReEbstac5cRcxy54/Ou0KGuBydjufmwP4wzODGstsgok
6zpfuAOvlhu20RNuwhLm1oB7bbx1Kbi036Hm0ucJwGaPIYFwySgzuVPkQh1oS9qSlFZyNMYoNjCg
4m0VOD4/JUKXWrU3PzWYM4DUtHJRdh9A0q+KN8OQQFF6uZFUHm3xBTOuXwAYEaU+OrN4YtXug685
lqYFSbeXmKiV9gXvoBqZ0CsFQAqRLeTP6+DtA9ggPdkczU2khnpJoBfTHxmcIw4j/ENwmufhE7ko
shS4/Z+JcxmCHxpV1GLRls+Edq29zmFKIXAAQTyNLCdvxebSTpeOCD15V4RSLAji4vpEYvMVr/fn
zEze89mucKE2W3ByakEGz2av4zVQSqRORadlAXqPehozIQ6mvpO+Y6ifQ36iGu1oqiY124E+TQ7m
5273CbyNeuNN5LEQ1f0fxzJ5nfJxLkxgO/fHQXbTijqZDgZSnz+xyb73o08i+vSLk/tMBgYMj+q7
YfRjueXUHrtJg0V56JKcc09vxBmO7rXwgPaXVy8eSL95EwkXVgu1sWxd9Yd7NeqayZWQT3V0bwxN
AezDa8wWSeruC0dxsCr/FmN+NKLeRyYq1w+OYWzoS0pXkpRsnYWgvupm2YzYZTAqjuyXRCCuJVLX
dFYnCIM/C9v3UmAGGyNCIZQaifrZkuwIoOziCSrtuG0yVwft5an0W8KmGqAP0hGeg39sBvA31yzF
aEuudiF7jSLPZoSeq4wSO48i1EJEQuzJHCoqWCfg79QIIZq2MYYJesBJ2R62NZlC8ls0BSH9nqQy
0HmQS3oezBk/PF2VfF+XBc2BacbvXhJiJOiT3W6aL4UYoP6PwObec8Gz75g9D3smFJnOO16f9pfZ
ykxKf8YHBT1iVUFUije536vI7lCj4FCkgBu2/xlyRI8epJfPMWhdj8AxBAchM3QUUa2yVkTeCjXi
8IDwUiwbQD4Dhcs5FA8aszPWLTsw7b4jbyBXsoryQFkozk/MiDEckfaEohWzVnCD7Wgri60dca/4
0rqZ2+8dacz71QGCk0VYSdr2MK0sDCbTeZ2dvMQLuewMLu/tnLbI0u4B4Yy1PUwJPsUoQ/6rVZrp
mlSPNg/23vI/4dOTYl4VDKa9QKiRr+T8lWbprt+79tFG5uUbWVoL8WQsqlgUETzYj37S3BFK6xYA
ZdrEvK9ltFbU87sYFbtQzhgNRD6opOB6iscdAaFns9IVpyeTo+aLKdMielxt4MlvrqxHwuAoTEWk
KWQTYIZ4onMtwsrbNCHQOk0Wn56a6ywGY4jYbroBguLO8y0mzNGNg0VBDzsErTDBxFMkCsd2Xhrz
eejwOQlzqBVGVdBZ8bSnJMcAbM8RgRlUmq2kwjucoidxbdxk6Vtzb2mS/HB4HNZ5wiKPcDYquzxv
YNRVd0IilmtUVKXD597o9pjZlFJka6gxvXadEXoRP0q4R3bEMMg36vqjKBE0N3OCYN9UUmoDk6jU
yGHXyNXui/Xllp9TrT+kqcR8qsJA4U9AhGsuZNFRJnSUPTw3hKOk9epLTsLzM4Qlu2tqZUMtesfk
W/e04Cj+eIBcCzROZ03/7scOctXN4SJSKpDVVIBIKOmAclEzoSTJX/3npULxzd06zeWVQ/mjK1y8
kgPzEjUnlke7TYUlE6kLx/g61lB0z54Si5ZKj0wrwB4y5NK97sqC4eyYuFcgJPaiyFRIizBDor+e
ua/IY5KVKQ5cYqlzGn47CHr0lkutAlrzdKx/2f3Qbf0F/etQKTi6Nz7bChOD96z6RWvgQBeDCms1
4Ml/ymzee87JOF6WKylDdwTJcdBJ4MhsGMa+RsKu5darPhnoezNaQhWcfO1MhNo42GkW2azivc2c
+JdNV827XoJCTGNHhQe6o1av6v2IIMdLtr39e36Yi5qM53fbrZGRL/U3f/kWXAh8R8LeXQO87Urx
4MSApMmARWHMeTWR8QUxuL/dN8nt1K3WGnybdknUcbn1HI/cJQ8rsxRoe1Jop5WwqkIZsclhH1t2
dYXmtwTJc4tWpkFLwWvvNlkFFoYLeRnqjaUbQkp0/pLMkrJ0Lajl3lFm5tMVTbFmn6KpDa8i7gqL
Yxc2+Rl4R3wTVArw3EDP72ms1kZjxT4aHRhdTyG87Ccn6PeXm2p/qT3V/vnjyPkd67y9OEjwQHH6
OpxVfn/kLiJwa4ywngiELbDwCMcQB92axd8xPJDs2WsSHCjSn0meBJOSOY/hqZ/YcrLEDWM9Rby1
cSPOkceXobUGzHFrMxe4CaJJNYh3zAkpc7+0EB3WjiruTt9FQbkn5/Id5y3EhOIZR3lUtCC3EgVj
hKjkzzqY91j5HD5hx87oKK7BX6Qaix3WRGWRMUkw3WIoE7ws9xSK8rnFWtbMiStBruttlk1Mrg5K
EO6oNqDdHxbmkgN9fC1OxXFr650BgoOqzP6C1iHB0NMC87InaOV9gPaCC1ihX7rGzMY2DEKRJ7j0
/ZHa30YVDqm61v8GKJXxdl7PezYFmIGCSOakxlUlADcrtmA1i5L8RydeAQiWdYzC8gtA6nimZw+/
5C0S5Qeoh6xIX44/Smce62IkOxgAEAfHkZBf29hQw/2sJLvtY0uy4FMnXOUzDx3t85YVng11MK9m
dSP2wQnz8M84lVtIExzEcVq+bnNBKBGAkVRolm/CEGY+bicDLQltGh6TJe55/DyZ2ms7oHQRojSc
1UtNuqyz7b7Vq+ja3A+jVRYIsgYpzbKXgjL1Sb3NJHyQqAv5Uoxvs/jasYBWKGjRMhj3rBJGDf5o
rCUekgb7tZnLVIjEt1O2DuqkEVcee/rV3d8UgaedtKJatVPQoRvWrOfSz/awBJgNWYH5u92BR2Sm
ocQQRh5aD2eGsdiLDvdUI4UzV71Ir3KY+Lu/s4RRPUupjAavf1EPdcoZKW4mNLve3OHyC0jHTm7j
n1P0YKVxiz6XGiHwtlvdwj79x12SCdoQFXAEITUqhReUHpF5YcM6L5d4Wz7St9l43ICDiIC+LOXd
S8WgOVBiY4sbeI8nIOfQRZJZ6iMF/qHHyQ2JyY+Vd3dONf+zEaYPcKh/x+BkP501yNyd6VYHA2kN
cck/O46g4h8VbPqrGXIgOI2bwK8ETYeBhj6CMeViFhZtwBrIvW3Ypg9E/sB1v7pp1kr6OEK6P8Za
8sgHcE2r16rKcowFMDDkcdxs3g82hF+mUdHPJJovwtOaAK+bfb/zqRAPhErEHWVgV5fi0SPgQ5Sd
AFRiakWp83bmk/UFY+cVcYI7oe6oqMhlIPHq4gPdVWxo8i4CEkP8NH8agTlvyeqJ2wbZdvXhqZ2b
U3wK7bo4wCx29jH9awccL6BkB3oirOqOEmV69SuTyHrJObRMFmiL2lwHlIn0Xh0q/Do0R1HOy1V/
+5YpomzT9Sktuny/+oBOgmc21yByrPtsnAehuw5b4GdK06YMERcRyRY3C2WQEaB9Dl97+V4LuCFF
uHphfBQo3U01JuNt/7ooR/+DOizkRfGEw5jkmsStaX0pshNWROqKLzvUfUwV+pE/gq1rT9PP3lmO
XolvbaRZsxXZduz0Q10OsVE7PQvEE9Zwc+LHEWXqx2e1lCdY1uhKQXqgC4MYDjlt8Qw6bCLb4hcr
TskuhgOc+jvuDO5AOEFDx4WGKYRWmMIqLAuQIOXOgtVT/tj5kDktlgMSTfo+Tt1rs6f8flspT4xE
TRM7Z97+WtFJNtgDosKaLE+Bci168+jZ53lNv8Bhy615GS28yRu71sANcSnVlbnjAzzPBPOVYAMQ
XWlZC7wwwH8TRCnEsHfGXbEbo9OpXPTXkDq4UijX288B52NxBiQYQPSH7+dQc4CFYzWJvGowcYsD
VZ5zESft+bvno0ROAYOyQA19DV0aeYsZYHRZVdKUsISai88FrwygkTt4Hp7wEoPen5AAGh0OsYvV
Eg3VoZd0l/6nO0A/zM2zF+6uwhfhZ1al053v889Kh2CKTaY+s7sSRSKen0c4Uh0KfKC/ka83ATIQ
ljOsLAOx6nHNuCclH2I5pdSSJZjLBpdwryRmut4KkMDYnQwvUEIa5y8O2fgn9gIAfesUV0z31nnc
eHERbYBtYrtPZrYfg7mEws5ZIZ5kZB1A3PB2NP07SL9LXNXsjAFkOsmcfyCcq2jbkBIoxRqaQGz0
fj0C8PwTZw0uh2H7T5ccWItcQZY2F8nn3qZvHsbnWCIlLvu26019qPh3vQxFRkoKccnoWRJvpxSj
iOOC99ZoUgB+FPNK4UfMWxU8e4vOboVkPEVooYyfP9KWJnLnmdzsSw+ikGPj/b1nsG7HQU3s8gf1
xLr0ux885BUzwBsTyoyyoCZK1Kxp/bEWxtpBGURohL0ICL/qdgvrktEhnMcCjYDYLc5uLMleCWTO
hbuX25wBhmbR1kEQjt+0rk9v2oJEEpoUsp3e4V1o/yONkhQd4+p6DbasHus++Y8ERgVuvEOpMcAR
WM3C9iIUkHbOlp5Tuuqgd4CRraaqx3sRH3D7RA0OVygyUcOnRe5cJhBMb7zAYApd7FYy1DmHtD5d
yLOJm3Md16OcXVioFWHXw4vsxy12c+BIP+Aa471QJrShhrE0Yli9XhEwDjknAuEp8ObxxoE/Y0PJ
xz+mYMg5rVy4cXnLRe0o5eTLvH341G6dLfdKE1g2rAoXpPV9kQ/9Eebn5Cq9xCkkCdIU1GNjgtjt
KTOHcBDaEyQwaxhZMzCrU+BlsTOm+lQuZ90cAXX9HpUU0OWZIKfRVQ7AuiYSdtZ557mrOTqhnbrN
ScSzsnEpJNoQY8JQvSy+2cbExA9iyGVd12sJkpFw/Fc67a7M8C8po/eHX6dEcGSNfz+r2NsEOopF
qw2MxUfMO2/kXqMR5Cv0ClaZh+MgEcnc2mh2ipiQsH2+ucNlCuIURwNGZdSBKzcKd2+Sog5AR3ek
YIsedUQLgChUvudZ8dfQ4g5U5LiXnJBe22VS8BOowof1soZ7MrhaeLvfEx/P6Og4uau125wUZZ+T
QUFQARk3OgrMiSG+JbaArOY9+Y+wbSVbgSKPEC5DzfDFlIJ1q1y0DglQ5I6GxET+9gvFWbs7dGMp
P1jfRNV3S2mpZ1ACYg8cnwCUdMx0XqJYr/7QKZIlHmn1xP6R9Zagx7/wHmjAPe4O5xruHBwteemc
OLxKkiy5siCTTmDYAFmqAfua36imB/wLDctJzbmhtY+HuVRz+iTzsyBhE3JFV6UAxLgXZ/7RFtiy
aBXi97bNF6ZfvR6TzdyhuT1APBXxChTsVMIzkcAAJbJhxCYGV+zEJMqnRS2mDXd5vbu+FN4RAtxc
TY2XsKNriDVeMOgEVxR/xxSEMOO4ejpr/7vRc0w/qGA3IWKNL272q9AEB6Qmd0GDUxNikBQk8VLh
1/kGJ6MFQ+GwM+bmGMUfs6h+VZdfi0XvhKfcpUm/cnJy/rfx9TGhOVZI7Pe+3sD+yee4/7kWkZQa
Pl8ioK8TX91nZ/45gs7CmUc0CWXYUJTPF+dFi2UiL4dbGMWFf32TIqSjuxZykA+mkgJvpnggerbT
sjBurmBmVJ6UyRyj66TiIH+pVLUNcauH8QHNw1BF3UD/4ItCc+DbVWQMVHHp0MHeWiJmipBLel0y
HZDqOhs7sOiEkpRDs7bhAERB+7uX7jl5oEkcb11Z/Tfvo1ljnaXJbtWyYJR8VTlaWd+YWuYNlv/1
zy9q2vlJpv5UquvG4NtpUTzQAGX4pfXQU+/zfkOcOVcA+8WxfhHitvOa6SCckVGaUSBks+BRc+j1
5m52nnUuZB5BmhMMgTuhtkyeSV5B1iojAY8sA+28kSULPOOojweSzrmU6lW06QXFr3jl6ucFZRzy
BBz9ZDyeQ8aTp9I/6BbTriDNa8oqdAn1VX/udvB/zoPG3wI6HioDdk/ibLflPZ4yxLeWQXhCDv6x
klxVAR46Ajk1bMHatUZ0taEtmxlD6piKmPXHGBUFDV/XUAKuzbA9GoUA4MBQtpeEGFwsa6xR+/Hv
0PWr1bIFrF7cQ8uLHr3246o3rPsJ0TKoNl1nx6Y5LtfvZmfpxWeqMLkCNn5SwQzsZO5T49LzOPGw
DvcCg0MD+hh638rk0p5aHjugdoyv8HeBsOu9T9dDfYxFj3iZJSWoxCpq8UMg9ZYwEHghN2hzs3vd
h4ex01YaDoPEyS/6ADam2cSZDAz4PisNARtfuvYyIuBYmOxagJAzfMhKk6dFYAdD+9DFVGVaYxWe
niw/MkV3EwCygmrMwbo4CvJnTbrH1D1/hxhEs1WPPPMvdyjZRLGyrwxeMVkl9h3gOBoaGhziffXF
XJcQ9Oz6+K2BbMj6EfyG82VlV2Qv/luW/O1Wd6S3HEpub7N2QDtO41qItQkZHKrvf+cRSAnE132R
jUCDujyW7Lk17YzFhC8lSnzC71ev+Y2i7dugzfNN0vucym5fpUXWYV7tfgj6rvQVz3dnaxM0xdpt
3QiReFqefnOtLMGeZipTVkDe9xOwYZIEAShvq0CGZw5rQDn1dkz+jHZ0IZeXIw4S3cxkubn50iP+
b3GMl7qKh+73N0IiXAApJ/rgkG2qNOCCQhF0YZklyZpd7WjsQpf3kdOo1h8DfoMLUTyLGNqKn5Oz
9urrfLCaAdJOTjDMEUsGTABV5kusulkcSy+9zo36wbFV0q7/85gwpCLaZvxyGBu4tYRHZ5mYJ8zH
2EpvAu8LWDmiLj/CsUQkI8FfO7fsGa/pRssBUaFehBJkPxodlXvxAFUZaOoBgBnvv8j5skAQ3aOS
CrXKFlrY6KVv0gyJBNFt3jGNQ8OlKCtz4e5z7aCNLfHfl5J6yQ+r5N9TnCCPyaF73sP25C7/SUkB
As8BzzBoh6UMlzQZxLZEDcTliaqOwwtmelYnK96awYwodB9XZpYcO5tZ8GkQ9Ei8Vz353apS5+e3
BGbxddL5mC1CUwX1McPwfYrxM6GVo2P6m0jAVVf3G63TPBI8gvlSYJy2c5C6vF6W2on+PmN5dCRq
cprxCU5vMUWEp7hVjk88mfrYATRKVeJaxE74rNWzxlPXS2lY+p+FBeRdTe4rtM2JDWJ0PAYDv+kC
9NrGhbBgq/KxrRa8kzB/Y6G2suQSxUIAtJzjA6xhx2iJ3XaD9+XlXCDIWmEpMx6coNeV4nGq5WO8
tQZLoPJQmbCDq51+jvd7ewdZTGZzSo3XxF+d2dFL9h6IHCSfn5V8B/84Uys2IR3a3pZCSJ6A4hbg
Bdu2JazyK9c1C+8JeHD+WU0KnEQJPjoCmnQQfMzwakHj2NOjq6SJTnkUUdKWFi8rfyEUfNlNabnG
HO12SRRYAUB8exRWhoPeaQSrgpfj/DDOrxXGVoUcuvcPqD5CQHH2O2ghHExpGH09CGZ+S55TwCPV
kl1bCwNper24PCCG+GNdxvUMdA29YwYtdeGciJqQqdLBdKxXJIuDntknJJGQkLAgPYBvZZEcCyuk
tlAgxEh0PVgfX19DTxQ6vV/qps4lpe69dcFxjJV8p2krJ9LlDT4XxT9SGbsZDEGLJSGxk/vX8J4I
7trQ5AlVyu8MhF45ajYhRqdaZNkVQNfx/JbL/O/aFJEk3wGMJuKn0Sp6veLLQaG1b/zYfltpxIJ1
iE462tI8sMow3KUUGzN1yIkeiau8PnoL3fe9wCzVybP/Ld/0OkC/zkthuUBmocOJeRjXWwwcI56h
qKzJfNbYf5H2r+t9tzkwn4CFTV+o4gKM0F4cQfpzLxVyqC5CwCH9iF+UPTYnoCUatg5ba9loMDAH
nMMVLE7Qy+JKaLnWMcPXKE5yTNy7aU3ZSZeaNGCV6fGF9fPffi2oD99om5eKERTlWNoZLg2xN5zx
xC5y0CuBJIzn5yURTz1B3ZWDYwjJdJiUWm7PN28399mw8W/tWALtX5sY8h1+7WAUmfDuIIphz+DA
XC4MhtPm+9Who+/J1HXd1A+P89XdcsDJcax2VCLbEicE4sTHG6X0zocke1HQrl2b2dTF/avHr3fJ
hXo9PBkoHWW2YB+JYktJP/wJz9pTwb5bHBlmzrdDOC8LtV7mvOeo9a8DpUkkzl+KJrSK4iMUmahp
CFoWm7hv2vFTUgE9JOoqynU4l3l83WNoCUH/kMJM7G6MvJAws/yoShyuAkHl9Bm9vViRiEKKRA6o
hIYFrN0t+7nVUEfxLqGpR+Yop3goWI0IOgRuhQrv24+hU6Mg4SHdb+d32HTXOh3ZJRwIOl9wK6Gm
YDlK/yGvmu22VHEToC8HKjczxCBfazXim9L2gZ60S9qCeHyIi/RK3vCxqfSRKUWXVyNMdBisStiQ
5ij0TeBFd3/V92B3AyzEAdMNnq8nVoe9jjfGgdenM/TKRv/ippD13l9kup4Zh0foL2mNYQqAKHbM
cAfF7y7GTZbcCk2bTDjrfM7d1w3tgvFBCMPBsQO7DmVB8Bmc9grUGIKf9OVelVwb/vyezOIfRmQN
3i621Govqy+0VOgzB99TjyqDUVCj9DjIqNL4aevJyiD/6+ocmePiDxr45q1dvADLlQmShf/ZSRTp
0PD8/N69bLnRqQaVxmQ2eZ4XKZFRD+qxWJ+pEHA6c/Bwx8MiRd7gSdm+ma4hpgt1pLYeEgwR7qzq
pdXh89aPMA4UeOCCdXCEqQMOsoGUnQcV2K0GfT7obSRJweYn6aWz1G31NMqMDzUddStGG/GCWczk
kH/xV5n21Z04lT8pq9huz+i+8HhPtRh4I2pIUCgyf3gysUhNYKSNgp5yb2GX357qEC1VrG9RiiOR
Tl6ceZziB6wwx9W+BptIa9BE9YtihDFd3QzNyO6kYbRWGdUq0k2RB/vCk7htkf/gnNffPaHbPqiA
N8ZCRHa6wXhZ0sa3/m4NlnhArErrItxQl9RUY4u3I3nvGkegRTtr908toKtWDVGvMlse2CwGA5Uj
Im5bvlayr8riHQCwBWGH2NsINsOFbxZwPk43DrXbfkG1VqoK9LV2oyss1MfGH0HVYiNHe1rgBg0j
kqD7Wc0saABSF75tG+1SVGMLMGpe3aiSy0myHnZYYA4WqcWgkwberSL+iNkAkoUUWxpntcb1ARe2
zVXbUS5FJCo47LgaNOpStbrWXOa76PTgtGR/bwYhNIivayBs/w5I2aRDFvhe98tamHqOUUaMVH9T
0pm3dPEnqzro0UbJlihVVyA694XUgt9qSVe8rEdj3l9j7vohvWgCYlmfvbE9zMPE+3OY6Old5vWt
LnBKEX1MoPv5vc6h2lC3cifGuWLjVTvJ2/3PKYE/clJBGDeVupQR5+V6+ITtRe5QcQHLyqjSfAFp
us7Tnjswc/NFyS3DnOx7z44x2tAChd1WM+safEfFYEJKoDg3WMDHWSbxeIsZcKiBDpcmq8KqC35/
bGcXIS8A7EV+8hC7cvorvi8OVbKlAduNn9Nr0NOmSpUsGcblZuoHXsZ9nr84BV2vNwgMIwaqJ1Fr
DBDfNBmZpCI8kYwy1jjcp0sLRFYD/ndN6olALh3SBVgHFqpNbY3/a42RU6706j5IdLp69VlZOJsk
WwYDo6FQVr/QQxVFUYuuu68ZODvWFDAUX2SgcjCVIffnwHnV1kfBHRjBe89oXqDK4y4PZ/fTgrGG
/h5N1s8IUjwaynefwPmq/OrhDSvsbbIhVlwaov21evte70iswRKkFHF3UTawefIFwk3BMuXfv/I6
4tqoaWSeefgQcPUGBBq0HAvhSXjWoHC+oz1wL9DdCkvZ07kaZbEuEjfInyHuifG4ViIxukUUciTY
qPM4FT5SHLX41kKWvvxaT2qYNdy3Py+LuaS3BTS4KjWwG5xl4ppN+QjwL2OiKLqO2dc0dMMccypK
uTl6U3d9ZLuvPc0bfxepLtXBEXe91Sql/SXB1MJDdRJtNZdKBV7dMENh7q1rihO+Z7/Cm0+r7UlE
PQNNOya61Dw9fc6fwX5e+UwKsZ6zQL/A/jmMjbz/7F7gk1ki/ZLwt2VVCLiWqvVXi+KJDsK2trkw
GoPStltRwg1MwqG+7rCg3OJ1IUuAb7TStdxHS5qnZFBa53Fx+kDlXptknzw0C1lGlk0BfpPogv/g
0WWsizq3WoRK0R8sloAv8x5LLmZ9pGVX57r5EgqkwbZmqaorcrTOpyJZn6YTUjOVB30K5vLLO2aF
plX4XeRcNjFG/pMl4dDy1vV7wuwKI9xmImcq6ue5qvK2iy5wHGC2nJ1poGJmznlvG+c4PMZ4KKQz
B2fwJM3cm+1wb9L1YPVCkl17Q7C/3YuENr3+VJVoZ3HYPRlTbPX8LRF1HaNZtd+LGd9lrgHDjJm2
4NOE/66/O/lKEOMx0YW3nxR3NoFBQVAgx39MmuB0KCR2T/bKh/8zqfDzQpE2w8vYv02F5/LNNDR4
2TIDxt2ig/Y3EYqH2UZwP9SACWz1o1juLpH5xmseyqM6Kvf+xceOUQd+LfQsSlj+taIdmvRLUw+V
d5ZUi9ize7blSi2bVcuXpTUPBhv2RkQxiE1EVVec9LvVVWaAy8KTmMW+BscbpETfwZqjqbC3uRuh
BecWM7C93ls5/fURKQnpzRqrZWkKY2LE0fEd5UEZcFKrr73GLctjIfoqZnopU0TYvQ2OuByL7CGu
nHS0kCOnxQYfK/pyZfW7RGEKJwVMaMFfqSUXUjp+Rc9Ufiz/DFK9rnrVqHSkG4MRCvpOJ0TONlmK
rUgC3IAR1M2neu4M3g+yOxXCMzXCMsRUA9hZnmp0c9lIo8YBRZJI/e0Majv7gDeanBA3zjgbYaIC
OLgwgV2X92Pyl+3PphE0XjPFg9seJQ162gccbhLH9U2pEiSMjGZzYGXabASO0gYMtV/EHynCijub
YYis82VbIrogmV5slQfEFur1AEtCT4E7LdvfWwM5WjnGhi0vfDLmdJKSAcJcOiyQeujTS4qQHGNX
fjSdQGkYisbJHVHGFEuKVBPkyjhrKZuV8UlqCmMeDEuRScikElTVY6KZBms8aI1X0/3zNuwo5Mdd
t0lrUKJK1IbpV7cEcE6AaQXFs57kvHc5B70JEyLoBsC6bKXXOnap1MZ8p5Oe4ucthvcQ21cDQAS+
3Ic5vPumZgw1IO/halF4O+rOT89IFpJ/j46iQfyddKXCA+f8Od0hYjEtjx8++/GY4GsoL1gxxcfg
S0RIJJF7UxlGeQDMJkOBWRLFEMcj0WK+Y//9Us7j4OaCP4dUVwirZj8ezReg0prts1vuhb9eAN6i
zSL07U/6vZTKch2ZL9Yva/kc1KKoWUp4S1yBNvH1AadRDfiF2Q3sH40zTFr0MIOPeLfY2HhVPbBs
Vpi1jYge0vaCSJTWHolTUSYcy9JDTb+zlJvviWdPuy01eASuMtiwAojLXVFe33UgMeMBmWDE0LXD
7JuLAO/T6fuRJhvWRe5xjIIh2FaesJq+F2dqAIyC/Cg1HLFe5vtLGh6T1Z3v+vQguSpasMJLtdV3
52uO5UbPDXBBTscHJlEA6N/AQKFX+llfqi9gtg/TurVFdljMi9VaI/FDRTn5sBmFR+8E0wvwwAhH
9PmhqMtIui1W0J3y7vTBkfi0S1lyQzeD6lcz/nlfh66B7OIPSYsKeIH9WhpYZmxEKO3D4myOmivY
V3pR4RqoYnOhCTk9rIfeKcLuOxya3T6O+ecvJLb6BUFSG1l20pxuXgIQcWAk32BN+XgxMcTEGnkk
C2rmv9ejISwU+8KvTBeLaF1kDwvfQh4MS0jgi180igziV+QFrTrLZGlX8IXPTRL6cQqKNsJZ3TaL
2ANUQ6eSK0lTJC25YPehs6TdWEB0HPMmirMjTGyI7kqNO6YiXq7VB4Kals7DYTnJxLBWQSq3j9kp
vWFOyd+jUc7x5vD+NNKRfdav2C/zKtay+/IfOmsQJyg8Kd4662FpRpi1AdSptlNzdHZG5RhO/b0J
t6qz6u0gfWmGH951y50rl16knldgSvS9y+oweIueL7v699vgf3t/JLPVvMyFJ58DymElpP7xFVn6
HENSHX7zBtMnczeTnm654/39VtYJXDUK3MmesAAzIkB5x/Pcu+OEu2iwHzi79T+IwtpqYt2Auw8/
2AyKp7+YDFB3dPhG45zfDnnc+PeOxLxhwvr1HWzjdx8lx8xFonjICXj1elvgyUum3W3grmKw5f0P
eAcVF/105K45QBl+Kunb/SNhjJrYr54g43ImDG6KBtexULuiKfzJeLltEnFGVN8nYrd1f2L305u/
86vtm721zlW4XW+0bLjQ6SxclE8dcJtUbkg6SCEbEcotQkKrjiZt9sUzp49xPZMl8irU/xAiQCU+
8prflT8fToYAskIXtDjceTEZpX8vAbEk7TmNwgMIMyAkceHRCTtCZ6nKe65rEGPPB9Zi1a3wtncf
QQJIV99eYIy+swyrRwUu05Y82Z4Axni/MYeyYoZRWbNddJsDCV/6LYrYH+YbCTDgM4TrpET6Debn
D1PevkSMhzJ73kohfucPil3Hqa7oAxqg8iL2Oc4wFxcbmNCS8+b1RtNCS9r+F0JhK8VBc3OzX3XB
zSGZ0vdGX/KgKfug++G0QVtICZuR2nqL6TuTjiUXirxh/td5QYffYycfZZ9/1Kq3C6wY6fEHnV3V
qC4ISS5MxC+QxKKGMPX54F7eNuAslGs0sKdu95O5b3vSBuNp41wPfmLLhL6JuLLsVx8pdm1YKez/
zlLecYxTAK1XituGJ9c8/Ndm8S/D2Vq4hKtzZ0MYOWIa4nvGKHysO+d7MyWsNolvk9M1AchSrBZe
PVcTjqybw2SPsH3G67vFLzn59WVjIe7oj0ENAVVNE8+03/kVN/8SZOi95TGm89vi+yV07k1Ci+MH
SJBhTLRHi3VMPxP3cDQ5kGKtfoxsZ7a4zEMBzDfeVNyRyCqmWLAumNqtXievkYqw3+e2uBM6OkDi
Q6q3/Ddyu31KpTKtnPJcN40HvjNb9O8ERP0Zc0BM7ofKaIpnTXWPg+pPMgh66lGeTCV/BtOJDMW7
gDQ8+g/cs+vP3Yhi1sPOcIVqfGzVZW3U/yX9qOYelX5pVKppy7ax/QTQkMioFS0/w92hTK0OdJ7B
lGj3oQZ3mDkcrw7H1ddVH5TdvKnYoJVV0Tt+C4S8T1SETxPyjDvTiEvpgFiMMhCHPOMOTyePvJc4
/mioe4aJ92UcJ6W3fmWVD/YNIgOzP4Qc3z4MY6eZ1MXJTPcf0L7SI1dR6dk+dVXblkdnTC7+y5sC
R90HNMs4F2wTqNx8q2Kpcjx2Nkxy9bCwW/BMmqQgTwQt4ykVh8I/7kIKvUPcAv7HJ7n7h0GU/G1s
Lfc48zaShBlVQbW2EGPsldRn7+pc+MCATymOQiU11Ge33VGWFBRDGeSY50DGEbXRRL0xnaWIadb+
kL6c7PIr/7h8Rne0iyo7Vx9TYjQ5tnMYfPb7uAGyj/Tt7o0/gEaJqAEvOW+5ITaJRFnQC2rKMO2S
/T75ktZysI8ihaDGVlV5RGJx3M6YtPNmEFKoLJ0t7eFZJUqzEYv3inejuGmeuh0iNMTJthyvSyxh
CfgXVkIxcauOKFI7opYp6M1E7lH7Wfdgpb4AsDBZvhvaK/uMVvPs+F0z2+v3u+gp0FKfJ68ivKBg
ocHG13pG3BLrSXjoq2d3grE9HYHG8Q3Ar3eMgwk5JvlPDbhwoNvR1yKrH6k+DmDslWlw6LTFC7eS
LgUchjIiXILMrht+IBfFmN7jL9s/doPfxlIdypripvJ7064B1gmkGxopiI0/5378zigYbMKDALo2
iIV9hlpQe4cEY4IHSSS3geGY66JeUXXNgu2iZtgeFB6b/R0qdW/nLURA5yapfnaAe3RBetqEY2wV
f7WkIFuJJZCwdGNdaWqBGPjS+C6mmk5uO/Klt9HvkiSf8ySrVzNEmeyGc3vANDV3zZ81CBShGOf5
3MY++gCldLu8gDcMkkj1GJHD+VX1GtvZvjPSIpp+zd0pu9M075rjDJEXA+VXBVmqH0hMvRM+RRYc
PMxT0wzSZMrR4tYiS79mwj1tp5SBLYbmGyR72rJ/JhflybZX96VMaIh3umKbfN0QVr0NiZQh46kQ
uNVfZp4LeZElHcjImT9YV3bjgTeH/i/fkx3a7L90JXEwxGd2H4BEhNc+431u/VJVmniV7IRu/+Ap
KRBhhG8W8pAchqyr5XGGltfgwl1MRbGtwF9gPQgr9oaPIYv0Ga61x6ZoCZlzgxzU+wMpUJmSBg9P
OvkDbT00KZvH5o0tDe9goeegkzGmzooyMQGejM4d5ng24JMF1RV0pVyyKyM7y6inh2kj3Nf5+ja2
KZX+S5Cgs43ia0OxOGoNJkL/YCDk4YyG/fSbSrZPSFxu0rNku1QqTddmWZVxpcTxJJP5PGcxklv8
OjJ38acIYhB1UKvSMmy3gBNNUsBs/McCDSaEsiTQ2PC9sxD6gTVgGVk5JiZHhtmK/iMYoF+1z/KL
h7tHENm+5wh6Z4owxbZ6YoptTvTlF4x2d2HDEbxzNm0hyif6MZ8NJ1EUySNUzmoS6LcPbA6vyxJj
zf+5VOcHa1iVNzhLYXnCeA5eTxW4aRBp20noA7khn1ud+x1eUWXVGw84QzaSdxGj21YCPCnzMaYv
b3VoHl/HAHu/xUOlXZEFnH8gaMM2dzsBN46njxO5frcBo30r/m8R/y68SqxDnseZOVIkIWKPRnSq
UoE3xEJBKj9tuRVUNpf8HAGZpuhfcZTJOGgyLOZCVyjA0cLaGbpLSeol2n5t+ksqDWVEi2Jnj9WR
znsJ3CXkjel+QHn8AX0DH59z9ogZegQVuQ5idCKhm7EAUpJWdc0ZlvW0SapzTAcmRIh4Mgra1Edh
omCIqaVmlLO5i+i5fGVujYz0MBryoUaWoXOtM/SI7sW/APDthsgo8/NfdWUc2Hpuc+SoRbRc4ECe
q6VpgsJisSmTEKu4qXF5SOolrCArkTqcZeQtep7TCScghidS12fk0ObdDUxgHrzxNUCzgBF3Gsio
Omm8Oe2YhwPLBIcV3NdYs9dfeNBXTFgpr9jU09ieynJ/s23iM4lnTP1AaL6J0mk8zijn/njS7thF
pUQFVjD1ot/RQDqpOnzsa9trZp44rHbYpEw0mUp0GNkKp26mtGN0TPhZXD+45reKjBAhsbPH5aZv
+mlqmZOlQ8rfB/3XC/m6qMydxv6xZhGwyIWUdPlMGaONeCPSJ+X6x4uVFpIP5IWiHMdpi1uqhjLa
BLMFVnqKtfyIomnTckAyNfFpNLWBPUfeQjs7DC68m6ldbO2OcEob5vg1d5nnyEQIbAOWeYWMh6qi
PYkzacC/xYKWj5TwZ+Kse/cXKOEXCFg6U9v5idXDzKnGJC09He+kD6S1MJWLWmKSb9iyZYncJM4f
FekCnLRjFQCaFMz/AI1IkaxSz3Q1G9vvtC6o0GkF4dgn6t+sgjMs7zAyNXOx0qjCqxrNl8/AtRf7
nz8Y5FmGcDZQACUfombzUi3ttt9yHG9FrVvvSiKJGqdp86E3SQiD+pAMMctZsEWIb9282tIr2Z51
bZNJ36FGmSZ22NNr5GkYO0/glEUvpCT4nHLUJvt/A+NFT+Z3wSqDdqNOEYr7DsnYyLxvTdOPh7tg
a0nDyX1te5OqU8Z/oNH46ygeiOHhCvKmgiy9o6FAOb0+xKVVYnBhxyp8hI5P1oHh2Bf0QvwVmQKV
frKnU8TICHDZ/ZaURcIgUNP8H+KXDu/T++V4sWG00gh3QJvZ2FohJiXr9XGqIZ3Loa7k+C31XMTM
p3ELLvvkkz8DfVLQixP7HZYyq/93m3n6C47LFjbctfCvLTIVgRJYwjHTQyuotFSlMMVZ7t3WjXED
C3LyoojZ2Mm0qXNK9QZ+d3PdF5y+LVE+NWhSna1gjyZKcErZrp5CFol0R+KBvskv5j7zfB6kSwpI
eA1BFkV/0++jRHq28db3kNO0yXdDN4BGtXvRrIlXvBO+Tw0kh7HU3lX5yj4zzYjqPv+qAAIMkRga
wmArdtMWcQlKpeSOJhHY7e6YFGhvEkXPkOYICA/BAzLHYDOyBtPZO6Y2hAcwbQ1yZQR0a9xNctpK
5/5sLOrmJKnMrB3XydxHwByqRJ5xsLXWhCCEORKrvvbblLXkIY3A7y6CHffQvgwwcHouX1o3hiVf
1r4NllAE7v7v3YWEWXAwpDKytWgvynrigsxP7+pm2HAFqWFhyma/U73uBR6KUcV818Mo0tWno+ch
+3JgsV+gQPf5QN6YPDYplQAi28EMcnimdcvlyuoeoi4fFyGi/8EKAacpRn9an2+63w4ee/q2UWe4
pcwtGmNDyuymLElmNTO6Ml8V3MKwbh7noXPtuGH8wD42Jmtpw8wuM0I4qlKyCJPSbb/WKqF9ivKv
9eRrN9IIPF+mjv8hDmE/p+7x2tvSwIL5VPmHPqSpehNWsIQQjtuRhBh8dLE1yjFJg7CY/0vyydvc
6ej3K//bLAPXV55PZTuB8ClCMNDVNDQfaUAG2OdULHoH3d036u0fHpuV+EEGY+AnaYMGWFrm6PzC
nHTGWlfcbsSVEqPEUiiJHXT1uEnRIaUsM6Uc9/DGayGwp1LSdK2Rrfa2T+xlefoRMs22MRCSgsoy
Y7AL32M5NVEyqlARWRtTdfgAnpcBGRTz6RUXXvoCT0cslZf6TyqoC0FZwHD1KsZJ/YRoy8jfPhob
JWNbanMbqqHfYKVmmwXlM+wYfEOV3B4e/WPh9aLI56rwmFrpyvov8RRLOe+B9NXaRPJn19udl+pX
7q0wZHH0OXHAXhUau4B5uGghV2kshuj2ycqlSLsMx/0Qpej42SblhLqe8C52qOeC1ebyGw0SpkRP
/FTnUG4D4MmMcuufgQmjeJeZrEdpa3aRiuutcs2RYqsdZ1X2cNhoaKCDmOD5zPzOAtanvS6Cfiok
s9Wki8XC/rQDcGKxDI8vWklZKlqQ3IRDBwlsymH69Duu669xOUGSsdEqykSt2BgwWfPLrecX89Hn
ctYaZMGzXsapF6si1O/aXewLAg0nowPe1l8jixLFhVWPVUeJmYKOutM1LTUxmkJFB8+P/p80XWUU
HNbLQI4jPP9AGMkq5u/rYkTQdkZ/5c9zaHfXS4h7tsYnMCrT22ry9P+f3+51u4Gkxbf+wd4sqIG2
NxPkcv5EFN/qRjatnpbiAZrEkOyK8u7k8AUxvPY0fu+EOsbUxTyjsAX8q4WXAqS1THxBD6Ji5xp+
xUM3l86PEi+erKHLCLYwSqxIva8wj5qNzw2A4XURfxXX0C6dXBPS1vswNxX45NHV2idfhZ9atuyT
BTC/tJZksq8MvWfOFVAVi7ZmsN8zQS9zT5wkFlIHyIQuif6jjOyl7DXk86NFnmYHhGReBwma17Xd
W+I7mjZP2P0ress5/T5lq5fNf0SLPGaTtyNSIY8dgJNJk83TMOTVFTvirwBlRXSxoBDvQ9JsE1j4
jliEpodFmB4DhpHmTrSDvfHeSGe9A74Wmqm8cHTnTHznVZlLc4gRpxvEVxhh5c1jK+EGlEqEVq1X
EsLCQcKPzsO7M/5A/0BFgVsM6erM5oV2OugoDigSPcizEvpu+xfiAyY9dlGHbNSmN8FWxiNty7j5
jaU1tGT6zYFvLEgW/XEy9KrezmwafjPfPZEAl1d8bzBW58kPp2Lv1I7CpQfUAwyHD2BJYeY5QqqA
JJkfM8vHmzSw1ac2muXUPgUxjvdHaBqlglAaAYOPVd57Fs/hWa509hBrLkqUQeD68nV8IPKj/7WU
6j+QXY029OKoEFRiH4pKCnsI7UlPwoQ9JUX1JPUS314Eu/9FrBcjEYIJ9042KpKYodbPtmS6+JUL
QXVKh3neNsHSXVcJIURdusrutQPz1RvZ7EdvCA/h5BrRQV5f0nhwVNjZy1jOXLATB6tzuxNryLXb
ZTsf16xBMDhj5+3Gh4IlpvsAjTXmTCSo/Y9HRdUrbtuagRa1GItmT40ZQ9K9hyhNkQzv/y552Zdz
4fmW96xLGYEqkTXxXiPMar5xo7u1dnBVZkLg7HODELIVyBBoaL79ZJMis7Omhu9JCP/AJdlywpaK
tGsFL5LennKiqte50SGe7gRRepbNqAJN6NElo8/iQvxkqw7aI81QzcjGMHuEVdDInFgIBeiLnjax
Y5GIF1MaWqHI7dzYwh21PLONBw7rkU4rzoRTZnKqSQqnZaBE4vKJjy1LnBpepMABcHZWiPCXIeuj
QA3yMLMe6uqAZMwp+laaufqyIHtLZ0ehZgacLoAile05E8BTrbyIK6u1J9J6tafVZnAhpyqOnEEb
wH3KGY6fJJhB7nOuqBzq8mfBCghh4W4vLBFq8VZX4kBz6QfGS3BMsWMzBoiNLJF1lkbIxsTNsgED
3U+TDtuulnJTBEiXMK9LKtom30bFfmRgVaOU7XjHmf/GOZxn53R/raHYi3W+ghbShrKF3/j23sOt
2qo72lEKoaIS9zmAcyDaiutV/M8GA237K66Z2ZdoDOP8hNcf+0YXywrVWQcvlKPHj0zKtFIeP595
3KOhiwEyuOqoezGKd/JmztGy87iq9f7jGUuzL3UeC5TtdavhboYpd6PWvuZSPEd5nsut7nK101Z0
31EcNHdijQOBqVtS7U966zbPbj/2s6KX8MTd0Zq+rK+WyobD6aI9dmoZmS8dMgcDJFI4IJquDx/A
ONFDp7rIUsABLjxhUKPttt+SJ6Kb1ACAquUl5ZyWMYqYvfJ86Xf915s+eKdeVmo5m8M/PgTzJZej
LuEhHoimh1WIsdGE/HUXyn5A2KnrraNRqZO/jDqubPeV/f5fp17g+eQac7sfBtXGzoNUEyt7UlHO
NUPZSgatRDXc1dJxURV5/oW+wys6EL39h5lbyWY03J7TlN72Sh6m5u1RcULCo084VMawi1+uXA0L
YKcUfLfjQGej1zL8zm7KFYINnVCQ5376+UDG0XtuLYX4UfP7L4fhVwiUJuftW4IhJYLDCOpg35s4
vIcZC/zzVUx/PLCIvxziWGcWhJVaxKeqHbWlNQ0cp1S45CH5ETraUZdhCI1nMUe0sSULtf2L6e/Q
/G7CXKqG9hQBAL5tDhG9EJNwBrisIePzJzGJwO4i/NT0jcLWqTYecak00Vjr8+YunLEiLmfUbAVf
OHDQPeyxaT9mGDCYf0sScZKGlqG7srLDCBTz8FG3SyRtNW20XrAPLe0PF9aGMVhbtWCkd5AiV+3Q
YLev/RjYMrXUMLXmz2zkPc+moj8+rw2zOtb1flCPAl5/achn6ZF3wkeVULmqF+RFOqa80wUWidpR
GCzhG9QBTo8+KxxGQgGnq10KJ+th3GgG6ckY9eFc93ldchVHJdYtwimxjQefAU79sCVcVYXfycwx
SPhAZ44OA+Dzkd4PuRWGw2mHFHSY8t4SLifxWl7FrG7GKmLejQpD8e9zJaed9vUvcqsWNfvAJqq/
D0nO7SeeHUS6WAT73Oum45sf0SKIYIZKnswynk4FdLjIy70rhJMGgwEeHy2j2TY//0KP3rUb+BJj
40sfcRm/xS5rZwNg32i/JdoCzo9lhND6JIczKKP1Kt4WuDHR0LetCVkD6i0SIxzuN0DicWFhYKal
wS0dOk+jyDvoIp4724GT5ytvvMCuPIsL8qP+JyZt2FlNt5ih2HOjbrK+RgRR6vyM2aepgUnSqwYN
DA5hXaD6xuMaOneTJoSfYDpbGw7GjAwfnLJdjdkCyyi+iUBwCJoyQJQ6CTu9IG53+gG9EXLVTQSv
J5IthjWLmxvS9Of0xADFUDc/OlSwgBVXdXM1G2MDG6+Ji2Pvr+djNUEZz3vNwPHSlOCcZc+jbjBM
B0MyMUbOTq6/mU8nE1wILMK+oFo8cWXP6GIpBsHToYwedA/nVx7uKvMCVuoxyzLIu7V98zB1yhX7
LNQ7MqYkSRwdoi5sw05C+5LgGkyhEfNNykiT2oB/mFNqQqBeKscNuEpPZRvWj65jvgAWA2Bn2bnl
BSibwp/LANmD7zvKyjQxWrBK820WKZUZGUi6socI59QTusmq+g4b4siTVQ+5sniPe0q24LXgkapk
wSRYz2Pbq6KJUGOaExjfYqn1FfHXIJdUoeem70yhjvCpXEYMMsRwP0d10K7Lu2qdZacf4gVPlMlY
u22U4Wa/wHrBqKUrm1jzLEIVZYAt1+DtiggUTWhZktx6tlUDYzySyrDoTW/QtH+NqOoHxQFzfLFZ
iSB/yKc3zUOaYQwdeaXJnpDKiC9iTRRlBfXUyzmFXSbe56uFr2ICViMgrdYzc7IWa5xufDey/MP5
VVQIYLzVH1pMoFE/76MdNyvS/fpRfdKnP0x60KADgjNyEI6KsQwRvLH4mimQb7tQK09See9Ap9Pf
BZigP1gEiV3mzuPYgLrDygjOsIXsCzVErgUjZg+y+IPb4/Fu+uvimDXxWJb7CqaJh1mBZ8nx8Abg
diznuuY7ZXSMRw+HWweezBYVDk+z50kvKm3Sswobp61N/qorjfaGkt3z4b69f2GGl+/XB5X1Vcut
nwsV4ixb8UtqMJfi8KRvWwVXViMU0aJdQpmw4hPvOUHGR3VI9X6Fon68s8dIjBVty77ix2Mo7hLd
AadbuglA2Aujfnr/HU7P5G0mhdJYQ2BBUUqFLl9xUU7Gt96AsZK+U1xbT1P0XH1hOhrzXrXcJkym
3AAXm3B/17Yo5gwvls4LxBQwoRXVbymk3pUuqI/e63rtNOjdw9ldSoy5Us7Dc57GbffrG/EB5WiO
00uYrLLOyHYQu5TSFs36QXgwfoWgoC5lASTsKcTdUTkyecGAiMF3wWpd4Ubp6sDqhwVAcu9EbeE8
ouHHXJyJwbb5/FYgW85fT/2G5FMiQlFqMSkmlvJzV/0mYpJh5RKZTJCcVu/Q1NDHhtC2JrXSH1q9
jlSOEq03rqJBwk/2NPNb2tPf828r6dM9k/KiG8BLWDoCmkAZ9Gz09n63qXw9kLIivXn2HKKlYZl6
BjzaxACsZaWfSgEC9M2cyUWurTxUNl+QzI/4+D95cMGkLZFe6QAKDMCmFEchFYZnY9Av06CnGwsc
YbV0GbN4JHgNR3ymB/xKsedUYA8dq38lglVI2kS2VYQqIxOy8l/khOtA2tMtqmvYKxsAusvTFHGQ
xjHFCJQ2dnbXld8g+jS4d0V30kHacGjoxedwzRFyPPAvRcDpmf7j32GWrTdlKR8CxTbv8wSvA/CF
+MlfrOw3boGLOZHB12yLixn+cTQ7P6jr/WXU60rK5ad54Tr8SyMpO/d6xQr5PAw6Uz+ZUl3bABuN
R5g8UAwfDnuHvGyoyIi97Y4xKnxbR9Oj59f4P5QbNHpB7AlughWIRA1nlS4Ly7xquvLm08nsAsJ2
etqlOYNFFHvYUG3td++6fvt8sna2S5m+0A6CbMklaM/410AK2ENBnEyAlerHAU8vfPBwTqi01C8g
wNulgX3f1/6Hssuhk/hqEaDTj8AQ8ccC4Jbbpt0WYKW+xtHEgevVX9020imtzEQV6/WjQSWBP5Za
p18JKuH/fhlnX99RBIgemDfBmINO//ft+TsqT+CFCr0E/sLopRZP7GKCCdmibzlP8QRSPjN4aY4L
oFChzdQMhYTrOkyvkMge45cetVSLnXw2qP7GYYNPuDg17RFCwwgcZaRkh+QEtp/SrEVKQXotLJN2
GVBLM4S2+X6K5vD9NNu1ofqg//K9vY8D23Uqd/0r0r97iam3YQqO8R9qOF0oSp4ywLWebJbYDAyQ
i9B+5mEmUPsHr1Cwl2UNQyZsMZw++UV0zkrnvtKgGhiA+fDSKNmngQJju1H9R2/yJJNrh8Jy/yN8
N4H0B5lJyT/HbPCYqaiqxmAXAKDg15QwLZqlnioQWnWrZJE/ZdDiycElOM4xXorBVM19KAEQq6OP
LroAFe2SPm+Ufw5q7Ngw1U4NZq7CBsSCvrY1tTWqcYKJuhFsUzv9zKrXs1B99joUz5iATmgkbI+T
dVWyUoDBbhmla3KcVXFjrKlsfaS8eZfV97C2ivjjWuzxX027B808ZTGlhwg+rsCKXvNrs2/Zi9Qb
7/PE0qiuUVLpTPNBlMsZLuy74CbvoR7PvknRatz/aiNo9qKj5LpW3nqv3b6m9Zj/hsziVNZwK5X7
WX3nkRnuRjn19CL0mf5QwyFmffmTGq51UIS3pczfDw0wc6L7XS9Pc1MysrrPZwMu9ulE0Gb1zkD/
dz03NyE32+GDK41F06AieFcri7XjHCHssHY7YyOfWsObaQJfartQ1QxQveX66bSyTovsywTjN060
d29ZsfAS7Ld2uTv5diBiisgwR4rcPQ1X00I0tWvo+XloZqGyFwDrC7BGBdo6NdOK9RlxYjnSXOFs
4ufvE+S2rWgCOB6k6eI5T/uNQapBtXhGA5aMKO6l/oXkQweycEGg8GYN1qAFO2rKknwLexteoaMI
vKRimvtf+zLM6CfSk65SoqQnfXoD9TYL0sux08PUmIjdaH1RptPXYIGazlLNwWbqrvi4hMrpnxLk
aV3CUZwid9rPBSk5QHciRJPudvvMekQqs+lLQ9hWouc4jVAo+yPPxJ2hMnJWuyR0FgKSpJpgVce9
FwBDA9mgHA35YZ+9ILhQpgiu7YMoOlHpWuw+tpcWFD7PVKMp7Gec+DA3oO+f6ioS3hBnG5p3ezu2
e059BK9Sfxg+WT4B+VWefsYUOqBYtp3hHJTn55bGrwSJJZ6uR8RgW2AMbxvU6vZVJTCitaT5FDFL
gf2clNxn+aFIhmBe4ob3XaXKPM5XHkCbo/u0amoIW5GDBE6HI9RrnJ/wPc0xwNpqkXJNE/gkkjgi
/BBn3VQvcdT/ocyTySOj7HHsbuEWTUZqu9Y3BZKeFKYj5bonXbOouWp0ZUzigyXw7FhRhQgA31rT
qyKcmVqVYR/ktZbzTOL+OpRy7Z5s3iHHTA4TqW/Z8TbXpXmK9evBZChCcRTzYH1fwm9iK2B6h3PT
lTjVJfSwkiD4uMMaGFbwo0cDUgT5Az2u3lqYpciVlJFc5mctpyVqYrINRaPrfUhrJ+OmiFp14G6+
A1+UpA9DrDt6ywAjfTbcZo/orA0xB4Rz/r34brBTZcZ00VrgTXZcBcZ5y+KiJJOq3UdfnX7fr9J+
ivY0zF+OcgVyOTTVHjrrvzW3TM4m8+fj+v/bJEG3U/wXlDYbnRdplOZix/XgXo3xMEFuAwt5KUKR
3kgUDRPEp6hHNiQV1rNXyhjXd1FebI8ozUhY0wzdujrpHbPJ6GxzQg2h1XjhcK4WUti2zRydLiPB
ZV74MNjdayPRmlUHNK5OOAeKWeV9zY2RpA6IgoHwZ80kMxi4S5FBmFq6mCbsYRkLNqvZDiQu56Vs
Yf2pccjc0DboIQK2FRKu+92stC7ctfoehQWltpl08AB5VLLOM81t4XbbbHoG9rzDIhYdouERhAcd
K8jv93ZRUL1XCulGGX5qZC7TGQAXgQVZjx2C8/7WcsxbYxeeVlLmLXoyvn/9jgQnnQnomnPeaeMh
q5PvncOQL07tYN5jH3TF7dv/CTmpJPY74vhlIo/mkc1mIsrFXiAPq4GXep/xs3ZClS/MjP6MeVnC
s6Cca7Ej3iYMlcCxKN1SzzZlHo1ZZWMoeJRM3DVuj5pWUSkfLcLWJL48XTduPz2j5l0ldy2NxUt5
2qz4mV+DEGbPRmjw9MjvWTVwyq77GDj9xJQz1SUtNc4q17qUmm2I65HS94oqxOo+umgbgbFXOUNB
euoAmNTUD95WyoVUoVTkDlJQqDawIDHhXV+isL8YRwr+LVSmBJ76YrnewsKGSYcXxseBDYVLtm8O
+PAY1FNfiXxmNVZevLzp1fNdwo5CsPIlwf8NXwhmQGS/QueJAyVhwDPyAri4uJH46xSyrdldMQZz
37xsXz/nLWxPlqGGDyzx9mKoWGpjlz656xHyeo8X/zo5uwNW3xq2f1YznheE0i4Kmbi3MnS9Ls43
6BPy4KrQ4Q3ZTgknqItTlBSUTkE8HrSf4Y7rDV5qfWyjMUIJQrOZaFkw5eXAtJ7QAYBbXbBjEd+x
kSVBCvXt4OoD0D95TmT/BdA7XS6FgklUDE8aKAdqEdtlTBcUp6b/UYtQueQjCTjvq534mmwL6d/u
rRQHab95cjgmLCo23yseaW1mPIWKdJMOBM5gaEZ4v8dHN7BeqriKOUd//+T3te3AkLVV0aQqgugb
ZBMWwMjNGf0a2AZIv0y+tM+gPBSi5yuNmdWXZyL/38TvvfW1HbaLb7T2D0Mzl/lMRJalZbm8VcSA
ErphWB2jWJtz6jYMm4i/yFmpuYZhWppU5iMHOTP9uugjTRbqJyoVIiGl5QmFgMZgRxlHiK3/M0nV
BgRnoHJ4cwPPwOnjeCu9Ub7HOJvE3OIg24ZOgl86chm79zy3uSdZcUTnkCyo89JtT07RzdD0DjCt
q/mwPLtfBym3m8AfwzLxXBFti0zwogyxMAfvKf3feNZqv8+XvAwI3YGHk/S5ccxB8lcPpRSJAFF8
slEH89lMQmNpr3Zo0WNWd9xAO1D4d37cj3msfeijM1MNVsorecbB4UXb3P4SEIBqlVoARi9gL7QK
IoYgNR57qPtPvpMP8I6TD8mJKkJ6TKBXy42DWigJg3jrZj0TZO+RkrsWBnNqK1JfnDCcS8FL0FGs
YXnOXM4Sjy+RvsgYHoC46RLF6We192dMJFIPeVeuNIa/nTrpbr+RNcaZk1dlVwzUcMT8ZElRHD3v
IWTlS9iyxwzGWbEpONSRAKgjuC2DWN7Us/uYtOKT5Hi/1wxzGsZUWZc8yEPiPbeWNllbFuzX269w
4aFn0ZeCA3Y7l8MQ0BHez0LtKiSqmyVeP8278JuLK2KZ2Jz0GLikDZCzKUSOHB/nXpPFc8dZENwN
HY0fYBssX7P0j8qK7NqIfvXZoq6hIZyWDeO8aQZdL6BkmEUfVsRWBYDKHVAizqyEeM5sE+VOt4L3
I8C5MtYOCWjpNaRbatHgxtGQur93gH8crbwY5woGWcPqB3mkGEgQw3HOKEM6xNqHxsW3JzB4qgAO
kFCjOXXhlgzqKPIAkd/PP/8ymFOrSEaUTe86vwSAYdRFVd2zVSCpV47Lobm0jWUT2QPRKShYpHG+
jy5fWN9aXB5Yyu1aGltzC2dVs7E6wvo9gv1sYCdE+5RXafD0DeJNQ5os+kw5fM+KMlm9F9TLlhRO
cLf68LfIYuMuv9j2qezPmm9Ah3EUWyqWHs0fvF83Fip0i3S0PV747+EAAp+qeDI00A0fV9ai/SUf
/Vf71UWfbcn1bY53ho5zx597hedqNIC+k0LEOKhhob4krzz+ZDGJ4rrvVbLbFG3sPfhhgLJXluPA
rLMLOYa6frJLed+0os47HFQdqWyVSURnjTm/5yiHZrAo/Bd+whazSojvzSSqcak8PHiF7G1tcfzy
8miEA10Gr89j+kbcPzrTdreRg+mhK92TZDWfxNWhFQBCg+eoq4BlvUJrKEEcUjbQ/wLw+2dd8rQh
1Qt+AtrDcQ+FuTgXo7Rb9inASxhcLbVaWpySOV04WV443jDQNoE2gsMbpS6cF132dDWrncK5NNom
7slcCP16EaO6Tfj9yYDhfDaTpfCivalKUF+QmaHvMf41wEkeokjVsAUUWs35sBUoG4dX6HcL5nTq
zImz2M+QLeG0yPWh2tr+hjpfayLhBamcEgNDR1mM/tJ6gwqBW+c0oJHnUls+TupHqUUM6dL7Qr9Z
X6MZ7MlPRlTu67PlIkaSXKmmKegxy2I/0hGiROKf+dtgh6RQoPqg+iHqW4CgOnEFmRdDMs9khDTF
fgwBjt3RcoH/LIPfm+r+nQthQqUET5EEm7ccSyiwZt0i+AjuPzcWwPpT33MY6tdtLYL25PJn9qJP
6g0/6xT/EZ7k3wexod7/iP29VZ5U37Ry8fUgXzB/8Z7OKqgF0S7XECYtVr0HGhXfWWYJtIBrF5gR
YttBpUK1PlKKsT7nrcC/QfA8d4U2MYyyU6MNvJnMvBH9xbIEebTdXLKdVepFeTvEbcazcizZg4zp
2xZAOhqKw7C43ZKYPU4n5C9QaOM/SlRyaQhRj5MWSMDWdFvr338a5CYP4S4dOq4J7uGABsCoMALS
psQL4Tl1BeM2W7iC7Lpwoh7ByXXktk06z3hoVfWLmyE+1OJBzwoetB9jhX1K9d5StzjujVCE+C9A
zldeEiofxzRBxyWwANFWGQzBhMio+1iWvW4vjNPXaJm/Zkl9zzr4xqM3m49uXp3la+TWZTjys/G1
9niu1SPUAT111MAPJFjE9eJahodbezTSM6rEyoPfkJxISo2r4Ro+7Jzb7g+IkK96iK/hNnoQJmA9
IPBQqRrQjNocJ0bmfNVfm/L1N9mm9H6NZ0rGDnVct5aJ2ruly+xRMz7V/sVuMJqAOJys1NajcCkk
dJcpjUI0m3bCxbr+76vC1Ph4dx9Z6YTG4DyUN3x8lI/KPJ9D5+pJdSUxHV3SPGI+CnjrGFHI15He
ocbTWxm40gZZGpEVVwoItQhYIVcF2PAWhOVMyOomACJbrieTbDu0hFjcC45vs1t4iXTM5CUkzsxH
dvQESa8mc0MFap393bQGQDLkayg7hTBlOKb8YbNKE87HrQGcApdS+wioJP01a8OlAV2aRsG9Qpxo
VzjYgwKp+NxP+48UyOXQlVS0uEdSGx/3QL8Ienj6qA1kfGTNRAfSBYKcBexb0r8ESbltx/xe8aJC
BXOWi+F18PuVc1AEslPrMBJFymS5GtrIl+FedOvNpcTzaGm5yLoHnVXCNoZOu9QPn5txsB5LlVqb
Dat7Z0WB43bOLnPpuPGgeInGtcNIPoR40sj3LXe57zJqiw9P2a4oXPf7jJFjKb29glecN80aMK3Q
fZv61v37x69CBnMYA21gh6xVkTbsaeHWxIzW4I+zZwZ+9ivRQkM4mVV1tI6fwNIAMJfvXPkexFdO
qPVi5obUVWMFejnUQybWWonaUKsWNa7v/aDQO0m8WhRRO8ixyGvMlGjDMgPGIvvaKYt2ZjYix4hA
f5QvH4b2wQyqB496fdsCMDsBkb9qu4Z7Jp0Rqm8TqCuC97tqEUpnj/AIy1H/sD4Ds7W+5XbJ7se7
OxZqJQL1tFZr328Ir8F+XOjuPXzx+ooURj3JdRGsgHizgfyIGTt0HORKfDB0Xme+saujhguc2vQx
+BGSzDFeJTW9RX0dSzf87bNKusDkviT8vrh6Zwj1oIrpey50Mu17kBnG7Algzu6PAEQVa3PoWhTi
mDlDeuynpf+XdJ+GNUZGnjIZmQc9Gacm19jXzs1GMCqqqKMGwdBgZRFdqPC5F9URo70OTD4snN30
khJRWcCtOnecpUZ5qmxl98F4LA7RPBHjT9l9E+TnIL2Gxp0vwGZwYw+u0Vv7C4uGYg5lraMcOOgD
qtRZPzpXi5oopetZ70SzSK7ntY1PwN+DhjSKqpQcJBp6p/YIC5nu5aaz7Wmj70BvyiP/GZRKXmjC
7HOkr4ytV/JdXPas4thXzCkf1JjaaGG38Yt3uppH4y8tizGWFibXpfx9qTUAYntUZMRPrKrKYZJ3
9FzcIQaEBUnUbOUN32lctySvUieCbAk57IMG52RYOY00MduJs62//oOpfwO1z2ANBGqIpj+GvYdu
04SByaA4EmJbXwmYEi5/Y0g0R7/8I3/f9n2I9jH9N8LhSDQdyTrB3MtSpapNezSXo802GP+lsVwR
NWXeYsJ6V80B4/W+lAnGmpsrb86OZ9mxsXVDKs1aJ2gzwo3KCVPfHWX6S7llPzkT0LvfQyceswIO
kiK4hYV35+Z18vS2vuwGHkLWc3kt3AEuK28cTd5db4VBRk0spfI7k/EbZCWhA8P4yHnsHFd3NaeK
4owWjBr4JDeu2dYOLZCg3vsPXzI8O/5gT7pOvgsqqllfyZ6j7kHkmtvXi/xo26pUefLeegILff5F
VfUwAeXI1P8NRXYlVidPKxXU8+PZpeDztkYKmn/uH71V7oMOhy2io3Co0z0CRoEkyYRDTsFqCr6/
9R68mam1ujXeDDtFlMuqzcHbmUkxwqRvvbgrZnxQJox70QLfvTDHfD1YLlPB+bZ90NReRqzuDb9R
c77TuarUZeYTvs09oJcg0SGWfT+a1oezfHvyF/84AOK8H91Eft7QmCMRzw6cD8N3deJ3lK6foYoL
XUFAtxj0XWk+X8iC2YHSShtuKhpnxMO5skmMMBmhAohg75UV77FzmGjC+nHM8M102vj17EYjYFsC
nCi5aExALTsLKbglwU56y/rro3UqQUODIyVCId4PrsrRnYLVicXxAGsCblaBocP1lGHMmjdbMmVk
T4+NCyOYzmGjw6/wVw3/YLx7kRBl0yGheGeGPY929dtJ/ygCwsqqUCwNdU+Zo7Ih+kM4H7vwsrAF
1nAHe5/N95u3gSDCR6B/8ZUwLX7ZX/M3CPirQlAZrL2bVyAiYhErHAadaTpeeTA2jNVcTN/tXgzO
PLAuByrjEYLgDN2YAu6tMyyTxsgTt+6xoUGaEvD337XLUiCu47VjXdCP+ovGezotvPL9wekf+iV9
9uyB+mwkOHpiLVolKkOKcYq8CrrM11w01YbVAcKOgEcCpGYI8NC9OD24TOQSDHTKLOsc52rto9TH
S1TMSVrhRPQn+ECqSrfGZqVguF1xMwT+a6LdHQ7kDoXmO7Yg9Tnk3BvGHsGiImv4u6yCEJV6rNyV
KePaRxikt8qx1x25L7tasok0aCJzAlriAkdWA6AVwaVSgD2yXw1WN9CM0JxRmEz6kJ0uWVq5DLqC
qAmczN4pGyt5o6k+Bctk1uxDZp7g3GTzv5s/kDbEXbNAUIOwdPQY+DCGuZu0ikC1SrejVwqzoA7m
O+eLv1+C7qt5G3FzOCA7Ybh2jjS/bsDXFaGekl5ZhCh06FHbA3NmPNFiQW+vI6xSu329OfmV0TlG
1j+v34UfHMCXKM8ObC4+Z1g8sp/BQuSyuJCSQChy/ZkuQP1LEzB4ldgIZw99Z91ljXqUiRAaR07i
FmvofYMzo9VzTqdtpTfJtF/X4UoNWuZ8ZFTqAwPrh373iCxDoLz/7WnzQR4OFU03qbMojJ2ofd6Z
xPp/qN9Pkggw3oSt35ClPsENUb3lxn3VNXRe3JzoEUUVNQKxwgrmbkzRB3YsfcO+nfBhl18j4NkR
629OlW+WsANEI6eBOTHYrsAJ/JF8/Ffpt7A1MCeMHGTNZq4bJc8LEg/Tjb5/JYemjZTke0ZYAMo+
vM6tkN2xTf0+KyPf4AUVKI+wAvpZ4hYAbp5EhUyKlAYDva5ixDhkNgZUxwW+oNYBfY/6tXlIvFN8
DA1H6hR1HSqz4a9eMSq/mhyn2MAqn7UN9Wn4iVQCtQUmfF455FtNAYr5/T+dy2q8Be4c6QlSspW6
7up8lB4NwtuPw39Xml1BIxLYsGXYB7eGoDIyYPX3RNhotaLmc0BqwHZMGBdxIzLIK8XJb0EF7dKr
BXtn3a/UOjccS70milLkG5z5DAbH3MdoCCDDt+B6SifVd93ml41hfvvLGkGJOCQaFbgrgTGj4YLJ
628o09nyYlTXly9ZHTcfsdRNFigx1KRIaKlyVM0D4QtTVzFXnKs9sIGEfbIphQTvWEKRiNtgePVC
ZNeVzgL9o+7nQ4vmLvwcZgQxB28Nel+mJ8xNtGezdepfj53M0OQ48CogPQD+1IEbFCO7hmxptU8K
dmw6j7p03HM2o2PbPTMpLYJo0xOTmWiqXX+rLyZp23IJ6vwkvCl+EvS9q0UGlip7BGsZQUWVbTO3
tGKulkBMaBjzNrCYq2IZF7zFd158U4maKeJ268nm50gC5dpQ7PlZpRLHupEFIYAhQ6nfT66xyVb/
D3y8pnzl1ftjumn+lQHbGZ/JycscKLGnUzU3Wv+RpEyj4/UMocjMEH75BGoJIT2rCB6DkVFT14yw
GkdVi1AL5gcsllxD1WEYqvBtuqeS+FmwPsdfoLpLaVoje7ZkBGRleT/Bpyu3GMDBbazpgMPHPSV5
HmeubCxzHI+tG3LKJrW+wl4gXHcsUhA8cYLjT94h0yayKrGpSo3kUAhMVhK9H8d6i6D/hI97j7/6
UClW1cJbwcZDYBTLoloEzYJdeny2ezeJn5LslK/BgMLqXVhCDTAvy/UkLwu6jfZ6L0ACefTVRmSE
f/HtaWlPpok5grM7Z0xnKEsww5wzQBjEUsaEbvwTc84vjAygnQUrfdwNzNUaQNlYTOvS6ix1tZJX
B+Nxf+IxYSDb/2l5B8DqJEYjNFo8txpTEL3jOKzC3m1lmVY58LQjoKa70cTC6oruKBW6wXMnUeKm
eQ8bZqkkhTUsCt1cO5TiKGzVXbmhiyXZikTQYSkTzWO6oeWpc/qpQgeSnhLntD0Abp0caeVDGYSC
v87L2GERyZj0KFh7qGcOfdDimWOgRUvRTTHz+A2Gt3m44kPjM5ADyNimfcSWM0ozfrwuBXvhOMOf
Lqc07VFTXADn6ZbwUHk+JgTrcduIopMfBS35MQvfFATEjCQzHQllAug0IfFSJiwRJblkbAZQk2YW
qD+FZ0X7D6KI6XDXNhf/hywm2eZ+faxlpENQQG59Wjax3iT171PeWwe4IT69Q6+hvwekA5VMDTMk
2XcyS2frCFG72Y9AXe6ShyAPB8C5kA1MB4YZshcHQeSz8pdwowv/gPOhwZe6w0lMKFVbLRFQXnW4
Yd+mI1h9T5btgX6AETkvMt/3Ay/7+7xp4n8/xxxsnp9Tsn/KETVuseFcySybWs1uYXzCGEdS+WfN
SPqK/K1ZO3eBLvkdCFKgyjH5mDuVOfnBKQClo3YNBea29y9HAindwWO/f7BRi9x0t9i9z3P8nDqC
0S/dPtoVIS6ygBzi8tqCLCnvqbFGCiHdECL+/JILmBxVW1hyMqFXj7Je4O9FwFmQzJ8URJNa02b+
Z6noT9SfKfxl6s2y82bJP8KXzBl6CAj2rFs5BegAIFd5y7eGgw3Onaw84M2zkY9f8XcXl/1OK/Pz
jLnspn68q5tWQyaxZg+JZHcFrqE1OQ3ooTxKXCsUFwSfmgeSsCZYwf43W2LgDfcO+eOn9Hq2p2P4
avBuPDLGBcdgcfbgRUGLJQsZ/8epgYgeP/+/phkqhLCFpSZT/esp4bw5o3TaUnT6VOqzKHtA15IL
ZuTUA9HYSRm/qd/lIih9iDR9D3qEtLh1Z+YMCGRpGe8AsUrFi6xrbWipeW4fEockxeMewwMMMEKG
Pl5X67I84a4YMyaszSdxH75aJ8vzYckKnDGgkIkd7yikJDeNfoLlx1dqa56Mro27UeXD3skZOtvg
hp4FEsBVf//LmkhSj83/iIma7PBhpixOSH6scwemAjDx+VgcGTEXjAd7ZIArqy98kgM4Gq7mq9E8
oMfgsBMquJxqszrEpox9ZMkJPLh90VSPsR7IgHE9OtmJSOojNkAC4ys85ng35B/WHF0TjGCxj4BM
qPTU74ZyBbrI83q/CdIbc1yBp1PDBtuhkH29OZ/oxl6jAtLYWO05ZdakI2TLVrAveJc2C6FpB2DQ
P3km296bbOg8EuvYMo5tgzh++TIgFIo3xZy1v4YvbnIwUrH1PxThsh73jcg8fELsa6YbrSD/LvQ7
Y5dribqjrz0tZ8Yhecwp8BwmZfncSZu101maOkVNaVGqF0O+OAzZWJiCjDodkFkXKq99t2XklaW8
RigITv4QkNmGEqzS1f10sL7Fl3YaVEhrYwe6XLsDL8X7n4IjUURf6upWllRALZy5Fc++sBZBkIHI
OccZc6xi6qoVvUkR7Jp9rViKVMlYGmG/dnR/nnt76oN3wryp4X/6m8EOypPyiz8eB1OWSMFfLYFS
lr7YOumr6/6S0dhefxkJcNcyXUUHOQlXcz8xKPpYDqkGPa9xev5M/Zei1JCJEE0moFGRHMzIKbDH
Bdwo9zGvOMHCfEuXSSnnon8J0Mj1GcISoKNpxdkqK62Qdf0huzbRkZ6Vcotaki2/EAuAjzkQl8r/
tTXKbsxoIbl8RA37JQBMB/9ieON75No0p0nHDmVmfa9L6GF4bKYoLf759GS5EMqeYK3pu+HXJxsD
DGw1QWCx9jHmBI5JMokbNi7boPTrD7z5kAU4ZVmCqkjg2uQVzwBWkSaFtx11iMlPXw/fBEjXCS8t
wvAptftvkdC4jkcrJIafsxbV2S7mRBK88fG3WEJk7MvsaArifjdfLi7POvgn3m5vniEi3uLH2SIf
tcxRGYfCJl5Th9PQjIDOpGtFxZ1/+OVhFZuVQROXLNBvo3HRwQkhhdw7vj5K8fYm+JPLssagvEji
oCYF3NYNoZJZn641eJug6A7c+JR3tMtyZ2xs+rPRuz9Ply6+pAzioIN6dqYKhuNSLpZoXAQTSTzp
4Cyy7x/RHjsR1vFYKYGoJv73hKQB4mRlvC1xISkAPIEJvIB89RqaAevPMlKuzX8M6B83Ia5P5SAS
RWQjbt2IMZFPSWiI3IqfNjDXx2g0UnL+jGxLUv3P+JBkU7+JB4xLkCA4qNoATLNdid+yvy7xw6pz
nn6rAcYsqcOHwiLMMc7rxDaEeO9pbeKENhlHdfKx+dOE4w7fapnAV9iHbBdrlvFhsVucAWtPAMY+
mME4zAmXXHiESftgkvDzqAhQWaU+u6BgEUc6U0Mrmzc7iD6ZK5LwJr+vXG1NL6LDSZJjnOWuSWZ6
JK70hT655GKBc+jvol6B7qwUTl8Yympawb3HNsOcEG9tCqdQOrmx5D2JBXyvzCRi5nkbSpeNKWX0
xpbtfspGfLyT1DG6Z6f4bKbBq7tt6G/Iy6yJnxW/0n+iS3kZ2S/uI8UTqdciC2NN2CDFSEGSsprH
D3b10Gokn7W6DCR5rZ4e6vTautFatB87XJo0gX/xfiWeQzWkDySFBIQSFRLHKfpMbTbD2TOo2QAT
YyYaMEJ3EvX1Z2b1ae2IQwUo0uCkR2xt7j3kt/3UI18OvHmPAtZo/J3QCI6CYoMX4Ip98A9O1fwh
I5nkVT2c+cVvNOj1gyOcD+/4bmnlyFz7DUeh8pEALoFyCL020e67o5j9cCr6+UhcTE/JIIe+Lzdm
ddxigPB0CaMyogR1QMnburOYDs5bQ+r/PqBgDdG85W+du7DAEg+2WwBceGymbJxDPDeKyPRLk3tK
qi2OzOGdkaWxuXqWSmoU6KU6ztG6mZtvU4ZPa6w2ArRK/yA9va07vekj1yZAWcas5ei0T1Z/f9tr
O3g0ghMZdoI7S2QlskHwuN4VMM1sXVIUPLXX6E3DZNjhRRsZ8iJx6TOi3jJQozIOgNmhk0gOkx0h
MgUzP/9yLiln2nFiNsSzwpd06BK/2rAgGHieZI0zuCW1ZwMChKLuKWG+nzdB25e7w9zUURPIYveD
Ck++8Dr+1NDOun0pTF6Ar0tzJFbu5+TwKqEw4KyQSbBvhpuuu+swEznTTkuz8WcFtvTNTgbPczYZ
DfuuTc5KeDN2SfejKL+MBUpOox1ZK6oX9PLW2PYPc6yqk7dEGSTXHJ5nkYdkwNnNLAqoNSRFrcoJ
Dhg7HMoR14oLuInquMOoRes4UH6pWO4MQgn+ang5y/v5+OopchU9Z1vukeZEt4FPxdG3EMpdc8xT
qWiMh/XkesHeX7mY15K80yQBvRE9SDvPhtKWb6sI9vOsSEkrPUAgIT/j3Uyidxfhg6mKdoPyYviW
GMl4QUyRxINBobOvxvUSkph804ozLMQE6AF34/nUHKZjczJN99gLb7DKaIeYRd9jB6PxKANc0CpF
SnTsRBdyrHnOHJtVYWnE4OfmnZO5/IM3JcL72VCvY8nvAhqLuTYUCHv9Hf/9cBphNaEWTHb84DVL
sg+D/6Dc/mkbKPFwiTGrxdpNipqHEzJ9G1rWfKa851Ge8igc+tkuJm1nIuAxpCo0WFBcngeCbqTm
fGeQpuF8r3AwpFJ2+ztuS7C7NVRCF09uKhosMDOSlZPnwxv5ZMi9XVHIs3OyaEjn/ZSqpkpIenqZ
OowR5EPK8RC20bvbLAwoqcA4/G46k5NvjbuklbGAijNO+2O/ZTQGTDtMwDPC0gX7k+Bs9Si2xHnS
dIUGZV0OMPNby0pcLSfBUKxpw7CXs9aS2xqdEQcMa48NsNEaRvWCVly9QtSlrbib+4GEpKHQwExD
Q5HVsm6Y5Zmunoif04kjjWe+ZmmuFGaZnDptu/vO6tHzyqCnzRvhAaCY/AdJHqpx/S9H1bJyE/LT
TY7yKsJG0tcHHzzM4JkKNU4bl0+ynylvt3Sr2SOg2zBLuRIALKfrwtZVxmnLJ9XCgtcON10tJmV6
Sv+k/sM0KqtjC1LUSw4yM2EakZIbpqq7+ekyUDP5NPSmwvfV6CvKBd0FQWwHrUtrjRgPqydCFiKn
fo543ODGN7+3TU/uNitibcr/Z0cFsmzPKH9Wv9cKR8c58hMuQ6Vcla+xzWc6VLJhAeccBrU0q3OE
7KvMBEFqxVn8QgVBHyZCyQk5K+Rqqw50V/80Nsiwjt1hRC2GbQYwWoQqDeo9FI6lx8YOYpBX5mRe
DLwKiSPDwGU3W7RZvtAdi4i7slDtoyaFkGmKA9y6T/AxUZWXr3wcI5dzCezw9Kf7mGrFJwKYMkbt
kknVMzQ9SzMaVFdow3a9Jhrd8HmQ2Va2Uw4+6UiK1mIYw+289fY1XB110kDh3/aHglGMOAdFj7Wd
dtFwRlKNpcPpx7Gzb4+hDTmBSBTABL0c9aGBvaMO7xBBrMBBMrLej4N2L0IEWi0Bz1iwjcBHQ12o
AGSyf27CZJc+QkVluaCYc2s9plGK5G6+rkeuI9MR4jKEARfmoGWGE7Wg0TOOTCoOJr1ZXE65Y2o5
nP8kuRIee2NayXuhQustuiGQyoEeUa0llcnKu/5afKD5zN/z5870dupbA1fuH294Min0mn/f8NRZ
rVJdL/rJw21b0KX19LEkwg4Q0XXg9x0c7ciWD6tF9z0VRyWzc5qapWqZ0k38yqfIzF59nur913eu
yB79rNnncKBV/aK/T2r9eCdbXcYR94WuCEjf8AMGl6hodgZg3fGwXHqyX+2c7zVmINr/6gkUfhBL
HF9iPZ0Bt/0CmuDlN4hrQY++a/DTO15BoKIZ5ZycoNL4LXzkDsrSiagJMCOrdP2b7tcsnJxJ/OXX
hQZlhhslS9gmXvHWYiLX5DinfMPKBNC+Ruwjcx2sAW3xv4l8/Q0+OkJh5/RhzFxwvWA8KFQdiy31
seGgfYANcadkKxJs+HmZ8zTW/m0a6c4/9WfX3+zSe8aUYc3EomjXdw79Qb0I0ZGE6Sm3qYkNaTAS
lsSRsvF1rRZx+fD9qk6a0Hah4s9CEKsYE12ByGSjE8cUVTlS4VxR9+GAfiGAoPTHGx21UgB8DZen
tjFbYCoQmTpkzIDCKrzllZwjQIQz4s/odz3xT9ev+U5ja3/x+13kEHSe2uw5P0YFwjMZDIxlVs5q
zcA2MabwMQXA1UZHV+u0Y/VyAjmp11XuNphcESxxTeWq4sUhPglD0cTEOnuWRSJSmGXb6yYmOjhA
LuysbRBrpWEqKFH5ZnIgYL4dp/nl4cFryGHJ4VXy/WobrL1JQAHTeue+9R2w9VBf0KUyumP1ktSu
A4u6ZuYHcbMS99yYfWE27wcP62fxlKbbMkD8Y934YZd3GJZtzxBgHp4rAmS0GO1yu5i4ZfPsWeG6
UhMy/h51G2l+o61E+KJokGNA9qNJF4znIBRM7BqkKAgb609rhnOsArd1xRq0kS3y3F5ZKqH7L8Zn
ZLhsip/NZ8qyR+T2RlIyZUvjTCrHfS6zIrPzHd5S6q9phPtMALJiRsMsethY1D/5sF0+2Ksi5OZV
cVuGTBdJxXg/saqHSsg58kg7vE0J72oeJkvbO5GQggR7xYmmbY074MO8Q8qE7sqc70yazZhJhmi7
D/zJ4ZlUjnWDtXHuRETU3bse5x57IGGoBdB9V/WR2N74jnlNAkWzM9y1iO9/aKl9eCWbJHjD945u
44Mh3LmjljarC8/CXB4x177rVvIZae9mSkStr3Ldo437KeUxNcZ5L/0DHrscWTwuP0a+dsUIiAhH
YELoJDuEahbLujwDvv07huCKkpNWSabLqChHvksa+HrABCeGCEe2MM4ZwwFdxO1zlxoTrhLpD9xI
NafPg/rvXQAnAGvuf1IqwhjtIAKLQWG67yKZBqAghq8IQS4B0j80w5fsfhuxzYoWluIHKuFST4YC
YRwMcMBj5UWXpM+2zpgKL5qZaELr5Ak1FAlqwiRPEWPgwo90bX1kqm7fvUGwRhC0W/RZok77Szuv
IZT/aw1xXWbXL/p0IzVi20qSlKBQVBkuRNIdGWO/PakqTI92cQOv2aFZ8cX7863LelmQfOLtydAO
FX1XQSMUkH84T+SuCgolzvWXULdmjOmwtdeQA4056gj55sj3zXlVz5c4UiI5W5y5b15olOSHa5jd
uF5acAQcd7oWSD6MrZxuDuKDKZliH+Zvagp74OzuvmKeiDxk5CPSIScxZ4To6Kl5IgVz2y+PjEaq
ZeQa21esyQmEKED8IPTPjBJMe1KWT5gFVEz+It0248mAPq44TLXYDju7g5RzsckbGb334DVWfv50
FS91oMyzuIlf72RyAGZ1hjRv3YSEMuG/2QPckC8HvyDf51YYYBWp11jvajSKmpw9L/b6c9OEE0q+
g/LBNoOAX1FCYd1+7EXth/4AUWdmXD1bJEc/rkHQdAoquW/WGuaDyjmtxUpFB5A9wrMj0vCFb5cf
GKZdE7Y+vYpPVbeQImmDu86O6kCDKqGqKjm6nxmTA+cnJf9jmquEAaqvOt1hJbSXMIgxe7/tc9ZT
IGuPCuXbIXeAPq/8qqltA2DzU63ZwwB+uxh9hjTLqGm7AkQWiyMjl6uBPHRa/UklR1rNT5qFGH58
JIFEfunquUfq0h6eiLLybieDf494iiErFv2f2jKtuC1YUWOhf3jtNzX3L5NShkAvlSYPAQcsIhx4
KGKYwSTbWwGkQ4/j6RlpuEF4Ltg7FSuY7dWw540kKm9wWEek/Fk+9N93n4ol6dFj2o/vbaMWypyl
Wb6JWZOYlJurb/3gomwTynz4pmBS+AFbkAwMGN8rhiV+Cd6WbfS/R+zsjdYUD6YwpxOXPtAVqNEJ
5MLZPXG3BzN9Z5OzAdd16qawEM3vv4GLfY5jSdecqANne1yddJ3rxIkJvy0ijicRRbU7K9sGnE7Q
wJ9zSANvvbxvK5kBN9kNlHQiDhdINsqlj+o8FUZEzPrw9wFhnI3LTEyAYgsCOrrOGInSbjS41QlQ
bFWvglt59ZeEOB2mt9Jkqds7oJxMg+CK2Kx7Dcex+uhsqEhtaT7jCw60a24jZFxOtawiWfc3Zck3
Vd6rsU8w42mLFvGs6HWhEsNLztfFa2fWC25+gjw2CFUn7yW0bnmVrfBBZD+AXQlOfuGlS89iJynt
EI5lPfm/EA+tk3mgz6rCeQzjBOff2Oi8KTuH467RZldn55sIrjXc9dhDmv9w6VzDTGLXOp4O1HYQ
Ry+SQqcWrTlmjpT5ECvqOn/hKl3WaAj9azBSrEYtxAsktbGrmr+/tccoO6IjlCHzptTbbfH+GitV
omW7M0wp1JzoL+zNwKwA8B41Y4+HPChd3CQREpJv5sfoKe7dFtRthLnP7esbgVAmy4DxokDc69TI
BBFJJpZ2u4ycFPWQCWeL7UdhZOk/dHSHFysShweP0Q9ZvyglKBuQeaHER3mnLw9wNqrTkqsaHHOw
+DGEYXQTahVoWRHtbQGo9yakBI1O/+rW3WLnAVvCxvKV+7z65a9yJpscsFJ49cKuEnx13Ep6QTm1
zZjFgImFNFel2fPlBmCfrFRV53J0KBIiWcOR6D2iKJDH9mUFJ6DU7ZSKUiNg+96Wal1LhBxMz8dc
LcIyPE3nubLQ2UYvJpD3rKNaBci7+0YXhmgXeMl5VGtrMtF0jE1e+sYzsJzHsQuoKF5b+ktnsXhe
4I7ucJhasxYnsqwn8w9gjOL7IiJyouOgBiiYEgEJCEfXMrmuC7ogkGi4CZerzDjQsIAiEpNl7BYV
zbSIrrMQpIvsnVtLPGbC2X/QqrUjgDchOTUleWtn5hgKsO59isX6hkj9U8Y6Rgys9UOYeIbKNTSS
atBLaP38P8ih8q/EVA/EU9tqlwaZyA4gBwZ7qumQKNLQuBoGDyJYUAmCcLxn2BSubfO327f4XrQG
wHVYq/MFPWNqvb4GsYABrvbboHOCTYoO4HrjKtk4Zk9mheZLqK3cE+CYVOpm4iI4XR9QuHfHQ0XS
jZLDTses89kZ3DfvwbKvamrBMMJhDIkD09GVONYPQeoq+M/kHdmzljJKliEMSA1n7sWvGNPAJrMt
9s49Mas+gSHPDhdtdJoj3RTEZ3TaL4D6YzG90ypRnbSafPGUL3U/yyi3IVMBki39SHboMUgvXCTV
V6wYgFzhhrgH8C+Z6jGltV44thjSNZurlnKz0vFTEluF8ZgLXoHtLoYR/SsiB1IQEz8Fl3k6C/E7
8Wb6y1Snpx0rgsgF4OypcXT3F7CPNtJXIpDuIfY/3eb0F51Rv1BEX/DB9W5wV9sJWS1+6ja7MdwY
4iVanm870lFPnI02OhVjtH8rhtfFWOs7HXcPu8n7h+8GUpkUyC5QY5CXAwr2mjs3XXxY/1TmwKlD
ASKPnTInmF7IK8RrBazowwgF1NJ8sLSwEeUGsBsjYspJa7aoEc7RIfBZUrxafHtADHOSlJIPG9ey
2ljQ4l9jEQ/2AaUWA4+HIYfitc1yLxCx6EX/rnNynygclCh3LAF7Mmbomi3gXgJOwn2JKv2ChwXI
UAyVi/2bz4F81Tk5mazR68VfQlERKRa6nFnkt7nS36pIFM3QNwzA3gBmh3UQ1QZ8jbP+fHDCpl5y
mK5p4FmjKEI4SLhqfZDWCP/E8ShNWOfPyWrNdEOYHOViIoLql94SKp4cvx021vIbEv73l1cpdjrL
pNwe78nBKwgWoX2UQJLIc1PM6qjH0c8FfjutsRlvEJONNZWiNIzM4BscuT0DTGTZAsCd+ir9a3ek
jr+by2kKjEAfxN2/8epQyMDAihDyoBZL40l0gLM5r4w0rDgwGgRPnxHp7AuWOFDOgngvy/Obo1qq
o6ynW0UhB2UqkgOee5bauvX6LNRajhvmwTjxqDnbvdrdh8vDVGONCGK1CSMF1FCMTCVgmRu24VTp
JAghRS1WYBl2WJAwOxuz5Y7xdx2yVVXuaODIq/axQRTpdgLW3fgX/C0BJwzXNMKDUgeSxRiYiPyk
uUHVkyXL2eM9BIbc+Ka4qfuyW1c4OBsaY/jxdFuJScAfi4bZsxD9t81ps4YGVeIaNIoXymbjKYz3
H7TqQaRtaahxDrlToqApCjWapIYSIr3cLJ6MOglQRgEjZtxNkytBhYQA16dTl+vkF2jZj1qXWoQi
dCvVNmTyy36jH+wb37FR+sRhemu36mdda2HdeOPLDv4n0ptbKJnQwDNumkagKlxb0YhRvDAqADun
1NQXfpghmtgVLDxt/65rfo75vOFRevniNqQGwHXcgeIZzi3oFpIMU/hhUFpqoYbjFuPEsRnym8EV
vS8ziYhrSMTUWLEcdK4oCDA6dfofzi0aDNKxB3alxJbUCcvjGZCigh5Q2J4xt6z50DP+l815HzG+
LdG2tDk4xmnhny5QD7NtPW1M4eQFcswEK0oVw+TZ5ZvptOkml9Ei6UZt24okHMBSc/mfcZQtJQk5
TW0Pn5W9MJ41cumBDG/huPTbgl2d08zL6iTQLQ1u+rpZvDgwjrtdxKCaxq9LmaSnLzDRf1qDFGN8
Uv55Zo+C3ITLobbeT73kEQyxAhn609dqt/VmLRdc49XmydQhnMz9dwbWjbLDAMwjqvO7mCXTstXP
7vl0P4uJ4dZroXMgMS6EcMGH4oy0qvYBCkxI1LZOgO7JLZgME0bHQ+MjyqcCpBjjEH1gKYiEhChG
p1UpRtfsOU5MwTJMNRqz5BhWxAohJfLlby6vGNKFrflyUi/HDG9I25LnGBvr6RUIAgtXQd3B8BTi
0Ghk4JgxfOYwSssiKrlHcjT0hPcRgltoHh3cxY1ebDoIjUkSfxlYaQr58v3kGvRrqBvXHYkMyseS
psPWi+4raABf8uFg7RhYyzBk7dCULWu294K8Rpc0NoILN8TLBlRzbbvfGi1angrr4RAm7jP08XoY
3NaBLbiueSyweOwrZ/QsWYBv3Ph1WS0HU3QjrgnfLZeuvnQ95OdG6LMLTi0E6N6tb/AMZN8z6exT
3QWMAnAKUf1o2BUspcMLh0GSPDDqITM0KqqtUYWxbz1J5lGkg4lhgDAHvpgza5ufpyV6A/C3FgnF
ObDmNA4h31ybvWBFAwO+X7y7qIIr0novsR4o8P7LL2QQqiSm2enFTj+I3J2b4F1uPDSP1ZjsEqRZ
sxSuaOAzGosRx85i0fi32OynT/d/w1wVAm5F4AGQwhin6edpGR0QOE27NDaPXmJjs6x0Lct21Jdv
JAkvbxZFpQcZy5yvc1hQmPYtJgA3QuGEOHqPGFpHfq5KiWxu86UgeRZ3aubv6mxRbPa8QM6eTd5L
LlOJtRl1lj1nozVz6Z6gRyfoW/QLA+fkxendL0ofH9rn6lAv7n3B79nQfhOusQ5tJU/lTH2GJ+1y
emc3VPsRqSnWxoEkCkd1pSyolpl1FTRgqJzXmAMGhOJfIdGg4FZI2isSQfQQ41xVNMjp/xKCKc1F
IRWhfFbpTrUr7rrpUW9EfBQAoD3TepmARj33bxdiYDHpDK1jwNSDucStDdFnRyRBh8QjpKyJ8LbK
cGmrQBCjVOSNAr/X6SxPAEqV/xTnN6PLZG/gxvTNQiKp3Snn+E7DfI4JvxoFnUrsG9y2CiWIYZpU
opIZyHEAqwDzaEVSY+UxCwXh0F25AY5buU9PhnB0kwWKn7o9fUC0cB5ErmGgJqgFdhAB91IiwQpt
wgI/bLY/ZMM9Wcah0kpU0sAjqKnmxpWMhOzhKgjzp3DqbMtYT365GIo5eEc1zuFUJrJ9EWmbcCXb
5LzTyamTJnXtSmC7mYmEmWaSOAa2dE97TPhZRR/JVnmNOO7wT5UKXUiMRxrOcLi2DAV1iSN2RZNm
x8/PNXWL3qjPlW4JUGxyX/mg4U9TRxE376A3rT6z5DTysRyyXMB9v4Z/KlkcuV7NFYrp5PvpgrOo
v0xT8xFU18SMzMsulfBDKCjOdReNsYzMOtctH9Smm02sG5+QwcwCRHCuzYhUYMJtacLN+TflFHld
WBBXUyuPrcikPnaryGgIt5I98KwXf+eWKYt5+AcLfy8VlkxQiZlGO7rPjEWi4gtwcY0Hf0S9L9pu
IK6T3qOet/TAmRgZP2uu4XnfSx8LGhndGF0HLOHhHcqdIWcCRTMFzgYW462aGVC+0mwgAOAL4kir
9/08rxhACVtT8K9r2vyAAXKZJTX9XUzmL08zbw2MV6BGhaQC8mPirON2raasCb20lydz4UUlzXV3
CPjwTl0gSJ1Hqy4vtDVNx6ROODXsLLWSHApkVJ3mRR5MIb9Oux+RmVDIeQORLkxJPGYpefb6WzF5
WKFgrD3fd49RcIjir7nmNyTc/Ometq08OCEj2mtvpEvOyRXJZ7XkIXagnNXkOharZboeiKZD7NEg
Ho7/J40xEqBz404WVgGt/CTOm7F6DboFwdtzqDREkcfU6IHF/+qbY+svYe1rb/lbzMExkKg0MXvv
OPDzFLXK1IIGbTPkVXb+SLncttQKNmpwJADz2rbJQmf59dyqUxKWuVb6VC8xPox4VF5wgUCRfyNb
byaggKXvXzu9WVY5kIGUJDfpKhhq0uzDokVaJcuDbcLLbUunRWGaiXiE8rjIVSMoouIP/zUuaXuE
EpTgk/Mz/EVPDfnltObXNIQzbumuL0HaG5bR0ftFVa539a3Yt8OMCevih5IPFnc8g8YiGmq5R1l0
bDVDbDCu0deS/hhmNUacNbH/5EGYPpG5MuUZgo+++DbehkU6DhVBkq2XdGlskj/l3nnYsgbs8B+Q
gTt+XPS224QpZ0eRGG6Jr6iCQYqRLnZMMXhk18Omga7BLRnV2EU6ZCtsOvFt4y6uSfljdlZUV2b9
GuknHWdekCCnvw39U0pXCfvxyz8WtoqKvcP6bYwIVc2RFFeBp2Fk1/uryMVIty1fzyUZt/FZ/XaW
s6hS44W3Jk/+JFicdnbOxN6ZlQBHGsvWs26a4gvTpHggLZnCy0HASZKTHSESFMyF1KjncJi3kqg6
NcckkTnmvujP0gdXnbpopc7RQYAqcfOyAzxvY+c7mvK6qBh6Sve27GfNbA5TI8+qtmKG2pSsZDPZ
UE6Qt24cTRrrRgEcdRKqx19b8EBKV2liEk7GRzIJsHn/LAoxiQubnCk9evS9GoseFOmyS4jVxqhT
Lo7tbTpPNTXxDwUUuaP+ytugfa/ZHv/a8Qp4Or7ZN9/xwxcjhSkTsFpKq0gWln26q51Ghqw9FpUj
LsaY4BjD5OYMoMe//0RMtMMZCs9VhFVF/Z9Pw04V+qFn4RX8N8L64PFWjv0+LuB4fJWnAqYfZyh+
2QQw+ZM6dA315vcxLYwva41jmO0NvW+TVCWgigv3bwTXnFqI4464DF6V5m0LUykglsSBIxZdUcAl
kYsz32ntOVK5kTEEFTrPuhY/zn7MC3TU6sFajmTkxMPFkJrV3E2r+JiXU4UmFRnD2yUteGGzUubg
VpgWGmB3uI94wsf5qNAIytYqpsnpGT7Dzd3ow075H0Wbtp2otsnYEhA+ZdpE74xKbcF82rWMGI4c
fumwYfWZFvQTQbyp8jN627R6EBTrREbjEaC11POlHBkMpCQCKGZm97U6x48zh3K3A+reo07wIuLV
2q9JAZnhFdHnQl2AA45qFuS4ZngYXf/uPzcfXrrKPqyiXWzYEhb/bNZbFduy9th7a5UTH37TVh+1
heBdsYSZ1TvMR4GE9styBNKZYmyMMaae2W8niPN3JH30MLBg/Tz+kN3xekY4+kx2nlN6hE+JmsBw
l2H5BYgp96OCp2b0XcBkk/AgBiHoUrIoQz8ZFvGF2P1U9hcBFIjlupw6w6j3XYEGR/7FI/34ZJlm
vsqBe80mDP+vumbn8AOKvcmXj5kAPmxTxgDtC46HNQ4ghBaqYKhzooPfuA0hNXNLiK9JLLkRYgLD
LU3VPQYd0SoF5YUMeNbN0MoYb1XCQ2iDj+FN6hXm1d4OVMwY4cMKUciKSmaaWClucnbeVY/BDZDy
6i5NF9PF0rFKG6yyMsWpOSGg0Z6YR8StD2AuXzm1oRETqPzJRFcfBZepJ8E4TMRaa5rLUlXlbIEO
Xwspd3lQGgXEO/VlAq4QeV5/36wpa+W1HX4LfbzcSgkJWe0O3l9MUfGERh/2g8XE6qUoNWXiFGIA
PpCufcP2wnA2QEUHaaRIiB7cwtibHiLF7+Vc2xXfAnku3OFkJ9OZHTrm6u6X+2TS/eiPhW4de6u4
pysst2zYwnR3aWXq6HfU1vSUSQiRSxLlUOBBiZ3keG9EKzq+myLEcKP69WYl7waVaVh3olZYBHKe
LvBd5XPkjyOE1HOVJE9Mq5CjpD3xKpG9KTMG3CLwmodcwSYKK/sKwGkvNq/XCT36ET5YmAhT8QrC
p89t8e2x6hxeHEMQ+RW0dEHtRyjI+JvKlta+UOUQnQUY/N52J8zWiRB5trqTbP9E5gYNhPbGZ0Q+
JVVOTXdDepHQ3yWCfPJam4rX6+vfi/A3qZVIEZxNVBckP03zsWe45+MIEr2TRsbpMhQRd8IgMu2f
Tjwj9VlY2iNXgQXn91YMA6fE8v3muEGIhnLkPd671uQlKCymVCi5ZpUg1GoscVOVk+cGtTb2sUYe
KyNWr7XwE3NdpKiya9XoLN9X+EOQGHoDPEps0/RpT3krRbLM4i/SFct24Ytj3dHzg6pFXL0cs92f
7mBry/7ZG73ptDzRTnmZpZE1FP1zP11c+HsYZq9utYZlHI2RgXzzxkMOEc2DITpkVHboHOvjykhV
2QdnfB2RPj+9txTqVUIAjiSE5kUTaf/1mBc97p2CuzKlPJ8cSHXxSrE7y9eX27QDMOFd4h2FjkvA
c+eMX5ABQr9EAdAXTCnjx4HwFoPd6gPLDBlBOuj8vXSTw+17d0aX0ILf8pC5wvgPjr+opMwuUYAe
fsyybnmu8D+E7jbYmXNASdUxU1oAPwsTcSnNod9lFc42fnFOwT5yB60VRn8RttG+aIoqhMaqambh
vTYRto8yuIYTY09RtEz6xuM8BflaNwSWE/OisJAL7sNcsM9zDVZkpHAuCpBbl7/fvn3y1l4YXVTw
AaFikTXrbh+2oybuft8o59wkzrPMUJQFDf+4XDk2pDCXKv4V6wdl152PJuwnR2dybHRCr7yveFlo
Iw2BBEuLbO65XvUklXNerSwF8RT5FvA0hQFK2qzMxAxjJ3xidXHaAyMvgLrSelCoVRP2gFUqFiXu
ykssR5ZXDHiKDdCSLnKPqyxFVpB3aqegpmZxvhFmYhQgmZISK2vD32PQJ2cfx6vR4yColPehmXzR
onZSpwJye9g9WgLsRlQ8dYa1ztmhsYcU79iK+fmjcLhzLstskArb92DWnBeW9vF5L0BdlGfQGN3p
4T4gue9e97dsjqBEugoQXyMyTIqqUHVNGYjJsYK768MKdugkIvDNgBgKv2OpNIvDex2pAZM3puqR
foTSnePviu2UFkcPKA2ZeGPQr8Z1YQ1jKXbULoar0JjS6p+EsCA+0lOLf/PdOaAAGEIsvd8hyQZK
1rgwafyvbAb1LGNTpGtQWkDtXYWHFZ67dpFNy6/QxZajWGeeqA/1/ELldZpXZcrFzWBE7vDxMxrq
y7ogFQyQTx26jzWjH/AHp1k7khlcFvqDFsgViIKTmyhPgdKduaqSGpWnkxRk4k2jM5wLyNGF2xYu
lpNoofJQKImIjdu0AXpyOvqlykUgidOrYduvAH8ztM2T14LEQlqvInXWero4jow5adY/4/Mpy09I
JvYEJibyhaG/txlcXyOZiHhPPIJXeOQacBdy/BuKux7mazk09fjl9ptZkcrw/PpAnQdtbwMKVGBf
0ZXvFtSFXV6EPWP45tRsCKTVV+yb4Cgf7Nto3jIVd/47Ifl51ruxKQf/DVHDvgrtgx1iQxTDJtp+
kynWNT1YZc+23pABADBFD6SqpSWcOvWD5lKRo+80BRFM22RP9kh0hdNWbQk/pwAZWOG+MwBZKDZr
VeDvxfZjjHuYoLR4rxDI8QKiqPdO+X9VkvhulHW7nxdMlqZ9nNxdutBef6AOS5ORjl6jgk75Yg6S
eE60dLFAWB+ZaRrU9DC3iENH9XchIrl5aDVhE7NQXvndb9V6YU59w66MF+zSrIc9pvtFbUJ+qoxL
MsKd97MU055r8QkD52WZyP/Q2H2cErxXN77ubjf1T9j/NnMaoaOwd+zz8x1uWPFE+x46rd/3l3uq
hLSr76hz/7S8bJGGtHZmRtRVpyyMOtiOJ2ZV1JahoY25wX6NppVPTxw7A95edNwczWYH0bMzAMWS
HUkc/xO5O+CyxzWU8KRJhEFTe6pB0Rn2o9AYPAeE3TpCnfTzEeXDIDlVKCcKZEpt4xfh6ovqkjJX
osWL6tVWYcUXfqh5D/8YnQ+OmUpFlbzdL6eekBeJD+WB1F/MNzIqvlquXDCXzDnJmczYy7R5t6VL
WaqGaa1hpx+at0mxxfYnP+bTu1KkQmnqTYHOubRSr7WlaGpavhng8/VhupNj5lDsPUELKr/KLMOn
0EoHneR2smDJsiGl9dtMoovYS+rBlZ0RnyTvSRBCJbmvYShCyR/tIQ+OdaTeu+rTqzaWAQodp5Dp
kUR0zrz0Vjky+GtDZSmEawYLq87OhugaG9f7baszPheMzE2cUBKlYx9DIWpl2kDakaLZpD6qPDtM
IiA/ZIrsr2gYbCTkv6wKs6j2ebMQkOewU616VGlFZMCG4mzBYzqxc6AnpUNkDv9jaOWcIHbVTqc3
Mgrgi0nhc57gZimxlfGA/5uSNu1vwNEnuyWGsQw0RHa24XLTwN3rrrMcfPmVuWXEMsLk6+Peqaqp
J+SNf7z78rqW/J2GUUCPrV+JcCY4Xf/9EBARiIiFtOndzoHBmiDtPub96we5eAh9moRIsvRAuEEO
/uHeAUGjSfPzmvy8VIuSAOsjFsNswsIE9+LIXzyqf4l2nCerY8qf77yoN5hDBmcgxW/QRaez/PY8
VI4ROuGh+t1KQNSZDzumCPSTOn9DkQskRis0WABW8q8vn9o7++u7AuTVRHgKTKrF01u1cjhGbkuo
2w2lNa1sH4MbF3SY9xv1tfvPFMp51afbAMVnUSLyCjgrWK0l6xEzzS8atLjX8RMMoPoM7M+8NPkS
9eUCtakO8UhxKYiB83sApVFwMWAvHHpw/AnSyVCmmlO5hcy9bwAj2Re4BkZRZRTCc0KlkZVGYYys
rbYGUAf/BV3M9r7BvXlReATlV9VpknKGfmo9JI1ENRo4Qsm8IFGc/b7N8uEawqpABO/ZqS35oaic
1zV6GrPiikXPuks3exlHrcwrDklmqelLvgX9ml42Y59oR2ztNfbe9+h5FrwOlu2aJD/XPRP1XGIA
vMbW+drepn9H0SJyw+b6qR5EG02lYuwl+aECiLNP8DSMH6gMRIaayzSUraWKw0Ii3vOkBAPvG/9B
JvIYmLZbG4kunkPOAOIg3sgjU7mOZAub+ND0LYMmMdNfwdFO6gyv1Fbyy9avpMe7jRZKY+9VtFRT
Dn6jTWmaHXqAoL90D+Amsfhp2Fw3l/3JKNbfsUfZCkLFWt+MNJPs1dh02/4qqdk+4HjoFvP1C50f
rtZIhXDFsmSeWiUs91Svr/C3DI+INgivTcy0eJi5ibaU83hsdFbzilcN2F+Ldf3cb+2ppbyIPjTI
w2w4as5RHMaaIs2FpTipNOSr+F53WgR3Qpg1h3p+FoAmaWHvsy+2uWYW2uQtbWAL6+hR3f2MABlZ
KLmnw0SicqRZNjeLVnKZozN5kH4b9OWQ8AUMcKAyCg/kS1a2xoWF1zQYgA5Z5Fda+MqFZzw869iQ
iIhr7UOaOMYqeUSOGftHbIoJf3rKO1vDuQ6Y2vJrMJDcprlbPgvOFWsB/9Pcj5mhUgFAd+QKa2D1
WQB7+4vqp3Nxtkdk/9oSkVpHpB14ZfJebVRaoiHxxpQ94LToLDTNZ6wJzsSR2mLnDVxqcBAOyB+w
q5B8mWAgc8I7iie3Jck/xmVm60AG139ca3NbpSsYFYXRifePXa6pvHmUqLKCkqy3y8sNRjpdQgfL
hoiWqOJQ/IzIsEunpCL51dn16yXvYlcI2kcEshrn6j5f2uxPwtQh+ghqMv1jzjkGlVFopUdkIZcd
ORMjWhKrkHHt23/AtdhQAntrKBLMvfUOdm1+TfTURAyX3uea4bbqYx0U631W5Uy1X3bQhYB5/2z/
asmaE8LR6bfyaFT5/DfoukBv/2p4gBiasR+KQqBkAgJHhCiVLHlIjHwq43FLwt66hTSFTSS/15CB
9Smy5DOgpolnY7kc6AhxZwJXaRrTxOdhKtj7OxdFY8DaZj4FyDJahWnXk/oO4RpEfjrhN69Pkqwv
he+qyxKdaPC1jqNRD5MKFpwFGmyqSr0pKhkC8kxdh+7VDAjgv//jKjiZUOsUZRhtGsR2ETArE6Bu
rrYa60copoMhRW85udzBygiqzYgJI2jYiLqcy0OjWhrB605Kjr66ijeWbEHABRPxzMxzg/fkI4a4
/VUN94KhRTYzQNZxWd0jKzQpAXZlBuTn6dVWjPw3kY7xy49KZjoHH0ig6rTtBhn1ARL0iHCC6CHp
X6z4AinGSzjcD0nKvfvxV0fQHgMhjAfFZ212N8gANceesdt3h1wbPZ+YrdnoGa8raVdt+NPOLdUK
QyrSMUILD0HWyMf3a2e32XC49HF9vcmuJW0cU6CG05Je6fKkPNfs5/ky3v6NfDpCG5PI2xa+07Nr
wP+FX8CuBQma/w6E38Dr9Pv/WP7EqyOUjEzR9ule8H00dvgVJk9HceCIftFMMEVWlo/icRcvSJEL
L1D4XOHSxYGEGBVmEeD7e0E7SXyz+MqMvO2TNoXj2pMfG0dzCvDHtgMVLE+14jlqxRFp6Cpn3V6E
9qIEHNGUjHSHPZWR3C818Q7ePqLyksBGrav9flMvx9aVEBF2uZHHmrnxj+TOjk8FdW6KGl0fOx3+
j1BAN6qHTsNWnW9WAUq4FZrUyBGtOj5i7rETKcDY14zxfbpW598Mtaf1uiYgsdrsYjxf/y2Yl21t
n9CFAYcULxuoHrhnP6ngZ4SKjdPueu0fic77Iw8yGmjTNDpHKimskEUmpLYWXjY7Q2F6Qe+40VbZ
2LTDnu8nG9ltS0LU/lRXNELaOtUatusoydwqZaxfb0VTRcpZBjWe1DTBDiiaLW375BiFw9NCAkWo
bZqkAPmcaAVX9WhwB5fPSxruULKJQ3jUdgRbcWKkO9rW5gO9rBnDgnUFXqMYwVnnXyNan1tTPaUD
lmPnIeGoy/PF/z+iViVQSbL0trlBTpZiGFIDBmfeaNZJXi1TKm6/ko9mft0QwRuzcYaM25yEKS9e
afR41c81m89cMOwPoesSP6IPxW4EFtr7jplhwC+/jXWVLvxCiVpMvAqh72cE3Vs5q16rRENHj4cz
9bYiC7y+GqculdJyPLk9oghe3G7mAKI2zZhLOisV3f/8JgBtXfMB+BBfz/8HkMARYMvlkZoN5Tcw
QHMdABv3m6h53CvqMjoQOK9h0U08tEGI+UDw5SE5yD0zuQO9WPDC+yvrceR5iEoqNd371Dt4Rfpk
WsJQoSTUksjK6J29S3jyqGk3oj+Kldff2pVTbJ46gCGDNCIWqxRz3byGOsY/JS/m81xricGXTQrS
413rH+8OD3y2ni/2/Zr3aS25tkbq1+8BdPrHUqOyIbji/CIJ0V6fhcYxfjP+XoIF2b0Ck0ZLf9NI
eSo7t60ROXZbZc3g4iQ2r5Mgzo4U1Knu1wcO3jF8riJF6NI0AV9BmvJxm6D2yIfDmPxEZUgOqIdo
rzIeqAQQG3PXu5WM9LjO3l44JqdpKNoc7/R0E5WbtYRj7mQyflvMzohVqLREDYa61zgCkR+E7cSC
hWVkmNZ3IRbqtaGz1n7ku0R3a6dy5lSUmYImUJP65/jZLjdUj4moT5wIpZT0+wi85jzc0rh1u9GY
6DGtKjf9xpM6pdEMdyqQ+GGdxdeCf8lxZWARjt5rMQjLSiVGZQlUJAZOs50GIxqyPqEiuFFSu0vp
eb00T8ZGNEDHs8YsifxCDhDW3fbj0wMi0LJhUqflRDoeHB9iCztaE+4mDq+5sy9vR75lxgnVjNzw
NU9o9QMx2dliDs8APxWq57lSjqmUjH7a1KYERKStRbhz8dvGea2oZs5+x1S364saZ5Ls3Z5hzeQI
FhSfhoB/hyPEfubF+jmJM4tZJ0Y8U09jdVmtEkygwQ5CzXF/C+8Wva3x7cxIWnj/yx995I9U6XHc
gX/byVBDjnyHFS83Q50LU2I65Jr3jTR1ghasTfMvitMoNT9IOhefKOs7FUTSyioRxQQKH+ghfClE
/D4l8Rx5vHiUCJPXIrwbQ5kPN9wHLHKxi4aIwpbxtvHRqIh+R4ZrMkptJjqxc5G4Gq/vvH4pyFNo
Dfn22tlEXlq4UUVvExFfjWBIS+wB8gPcHs6YuqB5dPGpi3HPvD3IKN7WrWaGLNSVKl56boqB3XkP
dh/+cV3vnkF+2b4IG4Z/oFG/FjRh6053dEVyxXXeNrWCMcMg9NtvmMJD8YURcWWIC1bPwkzpRZFr
IwHNfW7DJolpDEwusX6I4phdJPmrElFfvkuy6hItowNyutwAs7jdD3WhRuY1j6e9KvsYG+YUtPCO
e3YUrQ55moegxkqLniTs25akz6fpWOCZaoqC2cnAmm5dbBTL2ZOj8DDV/j0jZf6dqvYt/yTGxZ0T
z0Z57/9nNLZwWXAZ7p0D2pz6df+P+qnDmHZF6z/25d6oc2oVACTtJDNCluYXXUwTN2ArzlTnluG2
hWGUsLQS3D5ZvTTNymZ3xdWRnV2SRlq1aQe799FyQeWhuxVH+qjXEdHi5fXy0pHik+P0S4O76wLw
iRh5H1RvBkGK3+hkuhGnzLpyKJPrGcspCtMl7JY0tZtDS1l3NKaKT4zmm6l59sb6wD6dj6jWjeUh
TKEZJgkkfM0aOTyGpiP4iz486+SFHVXCJxTfV4WaI6QDVg25O9Mxx7Fp+ID2RSHLxdo3KCR9Z78p
sg2hX+zNmfIMD2u+VtFaEhbjSLWntfHDmq/jxkFdKwhTi+JiYx488Vmt0GaCuanDKGuugq3Ldl0Y
eT6WwHUIOSmS9a+zizojb6JQunoJfc7TEZN/ZobwAiB4HgGxfeD1V+m7BL42SIthdVGS3a7tBi8Q
g7c+VFrmPbwySE2s16r8pCoj5uqX1Cqo5Ov/GfAbQDIMti0aKci4X8uBKCfPLSxRD6dAAf4fRkcJ
0J3JNWKUcdkdSYZDuU4+fQSwqmYCjinjGzU2qLxfzLRf5WvcKVS/IMD2Ev6YBwKMoEBJSGmlofHM
2Ap73t8r2Nd+++jzVyo8/iIR+rA8i26t6Inkcb4p1XTa4A+HjHtAa4xwVIizAzFQBDblLgea7xBz
XXWBuRzj8mGUhMFPyvZUWiZETQGk8uSUEhvIBUZl2A1KlK1MIWJ2T0ZaJfaBGtzjia75mZpT6l50
7gObiv3XVlgu93zpvyp42uNar8D7Fqj0ceAxshfo5EDUr/GjeszQpMirUL72zFfPGYM0hCJaqEay
2o9eSkOVTPRVP6RP7JC4zMqxzPG75jhEqUq322WHS3yhSiusM3otDwchIc4cwUJTcOeP+PbL4UtZ
Ant8QgYSTNFjkIZXjGesZYWZlku6BWxA6sHoi8ZxWVSeGZNm/csRW4QlRe2ztXDyDJI/Fuz9A85G
TY+DM3hx4uPSI+ovROyRGi6wB3xYShlIy4HnMFgEWRlpsip672LBZ6xY7xS7RlSaYLku0ON7NaTQ
jzRCro0QifIXDQXJRM83xbYiOY5T92yByIBunaikUnMYiry3fBUQ+cSx/R9RUIksKpZypgK//Wz6
KWGy96gK826bPB2vBv4KX2B4SC/Ssp9MmqZA13Nlj3/qcErysCITvEAGKOcirIStVHeZtrIhF2L6
8zWOKuZ6mfnKdsMdmGdKyLmwY1a6oftQ2osxpWTys4slx19z1IZuoS2OgK6K/ZQ+km1Cr7xkVDP2
xFLxCFkQ52GGPi6mUBa6eWJ6AxuZyPpv9LFZKjLjSh1TepqxNkcF/YMHvIbnkFycCYRdXYlnKYUe
QtagFb27cQNfWilzBULDgOumwpV7Z4LaVEe+CglDrdeehcU+VOzg17lN4rSio67bhJjiycOaj6K7
SMy/hkvirbSL2sp8pbdfqQNVrkYovCucbcIfQCTtl3zMs16LzjSkoaNwrd8MJTvnC2cZbmvzLeqS
tTEESziXJq7K5plYmxS+SvkbB9Mb5Ge9wpesxfa+78hh+soxku6oxUcd6/wLFtDGhBloNwwsL2Yc
L0IMLgc8IQDEG4SwikRqT9IkmDrMiKG8FS4z9QHIKnkVCxmIF5BvN7KJDuv0hg73nneNaOcUM+tC
I84lTVZE2yP6UiVJE4NNs3uinAnA73kMgBhJpLisgB+0hyZpB1sKX1GHu4ds/gRUsqXduhuAm5nZ
W0yhf5coEvTy02X2kwpwo3rNoyk+dOSP9OF1Enbbe84fd3yO/wE+t2M3XPCuOmAFX3KFg4bGmDtB
FqhJF/mNLlTtVEwVNYDKSL1SBSNu+uijHc8iU6FiRh0soCdW1Ye83T/lFGXEqqZQoaSmEguORx6k
7qZIg2I+icqFv8vxZZ/+OrrTyvcSxhDwuVhyQznkq7hdzE5ht9ogV2uf1P0JI8Df80D5z26mRwrp
BTVDH7+B8FlniSb07PMz9qPVbtgfwFsDkgNTPeOxCdOyi+NJFmzviPV7AEqI2KUkyioYt4maK6WA
x+hVNRIXHXg14zpGKC0dN4bJMcGyi56IWevCgKB88kun2g5SGF81lTKO2k4I2/FkSrBBjR8NsnZ2
hkYhbxqg3i61vwrH7h8w+W2as9D+mgmzRiB4OD5awTAnL1jC7i8g3YiG1du+/YfX+CJ8vKV0dMDa
//Cf6G+eA0EYpHnaqCTopD7xDM6huEUe3vNVAS6rgU5ejL4W6IXpBAFqUwR2nMwz8ZQRQ/DicnKC
FSCWxkQRt/xo3IEXusqA9aYw9HERr2FXe0BdaMNlFdSXb/bAf+Fk7oRWrYY52ZW0mOOd1alhMgTZ
9YVIiC+Sey4y/zU6qV/jh9c0I1sSHLi3pv9bknRfzafWrelhtFo9zLa1XnWjsZf0kCGxaJS2eO9v
N7lCgZwJcs50R8wAg5GIqV/rKBqxcHG5GPRrXUVQwUgb2FseSMNWu2Xc+LVe7FElcd2zIoMcRpKI
WCo/nK5RkadXQceBe2TFZr7lhj5xK527OsLq1w2TQ00dBtQrrc46aZ0EcUn13HRz4jC+JTY8djr1
hB3Uw9Qa8ShO/sAYd9ydIzhztFBktBrSa9qt6ppCHCjVIZpaeVUGplQGJ7+alg2vLfViyWS2v9k/
HzoEC5pwPpD95RClxewHUV9qNxH0s9gGPTdg0Qbcrbjfknt7cXXb1CcIENc0VnvJr66hm0j7GI79
Yik5oC4B9LYVIRf16e/h22AGhv6vBZcAAv+Rdp2jGLM7zFpsuvtXyqGthCdM/iQAoIsGHR9Dws+5
tq8IOPcMtnYReYdRLGPAC5yjMPVe/zviBw8l5MTzDJ0JEihbUOQpHHRCiwAOTu5CWRAr/U4L9yEx
/4ypod1g6k/GGrLOCG8ysm5JZy3OmC1tq7Q8V9yMVF//n/MTbSO0znj2t06vuBA+6IbF82NGZiKZ
hthHlwhvHuAvs/p2xsZmv/8AHnqbAk8ytAE9ih2is4xLJwheXip5YtOYK+2JfbAA8UxKleNKubYX
4jBixYQeypSj8KIG39cezD34mZyOH1CFBnk6O6g+20mXZ4oXMHhdZBqVzFw5rjuLeku4M4qXOkKa
uannBMYOSKtaz6GuFe/2WhRaYW5DDJ1vmpMhRRkK8J0lWS14OGfIKOrZx2ZjM9U1+yi04MHXmwsJ
eNSIw8mt0DeKILmAlkmKAwKiJnX0n60IQ7Nowq4D0tshOo+KPq107ktBQeDNL+9JR0FgwKrO5Gms
TEFipuE8QaUScNIoA3VKP2lYCv4WueJBoxdTCqxAqgd6vS3Y1H76PHT5gXgELFDqwKL9usFdeOmN
uT/Q3NJ/c1w3F5CWcOzIuo+tvje9t2GvwSbwjH1tY/h5uEXgRGYx7WLdoWhhMtRvE+n8fXssk8Vu
U+U+x2xg67xIcGT3t3Jz/jR5WjbguDk2pKKe7abawvWFQtcR52MVXJlyfyY/Nk0Gs0qzZo2OFi6Q
Vlgybn1DEB4L5ZAqdbxvMHizoJnz9e9G7utg6GdMmMOh6YnRnOsUDIo0flKRNgfhR1vJqsd5wCa+
WlyhoxtVITbMwuR4ZbjuwGfkYT+bMzs9tEAEDwz3shDVwzH8Bb63gQRoIzwZ3hakPsolE9s3/P/G
03cRn4/qVyMDQOkYYoc5ifmv8g/rkBdDwzKLF+B/UytrU9k+mUu5cNg8HTA5z75uarwWSmoGBJaV
F/GA9dvPP5Lfghe+xcTAlvdBkWy7bPA8vjTDdbsOJH0iX8yU79KRz2sroSF8cweC9I+GBmjsjSvj
h6bCTvjXs7OG4j0sJxB6Ww3XF/G5jbqEnNNeihXy418hYZDfg4xdCiP/h0XKBmsJET5PBQi3MtVp
5iARkKQFANbuud6Y0MPNeclulDo7ctGSwoKHR3iie0mFfBtJCM25RhnRJy2jqENOUp+hIU5N1FFQ
hjOwSFl6YTbWK7wGbRuJYRyFyWfZgeDKu2yTcHFN1JU0tj75pGywjAG1w0ySISQHNsjIJMH/4qTF
olj5kFpM9h11EQD7lLZZ/9mEhZnX5BdQRgRNPcUZuiuwANovtc2CJfthER2NXasRbKaL
`protect end_protected
