`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25696)
`protect data_block
Xu64JJo/wm2IhbNWqyGVvlzheLSJcNBea04Tr093226ozyhttdx2WEvw4rJtAEx8936UqWlGwQeB
qRZ/OUiZm+0mFDF5RWU7G5r7AtcJwrjFscmXKOBJ//tD8GeFseax2vM9PsqjJckhdcpJVSn7CrdN
Hk3BW367NbkgenjSGVqRvfpCrzLo3tRRp/qt5WAbgy8l5BmdVuQr6hd8GyQ6vn/tsNXrt7INSOFb
7WL5yu1Tv9wt5Wqz0zjpgiN0qR4N2sWO04GD6dRstQvy5xECX2gMnsBNiYYQyo8G8zx5EfiXqUi8
jT2841j/zp4EJkvCrdmtTQrSLrrY2OL10FkS5KmnSMDIv6WQ+vhc92CVZC4eAzx7UMf2lF8O41l0
9W5UpR/aNc5jitSPoKwQAzkN7H3oI2e2svkNWDlTE9RDsPn5lEnkYRyZEvcIWJgdS+PuKFxnun+e
lmaD3XmgrtX4wTE3DIzTXsnoRcroUhjVOUO7cuHmzPg13o3nF88Cd4t868jhFFOKNFmv8810D7aV
/v+dL5la9Eodjn3SGXZPNm9min8sQFmKlU5K9lmNFM6St44iBQ0GHg8jTT1ekVzblm4HLebHVo2H
K7xL0L7cR2TRQubnhSAOcOVyrbgMoazCdnU+GYo4F61eMUcMmv4kQjYfN6Qcqqv3XLD7xEgbQaZ5
eYVONyZuETmkQptVBmD6me5MHEgjMPE96FjZ2EHOoucMBiYDn7VE5GImDs3pgFd2tyAsGa8/E2On
IrwPwZUl8lHeKA8Im4MGmbCugbPaai8XWaVzqrU1E17PBU9c2QtYQW/+/uiyn1SfMmYYFLy37OAX
+e6ErNo2zhqK8xQrG4QADQFlUvgJ/w7+mUl11QBhnVxmbAAb4lsfVMgMzYYdD4o9RcI0gXf2ixTu
Qne9G6ChUN8N3EE+zr/z8e9KtkbVavELRXiUh0Qd8Wjq86VEYQia7/O/DY+Tz6Lbqr7WJof2zw5n
Lk/zqJPtUQXZSLu81O/RQeUJLhmaZ/5x/C77NUAo580FzUmogFPsKzF1trRAs1hL2SF9g/Y3gUC8
Un81G4rwER9lK5SdnSCN1rKhhgvN6QXth1nGe5LJhKVEkq0hg0rhYWX/jyzDYSp+l32Q2JxX75Lu
HgInwDWl0A6dCxAInIqZ3730iSBfnQS7PCoPcgQjx9qYdRHVmXAtv+86uRYI8ZMDdLbT5YcZZRUh
rJXtuR6AiSmuThl2R6EE8fK6W3iqIttd/gJ1KHncNcU2xJZVPx/yPAx1Xgi6ReAvAjQWBLGXkw7Z
aH9HgOnx1wztla+0VRrNTolCiU4Ez6CLqrGHP4s1WeBhNHoSRvyIM9/0gzxCXX91WE+0c6bEYlvn
IeN8TgsZbHBcNhlnhVVcLzHeZ5Myve/CMhdtvrCjj6U5KVvoVSt5kdBhK2zapWB70XhHssOr0876
fEil7gN+j7CukaO4F3CUpzCWEWaASscc9RUGZDa8NAIFY5gVi1nTg5zLxtOzXwcqlCCWhoKnoH+x
3RNmetF3ph6kubcWiPAX53n954kp5UH/iKY0Ujf1GnawBUiPXsWB29DD6ccwQckzOFA8ce3fJI9X
qrL6zCBbHV5ZTTYh1Ollf7hppJYugRkYvumZhDIGC/rWgoCICOeyomsIfaYRV4lrqOCIl8nLz2Qh
hKYkFxrUoNp8NQplpblxSVMcBZXCc+nrGBd2QmVW3T2z22zhUDINwwj1s221W4n04PlStRmJuN6m
dU38t2RqqfWdjbX2AO17IdsQBBvmTGMPK/uemyM9yLIKWtBtTc6jmMFdzylQE/GVbO6MqJFaoy1S
Lm5NQvpnB3V7+uQztVWqYg4j8DBIvrQoTKOUd2AzYiz6Gh8JPZAArWN3IP3eNWIPMj/G9cHo7nqs
o/l+5iFy1KBmK3QFbsDDDCP/A78qkKSQe76eKjUE5AVZ9ry+H8QIuRNEbG4Lt6w4oBkGponR6sNZ
Mj1lXAuqYCnumpddbs1th/WezB5pcHyqm/JybjxZZrZcxMgQm48SWlrB0QBc3ugvBeP7/B4FE+wu
u8reBFNrvCOnFPSnkv3WWAit97H/qAEuBzZvyhv5XK6srOStFrIMuT+T7LKjOYIDMDzrflvyKElz
Rb3eX3oRbfWr6/mINF0xCMI5dfpAYVA99lPANO/C/Bq9FQ8xCChQ2wW/Uk2V47qbG/VYZyhzUlE9
y3UL8qYoCOrAEGbZw+IyhbtzzvlOm/yEEStXqgDyWn8hFrKKIdN9ubYmu1l0RkCnLzjDyh50fHWQ
e+t7D9G2JoLmR4C7qLDkKH4dW8rqu8qCoUCcrQYgj4kU2KjVk7T/R/7eqMsWKzlT0h5bgIvCTowY
dv9+IA+Iyloky6X3YIsxEKOpAsUmwLT0HxO97njk985cmRoca0XxeaUeZc8OKvd2rUIgoaeUy/Dd
aru78B2JO6KwFrUnrsy5PsUm/uscIccut6VPQlACXYmBL4Ti7ltqu4R430xeS+CqlZHwVDQ/Q6lo
97IAWKewVIrNYB4yKe/nUQXGSKWndrnlNbrnt5FeErgnHXSp/GPK7o4NwMLMwMrtqetDQGFHrwZ4
wWDkFnTWEB/dCUEyOzfXa9wgJSrfQmc4WB4jRxJo9xm2+6zPepxnsGtZDMjEZUau1ShJfiG+N4ry
boWDF6AxlD1d6tX1KyQTcHE4bQlXLNeEd0E01Asl9Ns3VphzvcX54d1sn4T1bVYjYh6kvym1QRGM
ZElAMRWeBZD9EhfR9rJQNeeCO4A1y5gV9+7ReB7yFlspeq03T27ucUb0K/zfVHR1BnAXAHqrYr+i
IjJfx20vyQtuPuyqMaMvenTX3yIvtwRSdcSTq5JL+EituOVOAmqeVRcm7o2XCVuJkkEkMQiYyJ+r
mhXq1bTzsa/Km66JMZj4rg2ao8ZKXBzuXazjbqU7EA83DfObiHB138p0+9EQ5Srsb7GygNHb1u/k
AHGCKA6mBkxDr+XmE8jkzO+uYQpRchEpQn78UNzaA/0FIkXCK99/MjVo1/ICyUBL2KOrAHVENMsi
itYW3wsMy6dGJGuSlZQ/ZAPSCnE7X0oA1myBveN3DwMX9etTJ1qxfxFiUKKo1zh9yziV+bIFIS+C
EKd7oA+2MEbs5LszcUBX0DePZD8WffyI0sNCWS52BmkgvrTmjvPp1b0oI9D485LrrgN03blKMXLT
6J57D6Yw0vWYToAJmnV5cXlmPJeiN8s7rsCoJRvcX5enIp4qq21lJIYHiYsQOdSx6iZtzDPiBuS3
aF7YsTTcpXf0FM6KQ9vItrhfhqgMuDahj1g4BFDtyJqJGnxEp0emJ3AvUvkjEkP0p7Z+sefuBqPH
xLosWOZVzSm5doUdqiguMT2ri0F0rn/6hM6FDqTPXGh5Dw5UlYeqGx2rrDJccMj7strK9ckJAFgi
sFvtSIm5ilGvDoZQFjssvkZAEehBAj3MbraTUc3xo5d9b3A9ttZnVvtqH31tYNMLDZSOmA3+x+Zg
+03MJy9RCK0dwlQTHa4WhqPvqwKrn9oG8qCktjcEM/qUSEPQ8/PLbj0ZLaez2vdiWIzSDKLAiMoi
acYqpSMHxF6ZP2+UvnXcVfkrmsKYC3beaE2REPe2p3onLC1hUc7SBhIHrRY0wBfgoR7BeufWWO5g
UiALdPxc80GgUJTz98qUfS8rx3YGrz40rrClvIfe+655klkYAYYh09kvoiz9dILZuahKMKlrEvZB
2KXbnDVYY/LrYbo8z0r/UNZb9AE9FzDOVTS6VFZZz8Rp5sF2ZPdxfTnikR+zMmbWGlv0c1msMs+y
b593UfPyW8NZllyJHz8jvGTvMuN5NForujwtE2Xk2MRbDCjx6PYTeH9qBUzD62j1iCy4QC8y8r58
MZwiofwW4DuHZjmvg7wsieAjiGVr8WXU6P6KeYW2AEust55vfI0rBHjTi/eilJk/UaATNHW+3Gu5
FgUdelj25LJS6LcfjImobbScLrxu30lHkG4vtSoPUXGyBynMMoX+sHovqaDeTnppXlIKPYYufNZL
SARHGVUT4DQLHv2XQ/naO1LQjWw3k1FQ+9E6jLFwGTG90HMQHbVs80BfhorMPbHJSH4MqzrNMT+E
IPBmnJMhVGG/U3OSZ6OVkSd+7kOZozEEkDWj4515ODdFLfeNbIMnBldb0DyJ96rZSydU2uPnkNWW
1E1DVp9RRp0JHZ0C27aMxH3IjcO76JHgPeyIX7zqp6WBRlsdPOUdJux/qxL3an9tMMoRjhT5CW1E
scpqtcHfFv8tB8T0L8/nSQ4I15Qt/3bVFvm0cI6o0a5PonLLflGvVcFIcE0cmAGnNPQ+bEdhRHhR
GiO0Y97Stm4sxeytDV1HDF98xsaZuGvfHkbmrLdZbsuydlPtuxTnnXKUkJHkJzPCxSQ6AXpdlXvg
FWGOufWxm2cG74e2LusqaBq6nAyCjdgyMUyZ2rOYgOIlEwgQ5Z0J9JoPtW4kW9t9T9F7lwVnKoco
aU3rcrbFiGO8Uh5eTuAvVpe8DXnWeO9GORxWsq0ejiZlJGL2dvnyhYR7SRlebdTcHACQk8v9P5pX
bzp3IQ+GcTOhFyF0WU265DYym4DLWCQlZWnMT+Ra4M3a7j3JC4T/F9c+GddSE6xLc+9PDPGtMGdO
36Im8Q1YUb2POoV89VCrZsR5KOboGowPiuafiXZ4MI3zpw9PZ26rOeazYQZRCDz42Bx0afwGLie0
jQ81lGkPc9zbixUZqTgvlMBAdSqi8XHg7foO30Nzqdzjn8Vv7vJQNxZNSla6lcVJ6GhxDpmzHdFK
Q7OroTbkYhgk8vBn/Q8fk6U/CBZuGDjC/OT0Y6ndRKGgMxOk/H2QTRXaY7g+N34DQdSVtssBBJUN
KWxIY4ULBXi/XTL3QJ51n0YH1ziXpCZl7ntUtyJWLXDiz3Af9ImQxx9nl6AnaPS58Ns+eAAzmSa9
Lf1O+O0gIslJcFnWkYdzIVrAcf8rOxv0dALgwI265CNT2GZt9NRoEUOFVexiQkRdwaiuKsfl/JIY
EWrZUbiFzdpkmv/Ue3YUPgpGSlwGeDWBWiqsKFCZlWJavXW6x1pw1ukOFie2n3tkmPjtVj/19yWc
g00QBZ1kkNuPvbm8y3vzJSvE045Vy2ezqAA0yeW6Po/fBc8Y+/42FIIeArv88HGm5xbzc6ZKKbmX
IUl6ry7Nj6kEFaDUxppcNGmMy/ffcsvHaNhlZYU2iTwH1X2edNsgPOfl6a/nAKcmCPwcy154MGe/
xRb+Ag1+3rM5uU0Yhlyqtbh++Oote8G+ekx5W1p3WLjSzmqt2TpIMfZWvc0XWoyW2PNe+xp0gwz8
DQt3hisuZGUvNAGhRbdm4xV0JKZKd/yKBjqhgKN0aUj6MFNu1o0wbBVkOCLExRu0ie4AW2HVwE1Y
feqtbpdtqRU9mBWqCSCmfLOneppP9oKEofrtw0oXZ3gKPu4uUGIeKIirtYTH+yogw0se/4YOTnmJ
bvXXNOxZMbVLkFJb+O6xFlEH+AFFJnnmfSgzl5ALvxRibJsijxyVWM9BRh8deDVSKkvm+SDwtjT6
AQIJjsCgfd6tEbNBYLxBTKRXftrr/OR16v7VLU9G/Z3XZKaBx3g5/km0BpYQUhMy6GPPi5353rKF
Ualu6AL2LRgwLsmdEeP5VBpRVCc3sNVbBk1jgKBiwhhLvuocGCJUThThn50dZxcYuSdXaf9Dl3dZ
dXDCMD6UG8Z4y/SXymXznt+mkycyFWwdTuKVsXFf8R+e6bzxSbbFsFrt4r+JDYuEkux1OHZOezoX
bKZeKPu4MLlQoradPg1RGjhnZ3SAX+O+xWolcfdte7MiqgLLQuPf9YweI2cvI8xRtopCxlz+kk/j
cOyCyLhV8PCLb24YXggrBVreaNA1i+qY/QTVqhgnlH97qfkOEEhG6MkPrZ4EvR7zx2ajtFEfLvpB
DncbkVMINmkJrEiK1DNoCqteT16/XKSJm9V48netsvgBPsWijrMLMBB2all56UuDjrMydupXhGqc
SsjzmWfhWM2A4c6Bvl55sM/Ig9AazL98Cf9sXGp4VKabg2V05oe1e8zjFGo/CTNXecrGhe5pcVIK
dHJGWO89wJlmZrN9LbBhqaQtRBtJ0zZ4B/9cBNMl2lWRWaQOovtKhADG2p7OqSlZnM2kVBgJWE++
eG5xyH+0GjyQibVBUgauZUEZQ5OEnPCezMHzVhEPmeUKhoUlWcNQAP+rjixKh12D2MAMM04jiV7R
siAZllc+1QWSpBVLln6QL1AAeprTRKh929mIDfl3hfMqsRlv9S5SfYi//cY7jgaYUCdGKaIHUpih
EEix0O+pnUmpH+lF66aW1O0sFm4aBS8i/kGp2dvhNo/0gTD6UVYt5JTYRO4XVj02zA5GicYK5wEh
tVbJJ0v2Ri5AGvn8zMEfxepNojhgTvWN6VcASO6auW+bGR21AxKEv5w4WX7NqGDrofmc5Vj/PcKc
rHFb4uciOP7mFsAW0fwbIS6ZZcazLRWAdjEE/u6QVQh6CSzVYxafQ0x5S2XS4RCJ76CFA53MSp0y
UU9LtgUKvlY3PluuWLeL6qHPUVYt1D3TiyuqW+cTu1xE70EWc5A/YgnFO23IvWT5qFEa4elJULdm
Jk6WntN5tWuFVyqSu4en0JecvIhxRACkbgHKSrrX33gx3u8EdNdTtCAT33+IgPCBK3y/vy3I42h5
74sLN9vTgYyBxmEUdtdP1rV/5ui+0ejwxYT3iJC9EeWRQ+G8EESycHTa2Ym0OGO5tc445k8Mz4Hn
pzqaV+2eXgsoblf3ZOm4HBAPwGmsELI3uxSecbVmYCq5KLeopS1oVSrsgH1uXl5H+3WFND3DmW1t
VMLdIkPSWYtHwFbJqQR2V0FW/fJmrfPmTb53YG6U2qmIThI3fi10/kuZlto/MYhj5q0s4nAZBRNZ
9wwIbPdvrA66piAoxX7muey4Nl/iAANFgA3CT/b1glvHCDhH2f8E+PeHlG6JDJa1jOz/6lzYA+zo
h8Ni5H/WufShTAWBZ+QJgEIePa+U935fACXLTdpAI57pEYeS68t+fA15ZYKz203HvHiXJDjzxmXm
9D9ezPKfGgaJJTFeCR8vYxV7VpldY09xXBh4p/buZ9yBMuGv0DWtXrURhdqYdnQhG9u6GS7ho+gr
TiiQqCCmtWhiE02Gzx5hUOAyMkkmP7kX+w4YF0OCZGIQXakvECNN5qTWa3yne9jV2iAwVeoD1zm8
we7O26VnBHuKo6SV0mNRrQZsomJB89EKNoJucTQXx7CYjfP1pqVqnUxIcKwHXMMYjYsBIFXnyQg4
oD9tdOt8k7O4B1lGYxr4tEH44akqbYdwnjPF3/N3ZnwcFrmvHgZcCLmQiS7PrTpRi+fWtWSL/uvY
fKjF1aVDbO66SzuEe5VztkRdLROXjuzLolkWNW3O6ahik9jQfbNK6tb7+BOl2QQN15pNRG5bDMdr
GV4uASVTuzYGvoh5MxwBdCx5IwzW4zOaVE0vUEBgCp5U6TP9IdelDSeFgaCSdj10AieHpJQHcSje
DQSILTTjIvmINN98cKQli4u4MDpy+CptgEhgBg3BekAVWWbfcRb6ixwVJL2896ms3E+x7xJHdgJl
+RSNUhGhCIc/wigW0o0BRnyUH1rOTrflJbVC8ggiBOFiayoAxs5flJ8g/lz49XZXoEiW9cE0MIVQ
IgeAasMVjE36l79VK7+jvkA+B4Xc4AX+cHr95H7vwpVz42LT5jRqs7SBHzH/Z7OaKWoYM2JOz0Ra
tr2hj45UAx8GYLELZigfuwUX9cbej/i3xl4temkPyqVbzAL/RPQsIAZTPmtKh5JmHWBsCT8M+kWH
xfDqY3GVy5IvyPiU0DWoeKvd38dnuse0gZwVldZ1jSc3u2IE2Y7a8HMFTBevBBJDq3ap9tFAcHAg
B27BHAxfcvS+TtYpYguVqPIUjYI25ordC2YoryFER2o6SEPPF7T62+awGmzDqi11rrOVmpOemf4x
98W/CCRyyRwLqKM1fRjdy0WnOLBZMHYuaMaXc9kjy18OzQOkYxwrbInzcZyny+rjBoORGTxoNwCi
C+E9gQyNKa4d0YEC1SF2MhBMebWq+B3kP6BvKioJ+GslacitaZzaOAM3J7UcxqFUYg5zQJxl5sQZ
r5mo4UW90rXigT9kRDkivoi5x84TlbOwfDw/+rn2x1hchcj8k4nQ2PNWiZkYDIqryHFbUMeWhdfx
3TsgNDSl3DsFKEhlDJdA6nqr/NyNUVm9kYrP0Uy4VgV+d+I9iz7p1IB+lxmQyM6rOKjDXGssIYhP
7w1mZz/jYllC6uzuM/pGMinnVsRaTg74YwvHu5gj7Wabrd0P31zPc7O7IbGXrKCnwA+vwfO3hVAQ
RsR6Z80dYC+QbSq0NkHqoRw6F5yXKGliayTFd+dSMjQ2wERenpKnEnUefHxVRkLiK1dEKl/Iqh/6
owJUXT3aP1z3K+RqJnDg8BtgdGxwmLIdMTDi26o3gVwRxSCLjx/ZJMeDBdCtZH+WA9jkIGrDyUf+
ZiSnzJMwooplHtRye4Ip5tEIZibs/SmR96mx4s1OE6kgTS1prhIqR1n+EKBNhyGiytenJp9NQwWq
+mV/+tVyXl3kGhGNFrC07GmQu0/MkgiMLpkHNx9BBnKUNSMjON8pX3tVNtA3FDVjdwxSwSIELPQN
LO6bA3skx2A6UXCx+T4Yr9XB2Vd25AEglfMTZgUw6YY2+bZPOP62rB19j4c7vi0SrxCiFbQmt04T
tek65xOXT17Xp5E91zlFZ4btnTA9aa38c7m6nK8pNZXBLIi6bogvZIDJ12dnXDO2+97REU6iYdaD
5/y5f9Sgf/ZLmnPYo/K4hYdjlOH9LQnT0uBC6pWd6vxiavbAFcWY62L7wJvx1Ysk3/yxlMfhOFDc
wJk864NK2DLaH+rKsbTpSbrlpDd4tntEbopLML2qa7C0P4XnTRCsHOEoZ5txWj8oYadfMLWaVjA7
/sqL4beE462/UEIT2wbrDgYSH/eWV5L6HWD7LqGla6guLP4J/ecSGU+s/X9Qs0hKe8ENF55At+58
9iKZXbaqztvSf8ZpWaQ0R+Mrevwc7AgqCv2eXUtDBM6+a6seClaXyQOQBen3NGzGR2BB5Qmi6Gz6
/x7+rbzzVJy7IumBva2ymddk+/ipioEugGhBvmEGxmjyslAwHpER/j53+2mdh/tPyf/CGdhyZ8AB
KE+/pEH4fYpsxTooSdtaip+ZktI+GiCmWXzUor6nihmGObGrZ3bUccSt8cQc3OQq4WfERPei4QHO
q+flPjsFXV4oiq+CM1NQ+vrlAbv1yK4x+wwJ/IBh0RUXsv9O5ElbB+7+LlGC8wFZuvAlZ3Z7naqW
91oyV+EtXUxvkMHbRWI+VuNNvHkXFNy9kDTvC3zaHIamN80uYW+/RSNwwSgHDFJ8OTTOLszprI2l
VVjgZlK1boj3uP/fKaZP5uK4ifuXQacDDQkEF92JOcPmHtJkrrpUL8Razhe2f0WfrmA5EKdt8Cc/
Tmn5n/RzPV1DETg2lijm34ZSV2ociPG/mp5+cKfodZ0kb4uwUxZtBiTEnfKM4i0dZT9urnv/ftpF
VRabfk14EpRsfD0MrLjy7+pVk+C6UjP2AR396jdB/2aoOr5v+BkimJxlAsGudYhCtUTmD6nUD43v
ZJoxPN+vVRGc6ZL8odN/WoY6Je0tEHUd6kdP5VN/gHHBXvvuKGwT+qwGIQUqeAD9zoSAqjhkekNh
OQVpHQiej6EcQZyXBXltb1StXqKCaIjZZQPA22WIKOR29k2Lrr+kgea0Jfht4eST8Nph1Pen6qUv
MG5AGLOIPcc783ET54KNNEyWxboex6yEn2iSRkhAEeoVhFtjdDft/WE3vRFpaLCb5lkyI8Fd37zw
DhYMtrqXGq35Nm/qBggcSBm41MNOALpr+h22/FBKWD2O7bvyk3cfH8u0qq3hKJHywGBMTxkl/5XN
kZ04fhb+VKMtvntInBCZRSJMTEZ8HebVC0fY9xnsqSj46OLQDzWprWfYK0GxJM28IkH0dLBQUC8r
bp6xdY3c6nYcphPnFkcqEY0LdVfC/e2Zu7eQPnOQVz60DFWvLTjAKGRoXqO9qq9QYhlucF+HAi/D
b/FQBDb03AhBJEsiij6dVas5vP+//sB6HS47FKlMNwcLuEuuKiDUmTwAzYEfcTnyVX48wHH19RTz
ef2FIYl1a+DheKHe/GrVGksYPX2pveVmLVMPwHd/WTurlFM52DfuCiXbs1MjhRrYV0qyaxk33Kk6
pE5oJ9t+3EOorjwLx3claJyaYTF/ULIvundbtaWRkUlNjCjTtVu3CFLTnzb+rC7S7AT2UnxLaD5N
k6xzjr3/wwJo+ZaYP/1h0kqnp8Ly4B7Vjkl7wPTY4cE64jYpINcpaE63pE6oUqgprJy/dZcHjZAo
1zWlLZ6W4YN2qPAF434zRlztxuMAmEdZb7uyvEEZwwEpDipJQBbFC+m3QP3MCYLdPwmAS2c16C8N
Cdati4obgDZQe7H4j5gRKsZgtCKhnN8TjZqTPkCZOXOs7r1C8psxP51LyqYrC/kPeiiqjPmSMyxE
P31ZoaWILGzMTDLHZQ5/Z64HaCJOhgyTKgAoV8BZd/dI9svEKwhtPuzV5uuvbloQByUESYxZ4rk6
kwT72TZSvL+I5EBtU8jmAu5/LYoaXz5o2hnEOJ87K1e2Ku3lPEsU0IQ4S3/DUU4omizSY3yobtcW
qIPsS3n3i2c0jqquwrgsb41yXdgIHzDHuFG8WVuQOFeQlozKCOC24af32Z+JXhenExGepo8UNlWs
T5g/aFnaj7DFIluAP5IHKvHKPefoVGNuOZ8kWRz9a+eTHkq+UblNk6zpL0yMK1nwTXUpb5GlCm2u
NmX+hIqHCwJHuBctIDPQHDWe7Jnm0lFbJ+lSRwph7C1PgsSqxxCcHmoQLR1A+b0iYrKJcpCljnCZ
pkzpcoqubFoJlZxpb2NyvDgMOMxkyB43d7eCM/8pVW1SViUFhyYxreXDMNercY8ASv65PEl16ZRM
BRZniVtjUG+Llsd1UABkHh46xGtRcxNSsyuwQBevfDV7J6RhMTdBdNRGzpNjSu/JircyaZQJr71l
kUm49P6y9YLJ5siKxOAZU2EyP5zjiLGnAze2v8dBKODzOTwPrQdt+ThG69/ZW193bgPCz1nxcruB
FQDFTohxWAZ39Nce1isoisT/Ut2BiYcerH8xJJMEHM6ikqPv+QFrwQjK918ZJaJSBJWujEJ8ofbN
LTwtYQnq1K4euWNVNZg+zBFa+/H//2ldTnODIeLOuaRpYL7gf74883Z51PS5hVfG7ioP34/AqSXH
QkJnqdECBUX/rvEv6Gmp08Qpkfid9ghh4eoWUyPVmmkB6KOwbnmyNnBSr7z20CFquHZnpUGeopWA
T1ox+w+YZBAjx6tFoOPZdzYG0Fpc8jq3COFqE+vKj5yOqX6KPUuIVgdwZZqtE16l8Z0WVFtZRlQP
tWU9ZZbyxu3mlTaf0D9dLTmuJkA/g3WwuzkAI1VikEKumIB1CXW4nDERw4YICs20C3uEpEdQNXH/
bSoxCaKQbMCL/rvc/O+KgQfgJ9KFOVCPOkaz92VZpAcH1XlX3jEatvOq7cuzowLHEjP+dMJjFU0Q
dTGcqXbD8zFzHEXzKOSqKeT7op6B3+z32PLKNR0qJQwMbh/Oex9ZSo9oG7wSwNT+wAkVjQJa6QSC
E21YH9391r+tS/bxnFvNXS2nHMteRc24hpJgammLKFmG/mhAnXzPlST6s+1DFsPLzu/O7D/tbdnQ
AqrHwW1amtg4/wIwqTP+3W0QCowjQ4Gbia6qFme3/35FxMsapZ3pGz1XkOoDBZebKH9weVQrtHQX
LEgIRRiMs/ISR++mN/pSBLgdLOcZmvPqbrz9Ns7eiS90DkbAx7qBX+BTrEH2CgIwDMJRW7SjU84W
KWOzPjtoRoAF5hyvQa77sR0zfNYQrmAFo9R0vemQ4FvWqsaiCTd8+Es8blXOI2Jv+ktgLM8jwsyU
xOF4uItarKdBD3oYVIAnjs2stqMhxsAq8ycu+8b/8rCPghgJpoQzCfs//K6wKn0jJoc1Cn7smSSA
TpwyScnPns3QCBvCiyC7/NMTXaaA8qyxlbMkuxyS3Oo3sTbd/dJwFL8bFgdaqKRP4j/5j04FqUBG
cKNsz1xHT/jXNd6OW7cCQr2e6DmSwMQBnNLcRDT/Gl9cqoccmYsriCPAo+gjhJp5aBdnzhyGNiND
7xyFa0N/770uJ7fsC7AMYypFpbVdsfnKT5oDQI4L5i6/hawH3vdhdSAuGpoJwQ92P1+cjwXKYlxD
3/7uZfcuTimVdToVLQpQ8zYNKDJO70qZqufS4DbZKI1HosEeNkG7qLUrmddBizeIgMXsyZ+7CBfj
fFQWm5Qj/qMLO6M558JIYTcvn99H7UxAGeYF467mn/vf/hxRVtjvNhdVkEmpIru0N2Pubxt8jfcE
k7k55+JOhqBiPI+BvspdgENdFIqrbFpwZLRiI63c7bJlyhwxdS9LM0b7l3YCv5WaiL7WiwcY9QSu
YXaojyWYu/RfczJEcvu5hFaf7Un7OU7uyceXbYux4IBdLIklXPU1Q257MK+7uqkToFwPlabtRTzc
zQHc1yWdZPFusqwUz6nQP7azPio5HVCsJlpV5p+TEiaytzJVP5o01Dwxjc7wum4cRP8ftgIfmpra
A74bQOIJzttFIqrpMRsa+H4NGN9WECCjVXRYIFySMz+DflB2KisKoo4b2vU+K2tgtYST8VXynX8v
eCCnY1LMoWzEcZF1q4c/JYkcbwex/wHJqTJlPnPNHDnHZi+QLOliy30NGy10phiQsi3ZIu5cIHxD
7nQY83plKCmD39LmFfsb61p98Pti27qdDbaWC9BGWquTIg67F5auxh+vdAvzoaZsVgP3fOerDzdF
PKYZ3S89MU2r1H11hfcpWQIbuiUmMTiszLDmmbQH+kdosmSliNb7VBl9BFGGe1XPMxTMaSZJqbCK
VnK4QwQi4sFGCHzyoqrXFCP2A8OAGpk3rWezs/rjjDZRcS03YE9cUdC8QCCcWA/v7jP1QF6GMMiF
jSKtNGceW1Che7/DN6b8CkQciWnK3OGXzl8j2kD10G2i6bQwv3224ucl5HohT0h05E14WHRnqmA0
XsrSKoNTTH+UEg67AHKgZtrFYBn1OFudXQaxPEHHuzZfxdpj+UvmVENtNLv2oEh1JODSCzxqqCRc
lrd3xmTo6AnL6nqDMGxDfz4hnLj+ZJvm1We+PY4/pFmnLa2/65rt6y4ZK5zI19aOS8g70wcFC2L+
clgrWNbhRY65L1q49+OMQtCm3mguVeQRrcF35ZjaNVUxfBT3ZNy0AuNaBwaJQHQEbFhYO3+R0M8+
T/p4SKBrXJAOV+n/YIThXyrkyXzTP1+O61Yy0rGSNWdPiZr/gkQ/5Fx9Ev2M0/36M5RE+EYv1slh
jyT1SHZk0trKEww+jVS7tPVdk5dFY9AWzZwEbItlvnIXYPV/RFndQoX+acFhDwz6RLstNrO5ZaeQ
KAUmWHJnsM/n5X17AS935S6mrbUpoAzDaOjHo49XDFCCtu65fDHz+c4dpuNUI96Oyjg18iYzntqv
4wqmiVVNYNLN1uWxwX1NwxOwPaeUZdq4OW/QUGnKAoePNZRl+FZvNlYYqUnLUTLJURRxB+gS8Ves
S4YoYCh7O7BhRdsCNy8YbOqryW3iAQLUjGCQXUTMgGz8Xqwl47i/T3QmdXM2Dn9n52MOWIxZOYz0
fuka9tMHOTNhxpw3ycvzSSQK6Tq0Oc7WTdIDw/axzXUJaDen4g+qoiLuDtySedoc6I8+yoNAB0eg
VO3cWfMfiFQXQ92Yd2EpdQbL5gxzsYVM6dnu7/gn4/tozHcDcn0ZgFIrGBkGJI/TzmKP4uhNsnwX
cqug111WzTdFcAV3zdwVnCir1PeV+fV+6UBz5He7tI0nhEv42Hhl8WAKye64YAzwq76QWe5hOON0
B6WSZyXpluv8PfM5SvhetBKtJmhdyCD7qZ2kwct+RUTU2kaKVkYpZWI4yDYAs6oe9TiJptwRcQId
I2MeooZ8yBHQSH0qlqe5YDCGcqGNSINyNYarMyklf7mivt+u8ZdJuuuLzeF+4Kc0btS0TnddgWjo
uTtEA5HAt0ccT3GajWGZEGDrN6o9aDorT/ISQnUqFRbh4aoierR3dRcvrtnFdRAE9z0/MIGVKObj
+hkvhEhrnZQ0mnHQWQx9KDsjE3Q6h9SCHcviEQdiZdoazSdQkPrUcGrQx8t8Y1xHsuFrKmM8UMxG
Fi2+BHD4BnCafKsJpy5hEDnZLQ32I0U82YPTPCbK1p18GFf37FbwP1qejH/0UrfyxdZfyBiQDIcb
U7AfaShb/0TvRxzKy0msff7lnfY3JFGo1GKsTEbz15gn0U8WnD68vWs+JEXt4KFl26MOZiLVpL+N
Q7iZBUizVHK02XdSsNqtZc+UNOrsWL1hM0No5MGhjwG96E4IqYu59bc03hXeC3rkmMn7AoUF8mcu
J7XpSqz/GzUW7TUAPHaUAYTNxODze16WA3em2SeXjFJR4iiyI2RNmUxOFXhmnNEZ8/iYDjnJVQO2
cADhgJVuICRas7vNczyJTvYehHHLzhxrCKYxJl46+pX1Ome9xYXgIsNNt65gMeMm8BWIElNI/UMe
DIBMUi670/AXM2YsrRjDCbq4a8nz0wJYBppV/TGBhvhce+vA4QokCmkVZfmcr+dWRWJEl1M6nfkJ
eBLO+14R9vURbZJ+rySfmWwq6sgIjkuTaSSQTVVoxOzcmxV+97+d9xV2xqwCH/5DhFZwA7RrZ+DB
8D4Ll231EW18bbuLyi/RsbhVc19N0XqZxCCJ5qMUNJBTxKDxWEFSdJsTUatKn2PeRgqwjDZYXPsW
YuLWmvnGWQ9OBx13nRUZdvRUxlaVvBTr/yCpOYWpUwBUbh3g5utpJVjwTObXjfpsorl+frJhihvU
T2KornDi9rZOV8B+kRILW1KtwCvZg5K+FgykkbelnTQHjOrKyIGjYFGqbj9OL4PFJcFac6W0BxY0
DQw7+xDzjkpUAHIg9XkG08IPRJI+pXRMa/5uJf5BLZF7hZAhCKrV+mmx4XUost8afrJjs8rX0tan
HOF+4hy5po4d+BczXukZ6gzZNGOS9G9VkeNg+Tdxpt0ky0hTXw4vwhdqUPfHE4nGxxUiGVCQ+qCW
1k4qPWExG+i47JIu+wBujzpUMmbPhbGz40mmsM9aJZRk2rtfoGZf1oDYGZTujgc4tI4uhAqN5b6c
56R5xdIifK3NzK+wpzcNRTxh+T6Ee3bOFlaC1MZBpZVkZAqRmpLQMbAs/VXR1kpStzxpbsyDmHwy
NIAQ/hHxcDF8CA2ewHugv7P4Fzh9+O6arhVdFruKSiYIgr/a67V3UVi2GOdwgQmctV+nZw9Ivm7A
MC2K8LeQewZsfRHzZ3r/EyU5PktLX39SywtQwIFTdLs5vTiTEMetUqf1/cS9O0E4DlJ2VC6z37Mr
5YGrwdD9AD6aY2TULljfR3bSuX+xpSnpmY6eo6tb3E1rYX4lnCghF3KTQuL+Ngh9toAejGhuJnk2
4UlZmTuF/eLQqvDsPu57MVJrmmYVixcYbM3AgpkyLgG7fSH/J8Q0Scv9oq22QSoi9I6y6N6EECyb
6eiklDaBoc0xLH2u+UzcoFYEWyxYrgePGMdov9T0JRI2M+z8GkbCSSz671qzFY2Trl6H03Xp7vSY
69OhkgnjYCWrEYiPk78J4rvpQtXv5gFtCRss9FMjJhkLqXNLSP+y2SkT+sbk9++/TIO380aCmM+E
C/6j8qaNn0CNGVJ2mz6cHdU9gfHXV/A957brpZyKckT8GS0BnvXyZoKR+kF2fKVbY0MsCSK80Oxj
rhBmZYQikFTjLBVTzit4cwmBiQLTWZN2G8qpJqJfbvhNJpaHFlraUSDswps1J+jX+bukn85xk2sH
WDlVyBLfYj/aHqgNr5u+EIaAz0SXHZYmC0A1OiTjux8nRuq8jmO0gEvydkryHS8Mp8xiZBaypc6D
HZeeH33yXqOZznxybfOy0GxFFrQMwnkR6+yYyGQzYlECN0xswwhoMsnzRU/OuWyxc0HP708ao75e
QTOoQ6HBzHEFrLs6pwfSr/W1xXDNis4cwRC83wgrQ8G87SFYesAv+YJvvPwVo1MVfx1n/fdmLS+Z
r5vujkajmTUKC5pREBC5M7XP0qcukf/BsdDCa2ETBS5JMwTqEA/96/34BxKTiUrLT7elg2lv/3ln
a0OV/SLDaD5nDvOTOnNDuHJCq53GsFLV3bxSb3FsA274uLHny1FkNcNCfRKqCOKRnnXUmT3fOyMN
pqwJI1a8GzeGY/WO3mFmlcmkbf7Bj9lmyOTxoejzzEadFj5iQSD/9j33zpedaWiP19sOKgxnwgeo
t1dtw4sbWqb53eWeOAh3on7Qo3eJTDtX2mmPxGyfJhBmKFcJ8vXxy4lRKJPuRLu+sMi7b2m/HioB
gZRCkjA4KdyeTR/V4JBu5aCtrqKnW9GPYJvv5IXwk8W4LGbHAjouLkTt1gW372tUVr3HFxgwBtT1
gbpRHazR1HI09p3nr7DYYQMcesOuN2zlTnUpCVYrH+wUYh023tU2hf3lUg6es5ydGTjsJPZEMJrx
eYshk/Ueli3aBuSz3md62jBBy1LZXAQXMxkay3dw1VKiJC6HVXo+pqySsUKB/gk8djc6GVmZH155
0c1T4YEDn+Y5ZhtEjQhNgO6/Qg0z/+C2TowlSsSBBeNl7w9AbPJxNjWXrEY9UTGMWfKqJbQKE9Kt
AnZKP53qIE1fRsVBwG7IGmfIZn0hcnL6J4yuk0W8HSmzoym0VpITJ7QAGuw34W3SUBdPTXoP5H4i
KztDw7OS/UJBDx70tt2tonyaXoJ4XinWL2tblh2u0QvfqN99dEywsIWjhNX+qY7gBVenJnOtaNJU
lbdyK+LtKW/OS2b30a8hvqQOcPnI5D7X2Rod0arms674Nmbh0V7b29DupBrizPGWxNOHaa9Vy3N7
JdcDWm0idkQMnLxEn7LgkDyVkw9yQrZ8GHnIv3wBYLU1sZ1P34x2ksanfDZ7aD4w4zzL3Lo+st1E
89N9IpgWm01NdoAAkiv8P1BN3RRFiwf6/cP0CaGzibyX+yuuT5YuaRLSEtZUHrVZL5S0yacGlzL7
b4MVSitt0IHM5lZVpWu5dfMZFOEBqS9nvscHyN6CVv7pBkmLfkMhpgv3dbkiQWcrTYgjVkp86uuy
6JUJv1nH4aksHOb+K5mWYyvy/Sku7S5r9Ign2pDc3qajalqhFcYFmPwvQITVyjtAzRwKhZJlsm0P
H5mvZPIMi76uG2EEfRtY2B8m++W/h6Ohbpn2JbRvAAqJ6G4HRNkoPaykJm/fJ87mo6spbmdFMctG
J1AMHFTevUhUSx5PRfxB/d87TmN/MQ/xoaMBXncIuLnzi1kkBJRROe/80RC/4+2AGRywYyG83rdw
GmneHPQAO21Z7HQsywFrS0J5KKgPWV3E0GaRwBzp3HWzMMCLFq1/VLfTDQRudTJyFj+iL+1G831J
DUibnda9pk6NVtaFZpHtWv4aUL8CeF34cxXmawhcWGsY1Gcm1SZH5BIt5k0Pn93+Pixlg4EBBgVa
GCWPaE3MR4ZdbFqebgQgBy6ygAYmuJKwvrd4s6WYgGHMyy1+V0R57Ey2xoIJo2h1LypyuFebDx1a
GQc5aZldLYluERHzskJc+g8W+nAE0y+iAwPHxo2Y2uEvH/QKN80851tDrrURNDaxFU+e9gWd+2fK
vqY/zCNDE+QGGuHhfo32z3UlEIKp3ZylhWRnbVckZn1CrjWlkidvR7CfY0Hhx6L+GguwI2mQLwPE
o+pgIF1qG9STb71U5N2m4UIejsfzQh3+cFxoI4nMtm6T2X2prN2T+IJX8t1bFLH6D09bh2pFYMul
BMkP+z+5CpKh53On40hHcPRFmVfn5JcgRlJZTmgrgKoSZpqKEmaiLTaJRwtLfTfF0+JH7u53lgOg
eqnweJjvGYPRKSN5d6YfNWnuXlI7K0HKYPAk8QNjixGQvBoPHRckQPrsCVVd7qLx88ZT+7lPy8mi
wBDILURuMHlFMGBCKEbf1wXpHgEpdfvJEH8IlTqey+cHy/xrOKckJTVUJoHfmSmFez+hQQ82j6/x
ER95+egEar2+uM86X5I2JFJ08oIMOyZ6zVGQfMSwJn51REdVXjaIn4kzTItk8UOmDLGUdDT0Pudt
yV1I3GcFqC44QsMUJpqp5pDne5p4fAnIdPgYY4QRBuqAf4LbuqhqNBZeO1Dp60eg6BSkydZ9tBvQ
vvrilb6J//sPtQqcFINd26f0NshGcOFEG3z7H2z42oLLTwgQFDiwcTz7LgyV+loIYo9s4wCrZtgu
wXbf0OT3R8ntCCvBImbDLlz9bmlnxPNXspAVzamEkbwJANaErZkUmlq/00F3pQv6feGBXle4xHZP
o38KpJi77bJAN99bv5+VcIpUKcZz+/ZTOjAefp6m4eb8wSUA9oLSsmeKe5pYx7l8I/licyd8k/sz
0+a4X1UuvgTmVviioPfeb7BcfGDUswdJeYFOFNcoViJP2Di/23lB4ttMXgtyodSZw84SeM+dZi03
KlSqPJC9xcYQfMmLGx47anTiurUg//n1fyWy1iiLlpeU3D8QDqTREGmGCI4QLqoXOBGnhlFDaS3z
7EXQ8uVNqa04hmZh260qV/9qmxq5dBehj9fXKOLXgt/+0uS/z2NzzoKVXrY/cJdQQf5rku9xFEkt
I7POyx14twACVqwaJzmNplzSjpuB9ty7Eo/bG5MEhg61ZNRLbo/Zn/EfxjIUUTHYtoAEJnPLeGpG
pe3+g4M29f6JH3RpWagqlNIQe1Ag3z+KqIR48qzRcCt68LOHHOvn+m+aMffQuWum9h40M+XjAP7j
wA0XxoeWXXn/6L7eq0Hajt+AID1q3+I0VwfkEVauXtiav3eNA+7hsMblw8nP+7arnGnfrN2IBn4s
7MFFSxys2Rm5KyCmTXInMVX4sOZvglWxL7tBUX3wQdbQEDuvFaq6JOPNTNRPqB1704LNF159KC7W
utmmrcRM2vmvojVRCv51Jot7CdrRvdTWtq67lnyI/Gtfg4OMXbcZ1fi9M+8IKQ2xItNyTpLQ7OPm
sC/+qiS7Q/fj1C1c7mDA2UOixEN23jeG3Ds/K15O5HGPbn56d4K3Ub07DZnS+83ej0fUjj/AJa4C
QGguNIKBqa4e5FEy2AHNADtOPSHdU/zRjAFBG40FDrKywhEEGx3iZIAXPfXBT7ADlCfK0QoXV8aE
VpATYIVZUMD7uOme3Nop8YQtXFDaJo1Jz0oVUd9tCT7BCmBIn+l+7oNWJMxlCUyEU4UIR+gM2SBC
UM3ZP8vcJlDfwnULcAxlnguX2AQuS2Chrsf/aAVHWV1VoHgpI6G4K4j3FpAf8IfWH+ItK8d+F4mc
PXu98EE4pAHIV7RrNJxwYwSkd5uCHJW3yLXxblCfn2TYwh4szV/TMufeVu4xiiAyyvm5PmSOdLGW
WtbMalB96I9HkQQH9i1k/k2tCqb9nYHDIRVAye0dHfd1rqoUIuFzDISN97OGJ9ihjBnIytSypIO7
61hB+WBEITprn6fq31U4o7AScRd117AfLLiis78L4QuRMMwXDkri7ttwt3W+0lYroKjxOvleDzmH
R+lKeKL2hmYp2OwrrMIjSrBozMQrj9xhufjS0+652krCf8jJI9hNFkTGo+zHc9hGZgZ0+8Axz55S
97jX5udGW7gusj43lr6sOv8b0j2vjUkcMXii9T11I0a5F3SgYelZ8ib7Enj8s9rfS+YTdQ0DTgkL
xNdvR1bf+CMyycJ4LJz7xTtWZKCYEWPUUK3FrH/4n8HyOu4Cb3Ys9ilu6KbROa/FV4QuTACf0k1q
sH1Zf/91r/UXoBuKdvFNJb3P6OIMX2aZrql0CJ0skcq1n9Bbycb1r3jp+ThK6aOwqgAoefrZG6uV
CW4IZpqJNAPdnM/0PsaTk/XXDCpb0o0UhZiXl5oGYYKjf/zPM9+u3JYxwn6gvv6I9lNqUy1uAIw5
MTPPVJ25Uh1Dr9gGxjBZteqAb7YUA9LnlGZIKisLOvH/sy0Xzq7kOPN3y3vfkbLfpmHRSxaZlB8v
d5Em3Vj6wOKk/3FihWTzNw2/5vdDorpE6AxclZN1Rzn6+7ERwpXDS2TXDNw6WMUr45jEgzESg4bE
rrd0j8HMzwzpuB1ybBnD/Wnc9LJDOdxfcMXux0Jk10jtqx1zoau5Kmkt4k7CDZGMGV8sDz5iDDDQ
hyjacbSfwhE/zYmJlNjxs4V8M+gJXRD09sVWujhQHxMj+cucwOVC4++nbfrlcm2tdueAaQ+FlaOU
0QmJudQGELC+CE0u7ilv5+hpGdHPr2pW0hg5bH0Ats/Vn8IhGYmItKDFL5aQ6uhEkbbbrc59aCmQ
WEK3ywGIWReqR7tavGoFqF+YWY33cQNZnbZPb94Yx88QCLjKH+bOJygZJVNXKF8dscuKDMPZBIvJ
Jd09WDvFCGW53IzZ+qskuuv2KZBr1gsGEVLXfK+iKGzzqkfB1x547w6HQ0pyGWV2roxUL46Jd6wN
FtljbFW3lvRFkLvCtl2VnvtJzELJoW2FdTqzwHwlH55pwTngXgqYtOuYb3rvp+ZmTCF8WeQhnfbx
7/0eBz0a2kCBR0gIWfrRPT2P6W1Fqrfqr22CbGRcx56lD6KgdjsY8EeDUxe2RpUuzBf4u87B08xX
Uugn77xtGK4hmZRoteBtELuxpXJ1yEJ/MxyUzIGJfp92W/xqV2SZieXSN9KEV3x+sZ/IrkfliIKT
ob558jAGJAJ6FNxDfct1dV3xiDYVoVW5QJ1qfupSA2+oxtm9QMS0iY2+bU48aCGagAKeHZC6GOEu
Uw4HVSEUorVdn7pYQDHtJNhzE4/CrGirdRRDAZhqzt7lDAE7PXASvfBgKDz5UpAWrPyFQkNakiwo
Oh2XANQ/0ZCoLXWaw8BvhqgprDXiCe1ibgmU1PbAjwaMoF5fA/H8a0CNotAdtskrrBwCq2Tsq8l/
VtV5/Q2Db5kXfTDQAadGBwxBZuVysE9q+XziP+o0cX0KKNlTJsHCQ+sV0Zbbt0qGgTfwrv6iCy9L
CXJWQWaFHOfSZsWKYCr0R+AVdCmtb3O1LWsFjt/UI7K/bVrZUOPVkI86RPAq6/9bA5fj0yabz3hU
Y+G+LgJmA/bpa7OCu4XHLJOLku3bMPS6GafzTu0s7gyge0PFWsZa6zLaLHFOhMoZBB/Gnp7dzTvt
+qU4mgGt963ecDITqB1NQsIeHNdlSnbolCuzsRgM+KM9MgUxvnnSRNjofSG1pKNrQG9J2FI2OGoP
tEjNljoBuR7GdOxU3sisysszIxXCkd4vv1m4yWYGVQtCBwezJbJcnAuY3e3FKU0u+vWq/ur4zxXh
Q9KamgiIxwPZgBb+eVmcR4KTaDVK8taZGbhRXAJYMhTM/WKRL2JqdZ9Z+ix6ff7aCb2xbWtwV+Ze
TgrWMqQoe/AwDoraECAYcyxZXFcwEIckNwJ0LPXAFg+wTrJWDRJFyTEnVHU0aAPc96myay2BQ9RO
+aL+cN5Y+zkj3JdSdllDo1bh2xcL+w97xHhDlFqBey5fnBNqr+8KwGJ60TQ1VpIVEKzqM3Btqkpi
PC8vJpv+93UTGxRlUd7CehWgBNwsiB9JqAzsLQX32e/2sVlnM1EA8jRBgagPHUiH7zmt8muY2e5N
QSbdR5+LNw0T3bVGfun/V13/A8m+9JiE5WvJHv5nvrcp+niEpPoBz+xbCntCYeTHhLcflb0MKmI6
Ow1B99L3kCR7xgSiAUQMCo5nzEc1uAmxO36a/AuZgT8XvY8zNGpkQrLf7eBtYeog+86/Jjjw4cIZ
1q1MvTG2TTHi3tDq+JJ0h4befAIE33eCOAvFGTdwlCpE541EzzqDc5eCPvmFFvZwX962q8kTtPIE
kwePXB0vaAUn0X+b/F20lTy9y8BSZIcqUIFSme255p7lMzaxqcmC/0o83uVLzYUX+VOLC+0FK1y/
vXV1cW0tIU0e3Xqww+FAjngxB+vdkQFvU1U4yuT8JX7LqVdrnB8Ktn4BaLnKCOzh6mV7i01WCYwq
X8u/jolqGOL0nUGwi62O+qGE5cubxKb78Xl1ZKUSLoNUjgXMRcq25U79D7HESQu3LRogB7Es70ZQ
sWJy3gWfpgNWFcjMKKPaAJN7FHHo/tKlMfLkm5R98hQpVOS9XuRfskAuLaFW/zVWz2nx4C6mBbPM
PKo1xmFSuuJqY91KeDq2ehlqD/sueO+nb5Mg3vm4PToIq1v337jD7lmM5IuWoMsTJ8Bq9uzo4acS
LJ2hB/E/OYjMfWJohxJ4EtnlcbMCsHgKRgYSWc+GGjTrh1k6vlQRHcDKhfjdnAh3UTL7Rc0/Q+QD
nrF23Qx7xQVg7y5ItwG9ywTf2K7a3W8FueNDaqyX80oJ7u9GgQdvdQEGOCXKfgRwTfivdzh0EI0y
YLBDRuY3vdoWmkj5mCdkjn6xc1/SNdA4dMZaK2UEWQrMGJuHTBN7kCGZgu3JXGIChSjAUA1VQYTN
6xeY1C9E4zdMQv7Bxx3Sk8LVXFul4BkjZaKZ9HINVWuU5sFGr2hmr7Ik++1QU7CzEXlipl6JxeJ/
nK4wnX6icpkXHCaRz1B9UaW53vCasJ7aIPxNn75mevIyxqejkCebtKhKn6BUPGaCjlJZQElGkiBI
YmaeGxOtK3Y+c+ci5GIGeNi9suK4LRgA7V5ua6FunCU+EtTS4loUZljRj47aesro5Q71MH5ZMXiI
P0cR1K6MWZyb/YwL70g4zGD0hBaM3gSPkHeS+bRk3Hezx5XpHiWU+6zWCmorCTiPRm4Z97v2bYnR
84TjVQYXGuZ5ITXP8oumj5bDWNruppcbRJyhw3+RlObAOIlyOVEcB7Leefk7fZAi/XmixB1etII3
dUCvKQeSahJCVg5Nqit+/k4smmo/9oIMl9kJrxWqFIlQa9QzHkU1KCpl31tygUa0iiYJto6nrOa6
PLORkcZXUNWvzsgQiaVuE1E//76GG730E+Dyc89yFWR2A5X3c8/0UK1ecMK4TBSBbMSQDKKkwTxJ
h3TO7oxMZlB/fIf5sxYg0iiGzJWI0vS4o3IVYtOg+f2eZB8uGpKPlRNNYrefJEd5V7QTtWQewkEc
nvyDabT5lRYI+XE6n8qu+mKZIWCRKe/TY+51DbuEQcR0Ee0yWDPN7o4yK8vETPGHB33ckV4qNboc
UweVI8pwNI9VQozVDYrUeN12e1RDMe7Yz2sb42cox4KqIzqA2ZFwuW4EK/cg5HQ/3FGcFYeKdVSW
6sTECi3bND3yeYT4FfkA+GvzLVefGH0cUYh1aO0gTgLNR9Dlp/Wjgix4AGMcZf2iQWQtQiV2ejI6
gpy9e0VuoTjuelEaygQQHpoaf8o3Z23kXalxc+84LWZjLHbPQDyMQzzYcmW0hkOSYKUz/4IQYd/C
UYslhUPiMVsceEJEs1s2NOX2GhtPOk40k39KZnPuxI0c0qD/lyIGnQ1nla/BWu9mefPUIqAFPwJi
wQIgB+MbbhzKLrKoQKm9rlkzVl2D/Bjw1VdPraHY5BwQzDLBbxH/51D4jrR/DMTPoWAg3qTzutTu
Pc0ad1KVILD6MdkkcNIUkVsXHJ8zQsbBqERxj0XiJyliOxgbljCer9RFgcWSsX+/jM6hGp4pgY/D
3bxfmVUs2ioMjJYX4FHd+N8Isnzo4srDOhjW6gwvoQwSO4/yA8beSaQvYRmiR8dkiYMAL30XnrzS
oSAqeM0odcCgtwARx/jTTUd/Pq/uFB5gbn5lv1whDZ8UvjZyZtccgdq78V7UBuxfTmTeuq7BU1+g
JfRQZcP2YrfHf26kf4wTveHsBJqYAtIBg6pMlcKeOOvvpBBGpBoiIpbYB/MbC2zdsSkTZdpZBqH6
niZE7Q1p8/c5wO8tIjhK2KY/nbxX2peyaBIRhp1tNXJZFIiuOJyDcPZL3yvo0rAZ4ONGVnXKdDQN
4/ok/DX5t0Oojs/Qydl0+xOqPmTF5A6xauyKjzMHfInYOuKiUT3Uvh6jzXCPmivWWNz8EhURRkwj
+hQgJpK3+GfwfGDL2fVwC8exRBnFD3F2DZ8I2wxGpsK52fraJYdJpSfvsyUA+LVwQHq955dGVGXR
zfcfm1GOUFVQWIuGZOJp6kekhZwsa3fMbIoJ1VG7N5Y5VrLfwplS2QxEt6M/6bGhznkJlF5sW8oM
usyaBCyNOEjTosbzxx1yTmdNWcIRJkKhUi5nu096MwYK0Ib3uWaPKP9wGhFgSAyUZLZjhcKrXI/C
9oJgu4LJDiH7g67Ouv+UJKqsExLJamsOSQLozcxebz2o74Dv5AgnybVwlxhLlNxThnQDq22OGgOH
8D/LvKWy5jneB9p7VBnabSXul6zZs3zxl6tGR1WqRIj4sOnD8gsec1jWM5tdaYDs1jYC3frVOFpK
l3gVSc+IRMWyL3hfl2ZNr6+4Ou2VJnKLiP5NfAr0Xqz1bNAtgo0YthhC3F00gK5JFen/3aGQFMtm
F0Mk2Cfw0oq8eC89qRakPVzuQ1OrAS7VSTq6e0CxIIJzdFFoRFOhwAZzrp2SSz33ByiX8stXopsT
fKBI9YfymdUgnCQXHcVfu04f/BQFX0ivAAEfTtBScvkJv1NySsCrN0kdRUyrwGXl0bXrkMqD8nvZ
qhhqlJFBbai5Fps3VhcO69F8sCUOlf/h3eMRLjcq2X9TM0rajoLJ8GU3WaolyufEEHvT3JtgGTSI
jqVXeG6wpKCOFuNheUvKAMhhtdcH9NHlZm6PpdDJkJodU8X8E3teX984yNOHNzCWT67TxJvcLBh/
Vz2Ur3sFgyHGY/I7OhWPPSHikphMC9vCnjehjA7B8x7QqBKtr5mbn7JKdAeDSSGrzd+3pwBf2AF3
ftl7Xe+S4qiI0rPDG5lQaHEZBERGFK9ET23uhDvkXIcu0COyMFBbqDB2u+2Z3SNDA9N9TZEBwHD8
dQR2xRfew+THYdg5DXTIKhNy9ly/fTY/ifMMSl/oGN6omPycUaosHk4ya2CRbBOS5TDPfNq5qzmP
JyT8aFr8ChA/neJtFoYEOD24vZpsQpxiMQQSNVKkp+MNlThdr5hnD03Ljwxpc/xyBPTFtS5Pitfa
xMxDalas42hPmt2fZU9nsMmeYzkcsVfie3i3ElN7AFg/NYuyrXL0eVRs8/8mEqIWpJjSV1qmj0TT
f1iXnt0LfPikGPhe4Ni5Uy23BH+9hfylLlio/ywtaco32kkcqF+/p+R7650vuLpfIYtp7fl8ffBn
HUS1jR2HnHVUNWvwNQsJIYCEAWnhTrWMuR/fT2T+tYikec6i8Lvzjs0/vxu+iZEcRzc2Tg5/DVm3
gOeJkpkkO55Gi+3pTJpTcVfYzsFMErq1cVTBrSGg+goeVlHTKnLLSG1TgKUr5E4DqgRlJW0ksSG0
kS60X520RU4aDX5dn9nhJNQ/lHgazz5ZCsn2YIlueXNDlWTwlHGIKQN3lswqIsGsm8XIrAy3CaLC
ky9CupfAOuFtG8WHnqPKhELVAVLoflqfS7UbEDfSlZqhdg0IISgqYxsv+QQ3+0SAIU8EsKdg5EKT
MuPRzEFQv474qN0BO0Ynq+V2p6fxpwaGWkvAiEA5vvRyK6/vNoAy9Haw+PcBD8NnEX8DKEHhF2M+
cI3S49FQ8ggE2T/aiB5KBRWoPyIa7UCpEyCwzw6XMYdYx8bYSqukZD4FrRCuj3VWurH9nmQp0zbu
dLyJqGO4EyvGmcR5crpAZOM64x722SapJ6e52E7mHPKfzH8P0qaVZT6xtn/AOSu7mx7iSzYjrZsL
MRR5VrPtmO8sWEJohkTlipJYLal6E4nhLAo88/CoDArvBbOrzSdp6uhuViJBGRx+z8GXvrjfE411
Akwt+ZF9CpW4GshKU0klpkLg/hndruKenZZrT8kjwwakHPqh+USrchhYONNigGCgeRSWFmxHIn0m
YRY0oaAfv8oobKfHuwnzqdDG+c/eSW735cPMdTwA727rBwUWx+zn16wjc9vzWLdR56OUuTXATrf4
eRhLMXH0dpGF8jfPqFnH8miW2VxXNnCEdY/A+fJBfWpxb7u+oCCWu3kwN5xb6c6Rh7heoJ4vF47T
HE/+9RuusPfcN/Mq4/9l6cESj4ZrWoE8uNhCxKm5NxAqqZzGQ6zHKAodJDhZJCF2MjPx4/vAUm8S
bZdYc6N7CpWS3MlHMOGXYtbBekLX19Mnnn1xSMY3gi88dev5VImWuh7++Sqk708c0BM+Sw56ists
okjeFGl5lkiXHz+7AGxGjDt0B+VQGfCkBpALUVluagFH7TT6YUNwNno27dgYPs8VYzJEQp5bd5KL
3Q8osQ3d5aCidzFuSFMEYt9buTqaPsp4ANn9pB/6WtOawd7YkcH2ulwZTpcClJw/nFuBFOL98S9R
PcH6Vt690N71oluA7uUCvnSZZsYNgpI52BtauiZGexS28/a632q/yq9rHmuJa4BD+wHvIq5uNEaE
TtiHtQSXez4Le3xcsGAXmNJyx9xGhXTIjKSrbzr60QVs04pPnDkbtcIlyNONLiG4V7OChKeN/B2J
0i1qLChg2Fl5iRqv9B0tW4szB0KiqpQBwBTv9bS9cOO/OfJtN3kQAtDL/j3iPKgLjHqZMGa5G2uk
qG4H8S3gKuCUeKtxQKrMSc0XxjidX+uGn/E4ZksgjFoHnGGIWKgcgDlKdTgWo5Y51BMeOHbJs1fL
Xu9C5g98xvPAdtt5TvsiPrUCgjnuY8G2C63DNZZH95Bs0tvxiRcximjQQXQBVzyPVVXvcqybQsq5
Uby+wF3fqe27wTvAwU+lKE36RmrYXf3CCrbVJCbLw2OKYKiWC04/byCSFZ8IoBHTLDALn5HL9BYz
BKRgGZT/0cbdsUUmBf4hHIqqyhie7KIWbbppTeJqsulmp9u0CPaMG7/i52nP2KehS3qM9TSIdbg1
aHc0YZoRiRXF6X/vQssc9THFokyRDpJNtJ8yc3VDV1nWpZu9uT+B9rfne0REgb3cBU6Gu6e8T7c9
C8VCYd/WNXZyFHnJW6YTd4TEEGgP9REu1WeV+jIDANiYt4VC/jc9UgO7rWUMVuZWXoJvyY9k2THp
8hfooo5xizJNsplG1SkkXwB7S53TEBzUCVsNJ5B3LBNbwbqr2cPlL+UR3kP65fMbIyPgdgq5GinW
r8s9ztf3dDpitpZxW/DzMMcO7y09NEA6hZ8rYTOV0WIpZj05F91/DHlzWaclcLDahHNQdS0Iqr/G
s7iJtbJCDwjUYI7VaaP0DFguWwVgFQfJ/ulDzBLtpZWtO+4PLHVvrTkRciQjb5NO+UwsCgR7J+NF
D2pj6RFo4zY/zsUXKm0lkOwT8h8qiRzmPI3pPk9RDgGYbmhIEKZmIhCYcDvJS8FCvANDJ3C3E1jD
N0SDMkHBGgfaLYC4pa60ljHA+lONJeOpDf73BBpB8UWjHZS1rw65F/Rt3fyQYrGZLMvA/rllpUxo
Zp+7Nu8n+TiiqxcyEFwMQEJDzjldgbYwX45Utj7JytDlNr1pBxRsh0II0d64hkyr3HVVhuG8SqE0
xDe2L8MQwsIO22x1ocEWjorIN0y1SoumQ9pPSN0BEiVf0Q9onoQoY98KIOR+sskYkH81TeeqleaI
QLb2/vvQN0zAwnvpG9xyNlFfm2W8meU5OumPv138SSd4kgnB0tPTt0RgNwPMXG2DNgkUfOgRgpxR
XvPGeKANGwi1ncoks2jSSXADk/tqwgPv+pxkhbpXSWp6B85KJciuHuR3zzkm6+45hKcFyiJHLkMD
jbM3JZmhY0Pa5d9tu5JXIFoiAGjNzf4cIDD97mD0ndqkZp17yfA8C+/La72VUggrgY4UwnZvHfJa
xK1ZvoH2UMPtRjFyoUhmNyvbGSJMW/tjLSfpzI76hjrbkACOT9Ez21gqzoGV6an8EgkfcD0vkFCb
cEfb1quGKjEX3LIGq+LahiGLv+jjBqbflHMsBXqiODFBosIn8ZYh+LobrlPcsSuhXRv2hXptAeDK
/udR1dvxmTc2RLzJAK5XAXw/2TeNJcUC8Yibk/JuIEsGOyRY+GwHgrdC/ldvNywWkemSO8nwbc0H
RpOD3Xsw6pQXQQHa+Qi2XpLvAMld4XdXfpocFTcpPzbRm5rjMpauFbDRUQGJEKIiGJ2K6Agtt+3z
mqgzvHAByD/ERAnD+lknjG+LlvXlM2lOPbYZTLA5FbcHkgFHLeYajABUV8sKeOlXU53tRwERZpD3
IvdstJbRejPcgxj6I7lS0p7WZ70GkcgiBacUx6Y92URs4xYxGzOkxE8EwdBVFmVIP1BL/G+ooTBf
LdEs5web4DqjkEvIYyBTXctgflknGKF9GqXNquIIQm6pkmqm+7W4On6NjIuMsbQwOuGH+AFMGMMH
ePdroSsVGTZJT0FA+CgBAwo3FG2GJF1LQ8REHVHWg5Tds/phLyvlAcgmaquwWQJigdPIfDhiJU8y
A60SXCnnVpBekk9GgPG9BL/WgCG5a74/YLGm018PqWIqCF4Pkoch5ZINP3JQ24paFAyVfwfW6ri8
+5ub6p2ztBU6ewq8PH/EZAv1i3qZS+rbod75qPTqY+ntVxYYSL3KPkpklCCDd+ZjfLyUQ6ErXRh+
A1Hk9xdHwf0JlFN2sJSBZkOAUh+5KetZ7PzE3EOmh5iheRAd4po8kDJKt3y5eALBafTpuF9Q3clA
1i9iKZr1w3F6dgp2C8WwQS33VpZDdcevezyGCb/9eE7zW65gLzA5LRDz/v3RxK9oH28fKCYrn+g2
Wleo8s+gI7BraYu94DeQZMvwMoPI957Td1RYb4xwBPjTOoAbgKG5cJGOvKLyMslPq1Z8XGPo6Wo7
IAHG+lp2mSHd+yO+qTNmDsDdApSsbBVihnDqgr0yZULm6USQPgDYfNwDUOhxbSACxrpNI/GLQGEn
CWtLe0IH/x324w/PclQ4r9OpywWun9vkewpg2whUffm4133XSBYpQIr+CEviNLawoqOk3bi05gov
uhzpXJ2gACyGccZsDBoQD4t+6OKcKrVNagKkSQoiuKg9OS8cLtkbnC1/DuP10T0RfB7uFcRtAhU9
Mi5LtoQ1FGdmA2Q53eYhg97HWn38GLO8008WKzhSERDKo8G6vFDp2bbd2loytS6yuieBTvMhWuS7
XCMES3K3sFCc0VotrjKmBmgPtfTzobKTdiExLi4bYiucjrVBOVssAunos2HzyiESxvABQ0+pQc62
xlYuMF2Y2t7hC6kz3IEC5gQixIzKwDH4GzHj395NW9ALGl7VP5H7qFhjDdqfAmNMCuWAwrihanLW
3cPjkIXpHwh3NZtVib+uFY5g+G5Cl7QmWcD2VefI17B574CKr3+uRWolKY2WLgEDlGcbnh4wr0/5
ar6j2ypFMGtq/orWa3lKim/XX3Z9GDliuzfTIJY0rvEwly/nHl/+syY+eGGm3M9fNG9kCGRaJ7nz
D03dDuwy0cIVeR1MeFLIIQpKqMifr57LAn7JUjbP7qAgfPoyHf5PfJrsKWtsOiOk0Xa4o8UtvwJr
K1vlSI1HrUjjYo++YN+qbaq6dBztRSt4k2jfFhvhf0aE51Ue63Z1/HA+fIKq32aLOcIF/RAttGvZ
5ypBA1hrxnRfBPtS5RCPqhtsTxESfe8ji57v202xIg/Oo2MErRQxcRu5uuIgFplaaIjUHr+Duo03
+3mn/TpmCEV5XlBhAbsOxY9FYpv+xfx2l9Y6JQGChvJWK9bZdf3693AP8wqWopAekSd9oTw6SZhh
XJ5p0Z4p0niCLNHQR9TJ2o/4FtHW3qQRmwXEtg/Zn9eQ4NJDRq4+BgsLBH53n6pggVLF7FKDyS1b
EGsp8mcRjKTHOTkx/tNOYGyg5LmsRzAhjCVnpUj1zOlmr9Gdtha63GFfkG0Q09nya2l4Ar1eRcMb
z8W589nXzn0+Bv2Kz0VjLoZ1G9GapoidvYybqtiXPeJsycNd/w675N8BpOebZ/gvrm3L1t1zfmk5
kyAQ8ukuCbO4O/3wTdhnz7juOwkRpjMTOtaQsne/7Sbd4vhKMu+oyqJetQueQuCd4lTkZqlgM8FC
lKhdrXdilRFuzxg+YNac9PQEmMSc6OTquUG6cliaz+gRrsc9C3zSGtEssgLNdEE6Rwffvs/tN/x9
1iDYSM0ZF+0gjzAueO/TFzvw6EeG6QtXZzBZ/wHyP0BihYv26NE+eow6nJUqSEWYh38yjOn4u7TI
28JqyqIu5GVSh88YlHgzFzdV8ptViYVtrYzMWWs+XsksU7CY5eu0lC9G7AEEnLxW1aOp0EHUFPRS
/mWhPj8Kwdes1xriguEBt7F0yirkXjGkXgNjxzyE6TUXch+zDgvixFkZMHXrfZ3pPSu1YwlvefDx
68/18Xdzx0LBnwKQA81QPXFMXY9OjFiumu9QSW4K2gcc3NgEL70BPA9u3eD9m0UusjFUt5VPpz9z
MVUqqyd0+xOGx5ApiwvCUKEqVwhiB/ZIeC46nLuumw5WYbSqvrwc56BrfSYPlIQizU3cycqEBZeO
5RsBNBF54AEO+YyOxZH+jHEtVrqkicQIovxe4wju96IvKLwVg12YJVHaHuGS1HU5Rq7BH8Vlplsn
KCFIq5YEdcasP+upbQr0Hzo7CCMG3VVpLlAz6Bvlv+jibCuPeCo40POxY1RLDS4+WTh/ac/f3BjY
YWecSHKNIDhWYr6yN/350dUM+9w3xqDFhYxUoH+7IgM/Y6sk8kLl/GlYLoD+27a4V3HR4/EzwViL
sIORxKUGEUZveB26ttBZSSRjzHURMLXnTI2KCHL316oFP+1TIcplN8NE8CGVM4K1l64JP0NXa0EB
TiEZCaUaf/FxIZ+e6oe+rTY6L19pVkZhrofkGe/Jbx5OdhcVdiaOXaghTU1y1pxDKFPwVVlgcX+X
E1HJ+Tx/+5IJThk+/uwEBvpxoHAhQnSbqN0zQT3cYZo73R+5/ZAwwE0D3n5ZJu3fvJ2vn2KOHpMs
Y+sA70GltXUjbor7CN68zYZwbYvagqwBXUWe07qALgMmkP5RplQnqKOpM5MWPjXzgIFlEs1OKFbM
QvRlA0iU4Ajvu3cwrZdxloniAFt46kvRr3YV7h4/XvBH5jerE/XLvavV4I8Hj2iS9zRMiP2UiScu
CVnOqGeEgmFbH8kZb/3/Tf/QPdeP28SY/rE/z3kK7VHKzeLMjjuIP6FJ+/qsY0+JDjlqL6Dxj0iD
NuMv9mba7464O5Muldt5/AMi/n8YoMJOiDF36CtW8sZYsVOIUcSJSIJlO7E7W+cIPqE53bsYESVT
ywynTzpcEKb+Gb8aEkYZM2AbeYtMhfNeqykK3KLUw8nDVi142FB0WBoNyTuNE7gQZrWIYaGtnYrP
5keRG1n76jbU+CyOHD73YJKB3pmXz7DoILDOZyYIkdXaj0QEWNUd2RkHBwlpdiqKWhtV3ueb3daa
aJJbhMlCyWdmjWbnkVurFkq5sLnfxeN575Wbq4QM2cxw7FVfiXIlTOSr0w9lvZaM1/jSwV1YOW1R
2iI7mVGyDiTdFNxcI1WqchE6X+TBvrhnHCd46Dru8/QTsCfCi6QYEq+IdQZIOTOHS8WKnpV2DcDV
hYOOyHWn/PrVso18AP5P7xpryYfi0yzHhGhc8J/JyQnsViK6UOjkxOC7aak+MYc0/KLuqVCNIcCi
hM1oCvEJN/AVVLGuWwMNhC/PBCk/7Xl9Z30QQ+4UJG1T63pYNEb/eLzUIfSlAGQ3G/UFb1VpzgVJ
suLGizEoo5xuhsKGASjZJlFgaMnW7erp+fnIXW7RmTW8PD4yA0pvwt3fEbgalmKGB2D8aJAkcqhP
e+gsXIIc6aZAnp7XMghM0TxX4JvyqtUutAHt+s1lZqO/yTpgJ5JbkjZR5y8GW0MinUvj3GvsyTb2
mw8d0vr0GnV1jR40H3U8QgFIvabstCewQSRr4iJ9YH5LEfGw4xKIZWZXyoe0nsGNcEAzjzNlr7Pf
RvlPcv37sVtC/LtA/1VFh4mb/+5cN3mzQWZS+eXOxE/8CvyOvdjlqHcCXRjCR9+4WC4wjGDxGjnF
SJJrCVEwWwSpzXnFpQpXQSyNLpvLPJfFdSBIbhUQqE0qdXpvpWRkxVytOXJQMCW1I41RxHTm1Gb3
SvyVJWk4qJ6lcGgZTJMFAQuXuDROvay+tyPvqtoa2Elsooea9FnTw4/Ekc8zMEie0jVex8ULf5cE
A0adhFlwcNRpfWVRB/g+9XLBFBBgKj6M2Utk/pmLnhFQrj4+jDlHmj6YfI6R1jgUCe5jZF2Afjml
imAfAwWHzUIR1y5Ce1p1DZPnk71R1AZayJBJinVcomGahU5iYSnfW0BNjDwcUZTz4IxOvDnnvnFM
NcKGEZRvtAXKF7I3dP+BMY4RUiBsS/nImfSWFjx0ardIu4Lcg0NzYKug+kcAwTd/1oeuOIrasa+3
3TpFSt8IoJf1nvnz+zFAmTQ+mlgWMMECvo4/QvDTSoSgGGtlcMKB7O4m1647Azmn7acM/q3G3VaQ
lDUg5YYXzN44tj77o4wplSaNiV6IDkAyu9uQnUUGfqbwldtwvsiIicAutdDNR8UbarkOOXcmUGGX
BHR1ZPc3/6ePrVzvzxi/2agDGvZ18Zwt0utsIYdECpFe/YmA9PM8PBhjbazVpHP5B7Yial/XZLY9
nnbXnEeBMx1XaSBYAnhWj75zbd23WGmJ8O+1WjWID5IVoV4U/VbBQrEzaqOS0WB5AqUqCuRI8s3h
ZJLQAX1LznOAZtQxhqS7Yd/adzElTP/DJUjhA2dXF1drElYL7HVn8xSeOyCvoFUk+Uj6ufgTnGan
mV0jiYRjCPPkrDjUO7VpJEuNfha86KSRejN6Kt+EaTcdYyp4VJ5X+xgKrljCGtOXtBVnCy4Ycll4
vlJn95IGnFI+4h8C6+0ZzaDKTRQF3ijFmtNNcSkoK8LEF6YvEeVh914uzN5DMe7F80coDxLhlAPZ
FzfGd6wBNPTjNlG7K5W3347N1RmQnwD/fQZOB3oPfxHf3Tm+E1DN4ubzA57DBDt07XPYTqQzF9Hp
q53+GkVfrvi0mLn6jt9kWJ+yyyY4cSSpH/ABYzJSEsZ8QNfR2AQBM9N1oPA3o+nCa2i3HPaSh7KI
VQ0cnVH1w/FT6Xa+0Y7hSCuf53rP6Wj5WsXD4HpO0DaNvx/O0lqmA54o2chNGvy36Y9UCEfd16xu
PQnZWcV03i8blP6rf61WIMSwUf6Xgai5oSdTMf8ZcA6EBRYVX3b3+WNzowHfo23bFXiQpojG+wd3
5SKudgg4REZISkwGLMnt3aFwl/t+Zp1Zj/jCUkHVAV3cRPKdF/DAIQulKXdSeNUZZzLXwkiRlTyU
jwqWQ8tcdmQLH3jKZWFMrul4tygGau646AYzqig1IoeJ/5UbidfEWSU2Y/eHZK7/kfd8I1ONAt+3
9/O2p5CS2MlpqS3B0XUn7HvOhKgGD7NCGj+XIQRBpFCI90DjbQJazKfRQ7G2lBg+cQK1TfXKw8Mi
0tTGFl0HEf4I7icy9no5IHZ6YdOvARESA/GuglI5oKsa0Q0XP/qsBimsuKGMVuvjt/Yys5QJIdVo
tP2lM6YSrb+VOubi0npqhb1PwNUBzvP0YGLvhCCtjy4FbFN+eiitkRQiWlElTM7EgpXdZ2NLxK7b
o6JVLcFpeilCrR3DIAjlb98lhh+cfgrDFoX4nm5831khJGtq+veO2t8FNSITLU3U/FHu73Gf5Dix
y3D0Y6tNZZsjb1YMRDougQRD9astl+/MK2hsvoEn6r5htGDWCOPAZG/HT5gXeghHbpQy910Wj2YE
mTApcLgjCl03XlUxI5jUEzq602tdwYP72CilQWcgjs+sgUabecJSJg6+etixm5sDCCgMmDKoauvO
/Ii5NKhW2VxFrUPNN2Pfkh6LZC0u3YgmCPmntHKLNY/QOuQlAzNAt0uMG1E4qPXaq+Dz0Jx/f/Ex
G+tc3sYS21mhrxOyoiqFD/X+nG7qbB+63GCXyA0HwNg7dhIHtZU7zJUlOUU6Eg7bUF/8KO4TwEfe
MgTDi2LQnbw0K4NBn682lqrDlyiUXH51taemMD5qa75RnfjduphxfTMebX1Fw2R1FOMHDxHs/mbf
SQc2eQIUgHiIfYknjaMTbzfNhLt0wYTskvClksdZ1xcN/VidjDoneAoqmlVnLqc2dOB75XwrJ0AD
P9IlXrbBP5DvRAYgOP58rTeJgqUXQDDqdZnuHvfrOGmhPb1Ni7EKpXLGJJF/rQ==
`protect end_protected
