XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��?R��+��Tv�Љ1�J!34�w��8�Z�k�M�Z�푫p�5S�EM��!��l�'�2{}D��Ѷ>va���,DH�1�&��y��<�$#4��d�
��VA�޿��&t-*�l�c�����H�
�T�1,Ѣ�߭].�����1PZ���;��&%�:XW����+�2J*pR��!���Cw�&�}�E���ĭ>�!���\��B/��Q�wU���_u�5M����;Lhq�.l9�#;�����ze��N��=sv���PXS�d�H�S��� �T�Ș�
��F�'�Ԗ���,]t��z]fq�+���5�	��@m�k5g��aF�IjA���؅L��l����j=���?]vpkq��[(�)�G���Z���P�lQ4e�.��S���I�����a(P����=�
�(����ܯ�.�t�XYU��,`2�pҒҔ�:Sz4�}�5��"���b�.��|W�[�zy��
�n9N� Ό���E�ǃ�
"V}�7Ł�k���_�$��o�����ڼm(�o����Ϸ��e*~Bz��D"��^G}�+�����a�>�F��ASˎ��,�j���/�"qGC��	p�ne�F�7�LR �>��x�پ��'�!/�)ȏ�KqࠖsJc�Xz?�wV1�9gW� /�`��`�qo��w�d��q�1&�"�J��~�� ��a�Y!�;�(�CGw(&���C�C�{J�J�����(�Y���̱(��#"���^р=H��XlxVHYEB     400     1e0�j��%��V�ԉ�Jl�T���c��_8"Mԗ9�+�,0ns�@�$��(L��<a�	%���̘w~�z��3��lܪg�If2���a��b%��o��ñ٬Q%�)��^�E�˂t0��c�IWX��{*��`�գ��օ(��٭��j��F����m�� �������H�r�$Ptv���2���ى�r8���1V ��b���p��W�
�ydj[$9U�ЇE%��i��tw	�klש�gJ[_��}��LJʲ;jB�E#��{��ơ���2G���.�}����M��*[����k�*@ 7��ߺ�t�H����y��}@�����2��\T�ZX�ۏ���ה�hՋcC%@P%Cf���F��&���	��&��/�Ki&M|:�œ8���j�Άhg#�1њ�����y�z �C�q��'|�fP:Ҝu�=~a��zi'/L���djט�dux�<�>���XlxVHYEB     400     130�C���4�o��?{�S�ԯF�Dm�����z�<"��&W�	q�7�����RxW���gKWve(_�nY�o�J�I�+���زq	��%���5��er!H������?��QA��V���lx,R8�&y��
�W�Sw���/
f��`�J�6�B�Lt\e�,���G���J�'a�(Z�o���2�'�Ъ�2��ltO���i:���[q�x�J�U�ٹ�q�2g_H�w����į8zm&I�����+���ff(����_��LUt���$N�V��f��o��]:Whs5��;`��z>7�>qXlxVHYEB     400      e0C;;7<3���C �}�?�x���7Pg�N�H��Q����.�)�s�3|6;d�)�ns��}�vz�08y��	���wp���{�:����ф*|!W}��`��W�eH|�È\����a�����]c���-��&=����v+��Ioy�]C��_w����b$J�R���ŕr�N-�<sR�|�Q�=����i��H��(�6���%�?�A�Ƌو�XlxVHYEB     400      e0'с4V�ͽ�o��h��I���K�ڟt7�G�C˅4�^hq��Y^��lB ����$�����<�x�2J�(��"�M��z�q��2#���ן!xExyK祮�����U�B4qEx�1�$���E��K$���Ɨ	K��@��P�\�SG���*�i�'��OH~~� ���^��9d��o_䟡p���=�� ��~�S	�&������ӥ���zI&XlxVHYEB     400      e0�|��p�<IQ��Y�:)��=4L���Ջ�)�H��2� U�nQT�ZC�|���E�X�7�#�_����g�n^P�򆁨`����k��[ڨ�R�S ���֓����6m���ΖARx����\FI��K�/�P&����Hs�2ߓ\M�V��	JmX���p�}��*)�ݚ>k-�J�n��>yL�$]��2o}I� ��cϯU'��R�L5-YP��w�NEC XlxVHYEB     400      e0خK�0��[���^�^2".��Ό�7[�V�GE���KX1n���9M&I�%�&�6�ĩiӝ
`��e�7�4*Ծ�>�P��Pٵ���Q�j��S���+2��R',��~�LV����M���?��g��_eH/X&���.U�U�>5�фXF�P���Щz��t�n����n�)A�ĕ$����/�--�u[�L��˽�/D�>��ޟ_�������XlxVHYEB     400      e0ax?�i���9�"�I���+J}�KSˎL`��'��F;/��}�-}HC_yH�Z�/�*��[&��|gI�ƅi?(��H�����ṄT.��,}��UBo���X��(��IR�>Y�zA�+�ιt�A,v��l�v���Y�3O��Df3~
�_F���q��g��g�Z�i�K!e��z#Y/�v!򽷵_��gjťE}�\c2p�OA�xRϠ3[�᪑۲�XlxVHYEB     400      e0��f�6�R_}%�Ji�����&��+����z�L�Vsm��<�P�H�v����R,�����\qV`@t���#�4-Ҭ�!MNQm/׿_�)H���v�N ��w�	���O1��";��L�����!�X��79�[{�z��y�0}6�͘�9��s��xJ�!�����Y^�Ȳ�db�\���B	&��FTR:��!������lߛ_�XlxVHYEB     400     1a0).��ֈ#Jz<��(}��|��va��'ҧTk�j�_	�]����/��m��{��jж��صK{#�ـ^db٬��=~j�Q�V�h�?�u�"q\���N%��*��ն�6ڿ�2v䙏�٠�t��?=��Ox�3��g�3�^1�QH�c�\����/�eC�����U��g-�� sH˱���T]@�����ʏ����L�M;�A�ћ�~�~���\��U�%�OLz>n�i*F!2��9a��~MH��q��;�,Y���:Lt���C'�T�?l1 �i�����6�^�Q��yY�����m_�}�Ɲ	d�s#P֋O�yk�h�J�7��DM���79S��=g�!Х$�K2z2l��'�*2K�P�خ����{@&1�d�;�@�>��l������Ӽq���A�1n�XlxVHYEB     400     110��/�5��y�
��2�z��N@����e���?"K�t*C	sQZHnQ�?j���\k_�z޼�����XXz��D4h�7�M4*X��l%�[�������V��#�pP�ː9av���S�������<vjl6Ty���tm�&��J�����/(�=������
4�K�b\�yWH�5�JD�uC���<\y3X��x@�9.�
#�
�f,@�$����u�;:6&�-t��GZR<nͻx6��������B�[~T�),¯�ς#�-� ��M�7�XlxVHYEB     400     180�íٽ?O�K�<ѯ��Z#M,\Tqr|p	T,9�jGzgW>��hH��\�nB�#N����q�G�p�{p�&����n[������7g[�g�ע��G���o��ߊ��$|�N����P�ze�q�^����Κ�J��� /��j۽C��+�#��*@���ͨ�/N6Wpk?cӼe:M��㕎�ysVZ\�I����/��u���󽼒/�'�00��M�wl�����G��	���#�6G�_─�[�Lƹ��p�y���F �Ġ�	�ܓ�y��7rAX=�Ҹ]�T��p��N) %��7/���v�X�&�wM���ν[���^r���a��Q�PmM�^eZz
�p��_Z�'�c�q��SXlxVHYEB     400     120"��t�J9;L%={�7B�������&v��zC�1���	�5��;7�oV����B�E&�d�q��M��n:�v4�;$o��f#�Re���|P���]��q|j��`��	$�tN��WiH��I�Y>�W-��=��2���0:wٵn�
4Z+�ܜ/QΣ�|۾~���]�R;�K,S�7%e�O��Z������rڍ��e5X쑕���&���CV,+�I�`�uzS�����?i��9y���cS�Ҥ���������#ϝ�%+^�y_ޝ}�XlxVHYEB     400     130���*���e�D5h)ڵ�E��Ɓ%s��A����R��Z�;x���?/�	�w7��]U5v�<�,[�.l�`��'Mz�ħ�0ю�:��?��MUa�����D������H��a�4��򇇝�)T�[��`��.@Ԣ	�o��)N��'�\l����ro����X�Trxk�ν_�D]I�x_n��� ��������l���dCb,1�C���c��$�9ø$�6����3F��·�Kbs�cKf�]�7&�n�#����1�֬��g���
b���~#rc����/��G3CEh3oXlxVHYEB     400     120�e���0����d�f��	2�l)�o�]7����='-��f���������Fk.�����PD��� ��B���{RT��,�ƀI��mH���Q�בj�8c�I�BJ���'���a��ʨ([:�r,+ �C����[ć2��2r��	<����f0����&a�T�h����:�.������������.Q��p����M���'w11}I�_��e!��d2��`H!yɦD��"�����څ�(���m�&������d�Ƃ�����3R�XlxVHYEB     400     140YJ�♓���	�����?�2�+�ST�v�r����3/�K��?o9��7��t���u)��iLmq�I����2�D�:	��wg?��e�x��y�U��E��0�Ě\!�p,�&�_��'$"[�q�����^�?�+n�)RA�	�'N��d�@���.��.x���D~�,�n��_�ߦv�B�mm��UH���%<@���쬱�� �$w+yQ7��GK#JT�q2���C�|��!襤���.t���0�H��A�?w�&�&���?<%w���b�����RMil�������ϋ1�;�p2�*x�3�XlxVHYEB     400     140��@�&��j�m��Ζ�S��r��8�s�&@Ä�4�g��ƾr�I�I� ���o��b�+����� D�x*�O���*��i�\]Ӈr��_l����L��7? �%�C��I����+f���gb]��(7�̶�m�U�J�F<�T�[w�>p��BbKB�KݍSCt`�0@~���lV� ������S9/�7�#q������Q	���h-�����[�㨏�R�T�9�S���3.rn��D�l���m���}ᐪ�L���|�N�C��a�ER���|T&�r `�ʣ��0-�z�
�XA[%�4XlxVHYEB     400     120%g�[xN�u�3�^c\�E�s�s�6����ad%�w]'�4���������Jh�ZGoH�0��\��b�??���%��	]�p;�"+�1{x��!��1�e8Z��e�-�(�\9�4����	���;匚��7gц� +����3%��W8�4�6}4�Y_:\��v�B�NT7��[,��Y��J��ɘK�5ūA�z~i�8�~���r�k�Uj^� 'M��Bv��$��o*��p|�/�*8V ���#ue�n����Un,+���������gw(��P�ͬ4�?���XlxVHYEB     400     140Z�]�.��0�R��X��Ǩ6�mQ/7��|��)�k��O��U2��`#O<�����Pb@6"=��)׊gz�9���Q��'2���~[	vp��C^�����cD�ٿ�ԯ��yӚ���ƍ�ɯ�C��tO���"���Q���Xzg�[�mi�+�;e��&���o���(π�P�a�kC|����{3�{%�n��y{=Mg�-�層��@�d��r��Nr�/l#�u�^��Zx'S���OK66��H��d���������+�?�=�r��@/6n݃'��ę\M
'�.��� �\x�A��XlxVHYEB     400     120�ЅZnF�98;���������!82�l+�
�Ȣ�^lY�mG��)/�ѻ��~�P�םJs���\;j�/xMtQ\���G�b)���𔈆�$�@Eo:i�1cE�{��4)ڥ��`m
"�]҃��1�����m��Tz��,��u�����rx�����gI>�=�D��,>WS�l-_L�G�!<Ʉ�l�BwH$]b���N�r����3?�\�dܐr�w�EvT��O��增����n�?�����6���Jq�@`]Ė�wH3iLAY�z���*�'}wd��l�Z|ș��XlxVHYEB     400     130�|�2���{=mZ#˔�^6=f��SH�gR�U�~�4�?�3�Z��1�"Gؾ�"��6��+���fY���l�:�0b��|���h����Nw�n#��'&��ϗ�jZ�B}��t:t"���Q^��}��4����uD�t�L'�i��3��9��E(�Nu�<���l����BDQ��v��(�r{����o�n�pھN�����bY��TS�a6I��-��D2YN\��$��^YV�}�7f�3ܴ��O�+���T�9�i!S����(�����Ll櫲���.sAџ��g��OZԦ&��XlxVHYEB     400     120�@����)��`�����)�:)��m������d=}L��fo�^�J���A:��3���*~Ҡ�$��S�(�3��*{E��sjڮZ�kJֶ��sS�qSDK_��=�23�N9�K��୐{�v�,&���n����p�R������X|ρ%�&����VMѶ���D�Զ\P	r�)mK�;��Sxz�wM�1�O� PӞxj��j�u"�q_]�eëj{��C
 ~
��H�����Ǆ��,��iE&�A�����z�����fg�<�S�slr��8�Q�XlxVHYEB     400     140a�����)�
��r�d � �J_"0�-f�>������}s6%��}�Ȅ?4�����a5�*�-2�	Ϛ�C� ��Y�@q�s�ڑˌ��ҭ�(XΒ;�,m�#(��b�ʾ$��z�<<�%��ȦD�=� �Pf�Q�������Xwc�)%]K`=jb�G̣rE&���M�=�V���G�_3F�)�e��	}���{|�7v�	�L�!�x.�Tӈg��7�q���%6`2�vGiMO6�{�pZXd���k:=���B�_���Л��t�j+��&��E{�d�ҧC�+�&�v47�MJ�*`"a:I�XlxVHYEB     400     140��@�&��j�m��Ζ�k��&���s4�����#7��Նp�l��=��^�Z�����d5��
l{y��_�k�B *L�Ρ|�,�"�i����4V-V����|�C/���G�ŗ���5Q	���zR���9�L�vtS2�%�4�.[��m�)�Q�&)}Ee?L��Ž����|]�j��:-�.�����e"+��X`=N��g+�c;"��uQ�~�-��zǚ$�Qc��ϫ��߽q�?jZN�hĥ��^�}q��"_�}T��t�"急J�R,?J��qK�i������1�㉦wq���CT��V�PH��s�XlxVHYEB     400     120��[�bzK޽Ixk1�(B��D���5���0�]�N��$�Ͱ�� ���3s��
3����t!�'fW2 ����S��d�a�����e+�)��Hƣ~]'e;�V\e�5���=d��@� {��gG�챧�1�S��:��ꕵ������
�%���ƨ����kϟ��X'�_�>������.�F��y�L԰~�7�0JdeK�P����?n 79��q�9��-7����`ՠT,K4 ���[�	%��R:��sۓ�>�#_�é��XlxVHYEB     400     140��������:��,����b�|=++��i�"����QJi��2���ϫ�+�}}Ԝu�1LE�k�b萵,͑��9���N0�ȓW
��L�����[�˺&J8�N��`��S��m��@s���P����	/�mȢ�WL�G�&7�w�9bn�]�n�a�f6+{�[Nh� ��Id��y��Fdpil.;߿�N�+ ��Bz���������@�u��V�;3�@O�(���\�j,�bVO�{efo�}�I]�_�l��W����3mu�O}�q�"�n�_3A���f�Y������.�U�%�T�cWZ��06}V켷�hXlxVHYEB     400     120�ЅZnF�98;�����*�%��F%k���h���	��gC���>��t[|��A?W04�n^�ޣ�&'����W�AJ�'�@�h
4ѯ�eY&%�_Z��>!�G�2����1Х�Z_�7��pKJ�ޗW[Ԛ�&�����Vqh��s7�:ѹ勵�8�1?�A	�+��܀H&�캆e6�8��آIrP�[_��y���ֱ�! ���.��iu�)R��{��ZѶ4q�h;STEA7�һ�nm���Qv��s\�WX��?�;k���((@V��@�X�z4�|Krh�f��sXlxVHYEB     400     1304u�^z��h�G5�7�~�]��kOu���nL��ô�5i2A�~
R��CF�^B���8�-<�$ݯqZB�R�4�!��&7�WA2�g��ILc����{�x�R:㝨�e��|��8�5D�,Qt ��"���W��A�YGO�ϐ)(7�ɤ��0�LF�`�f�������T��a��2���n��4�q�GE���O�P��bD}�Q�G�����[}�uo��Cd
&�w�=�_��t�
��S�X�,���4i���=�Vʩa�z%���8V�~�d��v	@�Z_(�դXlxVHYEB     400     130��U		����{o>[h�.�^����^Io�*�KJ%˱�l_Mg��`Giג�6�F*��x*�Nμ^%�Z:ٗ���T �j�&8�I0Ŷ��<b�U���B��2+ǀ�(��� 0:e�v�T��A�J�E��ӆW���L�~�p����t���WszPO���i1W�b[��>2�$j��7ߒj~�c�QČQ�Ut�zo!���ѐL��b��G����K^�M��B{��J��ׯ�P��&;�4�9u&� 9��ܬ��oa1GL�@7IlkKo&,��;O��>w���XlxVHYEB     400     140�\�3z,��!H���0X���
ֆ�*�b"B��=x�^��m�7��\=��@H1m�9~��������'�Ҁ�'�'�<����~��͡
�G,�葖�sZVI0�c��S�wD.�p����������|��b�jSQ�$c��̓�u��3T?a��J����sD��p'�X�o�6��g4��}Z8���e6�N['7��o}��#�/?	�&�������nD��b�h���P�c�J��+Qt[wCԖѡA� $ٍ ��b� q�����Q]F��Kq���ah�����b� =����l��KvQ�//)���XlxVHYEB     400     150��@�&��j�m��Ζ��C�#.Zm�V������������Z� mo��n����8�hl W~\�Ĕefg,Q���P���	�-&~s}�mb�bz��BIo)zj|��f���6ݸ����#���N@�
��Kh<y�	F����$��o�� /�&z�V��:�}Y0N� zCI9P6����C+�J~��	2_�qC\��n��אU�0�ڱi�y�Q�:��I\�����j���4�����˷Z�t�pm�TT��Qz����fW�d/��{��G� ޛ�ECJ���Ut��-/��G��X��s���=����NN n�]ފ;�XlxVHYEB     400     120>���e/���4a�C��ޟ�Nz�S�ғd�j�6�4��v���!�4JV�ܢ�/^�( L���12��t��ɀ�	_L(g̤A�D�6��	���զ���^�'�Ë��h�,{�6P��2pw�������Zn��ZuP�a^�cj�
�T��p�O�t�m�����P�B��@���s�Jh�f�T��������a포�&U�Ւ�9����gbok�>&[� <k�d"n	 �dm�r��QR���a�[�X�n'WJIϪ,�ta/�7`tx�%�trXlxVHYEB     400     140��P�%]V�W�� ���1��z ��̨ߪ���~oң���T���Gx�m�ƕNJ�Y�@��=Zs��*[� zT�#L�?��i�]�+�4�Z�Ν3f�o-��S�6��	 �S��INy�mKP,�'�XRu ����@��ħ�hZ�2(m� zJ�����z���T�|A��E�=GF�wS�7H��r)�=֡�S���-i�M��2�%��ٲQ	\��F�%��`o�t�,C6gbQ�gj ^�NF2j|F=!�s{~�HCOE6:���O#�}�dFe�  H������7�|������g�U���IfhF�1!XlxVHYEB     400     120�`��ͱ^G	PD�<�]�)Z\z��X�hM>��ХW�ǁ�-O�*��d5��&\=`�h�z��=Q�h��f���%`C {}J=;\^�/�zHl[�:���	D_�IZ�C� 6G��0e���7ϲ��t!\?��f=�U���eV��gig��[s�G(��`i�L;�e���a~�˝1��rX�=(���D�la��8��>L��Wg�����	��Dz��p�ޕ"*AIu(�)3�1��cpF��h���|�gy?����@��@v�0�0\�	~�!X�J �XlxVHYEB     400     130�|�2���{=mZ#˔�^E�>�0�K�G�-��`T��饁�٤by�0;ᗗ1I�e�����u�ͤ�6����b�\&.����,v�j7��>��@�4�P��2�J��UN{�@�.�`>z�*AȈQf�x4'Ӿ�/���ڳ�߭=KO"x���3��Z�4&�H9b6�����1�]jUR���Ш�>$|� ����5�qp���+��gf��=����|�tX�fs���R#�ʿ��&��y��O�����Cuf`�4`ď� �H�Y�H��gh���b�6\�9\XlxVHYEB     400     130��U		����{o>^	zJ��C[���	[�Q�)�Q��0r�*�!晼m�H�k("�Nx?��������x���X�������e��Z�@�IE8N�-��ڊ�Jϕg��
��6�O�VY�X������Y���L`��uъl�)<�,�R�*=��:��r���.$g+Ƴp>T�R"�f��N�E��?����|0poš1"���Q��X 
�YV8�D����eȺ�m���B�D~�Ɇ��X� tX4��pQ���z$���It D����$�!�a˳LRd[�$��XlxVHYEB     400     140p��G
�1�&��z��$}�nT/%Ҝ}��5��-�U�����d�Q4�<���d�ZHD�V��#I0�VZU`��"U���C��bڊ��{�
�����S�T�e����6�J��D��h��H@zq��+�K�h��
�Ys�5^v�8ʙ�#(2m�i9�i]���mIbe�D{�?��[������כ�i$չ�P�8������A�'��JH��b��n�vE��g@�^�D��Dt�Qy����R�a
}�ڸ��� _�g�<�j�7�D�́��`�K��U�$���x��ފ�>��/�u�������N���XlxVHYEB     400     150��@�&��j�m��Ζ��}����k'1|�/ڪt����#��-��J�2��[N��1k�dr��}|3��+�ft;h�t�8�YHXp�ah�9���>�dAN�;�)��׾h4�F\ ��w-�Њ��.��o���I-V�YxI����ƱT���C��n�?�?�N.|��)�Nn���k�\'[�ܿUY^]����^���U�c�����tBv���� �֒J-R��]z�o�����_c?��[�l��+\��e�4�h4��y�Vw�(J��k��Kd�jɢ8�;�Q��S�L����rܢ���x0q�����:)�g�D�`5{B]�w�6ޯ��XlxVHYEB     400     110�2���Q��6(C���ܸ��
ۍ�Hsq�:f�Q�k���z<E�N�px9h�ƛK�2�B��^D�e�y�q\�hL '�u:^�1^61��|Zp�,�*��FTb �p;	��Σ��M�� ����BG�
�X�Z���@w�{y'"��2��+���<|DH�]ґ���h:¸,M���"zp��W���;8�Kg�y�Qj�D=�{�����88o�+����0j�P��G�(��g*+7�������k�0���_R�����c���XlxVHYEB     400     140*N���R��By������X^v~�_�y�_�V�IY�Ǭsq�Z�M�XpV��^_�Ep�Z�A+K���9��e'h3���~i�h�
�hǋ���aR
?!�2����bд#�?_9m"�9�1`�����!��骐�d]݇<h;]��U��ui�m���8am!åb.�(���»����S5��G�J	���ߍ;��
q�1����J�JI�~�cA�3Wi�8=VT��=e=I�9�� ����t���?�>�;w�2[%�	�
��_��ƛ�>�V�y��{G�����4�}0s~�#�'O�XlxVHYEB     400     120�ЅZnF�98;�����t��!�6@ڳXzw=~[o_����3{�f�g#��d�H�L�n��kz����U����.j�=J�~�}��n;
�^*>���E�ġ�j�.��P킑� mN1��rbt�1h
���!]�>iE�׿`?�����h$�bH S5�iy��Ţ�i��v}�\�[�4XK&dN� �9�џcgS�I+�T�<1bVe���#�j�������U���yX븦�S���s5ȮY"1Ȳ�Kmk��ߌ�XSzEEk���:��>�+�S��)XlxVHYEB     400     130�ˆ8<����9|L�����f�{'8d$�-eص�Ϯ�]G�m�p�b�
���&�	�Ce�.�Q������
�U��ں&J�G�L�K�[�Me�O4���6k�~���8	�mK �}���8ɂ��`�|g��(q��%8��ש��7�:�'�F6`�����}�NW�ց�d� .�_ùz����*:׀�~|��ˇ�V�o��fm�]Em*��y�3g�s�j-��pC.˜p��J�r�}$�Ji7��ɞ����b*��=��ѫ<��jm$&�ڃш�0~4���;�%K��������{��Tu���2�XlxVHYEB     400     130�� h��87�-uǒOC"��>G��/n.e�;��L.~�Z3_��b�cEz����Y9������I��I�T
A�����.����^���W���;�eg�Z��o>X��G�r1ځ�)8_�g��[���e����y�Ek���<��-P�z�-�-��F�WAr5"͌۰�:�ׂ/���i��/��6�'�������ֲ]��A�q'K�E�O����J�{�}�
%��L� ØZd)��A���z]���|b��y����d�K��x�0�p$�7��
@������XlxVHYEB     400     140�_%KT�[M*t��U��?f ��i�|G��������Y;`Y;G��R�qm/���8��8�ܸR���L
��L����g��l9��K>��k"IR~*�4`���۔���҄|v�HY-xvb�o��dC6>�vߨ����AK���~1��2�� �ivE~s��p%��k�"��G5l���~��K���[��C�/<�A�
h8̉AS
}ʰ��T+b��Y�T���;��.\5H�x���օ��X�YK��}��^��B�������hG��?�ä��i>�&G"Y�>c3��Yq�72���`����}�o���.	�'����{��XlxVHYEB     400     160�n�I�o�W�@�/(��	|�V��uv/�VPI�Q8��蠩
��gg�u슧�;�)��ƃ6�L�6��2�_��Pǋ��S��e����|���������p=��SrB%ڏ��vk����;6O�M}��z��	�t=@5�8�Z?O���8&����TQ/�8��0��l�'!��Ơ������$��f�$/�i�1�~�u�a�KT�m\[mt+������D2Κ����8:�P`Ę6�����R�4n��5��l��4V�c�ǿێ���7�#�����鐜� }�L�d��,;6,�����b�ۅ(�;L�\��w�O6K�{ۇPP�7���o��b�XlxVHYEB     400     100�:{aPĨ۫=�b��̓;K@��P�f�Ԇ��25�6{[�~\sOR�����< �h�7�T<sf�ɲsg�y\��;zRk7#�חu�MU��O�]Z[�6<T��c���j?�mŲ���<ΊV,:��LB#�A�s��1��:�����D��Q��K��ub	���D��e�ǒzg���L�(��*P3���ui5�Y����Cܵl�b����$x^��PL,è�X�F8�/����߮�J��7>0XlxVHYEB     400     150�?v׳r��h��U�����j��ڪ��fܣ�;kb�;\:��J�/�F��e��Ho��5=��Q2Mm0�}��W�kosܱ��ޚZ"��(��QΔ��3_@�x��5��Ҏ�u��Qfb�����K,5�=�H6��8+)��f�T��Q�o���"��1�w��B}=�Uxq!��뱴�s��Tr���xo�xH&���=��� ț�	� ��K��N�,^p�$����x�{����� ���j��i<Y}�o��`�>x�N;o���R@"��C��`�tp\��z��hE��j9/;:I>P6�g��-��#. ��@�GB􎦯��%�~���Z�Y{XlxVHYEB     400     120X�?�~`�����a���f/7q���W�!at2��[Ug�`? �{=�{4 _'Ū9����GI���>�]��?��-^V�,�J�6󋗚N%V8:����(�s��n�΂��~��|r
S L�%>�`+>5�>�''9��7+ʔ?��*�����\GX392D飦�D-�Z��(4���y�~��|�+nS�h�����z�:T�	Tpݍ-m�f���v�i�]�Q��Ձ��0,r���M����dB8�K�j�[�fY�l�.l�XlxVHYEB     400     130�2���%I����Ǖ��O�v*�mY�wYj�e�b�Bd��%��5����L������h�̑چ�R���BB�Su�� �~�uW��#aųC�������j�X�~�� ]��u�m,�u����嘿�E��5��Z��-�BN��1O��\��(�<F����69�"#������#����#����W@�]c�3��Q�|���3Rr���3�; �,�1Yj���T�������5q
G_
��wz�G�C2�J��y��/�?hĶ$�8Ѓ� _�����&����,���Uƾ�=XlxVHYEB     400     120>��¼��պ=Q�%l��XO��lHG>P�%�Rk� �C��p��b����}M�M�Q�g<@�"�-�b��[�K�gF��u3,U�Tr�S
��r$��M-|�dq4��nH>�ȦM׏Ý.mx�6@��>���\���'�����΋a,/ضp#$��L�l�>��HX��$��;$�$�!�Ǥ�7���?Œp�,j�j΍.J�`Ʋ��N\��K��#�ո�\?Ek͆�IK‖92�5Hq_���>=0"�)$�#/�V�n�;��*$.XϿ�ʕ2��XlxVHYEB     400     140F;~���`x�j���1��Y�v���a�yz�R��E`2�9v�و�U5�������b��D�Xx��(U���P��Vq6O�L���V��W3Q��$�2�p��3hE<��:hN���8�xdKS�U�w��%MP��6�$ܐSi��vn����|/7����8�h��PP<�\yʱ}SҮ;��/դi
�:�bU���I�B�����ǉ��L�������	��� t��{#�Z�ȗ�tR9s�$� �̩�j����e� ݴ$�|W�����ʛ|�&����X�rE��<0�3�Dۅ1����cZ_��RfyѴ�a2PXlxVHYEB     400     140�y�a��DF2#�R��X��_.	: 6��7>���&7$b�mʞ��5��6ĥ�ܗ����u����c�X����X#x����ʤ5A(^����DX��!��Q���P;j/�o���B���F�Иf6k{E�T��~�3D�+A� _u&&{x��r��Ov��]��q�9�t��!��zG��IߖO�nvMt�0ZެL{�')��y6iSt���V+@�b:��iJ7P�y����ۺ��qq�D�l
�IM�G���KN�<�Sy��2c�Ҟ"��.s�����BO���D3Y!�M.';�wZf�EɃ�үCXlxVHYEB     400     120�i����}V����H����0!ӌl���,?��շ�����Z�����٫����b�N���W�#�[��*�o1иಈ-���7���x�e@,�W�j��:Zw�ʕ�e��=�X�F���]Ou���EIudl��χ�X�Y+��Bs�S����B�����:�V��bx���.���yHf�p�áf</��_sÎ#P}"�q� .xkTw؄�u�ws3�ZA����8���	[��"�x�YT�q:�c�[�s�n+���rlÔAE5%B��,h��݆�XlxVHYEB     400     140��g�m�/�BQY��d�tJ�x�wD�J�&�����cb��ֻ��_��[���;
�a��4<�� վ�1��`?dtw�'I�R[���<
�n�ภb���n�Q��j+�!�}_ū�Ą�����Y��K�_<��iRv�U�A-�B�� ���*W��r�ř({��]�!�����7��C�8�أ<�pߩ���3�k��=���z"<�g�K6�����q���|0��R��i�͠MՎ�R[�F"ؖ3��	�F�6ko�֋�G{�1��t�����#�׆�<��NQ���Q	ژ��*5:]#u�XlxVHYEB     400     130X�Ϗ�� ����v��@p�N	<�ˆ�1�,ѝ���#����+�8���ב}d���
��f\�/�Ivh��5:v�=�QOȢR�[)��8wAH���[���zXG�~)�O�H�|M�ፖ�i�9��]=���8�������7qá���h̜����#��2�< P�ȭZuq�⠅q���չ\�g[LX}7�w�4̼���ǌ/�__�V�$�n^��� ��V�l���:�ťR���N��Ŵ��0s�ō�m9�;y�:�֏0�,�t�����-U2I`��z�U�������@�K��"�`ߨ����XlxVHYEB     400     160��=���D�C$!�߰:�Vr�G�s�.:�EUt݅;ohg�k�K�����ݨ�w�q0Q�Թ�!��Z���O
҅�&���c��nަچ#�2QVVx�B��N���CIN��9̖?\y^h�M�/Y9l����|��ʇ(�]d�Wk����ЉT�Yf����spF`��C+W�(|�����{&w�&�X�����N�2d�j�g�������Z)�Qh�.s�`���C��d��a&���Ҍk�q���]���In�Q���(p���>���56J}r�Fת#i�,I�S���ǜ��_p7���f�$Dl�0x�,u���Y��h�VYʹ���-���*�J��.XlxVHYEB     400      e0?�4ly}���r��L?���f����86N@�w�LRg�c���4{+
�����v���\j�;�~.&ue�_1���3$*{S��\C�>t t�u}ɍ�Y�a�j�.u���˨����4��|�L��f�uE%��VHT¶*G�=-�E�q�����]3J��o��?�������^��VCa�������P�S�2p���;-���7m9U��oб�q�w�F��XlxVHYEB     400     150���yȂ���^����@���BZ`���lX��B&m�4�&ͅLHZ��ؼG&�6t�ϟ�!�Wx�L87���$�'��D���yi�m~$�G�	�_v_\M�1VEa��]n�m^[�|�9��S����M���z����{������iC/w�(����)�^����Տ&'g������P����x�":̺�x��p�[��Wg�B>�� ����5�t�B�˘D���)�dp�(;v�^��&�f(� ��`�j��fI7�9y�zҶ.�L��#���Q�L��_�_]���+�bBGD8�q�$'^�
'B�m�qÀnM�.��ߪ�XlxVHYEB     400     160Q�P��˒3@�$�A���9F�S�;���>�W,Iٺ��އ�j��$����M��+w��Q�� zCD��9��z�Iz`/e:���E睦I�u�_A�p����q��S�Jv#�hl>0w��'o��S��
�dř��N9�d�+�Mx����݇iv��8RvRؐ�� /
f��ڐ6��`�nkC $%]=����c�����S�g�f��s�s]R��yv�ϔㄞ��a4Z*:
���+f�1[�<���9�TH@�{��Ҟ-Q����%���'�!�vK�
r�C��;hz3�`��q�`὏K��j�@�QN��[.&`�<,�5v��Jw4�TU���Z5�v;}�8XlxVHYEB     400     120�i����}V����M�.%e�/�3����� ˉO�^�C����(�����'t}�τ�'���8����W��2cG���<?����7�rt��<�zY8�TX�H�2"����<^��02����E՟Q�~�:�Q�W�۩�f��ƨ��y�Yc5�Mo�2�>�]	c+z�w(�d@�3�\ɬtq��K��C)	g� ��s�� �.���ƍ!��{꿺�&p�A���@�I�6O�d|��V�S�U��&&08�l:����FxE����XlxVHYEB     400     130gk���{
$W�L�To>G�.� � ç����p�}N��0�Mu��ä���p����[�P�w���W�B�(�9�����@'�S� ]���J����!M���<\.v���,e�5�O�(D��T=�?I�G%j���s�Ϻ�,�-X �p G��v�AF��N2�5�L -J���j�S)̾���j�!�Һ�QJ��y���Р#��(�e~�\���(�01��kT�'��PY��u<�8HN�7n>罂.G�T��ľ2�8�T.��胧�ʍ�6oQ�=!�<}GsfPT���:�XlxVHYEB     400     14025��E!���0�'q9�1�5%\:�PU~9�X�|1�m;~��An�c�<&�	�쐷|l>�d��14{WO�ݒ����iy$��LxKn#P�����#o�����xw�����޶D��`�x�t(����jg��!o3�`�_37g	9��G��&s
&~9�N̊)�E�5�h�,�ƹN)LHڊU��~g�}mG(��Êꊴ����C�}�3~�Vq��∗�i���uJN
Y����!T��ч崹E�7�1c$���=�}�~7&�0�t�[G��f|h��C����yU���f)Ҏ�6i_�[xK��j���ʹXlxVHYEB     400     160���=.~�U��:�=��N^2��h�ؠ�S[�iB^����q!��}ĲON�3g0��p���~�{�<�}g(L�3$����2��N�{�)G�>=��%\����w#�\��'$�y��$�O�.u��zU.�W<3Wȱ���n�o?{��HRL�JgetbB�bȮ��"oY��4��+P\WHZH'�Mن����9���2�Vg�M�a����ϛ��k�$��E�$�1���I*�n��U�&�u�PMS� 2��q�p�����ٌ<`�\�P���bX� �+�(����wd.q`��x��i�����ꡭ沾S�˷��~0O�I0�P2qd�u���M�OƁh���*XlxVHYEB     400      e0���)�0��Q��C��A,�=1� �ь=��`!E5�K�����׎�}O`��!S���p8�BH֎�1�#����g�#h�Z=����S�5��W�L�x)l���u�F~ ��ٚ���9�aW�V��Ś͜����7��ĉ{%K&rÛ����\�h7��@�O�0,݂����O�����B�*�J�#���v����vf���4�����-��XlxVHYEB     400     170�R�;h?�w�q<U��_�Ys��=�ܫ�r�@� 2�s7L�� ���o����X�k�#p�ʿoQI�]8��Y��V���5��|&�_=C�xObyv�(@�ISJ�`l�L"��_�aLfrʈ-��q��!4��W!|Bs)�I��y����	PK�u���N�\寴�,��${����I�5!�m�n���)�<Z�&mFmT-�$m���U�&���u�a���gӔ�;==�ϏH�G)�dP󒧆3�������OE[���|�˻01��0�6���ui{�ێ��zi|�f��n����Ώ��1ԧF�h@o�o�����H$'
�����ⴸ�Ə�K�e�ORw�겂&]҃^���XlxVHYEB     400     150-�&�L���1��=;;�]D7�|�\�Pi~$9�����3�/�cB��Mڋr�ՙ����'���-�-����!���t��5�4�<���x�Qr�{�y�kǌl�&��T�$��t���NSV�̏e����ä�I����bZ+o�/6�����K�k
�
����j+��ڏ[�˾m��D�Һ�'�Z�ƵSqz�;8?	[��[c��k`{1�ک-7J���|��~�;��B�[d��#�6s��&�X[,�h'~��4ew-�a�\������	OP\TM�v1�<�F�"[��è'�-�NXe����5�К�3�9�룄Q���IXlxVHYEB     400     130T�`򛽟�ߊL��+�0}������~�t>W��	n̚7��pگ���Xf����0�b'����ٳ�I��Vsg����%byFQ�*g�HA�#��0�E��W ��r�Xv��
�:�a��E��hb���=�Y�4��9�&���a � ����C�,���C�w6Z��n,@�+���E����ی�Q��w�f�ߘ_�|T���ı·�K?0~����PQ���Yr%t]��V f94/���[H��}�Q�<�8��<�
�V���\��5b̴~��t�e֬�^l��
��:,���xXlxVHYEB     400     130L�m�m��n�A��y�@��Kܡ���;��Mo��n��&#��(7��DxƱ=Q�����Gv-N�I�ֲ%r�K�O��+��>�� -�R�;>5�jx(���t�D G��Jf��U/}�uk����Y~I�?k�������3�x��"�ɀ5�~S���4P�/�7ht�_�Lk�So?5=`b���GQ�i�e_*0�VV/3$��f�A�١�|�;��	�.g�\�.�2*��+��jI;��Qg�����!:�#�n����~�/�R�b?��1��2��v�	N'��XlxVHYEB     1b3      e0�mNj%�Gt��EeD��V��ણ�|�n-�Y��>��'�1�v�X�n���o���-��Zp&F%�Ԙ+(<_6-�����V�����Ðt���۸rd$a���U!��D�����LJ����#PAUzo�ID�R�9�!g፪�s"w+��������'8��7�seW7��F�jft�����h�.2����%��yT�)2�#�_�n��$��T��W�����Gݸ