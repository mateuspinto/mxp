`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
tueWitJtUMUtUJRpnWq6Fo8SVrgdhTrEpwJQkONUYv6JVn1ye3BRiFemwGgRVLBv/XDfs2a3xrT8
Xk/YitkP0lZifn7dBjHeGSLVs2cbtGMrBoiQxotemJl6e7fySg1yKWYJAqFWV/a7wW3jRD2DGlnU
XZkLeBL4SslMiI9SOkXjwvEv1mScFV/didCcybYz3iP+7JK5vJC8OdFouL6DskjOoYqTw8jLGv+9
kO4ApisaJh2S+mZI5Kzigj+HjTz94P3q4Xc64vHQ137o/HT+v7dLvszSCSRZt0mXNT09AmIA6Ud2
Dc6RRE2lFfAoCPcIQ6GvItoUj3x/SEPqo9PVSw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="wamxerXIBbfZ0CRMir4924bm7Vtg+jihJ/mWkam/lic="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6512)
`protect data_block
WTabAwo7rHmDWAszcPjjCSuq9C0erV9U9RSsP6vz8PV7m5kE55JoVEMSQPGuOOTMcomvM/31RsMm
rbox6P2aSd1PY1zX7jnngxROpqLp1hM6EslyDlEhGJcXgpVrkiJZ6cFtuGtVDD5GEXXSvs2Cq5wn
NuRBh8uxzTkHoNmtrekmwZpdKsEpKyI+4JXQrFoiRtDecEZcONRamzt1s4kIxkIRQoUffXOdGo6h
BriVx/voX8UpwDua44tBg84tTxlqEzoHCLIByZWWkoAuwSePzPKR5jpWG+dzpSAGfNe2cGk0zAgO
6FE3Z5GtcDUjwUrNm0iQD8lSGYMr/c/RrcuKxJzToHg+6tfnSYDJ9jfzxHjj35mCNys8ktNL+liZ
F5jr775GlUhlatmiHMIiueHFs33Az84hu4nIqMd3+vA6HZH8/NN/Kkk6/H+uOhkhka+QA8TzQ0Ix
4B750oVgtEecuaPYXtxK9rBgrk8oYprewScGUATHFM6NH/nbAOkG70rG+mYIeraD5Z91uiEUVqRl
6UAG9R5VtqHHS2DUnor+yhVit6+EHYXose5gIK50xhKEJP5FtJYNtMq52truivax7McdEntNxPmO
3CqEGEE9eLlFBfMUgvqmfGPvQflT5cw5VdqsCfckaUcIaWZwMi0fB0YkLEyIu2jKw35h1wi7MtEi
NWDaHTvR5O2j6QEqQJfl4g6fx/qSZI8gWXGHCJWMa1Za2ZwEV73x3Tx98JEBxIw3EWOjpDnzzYkO
ebKOlwoOqvD3CD82J0XW2DowB7WaMFYTRtQVVEZ58vBIJ04sVXkVlIYYrmpn62xcMzRqKbtHDqaL
KDxMnV0NXXpnLDiRrccFIsSGtTTCDFzkemo1XEzhRcOPxzHVGt6rgZ1b7r1wrWwQAcP7GnfYPL0o
TbtlWYIB18kkEAyiZ4mv0SueIV+p5MH96D5gAjlOC1cjhkTq7LNG8GkvLiI+Jr2V46qrplwe294K
LMMlinF4EiAgmzgE50xZI09Hw3Zl4YKt2BDLcBmcyaedwlHq5eLSqOjo1l33yok/wUixFZH8vJws
9/0buJy3Lo4iJ1v7fUK5uCrASLTdLZUr7n7kXuygWevNdhMLIwJJIbcQmuIgqx+ZDmak68DrV0hc
dqmyImkn+yrFfLpOQA4/QF1i2gEWqwkwSuKJV5cihVmB0GM7nFpTMhc/8N5RrhJf8sL4aSI0oLN5
UFIbOSrodxQgxgkD/z8g5NODB5qYrrskDjd94LNGqlWmLHzPP+19J0glHnE0qjbZdK179csKRZjp
cqc4dd+k1Hlcz/TMccMOUGBJibLHIOJPG6zuDIfqWhhA7OC2hKXgmkvtKEFw5G7xYfBu+5J3c6qE
Iq0IIROxkmjD0HM7a3eVrmw27T6XndWbwulqcl+a9SvDu2qLdEIvSwQMp3VDsdOznUykemTDBTk8
b/bWNN3Z7g8U/91Kv3PScc40ytwkAKtFFzdW7Dh0QCbsIS9MxlX35ew5wVVjTJ/FbZctCJOncnAR
WGuLMtR9pzl/k59CPIhSv/Wq04z5WREAYZZv3kwveIPOkSmZHWfmjQGlqrer72FLAmM9z22lLnnp
76IFQ9JwSKcvgjT0+s+rdMiAJjf9JJe91cHfW07fqwyV9vbNP3mFCqC0v8mJA0jnY/AVzHowhLyx
eVESqzd/5VMIxa0Sr3x8y1MfgGFRyNG7NwsEpZzyXCGC0xjO/6gUwAeVSuBBumZcO2IzciaeT7fD
Cfj20wJH41oFMZgEKrbSqurTXf+PB/5FaMFtG/IeQGfSlFTdziELv3sghECEZz3y7L7g3uTwC4Rt
mDqNjhgcZjt2/aB+GqlpwFq507q1/Noggl6myNRCdx24S9DrlYDduGpraScIF0B9V6DCwyIu2hOG
xbfn2bggU5nmmJq53zhTT8nXhXPJt15RLqtiApjfjiTlrmd5vfN+OOSNRLcBaQC17sGNvJ55Jksw
SPZLORZLdPaAXDNhm2szR+NHw2qoDj1Hvlj6adi34nPCS4bXif+vz6mZxe5MUV+zIhpgXKXoHLu3
KBVQViIIU+UezHEJW90DwxQTa8pdgeDHT1gxXRLCxZd6jyBd8hNy7yuEnuyXSVRqOBVVoVVYu3p6
Yn2JiDs/p+5qLyE6ZdADncDew9leXethYa58HeVfrgX+pHoUzRM616gx1KDnxe+xHih+credE+GM
VXQGPALxmNrFhnmcxF8EEcQYOevm33Dlw4yF9lFWukxq0BERKuaF0yZOyjjWGPqDibecEAJLFUzN
AU+nnyrk/XPs0RInF3fdCQ2ej9tqa95j3lSa7hVhqKs3ImCG6pftlvHsLIP92K0UIFSshA0AMIYD
c6SE6HgejZzbB7tS25bMlgYXdedDszMdyOhc7wH4G3fPE0nKcVb8wajfXDrgZ6XxCr0St0WbKzj3
9SbKpSxYyYHsFgOeuhkLp468cob4vfq6EoDfloEMMSZhkT4I1Ij5mGcDmmyU7W1daedr1lWOkyHJ
sSocR8IL1iupT/teElQMos3hVm6jmbilurWV1ninq7Wxme4DK6qw8cID1vk0w6Bd4pDaJL1OArnv
E67Y9rZePwV4Jqx+XVVMoG7hERwDpkrAte+DxvYN+ioMkdH6PVUhVq78DvpmHbxypK0BruVRNQ+h
vSB0K0POQW5E+fzTOIuMmGCFR8Hif3qcXOIZGrir8+8WKcw2lL0S+7uEwVOr0VWRQRG5IUH1fv7N
ueZU5UdF2qDUglICQFbtFw1DPm0t+eSMRHvzyvnySTchQpp3N4f0ItGIcBAnmiu6KFObDg7KSxIg
CwjgXxQX7PSNy0fRrEZEuGrth9AyDmAsbklCKfDrJ8wo4PHHC+ungnBTEzESNjIUC1+WBWdbYBVu
chK0RT7OyTQVOPrvoLA4XUO1YXEGSiCcYYEN7AgxcbKeDvsghCLbilVa0GOc8z/Jxj6yylovNiRY
M5kkj7s6YemSgjaDAa4vpLvcIr/JpbBYumvzkuibKOEFjUEtiMCaizf8Rczt4aS21PbRoNyqc3Ey
I64oE4FrfUTTEXGkB/4JNt4TcPJ+8NFV9L4FXIf72DSVi8lXNYkJYYUoJu+B/XOghKOLbQ3fv843
hkPtVKX8eXNX9dQ36NbUXulPJKw7Um6ICT/K69FxgCuWyqHfRTDAPXMgi3RycIwcawANdFBMDQlK
Z+A+wQboK81VvNyw4X7owI/G/ez0VM8ar/OXZCBe98hPvys9ZNOT1y/ezIy4MG50s/RfKT/LYJdi
QRP8XeZ0bLjn/24+QSHQGjN+ByhcmfSpMHRAc8nsSSkgQ3Pu+3F814QlTWwwzcPgl/39cX7oQT2l
lkns22Mm4UhEi1CCZEJUkPTpmp86hp/xc1GkF38+v87KVYrpUocpuW3cNL5GhSN4eTMXFIDyr1PB
Ti2DfcTyRZ6ffg+yH1HUiefXvuCtPnz9sgTtUriMEF3/dniGCoXQDX4ksJFbkdh5ngWXO7+DqVRm
NOyGdgb0BbxPWysGcwoddZ4hxITH5Q4qtMcuiaRRlUpwb2T+0kZ7wqyz06V4mAgQ2zS+z9CZStBt
sh+vImLgRIIYxLS9NgJ1wTjOuiuDLfZE+B0qI9XlvmDp3Ql24yyu8KGtbI+ADXFHiYMdUN2uHAmI
E8Zjf7jfwppTWFNE01wFQi4y2so2W1vtzxybhEVz5wsNlrv9bVkfcRlEPVbYaNRooUEeM3fMw/2h
pJhBouD3a5lvAWZotbLiGneuz67lkaG42wm3N0z3jl9fkYbc5uEi+pcu9JURXClpwd/9KvIH4Stp
LRk6DT34Ku0JySTrVTF+jsusZeo4XgrWN103GvNIDI05qfs1K8/lwwq7Qr5r5Xcz31UoaC1tdh/1
2smvvWQq+g1H/HdG3fVqwZBjTG4bwBR2JzyZpFr98IT7jFIzxGFdVPN+i2voEje3NIS/qpkVW29D
OBFTvz3hpF/Hh4VSrxDrO93TNKeTP29rGdZ5pfxcUGPe23x5qIXj1axmLxK4vBmJ1gnsXNjCdUuE
lcydFeTHv5a4zER5N2AKygInpghhKTfYzzC0kBmilDA6bc5ZDzVZ9p/3xbswVl6/cSnsiMS7RUAA
Ool8rXLLbEENyvTdlP1Qj3PbDzdoLEy1oAFLY3bXtOH4jE4ePnnf5uyUysVEzbbmBAdlIlXnSs67
BakSSY2yCYChbAK1c80gHD7h1dNILdVAQmfGpbWuS3XBIfSCyrrDjkULzKjvausnZZLbGcgL7p63
KpOKZXMoJMB5krkGIP4BXEtfLVPSBcBno8zWoWq6QR0HNaYHwZLIHIrCCwslCELl/qdRB6CiKS52
H5jFuFLdFObnOQBQfHN1Hk2dNmb1ASwwjFo8MvAEbvdY5CidwTt9395VRgojvyqK7I4pLrZ/7VIi
2A0v3TzO1uopLfN1tmj9k0W4VzBbNs0EYepwr5Oy0S8pcKfONNgWYMqfevIh27PkQxtAivVPL+K2
5QYCXoD9dQ5ZVC4frWiNgJpzhFM8VzdPIDCMZkURmJEBV4D6VD+uhrw2fGvEgNCnZ/s/ONN6P3p2
ppPcQ7HWqXnlaJO6uGS100835xYwilEZrpl9hb+iygwXfe/vhhJLAKl1fOPO1KwJW61hgFz3JHB8
V+ETESBGMCCMBm2b1koQfbTxssT5a9gm2ZqUlsoUjkitvojqYUb8Ku/U9XDHoRp1M4l0TXR+K9w6
tvteAsfsbTjsK72Zy4bmeioDENWpP5FgAj8WRWE9KZsXsSOqO/P8QhwPogOsHJjOTnuX+xDOcpKA
WpJwnwTNV6p5886Pao2X14gzLfzfEaUBrgf9efl09CZxDz4INwXiam5mVfyKWHebjjU4jOaxqWa8
H9sz6mvB4RmMqZ/HxEeP9tFjd5Nl3UE7E4r4OqSB5MkSRfR9gqtJW0eOuR1s3nGYUd+qNx360wBJ
rg62VSfNo4BJJyqJpwGJp/Jlayi/3vh2y9tkekBt3mQ7+p/dZxhem67Z7cuQbg6d49JVD5+DPTWJ
c1pNVE+y1EjXhmkM9+cBxKzN46uvRwTeH34CWZTlHLgPatpTpLj7ZqIzxBbB2Fo19hBElTBRqRgX
JdLsxlictKJNnAwWTwrH/kxGhvqhkW1CV74dWYGF2x0CA+IsAfzJfTWcfWa0Th51mWA+thMGw5k5
F2diHpfNtHb4PwtKIkvvDP+piMaC4pqLFi/leoEaJEanlg2TjJFBmQX1a/GUdfi04ASirL2pitjK
iB/RNp78OqLhG/sS/9WWfWVCnUt2YudXHE1rWopVpQlWegXDC4cNYWwAYvWCpdO8wXAc2iLCunAa
RHkeBq1avYjHImmf7in4mIQOs0589no3jqmI7F/rzKT9evw35YOpCY/RGBCqC0PiBnSVH7ivzx57
yiPLbEdGqp5FKa2OiaRqzSeowHcMcDWkLhYDjXyhFOZADeHLbQ+JRQDkXF0c2KBvNxjbe2oEYDOY
L1xxFT6rNDEbdIMVstzRjA1tyCJQgmc1ytvsQ6ZyVMDEhImTTucuymn+5BIt9OALEoMaVQq8cMaH
oPceIBlfCk2fG5Xaa6hdoZLoy9SolDBjUIdJW2l6Xyb2vl2ckP8tqm85PO2tDULcUZUASYqf3dgK
Z08iIKxm6bomhviCdrGJa1mH1t7oX5J9mkjvLC3PRdaoHfpjEemIH03hZexeJtOIoMUOZMnu2+ZI
/dVsHYY/CFrbsKYhEG0XcJojuvESWI3qMV1rV4cef8YqjsK8ELYV+vxYEMFr4Vl7+kSqCVM7jam/
/krUxHo68Ok7T9YeEpIIzXfstxnyWvMXs4H7xucQ5rqg6SGbf0aMdAts9+aGEzq1vI4Dun6IQ91L
BSDU4cYR6USDhWKrbrPinmC3nbKRhpZNI5gYph+U3Q/stDGnzjh7Kg7AS5xlHQWkZl+ahJ3fH377
fpLVSxfBl0hzxbR1xAjWb4FDqxegyte34UWuc4V0TF+nNyeiTSGs+KH6HQhcfrlpLjXOPmXI6z3n
MWxoTFoaFpsPr7r+NMvOroVNPRqsMRIw7LFUV7JQce1pyGv2zYUdNUFrGK42DEJJpMnD6bvm1RwA
TFuwuo1x4EfZCDa8CWfwfGH7zshgQkg0S8DFPrD84xRgG6K0QPYAE/nCXQAQMYsa/Hw7zxD7cA9O
7SXNfpWjBAJxjRYHdlpUHN+eyMjwRYx5OEPFU4ul3uta+V0IkKj2mTONlMAyq2TYH2zwXr3OX/U1
8KX6PgUd3V/k+u/2KE6v73aZLnkSPauWHUQbCoZfFo7tsi23W4mbRk6HNWO1rx7KwlP3EHdAjj4s
he6JVKexss1hZBBtSNeyzRoQTydrFHWb/bIy/r6tlZIldbnCi9OYu9Uhbe2IBlFDSOjJbY8dwm/2
9S2zgu7FSn/9J0pBQx4iR5TiKV3YeTORkNUetCne9n/h5JkXa3Bpse+rLsQTPFv2fuU0hL2AThWz
YFNVLlmVkLrkl9idqQtMcDn+G7wptgammMLzMrbQ1Q6NnWAFpUTzEhIzOaRuGqJP2Zusu3fjEDox
m/6RSgFrMavSStPquhfWW7kWPlxm8SuUNGOxqcD2sALqUvhOzlQ7MbuToXCNTgOpNcXH8RcI+qIP
tNc05EjIs/8ST3WdOZ4tj+0TBLXBXYB++66YA+my63ehIlwRxYBszyZ7BmfUwN7OnyEgvswNTHDq
XtWwK+lvKBJzYdPGWaF7kxcI1OFt6/prdCAfuokW2G7ttxHUmWzecMb0i+A+7lePkqHWMkwaOGp1
IqCejP/YRfQTzd89jBtomplwMF8PApJhkLrCXMHyFP8ScHUSNsqfBLDAXU3lI1EXD/bsyOFI/D50
f8LbLLVanXRFtO4q5Wl5homwn9vHgyGxASRWEeIEE2VAlOkUgTZmZJSmrr9vl5aKEeGBHFxqxxrq
FLn7NS5uo80TRm69dsjXPrnmGb1vCXmqm2TFfR2D7GYTjUFJ11+tmHcYHyVTzulVXmIdEdnbJcSU
TzDO/HNSg+as0iSuWCL/68ljmNdLpxkeZO9J7kgU4LhQRVPaJmPLQt6bNf+FTv83QABA7t3bv7Zt
x6bGKe9geEU6Hvw8WSis1vyNHT2v3OckaqP6c3og1EazNtcV6jI+ewCKdGQtT46QaJHWWS9MZDbS
wRF99G2XjTTqyyK7VPEP6Yl3hewEwAAjgOXot75l9sZ/BJ3es+PmHrG1rjp70lnrqR1lJVnnQ4zz
Ks13MTfsFA8emOpuQ6nZ1mhb9Raaga8l6XeDqlGGfTBCc0E1/QVuW0ZsCZd+7Dt4JRmiZj11OvlS
Ud7/VTRoDegcXzV+VUFsMb8QXVqLbizjPdtwU9e7E9svLm9P08yQjDNOPBvUNRZXSx6NmZoIvikN
qiLwSaXCmXU0lvdXWFFD2g5SDD5vkHPRdoZtbv4AhhgMVevkvnYsmCHBBorIr6lT3XVyJxvgj25H
PzFdGpAh25B2xJc5o25J2nBrHxBiXvwE1Yx8mjtVm8wkaKbfJJ4erV8enGsBTaYbOVidK3mESPOm
OnxwH15BjykKoaEYsYVjHznZPQxRQQbKpP9O2gzbr8O9nfIHi/QzV6x41lJ8mrqoqV5qMYsruyf2
lf/Pnu8cJYvX5hEaP95/KY1Bw6zDfCBsAiWIvkBd2n2YNXPZc4bWylsdvQYXbj8kSGXUzAP/lRd3
k9qUkf/JqMW9WGtN02Z53Povr0myQhtgrEms9g1MGGHDWHFZsv2Ulzx1UAOOSEePhbuMqhZy26gT
fwtQi9AnPgaEJxEhyddlN1lUvitfYDnWc4veofLOLRitBc2EQOBRYryHPilECOa64JVIO3ZWaSa0
grofPAvp+1zK4KjbbCWT8J2bHS7IbFvBCt9Ge54m22kRNx8USQGLjvAmpG3tVyWM+ZmqDpNU5CKB
TJbx2darICSOVL2OkVRN299SSZjukZh3KsWKiZR9YKU7U0B/toqdOoeueDntH9nLN7JMZ5cpb0Qf
MV7rwj7Z0KoWW9Ea+S1fliuIVj4Gr5Fc85k+pND6UTO6USx20IIPuIdcYt0QbtMnhgYK/4fpZUO7
t9KdmK3P8o7usDHnogN0C2WSK7uHIriAx5rYq/7Bvn/JktEyGdwht63hLMTnbwI7q1vnvnXTaEyR
P3HyxnZCkXJn02f6NJ0xbuB+M5eRKHwFohjso3KaaIT1qbyWAQx5O9eaY0ZE/HmK2NAQpegGGLT/
SMTZIwONb43K1LuDroSyIwKcmt5rzz5jb4F4nqqaXdX/cyGWGFsSh2G+NVLT4MrbSCJelMdzuwT0
fLCL3khh6Wu1RHQNUc2XME14eaM/xUXtJYXtrvyGNRaYFhJAzLXtrErnMIXbc0USJK1AKzTk8vqY
qTqckbl91TEwvoT+ZVzYPJfrDXxsijpp4SE7s7SF/0JV4y3bw8Ex/CtZwHFaHHUfkbUm69WGKpxA
3xRl/yivMUe0Or0rAbcwHlsToAmSGGcIyAD5tI2UOhG0+y4VeZmLSAj5c+mZ0XMlwkl3tjb1ainS
t0ACf2uG5tzRqm8on4Cnx5Etw4c4sYpP69QQS6B6ofKdVBe721IdwXUk98nhAFhXg9R5M7Sh/rhg
PhFqq8fxAE1qOMNAhwlj3P7ZDCVZdlqdHAyzi+dKGFIlZy3K4mz6EQIVOkMN6MOJoGawhI0CZgyP
aPhIVdO/LY6txj+/cc8=
`protect end_protected
