XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��jpB�.��T�?� ��Fj?&�QPdu�[�(�M6����#�#*�i�:z�E�͛+ڊ¯o��F�G~�Y��id��z�����91H��x���IW�0�-����N�@:&b����a��I*A�j-��&7s��� �h�Bf���Uy����-����Re��u��"��XG��B����T,m.�9�m�u�TP��CF@W�К)xt6cU2�\|8����ך��&g��hލe�����$��h�sɴ��s��FJ-��|2� Z���h�F>�*�i���͇�1�o�����D��.�p���c�[UB��,Ho�3�p���M�����!Y���D�N��9�Þ*�6�8�M��S[j�^�_��5^)��{��_�ޑ��,Tćq�7'֘�Q'ʛ���m�v3YE���c��p����i"����'�����0 ��Oа��(�0���A޲�d5��#�[\5[��X��SxCz�XU݉�=CkO	��`�Ox�#����*��l�\hd|��Ґ|��]أ$]s~*:D�H���;�JƊ���G����^1h-%���Y�.M�7!E^��ft5�ǉ�А}��yp��=��w�Ja
�+��mC:������c��Bŝ='8XiP�,q���	�	.����L�,��K�c�f��N�`}Y8��7�ݐ/�������0�E�7<��2_�M#�Ʈ����s�L�$W+�Y~���+�43���6���U*M|G,f�+��ff�V�x�ns��������kXlxVHYEB     400     1e0Tt�ez6�m��8�=n+����C��88��I�S2I�~c�L�Qޢ0s�2���%�����W^S�j\7]����X�V���E�{g> z����f3b+𯸉k���������q�۵(1�h�ct���R7�&<�
9��0����&�N���za(� r�#� ���X��T�N�����b�>�W#�	o
��G�1�X�f͸�e�c�*��g٥{��Եw�
�l7/z\r�F�C��TTD�Ѿ?�&z��r�[''��V�R}T�;V/�mo�^����CIX��EHƷ���x�%�����0�Ln0����:f���\dĠ���1��������^}�~��Ml�	%#�"�O�2�=Jp��|z�'&!՝�t�_4��'h��K�qt��Ѻ����ˬ�f�M��mi�GcI������pL��f#�Yȩ��tCiI�	��ԓRH詄]�ĩ�t+3�u�XlxVHYEB     400     160#��qU�0�:�hN-�Qo�őZ^�#��cKUqXb�˸h~3�dE%茑��T@O��U��;`�JuT��ҽ�'�Wb�i>�d���#�e�L����p�S	�Cг�~��K�80���r78$T�E�����"�q@�oE���#1#�����w��n�|-��~�W̕�CVO^��H�޾��,�;�v�+U/zh�o���v��V������3Dh��!�`Ċ%�Q�`����;9[�W2{���΀���=Y-A4�u�	y�3��^@P�~�M:��?�'BE��ϋ	��c��ý����c��Ak����`?&v�w(��!�D���7���hN���<M���nSXlxVHYEB      50      50���5�sn�o
�s �VjJ�g�u�b�1�A�ި01GD�3i�� �#ҏoz����Z�v���ws���"m�^�"���