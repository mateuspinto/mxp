`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
c33kqhSXknbEza21bFEiTtZ7/lVhjlEjdr3MbWKfo8AUiA9vgev3a4ybIsXFFu9zmW1ZnXtqxv2V
yF9MMDyt4SG9Sb0FGxoNCWmYLyPHmSZJ22B+QA6+dyaqogDQ///ZhIWgC57HO92P0i5JFHm+3Uww
ukRlKOiqwvDd1QMi1p0inEt00pkwzHL92+VRJqpbKHReaee2yrorm9qBBoet0X5LdlwlOf+MbpSk
uG/iLBvyGFFW+KlhDYc8gWrToq8L8DqRHOzKRz//aYnJG9R4FEVzP0F27YpHMiRZz4g3aSJ6WVwL
uEWLPmtK0XzVu9mVNzcj2jhhwjcykKexvn9QhA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="oXdk8zpPfvjcpiMHWZ4Wdr/zbhR2zPL/r1Fv99ArOvI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2800)
`protect data_block
E+xW8EGx/IUCD1/syfU9jYFevuLAz/6MU4ovlRpSxefvAkz3A+41XSTHBsyj7xcVnx/TK2PLvYSB
eYkNpR8FKhvjM+LFn8oToMOhNXcoMzRfsqA1An0kx3tvLqFYyqXQKL5nRt2SEAgvZlhdnOEion2W
PMl+uO1g8v8bNNkz01cbnKQwcidYoCoDrJd0yQDhww/y4C7gN5Ts6dukfxnqZaO/PBkrIkPRJ+Rp
n3heN6/xfLQ/0/19laU3+XQbWtTYF03y3KL7Fhty4Jb9gQx4beVUCyjxxxBp0GsaFLruFjy+OZS+
7lR7E1SRd14j1PefG936opfzKXMox48mJXLybhAd7qCTFMyyO+cFWrCRnEJpx4deaBoiSMgBlvr+
J3uMOT8sOvIqMOvdAnE8+RzD9yYavvZcaz029MOAQwtQkW6Y9+2orI7vIFJD6NKzVA1aYAFavBL0
n7599U9OjIdO2dbKI0+oosvp2uU69kGcfRWULWEJB0lNeslPjESgYc5Ods+AzJe5kbbu4LdqqDf8
+nOcfzUROW5EYN9SKNZ42ajNMyUsElaBStsuUBTmHoiGE0UCxdDWou032QMUvZ7Zr1QsHchpfFuH
Y7dfQPmddh80ImDwFl5Xys+FvrdHqAQxsJnR7ZGgANovdiZ7Eww5hfzMCUu7bZ+2hbdwkfbaCgl0
XbZyYPiq/mTZHU5YTiMtK1gTaZVVpVOAmMl5ly89uwIMjmekC7+Ojn5hVg2xFVEQ5J2Rhrm5nq0B
2rirUz+OI5u0WlxgMLFRoq3TAa5YMKg38Y6/xD7iclTPNDI1HCY5s/NXZmYuyh/14J+ysWzrB/LC
K5pSeQ4fYVgRYUAfbGST6xWESJgOG8wsDidmSqmCeZgGR+KxB/er6SQMiGK0GbzHtcxrZup1etAi
KrZqSsnh1dksFddgIvQ7SrSRmxiax5DQYOV2YGFrMu3191Bh+GcuEiuOJLFmVMchUMYQ1n+KWcZX
bPpPJSOa+i/KZJPdWGRN2Bo+kcrNNRR4yoC0N+p7bNY1BkiFUUXClqt+ojTOeo3JHXGtldRxksoQ
RT4UHTpDAz88QAl907mSbv96QhfxVw8iWdxd2ohyjMYKPaRF6hGgxx/cgvJy2nhD44+qVvTA/UY9
Rh6WQFcFjC9HPs323ikifqje7GTnPtAwcvBslepVom2MyEWDYeLijYhOjbZJVzPgCiuh1FvyAfxO
wQc5uDb+ATGFVwgYqtdM39W/lOSSnxyKATQgDxzNfEO4gSFkljsVp63L6A2YmeJVQnM2Hm2D7u48
v3rzw3SgPH/8wg5oGgnGj9qpuepg2zizsyHzLrpq3ezBK/XGRFyHdEF7jnpZj+cldH33J5bb6fhs
ZEdXIaYhbvLYfFn9PJLWsKSxcc8LJYkhtArCiLvyh3/XE9xdZfTWflcfpnfQ1bd6zAVb8j3w8HwF
uOnOip9IXnSkhbmbxswHIruXm9ma1LFZP8j45yAoAPUjLDq2bIsYZLvcdXbSg+6LvjziaGGQSk2L
7wuqI9U7H0V2oiphoe+I2rgxr3PalIVLrz0OPk+AGkd2C8djuroiHWzLtA9JPJT+5OJNTtAvoMCQ
/4T3EF5B7lKWZuGlUA88eit5276BryUynYdhqef77hZJ/ZQK17B9Up6r7iMoszXlE+oFZL16NBfQ
SyKDNu7TLzkk53/K4M/fm51tY4N0ujVKqQWesVa+Ef6YU+/zqfBYgpzGAfBCaSzmddVlMIoSM2an
eyiSwuxN5K2CtyQ0btmWQWCTa/Ba5PQtvxDCEgstFk6FcfUZZM3HA53jT0kuTU7qoGNx98+4mAHY
tB+cPZ/Yej1/hm5lpHiSBJeJq9cvNkFXEFrDt0MrdY47r/zpxlAkNNHJqREh/wr1C4U3+fO3GQG+
Z82etU75AwhMjpla8VnnOiGAJSySrznjz6YaEoQQtHsdXTQLNBfJM9gl5RREPh74rfUTzea+fsnI
DAzVZ2OI7jnm8X6MZZkKGim2zbKaptXBrPIxs97qwPS4FWmn1Z+ECJtA2pNxnJrHjxsHcTEtIvk2
eu8FQdrBIA579zLMOimTWc9ID0H93bcR1bOqvjn+TFAYaiHDY76shXxPAN4AAHz7wWJfHPjTM8yG
1TyfnQ6h6MBjySD4AjU2an7IVRoEOZVvjmYRPDrHR24VnFBjdgRSKjDqYJVFBgGYsLP6aalSypKU
3V+Yd1kDWAjoNcjNDr5KQzyHdTvX6+cQH1udJDMOpV6wTbjPTxOAivVmtyy5yF/xvSmCHnbuTcHe
wt0Y50yjB99dlQ/f2emKZgWhtmQgiKgMctBPHB+vSqtxUJ6W5SKg8fX6To5i3Hwmyd1I/rQNMG/G
3jOwHoO9oA0zaRJOixQSffci6S7QwXwqLkAtBQq8M4ZamHzpxGTsEn5or02tXpayY/QmmMWH7xUg
ub4pmoD1Qqhicuhig7+qrzkxvLp4NcTKRAE7p0oUSl7/p/yzR/MXLpieHv3s33kRHoQDrDzfZJoL
VLopPPXDCoVa4bVFTxRj5m0UVK73As9XdSaddfFIjxMlNYx+bzMMqa6Lx2nUQ9UnBjzFzkF4ZPwL
/3H24qWjQl4X8uLg90AvTwL93s7PGgOs48AdfDlnjWFiouEONbbKI1tS/A6slK0odP+zX5npnwzT
JHQBDre0s7BiwQRHKT7YeUa1+La7BpV+u5CwBWVkpTpTZGcO26hNlHFIRTVZtAP4dL6zuppXJeB6
yUn/B0m78whwAFGipFmrXv+UzKruo4AbcOb6T0PJkyCTC23aG736NlrpeaTiSxfDhZT2q+Z0n93D
mI/VhxS8JLDXcND6nWjxnuWA1z4Rl3dX+XyyZXhVi+NcKLiaCj/r6SuSYxXNnDXeIHPcQQX0HlGa
Wq+6ut8xoB52DAzslPLhw3H8QfM50any6s3htX0099FTO0Tt+GjmFT1TlmCv0P4bF05svo57TG+7
+RNkJd0yYU1JuWn2sIRI3cTWfH1QWfCz/Rt0unosyOBaqTxmyzFqwh0h1b31tgl/w3BtyZaACqG5
rdGz+DUKlDSIZee8DKHHDg1T95sCBoam0TWNnIPHFyZ54eTpBpe+vAjnB10ygo0SFsvnCiXtrytz
NUvAMjoHcupain9b7XqN9G+Mu663Foaxw2WjZLffYJdD2EIr/54VM4wal8lxSeQiqcHsr3j/9d5A
HUhAzprohu/nBtaSI36sonY7vOC7SZ0RbwdvF/UlhsfS1m9Oy+mXSTuNWG7t8n7YSk9wNjK4Jw7A
ijQxHLCCJXqUaXxPIIQODtwXxiu8nvaOubWBr4QTMMes1o+/CNg3zFLNz42wx7kJRVh04oe2DnWZ
7bBPBFXsknnqYCnFHglIVcJ6Siavb/JUpBcAp+/TeV4w/ExPP7+UtCRHyhUaXuGLkzv3sihlLrTD
DQQDzVaEWs2XqZboQNX88E8PRaPydrd9fEsfGBVi70qJBppgR960gQO2wq23y8n7r5XBhYyAhTOK
aEXJrc3r5STXzQfeK/jQYQJkwJmiRcqGBndutPMs0mGavLtgCfZL3x3M0aI7x6AMprrGOeT9+5Su
sMqWoAjrjVmDgTaM4XAM6wKvMAcCqm4H24CqYmpKLM1OR/gYj8qrrAmSuxfWgg7F+A2izt2RwBGu
eGYxtleGCKBX5nQmiZEZ6SYHgAU25tpA7XCVohXR1kBsPva6DLC0WGCkYLiVbgvJw5oQV4pWY7Gd
LR+IewGzvA==
`protect end_protected
