`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7472)
`protect data_block
esMTwiSnnLprfNVzqBwyIG+RHeWRt/YpKchj9LbsTzseNZNat4lDBUxsFq9DlId054pxnUYZC3+j
bJ9XoC5z6qrYZ3gRsKpRYVmavhQrkoAiMTRDbex6d/v4SZeY53SFfYsjUNuNMgLQQPQXgTKFVpV8
06m5nXbM2id9M76mc1BXD7yFwere6AmNpobqJh4sUQSgOhwmy5YJVZ3W0yPnRuWWjklSoJHBZ6i/
1WK5qN/RnGCA3qRYTR8zTX5OwPVwlPB1RD+qfxVSm2Bm18F6YdymXGlP0NDI5VUvArmAs3GSFp4h
/jRn6+rW9aD+sVvuS250FZv2v+G5Rqe3aNmtFINJDIpYj8q7VwSeoDaDmBVvMgjuw3RhrfJxtAiZ
/zbSqKkzXt14Kk78msb6FoWe50Cdy3u437/DWWUwB25E4gmk9pcOHS1EdFfsYxwyH4guNC4uecxl
m4u/IA+oaZaKFl3Dxb2TV4/SE1/0P9AFCbRWRi0PG2ess0GGTCTXs6tlUnFNEBYwanDXcHIWfdHG
PC1CyRrbIuEQZHn4iHnDijlR3YsRU88xJNyiXbqm/SgA7enBJxNmhqVgXiXGC4ksTvGfUwPH6Mp+
pmlWWqPGm28dIBXsmGD4DhBPoamPiXgWSWYa6yTp6uE0adsPqFMcDU5bhi2OFtiWUukyWzdOHg8p
smmyqTIGkUm9vZiTR11G0LqGiz9hrs+dDe69cXjEDiYrwo5Mc1Hs1If5tFiZpc/GAgQohIcgIRVx
j253wUcDtnV7Ua7JtxVu542YzXrEn2KMJlaBidtIc/wixCY/lQn0Hfnmgw88kAHcixG448+gV7S3
jNb5yDexSF0WbZNr7AphG+b9OLBanrl0JDO73RxRLpgrLAY6U8NMiDDTg/49aRNLs+PYI1geF85c
9pzeDTw5ZiZGPmDGmEqk5ak+g/V0Jjm0P2S8xtYOgGi0buY6t6Uh5ha+kAWEpY9f2t4jTzFC+Q3y
gjoh7Ew1dfE6jptJwd/fcpfbvu12E5a0TVyyhFfdkhRTigI3CMSWPuweaFeVZYbgllmffWvyQlTm
kTs6K+/4llOoz3pGn7zXEA4yK6FEkwZrNg9VCvmf9Llvp4b1PUX3oX4B8Yl+4ppla9zKwW2euM34
gGyixk9H0Ky/vwDUBuiU6jPAPPRCLy/2Bms7NcQYTiP6SwBXkemiDm4+hY9ob8dalDedy78nmPBT
I7HP/fURF4f0kclJt1MxQhbVAzML36ghaDqFJAgsHJKUsBxg83FKcrxTLeLBFJ3iuicK/ZCBxGhN
8GEw1nWm8H0inZUnKSEqkko0wYi9noqzOeEmxi/7QAcbd8IrZVAFNxt+9/IyI3hZxXInHRMC3RxE
KS6a0XuNLohlW5TvX/nh+j55Z4YAYZMZqArROVuaVi4F4UKNZjbm6+RS4mvYc5UE875jGRnYFTCL
MDTp4yW1LqHMN3WJvALC3w1t7G16oDHFrhrBxXEbFo2dqDmUj0Q7ezZLQ6nAlppJRjlL4ZctUOzh
7wcd8WycrrVruVe7f4/3qCOJjaKad+tX912Yhzb95BwaGFqN7e/T3ZwP2TScG/FY6SorDLyXwhpO
IaNVIaywTOPW1InrJ5BsU7yJLyFJEF0jyJauQ1pk0LNjCbzzYrklbfxLWta7TuXGn+FCpiXsto+6
2lFKz7ErfeH8yTC6A8X/cS8Zo2SFeXxnPiWjp3bGxhfbILUX4my7rVEdptxb12mqV3kxxPjjxvI9
UdzRohttApKVlf7+wevRtfEMySFpQc0dWeXTkFzlhzYS0HqRAIR4h70QT27YGum7WAIcHXy58KOr
Z5MmK9maESnadTTLShm64Ah2+PrI3dlNKSpVD4DjvZ5EAuVdXn6NuzKZXHDtngm2n9BUbjrHePO7
+X5cVL4XTXi7yI+CqEU5aFFZVL0bLE4VxHPz3/KHCMN89ri8+TxcPODG+z0LXlOje6zCMvAcL0Z5
TZYtvB0IQXcKHn4CftRQ89aDdxBn2NIB5oaOeKclqCbttpL5P1BzRFwjQ1fn6n0Tc82FVoq4V8Tr
sP2YbtHuYS7mIBb3evay+kMMGtP487xGsbZ5tqciXhHDIS8/QLSH0mV5Vr478uCAJq9UefNWpz84
JrsKxYbbxIGadFEmTDZu4fjj4pMEOVwLGp+/+rQty888DuUysV9Ud6f+WAfsfjl4rwlEQvaM60/i
YzIou6BtJ8LFLMh7LIlMw+8vQnZNimEBUEVuvepypyN+LR9L1qa+44sqFAApN/fD7pTLy0+CWxQV
8Btr64RFcAe1E0VsGzwsp729nXMgroXCYd0S9XmUi53sCGXDPUnl4nYq1TNCw0hKLwJYamDsgQGo
OKCqznmnKm2FakjORbadIGl08G7KyGtbZGJXLPYBUS4pnnc9oL+4lAf6XH42xBXWeH6vhYQs7048
o9/H4U/eKQXx6ZtXqY7rqQydyknHTmCJfyPEDkLw/FCwQj15ukE5t8VgvPS/ZMlx9yzOKiIBHyHk
qDIynG/gW2tAd06bkNpuJHWjc1/cNdE4RI8paDonpO55Km0g47uNddrO4esSYoOwzHQef8D6mjwp
oLo1ClMGiioev0FQ7SOZPYpTMMZsIJLSUx4M9lBRXPGhFJnqjtX+muBd7eY4bZblawMahH3sUR6U
PnB4GG10l0Y5Sm386yqSD6J9jB576nyNl+eHZa4ZOvh+PSlTg8x7B4qyCvARwalgjLp/xJbJzhFL
IhSJFRYy9TFnf3s7ToUb1CVN5A8fnpvkEwgrDnjTjlAU3PdZIvEwAx54Kued6xycQvPeWaBOoStw
iQ7r7IAwCJFj+pMcxbKCFP+nzjyXe+e8tdJn/VaKO/pPIsaN/Hb/Zp02C+gO8g2wGkgamwD2Xl2m
S/uQKvqQr/QSTIDeCLTbRH7E1a7Tp++rBy5IzYGfFLD8hjJYfCMsUYEgWEIoeMqTVggdsw7NWBKo
oIww2t3qBifEs++pekaYyULlOlsWDNGw3eLY8taZTWPy53XwNvOypCGF96OF9dQolJyYbp9OmX0f
6Dqzgi1Ob1zkXmrhQBF7GAYPGBxVzAfVSIl6iQb0dqNJKrty73WY7vEPisTArPH4ECJ6hyfKJZ1P
nSvLjd6I7eup2GcznThbq5WvsmBmP5BB9p6ysAOCbf58cvgse7nRi02A1dOCUBgMAJ5jvSrJNsCV
vrt8aicb8HRpm7lHaqHAL0irkTW83CzewrMzT6D9b6MZ9Q1eoBoZ4sf6BDJ/AmS5Pbxm1wfOgfqg
P9pAkEuU4iMKa0Zp+L3yAhXVLcSbGVDUyNz8tk54ZOwyKpqsVeb2ewy9AuQ1rQNfj2ZECRIgREwq
CatCOT7xYUY5m7Iw5XRDDanwxFuGRJHZJy/YxmJV3qjOTa0OVzFQ0+VfL7c10FUIV9f1o8gWeP1B
+z+4wMg0aBZ1VOs5+niH9eX7UIfqym3gZcsUFfbWox51uK/I5pt5A6vsSfGxIb+9wIa/58DktDyD
NYul/8pY2fy3Ai9bclkoQhGy6fT7B6oVOrXCIXbzPPbHodABu15YnH62DTggWdDebTcREcIibOe6
S3i/dswOZXbn1zyQQ+by7iYEmG85kH+IHJHvmw1X3RO8/qQMY1TTA9wFfqB3arGIvJxp195JtxJU
MHWZYcdeg+NsvrpdKpIcXEZxSGLy3R4de+h3roMdSyykPB1TgAXNhcsrjxp2g7NgX7a9tWaRQqs5
BudvjjQcazXap5Dqgj3THAXwaiJ3hpynInu0J4oW2d+DZ4zww2eWxi8uPTg4saKbzMoKalIcFZ17
kcc/rvMcwSSFASEofFM+jrJ89WCOm4jc+GflJEscQFp2EknLi/wTsN7aZipWg+dGd5ltxKCF9UKA
ixZSTQCMalbcdhKEx2VMnV60s5y3LuVO/iSu5sed7NR4Eo6elHMBnTQp6t1E/5l2Wil4zwbY17H4
vzaqVGJDnr3iLjyyOqoabKeYdzUeXcbw/4H9XEmkCVjUP00eDYnv/BJCEW6iLo1QdrO1ikKKPrYy
r4Pi3no3BhjV5fFoZNKSF2OTF93b2+rdMUB1zqVGeNqdVY+PTH3mEU9z3M/AzwenxySkibrY2SKQ
KxQLQ9pLFuxrCwuIv49Mvarqy3zv3w1b5pmxGDC8OZvJFRqZmlKI/giem0PmAzS8OEiT0GjPPCkh
ZbJDqG7VsGN5y5QZiKS4kzjBrmfD2eERjMaD6dunedoGLyK28whU5Z9Z02AIRZBwnnPP62l8X1mc
kZe8iyKhKD3tA6b12hEkAD92fYKAaobWTy/VNPRFfiud8HOCdaZbGrSPbXA3s5LZEt22aP09iko3
QrNKWYV4E9/1OI8J9yUMt17g+ucbsbWSy4lJbagWtiQdYkthJjoUR46Q+0/XmD3BfBdWOW9SBC/j
zqGJUanq7xFjHU8CPSxJkPa6r4FjBUuiXDqMAZ2qRgUqDbcuS5iwaNsbKvMESP3vyolZ4/YjCBSe
4pATgSsuqmvSfnTwzGyfYdP6vw2GAXicFgGUbPng+k/D+B4Mo+XLHoWnJtPZDgqCsMEV2i/tEk3n
fSowABg65gGaS+5zRMxCDILeRMrToiz69XtavZ5ZXlLK6wXaJuI9VkVAt4BApl4gSXZ9HiCcutap
RT6cl47XKnc+Q7vr1Hnf470QG0gSy8m759z+8QTrW5rbp2H+FujF7TPGhpGZ2KCzzKeikFk7PCwq
uxpJH0G0ZzHYeE7g3cHfF3iRNBZATqsaPEolE2Lo7A6tTLuAn0yyUjqQnXfgBCEyr8dx43uhphF9
fhwlw6pUv8GU6v5YPDdHXHSneX/afAplM+av/FhW1hi6q6ONpYqnQ8fkLdKxDS1SmIWXNJ5vtnZi
kf0SYJI5sIAIM39Ap33PJ4cb4IlUYOv2+7pp2bW3iZ0wLqOYPQFnr7NXgAFEnzAFvjmtqVBBJuRK
gNEJtCm0hQ4c5GdaE942l80Q/untZyjahxK+e+LG1N3TSLfxV5T3XHbVdBoMkLew6M/ZMWis2u9X
ZpwubISGOB7SucO1TKBKn9IV3yKy5kBmJQxQSGF16lWLGeeTP7yzSoKUtK9qyqeOyCeXUBAJVlSz
Nj1LjjDJlRxk0do17uVU78OmL4LBdGZaRqEatx+mc1AN1/fvLKFHmqm9p/03kA+HYv/j5onAmG8z
bYnmQN4UdpB8WehJh11wllGnL5Ko5GICxKBEm2+7MaImalozXv/+K8/yBPfCYHYdlrjRmfk4AAKm
9dhaHksWzCpCJhY5NHnhJcxFSuQDnDHg6+ENehFm0ix2JhIwk+yYQ7Al0dLB7YzBWf9EsyXLAZjo
7oE7WjUeKDA+Sk2IRe5KPcaCB3rorIl8PWnIvj3SgunjpUBFijWZgyQlwyG9iMf1JVuBVmuGzMJm
ScX6tW28CeorkSbmTUsHh9lnPkNcP5aX/ezKW1ifoMCygkhO4JuDeE9mzThRJG+NhUA9Jf7s6Qju
+kXOKn8B8c1tFxjLQrZtAXgeYbhfzfRY2nX5P9mZv2zGBWXHJ7K8gNBGPwyOrrX9w9dPr06ITk74
rcRgv1wjyLM5hDVqrP7MUqKxND6I7Yeg1tn9xuosHnGvoQDD1O5o8CB9xmzut0Hm4tZpZzV8hlzA
8s52p3NfrdjOv6CtqavvUAvx9zb8dWe5hNSAyABoS/CgYqdJjv8F0y51vNF93iQXn+c3q8hCIauk
laoL1F8E6tFAiGMrZmlFvPqNhihCdbX7iiAxCKLh5YGJGojdCB4Pv0CQv54/l2gt9//YQe7t5HcF
uwDIfiz1jWwcPSsoGMo5Q+wqHSvSfdFhvx9s9WTzozDAmD0YfvCCUIV2O8iNeeDp+vv5w/k+ZZqI
rkUuQX0EVRGOM/dVlqlJiqECKfv7J6rZvLTNLgGgZNHpIcUjD22IBzdplcUkHVbgq9LEDmr1LtDe
XTc1rrS2Z4oc/VtjSFNepaf959d0COuvVUeUIo6rOcrGloV21bVXSlEb3kNHqNOwlKspWAAcZNXu
iIJRwEypDc6EX19MMraaJb2GWHrae4riE6CSWXpyro/3jcBa9V3DY0xvHnTRdoqNmrWYXq2Hnb2p
nS9MbfXgYTM6/0xekAnoclGViNQK8sDRClMrp3JF8JiMkfIPjbrg5f8pI9mVY3F8LlK7yoJGlILP
UxSHC+a7CEuyuADmejXSqt8VgbQ5mWM0gOevJXn0YZ+njcV0qZsy8vLHY5+yOg1R7MQbSm0F6Zkk
aheuCnWeVImADpjYPsYoNOoVLI5kYQ7HEnO28Dyi+iz9iEgpRUe+OIy7LtDnTN9jDFYk6ZcG+UTG
nOHqWCWkESrWih9FNoK7ohgSfynt9xK3auIGqKXJ7g97O8ZAik+zmcQkfwUu0qhs5e2fyzCuIq/K
gPqQt0Fz72Vkys46rEhNUtY2Ccy/M0IPC3b5jUyd0UjHAoOEejmqwt56APjalo3phFWf1bs2W0Qo
Kon79kUq+WxY73maC4WlGIWx1aw7FYT+9h/LfKwKroAwyWzG/B+B/oehQWXOTQkmvn3Icnj8FkUu
B/sBWrzReMdul/9gbgVQsmyYQjc8k8aFxNG2A0OiWjtMBGC1nsBgyImkEqJdOAHsIYA0AMqdlWgT
6Q0dv0ALsDLGvDEfAKmDnDaMmXBgOcLpwWC6Z5ODyUoirHVtqSc8cft9AivpPFW655aiHBSK2O35
0gWJqKxPCs7S/0ty+tv4KeboPH/fe5rk0p4b2fgcBdc78oejAzZ039BFApNFapOHjTnT1uyc8KV6
4HAwR+P7SyV9PRGGpS1HfkESLR7mbP4hJqCrSeKCFCaa5HLbOof3wUyS74v9riroAfZONEtV++M2
V5d50dDfAlSeQeZk3BM1f9IjMUwthnlBVc9/By5JZAf+UxIxn2Yvyg32F5UQIGx3NfwFk/TPAPHD
ZkFA5heZtWjSXrGrBEn3yRTVnnSTXgTWKn2xa7hUWJrdgqx+I6cFHE8wOYldTLQ54ONMLIzEqGS4
+X9zbVx8quRbLvrmeiHb34Ktp/j9bLVxMKUSSR5PMis7JxiEQJFSYLiT7NHQcRvdTl8NbWFG+w1r
KTf5trX1JB1rjXH0u6IQHAb83JBADvV279cG5vXc5y79BgePNQ4uZ2AEp6OVhNdg6oTvUAa4tWN9
KXu8Km2v+7L2yHnIia3LHSQOZPzRKEYmxT0hXy5yg6pwkv9qQixf3GF51/YHj9tLnLMBpAqr8vcC
X51Lq51doKLWlpJfql0Fugrb33qx5Ea1eEjOoROSpdu+zV02GYC7DJg3AsOtKKOkvchS90c6ywV/
LF1UfYs45o+6Ukc452Lizz+QYptouZjZas4miJEJI5KpYsLESHmIlHQqSX3xmxLTcxyN5/MRIAfP
ZsajfjTHghPYL9lGFdh840wza7OJdJ/KmJ0xio+fGmdL8Me6zlQNgROL5A7GDvpEX20Q+FtDAvZR
CyrbjIuGedD3N2u+yVZz0KSWCeEnz3OsmFScgpJeGTZKHAixGyK6wSmaSXnpNS3d3ru56OYyAZFr
JosKo/f272vysYeaGD8ckGI8U3XwfW1WbbCLKjXzHrQGlrFpO4CdiPKiQ1pPPlWr7JiRgsc3Rjjy
S2+P6ZyaN7BNZ49f19LPiAKzhYpujPeJkf+swS7PU5MXauDQVqzCprsX6e34RBeA1FRQtQ3xayDc
z1NuOgrrE7DTRpljGSXm3ASuQ+5nf80wenu8t9DNYLdSDxHlCZkUVHOROCh4PZxBTpy6k0uYUOLz
iCkHlWUg2GBxaHMT2JzxbSX99Li14xNCu1UJXG52C6wNyAe+iiZphN2a16WNclVjUFUJvD8zJ3Lb
R/3ja3+De9dMW63uWKiJ+pGZb1h/EF75B4uRBUMPVEAJdeaPkyAliy32G3k3dTVj3HZ+3Tbf3mlX
ADDhp7yLwGOb4dpmvpXuBln3kEgQD6+t9dBOXrpuoUbBO4heomE1rXKnX0EssvPXsd8TjjlDX2S0
1fJpK+dak5DoiMQtVzRHk872BnjVFMAi1akFci1dMcKdcsIWy2CRF/TB3+SU6pfYqac/PVqWqqHK
ZkkgFKp/z5AlDdYZpzifTiV9BpDWhk3e4ETOlJqtDYWru4jz6MKMADOHQGJdwOLV1bDzD2qv1Biq
F0H50O7rCnWoPNG8rhQ4s8uk3kbRv4KifqNBkx9peZikcwonEvk7qA+dkOSBDy1YSMQmYAfxH2W1
rHxX5ETrrXIUvRz8iiA0YqMqGNsSbuvbfN0VadMGfL3DfM/UzNq5/XHO8BiOsKo0xWfi3E8Utonj
z1T1LldZd9BKLbv/OWkpSwb4AIrK+QZBbGWYUNtwVeIYbFP8xXrcN+mAoIVISkgJWl2oAfeKvdIl
c72n2sPzy03tI6o8h6wnLZOv9SQ8IQO1owmOq79i0pnwUfB4wosfd92/+BbAod1hqVvKWpttNaGd
LkCFkRtNkNfDoOeGCoypn9uqa597e8M8k5Am1krsu5NIbyQqRudKJaZ7jkumZ3QVdaqvoLMGqNxU
KwtFXUlJub8DBqofInUwv/v/rXiqusLm7OzRHGIqpVl1ajz+gcHsVlscmRcijBNAVhw1BLqALHlb
FJdTPhn91MudbmDrmCeZKOIFZ3R7aI05CbFRUptD6mbhRiY4TR2Pgnb2KB8anoN6HpNmri96EswT
2ScCZhPWM7NDym+JpIr7T0ifon1KTi8aWNsz0cfD8mA+36UDD+O5GwBw4GDuup5p66RALMob5Raw
q6wmClxotsm+nVh1c81psKOOtwmty/YDWRBdxSsx+r50eZP6UearraE/cOpydPH2mn9p6ewN/3+Y
ImBywuB4nv53jqPx2CEtjmFyQCpTQCv+EO8nMfUifflTWct5TqBVwyJYzfBS4KwNm5epwyrCMLIx
wBu5O62gqiXZe0El/nJlYCaJdIkZQ9b3jd2nGN25IMZVsWJCC0esI7ffENlcn6TAnyxZqk1BHASe
mETJiaNXwZn6QxJMp5MAkQ6RXXSi8qYUK+7StLGgAkMS5QfWKiPheamUkABGlfCH3aUZWHrrHHx9
w9pWH+HcUwbCnYGvLrOdivNx7z1TTiVzF1WJ2joGLK+SohBU5+CDdzpbm5MaHEDpCBve/E2rC95+
qvdl1PUdOTJ3C0wXWvQh8orI9oHwGuUqFcLzWcWfUDiVJN2gImBDci9+pGs7MwuSis3a59nk3RcN
Ld6gKydOZO5YIh/s91e8NmCrdNkYO7IRDDBwfOu9KrLkmjVaOIMGGHQIqK3OBFW95UCTJJ4a3oxK
v7WZ9eRFvQaMTbIdTOjBlCPOWvTCfmFEpuo8hBG2uAKl02JGWaFMeSJjJ9mQT6fY9gv3KjIwl1nw
VLUr7UP8dOIMzc7Wh0BwKbop3V47B/YFUC98Kp5noUBblHUUveJS7sOdX+BX05hY3b3kVu9uucvj
LHh0xOY/vRMeTTi3cR+HkVT44o19ooh80gc1alIGnCj1iFekJn7Gw6SfrWxQGBteMvRpC/pyHgFV
x/wUQnNcuBeRCgT7FPLpV73RJNtNOkQTPDyiszI5mKd2NwEwnp8spZDXTuS9NyW3PFDSdHinuh6T
vNcKM/67ooGvoSBSIpYrCbry0bkDgH75am3I2ah00Xqs6MiKV1gtmpQNbmqpHTAypqkbG1guCltV
8O98gFT7gcOjW5hrQV5BQTDMr4grc922CT1MMG8VNX5tpsRcGz3gUu2szBHmffe40tB8Rii4AJi0
2wnz7F48kLcnrnQbaCoFacrfBD114kqBXZfS1D3Hx8FDnKd6+Hfhv4FEj8D+WShm33NVe4yRYrV0
RoPo3DOGsyPmFjnH8Ha31hzq/VN5alTj/C9YRPWu2G73sdiTMIiD88R726en/R9I/otm+2aoHqaG
GrScVdEoCYzkv0JjeAHHOv99c1MkoLLwEriPk+ZOC36/707V5MYYHkprPBoJJ9jYtOyOt6XcJ8iq
2rNks4k=
`protect end_protected
