��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���?�;ENU��ڽ�/ı��Hb޼��~H��.�d�g��voԼe��H�'�����V`L-U:��9�0_�=_��8���rK��}e큇���un<o���}��vH|�2�?n��r���iq�K�Ә((���o���Ę\/��X=]x�	rS��4��1�<��F<��/}��+�F�j�v������7k� �{�Y_�=U�,��93��.u�̯J����3J@i:�Ȧ�O-l�4��G+U!���xH�?�V0<�Z,1���
2�g�׫���%n��A�� �w�0��i�E^;b(|�	���� 5su>r~�=Ե��a_�RxZ��X���<��Sr�"#�t������%M]��3��s3AQ	Q��)�3;tx�G3��)a2�-���_��^[N;��yC�{;e���N���ʐ��
M}_`\�#e^�8��L�2�+ﺱ�xѧ��z�Zs���I(�����"��Rat<��mM�(�}���Q����e�� �S;��=��1<x����<.3�����x��i8�q������X��=�y��y�\�eI��o�E�D�b�1�ax��Aq��* 6�G�+9��_��݃CV�NUȀ�:@L�Ѱ�`����Z#��?�/�ϼ;�δH��az:Vuh��6O�4�V�~��]v��&a~=ƥ5$�8=v.����/;Н��!�Y��y��eR�5���9Xt�jN�V�oށ��,� J����"ro�1������O>���f��vFȅ7��@�tԸ�"��ꌽ����O��W}*�o
��uR79' �m����\B߾����o��&[Z�xK���o�R��Z�j˿�Se�4y/xY-Q�1�/�Qدk=mlVO��fO*T��a��F���-��7�Dfy��z��$*�0�����Hʳu��kY���U�s0S$������;/��pF	`�4��$t���/3+t�+kF/�$Q��
m&2'[=a�Ýq|���c�q���ҫ!̺�.�����66�c�aj ���m��at�gU� x����{^�v8g:fL��˄���H�g!j��F�#aI�;�b����g�n8�0ԧ�#�DK��K���k�O�g��@+��R��W*�Q(����,�&L�A����\�t
�h�A Az3�-��-l�&Q �l#L>f��Y���Hz�S���H�P�����b\�R�����e&q�&��XD��ދr�,�=�%)p^.�����&ZM������^��	a'Ǟ}:�j��10�s�ԝP`�Uh�"#���9��kRe�Ƭg������FOf:�>�>-���se���je���o��v_ŎP$��F�UJJ�ճ��=;�by���X��E/�8�5{��t���C�A.�s�9�@)��bz]��~���W�$r�*�[]�����I�i��
��hkd|QqY�k��2�<�®��2�h�}�K��5�Q)8%g�B0
��F@��G�kg����AIF" ?�z�`i���^+�_Z�ǙT|�ߧ!V�����3(mM߫s���޸�������(3���֯��}���q��;�b�A&.h'N�������"#����@�7�X��TOp����+BԴų=X���5*�>���<�8(�O,Y���z%��K���bE���!�d�4+q8�����Z�響��13��_�9���u�ü�U���J��r�`Q��8|_A�F;�11��yt�T�GC��ŶȇA��5�mٯ<��\�6d�ȥ��sY]L	�p��j^��_��RN�LЦv���A�-#���{��C��'*�X#z�gh��GzGҍ۝4�M�F@�S��|9kq̦�m�/�;��A�Ǵ�Hd��VF�-�E�����L����XT���o(��nh�jGR@���n!�_d�ݖ�?����/�S~_&������Au��V�e�R�P6�{�(�>��u��XU�	#\���{i��؃�8��������_��O��%��C;�P�\=_�h�@��!DG������r�㺌c���%}g����E�<�7*�Fz)ԧ,/P%�'�Ǉ��i�a\��R	��|�
ͮ�Xح�8�K4"8A��8��=e�:�}�i���I�f�u��`�0�d�AĠ�p�A&��CE��BZטUw����ƨ�����[�k{ݫp���A�¢yyA�J�瘰���$#�n�����&��K�AB��J쒙��Y8,9,am�Ø��s}8m��*@�T�p��~�sgJ�1�`��)WV[b����ř��l�g)��?]���G�q����'�����|k����U�>���FZ�Wm'Au5p���!#�zW+��/��<c��b�&.p�R/LO�(4�]x�bc
����395k-&=-�?��z�׼&�.9�&Z��[�