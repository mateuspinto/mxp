��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���_�Z����,��������+��H�<h�����=�'j�;I{j(O�yoZ!K����J��9�pa^`��.p�	ߥ�7y�,M����贶��j�yC�?4S$V����@�SQ>��'�H��,��O�N�7-uS��_`�^Hj��5i	+��d�ze�3G���dpu���[D1{eO�4r`q
���
��d�Y�O�Q�"[�]y$�CԈԊ�0�?_�ޮ�>Q�gxtƫہK_���8��pwzMI/	>#4��/���d3��L��v�%��~��@��;��h߭�*87E�+�#f.��@kE�ڠ�oF� ω�������9W���[Q�b���T���} W掓���Aдr]q����xG��I�êR7d볯�{X��N�.�_�Y�Ob�F3a*�Ï����PpW���NZ�k���y*j>O����s4�d��5o�`�qΏ�rx�0�vq+�0,M�D v_������M?OZ����FT,8b6�F&}��W��;x�yg��Pno*+��;��r/�He>��4�d��m���&[ԯ ��	�'��@�3�LC�0��c~�5ș��p�~dd8
��c�1J������8Н�_��5�@�%CІ��ߨ���_�) �4k�n�% { ��,Mۆ{��Q1�f��\�|�d[}�>�ҭ2|����YMa1f>�UC>��Ot�
o��Ğ�q&.Aq�M	�ssA��ri5��M��
�7�l,6����\ ��^�����������>�Ӈ��p4��  L��d��T&}qK�or���j@+9RFx�'nM�y��Y1i^ۛ�8&Q�}�n��l�\��,���!��"�/ݥ���ф/M���N:��	D�hv�-�?��w��3�W]��(�]Ȓ�k㜀x &wH�=��y�����Y�@C��i�}{��qEu��[�=��}���!,^C����v�|V�'�k����߰	L��2��.=��u\��a�E󂅀��U������>�%#� d�JqFOo_r�������E�uA�nj�P�h5OUE�}����`�ܪ+�:]�#��ݓ���hT����!�e�Y���孳���=��_]���Z���27)me�Z�+}�����5�M����w����ƔԴYC��iw�:��/��\;�/�<yI%�x��.�G��l��QTX��d�F�J���|в���'�M{��=�@�;<�%N3�hD<�,2<��W��L ��z��S�{3?bٔ�}�V��|:�=��ѫ��uUY��B���R���$�l18�cl�������d�N� z�,�ǳ@�&�;a��)[�Mv<���q�ʇ�'�+Bhg�v:#	�ԄQ$����/Y_����#�y�~��Tm؛!�+���DC�nflxm�t��7�C���������%�3��Z���ۜ ����̆�ز�mL���t@��� p��ܡ�B�;U���;�ʻ�{�M�܅{\�y|���=����E|nN�,�6l5ws�gMP�;n��w�&���j��:�㘞���ݪ�u�2!��lW�߷��"Ew�~Q��v=T��e�x��I���K���#�<��Ŝ����o��][V�S}/2�T����`Ψ�IF~��2�	��ц��kR�dG�vt�#Q�/:)+�I>���=��T:1���劬���l�� ��� ^@���>��.�,\)>T�"�]�Sh�$c��⭠�U���=��wզ�<(��f;�M���������c=
@}B^�E�������郃�����/�L���U�/��v<��ġX���v[�4|��/�`��xֺ���H,q��Im]T[�m�ڎ�;�"M�<�iy�_A���ss���
�Dt�Y�iE3f�/��E���lI�)Fl��p&wJ	�DVg�2���ogӵ��KH�=a�V��3������S.:���l�`,o�ٛ�,�J6��
gZ���J�[����@�]�4?g%����5fTG:�{*��;���vF��_�D�����g��TLs\����.�`��JJ����Ck�h�z�b��K�▼ҼF����f����5��g�M"]�L���L:]"��CК��P��rEX6R��M���pF�֏g6G!>����M����ǵT�J�c8��)���N����!!'�a��q5�W�j�fw<�Dī���o����z
�魱�\��=</p�m��U�^������!�ؓ��P�ؙ��ˇņ��'.�R�m�\*FX�4P��7�J!|�}1$bZ{�1����,b!��\8
��������Y��xg-,�7Ԭ��o%���������#?GR�m~
Ě,].{e*ñ�ƣsHn��3�G%
�s�4���q��y*aB�'�Jv�o)�ɡ�g%���J���Xp� ���1-ޤl�� ��^������a�F���?�E��>�}h���i�Q�87�;�	�YX�Y�X�WW�S�Qz#��I�[���F�H�1���7�#��:ޖ�$du�G�Xkηю�*O1�O+�/I��oS(FC,�[h��r�p�&2!�A�)�.M���c� ��+�c�����-�B'�F�T�Z5� ZW� ��s;W�|����x�����.3��Π�+W�KA�Tk��^3*�I��#]���
�UXڿ�r�|�7��[E%L]����aw�^�h���U��}���扻m��vC���0�Y��ϭ��pH�o؀U�4ERM�m	�|e�V�{�H�@��ecL�Z��*�>i�7��8'�M�_ˏ��Â�\�Q��S�ݞ�����@��h��%:3�diս���}m�^1�ec,Xo�Rz�4���E$$[6..
�1'���I��zs�BM5c�^���B��8j��<�F�p|���{�;/��0�eSx����I�'1*������~����е�,�v8))@ �/���.�ə��~8w��Ww3�W���6����վ/JGP\�rM�Gw���u@#q-^���f4^=?����u�^096�ن�k���VK�m��6hGE�K�v;G3�-��M��%��d������z�1�םܑ��8����):��P>��? K>gq�}V�D,�6�I3N��'�޲̗�!]+(��&��
�3�5������L�T�R��ы�'�BkQ�S���We�MZ�eƢ�� �Q1>ثٍA�������-����܀EA4ԉ�Y�]ʟ�ƆP�-]�W�⇮�*��v��~�D����F��0���`[ߦ�U��#���e+�'�|�S;����I��/1p����]�+nf�[|���f >����B��U����频E�A�'�k�r��*����e/�&���ۍw�gP N,[:j���� u�S�ڔB(�����K�F\�~1��L_��3s3���	0|�\ٌ�~6�����,���"��b�����@���ElF�Ư_ZZ�����s�L��vA�B��ҫL��X��!���vsQQ�ӓK��ϩJq�I�����o	+�A���}��df��o:�f�&�I�r��O
�zO#�t�� ���Y5�˅$���:9\anu���i�3�^�=����G�d��z�!65Q�G��u������14���_��G )�W��6���yP/��Db��+���!*��6��;�����
[�Y�<cz,:�T1�~^�8M+=�q���2�=�K��YR<7Ýo:�ɹX�N��QA�r�z��1
��I�3mߊ�b4��yw�rT{ `0����>�՟4
=e���vA�B[+p?/C�	�ń�-!_E�:ڿ���ޕ��4���5��֭ �T��]Ǳ�����D�9P��WlF�����.]=�a��z��P[���-O�n��w��eM�ߊ��H������w�u��p���WG55+�F�1X���A�H�>�->��$��Ν��}����讴7^�q����1�žiO���a�q�Gf����ޚ��1�M=�.�����|�JY�l˕l���RKX���N:%���N'�`*>8=�ָ��DH׏Ι�j.�
߇ u�X�]��
�@�l�4��.��gą�@�-��>�U��?שL#ո�P�V��(�<^�~��*V$;��SH�	1_����u�=2��8�y����9���£�,#N� m�ϯ��~�&��4�;I{㘞�V2��(�^��|�ك3V`�g,��d��'�G�0x�g
i��F�ZҘx��B���T�WF�'H�4��>>�Y	Y�tU�׌�Up�,�G�h���
���o((IBIئ�{� SK��º0~9�o���j�v.��� Q
���m��-Bp���:�8�sɜ^��":��I�TD ���}�����G�}5�W=Hdz�x�^8Ğ���-�Bt�-�����̹Aod^l��%�VNod�E��N<j�b�au���r�HfmD�`�9�TN��X��J,�*e6��l�}�ɤ�Hw�!D��R%�^7�H��;�g����G5��m;�${���Z�iā��]��3���-Z�C�0�
9��p�܇��1^��{�lɒk����I��@X��{��O���)��a��E���tH�{�S �"PT��)|@��qF�7_���j�H��d��[���x��C��~���S��Zz�¼�*�ĵߤ��S � ����8�D^�����è�ӠPe��IT[�/���=EF�e~�k~���|�9��g�nt"�Z�G\�>`��l�ۚ<���%G��O��@�%����Ae�#�0�a (�%T4h:���A@�HU)3g N�{��lW�qfF����ي\�q[vIb3�~���\=�Qu��H�]~zoIJ^�e���F��B/��c:�;�сH�O:��H{�]� %r$����u*�MZa�bv�ūhГw<��~8�����0�j��`y���Œb���BLG7�,�$�M����aF'��R�7_"�<l�;�Lh�f}n��>E��d�~�E�4��TBf���k��'*����%_�{�C�8R6^Ld���@�#����眿0���!��l�Dʾ���� �����f�<��<�&�or�G�jF+�0�4��=#���q:��s)z��/�U��T#>C�뿅����$C���M��1e��q��x8x�ł0�\6��X��=^������/T�+����/��fp9 �w٤��Z�Pz��6�����R�o��Y��Ptȓ.x�P|'�6O�%9�$��8���L;�ؐ+Aʖ�Wń ���!bc6G�U��<��YL�68����D!uۙ�M�MyzG��k
�����l8⚮u��A���:�!��d�1��_�K%��wC�_Y���oƥnڜ�&O����;�bҘ 4����/ ��M�Q�0Q��y��$���^���iL^*�7�������hֈ�4:�%gP�Ԏ�EK�e��Qr�x�:����pg���o�7	��i��G��$Ep`�`lr��Yt����g��8m���>H�
P4��8;��P��\F��Nw�NR;�������'S_nR���G���V	�a�ё>�K0<D��4�#���K��mE�2���*#Y�$'��줉A��o4��V�mN�V5��?N��r�!���W���FHUG^E,�Ih_��I�ϕ��/>a���|������mY` ����!B�S��*��i���S�p���x*:�'Ǣ#9�5���n�rlC_��^n.o�$p/V�;���}w㷕_���9�Nv�Zh�'��r+���y苃[��2�㘤����1ԏ��1�-�7��?q��.�|��o�f�h���C���<�ѧ}���e��V��G�We�5�/�0�EN:H�g��OT&��:8��a|�H�
��tPT�����u�7" �Ɋ�ݔ�8�U��<S(a��]>Y~�>�N�Iz1+�S>��~	�p[��b7��!��ùwF�B{���<� ��m� х���Q�081q�mw�������x�]�z�S������a4�ce]��g�Y:�Mf,�(�by,�gbHG��n9��.�"�+QK��4h� ���h���S/%��ݝ�:��BN��1�?=
fN^"�)n�d���|��׸������?r.�*V�*��Sgd��Fa��@����mYp���q���}�J�2�htP��L�姮B���Xh����Wwv�n�Ux�xHIo�9F��a��=`0�W5o���$��a��������V�H8��J���U���FX*O