`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4176)
`protect data_block
Ds4I42tdYrbq4x7SNtRe9+INTH3V4aJAteCi9mZTQlZShC2W4yzZXQpotL9fsQUWA9G9tIQjMCi+
DLj3aDY6rRRwKQ/a784E6paBAoh7/hovUpLJICWa4tbJ7r1g9/tI2NRINI75h+60w1Fns/uDyhJh
Bno6y7e5P33SVj7zyYfn9qVSjeAdx7nGJXhY9jGU/QXNTYDnDcTlpG4MfNYgpzzT3QdKrFD80YZ4
YVxv81EcuUSSKEGo2UK+zg5Z7W7wL13N/iJ2OLx/tAoOM2CNEWe/1xF/Zpxh/zpa4bdgE2xdoFJl
38MSSaTDfMyxb+fTs1L3dejTrXH0CieOpN3EZWsGeUjWsh1Q9xWmC5foOTXeucop+uWj2T7YLjSD
DQn0V92XYw2NoKAH9wh8/RWT3S32K3PBQ2o4kWO9LSuMSSA+NoEFz0HHbabKM6VU8nFCiY68JHbD
JUuUR/XmttiVVBO5QYp2soIoDUAWW5hQ+EgdCLuydx0zX/DzpUV82ULEy5WR0vYY26Z30QeuOeGF
1pMM4hm96/NlFypRQyYI5SJ72p5TqWZp63gI4fK34MCw8Iwqn50B5q87toM8RWhwCCYQdJPrQs94
LcRa4JFHyKGSHrtWzIMgIV51gjdVI8xr8nrmWWsnv83dGiJdvV80ulBk6ERh5IpiadiWTp52fTp5
Y29aXC87+JS2p3hn768KV6VTrf4qeQ8GmdPkumSwyPZPHKD9i2VU3+17E6V2r/I/jVfhxr4+XRhO
R2xzoKifQ4O7ZKlqsmcoFEjSZn5jMkHcswuVm9C4Koco2cttNW6ZHWtJ3ivGf3E+M1IfQI1OqiVV
OGcraxdJYLOujfhIoS6UoHgqu4YdzG4+/9EH+MZ8URJypSQPm9E2PXxyP3FINyrlxzL9Bz8vAuaa
PpYIAuWmkD4qqSHo7RJR4wrOSGfN1O14cBy+wECJhapfaDjmklYXvmD4QOB+najLQFwJyUAFC9Bm
Sx91MHTDjOJLR8jXR5ojHTP7ocSeakLYXCZ+YFgANJfmVRtExIN9LsHCne/wTvH/amliJevTn/mo
430fPXuCSg9+4wMDP5nHe6dCQK9gAlkPbuebJ4gidhyGsi4gfHflUZOMGpJqIB3up3U9kbn78iec
ZN5E8uQZcEdHPZZaiCuEaVQaWm8UtWzVmKhIelX/H4UZZsJf1OlLYH1pXZyz2pztqkDOjnxO1tz+
Xwu9obgf7MYeyod12ZIK2n+udVddA0CT0KbYHi/+YHpfgNtfKfGwbqNZGzpIiRJ4bLNMiavfCOdX
2yNoBz+wHnCmdzMWRCc+xYuSO1xvrLyovNGeMWJe3gsGb0Oz+Zo6+h3ARdR/aRD+1xhGtfI7nbLB
vDYOLIR3Ceo8jfdwba79wJcpI2ITYliG+t6jdFrB4wDgVM7sBZXYj1WqLqwzovd9UTbM4lqixXQY
SNb3m+oPj6gQGQS2wAmSdhXzcDDGwjtNMRsQ6oyaTStLkr3qrmOSBS7dilQnG92ClyAHTBl+DIfe
N5XXfhwBAit+sdAxUunxmyec0xhiKHcE6FF5oh2K5JQSjZku3ljXOcuPVjC3sZ6O/CwszdI9hYqm
CTmfqgleeCUf1ib1wJstnx3CJQkxgdwedkQKbpXxpTXVDAY62EoYaro5XIp2KIRHIwPJeUy1VKZU
4ZGhd+20bVhEh+VAF9woTV7B70CGiPHSbh/7416EOb1YxVA3+5DTnsTH3iRUevIHeZd974gnoxME
ldmEFyiFbtfY/1WUXeq7SwgTaiiCzH1niXdykM7CnNFOkw647h/nNOwE7OudlHlnFKGqvidS5mG2
0V8U/5vORZKElEUn0uEePCkMr3wBNWYUEmeg4QAzp11Jr3nXqaqo9e1EyRzVaPSVUJUxSPXCWH5y
77OiZdrVtRL0i/ULqGWyt1R7J1pIsqTDRfjWkC9xuv4p0C1kZ1p4DUxZ5BcP5MytwBWiqP0WB2xE
ciaxdiKOwsZB3hSj5lurFpAxQx0+cfNMC3Mcjf25sz4YnoY5Pz0UdvOq2UJwFf2cNj4IdZNUGbSy
wKUJtQQ9nibIWiDRDoKe92Cdt3xjBLStJj9EqhgPKtwBgAKlvq9L9rOWRpdz8wwO2cuEKzJMOKLN
sPpXybC1IPvL1XL0YJjl2ub/oeN8DM/jvMlNZ4Iz6W62U8dSO98OTuI9Wrgwd1AYYWR8gTFBAWMU
4nVe/BjcyPeL5Le247SWQMe8Trq/PAq+27I2Zyd+n3Y4ZYWvJDJ6oK9C7nqqMv9DJDg4r5JDTn7T
CeVjsO0viS2b+myoLyPrmnsPk6i7bnOityfOcY4+Pj8mBK5VzqlwMhEuR7MwtPDqT/aem2lMY1+D
n6kM+NZAMEGHfvbfp0RCN3SwQYZgpwQGPwdjJC2LzKm5p9uIP/mjDDF8AbFrET9ZOY7G9MwICXZE
QWzjZe35wZY4kjD2A+O/he/i1Hm4/htKVlmpzunlc8PLi0HE9C5t0L1OKQYf0ti7ss0xGlvQ3lu/
8HHpSgB3GP2y3yWHmfgg2i6Z1W69HKoCSwsV0rmegLCWpcBGHy3tZudxZdU6E+zxKZJF76u3rlsX
Et1vPCmOdYyaFTJsZ/q+hHi1LKqJQLMgwdyJs1aMZtEcVhs3ZqEYccQTV18TIuyXIHUwZqTZ9xQm
nOg0RihowvLezGdcJSrobdfcDBH9oykldr7Sed40Lh9eKHNSBy2Mht+6YCz9gz0mPZkxUf4pOcQR
1pPXJIBxuOWJ/dJ5UtHbNQ3XT3YcqoyvTV2AmtHYFOtRpxmCUuvx3EErQ4buSADW2AHRVrEmTFxy
JZI6yyS4tMufUwjDlFEIRndk2wszSel0dHo/T+smTDjLkMdIXc7dz9rLoThyQQLeKVIUhCpZd1zm
+RDKpIdjP4vLw1hmwbgPkJbKd+jd3diyQZMME3mQyO13ZKgZFFOOFA9xL6Y7PkjRGkDZJIgkEZbY
Iuga6ECzJ30708EHaisrGTPcTsuJCpL4eKWmpWcfSj/PnHfztPHkb22/190y5KLRS97v6QHVfd6S
tJRRa8hYYuPDkak6VzA0tvF3xAOv8IAtd9YwUZoWFvhZV+z23HoJ17UlC4jV0o2PnvwMpXzkoiY0
AtfO/PknL2snLQfoHJ8ZVjWijPiOu9Ws7T54q9Bh+P5dJLglyERN05pRPi5aO1J/859DqPXbPeim
VE6GReW1S/AHVh2cXwcZ7/xycC5L3Z93r9ctx6W5+iAer6ZWkXJsaXQr6VjuXW7bo9FiaVgzHqt5
xaBMkZ+VfjlkFOu3O/T2j9ZGprc37KnxRf1Hoa1KJUdKvfa7RboW0/eHcZIC3tRfKh2R7VeMwVAk
ujfxTAA6hjmOSXrVYYrtIITEPxznCi/nTwcmpbzLyLsYfNG2JeDDTB+hPnnENoGqT+2++KOFfd30
+6AB5Ruanc0ILPVRP3N+Zj78ZvjXXm0twF+he+2Zvfr32s6pv3/wEKDhP3/A4jNAGg1ocfLtlzhA
yYVDfwudJzsauc26QROiwYa7E0fur2744p/+EtJrqCGgaWmhiKdgaSA4/dCYeStjFOUZWYxcHWqf
dqEDwM5hVzFjTl/PcNp8y5WLNVhp3wdIOQwVx5ktM6IM8Slsna5tMEwo31dOOTz8nTdrLdNls3oh
EwxTLrw7rDxFNiCGTxgFIvMliyLQiCIywd0+x7vDIMOD+Cb2xsQnKueqCcRD/w0xzFbq6/ZKojfh
thfAWWLRm8OwPH7ntc0Cd+j3RylTSvaU4FEvk2ihz2XT6UICACe5CQA0M19iotl+3q0FPL+CesKq
Zy5HpllI/2Fde+7meGwfKR3yStoBXwBFqpbzZySLQ8eqrB+DjZXr9W71jW+dJl5JOI/q0GTbg37n
9HEK+UBuxhEVk8877Rp9YJ/tb3mslbCRYk4bbIGGhxSz7RAWsLBqM85ib6mZ03M1hqS9w+egkfJr
PZxskdFVjlJZDnZYxhOXXuKgHbb+A9OizGjqkOXBvfnJ8+5IBcxGN4P3iYTxRVzFx0NcRXHDvfP5
NOaFvZUSPU2b3ta08pels+zWQiK63Yib2LspgjeA0niz03ltAZJ+m3h92Lw3MWq117drF+Lm9fLe
ydTz38684PK+BF69J0FhstnDwz6DtEZq/4VR9i+r+vaw3vL2o5L6B/v9V8bQrA30tHbRUSnsXjgm
m32aqsjytJtDh+kkuZqipglCFWheiWjOe0IsasslN7rqPiZrY2Ob7i/LQdhwVUXoSckLAO7+63z0
MiBNCQtCfJZK5HmZWOZhsNlwG8b8zzxKbmeBx2Eve6QdorTkkwcpV1M6SJ5Q5VpxWqjv/qNpER1J
4tOMEYgMUeGjVK3uNy6bWCYbUmoP6xAOHr1ErZMF14r6UKnUCy4DHpOsOtHaUnjACMzbCEXhXjRw
7A8C7KXLmaOvUUSmsDXGZdgE5QIQ8hW3HklbU2sd1vuUCSMLiq+O/2c1bexmnA8D7kPJ31/dcCd7
IPPSQM7dU6KSohgdFoYCtJ8gSQ3PSq7fo9SiN6iDyELiDpQnQIq2yzwQOhAo7+mpEGz3auLal9po
Qh1dxjvgZ/6cNDeXRHG+khkcaN83Rnk2b07IRu26Au8i1FmuUqXlBAlV1JpCYeW+qf1lSaZz5vmY
OdrechxTYgjkvqBboFucBInRDSbAFhAzHi3MtI2qwcbIfRuI1qzbM0l8tBX1fOoRcu8ta1CT04Sv
94JPMzg3G5LvISTY1/jdZNV3Z6U9P6slylSrOhEqu1i0yMb6vFe/k+cL5tyHePOuLjjWf/zZo6Ig
YD757JBsH/oUqmIZI9WPmGyk2vH4kMqySSnWTYq7MqMtrs1ivANpwCAz9w9JYNArNYsCKsth1xo2
srkRxDkXCMIlKPE8n890iHx7Fi+vbEom/qG4Omrb7O4UVoMWeNz2w2uPcbx3asGPKodiEH3Ta/9w
6rN8+H1DNG71z4HM3iNJSWRSpIBWh5cCJ6UU/0QV7+9lFhSPJ4lI1FRLQ1AZ2dz/SpE2tDFh/pT9
bk+TNyzZ4+EV8M9VcLhtcGFrYjnnVrfs1jUYjMJy0ntOcqc6yR5ijuXWmST1WvnTS0TC4Peu1yEH
WnEXN66r1Qo32nT6GkvQt4kzHnxlflCCW3lsZ2YVLs2go1XmT/f0RtPVJmO/tp56J24LXkPpjwPt
9P+GM+ktwZgm12RUNeearhLpxPkbLhXsgAyYCKB/FEtRPxxQcVtqiYgYDpsbLk89fE1aPHwne1rP
4BffFVf2wy+WOX4vkUC3w65P9dMy2ekXiSpJOgdfDkZDDSaBk5CdJ4uIFMsmfHNgbCqeOIOxcbhD
WZUITMzvW9zc1rXE8jMSAze8wZ6k97lAWM4uFfO5HRzx5mtxZAwW2+V+VqPo7SROhG5slKJQZe0E
NzVkeQ8tD9J+1FKBoXRttXDYh6MjrEEV6N0csbhgmCTswppaI0R7D0fsVvePxtf+0GGpkjE4PqLH
pYrn4l0uM+obPN88lrW9RrIKeM62/pyLDk1iG9+aaO3RsgVwLIAMebGnrduwu4siAqr87uuXeXau
HXKk60GUnUHivnz8lvwp
`protect end_protected
