��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���=�:~�R�Ÿܱ�*�_3���Mb`�5�tp�������K�w�k뺃m?���.|�s��~�����6R!���j�x��x&��S�j1~bD����*��@#��Ay��Er�ĭS,�t,졃oi�"$��PY-t�%/�m�L��^*�N�9: m����3I^΂Í�����%9KO�㡎rV�y�Б��sKS1E	i���yH��y'e5�G�_��L�Np	�7�q.�n�
m�D|	Y�5����_���v�E��8O�5�SƄh�覮���ډ���Y��j�D�!�nWm����0ζ|54%pG�����)�$
��	z�y �}g�O�0�2��٦&?�ov? ���g���S:9�I_��6c�L ����d�5��bEz��N�����/]V���%�<O�ⴟM� �5ڄU���6	&��-��-��@�χg�I�N-�Jx���9��9���n���6�5��y%������MV�Qu��R����� 9�x	�f%W%/�.�a�0��-���h��'E�W<��.녉��E���aE���YC�bWp�>.H#*�9�@���_�HC\�`��8�,�+�7b�N�w��I�c�1'�X���Y;�L�4b{�B_�:�����f�.$ᷔ�!15����G^��n�^<�c�C҃n��<����)��hC8 2"y��lT�Tk��za�ɞZ�q��{ՀI#���,@����o����j*/��0M�������G�I�tʿ�_���{bl�-v��Մ��pܕ�m8�2�l��g�ʵ�ݵ\��r@��K�����{͛PAѰRc|��sA�����<��s.2�5 ���B;ϽDCoh�����;3՞��2�q�d���ǁ��ׁ����˝_K8�����N�������:��9�UQ�i��"G����=?r�O��ٮˍ��Rr�m*o֧�����8�U�C�"j��.�4Z���j�6[�Ol?,�}�#�M���#p�y3��_3�Vu�����5�T;0Z�U�u�e�;uU�b��Ƃ �d�r���δh��]�k�����#���pmʍM��vW����i*S);����.�T�5�����U�9C�)3�-�~�d"osx��J���-D���ζ���#&�^��+�UʖG	��N�?����C ��~.AJ�4W�ͦWki��ϯ�Z1&�s�L}g����'P�ݴ(�DU[�~㨟͂Z�Vc"�L���Ӯ�U�g���;��h�$�a'�t����v�o�m�5�ȣ'blvG�Q���K����� .xZ�i��c�^���ftX<k�愨�x�\���lt�\�8����Ad��g +C��Ga�/L2=�O�ӷ,�����S��福*�Ae�V H�5o'_?��Õ����x"n���4�h�<L��I��Ѓz��3R�+e1�_�ϲ$Ƌ4�e	8=Ҍ��`hݦ�;��k&��{����g�Ɨ������k�qjv0�!>P�3��FG���ER�]p[_}�T��P]�X�}"��E����e�%�EhH.U��*�x����-@}�O��i�<�M���~>��d�g�f�W��Ķ 9N�1���j����:�P�{��7G�%1!d�gPȒ�]����/����U�� ����R��8y��J|Za�.���MY�G�%ߘ2v �ۗ��R1dW� it%�z��!iqW���:�#^ �Ef��ma�V�dB�� bHipb*�;*���8WdL!���v��ܨ���*-�`�LѤ�B?Q3���@	B]A��8��\_��ex���|���8��ZE�
v[�C^��QA�Dh��7T#���Л�D��qx^��z����t�Z*��?m���% ���i���<D�m.7��R��@/�y^�WƅS�j��zfq��\��pxz8,�� $,�o��XS��h��9��{��Q�k�m���S1��ʤ| 5�UX��q����\d���-�HX�J��b���ǹT¦S��%l���N��q�#8{���5��U��Yx#�z-��� sm���GR����ϘRFY7��0��n���D^���Bi��[م�>`U-�<[����
�����B;}g:�T���A4�P��.��nP�!�32��d���@�hn[�=��Sr�T;�n��/��t�D�C��f��i�g�����L�5j�_�������� tH�aD{��?�c�6�v���(w���|�9�����5.�	y�{��&���ː�#܈��F���
���J:�axu�����~��;�/��I}B �Ϝڅ���2aǄ��Q}���'������33�K(��ض�TwH� �@:�^�j$���w��������Q����҅3�fZ׿�u\8i���Mk��3�(� �!�)�>]�{MW:������>Y�$H���aÐA̱P�V���c��O���B��x��`�讜m�jt��d��3��tpM�g��%	i�8�ܜ@��Q���{�݆����ˉFZ�(^�8���;�������ʭO,;���P,{�2QY�*��p?�@�g��%z3��w��@�������a�߹��^�\��:�FY������yy�&`���rJ� ��eX뙿"��2�,J0n�!M0�f�hJ��p��/�\,�UB�hu�߻�vVZ尾�*�ؽ���Cfi_���ss��6?�ef�`p���H ؚ<��\��K�n����}�O�˂�U(�Rz\�A��r��cJ!	�Y�Y����I ؑ�Z"��T�?��*Q~,���HE�}���q�jc�� ��ǥ�8&ְ �N�1��y���:qi�j��
�Ļ��K%P�3��MqE�@�������0@0,j/{9lQ�W�Ec��P�8�}��N��es�	�9b�M��C�L�0BĪ-$���	�Q����/ GM�7���d�z��������10yQ��� m?�q�����c�>�\��o5s<�^�I�M:��{��fnDUΜZM]�y\�|�-�6^F���E���v�&=�{�t_�8�X
�����ݔo��R���h��Pأ"�H��a�YT62�=-��_�Y�����A��ۣ�)�Y���?iV�!���:iXA�<��K��\�P/�z�؇�YX�����{~<��ۆ-n���_C���x�tp8�� �x�(��H�i�m�����ܓI� s�K�`�&b+zƂ/_����;�_�&pt6 �䏲[ռ|�آB�LH�M^*닛��)���j�pV���{qC��)TfV'na	H��Ր왛��^6��v�1&2� �Bf^+�D���6��0Ƕ��]���\hFT$�6�gQUy������g�x7�e�)��f2����oF�T�[ �*?�,�xie�H)n�Ɋ�K�1��.�J#��M��t����I���
�[i�2�3lZM��P�&5���B8�^�^�j!��r+��������T���Č䝀P�5���E�bps�-!�~-��˲ �^�Q�]�Ud��N�:bb��iϼ �/��m�߻x��gᎤ��ˍ����0���E�Q}��K<`�(��� �].p�Z�&���pp�J⏷*�v
J��l5*o��W�	�AJ��R�*,*������c��`嫁#�ns���g���vR�Dw�;'��a�]�9���:��v�m
���`Rl0S�9���λ�����%�����+�l��/�E'�&��kޝ��P��_^��
�W[A��5�����n���?#.E�j�f�}�П���ձ�4p� ���籯����ee�H[�[V%�Ӎq*+*��:UXDj��~��0�.uMs�<��#�X�ѧDT>�-�O��tI�^�9㌑N�Ă��>���0d�p��tT$�[�9�P�.K&N{9f�f�l�}�Ih������RW����b�ѯ�G��oYL�����]>�>{!?߅�D�L9ڧ6��`�ue��pf���ݿAư ���n��+ױ�H6��yO+Wz�q�h�PP���H=r�{@h�n�����mŬ�ܩ��/~����>�Ux0"o��_�c��Zn��E�G�e��`Q��!k����0�v�ֲ�z��"�j����lâ����4�|4"yOz���9�J�o�= V���(���R�.�K�sF�׶�Y��b�5�pҥ�KeZg��n:����!y�������!R���3]���;8��)�����>��,z�������}<�~ۜjU+enS�og��s-�:�k��B�� 'J�=�����Ofw�M�b�Ф�t�r���$�Ĥ[�hc��L��{j�(�?�^��G��������B���p��Z�p�9j�i�![�X�������ώj�w���a��w��$C|��[���e]A�y��!ʹ�Ǌ���+��ڊ6QĴ6����_E������.�^�K�"Eh����*h*��6�/l����������>6B�+�� ~Bh}<��(o��	��-����B��1��;�ިs����A����`A�`2>�k���>��|,
g?�t���_��D� ]m7&?̶���Ǣ�K�ҫ�HG�Xx���Oss�ؓ���e�3���97�xP���j܉��Af$M�T� ��T��yE������'����l�heLI硢w^H(#��6�R�5�+���n��+s�?B!V�^��Ղ�1���W��@B:�Gd�ʵ̙;�K��� ���/�[L�{�v)s�{��F�u�+�^L��J9ӓ�4�_]�xD���%g\��+�3,��1�}�J��Tϲ��j���<w]�YX��C4�.$���v���uE<�d���/Q��Mj�J�[���6C]Q5�5�����kd��K%>P�V�_����a������T@��M4(R���J����E�^�X��Vpɧd�\�fT҃��p��;
ߜ��ɷ��*J��ӎ�E�7ո������=W	E�NY�'��S�	';("�Up���<"C2<R��o q���9h�3�	3q��=0F�n�P�<��o��&��N���%��y�u����0E-�M�JXXrAa��l�ڱ끱�c�S��D�)Γ`�/�h1uc�jÕ�!�r�#3\�ڭ�)���k����y���Ŗ�;�V�-럭���?�`/EJ��'&HD�2��lA��p��O7!���S%��ЙJ�O�GqK��5ëa�7�U�z�ڲ��8?f7����4?��R`����K�Qm�	M��#j�e�_�V�Qib(�0��uV'�*��&� 曹�䭅��QF�}��҃}��89�#{6����zT���"qo���<o��>��#�IqM���sE>�'�yĪm�[��1�GS#QAD�Jp��d�Ƭ���J������_XK>����dMGf�`����(A�j%�*��#Ƣ���ilt��������b��zM^����%�YC�s����J��`�;���v2.���>�JsC��=Y�5� ��b�f@]e��Nc�}��y��N�
��ٯ�3&i��`[ �v9͎�"���n� ���@ȍM�8�oI�ʹ�8�x�+��Y���fđ�F[: #�g��@�)mҁ]��	��-��{y�lv�|qY�I�"���� ��jg�|�E)�vq������ɚ<m�hL�������f~�;Շ&�e��)�*�H�����,"��������ٛ�Ϛa�|�h��1�c�Po���@�7�6�w39�M��[��R��~A��$1��t�p������J�ir�d��"�A´�A	�!��6A���F�Ķ�hH��U0�>�wn�X%z��A[S��۩�R��G'ʴ.*˹�-�	W�jA�y�������U�/�������O���3!��7ۆb��� �"?b�x��Z���7Oj��?�<w�cO�qR��gƧ��"�D�;�<�=��s���Ȏ�DD��C�w{�~ vZ��y��b�K��멨�F�����3����3��"VR��([�Z�O�1�w�ք��a��09���Kc�<�=(�S��i���o_�Zf2��=�a�>!�U� sb��%9��_��L�Q)�������I+>lk�W��n�)�V�+\�̭hg8\Bz� B=��l�����Rk��/[f�L��G@v6��7���#�R�a���M�tNEW`���"�m���|ja�ג,C�*�v,�BD2���d	����f��͹/)*�=F\sTF7n�