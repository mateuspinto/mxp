`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7104)
`protect data_block
hhsISeZ/xvB6eTe7fKqSvGcwZAaSZb2XNuKmlHDfPqKbzjpeKDyBI9dEstcj8ktYKB8EGIkLjJLT
xo6QAbz3DFI9uhsUFq/IrfDgLKNHAVm2YrC9pb7azbXgnrClgJXlclASXSnClWEQnoKc3h7PjEL4
Jn6h6v/zRbnvRO9d7s6/dJFc4TQQj1wD1SaPbQk6ncDgW1+F5ypBtWH+aYtRhsCasqCd/b8R66sC
aRnQ8nKvWT00qHB7FN69d93346jIsGQsT4lrHlof0rnJmv+2awbzWOOvKbrF2CYNszOrqKfm+ITM
8LgpsiQxE78WADljGN1JJWr9GvIFhKEO2mOJE0n9ENrlcgmRylMtGSX0DslHsEtY3LysIhGVEx6t
53ajbLCQXSDqe7kbOzX7Npta4tul8d8CrnQGkoWIoZ+/ebLSxBykm/n/0Grbs7O5qLhVUgByEzkY
lcHdxcaGX994M6bbfN8SitU9RGOb1rccGhnXAJ2dwbh/xSEfH0NXZaCDjWj2crBae1nJNe1ortk/
lzHS4OM/TtECc6Nc9Bo8cTuhNT9AWNGdpCaO6OogNeVIF/jisVXuGrlAXp1FLCQcVQiRpmwi/jS0
vmcXKXunzmJlwW/z1AbXYwrmpLfILQwvx/Wjje1cYbJsBDcqKc/CLixvlYCG8Eyg2Z5RyZHpgEzf
YxPxZyFX1mlvQ226BlNGy/TI4ykLbOPrZqaoE9K8OWbpmDMCiBssJaF0O2pcpy97nlhwDLYw2EhO
Gaw1i7bC5opbA6l/PyZn9pAUeZbf1HDkO4cU+Gnc9wGrtVGaIoBchgjpi3OyrUcp1QaphlYkc/GV
KACaRZ5slA+7wZlLFG3bMTJwrFYFq/kxNoTU5CxAi7wmT+xdHH4vPV157tzdaNP8rgh3kHXtIOdC
FECNDeUU444yD5fDBY4sxhQMW3GOwaz7ch2+RYOQ8HBWcW88cC0oKsnB6dt5DiF6olt7TsDIsQV5
r4wAIDSXCTIu7rhojL0ny97T09hK/LiwF0XJshBrTUaL6riiA++6f/49uDKLQYZJCaA4PPzxsr6y
s5tUecZ5/Rtn4rfxND0wJ6dz5rkQ7JU0OniO2/fUnMV2M2W4EjaJ1/0I51S77jOrfPfB0T3sqxPH
LLImPHxgrTXD5W2F0jF9QlHzSKKfIPTZrTzHT/ntqqUi6lXkcehea+Yxjoowqf2JAnUdu7TRCQCg
qeih4NDYOkuQjwEJW3MozUqbK5z/CqJl5JZ/bq69U4NOJR5KhH9m6tfK9GALlL2ba+5GrOVw6ih8
TsA0Uy7fQnSZqka8JR5kScCQqFQ2bF9TVc4RaV+KkuBhb2fdpmRR5kOhco3kOKp4Y6dmw1f63ezb
ZKHH+5PmJwaKrl8PEVTiypqfgBFBo1NEihF6qWHprN5oHVPa+y3qIsy2OyEL7aaAm89WzvPJ0jzu
GpLk5UUcAb9qc4agCsbc0UpvV4b1WhQkVonSx6Od4+jcI6cyaGj/qOrZqL7V6s2rwM+J+1W5QMix
pPvKkzc+u3vNpFwzVHEaE7Dn6W668dAB7pkHZYARQhVvymtGKURR05ZK4iNJolWrhfjd/UmuyVKS
04x4hJgzYZ/MMQh0t4r8w2YkMFXbsh84q2ieBGvfK4tQpPYXxbsx6B8j5jvWyFg0EaI1A8nbcwVf
XBJbsHAS/MRATk80enu1UZ6Uwf8T1jIYwbqwPybqPZhry6Ot3FRWoD84f4GYhD80b8lr+/y66s+6
6S+ono+JHqz1uFOvt16JcyeCD7pEbkH5AsGA+BP8A6NVCpWIc6p0Mt7U08N/EBk4zM6wl5p3LY8n
z3RmORHnkaCnSHgNcAZywnspfBBdc4e8NQDwBhqrYPEJDYPvi2hpjvfvX9D8Ta25rnt/jPd6Jue/
6nnMBxsk+X2srUwv744WKGOBWltPkOSW9a3C/dGwKYmDGzLlfdmgWG0vhEIHZSXWDwmyjk+ewTUs
zQQaRLeBxVthtdySzfgOYm0Ntz3PqDIDC/CCg51qLlRr+6uXjVmbCJhplN6QBTeaqZt9hPCkXuMC
EVfnsEP594QEJoZU+Bfrr4Pu0P3Q44MT2oRpA2YFQdh0BzKyUdTtMF5+Ma4Is6k9WQMmEXN1yyw0
hMMI/Jl3LIBM4geQn6w2xy7UuaI00xlaBh//Ms4vfyMIspuDEDnqb5tjQOBUppsPUjZPGv/yFSph
5s5jtUzKGJiZkG84YUR8Lbb/4geEaDCMRVJofFElpPGMaOUij3d98OLImViualh5A7RCiRZeTSbP
p/+xosvXV2sFgAAvj3gBXKKk+/EW3FqWIsqNOOV388A2NyvI4sr6lfNH0f68EcsD+BPOaDtcEHE1
bxZwtIgS7BUILhEd8p8dTeTTgLs/iLsPbETyuNTkobJqEgweioauDWneOHiUODEHNpZEpMAuxVFX
jTWWvNi6hZ9Inh3uCbHYb/mkIf1In1/yE8TBZG7vfKbMeyAU/NXXS/RAKQMfaDshbmOZlTCfTNam
a/kbp0uWbemUt41JwYzn5+v2y++ZOZGBQuR9VZ2CA3dEpmEqIC2AmPLD2uQiJPG0hMWDYt1olecR
ENZotVNYE98Ro6uAuAt28JCzHL4GexBgkMhO8M3SPTWVm8/7k0tXA4h71d5db5r4cW0mYyZq+bSn
l86DpiOAqco1siXfZZD4B2egMrid69hLRUgw2atmpfxVm6K/MN2L59VZJoefirscZrSoCD+kkoPX
X0L9jvNkM8jLdiHpQW0EiJAREbbiPB8hN1JbdeKVAWZlhk4/khuma6zMo3aZHDiDJoAvk7XHOVyh
lSiY1xCY8SX8YmlRDdOqkQkcAFmhPktEmC3Nqb68Xg2hxy7TJATc2Gm+3tS3HclaWm6QwKAH6o/D
YbWrWl+AcpBQ+pHyhoAJop+/PmfVL8XxKsGsV9GsdarXHsFMy596Wom5DbAYtMq3u+hT3dhg89j2
huHwz9GwiuSjwec9/Ts5xENyZ9f+CKiAZY4BSAQoARNiAb5uX8EK3TyPVJfY7Iq2VwZmsjjNJBAR
B+t/IDBFgkjs3HXMck0KsBHVqjick20eQHnq8fNxKcEWWCI4ELCxrswIVhDGwiVaJrb7pjIDYF1h
ZAsosY0iLbE+b2XHC1za4CmfHfzMhfLCkF2uHovbAzoYkKk/jGgGMsFKSMsVxUNFcfBy1aQ+LNWh
MxwLQcenWFbczTptY+BZmALZKQTCrewAxsqtFyPtFzh4hDcE+JK9ryb7/UcMj2reb1Xk4zs9A7fz
HQ4YYocmjM+zzSLFqe/B1NVn59U26lLjOwhfu8ECPEpBRvOqXK5R5ilzUHYOUXN9PpnbdLB1D1FO
h0oDK4ZZZgn18mequb1OTe14MOxWrijr+DpSLaDK9Hp/w/fxBh6nXueBGQkBGQA06mzlLuQG5p+p
LJQNesaPV/Wjmuj7ZRhyWU5E5gW6ljW8C1cIwJma3koIkgXJqz+tE6yR8CZcsoXiXj3IN43uxPhd
RjjBdiwp0orbU1MnJPuyWcTBqvNZXCC0PYsi53HhYdOWxWwU7RM7gJq+LQjYnX7VhPJh2FOtgwKA
rHx6vjM//niwgbuHnNEX2bWjBMvRb+H3ix53dpFlpjDnKp93hiZeNz5NtkjLjvtLWMKI8Bw1IGPV
ZlSCPhVELX6jPBNXkTlV+/jaKf4rpz0x2925lO+2RKvjKXCFsbte7ZPKKW00ij1Y6Ls0HtbJs/a9
X7d1TyonP7U2Y8qxohuxa7ka9bGiDoijJlhrV4ITrgTaF/A+b0l04I7+U8vb9R+uJ07fjv5dzae4
9Bt3ICWevmxTT9pLlq1C9ZT/5TTeIVw/RTx2CPJU/bKPQDqZoz1w+37XRLCZOWG9WY9u78z47Wt/
m4wq+EJnfiTZyu5XTSKvD8SRG1jV3eyRKLeaS1LFwjvKIBqBqYAqCuS9b1DWirNqLe4E2nVI1/BV
YcNCQLPUaPzMFE00PQ8xa4//oeNi5dCpVHTZwMraBdkebRDMM++LBBwoZqcUumZpht53AC9zRW1P
rd2caLqoPi6XjtsYEsOobPi5S70S1/rSiCnUZAwSmOdKfpsyBiWUR38JFtTDkazLUL4258QRwtHW
1Fd8RDSppXN+KAHWM1mxWvFXq1jztBnuwjVGZpWxaCekvYqk7fkMjmtOCnCPwfwIQvwBX2XSRYjI
FCSnKFfVUpibtDMpTR0hRydo8wmRE9yzaAZVC2K5BZVbKkILn59F6RmDVYnx4mNOYAlCDN2NKYE2
GDhWO/LOQIo3LF3FdQwNV435hSEPMhyrLzvAMjqgP5xA7ehKBSiCTwCco2Q7v5ZLHJMaWUIrisI9
e68qir2HsyInni5KHxBKhRCjJ3RTmZnrNDV26WXbOkGbk6lY9XITZS/CIv1qbVTRNDq3HXU61p6w
FPcJRUl4drFHUHWyCXmXvsit7Wfhwh4pLOIimcl9dVOp1hFfUn/pKOZESR7ITwiMzeHcHwZiUasE
nfNCjIX8RG+k0Qae2uH825wH5LnmBX2YHH6o4L139hyu06ExcwfnaVSSz2WydarbDKsEdDg87Yon
fS3MlaWcZVNrfrYbnhigKOO3S6CjXOm1ojUhvNBwtMwTIsRscfsJiJqHKVp+Gbsma2n+o4/GP9RH
WhXWhpJSP6hrkPRGyyWy1YsQRS5m7Ft42rdtZEyx/47gOWmccpB6/wiv6EtutKoiRUP0WP0XQTqy
acz3mzB1YFBQw5SaGFggkCqWqIs97BViWG7n3RLaoHNnJI2cJIWBSndtapt1dRpnUUxz3oNnzILf
xwMUNsmoYENlvKZBdYcbnIGuQhQnPuCHTRJHRhLbK6e7vSAMRYjrRX7h2ndP4Gmh6kwVErWaanTH
jZIKHOXz3FAIWJBqjDqVDP0OdE7zZgB+o3bCAr0jC79wZCOnEX4VnuXgjT2uR1wQp4dFIjCVWHrA
dl+t86Un48B+eDsDV86gzoyqYmuxs1MeUpiCR92iF6NKLphCozAAliAuVfLymvZ1sYZ6l2NTiL6G
C9VOKZInewDdKuDy23SKnK5ry3iz544g1HVK8tT/iQCstjOojp3cPk7ha/mqyhXzysJ9JY/Xgrif
/O+zXPTUaEek/SlKxUdAqg4CUtuzs1ewxeVQoOETqbfkF8/GYgYzem8zkuBeLAP1WLQzrYOU1WDa
CB9ZNCQ5+sbZSnSEFpRg5MAevxr1ulvkV+7gaF0HYgzJ8AlUruAYMX3fC3s61W/OBJAXg/la9fNU
giZRL5/k+PV+NLWlcLj8KXBM0G12m3zX03QJLMAkQcBV50BjGYPXMhW50T1xkeawRqPrvrmgUe7N
UXVxa3QsUfJlxGGsOkBokNdKsb91UHnGPtV0xJ8k3GH9XUr3Z/EileXsp1sJbo1KAlAhxOaKy6Zc
tCJhdbStG94hNVJTZb7G3PLuSAuA2UL7S8eL29w3QBIyKFxUekU0CamWJrga79kZW5i1ASMQBW0b
gb7X2kBTX86BOcuGMRA5EtYiaBk3OHaH67JB68dMPrx21aDGeV+ucF7ek1VC9iowLme2JCqcVbgQ
2lGbAYXzabrg1l3mId3GM4v7+PwAwpZSQdk9ugaer77KKU+m+9uXFhFqHN/24lViWKc4nWDYGrfw
6/1UUf6TXsvCcEWQ3cV75Ti2AFF072XJ9f+UEqWqjZL2Xo12W0dsg+P4sV/SumFTc4rI3raVmwOF
qOWHbTX/MloiSl0X8Gl1rnk/NdOF9MkKhBKlDbdXr+YUyTqxPRr+Zhb2CbGuS2CRwy7YpI5yPJIf
Hhm/Hyl3O/LPiMcfqMpzH8rsIai6mJc+QNLxwsumwWqc84MTYNxUzfK+rVJT4kw7ur7HnzF8UCM5
khWi/3lLD5UMgh26VRecAy6Uw9daCxVbuWv4WAoZRsQ5Sa6KNxDY75zxdghKnVwy7O7ziiV/yAAa
eQAbUDbzIt12C0WPdP3FW+PGyetDczwhr0BtbCrq8QJoFrl8plJZmRjn1w4kQ1+X7QpEV6OhM6XX
4ssRPwNQ9WEVWaGVFvZn8T/iTGyWMlYgAsYpRk/uasPv+QTpGZtl421lWA0Vil/yxwVE7fkgd4mu
VZLqyIDVk7dPTjGm+m25zMlueahXnfFMh2v9E1vzDbRnMf72oIY8/aV5M9GWZWPO57qvKFusIU7u
uBbimwqIplECeReuKGutG4OX1RxkZxKaLC1rpdl5kACoDYliyLTHdZBQeRe+vT3xzpz2oE/+gtb2
sCkoTcbHX2LkqHxjMS9je1ITPyeKbS+k1MyC3vQgUHlRi3K8LkDQO1adtEpkVOJK9BbBN/LKI8XZ
l1G7bKa8QtIxFuiJBlA771fsUgNkj/IZNVI9h9AN4VQ1yHaPROpcLin4Mo/SqS/IQ6iZqxxc4DIz
KtgLdbQrWG7ZjA9ah89n1oz5HsTpIHvBa1vg4ImrbYFqknPapnkfzO753Bi8m0xyJhXXvFCFhhPw
QYU1Ef4pxsw1IQuqaAd62HNKgRaJNJsTW41poKXb24K7IKngilHlcgsJPiP1tBUtV7eYwazTfJ4W
ArlxBLMgPu7qimwVtGRaIRIHT9A8VR7fAvmqp1mf4f+J1sR7gtn8d4ekYSZmMk7xXBPQmIMw7PBf
WqEcTDJMFKu8mgcm+t8Y7nAOOEyhcDCS4YlflwWndFYQm72I+Pv7HCsFazV20WnYZmNES2DL6Ln5
55l/FE7HUc0bzo4j10Ssyt5ZTWlRblFkVGeK12jrsJwKvZADGRWOJh81geTmtpx8lbJ+ikJkpli/
pkQi5Kkw5bcZf73vZP0OGhNPZ/Ib+Dhgc1FPsDXKRTXgD3IoP7caJeDYiTCJoE/EbByCbjV9SHGS
ua25jIpHvtMzfMyKS2NyV8e9qsItvcjR/Tl1SPyVI7F6TfuynwtXGiJnjyH2N+ds3xI40tKhFVc1
jBjeXE0GGbUj4/+636sVWQqw1r9sQYV6K2YfwYUITZbTIdw1P1ZrwSUbBSSNRiNPY2l6gjaaj5EH
WDNf2xBNSSIAy+DHYJ+GFfrdL3viXZPwSEsuzgZzoW2v3yYWYBB277w/L6yl5By6ZwUg5Q2JGr6B
8B47bnXV0U3qdM+bln9y1SJLZ/y9bXzPfzoLW+igzKjZ6MKFVDCqNCwp1uTevAHwQ+bbwL2c3N+e
qBZCpNNOADJ6JfC2XaU8Gn7aHR+HCzHHFGqUYxdpM+f48m3i2BmyoWAwf9R7HFPMV722J1HDp3s8
4E58wwc0eg9uRksolHu6uPR6KmWugPnFIbl+y+rwRnKKrbLSpYT0AVVom5OlwFjH0ct885YtiKyl
I/GflZx1y0TfN/3gJ9I1qzLoB5rQCawWJuUayIrJLJnnUypXjJIZcs0YMfsQDhZCRfd7Y0kqQmmt
7hXJgoUEE/q7LXU86h5psdVJDGybkGKc4uJpJL93kpFSLRQ2trEJH4bSQrq9JA69OxtHhIEbN65h
6/8jsLQ+jzPaRrceTCqKk2sS2TcWZmc82HeoGMejetKBcWYDLM/tddCNp4TAW+3DAauViTNBhnXT
B6cEcRU6pnaEFiQgKZnqhPE1QEZBq1wEehcB+ymcqBG0tkAJQkqQoEmC/gDJ8QKEgalTr6LsJfaY
nuDfN47DrbuWu2IM894LQenxBuG8SkL01lyUiEBbZuDmJ587lqZ7fsm3kWk0tAqLg1fpQ5bwhA4D
F6VnQT5uZAfH04A7siRda14hoQIFLlH3MSSfDWvqo5qlIYN/0vITsZJMksP4o4nsG0CnFv7rdNeC
YBkLzRxXmNBQyMOM/jmcbZ02zyQbdMz3VKrMHmFFKL9G3foNccvoISDcG4lmUEIgXa7266eJqr+D
i3iRAaMSgnHJY7BxQy8QlhyViZHWdIJeh6S7JrgdETY0nNMCKh7bUW5fcL53lbghcRVsXyQ1jSYO
IUDDrzHe2xlrhoWyloYDtPEFP9ofcPcbxk8LZnvTM9wu8c2hr9iCk19B+HlVRTFTrVxUdRV0nBwU
JO0nc0dxgYT9oM7M0b9tbaCljzr4DvaPPmembVCbxg9r1P+s/S5dumyEV9d20i1NZ6lIWv8eOEVh
qhg37cc6LTJfHwG+Pnyb0Lfxj9QZiv0/v6uTAKEUpHj9o+T4Lt14XK3HALxZoWqIrWZY6qtfigI1
MLucdoQKRDNHqRVSDWz+q3GfNA0QL25ffvGRJ+lyMhdg9fbQotD4m6TzcGkvviDhdnq8LURPVYhl
feFKmE88zuh/ntNki01i3FneIrdjV6n/YRVkvy8TjHKtEG9UrhJpt1hzolfdlNpg8d6V+lnwyQdf
/uyZG7VvpUKDm+kGv/22XP8Mp3Ynqyo8mQPjmBAIwT5WZHZXp9phcbNCYDKESwS0+4tJ+u/3ccMX
3WS9u9Yt9MA7f3J1ZZoDuW/45h2qVJ54cXcgZ89ImcxH1rGygDY4pdnsK9jWAaviLGW2BjSgx21n
kLwCo8ksaKCzR9iXANl5CPSIF2lhagxHb4QFsaTYpZQT8wVJQh4DuRj+9Invz9xBYgJHliiqmynJ
b9mrcOS9Cvtq0zGhB3G/RdRkxCE5R3796NfCdXJRi7cWaudheS0MGyD3LjfhnLQa0nJuxjREb4Fn
ahd6gMtH7u37TSjiY0wc51vVJ0F+CLCBSimqzBAT6STi+SuPYFmmwN3vUxbqXGvgQQZJLQ/7g/Re
QG7UmiAG9Sh8eunZ6kJiJceaXBnsBXDV4TxTKHsf2hdULEb8z1N0CQu19V8n/fVIQ1ARuKKQq9c2
WoegaOX9woDsZhSxz/PLV0vWHQR70unZd5CXxzaCTFn9MT4BFX/3D8x8RKdZOL0SKr4b6tqmGK47
s3v/ZyDYPQuMYDPT4wBDFd8M2F71a8mFUmNO8SlIXcumGQ2cC5cBlWRBOGrF4DIlchT1ZSdoTbYM
qnj6E6uI4q0tfmZ6WPhTJN0NHXeinywRpYZecES7jtZPrbmwnaRim9t0C2JhQyFqDJTdvGVLjXXB
LaMOKdb7nglDbgZPpnIP/HFYYk8ELepnT4DKtwNlrL8ouVZqDVSEabl0Ckkb0Y0xvX0RHeFxiaTK
y+E7QYf/ThcICJsf4T7tATF7scayDWpDg/Wth0LzAxkfA1kLPfj5ustr21KnMTefeoNG0nQEx4t0
+UuEl/wAbztfvcp6pbqtCTpXwSZbt41Fl98RDcNKmtmrX1wyRIkF/kvEL4KPLLcXyxqBZx/7Wg78
sRVG417X0bnTyireMXykzHjLPnrZAOIDAweAzoQ9p8T1yOb+qZwASxslQ0PjvzWoJnQsIdzSSs2M
vpEt9LdQ2XQGax10TD/0rYMY2NryUTRWUF256n1j9r9iMSqDM+G8KJGF8Z1zIAmLpm5P9CPq3+VH
VgeoPAaULbge+SURYRlbTjkKFRgtfeCDoqWyW4wZpW2enAzrWWeyl7XoCqb1h+OuG13DeuY5GFCO
J0uH7C2su2LMq2cnpkrFUr3L2qjq/MKNiwOfmeyR1PxdyvRN
`protect end_protected
