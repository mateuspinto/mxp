`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 928)
`protect data_block
+Dt6IcmfA+XDe5A2ZLWBYKlNW1K7bx0+CUQdRVkHrZjGzWL9YYEaVFGGOE1w06UaseWK5UefK5Wh
ps3qso+bkVNR3mdJ1zkCpIqlzRwkZwCtM/NSUB7GYMkBBWFKbMQGd+odJt1QnF41u5P4Jn2KfisH
DhS4y5xB3rksZMssDhqgqI7R06NhGQh2aBbPjOk8QH3kOHmL2Wuf0VlnpJbPAvziUh3D6b//uOzg
31UkCfjOxqWnsrSKDBQCKUXfKPZbrJ/19Ufugq9OveN/13GjpsCR1rdIQiqtk1c6cJBSMpkrEOsj
+3wP5K672ZTqlN+FovqbC2xvAVl5Hm5yqtGua1GTiCICqA/OUvcpLIY61HFzI6KpqOzh/RJ7C7RZ
ytmLt9i1jfJ2y2Xgn1BXpHjGh4Ldf/tZlnEu2GYz36f9N6JWmOctss2MN8GYMao05k/CUIu7af3G
ULQaVF/V1gBGdxb5NAnRuxB+Mpdr8eCyCn8bHVqnlzdUQgUittBeAu2L1sJQM9tFn9T5DTF0KZiU
eo3zWhVkEdz1Bo5IOLgqj3jpMfQzPsv1jX1p6Wt3VkpQ3KYAZMPcmDwyKsnMx8/BeNTNjaeoU0m4
M5dRwvyQ9ZKc3mLObE43wcS0vI2YgmUSzRbpL49aepp8nTKC4r9GMKaKW/RJ4LLm0E+f1s8oOoVJ
6VdwHVAtbwJ28lmNSWFubq2luQKXzGDAKmTlGUdKkEz0hzpSb6osXpAM6KeXyH9sl7Hq6xq+/TfN
4GJ0zBabnA82VEuifIJLopKCRjv7Aaowo2hrKzD9tW3fUkavTdcr0Mm1PRclnQeN/FWyJzaEUzA0
8iW5Y2TwgGdSQclI9+/OR7WgCogp5tCmXLS/NLO9ZEibv5qk3py1eof+TMamXbTd/PQ5EFrdessc
XqSN+onkfhQQp0cY4VrOFi8JV7xKJsunNIOWO2I3b/dj5ZL9TE5840L0Y0ejpvZ2vyUHjmDcoScU
By/NwnnYmFruZMaCIiALZZiQ/l1if1fGD7o6D1mrJY7dR0XnmmIHyQEnj/bspIpYlvvrMOAvT7P8
0UHVLVTJ3wv7x0+JXG3/3idR4Ly2p6phTIQ8M328YLAzyRG21UyoZpKtqs7P0/ojicOY4y/b6s7f
+iSS4ipVITdqOoEDbqS1279/b0xldmwZSNUTV9s9p9RKqHOAX40IMr1tpIkUvf7oURFLcYgaVO7G
JP+ivq7oTt/+7dkiZwqAeg==
`protect end_protected
