XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��QR��#����5�)���R~��+��b~4�=[f<
c_>��t���Av��lR�_�-R�H��	y�����#�AS۩-up���^Y[b�µ�(�h�f��~{3�ߑ��1?X!}W3rJج붋����Z����S�ؗ�EP��<��_��䤟�"�l$eH�<���Ͱ��3m+�-�\����HMW��I�3�F�"��uuQ\����|�l�! S�zۏ��;j�����lV98,��=u�D��t�^o~NT8F����a�����B
� i�;ŷ�K�jd���%�6d��ŘP�tT���`"c�oXUt�n��$�o�1���Cb8�!���g�9aK�Gf R
��^�$<��S�|�O�
4��K>���R%�F\_]�F�$A���Gw�{��o�7���G	#���:R;v�>4iU�I�@��DPf����~�$?��>	��r����~K
���1�m�{��[��s���X�B�Q�����$�7�o!�㍾��+c����@�}�JK�S(��%��d�ڛa@k�Ȇ�����k� ���$�e�?E��>͓[��RT2p���d��A����9��G?�0��|մ����2�H͕�x� 
��'i����IO�� �3��p&�I	V3k�]>s	/���$��{(^3LP��Vhz��X,��%z�L��"T�_lJ��qd�o�_7��d
��w�ؒ��hZf1�A�ڗ>��T �8�:^�0|@������G��pXlxVHYEB     400     220+�1A�8�۾���ݪ��t+�s�7�
��aU�I?�W�#��Ib�t�JxԦSlv��ԧ,ݛr����q�XiC�V�~z,#	�S�f��#�K�)�dg�鱮u؎�
�j�?���`0!r�ɍ�I�ٟ�гZ6�|9�~�(fa�ju�S,Rq����� '%�  IX� ��~�7b���}t*�/m�}E1۞U�u�����H���~r2H����)<"�UL	ɉipHڭ�s2Ћ2	S��E�ufq�Y#���g���O���!�Ѩ��W5��aȞ����5�$:s`�2d��Vb�?�^V �ű�MVX"�h�Q�X��1d?Tq�[?c�[�_k2�Z��v�8�iv>��	�:�8!ix�/� �9�x�I�q�p�{�4��p��?W �dU@87���ehC֓ �_xd�&Қ�䆹�"=7#���5hE(H߱zR� ]##G��H[�hdz��ٺ���$K݊���*V����64R�e��{~���=�c����;-(8�.���XlxVHYEB     400      d0sK�$�٨�5XJ��\<�G��#����U��Ę2�t/�X"�-U�XZ�F0�6'
�c�Aw2{q��7饓����u{�C�'u}����ru&��x��#��)0C�� �c=�����{"(��$H���w؁��Z<3�8��c*}�̿�͓���(p��x(��}e>4.ڮ��񩒑̨K��f��pX��١I���;XlxVHYEB     400      c0 h�#i���߫�����.�=��44'T� �)�wYz���~���}a���Ӆ�t�DP..����!?Vr
�l�B|^0t(w��C��\��?�mՒ<:8@��_�2�D��H�Ѭ�|��P�S�%���tQ�h�9��S�fQ�.RŔ����L�$z����N��F�/!L�Qe���L��@�IU�|m���XlxVHYEB     400      c0�e@��
�zhuv��;0�$��K���n�y����z�`��q�XcWВL��s�l蟕�ԙ3�UqU��G5� ��Q����ıSٮU"���ղƺ!
!���6�F�`/��'���<���d��B���
R�n�һ�Ǔ*0u�p�4�u����RN���×��_�
Jv�?)�j��
�n�h��hXlxVHYEB     400      d0)5L�9Km���/�� �������}�	�@8�P�:���dԛ��-M�n�����[xr���U��DV�4XR��F�c�baVo}���,ً�+eo��v�E ����"6���uȨs�ߑ>k�.��#���g��*��U��[�����7���#y����I��D<�q�6E�"P��L^�.KڃYd�Qٵ�<D���:;�XlxVHYEB     400      d0�W�-�%G�>婁�ޑh�P�Ǯ��D�W�Q�CR�M��]�L�
�PBC���y���u/�'�[�����D�" l%����8�"l(��V3�w��&���82[!�&��S���X�`�g�lӛ�:�T���Oz�.��ݐ>,�D[PwCf��"��R�A#ž/'�C�,�-��Y�D�a�P6lz�&���5�rXlxVHYEB     400      d0j�7_E	�ϲM�z��y~Ks��	%�7'�A2B��8���p�'�����V���SBjb�m��H�C��G,Do�+�RLT�Q��ӄqftX[�fk�d y��I�O��v&��s0B�cٍ�CЖ.^u\p��!�(��������բ�mhX�!�|w$Zv4Rre��^5�t爥]���E����n	4��a�T76��XlxVHYEB     400     170l}B�6O�|�����i2� ʘ^J���L{a\����D�z�4�~ߧγ=��C\�>@���qE�n�%5D��l�JR)+��[U���p	��Ե�`M۩��/�#I�N\����ɬ�9��&jk�1�R��_�����8�;���L�Jv�b[X<�igy�}��~#��eDHo���-�����\��P���A+L�,�2&�(�ڍ\9���s�^T5��[��Z�s����		#��v�Z��X��lM�}y��=��S���8H�z�ǝP
�����HX{�?�����)�dbu7��O~Y��,OFF�3�į�)�CWܻ����e-���	ukG��׿����e���+vSXlxVHYEB     400     140������������;���]�ՎO�_f+7-eo��*�6���e�]t>_PX�C}�JEn��E����U0}'��pa����I��n.|\V�:��20*����ᥱ�KRCm�vf�8� �n�����t}�.���ȐS�#��z\��D��R�ɗ0-X��X^����lG�����2b��j�}`T�Qpmt~
9	�	�
^�ر�D�)�}�q�}0��&$�;�$U�S$R�"�7㺔6z:��HKՑe���M�7�u#c3z���7��J,HWH����f����ۉp�e����ofϱL	V�2���XlxVHYEB     400      f0]�Z���z����x�%$���
򉞤i㢆j�B�M*�~W6 Jb��R{_�6r����Ĭ���Fc��!<-�CZ�����8T���E`��.�a��$ώ�1烤��Z89��v�t��!D%��K���#�8���r���#�0L���1�VV�?�Xz��B�e'X;y'$�x��T��1 KV���6i
Á�)�^W4M꽼"����?�z�<�V0̮�J�C��T�16XlxVHYEB     400     100��&D��e5�������w�v7�����FWZ�/�	����D�y�1C��\�?(�&���ۗzX�)��A�0���.��� @��=͠En�׌��x�}���V��2��­'�}�v�����ɖ�kn���*o����%�'��g����*�%���M#��P*eԬ@�� 5D�L�1E�(��.��D�p�2	x��+D��k�+ɞX0�{- 7�������
�`<3��1"�!)U}�����XlxVHYEB     400     110~�T�"��u�9B�T��Y
y0�����Q]��_�D?���z�p�9�{#4|p>�J#  (��-[���$�#g
�߳��=g �}�,$���6�+&=�;�z8V�f�y�LY��ʭ*3d�C��ܒ�.@�+"�k�F��.�m���c�����30�ɹ��c���y����x��?���g�դ|�������$�z��GTb���8�NE�@��i�(�#��9}�
��8G�J^ؽ�R�;2�P%�#�w׻�֗�%�ZWG����3`�N����XlxVHYEB     400     110���K��3J���N��P��І7ErE��L%L��#Y�lC�P0-@��N�sf%!��c��X�	���1�5Sl﹤��@�����L�D��5����q�!�1kH�O^��E���Ot��c�ɗ�H�8�¼d4L �ԍ�H�ۋ�H34��V�ŷ����~�J6[���>�[Y�v7̙n��<.��A@zd�R_�����A�3�������'T��FN3�E��pr6S��d��X=a��_?ݤl�3�����l���G�#�`ɚe�XlxVHYEB     400     130��W�:Ñ�-U�t����m�5�Q�OZ����Ӕ[��H�����2�z��:z#�������aW;{��gg��_��a�|%t�#W��A0w������w�M�|sO{1H9�?��$�~��l��i�:���X���uz @id�\�t���X�jbS�P���6ڐ鸶��ޯ;�a듥O��g>��I'O��t�ӡ���I�8|���9;Ć����<��+����p�:Zy�3mEO�=�z��X�08-�H�4;�f�Ęu��Tr��RU���w��0�2��Y�u%�&~��~XlxVHYEB     400     100j�K'Q�p#�,���{��3�b�Y@SѰ�)!�K9�<
���?���ˆVȁ�v�켎�L�;��ETA���O�����_�_3��1�uOUY<���?�=o|��2*u���X��:I5�wx��\[���ը`ɋ;�ǮX��ҟ#mp�S��#�7�_vSK�I�71?��Q>';$
2㦈!s����`��	�I��Ā?=�I�n���@��I�%�ux�+*Fc���r�=���Y�OJ`�]�4ZXlxVHYEB     400     100��F!�#j1	����Q0��r�U��6b��m�g*l�D��~')�xb� !�S���H�o�S�ȷP�wG�B'�Ri�sڭ��
��Ăx!�J�*����=��_�wpgQ@Y����y��v���K h�,�t:��Ske��󖏋6�䥀��Tk�.�p����O���oی��o�p�"|b�&{#���(�+�)�Q�?�����ck61>݋X�Zs?@�rS�C�C�}ΏA&�I.�%�X�XlxVHYEB     400     100+2[�q�@Q3�'����V����R����\��$��?Ka�Y�{�l���!q�]���o&�"D�Є�;[e;9ع��6U����5B��-5��������_qB�q [yxH*p�3�C��Z����}��yM"�����?��?@ꯃ���bZ�߂.��/�J���,X���Jn��,ёB�d�u���nH�q����W�r}p�g�{Za�&D�������� m�%1)y��1K^6�dR��XlxVHYEB     400     100�ʗdA.�}1���YH)�m%�G��tӯ�X@̈́<�{.Ș������ݲ��2��㼵��?Y���K���BW���a�w�QG��uL�dU|�Ћ!l�d�%�3*_�������1�� �M�Y�\j�{��$���|2K[�?�ު��ЏG�c+��o��"���J�������e�9'�dWPbɒd�G���!�y0�K[,�
�C>�$��
�	���w@U⒴ޱ�#˻il�դٻ�?iJXlxVHYEB     400     100��M�̰��v����N4��1ٴ��g�(ܟ����kh�p�:ܰ�ң��a�(=E|��A��;3��#�5�(L�r��G����fluAe������N��n�A?���kR6�ms�S�_{���֕]�~�T��ZNgg��<����Eˋ�Rj��:#)ɜ��F�Q�t��$�I�H�dp=���iR��2@�o.F��H�Y�5��7�p	�]������g�J;d�	�ץ!s�{��q�JBMt'�n1A\j?XlxVHYEB     400     100jّ�l��qC��g�����8�҅�O^Du��l��o�����O3��SYy>���X 9#{5ԝ��Q0�c���Eoo�=
�WY+�j�*��6��D�|v�uΉ>��n�=�����C��+��=����U�a�mB��_)��>(ʲ�S���
ۃE��%(�d�,!�%΍��ٟ�85��� ���q��>��� ���m���J8��S�NN��ω��=�GC�9�A�c�{�â�3�F��o�XlxVHYEB     400     100�,"*�RAn<��r���m�@I�Xlf�)M��!/���.��L�W��s}	_�X�0Xf��3�'��EZ�0g��ű0����D���Üv��~��:�K��Q���iwu�3��Yt�Sc� z���Ɩ7U���\��S�r�~��������j;�l�L�7Zv)�y��e{�h�ۤ�4.��T�י"Ɓ�����%%=�ϡx�Z�����O��5�W-�t�Z�%/{�K���̉/� �O��i��g���XlxVHYEB     400     100$o�:��{���bJa8kS��ya�
A��ڳrgn�q�YD��?�/��&�����p��`�z��
������}ͱ�{��P�RU���A�r0b�d1��3@��4^]�Re3�/A�q���Gi�L�~p�vg�&,�JƋ'TB3��3V���@�������9[�@f�Ӗ��,ce��m���|ũ6�������7`�=�a8�Gň*"����C-�%�l�\cu�F�I$��@�[�F�.M���(��BXlxVHYEB     400     100F5y@]�� ���V��t���%F4���c맷$["�k�}<5J�՛Z��f^%J�4��|M;��6�v�����w��:ߡ'�y��h����ce����9��~��X�>ĹI�
�2k������l]D�z����,o�����i����3"􇥜߭��lkS�� �8ca�Uaל,����O5�N��_/aя�V��w��$i=��._.��'��T=����U?F%U�tJ�C��Y/�2�j���B��!�XlxVHYEB     400     100������쏙��N�׆�oa�Y-��P$^���g9i�PЍr3n���},��J�;si��a?�3��=ˈ�M� d��ƚ8R47s�
���\��%����ђ�5�����t42|#�':r�r�������!�V9ǻ2oG��9	.����M��o�X3����r���l��A�G�q#�"w �D����qQ�,�5�w������V�����`��U�wi� �>���0"">C�bŨ�v����3d�!vB2XlxVHYEB     400     100�ȵ�����D �-�*Ml�`�<��c�0�sM�7s�F�� ����8���h*j��⹈���K�Q;/��Z��ap�X�[97��-�u�s��%�$��R �J��)��J0�w���(�f�(pf��$p@(&�z��%(7E��a��*9��Ҧ�4xT����14q�H�1d�o@~Q$�\�޼'�C��& ����ņ4	9�|�5]���@��J��Ŭ�Ld���W���!AR�g��|.�p�V+��C�jXlxVHYEB     400     100ݑ�����ي�5��M�r�?2k��s� ��<�����ߜ���1?Ib"�s\$�E_�3�Š���$N�3�h�U�ā~�	��$a gv|D�%������PV�n�u���B������[淎+G!'��cZ	�r-˩@9���"�;�w����N.�%j���g$��g��
wَ��!�TTP�����zT_���Vi�}�`EO��Q�Tw�� ��kG�I�A����g��7��%ϯ:\�zj9�|����.��XlxVHYEB     400     100=Q�m�@��!RiHz��p�#4D�2�H����y�Y��0,gT ������__�
�·����H��T�̦�,����K�.�t�������ͅ�����B��d�յ�J���`�l��һ�
�Z.��(��J̆�w,�79�>��~k�2F����%GW�Pg^EFk�5���K��ͭ��b	N]�v$zN���� ��f(r�&��A����켜������`���r��� XlxVHYEB     400     100��:z����b@bV��#Զ��aR3�뺺a��Dp��f�b�(�_��b�~+<���a���@`��F\9Y �)+����2C�ȁ�a#��6p���ɦ�.���Jد�t��#B�� �F�lC5i;0=m<�
]���-#�OR���Wm15����٥���_dF�~�"�^V�G3�ي��_W��P�P<�V0.DL'��]П�*�;*V#�R&��#S~2?��BlT헆�ʇI�1�wtXA2)8�^_߼XlxVHYEB     400     100>��+�t#0��� u`U�����߫�n��2K������~9���r��bw��%]�N�-���>��u3Z�"̄�������Ş��L�ȧ���~S��ױ,�(w�Jܞ8G4NSd�V�ܭ^r.���q;�EfKvi+R����"����9D;d�UF~Hq��ܭ(/x�d�it���̀�#vm �D��G���괱��p	(<�x���:��?��of��E�t�v����`�@�x�����~XlxVHYEB     400     170�et�C�a\�o~��U_�-D�ݛs�Y�Or??��&	G�P��4'j1�ʞ��D��1��x>D�H�j�\䳗�H��9�ДV��o�
jPҕ����t>�w7K�������K�&������95E�;�`z�Ǚ7�1�����Ĉ[��X�ӍC#�e'8+�a�SWn_;-s w:�!P�gDL�>�����_g��m �k.JU����&��z��J�#�8VcM���\�J���$gS�93�ù�?�_��%���P����U��[�
��M�:��S����H��_/	�(�O�)��_!�����M��#����ҶQ�U`B��{4噞uj1!�Vڎ��I/M��P�2f5lg߬&S]�U0; XlxVHYEB     400     100�Jf۾O�0Yc欑F����Y�C"j��C�-P!��@rU�^���ǂ1H	�<���[�D_��� _7����СJ1L�D������O�ؼ�-�öp�X��f˽�OݵЎI�U��� ��T����G�]��A��(� �h�c1@ r�Q����C̥���5L�-�a-_bDUYѓ3�6B�
g=	�p��Nor�"]O�0Rl�6܁���0fɐ/R��V2Ea|�daPf5�S����}U,w�)���~(��`��MXlxVHYEB     400      c0Ҥ��d��|�<�y��H��x�;�������<�Jԟ _�e�,=�M���;���Y��R�M8�8�t���l�mg�*�1��ĸWԱ�8
-	����2W�/l�?}�a Yϓ����1��`��5`�:5,�i�LڄNPT����Ǯ��ֈ�7p��%Ф���i'���F{+���_}��n��9�	�IXlxVHYEB     400      b0Se)�P��f��È�=����f���JW��kN�r���b���h[����� �V�i�����sNy�X�D��w�2��nR��5ݰ�N��x	������~^�y�6x#���	�m���8�k}��ORt�517R�ܫ�z�JE���k@+C_�JT&���������b
����XlxVHYEB     400      90��	槖j�*D��{�2E�)�j��K�>x�ڏ�'a�u�&8�׶�[�j�t/Z�bg���ԧF��Q�E~W�p��q
��0��.iQ�l���-G֨@2'�(Km�:�] ��̅q��J�Qw��*�%g:N;!��o��9GXlxVHYEB     400      90�/�fd\�f��sƟ��Naw�Q9fRvjLpH5� ���z�נ6 �)�t����M���c$7��H���^R��s��� W��L�!�]��܌��r��3���K������E��P>E�i[h�2)�R��\��'wf�єS�֙�=XlxVHYEB     400      90X`��Vf�~��+{E��`�G��"/�c���U߀~L,������BX�/X�5TYz�%��g]y��A��$ܾ���]�����_�]���7���K�>gWKN����e{у>pЗfZG]/�Џ+,���Du��A@�u+g�DvXlxVHYEB     400      90����e}�'*�� GO�$3�3���i��.��
L�!F}��k}%��ƃ*�A���c (�O55�@�Ia��L�	$�� �}��U�ǧU���T���η�bQ�����!X$�B)3|�wԹ*[���F`��◶��-�>�<�XlxVHYEB     400      90�����Ȋ���������Y��Z���r"Se=-�Ek4&����	6�$[���8_�p�8���tZ8��S�	������U�G4Ģ��R���s�g�&�7n3D���8��]�[�a1���-�7��������\-TXXlxVHYEB     400      d0� �{{F��=�R��*���&�8�[+
��L�q㫇��h`�K����S�����JX�`���y��X�n����I��S�Q�x�pf�΂p9ZCE)<��c:<�6�Jn�K�aDq��Z���PI�F�"O��h�P,G��l�(
��_Nk��P�[S�"6��#���)�P;���>�����v�xw����J��	FP�XlxVHYEB     400      e0�JF�$\#�N0���r=LQ{�2W�
`ݓ<����AYH��Oe*ޛc	�ؽ���n^��xJ�u��F�]U�%e����9�GBE��B�����75�R3�w�56��������R��������|5����Dc!��4�`"֌Tg��B����iӑ�H�5��_�-! 1��x0U	��SkT�9ބ�;�g�k^9]R�|p�u)�i����2�q�XlxVHYEB     400     100.��1m��wzF�k�Ѽ#����#/Ÿ�ĳɉ�Q�/�h%����
[t]�Үڂ��"��u��P\(9�K�C�dn���<�JO��T�g�u�gţq�O��4�˔�ϛ��	/1�CBn�o5h����H��73:^?׎P���)Jq3"�!�}}4E�����q��aN<nH�/�3=���<�����U�2
"�J�3�`&Z�R���P�d��W1<}���!�^��1���VS���(�4G�`�)����K�TI�^6�XlxVHYEB     400     160�W9�u)P	�\���{�o:*���G_zd�[����~���4�Ҕ�$�㐑 E�8�������������lSH�ZD��a oى�uI��#�oOH��'�d\&�S����|D�� �������o�;���nVD$*�E��\~o�qs��W�ʳ#�v$En�a���� JFᗁz��[q�)��P�2np�F���!���1���L�#괭���g �%��@&v�Rp��:�b�ȃ�ҁ��4J�o���
 �gT�n���=���X���A�
k7"֗�,�N��=�]D�M+DXh�!s���#��Dl����|�E_҅���%���,/03��� ,P(XlxVHYEB     400     160�4�k(��G_?J�˦)����>�V�/��ɰ�M �^��_��A�|�|���+�|3ါ��Z��l�ĮL@
o�y3S
:�"m]�uG�A+��lX'Tbt�6��M8��Q�����y�	����W]`E�o'O�mNҰ�"W�����M{�����(���:��As�,�O������
�{�N�Q�6e/} ����5�h.k�G�)�?+X��_�����U�73�W�� ��>aR�\��"r��;�5ѢLѕ3�L��9�d�t��Ӭ���nfh5���[]�;Sr��l*�L�B>F�ǆX�b�c�M���}��*��9Xs�����۱���.�����SX�����|��XlxVHYEB     400     140uܔ�\�!2K`���T72SPbLIh�U��\vM����f�pc��L���S��m͆���`l��v��1a��(�u�w�Ǉ�GQL�#^���
D��vgF^�y�֊���b^7��x`Q�GQ4Ar���8�M�����H�"�7��0sx��JC\���ފ�q�R������Sk��t�"O�'��]����sO�u��p�r�Y(�|��8�Kl��ʈ�E�'���ޟ,w����W��J�ƀ��nwV]���A؋0��E5��^�ig-Q,����q`9
���A!�i�9����c&I��K/lA���u��c�����XlxVHYEB     400     170^U�1,���qh_m�~^F�J��.H݅|
����&MO�ǵ��^e:"'TV<v��-��Mo����cǲ����3J@K�!���+�s�7�l#}���ÊDu�L�>Q,B5��q�9�9�x<��"��0��2ZC����,i�V�g�廌&���{("�/�%���D4_g�%{k|�Y�s;��/�T�4�5=��/�S�8�� �c���C��_��ԗKö�z��C��ޥ|�͵ 2\ .`n(F/�:ty�q&�j
/�D߼ڮ��dE ���WNӢ1��I]yW�gxa��K��׊���q��o��n:��J��R�����@N"$�e�2g,��!{��։?ێ`�9L��6O�_6g_�bH��������=XlxVHYEB     400     150 6��B�!_�1Xϧ��ّl�-sK��î�_�h�p�8j<���օ�f�'��A72�x���.�:H��2��o@��i0=���|�<��M��D9oNu��i�j�D�@���(�$�1���0�
(,�UW=h���6�;a�itz�9<�������V�� ��Y��%S>�ŎoN���V�;�%_�sMt�r��4�mw��c��x��T]���})M]qe&6���x"�yX�@��X�=FEaO�'Ev����E �́�HB������5��ߒ������ �*cqmd�*�Ny͓g7I㩮�Z�U靥X����h��	�%�Z���ۀh@XlxVHYEB     400     190�qkW��9
���{*Cޞ$����U�_|�~�p�Փ���h5R�2��ž�hk׈;���l�Vw�"j@Z/Z(��v=���Gsv.{4�*fK`dUob�C�;�!��@�m��!-��Ě���Q5R��`���<_���ZoA����1���,\�G~;�Q�$?A�5N:,���s�b�ԧ'��Ѧ4�-�zn6�/vyb
7��:�`���vӄ1	z���cB>��!5߲S%���)r���&]�<���K��;-����2����&��D\)�T>�aJ��D���
���� wuN�<��U;��w7H�t��@�ʩsv�-��7�NF[���B����犴,�f�w���DB�1w��o�ғM�Ϧܞ�|�$
).��$�b��	��@�;r��@iXlxVHYEB     400     150�L<�����Y��O�[�q臚c1�&!��_is�G���o6*:xD�AHʤU�o@�6���P�V�	�}�9����Z��~��+I����O!�Unѩ��QҬ�H�iv���Л��̽B�q6�Yk��/�ArP9��Ȕ��j��]���~՘��ve(���,�U��
g�	8Ayy����"S�	W-�N|<�9:��A^�>g��"+�.�Ŋ�$_`��/d��;�̩�o5���*���������3���Oa,�UT$��ÿ� L@���n��h	����H"�s����b�iO���y8�LlN�`ϰv1ݠ�q'�9O}��w������XlxVHYEB     400     100�V�+ܛ�k�Gi�2 P�29nU��p��%(�b4�6҃�Y�;�yi����i�����J���o`N �Nr`�I!�R(dT-�#�ӗ�x���,?j'�"�q&�����ޥ/�m�ߤɍ�`�8q�[)C9�Jx�G(j�Wɔ4���qdW�I�ju���y�y��,5�(��*��ݪ@Q���B��O��~�Nq{0#
��ȈB�c_m!����������<��{�u!P{t�[�5aXlxVHYEB     400     190��F�SWҭL�5�]��
$sy��}�h~x�����;͊m�\��x�N{��1���	��B!�����g�*���w�f% *l�Y��?�����#�l0�_���"TYȬ$�P�N�7��e��>�d� p'�5�!�l����B�Ц�-R2�Z���@��_�i��;2:�%�)/��ӡa�D�#��$��"uY��0���ܬcv�lTׄ���҉ʪ�ket�����#]E�oDֳ��g�(uupP�޼�RQ�_���y*j��w�����)��q�ꝟ�%麟�i�V����K^�\@�?�#$�l����+�4��ǉ�_���$D�,���{�i�r�����]��u��9����c�*��s�2i��M��T����{ro{|	O��RM��FXlxVHYEB     400     140�#F�����Yz7��`�?�Vy����94y���M��Mڗ0ǛS��kAu�I�ףixՂ>A���,�(A%��_��8�EY۴�Vڒ2�������������w��� �z��T�P'Z7��G�&���g/�b�E�q�I��B$���s��B�>���|<F�=/�;����v{�A,2�Ҷ}ζ�[+�%V�����0��[eɚ69�:3߱Aמ4[Rt�zȝ�G����P����)�q���TJb�Q˭e�
���r,�2�F�jo�]ݵ����e�7ײ��)������A�r3��T�f�XlxVHYEB     400     150z��X[ ��x����Dh��렓~�"��=Ro��twd����M���}���F�0��#��������n���o�脹����o����%	.��t�i��u�@w���
z���3.jd�y�E�]z�����/^���DV�/
�X�r��=��uOϙ�n��Ӳ�����w�!��m*O窝bFۨ1�`�V��*)3~.�<�Qs���-���t�%�6���e�)�����	h�V��j<,�`%	��q��i��L$!�[8(��~%&'r&Bc�NXG�sB��gg�O�T"E��>����M�Ϟ�ӣ{H�ܢm��XlxVHYEB     400     110��dp
A(`�n�E�{�EX�d�u<�&7�4rm y�6p���~y��8QaB��2�@b����YF��� Q��]G��c=����=�p��b����QV^�c�VH��B�^6˰X�!^'��<��w�jkf��2�'�S��]ܻ fG,�jX���9�~��k�9)��F۴�Tӛ0�\1��N��� ���j��zҭ��m�h ��Z���n
�eV�@�p�A�z��"�-%!j��G�1�7?�!t��������,�5Q���l�XlxVHYEB     400     160�n���Šr�M�Z�T�5	C�>�D�����1����.��e���;��:qЖ�c�#�"T�y����\N-W��@Pv]���F �I�Ee�'�h2No
j`ס6,I�n'��ޔ��\?�Yڣ���Ȫ_���3���S�ˠYh�0/���#�K1(��9�����~	��'�_�阠�Mt���łJ���h��|O����B��<������|i��i����4��_��y��Et\����	��_��Ifz��:W%=_�H4�xȁ�@��l��9s�GXuN��j�#*���&ߦ@���;��qײH1 ���x\����=Z�uNPF4Z
�L�]z���z����1i%���XlxVHYEB     400     160�!�Ǹ�C����Ɍ��@)���c<Z\v��V��C�J�����������e��?ws3,��9�B�N��'.���L6ӂ^@f�>'�m����i�,�2��qՉ�s���k+c �{C#���N3�h���$�qΎ!Pn�tH�3�.�e��t������$Iǃ�#K��ԝO�����+
i���˸Z�� ]yy�I2�?�{L̯��N4ܯ�����bi������扖g����y�brn��f�k�Ჰ�����@�sŮM����;��c������v�x�ǽ�Zs�b.�/_��8�w�$���D�����2���v�dߥ�-X���XlxVHYEB     400     150�ۋ�#��;����t���U@�F��Y�Ǵ��@�>g"uR�6�eC(ޭ�wzmU��s�8c�2�pδ�2�.#�MɅEg
��
���������_�`���9��8n��SFlݠ��>������p6&�����Y��t#��3`Te��]õ!��Z`��`�\�7W ������1u.m�Ll�+��~	����t۶s��ĩ��� �籵���C*Ƿ�;.�/�>?�ɻ�/��i�|W���"��BK��l���ߵE��G|~�q>����a��m#��6'���ա_H�2��%�+-r����L�d1�	�������pHXlxVHYEB     400     150MK�UU³7�c�� =C�Y�M��PV*U3����8`���j`��%O���ˀ��*�@:6���ǟ��#�=z\�l�C���z�)4�ͯ�,ő*s�n�#Y8���?�bygc%��R� P +c��B_��~Jvl����>?����d���>���9�r*ϝgcrL]����� z�K��E�z��m�ílA���w����M�q�j
�mZ#���{�Ұ{(�ϟ!�q���n���<��L�R!'ʋ������r���������G��X�(:�rI��AL��ƴ��(�u���w9>�`����)êL�)�8�XlxVHYEB     400      d0�����:e��z�%E�QSi��!�OC�'%T��"G��7D��7�7�Q���[��Z�:�<7�`�g�ҧr�{�}��f�aX�0	��)(i?������/�7xBa�Dq�.�
���z��\8SR�>bD^�o=z��*��^n4BڜC�Z��~T��
.�S���ը�d`����W�,Z&�������ȩ���򷦒/�k� Z2mc�XlxVHYEB     400      c0%�Me��;S��"�
�S�6bm�
AO���L�[C|~�ӱ�y.�R�M��ɖ�
���W/TE ��Z���)� _�2i����B9�~#�{n��F|�V���~�3"���L��±�j~2���7b�b��n�4�x���;�%����Zl�q����Ee��W:W͒�HY)���8%�n�?O��XlxVHYEB     400      c0CYT��	\��f�O���qg�g%2*�P��@���%��t���^d�Z�� e�z�d��t�8��ݫ�T�]��b����h���q��������p[ÃE��8�/G/�:�I�%�D�`=�J�	�Ԉκ-~إ��9a�p&�s�PA��R�	��hGYR�3���_
53�%��ְf�l��bӍ�XlxVHYEB     400      c0���.Ư�:�_����/���L�����h^
҂��t����a�[��XA������1�^s��A.�"o�"zp83̎���-}��w���nr��a��ᵶ5)�����ṙzt�C��5ҋc����mK�ggT'O�)*[����$��R�;ӥJ����A�Hj�v�*�eY2?O�����#�XlxVHYEB     400     100q��o���a�����SFed,�;�U8�<���?��W��7�����r8<�n;�m��tiL�ԮEd�����ս�F'tE�֏�;��!�������<[�/%��'ȼQW�������3:�$N'Vgwʶ7W�ޠ�ۡNe�	ևY���;%oQ·U�w`J��!!7d�c�@�Pۦ53�j+�<��k%���QdW��̂a���U�Q�����B�,/ƞ;�1����,�����r�{��L)GxUF��N�*�XlxVHYEB     400      f0)]F�zd��gكi�k1Ǩ��6�XC�imacc���&����ƀ�2DM-uJ:��V��K.��(��[��5r
n�C�E<he��ioC��Z�W�1��rj%VE���]�˂8���s���D�U_�M;X1B�J�!
��u�u�j�V@pkq��糹���2H��bPq��+��#�<��/�n�ett~]Kŧ��Z��j�R�c��2�5p�D8�f/����̀�ɟ]XlxVHYEB     400      f0c��໥�g�����k=�Vڐ���N�lE(e���Ь�������M`�Ԧ5Ͽ���T������ۥ��Y3��^��zI�&�����dx�-p:q_��̮T,��RMp\0Ɲ�C�-JO��V�(�3�·�����{���گJ��ڿ�+�z��k���yFʲc0�:Q7G�T�W�c���B�m�C��0#u��V0On0��ڛ�j��j����ş���2q�XlxVHYEB     400      f0-�C�]�,2� \�V,�����#���\����=��B	�<��z���YL�D��"lȅ��Ǎ��Ũ��e���$�cЀ'9C̗���&�K�����Wl�t������#�}}�$�E�y0a��J�3�ߟ �}�H��8.�b�N��RF;0$�C�q�z��͂c.(�y���4!�<����m6�Hr��"�����0�SL��Qwj��ڲ񏝟��g�A hSL�,���&�h�mI�"XlxVHYEB     400      f0^����r���,�y�=I�-૟� 7�Xm1�q�v�L�܂cz˸JJ�"�A�,"�����Z�1DߨW�J�����S����2�c,uYF����>竑n������O�CV���J�FM�[��9p��4����=s�cX9jDi�+��`w��R�`p�&� լ�m��a3C�K���A��U�A����X������}�X���p%�-�&��@Gs{�0$JE��=�T�XlxVHYEB     400      f0��*���˙ި��T�xgs�����HР�0E�&�0�H��P��@Ҧn�
��!]���qw� d\��C�M<�ۓ�`�R8xIr�dF�*`FgU�ɏmڮE��u<r�8�K���1���Ъ��f�>�IT$j|_����?"��v/�M��k;�7�����d$�N��Tb���/XIϔ�f�{�w�:5�X��*L>PN��Yv9����K�Vs����pޕ�>5ԃ�' �_�,�XlxVHYEB     400      e0���D�r�a!�Ϟn3*���r��]����`���^�P��֌e݉[�E�l���LX�-L�7�@(��\���ܑ��j��eҲ���r�hȇp�p-n9����lb楷=��c�ɯ��I�S=c*&d�\��䦾�N���H��=������!����2Y���ЌH��E̘��v�M��� �^DY�;�d�LF~[!�=/���8��9@k�,XlxVHYEB     400      f0btޥc�Yf&��j�:p�c}:�����e�զ���u�¶����G��H�
+Pn�#�K�s��
�V�&n����=��{�T��hM�k��o)�u�Oa�} �(2z�5]V�d���c��� �Q�񙫑&�5��UK��5����]��4Q�% HC��cXz� �'\uHJL��	6y2�e ��4��,E!0/�O]V2�6B�zۑ3�cG��T�/*%�R������8�5L�^�\��XlxVHYEB     400     150+G��tD�Nt�X�4���֐���H| �?��ݓ n	�S)Q��Xo!�Ԑ�<�F-�]�����X���r�w[o4C������ªϬ7XJTXOь��X�[���u (�j�̒{��&_�y~�G���PL��쟾B�����ŞG�0O�+<~g���8���`i�9�턬����"v�52��ȳ6~a�)'TF���Ds�58���S*�K?��vUD���z�#8ٱڗ�{���g����<0o�u���<]�����?����g��TxT�푥���8��_�.r?��.,�@�����j�G]�	c�@�P���o�Hk�R��n��R|0XlxVHYEB     400     1a0X�IkJ��TS���=��~�l�c�.$��ǙJ��p_b�Yh��/~|36$��K�d�af/�̅�8!�"�xǘ]��!�hp��o�~�.�	���Er=��^�9F�M�C�)?]��B}@��C�`���^�tX�^
�#H'�=�E���$�So����_Kߟ�@JYr�S������U@~ZE�_��}���	���I/�]IT���
M5G�s�ys�6�Ƨ���3�!�`h!*������0�#�K����0�j����'�}��$~�F��-f|3lT3 8N&ݨY�_�O�;���Q=E�3�%�����	$#��,�x��N}?-���N�e���؇������L�{�g�~��o�d�񐎨,�<�$�q-@�����D��Z�L ���G�C5��류xl�T�*XlxVHYEB     400     1500VI"Pve�����R����R��B�������g�(� � ޾��<����&��%�R�����c
%@�4Ek@���]�k�KAW�� �����ZNe]��	�B}�2���X��jm.D�3���Ļ�v��e�������vz���d,��xt�{g�x���5�n��{�E�@�C��R�#������NX�����~�g��9���5t]�u�Jfߠڋ��y��es�3㘤�[`��њϏ_	�bK��ﴬxmF`G
1=.p��|�\��@_���c�}lV�.��*w\*���#ݸ�M���ۇ#���X�'���v���؆�l&�J�XlxVHYEB     227      f0�jrPp>��D�E&f�:�U80K(n�Y�ҧ�R?@�s�(�����O�p���������ϻ�_��M{����x)��Í!�Y��:~{b�`�����\�@�=����)���U1�Va�Xp��(��@M��n(�;L5m� ����F�q��䰞�A���B���X&ڑ�/i�\,�3�����>Q���k���I�:b��,�i�T㸞Q�m���u�&�����)Oa��ݔ1@