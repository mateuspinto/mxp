`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
CHSZsjlcQocQjtvAiF9ZFB15cfpGxJzTe5Z8HuvaBJl98Dlp9t/gIaKAzty88Neaf9/Ic4u5aGMA
Qc8E0a6sDEGsezZFUjZb/LYNiGxbf6CqDfn9G5EvuXiIN+r+fvF8BnYNeP1rEfI67LdnKRzvE7uh
iK2mSULh9JE2BaI+CG6wxCeO2bzM1yGgcSOtnoXKxJn2W1MUQLubHRyoFQeH2J6WdKOgW9GzeTXJ
/xcHQNnKFFn4/60Y2Pq2+WB5f3Iksagvq8cQ4W1ZT/uGPDjE7tNhNSWQA+hc5jM0G3xNjl7shWqG
hArz/hZ9Y93F+eQWyUL16UqHNZZ5NUfKSoUxsQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="koSkeMZzzdLsaTOulk0GwrctEOO2lhJ81UI79g8FJsY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23040)
`protect data_block
Km3X4kuvanKKZR5x+pqB0CUGwWHRhWkYm/zcSjDijeP7WRiINujuFbOCJAHl5EhotRHn+WwDTKy7
LdCVfuDdULaIzLznf1z0uaHh6r9lAMdr8jhSOcYH1jhfXlVB0JkTB929/8UoXNL2etu5cBB0wvy0
YI8RzvhdSiXKocYEqZVhR36Ua0PujNnQPQlYdJytsVLvGjJMBOzBRYyKjrIBs4xNpgT4Mqse+GNT
IBNk3brr4NPVn1BlYvqmevFIl/dptJpktGwhOE1umcRru8IJBvs0MkiRj4SFqd6LBlHgPQTXQzSe
li3MkToGCkKZl00jMkUGGysmwM+gGamUVGaS0FQzzjtAshIwTuMXjBgju0mvpBwWTT8KS3dn3FVA
/Fz0CFGEL1C5/Cw8ypmZHYbbFrLdwCp6Kz3GFiuay8AzxxNgD37k2rR0i9+DNTllW8Qcnfm20c0e
jb0N6q5rxX7FJ7tw4dMUR0l7B/WjX7TE4hl11m//i0Ck9xDDyMcxGpWg4aY8s3adS9/bAhMOF3H+
y0yqAoiBNuoc+caUUkWJaFJI5QMfacZGbby83Zt6qkMf08G7wFHAnO0K70VFKHtw6Q17aac6ka6E
1s0S/K4u5GXXyf7KDRXi6V5RHNaFajri3NoW7SvGvQzxwip4nSZDrv5btHkSzTGkSIUXVE8Joxwt
KMzUOTwfouqZTYeXuFmsaN0rxK/X5eBbIfxbXGW7TWi7VLq8iiYad/F4ofmD9x2geP/CRoVSgjnw
fEtdje+jP7Jk+JtXcSp6fQ8NVi1xXoWRqTRRnj2cJ52F47DoA/nr2F+Cpc/lL0nglVvTRL58sDUN
g8/tr/ivaJONR+p0KCk2PIcOOqQT0mzvQWRMWj1IwX5cleoWb7VgAAovvVN97+nMzdV+sR9t2FA7
IXSC7S75YW9CeRMakj27qoZP0UHKZb9OEDop1/HLsKucin9kMShNyiWkD+zzj40uKzZBUTmbe0Ot
Vn/clp3+Jds9HVxPqkitSQbnlOop3tv37+KJpZ2zC7PzvCEGUiY05ZwO4M9s5y2AkGTn8L6pezK3
gFCewsrd2wz9xKTqtWrUKTINDs6seughBOKfHM5UE+Nq9fvUgkdfTjYHyh0XqY2aQuuniEzrxOv9
bvK/cWrkOAoKJyHqF2gtqh/bJ59sawdxiWJLRVr8jgmUfJaGcqHtT2A8oxLir+FVlIyXhdMi3SBr
551mEPDqOrlo/W/OCzqmV9idL58L4xNiAc7NooXo0N2PuSl5M8xx3cIFezD0quw5svQC1GunWGzs
UhhvDkB2LWDd9N8vOBezIbwW8u8IRuT7ikwy/dpweaMPfIS54QNaN4dQkB5e8iCyotn4hk1ikeRF
Xc9677nOksNreUJ7WK/zMzVQ/j0iR2+u9Y18M0Bc+tq/JX7IcysjrW1FZ88wq63kAoI9IB8+A64V
nuR6+73KaeNuK/+X7RqfS0pHAdF/OcXpC/l7enh6/ljzh6eWXPCS3mGbaQTvSd9hR152jS/laOm7
Ii4KGHWPcIW4/LwJXNCpb2XGm8cRGlTfmQmXDRYnsAag5aVCHnCFnHvemRuxVtKt7yOvtd3z/LD9
ZF0m8ScPp73EOkBxwWtbl/Y5ABg2Hjj/xUiNMPpocheAoxmz/rE+iE2lXQQrsDTsCLv2xsvrLkZT
rJ5wnzvHvI49Tm8oanskjCu+4KkMfLmplETKy2uCx+qmqnAkNimx7c534HHvcVdF5kaYoR7tEvhZ
VoXGjxC5g+nMa25cyktV6m38a/IssiIeQMNn/drQRp3SflcGdPxKjAcD6S/ZLTTqRRO6FvSEWVwN
AVshiBieXgCdjRAKA0w/Dtbx3AqnQTXZunZZES3YJF2bKG4s/4bx2hmDTNXgVmE0SpBoCNt4BAFv
obyIdHlShI1NhN2S7ddtVFjpdntiyVF4GeHIPyHcvh8s3MzTqkZlaEoJx/2fk0bvEOhOqeubJuRr
meyh3+dF642OeohmYI/m9PjREb0puopFu9nJlXx/pqrjE+wAFSKfzJr3vQxTSL+Yj+fcSTqBGmMr
rVPALTPnoOttvVaCG3XhAJfwgmzmkPYI4daGPAAq6JohZl5RrNfbNgbAUFmgEZ1SVIqlHz4phDpP
PeKmv92DVxq6yQ/IQqa7qlKSsLclVEF4lxu8GBnsBlAKRZPHvK3tE7KN33MsWQ9fsT9B0HiJfvUB
HB3Awrye36D4G7/UnSZZy3hxCq6ErCiAPa85NOFhTeHpnhwZRnHRocm7D3gr2aFDjR2rEHc02wrc
DcXTcMn4ENdBq3H7bwy2lbmgleg9CLOPG373jWb97ioUMsOVu8i0Jtr9XgTIXor0dhzB1g4U80jm
YaaH29MOupErVRHtXUNYr6zUwS/GHDwOXLpd2MpoCodoXZUVRGZvdMpHoIi3exCmzah+yRyJVBAu
gnyl7X5w1XLlxf8H0TQaEo2FaVzSYbWQ/MylkjHSKOr/thxtrib7Erkr7zIKiRdEMiCV2WhAjOWw
GTBgacUjqggAiYcfok71BEkVy0lF1d9J/Wb9FGE9keKznlLvf1UmT1CaQm1c6Iy2xSoC38xsWVa7
uGjQg7hgmVgnRUZvyagGXDrGm5I5gNeW/SSn1O0Gh++LuEfGWdj5pdSQbrMerZNvea7Kna5lLa/+
ra/vZLPMi1pjwo7ZhP8mnfPnp7v87Krn2zwizucyojNa5XOAxfpY8ncEMhIcpVMcDtgH+7yTU9/+
yK7SWh7JdIKTY32uxINsZvXNdiIIiHryoHUSKIbGCcGYgyEevwrz+krcyoMCHlKDI89EpFUIy1lv
c8vCthadgJUsaPGEQl7mgJAZbRoNH5JpMFGRz+NHG3SNB/fVh0AITz7Nw91aJs/tP0wdWP/X3Bta
vmBOyzJ0BFatQtTgLki7/Fd6MKXVkFhlxul1ztMwXGhg+5poLUF5GrmjK7zV9PLzngN9LHLH/GN9
ExRk2eLxutQv4uxWbM/Q/NPWPizPNBoTCee/ZW66aJNfTpOS1HMUorKTxObAC+XWRPWvD6L7scPD
pMB25DoNMLEBw5ZCZbQLoKhGXOdWCwcjbLNoD/0eTl7lvys7NR9oI7yam2mtS8XJyS+bz/jjxO4Y
qc0CtLytl98BMHQUA9mshB2Uvmw5NP1IoVqy2NX0HvTpDM49Hd0g1OBdRHlG1ZKEEbWHXwlDlJ9v
YNhMPhvhJ28N0LRy3J8g7+1dl61Ez2qIYuOGfJ6CWd1DuUQjibcM5cGlxy1ThtwSlqf5iTmTAMsG
0OrVm5TQ0ga0cGmUhCleRS6xfGw98CO+MGE/+xDhx9OEiAuaP/I9VNh92OZRS1qZSLy7N9LLcjQ2
SCcZySIoNrT+H19uekuOkEcrayB6AgEDlnZ+0WaTPDYK1W70+5cLjuE/kGCd72PNseNdt3FSQc4Z
SDqYTBqwkQ1Xntytzn3PbY2LBWh/a7xcit4Rj7eXHAsVQf0dW39wWXzqQTNB+vkKKj9Q/ItxizuU
QijTbvBQEUBYOA96kFUdpLX5mD8bEjpKMYE/23aGlA+wxQZoLs5bFpnnJT8syhl/QKal59TCAjJb
12/P5uuFuaafqCuUNYv/bgPVQIGJj/vLc22Jq5FVTbtPXtUclMYaLp+Sfa05gXmJmX0nJxRUQs56
L3dk9hLfpYxv0fs6C4VtJgdvaR9e5i+ogjrIS1B1YSM5eyi9oyRAhsN7BwXdfD7TILWFcOJ4mFnY
juQ5gdQuyyvbsZ5PWus3SD6VMWOeYJbGZ3qIjePr04alOuwY+s7afpLqHsPFd+Y+K2VVvJ10s25t
A4NpbmI94tnA8n+0cfDHLrTBlKc6JU9HpRFoh4cQ/6IRksbgfdtF71K6eIp09Av8jzyIgSpj2qIu
4qG71rba49VYehjCsylJAhee/vgRyimm4L9FuKjcVB+PpZt/sgDTmiR854Xx4hHkbh20bJVnikhq
aISUimKo77XmLhsadgfjYeG+qK5QWs802I+snv7vCRhS3VSLXFgcHvidYDxDnVMM+TsXfJaIgQR1
cdTNC4l7MgPhHbKKH4+0uWMwbOuM3njtsICLp3zEQwMFR+NLd9zZJHDaTvFI23axQkC+FOaJftXp
6dQw3MVdACJPW3rCB05+fW3vY72OnzetsMmlD0JEbrcRoimnc5EDqVGUbTvbEG1phvXm3GrFhSkB
wpMekwVlltkm6XBMdIvpO/fKAZu17Nv1uu9v6m3+fRIWXv7wJHXIqqBjU7OwB426D6+j4s94YO5g
W1XJHq0tArdl1c0MTHTz04IUOgXUNjxARTdepMOoNCRko44ww5EClLX806IHiF/AV5ba2uiUOv43
frZqiWIsda86R1qWBWbS5aYkYAjyd9cOmHEU9B2f1GwpbJvKo7byH8U2/YSTXsBFs3HVHMg8JY63
PeMCBNxBovq1hr0XPweJg9ANVleLgAjNAuhj0YMnlqsMgE0YhYyF+imvvrZSl0ZMULbuJ7vyhaWM
df+cST2EoWBrY69MjBaghY/buZ/lKfoeCxWUDyWgZ3osUhXNLDHX6+eVQUTdgOv4Go8MJ9I79aVb
tRu6opYnwgbjDK+de2TIiHL0VZP4tP3GDRJMQp7gNOo/Ad758rh91C+paCLf/K90hTxaJm1d51jv
nR1woVRkfTTr/4RuFnlv1OXioKRI9+yh49UCrGAxoCd0cw2Ymx1DURvRkDObCwuBLf0CZjNu7Wpd
P9hyptcJ9WMoHniRK/AZyKMMNJ21gopPVpvevOcAHH3kqqf/e1X8Cq+hgB6I6ViCB60YohX9xsiE
0lZ27Cxi4d3B0yepUK0zjES7sjDr9n/jmjHP1IpHYn75Hr7B2e0/lmMrCVKU4mNCTLl4gWWbYiS0
mEzAxlfx8/Q7nqXNiiRmYW4/UhKWl6t0ayNZ+ootSrXVNd5ysrkqljB2Q+Ee8YGuItkzBQpO7Wkp
zBH5YwUDbRjKWbDQXnP04pAgwPwRqUpolmFxy4EoYRgkb7UqfRINjFjyu2lTwW/x170PPGNGadpH
1mRd57dvOfK5a4IqCvD4BBlgmgrCNBE0TR8mvCmfXrYwY/4+gxFxMi7RrVBYvkMS0bW4iaKnFc5X
VWxMPv8qNmnTdRKodWrQmNFB/SsmftYO8/KRfxVnez2BgYpbMWE031Coy2kH9u1lsfurLCFPHMeG
82dnTV2QSp2UasSjavEwgm2ldMxT7C7UB9dYie4Fhppn1VyXWskyP1HfQgNNH3C+DR6FHIBl1nq5
Rp2cN+GqH9LmF9WGOGhbk7hYNe7cU+9G105+aShU3enMseGYZe+pff5oGZ6IB8qM7zZfQtLPVpto
oAsJ2hhGprZkDCzt2jhgdaGFwtIdTogK/5EePlfGs2TvAt3KWrp4OxA2h1foBsXe/jbch71WihCl
9SNkE3bgEGfRBraLG8GyjigT8h2pJt3aKINiLvNO62jGxhCzBm9y8vWwtNmRvB4OPxQ54oyzEevC
awoq+FMYhDCLevjKkf8FkIwqJuU5n/2h8t2j23AKo391k7XvNqbRZte+lIffpZvo8xNhFfZJI7Ox
ZltgPdyCnKClwchgk8kyKDmNKoALm/sI1bhIzsIwdw7BsszzT7ghk9GvCL+ZER/wPapN6xLQfRtY
ud/KbYZaex2Xatxa1VQGM1kYzVNp1yi9xheJVewvsRcsdfcsPuQGWigPLbZHv1rIlk/lZ48a7cqC
ecFXMiBdyqQQciwXltwLzB+yCiLqyPNsDdcX8YvaWzeOgCzVzN1W4jVDVYFnHoy2euA4qfdF7K/P
/FpbvUvP+dcYc8zdMFivAWA3aAa5WBKCSlDVkr4EM3XEsnwH50iftqnGHcamxqeVvCs7/Vzn+RuY
Phzi5BMj4sN5iUXS7yu9R5razOe3gGzb4M6Xi5W4azEprxmltnjmPM3stS3bSoO4T5DOpHRGF511
CbiY2pNEb6K7/UKxLopPuJiAEzQjfTxTEMa6hf6e0W8jn/lyZmk4H+Yf7dIRWB2RRfw8qfBKgGOa
Y33ESTbcHwHj3i+nMwV7VUSkMoitMC6sMmHAG8CNXIwFCt5CkpDeIUdFE/nNKf4qUQe7po6U4Wjp
alLhITiJPY2KHq10mRmjT73gpiso9PQvExWvR6lzIYlPut7EF9d9tFfVfUS1rMp00qiWyEpj04+q
l5+IPkydhVq6OKLTmvUWU4F4O/pReQIWxZaQ2pvlmMU5cUY0Hb6bLbWjjHMeKPcLMbCwcXRUW9yH
dcNU7lj6+SHxGnzgO0bqXGNMCtFBMJZXvO2SBOJ8/iyL0sELW2Ecq8fDcV/ycvE45YyZgGPhFrUd
8CMEBmxnHndKA8dck6wELFJ16MtW91Xq4Jqfki25ZmgHPaqur4WnHD19zapuqwQlhnBTqkBgqx5F
1tKvw+7MGlIoIYklJcFQvpdSIVCUUJ0DaE4duzN1aONiBpovaJNxYBPKvtQLZsFrNLPuPXcBPyGc
dqnDcgWm0gQxN5sOzjqF6I43y4d+YKqofhu4tY9f4an5yI5b17y5EFHz7Oe3mkxr8SgtmdAOBwyI
YmWAgrpgOMiv4ald29wFgfjrN10C9Ffo5OHhHq+MYqW/H6/jvvzU2E2BP4d0lHlbcGH/imkeyv0n
t6WR5fU2zDC6J1p4sa1SnDQDgeWLw1nCbRndexMrCdZVT6YNakv8fIT8HE70rJ/0Z6vZlE5sDVvx
Qu26IMaYyFaE9mpT6KyY4am6nHk7VISHcRfyrN/9c1jM55qYlUFL8WpeVWcbgnfsHVtHia+tGWpP
e+lEa4DHfnJeQWbWDlBTJdVatw/4fdl4byyKmLPqK/BCmKPYccetBMx/rsv0+GlIdMpJ9GaGufNz
Xv5fyqZk00pG4ms8wBRMBq8+58ntiZ2qPAjStfa/d4PNY2hG5YQlvs1oR9cxplYu+8RScXQremmw
qtd3FPZJYE1YG/uH8haQSUSmwe/0FHmFNtq500sSv5lt4xJ/fLd8GXSqTDCBc1tiXkMtWsjKAlHB
ifvaXKNACVIn7NQOw+ddNOu1GtVKPIVSQlfTibkY+o6jGgF/1JX/UYMie6E48ciaAH8/fgyQJTot
2RhtXyve+4oYyO4//N/DNnxYdRg6lkreflka5f9h6uf8O8oJnqzmddhcYOOSa5uoZ4tChxLgfEvS
ZixWZZpsXPUeV+EQNypP0mND0Wm5IKfzDv7ym1W84yQEWr7TJb3v0gxPpy8AgJmy3zdjLi70UdOT
BK3gCQSEFJSlKLg/Kl2c8uEVdTDVNVZ2qVjd7ue/3CBBsU/npMobuAuXKU+LEahs/V52TyAG6+Qq
XcuuCG5ySfkfrnBj/ZdJML4eHISasYPFYw+ubWF9pcUKEDkFBCZ1pbmwef1VkBZ27I+YBml1RcNf
SNYF6XItuHjhVlA2btDx+/3RwF2euS1N8T33K+eZzg8cf44TsqDchjeiUfvRC/Ze/2bzMfMCl9lN
2A3T3Q3c+UqTIGeC6xmlw7Nqqmi4bc1oBXiQuiOkXZBT8crRe2GZbRz9qDqw+7kr2hq1xqUvrj+K
RwoFWwjPedHUuggIPoaSksprBEv9L4hZ5RyfuZ/BwXt3I5bC1UBoAPvjebgm3UbPxgm6zzM+rNM9
LPSHgV8dc2lcJ+ZgJ1hGkVtvCoJi4SP9roqqA9Kk2wG1gmZXKVuvRILtHpJsqDh7z8wQXFoaa1YG
DBZe0m8Hd2xZeTqrN6dqlvz+lXb4IT53sCp6w51eWeO5MV7LNClbIAqICOwE7C0M3Nrkxa80/492
WB5Z6eL5uU6TzSlccEE0/4nbeM9HpBnQ7lLxO5XWMxMTn2y4yM01N0hS6mtR6ARs/OXvvgZSajuD
X8LpBRxophvu1mW8r8zJYdjLnmCIboFXubZ1W+lWIOMQamwAUgVjsdNZu1b6bTLACS8j2VoY19RF
/CsZFaYahXKRbaaA36BcwCj5DKsmtzbQ2z69+41tOcJa5aANPuHCvsEytC33HbUNtv9zLjFJapOH
tSy9sKp6qfVQneFEZkImitn7H30tWUuQ1LnPqtkDJ0kcLt7iyqlubDQsTYqQB8Kz/gMwEEgfsjg/
/RCaheffSYocnExQLwYNEE1GffQP/G5lHkasKcHdcM4sbPFtyMRMUdnpPr0QB0wbacMdOcVW1GcH
schXUyiKzrndAAKymMsnyUUenmgLmbezksNf4qKpp2yjADvLeJbWQHaVeI0JtlccUGfuHa3JK2x5
tFzpu1hS5+LYdMe0fp1iMBRuFwVISTc+AgyWBoR17tfQ/aq7Qg9tCNqj4dh0/UUJ3domh1VD+L+u
8qJKAl5OgmUE1SKRp4tdaEAn/HcaQFSEsnLWsRBvCrEStmhA/gpf56bu3qOfFYu//W24kGS3BBxx
1dv32lVtv7xj6e7/N1iQhit2vy21CckcSixDFBuMDhIp1TEQMDvXefYHgtY+GzSAYQRRMcdpuhtb
PdaPvJ/Qf/4+Rv6yhPZQcrqnHJyk9nx9eeIHkjjmrgj/JIGMw4K7lCBvOT5eguo4OGX0iQGav9UA
ledR3IR71xquNYIVLWRxQ5aBf7C42a//6Wb7l7baTe3zzyuXeFJMJaJDRqT390l/kubZNWC3L8dj
Mat3IIQEfAa2eqKo38Cj/RR8vkSSG9F5/MvY1NFtdvr47KNmFWj1Ya3XNl6lu8ZAJwvyAHQ1YeRt
cgmyXesTCVF2rjKiytVSdne4hhFccMzB20YULVwCjGwdbQ8CfyGToyWkv3sslkPkXfS53+nhIgwr
B0egwFPuiBx0CKXs9EEZ1hsvn9IOvVqVdSjyfEf26dbtkFu/m1HKe9Q4V/dxfckcP+SC5TOETBtP
FhOn0G2WC4O94pzwIVCPObsEmD9IWmNmra4DCRyduMsccDVvNwlKWNG2FDnCkOddoQwWhfrGGLzH
4C6S6o7gWjg7KkiSSzcvaKYJfUsAKJBhJOdUX3DMhtmbQ/QaJnXY6WkmoskJkcTZkEKIINVLQ/ji
xvvHtVtUsqmuKkwR2IXCMDf6zJFIYWBI4KX7gMJTZX9u/v9aq4do/RvTZUhNUsB6+KJggWj7spK3
/e3YxJfgbZm34jiOkjlO0o0TCP+QR9IEgt8W8oUGz28nseYV2V2Mg3Kp1fQB7/9B67eJKaWPTg9J
5E6c+etP/t14KqrG2eVOQ1rCjIc3fvYFev9z7qKXGe8kKFFOJIHinlqD5K15r7PZTc4wlKbAKYD8
NX/RhFRCVU6chtRCWX+rVvcFZUY+MsMWRyGGdo8UQr0MOMLKQJ4nEGZJG+UeR+2fJr44wwfylOJm
D/CIALqPMDYYLSHt90LctchtI7LVLcZl2hg7sQNlmixSj2AotHJ6k6D7SJrzQHJ5+KzMcQarveWW
7ENRsdyz8+h/6b4WbXLQVkynxxJNAnQEoR3aD/mBB3I16wTmSrakAqUJ2HGiKyqLkMbhX99Rp+yI
xNhKDUlhutHhQev8N9vzQLAYc+EwirFg78zJoCLPRneeETfuPFQyjhd3zFgwcxtfEKnHVH9r11qp
zuxZTiD4h1DA6JQB239KUYUckP+HRhiOmWmgp6PLERstMPSghpqg3e1E9fRWAHD8fPLmICsyA+H3
1wNcAp1hztN5oU85/BEwExVJT7j75aJghf6UopklXThT++MFx4z6bhekpuN5zUbx3DdMXwaC3Fgi
PJoQGuPeBbBxVgQKlSUvgkrDwCTwWUJI0D7RcdRPj0il9OHufMRMqSt5m978jV1mGTWHDfode02o
s5vfFJq01SUq+0t9J5KJ90YRbsNjgZxTMow/ZCjI/rOlk0oUzdw4UUpZTC+OP6zKRmvVzOZEOJHw
u+T0KE2YN/1Ck5HqlM0RoFsIrP5jbtEw7zzzXP+QHDxEdnIlCOpRjMA4Hd6hyKpDfdEB90kfZmyi
5ibFNElreCYALPIqR5+SsIxhEutp6GnzjLq3lQDH2a3EBq4KzxhNajaq2/iXeUtdlxqjFQj13evU
9GPG11iDvuewZFOcn1/PARbEpRDUVmmYm29y/Hf51Z+J895rpByIe0kAIDrR9313/vpuI2/mWgmD
tdFi1OuzqTq4i/W4+k+Vzwe8Cj5ziyWVVV4+GJAtY/SwRxOKTokuaKuoC8LmCSlBtpxpivmLD9fo
aV7UlHGO7oZv3SfCjabYWyYl9U5cl9WHqkA0IJxoEnT3gSaih0H8I5XctyBGFMHwjWtI27U+qXP9
D3YuFFNm7qDGzYSw2BqztHzkRFaRyPFF1tgtPYXR00hblW57D7mXhCX1kW4I+9Eqb249gL8rFlbc
jV8XkrYVIynqueRVBW8/XySQoyAZuxkdAvgIEn8DzLiS3VeZZS//72aESOXhXewZmYKvXyV5rUbf
eRnUhJk9NsjbyxaSCy4CK7hL9YE9EYV8uBZUVNgmsR4+zpev4/kToa/3JQgDjn3bxb8gxmMWJgs8
wC5d+E+Nc/yu/DJeHSNz3Uu5U9Hk/HJa3unrxHOQjR8d717+EVM0rwCTrJbRj0yLK3Vnl3MLNp8g
CGLVIwqAUpxR2/Gat08F6IaQeZUSAH0PyHEAxUJ1xOYZ2dTuFeugbGtZMWceZpbryqds78g2eWSI
QZ855D9Zk46qHbAH3c78018GQxupAr2ngTikKHMM5bvP9mrwDbVRd/ldnIs5NDL9MQkRW195gknm
80r0Vd26OLm0EpucVRhXLdnXSgEYLj0diCv40HuK6GMkVJdGXJtw2IMxwdejVEOY1iIHoB+SIpkL
/AodxKYxbnkP968FAyFjAwTp1YUKDmElitu6UN8+Go0O4OrwAKxGKt9WFKI7KA7prgERdPOA0Dqk
aoBHRlW3ZLtO79hYdQpXR5YE89DDoobiyOT4xbQ12qvkGMrOaMo+sG+ef6kCsGLobM/uHi/H6Kn1
2j9+L7D5sNZKg/5gTuuVm2rhlT7GABdSUXbcPQXWlDH968qSJ1opxp+zwvzd+0DA/RGoalPgGvwf
kJKlm5u1aEuXjz+536KvijsDNCWap4BtkB3Dx+gKdTayl4cxwlW2sbZzrFBi5x+jDLlzRzJ69UsW
IkkzV1XoX6rvQzbbTArYFBY6pTIIYxeFHLND32JzM6uHqHH4y+WcSpyn0GPA8bZ6/NCmXcwLultU
3HTypbPGCZIgHdsZkehGezH43QPbpYkLPZ3xgkZSZRa8/BGH2eYIZe/CNDF5mgfUlnkQlnaIfz6T
SFWuL0H7GJEeiGqe1K5qHuInhW5ks0EZAkAAHgvoYwti52iNl3BCju2IxZvgnSZDGGQxHz7LIGrS
lh9X0qCK/Ja7FLK6qECyBQ17ZrJ/lzf1TUhPi0loGh7Dl2wg6F51ddL8e//mWfKWjNzx1z+zXfWv
Rpgj03mPZNQ4A4dXOCKER98TUgQPry/azc+Y0bX2+wXzWZEzN8B0jVz0mcLO6yVZ3AEshk1yT5u3
L/yXfTTAV13TDqH/6dnBYYNtceerjK3MMRhwiaWQyKn2rYld84pNoGmwD97Z7t+gxJ12iY8QMTU8
6qvLWYq4q5Yj59+R/90AZohjCfAdiiyxcBBzxs1KSClcigTgrA1hto4gqvKDc6c+8v3YBm/XDCZ1
VfpVTKHGD4skppCu7dJ6n8Wi3uGArC65pzy1ZBNcEne4ZkQDSC0Omlp6kQG5iNVHH+JgxkdfLu2S
aNnT+gI+uHfq8ACTwhp70/bmL5MpVHl99zX8x7iP5BAiQ3wqa0/iUmfyBY7x388amz249XtIaxv3
7Fwvs4JQD4LmbsxlK7tpfDDR3L4gZ+emX8F9Rt2bIGj+VPDGYpfj5LtI0So3wmoISnlaUhVnf5nY
xbpTc7svvwnmaKtu3SiRNkgY+pqXYf/Kf4ae+LBMyQm6HIhkr7pbh4kF0hUeP3aM5YsSFmZLwcyn
/0yvT50n8mhcegvW+3xjWE8yxApBQkIgXxAFD61ro4Nbimse2gHZ5U8jKIz273sM8rG6QVWpv1e4
Es9mGmmWjoO2LnjTMX5+c8XPVQcfOdRg218ty6UaObX2/jsW51/UHy1kmfPbbr2PBiY4hbM056AL
OGbDkYdwfjjoVdNl3mVsP4ktK6oyVfKgYTRHV7fn3k3DLe1/lzN+qBCOw7l9Z033JxUYmqKwHt1B
eU2uZ9h3tC1IPGzVN3eRAwJ1Zj+b44HhmG3RZcH3ftVhiPO43b+slTtu7fC/5HRskqct+i5UIFSH
LLIPCWzsiB7ANlQoeH3kyduqoA58fW7fLIrtn1TP3F5+WKEgRVH+jJZjW0W3oqc8dpwcyhqvT/a+
9NmjR+hkdcWzJkVREsSLLCc4bS2fz1DqyiBIoNxklGRFCT0MJK42vVKRlg1qG76nraZTpLElMxhU
WqZcyu2fWqmJLWlhcg42PHhs730WPoKQGkHGj4Te78Fqq+DJK77JO5ebwN7b0Bo0uWTX+JYtaYQu
fHOU8z7lvVX4ocgAt7BzHhxCOhj9sPOO9QY2anZlWd8hE5X5hFJQZr5DdR6r0m9oAdtUxoDi5nMJ
rRqh02n+BGy3+88GKWOb+0qP2X+DFE3Xe+3Dc4zHWPDaXUhDpyO5ydQAYW0YCR9UVkqS1I4xkku1
OBTUmSGvDBVpj3nknM3RexON1IdI6PIh6RSQVhYzOTUTzd2eZc7++WvNMl4whxF/qB2fFsPywC5O
1YycMtFB5KO+q2z3drTp5lv9KC0F9MsT5t4YA6b0/EXPHS8LIRS2ZuHN94dGV7o3GnmvtuXdod7M
q1zb/w0gn4D+F9iub1y5IlkZBmtpKPnmqrOpabYcvrz5GwnJwfpch0hoFOp0evUJdgvTYHYAi42g
4cHcTs/ASjErfbuffW8l3vSUW40aB/XowZn8DKvZooNF9kzlxys1kt61KiptsbP0pf/3wfaeV0C7
qT30cHQEzE8B1fxNMMikjVDk9Q+cuSkUp3Pezdq8wm8hoZLrr3hjHN1IVtKB7P6F42Op7efLJOMw
N6sr737sIwh6W7cWOyMr8aUmW2Rt5uzteci7VdocPxiYBs9XMdZm5hUfo0f66SwZGCzUJG8aWCcJ
mM8B1QfUUPJDR7d6znvXvPiveHB3pfEBhgE0/tGEsf2v28bYgdRw83kXRuDxoh1sBSZnuYL4dlBi
2ZG3mV9zukCVb2irdRpoEhAtDJ1xA80gMqw3bn/wGuSjSgVoLwqARxKHBMlPs3bJUqBJsDSMODj1
jFdOkOqFhWXTPJUjo790mKtqor9siQ3npmyyvPIA38WrPr4UUVrYh8P7paZ3juOlHEDhtczbFZEl
ZJrRwHmrrXnXgmhCoirQMKAUa7nJpiOm/Q7ZnfWcRwQDx4XSTJpODqawxQxMlDy/wd8L7VPSY8o6
XtEiiNyzGDLoqp2WhX5InTRyD3j9QeB6EB5z60t57W8qDTnw5BXvOb3JGsH1WB6spEUIxNlmIXku
39/sMcUWjHY5swDPrKjNJWZRzIaFztYWAwCDiCw5LJ2zaLPKOQMi4cw+gHYylJLseNh0PNgJZg+1
AR95XCPCRA9z3cvlsiDs2rwOJwccLyn3x/ZdWLX0HfIqxBeUkOyhnWxsgWt630ONG4fX51N5Auec
SFv2XXMOfs1PDJy+anFUR32zR4HaCFRwO+f57Q7Gx0bkw159OCa53Masffbji5VCRJvWs6Kv6B6l
HmgL1shEg70ojAslVRmk+nYEzyqwGoKw5tUPPUVlI1ojnn5Wh4yTEJpO0ncX3TjYdNjHlCWwtSOb
aCqHr/GXPghRCxm3J5cUrguI++PNyF3NcULpu2i6IBHyhzp3bIXpONfdrqnKtxkkTivfttN4E/AP
TANfXKnpEeYCQ+egpjqb9WENDieBO+5cxlW8+oeTW5nnra7qBaoQm7ZzAltPsvt2uTALPeKxqZIC
B3CkDUBUMswxBmvM20bVxBVWYa/46ndBwGkasAFrjzFAlZVDKNpyUnx3KwA509YFUlJwW0XChiIl
VTd/r+rcLqBrbfExDi+FY2FyeyxI5zH+7AwI9s/qBTo7L5sq5NnqQr07LldWTDrrEAuD5uRKyf0y
aVicZ+Mq60R/q6aPlYNDFvCDjhijhWwb5tQUHoXH+zXudTxB7zWoYwZLKhmiKNufYlCeVPPL5902
iDDl05lwwfLQsaESnUSOGm6R6KhOHN7FA5y46SvLEcAgmRIRmS5KTlzGhqE82RhhCjwC+Y7o2DAd
EJk6mTC34AQzcHbmzUeiN4lhm8DqSN9ZiN/YClBa1ElFABSekfglT0rN3bz4CAT1Q3AbbQI50fn/
gyxbaKGLFlL55K10l8bD3xPF2FsDaB+AfZU48anQ57A15ZCe6ENVehqZs6d6WFNt5OaGdMJgGZLU
6J1epBuUILJr7UxROj/S89aeQrEZXhWYLBZSSkghr2yR0nIQXTgxAIYH++u6k274411A98QHaOQ4
hsfMNEyCql0954d8sV2Ek6hVoz5ON25qK0RPuafXmF+docLqrwnGaWFmJ/FzQQC5sLzIcV1vsY9g
BAL2uxkrNh6DRktLISzuSKqCGT+hIvtiYXl2DXKUI5J1SX9jN978bPz3bkLgbMaIliGxkjJwir0J
PSzScYYWLnXoRCpZCbTtX5t+5xUGYO3jRI09uUimd2efOvmIsM1HS6UIW+4jlbQdZdB0dZs+Vqnl
0QBvrO6N2xZMvFmgMRFA740Ft2V2ikB2eilHmF7UI8ztoWgcE98T5uPf5oWZA3tfFPtQE7zP0XE2
mhr9aHF9kOji0C7yYCkGdotaw7RVKd2u6ibwazzAkYNU+fQNUzY9HKALNojMaiD+JG/ty+canl9D
2SKKB+u4NWR9TdHjxOE6OiJUY9+PJJ1qY/7qqrmEB5CR0wHrjqelR1zCR2ZzA7JNfJHTPlBSFYE4
i5TdEPipqZKrIQ+MZ/HCPMpPs3EE/epTepDOTfp++D9hzDwz2xiohVSPsyusSO/JX5gn1Xq/LmUQ
MLPko1SsqujSGQzt9nAaxORrv/uMHAeN7NpVcvcEbq8y3sp7OsQZ27q1pcURbaBMiPJ5LaIQp7MV
prJTJTBKLWhIIOhuz8RIg5XzTKDenIFF88p/0ge62B+Qp1OwZIA5LfEPbAN7ceQlms3aw2XlZN2k
CYoDrWGB5Vpc8BYYsjFO0BwvDE9ov9SGZ7PLvLMnGv0fRajJOv0R7uhwZTk6Z3jNPe8LdeJdbRYx
ieT5M6MLvahbQHiEW3DS0RCzRBHS4IjDVDLWeDeRYikSLMhV1IffOXqLp3qqVlm/McBFMt0qfIz0
XUP+1ethrwHgRIWvGLZnptNboiKYgN9vtN0SYOpq5X4H5R9uE4HiZtd++QAzXa9BnJjkyaOuNXZH
F0arGIBEPDx64CDOT7SQ5MO30Pdt2mUC0A41JBATU/HYZJ9WtOhPeDtmjhAaY0u2sSQMrMu0twMs
WAlyllBmB1fr8j3gtLs+daZL7sS8Cw6ZXefWGClIEUunj1SyPJ1YJ3mbX4NCzHzC+pppOoCbcFQs
PWb+NOSgDbyfvT+tjQY4B26oGZ1zpkMpRp4rqYUjLEIloFVaw3i7TCI7O5p1ivyaFF8QPr0Zbp4M
uCoxH1XllYTIukPqwERLq+Mo2GC84kX4KnaqEKvowpJfWDP8zajVboPzhcRyIcKn0Wps5cUuUtWG
66KyB25JhHu2jUSQcPcIlxudCT9hofV1Mk9fS1O91ry0IgJYPm+BDLsz4lYo7eLcHWWhCbmvm6jM
SJlBcEF6A8nZCfqPBVpSrU/KnIv6ShzO5YH4Lo5xfTjun3ybWTg1vgQ7gadgEmqFMCkibizYjC0v
fGdNmNdZl6IfQ7foKWn0DE+NAh8VemFQP0V+uMAL+bpoGal8J3p0iyKlCV/fcCpjA3g1//NDYM8X
dp2nQDpC5c2i2dJgN0j3zvINf7dNVR2Cn/C6D+HRE5YNEoAIwMtJ9N6fsbueod532Wvki6h2su9f
ZvCBuZAflwNfwM9emNnpTuKrBu/cg7FvZcb0fbGC+3bLlj5db5c/cTS++FHlbOkAsQ5adQR+biGv
aKL9aSPO8ln5ziHEVp3maQr37YjDQ0nvt/w+bqSkYjqomfg3bNHJEnOe/xR0MxviyQVDW6fyg3Pe
avVRXlYj2DxmLe91g9Jk9/l80w/i8R423i3XFCZy2eXgTjAHBdxT/8D1hJhPOTo4RE9k6mdHSqNV
HElUeZbyZ5S+mN2Xx6POBE7UMkpUnMeVPUpkdQpW2Z+WHKn4f5WToOr7iw/Eov27fSvebrAs8Uit
6A5ivJGFpen+BfLcnPjiMp1vdTVxNqqxpnQ/pxZp1ccVN0FT/TwiqNpeZO3MB3Jh0LYEWnclptqg
7GlFeeiWz+dJYTAVsjnD7kyARYq5ej1gyIjhhWPI0VoxCx6BmiMCtDjHKTyQM76DcTURHfYdtMSs
C1SQVjHWyvTbH53qlEBkLWIMWH3JNC2zye6HL/CqW3XpGg870nHO5p0RjjhWKD7cP7kjRE+oXGpw
vye/dAvVQcgVl0dyp3zedQbm0ucYp9NI89szNX8k46TMqNfKLMSDrxdraI2GU9T/WdfbsaGX6oI4
K2W6w4BtsrnP33Lg6yMc6IlANlXZlh+G/K3cZyC+EbkgBgsUPSKSn9PNOHenhWUGx71wkrR4vRn3
P7S1BwrpzeFTjJoNP2dFAyOA1OS2z1tkigUMWcNvo+fAucz0k7juOt6ZrHxRiiXEF48GuElRoTNf
eTLWWI3+eOud614nHBztiZD6DGnR9tYBx8wKza8gpr+8nu6hokhTnC1YVIA6QfKHJKrt50aOOifc
8SfpD2c/AM9NKx4a5yaixhfGG+wJA7V4ZapGT57/LZiL1IdN0+W6oNV3Uw6K6pcpcD5e7z+umUX7
OQFBAT2jVKAHuVAV52LNt41y2TGqjhCYaOwloduZcr3Gka/B1kUwuNC02vzI9K/LQc7Yssy8eQ2u
jH4geew0biA29Ubhidp0YR7fQ1+ReoDGcVKUApZZNz705wQ5Y2xOSzqaPY6SFLRDAvBJVC6PopKy
Vs5lyRDt2+0pO5xRphOR/EivWtKqEuCuNwkCyFBC4Auv3hJ3KC0LlvdwzL+XEw3xd+cUfI0U5suK
txEcFeq5MLJX95wt61xH7E6B0160PKe2GEsm53L5FlF7ih2mb3soFBWPDz3iO1VMyGHYlmRItUE0
opI9s6V6R2m85C7yQd1vHrIRZW1N4bk7iMQouSJi1rsB+6IcyrCYCJaeHZK03jsh/RRv+c+h7Jm3
h50+365WobpTfpfaxjlajGv1qk5QDERIERu9vFs5+HcI86PG8SLMsLu1uQho2o0wq67EUu+sPJY9
t88cSOWIP86pgRrvO3yTq56n+krNOncTC+28Q8Ha4+6HfvzX2xHki6S5Rl8Qv3MCrbj6zfRtLGgg
tU0SYueS4sLdF2YZsVkYNkb+ZbLa9wou3PUlbd9Dufhpy7dxY17kdeHAXM9hc4h6Wp/d6bwPlPu1
a+zzpArMVvlDRdV9YUDMY0sl+Zm1tNOd/4sXlsrnUMMw8nlDele/PUJFNO0VjZsFThizg0O5PK9g
KTifPamhy8+ha6m8w78BaRVrJ+w4HmXXoyadHybINc4g8bQS1JYErDg1SCGdqd8G0NfSnf9XpSh1
cgTevqHI+2h5uI7GCkDtUIwTutmjnFHxjOO1WBG23HlOyhdYDGC1uCdHWkNhJy/dYIz9EvljfZFl
Sm6k4TsW0hNI/BMDnHQ00tYrSpK75cY6hnLq0yEhXCCq7M7xz7IK0knInfDpSNh+MT29FYcBIZSD
Mecbp7sXBppWAAtOxIVl/WfqMVcWamodw3C63HMk8e43d65vcs50X+J6uLqLp+P4zXcfuOi+HdFx
lLenvirfGD2DYsKRxXqF8jDBs6rJyAkC2PnB5BAZBOLoG0gbfZGQpGHI9oq3BQ6BHb42SiftMlq+
jbRL8bzXpKQ0ZG63FdWr7xkbuKTXxyA0oS61a2/4bw1GSMYIWjl93fAWRvCY706PjoSYpICWfHj1
9Bi7X8ahsfbEjHm6d0MPCgB2cynltog2Uc1RVFAehVcW4vg/zONwBOt5JiVv20Q8S9liwyUCYto5
NThApfMjOz1RaVxRAPezl5zsFS9Sotgx6uckatn2lw3ARvlWdqzB2I0XDSBL1B6/4rdXInSf49mK
gPb3EIcQ44alm9n5ReAGvcXVUm4leyxzKsxxYMEHGFDGzN0N98cwyi6snd06seanEhmsmr52ZlNN
pfWJej5Y1QRAo1hOHhr4htHqNFlERUL7qXn1vV4TvsCWwCJN5rdhIJyS3kMIBZW6VMVlng+VXlAv
X9++5Kmi9+LxeuUOV3OUKbqCMCb0yFRsCkv7pXMGjf2bRhFIxuAlGGTB2yNKFsBvxSW6Vamwdfiy
Ksa/yktjs+OiOWYljMzIa+MPzAj3D5HGIJtdjlGnWLPkaeVMUSt3pq0CkpmLBzFHB7ajZ9ohzfft
NfAKwlbzNEIkd9jQVnglYud5lHLrzpjs5sLNp2DUxxNObY0Pnf7II17qs3KojT+ko8WIuGipKa4I
VvXR8Uy4e3LLZ8zbPdv/y007xlJg+ZE81mUWoHisoJQZIH12JXNKNzLRuU/BqGPUF/BczVpqc+Tu
KKif/1VKm5kamzXO7ULpPes+KGd5sZGDKvZ9VFW0FSu8yBCmBoAjiZGA50Gp2p3mNmJRe1mMW7lw
B0H881CjgCWgBVd18Zx7sIDYn1m6VhtXq0gsHplHyuZ3OLMEbF034Ywc5xG+PbVvtTAKkhzzueuJ
mgzRdEurGXrdaKFmvcC7iYw3bEFRRhcRWz9SM4tao/48lCyepioORdxeYmXimLHNvzTu3nRpAmSa
5i5YzfVV69aMXtHWu66LP6lpYnNDdtaP4r/5t8lsmBHCdp/EwFBdSLrZsTKykjTn6ZnwPuYDGExV
N6roMWEvEtSqrO2kkeAWvCoM4a/3iBo1bzjUVouN4gFIN0goaPgG4VDrxcLzDUG3V6FfMTEamLFN
k8g2n+sk4u89We3MUeLr3ljQerdA6jwk74Vy0wzAJx8eq5ANtFXtSgW7r0JJvSc+T+qffhkWATag
or/SuZPngiYdUCifX2Fmf0LLeovN5vKwDlt6fb01SoCeIeZHsLC58FKxjj839UwJm6DToJZaZid5
tLmbhMu4ZABt1vhnbJDKTbk5LeQ3mFo72DSsCwykuMyV2iu+5bhpNf00UGCG8AOZk58E84F7oavl
z0XMgq+JYQs3El788lISh3gJR3xwJj4qrXVWllQaFh3QJSuuKQ9gc/6q917RNK89VGwlqD3jmubN
2gXaBVXt5+kMeO9Nr6INXJLaEk3EN5Et5bbOIzF2VRcNFphqxGPydumMVuB3joNFXPWmgY6NGhwd
2+GV6MChkK6c6QZ5V+n99F7cvIa5Q4Qr7zJp8dv3hR5tODCyHK04g+3yZGNj3kE24/EvGfKk44Vj
g+S7+WM+m+aWp5F++GQhoDKLQllj8bOupv9qOMha8+ODcrZ2eu/bAD8HmxB6TCmTSGjAVajrUVNu
HBS52cVLjGduiS8GPtDyroLwA2A69xmL9XmFUXfHwy+2fyAvs02QxEYCF88W6OEBRae6UDnnE1jT
+wEOXrfoPDaUSrKPpVur2tQpGPaWmGkZCTzcEbU/DUmmo1ac0J5dINXGGkIbBQ9X0UCb/qauCjST
G+q7JCI3+DhockQDEEv+soLnN0UTh7EAMIfbOUXmYEiyg0bKMsHU+jbciYLKGbJOzSTD6mFhrJiv
MfLABo+FsPG9QDaNyi5zLFrhPD7qkWr7rMdnUStSIKLEEsujooZSmzRWhRRwWAe+6mV4yQrtjMgg
0Rf5qSOgMRL8lTlQ0QlI767WFcrQYdijUSCHRaXIz9k3OdCpYFVap5C/jUwWR69Nk4rhHChzccFg
iWM32qsZsLoGSb4vEkvIDIf0Iq4d7+dcrLXL9pXLUuU7n89IuxHFAlZ3KEkcLJItw+NNEQmSB/eA
QCSI2TZQxFcI/HtBS05nfb/OpjN7RL5GglmQXj5ofyB8Mjo7Ky0Hgr31cfk1BvjSjvSrTMR7fteG
VpKdAnZkroP5A8QA5UQ0JnWxRucDQ/iXfeKob8Ml4oRwXPpxQaJbBE4fHUPw9uGzD3lRzZ9xkfX6
d6nOrSnuWyPk/9V3X81HMLzzjfuK1Z4zJQj6ZY7Uf23blpWz1T5QJBwUfYUgquAK5MCNTI3WpHLU
jM/cnMC7CaMQiq0QWQdwDcujbv5Pdbf5X1hOjs1uzsn2s3TOziMa3V63aKPNDxYUujeWRulvGUst
lwzx4biOFJGrNFK8Ozgd7csVKHFOZmyQ5lb0fPV2ln5iXS/U59iS58t/67C7AZ4hRnOfkje8ziDq
ILjhvxYI+6SIQ9rp+snOvmdlvX9aFviFYPLQ2mYxgX1vpcvz9rGizo8EZIeGF0Z6MwYEaUPOWahf
frGT/3SFaPIOWwRtbGoPJeYkwtn6tW6XAZTW8gOwnLDWO/FLbc0IG58dXTq2fysDhCnMdetX+w1g
yx+ij4FHBvp51cD+UgSMrGJT1wLQYeSgSgu1aqtZBve5TizdSa6uydqDNWSTOCKeX5WaBk0hU+W5
RJEQC/UAXqaWN/vadCvLI2A5x9bibQ/jwe+TdstuDiZIjyUDpMIhOHWkUgpYkKIurpQ0vJHkE/AR
ooxGhsqgcti+4pilSyiJmAAODR7SuHCkMkPA0GzDB8iNa28uefJr0ZF4b5daH/Uxkn+pKJxBg4Xa
x317a3B+CaPxKc7cXvv3ym3OsbiOmL1Cb9Ny99xNT6BSETbu8qwSh+GIJyr1eWeOaKhR+Zsn/YT7
Jddv3gPuBTAS5/Irq3QAFQHul6ilkusnnNQwYfJW5gDvOrbh9E4ZDeylxN5HnJ/hQzjYiT1MixeZ
a8ufEGBD17XySXknlXtWv1hkDaUaqsezsnEqDRg8S6VRgSrTBrtX0tRwYcJkPiK1ipbgJ82dAcmo
iAUOpU4jWQGjOwXAn7G5Cje/lSDgR6h/p0EUfar0k6MLOFlWQNIlrYM0ZwEVNJAjkLhmAaBg2jUa
AvoHC8LB+wzzToLZcIrHrZUiKK7iY6AhGdVSk4RHkP7TV21flAL+aN5x5u5LAPnc6zD3uJ8QMUFU
7vI/q45x2Bnrz78PxL90j+RUqoKoj/ogHtYDtttovPEFC8Lw5nGbONgjh+bxYo51Q711+9BH5xz9
GYXu6wy0HEi1RvxIX0MeUS//ENltdyn1IeFGwNfYx08RGfQdQt6xiJPIiwWAneo22E3cjGE53JwY
34buXEbTJCD/CNkb9gQzq5LAPud6tWHhsrbiNT5FIGmu7lCnXLZgQVZHHAgWDdL0GpqH7EXoEYJs
PhS0xDKIj1KnXZIzm6fbc1B5w7vMoodrnPddIOGXphvGOIqIXxfl8iDJU6iw99fgeHEBQ4CJT9Sq
mfcQPEIY8Vk/QEASyRu+l7H3d0r90mtJBgahzX7nF7qH66vZplwMfuKIW7KnvwCZDtgdmjRF/0Gz
HGJQLaUSQO1SF6kZpk5MdqGgymsqd8T4h2AQkDvi0MNWpdSgm2J6sp8IkhqtuxoAprDx+pHhr+7s
zPi756Yq3KYP8mCViezG8TwZHoPgHCAY/1/wqFd1dJvR+KDAUY9Q+la6fCLcgJjDp0p2AZ1gKzIG
HkOmbJjwx2vyr29yIft+GHt9eYVdJktDNDyfwmjKYElg5KmIdwJ5TwIx/i4GlnZPNKNOOEdajpiw
Eb5PRp7zK+NA4khs1Ks4FtsqICuEPe+ZIx1Yobfmd2qhHsO5ze0ss06sXwFTCrE5IDhveUW+lEs1
KM83UMv6S1rzaHrDN3MeBf1d7vXyXoH1qK+d/uxQtJLAQqjavY9X8QP2oLRZnHbGGWaY6AMaNtwC
p/F2Ayk0WS0hIcrxl0bHDI2ZhXoJ9JAQrud3MXsG9nt6Fmv+W3kWJBXQMQ03lsZ3eugPA/jSb77Q
w8ZaBVYrHZcq6t87rw54xxcXTVCnT/NswoLKLj0bvrjimsirjt6Cj7oqvhNyTLW2hVX4kd+6Nuun
Y3Mqh8maM1DIKo5jzbnwEwMbkT7s+sou/Klr8EIF+0Jug/GmsmhArLo21k0VgEPjFg4HcRkatdmL
+RaW/jo9HfsIySoF43MevyMNVAvWjNM2euGQEXD4xDv1MAjJd628ycA6r97ewYL+r8/CtCgS/91s
0weL3oVb1p/9XTKsVZfxesbsOU6Rv8CDstHuvxIQ5LVJU3o/mxJifJgvUN/PGtW4JFTsfUbxmF9x
r20xRMoOa5P6QUsr3JFAmF3CA6oJAgcxq5Ms0FOFgltZtGa/5ThfPBFto5y5Fw2EtEuOkU/l97ic
lEdZRencvIwOE6vvu31JmNprRip7gMwjsGj/sJ9RxYJCDtVWrfOtceorlAL1mKKYSprEjNfA6k3W
yvdBRPHSE0IR7r9ZRn54rQ8O4aOpm2IQvOxMcCWewjtvAq0zRG+gFvVT0O4Uf2Z0j5IiMQUChsgQ
VFvzoJ8kwIQ1ehOkOoYfVwc4SFLx9xD2XfKUNp5eYJiFECWAb1KatmL1DHOTDmYNxqnxrgfe5M9t
TNTDd5LfVei42kcNbQEZoosCFU+A/RBTmw3WaKe20G/GYQ1RE+fPsrrfIvuOEu9L+5dekWlSKPX6
7sEseOiaOL7hUgbECNzhtw/DUS473eBksh571N8sxXOxSVEmRpKSwt2m1wi9tMUcRbPUjhj202Oj
onSYaXKYpOJSjLyBoE8/aQF2yr6n2Fj0kn7B+JdxSvv6wImJKkyix/zRj/Ylm6/Evfo1PNELIUd6
Qx0Q2QFt2e91ukoYXzDnmCi+dRvD+q5g/RSbk3JV03dWnJXwMRcdFtD9+6SF/AFmM9g7S25qVutf
TinNGg7xLFtCr9XOYbal2rWf+LTdH9Y/+au9e+HCjVSpW3XVgV4gNjVPxiKY5gfJsN3n76ZLvTvc
GFDxKNsqgrOKwrEAubDnQNF2158ShHEjlrubH4dkdoHLf9sDhBFwa7reKnjkzlRhlfZEObZfBzAX
Zs/MnORRkHv+MtEmuLetLYHdBis9l0cnE4WR6UMUQWz4nsnDIalV8NYhSLaj5zROdr396xM2nzAL
aK9T4NFs6oeElzdaQLjQ0TYPnHyLmf8q1uD6Bbjq6DPuPY1yylcGOmLI9+C35ewNC6kfZPSIWkkg
ImdlFIXVzZGRtc1nbExXKW8lkd3WwkDn935mwpUjvsERxvew1luBa80tD7fXy2WZEQCCxVHcGoQY
OtugIrdfFKfuq9HCqnNupo2UUsKx4oYVmI19rFOKSAIyR6I+L4UF0LOuccE0maj+cTYAQDxYzTQo
T99lTz41W0myF8D66lmpds3D0qNLquJkMpLMS2cMNVy0R3cBPHACUxkvw0AQFkfY5NfoWId73JZw
gpwr9MCntDwl3n3CKLeX2SSlgclz8NoYSpZM79eF+htpT2nNHxeHm6OawcGqzz/bgb8DgwkwJsA2
S91X1x4zYTM/pFfmuiZWyST/0qzJqD6RR2JRFoUatPxbflhxGo16aFQuxHyqGmwYf0xQdSgrMGVw
MwaQOXJxWm2SmX83rylUs+dfDI2wZdxcBzhB0dt25LA4i4LhMhChMzayM+iC3t0hvEcjwm2+A6Je
qlDHL0W8gETk+iVoSPdJHnGIR0oOZzT7UwoaMBfj4GODq+UiQbQnblNZfLAEt8V/HQ5eGuC4xg7d
rCSPavGeWPYTzYV8Jk7jsWDgg3kW3KVAa/C/qrEI3634D+UQeM/QS84FHLn72Mym7IC9A+KczGSD
ihjxeLcz59NgXwiFOW1rSxnUHsUUoFjY5wrqz168cjcCvM5VWdmx7isUu+TFn4xQImmRkJtenh82
t8YSTSRW5VCDecvwjD73PQnlD+ZSYTZGlI+d99DP4+0GeNcJaTFMOzfTpZkFEtKps0Kngg0kPCTx
aE6ECj0X0WZu6gCXgRHzEPi4KnNqqcjhGUmcLLXxWES8NnrX5eFhYuZkczT/zacV/Ak8CY2+2gTm
c6icvktw0l++W9PDIrenmYHZHFRTN5g9UqF3ooL2nF4KuyElRLDv2TaUjjO07csGyItdJiIhljup
YUhoC6uYVu3t4xkB8FNr69YLmPGYLSZKxmavSHbK3yksK5230YPCDUguRbF77SGY+697l2ArHc7n
DuTWs3NKFvEPZD3z80hcMV0LCWVsY5fXDF69uc7NqMVeNCnt34rj7+Tiho1H8tycWgLAffylFCAt
6mOsemFIh7oGhS47ChllSBsIDBHpd1xOlOoyupm/mNllrGn9SigTLdeJ+dF4coYp8j8sW9xuMiH1
f+AizKAhKJgMjQA0ssfjh8baRgAA884ZQN3IUaU5eMi6sDXkCIX3wxZMh8Sf8ZJIrZQRuU5G3yFl
S11Pb04SRjWD0Si0nxupzsRCOWqXlwXBj7hVJjd1ECdmPDfgB1bKgz8os4x5niH+b6Rw2DyEDP3g
No12NMD4rNNm1mdCYknCY97w1qIRYXHknqWA8uUNds9WWNKDDbXLnsVSa9TABlcw85oU53X3/dW2
Q9D2jMA13dz1HhVhS1L8v9ktxmMlYjLnboWwEiZu1mndFs5BIlyu1lrMMAsK7JcmO06pUku00Wa1
xaF19Quro//q7F8j4BO4tE1GTXW1EIxqAn5kxwurhhAv9reR9Tqy+Akz3WmmE9+NzhX3w3PIenzA
jSCWIyNNACsEgNp4Z2XsCe+ju5seHhNMtbZDm4t71CpRu7fjvDJC8Vgk8/H14IzgUekrauBtb7ql
9jcWnOXzRkBSFonEHZT6JdHSO9N6vUEfFaPxspYXztTl5mKQfVliuwNmYYwpgvdgiQvgdnIgqFJn
oXz+leLKmxQqnvQQF5Q3RLH9ajQTNmtFBOaE2oDHwDITNKtVxAnukHNN66lMD9otnk2LgWthGyjI
CAYqEA87kUzXaLUfC5/O+5hqy1Qh3G6EWwUr7k9vufQIvYAtPyNF8gHbY8iuxEaoRgJOi0sQAiZo
9EhpKcWNDO8V+R5eoMglzlMlZOfkFCnP3CeBdj2/ph0JXFX8l3NK3tupbXHVorK9EPf5fX5VkwKH
axNd8uhBk9LdZtxIqRz7Y1SaUEwHfefRxqO/ZaF53nMX2+b9EKAt+WecAPGqLS1/t619V1H0WOnY
STTyZrhXXbNMSUbMjlEgzTiPaW5LygpuzB7QnFos9LtsrIapqhnwCJOp0hAMwYZGvlQcwQ6LNAA1
UhsuR+7sFsZFBU3VItmZK5m6rYeRB3XTBUgrMTICM8HT3v8zIJabqAqX9JVktDhy+C4s6B+tEZ/8
EHw3sAeWf/kjAmz7XjlljygjklxxTWMdIjNb+b6/V6aE+b9UOaetyPA1JIjxSSXfUUkAGccsF6kY
hTHjY106OYVLEN1YyGjqe+h0Xg33cUtvZl2xUnk4u3O4FZuDo7z4ihYGXlh6rduXKUnifaJlQMdW
EUQQZiBklXBKrdEn4Lpumchn7zDv93s+WSKTlVvSBjEgvPwaNFDVUuAlhGrO7jmay5WQuSCxbYzo
8yGGxfENV8kn2BtdmZKniGA0NWnb1E3Ng68aYF/er9HsOHNFFRsuKlDaC5/2kH2DZ2qRAsZQ83Jm
TR+SgpfI5jeF40YHVFX06S0wlEBjadHkActDE+CI8OmCn6up0aJ3fRL5SWJxKCmzXWWGUEIB6guC
HkOo+TqH/P0fF/71ByWHV2HHQBp5Fy/EmymspdI5l+z2jROVZ/MsQBT3+8J7JgioPqoKLnwUOZnN
2RbFxA7OY2S3E6DxNPaiy0EofHgmzRqXJK/MgFDh7WL5Q0QJ/kHR1xdRiidUi7oq7Y8oraHjTMCf
TiQAJScungpWdJjhdSnGEAeYh9ZimCFLmnYVF27EjmQlbvzXtJ8H+dbMRJ5YWyUe5NQtyEDTGnPp
8P7NiXTW3ZO+170MdyGGKb6SNTp4eikn5Yq4b0Nl0HT/mRJ0LuDNIlgS07+XGXBpgcXJ0gDCllpe
0mWCzl8L7SHz7leAmdb4eayPr5utVqUxqW0QO3FWEn4v6C1+z04qzalby5Kd00a8LJ3AK47yb5zW
oSuL73PLhSbJwI/wLtuKqlYMJxBvlQK/Fpl9Wt/0KhfYAMVM/HW72ZPCI1TGhEFWRKswCvoF7CaH
RC10rOzGHd8iMCWkSrdLa8nQDj/OHBteVPhNwXVqApcktLq5RRli6O6a6wXypX3GwxQW3ISP/aTW
3Yx2NyEvaJDX1Km4ry+zv6fECm2FeHDPuxP2HsJDCW0M4aptH1K5wnOjQnuRswXH73cB04hycFtn
aKiNTS8RPYuN+LNO/VTxo1hfNiTLyd7MWtEGhHilg3WwakmL75/7xttWXpHGCdHcNef9zfxht2ds
dAVq+b1FftOGc8NZaA5pXlFofeg/zbkUPujPiztFXRA6IaPcKyGCuaM4bnEF2H1guYkf/zEDdrc2
ZpPcC4syc/PScalr0AW4dRQqbCtBjVBjeP+UEDPQXvZYbzKCRvV3qNyH431Qa/5IvP0hI9UA8G2I
Kiw724j2kbkHwUDaxBEPKX4zd9mnH99AQWHvk7KklpdweFZ/tncK9LRPTrTxRDmKnBU3kaoOQRvf
69MCR0v1KwJoy8jKQ3C1rL9VmUEegtQ1sIT2MpprXJd3aXrD9YX67qTTUz+IXhpdnmxymRPYc+Ud
Ow8IXpHHNzsQs9d068Fjw6cjvKKlSePwp1fAbRGmPNHYUkyrGfypo680mkvw4yIGCbyMHJ5Qa0Kt
fMgtpZ16dMcTYQFJk5+8aGzd2BfcKET+hpgh2p92dVF8od6viG6F214qJgOjiYZAp3KuzgkZJcXR
9Hdecth397v5orflp3EuEVNLHBHDGfdMfkAfpwRqg4SMca+RJMRlZesrbHesq/7pasX1+PyzGLqX
Tcs6/yOnxu2p8WGw2Jajwd/642hYkZR//JEFdsYJWQ/FS2cBvuji+qpHwFJTsxs50DaLZUTUtplR
bo+YQzlW4EZlaEFLbc0pQJ2WfHhBCfhU/uWu+VfH6Ee2zZsEx3u9UOllDYAm4/BJx4mVL0KHca0O
7imiiAqrLvYbxXNgvgEYqrP4yvAJUwh9pUHZfSHF1dcxA8C8TNDVeH7Z7wfg/DzjGiu3rhLe2K8O
lsHD9xSij6ykuhb4YXWpsPAEG+mOLNoLyUJsJx/LcYdFA1Jr53qzZauexthQHqTFykAp0sckpMlz
p9ldvHCpHQ32IKPu09gQDvb2whaHHCYjDwvY0apf7WeFUBUPQMfhzUe4ALvIwMOjYxr4NoX/54uU
ttwvIySH9Ka4rtB5iggolb8EMq6bc1yYsfDBY9T3VxDSF3SmKoqyc6ubepoDxCK8BjtTi9SI/v9y
G+yxZ+bmrMcX1DrQSBnH54ZWaZOKr8hCRXoRkrdvCzgmv4AegAJtdyHUYjsIljHCJ5jQzCsYJDUF
7uiz8muAXhHH6JAAi9C0QCOfuEjxOhOpeqlb6w5w+kDnWkgWu100wxryoUmtymzedj88yJgjO6gi
DgpfzAjCuQWrXOXp41Sz6KibSvIP7KJF/lMdAWaGb0k3IZ527uJYQE+WPTui/iyjCZL6hQqv5Ja3
o79OZJcX7FsJ6Wgat08ijJ3vpbGlHeOs7OmAK1yaf58msQEx/dbbtOrHrjpQT08A+L1Bn/dnmI+9
ShMR9KAqEgFxfwifra3xIb/gSdU1RP3S6sDqhWEVxf0Uk707FL0Hy05CQwHNvxme3G4n3dh9o+s6
B4bNOxPWQ/iwkaTar2iRUpsksn2sz50vhFb8AwNRtkaLskejIk0E9d0DxCOEbOOXz+LT1ZLhhZjB
Yo7IWIGShQwPEGDdCN2j4QAbsvZW4hsJ+fYHBhNFodAJFZGJxszYaBK5UUP+16ifsM77FcLbY2ax
UBIMirWRc4X/6v2Aev85p7RKdsrwRszkYfHOfqMC/iid+e5iKUxgQoPSjVwdQ6O2hPahi0HcPbck
WVquKQmh9LWhvyyq6BNVQt2ZH/FuaTd3wuMCcYlwAX3jj4lPeZqOZTp7Iv0NpAZQr25jaGlBZ6Av
SqUgHwtAuleAoOiZSgzhK931ye0/vEj3raJpumrokqIO/6VXgmvuEZveBL9Miw/kbYl5XqceYVr/
dgJL60ImKXRQNXa0lEUndxz3WdE29jAwidOIY2AJ6h0CTdOB8Vlplj17KiUFu/k+4lwSAzhDOJYP
esOsoSMCVw8amxn5JqddLFQLtYRCAXHSbnvsTaVaKS7AQFmhKrzglXRA+Z9+W+qyTJTYvcKNBj2F
i24wEviVkwp7uW3mpsNOUrt5fijAOn6hK4w18LSWBszWCsMSz/JS4GNoJyfCKGvMcoa9yCBcFewJ
8uaX2n+WRh6VvJE0i7iTJ5dYKpFAVpXuHAO66ZJUIskvC5eV5/U3joBnFyWViRkbScK11v5qgXSv
AxMMhrfpNs9lDxBcNfB2pd77n060sBCGFiRXv63PoJfZb3ETTYOpCQdXa4motsLl5fvtZXs5wBYp
KUz09S9/7ctI2SeNllTxkcFjYAC8KFXAQ0Nrh93AMvXct5zeoY1VQ9kZDtg3aHPb0wGKg2910euO
PZGqXXVOtq+PaAbmjfm8lJtouymA5+cRLxIMXENQRGV5DIVRp22g5jAeo0n5p6GPNWARwOEoWF4r
7Qp3FYFyx37l9aJ6OAsG9QlY1xdnUoj4oe3Uikb30JRmwcpUtFkpc8xMCS/nviVDxzjYxcF2OnO/
sPk/PIBE3PApQO2oLgUMMIm4c3SgERQpK0Gdoia417PAqy/45+QT2uKq0tRnDtJoSFlMa+S1GOGe
h3ARjPYO5t/rUUYxAtOxMCx4RO3EbwpFfdDkOaf9jcERAyc4v1IsRLWka/xp9SSesHABnnNqSAkF
HZaGws6d8eA3zEWLoFGbAeeJrYgx7Lma4U08UwwB7QJVU9Wy0UkX72dAFP4VGqH0W2AvKsZ8ArNv
oj8WOaaJOooxfcMTUNcAYxojbGjY/ulzPgYU6MzxxhBmwX4QOPNo35XYrapHr/0fk2b22gYtT62A
G9kF1eKRoNHyAKPOV3YG3Sj2dfMVn7qWodfBHRKERQZ4s2BdAfuZa4WNyIBMsjiA9KYji1DPChZi
Ub98AmrJriUCmWJiRNDRbKnTp1J5EgbF3nC0hcCha33ZtDJNKAaMJFMlrKsaXht2vxiIgW/qx6Pj
XQdHz9tZZPg2YCAFFnfdj+dNMsvyVDW8Nx6KkYKtbfzJ4K+t2KNcpyi8rlM5noZd2CqZks/wfg59
DCdif8vXN4aEBP4gJdeK591smDhE+Dn8e/ztVSa7ERwso9OfdGd5N9CAqm7FNwPngb5kv+e67pHu
ggl9oyiFErygkQNh9pPn9Hgad59VpCOO3QVkXzUfhJfdbzxILozGhEiBuVYY9JEfO6mnHy//iADG
b1rPeyQkuz21sHe1cxi+Ru86zJxptb3c28ssXKdgwNWcWo9LNoOylwe1rFRORGFSZSRSim6g/Nsb
K99GnSGJ0wdNlUccoD7/nToYtoavp6ugBFNmMVCVxFLMsEhO5szRYgXMYqiMpXOW1CJo5XZ37VxG
e46KZO25ol9uh1+21PmxhYJg0dV1JB+yojWbwixDB5L4hEe5+NhhEagMrGLxCPZFIF/19OmhgSIi
fKp+TUC44O7RZCsRxrTMwvi9oFyEsNh+TC1YHGj5SnGB4vAptG6KwYXn4W5vvP3BVwJRUnHko/oy
InDsWjN8G8k/2ldA0bm/BqzFoCFvBM9B39f/bhEfkAqtBJQLTHmh2qHuFC1JLJKyqGOstXw9XyIk
F8Z+HOEWHaw1KoKIkn/o0Y2LgzvD4ebsLWeTV7LeDjO3q3tNCnRidlZZiGeIoMwS663nXgipy4mA
Qg61/Sqc7e8i1DHBdnY58hVTvCZtjTvWATHO5Q+/QGb4nKl6Q4GJMO7fuCb4gAihrebrhAl2Vs/W
4sH7HJnE4xMEhSaCMdMhR/dexAsjjw9j3m+ixL7tHIMs3OAPoK0DbLMukJ7p/yKHn3diCNPEd4n2
+Hl3UdfNrd2W88wQ5TWy/6uNZtp1Ce7EBFFuuT13/M0/5VoEp+a4dMl9uApsegmvalfeb4UjV5zm
OLidAQf62hqFd7gUAdkULBuhaRVYIo8sZGa0AA6gpSyBlxgD196I2k/lw59s26bbjtb2/oFZntAv
cKHx7SUp0DpYSnfh+VRpSB37rYctYpvF6FBPA2h66MJslLO+PqAxNto9qZdvnR0YT/gF42aFxvIl
7gxuRxN0hWRkgV4T2K5Fg6R1sEEpHerodejk1szYjhAI+Z48aOohPgBe5kTyfaed9YihZEg0UcQ1
Y1q37d3p6ChKFQzjThoiiHMTlbhJLvBDla4rB8gijQQre6ik1/ufXplYKB2MmOyB/aelWRIduGLf
VWbDKU226QtWoWIE8Ns8NBjUf/JZux4HxE8BnIJshVf5CogtojXkwvQBsDghJs9cUnX31TaLHe7l
2NwTFwRP3ySZpeSkjPElX5EXvEtWdwnCUygeD2/R8og/TnSEJWcn/CmqAI7RDKGyDOnWJK6bUXz0
nZRdL/CC/LzrUfsCshQq3kZft+Q7NYr4DY+Tg5GZjmsWnxrOt6OYdAxJu+tJlEgZ7tkxJPsJehsG
aoZFFiniD2V4+iTYOjH1kH8gb4PrVVwk+eNT1PWCVVJ8jId4j4Ldvs46JGqMxx4vMsijoO3zAKsB
DFhLuPXGDYHHts105zCToSsjJgLJ3aGlQE20xKI9jdVLH8vP9/RRa9T6WTuwfR/vPiuyqXaoIjoQ
Doq3JhFy1d0rfM9v
`protect end_protected
