`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6256)
`protect data_block
JE0Kb7NyC1BoeeVzbEW0uG/toodBNpo5972VYf2kzJ/Dra0/T69FARS1WwGywxF2Hap6lSjC0fMD
k3KrvjhnYWneovajGagei0dOVN36EXcgHSc8QcfXb7QpaVKbyBVtyL7sa1raDTYtX4RdgPWI3AEH
0enfugjnSYR8imac1cWcVKT/Jprgaxnja5iBM+06jM6rLxUcQNAe5kbxX6fScYY+CmQ1ZiYW3jqo
iWTwszK2QAFik1RIu6VVBc3i4F9pn4j5ds6AKkuoZcFqIyyHWYy2yzsoumG2Bgi84FaeHpFL/DCJ
wDeb+utNHb7cTaAgx7N96k+EmGZbH/YUJHgkd+YVjMdCkWhEaxzd/Zx49vjYRtQEZMCEJTGo4idG
YBd+jYrTCV6nST5csSUNRm1KPXgmT4znXQwfIJPHbDf5mGLDAhOQo/wdAs+bNHRzYERBG6jocq0R
3i7TyqhCdwT31MYpm+lHTakLj73KERWmHtX93kJo53vClhSOq+k1SgjnK81Lqvh/CoU7ANwMPVZQ
NsEwrcZotWIozqj1XTTgU3IfnIal1LEDJ7t+1cy4HXNyv2Y6ru/7XD2R2clvP0f9K6l8EAB+Dmqu
FrFE/XtHLMZlgA0HpxkAzokQXyb2piJCjv6Y5qE74c5Eb9mJEHdTjTpR46AulkIm46hm8NBiEXM+
S0pP2pgIc3DHwpOPyytC/t3yekYXKmR3/Mvb/th7y3oQVd+Zqwc7s3PUnXF3ceaFsbOOW6Yry9l9
AabmR4uRTTEUtRGB42t6OD80TIWQOmvUuoYYm0xsLyHOAmIrXHn6oUfO1ADjjliYb/3lLDqKHx4t
DEh0urbmPGm5G8L6qv7/1CpMRQHjlNqJJIh4Wqo34Y6sToZnNUJj2keDG2rQvjeMWxxjgHAN1PAs
T/3FbC+ppVcdObV/Z5xx2Bg1STh92pFDcvJKrzccXXlaJpoe1Ux02vOGiclOajPJt4Clt7g7gCsR
JLe8eOJXMpR1YWB2MgTB6HKnm4Ne8jAo1/rYfMrdiNrgdmR1tosaOU5ggwHgMzkOJiJHDtZvWDUC
McdnNh6kpcKuubU/ZgKJnapLIqMEXASKdiq0cA77sPL2ldC4s68R/8J8QBvRSTpqzL+PLUMlhFux
i/dK3pn56BcScR5y72dlJmScVtayT76D/PhBCmvNk1IhZPHShqCpGdeCyCAKa/waZt7f870jY7if
79lNUeLx1pFzyYwrFCqCadBnLAq9H0MFGq9UyGBTvctz4iDiX6fS8qYPTU/GvmxvJsjpDruq1Z8s
+OTTrLeTldV6tIhJxaMKM4YqZOnJoOjVlYbum3CXJWgBt2WNm7i6ZeWQSSUzIqsMFYp6zK11BbGL
5BflHwJpsEN//Zly+On3XL8U+fJd7mrgpb8iBHy5Z4bpIG04RPD/m+/eVEg1Xyknezm18tjrSKEB
sD/XkLcvz8Hymq2mCe0//B/GfVq8xGVBqz9zT13Yidh20eF3bi3yCCGRwwkXxUCu2ThszdaF8PNw
B2fXRJxYi1133ia1opfWp4n37V8yIdfnb8FiMuULdN+tq+eVgjlxu5TCkDe+cItE/QmLpfaFVuuE
EqW9+g7aTu7dzQlvlSj58AZ73aVk1fBLDcEn/5jHuhRBVOx+7L8BiqIKaoIBmOatB99Ocmz01JQ0
mPGt8TfSVwljbHgZFi7dXw9FI84BZcj7VB4Sm9wdWcEcvglRP5MiCFAJeCpMktRB/MAE7deXIQyq
Z2sLKchoByxqHUIcLMk3efmSyrbBj6YrLxJEIuyKMGK4kJYPQCNlddCvKlf3jVdInNdJ5W2ei0/H
oWoIsqIGvy8loNoVVHJo+52O/JPg354E3vCC62uY2DsT/eydVJPslWPlYnomOWZLO2mo35ysbLhC
COwrTI+Ge2fCUE5w9jrgzUAUOO1Zvzt/rhoMubFroW0iGAxc+1dOBfNDUv3iqIw9wDj9XFXK2Gz2
qD9j8PgoqNToGcecGqwGC0/ng5L4IaKCUk754guzc9Onno/+FRsl99/ic8hScRpygV0siJLLlZnm
d7rfj/Tqkp0pysydK2YCHGo1noS0/tv+uS/VnXUaWDy7Doyh8P6coqNtH+lSUsFHXTtJrvXYOS0E
1e/SUNTFUH0kF12rB2Z++aLIaZJ3z4+7dsbJ3zz3zlKPAYnC1UpzLqzG42JwNj7h0aVdIziT8ZU0
fZbo+Kg1gWgAa9KK26WXjtaxkbMUQxEVXBJJsyQh6PHbnzlx6wGRH5DvA8uwPo5c12mKJbwGq1l5
HhOiXKGsKK5niMtmL5qo+GQ09BjStleDbVVoeSLWBSco4CIbqbFRY2AaIW4s/HZwiSrcT937ybOD
cv9igTbHxJ1vBtXGDRsOjkyzhPUksDE5I6y7P/ulUDC/Jbrvq03OmLmPqcxBV6ZbZERgmU8RM9MS
ADvE+ldpXsaJ11Y4nBZ0Jx5UtWMZwCyHMQgzv4PXEDV8/yn95QaO0Qi6Yissl+HDuo4mqcmJoHx4
7JhVW3ppthE2mGagm7sXdeI9R2eIlkO1s4cTh2Admz/RV8EaUYzy7/13weELog1FhiEOopdzJVlm
hmfq8sNJv//tkmHYQ6t6kJREcA00s2PSr4ugtqcYD8sKK2RWU4HFl7xKkWPhg7QUtsmC1g83Skwe
ULy171F/RPBpVdhzZuP40PcOjOEH8LKPZySCoqc2M6S4uSJefpUPd843TeiH2L+5Fqo44iPgPBFH
IH31u12SqFo98lQA50ytEtYejhGpMMP5vT2tzLWruyC+YbQPlYz6OAUR2MbS9rVDocgrJBoWzUJw
BG4DVn69R9W76PmQ0dpsew4PoQQ9kkX9kh0odTn+vFEK8OnhWN4FjhO0PRUUseEjsOygX/hgnRAO
NdiseIyarGNehTggo5J9NA63FROqZt1/Rs4m6pEcDYDbKGEVGe2ds8APP8OK/TcyzHovPP1Rei8O
F/nG01NhgVYQbPkAAkJW/QNFRtmJDQihPkna5YTjrvWHEeKt3i5pJHdAzylBRy12xPhEhtzLBa36
tpId9ub1vD0b1xzWE1MLZURsBEwHeD93bNkF6hFI7SQd6VUuH6Zaf9uu9PnnTlzfdOgKFSrWMSRc
CYKOvb0vWgriPSqRGLQksMY/emeaUfspBp1L9we2ZY/JqODfStntT0Bz/R24ZcDkRmrCmh71s5d2
XWqqqoWHgc4obftIQl+cEXynh+AjPmj2EB30L5sdKpEXU3nGC9y6Fl6dyRxozP9Xz9ITGbTVzcAA
QGDZ4mq7N1+RQDyOS+DAQOM4BgexOk9oxvpZsKkWiGOMM3HQ2IoDaV+z7IpztkuLEOv+UJgYW9tU
iRv8gzfEZWv/eNWaSnsoUVkda4WNYo6/WooOSpcDzu8YLoAvjLU4dUl4gM+e2TRIqTNx18mPe9q5
zmVbV5nAsHJY8J4aV+f0sdyjDLA+lFgNgFOMm6Miic60/yNsDt2IgltQDibk693B/4JoKInazef+
gITrZAOUdT7+wiCXXDqCRjbH9UjZZT3yY6GQ9fEzZrHSibYem+fJXT1WYt4W1OBhd3q2V0xnRo2z
IvIqp8y8EiBiEpz+l/kX2BkINLZKEnMm98Hk1SFBayd1GlyqqRw+x4+dXQuSWaeJnQVP2ITw3Xi7
u+TPF3hQ7WoENyNbKeKtkn9gdahjQsKyX755ZVxFLeG6QqQ2n0MFJtYe7wHllkiRL1mqTd81O2uF
8v1HngnsrLUr5zqIMVxPT1ESx7DjzU5rhx1RuPkf5k4HKxgNv0/Chrkb0Ne74Tb1TTwLj9URMpvs
dPtdZj6uRo9BJ/zXkRIFTODoWVRVbSxagT9ClEnuvS6u9pSLrTdmHmCckbdz4ssnUOlpCcrVAT+/
jUeWxdldFb6v7huvIr7T040fwy72Idrj4bd8yn/z20bJeDvVNT/O+b2UIjKIDqs8K4AIAQtZWfo/
zcUwT/DWRaYxisjhXtAfLOFOku0s24pL5/oAg0kMcBaQ36cBRBOcGmeHbfTPW8PPmTP36vAP+xQ0
/YEyEafUuFZdiuEprGw/q/7yWpWvV1rdECGaEFvKyalrnJmAmM2qt0YqcOfZfhQ2uCmTuBCFkQDS
HmIr/x3+941HDrNMLsgNtz7S3gsGOqoIjtPH6r6EIPg6G62KAlrlWgunkuuzeuhbpTg8Cv1k3GaR
i9yyE26+vrXlHLJWWQKn1ktqBr8JNb67MDCjDECnG2RL33PkiF82mSi58mqgQ89oVw4+ZTIKAyn7
6MXJoxa4bM0M9v3BgCUbkiTab2TWBM0ORiePqdpYxw9qmqKMR2kxiRbEPajnBihOrSwgmRqczHmj
B4ETC1x+wjiOn1X5fVjL2V9whNeepCGVH8LsC5qm4/Ar2+eGzjMcbdrfR54ElznPWn6oaevnuPfQ
xhts9LivfGqVioic5VSLeW8EpdwCsgUYEpZNW5g5zu3kWfzS+usVbhK1QK9X5wUUoSRob3xT792w
veNjCwhR/0Xc8W0tZq/AolI5Tyg0lD1RcSE92tthXS24vvDCZWw+ylJLoJUXV9URc8bcr4S3WQh2
ZP/6k7DI9ow6jIUDb4+ClvN5TjgcGmFhHzDeHgl3w22PSDiYj5m/6xoUV+Sfw8Dsj9rMiYgQ0nRk
1z50ptr2YiMTZbgNTmb4xPZhG7R6l0e2OMDVUHXf9whfxAzXw+PHv/oPXOVcINOh1kXxSDcgVlYn
0mhb/pJI0RF537gqArl1ch0urNm4wsLiA2NZuupXr1u37L4ukKejQ+G50Uj/Usdayh6MIhZj6tT7
9icIaPrqOcBYkt405OLoAJwUQ1Hv0FyabhNNpIVS8KELBmIV/jY5UI1Z/TrpYWhsVYVZ0f9jk279
IEfJEwBX6yAMgprgC0colX7z0MHCfBCPPBS+TBqhRBRigpraoFjyVUYNM01DrpXzm2ReACj1CQ84
nx1lY5gQn+TYhRorv7X9EHABA5tpDXFtIcPX5kyVu7wolQ0w+x1Zuo/fVxyzTTCJP1jPCrbLAo1o
i7rl7cR9k7e7NNOmgrMY0SuWdN7cwJnVh+uWURwdwd4vPplmZYyTBqBvz8QHwVckt54LrrFUJqpD
WyNVazv9wah9d38Xup3Si0IOslQljVbI9vhDxLYSxJTtMMS/34P2So8PHVmBcx2/mEJCGpF46J/F
REOCmEUWptp1471RK+QxZQ/Wabh/o6RzLyI3JBfc18hLLhaDFLaZpL+rXJMjKOd8u4DN5u5FcEON
ztb2wPHWvzb4qxDn3Jwl/OL0yMDZzOcEYw/axAJJdAHNGjf0bkPlgdIAQnLyh54ACIBMuvun/pRX
hPtLoA1EX1rvLBTkPLji0FldjFLE6z2UuR2Qpg57D3XyFu5rGAOA1tea9EFOkA3MP+A8RTgW2GUe
k5igh/wO0leLYnehe7RuCkSJnotQtpFUFmO2wMsNl6eA+kgIsZd2CaoRq4WbwSRKejzzjyOqi6kH
ULnfFjLlNBR9cvVBaIfF2zth5ej5r/czFzW1E5ietB4RS/cDRv/z0pjg4kUeDqrNOyfBaV4+Oz4r
HrLbkaDZQ2xbXaMMPjYpaopyNcaLBXo+AMFUawevmfcGovtBmCJbvavjtIrwGrRXNBL8XA5v3Zuz
aFUgWqONfgQT2JYWXDd2zZ/SoPnj2baWnees1PLjXVqkFd8tEKyb9WwdrfzdL5rpzJYMs/xfAoOg
RfDRQyNHtIjKMoyWjt0L9syVWjHj+7Z2jQtZuUVkbNZl3WczqDVB5qPjX2rTk3zzhB2hnLorkBRW
D82GYNyzmgMswGW+Sg4EHfigP46yIhkFRLZ5aj59aTFgo7zVbEw3eMj/EplAcB2IT2amRx60sDkg
JraEr3F8N/PS7USs9RQ+/CPhidtjrMc6kDuThfNEXrf1XteKJ83C+9ESxsvEB5bQafd0JnORt1r7
00Qa0OrUo40d5jNEL0+qElcCsDez0e7GSpCMBUEZ2weY8eJ3JfHfQlKFNWOEsl5UCW7/Ruhwembp
ssGwY7OqL39qe4ErqJbg8ArxrSUJdrWCeC65m236dcD0DgnUoPuy6W2WhW+dh3XJ3fZrT9fnfcg7
/dsO/qgGKecc3vmABVCp4Etb1H+wooA5o0nevOrsmBHNAPkRWHehUIRGEoLuRZP5uRuRtCCkqVui
HRoyA0v2zOtI7kWUGXd8o70pxf2Vp4XwQVUNbjsZZsbT4BXIX2Hta/G9OD22whudWbAyZ0ucI+Ug
YIRMUqcnAfXhy8FBdclBG5MSTXb3323AICnYyPVkPXAsufpM+gj9XR4OiYBUj4eujYMv/GmSWUCP
7vgn12yxFxQvxTO6XQ49C1oEgne/XeiSzkbyWgK4BsgO9WONFG71hPOfSACsrjcI4H6CLRshPwRX
NaaQXHkqti/PflxepG9mv/kL+Lu23Q9pyhpBnuS4UUGcFKSc3/NOv5uwhD/BPU4ir4VKFf0hHxh/
qAU+t34MaBlUXivGKRjlbTVFJmiRDyo1zCoPGHiTKAYoP7gBZqYMwkbqgcczkJOhnqRqoF3Wk0NS
IOGggxkN2xyJKqZjo2EbFdv3Y3Ne3iw487EqBwiVh82+jWY5/Fr9EQJ/vN5NyYONg/71byVYBUUl
gaLdQf85+6MJaaCT2hs9HGTw+1QcEpeTwxcINlnXEV9SH1Xfwrf2DAmhGaR9cJ1Z1zyWnqiv8bW3
zshHIW2qYJ8r2FKHh4AkeYRuM8i6uAZ7HCppJGCNqweZKesxfem+TVX94QmmLZMpe14ffV8K79gV
dXIBdA3plJmF6MYYVPFlu0j5j/w9CIBM4aqlKtt06HaBKGrQI3RldKSDq9UzyV/AQTaxiGp19Hyc
OceYpK9c16M0zQ6CTMwxfA7pm9TzTTQsenlo3ZCyXlocBLRaN72bkyeAwGwDMg5YjDV+o7o2IxPt
qTV6GSPy6yvGMDFr+BfMZuA57RnqCJ8e5PAOsPxcQ5EAwX18WUto3G09QbRkYUCoDm7tZn6b+69U
IIn/cTS2u45R1U1dRkSb9o+Bs2KyubvoWE/OFE302Y2h3DHr81vZfeYq6VA6R9YRgMbu95RPrM1p
C6hlGaFJZIC6AD7oy2O2w1SOAFsYnNOsLyAwmuL7DBwiVbOpb7djpl/WAnP/lGNXzjreynKchKBx
0IjBPMJSYnFsFF9l1ECSs4p0IQDu4xefXHoTy3cLYoL1MvWNld5SX9EemgJxx9GsJTKe6GoBAnXG
5orjeJRvsoG1PP+UbHewY/2uVcCfFU6tkM3rY0KL2OGqXqUOuOlyheRgRWGeQlupDsWOZiSosnlj
caNU4WPu7iqoZPimVLdXKeqOGTEs833er3RPsNaxLH+2CY97mci6juLccOC9BqAPIBfkHE4OFAb/
uq2nsYM6S23lTpkEfsnH6rE84HaIEwu5ZEphWXxgdIeSjhLK6yhJphNl9Bq+YZezP6p5hC5b2xTp
kg4n5+MJNwBSQeW2s5eypmxt1HpIuEXDVg8g0N1TFZlq4f0qCvuf7RA8kJUB+PyZ5K4CCTPu5Ubu
4cx6B0OUiyZ23ygOEWba6zqmXsD+XwgTZKcDQBSjg3jO3Wkyakbcq2iArpuPxUD0Bcdl/HPwerBE
sDtHRq530Qnwq1btTnM6LfCHeKaHhe9V2wXjfxinCesalcBh2oPdCkwrL+T5sow3V5l/lNIkQUHK
I0iwLKpaqtLM54lze6RXfgcBjiN5jWI9ffLulyXbUAGleo+4xqNwdhPYAMW3JxrMWiuslLscFnE8
6b1FaohZmgWaLDUHpzPd8ZwCK0uYqMIo6K0YlO8oPq/pTkaReA2Fy7lFygRC+bPtwKUh9bnJZRAN
iC0z+vrP4hnduuFbKM6a1MIGSpd2wk2egA1S/dsyEct6e7z9fcBB5BlwmByEoHWi0vlD1LqJHC8t
uiqWvLCZ0yv15Tcswvg4jRtUwft+1aq0jBtqbT3ylqnHpqn2meXfjtshE6S4IIP4LO3mrvsL2CpL
ppiy+jO0h5BBcDzI3BXTouQBSBHgEYCQXxXnvI8EuZHUsdb/UC9KbbJy0HCnYRv0VbRSjSTsOjSq
fY2GNpNG79CoL6+G43A2I4BjFI6AjQznngxCCBn6rK6pYhfH5D5brZSaE+3SX8ApHrI6eHhdT0Js
uN20WAoTGsB9p/p1tfOt8xDDNRiDd8ZX4nZaPoHGsHJ+ib6IHskgJ2z2BQr3ntiwVf0fZcB4wH4W
F1zr5++VzMM08nLpLgtMzyKQqvZFg0Xp46vBc0MlMOUUhIBfwcaMZOmhjPFd7JFYs1JrCkU6d+y/
GYFRlumly3fsMn0TvvZMt0YXsDFP1PrU7lJkuBE4CrgcqbdeOSrbhQQdWQ==
`protect end_protected
