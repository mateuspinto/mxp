`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
sje1Qd3NIDtl1AGNZY2um7tsxRmKhzkZmOtfVK3RceQNPLo+oEpkhMb5eJ/XEFHbpr22ZVdysMQ/
32Rjuh1Xqw7ScevovoNG/qScNbkYu8vDlWifyBZFlNZBQZ+BB3TwKfcm1T6rbEI3ht2qGwaYX1hI
XpT2Mkd1QA8E+1wip/RZuL43WL37uYbHzKVGX397REma2gRpoA5dKZy0bSxf5dT2YmjMyjxP/wqU
1LL5nVJLiFSgixGbKQizNiBHQ05p/P/tqFYTPsdV+sqS0Hk4edGtUh3xjqFFy1vHkmrC1wJlTxwB
YqYdCpm45/8nA4YcPGBVPDccVCfOeJyavq6ufQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="U7E1kuW18QHaYT5F2/wKl7lnppEBl5f9pfUIgqBOi7I="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4384)
`protect data_block
5vu/waqNPnDHSe1hcjQqNQLivXNudbVXrKnYXmTnh10AtrOCWi9VQv5bAI0yWvV+eP3DQClDSM03
+viKMaidKcw+fGLdu3tHRDQXp7RjISVx8kA0vVCQIHQ6aaNzYD7vyVwxFLsfoo0X3kjdds2k55yH
WE8CFJDlIwU6c8FKLS0+niZH5r3wvVkTJNCozpH8CydwN90ZExrwVueqU3eZt2XJJrVLzqIUeQa2
w0fMga24dvAo2M9m4KrjbmUFej4ND+W58SLEUbrp/nimwQ8fFX7u25mCAgjzPQtWuc2raATi/Y6S
PTbEJFY3r6+nUFagHOoSvrZRDGs9N6bLmHZ2+PflHCP/hnESkd/xXEq3llXDxoFL0E2r8ow7X1yW
7jYRMK5uEYUgGAvudvL+xHf3UFtJW4+jyopfQuP/s7T12rAhrFgrdQRJ6fV7m8WEn0p+qfO6Ukrd
In180e7fbDlVkmrLWzu39XLh9L69lEZpcpBWN1aqmR80xYw2B0IDB6ygAhIdvZSsgribqsDPPxyI
SucIQPF+WXTuvk4Rn7ykObsXuqRfkL/jszwkFZgi0k3+kevIjydlJ24tUeYrdLEDcHae0+OMaN8G
Op4mpFV+7JctH5IhgHu9650Tr0jb3zzNntSH3dx4fknfhNrat97eaot0Jrrri1hztAT3LgpOF0Ul
/x3C3puh31XReOgA6HHgNn/tCZcfe9VwJjM1BMDlopapEJmmbqRCJg9z/2m3PZfg9+wxWK4h42jp
WHMJ5rbkXmixTjHrpJ21lMDORO2QVFcXIKjR8g5tt2qlzlkv1XuyWG8PcD1lfWpguR1hxmo+Kz/B
wP0SLpo7CUcqj9bZPpNCNe5rzQt7KbK3zLQq5uDVcovY4KpaFXX0Yq3GsT+uDY9qY40vra8jcEAJ
cDbhFh4/HNT4b6PevhfzBH2o8Cai2ErSsoUG+UkrHX1jy6LNO1ciZqinp70cWwLOugJkk6Pf+5Qj
E4Q0QmzxwyIKUU0PD7ndtABTe9h9RmvXpwxlClni3Y75B4d+ukc2N4G9pSXst5BgPIo9Vn71w9A/
mulIVXp2hHdOgCDT5pWYy9B6eN0BBREFHv+7llNEUBhr5kZf6+9ED3p/W+BO2bLDf1C9vdv6tNFr
q94iZo3lPj4d16Y6XWw3e67tuOp7YsS529dAiQi7lIFnY25ao2EHtyHBOj2oaE3t8xBevN7OwJr0
Emgth6iluEe6gvSRmwm07Z71LSoqO6WpdgsnOYOwmTnOClcUJMrbhDkHkDkIkMJuBDz6w4KRd+KY
61iIwt8sraAt6AJKPgP3JxkfRxv2bweHxkUbJYmAkm4qqieu3MGoAi8Z53934oOGRNReDbfhSHiG
jhqKgqwNsVH7AdJXDvuG0j+ZzOI6P9W/7tjVWKT+IsdJfE0rLZKJXGBiMH0ZTMNQZ/we0i2igDMO
+Jg5FK4C6q9edSSQGAmrD+MyTWU0591K9B3Q1A3QK6+dpn/+OUmHpbTM+blzf8LLSYNWiY1gkreI
UOTRuRa7c7QkvNnYRXVZds1IUfO1A3BhKj9kv8AmMqHOOVDC0gYYU5KzJQrHDPRHsN396HvjP9+1
2I5/E8rEkFjsRg0824ltjKNHB3+ImGereSIWTz4Xl2tj7jLY15qBW4SuucolvfcQt3NcaeCaR1no
YkJzVjzW3c0KlI8O2wxj0Ubv5ie5Bb5N/40XBFJJm1CRoQLvQ3HbRNYmBKRl6Y/qIp4hkYzecM5o
d6nSu7vafFSVDgSUrjhALbP6srvhfGdDwNJCltBXf6Id7beb/iD5IVybK7I814Nafifia+Awe77/
4KANeQij5g36iVPysDTrIAspaoPwHuQI1iVITU+WTiy5I3fNKncqxhwbrA0ffaDyMyeKjxsC4T47
bfI79TSgnWcwCLvBcr7Xsz4UVNjJs7G72g0PhKjoeQjWMQ6BSHOwf5eyn4oE79ISdkrSnY0SiFhg
oyfAl1HF4Sn6O08PcrRI6ptP53qpAbR7ogICFe9aPz6wIPgs2QBsbbwl/GjDfWVx8Kt+R0zbQJQu
073ASGTx6mpkj8c+X8B6Ly/rubGLbkXqDREFFDk86azJm4DOT2xaA4jna3P3bGRPx4j1grco1Jmk
6vOqxkm1oAiye6oeOIw8l3TQ75WVQLFYPHN/kch8wdNdjbyUyFolWhA6rgrWC7QndD84sVsr5Msd
QoJAAh7JQE0y6jARoCd3vXnZWPZh45iRyBtjeGiXWFPpnJGpNDqyNtNj6FykNIzvCPlXeq18kR3G
YybHteKRLjCcOsNEeh2on/d6t6CQsftMisADxmPPYo3tjRwRR+F+Rek8vrcz/lw7Hv30Jhi3bUYu
hgkIXXAkn3gkrNNHVLpsMgFXX9O0iSXO+pa6k9hUd5DPwhZ2J+XkPZjphCr2ZaDWQx6CwZbGhiEB
U8C86NMxmJnJRv1wQnjKcXAi7zxFuE639Z5koEIEEd2PrMSDYEA5JY29LbTU6oBqB1rjvey0rPbS
1swIQH3/3OB2UZ1xYSkDF2KqXESADefatNo3TT0UUrmGacP81xG93tHAjSxg4pWG7HYRnkevhvky
pMosQDoXQoryblErHv7TwPHVt6qMu0bEU8It7HeOkiErHfmILWWea+xBzpXt6YfkffcDQMFu3Oe3
8qkA7NS6VLK60ZwNA9TIHenUKfKkShkD8Bg6TyCrlyEgigyMsu4ZxgPObkGP8LecHFu8fNH3Vc9v
gW9avldJJLlPSTmcYDEzXGHwvTnW6/pfVXU6ElQQgjqF5wvH6X8+4pEHY5cQgOIZjgsQQtwvh7Z3
Nmtc9kB6oYM5p5cKlCi+XpQyX/sn+dbVFicRu5mEj0OJppg9hQqRgGSaxvvWA/EaG/AtALrzOkZg
YIMvP9UteOpbp4qbJBWAYuJPQtMU9xzWaDrK69r3vaouqrzyuxfGpljXUJ7G+ds/G4EDBoP2JkI/
wL7OVry8RIeEw7achTHkYzFbHj3wc5tx0IGHCmFyNLUdgZjZeHX8+E0LJTdcAKP476EmarskFS4i
ZtzZV4eiBnljazO+wlyPSM+A3yEPpUtXMMUBgPNe/VNaf2mAgSCKOjxmjQAi28P1Rv0lwPepWnDt
1UW9KdaLYzx/tdHevoy/BDL8vuj5uAS16PC+rtnxJUg3eePzWkgwgit6xAxisu8d6tq+8VkVp4lQ
06wpO2qWv5k4JeiPNtcABkOsrAU1yTaUObLzLZGuTJZD450ZrT1JYIm/orvXQ6FZuBYR9NTDpcvc
gH5sDwsvPfon/96aT03XOHpeYYh7KhuCVMf0tj0uAH9gpfuBYla39yF01VtHb2wwJri0yfh/lcYV
DnZN5FQzoTBu/OoPTGa197E/v2xo+zjXQUdSnTq4fVrdQpr/ExlLroK8EOVySkPXjxAD7aLQ/jcE
A/wKXePcjtlJ0pOsFypxOKnHdsJU6xzNiJLwcNi+PkfP+oxktEctm5mQyTsZX8b0l746M3g53UlD
lflG1CVdd3AAR65JiWoZh2gZt6LFXxvSoDFbIgfM5o45bfFvPBV4WEOMCLzRI7GqajputRg6Gdmn
GGzUeHVBYbESvMkfg1WsVsfZEh+VxVFGlexuTgoJ1M0qA93L85TlCy6ss4Jqq3U0dMQlREjTLDHG
8IgAYXIRvcBqL1jY/Y6MkFUdIT0ZBsSnahNWmRV06yl4dpPHuATP4LFNfzaBXsUugTQJqtJLSjjG
Eo+GGsM7ElMUAnAeempWZbNhwdRnUBVwyXPaBOwoEMNbfZ71TE45RApzvwtXRhS+/30HXDleCwkN
60Ma6PUDDYzRPtBij1xg2weNbUi3UXtuSjr+p4ASyg990r8syOp9ATEgGU3KjTZQGGmIuGIt5Okg
5fTb9NCNInen4b1AVJ+94vmsOTEtFmI9A7o7UnzDS0Pu3V3F2fPdfBJXw+X4XYQGQ6ryLLmHdSnf
5Df3qlM3AdOsO4+/c17EUZ3th2OzpA/LljtTh0ec/4CeXNyvnN44sUrMhDBkEGpTY7p6O8WRNN3s
vA/Hqz2zinVI7lfGQj4V0cafTDVmhMDn2S/vcFKCMdY6uOJ/klGNBpuLXtS5WN1HvoouU4OkHq4J
Io+L6+hP1sMNh0gyNWw/oqbJ2Oev3EisejA1UlPzhHgTBLrDwj1HGKusAV6kdmpj0EZ7wziZqKJx
mlGilB4H1G5HOufr7o+uFATejr1Re+g+xvv1GXRdRVkfN/fhbvc8X2tF1Yf2oj36QnbxG+qEa1gD
QDAb/KneZGmOqlTHCAohmU348ZdzUDSc6i6vWtgnPSA3B3tkryKx8FxNmc9O+AOOutwzg3DyCMmi
Nj75F0m/UgAAaxcQt2Aj1v/ws9SNK69I7FcDY/YfjRMbmeFgv6Y2tV7bldNGY7KNf784NaUrZAWo
URDK5nSO5tXJ3SenA4lgrY2ElKSFgeubRXUY0GliKwFluStOO+5M+JUVY8aM2/XYvZ7p1OhQ2B/L
vVkKRAlMqkwHb0ITGnkoG18PTMfKCoH9Ol8xLpvhuPaVKbKqaNv2Ck08jH5Efb64CtPA87saX2vT
NqSyFcMXYasUT3VFih5BAHIV3WXzv3FgfstdZD8DFCVxYn63oAoQQbb7lRonMBuwdej9z8AIAaSg
XkRgJ1FY7OPes5f3pUvibILDhjNa8VtyRaYD60FakTAw+vI6XnL0ZQ0gvLHfj6AvVo/zkmiMsiY+
ofwtSU3y0+VlNcZOSByxpw5RcJjYJ3gsckVH6p2yBa8JsnAWC/iDfgeiSiWFdmYJpy6AGEu7lixI
AxILFQMYq5C3afuKFCBdJxZeINLwFIBpnbhekZemCKtUu6FpOQ3kYriV40wGZNYQGgL3fhP2bQcM
zDs1LZxO1P4mXx275ldPwwxEMGhi0oKRzupF0CMZxNz/gMYwsY+QtJDBj2JtzBZzEuvkeZBl1YBl
FxQvadvoc0EQEIEj2Mg2EDXc5eiZlfXYIfirwYL/7Xw/J4QcTLmn3rZTmJBsMyUgdKBXASC5fKMJ
RC/dHTQ42LoGjrjMYI7Av5SPA4wUqIMJrm36iJWEvkCGqmHV6FwlCrqyMg/yEMJTe87YrZG2eZ8+
puLIuIOsEqzu9yQHr7Zt5Exsj86uFBoEUMGk3U2Sxs550yDvKMaEpPVmzKp0M8Yvf0AAp3C8qEOg
bRe197sq6GcRNUWSRibNyeH/f6LtQzK+DPzVPp4PO2BKzGmOygfs4TA1PcJxoYRYRuatzjjz+tXp
6TPymn9qyJ0yuO4OItWOfnSg5RUUrA1XenJsgSnkAEZ6T3pEfcHNuFMoUP6xwAJZ6/4okbTnYbkx
+j+q4soWEqDIcChCPoKsLL0LgsgK7EdXKWPaBc4lkhR8yoZNpKBVjoMqior6Cr/hZW9OePDBh3RM
j92O4ViqhALtO+ZBYJmvpLMhNhXkIVhG0ls7S03LCRMRFT2d7/c6EyWN0PbPnMirwjjPAm8OCAeu
bukhZ804r0f8dE6mw4GaY3+6xcWqB7XXH/TTQi/vt4CcedcUpEGlr4M7T2eIWiK9lTA4IJ8RzYUE
FaiyhnVAh6x4A99gYJRONWDff35FrwaZse0ewzyYp/j5tb2+rnEMbIFnVE+9dGrqgsHlzWVQArKD
1eb+b7aBfLH9MyZb9DWTlhe6sw73WXrEfv8as8rYMHmmXAUCVSWUmShATm8k58MOm9WrstdI4BM4
jbA9Awm9fSrqkD9ntqYFm8c2Q+7zmUDbHdFMJylFIwMQnsXxiDTna1hQ2BqJBk92p97OLWcxuDH2
abLedSxsz9Y9Z5L7sZvNPYFAdKrojNCFvLU8H8qlqzIzTGJL2y/HTnSN9qb16chlrGH5eA==
`protect end_protected
