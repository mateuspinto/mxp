`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 73904)
`protect data_block
9b1LEQ03O9V0GZ0LDoR5QeSJrW+h/+SSGanA+YmX+nQcxCYEcYsmA7nL36KOW++DtDv61aRSQAWc
WRa8YJKtB7+c1YC+0x9yoQpiRLFRcWzxOd22uU7EpV8vRdO8XBq7M4jjlKTuDvz2wnBJjfvqo49i
2jhlcdbxEibb/3lpu+YQgU83tEoWlv9A+WevdbPwP/zebWAomxjhMxRnxJFdk6tRsE8VaIApHH7q
7/fGOzOAurdtGx9b1xRJddpTWaILxlaTLO2z+QHwDV1ug70ZnB95xdcFtV7eCoAArCahVxguuaog
MMCD69aB81UrWL+sjZxQvywIOBq4tSbrEb8oVdhnvvtGAJAPNhihz1+re/0ZoLPEUW0SiP735m/S
IG9nXlFpWUZP+LUOyCXbR0PCP4BNfzN4N4QzWUs07xKjhMwBTl7q8XiQACY+xgvPr0cYryLMlNLb
2FW0aPz2PeuxVgWbQKlQ2wrxpn9wahqxM1vn73/64cvqGPLBPu+0PY9cwDt+ktfiCpUlV6YRk0ZB
8qfnaXMPFAJmmfCvwSBaq7kl7kNEzW561Pt2EIsdzQFcSNEJVQj6E63L57knkhrMXwz1gakgTRxv
NHPPeUtkqoCzj9QpX6UXGAf7sQJmbCXwFqkDrmgjciWsI6Hggf3SrBUs5/lfGCKzpeZgHJ81QvxO
sIKDV17JbEop5BjI6Yc3OqYvGI1fxu+CjY15aKuMDbWnFQJfu/hSi0Upg7TZjx368SAQhefgbZak
YIN/pRRvF31TVyCFbS72gb/axbBVVrLt/8TEntptnxCZfbgw/ki37FGONOAR0FCA48cDcieuqMys
q9fTLcF34whILtS+pv1JP9z9iSsAiJRkTmJ/crEDZ1X3sxkgXerubb2Gcy2Pqmst6mBUVzs3oHTW
iYvY7DkkbJrX6QU/RENxq4uRfEhh0uMMZ5bx+MfnL3DGyf4j2hC4VQsQJvRy41m1KLCgFtg9nA3I
R0G+HvXIioZJzD40zBXyqH8UlfpS867RvjvQJwVIO0pbfm8hWfdTpZ4B+k7uCtokgOmCSkaxTkwn
NZ8Al+SsGW/7bi9OUfpFdzfEgpXkGVy/vxF/K31FK34yONl3U1uaP8NFW3E+WzgvQz/k0q6vzWv3
7B9g+P+XvomJrMN9WjpTr0s1VWM0bouvInFJHmKVjZpDhHhjP7UoSXD6xrz8zdeCA1+CtwcHKZ3J
PtVzP+GU9iOjTl701coZkHL8uSDEsi3zzpAKi8Mlb5M/7dejoWXnrKO5hB22JvCCgKOdwpcCKUN/
gXMKyR2QpcdLOa9Bz+pYLcVR+v6eBdK12eQTf2vyufsr6/OfXD6u0y6vQAel1s2RWu0I0mJHNzKu
tCDP6UVOdkb7aLtSn+0Z/rSh/8tA0BSqPwx4y8yaOeJV16fOvLLmttOKtMPgAEk+rIi42lkYRAzU
pBe9oNEdT0klvCGCWMA6MEzbeoZGGiQs3+RPAVS6ASdW/0idTsRc9H9JDLUBFCSJ8KJk4AD45ZOp
A02Rfo40slYBZ3ISAYJelRLHdAwCzDR078gQPoOxQdGGCeukcMfLY5htDRFtZc758OIF9pa3Vdxj
4VwYBQ8lTZW7mnrAeMXmvMmP8gc/V5EhFM9HvZ0jMyf/z7lGcFZ+P58S16X5dhWYyph+z8G/VHeT
I9Sw9Y+iYjNWURSyP6UBvB3FaL1VS4mlF6WNoIHsQTbwbex8MqCrQiQw//7l/OppUzlw4MZx8PIP
t7noysfrs3dLMaQeA7GwvdI5Zq54jo4xbAtc4CBgc2oNBv95yUY0RGv6o0p5LO5TKFU03oOMarsU
JFUH3+yFvK4smzu0r3dKksKthE+YIfEbYOnScjBi1QCheyRtpYHIITKFrr9yACO9/meta7jhalpE
m0UKkZYJyjY8qI/WyvjHStfiwao2AONRWH1q0He6qBFLUR0TWw+VCCCDsYEZRhG3PHk4QrkvH8jm
x/DQiLA07uBiUs4ewhN/ZrNJXHwBcKIt7x+rDBda/4bBtw44IL/fjX+6C14cLBjQj9ZfzbvjXMrK
6mciemf0ULy3phBUb79A8GMnd27WhBRhKdhkDoliHwdhHFURN8/8G2KRMoHUecC1F78NbkRagIIS
uyvzoVR+AZIe5ovXbvLVf5dLM4D4ULNCFqVdqC62ECeceN1FxHHuVWawxAaC8wxajG4C4yzPHOCX
cSrmXwMhAwwUKcduMjdrEBOngRE5KmH/v+wwL4IN7goLtpkoYol/iKqOzux04cMTapuzBu2cve8S
4MXAV0wxgJc0ATOfIyE1qOE+RIL3HwnEo0eMjHbSy7IYHSBgPeoOor1bhXKZm0UftdJVxhPh6h/D
rMCpcluTGvlLY7+dZSiWNEGxBrsmK7ahOzjEmI6QW140XG7QPFpUzFxvJSOuEX4nbrDAbr3O6Gv4
oHhAzCmZlo37m4DMX1//Kah2r3yLvxUaiTViyfQ0Ll/poXebKTWFAHUG1dTc2Lj9+wt1rG/rMmS1
DoxthbsRaePbI2Eze/I1NcvzNJU7hRvX2ytboBPX7pEmsU1fUeK0s4eXStauedOp2YC9hVSl2Ek2
PM+rR56cvYIR5lqFYiC3oaD6uFqKew3dLYqzG2mZQbCfV2KIBtHINE7dHlutAILwIL5eU+b2Zm6+
RCMQjU/lOH075/wcSrmJ1CruEGU59MPyXtQWgrMM9JcjQizfqOQjMGKCT2ttBI/g/aAV3X4yHqnS
TKk+mMP3rq35P7x/cqovSO/BhIuTnqkkpMUe9njMr5m8lj6rZlMAaCAnDDndgm9vu+8GLdnr28Wd
o7fPtoeyjCKjOq5b3C+/NQQcYLKhlG63badtsFe0hWeKtbgcC3hxpKBWBPicifg2Y5tvhbG8S57D
WNm1HV6Og6scDVcMUAkoFp8KoBUuQPOvJnH8EwOBd8H5pPZcs5Khr6wXE8rWT8pUexWCCjP4URH4
J/LOdusAejMlkQnTPu6d5xpBae9Opy04LSPp4kjBTM8V47EqgN/TZyZ2ACJ1zqRDcavfDdCxqGkE
oxGghCyd3n3rsQEKVqvpdGmgeaRhdGqHDEAL6NjwfrpWREZscXYoXQ8LVOSoJw8HwWNZKiJkghRa
jGF3U+BmEQCm8b8KpGSzbZ++THz3hHTqjrqCW3g/OErjxcJqRpaxTDx4rU9ISOJLvdFcyxUsthTp
xZ/d5JFjltpsYpL6ljlMxlJhqxddXEL0n6MiPrclhg2Pa/oLRJwXgHbZUhdRh8CxBN24DujPAVfQ
QSiPuCV6TvmFdQ7VzrCA8VtbjdC1fg08eo5oQLEOL3rleH4nzX1lfwnePwZBItHBep4db6IOzSav
YVXgwGACqdsFftIBweA+rVYQ/Q1wmkAb+Sje2YndCHw5rrPZ+ST0rL8lDZSUE0p71EdKteC9ybrS
08P3AluFk/Y1+84jEDmrfP7XGf+IkMWA1buOYV6vMfjRKErtdX09CGLKdaHxVDWVI3vMddN/KeU/
j6SrNcfKau0dXtWSXXfvIcNa22zfGhy7sIO/BCZGqxhkmxCLOHQGCF38NpbcAtS9i8EvecsVclv0
Xob3WqDusY1jyqYXHYNcdarrCIRrN3iVtpbf9I6E7uspE3fKe/R/phxFYWHYtMXCKIf6/DdHPipr
/9WufhMJImCCaj05Njyf0KNmR1A8ZcbG7x780pa0THsXGekBQWVFBnvQ9jqNkFlVT3SXS3bYe/17
2K57GMmybWs5As52+Ja3nmnR6uFGkYzo6m4ZbCQ1YXqMsFX5UPROroPP2LDPTiYBsN43vgA05aLq
T91ouQUjhXhyg4xaJ7Du4r3bn2ALmUZwVPgNA+r4sEu4uJD8ReFxPMhC+C5WO7HW1t5RKkkeKZKC
wV1rgUJXQnOEo1px12rWc7X4MP4rfSXfAVjiWedcGbDrUn2sDX8ukHH+4HcB6rJhlGcdhNn3S23V
MqoLjRNCNYc5jR/e+LegdVKN/ixDZ3DJVN1WVZrhxEhN8nrsFZ0SqnWQj9VFtY5P6eeu0bXH8Jnl
2gNbr8KDWWZqRg+wKkab1iMPfwgKBoEsfX/wFLL0tQj2bfEg/wJcNSa2d+BRkjy28WRF6lnm1aII
2NKIHcG2QJwQ9XHMt+zA6lJXrn5MnohBP2mMX96oOBfCRdO12AMYPXYPtERGIQivop892MzIeasv
exLBiyopNXPdKXU5sDpqhRfXwz+6e9B1FbNp5gWoXBK4ptQ4bCcP3pe67LALKt4on1za4cGcDdGc
EV+sfRXONsy5XX02yNLgjfX+ar8y2D2mP9UTwH65j2/DDc0gVqLDRzY+hcrg9oWQBcxyxRxGakYh
+etOY2pn6hmaoN5zs4GLRCwjewaeGekPYuD1Xk8obEkc5TVNv9k2/D1K37PrGFn4UnyIoWNd7XR4
87ayJBXOHrhk/AhFYjEtDFlQB0FaZeWiRv1PSL34tdrJvmk9p6YvkSFW5wUr9p99P6UsRW3gVSv/
k0gACxP6PU67IfLtQefgnXfFclGP6K+eL61isxxy5uv3p5zBJBo0ZocVeljrhXxvNZzJe1sIbBwW
bjxawEMOYukm1x4GVjmODDgCc7Ns9ETZvbfsFdbgFG9poka2OfqMFWzWmHKxeUtAG4pb2q1gOiVI
ysQmPzWnaaovpDJ8CfRabqQ8JWNldRxkflQtzs3H/+HJJIcCQn3S03sy9GXApLrt4L2Vl5/ALU0S
NQ6DfczSvmRLQHqmveBmea1F8MUxiyOKRePHBhJ9bzCkKmbkcbbQLe3k0lpOjs5AZQBY4kHPgCpo
wyY+JnbvW0NHFAn4xCDIbU6KOW/kvNqtS0Vwo29NMpLKMV3GUOQykyGyMwq/mAYoLpD+NEu5Hetb
rBmeX5LebZHgDJb/Mf9uMl01zVShpISfJ7zoqUi++F+qxf93EJ4wgZDy5ZTw02UY3yzh8rOUoCZ5
9YSxfPvGUxuJ3YG0Lx5VsaNuXTl/E9aNJM8tc2A5hQ4esnevoNALrRBfeJvlS6Oi38Cxl2eyfvIA
YeBwtN2mpB9maQuu/o8x3qB3AIomM/1jE898ljj+7yB771od20DBHOwLjZ5wZS/52CvKs83JWgma
SgPjNrhji+W0ohfQREFTpqv41z68XVNNVNWjvMukdzBL8M8A2kNKQxP+1pqV6eRF2UidvYObe7+k
/8WCbeVl1/CNVa27U0R3IRFyrbtZhjjG1StXx1Ok9JboP5iYwG75EdKfeUjbshlHQpVU/WavpZBi
EUO5tjPvQOu0j0bq3F75tlLDDm/cNTE48Skbhn86yccH69fi/ITrxuMym26CF3Fi0y/sD7MgTD6X
rJgMnFQh/KYucQhqVfy87MYF0fVhlBhGKivRZw/0jk6JQ2SHZUjhns99z7aQgr+yu9p9qkvNLeBN
TcdAOdwMl6EP2dPwrYxkL5JcCV29olFgRwuMKjBU3bGQDgCka9f3iXyShuSFoiwZvwxqn+/6BlI7
kjYbed3IpuhYdxI8DhZ1ToC4jzW+JNj20Me0iZYzSkPgkgOCzOfDy/cOUy11LNI+I0YT452tO2Gf
ueDdQvwiMB0Uzza78elJtZ5yu64cpcsmfArzXpjr+McqeQT6/s+P1OBkvM8RNsBCR/QXd0yDv/dk
gso6mxKYvVF9Wtq1EFoC/py7BmHUkk9plb0S8uhXWgU1sLgmT7KBTTDs3G0LQQt9zVpy7xs8C65x
oSN/UFq7qFS/UHBAk+vDYLpCwj8yBUYKHiUfNjGaVZbMPa1spezdhVnyNf9vwhILRHvwZX7OEtLF
AD1DATt8LXaVEAWWuLK0/OUSuSezojujV68dnvBXdKjkeSvZgmfLJaRhwKHTi8iWL4iwZX4b1zgP
49WegULLxwLvnIaF0f6kgIAdO0O+jn3DScJFj88pXOMDqxSZS3FcVoWUgSH8YxNcFqCKoIvfkYAL
nJSVhvLK2jCac/JTUIhBa2CZ19R3oyfQ0qz2y9YbX3JI4ucH/oD31+LH7xQssD2o4JiUqcM1D5M/
qqDA+kNBEVgzTYWhrbFEK/oBR/zEhQ0cAQ+1vcaCZNHZw3pvZGCQW+n8MgRCmLJBpGVETCNedX2w
9LxPHbfBc2FuYCGiqPUSKjMdNhmD0yfPgoQWH/DRsNA8XcWaXN80/3r2hYXoPS1RxU5t1jnXAQAP
Ih+oE3frw5u7AjK5QiuWIrDpnoXjycS1yrND9fnmS3375hy8hq7ffkAFCP4yHJBtlxwyZiliRubi
vk+z9jMc8BzVlAM2VZhI+vYfnBniYNE/348SUC+etM4znO3zugJK16uyehcZD36qaehOiMUlWm3q
KTS4eXB4bRuVgh2WrNQZC3wPxAQjcnOq3+/SC39oC+9/NXGmLPmvdfn0uidzL8GOCWurTe0tW+3L
W2k2D0XApvPZAXFMRhxdvSuhhniBTbr2Nwyz2rDumpVcM3rjj1NIBL2xNvgKXkVvRbFh4fV2wbKP
zdzD/caq7D9Bcthd/gKsvMhNZ86nePyGktDQ4VU8fIg2f6k0TWamMMg85ypOJ0RiXp5u6OVQRTdl
xvP8QkddgXYCxBz//Bzgwnr9STg/ZR0mFzF2L5Mob5yUrDCqHI1RVm9/i2yoMTRpwEfAYkTaE/e5
1YN1JCFRGZ7u/MXa9f8OEhdxb8v8M3Uk65CQQwe9N9QQjnVFfCcemrHV5xl+tSxuNq+MGDSeWOlS
+on8f6IMuOHD47WHFHzDfFCgLBsLouIdGTwHFM8VHIWjsOBueDs+WCvBkTnfBm3iLslg9743PjD6
ugwccpz6EMNqFzovxGG0TzSn3hasV5ZbGxS26pLwYh7G8vdIMeJ+AfB01lPEOcks5Z/xw3dAtkPV
cdInz1UsGvAt1WOFu+w9ARQ1gSPCErNksylN9SxWRLCzsckd8OxfO7xwrNBtpxYCPafjRp6geqKd
pZ/p32LAnKzcb7a813JGenTBgk/hkMq4J7RCl0r+4M2L2yv2DmsEuDVaxouPH2bJ0m9I4SpQOmox
/mGkrXb2vy8k/mF/Z0o9eySC+OQPsQTZzeJncKgLVpIgz8ityK7fPAwHOiKJBlPiJqOVNkfiWh2o
Flyq+f8RVHJl6sL6TTAyO7CLoxjKyfF8cL74P5oYakz9IjmGfSn31+6KreJM1a1M5a2bHgnP2ytG
xxmeVD/QddG6c4hxADyWQYr5yFwZ1fZViVIkacGz1ZaQDLRgpOj4pCmdK0oWZQhIhQLqt8OPKMYV
3v1MusZAEnW0yoyrczcOvzU7EbDnazt+6POZWPValLMDvzHlxn05b2owu+HvlWaG2XYeCid7uv/s
IdCKdAMp6yO9RgBL2mbyMNP3lxOMY4JPXtbOUf/ZZPbs2Wb1LdvNykekzwHe+/sSsfk4MF7Hh5JU
ySu+umLRxkY/8/lYQ8moik/Ibb0VrJWGHpLOd3LaGKw2sY6KO1LWgwLtSQeK4DhV7ZkdBtZFnh9p
ZETzBKnRxVUe6TvoGbiWdDHrmBc+B4sTkUzpMb2idbrLPET+B8WH66J22c4D9DGwCWQIVEotIwNm
kEBF1fPU516ksnkxrshRgo8U2znt4ioqGxpSUcat9/d5mKGcQuSMvxlHRONTdGpIKZTQgiyhyCxf
ItugOwOH6jA68vY9ZCNG7AVQw3nJArBOkSRMHUx60g0X3QOcpVjGgPP8WpRvbB0TtLv8e7CJeZ+h
dPTASdRYjNNHZX440m9xFWwKD6M/3tQiUzgiKvdT4vT+zQ6sk70fsnl4zn+3lTiNBSTjybFHFHHo
Hi9+7W0Pevxame4x6Bk4+ZL2+UtKslgPd1vKKme6O2nVM/EI+K1Y3O0RQah75Z4gWrjDN7j0Y5Il
Z+zdD2wQY2Pq9GAOSps1I47dwxpU06PZ5AVyt/QXQyJn1sN0f38d+FmkZhEe6Inrj5f1sB2v4cuR
YsIlc/rPAR4wLj0OHUvhkQUlsxFK0NyA3chvJP2Y4V2k5m64qmbfZpEu5hKaViuZ6NMqvkrl1pad
Sg5TQ3OduG9Lpy2dxff7sEjOJdLl4hwLN+8XDjYfZGD5DTT9e36YmEVGzLzw1BncIlhxqNqn1c4B
Vs93uPB5/6ekHmypvaj4sZPr9J+BmpaSPcRAEw8eiDo4wFcyU4+6SqMfVS/I1RYrWuTLVQb29KEK
vtxl1Oyv7eSVhKRvClvhkjy3OY9+UZ+2gSN0scNs0ohnfvpfSr+P3lhi9PQMsNIe16MvhUlAKVOk
rOPjagNqslp63r5LK1j9rN2zbDgmP2dDur3In+9UKMP9B9lD6owKxjs1ppwK7HIGWYgIdcRJVpwf
sK45eBNCJ1Cyq0b4Ez36wqT7eKz5U+J7KWKEYL4+PL0k1q8S05O/HWotg8qLEg6+O0XXA0WaM6Iw
9fN8EzK1YPEkD3l/2YM4J7rY/BoLEoOAI4QLPoaMb4qXpTdywuTXoT9gFllny9nJcuikd5C3YKXk
jJR6N1cJsGQqRzpQcBXAKT4SsQpN0PwDb6wCQHEDAm1MQkuKXzsP9y/ktx0Lb6Gn64JXb48NxudO
CBfd0BOuMur3UB2oYEVlFQAIDVLzOCDAp7a/TrVGd5XJ2NSmMesy3spPl61Nv42XPhdedjmF0sE7
agA4TPDl7MGIZUBXxlk/r7bAGhOba/BDodutGCsVEGzkHTt8z7amzNwkbJiOOGPJNSZsmgz71squ
lRLjQiyETtAGSGJgVqWZQG5Yp63YPm45ZH7DKPSxRcbL1sg25UEi373jORBK2UMMyV9ueunG8XHe
zIVr0HqW0RUmRJfZkrT4QKr/8d3Rysmu+NmlqEc0UUnxV/JRS3u5srlRftsOnCC94eU/5GUwhTrw
UWB+o1+LG2ajuXAX3OjkcYzw9hmPLh3NoN3t5vmcjGchRYpeu+VY2/uHV6EqTkwckK7QBfA/G++M
e80BNugbXzLAp3B/hhWGL6uQjPan1kRrrWqZC4C4SkzSc5SmNPxLcyUkpouNpuHtXNjr4SV1Muae
yxM03jhzDt6m2i2+poLuO/pQ6dr5EhBqn54ZsMvPH6YpblG3iu3UFB757LH99d2pMpdcXKPVoG0V
knJlw3X/8thhzv/VsIVo4hlyLZePWWZhmlKk6ashGYcG2Ow/YiWkUdQW1yrfc/iZyj5QieXguDQR
7YCvqcKqM5xNF7W6WpSocBDzE7RWSknl5xlIxsO9b7L4OTwD2hjLi5gOKa/Ve10MXq6M8ypHKYUF
6BMDVKKawTpjNUWhcuUE2FfyxBQheqhDRC/5i4fk4FGwXYDh9BUgL3ui9/j8V2dNARPwh3YPkuzK
sADus+35AQUYljoE9CgxLZEmVFfqJiEDA0qGNloLjYAzv4ucDahkSPplm9p1+uOg63OdyVY86gfn
wlWpDLm9jFFIhLMEtZVaDIHGj8woWYxxh3N2jsubI4D74iZsFYCP4DqV5D62fXyUE8vR7su8lq6E
cgoKiCvSXYUqAnvlt6YCPxYuOVZ26hRFkq+w1DQtNheR5uMz5OiH4rMfeNsoqsNtpVr/oUZDpGvl
r1kW+jFRYVSqrwbmcOz8XzudA8UQHu4ThC0vaMC2j1WX1HAA6BK84a7hR7sfdkJVnXdSEhaS4pnQ
m2+idxhczfqPX8X9dIui16AYIHUGrfklwo9NQj62+XDsPBAO+QmF8MA6uqL92qmx7hv/xuIXrX6u
+iTpLGjBsP1mLfMe9voKabXGdElGaM8G3upmYB+XQvTdqhjm3vY0HtMxyX35vbxyOZa7eJ6+PY+P
Q9E3+1mKDMMMyUpdMWxAq9Bg8byaVdPceEn+6SA3bheDfFTb177PVZ8R7aMjNvdEKHxMlSMIwu6M
1OzyzIvRi5N1+JytYkS7JQIOTsPffmrHilJpes341XwTsRJcpI0roPZM/Vxzbg7h7o1n7156iue8
o/DZmtaKKipnSnIbvKSs8iJ9bEv7AOVXsE9CvDF1ioRNilIujoocQIMwOr+xvrDUF1EGZoFIQTrz
gaK/9OKusGfo+6TnbszVAzM6OWtX7VVQtt7JHJtDNd1vD9FAc3YPgFc+N1ySkfRrvKghsKy8YcxW
NoyELpI04ldLu0kxA6j8/62mBaIkRaMwwJin9A5p1qozvTL1OlmtNe54t1FezP9CjjL8hkhaZTNJ
vcfVSbNHnhM2faBFG5CdHL++gadClWbpRxiUWLkDGletzxfq17YyPKwsgc9yzBCok7le6T22ExVW
z0cGLVTHfz6HdQbu1DNXuJXb7xwZurVwz7TKAgmX6fuA7aRWoh17oVYE1yx6qVqiqg+d6NSgoZNc
phXXRT9PUXxkwirJ1/K/EJuor8iKZogUrzKzGpEdyeB1mFagrWM4dGSvbUBqUyjttBNSXf/D5iJa
5RYB9t7ktoIVemkzIUzTDOhJ1MHXtYp3w5i6I6KRRHHzhpbFGGyXefQrwE82LxA0v8Ywda/ewSNX
7CRIQkFfIimc8+R7+r39iE87tvHl9a0uIk1yd0GQbvoVwhrHDKO+++Njqrfbv44HTNgA/69wv2tP
mC027Dx4yn69fHb+qN03V5dQtfa6r1jzMlun32/hZEODuZ5uInDKk6rdxEThv7aLIeuqazFDa+2B
6aRIc/AYjWfr/3iYdKEZbVu6PEw+7wbOouIJoHgEg4fA5Di5ty3mrwARE1pqrYhqHVd7RLonAibc
XJYR9WGC2bphFi1SC9PW9u1WBIvy98YL3jcVZjzvXTLYoztmG6PC5d0ikXkpZK5rq8tCoSjcWxcs
fjWaxPI7C3V1Y3D0lEhbHlxMWqhGEbsBJK2jLuaR4iLxK6H/HfDr4Td86ydgMTGklc2oFwhnCWe/
cwoxwQd+3vKEEJr23ILofVuVQmDqgUDbFn4ZLnLJNBnh0rrS6aiJnpiL54CsT1qqNnLEf1+I3CoU
CfDE7hhjAwxK+69+ZyDwbZFLMwUUXaxkJ6M2Vr1MFpTDwzDktK16yROfGNkqXjpwRQuAx5OsDIG0
MNgHFl1EWhjZICpJLJhhSZ0VtmY2owbjj8/SYQ8151iEkgVyiW5Ctf1Rybu9YauPPNp/SDS9JlLr
qbmXqp3Du3LngLDsdzjT7CQAeeGebDRvUNznCksLaQVIydMi/hY/F2nZ1/vMzlh+qV0agZrS95YH
EJoO4dD2c+Uh86Hw9gnZbOEdTqUcwjHWwKML+zPcyuy+2+qD9FGwwdxP6/YBtyVoOqgg0p4GlW2d
fdQPrDtIJllZABdtU+H8Zmwu697n0Zfi0yqYMw+F0tyxsBUAYYzbAffPJHu8ipbUR0FKp5ObMSsi
BSYLRc1eJChNX042uRTVurNQke8KdJQ3xHyrc7jFNgugh3ouBaGX0HCI3jJjffV3OtSm/afmZohV
XyhIEphXDZf4OrgfXKgr2mK26+ZlqUEU0jwkMeYpEiFf/3GaeAn3T7RvWZcisQXt2JL1DWXxl0fo
Bu5bGVehFQWfPPDfcouEpH54M6cMTGCS/TUql9aQFwxcFWOe0yelURBjtts8VXbWhcNeW5BJyEBm
oOCDsPX1JxYXIsDrbOxc9oqmEIKGzToiVJObXeAfatijJJJaMuFXOZNAC0v0U/jTl0jnhxphRB+H
5lV1HqHOLyfOSAD0MlA3OGtFq4QaVtp9reLLW4SFHswo0tgrqPNUrFPkCYxBR9iF4HowTCtPFjws
gkea8RePcBqV4fGlBndrRPFNLWliXFLaH935btyGn07GdnsKoJ38rzEf0IB5fCQ2zBKrgWJdQ8PN
V3wdAUqrdZjtvyFcNwjFmhIts3LiJE4BW2xoY+xFXQWj0IXmv1deldxm0RdyUmWYZENkbQajcROA
J1fP7YDngat1i8yyxbQH5JW4vZzqWOODS84tXflXB6TPL27/kt8k7lFeNlHa4HmYGuL+a6A5Z4xD
/CCYicUdTOWkvNQvGAr2x/9tMNjattuSMNa9WDJW5RadbFtOwLD01ejHPEfEvAMRAapgSyLuAs/d
2HafzgCuGL1CpcKTEtGoQz4kEoQx3v3SWpAt+SLS7jKHk67AcuZaOHTua5oEehKKVKioBb2CyMdv
AjAUFiwajAbI1KJxWo3kPLWZ0N7/Sg0ptC3Ry0TWJJxdJpVbfAigdkEPqeZn/pelHNErVzAD+qUn
CO5RdgYt0teK01jlNo/uSgcmPPbFe84yTKBcup+jao2TGbR4S551fkRSgwiwVyRpeXWm1WnqOBIy
Mqa7pQZ6URyzdkHku51XoNrNqlOMp/wPvFUx1uo0WmvPLaZ12XkZsfB6n70m5pUmuOJH73cT3Z0b
JSwJX+MJWYqsaKckz0UYjAz18B/hNmLkAtudHJVhNzR0j9Lik0kV6rCuZClHYd43NH/bXDGBxDYF
QVbVUe1jfXRByxljGo08ah6PvnoNb0zH6xDlX42ZlrvqfXLyYP2AE3sCwFbyW1IlBqheI5m8jZPg
piYqi5UHCjkJzKdfNBqqF5U9iPxxKuk2dcSBAIbx1ZteIeW85D7FuWjqKjrbKU0PDB2VWfFtOY5i
zRC5jXORsU+B6tyN7f0LXA8vY0TmKoCWCKaUqj/Jou9Az/Fys4XsmxfwnI9opJCznaJhXfI6XVi2
nsjquwKaT9oTlu1Hz3ja0y+QVfdRH694Y708F2RS4C0aX/CgxipdhQQpiVNXrsVum2+purB+hEU6
NM2P/s+DVWgZVXtRko8ezCZePyJUhWx9QNUTqI06nF3SSKMRKveJHXIqndIX76/g0YgVjLKI9oxy
8FQnYUnyXMQiAU7vBD+l23+6lFQDQzFqII7fl7p2WnZ0luqBPDFtlQwosg9TIjrSPKmp95lxcPB0
dTAzOYYpJgy5/R9YdqLX49SYdUXFduRGZkNWxLFEJpMTEzQ8osThACIFPlwcwo36KDrua+gH/sM3
UXzS5S8+98dzI6wN27kwlZ7SazE22IFLeCkRRCAug+A0uX5/uZmpNSyLX5ChBM03X0yDroluJDuK
BNcx/LEg5XcDPjQLbGpDoBX+h7XcOdVXGWTyivF5LHmY5y/cwZLg859qVOUttzWe5ayiMDFuydxA
aWjvrz/Cph79VIHRox6Dra400ectXGIFX4lHqvj/5Z9CzZGYjRvOKkgyrEQW2uBrFbqhj49AMFcq
lBFo8SpQ5JayB2XXnvrGjGAWwIi00/oQe+hqql6oh7qb7Bszod2yiyQBq0PUO1e2Zyz5ztvGVBup
q/FNXqwFYG0diEdkvFtD3tPqanIuc7WWHLW2WiWVycYlG495QuUzgmjkDOejSpSY6MRnn+f5zOsT
I2MnG2MogkxQzNjbtsrI7xX5Xp+1NJ5aWOe8Ljv/XA8rqkhZ5wXVTEp9/WVnIGSBaJhS0c6XS4JE
WOmMuqUuNluKffV9K/MFs7oTJuhkzEMY/MmNA1Nar8lVfbkjLRbWZUq+Hy7Ae/5coQHzQHB9iOg6
BSf70vfsN80Y5oYVuYWn1Ml6aq5a27VPTYI4V/mM3kwK4tmraUHP19gyJglKzIX3GkotFIrbMygK
V4X4Ub5013l6b1ReRKteL7ZnjCZHrBBBSLzhE6leNziI+YMn/3B+qPUuMQbFsxarwTx24jxdth+5
wMwTwtnTuK8ylpDwZ7WGmiptc6tKP+cSZ8uEo/updIv5Wax3HNvrfI+QowdD/1gfONMgZkYFjmod
/1SY+q6mtujDnn0wgw+G1tfwqP4PJVZm83x9KFem9b+YRN9nAeHTzAz694ZxFvkLT6KN510UNK8c
/UGLKsSnFdhMBXANMMrhX+XQZPqAW7k9xvD5D8x2eDFHYo9QdzjC2mnwX1KVG5m0y8R0hjEocvaQ
WqSrDDjU0waQ3SwqvXxJg4ONVUXUPy3F3wlAzvBqq2KDS1a3EiQqPsTFetD4B1X1zatsuq8rFSE0
ZEczodvUDuqZeyPxiO7MLiqgSuUjdq05m1aPPGrq8WwIwjS3hp5UBserK0tKqYuzaE6YU3ZN+9gb
JvHarqTC2a2oP6ljMIkUqnmYpgvh/INWU0GRFKjjWTwNVTjrflfl/v+A/TMlfAnxbKi9DQbsiNeF
JGZVBi7SIbd1qCysgKkeVwvKxnLqAd1MZVzbwfPnP/Cx4Oev8RabtoskFOqlJ6z3APpDozsgJWTB
YfqcJGOVWjcUkYc9f0gyfPCYnQhtI75eh7yo/bFiKFXyrKS/zNWadRC3mzZ51cd8dPvR/jhDlCEj
HJpNUebE6aSMJp+01NMkYxFAil1ZBBGuhXDCk28zyJF6hVFKeRMsg/gPlrZZv1WD16Dc95rpz51Y
IQr/N6bmbdS78J1wOkf361pWgRBhZsZVlyoYhwQb6/CfZk1Dvw5CkHHrs3bOVomMpb4e9XuWeFeu
XwwXHFTDCgaR1sdtLpQSG2dvkHI1appxHncvAit54g9jP0fmzkAOWDBQvAZMko5KMwta2UI9lgKe
oFQaCcozbDDSFo/KO1FTcIWAQ2n43yhhJAIopzWKVqgiOR8ubAxcevU46kbLzRsJdRDG+q/cw0NM
gJHJbn/eWxN/WwEg9E4zABLdeWCYWkTlnMUAc+k6pH0n4GD1BCwFvEXWA90ibZDEvqePDyQ4fD2T
zeIwCSxXAGH5q60+/ds673lTUyIM++VbFkU5qKYFSlZjyYMQ3LoiZ1kJVSHdZUICEu6kmtI1SMPW
p/DNLCOsaqxhPMSOvCL0ugGxuD+XQS3Q/gePY7C5lL0RXWnPJ+S/5qYX65aJ+M/7IFdNypu/xKX2
qdJgTi+ONI/d6K+OOSCx6N8c3WblsPd04a6UFGVFFH03KckGP/Wf9Sfm+lkdFqxDqMVrrwz92XoB
RYbj+ZLO8/Nc4UJlFHDxFGc7DNGcMuT5mmjuoOdROf6wgLgHKkNvJoaYiIAqfeT5aqCn6vuE5Pma
2QtYN8wQQzD+kZ9XxP5oZixkKRyN43zdGhGczGZh6cwNq7hPWO3LWYnCveYoS10mGr2PFZb/60mz
UnvtHserOw5ow4bTDVkuGrw3asxRBPkcHhXB9iKcy5/y+WcATGqBI3RH7BQCv3Rk+XaRxWo5sfUZ
5nnrVVmq99YRvKKvTzDNDqevxVCPeE2VJob7+6rqtW0rAkaLvCxSCamBTSnA4enD+uaH+ZQNFFTG
J0EBOZCSLJp3t82XtuR5L0bP8amJ+wOA/I+HFfhSJ/xmAp8DuSfPEjo16jO8NJa77Zef5xN3sIY0
PRBqbtDzzqOA5SGzC7hJSUtPMm2agTPHIDUSUzORwc1ZidHTDp3nblyeujq/IF6WqgFiqxG/v5Vi
xNZFuFRMhCWfKF7v4PbmzqR5ifi37uWNx8Oye2XPHpy8fgusGLwUpoLchzgM/abXvVC+olXVWOkk
5lFyVTptQxShZt3oJ/UTmnVtlc083uX5KZgqqahJLK62waz38oHNFZHQtfGDfCWWEe5SAzVybdYm
DygMgLcM+OYsZ1kdmkM8MvWm6aQKu60d0pcNHiy1dDADkHSbEZjue3K/tSAliDuN8qrGKjHaWX8x
BTJgvF13I6kr/k0ZGjXqtXngPfeFABgbCo9rDSLHXYvO0UYqZR93+tdF+rjohMOoGx/ctlytCs/x
tKXVer/fMfbinhM1IyIZB3kgvCtQZb/ttVYD0UG7MbjVFdIumZSFijXXVqaN4AoMqDmoBZOMzM47
eKNYrqZb/R3keU39YWWqk0WpMlNqpVVCW4qY8e5ttxf++IS6uoR24j1b7cA28kE4ZCUb40aqd+Du
JJkR4/r8a3yKh4logb1DDqTx57SaYpNrwxSo+LMKS8FN27z1QB3BNRWDK4mRjGTItk3N1RWwN7b8
/qGgPaNfH8DhMjDBU0DGllujGaUll+Vno7fKtTo795H4SxNH/ByM7DkRIUOeF9WT1slIslu6zaNl
5/8Hjd/g1tXBszyRz7KCc2y3iVDLXSt1kD8ilThZ/KKHn9WGFnb3BpR34EWgc1JB8wtHJGZNC7/b
TwBevRKU30/l/1q5G10xRXvHD0lrwrXIX9wOSkq8ziG+024qCuAQ/uckMlh75Y6/Zun7MVuCVDMx
i4I2i6tEkzqwDaHXMwrUiF1utfVIIWJ/gOu1QSbyaGxliHu9mHQZiBpybNQpg9ymg9q7NxOwnngg
NI8eT7cCA5Y8LRZORNDXkdxhi1h3dZEv2v7bM+9ZFNkCM5/O48iVbdBj6tF5QGyv+4s3X1LdoXpP
k9kQuWRbks/0fROh5vt5MsRN1T22IgmJcBLgQp97qxC67xNyi/PUBzXgg4gcNvqNsUGBB9G9VUSF
tvB86FzL7iO62+dWNDSXA0rGge5oEFqF9RPfu3ogYvWIZ7sS38yRPPrEoxQuoyUNiHo7O5wkVvpF
4CTe/HFfJ52jMv4eioIkYk4/1nYvQtYzMH64zVJGEEyepGPNz0nd7L+i1y+1kGMK2+Mk6HUmJJl+
iGKx2GbD04dhEELv9G5qq2dRt3tRn3DbPFzqgB5SZlGkbHV8WJ6jREIsAfLBHNScg5eso3D+G1DY
MFncD52aKGGC3FPmq3CIfBQ+7sy3o9Mi1gM+3Y0a3SFECSod4kq6khjZmRAJhdQNLNWF7uuYmV4d
+fEmydjHkxHBLOoV8D8+TWigvnTs8rlO0QM3VUSsjs1lOwe7KSFnmnzdCwy4Jns5hm/Q3ylFjqnq
z59siVWoHCeNLPhNBrI3L3n2AGwfVvHtmk8EkUeehvTHGakfIGgb4pNI6TcfKKj4/H1o2eaV6E+k
ZF5MajFUO6x3X+HoIkK0Myh5ixnano0lRXFEwF0d17uoTy0o1xKcilE/FCT6zbJK/xG2k0YTbjeN
uDg5l/Y1G+lSi0E2vSqHsyk16vxAIOcruC33nQCu5IWJXFmaGUJDiZQ90G4P5lgTpoDw6qB8OwTf
Dw/nsNWqjZOibt0tZ4S5IGFFvZ8APqNXRwVvMd0qd9w8f76PL7L0fZ+v1mli2k1VFIIgM1r2aJNS
7iGyW335pLmgBkM9J9+GSYcKcbFJJi+7B4rVTr41fssFOCRHD1gBe2WidGUqhS0pgbIZkvR6LRPr
HFno84zB3LI67f1T/Gh7qfP0PymmKNi/1ksMOgwdD5Wtqrbm9e1Bj/58Ta8ZL/GkYSdrOXLkpFKF
KnLihEBNl0I2qrrozUUuAZ/o2FkjsGlM6SVHg8+FiHYlr9NjhOyDuHqR1jTdy/Nrvty0aMwfLetY
VPKpMDCICh7xwYv54wbuRDKklz79GAI7kpTfVhphDLJUXmNeM4FFwdqWDP51zwlcMlymO984lTHL
KV9UYrfK1fUKE9lRKWppi7RT5kS1j+5OOZKdx8g/jp5lGto2c+9qQQrOrcwB3/4xGKr5lor32/k5
rw3AHZi2L951Sf98Y4XpABtnOkWixp2grWazDAXY6EeEgM1hcKXZxz1ti7tIdnUF/3slpDF7tEAZ
rXRtjTmOfP6zcRmVzK6Wi3uGbW4Ln3OVSJXjQloqhivOIkSdckCyMJeBEjMmkcriRnWKIW9tRmmW
TfPf9C1fYwA6ZtzFwe6d12THcN2TrWlUkmYPPzhkKKXmBroe0TaH22U+5dwPL3lE28ke7Bvgsd22
7mX1NHrQiZ/KHWahV/AEA5lgfY8MimPUquprlFmcPWM2MtwUMrgHvgYOljl3V8eJRMUsgodCI3xk
b076FoNPKCugnVBTs+7YsFutmYikasZhJ/XZur5Iux19N5kCv/HIccwntA2z4HrAuOs867Y5ehvh
+eErfFY5+WVjj/N6lbxYie5f1mwd6LgWANazPbx9a8ufAiHDnwhn9qLJiPYSDM4Jx0kJ8pkkmuyE
cUSWrRbtvRJOPs02JxYB2T47sWDl7INXfJwP0tq2SdDLnf9cdNgagQSyMvMNnCvKK6lbN5y35WDP
WIvgzyLOafZYxY4sasat3tVGIXoYT0BvB3qK3PbnFRol9F6Ydhpd5xgOBf5FERkGj3mN8iDD44yy
FBxWxNwNneKgSkJ9YE5Z7Vjf4iN5xFW7JCHTdzY7sjWuUGy7cCrUUOnLD5+uk0JAwI981Vqk7R2t
bIcPDh54BAbymxOqqpnQn1HO8hzQ+L/pFmgk03OBpo5+B1nAm1bBWou/2CRNP3k2EL8VfewIg0su
4pxiOvKfpwcwylIFV1LSMyMHmfJIu9V7Ci8N8lLQLLJ+bGREyeELq709AQqOcgdkfA16grDJZlul
qWYAYZhDH6K4fCRUOneisMYt/xHUFuhBNYIBgQTMtic5eTPCexNkDxQABgc7oWVU9Lb3UycGD+Ee
wMbcogP1fKYCGa4sxLCegt05jauhCp47HEdUclCQFUoPXXOLkuf1CwS826+FC/vPX4wJ05vSrhRC
hZH1COiIKu5iHUQtM/uN7H+NaB8lRJ6QUMF9ikGGCpQz8yPfIqAkwFC0bo6QnJ/lwy91XQTIGtZU
+ddpvacchGFjJDFWwuCIEHW+hhe4H+j2f9pZtcNrfDsFjQa1t8eSMHH2vOa3t49cxNqqQ/4z8pvp
mygc+hMawBIaysC3TGRxuvjhq8IRp0INZ2fa2L8lcj8gCx+8OOPSE0wn0FQkE9t/cbqw1zE582tV
gqhazNgua4J7cItvDr4mM6plBkzEsTf1oNeZAX353B5kGaYKVEpehY8vSD4MrXR3u337/TGEpQIG
ZdIc+QB5GVCqis0f/JCrblAkI692kLVsIsX755+P3Z+X0ItNAdkOs3mFSJ8I+N+mxk5vJ7/j4WOp
Vr7K6OLdiGZzmFQMlqooaRI5cu1GXJdroxWrbcvBBd9QyUu1B/bYarS1zQ82nYWaSbnEpOeT3e7d
DDGYNDH6EWvRg92Qcx2niP2Y38OXEh7GWizNv3aZJ9wPbBSpOb5wzV2fxS8zoGUShQHh87N+GMKA
xGGeYxqZGFHpo5vaOekDEqH7kGZv5WJdhYQGuSZe3xIWXXawk/l4viUlVmDBZZQelrBOJZfJZMUq
cmod4SxV9uR+BwSthVdVwWgssrw2ObKRwxx0X0IMUtbHedXw3NXT1yQKqViyt7BqauPxhD2zfGDG
/+E0XeTD5xDpbu428EeqbBs48ni1bfl5ELTyXzuHFw0VW3+pfMqKBw57FU1+oSMw6+keCN7rHFgI
HYVIIXqEXGDkL3i3V3Z+gsTRMROluR7CuqlWOjn96Ld6+xLM3blfLBPFOzOej8qLzMtkYyYY5Eoc
0s28sp9mM4+I4xVWzpK3XZufm6HTUULQGUsSM97CK4RS4/FgEt87ip7gnxavm7jVw8rn6423dBua
zWnfq26fro/11pQl5OvTdz1L6ox34/f/BwSwgkLZlCwn06MPZbIMkwGaOAc34WFn9ctVo+vignfL
PpAgttZNHvYSy+qUcc1BShTr1tUrQ5stVFF9jdis7b4K+W6NGveIhQTQDhZ/BeqkP1WotdK4+3P0
tIK7s6OfeyIFZzeM9FTSlP+u/z7BjSq0eLSTakUWmOHTCpmgG7gll/SwtabYyWcGj2GfPQWzQaFb
t9DoAizL23wXzk3BIRkxBVSVsYl9eEX/eTvTwDwH4eFsubWUEOVQe1hYfhR0RAou/E+h9E2RoBdM
pZf2n7QgDqiocSybTTjbDSIMyzW+roqHIguF0EmhSQNKT0gdEh1ePre6jExNCMZas4OFkJZp/Ir8
AjU+jq5dayEiX+t90de/g2gGkJN8z2FO8/fr0q0FcVHeoa6iXdZ/RS0A4wjLyjVdvWn1YE19ptMp
B3oyJ+2E4dDgzETiiL1QDyehTkC9809/wCSr/+KH2hmcmBC65dIVgdNof85qCfJQ20sAGLuCo06y
PDFG1Xpwg0JJMJT+hxNi7udlxowbxSn461nPsEnQzBgOgJ7DGH8Xbb9mXmsyLpa1wafjg+7ywiWv
Ay8aN39q+dAd2KcB1W7yaYQ5Vq72jXM03TD40AcTRWU1uiNamjdEBaK3MFHwTE+NqsrrIwxQQq3d
08oPVTskjrXMe2ekKOnTZBZ1fiyRBLZO08Oedyo7XBUNoiBPdLnvATbSmT72XXTXW/L3ztjRX60o
OKTeIIIpLrAji3FdA0TaMtTPU+3bRTyB2zfx5GjL8JLFGrKxT51yDJVRZ0d54IMG5nZ+My2OwU7l
ZVQzZUlGc2S+GtDUV75ckhjXA7P3BxyD5I3iDlbsyhP6doNS9cmSsvPbF53rwreEMmIxv6Wx4q42
tz/sD+VXGAr2SNtNl+eMlxGYek8V/40flqUkYxcSX2JxE1JNYrcKL90vutZBBSAPKQjb7PtQ5GnF
ih2JN/3v2y1hMkvUkxjkVQM9JlFUi4ixFXVhhlSoaKqOIfhrXFY1gCFfSYSPU7lDEBLclWnUXho0
1a3kw1qh1AJZif4oFUZt/gv6+vqNkhCLMLSnP9/j1d/2V1t9bBZ0Adf+VK3QXDTEbhuoT8Zo0MXE
Nt027HV96EJ5RHFSjPj5Rbefc31kPG5FMT7wXZpY1Cq2VCQh/BmahH3UmAsvbY6fx5wFtaaL1PLf
rH8dJmjbs+2Lp1AYNRVqYXkve2a6S4en/2W1MjAAHW3OnxPYmlxii0NFbeYKZGCLw/fiQ+Pl95x7
OVToEk7wlM7TnAxd7qcLwq2Ee0Hl6bV289xX8VqAMsKQtZAPP5o94gbroSfTJH2hZWgy+yrxG6GV
VHEa9Ma0BFKd0oTNbCKyBaGtTgsBAXKvb7YEd9eM3MBz/vui1iDVtucAf7D9lE9kgeSAPdzIExl+
FwFARW98QLoi8h60iBTuigK8GVAZ7tApqsjJ5eGnyD0lj/FE0Dj3dTwWvHnLnEbZWIThNT0L9scb
AyCNZkB7DSl3d0kjAa+Qb99bbffqtZ3GX0vcAR2DUBNII3XLyDov1HOuiC1qEYzLAGwNC93Az0wG
rRDNLaBomCnfRKeZAGzUDSI8Po1ke2FIws5VyBWcDcKoekdjyDrYcCdCZRM8kA091ljtqCPlbGFG
s6vSLSjtbEWNr4Q06RzB4KOdabho6EySSQyUhTDQjhF6sMOsQHJzjjULn9td2iDPXbaPFSXkzzDL
twxWx8rUAOx4yqWg1cFa1ci7dwoqTf4xJnLaYehN513flMGsThlGEB9dFM58SDFKJVu+dVXFMcrH
qfy0gczMR7QEe3PCCeV/RLw6nWMEbG72ALv//HJTAYV+yoO0XB99gMwPNN8dHE5reVcoaia3eKDH
N+lHajpcNb8YbVwdHLPvUrkAq/Bnk4mkT02lM1x7bTDH5ht88c7xGNnyD5ICOzQfM8CT6DQ/32wr
J4UpE7O3l7ANccIRNRUwg11tPxBOGqh78w0H5TvG3J7J/M0owJFgNo7XeoVPGw2hh6krFGPRa7z2
qUJEtZDPzWEYcGk1LUr5txC9eeX8q8LvS5c2Jhbmlt7fRF311Dghhr0z2ki0pIzVC08T0xc+aCww
8fZh1uWRe+ytTr9XLaQRFUEIkVULJZ/soMyc0tC1jNtpNBnriHn9irS7RC+lUu6/InYSNxP7BcSf
SFikfpzCaZeWVMP47xa7eJsGEqlgCT4WwRUYsiaaBrsKDAgaBkGOz84FUEtJJxPsKHm/2nu0SMU7
fG/wfkc81THSfCXIs8ayt/IniaGbbWzmIzyGWW6nXvAPbWY48JsR1sBg0C4c5sSQg7eM3S+OCZei
UgfKVFlZc1n9r2aA6jHHhHB1dbhymBlxs8DJLf31ffQ1YTL2Iv6F/wfVXAoVgWrW2ODRz/9md4Ao
FZCb24GJqjR7+1STfKGV4zNDKJ4qeqx/cLTqzpOzY881vEOJgmhMEgCN+N2v9LImjBya/ur2FFK8
YKidxj579JM0WjzugiGD+eXNMVdTuPAcV4rIEC8y/qDHj8EJFLCeD5NI48X79e6/WUoGEOTNi9FW
e6vuc7HGwPBICl6eqZwyv6tgTtT28H5uroB5pbhD1Lk+vOaxU0JRIz5v3mbc83R5lA/yPAR37U93
/ghmyjHU3ugIvUJpB7YXCue3sBPZxoe2D/aGul2h+jIEhNFgQtSSEkj1MZJOON+e6MMq7oXeV42Q
aTznRiqZqJgHHBfSxAKDQlG80fiERsfp/QNqwvKmRY8OJfklZLgNvMU3t59XuwNNy3Ngm/3/VY0l
VCljuydzxxQ1ylYJukbS5mgdUsmb7AqKk0YzY47sVzZHjNGTOCoEVqttSD5/OSPzoprJ9HHYN/n1
P44IoZXQ149W3ymvjRvf44qmUtzL78ccLsIuJ+2t39CIRq9+/wwgElxsdWus3w+KH8uSdFZHIozT
jhmq9arjj4gUO2xZZub5qmtb1DgiqC652vZPvEjuG2JNvYN93I+RePHqxP6gy3lTXceV27UsVcXe
88EaqPXwxFRAXDOusRTpbAWN17VnAwOoAP7g5stDDUP5rEUg+AVXd8YAX183jovZlU35ZymL/t5C
EHkZ3/PDxATm4vxg7g+NZy+SqkFMeHMw21/xx5OsQ2k35GDnTAees9ZCE6HlJz1FDt8DZc7cBF1N
P/qtW+AWuhz3BrFhoc4DoJCVIIsQNmXN+lzccPW+p6By46gnVNPpfP/Xvcl84QbnD5+MdGPwY1xz
WL2Dw6Oi19lk/FzuD3hfPksaiIQ3uYz0Zr1gO1UE9dIAMcStVoSesw4aQm8avUqjYNxy3O72lVoL
RFRQEIAQjpXyxS2c5hySJy8C0cw88inAdMQmzUPdt90s/r8JiN7Zp636B1vQg5LXSheNvwlhD0rh
oGjWa/MZIC4pVEmfzIudKcQ9TkvUrJmXqHPVHTprMe4oyuJJXs2YmE8QWBkhzOznOSq66sHrk71n
9ZZShxZ1BurotpindfVF49OiT6NvQCaMkcmd3t5Qs7H9d7/jX2pkFQ0vkVzgrKtZ9ZsjDPlUFGZY
ctgMZOBDh/8d+ufkmi9tSIh4Ie/cofMBqGOgFqmtXIaXBi7j9EZtsAl49BWKKE3u8B4VJ05/EzW4
YRovlKzbru3HYBb7cMvj7vTH26Jndysr10/dOzt6OQsC7O9m+nehclWwxktfOC2HebgAZbYDAS0l
1V/vR38wEV2ssOiIuvCOxFIUpLML4gdkC7ejDfMRBgUKRXw6YbOnKsNw2PzWZBTYcP/ghXcmeNgU
LrQaTnS59s8iZ1uOH0jICw0QRBCDVSxK61Qb/f0Q5A2EIsBW3I5YRVJ0Ub2yHYVvi3w2cBd14FnX
Y/iYthnTFzSbF6pR36MHydPc0cAAmWsjM/c+ZI4aoYMVqF3ir+gRDQYq8osJXf+GLoewompUHuQN
41esb93yck5rlaMrWkwHZDsV3PJOIEh2awi6BaedITv1RmKb7LV1U/2r7AU5wL14JJCRdFQmF7yr
FioCaBJgcvo7JnkIuo9r3sfd7FWfNZdV+GM4+6Tdnq43idIcGAPdX0HT9Dc4NbCktqFKwa8pbCTR
YP4sS8h7gMAzVCY4ZNWoYaVaJtdcdCSZBoEGt2441+3NeFB78YSOJANfxLk/25NByJLLT74/ehl/
78OwstxmOW9/ipTm/FaE2QyotHMWu+RtaVP1juZlAqID4gG469GcPnydHjsjNuVRZ8EpFru4aMx7
u0dovCx19e885p59BhBGYnVE0TvcbvZH4ZEtDd3P6vNP9WLsMm7WLOj94EPugUHpuhGDyWLcmOOF
I2S148tHI3JaQbXvCYil/VX2co0Q0E6oCKChgvFg+wLvHhzm9ISZpzIfDaycJxL46AkLKZ10HkSa
UaiKkLSi1eMmw0OUintHMi2Qk2odGuABtsK22EjNZO8Wcqf1lEceCqIEDwJZWHHeMLGSHc3v1lAQ
PQaLGCFg+l8jkwWZV5UQuZCXSeanEXN/fENV234j64Ib/HxSt34C9eUkm0kBFrso4Yt8vwu61+8c
pRndtKdlfKzSO2B6tzkxwf5/QP0EGeQAjQewIlINF8KsGthR9HT018XI9HNkxraHmi1xlVUbdQ86
OlQsuDYCH21ICBTCGEQmuapj1ABEX54ZcATdlgfxRSvqlqTZ+Llq7qAXGQYlDX0yyP9qr5sa+sM5
QVUqQ29RMdb3nW1vGo2Hs+mTxQdiU1FlXrFSnCx/L1PjSvf6beUn3WgZwApRqr5jnVoVdxEyHfaF
ocODSBLleclAa+lPNL0S1Cldgl8AVm3wWN7W0P7uxZEJAzeZqL9uAE9LlI9ekS5+s3yj5ce770Yk
rJosDgBhKG07GjCet3l2Ojlv2Ia0XZB71quKZ1Q13gv+fqlQ3oSGj8zjoYvS84OQlbwwtmsvRI6O
yyUoBf4/flUFnoafVSSQJQJ1D0FLKSkm4btatRa+KhpWoeM4NFS0pxn0tz5zLwgABjsHBEOKFA6N
PkZ/jYiANiZI5tB0EhmNxXozRP27RZ8psb24BzRdS5umtvQktKlCiU1ZnfnDkU9xOV24GOj3ELE2
QUZbQS86Q6RQMnxV+2Of9afwBf6q6qNsPR8c6QFjJaggWhDWnbm8iqZyYY2DNztUEWMAPc8qwLeK
zoGsLOHgIE2AXOjELq8Kzso6MawfyDM0wKHPve9afTMjwcg275icQg6eXEF6OOtTZi2Mbu55Hh+0
47B5myWYdnzJivzDVlo4KKNyusRdyODDx/FmO1ryrkzXPn1Qimeh4kmnjkOSBmybmc7or9abxiMJ
+khsyElmon/MuHQdOkjlEhutAY0aQsRUTUfEyXy5cYmPtLLjKzDmlBv12/xCTI7tdcVXYzRDznhX
5M3gSxqKflkQeEW9ssvAPdxz9RK3qIKu/uvNm02opIHlkEY3jnmFoNTKZOAbfuscL6MIjtJsO8e7
UGIuJztw2SOt4I/6Nur/4A2aK8u8op2YCL8eP19q12LnQxPoh0TR7OmNbisYry4KnCT2u9IIsDeM
H6IJqiHX3cCiz4YMbAJU0593Pcl8IYrTg43Mh9yGD0oJDFfpGpb6UCZJWakN0ity/6i2AHEtB/1o
HUco2M5hzzNxs6XW+KNGGcVVDu04O4bPCfF5TgFuBNKnPOH/Pc9ivKc6VNfhAiz5/8C5jWTyEPFn
uincOH5wuso7q/YEokWcOpAlb+ets7LHXvefKqd8Tg3U4gTWsX+kUhN6Z5vJqTCYqdg1IBPBKtYH
qRbVIdVSZx61tLKM9PnLq3Gn16V2LW6TpJxQU4VGUYZx1q/7kMTp0iHAA7KRHtGPzM8o5EZUirXG
CK/SzLFcU1Pf1CeU5HMhS4c/22RSIN/hJTB3luGeBr6D2RTSiTL3gB2sR1cYEc8II7L+2LCvTWls
xExcrCF0ZhBbw6XjZYPmbcN0KqRsMx30p/uVZEhsftbYCxnBCXLtM5k8PC9qiQ2Tivj4WrOyimzu
JtCqDo9FJfkQRdItblGZhszWaxXKllGGFIUuzD7clkV+H3Tzu8Hqcprha4NCNko7S5oevCZy77QX
Srt0P1j3t3642fa7dX7PYjnEN4QDk2hh7wpw7AWWSk/RPcduEeGzClu5ZoR4KAeRQTdQGh0aAJ5Y
IavRRQQTi3xyi+BzRQkDduGvvc/X3Tc2FVhi/NZqaBHmQHDoLixJ3HeboLe++sRAf4cHXpfrRZCh
I4lkpdndWLhf2+rZ2v34K7XqXRKYR7V6dZHpEEjq1PIaiT7M0vsPH3Almgh++a0QQsS10IJEDqYc
dbYMRvFlG/M4ibQhhYssODOGd5J5zzdy48Mh+QhhU1+y0isIZu7zdItGPYPoJIOvd9Lf9upMZ94W
yPLH+sWzaT1qm1L8G9Mouv1oXzPku0DLRl5ZF/qc0r5y+XbKYFAco6hJQ3i4XPdgejWXwIMQ9Nh3
vqosI1mxuO+smvoYopHhADWhi+DftXu75uHR27Cpik/R3Dpzb7w0i7aWaTyImFpz0jf4sPP1IG0a
javjiWDnJzsAolIiWuRxpUfwQfsWUO78ifWVgFAixNqk5PHBnRZGWGupUPq1Z7kRXrQclGCBJVTl
1GzvXOGqdDDNly5gYH/HTkkvImv5tmiUlikubeWVECK/t93ADP8sJljpl8Yjs3MtQ4cWiTE6rq+Y
bATVPZ1jMUYJt0bgYQ84N8L6InuhAwT4KjCWMDxOY3ae4WsgM8f8639D1KcouMq0WZuUMSuzQVcK
EhKNL9k7aFASXXwViBhqOybmEzrJ/+WJCS/saW8C0yQBOm+QhwmkiOlwLMmkVVNoF2hPnhzKhgfB
BSwBAScQ5mkt0S2gQOttC2Rf8BWXb7ax6dEbflFsqLD6BFu1eTWA7v7Ux/HyohMjP1ml9ywYbTxx
+1V70C3pEBIoff6gmgMgLM5IkK6O4jgyouUn9X97DRqc1pge2tpO4JXC2X/lMQGrqLumto4B6x5/
F17gHqGOBGEYBUS1/fQyKxIpQwI57mAQGFtGev7a1hUvOCK9+K0UNN7/jir8na/mxAN6ll4vmlK+
YfvOY4ZiyGJqG3vEIgsCn8zNsgfJ4S/0639Jm1qvdoAxas9XI81gl3IN2Cw24Ih/M2fLbl2L4JlE
/KgVtL7uqUTK0rQsIpHtaDsSoihMP6nUPr8JuTJ1JCWGknuH2aFr/iPpGachB4JphWqU/Gj+H4hC
P+EZsEtVomrshp5ms4Q8Pk9pIrzMpmwUUEjom5La1WX+Vg+T16KGBrhVtThaLSlX2DulAIP3X1P8
QhI4evCU2VOy95bu1Z8iIhNxXxDTx1a9XB30VItZwUjKjk4iEXfV8pYveILAqccUuqXzm2QthpDe
zdX+J7ODhBfE7zdfdJfcqbK2aBZTbwtjR4CoPBPuFV+j8PT5s8YlEbcxkT71MkJQumRFJ+LN+yhu
9TmQXazHMO8dW7SQsmrK9JoGSSATCKKlO/JBBkUoub8ooQxq7Sc86IMznA0BhFXouQ2HexYHiXKM
fWCfq0sAxieUYxjTmWZ/68CSseAVztFTe3JzIIuQn6t8Th5FRVQcQwmC70YvZFtb6lyQsFYzFff9
as1kk4wyJmQhBaY481oMEy+m0xgXy2qYtLMj1i3fvELgaK6rJqHMB/tMd+k7WOtdf1OaFQpTIQLJ
Ujt3GGrgIK3TB/c4ZqY5QC1u5zmm5yLVPD3SS0Lx7nhdhBiO9FDcv4mf9pB/qNiLmrINdYUc9kCb
iGU/MoTyHGGGCPsd5eyqIKAYFEGvqwDZyBbE60TVl6w3vSm65Hz/m0pcbnhKuKHhMfHu45nv24G6
qJkaaSqpTC1lhpkpBsi+fAMgg4mqwKYpF/6RtkSfvJ6ivNJ1qygOX4tOMfjaHak0uC1OeP6CrNM/
A1/3nxZT6gaUO13+1FVF1QAz7iwLfvXGMSvtK+akFKz/1DQdYE4SCqKgSn0yLgWLlOuyKvmebI31
qeTBRsmb/J2FPJO7p4929c2gJPM51lth+8vcyxQAptvU2PZkZlimkrB/lfTVmmR+T/ZIxdm6U3cp
jqGPU6KdDgxba9ntHUsnUXiz4ai/OLvxJkwth3epQlhE2jmHSt55M345h+q4ojnyjTC5eZ5pFR9x
dVZ//lRdMzlrKwSBdPekdGc6mRnmvMIcwh/aVPoP4SwuWH7dUdxVKinIccR+9bli69Z2wQXVblva
gBWWXR0KW45QAeB8fKIrp3bBVT0inKJ0yo6xy90XO/77uRN5yujINR1VwBzdT7mEipN3ZLIzog1m
MI4BdOADS+NQpaRYr/bp1loTqmfMADfwuAnVdBAzc/r5bbw1Rf5CQCsrq0Oe/6vS2oYFPmIT0yuL
esQRbeAknoWZV7xFGYMUVmcsAMDFYuty7FJLMgu/ytUv713niumrOjBf6gl9CyYqZirymTsQp1F1
W/E78jcGL6l7kvqHntKvgpKhfvDeshg1Mt26hQzsBt6+PyCPg4NNj4Q5ktLtGfhoZN1ZwG21RaRo
eFnjGwkyLhd+wH6CvC3+Whcg3QcZh0T9TbZZEIcILIMFhotNTiycYY5eAtCGXQ/8vuXFjvV64ll7
JmIBLz0K8eRKXdLxyQwZ6MgdEbY2XD7JYLWo5hub+9KOOjX8r7kQeM5gm/Mu8n3CWQi4VUi20Owg
Xdvlq4BQ+iOIxM1daSliqUzCsBWDQ33TOz0K3ceATWNDXAGeclh1NG6irP/TSuFOgMFOLTdg35se
lcfKJfyR1UAlkLuVougrOJflA0blbfRV7Wofh0z4ZkOLQCyMYdpJZFPIIvH9TD3K0xjYedvbn4Id
Ng6fEgPiJoxsvCasdbyofRCCMWXPwtD4FntxlFbfosoKc0wK0duM7IPlc2jFxBOn0nmEGgdr8DNj
v5IBZILWwmuSeaKONCJxAux0NUB5hjt+k6yrAk8vqe6y2UF1gIsq45EFqYBCR4Hnn90epfz/eX39
sxkb7V+mWXfP8dBovuF7eUKGuaAtf4sgw8s0jvJwHMvevZfibypkXW5dGX/mSe3/k+b3CAr6At7n
OEv7xZarjwY9RYg0xRvI20E+rTAyZunTJkD+bYpR3RBhDoXkghf0+8o3gIQhjz60F6ryTMAKJphb
2txSneEIjvS6cZDvCEJI2S3yJHJSv8PvoR73IiiYbnYrWND1R/pTJbUz4EeRCc8xNlwBILUf1Cp7
rQVV0BgdoqUejrAHslGa0JP031IZav1iWH0bsEAFixWQiCfbBM2mmxcqrxlpM0CLWW7mc++CdEbY
0++9GwwI8GQ2yOOgVi5BUP/WRJpf+RGwFcxRU7oOHtAZT1HQzXSRHajp3VahQMXEh7o2tjmnTIhQ
BHPffK77c5G+m/j9E0GE70IRsKd3ZaRX7jHnHqU+9xLgzel/AlVf0ZyEf4aGK7oXt7KYdfTE+6kB
GIR5ctCh7Hjp838IuIgsjrwWcGbDXOkoX3Yimr5qf4KO/cG1AoUP2KnCEuBNGzHRA59mjARrbx/c
MegsGGDVEWn8WlBwqsrLbeC0A+bkAzfDjAKeo2VFlNIGVGyxLIpUIqi+PQOCgDgKvU3EnapIe3df
r424bcsnS97Iu54Pqf3YhUWzcGePHDQ9F1VcgnFzyU/KSHOdyvH02xRyxYxT8QpOMCztmFNr4M/e
pXC8W6R/mQqYYI+rTEgCLk1XT2s7PFL9jdA7yKVL+pwVIqjZ09mM1MBEkfSvoYNnmq8rhHKhwclH
OW+xDp3k7Heg8sxmkMBSYDD1/IQgGNiSLsY0aU8IHOf2CFcj8Nl60KWpHG0JYF8ZFaU1Ov6Q2Ws8
pSNiZLmtxfoYzVpHKEjA+e+pbwEW8IXyOPBox4uaBiv4oCUeMl45nckjXczBIR63ySoiHKeXibtc
eZEHE4X7DYOfwLhZ55Yd/Ci1Ne4IjyQNs9cacW6kRPyR29cPgINsmzVJAImdZs2kBFlAGW5XztVk
TmjuKOmOFVPOlkVXlJvwalkVXOA10CDqfFhgH0p9Zt+2IMtHCaIizwERmtwHsZrkICAebG0VdDhL
uitYxVNWygrf9YjTNKf5Cf4PuGtI3xFUMK1mlU9wXCC7VVmSJ4x3gZrV6YJuNPm5ZUp3Qbh/1llx
QULxqeWLMCDLRDLnQQVP1xtza9rJo7EfsNNK56SQYPCHh1/3ciKnB37YYrwkjLvT3DVOdLuyfElU
HBCAN9jjN6nUl/y35VuudWjjX4pHQ7gTuLuwVriZe73fW0XUMtd2/VJ37iCHIPwAERUSGTaR6zPq
Izp6QwU6xdEq2Aifcp/XL4Olj1be+1xzl4paUCiqmeijsxYETxz724zHcifMae5jEl+rJfnmMfKo
CH5k6kLoDtPUdNCgBOI9vIu5+bAUw8KJi+oCGEHrv12XZQFK7bIRFbhvIxGLgt+/Etdz8GShM3Y5
8KTBFQEHDr7l6wCOXaGBfiSShyKnd6gYDLGHHLlgorMzBrYQDpziRLfm/6YU/K36bo9loLL9LoRT
Bns5MNk1cUSAeUrpm4UvMjL4HH1nKQzic8p7V1xiT8xpBm1IQCNtZtFPQY6yFbCoQ0gHIvnw51ck
7rac7ec/3wf3kml5F31Qng1PzFwRxSoqot7232eKypTzMZdrJmYngdr/seZt8q3b1FJFgMZEaRiV
/2USLKzmHwlK547ivGQa2TksOTjpyXZ0lppu2+vqFv+QVZoRabZD8Rtuhtgv/F4O2Oh153+RNpQO
PRbLigfEO3r7a71WZunNrHcCoWVbFDAGb2qqXiBmAloKJXYztqY8wfldyvZdAkJXXuijbmOQ21wc
ZdnAH+42zysQMpSRXLHojtzNJE9WK/Fc5PftO/m5PnwwD9YHbUxAHTstXa9AX6XQq3bvxLxuEgqJ
8SjjeWiPtoDVY5qz7lqYZWDU2Y0hc3ODwdobDHqrMeyKe+eWqQxMvupCK6TqfJq+IS84LoQpj334
+KNKDGPo0trKfhIAdo8upAJdy/rY94Y0+s+nkp0n/XZO01DnJYrp3uHjGLPNA7oMjtCmzyEd52Wz
wpcECLRra3asledF3hizqMskpN7sW+33h3uE27nU2W9NIjUH6bZPUCiUF4cFm5VkEUS0a4nPz1sS
aQG3ZYUTbNmc+31MBMSxYLv7+urBdTMU3Cxk0H1LIIL5DW3k2c8qKQhYyro9oV+BRpeYiJU125mI
hJgyanGXBHmOT/dSisunwEUjXbEsPWQPGjITecUnl4TnQdvU4+YaUhuYEm9c4qlf0wCJgdj38H4A
iW/JMFWIqChOEsRHhZJ+kBUaMvtbVPKgVV5BJoP+UhcUIhzqx6vpbgj93EpuqyVBZCdQGPQb2Dto
BJOrXYHE4uO9GXzVlGpHGwsd4U6AoSHkUDSpv4joE5JiX+qc5BWR/+7YoauhzmAoAeab7W7t+OHL
47be2SZq5cYMwWEVxxgGfMLavnYjdNllJPhziyVAcYrKj+O1sSHbEfa4+XIpB4rmjhLyQ6aKvVMb
orh6PcvuNe9vCoYDpIgC2KUHQh8SkpLZZFFe8BgR9Viyj9MtrOqQforLiWQjQ50iGU2mm8pRORyR
vgdqvw+MjLi3yxWL49vExFZaenLTg8OxSuxtm0YuYKdJhsqWRNQK8XytInfvKlKHnlKPJOshXDaU
8nsGVXZ7a22C+sw8+an4d93aSaoh5HMN/Zk4J8+jx1Z7Cj3qn2J/s0q/1oCdVAH4gue5T3LspOPL
kbb5YkANKD6mND3645jzOhoBnwxRrawCEyOscJEXmg8qdUq2XvUFnRrivZG2lU0cwjmpSI3Sw8Gw
wPJ1xuQ5rZh+MW5UFjING01rCmFDHs97rgHkkiXeKIvHpIbYJX2tdJd8eKHZwZAYaYcuRRu6vmLk
bxsiqzYnAvcFpc0RnoJt5ZEnShGz4iA5DL8bCo4jhQqNCBmlIHvvyDqXPIYGQOF/G896chLftQ56
l2yWIpQV00oelbf/ezHQRZW1E/ZtBUZd/FGHbBPnvFRs4pyZQBlUaCKVdZljLaEKJnp7zy9HzluH
j93OV7GFYY+vAcrAlBxxYswGsnd365z/PPwa63yaqqWy3WKxQCQgKPkzReP1JkCJVq0DytZeL9Z4
k9r9EIB0OPUTeOHIq+lLqgF+wg7Z75yvYY4HeH+HidNbz5LdiqlmIAscJ8o6/yuBJGc+iOhkE2GM
6VOMUXGgBrXJycyjHqPjFbV7qgVw0itUSL/KWCsbn9Y/iT6X+IdwsyObRtC5fs3q5zEYO4IsG3Le
r6C+25825EZcHCMC7lcsGyvXCq1SlJCpNvDM9qgCPq3nbZ6GIsnedgQAyYo6NhSlARK13ZeAjNNz
G2dD6OmPp4pmlyjX1c3zrccVqCfMy56M74/PHE3tFgOvQz/6gJ+qcrKlDIOi5OYp5QKAov8zZVv0
MidIEYwEXdc/7Tgfp9pUBU4VJQVOI2nWvYwCEcfnA7dxccAzD9IP2+UnWsVfEM6LMxDspWXVvkEs
keAzFr+Wv1qmnIVrlhie+hP75zgGghUG1odLUvhvE2rBBSL1dv7A6mkmGprjrBLARYKce3h8k3wf
6Lc0YR0inAhXthPWoAKkmg6fjMcgetG0PycDHymlGIRn7MFx/iWcuO2WnG7sWAYmk2mYE29roBgR
5aNMciHT9eCNaamdPtGuEd7F5hnbI5+VyuXxt6Offl9mMeSxcKi7ACMiiy9OlIQ2imIM/w1vHK2h
tlGIJpWWrtUcO0DVQFAys16+ZEtCuxFb6urSoOxEtbaCY1JOmJ+kr7KgrqONHeIxPVSiWHBhSiNX
zGvFoPVLhb29idnP+jN0UnF8jetj1EbbjeXz/8FzRL+1RV+pMHtlHvsNdADe68ZKrAS7irJVcM7z
1ziYhznhzNhfdLX93XAY5I/qLcFK4Il1e0dpxxoo+JzbuBIMRijdxU+nFSbxt0HfhHO3E8FFzgWH
AaDh0DPKvC2QCI/DGl2nCoFl+Ba26vtnBw+yrdhumqL8Qdjbr/1+g3yFso5iL39wfNa1QZ7Z3y12
lCwFFz4TmeAPXDgSZaR/oSnqdYjRL5pa6tbRFn8WLTLpvD5JKdHYtJdEVo/JmLJSXcGiBLcRgb+0
s70v5ip/OpDxKND6J4P0npFPT+j9Lu1QcfrLHKkIH0KqgVgm+jsPRqEhtWnLW5X55JZiP0fpNfWn
Y9be1n5YYFokf9bBX7pqGZLt1cWEywPb03V1+LOWNeGUkb1qIxviTZyMztYJCSsyNgqC4BL+ZtyF
kQCYr4wbp9koJJnWek8zppOFgjmDsK0bTY21G6iJ4eEkkrbJAtBYIGx3AihJRjmRf+qrfPARcLnB
4yLQzgoOyzgX+wOVrJrVdJv0cqBXSi7nQNSonc5U67H8h9CmNV5+PjDArSNYwggCOtX7y5VbIpop
xlH/6nzxTPHOkAPdaAOLX0cYOML+yRd6oYbEqjCWt28Q0RimqPfrKgOAq/eZVV8ZBrLaLGsLpCob
Mi1hNmRxZ6OMRQg5CX4a4Qb12WTEEPn+o1/PfEnMUlEfyCSld0Eds3H37yaHX+jS4wq/ETWhRruE
a2xIHuBDPNA0lbtMCNVU1xykMjevcp99m+TCjzMccUY0GArbXlFdCaLVazZB1hwtBTmmLlQ4gHjV
TpXof6vBWttreYOthddE/VONEhNsTrIFrgYSxZwJcgPFhcBwQwICkq/CWeAvf2iCS195GIId5Cb4
Ea2JTPaDsasSiaKoCH7xmvEcGW3i9Zu99BfcRWIjbm65qG/pk3HS0pvcDhny+/gcZqUXx5wh57z+
yipX/+1ADCQfjnMejT+FfR9in+ABQ61mG4QC4/pVltb3fg1ES6oZsMmG3Q6yvO60YtGJYPkWAxJh
kHCv5WnhUJIeegzs9hkRD6iW50AVLAnQWcgCmSvPHhPuIy/DdUng5cBVCPXM/M797mJZQLXYNbnd
iDk9UsQiVmtcHs1bfZo7vi3Is9u51iIXfyagTC/CtVUIA/PFKacQnMwaXNjIFXCzs2CCfHi3K1Ny
snpds3SllmoADgWYxFS4mBfKrgVmIHwUhI21c2yPpVU1S9ApzH4Jhpe+Ugdd6pyfRVQ6IMw/WvmP
g8iVvtRmYz6UqFTkA8E7YiJAtAqI6Ks5tWQekAH6mKRmeNJUMtz4yGHyD3QyYLSXqrb4YAWK0Vbm
oxdcJ1r84uxW0kad/tdUpzR+u7d/cTEfVedL43hCHj/Rm8w44Wy8Auk+8j6L4lv6qzFwV9zqTs5I
7SKTkVSu5JfAzBAR82MFBOat/Te4vaFSln0uBGDZwCFH3D8ZLZ19vCwcgMSwISk50QMsWNhXtt7A
HAN/t0qfDJ/3o3snYDHB4RLPEKFrwcEbkn2pETdtb9B/TYBOhGlGRSnPNxxFx/PAb8H/8+i9OLQp
DKPQRLS6snOdjvkg+d5bt5nKJRXsop2U7SGuFqlIdPYRif5yFjGPehKhF4MmVO1OY3NzZ5e//7ea
ILeH5U1SciGK4IHbkD7woGwjMecOhEFto1cnpw0vecyrBteE4whMlaCBU/YBXEcVBmZ3fQqbiY7/
XULaA3CB3g1SYz3+1U8MBc+BVPDrInfaETrFhJaSuho0oHN1LyjzQZBn2KnurGUu1YNhnSKErIr6
pYzdbCmKoi0muDRsqkn46qDmV7cxeSPRJCRAIFn9ePL4iTLz+4jO2N+IesNbCweu4HXSWjXtvUGk
mhc8yv6zehPOtoZJyuZXFlM52k+1sGvIYY1FtBHvrel+rQfjU2uotZ0XHZWpqPkJAGqEViFY5CN/
JJNQ3d0XCJ4shs4ZaxCE+KQBks5YzqZdcHsu74oZZgWVEw0H03BX9HCUgkCDrqP7LtuNWyGcte6s
KWkuwapEQIemUyg6mJLUvI4UvcqI2esF26dyzrzMo9kzmVQOIVtIi8ZXfvbIW64gkoyO4j7tllCm
Kw6wDTyaYzJG99gALbxRIk+5TYFlzUkYa9ARVw04nQicKmGj0/IVtxO1FTad+73cBWr8LjKK6f5z
8su6Gc+H+Bu238vn4fz1yqiliO7omTbDerFHVKGWMnZc8EnHP50GF1Uh2O+KPT576iiNaUX0uk3n
bsM+qjCbTyAEoP319bIblA1yE2Z68iiynf/wFtCDmdppu2gIJUrvQ+cYlGP6oQhlKNC53UM3yKPF
K7r6diXEc5a6R5hLMJY82Wq+PRGFqZeGTXmJO/xosPUwSj51BoEe0WPb2PYKP/5ZmjH8hC1QfNiu
yQHePqonl394T6dT3jagsntji0qPfoLuek9DbbJEc33D3hLwkY/fECnZpGdwvasUcf0+VMs0NX0/
L/ifBmp8LlcK1KyQviPdAVOrtwL1/mVtX1oxIXPeV5EbnyCo1fTm6U4ePu2nRhDoubQdAAmqGkRi
xcxyq2Yw4OptrQ021sW7MvtINR2iMTbHmQCWSWQP+4qJyHysuoYpEUfyP8F/XnGHUMvus9otR7GX
lYSuiMkgONefAfZR4dnlxK+YKh5WFYteBzHsJumwxtfsM25ZVNhil1W4aWV+B8n+mmJtG8P+6hxU
VE8kC+A1UzscTn5uJeL3G7AsatO8BfJR9IShLYNI+jf/hy1b80Ef57/BFsbSfoNpNVqfChYHJbgw
SddrCbCHjzyGB7qd2UhQgFfHcU4kIlRZtUmxJmrcyRRoQNcPfAZSIlkRkLdC9kOZszVAQIRJBrgT
GvDwDa+8oW3h5eye2snsz+diUlW7ukRu1kycFpErpTsYY/RdEbP3DsYHMZE6joGSe1tGroPvgE79
eOpQ2LzSoS3JdsB09F41FoTo3vER82yjS/umsz9RGvc6viXJ9zc1aOK+GEsbmi1wdSeuFARX/16s
he9af5lpC1VtRq93HLm85bAUUeC6NyzdJVwJOSpABXXEKFirSj3m8CnuGfMa7ojAqKLY90I876S/
5Kvy8WbX1WGvjJxS1EN28PG0+Ky4MArva5UxyokUTISzo+6jwacn7LUk8VltOdOi+uM/uv85XaG4
pZ9ExczE9mth7nH56FNGyT4P5dlvAfF1/zDQMbm+xImNcd1E0RrDkMXFGNu0v5MRhfF/wNcvSwAk
1g46qzu+W+4BA6zVyHibXdroVhDniIFw/NUW9rrHiVYmP6g/IQYw5IkIGmoOitBFl7juAKvdb83h
+4hjnk7+zNkQ13VxQr+W49dTvhGWkVln0gbP1WXS/JCnhuDYVpWw8L8+LOq5cMMeY1UEKEPd5AQf
pfresEPBldsM/yIcVBES/i/vvdkKP15drlOiAXzJfAd+horexa8UmRRmFo3cuxaaMZ7tT+DLdoOX
uXJawB83HJvWoPf61NhUPe0OFN05Y2I7Pjh1KIndEmYHDEWar8aL40fUPgJ8jDvGm39rhkmbM9rn
zI9iE9I4cykO+dqjgXBCbB5Jq9mr/DouRi61sevIVJoXW8CRfKf+IorAgYFa/RLE2DwADen8FCmZ
BqsZYF/HKTH0xiZp7NqdDzuw8+VjP69zz0YGECiZX3WzFXFM2nlBv5vhiatGKZX9mLKEs/pUOpvC
i/4+Nv7/UdXfTycqUKDQqyYC9hdBGBrnkhZn1NsD9nTTTh1ytkyYHJV2rOZDiqLs31EUTRrIMZtl
s0grkH3r/7NfnxvpCXfWihXTM6m+Zyjoj8UOR1fZz1r4CJufwb4+Zu4p+2pieo6BKd8oSk13McTu
hVPyfoZvWrSypS6dg2WFhUcESpMxHrcDvD+qoVna4s95kmi2neDGYthplN1xV+kecPH9sGNKDH0u
hcl2CLawLTZaGRlw0/AMH05br86hQnXS02tzDZM6ndnql5CYRxgzPyYtfLggpfVPCj52KXJww24V
uEsv96AthJesueHG9YpG/yFp3MBZBGGHfDKaJ1NKyD77SYcf+b65oXe5rOC0GT8/ID3Y8lOeJnyx
k8TvYNdd0gTVpmdGGqn0N4m4Sv57qDBc5RSDX6xr67E2uxizy3O/4NvR4rrr/9/WewcxaN8Pu6wt
PPl3lF4Pq++Wv7L0VTR0tjkqKeF9f4F34EK3lUXzNrLH1gNXErYgs+8n192TLNhX5iYvIwRhrSd6
/OCIVIt73xxANyPu33NirHuOgsQDeiy62DjHYeBT/lpMZvfxd53fw/kBp0xvH1BHtrZhROAaALd6
ea9a+ISRpu0tcdS2uo3X9E1kaMGWOmwjAgaIllA0XD9QatJDEvC9YqaiFUu7lUH15yBzCWzrTL/m
0QRFtQtoJgpr/eBNwt6hKEExEbOCKyLeY4MgkTU0ycap6RJN+P3J3qihvPdM509J5dkH7YfB2E8Z
ta8rr5/d9Pze32Lkfg2TnjClE/fLsF7UZ09cKEnqrxTxmqAwhcC+I7VVJEgmqxjCN2eSPrAZAk3f
JX7q3Z+1yqM7EvqcdM4Nz4G6j4YupHyjb8QPQTUVvTu2vWrDWaeWtCofQXCSIDvQf3GXqHyrk4a6
woydp4Q7JaPqYvhDqF+ArZkKKawONY4UFseiIklL6LI9cs2fuWWv+kwiw3OJosKU6ZM7ZsZ3Fa4F
swINzGgJdvX4c4ogXZFqiBK4nQ+Fj7i6vsc0WhAsYGw7cEaPFmX07+Qc6/miakgFZvJAmt31UriM
YQlt/A2XwGcM8kVbopsOWA8YLUSD3wQrmNaT6uPe8TN0femLA7Clvk0ZzxbFrYtQXP5AjPd6O0o0
QDpKLakRq5uP0/jRPj2PwU3AEolIHeg2KK/HnaXFktE0yGOcx2wWCMb7rCQXZTuntbgsGyPCEdqt
aO5t0RDea6KacNmdvh0ckWZrC5yyuNf9TsIpJuDnlJDszEI1/AaF28A7bhmh1Ly2OYmOrH6rNeSX
CWUqJkqMSbe6pCfA3JGEvv8bd2YNauIk6zRm4TaFEEMJbPv/f42+rLI+6iNT/dXWyvIJqc7X/TPt
dhUNKOMDv+33YUWeJm8cInh8hqaC0v0UqKNTgAi6Gt8ZLoJiNjPHIlFncDuUzIkM4S4j3VgcO8U6
V+AEOImQy6diH8fFNftdNCC01zcHMdvgnMs5tuAYa0ZQ62t2buN2Wg6jlcttMVuP5r83sM/IhbzP
2Esk07BH1moiXba2jJponajzKgKk1MK2PwgM6ZfGFa0DdOHZ6XS6jurCPLAtolrtAYkPp6b0w3Ts
ORBWfGXJiagkgJD5tmV3a21d6Bqml8Kd6oF+rg1U+xsaEURyoAucUzKxRDtGvtVmD2KIkjBjfaSv
syDsCRrJk/zvgJfMURTqnh24sO7UXwrS7elWb4VXatc4bYgDGIAq/qOI02kYndLCTaIzzY3MF4TT
WZzKSN1Qe+UMK7qkA8DfAsOUpO5mmoTpQF/ECGMZ2KxpAvZNfqbAyfMcOpX5AyEIDZ6HKpXmxg9y
J28vNZLK4eeMFLe0ZEP+WgiNP8zfynelZXRD/L05IG0t3jtXGygaV0DU7yFbRpkEUn5T+GTbsAXp
qkbQ0d+Hw87WtK7zDeDlFu7+35ixaa5XJTBgN7MesTY1uDYupeREuP2uxj11HVlRw7to1yVxASrb
zf6d+udDIi3iJi+18z36Q0J2sEPnMrG552XsWCh2EUpFNNCXHGUuC5RpsngddxqaHP5XxvowvPBv
jQuhjFBEB5xob4EPDPpGnXxD0fcicEUHyagFmrID1nMpOyfFxARoXftYhZzHgnIL0156RMPjkVmI
X9YTCiFpgdxAu7UCLdLFEtRESAvJ3pq6spgZFw8sdP9Xuo1r6nRkrP8JTkBgXKud1FwhoTasxYAS
HFpA76M9YP/yH6i3YvQcANavo2Qi0JnK41+g5R6dMjW54UpUtQanxloZRz/2U2jblRrfoB9UD6Bf
FHkySwk4PVUzp7+TjLZyJbBifkyQ+5L1gwqSs57pKeNXZn+NEn08/goOM9Zuve0hhxWhcQ8pf+M3
Cpwda/+IgYKfhDBCWlpLUIyYcZoa67ACFFzJURKsn7hLrOB1rZc767sLfEYM4yqWuj1V5kyCnzAB
NRh48zdqHpSi9ZPBh/Srjba7TVuWveU5TdsEXIwlH4OT8ckFuQsrndz24D+SXxmxNX9V8ryzZKS6
aD4At6rJR3yRrUTvV+gdrfPvu1E6A6MTyDmpm9zyUH94EdwCCfLBYI0OZTI3DS/T5/2RRGnZAigY
QWqpzYN4zU7huUdmrCTiDT2knEjJphKLZJwdgazeKbRIgexd81zUZx/pVV5WOwOqNIvkL6g6tU5t
UIklYTYtcPef4t4WuhBodcobu1wpBo6HV6tv9vtIZZvVGEvVSe+h29fhPcxLx5Snq1aOxb86Uh0Z
HMCPADo5K8/mJkH1UK0QYXBK3b+y2ugB8I5Cuxho3B0Ed65iOnQprfrUxAfhKmipg9tZKZxVWp36
/qAJ8Ggu7JcuhNK4b7JH711RvesLC7n7ghnEvrWtggTNmFtZcqr2zyj3kexOIHZA4xF/A0z0beP3
igzMKf1tMczq05wgDho7DS0sGRUp28nWZtBtOLH7mWn2/+AvTntijxdNHW8SrLK6euaT2zahlbwP
4lbCxUAGErg6w9r/TnS7gN9LYplIrGEjBqrvEZyGmrpmEjFENE4FR5EIy8Bk3aHnRusWxTudkJPG
2U9SDIfLcs03JTepW4jN/sW/l5sQgV0lvskU1UTmMln2vUnj3ylegT15hG+vOEbtJeQ+R03SOFyS
Wu5D+30rk7AflkjAqHccx4Z48Wc44FdsEjGO3d/bRmqAJ1/ip2s4Tm0BWKzOt3iaNAVK13EkQpAJ
fTde91VlZJbLnCwlQANGDDtmvskxq/xlxsB7O6xE8xzqAFRU/oRYX+B0sV+qN9mh6XxoaV14/szU
XGiGJP4A28GkD6YuYDri1Yg5527WBuz2iE9xYKrJOxrSl4bCM0AVRjk1ueHt+fmLrWSFsYI77vW+
7aiyDAwKqJB11i6YPOk5PlYNqUj7xwQa8aTuySvRyO5SJVTke+Kj2RLXXjlpnXO5nc3dbvB1zamD
8Rotx3R6FLvzgNo5TLMHb68Xc2TgZPa+uRq67bfGhhneX/JkpmoHnrSipVZBxO8JXfj9RD+gE1fn
RkD8fXJZvNDxREL4XoJWS2Wn4s+AMadXmqKzcWyRGGANYLYQebJjLhsEyYY3ZsGO48ezxD/OIFgW
MFfZIvCyaIKekTBHdWOF3AYQMRJMCDp7xpWiFGmmMog48swpk9UJmKBTAdqptvh4gGURS8dK0r2h
T7cfH43z+eWeHdz2BKD1Ct3PcW4XN08idpunvyLm88nlulwWTwHxlsYjPIuwuzROzMXfQblM2YG0
3Eip17AlLBF3duhlJHlS5havrZs3BRvkuq/MJUNPk7Q9EhCs76s4bZgcMh+B280Z70hy/1VyBurK
e8hb857exDiuWfpHsDKEBBK6IjRfk0nHz4lYJuBeshBXfWXU5qNAdITPGD8gj289m0mzYxkaqj+f
3+NCnibxYFAn+tPO/cy4wo5sP6hkdKHAO70jeoY8r20s0+QgeNFAVDHXhvnJt+o3PvBoFg6ee/va
8QykuqshzhhZRZUxvoKnm9q2V1fnbmpwmcniarcfs7/+eFF0QOfDUGklOL+EpvFfNygRyraeWFOB
0RQ0XZWk6UhWMlOdBz/hvNsEgfMHhNHfd5QYYU1FWZalFgZWPZNgNQc/e2drFfvW1XeigloT6Gj1
zBYd2f1pVKgmjdTccMIbJwifeYgPqfE7YFOaSd5uch3rcOpWNmMk2qMuhC/RPjwnmwVIZSY8ZEHh
KGYm71jDNSfr7r08mvVfLd4kp/Km7Ae7PoXhz7nhuW/joo4zk/zID5SCCZk+WjK1mbZ2Q016Xyxa
93wSnJzCGv9psBPPFg4XZwIO13zfv/eXlRkW2UlYdCZOJE1LK647h3IEjacZnUc7jAq9T03qQ/18
LV/qrN7+LZOxcT/9fYrne3j3CiR7CY7JJ+mxRULDz08RcOPJbqdnB9h/QzSkOs4J0wq9aYiFzG2J
+PzjjYDAqtdYxU7jIymRDv6x+n86msUMl1eCJN6+JsLzgFGqdS99MsgwkDS4AjqS8clCLakWW+Nj
QuXOK+IoMX9rHrhlJPsxY8sxM56I4E/EoM2rE2LR7hYGpNFtAfTBZ+iiEhgISo8aPqlKZOiZHNOC
VQ3m8CiOWlKLvh4Yo9/aCgdCfdggBfVNkH/nd/6dqJxy8X0ImuS8DDRIZYLCgyJSzURlDG9wcI6P
3X033SL2t1dy12kTECLwe3VewRxMnfXCe5tLWgHzSju1T6aZ7Xy1gG7ld4/B2h3/zL+UjGrM4vCG
MlZImFhsUmVUejWmCpPhUNqFTgsyWPHyUrEcMz6CFu7VaBRIDBCL31fdRsM9B0EwfqbJ8R1VSVlp
gzsyV1gGUN1Mlk1FdVc3DED4C7LqVogwITB2rtitAEqrpyI02oJZKEVvrvraCvtgLgX2oE6T6/pO
U+00bDiB15bOSD6yugwazznS+FXzVPVJEklB4l9TGnM9MnkDQJSjWxC4z2pjk5ujEQFz3wfOgBHN
0TKrgqiuamAMKQe1dotC/sb+jBi7HeTG0tA2QP7AGZgANI5giuQ6M7JesgJwNbcyheJT3yJZ7toR
n1XTkjRmced+TKv62b31/1PF13TPUdcRKhAhXRCxlf3ziWkebO0Z3qaBpgP+ZYIyTQAEQru4S+ph
HE4eN7/wMsB3oZ8Wpq34OiwKfLRGJFjYgo47c8dEubyX3FcFraWM22H+Nm2OaS6Hi3mSP9ha2sbZ
gACmFX1jeW2c+PP8b4uUdKXvMw6xRqo9JFQPdS3GbdACE/DUwYX4klcKX0g5/NKeVc8PU/jawVfN
efOuVxbn5Ybf0zB2AgyUTdCY70kLOCDWxQyW032NndyGJWbFKAcDF2qNzrgnKg5K32D/Shxq2WZH
SyOhuCXrrTT4/6xQXTJSe2LIe6chWQuQdvcgIrI4NRJqS5MuwWy4kQmfWDtbjZptJ/GQRwKeSfCK
fPAk3C58mmwvSxwmlz0q+Wdhn6kxQBSjFmfboFvH4KPz2g7hoZ39zWYWUbTK8Ne7Aqn7BLgMQwrD
V1SBW6S7/ekOKrdFsBPcnbtEY395+4LF96Ee5teFd0d9x5c0xByrH4rPvPOmV0CQmKCrElXjdvd8
Mzng6jIMg4o9+v+Pkxa6+AR0SjuhGtu03J+b6nzsQ1yTFVLg9/kdMvaidPs9DCmJt/tRf4jE9sqq
Cqo32rkH5g0REhgKgnCtndjWFQ5Bfdemk7pUm18aCNrv3Ie1AmFmvD9m3VaglB03XQmpf1xSr5z3
E7jweDbDIwHKHRrP1MotvNg73oasrbzdhrRS2jbgr3cSs+pa6QH09B5YlVShoV/2Ucj8MDzemLfR
ESI+F1Nwcp13plqqA1egVJvSS3QsNfajUR/tyBUFIdzhT0uk+/Jf6XFfj+AK2oayE3+J/YSBlwA1
OL9D3Q/+oHWgtlEr4Y7giYXJid6pyy+5MWKysmgRu9mvF0OmC3okpiDtLqdUnMBj6kPBG6dFCj/0
CUb0DEO/niFAiS3TZSL8sxIORtGNRqFP5KeUXoP9lRGaZ6IES8GkFLseBMz2hvpUgIsiLru+sFYA
lgxQg22AixvubA4OlsOzQCL9HAofxo/xUHwv2x5SloaaU3a9y4Xd0FWUBXeNRwsklEpiG+YTiSw6
LibwsfzCPACVoAfMHxt6mGSw8/3vCVPtMt2iDxVPe5iEyccGij5FIHr35WD5EGczt8QWyiel/svN
5091tz9zjgzfI958ufOFMzf+zzY1NDUjJk3zwdr0NtliHM3DahV+50w1Dd1PuT9juqE5otDjsAyQ
m+g8y6u/KUsKqwsNXxLxULeUsXXSKaBKxvvHmv+o4JENxeOP4ryBU2Il9Tj2z85U330lHhBFiX/u
OIBtoRIeU985UVQx2u8fPzAi2Nh0W+e6px+svmUjR4u/U8GSar8AiRZAx3CNG0q0IFJ/BHV8RwrR
/U+lbqk75L9nVXZ2EnFm69E9OVUVQfk7uu+5Wtyw/lihdDv6QRhwwZaNn1oTTN6CtQw0i8EbsTbH
S3KrUE9BXPTN53FKjI3pzSC7mHia1nnya7h9kNgID3jI8yW2n+JlBehfqUaiS5OJPb4tXzilNHpj
7nKZ6xmgO5X0KGHy7JdD2bYSC1KBXqbomr+GQ1RoAKQdQE4IWAlKPXxax+62KazNLkctN0yizolu
6dgyMYID/j02EB8+HSAQSWi5Z6gUNRfZrioCV2yphsZI1EQ5KRXG3OkKwFFw2aGlsAaDIOSfCzh2
tbBa0zGvu1qGjV7c2pUARkma8h4at3NbfB7g9ZQGjHP1bponuMC1Mvmb/uJYeb0CakNuT7U5/99b
UHIEnB8Sp7/yRBMWdbtLynMbWCqxJzHwbFuT2UE9WXZhAr02wONMoOtpUwhrmVRWjWUVT0tmqhUQ
V2V3TOMNZj2Pi5JB3rVz5i3KmWNeLEpR2yQXbCQUaTxlnrcB1fg8u1kXdSN6cF/rwpWClDkvEQXc
fg28g26aD1eTVyp09r+QTENwP3dse0IwHXGL7juk4JPXNfmSmB843Ypb+pFMVMI5TaApJKpjlupJ
tW/4hpjgmr65u2Fhiia8Il7JZtfcd7P8dEpAapcWKciWlZ1ASczyIBibNo3EVfDS5ma7QK4HZHkd
R1UdxQaHo4w5zlywvW7igxpHAObQzm5guZ1oQDuiZZvt8+mHQf6sTzcO+GdVVuXVulGjfRhvevr/
vkg6QdQjGC/iRDsWgSuzAysiwmhWS6glVE1ECQOExqwmvzMcY2pfmznzBf9HfaSueGKNZf+HDmrx
iR/wJXmVxGgS/M3xX9rqvt9JwdeIczYzmh+klUeRC33VvXMYXbD5jnGKNO0Jvcg/24SX9aaxnvc5
5jSS1XKxn13ELDju/mwcEMwVF5kd3a/sTeK6tSyjvYwg7hMlJH5+AphFQelg9QJgtaRzJzK6pnHn
hJeDC0+ptz85sSGkL0C21SYFmwDOsJZ3iMwQt1g9t9kYMCJJWQ2SCqbRAIgYPESYl5+qAliRrQ6V
0RePPOCugXjU78Flt8CldwkTEJl1iFptaeY3HBe2u8GZL9DjlKVBlg0XMOw2wSI5U5pvCrB/WNfb
H/GuqX8kwF7V1RXrvJGSHJBthIzCZ1hq4LSRy6/LdKIWQuFrYgSdRpk87zuXMXAUDbOSMx04d1MM
ChoPpBA5xPcCOhZchiOiWJCHZaX3jdsY3qCZozk88eNopWJ76SVsUatxuyN28bOB96hWNeb+UCK8
SZwti0BVd8/ninoI476+X9kUwv7yfJBXTgXdC4c9cS8747O9+2Ricqiolfo9YnAnUd5lhktObWbd
9TgvIxDYm4l84bsHw2Ijwh70a4n+0XTeSLc3SM9/ZJDhXRS1/gUfQPDm4rayXKbXHAHMlnzMcNex
M8YpUe78z/k5y7AmUNqpMIk/YTVsK4zfvRR2qgMPU7wGynXupgegeBj5JTMzpwNJILDQKzQKSmC+
6zW9Xpy4tYMeL9EbkXBAUQja+rWjzQwZ4wJr4Y8/E4+WKXY41KC8ZJEiwglte2avJTKepJgoipMR
VynUowge0HhMOpAsLI3zBQim0ZbUTX5alI2hBMz5B8N77UYxGQLE0fRp51yfe8hqmvE2SJuXqjQn
OkY2Y4ZxkCPRWpiFnuTynuNvp5vqkJfzVHZOgXhxi7qvfjP8K3R68qiVH5UCGrFJmZvkT3uCYUyM
GcYK9WN4/ros1vRhRd3wQhDMrvjTT2n2RLob1AoiRo7uus/zh6iBr/XiJYXRJhuhNhgp1SYZ96Xo
Qu/Tf5N3kP+PGUdEujSbwBEb7Xa9bKxVbqmAlRxo/CGb/rW4+pBayMKsL/sb4x8XvQq3IGFV6KO3
JLBzGcdTOw9xn6P8BHE5E8ij+oFTaKUV8QmuB8SaT0vjgt5bhzeC42sB+U38UHqvKftMvECsweDe
zA4HJv7sORBUreEuX6D8eroVffKch3Fl0/bgKxZOFoWscscR5orG1lRk7tYU4HAsNGrB5zZfhWt/
id/yOSH5vi8SrstKm6pa2hwrGrirIJaN6BkF2BnQ5lBau+e4mpUMjieGxXsDlrzmQjm0DsraQq7e
3xZaGGHUSjIinrdsgPq34L13E4iSV7bLhzGfGNpFGugBuc16TBt/wV+q6rFGAi111vRpkngKvCgE
4/kue9qz7/BAkASVsOM1rIyy9Y7zAZKYjPPhw3AwNZKbAavaixBNJhrg+ZKkWZsDCWg4wEv/IpHt
a2olfBxu2g/heBBOkq1QrSuqFdKeC5jJBBXVdW4YsLmZIWx5fItDl2Qyftrsr/HvjtUlPrVcqCsw
q6d1ErEm1+/N9Azhl8fnSnFf6NNoFOp5OPN+BimAuTCC5zM7SeQHsVrxxqOcvJvWXRyPpCeznu09
MWZvS190it+MEqR6b7ha+TciJ5HGNBpZryH2up2PzuKO4aUaQ3rKFqP9fyRjqbbolgOjWEG6n3LP
hyygrZK9igfAFFJeKUNlgrz1Di+jCyJCCIr635TMWGf3Cyk4jOXYP2jCysod1UK1I4H/nz2RSNe4
Yg6LyY5NXgyLo1jzdKiFBLRKaJEznearwW8FjTuiqlJqUEZEmuMx7w5ioxklIqoaC9pqN5YDJ4L4
c6QJ5gZcVtR4gMpRHBPfzxWbPmLlV/tT/xxU1J71mKWYWb31uBAhaxfsVH4TgO/kbPYHkiprn5Uo
/omT+XSy3DKLyRT2Pa0uGQgpt+m8Hw1jBhgFBxxNR2Q+aBzMnMFYvVDuZhocFAjhDAX//Y0UqoH3
mcCIokUKJplL4KSkxsMvcUxd6+GGHa916MaPjC6eT7wHJqLDa4Zlaw/rQgdmcMtss/7B1cn7QU4X
lq78jBrlhAPcbQEZXTd1l1Vn0oQT1UYIlRQ9dAPv5joEyhIocCjxnFBuyScvNYn3z5Q4jr5DIhKZ
WD4eQPRdKEMZ32xEhbEvLX6hIQdT9dPOdzmw8DhhRh72AjflvbQeG/9iWTRfypAEkKJ0ur7tNOsZ
MfZaSGFQYeaeREyr/5u3ZF6sN+ICVzvq9BUghTrVGSYNGOJd1hRZvK8EPkKnj+T/4O2N5mJPThQm
n2HIRA6iiMOPRQxMYN1HbXX2gLjtlcApJGoxtdx/fO+iRD6Hs/V+of9tjNBHdD+K3kCHPpNsv40K
OFKZH+Cx5+7TfbRwiC+kf7/A3QEdQvHncIcRsDWDT/6cjvoXvQ2jNn0B8Ft3U86svRkIFMlq/YBj
vp3uaPxI3l9ErwXs4qczPhKU4Ig2KftStpSW7bLVqKIZTru0S07Mv61lV9dxFdYwMp1n6STRAn8I
eNHElvfGu9NkzcPrdiEZSCnEuhY4Detb10J0WK/VPo/EGe/7O2sjHvM+W4KD9h4TVSRtdYYQ+uaw
QVKPw6E0GIhu0XNZPJpZ3CkutMwW1cZY2tFcxvgr0LH7fqMTCZY1ZUYhAEOZMbUtZubWjMa0fzKP
RLi+y41uXKkcq87O3ZeIul4s0KzuZGUzClFYGDR69+LP8zFozzZtdLwbyyhCQ8X1lYOflK8nMb9f
0TDATUVB687vKyFnB+i+21mMtIfK2jd1s1XAoC7V5xJ90XkJFipFOQVr08wPFTm4iUTCzsmD3wuQ
OOUkvpkt6kYmgoKyyJyyYwNlOd7z4z19e+TKgTypxisYZe45CkC5LKINRL5LYcUBZhBUg8HU9qRN
q1YI59+VVMVclBE9LWRt3nQd07XuYvC1hEr9Vxn3OTg15PmplK2aM9QO+AvBbg4S4YadGlnFPjYp
CPTBwSHPnGccDawSdtsFvQjT5vny2xWWmkNfUUz+Jka0yaoM2cU1hbKQbp/OzEMwovtDjrHvs9xO
IRd/IeVZ+G28EsuneBxtj6IEdWe5voM9vQluKAY7Tht6z3B31UNWIlUkLKi0SQwHf/2zh37/PFgi
HlT6z8k7I/Zw+EEIXnuswhICVZ9onYhHIS6W+NPtl4N1V1e+D9sX+OAmnjL2UNGUmxEKUal/b+jI
FcY3ggkXzR9WFtzCVUti4UBBXiBiI9AMvTMvN+t73t0F181i55IKwkA0FLoxWR5K+FaF3XmiR+2x
vnAqOCCGlthVXVg8uhUMkZCNc78/kvY3wsvpVy6QhOn+d37CyNau2C8ton2DrjP9VyysnTqp7CjS
N+AYtm9+uuha5LQ/Pl+j2eOKY4mWHHZMVeGjyH73w8lkdaQkv/QDlByPvBPCrRo/ruU5j5gbRyf6
tQmLqx9KW++VP1CeCeo0GKnsvdhWs57eHD6+307O8Hu271CrKp4rexrgwqqwrDrodDdlgXC7xYDV
8eBZlw9bBNeiSwM5boNesUq0KXNT6VJJ+ToJDkPWbc9ozQTvRU1hbjCZdLbTLZjKCgB71nXmmuDH
pP/5O5f6pz7mcZlEM2Q3DOeuvdS/aDbRmMhXwLX0C7OINRiIpQnSlr3HwB7GJOv/mK8LUF1cafCD
Wd7x89VfHIaSEZXRFhAEAnJ9YsK3IGWglyh0g+7NOxxfmZHI3sHttIxbZpt02Q02Y3fMtRyMOeGB
18+f+clK5v6BciZC4AC+1JPUTYfMY87bTiF7UONLvDiVB04veK8woM+WVTBaBK+wzX+b33IsNkc4
P3hsVKg8rRXGvCWh7CK9UOdPnMt9y06ERqUt5VDR1QFFot3J2ADr5s09HNFxfhTub95VdwuK66MA
AnYM0YJSfkGH8djcR340Ks163t2oPpKSu3K1K0oJ69/GUJ5d6KKGkHDdBHCioGEdTKlNIY7BlJIC
77vvSLutJ6XuYIU3cDb3/WXa0u+zSvCY8YF86SMc5AQuWM3NekKvm8zc1NQGzUK7alD4CWWza1/N
9P/FBpwd/HCj2skfDkgDPTmBHrtRsBpMH/pz0ZPnb6264jvgikarFqIbfxOyhRheRYWT2hbKD16b
NXL79ZWziMBAzgWhqKnF571/lOIwKf9i8+C/QowRPKJMB8quzJNeKu3WaDqk8BfgWz/UbVhQgwp7
YZYvj1HeaaN8GowkZn1dhDRCrel354WsvxU+2u60B+v0cDvzewuSALteVGedrG1E+U416A3zLk8u
mKHAQBsE7x2afZPrOvp0agcqRzCF3tFAd+sextpucvOj2CFM8KlgUPqB6fqWsP5TeCnIc99ZO5Zt
WurYkmRw3gma5mAT8AotlbKpRe+0WMUr4ZBCP/kdOhvfLD35whFyVsnFzCl5cr8PjkxC8W70fKid
RRGzFGyldyc1TbP9ZNcOK+T5JrEX+vyrTpZVn/GOjvUQfcuyzDmF6gun42ao8mP22DiKCXLhYixW
RKYWkv90uRet4teoca81XFT9i515SsYV6Pcc3gJejB4NLAnbSZaDgN0cWsLQ7w5KdFqfGCkvvoWA
HyFdmB/dgY6QUBNH0JTNQg/6kGrChuFEdkQOAdzpem5tYoEl47slKSf0VHZRQ9yasNp69hLsUg0H
URLhp0N4UZ25O8AYCZ6crO73boHnHkpgV5aQ3a67hSNgov8PgWncW6038yH0sISAO541x5Sp4Mui
Ilwicg21QqVISSeMuaF13jq6C2QbHmNcCYXbNrVQ1BBQnLZbjIW3kMU1eJQfCEf35Q0bRvrjcKG/
OzQ829K8yIh2c/IRJ1YB/kluNYxAjGNgS5TElP8VMIIOKvNacVWSGgaJnX/7YmtRuHNnEqDYrpVu
P0Ii+Zq9Zlj/Vi/qgyY6TMBU50m+DA1t0QbrCEg9cn0AjkfwKFDQFVy//Uai9khKpVnos2AlImHl
qUKeF/VnsJmrmLo0Sjz78CXeo/LvAX6KPAzAE0kbDqkd8Erz1p5GU5Xm4bLjVX3vPqCkHMtiyKCG
mIpT9O/+LRB2afqFkk88xN+mrGGWIiLhUPx1F0reqImS51M32ubkuGMcuzF87rXkmhyHeuSzki4g
PBGTspdnZ668eFQf/sVHtf7T2W+yVwXuKCyLd4Z4S0LgT3fHYHTwWCtB0EkvMBInT8iirBbhKzuu
Njud3JKdaZqXCYnNPij2PWiv5Mj+An4BrFcOFE+cZZoMCCXh1CvZ16q6Vu2b56DrFxOlyTB1cn6N
Eyy5HGjQVw86/2/6Jx1eGVEgcyAQR+YbCNAADwFBMuTbK16/b9CMnObtUXY+bihMvtJhrPNoWof+
xus8et/3Q0Fa2O3jF6J7esO1h3G2Lmg5yvFgB/ZD++K0/PrUPI5WUXs67rHqJlu5RWeTDXONLSR6
cM02YfS8RMs2E2OpuKotLyGvYQFL6aFRUbZzmWddeeIDb/On9SU6hEG/hr0Q2z51rA2UQNY4dVJu
uiG0ul7NWI6pkF9kc/edETX4eBnXHZ/vRbcNUdT0205EyXUs04xGouiiywNpfAgsc2PjmTWWwsHE
OqUpqkxXfTOcrR0F+/7VwdgjyijvaS6P/sHz4KkqWpAnu8aGuJJydj2TcoIipeVXOD/CAcdCIjlp
7hjyI/J5yDJkAK8HQ3kibL3RRatzd2W7X/F/pTNIItjQqNtHgctOa0g2VAw0TosIZCdPfSOTmF9t
nC6G6GUsm4kK2F4AxQlHdBz1n81DqwBLIzHCVyVFyemQdr95xQEV3qpEWu0XnbQpH+W+k9B6VAbF
XOGfQnGIThd1YhOwPDVPgicAnJTcmUg67cgO1bLJTFEecNij/7r0hSukeg6lyuTQXDR2wO66stVZ
G16jqDkm5L0tqiLD951FY62sMZKO7M0AUE7XPeH/fGrmTpZkAXwihDVL9jyk1tQgoklxvXb3wYNh
K2RECL1b9lg2bRbFo4ApuyYTJSPGzBx6WI2MI0N1URvFw0KzYbXCIwvbwAwYHlNm25cMaqZsRKv9
/Kq87XQCaNHlTq/efMUWwPrKDuBohaqfcknWS+qa8q8Gl2haWP0meBWY85LV7BhZnrvaECdGx2EA
eck+sE3xvkGhJIrnHj4DF8JiAUxaSZnVgug51AXyw9AcQtuwp2KHxUc2JhJ/cLzbELZ47SGSPQ3Z
UUdGLFoxbs5mr5OCrU7SohpFyL0NRY0nTiInpp+2Jv0svLKH1ddtp1SEOTcRe7YnXiagBld0hRYv
cME9clGTHGstHQNbH7GTiP+8nbg7qQi0ZTvKo8u5R+MzOeHBNPANkYvcC3NJHOew+2GmdFep8SWw
ZGtkXJ1pPagFNl0IVkiGUzYt+lW5kSbXz15bsy5EuDhmvX9XARNotw8UROAlzak83qcLttTD3acT
FqmKTPycdvk7sPKR6Ggz/HbejIg2/m83kDYjnw8KZ89H2aPBwp67z9nu4E5MB2zMharxaEjI3AA7
dmQis40x/FHzDZdbd+EQmbYVfRpfkbDnPtHWnK/o+WU7cNWXi8QBQ7u9hw/kAW7oZoEg0PEJPZVt
mG3faWPYRbTSEW76f662+XUTcaCQ1mJYpVV0cpcX/jKgh+6/oV/+AlkpokrlhvpiWBx0tIQKrExq
anj3KbTB6I0AM6lxKJ6wOZxr9WL7/XKZ42dlzmhW2AVgtc0ZvCwMoSY92kjO1pTkXvpXg434OXB8
ja2S+r+CZydAgl6Jx6eg0LZongyVBRnnotuIm+LJts7P40AQXVTTsbV0AykSbqsu5IURay6w9TxQ
spwCBAQk3WR0FNZgaoKiaQt6idXqyqAeOuQVNis2Qm7dUURo5RNVY5wZY6caceaFJkxP5opHt8WO
YcfdS0iXOvPPGZcO3kOHU+CEBh/0yzvd2izFRPPbVfaN1CvZY0LFGmClKa54GKbKgpLFouM+dLje
puGXzSFEfPnmqr6z1OCohSXWqlutPEY5xas3GysKTPR3BZ3DtEixcxTbXSizbRH74nwhXFsvP/aN
+zDRbcQLMSd/a1fBwFF6HNI1kQ5llapQavKaGyHtUAlJrjaZPkry/QF/+yvjflOAlXerpgM7Np6G
fU9/tBeW5Dn0niq+tWCPlDmv+0PJjShKwwXY+kBd0FvhrIMHJTMIgv36Kv7o/cIBdUNlAZ1fxf/p
BhZS7BpbrGAKwhvoheISYoe0r7f1HAKsVfYKKWBhJf8c5tBkRb1kkt8HQchZcsPyt30Nh5OfwTea
ZzfwB1eAG3j76bFHIQM3P7IoRUVj7SgqTYq8K9mNvPJWRWyZjer6xWojlU7ULMBUS9uxQdbOm2XB
HV5DkrUuok/zwunByOOXxwB5DXJbDwh07XwstdddYfMD/qAjp8tSL6A1cWWSFSzX4SxocU5XlQMM
0NPEnvnmkxowSk0ErIUTLZXh2+csT12minbua9fmZhQUuxDJFe3hkN0SNP8fqMbbxeJjDlEitbJJ
lKsHwimaCklc8VUy9PX5JykMRUoBEE0RN1rPIFdxTyxNKmfqCyfidqWbuOUkJ84cijvhfBLuBSiX
Dl1Y6tDXD8CXPtytOkR9qSUuJNCS6iLoKRAEBFgSorSMudOg7HW0HzIDPgNUe7Y7YgC3xeJK8clJ
eEXfRjt2D7s/Zf9LP+s2ihFN9IA8cPhEbTjviGsefaIlm1ZqtU2JdgaVw/PBK24/i+hEEdFQ8mxR
M2Yreluv1SYIGoxKg6qtLaKyx8MSq8IJk6kE3YyFz35q13bx3BFdAUGCt7T3LQ1moeTZj0P7oy/4
Ov4U6B3Mfg+Lb9aPNgQQxvz42dmfhNVF+ti5wFm0u0+kHKxHBzEBgQbqM2WGu7+Nevn5jMbwlAqe
kB0Ve/hedRoMY8ITk3q/9R6XQaunqKkIwGWLiWwL7dMA6pPn5/8Cq4qEdlem332ieEmUvYHsQ48F
NiKO6LmUTMwTBW5O+dZaPENAwss4OLjAfe92pDTXbwKTpPx8mHfT5n/KBcdlBJWhkpsKGhvtvsUS
MwoP3r3+YDVxQ0e6ueu+cLtyNwTHoDpm2Wyd+1COMeQaMUhfFvcb/NnCnjalUP5fevg6CqVY8vP+
ZiEweeilBYOGzeNAVYP7hPqmhIggCj1FEZ0O/SqX3QBQIhOl+i1zT3WG4XrPfR1Px57IDuwyCzSr
Ti8/+RQnuv4OdsM8UnO0lTZdn8PNAMFrb7Jg0ne08eBZHAFZkDknOaFzApOLsfsrUw0bX2UCX7wS
h4PDz4qPqzdklP1JMQhuHNkjbahLxpSkrcUrvKIKdK+F0Myc9Ni+AkG+6IttZJVcAfnbj8co+itm
kVGYC6KUr6DDW4awWJjJ1hZzTJPrapzWlDY5LpVJYUTz1Vs1ZZ+spwa/ERijqVPk9vaI1Bk3jmH8
8AXmzx4pSzg+XwHIlbK4ArU9Sn/PtBhqw9s+6SycQ4ol5PRk/VuWI0/P1oVr1x/cH/E/884phZvK
Pa0X21wV2xfjViaFiA0R3SGx0UQ8ZSgh/7p4qqCelQEhUXT07Za+XOgGi2L4bA4q2oDi5aL8zZuL
bei4lkJHvFDetoV3wa3rj0did1ls7jV+2TCqmb/Io6hRdT/UyqRBFqEIrKZ62USp3ZAk87PIcnzH
c8KMru0EBRN0ZREYQ0y1ErPSySBZ6jHfzZcG+Cvp+ZnR7C8QSpXSjNnohGdIGjYHgYJMosIlAOS2
tPhzzybXIbH0qx/y3o6EdRA8+buaJxa+BYEAbc9B2I0k1gIREZLkkzvh0OTCXR7COhbmzJIBqmm9
aoZmKrSKYL6FX1VUd8CGDq9pizF//4eHA/+5d0DtCjU1tdBTAyvU6U4qiQDbRtMnRJ7jyGR5ZCpC
vg8QmvNYiJixaqrCueS+qQ6ufgVwpBOllo01Kpj1zCiHivsZrYYkbABTLTOCxGvUAApBvYoY8piV
b55XZgCwgkMCkqBkIjPHFh8zRF/A9XpQa/Lsbzk+jPZayWB4zuBj2Ij/2gnqOgaVZOekYc5qm9ie
EJKWwbwLirVW3sHGbalC7xvTbd28r8iNtMlNSgCqD9uuxZLumdPIQE9OwsyGskbPB0laAG9mPmw6
E72CXi2hIIEInTxcPi4rlwZu13S3eBmCUBGs9Y0sKQRxY4UhVX9uO7IoSjqT8209a4mEwVASkAKE
bXSJokQrdBQs/19gWAfR1XtDi1gR4+p1oqNwkSCxNtDNanPzbF+RAq9s6mK9K0tH5iaRLBrU4le3
lMwDDgaqSkErTlLrMGONO9yC7bh6RAQAZm9zwQHQYy5F3tTaUPa4c/G20z4EIq6BOj34aV4Hbcar
lU0I5/GrKRPrJqZHyzK83Yl4OQ+mL+KagqAKGpoUxPrsd0/ytdArSrpo1Zr3oE4zT1oDh8CeEOBD
6nOjrLxR+He3zMwCNPyDIv6MuU42ENCLbOCUNKW5/PDVtFyreNQw4ONiM1HU8xsfbMAzzhCk3J69
Vs27jOJa0B9aE37A6ae52XPycImbmUr3ZCrJ9d01FC6JNIwN+26D2ZeIuZ5WCq4ty91zJAUSj8pz
2wbTEi0IpbxgUgWkckyV0ND21kJ2kyuIP/8kw2MUeTLhFFRRHnJ1dGcahlEgaoih7lXh5G4yzFmG
INXBVqKZbrxazP9MrAQLfaqtRuqOUJVZwgfpAaubGZH/eu/p42/z4srmLWekJeaPFK98JehCS/R4
dBDqSV55DxezcKfsw11eJy+y1D/W3U+piq9e0zNjUxGscTCJSQ06DDUGnzgglRhLYywlUJsvYleE
0ra9Z2Q9T7AMmprMWIXesYM5pizTwU/yG8mcp2Q2+w/rpxJrspVxM4kk4ic9z3FOuLDLkWelGLh+
4bkCXEz7+vqxHvLEOFSSvzXn6LhGefsuVpCvdvc751zeHoZoENCkqHM6SWsqOYfYCQGlnZUlqHGD
TDKrIt48FloU7QOb0Gb6k2jruW7DxQf+8pKB9Ma+eLz14Ohj4jR2p7QQ8oFSXEvpLh+Dw4d6tsMf
e6RvLqxbnw5ey/T/rn4zaAbld9V4Y5xJZ2yrTAfySPjF8WgdH96E0vdYva/fYsrZOlKwKFUbpU/l
H42HbNqP+PrnJpJV+V3b/bbHHCVbeIYPh2pSd/asK31dPk25zyxqiUxjOVrnT3o3gfSWGND0Cufn
06G/CaCBCYEfrv5H74wULFoji80ozimQP4q3DwtEZxIuvwdGFb1XL7FosG3yvC220ngar+/xnq8d
pVf942q5YubcGwoVw57VxPTQdEyPwC7R3E7FOMGt19+SkAvNwuWImqDWPLO0StThpp+3K51BnAYK
eMoJ9dK/XzMEk6GOmG8y/85tCOFSIqZbIOIFAuqP0bOSaopWAIfIcppM2B/Bbhjif5SNzzF3nhPT
3EXyZnFXmPoqDHgzJcV0+OZdNddgArS4prKTQia2r09Q9vG6PVL0BsoVmC4GebAxqvBKB3eHQxJY
mtzlSjOKU5N55bsBh0ytAuEHbPo5wnOcfc3mqMMtwB9X1+VSoBwWnw5HxfNml0vPKDDObXso4GCw
OQj/pgjTI5OoowszBXwRh5sEiUU45QWoXg142OeGx0DKenlkXFfIfOz5TF5Kxb19u1+XsBbwL68v
xTsW51ObDBmsX8AnIR+GcdRos/jANQzfmg/kb5m5MCjkSoKADM+G+iy2zVCj5QyHGIW5NYL6/2aB
FZyiFnb73SrS6kfwkcT8rCqDm0K9u2I1PKFgsqG2VZnAwTQRc4+15wm8D7P9+pUpFNEOVKoNihgx
2qffuGt/hIxcv+Usp/vOv3L2AALudkcepNp3fOhEt6xASc5QpcBqXn2uSs5pH+2AWwJ7f5w2Tcxu
atNNW1ttZNLXP61WdQ4fK8J7TbOlgFsqpFDVpZEEtu9aanwT4j3RL9ROqZIiHdShHjbaECH5RNWA
MHZ8azZnc7J53rJrh+W54+DtUNa0zh2pysvtY25h99Tu4KXs3bFQlICX8CoMHE4j4fJS/NqHj6II
pxCPwvkRImzDRyqdETkqac6KZ2OSW6XPWzz8L3G+rl1LMP0GBv0RbFf8fW6fnzg1D0UY4KToAN4s
gkIFBdbGSH5QEe4+1JHalv31/JvJ6y13bh4Uj+1TbD97fxMALkryQ543RyRJb9erjVzsKhP/94xA
zONu85GFGFrqgCynYeJZwSY7gksTP2/6NxULBBhHNGebZbnco3TUw4ZpqUxKo6uYu4NkjDqXOYT3
XXitAqYMsjXi4AcsddQ4UEvcalxtCF89wIuDfSlCbgvtE35HbytmDIweJHFLHViHM3TDKh9QjjKy
mr4qapheHSk03pFk7YRTf1ybb+mEDLiqDC3qmZXfJ50ASANFiSOsBbiI06bjw2Q9dpeCg+l1LLkI
C2XhHAAOvuVshA14QKEmojmMEKsVId8x9AqM8Xl5h2kWwbTXKhGFfL3SstaZktsfTDNi2SyWNsei
y3G/ifMhtK0ry02kLG/1tb04fUXaSM4Tvk7nTGLZX8hI3Eo1ZUEIJnV6aqcRbX0rCs8PYGLh9bub
uYJ4M7i/ySMiaykomXR1Z7CYB1VPZBs+Q1nmgS1SSomEQIhLY+Wg5wfj+aUmSKxJhIhQBQUzSto2
D3Xr1ArlwCt8HQP4lKKyMT1ou6qEaElA31X9F2TxvNmQp9rcvIQPEZciJdK5bDdQAIL0ZTnYi55q
WiQYYApl2q0i2xhrY1G3eW788Rrv5Dw2Mg4YwenlzlCa+4BqK3hagXaHuT62avlXG/O07/RgYr5A
au02zvV4mf0gvmodrAU8pm7IjAxOU6EIe//Vv4O6VSgueYJyW3QtzrW92vXOZgMIkEuar7x70Qxf
+6QM+bjHfx0WHlCg7yzcYoHumvLzwdgIkUligw7j0x3tAM+BpcXGFQOLgTrFlzC4o/TwvcMHgCdj
TpHLXP/tDHpmQj3dQ5zm269+kwZQZpEvxvt6dNYpP4a6Gqa8j3mQ/6SBVdVXbZDermHV4gYyCPN3
gYyCnR5fLSn2WIO7zdEbZ/pJ2k4wnKUpOVbCyH2sYmMl8/NjXJmyOLWq4TXS9pROWcc6EN8tqh7N
IMCqe+mabQ5gzdk4ZY0JSb5miibjTt7aSpp6m3U1zWPy67/le5VpluNemZ9BcYaVHxYRghh/LPRg
Cw5wgLEbUQfarxMJsbzlIT3s2gjbHiCb20/g8/Lktw0Q17dGA5FTuJbFQtqE5VHabGgO/xXOM25v
qJ+du9iiZjwq3+T+E+CjnHk0fVmGxOeQZqjhvXjYbBLnM/ddZtvAgGGYVAMlyyDsBCXIwYUA/ThZ
13I/O533sqFlke8jNt6DsbMxb9EeCJbkJF925Vpy4YnuB6FC70GWTI5SeNX42ACIIRDlplDzSEmS
PmoJTWX2iz3x95tZ4Inpcgr1Cb6Zd7GuNFOq+y9xlFI3qMnc5+CNJix7z4j6hhhggO/3855jizKO
Ym17iOs6mlv6Ozr/El08vC3Qf1sulJCELbSfPtZB5C4xDJxPtaWDho3Uoj18pV9t7lcymhec+GPR
Vj93LBFBNzjl7akYysgowVHfGckNW1n0PhKeC7OsNuuDVdiqie38sYL2eV69VMgnmRs2dTyAEzES
AnTUt3fNexSRkMh9v3/FdC+DPC4HhoXXuh60z9e8mPrexIFDK5zepeneJk+aiCD6YhS1LtMydS8v
G/JHQpJjxtaMYybY++3Z5SMxZQCOMvZGe/MUNH4npd1aUtL9f9iRnj+LtqxzpsKphh+Y6IAA7y1W
5U7i1q6q9v7pgsAfUw8NwHuZSuKrZNTrnDQX0fBrxS8pd92sqVTP48NBV75tsnrInPEJULgigkAT
cVftVvdK6k/2sSQwBgKDx2B9k9hDQRgsmgs9OeZIO4sxE2rCFs888BF0oTh9wf83yAtmdFYZi0Rn
sM5uQ2yBxln1d7Sd3y3YkCPIXnppR6AJPZLfhr66aQ9LQ3XxDPm34znf4MFclrq191NIfWT/pVZ0
2PdZYhO6Y21T2/m+ZScMp/E6P1KjQNWMUzB6PqLyyYkmg5L/6mOFw9V8qtNO0CJwcBXkObezJdv2
YG27YgAVJ3TARV+ulNPMR/0LHF8MSKjFKPwqgM+nY5R3nlGjg5Y+56c+/HE3QUUJD6SyI3IbgIab
bO+BtJNQqhfp/wSo1LBlpuv/Nq7GGsEUrnC7Zk3FFC8Wnjj03kXPBS+bxb893/93l+0+nOJUuqCi
jZJFuBkXwMKKovkDGXx8JjPkHo+gIBMkyAbby8crbud+4rtPkj64bhAibOV7afhB97ZDNvofSEY/
M7Ymwf2SCdimrZw0C7KdiXcEqNWVB9aNMLoRExgA4F6zAtv6eaMP8aDWC5ojpy1sxgVtYrWbQnle
nVX7f72/N6cxilUvX4PYD5x0oxfFno6Q5FpTKw3LGM4ZfecOUT92jHqgdMbzNTk7hJUre5dyCojx
fUInlHhSr9NRqBEB2UwNP2KKhKVLYO7gRzvIWxfc0VvDPryGmma1jQxMR7yzrsexeMW/IJmcjjs/
TQJf0hCX2NZufAiMByjphJVEZUmR1DKZiwbL2N1rzG9XcSAxCSX/kcNQqh+BX3iu2rIu7axj233I
9l3s1HcC+JOYWVycn/lTXatjex0vWe7C8//YhDFXHH1/zvcis7+XGdqhrGKSYid0keEqvFSQnzOM
B7E0rBSb4+DnlTysnqO/Zvxk2zpPge7q8c/n9Biyd+RCp0MjW3PJXqFW3v0Zum+p/IGBK2nBThCQ
I7r0d70X8ci8WsCVcLcE3qxsfEDYma4rSdLYeii4RHJn4/ErSntb2Xk+I6VZoqzaGrnNPiVbsVHP
K6Hl8Uh/4J3W8Gft2pQD4+T/LXvUNeWbbD2qEIeoNM451sDfAG1GZxK5unSGue7U1WRN3Kuw1FRV
vqfbdJlOZ4I/0TpCui3rGTpbXivH6ep2ciGiV9ExIvuklwHjy/aD5nvJh6x2mmq5ZP4khUe/Iv5M
QJ4Edos4ycpZYGuhLb2WnliHCbx+dMnki0X18inuQkpRYCp2bESfdquJx/1qLbFY/a8rxqKtb/4J
9zOA965Lk2KlxEq9EscFw8a8wHDsDUF6pa9gxM17SLZLvZIpdOheaeTDRnOnGQG4ykaZV29tXVrB
1fT3QmuUGuj4EE2ACZzYxwcmeUi315GMnau3KoqdEFo6hatLRGBn2MbWe/+ecjbZXpr9370cHZ4q
YKEgmgNjX19DRKJIZEkUBOZjw9L0o1L3DvNkpMTT9WuvM7aCyFJEAVSAMsJCknTYb7szLEeU8HJB
te9xyP5xmqhieixJzhinO9fVT22j8vefVZxToRxn6s6+CydT7l+jUWPWpu2MemyRxY1/YXy+GCmx
XDn4TsGKga0RcnZRE7adhy7sxkKqQPHpuY8QOmvq31115cxSfj/MVOpOxepoKYAsTsDIM7Yde6L2
COkDYAXg6Ace8kS+MEGNt3rOW3pBQABbwNJdTHquaZ+HZLS4XYWf+6E7ksURSbbqxKRh9Ne8VZIQ
CD0XYOMlQtp9u0nHJEXx+Tw0lCRw4uhnsbGkG0VLg1uukhUMoKeIx4tQPyOgLKSbOZytE41ux8j6
QWMYjunMaExv/whxx2TnpEZKDL8QNRW7QTVLM0hbaaDUUabTFFOIXdQyBUYIUGTFXOeKJ1cL8nAK
gueDPXgxgeGZgEaz/wO7qzYJbzzdPlVNNTixWm+Wztm3cT7MsjDE/sCCPxyZ/Nm0p11vaNQa5kpX
7N89ydY1soE92761gSv6iT+8EwtZ5tXqHluq5oABVzFRV7fAnu7D/o4uA86B3b0045je4PDRrwji
Pv+UTt9SFxaJZbtH+FdOgKAooMm6XhjNrmTe9wGG05KucfD0B0SO7FmAcC/dWcJfUJmuhRLdSQm6
iLTAqvU5MLK+zQKKhL85BqsLcgTAZPTyVNCJyPI9DzTMuMg/wI3XNxrwVOWsDa6miYQaAgF9Wi8N
ujcK2otFz/ZZvyD8Rjsbgm16YuDHuDhdAdVptgGQyknNb1Temw6pae3c8P6J8W/naop5ATwi9h2k
YISvaLf0QNfKpOa4J+DrNiy59ILfYug6WXF+CpJ71Cr42kMvaZ2DljirqLjGDlYWnHeKIyZNPZIy
FmrB5aGrFHKipuabIknsD/o2w6geL8Q7dLMCxrm7Nj2YGm9N8axTwyDvjWuregZBYGy1Lh/8g4js
2WKdqGjsyOhJPhqlqpQu4yU4W+/Coweddwxzy08kOHamm1j20dOuGsEZTPvO3T9pBs18KyxA2sYr
bb7AP+qsqPSf4ElRHjQg7NR2HepbUeMk2TvuDHiB4yIQcm8ME/H/VXfXYTsiNSU6zTQslaKmSCS4
v3aYuOcuFWh8tizMlrQ6gQFQf6MnXl7qczGOVc68aI9/tHC6jx9lFXFBL6uvJ3G/mbo8ySYXpamZ
7KL7Dt4TyNp2ckhvMipTntT89Y2V/dF5Y0BSk9qbP/8v2tQzzmrH8DRul7/i8m5xOyVfoFOyA7Ns
F0z6DtcyQ5+MA+m8kOWI/4JLBjvcWQCkS58W8u6xQ4wT3Jzb4zaVcjRcVuc59CTVuHlrTA9xWsBN
j75cThgOWpx/H24WhkMg0abw6Y+fFhDrtcv+jR8zxIf0IJIsKlq7QewLAfcCGOYD0PrPKz6uciFu
GiZ1hYDSdt0TfiAIyHVukXwMuxCL+mebgOC0MVfo1mGj1tYZVkO4g0H51csBuwxhlDmOzm6kmuBQ
G1sMPj6bfAqrVyhwhQQfxNaxQSHGmwxWJxsmDz6QzGmAUcWmQHs2Uud3HUnIkZiXvZUpeXvGix5b
h2wl1UI3euRtyai4nuYcVphMcqTpRByJlS0rgzczVzsiwyKn72QyFcKZZzEZj1bFhINrvlZ5ZMTi
jnTcViM3pDvLdMtizgIBzAAhP4ahdijqJSNG47NMs8IFT9YxFUyKHKj6+vl5skrZ14S013W01vZD
+0xVMb8li4n77B7wf+vIw8MBjt57w0gF3krot0/9kuJTXI3CBHxKFNJg45awQO3jjB/PVThfMFeY
LgToJpT1aAhqChwZdSmCyd/G1Bgzh9JUYXHUoCjADOtLi9Kd6C3eZ7Mh0wERTJnY1J0GvezBaGUh
NX12XfplWiFfnXUkZC+iVbU3IIynzVPM5PkikIB7rz4c3Tta1F4Kvd0RwOipo3wV12v4Jwt2AQlN
jXQI8zOOD6rpdiIVFtYLFFInOZCuAkcSoNExfAqpLjxTOFKwgWzuuy9vjM/7A8rFCzSb0Ggeni+w
gZPaoTIoLqeqHAxjsenWskAt9sLmmH7UODYdgaVX+dQ9bKv9YbZCibB4AQ5YBh0bqLZtQQgZoAtW
hQE5azo1xknT8ysqL3fiQyzY/OFQzOhCJf2bG2c8hC5oVPq4BHUAcHHFfQnbEtjnUylDQ/dQ/cdv
LVMCzTakPx7h/c7mINfVMacMCYRyjwzhYIKrxFv71svXe28BatzutD7mRzCgXsWy3ngnZm/T/jf6
moQ+soJEOCpHgBq4Hl2uNgmk5jPyzl7a9Q8s125OBPOR18xGZWoFZXW963fv1RQMibAdWL8ig/nz
62sm3ZO5a3FWQFgD5EPez+G+W26o6POvlWpJAYdVni8JRO1aaRI5qgH9l4z7LR9Sw8uSHLNLdpM1
FssZkleyop5bbU95Ofw18z4y6O/WZdd5wRBaS8rxc5YfSK13mkEVLcKQs+okK4MgFnPll37x0oVe
IgE8KqHBchpXEvMapY/SwVbjtM7cQ2ry00E/umgLpzkK2Ebkr5TikKgCwXrEgNUj/M0eh0CJ8u8X
uDD8t6QM20IJObfRoYLJ3MOLgl0YSmQccphE3WDwBy3opxOCxKoYg6Q7tHwr+PllTlWwWbfW2e+S
2lHs0ks0JXWgfQrQBNgi+Ku4Zg/H+uRK68tpW/tTaf5WILy4fgFx+xO3UviIiz/9LDBq9A2MY04i
0/uZM5lzPPiGBfU3a4pAh8Naapwk0m3YgREhqBFFFOvSYS/77A//ovFIN5O1IUJ5q+Cj8PCi/SGA
4mayCJFeIQFrfgde+WGhTcKIvPLCkr2nEgN1hF/YUaeorKowJyrh7ZfcM3V07xQPEgqdACe/I4Ql
IHk8IuGtUxKFI5ZWHtaxHD2Q4G4irZf/6DcKKqzBtiZYZLeJqnkTV4x7uggl5yd4XCOTK0U6EmwX
gQvj0xE7e8xN+2zZdbmReCKBeoS4nAuPGIluaVB9swDuYn+x+1QCGgW0AR23qDV02PPfrIEEUqM6
pslFn5OScAw0FwypeHyewF4lagsgXQDAyFcnGVcPgwhdrkAhZeT9z8tKgm/8sE3tLipbJzohsUSp
rHajxo1hkiMik4V80EExCCEJkXOOC/W/ucIM6L86ueDekHO4zBCSfEnVii0AzJ5STiWBiypPm2KM
s2d0ojI3DsjLbLnpB5eptFYFtTI4YMlJT5MQsJZRF9sEr+wnObU9jZeDTpIlJ8qUo4PaWND+8/Ig
6zfPoTFaIqv6PzIqW6eakjOQy4pacMbxJYV/lt6yfxTbxYTQRuV9PPzIYyWJN60Jm4WcSEIHCqhA
bx7xyeh/W2jiPoBEWLqF+BVxnu4c+pigj81SLdy/PXcDdkrp5yM4zW7BqEfeowGpJmWWnvy0UFA5
+G5HTFjFf7z/bbGbRs0g4yXn5dEEjqP7TgsjjtrtC91k9sorxAxLkNCV/2g1m3U6Rw1atiVQF75x
0Dld8EP+BkKRz0ujCSl7xJ134Z+OPCSmE6hjOUYewAXMH5d6aUyf/zKJwCeQj5xyPcVSwiJf69eK
5hPurHisdTfxtgcGaznRgBCOpVO+t7+GPxkY7inSMAKMpXfvmOpiSM1ItefaSwtPUC/wgT2k3rEs
vwVLLGEO5gkANY3cnU/kehhyfET2sMroTWQgY1WAusSsFu/nWgG7UE0D+mPt5c39RE6ztJhyXK9d
aLRVgQIhJXZQCKtYXPw5BAbrrxPewLU3S+hufgXPaKEDKPmca9Nr2kK2lkrdhrAVW6FHKV+vu1YZ
PVwV8y+MoOzRjk7r+f+ZQuOJskUllkJLLcglKMCbZtT3e1Sg3JBv9CX5JyRwQYQ+AJ8ZXeXsvRcq
HNlcR963is53GXEhODkcuTT40JyCD/eun6dMm/vvSewok6j450lzz7Vqx31WTbflbRk6bUD7Vjdk
VpZ2sopUSZpTcOZqVaQ/7tVPt5XQSGHS17OHIt9IIWA0BeyLNWzwGp2UlCJAnszn59B2a2fKb4Lz
D+tuBvCsf3fmw1s7cPm08G4d5+9ixoltCZMwYzHPB+PYrIFPIEGF8egE2UW3+ekJuoYKBKqH96j6
i+zyBZ6b0gEITFjhpu4OlfuFYT2vYPptyYYbY92iiq38Jw+Q5G2rtSnJh5wm33qkA4GGA2sUPX7i
hIfVTy1FPOkg8UGBoqAm6I/2ZysBNubxo4NRRg2locAgTk3e0JxKFq89M0ESqM8HGzfrEYmpkNGt
zvNTxAnYM6+/3/Xt6/feAFb5+J0nXWapYN8vXAWM88+/eJq5BdxjbEPmDIZrFOILqWxPavoooSPM
7MV7Pu52e5d6n5WAs9FefkrXJDXv2BvjhdluyP9ihJ5X7uJHIgOwHn8yR/QnL3gDaiQFPLXb1hRf
zGnxOmoUVJXuHEJE1vSKcPlweTOYQXRPEsYv0bLrxJDp/KbvGL/l0RTde7sBYlPnGWOR3hRSySXW
Uw7rQSc21cPzHEjv5RfHjtNLcf4NoB+hs0jNAfRTtpngVY2vZ53WzXQQ8txbeoZKRb2IEygA/xed
TStnjjLbLD0fuWGtlFnJes4z5tPCWse+2qtxKKGTfCBKC+9J/kniZN9udhiD6o6Xsk5trdyrXoA4
dO57tki1h8vHFr2vyje5vdwQV4XKrHakzdgBC22GbK2oCTBGDYokuG+TkKgtSospyAJMGHevMU0U
VxRIeGmC9/iqe9uqSrAGQvWWQQtby2c4NLfPuBlFIRyMxY1TBa/20l9CIqDKrzfoL8uGT/f9jEj7
tyjF682huKCRt5Ri8PBPHv0N0PfHGli7Dl35K36vTKqHRw5GIEcR/3PB9jQGvqLqBBDHv0roWU6g
CddGpwOEl090bmctwHz2ddbKFmxTWloIiQ0zxGkv+Lq9lkuo+jesiiPpGRPPoSEizTDpeFWyfb+d
/9WQA4Si3nKpS66Tkw1ZF2jaWCzkFK9wJdFDwTxWHH1FWSaA3e+SaDbB0iH5iiulZkFYs4OiK0PG
xxQYP76AryDDIEAJsPfE0oit95+N6DG0KBvUfizl7j+2ufKYL2+xMGoaVeU5JJiShqa0hDC9QGzR
em7fLQ/Ibj1Qi5ncgxdUthJTk4ShxZIwSMo0ALoA632C1q2zkhAkEmUdPnUW3i4pWxHClnotV/HU
vNTb1me0WUKkvxuujO1ag8Zmxsm2dTwA0TVdllvUbKRdNq5/CLxGfXxWL4n4mqXQhmyTjGvposfa
qlX3e58K2poQbaYesNJVLSWxwdrcKkNhaSqEzMjIUIcMPgloBghLPtkDvmP3NhtOMxqE9z5jwkwZ
C0L+hy9gyh8qgSZIzWbgGfiQhPHcnhwcoH5g323W7ApTLWwWRx3qpUP0RoITZo7WhLKSTJhhkivI
HdMDNvQyYjFbOsQptE3cAIFO6z3A6Zu/rzmW5s8zfGDbvfY+8MzSTkebD4XyE7+wUFto9iLjQnkp
Lq1ddkmZEyHJdbFFtjP0wxjbPN/76le230TUeVdB5WVfBT+s7EPEEZKVVXUPI/qQ4MXS7cc30chM
WKQyLLVn3bm5jJJqJy9+l4tlgPDawk8dPaYwAtpWf825S1Xj2x5y6NkYK2+GjUiexqbXB7l7YlTL
muaW+kykYN7e/NVP4YNiK92AjCdUvdOeSFpbvBA5E40mY18pMScEc9PabKZ2bzElglMQcHS9Ynls
UWd5hbvLrdhLxLm59M4tNai1ElU848TnrlZacKoPz4ILNJ1o5bW0kYQ6vii/2SAOmBClCeYSl6LG
G3AHp531cUawYJ1pwOvRLZEW6nbsqZbNMPtS/1pJj8+Xsi1nXUTFz/uzHH0OSOUNQmu6/0j8yCIn
361bvSUHIescpwaOMKpX0NR9poLIR4t+2zJR9eaCtdJughae4GzX3aIalCeD4s5R7pILXvFioM+r
CBeUP9M9AI2Se3zvNKQ+44NhyPY3pVreZ4yk+Johq2uGGcmkStYjTNlWnpmdepv+CKzgdiJFj67i
SayM/7GpLwsXRrOADW4SAIfcmM7T+JTu/V3WkhrgFoPVF0cnNgl3KunXs1uj1u2qq+YlxsmCWeuV
jsC255LWykY//js5gHfj+/nEGI14rZU3MSfUEhloReRegLLrYZCeiUO77BUo8xQBNeqsptzQRxwS
borMxEJP7EmfDsqIHicxMHkN6ebIRPjNx3+6lJQSA/m6E2AsiOJ9KyBWJsEELPAl/F48kCEoTisH
0ScYupTR2huN+/lyLHCg7BlVwT1W4Hmmgl0s5K+ZDao83ln/mvTRPcRPvGDC63qdBT+Y5yI3V9tz
nkWJy6631eEF31sCFJp3jej2w4STtMrJUxzGI0k6hSCqv6RhO9f5LXCGDzbQyNC5OP+Cel+oiIjX
U6vuwIOD8LApbdllPX4tBJ1lnU8xWZ0kkPRWhPQ1ubIaRyIH4UKpRxizN6hF/NJGcbb2iaSM6YYs
u0FzrvwthDu60qYOGtubVN58yGjUfE83/gp/pPfNTP0cCzG5hPACLP9YCDJDHpnAIrPzPGIJAwHV
tXvsq9BAV+xkFYu7+DFD0omrAf+yJc2ZCUg6bPR4Ka+DJqYXCt+717CXxNrPcOThzmKOn2qX3iZm
hHlEYcYazlH5u5n4/JL7O8LazAYVgDC96oNnlIl7IbqvV+oS4sVsj9YIXwZfHt5p/uGe1XI1DkgT
Q3PkfC3RKSrStbac0o1Uaztwb8lplJfMoc6VgruJQk+Rzg56c0ifL0sYyJ4U2163CCmtp5GzMerz
9p9ZKuzm996z3TgRe/0C1sMFLkWexICvmDeaPnDeWY2tdXREd3c3vVOP5unKTf1AsxA6g/qzZ+No
wKo0vED5EyYRvQusXtcWWGbacyPXO99WN1O+iBPR3HRwkTG4UZt9g+CH2rwrF0ISG+dlEitCDkZZ
sTi5qjZibBXkuqNKcgYo8j8YmsYZStDiOdO2xpSB7u0slRo9EG/qI99SrTIeA2PEM2U8TRv+BqE1
N7h7y3p8x/1+/qp8llOTQwdZrCClyEU4zcvzoIxSraQOIqj5x086nsBNiMJTFx8ks1ROnE9U2nQj
ZB5qMAVpGr7skLQZDLWqq2fetdI5a31r5rHTJeUXm0ybAGQVwQqt7LNH58qXba46GQ/3xY+RcoXj
qvTGe76M1ZgBa08/Wf+AOgQT182HHlJ7lQgAzP64elSFpI/TBUarSVlCuYXbnZKR2UFf5ySEt7gD
Yy77ykCx3tE2WqNXYNplS/enICuXOpb5xG2yJ/aXvljIY3/V3ZIJ4NvV8sEFtw2NJR86ZIt25shV
dk/EKoJdhPI5SpRiOa9Lx20/YQ97t4QpTWTXVyEJvfBhFQ4i51+SyRHZViUvvpPe1lS4hwXwTCEk
9eeC+b9QWk5FN7wDuu5SVTv5wJC3Nke9ZR+iVxp6RJMQcsrHS5teM12iNi39pX/lDijCXWiTyZ6Z
XDpG37fy+Z48wvCamlyCYUKfPko5byuvuwndnsV4m+GX9bXmJYUXxcQcOj4sCNROgz/UByCQHLay
Whi35n8hAmxBdNvtRT8/6+m9L8fDtIt+MvVaxMMo0ypbWZdGneyj2Jzfc8Vaus3Drh1UAljc8yFo
XTTqkzxs3RfSPxzIellor/HKOkFsb25PItrBs7ijX3DsfzjX2qaSSVDNQUdIHDMINCFXKyuIbtkG
CWpUl4wkx343lKAm5p6cd45x5RhlfIGGkzfwgoubMKgeSr1DrVSk3b4u9Cxk9e0BQACUF/aYzgrG
knvd6V+r+ogXfUFJJY/NM+iuwpmEa+rW1/iQKkF0zV223vi4X6mOmWX07H2S5UKum30droVjXruY
GB8+tbbig68HQLvBDP3wmWf17VGq0rch1UxEz9M7UCSysygOYMPB3/g949E0bzRpeYQ9H1YPXDH5
ugqUR0Me8GRZwQFRFwq6qOlk2PkxpcPhnpC8f7jlY1X9ReKnbWZjQBUsJTCTKcLIcY1jH/Yua8H4
FseYXthLULw0gRVPMtBHe0/s8YrsOz+R4JHQ/ZhyZiIR8OGBTvYOV2Ts5/PXIV7jRKtiddkwMcnb
onu6ezPRE1GJbTmHV05Rud+uN5C2gElGB1PYCu8wAoF4kgXXEmOtIBbznfLWuqKRLHczb8DA7PTE
5eBDacD538CbRpmihOZvd6ni4pdy0muaiDIcfVJihKK09J3xpURlShZRu+PYupItCxrkoLWue3Gt
F3NSLJzOfbofAuLfpdTL3XoXVvpBuL6m9p6PaWBFMIF6MEZHs9NDhyNftQOXyFVt65y4wv2kOJHM
xzWv2cl42MV9nrthgAXf3l7To8ki0yCFWDZ3rjKwCT0C9H1R6mR50Wr3iK3t9gERVKuLGucxoGlv
hDy2nOBOg7H8+PbtANFqbFJtT0PWUf/KyG7XmhfBcRocXFDa73zyjfdk+bKkB5mMAGtdkuz50wye
FnEgk5lFOrc+qwch4MmDN41G1+3p72dqGDHNTz5fRt+SodzdYWg/nTsb582gEhbb6lUh3NtObegm
f3wH3wAFICLCexaxZUYV9zKRq/kDh/u0ILc+giEI5M9EVB5PLQrt+3Q6v6MCWUVXPaBhO1E4Dhe9
IukmrC8647JpU+N7u+sd73OjH1gwEtF1qYtMsI3Ecltcd4MS4sqXSJA5us9UyoGPAW6H9tNBRyQk
Wljd+nsHfSBwQa3aW27/k/9N/mZmBrzcMXu7HnOgBbMSXjyhHQnQdA2jPP0Oww61NHynqDjlEA7f
RvqGmazsDcwjGJLCdkoE37rrK04/Rgz9BNlD9Pv+QL0b0N1uNJFKF6nKECmwMxXh/03KfDpD+dGV
ES04DvtGb74hemtf4unX2d3hgfK4z8kDmcSKcCtXCibWcho91olOJUjrPtQ4u0oIOC96+TtTi1M2
nse/tPvhuQLqtY1iTmc0Eps3SJkbjAosY6oyQs5lepJDFF1l5S5rWBY17yRbJFe9wJ/xEqKSYs/z
ukGPfCMZpGYL2tsJjCb1lxN9FftV2xHi/lvZDgN57dEba37cEReGjf0/4WZouqvfgBKTFRLuNX91
0RCaVQnSUmf8af3yoAhIZ2AFn/ANz0V1WU5sErDh381nvsJYy5s8XPae9niATLEedQRES0nMMYte
NogLOcMjXd2wpht8ZYbyPYGxiZ/v549PzXAZ/RvtFeubr5A7oIhoBT4q+GQ2JD+FPdqL1vNueuy3
Db7hb9j7lh/eHsXyT+IQAlI9rx8lUxxUJJFQSHmssGBf2u9wUuwM4paU4bIfRH9cZxxKkaO+YIh9
VuGTGXjmSTSw1mBQXUXnwomWbbWbb0ro3RzM+hMA+o+qeKD6A5u96N1jgZz56xltdjR1/W166Ke3
JHy3TXZ6OehC3EgrvQntj07CnjNS5D2mKFfdrUs91XJeaj2QcmI1ZaqfME5OWqpxH60moBeRzq4Y
1c6yGJOqko1m5Dp6yv5ZEzdYZIhvGL864gidKjidRWX0AvsoOBD3ZBM6kuM9INDKp45iJNkFXgvp
UfROpdJ9rwcXrnhtqf1TXwNXlhqFQW2Js/EvXvawZT7bNrALmVTaHMNiC8uL2okS6akDjTLBYUSp
veDbUCKQgFwRSODpmLcn/G5pd4xQjAhq679XO0QF5K4SQV6YNBRyc9/A1G8fwvWjGOIdKHK6hYT6
LjdS2kG8W6pYAmzLyZUSwLBWdZZVvWfEjztwGGuA4IUsUUSzvc1ZOH1clWIaBpLRn3mkc6FnNUW3
yWxjTKf3xv/aFzU6p177/98dD3XAg45Wbwzlo76iVytmmEpDDUbvCQYrWqDHXoFQ8X1Odz+TKlVU
uAdiR4W8hmOVv+XV0Huvoda5SqicVuKzJ2HBEdmpj/AgEG+xJds1CpfDgbfErLZMdtdp63lpKdRM
ZJkcyLv70V/14ZM02vDVraJtW5GogMwibRuAasrrKf8OtA/5GbY09ZNjVxK3/I0NnndCVF2m+2BE
WT2gv8yHv7a9k8QJpZJZx0rJKPoxoGaspO+TCdmCxh1J3E8zuKd5DV+SGX2mghKBTRecPfr6lamu
PvA+vNqOCBpUjICe+hgwyUcNluRqSV9q2mPvbSFy3573eBZG77AdXq1xQdsQS8fX7U3NvQ4ilLI2
vjGm5DCOubx1zpUmuBpqOaW9LV6pjunvEGNsX+4AJ9GNfBP6+l8/HVSao7P6nk5oekEzUqIhmgQJ
M4NCFeubVZQNrlxnQHcAa6PZdBS8lfNLa63eoSFHpDot3iXDBLAhZ9z8D1V6TS9i9Mql1jGSE921
/st10i7oJo0NEdYLkvd3i0f8PKbL0pRWqrQ8Y0ZT5/j9jYIXsAMcRZ2wXSa1lRlBkVPHtIwJq6Bo
xALV4zTkwPcK/vpBb8qqqTC4VTiJy3K6fb2PCtFnAMfXkXGYoRQ6BZ/DYkgIWMbui+uQ/iOyGkX7
OcfalK1tTP4JYptu6XipAgbj0FwJeK2OO4iIGq7TcPprI/sIufXvHYZr1RisOARbCg/lMv3pE1n0
mbFkl2KqqiaLEWMrvQzxcoCHP/fAWDxHlUlq64DswsEkx3jqBQDodnd/AAQeQHT1oaBV1loZUzK5
RoDBBPbPi138u+u8cD96gS70mnv4aO4tUU5ZQK2cpmuKFxh8xBQ8uTjKLv2VGXD8ZBm0X4NPkZu7
KQUV5cQNDiBNOweJahgVy+vvw35Jc1xv1Fdl8beZq2wOu9K/ls9S8Hp5EPt5Z6CokXCZx7tIRuXy
oI6V3a7eOYki8mnpEzyU9qgPhboYtw/4sp6B3j1n9wrSMeEQE+gc2+nnFlNkM98/zRvnnT0WIDO6
ys0pJohtauA8pArQzl7GIseQ0Tv9YIbdOyJhe5e3RBiPeXzcdSZ0984iuWJJTOl59AIvQUr3Eax7
8qUZzIUu2Zco3vPtuw8VgsJiQMgUGSOW6iFzseuv4pmFzBDRbLPm741csI0s2wbp9JgtPHVexSnn
zJDlR9Y1brXN/kJ/fp3EPvSdeh7bmvrKBAI3G6exHmUl51LtqgJp5kMHt+TZBeJ8RhGh2s0S15oX
cDoXnWQrQZfSMKHefAkixvXP5C1o6//3WZOUsjJEy3aj7TMzV0wpuCqgEq5LEksnyNu7RREfFRwD
+EBFVYOZP3nrMf93Qp4UWKC2gAqZ3I6MIjgA84Q41DUAAbB9mZMUVbix/JRgZjv3J3wZdRkkn3iA
xuFI1SgUWPqLnNy5Sc/AqxAvZ/WZZ7Xyuk4jkX/UCZcSxV9AK6hebFXhNwzMm8TbTrJ2o/moGXXx
5wPV+DRm/+qJbnWCjWaDILnN8GZ5KQORHYTdsg+Kc3oW13zYGKt8a6B3eByJK1SQw+x5DJ8yoDGt
vE7zWuyHL3+TzdrjGd5gcFzcuS/+8feKvMa9+C+xf/wMcGgg/FpOXeK3zhmwJp8tdD/vmkoO9wOj
zfk4n3pH52DX5ZbJWQ0v0w7nFpcWsdFffpK+oH9o7bCH5j1lqa2NC5liV4u8/TD+OHVM1uxHIwM3
3iqZ8azYQraaRS6ihqf3jwrku7vYfkER9D4FUydp5xs7cFWkrfp6iLtJudk2ysx2tht7lOXqpRWB
HrHWB8iBew/jZY/9Xo4dpGusmuDw8mYN/WtsZzWd308gOMAYZ2Ygb5roE25eFNYLJkXh9gOFegJK
bQ9/96PI6DZVN25Tjr/Idse05zZuryezZ1zDF43oo0s6wEugDsyYuJXqg7ZY2N/Ds+zzgau+tmS6
71VVMCwbMxZo0pepMtQkLLSxRkQ9IAykjnnLuWa4ruacQJ846OA6XkDlm+4iqHiFbfeEyw1tMsIK
xw2aG+cCiOfG49JPhmSRrXLxjyKEPoqtU9osxHYnWcmcWHZAsxLoOMc2hJ+7Cv7+3E08g+O6lO55
eIVC3wsNiGtWIAnek1rRZZqjb4p85Pw0Gx8hDvGdAP62gNWj37ZJjAQ6DkQPwnm04IpcnnJawXIa
BsuJv0vNC015z01ndrqpXkNS3408KaanhFQA6utq+HVkWY8FM80xZa9Z1JEL1mADHCZCl+1I5rNq
Fm7twXjzMihpPVe9PbjTEB+KFP87EMxYHqeY7ZxB9Zp4EWYU/fUMzNx4HItBrlXCP9HJYW5sKP9x
MZ+pgBPITMRb+DDKlcEF+u3CO9Sk87cq2R82YKjbD7QAwwl3kVQNW3+kXMxn5ZMQD5wmOTmoVSEZ
+1uGmF+YJ4ip8qGt6vGRQ3Wp6JVxqqU198AGF3KhJKG+4NeEOJifIs3owrm18u96smAJGZHezn0k
Pm7oZbvyARoKNB7xxxK7W/kUeTWNpIt8ZiHil1KrifuIOroGHhQJANC7hdvcRx/d7Z2RZzvafpym
sEFm21Y5mueSeOjdppV40j0NceCUzkKp1gwemZCSS9UYjEWg2TKTc6WylerGX9Hi/iGLdVEksnDS
BBIAXuTIZ1aqNDOEzDhK7zAPoZZyTcUDGwC6UeFJsjLqt07b9ocwdhmytabN21FUv5h9x9oIpCSa
FQ7kaqTbxg3pD+BregiWzl7Bl3J5YuDd0QMEttMw8IHwr8UoIWyimitlnfJmrHlVTWBpWIy75bJF
FGdOgH9n9250gRiOrZqeFpMpFbajD+fj/ghvYo38fJjnpoo35c1ZaHxDEbdKr8/LlYVnVfWDlR+v
WlMNcjj1VAIiZ+Rn/wsenqqS/fpzDdh7OzHDTLIj57cn6sRIYUihHtGvume9rEKSWqwRnVmtmOlm
YCgew0dot7CtjEpcdcQI1oFJFqnj3IT9/iYclT5gaS9zyx669Pn3qhxmdtTS7tPlVQgBMl+u1xz1
2vUcBA/XiXd9hy0WMOkOPWgH9uSz+HtBkMOSQ9y8fWGmh+qaBVBBQiWQftiNKGIgPX35ikSSIs4O
x/NwLcfSaqksfvzYSNmaRzqQxDgIwTSjTUK+7DeOzp6WNvkUk34EB0lNmcUqK+ZTLKRw/PPBSza+
opUC6r40Ai4st/bW7+yzVRBiDCaO1cBB8TSva4vdUtdX6tySFCQnFy6jdxUPQuA9oW5JNi4MT6+L
/IDogWBjWh7OjDEuudC0aiMNFm7nYNZ1f1mL1Mw+7T87Lgfs2EBxREa/9UvsxElTdEEeIF6dc7V8
s8A7vCRHzXKJdmETqIwPGPviJAAq5lQblNgop7BEmmY/WWGYJXD8MoG9rwEtTLgOdp5lAC9FtJHv
0eOVunJxte4dtn3U8VVGiJ2Oqq+vQc6KE/86Qi6TOxhe50kzUwRT4kPKuyo+1BG4ZtQfWUO2KZXo
UJQtlwdFPjQnm7iVJHgAybB+YYEG5qhZqunySANa9opVY1qP9fzNwQncDbOFR+GcqAZpGCOhj68H
sIuZdCSHoRb9NzEzuqFsgDBtB6C9TOtGfLQNOsrNIX+sVXjHwQI3IEb5wMR6NAFvNCSgAY+OrQC/
12Zl7a10aPSE1mcUA+/0oEVB0UWDbeeubeV4YdymTntqTt5kdwOVdkyId4+u5z9HpCSMe2JfcchY
Aob+WHubO+hzVPeNsBvTJCDCEdbcKxPQGPoUNYGWZ6iGMPIajnLAkm6xKsZ5fVHZ9M2XphtNrNLD
9Lk9SXM6z3GhuEfCxi9z0tt05pZrt+3QFerOY5mb9Cttu9cIhUawMfeZL3FqtkdbBCMwQn/4CuQO
NBPtQP6rDVB3Tb9hux9zg1l+UwS9APJYg285JTxdMIrwHoeDl9H79AuItyHS7hGLb7UndeTFLwHN
DijF+MpdpQNh/VOoh0mAo1qjsOK2zipdNNbClAmPueYbkLtCCIuw2SrqY5UPmK7mmtJjlRMerldO
/WBI52azppnnpILooWTdW/zgyW7EFm1bD1bDXXpm0qzx1T1M1rDGktI9QGvDrsB6q/WbWOmB7hgU
4I13WasSmjSVpesHi9vi0lR/bwtg1IG4i51k7mPHw5jv6GdcDlosdu2htdVsu7lGHC12g3byZPnm
ddt/AzH/GtSFGZ2OkqZck1HD3oSpSSKOkUY9+cI9eSZhlJIpmQOSGUN9hcgTMODI9VsMHF+Gi5xB
Mh2LDCbvxW9XueVpd89H7fq8utmKsF9zNkqtsqidzwB7HLPvbkX510nv/l99Y/FP1BrhshyvjmMl
+RhTioHYciJppgtZsuX9MaWCFI4xYsoZOkPRyIaCxH4C4SgAT8hl0qG6KjwI9lz9/yJ82dlJIVQg
dzrRTJtXqGW0CLrZ+5nqUrygjcCOPklbbkyMvK1Kw3GeKGCHedKDe607KcSeG0FH17zORfrlWvRr
S8LVmZ+WEBFLVruoeugFrer/G3trSN2rjR320Ach5X3z2Ln/kzcAqsrdK5rGyGMoyisTHzSerGDH
asWruzdSCcMQuurq5fEBztAENj5JzLL0Cr7aL8Wsq0o8Mq94oC6AQ9EbEVGUH3B7II8hJJ6pj0bB
OYjzEBUBYc5vL1o0o2IoeMTKJxCTZkC3oy7dsrCSets9L9MWzlduKOWYXy+n9yb+Ws4Uxhp0h5gE
9SdqV6sTqLO/GfFwjp0mgCdVYl11OrsOBLkpUJFi5aIxJM/urFumumvE8A3Byvbz8g5RanvEHt4Q
KJ/9SolqlXT993yGi+7en89d71puPCwB4HXFxWhMcUna+E0zgJQQROFcMNGMBq0AvGGpoX580qUt
WQUZVETekEz+/sAB9WMKBwiVg/TsBscdjkUVYhgH1hs5rOcMdL4+tN+szxDtpVo8KHwoTEw82BVl
JeOhP+1itxf1fYMj1sYYxxnuyklrf5FYEaJzLu0lWpqXn8CLgLPX+Rn6cxUvLlOXQyxwooXeqLHx
sGI4LhTFqUb37RpLT9K4WEAKswWjCKk74AZcBr6ZO+w9c1TzmiXL4VTnfhA6DmP6WOxpQw8wYL3y
CA9b+Jj4So0GtXKzVSquv4GFDp6rqyMJB7J96tZUfhw8fgYaP93IxAHiuLSfp1l+17j/AE+XROtF
DRxy7kiuTQY4qo77jIkDIqxZaxI05wX2FPuvzat5FKbCYFQFTDiLQidjCKKuOU4/BorgDy37p4Og
pQ4OCAcaiwntBML3AVQxtTqmKO13MIC+I691WVrgGR9MAZvVDmCgkFxzlU0OvOv8gNO+kTGqGRLE
YOxr6Y0YaLb4xIIdRkF1LGBD4a81fCj8U63t1QwLfWmcUWRRbK7Im9Uh0K6s6snyebTwvURMN71m
38Osam90ZKxRIFtfaBJzCIj/ld0PfPf9FcSDvLyTe//a8XSUmV+WIlKnVGx8kE4dYjw40ZpRbPch
339kC0z7hWRAV3AoPJG2sLLfRVb1TfHv9KZDYrgn6HYglk0dFmWwrXepUipx0uOnYbxqOvuF6B0V
CLrsAmStsNKvSyvStRTCk1aUkrrWe5HpyGycm18ivmy13Vn/eRSqi4Vxi697cKSmT94vmjwlOM79
iUhzYwyVoJB48BxDv87lfNwwtSxJcj9iz6pakcNDLJkPbL54Lvwk3tYYLZ2BYhcW2C+vYE3yIp2/
qCRyjM4Q1R7dz5Y0gKZwhzRXxyss2QS/dbf9XkQ+1jpOSVGxOqRVHFDeJecsb0SNQ0INQpz6+fnI
rFF5EcEd8tcaaodCfAmQQk0JiG2TpR+St9MYjDp1rH95+b3QrxKjE5UN/jISIuCOEftja2b3Iw4w
G0owxwdIxXY0lkghLgOdP+cNDe+7FLPEzYkVpjqL/YHEm8/7ZI1WsZjjg4SQMuMJ5583mcpprqcF
/rG9U9DfDZ1hFAjJXbAQQTzNcvOUTjCUu0RBYMgCibwjd6Jeib8jiQK8SVe3OiKEhOxsh4AZih0V
PkEttU9EaDrMnOf4MNjKhtKApM3Qp2WWxEJ8Sl2mc37+cZJW8/DmH8DmXiGwROVGmCB1BHK90NQv
ORvTvGIbtd3zUJ/JDDruFpY8Vw3N6qQhs0TrQAogF51bxIOTaCgdFLis7xol0lpFng9Itr20maOY
hiFESejS2CbGIa7byT+OSYNMJ2ZAoZk+pY5VO1EdG8ln4OKxQIzpNC7hD+FkPsAKe9zdXAQmWgaV
NmaFrwfbgts1nTFlrxYrVe+37bR6361L1W2I/pMmegpq8QLHCLxSWicA2xV54zTT9igkPoDwtdLu
K7p1G6UZ7vVZjYnmH5K/uutqwVSfekHot46dDlg39AIq1g7WBCIdpqJ7CxUEOSN+gzRz5QMdqU5n
KM35EEckl1/tHE9NJx+Dj5UHk9d6BNdoIYO/OU9w9vQTEbjRSOGZhfMs3aTpUT75o5t5yJVYvoFH
RitolYcrtXop9Ev7mcW15UFhAGhiZxRgcq4LfzfNjHkGsMowsqhVqw1Hs44otCF9JuxedHuVvKTd
uOd8AtJHDJZyNx6bzPTPokoV7r3tIJeSE0i7NAUYS9GzLpbqNFVL8Afv9zhnuEDMKg+36m8KzhOf
Wo9iU61GASDc1h1iQSVEB+4kRFSE4rQWwM8Ga1m229zmR1MyU4FXF6RoZv9x13q4d/5GkyxUwWge
fRihS+yQbcYBPGEddf5Le3e4KqhKfNLKSsxrS6oLoHFy3aWCGhYG7h6p9kNjCKu6dD4iYToJi5Qr
SSf5azp767E/CS7YjJQHnakci75mzwfR1//g2Tvl131AWdo3P14bd+Tt9T8WVr81XPkpZXq3brZT
lxeBI1ZUrfJ8p5WUDcMYJDaRCEM1pv78xvYSTPZ0dx0Ufmj1uSw1gX4FqB7smEnn9gF1V/8Fbi0H
iwHo30Xp1/n/iJhxtE2obacStF2+gBs92KJ+T0U6RshMhtNz1M+n8jPhaoKDW3guUFXi7+px4JdX
omCw8K4FzPUL+nTYD7X4fDlhspkib6sga24IVJQsYzNNKRprYSzZC/dmguFZz5WpE9ysZ8aSbME3
JN86AkuMGWR/G8ls3UGUk9YbLBvkVxxZPUYKzjsIquQs6RHY/mGCfrD74omT81zTNW/7PDpNJ3Ao
L1IqU+KApsJmyw2GhHCRby7BwtewRwOj9UnAnmU+vVS3Jb+yc+PAEp1G1HHSv9jSWSt9TdYcrZyN
RTbMOUP4Bn2tX3Zsyzg/41g452Q3FbmM3E5Z7VptS9xOknS1X7vC6fV0pp03W9PKAl92yF5Cweu7
8TBsn1gmaVc9UxZURdpKc2g+LVvge9/Z8RDgTPdWDbjCjziSlqA+8QjR7uynbUP9nYZNSlRg8H1h
rVp4xP/XKYt+8QGSK6aUiwWWRw8DRqHDpeu8oEYb5wFY/z+GGxAQOBf3pfkIk+/1TzEnvI3bGwbo
R1YG1YXCJs6VCn9M9kGl0sIWoIn/DbX6pDNRuwIBXRcXtWqfSbZVax1mIium2uejqGP6vmDm8AZn
Vhq/OPLk4aKKno4kdxqkpDleALwMTxldlBXWerEueZBAqJXvVlTq9TU5kpAzYpyxnt9h3dD0nR4w
mO2zy/aorNI2MD0kiRbif4xndxZ4qjDXAMAuFqMu/3QohPELU4ak8Vv7u2O1N5dfLGSIGtnLlVg8
NN4gJhahv9xbUzInMP9S5ElAqeB/Dwo/BxxuCQ99TMackb609afsdk2jrBT8JCC7b9wREovtsjfM
k4kVhuGrqfoCWgif6iYrrc0eWFTqztXNzMcMY/H5N1lA9MLCIRv8e3vXW3kZc5BH8dCNc+ElEhnq
paRrf7g5KjOIhTA9BkiZr8GOowKNOpsw2UOM9VMbiKNWtOsJLLjP5OwtrmM/hVPdBkqnt5GVUdks
eyrxYEti17P8yZQKsZn3DD9GIwftG3AdPO7EUDqFE/4a5YqFsvOAD+0X7XhW9MtPr0P8oIN0lFZa
j8UA4bH2zxLV/Lq1GMXzoKqaf4wyJYy5fX1W/tcjiuKEJV6s+6+7Kgcm8HFJIEd7jofaBVn0ExGj
T6IorWoBLJRJHZgFE+jw6mH/x702TqJTKOB5Og3xrSzKowqtfLGvp1tmHXlZ1SF49nNS3coC8yME
NnuMX5N8RRTLVw2VH7Vg5by5hM+cGHmnIXuw95UGbtUwDxlhnGrZeTFAV9rUF74bamBHNfdTvKb8
PAkdkc4ii+9/Wm+HNrNNuYXH26pmDIHTOITktLJWHRb8zAANrYPmsHSsHjoAZS5v0Kslo371ul8o
9aj0CH5l0maXxDC04XgwOGaUa/S4911kQvOYQxmvvk/Q6hM7TZQ/OLcosIhJgx4m7sHBUyc2I+/p
Z/iRv7oo9SR32XpF9tF/nC7rp1BrCXkdDV3xTEjz8h/0ClGU+qgs5+SLtiRov4z16Q8NH7K1M2Dj
8rmITVaYItMugqcRo1TAeixAOEt0zdxvNiL7YX4Imnw4rCNmkEgaWdXpSzsmoRw2yTGuy+3Dq38/
8Fu4Sq9Kq3V8lNL/ShJUAtEaIGQTuKmZEW2OFadWLCDqZreYag3n65xO7HREFa8EiWLGdyE1QWnk
z/dTfPsoUqQxlVVRQIC43nL6iG8JLghKWFET7yKYg7WYXCO3kVBYlG/6vOBQZMLJm9lGuTStXdlN
MnBNAsvZBJh34Ze9Xllyu/vD3g/VYtUPR+wf7/tBdL9cBCjn3kYSXyzjJVKZKYcPFZP7emvARFE3
AlAyUK5sJu9VevjpmtW+36SDVguImWB4l5xwZLwAgGdnQM29Tt9qpUekfS2c7vk+2wg7Wg/lGAoH
T0LNRqQwGK5rXq3Ny2CJ4N/KD9Oq860/7KK1hOSeLzRAnOAoNA+6s/xlymDjffJkT4hjfwYERQ/8
KF56gk83xqWRkex/aQqUbwBmmjXSRpjPboap6MfWfagcLFUh8nCQcO6Dx7qFHqfBPSGD1e9VJvqt
SL4KkCoXHoS6LH3YbluLA+CspyOvtTj9mH+Wd5euqBzNyQlHPoYOA0A3xSfMPcR5w/vqUV+riNvG
KyzdUXhx5DQCJx65yiqfzE9oGjkQ6VUp1qbHLckSNtef6xkCMla6FZg8FOk/iq+XxqtdNIIGF5ns
kcdezp0fGj56KHbTFm0g8ugXHtKuyO1U1YLNISlagKQkF430wOOrYYyvCUmGRh5e2XS/kTCUrN8M
BCHYQppJ2GqGSdpuxfHG1fEvakDEOQ8PlAOLrliXRhbFK3q30cdP99i1QjHwyYorTdvT3BBoc3aV
X1LRgBPCLzw472NE3/9UQDmxm5UjS7mwBwveN3Vnw2P/Lqz+FCOf1X96Uh1wVD+iw3Uhw4PKpX4Z
NuGIkF+aWYOBSS2mEs3PYINUTiN56/kwtfwxeEyrYdvOz3PNfwjzCY9YV0aph+soNlKb4eN9GeCY
/PK7RGcktGG3/tYXd5oa9Kr0ZAWuGNSWmLRiYzoSvRkxbOO3Q85GsLmO3s2CAOj1vXtC9T80SHZF
GQeraLfqvOM4E1q1Fx1GTXQZ7JVyF4yGIFnLZG5asIq+5deF0vto2QqMy1Prsb7/ZQjtqFaHTg2E
sLagDCx6aUx9N7qFzRv9YWQa1R07Qi3ujTIa3xAdLVaBEnMpxUY5COE6eZRuLUlwhEeDEZhnRAkH
6ziHpxoQLVeOiSXlBUerhWoArwxbUTSKNE7hDnkhxdDLMpZdNqslMn6ECRpJ3BY6eI4QnSZjgZZy
D/eubSeO0/sSvdfH+k0DWlEPEbhBkjqf5rRFTvpJ9AAjAKcjy5lK45r1nZP4+JAYiTv+jesZDGCP
ZiEyRIG0Z68LFlOSA2ZM0aSl4emD8Vyd51igc7bU3X3Os7CbaWGjL9ccMZwHb2LzX7q6DtazLzad
WefdViNlUuXgbTU1bx5CFQm98cJHuPfzGjdwjgzXDPILOO1VbmYI6OSuH3IhcNUEKETxKFKVzeQV
yhCXp4Zb5pGNj/HAtcJyWNVrhSFMeldoHsJ6Liv/y21IX8bps9nIsqJ9C49Z6Xngl3RH80wodV4R
uxv9wO9yshqdxtTlg4zQ5CEtomNZyL0nLJkIaPPKVkgr+XN1l0mLnzl0NS+eZUinJueBQwIaOo2Y
4J1q0Zt4YE7CGyk7OCKszXyDl1Z6SAP2QJSekD3T8U3JGZd7+KpYkn6hd8HZp0GI3VdpHUBBLLg5
OeHxCAMw23UeesGdOm7igNfMRUCHQVBEP6roFZqeMpgbeb3CqQCBX6fxh+0A9WtnFEoesGX/fvYY
2sm7ql0bpT+rA/pWxkNRSM5I1VJVeVs0SZoOFUfrGLIzra/HEiA9gCvWsNiHybB2dYGSC7cA+0cS
N/SxHI2/XBjp4Ti73owpgPSxieliulTYsW/1tfGMk+UEnTo0aRQBHCYH5En+WGfLODV504tyvdfu
XPaUSIOoCkpZg8NjawIB+4c3COT8eJ/Hn/FCZnMEO8OXj/bAAn4s9x6ZkQ15GVjX8VPJl+81+9xy
sQA5n6Eo48AXoWXU+z25f9fFYr9bmlTGKFowbYydtCrkB/myKeqj0QdCgbgDFC+pJcfVYJbKP1ZV
kMD4HhWoOaYYCLRY9MUPu95dsCWfv80uVP4ph0huiMNSCL3rLtxHMLglMMwo9A0b9/IaGiFHupQv
ghZCCi+3irrujV4rjkCnNh4/kdzrjqfptmiWiTu0AymID+EnUejZzol9+lK1a36YJzvp+2K93x00
MJ7eyPeXKYCod+yTd4uzBBO4o+W4HdANJZQI3RmheUwE2q68nVqesDgYDjxAROGVnEvGw0jATMNb
gdw/8Va6LXPEdlgz/upaBx11P7gCnPij1bG/xhMjqOyyx9M9t8BpIt8J8GWq5oAPhbcwjDBILIUY
XcK7/xbWCPBVjPtqC708KAEgWxx2Kq44Paj92ZOM1sTph+KquuuLVLD8hS7sDkSIsN2Wr1CJAvnN
wkD2GlUIizN35nrcQKRymXykKVXkKwnusHYd3KhPWN5MNMY9OoZGrOAb2wpUS4OFD9fOIJngfPZP
khEEER/D5zpFsUpcVcr+00FAE9lTUPTEbabk/Gz6cuyUBWHhn4nBd6QZWtvnfdF5uqLLfMd+jhTy
QmPcY3e//Brnsa+2sqPlWHMrzWYPSh+aP2Q83C4BaDZbheOwo9sSBkBHKdEnJ8w1wrfHxN42Sq/H
hDRvWp3SVZ/yf2U1ZO0gYvNtV3RBvXjqLUPqiJ6BMPM7aPKyVCfkfD1c1NvJ0bvRQbSPgE7HdsnI
h+unjUuXFl86moQ1TU6PvzFFh99BQ+3XEjA36Mg571k6vQNs+ThMr9IjXoqbMI9V/zbpCPzG8/eW
4bOSj4s1unTjkivczT2DCxmrTqpqHkQOQ5bYjD+CSA/UVmvs72tLbRJf6812IYSHtLyPiIU60Qfd
PLr/DlHO3ukmp4ZiRPrDSMQbwGMfYxmqWxYsPxTrZe7ktJB65ZeBLYskDwhWvYQSCFZbnxMldvU9
GE0ZiZ0RCAzqA3zwQDfP3JPIYSOprmY9hLRmBdl9+eUcbtR3O4lDKoeSRvESAALYjHd7VCWqgLE9
wDnWVgByl4yinn/D6Wn9LhVzmEaR0/d4ihNgCVRl3LRbAcHkKCBGPj/4xw0M6x2uj6XpqsvENSRE
lqVNzyXut7P/qDiQv8+z2shtNZZn2kZ7lkQCew43LNlSQ9FxhSKMJMumPhGSPGHfeO5Bh6R2+5PO
nLLEzf27IP/08ik6TMPdKnq0zGUPe7PygD7m3O2strLT22SZ1HkdKJiL6fxB/BUiIOU7YFe76uim
XYjcrZu4O8S58mnqpQB9ekCwyCYnPefLe2ZNwuCdCvAiNseqtT1FjC+ycW11EDYJlYOEm5oSpZ6r
Rrd2NUvupL56jYNH6YaMZ0mvf6eqbs+j5JrqGsPcEsCwsyxtP1Y93wi4fPNlzGXM6+gocoDsZSqw
nVG1+oY4uHoeWl/kDoyQsEDiM4lR8ENw2evZCSstTAfJe2Nrl1U/F7CScMoS4qPFDMNKb1XntxB3
5Cc+1ltfM/1zTfr4pq4f0CyOkW5e9NxJoE6Y9eJKIGf+0tIr+VeI6VEyStCeB1UnPCnsW3Wdaw8l
hEQmJG4MpxE8C/RCRj20IIjHTc92fHIjb+yBLoijsUIA6G2XoVfLequ5jjuo7Hz6Peh/E4SzEgBh
6nO+qoMGEiaQDZYxWMQNJrNYqCiIPTTZAWqzx14CblpORgZ+68acA5De31ktfPzA9sbEbjDPxJTJ
dZbVSG284s+5MJnVWeLQZdsM++RqZDQdVXSmojfhrx7FEEFjW5qyjaqMiTsvQDABKpfH3/+PMpDG
jn09eEtv3wbHlVx/puM+1Fo95M1//8ZN36n1IV1b05Iocgp9yuLBWYKLHRHUDI4i8XSJOd7eUb2W
RzJI/TnbShU5X1TLRNFF4517N35APZH/lQUvH0/Wv/7gWpm1rQSHYXYd59aMiLHXyIUMengtmxOQ
rQwOxdzEk5LPrPQvsrb/21tUI1M+JPNCcPTDmXKS6JVh/tZXZ5+k+9yn81IxPNG3Hx2fdljoPRmP
PQLdTijikjXbfDCzBI3oHlRnnn0WaYubAcT6xp5dohY9wXPkC+0dMxvtesASLeepGNcvVpr91+fR
IBnkdZvC/WiRqgPrd8E65+BKTaA52vm2ZrVv4LAOnU1ApA+i/Qd5fGAPWSgnzY2A2X6bHgEo1jUf
fXxao0ZoXR6SwuMRpsz0kD5uchYs375q2rENZMqOqzJ22oURFvPeHS0dBkPA6ZTalVmakpJVNlOL
3LVc+1E5IAvVx9oemVWfb+LBlBkfb6DjblsocALTvn/sP401zik73r5/iFiRDnyOcRIFaa2Yc0Ml
68KRNm/MM4aMwkVg7AUkFVLV8gaWDoERr/p+ZieNO1DBRPeF6zu2oa/df8ROMP7lSSRa2KILcOP+
sTsFu0nnfpt1/tn30m/xxQO36WAjmccxd8GETUsxJMGeamkp/7k2jS5BxJr/bubYpL0YrbSVO1Il
6psjmJsPg8iBxMmZWA+G+2jeNfPBZzEIuiqRgsfa9MPnXHFWjPL9LPfmLSJvq3TmWDgyEDO/i6zp
2s67wHMvhcWnRksYHvq/dZ+eKhgxZNE1Z6DvFDy4Nk6K45bvMNEv/FzEgfRTKmV2OVstpgtneGyX
C2eMN8zb/JAvcN6nLdLYEQ5YhrfcNYT+YeNMMohSR5f7+MFyTv/Iy4htbT6a+5eKTh1+VGkR+VVu
gh9cblSogCPC7nKirqguxTJB/vZvMpOV84sg2Dbk4gdO/j9cD7QavhETBbTMbhO7F43FCgGVVNDI
j3lltEMRn5Ol//+Ni4gcaoKYmBFSHUbW+Tc+hE9CrWAb8o5AudFO9rtvgMmJf3WnhTFX2h2yMOZA
6pJT/iCCVHO5oBLh7SkHgDxlaTQ7Dz4SHEJAX4qorWCMLSWVabpUQGs56SGbLUSYZmgra1B6YThV
t6YkSLTCnVLFjUI5QAF1MS5dx6P8x1c+UZ5qi+FkO+t3ALYWZY7fi3yhQAEq8L76FJ1ZSrX4aCXL
4oy2MkCLlBjBvZ1R+wEcyXlp8fUAIUE9b9s2gJ0HoIwegPUY0b+sl5mEeQtR6Lk4Gkuj5J1dfF2N
Wqhwde6rmjg1MUrgnjDIDhU2nvLDx0K+cwKlBMYr4u2aRwHgu3j+fLeXtlQ55PEDZW5lSvpwmtXu
y5qZvF8tDXOxMOeGisq84YADNAM6OL+1O0YuhaeFN4cL2xdeVLcHYsQ4+EAu6T1uMgL3iPLhmHhf
W7teMyew6UJzLkVA+zjkWrSlIj5vNW6yR6CgoDaAohugCkXaJj1FEdzwfKqMIlE6u73mVnBuQuom
ILi6LWfT7PGHvP4Xi1VTGYs/qPP4x1EldrCH3n6F7Rr/o8W353I6hNlnPnxxiup5wP/jgaCjvLMm
zWJH44ln2DTlhqdgLxxEGe6QdtcHPlynY7RFzQ2aCxTSribYhp41P8J84e1vjWiGM9itOyKi3PAw
OTesbIXM9o2DjxwCbei3YTvBHACIZNWMQMejaGlVgPZ5CMRlhaxeZgvhzPSZKpmED5XtWtQAAQZV
xcPPd6Cyb4+S/eq9G9Q5HGDjMEpX/W/Qph8H8oGxeDhY/K05A27xUNF38MVKtOPGMeM0zb3jRuV9
oh4Ds4L320dx+/+fn1HPiJgoOqcdeXKwzNl15EAchJN/PLRs/fkTwT4g4rOlRZahZM9TaaKFof4S
cad0A+lVkrCx8UGkgPzcZuYoEjMwMpYcQzwCrelyUvvoC3HVzJ6ExGim3pgLtmwfnR5GoDajSzHC
5okfiugp2sJQtS+l3X+5Cvk9iPXn+qGyQL+PW6v6Ji4j/fHKk9THw2pW2MOQIdD/rTNiE3nI/0p0
bTa7tN1ILFqltSssYtx47ETGEklqx+xp8tbmClbK35nfR5ubmTzzozlYSUEoapvNgIK9UGV5YpqZ
7X35px/41o1ZAqf2N69e+cdvHEDJO6xiHbe1csrm11wFyfz6qYAYQa4PlPmUCMvorTUvr6s3WAh/
1jYaoJjYds0eoEjgs0aYSmeyaq9A+rXbo9QK/3Saka4LQF8kczo0A8fefHzshQRpuPK44nCX7MG0
h+4+Z8/r2yf0ZBZh3LFt4UA3/A9gCKPF/hICT35SMH0wNC0Js5aKqyFp1s9X5Jbh3ZddvrQe1G8+
DkvHr9fH3KLRsnGsWaqXZpQyZdbkkF0cnHf+xw3TBnghcQs4gVcMQ+InkG033SRVqa7mK0dt5D4v
QUccjSt7HHZjfRT/7e/P6plbhELw4fZbet5mDWXq3DXND0jTOov4K0vpnGVRpznsr4PXTNE8FFw7
BLkZY72p902cYFZKTaERZu9oF4faegz8MYSCFNqrBohv7XE5r/jw+/mtdfmzWLIfEnrss3p0nEEY
kVMNe++AtS5CzGt7TkAMu/UsXf1MhWpJjhEsEkt51mNiH+pcbuCfP8LimqqSxnKjw/6ldgI+BfQ8
Y8GhgPfcT/F+F0R3/kjWnlEgbWgAIQqxIf/5/Sv1VZWW9ZCQwly8aPhPlEZfdAW0rTkvxGw1mnOC
K0OV6cedclSND5twVKhc8B+8HuChFcfEVQm3GX927MkffRGglIslvguQ3h5IZUzwf41Y9CCITdMf
eleh3U3SbK2WYpn9GJsTUBIWQLEKFNxkshSsmwhQp+cuQh4965U4EsHLgibPG4vPf+SbIO+03/gK
iFbJzN0nl8Hj7087ku8lP6ZLjp1gpTKd+wKlGSiwWi4Rdhf0Eg/pKxJYMQwtuvUvLUzlH6uBAHCN
+gPwaoVdg6q+WZG84Xy4jAKuu/yw4JIXxnVA3/x+3ZLIfCfdgLYJy+yoAaWU/JUDrfJTDq6/u7oG
eb4trCEquK14nQonqr9ENndJezt45CTyoEyBakbjv+Mv4ayfd47hrTpsm3tZJZOl+f2rcD1IQu+H
Hl2o79yW34LJ3ygzTlyDt7DvaaWHb3Lkj6JiBtui3pnFBHY65bTanVZ5QpYGF6jhp3qq9mkef4iy
T7og/CfZE/3Quc0IapdrTp1FXg6v8bO1549JgO0gx2qmq463F5zzIrG1tmFE+iGcZG2miod03Ud9
MLEwYjVZlfjiWQZyJ71blthHn9WWc4IK9mH8tf1qGYn8uO3o1CgGdqN5iQQXpE73J2RNLlzBJHJo
RW96RzoHe+sl7g12fI/9vuVPr43+BI6tkvWJTJ7WTQVOZKhFopHiB+XRgER5YxiqHAoJAEkfQAn/
JCBbH++WzGpo+B5SHa4xM9IfdL3pqb6TS45tLTyrcdf5njDlZtvPWv6Xr3iC8fdwtgfq8tn2c56z
pY4OntZ2PkAzy4a5uO+/9RNOoPoQDNCZEn9cTwP6xCGbO3W1scMVk0CZ3mNpd0Dzib6KAVdW4Ohr
U+M5IHgUrhQIv5EJsXY0YZf4keSwpgAD7BFpeKvzI7LrJjKwwKudBp00mW2go1GEAKSOIwN02D31
tT9rM5aPdNk65333ZnBS1M3wE8CBgKeaAnTGD0XVSgfFrBs+hSBtCTD6d8Maa6EwC/VJdjlmkMFS
rK7eXCozR+lOMU1zM91avdmaTROluUUPjpAUezBDMpYU6h/VsvrTmkmPOYQiTg1ReudWBxDZ4Lir
5ZP7Y3Ud/YhfoTPJA0LhS0Wc6KLxSy1K7+j4fuPVaLav4VcEf3Dunkp3nwLiqBbQXe6kjolw5tHT
TxpD9RzByTIf5YXCgzJv0rBCrUNgeFTilYanchlbBgWcXib0Mk6MwigVaJyllvvwzf4ZxSrW1ROx
Dv7bOyn+yH7x6XRg6VCqj8rWSQBi5VnBmJ0RxpxM/vGJPWg4aQGzyfAA2mu7QiqmmD78VX/+qOLB
6XdIyxJ9uk1hyyuuaq3zCA9ed0UP+lelQ0Ng1H2KK4358NT0ac9XV2BMn1yAOzPy+PmM6DnPX14d
Cu18FeLr45RoR+hIn+Tcw7zSUuYZrtDeU5AydF7IYVo7pthisjg5XpONNux7RXAFZ5hrJhLem4kL
xhNrHy4ahw6ZZHS9imqQMM7aPrHQ03AQMThyj6Q+65IZhHy7EW17ibt/Xe4RiVmYTuE7Zv5k5rEa
VQKhN7iDMUEokE9cFyJZaTPMwD6jOvbBu5hi37eWv2/vo4EVTrsI3sttuZlI/ZxbRa2dJQsLoasi
+jv7fR0RY5nvC4EwBONbTvb2rGTf/U8riUUoaYNRYP50M1CRiNhDiEsKsRyt0rpRaByUQSSaaqra
ERn4YrcSB3TeBZAWXmSvF+eSxKdcy1Sqi5f2fQYG22rJk4CaeTV6mOaWktOGy0+uQMvG2QuuS2Ea
g6q31KLx85OTQpHZ1ShRlyHdc57yxWoFx6OguY2s/V3tT7l1tC18lqSNyuszyiH8HXcpxMdwiP3Q
QxZFako1EWaWYNHTvmu/x6mxd2lxeC/pm+r/QlKw5dJijOM9JmC0RAp0h2Z29mdkpJk7XsswaQPF
nbm66YJJpB0i4SbZdVbbT/na2eTve0ixH/s34HeYC5j9nt2ZVOFZIc2WsNa0ea+CUN4yoQ9ECxJ1
xNJLYXNe+gsdKDTsqDYcU9dqQSb+G3PjgzUwV/I/XYa4syMh/Ety8Dc+KvbRA1sVdxn2XxsjjAWn
Sdeo5Fao6LQGlpwvqZcr+lBn9Tb1zngNawCRgTb6wwM8Ir6x2U31GqDU2uoe8K/+ileLorSLJSco
V1q9qfatf6CikQ2rjAt9AfAydzSvm/m/XiK+Tg9M5Y3R/m4CR/vFgOq4w95Z1ae7lIukwtzLWQho
E9Y5ESb9yjwsFI8z+fNA5d690Gm+oBHWw/XojlF2EyX2Ht6NDKtcf+5trDS7K8WDkk5EvWmPjnR7
JrBIWV4JinPb1K9h7ie7NKCjGTUl34C2/bzE+5G+a/tzlAf0Q1Z2ftlxqU6gUq2GNoHufNkcbbZH
uhzQn/15shAKU5JO5cKufoSH8uJEeQLGmpzHcwIFQ8kzJpxg9ya06jSf5Gl9L5GXCHEWSJs0Sdqf
3A0STucgKD67W0JFIiOO1zffne1WSclx9NvPCfbZtiCvd0Wt0EVyBwpBqEd2ORf+CaQXQkOOGEAB
qGUQu5JdYly5nzEGhIuNNcmhI1BC1qILND0JLPX3fZp+VKwOpMPQnGeT4/Lh9J4nF5eI8f6M9ymj
c3DTYdZSBSd0uukSB8ujjsGrI/yeJTm/2LWU9/2WSq3OkfY1/NTs2XxCtF9lN/5J6KJVhVEJ/54p
C6/ZXtpbntO6u7qVOnNs8WP/thwnbxSK5j2eTRNujK464ChyuZuaofyFwB5xKyArmY3P8Xv4F8os
8DALpHGSW1fiID9EW5Ev8t6B/xvtldKQLI9uZiiq5zqG2NJUo43axxvDfmTDQ8ZmWF67OjKForJs
mqnAY4fkYRn9eqfgwkYSRvdQpJqJ0Bw+dA37Y/fKYp/Dvi9i30SlzZkLG3cyh5Q2UfI8gSoSXIFO
MBdUdYBY0es9Z61QxwF17gGKBmgNfg5c3P4Wphsy0PgJOwsBV3lLdnt7rt9TnzZqITxsqHrGCr79
3EUjBpcBcwEOjdPKPR5w26Q9ebCoxXr0NfiTPkoeUjA/y1sSrxSjhsV/+TBk9sBokv53ZEaMFi2X
XcV72EKOf4ep3JyzhHa+1l5/uscAK2BujrqvpZUZioyzuckqBfUY5Y9EwGD6MM3+XBKYrEZWi5sX
B98XePCaTYsSTtOdy/7qGbHjDNvcniu8dgYPZJE9xQZuzGUzZuwTGTWpdEss4K6uN+Mobu9uL+FK
Yc8ca3mBKxljTKyofrRBtm0107pnvPVH0Yn7xMbc5T93gYkbd1IE+vmS7YthEbUyNs8K+hQuiO/M
Y44jwuUXMUM1J85f4nVFppPG1Hg0rkIOoUYX1SL4/oy6fDchc5vHNDcWgR4VmYEefMQJip9K5stc
JW60ZjEzVX2gNwkpqJtgyEVtrspw8ura3HOQcUFAJGvsKvVIMW3tDu+oX5MDzyNyIubySHIy0tv6
is8PJNanMrhtJkSbWxSpdhs0sieToG8MI5vhzF9H/V4FLYVjPYRxnnAvjC3KiTzKPw0Sbm+7JT/S
MZXaknd2GtJg8HWqBVxKfywAZWJoWjLoVNShtg2vniC1UFIRlyZ85Wholyvl++oSuMYCm/YI9T1n
bK8HHEHwcKMz2diezuyiSURK58XTbUYI3BCczC+Aff4hQMR8hIqFLQHgHCR8t9YaO3S6Z6ASMMpC
gInOXLzCKDpo+k8Owe7g1O4Uhq51Ik3FgRFky8eC9RDgcAWhhCxYGeqBDHlQVj8FqrQuvdLvb99R
QoLKVDsuJGH8I0IflvlmEL93dYgZ5OIITPX5EZ3F4O+9HbxDeFyeYdv94cmKPTVoo1vACcUNI13R
3RfVf44q3v8CCeUxQbb4LRbyqLxzNUpxbrr6FuZixnF7tdD7GefVUBuL01outNS4nXKv8oCinFrs
KU2CoNI74yjpy+A2+RjV1eM0f70MA7j1wMOINDTUuuxF4d1B53CVsBzCN4+ExJtlidsnRb4sUYSn
6okkAuunPdi/1D4PQCjvazET0gW8htfro2hC3Xk0Vs7eUfNExNBsKq39b9WnoWGtM5i4Ewq5N8hZ
uqukUym2Z53YoxRBXnumdmYdtU+OxoTU1FcX5eXazN2d3VEntV6vXv0MS3AjIZ++8Zoo6ZuszPSx
tu6Pvb5qK0XmopUdW/+6O+/0wDKufTcNKrjh/gmSOndAo++bJmdpVS1Qb0UDR1xIcDKqWl4I6H3e
rDZCphbxqIZwYwy1wBifYAZlozuefFUhJEIoqONTq8l6VIi/40HB/G/Z7f5pZkAOvDe5G1H7ZSRZ
BBKAqXpuxvYtrMf3tTqITEnody6YkLvDvpJatqIZCUgiOIRMK/o2HYgYSQj7gDjatOQdhjZ8jiAR
9RtpzMm/ulgHj/BHI++ehyrxg+day5ep6KqhkudaZGEpS2n4oVE/PPmunPR7XmIJc8xal+cgS+rT
nDUmKR0mLLK5a1EO2SnSZMNVYAnvbpASOjs1JEGLNI96E+i84iybpMp7Ti3/0E3IkkZQlXxywPYu
DO+zXiNVOlkfpXiixePmewHTnjyWmiSz7hXRGWE2miMALJC6EiHaqMD2YFHc6/RCRt8nYi7sEpiV
7mseRqM+lDpcdF4xZ2ISSyIXC7FIb80B7ARxKnh5bDqssQZtzboqCOA1MTijCvMgdCAQQFvoauZ7
LJ14SurZdmIGroUUkgCvNps4PFx04/3l2WY/PV+Xpw3lc2yt+9CId8HGF5htmH54ntp4si/FHD1o
q3pb/KeyaQ67K++QKFLqu+5jh33EIsuph7b/Xe2WZtxuvEJuJfPcZGCKBJ5Y1/BvoHdAjPWBaem8
pTI5zzYkJU5gijmAJoXe1ba/9yaQ5GJ5HGs7dvUoKqibE7C4GI1cMe7ucxCzPlpAi+YiAgSaGQbY
l/SOWuN7RsRHT5L8WaYhSpQxJLZeseH8m3KfEG7qKAt5JMfKCNnU8wilJzB6A3MMN03A8BUEgjln
vNGg7YHfcIi4UvwvscZNDTd0hAp3kiTyoFcYYdCBK5CtnOotOcUmVjc/FEG+baDjKil7/bSUcIAL
RaRLLlGGForo4aHjjRaliPvqRQRSmtJjHSXcu449D2ozGxBEotivtX9eMnG2hmFSceLXGnnE5lFH
LCWJx0/JFpwP2aLZpZRE4BlICriv7QaigDEE7yeduldabbwZ3BESwNJ00Ac7SF9emtN06JTegWOX
sQ2D76XkiIaBPm2bcTQqaODnDCeHDFa1oSZRJbmGWGLEhdqiK3sZXNDui8PZcK+NTHE/bt2B/D85
Th+wR5IrKTk2VuG7WbASLYMlSf+Rh3Y0JaVAC5LeywRYRm+ZiAw1ShL2tWDuqUMb2RjwFchRq4ro
8wvK3rUOl27TV8kuu5mR+xi3QYw7yoKje36RrWY75o4Z1cz6dh26xB3BSpu45azcQNzmIZlo/cGx
dtrmuxFrubiHC5fHH9xNMkDzsePQEldAHy5iCrLLo84KTWyAk+/9UForCT5cw/hl9b5S2zyf2ZgQ
522DPoMHfQ5TavMPPDQbm+u7QM2iEUmbZ/Sj6gjkQpqZ8WobvPJR9gOmy91c4VYFtE+BWOWefyZk
cVJaONoMqDgsO78JtOmXjAbd17mposI1hoUCkohOSol/FRuG9Tt3p28rveJxk6xhYujW7rj6XDdt
Ak6scwgZSdNhRJ8I4r7/baxPtOlEU5XhwJtnY3PNhFGmOtLyJCOZ/jrMK2wQoXwQXr1dRk0oRqj+
Q2960J5KIikXp17e1wOh/1MCKtwNexqo6V2pm4/UQdsqkEhHu8mBMEvFtbzERIBBd9M8eNcai5NR
R7m6eMzfF9qZzLAPt8eEoNqkBbfM/Pe4Tx6pV4pXLy5S30z1HnRvI0FZExm58FZJJkvbhmFCyccc
ApvMEDeL5UYAFu6qzUv96V6Xbqb6b40T3ObkTnBJmECGebhQJbSNsReYfj6woouiby4AY0Nk7NnW
h0gJEy5wXbcde4ZqdC5ZsztWhu/C29vwiaYEKr3/7wbiV0/SKzcD3ujFWWX4h/Ej9bJu87XpxUD3
Crj7YGC32CTJT91QcU7jUh2Fb8KZziEbwcK8b/qTJIiGQNe3rSSFZ/C0sXU6YtdDWsKfArUJ0+Bx
ILD7O8GFZDdnJwBTCwzdnhfoMNFt2TVhFaJboFDVGkXQM9wD0mw+XcliCjebb+OoP2l6suCR1e5+
Es7JMImBG6+MN76Rfetm1G0qUN3BblAOo8GqNynCkdP7FaKv1ZFq02SJJJjfAgGAosg4nVE21trt
s0asFUbJX2S6ukFCc7L63NtPMPvNQpGPQiBGYw7MpXLqbjm3LXG+TVN98ey8VMiO3/5LjhXdrWoT
ersFdJNygyzS83zjE4FXZ57fOSJUf+PkYWCNmqxrxShmkZQo6eC6PjvMP4WTuUY5ctocyaDzabDH
TEWfNAZTrMSWRFdwbX1GDIOeIZAN8lBuuI6Me6VyZOc7QYEl5yLO21Yr2M59+TFtTuTRKtzIxOzL
/T7jj0GGTz+R+8AIRe4HSLSvxSL55y0EbMnrSf2Im9L+7ULgkA1Tt6wYDOh9rmM7tEqe5782UM2A
Wi9o3vttl0oBOVDKFD1bZJk0dcJ1TZnELVQD4rlY3asc515jwK6oDuzNH3r6ELN3cx0yuMc5sqsz
05lixRYioDcXnCb45D2ZDXyL/fnx4zX+I7GIi5LbArNQ/kXuYWiHvR/TCtpC1dPN8bgChsaShKmw
fWw9c3523nGxGD+lWV+r7+/9+NyPs693M2no/mc+c5ia/QgBwZb+Hw7KQgXCIzYItNAzDdE6Czun
lff6iJqu0eHUyrRKynv0lN5R+/OcXPRakgC5SMGNBvCjZ3oDY8NMCpMDoq886FZVTtmbEUVsM+bd
NZgXid93nIDYLK/tzFO/OAq1Ijr23yLHvZ9zsoQ6f3MFwkj1OKHDzQx1TOMfJFto0Tp3zRzJOIGF
NdmLWk0iXppXMnpILTZ8qhhDGXK7tGXchrmLLLAin1mg5ND2s6DkDUs4M5Zrt3H8w6M+FFahsDcZ
YoIFOKunRf4cTh3oAOKS6aECh+PT36vb0Pk71G5eATURNL4ko/DmuQyXvG4Fkwe6/nSzpvvFRKmg
yGsFw1eHZl7P88jwQEMKT3FNCR2Inyvmy80B8diV0xhpcUKkbMbgXRnzEz6WeyYOZSVksmY4csSf
ETyfN696IKHn5+5pKlCUMy3gz1Y+MhuzpapOjsnm2AOYQjHJx8GX6YIjjcLxoPUin09GKzYTbyoS
k+Osv6JV5fbIeumzQmb8M3QECQIgHOHC17PdM8n4R8hJsDwcLoN3gbrd6UEwn1oBRR87KmazYWB7
BGgM6E5vg+Okg+grjV12mXoZEQ++S+e2RCdXbZD3BPAa7kjJwzgN8C/RH7bfU1otowqYR6zSARe6
Q14qMdeQAGfcUYC0etKJ0IDr8zqSF0qAtIGsGg0rZO99CN6ZoBQxRFmxYoxD2/lLuw+/tG7TlGMC
y0Vldgry9s4UGKOw7m6AkLQB0PH+820nuwa4bkVqDUv3sOKmrgPqBf4FitctjYzOhQEoyTiZP4AG
c2Kdh3kUXabuww/u7Fwl0ul0/V6y8eSfNoyH1gsCJqI7vGrRTJd0h5LxlBwMUXfWDTdXBrOj9+zn
dies9NldFlrvVMlKlj6yy2us64PdJkCJx3eme50quofbktjVEB3o70lbZS6wY69FndmbeuvlmrA0
Qz6EWPQ5/fmU3v2sAN8XBXWr4ULJWo+B1X30Qt7YWxkmtMMAcx+wBiIkn95ZAriskPQ4xP7ZedKF
qoeeJSrQanNx0I4DiUDsoSEZp1PkCovP+HZXvu1LtAbbinPNxxVRVkfhIMfeVNeUHw+NcomumLsv
ZaQtRrlE0ZobyQsDCk/t2UDwFi7TuMHppGKwXouBAzgag3lB2qpEC99hv5+ZDtmwmtfexZk2gQV5
bsjV1KpHbphgm3cw9Xz1OXs1SltxH9Fv3Din2UjYf7OHhv8pb86DzB0keEPXNDSWzFSIO63WEnsZ
0i1DucOIhOpvBkAfBVqw98460EK6N+Xg4yqYfdKjAPTou72i2qyg2CjMS2bBX07t/K5tJmJ75WnC
wJqg+cF4E0aBORrTMHaOGB4MVxL+t1F+VBLY/OKXJInmDtSMx4rUjHyrxBgHjZsA4+kyfBk7vbcq
yf9tVT72lL3al/mT1NGIiw33FrHtJXCfKZfNxiMPWu3nava2v32LP/E+7C2jpflnewXC1rkMKe3U
XKj4hPH2DsX3Ju1PA8w7uEKGh8GysZhTfWGeFBFhnDTqfBIRDlvuseky3iJva88m18gTCkaajBgd
t0Na2hzZ15e/9+0Gxv2poskvpa8bleDkF4B0i4Qs6SyUTpMFKTrxuBgapbvMgadFG+4P2eW3GteY
g+nAyto1/eZAIcD8TEIlcEEee8K+anqf60YhEt3KTkIkTcerW8Ua1OLclyPZl3VD7tWPFuXf+g2R
v4xwNqomNXVs1CreAYkmIkJYvzE9Gyce5dMIfxnQm73CCCnr39b9MXiQ98UtV203GbM8VWaUoeCC
KhpXOysGV1OdGDug5J8LtQIRsWyGRpmn+BLq+2nOTUphNLBSjQBQNBwl/ELFBo31P8LrQPzuZF5T
Ze7ournTa4jeAo503uxcq1XuevwqZbFSRUGl/wnzoSs3ZorHq5zcnNl4HRGNL1mPQq+zzKFSv7uD
xt7pn/JAvJF2t55+tK4cpbIIQ7mq7Je/1Q8n0YEEAEE36gp+vXd+bp9ercT0/1lrhsHNmT+MpOXB
1VvLTRXf4Ey8SUhIAZQJejV/z/Sw9mj94hdFB4+0DALvnlQ8euv0D1Qo17/aTPU3KkHBlseWeJqI
0S7TNIPHZvNn7TaIOEL9n7TPRDXbe7NTeaeS3nSA0Gk2jZ5vn9JCAHNPNrYMXWmmRgXac+MYcvPS
X7KMD51iZL3lxJuMKxmqV2H/jlYXvr0cFs+Efkd/he6d9w1bMun9DQ2gqqzDeCf6cQLiiTkveiPR
MT6L54nd2EP2v4CsEKZ2rkr0Hsk5rU4KLssccX5LXh9xMwj/9EAuy2fgR5fu+wAJhRrVMHaUzKOH
2UrPGpLnnxJJIGdzYbP6ZAX1ZPZD0mgQrgrmC2crC41e+6+BM7ZPiA3StTXUiGv1TH8LVIbQowLu
lDOMBGIAZXCyix6AZvUoOnUYLX5DaYCnyx5Kk88SoCiDL6LPMXFjPgyAVWtcPvTmBK23kIqoVKlM
7h1vsA7JPPCjhF+yJx8mnDiPEfxfiYb179K+j99hYdMmCUjrxqBp9PgPrKqri+0uI9p6dFhWGdSk
8cVqW8E1b7o0LMppAoxoS+e0sfB17MczrFhzgwHkQMrS/UABC3QImR5BxA+TjHZDaLVgslFsf+ol
mZBBHGHqLUUGeRoNbrEnhFYAf5+ctrmY7HBppTpgYTXt1mZja51KIim04692kiq8852HZRhazjaY
TxGHFe8Vn4fp+vEFRjgHeP3pxemJRhilAZQUsG/0WTnBNBd7p/Lve25NTe6Pa7cCR6n9ZG7JQAon
r6glj8Xv590O8t4A6xgyIU61wsLfUgr7Kw8xc1XB9LoWvFuL3UStKyIpQqrG13vaJSn5T2XamsG9
U2ASxRpxwZjuqUv5AGA4y3HaYSbQbbiXm7tlCydEYo0y4Ehuyr20Y46NiSPRIWFT3s/KdSYpYSPB
slPFX29hReImP5tAojBkGbQS1SDNrSjDMqn+VzlJI2GM0um4ytmXtzGPadRBzxlGpSR/aofeNGBx
wRxgKEX/dWoO4zfQrIePUeLH7qNvmjGVOBGS5+m9h8taNxBtrIfWUW6dFEFVoYfdYxSHMEzqAozs
4iQW+AUi/K4F6IRrcdBjmezNaOW6EYVCo1sf/LcNEnSsVqqKX0lx2yjuJtnuXKlyH0Aq79aHuuLK
bej0t4PxN3rpx2ppnRWD+EJ1jjhfR082WGsWGYr3WxakNJsFNsGYlimfy44O72c/+yC8sx6AlPXB
OeARJ1zxli5MJXA+n+X6Rqgg4aQK5cvwEXw+/0o8FUjPowT57MsnRSQNVwr8JiB+L7iSACIKQTam
iMOZtLC6EMEn3p6pAdeoVQLiinxxxRTgHlh8JXk02AHHrDvO7YjwlStWoSwGVkDRd0wO79OBfvsT
TELko3qAt3iYrZ0a/pbuXgorp+BZEuY/QR0q4A/UXpE4VcT6i01ao1mkuygvLU8qtYqEUsn+hTNH
/5LQ55al5ERkLMdmtHrxUqV7+NbZ96WGZK6HQQu+rXCulGDp/9tYzqMa3/p57KAM8n1TudyqxlAs
MhfRHdl5bAUNdUhtKAs+E0lRL4hhzREV3TCmJHw1gitpPNvXeyifl08Wu100d+lvN4ji20vyyxRx
u7++bXbDBVxUzcrfbuQojdnCP6eZYYAB9BmHhL+w5deJmEfEwoBj5MKvVaAQwTJvs2OpUQ6Lo2DC
CuEISspK2z7kTVn7CrFQHwA7g0P8byNed51TVImpalhCesQXwy4+lLQKrazR2uHVbZwwCh/Nt5gh
lu0QBxyN70Q805PyeMnE9At1ZS+wVNdAsVZb51YF46uwbkqnnqp/tNgBnQ9YgRuGI885nz1/c3Mn
wq+543g/IJAqWpb7tViQwwNtpdpugj/UWR/Dh2MVJ/HSLm2NspWa92aIsld1yse5+nhbzHHUZaBX
FOSFxb1BjJPcGonJIOXBUjtrUiI23W5A+sGrNnvxtjl+8Ws4bSbvVFkrqBDH8SB6wmgxQYeYaPpk
zl1ahJAa/YxHgDNWvJHhlihBq5F5wc1ag0ZhVKOC5I/MkhnjvWhsT8J61zksn3WF23E29Zz4q3k6
nksXgO8ITL0mjSTuyotQLUdoULFX+pJ3uj27V2mjRps5pqy9OahV+5bdOKeCN7e/ukczVgwGihmf
F8DVg6EWBefGrI8tXeObFfIYEsfc0bKN6Bo977GkRnei7Ctx9RPgQdg2HCjYAd9nk/8+B8vn/HkD
D7+GkUgmhsgM/attffcDwcDmkQbOZHPlmsFXSUhCJVzKUXtBTRiUu0KbzOJE68V6NOGr440cJDkx
/WtzkQIw4LltgSabn3RtloTonmrRRb2kzFgxH26S3wNHBbBfEA2Oz5Gh8SiLGxYC8h+41fxQ5jK3
arzvyJShWmi1PuoZNdsaDYzLNQCMHlPJPtP9INrgNYX2FE+AkHJpochggTjCtrE7FndaZZQy4Sh9
O9va0dm3dfLZ50mi0mGcPrzPJRpSxlqRMHoP2qJZ2/Bad5+6OFewVd497ebBtb4QEv0Lt3OjS+Xn
xVfveD2ZAEJCgTi/uuPgS0F2FYCSixwkRwM5F5D4VSjFgltmQScZ3Q8tDm77gZ2eIjJc+eEt0tmU
EbRfzS3VF1tE1k+BpZsQMzfXJcbEidWgDpYjiNgKVHhTQDQ+7dw03NiEA4qdzpms/1CH0xBT1Aw3
TvS/L3w5hCdvbnLwtgalAd7aCp4NznFIEU2xVBvqs295ZVJ+DaxsXQouHQN2dfJqeT+CW+aMN/1c
4j1p+lLoeNMQAmajZz8Qi86Xahq47gZwqUFVqcZ94iYX1tdIBtrLZC6ef1UISxomcBZNZExrIF+d
D03GQJ5C0WfxB25wLWLzz0+nw3ZuB0FOkw6EZGijPqqpK4YILZn+o7m2g0/FRlScB8XFJLJiTcrY
hDyBJkFyzZxjA2k07IJfze51Gk9dhkPwZe8j9LBc/m8HbUp36Z2JOQgiKRjhtcezXk1G0DW0wWcw
HBP2+cXk0UAwkRiQxrU6PgO6QHyxSLJeJ22+Uw2aOF4Bx+HsqKjbqe7f8EGoynB+UQrVdBYBYBvO
5SColf9e36wX3fhKteh408N2R+TFaiFNnjZ1xcYYFBWVBBYeefKzJyJsJcM3C46b4NEcMzx3AkjZ
aXQY9ABVt9RV9UYgBPP6xXP+aYlKOdMGc6lM7QlDSNyrenZRdGrj0noGlym5chU3QNNd49qM20fO
u+0hFkpnzBisPklYDlZSScQ6TX+FBnoRmwyrSRJyP1tb68FwRNnZCQ+weFxTlR2CIcmFs7rV+ybg
j2okeSW07Mouw5cldEz9lPwLo8mh5wbyZ4SVrA8jcvkuqifQWLbQgBc+gn2b9rwkTtiCH3VYKMxO
fuyrQV3ascB2t4QKcyoFqzY7ve/+m9QOFFMeXLw2Yq3njOENxpvp2OWwKoL4TxkEBCZcKFzEj/li
jR/SserjCwQSRAxVyxDnko6sVhdMuq8ayYbQf7RnnRAZkVD8PQ+T1ZPd7XNTkxHIr/MY4mzPI32n
aWJrVOxqINEFPLxGZ6cSmoxaZ+z7D7hLWKAvENHlI5nJGVmNaX4j86fBKe65SeBBzEu31GbylpSQ
vrY2Wfs4srS4HajpSFJgDgoV10I2P0+cbisQxzP5eiHDOEVA8aw0U3Xnamxqcfc0i+3CVoTwXich
7PZbyLAC+8deX/tuiXmfVvej32H96FFdoSlC3vLYMk4s/HrOZAvAjylr96YoiLvxnpuoZdQK/bps
DCsPT9/OyapL0gCDMT3t+J6HSijm/kSMe1O5K3IuO5dm7+u1bNcXaucZ4cBw06vSZAkQTxFpUdDX
ia9dFLf0qQzI2oP9rp4H8J1jccGyxTgj6cctrsBo8Kg0GvODDz8faS4j02y3YNV+Xs0zkLYwuvOx
0InaJXCYjf6QqhkfnyQA1IEWfP7vKJJ6VUqeh5ZT5pt5jumwYCZnCmZ4HhwqIQjb3H1uq7T9GUI3
OmEA+OYAh8NBapshYP0rFX1RJvmJL/VElCjIH1d5VPgS7n6uGN4sjQJKLxkHzyvpKcuLut6XctGj
K6QOjVXoz9KUEkDk4wT194PdXzjvUUVKbNOC/Q6XzBDiHCme9cmaPm34Lb5Dl4HjtGa8UzRPP1LF
PakDUvcqT5DZZ1s2so+tyIbwVbw62yVhbpGjVNU3K8bHxPWBfOpg32Ex/2tI3PSJDzdkm54q088D
ezpI/0uSqJLDUztlKUxq2IYAILznCiZrAudasT3Th3PcReYYLDqaeyv/lQOrHeM4X7JVmw23HCTa
gOsPM4yA8cW77jdFIvm5Wr4kFU9ARd0BNalUtGUPRwv6fnpYK+y1XFEHOWdNtVR1g1Nof1L8we/i
mbkM17689717+8J2FtxDzHEkxFVR7EVHhnRFHK3A0lgFdPWNmE0qDiLaiaX+CVsZbYyfzHlBtO2h
au7cR2yfwX1FdyIvzHTbMSDd8oKdCEGxiDw8WwXxk+1/aV0/Ah1oDbfNzhGQ7PWBajt92Hhcva3j
FwIqoLDsFuUUSRdq+Igh6t9+d3veJNeYALfbbREoQip0j2dbH/elw9QQqguaHZ2ySushWcKtJvWR
sZ5Jt0Srm8c4p2exC0ThGDbKIrdRLyyYWr2AktOTWmUdNEuolYgZhcxqAFchu78ZAMAYDwtbeGSe
xoFoFlInAqZKdfSEBoC1zciatv0b+2NE777ZE9Cb2gJ4l9utvf4+0OvgqLnuAn5SaujyrlBoE+Ey
4Md9f/CvBGgbKK7vcQXHHbG/ISMOl5A0/X0k3cxEmWJYhiZ3+LoM96JYXtYX6d0EyBlQmHdOow8p
5M4bjcIofUj6pkxAlXsFkHmmcKDppJIpAhNmJCG+1SwufzKvYewxEePhtFKbOHp7EBG0UpwxtPz2
ibBV8wJ7dZL3J08ao2zFhQ55g1xKEd5sF7ZzrGXY+mv70IEFCEyFzAC4Ws5fJbeM6Sy1CLgBKfhy
LKZii11jvhhLVc/hhso/J5I6ZTZMCG7fk1dO4BpvEck85cO2LNkbPq6qUYil+4GsMEH3xp4Zk3za
8nvC7Ei0aXocGOwG4IXh2Oe75L4VJ0chHdfIMBikWMYtrkA8MVP889SipFjCl6eInl0MQuOf0QLG
OsyKStnxc2+Pes0FFCGGyzAO0/6URquF4TrUT9DyegWDhhsFofteyldXB4G0VMSkPfsIm/gxkKkD
vSQfZZjBfjyCVjutMFZa3PYZdAy3Zz7w+JsWp0jOeObRoyCUnQQ8eheqlranE9jqLbyryGJeU6TK
HzXsHuhqGoKRUGCaschBnObE9YQrO4sU0e6IqmW+VyebLM6IoQ97zZkLCC94h/iTbP585vSQAFc8
HOwDPdJcovMvQXeo+s/4VkxYB4YZSZWQ28iq8Egu1GyQ3b6VINEe/ukjhR4XVufZhPr5lXlOcKzv
VurOHfDeGw9bMpHy+1TpW5nNxSAvUzk7JN4WrwnfPn49IMlPsIV5PYE3K9s5Y8kVR2RFe59jYvfp
tymiwOlsBwN3TLmO8YR9vOHalhUqIm606C12XmI3jeBONWnXxgeH45+axNkc5UE9z8i5kiq/wvdX
2W88f7EUaAz9Sgfm9j4j9PRw2DDFcc1jqvsmEkUvq/BD7Zl+PzxbadgSbZHkjJL9cGqVoW0k3qF0
2KJZYyefq6l8xe1CbmbyxAVYeBpbVThxGnc6lPweyYCXQSe/jmFJf9XsEUZUjh4I1Re6Os8AUS6U
0KGEplgK13FoB6PDV8oWxTTzFArlgC3LGi7YsSfwPRSFlUOXjKl8B5/bJ3uFGyORQE/G4QaEZPsh
UFQ02Dc4SrEk9A98von2lvSi/cisQ3Xcg8IIClXoyziW6vxaT4dmxUX1AkMVIkqzvAk7QRE2gA5G
a4vTpYi1AqGXxz3EzB+ajrvaSwpRgbo71RUvhorBUOmZuf7O9C9MpWTm4NCO/0pignPovPnjKQts
YHs1XpyxRxDzZnZtEJauuUJi5TfkPigHM42uj7OIDLVBloPFpbqE/Evj7Oq5dfKTmUJcqc+DEdfJ
6V+ZlGS5PbJLvwCaAxUc5F9xdO4MWslDkGb3CSi3mfQFsZD+a9w0Eh4XKeKA+sOhByacsBaQwbTs
BhvdGeVQswNtNjlWLw47qx7aun2U0kRcxpWirt51Zee1b4nXT7EJ8eHqLRBjlQG5DI2sfLOB3NEx
tzX7a43TolUn0XAcI8fS6A3DMG5eAjQUBndRsO8ARWvg+c/9IE2LoHV6zLf2c+V2YL0Cvz+TNxbR
JixiZ3tEzUioUSy7jo7/aUZi99U/KNzsiwyzKFws7R1dpjTO7xLItQf2zDqVRq/NtWnsOD12Iy9a
N18DN3jBek9Ka/oLR0terGTXWhXcROo8wTXhuV0VVeYZ9Ks+po0qgSp1hPdShv2wSmm6uuvkpJva
FNJCp0pxWYWLa3q/BkoJRHbkfyiV3f57Jbmuzuw+wBl+rkTOw1fpyk/S33hk2CjUV2dCRP8Yossw
8iEx4ZACz8bIk+CkFVldg/4Xkhkp0smcHAvTIkA7l1DzXxxKqeyH/4mDaMKetwdY5HVCZUjC2hiw
t8nFqzpI4BbMfqgcyO37R/sdiHCPCOFouJcmN2V5mScj0g10Pv4EBTNfohv08rJzvSLwTFNCBr1L
5eaH/iVp1zJPHHtViFy9BHQ2LdiOOtcOCNoRBmosUSXXZUmUaQPQrF9jbDnZ7W2a9dluD1rGNTzJ
8HRUN+FJfq4P3DwbvPVLt1SH35F38Nj771Zf1H6BlhLnemDwb8rBhnjO1dgkxw0ieZy40BkN3GYi
nwXCwICY9ev+rp0qxGqo+bYn32E5+G1J38Q+UzileEDEmxjWSpE8MIOxxC16oZMGNkRPU2oA70np
3d1GtIzYZxcUAa6PubRW18Jt1wD0s9YvMXR00iBTI8I2ceXF+al1/YyurqXieMXdE+X97Xyo/LGF
DnYHWldSkEIZLKiDOwWznQds6VLfefrOXn+JfXeOQlijXReXdBdaapk77oXHNaneRp/QLfggVMvI
chlJfzKS0xUHetIjavRSqFPmeEyeqppU+ZthkLSW0oamRSGZlkpMWTUStkkMACAXh4J1eFfLaXoP
6FiAINw/jpn6R2DireLmhvQzjhZRXzQ17PNQ6WkgbOiBZQm4L65xujcdcSM+7dCdgH2XVFDm5gAc
QuXknFNazdUyewYjtmigeDdhPP4frYmZDNrdbxWHhUh/CNx54NkT1YIm23A/WjvNrmebHt3M4mOg
VS3t19gO/tX2OCz7uROadMw+0rvoQhuJufqHJ6V3NmC/aqmZLT684sDiwRq6wS/PtESB0e7uMgbF
GDClKuXVrUXllj8DJH5VntaGEUm09sOc29oAbtLyneaBbYVLilvN2LQD2BfhCueHnJyrdoyRRgIx
kSBs8/typQSVN7pUmvwz8/3vgzzPZx/RLPba4SHyurc3WZcFijQ/eHyddcVWhKNJ4PhWddX6t3ug
F3ReK6nbDM4sMUf/uLlGi3llUm8yzKgdUHogK6bDyhIiZmiVtGvzj+Loy1WOZyp/DdG7ZZ9PoTwQ
qluhILlWgtnGckHxuKG4Fqq4i9tck5Adu80p2zzzp6pD3CyWJpIyv2cjZ0eIH04jdTmOzKzyZaAe
utOZDXYhxwOol/0jKLKTO/5NuC5zh9wnTvzY3kCHPb5zHG04DFWPYCuIfNHixcWH3LiKq3hEhrTn
PJDLT2+6w2XenoisWNTgc+/ocboAxUbx6hd3sL20TTNz2HErCTm7mAXY6+ymHNbF/fX1/XysHpS7
Vze969i8CBuAw09TbXv/yeuldqqxSsZ9csbJ8hOdhhBCNUX2rhpuriT43A7ROo+fiwkdywuPu/r9
P8A2KP5E1fJBvOWi0YR+tc3u3rmlzuAHdPq64+B1yms1z3bkL8dWtIVeHlcygEO8fectljjugjug
aceeYhBdbajDw4Wh7+DRKNvEoPnwDmaH5vbV06NvsaNwNDqWcC3WLzirTKF4OkvZhaXJM/jQ3Xul
PyODM8pdBba6ZyP+B52Jv+D5+FBTJmnp/uw9FANCAfM=
`protect end_protected
