`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
sZ1VQQS667yHArlISgVYXZFY7DMWNVgJpwFqgwpgJIJkvO4jajBmk0Zq9HmDSX4xuPuqK9vqpzkv
oGr5zOGahJMaByLEsGCJe1X3Us5O3CQknXN8uzbpT+bVCDsYn29lzDtk9EC7U08Jh+MOH8xooF8C
rEi1rdDctDk3Ad6Cw3tYaFhlOrftyjVL28FWreOB8hDVe+hiRG9tOfTruaDXLnQXCZ2e9yJwnqa1
0v+5O1jOzW64e0Z2JUfJiKAV1dGVF2RCzuFMgETn0wLCooLJVGRKQ14I9z3BqcNmNB8JHSPE2/Ly
pk3DnqkNjgK1olr2Atzq434fayWgZxrlQrDPFg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="2c8kDpAj74/QYaojFD+RTelp2CQP9BvAwz1EBOEAYS8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1120)
`protect data_block
+tbmLRwNaRClLdY4/KlA63ZW6iLu2TUJjJpBlfT9UQU/0Gtvh8NnkhKO0axl29tPE+Mo4C474E3B
uSZcbyyxdf8gNiwRbkMaur0oaEEwpvs4RyDh4FxrtMibFNQLhwLws1NidwgP02c8XqRApoQKc7D9
3Pf7kqv5c1CuudnvoFkoYl4lemgLYd5D62n+irHgVk6xhgbu1itfnA3e7Qc/DPIHqmzQQVikUKPe
D6bZ4NJHC0VZCo1Ch/lWGBEPHaqfq3m4Kx0dM3T7cjJIenOoALYq3RAGULVS/OfvTCsDXO2PhTdL
oovDv+36WYC6jPHcDf+uuD5R74kVPzt/+zKF6zPhM1OSCmxOWvyHxSHHPhgK/xZVGT5PlQKCcvt/
luJ6nBep3TafvSj5oGt5I0N3kvq3778aB8JFFO6iI3IMiqShUYBqkSuIKgS5bEYiQL5iiY+G+8hY
CVZd+gnYgeHw9RKkhyWOb/zGtOiSo/samJniY1qIbQ37JfxJsH0uXQClSYhz6hC8zh+9W7XACV/L
/0JPzvdtcxmfMmPabNCx/Ha5xQYR6pFeeZg9OWoHxbKyIsQE0oCVIFXiRyVlKY7M2iYeJOPK+H65
JIhWdemLZGJ57J6J3xQUJFcic5MSvo7BMyvAPJrme1/UCOt4yZQsMhhiII8k9pRdqenlQq1aYHnZ
sx+NOggfYwukA3VozGdBX3l76Ig0w1m1RBMoiukM08khGOjSBLIt7febBtSPqyErwVPs8R0by7WP
Sn5uGTAYsO1m1tKOw0Mr2uhOxT7/IkiOd0vQeh7imc9Uq03LAP3pmR97RHcPpaCqeODLRgj1VLq5
esKOl9WSjscjaeHsBKoUt9fyfzd1KNSHBmUcrTseLS/DUQKlWnmRG+ZKjW2THFNBhMBcdhwNE/C8
A4MaBzPHRHJurLuymU7IolPRJMmNqLdQyaHa+i5KM6qW61o6pvkUkjQiZzFhWra3v74FX26568+0
1lJ8f/0l05Djc0jg4E0Xw21wvpjehtZEVqEKmXoGgyjMMEcZkvZ4vlAesQjq6gYhb5cvXtpTF0IM
HBHwDZoijyVTKhA5Fu7tt+B50N10/qn0jUtoSZ6dhiiBPWdvbDPK1DA3vThNxzqPnWL5s4sKmvi9
IueZeFrbacBjDiDbGKOusS9bmfBOCYDUYrub4PPTawGdZOW/T+Stj4IlcnrDV2IQT12FuwKfZGkm
JXUJTG43Kcj5jaz8X8Ewuo2HVJXeibLHhRejUI6bsiWJd2HyFd4YBEYJmgu7lFaDLnxC1Ex9KikO
BzbZNd5tscCB7t/XavRCh1uoCM+hEmSMdutAoWpXZFbdU0QhmN87XHzjK6GGpwchjIxxolsH8Omh
FYyCOheW+yQGAhhs1PRD87j9t/bJqra6ZyPnpWTbfVci3Iise5Fv/kB9pqAVYzI4dauOHVUs2i5+
s8Sn0J6Xykyc8aHWL1ECSVwjmzcBrqVbvyw2yAfQrvND6qYDUw==
`protect end_protected
