`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17472)
`protect data_block
KEvbFTfM82n0aNs3F9vXGOXN/twtSV8kJcMO5jkSZ0CPmt9z25DpVpj/cK1GBqP1blVx3wopd9jW
5dq0CX4tX6Tf+qPPS0evbUESSoYJFO2T5N+WIwP9++v6mEHlhhHiugQY3AkQl/WQGhLizNWsfgU3
YjieSkXcqxE343y3Sm1ggtSf6X8PGWckVL3wluRvbvMhJ/JTrlQfFl/BeycHF0wIKxQucIHmCE/n
hViRBvgRDzvH4YGf/8REN0562MJVsne3UwgDwijbAIldu90tG1cGgSF3ZLzE1oEXuZynFBzZMWbb
WXdE/44Jwvk7wMO3IXQapJn/BjoVmylNk/fTINqaT22hAtuCEQDw0CPqOntYFcnWG+M09uQv7LL/
PU7C94K666Ec4q8wRhzUm20zlMWOLhCTSGCfc1osgqdvXnNbYbunMb43Rm1Okg1vNRjf7IdJCOJM
vSj5e2TzkliLJJFsNohqbF0/v9/oqbP19cKeBdq0SPxoaQ/8h2qutMUtdjMXi/qcr4cEPqc9yDZH
VM2LoqvBNVC08OPx+fWX86urMa28ndmwQPrs1T8LvddhMgWvrEWbsAgZ/jqAOHl2vBo3mbo9Q9BF
geuDebCpsHvMOKz/pjsFWSh32WBh5jT8/FHZpG/hDer9H9+S9GR0PqiiVW5bAqiTqyS9u/9ALWve
qgJTgpV5BVm1wpnY7s9BKzSfi7m8W1GrsPE1ipW1mF6fXmbX82PHHNztTzabj7pbxX3Ay4d6Wd+S
2w4d7Y0meiizIH4o8kIAVv5/ZIFNP/ThfzOP3exMi9ZwPrLYDNofZTgxenUhGMu8M+tRrZOU9Kjm
5yTEmqLdhvLOEKxzLGDqeziwIQjzd9XRhH9EqBAYwcXUl771iqnNXU0/K9ThH1alWXrD3fmExPhI
zMe7qCWX9DJcOPcSqZzDTdiP9exMwQZh+1oGLMB2vtb2QccU+aLNT3XUW4/eRCZhiuECyjmzsM12
eKordaCuzzjtcEYGj/EPvGgcyz3GKWS7+n08uNNYPLktRrPrGg62vj9nlKJxtuZVmLFf1Q83sAJN
kum1DSW/eghkwHYvKxa5I2gpAkQRWsPKgyPrB6fCakWQXmqty4iWwt5BUnP9TYxJYNFVT+1OgM/h
8WrA+jnNzX9fxpBvRjtgtG7Hum0Jnwv/k4F1tgtlCWZrMlycsxf4eRZzy64qpLcBXqomBO8i1KbT
cz1ntOUqXakCYPo9EPjmeVSvvI/hb1ewNdDxU5e4WT+hpeIZ1DpR/P08Ps3uW6j33+bh6aQucs+d
RtH4gpzF6wcAzlBJK6vGK+K55U85v3MfSsQsZUVISnbjJx5fooOJBc85ONElai/GGALHyMUzfPsQ
xeYe3ETAwRjgvNXdkoKwkRimYKqYU6/dsNTLz9No0gPZytx2EaiQUmJHbVdLMm+SOYhr4M5j0TzM
SINEuqQ9+0N7PNWWzWYfW7sdMjkmp2ZbZGE42kh1NnCRIhJSn2bHeoaNAWv7IZ29JbUwVfHHqPXX
fq+5dJOb3DE5PARLpdYmo6vIb5QJGcq7v256CHSumGcB7tITKVr/6h/dVDHW3qUHrL0Un02usWm3
UtlLrr/k+Ogo9eRPA7eQOi1BoYFXBOn9PeN7x9HOaDjOBVjGjXHxXJS+SDziuOHKXNXv7iyPQ0KH
ePaIWPxRs4x/dJX59Tw91r6x6TjHpxLQLPZ6gkmei8YlE7c4567jecqk/VpQnl2e8Sdn9p3AA6ds
3iD1LNpoqM3l5wMCDd5BXbkvPAOk+JUX/Nv7W3eSzYj4xB0kR5WisLTYw+xYUCor3KWUJxqGyaNJ
9cN1JYbbMnMvHGO0143YkWL3FIbvSAuSRsUx7voTHQYiCX0Fa4hZwnMrnppCCjclvTi8yU+ucLiJ
Wz4yIyw/4vf40FY0756LY448JCv/VDv2lu/HP5ir53iKHmH6CDJNQ4Ert84KtKV8sG0CI57RyaF6
IHXycyqb5Y2jY0QY5fFSZgPkJwP9wOWXXJU1SQnTNsiJiWI0wCq1fAt/cAq2qAIomIflukVlXsw1
H7EpeGdbUAIU3DIg7DIpkVHRH5CSf052EvZCMZ6lieUhBlGSCzvTpbamYBFxQVScZvNmREdCbbiP
MiHbBZy8caY/xjz+R+mfoaNo7uCFZcfz+fGlBgYaxpTYLiRkgLamiuFZno3akXB6J9NfGfCMnLiS
hqH2EFycdDNYtQCqMucPaNBEXrz1SzjNJ/b+duZYvuzOqYOaulBLbEkEgfsDFFa1BGWJWjQQn3pF
4BoHUnuGeM12Xwb9sLBC8ui/gWrRcP21srnaSZeMSQ83d8u/FwLGdJBgdMlzJX5QPIGQQHFyFr2a
mQkpqRrshHlVmCuyQH0+yIFnvZtHXJbuVbWWWNc6o7K2wnpLSSjVz+kn4DkEymyarwmEdxKEKB+D
zRyTZz6JXMn8ViUgrwMk6/2/HHkSzNtdQkhOKGSUzbw1vHX6nu7YLv+x1QNP+hvPJKyqc9CHGcTK
MFfqTZE1Kw0OzqHzTb8T8ZUAXyAS4NqN6I0aRha/Z5vBAh3frA5O4utAihLC1CUcR3F9/W11MfPB
0WH9hVsmn3yOYyXXIvc62F+rUv2hmqh/MAv25B0XkioY6j7nZCKan8CU3BV/kkcTy1RtBpQzlQgV
b1EaKs6L+5JrMSbDAvx38iOfkSalBOpTC9QU3bXm+j2ibnPy35NP3ZVcK7E6tzykF2iYo/blHCd4
ckd3A4gOtDhirRcfdtbYjuzBljxpfvxNAkwzdlHdByQkD7fvGNuf+oJMVQTlGMFWN++HXDX0PPWw
GyyL3dC4WkySrn3KtoVeyl4fFf1oHpAYJDlb6cTDb34pfUW4CI5GgMunJ18n/GRngjsB7gVsP/rL
XAQnkjT7nU4oeOTDOxrKO6i7SqXvRJAeDHAHPlAvKE/AEQo4um5XVnGsRtiWIV87UVG/g96VPrdQ
5p38UhlSlo+pQIW8oLFbPUfsz+SBjugpPHpPtIhgmfVI3v1cmOItzy4Pi+U9rzXksLff8p+0fq90
P2pwTlYT3I4HqtYN9hPjldJRHzNle0EI6wpodQyeW16yfQ4krhddQoFnIkOotGiPJOID7ZG+PMBY
4Ya+FCAPH2uUc1KSYPESNGaf82glIjtOVBwJg49zkRgMDtrku10V1Cjn7iN1TrLLWizXOxsNg9i7
V3WyglDn2WI56qYMplcIA5KgvnG4DWRe6iBlUxRUW6n8RDls9W5HxKFqDBEso1VWP2iLCMKg580a
13wk/SRhwLj2b2vS0Kjb1tjS/AWq356PGpFveHw72qlQXWypIK+IoOGgwAcLtyNmvJgBUDTweFI5
lLg5AVMPok7vkBmnwLFdFDd6mlLBsbx6+vDDAvd26vTRa7fQpFnIerI46lTy133bANwqu+NS5T4x
eP2kHcNW0e1IS41336ChAvTm2pHcttDzYsTbBjdZpLsmSBsVhe9f4HNigJj5Op5zJSjj8Gz0O9J6
iHwP0mIPmHBxsFk9yAVW0sb1p8F6UfRkb6/53UD5U8fMr3bRNj/RwqVy4pep2li3WS4r2UnryHq+
EpIDhNexrmSyNEiixPR6v4fQ+3lv9ATw2LjnbyPekeAK1+DnHbIJx0ronfQSaxcUEjPv+d7viAlT
NwiorL0fWxFnDCy7iiinObNF8/ACDvZ/wGUhtl3pXoHlr7J6ikKh+w1LUVs3tTvgxzbuK7izopUc
Kr3berqxBkQPq6/ayhsBAh01ArHLWx23hTjI0c9MtGfEx4c6JK1BeD3A2agOMjmYZhULuqP+9ebE
Uy0CGOlrGNvXh17BlJo5BFFUnN52gUekJraLw8s7Qf6JV8pI9ojtifsylBNKj7lENMFeSEAGgWzJ
XNvoPXmxAphikIeq9cZ+6IrgzhpfvdOLbWYAqLIkAiIDH5pDMa57pIsNupiVgbPhKtV7+bdPqq9X
Iido6WkTcwpisxBQw4NFzclDrZ78eT3FJCKV3g/h5dFcXKsNmIY24pZ/gr3TcBvm8uIiK8VCtdVg
W+yhhIrxSbHIyoDTqqui2peC2+UaZ8n/qLARR6KWH9/GIsoPieIBxVr7Id024XB2eR9Yp5FdgYwc
DOpR3dA8yDmKqQkBWwms4k4Ct1OtADPLVMG8wY17C2i3k4EhR5uGgshxvfsRLhnv8UpJaVqpw9OD
IUXS1ZO9BD4tOrQy6xi6+7jYowUZS5GT3k0GIwiRHYn3+Lop1K64nOyGo0dreLeFyuFe2zMH/q8o
ZE3ngcJSNtIxSNDiG20zmLqmR+ZBPILre2mIFEMvcMirKJ6s3z7R93ZCEtIwN4zNnPhKUuZ/0vg4
Iq4m/QFehcDXrgocvomBcAPOqwI/5cYtymeYuIhG0QHa3+m0YDnYRVPWfEmLkZLcuiZqFr2Cjkrm
zdNuL9Kt1KKe2ej0agCwD32gIG1pOADd3H1D2MlEdS1zknCHhvq1fmTz5kFsjWMiLCmUdYc5OLKh
zZw82h4+hjUgYHtpXZsX2VrNxI2W/wnmwVBVI8lhFagWDcgCXyj54quVrGFKL/ep8QqNHBqyai9h
Ib6lfYviBkQYY3ykJXDggc64fQDO/+RWGRIVPOAQq2W89yUgB7wg97RBpkUN6hOjgdd3vCRMGZmi
I0pdo4ELPZn+cvxj8g2T0n3kDJyIq7KqeQpsplIeWYJflnSph2Ipt1Glx4q3/G9sgqYfs7ZiYN5Z
eonoUCJcVcpazZqlBnO2SSYt1ZyDVKjMSPNcY0GNWNv9AguqGGaX6Urvj5mRGPynXOsdlW4VUdAS
H+WzBgf20lo6pTZHKziFn5eVFSYcRqb2gtR+yW2FWz5FFZl4Sukmc+WYxKYIhJY1iwISwVJnxTmf
0jfTtzsa9My1DQBqrerCyGsthA1LEP6WFjNNlvp40moK5V+ECeZFeWJcZM1LLHOFZPULAngUBzq6
zahu4p0jN/gmZSf2lD1nCRgYTOy4w2iDMBJ72XPp3fz48EygW7yMT8DsZsYpb6nn1tOhs5T/ZUMr
7+5sCV2roOHh5TzoHN0jC4anFX3P3/Plnsm59RhA599VNZWNkN5MjtV+SY9a5MdeKd/urOeDM/dm
jN4dzfWrCLHlaWMAuCKRaMzTv/YYuOCalp1aj2q24VesiZFsZorm0CXl+CG2Ub7lOXN9xdllX51A
lK8iT+75APWkE9Kw0eS+nVO0phatF2/dgqg1xu+CuPXRrnx0p5iIh8lvpsZcAvc8l5a2wV1yZ6rj
x1b9iY3mFEDzl/oVgOVcxwP2LafCoQOwRlMG90UQOs3GIeef1cXKXuF7UcnJ6qSJg4JyyZhxc62Y
deduTXZ5in1IyI8ukgZl7q5jy9i/KCfA38103v6I/gnqoAWCPR+JBDtokjSnEnq2GQduL5Dakz5G
ge0dYiJRZ+yskulaqOmmIH92mRTOBQW8umPrrZcGp4n/P+3A9JR2RgL4US60t//zczHOwzgkK9Pj
G3+4XwrVxUBOH7aqll0CWkaVprQ/Gu4/qeatae5PUG6Ms233OkFF2ZkXt+06wAVCshC4Bp1ApZml
ZySC3XdqvH6lRCmm7niT0sJMGeaPiNFxxb2oemDfiGkZumMh/2NuW6TzibwWzqqEE3hmzB4db1IK
iGQKSzejikfk3vKSOMYzN+IlN47xyRbTssSjjdz6drXGAlqAugCzcbf0DdpHblnUM2F1Rd2BV+9x
mZfhVbu8tDp+eVk2NyrzmtbE4FJZFpsaYqtqT6EvtqLvh+zDsCm5pcoM0/B1sDdYnh6tv+n3+1vN
HytQf5N+sCmDr/RTw9iKVFe0WdKMNeTt5P1vmUthmmaXWCrMQmRGd0Tc4h/soYs7RIW4xwZn2NGa
A8gv7e2DPp4eOn/onCWzAWtREFkAWqT/AEeOjLcdfq8+Wsrb3MaWeKr8I13DtR4l1QvnYBynIATV
/iDZpR9LZuUq8GeFuXOnpGln4in/Ai4ZBhyQ1A5o6HJELS6BaMhUXhve2Xi+n4SdUGwmJLo67I0v
B4oVAD1VAs3S8eSecQNJYEIxxDKXvx05ZIrEwi9EYDrcu2aqUhSU1ify4GOspI138jzHGq80Ieqz
Ax+79CXV4W+VRt1amsPStIi0uEBnB0dWXlEdTowDdVlw5DZmIAtEvHcGiIj1foSbcyuY4P/PlNKb
h3frkN9jME+6Cs0fMq2mTdBrwzhGO55GQ84ux9wfDMNR5mkZkvDxvgXqn63soFzCQU9HH8UykJmt
mxkpSFqIHtulE8fA/rXkuFk1tcXRCIMqKNPuACiaOJdQ3mgDI+gJDufgt0kn2207VBeXY/L2ZobL
iXVJ2V1QOMxStu634rjViqRcTDJaoYc4JL2yYTfX+4skLUtNh1pRkK/D5aQnaQu/ZfmdJY9PUeqJ
yvFJs+olYYRFK+2I7wE1ayXsFJRT3+1+qIwnxEbCYlcVHACrX5gNdWYCbyilJFSnPLElz1JvGnm/
JUxkX5CNCnN8P77+4eEHy+L7rC621dpqF5LUCd37utDgHpulaKBpBoIgpdor/J1FTlY2/G+NzGEL
FR2Wsw1aDzw2ibHLUXuM505+qA3kSDlI/rdo2jBWD4hkqPYrkDUks86yuxkO+Re314Xl96pKJIho
QPilVD10u8Zysbm/YXNuIUuHg0KGGItcNQQhByYSX0PkLLvt/1pzS+TasF3qsHKoQ/qEyndCfq4H
bH7adl0hVysksGTSH4pmQZs3ApLbovX52Snmny8JgH7Ga/VmAqQrdQF9Kd0yWhiq5CwhGS+mpEUJ
/0coehJtaoiEm+6GS33l9Dv3GoQxQVczFQW84GGUvjctfBlb00YnusBHuZNRdGbJmSGsJX91LCcx
e5Z5KU2VoBfJz5mXwmPdKb+fop932xE6mUdqQnxnW8NPWCDlHtaFUIkfgfykt+knO1FF9EYQl5Nk
6qXqhapgu9t8MG9KQVfVZBQvz2wEaEFNrCZFjzD9dRO05/FkclGwHuIxuZvVi0Lx/7xlXvKCmNLZ
jqpUNhZKFTtGb5l35ZF9RPOy1cNAvzs+qM084bKQqWMu/rxxzLph6lmZI1OiJADOGv1CiQHbVixC
hz2CGCrttNMrLw5VTacCdZIFJJ3GnXKfD1AzDSadAIOwKeed47hGrmSK4YYul/uHeToRAnt3gMg5
pnLS+5RTHKQudyptvZzjzP838NjOLDZcQ4bcg4kkz7eIucgYMWQNCBHZDjf5JGG/LRyPMj/FThlE
PLoziNL9QdjE8nf2XpwqpiBeDxbpw5uvN73CG1VJc7TnEuBQa+VP3FYIBdoYC/zd5gSbMV44/zUs
jHAup2C3Y3VWVdVz2kdd+blR0y05G7l/2J0ALXXWRzT6GrAJ1XhlSKaofjniEVNT5tG+0j5SK/SJ
vX7+5z8ruWz4D5Mw/Fe+hzc6G4NqI+TzdtZtVlMqm+r8Ml4s2k5RONNht1iBgcBmMl8KrPMlv+Oc
tLGG4litVSdn69A9D3GOwhMxe2TP+iPgU2CnsGNLDOn7V/Jfv9rPd1vaFC2ZVjh5pmEhv1zNw/XZ
euYO+QxCiEhcJDwJ4vpRxXsUMWivz26XpfbOXjMILqYyxOdlmUideUyWalBm/HHlfdaBnTmzNab1
JXUK13gWfbpR9hdEJgRu3g+mczz7l5ozQZkPBGR6hQQ97LVTLIO1eoLCEK3ceIDKOuEyLri2x990
l30QHLNCeTcKgJB9ipCIJHe5nXC9+hLSwAtJzH+zSV+slS4jmt4xfM8HFs/3V9GnOZAy8wp0qVPQ
OafzuQW8L0ohvmYvRfKJFjv9yzZKUxIwBpluoN105EzjiVErgaF8pss9OD6SHIjYmVObzuit9Okj
JPYj7GJvbgtOgcCIR1a6/cSqUxZxIojyKen+OGVovG7pjQUdJ7JnZChiPugQvWB2Na4R2cMucciD
KULqS8Kg4V+KxWMBIMm4V4+XRAbIR2z28tJh0Evuez01OWPckz2pFjpnFBlKvCu8vrjNHZgR2Dec
OYKwxc3O6IAZhZLA1Tdnv/G6MsbUXb0sRTWo5TwXIL9Nq+amRjgZM2inQursIH+gQMfTFnoMkyhy
dzDw0AG7vEeNPsWKL42p54pvIUwGeT2+Kud1xoyEq9yxfWhXM3QaLgEL7T8o0II13QvoLDlbXoH0
kFDabJ9CuRBJGseKYfvAr8CfTpZ6ohKZ9r71UChZdZ43+rHvL67Q1aa3Jr2TvD0W+VUvwkFBlDXa
bALzDFkWyGOTgzDxfwOu283uMPCQVdV5IjOohsFFuQJNyyv2YCvr1D2y3s1kcZRk/rlWWeHwgEDm
upm8a9+M8E8Pk0MfTmwMBWT4QEB+v11gYDKiJM2+ZTRBJvPbTlKxAzsRiP0xmy10uuKwYPwPt/OK
ZEwbFFMgiGj4+RmrRKJP/1cB6vdToTerf3pSIPP6zkqrDiREj0JE46hZrNVoUYy+artXFiHOYuwq
PeSbJcybrfbMwgTWf4oRREP8yWKA5yt27TAmwZWGcTH9ClpoBSJ/FgAFwZob5RV5+gBfOJhpDHYM
EjxxWI2PHYeL9O3aY3C2+p5qHpP/E3xqbmyC7sADDZ6ECWeEryJfUsCk0vqudCoVJ8GwNRkRJ3LP
wHv1zQx22ckQKFAy32mWPG//4DBh1XLDuEooYWXd+sTKWomnwm3Hp4Tdm0xrxs9+Bcno0Yfxr7P7
IiZPpUgxQqD5B67jvPg0rjExTeZ6E4a/SK+/FbHK5XRKtaYylScgU8JfIlX0irOm0E/bsy4WDclV
TPT9yIZZLI28zvMmdASXVv3hWreKV8yLIivy78ikKAdSqtFcwnQFM4FX/L2DdYKgP5izkPwtip1k
YnH/uKsTbvphWy1c4lJ6cgfYBD7TS8KWE4iiDRMfa6jVC8G8KHIq/ev0AT+GYaLnarqbZ9uKdjIv
hPaLXC53LR40vrfviRq9rOr9s3QIw1dyVqYp47Jke1bqlZUfJuuWxvCrQHydqMHLDdaXMe63YpMw
A98boSkkwAhHDSgWp+le6QqRshtywOZ3zfSsOYiTj/x6+j4mgEv4CgL/kEkCvCaBB9D1tQocXdbm
FppJ6tkL9HxnTFQvNt/wrIhfFgnYHV49T8ciBu3UXwt4Ei27qHHCq8ypT3Jt8GmKSLSnan+MEf3K
h/A2xPipkN4F69HaxgyU6eTqZmVDcYqRUnChNawYQCFRCfl0e6cE+7QJhe1QnFu+Tw7p7PLgzkEr
RfGLfLtv6ds9P7SG9H3+uAGU3AWCbuqPV2xVcFmo9R9tW1zZXujcx6QE6gej6AO3L67l4t81pdvH
+XIsG3rcM14VfndMhXhynxf05g3A5zDebgdJzs7eYn4X/cp0WUlGCagCYbLaK5GCKn3zMgcrAd3i
q3++PorYCtSYnnuKdBKR6SpKfelB+aT3XxvDyGkAEXGM1vcsXeerP6XIff4LEGcb65wIM8FirSDW
EDRbhmdIejm++WUKVJy5WGQLwu2Q2CdUzulLmfq1dHz5JJTWKdjra2iW7JcL1DbaP6nem1bXHlgk
JDS6xfeEcCiH543V/QC67cRSVyTM1ChM+J8YqMhKVQdAvvEcBgC408YuuPzYmVUCHbM+NGDTSYj1
N3YDHSUH/ivbJvRQ8R/5OyrZiVuC1w/2tc3TE1HNZ+8f4O8d0A7P2J2gk4ehIhqlQRMtbDTaQDY+
9tEIALRF0RDX6nd3EpwJA/boEEnMQmJGBKCH7hWYhT2XN0y47KScXU3iW1j20s6AryS7/BNjuHSm
T1uJwUPL9LMrcIvF/S+Sgn98LLqtjoODSaVsaM5RYcrfrgIHC5v5JG9MDDq+c1bvldG27+PoubRZ
ThHYC2V0ynM2q+k3n8UPdrujmGIs8656mRtXSMjmEGHSHTjQEc3bJ0L3O+Kgd4o01PdQ9BJ46zgc
EvH37Jc1yTSpXfhZOy2WsI/2AoIvjPc9qbwlLPmKuWLgsX+QmFhOXPVfnxetCDjZzMe6RmxzUYFh
elX6BPSssWjhZxGZpaWg1gxhwhsKvpPqNQtXk8oG43F4MFeAuTl+j9TZqzBg0AnLzdWz2Jnw5PH5
DcVUltkgQL9ZIYtWhKw0a5FmR5PvJblLXPM0ueXZ5Le3TrxK43ercR3p3J+gcZGw+ZYc/+YCnLpv
ZrZaImIZ1PHONTt7tes3iEAwQAfp5dzu1kfFHloUCIqiNJWvoFv3O3ymdnJ38/BrLl0/OMMwkEzn
3HhyqcdH0/ln41qLh+NR5Oe/6jWAejCSnpJym/h5+VuGh2OiycK0EnOJ8Sx+2R2C49pmZvrTTKzI
iINTD4RRWgxSN7PnUTRAaf0Ax7R2XgG0WEDMve61iYeTERXYe42kEPjLHCMBbtajnejzRZeUnBpi
G/eOguPBTyiVsN8WMB/6E9s//Vz8ItM+q8ZTwHyYc8fDq0LuTj9tOC1syTAGAaDKiaBAl7inmKia
ImYzlhLGnozC+NRbgLOjCCJWgv0fESMqG5GrQJFORVg2e2/B9dRjpz4Ha/+CXXQtcpObWYQ2z5CX
httz7tu2fMpDmAaf875VIfnREwMHLtFmjOLzH6SD/uimnf5qtWwugPH4pXdABAwwHpdfpLP9akFF
TsBiQQB3qPX/Gl+IYq+u2Ovd18Jx9OLyEWkW/UizKtoczOpPXhyDdccBnIgw3B0RYuNWnGTHzBSK
6vUTstGKxdWEw0QrFw77q8MPhz/NBODfo5ldxXNqIJLKXxe8ehl61jXbQC3ZmpLitAmG+Vro34Qc
TFcKsKMYN//Rh0VQPhTbUgcghNKJMw6SljREMvA8+MQUVq1wVzqUFh4GlJ8yZ94XJ7u82CKO2nOE
bq3b121m/ZQ6vQlqtoDQwU30Y2bQd6FCHZYjkZBUaCajevk/amsZTFcW+JKwGNfpXy8DJ7gEfySq
6liKAjLdyOO6WQ5QGK/BvrZwIJkGY3n3ItpcP9Gy4HUe2ivH/K98hEBUXKfMcbW6sVAhXt14/Ygw
eJosy0+anYR8tEvZ2giLeqxOGk3nWEXHkym4Fz8ZO+OVf+Nk9rCZ4RXLHh74adIhc61OA2ls5PXt
erDrDEdDXf09WYGKSnn/VUru2bIQnmQHprMduzmgGvTMEcL1H9xAfu3f/KiJEOMIW1a9uvYSjIhm
uk5EONJUqmPOfUjoEHPZUY4JNpjOmSQgp0Yb1I509qkczIC1PolyipMRDclMigwRpknkG3VlO6JM
Q5CUouSapufXeBCYbsqtARIxJdwmlD76YdBHrcqajCu2qibWAluYgcwkdXBLiuVq292Yrx6hBrAj
6SlxrSZSK/FvnZ8RQhjoJTF1T/Jdv/mLvoBwbDHC+EqiCi9YldMnJZhsTjlNr6PrFrUzG3l/z3As
kC6mnFmm4smMSccXQ5Im1jOSs/ZpndasDjLnWHWOac6VLBe+fYlJUE9w9AbPdpnH/XJ1NJQKqkoa
aW+0ebwShC4L+i4gPRWdG4g/VTayu8AM2Mx67Ghgp4pbuwHbq6MclKr4Rnn0ZntXKgf1BP/fBXHD
mGmLimx5axNm59ixgiBwRTJnsW8y/SZspTUCjGOkh3dfExj9ryRHAbPXdFbhnavN+XNqHTM5a3R7
Z1gWnwRg8h56Mvn88RYSn8cBel/U6CmQzvhiaYhAHkgqfA5wNla3lKS0drAY80/yyR5vBv7BqDDx
KtHVygicmsEWklzSFMZ6co+eUiaUkLasXDdxGaCby/a1M2LJpiVskWLTo9BR7IlgBCYk9cG+NlFc
1cr2WZdoqak6SKPHMBi3K5DDlnGtef6WgwW3hKzM0qeh5XsVgSZGr+y4ZSgBGtGIduJVltQ6sOXf
/VYG9rJcnos/2rH64S86aQtri+nXj9jgQ6GLIDsssCMM+bfjjeM7W5MSw6VhuhNn1ImLT0QgevyZ
+fzjAV1QI6lH5g6THQMBR2ed6/b4yWqWsR86ZzgnJycHnmvikjXuQTHMOBf0M2kKieVjQmKVtwvq
V2o2y0g5QfofUeFGcK5wLWOUWo776GsckuA0CzbkN8wkigjIAZFesuRp1IXzUJpFLXjf4owpvJk4
k0IIkC4epcaTeJRBo4nvbVwJyLGlq+dR0MB1ZQhnTuD5PlndkUpUfuXu5y1sfrDztHQh1hsU1evA
Z12MH4yzPPOqsWiDr2KdUtDRE3zuDwhUtO5hd1IeccyyTHE1chpZdVh/EpGN88aWwadKcXBEkn6N
ANCtqAPG4Rrcal5g+xlAPyY8EeQau5N/YR3BghirEj7r1nRdVqqJ5yJsJThzhUEDSmNJc/nAyW5h
tFbuyZrd/tG1Hcc1GzJYJuOKdj/DYN4EFwOQx1wqDMgkWyV6yHX7FbaeWGR66R6Mm/uBcwtLUGF/
MCWnRpkr2bafLbvT59M2YG96JiRmrpjp8kCtN52E0iS9yhfbBW8xhk8eVXFV0HNmYyJjFvjOexq6
0nLqVNr+jCZlJYP+m2xH/51tAMsMBJbVlXcMcyfu6Zh8sOTlINc1+MqaYSWAU8ZSfiRTSo82kDjY
lFoFnDacYtWzoznteBkCQTNqBVD/HhC2pd6EjX5JW9Cdfjt9UW56kcL+waUIgYbWUEhNkcp0AhfN
5iYD6Gey1tcHVm+w9OU7KzfzxEsUF76xvdjbdIeIp5cvTB35+i4Xj5942RDfM8K1rJEhMbDsPg/K
YSnIMjDNqXYMax2CgrkBdN1oxNWgJqM/aIXgbMme4CYymMVqdVl9RR+ikpLCAGTTZ5XTql0mWFAq
1woOWdqh6wnLUEJaOKx2/F5DrfCxd+79oyAkutsi9/vmPROL9JgOwhfs5EcECInyVGOUPs2ZUyMA
R56RZwlAhjfNnNcZB5Hz8907M0nBnUCilrhISpImQf6j5b0+yFuJgwrTkqorS54GNZytRQx7MMm/
bhbGF+mozShr/1iWgH50fGBooxiw7r8ENCbDpymcqlZ8q9mBt20bdt3OzIVjDcl7gl1UPHB/m+tu
auFTDGsFeuzRcOOHPN78F8zGbH8sSio5POZ8vbGsr4Slti7fCYdDFucOwEqNKreJZE5Q6JH7+D2A
aqW1PCG1d+uhlfqjzKc1yXlpjoLbvgX+esTH73Yj3ScD5k6hOzI3qEp7UrBBrhDUSjHyiap4J0H6
ELOEnBQAsqoudn0bAAdlelzF0NxTHw0ijMNBmNMoNA0tZ3U5OwQJX5A6lkVo+YralTbdyrxdQd+l
u6zLosWBXXwq5zPHpjRfpicTTv7CDPFrUHg6m+y68JT4I9IUZ9BCd/ExUMEHkyv/SLrz/W6yWVPj
3/tNqElvOBZKv2AKBVFg0Rnx+PlmorrCOs5E2JUQ31/30AR2+TzIg8D4zNdH7I6JXq7A1YyuzBCd
4Ajwch4Ywqmz5Hb2AVY3iY29fXDXrBRZRM8UV6Jntn0rQtipZmPnB8suPcmh9xcyGFi7jgeLGrvM
66UDfSxhXDXaADA5HHteouDL84z/g6LrFNGD7/7PRsYyc+VmmpXQV2v7BDRQEMKcCYlMbs8m3zff
YKWNabopRdNPDPSviqmqFPeLxufgNMaHRy6hFLEyp3bZfdcOOlNBFMAEophufYF0BlrwlP0Qg8O0
5T06euUxIpvL3Ej086MOgUCaGriEdBq+Xr2o7uOzXdvT6wWdptMNpY3ewyovvcnFbs3Ryy8BKlhY
zQTl1YsGT4JZIaL0pKEfBwgYNkNVlFm+kdRFUboXcAVR38QtgU6kG/aw7yJfmzO7E1Szy6CXYuBe
YdBTAtQjf+d+Del4Rso03v/m0IMEf7hsvqS1g4Xp0B8Kti5UkHvNaxoRhB4mXW0zrm9GaQaFiVyn
avb8UHGNocf0pQQymYfU5smKOn9H6/Z7UGJrFtOciatyqhi17VhC6x7XVaZ+bWO1/1MZA1rTJwtt
cBwt93TQaSfGcU/6hUdzjga6ne0vTR86NQmZlAm00VGdI8oGWIp573mRO2w7es91/wDW7PHMujm5
5rXQXtChfNnj1N5xlPyqom6+x352EWmkxzNpE5SJXQ2ZeFsVYx9THESYE0pJDAevqV7hhNr1ZHl8
zIVnAbNjq+gBHOOpRrJZGbAX9Z0h8dUnv8SP7cPnBRZJStwKxymXCDoji4p92jUjsUzZdH6/QILB
0SCRYgo5tQOPSBhhedzfcVZqG45ZthAD5Vwm5n3kSqARAZBSTOuGRawDwiswdpqdKk8uIfG14nZz
QEzy/VGkmkDrHbAla2E35YTLycQB68+ytENwSTMYjrZ9h0SE4TfdLTdRcQkIvuO/8dm6jXeCLGFV
YdoUNG28DgXXtMccnaAkzG1XqTMLFzWvYccmP+mYbvN3BlEoAx+NTQqroBvWXfo8gi/qkVLyL51J
fYvAIkzppEmIjvz12s7gZW403kvOnmpGepRXubuX10WRZOTw2/RnVAi6qWa9HcaBTGaNE/6xDlkk
8aYimtcsKX5PeOOYJAI8hw4wheT26GOwUuN6Vh7L5VZ+fpfzNvfyRMcjSyXSZ2ECdbmMezl75m76
MUv+sYFF97IJqs5DW+w/NGoPS/QWVLLmLHvr0R0YQtkv9bBgX0GzYx3nVN7LBBuGTgLIS/jivchN
hkyh8a4ESqwXduu+hoeTTuHuEvHh3J0pOv/R8QdPEO8NyZPnjJNP9iemsoYu5nx3dOEiqACV1kHe
jyrC05oSQrDFa2rdLUvTn8KTPKSKhhX4JYh1qR3UQl37xq0+zpsXA8l9OFyc9VfRVp7AGr/FCEqd
gJNfew2NLsoI9bNB6sJF0nUIigcbD11Gm0z6eK/YA+GPlWTKpjupkEiz7+Of41zlUQXRZNZXv5yJ
FC//eeIML5gvhat/ttty0heCLdZpSqHO/DxumO+dHHx9ajo8zJZF6BOrYwiOp9JQWidhStlnYKYp
puxpYE3f75qvuV2nq+IcSeXNwjW9fm8iN2HQBkroLR18eq8bLsktG2mKNTYB+84zfrOGZ09x8rVo
paqM04OXhJ1iVNKcBRN5GwoAPe0DZt/K0V/4XMKjYhSsFxRH+MuOE30pFcdXFZGm62TFg2GxLv9L
VTAM2sEhqLT5KIS5Ni1L5YlanjgGG7flpUsac7HcBNW8EJsY5bphoLoYa8QfyyYAv22S9tmLkQko
2g2+46YLLMSVaJVBt+H/aApBkizfdzngrKG5NuNMT6LkbURBEC+GahuzzZIcY3O+ZE9q0mHbd9k4
66TRJiqeqQPZmyknPsRIJB0CHP5BWT70n4F9zvPIPxMrGt/p14N93xGr+CwB4l8HL/YIxSYfnYQ5
/3GQlTDLvCSGFMd2uz3C4+CvP/hySpNH6bRmmeCKT/WVy/gfwWAENvUFbedn0SjU0KULnw0mSKeY
+NQKA8MHa/uY1VPTb1KwYiVedUMGuIpjVFUd2y9zbrCQjFuSklMumm4GjRE2N0ZYiA9YqY1ZNImV
OKvQfsibGYb5b9Y+X8AYCBr1zl7BGf6ZwMguuRZA5rpmLw81s8t9mPnVxPEa0LN6xzLqSb40dpy4
PdlqH15wn945mnT7NrKvlGJ5izum0o/Z2ckjcTiT65ufQxYeb1d7/WxdM2WyCFanDB94vZNZbbP1
NBJYDLZ6SrdnvwPVfLTD1dQS2MfDeOPW+kBq/i5RH5cp2jMr0Rt3BkLAIp6eiGnruUtZb4p50kiL
neMwMbwnNKrHCiAzoYYtu5E+k67Ft4I4/4wykj1/a9lkq4ylgKj14gyb7sfDJKLH44KBToZSRx43
rRtRrc4yiBKpxzJGtkrM/z1mAQKYpjeFrCn+AkhgUn7iXUb12FeCZiQk505h9ZQ1Zf+wiZ+3l9bf
MjQz+j0IiOcYHx2y9nLyRWkvwHeevjLWFHoVetknopivqZTVc1LGVxocsiuuxNvybG5NIG1KMS2V
OIp0sAgtV4bUJvbBTRDDY2HrjhofQSErmRkI/BJc7cYN+A6jOvN2TfkD585pcfLv0HhrPUnEpaiU
uKRn31Ugu9o8k2l/9J87io8TbNAreETqQ9PhNNw1zFlwmoDWMdxPjNzktvLzqdPWx5OP3SBX3jcj
t5lfEB8WsOeGY67e0o9b7tz2sp6YFgB948VrufOPW5B+QstomUUh6Rns//U4IyjbDz9fWKXnWdP5
2DxHHV3sEOXQQu3KpdbYhg6y1UTwX5Ka0VC2+KqHPm7tKVtdwbEagXGnj+C8zNMexAOZfyFiov5w
dcz8PGBda7QjNCl7lLtTkJMsjNYXc76lY9JPah7W8DFB7MJxw+2jwqNCYY+FI+U8C/QHihP6r82G
AgiHahOitWuk78zHC88KWsBsICrRgTWwjcTwuMl5e28QUktoAQDeOk/p96jfSu2kWe9fx7x78YiB
mb0JoBm4/4DyzVyRKvlV0gpS9UFhwadBfZnRqSM6WOnmk5K4ZryAXPvD9RLQ7zhQ3Z7T1VRAqSpL
KBzTrPemw40a/65hba9cDPwx6beiy4x+C9ueoDPVCsbABAr4x3vmsEhkUD9VH6/kwS+jPhbPcSNb
E6TVsVcL3Pq/SHGmDvaGQpTi2Wny8A6UolgXITExWHFkIJhLBkPdRcyQYnulr8+1Q2N73gMTaUf4
O3UPIP552S8dkCVSp9ESBwzLXWJubwDpndpzWvVHMqUnuPSWlFjQCKG2MQPbZCKC23lWW2ZHBTLW
/8oG6ihdvC3Z2q+XrKZkQwFG3J7J/gLfJ8PR8P9MtS9Bf1+wg1s0lCZUWoAhwJ5vqZRI8vQ1jxkc
sMKGhklFDmQs3l8+ym0qDut4BgJj+K/0pLqyUoNlW8zgfmWPWNK/Z8Yy0mA3ukol8eJkp/c5k7sJ
AsF+qWyZfrmx6cCgLECMSwkQhGYZEnT64peke6FHXs75oryaYT/2ZQ28UYIGueOOXKXt2fMmMKON
oQiAtNO4nKemBBXB1GL8ge+1dTZIkoCxuprvWIP2z1As2rf79E1DDdvvbo0QngKRQBsck3y+dFv/
JekHD9QRbCYvhQwxYcpKZzzKbRKQUW3/ETaBylq8yn4lE7WaF1sTgOH+jpUE+GjKbNly6/zSb+Yr
+Y6rxHuuTywYg9DscXzROZsq+dq1lsmIagXyAFVBpLSYuIdHX9jZHWGq0eVyiAHUpRaca5abbgof
3xSrJqlhwC6W/f+zjrvaFhqro96RSo9uUT8c7PDMqjF9mwrZwy2C21CY+sCJKF3la3X2lPYySkJw
t1rtpxFmMAU//yTJ6TwL0d7qGJzKLbu34f0hMMg4DZSyhNi9zsoFkbsQDeXaMEkOVAwbxs7LZsg2
bKdmypellhC7bCen5RJP+cIOGPoMxajbzdFwCeaZkSPxzC/T+c90V2cY69WXgAvkMh4KMIZTbkt/
vYrSk5de9cr5AyAylaMbKsUkncBQnAStJYZ8u4UsOlGu0LF21dqKgmLVbjyqAH0jk/JTaPQUxrJa
XypK6bpvEkJNcfOlF4AExsA//BYkI8eUimsCMmt4vAkBrXZ6MftnZuW0ySWoxRAnVsoatmUL49ES
2lrDVD4BU4mWPI2fwohidUQVMLgFCF7gebfXyZlEP7Ae+TcOChMwiJnvrKY4ZgiHh0+dsfG/Hu9+
CojYbeDybtwLoWjN24qcbpu7owjPYfAbijl+HRwrAbX+IdSsQLUxAbKCmzmPU7jt5JQqKgL2BTCl
ZnBzChNF3fGgGw/aZZr+2SbB2GvrbT7GknY6UPPw+HIJAJ3JIM8G05KeZlZifbHAb39pMxym0BOS
XMbpfd9KakH+6VoOuiYIbSOoztqpfXw1jwKmM8GMctsrEJL2GVJObY9Q8FrXTT+GnV6HQn0Wshsr
0NyKPWBGwpLEW9ElzTfYppINOFAqiGHxKHCn3Mk6qJW+s6//DU96EZEcCJaB7FmgAUa2bMQ+1opK
GxPE4kJBRG4V8gd7z4nVCfBWHx8JFj+UORM2DItCbEIAeAa07uf7LtphfPP/WQIOy5daD/hLC3Ng
4F+uqhEiWkr4Qf2eKbjEYqyYzK5hC3/XpCeT6Bd9RDsjoU/EAfObRiLb8MgnHISisLxpMCS8QeDr
npZKj7ph55QryH7PWLV4AtvOjYpEKSysMnSwI5lkz2ReBe/qj2P0eskjeLbjA71WF1Dt6lx3rQof
8aH9Kn7WolpK0XJJIuDWPvICF6uDxLSpuqiXOnwYoXjW7w9h0OS2Ir1JnH9J9FPxhwtmB762di+K
I9UHElJSc5oEa7/j3zMs8kapKOIWKNMxnacbBB/ljslGqUEV2kJmW+u/Ioa5AXWdqi1GSt31gJdQ
oX3oEy1AeL5PXHN16b6TVYPDUKE52kkoKGL9hBWIjKBh1JvI2uqAE+r5XzTW8BmK0v1ImRDtnN5D
soGzEd8bN5n6s7tp7GBwc/oJNjPsOboXxg+XwkorQrOOUPc+kpWqIG9BgQ52K8BoQW9LluYwYuhl
zeFHhFKKOZ7dydW7R1TVchbSQ6gY4u6yWjtbErHWQvTmd0zbz/UUW/au5VpnX0RVSjR1V0dgEzfd
xfxGrzjtATzDA6/b52xz24W1Alm+rsz9FJJxFq2aj8fXv76wxJ/Dcgo3cs8UBhjrPT3svqpGHwvk
/qG0HFRFj6fslSODyqlwslPm4DyTAabGN3XNFH3GV06Iqah5LIyEyJODe9sebr1zbQR5aZvh90Vo
vji+R7l4HlrfrmMEmNs32BgeHYXeh2jTvw/xnwmqzXpsWGhfZ79JJ7wKXIpRC9JW9lcwvYauPi+t
NvJ/xJ2wdDyKJW99Ch4/du5LZxYCDkwTHUU+z8Tf1QlwJgyHcmrNEE+nda19MSvpzXRINvHawPeC
zVNlPgPaeNMty/h/8shBBmi2HWrAHPA0kusSfJP1Pw+Q1GT4QzRQ/NPkIgc3gMrmm7HNUXxLXY8f
jntqgD947WyqcVh3b9zHclCzgMmOCBRWtm1N1KSlJeEnpiWolGEMorcXi0U4z6M/rFoYOTWho6x0
wvJ4aPYPt/M1ZjXi2OpExcOYjxj+4WdI5UCekB9kZAJY71VpIjO7RFweB+YPKrjN62hImTjEpWOy
C3wPOQOIQYKEyajdvA9uH+OWLXOjJfX22gVg/hE8qOOKfRdcs1UEZoIRXQiUNVhP/cmEF67d1JI6
L/NSP1XBSgIflyAShOBZ4STEiibZsih5IZePUcr3mp0TfvPKEjBJjv8sbeEEHbIFKAbYrmS6+ZoI
mod9qU2i8Cg13FNOvMkdFz74MZP0H+rMaR08H0VVxLdJRYYop10GCVP874pvolzppIwoPbvnW6dQ
RPFBgfV1tTbupUzsy9EyKV0eVKr+DwMMff71g6JtMlJ0git0LQT20rIdx+o9Xl7ISu/y7U4AMl2k
4dEFjvzvaIZsr0x/0GacaFFk6lb8/868Pi95jZILI+04zaXl1nSwAyq21QPbKxu6j7c0mkPe3uUm
5PBwxXzDZA1wfOpVTfUNwArKB62XYZqJzPh7702ocJPF6i6apiN7l9lq9cTvbz8CO5/rsbMkMSje
mYaYNOzIEdJ5st+2b4I3i4nvzI4XeQ6+0Q2uSdYRGIZrJq21ci+rp5MOoE1cN482oWC78ZtD2pUe
rtos+t8IpkY4nc0tZYypUYa4stBwMbHPhXvBwsDW7LfRNF221jas4/AZC4PNeuRQXba02ueuIcLQ
DietR+LAFTXoKIsFClJxdyfzSaT9Jtc0zvvmgX4oGyAUQfdAvo0XVCwpkpSoXvce+1/NYtWWOTH3
TH+F67UROCwY9qxjmuhZ8FZzEwIU1sjOSKQgndmKCrGyklQtq+eC0CqRCiodMkxjviDcK4+aBYA2
pdAKFvEQuP199je/gHztiFIdqq7gPU1YXr225v6vBM/tsAdrufRUGLWYFmYO6p2PXEbfusG8h66z
xlklb6/ls5HG/yjXfEPLcibT64KQlwmtW4kcmFceUZE8rYsNTzGXdK5QCzEJpCgK1MgCUzLgs2Fh
3ia4T5AM+1IDKIj9+LVA6rvvFqL9eaIL9EsznedxjnzwL6+azbXbFl7ZvzKahWFMwUrMNJfta5jG
gnBOonJ6r7+oauWRknjKn3k/wnfXJ47Sud/2Uwncru5mx6Ja4iSydmkTcr5Wn34/xW9Q4ykNWRLR
93M94o/lcXnB5ix60c8WB+vk7Jr5AikMPOMsKlOxW64RadbuxosNveJdIQuJA+M9sRtMb4bovrH+
7mTLIsXHE/koGeJ9D02DkjwZtWRORjq0fpaRcnlN/dzeslSFHOU/YeVI/djKeAj0eeo9QTfu0kLG
59QOEoNw/z7RJ7EbqDvT02GIM9U6TtibrsDggbw4DLp6no/utrgEuCOndXNYZUUpn5S1JlxWninI
AGQmVwBAc1pvfcbFJfuXfNlpoJO9yu9jZWhi9isnchw2L1mBofMUiNy01KCHJjG3LyR3mwevK/Pg
71VGNCYefU3XBK+4TobztJpCIsBX8oGFk5Ps3gOVtOGDxj1Ds+ecEOJkG3nQDRPUN49Im8Fvgf2u
iz5Mah23Azclsg6FY+oULcVeoExGuMlfT2kCK2VhBUt1dgL0xLcwxKugpo3o4SagUYT3lMpV4LKn
Qr52HR+d7QL9M2hQPD2B1eINoXnte2p3xtXcTHMYeIYeVX2gHjr3sgOvp2v3AIIuUDFSVqgQ5pTW
FM1IlcQR8PNpyy7Q1Yu5MhLpOGIsIGcydQrKrraVQLF3y2UNe0D5UGMvrE8d086wDcNwo0kM6enx
zJG2B0Mtn5MITr8EyNVED3ISo7kgzEn6Jc+dpiezRfO9VhiQq0vhRge/9vywJ8JjVy5U8oL7GavX
hQiMPRhgtENXdPr5ULRMBbKVbNdhyuLb0B/kqH/b9jhzXUhD8pSzxB9+TGqq7UyWwhxJjrwq7HGZ
TzqnAWo/+KzjgiXwzH2v3ddSggzzV2bPXD6Ziu95kMN+tlWOudSYQZA2bBl1zOCh1u7bWqCurJ+d
fbHM4qbSILv3lj+lzviO99yff/c2jJGiFABoBVMDTYENEe4NGWtLomHfSCJiOuHtOWz+FOw3R9lS
2tzpbetef5txtZ4FoXOr3wPT2ABZSqoClisxe/0z/Gv604dT3yoCNVY+4Eq+E2uCoIW2vUtPbfZy
+rhF7DA2HpbAbvRWxTr8tPuKn0ZH/KaAm7HtMxy5wMoDgXFbO1Bw81Sga/7S8ZF+minUBXrbZlIF
0us1LlESB/s5SKmSC6w+k53v+dz/Hg882WDItMmGPlzUn7R2vDHJKgra+txUQmC6QwzvxOgsJZUe
+XplbHFRF6dabkEZSSaRKzX0VP2t5t4oDdZ5VXQ8XOfTv7Ou6cpWrJalUdrmoNVpRqXfAqp9lwHE
Sy/6+NrdgVBWThbJqrLl+fUN2gH+lmOSWvGdR7/qeICeZ2LtXIsRNc1ewDj6fRrSf1HWDLj+ft0J
rKN1G/nHWQGQS6P9cNgKXQCFQtJ1WRGitCBPb7KNlIQzSsche6DGtWxGsRqwSdvt90C0aQJwNqm6
6gvWLlRoU5ChmjHyAgifjvrLgw8GEe0Mc5+4evd6nwomGcbYTR3u0S+rcZocKy3kkY5NKtU4kOiO
1cJnifbkV4xsbPgfadOwyK0CZJv7/HZ+TYvFoLtYu14X2SstmCJvJZHkChqsYlEjjD9/Bal5Nwuv
Eq3EeHE24jeinaJMbXegxDy3Ec2cKX2eVtzYGggkKA6BqpE/A3YAOqVYS9eyLmAPvOqEPXR/ThQ9
CNMpJLw3Lsy2LZak7UXYFtizhOknSI0TKrVUlF7P4yJjzxMQhOAv3Ot49YwMTE+YodNcbf4KKCKO
GiraBGUUKcmfC9BKLZRXfrAqUOeiYFevsXYqkrzFAtFoMNT1ReiYV+c3OyEwxUTffEnx97gEsOyj
GctHLRKMLMfPCjO+171cW+8EJC1A19s5w9y8vcL1+YOVbw6ZJeHkKB5XIVnsG3/T9ZBihajv/dPT
7PQO+JbXj3m98lgor+EqW9Aq7nWnGDV8NcE/EsmrOp13dW8VKq0VqiJkmD6u7VFI8GsNpvpguKIG
JBT/l+ZmQNKvmn77zhkw+8mIE7F2QSgPgL/fESiNlSDYHx78u9uxr4zjgehtbXN9fZAW8cSkCzdJ
LovIF43BNKXQ3rCOvGCxlrrCcZVyLpt3Is9gAsh/QzjoXfUqYMmF+j1w1YYBn9dV6/yLDO+MVznO
niW8yh5O2XkmCJHRXxjB/gOzBKk+H+kfhe9b5XkG2tCeD37TJfjKi3ErdLKpBTZTEnizTG20fiC/
hVc3EBkElxCTsgzY95YyiUDr0xuQ3OnkcjSLlhGXZD06mLpIM3wMqB85jkq8daZIxwgZ/DmApHob
xxf3SzfStMyU2Et3ybRqkn/hYRCsovKHIJtocC9GOcDq6vZqZ40803kMTt8ySfuzJdKCh6pLHzrZ
eP3atfvYOUwYDuQf+Bq2HOCBKz/QL3qxZO0PFjSRmqUNabd2gZT18toBFAMIcOEoZx857Nt7LaTb
DlZFX5rR3rvpXEC9UoIVRcUQAOrbkx+5EhK69fYAQzRrctphhH+7/gK8SbDcPAF9pmgIGdBjDKDv
kE4y2Q92TcQipdnxzBm4VQ1w2xtbNJc/R3uLyywg2jxnlIu79ytFgv5Wv9rlMaRM+DzJd30WnUwd
b9vFoTZIwu3UoN8LWMaFPYGPtQZ54W6+VySlcLLfoMDnuXyHYPFDb4DcRbkkIFylKGs6eBNTEmQB
4E32i93Y8ZseP8UjPztZe9lvfgI4o8eCdg/MUQcA/eePW8dvLiWPhLNvmcMUXUvcDGcurxM6uv8P
7Y+ZHVO8NjuhHPK1fWGpjdzbdcFssgRosV93dWiWlq9OtMsYtAJFp3iNg4SGFwRF4/t+FVDy0oo4
C/NSAyXZ90EYFD+aCj8BmSBa41SOfyhaJ3lk3y8G3CvVmiypNeIzkcqwfTupZh+0lJsZ1Q03DjzV
DQM1HqnMXNqH+85jBkfqxmmf7JxhqftOdXXzy9z6xaTZPfygx0Kr8so0NoEFOnlOFfK2xz7e2b6b
7Pc2P1gnHE0f+nwjhHGftnqFXW7vGPJtY+6yio3ZSiJQvEokQzlcS0im+F2nh2HHMpePEdaTd72f
DPv2i3pEoNv7WmC6FAoiPADsU5m3L+k//9s/Pxl37yxyW75O/Z0fWiZFnK/nmXN9LR9pmWjHxvMS
kdXbBBdFkkvt2UbKFFu8V1vcQERl52I4P83gams5i+hWD3KDEvJLZVzr9RgVgGdDPEppRiUhjDSw
4J28oAl1MqIrdYv/G/BKCHNh8E1E0XdUys1lDYhzB2MnoDzPxP3zWYcCqTzkG64+V75XYlJ1yZwY
BWisv8w51JhXghTL0VhQcd0sW5960ygaAXLeRo+YSEs5k+Wx4qkgNFszzIKxNwdsj5taFN6saWe7
xCZcH/6JtvFpAWOwOMq1gUXMZvGPJUKII+leWJSL
`protect end_protected
