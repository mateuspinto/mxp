��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���V���hS���kAk!�����tB���g�s��9���AzP;�|�"Xκ`���L�JJ���A}�Dg!�B����$���p���0|�:\�#�GcpqO2?�ȹ�ь�ѕu{
�l��>I��7�m�]���WN#\�a�e�~�"��A�����D�I�Z��
w�e�)��^of|3]|$Y�1�Z)>R��s0c|�9��6<��-�H��w�4ѹR�vٻyI���~M�.���>�N�̣X؇��ؓ�f���ԃ�$nAɒ��+������X��1�zMi<�@��[	�׾a�u�F���UX	+'����B�1mK��c�����=�݁�Ǻ���o��^B��'�,�"�⊶x߅�}�/\(Z[�D��!���)L�6�`�����Z<���,��P�IV޳����J4$�8����)��3�X���Ϫbɛ��F����|�i�'Ӈ��6LI�WOQb_%$?�����`�Z:�:�� Jѵ�e)��(������x��\o��C)a)��0#��t�l�Z��2�!w�f�P�F�u���n!�xJ��>2�X\S"4I��Ңw`7;��<�]�d.X
tR��M&X�^�Bt�ˉ㦄�=��AҋV�d��$᭾�a[�şb�j >e��?`�N#o�S�v ��1n4��7�"\!{�I�@��iT�p7w�Ҫ��~ d�q�ۯN1�M�膠.��1��}<SW���E�fFdi=Rdj�w[�C�k�D�˥��r�����V��ªW�߀��w �m�2�o�-V0t��C��EX'�,sѶ�0}�Z8���P3ȴ��.�qp�6ݩ]R�i�P_�A'+��r�9A�xW�F;L&�ܤ&�qbH�r�X�dҊ�@HW��F�>�KQ��(e%�c#kv|�r����B��V^J��A_��/��@�r�VY4��G{�>(��z�Տ"�f�>�>�6Q���w9̅��޻���h"l�|�$Mgva�:ݤ��d�%�\Θ 1���������)r�K����	k_�F���]EC��/j�8,� d^�t!�L��Н́E\3 �˸�P���an�Hm��z��jG��6��{d�ˇ���	�l�	,��+F��[��fD�!��f����kQ�~���+3�i1�M�94�Kgﮊ�,���k�7��B/�9T��lmcJ0�G=��j9d
�*���-��^M�P�;b��BkZ�	���
#���b�h_��ٱ%���Ȉ�&g_�6C���-�):Hw����@7�F+���|o�A䀃�����0�O�[��ޛ(�A�\tf�v�(9�!"t:���'�r�]���q�!�iΫ6���po&-/=��S�3�3B騪�]�J�z��jͮ��8�ʶR���	���$!�^#@�����^~��X�o+|��F�j/Ru�� ��(T��+@+*O�9]H�q����;8\�t3&3QF���	�Ĝ^�H����u���3)��=�ɼ��$�����I�̳�qv��?�R���U[3��M��ι)'De5���n�m�� �9���Ė|�X��B<��	�����*ܓ{�[��H���W7�Vz)�&Y�0h�~*�ʝ��5��P��P�@H�;<!��� :i�	KBZaL��*���\��]�4J���9q����9��M���L�9�$F���>����W���_ۗ2�I�R�7��Ê%���C��*�y6u<�}v�
���v'Ǣ^�Y�c�h�q#Tɇ��&�-K�[���2���!�|Xq^��dp����X̆qz2�PqR�7������&�}��Wx�w�N	h�5V��ǎ�WvDէ�P�D���8�텟�@��L��oz�3(�G����j�C-ӸX�c�g̏�����>a�PJ~9�j׹%Q�˺�E�C!�S����o�:���љ���ȓ�c�	"�����ILۄ0}?ܤ��1q�/gK���ӈ����5VN�d��A�R�-����%��Q�?���K��iOC�����[�����u���|Vġ)���\c�xE�K��\�( �(��x(V�9���2鿜�)ߑ��� �n?
���I���Z}�<��n@�g��Am�[�f"�l!�Eg3_��d��t�����hӋܤ)Ի�R�~C�n�Y<�yX%�%s©�ѿ�S��̀��(�jr���hi����̠�u���;�4���#P��"��tm��oұ��XC�KoO�H}��E7�G�S����%QʲnB�y�y* �b+4����r��ۜ�Qpj�ׇ��ئc4��E��3椺F�
u�9׻
܆��'�]��t�tV�*�[8-r����D\7�L��'E
�����N���,�B{��_�:v�����PȞ�5��j�] Q�:�!U`�p7i�$U��?�N�����ab�����ů������>��Y��P��]�ީ���G�&�̊p�?h|#_��v���F�N��q��Ë�<��1�Qg��:u���V2���bQ�Hd����5�m�2���Ү�$���D�tQl�ۃ��x���=pO�n��oC�=�3����PD4"6�:�����)R�l&�8%��n�˿�~+*l	��;?�4#�� dA�[�\�=��F�S��n����P�1�8tIc��=m��P�ь��
���T�l���%�E����*��f9|i#��� 0�0L0�x-;p
����5ȅzv1t������uB|�r�3D�g�Ω}I�=���D̩aԾ���q�?����l�J�y���m.�ES /�Z�"-���pZ�@��<�5�:���ߗkj+�u��V�^n�n���x �Ga��[�v��,ܾrY+:v��k�|!Ct�/F����O ��[��F�y��O��'7J�>�D��q;�1��z�ĩ�A>-UB�4#_�0H�6F���)��%�1����HWT�;x@�j=}:�+`��ÑM\N���3��NDc��j�vEE_�'���%zN���ϋ~�BI�Q�}�T�L�w��Ra.c��r�d=W����o��m��tK��(J˰��\;��[��J�7{��Q���R���ðm�����?@���7ǌ ���w���.�� ��"��z0�k-yM~'�h
����xU�8�7׏w]�ޙ��ߛeC@�/�{:� ��Z ��;JP?y1��6����ӎ��PXQ�|��5#Yh���c1��RJ�����Ng:?���Tf�c#?CQF�s$��W�^��q6W��Yi8�|هN�*����U��O���a4�t|Z"'K*��1{{y�v��4	�t�+iۗ��g�ݹ����R@�O��-��@��� ���Z~�O6��� ,ri�Yߌ��90^�
88j:�O�ӄ;l��^����[�V �TI��O	�͉l��AZE�ehE`1�C��;9(��A�e�P�nč�g�[�dV��т��B���dguI���+ |��1.�᎘:�����T.F��=�ӿ��I�C��Jߥc���Cl���yz�j
�C���9�6p(N��t����F�H(��h�!Ձ�s�ӛlG�h�#�u]\���<B���%B�5�n�B�0�t=�0�;�Y
2�+Ѩ�{���#���[��<|)���#��<���fU	�|yS����˂<tO�š�z����_"��l����T�8m!���� }PkD4J�����u}�M���q�*	�C�Qj�Z�a=�_�2!\�;���ԧ׿��m�����oi�u?��9H�U�5g����یGص4��$I(��!۲�ۘ�]�yd:��HY����K9����v�T�w���$	e�58�����^�7i��$Z1e�A�Y�.�+��GC�,vFFk,����:�ԝ�}�\>e��;d�ssB��Z �o�Gxw_Z9*:�~Wj�	@X7����v�Du�7<je�9[�	�);J��d[�>y�d�1��H.EX��hD4q�IyL����GNl� :����ʭ �,(`��'�.s�>-;�<�%#���Xr�}3��P��Xr��"�g8�GY` -�ݍQ��M�眒b �y��<�D8T5^�%��κ���ȴ��4Ė��h�)���ڞ>!md��T��,���߬�u�LH0)�ٙ�2���9O�!�`�m1���I*��@T�`*]-�"����Ć2�汎22��W`ӼU��/\�$ZW%5��y���(x-s���NZn		��z?���+�ϻ�.�H�Qs�G����i�úYu�˂0�k��q���#gB�Gr�V`���f���$%,ro8.��A�l���j��\�%R��l<'_�X�\�����k����R�1����9����2o�de�a)f�����P�]J�[ѿ��z��w�f;+�����<Є9��&�`��O܎�x�wز����]�+���A�V���4Ϛ>P��x��m�gv~h�c�� -�/`̧������W@��"�ޕ�f�Dt,+�E��~m�MV�#6 7o��(�;����z�G�D_�O+��k��ꃲ���	��{�������b[�b�u��-s�H��:����[���
2�..����=t�ᷫ1e*D�ǩ���y�1�M��{���\�%�8ܮ/��_���u���L�_�&�ھ�=Xً�D�v�y���YFNˡ�������ɀ�64,��3ğ�kO�%���ޜk|HѻL�:[o�Y��<TupB��?�Ӎ���ʔ�7����onn��Ƭ�a@bC�fHt�e�oC	u��]�T�X�[?�Nt�����`���ҒR�m	��M!+�����5:}�L`��AF�Z�v�q�����ΧT�Z�@��$��,['�y0f;�Z[Yj�:Ũ��B��Q���&)Ufo�?�%�Y�V����Q��dG�L�~�>a"_K����V����w��6| 3)͵���)_�Aپk}�o��l��F���t�1~L �@Z�J���8�p���'�}�a� a'�86�	z��M���fų˄0��6�w��gꂉɄa�nV
�=��"�H�HS�a�A���l�Shc{P[�8��B��x|��}Ҕ��˪`����l����[>� ⷀ��$`e8X?����.���媣��ia����^I��%=��9lk|"$[�����wD����a&�:p�.Z称�S�W6�Sm�ܕ�����6���;����I�qG��
"x;`ʶ��lԓ�9&[�����8��AFZ�q���LS�X<���]Ud��<y>����p�r��A^&&�aI����{+��1C��=�Xi���OSfA'��5A���w�<!+�7Ӣ5T�d���{�����0KFY֞_'��z6����U5���-U��e7��uI���r}� E,@��R�N�ib=�감*����AM��pҺz^Y�nMhtV�^��	���6`��m�����s�VO���)|�M�t�"�%=�o�`�R����k���#��<� b�3uζ����ɟ�?�IDըُd�7I��ǡ@���N�!��2y�?8�qj���n�l�od�I��ORX��@k"*I;7�uaZ\�Ag���4M_#`��`$2�0�&QƞXK�M��!�>
�IRc-�c�b��'w���k��<��� ������kLsO=����q���>�t%���z$�DJ+�/��NR����?o��$�n%��1��NJ�8�;�[Ԯ��I�[�t��+1���D�/C�r���
�|�6f��_�x1��0��#�}b�ǻ*q0�V_ KO��YL#�����《�wuo�w,!'��"D-�)	|Y`cz.!��:?cwm��UԖ˳��3FP���HCb2���T�ۿ�ˊU̓���Ț9�X�(��>'�@(횸d���.�t��h���9���,�V�o�sB�R_���Z�(*�"*S�1KB+D����4�'���b:�Kc+oPiM���1��lkeo�)�#��H��K�S�G��(5���v��Q��>���M�Ū������b~�8�p0�|��ڧ�Y���17���s��q=v���e^�.ib�,e����cS���Nّ|yh�P<8
�n���у�+]������/��AK�x-ӛ����x0��(�oȻg7U��/+��B�G,:<�y5���tu˒�
Z�����oO.�7��#����%+��ˑj7u#���1��'H�Tx�����G/��D��y6ZWR4r�`yWcYϼ�E��;Y�>nF�┙��:o���
�۰�m����I�_�jY����>���&����/<�%����E�H��uP:S�B2>��G*�5r�/���w��{�З���+_�,��A�u���O"�/�(u3�IJ���{��bki�^�@�u��i��� ���B�y!�H^o�Yq��v4QX�aX�B�G�����f#Ӛ^ַ#���Z�ă�����I��m���(Q6{�����OJ�k�96S�\y���h�_}dG�o��_G�s u~f����';��@ޱ����	̍o�@��)�`��ޗ�q�0J��ӅA�Ք(���ΐ�l�H��ymQS��A�CW�b�3�]W���|��>p�	�UD��2zᨷ ߡ������	��xM_}��!Ƨ�rB�����Hٷ���w��Iu�f;6N�%<�?"�j��*� +~"���9h���ǻ�Ÿ+^����kY����q�VE5P஍n� pMv�����]�dk��T�֙_���9�^��N�o6J���:�i�D����0g��>�)Y� ����	��м���_�{y�<(l5��gX�;�:��@�b&��q���i�YR5�D����Pb�h;�&���"��5|������3=r�yʏ-������Era�24�3�@w[}ˬ��;���]`TJ�0}�`�L�6g�M����A��۬�?İl�0T�
Z����F��M