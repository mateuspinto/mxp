��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���`G}Ftv��1��rN^đO0V�j9nE��UQ���2����\*�y
r4! Y�����{a���6k���m���J�� ����Y�u��i��� �|��tv��_E��I��6�_\0}�
����g���Vq��$��Y�3|** ��Z��}��E���GH��_�L�@�@����,�V�Ǔ�1	��~��z��0�� P�Q�!�p���&s��m!�z��r}=(�;��JZMՋ�5 �����	���6�ˇ�]	�b	��c���:��̉�?P)���Mm>��x���+[��MݮD���Z=�&]�Z����%N2G='�j:,�7����\�)d�B��\93βV��4j��{��2�������Iɉi��Z8���_{���3�:5{��F�*��˅%Iv=�e%�������������h��e�?0���e����B�I���ly����[C���~����������o�!$���M�kb����D�1�	�?�l/�NH�>�B�U���5�Mi����2���� ��q?~�}�c�r�D},�AGث�
����ԭ����+2mr�X���y���P`��W!��!�3Ǌ��n��ժ�u9��B��3����A���1{)>ŉ�.|Eq#��q��=��iu��~��R%�0�R�#ō�r���c>2*l��ѩ<t��LC�3��m
�	ԩa��&�n���@e-qD��r�]:�W�����j��W�Z[�&��q�&JEhL�]�	�m�$�(�@r+K��ˉ�B��D����dLJ��|C ���`��*�~���h͘��=7�hx���<�&��*�hh'7�����O>;K�&�wcƐ�>ӂ���c�*ˈr�%��� u�=Y�/�@n\M9B���8-Y����ɷ�',Q$nb�#`A"�LgٕĴ	�H�by| ����Q>���ʈ���R��>�``9��$��(�s��_ѓ�����f�(����\w��}xy)��Y��fp���0hHzz��;��x��ԻI���p�I�:�C:���N�U6���^�"4}9>~u0C$�'�� �$�Bh���}_���	f7�"��`U����y��a���Yd�M�0�F��h�{ųm%���X�&]�o:.�m� ���H&��i&�F��K�H2��q�?	|� ����{�����p��e~D�:��s
q
�Z+�k�'�V>�Q����m���r��I#7��Kp�:����D���y�D��Ò�%��$>�˳z����Ň�I§o6����� ��=���Q-�|�NM �s�AE��N>7�A�W?z�%���L�����˔�������=�$N���?�]i*#�+����;Z����M贳jh�2'�g��'L���^=���$�,�&�����֊]Y����q=p�����TK��@ڜ��hؙ��Zj��u�+&-m,�4��v=�J�+�s\~����R�s�FNPe��fՈX
���Ǩ��d���ikB����G )y��5��"t崵�)�91��B]A!�k+�"�g��O��n{3�s�ʣq˯�N�o;�IP��{l�s�z��J���d��#Xf>��O�.���3<n��W/��Q�$�RX��� ����.��h�Ri9w�ݍ��x�����(�+�E�8�1��)^����Htˣ�����(Ͻ��)��od�(4���!&I���Mw��䒠qY�y������z狷�?53�M������l�Q/8�M��A$���-��
��cQ�W&�<�FZ��M�?��z��
�QC�HL�#��'LX�ۼ+^�? ��1�;~H@)��>����3�]��|-ሡz��D��A���&�P��N��?�Qd�Q��S�����b���p����䒑�b�2ZN�@L�/�KW�>�T����O�m<�9�7W6�7g	��b���h�e3{r�k��	%r`ώM/\/����J��=�y���8�;������En��Z�����cu4��_���Z4cQ�c���i&1(䋪��imà��T��p��x1%N�@QU�_tڌ�*R��+�v���H�#��4ѓ�U�B�v�
|?�L��r��Rz|6On1e(PXW{�ZR�����qf�j4M�!g�*�0�!�,l�뗨̨�R�;��G� �dޣ������
5�Դ�����צ�ye��y��rV'�E�����(��'=����@�1�L���X���ӎ��vw���͒��'7�*�T��5!o�d̐e�v� x������Q�2��W&�;��R��Vp̱���v�����/7�Suq�蔍U��R��|�Z�2q�*r� �Z.��YI���m[_i������|��VS�wB���~�\�L�B0(��В��T�_ۦ��������F�n,YW_��5���)�nJO����׌�g5	� ��-k���y��N�^����m�G����<Po�Ģt��m<GOЬ��+t��0�z`Qb��eΠ������/`��F�<��X�
�(e�l%�-|��X4�%��-�֣REIc\ڎ∫�"O��{����I)�F/��&G)ؤ�T�BL/y ���#�8�.�����/���=v?�{���쵒�ȴl6�a7�'8�ؘ�1`�M#ʁ��|D��fW�s����kBKD�+�[\�G~߱�3���d�[ aS%2�)9V6���}��j��i�	���)��W����~�]��#��ײ�2�>���|3�n�n9�������7�E�m�����Ґ����R�%-6v����� hg����M�/;���+�et^���H*�j�=�'t{9��X��;��4Q�A�fI�d�;y�k���2<����N�rM��g�_���鍿���o�c�
��h���ےW���.��rb��2�&�7.�$�v���KZQG�.�&������7��[��lfٙ'֜��_;��:�