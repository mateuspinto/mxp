XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ߙ�|z�ubd�S`[|b���d�u�at�� m����(�Ϣ��|�W�/X9����B8bd�+(�q�B"�z����Y=j���̻�)ZP���X�Wf���������5���l���ݣm�n4-�2�n!�z�����t��auZ�$��ka�W^s�A���"�C�`K��L�7�T�a�r����P��}��y@?��>���x���,	�Gv�w}����&�P�ϼ �yN�Mb ��W����#7X��ԯx��j�a@q�V,��Sҽ�h���@({h*Q���v1�q=�;o~wW1�tX���z�nܱ�7�t�T���o`�^ �z�Z���=z�WK9����K3��A��`^+���u癪���L���6��`�W�1n�7�j�b��g�%�u�(z�9-߄T�yg�:�Y���(U����Y	�'�yĽ�S��)?w��OD��o�Ss�"�)�Y�gO�G�J�d8 ��j�"�Yx�����cp]Wm�|�9�	�`��F@e��%	\5ZD�w��)-�p�@��0M�숝�N/�ZR9}�Et�*a��V,��]�y~�+�!�^$�s+��Q�q`D�k�����ݿD�)�/1�ՄW��Kr��~I�V�m���Aa���-cR� �e�p1/�E�t��si��ږ� �:*���I깍�H��́��խ�G���(P��@V��cB�ҽ5��RS*[��K�۝g5MT7�_No����&�!��j��ȇ����M�F2H�KJ���̡�\��ė;XlxVHYEB     400     1c0��K>h���.��&�V���ȗ�����dV.VU��i����
n���h�
V�+x��d�T�R����%Eqs*	�kT�hz�� ��s�!*uw���}d�4���x$&;� �	�Us\��z�
�uD��&�6UL��=X|8�)�-��՟`���B�' ��E(?�f����63tK)�|�v!��f��7��^�Yr��w�BԸ71N�(׈�q9�M�֫��� \�.�Nڝ��M�"��7n0H�G�]SW�/5����!��:<z�M���R�#8�_�(-�V|����q.f�yVVNg���0�����V)ɏ�����[g�f|�Ȥ^�yH���2���]|}�h�7O ���8�[5�qH-ؘ����~�-��!1+�������t��v|���?����.��8�^+=ɶ3༯�~e��B_aXlxVHYEB     212      d0���DŰ��;=�ƔZn��(�	M�R�Tr8G��������^�W����J��{!^I�J&�0�e@��^�ť0{g�T3��!����� �����A��_J̉.�8�q(������U�������O��b9E��+����IO�4B-i�a���kJ��}YW�/QHaMQ��&K�v�hP_}����t��wJ�e�+�/�%��`