`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17472)
`protect data_block
/sMJpJ7bNOJrAQMkvJHHAmDOicJxAIr3XSaAOu4AFENjmlLWyOgeSpeI79EdSGVQnGoPQROZ1QDC
yK95RIL39lc1WuUcFPvpGgNp5t8N5pZ2RXuap0F2qzX00XOQ4Uxhe8ffeLPjyn4W4IzA5ngTK8oi
O2DiPgZcqss+jItnjefvK3lusQ2OhZrcw/ZJowuldmBEH0/imirB8IJudf+xoiIZaLHNkmPyEr3z
gG3gF8Mjd1IUyESGSkec0OC49I428DeIymuL2CqquAkgrCUUhPrnKbRwdRU0yjDoiQRgphP49FUo
/hjmXnT18RJTOKzm6f2aJUkFPlTAxjGmBrdLBuHKKX9SV6jLxsSYQxyFGz9MCmbWovHimN6uEQ6a
swzZp3e88Rbc7TapXRqn1OckkNFuQeJcMQR8W8S/wUZvfBzjbZxrCWQGKBoWwKagP287CcIBLBLN
im2jbiO91llYxpbqD5L0s//B/ApIW/+yaL23qAiOSdWVkdkovntq1di9CnRhx2t0ZWdQLKHtSzfB
CX1mOsyTyGzDErq6ZWH9mV5R/O3N8VwPr1PqvdIXCLKxeNM7J1l2JdfWBfc44RSke3Tp1nl1n0AQ
Xb5K/+eolPg6BFKfBFFEo2QqPXUyRp3tr6eMl04S7HauH2cdHzJOofl0zGnTR02Az36SXZJMgRu8
VDEpui/NGeMiGQcdYnPUkYMb4yT/BGT8co9xcGc4iOKxat/TA+Wv5w9BXbm5yOxKA1ZEp7ecMrds
rOsTpE2MOv3dbpMikcDA0rS1o49DrIktceon1RiHNJ9MpT3bGgCjc1jyF854SFoNM7E5qlf+SwjW
DySUxFyOkTx2wVm50OKSzXilN1BuwgmdK7UJsL5yqb/FoulzwLaYbc/AO5IrOKPgURDxKHfAjML6
18cuMSY4TfcWOg8cEFQUq4BGTt4u1Jdsg8QSTT4R7TXB+j5ANvrWx5SFOlm22OIX2cBxRgL2Z0XV
4lMFbRdYdCdWtKGz2l89mXNkv2OWYNEbmxybSvL8+qHgD2Jxf1MokaPnYEmUTkKI7LuVqd/yuo3/
OqMZmLdEvns9ZcbR2c+PxRYb/N3UEdfiSanHJyYhNtQMF5couVIRIt3pL97A7VBgUvt9IvX2KFjQ
/TeJYjsvdZlp0ZvKg5Ra4D2yOyaMKFnBHf9n+4n1nnJLRQHD2jkdMNWMI3eYjWqSxWJbBYF0L9T9
TfgKptcBR82Yb2y1UJnFdjuRi/Xq7xJseXsY4Q3N6wkjWbWy+1GaDWweFn7o4EuVJL93FEMKdcG9
azGlDFObf0huCgv5gztaSQ5Wqo44Cu6UbNUVJizrBlM6geckh8sOoL9M/1fZMCM/xBi0H8AtECqm
d0yi6tdi8N9L0xvTl7ZoMCz1NTtUobWlLBPVZx8CLLiXPHRwSPLfeaj1wTMJgUm+lGMf4Z+OMxJZ
lm7i647HMn5ol3+8NA8zgb/PDjDmSmacAxSutYKajsKGvartDfhYBdn6pV/8E+tPaRPnbn4FcUIu
lQg+uOgQONB+SlQvbVRP+JTW1D2PUqhlY2qN5YLhxbYQmaGaCpxrvPYOd0OjNXAXVtabbuL4CuFS
Yj10nZPgLnMS1NRjTvXvG2KCnvTAHZaRYIG6d+drNsWeU/fcnNwoVbsfYAsLszC4r/pG02IlFq2/
L9wkKoA8KLkWngsm7KKYZxjCg+I5VMpcVZpfJmVDUSkrynY9097LJDzn3jmPS/rOEL8SyXTbAlaD
+XoYKTzqZTFeI0tyiGId0Ufmc0lBW1fp9+AiIVwkFelN2zBHb0mn+1G5RdZn35OMhmk6EQ+kV3A4
NFqirzmCwO4BGG5mh+g030sLIfS0mUT8NUTLDyZSE5KdhRFEAANC+HEC6LrcPNcMq9UxFwy/Q4mR
UqsjYm0gSsNRhhB60FIiN/5tfNqyjFVKNor3fN0QpQ1nbBxggd4Ba6kFjhyh+bYCqS15Sm66krM9
7A1C+M0A6mK1oalNU1P9X2IeefUiu/QgyAgXB+SmaGplPEY/ADk7ed/uTcv5S2d4FZRwsCV4YgFp
EJ4mDe92VP3r7kRmfuqKAiegdSLcAGIzk7CJ281lrThw/TptI/rpG2kb8aQfhc5FfNBL4242n5Ey
7E5KOjWbV9+ty706f/+eJlwaEHiuau/WA218MKxN/iyapTR6iW9fJNyO9/+IWQ/XNc3H1a8lw+vn
C9EpXBrFT9V9wG0oFMEvBRySNc/jz8U5+OlInjt4tTyX3qmZYFyWf1NZSTgmVhqoyBhzSfzE8/un
iYLPYCw5TGZN+s/GOFw+qLWw1zzVkmwKOaMwqVcUo9kchCMXuwRxe7rHyN/y5VdzehCdb+IbLcec
UyCSziVqU6lnfSOj351EWu+NFpq+vYZZe0jzT0CrsIZu45OeBZaGP6ViE1An0GGe6UWAmgSOsF/5
SSS/11EOhzYYeOo7f7tayFyIkehby2KNhTMpSrMJitfUlTT0S90g2MIrK2dTRahk9TKNaNcrfg/+
BCPDlQ+rzB83UeYPQ58/56v4pxb3GkgBQzLpHn+eSiFi3PCUkbsPqSySGkjG6Ae19OL2fdt9MlSV
mfkzldaSLECRG/Da32HTpYVCkiwb5o9QqFRwcx+OIYC1aDcOzBrp+fr7BfpL7x2Alqe320RKa8e4
CKLmYDKs4Hq5unUt6ap+C9kj4AHmLhO70/QWKiVQq39pYSHE/asNwnNplpBAbYKiY038Q3VxrCXU
yBKTGzefCJVrm4Jz9Z293YAvjar3bn/xHF1IFaJy2WifTYVyH89fZGIFTE6Ah0+ltP6QCaXYPOgI
8J18zLDovs2x+5nFxGaZ9pvAUMFx3tAbwaDArY9aTqm5IqOt5gMDDdIT0TlW0ti4CeZkDIEXTYnt
mo/xB+doXx8wDfeFmOsBRM42xnOcjo7U691brLQ10e5l2mdQNANlD5BD4pm1r6Ek347qskrY6h60
J11nwyz/nkUvskhZbUxEd265tqtTCiPx3dVd8JIZMetMmxhH8QmbmYxfJvteNqri4NPqbCJHf0T4
sUVzb2uBibPnwzSMF+SNWKAicyXHtfSibxnCYOntOVy7PEtdnFFqNNAYluDX7zLgFd29Pq7DKqYD
wZH3TXf7uiF7LLhtHohAZh9PZzrDfAIhLRYVHrhRXh/y/7DYKvs3ytS4AHKHRwe9MIHGHj1WWWA3
uKTYIh2dxMguTrVZ/vCoXiQ8PzaqwfHow3qVb42XM+2Ga/rBy/y+WYvPEFclm7kacaUhjFHEJlVc
REBYb9clEasyVQiZGz+V5EvTqXOdEE4P/URWr6ipL1J3ArhqhXWR1IvhcfHN6LIz+2nMEOooK3lx
42tG0HSiENZF47cSN0Xn8kVYP8XtIINVaaiyO3X1z3Gi4A1t8ClCF9AeVDyY1gYlB4goRo+p0Nc2
FIksOqbcGQgxZC8+4Fbe4ZP96GAX4tamoBwVHD3sWWRsGUyex0s/sJeC8rPvfRLJoSnaEeO4V98W
8AGl1smufElgz774q4vcTIFX1kz0SJqHEuXBnKPcNJlU8xH2OzQIqkGhkMatCXbQtJbDwV9cjk0p
E2XJOKwB/hwDrufFKEdoGT2QNtlHruYP34BtF52Cq4Alg1jHcDa/b0HkAt2W2pgWHDLJFPDfPkSj
swnvCwYT+ajZHvoTs2uZHFasbrWnJb0QmxIrJb/tL8AeKmfIfoj75TxJywyszNemJU4Kavsnjlg0
sxE5MpZmyJxdNqxZESHPsk846M3o7g0ngRay1KT3qZdx9LumWs9D2GMxNWvULNgkA/Uf0d/8s21e
OewPQeYAhv+xcMbZE2xjgwGz/2QZwaqeMhJ6pnqKHMZ/6daBTv6aKAhgez0PXbfdEc1r98I15DQp
ccEq3MkRVMDfZ8Ya8KXdeVuYmBLoKLu7irj2ca7QpPzkfML3P2d4LUBxrA/rev7gPEHoI1mlY2Ae
iw4a56jPisYpSxQ6RSI/Hv3q+LsW4wObAFepXDxSPMk91DV/KnPLRxr1lU52dyCsC8L+NPXdUBPR
F4Bbp0z7xb/Mke8Mg9o8DT1szTlUGZUc1c5JUQ0O3yqb1NM+62WgTYf9IQ8J5yy690ASBxMSJw69
q+W1nGq582cDqfmcKYeXe6kDCSkC6Z0HfdHeQWSQ/U2f/wMmxsXbS6Y9uZ6l4rRgcMssGEI7DUwm
PAnyYvBOHQraz2GvdkcC+WIADCd0LwMx/X2OiwYjDwXl9Ff0Em/NP9IgoFUF7L2eXOammgi1H/39
mbeB819UY/aC/fwB3SOyZWOmIKBZ0688RnjuGF00grI2H2l90e8QeSoy/Zt/I2IwcxqXmaTdc/XB
GLESQBCNGTnsNEnL+Psk7lPaiKLPQR8u4ejnPYfTv4Jt3bB6BEkOhNLYIFRi+WKj+pLSZRCt0+za
IcaeN4trwhzntMkG8JnLMwNSMv+TKb+sX5uRWRIhzGaGTHarHpKSh1ofc0DVh7i50AqaKnlu2HFZ
uJW2xVe6SANeAqh/3q7h1Gfu9afklbLLP6FuHcRcwint+OTIhDTD2xHQCWHnDGM5pPOKRczaxNho
jg/8DxmLft1PVDkq9IIVqXkGogXd+7qrIbHSo7tQfgPK8+NRt57ZDF8tt3S+XF6bYDj/URW2k2R7
pgS9kjloAYY3lMsl44xSFmLHlz8lv0yMgPlgOCsdRR0oliCUA/TslY0MWH5CEEiEuw1CvNMJMv4T
jlklx2M8GvcysUCUi5j8+e8WY/6CGom3MTVFjFBBzfBLVc0TMzrutrqf8cX7ma75U0qczfcW882E
8qU0ENlxAyJ3xn+kTKQZf+KjYOMXCzdjJZyOnV2le3CPu5TGYNqJTa+VJRswqceehIQt0KxsfUC9
gDT+eegItHZKC0M4ANLhdJedHchnXdAvxkR9VbViBXJfRhXcwi/EGv9jRE3tDkIGZ8J0aYzDAHKQ
FU7w9Bwra+Z/QH6Kd56OCJtL6sKCghr6VQ+AzsZR6ANNByS6UFO1Wa6pePBlMy3RevPsYU0Z5ZJd
txPI3BPKuVg8aw4RcXCo11PkR6PR/2UksRsHlXO/uGinuoXZNvWrsFLsmfpTynwbHsfsz8bkVmc4
eW+FKMng5pByUxozCBZPs3+/QojhQIv5RKeaeY6gEDsf2n3dBsSy0i1SktkOdX0DdSGzdS0Xz/Qw
4kkbzVd3BlCxnhPdo4ajiOBl0wIu1zJq4N53ekayXQjMp9JTofC8FdJPtaHtDocUpw+XDwlnf1X7
h5PGWa1Hp2BJulE8NUx4MI3jYjsavwSzDScPWfnQtazIbWN6eh85VlavaQkvMatExhtEvTMXD6kF
9OZ6rcsJiZG77y8/KahSGr10CCl5JwffuAX/TDbkI3jNbpDb32IKGngfULBlung/0NpZVydAQYpv
gBwlr/b19lsGQYOOp0Hp/49Rum8pMy7bRxOOk3bZyeZMKIphqmGQKAXKNXamVFz0HLJUt+Zn+p2w
1n9/Ldk00fXDKkgZjQQ1XV3nFm5TYrccJnjpnELpMic3QatSoyz4RvpD+Y2F221yQEy2JGCe1apB
Jp+rfCPxorEHRUu3jTjl5ZJhLP2AhpP6FeVNintHxL4XfuWZzkviEAv0ERijkZQ2WEo89/+fErWz
yF6iCoY7NCpQWzWAvrD9Z9S+J1leOc/lNNxw/9FHGD1K/ccfv49dXig59BaPYgpXt+D64+nJ097H
iQqjK6WQqyOd3sC4rc+45nFhiDc0+KR76JdqEpqB/6tm1kBPYrb+g6g1a7iVR965LvvWywBaSVkV
TeJFRpxJ11zMkyKWX1Yo8sL+OeGrA7y2cWC5U+W+7iQIo0AETlqnXiXilQPP8XM5d900dH86joee
+N4uVrokXkd5cXNnFLdpgU5KMOu5Q/ZBYiSsQKIbq8iLBuXhliRZVnK6q//XF6UHdR2h/hx7EBd+
d30P98XVMouSp4W2Q0YyykUCd/crK4NflppZTzKAdisxDA5uRPaWJR5ZwgoWAmp35MFSny9aE96e
3aQMyxWVykqxXzWMG4bpfWOyjbEd2KzW8o11zIZ4jfn2u2OKzDPA+JiFksQ4uPpLficTffODjUek
MZtJjgxqYd8ZG4Hxnd7doYNaTT8A4I9A6viuDTqoz2H7XSpxDKPJQHeqoI+zHsDvBsKnNVtIShil
FLEHf3p7ZPKFlwY93/jSbfwps2n6cWoBliO1D8Xr0EWMgLcSZGa5oOdQwcIN5MCqM1mCsVV0jYD9
WAE+GdzwF6S3co243C7A6InuiMu1GtYOHGLdicWqxxioeAnM927We4pls3HZMILzMGCOzNg+2hi7
a0W8xuMZ402f72l7cIb16NozJ64h9Juw6d64mPYyPDt28J/NrirPqn/ahKHrkBNDJt3+x34QfuRX
L18v78OeKlilwFnGTUfZCzMQv0XpgAfvlxxuSh951zKjziiwbXmY0TdD707HAJnMZRptP7T9QxLx
eQ3puGB3vHJ/ng2/1dGI4OEIkEcV2jsh7B/7lsixuUgHtT2FH8EZkJb6zOh+GGTWVse8qTLWW4AQ
pUQ2AmeGSiG2UlI0nxDk/ULDvuGFsE+D7fFGnCwR7B42Hvnd8tiOdWbrfH7UYLAooTjh2FmbgYVz
nivN+qyM2oSoM+lLEJhyNr9itZ4AtEJZS9l6liAEc/tf0K1bdJ8xafDCPrRRY2iKro26iD7w/fsw
8V7IFJpEeBxwiSvVCjYlcKMOHsV5WCP4cdz0GvmHcFwMe/7GdzFeIE22nobMgEQCiGNpWBDvm4sl
XF7qW7JiT2+TFz+HkDDgo8H4LwaVJoXP1Z0yWXUf/qiw2l84rmlSHV33R5pT0lV9zcIov2UC08LI
wH6K4JET3/kXRlA4138d2ESnN1HsG/G6fmzr5dKxcSpBBtjQJqFDUmQ6FfS4nI9DPqrpQ1WBTspB
Rc2XpCcRNGzlgNKFgY4SRb7kzfYuWU5Fl/OV5o8owL626bmkO5qJgZ3FdmnFZssgpryBrOOg/Vbq
d5FSk9x53Fuu1zbWJj6Fj/pQYYCGIM65SDDXDbww1hthp10dHYaRR74FRrUvQWV9LrG3OkwCXrrn
DHZ4+jEwwbXrScbqyeZJ9joRsvjFxhpttpr1PCuYiqhto44XD6QwWT+yNjctNK4ZcJrXTPoImCYe
CgLL5ZUbGN0sr/nGM3rriJ5JhXGjN0lvBoKlWBGfsmuU/1JPYH1LAOi3igQNFJzVUejEvQMyiOY/
Anph7JdrsOuC3hCAzRzSkpWH4JyZiinr0aUBT9aayGVXBrlMOcUS11GKFrZdVIdStznidonTDZ5p
Ia0waThUb11ISVixSLLsho78slT04ILCxBPxRyPWvNxrw/Fd2spoeVJoMCc/uKS9aAo2eaI6eWBL
o1ih/uELoVAOYObMV8GHOZRizlCUOAJdnx86VDgAbFss2wMrnC5hH+ZTZFjlVZ78dyFjW1E/nC1u
x62foqD0KsIOQulyE6j/+MZUs+lk7Wl57bbiGqC05jieEN7eyvLSiVR0bN6399/+pSWOpVFYTh0s
ar6yVekGvGL9qlI3RRha9Xl/qmqDbQlcIQ+naLSO202d6G0+SU1YfRvl7dImWfZCkYiBqp7BH9Dv
2jHHQOELdBjCfVU88JtyZVYniiS0y2kYB/XmjfCCyL8t2Ky9ULYuwWNzOqdD6vQ+u6rDsbJ2h+6j
OVuQFc12e0aa1wu8i1Bv8zyhLagip0b54lj4ieMpxL2bZPkpkPcA8SCGs/Po4dEpkov7pCKQDC5x
mWfGvWvamOKF38nCILGdIkgTsEzHXUzKU4mhV/Qblm79+jo1y8u3rLJ1oF9DNy0l7KvxxMTY0qJ4
E2dhamwe6tJ6Ochm84hEeZCklnnMz7a9TdTyTpR1MS4dUBOIJ6HQcGpmru09sLv0o2BLvtrolV5q
cqP+D9GWWcfPx74vQZzXwV7jgjxNUabmtjbpLY+hKH3q07nE5S6pSgo7SzksGiQ6+bm9w84CLCsU
0hwzfG/ocm9EVqCzVgm9jhZc+aLAv7L6mKnJb5lA+RddYU8yFqA2UmO9E9YSAlWkRxoEGDRC8694
2PKFm5FlS7VXOm2q4uHULh0OlJivVDd/ZPPedjse3j5Fs2EAZ7XWEqTaYn2bWvKB54GaDa7dghgj
C83rzESZCT96HPKth4ia3nQo/xxzOo1RWH6dYpmkik/9RxYqsSqtJXLwp+KOjnvwrbibyJ0Z589p
nDe0Xd+pUx2d9e3hqpLJ5qnPMgWxKYcbXnGjtj2ZrZlegV4o7VUrsqC7FDRPgHcV6VhK2nDaokPC
yMwH8iFYmPqGG9QaMV/fpVbJS1i8rjpyqJ1zd7Z1xorV/VhvO5q+fHzpHwbtpjUDZoUI8e3f6UvU
ReY9zmAxmocOVImQ7BYaqIgpDXwzeQCvCOao1UUxvlnNSj26b6DL8mkkir/00PSREVaVoQyfxBSr
aRrCutKnsQiqjZCDCe+qhonhcAmQ+vbs2AR4LInF3ekfHve9YoFKb1N2a0aou1uM6l9G1snyNQxb
yA6gjl3YPJIzyXtxuR6Afm4IEQyTSE70Egxslt/Cb0BQ5hZ6aczRenPTNfowYXcr/HBuWw6TkZkn
R3Pk31CJLWUswFDvCXc7T+++RGqPNutvca/b7WD2LEPw6+tkPy0IhxXY+Xb3C6wj41pZU5yvGfCA
12hkqILrXeL7Nuy8gJP9gkfQVBg//KCF6vRNgQKaQV1DSXrxzlPwLTuyW7kw4kjtdHEE8RC958l5
EmjWMzhvqel4qFbMk1QCoPulG9dHFeQ8swR8jXKzRIaPimsznGAVFzRsq78f9Wo1hrXWoz0tCT5H
MduuKA6S0iTbtJXKuBiVTmrLX2BUtDeH/XhJw/9w0Lj8c0tb4JaM4bNRvw6EUEAni/q8CxG0XcFj
2r6zypebjFkm5OIKz+1L/LmFWGLsImLj/0wPgbvnb7wpremJN+JsX9UjHCXiXr1Cg/yEFdazIHL8
iAkALbJ4pGmDkAoVKcXpTTpXFy6zUTYrn0q0A+ehk3TU297/GXQTA3DLZRlW03CVTfhGmBRmf83b
Cms487ivf8l1Vv+VF0csEbYUz6z4kBjYU1t8fCF9+/1tGeUeEZDVFiiFJdWP4ZQdhYWnSbuRcy37
V6KG8y4PkdmfC9bALaDoivbuTKCXBBnCHFByVcWKiTQifIVKyvdVmbPa6FBTEKFXb6hmku6q3zOP
Te0x1NrD4UmkTvkAni+8L1pFckuF5286jao/8NoOlzmF8fdEqucE0MzhVxUsVjdm0h5azJg63+id
YiUgqAM57Xp86oPv1xsOE+uLVpvtOUGAlBHm3A2BJ08KGFcUfe4zHiJKQcQyXE06+JJZrEQ4GIQ1
RzOqpdbLSJjLCyY56pcoLeeG+xKo8UAmjr3j1oltTtRJ+EJism2BY7peOMXaSfgJjZiTYBwIqDrx
mBGNBuYs7hmKKEqcDO6GDICLVlgbOwB/ysQSad4L/l9op8sytxEO/nRQ9d2VIgqRJEZ4SZfv+5ld
FzDxekOrMyVx+R+qJD+j4UTq5P1/Tq/9Nv6PwEhR7epKs3j/gw5DeD1wpZ4TGBzpAmLcArCHf8E8
a0yUNLvMbG/t2ORsfQ8f/qngQDRFam5vMMoYRDP2wXdi/UKBntma0B631dccAaKZvP+kijWCi+7r
K45GVqiQIiBl71wec07H54FQCbg/sHlYgWyuDW9/6p7kbNG/ZXBqYPMMF3CbHi4AQNX8kk0RCbgG
vyKwCk/PvSCXhJiCyYaDHP27GXJidfWn5TN0VA+F8f/hsQZ3cNEugsOCKKKz3KLeCOKM9YA5a2q/
suGRuKO43+vyh6e2b/QvTq+kV+Qz8CAOiXCupHI+hPklhn1qAQSdL7RraUutkRwFU146XPQbzk+9
533jciA9S2NsAfH1RJSV2t6wY2c6D2c9a8NW6Ou39gJnWEstCrj7AyiD/Ub3e429SY9fQck20WVf
IN+/NwghiF9f62CQ7+uogPOzBx+dwvuWON1iPGmaol7DiDFmoJfwKTMUMVvAV0aHR+rUIEvOKQj2
+hjQKdsibZ8u1VjBbvOlNvxQg2NCqsX/g5JIiXZGSCduno7R9Q5CkCADu//m31HipcwyzzwBenHc
+UWu0e7tAHETf8iUidcWrPJ+ZfS264vV1x8blTAiPt5IW+n5d6hV0IIhXuknpeBhFBTZH/bHzgQN
KaZ7MLXmG2Ws7w6MFx6JM/F1ZOElxBBVkBYJonQQ3UydpDMwbNJlSUU+cp2jqV4w5BfQaeKQGdg4
ObvNy8xjH8hxcw3l5jC9NvBbVT2WD9TjqTCWLIjw/EM3w5ZIPjGvt13e2vFZEMytY2DPfGNYumiV
0bZ/VuUeQBdAbmeZmtqk8bcRWl0+9uwiV2G8iTfEf7dk9MapoQW43CnqIgpvezZ3HzId9aSYpBHs
rRfadpkdalvGM/NCxZQYXx/3VxobYg4ZcqkXXU06vcaHUy2OyYLmanF92uFMWvvvQ4sNT6ywkhI1
dbc5y5+N2zM1kHrlfGY2Ml8eRn4iveQ287Hg9BXt3VFqmGbnobCx4fU9HCPUy3VLjdZ1YjORHAwk
gicY/HcxAujNbJAeGvWXmlN1wgw89ePRYertgmSPC0HLON8ghYFFeETeybZHlN6ZzCAXWiJgF0MN
Nj7iZogLLX+1PGtsz0YI7AugU7URpI3nFDiDwBuxn2LaWlzExzTE1cHDZa2kB+OasJf43+eka9lS
5btk7Norusw2krpUwHbwmd1KzKPsZV3zBg27XmC1enlSCn2Ab7KIRfP6ayA+Aac7reyn2jXEKg53
tus42TskVF2GZYoXOgEltpcyXBwOJTyvekQiz4NRnnk5XWuymH302OLU5dvQO/2FcpNhGNFmtJ3D
HOd1uWVZLGSO58Dgoju0yrgI5P7UfjUgZdL1vI7xmsD7bC97YkKtoRtT7QN7gLSPemv6wdpFG3D0
nVWO/aoEOSTd3ESQCb57Ab+iWOnOjVJKQbSrbxN+ES5G1UEuKt0Y/SEQy6aw4B0G6eRDUy3Udhu5
8g4waMBa3FlM24mwWIsTPvHIFQ8BT+Rz+wf+yPC+BlvZeeJLRTHBLnwD0bN7qcYCvHHFvWOiDzLJ
Gyh/G8BflP2r+abu8wdm+J4cbMaK76ytO4Ijys3L4cOLcZu6Imh3MUOJtxWyCpWQTtMV6ettUw+t
skVXYnbHuPx80qzcFTxVJ7khetk6/OIuK1rrFCDomio2K/iyBBJZ8vsSVBDQWE83KSGExgYXeGS8
pdhRwHwXe91Z49GpGjLnqbGf3O2vMRQMALZEyZR5kMynGlS5Wox8yNTwChqzimnZUnmbUg5Twelo
BFHLFLYtV5f3biDlREazi1c2btgdDYswHbGeZRH1cJHMZgpGOPo3/20UWzh9RMhjcAcFv8Ae921R
ot+iDEVK1mUNwak34d/4FO/yZip8e94T3IhCZkTaEfYoeDzSb6BgQKOdV2OujonPziWVEOKns8Dt
Tee1QjSoPnP7lBdc1DQBxFYyO2vGciQfliW/zyIIwr8MddlGUl5ZW16ThvgYp+32NJnNCqQoDPZK
YdPJQQHepGGns2UL81ZRbx91RhPcJDoNw6EJesb6Fi9Xu/8+4ygTsXZwCary/AHFvOpyzUh/dDn6
xLHv8/WWK3I8ugFWMxH6t2zYW+Ov9L8+06AID9rBPFHtzuoyF32le1+2DmtpbAMQe3+wzjymvZtv
9L7H0LHHyciHMwcVHx+Yjr9VIvTp8LE2G30+QS2YwLrMmEWMclDPWSqoCV8k4mPuU6TATZu3rRxc
hu1P6WpIXfA19LDv3uh7m/aY5PYTTUvs/uiiUnK6gjM7TXm4tT3jj+3lLxIOhjqJwJ4RO0cnzCT3
ux+uA6yJ7R85lRccRVeEyFnkhLW49SqrICDvDbO6q8flxDx0cPNXIXEIB21nGmiw/ZgzX60a6lBS
lmfFXlKoGgSR0ltwQBxvIUBK5BZMsWErLGjULIxEWtzB1c7yDCQRUYYY27HS8x01ehWSkzLOkgg0
Q7qnii6MIC5QZu8+cXeYWgQCmmxCvQfcrsbunizKDtngRQtrBWq4RTmJ/oYeMZc1viWcsSwWRlZQ
JgJRmoQCXW4kPFcPoBS7pPT1j6gpYPpOsCdRBfwNf8WKZOtIm6bybWtTt6omLeQSbXWcW3t9EF2H
v2Hbh8DQuJdTAunHRqa/Zj8jqUtIvJE9CpQ2WxpfxTBX6z7FL7j2CtlpyoC82rNROAspp95ZyTkf
C3PIqo+CC3VUDZNagQdtZGtCVC77iDqWzocb4NnqlsEovkHjZ0I+ab+dcJ1o765tYJyBNIr7SiA/
5KxjqXbgG50i5aRQ+OK5qtqeZOWHEkdCQDLC6VtONC+z4BRmeAtdfktrlvLd1B/rJ29cbjd+qQUG
StREhyu7YbQl+BjRQAjX0Xw4yM7nukFZO1LCwYuO5C9ng/jauspPviWUzSHejiv1YzzeUUVcjFJa
4rW/tnGQ4Qc8qfa0kjtw+uYmOlB4B34XZBAo2A93qdAaYuC3fWP4LC3XmGCZAvCd0kzam6eWLwRp
Q5OpRuV43HubdM2fUMcRniLqT9ULAcAmsNfvQzKISRx4Oq2ARovGQ1MqGbGIHIVVihHFAzdZWcUy
MNcOb0OpPCl13FKE2YveoLuZ/lgVTFJHA4pc+H2VLHzHyg0mHMZNps/BeOZEU9ARHichqksL72VN
HL2QEyjCLZavtKgR8vkVcf42kABElbCrLjDh0YnVAJ49VggHzeLZkx1EAQt0VLrkJ7oo8/LM1aw5
/R/D1OCOGVx2/UwqtLYPlsgimKVqg6sd6O3Awm7zrPP+hQr7vke0HEFRlzODa2UHiJCDoTh/S2c2
KAplM+PxXqyd3z7v0QoR28sBYlwSoT0LHrHnGiHWyd4Wx/ez3aUhqN2BR1Ue1ZLgnivdD34wLkH3
LGPtqROPXL3goiKJDkVvh1l/VwoOCgAz/BbHwBLxiUh0Q+1rR5rQzpe00fziqg2qhYItRwsR5Wwf
TILsG+roOhdEAWJjljYmqhGVH9yLvoP1A28KOMmpr6kwgKX+wy0YEs3W3ZEUPJxY4M9vJ5Iw5zja
qvQOt/ne9NZ3OzNvr8eM1mkJMbRg4TaoJ3hVvbh8YW2Ki54nmKAE8wsIo6tHGV/xEDhKsoa1gyZ9
+YWGsq/xzJPRTeE96ehSVxlO/x5kM2q1L6UqfHPANb/fO7btnHPMi0Z1Qe85SUukwVmd9MrIe/NU
i1d0Edtkte+EXW4zdGOB7g7pcrvBBi6L28L9pDDTGyJV8lH7XjfycHwKkak8ws96kwor8QFVciEd
cASO+RYY1j2qRkF6lQva1ssliiQdxSDBlvE/rA5HCT9oK1eDaDoCmFQDfLGe6RK+jg0K4zklr+hG
Fknlg217WRc8JeXk1tgawavTeVahaRBc0J9MS36WNHLevPFUlsdNxBpxUlZazE8XEZkUgoXvylgP
xGuhGRJql1x3MQT/iefRCyPLOYzn5nukOucoJHEdFqgfk8/nug71CwL3o8CLgdwfExQF1+HCjdgm
a9XOwpYq7zb+kA8fN+Khm7PSgzXeHMOgTriTvs5VDmzKVKjiAc/sicrynLByZZMrKI/KX1FBjhrZ
EuZ/o+cxx3W8t9296o8w2vLhDDcOZqLhXTVkRp0fDd87en7bzQw2ubIzMAtE0UwwLvO5yMow2r07
HuZTfKz8y0NaGlLksfY5IVx0sigHigL6UkTuBA9o1sAN4XX2pdY9nRbbKON1G4jVFice2ViaHnEk
qhvF4bmXL3WezC2HrB/U71C3kwcMzAYAFvyt3UWbprsRd+Ce6hNzqmCo3dEc4W6RteNL6ELs6KeO
pd9vZ23NAkDoVDm4b1+0AHSguNgFyMvjb2kZyDkpVzeKI8R+lI+T2yx4Pp1Pn9q7PRiAyRLQHzDG
7iE1MOohdXMiF9jFXetEPO69pNvd91YAlt605Jj+/dblDs+XIHgCh4OPPZNs0thKZO1/w3+aapzW
g+XjAliiHpQGOA+gSo7A/iT9zqPO0zEU7NtHVIADbXxD8bPGIJPR3zBXdULOmc5JO0ZC0dJ1ZjLF
r0761BCFwiOY5yGFUop7p4ATSJT8hqZ+dBSpy8jX4+OVVC3D1KErzxCa1NPYM5SRQPrElFPq7qe0
us7A24WlpTA3HisJ0K+ObxPgagred5ET2Bu1QXoAfD6QH/sDlNXfguDlY7phsvcC00Mv7eeC6A7W
qKXXlEB9RrJlJ6QrEUIr35Dd7GfnuPhfjHVZ2+Ji14EVTxXOtK0TzqdnxmhOl1RUe2jaAO0moMPu
ongdTfl2VGIRVxvLXs19tqlHLMqbmUUSPY1ov8QKr3t+QSs/FiqslEy9IV/671ABuKUPZYH9xcUy
AtpG33zVVTI8g44CGYF8djhtiAsrKi6Gaft+DxkniGuCFRF9verOPDK3gx7Df2rBGePL+R0T03S9
/QK9FqJlZG2JnJymYMnPhN9BIazK4ZPY+xjTupakKL1I+5oOVgpHArV2DLyOhm5go+Fx+T7JQIyf
V2zD+l+/tsv+CIeUlyayY+wY8irG0vh/Vzs9lQXk+ITR5deXTX6Sp2L+M2yLVkK2U+AB5ubA/KL9
PwnAemmSKy7UmXUQchhbJY6hiiyiE9wfI2fK0ij+pwpDub1z74dzGNw1TcADGuThTGkk0RJONPk5
C+K5CbkMN7N4srD1MvH9He5d8BqQdyA2g8Pa5n4cNHShVQBKTXg06bxvvUPgHGGeTWU3ax4FBTRc
KXzAyZDi5KaGHuUtb1IuAVIzEuKuROPmsrcaGYvUWq3dkr3z8T30YlfPA9q8ql6WHM8Dv0qiqqoB
Pamt38q/Wxd/BQUAYE04wWtCqzj/DKypeh9+jx/8yd2ibUvWch461JvRwc0W1XnZch9IJb3EiCkm
l/73wzZ0zgHkP6mF7ODbSDFL9fjG8r+CYfMeH0Ssl91MXRT3J6Ouc9muhwn434IDcxx7ghXyCgwr
zRbBY3gk3IPx5INWCw5j0LtiiQ6qSRX24WuTxP1cCmuUcxJfeRo8oLZK1Lx9916Co7pepB42HjEh
VhN9pqxAB5bQJ/1s6PYS1SKkanbay0ltYmGGXwhqdwTASGjrJ4XFPgfkHMVBkFkeFuj/r7sRuBws
h5p+eHN1US8XSGvUmuI8xz1YQ6JTbXd09J9+bADiIFFLW5rXLZjCry/3pzAiXYyGSMHvVsmWpR1f
5cHeNuhPP6wpDXPXidDpHBh1bvRvIc7QgSDrpQsyRJTpS4456j7B2BZ6m0StXenz/P16KMxlmtHp
7AYdRR9JNIN1J8uJbE8mMW6pJRFmG5mNK5bTh+ZzD/KAjpmOX7F/WR6J/ASuSzwhVbq2tcSCYus5
XmbmChcoqWmnsjNBxQzDD4kqBqIdRMMQLDFPYctTfgGSSUU7rAkKKof50/cXGUHMM4F1quojj6MG
xZ7sABi7Fvm2KmDg+QdDA5mZ3IpeDI4N8V6pRjPTPJ4VHhHx3jvpIYRqIamyMUtCBdxrMUrv9XSi
XpQshK+Au8OJcL3zijVGo1ycSBPFquJP2kZ409BYkjLTqCJtktU+BMVYIDdXSysqaBjMG/RpUnIs
a7qr11OcAFcavxOkOMiK8o2esI0qpPWlx5l2kxpW588g/4bYsEasZsoip+IxAMJzBT7KJ3aS/aUA
qZFo72KtQP1/zBP8W8m4/hvqG/6TTN7AlvthaVAZhGJNNi+K/KbBStb7bHoDB++nnPhGvYNHwWVD
8BH1OSPfti/aWJtQ4i3Pj9LkONe+uIL5eJxsJRD5ieijd6NpySxN98XxBZ06E3/Rd7F9YcJtSwTW
lw4/ZZFKokiUvx57m8S1pRQXNCPHlWKITFZKpE4hJW/F2Q8Y4xRQQGkg8kmuHXSknEtVIj9q6gw6
kfiC7FTS/cUlATO5jjQq0xYE+vkIAhKTGakHIMfuVLhGXuk6dnc+V3HbPMvaYykHC+7TACcjwkJF
amjiQGfC7C9wfPecfSghMcihFM/TNe2SEwxYpuvuQDd9MVANXi7mZlehTHtvDjPTyJ85GNyzPAVS
wb6Q9gOTXzN+kICLpQbxiQwByPelrXKyhcbVVf2vf/XjKpte3mpxtat3idklF+2J3wGFzMRsheUf
kZ+OZCDbt8ZU9DIz5RT8aUSUzpbhNAkDf5ijUNHXVwB36+YK+ymp75Wf4Hrpo1hgTsgqSD6Qx6jX
U3CcB4rMlkAJ4XVsG3QJ53De6W8UeZqDEX8cHd6+6jjU3OKMmtOnbfFXJCRxLJqfMjmg/hhnhyG/
YXZhDlNb+s8RhbRUZt7MOuUfXuxZgqzVqdJsx789lzaJRluSKB2R/rK1x9gzugp6eiCHVt1EMDha
4B9CaELgdYur21Ik0uQo9DhnOps5guh1wWTzW/UWhmNun76n1IcnLutnAEUHC69YqnL+ergyuRwy
RDluxxURQvyyjIig7vaanc0nMC86c4yljIpULDWFrJBCHwfH5bTYFd+ixI9PDUB9UfkubiFf2zrj
slL5uiw5pXVOyZEdqmE8U5LdJtk5O2Qn32Yc0vmJZ+jvy6ChtUaPk9uE8w+hLZgWyuQTNfBxddOT
1MGcm0vT0gpxgklFjUBCT2Lz6ysGE4trc1sXT4fMljuJRW1tiyv+UyAA2lqKrgzX1UZYHPsf+G3+
SLVOTuiQ3HghH8aafwZG7zHQiXkqDGxMLHTXAREx6JbhW6kTOBO08kgG1mL9RnErhAucWzGWCg0j
6MVhRZLJY005W2I4BtzsPnp7Rg40To+KK83RVKMTz72c2vVbqkQFpkZ+ZOnh8EM5uTlX6j7qjbC2
5NFP8MUIEyVqvrIt5g7MlMVeNmXhbCEOcQelJJi/pOdGdl15Q6oVnJuXz61O2jfVc0BV9Yx5NHID
r0BNhFjwOS6t7xJBniYwPpfAku/0vfKFHnjZxPC/S/KHCOFcNh+glYq0d/i5fMvFjLUaO5A+Zw7Y
sdRSGt4vGAH3BlRemWkjHJVpglu8R05HzT4VYEXERm5OObJrhLrYk7QHy1yy/An4OfCZ8wbQBYMW
HdNPjQtfCBbuu1f83nY1L3BkeVePN7ToSGRiiTUdGjQgl8Zb9PICnxdm43pBw10Yg8RmbaLkOL0z
rhngIluJy4usd+thGpBfJ2xv9XTI7b0LtUVZcTK72+cOKbFH6zHeTFMr+LMeA+NIk4bPimSamuOM
Uwiv93baWVBN42NIe+bIifptLcrObbMwumwLh24MnoocX9I10A9qjYbLByl2nJUuog0iKPh7ZaQx
0Lgr8XDdnGnPNlGN7/Q8UW20GZ8/JJK3lvJ+RGItAGUAOY0cINPxu2O39sSXCa9IiMo8eiSD91Vh
1OaVdEDlolhG2bK36KHqiRMLxFGDc0+jmGGDD/uo8KAvtSq3qQhpaBe7WTgt1EQ/JVAW9FDX+MO7
KBj8kYHc5MbWjHRIfGWZSb79BhvU3JjxPMXguFiRXvSknLHiM0DYblPO+Nw2YUaQg7OeUrz6sAht
PYTK0TXazNqsgvqH4e8TDBQ+rA3/MLF6LQOd2I0m2UYUyKjGjFeEKsozA3RlrDMrf61vOb7bjCQV
DZhJGSCmQa+WMXzaJgyAfElyJdRU6FyGbc26tv6WqTxWgUqLK9zlHCyws4Qx7BmQMW0qIOfOpYY1
na/0tJ1u6es0eSb51DT+y7qdWckiD836Mm3nEzcanhvifsoEj4wjjtt2ucuOhnguhTekdDZ05ri6
N4TwtVHDlNAat+BA7FDvXmrAug1LOOO+v85N7MevX1pOeOeYjLccKjvFi39PT2G5ellsy5qEpECN
j2mMa+1f+4PNNHqDkho2gTnhuWUBTw1Ye8FbcUqnkJw9ndosbRAO+gKIohvW8V/OxrhiCBgdfeE3
2GSZ9lwc7WFT9x6Ekd8KywhPe6igeutxsGGsHXUYWCDmafVffbQ6OajrlV7UV6qESKmEdjvEAwtL
f24/iW/o3Wt0IHf0zZ3S03i6EeRhq9ankTEC4pPYYsuBT20YKbwlaogZNGF2nLSU2ex0Hrs3iDrH
0esYIzp5wovSZ2dNqp+8yAUI3p9cRj74oyn+DxsqkJkjSas6jMsfDAnDXss6lBoUEnZnmjk4J+FX
nmo7yGXcw6rNLpNnRfbWdqarJn+xA7LwsCgd8U2PeKa/XVO5GGRfKwsMKl5D0Zb7SNOOPHhNhHgq
lE4urQ9Fw4/cTwShdU91JO9Wdfzjt9cLZngqe+UAg+tt3KsFYkCVE2QSITTpWgFPmdscAVtG6q4R
bP2QO4Ftv4AMpuukYz6tQTqlzfsj+1rpL50sxzU7f0Ydxxq9J+BYcK8ggdZxYShn9Jv8eiXE1rmu
05I3sPUo1ukyW79ZjX4df2LBj/9hehnBHFjyTAwvqwUg3t/mZiR0RhJ3QvBC/o5F8ARgLVpdcnxi
Qx3vBqgB/PPaRSbi/1LtFJ8mowDwQtl5sigNDg+50KyaYyXKGzczGXHEY3aondFrbWXym9cyeZ/p
oQgvHKXXHhQEpYPkpk/I5cfzO5VSp6VO8/EW+eDsy6Zcg6h2KK3kH+KiuCVKwIO0XQYtaOH0QTOP
u55q599uinEFdyG9hOhUrKApMn/Zet1xWPu6Wmoqw4ZTMbFKb7KdQz8m3zToLPNRfd+SAHz8D1YN
2G2LP2yVCllW5np9m6aQ4RMBSf21/8KPk+n5kUYTuoDHsTPWFv3ssnOHRYJEdShwDF7P55e21Z09
kKoG771qCUvT9m+s2TP7LrEPunbyslAgwJUGaISjhy1C0DQvCB3UD03fWBuHRtum/oBhUdfaRtR3
MmfiW7HRvKUaO1Uz9htUTkwCAePVAAkjLVL9RdH6RaW7FDjpMHi6poRM71yhbLKkHm3QLn2Klbmc
UbtBkuE7rdYT/i2iPVunZ5uPkaXljM8LYqqBGEGG5FBEoAi/0PEZQ86J0O5FgiWYUVSDSpZ6mIKZ
UynyuES5x8lMnC2YAXbw6LeTlpZvzVqkv9sjwrx9VZgWVAI5UeA9mrFbAkRsvF5hlHd53ZxQ4H7C
c7jqEr6CWmoOHPflmC8PUkCoGNa+B5ZwuDkzk3EnsrPPi3rymKjzzSDSBFPKdnpvGEHydDYYxXqZ
UL9N5CpoShpSQ54x+MqMtaR6tGqN/4siKax9U0y7bOPUP+8Le7wxAx+3wX6YJHFEJ7wjQiELA3bH
BEWtmTM3406ZmDgOstXjwL1nuEDM6IUGpdGGAbLHzJHNiVKbPX2dy7HYd597u4gq/RFlEZGp1wIC
BlHf86SzWj1DPvwj5WtHWQERCisOHWMDvsABIHnOFLJasWOyWjIwZW34uja+RIq+wJGpb/DMSLjj
T6fbENMdRIFt9u3lXI/g8VD4b1NBRHt2lSwrJcTlr2BfjTujJuaeqDdgpTTvIjjr97ha0gLp2iv+
hDH12/wpT57BnV10Wrsa6wtc9DhjjdG56TDD8EsfDAkyaO8kEsxoNqeGmGUCVZD0VOdmBUiDNXJf
Oe0IzBjWXP5yn/bKLfJJ7McwNSepQmFmOMuKR7v55O6iHf7+HqFLqQasswF5pfJUTIR7gqMN8I0S
qLJkj89PF3Z4ONIFONIR5OECLT+JYc2HHD+Xip8ePh/OTSZBiItmWEqWdWRHPucIpfyh/8Nmh722
CWiVUMLBQWdwyZD2zr09tyRiR2+jXJ5+t5FRJg4TZ6C1ptduGm6nnzlNl7btYrI7JVSk89rI7IO/
1KPWphIKXIMAnUntsZBi/Hq4/WU1SLmHW2hrK4ia76nkekvGwOPjYum5Nuf9dQJKmNl4UzbBAbw1
rtwgGNomC9Ye9OaQaSqMT098fkPjjkkAEgtUiEWX50BHkAZvkYAKvkqLS3twpP9S581JgwvVvZuO
+3HzBb89fgucseEDQcnu+0cpxMMAk1qSSGqoxXAxyzP0+oVj7wg5DPhBzALbh/6rYJVI5kgdRpvO
0eTjpJN9C/7jYFh3XbG3BO1Xbq2BDnhhBF3t2VUBoSjOt1EPx4VcFlzn8WYA+mnS2wupvaLtxiBy
W3moAjgOnWsGaphVEUNiIZu6Ie8bK8rQflml39F0qVNJiIpxeBessYyDMx1NTt52BvM/z8n+KUCA
Wwv6onheL3+XlaBl0HBRMx5nkYq7OU/+9NkvIKgZfRSw8QwHPfkP7X0vpjvEXjxHcO6RvDNBKsbY
t2nbXv3Qzjjeku00AHYuAkP0kxtu8Vu3iUTRYSyiIaQkDDU8cBtqT7p2yf2Mv/jRrXNbDeIIeOnc
RA2dxErUJFzMtOkl52yZusaRhuXCEzJ5Nthr47xi9Z6T9f5DHDx3ZmKun/hVslTMXyLn3JpGILxg
Gtmg9ly3F5MgDM2HrM0YHMM5GhpD9U8uW/xc7Dlora/fxzkpCvUrXNPj7C/kMxMxdPDzjJxXN4x8
/ILEB/Z4ISvjmQOv8jH/RLC56hyzo2HPduxbXiHaBypWfbN/od/TCXGmuDjR1ZmLm7FAApCEP+v8
980vSsUIok8rO6w6xln8c++ejL3RYRmtkDjJdzv0bU57twJn6fyjsOXj9g5GFR59APIewUrRbhH0
+75Vqz1eB49n4g72uPJK0AWs29alX5VNtgQZCJdfIDuPIq8F2Nlod+ZGnKpA9kaRLlflbqqthWS4
1kMv4Vpks3SCrvLIaSy5lR0pdOUlBmjxRVqscMKoAz9/+ExY2keZG4ZI0j60uaxVGw/F1wUQOqcC
Hx99eKa82edv6tN0aGB64BRG0CniJzBiBLTLS5fh6pDDIg+79tYSOqau/plAQf6jwJfuoy1zdPgj
d419BMLVCOT3mHLyf2/pIjjy6TRjfnYhOqduN5C/K0Obp0LyVIRwRxImdynZKSF6//AlXDVe2TMP
TBXulUlDqLIXpLdT+vkI0FUuQBaydvM/Fh94qj/N5tRHFv5RHStLuuulYrQSDgimtCN1C8Vjo6pM
dvvpiJBR7eC5ZB0lyTK7UY6AJPp6Xi/CxeN/BUl6orW4rKv5pDrZG8afiPeWWBRFjmqwSg1hhFk5
hkukQXLjkxdyFoDwkYDAesuFQC94EjZSPAzvDJ4BvFZ5jN+Nl4p6LBGLJfr3vimfmTjkdA3Pidwb
5hKXp+QkSDiKwIzYS4Uc46CMc+UOzHIEwY0M6YMYM8fQg/SGmBSl2OcjA0ikI1uzBQEgZ5jz0PqA
MBXaZm1bhIbb4t9fmq/1opqTJDbDQo7xmOkFDNx1RnmpaK69nFRP/rn+u15dooSjnexi6OwFIceH
62L9t/0GaOmgrBOrh4JRUjd3tIgJ7eth7iUQnmY582ZSJTeQ2shF79IrXbtwFUKV3VpCxzLqi7a+
m7KLNKNutsYx3Zl8x0zPgAWh8esHBz8K3OKWR8KmsBXji+DQ/8bKQoqlvWWU5lHBu8ciYWJfmi4h
ebVCIMzu5wMTDzQv+zpcDPsOEYngoc+uB4XBHpXwJQaijTPbKeG1sATSaZ9VGndu2SpVLQUKSU0q
waIHqPlqdcQ/wy096UdW1fxTqccqCKPVOYREvmvW//qXIfM1PTu7nZwL7uauIIl1H043kGslOKM3
qt4wIxaVQ8oCmnLtJH9whhe8N1t0xzvT057orLzdeYVIAgEkeR92p/mvpgjXOQWnYluCPsZ/pqiV
bF6rSTjnz7KL09Lyv3cM6OPycTdhhbCnxnFH+bITyIGPgPlcX3GD6im1i30U69hU/d9bhBlE5Tkt
lqAOzs/g2FDxgrYNOWCUxbSb/8F0xxU9KB7+g6y9eXdZM1TnVD8LMTHFpu7qJRNPp2AIBtJusyD1
OmKtlhFjYrXQBfy5OnCQoXjyflfXO0U9+AmYvdFDS/cB3FHqs9R/hS8WjdvgmPq2WrCmo6cNRKfI
TTGK7RKOPgSDlWTir5XXoWEdL1HaghxAJ3DE5PZTVOKJD15surARiCxmpERhkPJ6wVu6JqCTje6W
dIIpKA7RhD02M3tvm6oegsmZiD9aOmtTcu66TyjXp/TIeGRgvgvb3ETKDquO3nLLRS7g21nvpHFQ
W5aGmsJiFxOGgqPzi+nCECLaXjJqcT1ZR+a1ctkwWVQaCeAKHHHcuseriLzzeRSVm95AziUWuWyk
M3QqnkiETmOJ6MjKIemjC/KxXljQ7e6vnQWGSUOOKZiq477MRnBEwuC9fbDrlpz9TpJZMBnfFQ4O
Nq7cdB2JvoD+dc61KyDrd/70p42Ao0/hiLJyA3BSXcr83Tj/9VW7Wfa46puMo9wb6hMDXn+yNb84
ItiO0bLW3qQYE7Zh7UeQg6uigCthoTKURvz/63y4WJceDTEmKwQddh+YwCMtDbvDpqqnNXUNYGuf
RyKomWCPB/6pFZj4tLJDjGImiScS4RCZzdsHnv8XSSw1S1T0+RKgEFsBBZRbgC5wVaYVCCKaGi97
XWNpdIF5z2yMgpCu5k/lQyr8kXRzI7HwtkE9V0nvBGiuPN0AqdG4yHnmX0dDxuSZl/I5geQ4MVdx
8jYeUumRZFwLJHoljHi1jiI3BGr0ca0TsfErEAS3raeapH93wnVg7/q2d2Pa/5eAuQ8R/GKK3d8l
CPh16g9Wx8ToVJ4OOK2/5oZBY/xGqxVjMBx057//+PFyYAUyLgh1K/pLpeUeE44Uiox/20sVcSnR
lEHTxr7BWhn+CLQN9Ch1d0+Rpxh4sJw3kLpH5jUV1CVnsSLXus0StRh2+9r30JAC8Ivn8bvYiNjK
NwLMNMZpc74uLbjwh5qO13ZZGhExG1triKDUkw8GNnLS0k7RxEA3bczRXjE9FxqYhfd43SGbfdYQ
5qCF4Ph3fQ5uBqor+VHoULUabNuoI3a6lWitg/nFHh1tpzM6FFx9QBLC/+DQEfkhEOuJd9sX2//C
TXP9RkPk3JRrkBBohYlw7cRRrhQTyEHcR29y/48NLKoHshJ0LI74kPDRJim6bmrhhEyq+f6tqP0F
MCkfs28aMPllRWxIbrKkOTd74zYv96fNO74c+fBY3ELWyaPLY5iUeotWY0Zwe2iTnUhQZ1i9YOCa
bsFighHUe0pSZHj8HlInXXjDyu3+1+NJx13cFyTzFYUAtnzbnTk8s1PSctsAurDedydn6psH04qM
1Lsq/SLvB+ZzqEpV6RebRLnDQ7lvXM/dW5vjoBsr9tbXFxcog14AMJU3VzaTdFvrNfLmV0N8P6np
hJYhlZAZxw1JvHxWfaUe6q9BAbFPsfif0GaG0WXmNbS+d5++EusMRZJ1MoGE11TOVfSwpZCNysvd
xDrIMTZd/5DnA9iZLeHuCuxgV9uxmpoeg+O581E/4J2ZaXjWsKH7pD6rBVBaBp7EGUAhk8d12ZgJ
m4Lx2lkNJHQr5GMO4+NQ5sWcI3xwPukI+PBzvl/f
`protect end_protected
