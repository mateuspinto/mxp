`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
d/7RgL9MUydeTiNfD//J0bV6NYxelJlrxDSWdk0jpqyXmNoF96W9e2di5TaIE2rHZniiml20b4xb
Fd3p+8AMdpD0Wt7hTl4Csnf2CeAHR6QmADgQqnS+AFFvqJtoI9mKtBOptMCnafT9Yo1/R6EPu+0i
U++RaKQFogYEjkBsBIiPCx7fPr58HLtt+GUeaQh6bgV4u+KFBZHOi5NeFhXZAzDxLttaU3aPlHvo
8M7E6AlGKdyONO12Hp7R/Tnmt8HMdIJ41bmmA4CbeEWIirWNFOpZ2xXUmSHrlHmbVYaEFXDlqFGS
4LKGChwEIkR/fF4zWI2cx9x9b/n1S1kyq87j50NtjyDOid7vYKTQLcK+4XD3UdBjpjjfvkgAnOpl
WocUN6QKPiBfN0wfIvk7kagRnXLlJj990rLFCCRCSuYSc18QT/6yJCq3o9XRG2HC9gbsU+yhOg6L
qQnMuC4S1UdkAlqQOr0S5mtWTTwyzNYYbYHVfu1tnD5jdSJYlEQdCDgYYYODOxLhknvXI/W3PK4I
xMxVTQb7C/ruTFHrxPle2039a55oyivVD5vJG81E5TesCzSRohE6Jpo/vpwILmpvnJfatjl5d7Iz
Ti705Lgn7TcXApoSKoahGeoQN8hd+ZXEDfbBc3nZ1BHQ5gPCvp2PeoM234Eyj8Gho1nN+v99Gnyf
GxRhrqk4U/XnBmZP5nChOyEozq+NDjzjemec/hGF/WXNxqxs6LfTE6AHmxIBIi5JWB5j830Zqlpp
Sy+JTjB+VLodZEVrlHRLs8/kFsehgFgis+gyjz6QRo7mFEP9rZ2Cba9w5uWZ91aR2RbmyZ8ngTtV
JyROyyxqbu6HVdijXJXSlUkT7aJntuDFvHQP8jFIFj8BIUiSxuwe8jaJF0hyb02uPK+As7iFB4Ji
myI9ogXhw5Z6TsezdQV/YaK7UNTQ2hyumgymigXsOkSXDVRvBZpeR+x+g7V37O1PMTtg9pFxx8BX
GXE2TXiQCiRmfqDW7jbXRd+8thvoY4zTtTGibJrkndAC9EsAwZemxm4kvM4zy6vMosP9+VnD78DP
PLiwBHugSd74X+Y/NIh0FO2G6iYAH1PbPeyeUkXZAU8jVOGrJ6w/HGEinfG9bw8/tI9XaqNO8Ls8
VC0Zv6Zd2ltSiiW8eUqlhahSVC1Fej5+uebZtu1tqG2DTUIKo2UCaBWk+M39Z2ApluJrTFrV/B19
oNpZPAHqzdhpPngTyyCFFs15ikGWKz9u76MebYtmCJhvNlO4HBE5lJ3UgoyCBOnIrFaqYoiSXAsT
A0FhWN6ZGwtEZA2cuJCBeM+aS8EsetTW4kPC0mf5dZFNXZQqryndQqoP7VrFPLAYeNeJwRqg1Ua9
SdIpkUNyCm5k/w3ykkkg8rcSC+OURybI0JmKHxdxH9fucj/Tmu65ocSHKNaZD7f1BYZ1PnhZpT0Y
xnm2WMmX7+quhCA6YzgMb7tjX0OEwQDk6zcdiUwF/+7diUq2Zd0urzaYNjD8RbBjSCez7Nu7VZq7
NpKXiSWuRKsxD9EJap1ubgk2O446lgbOyLmdWzLFbsIfBEA77gIjAx+CP5ruChsbqjca5QXv7eHa
yKY7D4ASzHo5OqAyK8Xi+uJFraA45LZMau7OV1BbLmEuW9FVrqHMS0dtOcqQTmFzdUQNEmQi1Zp/
ITGD+Op2OQNspWTGmPCSStDfEKXbAhUaWjReTEMYQCHoS+VKkomwuMNcwOGX4SX5vDmpcDBPXCpM
v5hdNJtv+crOs+iPDZWFypzTWk2LcBHYrOtOXYBKlR1k2xy+0BnHMnRaiKSlYMnHr3pj1c1d6eV4
d4ZfK6Oi/tV5elrVGVDee3PkYfhZRp8DXo9LJTK+kydvsoKsS8RmN3AcUxFR+M17qK2Dk00tliK+
1N3+Z/g3WlxwBwHEvZXQnPTQX5n7SbtsIrxJQk/+TdHlvmm7qUGAIfYiNGsQORIml/Xu6Y3IHHps
DvJ5Kx4bGg1wnvwoLAlnSJRqgj5ARnDvmDWBc/u0Xdo+Kea3zW3tA54k2AG0iiaH9SJBeSxYSsLe
pkQ2yYi4Wm2JhxQo1MEZqEVsGh0a0ZNk217jn6jJG2D1HVBAZIUiQrLODfdnaJYvFPrHzpwc8lmK
xDEEwwH9nSxanboQJNnLY6k6Hmz6h74tTLIEiVvzUnMDFE3EI+0U5A4vAp2npxbH+JDF7um7NdBO
ZPbd7PyGBJabWMfHt+EB0jUDsBJSMyaCcn/83UxRIb7dRuG6B/o1HNtFULR8YtVJXyyRw6ldYG89
9vXFC1P1uoCHzARolxwJZpaKMaehnUEmzM5KiqHXPaDc3MN0GvKxoRsLCHsKOpQziygLAEjv3ak+
vqt6MUmF0iRmV1MjBVkPBcBkuVyjVAPAAZo7iMRyNaJlCApOI3u1QAbQCYf4HR2AD7tBebpCfr/R
H9eAA/w1vUMBW3cOwvyQzS1GNG632rtFF2FvTHoi5n7lQsDZc5mRsU1qPMiM6qTvx06yV+dAqAze
moP8T+hI/89+NBaBbGnolG8Xm0HS+aU54hIDmvyIm5S4kKx6RrPsqRf/fGhMPq1wZSVowWGGbMvg
3zOvteIS0olL7ObUfI+/ZpDxQa47LbVaVtE74TYeOswSA/IaqRr7rV8R3rNyvPQcuWfyD6PeGDKe
1okxB3g2t8eCE8yL9MFeWldbfwITfwZIchGEHyryrFsweBijjYsiYEZbFeY8GHuNxZCqAv9Pw1QA
px12rPnjYX7/HFaTng7u6hN+Ojloh7vTSYtgPY4QUgXx3y5FIptW06VoIWiADeBzWC5ghSgXVm8b
NB0JVT2WGRN0Sh7UjvH8X+fWfs4zWSHyQvMWCJSDs7wuGBbTNwDJWcpcoYv1gHBJvRqq2GvIogmy
X+FSRmTEKn2tZAPNFcVg7m3vUbsbfpx+0CumALxUTYjxRThFLdM86UDendjBs0S5oIooKPcdlwPE
ICCeUuRqQC/LJwKEEIw8NBCVE7m9QLG74XALlXNHgOjC5RXisW9Sg4n3nKUvm6aPpJMBbY1QeqVE
dwcC3/7VFJEljXXWc551g+Uu+87kf42VKuNwSxEhIifMhnFNrt8JB1wz4Qlgw9gWixoASU/H61NN
P9PtRdK6atK1QNxbyW+lD3TnUAcLVlNcl2md/09etYfRnIN8k06Gg16yEcqoGH1Ta64x6j9Lbdsj
fulaqBzaZwnIw69sEEoY1+V/zzG8hU2XrzOP2MJ18j8frbEl5kpyS1+OimjmTtjXRlZpLIlysJlI
upC+kAg1os7nUv5hshlto3K4JaTj+iJOswwEpuR28CA3T+qgdQcIQL39afFuCYkvCd3CTam1blo3
aXl9+7Xm+XgfAKkseJ8EKKZ02EXMcxpARuoctHISXGrb784Gja3fNxQaXcY+vbgXES+m6fijv8fi
3GoKuaiDTk3ERIlLlO3rGGDf85X957t0M/6dn2Rr1ZTGhqoOHv0cxYeYHdHZw8Dc8h6orsebGgp/
Bpih6lq4fn7KPot6KbBui0TCfSNERKaKPU/CkpbP60NWvW9OnO1PMzIwq4um+G4aP3JFPdPhhv85
bgfk0hiIJydDGJR4dOtYpegd7It3pMPHxNc3GDGAVR16v79IMYxLzHgEy2Qwe2e/B+Kf/d5tYOrR
wLN/FX50sPhZ7psfmXzTpo7nAT4JYVTlMxB5e/eyBXazByPQX6O+kdgbud4j2mCmCTqr7Kt9NoOY
twnPyGZTsg5FK+xicMw01d7+bbzgSelh3kaCTcIq+oJP4cOVFwMo99/M0uOMVVSEgcsDVykkM8Yy
b7t3G9M4Cv3x6IBQ0ZtBFxQzs044ZJErtT7RvDjf+945Xiqe4p9RUfox/SV1RUZlsudXibCrH4+0
2HRw+Wpp5iVZpDxnmqD5turXfz3/i7dSNzOOJeT5EAQVfVFryEUryUbTlNqSdyDO27EIGG2Tmgyz
FJ0E3jaZL/E7i7fNK1RvqpBV7tZfoQwk1zaND8XMeROhNTyjqOZ7T+Uo06L9SYLGRiTc9xJ22Otj
eKhnHv1WS80EUigaClHR90jGseoB5SMZUdO5POznPAHmCpanPLG9DwQAF/c/s/dIZEohHBSSwDm9
XjQqeSnavJsr24Ks8BkF5GyO6jWYefgU60BrUnI8o4VTf9yJNQGuxcpY1b9dfa2xBabEhRImEonH
N+z1mjOIGRIVXHe2dRNvkAtk2gCrEIIAvBtPZTmk+7IMj1fotMvXLfoK25fK+LAHvHahCuLnoH2v
/41CUBJjaF70nnmrWxk+Zq0Aol45iPtMBbB8RgnxDLbaQ2r5TcSm4KoV+VXzDTP3SQFLYxCYpc0R
/eSYYYVrj1c9lSysHhyK7itSDL8yrFuWwfi+RRElmUkNYwBUW+F27aR3eZPMlbD7EeZJ6Q9iJKXr
rRG7+NNONA9Wx4eSj1vxugPx99ukLqYped4fMiBNMSxFEeeyEuOH+OkLb6dzqEBwCjrZhCvpuIFJ
fLXnbblRNJGBAfbQ27bz7BAh4lPUcYUzv531lQT56eZJPf7+e703lqfRPPHtIqkwpFdaG6AH7rTD
VQKI+Ih2YIaqnjaMZlwjNDRhOwdwnogjwVSxlDqb+FX5kooJW9ZOFyFYzy0I8gg9qOeJqPYeO/Rq
RXPIBZOhRsOjLTZW+jOwlZnMswPP+cRCIs/Gzbg+DzrMhhQ6cergTB756jsvjriVy6ZXgqOvv8Cx
Pre4Aq6/IDl7TWDYsBO6zWGeDoUU+ROXvUN58VHUhzCCMo+cB0D4SHZ8Zr7RvdmEwgjYPpLnU8p7
zg0T/MGvh+0k81ofFjeuDjZ4uFfrjlbGvdNmgPZj93daU49xT5QoZEfOWTwxmZAKndfP5bsFwQrB
q3M3feH/qrGFCbG0dPQYKVhOktJSL+knlLQi8l6BRrjz/SH6ZxEstb1+fsTQW866DalE55UG6A/m
JxgX25AW1dmicBzdPCDz0WB5SK17JLI5sX0d218y9geSeWKgpCv4du2ko3Fbv7W+WgAbyKYtEQHq
a0nZ3I1KIpuYKRJRr/8MxmwoVofqxLe2mL/p+fv/Vehc6yGXm4ghitlIoiOklzUrD3SKJCwYB6xu
kGFmrh11maK57z/w7v57zsgtu80euGZsnzmBNPH/svuOaHdyneSVE0bNfb9y++CanjWeyOTyRzEi
eofT+3XRoJt7TQeDCjNBXjS2PjHK2XeXdkSpEBBQCBjOeUZULsYv7g/imRz8RLqMdPouY9phdLS4
J4NT5/E+fRqygGSUibik2jVERNX3IMSdsxsIaLFdDnPJJuljVXLqYfvYUUoAKMFzrJxApQjYNXOJ
TPKW7d82SiWv/w0afIQvQlnSdcL3PFqG+yQZKzaLEjbrojhdEf3K5e3cZKKGDIYEvNOkDh/INDD4
SrdgF/eT0WcyZbjObpgsqXnvFPkQZv6ULy3E3CoHkl6d8VyLiZzgdkHWuhi/FipOtKezlsyt1vum
VOYCQOMkkIukK1uInx5QGxZYi9nmix4J4hsj4n8+AICg9+rFhqATP8uaguKw65MnvFLaNOwRCZPq
Ec8ag2Hh6K6FKf5rH5BN+EzTTab7w4LVqtB4bvJ8BRX/W2gknMzar6hvMOydGDpTuNT0M5mZPWzS
b/Nu2Dt1y/EzRYClG1o2EAPlfw9SAfxAlaI7DCM8zSQIk9xHwNvnwNEmgBSK2WqYfMyPxN/h5Yef
bB+sU+rClHt2SzkegLlWMaL9AEqeQ1vdAobVQjDz647YDozAF2BayRBB5kBYKw3AHK15pc3wYHCO
T71nhEgnr6Y8jEEfp2wvcuHm6xDWmgkvzZkrca+fU3j+ZpiW6/c3Lvf1Y/V52EExAbSA5Q8sLNCL
x+lGair99J9mWOOLEzg5OUnFYcOGgFfRK7LvPeOJbhbOfqaOkngaegJ1qy/A591zveh7xNT/imUM
3yTZYP+2U372umrMwEX8FutO+hblUzlfHqhg/KG0YXC/oFAKObKkTbmPgXbIVaH5jIaw9C+JzQ3z
GlUj7ab/wJ/b+2eP4bOLqvOKObvCi+Eoc1oBALCjcflGgsnMPmz6lgmuuxISdGWbOIgeqNtzmCBd
lukvts9vR4SJxGD3dBqSUOo71P5fRLg+CcxA/W5VUElpfHcMZaM8Vqk6S7dGfjCixPKRtk/Df7cp
4l3r7yGvftfbNfKmmmcGYCPoDK/rqbhZWKTcqH0THoBQXT2P1XsUQCC9UBrzutjWp8+jHNUGUYKQ
unUzAqSfHBh9cYZ9nVQL22E68si93B7KzlvHhT0Qr8cg1LoA2OvQcOlAXs1RmhAoJbxkCf3TKWWU
M+8u8kqljHMmpC8acDK/+zzROjGiTSOZQqzvhcpWUpunR61D/UKMewNhnvGMUaqYN+1aBTPAbSrH
iT8iKFLWBl1yeD+7hRCi+BhxpufbKes0ZmFdXkx2PKwPD4BOhe5DLAXWymjxvfQu0SA/WlLWfe2Y
wIO+s9zT5vivhPFqR7m+9vxBK6yoAIEITBZ378r0w72cB2YjN/3p5W/MyFbWN65jQDONDxqiNvJ+
ARXtPjVPaIMC0RgG2wxGo/7CosewPuAD9AaBJ4JAep+mOyo7vhAtQFk0FeOpzq5q7u9cG34Vizpw
Jx2sE+ki0cWK0U7Y324rGyZw+gqtR95B9JSfrvhq/msx5hucbQG5YUz9V3XoJPY/BNMW0x2LWeRW
qb2onF2u9wVxn+oYVcF41llQN5JPoFR3QkobcxA8lTowxgFosd2S1duakZGMptNyuj+jHm9gD+Yb
lvb0b2TuGPF6m/ifLNffkwC2VEogfG3HAXExgLBG9YcCw1QxG789AyHWnTqz1rAGy/YYKwcd1sUi
7nEWDQd/qrgKImsiELwdD/MakLhLXn6txPuloHZEDtYYFrE9e8hmS43x9RwcpxtOoKNPvPAabSaK
rtTystebVKXurYQIem8kezfrvYL0Xs6rqETJ5cXtaJ70VmBHN0qxmqx7sUHJDC7jWLli8ZoSJ7JN
X4iElU0Xpxf3qvk6ahfHDZaKxZXEU5+Rkg8l/l+eb7RoSq2SghHlOLGh/7tCtRV9uLma4g5ugKTz
TUCelf9pwhDBIMIxMi9g9dVfGhlWUGSzOl94cDoOTh08DF8KrMKAfdHww8+HimRl281D+DvNQWfa
jYcNOD6K1wDPi7tYkXlQN7px42MNAh8yTgDoC8KYEpVQP1Le3VYxRj+vZrLlCIYzN026cRu8P2sW
pw/MGZProddj8AdKIlpsNGcYClAM6bjDRmLo7EO5vlQCywND9KRGflcXCGgVcNK1G6ixHwtQmufo
N57ezf9X9ZexC9BysslHmVXgqryMAlWJd/bEJ8iF+KzbI6vKw1Fi8lUgXXnu+H715dnIz0OIrirL
qbNybEZ7JZv6ZS+sz2Bia2VN8t4WzkihPYQz/pDiXNYr+70qzEs6LSXtZA5VG9Dgu0v9iwCz8ICb
GjvHIR/x0fFS55adpW5FCT0noimVkKjCB/rBq3uhwQEJMzlGsxIoZEhIMqJ6Otz5s69kycY87w3E
EL6t38cGUgZZbMxcKGxnpFP7vZ+66b+ght3UQsZ7We6JuP/RZFMCeih0HopOJDubAisAQHzW8rYo
AyLkB2Wjn7pEdjHR6IEh77ruSsxUxbae0q4F7j2WyQklrTOCbTf5ba39ZOXlGsug0CRxVh6E6wJg
hPOqqhQNIuj1zbACSVS/EbLqh6tHg7dV2A+WRTmRaM/Wh+CEbGDkJgYyelFByMPua5cHgAxtE5v4
mooo3nT7n3SfzI23MVZm6d7Fa8uUiEgEryxfUiqPyhKym/Sa/nzFu5E7paaxuzbfm4MyiENQt8lz
wWTt7GnCH1qyX2TlwFGGgAm3fS5LakgwNGJ5Ay5IbeAza0/VwQ+ZFC8MwRefjnZ/ZksJDmpoPRDW
N/HpiymH9bqtY6eGAVx9e3VFWaoEfe+jwVXjGRVyC13qaNe3wmsqVFIJ1NRT3OoblsG7Ldqb3yZ7
WbVvpi8gD/sz7+X1rx43FW6k5kjhwDCfZxk5Nkl+3bL/HKghjiSuX+5Y+xBjDK3xZpkEfbRgCujk
1t9uuQ8YbLGx6NWuG8EO+5Swk4U2h+Xzo7Ore3dSx7rP8YcH+jchJlXppssp4eSUDYfRTzLbaqrh
EZHI1e782Y488/2jL6YleIN7fh8QeRqMt3dV3TOz/vNy1nLEwovSIYrdXh099sQRohLOr/0Uummk
85Qn7vPggdaoj4+1Pqn5dT4l/O2HQzYaYawNE1b42kr9G8BwhNIEEPb+zRSjguZc1ANSuWzx1uvV
bCu0pfTeG0lXSlT8cEQK9V5vv75t6dY4NSVXuIau0vuTGEsy65sFDtn1nXZY/PpFB0oORkCdRVOQ
pazSQ3wR2gawDWJShrxzErU1APjAsJSVCbL7clj3d/yHI8gIxoSP0+/bN6vao3YjKITOcxZXj6rH
/mUKM2gLNj9DNGKXr8vbjoVqIJlvfsNgxY95r9RcsWIi1OuzFVn2r5hUQ6AjJ/wo0f2BjKgF6d7W
k/kJWx5csCwvk+FiwQHHWA==
`protect end_protected
