��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���8ĥE�ZჄ�%�ȹR�CW�:��%�,[g]�`����_�#@�3�A�C7A��*�ۮ�moz���= �l�y�����_�� &���9O��UpR��/����u��Y˹�%[&KɈ�� ;DR�������o���`q�k�:<P!Lm�!�&��!�H�������xi��"�g��چ�[�b����cRn/F��q�R$�ׂ���_��SHxz��j��I9��uT���U�l��bk�m�8n�l��\7�D\��ܥ�����>�*.=�)�Ø��:�0�2�K�Y�_�:�+���Մ�����e]q�l����g�1�hϪ(C�k���HV��+BT�L�Zx1OR�kB�Cή�����c�d�L��f�zCevg4�=&c-!��S����x��D����ٲ�OHo�=1����Nw�^��W5��{Ӕz���O^�C>'Ms���-�e���rgf,��	bJ����@�hq��68�b����B��&��LuMAL(\��p� RJ�Uw������$v=�I!8x�j�.]��
$ړ	�#� 	�s�J6#+~�I�s��N��`�BMT>���Rݳw��_�����?pP�ϽP� "�h%��t���#}�%(���zkV�)L'Qz��-�_"���!<�W6q�2�v1�?��y�۬���=���K���̏L�if1�N���w��[�-8	�0W���x�
��t�.�ġ<��N���Z�;T��˕����D���֐�Hg�ňd4"�y4:���-�dff�eNd�L�`j6��7��2"#�l��v7���-@�*��%���V��LL��z��?���i��=z�SC���q-e�|-~�@�n#�H�d�f\:��I�q����J�D�,n@��0�<���/e4o�V��3�5|\�(u( �}��!���K�4�ȬRe�̸�ǒI�.Z�KP5�&��ED�L3�,%��(o��'gF�ڙ[���[pxı�{XRN�[��pE���j1Í{�^u�i�ea�!�|,�yD��,>�w�Z��X��gAp�V��(`u��s~�r����(2ӀO�+��A�����eB�f�~Y�b?8�r���%K9��|6�g �6�"��{���Ԫ���h��d+Ҷ�P�܏ӑ� ����P���3%;���߉6&{;��ze��g@;������5���yR�8�z�����o�C���P�md�I���N������s�-���9(e����8 A�⥭4y;T3;��~�#=�̬�]u��X٦MH��7����31e����yi�{�\� �h(��qbL`�C<��b���K��i�Pp\��u؅�?�sg��l5�\z�t|b��p����J����R�*f첖�����=���)����e�}eN��㿤ʶ�}8d��8�,�R3���o����X�F�z糺��H':I������j���E�L�YS�غp~�N�{$g�ǲ���n{�G[z����
|e1����n�~������H�fG��Em���^m����I�P0���������8 b��eP�<J/+R[�vC����f��Dp`I�_>�EpN���{�� j'�(�5N*x����~&�X���0��Jζw�����?��(�1���Vc�n}pf!��0~[�J�w� �`�E�����l���	�D�@�M�Ю�hI�4a��b���i �W�})���F9�K�sی��w3�����"���w#� ���-x"5��=h��0�@ �"{|�nbze�u�B�M�I���X��g�ߖ�_�"[����F�X4�$��E1^�
���=8Cr)��r���<�W�֪~{E�|3]�r��e�AM9��r,tr��6^>��\�r�go2����0���H�hE����H�.~-����&	O�J�t��q��O�!d�y��G�YCAan�j�l�J��ơ�_�~<nD�i���A�2���e^���H��>��d������O��N���Y��9�ۭ�*`��דT�ĥ�Vc	�k5��+7*��(��m0��@��9�[4��"^{�*�|�+�2����x��m9�ǽ�պ�(n鋈$��N����<��Ś���VsPMOz�?B1�qt�>� �Hq��`jݔ�@���;W��p&����m2FĨ��z��B8������-O�ف8	,=pX��/�d�-�X�~�~���Kퟨ��׻�[��!Tc�ā*��K��~���1��	^W��G�K.5�<�� ),A���z�	�lyVLI�_|u*Jռ�F��b3�ݟ��;4@������Fb�,h}AɅ&R�Ϛ�ŔaV�Ӂ1������ԗ���c� �w�NC-	�j/���,xw������7�*7ߔ��=V�S�E��Ǆ _�p`��K�%k���i�_E��h|�߈>���d��>��Z� 4�-�'t@�uW' �®⁉h3�Q!:U�~3id@�
�=.|�u/��H�;$"���r����ђ�'gPN�l���`�%Yt�0��@A8��b�A��V���nW{j:�o:����P/J�ō�������o5�+� ��?�h
z��d[�
є�D ���N$�GM�F�$��2?�i]����`b-�#���pzb;�teF�8|�	�9X0��*�~���k	��$�(����,|�'�`S�-�	NYߑ7!�m�w��%Zygş�օ�����zE�Pda]X�Wu�<��<�5�A�V
o����;�3��,	M��B���ۓˊ�4��#�SR�i�OQu��st���y��W8i���<"�x� 41CoX���?E�H��%h�D��BL�٫.䩷͓AA�5 d�e�h�?e
c�cA<A����B(nA���Z�K��r�Gw��B�#�{�Q�`�e
f�Y�mQ*�?R�rS��*��k�����G�Uc(�Iky��e��sMU�<0����m�/v."��������冐A���IHN2L���/���}q��
;\K�6u0\�,��Ğy��(A���j^��>B*)�Ǚ���T�qh�$�xa5_�n�C�lM���M��2�Y��dVn����!X�S��-NF����S�0�4w+ ����{�+���`�m�l+V6d ���Ӈ�S��dguG���E�NV�s���7������'ĺE�K�+�sa��*~VO�}�S$��Ɠf�_"�'�X��y#�{XWJ)�LqX������O�.���h���D���ϏD�BG.X�Q�U,Jb	X�h�n�"�]'$͑<��~)�[�W8��vBLC�@���h
wȴ̡���0Pz�M̵d��T�%T R��`;;�����6������;�X��v)��'����HI��mX�;�2��XA���R.
.��c2��y>�y3��G��dNu��$*�t�J!cpη���p�����V:��G)�W(��i�<5�C���'�|5������l9�x��OO)�
qp�� ��~��bvn�#\0��S��T
+���G(���9���<��Fs�J����~J��y������yBU0 ��,��Q�-?q1�,6��n��)��3IzG��~�u	�ⱟ�Jwb�I���cI�5���8�C�⛐�h��6c��������)�O�=��\1c�F��
R4�UG6�g�a4�����p�Z��!���u	�=�o=�\�B�
y@�|:mV�x�r��cd���H$�	mf�6��K�F���Ad��71�����8�"��i�p� ���0�����`��P�Rx����n��&�I���IY�x8|e�qc����2�}��]%i���DW��yD�K�t0/�
���ش���*�)G��#I�;册���J�=�w�0�ә3J(]�9�����ϩZ9O(@R�K�B�,)N���1��=+-ub<�C{e�ㄠ���e�&��ug*���Jv�?e�v���*�����R��Ҏ�nH����q)�9�����
�:ѨR[\�s�\�n��g��4r�Z�ŝ�-_�Kơ��MԿ�~3`+@*`L<�.^Ƃܤ��D$w+p�I�^�O>��6\MKM
�*a�Q/������HB���_;N�.��.j�r�fg��Tt)����I���� �0�i�f0�8��^���	`�C|Y���^-��U�J��x����C=�yfVO�e�^� $JX���x�(�r�&_I^��\��}a�),S멁kLJ�����|h���\ �R�O��2�2q$>�`�v)�M���"�1iԄ[\�|�eW��荺��AkO�%ޟ�)1���R�9�;��G��h��RQ�]f��j�N1-iB:�K)���T�h�(��BG��WOb[S�jo*ȼ�Ρ:�d�����P���G"���H�Ӏ�
�����r7|Ӂ�o�vP�־hD�<8��!�o;���l��'I�~6O��j��)L�B�����p�S�/8F�,��=��*�v�
B]?h��¶sS�L#���@�/�>;����>l���H��a��+����ݐ�������ܮҕW���\u�OwP�g�o������{��/s�'�|� �q��&)Ac�u&�,\���@s�|��#JU��ը����D�Ē��3lv�@�����9W����<�[2�Ce�.�S|�b��+��bz5� >�Oŉ�v�C��U
����K�+Vԙ}�v����0FU��s=%{.�`'��]M�3�*{�|M�X��%M*8���"��\���J��zM���&23I�p�=ydɳ������{5�}:�;�jm��H6���jq��ϋ�bz���	����b����P�=E�������,of�@ �|
m���6,�E9[.L>�2�7��U�xM��4��R��݇����z僜
����
4�����u��,W�t�|~r(�x˓��e>6r�v����⫱oѲ��{Tq凜�VOh_����o$r�1Y/I*�'���.�k�Ejש8x����Hm3r^�b�l;�� 7:��GU䊰|P�Ty�W�88X�
ہ A�ŧy��P�FPN��c��xM����1t�m�`o	UMHך��D$�.%�%�f`>N�9Mo��onz����q1-�
���9�s�r u�bU;�>��f.ݫ�i�,$�t�Y��c��9�8�ɹ�L���9�	�*��*�2,w�ִ�F،۲�h�b��[\�n�i�h~R�A��;w��U���N�9~�7PPj�h����$[5�BJ@���w1NDQ���{5�u�u̧A����l/ѻ��wU�UI'1m[���1���gqmǻ�(������t-u�m�*����Jm`���͚ns�7�r��9�[�A��*h���z�cl}��ѡ��:5c"���nV�Z�v4sLC�&
��F�dOT� �8N��I~p��<Y�%*BLsFTK/�^��V�~r�I�5�Z���]�"!	#��սbfZ�*��QN�!��f��(��m�qTR] �R���%���C����,o��?`���#��x��d@?�J�cfgx>��,�h,@�>չSN5����Ѩ'���eL��oݔ���D���-����+�H��pgfR$v��5�/�B�������E�_V��^s�S6��)+Frz_�'�Joi��s��\񓋸9x���@{�%��O
��I+{B"L�b٫k��m0�{��*v�s�i���=���	J���hƣ��|��
��f>�靟��%�+)yV������&X����V]�#*V�UԾ�)c_�6JI��E\��[�Z�l[�2]*����������X�CA�4�]���f�ʝ-��}M����([2��j?1�;ͬR�����Zg�T�-�1�9ã��t�������_=H����rgI+��$X���ksR� c_�Bp��(I�\�*
���$��[�:�d������RKo�st��s�2*7v�NCXIHCث�}sĺ��xɊ󯍁�dk2�Q�y��6��Eod��Y��*"i5�&�dZ�M����|�< 8b�QY~4�'�4&1�����|������4�5����y�%,���*�T_/{�cLI��P+��c�)�G͐��A��(���y��dR��L�E�;x+��Mv!q1��=��2^�����5�I�hH%�IDH�9��N{[�%�r=��/��hFBl�I��_QJ��`�9'0L��m����W�$��߆f
|�#�Jh	
J����/Ʀ� ��1�&v�f�@��ɟG�%
� 9�������oi|�0Y�j��?�إ�~�//��)�$�7w^1��ڊ�P;�����^�xq�5Īr����U>��;G����<�$�DBU��m1�D��>�$�����CC�]�d0��(X��幥=(������6�x�Ew�ɖ�Q��M��xv�;���'�G��4��^t����u��e��/��1��Y4|N�	��C�]ܲ\�r��Nɓ��_�`����?�*{�P�J�����lC-v8�~��
�3�P_�rS7�
]A�^��` E��8W��IUx˴|e��/ktx ^���A��^PH{�����L�& ���#�Q�ԯ;~��Qk��Gj�`�$��JvRi�	76X��>C k� ���1��� ��p�22`��j?M�-
�h�ed�yh-n:02�Xt�ɐ�MC!'d�-9b΁OM��Z�d�l�����G��dP��^�QQ������s������I,S�b�T�����B]�P�ʳ��5��c�{P���	�9	�z3Z:������̋�-q�$V��O�
����<I��k����Z�Fì���O�l0)@�G�x��O㖩�nPB�&�eme8k�u7MI7ǜ����������e<ϙm锉� ��8��Ǫ�u�(���4��đ��(@_L(qQ� }��GȆ]�"� ��ɣ,�1�yԓ�~ClJ�Gz�#�
���H�-�f{V���V���Lh�E��.���F1�Ѓ��O����o���]rg
��٧��y�~�<���׳�Χm)%uaa���u��J���{��ɵU0T�@�����i���ß����cv`WWt9�'�ܛ)Zp��r-v��P`~4���Q&�1���~}�g�9���G�͍
ݏW-(聢1�}�_!O}����e���gF��KX*0�����p�V@r�If�b����wh`��%��������<Y�P?Q|I�`�XT3����S�؎�w��h޸�BZ��L�].�d��m+7�	>���@�;7�c�H���O#�����g>9�ZNO���Z��t�C.(u��E�O\����"[�t�.���C�k�m�O)8�f�GOnz�t�`�rN}���<�~�o�+k��vḱh�㒟�[ ��}��2��ǧmq�[�RX/�̀+}������c�˲16W�
�8��^�?�հ�����(����]@s ��j�l��-�.h-���u�;oD�l�?��$�70c�kY���� ��/���\���w*�|B�EX'��� ��4Hk�n�epտ-�k^�q�G�〗�$�,�sb��j�B�􂺔��Mk٠3:N�f)�W�1��$�ʸ���J������P5U�;�.ȗ|:�ܻ�����a��Z6V4��p"{ؚQm����.��U��+�J'�L�/8c�u�5(�\_,�5������N�����s��1G�#cͤYC}"�k�2��T�融i�;?瀿��|2����ѲZ[d��k;}�C܆�	�Ȍ<Icqw3ͮ!x�A��"�ǲ����S�F�k��
p�>p(��ɥ�FYfڋJ�&ܥ����Yg���EEnn�Ex�Λ@
SE!n�/'�&|I}�H� �	LOߏ��!�B?����*,��ꎐ��J@�nZ��
,�֝_�B3�G]�ұ��*4��ۢ�h��I��\������U%�"�!��jA~
���޸���:�ecmv�p���4W�:=`����x크�����Hf�����olqdj���vZ&�]<u�E�����'�<0_�d��>�0��B�Q%�%��MJ��#���Ǻ� G6�k�Z���0�Q����[�L:�)؍"��8i�A�d.w��2���7s�v�`%��g�v;�("p�|�Ąö��a��:�"����	�'f����*����௥kD�ϕ��//c=w?���#� ͢(�(� Ǭ���p%�g(`�tә�*��#?I=��r��	��1����a��M>�㟗�b;`{��]��Һ�H"���V)wL�Sb��jI��Y&-��p��F�F�k����	�������e��"�K�:����3E+iZ��~�:?<H^�Wo�r�`�KO�n��쌔��롗K�a���},�N���0ٌ�o���AbQQm���p)��M�.-�MD�;�C ��7��px;YU���6�%�$=;<}Ӿ�#�ɻ��L˒�`��ϳ$P��'��Un�����,���3����v���A�U�W4�ʽ?+s�e �C&\�9(W_ =��~�
��QbS��X�d�/:)©p��m�Xܚ���������(3��Nj~
�7eC�S��~�h
��f$�DUX����[/�h�"SM��&��k� o!��Ps%���c�������F���Mɵ�d<HB�)�hV8|�D����Y��Һ�_*C����� eT�T42sc�8M�Ϣ��vm/��|����vu�s���a@�Կ�O����z�l[�H�6���U�A�-ғ7�M/�� �l��"�s�'C\�-�58y�F��8������gʣ8jh�<��6D[����,�lh��B>�$="�{�3F�GF����a�ή�x˰�A�%1�=�~e�J��ڿ�y�ޟ��ÙϬ�!0-� ޛ�SvW�k#����B��y����y7J0���X9wӶ��d��v4D[-�4����w�c,m��d]��.?��i��#0'd)�S'%�ޔ�(ꕽ��	@+�%�3-(���!O}�v��&�u����G.ד��gј�����i�\�U$.������[�r}�e"J3��C�P� F[�I�6��%�P��ͨ��~3�w�ϋ�(�.��Y� N�5�r*9	?�-��CE%�+�1�FmŗOt�=��Ns�>O�P�Ҽ�f3'��{l,���χ̧G�:R�*P���=yl@�tD�X��mIG��
��մB.�NK����U�8 �:�uLʊ\W�i3���W��)�W:�X�|����E4k�@�HA�r����b�.���u`�Q�o��p��n�8�i{��^�'ިl)3o�i�J� ���D�nl�0~0�]�t� ��pPk3A���2�0��"��*�h��'��9�����:�C�Q�,�O7e���N8��i�G2nOHU��AtXkL�x<v�9ֹ����J��˵𼼹M�`Z&I��.�o�&�e�
C�!�O���^Ə�M���9*'�J��b�M:���)����(�x��̮i���gW)����uE�%Ʃ%4�H��%#�[QI��.01y�^s.w�1&�i�z9�^�tb
-�s��M4�u������b9ي�kP'��rH�o�Ug���������D8�1�V��>Yt��)�˺S��(�Mc�g�?�kߨ=i�Ć"�.��h�����x>B�\v�?z�'R��a�^��KӀ�P���|�̄:�Ue�,���~� x�}C�?vC��
/�-vd|�ka4"���,X��}^���KLFT�s_��_����9V���|��	{̠�ݙ��5���R����Q�]��5�}�
<Jp������Lyc6k-��cDq���T��g�(�b���B��-��W@\,^6�}I!8`�Kb���=&L�;6�w:)��{xņ���`K��`��C�E�p��Sh��vm�uUk~F������g���/߀�܄���s JhsW� sEH�ĳQ�Fl���m1�T�9��l��{j0����%l0ȪQ���,cDȘ�/��䷼���C�u��nV{1�6�G���S­���Y"rOC"��mcW��+r+x�B�1o�GQ���b�V�&*w�z�H�A�W�\� |;V�h-y�^��?���.�ۋ�z�����;�V�UH�FK=\3L�;�Y���T�@�t���_**�7Mf�x̑��	T	�PzCݱz3J����7��-�K�8�d�����tٮ�l!�T,��]��v 7c�#X�U��
��7��d���?r�/��r���tA^Q&�������ˤ�l�M(�Ԛ1�}0U�ڙA��)�����"/[���. �xW(����}��� �=x�c�`+�#V�,8���ആ�:�d��3<�%N%Fo-D��E�犮��צ" I>��>v"C �1q~������B�e
�14t�}�R��]�����:z��PՈXO�E��䀵URh�p㉡"z��
Q���-����&��7ե�u���rj�*qf�����g�Q��K�y��J�ܘJKT/��&D/�n[�l��`�
�m0�o�Y0�G6L�V��Y:��}�|��D��Q	�0T�u�^��߿r?��Q��n��Zv�3�Mc�	e&�]�'�|f�a1z{�Zŭ��5���O42h�H��o��"8���`k�:(�J��{'�7��܏)Ǧ�ײ�������G; 	-���-囅�Gb���LS+v�?�h�̗Ɛ�Q���pS�n�*�U#�;�����2C��]XFFy����F�n���GY�@U�Od8���+O���R��-�R'���P���t1����{y�C�o(=�b8��T�����{)���EY�K�����Ͷgx�D����� �������[՗������#"�)�6������[޴ick�Ց��g�;�)�v��h����1���C�)n��ʫ�̌��t�T!)G��~o�J�ݣ���I������o/����MoxG�O������F@�8{Y$�t&e ٗ;b����x`I� P{����-���K0��6�Q����?��>�'��>U� `))��.Xﰆ���R�8l�v���kB�s?��~��x�\҂\5[j�'�2�5�m9�=�Q�R�b9�0��j?G7�wGg�ב���q\Dt=!��X�#�ޢ�X�}���M��R� [��)��HL?�P�J��" ��0��_�Cp���c�8�
:le_|�{}�i��{��㪐�XB��I�	�/f����)�]��<��.}��u�H�k�vh���˷׳�����F��Ȓ�*�1�qqw/;p�A9��(��lE��<����1f��Z�F�_�W�5.>ʨ
���B����ũ��db�6�\��8�M����7�����Ă�)h�L/������K�ݒ�z|&��Kde��;f� EA�x���g�Ǖ��³
#�� �2,.������ȍp�g���,�
���O.R���NJȴ���<$�c�	�v�� m6&mW ��x� ������T�h��O,�<\�p�k��2<;�߯^����x�h�Üt,ꮞ���rq�ݳ���n��87��e��e��d��Dט�6�v�v�
�CL���@��Lݥj_DSCy�I�����D���!���@�͢���~��Ŧ��S�|UD�5ի[i�ͨn�2Ʊ��S�l�Ǫ!Qi+�=2�i�j<�9��U����4���&�t�W���9�y�\�UR��P��i�oO�����0af��,��&`HIM����:qD[Iq��������g(���*��a�N�p�;+ �B�_�힖����;�!��)����I��bu�ϙV��>�H�M�T�3 &x��l�1I!�F��Ͱc���`����A�8�mEҗr���n&�2L6�1�8K�Ĝ����{�-2��5��D�)�DW����4�;w�i��<H�Q�`�w��@�Tad_�o%�ܟC���k��&�za���(-�(G�:��[�M�V�z���CWǛ n�Mł5�H('D�JQ.�¶@|�ö ��S '�C��Z-����ߓ��������ҷڌ[��C����-�ayu2%��ኡw��Ni(FlQ2\��ڢ��+�
��*��]r��@y���IA���䌜��)������ ש ���%�k���-�K�>��B�7��'��鿬��KH���*�De�VNe��w�_����jY6���0�<�TI8,So:av- +�؝��}VV��J'a1�C�i傞�k�G�jO���V(P��H㛚�t�j^AS.�k��K�}��*R�`�����C! ��t�������@�P�hx�x�1?/nbNh���O�N����;Ε}CX�ŗil��D�I����O�U���F��7�h�-��S,0�9���5�+6�邠n�1����sk�g���uV�J�di��|k!��8k��77�Q,r"/Q��,]/���L(��A'�c�p"�e��K��۴�F�ūf_&���j��'�zTucOq{M�xcS`�D�����:�����I¼ ��LIhô���kd�G�ؾ�.x���}��iؑ�0�yU���6 >s����As;��g|L��$�������~���'N�F���x&���[\������Wz��CC�%��Bn���T���_E�[n ���d��`��ծ�B��C�q�
�� j� d�#ь�$h��[��"��ߐO �
?Lz#�#,ǵ�Y�qp�C_Tu|S��@�O�p�bKD=�Y��q�z�����w�(����w�ϗ�|�.���R-��N�i�R)_�N�Ј�ϊ��#_tצ-#b�:��!pR��s�}�������Z��Qt�������̾���]�
:���%I����}���>`)���۰[��VQ���u�6`u3��|d26>�P�)�sul:����U��ܲU�V�$U�sY���s��}`0E�ҩ*=>(^�kcV|����r���C@ݓ��U��MW��hXHs~evYI�+?ky��N����yC�s���Ӄ����Cp����<oc��#�s��߃rS�pdN46O��DD�R�5 Y}A߂8���.Q��cԌ x^�*�[[��_0�r�S�r�ʝ�O���8�J(e������AQ.����N������v�	w$��Q��E���>�������[4��K�>X��A*�-��Tџ�uxfA�5��k�uIR�m������#?�pk*\����LV��������J��l��t��@Dba�=�䟬���V8Gje�,�:	��e����)_����.Rg)�
�99�.��T-a�&�|��F�R��?Nl�p���כ�My˔���.����B��%l4�R�"�.v}��,kNk�;��o8��$�2/)\�v|w+>��.���=���mrQ��~���A��@^��bo� �+h�q�e��E\��GQ��H-r�B���q��OkԺ
�Z�'0*��r��*}	���t�|����f�����A
]��}f��Ғ�Γ��������z�d`S���u�������%������#5�q�ͺ��r^\|�QQw�L^�ӭ��~��l�&?�17��^6Ƴ���RP����h"C��'�_
�+����n�  �OEDw�;+xY��灛�y"�v��
��׻��N(޳̉�G�S���$�9u�@OY���0����|?�z���.Q'���,Y��������LD_�C��.�Do�YFq������Yh��`� G]�Qһ��Ty&���!X�r����n�L�/mɹA;?����?�+�eW�&m��o�b�=�e���ݳhN?����k{�W�s+��>�� �eՌ��a&!yc$8��~$�9<fG/��l�y7���d;#�}�Pt(ߺ
MOh;���#����E�S��
�Ήa��f��O��3�?��U����H<L��[~���:�?�eP%�0<��cZ�<�t��)�L���9�ܝ��t�����X�Z� ��O���	#�4�� s�V���Y���N��AZ��m�C�5�*�n�!��~����Wn��4n'�����A7��, �t=8r����jKaח��15��<�9@���al�J���Ȑ���ʡFN.l%�T��g��[�0�jD.W��a��IyONۭ&47�MM�6���f�e�df�e9D'Bk�9��^��ո�s ��˝n���k�wC]ל	�\���^Q�u�s�T?|�i��8�x�c���E��N��-��vA�捪�qP����ĥt�yȽ�_�t���Q�+.七����2�۵����ψi��:��7��Vj���V�Ҝ���"@M|�k���?�a���f=9唼(�C��R{�Qc��!K ۹Ի��l��W�1C��d����Y��觚|�����g�p��v>6A��v~���'�ѝ	��#1���X�eM� 瀋��8]tV9k\5:���_C�&�,�yhI�.�|=�j����9�1& '�IU�E�,����u[f&W` A�����Ң���d�5+�!�&������b2�3�,��q�~�{��wq�E+;��毃�-rq$S�h�y��M�rg�β�Pɯȫ��c6׋�"�tRZTv���|R��޹�=Oҽ:���uwA�]���� R$��#� �l�~�����`��k��D�;�+�Ԝ�[z��l��C�$ba~��:�fv���gT�m��6]Y��J\�������~�/=k�'��>1��ǅ���Ʌ팰�U��L"p�|-?��B����}_XI��k^���di��y����!^���8w=��N�v�,��U��0����OLR����c������yJn�$��<�VM�y���O��M�_}���H��S���&�[xt}�g�?���{ץ���<�
��*��^a7�>������C"�,J0�
�[�baN�τ�9��Y�fȨ:atB�$�����i\қ�f�|�c �I���1���k5@`�T�f�&��3�b£��r����0���pG���<7�DB{b'���Nf��O��[
���Mt/=��+/eGfL?y���G���(���-Q�b�y�!�� ]C��TLR�W=�e
�"RY,z�I�4��/'&�� ����'��d,<���~�_�e���0@	llޯ%S~�p.�q�����Y�:�2���6	���e�=yŹVr�9f�A����љ4�ckyIA�(~iЈ��3p��<�M�����f/�{�3��4y��G9 ��z���'y� N0V�cyS��aC�:��K�\s�n�BR�C!?�]�0�9�Ǳ%g�����A�����}D}Y�oK�_�p.4��{"[��礆Y������\i�E7xvHwS���-��U�C�d�����Y^1BF�����(��k�1��;ޅ�7�*�@���bOh�+[��.F^�T6�'i�q��
F�qC��D67E�Y����7.ZԬI_1#�KI��MGW���I���̡u�yi1��%S�4�α0�J��왽:��xm�m9(G}a_G���F9]^_���[���l��%��}����_�E��,��'�,��WkG����Q�P,UPjxx}�_���I���&�~� ����(&l��)⎆j���a����-<;\��<��2N(���|�����]Y`S�U����1)V0�M�M���{��!��`�'��lA�-�� Ҟ���ELU�7$��98yQ�)[�������bQ�������L����(�o�?x��u;���=�N|~ ����$���N.�˝h%��4Y����ߧ]�����	a*�%-Iz���u$��҈6qKM��%��-�ɽ<?Q>)��r�'��H�θ ���=���?쯕��sެ�l��>�'e�̷1:.w�z��2�i%��$leU��_@�D<�����Q�O�c,H�Ax2nB�Z�� ��ER�\�
����>���6rx#^�(G���	�o��&��G؇s>߉6\q��F��<7zM2����σ#!v��V1��b R�-�v$��q��R�;5PD#4ԯ=�"��{#g�\ث���j����W��I�����^̾����8�a��L�XP�	�Ri��~�&ca�)�>8�@Qg�(ߙ��,O2L�|&/M���]7�[�?��
�kN�Iz
z*���j�7p�j�Ξʨ<l��Ʀ,pD� ��Ԋ~�N�?�h�NW����c٨��f��R��0�4mM�/�Ѣʈ�c^���R7l�=���0R���5�L�,���ari�Ֆ���Ё(��ܻ>;Ĺ�F�zQWt,�������A� w�v����\��^�nC��J�*�i��	���P���|YOS��gR�iO�ވ����릸��k|�`()f�K��+:��;7 ��@��A�d��1�����VSd�ۥ>��<ZL�W�\�Rp��%&n���%Z>�~��R�����D���h��=���*����Y0:yċ������9�$�<�fys�+��_���Q�VL_g���ϖ���}�	 �i$�ng��5��������2���)�Ė���-�4G����jRO�P�,�ng�(�w��q�G�0��,��8���������t�F�=�r)ND���� ��~�j��ϳ�w:���Ƒ�4CE��ߛR[B��y[�[��I�(uR-�\Y��-��ƌ� �ױcg(07Ď!1S�P��!�9E�������q>T�gǒ)w�5^B(D�7<�/��������P��Mc�$qGw!��xCəj��UټG�-'�i�(l:'�\���1!HS��}�!��&��?C%#�LP��f�k/��S�x����Vg*/���t�
���F��!]�*��_�B�� �`��q���]�7�%'��1ڢE�yņ�Չ�T��p�엃8{G�g}��Z�vș�@R:[��;#�*�Vw�*��՟טg���ۙ�ɷ�f9������ ��i��vUHm�7��(
��R)����j`�r�Pp)�m�/޽�]:!�������%I�T�%`�YY��z�w������8�2�tz|X�Ϫ���漤�	�/���7%`TN���"��1y��|p\2e=�O��f3� ���¦��p?-�.guOʠ^�h�H����2�n�Ɩ�0O��
�*J
�Q��َ�=�60�X��S����SӶ�tZ%=Q��[J�o����%��R����i}�Q3���a���"�ׂ�m�+9��7��r������l}ٹjNj#{�	52ʁ�"����f��^��1M��"�7�YZv搡%j2j}�o�I�6�Ys�Z;G�1�=\�l�E�R�烌�p���B�e붿��}[ad�����L`��d0۶��j��z�M��US���/��X���^&������{�5�R�K����%������h�E�ҹ��`��h�48�bU��~B�1/̱������U�	�@6^R
�*^\'V�/�#KS�PnoK�z�<Ia\���)��a�����yD��AI$p')�>-�3:SX��д��ʨ�vha{<����x�
k�vl~{O�T�[i����7Y�t5������{�*��n����B}��p��x`ݨV
�8�ХRb+�J��wĄ��6-��:H�8�e�z(4id�|�C
S�_r)�s8|�7�7n_7�	���fΫ��/v&��	��W_����!���"���>�P��:L�iN�[UK݊�lb[�`�I܎�Կ��m�G��V.���y��Ǧ�˲��i�/Y8��eW�Y���8I-�� s�����eYD�-Y.�B/��M���̲�$�$F ����Pd���/j�ꓥ�Aҍ�m^��=�v���k=]��CV����!������[f~"��шu���,f�
v�&�.{����a��
L�y(N�ߦ�Q���f@XA��Bѐ�jF.p��s@_�-�"E}d�g<���s�0�zn�d��c�v6�h��hGݍ��s����&4�s�D'Ɠ��n΋����ߛo�y���ҩ$E�n:qÔ_H�
t�1Zv���7T��֪��t�i��y�B�s)�L���C�ݐUq%��V���o�ys����w��Q��~c�q���X���V����p� $�.�bO	;.���z�J"���y��$�T�9_:v�����vq	)ִ��phE�inL�~b��#�:�A�g�L��`�wϼh�T���jEv%�؆a��ڗ��H�v#�@N<h6g��~쓠l��:�x��\�������^Si>U.�5�7Fb�=�@���?6���>�b�bd{Q�e��?��Dt�r�B�VEO��b�k|��M���#�k̡��e5b�0���G4��C��z�����f�j����X��*.sͫ�����!��L�	�������=��6\Ů^��
�Ks�������V���o�W�*��Q�O�T��(i�Vd@GtinM���9,ꄙǢ��5�O+�bj�n����n��bv|�dӘ����"�:府v5�5��ݮ�w�Cq�Z4��&�\(Y�>k:N���.+�xvBu���B`�%{XYnM�!R52����|]���|Np�Y�U�2�IK���Le�Ĉ���7_޹h/T��z���I�թ�Q�U�+��ř f����&�WO��G�C�"]���C��f1��C��(��:��
��D�w~M�V����q7�h�	q���z�0�R�F73��ђ��2��3����6&9��~�+O�x��d�ٙ���m�E�����_EΆl�������4<b+�l��͌	����B���������jDd�&�H��.�n��~X��u�\Ȅe%@��D�	��i$˄�P'kN����c�IPl�9��P���?�����Z�-�
n�w�1&�P{�60.�1b����/AMT��u��V�尷<d��/�3�y@so$�n~.a�@L�{�5�C4���	]�B����F�Nv.�AnXl��]�n�\��wOiA<U����qGq/�0�ᆣ��3}|�Yc��N���9�w�)h!���bg�Y��*n��#�dX*���?�M��01+��Z���0;'��jq�l�X�
���A����>�z�`j/���A2��	P�l���Ss7�KA��C��W���ߵ������J6!�D�΢�36�O0�O%q�.��+'mD
Y�s6���Q^��
�ٵ��؞05���$���rݒ�hU�m �	g��|�!C�� wEM�=��Ǡ��g('2i��s�)(*m��!�@6�0����п?�n���H�iU�μ�A~P42��𿜜�����i���x8�JE�&ܨ�%5���!Ez���,�F��e�䌍@�<�y�h<�U�'s�����
�m[f�Hg���g��������4Rh�l�'iஆ���7�q����g�qd���#�dE9p���,�x�K;�$jl�rpԴ��Sw8�'�-�#5cy2wv[\�A��2��8cs�gQ�������X��{��-fm5|q�%�~��7��'\�0&��+�ЪN��@;���'ߗ\�����v(��_�6��}}�VF�б-���k��U�y�]��F1��@��鵜���Pڳ�5���^'�|�{3�QN�=Q���d8 ��7�x���h$�/�K�
�^�̀�p�e�쁣z��QU��'� Ԓ��B'�	dM2�0t������z_L�xo�����Q��X�]yH,����e�E��%���Ө@��)�d��JDY�D+\<��E��Z
+�M�>�
�*O{=rڳ�q���pG�oq�qۙvO�iuK���&��{H�������tV�Dc��/��lۇ���$�S+��U����Iv�t6ٞL,j����v�휗ّ�>W�l�	^��@>���~&)����$9�^W�+��15a' ��og6�q
���V�BD_}^�d�$��֔���� �jfO0o�/���ظ4%q���s���c��\��9�Z���'V>����)�
�Ef�4M�U&�#�~ ~�"_�$�"C�~<�h������lVޛr���j%C��R�+1��"Zz[�=;��"{��
iW�����gZ�s9F*���J�:fl�RFYC 1[,Y��N2v��7ؼ��׶v����M�B
���c
�����3��7�eْ�����i줏��?Jz�B�@娄|�J�_���-��{}�@	�I�����|�#���6����h�@�M�
���մ�JqܟQ!��(�a�6�h]�ɔ�ƚ�﬛a�,[h��OX@�L�~C|���2~�Ġܥ�4X����� t��]q��O��<��%x?�ƪ\��Ю� �h�>�ʷ�����9�V��UČ7n�b��4W 9�@��'�id *�ygw���=?��;�56Ԙ��=,���ʹu����0V�cR��`߾
�H�l�)Fˌ@�x?I��{���T��1wb>�H�*
�O��?f��-��V���^�+�e����m{�(F�ϺT�[��zxb}�r���Db:IO$��Ψ��V�EcoV��eT8!}|�S��@@..h��V���_l�F� ����[ c��bL����-�+���~���1i�D�Y�-&j!w��_�I�$z[�Ӝ*�|����#�J+������r"�Th�o�<~������8~����?z��T�
񍸖HEwr���^E��[<����k�����2ǻY��o��+��B����韧.9��*�$�&��1N�4��o�O�k�F�x�S�z�|ܠk~�LY�y�_%%�vl!�{��偻�0η���Y�)'�)�4>ipb�F?E�	$�[g0*��Aw�hmvV�q�,�4��4�q�0"
I��L�t�/ݝU��p%*���`��&�����A���7Q�ѡ5 ��-�p'D���T�QQ��&V�j�T6�∓D�]5�n�L�<�i��ߒȄ7<jSxX��)f��"٫B"i:<�r�(䣪+ ��ȷ����0�C����e�W9�Pl���^m'��]ϺH�A��x�^��Uy(���H�Xc�!!18T��ӫ�.�,ͮ�dʨ��j�r�M,J�������ٷ�ځ�4�Uzi�{��^��*Wj��(��c	q%�5�+�!N�w��	���}�9�=/X��Ob�T�%���7�Ճ�Ej��iGb��+:�!��o��b������~ڀ�bO�����*�VzJ��T�7��NK�2���x��@'s�&7(q����k(��N��O�͊�N��@j��w�]�M)G�xr��"ds�w-z9����,9�����C���5~��q?Nm�'�����.��H��r��L�b��ǊuR�,���;Ѷ��#�G����J�1d.��"���>��Uq^�;�� �J9x� #���
jv��2
G,��݌3�;�f��*WT����� �[n��y\	I}A��v�K6�^���[�D����M�F��\�t�=��dz�Յ�� f���5Y>�G�;c�G˒N|�6�ڟ���.���t������$j�4BĮ ��!��Ń�����/��� ^Q��%�D���@gjj��;y`
���a���P]]��@�'rEs��N%�	��=��}�w$��b*^��/6��KX"yT�M\�P���1ݎ�>�	J�ۊxh~�e(���6ֽa 6w
�oaE5p��T�Ƙ�m���R�j4?(|�?(��K�	����>O�\@�R Q�����j	�3�^���G���a���p%���>X�%�-8��s�O�V+hm��L�gL3�~	�&Dt��ܛe�7��Qh+���zi��^>�ud
�Y���>�����a���n�@�z�Li�m?Ѩ���0��r��~a����Ci�R�|���V��ג�ӣ��yƫ#џ���Z����_�S5��_����;�t��Ps�:����I@6��!����j=�!y��LR�)AVp��p��g	�YM������i���r����+\����h��dt�j䞸\̹��ѣ١ýz;D�4�V�'X�r�){_���C���5䝀�o�G��C�m�!�ߦ,+����-d�,VT6�^5�Q�� a���-a�D����P����[���� ��%�z|�c%f��S�����#2�Ӥ����-9�|�H*��!�6ׁ�T�����'6gGR�+�N�8A��;PY��X���bx�V1�_rbѪ���΄4�#�+p��J��4VQeh�buaw׬���]�I����2>��M��9ր/{t�G�kq:#��1+��MG��~��X\�,���r +��JZm���Dl�Y)(G��+�����8�M�g<s`X�R�]�����r�K�~e���ѝ �z�w�뇰���g��_�a�L�p�����b�P�tb�RF&����^*��h�!�z}�I��d�S޴�2����M4�Ia8r����Bݘݫ7���E��B�΢�n�"C\8X�e������Α�"2�(��(���a�J�rf��[D0��bJ.��cUP0n|rwK��������'��1��C���=���=�(Tx���H*M�E�����Z�+F������W$�O�z��C�u�t܅�\k������E|� �R�Y�c~:&������k��if�N�1ӣ�4RaG��i�P?-�n+3���T"���;x��[�/��i�H�@���{��qY^1&�_� &���Y��U�&;��x�m����c`�[w`��X ��յ����S�afX���������#%�f����U�$�����er�i���[N؛�V���7sm��_�3 �M�\�߆��!�[��a
�Tؿ�77�RQ]kN&{���#�E�TW�zS����M������hQ ����ίb�����Iې����D5�<�V�m��]�(�7�����޽1ul^�裚OH[�(E	�ݢ�l�Η������ݲ�)�#,�<�{�%����v;Ų.��<���9�k{BFq�*0�{V�yQY5����h�v.it�Q��B˫6�?��Y㽮 Ώ���u+��ts�.��l�����v�<���X�Hu9��+��QU�A��\��ٙ˫�y�-(��J��7�7��tsn����3��j���䅃���,��P�}���χL�F��_b�m-t��\ai�(k�'���-�f��7�Y8�@�
��ڍ�<�`�"3*�V���lіu��Ʌn��$�hĽ�"�)/*���kS.�%sBe)k�J����Y]��w�����\��I��#�IKKV��f-�J�vت�'E��w����Y����d���)♗�/��^>���}�b��\u��1��j"�K�#���(,=	�:$��Ё�D��O=σ�6v��`�0&~�JT=���z�"���
� �ʠWVh��m��	'\f�(�Ti8_��L+H��e%����@����h�(1�!��WX���bN�Zf��g�l2�����L̡�?k�56%	.��Zp0&��%Q ���li���B����$K����n�n�+�t>;W0H�V_���O��ˆY[�Z�u�M��Zf�8��c['���3�b�X����𢀐F��A�)|"�e�
R\!e͘����� �����0�4� b���[��M���+�������<s�'E�~�L��NXM������+^j-�R��@��o*�|�И�uN6�Ww�!���jg�;~���3(�o~ѽ'~�0}��U~-�Vӈ��)�v���*;����+DK����� }����[�����o8OP�er����4���8�J�uU�zӦE'�K��(j� Y��Xd��Dq	y>!��|u��d�M�D�Ӈ�>!����PW�'���r�5C�{�B�����6��b��z,_��ٚs�26P#��Z����t)3*��}���ާg��D��W9'��WZ��'=(�O���71_R .�>$�����O�jߜ��	9"��׎���}��{�u,Iϐ�,b��2���FxJ<MpW�SաSjA�QJx��}���YsT�w��DH砜`tE�Ҵ����䬺�a���57��V�8��V��S^Rǆ�p�-S��:p��Ax<�k#o�ե
���76��4֛(��|W�_-쥽�'�̝�8m�ȵA��2Yk���W	�V�z���I_x��p���麾�4M�'�)z	�'�Ӛl�<�`����a(���S��Ťbs0kS�?��A�l���=�2�q��J��\c�:�V�a���۝L���I U��ו�iD��`$ٿL�M����
�F���	m�_���,�I�K�d���T�!	�gNA�5nL�C�%�*��,ĵ��?�l�.�\X��9-��Q>�j�)������0��].���]�,�:q��>���OaD�ʊ��M2ï�jk+��v^�4o�m����_�;N��G���q3��>k{��,�"J��B|�V��ǒY�X�'�� �=�������C���:�UB^|����5�k�^K�e���24$� �)�7��88����@���;�)� o,������Drk��=���{�CN�-��r�],���' zI^1"�+��~Ht�k�(��	�)�&'@�C
�;�,:����Kn��R�Ǔ#�{����;����ih�Q���̋�G�<go�Z��F�1ȉ���i��rԵaUX�KF@F������t������P�B?l�����
�&Q5	m�h�r�̔/{��a���������*@��Ko����W�К�8Ȼ�({=+�,��_�� ��)�ì<���r�o��o�e1^T�=�F7MĜ��u@�kx���N��H�	F)�բ�:+m��"� n�{�c�y�� J�0`f�x�����9e�������.~��~�Ў����r�3�U�H9?�_�Hq�X�\�y���#K�Q�!�2�!�XrH=2���G��r���\�8���xᷯ��Oз��R��|����m�C[��h���<��m��������'�����4��<�W{M��d}��qڱ(���l{�V/��*�;~��=�K�ه:���ƶ�����P��s�0,���Cj�+����9ƻ]�����|g�ayˏ>��
~�����'G�ZO4΁O2�X��h�ب#	R����0���"S
�8*ڙ�W��#A��1��Sz�=�k~_s�:Ca��8�z=x�\��r������+�Ra���e)cr�1ۡ�>����?�G�S�~�{�88��ڲl���g�s��3d��n8���#�l�/���� ~��%�p1:113�<�|�C����Z�9+EP��q�~GFǓ;Q s��T��T�ZGY\a�F
f��}���K94��I4U���&d%��n�[ŷB�2j�%���&���i�Mdi��8W�P>�Hr��i �E��S�\�VV�?,ā��X��|)��눬����i��O�,��Lz�w�����Ұ�'ǲU�ﴯ�K�4��@!>�x�w�D@#9.�nx������h��b�y�a���q��2���(��?�ձ�g�׹���%�=��
e-��Z[���#�aO|Tzu���y�=7�өq�KTv=�>���RRˏ��Hr'!�dnk�И�U.��+qX��C���V�i{����} �`fK�����i{b33 �\�0'�*+���Nl���;ǅM[�"��?���;/���V�\E �a�T����Ƹ�A�6֔������$9�i�����"M�m��3|��H�/戋�;#�Eڿ4��W�Jx��[���n�Ձ���|�^?���~d�O�.M�	/�'���9���}�����4��z�s�%yLD ��A�v�҇�;��'�R��7vy�/ݢ�.X���J�4�IJ�9MA�ɷ�R�A,^�,�N-����>�����MOl
-�?��&M����`�����h#4w����!iX �f��)��Ƞ��$�u�����gץJ�"s^��F����X��i�(��X�}hg�TFQ\SS�_�����))��J�h�Eϛ�EDY��;i�H���ڙ#���P;���<]_B�%�σ�T,2ٲ�#Z�D�<���I��_&}�%�^��Ű:��O�����t}a���y�$�K�<��T��e!��&���o����ºZb���E����b9�`Q��Mc8�V��s�u���m]��$_3��g }tucY��ڽ���.��9��A���3�Hu S?���˺m͖��S*n ����I꼐R��W�zy;dNWϲ]�-�׻���5j@񩰂|�+�vL�C��UuW���.�a����,+Ы�C���1V�����a�l`y��Zia�4cM۸�gb��pj:��QJ��^�@��Wee���3^�
"�rݘ�>�d�L�瑯�	N_�E�� �� B�ɵA��m��JMik�A����J�>D{�B�20f�#� �Y:@2M������!0�P�HAc_��5�B[~��&xY���z.�CO3�����U[���_p6�f�^�b~u����/��Cw�Ƀf���`��IL����!%�N�؞��7��TR �r�|��M{�]��\W�"�� {���%R�|�[`_��)��U7�7�K�Qa]�ɹ�Ɂz��a�S=�Jǧ�}A8�J�f܅`�2<�����XN�8Yv�	�t����s��~�J��qz�w�y��k�*�fH"�P"v�M�7��m "��n�Cƺ�ۢ)�TΝ�����is���&2R�^��_:�Bm
j��I.�!���L=�k�z�{�G���/ ,*�<�)%~��G��2$Ti=��qy���`Ե	.`�g��(̃H�()�B
T
���}�����/�ݍ�@��폠W$�6!��L���2�M�o}H��
0�E`M
,�=�pv}od�x�Nݯ�9cC/)K�W/�Q�ËQ��5��˕�RD}�h�6��\�務O�+�\Vr$����PJ�t|$1uy5�~c��W��V�~��f���@5�ڗ� 7����,��]� TMM��;r���^U��ID1s
��ш�e�=_r�Z�i�T�%'7n��m^�)ۤC#��Aw|�������"Z1��c�m��o7���	�\�j��ơg�"��(tD;^����$s5�7̉��F�J8�ҥo�S��>AA=9��˨.��KW9]1x�<	8�T^�O���n�B���m�B/pEj`�0J]�{�7�/b�o>$��<�Z?$��~�-z�0�L�+X����&�"� H�Z�y��l��
L��G<x�s ��Ҵ���Ӯ����4�e	}X.�ɺ����T��j�0$�	!1.�t꛶"ԯ$2+�C۴�#1�� ��� O�'��GdD�;?vw��E���K�p>���#�ܩ �~�D�s�Q1k�9�E �#x{	��{t�{,���{pl��WK��b�Po�@v�g,�&F$�Y>��(��u�Rf����?��g1k#��ZDsiĦ4�k}�9������C R�ّy�J�m ��BQY��߇ ]�-���`/���]x�4�ڜ��`�YŻ0����t�W��H����SPg�ܐc��T� ��:�&�=p/b�;�W��w�_X�?7����d�x�L�c|���˯F^�f�;���#,���2�G�C�ڳ/�jh�5�C_�WuN��`��ߺ0�p��=e�*S9Wg�*GJp��jS�0=��&�_�]dΪ ���lx��6٘b��x�(٘��	=�)�+����
p�
7�f�C:h'��~���0 �K�u�\�qg���4CB+��'ǔd�Ne�����N^���0�6E�rS�v���WKZL<�ޙKI��%�Rc�?�0����_ύ�<�:�}��ɹ�K�<�h0g���?�Hg��QwZA��&�\o�k�����ԶZ�V���蔯<���ɴ8I�^�����yh.=EM��J�tYϻgR_a�sVM ��
>ՉI0�Xk�����e�>:��h}?�� d����Qx�sH�q������z:�A��>���O�$4�d
F4��;���)��A8�l؝�*ag4��P(��V�,�o���x���w�x�ӷ62G���A�O�JbK.��"��R�(y@�A��p ��� ؍���yN�jO���*@_�~N
�j&���_�q�ނw�4i��9Oe���7E��A��t��KtF�:�0�8^g�!*_&�����,v,�	=2+;�b�~s"�S��~0B;#�������礚��Kԃ���;K�t�i���`.~T�h�|���ky���d����z���,\��J�9�jux�8i����t��g����k%v�l���Γ�>�t1������s{�C@!�K�3/c89�g{�����	��^'t���!u�%�t�b�6"u{��B@n��˄i��gK��_h
�-�o�+���"��֕�'h#���K� waƻj�"_���fgn�l�L��\�p���n���^3�B�oo��>���	�1�����	~��09s��,�2i����b��T_��i��g��>M4��1�Y���gC�£�8���sV;h���F�='+٦�A�`T������GCC�ӰG�ֆ�c*~Foס�:~v��6�[�/͍�,r��a!a, 5��,2[ę2�jM��	o�YtN@�X�$=r������V#0���*�&M�꛰S����P'��h�a�%*X
�a�i"�rV����KY������J�Y��M8����c�[�[��$�c���`���X��UI�5m�U�8E���l���ϣz�bn�%��l�?ҋ>dլV&K�m� �?�7�}�|�Vd���5�q��}5���#F���R��!:A��GB�O\\��ǝ '�qg��f�(��$��P�X�S{B�Y�+3�}����u9���eo��$�[�p�u6ň$.��(���l<9�-D��38_��3��~�=6@���}��QC�T���+��������%��x�{�	c�n��)�i���K�y�d���|�b�{���/�jg%,��Ɓ	`��`z�=�@&E%!G�#�0L�W�Ӝ�����J;n\���V�2
�&ƻ7��h��|vzi]��������E婁��� �؄�;����-B��K���}0} ܾ���jz�Ê��a;8[6�:��K[��n(s*�Rn�=i9HO`D�7X��-ޢ&����*�U�)�A,0�#L{��/���1ZJŐ�B�jt\�1[nJ��|u�ԋB�B����!f�z����� R�o�40"�OO�=� Q��V�eɏ�,���M	'9a���Ѕ��kd�G/�,i;��}#SH��߆��V�\$<�	R�ޣ��:��H̘�����-Y`6���
q���}Q�9���%����r�ȼ�[ �	u�	6��<_d9!��y𛟻��.S����6'��.o����J�3T����lRg���ʠ&�o%��c�X�0�y��G�a5�����Cam���c��-j��M��K1WL	1čz��r�a-���!0P�߱�vZ����ǝ,��x�w�V�r�h�<�a�l�����z�߮�!�7��7~3W�hy���=|T&&�Kl"��_u�.��A�+&3u�=�2#~��	j�x~��uc��r��' ���8`�E�&,̸����R&�<���¬��C�����·Xd�Pd����:0Ȳ�����%�Du�m��kMr��笠&�ϋ�~`QA���������/���k��@���@É�п'i�95������+�-=����yLى<�Yew(�Lw�G�Se�\����Fm߾�.G��cNAM�2D/憟t�HH����c`
T�Y�7l��6�p5s��Ցx�YwȒR��`����:n�(]@�<*Rjs�fۙ�GD�"�7�}��KS�2Q��
�˒VO��i���V��Q >A�Ch�'��y@V`�nF����c��0ѵ�)z���|�>Z3����O��q`�,��
�-�S�N�Y��2_*����]8\��f]���:E:���`�!�?�4�ѱA��Ӽ`@2zuBǠFZ-�	3!�U*�c�tGW_�E�͢��k��4����__YһЭ7)�e�]�C��h�3�m@�D�	��ɫ���ib�x,��
aʒ |`|9�@l����O��I����C'ıaھ|5B
�i��\;���Zuq_�&�͊�� �Z�J��4���:�z��_�������t��h�l\�1,	��f��#J^�P��V�2}��L�	~��f����S�b0�W��O�b^k"'�u�f��^����?�m\T��
���������C��GqL��*��Z&e��]�c�x蕵ؔ�R�1��F�U���!Q�M}N��g;�p�˖]�X)U^��fu��(���4�H#��Bҍ��_(B���Sz��0�#."�9#K �)V�&Z�&zپhW�х<�??v��<�9��?�5�{ϊxc���d:P�/� ���y u?B�i�⤜J�ȃ=VVx�O����'v'���b/�����R�?pf��;y���t��%��Fk)Cq�B<l��m�S@7��NV�M#@��n]��ȤeG_u��j�	����4�*:D�N��u�h!��[a���悸}ѽ�J��2�k�v�3�{ϯi��t2�d�3m�n�F~�Z='9̂ѷ��'��߸2e��e
�����=^������Ϭo_��a���bx�<d#Y�����F�p=��k�K�v��@�%);Ucw���-��t�F�u�����S�u"?�j�v
s>��DXg痢R3����I/f熌ҷ?�_����,� ���KP51K�j�2�CI?�ɰ�wG�0�'4[b��	dڪ
������<��|����v�g46Nϝ����F���(�V�fR�CT5c:���*K�E����Vx�����xLk#�Ú�,��Z킃��Ʈ�ŉ h���5�?N���#!�hY �{���]���yܼ��Ef�C�.S*�fRݘs<!Z��}�MT�ѡ�N����]P��'��fP\��w�����~��C�kp��u-O��tmȩh� @pf�]r����@tB��6=sİU&�O�;C�-����S���%�>*-��8M������@�� /���7���q����2�Iu9�����`^��CV'� JK[���'�?��A�]��.A��q$�t���f����IZ.���wD?��U��Z'��xL��n3 ���7�lo������+�gyT��.�8���d=ح�w^�Nc7�a��-�P� K,�'�)x��ֲ�>^ptq��z�@H�{_Q�f}�:�UQ"R���.u�����~d�͑m3��Kz6AaKd�����Ѩ�t����~�^m��W�h�
�V���l�"�Q�nP1�;\��p������O�����i��j�������xn�<S-F��M�h��^��u��>sfÅB�|0�B�Ku�
F��#��(���̢7��/�~IR2XH��2�ł�u��h���,O�N�2:D+��4��row�s�?Q[��o�0�V
��� a+�&� g��ݺ�LAO�����D}�pL~���ú��!�[!�Ԥ����E��=��~��.��)�}���)�t��@0_`�%��R���PP=�O�@�>��r��L�;2˭]K;�@�ك�Ȝ8tw�ű���v���,&�C_��b�;e�W���y�S6 }H7B��ʈ�7-��˂�47�.e4��˕~��|ZKG�����h�Of�gĩQ/2�K�?����W_��������c��a��@R�ZF�H�-U� g<^��� m
���=�����M�����zf�̘�;j滓I�3k�`�p�z,^D/KH��N��wIh'Ww�*}���k�k�7n9B�>��!�<:X�nV~x�v�]�S@.�t�/���9����6�(��t�Pz�4D�x��F��)�\v$�9�4�e�f_�grw��r��2�ʹ5J	�է����B?������ ���jÇ4?.Z��_�{��f;HE�j�D��j���� �Øa�^/�`Fo 1J�n��0>-t8��_�>9 ��#���:�0��W������<rg��`&��LN�X�ԁ�}�C,ԣ�d��f�w�!u{e�Xk�;�����jNT�e0�p/ڈ�	�˷Cipq�q��l�0�����.�O�e6���A����kK�w��8�j���Ì����%7���t�Ghj����D#A����Ib���a�Y5uY�o�t ,s۾�K�>�5� �D)�����ɳw=��c�Q�`#9��X"�j�%�s��9�el��]~�t������j�8s�S�)*���,�L���=�k�(���w��ɲ�D�.�DF��]�HY�{�5S�T�pKZ���h�ʧ�6�#�P��l�p�C;���P��Vo���j]]��pl���H��_c�����d�91q˽��_|�7P����%����Wb�-�%�����U �:m��r�����bs�V��(~�a���w�t	j{���&d��������3*X:�*Q�vb��^`rNX)��u0�a4*��e���$\0"|h�]���Ztư6�ɰ � ���X�kw;r:d�OOfV���h$��E#���$^2��0����N�yn�W�����w2P�,��涁�)!AT�|�_���@O|��_G��7W~	���"(-�8���<�Z���žc^�v��B��&���,�]���6���n+@~L� v�����+�!�0�+���	�J%i.b�~-	�(p�n�f�c����y���^aN��(���#�^^E�P�-,=�)M�M�cc*J�?K�y3B���yi&Mj̾\.D/�`2��α��j�e?P�A����	�M���m��v!���TK|��X@b���ˡ�&]�Ѐ<YM a;=Z��-̣(����a��ayo���v��~Vt����D�Ѻ�(R6�۽5�V�i75���.&`R��
��.��YD6�X-ݘ>mxcl�ϹA��a'��]y�K��3��	��}+l�8x-�o�aD"�ç"���5c�sHWU�/9��c����){h��{� ��V��n�P��HvZ��Ix$��,�@<o�τ.�$%��!]�/(&g�c�*g�_	�xE�u���;����0W6�-�$���(�Iâ ظ�0Q��1I���Ʋ1�8pb�-ʬ��o����1�྾�����	K���M��e�ﳺxk��~/����)���`b�.�P%4�S�2i�rt#N�ڶ�BL�C�o��s�\�k4��Y�k��ܩ�B14B�������$��Zc�'�j�����Vօ�(ӼH��o�2����i�A�=ZO��^a3�h7�e�7�^���L����"�T z��I�pfL.��임�l�-Pf��O�J�R��A��9(���8��MfJ7��©�}/]�2�t?�g1�B�F�%ypL �q�s#����֢�X��cu���ۋf���*����si8��v�*50d��fE��is�*O������D����$/��Ř˿C�Z3"��F_�(����?+�����]�~���"H��v�R;��������cY�F��G���J������k'(t�� T�[gᕚ�e�[����,_�I�?BPPmi�(d-���E�mmF+�)� })��|��u�K^L��k���2��߄�^q�;�*���q!��q̉R����
��B6/���?�HJ�e��76.�m�E��:9�Z����t?0 �w���	����'U݊���@i�<f����c��`%{>�-�a07R�4�e�K.�w��׾�z{YuT8�\��W�-E�&�2r�-���!�y<q��H�Xo�'�\B�86^N� *\)øo2�m�t��)$ƽ���j�̒w츯�YQP�(�:V�_B��q�$+6�͐�_��"���#:�����#�_�!�>d��"
�H�������[Z����x�L�f����ѧJ4�K>S��Ĭ�E��28e?����#��Գ���.�T��cE3��ğ���Z����cq��J�p�iOs��y�~�"f	��!��w�{n �� �l�-��2@;��f�{�����8�P�+�ށ���.�D҂���t.j�) �$(c_%m<��Ia\3+'Rl;^������C�C��g�����B���6��#�f�[��AQf{�nAh�͛s�%v^G�>	|8�	l`�μ"ˮ��Dr����M���/Cr{z%���}Dy.�����]�Rϱ_�z{LݨU��BVN�{��v���qH@����a<ӽo/	���}���3�`���[.�\I	!ř
���?� �TD%�f��i����fY�3���:1B�~GҸ��� ��om���N>=r$,z�Į�"�~%5������BL���m	��_�
1\���83��|�ѥ>���q�
QY��LK�]��&c6�6ψ�����GR�$=7K�oZ����������+ʹ, 2J�?4̮ۈ�Z)o��[++�-PU���bT�I�tʤ4M}�S�<0,�H�q��ݫL� �G � 6��+���&�'��g��M��Ș���+z�h�_��O�-��"���7��>s�"�SjN�!�@ϝG�2.0خA	��WC������:��/$�.6aIT��oS|-:^�j�I�SV�ԯD�����K-����(���33�.)˴9u����_��\IC�<7L���i<���0���(f[���y܍��Nn��{��S��D��B�i��h\ؾEh�����Nddj=�_��@�nq�BH&�m��L} z��g�D��"�rm��oO���z(в�T����#*jv7
���(B�Uh�L ^��Z��!9�t��DE$1�4�2��	A����s".I^ڇ�K�i>��ӻTR@�N�j=���a�D�M�Œ�B2(���:͠�6�h
VZ.��:L���Wcr�"���=�q2�(�����v!�2��=��h�p�� ��7���h�9����t��ϑ!.��}4׎�m��� ���o��@���NE�z;���J�}�~s��V�͆�Gs,�΄����ͣ�,�R|�^��?��*W���5~�|�ە�xJ�Gd���������2}7�>ӓ7�o�/_��.��V��d�?�(��ܹ���\�.y1�f�(���`�g^��$��"���,*t��H��C1mT(҂�yZ����Aa�x-u8Wt��k�^�hG
&��0����x[v�����Ẁ�So��%�J҅L���6p �-_*9"�Cu�]��4��K6�7��� ޸��>�PR~�K���p+�����aE������>��F���\x�q�������U1hF ����*�_|6���n#{����!���}���8����n��O�B��������R�Kh"���X�r வ��6^z���6)�c s���V������{.����L�.�Lj<D�86���z:��?�3D\��T��]�L8�z��os#wp{89ʴP�_P�:�G���)
�_�Q�ݷ��d
��GD���$Nt	��_n��R*6������ѝDv�������v���%2�ݫQ�u�2��ġ2�-R�f��{=��T�g�4�J9	��c�0i�����bZ���s3xh'Xc�`.W.b�1��~�! Z��AT8�?����{�E����ؕ��z.�	(V����M��9��\f���� 6�RN2tr'{�+�_y3��6�I�܄�.�r��=��A��J���b��,���,�Mo���B�i�XA��q���bLT�pvB��PsO�S&��`lhǪv���[�ցTv9�i"�ò�	�������ڬ�~J�h(�@4��s!9�3�����	 T����u�2���t�������9���^1|�'���2�R�G�u+�����%R��Ag`�ѓ1�������I�#mXt!񯆱K��hc��/��T����������G|_��pz97b�&K�#|�˲Jbg%�+*���qF�4m?�N��ĄT$��NG�3���H2����=Mi���*�C2��}:`Tjk�~��7�F=�|$Vt|�r���m��O�x\����1�����?$�}��E�o�0��af#��.�ء)D�ξ��G��T	
߅\B���j��J������#¯���+]~6�L���Z�@��IYT.p�����s�&���/�R�����U!���ξ6I����}i��_����i;V5�ZD�kb]q������y(R���7��jk��Y�ݓZgg��y�T^��JB��O	�.>�Q�P8�R��'ө�v��!�.���N2��m9<�v��m2�:�1%_�P�D��<jw��*յ�=�8��3P��=�Q�g��q6pf�3O�C�{�´t��*>x �.S`��������uɲa?�]�x��w��6�mԣ�����d���?5B/Z�� ��K��@鞔G���)TLU��x_3��R��*���d ��v0���C��}؛X#K�Hm<�!� �����7o��4�襇Ҳ�ڜ�|dr��2b�zt�ق�p%PI����:z+���^ �M��g���T"fΑzG�͌ajF�x<��y*MQhM��Y���	��t��"�6E)��م�p*�ǥ���[m�欑g�ĠH%'�Y�Y��E�z݃BIZ�M'�!K&�JD������D��"�KpI����)M~�B0��C��%~C���e2f'�=0!&���������O��[�������zv�)d^�b�,8�U����;��:�����3�?b"��C��e�o�nN�g��4�:�8A�i����͹K}`Z��������!v�Aj�x�����>|�KM/��h�"��_����*�~��)U$�L��sW���۝;�#�����̬�7 a>�\�_R��Cƫ�{�#�Dz��`D�MSCV����f�f~������.a	��n}�1�M+%�8R�����y�Y}�����-�o�K�m�D�����'�.R��	�5	/$B��pY
z��#d�Wq_�ߖs .��!��0Nq��D�^��m7��rq3R�����[����̴��el�ա�#�0�W�5�x��׫�ѿ������"�+�$�,�<�*�"��e��,��{lCm����=�"ʆx�G�cܡ�8ZuX�M|1��!'ĠyR��~U�ɩ�0�S״l�G�]+"���ݛ��T�wy�ru豶��_ l��sDH��S��W���@EGn?��emp�"T�=���1>�oP�[4���>�9�	�>	��J�(;��V�r�PR�@�1^4�_���?(�����`n}���Q������|r���X�蹯�r�k�3����h�^���~�&�i�f�sBtk�{G:Iw�5;�ω[����p��<;U�5D�w$
VG�pڊQ���jЅ��)�G����G�>T�a�2*�� 7%0��K��uVE�b��{�ֲ�+��HX�xs��X}t���@Rũ��=����ҲY�3�TK=�B�
������-�Ֆ�G�"/��=�l�6	������^��m���ɶ�h�����*5�T��O�a���l�F��a�ɐzY`(FVF����	y;N�p��u��ߡ��Ȓ�"��[Dci7�8Gx�D�z��,5g;����QwQIz�g���0�V���s⽥R.4�-��,ʜ�X\�wP� ���+�=�}�m��$�
�f	)�->�M��R�9nL)�.�3h��M��(E����B��}�� ­�P#H��br�e%����.�%� B	ئŲj����w`WF�3�|g"w����s���l�T� Jt��(���^)�'
�H������0���R��K1�W
|E�ޠ]Mv�M�j�0��4b��m�����&��=�ӌr0J	��\[���
#BO)�%9�&]�1]��e���3S3~��㲑d,E�T��܈]ʖ�댗��JDwu��t���������J��JT��0������ظVÍ�֔=)���[����⬹��S+d#�@=S����$���Y�}b�|���jM�|�1�1����������)s�%�o��
f�D�f������v��Ӗ��.k-!-(}�� o+%��l�~[�M�t�fPEG�c�.��2�jf�+m������2)��L����_��]�����66�x)%�a	�� ��T%xC�l�Zu��~Y�'<�Q�������q�KJ̈ڱ�=��zߺ�B�A/<��:�[sXv#����ճX�i-�8�3)�o� F�3b����V�P>p���4�Z�y��>8����t�8g���-���}#��3"p�{b�<X��x�_�:����ci�^KV�Ts�_�����l��U��N�<�^�SQ D�ȁ�n�)]�X�(|�ƞ�� ���M�x����c9;Q���*�==�˚�7�Kq0�>�-U=e��i�SW�1�]e�Wa�[qS
�8!Ɖ^!&ޞ�y,��a��p�j�[�����S��� Fc^^��6�լ��˶m��M�Ya��pG�8h+��{M�1��e�,���D�:� !lL7~�p̾$,�5�iw�?�qY���ޱ�x�x��ğ��]QW�� �؞����3b��/T��CEi�x+V5>�:�p[���J�VD��˔n�"���R���>�=���b'�Z�?��Wמ�x�r�mV ���|900��,�	i)���b����-[�T� ��S!k�vG�������m���8��"�@=�!�8aI�8�^��&���ߐ���քXNc�I#&z��\�%��<4f�����s��%��7%��]m�*[���[�{w�5�>�)��ac�R�tL
��E�������8>����q�� ��@`0�X��幱�rp������Y�rP$��D��F��Z
%�6ۚtͩ9o����E/-0���/>��oͶ��{��˙��wu��u�Y����Γa�Sc��<5�'���aZ�-J��Nm��X����.A�Cn*��;��2�)��p�J$R{$<d�3^+�<�c�n�o�
��)��;��0�E��n�rY2��-�h_I:}�Iѷ�x8Qi��֞	ol��ư�hA�$����L���@e��z$�ǰK�f�9*�ؐ�.��o��p���L��X�fI�C�~2�>#B1l�͔1߃�5�,���,�1Y�;6�w��oȃr����ɹ���Ϳ<��| ���c-P�� Q�-�6���@�r�V2ˆ�!Qz�ع�ezɭ6Y��uV��a���ͷ�}Lj�ɨ��)�xE��^�s���+	/JE��-CȔC����h�+���{����sF�d�^��J�P(8|5��,�`����Us�A|�Ez�DtF[��W���J�wk���*F�(�虈��:Ҍ�O�M�G��Nx�jҌd�K���N����j���f�6�%�������|�F�� �7���-���A�6�̋�u/A��@����:�Z�aw^���,��]��K���c|�<`�n���ǆ��4cw��������L��-�h��q
�1F��I�6pm��f���x:0��	-oW�O��Di��EԜ?�s��{eW��W��&
�V���_7��,l��5U�w��%x���!qZ`<�����`�Z����LD�Y������M˶�_!��v�������	~1��o�#��0�y��b�m�IW-���A��q��}��l�vAÈ"Cl�8��@�����^<=��=E(_���������e�@���@�[
C��L05b�� [�ϝY���&���A����w|�K��/���A`�Pc�m�s��q���̘��c=��`���[�mD����;!��4�*���*�?��O3x�mq[#Z�UMuy�������#ȍ�L��h&��t�¢�x�~�GT�jS�m��[@Ɓ�pC��r}׸	���Ч�ѽ7}��i�	�.q|�@���>��$#�<�^�&��V��)�u�U�{DYc�
��:�g�=A�:-���M����B<t)+�H�r�|�s��Х�)���鈁ݬu2`A���~"��sNB$A���G	)�eiof�E4f�CN�ҙ�@ӝѭ`���"�]�JIi�6qR�`�(�	)��c:��{�ऀ���	���ݬ<��Eu����(���m.cI=��͏�V�)0�����'���%4c���ڔ��Ų:Z�כ�W���DO�T.�'����26H@��Zow#�Ę#/��9)��j����p�Aq�@"�k��#U:-���O�<��R��%��Z�ϧ⹝mr�����i��s��r�6rw��HHY]���se���0���A.=6�J���㼬M2c�1tm9���	���S�q:F>D�[��,��SW��t��*������O[�(��N�֖r�H�p8c5H,rчT�=�����������xҁ>tc�>��1���؁��>�iL�	��/��Y\f���Aʁ�}ꫝ<�V����0g"�8Aw��E`���jgM��ڐ�85PINL�["[A!w�$ µ� ��2	c�$ �ȃc\���N�����
R��/mɛ�k2�em��o�J��,A�X:7����s
]�v)����x�<#���^���G0�#'H�T^�$L��Y��z�Z�F��t%����؜���󩺻�U���^����k%8<oXi]7��w�( �k�1����K��M�z�/�`��Qw5s�?����N��K���$��ո7��A������}�=�8y��������]*�S%j%�~�	Y��11Yтy�@�Tr�T��7_Q�x#mܛ.�ƃ���������ȉaiݥ��_޼b8�n$���Բ��OM��Q���{��W��l?q\��͖�׿��?�"	�8u�ܳ_5ሧ>AXE��5`�/
���bu�(@{�ГnH��>���� �8�~�΃ۇ'����T��n���L�$!S�QP�q:�4s��i`	�; ��z�\b�wB��Mub���u���?Z�����l�͠JX���zs�[PJ��,��Qw��:cxA�:�sN�v&J��i�,��8aմ@7������FUUv����dN�g�xZ��.���h �i{u��x>*`O ���4���2�X8����(��W,�RW�c���d��/���#9pJ���Ȯ��s'����X1��y�2�*�.�� 's�?&e������798f�#])�N^����~S��al�I�oj�0�F<�N���oxA	�ٶ9j@�ƕ��+�8�x\L�$N>8rѥX،��?��8A�0���͈����xj�4nց��̉���YTK��*C~�Sj��'Rji6���#��ZOu$���v��P��G^�:OP�e��T�l���k�v��pL�e�%^A
�%j���C\�~�
ele�b�<>��C��6��P���Ź�,�/�x+����k�
� ����~b�H���0q;1t2����W��G>����_]J�!���H����ߛ�}�Z��iZ
��=+M�m�w�=-u1�9�kx�+ �ŧ�K+Ĉ`إ
��/0�-��MCRII���tF:��S�(�5�{��W{ŝ�q硂�P�F�IIX���h�b 2�*���F�Wʶ}�2%��Q0�����C׾,[t�׮��P0T̋k��Qocr�2�~�����oC~=�؀҆��{��I��J_����S7�[I/}�:�M����#�����)�B�qL9��q����j\K/e�s0����#�����~N�ףK�ڰo����σne�)�ݩ���z�\��y_K)��J���˵��~��P7osʗ�|���=����)�=M:O�?A=m -kul�:۴h�w��DAEh}�߀�U�^1���ɀ~����c�NF��gX6٭�_���p�i\͗�{3�f�Zf�k��t:c�>���
L�x���t��7E�B�'�ʉf	jKP1y�K������8�uo���#S\u���� C"Y �nݗ���#_�v��9�G����B �����S>�Hxj�K�r�2���34����B�_�Дm�D�Q�b Fw�SQ�5�{d�%kULF�8����0�K���L��Zh"�*&�_�݈��n?y�����5,hŔ=DgNݐb�u;H���ظ񹺛o�i��E'm��G�;NH�z�q	&��Ov��Pq ��X����ٸ��Q���3b��S乤|ͅ�]����jV)��>H�4`�q��l���n�����L�ˢۂ5Ua���ac~Md=��c�9Ǖ!F�� ��������9x���uz��}���c����O���,}V�D�J$�D�tI���fZ��7t{c]V�R)�B#�.���@�Z�)�U�ʔ��UKm��3Zy��g��3�^��ă�.*9�H8S�������*:?$��c����L��>�P�:�H(�-P��c��4[�O�k��)W$���������F��dqn1��i��=�q��52�$��uW"M'*��G6p�˵���F�Y�������>HY����3�nV��D����ۄ/ĺ��ī��~$�MO�	��\���(���ރa�p�n(-�������avk+��b5�'-�t�E�g#XG�}���l��І3cK`�z�C]s�sN����V�<|�F6ܣ�#�#���0~�EzE���Z-��BZNGe��[�՛F|F�k��[�������	~WU��w��s�O�-�X ��w�I�a���{r'���*�|
�˫60�Wf�y�Fh�M�H�t�j�T}k"G��@m�6"���žBs�,��Y׀��_�QD �7����/��ҍo�uJ�a\E$w�\���z��@>�%u���U�`�: ���8Do�2�F}KuMD$k�F�`�c��\�lD�B��������H���Π��ѓ������Y|�a�_��Na�0�-������t�˶�� �*��\��4��G�.7�����54G$�g��PN���Ŕ0����XA1h���}p��dqy��4�i�qK���A5ݣ��pXr��78�ЊK��(çj�E�0�']*~i�.���A�@�
�0��;Y�����G7I��.#�6� 0��X�/����d�C� 9��/S�Ȳ9�u���v	)D:f~�Ӷ3���2E�6��V�B��t�|෉�H�}q��,�	�����;�8���^oM����D-�6g?�q�2�,c�`��噒��t��V�G������ ����È�qC�iM��cJu�[� 9>��9ҡL�!�����tl�J�v39(E�ؚ����o�e��K���r��ɎD�#�	��͖tvɳ�oL�L���^3clߏ�$����nX�~`4V{��K��ȳyT'��GQsms溪4�eQ=ݺ����UOK"i@��U[�sVb��c��
�>�8 u�2�dr;?4bh��Qz�Y�=�2�>�Hs9��6�'�O`�#6�.Q�����/�sY�@�i#����G�FԚ�p���e�,�:��?}�;��U�̳�E�y�q�����j��q�$ݖK,<�������QX"����?��-�b]�f����7�#�.��P<h�u�����uH>�X<#^��c�O��ɢX���Z��o��k0j:���q���2Z�-�B�%cM�t��� �T#����ju|�o������cT�����uj2���S�=�>�WTK?� �g�W2/��C9��hP|��Yvǳ��s�mdTc���?DU$v�F��|}x���5�ɥ�T��1��<,r~!?�C�Ax�U���Xf'��D7�H0��?p�����Sg��'���R*)i8W�
P���o�$D)XoE��v���h�<���L(7�tZ�o:�O{J7+&��~3Q/����ͻ
˹���py�
�S1�5�����+��/b���:���˰s������EG	Bb��͊-��@�i�yiuІN�ܫ_+���RQX̄�!"��-��qG0���S���Ԅ����[���.h-�+A.�܉V��I
��  ���js9�swsR�.w�ć�� '����t}�=�u��勣x�����`��<M�L�f?�#��z���� �jT6��9Tt4T�" �W�Ƒ�GϩpԕT݁��rޜ����
8x���v=��4�*M�6P*�P�v܍	=��/Uc�%���$���`b��ڮ�w��G� �0����9�[��&�����a����|������Q�R[�r���a�Q����������]����~��VQ�)ռ<�$�����eoU+SM��p��c��j	TУ�%�l��i~��fo�1�5�0	E;��r��A	�6H|}8i#,V��&{�����4�O�˪o4�����z��nTc����]�}	��4)��c��FAs+�R�	[�|�6�}��R��i��ӣzO�1A�D�(���ʃ��-��� ��]�S�Aa��"v%��� r�Ccl ��0�Y��n��`�����g�@��O��(�uw0�,3�~���~�b�,�dtVF��������>���,�����3g� �k�*%*����~��.�hR�������jb y?������'�2�
�di!s�o�w�?p;�P����Q����z5=�g��h��U���2��Z�{k�6n8l�M�~8�b�L)sW��L��7fń���|r��tL;h^�����U�c���6Sc��
�w<"0�O�}/ &J`��܀�Y~|J9L��5�rcD9r��2�8�.bG��B%=8l;`�ˉ�`o�46K
��poe=Is�η��'�l�9�.�(���������W��OEM�,�C��Fœ(a�僕��Z,_$˂:��]M�y!8Jre�^����&�;���*�<��v����A�+Dq#B(0���A�Bė���mt�Ut>)N)�=y�?6|+���>�d��CUA�޷�;c÷���DU?6���\�i�u���F��l,R���F�J��.L�t��{�.��aD��~yx��;$f���1ˣ1��Ih�uJ���Θ��a�#�8������c�ہC g��A�"�,�4�c��}�'2#%؋��c/����폜v�{��s�;��=HBhKˌ�v���4�6�gϭډ��E�7�!"Gw%<�NI���z���(a4#T��|-�f����юF�?�0���
��ڕ%�x���\Jш���%�C,��%Ʋ�6Nȴ?��6�`�c��{�q�d3+\���-���4�������`�Ҡy��w�#l�3d�M���7�i�\;"�C�tzq��u��fa[��֎��x�h�VYȣ1�b�@3����KK�h�^�-��Gr� Ӳ�Zݸ�/dE�1���$;���e4������v�z����Q���'O-|`��02Աh����r5�]^�h�e�r�w���y{�LV�=������>Bkx�|��7Er�!:AC�lj���Fі���?�S�w?�~�)#Kr@P����F�n��9����zM�!fu��=�f�|a\��6u{L��/[���R$�����(�#��g��S$�u�?/'m-�J�������luܷ����b!�X�W���#R�t팁&��4o��LY-$���N���d�J�f�pu1 �ZH������O�ߧ=�
h�!�c�;�;ߚ��/P!\��ER�[��IY�z������������~u������<J��hO�ۣ�Q;�V��)�k>�W'
]�}�bE��fD�7��E,�Y�[�i&v��R�ޮH�3�2v0�y���q�>K����M�3e�P�6��K)��3L#6��X2o�?�4��.�~�ͪ��"�r��b��ۚu(���f��Ŕ�w� �v9cVCŃ���4I=��X��|�M�Pn|L8�"i����o���̣�����ܽ���Ȕr�F ie¢�� �
�Ӑ�G^^�E���ݑ��6��t��P{ܓ�;,^��Z!�|�K��T%[3y�����{=D�a߀�}�gҷ<�d���dƂt����C�r�<�']�#�H~�o�w7ZG�T����:֚D�V+"=R��*��9y��M9/�!u�L�4G�)ͬ�H|�x���*��S��`�x������ f�A�@��cYqY7�dyUV@<�S��~8��䊶}"7�ҶeY
�˷Dd��G�:J�h�e��L���a�s�u@˯o�x��ʣ\T��W	�\����<����)�{��b���l9��� ��t�"θ��!����+swL;���r`�TL+���t/���(s7�n$U���@S���c��,��/S|����� �	w��6�ű\O:������:���C���O�@I��@s��]���&� �ߓ]$eQ��h�N�E����8ga@*�<��Cg���5�s��vڶ@�=vZ��yM}��+���@����针����r
sU��w��W ��G#����qH���y�Y� �Wz�\�^Jǝ�p�D����o�6�Q��_��YIF?ϐuXF��;3u�CG�ϟ�Lx	�A�7i8j1:EN���J�Yt�O�Gw�۫O�����O7��jd����_������,E2�JBg��D�4��OX�����EP�󼓣"�(T 7�k�V���P�.M���2^�Y�W��SÍ�`�(�\W[g�:t�|�rX�0�th����ɱ�'Fp��{� sb����5&��x:�p�2�d��7K��0����RU�Ea|�6������N<0��@�A�:�ݥ�tL�����s� Y�w�89�jOyA�I���ˠ�Qy
qrN�a X�p^7�)@Y1��`������3�QN��xtGA.Q�phy�b*`��F|�]� 6�����	�_
�Lƪ�,Τ�إ���xrg��'�d3��6�e����U�J��y�OvdT�.���|	�Υۇg`���}�Kz@m�B��Oeᶰ���@p��dʦ�;��H&Q_R���҈ �4s(�!����mK ��J��E��bV4�gJ&��^��]A�9��j2ռ֤��GƝ�z9X;�Ejv������Q��uo�=��� ��\c�E��.�!C�����}mҋ�L@�X'��j}1ب��1�H��L�����H�b�W�_���
CŊ�۲�h.�E-O>�?{���2 ��ыT�,�#�~91|�툠`�PD���\Re��պ��Ύ����J<V�mz�d���e��u�w�!�⁧2׼+�/{aV��H����mδ��R�@��!���)=۾�%�)�e��a����~tw[$�yp���݂����2�OƸ;�n�O�O�y��#msq�y�-��UmP��@A�K0��"��;?�w�i!$z=x�F�����Ē�uf�����F�w�^�n_��Ô,�
�\���.P�ӿ|����x�rV��" r�'��X�u��b6�ϸ��˃z����U�?���T¶��1��Aَۢ� �<�e-W
�&�,}�����t���{Ø�m�7e@����c��*hd���֨V�zR�)�8��)�8��U�}(b$��^�k�gO%r"UT��k���W��*�ֆzU ��Ʃ�Ռ$e�[�!K������'䚖P5��+��lj�Ly~X^Q�,��r�>k����#�7����~||s|��\�'jPX�Z%�S̞1$����Ņ8$	����υ����i{�<�	�h(��_�S������.'A�*꿿_p"!һr�/a��q��]���|M���:�9��a��:�w��`�]��
�ƭ�N:�勷� G�qG<m�O�INa��[�Â���������'9�֮�)(�z�j DҮr{y���l��>�Ķ��	ʀ�^�A���+�g�]���&��'&@��%�H��TTn���$�|1q�K�aƄ���inT�<d @}ɄeUM8@��dP\D��ߍd@�/e��Þvp�ff�&��E��.�8_���sY��龹�ߩ7���+���޽R��(��?�S\�p�=�ZΙљ�X��v&�`��������X��N@K�h�Qn_�.�2:��à�`��b�]��.D5�N��޳rrh֤�>[�ܔ��IMphb�/p#�� ����O�nl�Xq�jz�ٿ�4<��՚��9���C3_Ϳ����n�YL��Y&#>�	X,�Ѧuj�����?��2 �]�M��t�yd��N^�1�P�>��z#O"�ll5�M����T.�7'��**�YÑ�ߙ<c@����)`�2$&K���~�i5�vea�<FE��eڟ��ڤ&��G��#�y!��G1���c^�) ����,�a��Ɠo[�z�]}�EWx�!��T��Z?��$DN�R'����ؖ���.�����\�Yu��v㏹�*�.��0�?��3ʶ��2��%Ǽ�t�}#�m�+N��b2u��X��/�=���en���У���������Q��>��(
IBH�͓tw����m��<*'�<(T�Ck�JwLʐo�5��h�Q�+�
��Q����\1Tu���4��]���' ��vb���1�N�+�K&�;ճ��5�s*
�o����<'�y%�6zX���ē%Z�3��=����y�e�M-w���u�����&�E^<Aر:�$;{R�ҫ�H��ݖ����_��9I�5�bGu��"k	x�[�U�+Vx��[��[b�C������vg|�J�1+����\U�{�x�^p�7�K�b|rs9H���=X��k�"@�K�P*����o$P���ΟWD��.��D	e6�I�H�k�e��·���W�cF�9�^r���Q�7s�됍c��Y���\�{�g�;���s�T)�Fu'�x�� :V'�T*3]Ѷ�G)�O5��v��(���[��{pDsɮ���gW���pV2`D��@,�TLi�nʚ$3���E�I���ҪZIQDmJ$�{��|�]����+֭"C&w#V���X���wڳ�oJ�N줾t}����F)��!���D&X�@h�1{U��
Emi�mv�r�.�����&��u��TuKj�w1q�S(�!2�'�?�E��C�m�B^],�{��/u���b��{���|�B㬹�o�� b���{rT���m��t��a���J[KOg��'�I��/KՒ�ʹUO��L���;�A���)�SF%5�rr�:&b�r�e���<���TU���ǈ��k?`�I�;C&�Kb���m<���2>3���*c��5v��U߳W��&�gVҐ� b�TV�U����t?a��+��y*|(�.kz�H���0� L�sw^�}���ՔY!�*��ʫ���a���w�ߺ�U6)��[�B���ki�q![�:Y�#&����5�V�Ղ�v\
WJ�%󃿙|1�}��=� 8Kw@;���i-��f��i��f�	�T��vi)f�A��>(��d�����ݤ9���_�,�g}�/Ϳ�V� �}>+Ȥ{�Z1��&�)鿞�(=C#a�h�ר�PHa�'hdۗi�`o�~�=,����xL;�;�(w�j�.p�n���TCk0�W��`�g�CL�;��51�(?A4����Õ�+�8�/T�3���C(�"o7ƘBi�N��t��!b�pB��1����ܛ\�V'���"��2����Ov���&-�E� �W�ih�5�,�+@�s3װ�}lb�	(��M{2dl�~��QQ 7ƴ�E�3����t���2�;��Js��&~�A�r�Ρ�J(���� �I3�^C֔<_�+���e<!&�f���6%���X�U�EZ3^3�G˷�����j�/����/M��O��:.�L�31P��P������6�!���2��;RmS��y�el�46�m�x*�t�s�|���dΐlb7z0�S��Uq"�i�-��`%�7n�R{	�:G �E��u"��g�d�}��BVѳ����u\��T����v%��ra�d[?�J=g:�ҲID%�����4��f�^�MCQ��B����H��y���-�2��.D�4��������y8��kI�#ΞՓ�	�4lU�w�ϊ�4ZiI
���~iϔH��ࣝ�\C�䶐�뷙��tA	������W9'�f�2��׎�y_�X����]}׭�GJ$�aĿm$W�vo$(Ғ[������]K!S�;T'=�K������8P�$!QYX��-ӛ3�L��X��cλ}�'3��R��#�c�pG�z��5k�"a�܂ۗ��gw���>�u�I?|t`�U�7�� ~pia�W�E� ��qTs�}��b��^4���Ԟ�AA���ɂ�C�	$QV\��Y!�>�df��(�f��#I�7DK���f4�T\gPi)+�b��i�I���zR4��T)_��\�������0دꍩ��ߙ��|��7�~ 7,�Ow7���G���k���j����-p���PPK�\	x���	+�|GP�5���[���O����GczVy}_�*���m2���k��0�߯z���E��x��ڣ��9NÜ��P]�<m�������SJ�/ꬱ\������^D%�
�@ݞ��;ytvaYS�Q�i�h�����������%Q��n�Rp'��_�L���H�wh��a"")�au�b�8���!i�υMy��U%Ϥ;+�n6�!�!��}� �s�����%��Q��V��"W%�ݫv���K�N��^.6���L�"�?�a	�jU�%0Cc���z���l)�T0��/�sް���
9M5��S-�M�����L)vf������9��s�H
#ٱ��=̳'�m��D4�
|�j��W�Q?�E,Ni_%ۙAq��:?��L�r�<��sR��\s�(�]"��]?C:�6o8��_>�f
ǋ��ѷ\Z$�h��\IRZEd�i�>��=#ul��T6��6.6bL����1�� �Փ��<^��fAiwk�xJ�tǴ�
�m�h��f��u���R���Q������G��iR�a�k�l[����J���-c���	����Z4����[p.z��>D
zu��B���IF��:�����q�"��]f����հG?�n����,P��#���_�[�Z��wWSU���<�;�*ޝ����J$�$�� Tq���|�#���Yh,�=a��d�1��v�#�l��fu��˓���g�#K*��I �ed}�=q>��cB�����4��A9���3+.U�[��`O��� B!݇,_u�����{VƜq)>�Z���|�^:�3Q6d�
����6VR�5������>��C�7�󬫰�H��DG�*(���nM���t�<�+����N�Z��.�t#�^��d<OB~�Qʘ\϶ł'�kD�]	wI+'T��}�^�{ ��!�-�U���3t~��Ilsp�:�!�KhN�+�]��aU��:�HZ�؅��{��PfF�A��S�NC(��{R���ߧ Xl��&JRT;�׺ǰXժu�&l�J"F�O���:��s�~�����hRu)5������p����?DGh�tr:�z�o:�r+�vڬ(&[�'jtvL��J��#����q��22IR��l�ʨ^]Q�[�TC��LOo� ��pd���˃ш��X\��e*HX6�g��+�ƣ��05e��f�|�^���jMÎ��[ݖ�V7�B����z�o�@��1b�p��["´� �M�"�ܳ��TkWSëʻ�6���
��h�A��`@~h�}رk8

����]�ǁ��U��YS�:�J�
$\��K_�zb�S'����'B㙜��4�m��p���~�ŏZt�ν��N費���9
sjO~�l����H#�o<��Z��ΰS�8�u��xK���\˦�J]F�������8q�P���^�wЏD�kn�Z|/k�O��B�R���õN/��"�q:W�	�ՍZ�0vf2V��8}J$��^��6�J�!�l��]`"1�� ��?�~V'r�j��Ƀ��V�x�Ku�՗z���eq�^�l�����˲�8�O��%y��{P���,�i<c���d��# ��1m�ݠ]O���7�@Aō��.GH��W��+��-���j'�K7��5q�S�n;�G������P�'Qej���1Dd�AP.�G���3�Qd?��,�J�����O4C燁���>����{�q��1��f��/q�I�G���?��\�.�X���B��H��.*zտ4�9�������ߋ����cF�P�����RC�3$�{���=�SF����]��W.J=��Qi�8'�V_he$���>|@G��M<���I�@��3����|A/�j^��C�[��:�]<Y���R��5̘�1����JU�6��9�;�M�io���e�X˭4#�$�!N s�H�˒T1�;��P���@����;�+'~���j��~��w{�Ӯ�us�!Lk^,&'�<H��/��JгS0s���ҁ��z{�4�YN�*_൉�N�-I���4$�n�Zp�a�Y�����"Xh��>��z���Y�^�8��l��Ro�]d�.Osjx���W�ȼ/ډ��)TIn��y���s�9����d�6�ߖ �����TE�.����2���P۝�t%Q�(Gĥ��5�����ϑ�ӳ7Y��T��X¿T��㎔<��[	A�&��9d5�~�x�����R��)�4�XL�8�U��ox���ڶ��	���ۚV���3E����{߰[t׻�֏���QI4���IsM\�B�~$59 �����d��{M�N"rցs	M�-00fE��xn<�i6������8/[@�f�e���Ч�������{�u"*�S�8.���K�]������-�E�#�̒M0C���d��y�* z@��F[����l�!C���&+�C-?�2{��S�j[�LxG<�g�'˭�j�2�Z�6�J���km\�Eց�"�G�͍P׽�^�G����i�J	�����!I>�n�W��9��� ���%��}�x����v�9)�#��8�@�'j�ܘx�.�h�۳���?ڦ�����wѸ��UI6C)b��i���Ya���m��X֡m?!�����3
W
L�10t�KF�}R�je�?�5���^�%[�<m�#�M ���GJ@���i�0�N�z�Ԉ]�G��A|�#y�l�z/4�R&�r6�JĤ�8\�j��\3P�i~��?0���ޓ���M9�o��f��w��c�Ε|h.&L���Mu��b�)ݕi\N�6ك%�8�����De��o�U{�k' ���� �[�/�;��H�sI���D0ګT��s C��=%�l_�b�5 �A�� p����S�������S�!�?jbtY"�Q<���VQ$�k��D�M�Y�����Vɱ�5�5�ؘ�)��jW�b�i�z�
l������KYu���}��0)"&�Z����'R�jrL�����.*/�e����]�R�e(,,ztLk-s�d"*V�ܥ[G���[�k���{}�}x��2%x��NkZL��A��UV�2�Tq�N�m��~o��҉�ҞW;3<j��j��9!�Rr�p��B��w>�@���y쒱$3'��������>��)h����\�/:��K�������1�j�?^9���ЧC���+Xe��j�+��}Cp5 �����D�RZ3}��?�f�ïs��o���pV3�/���3���ݔ�mf���xt��ۜw&��"��G���%	�2�t��a�%��B�����A���K�����Rol���	3GGg5};�?�U"X&3�Pn� O�4����l7�.~1��`m������(�٦����-8"�_���}뺬�T�^�`.�?Z0dC/���n�B�Lf�ihʸ`i5}
���O!�N��a��8U�N@��v�:�<�pS�>=�0S�h��(l��6u])=t	]|��#(���8�;���Vy+�#n��RG����+TN!�$'��n���6�
��;l����}��M�e�����tJp���.ˣ4mD��\�=�̴	ĵC�n���"�EhN��s�=
ׄH?����1^�	�,�s�60;)�����d�:����,�61�{O�S3�,Q� �i��jeB��f>����=?3��Lw&_�����۟�=c\N���_-�gk)����� eq��2R�(��.��P.��{pu�mֱ��y����?x��Kf? �t�>��3f����s��.e˱�������Yʼ����Z*��#�A�W��$9�߭�ٮ�Y�����(�M�1�o�<p}��n�֢?�����j�*Q'�"��5�iB@���Ϙ�Vt\�[ï��X�&8�a��X�&,M	U���^����x��22�^mV�&�*4�� _>��2�@E������GϘg�sq)��i�����C,6hP\K�H�C��9��*.o)��r�����rY�CS�׎[�q�jbe�U�?��zA��88-y�(�iJ�nm}S��V�i$�;2ݳXd�{�@�XD�דC̡��y�g���
Ĵ����cHm�kW��.\Mya,.��^b۞�K��9��qp�~�V@ E��~=Str�l<�|� ��:�޴2�A���z7WU��"�T\u�X��=�̿}��K�M���ϐhO�G�-�'����}աn��Gh�8K0�����Å ���}|���/D��l׉�m5L���u� B���ґ�<�\��J�ʸN�?Hbb���0c�.�qJ��zQ�`����>f�v�K:�\[���#������{ثd���� ֮['.��;�y�P/,eW�A9�G�(zg+`ۥ���/<���^�q[��2%xy�˓�� �4��LS
�z؂��	bZ2o^�$��p�C���Ba�5X�`Z%|q��^i��_Q�)?U`0�IL-vw�����H�~��'�d˦T|���|�x`��k���%g#�̧�FQ�F�;�?����~��J�,7A��� dw9�x"����p��3q��ubeu_��O5&'�5���A��q�����.+�`Y(1d����-V��D���`�����n��(ITad��A�k����Y�:'���gu�H��N��3�uf��m7��
<4���/��G0�6�-�J���[�1^B�[Gsp ���S��"oh3��b7�ӫ����2.E�Bv��#�U<U�A&$u=�C�,��g�<8��d`��d�ev�qь0?�J�qI����5*_^�ɥ������)��1�#)`�c6��;��KD��8y��}��s��ޅ1C�d�u�.zi]�A���H�JϏ�F���xZsWAu��ٙiFVY�uZ��D��K�{'t ~h\�v��V+�Fmx�l��iB�����l��4�!Y ��eT8ߕ��J��-@��y���B����*ѝ��7��wz�X�T6�^c�~Jj�t�xj������&�J�]k65�R�����̺�_t�E$��ٮJ�Qע�)B8=���;��.�U)�3�҆�J�Z���Ew4	���lՁ7�j�I�(7<��	�o�%��ju(��#�O�&����@W{��F���ׄO��Y?���+��(�?�� ɳ0���
��m�E�7=�"�Kjב���Ƶ���b����עj���d��f�&Z�Hב_N�J��~��tE�����
����nY��ހGf�f��[�p��EÍ{��be>P@P�m��1�e�a����D�ūҦ������|<� #��S:(�Bӏ��#i�?�`7#�:�a��ӟ�H{�|����l���R��x������0�/W��z� ��'�$�	1���/E�Z�P(K�y��}�~5�5���莨�*��	0҃|��_��LS���j!U��n+<�>����e����P�h�g���S�{���ބ����jYڲ�.]5.����r���w�d￬v<'�aϧD�V�lV����Ԁ��&o�j�ZD���?ɛ�(`|���g��Y�� 1��[w��e2�V���v����هt�h��<L#*��y�Bg\�T����XT�։�H�E��}�,���׭�Wd�m��w�T��*;� �%l��3�!W�6���o4�v����@��L�&�l�c{@�|���s[c�dR��<���ex�ֳ�6�~(������.��G����nO��G�T�C�J��Aϭq�	l�pm�)��AU�EX�aS� �)����jە�5�%.(=�9썸�em�P�}	p63j�zQ���l�n��"��i�'��G��{���J�h���|��������*��w �[��}��)��당�� �a���F㫰�a1G�Ht���9�q�����²�E��*�P�1B��V���T���rk��Wڈ�L�:����}��{�9��M�u�/��(Zg�ґ?�8��1�$֐�1f=�z�d�[�Kޱ=fBʕ��ؼ���	�~zi���6��1ǰo,����3F�W��oB�G����J���e�8�3����F��Ȏ���I���Y|i4�k�y��H�YU�cQCZ�W��+Q�$TL #���6x?�1�ׯ kd�f>����Ve�ZU`���Y��>I�e¡U�<�G���Ж�.l��s.9�����?	��P����=�VAǈ^6<�]���FH���]�^�v�pچS�W�`B=��؟v��-��J2y����dw!ښ��0k^)�!���tz��EHN�-#�|��g�!�k<;F�/��`�a,�����m��uR�����[X �l9f��m�L��
f]��	�.�^��&VN6!�?/��<C�r����EB9��=�j���p�<.��ci&���ŉ�e�f���S7bX/��cd��YL�Q�M)������n�Gi��P�E��9�="tߒ$b���P��I���P��V�k
�3�Nr���Mͩi��V�Ǿ���E����jH��XF����D#��ԟ�V_j�"k?�S\�۝�=#T���	|��_|u �@��_�����)$��/:}�!����p/�1�Z$|�������=h,<��Ķ5T|c�Xt�Lm�m[�ǎ�`6�>?��;�k]����[noj���CIV`���1fMF�Є���z���{�	D&���1+���������9�%v���4)q��.f-����K�0%�<�r��?���T�?X�l�h�Ĵ�iq���cL/�U&�	U�
`� ,�;L���sc�s�Ea����_�k�l���H�蕍�Ŷ�_ �e�@!}�v�t$����悸}R���>"�\[�(�P��F5o�k('�/�tēkA
-氫�	o!�k�>8D5~�
P����&��y�r�$^�3חM����>�����w,�]=Q���f���C6.xz(l،�!}�3����{^�\��2֣��rj&�Ϯ�f�QgӃ�~x|\�+�~ AM�n\!��8mH9�V��@�� @��۶�qcs$;��/�+S�q�u1�2 �_�! aq�NE��Wx�z�4d����i���E��0��?O��Ѥ�$���ԣ�-�,���u��R�F�l`�s�(�s|l��q����F��w�����y�ń{~�/�Φ��Iw�C���D�̵��� ��ʟQ�����M���Vp9�	OnQ^76ͭqo��)E�	��^�0��0	\��}�I	xv��'>�̫��#�C�-��,#� }���tcm�+�4��mo�7d�K>���y褩��e��OV�%����^9&�R�_�;L
��S %m�y�?��s7�������ޢ�rXQ�HWj�<*A���|������M�D��8����sca٤��g�^�R��1�xݾ8�|�8E"���,�K�_��&S�͝V%Ț�<w��<fݨT%d�x���|�x���$9Ǐ�Zn���+�r��J�0� ȭߌ��vM���@`�N�&|��s�Pe[�8�b�pGkв`���U!�#��(����s�b��9���Ʃ��:��6!j}Z%���Sd�z7�PoO���E��n~t���M�]y���vQ�)肰�� �୍��k�*yƜ�;>q���`�۠ԡ�I+wm������Aϧ�m5Ú���B�)����ii��K�u�[L����wL0�*É���V�)A�!�6�������΅p^4\~џ�?��~�}��YZ��Y5�G��|����3v8y7#^�A���v�1-lଟ|&F�Ab�^�Ɇ����N�R^h�g�0�ԑ�o58B��,�tea8�0�~J����`�E֖R�����s��z����K�h�B������O^%�I+x�]�
�P��a(h�[���(�)�*��UP �0�c��m��{����޺�~��;�����5�B��-�o�K�peAޱ�4߾BH{}"���r	]0��ss���"�Eg�JY�>�� 4ǯ�}r`����oL����>JU#�.���Y;p��Z/ynH	3P���4���U3e#�d�F�B`r�������p�֙�ђe|ߖKl��vˋ!
%�<���a��Z�t3GC�̢�W39۫�)��c���V�Om�]8�D��=���j-K�������J�!��_�ST�\Y\��V���_+o�r�1&����^�L�r�ͩ���I-?�s����}���t0���������!�D�f�j4V��X��nʼj�5@�W�_f�¼��*�4Y��H��H�V,oQE$��a74]+���}$.�����Ъ)>1�'��^� ����Q�Qo]�G!�d�U�����u��4��茟��1Fg���T)��A#�T�%12J][�kjuJ����"�����W:-'�)�u�l�%�F�L�p�a��<���J�E=�D��W��m�_4TLaB�b���';�O�YU��5N8(��4�,�R�z/���̬�,��f
�ݐ��~�f��4	�;�������"�y�p3¤�`�Ž�m�X6wZ�n�W�q�
]�-����_�-���X7NTQ��c8�#cČ�>���MY�Ზ�����Uɥ�P�с��\	կ�ʉ���Ü�����#/)]gp��t�7X���.١����2��Z38U@�����"��zK�!1�6�I}ͽ��ϋxGq��^�Q��a�����6�4qy��f~|�G�̉�[B������+����Gp��6�5���o��לhI�3��L�}v�t7�z�Ig��r��΃��m�=���!c����1BJ)��}�Ƌ�Y5�X��j�	y�se��a	*��+"V����L��bs_(���p��8/�
�wf�����$&�I<዁��o�J�i��[�����4� ����ˎ"f����;�����USuV�)�~M
�h9��D�	$��F��
7�V�����x����W_U+��ſ0
 ���4�t�s-�bWIL)��a�8,��_��*�IO�l�%���\<L�6�~���˓�p�M��i͏Y������KKf��o��S���(����I|(Xas�C�K�U���E���L�AA�}h+�;�Կ�t�9�a���.������+�q%��A�0�`M�RQ�ҥ�z))#�Y!�N�G��bqQ�|Ti�6ߢ�!b�F���ġ�Uv�2��잏ҕ�Y����x2sS��՞�W`��]��ˮ�r՟8ͫF� �.����m�!\ ۑ�Z��"�o����%��� ��Z��@���$�N�)���7 �Q:>j3�� O�g�X��7h����2Lu��웵�Z 2�I��͝~��M�˂��-���d7^�}H,�}m^�����V�� ���pc!�Q�N6�L�ϔ2����s�j%��{�U@�~ʿ�9Tp�M�X�e٠k�"|T5mx��� 
��OB
nRslGBE�'��\ѕ���Y�����~�{藹��GS)J��r�E��55%!�H'R�v+1sA{�T(vtR�؟��n��$Q�>H��]�>���[���6���P�O�u2K�u���q��r�Y�K[��3 ���S������w�A��>2���;9����ݡF�#��žo;l�����Vp�~8v���SMbaÔ�Jf�����d�NI�O�[jV��CȤz�6������:�R$_�EC�?���/�ަ�{	���m�S;�����k�~�C�n\z���HV�e�|�^A��z
�hd�{e)F[��}��:�b�����
9�����ҶW�#I�T�r�=%��%�� Y�"�l�EG ��)#Ν��r��ڸ�L�+��%�g`28�"8�%��F,uF�X�q���ی�ﮁ���B���+��CϏ���U��l��.�a҉3�d4���Ap��D~ڋY��}���_HB:�w-��g�lW3�H؅��lK�g_���ަ�Ȝ���q�RI�m�;\%��j���+���t�S������V�������;�B��ܽ����sh#RD�1wQmdB�� �>�?���%���[q�\~Av����W��x���y�L�[���]D��6�p���7,N�~0�P��7�b(V����dʏǇ�vG��C�C�,���J��\�d���ġqE��ĝ�7?	��p�b��d���Tg�0�TAJ�^(7Z!�=\�b�ဇP�oq��mg�����S��Ж ���xWH��$�/AO<��e=��h?Q���)s-:dׅ?�������=���g�Qx�`�'��\YTzc��8�ȳ�T�G	2��e��({��	g�X�uP�t8�AE�s�vy����	
��;�e�k��V�WB��*������&eͫ]�����R>F�5!�ˆ���R�S��Q���]�xm㎱���|~����%m��!�L��2%��Awo�I ���W�K�,�{#�x~xS��?�*E����=��/|@�\7U_��JlЫ�@��J��Ǜ������h0O����,l�d-�������A�i/��Ǫ�E�����Л4;Ҳ��i��1oècGpy��A�y}�:~�|��A���V���^�3�@eE?^�P�nBs8j]� ��7�\V���
����˔��(���OhK�o��p�M6���dXc���wчO���m�e*�F���֪g��%]�1��!|�8����.�h������Iۘq+=������~�w��6 ��M9�Ɂ��at>������̹ƣTv!f�.%N�L}�q��4�F�?�]QwOk*�R�w�#�v�+���(����j3�Ӭ<*5~�i������Zk���L����4l�q��3O��9��`���o��]�&���� �Jo,�P��C���Ä�1�(��t�*��P��0����3���E�D�g{ۿ!J)'����Vy��
��4��"^�9���G^��t�/��+N�K�~��?��IzI�x�u���� �~p/|D��M� %�y��K���La <�7��P'�V �o�i�Tt�%5��KX��a����a��+6msx'���9����eطI��;",��B��S�"���wꏿ�E��n0�"D5�r �w��S3E�0��*�.N�G�����Iw�Di©c�u=�N�2�8-ha��
�G�UE�Fa���BTv�A����zOB���u�g��������!9�0�=z ���p)k+-r��?%�N<�^�L���v�>��ul���i���'2{b�dp���S`/M�)��?�V��S�����x0u}��QI�,�b:Uz�E�L%�z�lK{/;�����L��*��2���|����5^�� � ��so˺��]M[Bܽ� ���Ȝ>@F�D��_ecA�~Z7h���_r�chmU�2v�������5\�+?��Ԕ�>�ON�^6�HC��uj�����s���y�yo��s<�o�����a�m�@�u�����By0��U^A�|C�:�\�!�.������&�����bl�n��e ��sK&��o�ƹ>[��:�qP5��Cw���*ߕ�َ�}G �l�Ժ���eF-�ђ����e��Ht[־���2*P�Q��kKH<?�
?P���pq�q0���*�z/�2Pw�V$�`#B�S��&(;��BV6O�$$�Wc��Fj*Z����hF$�|�n�@=,Z��@-zͧہ9EGT���}:$:]W����~����G�c�������;�����K�!�ͽ�r������� X���&�kO=X�`������E���)�xCᛖst�P\1]$�KO�^,<zە}�e�9�:m�<��z01��Yus���l_}��i����0bZ�#�@8ԟc~w�3�L�}��ϙd�����3̔�Č^�&�Z~v�N�����a4���IjK*�ޗ�����Х�e�q��)�9���Ym��<�u��˨w�
��:Y�Tw����������2<Y�� I)y&IX�#b�I�w~�������YW��J�)�H��<,l�/����h�O��m82q��n(̅F*DTh����J�J'�ɻB�?q�i����5��2z�2 ��>�נ��Q�m� �=�>ʸa%�>Jf��A�̎c�����E!<&�!QIg�k���T�}��ftQ\�����r�hc�����A��P��!Ϭ���9�+3�I���Z�"�<s�����ZC�r�ķ�U%5�R�����ܷ�|�A(B��d;�>0���u�E�a��n�zi�}xϖ��펱��m��6������7���h�5W|��!��a�N@!�+��?�z�e,ԯ�D���QE[Y����~���������ޯ��A�k�$(��S� ���*��f��.���{_��[�vA�8����X5�!DX1���	�z����&ߏ8K j�,x��>���{+ڵ�Sk�`I'�;K8�]l�����]P@=�c7�y-�9��.��b����$��p2~�C�Y/���������q/00��'�1�ҩ/"�N���2�N�=I+i΂�*ć�ߥ��֊"0*�s��z�	��׬:H2�m��N`��z�v-K�з- �tdwM�����co��v.���Q^W�����r$nH�G4�MN�����`��������!F���k<q4��-�n}�g�rMI��ʌ"H˲b'�wh��=�JY���G��b���(��U�K�-_��y����tz�JW��.�u\���D(*���
�
6}w��[�b�*��=�̃����כ�5�{v��}��TH>ܢ8��1O;�Z�;ѐٚ�=]LeR� ��¢7��W�J����ۅ q3E� ty�0r�lc|jyn5�.��-aJ$s}՝�-WdF�$#Hg>)G�ؚ�_Z8]�a�
�x 
j�!�"�f�Ė+�3�sŽ@4�u\CY�f%��������o�a�#I�	�����R�oWw���%l�$}d*�H�t�zDiexL방�r�夕�%�ŷY�<�6 0���>��H�H��a�ʝX�{1.�A�:�l~��P���;ñRӠl�lq�'Ы�� 6��"�<z���P9F��a�t���mZ�(ԝ�%g4݌s4c@}q~|S�| ���tK���r�I[�W�x���*�vl�V�j� �/�@~���H�@�"����=��]����|��*���Q������gm�h1���g.��뻽�?�TϤ�|�c�9�V%��fX�%�1���w��@�����>F��Rh�X����Ձ�䜷1�5����>��b�!6�x�o��� ��Oa�m��m��_�!�J`�[v��l�#��qN�EYƸ�}[�价	�:��,٬M�8B꯼����$ƳApE��{�bG��(�#L9 f-7�%�\����{�N�;(�*�!����V��׼��k���5�h����y�01���C��0�6۫5.�Q��0ojqٮB/j�ų���#'��6�M���$X���$	����RL�/~����qb����O�v�&e"#�/���Em��1���0ގ�Խ�[ü�����^��Gl�Y��ɊO��?M��Q1x*s�A���]��e���JW Yet�<G|�O
����G��IO�&2�!l��
�˒]�׎k�W;�)0BM[>7�2s�\�n���:(JϋZp$)G��E"`��R��gek�==�`��:����iYF!���T��Tu�:!���������P�<D�l����4��Dk?�wFM�W.o�3�>�^[�3��x	=܌�Ύ���56oj�4~�S$9�T�oBd֊���ZM'������GI�,��\`<ǕH!�I6�kgqPGQ=VZGڧ��v!+D�����.E�PQ� E���Tba\�o��/4��܂sӀ!��pR�7��K#.z�t�H�c,��<���X:ު7�Kb���!P����:��\�W���M��.~p.Ӆ��х��iSd�����AV<d ��`�δH��lF�!-�}
�ܳ՗tŉ8��B鏋g>4�ѕ��r���1y������&�C�` ڄo��v����v�D�_[�I��X'�ۜC��%��S �/)쵸`�-�3Ca�D��Ii���=5^q���t�E������v�@9���w�U|�g����_���6�߹H�!�hܗk�_ y��J}�=��6���0%�� 4�PYf�(}RT�J����`_�
�5N�/�~�G"�>#Q=���Fs�>�ao8��dB�4v����ZW�el�9GP�ĳT~���+���$�����7_�Bz��r���/h���<�qO#"��eذ��a��EK���Ч��,�L�|���~�{��\vr9�~���@Ս�l���l�0�Q��J���*3�������)i#}v�.�U,/��:�\��:�'Ĺ�zw�u��*�����wNv�!�y���X�H�W�L'q��A��0�6��YW�"~:W����p�e���@Hy�x�8�4_��dͮ/2g��x�82�ڻ�46 8�$ц7}�~5�W�����kW0r`yڄG����ٺ�c�nM�Ӭ��=I�B�:K����U��ȟ��N����vD�m��%�V?�����N�_1����yW7���.kc�1h��/_E�L|��@�B]�n�;����w9�s����[ �@��,�3�2@꭬��:�J����]Pq���T�QG�@8��X����M��ǡ����А4���������xU�\����L�]��/k3��/P���w�E�b]�S�͏!�MB�/�y�q�C(q>��:��d�ڰc8�ũ{���mtÝ���7����&���\<ۯ�8ǲm8��Q���C��,I�>j������2��iϗy�2� z2Ykq�V�����᳉7��_/AI��̩�Α
���	��G�W�s���]��4h��k�� py.��b]��P3q�i��y�H*x4���tc���cgJ/����m�g3ZN^S#]kmL*p��'A��w�l[�4�c�:�z[I�G�D�#J���g�P}.�����y<M�Zֆ�\S�9Y�-R}s����*����ũhU��B#wi�ٴ�^d��('�+AoJ���@8k\��N��푕���k�<���ZR8���#��a͕��)z5�R�4%&7�B��< ahHUa�Ӓ����	-�N��ywy���vׂ���Ȃ�;g=KL��˿��k�yz�Vd.��I�-��	���vQEڵ��S\yNؠ"Y��Қ�X6�g.h��3�%����):����Qw.a!��L�
�е`���Ǟ�z���6Q��vǈ��-�R��;]�ʟ�{�S��tr����̚M-$O��-A���]��$��M
U���m��[���)�h@���`��x4�x��q�z\�L["�3B1o���	gΙԈ�tQ��P*~��1ٿ��ҥ�d�`�٦?�9e�Uh}�a�R�&a���'w�B$2���c�gV��ta�Qi$ד.jXN�ꢜaJ��@��S1CE��N"X�%��D_s�YBp��f[P<,��?��F��x"��h�,[ZJ]k�ĵ�� ��v.���G�N��
@nS���I�x"�����X��*�FEEk�!	FV�b�=W�<�Zz�m%�х��`�U�^�����,=>
%�3��r5��~�����4�v�� R�U��!R�P@ ~��n�x�_Xx�#U��'�߱�e���7k���������I��[oX�����B�;��5x� ��(�$��|��AI����lT�2�:EחQ�\�M��ŀ�C�s��fN���i\~�P��l�V9��}XВ��ڐC�ʁtl��9Q�ǯT��D�9��nn�^U
f?^`�ZK�EA�>�	5���Ȭ�����x��&4���j{�*�t0�7�TWLm0 _��t�|\�����-a����1	�m��j���JJ!�
��R�/Z3J�xJvv��=�C	nfS�]ݴ#����_�݄�����Q�N�%�}���/��msGZ��Ʌ�g&����<��k8�	+Y=}���4�B�S��2O�K58���4Q���BnG�2c��#���Wu!Y�c%��}��"�}�R����_Y2����'�,-��fB���&��]��+���C�j�>L���,���oԀQ�Ai/6#a 9z�3������Tx-�k{T[�u��3z>>�Z���_�/A�������	� �ں���̀o	�je��1�W����9]�tgP�����o���������{��u:�C�(��Ⱦ�/`?y��G��,��"�Q`4D,' ��(��멄۹x�����_���H��V���'��Z�Wqi�46I]�@��e��Q�<��\���ɿ<gd��N�8��F��v� (�E��u�M�1��K������Ɂ��tMlX�#:8NX�hE֧_FUmNpPL����a�0｜�2��}��U>�	9�]wz�9� h<D�»9�gf�@;,�=atO�t�~���T� �J�G�(B����a�����xTZGp��Ba�u�����®��l��/R���p�sr�N��@G�6.-��C�^�3f���.�����T�
�H��S5����I1]ś���3"�[����X�c ���󫤏�Y(��˻W�i�P�B+�J%V��%�����c���2i�� ��E���G����i���qr�>o���{.r�]�g@��8m���{v"o�6�6�k@ٛ�d�F��$���c8�|I�q@x�ۚ�<ha[�[L�0ʹ��)3�ZpGAQ]S�0l��'HN���;+$VK"�D����E ���+QD���=G��rabw�9�@7(<��;�t�ή�9��₮�X�Sx�̍�t�^#Q��L�5��	��i';�^��\ja�����f�"�s�1��6���M����(Y. �۝o�c�5��L�	�bn�����3��5���O�K�����˙q���a����味r�Ɋv��`��CR�^;G���0Ep���R�P�7u�|��"d�>ԠB)�9|-�yx{�ܺbQ��#E'�/�e5X�.2t��Y��1��v_b�|c�RSwG���w����r�D�a�HK�~cK���a�:�-T�)Ŋ,r��lK��m7�XB��\e��-�b�c�_ �o(H���u0��m���1%��KG���Z�yTYk�ٳ�^�,z5[���؈A�e