XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��!˼�K �*���!���ϰ���<A��3�-�Rv������^�;c�l*��J�r��;e]V���y��bgmh`��r_	�TU��F��H{��{' �M֔�B
!�����曷[nsn��.%��s��\#�>����hE�^)v�ì�ĥ;��Z�����sN�I�����tF^>!T�ǫ)R�mA�nE{Q��ԉ��Hɢ?1(�0'�g��V�H�A{3mߟ�iW�2� �n�gՈLR����!F��oB�s;I*,_.���^/2S���#���a=}p����^J�16�_�+�׬����t�����O���:�����!�Q���6,�N�.�vPu3 韰2����gۚK��a������7:%����$Nq޼��a+�X�3gf�kJ� -���PJ�K���-m���:�'��4Y'y�z��|�3��4\� ���l����GD�(@X����ȏ�B.:1~Нj�˻����w#�X�rB���+����`G�p����}	&��[U��TQ��3&�J�U@C��A�=1�my��tK���	#��fWI.lR��>0��Ǻ�^���$�3`����[9����~Z�S���([����G_���M����/�J\*�z�ج�<�pE=�fP�,�M�&I��X�A�ϟk�o�I�(̷oIJFĕRգA��S��p��"d�����|���@$�>/���3��V�������Q���$D�	]�4��'gB.T���}p���-6v���XlxVHYEB     400     1c0�
\�%�	�ELHwY\L�ahے��8��b�J�1�!k��{|׮�D`Ep˱;"I��K���g��!����^A7�eW�TI��K	�{`���b�����i�|�e�۹�.9+V�V}�&j6~�~s��"� Q��e�Wk/�h���u�c��j'F���*3�c�C�dd:�*7h���:
Whݯ�n��@��9���"O�P��P~�U�>+�G�"�o�G��3j\@.k*���o�"a�P
m�Z�O�0�T��w� �=���n��t��^5����D�N����-���W��O����u7��˃b F�]1b��6�~�C�"�Q��ބ�]i����_s�'�A�ʂ��]]X�%�'Y<��9�D� U>-�=��}�5)e8��V��C��gX�gi@��y����og�1j~�.�<��fXlxVHYEB     400     150�M|Y�b)�'9T��g�Y�?xd�ף���88���<�8#W8[VS|�ֲ��$�C���y�5fk�v�
a��-f�7&T�y���=��
�ٲ)�F������,_������W;���5��(U�g�!�@�y�W'�l�j'���i_ZR�#��
m�-�	�O+y�6nݪB����it��[r��L%�-�cb[���P��Y� g�tͷ�8��z��[�'�,��@/`�"++���������*�.vK�)��5�p1��N�|�z��%CQQB��������8���3j�����:�3 �0r�V�:N?~������|�T���(�����XlxVHYEB     400     130a�u �����KF'*p3�)�b0+��Zq%}z��K�R��mT L!y���6�2�Ě��Ru���?ګӽ�O�HX	���]g����p�����9���-]�?H�פ��,�8]���E�=�G��Y������:�'9��iYd����ןL4�\�
���?�Źݷ��ZA���=+ؚJ��]�
	�o�|G�A�	��j��"�ߛ�GK¸�o�������A�Q��t�J�(���*ld@��'�V6R�"�r��l�A�(8�֚��@㏽�5 ���Qxx?̝TAt��!m��f~�q��|XlxVHYEB     400     160��l��:Q(̮l�����ϲ\E�?�ȴx���6|4Fp��z��8�_�|E�rѩڦ2�C#R=��|
H�a��ԯ��@���=`��)Bٶ?��V�UUP�T��4�|�*�m%�p� ��	>)%GVb�[[�z��Ip��]�s����=��}�j⯓��� �&�s�~����H�ݺ5��t}�����uz����|�����v��>�bNJ-�.�"�g��M��Ժ�z�̓��M46���/gdߡ���rYH�&j(>�>����3�3K1 ����H{��,{�+my<����#>U�g-��V�Y�߫�iv�C��N��˻T��z�lW�l��7,�XlxVHYEB     400     1e0�Q�7wR`��OPH$�x�]�q�wn��SA�d��g ����o��N=6st��;N��6�������o�K}�_�M�,*Gu�#f�)�I@�sR���p�}��W>��(�:Z���Ph �;�*;�0>�H� �:c�c�/cǾ���ܷ9�4� U�잮�!D֬APdV]���k���;ن�R�ɂ��%I�"���g�0B��,/��̫+82+���*&��\p�TQr�8K߼��M���ߧ���*���O���
�G�wN�(D�L0��2���p��G�VR�+B��ȎF�7���Z�ϐ�Q!���Py&�.وy=�V��~���8��{��t�F�ll�"���v�o�hh 58<���WB����hc)V:�]�L��ֶl���d�d��Z�K��;�_ f�MtɲuZ2�zu�� ��hM��ij�)ݯ(����5����q2nP�[:B�po�ҶXlxVHYEB     400      f0��Ba/d7a��e2q�2�s�����V�"��;hS��i�6�O�_��g��4%��ë���e ��U"�)��n&�~qPB\�q3�}���X��W��믂�\����,u|�["��H�Z������9��*�@�z��)Er�r�{���4��ȣFN��/�I7^����Йc@5e-���,�Gn�7����i�:�S`�*�u����.8��"}p�ȑdXj�PZ��(��G��XlxVHYEB     400     150���yJ��_�]M�I!~��\$�j�� z�3�������y蠫9�PX�E�k5e�J�o*�-kh���@�j�o� �%�0��bS6��/�_LI�N(6zf�}H�{��Ү��NK�0� S6bʏ�w8
�ƛ�U+��J�hj�X�+b�)�����Q�\`If�{�U��RT�S�;�d�B�6��s�/QC+�8�J"Ѝ8̅�b�g{2+v�U���{��ALc���D�¶� M0w7a�n���'��������K�_I��}^t���#�2I��B�~�XM#>xZV����mRהI ����=���'�hI��_�{���B�XlxVHYEB     400     170l�\��/VnT6%Dt-KI�0(�����I1jB��T�^[���?�K�.]��V(�rW� �V4	��T�8���M�"t7�+�Vls���coX
�*y�_�S.�&���@���b̂��]7�0>����"@M���0�4b�|t�;3S�o-�#� ��{cT�8���-�n�^f��+H��*|��7����~��R���m��:����V�}W�դ2����܈��	�0����o>��қ����[��ӻ��)g��4tٽoI'[��ya\ܕ%_������!~lGr�i'˹~����9Q:*	��3;�Mց�n�(	B7���;�"}>�����J�՛b��լ%���AXlxVHYEB     400     16097����\]�1�	(��~�	�U+�hP �ܳ���8��ob��i%�'ʠ:�A�^f�ӊQa"G#=Օ��j�{z~�^���]��#�u����B�\�,��S]N)%9��B�=_']���ª<�o>#�X���}�'D0I@}�{��`�+�R<�X��)�����T�p0�dUw���5� ��
�>�W��v�g���L�B���<�e�j��X���{e�%V4W�7J��{�L�0�,�x�n���9(�۰���"�}^�����m]�/��/,L�#�ͻ�w)l2;�Pս+#���j�n$N�u�Lĳ9v,:㦊<|��f}���:b�T���n��=@nXlxVHYEB     400     180�Q�u��9~�	Hx���8c�}���h[��z�zL���~�۩1��U�o�XB���pʽ�N0�>�/�ȋG6C.���Q�;C� �����{x�p˅ֲ��LJg~��;��3��M��mN$����
w�1c�댧!}��d4}|����g�u�:UGi@��c����L2q'��a�W}��6,�fϗ2�x���h�a=�ˡ�F�i��A]���@FZv{%z�8����]*?�0�``�$��B(�?q$��}�����O@ô4������~��FC(9������X�[���q�o���Q.���p�e
�~���s:� �V���tU���c�.wM���`�1\��;b��|m��j��~�C���x�XlxVHYEB     369     180\���k.A DR�eKۅ����L���v���{_��3>"ZQ�n����i��y�-M"�L�Y�o>��z���� J��b�Zc���% �lu����@sFɊ���qf9�Z�2�M~y���fU�Ȣ�;0Xt�M��Xy��x��m7?e��ʚZz؜������qP�[�����j�^��A�sKQ�t͛�cO���������QП��<�'HF��{T7���R�7x�������Iݺ�{B@�4������8��/�VV���~�5,�O�ź�4�g"H2((g�+�nԷh���!������S�G P�{�eל
���a7<�����l.p�h�P��L���f�~�t��̆u�!���*���$