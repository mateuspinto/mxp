`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7104)
`protect data_block
9CgApHeRnBxI9O/57znfVXVRe/WHfpq17Jl57Amk6sF/OseWwyku9LcTgzMOHyHtfyy8oQ6kj3qr
t1xtJ6tszewboVMTLfFbTxsbRxC8CCsN5F1qeuStkI2UnqoHDxYdsdNCts0Z2Ck1OViH0/bH52Eb
RfGo1j+HQg69tfg/Fe5ws87UC2ejk6oXIKkxP1/QySE2EFL2flrkvnNxlo0S0kdXsSAyMS7WLt1t
FiXKZ0T1RCzIi07E652XQqIpFn/ISOdV1P8jpY0a7JPBue1h2XjnKxjZ06I3GyN+nOV93IaOyxV/
xkvo/gaFeyM8uk5rqxTP9uSeGEgulXB0PMaPwwmbGxkGGct2BK+r+szckYh71ayFpkgZ1nIhwsrD
c//DSFjZY7n6mEmmBCFCilCXq7n/dISWM8kGpp3TzYV/DNU8riHmFauVRms1ZkWIH3fbWlZwNzrx
eValNTVnmRdbcMzPqHpzUCbvaJocfcDvP41x3qvEJU1v//ieGDwOIj1NDQxRaCEDt+RuSwgJqYbE
u0wRc7MO4/gFjad3L/3fWcwh4NTrRBr9oFsm28OoBuNWXVMEtdPIbq2NjkyDPRoLq/eej7YuDmmT
MvDVYYgr2q9SbwGjAn/nDBnX8Pki/nl/g7nw10LkBlxKO8k3bYEXlkJiVM0hrxZq1siSwa4V6+Wz
sxOwsSTzVAY7Q60sksB4lnGd8UE0cxCVvLKX57orYmWsSoPNRZTkz/CXYRihi1drIC2ptXU717ci
VrlAOIJLjaHbugOHbszDvA37lS3Iy4Ou9SoqdRil4Ri9HBG0cctioc180g7/r5jwXd2LjNyuni+I
n7VO0+kb/+QLdTy2gniTXojo4+nfLBeD+TBL2XcyudR5f97A+vfADc4s7RA1eTnGhDKyH8krNARK
se69wz9P7bUKTDXEaJKtXYUza25UPqIgXRHIsEWLSaZYDVABagNa8vU6127ifLSKGHa+FZwpOA3L
UsEaRgEqGRBoaoH2TYpqm8FrGY5WHvESuJUfilauf49T2k6gjy16HZEALP8qTid4A1PzsmuKQmX2
Cbkjsv9uG3+or+XgIPgboXtgdtQbPHHFTTdURs4zmJTPFN0uCcTCqlm9YzwcZo4YwpsryZwD/toz
IPAIKkdeG1ZeBJg0zp+Ti+8dV5h8sx/HVM4IhCviY9uu1YeTcB26RUwLaBVnvGCWrSq2TIvy9Wf3
PiaYt5o0i0ZcB9Mgzd23Rd0DbT45V1pXYKLtIPG+MMJFYcDcQ2ofNAd3i2WW10E0/dfssqIf6SVA
l/xnjMFZ4+0FWPoYh2JjG5/SqzNbVdjJJYtVdg5AooYWn8Ltcu8PVzwvJWXUtDyRRQLrKgPsKefo
+dnFnaFGzNxv6uh2ztDglXKTanfmS0vgj4paY/XklMH1slBxIkIcO0OPk3B7g7O7O0IEedo/o3jI
h6ByPQP+gQTKxLynWXchc8Mgyy2JmMpg8aeRtyFxYnZ9zn3ykjag41KzOMaLUfin6yn6wW3yQDbK
KxpEWkyAiQZF4SbH4MFjGDrrmjKn/iv3oabW7yvcM5RCFh+/R6GIXxJEjhQ1axLTv49t8cB4u+T9
IgDrVm+H6t73pR6RgbMlNFgiq/dMm0PtVMzXii1+5tFyA5im6VOT/5Dm/0xErJwy/Z8UaT8EdUJc
EzSA/Z8NO7F7pe98nCtoSwiPCMZjSo16Q/pOXgsq0wu0T3hWh8Ftn2AQAJ0QTlXBQGpePtu2ONZv
+TW9QipAlra3NNxb/yrpQZX5tbPNtWS3QwzPsNgO8mNOHQH+11dLduYF3dfGJCh5bUWlBmQHnn0z
vm7bHvMwlz8aXX1eeJnUQMaw15UOi7F2w6t4R25P5pMwIEuJ42BTtQpEqkJskS/OinZpigFNEKhk
5A9HU5UuQhZB/FCkRJlvyeNdKHvHEJL+nFtoouN2rxbdTuOjSplpkWTGJbiptfRE2aI9PWXprMZq
evMYcst0dDAqK2Sbs+SUNbkFnuyLKQoTQgd1WvLkhVzedXfedl/6mgpaByxcVxNDTucsXdTwBjdd
A13HjUVlM6S/h6v2QzzWpkQTyIkx0LS6zrNc4VWLLTGubH27DAgIXb7UiDmukAfAYuT72LBK5nMw
o7g1lz10Tf3+06XMQmjCp7exCnDoPa/WOs5lJ+vVrn7hENIWfcy7Y/E7yNr17bgCXv+mXreZGzDr
T6RP8d4ER6feT+FkjlYCBpf8GaJ83/xdOWDf5ewISFd/PdhEaLLCDWhr0owXmspj4wIs7Jr7zzIy
0wlyY/gHtnU8TTiRBtH1t08io1LYY5jpnH7C6Z+PQbIFO39qLSESvRtrgpuzpJVqIU+gweWs3ZDJ
zSf/sk3FcLvNdwt9OraxN9TfhYg2xcaoKeXLTaB9bC239lLzorf80cAQD3IILJiznIqM2lZtkB3P
LbkBR8tOat+59lzfJBRd1FKEfh1FpXNjrcTM0qyk5qOsvHVb2sAHja8KxWRm6swYfihz0JhGFVLb
eXJYB0hajFbX2q7nJ3Q6N8dG4iKvslBmuiPNELifNizom1aTgQk7sQ2VsdfE/jUadYYu+LrxZnsS
pactUAdbjOmsftU9BMcX37nnhdoKQjyl/jTvCQ5vU72O1Q4glIBJ90DpMuIlPnXmTZNH6LxWvs01
NK3ozyrCZ/bawtuXBDH75PuCl6Xz0aBIqi4DCdKn7gNddMXKtMtNfGIXue55FdgHy56AL4LaQ+0D
bo6KZgA/EdZ9Rre5PhQe8qyPADj8H28tudGvAW6CTmnIXbqaheo6bXm/kU7Dp2CS4PMjRx0jle+z
mU8faPuN7M46/oAgdQi7A4a+yNaoGmBEfx8I4S/OaD5MZxD7ZUrr3iJNrQkgNgtY98rbcOGctiA7
qDHi9YZvinnOmnO0OC2ATxlgqY2Vp/LF/E+akV0sOeO0HP47k49QHVZ8VbSCmDxLzMm3MmTmNAiC
Z9TYFzDtrzbyP/mRMi13xXzyWB3qLTEJ1m8XSxZeY2mxcpugucSfQSLpHo4cEFNYgbFmSBv0xmt1
YVOnlzL6N7jO7lNyGvOJvjMfcUvkrmdvlWnVI1VSGyytRd7OawEIXN64CnTSzCapAykpK7GboCq/
2ZWIhllUoaMPLmua3f9bggebCDNA4D4JdeuKTuNt5FSOkkLNPmbkhW+rEq4mUmLWXBJcKm6u6Bl5
XfnvYCJFE+lysE2AS3/GcmYqfXJk/9kWlxUYw/eHr7P6jQj8jwWTZZLuYCTHCc3XXGhhSEFNhRFl
fihVgj6o7YQEdYu2sTrgAnSXulz3BdSHD1vpOSSkZHUJlv0TIeNa+AH37eRkJuYMcEEYcJ+2tgN9
9R4YWe9j18rfBGi+/0sKfkEptvyGjaS6u+3EMRPZrNqmHfer3SSlYVhsX3+XEhwFqz5iOVPmaruv
eyDlPCj0jAbL2jZrETwqt6lmLTEddW5IohbkE1s/+6AtQEgrqwBNMib9EWjBmqE1SPGv/B1iJi21
Rkd7Sz3SfTGd84eLY1flzCjDYxV7KYCydoMLtaxTWUZ7GljgDNQIu6FUkFj5OcLgUnBCjQn677nJ
YFAf9dLbfHSCVa8z9VQT4pNB3tiitY4DaspmugGW/uFCUmi4nkIV0zaQ3NDbAH+5keQI2XV3O9nt
0OGZUP9Wh9xW8/2tUmqO2axHIYcqT1/hwM2fkkOrK0iYEt+T71/4O6Cehf3FCaKgAABaC7rJanBD
AvnHpSIjt/N1F6tIxaqZXty2Ra453+fUVSwCXjJRkX34REShSTpJavGiNbxWlx2WJL3u34ZZ73HA
G9rzlnW9poz1y01rE6gdxMZgTjgl8j3RKZIZJcjafJ5W0RlPANywLW+ewWAq2L9g1ipwXlLq2WZT
vkojgquBuKplwEbz4N5aP5VyYpdKykEZKOsf6rTeqj07C/la7tGsfdH/InbaVnNt4gMMt9LiX0/X
LIciInQCr/MakM5WUAz3rAU9CnYuLJim9SxBuqVzCsiKc3hnLKQbx1+iSBOIsEaLI/4UvZLfLnf8
f1MX0LkcqD8Y/Qkv6AFVhVnidK8oiufHSPj+oZs1zD4B9h9P5CHWlvY7A1DTVzcZDSOYaSkjzwY2
DYGqdVgaFd4g4zGX3BDc3wktGlWONg80VEKbblWfWh7zyCBcDQNdp+o55XTnPPDP1DHBb/ggLPqs
gy/Yf3Fam/5b8R7ppAm9nmTuSpROEGitODavPA5y3xUe8RAmaayiUHcme4ih50sgfklLYbuNeGox
8ceAhSGDv393LMiMGHR2JTpSm3VXbrvdSSv8s5xXyyn31v/pehmnlOnwOjA5O+STASztzpjxLHE4
fecXXcDMyG9+uIahCJSfrrWVJtVqiGI+51tCwKtZF5XaRJ2B3aO5VLS/PRr2HI4VSY96cxfJw2ex
zXJDuVL/W6ztxDMA1HSRyaAwTnCBcVXWRP9pfJvrkCDSRvvIjTCOyPeiZnNGyz7x5jBGFGb3q4Ex
AW8ETHte+rhd9MrVr1kkhOWJK1KfbO30G9fn+XvaYcuqbb8b1RHwxFQ96Uf1GP6Bnw2W787dLYou
AfnS1IOTqMJhlKACU9Xx/Jo61pvRlq6t5vrA6nLFMXNYDw0Xti2ScC9Cike4zRKolScVNsnLk+Pc
3AnJcYt/5KUj26NbEitU3vCapUSfM8a70lrnpHSD8Dp0of2v1afNVmUHnHCrcy4PE8Pp6f46HACB
XlJqUbTyfL9CJ7ptYlHKUy6dM6Q/+27Z7sKTX6+nxgDkJiuBzL49/0Mfr/WmRlIcFrhSBNINZFPe
NnUSKdtwBwiPamiW+mI7ttQiAdziN7R8IFrq7j8Id3cDRQmnCpr/NMBaM+PmeMHoBOenV4SdVyk/
yISB5SE47fQPqxNqAOq6lvDg9vbp3qMKLvlYxzg1IGyqJ0EkyG8YMds61r6K82oJcuOH3BEUhQhm
eyrRTOOxtyv9JstfbtDlkOFD6A5UdA7y72ON++BL7U0k5CN8IIkGqzRKgABSfrashRj6rtul6tbj
kwkZ5QE6Mx6tzHj8uAxYsXoM9gMFuUMLWe1RfVctGxWRCQXenkq750MKLCX6ld/GnbDChxhI1J/1
wJAqsVowIruxp/oxgAqeGA+Uy1qBMHDKXb+bv9GDbFX+ZdqsVzmIBULYj5kRSNM9nLzxksdpJxgW
gkW7mHMklNe/d/Dho4ggwOASZiohNj0kLkFN8zf/ZxgCuiIBV6vd8ate4h2o1JsMN8Y9sxtMG3O5
7r3K4qlD6p2Lna6cyMuDH+5JMsZEapsgR+1FCzu5ZLqpCTdPHAS4qUktBh5aWp81/tjdN7Cys/tW
2hlSUG5HjPSaTaw3ke0lyuqVSSXpckystt/ABmkZ5s4K/x4/SeeP39P4RLYZsD+QzTdVuqgrLZIC
azjVd16N6Ry1CJ6DZCmXFwhEAczl2OQCjerygE8Al03GcWPp4LOONJno6l3J96FQIUEfZBNy+Zzq
PGbgfxGLlGWnm6ZJ+eeqg6abbxOVl9X9dUUwIV8zLRYx8nkkFpN+dKLE8cGc+8XHPQqVUQzPDC+D
V0b9xPFMegmwfvUaoefJT+YRZowQsJI04u74MpzY9dNGEZwUUpascQFln6NISyW+oB4Lt1J2+qWH
iMste7x7Hd2etrcMMikLTndcaCgrhYF8RjhtCwNIqqUym/NjUvR0m0BgynNhH6UwiXzv+Q69x3N6
LswhztrY9IeojVELLLmCVwBQZWDBs//r/bfJyffYJOCebFYHgGEVKazTtgGueZrY4DOalXvAsIO2
O02ifSVVt10T8nN59uYkEdD2mZ2/iv/kP3ltnuXBMpKzAYZDD+hKFvan9xFZE5VNQigGdOiYUyNg
bxSMsxv7R7D5C8M89IjIhTaW2JeiqrlyvPVqufhKmmx/9Ml3RPWHAupZyb0ZonBVsyWFAqHmG5+y
NFOfdE3JGa6Gwykd6GPwIi9mKQCqSCDRoTpo5oA1nByBQPYVIMnt/M/HkTxpno1NpZE03QeQVVLs
LpJTVMBp4pJoLp81M7hMkT6MW/wopdcGEkupxjOCwnjz4v42dZNvASuaDdkHHdXog3ZcupislKdp
C7bx32ipVwBfDs+XHCfK6r5TnqZ88nH0Hs4WCWTt2lthZJkPYe1GG6pvdpStIyiVsaAzCuumcnXG
MhFn+isY5g4cGXjvgN0mUU2csXh6tmwLjDuh8NwdvByDEb6GexVW3dJUotchwBrConreYxlJPx+Y
M25/KNrWYQdb3cTP6ZQB1PezWq7koc5A1DUKH2e87UZp/IHGgfhXxY+wb7RWqtQKbugdqw6SgaYZ
YWxEFGJmQMZsbCXftnq97i0Ukz6f3sbXR8tYC6erMQxrES+cQDSxeqnk+rxkpQ86/678o870VtKP
2WvzO5h8EZ0r87Ygb/81/O30YeLq6WAUfBc1toVmBrFsrzLn6lJf5gEX8SmqUAuGHc/q1+fgcb3t
I7XbgqgNx7FKrENurPHx4Sv8TAmZdrZYYxo89P85xes7OkeWUK7GWu00o9tVD/9mqz0xtz1L8kBg
F8AXBRBb1YaWDOKPooYwBrBdsV/1LyH8vqzOl8KAyoT9P/mWLKcghPL/FhAShQ15BXm18CwPwdyl
bZ3xQP+IhVyRmJEqjsDp4P8LwyzoO2MpjuWEMsLMFXkQORQrVDbGuA8k/rpw+qAt3wFCKgKpwiEj
cs17qegQGY70Ft4BsTZtrJV5g0fMH0970c14vIDZTO9em4rYexqb9RGsVjcXp3uERrpsmYdzIiKK
HMPYSe/gSp6j4nTz017TE8Ib/QJZksVoxaHeyTLreBejzSJ9Obul0CgB9NP+thDvInIospR/M8mq
wXjFdhOZTdEW0SngUjpWMgHCifdayW3YKjpBmIrEkwS6P+Ct6ke343foGFnHq8iNqOtDHweI7b5N
qDjN5RThujmx+zWw8lu/605w9niWldc9h0nc80X5w3Rqr/6Bmlx367PW1TUd4TIpw3/qryBqvX1L
sFgajKhbbYwYDCA5jdJsr+ebkgdOqDDxkIgqePfWjvV4CxfwFmobaJGVgbXyRJiUMAQb/6UdhvGX
8K9u/ahRx3nZbDKnjp+gg2IQ6VKuJTPqCgABmHnUj4ooLavl4Iun7VApLHzInnBCCgiNa56rFThT
I5UMl7mwGfhY8JkgzUIbo+5O2nxiWUFjnj9hDkikelWOREIHlJ3bX9GtNc3cCufxGO6fUwPkwmZI
JlmfnygUDf3HVcoDWHvK+GaRjuoFvUUGRa08JtG+75QTNV3F5Yl9mRh9yqFrSWXA4bHMlGlv5z1V
n7TfyXuxgiLEwPv3BVtRJPYxKQ4kNsk1ExbBtp83Q6jHbvpNVqXgTpae5aOj0Zi0hK31/xS9e9XM
bjR/wp/X1a6XWNySjggKcF4SMwL/qPRH8dUPv/pJvYoan7MgksCBAMwC2dayc+vg464xU4q2lGXX
+n7+qIZ0gdlJLSH18F4mm5aKC8M//KA8Ti9xxi9PO6gjueSTdQ7uPpMzFq+HacYCCmPLloYoDZ1Z
56GLWiotkKd6RK0RAAtV9T3jN1HIEqEiNMX+AoB3+N12AtvLxJA13OYh1j8N527hJIk1C4jkGgnQ
hOcyGCbEWZ05N4VZglVX7GB8Qzs+zZ0xNxsO5TIi3IfOAu3xhlvdPFl/UA9Jxq6ymHoUbR4tneLe
1AQaY148ShPZiZHde/M3CJVHaM2O3vBKQq48fcJOUmvWafx28hKGsIdzu9OZMD6NjsS1JKlG5W3O
zwPpV1jk4zbGQHCWCVKUn/bCZkutQv1DOL3+E+hEnqBFBGDrBl08CuKg6QRyEumPLYQ3L6355vNX
lajYv6R6W0b3L7uGRtKkNoyZZ9RwPkxJJlpVw+0yQShasuFQd1z8SFarwV1vtnwVT4JJPy3+uu8r
pvOTjN07kAudhKzeKAwlOJqpPcc8zS9/ZeXusx1Hfc6R/WPNnjgOYvRoylTpTXgteGkdMgA8nQkO
rpCKiKHiRKR9m3U3j7PB7hpSwnltaud/e0+WdFboh85cdClTv7RxLyMQdr8oAY1nI/ZeFX5eGHNA
Y1WroivjPPCS7zZJpypnvtrtnZMwaFtcDQ+tAPYmZPloY3OQkdlZ6pA+AWi45IV8vy96o2FlvwNb
5LyNaq/d8P+NBNS7KqBF0xZq85JZ4w6/7GOboNTLrdJqqLtDgyjKDltVgu9RQZmMvP4R60uddbcC
VdcMDKKD8FQg7Xe8ZcQ/AqDtVZBHs6+IMRlqLFXy64vxe9iC2OoJUU+OEw5ZUKUxmufv+Sps278K
qnW8oXAWuUud0otfD4yn6hhtgzwDyRfUX2tdFhvpSkP4MdgUhgYSc/xqAYCq5MWrvYLWmrm6/KTj
RVPbaHCuJ+osLRkoAfLi6Ci3zPKT72Z3bW/Qwjk9HV8t6i7un+UYxlyh7KIijCj+vUCCa9YzXEQF
RU1UwMPJgquWN89UVeWVtKFLVsHechV0MzUzaa+SBx/1zh1WvyoSmkNutmcEUcIYInV7BMkkwiz6
GKz7ju5rJrSzEmdO5eJ17P2uIfCHrM+56XV6tYdpyCaUMaYd3OQXjBErrF25f424I2UUCeJnhsGm
jzkoJVjR/6kpaOJ9ADn6ZGUz/oCVseLxDphPQlAA1GcmOVHk06VIX7GU+2tKkZ7ymu++v4+Nqp9Y
xwbrPrrDBVVrWQ7dgUfpCgz+1DVHPCb2HVLZVSV15kpcWZDOIWjolWG47BJyCmjEmux87fS478/i
f/OQl50NmJ6QZCh/HnL9QtelrYchY+1CHQMoFeKlCO2EP7IwQE2NwecplAHSMSQ9FYgsOAC7G6vt
zZzsNEO5nmRq8lUQpLE2Lx5DPdqtHLGpqUwcbRLaSnBd2x6Ybgdo2QwCMiYeZv1cZfupaloZ6yEJ
QqoDV5aICFzNDGEUCV3IvD6L9cq8tKdWAEkhwdGX0xpo9javmdhB/zzmngXMpSzy6+VIY9LJPkDL
K3WWOaMRIadsjtVMu+MLw3OlDTbgZP3J0OHDU9/yzXJiDvrABIMtcJA8LzcDm7hq7kj3sHxLkuQ+
pIMjawOQxjcfpkhjydRqXdHJyufidyBKQYMg84Xr7NjxRwUnFqucOTOa9LQT1VMZFa9K7IG/qtFZ
Jgi+0F2ooEP8zdsuUh8U35ccR67sL4r2SZmlSqu2ts8IFSvzCl3Ftw9tCHA5rh/I0RAfUiQCD6q5
AWzKiiGTRVl3yVornOhM8sV8mdGtppTP++rnc2stzEa6BSVJbTxssShk/5xmZ+GQxd5tk5dJZ1Ad
uSQaG/uvz8Qmgk475r552BZzEbq4l714V5BCyRlkq7N1dBdEurF6NTrkhBlKdLHe3gGWdz2AHx03
HI/S8QgPbee71D3lHiZtVsiqloy6tfAoyA65YXfA4MdTC2eln1OxjZsr17nkM7SiRLxh4hAsDX/K
8aWG9vwA56N71Ux31UXr26Y6FDE3NeCVmkPr31K0gTPhvpMU
`protect end_protected
