`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11824)
`protect data_block
0USWSUGxovGsyBJteYpEoQMYe57U7EVv4KgCh0gNmqLndd6GcMFKrysHERSf7SgCxFoE8wfI6zUr
26GOa6eQcN4a6kbEbK/OqvX2+AF5Ss9ZqY4vrlC+bupvRd4sT3N5pQDUXR8CIThtR1TUE/FHp3dY
tBQkQ4UVznzprTeOqDaQ65+m2LxcIR4dfxa70vG+fUWj/zS6xyIKEMZIFE9NvwG033K3oFc4fVKp
XyWJNDUHJKOrtqWNbAX9YrQZ4a8fxRNDdEAXceGGWZL7pJQelRuAo8ub3ma1S2FtddkKEqT9Boue
NIJLW90ZJKWDgNV2vht9JtIbpwuD+PzUoaGmp1AL551Klm55zSdbUPHXrnVL4wiF4XiCm+zFjH6L
pWo9qN2HW8ppDSyd3ctb+ffpxnskEEb+4PdEpjioERnXhhCYHSM1JRWqloPV8cvOPdpTC+BWOBAF
TY72Qiz8B1u/lBWQfoWQ0WLFFpgJQNDp0CHCyY/nNohzrnWVTSJBOm7wacZKzf1AHlVUC7/qthZW
9Lh+xNh+Q5mus1HJTnFU8Mt5S0/3sYgDhJcXxmYstjw3kSV956xrzbq2dYaKj1PxfRyXCFe5nRPh
DNfLTNX8ZTCTvcMQfM+PHFL6lJ2vd+6rBnob7IgiXyXyjgBVRomlIGp69Ang5ex11qUTN0bS2kp8
6drGl7MGgT4AsAx6oEsITD82edFj/bubEQWD+UeYWoowIyuEZsw+j0MeAxgKXFzS6IdpRQB7Rov5
VreuMKWOfb0C14cBOOzHfVTW31ATuQhYs/0umS1RAJWgwmsL/nArDTCBDuWRjiiTordEQflYdPrT
rtAoj5pkWQEe2hOhBgODNsnEivStnNEH3eiJhEhGFZQghC8PsvapiuwIdfKZ0LyK8Sizb4wDMUOh
sZC1WeuCqSBJHoGbIofIblOVakW+/5mVGvKOGfNA1uPxzZ8MriR7oG5tOeJSjDAdgnstykf2E8N0
O0jQ3zqyxUG7KHjI3dxJvhL7STcHm8a1jFil8fQ7p2spFGZkugQCEpRWtHzX18cysE4NZXbRTNyQ
IlNDd472zkCqyPDidD78bDwbB+1vz36AE2ZeXmlOIdMizuLfmjW8wYefpuLrfbhKiCbXOoBP9Tc7
kMbf8e0ueP10yYRPTy8n2sl7gFLW/6cB+FUWhWIYcCGe7RAHiM1IdkReF8A20eNwSpZcSpXyjQBt
FLeWQVDLTDXxrMbK0bceytvExyJFp44bQuEMOhXik3C44AN6KYr5SN9YxZi7A9gDAJSrCqsrFsKN
FC/BakmbuDm9g8uM3VVqNiPdIYbvIPqi2mdOuVLPfTnb+wM1fvK9DR05lEOJOWcmOrETmf54ntxL
NlhrVf87nfz1R+8fjKvmoiizm52hz9a/vTtrCVpWA+OJZZxTQpgpooME3psYmc4WEk3ZpqOydsUm
XVe/lswGF6fA5pZlgHO3j0rT+TVjOCjA2WiIpX6eTuTEipywgQ+GrgiBz+3Mb4k/JIsQ3qroEJcU
oSuDyhIn/3jo4kvCP214Xww2Q4Uc3ESBmqR/WrMWsLRBh5KvQJgOZIFQjnCeU2A71KR3Zqp6ftZe
a2yaiWQhO2sFVf5ycEch60HQJYxI1mImI+bw4beWcg1XtXfZ4kRVwfRpf63t2V7/uZ84sw7zkWrF
ZD1/ZVyWhCVYAF6nIG2RQz5RcZCxwWws+CB9q9NziKuLV9Zl3hkDJrJt3H//9VL9IQz0x9IpNSIG
8Roq1Kuf0kwFdaMx6N0eWr64pTOaufaWHBfmz4YKGAvG/2c1h1XliRid3GzrLGZWRB2nTG4T5/C3
j1/sWo3DqnEv/ld2zB+7jHBYWuUyZQ0Kz/NKHLcWi3TGlb7MBMIt6JEyOMUr/YbrSBIlLwpzYBsA
/ogcunSVTdiYYT5qSCrHJCoLNT+GB+m1OaNw20oYY6UW8ocHqJuJdxWZSMTPV2UYeTiFrkkXJTMV
YqemjoP+0VCbLbSKlvv3i1BEm1TmUuPScR2oXz5TK8eRwYLysYClmBba5Ni1M5ulylBmPmNYPCq/
0SRWdriJNAVShP2fF+9XCf809eoVhOnq1pLYbT130IX+xKywO/5DPz6CzVn7VyK3jrgbrQePKZsg
DQpZhpMta5Ifk++yDDvvBmNR86IyrZJflIZBuGYpLrHU72euWbtUBXQzaeHUUsMsd0tX5T6cOo+K
5RElP8OBFLk24HtXk/Ggk/YDnn5npEIDDor5k5qU0UWDZ6ffEZJDLUizCfU1Gw0ii5xvfqol6RMh
lUvWGiGPVSGf0dt4zP3fQ3E2OwPjrtGapZZPTRBqviGVLcdCMU0UipQsX84Fs5htg1CM5HzqElbi
O/2RIfj0q/AbVg40kpmy1smVvnhLP7p16GAQ4DHwqnQjvvSHQ3tW6x1l/YsUfI+8tyc8w3GoJwUT
uFh53g7xtUKmABBmNQmNppykEIw/a7CYUPCIRG23pAWrwWA/yPtHQ//fPkua+NYD9p5QH2OmeiQk
bcZiHoPS2sIvFXTvd2iBbPiEOGEhC53CthjH3wavQeCrQoSk9bhyZErPR5G4OqDykfIEPj/DsNjf
vsM0OSCD7gpBQE0MU/bdpruxX8pGGqTv8SXPZcLtbnNMvUAZDzjkaJ5bq5/5enp0sToFNdVASZwo
RKeB5bqTZQAWt0fSNnzmsZgbmJXk1tYXU/KiTsteOUNmOdCgH9AF054919/jf2UAfQm8pFpIUt+Z
5YTllAqsEPDFJitaHubs2mM5qSgbSqzdVsFBgD/qu7M0wb83v3RpDTUOvaNRuHoenSPAC3AanRA8
pK9mhdTPsUHsOE+cH5NgZCsb1WkD3EJVxujCVemncvkITtN7F5OgkXdwaXSWfTGwA4R+A0sv2o93
AU7NWWUudXqm100M6QuImQL18EmkPe9iILXJugoKlpoRqUHpbvs908B1rEuw6CYs3abw9K8y116u
j82OvXhqsgutIpa/uiNJDX9mF4k1xhmI2Lopg1VQleQSd26JVt5u5rgz5io9DB+CbxrwG5wk79AV
K6W693Jw1FdpVOdo2h2xVgmkYi3PMoaGDVlrjP8BS+rdWtjvPhPn635MliurhGI0KzKGIcW4q38d
cIZQUXXeFAgcv2RSQl7V5xXL18BG8fqm2RiH9iWQV1ZytVd0j9wTTMPRMOnbSvL/4p5Oxzg6nFfk
y94Vu5esgG/8GwPSfQshOIf6fecokJ0tNdO427b/hornNCtxosH0OdATWXV4frWPmTO5R3zOziyf
oRiGn0C4X8hk8Bp2vac5SpLGhCIrsz/4gHPQHRqhLZex6joW67ia6mimT2K6V17IjsBzfPIiiwM6
G0mFFxS6UW38NLKAe18Noc9YZ//5NjYvQWMc2+qRPtR1wXaW8Q476aKmFwktkB0KKCLIFkCW3XXw
CN2uTDRbSeiN3WhGGjhtTeF+0L8eUfG6QUIDl7eVcVY8HEFrEpngtMaXccX5OQ8R/SjniKY4UAv3
2klU2rexGjd+D6UwhrmE6BQSYLYSvlNR2UeshsxugfFiLbHmbwJ8lcR36UBRpQ17sYiFMDZhk36N
WcrdhpJjsfU1b98VXyKamhPsEYznSU1JV2jrCiSchhsQPTbBKG33QvesrflKsuFtgN4QslxwWH2e
vwud7vgUmyEYUc8MaiNS3eVdyNk5j/eENoSXI4Az6cL4sAiUiuRsipAfjlbLbF53E0xe/fXljkjJ
Hr8ixx+Y/0yosuTLVshm0N7CajgvMpeZqZQon1gLUd2XQmg7dYAfO51MkDjJIaArbn6suRVkRZGO
DTsja1CZmIMOhSFX+tOBFkk4wYVztij1l9FVY53gMNcgFHaIUMoUJ1zyJjyiwcTUuX/wWkyZkKHD
tJWt9dshW4Le1ovzw60eikcadaxjqP+qEPYg/2ZAb657tWDNUwRucS+YjZkABo0AG6KX4n41lzu9
1DrBD7x626LslkK9Q4DRAwcZG2/BhYD/jaMYtwsFCbeojl8P/6935iJiS1o0+LN7YdFE75g0mBwE
mlUgsS/z7NMbKrQdd58zAPl4kcjNJtpFXA3DXGR97CPBNkf1IidbSy1rViFuk7D8MiqxioNnDThU
ovIDaJfTRSAAfiF00HwHG46azNQtUlGraFXOKR1uEMpKE7y14FwkRv4JqAb7+Daze/vjGc4ukCEF
WQhUzHCBDgtOgdOAQRaxU+ammmlZLfBydFcs7BR6QmL94nawcd5HyX00FbCbS1fFDzMtu3Q0LCIZ
95/P0QgDvQNslCrbm67vGVytkpN6levYiahOqiXPMgNyNDvgWBVoCvGbatJEEfYgh0bZzC9NwmU6
kpDpxBgjEIRgUTlFVSKi51+Y+n8m0E0uu6Hoem0hitUxnc3hXaADfTKdI+1RFC4sylJL6cZRsa28
tHJWe6dgdzbbJaqi3XFsZdaObF/t8Er3qJ2TuIIjf6J4NvX+9Os2ZWrKhgJvblkKit2EurP6pfna
U8KuQM8fdbiyFp3SkBawgn2CAc1yL1BPzq/p25OAyNTtItDrmQkoJeNVYg8Nw6hfguG1Eoe9UA0S
TSLXNS1RwY6RI779Vl/I+SJLbPLmQQ+xzfh7vfl7JROxX9tqJWkzzwulLo1cMgw2zZQz2lSU0/CG
23nfrfh1QyoknjCXzQPzIxsAEqUhZmWrxbD5FHGhAqlEzQJtYoCK8rto3EpE2zhwz3oR0Yesh57Y
mqeroPbqNj55UBoK4A/JRruWgXCyvhLJSpLh07HoaBslbCv4udE8JiOiy+IZV40aD2r8bMHYeIcK
oP7l+ZE5Cd6i2Ws5RrbSmcV7P+Cuz8PDsIloHVxYpqTTKvlNLc55M/e0wkNVxkb40Z0KhSelkc3B
6xrQsEuGik3eYXICKXbDIBuzwgLu83Q+WJZ5/3yn/BSDvrgL2kjOQE3sFILBuQoGVd/aRL2+t5rh
/1Qahv3lYhFT60vOCUA0hNuzyx/Hrm/8HxKurFKySJ8E1D0SUQKzyhyCtNXd4Z58gN17doBEReZO
h+f75htejT7VIe7EnbZAR+SZ5aYiILcJn8TqwhqIijdCZBoiY37qThf9j1UuhGYStNjZZtz6uSQX
KvPCSxBqOqQ9tGfGjwYXq8ZXe6gFSjTAMKTl/OLZshmIr6irZxyTed/AezkekEq2ZWL84sPcE6x+
LM8QHm86NVLcbGZH3wRvZ4bPSAx4giJIC8hG28yqDu/I8W0mYmv/G5R0ykO0/UzmuJ1x3nhnuvuk
csh3Y3ARZ2JvWDcQAn8oL65rTQaG7qZ6BgRHAQss/1h7bp53a1DjUzuiOep7zuddsU2wONA3X4pf
WrCG5SenrE6sI7LGNY7inV9kg2W/nmmmByExCAZ+KJsPVR1n5hI3m99bCOzL+CV5KEb+TKFVeiR5
nbsJWhtLEojFa/WW8UTrW0v8WrHLjVh3fY7UAPhNTGli5JnQjhmArgdeviYs0sQRsp581VEb6Quv
ucM2kFS7Ej/0exvr0oyOqLfY3u2hND1Yu38PWAUuTLfcyQnMLjbdmiC2SuOiOQNe2MJ/1/fSB9zV
CzbKTy90moy6Xj4g/xcehsGkXp8CXKarew1s6yp8LrptOgelupwNF5+gLJxFs8eY1EAaIH14MGOY
FhDvrxM002L6d3l3lWIpXzPXBFQRszgUEVrwjIRyFZO4OgGtLVaOfuHOf8fCD+oFWquDbfX0Gb5W
LaikJ0GT0Z31xWhbW3nyvAGc2Aq4RIkltn6Fbqroaw6tMGGQGUtl7775DmWdx3/3SU7+mdCKRpho
w05H0Gdhik2RdNgzZWrk+jDC0YBsJJniKCTdIKTZ9FpIA7PkF/VzCDM9Qgks4RUYd+3dXxIqb/Ro
RMXhWzNGtK0696fGSZmhX2riU7Ikd/DtxeLW5UGxHgoFTk6KFYqofnMc7WVr+Z8odB6CzPJw33JQ
+lJqCwgxOmaCikgrR+Xl76iaYSfwZ0JTBFLfkYwGxtBtI4NAUOqXWswq/7Emo5t9dcWVNYkV1z79
WIPatr8Kv9LTsCq7Ymd8LOYrIFmLU2XpMyx8HZBrI6Fa2fSjf1mpIbzm7Q/NE7fNKlJoE6APgPWr
mO72CzhdiPrN1Y3Fgdnsqu++5rtTxfVvkcjVHEo6ZcjWoqG60iemGToDHPVI5fcR+VcyebfMlv2Z
G+A43WXwIvnWsGaxn2g35zWSU1Fwp869wLYxi21hxd03TrJzgl8w7ZjeGEZhzM+Jx+8rlLcJIdVX
j5NmQr87LFNfyytJPwNv8UIBZws0YOcwCaX70J+RR0rJqTuOm19Lxjx60MRnrWOQmQwQjXAi8zBf
y3Kl63VYkQo8dHsvj6a1wg1OP3/RL47wnmozOoBJUP9U99hEhjDTchIZDVn+yp5bq9PG4UKD+zXl
RmYN2YcpyDlB8D4Qm6BvpJhqSPYRXspHRgKdG43Z2yUT46O6DBxy1q1tKTRl4a6OU3hqJ3ezvPZb
WTKmL6IKTgjdAMqTW24QkpLeLiyQLgf3yq6BZyQ6JmRHkpsHig8Q7zvEgstngBn7XqSewRlt9dRi
HUq0yXyleVmRkps8v2ZdFCJIlz66dV6PDpcszuSfO+w6BDnkPSQvEhagVocPTfyARa5e/c2IHmgW
rK0je4HUb4PmyKs/MVa/167UZxo1yJjE6Djz/RlnaswV8C3MU2veJThOtowqjggxGpEB6BE83XfS
7CHC3425WMzDwpJlopyMrb4kPOu2Kl4JwSghdxWs5E4Gf77R1TOlIvUhxs0QYQsIVZGm+6FwKM0l
woVhMm7iW6wsBrCoYm49EkarjdB3tYzHURgARlItT0YlVgtcJrcR3gZZkONXiNUj0AXvdnYWixoc
XIQZFIlY44vlbW75FEJzQzZtszlmFUeJkzWtqZyjvFS6HFSiybcrDCfR7/rG5+Vsgn42A7ZxGRrY
EXvW8SHHc+YDqPRcnLQdm/CAeiPl7cvtGnCmB3hcJIjeN+qM3PxritqjC8XGRJXDzbZfJzPq0+jO
OPEim+7jLTp4UdIXoAceodvPFNrODt4cx2CRd6gt3Havs/hqPKvrR6Urs3Ux1Pmd9td9lbINZ3cr
5L2n2b5ROMIjkMXF5lADK556Kw2cv8upAidT1Ii9yjzFaoPsBhw16mR1kqFKFfaDSl/s/bBw/iM6
7wfuaqvUOvgrohO7VidqrE+EQOwaL2aleFNHa1Cy/JBDei9u/YxiKCIS0RW2CdQeJMfMltcz8+Af
qATT8pneENICXaXH0JfASCByW5mk0CP47w7RNEUqt5WVWwbsO9mbrz2Fga0Nrixti1Ycz7ov2T89
cmVMPWeTG5HMR6QvOo76xEK682Y9aB8teUsepxCSuIneVlrYSnYrihWaTgsms8La6D7x5VoeiRWa
XyqjTpNT/4b14CYQOMlLgBecxoriNOen2da5pd6eQjKBRUvnJFJi4nJ9/itEnXhX0JYsVksSBbky
ujHExLsj3PysbxpydgCXdj2NTEhKPTu/RuETCd9R0aBUJPoSnGc+Bx2RG6seZBvCi6lM45Q3hTkT
BI9CcQbYcvLy4pVotkJ7mio4dPyK4Ywg5VKdsWPLTvXTZxvkLX8r6RAqVOh5FLLyMvADA2Dy9Z9F
CQ9Bomzbopx7RXHpP7Q5ODUXBebK50UfOgiZjFPo2xVzSXY3oxFrHTEMEvu3y6KpC8jzSPTMgb5H
PhyGuFWsZJGJ080kvnxidFYG5/gxbGpe/Y2dW9teumdmf9IjN91NoC1bs65An511pONDspWGURsf
0Xeln9EWHpvNNqoN/C5LDQ9MbLgoNzySW5GY22h1EKIjDwlhw/7gh99o448Osrc0FGgvKcrvYh+t
Z7NDWjUdv4fctsLgu8RwosuWJJAJN7HrU1lPfwe0m4dh0j519My7ePECn9kPxG4G7vMPZ+Z3GciL
Lfi0eljO2Khu0eBvVi8rU79ShbZ/BUCa3gXYBBZ08e836TNQULMD68s6d60cCpHxIRliaAoEYUdt
Tb0HoFiXYrpAyg0daoC5YuT3d1pUnugTNZyaK8EFNmiljTCFiX/ubG6cTDtG62BRDURJtA7LkL5L
zmaSYzBeCUTnjpY8ug1P6di86Duf3kObLgRUNsbPWA4UatJ9lJmVsqQDSb7+8gWYTq/V2WJVTc10
L/lNyEogtr4SxYvFpu2d2QH7gnbleBsD0Ld+iQeJDwEAD10ggC9q4rCZs90MKeRmhsT6C4cEmfkH
eCHs5yvr5uZpLSPv7xbdBkcBbtvphDKT/QbD/89hbb4Y16kcyYdx2JSyPdUgYTm7uXQ1GF5iVD4c
/RSwzItLNPQuSCWtfyI6wrCJ0GeK1K5W7JR/LZzE91HYJp+FtScFSa8fKr5Ur9d+DelEuXT0USSD
YcHgBszcE8V43w//1a/BIpbl+t1WaVa3Uy4qWrd+fhuBWSGJ3eyDxWdE9gxsknrXcnDxdaHSy86U
hYsB/I1y2BjSgZ6B+TxWup0SZ30X4PXlEQB5fuyI9iq+KsnlvFEZjCEd/w1e14tinKlz+FE9sEgw
iDzkcJzOp3wTooXpiERrwt5UpUMucSGNyg21s6bXHRODQi2iYJjAzqueLEkVUnwaYtWpbYMVEMN7
MUu9O3mKv9HFut7+5BTnLRIsvwDn1x06WpHjFAYUmhotBchaCHsjxPbFoytf2GUbu6lI1IsMOA2K
dBTPRzxNDmMMXIN55EvqEf+Fa94PCv3bshlWUP4pnXIg9SUZtsPmtdG9EreefJ0Xqln9lccrKk1v
iaY0hMIYoqcpjcLGJZ9AoDlet8DbgeJPjz8C7DD7p7Z4y71sbBmCUjjO20liZsIhFa6wxHJZCI+r
Ia2Fm2i4Vt/J/u48XjPGEBBWQD/4k+DSfUWGcZH0jbZN58XhAUjEP/CAqcRXyl2PZX9262FtfKG1
g4b8MQoKWywW76XlpIPeI/N7ECP54wEQ6l5YneYnpR7exb1kNSqVDbR2jJ3Ki6uMK3RVouVAzyW5
cWDSWxreJ2G7H6ebxvA5NAKedowXrKE+0FHqNr/y7iGfazWN3nXMcoB5PYjKRSn2B7MMiBUVYgh4
aTkOsL7qnnEMNJyeQEmF91+sgTiDw5jCe5Ce5ZLz1lVxN6XcvSfTgd8id/JfLNRDw0U6/8xci1i/
cpld9t1+qtEhVZHzpLQhT3785FBBVP5jO3Ti+MeVyKPfbA+zCzdzbEPsGGonGGhNQSERdqxiU3Za
GWDk2KUyAAvV4m+c/oAMxY0MmVD6qNcVGjj+WP5VMasmPWuGwA+AJ7QrFutIoyEJaLSAXxJBPRAc
ahMD1tMpQaaQbUW08EtKVYulr5QTW747CfNeESaPTPHlu4+5Abu+iHHeaq1eElsqvashuExLTTkb
deMyrucUlhDSCbEqryX6QFay2utTpRtSP18dCtHh7Dkive9EXzi944U+A0CMjJ1kNieMlCzfOjhQ
bmGC7NwC2XPocqgXJmiTslowxYMWvqDB3XJhueW1sT4/u3Y4JSs/9yG53yu882c0Kl3SfcbBD5mj
fsZNXB3OaievLR8+L+Kdh3iWelnvaPYISVpvJDlW5rLMlO3HaHNZOCv4oujeLEghhL56IAcDCvSF
KE7jGpyThcUz+w1/srV5/Ztz+DdgUnE25fEXwIQN2mqnPHalGObEffQqizb0MlTsjqxXnVbPf0iR
X+vO5SiU+2nhFvbmvaXIdtDTQYXDuiWuL266w+D5nSz1zmHpInoZcWfeQ0pSVyvKbbXn0t0hwpKe
gttVtyv+CSukainEmKta/POvM/os3KQLIbvXCrkUdOIutH/GVTl+BvGbavowNfSGT7VDbqV7OKI3
3knKYWvSash8FrgY3jiLn3P2qOxEcclkpVnJZLeiUtn73y0yMLDyNazZLVkmlzXWqTgG4YtxhLiq
lxoMW3fiTiGC9sGwG4IwRiuylGFS/D1xeQJan4brm+8AUwufmUPdtZqFUD4SojHQjpLT7WgVNObM
nojzoRfrArFG8nJubd+HiNxQO2JwQMq9cIkiDB8U6t0O6A9NRhoZZXnTDszcSWgqeE3FOU1oqU/m
xmgE3D1lq7uisKivrlB/z8VwzBKmOcDKumkWxkGS7/7UOdVM0W289HTniGO81/a2eqKJqrkk0V1i
yB0RNIMfGD4iA3IxO5vZRaFEgyBHiuTURM7pko5fkS0U7ZwDeY/VkuvSs/XFFiI3ggp4j2rOrsXV
b/kPiSKWLzjc3QXqf+dFGMKwi0Vt7L67bXG//FXBfg/wYq2pDlSVbIMfu59ysSAQ35D9HEBzycE5
aq/rh3y8VlNT+7Ky0E+/bsy8+O/sb958bVHCqxlRRyuobYv5t/dqgCfn1oJgdZjJp9S9diGPwn/5
RAX5aFmIUqcZDZgCcyismSFHTWH1OnwuLOQLy95Op1jnO33IzwR6qzqBlt6cLHiFM7J0e4uxD67g
adRR5iXJFRC/cdKzsjoFolgC4Pv+gTwCLjmuDUp6PDYq3zuhK3fg4cn1LAl4dvDAVdMB7kazqOQ1
uC776gZxQ0KcfTq+iBabeDji8xt4f7iWJVsCtNLi6PtYnrc+wRgatJ7/Sn1A+VHJN/YSycSIHSz7
dvWX8G3GFTXosPjSZtKjdXazdw5XvdcGYklM4azRNZVy/rvommG4qakgx1uOr80uDVwUyjlLRYtd
Yq432zSqpFiCzc5O/6mUGgT3Rnw6hJgnsdMjjoiemNIVpQ7C8y6lp+uCcnSrNhu6zH/TMAQ6SCFN
VktOOVZ2y9d3RgO1ZphJ4q/Bs9dVPf3C5VXUz0w6aUIilD8K3Vn+7ZPCs8p1Omy/pNU/Gkz1LDQv
E+TYvpH+MQ5zWEyPkZQW2/CkWGNQBjSSnH4SmC03zGk2QZEF9RaT+rWFvZm4w20mQ3X1oJTAFtwh
aBk4YmviMSX+1GoKwFTIO8c2PCbMH3kVSAJsqwLr/+D7NJWliSx5jhGnUTcEA9ZK4lm7J5ip1kih
OrYvdJ+l44w8ptDcs4H1xCkIhjt4wkDe+3nKN1PhKRK1qJ1Lf5/0+ZS8kbHn4u3bXNyIUFN8tHRB
Kf5c8thKc8fCwjLkw76hL64zf/kTHuxOuhmd6sSPSQBIIOR6md7dmjwD1Ois2FlaZcZpXHPaxNZJ
ZyqWLIsAchmPCSVMDwhIoP+5k+JrdZx7VgTFfn59hWenKoEv0CdtZB8GWij4j8JvgL3ribgmYqxw
m5LqPeSzh4uf6Wsd12kIHb3YZC4g7TFocBTZNBe4nEyFVsbjT4XacGapgRLKKR5kyjyUCF/pKSQC
jqP8nlfu4ILI/d0UTFR7pyZpoUcjRKqEbt7sCRMJG0A+UBhJxrss8arIgeqE1jBDbv91Q+wZDQw+
wZR0sA06Gvmg7y+MO2oHl6y6vBBzJM/BosLUiv1PAgeqA+4DqujmAAHZ92GcqF2qkscgcZ4NoTmr
OeZ7pDmurBOnwbsr6FRhGCuAUL1RPEkq+f3epItEoqMX0qr2jFZ4Yr8hCea3gmrjbcKsM4cVrVk3
rOzSgnNchuLkDvg+T7ceKAGHTp8h1f1TiutiNrBNAnWvPqlNMy+I73HOKpLnBaRj/dYJPkG518CR
kpNDfroPYWMByNeAyPMClIV6XhEm7SnXtVpw/bhmX3MkBc8k2h/qpKKBArJMbSBq//H7e5dxc8Yj
UN31seL96iogy0piWPJWcdPwEYWqn3LO/464wa/Qqr+1KmxYgHgYgnd0RKb//hiBMfKD9QlDzMEs
GEBtjjJKeur5JOJYM8zciuft3PznQXrBRU/doa6xJYdMoWsgnh1RBFIuj93wUlPJfVk0twAVIir5
kvf9lqVoXwDH5PeqvJYJ9gUufZYJ6SY3+bAHH+IHrbqRbw3iv724jXer59r7n37xXBK/ge8RyUDD
nEOH7k/VMSC6imo0eDClZfLnky/vqsjf0svJrtzMvkqpQLwg6rAGSOGn4DTk2rEEAbMdXLibFe2d
OWwDR/pw5aF/BtSZ7AQF6gNenmt64i7HjodLYgGAelDrayE2dxpKaPcQbiIIJw/zvaRwZfDs/s+O
Vm+TGmYFO5naPJRo/xomiogkGZScPrdpJE/IrhZ5I47ijJxt55doxYWsHthbX4NKt8yfr+FiW2e5
JJUdFcUOlHS+kdZdK4mM/vtJR1MzmtEirMJ+Zhwj/rVlwmAT0Bx0ElsuoAwOhxGdgvhyO2ccAchv
HYQo/MxjKFErhO19AyH7TzG5qDCStVIq5QkhNgrvkeoYhkJWDG2A0VnHGaZIzp8H9jeGXWsnBLzF
CCwgojD9o1HFO7GU+p3BFCGGWO/AQR1fIvyjOMXRsVidF+yk7oeqPO/IkXqREQluwPnnWoWxPWRV
nM2gJM7WpZdLFinIGRYntLbE8UgHlG+niW+7ROR67UNsz8hAOlPAjLwptoG9nKFh/nTVoR/Wg3PI
naIYYZKZ2npVU2BHlnT2LMszt6orqZtXPBN+lLMbxxBTE1x7WXNH5HobogzH6Jk7uRFp2fkDjK92
QaK8Q6G1tHPtK5XDGvNqzdNlkfEo+ksTKJ436plt+MOXmHe9pN+aNgJU1JX8JWziVjQxjq6Ru2YZ
czFGpJPdJ0QL0fVC7V0Xl7EC1RH+5rpuiYYxxzGJ88fMqyfNlQcF4IEsqJZbIWKxQCOxidErr8Mz
ViyVXDEP+YU3WO3R+xSmPpeuK0mmkompsTsHSsDNm/O1zqGIh3cs5K/HUPxgnmh9aCDNaL3YkBea
OqnOZzkvvHaMjCFntiZYXSI9DO1eZc/XZHsYbbvzFOy5mzpM8yGMJWxrIp3PSITXqqKeekj0jEpK
X7C11XwoIiSr7CAEqDRRJNETmOMnE0bPNvdj1ukTosm8u4BXPUL4XNRN2sEP3zhqJOBc4c3G2cnK
0OrPlUzjfJ3zlKHd1HyW/8B14aURubRNCTcl8LWvRMurTaZ8jtEuMwuisTC68BIJ87Iwo7mYzuLY
QCD/Aj5PDtYSrvGqkNKb8D9uwzB5op/JxZ5sqNFWVWNEKKsspdHI3oMk8eZcbKbmwXCIYzvxAIXZ
xno4pUaucvzMAOq718GUxM56bsqZbLxHgWzn9We7Q65QQQyJ72V38aZThyui0AGzZMUVCvPH220r
C1QTPhe0kwL/kp2Ym8Vjj3z8Q61yMfg2NU/iZwR5BRNXBoKZ+ao4qFFZVDzBsl1orgFQg+szxRfj
QOhB+vA4S/cgXn5DL7JkKdSo1eWgO63oIiFUY2j4lBrG1IXskPa1VxUE2P3QK6Ll3JWD5ZqAebK7
Mc2uzr+cGC6ZncSzEmtO5XDGK7YFoRfqpiNKL1/Lrhp3c9JU6tXp9CoyzLtE9yeNfk52xGLFw2SV
TCIPHYE/S0fkyq8ulYfjYXrC+uIUC7nYx46WDQzSBrXVhokpcbGO8v2ZPiZAN5fcZFpe4Xwe1iqB
TW/MKRL61SEn/m+210qN2BACyyyERWr+Mk8izUr2T09K4j/O6C8Ymr9scq7oHDMs8UfKfWr5hzRE
SKm6v+nTvJpNF0wG9JccvRBZl9b+JXlF8x5C7xd6lPER9Y4kCLDT3t/74zOmWz6uhN9J4tHjCw2K
nbKzWjyabaOqJPwaR+2lc3qLVYjQmEjqiUqqOvLa0O0XuSLgSEtwh1p7su23BCS0UJwhlx0xfRcY
qNbIQB4maHLqg4H/5cESVRTNKj46q5MBtzXvFmdCl3Ti0H5uuWiH0uXK993TEtVg49CG8piO2h4z
j/oFH8vtPOYjBCEiWs1rgiNmnGo5lSXBbNvjLlbzLj/Dt6H8mbQC+NZTTWI/l8h2TG788rg4Ka3T
QuJF4/0DvijBb6zOSQltyxppraCBCCdATLlHbCx7VQqREOMOXp7spmbd8D7AY+syKEQ49r+6AioD
HntwYNKGxXPBfc5OsX0vGwqKiGUAROE+flgz1j+p6hmhpK0wxYm9JDhzZTvGlVYCnMSGqK/OD85n
bMIgxiqFFptdjGvu7ZgKDd0X5zAGDAOuT38HK0K+ucp098vz/ixg7kSq2naOd83vJPFbsdC58r6U
1ftmUKeairUglPfVXp4jjPy8FuJ7rg6yTvZPRDxKQMGYYIvi1zQZxgC2AuTIOrC9HDij4PocUecY
8o3f3/k2wX1I6CH+zZ8Kboqao4XeD+smxCZv5X1vfTzxQ8b6Bd/B1PRwBx91mAr/MOmbKzkOmNwy
rmqhkJu/WpTo8EDj9k3+z0qmzpImqhcuErmYNUzz1yoSeE0dS9ChxdBNSdGUMHM1c5wKp7dN7CCG
ixvkH4FMeyzC6gHHqwCz4cG3a+c9BrIZHci5Yc2+DuH1hx6laN6jTwVKD+0B3lo2hrA+EkbYIBcB
oCN/vq63LqY3wG8o0N6yovquIAfG5tg4lpgLSyFzYW+RIfV78yeW3z21B0o0FtIHJeTDtV7n7Ehg
HD8lzgvk0yBLWEOJWvHbuFwTk2qic84i78SnsIQnpJmBHR4DparhSQ7/wl5BSJO0kSwb1dkzlLDF
UEjttm7pFpn1xjq9UGb4gjC5IAfopBcFgaQZU4Sd9zzmAp6ucuympL53DCmxf/jwM6IhNXg48CTU
GqoEb4J20zYVdN1v2Yvvr/9mspDPm3NIrfVIFhHrTkIbynrT3PskXcOWQvRkD5rsXKi+PZeUhnfI
8Da4scHtoqoWZCLxiF0SoCJoHLQdWW/Ia7kI9uVEdgccbMVVVL+xYEWGX5av7DcyX71OX5dxvW8k
DGd7fAh9pMqnKPurk3EygNXR+qVGavlWYpYbv2rCghsZlMANr+rpNvDYBioS9Ur1te/HjyU8DVwS
hdnKCDyGoukhOiq9BdrE5rDD8dIssNEH0UW2HmXDbOc2mhCxxLiLoFP0O4/H8iLJoc00ka770SLj
eV1SoSo+6lKPVkEU74urLNbK2gQEia3eOnOPCi6gF36B+g/aDjQq25w1n3NgVe03DMrSZzdemqeT
qSsErFLtN6qDRajQODNphJrlXgx9gFiueuj5mobNmI02At8kO4cRkmkwEMvJy94f7elNza5dfrsw
36SWpZyRk1BjrynTBgRhnmJ2n06XM+BzfDA6jiqXyDzK8YLom68Lm1g01K3DRfxPmEttXEIF3TrR
NV/m+ehPzLermAPSAKC9sAQMts3CswGQ/6q49hxeIIQEzToxZ5jt8PzBPPA9zh+726rQPtO+4oyM
MRKfS2EUUmo38PRxbxMnn0FAYRC7nrPeQ3/FHYGkIX1jfklhtCwyij4PHUhQYH6Eo3v4ZKKCtEBS
tSbX8byWSUV1m7pfg0QWjYrPDa+tXju+EjcqK5zhtq6w4g9aQwUltfOxn3jFS30UsZIbO/dZApxg
whItvg9ZkpCXZt9N1ePUpep9WCg7DkhdQyMgdy7ykIv3EUK5ZtbHI/gC45O9C7JT1LI9/q9/m5cj
A1wCHRg1iy8KezYV895wRkuiI4i81gApFd2qFppPzFxbCTMvCerMHh0AEtGOlg9OfRtJcS9QAdtX
CKagQvQwLWvOL+dmOLOemjK/4ajasec/17zOpcsdZYpTc3XQnP8dUMfw5Vxym8pVmHfbpvYqqUFF
xvPy3QQw3I4NCGbouYxrb6IK5P+5roK36Oiw2Bmpo0Grre7dWNTW97bU04xf1NtMJtycRRUz35FO
vNZuvbUA3foQeH9WIBJb+/uJkpoDY5Yjojbt3U7OCcRDd8pCSo08RQKMFHBSRFr2/9KYUnYVN1+C
J2ghkTPFfLuuWPBG+Sm6t/RwhhNAh/JfoM8mM8g6nB6fB99eEe5WgLyC9GmsvnBPiJ+dN+o5HMqD
OHmW2+jgPx7Xv0od4liieUMAKVuuhEcrZQ==
`protect end_protected
