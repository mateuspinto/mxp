`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 73904)
`protect data_block
eH4z3oAaGCcxMDjS3y756Xcd3B6U7bp7jh93/c3FvCGQikRptPOvuh9K2LQAvimNsJRngx7/5hL8
MwUamaa8iP5ivZGguicS3BWtYsooH/dYpom2sAIc3lNSVjvlTMn2SG2o6kcDmMxJqwiRoo0A3I3e
AtKTRnajZNUhVXqL/vr5yeVYzVrobVLaSTJcPhMrxxqaBTsIfn5L605eYRa//h6rQKNE22UeNbCE
DhQA6ygSFzq2rwhc5vnknBTCpMlCOrFEgNa813hsQ5Q80+/rkJPLP3pawpVXPlxLE6T9G/8/0rF8
OXBKq5fxiF4rATQx3XWGlvaqFBx2SOEQzxWNZCvmc2taa+IPnzE4vrd1Vs5C84/tyl0Ze42xsi6D
GrwBLV0bDoChmM5HRH3bWMhJsjKwwCRNheLvDvayiAjrjyQJdHBNP2yMLGCe92ZZmVoLyw1lgROs
IpH6qLGsWRyb8Kaq8M4VWmF9IhHIxyi431tfUHfHLj8RjXXxV/wq3Aky0mT+yTpBx2gg/G3GKhDn
2VNsupUcc/y/o3cddnTFbzgEEpZblO6e4Cv8xYzsfVmk3TJ5YDyPcD+qBp83stmVO/3beQGwjk1P
tegQxZ9tjdk+dFeM1OsaR5NFeK2xXmTWYgpx+GZRoU2yuqOcUmKjrdKWrMV/6fFvtDnnr98uDd+N
T7dwgslnrQjZQ+oc/XCgDZxndWCdRW36PKs58Tm5dkwGs1HhJPtLLaec6uRvTrzUkMD7HBEr3TPX
FInfH7K2qFP8mQCwyHsN8p6TGudFWz153zPfHwsVQp0t2e6vX0LgzqHN30CRfJ2ybFscGcZzX0A3
PheNWVTc1GymUQr7w2z+bGD3iZfaUavgiDfGJUnmErhTDdKCDMKqHk1+CDQ/ALgWdRQgcqwMvvIN
AXZ/OIxi/oj6CzulCMNQAdb9TRT6DzMZGJ/7PHlmrsKd+KyRHbktesaLKvz/xnhmOH92b9nALab8
wn8E5iGiCj6SCVRNWdDWJ5j2UutFS6QZP/N/JL9oyBniovas6721jVHvl4ueetO3jspBCgDgJzBr
sBJ8MxSLm/fgZa4sKAPxi7UiZOUoGO3dHu9iRqxQlPMeTAfPFvGz8p4EQ4PCwcbWD3dRvwv942Mw
Zsy55HcLrjOnZkrjQkZy1a8ESxtsx0s4BeMjMKzvgvhvqYCMbN0Lf2RizvKSVz4Lc3DhkhaKHiNY
+usGYxXVxIwILea7djmZuXUDIgZrRCdQd6xIIqDmnBuwi0sifDYWpWwDSd1UX1l49qlqAw2wfFZy
QA+V+LewD4+4PcbQY6gV2VYYPqiYUhYDoDo6fXGEHUxDRDbrsLLeEnnwNTQt1HBiMHZUDw8EFwkj
LCr/64l4PvfkVV91y9KJkoTphnpNmJo9xisNpr5U3aN3ElCqEDRYN5gfDWDz4t9MlUEqTOdJHJlg
95JQUprtbQsnEhQKHZQohgp28QToPktJxNWbo+Kkp5TfLxSXZyA1v4YN7spX0ngHPtUnX3CDWLST
NZIQ5RbQrLA6H3DIXN9AkQ+AzuKJvDC+l5JZ6v9tyWddcw8kW4F23S08rQXAmiGkvZuFJAbCTOVv
KJKwlxpBkg51XKtvsfqi8oOO+5kCeP99XmaXO5o74en6J6LFMqoNIAb+MfkU+RDSvyH+dFoDn3pH
c9BUSTALREY+9kJ9teydkvyXYZRmp2L1S+YlgvCryaU9ZcVZMOkpA5FBLdlo0QvHTEcV5W65XXsE
XoFq181zWH0WUxawss2Ah9BinR9HTtW7K3YSIGOiz+s+jySFb8wVTBTfwp2LiTrwOqm79ujArm0x
hXI+b+42zNjFzHEFKnbtAKXfAHCgCWsmNP4OhvIdfQCrTLrVBnj+VhYVfo8j2X6FtdyU4VgfUjOX
SR2xinvyHHRObioy49JBL1RDtrm8eKkOZzpkAB6bForigydE2wQLe7vdzIxqa+qjAmfocaNyewSw
spEMyxEIBRiAa4DN2ytP1a66MSDJcwpscHOk7R2UYbCyRkxeNYG4qRk229JeC8g9l6zBhSDBrwry
8ARSuf1+jSceuZi8AQXGFNUbGBykblSkJgNDj2NPuywAIjL2WCiEd0vgH2bp8K2fJfIWtUU4LACi
L+ClDIEE6rSt8BnLmxKW9liU/TZ+LNVcqa9Zx5dohGGWyMI8YVp82v0gya+aMINTM/sLDv6wgpSN
1TWi7OASvQRYbWbIP3GJhPyGpUvhbP7TfezRGbDgeRUPTmK4MwYkFPA+HRr4fIs5ybeBt7CfDGZ8
GlsK9QZah5gLNkAAraZlJosxiNyZPfdb8OWCHyocNCJAiGKebHCivb+hTjKVxjgGC2Ec/8cn3E8m
FE4O5u+guSgcBatjzgDWJqK8cm5I96sTnRvQWFevELrT3VbrmaSyG9kb9w/x3itb1fkmSAihWYJi
5bo/j+/iNT9pR0w2/FWaycGxRPETZI5vItdKpAu8Cr0BJcYbSsgzlDBkpWaL1miHbk/wvm/73bj8
ODS6Lbrkx43HKzFEL3aSGGgGxKpN99z2MY0GyvT8TWF3kgNZehAWSzU1h/qYYvkA1gLRyP1FcCxD
pCEMP+mA6Rc7TAJu1ISCn/Ou5gpov6n2MTsWCs3xhAaHCDyUNvcvXdDer1/MhGbU92sslP4VrYFP
VXYnbeiJO66h2exd2pmyF2ylV+1GGljyR8rQBLcSG4iVQ/o93B8vzcAFZFJHu139Jg2Pfxqq3/sT
Cxn6eceZZ6K6lzjnLPbSruTptmt48NQCguD6WFu1W9IgMAD76Fb0kJIRFk5/Fy73xK82IxYGagvw
3+xBoqsSTnVXq10VTcJ1HC+jifwPyGM65s704XXEiL6hKCBBcN4MaHs0lxHTgIt//I1O2SCJma5/
ogQ654Ox/y9iBRdB25NIZ0iFuO1DlQX6m+rrPJHJLD3gDH1SMemva8bH6SeQQDyC74vyoz0DjF/4
ivU4w2hOWSZLMZuCxpXhcrgTakMpBLTLMdpuWX8/LbaYJCPx2glOqHHqiYb+Ro2VByEuhnxjEbxe
OTemqLzHmvV0whdqt3OGsAs8Xpd5VL/0WJJ8yDHc9keUztCO9fOroqvjBq3na4x/Mgt/T4fgDYyA
73ETS06djWDUxqeA0eWy1R+FIDFFXeSnCvq9O7qyiE1y451far1b+QfVqn3lKoaafUVgOjh2uhe6
Gw2HVBlIyuZNlcryWnIaBQl6hMa535RgEw4khX3bJ8Ez8o9JTZ7vB+1BWdG+8Ltyd2z3CBdYCJEb
xs61EgMkBL1hHk0XFbAnYVOL0xFdlSyUxlbWj5/DJcf0IBeLfhKqowkzyBlpu5AjyXYSEQByoQ+x
zG8Un1/RZZsTI4m/+nMSbCCX0x1gKXgYGn/4ZIpTaGJiIr5vpbLCaiXrOhIUvsCcgNGhq7gljyGE
q33qVMtfUP9fz9w0bI0a9/5RNRVmxbXYI3gp1cSVnggIW1ZnsVSKPIarc/JHHfU/GIhm0w87L9GF
sWqKuCEST21s1jGh+aS6E66qBb1ROzBHuGJquz3KzW/0UBg1zKDr1F7eJVS0TyH0rx6DLC3+1tXP
D/lUXjJhU1IxmTBkHUGiwKMBp9fChGtN5TH/+5JFIsQxMPVHACR92z6Y8dnMbkgYh9pxszd5TBrP
O4++i5w5NNloDit8xLnhJJ3JsL1Y24qEWl9/RuNemzdpB1dgfS8CbtKj7mk9/lcLkueeqTJMivLC
Q3lHg4XVk6uH5fOH/xVasPjPxQKPSEEjW+BMDSpC3n6fxztJbVhBIJM0COzmn2KjIULjfdUbRbKK
/8oi0eZsnOWwaDYBUDkojA0FBgKy3TSIBeGQ/5o6fqUgE9lbxyYSIQanC2NrTs2vmZXbRMU5NETS
HYlnzPKhkmE6w7HnE7k3R3qW+LuU9njgkRQ0j7Kwf2xTkAvw+FHebHybyVlGdNln3FUPmiUJY0B9
WzsZ4q3TXHDXbnebne5kIpsqDW/jx5i622M4cQs3LgHOAnVV9eRzfJW9+DNkYGya+9KcAKhwTh6L
vqAjd0AEivodxAdVjdErN942aU1ZFtKhNGcE6+a2PTnlHb+9YphivA0jvl8OccqBeRpCDiXwuboJ
dDNi8Dd7zLawHXogh/3NjgMNf4Q1hUB3Weuk7tTrsbjewYMEaxKBM83f92vsjUvJzvm8dfssKwH4
S9UjWUxd4UJj2TJupcy6ZcaJ7Z9ZdeyMmfuhRF8GnH09TyiZ6iS7KDUnyMhWMjqGpxqHgtDufWR+
KRim8iYB4voi9qs+v8KfDdX1Ojjn4xhgYww5Nf3/vW6o/5bBUDXwMz0TUkgnwxi15SMQ+SSoHejr
rwMch49R9UhWJDjnJkiVOafsCsq4B0LmzZzTSGGW6JGUwoAAUmH7wQM7+n1h1NZgzQ2fZIkvNpt+
+CeVY66BFBO77rLqAHCOs+WFRmJbWDTXmmn4EO66vZh+kdL/9jo5LGThxTEoSqoreFBMXTZIxE3a
JAKRnNfRvI3ESprgaSqkZ7rcszccFMXy/KwLw+HEofHPHZ4pWWmAqkx4UNmctx5TTcSrpF5lHfng
4paqG3g50zJYqfjOOmyOTl8cDOHiZ34XvDJuTNmxIMU+x5fR4IzFq0+ea/w2hmk7N5nqcEyi/7Mk
SDFtkqxySXdvyRy6r8SbsahOyliNI1B/AGuWPqwfNF00o0z5esHUPEvzNl5Sgj3gLVb8bYqWyDuk
lSSj8EDilvLl/BnhIVwPNT0jTvnXCL7Ctv/CxYEBHTU83hDb9j2dRikR47EdVzFs4gzrO78atITS
LzwxV8Ks+VZm8PS1+PbMqNRyQP50RC3uRCl3QmxDi7iIy9p3T/BSckXKlgLyVJvwGp0GLTFwYrLp
zdQPBMLpsyqWSyzM0t27um5h6chgqG1q+vsnXs+O2Q02wIY7ItEz2gVd+nBrRCJSHt/ZOBdHFSZ/
X1E3K5yUOaXv/oI78omjBgk7fBBPPFz4pHm5MHwATZrNQh2sXFKJj9iYNQIk0Bx263JkR6/i1ByL
bTyLP0/LsYWlCSKL+zndZP/93FK4poa3B92oHYrD5/FkginN8ryuZ94SiyEGfvZAiZYzxys+0pg4
lVr7EEWZ3yG7BBUQRrxIBarGULoyyXkr/7iOTGFBmL76sPXL0QRicYgbG3MpkgHypsqapZ8SHO7g
cHWRLwNNjSocfRM/T06WhtqIuQpXyriMyvhRgCntT6V7gao2ed0i5kWKKLulM9sePPK01UIKTWWC
sHfrfwQ0Y3TxPP6r7tLfaaEUsYx2qkQwmZjPlAbMyaoAz/1Zw7YSdMjiWptWLhwpsoxzUcA9IKMg
/jUeYk7uOERjcLJJeLNykmDCpc2pXR5dtNkSHVwkKWOqcd6lV1c6Ao73u1Kkhnk5KVS7CqPG4U3Y
G49DufsXhPvlxGXwQ6r1tjtVZGLYv01OuKSsEJOzGs3JTmJ7pmab+lnCeM+P5inyk3zIFC3IiGTe
j3p4xhA5FV0wrzQwmUABNcvYwq7nv1k4xCPRE3Bc4YG5OovTw597Fs8X+jha3bRbZcx0Jj193S1H
dHA0bkObV4GfKhSiGmJouUHgteWHGGK4g5sGD7dr6Pt+ysLZ+6D9xDhQzN4piGfDI/jxtSlSOc40
/3U0A2v1ltKluhVxLcGEdj3cq+mHbSgeLd+2xt/JobzyEdcwcwuScdO3ZTp/NOry5dw/1dnV24TX
d1Eu7AfcFjVxLley3DKrD86c8QzEQmE5t2Hp5aujt76QLSJYC5Wgkcrj8ORRJ55YlFfiyc4xteMI
6As8jepRu+4tjzIRKTsdepcIWxTN8G/XgmkKftg+zIvWUI9UgbpYFAe2fKLMsRztFpxJQmExZK1Y
BRhPdSMRh02JDzKGg6pKBvplLCK2xdE0SkMdnTCbx0R2ndK+eThEDOWjJXqtk2YddBroLqvV38lM
gM9ilkZHApHhGcfG6Vd2+7hOV0gKrNqQZ+1LVhRqkDllPqghH0Y2TbEwWZmIPg7H/OKST5kcF7je
xLyGY2m37NZOx+/YVwAMudyd4LujizRScr9OskyF65O/NBD3mDm0IhCLA2G3QgC52TiPKr/gDQFE
E40HSSsnW8l2WNoAPQp9meYGq8QdZhOzRNCRrK6hoAHyOBcl3RFwIApAW0qQfoJ89Eap/+ajN/ei
qLsQZmz/m8xd/Ow5i805ajyBUw6Q4vWfDzfe94RBO0v6lCh5KJ6VdK8eCIK0f1c0dlszxGfoAQNh
gMHynC3iHYQZPeJS/FsO3CHw4qDNr6QXH6phIXEqAt6laJfjuyz3GKhFg0nvbKtQUBkAo3hIMuKL
701w/kXRrqvAC+K6f2H7b+IYZ2cMhw0FOQlISxDbkUcADVnSvtB15bul26o6EAqIMpt7E5UNiE5h
PunZ1ZNH79LNxNEPyRUFR6mRE1vDdaPj+jY6IXKLV0LwqczOVS8JpoK6I5LId5ETCeKY5w4wyeBd
eR5IZgJFBR4A7Se1nHWlKRMzqVlfrdP0hdIhkTfJP5RnCTJ35ia5n6n9AxszIK0oc4bQLvcFg2cA
xz95vN8OuwFlWmKeGgwm2AWDK1G47f+uz+cLcgaGb0sflGNKF5qW8YuqGGiHlRb7MX+L1uc23g35
YZ1WZI56WWjOT8C9Ld+m0TPMzkKSsLBWR7yIcXThcT0tnq9hOvlzwnLNSQJDFgWfB/2hNF7uoGOs
xmhxCHNvpH/3kC54BVOYWVjgdzf1DvJ2lodEXD1fFCzaDlgqZVDF41Si5HZrsmCDs+MA3yS5o+6t
ehQe/WxWKcEAx1Y7xvLbVTNRpVQP5pGNA8NJetbnBTcQ+YKjYCixRBqFAB+iG9yx1RKdJSHlOtre
DPp+TDszhYIaMechk7ogSlxGH12IopoTxLPnedzzGDh0VohFW4wUesUl49P8WWtVmtJKghjPFbki
mNAGtTKBU/+Z8uvZksK99/1YTPympRr1C5ZJ+zDh+TBOXM40KFPIKlb3VAqvL/2Nv9dIg68gVWhY
Mxn8SOetWbxyv2S+FmOQP6Fg0jf4X6AfbtG2xtNV8U9d2c3IPXW+0z6QhdPzcy3V1mmO/W0Bq5EJ
DRIKk9IVRoCOO3w6jqOTIwWpIEwk1ymrAXqEyWxZpRou2mR+onjKbB2UX8KrZpcgPVQv6X7fdnCA
b2OEkTj3EfgUnnVuQhJPRGV9JemX9ZKj9yTNSPOrbw2LhX183b6Tx4kcyxl2lyY2//lfzfx7fzm5
fSFoysUXFQmBr5gOH0eikDB9Fai+xsdij1YC23jWTZUlXO1p9E1MvI4e+sOmMUnMzOdjtpkNeJlY
hJPsTKfQB9DtoISA+EvR5rFrCAxsHpwVx5OPPdQhojwf42UnF5cpUWPPUGi7co7Fh39VMyYLlotP
XgdeVH+pmvjPSj0ABBT1LaHfiw/+ccwsLiKlrNqRIl9T45gbQkujXKv5yqaQafq/MkJz/ByhVOWQ
B4040lAJFZ/qqXMTx3bUWgD0incFoGF2E8rkSsN0q7kmI+NpyZoRrOh837y0yLRLk0kaqEEqjcv0
hPMl1Rx/kGIdLO/hEtl8lSUdwE6yOw3+9PKiGlGDOwzOXpepBJNZDCWHrG6ShUPRuTtqSMoaPTjw
npJpdTHCtEuHRSksFD8J7G2yy9RwZV5vD05cZuGLhwzxiF1niFMklw51UYYIHKzmuKfo9j7McWlK
wmaezXwbz+V/hW255ZFHV5eLTl+EjWZ73XN4ziXTCx9E/VTpMihoQGsjge83K7jpRUjDA71l4Wbh
eW3dU8Bj40TnDj4Pum/m3ESe6M9rMpbLkbMAh48ixK0f5Ku1DAw5XiuyMhYFi76HRbxMLn+mUfUZ
xS5jHel8eo/1xUrwYERp5ZhFizQbhHBd1uHlKO3kIHIimCSJuigHH9iUfRZsE2vQH28B11j04I3/
u6j1k0S8QvY1UeEiOHPpTJfhnrLAXmziIihupV76VTSZlD6VZWePveTs6cz+KMePTFU1R42wxQxh
Sr0Xh1dmm67kkpBWwERxi9vgj2MJhMvhxNjzv3ZSDPjbxfvHws7pkMe4t4S+SmFAPL4z67sqrZ94
kb9SoS/ZBDnmMMjmUc1Gip6QJfXkxW2HrYw9zonHnWOqetsyD5i055AFqpa0ja6AWouEpM9MQlYB
QMOiofF0IyiEnUWNKAXzzGdIUWcndVFb3TWfUYxG5Ic9VOUqfXmlEulgaQXZKodB4Zy4N76XJ80D
apV8JxR5CE6q3IojBUj4tWPb0L4hiykFG0D4M2i3gk6HuAuvMv3srsFazYjRLjuvCIdPBJllvVap
g9Y080yIeELeZLmqiZrehy0NelNU8FSnS87SpXnbD6yoCVHj78NB5iW6MttKFR15rfFxyzl9bJNJ
4NN4GOqHdG5QclNxU6S5q0BPSmTiv/ORg3rQA4wePCsDq5xdvwZBZ1ORSuqsRSM2i0m5p3iSCkIS
GOeV2kq1SETlOlKMzIbdVLMVb732bmgy9mD+gDPc6lXGfkeEVbT5xHT0NpHEmijEGzgGolzmnfBZ
uY66jUVjND/IYDhczsQEO6P3E4xDpctO+YMUH+8QmK+ZhadmfopMLji3bDjYRshvK9k+ba/+s/60
O/rRG2L4O5TZGLyAjPVdC1aVuIZrJyE7TrtPGkqWPV6ccB+SRI1udyyjOJh154q2dYo//wATadll
UiRv3a7rqBrxtuynWwffVKKfDXEmgdBbj2dFj7R/yZavSG2Ry2jQaQ7SVagctt3oQdZYYhS++LsG
pk5gD4/ZG27jDc9A2kmT4RS0R2auA4vneIUq63kVxC30B7X4TY58g+7s7hP8gOKzoq5m3vWgTeGc
DwUNSQ+raOqHbQGscDbyauO1TN5CXcQmxDuorTbpXLbeAMP8v+sFdJKfk9CSV1gpY55VHMj1zxmM
if35564dJs9DOrsC1gR0WuG3hV7NMt0d0TOCxyoYgh/hXC+yCqvwl1cVnRRdvbKmbCFv2BpzL2YZ
rLKxQxQkpY7mNLDy3kVFV8rRpgoyZZw3rHEh1cL0HvBQ2io+hmDPbY8FGzGsK/X/os9ec+wtmvZS
6rHnHXLGl9mghUVJI2xsy4O1O8PBU9ret97P2uJYCapjYC5ncgGNQpBBNro2hqqQl5O0/ndYc784
QDYfIeI9zRinGuqy+qazocKp3YT9NmbwJA9o5ZgAVeweM4PO+Bdjkx6yRGh/cl9qsAiaZ1VdKgpI
IL9gx72mKwNny7qhNFgHcBsYDtr4BbkPeCHQR3I8ShhkA52BcgAI2GBUkbr/wq+swrMveqhqiZYU
AAwaGR1gJGDispwdt83RTjWe0HMq9VAZda1tP0viNmCgNLaYz7BcWXTOL3h3ranLyDXwab/XDbkB
RUMMY+xTOxdczHFayGToIttDgFs1bEUhDLA41La0rLk2Ag409OG1HG5wDiKMMYDDNJgVl7TZeD+E
KJGoghhuX38S81C/KE7K8s9KFn3/Q7vpozNUPb6oDDP6y/Or85Sy0/cfsPJRlkKR2OCnoCoAivRU
T9FSPJN9mrFji48tGailhfVp/AzJ0qDaMOYW7rzz9Z+YcXMfXnErplnvmOUiT19BeBqGppJc47nU
xME2gbay20CfOSV8yX6l+aj9OmbUOy7IfdTwOwsGf3GwWjzqK4l79QrqR8BMoqA6epmkuYV6tzOg
vxv+0E5pifAUUgBu0IX+nFz8kr1x8/oxJtTB3ynNsTsCXYCsiPITROOdJd4WBzxzjv+itIXsAPQY
JLQxaY42ofzGIZyljACNTeZAzICFG+B8U5w4oBpLJcCfGOSimkpbc6YKHGRJIo6Z8jhtaU+5m3Gv
ASAIt0QFKIxacw3q4sQf1PgGJCGCUJCMWgL+9y2eWdUVNVnjRs/p2Ja+uVJt/dHlUWU0nPIFWG84
H2ce+a2tHmGdhmD9BKg43fQHChC2VqXqRyq8Xf+I0anxRmI//3OzvqCdWPVb819PQhrsByAG6BGC
q9AQ9VqgEEXwmyu79krwCIeF5bxBgJ2pHmPpG8A3Aiy1CgsA8r0uvhmkWYAwwg93iEqYQJbCIRD1
4sxxSvb5ZtSjWXW0jUB9kIqjXNpnv2w2/dnRcXbsIftdeMq9xiFn0RFxM0tdl9zMKMCI2HQiWyVq
CLiBbcXbBmW+Gu2i0E0vVYA+H6wnhb0fVBbvrD3qprGk1hMZp0B7XZ7hIO9n1kH1ymftv8fyDBpy
T38AatFRn8rFyAMRCdv8LwD6qlMi/vFGDDHsJb78yA3pbURspTi3xAoiMC6pHluUu9GR2laCW+hV
O9PC24bQ9TUpp+nei7EC0+xFd2S4dIwDI7Yq1tIbxMOQnp33a+vBtWnrImAKlDB/ULyAHawpi7Ai
GLVSuWCjTU55+Vv+WUS720FFF8So+hSzkjoiwwE6LZzGddS43rgeiQ03wbYJP+Qr/rYiavccRVSc
pb/uakD/1ZbDUw2w9X43ZE4NcLQsC3+7dDE4FMTg2Y6RZz/JPXhbgkUPOY6+OPex0w5qnjdJInkl
UKILMisJRZ4M4ufB2Aq8w15/yZKbkRh/DgEX3JPmQcMkTFkxbTJ+gNl/g6ZSN9cAPbefv70+5hUM
2907AHIEefIX9wq2rceHxHxje+9SZA2DJHPiGpA0XjzKWq2yhFDxduXeTtXA3oGOyhPBl26ewmmn
AULcrT/gV/swybMHdK1zKBgHT5yhtRLoNWUluCnHpjVP0EoadomsBJsB6HfpsAnOsLeqWX5nOhIX
47lMk6z3ZiUQ1bCDdiZagDqv9FuuZ8elVytw+/dM+H4EQFNuK6ICd6tvaV3y8aU3mwpOhY7lNtAU
R+MMVnQsWodiK0581xZMgBP5+y28T84DIgRfV3eoOEamWiZjfh9Y/9bxqLLUyL6/m3dHunIUs4Yv
lKn8HPhhc7NeUugNx5jFBlvhgLOVQDbgkhS4v2YNwOeeJt6VuA9qxUYEhSJzPGJfu3qQf62Zd2oJ
C6QbrWIR8mEv4C/rnnMgIrrtKipciDZhP2CsVGvHqw06kz5wtaIFiXEZSuZCyQ2T1pzWs5IQNflK
ldeg5LMKyXLkK4ZuTL4rTJqS629EYYNkfXxaAvqyw9bFTnwi5geGP6QuXIwJMDYK2pFYsGUDTLdj
BCWk6+IJCjfLPsv1Oixalbu/hVLDqb4Tp10VjKcVvPSGvrS7LwA3EPrz3y9Ijz7ijvRzKZNXFAlU
2DHCfz5n8kAuXYf33+EK50pQ3VUQqYazjXKTc9VJY8LfxuA6qgMmFscxi3KB3K3jUuaciGS1nuae
9hOuaBRDV6uBmuCSkGsK4KXCqjkYKz5TMXBrX9DClK+dJM04OLWGXBpuvW0K28mguAV/SE1CQ/5u
6S7B3jlhUTYe/bDbI5c4JGr+6flzN1Ege79vWj1tqLI8+Cip43rhctA7HU0qxxAzCK25cTeEpP/M
7bZ/cHy7lKs0uW17sLe5R5XrZ+MmsbbksxxPWfLdht8afkhmxeqCbUbWhnPMWCtxGW7ieLM+jM2E
fV1uyAsijmJZMsOv9I5eGbzf0lQDNk0uaJbzITJuDVeDVhDnQ5li3ZqfrgxxXkdfaLpoKPTUqyLj
SOyWBlRiZ/v2tUAv96lTtBsgLbY2ZAw7koKZnd1iUtW4xuK/bYIlf9R8ACNJacHF9fXYLJotM0Qx
J9DdVnr6HwtFtZ6UqxnLRK6WxutSaWAelmavt7ZvH1xje4vJf5kDh+u8p3zMp23g242znptljsVC
KTApzdYkfDJ3LakMADyhS+cLehAlh/MbL66M8uvjTxsXvipnXgdzixLlu1oH3oBdTbLy/c2qSWKT
+s6xU3l3U+skHI9mRO1h+PGibFwb4vclty/d6lJ6j9/EXKTxKuuRfLdwTjn43UycRLaCGM0ZghBQ
RnHbjXXQEUrI3Kqy0YcDCzhUl6xaixmNNrvO9oDPCcxNweVQtqRg727WxOfe2ZMNc+XlbpNoMNwp
EhmP5v2NZ2kxgWG27DveH/1Hlvl/cUk8IGWx8xTMQ0IuHRjaLuLtWaXqEUcAKUUK40Z+yfo/ipNr
AW+AYdwomNfX0d+Uy9YNHGbDLZ7/mY7BSJY0dz7gqpJvH2ZwmYonr/f2GCYDJO588eIBa/mV7xpQ
kJmd5U0YGXzdPs2QJGyGOBGu/k97BRPe3UETDM5caKGAgCX7BOaQuBIU13oamY2aM9VrgAn8fDFF
j8zuFcF8VCWOTLUm7K0xv/glqTV960AbG4szJBtRVAcalhJwQaPgQxUU/wIUnCmTKmVJlPlfRmH4
W89mYChW9LNL8apZurGA07AP2cXvmG+vCLZ8yB8HzTzYW8SXEJyx0lKK5Dl5svEdtr9IEiHqP3yk
hx8CpG3rSe9kN25Kba09xITGDXcgglR7JAQ9TRS1N5UjNTsABhZr5glpBPDmlH5vi4/qRKbnyLIt
QTm/uYjK1uXU0Exi6HWHzXl0ThwORRy/F/rJbpiJBY7mmvkYt7c/B1h3If4VCktXQ8KPIbRy64jm
54NZm8meuwoxOWqEz+eb8vNlUPKEOWGJVDkX2uccaSw2LalrG12He1cpvwOWtpC/MEGk/FtF7QWz
+oH25q1JRdmIZED045NxAcREXbquhGPcm82xZm53F0fCSaadgpw1aXQar2fcfcX3h8bGscw91lE1
Jq/1+EZUtNoatFo3OIXSnFtECvNbhoc2ZcwGkTvKXT9StqX9zqnN/WBJSjmu4Wz8MXJ6h/4MuMNx
XBmkA/ZKii1ccIHinBjWCK2Ij3+kr1RD+TfdrHEl1xvIbl2VTgSo0gjjqJsUsuZNK9LCJQwQIeGc
EQJppvlXXih/zEbLRBzMLKvwzWXHfJkqzqDVsJKWWnvHkVNaOBgoVTXU+1BXYFr0/YX+5h6Ui4Hk
qz9DzHF/ehejq/goxBtyPee6hPkw3wchUY49oUkKFsrgN89VtS8MEZ06Y/8BdeioRsKefrt9a1LB
pQPo0F01b70yD0r4jrkbVwgDa5P5Xw13LeIFLrmA2OeFIblRLZmMHG/omiEC8P/vg4WK53Pj7W0M
Qcj3ORGS0Ocy7/C3D189CBJP2UgiyFAETGdMPXaUEd12Jzonc746Q/UeKjUx5baZbIQh7UbCuntH
bCd6gWfKVVMF2W2L69imZbEUGDzt8Ge5kOKWcnOa6cu+99Z2Z17/y4voqkLR1MaFNqZRDvVkejwe
2/S0IhVg8pXQ+ntERkBuh2Yohjxd5plr9vGNcKxmRtRswFcHUnmKRgk0HVtaTBQ0AjN/UpRbQuVH
kYg1B/pvKNa6nZ1qqmztrA5qofK+9jQO/DYfJ8D+EyErvYRqTUIXYr8+inHCVxAcW/Yrgi/OV828
ookdLX8eK5a5sN8QxvfEuEs2+mPP4ajqNZ9IPg7mZCk30MDzvxDwQW3bxWtKBvC2pawHIXx3dZhI
RH0/lZ5YZHqdBkqIQYSBqzYG10gjw/GeMvfMR+ChDMDJKntfGvabK3FuE4nxO3UlDIjwSoEqlxax
PZPMJ1tfT9o/7BXFDRO2ECw3Ycu55xGCpUayBVg72wmF0gCpElt9zvXOs1VRkZheTDxpinyZcfau
l5gmD2Xwln/KMAo6wZzylW7y+YCf0xPqDaZEZy0v9/unWFugxVGk4lZ8QcjdYD0rs6uUA5SxWfq9
upY9D6zN6+z6VDwydpw/Q+Sh7RXR4JPsc6B8naW7bCrYYWjzDrKjIDe/ur0m8VWMl+SnH4o4Rrim
pw9QZH0BMTd66KwMTShqKL8We4aQUhvno2J208sJs0kgzzlNW9VXnDfhIZgLJrK1B5qsRLfa9cun
DtI5x0wOYCrYKvNEydiRyQDkux7zQByGCN4o2Qpue2Ji2T8afsoAptzKbshBS3ZnkpZnBXlS0q+y
mijhfFhP2WGk3WS6Nqf6YvF1pG0ZD80F6NoSKMkxKEupinDWBsc7QCRFz9CaKhOmxoRNGuo71/lO
b9+wanxPMnIWoMHQtrnJUkz67TbxMV+QcYtWSzHUjakLnyc/EM0po3EdynhCRBgEYFqPzNFF1T6G
jNwD3tYUNk0kreDtn8HY5sBnL0uEfcUVFGv3lmzIUz5bniad0hvrbYAt9oYc8ZIk/fg8EDlpA53l
O1NIKndvq7mWEvL8XY5If0a7WnQtZRBLQht3R7aCLD+rPk1WZT81AAhKxxHYbllrxEqa29CjT3iE
khf0RqgriF0ahFk6vwFLhXZTYo9xkwMw67dV5ahpyYzJOcGhR7ekRZ144z2ZHC6MLbGyM/Ws+uII
NKol85ge+FQY2nqMdGh6xFzhIL40jDoAbzFgbBNoPib5BPWhUg+v1eXrzPTXfIU39Q6+X/zkpSdT
7Us7JCFuQ17P3wsXl8i11AReTYteY/rUwl2VyCcoUffex2ZLyxSHemSjbPDBJuzIbmaOMmuj0S88
ioZG/mwzb9gDUVRBF79Bqb95KjNeSuSprrhV0lmQhM4FMXzaZFlL4SIBRWCGGHjWfjK/v+eI5CPz
9wwHdjZUl5A3yQon83b46K4k18Spb5p8Ei3Nm+RevX1eJgEGo46ZXv5GtzyYl9JZSWCFlWSpoPzA
t1lCaJKSiArIGyMDizNIO/c2N7DBCjbB3i80ZV4P2z+J65WHgikcY1sUZjYvree194dYliESncYp
hOEtnQqxikXoVZCYvj4b12L09YPa+9E+eGM3No5pWLX8ZJU7xRue6/fbcAFnIB25QD3euUNtr5BF
kHZzdNsxsTeTS3py4rTIw7wzyeTQw9aWgdf0V2dFquCX7t0gmyyut+9M0kpTpiPx5hg2RKVa+eMh
D948AI8oBNAI7lJqClVZ0wfRUuHeb7VAq+AaTt7BxlgiQUI29qnbvv5MQcZVluHf+D388yUjP8FE
+pirpjtkdS+MS2VVtgx08SbWi/1jBLV3g050rbf/MkEnr666EIMzU9zrHR3TViaZWIpeH3zH08io
a89p/j5m12wSwBL8LHauyRMS9cAowg+CKBQoDPSillU1sEGjD8mQT2XcLL/Oy8rol2QBLZKwBsBt
GHNQPeACocUI3txsX36Ns/pJ4LzFM7MqHOxtX7J9wstOvn+iPdaCcaqJCSH/G0R5AwY1AQcCT3RU
GoU3y6jls+scoYheKxDFwlgD/SrwD+IXaZdw3MQ948Y8X9Ro5d+85ELbe91bkDQTtuceiUeiGwfK
oKMGn0fjSl9sHYOByS9howSOqFmAF1mXVQZ4YcLakhtFb9OisnJMXx0yB4aW1WVEYx4jBv6GXfL4
QTti/N5qXjnJMpv+wGkacrVvqKMJ8iDBfTeLVI1Ip1yx4d1jDKB5PeqHX+Bq/mqLtKwDjkqdZwAt
+JDtzD012BGz4o4j8M2QLjYFmLgMR3JGarAPm1hIOoplAPeokgEXf6NPJwSiv7LpiMuUPj3LGPM6
nBAgK59IR1EBYCA+YTPPQY8haj9qk+WIXYKivXFUp2CpGQS0Bx5eW1KGE3AaAq1g8hO+37X9LxyM
A7OFqYRASEFshivY9kWrMhaMoBcE5aqVy1sYlGByxWtxhA74CtI3P0OUaMX6hruUjxSGwNqbgZ8C
nIZmFgF3pJSLjIXYGAlzjyi0wvDiHlsSm+a5toUU15GyvnhyRQIkcU4fZjUE1oaV7+TJDS6O7Kny
8OT4CrgjxNmvB/h88mZFMAa0XhsU2rYtY1vShbIwYT+xytYKHlwQaONso3o2sLtkco9CHfGzEPyP
OwJjMBIhdDCFEI83Hd3+LgSgU9ES3kyqO7wTpWCeOgXulWJJr4ec/mDPIui132cUxukPcOVHs191
TGvaJ5mNLxlMYTHwvVVWYd0Pq3run1rii6scDnm3ZeBGmqNqkLFFk6MX1c/35IG3MbjGjwpvNAhm
Txhp8jGmS3ZBIewsr6Je++jhJHlFnU6Ojfb5cg+qxsd8HZnuJAplDKsQL6mntLmzvMtcQWlIqpCT
R2KOeLXGQ2sNm8M5PJljU/Wuj1cA/eBDDYSSlMumyMiMHuRY53p6WGXbk1E7XIJ8P93wamY3doqD
8H5LHWZIXCp9N0oMLBW6cVkuelfgOrQs4UTR9bnvlCZPf4sPUV/zZbIFzy2xlcBFw6NFqtbTq8sw
FcfVzvm6C8B0ClkWlDzfoMgBBEFkZ2zpO/7J/hFonwL8pEi2UsJtcv+97wlPsNs8scB+t3IcDYOW
aFUAAPA3cWIvvGFt2twOgBZvS6RpzVY+TLIiRBewnlHECu2hoWmnT2O1p1rOptyJGgUehdiKSdx+
M+9oltX/WhTmSq28t3X/TKPGBEZeFcYPAGwZQwD+mEE2I5jWmS+G39BPYjiMJyStHl6bm5aWyu87
GSXJEbXbwgMDF1tK2r3CPSF2RrVQAagemh7KLFFLwKg+9x44ZWkxdLRVTdbqJIdyt7dL7qQaP7OS
cKtRr2ngBiBezaad9xqYXsQtRX+9WaArQoCo2mGObWgPnOnkwUKXXfNCLt2/m8Oi29hr7m0SNk3C
YpK7aRfAzxy2m7V/bwaJ3qb9gK2ZwZ8I1BRlsTtINfRXaL2KezHIEBaQmO6PhB69VKLRT/EMsVvb
eTMsd+q9sIKXHw+x2qtCInOJkmTinjvFh39BWpg3OvG9Ci795Z5yVUvIk+ux0Bqunx6HyBvbKrR0
S/2TLAbWjzsMc4j659rWhyWGeBMJnUOB7FXfVchaecntJA+saAWkvE4tvSkaQ96UsoHfWi20DyVA
7QGpYjcxX9UyDvVhMlDGsAKsOQ5Igor5x0qz0JztYuFktVmdijlgsmDxfZQsHS4VWNQZ37auUs8x
hxsDPtl9wXVN3hMPN8GZmm81F962ho/FWpRF6D6Lxq5HnzTAizxfftSUIMBbuwG4XJsoMk4shRnm
eHPNF/sRNR03zzS8bRohTC2jYxcG4tSfzbEKJXVB3jPaTJ/7hPi4z43jSd3ZEOvb47HRQ4y095lk
WpUz5IO9NvWplW4qgL1BhcHd88Zlx5GOftcja1iVQhsHk3tsUi7LPgp2bYLkSWH6qbpiTzp9F6pQ
pM6ITa0+aisX2xjOxuR1tzywzQsaz3uqr/u4VwGWPghf3R147arvZBAMswOZa3vMwEYNKUhMmTDR
NrNfh3UuO5rTvniJJXoqy4a1DpqNYQEbVukdPlN5JOO+Kqy2FS5/ssEJY3bW8QffQ/Ls9qAAhsys
jz+CFABRpvE3x8A7x+JlWL83Wk/ibokOKjJmqr+C2mzfBmIcRu6JvEGWEPL0BLUOPxlXUoQsVesO
VjiRk2ELY/yIsg+07gx7q6al3ZibNMjCBJBZqebTYSvdiNz+K78JHu4T1d+/5BC0tzAKEqfNwevj
l6HInHMUBpWEADAxZC9AJ+umtMiX428KGiR8i9c4cW+Wd2cv0EROhslLahLVzelXSBNJmEHhhnCR
tHZwQxy51K15zSMBa2CAFWoWEaWwuw0Hh9YA8hJTz98+Q7ttUc4+ymyh476niZo1uGtCfgzq1f6m
frnenPUJowT9bYCE2Z6XcrxerTExHJ6jkVyBDfeMGAdcVOp/NKj75hqr91Z411v9s2RMdq/hTeNo
PHaJHqiEINanEmdt/1McfQ2rcurcuOG5ui/d5MbnurdOf78tbR4dredkVlmk3ik6Ij+Pi5iPK61P
untv3x8vgXEOtgqf0eJ+Rm//JS7tM/IliQs5nHNcYKMShJii1zpSt9fBwLZ3137vjhqZ/uJvf6F8
oHP3rhHlSXd95FkZcXDnMn6Rwi8MgBsU2gf3/oWjcWB50VuIOCSIFhYlLn7dt4H4YU6gktGwm3T7
qE0Blrb4qWOehUOEbE9meQbfulAiiS2MZ8fPwQTkWSQOs/UkO0kwAUNq5xYF/OxPV0tMpXztTkmD
mhhNwsEXx3+ACfb1gLOaeZ241m4+PkJQI5nYMg0DdKJEAjEq7KjLt27/Dz07+P807F4CUDsRTvwg
p5FfZoJjXi/fb2TtVDkilX+tXrFJapI3myzh+Sh2F9Hk+YEz9TfzenP3vwVI+OxbBVQ7iAKTmSvC
LW2zggTJ0YS7HGBHnQm3IomTzyMfuoxitcnMpTn2/g7KvVq70PI9VjL0SQqOpzPyPNRUgwckcLQ3
gEofJmrsP5vwZo9zptjgoh+B/Z3tXz2Ba5ZgV5C+QaHiLw6pZeOCo+wssw8AxKOg5ulFpVAAIZiO
sU4a3aFYL6ZZvXjbYPhQLXDyejbwFf93z8SHZlHccy9Y7ttc1pWKQnZD8tw+TUy/ykoKFTeUYutb
JZ53pdaHRHubYtKpJAG2ztivJoEWYmr8y7KI0MBZf59aRWiE8vhZTCG2GnOpIPX84odUXfU8VaHK
6QHXfLAMj2ptJojF2WOC4jQMf8EW3NQqhxb6h7OWyrUdfeVsB3l6YxTIfFdVI1T/KWxdqWy7h9bH
247ulpyvt9ntJEHKUdGv26yRb5aoHNb6bp+w9aY4ODXNTNCwDpEfnBlvZNE3oxi0ePWkBh8rjfbc
QcxpC5bP4R/Un3lRMcCFW1IVDwFsl3IKDy2xDvj2xJ+/xR3973RUplj9SKZ2oaszYDPtWOI/yROE
mLSRYYdKmWmUBcs1eC5nsuxncRM7qwelMBbmyGU5IVCJwnejmR5bJOQSpQyjfdjqhsMtKPmhUzkL
GZvm5Gu13Xs9JQt70fKO0nXGEGHFvNMPvkItixtfzQxhQz6JS2Y/RDC153k5zhYkzycPQbFy1krJ
qghKRijaOKE/vKtCz/EoT4PAjbMDk/n0cB6rYN9qUgyoWgEP0K6iDysDSX1VKVq/MZg1OvaabL+7
yGtiucaAS0Tzvk7ltPYyhokknMRmnA98RAkUrkrAOCyTwSevXHK3zdjDQJFOYbCphKZ/wov/rJgf
Gsg57pT3v2kk+rCsHUi2mID1WtI/uDh2hixQzsViH8AfPemGHF9VQCHWglECgT0dsrlLsLxC87lU
eD9F2mQhZz+YfCThYNICK4Gy111BEm/UnUQoqkspFZ10GgTqLt/j0K3AXVzCEcy9UvFtEXth17TH
FzF8aLGWlKJAxFZmoXin/KZqOSm1lokw5i2Uk7ZcuShPXsVy+nyJ+FgYOHGda3L6JeOu3A9glTDu
BFcdu8QILpIMxE7ZlYVrxCIWs7I8zwXw6TJGNOyR3CDqyAvm+ynGfasOhCSJuUrW5PEYcv0AK5Ii
A9QG1hMJMPFaOlykHcnSZ9nuXzfKyglMnqEOXqy75PM3bTnkUt8j06sCX7e6K3UwSKpEv4k7d/Kp
+POJgRDs+VzR9EzPXb7NvzzPINJC+T3ErJQdWR0ujIYGI23HBRMnM/L17XuM9gLpqrWjK3Ud/YTu
Z6cgikXQitTqrqE9fvluKXsmAreDWiqBkKS+cTEX4IhoDbCZUXMPzVsolGuB5m0VMSyQfMa+3Ihi
lO0ZNXNym5JrfRmZRtzQgJzGy/vw+p2cmR/QuB5JNUHR/xDWDZITrLxrYdS+nDektVIZty+zlTgH
hHo1R++tAM9IcZaGFGxSd/kPQHZUeaS6fA/JCuARxjld+UMJPM0+LzBvTXCSVZkqXuisH/cpofRs
2gWipyzS1M0fEBnC7HSUwLlXsWs78mmmpEAiZKDAL30NV21BzYSd8F9RuxppouxJroxW3JiE83u4
o4Md9IUV3eiIGrBN9my4ibKfsjcuMOCMzv5pGxZSF52lghbt2+HD7G6rPkCGENoxmH2/6sHYz4lc
cMg+EGhV76e4RDhPV5H7MSbdEDCRIgy9ep092wQhAu9lmNU6yMGlhftGszmt1F/MjTDt2U+/HoAl
5/pA3oxGSMxvsrTsdPZ0OZzvFHaJw8p9imRJw4W1ck05iXZSEuRBNFHDTzlkwSrT4OM3tuoHezIZ
fk2sM6fi+ki7AvqI/NBfXidPCKJNYtJdJ3qDGuc1Ukpetid99BgvmBYV3iGYONCmJ9Xl1ObZAPf5
296evC+E6z79ooRDJxULBA5cfpM2EFZlHuVajgYdgJ98cM6FISqic4w9KSvEhUJO07AziBOpfY/o
ZgBxUCCwpE7TWjtE8e3awJFji3WptUVn6DsZXRCOGzjQCaEn/L6UF6zShnfMZkJy9COSZS7RkLrc
Lzh3mJD4toHywP6VTS5nCyzkeb+4BvCvOjaHB4HKj+EBylEurFVxHveLdHwBg0UNiTNCbYLTzGAb
NKs0b2HNjKQUkolD7gRLdSaGvMeyFZA2n9J4kRgjlw6D9QZSx26RUhi0yqsxwnE0/LQK3ZuMgXIM
nsHGBGA9CntG5MGkiVjDsvWWPpL7aX5OgyO60sJZ3cgSL9ew/vLhhuod04eBvvwh/KZJR/8Zi3c6
asJdV5xt42t4iTnmeYB592KdiXxcgeMTGSVCs9UO2m+IHlwWLCMe2zSczLrmHsidgJ6/FpCi4v85
cBwQ/BnyDzkINXYPjbAMMsQucLWTwUPjW0Rn7tQzB9OYny+UjLGrcVn0qAkZAwddV8XOukfEs5Fv
bDci7OeLmteH5Bvjf5tSuxvVBwJFKKOO10NJsnfjVEGxYcxnPyhVS9Giopfzsv0u0r2rCc4gAYhU
HHXdBP08Gy2gcCjFudSdl/bdj7dQWjHnrtDUhA1RRTcLDmR5RTXWou11DGH6ovtIL97d+9/6lnOV
tPholYqWyEcpKglTpaOrRh9k2OmAKz/SCIvqDp32ut0/iycDzKD2mY7d9Chq8x0JQj+EyADZvJ9h
HaV+b2FNGwXzQjJFIOy4qaG2WZMJSQVMsWBgzEdf2tStwNAOawUsloiGhi4mg2LOdjmK7RkEB+bL
i55GJRyC3DMP51yEluY17eE73H3ItApOwtinkBUFfGSkW+aJE64EtvKD5uiMfpbDrrV/Lp+zlkkb
Aq2GL1k04ujZ1+plLVqUFb23h0qs+quAB4v4j7Af3ZALpFFS1+TJcl7y/jHDgzFtqnbpahFFnt/2
oRZ7wVikAszwrNd0F/1CQ3uzGhmKFIUI6WyqFjC8tde0/7fcKfCWskpcrSSULs9pdub4l1DHCW1z
6tMukbuCpI2dREn5NouVFDBQatSj60eyENjwIblpZvFd5mfndN2Dj3ZAyYvuqa/kfcxHRYMr7far
5zeEZUOAQJFjOq7c6TXjTxu3QsUHAnYr0mSjZxUN84HCyy2X16EwYPIdDllodMUexr3Oydh3N9zG
4v+8MimU5nPTKBzhMW3HGmmTmb4ulmVzeNtM/zdnae2IhiY7DJlR3d08qHTfxKXUrBjHs7wzDHCu
JKkiUrT7P5W0x133kmm12ASxxfUXL01RyyHetRtp3mRpHYJi5HueSk2JDVI/lXyFo+tyFwWD9Hyh
5wzESQnJ/oL4DBd7bW3mRXRIzeADx7cPbIQKYm8xPchrMJBUKtMcSmL53hZbWGJdsOQaaaqGbNdO
IZSIAKyFTt+MWeOQiO3bMwuPuAfEfRwDFQW+oF9SlOrluTAJNh90UxmPChtB+KPVeroX2nFNcy2E
GWOxkzyvGatAA4L9EZp+gUO9yMmidw4YhB10xIrExPTMuFXZtQDw+qMfIxvJJEuFbEx5+NniZwys
91G7FeT0pM+a3RlDlPjoNwh+9rS20CrBBX88ChcQ5Qo/1rQbdEyFODfUcZ4zURy84TGIdDCSXUOo
eO5qNo3gHvB2ypvJkFtnzXlNM7Ipzaq+KRjqKDCDAn0GTOYlb26k8oxjBdxdlxHdHhGe4WHYK4iB
rsb8p92KP+A1zf8uhucQD4mVc+j5FHtI+uDiWR1VQp9M2KXncpzKPG668tquJGlKyt5x7afqy987
3vukPpbUPmHjbbdAaxV/MHa1ADRPJJhVvtT7VeKzJ0HJOwaJXvNYiIn1WzgOLZzSUipwaMsmGYZP
jWF4Lw0uwYtzjJC9mchJjmWxdQM3ds5QYUWZRsIU4Lbam3l0IqVelpe1qRX/3IMM6NfaOLbca0kt
0+3A3nO26okRG8AxjXk5JcNM+U5APN6EP/4cCyxpfOTouT6MwPfROvVfp7ayNZxJcGodJ27RCSXb
S6U6WbTdRQRS6w8obO7M0vjLi8g6yh5SL4c0AqEXpxFpDr/P+O6zq5nwi7RhPOApepMkLJvWRBkX
qkIEuU4Q/J27XPBLe3mwPWjModvwh93F7+nCZjg+bbia5X/k+XYGxKgGKR46hSP8Nghlhs6dVms3
br3jHGdDUEPFA8FcqgWYHkonDWUh+Ac6hc1NVLboD1Dpn9Yx9pN+gwnd4RefL7Nv+wWanvbaimN3
QPbt7xv5x/muqGM2jcOVxoHQrIiMnUG7BulUvh+FoGSE/6yiV36GXoXSYzHOM4CcLPD7iMsCAxof
BqjphT3o6gQXlP1TT01BT0BhJbesF4fFU6UfyomAYl5DZsGyR6hBqzcC+tPRuRo10ufLF6aqrdJl
miGQuvbJjbSSruPCUKI2eGPTyagrCW0GWhZgGmF+kTityIaWmUVA2zqT8jzmUtI6X/SXH2LfUqZ4
gH3hQgq/7Vw38JlwfiFbCEON6rOIgh70aje+6W6EFZerMZZBXm7vpo+B8Gc5emVrAyd8gJtTBNuM
HjGPtgEpSRR6xhjfF4dwHHiQAjEtjv0fUX/wxO9EGW6X/2CA/dP3QKokaNlgmrQ8Ix9ZA8n6sFVz
V5kWYdl0JHpMUt/Ewkz9wTIp5gvGqogwkludJmRELLvWpQXg2y3da5sCFzAFAV7m35Yx6i2PqO9c
cqD0pRWYaq3wIpT8kQytjQ6CSbNt0Sfw2I4ceZw1ldfSmC18KKP7eFn7sXv9JHaZB7frrRaiGdZw
vZcTf6h+WMwslSfotLDn6ySwkDEJOMCOUaxn+VKUb6a7oY6ZR+Y9myjln9Z9RsEJNpgTh7/Fgtvs
Guhj/EqdLwWOi6K+M2+42/BofYIbGZlJtXkbLoyz1js9gPszqHujvkqzx7ndmIydXgWvv+iaova6
EZBTHNajjSnwJ9z763XbTDCuDQWvQpjzpIT+vUrT+qniXDxuzurcv6b09I4eJ16O0+mPFUlRB+c4
vGNq02RrXCOHSEXGmvKSHAkk6JSmr2uq3znAaDlftAMzqjQCOME96GjcI2eXSgRdZMH4x5e0jRKY
SNuZFwoT1lAdfmcZrkYEyUR/Jjo1CKaJlXEhTef58WNR4ocFyui26NNTzIRbWssBuXR3+TQkny2B
O6sRA5n9XAjJ8VDPGYdTC2tIG8sRgcXAs3Wr9BzjDb8oL0n1Pcgk/0QsIlMW+sMdRIANijKpCpdD
3dJIQ3W2pO7sFFK8hG0PQNxnc67hG8c6PHry9uyTyR793Sm7AGkn3SRwSHr/EzEDqnCbcf4BzUoK
xAeWfhzImP++RbeMLOiop4/NipcqcW07Ec3OJT/7zlbbA2yyJKdhgEjvM9oH2IaAEn2t7tuXmx3u
E+vIopPimsuVG3BqjpEJzu+R+dej8MhbULVpt2B85XvEEKpSVQ22FSOdA4eBKarcxstslyBudnqU
tksz9hVhF03Fix3whwRmYHjkRKOBQUijl5f4EDAuztcb+2HZ8FaOiVqLLI2kume9je3x3RPMQUIV
fdxTeMeUtcb3vF5V5d0OiKx5M4geS6SGmHPXSACbOnF/HwiYzOcnrciMSQL+UjwX7VBi5wTjnHaH
sl/LC/ps3fq2Yuezkr3SkNgLcsAz641hDudatNP3qXkr9/iMQDY2jvg29kKTlUgsGgHLqcj2+hOg
xWrSGn8GW0r+q8NNHwp+B4Xdx/7NEgfKQE+c63sbo7jnbCDsGsHtD/UiweaxnpmSi/uCjOoPlHNw
ikeybZckY1Al4/ziylTkCfnSX2UAnTuzJQKXQ2/S1e0tz6emKY1nWUDlglZu0jg2vpN8qZqYYIda
cypZ+dyJwFRUq+eXWkyk211atAVim15eUJf8AXk/UgfwRgSHMkyqN/l1Bj5dPB+uRzZl7e3i7M8o
p9/2FxjtbxLRocEjE2p/hOiQHCW2GhUJsAd9u5Xu8gFACykegSBQvkWp8KO0YCUSj7rzwYKwesSD
3PIMrB8RAZV1V/4YjVVhBO49323uBcZp69AoJy4u9lbDSukF0JsQIQDjZhQbvANCDbYb+Swd0Wcu
xQ5f9Dv0HGgUrnAJyxKQtmV6kjdo1gVnbiwx0wdx3sXq5NijEQnmYt8KHUxghzLacxRO4wFtWi6O
ofEEb/Jtd9VsSzLDLr8HKKFv156I90Q4Fe0zSq4Vn6dg2IfgrnW/JZF2xTwsFT/vUvV94rHpW6cx
L6+pqu572aXGmedhk/qZTzcWTfGXnpNcTC3KQYOLqpimYbXEU0o7YYzTfKck+tl4wIimQTChNrkc
IndfthiTBPbEXZ+L4Kxs+O8yPDo/t7COnNMjje7iqzfDX98dco1e+fdqITEWohBXl2hJIKFDM0jV
tynnQEPtaO7l72IidaQB9A1PoQ3iSklTXyzrEygPvo8Hjr2RyNvkR23GijdjJBeIvnVP/uOqc/hm
vzfb6oee0+VsBcGsuLKHqBhkNw3a+n0iykTheyOnJeoPXZ1+PzOb9Q0lXb5Lz0QslXjBCpekAbZJ
AkT5gcB2wNpCuN3T7IEEw+QscYDUnfL/lBFFdrhc3wR4KQ67tuSstYiaQ3vJBE4QAjQRGSrM2uwH
sDCxsdI56GGLzjyCalI+aL6/Xtdn2Z9pzibPIOIAxJS5zsZPTpcqKwoDzPwEQkfyrM4ES0fFeaS2
qW4/Zd0c3d6jynE7eFEQYIg53Q+SC5vLfTEFRiSsmXzELY1fHhZ6aYrWWJjtw5NE5M4G2ChL81FK
Akk+y3ht0J4WxVREcMjQBdh2MNweae4GaRFwHlMwAS+B2WrBFZRxxVhcLGLZgJnbVn2rfxRJaIhw
1lfsOdVilDxxhGM3r19hhkAIEFNEgHwcM3XTdxEkl1RmL9gas5oGX1q6y/qUGyEg8mpbs/l0uVCF
+hKKFyuUUSRNGctaVjvCvrV0+09eJf/vFw6OZc0KKmH8f50NRJRblHvxmLgYPScXXY8pXupgImyJ
uCSiAZvKNNudC1uVPeomJDGrpEDjeCSgntkICvdd83TitKDHQvLwZxwXbin86W5poSDHpmx69xd3
8BG5DzcYJYmVBRCCBG42ilV08Ip5W66NS8U7Q0S3bGEiC3gpajBlAbSoZ60/76+MzTc88YABl4j2
sGAMw3UquFvFjLAPXFET2zB08OecGyjflUJBvUVOyBVFVxnCv/y5c3cn/PWQAZG2Co5goeopUt+P
fJ/CRs/HQh9BmFIhBTUoKRr5bU9n0fCbGalr14z0cBJL+a1KIJ6i5l5PheSs/gpjIlqyrbfC6TzB
3XIsZfBh58y1nTJW/HCJZ5d2gFldZVQ9qzABbFMz58GCGQBtvU9zmkDUYSis6/VF2WG/rGJLmO7E
24FrCf7M3myYKoeaaJf4IfEgCUiRGYUnWhl57dEousjBC/mu51n5oKaBR+bxX/fj2ytCCgHpGslp
STAcJ9w7WPebn15OSgr34q9AfXkiJmrAwvqBXq/Ep/m+0GorugPgJ3GORJMaXgPk9xVkXaYSQwKS
MDha050aVeR4DmUuOF3XxHZDAdPYrgWDyTnvcEHDKY9sfObVCjFRkOHwx3o7iSq9E84jawD7W62a
IAFUPtLYNbT/ZGN4prna+koXdjSgGDwnUW/2Y4f0dZ6SfJ9yanqCpCibVTCVLzapiL1HX6wvOJF5
sNZztIfgVhQOv+hvpSEZaWtCQPHW3Qs2hDF41ZQdFXLwkgjtMXMKelMYCtU4nB0si9gQNgZRLAzT
Xh8ZAAqpXOnW4cbZkO0Q+aMR59MYqT7SyfUquMvrJ5qrD3myWqn57rHEkJ5GTubNNzSsnnZY2Jlv
uXvb8VskS8GRXvda2dsg0zAoedeurYe9+tFJNuSzIBYSwlYu0cCQmfBUIHxCcZIyN4VrztvIaJMp
VkpvQkPU+gl5FDS8abS3RkHiz++obM9mF2FY3MSq82rrpui0LCBG4JV1LfdCpkKB2bNfxExqH6rl
Wk1wex2oU0aYfdqIuxk8W9fRGmYMwW+zxkCAcEoi+ftLkROncgh/4GnUezJWvpdcD+KbuGaA0qND
+C4Umgte7glDM6oSn6qGM3Dk5oUbv9kNWjkf3AGMQFthMkrlS8llC/DYgYYmurcy+aytkRjc5V9T
OOZTY+noCMB0apV1+2CLPAWkueeyh66iMFKj1EgX7Rscu6u1aC/aNNdy9cbFs8Bk/j2GOX5MC/Cw
BSHS+XJrILVxdlKpjBGVjdSxAlfGT3W+qMS+jVUkohsKj9PJWNIhji2S+en8aP69p4OQZqZF7ZQz
gOqlFttsTdWMnocUPF1FSq4VzDGMyU4s1LRAXdSenmw68MIQE/oOD2z2tEi1dTWCBzh1s+zUfBOH
1zv2nR5kKM/cjOZNRJnsq/CbT8X+mhOhouhHAStvRRQM4E8qCiJ+4ENJDl2JtDabHIkDp94rEE1H
enJrvbzHSgCDprIrKtDoEbvHC/lofAl/c0qpiRDx9Lx24ex3ZT7ksl/H2z+dNxNHNdQlCil4uAdW
gJ0TBTizmrw++F/IRTxrONrWOErFU7v3HWZYPHuCtSw6hTM7DAS97oUuONqzURZfhTlzZYpp+ypN
bw2nwdr4YllS4k1GsCSgPxKQntPOZOwreT4pT/FaVcnffrRnk/DAM822KmglGwQwtoTKmAQumJlJ
YV8yR8qPIIpIAv7v9SZ3yZHW2bJOo4f5QFXUtYz4A+7aSlXCjv2fC444cPf0UjU3/2t8PyeoaXQ8
cmOJbJNBOy8Pl4BNKLlMdN/xBwiiUOKOf3aqdE/wIZQ1oXfr+tluzFc+qFmLnbyrLhksKWELgDVi
IiYF3dxYxXORHyjBbDxPjV7XV2ySULenrqAckJO5IVsU1rtQ/72eSMRsP6gFG/ByPOlddnz2qhMG
ZPsdk+Eix3WA7k7LUvEVsYQqUFbJ4btMLB3dtYsAxmEKGxA4KRUXWaISlyMdX9DKYDUL+Gy8z5tD
ZOumpqFvz9n8kkniS8+ZfvExQoHLhzKbov+AOo6Uutyhn0DCkyuVQvLt1U/Nq98ur3+DenJvTHwH
54ZJX0sRou8vd3ArXpL6wYoRTrdQ/iN6LEaeydok8vjF8nDmQei+fZ6WLGNP18ZmucmrFl13tpcI
8eiZwqhdR5St1km/uSP6RBVL6DXrXObhIR3RQvDEFft3AY9Ahzyp3+pjTLmt8gL5ENHtdDBaalDP
xvarI34ntHWueG2LZeXrBwRqvasbpsFV3+eT+WZOTbJbaT2IhGFJGAbl9j0Cuojx8wdwd7D5cwTe
+dMP9dRm34EDEPH9pzAfiUDL0Rv4MDqGBSSCbQDsUOeRKHbHmlUKF/kLv5yYXIcQ7Rt11kmP+aba
i8GM9ZCDhKC7fuAG5Xba1Y23YfpF3zHvd2yotna1EQgh+Y9KFSHRECFrYjL28KclhmrQ2MUb9rvJ
WDDkOZjmcLOSqk7ttCafKt49LNHfaXEuc9B0AB/u3MGK0zI93MgoV1m+IT34Ysb3oMTnlvilZ8d+
7+nT6J9+ad9PsPoNJ09Uip9LER5CLJbUK4QiY6LA4ouOzy6fv0XBxRUQgXyIX49fik77jhfL6DjU
Bizg6ZWLIoEHLQgltpNW9o260mI34cMHLezBNJHPVoKRDI7ctAa+obO/NVO4rTAmUeGGln1f878p
rBQJ2gttUz9JewFAVxbaarmOVUp8FVcv1f6tM7gpjQWK/hAUq8dQkiGdOtn8tnG0O2smEF10JdEp
Il3exOBxIGd97zq0mLM51hdADPtAF1/jPraZJnX72BVVQD9DWkLH9IUBLp88YyKGpo6BRRctX9NV
pxi8Ej82Rpf7fVyMRETP69yey52sq7vRLzwT8ywW6n2YBTudHsWEk2n4TEnyS3E7ZxgvNL6ZGFWp
khYe/0n2+OS/A+nlXYy6khHDSezHGoYNkry8+l3rmK6c9LXJb80CYFlSBkvyVCwsNKKqBSWwygP+
LwEv1IDkUIpSQzLgDAmwXnqA5N0D1+bnM2zGmFEnH0HnZjQee5fOYUgFSfRdygjCCM+4uCCL6/t5
0pqQlnE6/+I53jnzecR8M/NArnhuL8K1ZZMkoo7r5qBmbOPCLTlJayr1wQz3HuJ95qXzIzKK/eFY
7oWpJv0vQsKr9lnwFvze5GA3Zinyy6+oG3lN4HcMXSK36+Ov4QmykAEyTQotKnjz2ID1C8xRLgSS
+gMxtc26/vgZwzVqZmfZTPa+BB9ZsDAavFHEZ1kd+nu/wl/BgzDfDKFajhzP6gJlWzKq4/XqnzBF
8A99z0ugYF7QPkTucQAeraK3eFte3LO2j12YD6mU20cLKM8fV/3OmxA4krn0teNiyqsc/fmGJM+L
g3qu4Sl3dzCEjec27WO7kxxfxUvMVVZReE5zLvSCYd2NczJOEeQXV35KI0pu7+ueFwz3qbo8D3kW
daLaufiAlTHerAErfkE3LuiWvR2kPEOw7ix0/fdIwM6xPCyV6FL1dgWVN91PkUtIyj1gwsdZBvnc
UGWTxgEEde/qOzgbQUqMikZCZtBktQkjqI74dr2sTtcYaJKZJKWKCfLC/XLOU2N/SQlXbWYI9/2t
S/Fwq/uKGGRWq78es7nnawvbYeweXlRX2q+gyj8RIHcTTEDOhM3kTO8UKKy9EZPgM8prSGOdXqTG
wGYLGGT7YFBIgdQygHzyhYzuVaVdUtnyRkRx6UFILr8Lz8CpwKdkiOTCGcls32ojaN95D82kGsBm
ySW5+1KNnUTMMc22LwllK8aohy4QFvqslonGHmn7sUxXr36nviAUjHB4jPMg041cPlPTYl7Vov9w
AAbWsvSC13ad88n3wVa3uEAgqEAG7JsvnlizqeOUhapLfQEUO3cxOpYTkQFVrTKS4Xw6sfGO7iYX
fImu44QnroPgGuJaWw3oKIXySooxhZ/BfJCs78axNK8VY0etCAX2Bi8iHF4IwuH++umB6w29HGuF
9nzvcUlm70wWP78LdeZ713JW5XL0o9w42aSrQAzNehmSibKZklO+SDx7/oFKOjJg6InTluWc2fPa
RWHh7s2T6uiduDZB9E8urLN4U6CmTpIqEBQc0LKAOAVOyhwCXAeBr/j1nZJZmpOsfgXGey0XJBbA
NFA1U6a3SnfWKPROnJ0sqYKU8VisH8KqwTMdXrwR7DkS+rctHTXQdSzuPikv1fTLnwSz1sUz2DqL
J3G3ZzEDqsZ+0TDD2j1VOACZys2X9I6DZ1gZt0XANhpoP3CAMhxEzCyAclru5AnZzThCTC0p3Jur
SY7dhyFRj1Ls+MbLzHWbeayXHcev+7pXhCOdCpilKIB5JvhlOu+/+1PHJJcgwlwOzn8YC1m5mBoV
B9VkPxIO3yXWukOnh+nh+WjFfUNG/rgFsnfXijK4WDnoxZRhw6d05Hz77uCN6ws1VBn0NcffuiTh
unkKjUANKVU97YBXsskpRMRxWJlt0fl8An227C5wvmzPD/8UmcxIIEDGPBP1gAv0y3BOMJU/dUMw
QUxx8FimSNAcun2K4N7ldKb06eDZzJSbHkue0E/7nJCZB3yKsORDcT3UYvfGpp3Sncwca0C/p1MK
pg7fTjgO98pXnLOC3iUnV+ghtORz+O34pYpy10ybEi/1kn4/CZ9kR30KHktALzbWtRtgVlcuaCML
GIb4s+9hfZri82ZL/78KPSfsXIeK2CyIm03VuEREX+7s16lDkwfQRGf0x95D/XBV/cMrwT2pB7rh
iVGQ5l/sZEsyDJBxrtvyge3N23UU1ef+8LsYce2St4KxdL54qmEcYx7j/xktQ9VaJYszwA/JkKB8
myIY8Q+kPbM0/eDdLQ2snW5yWzHryhYDeGwBJJ+NeC664ab1a0As65BlsugP5paSkSljhhCXzyZO
kFCOMpTqt3WPuuqCvxpmenkQj4cpU6gf095j2GK90ptKjBTYXXn8VcYhxn7zHhHS+HeS4ZbhxL0M
/jwcMaUSmN6dbY4k+gRii4TGubeSR3b1qne/F/m14YY09QJPmIzqFUFBt+846XYTcnl+e6NwA77o
E5aftRbVFseF/01tpJWByAmJo7FfJ9dBmRmxYftoRXt/wfvGrMZVodAUE4+/SXs8Jj38C7sWTTPr
QCOFc19i+l122vlQfGo1SLBe4nHkkVUO3miwzi7T4bsHsUc9zIObEIyoBjuESYFSpwPzn0uNhyAi
ZmigLDISXZ+4kiAMUIYj1aHqIJeSZxAtxdJpM3IJVVE7YGlPrilQUIf/2zjIoulWQb4jIP3NmINd
VHeRwT7svhvJCG6PaU0z44UCgX45Jy1zK7BOFqiIEUuGXXdsyEFyBybcLNP+cfI4cik/C7nxjOK9
Q5Qgb4UIVdE1ievPqWeKyL9OgfWTTnzx6W+aUcB3XM1FAffeNakmYoQvkA9yENx1/37efrI614Ix
ucsX1DnejCaCNzXro4fIHXrWS8rEyWp8PqufW8ei8a79vfEYR4Lay+EtrKdp5k1kdeR34l8IkAYf
E+AIlmVvLVTkbQMlOcY4CriC10WD+vm6JU8H22M6Pn3FG2v9nbtuB1rFWz9YlfbAZpV4V4YIg1/4
dX1I4ruPPzOTe4e7Z2xru/l4aP6DtHoKYCzqPedlBaOkspVTZpUIUS9WWaNgB8EG1cwBxCLxthWA
Ht7vBl2S9Uwk9yAg0famGAmucMXcnxZ5xpvqMGnFusbMywNx/jEwG99OrG2tNrthpT10zL061jTN
f+7vHn17G9KKRicigPYINMIPVPFWCcDuaXCh4gp+iUUX/41iEgAbK/epWdsDvSUCv68K6WYwa4RA
CL+/QXLGBJnNLk2As/iMl5ijryoZhDNSUwlejCPw4r1d9GwQPmOhAO0B3vxA3JxS4TYp2jfSLWCp
5AsSGAtz20h99us1MRsUY4vEyVf19MlDO6YcwExiCKSk9uvRsXqhlkFu4NaQGzdyl1kRcP4MK3wA
V4zm/zYCGhBX46CAOJFt+TwIjXozHibv60IITq420iB4ImI7V71E2sB7fGKtcN3XtSt0t8z1MLeZ
hI1A/pE79YI0b4tLCBIS/XvdPIPKT0DyLzhF1kO6NbCnNNvd/XzkfefRoxbTxkc80f1T8OWoYod/
7tO8PC4ElPeL27DdxQ++48A8vMZTvzbfgrMLUCPt6S5AZ1q2h4kguNkXZjXCl12eZDhYjJrzKKCh
1kvGoguHc/WVXBz4+gcLLYMJ1UWt0dbHdV6kydAs/G8f8kaAOdSK0jOeNp5tATW1qtYTZtvTNF7C
89AlaIg4YIrVYnWLw795ZxP+5EfEhOT4Crps8zbwmBmIJmMbYIxtX7zpspl0Wr4ehnQHN+Q9S7Nk
SQdTfeKy/mjGaQX1KjaQU4HvtdYP/c6ZWEOtrC6bvMCCXT1lIYe4yXz6miODw+Y8wympt4wAjBhG
Lw/IDLrgStlhGI2LBcTNKLIj/+scEs9X7j4i2qGG4oEsH1vb+tMu/2lzmiKFQq7HQiYLosptiAgm
hPSC4C8PNBmZD+9lqj1JMsjVdUh8QeGqEYYV4hHoN9+6GerdmNV/WeW2UPxT4ZkdiOOFbwRAnDT2
/MHmZYpqbvQfnhOkzd63Ludi2tdQPTGyxkCyspr3YyDFgbMDP81vabzN6XI7JJFJjleHqPQSMfEV
cQmaeo27xo8+eoTqo0qQand3F1IcOFYHw0gmWDM4iDtzUei3AdAni7tpikbEpEIvIluf/EV2hH27
6BGCSAxx8tqQVHfJuphCm5TXLKJ96srt0atNmmVqDWsB3NJwsSRnGQD1go9KZBYFQkSFpZ3Z38c7
zsXB5A0Vpeloedlc/P2rNhOw/mP5hm47GfFs8oFmcdwjVGtrIO5slpYiscfZKbw7YCAHoXtIWiEo
t6Srb2upXb0EvV4SkVTeggar34zlZDYb7lnOlGm6cscZDyzlpqFjjVScDMNFsXBAmMH3uIAkCM0h
35rtdWJmpu9+Ogjnh8EG918Z6zLwD4qD7VM8ztRWqLKQTXyrq28py0uyzJpC0OleaaGHogip7EyH
RarfO+fY9RlE80AqbJwKv1K9jkDBliKNMkbrRR34xoMtGYl77HkzEa0DZ8xmr6+wZuGh8WlcKU0P
vveWWmcsCbM5nCSB8QZJtvRvIlgLVBY9wBnDCjTY2vFAuYCJqV6Ae6haOUBvgLdkVvREQR47A0Ei
JgR0US7viYpdzMe/mDzqGOrtCCYV31wO0zePyS4BZuBZvwRUaEQLNzQuLSX9QdDlXPKBU+/qLe1O
x42YxpHaI6zsRvtxYUTaV/PqSUOdQbdfqa4a7hI0qy3Ixk1vaXv5gVHdEnrdVQvO0sgyCzcTJGFg
srNhqD4OGsHlZ16UsV2pmvLQED9iEjQ2rUXOqxEw6Hhj129Qv8UIXp06QN9YE8WJfsx+eJJbZ3mh
3IhKbPSl1VLS/6ru4SGTP5MQYHTDbHJ6NMv6plWN/G5r0wKadJ8bn060f4yD6DszIS7LlOkjSbkI
C4aXAK7638Q16wr4VnOOmhlUVLjT89O+Mwr4n12UoaqM6CthC8dTN6acBriSknLikat9yf9PvvZK
TaWI1jp33jkuVEYHvqgDiGMnJNXSavvaZG/SHGLrXjkOjMHI6Mr+mw7VlC2QxwTHPhEsYhMeAkFL
faFvyeQAKoIZR9wJMJjb/+qhIlA8jnn1NhfrLgRdx4VyRy5P8HwIcf+bpjq9Nr26034lhSi+uTuE
8vZ0HbtMhAlGqTmhbWy8nwfkS7XK6d43HoS9e7jtzxGHMyRqLTfYvYVzeFvFqYHRljWe1xnz2/1l
P5VZvmFYK8ndoDxya1ou7EcSP6HLXc90Pw1av4LAvlkiLewHSySDkvqHX04FuY4sPCniUl1o0xQ7
lGUHTkGcJl106jnI4JFiIjud5nOl2xM2YC80dmHRLTv6DQpQBYbaNmLJqjU+fCT8xW76hvE2fk1P
TnxBJXporBoTMcRPEIMMkpp8eEyFt87gyANPRqLjR8J0RduCrrbrHUaWuYVjFEwdjTvaLSIPYH7G
O6+jlvl1IgoB6rpWCR50H2+0rkIEQbHVqUxsdA85LGrwBOgppOYpIP4Gih6l5wue4UzwR/BMt48X
jIt6Z6z0ZdrXZigUSXfKfraB+QCdmnuRE3Gzri3E94HherzABUbzmAgWSx4Qf7e5+g7E4kgxU4aU
Tg/8LUgllBmG/8SNL3KzXzIWl57lzUIKLvq3Uyvobaz8RhlFGugYgsZCaVRevwAeHcW2WN1nUWEv
w5BxF65lXrcvPPDTZ76PJvqlnPFWWLwRD6d0sF5uu5+Qe73zGZZynXBAaNvdgm/ov1+trt9ietPz
sXndE2YfSMqitUieckjuxQEm4d7yvsQOMDQ9XNool3EcwEsHnIJWxjOoRfyOWbhvQVsbk95BuZ+a
2Bkb0W1GQrvvhzZB60cRBmTq4kiFTP9AOnpMLGUTouWhWMU2MmeQmiTlaKmYKqRG3tdB4mRUREbv
+SWoKo+IK62XnyTl2fL4Fpzy2U8DC78YaxVoK1uLYcPjLZpEDaapOPXejMeUJbTFRH/Qq1nBg/Km
RMF3U0vZ0/jwP0W5DozsIe4lg+rZWkXCf+oEB/4QW9uiSU3QMSfms/K0QEzHdkYYMUbDN6FKVrgi
dz6c4WMxXfKNBvzKUKtglHKuL/lg/n8Yj9ncI/AoT67svMtMvBZycHxZnwCpO9V5tqqeLUDS6EKo
jm2e+5a6liEW9Lggs1+l5yW09DdArNe/ZGNKQd6YugNB7zKH4/fiWW+cMlkJfqK5LBaF9afMGGxm
7zVstVagrp+AqVkOBgbS+qJduBcRE4g+ZajWzHsEYiiAy7ohlECbk4nt5WUj8b8pzr1Fojs9P5lv
76CTsHHuMsg0i1WuXHFuxpTOff2X9fFMHSiGuJK8k5bAnllms3AV9d5u5m2VCziH7MRQKtfJZ+jQ
8pQpnd++yw176JVKlmPq7zS7H9V8ZeBcBDTSP0CmT4NG2IrMzrTGpLCC42U3FIyng2FSvVSpAb8d
WG3dU4TlMUAA9KkZCw+KzupX6TpN0rWYnT2yUAFxhp9pj2sl7QGBHkuP2NR9FrsyQBexdzVmCW+f
s1dRR6KLutfArLHnxLt/w39JLns/LkyMWCONDfDpwI9BCCL+46kOgeYsBEMsPOU0Aa4IEe1cFepK
qC0q7DwztEAaPxSvw8LhH5gu/J1qvyDo+QRI06XhaCTo81Kh+Wis8YsYxV6sdjm9PsroBIkmENik
R3s9m1NeHgi8DPELs8RjJ+Xov2rFbV8P8T7JGdix2tFho8W8Krg1DpyDNrdniufcbkCTWud6sd7T
G7VoTNt7YNBrsMuO4L5aevmMRGzcFpDosh28H3/hC3WOdfpKW5ICkRyIhS39NfgtULJYn1MdoTmq
VAw4uE2j9VK3yjQ+kcbmsOiFn41O3N0CfCL8Eog+SPBK7rcVu5YBoDASWwFyt0O6+6QbVlHt8GXj
f2ZZF8Ro53kQXXzoX2gdllgHRvUUWnVkl1Aekr7iChBRHLcyVEd+dGWNvRslo5WlQiN7JQr5ls49
eqzx71BVNf5iQCWh0qm2vWSORmKN/PN+55g47pxmUd+nkn+upkRYd1l8HcC6xBeJm8DMUTq/j9MB
E9VYxrkafaK0nECGmJQfrOlsnTbS1eDAnouIJh689o51cZwcYDBmLKHT9bKIqptm2broY6QsWoYX
NNHfZc3WnrufFmjyCgHwtLGvD5N74Tsii6N7v8oF1JCMkOqfI+PWxvaAY652DSetN3q3apjXNCPJ
z1b63kvyuJ8SDdioSeBgW/t1Mn4GqG3keyhYZmFX3c5H4RL3pw4mxQ2O0f2SKZZRWZJzpZKZ1Gno
flYMk5J/NUzrwUBfxFht5ceoox9Es1z9b8vzVVYeCQbZC1PhD8GGsQxL6snzXcbSZC/8rHuUbo4v
NwLQNmmEhtNfxKfMgs4SA3OrdZf8F9Tm73NghUWwXYgGXq7tCWJ5ZG9kRSiW+RI5VEZyZB/v3Hk6
FO0fvYMBfr9Y6PTmFuI+dHM20UoBNj5py0zO2+XQ5bguiDhCGETriTMeCYEk0odgtm9NH9L5ZqKc
JzRd0+tMG3z0OS3SYJCFs4jCy1poF9xLUKVJ7cFUeegpnFQflicvHih2F3GaumA9eQ+WKdx0IpKU
asrn5IeyfmexJSUZ63lNUUZ2Yz4fjSkd3mDFahyIBvvq7HjCUIkyB/G92g8yvlzzKPW9aOs5gauB
H8LT3XTOYCMcfK4s0I5m7DJTR7v61l4UTherh6FwXU+tAzlwqmdrg7KqO0hWYj5jZXozUmJSUeWh
YqWtDEGN3wOYBY9P9QmWL9OPkp/+c8YS1K4MtUFOcbUn/IaB4+5IidbLbe4turqCRqzMc9uKlBYS
ems3Si18alPOh28LeqzVvbDWnIiiZCk/kh15vVHzzjayS4ORRe9P1KQrs6maeeFaGVYP42P6t2iU
/8ls/5D3bkwalwY53cDbk9tjVbf6778FHsVLFiSh8nJBzDeiMriKUosUNHYzRMsfmoLya+wa8BeZ
bqjuEJdPW1JimoU8UhtvSgC3riKCG5uOnVHFJ5kXbZN6gQj46zMQsYMgvrtApiLZKoXuvsP8WKY0
9IREWz30z0ZsFfFcF7JEvqW0iiLoW0qiifxjkMGqsQgWFlEzoYkuOCjJRJSeqjucxo3ntaBYlqJz
TLXwi6nEaHLOLmV+96Us47HkL92tfJWeyIpRac/P6XA51Ch05meRs3nKFAsBl/hZ6nwGMfTGezEh
UvEmwXuLnI0Ft++yMkyBOZDQH5HMGKykq9GCfdrotH2WPbdcOT0xi4xp3Ekspr38l+E8hK9ddaFB
G5c7kl/PBuisTA9tOpOmbyg2bIW0GK12z4o673L0tZL8UY5YXs0pKki84680k5m+XcxbhAs6PIoZ
ax09YAzVSyh7omzStadXlutaZuTFa0aQoOvBCfjkdWtcL6bxce12cVZYifbfA8V7qTXIziyQ07ae
veoOJmV9NyItNsGPZiwk6v6HzHROOFs27NzZj1I6Hsow9CcfShHWvvaDrLZHe+tJI6kSzmMd8LlA
YLGU+0BoibdAIeJkeQrADgTTumYNaZsLi6sBsBk/1uowsqSJPooooXf8OvZTJlJzekiM5sId+ZAn
XXbfFiqRJ9YrSj/RGEXZ5wv0nnnbzCBYt4MUUx5tcVPGaFu6tWstTljvySHM9G1mS4MQidA/c7VR
ihspfk6K/SaQc3l70I40jGuFuX8YU6Z/aA0YWuPl9DsWrnC+CYYuJiuojNLThEK5z8PjbDS5yKP0
MiBvICzTN4tqWNq3ArfYPUr+hjoV4qn5tU7TqslsXqGS0TZZEeKiW0iOXbqjelofAOAHWY5jWnq1
bsINm/yEzLltwH3LAic+tErYHI27FADU8XymWTyf/CfUlJwLfcFKxV4+8d4oPp1gJly/bpFimSfu
xxNqKKpLHGuYz/9Hdt9HM/ijIRu3zgAaaqeGpbyv/LwY3uxCG4A1mZiLcDbSNUMi8on48+QysUFJ
CyYdmhDHQrSnZvalaOnf4mIz6sbngF5rMJx/OiLJRSKwUgIsgVwHYboxj8HJspcTM/VFpsBvN7os
ZJuNbJ8j+dbaFtYKirYWg027pRwZUIILS8DWzCfUx9OU5Z4pi1SnTvwavSPtj5LG/lO1j8Ky6GR8
6w4w+K1RMq/64q8AYQk1cKfdE597L1f1P8t+Bxrk7n8D93N2WegUt7hNq4fy6qGD196B6CM9Arhw
aRXkSTZ9ftaHW3S4UPMlplC0wI3CAa72ZK1OZ9+2uMxHrVIag9rLQqctHscHrjkiIjmSq9C68W8a
ZMM8guK92fPL9leYLNl07hVFnGTVQuerJHKRFf4cSkvbuWTsTkQSyn108E6HY+2RMODWifTlW6gr
miMFDg8YN/sznvbJBvl50NXaWfmlolECNvUD6FsRTsx+mr0UAabf7vK3OkEepPmNVqEJBytG+dSG
DgODrTITveBfpbqJTx5r6ZQhk1UgiRS3Oxfr/waW1cQ7HprSxgzkxX3mLaRxIzKeP8pGqihno0Uy
spkKRD+pSRVhVvEKhRknqhe7G20bpMbfhqJyvSUYZp9TxZvlj7l0dXCsVtPBGcs3RRjKZcARceQS
4fl6RywNEZ3r46RC4KqJCKMC0F0Wc2fOG9C1BMZ77sgUCuS5/yRTp0+tEEJWHR5yTjn2tQ6rPrEw
pMoeAE7QWwqe2inp7dUK2CN/vKMEeKsD0wYZhOb3Wo9ATu8jxPw6iY5UQTv9arhfyNUX4DuOGYRC
tNyfPLU8I//eZSympkZto1NZkFCpcShgVKrUi85tVUtfSBZxti3c5OWpzgwlMElyW95KlnC3/TBo
ckXd6/+1jOsOy3NP026Wvwdf1LHwwwsQDDhYE7eF8Xzwc8cjahc/je3DKKJUfY1VcgexQv7harHk
ncscgve+2zmgHzQxu7J8P225nWDUXisgNpZZ1W20CKnhA3mNlUHo8ZiIsfebk26MPnT3r1NDjCZg
gLElEb5BQiF7X+s6W8K2PoaBgd0toSUTzCl425LVSbHDP8FWbqf7m9F7b5i5WL4d9taxFGIZ32e8
DX2S+5fTnwWE8oYyv41eMfDtihYohKRpQlITQjJL3XS1PnfzE1EIN7OMNWLllXJMzDFVszaeUdbb
IpK14HIVYMBuZJmQ0uddY8cIQC1uYfuoVBgEfrLCd3GGmsd12YXeDNnT/NAfItC4wuzH43P0FAkq
oYPjysrCQCKf/N5LVNmfAFNX/sjx/uVhseTKGKZhJJQ+Toif51ERE1ayMVS08WRq7a/PfUtNjSuJ
RdFHqx/7fTpprNYLfo5uVMhuohVEeU80OQlGWD8pTk64Pt9JkgLDON1mzDtw+fFE/Wcx6yD7pYWz
qljXmdVlGi/OlRJE9eJ5DLquPxMs0SaQXCOkqztOAug7eA98U1YDS3MOeqDuVkZt284lC32woi9K
Vf7VUmiFvjKxo8Js9ByuJ0OoNNYlB/Wio1Atg0WNMzYgFbLA4ne/WNBYsmokUdg7WfzHsCqVe05s
Dnyx4lJPP41sUeEMie2uYQ0ZWELqyrmrGzlijEapEYzQlKEOFRhJceHzXmh2ZzHO63/mMLOT/Tk0
uTxCkxiZHRotO3IqMPMPNImDWpAs9IcHklTPczrkdbugDiYD+3pJqFt+3g/qSNMy5QLgV1+85mCK
9RNZPKRsir4ATZGJnhzDlCXJ+jAP3HUD/Rxq5pDvs0dtSwFUUmLmA0eyJxPnSp5cn+8mu3HO+AyV
sCB8DT63k5fvECGK5BI+L+SK0GjvEXzwosV84t49+DxvRmu8GPRH/tsiSaVobIp1regHpkUUUdqs
SbdnIm4gFL0eCaxrZ3OM5rw3397Ntu5BNj6N/G39PF7nW3I+BFOqu23MvTh8/TzQ/3rJ7rT1vBGh
lZVGZI7GZnk5v/pM5BUC9UrVAanBlLIMUU2td3iY8Cu5Eg0UukJDrkfnuUwRc6xf6jeaB4k2/Tds
aO9yHlLhhyzPA1ucQ1VB3mHeWI+oYEyGhyWHAofMIiymBWjC1gEqywfhyk/smkf3KCJb+nE5T5tk
U4OFzLWehkJmTPswVelfxviXBlKRdYMqm+pmiY4BVanH+WunBI/pAexI6rRiyd4lYI1JGjANP9Pr
WT6inF6wsjQWoFuOovOcOEKAMKnUbpDwd/AnvUU5lqoXcsPpIxun/5L5/6Vf1XWv5CRSvT28weBt
kwWB9GGv/KBzR1NGt0Fa/IWaKbWPgJIScrPNdmd4lMRw3IaDq8t5kLN292oXmvFXq7tJdi0+y7a1
5KuqY+YkZU1Gy82lzLmYCvYPmjsylZVci3maatZ0MzGNyKyw2vrGw6jtOGSn4SPbD3/Rc8J+xsul
mIMhRkAKH1vKRAjtUZgepbsgVDw9xs2daLlU3QZyq/HixAUmI6wxvAP1cXoDx3dp37YclhJ3eecr
xUJTD9b1a6HMXlqHhC0E95KroFmqbf7ucPWNkBoGSBgFNkwMMppzlfSmnUokMKp/gP7V7Gwmg3iq
SeNHvuwas9wAK1StaPowdfCHZKkEV+Pfwld7FdMajdbfjjeP/ahcPozDjiINMz4xPX354vE0XtEO
XwJPTTs1PqcWfk89d2+UDcXYLWE9dZoJyDla/zEBn7VcfXgD8WWCYohfNGkCQD26KLCeUjNen8Ca
X4mT9Ai3bnXNmLHu56FLu3VwKII4LRCGp4ll8YJ4eyU1NUm2oXecTbAz9Y3rGxjadcn53z+91iV+
7i1yaySYnli9Hn2m11CONdb8XyMw813+BzJFA2Bl7cWbbU+hEtKuz2vg17zWQZTA8Mjorcp8yohc
H2UIlPnxCOm1Vn4VPG7OfkYvh3uS4yXDbpi5fDTFfoa+T+nTjPJ93LAmFxRmQCAt2pT+5v/F45Np
Z1uQCmKX//Tx0kn74MW6JqZbBEhNI5DFau3zQPu/EbjJOEb2FNBYe4N8dl1qLRO7IlqL30vZ3vHS
nctWLJu56KFU5F6y/6cOlxub9NdQKZdA19QpptxIXUaz3rIbSs5q61V31aYsS0/TdJ+2BeXjSnAg
fxbPy8rKdXB5h49FepROO0FfKHcRPEA1CvMxDW/acRDT0RLsZ0ejFOcGcs4fbMOUVwlhUBhZhSZ7
MSldUD75MyEAYlrmuenj/cOXs5WREdWj9mNhvJ5NNQ2YQiYA/U3fydq2IfjW2VDXvvY7FPQ1aLih
f1iyEpDtafw1V2JUuNP366pvPpz1l+P2y+ehEeoNDe5cGSNg7pKPRVszoqUw12ILDd4wVxjt1nqd
JSDs4Sr0farRRVEO/1w3UHxdI/LI7P8uR4KEht+aY4z1hZ/dz744agZCsby3GpIx43Fc15bxKXcc
rgo5CILEmGK+SE/CMPJE52+11n273jQ1YPouo2TsgxTYSKETe3pgNUgU1oLwjNmYjtB3Kkk+G3rb
lYID5T42IjbQccfMpif+KO1L5nnTYtwLhFQttNBtnEVbtTfMwpEY9m3uFKEl2RcO1KvCELv8k2sw
e6TA9nqxTthMPGjkLJoFpw1kzLaDTZkmqlfmS7Sne05uI9lvHY5HbKWYdkRirr5Ijen1UiIMM47f
yDshNFIY6Who557EY9i/DcrZJZ1dX7GbSL+MDaysCgwbYzZEF8ir+S/GeV/2TfACWFw8mLTT3N/D
IFP+mvNcjgaMdpEmMYxWM36fOp/mIjbJfIwRVSgN/bkWhTT03oDmuMfnzjpWDM21d8pDB1hu+4GE
PXfPQaWVjoYRiR5b2jyOk4vIvDTIbVU5F/OciV45pc1IXmrKuZ5gaWxJ+7LDJFDXjsA54f7k0GO+
ViDodaTnwfATHl2tgrqnTrqAXZzv8cx2LTAcZQgqzVzrZEBrv72XqP4zmP1UZ77aJN2bP88V76P0
BswHg3WgH9vCfc0p3ne8QWWfd988zb9n/7TxMNIcdjSVRDSaT/AKv5Fn18sahK2hPq4/4Et6QMpE
KCs9nrwOHl7BEZGexvnTn9X8+89B/kxLTYe4XASKVz3RXhQA+TTolaFYx2cjOAnXpBM2fv9OjEzo
AjnJlf6JYeYPx4BAdOBGFrGlBzV5AyEs+gCiQKKZ7Ie8AYIFt/btR9+KwDeqYcsOF4TyaziMcPbr
X7x7sITZNDhnmXxR+2F7f6aQDP/zNv1rFE3WObUs8dNLdASEVzGbpo60ct2A9TvY5ritWLINw4qN
BOGOjp8Dyjy8amSPNOo95qzR6D6Q78t/D5UoVH66m6L9e7CN0T5fAS7duo9KEIMlHHrh9WQfDQvM
1TUmIbdnCCl6pfVkBBj7cKifjFIXOkWTyTFlXkCaPC12owe1KHIsefFxHU/ql/bPCE60yipWdAhZ
pd8Dr4rwhoGBtAW2m6ibgfBEvQ/nP42Y+N+KYqRJwt32ifqoM4DovjwWL1gFGIbk2TF1FXGCsfZy
z3/207AAujsnx56HGX2ePnvFBX8H6mt8cq9GmP1MESOnuPWAIhXZHvsW4Ocx9RosD3iP/19/4EDa
fl4J400BEVO9dWICCTo2YWe4fA74bPwkaY8cX3dMElAfvVrgonsgdZLaJjELu3Yr1ETHNeeAq1eE
W1daYAPO1fwF1aHhXeWuxDmIcfVW8wB7u1b1fm4xKgaXBUmVbc/SFDncscLAH9Gylv/NZX9uCc2A
nr0Mcwa7lBwyRRttPVS6RQ8iYNYwhtI4d69TVNfYo9m/YeIpoEYhHbt1nI0sx18fiUrt8/z43wYp
YcPDP15M1pbwd32DlvWnTttOson7f2mWAJDfuzUf60kah2nUiLaTVZzirFRz1pPV5P2q+fy4MDCx
0EasB3YBM6T8zUQNeDNdVeoI7XZr5yTZwL56ggwSBkOy1hsk6VrpMlu8oi4lYmtrBIrc1a1covbI
WGTzy+GfSSSLNAHjgHn1/6ll2FRFFSFET0XUKbyYFZT1+iC1zwfweWeliwcfJwvguoRDBa3tiVGh
y/3WuwZmATbcFdcLRqqX3dg/4kj1WYX8f0I3ybLPO0toGquN5AJIXDrEnea/LQ2+Sh/BuBWYAmXH
i9yO3t8ynPlt4Ont9D4/StlQwge8eTsNPaobhn9qxm1Cv/P71MiRkhnEUjTAGmlVuXJxsXyaPC9K
n0xblW48kRMjV4jM+s9Qlsjzc+GaNye/eHR+Soam76SwwSkAQNu0WBlNus4hs9ZF5+GL9cVnO9wX
7hPCuRiVzu3bJL/ni9L5koHsDI9Vg4P3INCXRrJ5AaAWoycb+QvtY6rXt9Hg5/N4X90mmru22ZWp
TKRFnfWNISGbsR216mMKe701WKPGAYRj6w+E3jkxoXUuAz51dqoVwUy9cSP4tQ8PS7UJ9RrQH3IM
B3qKDzylLwsxeExbeDMA8x8K0VozBuJ2eAeCXNFgSvIo5UYU0TDX/fuooLvDCLiPdmVx3elVph2j
UMw4gOTwWg4ijLix0TQjOxC1Ufqj0jEHHNAjhsCKor8QvtiGeiCPf1Vsbyqjm8JYpPJ7i6KYFlD3
kIRSuVXZOQ3x9q00PsaIv5w9rVIpISYjY6I6XSo6fNaWyfNa7s+yiA05cfwO3+d7CXvzo5kuakKo
HPT+o6fpal9lXVkbsozfBZUxMt1Or30zCffhbq2wk547bep4mq+k9fKEulWHdMlbHi5wNJm7Q2XU
BW5dLne8U7p7nLGnwCKsb/xhePmSYhQNnvFOQz8bO4rqWr+Y+tPdlfcmXTGkzC7KEUtXRgJcD7jq
nF5fzzAGfMbP6bp1r7pi8JTSQsVZgIZXpd75OZ7/EfSYJ6JRNi84gKY5qU6l/K2DN0I1YETgmcCx
UAF2Ifny5f5iZ8eza2w/oeWSCjqLk5Dz3YfgIGP9eg1My+FhyeJx2RhxNJruXoP+jBRLUh/bcSTP
/KSM1ovly04mXLBUNAJ03yTiJh8GpDh9dD/W4xvs6Ix7ufvWwIEPtO7Ip3bQo/Ofly7vMpcXYk8l
PMrGJFxBjL7iPeQOJFR85nadqFN1lStWSectOR6oq1MyoUFoGvwTMLJfwrDBfhb2uZW1HDpppTHq
LGGjmQ5EjrIy/WH1uec/tMyKItb09fGX8e5Objw2FOVdSYT6TNSjZTnwXUZEaxoVnW37Pox5tof9
nvQVmJmahndpnwL/OdHeNFYIbbF1D7pjs8w0oUcmUrFf2VSGZ5Y8BwBXWo5QRIx65ACP8iLRSkPs
PvSyw5BOcxa+IHPj1Ki0wg4yaGa10tPj95Jq1NTqojCNHrPjgDo0EWtYXj65Eoe3ZerAVOUZaMmw
/QMymkd7g2iIf4fM+tiXPNwGJzh01SZ15uOIk16bUD6CoIZQUntop5kLr8Iev0HjnusW3MrAsVmk
2yP118Z0WsTMKMGbCuvoAJpaMOrj9HPxORQc78tSlmOZ6jkjCK96Y1HQoFQsYD34PhZTI+NCfSqt
2oDmVKLa7IKYkcHPkii7fS/w/+lSGLG/eYdBWaRNSo0GxJOuvjkhD4XB1Z8NEpkbrMDthQqw41SW
tASrjSed0orfW2KyWjucv7tGPAdngJLI6bZNVVFX8ptrVhSTuPz/7+x1zlM1vXiyp8DrbFAUvlrS
EIMfjpDk+xL6cEWro9Fq7nKEQsg5pCdG4wa0TZD8MZdnSPIXSUDPoRHqTWSZeXbrpPJCrqrvlGrc
ZUKBf3yuJ3/dLkXrbn1C94pkyx8jXIaWyNXOGfN26+/v0QqFKEZfixAiLFc4aFFXzQfNCKFcu08I
0LzcztmnFFDgWcJBbzHu7oMScdH2OclGboM3x7pdHWV65SDCsgLOi7SkCvNabYDJ0uCheEz3bWjD
R0kh+YCbsomi2kBDDmeU2IadEsgh/ONxo3C+hEhe74/T2ma8w1m+L7mqOTPzG69S/j5yCN2ZvZ4V
+9CeJRPU/ZxnUrIJJ0RzNCDiPuVrhY38vGkiDm3IEgJbVvX64bE8fOrtVyiqidTMHoM2775zY9G/
Z77y/sHziol/OXbOCUwPxLnpylKn4eMHqn08KVWZIK+QX+EAltrYrUCVIKM2tIyDK595yieTwGTb
8GZ2hzjS+o7fBt+X050zc7FnvsHCeLDh5RRILo6JW7DqKdfL5wz2Oj6ESy6ZCV+cUmd1vu3HS3H3
rdsmKQn22c8h+m+dxqdaTsVYilJa2GoCfuPgAbQyZETlTu2AQekxvqIV24LFpXmQUQl4U/kYuzxj
JQ+RYpAHm4rU3t5MLTNEfhfdjNbmCvncxf3ntBIYacYjdXl42EY975/D4cCbgUNBNWnI/0K9RvlM
EJ17fdGe71wg0/EdUTL5+O/8bj/1M/qxTLJ/lEVPXl0oCOjs6/MAZg0ue/DUWtSDO8y7WTsv9/RA
Oqlbd8UprJlV7Bmp0/vD9G9q7XnDLYXdshq0bQl8yacYxPS7PJcXhPIABFmu3wm5Ev6fUJ2rk3ti
VVPZUXuB+E57jrxZ2LYA1CUAkrsC2adw+ITgXj10Fjt0eS4AqPm0FTx/Y73uFx7YUkEzuPSTfScg
VfK2pz2yqEWtnlaQlEI9Py58IZyeuk6AejXvGtNfJ4kYzpWqqkJIrBiXm8Tv/L2gMtLJ7uItyDmJ
0UlV9aUyTY1Bg3+f3MUw/Ik6b6cRvcyJYh5cmkzZN3ZSt5Ut/Kp6jP25q2fIHVyGnBfRl5pjCdSQ
H2Eb1mR90VvAv+4OGna5xGbfIO+c5eZm4LToNd2K381MlaYtHhGXDZ4kJmy+zGl+07M+tf7wefVx
Ek862XVsgq2pSva7f6ecac8kJzYARwG9tVEJwp0nmwUMsu98PqUMEBOcPNHb6jhA6+28WHaWlc12
H+oZF2/VA40SmocOoyOBbCsLkkFalx8jfRXZAOIPrx34vJxUTWDvzGDHapKuTBvF1UvjypcySVoG
w7WkD30RBWfU/qQaO7bj3JlwCeuEJ/HPDYv7VguvBOk3DdzWzaObjLe4Cc+7e+WBLWv80wkYHfNY
hYjjFSdTIlD0Yq/910K1MYl7af1YDBlNy2+24R929mY6gInOCMKGWQGdDD5vBpoMvrASFR+s7vF5
MNpr1c2CzIMgd9t03qebfNQwmvlJmJ3Jy3Mm4gsf4qMiiPEzb9FTiYr/jvz5mNzsAL1Xr/c7aBhD
Y/LHwqJsjuJECpX1DjTflZZRlKDeOUy0+3lQuInwEqcQY7FgSLyzEp69YpzCcl07z3WCT2PBple9
d0/rCtn3s4KOJeIFV5qcWNzK1DVJWTwo2g8s2sEDwZu+X0DR7G5j3sKQOXqpPBx8IEhp+qOW0c7n
StaaFe4maSJBil5n/gYe9aGTl1DCwMfclybOWRKBipdDAoXxI1eHxbzji+2LFWsnDhLV/DU9LZOb
6fjrWxUCwOqUF7eSDJ4sKtY5FjUU9LUv5MO02ruguXBVWjiTbMzsyh4igXbVf+1cM+ZTrxwNN8Wm
Sjw4WBq0MXQ4Qweh6q7/kSCjpv+0Q5P4l6QAEybwnb3WDV2RRJ1lg3sHZk1VOgsRUzSABu05FMgr
18R/xJgHpKg+mPoJffffwoDcnKxy38lhRyNIpaS6x8yqKobxJmr2uyv389qovJMVWOjdGjOwgqLg
PKlTwtyqcZj+Bp/jMYwmmzKYsmpo3/ELthkWZTCuOsYAS0DH3cqOD6ea0OpkPRttkfXx9C7Byi1R
KNqJqmznLda01CW1C1QaVO9HPEHAdlO2kII1zG85NHFRDDhF/+9wF1yen0/G1UaYRYyahnS2k9pm
Z4+DKlJpaiwPUr438FjNZh5lNXl4SirDuK1d90G5UvFto5mSE10/zUwc63byD7Y8zEXehXg25qxW
dTgKoU4ogLK35JNy0pghw7/XXf347DU9kY2DVKpl9yuf88r/PEPYZiEpPXme8PeK14voAQFe2OoT
5t49lbagl9+1SUZqp2/Enb+C1STUxbT2jmd3RhqFtBkmj5CiOnORmgW21PRkxDEfbdWUojnDXqpF
NRckPae86UjIp+wVwesqt2tO9vbkPCYglaDSqQ9gL+7AgbCKAdEO9ugzeYn8ZY+RtOLE/FQiRov+
HDBhg/WNASy/tBTNGlUGgCd55avFtBBbRrPQZz+k/D3Yet5eBaMAL+kD77keFtvl+qphB65Gwz/t
EZAIAaWziZcQ4Jn25t7DGtxeZtOQJdKGHAcdydlarsLZZJ7iVpOhehr97u3KTx36caEYbfYZEdTQ
a7lWzrO53CxqYATlFA5bellZKjwiw7/Z7TLLc1ANzjJ7Q5qssxevZwRT5nV1L5ezzOHmMrCaw8Mz
ATgecnyD13a38AVVuAE3uxwhs7OygmV93pDbwPRoZ+upDDyakIjRrJ9nGqZJ/VIjiw8enopzDy9v
3RM/ipamJkPxZuGeMXRgBjtYdoGlIFH0vTMQdUp8E3eIy4HAW2uv5MzfErju+BHhkkD/gATry/jv
wOd5jcU79D4JXiTSiYeCCxaCVxs8GWFL5Ecx0oiOwXkRmLc+pBRdMoJTpzayAa7Thev8s5DRhruE
A0gJYGRLjGT8RG0Ae0tc9zZ/Z36q6UW5DQT7ZrLPwno2rp+zR0/jIYIwtp9KQBbgH5zEQqG9qg0w
bKI2LEi64Mikfl4EifLQVm+Dgg4ybtfFOOlAlZV7uYVdvVFNaiN8lXqFdTDtZmA7d+3jNzk809YZ
4rmbxzrN1P6YXc5bjPg/PW5rcBIiHCVarW8cMvP0g075Co4Py3VqiOJPOZ8PQ+HeuDI/l6bd1Wim
5eCBV3P69QIQDmVt+H5t9rTUkea2Ezg48ZeYJBcy63yA7W8bnvsqBvPmxA+8mI5Ce0A1KpTJnzdB
XCMByoDwx/I6UhAjtt/M7Rn9upPPDogt1nnf65HmCNgm6fLIRUW2l2WN5+Udhk/h4PVsvxwlGJ89
NfSj2oppjQCNfW+x15jOFGAYJ9v0CrXJCp8S+ZV/5pSNPVamRDz/FIa13rrGX+OAa78JVQ72mrt0
g9iORWFxbHs0sbge3utl43lHuxBA43S1zdQuXkbc0c7rSscxlp7+eNPDntXW4+PZ+k6jt0qglwYx
r7OwY6Myv5FhEqLh0Lts9Ss9w5hGVHhEkTjzXRiC4nS9h3affSkCmdPEGfvNctQy1ti7kS1LWuCB
7WhiJECEDJ9zkwk/Px/bspYuUbuusBpBzQEijsjUxjFiz3xsntMVvJmyBz0rqt9v+D0Wp0J3KfAd
oRT97q3hG2GxgYdHYaJGh/mqRMN+28JlxZZYrMABTRzr2ggPy2rFiB9nq4/PQR/ctDAHmAHuNLlf
5E82M9hXvS2ZJe1sPEnB1FpcZCmuMOQ+bYAGQQBDHwKsozu63IBp+XY2QM3oNbg1sCBf+mdRyFuz
zyulXgaO2nwtNzYbY6zUNidUgFGhMxGscs09BgCj1z4IlU6SMMCg2O1GbhkQau891uMEhtCbonF7
xbtC06fmB3CWaifYbCblvSS3OR57WFEaCQXnJ6X7EXrGi5CGX5hmH7dfwxar7uAH7B4644bE89CH
ElgV2479fC/RcHLjXzVYJ6ELd9ywFJnQL/xjOuIIG9qR4M4A9YMIBdo+rC08OZ+40bIewdrPBs2S
MvuuE2Uu/rzMxRyiJ5JxH0TA0EyuQbkgAnG7uHHHGxZy9tZRFbeSexUdYpa6I7wHtfTY0noiPu5f
baYsJ1FBVmA8de8scInAmFF13QkRO/IOBoKFdh2JmjIW1K3tn6mFGmtWhaIiA1dD84dB6QdDh2Qc
F/JWg+h1xv6FrllsAcrUZdRyuFZcKic0SHQ2gBgCPRhcrQOQlXjTa5ZDgG609QOm1Z7T7RvwwzPY
34ub+gi6BW6Eb6ql8xcR8wB2W3KMMd+J8Lql7nKotlQ4S6+AnZxl/ZT1/RTQGnIBWyXEvpfjXCmX
7UtYiJ8klS/2tXo6i2DLcFlp04SZLP3BmSDWd7UqIPYsXCI+Fctq52MeBsmhSwT8iYTwK7ttqHNR
YF9L04syvCaLfD3PNVLyLGVfz3NuQ9dv+e6w/5owzUVqix4CROlSnApXVtQPzyeYD48rCegvjXPs
s5KWaekLK76gDFtlii3G2T40U0VxXvqMLI6Bmvty8ToFFguW1nQQ2AMQin6jIrfFU9Oq5Uar7ZTl
XYHr3N5H+dcPAudrqIy+cQN8rBP9aD+jPfiq5Lp3Svp8w4HLEN8LcSHs6zoogZD4eHLuWHLKYzfE
hwUD0z1lzKfZu2x3FWWhcbeG1+hZVqaYEm0eoqnYBadxqjI2cY9SGfbyDqt/372MZ2Y33/GKpXee
zn2NPylqppKfan3+b+LqoDZyZQlVaNm8cDNDymeuv8rFW+oJaC+syF2AhNTxGlbk/TtBuLGN8P4f
zIIHUKZmLqtZFU92gfhpNiwA61bXCm/t4t3hHEtECkaD+pUJCw3WAeBdXVcu/I/b0tmy3l3QURBt
bTg5TkAIhtwwtwovXOLEsXZOv3FrCCjM/8uSSxQ2+zmucDJbZhudP6yfFlA61rRHkb7DtU8KRMFY
Sa8157/sKDmQgcGDqQTy14xq5DFZBi8DCK3Un7N60xMfqQPLCflDGa83EdLAe+vAMUw4J6CzR+ki
QFBhvzn1qS1MSZrWkV9xkTCfwOqq/g6i5zHTth8iO3qUtjaT4QEsFwJk2EAjHT339OBvVByMDhtn
N5GXjCb7s32KjtebMQSHcVTQctpluMIJR9j73HydUtiEDqqsk/7PmqteKiMEXKt5M86HDUGTJRbP
On/nBolCz4qw+Uw9/fZs1DRYtgh5UChboiWtRglOmYLMaWgxw/I6Cw56dx97H2q/zYLKvw1dPsAJ
XGNr1uipso1zhg8C1EBDrklKiWhuBirD1WtZ6z3fULR11iyfwzVNQueEH4EpL40OwrMvDeCceQfD
M3BC9ydRJq4f+GgVkypQf/JZQFZ9nPg6QUaL0T0SapxWYt2FepSXxq+zO4BxYLyd3mfpm2IW4p02
6Do0T/+6DMqay35PLpmzfad2IsKpbrrGrRJcBVUeGW6O8C3vXpYQIYideDBshz+eYE2fRopM2IM/
NHSPPcsCm+41Qlms8qWp8RmQ4K+BVw2WBCLoV2ucf/+IElpjoZ3fF8Nk+59afEUbckDRu8abMmx5
SsKN7PbwR5vm+M2SVDB/tMl0DICznPTYZ1sjWel46Pp/ajauXYIOq5tLR+GqjELmGGs90w/mUGPC
0moI72Q6hiOejxRoHxCtY/Q4Iaw0SbL5FHSIIOXmkqYcoVwEGy4vBBUN50nTr5s4iMhC3jWPcgfK
Yk4dfQE+yw43NoCCOKklOBHae589bK3BUvGeqgQRFmfp5ttgLAOxPjqBb4VGbMeokbPwUg9oDp4R
DvslM2/G0ZqJiZYwMRBYZ/U+YrqeCzRcjgFGy9WsUG0UoonRckGcPvRNmmtZCWautdJuzzEiv+89
yJZOBA/h1OIHYkS+0/bh3gRVUbLdJehSaNRv+dNzc/zE/BsF6xTmE7k/tsmNfA8qispyx6VEDrzJ
Wj/jD9ydAK0cpEB3Km+QM1iWlY7UzxGHuDzh68njdtgg0pyoQTBd+yFUiBRlb3abEeetPqZvAzkR
qd+/zDAsfVuVI6yWJtnEpoYm5CdqjQi7yiN0j+7P06UwpC+hq4U/DiQgbG8aMraX/bK8AvMfcZOE
jnydaNuL1AofMyYdnzSz7ygPisVrXWaeOnu5xoSOIbAMggms9JRI6rr/IDjwMCm0s8eAUOIcujdW
P0P+ilUMChUdVtIzZ+vGBSyh0C2Fvy0jyqviA463S2KWjmABlc4lXNZOlcZwohCHoFb9RoUPpOgl
Id+tJ5QvJtPnkQyIXSZXGqYHxN+GIGMuLEbKtaiBcoklYz6XsQG7ET4GqC44tvx9WpGucu3t8iId
ovArH7Jbr1ZMVyvCBxItqLhAFJ2A8qkR8uuyd+rLvBC/6aJezz7uA7yaehL2GUUK4ClgRI3VZiWk
BNJFN7/5BHXulk4oIfDvHCkazPP+Ud/L+z/xfIkIcvT4/xDMzXtd1IekmYCktW2ShAIA03IzgwIV
0TQnLLeD9zzEN3wkLUrHVUqMIPYNJcO7LJwbxElqV4lM/Avq5HnSkZ9DdM9LFyyTujfmtYLWIrPm
imyL8vpF7gd2PgC8sCbx9xCLbB2HPOpOJ7JgxFtLdMOPWZicdAJ/RYnnKNWAb8VWKTKV8si9NNQQ
yFRRkhKuS5KebjjqzWa1v4e96AhWgEFrQel6b9xeoRxMe6f1h0pgv96tceBqYXDPE/bcB1Y5e+s+
oA4HbTRS9zMY/MB0H3LgYnLnd4lg8/zzWUliLSfQg4BxUpDzQzMAF4yZEpPJx9WyMHKhB047f0S0
VH2LtIESZPBDioBYQm7SKwYryc7lj5kCJOzLWqOMxMwurWwdiyPfsGrdI3K1F1Uw2vp8GcGQtmYM
9nwKgAGRgHw9XqtxywRxlD3C8YBOOD0ho78+VIiL+Gz07rRfOSWRLwb3WpvJxl05J98x9i7UnQVK
ngNTB/+s/0216axxB+oUFOwc84oxqhn6Ncbbb6zPIrlkA+wWFRC78C6fNh6QGWuqdFZ9YRGcK2Aw
gbxwEJyqpvjy9q/wq0onDU5g0kBLtev0cth1I5tG/1i0J9HSKhUoz6Yh2CO7RuSXR0JBuBohnqnZ
e6rENZE4mL6tH9FgT+5Frsg+RVW+CPl9h0SeVvRcyemvZubhCK9zBDaqTV4+upVgt70LQ635pAOz
hAD8Nyj9BpvjrrC+A/4T38x0BsEwHBO5y/uMvpyo93Vd6jw7/x/9rRsO8VW0l0BtNdtERa1/2Yf1
g8YZaGa9GD7RpYVvQzLQ3JxgaFBWvmeBq71ygznExRCDRdj9sCCooKu221cYNG59oDBD8GeVirBc
SJs/4nWApORcnPGzZia92ETyZRyayksutSqmGl4mSdX5HDzFvpouh4gTUjW+hvFRBwasgmOw7xIf
ET+3Eb/c2PCaVhS+wmVveuDumC3vkzHKwbmzPQNvVJQOterbu5wjCuiOJxb+O50aaHE5DkIIj06i
iXY+86qjc1Dis816+CTDvoG5G9CaYCgjyRzCVdQtlNvnr5mww4Dcf3i4zZ2HcKLrW0wlNe4VR5fo
rUnpFBGtePskS8kQORbdOmSlYc6SieHagyfoI8o8gVsaEXq7LxslG/kEwsW2PaRdmzObMG/1k6r/
NZST4K9YfdBq4lw8HU6PEF7QdsWw1id0xFKy5+vk/zr4S867GXsSsB1lW4rIhWShOAAOz5mUp6Dx
fW5x+8YIkxu+2u6EpooU6cACrlsA75hSkNrpYmNfplo7upNAfpNQ2WYECpnM6lPRbgr3bS0l4iWi
Ndafo4AdZfw9yhlwCsWJzEmEKOeWoYrCryjrtG4JiTZIvgr0rs/bVGGY5v/07ueHwgYk5lFxP1Uz
r/U88zGywvQ2TpxOvoQ5XTCZNCbxAzRL5i0P/74frFz7vQDWuowZdmH+Eob/sQQZmPvWhqNZFL+D
joPtWWUJBeYUBg434Y1uYOLIprb4GjfcFYwhGnLsPx95ykpEaPO7IcwYTg0Pm+nJcCtX0vs/YSxa
A7iRxxwRrtOyKW5YxyYrTU1V5oCAU76eX3Nn2xh6iC5IpGw5dwl1Kkhu4tnmDMZvSgEVFtbX0JPR
HjB4zkeR0pDUW+bUiqAK+5Na3Dl3x/qKO74AYkrDYv0lf7OOvJYeahhuNMidG9L3bhV+kE8GG7hc
Z9nlyyy3W4vvPqaj8BmJxFE5plDV3c7L6bMVazB+pWGRBV7GI4KK8nZzPgEilWCAn5Vf78iNyCk7
vBcAurA8IMAVAieMaNkJOIYXAEEVj1NDC/mqqe/zzPD9prcH+67U13zd3AOWiwMmTaLAdq2gR5ii
mscPOwGQd+FrnjEsmEMmGzqILhCaK78p4RGkxVbfLULtAJj6lTVhhR+nAArcFFTBAsl4LBsm9ALs
MSChPxmwYYvIyg5P4WRyJPizSAzk2bposGwzPISwDqiS4OtdYWx0Fo7b2h1jSpbME5J7RiMxXtRm
e/KG6wWQ19Bay0e3B4Yd6X1mHRU3Um8AcOkKQfDjUCeOa678zmZ86i/GLjcgTU51NLOlkWqJOZ2A
gZXS2yy4M3oAdrPLLdN7yb+2fVdWSxXz0+An6hdKmRXaUa7XSkKhUbK51QgelCmbKHcPEHXMgaVx
+bn9lQu0ddNw/lm1giEcT+OEkXR/8dDl+629+xFSao6MT+Dc7jcrfrm7SlNy98OoMDeC3ltMn9jX
Ge+oLNvvZ2ay64hy9kNSq7D+6borRRcRr0f2WZ99IG/jDRGChzSOPpRUPhnWTkG4ZB19BAPdJxiE
AfBhG/6ORh6vdeDgfJDbXz/LXHcU9fvgAaNkRT4o3jH+OSMYdZdNOHb4cTfAlYdwQp66RKI8IhHW
DvU5KkomJZGnyya0mJ0K4dfr/JWpTB7ZgINaW/+lmMAD1M0Aw0VVXl8Bei6xdPkX0AVIihwN2gik
ZGkjESoJeIdnTo+mm61SBnSZ+94QxtDUaR4Nzx8I0BKurqSKrRqVwOFRhme4fbjVVVPTDb+m6s/m
6yZAJujstzdj0QW5VtfI3b5lwH/hv0MgdC+uI4a41T978wQJL2JtIYA4qGyY5mitmy5hMKcHhA1D
zonZq1oTHhIi2spqxK9JYQzNiZ/pjo/IYw3xc+H1m2+SYjENrrp72DOHemsdtk8a3KIpIWY5CZLM
w2q7FeRu3q/leCQ1n/3R2vo9OI4dVnQ4hOA/gl+uMwjCGx8AUcZY4Sqn97qGcSvcSy76bQv8P0Ji
kgFcn0FL5oqT2qdk52vKfoR38MGQcKjlqqhdYAKW8cjjgN0pXRQs3y1wxi/voPJGZrYBVfqKB4A7
cxTlL9dwMUgdKwgnKaISFzv7RqAZFLjFNYrbHL6UgtLj9RqpnHX5B7VaMV4NH9llbk0ulJbbiooK
zSV1MKolr8nI2CBfi3N0JpaBFThypZymnn/KOh1fTCxbYMmtwVZs2X+8CMharJveWzDC9oU3uwyz
ChnDzfgmcOgdm8heJ9JKeolMrLneljxbfXmwtdW97ZSwKeIewNpRRG4b3Ejv/cG+L/1dnRlr77UA
exy3s2sxSACHg4JT44X+qUtloUWVwliJXSNBcBzhb5ql9TBgqWjC6efEmSS7AOa9JDNT96SwqYIN
irRElo7LKLWctHpFyDxIjYCHPdi+v4GYbxAsdTELD7NutQOkaMbn+iZFek8I4ENE4PXZr9WvJtvl
NCmnrb2vgTzN4r2FekVs1nxOaIQ6oO2/zzFi66K2Shr6nE0xY5/Z1BZT83oP3fXJBuuiiyq8ozAq
WR8N8zP73s9WFINqwcrg+Ixk+bbXtQQM/P8K/+j7a+lzsGDrJal/2d+GNdFuLLEObmDQKOyJ0boW
j5wSx3OrgYVCZDda/Q9qRwdzDs+DPU1uXnxsZ9+lxOVZAs3cPL3Y2J3RJhrLHUZqv5gGn9ldsr8h
FZqJFa8M93VNxqgmHUcuhdm6QVDfgwdzzWd27h3uTlo8pT7CMXMUD4PQNFWO9K/jPNwjzmUePNyk
Sq2mwAO9p7BLA0zFdFIm7J4AN5YQ7XlNOcJmuXgedATOT0aCGkW8b1ELLjcbiq2vOhFq6wS6rU9s
3Cu2c8D6mKhtX9a/5BEgJ2mcattkyis6NeRjffmH8nxxKMfmOMUdqvJ3DJOCvKu/lSGScZ5aT45m
gbaJvoBgYQuc2mBPdyYAuZN9m27XNDSzs7ex++bPyvqE/+vOGymCuKZdWrq1GbplsFV83ZgYu4b9
nIQlwC9LNGwFZEcxIy9NGPJwfPbyc8hNY+3H2mwN3F9TvTRwfeLHkcbhvFiLs32UpjN6L+X32M5P
NIs3Y0TgKIO9l5JglYdhh4MAqqX2QR/Y2gyqxtRbJkBI5rLlDS3MX59J8aUVfFg7ob0lGvmG5tik
RpF5lA2Wzj74VyoBzx7sPmdxAKKddNMZRcJxk5dieD11eEceX7OcmsWHAupdXqLpD6XEVylcxfhT
XcxaiRHgQLOHFdpNuBV4gk1UKse6k42UIME0t/260ZCBx5OejV73EUGVaKHuY9d34b+fNaUalYxn
F0lDXt7U87w7qRt4War10ls+trTML6CbQF1qqkrKl35+isL+HFDfufaPT95lmhyogdZryngT0zQh
TuyDpIcSKpNFkTG4kBlprahflz1b4Ij++86Ys4KihpJenXnBh3zJvCNIH1+uIgDw5A1A+FJ+1dFQ
VPy4fpwp3lSWSvDUeBeavYYamEmsIx4LNEHdEomgYx7rtTHc1lAsvcjSppTmrDKIv9lklhesveP8
HClAZSAzMt+FHy/fZ97TUbBFz6bAwQq5rlHWixnY9e1jyJWK8VB0DDlHFaBn5xBw2V2s1XjR3lGv
byYzqdrNiDABapnkqX22EsPAcgPJDCE6sHqgQBhgZK3R1qEk0wS27Xa4ekIjxD4NLr6MFOR3qe8D
MRKqw78cjZue9GknDOiM79CNFGhZ6cJgNt60tumfKGWS2/kEwGBA2Oj7nAg2YNS2I3CC1RJJMHCD
Ab0MByU3cyVX8DoxK0wcTlUizVgtnR2kXyHHRJnSSf2tebSbHM6tGJ8uSXzljuUkrqy0VLIVIody
tYVMuFIDEJSGcjmnv6pya/TIe9x9L5j0/J93upKs3dnQs2lvPHA4VAr2SwCGdKcJLkBow7C3wndl
Pj3kmOpPqetarHU8EjkqAe681/i4t+FAP91e4NsJMoqQ/OI5NbgfTzRYNuPc0i/XmOXy3B4ipiZ2
gsBK52l21jWUJjdsCziNOyzarX1HijT/Rhyb2yd0ddJwjZibI0GbLFDO+ekRTDo8E3s3VAdkOHqs
+dWFHbAddxI8kJUEI362n6hNJPPOHMUIyQV5Q4x8BAL2WPBmrO7fCmHucdBZa/IQO2PRMGjw3vOo
8lKgibleCBtmlxaOsayUH7ArHSUiXjrn5ItCiXUVe9s7L8Zs9kdwqFaB2AoFTU1yzFC1gb+inCq4
BM2EhIE3sUrkNHAD4/Chtx/DKIWOWWp0XbRnoUp+V1xapYRLAEHwnQimBuePxUdsNn5chznziePT
MYx2LqLwsOF8R6FvTjRrCSeditl/0ugVaU/YFAqKL+R+0bc3hwMzpqYHQpMIJjFlVxJDVb7HnHce
L1z79VBtJVLd5Gd2dWo8uwZPcQSHVHs92kFzjL/gQYAXUjxPfBQe76O0vpNh5dZEm0+CvWgUZKg8
HyM9jwREAQzxmZZKaf/3ZfVEgx+08jn+kteh56BJiuJh/2ml+zcQMhEDvsyLqCnz8R+ROZeJMZfB
03BR+g2b5LmJiJlsmO8OKbyjd5sPB2Rm2YgA4ZT76VfM5XzAr4J9rnQxFzz86/C6w/0FpZU3/aJB
PEirF50I0cnV14mP85bcJxHhSzGqoZJuX04JjRPksi7/V9UBqratuvzyDsYeQ3LDckvbryamEIrv
Weuz9Q+yNGUlW9J4rH3h/oYuh9nPuaIJpb37354cwkpj3xv/1znxl6xj8zfyM8L0PGSHO1pkuhES
eh8kNEl/s1i4XwXJU9/XUDy/4Y3Z3p+z40Nk5jStMS3x7br+bA1S6fjimr/tD5Z5TX8C7+KPn9C9
ILcK1AMLSD8oUnOSk6eBgoce+wyZm5y0Am1v4iu4K8M4TFi9YLfRFY4ao8J2bP8OtAYg6pPiDqWm
kJjQnatKcFjvR5e5B2xOmSLleQBr723QS+AtnDIk7X9QIKpbns0nl1AqXgMt5mXNl4ycT3KD2m28
poHefToN1LBuhHLx2asnraHjY6PGhRSiodgMwvls7QIDQQfzzANKOaCc0g7O7/h2azPcQxbC3lNw
KS/KL8yGTv4xpsMyPN8f26xvQXNb3ih4bh7H6zkKAUvX4nr4XiR9i7tkgyfj7184s4YutfmdeX6N
yQBQZ0nBphcdHYM7GZLRejDwL7DDGl4z1MfiEJyVAiR8DOoVbF/RQngjU/g76Jb13kpw28gGy94r
q+waLfB7CLTNJ/9wkiBSNGOs2TQSwslPxadJkqBfwQSTI+50XljHu3Hr+wQeyO1jdvWa/Dy1l7vZ
ZMVRvcsp9BlI3iQLKNIsDUXpLyh1x6Z08yYIi+tfXahHw42SwUc75qe74BfI5Ivgue4pdglfOFR7
zWIF+crSaC91gJNBj+GEEk0/Eo/atHiF5WAUtCKu3Mwcvm6MFwmStWK4HMvDdm5N9bGxlHaCLv26
xVGFI5AmSIs8ScNanLRDBBvG6PaY9fX9HidC6fN98Zvor9/FHxcaWfoin/EF7ErUW+t5erp6Wzmr
fNQFIzUE+j9v76Lnd3e+q5jxvhD9usy6cPTA6OWvujn1nWCw3GpgZD6ISdOCkQVQxQBV9BFyZ2fS
oQ0UvDNkcLUHAo3NKFD4Q1zguID8kTKBMfqh28EgSPGUWy/3Xe1V3oAhx4P0SsPPYN7jPgX62IJL
P8rGD+PQNpmeKdlXQ/E0cjMOKrbRc6Qm3ivC7DyDfAMfLPpsVyshy0LbAPYHbVTIameQV33GZrv0
glPiEzTVWqySxf1W3VCX/KCnPf4M8jCDqe+YEphyTb40npbmogQLVkn+kHQaWfX6Ys86/3cdMmOB
Iz/dyMhvKm+KKqJYG4l9rBPRpANhVresi67HdBmaOCjKtnb4W0Wi7bKpbTmScvj4W/BZzj69Vp/f
4Poaw7ZrbuIKOUf76kW8CXvMgr7Apx6njld4wwS73SJKsmGd2FVr4kegjGfxc1hFhD7fhQk8Ogrz
VcMVvbWv+vym1AQsTOkItjEEXhowUOGCNeFEcz1fU5k6uIqkfJG0hCG/QhtORKIrty5go27jgmRZ
+gGabX0OMnVes5ClDYb0/UhUh4BrG87jnjV6CYxvHyMpiBd2eFK3CreXxOO6RWUyI67qR8fcF+SQ
sySqEqKBfDkbgJjL3T7Fm9h8FJ0zvkHis0Jfz04opdQViXVvAOnoOEVa9YUc2AdOji+u2vOuq+W/
niIOgmLYrEVonqJ2jPFqUml214FDwi/x3g5bD2/eyh4lhnZCd6yua01al/nQNyj1R6vsU+GCOGDq
DuwNEozL91Yg4Qfk3hZAkfiGpC6Oj87YsALgJa8HteCG4JhtfbBBuMgQDlvk/yuwZHg33cVrRZW4
gNAeYpoDfwvglDlDUjzoITILvxWEDooS8vmJ45TPLGMelUDqYv3wpMU8fYmSy0/xj4G8R1bO/+k9
6EDxXRoDV6er5CZZqdQLUGbMaUrPZOjFYL7tA2c+kXLqY/6D7MZmKS4E2c4i7kSPyQY9xfgAWLFJ
apP6O/4u5wwCDk7eQXOLNVpMyM1kk4/ZjmXiHIyYkVoKHKp64XPiXtg33Z7kdD4o9DnOXwLcfVC1
a64H+bvKubxkxTuI48u2UemAmsP066q/rXOwS8Ov5mzW3al20LTWAaB3VwYlGZpZyeaQMb4AOnjj
Y2Opqb5KiFUh+rHtqShBW2BkCCBFJo61Qcb7XBZ+TZPuINFjCfx5m817Mx8J2HngeYtPFlK1Fv2E
5bxquAu66mdTK5tq+I+XBurh63HZwWVN8RI7+m6JZFyD3hCMTvRQ8bOPVx5CI8r6b8JY7SaNbX7Y
X41X/8FI3xybXeN49PlnVJmd6LOP/ZcS/X7EB5NaUguHD26/s5NX3b0uz8IkD1nDEaLDEwRbgysp
b7OXLHLoZsp69F+rfU1dr3/mMQ38lAQC6XyWZ7SvOKeS+HXdiDK7cjEMTF2Y8DSnspS3MDmUks8G
U0832oQ839gz88ZXE5smGIwkAtGpcTR9PQRajW+Il1p9D0L1hvIn1HLwfFWHW7Tk2aRdxC/MkYtP
0but/GnkfAYgh5TANNZtMsXLvkmMFUwhaZgDZXO2Ed+tZ+D2aphc40AK7ZzeJDrhOz5SGcGPtBGG
BaTEikQKpFU2BLw9MAmAyKGBRhHqjhQVh96/aPOHD12YSFkkaNMcT2Yz2clnuxx0ACDAhoyxf0u5
PlVyD4g+K4bd0i7wIuyABkWLllrqHJ1AmIdRLp9bF+iE5OsziCy/yqbBuUNAT4gH90sMPIaAJUxI
pbOCbwkRjqFgEd3S0WUGtFKa7W+2+RwnMrSgsbUaVutDkP7B5N4UI8azAQCZH49pHgtRTRgbwfIT
vZbTHPEgrvsJ8B80mL4bqGgsJ4A1rmJYTi/quDGHQKpuHFccZnui715iCjkuNHjCKMrWMZbnGGT0
vo+QzOxb+UcxHRi8TlE0LZxkaDVZJRoA5NhseS64q/ByiXkoFBPhXlpGEYUj8u46OBZNRfdtO6rZ
qFojVSFV79MhGj8KTRjuAuC0c5dHu5Fe9h/2vkMieebkoDj9nd1P4OewonNWGtNGGhigdDlkz+pX
5HAyggZFZRvtLAItR/jYy6d1WHyp48EXOP7L0G4HLQUtjLNWI61c8Kcx4xaWZfDlGlXpPprfuQJm
JNxMoFeWh2SNoPPgxI2giBCSSd6Io78xzkdJJpd9/M/gvQwUG2t/xEd/ZBR1EKd5OmJFdjfWdXvE
eQg53XH206HlugTmUnIG0fZlDAhR9WHvIMggeqS8DNbQA0yxybBV5Fe8rEtuez7T2ihjHAdbec4v
S0/8gi290rL6JPqJs+QJ+W0SJOzZOVWidpkYKqjDcodlx+VxOZA9sI/Hdj7KoxcUvqAQyW5oqI3J
qAT1S1ql+Vf5BcgX/Zr4X1TDg2seXQ0ZLxAyHva3b2e0uuK15+Ilj4Qh6UX2NNGMi7MjICUAO3BN
x3RJwmXNGBJON2W3k3d010vrBCmmVl/TUj0NEjqM3OAFHyOpzjhFqj2pSUiU3ptYby6jdchJ4eJr
oTMBlOZOHIEINkJnj2T5hZ3dV6mZxCT2R9LW419Ij+fT/BJ8XDej1Ni25eJxMUJibX2FPwPpz422
fKZnRzZq1mHJ8M1XDFO9bCOiR4xnwcrj09bVxsFDFNmRY4nonTUFtmPMqKRFigPyKMPTK0Hw6hy+
NyEx2Zmsr6EwIu1TcwYORvwDDgBomn/KryP/4+nv7OG074bM2CW02kkjdV/B1Szn7IKXr7S55zgE
RJ4LnX/RztpuAUUKXx86pzXB48cQ/VYeGPA+5dBOvKKZ3DqKeQwxqZxEpFPm98FvkH04JV9OhGoJ
25Rdei7G4+C+Euy7Ofqh4E4VPuZ48HRN416HQRhTywSn1jWdXePFwJpCpZPgWg4Xtkg42G2As6uU
RWK4LtCH14bHIAvX7wHVSGCfUzbcexLdNRJzKVY8aUZmmPh0pFCiyHRL0GB0Ya9aguNkr3SW28Ow
4OZaJJr38kaTkMuZeVgKX5OKL//RCzd4FF771vXf/Prr8iOal1/BtQlZvo2dsqu6bLpez5caISt8
BUQSr/Yefx2KkiatfpGJA5Eg/OcU+ia2mwK1XkGf9vAI6Vk/RtBShCJeTXlvER4EMyftdoY5gXS6
MP0sVMMBqKXkHrUYafvswXGHzszYIBou4HhN2lPHZZvzaVdkaIZ4eVUzolWQ0K6JqAitC1FjUoA/
exy4u1M8OsBDzK4GRSnqMzqBlMa160+CAvYlaSomCfaKOppZKY3zw+0IbEB3L2OAr35sJa/qLTbi
iOOj0jpVBmn54F+8Q0cvec7DjMSXxkGp5lsQBx2+LTjrGa7CQlzjEVzssUTwlPhS1i0vW0BWQYPb
1wcCkxSkgno4ip1caM0wo+JtpewPnQdB+8GuW/xCou/6CV50twtVhjtaFatDLD7AeFYATG0/sgxa
2/gHK31nUIHk5/PPLlFkR/pKEIJjm1vKW1rAzMb6ZJj87jD6/SViGIPZ9L+2oRQC89CUJYD8ozR1
HRfPkGo78Lixo/B2nhKGQbSrQNRvqnKQTVF9YRHsa3QQ7XjIXDGLJQtqOYyP14juQZuA6atU5SpR
os7VBJsFh9rlnZ8tRMoqgFhm91zuKtRFYePoz8USBGPp1J/aau+iQUDHn0iR7ee0tpxYwrLscAR1
Ja12JkKcdcuSLJy7UrFiWelT3BOf9ls3BiNgFz2dDaGqsIjD38dERikPFOO42gf3L1I+Rtisarpc
jZtYi2G0LegxWUbRzKxtDehPcJF1Nf06pYH2Ye0bBwKjBqBHoN6aKNGjOAhktS8B3jbgLcDQRR5l
6fTup06zZKaHxaabn0Pg2gnH4Gr+p8ULLjnXoDaf5kpmV/rFFvo2f/OXgXFn3o1kjDkFrXytrXAL
8WTlFwEl1hpflQpOWfUP13SBtTkHDNL9s2Ws0BYelJhrvcZzEHeWu56nsXak44Lq31dKpHSbrEwU
IhWKxiXb1CxS4kgxAvcvO4Ag4nezGm305OSzBEfyhCW3QcjgpH88z+ImXJXoMMX/iBgWwLKlXTYA
WMtxNk7WEOKbZ0SkwyYU9BmffrlpsJRmuVfi6w+hn0lJ1fT/vf57H9gsIaCbw97ipLn0IU2YzgQD
wNCzB7+4qi+sHppzHSuaTS4+Yf32gYmjfdPlQ5Tp16A1ByKUQeDWwJyVFoe9B/bR/G26Uifr9aX6
lwRyPu73Ypj9hOHpajXtzj/zrdT3RUdicSzwEYoU/GvdUWfMeEhRvv7VMne6qZJXITeTe95FGSf8
dphxnfAE2NUkjIMk+BIcOcpTij/vhO225GvLPNka9kQrZQ+vnK/FOGC7X6Ub2r7HP/uZ/J8lxdTA
LpVY2pr8v9Zi2R5OWd5R/h7eYKL5SkAMKbovLLvGExy7JHKa+9jKOfZ8chF9a0mk/U+wMwdKt6R+
z5ubDebDGsf37Kr9KPU3Hg/W1jEPIKmvrXzcLWt9LmnwXNj5ae9pqEgJX0UW8t/baW8aOk2GWHB+
czF9WT6n/BQ3AMfhqFGA3wjDzzbZdXhTqWa8H5JQ9K2Hv2r+4cKh8uTqf33EL1rhnjx5JDJPs+mx
GU4fV6eK4h5Mwq/Nvj6GRnR7P+jYVXnB65VRDm4nMyK0JDyF65e54ekGLXkGdU0N/N625m8VSaEb
aUUVcPaITaQcLqvWyjPl7nLNkXJyVJ0svxq9n/i54HwMfRXgAkFmZCUBkRSa2QME6K/L4P07RyUu
MFNlY4sASTuksnSUBjJVJvqxTZkNzr/wEex9/I0ycpRXiKnFneq43u/ID6qk2t9ykGKnIaQ7IAF1
RB2UNnjKRutrNlhjO/DAJ5JgsVvdvknxlEccZAV7eIZGee6qnP7kRcp/EPpLd+ePUmzmUFOSkENO
cSXayxRja+gVENF67xw6O4vVH+5Yjx231ZiN0LTFZpt+wdsVOQVznxwCGHjhAeitfX0hf/z7reUk
oEEL9Omdh0eg5thz4EHg+eTFlNjbDGxEC6atdHbY1lUUnC8ErwNgYSdn/VZlCMQ4ljzS+Ln7vIjI
fSvHKifB9HLsItximLh9SDJ+Iga2vxx7Yh8fvVj8FdVt/jUnmN3hO3/6rU8/CqR18QHuWfVyAAys
/Wra4ZUdFAWs2FpwvNWEwq+WtIkHxNmLV+6Dkz4gXCliw/Ywq8xJw7ZT6O9KaqkxpDQQV7gSuYwj
4d/LfW4VCB5aYMZxPwj9lylzCjCnqfB1hIVhwhb7UbfihHaRRG6rFt5jBlKanaRciC0ZZbqMvbSG
fkHGToip3RptATj6kevVjM+b9dZhwOxauLmf17oHxHE2y/OGXFMT9OV8g+eCG6AH4XA8SMkpyJvP
gTk7JLrWyZny+4ZvGEjqFGKPAaoyNixfS74SwVpGgg8l7uy7ZvrLnmLvPP9VRVQda1JhkzmfrjcD
vR4Pq1LRHuiVQyz4V/RyyQJnHPZxlEzqPKIjmp7Wgl6JWdn+QjRQItYGI7EJ3/UV6KZAFVkBTLMg
4R12o3lUcIcd6937VLu/y8HX5srZf/bNaJUyy0Kf6qiq4MwmEBA8Di+NcK3+KFZhzffmMn1eObkG
NeP+p3+HZGH/77S2cg+HwVAKVS0Rnuf8pI4VgOek3pIOQQgyzzoRIdSmqJUkrSaCaLq5NljccNvY
6nAC2uItFo5u4rykSUng/89dSMLMFe7wzcsOx4FAE1uK14oZrmk9SUMUjkXzE4vywHCmnB0s9u5G
1DsDNLbk2u5xgfYKhLPuHXeLH0B+ev/zLLxTYF5jqCvIwnraHIuNDueLf1zWH9B8d2oIYs0PQf8j
QugH9ZF4CXPALQKb/fQpGlpydhrZsouOfVI/Nn4vXeRepw9rSPkUZ8l1V9maiM3y9s6KSZYoJ83e
0RJAN4XwVWJP0GCrLhCzYE7ADkqYDZzGiprPlbTJr8hpnmStlod8I+OIy5e9nN4dKP0owHDjIeCX
bQ49OG3ntOddJQOqZqd5ub5tRo0DwAJYJeztyVCL8/EkarKbdPccO1wSIV2St1S91vMd2F396VFq
dSl6l2dQPpSgFB+Ilyw2nshc4u7owyC7Uj4JixNO3yLP2jSX8s9X4LxgLz3fqW9lpJAuSiVcbydo
k6xV0z9IOkz3ZuteCSJBK/5Q9e3+aVOflbgCqKlyJ8/XZYHzl05MoR4FYaxHoM6jaUdTzTQownw1
l5DAG7eMlXUWawIPMYo+AVEfB+7NHzer/2YhW0ZYPFecLMAmiwHgeHaaCxk62DSQr58EK8GQhNO2
GmuNGWshy124Z1Bp5c6OinCcA4yLNbwFiXuHVqNFXXibRldUP6E7qgb19mI/SbYZcsr09WR7DWbz
PZDVDf8J31QINvOFceETl85slwhxrQJY9JZSfkQxYDeyjnvZXLlbr3zMzIIT6r/YA0vMxKSR63uI
sJn0KtXwPZ5HjA1BJ7sea2cNmw2DcgDV8Mk5htpw0mM7se9ZZbKZH8UCFmcUnp4tlQUZX5ncksvV
jEXL8r360pY0f+cmzooyzvKD5wj+G1IB90l7ymdj/RCOWwWvxPZvotUjFqlglA/C1kfByx71Y8Jw
BxF8hAP/gvdFmnvQqKmoUGxNKVmOQ+evxmFgWebgEswqI7FRNTR7A0pBHFPIf3Puufi5k9xZShhw
nufiLRvsWV7qI9tMRRw3LiBPSchtP+uHMl+3VTZvaWj08A1zcLg6zdi46DUnqW+6hcRsIgxiLQnt
YrMxTsj2gCsteqnYXSCgLn/tRibF/oSIv7wu3FFrLzSEoaXeh5T9AugYVEMs2OqRpXDE0qFNNQ48
0r2PVieP/fKZTWgShASHfK5GOxuPdUoL3Mrpe6Xe4vxOcGeKJ6mIWniTdqTzn2T1+cmRS/4NCuYU
KdRC9ZPH9KkDgAW4aCEK5VTMvCGIebTHM9wEL3CvTuuCHfTP3udTh3Ha/t2GQdf0CPRFdITymc/m
qhnGiW9TlzcI10rTBIxETrAStyxGnBQcrEL/3MkAVW9jNHu8MNKgZwLnLW5cC6yqrl+eaKiTbs2l
6IlTvzPhv8YAxsLu0U3qcq3M80EAyS16a+jPPWb40unFuWjGLHcCkiVJiBFa0SvmTCwPSPD46BBu
oIrZqkrBsrJlD3vQFReYtF7maEkFdRzFvCRBQlgBuMAZaJbdZpA86FdsXXo6oFcD4uqMjqe7AcS/
SMTOSSKdzzWUv2Sa9hL2jEunwLh9WhgqS6hqnwkSjuYGq/8796SisXWoAnnkaKP9swBcRI+gaeA2
wHadENdofqldAAgaUPcBD73Fmtl5ijt06OhuDBBdtpjPgxM+hsM2mJQhEIKOwuBGidfBBolWkADV
jyB56kEH3WkAfTQzhtMOnHNWT+HPPI5xg9Wsh9s3TTV82rvk+VPkYHZZW7ig1trBxYnuKq0jZ4a9
Sbe8xFkQsf6oveUDJmPxNKC2G2I6jb1D4j5lVoeSzTU5IZd065V8JRmiES8oXIzTDGClKWgFIDew
+84smW8QksS8CDQk2DGBXPU+uOGmmGqWD2wLDIPp9I3ni0f7w9+E5tTyRAg0XWS9Jd2kn+0wKRoR
+AfdDnL3i48o2+w2TlE6s76hxAS7bdYxHPGSTEDn/zmbwsVNt9yie6j75Behd1tIcSJLU9PRd8O9
wlQ/3Iz8mfvDws5m22A5l6dZvq1wOF83ILcZ6CQ/vcMXO065DQ5DYK4GsByJQPFT4cUaViswmHdZ
JpB3DwtoZy1iZQ5WBH9txdqkxkm0lptxCVMy+JiCzfqkXNwpDtZcuVQ5Rit+K7Dk2vGsgHLMLzOP
G+fLnQdUxOyvima+Sc35wVKY48IiNk5RpuzhCYzhlP8u9XlrkfLi3W7hARGBk28v49qRXW23LhmE
7L788mJ5vMnSO5RlBF/TVQCg3Nux4a3LEHfJbLNUu/FibPn813E9K8kfTZu7LTEWP+OWrZwiccYf
TnWxM+g4dfZcgMGrBymcZUMPKnKa+I7WFLilB+VNCGjyIdnp5FrRf4RJ9IXm8iXH94Nd/gKw4jSA
/fpgW9lnVYjHLRPzOmq1ZNIXDhnEae2MzRzKAyZK8bULZ5PMWUSZ4I/0xx4Tnymsx2UeUTJGY0Q3
jg4MiY4xaYGKpBcFq4hH+rLeFUDdJnAbV7eMeFs0ffCsvFqjp/ZCjRYDZlSFzegryv2rgyE7orMJ
s9vFAJDHv0GeER+3xSBwkFNhVCIW/q6tDwqxhE8Vwfzszl90JdyM9BZG6kP/CgTZD8wd14Mmoib9
IeEvAQdoIS6oyJS6HxrXt9bpEvgUX87pt1pnpGKR6I+8owi28s7hQTt9TiCip6t9teqQerHZRa8Z
HyXsAtUrMjHv0i+eTKadokLLwoqHuyxOUnPCjO+qUrIVgR+d98wJ1z27sniQjHyve01SZsNgeD4H
VQl0WvGCkSgPOZ127KUqOcun8s8oUL5PAv7MSXiNI6gmtG3cFfwPprGukO8IcFmDuPZUXeUuuM7b
hq906AoKmwxiltnoiLLAqQa/9fojgFYsJLPoLnsL6qUfAjYsnZBj0tV3az9LIBsHPTfjm5ncjS+u
1r5y/feI8OYKk7nnbT/2TBKMivqLF3DtyBo2RIhdQjRfN3Z/RtkrwP3P2PJNhhdqzvK4+94OhNIx
PuAZLy4wyx2AtMfvrgLwIC8gxbbG8jOGwaXTMjJ4l1zOyQEsl+kycqHfCNB8DS+wJZFcuOuH/u3y
023miNSGiSbwBh8X3+TheHFwhpz2S955YWtIoADRE4yr0hNRIyDI4yNjiP31jn2etqITqn3zGymi
Qquz/PgiGv7gU55ZathWn52/PnlaM9tihWrHonwyF7SfkNaKdWFYRBPT2GNoAEjyLsuOWLKgnL6a
U50zLnLqP6TJW7J9p+7kXsULLMe9M1vXiYBJZ98z6lx/Io8Ncc+GarJpERbxqIN96m71YYttKlR2
UYOgweTG/VGdZOsicjA38k2jGAB0745GGVKdHLUA8d/eVCYG9VLPiyCL9Xl+dwvLFgE9xmAtcnAT
UZWkoPU1Unp5xwZVbSmFEdIMrj6De7cZ5Q1efKq61fKY0466PTckhCp/SLgai/5L5pA5rx236ssq
0TrHLCL4KRAuwKpQM52Tuj0PdOYcLFy45Q/v3TYD9/2vSoDd3RxskumZ1a0HsYdnpFIScfXNy1D0
7KkJJQNq1SvTL0Zo4x4CdIeGMD3hP5X0xsllUYRL2VnR+fHw46V77z7d0P7muH3swQAJSOnXVCJe
ycvvb8aAe7YVLKLwvOOdA0GfdsK/S54l3b1rX4LxtBCK5cNjIMM44TLk2bA8UAsld+2ScYxuSuc6
iZmOix3BXUpceRdaejfpOvuDkebLf8drYbpbdeullqHMMQVCA11ohKP6VR3j3QULxgizXWe550+C
vs3phP6MnWI5C/ftdovtc8SdA/aw+XmLiXD8AIRgk2aHtp56ZmREcoOXF2yKeJwNiRaWzE2mLNUu
2abt+sI3vHrMG/5Uo44+nibdPsEiINapoPr0WmyzlfyNmVfY7idujutZ2TrmDumRD/VQTXakxAQE
eesXjFeJFAR98Mmty9E9kCJwqj1nQ/NtyyOdpXjsBMih1XnO/KF7hQRwFVxCgwMKz5xxOob+ktHU
V052BOrcCBpUpq1Pp4ONyRfl7CkZjq+kn4MYPuN092/CdwDA7SNZ10SvT83gwJoVLwPxsVcY0U2B
3+85nGBt2isitX9Oei0X9PRj9fvmd1A8oVXBTo7vr/Dyc0sWfDv7UF90FrPpzv4RyjnEY8vRpzSw
IShBd4Oy26SlFs8+pv86fRy4XR0xik8a28neeQ/AgMxplDrSVmHzUcrZEAPhA2lua/TlLEJztIQZ
/eaHutZhdr4Q2AThXV+y0Ck9UuP6mtqfi3bFuNRXQPG863JjJbHpqpkncoDho0GNqIVxM5W4yhZe
MH8+yY+OzrCa5X5nVgskeus89V/whBfG/icrCQFi4jGv3vPMKDaH2acxoivx3SwRZA2SKRowvDAk
Urr+Iw+i2u7ox/4Sfk4WoMEPTTrhQyC77ydXurG5zx08D1+XmFeTYU5J6wi4T60lqPt0mRFCz9hz
PJdsfiuQ9hPDBnb5ic+sEdSCsBV+C/HCo3B4IckZDfyQ0oAysUwWtRJVrvveovhWKXI8UjPQuRI/
sMcd/yCqzpK2y9+Emf4KMaHGwudbhOoE72ap6uT0hOEpF0rgg3flVp6rZJDrzRVFmaHGocUVniyF
94mhyzu5FayBXF7mTI7s8cwRkW4khOwb3DDYSncMEetZSBnGoAliO4uOqPzD1y73oeRkR2yWLE2d
LsmdPH2tnySiIM4Ph7u9hamQYCqMbbjN90BlwODLcuD0cf+g9VUYliUjnM25cvh7RKNNvHfOr1MV
kzVMMjwxtBpvaY2u3/DR2yFRs4MV+jhW5eEKNBVpqfQft+9BhfTuibjlGmthg+5ThU0gOWM0IHrB
oQyZ+t8zXKAW/MFC5NPET2WqV2TWK1FEdHZN6I4CdOeXmZOioHlQG3+abhEod8bLY6yS8kH8Frte
ksGS7sDdhbnJdX1/ctUFXy1bYfmiIe3iRS5so5uKKdgZ60sDh6vENpC4FUUXqmVET4LjCKOpkGc7
M3UJ1Cl98S7vuUGQLf5wqbyPzWpNMfx2+ETMbYi27pHlxLyuHvJFFo8pGhq3807zN/dZZlbyEYUA
Q3bXcgVJymO541aszDOH5isZ3JL3bGk4yvwpBcz6iB6OIuAg0SHc3V20YgZRpjlYgz1F+Gys3+ew
BP4UGi0/XdxO09lWrymazfGFtoKP2rlt0BWqnmoO2660rOnrVKZaRa+aIYY24CUUFOOUpLnFJowO
3H9q//r+yjY+JpkHk9dyloYJjGNj14ywr5g9wk5gd3GBd3PYQjJ+zVhNXiHKGN+9XiDy5K1RlcLU
AksPnoxE/wE/t8P1piq7eRPmVmfjqhNz6LCOzUCmmUWoVvaGaWoWfa3uTSz1HtwTW0F1uFJp5Zsp
PoxoXVHb8FJsv7y7+Skou2ergs/maTF072vAYH9NES+q5mKOh1cUH3sPfyFiwZTVDpYxDrLtfGTS
qVWDmRkXnUbcjdg64didyo9SoTAgf2hfwXHsarJ01BeMPrYEsSaSrZIBuXObURkT89cevyy+b1Tf
H9sECbUcPj8J/K2Dh9vDY/FCE27lBQ6DRxvwP7gFyrQXJDkE9Jt/T8wH85I6GrWPccIaNMJiPJba
iuLFvZ3We43nhjm5J482mvqqwWAQ83d3muTfQrFrZkCnpnGEnZRtIoi37YtLYnMDgBnmfJRXGaa9
o1p0qdjWe5VD2/qYbyb2Uc9uAvJe16zjTd0XLtyamW/YS1jSW2JS09+wejLIp+x2bBQGcFAiSeFM
ofqLnksoGZVj9vbPQwigemCXbIwd6B5cBBg1uMRzzDcBEm1RO7hG26UMGFw5ukxFzdysGyTOYOfd
KJQxZhRiE1lJVNUH9BCDmP4Qm4zSwBUaGrYtDfZbGgY7tAFX5D1ROu5KEuDrnYKJxM0ld8AoF0sW
uQlrfM/HV54ByOqWVUkz31rLnI42iea5+KvSmJVXpifmxmw/IeF0ZTmcm5vw/qWFuDpYzA/3KiuL
ntk5gZ4k0kVxn4ZJdxJY2GrJu/betA6tq4gqz6lRANkglKpsIJgKfL2Ri4zDw7Vw6cmSQUUY7ZF5
qWfB6nUdMBWBg55y33CxxznJ6+eCxnUWkmz16X5x43Lk/aNqhdngvqgZjF5Dt88yaE1wlRUT+/Tc
eA6zCBNnnwyD46V/cRSLFpFoYk2MBon1n7T29YonIgczK+gCKNr2R0U4aep/F/lKZ81FUnJfoOeF
p9N+gX1QWnaEiC/MQNWed5+obTGVgPaf/7imwtEdvQnl8ax//n45dYVname5Jr46hFcVW8+WsZCW
gDTZWa+UGRwkTL9oP5B6qLsB+ye/RKm5g0OoU1yt07xiQsWT+q+tLXoLfQ/eb+K79iawiTA9GWQZ
sPHZdkBpMN9bXSGBnS+++QoLwbsmlTxYExUYbNWF9vbMj8xoy1pu3g6M7LfWwijdsjkxhxjiydY1
eJjdjRHSV2Y3NnxDXee5DgL8kZP3CeZSu2EHiadZICeOgMToZZ7U/hSrEQQKYHfndT5yJUkhuB0o
aSDTCvb3tgaHAGpwjqeJJBkW4Dc4qrQPDSWQ+FzDTKDg1y6hX0QJe7OadkiQDxnT+nAq7B6ZJTt0
91anPvdM3PYezKNxT32Igk0+CwQmbLMr8Y/m1x0MYmSDlTq5hVnKKJ97mnrsK9e+pJLHn+bc/x4I
KXgfhHwLj1l67w3zXgn8NR8PuclIvFuqD1iNSOjJhxCzKXdPbjf2eRsBINgAUbU7LoyVrP+ALoif
Nh+R+Wa0WiTyhLTuPvM9SLWKSs1AQnearURU5/OmBLXT22sXlfDiIufCrufH4MgCeAbd5t2giN+h
SRGejCJL1DICZS49odB9TLvrhLFzRdjrRp0GYr5xFtEV8uzlP4FFJj0DRvf3BZ8KEy9KnLY26Z9h
auP4R5azYxUiksHNkab1+AAE3WwyDiprGqxHwG6IUX/BXUnDHeaEvm96NETavQz02WhXlevgY1f4
rqDmfBHXsVxi21GnHaZk60PudxeBQZuPUYlrqe1gmUr4RpB3RqypXH7Nuk8j9dBcZrFNbkt/UePs
SjaMxQe/a/UNpJ0cGiEcgDs+7v4qUALxPsa9iGdjqC6bJNT8yPuQ0sdfkLsWnGvuiL0xM5ajjppz
8B/qdy9b+Nfkfh4JjllVCs08GuD5zF7/0Ip0cs09YxCpM48yRj17E/J/uoqkblVKB8un3Pa4hf6+
pw6i1653WgK590t5CIiHMc85REDmwfmvmbR2WsRrKPwClrxNekOdD53sGDp5nRSBTwIvyiXWjJIi
LeTTHZPrzsgwGjkV7ADIAMAabmdBeBX5xkw+YrqrMkgicD1G22h2StRPBHgOv+tmDtf/La5SqOTV
QO9/03fuxxW2AJUQahBO9aT88LY2AUN0Tqrjz5DKzjDKDoYyltsKPHBSsRiyN8Ro5Nkdt265F+qd
8NzegTE6btPUNVhbLDWdkd8Nh6YUeDqnyl5xxymcj3f/KjpAeMqE2d461AnhynN4FP5q/copbHgE
V0xvrPOYXv5wlIzROkxSWh6XwfgemZXX8kThy43z1GyY0fFVhKDmWOnC39AcVFFT8WphDjUDAqos
5D6CrDTLhDQTmWPQybCqPdR71Gi35FgDdS1R54M9QVLtdCZH8UAZYq423h/F5AlPKHY6bqE0e3i1
9bEEDdRDnjlGQwSsCWu5MhEFMa8X/jdD3qbn5Pp15WhqpKz/xzP58TBHDFAWNaLTASG8h1mpaL1p
+Ab8snj0qNSR+9cjEbMRVypG9mLUqvgsQ7ZTs8Z6wmOfWwU+nrzDsbHxCDksVDWcoAOMIngG0eQB
vdsv2UUGg8U5rhs2IgS66YzxUIn+u/BfEgYn2Fyl/yKjQP811S69VZNFb/obY4Am+pEtEteRuJUZ
rlgj9ui0yN1r9JMCfloWJsGtFve1aWmvFFLKJbQ65caweGVnUYbgepVWgnOE2/nxnGZI7iI0fulU
ZYRF2ClVN6xLM47YfUj+Yj/iHmrW40ItOwDbD/Vc6dbtgjJ8CEdtxWvCBkHDJzdKioEcNhZWKMTW
vG2OAfhkaWffjrD8jFudyZAdMTF+j1FCoIGlfX7QwdZPzI1mzCHBNL29M2Bbb6hqkuKUwaG9iREt
ISySA9uQW3j9/ZzFbFRLti2Gre2y49MA/1d9+SSpy+X/BgsAG0M4oWc9AdNEsJf2hJrKRzrnm+5k
AKyqNNzvKSADLbmfRN1kVSfzYlqa4u0U+TLOJFDwyuPnjY4SfsnGh+Fis+KPQhBFq5v0cJU1OOcB
nRznksZpBZBiMkWYbkF5MgOUXraoJjd5Aa8XxpGxzZjZ9klEpOmLPykqOMYhYV7Qkp5PAC1vI+HO
AKg5vhqGUxXOFpS+rJRFHr9IpCGEC5iQFNf7FFOfaRo3WLzFhdgqNYMmm0GDzqkY2jwpS5QFJ/fy
bFvGv0VobRfXnbbVTtgL3I8KfciNhVfUp8trVugLUr8SMkMhTrgNKhaxs0GkpQfCRVVXpAQGR9lo
7OTkrIdg6/I3KE5u65+cEUcWQ/9gXiDrN0zsDVw/W71Q+EZf2UdJNkZJX5xXhCrJkPMmqDyUyDWt
EjmNf03ikJEFH9sGw0ZB8cF4xt/YD4q9smUWF9gRnQGBRjJGI+d9OuQip0PQzQ4ijlwo+NBI76X8
oRVv1tRBrfSspgyHrMZ88sal+FmqEmklG9SoQsTZwjb4mxPWScjiC6BnXYWwAVtmekWnMP2DuwCk
Ps3e+qTsxAzKwJ8Uta1ahIbbnaq90KJW6YzuYrtYxWPM07zJ8Ag8ALM9LjyRKwoon+9M2Y1+c7wa
G7CMgsXDTZb68fCwoJJMQFnxrjxyJbs0u1cWqc5FzGFubqg5wy0VqipMQUZyPa9+dXbIDulSfC5A
2raXyEzeosAIBVI1aCQ97ppE74Ph8UIcq+pNRCCBxmlnepkigu1nawzATl0ZxvqK8fERyYpH0Ei6
jzFDW0/0vTP6GH+bs5IKPtPb2qfm4mDwQ/xSSAoqLzHc6Nzy4KfepFz52yZ7Fsq1KCZmmruU8IDv
FyYGsHIVxgpJnjX3VNSeYgfk9/89cL/BVc9G3z7GpcF2SFEVHCK17ds3wHc+1siDrJQeuME8WQw8
xmNLCM6tWPMKoep7+CSXtOOoLT2eVJd96jJtoq95uE3Hw8dxEURg1sxkxFdywwQgxrQxlh1eewvQ
SX6JujlAxbnfdNb0/jAvh4qyBugIJT8t0OptmbSXeiUkEJw90UiYruSmsbWw/pYLfq2mdhVWymV+
SP5TmKUKrJNGr/CCoEFTwctd5dXqNqu0yfkUcGNE/vCWoQ6jgKST+abUJhJ8LILHMT2zaZxJEi2q
0nJXJvn/ofkryprhzkC7m0y8wZVoAvS/eqMvoiN0UUJ8cCERhq5xUGxDiOW0CprzJBphkTWgLBY0
xnMkys798ksymwsUn1m//iO/sUQyofTJo35j7GiBjnwWNcyFTu6TgK4jSIPmYbjGp2VFmxCXKXUR
ysY2D9QadzVbiL6IxKK6RcuHdrY2/QQOxwYANzh6cKlC4mxQ3tIc8BGJDg+gmWEc/gPXzGfVF9AJ
gCLKs/6raH1pTexjNrxbmwaVmqhKMyibsW2nB0Mgn/tzNlAt27z5RQAVbfPVyy+qujvTyt5OOERG
u/ibb14KDa7O3DvXphlUy1PGNlrw2NACnZFZ4UV12zXRuyQMbu6zFQuVYIWXnwtXZ+cbQkqE7zEV
qNhA6TUKDoy1syFekM5ZyHMFiPuy3Hzl+aY5Hyno4pi2B4Kk0SYpL0FJEydG3HUufHD9KVqkTTxI
4LIjB2O4I1S+UaL2sx4yfsD+7C/7Q0Kly/SP7JfykhKN8yAIX1ONSaakD5sVrFApdJs0a5Cw9kDI
IoN1uMX3CpULlyB3dYtTTDsDGBI0rz8yX2H+8lx9VDxAbQF9VdlIqXZVSaygCUhVXuxnT9DhtBY3
XoTwOnAKUJHVWh1V3QM99JbGefYzOmllPjtOLu5uuv3/56dK0Hgqd5sXiOIqZa8otxTgOiJrSbhm
n9r+xx+bxVFL/4z6+ZCuL4RStfZ9hUs/z4V5xtGt5fAJCncXg2etx66pqQ9AYhItneG5ojkJ98HL
dXq22N5d0gDirjp0gDrlo96zWOGbtvhfcMmIbbNzcJk43RAC0kLBiW5oiF5PeWkOm9eXsBfMAHO3
/8EK7WYg3dDANlUOm7gcxN8f6xp4k5Y0Vkptyb7nvC7k0NI/WfQzUQ+ORlXbIzngIQwWamNVfVrp
7sdzrJiLicKoNCJrAbgNV5/VdfDhoiqyKyazWVfRQMCxtLYmDjs9cBSM1cz0SRe/Ls8tpSQpu4vk
5FIPzEE3hV8q69RKSzEKSIe96hC6GzARUAMs7LAXCVGQDAsCBNt9d86bN8cAhqQwuNkSuB7e/SXI
SeC3K0IvqDzwQAWx0SjPuUaIokGYqD3QS8EbDiuQ8D3odRmfD4ydAIpeFmGhXxWxU1G9dKOX7Y/9
tfwXr+V7gMSruOXH5N6Of2D4jOJHlk3Mah9rQWLjkv4gIfmDj58uqQEYoK8ykn/jU/xlnibvt9QZ
peylgFnlvHUCtDG9RSwVm4Qsa8qNCbG7r1RmEkFwSWnfOHyT38Xu+KKYddo/cQO7wycvWXDJWr7e
OGPolSFTJZreFQohWzGOd3lUEtQ3Rb4QnC/n5mt/qv+rmT20R7mXKz2OEdDIEm1ctH0z7N63+ZK6
V1gNh9druobmLyoCO5jq1GoQ5QiCPcng6nqnCAWbo72utJQMM8q/FwXdg5opqXJvo/C3l7R+k1+X
LrGy1eoTupmvpig+eHGdC5sWwhD4LyrEjeyhEeXj6k/xOjATNeAAleEJDLuhhu3bRLGKnVv/WdKh
D8JkzsCa+HbwEVcZKcilG/nxdwG1mJzWJcc9aMrYIJkovbjUWuliE3TpK+jtQuYjFtq6N1WyJhNe
r5G7Pn++IFoXi2hExOo07g9MBLAMnMNb/r0tfm6VVYNG2aI5s3XzfDGrZHmBcV8EFqy4Z1EYplho
Yzw2SlBLMZ0WHyGw0Jwi7Dq5YHKFz6S+wngeJM0LpRczjL74tK+lHxFfigAnJYPZy6GaT6wEYckr
oCjXBxvYNW+VmCnqEncUj9ZLWhZ3yRlj924a5rrnx8ZIxXiUsowMuoJsCGSFEolaiNwExiNgvr6M
LuoIx1Vt2fTS15bhua5sMabrN9ZKkkEasAS8LqBhwWorwMPG2NsJl4sVdJ+5SaVvpZG5ljN1wvDd
02aLBKUCeUIe13z5ZoiIrAHCeo/QDgODfa/8XQquFnfkQwkWh3V5Z5ctVcUUjcMNS0CMo3MwZYv/
tTukT01wuJAuyZ+FTzTxjoeGxt0TgWXhlcCsqsPAfZgDD046VkGbWTn8Q+VoNgAiikYilY9frY9e
FlXOtOhINApR+U7lsAXV7Z1xcUJ1jzv5pqMRpOl+DBk3icyDrlNQJEojwJG18zON/dHTz2fgZAEM
2M1qhP95MY3zBFcFI1dr5KeT5UekUOMMbOQSjl3uhiyciNIEVYgV3MZTJcFsvf9zRAa820d8p6hE
5dXHgZAgaOiCWGddb/g3G2FLoVqkdb6OOlDsn6qtXjQhhp59dQaeeeSDPPW2ewwO8xrwpmyQYKSG
29FVWf39LoNsz+AEKREJh99X81jgJi3hgnVS5mYFUBdB+/hgo2r2rnz+Otrs3kQ/OWYayzPiG9vo
oRQLL6WONYWZqIQepPbh8tfnvGbZTfEzqMKvx7oc/qYBwhuCSy+kktDfl5Zf6HQ6wJZ6ikAeRI9V
9F/4pBBiwlodrYcap8y9FCF6d7w0/ae34SYnG8DtxIeRUKIsi1ebo73LC4uXKNWwtdBrv7TkQxGw
5eLj+A3PqrS7L6bCL83Aytnn5EVCjO7VDxkWHHs+QgfEYi7VRcM64JgyzNuSKJpS0UNbFWQOpSN4
F9e8+RpRDT3LtMXTTWX7YApbf/5SklggYQxMlnuf07kLDGRaE6ajosqEqr3QAsULuL7ntFU3UVAb
zSHVpBfIWdsi8AMkHnujBw3/2AFrRDOBghRvGRMenDqt8Tb1IOO6PV5sii4nMkP/G0ILcFfaaAJ0
zAFNETGIFdvuNqdLPI/AtZ9Yrm8Kew1mx/b209nsLXmuil+gqeTgA86c7sgbq8szxP8UfY5PvmW9
isI+yp8kaKld9JGqMSHtoQQ6J3HShryUczt5fgN3OtB2bLM20/XdyVQ3d6bxUspToVg9qrMAGSpG
FjSOBz9hho5J1ccQ5l1e20LsnlU7DdkVXKs8nAXbJ4o4lNpZs84IklmHeSQMaBLWyiHK/b5UphwH
zWo3XZlc3KvcgIeeJ+nTHhllLPQwkDKhnzexQfkopWaOQ4r6nQbMiLX/NK192pXY1Yoo3c26dyVf
yTA2G2X/h7mkff3CzmMCRDdht71R0uTzS9LrvjX/DVtS1zi464buv8QaqiIE+tKSyj+yjfgVYMHQ
lwdvQfbcO1doAhMmmoFs5GhwtMycj6oZXw9Sz1fjdJkRxOYoROAmsYqYelA5nQAShU0V3ABGQ5w5
gEhVh8bF1FNyOD8S2YIgh8qYewgatl5RpA2MQL3iK0cjEd3EWRi9duSlc2LlYiH9gsXUjhgGHT3p
Y4IAk54xfyutms3tayVm5MNbkx4ak9bESDGnR+ysSb5Qs0CBKsxZ5pti/GmE/8+PhiqOFr+mmMU7
kDe9SxFKdF7h7SAEvBh2yNqM4KIuhQKLJFL3lLaTFmQTP8rcYVEykTMBWwi06GQKp/dYZoQ5YqcX
3CGr1QBagVE8qlAruY65A71KxLeUFS9LpP332/DB1Eefj3ZqfkhnljQqSWDim/Y5E1TdGcnBaklN
SZa3LgE5rTwsXk9inxV9QTwSZp8WZZiQPHn14tDI4eJKlRP8jeJ/sxMvKqa/pyBr22U2MliytmxP
IUp2UntgVXUFo9Pn0+W2RjWN4nNMweMJaCQSz7SYOMa0sRhbwoscEjdcci+uRGtwYgH8ZEAc7HJB
YwfC3JqkSAxsA3TtnqpnMWLyR5HvZaK5sXLy1RFHxjZOILUKfQIAJwpsCrvicyl5p1N/h+LP3LfS
mh0LH0rxQG/P/Rd75mkLrfsi5xhTQMVyQHLwiriHI4fBBqr+LZGBj58rqzVNaMQtLedvfY/cVCql
fDsMoVT4b+IG4vB6mp4hSaLLsgHolrnAGeXQXB8bDnLPb8Bbyz6iuZHwWkdOgNflpDNldszOud8D
Za+MkewxsIcaVqxhBJWGfqKdWMEJdgGP5apRRsNVzpFBAn3c1+5SKUQCgY7g8MJIRGNKT+a4o7xp
PKAm4HsZZA+h2aDlluS4zTSf7YgyTueK8cEC9PSMswjIyEk+hfmE24HVbeDtRx+5wtA0KLamBgcS
ogZe/PnoWLmaediBnhz8/HzGajHVFGpjS4Z0dG9GMpvJXSnF0eDostfyEJvZMKl1VHHuFUTGdZVr
t8xwBg7NIrPTAJsfyP8J0t0NhsAMpuV/1uwMgOQhHUzB+7IQs4j81X3JnRMi7jmj7P0/drvYRU/l
OLQw6VxIA84NfHyBxnmv9VKRNkWbxipoTEZSDbwdtH6NQBBhexCjZuBUWXitJ80aYMlSYwy6ICxo
rUBWLiWDlipl8mcFEf0i6pEpPyKCQEuxqFnROrfrVg76L2fodk3nzlHQTlMdK36fPRV3wh4th2gb
FoIT2DvOgRjLux4TeSuLWKErfq46+h0pU3OhK2wBJcYXoSAvJHTAGZIeq9rXBH49CjAFED7axubQ
qW3SVmCntsifKHwhhcKNFpUg5CyhF/VKUxXZFZgGMSdB2sevE4pQXhprrQRSas3iK3wQoxtxuiDc
5RbQfs9B9jgvmrURxubmt0H8Eii/3FJNAKEcgMYDBOEZUR6F5TrJ4kztNbvnHPV+7sLbAcS9zRhI
74Ct8pOcl/R3/Vk1/9VfETXhQrnThA/aCsjPjKYyJtCUuQGx0qYfJPfIEGI64r0L7XeC4XUjXDw9
/hnbiX/KUT80WMkrQx7HyDoz6A/CuiNrs/r4HAjDBegvTOmGQ8rRac69yepNmNGtsHoaPxuE1lDg
LACH4DNsGqLXmyoqKceRHwEFak0YaK2VeQlPo9aBuEAKQg4wnlBMVXlLo5Mgsr0JSUTD4Uucb4+t
Yo3tlhhJBlYVVT2vlB1aEXare5lBZctat+1fXPGlLbuV2ykcGNMrcTJFC1+Qb55JqTHzNKX8Y5Nq
CFUxJj0Bma66NVvC25wZECwlQf3WC48+m3HsnznzwFgmY9u5J+SH6Sui7bw577OlgAE0YRMdQGy5
4f2jZOxyZQ5NXivg9rAiOdaUz7hYqRMXBEKH8RP6SiWCGwneF4ZaJLIL8dami7FKL7sGijww/5dY
rWEjOvkWERJpGH45Rh1jW7kzG3cBCe/MoKIjgr/oWUMc2sbzPll/CucX/krt3TUcVqif4fzx4UfW
XY9+y7AnpSSX4j8oYNF1UwlQFs2shxz0wCH2jkKbIotdigxS24r+I9rfYvdsRkxjHvTmTO1YST5+
i1H1wHMObTEe1FobVk9Xqsl8Yb4Q/E7NVKxqWBPx68vH9C7dQ/jalFFGcC68NVLMkRIxA7hrN8Fs
MfeUXl21AzhgpeDW5gVydAVRzDj+S09izHOGIygrCpJfDc/8t09Cbg1OaUSJ9k1kp9rOqKTNE83a
EA3RueJDDRubHN9SQTHJTcvmC/Xevs1Ur1D0nIRZEdKa8l8qobNyD9GKOtyowBNtu3dsUKLjLWz6
qi7HMqko1VAAJ9KiQzd7yw+OpoH65sAIzHp3+UWL8Px2UULawpxKI/Qjs1KwEMqzOWmEhv8kfY9n
RXfy6QSyaYkN4P8rVp9KAJQRu0emqPDY+9c4iYR5Lrn3cRue+O1+L958xxy7wJQxZXH55H+rB+gn
9ObcoGh2L1ZilKkwvtvHvjG87/qQ+7T2IxqRaagb5/b7O2hF65NU6AuKpTg9/XiLa6M9ny73542Y
tTZZAh6qaBuJ6j/probXtc0PIS1Deuha2k2R02yADXjddDAZ3sgTb9spMFcTx1M/FSrU5/WqpJYm
Uy0Xu0QJXdRekXZmOD9nKm1nPISDo4qj3+u9dCzUYv+5afRkOPZr8EPt11T2ISooSxa0PMsCjqJR
i1/PGVHLztwCVOMUPGi4xBRlxK40ajHDyAwlwxGNdglza5ZoUFjsgQydwtHudVxlIEYzpS3RGYho
1G2BA4uiAB5bm/Onz79U8f9HkgB+9hTtGNsnafD9m4hWkPlUWTnSShrdEj/1PmNxTVA+P7zrAJlO
mhNGuFdgv2sMzeCyZsqWW8+XdwCNBvZvyk0/MSVuhZ8qmfnUXfDzryKxUWzxMHjTkt1NjHmz7LES
58CK9VOX6LdNiKdV/8a0UVXlkDIB4Y7GAe04GWF8p87k3T0qAP+4Up0Q1IeR94LqVWsWmmRn+Etl
jrXBY0dAw5BMj0kWNmAX8O27jQSj3iPzCir8NiDEH3m5YqTBfp3+ANeowjDxvhLbXrUOn+BBPozA
tNxUWQqJFw3+7QOlJZwbyV8qjL7dwh84y1p9LjjByZz6BO5gh6CQIn3jD6/sa7hBhuHlDO58Tsuc
f5L3OvP7xiCdcjW/qFk5UMNuOovYUyESRpHJ+sTZNYpWqqm6+nU/phGhoQOfbQV9JO27yYxtjOn9
assD1RhrO2pfdpSSuvtrEj2lQQzzJBNSvl1nGHnwsuD7bpOW6hCpwrpTGfLX34UiiUPeWOIc8QQz
/ik4fosINGwog8OgDFEJ0oAu6f7Jb+1O8hHUALYzIZoGdFRvjbyK9Gm5+LDpqCR7T1dgd7+td33R
aAYFFBKNF8R7GC3Zt43oTpvOlHQpA9Gw7FWNUdkzbqL74MYvkPXZL7QwjxqpAc7wCIfQqHtpdW0T
TviYHTJhMsy9pxIf7eQRGN/BpOYP9Y2grKqLNVcOfMA89eRyETUW6doxneAQGVCL8ipsWt6pma8w
E24gYDyMwBSVjicPvEDTS9LACuMNnVfzF4HIfStUrrZwxh+SQghPTLDTmJ6HBRYXLRrlCk0z3Rbi
vk0UFKi7n7zzGcNeZ5UvtzDnIcSCg2YbpY+rF2MtYAS0qiIBXBVZOMaTPGbXdaOZFu76kPmI+mqH
sDxR/V7SAUhEaR7uHACLtpdCvkirf+2Hs9onKRScixLKJSbYzx9/ZttCPj8yB0810/np3yBkVbga
uroRasP7Te7BA2fPNpp0ppn+U2mK4p4FJWAILJcg5vS50307mfsZQYFa2a+2NY/eKJZmU1AdLLtz
gfe/cm2+3WzDh5MrTYYDvT3hkWqaKqTy7JF7TaIQ6FdIhW+0RwUy8LRQGn4jM/Wwf/DtYSAcl3xV
0Wf3IIAdoRjGUUYIsQMnWMXZfM/3D1gWEIvpKjtPMuSgB6zOlZDfTK8JHNkFkWoHkQeF2dlALekG
pW4DD3pvgQg7R59gElzLIJ2X2FhNMNpLlYR5edUR8HSgheYp4eYw+PJSJHEvKFZc5aXXUH5Z3eJw
TQVf5KjyrAkgXYRxoHpV+kEN0wT5KTx6sgkgO66+11nR089EgxR4isMoMLBawas9Wh7LBnSKl3vr
5oQON/N41hPcsETqUfKD74vHfhqoCa4j105I/yErAoTzBJ9mqx7fVtA96zmY4bGvr8sBnhFIvmU5
tdGtaoOUeAZA2s5rC+z2KHsPb+bI6mrtt9KfKn0TwoUFZCIZ77Sm0Q/7iV2nflqNhYHhFlVRq90r
FwjtzkaZr0ZCyZLqJQVUfBiRmPIDp2SiWAGepfdD2PLChrxsrsQuvaOt0GozWxQMAQXcBpXNEGDj
krVcsLKXaJhOZ11VAx/GpLDa6ZNwE2mxs5otJHbSTaGDCYCaHkahIxAtm7OIb45s+0QXj6dD9Wch
P37JjNKYyQhMGOEcSvSy4GyZcitT2qLEeFf4vSj0T9g+gM5sRJ0JPvZv3DviuDbouZGBw5NPaNE2
b9sx3MysVmAL/XZbpRMGpR70yVeCPpZdDYrlX5DMsAPmbFVTQRY+zAyCSWisaozpzJ5QxeYdYAMp
vus/JRG++dWT4mSYbIuUt+p8EzasciWlV42DXJ1iWmSAxwG5pb7imEdexkmXvDRI+9Z6RPkialuS
Haxq1cKosQoOSVJLa2hpnnz8+lCO1aqlE/0+vJcmNEKDomGO5CHz8Z0Awx3fW8VcdvANpy2xfeZ5
8VZSI0R8INkDxMNglgn+iTzqbU3p5EFOP7mJuwjxIgdEfp9atxFPpGlzU52R3PWduHxmrvnIrOk1
q8a3XMPwW9npTut26c2iEKzv7uMvZZ/EWP0qh4C40nLDkAy8GJTwDyGr4Di0uy3XmYsUQ/MTDZK/
ruvWadc0XB0bfX8aHk6xNtUtzISTGRhtd/6b+WRUugnKSO7De4hagHTMOQcsRNv4IekLJyJAvjO2
6Gp6rtW1G6KHlY9KAZYZ/srlm3O5xJW07VROJD53F9sOFj7uQRkZXVLnQhCGjxUx8xrtdzMG0tcc
a3Eo7ZRsIKWb5V2IX+MspVRiEjmmEJkpQTWhEm1xfNzIOG+D8FaeeTwDnhDxhtRDM2+mvBjvEY4G
/aW5UPB9+vq3bwg7NlgMMe4Q5QwuOpZoqZG9xiLCUEAignni08rBrjDpkfgsGFi2kNlFUxfMeudC
pIHZHs+eaq/enqWL6nrNUv74Gi1vxDisPboIV/cXeEMPX4HDPtufSFTRM/hNNIggyXnrtIhNHZH2
E3B+iiqyzBazrXgv7QDzUcjyXYy9cB8ScP+WCK6LbwvqlxQmwTQ52SYbi1OjQRhz4JN7L+dgLj41
GLjkV5GKQ52zSDQr0TGU0NRq7/gjKAvTpZzSi9StQjYPRoi1gO1tkl0mxvfdQrzbSv21bi49JCO7
lO/iTShO3RYKBTQ3Um9DbaBt78FVrw0lPjpn74bDf2wJUwKS2kwTCtT83t+aq8wkJezRonJkIMlc
9+BLRHHjS6xCmOwSx//DhOyv5PNHMgxZerz8dWipSEm1ZLzBEAUx1R/qUcj5hNz0ri7w1+Q/Tg/j
00Wo9tFA9X2T+uo2zZEyLS7/qdW+gaUn3apcFaMnr/u3K97VvpN8lP7/cn3+ajTXf29c6E44xeU/
7TMiNR0rds4T2NSXRlY+h5EBLJXjKt5lNxx1Rg4/TTBNcc4hbRO06rlRcgKQJjhxXA9F/G9lr+Nv
Of+3RqfJj0d4WC1keMl+o0nuGDqVJNHuGSWOttqV73SH01ahXxzdsd0MxPqBBjMn61tcmVnaPJ5F
dO5wXJpKcKdOeRdqAbBdREVcf2dcvn15i6GtZfxmGaPMkV4JAiqwZNti0R59sX/Fmh3bBeWPqDMe
REOr3jdWJM/AZIPMj4Xh9eLi10/rL/li1MpvGKuwec5xBsIqSjkP/krSuNe5saMkZ88VRsPwiNwB
GAilKSlLnYh7/yCovYtIjMz3P/peBPVIM9HiQOwKg8e4fROYhQwzOr/S/O7PNKya5uQTLjtlw0q8
tfg4Au9527MOI4YkR+70SUOPbitq22JmF0z8e0cc9yMiKlRAu2i00b3RLKkPBgwcztqdxuffANws
1kriYxQJDF0MML3YvKKnM2shAvY0bnZxdlXfU4HaIfxFL4MNBrJ4lkRG070R/CnZGQeTbeDjnZUr
yrjNtJ0W4xAj9GgoQU1j9FryRby3IYwcHQBuSDCXsaFGJJnBwbQxjWyQdd8WY3MHjAIBDL4bMfV0
OTSzTckldNkLxlrNt7d+NThi9zSVLs9uEgbxJdvEhnxDrACZn+NUoBucB7hZbukJSX8yjXF0ex8r
a0GLldLYXrM7h6pbNMHJXmkQpn1lEUux6zMnc8sXzRd0dMA962pn5M1cEybZCIwSFZYilQNKyJx6
eo9H7ERk+biAdIJoFvDzr2N0BKHVL6R+QNmvwoya8RDaQhKPCgaJY//3ZDuM7uZh0ROYVN6HQy8J
ieY9241k0dlhqqXvcPuIhp2Du3zounW0YuZobZ5nQfrrAbFgO3Mh7KK1wu5DfvwFzER81IayFzGi
v8IqUHI+FP5gw1an+JTAOjedBNC3jwrCQlC9soAkRcS0FGZFg19tuBS8oO6HPukF+vuvolaIMkHo
ZEqVeUqiaxkngH4XSV1TT4l+WCfNHxd6IrT3IxNPnFvsBOG6IoYYN4PkldcOJIagnphJwu6SNGST
mvLhHhFLh60OjJoUeB6mn0lhdn2VjQW40Az/PrzKrk3TxoX/w1Hsy1YKCFG6OikmVnKopKU//h+M
w1+Q6v/LwOr9SHskD+/xMMc/Tk01pN2zSLyq9mQeavbLeFtO+jWDOWr9TBTy+Q/ZYNM9dcQYmEI4
7k4emcUa6dIzcx/qNXiY9zwR2MHJqve9HUVQ1gAkXrYVUD8U5vYipBAXq6j0WAa0my3Nsc2jmAPv
pJqOd3USORsyJbHwnYXPClukQ6yHBDLWCxNREBk9ShJ6KNGcftDrFT3QXQ+Kgv3TXK4Wyh9CjUjE
oYJTsuxEd8RbIAD23SHQieflqv6WtDJPvYefakKQBaod3rhSPUxj/QeNNFpZC0qInuVX1wuGvHo/
GAdGxQYfyAApot825D95tmAH0Mjv9A6bhprOxFgVgAnKchBolAWQ4OCP3UqPiIC6nUNueISBxaOW
9fZHwVqTEiHOsPPRFK+VpQyomy8VZ8alMkJs3FpxDzeN3Kqo2zu5i8h0ylwPSAn8TuV5vUv1/XIV
7/dSgA88Jg8MgwxaVbNi29lyvCQY+bWzNhCMBUr4Hnw3m2mqFJ6LcWe8pWfkyvukTMSxySTBXjvx
+DHyX8Q8JhjEd30spGqgm2x/TpphJXK+Lhtl/h5SLYXMVgAJWIl1ZnBdIuLze4xAcscyX/+P6Lal
rE8OtHPApIbdUh4BmajVCzkPU7QtkgHx1vpZluzCLNjeno9vkaAyYZFCULiZ7Ffpm6Ftlpfjgnpn
RdNmLlgq/3sBpbX3SGeWJcS0lX3NUB18a/hfPI+i6CMadJktrV/9HbR1KWp3zetYjpjkKb7cbnmV
XCcpDyM+EYdtzN2mxf48qaZ2UFM+L3eI6FFSUrXp7Ej38rwFLtD30vyUGwjm06wXLPs2spz9FMvc
uS8bsSQqPQKS+Y1jC31aUpXtBtHkqSU9iIaI0nJ+9aodJ1S3Z7Y9MX6Ip21yGxGrFGe2q+Ve50Sv
ST4ZKb29dCkmuNY9KYNOejmsfj2hZsT6EUhEdLHe+t7qjYLKrEH+mLwcWZGIEy902fFFa9x7itm4
r4kAV6+AFHjsjN4kAQgMS7jS1Qg2u+/6TQuLNjqDct7pIuZmscZSjVXcf7CNjT1Q/vLoYamk/aWa
2kvfLcLAElVKUJpH8j1L/dovXxY9i7hSRniWoWVDX7lbhWBYRiLHzzdDZkcWBGqa1QIUYShI92vq
9MxrOqn2VbDUCw/BuI7z2cKz89uJ9Rv7JArqD5FmxYtLCbgk2RjH9aYAhGFlxd0qVJlicebZj1Dq
bFDX7vPCmthbi0XKvxj8aHJQ4C1kZaQIeZukm+WWOeIRXqA7B61oLqmJd7tv+hfbCaGVZxggzTJp
4322HntXxlpiKnz2+cW2cbRVS0KeweXDNKzGRR05BoPsBrK0oWThT0CDTM7FmMRS2BwY/EdrmUOq
GgSzRQqUCyow+0zHoT4B3G+22NDrUOkRBDtfLzWoWB1faaOE1j3ljhtt/5rIx6J98CNOaFgFqpmA
8v04B1BGvj0jzZMj/ZRP8rg+z2NzPpIiS45xZW3qtqFLfJHSpjSzs8sCt/4hFbwNYJR9bLZe1r6F
+zxFmudMp74J0b/c/d62yO53xACjf7WyYtLRXdsyHLZdoyBnV3szKhZ/NNYjJ8DjaP/hvMtjX+jq
/PkaPw+CAxQl/oUNKtfHtPKkaPiA2FClKPRGKOGGbunyesMwrmHocj9/yLkKUpDg6fRaGrK1eWSd
iUdXn60RY6O736Ihgjhp7VYJzc/6BE2w9neznQh6hVf5LLY3wSC0upZPxVZePa1D0KH34rqnN+yX
7wnXUzWIm3SKXTK6eVG3S4urmD/5Qjao/DF5x0Qy3fS48yUdlfqfRsCCoksOZzseHCyslYB3SRRj
q7eKWZibCq4ZejFTlwcLwnzY5rc91nNLgDkott6CzB8N/z4euihUCPap90OEgy3K3jFIwJKvD12w
Trw0STE2jGb5MlKDWZMbCk/jv79Sr78B1GFX/2MVEBQilzPSXKxum7JKRqfB2dHM75IYPHPIt+AA
8CR3cl2eu7eD5okd3E5jvnkGonHM79wGmPVaw/SHfknQMg8f4ahyBm/ooLFI9/Dg/VQPUkdGxx23
E5ptj0nzLD6OU8NrA7ammKUYl5NkoMTN8fSEdmU9aZFaZFeeU3/eJDfh67w5G/kRREKYHsJkF/3U
00dDxWSleG+YoBLY/QvaGkiisi0V2Gwf8FVedM1jukwYNus1oiSFto0e5i8s8YZ42m3tC5sMa/+4
b96Tk0ZYO5GuoOvAMNm7Z6symIbiNqk93ey2dtWYXq34NBP/0igOFyaV1ZqPHkLn0TejMbj4Y73j
7VnWRWgUsjQboKdzdBwY6pPqvoq1RRqQZnmt4l//mYQlfsSDJBIAB0+SPUkEAQV1na7iI8weTJsW
Ly8qxiAPIjEmII04e7vwFiC7vo7r6TGQdTFCjU+EZjaxj+5apZRroWxs5vn9FJv0FGRfIFa855Dq
iL4HrlfQ5osX+FrnnGVGBInREs5a8vbb2S3KllSsKdDFn1wLLYtIzRmy9KzXvsWZ8rJJad90bAHQ
w32dUOM0qU1I+n+5hHlFpFYApArffJ6pzI5SXgxh4EGXUoTPT2lBY7Co1jCX+aZCJMS1j+Yy8LL1
pYINiusZcleqGw9T494hgap/EakISXH38DS2z0WpYyI1zgYd6+v7RUi8OWhpZCYHXAih2oUGYp4p
oOcCbYM6UpSonqYq2ZzyuJaWM/60ol2+oRjSt/b2rE8jSu/xv9WPi6MV91FKsJv7ii1BjT1B6I95
6mCp6UycRPOGVpdS18ZEy+ZBs9MziVMND08nsT1B+vc30Le1uCHa0xl8kBzgTZUnJxGJALsGtJmc
UGFY/SLSuZpn3Yxfy2WSfpW7dvnW8r/8bXWgg/yOZEL2vv0GGx89mTq6qOH+ZAAhqamBq7VCe3uy
ddhqv/F+6c6gTqVOa3YBzIoJz4ZFjyb/WSoV8hr0C/J8qLTJNPACgMY1KNqI5kN9MtO9loS26uL2
PqLEjahgLH046HG8hY2VZbTjS/EO4tr1piGs9G9qwMuyjmnIaziMm+ANApNEkjvg77f88GfgkDSC
q0ct7e19dQUfT5B/2xcFp9ETFeq4TnIBANkJWx4mq7kPvx6uLevNY6d+9tqS1HxIYdtz5cU76+m8
Dq3Wk4DofI82QjItgqRzxRxZr8/f3gIXTAwojMi03Lon6j3GENhxhNCoLIbdfGOIS+Qu+RADX+jG
OdAuyey4Ssv4a0P/C9vslC6mnL/6DRkt8fKxyVNS9nshEPpLzq2qEVeC2k/PB3WSUduzn+yIpJp1
Xuh/W9yPvYQL8G6T8Y4jPbeROFXETx/YhEyzaNKbnfn/EK4q66zdJgGCMl0tf0l1fBx/FIEl8ZQe
gcyXPSEHxbyHsFGS5TG/dkwtPJUyjOpqFCaujIHa3Awkcrs6251EJtlzETkoT0Rh9l/kJno6qw08
IRfzPmlv9dqdvFXxBMquThU7ez+MPdIKtgRb2i0N1CRzMgCL9LSkeeq9rMlmrol4Te7WFmLAmGY+
K8AcN6YxujYw/UqtKNfyqwcP1BY4Xhsq1tidoJW5f4zwo2A9kWIcNJC5HiiIz1Bfs+P8iDOlwzl9
wUukpwHI4RNqRm0NW5BCArP5yH3M05frI5MtWcqysBPWOmNe4RIC6vHtVQ6E7w/666P3OHVNjGjG
BBvtL5apOyXaU4KukL41XyGgaC+FPL1UBSctSF1SVHTLME79SvwEb0sBJfnAyfHuJ7RqlDFtC8o/
nWz/wrTEbedqLoc9T2YYhGqVtHETPBg6ZNryb5Wdv3qvcdfAdGcB4otvSBUYl09YQPA0+X0/E7ps
deYX0sZdEwRAJtGpO66CCsAxle2Doh2xPLylkgeU7lwAqvwOmCvDzoUGeSdCo1WN5zhs8fv7RZjy
36JnT6lAHxxB3M/1ekTlRIxIS1kHFmOliE0zLQ3vIDU0xcE7qpsBaEU1xxqJjRAvhxPFxP92P6xE
sKM/dipa0MbjwGC/P2HNV4wjkjhb/1052MV26wkWbQ68lWcCPl7AqjGZ+qUikJq6VNTF++gRHD1Y
4Rzf/uU01biqT3i5dB/luYXAWtKepDfn8BYR99NXRIE/WaeWYb3vVih6BGKf3tBLw4Xumola2oKI
rsX7nvjOvoKWK7px19JrcNlOJ/mwI51lNFEvmtgz9kwa6z/ww9NFkgrFH2sGUUqoW69oVBylZNll
+/jAwJCXdJjtltIgQ2EAwo//ofsk+jU1cNkM+qvBRYoGtHVHjh/Po5f5tzMv7/m9E7ORGY+tAHe3
z5wD0I4QDfWUjVNZayCejAKIYpN04sjk9db7ZO+7pSdDJeHItZ66FCjiDYu0KcsW4LWHVDXsQcDY
lPiXoHu/3EFKOXcAwQ92UDChoDYp6WgZGDDbwCxwIrDDw8x3Wt0WP3tPnPmKh14As4nxJbJdFCO0
aAU5wBsVNo5T9JKMkIjdWTmmq4nbfQqJ/MKwMAuLG19ZC2dVcKJVz7FDZUXojguffSUCY/ddnWCx
ZaEDRF+2rJqxfYg7YZvieA/ljWXO/Orw8llt5HBGmaZ7GK36LPRcpO0Dq4vYykY+wXP6RwhT/jUF
2RnfbBsz/+32bDyyq4RHBI0h/6uJ2bN8+t+wcEiGLtoTCAXF0QlKsWPcKh905Lz6Mpjp5pwfbY4l
gUqAIaYCVLXhk2AP2LTV5ZQ0emEmAMF9SHMu5BBKa3BEvqPWSqUSrCW21YDikA80gomTKnHjTzTK
Bk/L9QrGBCSV9ltWGFK56j/BAPIVUFqjry/43lc2jwBtAFnrgEUqDBwNQ7SDyJx6IA9JJQ80aBXM
l7eXpi0RH78c35BrQkXWWqi82m7h8msC6GK1H9teHU9L4L3BC78x4Hg7mGkLDoPenAy6SJ9GH/jv
cOX5ka16+EBYTprF++t0Bc79O/TQTlnLkBF4Dyv0Zg0aMbroBGIklwtCaGqz+Vm4yfL8WR5LT7yo
b6Cc/I5mDQojOIL+ih2RQOcwzcSK19bX3HiCZR4ne8xYiAXjTlCPY2lPBAKcNl2HEX9QRDX1UMOm
I0BUWZRV+xVaoMOzHLtvSFA+VgZLB2FApDtRxS1aqnDbHstm52dYwav/fSRcgMQIo9xLUbmuw0Yy
AJfq8cUMfOEXSpdgRlDMLaPNVRDqbuUqiYcozXFjZLOfPvCg/mWge2stQsBoN0i65PZ18MFlpp8k
wg2nTOfcyi2VL/5fWU0f2KwatN98MWgHJvZ9SbDEQc5OXerwmXbme5rWZUxuZtqYSp6hLCac15ey
u7N9PUEACUOHsoorqeDsXcPJQwme6FvE66cmTZfeyhIB/Ha+V+WPU2SI3tbUuSMQOJNPzs6rinvS
depHY2a/P6Q9EHzg0gPzCUGOp5+cKuDCJbTD7xDj+/yEktuMayZS2tAfDtx8SJxcln34XARDujSL
J7aqqFB9Ecjire+Z+ljjzKj6vutaAHtFBPOcFVvRZNpd5p3bYb+iz+beXGcnQjl7EMFMGBXYHZUh
uEsYjppKxt1fANswO5dGD6CmFdyndw96/gOeXv9d5c8wLC/3YR+G5dd9R0RcNSXIg7iwSEheta8P
FfGz0pAs2osRRah5br4z3UAFs0VIYX7/z7E+dQsOftB3zBr3cnKFNNr+TSEZym9v23sGJteq9sEs
MLtmIutiNMOH9o2k0d65KsSw1v7e31Ip+3e2SBwGsCvwxV9qr4Qr2XKI1BOJxQaQXjvX95Uieg2F
diXLK4g9JypEKTkZukermXP4Wh0mdrMwUo9yo0TaBbyqrLTNtkG+Jy+mlbnEggRji0hH+uNOcrR+
YLa1++MHJb0EkP1sEwwQ5A06wv6Y1NB7uQFCVblcYEjHNB6AcelSLVkavutBZiasiZSuDbZe47SY
In/Tc9kw6gYpTbKcRbsOzVk1ye82M55UVKqdGG2gPfMjXTF14mepbTEKcP4CdbusNWosehK/9Svq
UjB7BR4O9XvxdvR7JGXEUzhvXbF7SIN6XvCq1PljZn8BVowzlkindjsxX5FjReTIKS7UqfH6kVBR
7GmVnRkgxZWvVQQm/oT1E8vm+az/nL/PKpFxsDIXT4Sr0PAzTfDowC+6zD/wEr+Tk0CbpVLLlYGu
qNjbTVYcR9aZm6NV8VXzOnHPk7OHsRAi4jDEUyHY9Wc2hv7IieIjfFCbKWrhK4Oagwtc3/V3oRx4
yxQUEF46wR4s7lYreu5J9QO5kt4Yk6SNfzhsKHT/qQdM4AeL8mZIvC1YVT6iSB0+RiKMzrMTlNrl
quwlmFt/Y2d84vtYpxMhCDoxK0t0W9ikHzv6GkTBCqPiLXdLrtOjXCXFkGL6FaLRlR2yS/m8DPh3
izW54BSkdbd37cJNP0eW67BOD/ccQzVYrQ9gM965YcxonyLcnLhmVcsvB6WOBTRjvw08Xz19Ypto
5cwVLKDF3L3RI+1tOJDk3LsRR8BWdhgJ9DIlHlKSHCjwfp3BYnZvK/F9Bj/n5jPDBVMXxMJ+RXO8
rU5/W91cxGWB8x8CLYK/JitFZyl48l/0ONmWEwGWDUCGSQIaZWzM3XfWg9Naz3HIyhVd5xB8cqLF
3XYShrEZCKu7renfBZY+hypRMXOlEnawKrMj0rzzQupjB3zbM1JScjdsCZvAX48VemanklyukKPF
2zwqze0omGiIbEfXAyRWNQorUp1Y8op1f96E8GDyaOb18s/+RrhYnP/amwL2VgAJOXAKXP/HDHN4
bLGOf9/fKqyfubw1w7cgcjpjEkgfGD93YEHTJU0J055L9zow+EHr2GgaRHKwkkh+DO0BmzjaSJcv
uv4OuQZAxKM4GczqNK3klWLxFb0iandd2m1ueS/5bfZFTlfCwk1vfUKoy4v/iE7xtAcMM7jir44B
zSA1MfRCPwWEhLP8LKuu6cJnPBkQ8Si0HmQbE2ZeScyLMMdTIhHZqgzMV+Owgh8ebxLIZb/Kf2Nq
1vWCLau+yeQs/Pnmtd6ND8j8qtDDS+WcEY0pTFH2We1UzYCdLP/tXjxkJHD34ZfX/zLHvck3F0uv
cw2E/irlQTBXgEAM9q2iLVBLE1XE7ggyeozYtLFMzvFDseOlnASxSfDtZo0++BijS9mZnK47Guas
5SZNQ4+nMjIVhb5Q9oC9va1pXB07TABcUl8jPz7kdJMCwlkXF+/4rxRo+2dVFupMW3lfrvsvrHRE
uX82fPBSa+LCYfVPoiZmQ7uIlMxcm+vecDIZD5Pea0ass2qJ6bUeZ2AOjamP9y9YBp9uoPMCN6WD
epQk6uOKILTw3nVBOVvdL1eVJZwq3RAmBeBePjEK30jfVzKSWid18RKsxSdM2UtnxOU5NMbgy9qQ
18LefWHMAodZnpMWbzoEbIF9P1665N67JGHNx21Le/cMiSxJkLLxTOCICBBqZKeysoVnK5GY3g8d
Jm4DnHdUa8eY7WGBqMZPKhg+fOZmM49Jx+yR3YtkPLbzWCAvFP4WYz4iZ4fg6q/v2xCugiB2h2QR
JHQzZUx2TDmCaU4yVXfeECT04lFATl9PJ6KTCRZdZ5I4R6iZIzKZXRfzrCP/7nZ2q+jRkZpH46Fi
JPhn91SXqUUpLVxMk4XBk783+n6yRJfoHQHN6GW/SS7CvThCO2x6qRacFgUtKwnQY+gQtUktbmx7
UFL9pF01HT0xuR/T1+4yw1sVQ3PNHuOCDC3zpANV1TMHo0HHvc9gpYYZKZjtmgpe5J3TPo0xNc2Q
0psWXkxkRp7t1IXTlDl/mhYH7u1cfaKIUNhL5pujeokilsl7flhGmCcGcn2SxI5cP2s8WtRzLwiV
S49ilgM4Ntu0JGgKNiutEoF9B46DHhqw2qUGoVRLPA/oacVWtdhemejhHZv01VbGB8Jgfnjj+BXi
a5R72NEODl811G1KLMn/Mfsgk3iBGuK3Tl0oxn9gI2NzuhOXcmx1wyofh9gCEOTwvdJBJPbjvu7g
lar6Eczbw30qP8raqrABGHqwOvMxvp7hNhOyvytqn2fHp95JhPs0hHcuKJAjQ5Z5HPptGNkAaz60
vPOOoC39PIaVH9qPX4ExS+1nAja3ZcZYI9I6Vt6TezjZqp9y5CsShncfKFPnfzKraG45/xEin+DT
5bSavbuy0kBFpe5jsz51CyVcUC52MvGUruzidn2bTzncxpmNP+jKsqLHrhA6+EWfXJ6jd6BCmw+T
oaeD3VODW3zTMASIvn5F8ixrMfcdxZmkKq1wv8pvNNZOfNOOwiGZ+preaH9CrHJcwBI5RVSfnMcV
XrxYOAa/dxyx+eeVSk8eS3zEv+MQ11k2ghQk3Kc3o6Edsa4QtRGorRzQWMASfqQqPnSDX3FsrsNw
1m0qSyRfkcaQvERmn9gkwyiUgbzv7PuYYggo1yv9n3jNRSVEI2xq0b7MXnir7T12OGXV5hIoNYcN
3BSJGPTCRrt/yRiXyqX7So8nppAG40VfZuOiykmEj5fgc3OKV54dD0H0dgfWaq43LbOgr2TYyDCG
9eDG8QfcoSJOWORvReEfq9KdkgGWSEzAKLKKnvMdVxX6vFLAEnpnnOOC2IvqOg1kMFZIKVV7Vpiz
L7GLSdoMlseaAPjH3dmGWhNH3ULTOB9fVRIQNmwQSLJIHINCZWucmCPQoKQ4HJ97R8XxHpzrWf8B
PGWi5jZtNn6USQJuhmkPUKTe2Vg1SUDM04dMODH9TUy3w43VPD6jJ/yVSFGDEA2LQ8b+qhcCfUE9
+GSCzz3H0o4r7kCRdNqxs0LhkiApxZSpxqqgyZmH45GoZuAILXumGliOPpp43gQX0j6sUHfQOTFP
huQMiAsdMfJcC1QAIcjC687MlyZ5nFPDat+TX6GXwbzFoLkbB9pPnuF5ykCnQyfGFpGaMbknFq87
DJPXkrzShAoMDDkIddgpLIcuWXvsJK9kG9nGnL4oGe831WaraOoLkTXtnZRVjTE0oHrdBrWrrjeh
GRiB2cYUxlgP9ciAW3MC0lVc1sahL0YgHRnyvjAkPa/OhS+Gs4pNVA2tnEQxWZ6nR9aqn/TKZwXi
3DDRYay68c97Sxq6riiWOL3v12HY/kvxJGAewmSGjxnifr9n8Hp6gUsC8Hzllp0dBmFCGcG12nD0
GOqH0MrvM0+1G7uEzwg4uyOp/Cbi8trjBDR6y4vrNPhXLOO/JFnaeYIcMju4POL1Cnv7nLex5PSG
lRmSDkIqjMM8UzJ//24sOtsIHZKrnvUHti3HY6bz+c/efGcbLw0pB2jkZYERES7MLqB+gUpEabw5
6VTC6oLlRDNePsSAR1cgGNNkyvMjuoVu2fOCePwuS5b0dM7oGTW9Wuh3tn1eLC0CGBZ8lUUgsnTe
rh7oJVWwLJtPPw7VOO5ho96AxGRLAlkKhwvKKuZqemtmP07RqoaVVFMLJ9d/MZfgkDcg9opQprME
gsI58oECrrTc0+LrzC55axNwjRmNmqqHXGcglzgmYh8JiTkhOHcucNUWDDL6kKmDov5zfe+WJfCb
TkcoYiCdUazR2XAK2J7b7VIWs6vFHW9GK07jO+t8U7F2Zx/PXEHUcu0SHrz8H/ehyG2oJnqGziGl
tV7p6JDCVTRh44OwLBnQYwKXESJ1FwU7+QcR/VlkBwp7AXenJjS8KzxebqoZUbzogf/ozlbzK6Vb
CtVQdD1HtHoS1ex30b/ygT88XmXk+dJvPG7PkRdjF1V+JNXF4/rZhkXG7CWb1mJ+/PWKN4ApjNI4
qwbYh+IKohfb9QQ/1gf6w9y1jl4izWpRfeNWfkAPTcsZo8rAGAUjbHXubrwE69h49vOyzg2T1Wq2
mU+iAtc8Otj9vS1hfAzsKzCdFDLP4FamTY0RRwXcYcQRLU1O9jX9J8uMJahBFhvd3DnfnIGxDk7K
dJo22joJ/6lS7MA3yk6ZGxJrFIDIKwMKXTXcJEnAnQKUZt9212ImG+uZ4ehXLzHaWykEivj4keXC
IxW3GKWacTqdbv8xxntA3C6IHfeUpsotVQfCkham10gBMP8ah8aaPD+hxm0GC+KQ4r2GWVJIes/D
qqmfDjajlVDRDftl6KZc0ENhuGhpntrMHacs/HtSNRkOInuKcpXIdYW7ISjM0J+/jWPp6eWHGVLR
km5G3IZjKnglRzs9SSJ2+IXX87axNf4fwSOg3muesDGBrC8kXimM33nNHwVY8xI5Q8r+1QFii8lZ
0QCsL7j5vuSQkS3JzG3ymWRNoUL2Ge4DbU+uclAgcJQXTcnLpSXoBD5IDJrfYaP2ilqEaPvGURd0
VBktChFv6hKFIbfy9ROGsYCh9AsNmF8kPncQLHvgBY3I/Lmkyy+9SC2uDIafwasVPc9UvqJff9JN
HkjPiCUmkf1fF46h/imPUPExxNjCxsjfr46647TEHlwuCxp3aiejSSOyHdbeVfLx7Z1Rmb48Ooz3
EPnSZCM4vuxTk0LTVsuJSFUSZUSxISMmtWG3qONg/qokN0mUDS3urGnDMuOxzFe8ETePgNRESL71
ikZV+syBQ9OVb2Kps6At+hcwLbV/GZRhwPqlGAFlgMon6t1OFPIYk05jhLUy+JwZAj36n7uOxXwA
yEdZ2yavTncRowcK6DvbkP9d6SoOtpJxeEsKtHZ5ajf0X9tGfcxUDetMmK+/kBr9YXe/bUYkDtvF
1B1h/HmaSOcMZbrzMYxgmhKDeclRMf1mMjJjylZyw0GPlMyeSoxMfnBU3I4a+zQsVymSnoUF92U5
uZsVSDtk+ng2pjBhP2XGI9qYbdW84uN/V/hP/aouslQ1i0P9FOcLWHlo6TrU+3enmYl3wivGVAXO
cFGih5AkotBuewKZG9lSVpNjx6AentoKWrL60TuZkPtxuBGejlgJBgT2L4Ja4iUOrbhF5+J9Pl0c
jI8+Yc2EGGFRpHTnWVSpYe29wpW3vfF0ERIPMUmnxVZumPFkJ1R0Syp1bM7/MCZwmeDxcWTbLexq
iL0rf0gI+nYuQVPvgtdUFbyyK1pUOnQGHZ7et4hCpQyHgm/koK3Xy3h6IclsLifTKDU6Uc95dcoJ
RFAZ5Cj0TnzFe6XYWSg2AUDObF3LzcsNyZe9g3wEV4gmrzhIO+i1YySM6Db2NlLmwxMDCC32n1nX
C/rZ6vStDgN+p5KccyYD0d/VS1zpHFuGfHFkY6yWxyEXPr4q4sX118iMRu2f2LRl8mhJN7qmCoEy
LaRKHvsmZpQayCQ77AnwZmWG/CdvF19R5HH0oYFM+D4bGacTNq5jkWRPVRfIC0W+Rg2BfgfNrZ1R
e3FzpQfutQkKevMHkKXzPA8928sbkX+bMEfujq2Z2560n2YtWkjFevpv7v2hkF3+emVfYpczTcE/
r4rSqTLwVHnGzeQNmAylAy02Y5OuKm0vVZLYeRInywM7lDGNppYAQk4T2OWRr6MKM2ye2UaZAVVD
Al8kvhLE/PMKgd1M/A3GQ464vLsla0bGMR/dtUzUXOcMcJXkXN+Sgk52g2xuRPtPrK/msWGpUDsG
QSexNizqeTTz+BDILSWJA29Ha12RV8Voi8pcPHPhxosQAK/ZTAV+gnmy7aqOQ3XVBDV5W77R7ivy
U/IRbo9c/wEV+3e3IESVXrTcMlUhSBkPmkpONabHe51oyv/C/lcORnB24BWAS8izUVlEa7tfoDRR
hGXd81Q5u0z+4XAFYG6a5mC3GG4+at7Bc3CGfGWvwnr+xVOALW3atC7MZflbuHhMBU78DhCt+oyj
Pnl2JZSECzA0Fc3ScIiaGzb/gM+wHFPd7Xh47A/Km1/ChPKSTMrSVCVE87UAw0ZAKC5EP7S4HPSD
0gCpej0RvjwKb+ExQc5yzZ4zMFufI3Q7UN6eCOIZe47I/Uufr09zK0e5kqoz81ZSMrPG/QbFzRNc
Fu6Z3pNAMqXtlrXCGWmAAE+io+nwBNwHcR7bnoZUWCtFSo2s8C3op/jgxZs99360AcKqyv7B02Pm
yisoszhAXfv0FghWGWpYFFRAJFF+MCfOCeiXxj3jRd15Obggo+jhYYh+2rgCMij+my6lbLuMLE3N
CyfPb5cAU0mJwkvKZ/Bi48wSShrar3GRWM/aIlFkzOtrCsLpbK8SBnAqXFNOQ791BnBlNhrRO9s0
2KT5gsUeHXKjJu4dBqSlXQvbZh+A81OHFInPOy5sPQfl4VentBWeOwjan1OFIM2icmfuUr+f/vDy
+2Ws4mMZshx4ZtGoegTLfK4Cmpg24IDpwRZiQLrlAXSwncrcuube932Rf/l5GrUaNGtfXfGYx92p
m3hnQBM33aLmALc3xNyiEiHqBnA+jtz6kWPlnJSfo5vFv4CCM746neUU0IgSjCHuUmPCHMnJpnKu
jcviGGDenSk1EEN4nafIpx8WFQgtCezHnIsKzgZb+pwQJeuVARQoeoCKbPoOecpFKdJE9vguuEGt
7AoJY8QGHKCTZV711QGPRd9LRTijSRU49FRVs5r/9K6owxr5NIHalE6enEblVyDJmnl+NN4STTfd
vcAVFa7ZN2+ZfxHB0MmqyX0KHg5FOSAlSIxioKik+sexd2LQOpaaZWdufpiunRaQ4gwoq+hIVpyl
ThR+avVImgbTtiEsaeqCm4u9Hkrat97d/OxbGzHEckICZSJsXWMaHxGjP8wgPaziKe2nCRSSqY3B
yfFPz4BmTjjBXPz7EsTv8vPm5/+Btt4GUFifcjo7cDWvtqVNH7nHMg/6ajb+xAco4T4cXrh1DpUC
PnxpBMcCzM2xnQUxKbLQMmPVhEe10VMJIEa/MKitZQUE59xvsJONdLPzZK8Dx7qndxasUSgWdD+6
mk0MbIlvC9M1LWGvSn8KbSxwGbSKXd/bOcMsUitdDcdmRF71dCX3vCiiv/McNhelMrtFPuO7W+Uz
LbYQnIfaWPqgKRjSstO89kvDER/nk5Evk0IOlFi6Hx0VvdkyEFUJl3TDLMahiKSXu9QmfL9AhgoM
jfocanMCDX7behT7YstRBHCsFZ8T6ob1dvqldR0W2aveaK4dFuKg0XXuD9utLTQojb78n6cAz9rw
Y2LDQv/DZEWp5z5Z9ch87FESimWw1LkksW8BQfGeNxl/rSqckSeg1qTCl+g59aWWHfc1Ed16WkJM
cuvWYK/SVs4XfSPDlf2saNhHynOqYdYrhR1WoT1sZE4kkpfUNDkI6lhLbl+o7CoLT/0y9XtefDjv
X3r6kdCKMsSLScrp71QnpmAD8ToXiL4n4SQEp1CpOtVc/R6sx5CTfxGZRhBf9XibKmbIKTkowHuy
LuNQS1D/ZQe9xctuKFSd8OGVQzLdPVerke2m2/E6ep4kXr/w//C/7VYIuUXHO8FSrMlMf4bCpxJp
XVSdZltfJ8m/F98gCw5Ghrf0RaWAQjnv8N1AJQ40ZOEftJfMjw8Mp4JiWSyInjjuYtW7I03WtnKJ
YYWCjOk6pwhTi/d70JTHSEFHBsV9CvCEbvz45K+TdxX6+aISkvJCnHFtIawZ0mcL0zz33rgDUYeH
I8vIM1XA+lDqGEa8KWxscHtVHn7iTvx0aC+h68RfzJbizsLK10zC+LESsX/pvI2CkF9875BGF1Ah
dAuGhpP8sRdxEYvOsZ3PQb7QycUn/EsNHFt4khlVyquTRNpjWq3JC7sUOtc53anTqlx0vHF9omHj
T9hfb6IPuWq14Hd3BbwdoZ+luZhiFxO13gKCD/2qbtReh03RAo4i2V+oU0ByRmyGgm+JnhvtqGYk
VppUpF4miOpikPHfWZRs6Mo7gq/GAxPUjUsIRsgwbrnQqgNnbT38Dj0RYURYI59SYX1Iz+9J4KVM
3WCJ+9sA/BE9zc9J+lnfuXej9JPkw6c9UpX0W7RqCW/cawFcNwtU7F7eCUxoud8t5ooGBHkVj5Aj
/+SG2PNcYNZOyyslcMkUot+Dak0B+iMMGMKTKY69zkQgSPFPZZpZ/sIy+T+USyUggXVzHi8K0pgC
+ByZqTbWsBYo8Iy/KwvytRuAjTLJPC/8Usp1R0YQHC+qfmFDAZ37MSw6jGU7JU8e1aJm/KnhIdo1
pqtPObFxQXMEansgIqdtFrSJn2M2+4Kqf9zD3NxfBR4UId0E5iVkMKl25YJOJsw3mKPjsIU04iOq
tXswuVK7xcr83AZuOCLbkmUIYg7I2pqWUeAP5Q3SOy7M8KsnY06uhknQYXyfEfUEkXF9dIX2c7V3
GPjxqvQ71PqFvmDhcgdjyyhDj4djil3pYoI1wec2WzlrV2EQuWJ+BHCpW8LQwU4/I1C0k/SH4wn1
vkoz95+EN4nI1hSr205UW5oxT54uY9RWPKd3ovUSvsHUNXfuwe3IErawk8eiBaeunQibSlcPFXuK
Vz16vdQ/Y81p142xlGm+KYipwJH49MEccPMn5iIT1JuL8v7Cfkmya2nW3lYPGhLn6rd/IpNgojKY
O3yRj9y/efSMWdkyR2FuGOU3r012XM2SdeC81jA+BNLPXM+ToK5sVJl2fhgs8/CFtTi4Do28roM1
5+B1eXFok2QJL6tyEozdiYgVcg+Fh2RlGCM1+EL54R9DadvuCLu9DlZ9grztfMG4DcSRDmSqF6t1
vmJnDy5LPaXEVciwXLiM238dsm5L06RSxqFKugk3a2GpL6lgcmbV/66iTaxfBtGyVNMhgxm84qzv
yqeGzsdkgdyBjuATwtirw9gr5RgfcthwnTXwBg1V88CM4VWpdfPoKM3/RX3p9SgB7BUJnADO1nPa
mMMQ5Rk30SVk7DtiKW533o5hMHJJkVNMtZM2eUvmM+TQGvB49DPteF17aT5OPRh7nif36XjM/bLE
yT/M5Op2OZwdZ+2QQp5k1302BRyp6ZxcK2ylEiIvfEzsZ/qDlwfEirPAef74KaorIHOTjJr1BPWa
nWY0QaTa5yGEj2siwG+AROWXI8h/F2Cf5zN0cRq/6iJRmdyHqLWyVO53+Hm9nQp2QWzTLO09SQRa
fLh4W3QbqNnBx5fklARyFINW9OSZRbqSb7G0akquuFgFDz7kIgRYFP1yrd9owWIhE7S4LqLusVT4
8vjfUhc4B4H0j3JYdLoGfyxUxIaZFQ3E24XbX2Y38JlTe0xPP+uAVpVGPlu98ZNzeAS7F17v1G9V
uqnBv3l7oFWkdBimtvk66LPv+qfa1s/L6QDPEWVHI/F92mfExhrxMiStm4fpEqo+YaPFtL4a225k
/88lB98blm6YDjlapoSH+SFwFLTQmNPq/3rUCE0CX2Snbuaeun4+PqWnPddT32ZUhN6nFPJkblx+
7rilrarucF1TBhRFRMLZRrkxrdrKM+MHLQEIX+WhPQt83iW9epINCgdiUWTzvQuQKgM9PLVuHodL
DIvpWUz3FxibHDJD8/pVBmzRo6hwnsTObJ4zwUiMhIzzQXvZMDX2B2m+3LEIKH9B9OueGsw/SIqx
ZX2qirFwcONorIt+bJ0kJrhwHSoUiw2WSjSuAHnd+s13IZLuXbQ/IXuB8wyNpLGOkLbmITySO9Aw
sVpobelWqXqUAdA+S79YDAiE4WOmG/oQgYcEC8PotsCD52VkWc5evjWAG8wbJehLg+Dl3T6Lqfa5
3vnNL/CiLZmI5pSL3qKva7Zcpvf16e6pDug8MucbG5Bcx7RGctzE/LCa3Jrb07iA7cYNXaw5r0h/
VBwNnL3YqmiRiO9svqFusTpJZToylLIW1UrYyyGXm9tmOFcwR40hiPgZOzgl8GK9Gj4N/UFZC8Kl
14iNNn36sRG8mI/w0N9q5ZIFfMezg0XjTKxQU6gYCTJgE0UWKsWlOrbtmNdl9sbtsy56Z4V3eB76
+1DcNuz2AAqB5fE6bZtHGGqAQc81aRJiFWDFddZIykwX/wHRAes9vV+lj/zfTqtkPokrzqoUftj8
5EgCXiCjfMJCP9XWEajXsBU3+3YrlgdHa4b6kxdA0WAs+6Sk0N11Ba9l6u+Ic+KGHu0Q+hHV23Xw
vtD+KnRfzUNPHiqzSIdpbhJBWJuM3Iv9QsqfuTGLtIGORpoEBGW8TiEQ3d2WjPhCvpyvPz/1dYdQ
/UOvDfpxFf094ojLiaHmSphYIhxZ1xSwNkblm6TFtgG4dcNGM8CdSKRTV4zC/KINBB4oSkZb8KlK
RPU2h0kqng8d6RRqHoYgwrJpv/2dyijkL27IWsDb5xg1To4iokTdJygL8n15Jpy55yVWwGK6c481
nyx5Qa3JU4ZxQbGuEd8g6sN85AqwU3gUBUl5iOFEI/S+2rvJq37EQJ5xOOzdlZsaS8tk/hq4aLHG
1GXZbD54OzDcqj7WblcK5gpBsiH0q081m54fIAsIOm8hJk4F0XUWt9SzBfuuqnO3IaLcLsGyjnrJ
/g1r6RSUcWeTZ5ubFnPEr/65dnej0PawHSBHOrHe0raHc8JwU9GDakr+pNBaqO7cUBLGOdezg+Ek
rNu5fWHUE7nb4CkUwLf6oEhZaJXlt19hTNsAGsKcxQ65fLL7rH3s7bHCY2QnN6ZukaRs55XkWQl4
UVJbRVoCHEn0x881SbAJYo4HWWUCVhKInmeY/pavov2ol+/BLLQ5WqkXo4y6842CNoyNd31LsHb5
APwK76DwFVOq64LqJEDBwLroC2Wn6BtGI1BXztHw0VlzbZUz/xz57H4Ftq+wsKEnIDY402cFfJHj
aZzHEYG0X2BI4wYp1CW/fSEh8g5Mc+ZtB9qh14vDGIdcNRAiClgLzyivKUn3yn1tJ5smltW4XPYF
AlwVIUm5wxYnl5jkPVPsYYJnveCeHhFn9W1mQgfXWHKMdYYSMuVtwC01Cfb40K7BB4J1TDLR1HtA
YRG2YTmowXwBnHV2bUbgQ6TnyTezzLJCRRV+Z4BBKV4/pzRkjVQgeWDjjT/C3DEaDg5B773ZqtJq
7XbEmtYcw3+KH4AKHW5MJ88KymZXU9rJ7S1HZUh0WU5Iy+91epKhPRtqqNVdvogAKYEZj2FzxsiJ
JTjoE1+TzTZGIvrxYr02KC7AT8SrAg+gEEn4QZv52SA36k2O7vNQWAHZS7L5Pgzr9BmtgTZo/mND
Ulowepm41ASfSSPtpZv0TSqAiUhmEkLnAGsacZa4vSH9bYvHJH1epp17U8lxnLek11VF/xRrHTsR
G6wEi8/MxtJm2oeFLtO22Mjk9Of/Tv4umteNTqYclG6P4zNZu+d+HXMX8OvHvHaikVW3i51XVIsG
J9xhGuOiaUQOJRT4T4diWdcQV3JG51cFxpAXhVKzBNZktUgfmVKtCc2Nj4nPw1+M08ZfJho3W5sZ
bX6GbL/LBazgAamLZAcQgJi3hB+oSnas+biqJ/6RSx8wrA40To8yL74Ihy/x5rgP3gp/CwW3fwYQ
KcrMPCJHe8hAuTd19zb6eIh/U3IMLHm3ecBmJu5ipHfKzMEUgSsuh7fP1TAaAYNMV7IltvNpBH8e
8SO32/F0XMHV3SViZ+5X9kyDhUecpMKINwH4y2XJIJ7UzqkkOZehWCn+Hw7gL7k2KcISD1Fr0Zg7
WHmL/hewsqIG/7RwthFpbgbCoVBw0iiK4zuT0ig3AOtQKlgPSCSbrYKQUefpfOGtSV3UYWC6BpT3
/GMrXDgKlPzVjm8rBMNDCg4vfdimrTKN4rjKDkmG/k3PaAJLsY/5plBduAuUSsLRSfEV6cJJUD2H
wM4iuSsfdn6creal4EaWG+sEzRGY115arToRnHdnyoGxHEiYm4QTvwH1oy82Vzqam2niy/3d8TMt
MDUFhyl3QHKjP73qG0Bw/ToKcdH1EmNQLeNHhqvVz0xozpfpT640tL8cpio3iexm9CNQABqUZ7z3
Ai9A6I7EpsY67RoNgsfLWIiU/pFUhXkHBVsGH+TP1Suqc68RqrJ5AvWSG6DO/uPWiYCxw+Hvhqom
mxaBLjntd/to44tg2JBYvhs4B9rqA55qpR39Mb3UcOUfOdwqUfw1Hyc3QqNrrBetMoK2F5D6tYRO
rdYtFiPP6nZc/sNKBMvEsRi//O359sm3hjEhG0yrCFBw8y8AGlbnNgEmNumFO/3ZjSvHHEuZ8bWg
loy4+spBJ9sZI46zpiMdrLjeCJQhhTZMpcxHI8E8AmAaEd+C78uzp+sQXiyEZ08wPbtiAWFQg1kx
C16tpCx43OnibhpzdU7Voh49JQ3v4jwtagcuwlT0c+hC/GUVw2jkUWJ6TTQ4r9LXbtQ4Hm0TJeeL
NoTxLH3lOTD3yvnCYcxZKp8jqUALjYN1eYxpTF7UGLAAwoLSyZGuzxsgtc3L/AYpMzBspqvrvKqB
uSEwo8/5rk5o5G2j0HJdhsanmTJ364Mg9UzzqneAsvIohqhy8jyxSHBlDNzVkBWqhn6UpgD4vZgL
Zb+YWWY6SXj86PVUR5EHjVyE0zMUN9ZLW5/ZrOrnJhbjsVnC4tiqJvuOwvwGMrSGmR7YfNH72jZs
ds44UgVYygdIihWta4a7G7t6qSmC3bUUzF1aU7d0oeQ=
`protect end_protected
