XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��L~�D�vHw�rY�6~��)�ȸ��1�Y?�t�$�y�?�����=�Y�����l3ğ�Zv὆I����nശ�O�B���/�j��=����2��f\/�ܚ[�_�{��s��*�c�G���V�WH��Pv� ��̦�*��fD��&�q����D��o���]n8���a7�JN`?9�+� ��Aj��Z�43���x��ۯ=Oj���q�3FnS��P�,���E�nB#!҄�����xm�B��&��d��V��r�G�`lҵ4H���߾��C:t%H�D��f|��F�1�VN��yH�Җ�9T��$��&�h�*@�p�X�`��M����6\5)F3���_Ȥ�e���������O#� >�l�]pk�<�ؐ�)B��c�ɵ��ǹo2�z�r^�(04z�G�;��N�\ؐ�L�ALe�}z�oHBl�c� �‧6/�SX�қ3�Y!޳�����b���ё2H�O�����E+e����-�����d��F�빼�fa�e�)�˵��+E!C|mw?���כ�J�`n2^,!����S����QL�����:�~3��'�0o�1�S�������݆~y��{�Gy�5dp�Xǁ>��P�Nw�4z�>�9�\RVvot�5/��>�~ �/�O����eop�5�Ο�4.�T��e�^�6����tဪ@��]�S_���\;bԘ�)��MWTk�..C"e�\��h��~?XQ:�{�\�Tw۲�����ss�XlxVHYEB     400     1e0��dcqj5w�h��^,
���(�����<aw�/�&�j�5�1��T���`&��������$u�=����h�L�n�l�;��T$��d�l�R��8x�h�s�u�8k-�
G�fh�'cIf� &��J��
�e�'�?=�˳�{���U/N_�鹃p��UrR)���g����4Ze ����I�2�ޓCؑ~��$��$�6�_����N�ٯ�W�P�;;"�G����/CE�u�������N�RI$ߟ7���-)+�Eb�����(��N��]R"T����ln�io�σ�\��~�i5P9fG��Ȫ~�s���\�Q�,�`�����ƭq�6��q�4�(�r��ɀ���Pڸ�/��m�'�]J��L�Zى���5u�ֈ�O�q���f��[I�sz���c���\�1m��.̶f�vpa��b]h';�Jى[�ȍ��h�T�b^(�E���$uXlxVHYEB     400     160�MCЕ�
�RO��s�����L�L���r�1��X�
U]�\s�������@ &)\DŃ%<�Z�Xx�z�䃺���M#Ey�9z��J��g��$�ؔ;�M��� ��3���j�{ z9q�c>AR�gH}��Q�5���������'��2FrΔ�����1��6Im�`�/m;���O�H�("Tߝ�g㺧�H����wV��
߲=2p��VuK�&��.V@*�Xw��"i�S5i��;1�/
�"K�F�"vQ�@S��D��	�M$����}90��AYN1�[��tk�1�t؉���ke(��8�L��q+.�6m��&���מ�G��s�EXlxVHYEB      50      50J�R^��ʬxn�՝���7?�}8��eˋsf a���<��?��%�7���4�AH��kdj��}�1����@j`�-