`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
dHCuy+uU8yXLc8VgJbi7CVYD06byihcnNSjNY5FDEtP77u4FUXSO1LfdQmgAnxH37MH49ygATeeM
g19VNdLOjXPZ7AoxjvL0ocD1Rvt+145Pu2Su6z4Cw23f1VBov8EbRnQlebWYTsXMdzNBNEKl2oCr
K3e8Rp7pOislSg9sjhCqcebohnjiaesMs4NWvZFS1lzE+apal3g/6iDqxCSc/b6n4JN4SCP93Llz
wN3wzWHx9+QZ3cD0QFusEJqcPaVhaK5rXM7dbpmBuNlpTkMrplhG0hRRANGW7h9fJSvXhkQrezFm
82CNN7lgGzMIJW9a6FxfwS24W+1WUsi8mjbV1Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="Yhr1bFqiqFHJugq2yglH35r69FXCI1x1dvUlhFvGLmI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18000)
`protect data_block
r+TBfNGCpRSaas7cWHSbG8R5SxdIiQgntuN5DPaCm+4+oqGXkRuDRWWi8j0ZSabWkqN/lf37D61Z
NqBheH/O57HCjQodwO1iPXMZZ4tlRohnJX/yEdTdfXQ+RWNG6cjB7Ui/mr9me/1xKhsMIYArKwtT
tN/PYciIds/Scvk94yx2Nd8ohYC5EQFjohlDd6tIhlnDRTurAUT/09HC/h5zQZTHXoNHsO4R2XXc
IwWU66sfQ2U3McISaTd1tMHsyFMVZ5XJnJSp/wjoA01uouSHbqStQRiJogdpsorSLZqjxB1ZxZe+
5/2+eOVaLnv+sJ/nKM8+CtYID/BE/y+agbtTiRkm4ZV5wHV/ILk/pxkKrGwALjjM/yqLyitqxTOH
seghQsRsGdGJWoHRtf6iu0z50WnyzWsh3O4TxcO9I0ufNqsfxsKeeKc6aanNChyst4XzL9QoWkpd
ry6oVs7jqG+6fT5wVMLK/oATv263Y3geIGJ/iQ5v38EodEcV1dVpscRwvImV4S6Uq3SfK1bjTVs2
ZGTyr2NvKegnzuUsEXJrL3yqqVpJm2o6Jc4kRf4EnyN5rwTV9qnF2/PEYADeINrkE1feRxim9zRY
rqHF1uUH6TLJcoUiPW2ePY2JIVSuorTrFZ5U53kA0aba4smBVrKuPNGOT03J2w9+fNCtBjX/BRqU
Kwf9SWRLgfOIYXb9yC+0RMm5cqWq+803o6uC5yUM+0GjMZCVyeQXClzhqZoOm/EpaZ3D1vxvQfrK
c4VB20xk0KmzxJeb5QVrzWh9nxBO7VTVgypco+ztBgQl7LKPLQ4Brhz5pQLf3p2zZxTSS5zG8Pwj
UkDVspMdTWHw+llFqCz0BqUtYAJ0hsuDVm6rVxn3zdSmAbc474YUbVPFy0ny/NeObHuENrSsfDhV
lqkPcaMV3ATdKLiBj2Agru+PGieM87YJCZXRWOpC02BugB12qq+dNs77A7NRBdRT5UM2lkldsIvb
ueyfSkuweYSR1m3UEKTSexyLmdKztqIxx+VH2ykR5Lm5zuiPktsazoXSq9nD3Tfyz1+eVhf9AGUV
SlxPS7zlxdVzG9daDS699UFxUWTDDA3d0fYntzHMLS7ASuTh+D63S3j5gbjX3aL32kAgz9OHmomY
LCUIvs22KKJ3F4nRbkCKBmVQIosAF1aYWOVyOB3XQ1RrTm2EkoA6c3c1m9s7ySuxTvwQjyXRaF76
WeE2N11Tr6DzpdDBErz+ipeP/5StcGl3w6vMAC1SSq0BbUQ9uWIKRQKFQHPhgLoS299Ogm3sWaXw
+OjlcFjpg/h+nUGGv1a0uM8gQ8pNBOI3wkjwBBPBgOTcns8QLW/0/N9WpfuITnIAl9Un72ytki/O
tZKC2Ow7lrWgoXCeL25MmWFndELCqnRyj/YORjAZLTajHGQgaZ/3RWyvmGVPphb/H7SzeMeVQaDp
phqVy+J7XVP33CsOGQ6ZFKt7/M2uk8ZqTzXCqEjx3pMTptMwmZLioCKLLXu3Rxo4C9tKBZovJoW4
xzfwQunvockTaZn166cVB2dA9dkzwQUZUwH+9LZ2HBLP81V0vr3R8tZ1/t5Amc6py1H/VBh36Cq1
PoG5emfeRrsn3qjjtVhG6/slTPsQuS1kT31ljColqn6gPl1XCf5M5ePc0uK+JCHPM4Yw6ZE2y1rF
eBXUmxKpikVVlwz7sj+kIbxfvvKKg8ehdi1TLb3t0elIVZzA2aGW7kk+5h8BozXsFxiG6Hvnow6e
L8dBmb/IRlP7RmElUNIDQLlfCKKE6kEWZu5Z2pwlQkr5rqmOIxfQ31jXzmkdzufZOmMDx1sTMsWl
cVcYq9hQhZU3RI2TqU2USsa3scsfvTQj0ccFZ9k//ygruu3z1rHGRBc2CrMFKI7/k2icawP5DDiu
SnAyOQ4Ok2JXXx02gor6R8ov7u6eHlpxESIgk1Nps7FL8b7y7g1UdDaeabWLjBsWt4sAqv7Lok64
HJjHkim4IvckS49nrLMtSPjrTWFQUKE4cubKx8p1n0TmLaerGPMYTR20b53gvN0aiy5lU84rQ4RY
kSV9FeWwlvsxhguTnup18CacWGndT8N8oqLLC9ApwL4LROxydY6CB2a387NjeYU5+awPjrZB4uDX
i7w4j5KWoJLsvD1nPy8TKjmvnf5LvWYUzcvoFa0bkrutILKUsw0aZr184O7MJ/4Jtr13+XXVNHno
272nLwdWcnf1kw/4dMFR7vu1dnrXvO1HUn3kteCI7POQ0RY5tlXLtgbqTW307IltzlaW/VdfFEXW
la6mqzraLAtJ5CTZcJ90dRwKxPBZoa6IGzEFdnWkZQjcu7wvLWnQEpkCeEhm/3J5qSlfIYGQZbbd
/fKUD2qsfUcqJ5mwhX2L8bnpcTPsxX0jo7yaBgzSnO2osKHh5dV1MEN6ZSlKvStNrU6bVPH97AGB
DqDhIMYIFKIPcDvxlIFctd+S3vAIjyOH8HBU3yPV7jd0u7x+fBJKkAWFzTWJfBNT0qyrVWLWLDIR
5UlJ8q7q0gSnJ3k3BGQXyk+jBbrT04wLTWatPnmoozmJzbuLdu3mqAHtNJQ9e+HSSegarxugHoJ7
tEno09DoBxw1C4yI/z0CI6SSM183BldGtOX9VkmzUiizt9EfkrzCTifGhPfUr6wuggNWnYgX2s5O
Qd8g0LAYNlZ1/pbHOcSzxSoK07SYZ6ykOgjDOFKJyNzkjex2llhWXLoAh8r0gEDgXPfRQf6Ejgeo
SXgCw9/fp3uCLgdc76SRP1872ophIzVkqemMUZaPIjUzTxCBxLwx/6qFFacS9YHZ09kY7cgNASW2
IjIJm2L2UmU4WDrSG/wiL6lp/GHWPsHcHbf0pE5XAOpbGDEKscrwctg75rJLmR24NBwhu3S7V1On
xqMkgBrZPPeJRd7+2AqwkfLJw7swRpJtdHb/FyFnvVhLaqNAUFiZZ7V4xGJ6KU3lJz3q600Y8inK
GS0NyUTE5ikwkcO9ldcdP4GnMAvOBV1IwOmUkEvmvjBTAyX3ofvpkUflZRMSEnGEX4Z6HoAZ5BEf
DRGuEeMvzWzEjW06vXKstyVic9QCeZP6IcE4QJsLxvVoyAfS0UGefPA/JaO6UIzpmES//y4bfR6F
9+vUiieCj6/os8pClYSioZPuxhiiLitRTVHR5SvsVjJOcJJ8+yhGELwmS1mK3XI03/qcLJjvRHgI
soxeZ36X9/3WCj04eesCOEquFD03kGwbxM1rpU8ZYNas3AkQt13lPL4ny17LIH0JdAH0ThjuMYbz
OkVQVtGUaTtsSTz3OSKAVS0WyrenmOuOUMyVjS7mXf6skFJVuygPptyvxComSo6gzjP6DxDfjE3p
S9EPKChQDRRqoTyLHgzxC+IYiuLhweWIdx3cr9+uJecRL3QfGVlLpBnxQns0Ed0HPU/GgrUa8Uzn
IN8yRVy8Tr08SZ07/ydh8BfpHVUxYFts/ojLFQDlGIiLtvsOIhreptTprWCOEA8bdYFkUgEGnOY0
5e3mO10F2r9PoSsdOVawrroDcR6OX79n69PsweIlpq+157sfJjR71EuKOUhmDz8Ee8goR6+UcBQb
1XaN9t/41L7uaPHObe6PnClq+FBKwxDpZ0mf6+SgSYYDWnt1oYBp/ltMNgHNOhouZwnL+xo9PULf
faETNH38ur4Cm/KLBt888lQmBaQQbYG/gaRrI3ifC2jKvgNQVIEakEyK/XzlLFR0Q5dH0BGfaF7j
D6D6H0VpVrdyEl6Dbul8WehHrSVoCFQ1rY0JGrmqTFbD/lOCq5IrlXqcYnlWcIkPwmfsbGrNSE52
bU2O04LRIV5EAM0roFJNUqcKDBWzAcb6aFaPga9GbBZn6Q+rw+8U6nHiqzOymKxr5C2F+UvVaRsY
+KO+1JODeNHs3klNMITSrIGDffAlv9vPTTujpi7qsuISKckgLYZeMyvk42AafsInu/Ff664rKpsO
77rAfsvmfoZem5z+j21457V1mo7U8eVPuPg4UIjVFC0WK+s7M/6g/+YAuz6lW6UJRENa3aajeRYH
QIG7LbnzE/Optc5W0sJhHO3u+lAmYDvnJs9HzsQZ9wgO0AFr7MHJSlO7euEc3XJCAHYq/6lCQRQG
fq16uSjnN2c4CNsG57bhUAder3fvXz44bV+HriY5YyApclGU6MXTmDWPIw7yeljgpVqNWJhweWYF
cZu6MNBQJuZrbwi3H2Keck3XzBHTq6oh46SexskPJdT4IuHSUSH09wa7+tHB0O/n75UdUZaNgwWn
QhXoft9qzR58FFNsql7yG8K6+I/aUKeboy6zulAdO3Ya92X+7i8HrNqWpVzv5XFSGpS8W9nzCpGO
/7xGHYxMX+6swmwdiQNlvdesEmtcobAa137qD5ObuJ3E2YM2XI48CfmPXco+1e3Flz7eI8L96dJE
ePeUTt4hJ7zOwatUe1EQHkIWAnoY1kFdSqtMYuIBO1xy0MnKK1470/GqM5ocm595YZFjc+qgmmh3
4wRSRW0fw+fM5Ze+1Q22yCIkV/AzqMdu/FOOsm2NIedv+F3hoG0oa6aQZ0WC4JZrxeyUC4Emfqtg
fUOaZt1dlnjQTiCrE1FtiofC8QSwgkx8Bk/5qq1BHSaB+ilY2bU6WCdBDjceNRmYFwT432OsfL7c
hlUTAiyk1HJRbAxZ87wGuiCp3nzqTq6TFMxN40j/EvxKj7I3y+tZo3AwdXpF28dJdftPdJFx/ToL
s5cHQMprijF2bb9TgTGCXL8FWdiRhFH09dgfU/NGgXhW/yBh4o7Vvf2ZZn5OQIY9X0SoI7WOj6Ii
tst7OHE3CUqU4aohLSXTE66hHwsv0a3ado4EGWudxrnAtskwX6PdefjiU3cXapdPn6FcvIKvsqHZ
KAqjZlOKXd/jVTid2PQVU+n7+VdKkVIWjZeFVFSLjuQDQDxMYOKvLU+9N0X0nSRV+5Tmw+ncDPrm
8qEV3s65cc+4Eqjlb/wqY8C070FGni0E92/5RX8RbOtp3cL5pv+aJ33bFAvNjEngDZnlOFE5rCu+
oZu0F5JdF+GeGko6qFQrGIdq17EzYLcR3Qw2cr+b6zHSZSKS8AIhwQlLuW2U/meVqWpIxWk8EPgm
+5dke6YVI0lVJXPzFEuTwuD0WQXk0ofxgfEoCBTtYHm0uwvpv7mU3Tf9WCZDET+hV+jHfi+pJvpL
oDvpM43bEPSs5rsO82KH43bip9+e2iSKw9J9RrRhZd+ygoE+FcORXmcneKGCRF/akgEnHRXBwKoJ
x8+czF706rhJFo/Wy6/3NaOqOyUZIBbUndN2TSOVsn/HPvkRbnGKShOSvmk0DT346RBcJ+jzlCbb
71p6mIeIVysM0k5cl8XOtXo9ZF0AJrSL/WafuOpOk+/HdExpO+3/msKt9MChrR9V+dBw2eD++zkg
B+jiAHt4qRWD/TAkxCbzjYvAtbrf7XkVtNU2tPCw3P6Gdaq+0tOy/wWliBaNRqCmhuOQJeIuf4gm
yiKjyhCm+XEOXv5bJ0snBGa3yYGHOss8Sm2SLDP1Ir5UuVtcczdlE6gjeMaI/iE6LAaEiWhUOsbv
6HW2Cbi9LT93RMAhNpIjuyKlOLZviyxQ7yjiln4LwnVNRJq30Qrbt+f9Kh8mf+sIvzOHAWT+RWLn
uFX8hfYMVlmCgQZebSRA30lK9heOhG83E5aVYJt2MxXBcP9faiVuaaLWRa1DGPAzKCZFuNa4q9jm
US+MTtgoDmulI3KrVrF0n+AknSHQn6lfS0gUVvSiSgCzztFZJloXYgFo6TuYUIh1TLSTKXvXVxGE
kQwyRyE4lGI5kl2UIrYpGubnrcgZI9beb5xl6PLRowX9QAKW9Ma2fnnZNJARCk47RNlUkG7TUTiJ
FC5/vbx3sJUU12jed2BUY7f4bLi/o1MMV3+Nnz9i0NWAoCqmkICvQXYGBNkbZw1NP2BnKLPQnxL9
BpfOGV+9YCGq5CFq2FDouyuPVj3U1/6Ide9if3TgJbLgasczTluiqUOlltjC23tADp9JNiTyAhJk
h+LP0IiNdZiQEu2QvymQcf9kHfdPMe9JbloL+xj8U7ZU52luCTMHfN39O1/DbQ7GNGR5jrr3eE8w
mARPeDBlFUTk5sdN967Pu1aHPhjaNUtdvmt927OZVs2z2T/aLxRlIx+tlSmGYogvYkbb4t8NeOrU
Q9Aiqed6FkMQK4cC2cLODzvKK9tkWnvbleDwX7DWUWn9ZRMRM9bIPGA918b9sSoBaKPeiRkKJwku
QuKTZ0bHaZ76LXNVvKTLqimtEmzMtV++9T+MOjfhDMyRFdPXL2OPqp7x3cpqGpv8X14QGHgYhYy8
4/ESy2WmnxJelKiH/37RIinN5aPhB58pIj6k5MVfCzL0Z+jyiyzdgelQadV8OIdHeXNiDn76D4sX
75a0r4bOdMG7FD1e/kr6FBXV9OpANdNecP2ILeSrsmOjp7rAyniBY8Mc+fYhxBqOykJVMG9JvVIY
tUHLXZVdmYZ9C07s5wR5pYx65SAtPCQyHfubjUyk3X1+FRSoWUfhC/kiR+unZMNFm2IeP/qS5UAD
s7naw0RYvXjb2FPGDKYlvtCjVjBz5l7Yhz/qIAC/sr5aEjgE189KCcEvJGzlcVik8Tq62Dktd85o
JWhMqfT2OXT0XtKBONn0MNnPfyvoNJKpkK43QZE/ATpOBK3g6X2dmP2+KhNKMvSF+BEhZCZ9qvyP
p3nLTvoYvrWawF2X+yhS4VlyJdeWmKFKGaK52+JgdX8eK03pSWQiFGzGfTSYG5rnGkC03jvZhh9h
WbAbCAIMA7SmILjMK3Z5Qr+6EfaV681IjZVGQ5NBBUb9SKiQFIYMrnLxHxm3uLFB2i/xf1sWLnaD
GDF4thFnltUhPMWKMoUDXSh7lAfFayEDp0idiwO/NQUiwqnUVoqIypvmQUHpcuTYb2GbAo5vS4Jy
KlOh2oLGAMNfAs575jgp6yPYEQ4bMvV46p0ytSpVrML4/sawFYKZBMsNcFRN54Az5b1VsBGno0Bf
6zarMLLb2KElHp9glwoBWVshNHY2mdunIApl3jMde1wbYnZOPVPYtziBO/e+lESKnzvdGHLZFpN+
eskHTsPCfqTd47m4iVN5TahV3EwgtbFp/LqCubD0xu6HerNmdnxxMiFa48u15E62+s4irCWgqxKE
8CS4x+JwaEr/RspJ9hkBSRfqio8D6htFCxsrmGiFyCTr6GxYuHxXr7bhoGUFx/eBjDvBVG8P3SmH
uADMcXwCIUskg7rZpvD+6iqLTLlmUMcoyschxS//09RAT5aPzG1me/Y8N0/hmxq22/loKZUDrl16
3guZie7c09YrFCJJBcXaJzKpHBC5rQBH0Ci8mu8ud7izKWmCMO0+e2X/VxKUPk3rguY5Z2egWNr1
/FwJkOuPRtxbNeTcH5lq5j5jDmDZpYGjLbSnKQBfnHeqau+oKDd1p2sWlLak14mW3EOiQc8YBDa2
APJXqs8X5Ixu2GpeA7Hh/yZEiPoDb84q6DXRj9M74Rl4gr8ypOdEr1zCDk3lUEA/EIWSSsCXvb64
gEBVCKMh+S7NpF/LFqunZ51l0GSh/PcVtwvRAjEj11aMP39g0z+a4g1b+E+WD5eZXG3hYsm7ajTO
Gh7d6W3AlRpTVvLKSaeMzqC9KxZImmm+QGFg2p6M9z4yHuTVjfmPnLr/IWDcFZTSn18YppEsWzD7
ZNz18tMbiE86xUZgw1zBwSy0D/ECogMAhSeGqvNaN6qlT/RZddOjOPN95JWh/ivB3YfPNC7AG8TZ
cNF0iuXScRI/LF+fYEYZLQ04CNz1hHx9MjXnSNzK+uXPLvEWTQ/iA6zOfWh8faBdy3lzV1QneVh8
fjuOM/JLDTOnWRx/IeKr908dQXlIRmLyuHhdARIGVS5diI8dK3Rjqgp1FWZKg0rsIXmuGH7ntufo
1q5P/683mUh8dg4686qOjp2w45DDapdAnB6wfj+J2wfAZrN8+iA1htnrU6OouzrKXx3UMhxb3J5l
SnosR4RXGiabZ+AsFy27EOpdM9BXNnghqMFgJQDThCocq212jhmXpB5Hoa0a6qFAmbvM+a1qhVDi
wtdzukYBjkI9/gQUuLaAWJ+zI7OsWPcZXq/EYOqvTJqD4jxe+0e8Ll8op5xqM+g+jHnckUj9eTQ9
UgIjXhBtYoznFdH6o+JKrJr42ne6+QxsFq/etgQrH7BHLjNdul1LN6j/FNWL9BIlzZxwbV3sX9IH
P0iuzrB4MJPpVAk01OYZYgZXr4fS4ps+Z5oOXx9mk7RORI+yG46dIYput1iB65YAm85MLzlrtmZo
hqDN3Eaq2YBomzuiOatOcjYoCbDihvz3OVKkDW2Efq3MlPO6JPn3upAFNkxogSt4GtQw9zSr9vNH
Jv6esxoFQGZfcUg9b05widVFegXPFvKC4ZJOOPc/2QBa7pgAPjNCfp0BGujvT0X1U1NoY7GqBFCU
1DEl2dEdpaeBImN3mD5B/GJPgvkzM6jCp/NyvwPuLCIrXi4/C+52Tia7urA4ZI4uzAZw4nTL82IN
FoDBFI+4wW+2Jdaim0LNKXwXjbZZ0/LUtbrEORN+iM21/ESbbESoa5DIHKSR1um7zOf/e9fsotQ9
EzCu29mha0GYGXf+YNgj6zqkqN9Sj9zyLbao4wlK7Or4krJh/9xi4tGdRNOe5cd5AMV2rW3F+pq5
55BPM+J9r7bBqnC8CI5n+3W7dsbyoAiK2vAgCrzVck+Gz4C5mJDK7Xjodnv8IkYpF+ZJdg0LZLxx
ev9hcnyqDitt9prNcDsRmxCyT7yZ63XS48cyIgmXIESW9E75wY2Am57V1mKQ4kqzCtSLrwRQPVAP
wg3kVC0dOJfXuqkuJPiHcQErQUVMIBwDJyHoStSL0FPhExctkpWJeQFMqjqd8LtA+5nHnKMaf4ll
lebqqgXKsSU1BL1hadBg93tRiD4ym+h/g/GMvp77I6NqAafZkSAuiJWiDItWSbnyKZsfXT3d28BD
POKYqHXTfcS3RGNZgwrMLqNJriYP2slVdOQ7H9RJrQ42flKJYZTKA2quFB1i6isknBdXWbxuD6yv
wJBFLbJz4RlPwtiIphGDVvOFiMuPbFeJdFzZQ5+u7Oke56TKzluZuuyJTZBpZD+8f1yE08mykfh2
czlm1ic9sCVg/lWhDngIb9N6EHeYiopLBmxZJfU6eJa88O19fHZjjNZxgo+LMYM/zVuNMNXbNl/N
z9RUN1xQ5LPYg8V618RwiA6yYyfxHePsRa9h2EOpqc+6dyb52F6wTg3rug3lWg3B15oyDyOsADfQ
PXHh8UymGSB8H3vHqIDTjjXY/1YILdn4pHtaZw7m/c0x9TwIS+zbiyaH36qOGt/AeG97P8vOuPju
GtnBIvcTlBAZVvyCfsaHTnZLJY4YjazVj+KILmt2D2MR7UaU6yFayo5Z/6Or+mXkSbv2QEy3g4mE
A2JZdRfgJeIxNhwocGRgzWgywwtmRmZQXMbW4A3/zW3s4WO+1TDIRsAu81aUI5w6tTVRal5la4U4
CyA0+XjIOY2jrgee7zRMkmfF8zwUW5R8+hyUz5trsWhxG/Wlb2hnARP3VMIk6IKHfyjdLFH6kYRZ
n2ujW5Z1abUAm6htEO57dtjQQSpUZAJHRrySRFfh5RKjI2We4oHsUAUZVysSF3XCV5bDTF13ZfnY
COB0x5CVuOHJ52IhaBzSxwl155hCjo4PDKjZNhE/1L8pll3GgjIyNGT8fNPjqJPGaYEkthsX3aLf
xvl1bs7Fo0hxYea3gSc+75SB1d8PMvr5ZftzhPL9hzn3+UFozoCKxDmoB1rDu2x8rWaxbyPDA7bI
ywyj/gKVBf+FkcqOo/ByG8pVHZQIv5XwXrs1Znefy+lcR+XRzOhU7asykOsH3cDj76/wf0Svd8Ns
9I9w89ChbDc9C5s7V2NMkQbAu4yZb37De8VkIE0XWa+2WIlIGFY8zmPfkLWfDUubrgOeY94HdDmc
g4cXFgsRwe9APjOVL/iTR2dHY8yZgkqWa8lsd8IKUSyLWNUGGxTVmI0KUDCylgFRFg/we+cq9JL0
U1NHzjyWb9OeyHxmO86mp5IMwWUhuj/7pmA/Tk1huknjBf+mvn1PWQQvqMAX6arBqIyxZPAJv5/Q
0J/FH1HLP2LIX8uMOzbO3a5QIRAqmMPHHXO2xpGIohNHFgffDGcVd3uNKdE5A9xjB9TXzrgVEst2
R5OyUSlmyyU4m/aNYBv/PE99C5CBgHE2sAYL4ozqBxortxzfownLXMtrvvzPdzrYQo8qyos15jbS
zsQaRckHftFFcE/4ZUuv4A+z1wxkfICr32kCe2EfB8RB7MFoD53UiLnkoXdc1CQnZixZOPkDlf+L
XMaUT3rsl20xfpGa5Hze/jKyW1nqmtTiWocyj5s/8XA4LLFqlZTlcNZXu1b30+FKkO2FJX+tkbQY
Jjry9IyGjZ5tiu2CMvaknBaAmwBPI3+M5Me/I1MHUKb9iODh6UO0h7SD8mADT3NIAKVxmN8KtNu5
Au8uYaBVMaWF1DVcFEtRnzwf2CyYX/F3Xy2lJInq9MWZIei9DqfMDAG8b8Lg9B4NP0p+/twKon/4
bhKGK3L1wj2xI0bEf4IxBZQ9ZDIKYAyYXTbVsS2SqycFzBVGAEc/BUsoRiKIahobFyZxtMANlk+m
rkvycAdtpM9jtajaO//U8WAUtvOhsGst/E1IHrz0DajGQzC8sps/ueBjLoDOtBbYujHJPB55NrBd
LLyNuqqcXqCKaeJ0qTbUHCe3vOuc66C1N8z+VUnJC6fvWQ2wWVPfNN02242t5pyolQ3Uqti7yr6U
eOWE7dQEya+k7ltRS+1pSfClPFRznzO4ZA81tIerug9DbL/Lwkol4acta23iwUWwEvCdzLwhcOS3
fNGFW20W4XAm365Y8KNmtHu2SBRKhQa4Z10xW4nkVhxNsggpLybBV8pcQbGDqTHE0dhj6d6k6MKL
R8/Bg2p7PXJYl1knC3QvbHoHdNs6xxGMkVSFwyn2DV8vLvWmAiz01WCWNDQWWEgmPHZD4IsUVqni
O7VBMCYlCK4IyqVIRY3Iy3Grh3VtcXOwXRz4IEixiJhyfqwokIzpAAoxeIYnyWTs8TecIuA7TS1X
Y/0DCeaERvObqk+KAc094gL4tD6XkD55zppVIYB2kumwMxkwqouaWHLdXwz1pD6HbP6AOGrbRoGV
0/fJewx4q7NCqa8Bykz9xzvThc7//n/uHHVWRr4jas434L/tF2rxs9LGaeW043CVBx3qKqXNuKD/
rL8PkYklcRtHOX/xs0CB+WumT14N+3zIBGO61CwglHmVopv9QpMcNdrXMsYP4f1FRXep+zb+LJar
kqr7aHNHxbzAt4xUmfz9Cz/UnjrLICylXzpQbjtKUGkncYoljAC1riV4cbT8tbfpIhLlD3f91yNX
Qrx2X5FSDKs5cgusFkoLpKSr9ga6QqQoV30uGCMgWIVkBsJvE2MVozIzeuUeDAW6+dOy6r8SavNO
7DbMzw4I/EhF7w6dOIK0oAYF4o3z8dskOAz3XnuWUHnBgKDHvyofOTWiFO39L8RAm1/Lu3wUN/6S
Km00NJUb3pbzeUx/+hfJpgwM0r8MHW7K7sEzPe3SZfEy2M7vMCiPH2R+1JLa5CTFeDzsJOMTkBTX
SCLvrCfDlktEQZlpo2BP6bgxnOby34j6Gda2SLv5zrv2k9c/bHLjUFUdBoYZ3vlK8l94DGfmtIj2
Ne6B0UvjdNa/MVJRfBnlQ0faTeeL4KOV+W2iwvRmRpALLApnzmIM6br6PzOpQHtRgkGfNdXVB/zl
zIQAHpCF1yMHUP3QtwgGNAJXe55+Hhvbny1cdk0QY+kzrWEZG1QkkapmDZ0nzwteacUdDSD0OB0E
JLDbb3blRSYkBsEsbRvlxTWPCS0AHJES5EOnBkyfSow2MbSl4bE8md08LMNZ6LaG2T2gB3SPsHck
OYxpq8qd/8Zcqzwo25y+5t0OYJ39y+FZGBXHqmQkMjx9YyxfcCSKmeZFYdEbTQ15SdEh13jWIdBJ
Ixj0f9dOjldK6Gac6dxz9Kcrlj1VhEqzXRvws4E82umzklwllyOsctwzzpmZL1z3fLIqLy8D7ZsZ
oz8k6vNnpkXyw9yTYs87/CSX/wYO3r0zA0gJ7NlHw3wQciEjEf3UvXtfK2uZGJVQZ9Q7amiXsM3p
jWQuIyy4A2ADjvHSUdb2SlWkHlVehZsTfO7z8KGYJBQ7uTqUTL65Dwgk2VfyYkyDCZjdgdxyiQC5
zkG5ubaaMMihgTJfEyp3rGZdPVMKl5ttmHLmCOugSwpkfYsCL8aYWQYjfG+8ekbqnj3CYMKYfhFR
l67odSr0lDf6c5Hg70ZaFl11smXXRVawbek+n7jv3mIrYm4iC2aLoTiVvR9OMKkZZX2K4ICgE9Yn
vi4lDRLhewD8rG0UUHBNJxRKlpaCcuA0r9w2g5Jebqydlp9P5BCs4RVZHLkoRIUFkKE6O9qeXvcl
HK2qYLAvFluez9u0Cr+FCxaa3Si920YVZZPeEv81gvgLU7QAmtYhwVQ2H1Nh2qWf4uYHDYpDOQVl
UFuZS10XwlfwXsG3NOqnKnqjobHmSFw0Ue7CNPYvu5WlIgcMqqczYcBtyba0Y589HjM6cEbqPcqi
yOfXeblZY7xdmggGuhu6DLTvelNx9N5h2XmM7Zb8U6UGqkfRXchjk5Vd3mYssVQQs6rxNXagVI5p
LpXWrv5rdL81y+XNLgHMW7hKyQafY3LOri8izFeBmVyM7JLp53UTAfO8LTMTC9C3cwWqfFjnjvZk
vfb8hkvgx8J80BQB0x4VJwSVQV1nrmeeIMO9a4EDl47BPTpzxl78zrX0Nspw40YAI3zY/vZmGgbS
BeID8chEKhCWmg24r6IRxOtTJcvMuu9hVdvYRrSRhjWadz/DJ2eBm0OhqcCvaRGQCoqqfpGBY666
Kb7jxD5rmDmc6RXo+EovJx/0Wfc5VQbcj17e6K39P/lTDeXtkTEX0tyZbjOevQRBbFjcCksciVN/
PcpRPGNChE4sj/rY4v6OmsjA6v54Di040/6DMf8exRKdD4RXoUTWsrkGsKg4XmObLWZraUugodkQ
eiuAFpuzK8nzSyLD8cXE+AZlfHb+WS4DXwx42Jpt3M2BQ8JFENdDm5Sl4FW2b14InUov/Mk9mqFz
ueeqbO9P6H2QNr89EUDscXZlnSdHIJhpVW007lWgtPlzzxdpfXQC8Lpko/U1v39stw5xEa16nuFi
x/e+xagCISFofZBeHCXKfZe6FzACGz0ZjwJ+jxyjCw+xALDg/CCxU424KTxVJJatGhv3qWxtzRJ2
rUlhjj5RHXtZ5BNYEg8d3qIz0YRsEevSD9YD173fp28qdNvfIii+u+LTtzgXaO5q9OI2mdBE5s6D
m5iiIvRJSCI/0AYzA1i5R3UXDu0rhco9xUlWBzh4NVRZ2kj2G4mqVLLBDSo6t7g/QFOWphUC/6Se
5Z20aEaDdfE7Ml0TtXasiDiiXEBoDICfNpKbBhgSGw7bORCjlDeQzoNJ1Lx7Zj5iI3WpaODCQgO2
TW0obcs/A0IKPYsQrsDNZJRS7Nie6cH6qQev+pmCxvqi5SNASnQ/hkl7t9vicOZhgq+CvStYjeOE
C8aCBxvp9fBg5IbHj9oFCky/9irpkEbLi50qlxgvxKIhcogahYW2fSPzOFkRX1lIitWWaShFCxCF
I8MX/3JC7Tfnjya3xgilhOH8sZ5p6XvC/0lX7pjb5w8FG6xdTAMh/q8SyhE/DNYZ6zZ4VvHacdYg
J1JcJ37F7OuievWCRSQfnZ2LexVWELqM+m5yNPDidOnMHhk4E+KydSbUyXlUgppA+4r046wf1rFA
9Kj+JybVae5upPS/g2gi0PI+lhh4iTbKU66sj5U0NpbcSPZtPJqy1uotsHTVUAO+y5AFZrALBB+U
ChC0SiaeINJzZ6jirVupdbEC3Gs/V9tOhk+Z2r5HcX9z6VdAjKBOOXLFpikTZXJxKSzKiLeTSrwU
E9PeJUdw24HUSdh4VVg/jY/Bzse6YFsxjC2v3A/POY87yx9k3Qobu6I0YsfuGzYPBRWb6QYTpwYh
qG0EW2freonfsem/fj+YzAjxKdJXzvrChO06KDZAUsDexIGFXkA+MlAK261LuRZFHHSkhFulKrtl
bkqlg4elpzdRw4gl5KsrW/Jwdi7S/zSY/lstobyJSsZAg6RiJTEKF5pmvZ8pX5rMMnzSjKnWFbgo
y07Wu0qZByT6bI8vDaPXKD1EAWDApA4luOUll66U72bQb0SCqvnKzwfGfvhXFgVmV8Vyic0PlE9y
7EaMmhqHiGFUIA9eotubfDmW7YFBSgDn9gA+0GC//IkILUcWWnNg3rMgxa6Ba9TfKo8u78CsoJke
a1CDBr+6ASobF5dVpfpDLC6vBgZnIFJL1ZK98xpQDVakrtsmO6oIDiib4eUO1K/OcWnzpmKHgWdM
tOEO8daKSEMH5scBPZJu9v3q5KySz4GVqrz1vFqlUQLd24Xx7+bze4CPw5MWCu1k1M588XwiA9i5
8rOEKxfXuWuDz9lAp+PBhpTQ/iJFL53Zc2Co1vH9RjILyHFgYUPh9Ag6UvGTzRvcADp7+rWvN1Fj
Ut7CuWs60G6op8Z8awWM3O1VAtksXiPvN5D4tdoZZb+UFZA/kIpLzN3Zt8k+uwnW4Er2j/M/XmxM
sKJTIim0iY2bWgU1H3Tz9J7FbEbVXvbzmR/fo5MUk9xbWtMnfrxsicLgTjUQ0McLC4hNyCLjf0mz
txXhVbne+9GjyFN70U0w6Ov5ea0ykyO1eqKjjopcR5JUUuCRcwNO6pLN2BF3Mlc1rBfAPkVimCdl
dLzZa1k2XKxlPTW2KE/fCNXZyF/qDP5qcZ9oF5FlhPi0/fLv/3DxIMr90ufTLWSvBVdsm+qce70r
UjKeNxBDFWhi5cHF5GMc1k5QmqvVqob4/WuWXnuJVvZgq9Apd+aGfbGyZz4aH/sTPkpTfEF/Ojq3
X9+/N7tVE6B7GZFx3bObAwUDz5KWEed7jUYUc1rUbyF4ll/skWjzABiEl/u19CUs/Wf3tRIiRvI8
3If+QbJqwnfjeymOm3Ab/lwkvYjSLe+LVikUvhYISMIFzdl26+z+Bc42nXPG4XU9Z3LGeA7171+4
ZCdtDg4YIR4xTMV1FyOazZ9mQagUF5/TAOMRD/9Fg0RUUk5pw3jEIgsOCYaYGdf3/fpR7jjBP7Fo
ksDDdGG1s2t5QRSAg3rYBsgD21ZOQeMQGAmdR22w66/DlbSsMcFHixY9Qfy/lTtr3lbMk7fiMtBv
B75eMFY5ripGFQMSH+r8MDGzuisOzHPDYLNo/pG/DUMCZcdBeG1nRQ5INd++R2SnVtvsXjXZyazh
2xP+Lk+44Jlw9Sx9oGoB8/4RVl8Kdc6pawMDNZpV8cmuXpu4rNTlxKpJd5kdSWDTDcvkr4vxXL5V
nNd6/RVwFBt0qEXwhIS6L8vrh8phxo2ox0f4z/jnQqqbA3/1F78yX1lYYKCvvMwWnwkKdEbuO3ro
zTca/RrWjLLfiNGn54Gn+TbKDX/9RtW10NcyMwcnc9tt/kcNX+lqGqjiAgNIzm9L7QzZ2qr3vkL/
Ss8wNPOsIr0WPaXPZcXqdCP9HEcBYWk0w416ZxqwS4xh8zkNuXowiCYr3/PIGrk59ZVtkIX1lx0t
tFhkL4ljsDnqj2QFjwlnnQfQf/3QtuV5wdP5hH1dizVTSaJUm5p6/CR/dXlgwDsHqx2KvGSROENW
cLe1xXk6Blq0y7wYIAFdGH7wN3hlx0a6cuJ93TfpUZe+tju65eIMDjzeVKuCNhmg4NkwOHyuLp5t
53RgnPz80CkK26CQWDHo7pZrLTN/V6dbdUQOyvYEEzK0MZ8ov0sKTu+ohRVt5fSfIJ63g4hzKYL+
7hCfQjmxNJgvpaPDcNGNi/jvTE5Qgbx2u4WmZht6MIojzuGffF9kdcofDFnog0eMzVQuEuz4Lype
xaQmEmsBeBNSTlseYugpfd9GviKYXO+l+sy6K9MwbCUeZrSTq5kmE6hZkcmaqkEpcdt0S7zyny91
yqpmOWCF02K3N+JawDdoudTMK35vYUttuQI2+xqauSlxcHxJF+v/qMDRbYchSSXJiBaYUXZ3M0uC
bDVqaLTRB7cw4NzdtdiIIWuOzXblgZRekGU3FOFzp9ZrkzJ3tJt6Xp+Shuv/O60V5U7YlDt6v3FA
CyWNhv0Ewmw8go6JzEjLKg/vftwlpOnnPvcXKqTF9hcBz94VZWl7Hz/4QASmqEmx/m5+JdOWoots
wVvozwFKMPuERuQp+zK319ZWQTNggynkUQuMfHAkQcX6rj7IStNs3yMm6ZFFYppWcsxpEXI4Q+4i
/gbyto8x+k+g9/wDkzawyYwromtMoPU2hI3XoHEASGuwI4zQr8bgiaeHM51GwRVbNWq3h5oG3gT1
vOa1OTBKZSQIqtT9aQXXFONDoqfNXf8ehyjOPUQD/VqniHZOQnWr7EATVQlUB9wMvvXT74la8oIJ
oRFRmrdMu/49Su/IXXjHZVUT0hl6p5M1hxfxk80XeQUagQ2LbNTjDUNBmHN8p9gmfL8p8bee5688
56cgWiNGeezn7ZHaKBrssWA1ZAbiaZ2dAh1vkcAwlriJns/gm8XgFe7jhSsFzLzRhKTx98qWF6m7
Eju7jgGQe2gcDXJMgQWn2ONwg72Oeehsv0iZp8njml1iwzz5Q2PXKQFjU8Xl+yi0chZwdX9eLtvt
VF4dtVDwoLEE9TUwq+uXfyhiGJtJiz/Pee0LAW+ujG7lSd18pcDMYDvTo3Vkm4UCiZI+oh6QFPgN
7erTRGTORX+XiEbd1aoikYN87Tdg0R+rLDSlDdncZvswP6ry3PEjFsddpO++9VAJ9M3UYMkTaA3a
2tiGLQUc3TSO132MnTNGP4eWV9NxpdGgdrrkdy7p7ys8Ed0MXgVrkFSHUDVc1GZ/6saB4j7MvanN
Z7w3ExpcnOftZqXsTkpVb/tkUqgga4sj0XD/DkiiPgNJz6Cglse/bIzuXQftOvs/kv+hJHiPXAUW
l2m3y99gaU9xQyuPMr/GgGSd/ZNVfar4zbWOcC16w7oxTYdR/3kDSj9pjYogOu2LnnApiCc0BTGn
oS2J6/IA3otuWvaGhvx4qYoJUY3cJrBFPhfWWS5OKE0tpwv8j33tfi6b8cdNdkWNjUxDf2i8+ZpZ
2nRGLMizkwxY6K4ucq9Iet5BQMRgbfCz7yaGsgGSYGY3aX16DFEQnnSt4Osxn4AdfEQ9uBwThzjV
JhPQIhCLN4BOGbq0JjM5QWS6OqE+uBzPD2c78D2RFHb37AjC9y1/c56DatThHfsM69w3Fi5M8bUB
wItAFivoxIbBDdGtJ7lZrxz7XrjYMWWM3gkWXCCrUW0pDEyuaaMBb9iwOI82dzsxTUTHDlqpu8v8
ZAU6dmtmPTrI3ADvwvOoIlh8pbRSvDtFSn5AkBxIMh6u1JtGFERMZYSFt7/w9Nn94Pqbte2aIz0j
WiDyf+Xf7pY1CEkYsA5DEjqim/Z4TkcCcogXPUDJUz1aIyqKGMpWA6S7UH+F+BvVOp25XnNOo5iZ
rFe8+RNKBEyyYRyy31XaUlmRU9YPA4oO8LL6gKtUVkNj/6Lcs08JR+9Krieg0NG3YhqV3ODMsmC8
HbNcsOSguK5TNVOYwRPzDy6o8EPm+5MpyMbcDDHcEtd++nDuQYTEuC73/c/WijDiVPCOmC12zeLI
vBVnQrSYPt0z+ELvZ0e3zQ4Rwh7P9ftwzFpj5h4z9WfCmGMwAaAHikGMDwhTNU0uMroyxgzNjhVp
5SMILtITuLLjRwzqvsJelBZrS970zY1K7+C2F+W7vrcYCSyhAIqYTjo2LiU74Z0ubKo/YZ9tDkNm
1jcktsgZi4l9PbPREwhjPB70FLE21SWPr+pn0wxZ4svkqMe5YdeMfz4Fdrmd4/WxAJVk7Ebxzmjh
yz2FkwtznK1rM5O2MW7zfqaxcZViL8CnuM2QNYbaXJlcyw5kR5T84mhkNdugZv95SouhUmasPLEW
+ntLxNp/lAjKArVEtMAguLf4RRTJU4piurWqUDky+wuLnLc6XLCX9rbbE1wprffTPFtBc3jn1XUP
wJMNuNV43hIiAQskNrFcKSMNXIKdIWdeno/tSir7PN1GHLGfFuz6z/PRizUL5IOTDQiyUm8TpOxc
PWkbg1ytBuQILGSCqlHxaGaMVQkDlPXPFhUKvIKp+iCBLnMOiTpZmpSzD/gg8ex4d5Zr2tO6tcAQ
23b7bz9mepeqC29ERml6H/Y5/yMZC/SNROPd2agUSBPUr0C0q5J6KbnZ9OrRHHedDZhp9k4DnwQW
/2qJpTXK9DLgM/WM08B5n8pbhflQevSgBYrfkQzW1thTTuCfR5R4m09jcz1B+roSLO7D51s5e/+u
VTm+01HGW8HOxHaMw7iSxb2z8oiH8zoEHgYbCB5yITJMuz2TG5bbv4mY4+7WXsxw6WbSLSQWoMQT
rWCKmjstupXU5A5xgDDQAxVJfgaHho/+BvnI8PyPcu+b9A1hICzlTr/zpuEQ5cv94yzirM+pfddC
+mp8XvPibn1nFdPB8SweFj6vMyiFlVgUHXU0WNVr+gPeEOUP/70+hThxKvxVWvW04pVs9pr0ou2L
ZD+dlRWDBv9w8XP96CjA/4HIMXbBapmBQzzkeUSqOCBCwlA/PbHlYM73V7i2h4RHkbqpGO7nS8mc
CEJkiWaEYp4w5JCy6qojpaqOp+ROuKeqrOJuL30iNo7OZ4byRbJWYm22KyjvONlH3xS+xfesxlPU
IuISiwMhl1ALbOROU3wTTwtQ6XR/2vYvlLvp1HsLuRos53cFM6X28NRILDLJJeOpMyQ+uBYo7IZf
rdmylISNgje2ftBBGMgobRDXmqiHiFenDQTl+5I+UOKnKe9X5SACLpSm6wphHaJ8+EvXoPGiTHxv
NCFnEWP+NviigqHEAU2R5w31KrcU+4fxwAdN4iFWxRmATfzs7pt495rPmiFnZM827aR9M9oJ1QnC
OGMpCsndDhmSIFD83nYz2r+ukPnRWNyLYebE18yWPmFPQhNfm6qh3SmrphRbikyEK8gmp8n5Mvq7
x6RMjp1qtLz0ja3LQYqg+qPdgFI2LBTiVC3jcpPlAHkgDoj98NCX4L5IQUjX+V3mBCeoJhSQmnhT
vZEh+2piWXQ413zGp25QbW/oP+VkDFFEt/c+vqUBPcnHu/HUwruEZ/ZvfWy4NhxmkJuCtdrJJhi7
PNaSlLTIRy1coNi2oFYbrBfEV0fm6WP9rAaPiUragIFiJSXeTlrX5LE7huRiKEKscbCo3M1JJwGA
zGQwOi7rJ5FKc+xc8EYk2o0pJwlu+xk880GAN2BOH7Ppz8Cj4OiFxD3ckdJ+hBgFbUuGGKYP6oPZ
XN9c+TehpNEv1q/NgNXg2FAGt8GU+K4TZla80SI0tQShRPKfA1ac8Jxtw3fC35M9hgGidxl4BUrO
JfQd/kNuFPu8p9xksGdbDfNIWcaxgV2abrDxXciC0FX1Bf4IIgKGzwKyuI5iLK4wNjZYcy5bMZfH
0ISBcnf4k42WhIgwj5NSV0uxp7Bdi8qIwlE26ThJXDFxMFW8D6zRNjxo9zkmfAKIcIegsH5qyjm7
1KDKOONluiPV3UKGLaZcxGXTYuU12Tywz0jVcnk9HRpLwIMvc6/lH3RDOtLmQwhCkihF5GqJzNA7
HOGH3TIv19I432fJbKSNqZqkvbCwuWuaCTLp3Uxvm79RUmXD9glmk65+jjgLFghiXMp6wZxrgo1J
MzbuhAK83YKl2Q2azQ6svDHsTbmitsBidRtGJOKLC4qrR4O8m6GgKcZ+K9gGxiSAvfDHaMrlu7Pq
XhZaA2KGdR6JLPktU55uXBZj/8tjWkNZRbJQTOWuCx218AcI2x8EH2WGYW19ImMb5Ip9Hc7cvRUo
dWTz0Odk4mVluQ1avHasskIQaPml6EzSp4I+eE3nLEzayr38flDMDfvrMtzwXCmoS892BICYjUtG
O2NtFzmOj9fupmKE94+Kv6wX0uBE47/ripK2t7JgX0n/mskW6zk+I7/tsWhCYbw2i/ndpENmNwO2
6oS5+1FGZ0vLihxjFUvLZ6peDgUK7xUjl77Ej4WqUoUSiJEm0y83EB1oY+KWIrGWqt92Bh0WvdlM
3jfGc+xLEFn8sNxD9DwJDevcnkz0sw3LFh7Z+RU/oiNhrloRVONHXCJdzcfGNPWWSQGwJnbHOnpg
Od6NgIBxY1zqbvQWiDTGeYA614yDQtJEcPfyF6nZ3l3/YQ2c3beIFmzyqzAhldjzBrv53riyyRwn
ZtEZTST6/5h5isKEqoummpXNvuH5XSAgmR/LcZ1FQOzsgsB5U4WmJNZRSZhOhYRShBRt+ZVmX01y
9WRzxAAW61c6UucgMaE5rjojPq4lCP6eFK5ZTotjCbWQ3DZzy8XsGTEgBhDHkhwF9XakSdZWNasd
siQNu89WL6gUU1sB/AzdsMXIGfg+pMsYASnEdMyxlQb+qkGesv+fObfcz4//PDwk3a8czV611sLQ
2lwAWB8NAU99u8O+UZfDkOOy7uzhgM0xc7QtVTA9imWa7NjxN3VzZ3j5xV8GMkkGI7SSG/dvgRoZ
2NKucVKoyY0lqa1fH4BabKUMC+TAr0FdcqaWCjqD1OnLxBfSxKUpOalh/eCvylyoNF4wbODWcCtd
96qFc9h4aOEHSGmdhaaY91u/rplfkO8NNYPawM6PptPy4L79QI/xCD/LJSY8pRcpoLterN9Qs2En
+raT0hzvloNyhH98ElRv8i8iZPVf907m2FZ7V/MdnUE8D67Dp6nJR/A0nRUbS245OmSl14GeK3s2
VHQtvINsCuyx3S1gUQZ0g9b40WFkN4eFhc1UvFpql4IF0tXQcnbHpXJLBtZ+hJrwiwwSt2lnmGFZ
b2rHxCo/+NpejWF+IqXlcYMmAR2w91bw1DG56t9Ul+rx9yKRAh21Gtrc1j74qcsSGHTff5T8jM96
x/6HxVkYAbhGO3CT0j+fr5s/eQ4CSgRZKkjQQtbafvMMF4YAUroxG54SsyIZLwjFiAk4vR9kNTud
RCOpR/jdw5T/2aWX+6seSB8udc+Z+Ah0zck0W/f6Qc6UoQfj12AQDuIP9O/mgbgOQZ3edemIckdy
vjGsxxUdNOypWEJOFeRqfY3IIjJH4GQl/uRbS6LNV0Oc1yUt7qfbXNe0heN5F6OmT0wu2h+ZWVwi
vJmGQFFMuN3cev19Cax/GEqEkGU0Xgvtqdv6AxMKZil91E9un0sHW6HtTvB1C7tOCS5hQGfhZBl3
t3GTQ+M480GnCmE2idkpoxOqlQ+8tQjzt0ZJ2+JXrJQo0Cf7D5toXtPxgnXYGBeucppdDDmrSpVQ
IAmexFnT+XQmDc4jRnaaY1TyJ/9JlR1FpJveWciXimm+E1wLQcIf7VSGkFI5p/NRS8Xx/80ITEgQ
9H+r+czToZZNNqib8/0eCaUzFMnR/zWPPuhbG6cGinaAsaJlU5+XzZL+X8krgiPfRtrWODhETXN0
n9ZrW0q0Z3E7oB98c7cY8ktdTvqKeTy9qrDparjoJa/ZWNxGMt3gMy9SON60ydPxnEcXjAHuyIEU
haUoa256UsIb8Sx8FY37g+IzHGbY6QJGUv3l4+F5B/ZJljNCLexFxa5b4e8zBDGDtv6JJEARDjnc
VMvp4XSNUFdNrBoYdHSEmw2pSseJDGejdGm659iFnGVD+N6smn3yNlhqUt9UJ7Nr7UL25g2dwkTk
6lnL9zOHX3Nb6j5c0GwfpDMBEXnHw2rZRHhSz3eyt+qZwvHPs5I/URa8wy7/pq8+9A1kd2C4MW2W
+pGs2bRxKfhQ2WaUDAEtPwstvyDaxPGvOrVXD+tRKGAGXl39ITsApb/8f9QnFccvyczth7Z+5kAa
A8zxEOTwu93xdTFF/XifnbYH/CZPrnEokYAT8ZbBUwBgCnFSQGwrdwtBzWRu2Cqbjw/n6i1cI4HS
8B1xRtQRlXNH6pH60ivbDe+7uji5gOsj6tFgF/eZd5k6NIc4YAYkFLSHQITO0Wf6H5smd3PA6MD4
W7EwE3/UZZp4yzNPK4OK4DZZjY8rocjat+9l6SomCchHhD/fFWbkF15F1AUvqvBJfmOly7xp2qUQ
YCcQC5cyta0qmfJ40GNDNULM1ix9AHK7MGZILz1bL+gBY6VBXBmstsHVG0PwTGDCCFy8l05M2e+K
6Asu20M9pGK/lDEYYOsLItqWzG/ctE7hF8ADmw0vfgbDSjy6XGN29+GkWy1ptoxPUuFw0/jb07S6
2yqUNtpQGR4WAiqDZ1484UMO5fOLsKb4LxdFZHPWmD7QtbfZ/6MlKT4hPcqPwqn39Ynah8DIqkLw
WJ36CChI6brsNbHoCWH/NcfypdmRIJIfWW+G5UFRl/biaK1IA3UK9DpxNC/PKq+XYI4JB4hu0hjf
A7ks6glhXv8BKAmUgr3rYhrojVvXnnKZ0cAM6F1v41yS5gLaCXNfTSPlDeX9zou1nKM03qaflNDQ
5NFxZ1E1s/savD0Bypu35rAni3v1VohfPRxHL+sOR8xRTtPiPqSTpnFX9ZA4dTTMYz8mdeRlbU1G
YJvxDeBJbivgqBH3czE/BAoz1FhqQ9n4QcOGY/bJwLmHQogW8LA2cWS3cOjHIkdGVGArsXpmnjCr
Wliwjt9EaRjjs6H4B8/0xcG84lVQI4dk0Fqi12Zk7uMxISPhBz2Y9WP9Min/wgIu3d3PXHvWkA4M
oCNFPUNuO68ctOvyi09fwd0tY/rj8oB2dtNuUv28xvpdZm1P6TneO2LHpmOW1elGSp3sitoTqcY9
VGVPjP1NDx+AbGmq/RoOaAHCuU1H6qAifcLAthaG566vJ6wgDeC0LcYDQqvMnMg3Xog9HNfCHtV4
++THqVz89JbmFavuC/JY7UfO5w2dTjt6rcb9FiLE7VF8yNGTSY1EJc7kh/ek2wMo/6sI3P+1rivP
Jpf9/oTnP7GXakcaERCdGEDeYj+lDpWsmhKWoPfXFaLc9wF9rRDRmuRCxgD93gpigFpVwQ7h3P1S
aC5KS/rOue8vSD/78uvTbRoTNEcyMpaJJkAhRms4Cq1Xk01P/ryUUk/WTwrmRUuSB0CA9Qihy19c
s90YVjtZAV1dhUYnjP1dfB4mFydFG/wQ/wQ9GqMgHaIcQk6lr24Gusg4TmCKPB2Q/FFxXPf+GSUp
6N0OzU9qdJvtQ/7sXCNOeLkP4Jt81WaTWcP7d+NHb5dYrcGFtwjEVvReG8s2EGQgvo+KIfYorgI5
aSDVMUtTwdfexY8xi94q96SfigXzKQUleuIUpl65B41XX4d6EYpePbU5+fhwM1/d0/oLXLRdNACr
sF9uRkcwZS7+oQVyDI+zWpM2o8RsZJCFaQJLFq4YIqHYDnb3Ek1iDQzPCFhb3qK3oESIS0Atn/81
ScIzU8r+S5SMjyAOSATmvzAJi+/aVYr4Vm6RSf2R498X1qSe3X985ZHuDjkk73+C3qxR0lgnpUH9
Qc4i7Kd1tNg2vSNQX5RJNps9ExuopYiauo+7YMw9zlCioffFubg2OnOtZqQaBTWEHvByA/nQCHxa
lOa5YGf9FRKpBc9Dff8IS6BOduAUjdUMycSyhvosnu1Qu6VsxuELTfqAIEXdKEtxBuZRcLqx9K8s
VkVr7HeXWFin/EJz67I2S7le53D9EnYRNJQpCwjkDHobhnd8cAKq0onw6z1ISSPBHFJqy/mo303Y
l+4tgxGERWPZ9CiT4fQfoI+raTLenSlPMBO4ZCJdUiyzGbhXQFOn9r20Iukl1CpFAe98eNWRqUVh
ECkU7HESThsb5d7rHMztD7JUXwFyGpx4C6HLBO6iCgxQEXoVQ+y5+9YgWuoPDh9eOXw56fJiR3oV
RwPZkgX1vVkr8jSxgAHu9gpuGrxnb4M0PwI5zbapi5Kr1GyiDrgRMklmQoSc0+5gGmCWixAFwa6I
rX864UbY9ot1WNGo6LKg0tnbGzY+6fgO+vONY7vpJjncEPzFhMRAahtaRXSE
`protect end_protected
