`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
Ni2NjBB81RMC9+95a8PdLXOVzPxNBB/PYZM3XG9aUK4kz6jV0s/Y1AfsjzdYJyJH0YXfUdPLnPSq
mEFCv4oQOnmbnxBYJ+MGPKsZudl2fZtbIlW37TEdYDMJtnI58jbBIXy9s3ODzRGnhgDchPu8FBO5
t657j/fUAclrtWBB5zjOEbHxhxZb2DDmpLLQPTGT0JH0YpVbx91Uz5F4rgllqpZqj1hedXjmgR1r
xFILEK+Ag9KC/wzojAyK7nJ+lXtNVDqW+6kE4337FoK9R2/Hn8h+4FR0eoiNg+cbZNq8FhldZo74
BnxZ21YymB2aSzND974NQw4uY+bul6n2XltEbA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="z3bZrWngS+Zh/Ya6ITXDtooqKa+DcPTeHlBsEnJpt2Q="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7488)
`protect data_block
hak+kDLSi0B4WR3uh8whcMdbikC9h6/rKc8OsIcEQLiAiIcPyU/aFwuzweFWDzvZrHP8qi8f7ggN
3oMQkiwHb7TKYIZEI/RvlDtG/BU1J5O7Hqs4TWi6kGPwtx1+r5cfMZBIfAmgqnF0zmtOthHKsDcn
bXb0epBE7y3FmFF53Q1UB4rU7gr8TtA4hRQ/Q8hSTGbdXGIsIMt3EE7lnp7vvEmkHsLfXWO94n0N
Y8JUvz9LcL3nklAOMrHu981E/kGZOo0e0l0ZlaH0H0UD2fSquZTKdjWBE6FXa2PzBwJZPBTZ5iNs
12uCPNAou8cmhxK7POqk5vIJEF6kC1DAHKkY++asest9Yx8+Y2SG4DOZe/0LzgWD/sxgKLEYrgAX
ntZ5gYEJw+FkhqqIxYdjtwCq5C0835JyhfrfegMgzx6sRR9AnaTib6V2IFJk07/QAweqH8pUNStU
1JPgNOTU/x6081dkhVejbKYpxqC12pDoGs+XyrxD9NsJrsPvk9Z7iSL/jZzhN23rmGnE8aU113Za
gMbTmp9jtzDUGEv1ASFFXS2xLD13fk/ObnpR1oWdRcwANPcP9PKgQvbTJoOvzxT6njpAj9+ouybI
UnPVfUg9KoGHDnwZr6g/Y5/rouQGsidoBPZUMwxaHV5Es5kGo6z7t2NapTx0vufnIb3Etiw/GUcq
6QBEsHw8WVkbwCDziuI67jqd/XpF46Ng+jDvwRUEG1+wG+AMkisdmrePK3vvCDy2kPGY3LvyDelG
iyx55YaFCuphlp+rRRNmanL7MgcJL9hZvgiMtcfYzW+YDBYhpTjO+KOT4tXKlQGLkCTyDh+rqu0d
AoDr5ifjv7PfJmagmaHNYlpIOB7g1Xen+nezNysZU3S3RuJVYDFSeOahWyzv9vHHFNprCQMIE73y
9wHV6ENtFq4GzeUGOQrHAfcQu5NSWvrVjAw8ycHsNjaXqntTk+dbUqgXZC5u9P/z3rPc3NfWAPxN
RfkHjiRrGAVxL9cbtc/vvDUtwi1MpcQhbtzIUY/TGsNb8XHvxZKO8+sTdQK2VbdAiK8YT8eEgIuw
sT2/y7FEqYphLV24DdMSwHwjuW5f/OB5yCFaQcF9SXjNpMlDIzmHoQMzXOFCUuCeMNwVPF62NeBz
KoGmFFARMeG7HjFh9doYSQCs+r2pnM1yaFVMao7yDOr1XX39cKxLudzE15shoDHt7cKbGO+pGC5F
iAT6wjhDnSOaUzLwZ884IpuFJLlEo0cIBwZH5qID+RrNoTGSK98AriwO6unYSZyysDapCFCpLvga
9zqxodeAvI6oAz+8JfdZZukDkW8AO2DSXqNtUTjOnQqoC8JQ39oFRlMED2IJvwggINNABwRun0Yk
ErIXV1F2RgHYDbU/jepJCYGd5eG/KJin5DQ9Zgt1rcyHzmuSE9DJjpYDBBJESOEqxLdMGQfu0FLS
qiq4LaEqyx/83D/dUmzq8PgTEEXKq+wO1y/tvPKIaDsE+bBES/a6pcjmEiG+S54vEI1woxOavdw+
J/D7yT3saryWAEfPrMY3Y/rfi9topLvHNQlMLtB0oxcr68IxiFy2mtqROgmzZbcVwN+F4ga+y6aq
0goOeYtOzY+xOPXn5Qx3f1EC2fSeqGaj5YRPcP1GGOVy/73fmGLE/JC644sE7vit1IGWHmzy/Ua7
EZUc67FJlsiFpTD6nms80XLEc0YBcO63YPqGOyjOjNTUI8YMp6L+mgnO7zN641+pSwEbbqNUXM4z
TMSMVHlUTLh3mL5d8XOiw6CnPX5Ut5j0LdUTiy4ptdbvH7P7nv4GyBOOGYMKhAJ4eCYeo+Rk1ywJ
N9qwC5RhgvaeMgjD8nc31jn3dIqBuJTpd3TITA6Wh2clNx5EzgJVJMIFPWKnnKl4LjzkSIIRvwjl
EqCZXteFgmST8o/BXqaLWvMJfA5c/vmWiuhESpZEYzV62jOjhlIQ1Fv73OvHPOutb9i2RRr2HlO0
f9ZBWfRJA45FNFC5JQhKC5hkdkhGavo91Y0jmi/fbdMi7eINOSIBTirhuxs0Lr8NEamfqllzWD4L
l49lIRQ7cpfBPNX0AoWglC/afJPenaRHk4SrDVafKVoD4NsWyfPRNCGJVvubglq8Ki+PKcHOOVaz
mP82gmRuQXWXyBciLXXK0wrl7tTi0zCMarV2ss/Z5wDWSnOyfnyQe1I11QYh/MX34E9svMA2i+rc
brDbduUEZHGLTyU+GrWhh66DRc4OW0o/MrACwA28SOsWxkCkQDFgigvfEDuVbmatFbiXilXS0bIQ
xgdK08s2Iae7gaaAg6i6TDO3lp0y3pwsaO0/iYOeg851NWpikLhGzSBKwCX3I2avHioLfPG+T5Z4
F4EfCEkh65ulE5TcBXGZt2752xEULCF7Ykqmv4xrgN8+hhhDQSXFiKmIWsZ7Df5MpMACzCF9SSsu
izc/tNRdDntOgIWTY8i7WPI2skYVknuAIap8tyoUxZ0/9ZluhaNrQ8BvE4RLqF99r0cfB9idnUBr
UU1/kVmgJkndMQ1UpW8GUgKyINd8Nt5lNImdjmzankA7U9LTfOZz1GM25DDy7wodouWpBfB+GPry
ewlgP4BIBNw9b1Fj2+fmM2erTKvRsLE0lH3JQyY9B6MR0BT0qWkhuIxJzHs1izF5Vr74I4qsM7vq
U0b3UluDeuLLPbvQC5JdwdrONDHSSnHxD43+HCoViTPAlhLvm0VIwefBlW3IpQtsxUjCwGo64OG6
94TOnLNFLrKlJvlfQvB1roMdlj6DYGucKnROlHvm0/wKS2bqUd0mxnY2caG0owzjhX1LnIAP2fVb
Epcbpdbi3pDyG6JGq8iOJP5KllTIzbX8hv2BXdaPmkmZy3Av3xKQpDWiQUBNAIPg3yAMooR56PtB
U8u0W1GMRapJ5AmzhqDiVnzVkbqI2Z2TkIovNtfsp8GPo1pQIqlTTvVInCB32tGXRu6FPL91VNSl
USBei+mqJnXGgvleSt/0DBSdQlMNcJ2n+yA+qaFCw/temFRGnqhIcOOzFzt/ZhNJpfdr9YSBic9s
UZ4Mdbez7BpiO/kbl3qRbaYSV1Rg9eTLy88ZqZNnURI4I6lgVlUyrpTvGdvt1x1y7rNOiWGAhuoc
bZhB6hJkUl+nuSrl+JeT8pRIyZiXu6ig9YfqfR2u7GWwSCc1XtdCkDPbvDkCRjqqMXGXoYe8h+L0
aIenIoFcj1kQkETMb/Dba9+6S3iJvMEpoGrgPbpnlzWDkxg1Q/Ct0O+0byPNM5QB2cJLQ2+vfzxv
0oRF3Aoi+VsDv+30Wvkp9CALMymUDIg+CH81hl2J7ilB4ZLGXdanrJZoVWPBprjZiiBHMJt44Vth
uv2Efrf9rAHMDaB7EHCIguXAguxUcYNPvjnz9R0Lx2/v9WekLMZROfW1FS8wk5+3CnlM3L9/MGAU
m88i4r+4OXmMg4l6G3MhI0wcKrnyxqD3/kByrLdLWKhW74HsxKn6BwwV0sDqp3OKM/fcVXPGbnP0
o5jDfHLKp6Z1N2F+H9skUAZ/aGmZq7rcL4n5DskE1LlvE1lHDTmbDIxGfIHXeuqqK6xyj4NKa4iU
Zz6mF4xp2shXlAOcaIa1OtUl90o8Y4AQTEMjRyHhDqgQDsEgloNiucEJFrVyictbXdlioT2zAT2E
uyNeSzQPdVtz4W7iYLMNe53JRwlXlwImnw4MCJUXX6iFMycf8ca01rwRbwNB//nP5SlmOEwdDPTE
301lIZ0JdKrrwcwVP9qrYDe65sBg6U84bOGVEOTW5VaZkynBxDzIRvJ9p+IZGDfDgHvSpz1Ldi1H
hWHwOEqXskFMidLg3h5sKtdii733avbD4obVac+gUKASiWUrun9Y4xbpASQcIb0mGLnEr/JccyMX
9nBdFbIHJZ77cM5QNmFxLLgknkeENH7GZBNepUaDYVAG4XcPQ52qthr/xuDh0++iLaMeYIYNX/D2
Awmn0Atz/37P7SoDvn7JIk4yE61NIgXaGgE/1/O6k7U6NS0NdldOIWmLQypQMc9kWXqGyr8uc/h+
s7BydEGKpdDwirydzDBPSOsyTqiSkOa5qBWoR3nADTunpzjgJt8OOW1EMGkPimbPUvttg92v6E3y
RKGU+Dt44eWigsQIgfTyAQTEPrA5s6q9Ys77mOLEYHHL3wpSXbWNPGR9sD/1V68rPzYlkQZy0bBX
cS3IrtH9iP8zEshtFGn5szpCAYWbQO2+FPp3L17YmPdUOwqIWJxi0fmt9tpEYCTAG00HUewBlHWL
obVJWQnFUPRxbivtdVBcf3WyZufL2Ub1CrJ8RGXEmLQwEmD72ZokIRBMwoDBS9B7Hq+1H06UpyTR
HBoYDYbFR3/EzNUoJKfIizauOV9KAxPc8rew44rQGZPuMOZTCkudz7xcx+pFimdb7uANmWjAHAQQ
RJNujSCKfzFhptOz/cZfCiVJMZUQnP4jDQ3RRDtJoTMzNjORzEoq51wxaZkzQxqR8rwdT2HgjGYZ
5psBdpPBT+bGV6MQThO4QWhUdU0ezdoFt5M52bOWFIT/wVz/11HIvJp4AoEiDUh2dnFOqT67U2fX
Qy2KT/iIUYR6Z8cAV1OLDBu/G+RAvxBUM9U9uYK60pbj+5BtbjjAbtIbM9TROKOiGrQROS5nXSaK
9bs1y9wvoI8qBKWuaZhtZBWWf42mbWLGveqhaob6t5tGSZYE7EMfK+gEYksZcA9KemYqPu7ZLt/E
Pdxv31VEd0YP3+c0SWWbQ6I6zp7YLOXWvm6DhBmkBNbrhiJUIUkkz614YGVCTCybMWvfTuUaSGzu
wdmylxSBPVn/pIrnEhLeFmuC1arfNInAx6h3lFFwpdh65vBq84UiVuvXp8nkKl3ItJ0c8I12kPzO
fy6Nh2t8QZMonXKAbXgGpWk3Je2uqdm6mPdPzuzyUk87JTOuir6uXJPipaTfIafIYu/D/gtVUmKl
QTzRe9bHfTVASA9giSKUv6v6LFppYVcpYo+VpJvEVPWQFT+4WNZYGVKqXMx8Ww1a+m8UEj1i0N7J
Y2lS0r4MPrY0k9EB96QW5V9WHtqNeNNssw9QgkdDABsdfL+lrEDp2PVkmJg65SKlQ+D//sFtyGjv
pQwib8AEygfbhs0Lm6jJPNVrmssNLvJ/vC9CAvg/Jlpx92GmhWfbhZRTcZMTZp6eHXKv9BAN1Jri
Rnlvw/fG1HqidRQLzgnHPdjJJXE78I+2t0tIS0qeI/l4h4axP97vBdOlHsydBcdnH41G7OePb8N6
2GN1mCsO6lPhfCPiUVAuDKk5tWhqtlnhd9BmXB/HChqXt0FsQk5zQsjMZrPMUs1JRJ3LU/Dea6Wm
UGfrbf1A703+GF+GmrLmVWurwO+gcTVYR4rXBJxh+WYgoB+ZfZxP4v7mxUCKWKeTPKCi8nHuA5iV
UKVKSIwMmwXgw6TcIm/NtcIog7e9KVrC76a1x298ygJMQ74p5NVkL7pgyjHGhVKnW/QOAQq6PE3o
tcQ3bilN2qmKRkvCre7KdCpSB8FSiNrB4mZ0ZDl5vf0aS1C6RJE3NtWyw1SoJVHT7/dzmvbZWErR
dvl2ep4/TzZpbqFbD1Kx5mq1zzs1nfqbHAU92iNYk3/uoi03I/DeZX8B/aUT2PMEYSmZAzwrnoE8
hWSMBknRFPwqjwyirWWlwEWJNWoWEv8wj+XoYzuw14cDa0mPDaezm1OpHmeSScV0dzJBGFqVkCG/
oV6+lQCAB1WpAA0nsjGOyWPA5xKYEOuW+b/9Rt/4vG1pws3gwhqIMUw5j2d4uFrTCdTXBlZy7JTL
nPHy74F147P27KywsmdFwybnijOkLlcrUg0EnxLTeKA3U/TfUc8LADjqcDXM8kcYQGGGXDHReCtH
9kwIU8Je3EZH6UDDldt665fa/93TccpBT7GHgZA+ecbmyFePtPQrgYP+cwPSuopUCWTOXgjiynlz
g8l+OUbp0gav2hkZ+FVSMK4ojKb3hA0JvtXwEfGmsM/bnlqHCc5SehiJbrlyVQHIKOpC4aov+Kf1
t2fK/wPY40j6IoCFaIwSZ7vnObZFgAw7beQe/pmbpRBBP8veVRp3rw7zdnW1ccPOXQViQbyLa9uc
s55gy/Q6CEvdggu4EvCs+fkIGC1EoTkgk/oNTUTDGZO46HjMYCwoIna9hd8a3ed9AK38heCxPJMt
fAihptgAW29nZ/tSVGsSP0OblLZcb4sYnJxE8vwm4q/PWzk6dBVHAe3zm4RvLMbu3meo4CScOtdo
zeufZa4mxBnliHKIKHdH/fjuLM4DVO9OYH3PIelFW738oT05sU8GLjUOymvbEU7DqaqFNBwRe8Tf
gBU40CzF+PAC8D5sQq3kCPsEHqDU+47eupKYOyOWpwVGcUM0QW2Q8alfdSZAcWHarMjrxiYPAzFu
6bJgdBkrTq4XyeaSlRQUlutr3R5SrK0yjEoMjMLdDRArEfhz+NCrlkLZHPhFzrnEe6BO68p/UE+b
3Ah4ASgUiAnEGZhyWediGGbAsqAPrKI5qSJDgF1O/kfxKjER7hGO+vy5pvvkeSNB7lLhwkv7EHdE
iC3ru0HuEswmXYlotNdsIZYwclFaS36x2YQIsBBNUeIAL61KYUoVevSUdlYSDShcr/Mo5ne5qwHy
pPMcz+NgWng1dBgSza5+ORfif3WkB7+2azNt41CKfVLCAfm1WnAjgU2H5F3bW5MTJ/J1ouPQB1Rs
K4+KplfIGKlPxSmxFfdM6MDFMl08ouQpVkyEuHrciGbaz47HTNOq/JjW98PbbdVkOjpOITzW8kO+
8U5Nu41rgLHQlMv0b09sAeRRuGlugnmKyyuDTgXyGJpUsct5vbGLzRB6Qci7ML/xqbG32KBowqnT
MLOp4/bociL1zWGIC7BOe6ZnErov5trv0lozGAZsnF60p7iXsqCrxpxOarzGc3/qFi5i09l2Zpyc
6H/iSBeZQuLFsOzvemlJlkP9SYt5bcS2MwpkkLaeCQ3Rg2Dm2bnbHQuehorblYAMJWIqYjMIDM4z
/MB5FeIiyO6J+xec+/FhcodWA1O63GjSL6mpOTp7CNX+ygkgfxrmsYmicFj3X3KlKxqbrbYmzgs0
chGHJM54NtMSTVd6ek5m/9C+23deN+T2pY6BhWvTyC7UWlXHgtSF0sx9XVdRfOOarRKP2nYnXPVh
0tnu+7+TAWWb6BlRzo7qiZMLsP2LbCNEfd5SPZN8pfIDlvVwso7MzN53s3Bs1MDUzAaFUUyfWZvn
4rNXarCSSS0vx9CGrkCtc91JqMk3TVYtKolw2CxvZ3ZWZ+uoi2bI1KaUFPTgO/4Ty/u+heINi+3K
q47CZIpA+YAKN7gZz7l89YGdXD84WZWwEKQxSwEVl+EirX+dtTpoP7igYUyf2F7HNbYu+3dsGCiV
2M21oArfAUMgbaLS4ExqQJDRf6mhH6SDb8xyTTtZfXQckE+Oe7ZUxK9wTBU/N8ceJ7qTPH/AKcy/
LJ4kTRWaS/Hthx5XfIduw6P/d9F5Vknp11mV9BqkK+wfxmvRFOjapaZAV9lN8pYzEJdVIfcwjtIn
yEGpphYOqp444eyaLraTLcPn9MwIk88pJS+aGqVfqBY0L3uE7hgaNLQomFNOEEjEbymHARfm1gKe
y/C3EQ4h01Uft37a2BMeV/L5DG7oyULDrWYGgTIwU+5+g+wxFA9kfShRI0SnwGeio8rmlmRWpvsB
a0lnxy5kwawQAZMu8cdXcVaaMXpjGDJ1HF2NW+iPcx7ll1T3CnwuuqrdpyDHmHao+7vbaK+5CTFd
OdHs2gUI7kewvtSQVmrKzcBzFAykSplRRCV1F102oEBTS+wQ615aXJbxONhHaL4M1z+L1cVTix15
zi3CvxAsa2mVB/LVemqX1jrxxAkDCRo2esjSXIOTpFQWkT3uIT5Ywg3QPybgPyIopOJmVDrfVItK
u6172Ykh17OQUDqlSQeadPfRbh2WY6sWQdaEzknnbwMAu4fhVomU+gd0JpxlytuXWUm1ORmgkYjN
k1PEkAHkxkfoRscDnEKpxHAU9sw7CoRqYVVjPLyKaf3kFulCAZ22i2heQXRyBAcZ8O9frgJsHruE
y8ZC/R8Cbf2nEjMRl/ChNlC9BMgEP4jUw9LCoP7gDo9M4XnLRA4SpeU9jjsZyBhh7+koyWXw6Wwn
4y+lwBV8Wmih+E7LO2PXMPei09IojucC4vDzsFHSyalBjHv8K+fB0dV/xr9DnSLAve6vNkQdBnZE
NJi1azvb3jZkd4yZ8nEmtC3anPSyLZGt+f9x7IfvvHv8fEUp+h5+FVTFJrjyxIZcObayXJ0KVIPC
EpZkkaVq5cBBXHwFQmiF/CrKIZKse1ZSMd4Wj9gXD/njSaD8mY9vj8CfbbMzAIBOFgVKuyckrXIr
2WiZa13jMlAmcpmusIMpzGJ0fvcB3oJP3doIKSeVFXvGrFg5mflY+D0Of730r4tPVSLJ8+arD/Bf
tMvDxIn23/iGsP7PbdhtVo1LFCy6A3V1d9sIohsjPfqhmIPtTFqsCMiMA8AKd3p4QKR/YOazr0Nj
F9owps3aDy2zrQjr8o8UkjHgWoEQDDQ4J5dUdxf5kSOgzfrPyEEBonDM0r8wNs+M9ZABpciWf02R
LaKhQp5pVPDuGKqV0/gjWt4Se/k4AT8OFcG+Vf8ZHIfC+FdFTJgV0PpFeLp7qgcji2GkkYTTIgG0
k+2iYa4NEuJW16xACWOdhDrdhyuPfVHk8BOy3TmcIfkBYMJjd0xHAvjqKyReu75oveuE8n1rrlHb
9VHO3UGDhO5DmLvG4uvQy0r8Ezj8cEeQs5bIA0dVWWUuDMxogt9kC884eo8J2ENdCObD69FjweiA
v6JUAvYrV+NDaMSWhHzLREp1m0mtkvmqLKyhW1ogdkvf20dBgdeDjCVRDcjHP8xd6HZWtslotOLm
NvfaU7/1cn3a38StGlvIVDw4n9uB1BpPdkrIaGeKB9MQQ2NSl8z0QiWnHLVOANrMBAWI7Ubdni2+
5vapDMS6GJhiGJ+iuc/UGldv5MotGUk7dIYygaaETU42NvpWkVo8MSGupeCcj5aQk/OgvdyU+MUF
Cnk+hwwmV/bNkaBJ5HYpS31Yzh+15CdUfaC9QtMLIhRH6v+J2vJ1qN70aryuLqJBOPqV3LlpFQTy
fpIO3/2NZA0R89PIVZGk/lK8nhYXxwxqa6QMbzruEoPx0A45WvZ7rcERSb5AioUNisxTrHcvjcyA
R2pePmqqi36MXQo/0AMRGH0lWGkZtygxmqXOvkcWB+JP0VTDo50OVbq9FN1279/G4M1mZNK4jYYe
UTL2F4lcH7gGwyf3EiNqjpfVFdkddz+fh5ASXsdgvVEvANNQq234sHx+x8c42eaQcVi0K4N7cQcp
rQls0ulFl4RFHXKpx503EgATX/ZzGW9uq7+a8rU92vwjmXza0NNLuzRbvXVoYvQBrz/9AqwEAImm
gHB8Pr2J7TCe6G9RJG2RGQcUteMD+mvNyo7MMOtc0VbP2xqp8HxO1mQN+772mEyzBQRqNKg4qE7W
ACQosXn44OEl+6Syx6T6xnWCaJXDKhvZ32M07mGSbKv3SMwwqrzU3/s8shTxfclyCxoZISx4Rpfd
a3FHQH1aVRbdqFq76qNGcF3/+NAhxokAdUq4VlHcXw43UaTuCOIi7Svp/wn0MV6se6Ea/ZM4RAMR
mM+PzjscdhZ3YvSGEARpFJizMVH+Zi3KCz7cYe9A164xCA1OJ3JqmLsE/aHAu64JkPepDAWwC0HN
P9nLJeXq1PvzFa1SmACUtu2+SxbEkzzfUoReobyjQjXzTaAhIaqRmYMcCJKHrdBWIEFkwutVYuPN
j1nAVgZU/djhyS1U1xLhwPJTXoDTYpAZcZIHn2FY2Jp2GBRMfqjkUrN9dCvEfpPz6TBzUG6x02ia
EgB8DjlGl/1DYoMLFI9auC18fYClSUNSLb7Q/nwWNL8mYSD+QiC4EZk5TRIgSbdN/nS8chvSm49R
rQGychOUOsvlLQ62VonM1rbk9PL9
`protect end_protected
