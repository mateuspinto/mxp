`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2160)
`protect data_block
lPN3wYXjNcIohU9zxOOHV0hBJ5DIIBcuSQD0W272IWUUTIvTVcE4IDSWQ2noueghRhBFC+o+HlwG
KYCZRyCk7AL/1NvjzlcpOEgiZZrVREZhEpPVtSmzmi4LWJfI0nAuDDWkAXvgUz6bNVI5c1yVR8SV
nwM4kx53IAqlL4x8XqXcyAyhnUH4uwaGOm1WmT4KdkR88f4/kj0c3FWa3rpGBiv/E7aohkRUHHLn
ZzOtUI1eD9781cjpzvyUqSaaUiI6iNtJA9iEfodA4cna7JokUyBbQFP6ifL/Cl4MACQMJAUR96UL
8ALBGAKkUN30cyt2s+b4erqmWmvFqBJF4pTyk7Ugjpe4G4xHsKIJTRAWA/kMrZQUPlznMPT6ftNg
W2ivX+Q0WhM/rTcOGAn+jzKEOrdLTCbM30V6NttqOgnyq3lUi5/XbGx6JK2esJY9vmARF6dSQf7H
eZlGxnf32nWPwWLWvm/2+aR6zfmqRe+eRgBbRc3Xd6TvNcEiRcdPtfU381zLh1pqhK41SIQCcijD
ZMu9RLA97q2DZuzcTiktc+8bc2WLJl9m8JUkCk9EiISBXcHb0od4JdkfQB/4F0hRKv4ZHiDt2qX2
rUXWiiHEu12Q4wzCyBPbOvP/BUa1JMY2xTHs0ODSND5Kexq9itnkJgvNccB0TBMffyvrPzQZ32WE
AufcC+UW87PbO/X5El738bu9R5ULyCzC+2amnzbNtpWRWf98CbWxjJmLBi54lio8ucUJR1yZbCv+
Ktca8cqkIa0kN+oMiNUMnuV2f+zpmqTR8GxnvOx/xhpXg3sZwNIIZxRO1tvT6VFv+8l9mLAmwsEr
MLP1EJG/FU/zH/cZbka0o+SFhAIaQhSo4NLm5h7GBpJ5Uvqr6u3/0KX4H1K6AExRjJTnSskD98MY
QqJFTGlOGb5s3hgEFXC38tN51eLy2ooglil2kg9x+hUrAMLcXI2QwGaUN4sLXn2pdIJNS66sd+1q
sRiwBVBVGD/Qf65x07kBB1iyBl7IqntqCn6Ru4K4yDTbpkCFnL4YY4LeDJpVuCPU2BpflLbLbgtP
a5Fozt5JN3uatwyH6OcC6tPPx/aFjsMwVLtAkd08f7sX2+rQTx21VsJHh0ThKK9unlz/Mz20XPKz
nupKk+Nv4T7JFF7jyFZPWDBkFJL856zeWTPgsczAHM0CV53PWf+6Ewtgdf6KsWc20r7f95w6Eq4E
PYC1eRSDpC42N6XGPHUdZ8kvu5NkF9XbGUWjAOrRxzYobm+HX1K0e15FVcNn7pC115YjxPn0Pomw
GFW7d7p3aQL8ElHXddCVTt4doCc0/gLVmhUc4FWwHbH7PUsvPa4TFKShnnbq+9JMDWiaxpbeDn5R
EmM2s4tRA9DE3D4Pycf6CoiiDXTbdWs5uKZmhULC7sbSP305ZBeOvrpPd8ZYskAqJWTKdRzQlp0P
xAPmguGQh9rhdNi3thwgLYirG9FBV08qQUTrqDP0YBJrgjlq5QMXECn15heMwfctv4xrcgkwR4Mo
lGzttmUUgZAhW4kmhdERGRBARgT87cmjX8OJRHaZ6MTEDONGVxyZe2RRvky6dYJKDQOosjDomqX2
jsPvFmbsOm2cK61zbjoXashJTdq02KEcjkBZj2ZKBh953gnibnwaITtGLKxgqajBto08OKcXo6rG
dph4TShxigEkRejBvlEwALuRjTxt81j2FgQKx6AehTFtLUh6wcReFetMsV/Eu2cP9ctmH1IO0VVx
Z4fah9dcEGnTmaEA3MEV+wbTbh/MudVMPiVgk1qk/mYrDspfki4FWwYFaI2RTJXLgpAPnq8jPTP3
2I0trdu7fz7U294FSSDS+EDsS9Nhngsv0Kd+pk3AzacUXbtfYQbNCbYAj+CQAd0bYxyBv4WwWQiX
IVgRO6R++V4u/WzNq/GqP92bUGdVQjAjwif5n6gkxINpvd0qD9RDwb7Oqn/0CORRD/oNGDr9TrqO
xG98xTywVuhgJTbnWYYPE8Orqnc2cpgK+4JtE42HIFgpiYQvXq3G3OWwI8ekkDJV7ri9eapzogcA
l7IjuMJKGsfLxpVSxbOQjIt7CCRcTIBMhm442nDgXC/SDEh5ABEgbIht2L8C9W2pPdfYvSazU28n
BoLg7WiIePUcSBQPyoiMD4WtnjdMrA52tQ7O4eVStmICPVtobhglpDKUgU6p6oFqgxFvjlm348+M
YXn089NP7MZM1pHzSFDLf31wIYah997Sz2e7Sc4bS3K3nQBvOj2p/PZocI2iVRh/KACo05eHkMiw
Ok9l8+vGygGpVpmxpg3JuFtSTuArggWdcepAmnSKkUjgp9w5j9LC1CCLpIca2DYI1AU4Sq+N9k6e
T7c6JHA3eY9m5mIGpamGWonzZCtx/H1ktlJYGG8vyAq4t88l64R3+gKQ3sGVwp5F62xt/UkyPPrg
L3e1+QSQh6ERhaW1xLceVoCCd8yed9M5EYXvcjujD8BrbSg8ElPudHK9iQOX7aKx+vguViUT+E7Y
uy4bby55rK8kFFei+Lc7cE9zyzQLmj22kqgusypyv+UsxdJuWIPFUhVv64NOVc9eNE2ge8sXeXHC
FUIeQcsv+Q7ZOWi4srHXhN3rOWviIDtiOKaX+lnZiGc3MP0Rmxaf4xsAYjQ6ilCrFMKyVl69lvFk
grtTvcKm9AiGbys2g9GlhDEzB4m04NjPUAHCx/qK6Fg5YnahflwEVKbncXVAaE4toZA1/Tmx5Dx/
aOJdfNbWD6HdTaDSZZ8dqjIwRUsueQXIl444eaXb+FPf5DiptEwgXs/zxvdAMMwIrHeDg+X2BnGG
XmR6ioXYvau1hdW7yk/HOmTXg5/fsNbhrp1ESo1hJHRXvfgs5vYmHxo4v58HbXwITrqh
`protect end_protected
