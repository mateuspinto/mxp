`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
UcokePcifKMqsWT3LgvAbA/Fe5vRGIKMl7JB0vP1TpLaiPiYs24abv5Kxsfu9z1sQEjvdH7Fgnf/
Q+HDQpeAEUjTHHL/g0n6Pt2Pie60Hsa/PjXRviDCnaE19zjd94d9EqE0sdGaG/YHd0wUrNsNFx9N
+71m+8DyC1mbLpvTnA95MjQA+ARykUxniqGY7BIrH9ZZjB5NV6ZurkWbR5ff80gSpUBeGIQb0kd0
bQm2BvILsah95jLYZCEju2MFR8qu40/w1Yg/zaoZJaJBpUJygGg03nkYbNEdi+dXlRXYCKt8UmHJ
P60O/LJ5mK+8Dun4UysPAkMCflvWZbOeJFPkHYkrklwxRbZXuKB6GabWPvNFz7x+sBr2EUL1aO0Q
y48aNCtl1uZ9DTpU3QyVEoO1LguFZlZoKg4m84mYeOpEXsD0aO2SMzKdrBuYeN+PgAdAIJwgk/ep
nDNUM5BKre7DoQkBShMq6qDwMgFpwUEdSN+/V8dNLG6rxAzvus9djEjHB5ezEHLWOhh/oNmG8o1C
gUWcTimENQFwhSBRHIu+nShGQE7nmY9M9PHlzj9s8Phl6B3iSjPDlPwPZOOAiqdU0kV8PS3WmLtL
Q4mdQyF+tJA9LfI7aNCMJNaXFxY7ww3/FAswuClB8I0KFSBpNp2gMp95dStuoB7T+McNnXNBfUSw
MLkhXbJpmtmYHuALv9+vwxO8Uu9fpF1rkYJFWr2wskfW2xmpAsM5MoRQxGZhFnFigQxXL/Sw5xOL
w2QU56ZGTjWIPaIeUXQKQEQG8cBAbj/7vV1FNXfhXw/5uDRgKt832YFotokgy81tWdg8/6Goq5s0
AUIDCn2J5Rg0R9GrisPtoD7gvGrLQ3oTLauGQ6sisP6bI/dRLWN8ew1PPmUf2PuNtujB22cbd5bt
bEhAa9RTqp4+hme8Z18IRV6ScmjxYT9HQz28bs70Kf7pvfeIm+QWDMai0TV9Ts34cjNT5p47PI47
MEQLB4opozf14FIpmx0OUBwCv0RAumMjOKUL6r9tfHCE0ukp/D9GtgNn+NOZOASQgEjJ0zDIoior
5Iku81rKChtzMnOkVPWm6+vwpxSfRPuVX2WyM0NkBgavg1APsR6jYlfgrkpY/OM8mrccqgz7aww6
WvVFVvCZvQhpLbKz/vFg2s78Uc3cuDHK+arxyCtDvBwGmMPwdNyssq9vtifzWWTqcxAwIC6v6Y4w
YnBy/exJQVqnSSyFPRHL0MKNZZFo1WzaOQDeEHd2b4/71dVm9yNyuNbdFtla/nmlIwizk0n3xxBh
+zWu2aFIGDRqg6n29e3DARQjxPsl4Jl4sb632vM0pcOaD0NnarJzMyjvzUczVJweJaLG15hG1L+u
rsq9F7AxPTGIm8czxPFIm0TP47XXBG0DzYA/qa3DksTgbfItl1yFJCKB/PO7Jh5/yJu5Ss0bUUJf
82cAKE8RlhgtjoO4UREcDkWAzRD+6Wv7aRigsa2ggcpWO0JvbNCwQ5ed7jGFB4A43gCQLrCHjt59
+zUNQxM/bXqE96pNhMLedRytSu1gJFPdqiPK+lk4i81IWSqYheUOADvWdy8IdLjmbXCFybi1o855
hLDuC/ei8SPVoue8LGZ1yXIFphkhcUbL48HP55MZS++Vpl02+Dss66hdo3cXMT59dXpacRBOVANc
Rcw7VusuWuUTSj6ZcoNeAqmS3ySX89TDqIjAfMbiJ6i5Y7Wl8++ySCTXdL09NZoNU6hIR6TC6E79
eL0kcUJO2AZ2PqmRUyXeJvVEvK9Ck3vPWpEjFnfAf5IBYk9clH+9fNL01sbEY4I+IEX88LMYReIU
m3RgYbzWA9sXobiIKynvj8Bd9A8zzd2SfhX8mxPhLFGpV+7QvVu3ABJSWjI6MyLiQss9XVXi9G8/
RYTjorMS/fJu8YkbtERJrdrE8n+NdbpPJO5QGN6SuxjuMekERS4n8BFglD3oFNlwFdJVKp2iqxB/
rx52vozZ3hEzTrft40a8m6b9y8/i685k0ezYDE8pH7DC7unBRWJp82Rnkrq0oIxUwcS/rocGibFf
Hnhn3YfZ5Gv6l8wWRxsORn4i1OJ7iAVewu+A96l3ahYtqzb6w71rbrqm8zDxWld+X9JKqqJ1Ks9h
TbVlbeBN8ohCKg6wJlOythCjA3qq8JXtWV+dHj9eajlGd5aoauJzCXxYqI0Wt0smWtaLA7wCeQ/y
W7sG1I/8JXtW7n3eDSBkrb8crQF986vGl6tNnZfLmw2CAdV6Vx5/s7dW2DE2KZ0mHjqeaL/NLem6
l3jQ9jQfekLNLX/8hB3cJBqkj+nUGwQXCDvkKGHgAeTmejWiuXQKr2c0F4HIAuvQqU8zyX5tx3wH
Hvwkvj3rdGLbjsOlwlUJ+uWEjTLBoVJHKoxtmN3fyestnVmYZN33CNlfaF/073IFPl/wpmhGXqfe
XHDjASkk+cMkdmh1ni3cliiRewrYsbrdnByVog532mXzluZNXsy9LLAe7kWVY4Zfwih+nKQ2g85a
yIlRLRkfbxFB1Uef55gnDU07lF02JbEhCGfxM0O2K02X1Y0nxS7vHUtK6q3lWkMGLVeZwI2Nmedm
oyjhnij3SECfiqb3X5poFAu6v/Uku547OHT5pgc60cjt/tDsThZ20w0t6fUWnkF3twsB5CRtO73o
25tO5C8yIZh5nXUBQTRkdpXuMUARR/sk7EoXIyme5tUv+gP2+RPhfT6Ytb0wijZUUmQa+zVc7YKe
FNyBbg4l+05mDwkOEvyZaztQB03ezXXrvEQnTai4uAi8HSB9MG8VsT+uruca0lySCp+sYikPx4FX
YBimqXR6+1sXoOIAE3f6V8pJ1F5CDJljxnFGlmWBB6iwYls0uE5DraRpIOiIV8UKcO/XiHsBpqSf
6vU9i2HdHgeIAoOUK3dCJ6UHoq7/OuM9n3vMrpcnN6ZMFdzAx2QnPkeRJErjCMSg6mrHUAN7pNSk
n8GDwUjA9sV711Z24k0cZWvpaagYydIVmLx809v9L92uMBNSI/40nzqed42p9iEgriM4vB/IkVpf
+d/ypk5y6Ly+XWfefoqQbh8QG0DLNRHlJBcQHtTNTyqJbXxPlUIiVOiE1gnYvhNm0L8A1DGpQqdo
Ylt995yWrI1adnxsJlDK/HFOsFUGSmbZumMibJOIsMpwqPZxdddb2NSFB8yrgxN29aMxzQ2KxBJB
gh8Tw+pn7kWpHm9lnLNX3chm3RDboZ+8nodz3BdOkHPQF17UPvhwfobzTAr2EAiP/yAWXPwr/hFT
zoZx1Gq/LtUA68e8VRoEG2+wPmwljkAGFFiKCubnvwbANgeCg8l75Px3GUeQ1/qqH0Swhvxxak40
HRMYtf2PFRFEoqIV8obNQCZUJRs3eC4Axt84Smn+lhie1LPX7DGWZ91LFZODc2f4TZoYT2huf7Of
chJi8AUDy5SiAlM4yqkfiskhzs3so1lxdG0J6tvfLd+dYSc4yO/p7rY0ZlHldpe0Y4O7FV5oI4V0
o4H8eOJIrTTZ4QhAK6Q6Q2EmhRvDjEwhQWAhpTGIkbM2iqw4J28KnytO91Djv38ulNEThrX4Vpa+
SEizzPzYV9gEjWMbPnbODdYmzH6yrmB7OmyMoSbC02XhGi9XNbS/+j5GP0jnmQXpA63xpbCGritk
iWqfRH3QOAvNMFUoy0pJjCeD8Q/sE0cbgBaGm8VatOruD6sssgEG2S/hr7DBVRPy3JGz2eFSVMMc
NB71Al4yStaQ1gAoyphjzyiqsZsH2PuF0S5SDrQ7djwoAV2WY0BLxQtrpOtjXwWw2dpG+C1Nyy2k
S2c4BLIbD9B04m2KlqyhlVFsS0W5yCGTwENVTuoMl7skST8VvD7DVHsHBqOocAXOohU819j1MsjL
d+3Hw3ht9pb7pjvZmkvkjSz4s6TUv0FEGw2YkZ0yUVxEyk5LTGIgyIGhbuKPbAroVhvrzs78rkWA
ewbMONhhBleGvplW97Uu/b42x3P36sqs5riV/vBGXkj9pUuUZYlu3IN2DTd3HthkRhATGtfxJflk
BW3kNAX9uc8+mx2+TQGJxMBhGTz/OxJb/vLDuhGvIyI6XxR5W8LgJf1aOrQz25GsFtj8ISHnxgpg
U9DWQoy2hdTdMgETW6INGGOeya161veg8hr/blsqLZRhT6FImn7HAygAiYYRxochd0DOSILJIAWg
vdFXcLg6aq3nhIAi2AWs5kGsHYRmLU8ue/iebC7WvsYtiF7UZhqqL0lyw7w1xiV0CzhouZCuJ6P2
L2ALE1YUf0XUv0MUTi2dbJfewFjuljoIDMIKkub1SIrEr74hxv37RKDVO2XshcOC5mTy2uL3WL0O
+fS/fBMKLJ/nrOHtWAx4Bml2OLaNJfLjUXyVllroMXx4GO9FOGzixS0YCGTgKRi95MQtwyopv2Bs
GM9HlxD+cmmNt/f9UAVASjqM8yXPpe3+cE+JlZIElAFD+6Z/QbuBHguYyU3wtwCXstroTarQxX4G
oNB3qb6/tg2Y6bXwRZzRp/8K7LlXOgb91C0U+Tm+sCWdh/OodRCNSH/JVxemmmT20EvcuZULnXc1
YSu5tj5ZPxtNOVWE01/vroYplQjijvWMW2dlnKqxh+x2tYYYaso4QrulFVZUrH4/4y5NMXZEM9iD
kBoviq+WItOuvNYE9lB9pJyz3/wsxAOQKdbBeSVbg/rMGDWy8sgvM5hcpIGC7FrhV7uKwJP2e3KI
oeo0Dp17XNWoJ3QbOhU0p3ddN31jMZwoAkmrHWJ2MoqcYDZZbLnXHAeJuxhuBm4UiYp3nuBlqHwd
tHubSmIXbKnmaZNUVs03i60R6RJWoDW9ZskwPzX1DRfmd3JPHUOBtFXVNpkIG+AnSJlGlbXOQkOm
6S3+EqxSBhExJe6BbU7h+cdrcTnv/j9oHkkA9sF8QZcNfku65N/0GuGlEIfJlTFlSHn/n6I4u2BG
E2E7HzBubkcuIYsmak/ezLdvG9lotHXUBWZ3fFQLQWOVdFjJyeBxsDTSsA135kGyC8VSXyNH53UN
+KwdQkqi+dwswKEVMg/iHoNOvzRWdpNdl0uEDTtz8fSVUUpUUV/36meI7lc3k2MKQIy9DPyOAnfe
VvoEIQBjTKPQWrQDpztUwfp2Imx2WBF7iXlPRolyIiuh0mu3N+2BU/YXUNXyhyBIrgF7UaiKiPU1
bBw7lMcchXyMgFdCSDQCa0JNF12N/jlkA6jU9DxRDmtLwB117xqHuNrnihae5/gDMwmRlMKr8fEo
u5r42nkeoNcCcxQEP+75dU9ZjvBehz2D7jykb+4KIkA+OVhHVdFUQCekcggWDitJmJfETktrG5DE
zDVynKXJ8iNJmaQU48jIP0FJTjOFOE7mOyX+xOyx13+YmZoFmH8CW15wbZLOsT396vDIOzbldIJK
p5gh3DnrsrLOShDaTYOxNWCVxthhf2BJ9+R02E72g7DomPew8vzVdYF9eSfWBvli5zKOlyCJgk3s
03S34wge841w9FVqcVn1olMvLWf8IfU+qVXGPSt68Bv1wDWK8yZrliY7VYaxpuPwPiJylWCXqsa/
rw7Mk8vD23T9QO/8wE8gGr5WiAEnoYPSSjhizHe7rYwu1OCOREwAAznTiKdGFL1p0/RfVWzcqBIb
Tm0zgkAhPAIKFv+scugoc90qecboErrwC5vvkhqjolAsyAk5amkiyuFTa4wPc6ltw47GeXpUPd8J
n2cY1B63caE6AHJpUIT4gBAQGRy3H8LqZjm3KyD2nNu5sO0XdCxCnz8QPoLhobL5C2GG7NqjTcf0
/X3im7WxE0J55StELOHUfrPpPsfKIL+8YxDI3Hg/E8dV3ygcYy98dREITQN5I9plsP94L6U2n+G5
F9R7p0lNqNLN+Nr4urTO2Zqcj+ns2rLWp/kdbGCy70kYJI43sH1lKPy3L2LcQBlFPDIf6qzuobD3
AEmmk4YUzzH9p+jYmjRC3HSf9Je7WeGZoJRYq/uj6Obed8FVZabs5ilVSEX7PYkm0JQfuFJymli4
5yniFyyXRyVDbnc4rFOQ4k7Uc9sKnQzLcNgG00EJEJIRf9ynnWOrv11nQ3eCqbiGqhOEU5U8ZWlG
I/l1BVBcMCTkiAvTj6NtbQT1bYp3TReXN0WaFhkDSnO6ZkMxvp77a748+SMwATeFA/SHRpenDcLU
Y0RuXDNlb7gFYRSP53zQNkf+o18rMCVDj/wOZln1NkzxeWjmUWBU+LmLvRGCZuIyzjumb+6zGr0N
TkpW7WtNQr+owjlecPIQp+/XBA7AUKH5JYb6zVQyBpowzYBnAoCpplGwG0nIkSOpp6wrxzPgA4cw
0nsiP5Pn/m3H9ccvMoOaBJGtwE7P5bbhXJecGaLF9GfhdfxKYWqWUYFY8ZQ7wRUcjX3JRn7pmDVK
aGH6NyOz379+k0Jok61qD1Di6F8HJnaQ3lKLP9sGcPWCs9DDizGUoW2yYgO26BnupKWgirtTT1ec
WCKuz+lKWGwXpAY+DLadglVkEorHwzR+o5EzGG0XvOuya1ZWnivxlIUeQx9ptoKB+9n7kIroU3wt
yfp7unxjNllin3GGKigh4DdC1r9ixHLKwjRQO6xqIEHDLjeNBDAJSaxka9NxL3jEpyH9hmKsVzva
8FFrqzdBWicX6+DMnCR5DsBqsHz4gLdgDy2uOKWIILJKQJiCSvR+0XapoX0VOOb3ysFB3Qe3Dlie
AzXt9p+i47S5EbBK0JedlDj3jESw0PlMSy+wFC7HiCZyLAGJEo7kzoMGpjdu4Fn7BI7sHczCWHPk
iwD7+lVAJibJ4J5dypzeMovm3+rK/neCU82rCcygYnx/bR/wEZdgMjbrUWxBRy7m92Nh6GU+i8HN
6cidYBd/ENWJT/4WkLNnQMka2f0GXTL/GYtOTC+RA/mDSe+Z4Ef/4x5VpZxJPmPF/tue8bpRgLfr
9GiKwFmU9A2ygjxBLaAAodOKrrE1BwQGU2esn0i1OcElAOt4TAwz3KxxIC/8XdsBLoEoJPH5mSDX
LbNN8NzaitxBffMwACECHhREtsB9vTuTcehRr5Tmq8hiFl8AhYaX+Ajkcw2fDNNsVFbCOoZcrUMb
5sHzOeqzb5w+w4+alIrU7dlLvdRUZq+kPwcdWznVaSHbQU0j4bhUtbFNkK3v430Q4HmaER2kkOQV
8hF7QrWa/UQ0C3t/iUpZ4OC3vydYzswAVGowRJODnn6zWbTlTcTndQAvQdBLApdCfKe4Ag84QHWH
qBMqpZ3toI2meti//VgEzl6+C2fRGapWuW6srMf4qwGlD9X70onOMdVfOEuQC29hmXes1ObuY9+q
RPut3BKOTRFyHPs5/kyqMPQFQ6ow+YBXFUftkNqecP9jHKimIY/X9VbkT3N90LYosJm6tkHZeWPj
PXjjXvZKSLNZx1+5X4dJe8mV/f9VJSj9fY86/KGWrgyFdgtaNOorAzQzoH34V3EITsAY+V6PyYtu
DmW/M6mfALpIoKYrDJ5BcjkypX0nvDvdi8lIbkq6RSm4LF8apoM0aEoI/bCYamzs+B7F3u2wYRmR
5ppaT0N2FQ2Ej95Bb+MN+DAwNfhuMhwfi0gIDgho/IJVYEqa+DXXlMZfVKHq/NmYHuy9KwzDw26C
pwb81JC5hL7dz1vRJV3+QA3NdXNjuEs1r/xwZ9jTG5q3aJdkzq+AQTUaMIYBh4xrC72y0HJkQ3vD
r6j9dnNmfbfjdkRIrjzdYMzusBfBdNTz5d30AXfLJd+GwCsCaibOMINi9XvjQKdWAO2IIuDcLUgw
0H7drDNRmNbwMRM/oUCS4QaIJTpZIZIKmLrJJwa705MLfnlYjd4lChnoeOdZmxSm5tn78NT0tyUV
ysCLgz6UaDK2RX+0qkwTbzOqhb0M8+kw29wuwHzgtyI4FS2hNM8XW5q2ew/FKCm66LhM11+fDYTT
GCPqEKDqhkLznaanyvrNrBha3Wdj8HqLlm+RtSgV2t7fssulEPabj7imfuT8uyyAs8rYUmniKsYl
S4z/4PtnzunzJn9VnOOqK9TEpuldRVKca+yAVHVoxkbjXnAZROh6wK2Rf8idTe1og8W4cQyJgCT0
4S2lF+jsLhPCPyU0eEMENBj1mgmEcaPXBl0e5rmbcJAB0abXX4MBq2OG3yUOBcDNu++eVlmDyfwU
WWGDMccsRqEqOItb2W0ENFMW0789IIYfvQYUBjRG9inKqBwTY4On6+AAhT8J1gvTCdCS9jXcSoor
mGitQhJH55jwsyYBPHZQ8xQykBCCMihBy3aZf/j1wtF4OF1cZatUQxMWfAvLsl85bdBJcvcTdMvH
p2cIswZqtjJWUfQ6QS7VA7IAPouCYe5sMldoqdzGORQXdoyUfVoIPpueL+DYTXJz1Cxafb7fzfxx
lAuuewXlYfPyGPywg16jUDOBt1Zs2NSq6r/AtlaUxR9mQyLq6QldrxTHeok1nZfxkx2PjZgTAO58
vk0Eavqgq5RNOoeCEGjQwtOBxFKVt6DGJ+X7CB7hfyXnygL3EzSMdlEPgxe7953KbPtgwgdIWXRB
MK3rFh8jxa0xrVODlNDKzw==
`protect end_protected
