`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10000)
`protect data_block
7SAtN/VybvroZ7iEaiKuryaoz0NRyhWCTit4L/P2ze8HEywECd9e8Lpbh22q2aVlEhuXdL/JVtup
hcXru4KRuAgGFmLyl8jvWJ5RhNW01puFku1t5/CjeHdW6VObBcQY0581Oeydkrdd6FEvMZaZfmdS
KIvWtOHxK1DA6+jzx88k8qUQJpBN9YLrnr+flE9JjBQ+Pxll+st10xI5t90Bys+LcOiFl+xMy5Xl
G7zTlqbiPbYLC1WaWKIxed2bBz2EEDfHNiIL8marQ2i7qEv5FqoFQYr2zX06nrD0G48qi2+ww7Sj
6pCeqRgTNn5PNjRQ0wYFHbFhe0v/1+pA74BoG+H/UIy6EVp/UdQR+YuHWL9+X6hIWjfdDjuV8oxq
ReNLFWILTj+yH/fASubasdWjrvlIU5wq4d4tNb/5+bz7KHKgVgVO3ff9Gvl32v6ZSSuMPg2MmgL8
2iooZCY+bAE+c07gW1SUsaRiC/NhmY9Br9IYzUan3fYld/L9D4m/vcpB/ghGI1C3zy+HygkKvmWw
v6kblloBZqLatIqXT76MA4WtyWWVX3Gmk9MboziZhTVQclVBLZedRNgewTr9yd2UIj81iA1jnp61
4Ji/7IgCVava230Ve1KhTSrBCvBO7lX+FQW5F+g3U3mNV6SvNyg/0qioaAPe9Lg5BhhGY2SLsVQ5
IHRA/ez0LoE3TQ5Mw3UmqYFQEbVEbXZ2f7W7mUmQb30WlTNUiMqcRalsp8SetmW/6u3Fwz+NwStE
TSEuHefuYbs3A3oQrNTJ+1PI7sCj7L5aXcWJopVx0T8RMPMNmgzm844WLusyJkV0N776c1zkvHnP
Zhsy+tK9A484hT25UxfkMZHuiDkP/7bbMBYqRZ02JDXVLfYHx8AvSieRQsELZJyuprXYwvkby3kl
xwLItYaSSH3W3OIIV4fhmDHPADbsw/M5j6CZAp7WQ5vRSMU8sINYyZGO8gQAdrbW0j6XAk48RbJG
ONiIFDMc/xohUvY7SkaAFxyrobPgk2YTWTTy6/2iBdTzE5X1tf+t+wr8qqHBXZBPRNTKeYwGLL3N
Vmdz4U7Q45fZq305rkF6jinOBa0qzqOz9y6aR4p8waCyP9xk/ZHX0/KlXEIEVa3gb9RPEO/hHXh2
1Q9L+9WvBd7l0HmZmBuDW5V8bRPDC4iQNQE4IZDSzPMJQ74kQwQJlpgWahQiOiytX5RTqMZuBKbb
lpocDdtpP6KzMi75P7KYpaoq7uBvHR7ksVZMCraEJxygW31Vtf+goNazTCQtMGqmDFz6/qihfhxL
9nd/hD+Ssb7Mw/jV9wgk7xDDzgferlhHvuJABjLPfkFfuKUy4QZrdGNbLP0tMMeZy8fGrYAp2hdd
IH/+t0SaOOdGZ+eUJP0MzCJkhM6IrMesEOMWusKY+1szEWODUuhX4E1LbfJL9U3Qdkw/5GxMjG4i
jXp7ypk1IuN9hLNj9eFdmKTWrUw6f+ifgqQq/8DydHUtjovsrSeNEch3eXruG3HapSd60Q+//hkH
fitokjQWnktCJX5ubsAi9kumP93WUUTeuuuICGmlD3/ObCQEerbe3KWF3cEomefzIPo8P/KNQlm5
iYRnpBrW98mgbSmcgcqFkJ67phj4P97EI7azTIG+aqjLTjEHV2raq+SCnVXONWMdM3OjhKdqMNJ2
OPySQn0bGWVZuevp/VFOhz+8Z1YqQOza91WoBOwObP7p+B+Ag6+a1QAuTGcauvs9VRcwh1AedFfE
2QCxgsQZJFPYlu/r5opNNPn1Ph11sUlv27Acf5bon+8oFETpKEJRD5p80S0DKpSobF33VfxnKXDq
KU+lmkr2XPHyHmubwP0U4V0+7pkNxOvLYCg92H5jNKF45qhyPI/19l8VkYGs3HyyQ8LIdBDD0s9o
T/v+yDUvorB8+xtoMRyAheu1MSuzOr6bTaqYE0jmeIsxIoB8ChlCHiP8lh+rJlRo4Wr9jSpV4tly
GK4RUVGiZrMuo/ART9x/SHYMhgo6JevDNoZBd3228TaK+bMwDp6PreXy090BMUSvjM85WzBUePnF
GY2gqC9U7NozK/tOwsJUfwdxkgrXcTItjlHnuj5j5NzAAi+N1a8VWsrlnKUeZNIUWrgUp00/VAVE
A7llWmpG2vHcxqu4o15R3kf9+qr9lp1U+YfTRY3+HeC/ivJ9Tc3bMUZ6RAltgMBO4cD52Q+bhaWV
ghLaKwCGrgyqAXy3b+1IAySVzxiPGIMUByJEzjLEm2HdQE4QtXkcw/Y8jVOzpEllkClbINu+7jIq
O1Fgg9KhdIYKVmQb0hPEg9aL/35ey+Z+CBAgGaJWOQLbUDFglhOh8BFTO+xzi/cyJY36xacg/6f+
Uw1zTHpx2mIFDx8i/oaGgJWHKZrubNLMFYbMhLl3c8BPXV1s0oTu5jbpHahYKsaoQDaI5x7wGqPs
VH8XoOxsBXuUxCAR4y2KtO32S9kM5SLQjbTXTCiQnCSONnaFVRdi50GGzuGtgP7D3uDZGfXC7Ggb
yU0kHC35yTXVzntRiPK2KyAitZWHiKbSV8tD+mJKCRMJJnf4YStpby1f128rPrxUgEE8jc0Z8sXg
ngnflCjYkErjNo49UeGAeR82UEpyFpV4zfYmEWkpLAapjCkzUV1tfUZGki4ihSB3m24mJS1nubb8
wO9N4N2QypHn8YYBd12eaiz1/V4jcuQ85qJ/IEc7e0GWsxjXfTgQr63OTnLNSA0sCAEGIzcZwYtu
cdhgjYtIee6tUSd/cO+RMpOJ3XOArUUc516o2y2DJFXVhMu9MGN4f1FPPJrcQklN/k9FCinDVcYS
hKeY8ywid02qXo0/JkDm4Z8HNEj9yp7mhOEhkA/EgYNHdYbhnuisuqfScLh1qiH33i4TFXACAU6A
cmlzz1WimGvKBqO+ic74HUfm45t5gqbgXWs5dWVr7TKJdd8S/kKKugEN8m3g4jvN26zJsLgOHP7P
aJqDyDh9UG4NOaJppwAQcz/wWdcSF7ExQqJ9vfy2VL/9QBHt8BXGDryzGgLcPG191h9GROLg50Cb
NZ+o3vnnmWck4c7C1u4sPo86UJy/LiNcJQpJrehohzReSmuJJUnRDH2D5hTHrfTrL41CwH0I7EkQ
iQvoujYlJNdd4fKYE+YJpoMFciB05yI1gvBAqx0BU7ExonVJVx1qgf4oIemakmG0iUOIIaW3qcN9
b5Ai75sYn7GdVnBDHgKfIsql/XpCt6Jo/Y/l/igY/ARffzmYNyMhELt2Lwvic+Snrbi3WjJIh1j8
vMm3zGlomnskIlaaW8zhUaFy5LTimG68BfZRn5dN9CEG//6nXpGnUBoCJHKZ8lPWoN3ZCJ0v6ft+
HoWMKV4180qzH1HxQl8gf2JgTQqBiEVzLeD4SxkHt3yhLR2Or2t6hSyOSIVzXksZ1QoG0iWeyTPK
NLWHPy4MgWs4vEjCskVkKiFnArbwCXbHc7+Ox9r7nrLFIgf/uHw6ko0+2B4hmoxSJ240Gya5r43z
Ih0/8CQD5ifHUPQfc0bxZnVLIi0PgA94L9HgfaqoEOPnsFLCKxq/iYxqTyCNGmvkRtGGSgUMDMjT
ubwfIh1z7co++bMn8qa8Tuy0AwBn9SmALFzsKexra1l6fZ6sK61sffILBsCBti1l8IuJax3yhPBG
q5M8h3NzH2PXm9P+OeRYR1A+rUqCPmtyBH0Cj8O4p9tGoJozc0ZPIfdWmlpVTLTgF0aT7tpt+DIi
CTASALaoSgIH5n1gctfTxR4ESgzNvKbkG8QfGtNKFuAPXxkQ1XtluRR+nZ0g6ZlRUMb43DRv+Z4q
FXJZKqywxKAJ81syoZ4uBqaFvQ+9FUYQqaFBK2+9SdYpRlJr2wBZlBQuftAacCGZL3mzEWmai33m
YCjuP+76Zbn7Sp/tnjvD2n0VcxdFggGsdiSrVBg2vB5QEIIeH2mETUx4TWP5GwFLnOVcwa35qU/q
ohMShw/qRj98TcOreh5LhCCY6WpNxX6db/QFj7GyQncw9hLGla5otq7e+SIZk/j55NI2rVCKB6d2
tP4GOOHZc/0xu/r6S4KxAUYLh6eq2/Ta/Ou3qxps4ZYBN6JIPzPyRKg4681tE0eysol+bjKydI4q
PQof5mXJLylP2VBo5fs8sNoUrQagnx0siT6XyXP0f279XY6tF16IuyrCA7RF02cJy0JIz84PWLrk
cu8me035ZOgpxr/BFC1G7TZr1v55ztp62NpXZinN6L0jWkvnQN39WU3zb3cUWZu0s9QpRYJW6zw7
U6XQA/acX9YCpq7Up6NC6FD/d7zCbVCa2L/XD+R0x5uGcqRK1zD+njiQzNLyKy7zBPAqVN7pOSav
Gko+9Qi2NC6/XdL1z3PVo/WLjqoxrU8kXHbujZjrKQ06TPTRq8WmYJfRD4/8KuW5+f7N0SaKAOPb
QI8yilfab7ivdISTjjuaMulJmkelaQkjKnmMD9bkZqAr6XKrEE84w3BaLhsHkL4ZO5I09nWN+Dyv
/qySBMEHCH/vAUd9XFXfNhEQCSGtkcj9H3uDym45jQelGqYSbf0O32EfAPGjHF0I77YbPKrUK25O
I1ChQPd7KiEO591L64D5A5jomFYkZJL9EkgP2Ty2aC78PwfmJJtE0IjdDsihV/oN/US9nx0+hjEM
PEa45d5skfL9BOPBj6NTpSf1AhPCPi3QmqJosmxTloT3EVpp45wE7vdXoeHuIzD9GLVgg12MKTP3
In9DhaH8v2+lQyfyxAmFtn716vrgU1EXFgqKuQEb8o5qHZpaEbDn/A33NkA349yakLgxkBF8ZdNJ
BLr/8sIQNFlHAcpNMXSJcwqJZYB5iqLgittDFs3G11BxhLTF/jMIRK93ptUGiA0HOcfnzUIkWUed
Ln3ri1b9iK9aDa7nD7Z+Wr3RK2T34N/0kkkSKbJeNRGOOyyEkmf1WH3fNcd1zE85STmlESLhntA9
4WLCdfA1DUPPyYu7UR3i6O4Oxsic7keAwC1WqhPfFm0eXe44TKw0RSA94cZ/xRtnb0KDYPTKX627
fhOSj0EyvovrVsYYlVtF7bHDjQS/g5Q5wg8n9w2N5iHWfu63m6fUd96fg6Wv65j/10W8KTHzvXp9
vSOXXf3EIigxPg/JmefwArApQ5NSVgF2zVyUmz7VefLOmQEiCf7Myyy8qpYJ73lcLlMiRoRZbYN4
lMN9c3KCGDLltrwd5zGPA7QHsoo47kOQYLXLUxZfwmu5C20oS8/rwWLOVI0l2r12zKsoztZLzg6d
4H9rcfy8Eo/jfSRn1bnN/TkSBSv3xf1bnd9fig5p/PTb3vUhjiLB2Ajt3fKSWrIbaFQd9SLeK8J3
YfdOTx9Bc1qwI8+qSG33Ude93cXNCZSkEHZTAkoJ6nVgN4KQI2WIRkMlzuF27W6BnFVn4NDs23+l
02ppF+JTDoEWwc1gaC53DQm4cC60zZq+SM45LqMTwYxbCH5aSVtBOlD4gUEQg+bafhBN7lvHstuy
HeKv/kAUkjqdOkx6EoDK1UH4+YUWK56JVWJ6D8oA5Ps7nKbKh47YKHyO5XG7iQx8n7xx+G1LOQp4
F+9W7QsIqu9E4g0d302tZ7Xcv40hdb6xygQ0XeF6ljy4R4Eedw578oBbng29aNOuGYGKHY6yuwiR
O2guPlFS9bB5dftJ7HDJmggvCEts61dwV0oMP5ORm9fI28cAGGDinSAPEG1c8nh1zq2rwiy/hQ/5
ns+veOVM32tD4uQpmbA+Sf6qJ0bpIud95VdTeIN0O92wXWvyJimRgkZsUsH+wWPH4mP0+TETsjtd
BmLyM809KrFzO0YD9elqdvzoo5eCe/1iEMZ0fqozqpQO0rILsuWLwiLpuMWLMaY3fGraJp+Pv36E
NYwOvXEWlQ99mkzO6YGqviyCiEyhQUHys0w68ho0o7w93FQuu23xn/SR4PmFpCoLDTMMqxLS8tyC
PDW6cgwo7Pfcx2rQv6ejaUAckAhOs7CYwLoGbjuLV7ZTWf9l2grdvUG62HGFzEgmzKptS/h8E04i
CwWe3AjVje/LFm4DbZCNXSkvs1lRyDZW+Gqmw9sEJAsBmIQlANgAag/DNEGaTEEUTc/XcjZNuP/7
8LXr+BZNPQF5ASCGTsebAk0qdDzfyY07EeSybCcDifj5FmjGLWDznAKMk4Ycr9LQeGG6ZK7Q8cQO
xzP8YGkBMpc3wlCmvPSZWARL2xlXYbHpITJXzU+qKgI2+fM3iHo7MVu2ffFh+CZEuEbfTP0Ast00
GgTRF2N+aBcx/bg6JBD6XaOD3TDgFUCuOsuxpOvx6ukS1jcjy/YXevIE3dC7rOpThoLcJeZuyJwS
reVV5s1hBogYbekvR2DQFAgLpqoe5Np9z1jGsu6H026Wevz7AdRbyTa4sAQ3ykeEOnDJbbz686Nx
dWp/OkdljvKDsSsQqEIklf329cHg0FH/D3q3fv+oEzh013n6dEuCWHfciJsYNICsx08vUYuMMF3o
DtPpSgkOK4kORtSisdb6npZk3PFfcvAq1aPfbVsZItewIRAwOZxrxPc3kExSH9GeQ33GzM00EXDs
YW1l16W1ZvWFvJztHk7kjp2AEbafJiWjSld5fKPTmtUcAGnZ9CzEqqz/yQ3sVmD6EUz5UZkvqegi
SPB7UhqKfBmsCMsxh6cNXY8fBVBpVOstx8YoKF5iY3nETkNWSb8hILzt56bmlD3E25MasLZCBRbX
FxPpxd1oVumQC0UbGeqSNsbJkBdvnXhdP9lpptxTx0JmQUHIDRt96VplXD7DUWDdgXRBkQ+4SP3j
4YqGWljrNBO1vATzotvyG7F5V1fA6qS7vAwkb5EdkqJP6MDwp4tHHRx1uiG6wq3KaZaAIKCTMoKV
Em7XXMymQe3NM9Q9NXY4aA0J3DeuWQrZ6BuD6aWlVYYoat/NR7e8Tz+zJXl4SRxCkego25zy/4Wn
ekFCfWDc7HBNEd51H1dDhQpVPtGvD5kZwQSatyVrNscF832Yrm4CichN4YGcvOhSFet8GBnPltvY
s7oq55uC8k4cXjH87UzxD5b/R4QrzeV+3BbjhNNaU61ADcYLG+mNBnWxPzy6yNqrvbpwKE9JkWWK
oqtmIHNvdfhPU79DzjRoLV2HHRgrgLcSfVrLEloUpcq2cSnai6aq6eKSynxvyY2u471XfdGqGSkn
9nrovn5ckVdgOsj/hA4urxMJvi8vy7n3LWHnB0kEsy07nwu1wlN60EekHyBEjXNCrCor7wZvtquB
OJzVuCgucBW5UzTcf1qmc+iXMoet1vICZG0nXgSV96JoWZvSLoGvHcqeFUfMNRxtk4+69lzYUYsW
RwjbyUJhDhWVtafVYjiVgdhjHKow6ytHVXzgoksRL0As9+BTHK+0pwDEO5zVpdG7A6UY5IZBrRzZ
3qDgE9nCsKAaM78KlteVlh7ni51dayu6i0UKfu1p88skRjIDwTldc+sXHD660MzGuqltFirdzifW
OGK7BH9akVo6hVcyLqigkgy10/2CqC1GFjfxkRwKYEd5Wr5Kw09nkEal33z00sSEFq5v0VdYsZdL
u4/FLfb6p0SKViKIsymSDHmkkGuAgqDZqOC1ALXG9VlATocXi/hfnkMO2sD405Wx4wwBwU3llbcN
A+tiQvYqXL5kH1adTqk0UDdUagWr8RYHBWbe5mIxWyzHMn9QV3+4tKmIJUFX+sura2ey8MWyVT1n
scqUFikQYzDYWzVQzAU7qQN0riZJNJUKAjCMS5JdNYZo0z601+DwTd8+tSluqb+j8M58RpbD1sZP
TXP5q1WXU/GA0b0FJFzUG8JvVaj+7/6pEupD1Voscq+dUbHOXRtvGyUs9itSgK9+1m3YtAku9Nel
Q8GacesjOTfgPcDpXQ/34NVYBijg7AIRtGvdkROvVgDIkuBuaBiFUCeyGR7oUOi3rQTOBEm7aNa0
SOJleK4iStOVVVOClhlnZmH8UFGcbwA6zX4wAPpzeRVAQ8RUNlo7p+iXtjaTk0i7pWNM/+OyzxbY
jSsUhtSVFKFz+zrPw2/U0epO4ZE7rkjEEXLTJGeEu8sI6DCmqeo41EUluKWqoeUxIBEoAE+XmzEU
e088nTVGsbALt1zbi6IYX2lLJV1pXmAjxt7ADKXLuqCeHvf+DH/4iWIyD3N79LJiDHOz821utmat
1ezV9rwdO0sMzQDl8LmeBmXan7y60C2rCeUS8m2BCMP6ykRQhJnX6r2TJW8wwh/pCtI3ZVNrrs29
/LDXSuXejHIGMWWU0K2OU4bkfGRfqB88M9ssn6h1jMTiR6VQ6f81LU4KTrat8S1LKOrQ+9TEJckN
UqbcyaWblsMdY9u4mraDnWoYvAJkJQh+dhyTaN+S+J69uaQgQz/hjN3v/P3j7LLabwP65ESxI90n
1FsAWBPECpTCY93D6DK+JeT1vIhe47dBIt2UdMQA0WUJQXhQlwkGuS4nVdYbZsMcDWN51Cb8aOs1
Sqj4yXR2jKU94szwdDhCkZVBaPPAhLA1J8KbiqnfcuwKTZAsDcGzAOdxBH+Ch1AOlcJQbzPf8J+x
kEi0sOimcDDJxK/aRTchKOh9O9wj9xqCq/jyYgAlR/EyA8AourXElPssytbCY6Wm+FhnXe8tsss3
PSL9VGVJZtfzShEit/hl8xX/mfam8A+LUSD+huPH/GkCak+85BkwcSeCv5bVk3v5cZPxN9huTRoh
4cWKEngAEf1+GZWoOIoXrh1XPQRmEDjZphIaDWwoZgAAB2Dm/ufCubATIm2orUB+3j3fau0gnemo
dArHiIrP6aASXcCfJy20VPK7E/wTzGtV9L+Q/+07i40B/Fwa1KdMeQ2LXmyDsEuwIJ/qAJGUygY/
lvnZzV0b4T9FYxMfvYOuPOpzvZuFGN6D9t74pn1kZpMsImyae7jESNEoRrnYCZm4a5QwBa9Rvjyv
pWrXORQGwtxahBnH7gQtswmZMRm3bffU5dCDVxc7mprO8AII16TKH6OJF2+dMBFE+ja7U1MRBFai
LESPZK7R1ZvnVg00FzdQpRDZ+YEJZ0SJ/rjPIRPuzHRm47G5Zi6MvReMNsdpe+U2wE3ZgCZaQM6E
F+60gDGoBAmd19F1tn53Jhh4CDJvHa1KSqkSDbrC8ll2txICb1Ix1ZueylyyAR8QOrTg56lAepF0
OUxaDc6pl68/Y2CtxoE6rllswSS/9oFeP2vn4avbJ3NPeNxs7IfrieBh83l14qcnypyGe2qrSjNP
e6nsnd+A1onremBe3Nwl0uONevGwBBGBx8yCkBryot2op4gdSvAVBaoWRUJnF/EsRIsJTG/Y930i
4CFGAXKl/MSzQpATJ1KsECcTb2z6wuCifHheJWF5U38UOLbOWmLcrgLuVJYxvVr8hn6i6dSFxsBB
zJm355kupqPFKPsOhp8T7MXNYEwMw8kO9NxRTMQ9I2I43WJfB8/+MaQKV0Eh63XzTj0kxiQ2+Rzc
wWfS28ypIhtuARgqsigJUUG5H3VB0IhdRF931j6ocYT3fdpahmObtcJQ7SzEHI64lVSPULImaVQI
+SQtZStTd7uGK4QzHfBqRrtKQ3kaeisKTLknapbD/8oGp24YlRlQVoSkyDlLYK8F9KAJH5MEOCY6
3mYb2cUDpYoeFJ1pXWkrEqjAARCXf6AX5xfDLrePstLAkF0R/2Z2I8oM+rzPwLCf/bMCy82PlJOT
aKmAhsYb+XEzY+0oLbsQAEqczcguqyQRui1OjSmlTXtL4csmBej/XuIAX1Z+Zdu8mpeG2/iYnUvt
RUzwgAYwg9Y4D+vXYOWlISGah/o2Zp9sG02OOyJZFK4U3ZUuABJy6IGB1a7oOgXIHJ56BoWbePfv
U4Amy7aIJ3/HgFHbhIaCl1EL4lFFHTWExPHDnkAd1aEQIlZDLe9amOD98GTya+EC2xexsMeq/wRR
W7mBrCqVa5XPGg7vhvZWvaXVAcoNKcTkQ/u18lwND4D1EnhG+anyUMwRcuFs6AoLZD71iiOmHdss
8Uh/TsE71T6GXcgRvl9JANyMIt70XVRul5Owuy8ylt2u98KlESRLHSjNoHKN+wVX4alxz7KQP6Ka
0b7oNm/fuFEsY+U7Akebh04oVr5GRrMWOR5iwRadfnA8ZyefBai69gSDt/b89SqUD9n/ksL3JmEJ
/0Ah98Hh38ZBS+lkf0jhGXr7Q94Xa/qUPCta+HOPdoK1slgufakztaAzbnsIO0nofE2t95ErpznB
XLR9/Tzakc464UFrWWB43JRfxLaHRNYXxlMa8jq//CG4ZPWX4+oUgUVNlHjheGdKIInSHnT7JKzz
X+RkGg9tgNvHeFrv/o4o8IhCceZF0gueh+K0nOfx8D1mi49PkE9vBWAh1QycE3ZbYfx9uxVzJWIk
bcfDLDqVjbmVSCiE1i8bJlb/1yOFWAZs8GnzP9CWwzz0qZ30mGbEb0AyjpnsenJJK24GoPwtB3/O
8oqJSyBEtXvWu+4Q7JrGFon5SGCIRyn51/uR74ux4UvqanBFMaeJAtKyrHS/6tI8XcTip2cOnLJE
zyasHVjnaaOpf1/JrK7FQrkHq3FmDlXrEnE9FGk0JgZsczoDL7P6H41H1xDpLuobzc3+PPyb2v5A
uq+SY5VUUlaMW3TSNx8KJxnLMLIZyavLFJUEkJ47x3SNnkBfV4kb3MrkSKTX/4b5VDPlhGMG+OLO
2ppd/Qy+CA9aRMaUOhf10kG/4Qz+48uOt39DUv6HQba+KqjO2XF+UlRH8dbSJVzrR/oka505UaFq
5FE7N+5z9vRs5d3wf0ZGTBtNyMtxjvuy3gHPCWJvUvEgU1n1Rrpmb33kChlR8AkHDJic6zfo8Qpe
FyUdkHLF3XMscE1i4ag81ciRJthY2DQinGXnkV/i5TAsTWLMXRbc9Y3bN9aBxjIM17yavt9fpncu
uUb0akd+vULNzheZl32V75gYz7cRNuYggdEyDjoAzU/aI69GezBqr8tm41uT2DcCyGX7G1x6R096
I/6u4jrXaA9QvgroVfrxq9VDdqztN1hY/RUeozIWZ23XgTx8TVfbr2/btiS4fRMscurA0jg9AQHz
NSwgPRaGpVvG0w8To89JDZLDYzjbnfOmM4OWdJoawHO7w9jI+zmJcuXzdX2ynKjmxQSHBeo2Qmb5
XEa2FlaihIDu79JGz5thWhrpX+k9hvbws4fqOHtq6gft744ECvMdw/8m8h/xuNMCrv/u4mwiFhLz
NsAMGD5hr077SY9yrDbuwCBjJ/3/L/2PHo5HZAKm2sQLs4JCmaJU+QbqSg3kzBV9FW6tJMMWZLF6
D+F4bDIfEljkVAgzlnd+PBcUUma3vqV48IUjsm84+mDsjQaxKiplTaLFQ/+gENZuT9XXDpA5wcot
LYEKVL67mS2yhbTlFhPVrrSPbxish2pq3EWNijR1ECUy8SLvkWKs097A8Ce7GPWZwB5OqZiroJGH
hqjt9wU0RvuGwxcbMfhlMZq5zAHYSwT3u7085kbYhHDclz07MV93+vX3z4nKSlGSuDFt7sVBjmkY
fwzbk0XlcB8EpCA58v9zn9thNoY+H53SRZ+KsEsuan+92dGRvzOVd0U88Uk7sH4w8tMTaQfgpK8f
d5RERhsDEVVxMBzCyBIMY7QUozuJptlIbm2jXfynnyYsAyk8unBZ1LHYxrPyemyAEVxw7k7V+/Uf
iwQrXj+j0hB3h7Q1DYoG13XOcyFT+kSAy8j77jOhnxzL8aMXA/o2rqi1jp3+eotOl9zI5anDzSS/
kXG2PMvWewl0r29yc0b+1j7E77AoBKeezZkCE+RsMFtAJNAGfpgzm9nF+HkQN6FDuT8NzgQFDpnA
lOWshJkSKKXdAydYS0hk64zsq+g5E/a7w9KHQRytFWbzt4V1GdQ7KiQdnHDrE+g/Yhqg+ICxY1U0
PgcBmTeuWUQUI36SUB32TC0JN4q3sUJ8G7BdyyT9RJJHELC4cDLP2Yf72TCjG6dmv7zhU2l8oG3/
6uLHygsHYTfYRANkHSvBlIxgaGtk0sUPv4JgKf/Ysq65DvcS/l9fA2C1iNFrNvFtp5YfXsMBWdyb
e8eWIAwPXizAKdBVS7ji1fOaKF4YLCYk4qA4b8UR6Zsg5V4lPR+KgS7/851gSJY5xk6pNYhafLn4
s9XmS5fAg89kK9lzx3hdFSHZpNgO8vZYULpnc6asHi7rFn0kXIUBRG/WHd15V25MT0jvH83Nnqqp
H7BZZgXvkZQ8HB554gg/jHLXHxp0Eyt057zFg0hepsgLVn9A4xBk4dF8x7xCVLtIbf0OHl3EiQbK
UqO2/TALAgXYfmfz6ghUJijoGJRC6S16v7JvjLFmI6EXpAbnPbVKCCA3pIdXiQGiCrCH8HHjf3ry
GYCwlofl+LMZK0u0lZc1clnvjiKci5yXYKpRQDTcz8lnMR8MzlH3xZAwiLa3NasfMyeCTdwZIcuf
cHNSM6TcQo42ElpiCTNq9Lxl/WbD4TWbfs+sN4RRH+x/LHpKLh0FAriyMR2te+JRALbfpVi+Wm2v
I/VUoQAPYCG/q2pzjcxaRHvOXdFRvA7loWgb02/qScVDA9yd8kWQcnROF4tG8o6pAdFgrd+2kFbn
FBoF8mqQI8m2AtIB+p9ebeupYfuoTlEcvTRvHA4B5F8DRbWSPc4eNvZ/OLU3x7dPaYA/9bav+nww
EqY+V1vfHwmizB9fVn2OhoK3uicyqNtUWwMm3ZBgDm/Wy+H3FnvPFzmSOsw+8nIWFPRhp0Dn6azb
uESLAddAXmIiF1CD9rjg1aAINaTGSsmgr5p2Xsk8Df4ARiQFEfJ+0xJVsMg7j3v9xXKZfrRzIWbt
ApFhZ9uPOUDLhdAiTtLL0x8H0biHktad4AbeIHHAiDWwOjUK5kpUrH//NbC4o4ehGuXGLTkWxReK
PTdCRUJotXuSH1AuFCq0DbA7HM90hiCGi6LmQMq0q/aIYsVeRRgBVfeRKrqR0bdNFUeoOgF6Frvu
OYAx3/C+o/t20uHDE/15pFUIyphJryv/W9nEhwDOMcz1SJtc/1xXLWabj9MMBFKatFf6enfjQzVV
BrHejTVZGr75DDrlEgVVl9h4WOxqSugNHL/jXd/VwyFMDQq20P3iKmAAY+d+T4Yi2wmrVPEfozlw
z0WLFT9/gdY6ZzMKWqwNReQnLq0a6TrA7XrZurOmOGfN4K0w9E4rgI07SbQrEZ7dMHE6RZhXn5J+
Wendm3M6agM8/lTIbK+E7TieSBxDlaByk+mcBOnRS8HybKjy0rd4NtFjI9Z/7HFtFBkybHI5/FHo
fTU6huRKqypwbBzWNlMiiaPymXOnUqmnvgYlVyRNIv4whbJKEfLHHe33B3F6GU4Nh6++5NGMHW8a
SB9SZgsTShyQui1ZOrEjV7QHvMdhgS0XFA==
`protect end_protected
