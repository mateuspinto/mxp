`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12016)
`protect data_block
gaTzVQ6Er1VGPzFG9DDnr+sZgf8yrNtY116qUZkW5gDb8YOXV0zbZAiRWquAQRJh0MUpFdRzqM9E
1fs08m97HRgnlcP6qL2Pe583qZmWn0bKg9sb9ZNT6BIYkLsayqQ1VRmzQLlBf6xURrCt01Seb7oU
ZvV8y6qIzXLQrjGQGH+zg45LgR9KkRFXTWTabEErkPOrbGcYuBst68htyRGlDLO5DWfj5RehLYFj
4GT6kZbNo1J3RfcvPTqb0x8d9bG4VblwpW8p1u+DBMc0GgGZHYyakNs2T0pkqBlOLotaavM7Wfiu
j2ieVp7biBPAnC0vPHAjD3bPPhwHhs7DCslRLl0VW9F7r7+nZQpAjkn2b7Xj34Q+PVqEtLQyytI0
tjk4GE0qBSp3SJUmfUs60bCv6HxN8Onp1+okf45ZRebGAl0G2KFw0PzhQr/VMICUmrcAc3KNdN4s
VNVFbBQvhGNKmZZ0YSS+p7vRYTkL0pzLJmvLXRbaxyMsDWdv/XiyAjttlIq2P8+1LBtkH0PvMCoP
o2dRMLwkIfJYqY8B+6jeWNSTAiroRB2ZcFiP86/wLPIHSi6RmQ0lGWcwEYdo6EOqcBhfFZRARMv5
kSY/TcZ22YjTjHxQesm17tM6lmfqNvX6KQNUlG+vVCNG2hZv04cyX7aY+EWViIcORuToYmvuHlFl
9yKVWp9Um1bngXeQcrtdQqXwq4wSzdPJRqEuqHz39RtawdYdZlwshvD9SybsBepToQsT+wS5tyA3
B0kdGQSUQp63sx6RlcvyRQvOQ9EPT/uK+wo0HogV3im09XoL4muFyMhV9gr+2+6gbadWyjqD5h1f
pZXV4Y0EfWhQFzAdE5n6iPvA+tKxh4n8GewaAYM+uc5Zebadnvg/oTj/xjpwG58iGrgJI+zghwWi
kTLVwVHU025i7QM74a/pDXqbJnTm0w5XIKWVf2wVA1p2QjpDWd4b/vQaGFbz7Wq2Cx2Ne8I3azzB
mK7mB9JMzoTZHcaiXhQrpFtzouW5j9Ln6RYnNf9dp6qKk+0TKGMw5eXUtZvv1Cbwo9VrZ4MnWS9F
CgVCGeWnuDQ1V3ML22CTFsxywpK80PJCL/C5BWZV9bUcFvdE6Km4h/gBxs7UJxXP9j85vefL1hKU
JDkqHw15UzRLaUDDheRYv8sqsD58lByCpKkDqx4uaikMcjCJ4LghBlAG3aGxJFaypnIrra/iRYgv
tGxZoBBOMCUZiZZ30MppfeUTYMje9b9UOMoZ9U4XxD42LL7S2PAUK2wDfvr/Hbqstvnag1WxINSw
S6l/6k5SPQJiEh+iIr7FNlGmmc3lSA2v4JDqkGHycNEgaNQGPIo494DzBm4YyNMQyeHKD4rtUBaR
9ALHJOCwM9UmF9dAJr4IH9KhFxYYkfo/eE6BaFQqjFTR0MfG9pVbri9fas1qXWvnZRwsCukal6nK
uFqSn5y0N5Ayw2p7dIi6BPXYRlXqlo8EN8X3mjHZzeOuboZPYdFoQCqgP2ruHYYRNRWwIFHsumEP
Qtaj7wBDDzFKWF2qR+X/urtw0Imj8NKpjWxpTFWvq56beIwpW0tiUS7ZJJ4bkX904H8Ew1vuJyeX
OegUCDzsYnzJP00F8tX5i1lOJFQI07sCP5j+XL4eS/UiM3ICyWOdi77+DPo/ofe7t9VfBcOxx+da
rcysYllmxxHhhZWg3wLtNtAebXiS/D7jwukFnEbCuRDJtesk1ch2/+SthsYU812fv04rgaUjlUrT
pA9u1z2YVWr75c3Sd1R9q4IImHxxKGLBNgiYqtHH40w5XbEn3XnaWHXd+gAaD9UsI8APSQZQTmZy
yqOn8i9mMbWdxGvP7Eb0tSH2SqO/aiUydMgdbICU1uRCfCnCioQjoVTBgLlIlWmgr2aN+i8HGuwB
KopdsncqTaDCs/WS2GVV0S3UthRGAcRCQb9R0dBYXNk7Bf3yV7OsKHtzZaAUZgjWGkzgOtblBHq8
FPWKXsYj54kPKX7esJj1tX/viI1B2RZ+Vi6Lsy20J1yP/GDT9OVf07mYbxkhPsKqj1ZnvepChRlq
YX7b8vT6Spk7uVH9AkU6f0S9QYPauhekr5fkpSCAxgbUKe/PSjen8FFqoGOiVNxc+UyaX7w32GA6
7UHqbYl8IP7eYEZYr9q9vVdIjmh+DnMgpJYN5260iqqm5QfdHEoaNCcaKQ/d9zJQUH05MaVl0ZO3
GHq0m2MR70gnU1QZvgs/pPoTXtC4Qjg3FHtRqZjFt8McuZqEAVBtvQxpkHVlQeD+vOyu7vJmyCjj
ZnIWhjuOYUybV0h6Kfl3EkSs/HbXkfpk5oAPEVe+PPyol/V+72/rRItxACdTs1wOSEgFEqfFh6VY
PCHnSRaOS3XHgJFbe7njhyfMQd+meabQBHDtKga8Ku1PgAnFZwfJSkTsc2oUHow5DpG8CyEQMqzv
gWPdWQA+L1hCMJ5pUigYfIzI3mpF7WPx+pHCRsDMaOsn1GXvcCu0BiFOyhmziTC03lHJA9IJydq9
PI9C1qKFog3JZAlWAqs40pJsW5EQQiksGeF2SSkqhrrIEbcONhN+gGG0shOJt0kUM+VMXhomrIDG
tcYcRzOk7lKCfDq7XaF27rf+G8ERwfrTZ+cv2wSTzojNOogvy1Vghlye6fe0SPdEiMom87syvTfS
78LrP4s4UNVEtJoXVA/az89yU0+GNX4PCAC+q1RlocSaQC0B705mwVbtnKCpj53lx3qof9VcN6Dz
d3iB+dX2cvnHRMTxn1eh6jeZxbAnWnteEn740tvWM934mr3O+h2GdG7A5+MU8K1rVJUkKKMKPpQD
8oq7jRem5v6xUV4maPJM4nzfa+n46zWDSbeV2ZZbdLjcXYQdnLuu+CTcnPZAKDCusnZJNMCAjYK8
WWhzme3ht6WFKoJQJmIWtFD6bVldi8kml/51OeVMgjmkldQuH4/4M8qiATVtkieHcUuopI8VP5Cw
/XHQNtSA3DnY2sceMn6zBPgUo6LJNLHStrfrRps/E/yq1/XvGgIlS/rPppC7R66GrTuLddhPzXsz
29espWXjygbl9eWgeXL8+D5XRC5UG5kzH0mDW3COp861iDxWY36ntu1t/7xXsR609RTPv5TRmKbr
pgdoRktyRD9ptDW/jRt48jX4Jb4Mjlc0+WtRxEcg9R6rH499ZnAC13W0q3KwmNfp3P2JUn+3k55b
VHGuMOSK0E3I4NdCzsgAy7sDr7yGvX0GwIL8PWTBHaz7Wuv9xOO7NS6/Jw6dShxX7ue1nKr0gHeR
pwFk0RqxFIVyfYCEZOaV3ZqPq7UABwOt6lze/EuFHQ2oiGPJL1laU3T5xYvzeb/1GpboGCjGZ3cg
dC6pZrmeXETW7fE9CIQIVTTlNb3xW9BPZaD3nzOS1q+b4qQlOIKf1JwC+V6iI5aCZIt29a17GmGD
T6F2/2BFrEyr8P22Z1kdV6g//MZmap++fGtUA1rYLjXI0UJ+mDuc9geee+Gi5cY6qC1scOV4COzG
qHUQdbCeOMzUpbs/nde6qJJYtWg7k0iNsXo8EBFnZMX3Liwz2Fi8ws5TpCcFli3sc1p41mgK6P0E
fCSiiRdSinUtT0CaVLOvyEMBYHV87l3gb94y1IuuVkO/9BnLIuK9rh0sPAG5sOZmpAU3+veGBu2p
OGH6sQfJnY5+fGz9WXVCBSbWiIB0Q7Q5KCgaXQpTYRi6CrNifLHcV5FjZ1A2oNxWPovY+2SfnFIt
aM973JyukdykBxWADyuiwO3cH2JqHxrZwfsfSaqLp1VqNtmJoDUBj/AtGAwRdPKo/4XaV4ZWzLCr
KauhbeA4+5JA4H8heWzbS18LH/TNhK+Yw9n/OV0tMAptfK76Bq2niirLm9f4KVDLsN8RJzJr35cV
3qEPg71uTOKH2+ngBMfwlwh461iKbz9PCQmj76acqaAUQBcowzorYqL4d5zPDTeZazpF+who0NUn
09smVhDKpRMeWiDNEGWZJL0mJnu/PfLk9dB2XaFhkJF9kYFXHwTbD+AyljWZmsv/xSGJGBmOXrmV
6n1fpL5jOqMak9f3dEe13Y1jR+RA7k+2+fOSogKD4bBkfyZpo4FMvm6tMRy11E90Ux9yxL52tFV7
dMl/cuqoNgulo6SamPfjO+59kS+Y9nGJKqEZPRjLWzzpjVYCIsiPyJxgLQEi66oyBOADExdhicDA
Ry0TkwaGcAFypUsjDrclonEnoR1wDIHck43PPZB1sInRarjghNG4MqMQnGC9hP7/cC97lEnQpzgF
J0OpWnlFHTFd5qkVlvozau9Vs2iksjU5ycAH1eVtuFyLbsb5wAqI5sveqA99sb1kF1Ai0TAvMgev
0gy3RdCKqDU0EavWl5mFwqvGFzDhii29WQ6gCqL+zs+tdAb01t283iWyF6H2KAD9nB+2vAaUp/Kz
kP6ODpbW7xNr3gQxNuy8ybgHvdR27clHsQV/q/bGqL9a1rtQhNFw+IUN23yUB0Fn1+9d8pbOsbQg
vUZoIadgvgL5AzmMIZwpy3uqhnJvrVw8y2lKm/no+oj8VjSc/quBmxsoflQHThmOzj9ymSkEp0bK
ZT2DJ2KLSO4Q4tKNHqz4BxjSqoYQ0rq8RWI34rBj3QD/sdMjcvyHJGfJCygl/pBkwZPCdjzcWuVU
JWaEm/PLXQcs6HN50UllztpYpIbEn7/3Dyz6KR1qx1hayTZsQJORf20huXYS4aQdWZ491Fc2WwNy
JEpWxkPhdzvjatyyC3h/Ug3ylvg6S68u5t9xx/RgJaBfeFAG03D+tykpTR8QPPXDkob1Ki1aHXWh
UYHLKSlbUPe0w8jK/0ebv3kLkPDRzt5SzwUGE9KRC2IXVSW8tbfzNHMxUyUkPt+ngd8IMWP0IFKn
5HqyepJ+gHdm6Imva6IWO3zQfIWUefYtb7r1CLU/+Q6ItvhL25LINbZdLq98dZdUfKcSIApjC2mn
82Z78i8haKpn1MpJRckEi8HiKUSnKfnTeVFe9JYV6momgR/Je6WRBGX0/669qq4SWhNg5acFYBnv
CSRk1EXWb0aN/TVtlbxoKPLJt2UXMm5j5VjqL8MANxUcKlSZK/xogbm14fYtnk0xHUDsb4wx61jn
24sPZtc8Z8QBcn/mNJ5BVfmnDHkIica8HIxSxWD7mwiOaM10jSUsYxbv9QICv8Gb57c1wlxiFaH6
StgZStC8LuSSj6zrX5600p2LSo8hnnWkAQfAalRV23+sdIESkqsi2JrfkYKK4B4VEv5+7fPL09kF
Okgkp7uJJFyVPiE9Ax2oU/Z3LcSF27PF1zmWMxjKc3XM7CQyoO66Hom/4EphfJojWzPz9y7XR9NR
qe2kydS0QNQ8ykFlMF5Q6h75n53na2vE0/djbOMI2Y/tLuc915E2utziwFXBVtv/aczlOCFEebBV
2DC+iDR+4KsyuphFVL31jj3xiCBfcwNxp4Sf6HsGb5W7/aIMhJE8pVLyTqYEwGfY2R/ZdM6uvEvf
vDq0PospU4IaCM/H7G44RHs1RmGC+ctmefNArDZOxyLbmH/eY0EpIC3HEsVYnV1IfA8yaITTKZP3
UqNFwMHeC8g1fZVJ8YxWkRhBH5fZtAt1Riskl1xnaL/Yg5VCHpO/NLfit3BCdtRAQZlE0TsjMgnM
yeFKKu7nnAHdZbBcO77j3G/QpX9UnRAIeowHCA6se+tgEjKw0MKvxDT6Cvpy9aCM7XE7ZNss3fjU
CxwrrcU5lfP+MRQ4QRB8raRnIhVT/XpQgm4NWsKpgFl3j7WbPvRkO4o1Cgd3cN9S57z/oLn35piD
MO+QnXNGR4Lf3MkIND6v3/BXUnor00D0g1lJtoMYTeY+EAbKIHeqZTXb5Ruy3UxKc/OVXsUbrg6y
hUmkaU+ywxXcHlDQlTwXA2fbjr5JhJo14mXkyRddyeDZJR3iBWc5qsV88gt8z1UhWkY+Fj8qyY0A
r525aOsG1qWqErleOkd6wwv8iasvlwSkloKipjY4fwlWW7nhfdA3CqQp4vDie7Rvb5KgEOca1NzL
zQ3GfJ/4nQf/pc8PKKPU2xyGNvT7Xt9WdUJGklTirlUX1AqlCXbCEgwpL/bTPZtpfjoqlaWgiuTJ
sXWdABXVEzIQOSIFGxpqEzqlzjqbo5W4veXKPRAQ7/HnlVHzdXN47UIfjzR08dJ0T5Z6G0kEsN+Z
1LIHcIUTofSdK9ulspPBmSTYceWTOB8UyNgA9r6Nc2z6FttE7y+PKEnIuk7gdC8Sgq9araRncT6e
7I0j+RT3nuunDbGGr5nrGC/urB2pff59kt6yb6UhuKsEODvA1LiLmTS6hb+sjqJPCzQ3u0dOnaVi
KAE1UCYmZG9PPAmHbG9t2hy0aXDaVtcU7nG8ESBnj84LoXnsFDEuFmgipLqSk3mfAoybw3/ZQhim
Kj1n1Orr8cCRreaiHLY+B7bzHPNLONTPSGJxwyFhWdTWhOtJlkuLjfkJKtHzhSoSTzPQTDoV7A/7
h8POjtrpjBbsZcyphoSPXcaX8568wbnLVv/qXL8VjVp0xUbY6Woq+0Lx31OOiRvjliSqkMw0iJCS
XsOZvbBrjPOBYRCkYh39m06yg7Rzo98M7Uiu7QIJdlYh3VAOHP821NMtghSWEIG/VnL+z5/PlyWb
zFakhTYlQJoWQOG67Su8UaBwfB1ojnZkceG+wtVOd9kmaUIji6hbHtatdllkY15Cv3n27M5DEtbj
umadJrEyp82iIqeQJbXP559lNFmENXLOuBQ917o5aUDaRVKNnouugTds8DBXgXjzQNzwKuE/XFoF
wvPkWbQWeJ/DX46ZBgrUy3An0tiGHixVrotniwLZVgBiFVHbueZht+6caXE2XBecojDzif5UKeT/
vPf/gVcT/f9irsY7PbgqFgvC9UBpSJGOkMNx1v96IS7PMsO0hWx1fFPDXZ3hTUWBzDh8oRp2M66b
prsZaEsQ8a5jJ1s7EZzu4/7v1uWEfgh+E31TDE5LNbZo2Moo0JB3RT47O4tvyS7Tbowr2eyHrqj1
7XFfqQCw9vlJyD98UjPXKGyAJ2zS8l2Zm4ziRxe/nT+wts+7P4WFecQ1xTwVAlm7ENAOhmXV4AFH
lB3AkxAfYuVOYxzv+bnXKXqe18aDP4WrMs5BjURa4/ZXxNdM0FraaKGPLTUX8dfTwWo8WKgxUr6m
qxrC490v806djhAbsgxoTPgjJmGGA3KJgw6UjdzcgFzp3dlg5MfgJzNfoMnpeCH7qqxOUe/l9X1+
B+mq52jojk3YozsLAYr6n508RWjsfJVbeDnd3gLy0M0j3P3opi9dCpT13WBgh91i63gOkLvF3YYI
DLEXGd1eAqpbSKvrYXZxsUbEL9XaTr1Bu2JJJ3IkZBS16K0CZoRMolh75RFrCcMqRFss3kqZtDlO
mRDD5dHM9slZssWSWfGQKGQgwSztSavlgpTfnecPbFA0AYo153z+2QJPzmgrACHFcQ3BzClgCdh0
P4je4oDoRP7rAQwG2X2F7n6nMV8LtbJCw+8nGHy2unPYqh6LXdmjuZH74986wEYnN830FWTDGI47
R0dAW/D9kYNuin53xjgYuEJp6aIwf6ozt755wzXrOXdNcJW3DDKjqw4BDjlr5myh+i2Fy/cksRZj
kgM6JWcaCjznuuBdSU70t0B7N+LFa71HCupyL2b6SSSCgHUHqBBLh6ckwciWzXeLb62lloRJKyv3
ejWq3NdsoSZg8gajJwNecZawjszC40yoxcmOHWyuFkKeJxjNOg4HYrMqdyDHdXWWHSBtCiZtuocw
Osz8P9B1WOsWM+vaRM2SMAYjbiqW1z+ekGI/v0FtcQFVmBk/TLAe9e9xVSRoD7PxEkP6whrrHcej
AsFkCFvlsgj5JEV95ddXjRLugmAGkGRnPtfqZ2zsbLVnyvfQt1fgSJgSKa3q53h03lY4XmUOtRwG
N9Mrc4MNvSukkWnYTqNblBSppoHAOShjGfQljaTKju4IVxmfL1qWm7qfhdMdyqFlZJ2JM9eZrSDx
QN7tgK+hCkxpoASoKbIHa9YGXTjMX7TJjVk5YjPvkb5rcmlSBmDfaSS2L/uCQIn96ZhrvJCaKbOM
+CP8PCSUAYdMqeryPKzlyIIYgKFUY6/V/3sJq7D+skmf+IwIJvV9BlvsruXiUZDAZ1W/iouc/Igx
2nbisBJAjzl87pdRgjh4iT1cB5bXxh+fW4iWDs/4zqNyHOHiSTkLrzf3mEz3aYtsY98zlSr2fskT
eDOyySr4pbFkJMG/x3pjTe6PDmaSvAaAiEOlQdRJVzQO4JYfMiQZe+hQI6592r0nl7t/CpHtNg0p
+Dibat0mkEwTieygsjKs1x9EKfFNYmTJH+rulRLZCgeF1T8KaOjThDDNT8Qri3LlSTgBxDD6koc4
Y4WKV5WsO1ea4212NURBd53qPzQA6XeqF2mCFh0dz94P/JZJPjzIJi0lllxqqrBPW698cZ315OK7
5gYW+Q/fbvMfmEDxNvaB8DteuRrN2jm7lLCNwqbbaQkaNeofXq/qAEgDytoEFNQVxwoUQwyLRgn3
oHzsubK9x1Yg3OKsxW3y1wGB0HdheCLM6pEWuHQb88M5J0tqty5sKtRZK3GtHzdsYZ17wdnZp9vW
l0ljCbMX4vqSaCvN58tZW+3pzjIip0rFPgAyQvvUfbvuVj3GeaRYLFEMDFHESOC/ZJrRmwcp0qhA
hxP7oAEzT1sGbfrVBw8Hl4NyNX4uqQ7ed49dvhDdPp1g3dzZZzOXeg0YYTV71HEfs9YfHQkAqLR+
u4SfnaUF7IeA4RL4nvNWW28Qnxd0CDn4Gv6xm1MOlfAwmPQ3RZCs6OrgEHOSEMEbJoh68GC7vwxM
ZSsCbghX2r4qjNNsJT397x3TbZQnZxYAfiuNLwRyv3KqRezrMvDQwgI30/fWFsK7FYnHN6kOQx8D
+ff8HHPhogjAZpe6cn3ZccXApDnsyOa53rDmYYg8MBEfGmYppkXZIvui09bYyssdTkOCE8QRwrJg
XLNOn1ucufYjqz4jp+n42HVG8G1C/3bR84IcCay7Z8vkFC2Tlr6tUljOdgo6HZ9ZBhvuXM0OiMs9
y+1clBo4BjlofWWBDYr1Yda13OLrbWJLRwq1AZq4ItldEL7SG4+8ij0xUljsLXPFhSEqqExX/VCZ
RTx1NfuxUZj7drXxfFV8po4L4q39nC8Enew6vgRvRm8B1vzh9HrG8Hk7pNSo+X8rDatBip5DAzpc
cusa1fEHJ9qGhQaW/OaIP/5RI1a48qCgoo2KoyZ42gNF5gu4gS5lntHDxyon/wVMsaYw3cU6pTXH
HLgNQUXsXsz8QqP6Ou3Zy/wFPMlXi/8V40N8f20TuST+3ZmyMP6oXj6iCg2Jqm5t0h0UDB56yYp8
JAlv7UGkW9WbaldfbbaQ58x3DldfJLLcEiPRR8yrU3LGfx98MfoLdJTvNOHu4SE7lXgXbM8plGMc
uWy8DMBmuSBw4F2TeA/EuLPsGg/CvFA6FgBuCc3XIFL8EoioX8a4+PIeqg74zRTPR9W82liBRSV2
Z13F6RF6Gvsmx2NdQiE6tw8G2c9UPbZKak45ZyE3RAnxoJ0VmaKs/utd5Goxy3XxFBAZ+53sJ8v6
eDxBKzXmHsm13mokWoz3ju4Ze9HDCqMYSg2LmzNGw4XHiJTpVjjlcUyutNT8jV6msbci1vlWnJ7F
tCKSgPtWWcFznwNPwrUjZP6y9okkJX84LNPLGdBJYnCuOA7mwVu37PmhK6UdN2+AS+p1E88+/+ja
n2ppxjbURlDec6OakO7j/RtJbRVopoHwzYRaMooOuz6kCf6af2/lGor7HPhEBMmv1Ur2bWVw4GPz
6ATUGckN3XMwdi0O0ySEUL8weO6wHizo00x1bYPdbuPZxrC2GHBUiC9UEuKfFxAg5v4ExaNr3Rvz
2D1p7agXHk8J3JrOrwLjjl1yyYNSOk5L0BqkGd0xHid0HFVV8VIA3Whclr2e1hDwIyp9OFhE7Wd4
AqNfAz6FJiy7ByI0DVeoUVq7BecJTahiqBmkd4YbTnC7TrzKp169p67+E23bkz9/Qn0G+D7Kkt8z
/tU1SuLbKtR75bRKeRCta+rzl0S/8fxaMN8Hy1CfJ0cEiQk345HPuiv9NyUcZRhbydnKt3Y0np7S
scFFZjScr05Ga+kHchVN1aBmrir3zxzxiBkHWbPUq1ansk31HkwlpMignHAA7rlXJR1bdMHsf7S/
lywrgvCkYP6fdz59LSkZYL1VKMNl3Mz8CO1DgHft2iC1jIoW54hCCfEeo1k01vDzPYZmtKbljds5
f5SMm0jhQTinXe4sAhZA7QalT1tHe2W8gN9sCwTQosDBIkBO1U5JRYwcDTOWlsdjxW7YMogID3IL
JeSpW7CnBGtlQClAPOi4poVktRpaO0/PS89C6Lg5iGVbD9TZtoWAsk0P59/+8jrvw4YMPKyUDcQ7
0MVIYWjzIOJc7pXEe83sBgMTQoOJT8dzoiVJjdYVvRzrdDuukSlLoufkshNdQD9adnf2P2zPCWH6
IjNHgjMxvsryJCL5sXmaJxygjJy6arjzI6SrzsRWhVv2WXOp5wvus2ROT8Seam1IIOHJ1W3DkwfB
jGOAayRM8p7GF/vXpQStRNrXzUcQyeYWvQ/DNjIbq3/tTc3RGOesvZXzV4L/I9vlsAGSrag3Cusf
GpBx4hYH9eLI2JSa/44qgYzxpL3DxOr4818eBTwkDINROecGLGxLC8sCLNkHovv1Q2vd4mzUCTmM
sWanC/rMgKjKu7Br7qK7niLgqhz+uRVKGhfaNRPdjIV2n7Qy3G+SAiFtFWuFITtaWfuuWV0qOrGn
/kmqh1Z+zWRC53M7zU9+xit8JOhh4UTwSfdtE7cKCzur9kfINEa6RqX25LcZ2+0BnkB76z7eDRbR
4y03rVeYW5CGCNm5LNFCbLdqk2d0xKcsgCRgVCN1GgbRpy/QNyXDdXHO7hw+zsrH0phb3qZ7s9gI
AbldhK9T/WtZcSi57BS5AVqY4wYTVQ38gJkqcYj6MWyLzm1O33EYjTPefYhzpueYvRkQrbYl8mLv
ZxQG1GG7kJlwuk5ojPjGZUim6x0ThtYjNw9h0P7zt+XvPKlO9nt+Ov1/1S1SRZAS8ikMWkh15KjF
GisQDbHhgIheH/NXBFCrHIkk0kq0ZN4dUAYp4pZ6C1AaKHX5MaYzly0p3imGN/chfqAS3cigFEGr
R5vuUsr7Am8A4EyR8CVhqu0Hjf/rDbl2H106kT5s/MCQuidUgQGQDp0vTDLexrGP6r7s4WscPcHm
k1w9sjfIKiRPDpughkcIpCr8tQOI9kBHcoP1oRBKwM8nztTjdhnZu4uEa4sTyR7u1+Mi0Bz9VZFD
A5EJ/mIPtHWQGWDwp5vtebXAeeKDMXfO+EPggH5VwcJ3aog7fGNWJH+rf1UEvpcOJkhtyU3CNHK2
erqnmpoUL9RGAYW7dLTqcmPVy2oZ3d1nl7wAvQvVJQsG6YVBtAkrD2QUuWdpfz4SS3iiTzkbBYQv
uFIgBUrTk/gszt/66UJN3OW4gjccsMQNYGxzZu+0SqtatbZecvc9YLUx0oKo8Xl7Pw/SGGY3Bbj7
za4qIHt/9rSFeJNVT44boDtkogBnWvlna/5roGlE1KEsxUHBe4juNFFQSoVO2y0lzASuyNIIEpFb
czeTMxtok/fzJm9p+Uf33xIg8UkaeeKN9MxsqnYG7CpDl0rwnX2SRSPq4Tn5rA07RJqBVcF1turd
U5grFUqqdOMGcVzGui+Vofhl2g871PxTEsomoEpE/OHSUvTgNaWaVQfEqUqeWF9mar+XYBmkqeQb
RMVjn5IXfvLAE0IaG4te6GVzxyonuCP8UiMLbe8T/rAttYmEVWmb5V1MzQJcsZ/fZu/wiMOusdeI
ZR8mqCp4FXHzFJM159ZHSLWAX06moXEzmWW3DWLuiFaxV/Iw7HVtGGB8eOBPj+2Ve0RpArGdLOvb
vnoA3B4oT59i6s4OHZlBzD/Mg2TK0YXh6USeU91D59BasRKLUFOXgDslKnVqKa+kmvdtoUeyI7MO
wDwMgSrR8IHhlLZXDqDqNCMeZiIoN3mXMhqLuqf2jj5pyVYjJ891yt56qb61in9/kMRGwvwClz0p
02CCBNI2/ypQr4kxkIMd6Rf+I88Sr7pbkkKVXIvmgaIRAGDIdrHrrCXUsIG1WG7qnpTOVQ5jhkv6
obqx4E9P91sjkooumahCsFmn4SDtGrgmdSXt92UA7VTMtxlIrjB/YQ1iJ/0uP6dCop/d2/XFdOpN
vMiKueYQJ46oKYFcZ1ST0j+/l2NCF1GFvcqhTt7rWmZPh3lZyirhcQhGJ5DyQahZSBodIHrKaNzs
O+VArdnILAdP51N3hb/syo0GS004BWstH8yBczM2Lmdw7USm6DlTEQQpRUiypZCJ39T4Z8pgQAPK
zPnADuI8mCNU1lkg14TFRKZHRscuTQstBszVRbHzw30puYYl8NyE6hx/iBcVzE1GOGYBoakt++Up
nYb98lw2Du0Dbf1rPdZZASXT2PA0u7ICtK//PQ4qO527cIFD8jnCRZeOqdcg/Icv8oHMuegJEeZQ
OHyLHaXnpVSNPckZA54v9VVQPEDcLo06jvLKWYuuF+HPKsfS+PZcEw/eELvonZ2b8NfyLl0d6/FS
EBKKZpk+z0uamHBgly3CTh6/ur2NcG4zuCspnnnC/tQJM8isKqFsBviBN2ZaNaZWuK9kZLMOzlqK
LRnvckI0ZNXbSe2nNdY4qKaFhV8oICgs1E7AbQ6+i4tOkMY6UTcTFVSevXrFnffZDwPsh18r5NOK
tDFWfjbz5eS+vIlrXXDBjJ5QM3qFj6YwUSULfrZ0iAWnrv0XuKu1NQjCjgvFueqC0GJOjUEWb5+b
ftXsxzJtFWgB8Khhce0dXZpSGt8LfXN8l91p6Z4tsnWUuMmBsFE5TD3JSBX54JO1miL6334eeWBh
egH9RFJsRKhN7eT8Ho/17aOonlcfJnOB1eBupg+uzp06aMEOlR8tUc1/q5uqw+ZYkTafay59rtoG
sJUy+gZMRB2C+hmtO0MkBA30B+QFMFgshjLUP5HDV7jECUZQglHgxUXlqFxdLtA9UPtjdh/BOFl4
UtE7E3UUuDkrWrZP1Z7wZuYk4jO9YterHR/2kLs5Z4ecd+LdDXfqIm6RKqXK/yFDOke1WH4l9Cis
NhhQG+3Z1Hq76yD39G8lCdVKtKkT2LNvpVPXXU+5AJSipODvXE7j9x23svc/oI7vxAy8MKRZTUnq
JGlIQSjDJj+HQ0ZWhys4lYZbDeThPJPkpAqme4Sr/vHnQ30F2eOhH1CXFOZKVbAUY5skslmQ47gU
mpVvSPF5/LRzaDJ80XQXRC6Bo1KsHIteffZEKO7QNLwicA/frjDlNnPYx49qVy/HfvswVTs7SOWp
dPBWMadRcfjdounpvbGuHkUiJqEXDDKYw5WnnnTgiK95dbOxNmAOiAP08ssueWoyD15ksH9Edqlt
4tf5IqSG6APa94omyiMKmXA/OwM/AbyrzDopSINcr8lXadGdKUI8eHQSc6jLiPlQHQMElWYeA3jb
zmNla0ZRyp/XbMc6LCpNKsrvGWaKlUV+oWBXvvFWBIuIjKYKNyznO9QuH7FYM1Ajii9oYc2QFSnh
G0Eb2zfJGoDOVpBVAUVRlTnH1c74VctDBGTWYh/8HaSbSx9bL50xp2f8e6CFsBBkbDkcqPPetwkL
GGJUIuHA9dcdUFXiFpxvTG1Cv0KHv9NAroMdICwy1HphDPQQbJGi8G2Ib5f3dlJpedHL1T+jJHis
ocwHf4R4Y4Y1CzqkbsH1zspbqYQCr2RKwqoHIS7tBmCNCa2jmyLYwVCx+K8tLS55mpcOPKCUaVwQ
U7uYSYMbBPkw1fvDmeRx7frPl4d+GV8mycZY/FiV9KWeNKsbodVF9TPBOGNMlcPOSPIuFa5fXyT8
06F10JncTx3+NyIEpZT1SzeYb+Kw06IqOW+zmBHFgIjACW5p7RWU4YN0sur0b91cFnqmZxC6H3YC
orcu+wxW1ICOjF7knsd5S4zK0TUJjf0gSaZH5DCr3SVK6wpS95fHFYLhGnMDxFkPeIIu+wDxgk5K
49AMTGDT/ujCOvfD7MAWp+cz044o9IglAsfQr1C4clEt3YSoq5j2u60FlMzOWbkSB5bx6ZAeqktT
iQdxA5MmFYEGa3jgG8XHrtLMU59G+stTCV/hXgDPSR8xcFUQ3vxvRnrL9LOvTzmC826KitSMtUXS
J5/sUZYPF+EpqyenfEm1OaLtF/Wa9x5cjVaLMXlRIRRh91039uA2TcKjmH8nzxFeczgWFWt+KDKf
ANautaEezcv5+d486iwY1O+PKeWNcnd/pfCCqvSZNcw1usdY7rxnxMFSl5CC4vGxYO7Ug2u4LjcK
hKLfgTUroenLvcdJ1sUt3ZUm42cP9B8lA6JCZDxVBCSYKQd/WOdlkYDkVFGBGMyj4EmJ4u87ZzQe
bNDMm8jHbF9ZhGPl6LJ+WrNqpMLwJMwMCGMO9jlib1VShmfCSfshoHQHmk8qiryaZeECNo/FNKsF
+d38kmiBqBp4U28QNatazkX+PbL8gT3gF85VHPv6niwcOpweRcGhqCqXHQAmATo1jhOS1bPpoo6g
lLaSwZB5lwBEvCjA5ClH0kNb1B0y3OPlRoHwRoH8zAjKW9JLFRAbQZ4PD93nBItN8l9VdnDNVjMi
bTLtrmJDE6N7q6PDOaejYw95JNepTmdLlS+VBxfl5HFLEVB69oAgQiAxrZp2vhWWEVlEeJkGm6lQ
n05mp4VrSZx0+osRh7MzOktmtydmJBYBjCfUM3Mj7uUNx5V6AsOi/+3APsbSZhM69YJfOpt9+Tso
Ln0rj8stmZHYWgvQ0lit4EpfGOAUQUKB2n142OFo6tiNDcEq09VSFhbXhhkDoGuqeOiyJ+a1Mdwk
MyqedtVCmNnkN6Rc+rgdXZjlKSZ/udfNRIzqfmBxgVI4zC7efNpaMuVDHP3XdGhAlI6c1jouEw2E
xZXWd0SwJIxhbYLVkGIogKRwFwvTy1m/ArtI59dty42js9g073IJ4kUTsMzP0gQPm0l+s+EYtn7D
JpZreuPH3KaNIzxKZqYCv7A/thk1lOdqGwlBr/7cThIoBIhMokGvRCquZXg9+v4TxVarz6r+HKBt
myJc7dzO9ZdHcc5bqHmudz4JjpqRLK2j1K1uoRff3NtsM7vF+8foh6AnaCG3tS2rwi+Rwaazkwzk
sCMDzbaShy9iGTe7iyTm3UrLwYNqItAE/kemwRep27d0mQDKlfmSj29NAMslGed49XBluoxsJSet
nv8FSJJyRn9NsKMFpEAy3nGElwKpVVD1rNy1WWaDil0ZOx9bpTjHR3P7y46iEStznFqldSp/2q26
QqypKCzQDOhwsIuAi0PhlNUeUOSZux+/Ye2WtJaftIN3OaLkWZ9yZKT8SiB2NW/39iLMUOQTMJ/v
UMNDw6v8G7gvwGU9/ogsqf7RQk85Cpzf+FzfHUL4zvaqSdxoEk2pO+cPpj33wvajqMWgLYqgKCJ9
vuLgX2SMZtvwaITNDtdUZjfT8VrreUBcLg09/pUhLvaIm/LSBA4c2kW+PaRza7GU0X/hwujkrJE7
w9TV6tPnlKD5WSUd15P/x/SD+2qACJOeeZa+WvsuRMHSTLgHKFtYim1j4SnVf0/vcTWjhwHzJmiK
pMs6BiC4LM1L88QwcJ/DcT89tROsDvMjK+3myTKdEIsaJmMfXfDGXRB1Y9EsWHX8tEc3y9GhLtPi
x1Bl2tvcV1+oB/ZCHKvsnY0i2u3oxPV68NaECo+dWVt55nR5xGQI3JF/Zj7mkzevBoIXbMXjYiiC
09rY4wUUE79tOfTBLr+AHSBKdTV+QYk91rIM+SErpDAVCAC7YRLmZ4zIGZTMts3v2KsQno4tEW90
2HXLimv6VePwGSw8i9RVqwgsgA+AhHIjksPcDm6RaLkZFwcqYcChwFU6ktZjQ9nh3aCi5M7r+w0v
nmBXAmtcG3YK/yAvG8yRiSlaago15145ACsbvHvsrsDaLScqzMPLAfSaVmS20A==
`protect end_protected
