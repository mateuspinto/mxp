��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��О�C�?���'G��p�q��R{�ZWn�`�ޗ34$ͫV��O
[j�}�Rzt�L��4���=��NO�D�D��":S�����h"�����-�M��K��QQ����NG��|�����[l�=�Y�Qs��ii�_O'���x��$U�T2"T�4�E���*/�_�-�.����Yr���F��uI(����m�N�)2�;��Q�
@��9����L���#����(C����^��� wJfY���[�ik��+j��V����?�xR8I	�p?���g���&�rA?��M	��{rnUD�.�R�舵���w���!e9ܶ�E�6�?z����PQz���A������=^=����I���2��6��sR�UD���U��$Q���ŋք�b��.R��K�\kΫ��E���,�<O}4y}8�Gx�.&�W��E�� !�S�C2:��U��qz�Y��t�3��T"tJ����a�>�7oI�!hp�Ņ����SD�x���1��>�mKlW�6���n^eᓩՔ宓�S��O<��!��T&U�^�hJ�b��������i��:�uf�y�5��[�������ƕ�D��R���]��ɿW~H��h|V�K
UiC�q��niOO��sٻ;/�����: �'k���H��Lt$��I]Gc!�ub�a���}r%},�.<�&�7��j�ӸԻ�+����}<󅋑���YTha�G��6fB4��� 09*��+i:ܞ��=����H_��lr�)�I�GN�Rd9�ɱSW���H�� �j|�ȕ-3M�r��(��*��<��ޯI-'�����X�N�-Frc�̿���E�CMU�D��4��as#���F^��}x��Q�qY
�(^D`V2M���˓e������a�b®��K�w���V���y9��(�%g��������]g�褓y`p��2	mܙ���`��H�`��d�<TX�A @٤���-�$��ӤU��c��"Qi��YZ���?����+�5��^{� Z܅7���"�wQf�(���VɸR����J6.�hm������V18�������V��#vD����r���LSf�O` n�5�6YAi������B�����t�Kϴ���l!��%��v�b˥�kg� kCk)Rx���Y�i���PD��E9A]%��b�z��=��F��1E�$3|P�
��ܛM��qy4>-�®\>�!QS��0��Q����tWi����RqSε�χ�\?<���V N��#F-<���iy�E���ͳ�UOꤗè�n�.�-;���?�N��/c�� �E�|�d�SˌG�ͯޚ1��� ����X2��+�z�� �uC;ip̼����gNl>�0���$���B�v����R��7��Ɯ���,x���؁Ս���y�o��}�U�"bm%�jsUM2� 	K+0�P��{<	�sņ�����̀(N�?`��̹��L?=�!ꢚ5�X�{��g�θr[+�Ɵ��U�@�"�Ɵtkm�IR���nJ��c{Ѣ��L�X���WcH�����$�-�3a�Qm]xF.u���	"�c�)1�^ۂ.�ю<&�����E�wLa���ĕ�S�or��n�kSL�ŉd�5�>��~� �H��\�ÿŖw�.��]�1���Kk�CNn����G�Nd��'��8���y��������)#򉋹^�.2v9�v�!',�<��;�G�-��Dy�
�DY���͡" !n7�@��O����U�S�d�Y�0h�R*���p9f+7k��]Ά~A�]G~�	C�@4��:��,4؂�3�'
�Ώ�=�#*H;��{È����L�f��CIo:Q�|�9&�X����z
E"t��A��}V*ut�J
��Q�n�'8�0]���Zb��qQ(�`��o}`��H��f�on�<�@��0�g��5�$8���}����e��������a�2�����5��h]m�&��t�R�e|�Dp*�cE��{+H���W|N���d�RO��GڥáF�~�� \�b��Wt6�k�qn�u�L+4��+�g��:*~d�Cl� S1u���������ݲa�i�(�ã�=��|�靀�Cz6��c�Xz�
���?H"(� ���VJ>��L����ż`�4�~�t������Pc�X�	���_^�\-��~��#潐5�<�u�!�2�|c�Rrm�!�-�2n����Xk+�@��F*t��u�49��c�ᐳ;	���ӛ$o�p�c��Qt�y_�4/G��?Lym���A�T�U��FeӽEK�! }륧��v�����D8绊���'��'��ч��>�q�" nI�UN� �|�,Q�;�>���84O�ۅ@��'�2:�{W����ȣ���%Ҟ�H��^�0 �)o���s����"g�A��-�RL����	�Q��
���,��NN!!Xu`���C�F�˅GN�I��Xbz2�A�,��Ą˱ٷ����V]R�ӣGxT�%J
�f�pD� �ٸ��O�	fD@��i����BlpP(H��gA���7��.]�#�?o#�ч@J@g��S̋��t nuV�G���m�8�N�!.��#б(��8�T��y�F��qW�J���G*�4(�Kc	)����B���w��:ʄ���VtVN��яP������*ߵb�Nm{j����c&V�����!7���O��QƏroJ"G�-���*��D.&KN�u{1�p6�(���-y3(�S���t�A�s&����H��}2T�!�Ϸ������>n�$�f�?!�Ď��oq\W���ݕb��f�� ;����{���#��P���2������1zNF9���ݕ�G��ܾ�q:�-	ֻ!�tQ�Q��-g���3U�w���L^��=�E����,N=��5f4�^0sp| .r����� �t�3q�'�~�:/eV2����8�������w�t�~���B"�sA��|��D��Ｖ&!���1�cuSv��C�*��upP ��T��u�2lO���'��X��^Q�B�`�i"�PZ��q�n�$�p(���\�xӵ#��_��!Wbvon�S�Σ��ZF������(����ձ�&N��,<����5�T��3N���_���`���ɭ�M#�`i\�r�+�և�o���B���!���l��¿3Φ��r&�/S��lB6E�v��jg���$�v��3�e�b�C�./�x���sZ���%�'�D����Z�s޼j����,�Ph��]l:�#������3��ˇ�"���Ϥ�<g��BC'_��p���_Q0�2�5�����+��&�{Uw�3C
�p�U�PC�Pb �t#�?̠E�<�h4��}U_(�3�������Ry���v��,�ƮeI�C�
�1���8�`��C��@-�f��PR��8�@�����c..��JJ��68�ȿD*�-��aߝ���T;e���ݨB�Zs���H�M&�E�M.�L�GQ�\/��ʲ0y�S����H㬄�@�v��uǔ�y�X����ǈ���n���;ߕ~�[~�o	6`�w�f5��0bԾ�D]�ƒ%s��P4jͣ��*�Y���� ����	Z�R$�E���M�X�F��Ȋβ�F8:��������?�0dK^���W��|c��{A��������"��\������*�s�\ �D� "�U�O�������HF�r�N_*]
��˾@��H+����tJ	54h�^�)�@���U�m�M�[H���Npu�u�%��#1M��SS�_���i��FU�����gF*��W>@�2��VS��^3����|�Dv���&�~Ln��aA�zvʿ��hWM����T��̏G ���Fz �k���0ԛ$�<-��I\[ʳ�1�/�&��Z��~a�<������|�yc�d�RF��'B��+�E��k�!*��30�B+�DQ��ҁ|�4�e���W2/97� V�Ok��b���܎W.�L$FzM5ࡋ̨J���ƍ�����f�Z�A�w�D��I�yi��{XmT��s�I�� ߾�6����c��톡��4�rp�J�B�
��՝�5�HDIG�Ę'����7,��x��/AvP9������딜�z�:��Qy�`���3�&Ū����I\'h7�d>/���
"���=?xƠ
˸���o�K��E�)�7�z'�C"_L��_�E��+�I\L>��+�W<��or����`�i�9�-'����tiD��5=M���؀��4���п���׏2��Y�iZFv�`_"���D&�`�4lφj�]�\���5�	;�W�W��*��0�D�=͹��c�C�g�Cdl��S����!�`��E��|�� ����u_��x5qr*��E��g��|JC��?���:#/�Y���Cif=�D�Q���*�DϭH��B�M�L'd��'�7V:i��O J_�ΦᙇPz�Ξ��Q��!��XGG���2���cP�O`�Y��	��#�q�����w����hC�oҮ~�p��=|M7�ar9�Iv�|yN�i�����x�ۚnWg×�I&�����	i���F���4���y�E��)t�y5.ɂ��!���љ#�|#����Z+��VＱ�ow�뺑�T��?qs�	�2��[��;����SR7xf��
�Y��GL��,)�?��`�����L>�>u*�5�����l����W.>�3������2q�?C|�F߾�'P�N*�=��B�>���2T�d�y):O{�Qm�0mb�f�RaVp���."D�
8����P]����� T4�^��b�j���(u�2xڌ�Ӫ/|�c�g��r��� lpDq�u��*��D�����H�M �����]w	��|SJ��h8�0z��MH-�>^g���/R��{���@�e�a����pa��rt Gz�M�[()��L����Hcf�B8k����~�ẗ%+uE�C)Ǻ���4�Ƙo&i����!g	%�g�u#(��"^�z�8yG(Ѵ��e�TDJ�y�0�Gd_m]���Y��lP���v��%����tB�h��y�����i��^�=͔� 68��v�[h9��A_���~U���C�S���e�I�i7]�y_�9�@2h`M��aQY�% Y�h^�3�� _,�������6�6,��#O�=�Ճܲ@�~�O���`H��X0��as�,`���3�*w�'Q���)_7Lȹt|n�rbu��vH�u�6�_�k��[�K���l�)�ߚ5y���	����g�
 D��<(a���;|�<K!�z���9�����C��2�r���k~��@�MݥT�2Q~_��(kɄu� �RL�O~�p-�?���o2����e�-�Y�T��6��*�kZ�*ӂ��[����@>h&���T��O���uGA�҄��/���N����7X,C{��",�X�\��ӘhTi���O�4���:�#A/��<Makq���!���C2�6��K������ɧQ�C���'��WM��=B��H��C�Y�Ĩ�.�kx�
�!�h5��ڱ���)�Y��W�UF7�������1� ���%�tR�j���Řq�"�1�]2����<͕�8�YŅ��}	�ӬD�9���57��fxG�ѨX�mz%���}1m��kϠ�P߲�f7GY��|��P�G�����˥��%��?���c��I�|+�p��y�i����W�p�44d�z\��h�B����6����ݠ��/��k0Amas�O�����ƙ��π  [��T��F�����M)�
��s�sg�����պ�� ��vu�vZ�T��e�&3��bp�ukX��s�g����� �"�,&�u�k!@����cT�Β�X�d�
.��FȪ��y�"�u�ؾ��W<5H1��#��T
uG����g���l<FF6����L�/�y`�f��u�K��M�"����z� V�J�7�^���ퟂVg��	����]߱x-���	�)�b)�If�c&Obn2ѿ��{G�kʐ�����זҖ�+׏���~��_bosΕ����~��h��ǲq�F�$����!�W��6�O�p�[��0]�X� ���,$:��˗����A�}�/@*�����(=�`e��Xq��ơmyT �sr{s�:���|��?��K��`t�h'���W �<�sDPp"�%�K3�Qb��TN,�܊_�E1��}�{��