��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���@�ct�: �t`��k�r�i��ʳݴHEL�
i�ޗ�d�X�iP- 1SC�M,&����1j!�5s�E)��
����� C������rl���[�H�@
^g6LZ*^P�2�0z��u+�����a��a�7��&=QAƸ�,ֺ���^4 2�م܇>�p���T���¿�#?3'��� Ǩ�A�R|/��������d����ꪐ��#��� ��m�5c�Վ8�V�Ji�C�zj�Y��o�kH�`�9�8M����y�jD��!#&�3g�X�"���;���ڹV]>+Q3j�b�4d�´Tؘ�!
c�r�ĩ��&9��� Q��0��k.��5�)����8��Z m���ՐՙT�s��_���,���$�y��+=�;r�J<�����e|턉�MH��;E���C|�0��d��Z���i�G�����m�~��0t�/�i��o��x�6��׾3Ʊ���@�«g���>��!uYo��@��Xf���M�>Yot��c��C���c��.��~R�U�n8&��I��B��!v�4ê�����CHĮ�%�A����χ�����v�	~Ϸ�}�=}��`�7�i�ls�v~#�7�Q�.�^4��P���`�{V(`������O!�%i����u$�V���"��[����șQ�ۣb�+dqQ�'C�x����̆\M���e��v���H}m�.����vgpFx�`�L�4�3fV]�?�@[��VA@�F&�ueIzF����!������N�oga��Q&2��Z��Tù����K'�s��!�b��"r#�H?�#�D=� �8�DU$MN�ʽe�O�D�֭�h��|.b���Wٔ*�8���,?0��朞S��?G6{�������%z��Of!u��|.'�W�{@ ��|Sʣ��傭8��>�g>@��DCj%�1w�����7b#�'E�B��o��a��+.�������e��VTUxS����(�ٶ)E�C���~��g��p��o�d�|���`Dа�b�o���ԍΤrz�܏�m��x8(p�Ո @����HX��r5,:�t��󢈜�ޒ7�1|3�(�T�������9���Peyv]�G+��Z��}Ԡ�kIZY�	�)GpY:}@|>8W�ҟ�oϒ��a?*�=�|$�kO�o�IU��k}����΋h�x	Bw@�*�XL67A3Q��髶�-Lui|�B�}�#����3d�`ċsj�����,�@<�t��`h�y|�@���b�J$���L�����s)X�K��9#?pv�����tL�4"7A5�xc}Cz���@�pQ?�&Lľ-��@;��E�Q���k|!�����\m��|��S*P7�����T���)N�W����FR�dLfm�@/E��@N<@[j��}5�4�6�b��¾��X݉&�Hk����1o���l�*�)EV�=q~]���Gϊ�
x�I7/��5_����"qX'���U��i�/׏����<0������a���b	^k�J�812�*�� C�f�ƈǾ�"O3Yۿ9u���܌ �Y�iS��E=�:�����<0֭E\��<:� Q^����f��i��� Z\��w]r2�7�_h�u!�!��:<V��`H�5���������Ȟ]u�~�_�|2v��6�0Z�gX�15<L
�4��3i�+($� n����u70+�����4Md���u�(��QZ��8[�"�=�K����8U�}��@@�!�%���	��fF�it|��z���facX�Mz�"��x}�5_���`��9i6S���[٪`p��I���zD��}�6�0`i����/��c����"X"�5�y�Li��$`٪uij�}���re�z� ��>Y�x,Lz7��꧌>l���銚%�
�����q�mVYv�6p���~�84Gp�Y�i5>K�R��[�9�E����y8��GC���|r �P �؇�dSׇֻ>l=3ȟN-:�0�J��̑K\o$�@JQ2��x�鬼�(K�'�����:��%�� �D8������'�5W�$%Y�|�1�5�+���Q�A��E'+��C/�$��k\k^@�V��	b��V�  � ��C�&��_M�����%}P!�7��(ue����gƲ)C��^�}��|YAx�A��eV� �����p��������h��m��ul�Y��RT<��A���!�]���q���6%��,<_;�A�-]���N`KM�>/����R��H^gX�A�c�ˍ��(-��7�&�7�A�Jx����|�	�j����46�Ǔ�D-*���^���µh$Qu��g-|W�[qB�#_���(O+݈���2�P����Co�G+�Í�桩��<?r�=�v>�ɟl���-q�OqV,�GU1���`�2��X���w~�s1V��C�Mѵ�<rV�����\2��-/�Z�6�Z%�f������w
E�tj�O�ba$n��Ji`�����wWen�1���ܘs0��\�>�q���Y���w�\�#�V'H�N@�I73�X�����vZ>WD�$������]�ncZ��i�7���7>'�=e�T�%�F�]����6�m�*l�Q~�v��[��������p!A���q�n�D��K�%����B��� ^\ꤰ��ɀ;�`�oG����6���c��u5�[�r����7���Q����Ȑ�"�\�q��y�w�b@��;����:Q��{���ܻ�Q���[��|��z
'T ~0�(�fN�%k�� �f	Qn
Rz�R�O]���@�L3tA�0�����S{"��;j%h�eʹ\�i�6H�<��I�'xF��?%]�t�e���JqǠ��e�O�WuE�2X�X��t��S�G�!M��l�h�w��T�4�?e�߷�!�3���S�;u�$vߖz�$��W�(�v#�`cQ�jJ�[��M�@��Ұ���uϫQ��<53ӆ�����u�M��r �����p�؀Mv��4��e/_I�;�F�hh1 �аz�1 ��Q�]���t�AG���b����5p�$T���B^Akd��\-V(�;-
��0xؑG�ט�x�hObMY��c�a.�?2!�}"t@�)|�X0fl}�\l������ ���-���Q���z�#��4g�9MYz��[��e�'���.�J����1�������;��r6J���dx�j�5�c�>ͳ2�5u���x�������av&�/Lڻp*�='*�U�_&O&��HN��ղ���I�!Y�����Ӿ�B�����h��4`�S{5�n�y��������j+�7�?W��H=�<��� �� �c!?6έ]��-�nJ=V�u�z�H*QqzGd��*�5������5�.n�4�K8���w�hG�D�l�/����9]���}�R[���n�f�r������'�	E��e�TOYں�?�<�q� ��ڟ�	������x�a�!��V�^q4:e�vW�^B8��?`��)�X@(��C�6�Ι�n:��=�Dm;���;�����c&r�s��D�$(,�
�<�ab\T��<��434��	B=ꊓ�V�ǆ�>ݷ0}_��[q3���yՋ���0�@qnV	6<�e
hiz0J��<�*���֑��$�sڹ�ߠ*��j�����{���Cy,�$��:�<�@ٴr��ѥ��#�x��]Ё �b�Ե5�^�>Ē��'��,��*��"m��e�-� @Z���C(*l��H�oO�mX^Ԗp+�U�d�̫q)��^��� ����/뺥c����H�C>΁�S
�dvϦ���&�X�eDm������'9?�(� *�@i~9ҽ�[0Н�R��ig��M���y��o梋�vE诺L��|�_�9�&���4p2i:$W��U������o� ,:|��p�:^��Z�v��)�j���Q^�d��Xǟ?��?�������
F�~��Y�q�ܚu[��M���o	�؏�8��\dfU��77�k���:b6T�R���P@��|1�s+ח矜x�/7�Ig[}���}Ӫ��tB)⊜Q�ߨ����LF�p�vK��Xl-	1�bQ�Px#l�/ڔ%��W��]S��V7�v"m��L�9��jL�����f��厇�S?�t�[AF��SuXH z�1,~����x@v�������� ̗�+`IA�����o�А���s�H5���o	C�T����^m�ң��_�qW�UEs��ڂ��$��k~��կ�E�C�=����3T=���8�^��L��R���,���|c����p�]��>����挭Ð����5��MT�yx�A�"^��/��o(����h!DI�&E)?���^�/� ��5œ�!�����K}�w �ūE ������(6z�G̼ॾ�Ր��IC�Ɵ7I��
�={b�[��8{�i�	>H<y9t��1��f>j��R%�HNz��A׿J9Fj�Q��P���4p:b4�m1���~F��[n��^ڎ��{�4D���Q�k�.��|:�O��Kyvȸt�߄��n���(؅�
�s%R���_xI	:��O�=b8�1 e[���Q9���	�j8B���7�&���ֿY�G�ˑ:Cgk%|�Y=B�%ͱ����)�`�G1/�r�T;�)�2�H�U��bq,�5��h��!'����Hh�Y�c0�xeҭd�\�	쒪��O�螄��^����r#0�f�������̌��KOI2H�N�_��^C�-�4U�����T�����l���s����яn,Q�}/"�AF�J��5�.�L��)3ʇpqX	M���R�S�6��xK����c����$�/��R�&_K(����mD���J��IoK�k��o���æӻF&Id�y%��c`{%6���#G��������������x6OF����w%����4���#��!���[�\U[I�]�Ip#�v�X�v%ozn�	�G�������χ]�D�2:`�vi4W�ut������f��%[���C�Z�5��r��x3C�@Yx�,���3WT�RVɍR����\b��ū��,�рn�"z1n�4ɪ��t/�As�\��Q풠�Ǿ�M����d��п�(,�9�,.Eӕ-���t�նi�즠V :�S��c��X����"����u��G�b~5��,.���<�uUK�?�B2�#-o�<��\SmL��b�:S�	X�V���55x��C�C/�?��D j�����n���D�7�n%I�	r`��A��*�'b��h�l�P�ː�_`��`X��z�Y�R�hY��c�jQ�0���
�|����R�,���;o�o��e51EΖ�������o�b�gZG�"�giP��|�ϝ�i�*�kg�߹�hӱ�*%׃c����2��'����%�U��rh�I����xɃ�s���v�~K�:y����A6Css�k/�(Cl�4J9=m�ʡj,����3c��uy����%I#��C�`��m�U�
�rV�2�/�7ҏ$-�@9�3͜�W���B��~�mJ_�������+�d7��/H�>����.ry��b�'I�<�@�J�%�(�i�x�ө�%�}�ŗ3���+��+�}��?�K�)��C�fɃ�v�Ź���)����sB����쒱�j�"6�Z�Nl�N�wP���^��H���uNŌ6�!L�G#����+�Yow��h��L:+_B��J�1��Y5�1�_M�b&��/���Sߴ�hڛ)ﳃH�ȱ�q	��ξ���\Qo�0v/;{������@׌U�>����P�
p��p����k�J�H��0�Q���|�ˣ�|�J+a��<�w����}�`h4�p
Щ�Ϭ�j%!�0P��
؈e��h,�ᘇ����4S��?l��.��c�*��Xq7.P(<�r_N�.�;�[5$�T�V��fk�Ǯ�wk���J���'�%Zh ��O5��fB�--@4��j@�`�\�ڝM�w���`m���6w��bJ*u-����p�l�#{\�8ۜ�ui�A'��~\��k�>ڕ*}�TƊ�Aw���V����A
����(�n��s�*Y}���a�`� �����~ѧ�}���2��O)|�W��T�:�S��g^��ۉ�Q��D�{6�n� )j\֑�!����zK5���o`�P\��,:��k��^yvvZ]�v���g�%���ݛ��͠���@��kfՃm�����׷UH�R���_*5!�b�ny�A��D���ܾ�خ���-O�`����Qر_�M7��{��K����o}�;,�5���j0�S��%�lH����}�������zٹ��{�"��+�G�A�?�sC���R�=����<�|�>�`��8=a�#�G��4�o�eYon��O�Ǜ�7.������`���� b=؎:��.�쭃�M_�,;wc<�rLa+�K?\]���Za[/"��_����FB�����W_�64e5Jf�)*�=�6��]ɿ�`s�EH˯��׍⼀ە)lF�7��@F0�O+B���D:���׺���d���J����L��,�n{�[i5���n'�.�k@l�	q��2�j�/��m{���=3�2P�G�N{�%�a*����3Q03A�v�#�q��-�>t|���#��)�A���d�4v,�|m�V���^�ͧ�a��ךD�~Cf`D��&��
�@��}���_�!��N�D�>�T��x1�'�C��ZV��� T��G^�A�m^ê;���0ܰ%צ��#�e��}nz��
a����u+�똰h��l����B�?�`^_�M�;�$�>6$�'�&�KGu��ܓ�-�m	�X�aK!S_2��,_K����/^�S��aT��uyl�l֖�68Ǫh�М���czT�ԝ�!�ٳ)�Kb��������0�����{�Mn�>�+^��ն�#���.�����E=�C�u�~�(ܙB;`9)�d�{
��������#\�B�ǜ��(���Mav�9/�O&K�Ð2<��ץ~�����L~�{�冷��eh�|xU�t���e�cXj(��G�ҎC�d�"Y��z3�P���[$U��b��%�����&���M��:�UQ>����(F�:���2IY�zX�v�j
�����F_�,�3�Q���K񂛢��p�a�+�D��|%�����;nJ���$�"D�)G�ªa��4�/Ʃ&�܃ �G���Y�J[*j3T�8�A�L���
VƠ��Pĺ��G7��_���n��Hxʮ#����_`�8�sd7��}"'����Ψ�ix�<-�-Z�脝c}2�.~,;�%a��uח��%r-���U;)�C8sA��aZ��ON�gʙ��r�:8e�Z��E��2S0�nX:���¤�ǣ��ޞ��>���@�Q ���߁.t7Wv�ny�̾�m��� <D\�'�p4�R����хb���7)Sp�'# L ���f��'�[��{��-�'��B\o2�o
��1 �5��j���q�W�_L�y-�Z�+E��%���ϖAo7��Q������G�Vכp��>۔㶉uwP�g�	��Wq#9R�&$�C�\̼|��.w�b��^{h���t������4-S	YŦ�����:��S��C�_�I�*�IX{����_���&"�GQ��p:����1z��+����D�̙sW��z�a@���>r9��?)�AF��fI����K��K$��"h得b��
�$P����OS�UK�cBYuC?R��RVCs�)�߯e�����(�7v���>����\��pP3����J�
�{���1F+W��״����J�Չ�3V�3p�T	��A�}���W�/̼��[t��4�\E�#T�7|�[F����1��l�ˌ�I�/;&�&�q�a�S6�;�������9ܥC���k�$�F(ΰ�0��;� -=6m2o�ic��Ͽ�t�ɠ,����Q�	u��s�i� }�W}����Л�<���|'���n���[']aS�I c��t��u�m�]��-�3��d~Q�I�X��uXH�Pe���s-O�>�kih4���{�{)N��Z�3Ofu���GeX��Iރ��ZRAd����sG��7Fdg���B�NBs�c���BP`�4���ٳ���n&�l|2���gݕY�B���2�x�����-<���t׾p��÷���+� ��'��P`U���2l��K"]<�A�AX|Ѩ��Z�a����9PX��npr���U�V1����4��q��>lC��n9|^�@��C����[w���SKP/��DhYpL^�*6�"�e�Lly���_7 * U��rD
�Xxǜ���1�N��[ē2�Ƒ��(8vN<2x���rԮ#1�p�e��	�˗BqpZ��/C�ԷP�e����#Cs�s$w��d�����V���qP�N��"�����kt�����5\m���H�m� ~I�0br�y,5o��h49w�qg�&��i��B�O����Ҹ֮a�7Q澴�^�A�,O�K���o�m�G��T��s�򴊁Qff���Y�@���S�įѝ�c/�7�	�RǼ�B�Ӕ7��JW�_vwrf`р�K)����a��ʿr�#~P�8��
�^Fm�7�&%q��$nL>s�d�2j.�|�J�򳙌ͨ�2�%t��s�R��d7��lm�Ѕ�%��?t1��Ȭq�o��7�P�|�����Y���-G��#��3)� �I�Jz���x��H/]�F��j�����l�� ��'S��[4�N��яӐ�X9TuۈO{6l�	�o{6y���¾�S���F��Ф�D>��y��*b�ß:��ǻl��x`��rcLG�G9M��"����"�3T+7��]�BΠ�)(�4$[��e9w��-hb݇�����.wt ��l��v�w��R�}4ь2V��o\l��J<�5Sm�LWm�p���n��6����I�2�hJ5\8��t�9���ۢ
+�6l�a���� ��8Ko���;�W��A���j"����%�,�h{��V��Yc��2���ܺ����#��f��د�7���t�<Ͷeк�.��U�v������(޴����n�[i}�Sc�ȪӉ�M|;3F��*\9����0U��?��
��-H����Z�?�ɍݎe z� ���	T]�S��
�u�qr��f����9�9j�p��0~�6�Ě�[�8�L��4������rf�${�<�fgr=TĦյ��| �k�B�����S
Q4���q#�b�-����J��f��� �9�+]�u n�y6�i�?>J.�0N�p��Y��Xڵ�ވ3�PǼ��w������j��;K�Z��s��������3���!��OhM�X�AT���ե�z�������07_�]XBA؃|��V߅'����Y�ۭ�G>�c��0)����4pT��'`X_�Q�w�kVN��|jwVk|A"�[M*U� l�o����E4X���O:ב�3n6�eu.J3�WyZVOB����5[8��*���
�u�'�����7� Q;�|�W�a��)�X�p�}ު�~���G m�.�S����Xefa,`z��l)1��r��b��" �$�R�74�s}�����߈�����3�c/��Ú�Q].h@U&�ǲ�ނhi�s�n��|�g�/H�&���U�F�
3�z���AP�N�h�S[��ED�Ier���6R��\8>
ޯ%�
���
<��9m����j���/�DJw	Sf�(�m����Y�ɺ��*��+8�s�v
OJO�)�D۷�� TVv���V;���-�O�W�l��Xr'C��s��I�{�����Eg*�)��l�'׺@�tKɪ���I��Wu�?������_j�{"yk�[&���QV%����4T��#�{@<��@7C�� Wo�C��[�`��WN���!���p�7���:�$7qgyG3r^���B�u?�_��5x�}�v��0et�7����߅���v��d1I�4�b�&=2@�%1�9B��� ��S�R]&
��� �����������Ձk kh�,���b]�[�iV+���츕������y��)[p�*M�n����� ��&YA��%̔;����j��C܄ap?�LW��\A�tU���|ΎY�1x��YЧH,��f2\�L��_s=o� S�!~��6A�!�;è��zܷ����{zǩ��
@D|�Wl��%C�g�1B�w	QN�n�������Xk�̯q~�Q=�5�j|��Zl�x]�CL��4��V�Q
}��r����שּׁ�?w��̯�� S_E�J�����%���b������I���ܾ��B\����@�C��-��{��Gw�n���4C	�?�es�X���$�zp��>��x�<��#�	z�ZbC$�RC��FiƵe�y��ڪ�'������`�N��J)v�4�L�m��e�͘�8�(m��������'I}P�Q%�t{��'(Z��U���G�J�'�&����h�:���;NAF������:.s��
��X���@�T��ENӫ�Z;q7��ȴ�{<�ic	b�,�|Q&zcўir������pH"�,O3,�v�]Uc
�c����{�-u�����
-׏�����<ɜ2<��
}�"�,|t����٨�Bj�P'.8�]g\��hзY3�$9�	����S�q���|Ouax"�I7F+	:93��=4���5�8*���L!ck�u^FC��(�tA�YP�H��h��׮��}�N�he`�˲��'��m���Т}/H24�A P�?���BkE}�i���\ ���M?2΅+�r�љ�ɓ��j�s�+�'�8�y@�=8G���?1��h���\A˄g �hY�p��Y������z~��)Ω	��]�0<�������&��X`	�H;�N䵔"l��献�u�%�P���:;�K�y�`E�m�4�祉] R=\���Y��4�g��
�{]y��� �M=��-��{tb�F�N�M����1�T_��~/�&EW�iy��H��� �VC�����m5�sr�GL_م�Z,�\���m�M����G5�=Q���?I�\�.��ܯ$V�*J����=Z����O�MT�PV��M�Rް�h>�!��!ϓ��bw�%g���6�{��y}��Ϙ�w�!���8S������\4�jޕ��z�M�J��/������� +f�Ԁr��6���Ԃa�3�b���w0�j�,�_�zY�J{yٱ%����0I�!|9�xDT�r%���I0�fZ�x���u��i3����6��)�XU܊I�ݦ����ڙ�?t&RޢI_��)*5�����?�\{�#b���L[�J��!��NUT�+�toG�����|�R5�_���x^����<��L���x��a��/���zv�����d��\���[���s"c�O�'�o@��X��RT���G�p�>�����'��HX��V��q�?-� ��T��*&��ӌ*ɖ�,�����w
q�WA�j���9��sC'��WՁAXE��w�p
��i��I��Ěd��fxP�+�k��ř3�S t)Sx�2�"�EƮD���u��'P�e�v��,�x�x�'�zX���'ϟ#�ާҔ���kJ c�IA�-x#�r�����
�߸�H"jxOX�9i�_2��t=ޮ�\/��>�� ��;���ϒW$N��ʥ��`y���4�o
��P����1E�0�\���h���R��$�s�n����1��d#1b)�9��^��, %�舩�-��e5�'+H�O���� ��xڃ��f&���Qן�8V���&,���9ヴ�c������L�cP*V`*��K�I(�8W�[.�lJ�j�-�h���c����L�s����ja��K��H�m�f��j%�I��Y����m�K��)���{yӟI'�;8-o��9��K�'f�a�L4�O��b�rLh�܏,�/m�&l@"՘=;c�����p:S{;r|��3 ���}��N����|$�}�����T��΂/m�G�
*R�!���Y����P��<�w�O����#カ����w0A�0�^�?�Q�(�d�fn��K9)pF�5��)a�@��Z��l�Z�"��X.+��o;��h��b��tL%$6}��9og� c�}�)���i%���m�ߛ��V�_2�F-�7�u�nA�� �%,��E��T�4�V��2\(��d���*W��}4K��S'��ID wg��]��bkS�YV��~ORV'�����[���Pui����P(��
3 qɎ�a�E�Ɠ�ZJ�e�^3R��9@Ub���c>e���1EϬ���J\H�ɠ����=ζn�v?��o��W�	��N�PWK)�?hsیoϨ���DF(E��Ϻ�Qh�2�U�$��81f��̙�R�{�g/�#A��,;#ѓ-q� xg�o�O��cT;ިY!y�$��j�� �,�	|֫�R�)�
�p !5kVv$�F�ř�|��w��W^�%1�7�8r�e�?ݴ�x��|Bt�1u�
RJ��c��n{�M�X	�(����5	䠚Z��Q
��~ � �?|���&�C*�ԃ��]$c�7���&�����ۗ��ٖ�o��?��'v�Ckؔ���K!��J�ͳ����%�*�2��&h�ʭE�NI�Тn_����<�!�s���J&g��s'��M!- N��ď���Gr���W"��o�Ɇ3�"Sܪ���Z���[���wdT��k�_$����KRuߝ��g��I�i�U8�\ip�;��!2��v��z���v]�ə~j8@J���qy�3k�
�>Y��:���8-:E"ZO6r�R^�lf.��`\��D�| ����m���7P�G&?�χU��ߔ4|�!|��uϺӁ���(�S�LRX�r�Y��&���Ȍ��I�7�E��m�c��E���4�饻��Nrz��cqD
��@��N�rc^��}�=��L�ƣ 6��}ߟ#0�l(�,4-�6w��Hp�!�%�8��M�?�x�WԾ�@�J�|���s�6�mҺ���X��	D]/{����+�d�#���]���Ve�L����2������9��$�Ȋ�zK��կ'm7R���*G
Y����?Xf�-����Rqv
��_6��W<��?U�f����,53&A�Z�A� �!���v�I�iQ�G�9�h
�����l~k��^3(��p_�Y�}+��?�X�D{�l�$?
�H{a�u�kU�^oO�P���j�5!�ϭW�j�$h�;/H� ѻjouM�Lâ�A�����3~')��"�%�cU��M�(gޱ(�g���ف�Q�Zg�&V���|m�gI�RyHbi��P�Oy�>�\�s�Ȼ��^ ����ЇzYҦU��-���(\���*|�@{s��n�ɝ�ܲq��9ؤ=[���𤁹8a��Y��<��*� ��9�}9�!U7=�5�����w���5��>��۠+���G��'U����b�{w������/�X��QLZ1pod���"�"��YLK�'c��iB�d��1�:�;Y��Rz]K��x���av��e�R��n�:�<���byl�I���8�mi!����N�b��d�)�!��Ɖ�"RMW��NyMʉ�z
���p��mCC����#��Z�Ŕz�W2��ih�/%���	�ҩ~��vc�ؙ���R�O �z$�2*^A��W�f��n�4)�ǽ�7ﮓ��i�eG�"�;�/�[a�Ɩ{\s+��)E͸��`y|�Ê?g%����0ŝAP�B�l�x���V}�ܶ��1
=ʠ� L;�eCB�E��RE��fA��;�š4�*T��e�.�?ٯ
j��˚��u���iU<s��{C�v �ޥ��U�V0�W�(s�ݨ��������+��;�͒:+�Z�\�OC<�_Q^�6^cKxbQQ]��Ƀ��]i���Љ�Ά�P�[`}4x�t���Ʀbn����i&����8�N���?�g�!�n�x�_���e�������K0;���k���Q:�@GI|�ˮ;-^�?
^��h�M�7X�MSsc��lh��"Tb�A3^6�J5P�h��PJ�cqrs$��[�վm�j��l*y��xsl�r��� �,�Q�� ��c��V�2��޷"�E�����,�j_���p��p�o��C@�
샰 ��:rD�݇��)��d����8l0�ϟ~ua��N$e̮n[�,jx)�}峁&��4<�Un��Q?�����a���/+��B����o.��� �\]�6Rϑ��}����as�B'lag��|�<�0(1��u���v9�s��0�ĠJ�r��X3o�~��ד��܇!ZӪ�/F.)�K8����FH,�I{���2J���֭��sF1͵;]ؠѩ����{|.��]C��, �on{���ouH��%孽�߃��w���9"7�=]G���h;�����P������iMz�I�w�=,�|�zp\�<
xC0����[�}Ë,UW�%��xC�/r�.��q�	��^�\�f5�c������Ʈz�hĹ��0s �\N�
G��ٜb�=����NN_;ZR��͛0_�sR���N�Ys�� �}�\~�G���YH���<����B�*����o�"Zq��\^�&��&e���`j��$�vu�2&��M�ⱗ�>T���
��@�� AdD(&��&`8�{����rq��˯�	���f��f�����6&y��XV�(�����x6�xk=z?�t#���vš'���m��,�%�!6|ь~/T�D�L�&��C�V"�%��hx\��V)w�����V�H�1�{# f�"�������e����?��m�!w���νr�I�M���.| T���0���4H��,�Rq�O�G�W=7\���g3����Ƚ�	�~�<}�2�w�ӓ��&�E�]e�|<��$7�q����Σ�᝛�B�OBWc���m+�t)25���T�=1B��Hgc���3����4��|:��7�#\9�lT�{J�����r�0|��OK2Df��*PT[Q?tY�vm���_۷�~����'ž�u�����!ᓣt�A�����׹₊	�lѪ��\7���G��c����#�v� �x�<5nV��v;�F�g-�T|7e5b��M�?Se0hU�Gw��<N��L��f��,DGg�(����9�
��:�@�K/:������b@_���y�����)��t�c����dhr_6Ȯ4�qW� ��rnz)Bh��-����N&�g5'�b��A�6���)���u2%Q�n6�K.3���+$o��7�Tݾ��g_�����y��=����a̤s՝yk��\cǓ��o�p�%��*����C��i�K�D�^]��)Y�ڄ��QҌfFɨl��+���-l�lCm�$����)�Yf����qd<C}+�6+4(�1�4|��L}�x�_�p�v쨉��r�_��}�DG������hx��d��=L�A�s��I�9/k�]�B��v�
D9�/I��3g;&�����q憮Q��9���z>z�Cw{8�D��j���m����eA���ñ蚢Ay0?��M*�kA���'�tU8���r�&����Am��;����w��}���Q�Eٺ�kj�9����jdv��ڂ��f�k����rGԿjq�5�8��~�I�r�Щ jqg�����a{!�"K���w'o��J��]m(3���|��UDB0��/�p?�����1���nX��I�;}�W����NjSR�C4������rz�W���J���l�$.���$���J�j3��H�s�Ƙ҄��
�I��K��g�M���ܠ�O�{^��@q\��T��`���#=Ɗ������с����$N��&~�u�-���3a��s-�|�x�Md�ܻ�I�.C&��^n�+]���S��U7.���C��Z��#�����}��4op�hEğ�
[���Y�vZCM�d�ND2��K�8̃ʧ�>�n�^�;�BmE[��6/�f%52K%�J/߾�y`&�I>�{ӣ]�k��W�m���$�6d?�1� �[ȵ���-<iI����ۦs(�r���Ũ�_�n	]�
GP�T���p��>(R���$�,c� *r+��偶p�E�S2z�|ـ�
3�pE�p� *n�$	8�b	Ȯ~�|�	���e���G�Ap���Hc��ֱ8��j�t���}���˙�}CG{WfA3����u�u�,��;d!X_���J�x :����G����SѨO�ω�f8��y�[G�air��ĉU��+�KĪ���2�2j�W�>��.
{�@}b����F��O&JF4ؔG��P|"��ؙGy��A�5P��lD|�u��0�_���D6�s���$�z�[� �����f3>=? ��m�`0������G�n7ĩ������-n��>>���n�W(�N��X�=�/8/s>{T6�&����
�ؕ�o7�+Ɲ��4T1lj��y�"r	��F?n��������
3݈�4l�s��İ��F�} �o/Ǽ��4��QŮ�L��jzE�yn(C�B'r51]i��~=R����������i�I�q��d8�%-Va����T��	�}� _��p�_\F}�5�Irr�)T�1��9-ԣ I��*)u�$Kw��X����4��P��'��*�^x�'�_1��Z��R^zi�Ό�.<��-\�1y/����o�i9�/"�>H�um#�A`Ƕj�(��!Q��FW��c�D�1b^�d�AIFy��5�@�V!h�X��d����3��2's(�F�*\�؇������?��]�=�*��\?d@C~���|'n_P�������I�����qrL��Qm4<�b\D�*�hzG|#t�!�|��\�a_����S&&{��G��c���K�f��}�d���!���j�pV,
��nsrv7�
q�����dq*yl#!Mt�������K%\�/5�P��p��rXs�e�7 �Cp�)��LAg��>2U抓������]4>ޱP:2$�F,��{�Wtb�h�03�q� u�@fڠ')ɐmb��W��)�*׋��*�?�
����+�ţ[�MU @VP	��������y�EL�����L�6�$$%�=���MSxN��U<F�y��z���+�<�ٍ��݃_zD ���4熀�@�y�EК	���K[�C��:�_�6��*RmQ������\���&�h�@�@5���'�nI�ύ��dm�Q��T�xpPyJ�w5��	�Y�R���ҔY��k|�`�nO���;����LF�U$����޷��j��Ϗ��V���?1 a�?�Z����09E���b�x�N+B�&g������vO�F,�δ������C�����gќ4.%O���w%& ���Bs$I_���6��>e��ChSjW��)d��֑*��vaJ!��E�����q����Ī
���	�)n�N�I��kN��M?����_D���w�6(���������_r�>�	��p_���ZT�۵�d*iv�?m9U5������E�