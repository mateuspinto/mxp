��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���6��=&!��EK��`������H	�ʍ��^��MV�������eH^n�̚�x��@ͯQ��I�gb���28�{m?G0�e.�������V��-�j���I�-���
_�ueZ"Q�ߚ>P�UW^B �"Q<�,� ��lw^0'����$���z2םjd�!���)�{E�S8�X�U�]q�)O@Z�@Nj���"p��~���C�<W�NuI��%+��>��[���}Z��z�	�m��$�z��޴
Ž��%����%c�J�Q�Dq��>>�|���S�L_�*��x��}'�K3$3t� (:,S���.x�:p��!�)^V��e�T)���~��	�THh#$"r0/��Hl孾8����EF�oეN���tX��gXzR�[CQ��v�]?CҪ�� {5�?��	���(0��{)m$p��X!%6C+�m�%J��k�ݟ�x&�,��AW�_-��"�RϨJ�e=L�f����̎��m1�X�u�;�L��E��I^I,�AI��ڌ���8�=xU�5�L"�AJ�m�O�_����T��4"�Y�DD�x5��	��<�k|0�p�!RF�~]#X�.͜�V�z��{��'}���>Q�]�!����?�6�r�W>�;� emb"6Na�Jne�ж0a���j]
�m�����Ƽ�t�Q�A�ڎ_�~��(V/���ak��NO5�+J���kt�u/ܚN����0�d��{�����oHWc���N:�s�����f*A�6vq��]����r7��gjY�3��2��}!��c/?�C����]6�ǔѱ��AF�� ^��1������M^�²���u�O�PSA��.
O~�6��DnPq�+��������%����܌���U*X�ϠG�%L����Lm\-N�����f�폙��{[Qa���Lv��%�bvX_/�d�?��"sf?��qh�X�y��%9���+}I�1!K" (�D[�$�qD�t[��1�|�����h��'�+���V��М�s͠R2	��	*E�+����qEy��Q�߼ۉj����B�V+��G�|�F��$6�*M�����������r��bd.b���]��X�0�*��~!��}u���Q�FSJA��H�C�~�C�KDt�N�A�Uk�D�4meR`hzۅ'��]�	;��f�{C0<�� �/�~��V��V�ᄝ��o����¤3C��8�EG�"�#�1��Fe���� @pIH�4��V�(�^B Fq���9�Qc�É��ݐ��k�m8�C��i�8s*��kw��;���Q�y�m�7Z�����X�5��X3��5O��kD�|�����=t�yY�!�֯[Ɍ���^��� �K����y�l?1�}�:!����IP�yg�ģ�W%�?3^@��͢*�9���� =�x�V���?���� \�&��C$�& ��u�H�f��E�8A�?���L�b�0�[�O����ih��Y�PAon2��׆�ZF}k�}��No8��[�\��$����X�y �0��Av���/*�5Ӷ^НJ[�OJ^ע�c�?�
!�'"�jM`��^�*��OI�w{�(�.]]yТH���MbKPi�s���tb�Ll ��P"�Su`,?�T���"��F>�m��h�U��.5�� �7��*g�l�/�aWN�T�N�
�IN+@	?�M�%��Fw.�P!���e�d%7� ��=F���]�\Fk��Qf�:�Z���1�+�[-/�V���F4Z;]�.��ֱ�?Q���׫��T�^�X�1��B#�)L&x��j���V�1�#X���Ѿ4�E�3�y%�,�yDY[����dۅ&lT�����Y��Ȱ�:$�G^<��[0&�K3�ǡ��� l���r�'-��b�\!��x�, $�ضh�3���n*�p9~���/9^��0gt���5��9,�y��<_���R��ڳ>H|��m��y�y��t%ߠ�wC��1_ϲĎ��Z�t��{�i�	|R����=�@Ҁe���٢�N�a��۫ �w��^+W�~�[Vik����K3�
�OPά5�㬼/.`���P�i��`ʚ}U�HiL�Ta�#�-��.n���;W�F����y}W�la�S��m���	wڍa�z���j;,Krl��"����F�ԐUu ���b�7X�Xv�(Z(O����D�0w�aj��\�
�� �z��	����>�e{F`y �'يAnu���@iX��<OK�ٯ�]�~�z�>&u�*:y4e�
��Z��5�c�S-tDN�çf�'!���&�M^��������m��a�T@�z�(㪬W��ʞ�`0�͂!b�xˣ2��`�h?'g�h���*��w+����f�j���`��B��~����d��,|̩@�ر��%�wi��#B���o����<\OY�p�%Čbw�Pe��:L���&��V�\w�Nll#,���4tƗЁ���YL9^�ܸi�A�i?̬dAXN����������5�J�I� O>XjEz�Xea{z�����9`\�*�M���+���& ��-@�D0�u�sT=����L��d���FrL߈9�)�D@��{�\�O� (��Eoޘ&r��'�2� ��1���\�|����6�L�ͅWD�J�v�1���B�*������H.��6\P�?���s�2�D�'�)�#�5�Y\K�d���]2�����5 {emzL_���a�`=I�)C�7)}��p��o$\p��T�x��N����h�����o�t9Ƕ��3��D\(=������<��N�c=W�S$��H���|leC�Gtݖ����V�aw+���3;H83ա���j@ytgd,�5��=�u���+��Bh���
�3�փ󫚤a�9&��v�]�]6.u����6��ӌϒ@�$"�D���l*��Hm�QK�[�0��ͬ�:��A4]��i�.~���E��K�;�Y/��i��]���:b6�WX64���������ļ4?H��h��s��QuI����#��f� s>�>!���Ʊ"��@��=�эű+g��y�Z�S�ާ���л��U6������J_հ�����?A�k��߆��c[���3����0!������vW򪗛�N������@N.Jz��|�z�lz� /����ԩ�����@ Z�S��r+s�F�����=�F��L�
2nm)ˠ\Ra��;�^�ʾ!/�[��Yy�X\��åC2mL��)��M�e����V���)!�ke����n;�B�:�F=�L�HM0B4b̎�A�k�{�T�Ц���!!&;���l(g3L��GD��=�*���~���_Ŀ���''��+���f�
�q�Wjւ����5}�,zk%=O �p��v�b]�}��{u�+^���{�.����t���% �	nGHQ�E�hy�5�knxO���]Ol�~֟Y�3���<tlMSx�����u�y�
EWQ��D\E�>��%����D�.�P�R�
1���b�pѱ�`W�m��W�@�Z�j�y�t�m�1�o��2���5v*��tz�5[��| ��-�Vk�������r���4�əA�E�C�Z����J	дdN�
qQ}��V��5Y�t�Q��	�{4�kT]��̓����Hki��]��n5��.�|��b��(P�4��/3������U������S�V�ds��=̓D��u��(& S��'�-^uǼ�}_ �K+�����|"�O�秧Kz��L>̕N�tI�Iіd#�?���sl+5�ɲ�?/�p�X�f���c>N�>6���%�T�}�Oƴ5z#�~�n�S��߱V;���N�:�����ף� vr�1: �߁/�K|z�Si�C���t4Q��<%���^��po��*4})�m(��VM�i��L���f��@\��oN�� ͎�g�PĒ�Wy���w��7q��y��ݾ�Gg�#荄��NX���9ђs����3c�m�g�׵F| I��o���e=�����
mwD��:/
�D�m�*�m�kEqu�Yǧ�'_��y8RO3wTp.?��!M�'��1P*�כ��2���+���w=��N�X�f�1{-�c��]�}�h�����r�TARn��W��_�^'bRQ�,�cJ����ƻ���פ���㧈[ݗ��R�'υ���f�FBKP��io��kB�"Mʨ�ԙ�?C�`�E�d�C^������LaB�A@�n��Tt.qy,��6I��O�2A-�b+�g��Bg�S���J[N~�kG�1T��Py&�T�>�O��T@��݇��P>Y��{�3R���B���pE1�̈hD�nT���X�T.�����1�o��C�/�n�Z��r��w,�$O�98Ew�mk|M�Z�t���/�M<��n|Qu����R�{Y?i��Ŝ�6�q�^�nҰ�䰁]%��_��r.�҅�zڝ����̰�|�5g`^u8�Y�rY�ś��� �� ~""%�cd��T�1��K�e�o�c`5wj��IX����.H���^�;�ᇍ#=�YÛ�j�V`�[𝋸_��9LJyN���Lv����G�������q��3�z����V)�lg���S��̑��>A:�I?[}��F�B`�Íx�g
�3;������掁uW������ZɄP��SNf@����l�)���7�d�ȿ��O	Z��}�����G��G.��LbE�Ѯ�谤	a�W�'�e��j��O�
V��
/[C敟�,�����ҁ��,�1B�ZlTa�gu�h% ��9�R�Q�Q`RÄ���H���@�_ā�D'���/)�3��>����8Q�!D��J�/���.����M��Qe�^~�����D��N����I���.��?r�� j|�;{��T�u{��A���1�~s�p�,�BNǌ������!?���u�0V��$��κ�_���z�oO���!9<�
>���Q�����cѬ�B6�i�k���)vx��m�-����1OA�!��#�O���zHn���(�taR<!�j�_���2_i���.�4�����h�]EJ!$&��QiH��vY�׾�5��f���Gu��c��i��܁T���z\�c^����4	�F����୉� [�|��3�K�zߔ��a^����R�o�L�i'f���:�B�(啜y~���(��A�f)H��B\/�~ fa
JP:N��ɩ4
���O4g����"1� �n9�.K�9K���e��Q�x�+>Q�k�:��`j��T$㿶"Nn��w���ؕ���f@���B[�'�MW�6)��t��W�{��|�#;�������UB����Ë�( ڢlO�n f������i(v��ѳp���=��Ѳ�/��͋+6HV �>3J�ur��-#����i��uds���'��dg�'3���V��I�"%��Ɠ�wS�mkTh���鲨X>v(<�z�0�z���F�'�s�B�%��5�\��re/�|�S��h��Z�ȼ��?���Q��^��S0g�lu)�e��������T2�@`@;�9����+����"Ƽ_"%WG�XD��n&�W�5�1��94���1�#�&��9�T,/�p*�(%���A���n�~Z�I������ 5�G�f�z�
�[��ъɥ<�R�V]�<�s��0���f���p��Œ��
����D�Px}��!6ms�qƴq٧f�Ժ4Aݹ�;#9�}����p�B�B��0�
�]M����H:y�#Ύ-N�ިB��+��@$���4y#����ԼL��2�5U�͊,S�KF�f�`�},�*N�<d����h�w6� ����tJ��ȗ��̚F6; ��魘r�����mSN"�m�B����2�c�ΆU�����,7@�M�"����$���F��ħv+��o92K
�B�����`s~��؁�FB����x�#�'[��l�N�M��*�p�٥Q���wZ���MZ|����z������ g��")���S~����g��1��P�.T��+�^NA��B�o&��2������>U�*֘�J����<1�Ll�<ׯ��U��Z.雝m�&~Z�C�����X���0�ƌ�.A�G�w
����7��z�_�L+� 8��ui�y@���Ds�UE|G�{E�A}@n��#z�Q�y�kJ[��%�~a[�Ҷ
4��4��J�����3�"��Rqw��7�|E� �P�	R�r��U��ު�}���:�8��`��|w��\Hؔ��TO�_yL�ۈQs=ΥHT��bPѬVq��߿�������e��B����!C���V���r�e+��&-\Ʊ���P<Q���ɵ�B&�O&���8!�҂��<�$����� q��>~�{u_�o̷�d	�N���w�Os���C�X4A����Ϟ�ȜB�C�`�*b��EPP�0��}��O*n3�O`��1=�"��32�+{'�����߁�р�6etO�'ـ�/R�3�{ZЖ�f�b0�@��2�x�[����Iyo%{���t�k_0,G�@�S����!�4[.�.��9N� �!���1�ET@;�iڂB|}��ipX�`urx�s�Z�&��r���Օ1 �-h� �� ^�O�0S����Ej�,�o[�Ӧ�چHf� ��,y@�:�_��l�:��D|v ����CKR��z�}^�/�<`]e��T�2��p�Z�"� �z�fXc�<��s#9�%��Kߡ�^�������K�+�F$����5g�j�#1ꌽQ�Z)��`��fkC$�VV�jp����e�;�Y�"���Jlg���ט�9;��4*�98��F�
��OO��g[5)��_����x��k��C�zI���GTؽQ�����&*?_Y�E#&`P�~����Z�Z�}�fW����Zj[S�cЄ��ކ֋�c����}]�����$�R�țO�:�~�����XH��^UԱ��j���\lm�����"�ݶ���5��3�'T�Nk���:R���.�	��d 1oD1���G8���j$�B�@[A�����Z�(����x�w������e)*�=��%q�ge������"F[y<0d���T�aǣ�:	C|�7${{�5�S{e�an�1�Y�&�凖?�������k4bJו�u��
h���[�{[M�pl@�b��)B�Tn=�]���N�<��[�� 军�4�_)����[Hې~�����.|I�Q'Qn��)�_�A�� j������C�����_�(K]H�S6{�ƻD���x&�]=��O�2R��>ֺ�v��x�#�I��CP\��?�ٻH}���TZ"��6 ���%n猓��8>@nԊ޷�q�ġn�aE���)�54�TZX� slc�,��.�^�a+�cR#LE6���.�ۋT�n;;��m�	u�mw�u� �a��3�X�! !{ 4������d񋬕���8:zۜ��]�1гۚ�,��'��v�K�r��z��Y��W�Xa�k��i�w\`Tצ�ꑖE]h�8B�����JD��+s�)*�J�+��k�]���ݯv�2}μEJ�ߥ������������M�e��
502��D�ݩ�J%y�墯��PE��4Ƚ8��t$�f=��U��[2��P�lh`��S��n�6�:���_��4��V�`͟9��[��]a����.Ǡ����rTm7/�?.E��N��~j5��������DՌ��'�m��OZ��d��J�#"�m�Z`8oiUT�"�8��$�	G�)�NL0#}ā�����Tᦲӑ���Lz�?i���a��0��z�xh��F<��A�u�*���Ķ��UR�%2���|���}[p&��la�B)s��v��$n<���-
�h
�k����<�5�0��x{�D��<B"�lTTaN��8�vuI��L�2�LZ�´�'���U�»�2`��|��nŬ�\Ш������*�f���\�X�T��-��i����.%���
�0����NK��5��������%��0!�RMҌ�p��T��-�C���&2��c��)Б�8��][D�`��bj�Y"~�)�g�r��fxx����0��_��[<W���.;��F?�^@�7D;�Q#sQ4ohe���AYXa$W�۔�$�����Uq��T��C��c�Y#�Ȍ���O8��[�+���=�]��|���n�Ǉ���KH9��ƀ��<(�o�R�4Gs]��wᅎs'�b��w?�r�śU��,����v��2�>�Ő|�pYrn����;�uz翛�0Xl�)2#��HĠI�Kzc�-C�/Ѥ�~;�4gg����Y���f!-���q�� #�wׁ.ǲ��N��K!��[1�ͳ��w���xe�K���5�#_K�ĄB�xv��!�o���zJ˘����sj�������E���\�h��y�F��Ȥ^s"Ԋ�|�Z��^Z�o�s��ʟ�@��0\��w뾭�43��"�j��_AgE��~�Jk���n{v��s>��9"��W��E� X�9+��i����P�;.�s����HF��ND� ��>?i�g�R�8����:����=�b�6�>v������t��~��%2||$�P�̒�L<�%����: �:��d኏� �X��C�G�U���4���|��Z)�O-μ⪛�d/mFڙ����r����h3��Q���qd�������FQ�;^�s�S+�����P�ɇǳ �z	�����y���� ���H�P
*�X U��q��>�Cr,��%x��*��-��y&ˌ����b�,�si�f|����3
����5F��|��s��`�fƊ�ݡR�x��]f�q(��`E��MO��������h�s�A՜���ȋDN8%�ɤ���B� �q�=�s����P=T�ت��p?:tI͔�ݓ�aY.RY�Wl����N>[3ա���'�i��	g=1�����(Tlc�	�I�7�i�]2@���ZR��b��\��u@���$["?k��yD���~t3$ߗ\�,0��.3��)L��+(6�*U�9Ly�!��	�0�����ƚ�e?Ԧ���Y,�+�XX.ѰH��Z�]W���u�-��B�^�8�����]nd i�6��H��r��Af���{�\g$�B�� �W���Z�pRT�I�P4����y�,���ъ�����Z��ެ����)WX7H��U��&�;�� �2./�s�e�����!��0=MK]9�䔬�}�~kF>o�~<=t`�r���(����08���h/��G0�!�(n3��{M-3v�J��W}�A؂��_Nb���f*9\oE!����h'2��b���A�.���<�D��W��r�̄l�L22VB��eЩT�t�vGq�lg���<�sU[�1`�Qj�;�)�������з���/��Mt�*�t*�bՇ�����񼌴%f�o���%�����cS��چn�K9�%�5�yNc�py��V�x@��4ߠ�A��=��4{����:�|���2+�}c��r�b:�]�(�!Ee�7��TRB~h���=�e{�>N�>�K$��%�a��se��'�� ��QBd����[�Sx<|U�/6��$����--��4[���۠ζ4FWQH��{F��k�E��y�yŰ�����cph[��=�0G\I��W�cv��Xe��f@ܱ����y��:z#�ĉ��#&�/xV�,�wsݸd|�B ]�(�����iHA#�^��]_K�m����{�h��8�?BZ|�(4\���nz�(g��Nq�L�\�3F�=�C �^MY�Z�6� � I� 4�
������X����:��v��dw��	��Y{�X��ӎ2k΢<�W���e�wP��	]�z�ho���s}o V�ි�e2�Z�zG���	a8����s�0�����"�w����V��7Z�/��\�� �n�JQTqdi74��ߩ*��@s�`�ZZ������/��k��,&��w�/K���%�$�(���K�]��"�SD{�l�*�!�7�������jV�g�/%�XV+�jӍ�Nj�2�X0�G`@��99[�r�iS�+�z�*9ñ�ɗ��0�ի^���/���b,]�D�ԯ5P�I��aׄC�  ��/
´�U��3�D�b$�:t@{������ �Uc0>��[@�*5l_,��/=%����1����F�~^F#%�����_U���&�j����l�{t�O+>~�s7�|V�PN��p�'��:u���w���h���W��;ESm������kN��x΍?Yn��P!���Q�$�&��5��[�9'��ۜ�Ⲅ]L#�V�%���1mJ]	H޶<j��xVN���4� � ��`�\ra'�豰�<��>VW�
�����Mf��ɑ��J.�G��11bBڹ�E7�-�렧���Ө���=�� ����!�s~�E[��-��t1Y�Q,]��"�[m"�N���{Q�u͍�^��ڍ*ְ0���>� �Wq>�^+-�,�9ۈ��u���Q��h/Q�d�E��@�=F%cꯃ��zc����L5�ͻ��2��4��4�.m~	�/��(���UOLzy���ҙ��F, ��O[8�A�}|JUZ�*����y�u��EFM YpW�������1�.[�ؓ���ޖ�&!y\��d�0�jyv��N�ޙ'U�g\0졿����)����F��$�v�u�+!��d��~���[���{���s���a��f�\�e��oS� �Z� fI�^ ��h���]:_�t��7.���JG��ыAPm�¯��V#b��7\��Ac��(�5��wA��V�5����FV�"��í��~/Icc9uM� 
����� ���{�b�,������U��p�n_�y����4S	�e�����R�YD�x�>=.3X\Cz�~�͙ ��yTh��{8���'8�n��wxXڴ�a��by@��W�����@Tk�B$A0m�֩�ڐ�)���i@�H>rLx��6Օ�j	���ó�3��'F2ґ(�.҇K�^͂6ڇid�o��F ��F�]���ޕ��{�:gqf�q5!����x�Kv]JN�9�������R���0����c�դ!d�V@RG�xe�/�(������"�@�P� ��(�G��ҧ�U�,e	]7I?���wˊ�13��O��U��0�ƕY�d��p?:������h�8��#������y�1n�I�b��OFZ�pX�����c[�-S�Y�8����)�4��a�í�����	���O,�U>ś/�,�ֈ����9/Ă���w &���LK OiX��+� &���-����@e;r��i�Ik���v��}�7�ͩ+Z���\��q&)��أ5SSs��j��)>�4�˂ڣF	|h�����g�]��:z~Z,$��^��}J�`CH�|9iy×74�yAmV�
dKJ:��f,}8/�z���؀0j1�v����=��~?6	�Y8����ɐkrwaű�2_�O�iC�JC�\�`��!�~ܺ񂠲,W=r����V�ϸ��������s
d�<#_D/���z��P�P�ɜZ��t�M,�);���Z�Q��=��snT��H�1>�N��11����u87��p�zA�7�?]��;�}�hI�x�]G䉔�ufy(�AID���i���L|�)���ۘ�JT��R�_$�p!y|��f*�br��Eu��'�!ι@�r�c��qCZĕ1>	M�|{݉�F�1�Wh2�%VuI�S��8��c�4*���ln��P8�	(!�g��Rg+IH8��}��;	�eDb������eG��G?m嶙�h�t�W�J���~z��/��Q��6���*��
ל}ZCp�b��ls+��M��F��g��3kԛ�P�f���0��r�
8���{�S�Fe�̙��k���3��dC6ln�Ջ߻3R:g�I\�(S>�ţ^��Oe}�^�n9Ě;Ah�EZ^����� K��/��>/7��09�����j�������qT�IT�_��l< �ڄ�����إ�[S���`2je��`���ҏ�[�l/��"���?lf�X�Wm��^
5�sKk�7+�nF�MkVͮ���>Cč�����,J���ʝ�F$m
�$I�����&�O�c2vͳ��f[�4�7+%�6�PY˳k[���	�V����$��8K&��N�͋�~S���6�#���&Ux.Ċ3EΌ%����Zм6L�]�o=��8��(����
|�L����K�q�Yq�XO��t7��/���c<�z.`�<#����Iz�A�����gY&����ڶS��M�@wjG�(v|D'M�Y���y��C�K�R�E�s����]�2�q�?p���r�v1���%ua^�'_�=���C~m�J�o�$W�(H��)��.G9?>~IN�僳���q0�:�����������l�����Ms6��b3�O��˱^;�q�k��j�*#�$�wF��ٿ�����Uk�6
���pB0:��ΥF� z�
_(�e��*G�$۠�z��H��ԛ�%K�yd2�@��W,zCP�G~�����+��ųr�����3L��	9���A~@�Sz|�g����XO�}�w�J�=N'�8��­K�m����'���&�z��$�z+�Rz������2$Yw>jpm�K��5a�閸V��.�����
�,�ꉏ�]*�Y�����4|��V2�-e�e�8���\bT��q/��S��nt`+�rk��$���ػT����Z�,z@�F��6ѬQS��]�Pw\���ˑ+���H�0yn�VQQ�9jU1јx���%��-�k��V,C�l�/?r�#ls������^#3C�}�f��x�L�˶�2s�me`�$�S��ǂ�t<2�DwL�.�iO���O���B(qLM���8t`~�#J���F/���of��m��!A2@Bۮ��%���. wp,
����4�V8�~�"\�B=t�ݢ���IP�Ȼi.1&2�}���0��x��S�h?'���� 9�h-Lg����21g�;)D�r��6������B~h�`2鬲_�Q��pU�k��D�����I��?"e�$HN��Y��R,�;,�eʈx�B�F.!x`��Y�CF*A�F�k5�����"&��P��`�-2F�4�؟y�T&��,qQ�"e��K|G�����D�D���yvd7h�ヤ�`c�'_���O�� ���g�����1녪$�G�~ڟjԹ��q�v��t�������	-x�J�[ә��\C�τ �{Q���;a�<v~��*��"bx�q�eg�>��ל�i>Ż�1�5^W�b�H���x9�@Gp�������^��J��<}�Ě�`�Ȣ5N/��N���ܖ��x"�{��$�O�'��U�C��(ɯ�~��DV�r#�a�꼎n����,`��kox���{�N���ᶪ��Ĉp�k���	��k$>Z1
*�y�j�Գi�ȓי�����KE@e:|��8�����G��en#:R�Ż�`��r'��A���Y9tv����gQC��쯌ͣ���uXW�f��
 ���f!���f�dxxR��R�ȍxʈ��^lX:2R�R������`R��&��������U���Ѿ}d�\�>\�����B��2RP��h)p��B[M�
z؅��)�+Ż�Z�'u�BQ�a�����ᚨ<��+�gI'��<�KZM-�3v��E����2�/z4s�v<��\(����T�[D2��̓�h����!���[v�������!��'�~zyT'�y���������E��uQ�>�&����Uړ�)�fq��k����M��5��Q]�#��-�Y%��ze�b��:L�\�P���WT����yw}�#���E�ފ)���6_mi���4W&Oz0�N���C*/�MH"q�ze޸�Rrz�b�2%��֗&�si����H9n?���f�]P���m�ZA�����,� O�( +�@��w�{m�/��m-�����=��uB�#��5��Nu	�)����/�d����Wv%W��1%�K�������q%F.�E@d�F��E�`+ϴ��W}��{ݫqfR�>��p�i����Y���$�q�ahz�f���+�߈i m�M��odV��[W*tT�W�����`V�bΘ����S��G/�p�a�[iˁu"_�-0���� �t��Evq�9(53�0�]3^���5-r5%e3�)�.� -�P���llD^"�TJ��Z2�)f��-��t�PbĠ�^YX�R9y�b�1z�Vٜ�y�oj���*�wJ����o��g�p����o2+��EK���gv9\�N����.Z�s37$�^Uxo1c��A�_Fun�uL�)��

&~Y��J��w��VX�Hb��]6U&;w���31�6QIFDEcU���t+_�'Lx�b��3�JW�k�	Q���)�x��8+er�/�~��UH���T޺�xMx�T�	��r]����W�d/���L
�d.*��0�H���"�H���!-�gxVRca��?��J���$��@y��uW$+z=(��^����T��j|{�gzP�|H���� �׃w��\1���x�L��{o9 }~�r�䙸�:�pO)պ�{6z���O/�����H�3�#)Z���"m����XH]��_� ���ס.[�:�40��i�Tmf��-sTq����ڬQ���'�B5��A(Lj>.˟�p���H-���F���z͊�ll�6y��!d��@��mAg�x�`�:���;8��h9��.��=y'��!1�Ҙ3h"�'�r� '���[�`z$ ��J'5�@�'�h�����EP�r���u8�Jo�g��&��g�3D�� 6͝���R��������l���O�iق��7�n	���,2 ��g���#���b����zl�~+@ ��jK���u5<B�|��6�w/�y8�&��K��� �G�!�ΐ�<8�C���#�Դ|�$2;&$����4b��J�@>�����loHa&����\�nHS&�4�&� |��Ǳ�U{;'��p�\I��VM*В3�s8+�Q��^�S�% �M�-kUeC!�b[�9����dg�xP��;���9l�����;�y�>�W;���9� ��KW��=��)�80�G��W���x�<]<}�O����晡�u�{wwG�d��tlH:��?*���)S?c��Q
��A���n}���h0SY7�'0�7���E��d\���AK�d��ne3�F�ܠy�-�B"�	�D���<� �?�Ze��3+��	���4L�١{F	,�x��|��������%�[��'�,E=ͅQEX!~U����f"��S���i
�S3�#�^$�G�s���]�䅎�w�5�V`��yDa���� <*�|BO@]e����̟��y�����Ei�+-|"�h��jtv�sd��k4Y('8?�?;� ��G��,ٞ�.^��sٞӊ׍����r�&9~WE؜xm��dS0�#�Ɖ��$郡��o��[j$�4�5q�����a��-��S�N��5�Ut�66���t
4)4S�a�hgJ�7�Qo��t�����d����&��E4,����Y����+H�qS(��ݖ@��>��]=<��#�9�{�2��aS�^��X�L,Ҟɏ��_�O+���W�d]�T7��~x`=!ogV'���z�u��l�E����%Y�뮈�bʻG҆ �an��i�Fp�(Y�e�7}0�����}��v��=>����_=��X�+}�b�]�K3mԩZh�!]Z�`�M�Ξ��,�	��G,����Qw'�A�A�\�u�:ߪB�咶���8-�0���.h/��kgp��G_����_f�n;���0��	 ��擹�BbɄ��pЋ�F�׷�z�K��^��v���7�K;��AL�?��!�������;t�4�[�l�`�g�N�MzW�T {K�����2��wj��K�#�+8�M�"��,�.��-5�����<������>��%{�,��`5��!F��l��u�D�և�3]�6�������Ue< ��'��^�F�t���+3(|��T���c�Œs�p���Y�/�8�X�@j��,�O,�_m7���3ֹ{����b�8��Fￅ�N����m��Z����>��A����(�<x�v;w��Я6��)
�LB��i�
Q��5�j�v�p�yxmy:/p1�N��<��O��N$������D����ȡ�������1�`�o�3�A83�ޛ�A��YsF�rM�cX����C��2�͒��{Doc���U��
�bP�?=A�Y���=u���i��jd{_�� ���%W�;E�P�83�Ͳ���|v[Y�+�/AG|�ڥ�(dL�]i��
��՗;�i5��Y�p;�^u��.�f�pw%3������*S�_�Ϙ�� !�^J��<�,8�)'Q�i�?#�\t�Yv�a��b��-(:��:l���E,�{%�z�Cx��}�v���^��)�n˸qoT�2��nvt��[Ѳ}Q o;t���
��,�٣� �1��Gc�ݻ�JQ��uS�e���N �{�5���憩9����z2G� ��(�z�bet�%#�S,��J̩c��T�sQ~��q,|�?z@�쎙DG	��-ḥ̂�b�m��>�&�BX5s��͠f�.�7b_=��@��j˂� ���%e[��6��Y1&Xuо� �+�«�f�����w_z?��>h�4��6�0���W�ԅ��މ\C�{*�� ⾗@g���?9�GW!>�;\�~s�@���W��'�L�Qyӫ��&��-*�<�~7�}'�
: ��虎ӿ r�k�'oD��[�6b���V"-K�.�9ĈN�������Z���Zkɭ��t�|Pf�����O��(ު�}�A\!��!���]�^���2�G4�h(�3+&��Q4����wz܋��;ؘ}a�$ `��Ƀ7���/h��y�V���f$gH;��7���{��Q��7��R�h��0�&�`L~�YG�sUFs���:�������Ö�`R[��E�(�H��`4q��8��uM�8�	�y�D�Im w�1in#¯�c�K0)��U>f.ؑ�B:Ve�L�fZ�-
�ׇeT����� �">����w�IF�
�3�py:ڪ�cS�?%�C��ROMnpқ��
�`C�zT�\��%#)p�Fb�uU��s=�k��;%&�)p���n���财�ס���lS-�@1	����/�]�
��G�Uz��g�~[�F���!�Үqڗ�uRt�A7��dA �#�:�i��2�=Ⱦ�+[324��tY�1?̵t	�J<�FO�=��-�^9���~���8�����AO���L�~h�T�zr��3%�G�?{^=.���)ӊr� ��f��� �Z@�AL�7 S���p�2>r)��+�o��tL��\g�Z�����D�'#��a���25��=4�,h!�s�g���'�K��������+���=��[T9����b���/��i�hq7\�%��t���əL�I�hX`����b�{���KKh5y�=*�#��t���0oP%b�P��Bm��13[o��t���G������>�d�����k+���=��޿�d
��+��<e@�<���,Y
�&�����HY��|�f(�7��`��?����H��{��>�OZ�JU��[kIَS���P����p���v,+�����G��] 8�S�fٓ��M�����a��VBza����#ؠ�t��諻�7� A3D���o������կ���9���"�]�b�q={o|0D�6��Kt������g�;�^#�"��˘�&]�}�B%��j�	ހ�>����	��~J|��dl��hϚ^V�fC�
�/�%�ݝ��Y�&��zH�ɐ|�� Oh���<\���Tn�L�{�M%c:�^ƈ�D/�?&{���&����3Y_��HGɻ�C֍T���Q��zD��^m0F��$������7-�A$�{�3�I�$��#����3׬��tc�	Wy�3���J˚�y,1�ƛ�0�'�:��143��ה?��5��8���XeO�*).�=�����8*o�S���K*'�z�,���;=�F�A,W���á������3Z%�Z��d=od�QsǛ�vfDu��ܩ	H��z	�p��p�ܞ0���S�Ki�89E���䶴Q������
�w���-l~�m��py+�x����B�R���5b#�S��b�s������x�,b��D�fu���U��l����l��^l�R��6���칯/�3�������S������H�K�k'�ʋ<_�-�c"��ѡq>$��iW��"�v0`���l��]{⪜�йS�V���x�+�7:�u�c��.(&É��]IE� ��g����l*s�_`{#���B~xL��Cm����8�_���+:o��7����P0���	�9��M�+�3��U
k
9�9�o�?��}�Ҙ���¥��J�O�ܛq�KE��i��:5�蛴A��5��'f�֕�j� OB]\��;����V$�g����fC{�c꬀mE}`�Y#�&�2͒��GZ���U��ۺm��v�q�&1U�o�	l��QyoP����}J������L�WwDʨ�����\��	�ǃ[�ep��Î����l�us.�%����ho�~{�ܗڃN�2J�X�jvaT9�T���EM����E�����`3��9]S��-��|�Lj`Q�"��w1��d;��f /��58Q�FC5i>��}>����{�L1<��F���C��ή����[0<�ƪ�� i鍞�Af�T��"7c	�TK��J��Sv��=����0�
;#la�٣*4e{8S�
�BljϏ��!n'Ǧ���A�^�	PXi�xv��n�˕���U��E��_��d+-�@(G�5P ~��=��CՀ��"��t� Y�g���|MKh�*�!gM�k=.��[�<wzʏ�������nˏ�+qN՝b����p����PR�ۆ�G��aGP��H���Y�}�KF<}���9kĭ�h�V�\��9�KI��[�1`@�0C���Ј`x*�1�˫	�_2��}����PǼwY�.	��ı7"O0���C�x�I1�\�10��i�Z�ARN�A��ؠ������Z�2Uk��A���ѓ�#��X�|��t���}Rڱq����E����BU�Mg�H��L��+�Rc>;���l��C�&4<0J~C��tA:��O�v�y���ҕg�Y9a�K�-X;|ew�	��Kƣ���j'��hb�!_Q�T��`W�qe�62 ��V��g������)�(4�g��y;�s<�
򯾞�<���K�{h=C y9�b:	�{cM�������Ot�M���o�":��7��^�ߤJ�;���<�2|������cE��.:&�@\e�m��No='2�$��ؠ��3+�U�?��D&Ɇ�S"8F�Y 訞���]O��؞�#�����"+r_��`�����XG��p��;��юhÅm��LXB�+�-��n��__v��-�<��|92;�A�G1]�f*���I�1=Y'$��#.*��U�Ԙ�}�86��p��Ђ���_S4�,�
�g+�T��RR!?u[L��ׅRF�G��+\��	�P�1	ez:����Ԥ�E�=Fo�,⊖���?H���7�̺2��v���4~G�Yj|�ߴ�N�=6#�����߁�N!�̱>�ؼ���C�%��^�Z��\���@�7��-9��ݿ�<g?	i��8�.��C�јO�nB��G�!����SC<�R����p�yޙ�W��"0Ǳ�d�]����t���O�H�c��4o}�A�<*
���8�x��P������1��j���w9xT35X8������,8�Y���[ �V����܀2�*�bf�F?.��+J�&�M�F�Sj����P_����Gb�`������:0����F ���=��
�7k���⴦�W�j$�qR|������w�[2,�mp�=j���\9��#��UG��=H�v>g�����;�H�EU(�D��ܨ˷�rzg�ڎ�se�ƽ�q���A��p(�L�g� ���%����D�O)���~��%����u��`�$�2�g }w����s&��c�Ƴ�������j)��K?yO0?�s6(� �9��?����!�[�ғ���W5Vr;��r�'�7�cm�*���W�ry��b[�����Mȸ.��Z��Y]�[�o*}c�i9��:�=2��@3�C^ūl������r��Y�UȒ�=�rh���6_엱�Q��C�N����ME�>���.�\)����[�}����Ǳ���;�*./�R�A�1��'�U� �%Pw.5Lg�o�K�e�p4����MS�}�k/�����6IhȀ����>���Z�1�!0t�ir�6�pk�)b{��,�qf
��B�G�S(���($�<��9�ɧ�@�D��徭���;�-�R���T���铎_[U5j��td�8N��S��&� 1�E����t�����R*7�]je���ًP�z����+�J+��̯- �ߝ[Kv���{(��d��g�.���o?4�	Z����D<��v$��!(%_	䟭/u�<mIh46�w��`��S��|���!_�~�Ɛ�=��I/\]^������0"5>�rɛ�^�E�����s��}O+�NK�a� �g����OZ�=bT�F��Qu���E��7��Ōj�ڨ�@�nQ�A����X��j���� �k١������]S��;J�۸"*�KMe_������e�^���&��ڹю"O� �iF���(^9 ��a�aѐ7�v.�����X�����iQT�6Z�i�p�x*_dl��3�QzhO`�n�;�wp�)��������n(^V�l�G|w��׸s��?~D]�����ȣO�`��s��ʦ$S�{�|6��d4�u�!:b��
�`���yn��B/ɣ[̴|+ x�gG��E��$���Y؀�Q����e'��6u�?s�Ԯ�;��ŵj1iG��b ����6�za*K��06�,��^�{�(�G���^�j���|�Wf��'�C��������X��?.�R�:�S���}�,�*Y��g�$�r�2���0S|����O˗�z����úA�^���Tx�]YX�:v� ����T�ȬC�;�����v�?I�`����N�!�x��A��|��b��6�W��Ҷ�ˢ��L�֠�|c�c�ަ��=�r�z3tg��哑l�.F�3g�>A�TS�\U���CA��eJ�)�*tx�x��-�+R?�łW��0dQ��m[Κuhc�g4&O7~gWD�O��T(NHk�]�(F�zah�m>K�J�)R�����T�C�d�Ď#a<6PL�UKx8%�i���k��m����I�U��������w��ȥ\�'� Q�p����Z��}��Ah��Vp��|~�SwN�KH��l����w���H��8}R:K
�u�|�`�.$y��9�6ޮ6RW��rw�����:7����>��w�}C8��x,❲M�bޱ�O\�,徫W��=��|�4\��L�[�(�� �e�d.+�au��l�|������	GhQ��i($�O`Z�&w��7VU(%)�P\	78[ �5n�&���#�(j�Gx[�b�B���e��>�E=ש�t'O,b���̙z}E���m�LgUǾ�p�o����;��O��I�w��uGy�H��+���P�2��l��������d9{u���Pim�~j��b�-Q?�Z��23�W�����mp%NK�������TK��(&�0j�x�RM�PD��G�ss�#��QRV��E��K���jm띤%-����Ld�;Glms��'�_��Κ�t���.y����Z5�Ҙ���L�ņ든��+Z^T�PW-0�Q����y��>8���N2�q~4:i��+�AA8��،�Q�3��{�u�in5�M�%6�P��-�۫tǲ��h0�t%=�~����k0�z@-�Ԝ>����^�	��~A������"v�5)�ID�.쥼f�Y@���ͪA>��B}D�޻��0�_�@��{������ �"i����,�;��SC�G\�e���C1ق&O��J�%�nU�SR���3�^�
H��?���V>��fvgLݩE�.�.��1]�/t
�yɵy�?Nbg��(j������
����=[�ݡ�Xe��?�E�v�f�?�P��;CB!J ����A��P�e�7Xz�}� |���%�3�G��J��қ�,�+�@YC?33:+�r����H?��ӈ�� S/�;PaF£�.=8�i�w�~���Y� x)��HE�#�/�E��!:��7��>σ���/*���EO��x F���K�+F�{�8�IZ��Ѿ���ժ�*����/u/qk~u-�UX�������`G���7�΃����B;B�����Q��J��[���w��
B�BceY��av���n���֝ht���UO�����ˍ��q�FH3�y`>��ɫQ=�EݯD�S/�5��u�G�V��,<s��1�t��BPgb`:v�?]y+1�^�:��x#����F���p�{���݌;�����\�0�_����8�>0�R�� \x��R�'L�^�2����������k|� ՛��r�(��BB��
f�9��g)���{�<:1{����������)(�y�72�2	%�9>�lΥ��9kr�$$�o0��S2B^�i9L�s�)r�}E5�}�ز���'�	�y��5^�4n�o�H�)B���k9���_
|B�{d���_������d�k~V��X�N�͇�,AF�j�ͺD�RR�/���f�'7��r�_8m1s+ݎ�Y�͠iR[邏��(m�	�M��=N�c������1���m۸(������گ���yH��a���.��(��}Ż���s�����J����8w��@?�$�G\�a8�x�`�B���*��kp�E4� ��К:E�^�=���3�/ʭ��#��>B��J���J���B��|_Xk��N���bQ�0�/�S�}g϶��s�ʖU��;��A�P�s��ơ�������Л�'�� 9Q	�����3`Щ��d��@�8sW�B�
��es"�|Q���ڟ�)�������ȅ�|��I���Oa������B@�V�J���܊��;��t�>�ِ������#U8�	���AԿ�ۀ��7�e�zЈ~��"(6����6z�����Y��'Q�%O��)�D����~n�h�[,�~���138��?�y���ը��֑��m'����j`�{�����\s�����y�JU�ܯ�,W�bJ�y��w(���O�,J�g��NS�p�7�I=���&���u�
e���!f���2c�/O>��4�q��y���>{~�$-P�ป�~O$?��$B�t�����R��{.�x�j��E��3؂���N~��L2���h|_���FRr����y�Pģ��r�O�r �e�=�=�& ���s!�*�-��	Է �2�d�g��aJ�9�\�=0����'�F��\�v�� ^�v�)��S��28a{1_,QU��
�!�����Y���ǲ7Wt��yp|��P���ݧ�5VȈ��'+Q�E!AQÌ��f� Q�vB�	3�����V�P(#�$^绂��֨+(��}��9{G��x�F\k4xLm��������� {�
�%Ż�1���Q��8)�n듣�.K�6
-�	C*a�B?,`�G+v�Ƅi|Wyz��U��u/�'Dx�|�t�h=�)��р�c&�	��m�^<��� q�=6�<���u�*�Oj �B�d��$���2]��z�a� 	�NT�o�+�^xi}drT��O����{p,t���e-1�O����~�lh5RͿ0j��O<*P���3e����rf���=���v����A�ʮ*f�h�XV%&]X�u~{D�����syKI�#���>���}������\c�m�B=��u�\���BCr�����<4�N���n�xX	���Q�9�z�?�6u@*�a�qg)f傁�,�2Pq��C'��r��rԾ,�%���d��IL�������M ��1b*�p�����{j�̮$����p��\n^F��GdpR^��9�h���WͽU�q���'���O�+�-�+�a*P��&co�8��[O��${�e��^�����b0N���e�C�w��(0�ض�!�j��T�I�3o&`�|��o�Ş\28�XT�����VW��<��`��u�׹m/�w�`W{���8,��pA�J��z���YL<o_|��"�7-�М֚�䉕6��%�5��P�e���E)D?�25[�� CCM.y���x�W���I�i"&�DJnw���q"�|�3�B�-Zb+�)����R�Yh`�H01�#����iy�y~V+�Z�p��sI4^Ki���\5�>k��L��	���~���o��5߱��VIZK�ē��8��@[�~TŢ�1��=q�BDi}�G�|���H��V��.56@rI�8��G-�)�j.	$��Ǹ�&,�cլ$vʣŘi)�9�(:��j��<:m��^����$\��}�H��\;)�Ty��\��L=���1��%,8�w��5�����4p̐��500�0_R�(#	3��n�rI��2_�>� �O��D?2��|tf���	Y;O�� ��P%�16�Iy�qQ�>��͂;a��G
�C#5���et��A5S19��q�C�� ��`�*�&��a8,{�}/06{��� �On�8����0�ˬ���-���1BAMH�z�J6��X5�m�{mg����R��ˑ�����ϰ}a�Rf���8\�G�� ���G#�v����L�NXǰ�z#=);�h{����ǩ3�
P $p�#��ɞ5��s�`b�\%g���k׷���Y��Z��(�G\
�؏��2���ݜ象�.S�)8�.: �[ڟj����4���A&H\��uܸ�]i%�AJ�]��g�;�mO�P�I $�c(��į��2��?|�9=��\��`z��ID�����Yv���O~J��NK�����C}r��@���^*ف�4lE�`|���; ��6�׳cR���Vl�H�@AH�Y�&A/!�Y�d�ya��l�*�ky��nZ�	��֌�O���89���̐�������o�"�S�����3f&L?������-�zd)���o|�Ha.�Z����Ҹ���3[��AN$�.�.��_\A��$��B�ۣ�&ĩTV�F�DG4]����9��<��R0J._�&�>�D�Mz��������}˶({�W]a��Ȗ�sDB��A���l�]pѐ� 9�w
P*3��3�5v&p��0�̚��*(����T0��e f��ܷ6S�Z��C�D5��p�Pl�qz�M��@.��?�X�>�r�>���/��eه�5���r��ށn�����F���2Ofځ\y�T�Ԩ�x鰳#�X~Z��s����(�Z�|��f?}:��) ֚z$���}�YF#�U��]���*i��0��G��s��P�}2��~�������v�2�O�q(-��%>�.�>|:������6�������y�PB�*�����mXsk�s�>�5<v�2�I݇	-O�����j�)���Ǭ���O��o���r��D@}	�'	��c�݃U_'�Vc�)�t� �Pf��4�_�>�,%�,j�������P���yr�����.�@ʚ�D ��U���x%,����Y=&	2w�C����<����}r1�(�*�r^H�=�\x�M_����H�Կƴjg~j1pqW9Q�����Y������}���f�D߮�D!�Mw$ʅ��l�i�+�H�"qXEF�;���ϛoՉ�q3��iL4+�@�%{ Ǻ�"ER�Y�M&S!�	�>���U{{wM�':�B��N�_Pjl�*w��.�k-2��S���Y��[�и�Εf�4k�P^�BJ�ĎL��/L���Ճ��<6 ���v$T�aר=u��{����LE�[�B�hy�$��v���zXb��ʽ\�'np��X4>�P�r��Օm{e����֔��U�<?	��F���z��#�c@��_m� ڹH%X^|]S��.�rF� Hy�Y�&4��Q���������p ���HN�3:��JK�C�5��4�&� )�9ŗ���v�>j^|'*C��q�e?�g�ʻX��էL �&]�Y6p.�������nxͨi�y�>��<�ꃠ�M�ac9&�BK�pMj	��w�P�k��ζb��Ws�\D�/{������𘮽����p��m�eZ0�����0�~�T���q�n��_�I��2���m��� uo���;L@}���Z
�}�h&j�~�=՘�|��C���Ē��;f��C�'���st1-�����W�n$�E �+������2��о����[��I��A��h��r)�ҪKO��HC�ɲ�@��t�!ʎ)�&NÄ\@c_��@y�/�<���?���ܗ/��V�Ӑ�i�ج�?sMB��H��s��g��2I�ee-��*�r
0p7cm��K@HF��c���,��Oc+��<�
��\,�(�Q+�_2����k+6@C���
.�t�F���K%�xk������=v��)wa�u����h �����EL�i	I������.�݌���	���|�2uQ.�-�]�����ҋbkԟ�<�'�F��E�1�$9�B3�uYX���!�UF����L^�,Q�e� �K,�"#�<�y���L�P�ӳe2��"]8}wc���#S�h�8��[�c�69���p�.��B�0�Z�X���k��\��ijPVlYj��a�|z���O�2���[���m���vyjm�Go���1'O(��������|;~��|)i=��w��H�?̵O	ob�b������ �T1���3�/��n�o�l<�0Q1����SʍZ�g�XH�ͷl���.��f��4V�7��r�؇w�9K�AZ��Y��̡�� ��J[��FO{�1`J���U8���'�G���[���e���тr�'R`[S�[�T�?�nJ���8�g�2V����eT�s�H'��=U{`�g|����4)�
���t��1���Ѫ�kVX�x����K���������nD���3%�)�r���_3E�4k�!]���ĸn�&>�O�<:�N�U2(��|�WObO}����{|��{W��Ei��}�U����G��C���B�3S8��>�����P��K{'T���;QD������ֹP������nrD��d�۫����K�D���_~����]ƒ�9$BS	Kk�4���Oa�`â4>��9�)(����3H�V㶎��N4��	��8]d�$�O��w0Ѐ�k?�9p�j�$�(nä�	w��d2�=�x�5Њ��EʿW�o��>H��2x�E�2�q���C8^�&��T���op�<x�����X���J*qM�d0�R��N�I��&[G
��lXH/��U���6���Z�4>�qM������б}]�����/cr	�ɢ�Ś�}����a����0��5����S������4c�+E���+��k$s�������OUAT��0|>���4�m�	˃��k���4��M3�]�{��U�弭���~���$�ͷ��~�F|��٩F�	i,�xl$�A;�-���d`NY�j��S��g^cX^����`����X���+޼Xf��~5�}�����<�)&�lx�g*g?R5F¥#�R`����
��C�$3��Nh{`���~_���*�:� �`��͈<{O��>�o��"��� ؇�^�α"yD�4}����W��o<Z;�1md7TR��tb�D,u��=�:���E�l���
d��֖l�ӶKar!�M� ����6s�}gDI�a�q��#/]_���2�$�-,���J9��xX~Z�+W�,Wc/�\�Jԣ��!VɅ�����>7+x��מ�������yG��Z!`��0���;�){����fu��N�Q5�{�4,������DQx�HMYfT���䉯<��ʀ�p���
�d����6$ށ��V�cӌ�ó�.a:7_Pir0Mj�"��~2�9�1Q'o�o��¯L�1�q�C�MI�ATB#8C8���[i����B�-j�C�H�5AKRc}���H�v^�7�B��ѓ�ǠF"�G��ݓ��|�|3�$�3 ǊB�ʽ�f���6,d���$���{�t�}5�s6�`��bv[=ƶ;�]��.��N�7����.Z���-�ɞ��Z���,Xǽ���*.�.��$O����v� �X�#_���n譔7S�5 dI��R.'���H���PW[����2j&��ռ'�n��{)T4ט2�x��˘�չEp^"�������k����:ՙ�	�]�>L��X��}���ſ��I���M+�4�S]H(��� �$��@���}�PwPv�����sg��~Ug6H���34��(	����e{$��n��hdE<����۱�#�IWj�I[1��?��~�]�ss���9�핒i<���A�9�]�/�C(���=.JVy��ۈ'����ex$*W���!���F��/r�K�G�g��9����-hz�Z���o��j��^��-�+��"9��9���G1��Z]�J.R#���Z Š�yȔ���`�.��C���u��m;��?,%k)���{���Ԡ�J�k������I82�b�5Mu(y�y��:���nǿ1�m�v�v��	�KS�ի�,5��&��Ń;霫�%Cʞِ�X^���|�٩���	ű$�@��m�8c�[��H�{eI&½�(c���0@�cn�TH> �u����GC��ޫ�S� !�R�� 1J��� �?w�8r�>�d�`��;���9�� �I|�j�L=;A-b��8�
͘ߦƺg+�7fx���BZ���N�ԭ�4�`�$=*�r��̶�?0=��m�q��y�s-�����Mk"N9޺*y����^��o�_�:AW�.��V8�������}�|˱�5����`�R����^b�ح�n�I͊5��ȃ�,����d�L�Q]+����n{{�E��[|�L�,���& <0�>	�"'��DS�[]c�nᅅ��V3�Jt�d�_�`G������ŏh{� �)48����,U%.��U�\2�k��3�d�s���_0�
�Q0��cX+�k
�7a�ά�gӥ3b���${��:;�M�ѻ?w<��p���HI-��L8���K��bZ%�ǘ�X�3��"dAط���7f�y�yŭL�/����8U6�u��p6���wv�Jh�Z���� d�~��6A�(��+���'��"'�y�� �_���V�ir9M}�Qu���P�'|�E4�ni�2�f���Q���fĠ8�.e��/���*-���!�}�F�hf��"��p4��X�B��ʔ��m^5�R1�Ա5�M�w��o�P�r`L7��R�d�C�(]��B&]��������*�V<�b��V�x�TT�ߨdݘ�,oayo�ۍ����V�8���0���5�O$��zʩ̵s��I4w5b��s�t��O
3��d2!�?Qjt�!�1u?�+�L[�0��u2���_�k�?'~�3��=�G�U��1��n��@$��ʘ|B�ֶ́��WbP��� (��5BRu4m0��wGz����\/W긑Q/��YE�x��d�O6�d�׹y� ~zr���j��5�ȳ�?������/{����@ֿ�Q�</�G�g�{�����8x��n�Ec&�;<WǗz��B�*&ƙ���H�&I�*w��V�l �����8��H:�~��'DioZo����O��B0���<�
z�����G����H����
�A���^�-��Smn��w�"�ǵʦWja��;�Ț�
ǁHw�}�����޴@�n�?`l���I���&��9��	:sݓ�JiI�F9F�^fD�x6���s?�D���dM�(u��'D6�4g�L�<\�X/�I:2O^��\'-�;�@_�H�T��Βk��r�yhQ� ��.^r��Ꝕ�I��6�,b�;pX�S�����:�P�c�c62��\�G�C6��|-�l=KTm4�(oj����W;�>���䖛�����A}������A2�0[.p+��◰<9׌���ٹ��A^.��ʾ�1��M���4|��Gs���_�\$��,L���=�\2L_�UoP�<�A�l�ȏ��K���xv<�ڱga��,��4X
��Zô�a�+�Y�T�9|餑�9bV�U�Zϼn6�e�S�P���JW ��Z�OfC���b��|Y^��m���^X���3��% ��{��Z�C5��{�#0��?= �de����iP okEΐ�O������FF{S_��������n�6�g`��]|��ܥ��.k�q(��vy�i�l�^.f��-�����_��bA��=��c��2�ީ��^S�����z��+�ΰ`>��\X��9*%�{1��^d(�o@K(zw)DB+�8tY�q�2;�=��������tb@`��'�n��P��>�p[K�뤚}Uz^�lT�b�-� �u�]����f���qYKF9aP�s��yJĽ�*>M_�x['m���y?�t^�yf2�][9��䳐N�2�	3��ljQ�/�գ���$=Ƭ[NM_�B\�3zO�g)�����!���?؜�o�h����e���7����<��c_��Z� �3 doᩜa3����2w��Y��js2x��	��!x]Sy�^˙y"�����<��b�^D�!f�Xm|Z{�ښ�ܟ�Os��+�4�:H��b�i���/=}�mO���ab�c!z��B�F2�c�].����,�9F��
��� +�
ݮ|���w��)���OA7�	�	������c���U=��=p�_;csF˲z����H���7�J�6�\^�/��]����';ڂ�`���7K�0�����	8�hS7�J�a,%�OR�x�MD��ʊu���7CP��;6��$ɋ*l���-�-l�C8�ӱ˝y��P*��f�麊Wd�.N>���r�N�C���z�C���n�-��F��p�����7��/5i�#����<"c�$ѧ�Q��J��' U��-1�9�I�r�i����T0�{��+�("���[5��+�we�5�(k�4e�D1T��s���!�o�6W/a M�٤n1�&�
��wG*�o%!��>G"����Y6V%�s��g?ג>U�����fݗ�,0٠+!|$)����c�����dt$[�RM���#ã"����r�l�vt�����А�x��t����	v�0�5z�F�{����-�6,K!]E
�Fr�"-��f/Q]o#�8�?,m���4q����Ӗ�#=ti\�Ć��0�1d֔-�y$)�ѹ\���(�Lu���Y�~��9�Z�����R�b	��r�c��`z�b���o�K,~`��$�	�R= �:�<%O+�c+���v 6�cR�G��U��[E;B��h!�,�ԥ�J��3��kTR`�4�=7�|�[�sA�C�3�یf�n�	A_G��ˍ��]|���h	����?��E�7�aFok%*ʅ�����.���Q����׀@r�L�H	3�&rL�rX�c��?h�6s+�gES?�F����Z�eϓ�C��R/��f%�E�l�|=��B�Q��T�r���Y��"aݥ���/!Ž�ꄩ��s�����҇��t�n�YX:>-�j{y��:�dk~�3}�&�S�`�|��g�4Vh�Q;]��w�����c;tшTk2���z��x0v�L�$b}�F	/���gg��s`)�5�Ƚ$��j��)5��;y���Q�^!a�Sm;z���O�����I��=�9�j9OZej���g�;�3��9�cg��@[m,@ϻ���"��շ�,I}绬r�9U�x-�
�l�b|����k���^�p�핡V��网�5�L��,o{i|vt�+9:�q��J����ȯWm�M���/l����
څ��l�6��D�7r�h�������pW�@�=<�k�$�:��ٝ�'Ѻ�r�0$ö��Oy�������+n���r�ͷ_Q@�f?h*=	���辕�Y����X�t�;:G�@�@be��El��tҶ�����뙤
�����k�6/wt?���h�V�e�܋ZȘ���� �k�Ź�U8��ԇ{&ki���{�r#%��RD}�a�u�$:k2���h�o���˶�n�A��펣�����T���S�(��-����I{�s@�be�z��S�<F̧�2A�N�v�������M�+E3��aQ6��g>�����+S��fyk��>�~�Ar�x\�.��\�*y���O�&�y6��gL�ݼ��P��p~�EZi�枴|!�a��ma���)�vt�'Fv�~.�XV�A�
&�9��W�.��!cDE��vi,�R�7E�+U�;B��';,>vm	�UQ=�:�Rфnc�$q����M]����ĝBy��(�Z��/5����X�)1�z}`OƃA���۫5������Z-Ϗ�g7Ŀ��#Ȁ�l���
#��}(S�Bt�=���1����1�y�1��m=MG	 ��������utvg�u�����9�����NY�ϐZZ�*Oȃ�ܦ_J*5�L}[8B�m����5k¯6�l�ie�"o��Z����:"�)�-y	���3o��s��!1l���(�zX�^�A@�_9S(��|Rg؊G :�������+�OU�M�o.��4�$y�Sߏ2l�@P=#��$Ǘ�)�ݬ_[��O���υ͏���H��(��(�����g�1(sл��/a>�\��;^I�K�d;��V?�q̎ar��h��08��!j���<��>��6�ƭ5F�<�VC���P+o�����+��#?�Պ�c�9���-��]%�W��?��_��Z�,{����&�'�I	* ��R�T��$���)I%�u`_�&����[����r�?��B(o`��)*�p��L~�Fƿ���>8m4j���=g�7��<Gd�
�<=��j��{kΑ�utc�茆p~�)�/������ŎO6C ߲c̩z��g�&!v��ͩt����{�
����X���vX��*��4��vG�$*nt]/h��mX^���Ŭ��s�AP7z[r�ճx�9m�'�h��;�ak �G�d�%ꅐv)g��F��"�m���$���jp������Y���9�k��چ99����N��F]C1�Ɔ	ii����;�?��Qʢ0���O�������<�}�ٺߌ�RhB/_���V0 �B�I�� ��n��v~V�^��Z�
����9�� V&EO��Ec
$iO'��x����"Q��J�)%��Ym�y��)�E-�p��4���1�>���_�4'PKu���k�#U�P� �y1�=�^�l�����y)(�/�&�f�&3 S�/a)�C�g�$�m�i�l�4%N6�l:��m�(
n�|>9���߅'@�����bC��L��������♽��8�fl�?4���!JG��S�0J1"���֖���>?��;��N?�(�ּ^�Ìn����?����6ӕ�q��bH$�a��ֻA?03(gx��{ӧ }!���_��D���u�M3��E�&k�a��PP�D@�n��%��uT��ؽ��e�We1�o���se����4;�P(�gk��S�m	�jR�@�❠ڻ�|�-� �g��ȼ��_#q^�6�!�٣{����bv/9��ұ凡�$�ra����D>�%YD��ﰨ�OR��;�DM�����	aڑ�#Z+�_Ws\ء�4'*��AnMٱ2��!hI��A�KΩ����5#� �*�=I;�f�8�LB
*��=4y��)A�^䶖���i��4�u���TF���`�%e@�;4�E�����S* �\�	*��|���x����8�}���D��>�ιur|4l�q���$ٗa��um�2�!O�@�|X���so�3M'�8/���?m�f��F;�3���9��.�>��UK���Ͷ��pZQ0���c�sh�E�h�%#���T�<ŲsMژ׀�R�������/�=ן9�#�H��_��*�҂��9:>N�\+̝yl��%�=.YI ���ǖ�AΧg��"6��i��]'
7zk�*��H�&���iu�"�냦P�����bVI������b��,�ē���'ܵ�?1c�ܥ�!k��gF��C	de��^�t�A��L*Y;%�?�;���]+�m:=�Nr�KFC�G#)��m?��~��Z����I<a�=��8���iCLW�r�<֞�jbkq�\�:�A.T�WU��#6
)���┾;0)��8	��җ7�eS�����uԂ����I�d]*��Ly�iܭ��H8�``1#V`3go�-�})f�AL?80ޙ�A���k��}�R����:���i�AUh��#KD�}~_�B�ԒIc�n,�F��ס0��Lmk�iNl��Y�w=4���8��D�!J*�����+ڝ
�`*�a����	?����d`ʨ�2�Cjh�[znc�6�ȷw�Y�YG�,�K��9��m����@]rΦ���j���(�'P1�K��d�W���ջI	9��8��/`���Ɩ�	�쟷���{3�NdG�A�Y,7��^��V����'�Y��Ny>��T��UZ�U�fHio�JG�7�8W� H�s�P�4��fGv�v�pH*7*�)\K��i?C_���rx���	�h^I�3�!���i��Or�ϙ��[�RM)/�p��Q���<۵�{a r�x��/�v�)g(�+}�� l��>��C�-�`�͚���Qsc�i�W�4�}Qu�(]4.P��Oa�krmWi"�1yp>o1��Yo�4J0B ��g$e����!��s�m-BF`��CM�h�m�����i�;Y��[ѩ�['MN��[[d�O;J��M�܆�|"[��A�G�E����A�$+p����1N�	�u�[�8�pz~!��Y1ཐb.�3j�C��6�ne��D�μ}�]�~����0]������f�	�������P} �r��*f%.���4!i��O$(Y~abI�L[�ja& ���Qt){�7Æ�{���� ���/�oj���)�η���ˎ(��O���ִ�m�EgH�y]�\<'K���%Q"�&8������Ѓ<�����ZR�P��߮V�+Z��T,k*�|�T�%\��	�6��R/����?&���fu�-���(�	�;妚_A���^F(����V��	�W�Y��X�\��5�9�mk;`�aq� ��6C$j�7�����)Ǻ��HݛOw#(�j�h�y��%O;2�9`FX!�o����Kj���5���.��>���3�(-J7F��-��17���<�)�����j!��v��*�B�����1�+^UQ���r��y|7
TL�b_ �}p[w�(���*a����fV�9��f{芼�5~7��`*c�J�h���[�U��O����� *#fhYsbެ]�/ڒ��q�+�Ǯ�X��6�t�+�\�a��-�n�W�f�D�!� A=���"ŘL���靠�U� ]��-=M4[��{�QSQ"�*)�'΅���z�����e�l߮8�oT���x)�=C{q-L����BĊVEȠ�-]��7��]����W�a�}S��@,I.�Vokq��%�m����7����@[�ǚ�um����eҍҴZ�#�|��)]�y�5`��פ?'��d�[���M�듂ݥ5q��\�vNzL&�t(�a���TC��Ƕ�ԛ9#{����a�Di��y�iy��s��/Ai�����=��(���^#S��br��h������a�⿥�G���L�������H9e�m�Q�~�^b�zn�1֙�����f��ƨ4��Cĺ�BLO'2��������=�J+��`R�(h13qɇ*}ϴs�e��o�`�K���}l/������f{=����Y0���*C�>�h�X�,˰���|͙BV�r~a�db�+��'^�72�C�2#s���54��f|O��{����^�p<U��d��`X�m�֜�T���հ�6L� V�d�z*�b���.�h�ל�u�7(� �����QW�"�q�ͯ)]W]��Ӧ�X�g��6�3��{��X�t��E~V�����Rʋ�Vl�>ʐ(� 8��>�&�"���Yas-�~��}�nۖ�IWR�ZV�{<��� ��,�c.������x���.X�Q��Ht�U;8�0�-��F�Cqw}C��/�����E��h�J�@j��V�] yc�mv@ݎ��OL�N}��ܭW�N����BgIM�p͈�0�g3�^�B&�w��T�:6A>he˰L�3��8��B�z��L.�OT����.t��6?�Q�.�e�t&;W�z Ҕ.6�f�@�<y�b'v�`#v��M�k�~��0�X/{q�
S)C��k��0�?S'T��dע�ՀƁK����y.(�*�
��μ��u�N���=���k3�d��}�u[4vU.���{�b��P(�z43�ebgӶ�3���0�>���B5q3o�K�d��dJe������cҳA%43���)������Dҹ!/���>[�����������떻��D(\��"]6�m2Yq�䨫�� ��tN��P	�o̔'S���U���_�O.`W�&�b<�c��z=�]���a�����f}�)c������� `���6�`N=��F)F#�ⶸ9S��-���A��[�����ڠ��TA�����Z�LK,-,w:F� F��JM�O����<�w�Z��*3�ߍ��-|��U�J�� K���_څ;�+�
�tby�v0���S'Q�^��m.��z�ۡ`[*�	����6S�_��Ⱦ"%(��@���ۯ�Q+�mn������ �C΁QQ�z�������oӠ�A�����jܖs��w?����+Y4�ԕ��"_]��D�����1�Y�Vf��h�`-5��%8����Q̛��'ͧ�������_Kv?��
�PÒ�*
O��b�b���]�Y�8Ξ��3�\�'3~م�֌6��_�n��M\S�3Q�4���+&~J���O����'}p�#�\\a�a����l�{D�t�!Yx��;�ӣR{�n�Q�ΝfS/������O�>�~f��6Eޝ�O��aG�u^1Զ��}�#���>�F���6��%�V�+)�e��� Ә�Ѣ���j�p����Hwc1���J�As	h˟�EAҮ h�����٨=�(7�r�z^�<�Vz�LƯ�o������-&�D.[�Cm�Ȏ�xL`�F;��dO/��-�����xq����S���-��Y�U�bh�KK*����ַ��2m4	���ׅM�G+?S�?��rC��^��䩻f>C�	T=ʃbW2������Ս��!ڃmf��ʃ8��HH)˳��!���1�M5U�\z fp���ƽ�GbcM�OuS�eœ�H�B1�E����W��H��`+�ʹ�9�|0�.F".��I����u�{zS���m�?)U;�e��w*���zy���+�
WJa�t��|X�n��'�;\x�}9�H�e�N��w�����P�҃9�_{�O�B���9ĊA����-��$�t煙���;S��F�&�� ��x{X�{׬9�2��:�2O���ް%�s.�+����j<7TV����T�2~�Vk���S*g�~���3$ߒ�A�wV&4�����,�B�2��I3���G�e"�6.@�N���NH��`�N�1�W���u��̷��}� �jk ��e�[�Zi�E�;P��;?)�a�8rDg<Ny�t(� ��$�X9�7�� �'�+	c�'�V�j�شڳ�����IoZ�˃Z�����d{J^�����ND�Ӹ�����Ձ�p���2Aa��������� ����}3�UѹvCG<<ƶ0��䫞{@�W-�ם<'e�"��6�18�?:��'������J�>�ʙ%���)1��Yp;m7�^"��#'K7�������}��^���$�̜��8V�ws�}|�s��P��8��P��!��D�'V��ߗtβ��MH+���z����Q �`j"�Q��E��D����#���o���s��EV����k�Ŵe����΀
����&
@V�FSm*%� ���݈'8���?��)��[z���@��Qy�NG��F�?S8]]�@H��Ծ�>.��k��Y����J��ڦ����$�~p!�r@(ʘ�q�h�҉�کC�,�,��P�<|5h~x�.PQ�S������2�ޓ��B�}R�:�����Q�:��!�WXQ����&�3�1��N���-��e�#pm�7a?\�Q��Nh8�0�و�3J)��]g<�R-s/�Y�Ǟ��T�(ķ���Aw���Pm,K�������ij&x�J�{�72վp����=p�>�n����O�v�)�T�(�ilʀ��>�q��jÑ�uu��Ҿswr����I#�)`o}�ݻ��l�֡�̣J=��0>	���r-,@M��p�h��Dn�o��>�Y������a��0d��#�Rv���E%�|p��1n��D��#̊���)]��W�͎,q�f:���x�k��R��N�r�]���3T6��[MXvO
]�7ry��#������:���7
R���ScNV>�A��T�p���4�Ӡ�X��/�047��d���:����@�衘��,aJ�Ǝ�5�$u�mYװ`���E���ɸ���p~�MyC*����)=P��M$(�B"9���~�-�kXs���D>g�u���H�*��Z�����&UNz;iK,��9���Q3�I��(5�0�#�`�x��Z=g ]�@K?���̻�r�5x��m�I"�6N�(�6�x�иq�ī�ϔ�ra�]:������c���9�2�x��,$J/';Ґ#&��׃� �|rԾ=�F�cMf��[+`w>��䔭#�2B�6v�H/�Oj=��%&0����*{����!�C��U���6���OD�c6� �3u�^*H��.�|���:�hl"���2��h��
�����<�s���BC��)R��5���eD��w���9�ZG�`��3r[l��sОט��2�!0�Al�_�	���m�F�I9ѧ�p��fѪ�ȯ>���n)�m��ѯw�;�v�W;,2m����xJ�o�
*�	�b8���'�]���$(O͋y��6n�y�\"d��yZDLex�n�	����"�����-$�{�Y(c���@�0����g���0��	s�<Nc�[���C��Nm��G {��*s�6/�����������1��
"jv��eb�MP���L�����)A�>Z"r�]��f���JDY+f�t �G�F�!��4�gy�Ⱥ�����l�,nL��V*���ۍ�|���$���כ����*IfdpN� @y�{��n�}se�������t3QIO����:e��uJU�l��]��)V{��)H�s\-��*'<��jO�e����M���4<h��Z�g��&_��Պ�Ƿ�)��)�4�~w/d
>����=���Pj���bHi�NN�j��������Vf	֗�D~g�J���J��}�,C���?���1']z��*)B��TV�3d�岞�N��h�(�X���	c�= $NJg�仡eQ��?�O��[���G(��(��eb�@�O5��"�=�}Pi�����έ�	nR�%d�q�+�D�QB�.<:İ}DͣX�6SE1[F=!����B��3�b$ܘ���mw�E�i�I�#y�O'���tv"8�]v�{�qHh��Ť<0�n`�=H[��sSj��2���sh$)�P)9_�iO��L�,����>���m�+���l�$H�:�c����`�q��>�[c��YO�f�:��7�:�}�c�i����p �E� {ⴜF���ja���WlÈ�i�So&L$�:z��BV� ��c�h��;�0��tE���}���'� 6L� 6���N�
�0�{�}�t4�w�՚43hn��g_j4�F5e�,oOL�������S 
˾r�m�!�g{�7ƥ7��D]	9��c�`; �HU� ��g�t4��F ��s�H@0,����^��i}!X���z��ȹ�:�b�
ҝ*8d.]�:�S��O����0>y�� Im?:�S�!���F�EM)�mlgO�{��{�+}Re�wxu��Kx�;K�u�6Gd�/�e��"*B:M���Qg�[��am�@B�!������v�ݨ�jU `����W�� �e�a�V�Q�n_Ӂ�X"��c������;lc���B"�W���������������;aO��t�*{<k�2��F�To��RVc��~�xzG���DR��,���O��_�Lz���K~ܑ�,_W��7{��P��˜�������5a��k�)Go˚�;�������6m2���I�3�����0˩��2���"61��*��r!%��=p��1�F�-���i���^�%��k%-L��	]��m"u[q��Ofݱ��?�K�k���3��*�{e_$U�;��oA����y�	s��{_	-���x�=�i� ����I#$�$N2�/9�vG�����/@`j'�W+ Kb�I�K��T�N������`�]���W�i*jM��8L�v	>FT��̊*����;9	�h�A���<|�*����u��np.y�N�l��^|]�Qp�u[S�6���SJ�����wh L$E��+W�g�.�����
qh���Dt��Re1������0��٢�7�76�Ok��M>���Ԁ����+h�#Oy�ӽ���8��=e$�p��� ���Y�<�i�P�������.N���ʵH۟�u��ж-,�����/G��#�jW��x �p�٤>���w�^'���͋f&�����VE��v���flY��q�#+�c������v�B%~�� �c�m�,nO}�Ist�.�5H*'�T�e�0O��g1ml���*�Z_H ��H�&ֱ���B��>�O�W�Q/��R�Fո���ٿ�[f@� 1���5<,OE��G�����3���2>����eI�*	��D5oZ]+���ۍ�t���8���ӎ�S��e�'/ �Z�?`�'va��s���	�G���w�;?����v�ކƌ��`KB���A���W:�H�+�[��d=n$�j��;X����Ϸf��^�=(.��c����Z'��R����L=UޗD�Z}��tX񡷸n���?�fwr7��Vc*aM��e9�����Z%�Ѳ)�$��y\f���/�	�RăwKG�.�q�����>����`�%�";�����}��D�F����*C�>
�[X�M� ��\,Jj��O5�����mh�gT 51~�����R�"v�1�j�Z�����mM=%R���f���+��DP�2���jP%�ސ�ku��#����;G�`㱘\��\�(̱�a��~�g��a��L�Ns�^v�b(���A�Q%��0�#�g}p<����7���wjZ�V܋J}�GP�0��|�@$*�������z�P�"�mN\�@�W#!�u"�D����'�*�?.*j@��0d�yd�-�$�z,<��2˥���a��x�Ӂ��Y���B���e�A���-�L?��Y6D1��:�P�fj���bǏ��t��1}�|���e0ͼ%�^�"J)Uɧ��m��|Z�D2X�΄�t��W���y��9WTzi��O��(žf �����K:RK�YFlZP~W�M�׾8dU�af�"NHxO��j�/
f��#$sPћ�[;f����~m���Q����V{��}x�;<y�-g�,aی����A\�n�#VLy�_��t�=�zT	lE��Ɍ���d��C)�@Sڮ�V����Xn�O_o��uA�w$��p	j��۽dǫ��2q_<sF�D�CJ�5��Y`X�g�8�>X���]wLE�@ U�N���J����rg�ET��b��AC	m��0�EOћ� ����G~$-d���HGn��, *�9�{jN��h�/�GYk�v�G���V&�c׎��RxV��1g� �6ɻ��W��tMX]��?Hu���\l��%�a�՚
�=�]�}0hO�Z2 ���.A�~�}��!ck�c�*�x�T}>����������/��_h�)�*u=�	ސ)� "<h��5�������J�T�lCU�4���)��5�6��cOY�9jU��C3�J:k��v���c����3�d�
e�_�;Gx��Z�b���@h�W2���<Tś&����Ɗd���~�٘PO1z���MP&j��8H�4&p����qJ,(̪��Ё�GtM���J_�D�G.�QL��7�J�Ǘ=�K��<�?���V�rY��̱���v蘒�1��U��?��"�ˍfa���^ּ�K�-�N1����^�D�ab��k5���H�� �jߓ��S�5Q	E2'���������oj瀋?p��2U��I��/��o�`l��f�4z��mr����-k-��H�ҽ�;"�C[c]kzln��m�ŷ�EU�����>�ζ�, c3�oN�p��;��û�#{�k��hqr��!gI�"�U�FvV����-�;c�?���l� V�'�%���pt�c�W٬Ӆ��~�O�<�c������E���XB�P�����>[�l����@O�jp[����mW���^���3}���+��f�&���!jɖ��1@3���V�aKs�$��l�I�w�����?׎�'!�����B�U�ك|{k�j��w\���ԋ�NN(�c���N�;��7G<�L.�M�b����`KB��J��!-�$u�߇�&�Dd%�5M�я��J�oTj�#eӎ;N���I���]6�3nN^L�a��'g�������8&j`'M�87|>�|f��2z�g�i��]u<8 `w�Z�)ڐ1ݭ�\{^So��h��	�^��ȱBA]��=�x<!��I+ϰ$�>A'[[H��O���K}�xʎ>I�*��M��:����� YD����p���/X-�����Q>���{�#I���K4w�N�o���vb�-���c׷�vJ	[ ^ֿ�HzJ_a�R���H	�xH�D�z���b��h��֘4�ޅ�Q�J�[�e�(u;_D�c�o�{D|�΅�IeΣi��4�,�8�-���#�:"�y�`���o��ߢ����ׯ�������Fx��a���8��D[녋� !�TQ^M@nw�Ov��3tӅc�RJ��/M	 z9E�$ٻ]@�@)���;G�JqM�V�t�pt��g ��wt�[c�x��d��3�}�`���S1�#�:���|���+}>
.V�Wk��8�V����}[ �'�lX������Zt�3�e)�ch���#��	��,�j���zp�:[���u���]�9���\xs%�e��ޛ����ź��1(��~W�(ɢ7����Z��5���(��甋z��ACS��9:){%���&[x=e��6����)��Z!Z^�67a�\\&�������go��g�1��Ϋ	ѻcT*�*����O���[�tzj�f��X)x������s�cYHg���r�FiL�b�v����F�y��'v���HM���v�v��LN��v�0�%����T�c��ZL�#L�	�C< ����AH�M�$Q���ǘ�6��ꬓ�҃Jv�ç1���lO5�@)9
����?��!e	�5��F<��Z�3,(�����w{j>:Vs�T��3Q��{�t3�"�3	?xC��,��AX��UKb	�0aL�q"k��.��R��^�p�;4*���x4&��:B��g�#ίL3g~p�����R(���bLh�K~���lN�����%��(1_����mfr��{1A� 9kt�y�؎-r3�W4Q�xb�������u�kH��_������gVQd���/�lЖ�Y��Ƃ��j&����X(.�x7�P� �+��a�Y
6�w�D+�x��K�i�Z�f�ʛ�aӥT7�^�Y���"���~`V��EW��Hg��)�w�)i�ޙg,�N�V$� ��r�N�S98�~�j������%{S��z�4�@3+?U���㥟�QY�*JƛS�v�G���:܄-Uu�Cn;��Ժ<6B�"���CIZ�����Si
�6Y¡1�8*^�R�ms��\`zo0cˇ˙~q��
���73�`����*;�b��c>�̞Aeҕ#���z;]�g,����HT(Sޖ�i�B_6�!�Z�\�~7��ܽ��T�4>���h*�� ר�R���z��<~�lJ�p��v����Cl�'vPѯy�8<B�S��ܑ���)�5�S�v� H�*���N�Ŏiƭpc�D�b�@+��pˎ>��5���1��c^\48�㲘-a�Ӎ��`��{Y�č�j��k����[����@��Q���f5�D�=�%uB=A-�����|��BGHϻ*vL��B���ѿ�B��ܸzdv�^�� �x�3��0D"��[;���,��I�w^���|g������9]�}��$�1o��h��B��ه���f# C;Y���$y P(0
�]-�X5>�P&���jR)�[����V���H�	���Nq�'��F�}�#��j�^>�_ sM(����y�0�;���l�x���U12���A�Ŀ�����9D*:+0+ͺ���X�*�\�g��Y���Rn6��8S��b����wp%�*��,�B�f���<�a]�&dZ�Nm!'�����f
��OJ��>51m��v��P�q�5�2��3�b>��9�� �-d/TSc�E]Ŝ�����Ra�e�lq����g/n�g�(ze�j�(�����7k�=z�s�,�����	\l���ӡ�6��s�W(�������{�9k���^�_"�]I�����]f�e|����x��uх���{4���q��:8D%�yb4xU5D?lS�7�E{Q_^ʍ��6X�33��@�������N{;�����ܧ,��j�$d�4C|�����5��B8*u����z��?�ţ���5�h��#�ǩ <��thX�m�t�/ev�l����b憱�~{����4�E�r+�o�2�*@�����{_gm�J�ͣ�]v�"'5{�[0�,-��WAWs�ߜ�;��-�K��ġ�LCzgp�ܧHG���Q2��%Wi.ϯ�N`[�b�E2���E	Ҹ�FY�Jngp�Am��Atn��+6��C�c��:C��z�y��\u�"߃n��R$\���Ur����;SЈ�����wG�dD��P�4�� o���ԁ
��]��u���*���w]���r�Q�®
0�P���<WسbG#���l��w�o�,��h��yv�_~���aEYٲ��3I9��Wn�;�\ī�@�1H��Ixb����A+�,U�Kא���С����d��w��u�����T�D�[���XZH�Q��̝��n�}�'��sI���jϤ��!(�c��T�Y��^o�f�Fjp{�9_G���j�{9�[�H�����%�e~Yꥡ��2�X����Wp	L��~�hN�I-��hRș�n����"�֌x�O�#L'�-{?3^��TÙ��Y!��pY)���3b|����I}�H�I��q��#JXR�N�̗���������e�'�{�j ���@;���s��ק:Қ6�L+�#�}�u/��f˷�����S�!�-�\�]տ�����o�8�گ7Yn���`����e��2G$�:����&�ҼBߎ6R�< �vP럤�./`���Iu)a�Ui��F��|�]��E �Ϻ�� �m�lМp�s�q�)P�sE4&H�����|��P��boH�񍔉z� ��Q���P�jHNP�U�y����� x��=�����P�
��� C�Q���5p#����D5�ƶ*<z|)�
`>��lLPM~4E���+�A4�4������(0��&��2��Ǧ�X����i�d���f���N[&-���b�C\�y�/�i��u+O�^��$Z�SQ�	3�xlpl��Ȯ@��P�|cj[[��k��.*�q�@���#��>�R9�ӧ����1T]���|���ڽͦ-��3��2��)]꩞�"-P�@�0�3�~��H�J�J��M`��� �BV_�nRG��f�_Y��ZmvR�R�T�P/�'bx���L��݃�q,�{�:��'E�iG:��g����R$ȕ�ҝ��}������4}S�v���~@���ج7�i���~\*��?����W����T�Zr㡂xHN�l��N&��ֆ�����Zߌ�2��@��
���]E��E���{�Xmjx��F���Տ���ܦ�.���dc�a��{�D��l����>��&��;���?�������Mhv]��X������?���>�#�-���9k�peA	~���q�a�)�I��:�ش�k�����-�bԺ�6�ü�uy�ج�Ml���&��<��"RX��}գ��ȟoȪNZ�og3x�uE9R���8̏A�.�}Ƅc.�	�Zu���jR���ˏ�����˒Rr�9�r���
 �U*m2l��;�xhhn�c�����%&e�4
`4~Kp��D�̐A���g9ֳE|I������*s,�����|k5��S�8�ۨ�5 �Xdi3�1���k���'�x\������<Ⱦi�^V�*;���Yƹ�ap�}�m��VӅuŋǸ]R	�:ͱƎ���=!t�3m���������.�p�?��I�E����~N!���1 ��D� ���`�_1Y���ɱs����]��~���7����
��{��r�r�n"�+�W<'�qi	6�	∐kpW�$mn�T���GF&H <�X��|�4��z-S���i�v2�x��XU8b�8�Ӄ�U�z�P>b�Ìw�$n�ȕ3 S�y���>k$���aR"��w������tps�V��S����7�<���x&_^����3_��d�����Z�/^�X����@�.��d��}j�6z� �b��z��k�Xa������vs�^���[����a�C	���Q�����s�V2\cNwu���:�v}S�fL�j�����l�E;�}V�ls�4�����}���f�'W>������Z@���[�ko�j]s���-T{���	鏟o��1�>��$����ΔS�V*��4wn:�R=�\�9Ǔ�K��|׺TL�W���4��#`?��Mu��qt�D]e�gfKk�G{̛v�v��G4fq'��e}�)�h���a+4���\��p�D�NL�	�.�J�MH+��3 �����'~p���O:'�'������,o��ZfPk�`m�����w�rOϚ`z��/�Y�j�<q,&����W8
ZP��HD�'��{��Zd��z�C�:���T"M��0��t]?��EvL�*����r(�, ������X!��d�[C�= ����s5�/�}'��x�SY�oܭ%H��9B�!���E퀘0[t6���u9��a{�Cf�o�����F�}�s-��!���X��RB���s���DL��H�t����q-J�<�*d����$�(��xh�G�e9�X�{�t������٣���ױ��v@���ݠ���
�/[^��*�Y��ZU�c��dܾξ�L�W��Mp�+ߵ�z�l!�7X�P%S<fԤ5�>I���N�Ϣf��x�C���_���@�!]d+�A$=g�H��b}m���%�R��Z0 o]�}�L-�~��UݧBdM�� �#{Hd����˘H4ԛ]3�y���
G�6�~]W��q� �LƩ@n9{����?�����	A�թ'v8���V��V8	=W��S_�op���y�P�*^{��榟1�V&b�wx~��q�D��eZ9���[&�z�̰�/��K�k�ŃW����PS��Cv,�nl�ħX1/f�v��܍B�RG��5��R9Y���Ѽ�ꝛ��O�s�|ᤱ�*��t	3�̣�k�M>����.O�;9N�_���eL��j�[s�-�5�]�S.�[�W��}xo���u���ڦ�w�Z��S��-�c�[d&]�Q"DQ4����5[W��Ş~>1�����H�#�����YWY�+�`�4pŽ���T� P�ɥ�������P�y� ���$ߐ� ���6����p-�l�'��I��]*�J�Vu�,��GߍU�0\֔-�0T�i {wD��
�a�?����o�'�����,ǉ���NLQ<�f��q��B��&�z��F$���]$X�3�f�ִ�?��$Й�j�����1�FٹF���2!`e������$�|�4����5������I���z�T�@�j�Z躅K�l��|6�n �GT�K���.��5��zY�0��pYk)s$����4���+q�)C�$�:#�4=r-������M�]�F��we^�ƿg�ko�FA����v������)���[Sc	���F����D����(����y��n��2�5`�p�b�1�&pe7ۆ�|��:�H�c: v�[�-�?�.L.<y�t�Mu;� ��|HR͋��$�0��_�HT�.�Oa�䰢o@���_w�����39��x���l" ���|��|#��{k#c��r�'&ظH`]�F��u}S�B�9��d �z3�^�Q�b�}4i���YI���@�������'��ތ5�'�5���/��=�O��-�_�%y�����_�NSzش8��v�o&�H�:�	��1�%�&��=��dz3���ۭ�Q�/��>E���s��~�/���U��|@��N��\�ܲ<�~����
�`������_���b,��"@�-��z�8-�~�۳q��&봘q���Rm�g��7of\��ɔ?�Z�Q~���ȶ���2�/�di����E��u����b��8r#~�<e<�����Qc�7p�+1����&�Z�H�����) X<��u���b*�*D}�T����s�9��W->�s�}��~.�[�ys`�ݮڃs�=�lu2[K8>��󩿘[��_��A&W�8s��܁܌��G��+��äĬ�[���&���V�np�|��I��{��tn�~�Q%*۸rV��׊���?LM����HAz�|��(�l.�.�v�a�3�Qކ$�h���C2���{��x�&��xtX��Yj��	b9A+�T^	L���(?ɐ�!p�!�)�4�g�SF��*]B��ZU*^�͙j����{�neV��+�h�(:3>P��N�y������U���[�螽��� �K��%g(�=l�j*���0���G5K_�²'����젉�!�;�rS��P���c�)�;�CFy�aא�p�4�J|.>�s�º��{����/�*�?'�{�4����U�\�\�M��])^�h�{e^��G9c�TH��L�+�v�'�g�� �y�p�� ���bi�K�%�\��@�Z(��W-�?�)�f�Zg�c�Pu]T��ڊ*���9�S��]�^�����Ot����m:2���!�]4�:���,c<���#7��D��g)F�}�4*$)"օ!²�52��G�{6�	���u��ƾx�����7�<���D���.�H��PO�M��fv�ں4��\�܌�� �;;pl�4k�^);dj�i��q�%��Nd��rM?�6�n���4���������{G�y0�o$�G�@?
H�A2���ꑦ��@�e<��M����\�O��њh���t�P'g�f��K빵��Æ���^����s�x�|uq�v�!�����X* ��Rt8�Q;�
�c���Zޔ�Ѯ�q���Mo5�¸��� -�y���N�zPƊ�|6���d����r�Z�#7̚���Ɋ���[�����<�ߎQ�?�X��M�\Hq�����C����߶G(xN�|�����O����ֺy��;�v�&��.Ah?�o��jY��+<�Y/0X��[�2`���w#��.;���&����M���c_�@�'�3!h���7��l*��e\[�ڐ�(�s�N%u��,�L�_PÿF�IKݷQ	}������n,ߧ�5'�d����D���MMrZ^z�N˚��H!��^�ra$�_�]}I�
��(ۼ�m,|�c)���5����[;� �V�D��`��_�%���0�.T4\��vD\^Gd�$��_Ի��t	����<���� Wj|;1ǽ]<(<�Os4�p����@��' P�#��D9�i���C�(�S�WYoo�>���GxZ��/&ѩ)$Y������0	�l���Ag`�r���5H�*��ǹv_E>�̣�d�ᖕ0_U?x/��X��7�������@v� ��ɕ�1�VQ{51�Y�9ʆ�e5q�x~�8Ma@�2�Uf����=�D�v�B!����wB��˱t���F�r�\���r�J�w#(��0v5�I$Thf�����[��R8�"u���#iu6�������w����.<�:�t�곛��i8hM6�;Ϋ~*��7>�2�[����=N88?}�������8�$>|
H�+i�������:1����6�����*ә+����\����P�����-0�8���'�#k���o:�>� O���l�+���8**�޸Oe�*�_>���ƛg���G��'s��>6�8X� �π�]��_>��r��ȦVޛ�̱%�h��A��]/ )���OK/�2�,�{� ���N@�����O%$Sy��gK��Fr=R({p�.�fN�<�y�P#-TԬ�~�c`�n��vPh���̩���D5FQ1׳��M���8*7��X3R��smS7Ю���8��-w�=�}}8١�����=���#8�:������?��ooLx1�d7y��\����O'6ϖUf�/�p9ЪP7q�r]Sm�ϛ��������(�Jⶅ�
�^ŅT��b���`;3DD4�I���fCo,��N �E���\���<|Q�@`�Hǣ/�z���}���
�7\̨N�m�93{����E�J�8>�u�����>��)���R��6�?��=��F�4������t��D}��=�'�]��D��Q��b=�5n�"�.�+BvAm���?��n���c4?OVԿ+�,��kM�0�8���^{�xFSf�HT�7��++%�
q0սil9�-�c��Ȑ�K]9���O�oT#�"1���̵B�>-�����KΈ���(�������c-�6 ^TϷ\E�5۷.���e����.������P����VǛ�x�����ֱ��㏆����$���nbxL�'b�U�7�8W~<��"����D��Oڥ ����m�F�= �*RN�ḩ�0Rg�q*�kIkC��U!ݳХ1xq55��:�R�\1U\R��M����=��݂�JV�=�졮ǟ�����O�ܜnF�ttv%�&���>M8e#2����ϹruGsF=ht��W?a(�*}�i[Ww��P�d�6B-��I�C�>4�I�2fEPڹo�5�Ƌ�ׇ��Y#��ʠ^@�O�;N�v�u�����G>� zM��ln�������lr�i�x�3�HSx��g0R[X�5Q͒��}������j�J�e3��<<�4�)-�#
�-�V���bo�'�i#h;1É]8#P�r� ����;:H| 7����pX��(N/Q5�����v��� H�h4�]���â��ēĀ���b��X���8�_�үfB����q?pd��0�Ͳ)�}"#��6�d�<��Ch^��o��U��&8�3�&��2���Ђ��bC}��{�n_���0��僃�g?b­j�����A����@��$��N>�<�ʀ���]�r%���ԟ��9�-�-ly-����	z��F!�ؔԚz�?T�ɵ`���~���ٵ&�d����6�s�rN^s`\v��?�3�3~�3r)�1@��+��<�`��gE�����S�v��Cf,���f����N��-K�a��E�Za��ϊ��Z�܅�����cj���FMP�ĭ��H��\ԗ����������x-A�]ǯe�j�Չ���@2������v���/�`k��Z&��4�zr��vg��R�O{��k�)-����^{BN�s�n�y0�$�G�q
j�ֻזp�g��m��C�K?�`���R �gU�Ao ��~�
��#1@�4��ԟ?��Пs������]�P����l�i�\�F��?6u�u�J�A��XBz����g����G��F���`���TQ=(X��'��L��
T�Ү�j[�ݼ_N�]b��ܚ���D�O����Nm����y�(����������b�r�M��|Z��t����#\�F�2-���/��C��f�'.;�u�%_w��"���_��z�̷�<�������+C�J�V�Ţ��1UlR��m�lA�|`����`��7�k��QM�'�A�����Q���`0-�_B�d^-��qo$g����/q=|bi��%�4�'O�)
\�k".W_ߌs�\�<n�3����b�@���X����"��	A��>�ӻ�w�����=��(�Pdq�ߵ
��`��K��w��Dk�-�
/V�1������j�2W����P=����T�K���2��ڱ��!26�E$��mJh�^�g�u�ǴS���lN� (��qy����>�nedO�~@�J