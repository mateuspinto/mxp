`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17056)
`protect data_block
7HEXQP+X0RwsWkxDj7j69l+PfIw73Zw3fkr/BcdD7mQKOpEE3ae1hwZqoGxz/3ZfmclQ4uwaVtmY
XIfz8z+EbmYU8q6rK2JG03SbKrJ86mNnny1nyfs677Xck3PCy73SPzt94vH0zw3ytRw1rejAIItL
cQQ2GP9cyAIdgKMe/grynZbG8hQ8qGrkNGNG552z6qNT2ql7LuTLJApJZ8qZL9FdLsnxHqD/OuVn
PrSfQHdwPfBAOrERNmNwf6iMJbWHjBkCru0RxTWSL0sqUa8R+NgPRYbbiBW6qy/xqg5LxQqAzDqk
XUjkcqAG0Ic8cMAfCazNZF4JO+3znP/whxqdBl7HzRmfhPZlc+svVto4raWdazdYVOqHtjTwxQmx
H9UshTAariLYRi9f4/YYbAiMlagf8gDrNwvQXr84OHABcs2yhp1QzrfiJgz9RXaYh0hZRs0Yp6Mc
ggSRsdTl81Td8OE/zP3rjPlP6Ko8oNap0WXZspkAtmvEEtnVwWpatSiRRTilWZIOgazqzvfo0wMw
QTWCUrdSD7gwJgUxJWuEswOSKssjy2twVry0kxw55/Xa1POL3Xizp+yKjKQr4qhb4v4ye6jXdlEM
neEEeyLulZkh9cqLj3vguL4STWk6tc/FRFlf/0KDtjYAc4Q3HRsH+BoABolF59Sdj2PC8VlYrBaH
1cZqVq98Wr06483QB6v+MD3ixglA8GVSX9D2ln3oFXSZxFmsVvpNb80QWJlaxzdr6bgs4Im+RdXc
qrYZFig5f8rYHNVqwLYBoV/eyxFsXCnyD2RNBTC7TPhKBaVH1D0pPXDVZysMSxTxrPF75z+/macw
gewMsnRlffE7Mj2Ha+c7IN/Xh/5/xIBsMaELwh9hUh7wB4T2ea6G/sjOQWWlG918F7DnIfgSZgge
cKTBJNy7dTWvwv3kXNZZ/NjbuldnRuwpZdt/2B6adpF4aVw3PiVq330aD09vw90QE7K3H6/GYWdq
1ZUr0jq/XBhJmSxoaCEXeP6zVdRpKT4UVB4yNawXbtaQvOKUetpP7R/2HAYW/kZl6h35Rry0kNSI
BICnM+dd+5ObdxXWv72dbY+0E2yEewdd7nCJ28VlKp1yS6+wx/+2sV6EP5VYl3+oN5s1pv4RdXpi
p0lIJ8ClvDcAZKTShyWi3L+MYiKg3vopZR3owV2FAgQmIrd2mkt6B9REmROByVhKWO6LVAGV5dMb
B6lZl9HvgOAItEmCoVdYUHeyz2HwlPVNbY92Sd4+WgxFS99dn7NlG7I4hp6XBl6gpN8NYfTMyeCH
5ibJYpPVwtlsqLWKL3Rf7mOf1Vg7FY3bQ3jz3KJRSP8LwUB6o3KZei0Lwtj1PBHkYO5/9H2tY70/
AuNP4y0hVdQcbYdV61cXcG8fxAxNrKu0cSe+XWP8RgA2P9WRvEUMjrazMRRbjHgY+5zotUAUpgen
5gdiRxZ2W5AAsKrdT4SSgRip3tSSeitIyy+uJMFH8Q2Hp81yLKX2fYJLQ3YzmUz+qE2LjNBFEKoi
TD4oI9QYVUDkppLWziV2OpdIv91F7LWjyRGVnMkTZ1rThTDWZO3t3HVA5RRnfq3vDHuyPOejaSl4
B+8XgMLZOcR4bx3452YQNqGAjSdZvqlbk0ORWekzKg779szPf6lll+IPhbUf/RFXGueU/CgMub1P
5TNjiZc/5jHyyXAF6enCTiIWO4X3+w1BlqVYV02oX+y3Vme67tKqNodQynd0BvgEwsd5+CK20vLx
9xeSpIR9cRPB6+ZLDb3x3yqYAOKyNKHQc397UPo4Bi7gOsIkNeWKT6/bQwvXRWXrEsNw3yDIRlRK
EjUUziNLaWRcmDaWycZhmK895NvJ3zr5sCrFIfgqKPsqOPcwCF01pIvgayT5altncmI1cH+CmTW8
BDrVri6JpVNcDDxbIOObVbHjbeXjRGwKHa0ZiC8vd+alLTx2dYMauY3UVteY/rCFrDJb70xODjg2
8Nyq0lzKEitrll4DBBHJ1plwQRIhh4Ug0t7ihDFor3WpcTNoqJBbIjmlIDFGLJOz37k84UHxYFD9
QjGhKIuaaATJ7ztSfWilcUnsDh32RaFrQFeNmKtcMB67cEv28WCTgaqPWzCqNbjJ+y/JTBQnbIxM
z/vgR1di2kH6iWvRnSj2I+G6Qchci+/jDzrSGa7/5Y2o0nDpKf1J5OgTA9s7NtukNzMtHGAHxovo
KGsZebwGzPBb3HRw4HuMU6ajJcQ4Nw1S4VDPF6CkbovC6iuTtCTSvBtL6pMr4MroCtNlO3nZIC6r
LocAg09OOJ5eMchY7M/4mpt4RfD7RQVeYbqZp8QHHxtil/Echo8XBs921F3tFGroBpKLlD15GokS
cS47NKHiGgnO1hP4xru1TWhCDQmcotVffO/r/xiCMgqewW1bPX3M68agUKKcDjv8xCYk/rN9aUTb
xexP1xoE7gdRhslUnkx3IkuNHpjWj4ij/7UaGc2oQcyxFrGy9SVBLBpPN5Fpp//NuNei4OSBujaC
RAz5BlGgXBRfo8J/fYFWg0qQU6GR3e4nAHNDTWuDzD701T/h2EQ+rRTDMUIpwgjulgE/f3WU/37t
Um3xd2K53RLpfmqFopIHUoXCguqKp/VdKJSlQd5wz74cpT9w7sMEiIeQQlKW5Giqf+l7A/62EEWd
VSgcYq2VBRoX3rMxPT57YrRkOkmODkAVcu5SEiLMn0JmQdOXY+0I2hoQ8knEL41qiQYmo3rHawzG
rORqZH+OJ1B4Yvhmio5BExAmUr1jbvcsObHF2Jzq47tSE4MVodpCkO5bq6Qp3qSNxUxsSUrfGEaP
S+bhSKy3Zdwqe4l4PqjNDe/hhz7UW9nsgrYL14M5yb1PT+3VL/WD1QHBmYwmcwFJ8ij6uQcpp7iz
VoNvjQ7luBH7wlHsf5u70Sz+5PCLVironT3ESDU95hCM9qnwAjLzDmehx8pC0eRLFGiFzm07xQkJ
XOuFt0Ka4lMq/v0wRq6YSCdRFHurwKJNn44FpGgPREH96lSvYY0hqys945eJE45sZDGzDpBwqmtF
Y31oAc3+Bu8KYsyL6A0MTeMSGs+eiD3YqqyMRwHvHZ5hbYuEnjDAinlkWV1yKRub8KG3cXcJ9toM
wDP3hrAUcuyyetJIMlrL5zKrTXFzYhI0LDSoKclNgg0atJwG78ro/ls+pNZaQmH91GgWt///zAAk
t0aUPV/Z9GDYfszr+nkmfbWLx7I3bAbPG/REsGQLDxJt3B4A7hLuBw22iP8s3zyjvzF6UYeePdt0
h5La8yc7E6GJBh7HFKpM1ae4PhxsQNzdllVf4z1KAYM+MjAHRwY3uPmJws9782Tb7NsVD7CzQyVU
3CeMIPhPCd/VeG2kglUfTIRDnCJ0nqb5jH1aTagSOvfAaqLRvjlgPRBxd7RZ7XvUUTfjV+BaRzCk
cZzARm3sojuDZBM4n3KJzHIjmhVV2cDQLNENQdXGDoX1su9VOq+4fkUstOqg1fEotxWMBrjV/oQ8
pzox5OzTGNCeGOhyhKlN01XrqKs2/C1A335yTUitUaXZsRif2CYk2RCmbJ1+h9+z5LYLEQcXwaw9
UX6D3LnGEE8KV4JvTihqgUVUTUx2y+l+NKX6bogoOKtNF1k2xdDtQgb/bddOwO+xM3dTv0ifQ/EB
aei30nvsMV0CKpJlmDejBxaItQo+Bop7MOGdOcE/TJqnDxCG/pGG709xSFOvQzKwxIHAfAbFZad0
69nYoIVEziTx5zmpAwRUP1uxmZO6C/ydjCRQ2zLtakSj/XKzxrUIchxGs03PfDMKwTfUtyvw6zPd
JdEAJhDp//6YBN4A8Avc/B1A188hxwKLuBpQqNYymIuCEdr+fT4+sofOF1vkX2GRBd7jcOZH5kx7
vrjomvEau2VGQEJvUJ11QxfNJGJOTHq0+ur2F0zXGUnAFq4Xvp9OlrNYQXNQ83Lnz/JPIEzvqg1d
9i7FiO6c5yQgzyTGUrD6HeoNuRAOxTWRBwStNZsUeWoeO0IsRyepQ74h8DpNTlKyMYhl94j8voLz
UjLjNaX21ixYq4Baz5AttfkS6XkmgbvtzIidtE50wnWrJLxJ3kvNGXL+Ry0CtdCKOBJmRKzZjBYL
5H8mvllpck6jHBAikHH/MisID+8aTDK/Fz6isLwru1ODx+lG6lSwzend+Mlpufr4zpYwT3epyHYg
SJE3azt/ggH4Rufz3Zm/LeCwXEJnmX0pp5TUpt+DoRRwXFokeRF9MB/GfO2Xx2cNKDcd9Zudih8R
HfJw1jtJxjD3ILatjdwEFxy/INRpjPukcnbAofmILZ/k0OkEv3XnNKXPin7LCwd5tf01nUBEkIPX
iLuFOSJcHarmip59HhRYWBBvzKJ7FZdvrPSQhKm+UTz0CdIRlAJM7mu0kibIOEbM0d+jouw8xnyA
E/WOJIkvrM3IJ/9JBrYKNWFI1c8qIcvnCDDwklpsE7CfEot+r3dX5r3XLz9BAo4y8LRgAKn/XMuN
lT3VjEMfbe6x2umdEqiCzui8McucB+Rwu+KqzILGYWnGzmbsiodVn0OdrgL48HxhIJXv9YbBtcaa
dMAIUx0JlJQhbqaW0GbVJByguc4DPNxzMkIZjC/Y2uUnFSOrNZjFbQtrTuK3lBRrYxECF6sLlp+1
xgtIPyPwj6rc6BcAWA8mHgfNaMJNAUvvZEY9LwgXoLZYVyoyUQD3Dv6/jv34MBJJeoabJEmC9Xal
aRq7MRfHH1i6NSXQehEjwQbge6gdICiRroTGCaBlNJjO3BDDt6Bc1uSa0BeruQiudZNudQJ+FzMl
Y9KG8jFdBHOYCuEBQUgJxiQ7OCLPxzwPhkdFGePDQa2k6FcBy4mzxSyT8FH1eNrcIMlpGhaHR+EB
b/dumDIu3W78kFo+gQ+i7HCkygQdJbRXGUcLodbMMpq/v4sHU/lDahWJr3CgLgrtv26FB8rlCCod
4BqGu4IpK07A0F45bSLd59j0C925sn6kV5yMS2H6NIruRJN+XW1YF2jPuHJiBK1AcMZDef2sl5ox
MJ37nUzDE8RnRUgxZurB+jYty4+s3iVjA4KEDTVAZiVIYQ9uwC3GjXXPqel/Ze12KaQVCcvPxcws
0TmTQRZRejlMCLl4boMW3BhJomcz2oMfz4srCMB8bbnw/ShYBoaypA9W8L26YgonwMrXQuH4JEb/
7ecz0aQST+VswfI4t5MpX4nEYM42LjVcABl4BwNKRI0pTOyLOZGkLetZ3ISLDo/GvbfzkeIh33yt
uKa5v7HH50uV5CMWhQ/1CnZISljnhtVnmzFfgmiRd/sfAQ3yxG9Ujjrj1U1sF+r96fNz5Lhxpqlg
rRsOFbshQnV30lNzGhbI5QhWapmpFcZ37hwcchvRsPpYPcGX+fwWQWxJL7/7myRxyJkdLSfOZbt2
mL7fHvgHh1DhmeRahr8A/fNpECtcwY284urAPxS5UW8L0DlV1ixfwIiHgAHbrG6p459boOiX5E1M
ZGq9wPjKWI0fMyZnqGs/RSH/ucnFR2WhWm473Qn3ClsSrpgPiT9DqE5sJL8+Nsj0AdmKiDsWrrR7
OSwtfBeE8UyIZAeEXSg4wTBU+Z38SDJBB4qsp8wowdQkVnsDYFzmGYnvU5Bb2qkscKAnEChk5fz/
MWOB9T2Uj5LOfDyzdmsykbRxjyHecVkriRDEcVl5oE+Qfh2dmIXusAtCCb1OTRe1oKRl+bB4syWV
GMuC4FIdQEMVXeqIk9uKhxFZyVzjZAKUR6rq3uyMmq9kBC2baATh43kMylTB2c7tQunQSt60TDDF
expkdieRLIdu8s3WZ6B022LakfVgmXfu1NKVLT55Eo7SQquCSMhN/aSo0Qq5WLl6fGoLsmzNnJ/d
tXfv6DxGOCwUYIA1aqTu/qIXIht7FHbHDIl2kMs9TeGOeElgYgF9OaWvmBOeFMTfzqCqAztOh+xj
G70Xi4a01h3yTvv1n0qYkwxLmwJkzea/Hl3raWTRvXn1M4iOb8KfRA18N4KH/KdCOPgbDCrZpP3z
y0gdfW3oCw9rEC8SeE6eTlvypNh2vydiFFmqoUDgCr1GbCwGGnq2OJJ93/iNnQS6SjRH6tFiWq4H
oHzyDmyNDsiwA3nk/rFCuYYelZHe6hVXtQaR87Po3O5bJY7EnqtosrTs9+9d/9V0H3hOi0ZYuaJm
69cMyzPiV48ULmA7fquJ298kM9gq23MztvRPm5YcDK/iYYde5kctN4e/6snVLfaFQV7I7hRtEF7w
W8/39WMRSoN4a8U+pUaBdKOv1CJSWZP88/NEWc2AuM1sDU2VWE6GGrAdOAhiaPxNU5c3ZNY6uEg/
rsS//yN4kXWEkTCIIU1XKmse6NEBtt9d6QyhDCL44DU4Sm0FNHrZ1quyKRrlWkJoQq7f/z3scmN4
T3inwC3g1ikhBrLbqfvfNU5EuL8QdiQHaUPuQ6eNctN9EVzxlp5khXRYMqIPTF25uOsk0Yn7U6wS
OrKk5HOBUbuNvbBrNBhvNxkVY+Ai9tfq+8YEybvgt8vgirxoAXQUx3czv/WjWQSYPLrOsMLEKNSf
lSL+CDQtOcGzoG67AHLFPbzqWgOy8lpgFIvq6NeRrZNDd4SgTsVcJVpMIZoxG/wELb872/PCXyga
W6FuWsU/V483kUa+vvSyvoXlZmCTEFehdCm0dSDrdQJ9THA3LgXtpK9r1FC5u3O+ACMYPd7MVWrA
Wg6OFWn0CbK6AB2bITYddrSGo+f9nOdT7N2h3y36a8+0dr2X8GEg67nZR/oc8GCWYmrIZRr1QLyA
ntxX4kOe1rH0gx0TYY2huHn+bN8Kia6tPTEnwh7LOFqjyECi46frdcuW3lPyaO4dOdmActZ8vidc
NLexHjG+VRvazrSVzWyl8E1+nnTIibV45VDBBgNi7cpRg8WwjQr1V7GNoyvW/ESthcxACsu06d5a
uEHvBzeYo+Urni8dfhR582YDpzvCZ9RDHrEeFiB9eL6TpB49mFBBOdCaq/YX7a3VPdxDYy/d1aPS
H8FcnPUFof/OMaAbWQamx4i828dktws15hBcL/LZacNZ0h1PXe96o7nTZ5kWOo4pFA8p29w6GZmA
YINnXPE29vUpqqIgf6Rt/2RshNFMwogBgKYHtn+aym1L94j3VYIeH87Ego0I5u3lOi+TabOiBWUo
lNblypKzqMYNXvAT6c1sdiyepVUeNJHR5LnhGSTk7CnIAILweZTGmyxfDsTgw7TCyWipvSb3VY8E
FbUDCvN157RcsCDx355lxbSCjsoWPkkUPkl+Ypwy8Y6zavYSDKghn23kosvZQ0wWtJXj/6uwee7f
3nPyVdU2CGzKiE931qLtS/5yxzHfuIYM0JfFEr4QPdgJKYwCSGpFyLuA1lV+7WwJYWNONTa7nH4m
GJvJk1Yf3+Bef9ZTNjs0QiuE4mpAWt2FNOMCnvchjErdz+z91DkwmmPLm/h3jYv9Z0GILeJvwhCE
QXwW6dvq3CVXhnkHWQGNMiDWFRhcygyMta0mDOgynFelTwgeAOoXuuSdoCn/bdZBw5lOXKLypaim
v3w0mISnwfCym94uo06S0tFLXe3kZmoqt+OHdGJKMZZHNK171PPulS/Fjzzy6qNLTx+JxFoGRHf4
iqdLmHKd4dp9Z5WzpLKgHOcgTP7EsRDtQ7wo5eSTV7ZxHTIjRn60Q7rnYoneV7oTW/otNLS43Ov2
AuFeTaWgeuqrqJsuuEVrQbNcN+rI8Rts1sOaymMD5NGWKAN+7qt06SeTNF7zioeV192mk/bK8FY6
kwQ0gE9HsHNqLNJHtjOrD5YCU/teXC38W6Cc3wjktyERiLnXB4qR3iloWBjObZTe+atQGjzLFkrZ
iIO1hSchHJUwC/LQtQqVxuDoPkw4lfoisBB+gqK3VT/JxkwUZFKI30nwvJ9tkIFVh/DpYAnMu/OR
u1ohuzUEqH5wE3LWK2Z0fTF84x++F5JugUFe5frNyJPKJuYrD1NZXccNh3fKHcNkK5iB1YJAOi9B
1OZfNscCdxA5EwnUC0zDwRqX/3JOkE3w1Q1c0dcaGq2my8KBfC7c6DAWo4Osr41m/HD6Nf/k/ni7
zlYE8GyUp1myrPjat5fROkQTEm3usruVbUTGVyDXmyKbUUCwDQ035GWspWhR1YM4jGDnJL+tbU2l
d7OqXBFzwiXZnBAbJhG18zqh+g9FeXV/qXikYsNOM0oVnKdndcNHQpMjkOZBmZOXFp/UCe7nzx67
dH0MmCm17HwfSq/tLLBFm4WmPG17+Ok8DplwGassrStieYuG6UsrPkwn52fi6r6GUzkgnHlsHlJN
+J8aF+bszIKiTmr2znrN1xdETKiiQqU8AbItMcCm6lhIUi6Sb4OcwLmVm1x5/RIOIb2yypMjMH4M
+XuqxL0BvfmMUSul5IKpf+ZL2afVXMdgJyJsCMBBKThAD1HXVaLlFhGOc6JdurWxK9Mu9K9086zz
785C7c8Z86AUMMouXZJElpgejB6eCVwGHzPjc+NpWHSBfyj+rEnNsrwYHEHEhcfJLgVX8lE5aQkX
vxXFdwm6GQWrXE6d+rrMiB3pyg+9eWec8yA092Ygyu9Omqfp5IsuL2RELCrkBaZ68RPsW1TGhuAk
Qe3uW6FY8BvgtXMtOaPWr+bJGd9Kgmqxv8WB+Pa90m/C7cYcNPKjWJZTDKwVWSOuvJvzwrqPxePF
0j5gfhr0httqqid3T3gTtP2ZPFx2i3f0fHiVvN1Kkq78IL+uMqZJQNIyIvV3cTJW9CHCKvqu4tYN
CMz/uj6WmbwWikRF2O0vDf1MkpJjZxm/2b/p6TBdkA+1ETym6bbmze87ZmjLXz7qYg8yy+7fz8jb
UGF+3+b15I1Ocxh2oKXCFRoSRccgXqIUtFT8CjzVh7rp3T5q/dN2A2ojX4Mov/kTi3hC/vte/FXu
Z+auGEHtAmXFqEHXlfZC1dy9iZBqws21DTJxf8/ViJ0PhzvdH7OeQQpnGu1bnbIfncuJYuE0b7yU
v/yxOw6keXBQqMY1YrsWX01DRUCate5HcUgQFT9s4Ym2pm2fdMy1lUeRDSBiaNuVeK9N0WGOALVE
YT+eaMkjAMm5QG5b8fq6aF7PadS6JcvCaCf/dg/IkDHwcSE7fQRe9P+KEgK9bZXL8ku1wGf9e/vm
8fPK/LefmOarl7hTSKt46f2Cyc01CqchoCpVx/qYvRWGYW0DmEc8udiMA3IV7aHtM4deE9j6glCm
PMQ4DS41E5BBmhHInn5TCoGFgi4VgSogEVmyWv4wFQ/C2i7qDAw7a0kSTsXyjarIsFdi2dzZoqLm
TgnFoZkq7hvPCZiSJ4ifVrrbMZU8/atF+RcC4ui37gvqoux/yGWk2H8LmhlgqNbKgCl0pEXWiyTF
Ulk+WCFX/kHRK4tRd3mtnGitUtD9W6XhA5YuXJKRmD/i4TzsVrm5pQp3c+1I6lH8Ml6MWpKj+evu
2c60bbMego669EXLchpDUiIuIdy1okBC74cmKCDUKNKineRHrVKOgAIfDAlvUQGK2OaOAsKyJvWG
s8vVie70YiRZ3UwGhwXISjpQgsAbIxT+9pNfXILtoBbpQbsKMC20iVbnzAyAKLGe1QOVBGjJumkm
WfML22XE4Cu3pD+yWP8UmEW8jfsCBz280NOE8TPrDTdIjSO9UFKygesxotoX2T4GWOrOO4laampy
wGv3/hAFlz4gYESVeT2ORD5tflNmPXq1LXnUsMgylyGvlqfvevjCk22wKOFor+CErooNhMJ5QwqV
UL+7Auld0p3+MWl+WonFcOb6fAyOJ+Xf7qoztuuNENNuebXuH7HwJPqeDKmLmMWfHQHmWn4EFNUQ
HFqTv9CjvzLvJqaBpXXEhngn5NyewcHWv/PoRpTe59LGllfnqSyIAWwRYbpa6A1qEdmr68txlXFY
ByOeSG4hYEyk7W6/g2D14gPuzIsIsUZBIWMn9Zxp4nj/A/MlFr7gFoCiI7DjezBj0aEtxmQSA4D/
EJcIFq4JR4oR9UmGWcVFcRdZ9b+NtqMnzKZekKvYXpIvcy31ggmFw4Fmpp9ALnvbrKuIaJ0tDR7e
6/kqe5tVOFDQPr5461RBvmYIAbGShy3kGNiL+xEuJfhLOYHanDu9sp6VdQUhPwdMicMDPqOxNRIu
7PJogj1D+UUGr5eLKiAiEa/dnysdgMF/DvWeF18+zC5roMTnfTsgrYqRgtU+nrKzpgayg3PgQ0DJ
DAVjR2mI85CNOQuEZkwTC3Xvwe2W/Dd0xZGH5Q+ET+mJJQdyApJ4CYX6iqm+W1JE1gIVlg17IUHm
iCjHBCs6izmKfgx0sEfNYB3Y2diz6If1Z2ckD+K3zLA+pU3tC9Zts/s0pHJ6xSoiq4/KmEv9CJsl
E2/INvaGsGA742y69PfQxiQ2dp4G+w3aTyK+ym/PrOBUglfOTtoTyLfMf3oZP+RlhhsECJybSwcg
JzpX7pefMDaRMRG3PrEW90ZhZPVSL81/8YVdBndXaM0QDryWAzkiqZlyzxNlqmltn6d/05F+p7Yl
J19wxgYM/CAgl79ncy9EdKcLzT1Uotni1ZgreMJOuNehNuE8Teazj1BJuiXOXVM9kBlAhE7DuAMB
FgHJYLTU7W76QV4zIbD8j5IkSsDLB9rKu9xyu5oXUgKERLLjOrJvLDS2PjhcMyN5uA5o8KOa9siE
3PdVhWWLG2k86lvyzvScjUyTxVwuvvdqyDQIDOnMPaOoRFnieEzMZF2dDwuGZV9013r8NonUm1eO
gTVEtXiUDRNN2jo37gWNn22/bU6TgxkXYSsDXabFrkOLnZ+lhR6ZlB3yUJcuSTZhd+aGFy3mq7aU
C/CgjqPdxPDJv5Z5W153sWJWqyHyF7IKl5crqm7uZUigQbMWXJbe6EHUDzzFGqMvG7wT+/4bdVuS
GvLarQcNh/7WgJAAFqjhqW2JTaPwyUYH7JkHEWSh7OOs4wWYfhDvFpPhM5+77D1nhe7hMSDeWM+y
xAzEdVsORsQRNk6Ro3YCuqfKCIWkP3g2VsjhkomeDDLGL9nUVKHQzHiKPM+cmsYiXz6CsfS4Kkb6
vDy9RwC3OlXan8UZr03Opo/Uk+ozw4UZDgBv+G71WQD3Sufd37Yrd9PcoReX6eDgKOZxOkMBErjN
RV9tyXvBvmYkO6Pem1sjuOA3HJDO1k3dXJWkziwFrLy6gg3W0nQPc9LXPSth95jb2skm5GnhzMGk
kVh1ve/ngSNsvdnrU3z5kQXafs4AsRq2abnvH7jjhki22Hq3eLIiWAFkCwtA3nEl9u0TrweUzKgO
GXH4mHMf6BvPknD64EMlH3KJLvh3pB+tTV+DgUTJHZzBQ1N7TSU1dZRNBS56vSNY7LQnGG+MqSNK
6lHb+v7ZVHB5DXDyENw2FlISXo3PCtAOATZkNbkXMpIqp8OKemAQrWYc7dAYk5Cs6zOLG/YpqQfL
MixL9kNvGehy90MFOOewL6B7QWLzFR23QCfINQgnccfGx6ZPxapRyrTzk4SrjrFV1W2+owvAJ0V9
R0BrhKqJYcPGPAEQyHUF8lqH6k5UwKMGAGC4vOCNpCIfFPvOLi6y8E31e3IsuTyQ0l8hPFaGLm2V
j1I3cjlY3VG+8R7zRm4+XpRA4ffQUQmMrjjT8sh7Un5IFH3iEzPldb635LR0hBSlR+tX/E4OTIML
+Q74tWFb273/OF5V+uHv9bX98+GCbw/4pWJKzI4tXFBfq1klaytm/xPDR9+m10YSvJX32+JczTGR
bT3r5+WFyMzzHhcO6kqew1midO8P/cXxBIjQHPxYdISFMB6yTWydaiaOKqBu3cnMWHlvHc0XX5rw
T8CkRoTvBCnknblGlKFfff7ukk8GVPpfAfwq9FGOqg+ugYf8i7gJWiI7F0eLD/sx9bwWxUoY7okz
vWIPsYKBpCwv5KIT4Zk6tEp/+PJhqFK2hL798LIfn/IJR27vyOhdTuuX9dafBQxydtFfZ+c3i0f5
LgMN5K+FoRT/+2O6n2PTA6QkZOhRG4Ixb3qX1uRtARdeUmtDaiOCSPUBoq3xr9/m7CSsIqHqRNOe
Ts4ddcbwJ8lgNz9rEkTBb5dw6xGnJVgaVoWTbzAA7tMD9z/opGTMnerVB0WpM3oyZtK2Fj2IC032
Fb1Sf1PtwHGs01Q8qAzS0Rml4sf1mTKHmwBQ38PfLdZS/gQF/2vJEkLF+vkAMkkco+p3BlGexf9E
PNS5iRdtJ0NGsVrbeDGlHw8Y9cXE/wvVQJWb4E+G4TprJQUopmLzLwvmeILlzj1s4LGIYPbfFDv3
HnkVKC1CnIW/FORNa++lWowWqLeTfBGETInGl2ST1VhVKTMeT7SSMS68ikxYZhcvBbhwjCtkegOs
DDnpuGP/oNX/StWpiqjKqBJhupEPVHwn287yUu8hIfG4vfiijd2/WM+8aYqFucR3XEFb9g9Gh+y9
o4vUwPS/8dxZ1NGiJCU6rLJ3DgEDo2dPD0oxmiAxGIYHbmbWVZEWOYW0MwhMLE/W59TyLz2KizgL
Q2yNHG2Mh9jxvBWpX+Stt5Wx1Y8Oh+FIq7LG0Wacwaq1gVhokELulr6CQKoLCnpLV7EQyV2Lt/zM
on09jeqVJ/gC8DIDM5ZTLY9jyndN1qvqVv9elsEef6yHy0DzIJOM3P1C7xdm4FFL2erLfy54mi9o
5+fiGY0dAGz7v9YnDHCUEn+2Lg1OLmx/ExK1N0It5lGWCLRd17rXP1lQUFSFx8YDWMv+fEu1zJf8
H0oa0Nw5QMnI/qIPwIAQVE7/TLS7WcFfeG+N5wk4IjKH+FlFBf3KC0PVWdN94fVHTrgqW2Zjy8gi
Ne3dleuA456GhXmr2dxfu7Lvr+UN77NceLMdqi6WJ2UcDNVkNzEqIsNQ0eLT+xqpfoUy7cYBGcz7
u6K+4myIEuZ1sVB9mWhNC3jaKio5gTl5wG6ctPXwehRxVxEumXMO3uqyoxfAhTpu3gXbUICwFJrA
qjAiobMzpXNmQqRwTKz1Cvu8Y6MTGLrM1TT7w6QqxciNHYgJV5EMBTjtexO3EIxWKTYjpz4QYUn8
nKSr7AezeNgEt25XpEmHtQGFCa2JqHIK34bTOXEL6WNSqQyvgeakQLuFGYUYzUbIu8vvR1vl5+y5
n0KeSGcLtYGJhj+ZBvpJuw9TTDjN+Cs41lp0S9SPoisNAuHgpHn5UXRtj9Rw13lY2XXH36hnWCcc
+L3dU0hEecdJA3ykwLfCAcodZlycOX12QGo8JPi9Us4Qa1MDmcdeJxn0C9s/YnqMoG1cK+Nx2zVr
JYQb9By2Z8UaCxnMLNt01kY4IjgrkeIGkNCPZ50ZyT+zbOmCfu6JCJ8jFLgMIq0oCJqm7uOwE/NS
FK7xZM1UuuVQg0Km6RYWvoKp/BGOudiKG2UKmE4DUAFSOb6GNmGWqHCFY+YfSF0ERb+Q+OomvOEO
q9Vk3z28sRAbg3cxZrUMA2W9CYXpOMi2zQllLZ5faNwS7hSHM91xzPb2P7u5q8QPuMkL72t7OjeF
69fKoxKo0UkKfhaWsgyPckFKuNeDGs7b6ETXhz7ryP51hsekKN+IZaOubs5G3CGnbHsl4qrWJOHQ
L1TDaY2rY/wgG6N7eTl/mOKhGkXpUKnYNzDkjA+YpyyUq0PMYxfa+/syzCgqdR7lwmN34PnMzJsz
AhRvxEm8MNP3hoAZYk4xt/vuX9a4z+hnGkwJ9HfN9xPFRJ2141+ts73MHJvKFQD/0XmeC+qxYhbu
b+ADjyeBo0fTaWrdY/xDr0ke+ZN64j517OxAuosjz5ZMDG9+FoN0xDNJggdL8PxIhqAwyI1zCFp5
gI9PnWruqfsi8JY9gzz7FjBuiIwIqL3Udv95aPBGl/Oyu8X1h+BIHyOlx5yX51waEvflp9CPjFGe
JpMQdZMylgb84n4DyWShT6EYcvpWhkXHvozaS/3x25ePLqB9UyS08pO/b0t4kvrVOVfAhxyIrIFd
4QqjLDl6ib9je9NiFDkA9n4bscBK3wILW4nCPT9ej3E0HAW1udWVu//vUk1N7YLilzYhpe8UrMbc
cXBmDcyUc7NJdnQlXAFFk3qAWyOjZPazFqxKgptilqiwAAQuptwsW20ZHy9mfSJrTUBlFZSjrrDy
Tyu2cT5Ipzlp/0FWQf2fhJrnc/x1FLlGJhYbFZ8VrtUQuipPw/pUa2+tjevvLAF85J7U9YHWuVf6
3Unt4iWDv8Oi0m/qac0eOjdav+zHJD5MCml7WOpIWfQxfl0RrZ8nv2tnuH2cMEs1KB/Z82e/zWgL
A+iCTLPNEhWhzSjEN4lHN/tnrkzTinCeeeksVz3dHDlOJN7y6/F6SgeNUVaEND7xCRJowKAPMy9g
8lMDUpDpk5yWdXMHh3LTzP0z3jJR5C/zXToA0hQToaJLu7R/kU/3Ik5PO4jygs2UjVyYi5Rz/TBQ
iyAPfwXojSbtUdO41veBA4Ux9vozckyp/E4auIBtjz0TZfIall8iL6XIMuNpYYg59GV0NcHg12ld
VHwpqu7e3QW2NRtCh4euerjbBrqc2gh+pf0Kr8zmDXsDvXtcxOVyoP6jswkeKAvGlLif4SEqYydL
c9JLZ/oR5k71LY3p53LuykiJcwkpGj7xM2MsDi55obXHoEPVdZ4jQimYMDYc7zGQAOIdsj2poFti
Zo+33hH/bU/8kAuHJWL1L0RMgCBPrlF8Kj6rVb6HnX91r1+4VV7BqWHs+ydgU6vQRYH84YLCuHB1
gWChwh4zPfpKNuexn42Qypv3AQDDERcY5/Xu+puPJPXIbliwYboEnkY/9rIN8mBbqQx5xbjGzWRc
21Es3O3wfNwj7BmVXN2k6GT+wEKSqi9r7fYx1wRMNkeTtlc5Lv9iQroHXzhIyeQtWkx+WNt2fA4h
TQV5WtwMc8HrbdhOBiPnJQqH13BF+oeRBzJ+T56u7J7JpPZM4v4skVVCIXXMIY7JLFrK/3onWgc3
uaQYTuXbvJpGIkXNUgrAwu7rChMx0WtErrYP2zzCyQFlx4W6tQgi8k5Y81D667HAJHjk3AoUt51Y
7Un+aHgqrEWMaKMZGskYkspzWTOTlrSjM5MzsLuHfBsbWfXgdoL+qHUpeX5T+xRtlNgCY+0Oc1o1
ccZTO5i7EmSuR0nNo8PLIMFjgJkWe90jO9Y7V+r6i98dxdjhzYa+6RLdqM41M643rwDBiegzEnrw
2fYiNsqXU8ihk0qA+0btIuINUdvjkgU9pOxRKnVpXkEGHzP8tupYb27UDrzj6uSkvpel1F4GjpR4
TXRjSf0oCsEuUQ6UGDRk2rYPqp0jSs3wusAOkop492WlnwRFc3cY2mkG/bur9LJ4zrxRyTdTV0lt
1g9GvssDy8ldUFngWyUvAh95V38vGxE10A79gNrKUqYbKvAqJvVifCQt3PgyczdwOzsbLmIGSzgT
i1znPKOV7yZUa5XpGkWHQCH1+9FMx0R1dr/MMzI/J6i0Jiuyot2RPIuyTWPrK3tIQJVHH7FeMJCy
7gAsoE6FkP10n7nFi5HUHE1/Mbfn/Jq11LvTO4PIFFdHYQBkH5YAK6nIW0UnBG3n6Ob+JCNlOl4I
JjlwRUaaJv9nYv9M9x0nKTuPmhquWrXfvP2ayFDRACxpTy2bH1umxd28ne01bSQzqXTnRmRbwsvl
8zYnJrj7NHxOFYWjVf50wqZI2Cl+CD/C6jW+u00PVFOTlS5RVqhcWrd53IY389Rrr6qlDiz3CiTb
3wwC/BXRiYmwxiTfE9mUm/ftrjNDS1d0V8ilnzx7hGMtHZDRJXme7MuS0fgwwEyi9y11h/BNl7Xi
tS9vzIQx3IkbDa0CfH/u0GI26uLgNqb3TO4gYcfbZWTCq71dz2OCFqC/Eol6QtWuFADcDvoyN407
lgXkFuvwT0J/qDzO9qLRtjtkVs6gc5MZxxzsGa5Df99wXstTcuxD9f8YKLUkgBywZOu2TdwcuAso
wpaJrXKCU++8FVbbNCyCyXqPads93RO0Q+tn7a/5iaNjgr9GRI/nd0R3AnHVCkcjqhQBrsnolBA8
91cUypxAeeyte4iVZNGmbzaMNxGLzqnx6p86TrsIXO/dH6lgxPOKR1gkXea1tiH8V2P2Ykll/JAk
bD1yOwIhqlik4OetIiQWzzGVBJn2V2x7Id4PuZSvfvApPZAxMzU7OOcg4i18XrqzOOYg6NVsWGCp
yPAIz/pGuCrIV+UcAtcLaWF+ay3SMWzeHPYvBYyxjG8J+GIH+TvOrkLqLEJu4HYfTIiAjC3WxGBO
+Rgj50OBqc6nLLbuMhAFXtHJoniI5H6vO3JgpE8zRLylXXLMV8Dp8HHeM03LOpzZIqJKcbacfCy5
jR5nOIwzdOs2/5Qc4ME6rQ/hqoZZVNOJghHwXcAUK3Seo04tYB8bgSaksnStUnsOOXLR/0kZ5YpX
o2mA5gnpaR9SXJs647t0VSE30jtAOCmFzMQCLULSVk4q+KfZUQxgHlqx2yLNTO8uoSJDf4Aj3SV4
A0eLN4gRXI+31a2azfMg3PX52aAc9bNUvkYkMjlDoaTMWdY0OjAwvhlcjYrpQj1ykFunMqeD3oW0
oy0itOfpu56IbE73TzY9Trvh2gtiRrq08rbePwZCoGGEqcQfMQngSNLhaYvnUyKxk2Vvc9kwoy8n
5j1JMW20rl9hypjTK3qMm77zcKiGMXitQ45Oe0qMw330K60ry1Snn8/W7yqa50uLvdRiWKGIN0w/
dMQXm0IxIXoJjQyqI1dXplLjhbrgaNgyTTJXSzYomTFicYsfI0x4/dS7y5c3Z1foa5g94o6/WbM7
AK0SLJt0qkZjTBiietV8ub/3Pso22wKIk4E8wkYj9vuM24OmYCV3hagw91vwp0/k1+myN3/xehRM
XAY4Nj31nz6qk3p9amiLBDzGHXKeykJpUYlDqTT5T65zU/drGlcVM8CFGIZ9fDrYl5ubLkXTgLfY
RRG4szOT4Ld2tuHQ2wSqx/Mmav8gLDdxYwEO3gvpP2c2oW76rZTonMjYoKed3iqQX12j02aWaco/
Zbt2WqjediuhDkoazXJ+hlvt62pIteTTgoADYqQdsAZ93wUjICDg+1vIgBMO1NYJck6GAtMJRvpo
D19LrNK679UpVrzLnvQcfyVqWDjUe8rcSvJnN3bpFTNbkvzMX646scQs45S0h3wzhYBw5n0Brf84
MUpKFWeNzlCuh1lr8Y24NYL7Zw2vIpeZZEcSOInxYEtBT6Wu7iJLv9ezqx0vXnDJyR6QjrrJ1lG6
NPHgHAlDOamkajndRXeRh3UyxtHzBYK4BlwDtSk0Y1hxKjYBH4NbLHBWV+4V47oqvN2enKtlVc60
O1ywfl2HbysGgwadTFxoiitVPh8X9F0Pz2yfxbrVlxU5BxqKOueW20P1/1wQ2C/jSPk5NcrmTfOM
RU0fcfjovitxmfybUYMrWEzPjvPFx3+5uHWcGRhlMU0dVucrdDDqwp6XQ8EhGMAguJfp5KO5tuj5
E6iHtlspKTAYGLywam9dBNCInytfxM1aB0yEtAxfB6giUAVM0QznfxDx3Hd4anOM1j5LJb58jOmo
oAsTBgnZr7D2asMo/dlxeOmOitrrok3BsWhCuyi3BnKnnbithtXUFb5uOYMhbfT8eIbkFuAIx6z3
Je8O0m+3rE6djiQTd02Er7/V/I319/5NejBwNX0tWJpptmzsGzdO7wbu5xm9z4wip8x9r0y3iHpB
tylVK2dQa8yz30jK/3pLdll6b6dZMpI0UnaC2MlsgQO7m4VCkPazNYvxQO8LVYL/KrBQy9TheaHB
FbOk0tzEJhQYoibjZLCOMJXVAiJe60wbt16Avmt89gtMAR//p+7XUZoDV2sA5gV1GDvNXiimcG08
XSlqc3JzhUrVzYyEvEWz1YpozU26oyke57BCJmvg0atFinoQM2c8eK88v7/u7ExClJtGQ+hzrIJt
piF1b+rghsvbll+LqFE/AbBrGfMgVVRcanvntKhqf+aKgKUsVQYQfrYPPwj1Pdc+69NCO9GeHhCd
eKrB6oc/WX3g1bVl8xsZ9CDaCq2IHf+fDccQfmyM8+3FqPk1AKsVwjbywtq7pkQOn69fqnQmcSGy
6lMvvFVkooEvWka1kkuvhXwJEcj6DTtGgv+RwfzJscxaqw/skdblP6pijIFJ5fcL7DXasoJaVZgn
FvFIg3cfICAVnclrkc9qBtpVlOqBuvqqs4UQprsIwHG/0RmZnALijD85kv6hfZMMkL0JtfvCzrDG
GVskOrY4fuuFQNrp5ufxBdtN/KrCaBIRSkiGrC89xa3bVLvqBd7zvSeTnHnOHIa85srxzWwzjrtG
A936HKTioQyodEmQCJjsIswv0kxzMu61zEIxTBKAnEu1E9PEVUIicz0r6cBB6mn/VhdVJ8xHuiTp
IGvApTmo9wMLk646OH14W2Zkb+lNbyXo3fRS9Y0wtP2ZZBIZTane2w8SLKlABTVUns3jX+wAj970
+B9tZgLuHoJhRCXIhlPSTWh9tTar8vqrUAuq6XRzHqVaKBzht577nrsUWlxbGhqbWE8Wxdh3DLJs
UmE8KKiBDvh+JRcRx3Y2PcD2y3zte2JjLuUtNr+tB7jn8WjiyvLsfStwbo/U0AovOtLNetOxWOcn
gtYK6ONF/448Uq8fE8XBJhZPQrz7JV5Agm37/Wjho42lCNbJgQt2n5xTfbIDWSfuwqP1S/kv+uRW
nkcx0BQbY5VlMYravhoQ9XZRD59r+0DwekuGnbuynwHvTg5coTd0n2LQ7HOmNAo/zBdJTVU+vUOP
GduTBcaEszGewxXghaA62bdzPLOfJUNQbCocqNX+egPGW3dCn3ItPzzWH5f2kmcAuCLJD7V/oxPF
GibXFJ/rPklMYRCLuQhFuynJAU6oT3Osw5JKKbf16GavxTRYF2u0Ms3LzH5uyGn0l9iT6qg9UOxj
sjcl1r92bRp3kAYKcSzb3Ec8g8gBRHfIOBDp78H6oWja9qvTbyNTZ0atlqLA919x+fTw/1qx5VNq
fdbdm0SkFre+SLdTa+qb2KFRFGK5hBGj+uLFgx/ZwcfBwvxBKLF4wo68vtdhiDnB+rJkdh4B95tu
GwscrJ/NNRKBprCFHLv6Cg1Knv5/Wk690dgjznWOI5Kl0EqCQBMApcUB2hFZU0eWmQlR5mw7EKAX
Lm3iU8MZk153MjbU814F6mE2XZWPRyxlcvN/vGbtfMCMjg38DktB8J36qEaUw1omP5h2tC1M6mTS
IPSuOlgMt5HSyN48qmDPWmTM7hQ6NzxZWqOVyeMj+UmoroCZvkA5N3L0OmI63xQRMFLKWw6Sjg+1
dOHRrx3bYF7zAI/FWrw2KMliBksWf2Gz/U23Pug7Uuc9LwWR0jKFaKV2AQ2v90DYmLmeWlBPiQ7P
lRFDzkrhvRrEoqlv/G4Dwzjj/YafFi+jPSixSu8tfFSijzXF4T7pCFhJ83SI4aGZeSqwX+kGAYgW
c/KZO0tyOhi8XxISZ8Zqo5lq5MoznMVhaeyiEZkhqa/znYZyZKldc23ar16BIdgcO7QFGSQbnjXc
0OA8fql0TaZsHIYa9pKYxEquPKtckgM8oIuPyiEu+6VTRxmEwS+UpvcHdgtR2ZQKT+IJvmm4b331
wKTW6NJIQbxxNigyojpH++wzAOAN6t94JlUprBwW6iqcieGfqFoXQBoYCgwhLvlAUsxa1YwANEcI
kZn1N38N3CWxfsaBIOIiiCIz3HCcB/YLV2QnzNmpnbV3FNEq9vCtr/vKl86mCxSnjfgSss6dPS5Y
seN/sikY8WulI5VewUxkHrGRYUG3ZY4taJaDYhldlLPxrF0XGFiGKKTp4odcwiogEezeagGdbMdD
PnPvP0P6opP4JRbH+3O4+imf+bRz8+VrvTBkYFNHXvJynw8DqWfjDwMRw2jhzyJH4aM1H95L1nQk
Bbx5fWTV8kUgbdPwtQzXejNarRmm+aBD/lmSJSXWtc/+Ikx3YxLWp6yNGjMtW7XG1tkyHiyC2OEZ
pQLAZ/CYOOWTTIL0dkbs+Fch2xbUgEljPVPFzfnCOMxxi3hZ8vdayQMsRDpp2KpPBe1aBpjKAnfS
+CFfBCJH8GLDjcFvciQmloxmz1hxLfPGt90euD2dtNUH3Lf1lxMQmSP+62P2U6VxmJ6DAba64sy9
IBTUrq/9NWc3KsX0fnwZjVDA96mc7L7Hxr0gjfe0ilSLr4JWEWrWmLswAfPvy/W3E70VCAaFYHS3
relmvEJEVJVnUS2XO8GuLRlJz+N2E1Mlj0q29oH6Rque74ix4oD3RBRQHpyC3agX/zLi3nGAwc2t
C0R9eUqy4rCscFteUR+m12GTRMpTZamJ8EleVVcLMAn12LgD4GOSeOoFm76FF9JBme1XgtbJ2fib
n7LuuWMNvu02DHemHtqRQuNHzSawqaaRyS/sf2Jr3YmjbxN45+8OAW2oKML+exShoY+5kwKXlcjD
IwPNvaopNIBENf2vgVoXrt2xkOkaODQJond8ObX7DaaeYlPfCQRWP5STzi1ROWJRk5FDlbWXzgbg
n0+WSL6VmIrwbIwYKbjuT1uN1RLM9WW5kNK/o/aHEAEZaLDSJtFSaE+AsPVRDiMBG4fn1qSy6+F4
dxb9zMxLzsQEn2N2G70FW4nCMZELk4CCFaYfBA4bixGrmP5M6Sh7nPd7dJYMbXo0Az20KiuJWH6Y
uCp3Zh7JfGeiKvcVgeK6B6HEFcQr/yb7F2bCI6B8c3+6FW0dqqNhGshuvbzh6Mh/cvGq5PR87wC7
TFBPxgR5J+B5uqTxLbXBkm4vJvHJbI4eO1o7KUJ5uV+AS+r8CbezXnDtZRsBEw53yncdo5CDZndF
2HYD8FXNignsNU83IoiCynM9qlXHfSQUlTpvTIZebMicf7bjSzXWhCP1jMYL4VfodxPod9NRMk5u
r5qceHTDL9cAcovKTYpvIjNBDTf89tSpki30/c11vFAdJ2qbUuh0GRx6/y05+fivn86ThEm0agt6
IDuZbgcKmRq07tKh2oM8A6pzGuSyYqLkeQaxrdfU0pRTxUxD/a9G736jfATz4YvVWFmRXxTaMCxM
NmyIrAQq0Y+CB9JMcpYs4FbmFeX8ErRIeDkX8Gu93UDstvtxD4UwMF1br4DIKDPUEQ2BGmdg+1W+
tIgJzudYhy1KFDvxbaqr4jpiTkbEnJPTe3Q1r1qjyHvROBvIrMM5jwQdonI+u68URV4dvkLzP9x+
btgHObxPVnF4ORBf85ulp8kxUXJ+yI2p0B/1qLxwcSDwOSjH4xdUnVj1SFEqGdtB6W1fZMJrvpNt
m+XfPMXx+0Mdf/PUuJ5qFMhkHl8rtXc8MmB70qMyw9kREr9GPRJtzXyxABxD7TiMZy08zkfZs5lZ
ZNZLgkhQ3nZlOb9ZgHAiPTdT7rQ+ReeNk5wmbS4jqfzqYU2bQ5lkk2lRl9Ai50Gg0ymD+dXdC6sr
DTyRTqw+YH1nZ6UDDwtHBhFnyO9NuI35I2mLrmJwl6s6lGkUsZ4ifTSOSFB8BzhHf2PSeFUXpURM
FNtcK+x9EqdNYAZxaI56BZdMFevdtIsNIjk3dfjJrsX9EqIOiZ1Wh4BaDAQRWm36DALuG2MjG6XB
E3eEN+62PQxYbTF66AJrjZuQF9jOdA82/UuomGjdUatn052nAZM1mjQ6URoBsCpoZhpTLWhZ6mo4
jHP0TR3P7Q9qqB5IMnTWCD8937StiP0H3w+uX29rYVe/kxbKRgZ+k2ENcihB+x/oDT3yqfGXwtoY
CcawjiXkRLOvYkzzPbMu+lVMZaAfk93SpXX6I6YPQJorQhBGRZZWHfi/NMyYTdtyItVvSwrFeUcY
FHwcK1gUea+tjQ/O9Yf1DL0pLSu2zO9AZiZzMWDCk7TUSPWZqzU+yWlr9DWOVCiJD8UIHkxAsby4
x1Pco8y9NGGK+XUGY3vE9gSNZbebdVEkQoZP2874FBO49BprLQWiI8N7yH3mxR9fabrvHitg4U5U
KxQXoqnrrMO7kIyMQCxnVMaZltAouXgVtUVsljZr6fFYMtDAJ4S44Z9YS8buiP1XoWAJ4XNP4tJ5
eJXVxbcAshgHLT/q01jcNm5fh3F9qLJZAH4lUdqAbT5pfnkx2l1z8XN2H2wy6iJgpj8WDBZJSF5H
7sqXmSaDjDG854NcrAFKJDHfivrPSyo1LSaXxGXhguyPa+LrMgnQSrwaSz0vJyJsHIqGEcW41jze
/mfxVfTJGHzUY1HNTema943jxNsIxFtK+BMJA+z0LrI/C/3KW2C2upf+IG63j+U5XAhlBGL/4tG5
VCAzEJyag4/tLb0b0Me/AEvMzoZ/UGb7wM/Z4soxyGk7HDe3bp3hZDSGgNYdQXcvyYKDmogf0oIE
6igSIO0r0RDBKbYHIHS3lfXfVqvirOxL/HM4nli89EXZHs0EgeLJ3m9vPR/ZdUMIvPM8xXeWlVQx
9jdVOppLU4/KSdoVX1mbIUAjkPcM+uYmh6raE1gb4PBgsWCdQcPdx15iiNpGF+uRlrqGkMBaWdPP
4U/8Mdl3SPrE1IDl+bey7S5A7lX0XmAm+sAacs/JmV5u7TOv/c6DC/H0sAZORc494i6IkIK3M+/i
6WSGHPUQY4J8u6gkXhfa/aY5QqZJhcVP//jmHGFM+uVbeGmh/TVpj0r/bvIKIk54XJ8gTtmCtG+k
xogSDtLjD2VgtbZuIS75n6V9gmyJGUlwZmNvd572DBSO+I1pYVH4GKWZRYS+659ubBnS/le3kOvv
LATs03eBTwsfn9EiMMP1b5ml5F5/sdTFjh6LrAZGQFCcrOSNto/fuv7t736Ns7bBxOdjiWABS0sL
z49WDnOOjGhdsjiEIQ==
`protect end_protected
