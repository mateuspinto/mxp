`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1120)
`protect data_block
0USWSUGxovGsyBJteYpEoQMYe57U7EVv4KgCh0gNmqIMNeyn0NylMhbEz7Q9aPPbVwnh19A+zPnJ
GV6MX29zfY0sRtJMTgHCLe7xS5v+rr91hEwovxoqyL/IS0irnoDaJSE7SgtFSp8WdDmswgukHZC8
YW9IJaInHng/d+a1Bw5svaGsIAhoJvBq0wnZ4QHoTCJPyoB/w/AzzuWhtow/jLEsbNMzZxqKsg8y
dgPZ//HFi3fKTDwYG3pMng9rQcXZYtu4TzTorkcDP3do5Qnlbe2ky82MSfqTJboIAUU4XyGNt9qo
Tly4B0IH3/f4RJ5JlcNRtNmxytUyoeu6QSNxwFWipAvcz1snJAyCTzaXViRy0OkWz7Qiuu1AkJhn
BWvVkt63T+Qm5zNLmhC8NP2mg5RL4Za25284256jteYDA0HvN5pllvBvPPhU1xhoHjAP9kpUpKUO
gFdxYYzIZwJ8HW9BGS6XCS1ob9MmR1Azvt5pehbq9AlB4/r9bzD2Lvpdf6ZXPNV4kjyGDvajID1w
CeadjO8mKDlVp4lHCWRK/+0aTEdBnVIApcB7GCqjz2u+ST5NwSEPc49tCgvcTWJykUUVOB8+cNVD
ry/ldz/3ua3uZUUv7Lav5A6YkTzVwZRvYQ38p3sQQdFecjxx3a+XGhcJU9iQIdp+LA401UbZ8Bv1
wl/khdsHfOlSUZSXB3lSWNcHJP6oYeWImhTZLo3liMlgGTqpKW5Bl59Z4mv08RXzrtIgyhZnO6ee
ArPVDgwmDxgKmdlv+zphyqNF+ZQ5ahwXcT/zuY3SLgnp0mt9lIn5OuqzoDNvB+FznmsWCmAc4YeO
VN0LUwBYwvH1Q+iZbL0UvQkZFJeaRlKUCsGMa7AV7RY++KY40Qitu6+p+AmQbOk0JSNGB6w8r0l7
gAbmzm7n4omNU1pN/iq/vtgwL82cp3QajhkaQ5KmWYDFKW1XcmJWJdx/N1wIPVfaI4TTDor/dn5r
HiQ0po+yN37pfqRI0purYzIYV7lTroxTaj3EwrKi+GEbi91R+6DaHFPy7+LVRT88xdWfoGOS8i34
dDaD7eNvifjL/hCpItzDyEfwpulIFiIe60hgjNvT98LQjOBr/XUjrPC++SksaItqzRKFhDKLCCbl
38Z2DyO/l2Vyn0JYs3ATx6ib9aZzjdcUNZFHIRx7yHa4Fsd1z3uQs0o8vjgvwSfFxq2XMfcNioOV
zRD0ffr3a7ESsLK3H5NUK6Oofq/CFZrOe3qFMEpc8fcxI9/CzTfAzM9G0DkpGWLgODMN+0/6OVbf
15p5k2PG79o155LLcKQu2ViDA54cEcArChtj8au1Prg7XLLEryhkQxNfVKJEOSyRpw4n1G/+afIv
uToOi0fwUElHfVh+jITB6Bw16llG3LR3yEcrl+smlAmu5aL57IaxgwVZNJamgpIRSe5h7WRqAEsQ
ukCDrtA5H/ndS3C+Kes4hGYeNFGFaLElntmL2/2Lq+SznNu2vQ==
`protect end_protected
