XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��p�Ӄ�p���͹t�?�-��Uuz�3f3�����������v[Á#7�<_�w&�᝗<�P޼�&a+B��	)�Hr�"�U�ƶ?9��w�w@���&�l}�`�\��X4a�8U"䟥4��q���,�Ѷs!)��s�i�(/Q�����з�[�1�W,eL�8��Vy�e�(ogD�s˾z�_��|���Fp�o��S���]��2������s���=�7��_DZ�?tk�C��V(K���m\�r�%Ë��<���;��
�dv�0�s�h;���fK!D�r�Zh��2s��[��L�=�s6��L
c����*P���ME�$��T�Z��V���LJ�/~�b�7��A!���
́�<SL). ��Ym};�����d��^rQ1�"��g���!!K������ʨS�.��M�Q��9�	�a�+�� �cx���Mp��2s��]��+����f�o����tH,Gp���P�^B��r΄
t��4zCe����/QJD����'�e��`��,����U/��T��#yҭ�t�"��n���_t�����\6Q�M ���n񍈿�7G��>�a��6��t���_7���|�Z��H��A@�,(`9F����[�h�(��7���5c:܃F���JŻc�|�>������y,O�������r83��݈�k:p�g}���[ȿ�tm��Gn�K�h/�{8�h$3{d�tMc�2�<`c?|"]�feN��%D��WD�XlxVHYEB     400     190'�	�	�2��A��	'�$�x1M�;�"�&[�Ti]M�@�+gAW]��H�7�Ȋu��ٙ}MՃ�$�h����;iv�:nU_�s�N,ݟ??cj>\��G?�m*ڍ�ǻ�X����D��R�C��)2.��%��Q����ZֆhGT�� 3��mҤ�>�̘�]N1')c���٥�����bAQ���j��*H�=��B�j g���l:�<�dy��� ���uh�_w�X'>�ݘ�_�pw��?уw���k-I�2q�l]l;s�g�\~�Ԙ�P ��(��k{6�)O|W�u��WNmf֟��{���L�,���o$a��w�Ede����GO:�t\�5{��^f�_���p�&�} ��紶+�7�,c�&,������K�)5;(�XlxVHYEB     400     1a0���&���Z�� �SF�<�C]+�$xf�R�;��yp���|= �ޓ�(j-�?��?�xY�ޚjv��yJ:�B�p`����=�!��� A����[x��2ZOcV[l�y�6jA�������O3�<%���{y�z�`z���>��<��N�{ VS%�'���5N�'+��7a�ۣ�va6�y��N����4U���<F��>��]�h�H�|�%s��?�M�h"�Ä�~%ӗ�PvX�q�6��9��A8��(�U�e��^����WP��������5h���A-������é$VU���*��%�;3��%�W��a3n08i��<0k���z�I+2Jѣ���[���Q1�[B���dƼ���cy���������>��&��� �KDpK��g�!FXlxVHYEB     400     130Q:��1��)��I�T����o8s:ognRs �h_��hpvU3�Ou�li��K�V�K�<�=�b�5d�r�n��7�=<,l�F���R�*�E���w���_�Fh5vTɋ�xQ�1��f���	�L;g&�]Ț�Sl6��F���lCʫ7*�vN����RO|�?�$�d����� V����u��ޮ�g��_��ceK�tw� ��2@V7�K�ޓBW3����Ev�[��p~UA{�bޕ,�K9�A����ʬ�u�u�)MGx�ZX��Z��۬��#%��,����@ժݳ5�XlxVHYEB     400     160�M��K�����H4=�y���!����Db9�?���R&�@D���&��!�J2�[!Z�K8�y�DkVQ�	��N���g��1����_�o;�܆_�;�)"PD�[��-���ܖ���οz F�!@�&=�>��u:w�W�g#Ʉ�:���	�����KH�+���'�a��#X�G�N5J�4=���N�G�Ę(���6E�i���8d�｀�C$Id�v�u��Q笒%�`b~����N�%(�u���Wn�G�e>�.Y{Z^����t�+*\v��ȅ����~��:��ם��-j
�9�a
�-�v��Z���N
/]&�"��2/�&4Iԃ���@�Z�`ߛXlxVHYEB      3a      40Ι_[�yI���.m3����3"Fs��?�3�Tœ>j������m�&��$=�)i+�V)����