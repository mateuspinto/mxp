XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��~�J|`4\x�E��.����P%6-��,9�C�$�6^��9Z��M�@�9T�>���"QV�C����y��^��?Ma�&d��l��t}]�VZQ"=�~@(!��0����r�0Z�٪疒��,yй6eu�7�U�0��|U8��ڢ`��Sӄ粸�-�֢{�0�	F����[��Q�l��s�*9{�3��|D�B�6b��
����6s�Y��t�b
c�&���Җ&uW�U���F6���]����<LWna�̕��w���!2�;Q⌻I(
�_�5���C��Q�g [��A�f�N�<�H=�aN�i}Z��4�Z���?.`��yɅ�mo4"]H���P��b��TG�j����ڿ��_�k�ç�����붦���r�*b|"�����L���MV�ʆ*�G��q*3���z�!�ŻlH��cx�?h1E��J��/T�wJ�j薬��L�J2D�g���I���M��r'�������3���kF6������n�W|�,-��H&�%�����m]���rI��;���L��h��eqd�Q�b]�V�NP�-5���ȶ,������F��dd�����)�dN7�S��v����\���u��<�4(�П��l̀Y�����,EF�H~/�
�Үͽ*���������2��(�5l%�膿��;���P[��%!е��I&	��
�v��y��Rǿ�7����d�6T��a�4U'~�r���{�͆-|���C�}\G�Z�^�C�XlxVHYEB     400     1b0w����X�8����[����m�[6ǚp@U���G��v]j�=U��[�����Cv%���ܯ�+K�!k^񋊓;mg��)b����aRe@
���׮"�F��]����X���cB$���+��AJ���ht*���J--	:m�]���=�с���0T0b��Ԧ����xk9�����1����u>O�R�#wP5�cm�1~P𬎏Rn�7�V�L�&��)h	��9��D�r{M��yf��}'�����>�I0v��OTb:�7��Y�F��W��=��`G*~��ބӭ1�#䤨9�F��9SE�Y�1�/_W/�N�<�U�z:�QO�kR�D�.JX����o�iXI�<�EW|�9j�s̜ ����nŏ��}�x=wpF<F���B�Gi��w�2vG��{_��@O����:r�dXlxVHYEB     400     150!� 5l�~�ne��~�� �h���� �E���;�?Js�\���Z��9PhLi����V.��c��O���a�b��I)�|�ї���1�5*�W�� 3*����M¾�p�_;5��������<P;HQ���kK���3�\���a���h,�����Q����X�AO,� �?�1�zWf��,}9��H�����Hs�_#�S�ђ�P� x��\s@���7w�3dk\KT��&�>�񬘴��f��hk��XA䩄eϕ	=�F�H�M	�b�o�,��*4�g#m�R�:!��7��C�4���2�@eE�� �PI����6l�bַ�7XlxVHYEB     400      f0Y��S���6�����)npE)��������cw��t��:,� ��d��9 ��ԗ����"TDFG��jfGN�4�h�Y�����2�t�s��o�C{.S��i�[���G� �zo3ؓ*s�C!nD����F�q��<"�^��{�$���V�Q�(�K�'�Wˮu��c�af�\�Q���X^��q����q���,��gd��o˷VS/v������\�Ul	e��"X�M5XlxVHYEB     400     130z�
D�繪Ä䧞��	�4#J�;-��4*���!`%����;&f�,��v��En�WmI?-=#�!�8����R��;�=��y�j������*�
���	!�]^�%W<�A���9��cX��l�4�d�@q?z���u��yLLeݬ����ᗿ&��<�vXY���v��j���xi�yN��yʪ1 ��������kǤ�b@��c
�����4�G����}ZƱ��3��|z�������(�����<v��v��i$
��%�Ğ���m�.LW�ZE��Շ(��)��~D�}�����XlxVHYEB     10a      a09�J�z���IYs(.�q��{Q�O͏q��)�X&�i�⠏I_��q�᩽���]�2%����� �o�9��� }u��X���<��D�$"��'ᘰB����V'�Ժ���F_�n����;�c37�)�Ch<q�Z�*gS@)~�ͳB�N��