`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
FWY1zd1PujFMKhcJ2V6ejmZtIdW04G7+JwctMJWS5h7iQuA2hAvCCSI5JHDfzbLmHzkBRmECWLDW
lEUjJNeNCwaWTMD2czkpZuxi6kjfDqWcR/WnTw2yZcOMnQPxI202urX7CjYLiesxGZoKPZCsj+4B
63v7T3gIpq9WBVhiHDSD5J4DSH9s7erjmp2M9PRs5j4AbXIRFYua7j1ZePQEo3KOwM2WLrsQiHji
b8T1ky5o97GDEVlG+exe6sNE+MK3DkaICFZSPkcBenXynwvGb3AlOh34DIwDar0Xpfk2KkLZDLz0
0Ag6z8edSDEAp6esJY+fa5AHPbvGUwKU8mmDdw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="7sTVxDeBRcqfpD+P0szwSBNsZZJVdC982uGL2jWwjaw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 51072)
`protect data_block
8aAMj5v/tGKcp0ykUftWYF83JKzaCxZ31kp/EeUbM1cR35bD+NGq7LuqNlUhoM8LhNo7AaAy1hUF
hsaqgnh1UOrV5/kbCrPlyabiMWSKkfkkaNnl4DgX382IczNgFcZOLzc8eP7oMmC83mJxiIn6vOxC
OGjxAqrcfX1lD7Ohak5KYdkZbtg2vNKhgi+oesQrr5d8uyIbWvKxSVpaTDZ+WGQASBh1KNhnP+Si
ks+DlAPcAAwlyfn+dklbTrwbbqXpyZoWWg+js9rpD9Rj4Pd6z+dUM8fe8u0VbDtnMDWYENQFdGdI
ywAOrIYQsy55hIxQjNgG8s25i/ISB2aRrYNwHzUnM7eAZ8vvWgfh+fTFXj2rXDCGyt7P8vmDLJ7Q
XhCS9AqPjGVHEHtZJTQG7puue1Bt+HnUq36uZSoELVMaqdFZa/D/WYjrejsxiomObRpc8LPA5/TX
U1khhezcwnjFNbKHzHEfU7bH0x56rv3w63o9D5+IOdW3V5o2NB31W+5qeJAuxfDPpggWCBkiVeTc
TVk2wbUx+5/WTTtPkk7dm/hEjzaXxD88UPt5XdnWRvCrRQZJaFL0pFuFiFCHSy8zVYVsLyNjpYyd
nPZsJKHJr13DVnPz7n26EwJxy48dAVU2ybxhMCQnpX7PF65qybJ4/VBCobQk7vbCl5K4I+hYC38G
e73AFwDrFSHXQCtAdy03WqYj347CmLNJ0BbRn6wUeJkWyxlr1pr+S4SHBinsAcM/pjMQrJFe2g+b
Y/VFIpijnlTnmO2RqTmDPJlfZ/E58PJeQct1QgpQg2AfVfj03waOMkYXeFfgjwMwiv95X6CO8Jo2
nEkfpH+lQt9nDCa1k5WHLRKijW5mKxzXLgB1KA2BpTUdIzR+0KKcpt1my0RgY7sBnqfGJ4KchZ7a
i/mLlvsQeBRXShAjo+431945i3BUbiJ6JflUIxRjkcPTfhYD4828vdjWzqJioA5jPjNWue8+/dBU
OrPCViD3LkaB1p4lTzs2qcu3RheMBOp2Ok8nZB0zuvff3B7RaZKpYhp5k/bAZ+0zmP3Vilq8GxNX
6wcFX3HkDB1517hp3ZoxGDY0eJ6fLAoVaFEtcQU6jC5hqZRkwjitYDt7oP9H5i4asFuyRP2y/EW4
K/qKRPRTWrqSmBpGUZkbIYzEHhcjkpSGqMqsF4hbQcPCtOD3FtyT28ua1QubVvIM0BYnuAPuWpCz
74Z4kuzGXEvE7Xdc9sT0r16bdUBm5V9FsruPbUn6D3RzVqhVk4oUYaZ9OdvWJwqRYfQbU4WIpGky
6uyadNPRBElxzlTp0TLjGPpATRfgHuT4eG0hromGDuND0xmFKAu3UXdCQfxB67HjDLTWOjCtUewM
0c1p8lI7g3FE4rLWF01eyzxwSbTUB+8AWv5VXYfYaAllIps8nn633letqtj0VdpNx4703+9iglL3
1CmSilyFL7951260ty+pePSUR2vJ1t4eb3nFBwAqT1pty7l81aFRbbY83M9402Hzl06tJmrgy8z+
yiLQYbecRwZ2Dy/H5GIpedy7DrOZtLVbcHTTMgKCGMaFJpv0eb9MJ1RhNy3myuHARAV7uePJeIt7
Gc0Tj5oHgVn9qnm5cCkbkpC9WkQ8v8xrN6NCsM5aPLr7kXyQ0NIhYK+S4Ib4veag/bpEuHyRaZ6k
RuDtPx1y/06vpE7pWCUwmuvTqTw++SwHfCvY+dfcVOcejPWLDfQyQIhc8dVdzyGbrhF4SEWanqw6
hzvSZ8uyAuePTFcqTQCO4ADERQBtRUtzLEN4PH5FjRV4UxMMvDEZXATIMhz8w9ixtguCeawF9Wtr
nSuazyF8aJ/q86T7Mf1gRLQ1K23KNYKWg+FjGE/F0RRNuXhYbn1IrF4Rt31xfJRO/XP61XmSXP0b
mrdElgW8fUgqQGko6RQl8n3rhwdGlJNuMRVkIlXIC3/axmDkBXgCr6xD7Yb7oLZD3IY0F8XTvcxd
COGhawV2d6DCZDhvgLpjlt1v1YXKcfAR6WIk9wf+bPAw2aDkD/hi+uiahs3sxzgY6h132+TuaSPQ
2SzF9IRhfrj60WNvaM7rkwmR1igKC0q5kx4yrsAbYUsNq5LN8v/QKZ7Lx3ruJYsB/RsqIkc4h7+r
3QQQfC0j7tHMwTefcZFlN7gh2uN5E5wlQOI3f5QaHm+zQeWKANoEWl+keS7Azc7mbRRJWX/hz5og
peByGkkN4UN161VOqVdLlYo3VBCqWfXhgzRFmLv0FFAtriGfrry8P07N1bJkdiE33LDZiht1pk05
mOd4MTudAikPxFtRy5bXPEA8fWGyUnUYYgN1DtTqUpwLiMxC19E0Oe3d6f1uaVYmtMAHgzsKBAM7
0zno6q7ZENlUvl4B9focsBG6iOI/BMEdLYA0IzRKgr5TldXzY5A/gNvXGXndB5t4iHFIdxFjGXXP
aa4N33YLRdJj82jTLnhzvf0skksI+QabXihTQ0I1aew4XtJKV8k4je1PJgYzsFhcx+iY2vHttAe/
/KZGSAyK3Xr2cmgQi8kdb3DFr338rfPa3dQU6lFZe1HovOo9enGHKjQGIZ8QDxSrbh8mVIktY6M1
f7y7CCZz0rCllqaPGUfSzHEZF3ZZeA/5OEgMTNq5mXWjSKud2VYWzQ/kqPpCQ0118FCYVEzTpCML
DVLl7hwlZKkdkNoED9q6I4dLP5kZWuh3CE+DX9oThPvzRs1EzZ95WdZSTnPit9HC16w24NsSvLSL
dYrb7lD+GlzBgax6mVXDZd3p1kcDGPUnqISuRpexeL/eJvmj5cVd1TyqUJqmV9chp74yMxJIKe4+
b2+hsn1y8MDoKrc9ePlt6kJHs2KFuxBf/MYrxawyIb/UPrs2q7wOTDGnQJNxdlHjTaAnC0kWXRc5
bWPTbVInnGBV+pieHDJyLq20e7EFI+W6rPOqV4GutRkWfQFJ0gu9dZhyvhBKqueUJNNLi8zQ+bHp
vZXqGjniVOSkG+palEMtqNJGIdMxgKhlgVAxyBpuWBJu0qfzsBIQ8GyQ/t2QS0jQ+V9U9CZCujS5
Y/zj5UUVq245d2UhpvCaLa4tV/b+85qWbjKr9etJ8QhSNiK2psJW0u32ZaxJxfImnbsCoeeOe1N7
L0h1b/6ECtll4uyS4h0jFX+BiMRzRBKcjWNF+zCtEKBEUcVVU16jKcaEwnu3eL4yq1U4wtlSyxn1
a3JTnnIYvzhc0hh8sD71Osi/3O+tB9Wlul1uQwm6w1Hbhibm20qj3ibI8/lcpZmnU1Ib3+Cs8Qsm
A5NIPLN4lue6iSMDtuXJ0GyV28Sj+6DNNPWVTs7vz2mmXPfgiPwW20LzGtqKdhNBq1p5TO8AKZu8
f1EKX5FFhtONReJ8cpUTgt57qozJxILq7UJ2xbav1+GyLU+zpKsAR95y7FWWdR6+EnqZRYaccK9N
NnkyXvpfLcV/0/e7wtlDTc7+YPDh3INOJdStI+zfMk33PW+y6zhhXijh7HbXnvS3WaVvJdhQyAKF
UMoF2/ppxU69piBBfLHHdiR7WuJSnLrtA4I1cWNW8sC2KjdPJHd4XBB0/OdUS5GZQgXUK1Xx4cGL
o/xLtVZjBJ0U2ajo/EW8EBPsOWS8Ysuf6uNhamk4oD3Gq1Jr9jtfDF1/6sDPYUGHEoUngSL8grI1
YwwiXJHD230Zf/G3iZxrPEoZ2yz5XB+oMPDiNpAZ64ff/dxMMv5COCpyB4NSPTYXBCZUN2oIxhLc
ornXg9XHtvZULDdsayAFRsJ2zO7XDeU9cIn0VRiTY5hXzXYg3mF2s1jBDbzZb+kL5GJ5qDae3HMr
EKjJ9t1MqyvGtApo1mYOGBLQCEiJJUKJmQxP8da0s6mNQ0eXAQFbnAHyQiIpvwFFdySTV9p9e/x4
vGeRWC41LdfowNGwJuqSULGbyQ664IgYlYUpXlLftHYaV3BYO0N/mHvK+SDHQWJfbLf6V4QYNg7R
g+Rq4B48QG7QDhXuldX+I0PKkwDMmQSyIoyvoQ8V5Tk/Nzn7aG5cENckk57rQbm7SnZj47yBIsA5
AJlSlKESoWZLZdZCyVnnpnbMQE5TZvBuypr3wgr+6rNskfk7qFXeEegnRFfO3ZYTl8GUVg/JfPJU
FkP+z0dEY5i0/nntdpddnxznDbKlMn5STbV+8BngG1ksPmmddiWmapHRY3hwGNL6fmcJKssiDjUv
9FN5tFz39TdeGix+dqZilaRyCpA2M0hjMHNCY4JI2qy7du3zcIofhL21f58vzp++CeYiWnMb3zI2
hCjHxR9er1rdWicSoNN+rPogq53G6oY8bgpdI52glFiYo6/jw0EFNUnJcJJPcC1ztQmqqJ5sDRW8
GBxCukp17UsSWReW+l3FFXDBwH1+hDtkze5a9sR9KTI3CDTXMY7fIEsgYDSL4dmicDnY72dOZQvM
CAiscdo/548UUEo6G63/I0LTQQv5nxkhRAdR3ab6O5fIris1c/Jp7907WvNytt3FmBrF/UmwjExt
vFdW74EiL5CgiLWRWgsl4MGgg7obULUIKxYIsUh9ZF3lCtwZQy3A2/Hsff3mtlq2yOfN20X3HGEY
5zEzzl6ZRRzny2YBdDEwQP5XU0niF0P6K/N2dV95+k1ha987DYqIM3hAroXgWB00weeG5yQGQKcj
Pnb3MEObbQXMOnXTGoH7fivfqAu/NzPlgdnQJkanPYPHr7fpluGI0H819VCasbq9Mwec7UTBHKjr
1Xvs+XfBCEcPlGP07w0K/YZPa1T5uUKnyIL7CpD/1GTEP0z50rsYcvr5hRrdgKKA3B65DKAgp5ZT
HkAtSdyqU1IZ/jd6zZTwDLZnKymlFBZYeGveebk5F10RKijz6FwDDZRolDuZdyKABUUHd6enKN0d
gTHGmYMuU/x4nhdCrKpIR6Bbhn7Jq/lxzot+Jx1Ndmr/v5GxUM7NzPt5kg1kM++MI4OWo3nUjcuB
m3VuXU5xDXheKopw/CT5GLOLdDLP4XNnvYFwfx7icebQOxRdJgshBrNG07a665w73ekjJqJ50W1y
Xsj/ATzxwuhWDA4AjIySdDMewPRVutzZLmbjpnnyqgf8Osfe7oqOAcvNeip/yVcsJrmvjty4kPcL
MaNS7pul7EmWHmrlHWnLtUxU1IA41qZBc0sZb096kH7jb4GQ/UoPsjS8FA5F46q+Bf5zaW3FR3Hl
qnBurP0AgPf6SM1ZSkukze53pwbzcfURZAr17rd1PPAkLEabXyDd4KOsabl52jrKC7a+S+T0qBYc
Q61xn1QBehyaWWmX98A2UlqcfgfesVu3rImus0SemqJyjJ0o9KZo1WqkdYcfC33GCKwVYBoKTfMN
yPj9T+566TkTTYpUAmA+QQFwj48nFbZjWxv8knV+uV8+KQOXQ8AdmLGdG9aJe8+bcH5a8z4S2eK9
shpfx46S54E/vik/xvX3TsJ45TwLhxDbEFMR8kd1eBvebHN4ien3P9fJ45+onsPclYMH16XRYKg8
f0eDLPKiYCNe0jO+Rb8PC1tZqNELX20eqgBIG0tNutnTuwzh6Xv9Re82NWBUIudh4qkJjc5C7fyj
IRggPeruqnwOK+/NHqPK9SCYnKBAV8szXY9GOjIDuhRyw7U8Cj7OyofL9bIDgfSqbjbxn1ticAle
qZFN475vdCbYvdE4Q834P6J4DufJ9b3mPPliDthBdeNvzTQ85UkJ/eI2nQnEZpcGwImmyfe4xd1/
aWhzl2/O2RWJPJ13cGogt5wUZ5Z8X7rKRmFcZerOVg3dGmWcUeZJTprUz/jBnVLA0CqXZhzrMaDo
EO9OTA3RIyN4KITBF9UKtLkbW9fPaMtL4VdzlpLlKLS1Ga6FGGuSNjyjif/G3W81TSXjmH2dA/z5
FqRysEL2kZWQLgamWEhlEVyvxD9hXZF0HKl7Lq8z1CuORk7Edpoim9hmU7KPL1Yw+Kinu6WmgkC8
WUOUKATcZbCba+Elyc4o40UokMB1UPDHr000j1WGKTFhklEDrYwIRnQLoVrl4ufBHz1NkW5QbWJy
hnqnwF0JG95cPNCYA1or/bQAglnkgDQxRlBEuC9WLxxrb2qHuvUpD5jMnv/0LVVG0eD/kyjnhYo2
HBN6WMSLnD8UhJFUDLQi5nGQOJbqexTH9LMCMc2P4jqgk6kpLp70MGNOs02VQmxxj9G8PCfKzITx
rAQY3HPUxHKVVwAV5wvxT5SpZN+SEXLW6OPTvXV0popKHSqvgakq0d0awcit05fh/8JQjvGnqYe8
2hLit8DIPB0K+p4x1vfNkUPsMn5NHdD5xn35LVbTKSuCisWhB9QzQ4XU7EdPZv9IYWSnUvn5uTDs
nb26hQhrr9JIo/KuvkOYwSBUpi9GB04vWP/REZaiX1yTZkTeZ2ZRutnQkehZrDT03KEdrC+oPT6m
PEKVPo7SLuS+93+C8C0KxJDnefmue2+feh9cNxbKhqnJB9Q2m5ZRq7dXmS3yrPXDfsslbCGoD4JX
1JQwHZK1J8MLqOHLzsjqQdSec+0EQuTdqWJrMsI1C7j9BeYxNuMSCONHkccDjZoGsutcHarNIiMM
OzvJbcDjXJ0r15TZB6BKEOKE11UiTt3t87PSeY5BGfKuhzr7X/zwCg4ZFZP3DPc3uN8jIlGAXPNR
1tm1bkNxOotzC9C5yz3A+AQSkXLasbbBwGS4/Hw8R6HEV/RLWkXQvHVa05WTzy5zjTlj0yy6E8Or
4QiO5Tv1JzRCnmcp/94l6bJ6/PGmVJhQtYtL8XPZbTmwXkKE59O7NmpQnJGRfh621PCnfNiRF2tS
c7kMjZRSyFPbwwPOEkXQkxcgvom1Sfo3mcMyxdybjuwrq6jY2Kyow9xSW7xcqEbmdEo4K/86B69k
b0bMiH72XaWw1BzFKquVCDK6FWuM+xmwbPaWIQz1RKWnHgr6b13iaDrZ+e91Im9ePdz76hQ15nTk
DVyRffywRL4BKMHK59aEzQik5fqqMHdXf1XuizOC/PfyAeCKppZD1XDd56ePuO1hjuALOTXoCpNz
p+RBxsGZPoWD5vgt/b3PHzlJTw44oZYYa377UgJoFti5wxT0hOmCQJ82z91S3RYdNY/DWvsTR0Bk
j5La9h+x4yhpfJpHF4RS0Br0nGwrxbx3TQOCe58AEk0m50qHx0dRGGU0P5lUNndiap/Rm5ewUoaR
Ull/LVDlmoWVJnUnAJo9dY2HiX5f4YLMra9+048EeSMXsaRtSkfe0xUTHX1xpINSH6f8piLT7m3y
hPs4/dVUxx6UgW8RbSMuS7ERMAcNyv3dnBNZXoPj6B3zaPPsZJ5hF1v7o5qQyNU2HCYTL5ZL/yOs
zBFvy6kgXYLPSOdcYu87K2ONBFfpU+SQqbZW7B+0SllOhuJiXkTbam5BncVY1L/q4xY1WIOK1KDe
zvt0J89LRVUvmOMhOZ4K+VleMhKZn9W9GROHrpllWuMkDGAbyl6Yz6VNCWSWGmAQtbFpd3oVUqAJ
ZFSusL1LS0Cqabu64E2DgEfyzgW8OG+g06aTotrwabgJhtdLQp8NGxYs3kP/V9bJ4QCFJIafz9ls
RrMb/6D5Xtj4ipNN8mSwtLDJosNRYmMJFuwQeerUxpRX8FZZcNWblFXd9Qc0n0dmi1RQhDscJ1Nr
8xHOo22R5YONvM2uytB/rfWxEdBes5Zd3I7Ek1cY7Q8d8RihER7E4xrQ3jLS+c3UHMuUWJnNRweI
kwjS6vLg9C8GlGMuG9xXu1IV2Kotk70Ca0SICw8ZFzzduV/cmWgQw+u2mNC8FkXt5WEuuMbszIB4
MnnihZDYZ1XCqBtdY+UaO39NmCwW5nL5dxxdIEAPP0KMhkqf6ShS6HiGGyJ306OOTRnDu6rBdl4z
Hv5gO0WiUkrA8WmIbyZKn0V2UNmuePQWLWOb27bUFovOZiYW2akez+ErK3AAihwsOmuh4DAK6Sc7
PeSDiytJzK48bVdmEKRKANURsNuPlzRVOSUa1/hFY+3MFkO53IZ6lfZEIezCl0HwHBEeZI+9L2oX
5nJjnY8IY3YkO7f1D2OcpAPLxgvCpNDqTbWOguTGWeGbi67uD3ZuPAI1G8EnSeROEdHYIYByy9U7
FcmEFlHLbqsNs9/48sy6woLKBtdotouQy75OzIbDyfvy+TmX/6digP9HmS8AsQp8CFGOZ+wCksJ+
XZjPMsIP1uVV11ShXOm5T1jttq1TztzRLer+iLnbsii3/gh6IXBRlT8XWa79G3oKQNew3CFZiyVM
oEuspJH0PrxIKmF4fs1l7mrR1TFz+rxxMEOTSYQukAkyx/Dbfw0tn36N+0QhHIdRr8rMoUmdqp76
ndwhQqpmUOXenDQAKjTzlm5ll1FZvWtXg6XZDjh13GJFZs9EKKJqt1ykNRxLoe2w/D0n6M6Y7vgP
o5+cd3Ml3DGuJqvfx9eWnJc+eFhzb+mM1M38SXMFA8qx74OwPpooIcHN9//yqKfr4iZzs9pmQnO1
zt2eY1MLhU8JseT6HcpY08Qj6tj9CXhzutiK8bDQyivEiwvZp0meJTXvS2zAV9uY3zKBA694keQk
REOizF3WMdMGOgISq6Wle3FRsWpCxic0+dbNyjTEK/ld0RNAY3/KnrJqfaoEPlPc1ly+5AZ+oXig
6nyAkcYyeM/b7L+YVRYfjxNP9AqtTKJzDvh+iID/VxSJEz92f8Y5P4IugsAtzzSOVoKljCnlFSRd
pqjVbETEh823TR0DU8uozChKmSIlo/lIaWu+ZOh3sGAmX5bvmyNqRdMXFlkWiDMu+MugCONgLk8r
b7VoPVsYrx4OZitBj74t89/3+j4p8zvANH5PwLff4BjxWnw8cXRpWX1uwgnzReZj7XTvZ4CMA0oH
Vmb2ILjTgw4n/4GXSqEoW/lQjZNCNiYJEEsuyFMxJYd3c1p3UZ2pOUpfOhjN2skZUNFxQ/Nu3h1R
Pc8iRUGsnPbfkU1BFkkKiw5isgjOLFesx7nvbfZGjDjqt+Yy+H8cXAzXS9zePNy/LXbAHaTCoWVp
EyUEcAXnd0rpLnljyOYkdJOrTcqXspwHsaJw/mX6We/RtRgCO/1ms2a18OqNv4c/73lMcTAHi7DR
wcW0tfasWXWVFWWfA60HsnmzVz5AnIbeiO0qfwXoK2JvrHb/S9aiMcibXBV58+TTw1uawG46sctv
layXov/QGdtUdmnusA8mG9fbetK2nXJnFs5BrLRH+PZzyBBTa6p1FaJ3IhjfUuZO9YdZj/reOF3k
AORD7MHXDnSsXNZZt60yu+qZ2RS0E1jsFfPCqCmMWxN9rOxPJ93aZS1tJZW/IyDHf6YRagZ7ugm6
avxzUru3jm9afhCZHZ6azdFOw7PgYgOlVsFugTYRZ4yoPJva4tAj3zPejauyfcWrEimX9bMplLsM
R4AZ+vDJdPYte3ZJk3j2Ogk0v9u6WjYtp9MZ51WTV2cR1guDz2B3F5CAt8TnT4ul2dGTWvW9S+Ed
g4lNpcPIKxaxqDIbvcxjv5DP2zHC7o/uNAtNAQHJk0z//1r5EB1drXDRatBwzYRlhwDlFVDB/Cka
nB41Oy4buLTPE6MV+cNoE8hY0iuISvPfrRZVw5G+N/3hY6fqO8JSb2EQw2tgGOtMBy0i0Q/gYmbS
z/oxEw1ga17FIOZnnzWJ0JymdVGpP16YMxguoWtudtz4tiyAm0A32il4kEU2q/XcE199OYAn/nUn
iSDZVbiPnyZOhFAwYwiRNh3Y2jBeXS4eZ2+UZi2O1ky4lWQO8wU4am/4unLDVLlbXhNW0y/B8OFO
Fu6IPO7CBvfwLcqrzDqMZCl94gSrSgp48eZYrHsURROXi9gF0Mj+BF8ruWI3ZZh2nJeD7gunRBiL
2PLtAMbopT6qIbEdEJb5kYk6evDV1pIC+vzdnGqmTTitymVJPG4zXXKY/S5LVgk/r4LpzpciwIw/
PprR6ghQlPxwy+CrxeVWIRU16jJbkWKZcxxUn8DpYW0Wkz7AFHs51pdNs20sHj7+vBxU9sS6Zosn
5pbpdZabACgkncnyl/DTKQncLYAM+fL2KlPVuOWbSq2TgvoUODBx3vQnHTRSjxSVG0EFexO0i2vm
2eqLxycbbzSQDRak5OOGIkX32y8iPL/l7cfvfzjfuNeFQx1PnPTWi6t4Ra81/guNTSEVSc8avVg7
MMiybPWJfV46Df4ahUts2jBoexO3CLC16PkljxgHu/jFGeMoIUhWXsO0rpyxgMx5VleJIIEGY4fW
nQ3KDPpktaRO2CERU1T8VnKdmnZpL9aY0ipsE/GCjXndd6B+tQnTgWGxdbmFKenD7w6Q4EAsa79L
Y9AfP/lc+NIxQ2ZKX9eqXdgvJn5ogXlvkaYPbVfhRIT5acehe3nJa8rkiGOQxmtbMP7ivNi5Bl0R
7+M1wEQVUscGiajyTJ7Me9zEDybAr8bAYBSu62+F1+taaNRTAXgHVDNtKE5pb0B/GFlYy0Wgz87g
1XRzMixx2vPBSAL2DyBmHcNP9Te7AXqHSKmEJ6pSPlWh+jIRvPRKj29V9FmsOHXYSiQsv4ZdZM24
dvuJBpZIYkIV/EmuCd4x6OK3XV1973hEQoz8cv+MfCgCQVSvGiqnJ3iC9AnDxpgofQr8Mlb/CrZF
3/VRVb9r8Vt5bPks7/XbllGCRTzYSg851PIk102Bn478a8blzt8QTeY8Bz4TQmesXozIeWvp2f2M
r7NqEMnW6cgh+20UDRVsQpf4Lt9qwwjjRK0HzRRAKAkyQMd4nlyEcJUZW1o4vcqWjgJLBkre5h/O
6i/U6rQ7A5zIoL2rGb5gmzYhfA1Lc8j2zMXH+5NHSy/WJLSHiosKgQBefC7h9I6/OQ0/sDRDTjOz
KYozjo0yC6Ps5kKFoEGTgbotAVLDdMmwo1gJHZi5buBCcxHZgYIXiUWYrFU7NnyCIs84wldOdyTL
rFkCOh/nFLUEOfg9HIFhfsTGDgTTg84iMkoIGep1ZqEqJdhbnQdskZ0OwiWOLrvX5+rr/0DKqTXH
+D9+yEvR1WwwQWlizJWsKXP7lQGGNeW5QT+wlvaye9a9uU5tL8qNN6LpHWP45SPhT84k0z3gkUjE
1WoJjLh23o3UgGbC6B9/mO57DXtXelDAIfnnzl+mTOnDZSFxGAkxnpiBfxwNw2EGXsCVD6PfEk/o
WUu3duqQJHUn8aykeyY+oJk1gXPuxQ9+tyW2/Ih4RTgFfc3yNUaaSC+4Ab/Mk8oxhv2Tso56cBGz
4+n6YOg4bTbj1kwjspjcxftq14XRxqs5wJEpQjfbPMJiJrNUthpY3N2RX4pN6CUjDpIU8unl+jgc
NMjen0mD8tckOT0x+V28DneAe/ZcHPcJir9zi9KSv2AewoY400RZKypZNxchWAEOKkQgsTBkwBbH
N3CSK4k5aOrA5vZ+3VN+hqbAmP410yhPz82q/Oq9OGnBZZz0pIihW3R1bxe9VnRqWYrVPGykWnTf
naFYrMKsuDHummcfcZaYqm9IU5JuiA4GAKH641vqYnUNu/+r7+J8d7YJOmkDCYLJ3qRycOvBVgdy
Aip5cf+wmaFQRXKgV/ikfVb8QhZz+ZaIGrfk4hHuTG3VdWM7t33XyrxKfJkdbXkHpKITuWNiZjxk
VRY7CXU1J5AjSgNG3RfE9EOdXcpEnzq4jY9hVivmtElIx2ZC1nquIHdgpfgT7edDuEYZM9uefuwE
3oNt+U1pP/DqSN/dsvhzNlJMIC1jLPucAl4/TTVeq+ykw6gB5WASM9/HmLMBgFE/+gEF2iBIT67J
uejzdLflNdOOF5tzqrRoyl8QhUkDETxcMjDbMk3psuuL51Cy/lB8S8AQPzs9hjd4c/NP8Ul1xyce
nZaFnRx4++zFJEj99n/O0mdYD8shGAgZGW4NrsjvDrpCnsoGHNHSDmi//zqo9/V5woH6Eys0pXFl
KehgG0vJ/9Xn8JaANF6IWq6jBw5BMEH5r+Tjegggh6jix7cYuKFkxrDIR5qbQC88RBSP8dMwq7/D
hIHUyGFoS+o5W1zFaPwTB74h/b8jMP/1dWkd+fuecblG8TOFmU1VQ8lOo9cU+Wac2rS27gH8HyZZ
OVW4I72PXtojp82gj970bCixWYiKfcRWgyk5k3ZBKRKJ86D3RHOxIJDVntFKKq6L/9hZDaNzsDk5
Ie9tv14pYvSt5lrLhRPuG7iCWju9bLTC/6HcFI+hSYFY2uDYS8eHNfzckucNExIvqkirEpdQHZLd
DTgUPwuZ3/1TM9sFtqz1JyFk6IvPGXI4tDtS57U2gUNJ6ST02UCA1HjHbcrxmsKrg9XPPbHxIzZp
dalUkA/jXx/mCuRrNTKDMZ6hvOCPlJpOnrwe1zX6cCn0QAiz/b2/WDc8hnGXROT3BYD5Bidexr7+
0J7Gj9ptNoSWXPZkI/ARVRsIEwntoJ+oEnX+FqOeXgQwRNd8dVpoND5tJjAukllEgPIYAaMV8puc
dvuVxH6nip5dWHuLE9/9WdHw5w/91S95mSR2XRaNMDJNrQJcMj1q2en5HnGExaUtFVgNupHx9EYT
LOivoGBhZI5nXpPVyy2rUdHBqYYcdHEi0n0fVDxqQ2/Ana3eJauFHwtvQgKXfwaPuXYpBCIl7pAN
pF7kgmkPA6pqjlw2TjZq0gd8WLSSu0vD8WVBMAF9gXXIXfLI6RyLnhIqSS7SDlA26EXjGk60DaBx
sqWa6e7C2aweAvo94yOLj2P70CdXaYE5RYFZta6oC0vF1zZttrjK/YnU1gODUSLSzFqncDKZvczu
RN+5CPaZADr8smgdjI/F40j9zhlV9U0U/Qn8NC7VpZjZVCGmujiJmY77iUbE9fUMMUp3m9NYZ/eM
WGIP0ClRrHpaRtGSWvS6ZGDlevU1HwMHsTMy2zzVOJe41E46yItz5Zgq0+QPka8JINnyMZqeACiU
erW7aHHMYVuCL9VWTjrtpa3pjOXKW3vKeaNxfQNE8EovL8fILWVkEEiiLEXIEqDPORZoDTh/4XNn
8ZGNeVOX8d8CTdB2LaROW0bKFpY99XBJmPCGaDBU5nil4wMIO+/jmCAgvSu2tHYKSrdhrPU1M86X
2YF5Y/Zj2fuy3ewzTxg/kZLBlIkgnIVckH3MC8PsdYfmhOQuQCunNEZidtZ0WL8h98DMoPKdNA0C
k1CAXRFjeR+BDdii4UYL9K3sDxW8fq0sYDL5MXB/RdVbzbx3zobe97N0Q91GcDh7OcagpSKb5P+x
Nu4tBrcHVebSotCm0zeT2zAnMZ+SmyGlHGCmumyIjbU4sTsMPng6ZCxR9nCgmhpHGy3xdLIw7yvS
ASRhYfNj18HbZLHE3RYSNVRX173Rq2T10az2Z2rVEUhGPkELXF+EPAcl2aKd37B48DHd4UlB7qV6
OKyAO+26xrTGTyJdgcMpLmicVib6jpY1pepJonxBqJtZSaC5ZDTWzf77g7+RyHqhp5nUuu4oF1Lz
JQr80L6dTgpdXj0dGaXyrBHwJx3IpZNE8n78W9CQtprklAZsEM6XWs3NZjiE8qLIkTEv6sDKarDC
yy/HrK9HfnEzNGKZREZStQCBjuGwfipwJAXxyY5D3SCRfBwytaIMlMv1KqmOKPkgcJAWOtcRzXUa
riDdP1tnMixzDvzYDnnD3tnLZLDSx6x2V9297Dw0dBocZpCgJVA33b5tuHSI5IsXeAonEqjO+lq0
Wrw63k+fSiTEVZFeSgvjohcwQCpGxhmUzb2VmQBWFXvg0YUnfk8E+Xh8uYjhjErb3k5+aQZakqwh
wPtFbfXjQ6qbpw9yQL+7wrW9oW2PbWq/JjmB0ZIFMvSlbZka1qOBGL5h8z6+kfFM4Tec2oBPnNGI
PAqAj12POkJ0hZQ6q7JSipJMcRJtSuIlGEV28LqmPqrkVmSqUJmLA0cM9Nkixgmfqu7JbYPVRqst
I0U/C7tAauMf6YDxCv5tLjeTKy6CzWFaqdlQOFJ5kAKWvh87BqF2pyfcqbAINcOJaPVLFBhJVYsr
Wxc4PAjTqc0cUbZeoDKjcviJPp9gBz63XeVjrpZIC9Be8S9xNONUOdPJfmFP/HuvA/mVze2Besqg
4kVkLVRMZszLXi42T9tubTni4jt7mZw+WOz2YSlIPn8RfHzn/Xm8IhiDK3kFwpIBogk+zsS0LpFR
Kb4BmFc9DhdhupOGYv21zPUJB/0ILr1bkfZcuUObf6nf20BsLBQxDkwfjmSsBq2269A8CQII3fIY
Mvtdv88UINUI6Y7cHRE5JZqkosFNOIA5ft4rpnpsYrkBRsrqoYjpwZprh5iZWLkIi/edGok5Mddt
gk0cjHB5IK24eJ5rjiw+FkrxrdXMBuE4YT5WcdlrpJ68jYt8qfSUxPOxYbFI/Yu6khhXn8WDD6cp
s7+bm8AztzUHWGWnLUcc+0QgzBAkZIQ8n/cMOOCqERy4AGWQviDTi2LAS8D4jSYpmepBQegGKXsI
yWU639panGHLbUahnAtM/CKNIhMNhB+efO17AzbEwbSbkdhVk6/7FhAklu9EEf6lqq0O+KDgSPDC
49k9vnQsdTjWt5Y3GqSgNbVsh7V3vKVvQxMX38CvdNyXD3srwu+ilRmOoSdAuIr1ijeIVnNmgx1c
ROYQiEMKur3ThyrhyXqkag40Ars4OybyXoz479sNKUgEzHiRh7g2AzyIjOt3rRm9boT+7V9ad4jk
QzaV4hZUVAkkDP7NmYqc+sE2+F9JrCw3pZ6ulCSsfWHwsSWy8mDxIblwM6IniepPHASU7deZqzoq
BJY8upOkv9J6B6TWRsRaLNd4szm4dwRgX42xbPclVX7XjafJgmwQH7d9hJ65jO0fjNMsrWQdlUBQ
eqAltDWcD6zWCZfKp6yoUdSwb/Yg+UXehu+w26u2K+AXz7wiBHfLiuZ1L6q8b+8lDP8iJVqmiPeI
SdDAnz1XBsp4CCJpbWfGSBC8WJI+8vhK9vV/QlIMRuzqjUQaNrLreJaJ6dt5nR3JBknYzIRzq0AA
UH//NkjmI5VnNxj7a5CYfnbJoZlJ26f0AiwZiEdg8ZV4/FZz8iLdu/M1oMM+FcwDz1diE8gJ1BCF
Vr2yaVrXVw7NIkJNF5z2pDHlCx70Y5L0yP8SYXa/2gkqrzyC0SpwEv5S7LXyFoTGXN7C0OjvJ5Ym
s4qnD3ks5Nf/LrrcDEZSiQSY3/CgjEe98AF86W2flQm4mYQYGL+49bSft6mP4UUBaOZ6uJYxrqHl
Fe6NoujFtlmIYPbfzbvs9Sc8JKx5PqwiHO4J6a1nuVVrVwN5MW/dE/oStoLRbtTbsqZV1naQss9M
bGrFoZVgd0TCKa3wZL6ID4YQMduxQJ2Gn0PRm5DmveCwGKdAXcfPN0Y2fGlSaweObcn3CtK63Cv6
+x8hdQcb1MlonaGJ8qzCUzfeNcKPBevrpqJb6DS4Ian0+rqkkLMEY5Zw2SXHLL1ZBweQ7+xFjYF+
/st8SDNIXw8Jnt/vQD9Pn8fhke1E0Jl0cu5Ip6RAteTYcMGGtvNPvHxiNuAa+dwqOthWp7MSif1i
uHsUmmPwkaSS6B5qS0zFOORytZ4As8wYAtl6w0XQ1IsjB94YCOPBEwbH1Hbkj6HC9vYsxr81vHh/
h3w1GECXuV6mdYrU4WoXl0YLl/rBXOzNGB0cCQ3P86XF3ZH1uWxjQK1EQvPTU7MGkrDGCoQq1xmj
x/Nnvd3/jmGGWFvKst5mzVxeVWxgX2MBDql7ZgWxUHo7XrI9slcrBRxk44U5Nhj0OhVgYs4CCPYf
K3zYy8ufzzVafeCa4QXu0hpLujAccwD1cdcBNCM2ldR+/D1fHBDxCfiIkoqbPZpVz/HRZGbrKUgK
CpIugfvLi7t1pu1Ves11AY5HyE/O7u18+DMkDM+jKLAtDPWotjsAvAcDeehL0m0tDnMQJcKx2B2t
2VnEVRoW6adE3N4+lnvtDKwN29Qp6qf889/XSGcnNx1T5ZTiM2kKSFMyCvuKDiRUhAI887SDWp0/
Q9DJDhMMRZCebfRFpi1xzRs6sRztCGp/tN9WaqvGRCt+GWwmZ33KC7o4fml8mOoUpPOmz7K0ksOr
Pq14uH+B+YbrP6Lfv33BRJm1Mhz9u1Dq87xYc/eI8nbkHImOdqAuRd0vh6Nb3yzIFzDw1Ju50FN6
I1janSz/ddMUSl9Jl0TqmOSYgLa9pzUH8NaGKxcJoT3T9d2akiS+tN5yx4Bi1eMSX7H41p0+Uh+M
ttX072cQL6+15Qj07pAwkY05+H13wyFx0lYNDOu0heUGSCoVSisjiKIX/WbiHig7OF9hZlko4qGo
/yVp2YfoQrMLEgLAJIuorlgAJmz3oiZHaB7yPtSep7avmKQvZ1MV1FchHJkp2HBS25gQYaNdX3MS
bybxIh1YVHGENiijNprK2AgwNZlusRhJzaFTZZl58uj24Nx0TWbebC3dle6nvGHGtPp7ruZwsJgH
PeICM7Y0ZrX1mqdlgNSk+3IYIB2u3fZ+7JOGhAu1e69Ab67VB7zW5fwndxxlonN8eQRKflgiH/hX
l6Fs0vIEFYuaGD8YttIqA92Q9YXPcG7xWRqDKnd5z/9T4rLJsBzr/l9lwHrPiC4lOnHhSFzkvuhh
geYPzdz+7pAxbhfobFJL0gMnyruYMqEtlmo0lRcLLKK3BF86XC/vafjW+FKgzzMZ2Hi3a90w2tbP
CDV6sx/ry3CLm6Md2AU6CxWGAcnt0h20tQVLrB1QYWxwyIFkqGagoAASmMSWSqsetDz+kTtEdbaN
XUKZdMfupg9StcbDM/14DsQT00dyFbvMm/8Nj8kIq9PzOJU31XdBSkh+q6gitecdx6NNqAVfJfP0
/Xd+5W92aOH3f5BP7nBlZOelZ4DjZrc60NU1PWP6TYUAey+OZqVgtY3fl7djIAdOlpO8OhFT8Yg8
TA8n2/jIVgonzUcU2gaajyPFvZYw7yKuKSRlB9JJ4CRiC2Rl5CWFVdKwpkim/ba4yt7qVksGL8/0
ZkwpquBJOLJWH0PyLf1b+U1WkIKekKMCqlBSH8t5p5DkzPw6j6slrioU2v4adR555lThmi6cNCIk
EIHP08Q/BOlYFxyhLiTfaH7DNjCbpgm35zOCQzLEts2Ad/LmYMyxIy+vWOwYrGFc0ZON2ORKkL3j
TnoZFZ8gamyRKZds+VyL7tv7EkjVnWYVY5f+R+ldzQF7hKrXoXLM7G+B8bdOg8cwpVCzoWAB/Jaf
KV6Z/VFlagxi3E3j8BnmDwBCyISwbg4soUFDzrDxtE6HHuKi5pHuQ0elI/PX2lvLPTa6PO7IxXIN
V7RrxspIvYbDQp2RNniiK8tOVUuwnP4/0nHZt/TuOrm7DHsXoGqu/zAs/sRP25y2ZP/IKLfJdDcI
xLuizZmoHMKLeywnxtn2eEip1ynYAO9NaIn5DBw7wkUOdxeQB7hLQDFcuDWr1Uc4PfJOsSyS0WhR
cvC+1/37hDqaAoLQdG3wp1nckzHUiw5/PWeYew2XtZ2rl/Z+Cls2gjbaUhTlTxFhG/hchN4EtrPZ
Ei3aNdVYedFoGgjORmh01+1UAQL+2JroSdRkNaM61jXlkkyCJ2P1FmRi6uS9RpWbl6El93pJ/nSj
8+I+lZiqNtWQwnfHj2sQepKKzRl3tgEw7ZCZ9qRFemGjEf9/Q1HHLt4CRp07ARakfeG8G8UrIp6/
Bx6Gh3eJqIO+2Svg641UOlEAQOvVLv+F3h7xiSe6MkKRd6X8dkT+mxMPnob4yVbFwYMwTXTJ86ka
/VzbbcWyoAUEHc832JZMlKEJI9L4erQDHy/ZfTcOS04JwqM/r8FkQejWuLtcHv+M4ewx2EJDlVmO
aJx/4acIjZBBE6Yxy6vg5WvII4PFON/tmvib54R6LbrdjIQLsw1xYPgIVEnJOjBP/Rh7xEfFHtNw
IF86iXOkq6oyZ8wWzubnGjrEY+ez+Uq6/jl7C0yQOOEyhddL/WbwCccc5p3h+JA2LOqctl9MXmS6
bWnpl1uK4o8lmwMlV514Hlu1u8d0SFy6AClWvpA9rhjhojfDzu7v2YdWuQbtF9NFBfDvxLsZXd1Q
rcyky6pSyd6lgKMzzwfBObCv7yn+icQq65doNI9KL6kraloKGsYe/20WD+HQFRoR4qSsu/LorIUS
3R4qY+sTfPE+uCTnwzf71t/Dmo5fErChG5eQaZw+BJPy8km6XfTIcKNSAQTM/VGu3KrQL+Llk7v4
wsj/wdjjrkCWlR7xNJUoE4p327jOTkhJF5r9XoOKySnvUKWOC03SE+jQ5JgAREz6VYBUqx15L2b6
bchzcvOGaOf5CyXEt/gFk/vzOu5+3CbPagTZ1kNw4/spmsE7sjCQnHnxNmDEvFQWsaHOAW5O3B+U
3YDQRaaFhFNZUKDhqkx7woCdMNygbhYrGEM4DWk3a0tS5CSG/bey5L4SWspKMJa9ViJaAoRSxe6h
8ZfrSjtH4OlBt27Zf60mJh15+4R/sCCA2+1d7KXWE0gMP/bVLwt5oor5d0ic6JWM9/CgwbrOciVx
1PE1pdvlRfZVeO9KSaUfPyxFJRg5KwZ4es4ii3w7UOxiMoY0VcqKin0515q/4i9ajUXQYKdalHGw
ZCOXOCh60SPjudBqzrNz49w/sdaS8bf3x9umDRCWSkrIZk4UyVomgLoShNdGPi0Q9HHU1Y80sf0n
DdgPw8lwH+aqcBoyL9XMmL82vShJ4U7gYD5U4DqJt3Aa0AYFea7rgfrDSdlP/SMsIvTSBywXCfhx
dZlcxzlhYKHzkpnB8/pbdRJN+iA19TnNlv0WWc9ErJL6kiTqtLs+IOJeQ8xWtYES7Bqi75+Gjjly
uzwZMzPv4yUlx/BBGUhsD+ZdMuxDCO9JOybMFWU/VwrD3blVpiM0kbyZ7WmZOz+CWDZTRezR6ux4
WcdZ4vwWVDdbzK3Duh1bIwwjMZw+5vb7M5CZxFr2rKAzW4D8fkDMKRjZ7zT0+/1x0KXY99QB9+OV
KwGAbFIs11uujc5gA9Ksckzif6kfFGm4k3pStGEA9Ys4X4j9N77olNVDhp6yX2lQ1uTZ1dyYIFB0
U9jZTYLFJbErjrTl3WJ5t5Wq+EtKN2IfNBaKAFL5LYlSCzB+9GqBWLzJLuty5CUW+CjW6tfjC5W4
945sXYik7fdfHjlqIAOGKdcSL+nqU5f+IkVFzTJk2Gjp27NVoEfV64t4f/e/Ns5I4nKVX91pdYQd
eR4pLa1CHcG6IAF9YL48qXj8ZwmrePcOtBSZKCVQvfXX8szSrlU3/BtDCavutGhdP+8YbgEfjigy
duDacSvW27aYmqkfs/h6uadLy97cP3ISC/dQoChe4sJmI4DefrNX743rBsAvMw02CeHl9x3bSIFO
OKvnJ5sHuvVDMe2IDqePNPZfv1yIKansCcSZULIU7/Z3XnK8wVJvm3EXvs8/Z2S3f7rZRP31lmM3
xJVDPCTFzB9OePqAmMMnp1bZF47j+R0mJXROeqfs8s0UrYP8HLpe/0FtJYkDywSOBGltIJRPhj/C
J5M8drywFU3XNqMn0YvKFvtO5mQLh7L6kvhATZtxm+jWA6khguqatbWJR3/cE9GZleVYdyuy5684
KNF9EQ1HNtdWzLUh9pa2Tb6KHzFH/V4NpOn8EpWty5/ewc0Ax6oFFhS3zKo8gcZhQV+xyLDABjjW
YsjYZWY5pdN5C4xLydxiiqPZ40VNVE73su5JyX/YrBV2Nexc/YcMrwVFZyZQpqJR7lWgDdmkKhvc
mB0cZ1qToHbLpZDPrwHz++EFP49+htiLE0hV0iGEgBCxZSPYpLknHeSbTw5XveOktHmUPULK+so0
o/wgWu/WMaHsTQUmghqFt1/MTwVXoCoI1E8p25xz3c9Z8XVNY6ucRVOrRoSUTMfvhEvyumDmkdPc
c/zFU6gx++p3Sb89wKh2jJBgIc2uxnD34HZjzSYgpKakGR1xPK6+O6seVgCxqQryrEcqUQMR/Qpq
s9qcvR0CnZHIcG9l8OzinvILQRtlZdEFVVy8ji12rNpyZHKTk/i2jt3jnuvqXX54gDdrM/k6sWw1
xu1KssS4AypOLG7wbwdjAdioxRkzvHQXe0wAAnysGbD5GKMCIFW8u/VEo61ESW9uYDhch6CJ0uUG
yXpo9R/WfTeZ/M2C3U+64s4zDxfau0QpSPZj5kf1X/Ep/+Vqqk3Q6L279vP/8JByom9r3tJpcYDD
p3j8NGpI9Gou0IaF7wud1PZ4X3Na6oYHy44TcjGRqDcJFarEulyhSy01HPD0LrOK4PS+6DRtgWBa
cRTFjC+vUEZm3U39MSJ+1RJng7z+2DRUDvaIsj6GhbPWFpW4I3xhXlYWtk5q4t3+av+77ODj3kF2
EyR1mYjrbwgHUtZlt9WLJ/7vWPJDmTRpubaTWNx7aMjoNdKKup08/Ky0n3kv74GFTvyjeVQxAgfG
HB+wcLUioAp0ChCb35o3NN4W/RlGYBsS2iUm1VTegq/bTG9HL/xaibwr17iACfRXjOlO3CBKDGnq
FQPOS6lbr2il459sb+Q9D12P6vRIr5wpfk/a5zXwKRl5K1ZRkQDX9/5hic3AwVQxnna3hJ3Kaeuo
eS9/qiYhIe2t+vXAckJHI8vmwVl97vyp/V8xlZia7fkHSZ2+IX/IiNIJnhY7apFYZ5l4/tKh4Nm8
FOGK1cZe8rXRD8Qh7ysl+KG5gTYc7WVg6Y0jRJ5E3/08LVp53o5/grNuJ58L0x5gNgQIKhke6cXa
+AAIM9a10sWTzdRns+QdqgGfA/RdfLdljGqwu9qjKmRF3lLxg2TxQy3Fu1Ub36h+Xdo7LLhacpYh
hnEQt+AcF6AkCtHMsliBKzHqa3IE8ip1U9pJsZXbGWNuR0BpFPHtCYvRxpyl3gEjUGVKaAPFyeyA
+m/ifC3Vs9+hEUHkQ0aijsrFIPL6nctDAHI7Im1MS8EQTh87yKjaZZwohkzmvpii+cwu6Y2PUhxo
HPLqEVzSvGi8bMDF/CqvOQ7wtTB1py1ONW9K7g0g2MM6E6CHo3GYHxOBy2nmqNnbvGgEYvygnasM
O06UolbRk3zuTzVzxq4RJjfUVNmQcTRaJ8TuJK22+dBwziBKyB0X76pHf5FYThLXr6/L4Tx1tHIt
wQL2LPg3nFL9aWSYEadM2kHRbq0u27vVpdrk4YvAsO1kmKMPWXELjO+PB5x7svhv46jhj0D2NaQM
+JYA47w+YPBanqnzQVmcFigm12sgoOgU+A5omNI71eLDlkdqFLK+lZOx+H0hDjKGsHSFP6B0YNZp
TLGYXAuWv9e2ja4zDGI9lu4bppI0sqiIEcmC8lyisxf6UFWJVxmR0+ybKFe8Iqf+Sqr6Mw5Uz06t
9UkTJT1Ahwu4vthnL9K7pcFGkPJUtj9XNFrA6zDjoqoi5PvP+IhmkFunHWe3pM2lg27PsoA8L5jv
GaYiwHKRoE9cIIi40RFfwWFAkbSjMp6ZAFm7DnOde+M7dTdaTgq9qlLbTJk9U7kcbxTWKVqkZPku
makaNAq2g/AthMwsjiZRx1G2liujmN99ue7Enow6pdGEi+KVSwH4BGmsHyv5XXjJ22J7Bu20Id3z
0lugX9IcW7WwwwFudG7KXl/aw2q3KgqLPjQ+paAbkIHOF3M95Sbv/ifdX82BhaJHNesU5l6BXVr3
fm/gyFFWE0LauIYXrfEgI3CeSMsfIH4FAYfRvE29baYxMyc8tcOBhBAOfVJRQT0KcQWBJzgRQJYE
eA4hHCY0U5vTvr4v8PdgylVu4pouxXXTWFx5I3PbqBhOXlrpIGm6qOTrJ8zI0qrfUdpJSPj9EeTi
dQaR3w+v9Q0qxrxRnZD1g0wkyXTTOeVU9q/fomR2Woc9fdMIyytKpWLy14c+QkTFlgYgtFX6Isqs
Y+k48b76DzITx/105vk6LiBH7wtxk1Fl1gfK+ii6vTqOXwGkO+0H7fsqyZWgTjSGyLpeTxjFnWQX
QEuofRL/gj8E09GSZ2ynUHhP8HgKrQnbj3hIkuVWlN/EFsnJdBRgRNhxUHHd59Ss2U+OD6VQ4vUu
O0jro3FMK8mEzZj1ZNaebLKmv9vFJ6ZWnAHtOeym81TQ81Hz+1qu3ailwENqOZGGIhN4x4RNpbm7
eg2nktA16TjGCKo4gpJl9qBmGalV3SQAvL3ZEMbbQEg3JhRMiXNMOzExjyeEYH2Qvi7zckxWWNAh
/A5kWlOA2/9V594RNm+P2bMXWmOj84JgvVMdRtONVKZKtO02A2O9pdzHOftskyUSrfEiLdyl4JUo
/R4H3ngQMtB/DPPNcZgW2PQhira8D7WEiKZSeBGlm0PBUrpRRRUxvQT+8byZkiTzwtJS70KMznHt
18zozP/cJ8uQSiMXH2Kojc1BELGRP9/Fuhy7rarOqedSJAywGTveah8vOma4GUUZyd17Y6zsxMn2
W1PxDwEEWSS8NW/Sxo4XIAiBz/bFpdwk7yDKVE7fuS2/nopfHJLpAbpYzVowkWyoIIwbupanTbSF
X+jdyVqpodCZ1PMAM/+OzxTeZfJAqQz0zNHP0nEBorRP/1mqSIQrJyGzElgexff8/uo4lbqOA/AK
RrlBhefywoJt0bWOg1wCkosxkhqeb/cfr9zSjpRSK38mMDwrbdbBr/FvmjVTfn4j+j1KQvNSxCE0
7h71eEOKoX0QirEul4iBqS3alTeHY6PEOUkq3u5fTZJwEDVmA1uD0ewiXUpTLfMavWNDVb4NrAVQ
YjKxjVGlwI/uXDvSDu3O4y1BxlW1bdOhTwnJi8WqwFU5brWx5hSXnpyP5A8WFRbr9Nhyv6mspF7Y
+HzxWFtbs2xFYn8bUnxW3/r1ah1AO3lBeOqw8MVGzgt5sle0tePMap+WwScSSC7SLLARrxHmXsu9
P5+QgdTV08E7ra176c1tDpi2j3G4rOfLPsC1agxTKtJBANkHBSzLOauI786aqisyitbLdPLKL9s/
NZcKx3qUedg1IfT0som7p+Ua0y3GUR9fOxVFOHx8NnjCS6TJdWopdSOLQ4+jSbcxQ9Jfdp+JAXxv
SUBgjYUyv/EZPt+R//oaIFGei5ha0Q64FmC9eLe7zrtItPGy6cUq8ZDQ6L1rMZNFcyjdTDFvj8dS
DA1fIUGGRQjEeX2u1hJI0j1KNXXicu6w3M6rl3X95zghDWG0Vk3m1+hcK7jULuiRm2aTipUInC/I
1I89QIotERhre20igsE7K2fSQzhF4eSUJlZ8yWxy5hDwtu9fpTlwVburuK41PxlEPQq7ep4bIQJN
bW9dISyJ0SYFRf6pFy95Txnr8g4hXf2gptRMYylpwX+IFZXwi5mON/2O6ZpndUl336gp1VXY5WmE
mJN+agK+Jdsm9d54uet+zHHCJEKA/CLHMhOPfPzJJLzpIrCYnx90WO941kJO0YLBiUfklUULCosT
VOfChIWkZkGaKTXViyH60EJ0VWb1Tn1rKiEuAWXnjrkrxFnr1VodSppTt5rUF38ZPT52BO+9hNG0
sox59nTsKF3EYjsSMUmHmjomUakvLVLnkugGng+CTCpmx6MPPkY4BkH60D9XjSVvsk6IYjJ8Ms5d
pjWOXl7CblOAyPFs2ql/hb6MYMEAuKRwEj5OBgdIfHqotAgcy/55bDiv/l+ronQ1VkhTYeq2OfUl
O9S69GMFy2jQzGQOtufzyKZQJU277ptLZErGZDwzVzv5+JEn9W7wAXMhLvvvQymWWHg4Vu0iXSUO
1mW2wDtlJ913y7S7ePAMFiG8Ek5xzJBhj9sBF5D86+wmGFpRfcm6hUT/qGZSFjzfj4M5wowkuRCF
1vOq1eSRVyoFrjEFecF9y2L0vvXlf2exNEAR5sCpOrMUamx4Dh4jyFDgjg9kGuFKgWMYlGvN74uk
/obN6U7kSwlBH8rZGLzEkoUjwJDPaiLoKSOL19ANBDbaSWmzxN0V133BHTBcHeX5ldXPLBOdQjs6
6PpQnUFLFHhCOwrsqwQdatvENIr3LSM02R3SOGAEGSBrAcc4n3TGFNTt/e+oprgL67IkRmaUlr4L
WWAJRz6gKacqJ7S+Ufz2RJ+C4nhQPrwcL9dr8jfKktaXBgAXaveBqjWHTSiRPrJMtqd0Dzy1pr9V
9Hsa01SnSsz6p/9VavNW5ab5RSa4PuqC36aG1D/qnqXlUtiyieFfxXP1DKi6LMaILMDI2hYWRbhu
+2oOilMJOj8ZxMKJyztQN8wCAFqvtr0qNoScUkAeqNALOaSKn++berXq7IopUtRyzN2AEQuUwj9s
H/ngwnpA9a4Cx1tMHD53HANm75vBuK6JqDuzr4viGvFhbD+qpK47Po1iC4Ba0pC2MtF3kMo5gw5T
Ec0h0hW4Cya1GY+xKltDsGv+9Lfs/sJIGNAkmSqqp8uzwNDHCqH+dddDn9+grV9BuzYnDoBEqYUG
fPNmi3Qc8Nk4RpOXNVWcJJN1Jm6Drlbx+IVNze5pXvLJQRfgi5o55Ra3s+Z8+BMJ1AyHCn1UwalQ
fBRjqGwzJW6ZqBgy6wBjM3xCtU76RfZopy6ot+qu9yj6uulHQ1e3U3PxI+B9B8Z7To4dvxSYxgMN
D3eL8NMmfur2mhG3wKD0dKKuWWwRVilYXL5w19L588nvyGcs9OVpwbSZGyQJ3nviOJqMgj7y2EdQ
amTRuS6E53ko6PyhvefncYJtIwmBRK0CDsgx9TN8JprmuaAhP+JF94OruqNwuEZtLlGLRmOZIsA/
Z8hreWsTSOojUDrvL2Tq7fwkjUEOMs2a39Z8ZYQwRYiSY3fgIIQDP8WC7Zn5BfTL3aLFp4wbi2Eb
38c/ToN5I0N9RJ0o6jVBs/WZ8U8h3J/iYPU9UuNUaZ+qsQYxg9vaCOtVSqPAVwtEQl5lpGfcFld+
vnFqGiRXb0A2zhxFvI1Ux+3v0bJNfSzdagS1fidNZEEaNlhWoqZ9gcAaHprVHoUi85Wdc7a0nuHZ
m7/m7Ed2vqmqyd28HgIZ/LqkAz1KjNUCs/rFssu/YZVRU+OGe4t5Xdg3xv9iSjMNZKYDiIjwT1HN
yyuAiwy7oJCCF3JrGPfTzigFUmRRT5uKS0t1DWiEJ11nggaziHG+fDV1kuQUoUG4qtILj8FpA9KF
PTUOi7+IkUwBXUY7WszN3dDrGu9NwBLBiOhSvtnJxl1U1y5YSdaLD4fEHtiQo0IOAHYe9P+Xdbzd
lLqVYDImB00GcPn+BKlhWI33jkDC002cSZ49JSC2TiKc/s5z9LYoRj/nj/3Yoiv7gmEM8vBAppTD
Nf2JNe4S5XMNb200S+JmQpferl0JI9lpBkSwKe9p1OwKy8VwpCJhER7rZeOntzYFPjiIUFz6kdef
aIBXIeic53zsHdqBjgwLI7/Qrgi1xW6DcqwnBYTkvxED/WdMbYqRb9YqxaWB9BlTGDzSrG6JAd2I
ZWxGInTBcREcP4XNps521xk4BXaFxslH9Sw9JoW8BAQBUGf6xU4fdehYvxtZMKTIvKoHpYlRwCsQ
Gq7PyjEHH9/StKrYfVVckmE6VCJshBJCbhtT/aRpyVRojK20jfIjddrID9pj54eP/kanzfx8kJUM
prd8jMMFUm/m9TVYOm9tlU/Bq7YtN7ao/W6VEcwTpC1n5HaPTJIbyQEjwmu0ok03Zeh/ZU3XVLZY
GlzhiG6j/gfttSmrg10lUsuNaTP4sbtbENQ+RGuvy/bdxXODPH8JwqE6kl05cc8V8z7HQgJHRGFW
T6GFUE8iVX0nEMsnZ+NxjwUkOmxmi2Qz8PKsUJApCYpYcpQ+uNEfgnOkSArJot27l+AtbOBwSwNb
PBrxWDYrOBLL6qk1dWEbCalIdURiBfJG8kTbUQdXY1G8fuogqvDtgoNt1KlS20ykVhbLy5xZl7nv
e3AAbMlKLJV08Iwa6Sm+Tgo90Ob3ANWHornE27Iod5GJJrM80M8a6SSXOKCt8jJ51eU3vFSLNZs/
RoT0pYmP2/NWdB81rj/KQgNHNP6Pc0JiQuGCcEkvJ0Sn3WIIEdUhbaymGDaBeQIhZ8yurALfQY4i
Vc4++lwXoOEz5CUQyMiNlwBeQcIRjdUijO/JlmTb76sdVRSIX5lG/OG/OBlo1OqdOMnpZFLGa5eO
AWt7LcGJb8197kyopymR5qbvD0HwOZRDVLYsFU/VeNftVOmtn3UF43EJ7TgU0gM//JkPfRQHsfSm
sy9ELw1sFhk2msDxtrPVdZBz7izMW7v4R1yFRGFFdeCHGiv+pwreloUNGyVfDgjLBlkNzvYifWNz
pr3w1UntZ07sqhTKxwER0BHWI+aUQSf7WOtB2S/VVbMAMyRaSMiJUoFAlr0pZrlYdqJSVVbhZBQ6
jqVV1bzIunStWWPEunoi+tzQ8NDOc6+nFymd0gjLjmtBJ5MlOBMBBBdsn86SIdbG0uIDdV5xghCC
xFNqt5dfcMDTCFQ5xaZn1e6nReMZL8eaioh//XbvZ7dren62vrru7uee16Jsf9en3uTGbHrCQz8b
PtGYTL5D22/X8CELJT7Hps/5v0Lxa1GS+pX7DGa0AVegNaOQb9gkPwvnHEgj++W5ErIzqSJBQQ8r
gNA8YLthuRREKL7O+V/M3H4d4vW7pu+FHLNGLKcwb/j+SLJEKoArgi50p2KQ/Qp7nr/CVx7K41NM
nxKoee92R7IpS1s/gfyxSL5kREu+EMiv/8YxlfIqFRm9wrMWfIS2rBDq+qtbtASwbnyYeenXWpKj
1nif9lwUfZD30/TQVNXRCOFQB/Gn/5qO3KGkDfVV0pKGEsbRgKfOEfe/UH3a1rJC/0bMzafNG/AR
9FTjewkF0CCPfWZIMago8v2VkKgeXWLyfsPTUpfozUkhDTwfWrYgzziLY0kH0p69rjpl1kC3racm
SXfpIRZvnSO+t7SbjRwAVgo40dp2z1492lkIJ/cWMI/mNKOpzu2NC6xpl2jDphWlUjmId61Lvk4S
J97cktCNllCbWi30iyqMH5RNPVJ7YUtn6sNhpeOqhUUwcDqaGHDTxktneOMymP9pJSVD4Ga6r1Cf
jciCMwY9XcsiMJ/HiBBOqizhmWAO5/BIQshzcpQhYHFa5XxuQEk44il3Pf7AI3cc3EAC2LWRCfS8
oKI+U4QlVaRxkx8L5WGjNwCHWspLj8Vic2HyoSrjK99AH3WE9RHcgnW1MXaPtTCb1lW4p/lRmyR5
0w7Ofsr0YbRWk2qTLsYCNDh3p3gvDuTtrEEDZMyPBolvCXJs2SkPak7vfBYVxQy09cde4X9vNB9W
tLC2fjROAPRFqwW3evVyjTFjALWfjrPxLYV8NHKGiHv8Q4FSG7iyHx3rwC6fvG7nmlxKe1MJSUY8
3/72FtJFdqBJnlyQvquQA3G2fTic+IJiJkTj+rcNSxMot7R61I55SvMEqSM0Yr+LvPl8KdBIpLoa
fPqTK5LRJ/Hvfhv1DoDluli1pFVtuUIUzsjrErv8im351EUdPPdQvLDaaMK7S3dCTRYkQdjiHX9A
ssjc1ktBAjgRSmd5x2uM8ircHdwq0qglhRXX7LBtqWyvXGNPQJe+MWDuxp6/68IL2L+pkmNKnZJX
8TtyiSu2Q7n0WVBVwf6bkIVONGMWB9UloTM5jRBrHECMNMWpKYnigOkqD+3VK/UMj18E/8qMqSD5
q7fmFXHiQHXxJTbvKeGY3bsaTywdolo7EzxPPN+VVxqt1WZqfvY/7pE6GxA3bkqzVKdraNIAhCo4
t5s4qlBgIX0GinRQPOPCKlJmW9fNIszsi2jVun8e0XhRiFySRb4zBZG2CEIJxVVgfcTQm86Poyoq
Sesh3dBkmO2t9bm1cxmF4OvhqGnNMRE9XnR/2yVRN4/Npplj40C3Cif7/9UVnH7Y3s+JoJ/JOWWi
FBRk257TRsk6u/lIHVWtmh1e07fcA/Jv89x00WiyOomL+fD831yMsuXGE5IsZ8pm9RZ9bu900Iul
gYJZfTPoSzgcXYV49Qb0c1//TcOVjtcwuDgGDWoRwNrbCUeYNsxucN9QiYuIgkb/lKlFrVxvq3py
t7mSAy6pCFNqfMEeD6bVJCeCS0NpEZmEADBrAoBGdLZKjNFBHfrX+z7IQgrF54G0NEQmmBbexhr2
oBxMFwds6QEq6YkItVm2JbN3EWG1dGp8pPOU/XdNJoF8YZXM6X0c1RPB7J9+ZUh43c2r+OkpiOMQ
00LxYaGOs/UbQPJg5YP3mn3DhBRF071xeWNzpfzrwM8AHJdePh1yupbhEJGmKE/aEDHZljLYUf7L
eHOF4cHEzrTKZAYfBcoknTMfR52aiBL4XZ86SuLfYLTDS3r1V86MkLW4oFTN4WyGL1Wk2SmZuuJp
bIxiuRyqVCzlSKewnyQoelYlnu46IAfEZzysYnN0XCHSQgtJeLVthIoW4bEF7KIKoLrteGMaelN4
m3je5uSPsEvAGeEfSD+EToSPK78QbJZxjmAnkoeUCdG2u3A4R7A3B6ikVA23Plk9qCOY9Pwm1dt2
UqziJtORh+aqnj9vhIUqUjOVR0ti+peeWlMMB1SnPlSwS/oJQMbDrd8SLemZkKGKFj8AXeISkwUV
cbAttCYfGl/xeMQb6E8nNWX+W6B+vfsvtV8lQ/aODL713Px97ZGXSUbFihJrQOmUYQTPIC+ziRRC
s5UJ9WdWSjuyZLuUaUQkh1/EyVbmAZDVVxygRaUd8TZbDQetUTn7mX1UUoSV5FTWMSEQFIrfadxB
lzy6rPI+hg+2IrN8fVjKGX5e5czLEEU8oC/OHW9DO/rx1/1L3EtPuQ3+hFbNfzY8dW4KCOVyWdbb
gGt45PG8VU/vR1W3z/YJMLO5H1fPH546umbnzbsoUcwA4lJOrbtTwEIdz277SW+vWKDjuZOWOIx9
J616BvKlvxmDnMQUhOotjuXVQno5E78+nTVcAJ2SZrC4YW0gYaCaW9b2U182UbTX0ErFJv1+TmGh
GREAi82OwzpLjWNr0DJnj58eXaT0zh3ZgL2/RiZwSekAs/7cWaS6F2Akyf+DgwQBywiFXusQI+cF
Dq4VXyd/3Xi4A/iyOKcuRIPuj8QPDYyueTHL7lGfdx/1wCvp6bOWntoKF97+QVCzoAOQ8QCObSWL
jKDrRtsio8m17sO2UITvW1PvPI6U8jcRXmGs3WJyt8bHDckUbg5/Mu5wsx84T4jIU2FGx4zlkkpS
AvRJv/YGBDDpXX5GZstB36gEZ6Hbqhd8k+bByiQpPWv+vkjDPC8ba5XN+znSBUsixByAzmgv6SFC
erubxF5tsMOZTx1qQ22/ScrfIhgvWRXVbG21nghK064nrW1l/wA0f0brW3mlwcl6EusrXUi3Djv9
qDeMHP9DcPELFLBftA3lTKOjUE7Ie2YYLx1fgR8GKtVpov8aglhTfdWjizQfQHDkh6Kf/NPn1vKl
fkbWFsZrSSZ4wCiopUryr588zHyAmv+XJmt9/G+GfykqChi2lLqFira/l4br4Mmc5+UY0ggjpnU5
cmqR1Qrdq3AcbAJMX6aZSIfh7ANMKeGn3nVHo4XOaa58/UqJnVkhy6rBQFMsW7DxXnS2MO8ocm5L
dwkfON30bnnvs0j4fb2JI/tFntmxsnXpleseSw7iMR00Tu2sy5ryOH1+jLHOTSwWiHGNl4fnUO42
ybq6DnTfFWv0cCrah9gZ0aeSwhIQUbSJtNArVehVtvZd+ThXRFZ/ZGVIBwLhPttAtRy2v9m0e9WD
iwvSwVikwWkuEExpdgB2uqMx0yBxjCdtBsSffjOG3Y1Zog2lKKbAiRCX8efWaxS/PawFUgiwl4wS
guIr2QuSQvKaWu44R+t5IRtj7ic636JzTj+a3hYcVwpOr+vDmTanq6g7KUS/V5tJH+0WQ3rT5RuL
t8f3RLAio4zJ5NCGyaWtgS+zc5o9SUP7HCOXZUB2SUBhTA4L+Hpckln4H5yImM4sGhFU5bJJ3KcH
WwLew+6sS6hVf8gETMXPG59MLEDcwwzDOXaU2/SuxLM/ilvbm8C+UllMRXWAJczekQB/l6c7AE4+
9Szilw7PlV2RcErDQNBkTY++ZaWm9UXYpwiy0mdmvP8BkLYxo6DNBoox55nHi72V8gMk4eGJ7835
A4+6SSvbADmc1doN/rzW3BIqAKZPR2YAtCJpyO8TXLBreHo6jfW5xc/eEmU0jESGBGqwAoZjKkfV
vQ75yo36ekLpHPJqrVwqiSqlSdSLwFBJwhHw4wDlXEfUNKMTxjids13NZkQSJWfQqYYJ7IAtmlh2
Cso/oJnsQdL+j6nz0SG6q7hdg4NqRANk6AcAfEXGDsOvoJtxo8+ZnmFkjrKL40p0GaCvg105tAI2
tYgfjXKadsGoK8xPHEODeHpwnizCe0HpNCBitY6PZ2kL51n9UGcbqOfQrJWM6Xd8pNYwHGyBxfxM
PPOiVRKwU+FgzYfYUrWWihP+I8CWXMpfdseR5tN77SvYKk9ugjWm1pqQ1qKl3yznHpUEnn89XISE
yA9QhL035IZ85uPgY0rAVjtA6OAVVNXPdGcevTUBaWBCNSitfgUF3pejKCE3vJqfbBVIYI0IdZru
SSbFGTiIbwwHYbucaGu75EjDLDJfdiuTidKRmabH4OvneFLBnRAvAw3axOmWs2cih4y4AyQcti85
Z/W33j0GnXuHAb46ewT9gzmZIchHAQzF3voHMRkIajN3c35Y6f8nej4WXt5stMHcB3ueWfMP2gRL
M3mr1DCdniK/GyuCJfZyuUb3/u2OapbTgRkNB+tmTlkgif0MwKOM+LiB9WyADUEglfwMKARGZUvE
1hRqLiS78JaFYKE1M9OM356OiYhC+9Kx99pwba/uu/U6m66jie77GMIyCT9ljSkUrw51O8Ovqvem
b0TixCSSgf/24sRghDTPNSBzS+k2RP0Y0j/w8HzvBk0zLeqPE4WKcD67JIJeGQKF6GmR18X72LDq
zEx37PVVDhs0/W8b3Y9AOAG1JIlyy2OW5g1jET/zUX3mqdNQUyRfXp/5A2k59nH3EvihqsoXHNW2
NHXjkSXNqoCIgycmF6yMtQ+QeOoZq6d/I+rjNyjljXiBbUkZ7YE4R7lRQWk1JI9wQFL5Blfg8RMu
Uy4lHCKstd/19bnKUpmmXPomqg8KWb/jKkIHCB4o8vp+7olswWvOw5h/D0h22f8SwuQ1trEGWrwv
MS9JFFnTmdKAYZiMtOfbZE2I2jWip66/BLDLIovG986al7dVmpRmLto826RJhb5NDvO7NJrlvPRW
086Yhzyh/jJ+MaUxnIzW5G6r/zc5UU4BOb3QaKq1zYmZPFYunY2av7ABU8tlFhPy/wlBcI+GQ5bf
uM3AiIrxB3kqi8N+w2f0hzoHPsbYCUh04tw08a03R9GB9K3NKV+nUh5FgpdCw2PVIuvhvSr5Myux
IEu3iygByUqhyL4eyZF8UqpWRkH/E/vOQVj3nJrD7tyIXH07atgeOZKKI+lIL+cQoT8opi/k/vku
08pjA3usau98tYVKX6GTKCdWPBUgrUupq4+jioP2/cKyVE24SvdlOS66gBaPVpr9HE4QxvEFv5nN
SGRvPS8Bfk77DEZu5bkD+ehP5K0vpdRMlFuMlZzJB4QmE1GYHrlTOapQyHohq4blxoFbtqjaZP1A
tdd2oBbXAlpi+w24HgnlYuy5fQPy4uPPZsSIo5WU5odUb8uQws4yMtV5GKNug1IkVnKvSk6ad7I8
AOd+aHdpmPVjrbXv7QJwTIIGcCTfI/w3vmXBiqA5j/XvYVcd4vft+yqQYcuHFiokH5W9iEd2bnAv
NotMO54jnW2IqgT8E9fAWk2whYc2Hk/cAIJfuk0yRFAldxCjqolYQiFow5SCmA0IoH8X6jiZ6F1D
rY+lrSUtvVfMIr0Mx9NPyhAC65AZNgdh02MdstyoaGruesvvzA8PIeTt2wqSBDH26zfz7gEuTNdc
DvWHmEjsT//yM0iukwxRK/QvfWTFReGu+s0+gmwnmiUtbXToTEfkErIcDKMVx1Sku6D9mAnt7G63
Qr7iiGNmBVn2jHhYJBFI+OVyTuCTsGmhkNf2IsqjNEDTSCXCXjHGl/VCakKW3KyLwUfXOY/GH+xX
ZBUkgM4avihn0WZnzRlra7K7aW9mSpGr3+r0TZfDprpPJRJpxGRA5ihkggX0a49DGGL9JtHQsGha
mrthx3XgRjOXNVcegubTIikZXB6uSFjcKEmAtVeWckdDt0L6D9rKYa1I2r3qCwVaoWEd5QOIR8iO
3qoCxVjQfXMNZokwY5niHEPZ66zf7+0xTjPnW0hb9L+FzMnSJWlicpRObYAm3+UAWy2g8XIABhEn
0lpUFUcC3JGFyDKp7uCpMdSSlOn+RDtB4VU6DKCBojCWkNEdg1ub20rkdXYaFEgPbEYqbDHqw7MG
BaK0BMWziULbBlThusYOuZjEuE7+BTkj51bNivjKYk/EzlRyD8g+v11goM5MNK9MfqixDY82Dhhz
qqA6A8mJJHIcAzZXAtFpwXQyScoj4wNPWL/Tl7VoqOUuBjdGKRihOMkghxGDS15rlpgCrvJ2UZAK
cE42FXkFoJdBg+aQAliL/BDUjrWqhdxbqf0NKzAo10C0tQCFdr2hiWfaYF16vQSLXT4ZsZ3LJ//E
6KLcTbBPkgFzzIBkcnS6Xijg17jRgRWBHsUaXz6d3StTGNL3h8yK6LJXeDg9HWxrqmTjc0aozqk6
7GSLyaUfPHlZZg2vNP6/VQMmXzw6T05+qK+lwnE3InEN/EhHY0prKu8gSs41783b8ON/LZfDXFba
H1vA9R7oX/bzRFiVdx9zLnbudifDhrXrcqpKBAaA+sP452JerWl3cMnFeD3/z5jGYVvSEr2oENyi
lh1JRu9pICc66dayvRKLM09NxECVoNsa+9z1eCYvY6TgG4FTD+WEsyZgSHcDthXEns30MdGF2wyt
BNrmWAGOKBZYeHAsP2JwuH7tRzBgP3oirv3pbrpGX4Y7SZKS5V2V8cGfTajEkDijNhpNoS8DzYkG
mpbJEjhwVEHV0trbVmM7Has6k/Gy3OLL+oHr9WsenXIbaU71ra1yl3P6n3Wa0QU1yJf457T/8Ktu
en1vt5akDaaPCo4ue1QTqJctMWoXEl+O5GsFYnv+1j9Kxjc6p+JjRQCBhLPm9HxOMKBUTR0SLbok
gJYmVEMHOOzW1pzkM/p3OaWz8cuMHo2XfsgC2sM6hBHqnX3ixG3Z2rOruTHWk/1G14+Mq9gEDU9S
yhkuN2HkMc5VHbhBDuqGQkbMCweW+2NXCtyQb4vqeBmR6cnuJK524eFrTyfgqkuyDwhFY/7DYmzw
0q+iXCkOHghsk4rkRZvjzzENSPjCOizYeKKlPbKHiNQvD0o6LOB9D1BNjg7/enWUKppcLFi4NBan
apkKLehNaPdWrssbQ1Y3gifoliTwefOvx/gaOhjOm9zi9M+s+KlEMMX8XEc75/DfWr7U+1QyAENv
rHjqYev0EVly3reMoe+rquVG+R3WWVBv2jcAmekSbp85x8228rKMvvSSOWH95P7z5mDsOdI7cvqU
u/PlpoJXppxZHs0E6xH+1q/uOHMeuWCEglQNT6hzordaJgAA6tu5ZjmXWfQ8pcMqRacDb6hLpbSN
oqtvOcIRk7uqeJltjwQ4vcWc8e1rTy7ZrkedtScDKR0cLfGb4exvXNzhTR53U3jysLBItIKpdtgC
xuoDDRyUWEx/6vwy1eNeBT/6pVoVNqrQ0vlArLR48dX+Unhd4yv2L6R5TaVc7VEhK+dBjYMwe3x4
RRZn8e5yuypcljSi9iYLYmoG2sV1pXMuBLvV0+T+nJegqycR9hDnFCLFvY2y+cHe9GtqfoCuhWzd
O72YOr3w6aCze/WxVoLbYqA9yr/7752vWchFx43a2v7+K1EqaKazS/ajhD45C9MMhqvbWMmg1dfV
zP+Ks4I6bHTGF1T8j6RjtkSCRpRuuJGTaua3u4MZSlq4GwNblH1PfE19R9TOv8jx/Tjh+XiGgHdg
IX2TGbj2OQLO+SsLPmMha6md+dzNzsi3gjeoBHoolHlnAix+RW4CbRn1qMqEIlQT59/NgHPLh5Hj
rzS0lNe65sXz3wZhnb+SX89hNQpl/bzTF/LNaTsnvmyV179vANnhjGTOPlTo+nSQu8XEQXq+d0yH
cIxu5oDv3EgmVUDw3zp0hINq36H26Jsc9hxh1/F59xTgrEHidEUmXFA3PIpiQ9pdOqxeFOsBgzWZ
MJGLbagfvfjjmlg1hoc0z03Ez6CgzXfLYr/GK/A4KCZOZc1BZSe1+xssOSpU4FOmgwly1DiYdhS9
mYmsgNWJmEfW+l+UhFfUak2+3fegbu0Jz42AhTNDelAwd1RWxSnFpbqjSOc5fgmKDE9dOwU/JFe7
73ztDzMpBxeF+dpqggzQl8EIru/0VJ3VS8L3aB2oWmWpmhmFaehyKM6yN9a+iYJrzTXsIapme+Z/
m4/2Kh4qjkZcARIpoHq4tTBjalMF3x32JkEC6R0JLbWeBG4cmWdaC00WJBWmkT7Z+cqWtIE6Su1x
vX/mHxaiu7+V4iqPwdWB07oHICbCriZwVxJ/i3Eq1/xNqFBHl02TFlCJ8ANdWr0AK7wN0ScdiXz0
vBpgI12CzmagucSKNmEwtHH2TsrX5O277AwTr070l9T2ojBCQZ4U4kDDiMs7devi/bxagPQai2nC
9QnkPTrefxievXh7t1bAvbsuyWUCYBMNIJ8ThiyIXtPNYEAaIh6VpWyd+NRnyKXLss6y/lEAKsDi
bBlfBAGxvGJgq6Y14szW+tJ4AQR+cGUqb6XrCMHpMHiVwtGlttasUpK2rsbzR/mjqRvLMPY6mcwD
/ie3JxEE3gHrPz2METVfoLSXLA2wgo4NiQTGHvA6l3J6y+aUZnToRCHjWaed90gCNpkJzE8I7mil
orh+mACwu36p8MPxfygSe37o/qPXeejPyFBD2Qrd9dhyfJRbrv/8i7Pkbkxecfs0HTPrJAaP4cXM
ynvBjSlvqZMBhWTn8brCw3m+9mQAsHxbMuYh8X9XtlHv4U+d5/CgBMT6gb3YFLnI0HKeyh2RO8fX
o4E4z/7/9XXTP9qNBIfmFw7caWfBFg65a4vAV9uGM5xYMj+o3vJTdaqlmuwP1PPeBBjbCI/IYgSe
nAo8DoPIHX4dq15wQH73gnid66CFhMHMBoxj4xyt1dUQLU+fZ7kV8jC/UOHd/flyJ8MPswqiGbSL
qp/7mDg3VSa9/5+t1/fYwRr05WIHNlABXVUXMDx9oygzAnoV7Rbxq5LaZ0KnDnbI6QDhpQsiLWLu
jZW26H99cnyWLuc7LG+nIeX8sMP063f7OXQufcPvEfzCMyNz9xm5Dxc84qNIirxzN/BdfRek4s3f
o1/3wj0QgFzjIOU4xroDrzapOWWyIeeCjVhFh77V9LoxAQuyPJCkuMweBWsqf7fRjSOHr2MX8eCa
anaHgOBIqW4lgc2XH5YW08cJVULeOHPX6WhGSQhoJOIgZGu85oixD5y8rwcG7ObqhE4w9yi1so9q
HQcfxUCf+CGmLrCs/dR6KC3ZimxaIi7KnxSWta+sZXxQMcSiviPOs4lv7Sq/x5c1gV3MtSCQo9wS
dHsxvkiNY+6e24OWagHqhc1OXSVjzdBewAgAIXSJlFkboDKiJvxEoCaAXZnKSEq/Exf5k2B6x/1O
OjzvHrhPok3OrDMe11Kxr8CxWw8yzpojKOp8YMubVNUPNBhfyzArY81Wsh9nLJ0xtti8eWiK9dr6
B4o09LdI+20rQ7HLsuWpAoHuAP4qfH2CmWDwoWzRJ41t/UoJi24BEbQXGiQHHfr4vo03ypnlPC3Y
sRqKBw2go0SICIw/et3Dy7Quj+AaFcjukFZj/Eb/GQRFjMkOdCzraAaWtdDHxL9C5UKCsnmWIS9t
VO+fSuP4xyeIm7RUk/k6nngho1uyAgwM16qAhBAvNSNXlve3TkJ8nc9ezppuus2eiGtZ4kfmqiwO
Eo9kgjjvf637LBFfpJ1gSgXKwWBUpM6a5NhAIdnt7KdM4QGV6N5YSpkFlIOb4a7ptZ8vGFkRI4TG
qq3eoDZGhBDJPZ240ecfL6+F8wZw8Mg4ugPSAC7hcfBzUGz7C/nsO5v2WEtWMlkM6LoaeX8fJ6hz
PNv8syre9jyOC+4t7+ZtqlvScGFSujKxKkWL30HQiN7lPA69Vu77y6r4FVMn1DQUEMfQEhJ2NgPF
jf6ZimUoR/G37CKQ8kgoVVU9VLRtTPx79qpbh51Z1EqcY/04G2S5NjMDpOh+klt1j5f4X7cLjolO
X1GsmEu7gnXzr4GjSpaF5mZ8Bal/ZNZFrEDVnnCGYK4BEPKPFbrfLIlbe4MqWbILrdmNPgTkiAKD
dv24j9kQx5SBAZfqFzyVF0fmh9TmEJRTi84drALikf9CzfkH8mxogAtRoHPg62e/f4UNlEgtWjSh
9W0HscEoNdctvSBOI4IxXfpmcoeRnIcbA2ysfPhQOzNSIj1kMqNkgBQ848hvHN9tg7U4QrBivpgb
Ow2faGv6MTLoKZhiY9Jzf4g4psb1ICoabOOAO2VdGyrOYPJj6eOpJJ1pS7UW17d9A+1z//fghklP
6SmfG7Jwch3+yjjXG1Bs07RGX1WG1PuAd4j8XWDCAFq0pIgmJduxa8FSfdJf6Tqs5x2okMoijZEf
dAehMU0Wi4aQGHnqez7qQ6YeObwxHs3IExThkZogQurn2o6tL2nSY4Qa0ArWIQvPtBUJVtMnjyM9
65CnzI68WH8hRvih8ZZX+IN7Gl8mix68+uFdOCHodwGGLiDyq2n1E9eLyrdMywgBSQkwXCkLui3j
yScQLrBnEUtFyf0HS2bWtDt9VdKJGbNsG5XwUCLaEMrb8cVXmOvUAyUMrL+562cFpQyQxafo4fVf
eTPspptPprMXq7sQLklWDO+choN0XY41oQid0hMJmGl+09kNMcoKC+vWmqkV87ESdvApB4tjGj9+
Nu5fvEsKxOPkOkYcZG4reSzGwlBmTtDDGQrfDF8PTVwpHt21HZyrFy9hJntaXJWM89EezdsI1tTh
gXTFTiaG3ttU+YyL5TJxDA92umkOd/TE/N+q/0vECb1MUjWegaUEFymzb0jG7DTIlybHwji+7WLt
f/55foun1wULM/k6Y7LRB1c0zn7jAvo9eGfzu9Sk+Gdb6VVQuzQCdGbaotPzktrimN2u0WamNWRa
s3tx2SvAr9sJ2VPg2XRnv0besmORjxqXuR4L1/ogVPKcmqwi7jr8f51g7sVshXm1WbO4tO2Q/fuN
WXamCWkO8sxsjuHYvuQSfG4gazMDA8yoxlSQDz96cimwt9PA9FRxpZIr/kgHWnBdxBZimO1UZUFQ
U1jCKQgHCfceTXraRv28weF+KmC1zlEjnctiTk0RUX+KjzPUJA3IvwT4Uz1TGCwkNoxT7pUXbWat
IR1hXYk8g6h2wpWpfMwRabGP8g1Q1zGvjC+reZafJn7OahMDDqWJGjashwwB9saN7ffVcGKvJsHv
eW0I4vBF+JLMKeZAyDSXFEZr/9itqy/dvY2r7/NH/zrP5zmo3hzKN4i2o3IL2SkG5o/SvPkxRVbi
dDR6c1gUiG+GhuGmlFrhFicTOy27brLUigbzg977AqaLRBPukmhJt+cen4zVHTAVCDi+WOUXHj4K
NE0jxNzHXNgwN4mNr3iOHm6IS/TUjs5g1vqVQB8Y11slTtFYoR8YndFCCiAWGOISnnKlecg8jgG+
VmLfUIpNJRqXIJ1FL6j87hyc+2RxFgYe0+hCg3YAgQ6wAA0v2L8HffVHzI9rISIMKjzN3QrlWeNU
OxpUvJRzOvJoOppMb3ZgDGwaI8qxNKCAXxxi6NSMvGM+TAMiJjOkaol0+P7wrgGDc/ux9oME2/R+
YuCZOLoJefl+MMsZBWk2WQeI2DlZP+H6Axn6Quah4+GMx8Z1ABWjZsvQcBTO0DRsY5/v/fg5/eLp
DJ4cqmWyR8lsD0gZYCzp02Y9j0/ALuuquu9D9PynpY4LFpou0xjE90OLOIuwMPQTfIfxo9zblpLm
ShG+Ht7BBWVJBgPKLP8W2wpOoE7Zaws+HoNKCmHxsOCyHbD6yEEAomxUdP1Zjt56rBlm6eKoLs+A
pioBQ26I4TJfsPLxApw9ySKKOvTRZWaSGqiIuGkTRbGa8fWwhPIAeRLlzFCG7XIW+4flKc+Ak9tZ
4nFoxQt4cTMzwYUXx3NzT0ODvP/+QnadIhAN0iV7AEEHRD689u4HQc2WVURU0shl6/i7NgQ2yMKN
ILVp5TQIKz3pVIKjiNXvyKzaozjgEsHDwotjXrXqvFUzwExJ9XTYZtrHvt7o5VaePj1t/fwo2S/b
j3p/Rw+GukRp44fdnsQWTrdb0fO9U2dcQUBmObWu/E53EKeQo16RAz1Gz/5iZkgi3rG2JIznmAxQ
fJo+sq6d+nD+iVphCtBARE6I5aKIoIblCV5sNTmYYwMRkym3igRyOcAdsRUIWnz0bRREWewhnVcN
eZItbeybqehJc0PPBOYYxzTn/Tcvk1QcslZRVKaUQlA4lWM5F8Zc8MiU0lHqA8J3fBYESwJDVDVr
3QMuD7+UuxfpLSBUnp9HOr7sdYVMf4PBT5xMdcRWRQ47xWJ3E63M0RXxXHANccTLIayd/7IQhjxx
icgTRPF51qv1ad4zwdiTA1djr7rclXKHeaIo40CK37OkXXBSIzvwWdfJEFRbwUDHyTV75ro14iFa
dDvt38UJtHUF291L10RgmzrcchMf35OVBzjcOUwYDqXAcAarBKyzm/x27wdAZOkFeX64/1kSmrxp
5zfzOo/PDBIKDi+RztNL1LmAZmGcmP1EWtvsP6ncvxlFaVAWv5thr2olrhvZ/uW5fs/Ne24fGRTS
6HoFM/py5XaUmCD+5V7O4VqWJXorGT7g/jYpARSkkTGk0BcT1i/KUL24tT+sXZTXB+UOMCNxrrI2
3w4/FlRnkbOKQ0P/r+MBd81K7f7Pdx4NoteowUPzsn0x44pkQIqdmaAsDRdIG6MSSpq7JE87YHnf
2rVlmUJO7YHfO6tTmawTmNhr2hNEauvrsqx84ATXp2fCgy8Q6rkDVpHqYBYEyph3iiKWKZTmOSeD
ste/Z/v2E9iS7vPi6lBIFSlXItgU+ax5nIz/piX2KrSeY6BkkNumm2CJVTY38f6Glot+2GniIknC
iQO8aXlVVWDpYtvqV+HtSTZi0cWL4Rdcs2lj37iIVfiZ44I7J4+1PgFJi2BZxgO1arhj35UYrnGi
2ra2F1mkhEB8gS4xTLpbwiCvXFPUnEFyNnACY7X9QeSsiXQUZEZ6RonNxhN16OZkpcZ/GUtd6Xrf
DzQmB8HpSncCQzzPoc+vXMTue5LviRXUPgSXzf2DMqO6C+FK0hTRE/5olWGdzbRUvakaSRjUDSTT
vse5rAuHZ/PLqeWk2rbaoHRK0g6nG3NSVxoUpCu7VZ/tNBVSgUhzeaOuLYWkiDfyrzqBYmlk25WN
pC5jCvWgkdb5R9jhQzqzmW5TCboIwtfgreZM9g5x2+nKwuDomftFrC38OLENyn0Q+W8UTPi6D77L
WoqBY3ZFcLr2eEv5WmCyg2mX7JfgwNe+vnN0eAK1XRc1+U7wEktAfxYCahaGJwN64rgoYR6ICuYZ
nqv0h1oaSTzEs0ztxyyGC8WRb25WGvKO53EEnc4bhn25l0Z6m3u9DDpHVPbiEXds2yNf7FRUe/kq
jjt9jFtOcOJjz1Hm1mdARvYlmRUWlD7U9yYZUOYax6e11fj8Hmczn/jvHxfVUF4XJpiA+AMAPa0B
vWiwh2CUYW0H4waIIBAA5Btp00cDVhqdTiw23EiAKhhuaiGGParhoZkkkhaw2X5myeKhecVLdvG+
QEW2YqqVu/mCYQ3gBuDJBrKnp6E7ETLldSw+tyiwMnlvdkOF0J79/RcNAsK0bf/6yR3REnskHnq9
6DG61xP+DiEX7677hZN+Xkt1H+r5WHZQORwNYVDnsnT9NhaBCElsCdOWFmNRXCuX74Bvpbregyxg
yguluoTdb6TrhFWNUX8RuSXFSi68PoXnQOyhYbPEObZxxgQybIPg/QgQ7PVOWH3fgYcA1jipy6k9
NCgxD1yRIAc+UmTIWM5OcR4pVZm2wTWAtt6gxOewQsT2iWNpRcqEa6Mb8Qv/t2kVUkpaNGpyJ8+L
jdGzC+1Ebm9oPq3eTqBGIuynjeCX0i48qHV2h28sbwUGNdu1r+VJbFfb35yL39JWHjfLAY2kkNOi
lMmM9WzX8+UkQcQIVhINKIqQY0c6FSutd6AskHWt6gWH22MG/q1ZI0gx1Q/30MSFbUUg/3Q1qUIT
Z9GYdjUcBvvVbOIOLllUWCd1qku6iAO4uTR8DSgYHQcxgWhEWorVSbUvfYA2LGhmaqKtbgTlTAcd
XolnoHVkTVH+OBYicpEG6kIbvptJThzPLwbKBkWE3T7Oz2Zq9u6aSWgKD/LvNyusmPM/0m292UmS
1gwdFW85OpUb+i3Tk8xDB/2bx0yM6xDjgevGajeEVAFIsZzXeTg3j/OII3fpljauB1tKx/u2NpGK
X3PXGzBMiskdJI0Fuj3YFV8p5ZKJQsN82DPpbwEn/rSm/uQfW60VIsCiM6xNTrsgJl8/U0iXOjMW
HETsM128hS8YFKlrYDi1Qw1Zpx9e4fqPG8DlID517HFLj59fryrZsB8CwtLLdOfp+/LET1lVsXrD
LmwmK5x+7Zy3yObJ2s9x7IoNZtae1gObkhCnZrYHeLeBWSbx28WjCjuPV7d/ngBrD/UjaxHKneJ2
0OhGxbtkeYNc+QzuxQ8k6b2aMViXWxsRR47Ljqj0erwEOTa2JVJtYMQmECfmRRwOIxxunZtnxWrE
feCugbzeZyg83dm9FL8m3rIgtIAh/jNq+iOyxmKbOrZmgz6B71xmi0rdcIpE+rviylcqwsWjrB5Q
+dmjEDCRmWX3MnIU2UUU7yOIU3Qwku2chYdyKU5dLkoyQPwNBZsltPb0BS2GRvV7Bq3xTu2qIqfA
LDa0mCZARwQbPUp57ypsKuxmx24hcLcddEiyc+y5BqxQrZPaaD/vpQvhIHO99/xBZ+EQzJ2h5/O4
NdN5Nlv6du6hE0OXP22hA5ytbx2E+0MDUi29B5Lg5deizQggBCoErkVtI/1dXBqFu93Yncv3Ok15
tCVJDMlEqSU5rPcpqOtr2n6Q8rIf/8u374pYYsrJOrnx/pXzq9rWj2xCbZHJQHd6dPXqcqg/BZXk
gxShmy/KzUN+vTWaNtPnug0+QVNPnWHwgESrcFTtU0i/rIs5X23VTB1y5NUqVuNW/aauzPI001oh
GFYBRDGMtIAUqJkWR4cPy960NK2pz6qKDNMQ6eMQ8YaeHUd8c82apWuSPjj4SJOA2lWWMfTTu4z1
rjYWN/vsHRfB24xwKOWtQcP26o1E+jNj4zL8oeMWOO2VAqaQ03Jrg4fERLIKpkye8/ZVCppr+I1g
yD29wrKR4L5Ia/WJgbszqQ7oBhfD93mbkn8Z0zADegbeURgZsz2LOHaYSwiVpiV5cxTl1adVqEoM
Q++UPoy03Yzp3xbDddjaZnZPe58J3NRMR+ixWg8TdtwEd4MrJvTc8lGGqJbNGPH7rSYBcJivhjdL
X3gPQUF/JigMjJJ3ao0vrBis/D40KH7kBHvKJablAVgA27M5V8cgYlaPNE0zpIpM4eNdwa7Say8C
amIg+qBPMoMIg2AGTKL43Jx4W4x1MhXfBRmX/Wtpk3j8Eh1tHijxQqA0C7IRIsGqgUB/aRuzlDg1
8up1BOE1KtM4siNLLxjReBoYJlpye968AdxR8s2qJTI46c5h+OxvezYehzVr4isj9gaI0bLdoqJ4
cULuq1ks0l7xa6e+J1ChD1Re+UMCV2b3wosYrIRgV6XjsH0oQdSN6kStcOnV/iE9d6OoW9032KqX
klNxeS+q6MkXo+wIsRY/BCxcbRpRsnuBa8p6gxvhHreuBPRK8Or2vCMadLsIZomlkR7MkiLuhxYQ
el6ztlNvKpPE69PCvHcgzL386bXTFVFLBS+PZ0a7xZzdHDFIe3rDWyS/nfgzPXxfyZAkzG6Doc48
nDdgcLpQLrub28qXBt7L6QS1yxErNk6Sn1MLIvEGpA9Hb2wDexXb5EmSCYjqgX3QuRVxf9RTkVKS
MJKO2zRLA7w+a7EvW/GBukU5/qJ3OOhCVRhsdkzRH/SaFEmS1K65wDCk9ZNv2T7E1eBsbIMo4Z8g
t98pA8shlxaT1EJ4iiURUl96WolKIWYqn25WM1jeBhCdoe/tkeaaDfOKondzbPeI7LFp2HKMg3FO
1J1ckvk6VgEUigUnRsG9ctQ8Vn21xCTCB4Wz/JDMbDVR+yi76XANwv1yhBfoOHjEgkENXN1j7LfN
kAxzV7eMrCS/UgBIQtuVWCg2xNkr8rHZ+tVwQHqm4y1rS4ZCuf5YNuKoUQPgoshLCSv1g/nYDM9E
HVfjA90hV3LXin1+UoFBp78vHkcvH0chIZGTBmMmrFnlit5LJVhWAEOGHVm9bd9vIjDC7F4G4jdt
Xh5CJDBaddgnatDLxAwKEbFxgtwz9Otnk30aG/Vpds6/2Okaa4AjniVNu0PDay4s7o8vWbdWW4DT
GCp0ZKpj5x6GMvYV4tHICGYK6OywjwBJACqQhJ5HVpkhZra4ouUVJATkeHCE15GLnh9//II9Xa5e
vm2u10NFEzCyFq8P3bK7/5b/igyum8g67jCl45QrP74Lx8K/5xozu60oIJ90DP4btor+olv2nIWr
JxN2mPSi/fAhbk6nTI+kg0O9SJj+Cykeqc+5C2+0Gb6joZHYKPub7iajZxFYSYEC7Qun9uN9C2VA
DoWXPdwqbRI+bkwqi61p/15OW32EkpIaK8ackrcF2jbUtPqvXoPXGEB5kOMkmFaNIEW2zN8fRSrC
8Gup0wriIdLnYXD4bhaQEToBogPss9hIuatZ7mONVHcL2rVLQDeTr6kjL+qQGieDfGg3zuiGTHxA
EA/4zRq6Q1jGHvsIi5VQoHAwBPloneHU/GOsWudQ/4LcpkEZWFxzL4QQphC9odpoStosv/RJklB1
56CBa3Ix2b7ybWE+I1HxsJyN+4jB/u0SNL+Vp/RXIkm8lfodYuKc5zXKO8uJOdQ4hSGkvdiRKeh9
8kDhuExa6IVhB3FYcEIAyDk459E74rsa46STyULzgtrEbbKbyz/16LJ82RnurCfcyBe0QK2j2mWt
mUuDb/ZVjiMHocvmZbk+7spc54tWUg3Tly9AyvrH7ueNSgPpjbqIjgSYwOqkb6W0emx34fswYh1X
rOeMSFpGFOcEUc5RfFkZXe6dJwb/9ba2+0VadWGLkfLGVl7Gdq+siuXlJi9CRSVD3ntAgTTKEW41
KJNgNJsMBKy083L9Eu3fW0LxN2jvTNAhgs2QfCdFEZkDlJSAGrsgGXdyvAI1iHF0H/HfywPeQOth
IOLdOxVctv77CpIsgyxHcc88cKnbSR8J/9vGKL6vJzLMgXNCdnEKaUghhM6ddO8PC7s0yWKPBVl9
dutxVRHTOzvezMbw52LAJ8l6WviYeh6fIq4xiiaBD2Jm9br+LX+4OaKvQ3IHV6rX37XnFKBOJoqY
+/FCc+pMTrgZ5+UcDitRUBn8aFdx+v4oBx+d9M+bOxV8vH77DSJBawFrFAhkut6X14AYDuLfgQAC
pv2BDEEO+33aNx4IwpT0+ji9a0VLdjpSK1OgrHBv/1UR+AhPZB3bYBYqbnsxlQ4nyNtbct6EUwaE
bCh+hPKEjveIfHIrt/sq8au1kEH9I5tpBh7XFjyWtGila+lMrlCjie6THNroPegYoWC6ABP4dQuE
blRUJWirDyQEnJOskYkW81Coi6MVRWNZhoZmKnSg1wySqpP/Oy6+X0zMViEsE3mzLVoTIj3EZ956
wXfBktJF3pN3CkLtNEc/6178N4jCB/iHgOfR8yHPaaX2r313pDsYoI2wydfRjhnVFBL4ogEgzr5X
tr2mfefZZA523L/tOgrC3q9g/aD3YAEVi9rREpCbnBeJcgGp+vPtIbnU98mT7pFF1Lo9OSCwIJSL
WPo9QqziRYxkcFVdBTPR01xPM8y4aWCY4l78CrsctTgADPAnQBxTEribrnt+h8f09VglT8ZT/g/I
J+UENFDxFU8IVYNFS7eyB2Tdb8/pn+NEQH2mDIlrc1P7KaoN/OnUIsJzZDdi6OnZ/TJjWrNwWWYP
2jOBv0zqz2l8wvscck/7LlQVQGNcz83rjRmWGGooVdVU0tqEx/Hvbk+tgb72tC9PJd/tSxs3ufrh
q88u2FTpqeivx9oCTloxHpSrTtsy56gUcTb9FscgyUDSnPfinTIWdoRdPczrBNo7N72GExKxvql2
W0Gxj7Bg2kjFVaBReKIia4LNAHiJCSXYp3ueJ+CgZ2fEABs0r5+ihd6H6Lh4EzhaW0NymHd9YTWO
E7ueaoYFkSQD1ok6K667Jkz40SWuzAf80Y0VzzFFm35pjQcFABPwR63z6BSGJXEwa6bafdiOTiiC
26EtnhltxB3y50PHnv2qRSMiHNmQoxxsgZRfl2CXs/OUK/mAZFInf0NeZiH4dHu539CalUfSe5tc
8rqvBf1O8bVcX8jY1xpVN+cScu7tGMITl4tqu1qxsLxleZnJjD+Ldt5UtA89OJg4gi2iIPf1Jihy
kKOrmX+q5Q4cpQep5Ne3okGQvT64DfqRleWL200uDpEHJUy8Xenpuhp59pVXTi9Y1nS+XEsWuHiF
Z4VQNQx8MSw+a1alsxh4mMI9n25pT/6fH6huVRUX71VuTzpWxOUnz8g87VDbLZmrtXdkQL3ixxIT
lbBYfgBPyDkkv9t9C8iKPKy7KtsbwkhqfrDpiWAPNBlFHSCrWaKGR9Mhh7ItUd3L3yFLpomkxExM
BbaZDx6ahHwHRbM2RI3BSnW9LKc/ibJ1i7FnO1phSbrZVC7ORJK5Yqc9ynuzgIwgyivxSQR6szGd
hPzR8nDvwiDMWURj+9JPG7+FIX4nCFn78dLz3SL+pOBTBMzaCSZc+YkiOoRfalxGxxnuNyoj3e/k
dyhiQvZFonzIvWmaLOC3Miuyf6OP+psNFzaZ8nb3uYL+KELSa1IhDBcSOKMwBGWFtfTknyX4Q6ZT
A1cHQ+kcUKfAaL/Vkmv1DD4x6hCLHC0MIpiLxW0AkEJsAMIB9fuSf+2p4h2T9d3MRHdFvJi1NiQL
yUFad2IXQfWS1W51UdtI+C/1Uif6S7BH5btGtpEh7gaNhrxQ+StZxscFZvPRrQ5PPZogyTZjGpjD
5OLQ4LTxH5mRnAgzfjztgi3YqvUlR67ZzTy/va6/KGZ9SP5CkI9qXGeODULzLA4nVWX8bR8rDdv6
5za4UIn6UnfHyAqEhpY8En1ZHXnGkP6s4a3OubcB3HrR3k/01rMBiB05OPfKD10yaxf2DhikkvCe
OpgL6wFT9g4UzDc/8krOfnJ/oEFfuy//1JbeZIN0yi8mZkozLRykTmRK5IlChg8wlXGZCW8OTcZL
49iOH17u7Uff1Kv3zl3+53/CbfMymriGQxrYI2Tk+Z4mZyJAzetS7Sk05TIx8nb+fDs+Mpv00YnK
4DNRv/nsMNj7UY8Q9ovBcVhW64b/GKNLQJUptTHO6qHOsoh1ighqzzp33MZEybZoqpr3+TDrTc0u
vowhQb+Y+RX+5PQuwNWC1Edc7AiVqDE2zDw87nQPnT2iG74iFBhcTH6IWjje5JuDkMv6tiOTb+iD
IfDWYQIrmwd+BJxEuPrxkuW3dr4EQ3Gy4G56xb+WJMl+p0WgQXpD6gezNflK5+/iCv8vSum9LO1/
sZocgR7hCVrTM7XiFNZVOp4+MchEPEHnw9cysXv3W+8TvIL91tsgdIdE647wTy5HwJTw4+vbYitz
o3G4W9n16LmMy1NZUHgBtxpOrrY0Yh87YB02+mzOhxQfdS7pBYq3JQjFXyvYwW16/4K6mdY+kws5
ZsIEWXURpEn8EtpqVqOcCKF65BQA23T1i5TMggQkxkZeqCIkxAYXpUBfCAs99GsLf/XrfhYR7TdS
VTF4hqkj3f+5T3idwhJ4nxrziSKjHBpeq30KhgFfvl4jmM6CIdFuYuBALAMN4nGl8kZDo7dOtZh0
800WZXWVFZsv8RCAe7fOmDXgJVMhN0Xej7HJYKRJfRvwO/gQR6JmfcGtzSdSFDKSy9mPv1/rer4D
KcvmgO6oKUigckwlFcyOxfPy5/7RZDrSvQXWkFa2XYDu/kMo17XpI+vDenVIOyjD+UKSqX4qNnEa
r0aVSDds8Efs7lk1XtBZ4gtG1PIcCIusELeZmm9ixA1ORDv8dTkJgNdcrI13rAk4Awr+wJ+jyJg3
djprsc+jyXFWZtsman1+0nGS5vm2is2YjDjDg+PAGBDa2agtltA9BCW9ieLRh4/cb9+d9Ho7iqe2
+vD80F/5IcyylIKM9xOtoPVYXQUhfn183ByCQ/mr3ELuQHPnrgFSneXqMPLNJ5KiBbhGErPUrjEV
95NRTyU18mnCJmnfxKE1rlGgUtdKkJhPAxbKAW5UUALpquDWrKF8mrwze3uoT0HCTy3i1AfGSeL0
6bZEJqDNEJjVf1wTe8mZHcObOxNBP9RSAESn7hJZ9JqxpNb7pC+jXJ3+izsKwIENfEqdczK7FFqe
o1knYSMVBaNNjxY74jJY179gtvbp4eJdhb/WnyLw6fEJ9FWMhOzKk9te75eR51OKFYIUoA1X6yNJ
1CnpuSDVM4Pn4Q9+E6Datxl80k8zryLpF4cfi6jTS/m3/F3q24iiKbv1GLj1SDdCceWthgGgK9cW
2k8SCc4eI9EEozItv/h/m5KRmQKZ6JBZh+jmMVR8SHsbbcVFD5snopfYxEqJrXiUupwEGf+vcaIp
5kUrDpkOniZMrZxoGxArzcu0xfJu8Ywhxf6Nsi+OyPFt4gHct9jAG9GTp1RbcT+AHpY0rhxDV9tb
Oki8mC6EiMgk30CyCcpY7bdNuvhcc4MRh1YIG1fcJXjqpEJs6kzz8Ymxn14W9t667OUffDY/+meA
Y0zf9qaOckKfYiewMjx5l/P8PYpJEPdFuhxGPfYB5dwYqpp2GsNvJS1MZhuFmCz2nth2LRA4sCv1
eDsJp4GYJ5PqzeJBO0dKeZelldNwSaIhdhfl6cg8lirVlJdYfa1k7GCSYV0FahjlYa+BuudrDzN2
WHaQSC/Mzsx+XFAR5o0tGTn4zLTfgsPOtU/0Qxz5BLVR0vDjWL/u2cfe3uzHrNLTKmzoRQ04Ifbo
iGNaR2tp4IYSlGa1n/pbzfZYX9fq8GICvQfjieQ2/N6SXLjr23Kh/e9PZuqGSxdYMMhA80eH/oIT
W4soAE0xCSIPi9fijZBVk5unrQa+UGsbrxHenknR55CzdnhDktzu+PY5NDv6//D9jD7vM8F37dXn
jNfWRmUSXY/8mn0h1IuaJ+MxtkQ9fnJ/FKdQ6sNog925v/KDo7QmdSttfsd/B5jzMDyM/MS9wYO5
WGRBLsBXFezhCXYAHNl4QaxKElupdTaR16SZl9RsR6GLPW2oYcRVThamhIP8CLuzZBybfCMgW4uC
3y74KjSHksKAJtlNW/SZS6xXOjdbeph0/pGP5mmt0sYbnaCZuDXRZpApeTp37lff+kQ6QbR3u/Uc
iDcs/6zkAy0H1ccynJ3Futw6dJWrT1oV1TDJhKbQaP7MwzzHBW2DVPdUUqR2MGV5dmEbsVKmV78n
yNhKLl8pzWoOePgauaej5aexR1xO3TWjYoC8+srp4nCyGaHNHvfQTtGkj4hIoc0U6AUIf6kboWUn
kj2YoPssFgm/CxYc5CixKY0pDvpcqeV/nrebkXS/6iu/9sldZ9HRsS1tItSy75yNqy/mtA+SN016
YTcSwpRcZjFW7nlytdfQHM5r01DNoOC0EluI1Q+pTLR0OBWX4P2olkewYZ7/CtuQFvv/6i12Gf4q
OIXDk7MuQbFvyoGEhhpInEL5oif/2xA+fTP4P77XEgJ9A/ApLySi2RUqvp5I3f+9m5sUg0F8RyDp
5Sdh7PpB39ad9keEHVTY7QvtPmOKT1oteF9OHLVn3WZVNiwb4UZRBH+7GbdaOUnzdUA+Pg+ASfNr
ws8DtVoWTQ2sjKGFZF0QzCpp/dyUL62fHftJLHYbrHu0Acx9kVIMsRe0vaFFnPaETfxrn6ad29Sz
UnoXQ4q1tB+ymyIe/cLG+rpo9HqaEPTlSYWHhWyRBGaudW2RlrrEwn7kppCiTFvEKhMBTM41CfaW
OjJ6i+nL6kbwMx1VRn6v6QEhbX3VAK/ZH1FWDiboYuJRnpIRs85zE1MY0GpKaftcqxybPm1A6ts6
cvMfwCWRzpwskM/XH/IPt/wMGzlZNytw+tQaDoN/yxPbjSwG+mNQCT/Xsdw8/AP5fg6vpuNTP9Ak
DwfiQIDqIJOlDrK06BPDn8ejqI9YpEJtpigczaNobm/NYB+94YdlAbqejIm6Ee6U99jqv+12qAmu
3BVi+iyWCJ98NNuH7QfOVPSzVECo1/V1gXDAT181W3z4BUypR7WabnsbVd2EaCkpGWL23uap3UYr
1NmM/ByD2MJq99XRQhk2rAaUUTlNHVvx7usNnUXxmWamwBobVNZCE46Dr7jLduK6oL2Zp1znrYPo
kyLa9xG8LbFH/c+UsWO804Fvm1vhv3Q3sGZDwcIj3RHjE/v7yds2XRg6NdQ/eE4weps32lQFscut
UYRUZT7xDWPjfR3Tt2/xO199cNsTltN8BYlC4Yum4hCKxIc6NCfC0PunZF+3Lh8O40n6wKT526GA
so5AX3eCQUW/02mEB+WbVzuuhXYQmRD+rm0v+SyRStjyCp5pwEMuJgsU/d6Gtcrlv9d8UFMnDFkX
k1t0K7p51K2uJs2QijTF86yFPcYnHK2JZwUglGESB82jXRhmwKzwOf2tf2qhKaoqYe7qJevjYwS6
lLTgAtFaNZrAKUIpVYf/7hBxsKEdFp2FXId6BWYiEw4iZstw5DVKFaPz9jga1sj/uYoKHKo8l87I
SFEXjqSOdxFcF+eo6ATvYfZq1Sr/CDtq4Xb4mUcvfuQqk4jzOVHQvtJP2uw6DlvM16yPp73Hevcf
HMD0UpQbn7Tu8GGchCV3ZgIw9KQieZloStciHSjM35ac7fToToSfrl1u1XIxGSNRISyqRhCZC7iR
ATwwtdHZ7TOAtbktEeLjofvDMyxpG0bv2R5gn3wFYj0CZKj39oZcmTGPBGbMsea16YP2JxI2iIPx
lZ4rD7mivi8Oy1KsN+h2sGNBHVQTvTMdbgkbeS/XkIkkrK7Fu1aMwYHhQKcdrWyM6S/ZnAZQ4jM6
13ZHQmHJQFUscCopvh4gmtpiUGrcazhzQj6l3LL4IeOdkCIyN6N+4EN27if3RxuPoI249nTjsD8f
N0hbhay8EbXOpf2outYgUGNlkIhiuf3HF1BsDpkqLoPsvjsvUzHLi/ZuzAU4TYmqJbGFVEJ1ZWZ4
fMO37qyVryvBMkkz8/bIJ2ZBuzN5EXr1biGR26J6M7pUOrcT8lVcKuug8ymVHVsh5VcziL8otq1N
BA5UkeIwBnB6U59+5SJ9SlEortif1W6cuP7FKD+QJGilobLwiVd3ETP4mp0g61XZdA9/zVr7vIEI
w4wSV6USrSfvQmsvfxzQMvbsBdXHqGXNP9JQRHVBlTIpbxHXgaeXLxzelow23R4bgj5W6oWxJKJl
51fLmlO/kbeaqSWqUD93/vmy8CA4DdXoZZ1ue8Jm/YkNH5mZ0e9ARZdX1KpjQue0aaF2YwZbENPc
Hmjeu2iyiolhCVONeQ+IxSCqRi6A5eNX8KSXGzUMW+E9tTrgM/czpW+OyTzthhU5F5CAqvouxu+v
p+A1QeIZPxvbjRc57p0OkcVZpFDpssPT25+pwRaeDFT3gPml3qIX9QCgGx50XlwGpa+SS8f9pgZq
GOEUF2vjQ7OLubCckDWN8U8Vbxz44ZVxUA8Fs8hApJ+5EVkBpaFo9CHzXucDXPZgBsEfH7jL6K3+
d1+pAplhXj0k7sJ3yx5xxi22nGvAjoedK8A/bo/fwdM13/CMEkNNWFiZZeAUtFCq3iHmEr9Ut1TV
TGwMBgKGaVUIRAQu35roCpH9xvxF7DbeZYNQnW0DeGhKMRbv51sHy0/VFIpSE/wTcD7HpMMS5iL2
NKnpXtDCu6E/EyE2FFQ8vtvj9wFo2isi8qkP+ns9FE2In1jLtU3QgIdfmhtcpIxVEUqVRaOw2ojC
wj73nPM/G4Z0zZ24Dmqtp8q7FIgaK3p6mB03YC1VRTqZA+Gh3v7QtJIWp9LSX+89MlV/72cCTQKN
/kO1+x9QkKiWb0xhoX7L6JQ7qWASzFzr+QVH6/40j8WzBot8aps9fy69OEu+oM4hV54UQ7B78b5n
ca1h3KV9VtKwmYApBLG9nOxb6u36vGCjTJDVRoiey/HbFw14JlRUQn8dkahd3gh3QJQihsBhg2Cn
CeNDONYyCWUIifaxdNTDbyTazTIzNu0Rs8ClPzk++8r2kKBxWE3/ZAZBUfedlfHRsPSxMJuYlrMz
yBHIw0Y38OjOjh+2OuiMmx8bKy5zWClj9/gVSyEld7Z8QEbTQGYIvNcKs6CRdELfFrwk6V+ud5AO
RxZjbdhM6aMwiXM0YftFR3XFRpo9wK0WLA6s96PIV3WtxCLlMrbTAKuSfynTNenLkQX69P0ApDYD
hCDznJhBmF8oO9aB/i5U4xmSjOr6USnt5cAVA/5y3aTljKSB24PmoB18IPkByhWoAkTiOtd80BB8
eqXH0vKn47iDTdhgesNFLieX58nqJD711wveiroSVsQos8jKlsm9ASfsXHX9Ctrwqrbrc3B1tuyx
BuybfPDs9Xy0cI769DbZHfHQbdiHORDKPF6uEw2QZvUHAlpzt9HbqEG/mExyp0APhc6HhevvQIQB
Au1+JGaeVmKBm3o+dtoLdOUApiZkUFanC9iU1LkVZMG0amtc37tKWTNvoT7k51SVzrom9v00fDyd
PWzAUjkaUn9rKaIRsVJMtdDf95ipfae7e2Xwopw/QObOPet1SQ4U7TXdRa+rR/wbrPaJLMAMZBgj
73l+RM3BFw7saGMoeZcqjziMKMnKDPuUVBkBQPv03iXNuXGkioJ8wDKAHlYlgJIci8miu/zI1twQ
B6XCwBEDwmIRSlokr3a9MzFo5KW7n+FYV5650uo7v5yRwP+Lc9MOTx2QEJxBOOSxVs176T8WccLu
EqaEMuajOnh2IsG41zBttGIBeqhOVFxERQJXvA2Wv/b4UfPR5Cj7oZ3Okae9k2KZ89pLtFI3l6nr
BgT1MICiXLdyh90M2WygP1r4vXk44Ek8q5/vQRQSJFA2UPJEb0NrjaZmyi+UNcYJVog/2aTjX7cR
BLUdJgaS/fFGZjmwHb5+QJe/4TIf/68M7xlgtHBKHIrD8yrAL7+a5rf2YGDhGRd2X+UO7kTVUjvD
zs7Ji6jXui8nAWDXd45rcqAZ+vPCepYS6RGfLBuWmL3t6eq+GuBDi/nwO6fYQ/DEvtR/GhR8fGRs
HPRZqWZgrwEqW3fUhYVcsw3E8K0tlrXc++8I2HD2/BfR0CBa2vRZYDa8zKzDHNzceM1OrP3vIgok
uEKR48VHlC/p+0vJGFNXF6VGH5mX4QL5UTB5ExsPYNnoTz9LXhAPzWTUCPQkS9qjYQfFyohQJZaB
ifMUaq2j62NMHqF1exL4GIofjrJ1XT+dWrva18j0Xf0fwYV71iuzYVDasndpOpEXob5G7G+A5iqO
DM3sX5PvJMFbRZsQGzKVBLvR78izg17BrrSulfJanUjqEpygYX+2XuVcl6QsLv/v+g+n/eGSlars
QhG8cZ83J5xC3V9sDryw3BeN0h3aiK2b0ueTA1ftmwczESLluE9paUyMRq9ZgEOICsWVWxYopno5
HEQ/jGk8Yk7uZ193K7RXQpbJ8crhmDvQLGZOv3+u91Wo8e7bCvEn9OULV63haY+Y1YlZgLrmFhpo
mAyi45Ledziu9dvEgTGq2PQqXvGIedK5rpYiQrP95aKHbrTzrkHv3IgFEcKaZX7phUaqIZz3ik3a
J9Xj3RAsA6ZE5WDEMyRoDeO4siOVMusjC9su9K9GJsEMTEw1V5FiwbbDxSRiVyUHe9OOFT3yLd0x
hTgdutH0IJL1yzMALnvenBjhmDQxiBGMU3KtRns9S67PFvTvWhiOJNlrRn4FiPP+nNgnGzbO8BBk
IJXYSN5hjiyJ0aJi/T6EX77hBk1bXnojIYNOC0j0sqjHjWZvHukhMkQogmerOqMPQ+0uxHaH/+NU
Qt1S2fRnLcFs6GIQujihyT7kNbVcbOBw1fM/DMCsApndabMBGDJiKBqHzBu1evUJfMNgu7S/5TLz
t2eVSk8zzLh9CYVA4ImTKr6ECauf9QpYXIEZqIx8AMqu5xWUYPCTagXOHQbyzwJnESdXOkjOgtEY
xmhf6/FRNR9g51KbA/OCV0WUEShTLK3HeOxp8BVdSXq8aPXOFKgdsqBp+7haUaBnjPEGBK2Gf0Xe
8ETrFY0l62eegVG+rEZ5KUutyO4d3/IiU2aIEK+koopC2Y9rXAIpsOAdVzRHC9uSaH/KBxmwNN6X
P6dEz+3jXVr953QRiTg93Huv/jv3XSlInLQhKaA99Ch0S6MIkH17pYGChQRnPrnOqBInWJDVtbAY
3C4QVZbYf8lIKvfjczDvcyDRQreZN8GgxDRnd72b2F8ilIYIMiMILq9Z4tRXwvY2hTvhNaqMg0jD
TdtHxfVmU94OXY2kTmtp5S8rlqG30EN209GOGeRBiZsgmyC52wLd2wT3zQa71e8KBoLhdkqT34PO
PVraaqYcCnaTCUxmd8RKYAsQl1CR6O4D0a0w3d9ofdYwUlLl5JU4NYLTvF0QgTeB2W6XDwIQTXU1
/f2fxODRpkoi69guUS857JIH3jICoqYATdw4SKaeaM8oSiGeImnAy6x+kLJAjarJ0VL8N2bDIlnT
WsgfrqVNOogP/JPDUtzBH7A2Z6OY9Mu2l06kqg6RlyJsYLrUJxkVucxG59n84LLfLmK4bz5WQsKp
g1PG17KySxwbnI/MdKyDqD+awt8AzjJjG6irpoShtAopoaRVigO9R4piIPonDlzPvW0V20fDT3bc
OsG1BaHb4ekm35yDyL+7Kie2rSVOaSg36sNpZWymlDR6p2OOkS3S0Uel+WqiuQeu6a1nPPCv4dL7
xxrGthJe9m2Kv2082u0mHXKDmRKF/q+4yTSRl3p20MPgqdnKLPpgTr2a1ThsCY19OgC2NnE+Ysbl
8jJv1W+B1R0At8MXOaRXflq2V494etVSyU0kgiweZ8TFMmsFiETby4nyypmzbYMqXtIxIO2s2yAV
WtafTIBImiI2QH5QZbqKAJnC7q56AB9oTWzzhPnOF4UHJk4UuFDryBXPgNPF5IIT9rdUXJjoplBV
7NaEUfRHbDFzqadoVy2DtQK2zgbHbRBhliRxnB+si1eVms2wzgDol3rVIPQIcl7Mxlbyux08Q7oj
es5Stp3eiv6N3AG6o1WgESApQH9NW12+tFhT6+16p34DQXdcfcORcUJZjqRGeX3zZRu4O4w99uIo
1KVGZfAZHWANXnQ/Rvy1pmz+IWSnY27o4bi5cK2Oc0LemfYpei7UkSe3lLX6kCafkw/wAvtDBpa/
GE8AUIRyNfmDvlgXuF9O9+FHEVxwODHFZY2tU1bM9/UG+YoyJfOHbbz4M7cxF5+TnDGrmVd0yBQ3
1YPQ/C7ZST9B/QkE0hjkEceTYokmYzTlR0sUPz0JqGTeMsR04CXdiB594NaD49JMiYV/Gq/SrspH
DxJXlnLAdfW/isdxGI35RvXKn91IUUS+HCtkSCXPrKTVm5NifXVew9N2+ZRA13iKh7I9/fgTtQ4x
EwLsgPcyWiTtQJ8QxyselWcqgspT/VP5HC94WgadL6bWk8hhutApMXE6JwYWdXzJ5ZMGWxklF8YH
j7ftj2sHm3+7iZLQIUZjZBE6XN7KsD5vaGKzr9OT94IcNFF+Ez+sLhOJBFuMrP0FyzFptPP5iPyP
O+A1EW3atjvGloFK3/+E2bu5/elrYD9Fj8DzzMcZOBLMcq6rRcxMi/aRPCd1L/Ac4QtPOcZIg3jw
fmtznX15FaVsFu5IhD5BQT6Dc31etK4Hqu8hi2t4b9PJQTIC45v7ycO8CAulDrMAf1XOlhauVdP0
NdKhTMAylmd8C5/oqyp9OJ8+pu7yZMJuyMZMeohlDfP2qn9s+7HMPPKqlgeD88+tuNHooUb8e5EB
xYjXrVqM6w2H4DNRHDAr7ubV7ypWBRjqrsQN/U3JHNg54O4P8E8GtlRt3yMZuCkQi2IYRq/WDe0y
M5DxDgsFUrxpU7qMIjanvyadSt++Fn6iea8NTRdp+/Q7uKIcKQrsvszI/t4qtk29TBspYYL/VG7U
D1UxLbSS/2zlhJl9mgQOaKYx7Xiy1LE8pvBKaOC4PFn7IKQVyx86t4GTlClo2+gSgmpTb4uPqwDu
bCIBqwpEnRmG7F1cLYn8MyJcSy0FaZZJccYXEnrvcc9ookPcjRMoYb1qI0A/kGMuxBKKdOsUXcUe
gVK/d59xKg+CxyRWrxpSmau84lrbHZaK4vvwuJ3/dg6itUy14JjJx3n0mmWrCnWci+fgNiMD0TBb
A51TbszkxPXIk+3wQnwTOtISylcGwpN8InvP7VOOS9UES6oF5Y54cT+iWy1PSb6LfiEV+sh6wyEg
9CjYOiwPJqPVKxJsRYipfZbMpuEcYuDc1TfMC40Mz+Ggf9Ean3uGAmbGYMVNHH8QKHTErAwdVWCn
DZj5jDLcqpSc58lIv9D0F67HbPaa4APKjfM+Td+JV7eRoH28LZQ3W/rhZb2Pu0DrftGnbgUPKWpc
8XIIUZOPswWRGATqgJrkVUwDWaxDP5e0xuHUAt6nbgEZ4evC5twKH36IcYhxRTNDUwD5GMkNsypO
entsZqPbql7hppQJMwkCgeHqoPTXR3d5YX747tewXLfVJwdahxwYHKaXOh3mR0V/u4WGIVA6lEm4
Z2ZYQbrcFWSI9aN4ucNmSqshjYftg5162kPe4nLjmTKgfeT+p8TsqXTkQ4bC3r+VgOq3+qNrRk6D
Y8z9pozHpXjzmOeFUOTovk994OgezjOSgBUZVygF/FD1rU6kkffWotvVy7JwsVYwfcR9SQwD+is8
LjSYqJQA3mK9Dc17OW1pjw+l46zdjsskGj0gLM/EwMnvGS6GWXmqN12R2NHNSqyoExBLRwww33n7
R5Xus2YVhbJF3St7yy27Clt3qgvN0RHh/v+XcSWxVE0JUm4pNg2Zk3UVXM2cbAdTHPd0KH6XcDa4
3vahiwD/NE86TiHwLhN3xkzFeh2nIuusc2N4Dr9JU8+OZXnnbxDXbvT3rTS+E5w98JlADunCDfl+
uYc/2QxjFPWHQ+WFo12i9v5iGDFdcnRkIQYkCDIt6MdtgRZQiuNlft2OzbivY/049PyRCmht2KpM
EKwrjI838X1hfWqrzFIBTUEpfyYSScZfGngQalTZ3o+M8ZE/7NmFTOPseowOwqFzGat0PKsCBBmZ
dyv+8EBH2sB2E94vErwJa7ItB5buLi83JKWnIIkhPX4TgmcZ0Wqlu5tJH21KQFdWuumDenfKjwAa
411PKbj2SZG36Pqzs4vatMq/gAXamkJwJuFIU9A9PnPK6tOIBWiRLcM9yRQDrgMWFVKLttwH6gRh
t5b3ZKgnEuMSt4ReObl7+7aebdb70cu3T57zcruRfxnTbH0JXAd15vFeEfor9vXyFmMnZsoPDxqS
sLCSrjtmHb6+VWvuLs3yie3j5gOdPW6y+gRl1Mzkh4T0ZzfHkb4KC/AGIjVcUoebLFeuanihKVC1
35YM+USlpJ7EoWHj0ek5pP+JAgw+pKtj7pwCq20jxMpA/3bJy5d5bPhGIod2WwgvQtrAB/VBX5CB
acAAPnbUsLkfcuk2/g49Ss2ZcLaTS8RAUFWx87r0S1U7cZ/VcxVEkkD8Z52r0uZ8A0q/0aYhloUZ
99884Vjbj9QbI1fl3J4HDlh/1SO7i2kobSHe5pGIIFU4ERKYIhygXaWk9euiHCqkjyUTPBLFxmfS
sD4Ns0J/cLhqbnY0pQJNCA/D3Pai2CcYY93yoWRE+Hg99CIAExCQNEA/Gn7da84edJIQer+ZVQTx
k3xIqgIhi5CUp8jmbDxsfenpAZV77aqXjvWvfmnwkzeftld4rZc5cfUcceGpAJZhIsM/2Zm7fANs
NfWiXUKuPKtIzxt+bwfxhXku0Qra4s3mH6oGDKaUj4Yd7FE3wPL0hMe31PFTzzQQrLEWI43IZto3
jBHcKnM2IOSoAhSVwJ2K5lsdZ2ssR+AE2EWR7R/p644wI6WQgUsQsx1ybgwTwkwsFEBJnudy6HUF
yW2jso+5BqNokG6Eaxlu+ULIkK62YDnBGkBnNE/eXLepSUSgSKs6oxhhXS6b6T607ZcUJFj7HZZv
Qb8hyZ4gQ2y+TG63Ig/nSoaPKPRdKT8fv89ZF/IZu4naNRRjDmuzOlJDQj7vny22aQRQVSHvw7tW
6k6ADWarEkUj2O2mfiiZL5rdwp9SAvc7bRvUfERSz29oj2MsPLNYDnnZu/WR5fzSm3iooONL9lkz
+p9s0UKshaGZ1v4GHUCPPzYr30dsgbuiUFLbXus2fwhHsmNcg2ZxOTx/y968yny0ydZKYPakpi1J
0bRwJ4hSQ0S+1V+FrVy7sLcC76EM4fQIBJ2mGbmN+yVR4/jj7/xkqQZ+2WEA+snaWSXJ20z9AL7O
AXzpfO9VGy5iI3aw5+tvx14pfAebQsB3Vc8dJaNUyG/lWbn14HXi2SGEZKJNTR40zJxCN42YE4Iv
rSxldsZMW1GGgxb9iw2+Ox/vLrwNpX/ntDQDmzkAtG45fw4YsO8GeILmcPI8RxHk7wlXQOGP/Ov2
Ptzksx7xg4bpxWz2IZlFc8oTbfv8Q4+Om7X7yQMiO48XPR9V+FDVoUGCJE43p+x55egdaDIy/5Ig
JKFvQUt/JeKR+E6lWocfgcSCGig0b8vO8pHMewbbL6ai9tmDvCR3z6hOqqnkPgjD5OzCu8dDtRcm
c/qubg1m9oQEphDvTL3KnYU0Dt4pK99rz2lLznXRi211Pok8EiIPc/B5g8PbKVPICVtrB48C/giB
MVEFiB2GjwEer0hHqIHI2Dp/p2wNCMjThHOHhoBtixyRVlHFilpOr4QDNWhWCcG9cCl36MhRkD9S
PyKGkeQAERZjJv0pwvUAb00ArUm+sMtlRe4h8uhXBFt0hhLYzjuVRFLienjvxgMKwXgmMGz7NmNR
GLLn26QlS19yuVO1QgnVLs12naMSiY548astCl5W9/qR110nZ6FWHYqw/b02z2/thRbwOuTs+NVR
It7YX0PpsZjLXxYwSAFiLLg2hTwKfKEjwL6aHb+o88MgkTxuUsLlhMDI0GpVC2+AcPj0Yu7UZWQV
SWk5CEm+AUQtjEuhd3ur770JhUyuW/oDgimlbh7/AhyFH+0Hr+MG1QM7IujiRtmFFbH5K0KQWLJP
45KZzqmuABcs6oFkFnI/PbwvoG71TBdybAHVRmneBfaNBY5C/Qa02N7XqI5I1INslpIxYV9j6vOs
rNcegMWJRDIh6JY7aIsA4XGc7NRKuU0uLx2CCcGuhtlu2gkmv3GyaMTiCPagPTTOYR6z7dXLz4jV
im5pgVt/HF3HXPJFzHVjNNcd6XzOf1XzEkU/mrOrhQzc2wVcsSSCFqoJKDj5nhG9kwe7OCogKWoM
DpCxukuuKCGKvn6gMD8Qx5vLXPaO/knTfQm12lI3L25YKURZWqRVLN/pzxefJ+2NBukOp6f3Y3wB
QYcLvfbhAeqnEZc/9iLlHAm3sMMq11jrEZ5jow8vKTPkgEXUl1+W5DqVfABeOlGoUEjlWtC53xH5
nTqKjOI4jXof0XHUjg3pJvNhSvipgI8pW3T2t+EFp6l64fNASKWVZjPAR1C2eRuIxQOpscXY5QQv
PKHivFoCQS7Vxj8dK66vAO9ZYooEXfiTuzSNnYqlKo/NfzWLAYMXbI2b7/4mGqj3J4YeSaQvqgrt
bOzqn93kp6P6A+qhfXMOwR/7TVn0bTdXV9VM2P8CZU3nF6/2w5DaIw5HKMM/7fBbZPAMEHYbThW2
Efy7iDoG9RJwD9rLQ1/bGpIHJCULQ3dodOYIEVKVqG7kal4QeVDOrmw82AeCLxzLyNEZXDpdSKFj
Vs3OalXXFkZQq/lj1IAk5iZ1PXN/8Ek2CYOpasLOS0j/LWbjG2ju3vpJ/JdLQS4xuArX9+sn/Gib
TaauhkCTNk0owiLoiu2j3FeoLKOvu9yEqHtS9s2I5dHN4rE6oVTcAiCSgRiNLtN7YguXt1817hdh
BDIYlc5E6rEpSSgzlm+LQ6+EZMZgh9qfujUrMtuQc474e3ujUfcZKnYJ5NQS8LyWFmp3E5vIgAVN
vAm3mhJiNRO4H4KGwysNOi8rmqzxsT9ay0OSztpLye/ywkpbzSflAb5lXxr/tBrW3sd9O4xsyVMZ
YHabw0+VlVk3UW5vx2vxNJ225JWg5i9FoTJZy34iXhtswz1ntC8McLyNbGQ07VSFWGCi6rYVz4XK
FZwQSTXO5xmFVQkGP1TBxNEcCb+XC+aITLA9ewtwWtws1h+8WC+g8/fdzMowKmIBpp2HZe7orePR
FhM/AYSCbUZjjdpUSoXTvPhbRdKHAphCjIJQkV3ZffSSdhyw03nfw6Muo+msCbLUn0DJ/FUE1M8l
pAsDz5LeAsZ8DtlweGHBE4o7EB+MWznEklQdGt5zqsf5pJZ7cxNzZAUZYDQVvS6uQxxIHy1kB39a
h+m0tiQTagubYVki05SwV2ALBXR3P/XHf2ONXF+yIISn0rBQKIzoCmj8m1COl+rBqCjSgsqic0TC
k9KWmNpc/EFOVWSyMdxvhNijg+oYcJmhiOBIO5VZWSt+MCozfPng2n9dGXGQdEu4gZr4sU5WeVpY
2IMHleh1nWSKvf/dPwB4eDjeuD3EvIBq4oR6w9aDudAwVRjxTqQCbgntfRfOHAvFyAAaTNKZSDhx
8E7gLqQTIM9lRxBNQ0Nyv0aiXZW+VVQe4G1qD9N0b8u2t/g81ZMgKlSZTbbu08/lItUWpf7yT9g8
BYDK0BU5u5du3IIz+Q+SkjtVss6bA4GJDGLwHHpp3fqsQZrF9ennNdyGZtHxmUkZGbVUbQMTOZK/
oB1YzCWAS1eJ3Mkhqj8dvhRmOZqecIPd4DQHzOoFsd3vb5be8qcbMI1G66EMoWsN7WKtx8PSWq5n
uvqFH0XN48N0T4gh+bWIR4rf271lOcpHX+CJTpbQKXCRx3PZ9CkX4Q3LHESDxdJa77hjDNMzujps
8846+SYuJhdv/tcsh+JrltDjEFAHBYkKfhoV0BpMIjt6HkLyun1r/SasTwQXKOjB6oJm/CzKi++9
z60ugluTu1FNcctkkP3IqjyqxVqyluPcnxPKe+FLBz6E5wZii14G2hAnw1LYtNsS5+AFF4n+wb/g
zK3bBk8NoWTQKccJSc4CScjQUmydZEwu/PXAHxJpwXq9oERABz4RTbo6Fek62Lw2geqN9i+AOASE
McRPFBWFXYR8SYhAhLru4wcjSxQmaBJKXB46PugNNIfgw2d+8cHq9IIhco+WSmY/aNLmULTZNP4M
NTWcC2RhbqRW4+vQ235Vf3RARN2v4Yz02qB94+WoQH0BjODnHlgWfD5sXk6sf9+ZPfuJnO/Ar4aB
UEqJ2bQuuwfQiVhvXV3sKJUR2L4oAGfJa2r2bVppL2VBpezDeS1kXuCp1r9rcyudbcoR7HDCxSo9
BpOh+N21phKPKldRUiHFlDB3QYebwXNZHzhRME554bELsPQeQwupaLLMbsl/yHZ4IlfFX1v7gw1Q
mvCdnCVToCGhAnbVaECtVGWLoUTwrFyKiyjZ7c8w0k/4/6juv0vCdmib8IfTGG4dV0OML9iIgDrC
szhOgNUeGR4JuKDM+6h4pUAWPSnvdhvTJURBNy3N1zDLyFTgNgwvjgvogQMDqB8x8tJpZsgimsfD
+usRZRgjhEYL2FNwIUpvDmO8KjUfI/iAlLsJjAZgylO6TT2T/lj8DHnsOiBJ+0NhGVqyBxwkFdVf
OdAMKhog/IyWMOaW9Nh33u+Bq2MbV3S2hgWi4/SdIKeDhraCb6nXG5r+DvYiY8RNck8JmmnNVKi5
AsVTvxkKeDaHOwh7rZ6cL7HQWZsAXBAds2NCOGceP3HS9Z+D8pxtiFbJ7nkT/htqvZ52tbp78C3I
0i/uttmxZdIiL7saBVYFJxOHNnP90T94m4I0ZD0ICCRP+J74KJmEF2Furn4OrIvIt48oAOKOVOOd
cRSND3hNvuQ8e4oG6XkXGu033sMfU92Lu0mrOUc3ChhUADeYRgDemfXLLUiTDdYeZ82fk6rNYl+f
UqrJaPbzYxunt8kguyIyJ7Ywkx5FzqFS40qXH1sKHJBd0SzcC1XnB5/lYg5WvL2/P9s/h9r88CVf
E9EqOo7rZwvzx9RNJWQ3mZbmkBrujw1ye2/d9wHSZ+vxSZuZgnB9yUrAnHrj5u4eiL9b3cKcpP7B
Z9FYB+IqSmrVr9ehQmUs3vRNpQjZg4H3t7K8jkytpYx0U5eAtGylfnJjgrXfHABitLX1nRwVxi7C
23uQ8+SBlEtv2fjeT9qid8WOi7Zd7bSjHgEqe6Xp9pTOhyMyn1Z1kcLgtCq1DLq9Xi7ENY1GjxBl
Sc95wZLMSBRiCEAaVcKUyEMY/ZXYGXH9xt7eIdnYsd9jKBTaJxcRRhlgZw3eh68cafHmRZblv8N0
35X1JMKpgXOLOTiI5uvup/dtYhXMa3AOP/qmEQ86vuPCFvtPB7AlQo+U95/FLs4vC5Uy5C0MG2bx
wGg9ADpF0qPHTTUgjVJV/zic0/uFk2BkdElPAsriUS0qeGmROuAq9Aad6KNSv72KbPKCTo03ru1n
42nYDSJEcP7UOXijIOLrxKCkob+EkCt6AJwK2Q72Zgo/S4F0oFiPWJdfMPWEadkTOZPdCVWOjtJX
n183qC9f0zaiRDtgrYf5/L3WZhZ9QjkMJn2/FO2HT/XJ+9BzOoeJyz2hK6NNhYhozK2rqPXQ7xub
E09YbCgn+ahgGMkdyA6wT5MPsyRCIjky9FFmj0Ogw9BnjCRhGuOtpJCQf0h5gHGqhU8sleJ66nNC
aIUxxfHV2nXqwePwP3mqEWqIJzjK/XJVbSapMfNGoGz8yySw0J7rbvCoiFAlNt/rccOETTSfUj8G
qk76PDntFm4pXPKmeFILG5z8683g2WZf64WP+iJMgujxq4Qp/v9+b2R8BuVnIXj4B4Cwtv0wTmPZ
mMG8JOlYI/SkyssqWSpXHfyPYxi/xqRVGCgaOfQqEiL6qlg1kTuJELFd/RaE9wlSZ8ni/Xl0EIyA
qbIgD8q/br0XABgQ5fdcXBVJYbNdtY/MAoDVy/3KCanly/BvqjbhBduaOF75plUt9m0AQvoD24Ld
q84vGVydQF9ofqyAcHdSrty73W7zKQAaxN/BeL3g/EnQNMqOyjp1Jji1fy7IBCur2b5iV//934b7
9DquXSEfMYtpxOjINSb1kMKn+TddHCQcUOHzk2QEM85WHHTkt+WyTuic10yAWT7myy0mweeza3pA
4yR16Z6AEvkVeytZY1md8Xjxif3FcrU79uxQDVV0nU8E8d5jBP2wqRmuC09mj7qeRa0g28oHQ1ip
szaTpfLkVa5/5IJccJ0wvyPq2qY9ZlQd/Zy90W8lT4G5w420MJbJgclNXnWGmcN3CMm0hlFArN12
7yGppLajQ49y5oX81ui3qLYj/gCpQtsm3gZ/P5Tle4dyCNSByLeGz2XSHdQJEN6b7iaL/SVExazp
VqjYGl4lCYq2YZorvYhYI0h9OA/28JqPJD5DnhPFdBre0R1kdk2o8KrrZ9AVbmQRyDa3W45/YyZu
7Zz1ybD6mOhaU1nLh0aTFE0z2S2RB3LmeEjEYz2TRJaX3A2IeMGW4xV1P38RjYV1a1pRQ1EnbMiv
2soPgtP+gPyQTRwRCtqn1nmtNOLB1aLjZ/ibpYl7jx3mJnGy0Nc+tJvXPf0okIbrk5k9IC6/x+rT
TeOdWSaSqTz14p2aHLw8I6MtbhypV8i2DVlLybBD/qmFUqSpVmI4+kjCW3loUO3NaBB55C5SBIha
a07BA6/neVxcJwSEThfBUKk2XuhAW9DyH4lURYuLu2e8ROk7jkFu6FWoeATdYT079GfFqygv9dSd
NTFmbgvPp+5ZwFIOWWcxcuZmqcRslki9NGCfrLslmT4JeHNepw1kzMvaCjOqG+Cq5QC41e8u12yD
lbDg5vQJv87VHxVM7bCSg4WF7cjJjjXBRwYsb0UHZOcDN5aHI4qDUbQnwICCC9qu88Ydc55TZ9Ji
BKrZ6vHcjWPC9sHnIxchq6/MfKZdXhEn2KAItBJKK3YgO28MiGPgqA8cE03xwMf4FLml7gHhDSUY
M08AMNfZrJSs6+MBhykOqZiR/Xws5IhGnsRT2o4sMHI8zz5xf1pl+3sMdKjhcTvLDPC0o7RCebMg
h84t8rVYFJoGIcQ1zYvT9KYRsv0lXPnve3vsCi6wwGMltBbKQ3dORwdtAU3ObPhgCXEOR1y42HrB
VFmLugLQJ22V5ns0qku5Xr5lGjAborzolSRl1nlPD7BB28n9t77CHzIhNkDoY1xCLuaTPYWRRe2y
N8gj9GeV0Q0fVgoyS0OcUa4lh22YUMP/HuO9CdAW71InFdVrifJoZu3E2p/Knxfvu2w3zQOZ4VKN
oTHUoCVROv2LRxdSsMmblt7qKNQrEKtmZdfdoHazLJVyce3wjOwoPnRHsP5flP18DmC0pVaYmzgn
RkoROfxQeZNe3bK4AoxW2z2Sjxgk6JkDuWreECH3r5sGob6szVu04W8xNMp3hy4LkUioy9o2iLN8
gDG7BnVQ9mXgsfBBHoyDlzER8PpxxoaaT41IDEC8m0GTA78FlX0rmh/3KrSv8CvYGRFfSABNskLo
eJFd6cCzjxDTdisnd98UY0Gjt74X+MyCfe54IDVujd8tWe1nYHerIqAgnq1bRqdxwjJoLZotR8Hp
IxP4BoTdc/dh+EaVNrc+p4lrqNQkJZG5/iYX06NqUMvzlm+fEEEpZiVNoFOfEYQH9W2wZjJ1ICbe
F9HOfkeOG6Pwp+OuLc3xcIjbnTBtyDddecl8LO/tCbtar/YgaSz8qeM8trDZJr387CSC5ND13+n1
dpFy7F1MWK0AW8HHBDRK1IiyDUz0520zqhgcgQ6gN2fE5sS9uEc6GRaNnVxOOg5V1qWdSttJUnLv
VkRPx70WwFrCNLhgmjvsGU3gcCODhp/7dslrQREyrmXB4VUmL/20crvhdHUCXxnQKWSF5lry5xXG
r+sD6XgWEVXkOJ4qSVW/jx5+V2Q/cLf8J54w6k9UtScj9lctOr0nL9NI8QMxTy3YetkA/bocLq9n
46NJc5BfN6gnhiuP77hxURIj2aw5frpQa+HZHejoQyuwkg/lqdsjBjnvVli4qJpnfaHa+S1/athC
qfL3lEx+ZsKV1L4gU73jGO58I0+k9UzJSs7DdJaQozNTjfNfIW/+PFTXai3DlsY3ZheeTiL/QHYY
GTy5TQkicLSDi+gia4P8xnNuZ1pD6YaAarm9Q660tSRmb7Ptwdxr9gqDD0UeDh0MNtnLCw/lSO6P
6lA5cc0ywcJxM8kGFj4vhaV9mO4F05Ay3kEXsvSusd57t1q3yXKcC7VnsrKmdmwMi8VB4bwwKilL
4f6z1baYiDZczIGC+DgWITS8kIjIbLsPS/eWV/S+SsFWLNvPo+0ewWINFYq1PWMgfyFKpvMZU5Ae
1TOAGh1TqNkuzEu/+Lh/1mwdHeKVJunaIaYnb0zCPZXutKRp+RNpEYRuJ3IFHoUo7Mc9UTCRsBWU
ShPDiD+2qj/3FFjphB3KXNulWDuVvLgqyHz7dmRHeTuXMn5TklIYdo/MD7Ha89jRbFhZgMA/WS8U
Q8sWnYHzmjkj8EufXnLJHrli3WwRRGpL1dM30nuxKuD+uLKZxfIc3+Eot/rIHt3koQ3yGgOztR9h
R0wkIjPDhIUWq/AOSxPJSZUdSy5Q0fX6WlgQPzwcvdVbokNF1EsbqYcWJ/NEe+Ub7tVkyOjeJZEL
Ukyq96aVEuoPeuKCHFHRt5F6DK2zVZBYvvymB2GDf9ZN2jRG00NjHAhnN+coMueDQ/ZYi2uVozEL
XaRjotnBsB/SIBr7EB1cDfSMhACo/GEaoWRWho5I3boxmSGemS29F2lrr+ak16mmNhrGTy0cDCUF
J2D0nkPyg8PtEN4Q/ryyy3sVuglUcvXRfYIt1AT7yYPGMgpTRSAEktPOahChflwbSPoNg7QQcWPx
rAtcaK23v0eryKOv/rF3IsVv3UlNBQwDYROCjqrnc31G8T/vF5e1720MdEik2/rk+RLSRHIuH892
6G0WYwdYgSqX8K9HeQFkLXkhgExUnlqwySdG7tZHpgcRg4yH97ybXEN2cb+9rRzp8mb3q6aHvigA
EaEy1wCvW13+axIEnFNfJOuuBJWcDkS+Qm/4C8AIdbw6KQ04tjCYm7gGfsB34GSC8GNEUAjCKA7Z
B9VVYz76HqEjd9EpAl6Kb5rgPDhvQaATjiowFIgCa4rjPFzpvqHJz7ihQ713WThQTnNB8fIN/Shu
lIAanw9JQxANfBxywR+Ej0hadn0HCVcEP47GUzOvHCCBT3aHLLRgfPWIdnR/Y6i48//93V0ArENZ
FJIyIMLM2LbOPV6uE0w3YqZlyS/Mh0/iJhSLQsAOjHRAT1Yt+8mBPqfLUtQgC/6rkev8hit70i15
XJmG5v/2HSBaDIO/CffbIFC4C2xyOlhyFxbzxZ1f4Nm+O/wsVy5AVoTkX8GIf4Uk1DMDqMZhepnK
YPTmTDDwGgnkn2tKFZ8Qmt2QgIrlOLMj3uSgGNt3j+e1qrCtXDHKdfrJLsN63EkkEjedGBeCv/tS
b2/AEeKDaJqoKSQFNSjweZPFOPFRqGHGXBcX+3BHYPt3dS9OKwwvA5C8jujFn89BOO68Bx0yWZFp
diZiSXTnJaJFweuJpWbszrrWKkgu404BXOBabq8kislPuTCrElhHx4HpViYRuuayzWg9V69FPKsQ
lVJENvnyfxE3H+hRRyKW9akRVB5T2HUEM8Sex3YQUuTl9InGGQFtw+wleyA4lMxKl0b8KYM6+vlv
5DZZe3oT/5MsE7UJZ2eQowmAH5eR8t0fW15xn1TZhb+VYyb6rBfECA9qwhXFHgdN6qpnMZAvPx+m
WODJtnAUmb3/WckvBQIuDxkiOnsu3KhLaKrSW4I+H9NbzIcwhajurUiRXKAoGph8OkVotFdGNLMR
WY3HjBnmNv7iX7QDzPSZtk1bd4JOzmxwHjDElRZF9kNwJ0AyKTTK/sn6kv+yaN2Q/Ayv8evIMjcJ
eH3aKsF8KYy1MwUDUO2wtTBkDZDvu3nY+qi6Js3aB+Lmkb4aVm1/HO3prJwBzJd3NqMu4c4nkNpZ
Ke6qSUF8GRN/kEM48IT3mEF+wjQ6jQNzZW3uP1uca4bIdlCVmBBXy9o/G2Cum3nrlWL8sGVytpbf
jRejNK/XcUXj0XE9/Rkfjz+1REHxyaPnrRB1kSG2gAt9KgzPUyg3xkai4Sd+s9V0Y0xRbM9B3cyL
FUA2hfzevXLM4olWB9J8R4Kv/t6NKslXVYAEUrD73qcRUCk7dOGmLT2Vze7JKqdgBsR0369xpqYn
qGLc5srEFD9fg6YYPeb86/L45jGzdm+O8XDUfyE+XAOTYbQ5+2zqGFJQ4ZfZJ0i06+GdLMQeyC5E
1OehoDavImAKjg0SMpdfPXmi+EJVxu2z19pTIaiar5Da1uk5t2pf/RVkNzOvuzlBFRMHApASDDhd
Y/meZbfFrg6o0p7liJ9VoNErVGsiu87qRyMDfCln54jRyZGgAIld3+9x2YvhsjzAuvD6Q34c3TI2
avSR+5ckayRLAKna9TBXc18PWnYpHj4VslyHFBauYuw5uBZtA2n4cxMWGeMsppzdk9XtD8tsHqFX
0XqH66+CYrKo7Fo+q+YX1p55gXl7xfxouwznXmejO3f5F6jQn9hg/4JS51YvFOVu0amjVy4xdmjQ
iSE2H2BYwdw+SLvnlivvACtzk8Ja7q4MZm4pi34PoLedHsq+rznpFc3fGPfddSWCBKZ1cXf5DanH
F1s0Gazz7lNn9QopwBdWUNAg6Ef8YcnWUzfhFpjOuDGZ7BPo3EjbmL9oBACeKf9wRfALs4MzCdnT
FFMUMK+OAH+GVFX0SUhPhHQ1BdVmuSjUNN7w03gH9MYvm7gAMSaR30fDUnLkIk5kXhWAme9JKSZF
29Z7xrssgCNUtrfDvadhffQ3Ovcf/W/1tZWHlbfHH2FPmI14XvYOoJP/c1+g2wXkaeWy94x39cP+
Ibc2GJxspUycnPRIo3gjIET+J0PgwNOIShiSSBpc0tvE7feInEfg3vA9aEnak/nWs+12HJxGfOXI
U9YBIwBSbH+jPMfcUBiT21v5jxVM2lQ5jMsCRLiFJZDY7R6FkSeJllfZzXHwZulizSFYhIj975a2
oJWrlYlpHB77t3mbPFpOvefa9RiERlOAF2fASVIJlCAtEJ9NkFxKWWm9+CZDv9WIPy5cypQvidmS
fP+4noJIRVcaYcNv66Y2DeAkLG5H5Iz+cfhWaQZ7c7yk4Okp7dMgYbCd3hVJcLoiA8/3e/ZdAktd
9oo2o+kWYKYwZnsWxP4lYAdgA8b4Skq1TayVzaxsclZy5n0rmZ8EnDLxN86+nUKG6el1AfI5aPhK
i1pVIKRPYoRIP9mRFi81QMMFgnV+8HlulrpLBYezt8E7/++Fh8xI+v3dZ1t710I49PtCXdVIExZ7
wMk3SEhaWkQsnCwcW8KPqNnfKcKY0WWmXEeDlEPCnNFaOwaMu0e2JkZItKQMhlmj8AZeprv6KiyO
iZtLp2Ap5IFz5M+YfvenElo2eIl+8rpC8zoJvd04taS8kvwY2ApoTvx090xIVFlMS4+zLb0LoeiI
3RVsaXxipxIDXpWFJk0l6/LN1owDPpmtLtBILUsHaCfn+8F3DbGs9XoNnT/d2aKcsT91Ap4lOTEm
8xkSJRTqAKMeC273+2lhY1lu+AT4qQ7AbAO5opjpIxtMM8Cyr718PClnA3vq0P0pGWPxJZ1vT/gf
bHP6j2+spD8plM7iyNLsTa8ivcTCQmEziMeleg2G0LhnCOABy2lbbai7I2KTiapZucVOwM9OKiUq
pOfsdwoP0kv/uaf/bM0XT4tjl+SKSWDyaBo5VqwvsywPbvCvUrUvDSY7KZEwDCfZw6HVq+CmACrF
YyRLZUcR5kIAnu/2Twt2SMTFNT1/mSn1hm8zIQZGqZoOaooMMiYe2/vwC2mC833ktFy4JpvWxyke
/xUsPn25sVLJk9fIb2qL84VAjSdTj3NqYmmA10RJefXdv7yLE0MlX2NxBdoAhWdGWdOA5YpsqtWB
Dz4gVeuRld8+EcQrYtNFfj49IYaSl5k7p0y6zbDTOmXwcschQuRHaW9Sh6x7cm5qcWceIyzta7aP
dC2j6dKLGSK45LFpM15FwyxsDrW5OJal8sRjNWNGYD59vpFRskiDRmPKCChOu5aIOpqRaQ5PJ6ev
Gag9ZelEqTgGr5KGOV79qXW8VRIAUxJvKGk1lXMX9PAms7wSgkwm4b4jmK2osxosZFHuj/jLqZmE
7t/NCSRoTDMpv2hftlr+fybLMgq0wYMLgOHe619GACJGghrEIb2LKyRIfheZqtYSA5X9LEOBoM++
JZmEQli3sMkxJ0rEmR8Uk1YZkMtUktG+Lctor3TkmTACt/Uz6iMz+cw/ZJGrHON9wxvytH1uBOmw
aleYDgVDzxAEWu6rcm+VmNOdiTVLqBjsN+sxKTyzgIVHi91QZRFdEalpjDkHjhpILDQtpvRTsVsW
27l9TVakwZFWKnKq5eMk/fpChnKTx6Hv0EFIYpQT5yQjYwRd98zFAueSJR3SSdVf3HQUGFeVTMeJ
meO57AkQTkdiyH8drd81xTuoIdrIEZh8Lp6Hq2eetf+nZuLKEBfDGB9ws4UIrDr7ZYi3nkR3Lu6T
LmquKA2gVDbmrpicaOBlP+EQAeKy6FLmZAZMRz0mlYgAC/juiOoHlxDKZLKETeJ4ls5MydvE6nN5
dep5o2IdJ4MpZte2ARGW/fnSOkPicZcR4p1FyOmpgny9htbpLifjGliikpOU8ECLQhKH/VcX6TBu
L7mSc85cAjvh5SVDmlZOQW5PY5XtTFSHiaunuB61vocKrC5249Z4gGc++SHyQ27W4gMFDpP8hBmX
4XweBQeJWTmS3N2pCnIxON5G2Dk/3wQ+QU7xwl0zMUE5yka6wHMSg+0AUWec+e4wtfHKpsGf6CuW
`protect end_protected
