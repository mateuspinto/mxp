XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���B�a�'�kh�Gj����3��ƥ���)�C�\���m��E��$ے��I���>�L��T���hR#n���-36�oM�I*�z��'�-`��_������������LH~hCU=O�䜷J :ʼF�=�� �G�:��q}7|��h���ZC/Y3g��p�Kp��)TǍ��B������%�y��ك�J~��A�hCr�a�-��%�9��V��Ό�Dɏ4�Xx�� ��Y2��k���� j�T��BF0j�L��@p+������-����Afd> Qs�-����?���s~���[,�l��-��f�pa��� �FȣԢ6�K�˕��0�� ��Ғn.�t)� �{���jp/��Ƥ��+E[���آ�0�ʠS�<H2��̀'GJj�C��O������\�f�?��V��o�LpY�G���9={���Ig`eC?x�{*#�� ��=�μ�L�jJZID�ꓗ�q�]�%�X�WGe�K�xܮ�<���'��ގ���u�b�������-�c��@E�ױ^ד+"�l_4-���n%	�$7���u��/of�9��f����@J��t^����`�E�6��c!j#�/��!_;��zP�������'�=�!(N��F?��m���k���e�(/)�A��}ҲI.���!}��Ē:-G�rǉ�@��ɍ�����䷙k���nԆէ8�Vm ��,k�o ��|DU���w��X��ǿ���:!;�XlxVHYEB     400     1b0Ui��� � ��ǩVF��2P��^�a`>�e�%o��q<�ǜ�A��-�JB��_�7#�\�9��{�ʗg[�I��9���Z�	��;�N?���_5�q]#Y��ʱ���ҟ/��x@�s��`�^��7����w��� !�躍>��A_:�b�*�FI��˩!|�h��K8�����n�=��#MMY�.]�9�ge�����g&��M���c�s0	�Bϡ�X��Ɋ1����Bp\`�ӧ�a�����I�S`w ���!a� D=�;)3�4�a5#1Tm����/{{��mm!w�{]p�ea�`�lQ�T�3��Ij�Q�œ��3^,2=7�6��.63�l0xt�0��*��gV�ԐV��B�36rܲ.�@k�;�
M
��N���ĕt��\V?����Āb��Z���+:�
XlxVHYEB     400     170��1��n�O���OS;=���b����o��3�?8g�A�Tq�4��;:�)v�i�63��:�0��p(Q�Y��4En�VtE��p$�&��a�z��&g�;]�`����y�h��&���QȮ�wӴDӣ�4��Z�%l=(by�r���Gb)��I��4L	�����r=���$�8v��0�V��JEUG;*��_یm>hS����dE:6�0:��`�3v�%�V�A���%/��a��Ͽ����$���z�c�FUN^Ҏ��۠5ŹR��0�m+P(�α��#��ޕ+0_H�(�;�&��\h�Л����GT����]����`E����ؚ��������U4�,�>��rF����1XlxVHYEB     17b      f0��a�z��v�Jd3���I��^�n|���^��:��}{�Q9��yN[iK·=�ߤ��9�_���\�uhO��1�O�lB1t���rl��RxːG��%г$7����tO&�W}ӗ�FW'�z_�1jh����wV�����hv������,�k摣���ɲ��P^*��$>b�f{J� w��;��A4|ğN��ܣ�T�t}Z�1��3ЅD�t��*O�;[
�{vgV