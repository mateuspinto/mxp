`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4176)
`protect data_block
vSYC4Raz5tVCOzlXierf3CGDQ0oXdnfqZ+elj1EMoAsp/SXRik/wSMDHGuu7hEr7u1ggyWzw6++a
KF8QSyOvjcH/QgnoqIulki1SyLjaJz+qLN76o3Hnfw/fscZEUgW0gczj8K7JJ59AC+h98WjYFTC9
rQjpizrIhewTsr1OZmDbqGOUGCS4TWAE/49hDG9BW/WAx7MRIyF1Yxa8d7eoZFl7K+A5e1q1BzJn
Kto3brD/cU/DIF+7XmcdKJBdV/ROi0oVtu9oZzpymwGUFthgvE46mGG/1cZRczi7KTxyEZFdUa44
vXGHEgbVwNlxasNNNLSR+lBvOzSHdoGbzvyjvMgPXl44Nqyqqm3W/T3MLDGLAftGAvHqGehaz2Zu
wvKATEIRZQedBqf0w1tf+i9kkkw8XuzEWkLdRBw5ieS2KLJWJPUJu7US2EhmjsoYyeMMh5USdDsk
0lvLFAfMAvbWj9r5JQpbErJGJ9WcIOnNlgbRW0SHkIbCzEVH0yfxGxjU6SZyH3H40AD1/UOi2HfW
1KDq4A9PVb6L5UnksQSWFU8tcg9na0v/6mRe3U3WTAuDzKy5zGPg4xZABEJDxDaUaypY0G8HZxyV
dCabLDYtlQDxhvL4q3Wkgb6jkGqTYdsq7iuWOFWF5swW8SGBEu9lIQRryAFXsZQmFCPQWhscMN0l
luhXnXBCeHTXWlo+v6hI71nIedqWIyOk46NLBNbdTNBNxYTf5YINuzpGq3WSAMbmeBfhCzv0q27a
51Os6/Fm32e9tLLRHyberyJD5pBykfq/gfzMFP9XIpTamyjUJaoEjj0hp/JCPjAbmei5AdJVqkuP
zoWRr6LRXGCd+Qxdcw1u1+y9Uaq+jHNmbqRpVsq6ruRZQhynl/U6AuNET465tFNpaR6BjP+z6Fqi
2omvNuYIy61Bq0IHTnjQSwlqGGze8KzMxxTJEHk2EBEYXdjsBxk1nX+HwYzV6dE/sQNVz6Wqq835
K2IOBCed7K52K76omcklaBg1yo1XnhcozLDHI+JgC6J6VLeCd9Tmb6o7QaaBLCgSQ2/XzdRQ4eJV
BeUSWg0vV43pYws7Xiv8aKPAyWtSpjeAbSSZKnMsKICquuGFVqbFfulCMAyk1booh/Ung8QRnSGS
KuNPs3db0a2pN0tTfntvOoHJRJavgpHCslUZllZClimJeXYeCFfow1TiDjHtQ3+tyXqzRE8Y9ten
3SQ9Q0Sh+apazFy558sQXi65kPqwP2tzPeZJGW4X6xCndWWzy2GwlQd7+U3S5kiYc6Uza6oeOGv9
9c8X9+a3RqObJPGF0GoqM457a0T9Z2TiLKhWG54YY6wUB3AOJD1LmMq0UhCE3Z487dr9elmVLX1+
WMGYlnf9xyfj0LMzegjCz1fY7RSrXumE1pIwAzFNfl8itLWLYHVjnt/2zGs/Buy9sdXF+to96+56
9lsFKrrGYcUFTz1FRpp2vBbJsmFVDYaVh+4I59q9KK81g6TiKYGvU9r7OTgKVHPElhQI5blDEILW
eitJikFGgklY/2lbGa+SC1TQMuuDj8QJx2hhuGeJKvuJMeH6WpJeDnzl6DJ5crMGvphP4MRfrrV2
emCo9eoTBEGlRn/4V7m660WlSg/G8xmmArnTzVjLpgGeDMoGp2G/NxzmvX+Wvo5IuYQuWC8YFwdM
T5mPQMiVEt2Nfh8O64BthLJ6WuAr+L6G7sRSfzFWVl6ob048SG7Q+TYMJkVbG0ofGTgIW7dhLsmn
pDIPEYZdK+oimVIXHCRmW2hCti0uggbAHjtz3DfiSBSSHTxHvNztMyaZ+P2+1L3IPczVoT7NVmx3
H6h2Ty+GsE1pFYT1w+WCfvJWhh1X/kROXHCyxzcqhvk73lKKjY/masobMncQZbNuSESEGWay7aTa
RozC9QHicr9xifqpyi9YFz+suuI/pIHfQIfmaFoR/2vlp3MHqvj121CmHVoU9IH5eHs3nnalbEh2
E7zO0Mz3FqRv3oAeLJdmCXsLmiZjyRFPgPuc3e2+rIEP+5mS2/OthPVJhR3a3TuJs37XbePYrHPD
/ADrdFDyTvzgOQjaSkKeQcP2GQOGRWSwN9nE3sAygvZOfavG3eUUgzEEP6XvHHvKYILbPrR2Ysjq
Z9Uj0H3zjDawPD21QlpEtQtkqveZXIhB+p07duOqvNEtDwQPIyyRyU9QrwYoKEPZwGadcULelIFe
Kk2IebQHRuNQzzGWg1ltyBSrLUoXttqC95f8SMaJTBlBPletu/Oakvo+Rn23MVRcCM8Lho/TvdRs
yu7nZd6rb22edpzidzvyesZ1DqV3RwoUIP+hRBYeadIplxpsdSPpyRfTYpzyAulggh1j0ajff1or
Du1a3aJGbLyfdh4DmpdDP83j5IMzOs1/Q4sg0YmXxW3CFnIU9e3LNhRaejH2kyolSH/E+ibRzwpW
N93/qhxFGCkCaVVYA/u5LOlfU91DBB2/ajmxlIR4cFleZtvdKUGlCkS43LlX1tpujoUnmKoj9irp
g/rFtVGzBKJUe70r6U1O5U4lQHQwsyX+YLFIpSk95PZL1nxSRMYr+B3EBHGiG8GYj00AkOfvoS+o
vjMwj6fDKWm3pbDMK0BkiMlfK1oCBjF9nPXXNg/bOCMNfxWGVZaBuExITvj49NPn9I68Giz1kWYT
X6QqJc+ceww79ZRkzpNZsoyrz6ZqFQtxQHWSGvAPP1eeFSQVAFcRK+2c5l0Vew4OpVDFKRdMloYN
+Qt4fclv90yW2nxp4FqwCEtXfQYn6nFkWj08Ze3U+uaHEQ7s25761ijLTn+wzWrR/JrXq3sK6Jze
q5EdcYdjqARsS3Gt1Ps0U4wLiZZAI6e5HhcZbXJTjBr2FaD5pCeBC7YeFhxDOCwgkmsSPKy6XmI9
rDnqxuMQR4qjH6apj8zGeava+HT5QcN/pMujzoFKRkjjXumDRpYgyg7uJOEEqZSMcqsaha7UE9gz
6zWy/vkHIpM5QgZ4iCBpQhPA1IYy1ALQdivygTH4PwBE4ZMHH8VAD+XyIUkflUXNEujkxwqkDxK8
xaHdAchu1ls8TpciWrlEobPnj8f66BHkefq7BHE45WnJ/yZwbhZEnZm6cQxGn0fQGoNUEcX2ve1V
5agqqSOcxdC/X1jvSsj4wgZjcRZMb5B07u5m+oGOgftu+8LDb5sjPBhQ8jsw2sSfrC7Yx8jw5XHH
BRK+M0GY1dk+bpEkhXYoQEDCzCxxx24T0Ojs9LkZ2lQo521MBEiua50RiD/DUsNCo1B7/qu4QLXe
3m2XZGjzjoezzFsavpX4VEbKJZNfFUw2h3Fj1t7qFAyKV1pD4S0IxsX9tGOAzthEnwHPVQXF/lUs
BqUjo2Qwl2bpCgqU/BtwXDaZX4ZApJM0wDIuPdjx8EdKQHZhXXAr4e8MwWu6K5x/nPLYBjERsZNi
f+MZmYorlynHyxDC6PSjx3u0IUnnbPwOQmj+eTBPlNd2lbt7XQVMNMMD5j8vsAD6KM0SKll0/xFk
X+R3J7ukRNLZyIOQlH0Iu/RsiDMhuHI4siG2gwb07qq8pbT4F5/XsCLSKhvPWpqdghF+yfZeBWSd
bAfZgY2ItCOuigWuZx9AlXLO8aSFFjIoryCteN2WjlYY1q4qQ1xxKG9GKeF43GNtLHj0bxjOYFy8
Q7rUU1Bn5QfSicotONCZmWiGKt8t7w4VJhH/ShXVyRfLQ+pXFS80pS+0RclkyG/wOt0Tw0OWYyln
DXW2cnVgVV34vXwZfpE42hqys4Tr1SF359E/6c2K5h0VS6MqD2owll7L6dQtuFlZjF/GFFS7B+pf
/3rprPG1URYl9p9036ZMm570Jpy6fjXShuqMNzDFc4D+h9dSLZOOiJWMgHA4ou5BdXlaNM0MTLne
KT7JUzD4FG8KFIRSGieC78Yx00dqoC8fMTv1R6vTVON3jJyDqeTepM591E8JWMXlFU5D7LgB+LzG
SzTrfb/Vj1st4Eurh0g6qZRh+n4zDG38AZZbQK2gLqo18fYwLbEoYVS6xs56LaIhUaZlNPwc8MRi
gw642kkxR5u354WqBwl1U/8pYkxwk6fzECTPxJlBOl0G75OqyMOcJqiPEFLmpZqPvIVed8Xh44U3
8dBLqo/jqHbd4y0kIrzDMbKny3TzXOqEGKfueNK4IGqvBJqxvINLEO1bwJkMvhauVp9zO7GP+e08
j4+1tQi8HQM8+5S1Cydu+XKcu249UPVzE+vFme0SfADGm+noAiZ0JhW3bIJ/tHPTaITSskQg0nYX
VcLuk7XJal/AqVxFYM+DOI6ocLAfDbOM6S1EfQ85ASUk1Ewq6y9Kh/y3kE+2pcoEnD36BXP/rEkn
o8f/nmov4BXp4Wg2eQVAEzend6w6vp4RvIWT1Yoch8+DLdPXJ0a1N60323VyvzTVkKWD1Htpg7Fa
kWUwWmSYynwoC04oZh9ZcFULvwvugvSK9bw0+7vKXlAYNj+tCd0b3DW0MXofj5zSa+Uo3hoiwTmE
4TY97QecFL4Pnrq7R5rvn47JTVdKBCSjIxABLzBh9RnuhDt3cYHZivMxHRMxeadIqM0ZaGTOkSwV
KJQvlzg0K7eYTt74YFEjz+4BiPEDSJ0BDMshdNhMwanwXSi3uxwqZK6aDFEi0xKbDWmo299qK/Sd
ZTHbiPX8UI1qKmclHoSAQJAzDQgf3p6k387xFo0qtH4XIUgS88oSU+WbZUqlPrDgUIu91dqVSr9a
PvR34mXARg1SUm9kR/QOdaTFUoE4UZ3+MuDkd+p62zIJlWJn+qkvTi/l+e9M2GQbcB6TqyZn9e/D
nEJIbK0VKGGoLfOKPO1CIj7dliiNv9pfPcSr77MyJTSAzFcXzRwC3fU9ymo1RbKHnwGYHnwGK/Ja
acKuETTZTw7GXtWUWinTYOeri5kb645ZLaYJuhLkydzJSDqnZhz93VPkwiFcKAcAu/TbVnISwT4+
kQayoD4yYgPR5k4wloOGXfziiSeZpdCwPhfzJ3TGGYFk95CWgpkpLGgkRQwySKoBLkZN5VhdNL5h
2zJtlLSAfyVscz1uiMpIZLOr13vnACYpNq8fPueUJ2cx5W6crYC0x1E+FSqk4WJup61PAHJAe5Tl
6Ayj1Yu6q+/1RGoJgWFGHxUOnoZH7AOJTlzV11TlYqQq+pdY3AkyOl3JnuUhA4K92dNna/pAMBN+
iKTSnzlvDPw7ufsPkLHSYbJWR6YjhBYjhfEK+xqS35aosXmgQ/79xTQXcFgbtPDTJGKoXTKiEYSi
h/FjTxAWvoCp92auEMwjilFOxwCOUxnVsx9yM7+LVNqD7izLooLSbBAd0IQFbVw410kItP0iRblC
KIvU72CXBvM7TsiQ4WXDwOuRChd9dfyOzHKgAWib1jTpfzl4Uj3Phc5Pk0nZvZRChedm6JdelG1h
E45RcbYNzCo4X2nbSkpvrf9syxtoyTTbZRbs4QShS0n/PKi0D6vFBdEM/WHsuA9rQ5pmL8rjwXKy
3iUKL3sOZx3EzXKSgKyD0iIxZYkq4EhrS+8ILnxp6YUgPVeDABqJXQGK5QQA9iENMAU/fqHb4ktO
pCIkgipzHyWiPmi3IpDX
`protect end_protected
