��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��ЎW����� 1\�U�
��4}#�õ�~�p�	�dH������M�,��cE?�����y������uz]z���ϭ	�q;l�n1%LF�᱙ޟ�1��;�����T\�|J�d�s�w��(�^�AzF}������aq��F�]�K!�j=�*7��I2m�p�̳������+Nd(����UE2H�4��%�-�D��\f]|`�:3:��/x��_���aSrv��J�q�p�Z�y��	=ߧ7̨n]�hi��"�Ƒ���<��B����C�J�&8Ua"���',��*�JxI�f��}�܈��xÂO����8G�4Ob�0��E��M��u�;^v��ݤ�(9�U���7(�l$�_��c+�y�)&�xs-���Oj5�� ��t\�5}kȃ�CH3V6��^� s��:4;%� $�]lb�ᅇ�Dʒ��ɞ�6��ZZe��<KͭB���l8v��ǿ�1�>+!m�N�(�����"'qu1ǟ���)��E�S/�`��2�����.T�Zu�����ϸBC��g�4=�e���o
���+�3���K��9�V_a���>oK�;)bs��>��ۛ1�2��p'7��ʝ��+5�:�^��L�k�j�f6�xFa�~h�Z��}�m�Ӝ^�=
�|7Ur��Awƈf��}U�� ܫ�@f�X���e�%cT9��c�K��?HSS�l!��$o�w>F)�`$��
��dJ�!+���<��h��Y��(K�����j,�~�S�$C�O�Kq<�|��$�m)��<�� ���7��^�&�F���S���%+S�5=��@ߤG�	��-��X�M�����S��*���Dc���0x����#I�Ԇ:H���T)O�ܵXĄQ�^zor��S�G�l΋y�x�=6��w�5�;Y�/l>"�:-���҈���<<|π���3w�O���R��Fv0&��n�Y�"�8o�E�x� �*R�����ץo�&�M4MMQ�'�Nd�L�{l��)��-fu)j��������CZ��515GySY',HƬ���V���_b
��4�1���!� /|�tT���PT��A��ЅT�P�y�'���ŭ� �7����b����Z�f?��>�Ꮛ��Ϡ�� Ð4G�ma��*�����/���{-����uɝװI�h��Is^�D�l��c"^O1$��J��O�e'|����e��b��CQ*�"+6��1u�uL3Y��BHR�F�ˣ�؄O$�����w�}Y�C�����,X@g5�/�+,�p۔p�Y@r׀j�Db"9�� ,w!�b��ʍ>gº�v�j��^�����h��l~t_����%����@�e�Uxn�F���u�D��.0/�&x����oT�|Ӎn2'W��:� ��&#e������n��ʹ��N���7�Y譀]�Y�p]���X�(�]n]�*ؤN�����
�~1?��3�X��������35����^� �#J�"��l�D����a��ϳ�9q�DE>G�����V�sw�\a�:?�r���j��}��1)���ן�:(P<�/�9���0��)S�<(3 �2��O!,g�Ã���Z�o����P�������-����$}t����3��l n+��J��i/yO�x,`ӝ���g0%^�u��\Y�)���,�"n�<�=�6��	��5���?ߕd�p�Y�rf�لL�v�=�Tq�UH2h0�Q{��.�����F�כ;U���Y� �=-- o*n�\W�y�/����$K�b�̝�x����s�V�t��ڽ�:�7B)��O]��H/�ө����X��(ط_[vy.��`���<l���J�j%�b3�+n]<��ƥ�B�xBe���8���K�n�ʾ�W�M�Kkș��l�v�ޥ�B��FFs���J���w܅�g�\�Ҝ������%�{�6uq/�2�")+r�.�� dn!6�>�&���C(���gI�c� �d>fw��.^�dꌩ骮e+�9�BD/њ��}������W�DYX�.��p�j �8���	>�>d#W�s'�/�îM�e��ךh`YbH�=��IU�-��1�.�m�Ry��Z��2I�32P��'��6��଼~,^ZTH��v���9���_p�ؚ ^yP��>�*j{��%p&��ڼ�����Yl�~K����k���*i���D����/H|z��6����;x� ���|��m䣷2�5
�r>L��z9� xT�4L!�	�lQ�@RVÿ́����|۽��IB�̀�x�{�ƙ�N�L�,I�<�g�vh&�ꖦ�)�g�z�\�!ܥ��u*`��ɱ���D�\�w6�zS��Q��Q�W���gO�"���z�|֙�o�jk��� ����$�\"�:g��_N�SU�*D����f>��p�ͮ�K���;��`x�Z��]1L�b���kX͋�n�5����d���2��M��D~,d�\��7`�@��o��ޜ.V��mQ5"�삽2��n�lmR��9C@�2����o:��X�ԦhZ�nx�<�ja��{�S_6��E�;;��b��+��,�k�P�j��8�+8o�R�Y�����5���(��q6����>o��	p���=��l�zVЏu>~�e��ox�6�ܹ5C\��VJ�:���xq*����G��@M��	{�����b��.��Q��]����j����j���G�e�@*�ي�����	�e��Q>A�����m;�-�XEίLx�,x+���#������RD��Tr�2����g A��x�@1x��=����9^DՎ�%-�n�b;���m�f��ǵO��a�P�GU��C��*(\{�M*��� C�/9q��kG����j' �5��@nY� VP��<�����	e�>�J�	������Qt����b#l�ɼ�;
�K�.��K׵��D���Sr�78�[�%�m�;o��J�s��ր��*��w��@C:���_�c������@���W��c7oԮ��$Lm= �0����J/i�Q0���?�r�N�VL�b�VI(�q�Ȇ1��r;Z��5��������:>�/-OH�Qrn}~"���4�"'��`�����%�*�g��j1��U��_�Vp L�G�������4�r9���#w�=yG;���Q�e�g3c�!���t}LZ�G�+�����Bp�o���b�#o1�`:����X��}B8�u ����f�U\�	]j0��휦�dg�[}����YyxG�g�����˩ph�(f��.ُ��s��S