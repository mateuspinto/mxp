XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��4����21P#xO�O��3��Ӑ�����(��=u~��:k�K��}*'�w��K9���5�~�{���m����V���+so������}z��a$��0�Ǹɓ�}�T���t��4�ϝ:�N�;>�N���x{�©��C)�ͅ�e��j;�R���g0��jl�!��4�v[K��:q�w�dT��m�N��{��N�u �����*Z�i��l�M$���9�Y�D��r/&�3�W����	�ߒe�aG�S/��Kcy�ѩ�nY�3��xD�-'�C�'�&��m�6h���d��2�4������O�C�9�4~����|��b�r��nmQ]�+/��&�~aH�mZk��*��Bs	Y.6�{�S��qL9��8ا/��nΑHQ�#�4ڸn�t\NC��N�+nh�y3�΁Ǽ��Y�P�}�A�����y��`v(R�X5�|�I;3�&-���Y6m��:�߮ܜeOݽ�U�{�o�X��H/�!v�ῂ�����\2-��YR�g^��˦� &�*���-�f"-�*�?������ѥU �	�$e���Ym�؂&d�"��4}|�ὼ�8s�r��-��VG,{��;;5�L^�a��@�Xe��h㈀g ��Ĭ����[)�cq�:w�~�Jvt��`�+�^���ߍ�%�?@���#K�X���R���VwŹ�0n/ɭ� �<*m��8�K2�̷2���T[q�g/�����̫<�� 7���T����	i\�Kq�_}�<A��26�C�XlxVHYEB     400     1b0�����/��+�� /'-�ᇔ'si��/�T�U�Q<���ց�f*GL��Z� ��4�((�==& ��.F8\F�|S8��k��6���g5��kL���~�����u�f�V@�SV���4�f]
y���i*:&pCĪ��&��T0�Qu���	eћ$������qR�ߕg����n�������ҥ/p����)�7��7�C�J!��<ĝ
m��Kх�LMhן�w$�hL�
����b��h��]t����0؈�#���8��p�f�X���5~��Tg�ܻZ%U꠾�?��D�D꜡ۈ{�غwFz���������3�h���?��@�hsa�]��-������3�X�-	'�����O�%<�K�^�b=��$��v�O��"��{~�[F'����oD��*ZN��a�XlxVHYEB     400     130�6Nꌹ@{@`S��஭����Z�mQ'\�I�j�騴HO��eh�����`7��� :Y��f~��-$�Y��E�LG����ΧD7�+B�A+�;IL}|��-V&�>�����z�n��bTzkAx6W*;�.��٬��,*:Ȋ�r�6� !��g��*��ܥ�M����B �d�g���1 X����!|p���ؠ(��\��U����G�	'��|�6n��w<��m�M�J��G�^�>N�1�2�7��
��E��V߅�Q�vs�`�8��EV/���	��R�N	�XlxVHYEB     400     120�(��Lg ,	y,T��'��]�<p�����Ĩ�^G�'���
�[�xՌ���}�����hh㟐�W "[���4�U�œg�Km;���]���0�so#���üۻ�jW=� *dDGݗ�HɟY���EH�B��7���4LI���d�FZcI���x�>�0���@>{;j��>賃]��3P#���G��Q,���Ef>YE���7ʞ��U**�BZri��G�n�>�0����_[!����tEh
����n�W&��a(�M8@*4��5���BP��\� XlxVHYEB     400     170:�/�)��u�2�x�~A�k��vT4�P�_u�uA�Ķ���6t?�9SY�E�?~
�H;-%Ii�e���܌���cI�4K��C��Yk*��JN����?�״�Iq%`N��nK��p�ݤKT<�*�GwҎ};�ʹx�����"�$dX'ycf 6^���܀����H��C���=o;��6
%NV�e&�j����Ӌ�@�y��rY�X����?�L�tQ��笔��6�T.���$�l5�N~1\L��ó�;�,qz�E걺b�+}	�u	�	Tk���j�©���{�(�Ƈ6M�x�`��	�o�f֓���܋k٩f�Ͳ�_�%ݻ��8��XlxVHYEB     400     1c0��:�T~	kA�k�[�.���˕�s5�<(3� ��JD���YK���QkF��BAH �ڦ��-�b��9h���w���pWi(+mǀ�	��U�L{"���j���ʖlEr�p!�70��o(��ɲ�%6̺�V}�����F�)Jf��e�	)�~n�0okGe?8��^��Ig�>��1���	4f�s�����`����L��-�/����7��-5�}��i˥d�m5�쨷�ƠS�����2?����f�=Ų�7��c[�o�e�f�VJ䧀�V����#uL��@��k�T)�z^�)�YK(�A	r������ɔCjR�����U,CB����U�0klE�t��ny��X�<tvQ%��'�M@Zp�l :fG<;�8i�HpT��F�vٴ�ey��hR�۵al4Y�H�<X|eM���jMS@��XlxVHYEB     400     170Y1�5���Ő�#Sj��PM+�����s���Ɔl���;Ac C�����P��ɛ�u�R��1��s���_����@�D:M��m˂���V�[�e=j7L�[2�����[w���7���`��-�Y�Q��l��Ye�H�qԥm�"ϣ��sH�בRz�v&e�����-�����/(��,���N:��8�����x��T�h�k�Oyؤ�A<'���m-p�*�-[� Q��\�>O�3l̴^y���o\�4��R��)��[�R����={����x�:��;����>�`��������|�zҦ!f����F��>:�xw1����l�ba��\�Qr%�A�0V���	�E�����KXW�-XlxVHYEB      5a      50�J�G�-?�`�'W�"Q�w���T��z;��ے��q(8�K�����|Q�l�C����J�t)�9LYE��=@�#�`d