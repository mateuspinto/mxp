XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���d��#���� ]!c%���ڣ� Ԓ'�JXpr
Dp�T���&lŵ�c9�GL��f�����A�_�sa�v�(�K(�>{A}�B,����4P�}��O�c[��s�w���������+�����0m,�o����!⹜z����u��B4ǿ�^n�)mŸs��%�Dď�$�R=`���	�s�Q?+�>H��32h�?� ��l���`�����I9�P��C&��v���@�$S������R/� o�2�[t��G��_�nL-Bݨ9i��,���\,����8�
kmf���b��T/����%�����/w����)�$�m iP5����%��o�,F������3dO�q��F�m�7K�'J	�-.2�=�#�:$��'���Ɩ���P���Ag���]9 E��M�TǼ(pI�^��/��I�3�U��\���3t.ْ�W=�[K���c�����Y\��>��|��ڥ7��	D���N���X�6S?����Wli�^-��Jq_n:�kU��i��auc��8��j8G�1�\�c��0B����_1����[ǵ:XF�;@�����M[Q�m�����<�U^}��a�*��L|�H${6�`������7����׫�	WS��f����ac�q%�ȗ�A��_����K]o���<PG�=�� ��wZ�q���1@���?UA�䊻p1+�۩,�������I�}�hBJO1�oE��A9[�0Ǥ�k��{K����5�;��:VP���������[XlxVHYEB     400     1b0�{���ڬ�֓7���/FϢG�# ��+���z寥�������=�{xg��s�N-7�E��=8f���/}�:�r���ՍZchx��2���g;�v�t�����6+�/`'kV�<$\���������[�K���	�E��d��3U6r{'�2Ɵ��J��@wJ�8#C�UZx�3�H�����O:�-�Z�́B)��$��k,m?R��'�ؚ2�b�<dH�u�fV�'���J `��2�BN��1W�o��j]��Bѡ��a�W��{�Z��r.@�8;��OQy��Eu��;��m���H����\�7���їZo��6H�.��d��!l�7M�QHr=�O�6����E���1r�#a[��4gس;TAj z{�(u��c��ՁC�lů�,؟��B�3������|�y�m0��XlxVHYEB     400     1b0�k�I�N�m�+�'u�b�b|ϰO/���RQ��%����ޕ��<U��[��3DS\��B�0[+ 
�.OG�/��q\|��=�PQ��]Zr<�����D����:	W�����%dì����F{�: WC���ɬ�>��^�c�qE���"� ��]Q��LiU2m�WBf�t<l�=9��d��N��{�{d�RsL�|7�<�c�nZ���_}����X\lo��CwOB��q-���ǵŎI�v�x�t�(p�x2�`�O�iM$=�K$;�W�I]�-��-a��q�"��_�ir�Va����Q�^�Ť�E�������VR%�������Ū9��h#�:�r~?*�lІ�����hm��v
�;��F���A�1g��mn� 5���d�I��A�t��-�$%{��G��*נ����XlxVHYEB     400     130R�r�����Y}�U<��.VgE�{#��E�sw��O��Z��v�X��fݪ�Ss���AȔ,� �ӱ�~�<d�̤/���V��-UO�%����M1U^(�_�h��b��6�8'+���.��<f ��'-C83�L�3E��	ܝ�ܩ�';
�X�DDԪ���Y@��Q�Y�-A-s�����X�F�SF�~�p$Z����(-4��v�3�1�4a�珥2J
7���!7C�B�i�	1avv�6d(�T}Qp
H,��ٱ��
�T���a,�F���.0��Z�,4�LVGXlxVHYEB     400     190�ћuЭVq�N������-���c��if���A]Vnޝ�A�vK<5��wU��L�jɆ��Q���3@�h'�h�Ɯ������S��g:w��2}����]�jV����vPa�>9⨊#E \hIe��7�А#��ɻKbĕv]$�\8�ĒN��� ���o��~))�T])��z������h��^��,�t���#��%+��/|�.8��G8��(������&yv$k)�<�L
�?���׋��{���瞼A@�mM��_^��Ӏ�Wwi��5z�`՚ �y~���3�6�3%�� ���[ֺ���N�)@C�\+w��c�%���G	3�9�IzWT`)�R��<]�۪�x��>�o�s�b�TY� ��~����w�u�XlxVHYEB     400     160Z9^�TzЉg�=UA�̅���3���yu
��Q-D�%���a��f��z;W��Bց��i�{o+r��M������9��=�=ٔ;ir���f��9�x�����O۞$�C�<iV����0�!��"���cا��/�LSH�$::֗j=\�<�xtVf�L����� �$fiLԻ,{@\y"�6�}Z��vx�m��-פ㎀��950�_��"
f�l�%����V���s�_�v>�Q�èy;�C�Q��S�4'�15�W�\[{��ȶ`���nk!0Q+N*7�g��P��r�j�Bl������.sz�<�"	�ܑ�*����?�B��L�4���
L�XlxVHYEB     400     1b0�&w݈þ<bl��/sn1����@̋��ޥ��}[f���j2��'M�f�������n��jPi�8[��ͧ�Ѳ�����&Ú��c��݂���P����׋��xC,6�: ژR�������-%+u�iX��(��|�6�&T�i��?�c6Fb�����Xq�����"X��6�JD&A �П��锏�fP<��1-�|Ak*t���{��_C�j�������sZ�/9ʍ@��]������pk;����ڵ��ߧ_$���!�Nkmx}R�S����5Wq��%�0)����U�'0���NG�Ld|�[�d�y�.Μ|�V*$: 5B��iT�a�<geI�j#��l!�����[kAP�\���4��8vJ2�&���R�9�t�C"�cDy�����#À*�&�����gv=��������XlxVHYEB     400     160n�|hXK��@y-�9��a���D��̝��[-��%U03�>�1���D��@��Ŏ��sp �K�D��Pm��18�4I �G.����d���^B9�,�.�}��4�@([%����j��ۺ�X�xqM6�K J'�Wy�j����E�<�������	���`�8H���+A���qRR0_�Q-5_f�>����j�۴V����*�dZz��[hi�����.�z��K@A��M&M�!2p{&�<���m"����!
c�9�C6K��v��-mR��>UӅ�"E�AT4�`��!���`����E�;x4�d/W�$�'�om����·rƧXlxVHYEB     400     120o�8+����ӜW��l����Sɟ�:�}�'��y��W��Mo�QC����ǎ�I�s8�.�����A$w�͍|���X@F�Z��<�56.�e��U�'���h~9�U	p��(�M�_��i��җC������K�]�/��sJ~ �.!O����f��1|�n1��O��d�1�53�����[I��BX��<B����(����z������/��
 qK��`r�qǑ]���\W�oxtķ�%�1�����AF��Ż��ӫh�*yȽC>��c˃IP��T���XlxVHYEB     400     190Lְx�I�𲽍)6@v�[��W������v��9�����?#{��&\����mid��G<�t�i/��3�5e�C=�,y�ə�e�Yjs�Iv���mu�~nOrh�+'��}J���O,C��C��m�U�� eJ7?<
;�-���Q����4[L��Q���[.���ɾ\������x���)e��ɷm�d����0)n�nt7��������ax<�i3�*	}h?�qg4!V4F,�mE;g���''lT~\�"��5J�X��֟�Y��RK����������b@v��E�C6/�X�5υ�0�� ?��~"/֮(MZcW^V:z�/����v�G�qV�1_�%(�Y*��_�[/#l�p���J�1��Pcu�&��� �
�g^�SXlxVHYEB     400     140/M�Pm���G��C���ߦ�^�glU�Q�T�cڢ���j���5��?V��m�v�ϼ=�o�X�I���t�:�`R�B�����C�V�]2ё�9�u(?�N5�� ��?�$u�m^��$�)�«t��c ����1+��Vo��֘�f�2��Uv�*p����q�}�pM�����TW������lj����e�Ѻ��ؔ
�U�9 l���<��WAq1���Z/�ط���g���_��%ް����g9�r�U Kgr��uc�j�g�)=��2��X�i��Vz�N���VC��n���z	;cXlxVHYEB     400     160UGM����"W��s==)�*�Ac�綿 9��zZ���w*&s��c����Ҁ��g<�lkI)�բK�}^�R���:�+�]A<	�7�G�F�/5���hh0���.$�V����(���E�3o�j0�%���.���+�d�5��p�n�M�N�7�J��7t���=��q݃E��B9C8�hZR��0#;(ܧ,�������ùP�n�I��^�Tr�ϫ#-S�ӭcy�[�;�Ư�vI�����l�4��3���k��;��,;��ұL�|$
J^��Lr��e��;�IZp�'rN�s�m�nm�u lNI�2��s�C��r lڏ��3��A(���O�XlxVHYEB     21a     1003t{�B�@N04.��hˬ݇���Yjt�,�]~�R�J�"�����K,>��a����u�려�e�u�Ω�n+�tEv|�*)�
n�!xO��B�f�!�<�̤<���ę�X��ʢ?������#�4���S��w�ػ���$[���^_?]yv�=VTj*]�P��=p��q"{�`�*a�Ae�H	�5���_ �q�syzG�Q��G��K:9�5O�79��I�Ѳ1�+(����J�/��j�