XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ô
�2?=g�^'3�t%�c�6�N�cd|���|�I�����o}�o�ι}��͢\g~ͥ�T$�ڰ�%���(������|�wf R�vƙ�9��<�!�c|oS��,�L]���8{ۥ���؅\/�\[�c�{�?�m��&@��H>�F��p� mZ������6����62����(܌�B�,�+����3���X�IT>�S�,�}��JQ<azt-.N~��ƽK<&��jVKZ.�lM�1�\߲�,�5>@�H���8�@w�T�{��F>ù���9U/S��m��s��S{�3�X��5["����R�%A����V�}Ҫ+��$O0�C�7����H"9<�9�-`�kK�Y��6�Y$�x��L��T��6������ K}�e!������I���N�x�g��U6݅ F� `��]����&�	��Y���K������yJ�8�tl:&�su���Ǧ_U�-˄+�G�1+�{�t�FY��h��k\�h`�k��
QJ~�<(:����������D	��+�}e��Q.�Y��������@[����ީ�/����
R�Q�"{ou�y���8|Q	Nk s�2x�:d���B��
���A����
�����rQ����d�������Դ�����}L�(�ϣ1"��e�t�	�-)�q��>3W������%.[�c���gbqT]TAm�Lm%�4l�.GA,?Ќ�����=�6 ���-6R���\�������|�)�ˇ��y$��A��XlxVHYEB     400     1c0B��o��ʺ�%e'F��>��!�Й��=���<��/AԹ�1"��`-��rs ��]2@o����M*]�E�mH'�2�2~ZVtٳ$q��0p
�'2o餬>+��Sٳ��w|�Y����V����oSA)�<�}���	T� �H���	�Q1;^N�4�Җ�9��u]�mW��f����m�|+V�؁��O�L����1�h���6b�/��ab�Z(q�ˑ��v-�U�8s�� �f��aT��q�u�,iK{U�%<��6?�Ab6�����ߠ���#���^��^���?,q��pAںX&�,�-������O枤�������K,��$al�
D�k��������F�f�߀���F�0}U&�L�Hk���P,"v��;a�*R:6˔�Aih�&�>�S�(Oǿ��?]LR7�б���̑S��&SD��uw�p��XlxVHYEB     400     160�uBG`q�+p��dN^�pT�-.��	��i
�o\�����޶̂Q��j;�0���P!p~!�#J�}�1�T�W��XY���	r�+��/8�>�~��S�9�T2os�#�+��:�C�G�
�l���`�ԙۥI�{��%�o�w�����vSz�H��(�Z��Ap�Q��Q0��3���8���7�Pm!�/ �h[G��X��3����K�C�.����b�!;	L��Kl��?�$����Yt����N&2�7n� �Uw�BR�
��
ʀ'�Ƽq>��o:;`����6	yh��g��"�(A���{F���ڑ7��q!��l���3T7D����W�'��8�XlxVHYEB     400     160P�܉���HF�� ;Ko\���y6�fW.��s����Ǯ>Wv½�la��R�k��&aA�d�� �6;C��g�h&�2z&23	z*`~����./ekW>��LՍ�Dϣ�G�K��Ҡa`����-峓h�e@�q��UHf����{����z[�q� �+]�ʃ � ��.�jP]H�h�&�8,�nɟ��K�ֱw7Է*���u'o��}�sl�/���\��ҮG�r��D̎�L�^=Av�_JZ�^}7��@hT2c����H
�d�6��ݬ�X�b �}g�p��/��Y������t�6��3JЈUb�P׼��2��Yo�8f���1X:=�u�aY�"�XlxVHYEB     400     100�j x�c	�\��th͜�C�>H�q�Q�&�.��ޡ	�H�ZT���{	7�5oЮ��� C �F��PLjL�\���}�^��*g�*59+&T�E� n�C5��D���ر�zB�wX��C�އ<ͭN��Rtv����z��7Ȼ��rŇ]�q~zэ#�̚iM'��Iaq��L��6/�A^��Q;9���\))�ta	�L��9��	�r�`S�-r�A�v�k��B��|���3u��x�����#�&�B�XlxVHYEB     400     1a08y��5�3�2�>������b��"�0,�Б�*L���)H���:+ag�1�\���ʻ�¥BQ�kF�M�5�]�<��u7�#jn�s�3�K�����\.����Ꟃ��M�\��c��5�0JƉ��fK���u;���T0?���F􌥇ZN@}vN�ۭ���a N7iJ�z���Ng�gh�L�8����1���b��I9�O���8��Z-�Qހ��G���3��J�&��\Nb����T���2�{De�H�-�gp�q�R�X5�VB���V9��}w�������˹��)J��� ���@����E�$������˭}��
>\�V��m�*�l��p�������UAiO���q2�1��������"���������"ԩ}˼��6�Ć�Q3"�+���X��)�çNڀ(XlxVHYEB     400     140i�5�5�����,2�T4/��� r]���F��,��x 9��Ϭ�����������e�N��%O��bH�w'�JJ�8���uQ��n��#��ue���:,m��jUN�L�Lº�Zoa�V�%�F�M���Cv�/���Æ��^4�]��G�T^�����R�#jy-����_� ���~G=����-������ ��"��B�辪-�yە��֏�_��X�I��r��_�4�}K5V<C��OL.���G��(�<D��<�����ˇ�
p�5x��bCH��p}F=�-wLr˺�w�hբ����coLc!�b[tiXlxVHYEB     400     120�kK�m�:�G%̊N1K�?��������`����)䨧��a�g�`q��G�8��\�~��1߱y{o91�V���*��d�' ��JXL[��u��&H��S����'�Q�h_���^ɜ)V0��{��'���[l䕉����+x�N��%�P�'\WqϬO=��L�Vnx���,�tr5/���Kװ?۠�~��Ģ�(e iڛ#�������n[7�R�_���	W��<_�ެ�uGE����gU�ۜ��3�{"�-W|�pFBX˳a�G6XlxVHYEB     400     130��%�#���3��Xb,#�*4�s�_����.c,�3�o���Wd��IԯXŅ)à�Ip?�Ag[ɂ��O�( ��5Q]Q�a���]�ْ0�t����,��k1�H�>�����R�S�rn�f#���i�c(p�����w���1��qQ7�(L7�X����>���R����L����~����i&�8�6�0P �\/�l��_?�;o�:Ǿ\�-�{�0�/���~�늨�"��ч�	���at{��Z	�eL�%at�\�+2D���0K*��8a˂(8��G���ӕ"��WR����Ws<|�XlxVHYEB     400     1c0A�QT�!�A�+P����Ri���zy1*� 6���8OC�^��5����w�S�R4h�s�pu��|(B���Ze�",�F>pL=��~P��8@�������us�+8;9� [Ů��\;����S
��5���I�*~v^���*�����o��,����-`%!+���K]�����tɼ�"�����rq`��ͷ�	<�Q3�.J�x�f^���ju�V�1�`70��ڟS��K���>''����JLg���]�X�
�G�/����eY�����(2�R�}Rz��RUp;Ε.�Q|l�b����:H	�v��~�[�
_�v<�h$��F�L)�N��I_�Q	X�1M��9�v�d'���͌v��JK����<Х[�h�h%'%&�$��$��]��>���B�w��@0{�<9:iy�l�!b2KՎ���BBȍ ;"&XlxVHYEB     400     1a0�� 6����Q��2�t"�e�ݐL�*���Jt.����@ヱ��]�5T����`m�GsX�/���t� ¼ֱ�Tg4���|�A������l.��[*�L�7�|�}���1��~��Jz�Y��f.TF�lH[����s�� ��/�-L!:E�&���ym�����ҝ�o���ɺo�����Nȃ�x��MД0]�	R�t������16�K �|w���������.࠱��r�R�R�� o��x�|�n^ ��� �[��\3~e���&~�)�B�5�P3�B��-�U��ԧ�aV}^�j�e�}]ڐ�Qn�x�Ӛv����xBޚ�%E�(�<�lш�D2�z}Da4��{��=:�Jbh�S���!k��k.��6<��˳���* ҅Z�� BXlxVHYEB     400     1a0���y��V�'���x�	���t%��kY:&
yL��rK�vlSmT`�D�`���������߲@���l��:�έ�UF���J�
��Ct���Z`Am3ؾj�񄪟��~�eZ�h?)��`?E����w�dl� �R�UhE����z�{*Ur��
h	Q���.K��9�����#s(�)�'��{WF�M�I�V�����\�f���A1���]�����G08�	���}���{�aV����+գo�R*�Qd�(�z#��R����n4�^���.s��{�_�����s.�0p��*{��_z���ul]�����$�e�����Znl��|k���ю���ȕ�Rb��<m�_i�%�1i�W~����%4�/��a�i .h�����,̙��̖�XlxVHYEB     2d9      e0��A���]��1{vɈv��d �I��1/sέ�5١l}����e?��6�Y�/�ྣ&`�P����D|�mƫgel��Msϑ*����ZK��G�4#<0���ȗI���a͎Ɩ��3��8�F2m��H����)	���t2�l�%���[�|S�7�/}Ղ���\�x�����4�(𼂤T���C��Έ~�n�&�q�e��s���(}����R��^�f��