XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��� ��:�A�d�X'�A��ͭ��)k�d�8yI3�sϗ��\���X�/���A�Q���� ��z���ӵ���}�98"�c.�%�vP޷�@c!���o�Z�P�3� ���6��i/g����BY��?\��p#�������o�2�+�[��<EVtDx��ŕ;��b�5��/��$r�a�'"��>@���i� [����n1��
����U����3E�[�?�	��Md���r��-���.���%�$�l82x�RRo�_��Ϲ@K�0]�����s@��>�)!����{Q.R�-�A��?G��*^y�]I�Sqc�oQCҽF��fn�c:<v�(R�D�7�9A�w��@�8�B��I��C�@F�HX�������o�n6X�qI���6�����\�^��V?�/o�����:�i ~�.>:,�X����p=��[��Ì��e�OqI���_^iӗ�M���zGt<*�.�����p�ۀ�F�D�u�U�B����8]��/eIsԐ�2	ב$,�Gl�z���3���S���%h^�k���edB�j��v��Z��m�&�@�#��B����;�|c�@|e4��`d�}�U�@eR��I��jF�����5S��̽޹��b|��k�F�	Յ�\��A�f̒��wK?N HEsF	�Y�,��)=H��=��=�k_�ޘ|�=-ehG�X�K�*i6f)�~���[�:s-��,@a�{�ɐ����e���o,����G4>fGi��տ�M�XlxVHYEB     400     1c0�)��Ѳ��#���،	S,O;Zؖ\w��6�eh�g���cϙt�y#q�\�"�)l
i�?5sCظ��JԭylJ�VJ��Q����֧�:IFQo��QY��&�p�C�r�.m�� ���#gB0~�0_F֙K���n��o��n�&c�b�<R��P�t5ɿMI��WA�[7&��( 	t@A7Yˋ� �������B����PB'�@�ܢ؇�����Q�Yk�j��Ǘ��M�w���,G��v� �C�LK�IïO��9��>�5sh
���5N����O�u����awR�L�}r׻W�^��}Q�Ϟ̝w�>�Uf�>��!����=!'�5�_����ʝ+�/���!��y�d��� ����Kc�,���~��k.�Ҫ־u�z=o��> �[:���Z�?�8�L$����y+<i�Q:	�[��YѧXlxVHYEB     400     150��"ܣ��)U�>���Hk?18�I��˺A2�&L�!L��b"�#a�f>Ct�Ƃ�L�rZˣ���`����g0�)��x^p�~S�}Y
z�~Jv)!y���@{�-o׹A�O>b'�~�����~����d�EOo �]I
Lr�Iݷ��,�����ɀih��w�	�(OC�Kեp)O�"�A%�xL����ȲOX$��{akĘ�!��H�v�9�-�u�>��5l}�y@0�V�����m���~�Ӂ���۰����AMgN���N��1���u�4)`�BV5���ҸjK�S��qq�AR(^�Զ��
V`Q��v�����He1��N����XlxVHYEB     400     130��Fi�3��V�4�s�l*ˀkD����Qb����P������U�{�]�Hߌ��7�<����)�Y�K�V��%�T�R��^q.��,���so�c���Z8��Z��C3��������d���E��6�F�i�Ę �SfS�R(yP�7G?��*���֎�H�h�͌�d��fB],�iMZ%J5����B:��VEy�ԛ�c���e>�XP=Q���NR]���Uz���H�{��`?�l�j��y\F�6�B[��|z�m��ׄ��o�O#�?��V�+o]d�l���E4�XlxVHYEB     400     160\	��F���go�ѵ(��?6�T���BG ����#��+�I�?�#ҁ����I�F�4���ȋ#_�Jw�n����_]CD=�9�;�v��]xo�p����Bн���Z�N��X�
\����S.�2=(�.F!NO���p0C�@&�eQ�QΠ�l�y����r)_A O�f��8+���r�*��������NB&������ ��&R%~�_6��f~�;P�'2��<D���L$�ʄ���{���̟h�C���N����Xt����<$�m�a,�ڴ˩�Z3��Ӡ2:>iw�r�O�
<�֖�W���X�Y�R\��s��SZQ�T�������R�Pe�JK�op�V�\�ʒ=��XlxVHYEB     400     1e0ȜC���-��3��U}j�o!�S���-�	��ϒk��=�M��s'*���'A;Q��M�<P�(�y߰��q���ȟX�iZ׿�����\�l�j���F�nD[��t"�G����J���k)�V�	I���k{�Jn��R���㺾W{9��o����0qҋaY�1�����{L�N��|�`3��r�g��RӀ����_�ym���(u�D�*��r%���l�E�Wl<5�˱t�m7��v`}�Sa��b ���,�9fY���4}z�/�$X��F��e$�X�H|	���Z�����)�+n����swW�@��	�bVD�'a2�g�׏�f�;���{��m1��O���vv���v\�A8��wTVKzh�����ZP)I=��Kw��ƺ[Iy��>�B��˴O����xC��.�F�M![I�r)rf�6j'ZH�%����[�����=C���}�����j��Q6aa�vDXlxVHYEB     400      f0]>ű�)�F�?d�G,p��2���
�.�]���!l�M��Т�(�=�ep���A�w�c2������׶򇸎m�y�����>b��UQy���8pBF
H� 1�E��e�� �Cǎ�6���Z#�[�a~�Ƥ��Q�c(m�7b�:N�6�p��5�^o����z�`����ZHA�1�i}��L���⫙& оQ�|8a*�3�]p�䰃,UI���D2A�ؠ���~��EgXlxVHYEB     400     150<���D��d�	�W�����mCY��/c,[Ng"ݨ�Q�(9Y�ĉ]����j㭶Ͳ|�w�j��w�~�GjBN_��"f��al�;)�ȅ�f~�|����4��hy�>�~F�#��~I��S8�Y w��΂d=�N^;K2 �tj���ӂV��gz�ۥ~r�C��R�ĝ��:�cN��8vv�|��v�^�!gs�y�^�b߳T�~(��7F�l�䧥H�Z�l/*O�\����&�o�*:#بH�U��:���Z�27"]��(��\+Ďߟ��ƻ�~$�JƱ���RS��v��H����g�5#��6�'H��؉XlxVHYEB     400     170�eE�b8K@�!��G�򚸆>�+�U~a��ښ_����]rI�(��D��k�PF��WG�����c>�*�rӦ5n:�c\�wE���
Ɵӛ�ʣ��Ԅ�����F*C����K�A��~���D�3Ȩ�v/��b�,����)�Y���6�h�SQˍ�L�﹄z\�%�D@�A���	�
[�4�^�'�S����p��(�@q�n���yr�ʟ�P�;�Z��?<V�u�_��"m�/��O�����-�����3�qq1T3Q!��!����^�
�Z՝�(�I� ���׷�����T[�b���D��B@11}�(��Q���ދH�Y4�@C��q�I�ٜ�5X�3��*����A�XlxVHYEB     400     160����U�-��]�x]���H�6?����	XtXL��6��t��)]�����P�����c�8�ů=�舱*�g<�|;+'�E�;���P��X�;��)��$�f����H��l�
��v�{�fYt7u�U�tq���au����5�O�+p�(i��Z-����r*����K��D+�v�?G�ݷ%��d�O��i<W�	��9����.41�	f~�j$X�Z��K%���(כ�R�1�(�i���H}ղKd����z�iS��7��B頭�%rx�qD��ln���+����دZ������ӧq5P�M�"��(�h�9!��[3^��n^XlxVHYEB     400     180����(K�Zɔ<�Zg��F�H5�IK���v�ϳ��?b���/l$~L9p���.&#���S� s�Y���h^D
 C���[$
��@��F�����p�[7f�z����Q(���+6=|'�IobɌ�j��-�Q`��6H��2x�8��x���aH�]?��9�Bf?aS14a�@�\����L�Tﵻ�<�l�F��d�?�8�����Y.�@ S���ꅻ]H���k}�\�����!I_Lp�����yg����%������7��6�Nfh���*K�l�p��pZ*3(A47v�>dQJ���[O\�gPZT�8o�
�̺���<�KLR{n��|��i����cm�(�C��1v�m"����#���rHZ�XlxVHYEB     369     180;u��;��yp�/8?�=>���x��ƀ���z2��4/ԥnE��k�������J
��%��*i�_Y8{�n����Z�DS���F���f����[frBe@�GG�t����=��\j V�D��v�_bA�c�@�����gE�D��gȂ��^�LT�n��}��� _����p��+rG"��-�A���HɜC�0����u$R)|�;�CҎH�:�h�����g	�ߦ��ܾ<��!��mӕ�C��B����qlȍs�,����>*���?����;)�Ӕ���Ю}�����V��~Vm�u�x�p�tݿw3<v&w*=�*&�}wZ���J�j�uf«��Q���es�	w��}:����2:��GͷFM��n��k�