`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1120)
`protect data_block
eOevkCwOZGAt58xcTufO21Z9y/lCektJxnsaUNw18dz0CVT7lKxHtuqPtgRtGJ0J7Mm1dXZpvV1N
pe09dvaW5WaITUMuNzwkC7y2/nVYnyLoqHtUh+y/vjh/v/wiaAxUzJZcOGXH0RIi0sSRcCv75LE+
DKDw/yN0Oah6n6K9mFaSivW1MCOgGOFpU8Ah4QjI2LWnuT98aJZxHjwg4QGAWVD30aBz5veYd7Gb
MMJV1voVjQH2fOC38bz6aFnDY+AwQzzdAgkjD49gjzIJxcs0Um54YIaYV5pjbfZhrFhsxkaBOj3N
nouU4QEFMD0gA54FgzlkEesGTq1Dwz85CbM1vVmAJoiv81Y8P5JkITorE1hpTzdnIzqp1YV8MPve
PHSaThcbeWPWjF9zVmodacSFtJtVFMhQrQIdga2TP/W8seTK20iROEYfM/dXO4O741GU7t2iDayb
Aq2806JENMkl/WgsyoKDsfL4EkJ4OppAmGgAYPxG7tslWCXEQZknnQHAbH7Esa2EcoJUOz3oJG96
KXYz3THCENjW/ggyffQQe9toVeJ9ysIUyDZEAiIHrWf71rFKFVOSkZAMLHi50DubWxu2ANozfgOv
QpyWR2mwZQnJ/RGtfNOizF2qE8nA1/tGLfKH4I5P/+VnyzJyqoXXHrbLs9n8nchHM3pYctRQFm/6
0SzdXrUiCq3HjV5FqCqXvHIjewVcTql0UXWpzmBnadfqw0p4+1ovbEeoGrYB38OOvmvplJsOQYqh
GMmTJFcSTAnq0m0gVEKdtRX3HdunkY7J6cTc3ZvfF8Zdv1SPuOE2Dxo3gwcVuI+8ucB62+inmeue
7iQez876p1ZttSrjj6ABbb2Aima9cMnN8hcie+gaVrdGNr6evQ21glrHS12qbNoZWx0Pp1/Rb2S3
DgAakh8LyCCvOzlwpIfbpFbA/ez0P/okDuk8x8rII7UYva4LObwafjVy/oQknm/uNoWSLFD9cH5X
7zhV/EKUWuJ/nj0nAZtCCH7Mk7JjMYR+/lsBngha8j+5JVsgxTCLXjfcUi3RwpOcSihutxjmrJvE
pXyJVFoYLXqC5Jz79G8JcIvaS1zl7VK55rEZCX559TRVPQXBCETVFqC2HoXEQZqZOd3rmP+0JGyD
m4QaXK3XC1NNmBqtbwFDo3ZfTr9WQjCXs3zURq50wYlWxeWzEVaFUOWtHiK+/TZPPHPITVYa247v
5gvTXYy0PzQIpLGikH4idrr4IcVmb4PlH+L5sHqw/pq7yB6n0eq7YiwcJ+5UKi++K9iO+awly1os
kvIwwMedyHsuGTl75MOBfmSu41Vu6OSFXeUngDqUhM9GXA4da+/1KxhkTIwZXfUS1HGZHOP2m/Xg
Q4eRFwgxehrPv/Uro8xHyTaHWTD/eWLcn+RrFyN680aVCJzw3xUFFpTaZXtwgZQK2l2bfxsdl/pM
5UBrzIqQn1CNUEaUVFX2gFa/Ak5+y3t3bAFj/4PEpw21cwGD7g==
`protect end_protected
