`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3488)
`protect data_block
jUFCkOR12oNg4P+eja87kkKRDLajApMsTNyLfk6FfZxu/pMwKFEfMTESq/BvinL7HY7vq9jCmFWY
ulvvFfsLPC+nJSxZ6dWEabmIQw4Bj29mFn2NRxRnohaRHKaEatiOEDoJUZV4VBuViSTUWfgmxZYZ
Pjeaz3FkdbDBuYzXp+WHBb3kM924ZSXGWl1K5AcbWsW4cGc1XxktHBzgQKZ3+Aay54xru3Ij0hu3
0dBzV1K5sJEDrjMCfJUt2wtBL5zXiR+8SMhSw3hWmrq9IfI7/3H38Mn6qHZmCY+H9hP01AN3Q+H/
cV4jPo4iyZmEiw/DL/BMbmAz3sEtrUN8r7zVatQGQn2XnvqPQFGQkRLeA1CUAe0Rw3LS+0m/iLnO
g6YhbIQZPJqFYSHA5YkmZjCWVRSJkpGVpKAFmavAXsg4usycrRXVESb/YgSYAw07VsKEVUDmU96u
N+jMlGPx6fCM25HIextyQL5eafyQSON3ucNpixeQbjoeO/PKJ2b8+EZUIEajvGmw7CTaNcwI3fOk
buYLnFgHtx3ERemQY8Mkd2ytnBQUtmTBpJbJWguLE/j0xBJE6n4llUHJZtW+dcBGabh3lmPiRvzz
vIOi1q5aqg+7nNMsnUvqWcw/Pnn8C/7jVo4llDN5RxMWo4yX6XQ6I77cXjkYOkRDPWNO1cNwUEB0
JnjCiZZcNx2HYFBDw3nU1cS2xFhgsH6Vy5xka0AhG0/dMjBakJaTQ7kA7NJu9hRJmhCtXL6VidPC
sjrkKwYzadGZeX1v+7yPN0cV5sabTkkJmT3zGPoY5ZhSjkLbuuA0xiFXD0fWxeCWKzwukZCff6Q1
QalF0IXd5VxatIyzUW2yKNgKtQWveaSBsWPP9OWqAwTjcpDS0SQvJSUmTWcU6gWbUHbHXT0bV4WR
Tb9429is3TtGndPhW/xDTSB0WvQE6xKn1YOWRNG5mmVHmaa5mrqKy6g3+dyEIFkOGXAuHM89158Q
TIgbHOXUa/9k5X0WQ70Ia+6tRAGwN4hDEEe4mlbkcB5wh44PiZaY9i5WkIUVL+l/9ZGNBsJaXTNg
F57ZKsWY+ifntwOz+WFBjGlszlGwIaWgl9/DpdZzfHctaTrGcAzbSGwUxehvBtNK40Tr/ESAQio6
c0l1pcZ0v3dG1gPNoT+7xAmg4l6dhDup0KBrWddCY2nBHlkGtoVNf42u9QEhtpBxxXu6kWQLYorf
yq6lHAsU2M0TG1q/XLWHSsR6NvzgQMKTM6XjMkihb+VAY3V01MDVMMZPvSDcWnlQApQegWMFio1M
TRMNGmEYQychQ8kMKHnC8K/WxiOz0+9JOdMeOAJrmMpro1ZNNjXGJIy1XfAgiZqkxh9ZdK8cfzyd
cW0n2HL1iSy1hq2VRQBquCKNNKXPsDEYulJOrbN4tqC/zn+fhHk9ZIXbPm12RPExF8FUMCogUaH2
XJcSBo07bgMGQ34CZ028wmrihZdTOY3QcPtZsGathBxbBbBtAGiaesVsXs1gKJCbynigMubFBQnU
b+GqB3PHpcqs1ynoTKSx4XDSoENOpjFaIZgIW6dfybxUr270ooBjjXQDg2zMip2ASYUGSHNt0efM
DPgbzvjx8n6kcgjM/va+EuUeWRKmdE9y2KXc4RmAionUvy0r49upaOMSuyGFvgVhG+ODykuKJe0E
H6pCLV6G0j0B5lYiEHF7FKrsLGgMLqVffxuP8JuOd8g1dVnb+5DhpPDrlw5Cm07iio6Qo1NHCYyD
AHlZpWFC38yhVs98sR55Oc4D4wJ1nN3ZPHWY3yqi2LAS5G66KrMAWwg4MrGxpn9mXkZPV4OFQ4bt
WF2p+6OxA+4Fb4k5+yelb+QqMe51q3BzhbDZqKg/bXAwVhdHNNsQAbmx3A66MMBrhdp9Q/Zcu+wD
pZ2z7J+kAdH9rCjtH+ct9ONhDDfNWxGLXn0AVYPtnODA11KAn6H3Ju+j5E2Qnv6H2/pJAmC657ek
M3cn5k6nfvVPd7CogDd11cPAkC5GyN1PiyXma/ERAk/s4CLylvUXGlZ7RcdgIgJTNWNzjTL7XiQJ
RDjDaCqum21ONV69su/FIsjUF3rDZRUesqdeVzigH93j5tu6iS44str3s+HFxDWxAFmA/BHS8DHe
+xYCqHJXX5CzYHbJQsMlAtAIO2OMgEdpZT+Qc0vWtXKVOKIn1Kje0+3wTtPGPpNcsGYn01K28v/J
DaCt/ZWiG9Yo3sbP0jS5WCywyqtZUjnG+MfceUbEJGF0ZZ+8eUqEGJ1Jd+Wa+v8MdkuE3x8A2ZV/
wZi69JIj8px1X1niEGIKynr840wUd3uV3Jhz6el1nnQGz19xXRFenA/XSyZ32fArXHtrMGft81yR
x6Z+q5YPCr7Os5osBgOIjGZy4fuuwaixKTbOcqDa+UG2LLRjol32Kr49Z4N14EN1OcpOOo2Bhkd+
IVAkE3XQylM1zVDPAtNoytww5H/VPraepl98Hcav4yNw8BjowYVnIP3VNDaQrJic7tf5crfT6Y/n
ukQnqNEtt7PHIryTIFCwMU7WRIrDQ1VasTM+OsZL1XpxBkY5cySSS1LMJlpnFvQD0WpHKAXezGLs
MB18sXAtE4+ltMdUqXZdqvazApmpnQOZzjUsG7A1DPvizmZDshm64GkbP5Mx4hpmESKojDkUjP58
mb7AszDYKaSKFx+/e99V9Xy47e2j8Z+WJOLEuXKuwzxiEpu/diNMkrQOyqBwKK6u8jYR88s+axI4
8Z6NMDpvFSd9IXMpOohXUX0BzJSX2Fq82T88MgBQWbyrIQO/FDt30noqLpt+8AG/G4fs3+8J8xCt
8TQDbXiTJ7zv8vdabOOzOSQCbeAzw0fZHzB12XHdkk8Q7LYzsGqSR7yR1CS9XGsmkRNbOUTu0xdx
K7eNH8xtB8nSvh0BEgOKfeXyUGHemHdSxwEqFSOzXHRitAoTWFc4hMFyU40UWK5jWpBS2c5/sU8b
LgXBDbUJX5T4t091UX1OeM22+OFoDBXpNDBrOeppfjJibgt/WdEcLVpggx4qceBygjmGoxi78PkT
iqbui5b1nseHIx5GY3p/5CSuTJ4RCw3cxiHwnGlRrgtf+oXKP69HZl/fEddAXHVyV9Hd+wKBtuJK
QB/hwCrCGgUz161mAUHMWOL3deSXMqpQ6kH/sNr9AfV5pxlf+3vFrvRMFPGkPYOcrLhMHr1WZKy7
4CnISXBuhBGEWHUh6IhKnu7oIkROSdihnC+yhJIEmR6CXfVf4e4JRZT6FDiO/w8onUM5dM4ZCFmp
GiZPbpnlaO/Za9Sel64ej95heWyrAugyUhsamfW9+UKTnJNPtQeJcgPUY3KwWs1pppynkTgMF05w
cACWMBwkh4Nl8FeUnubYAcnmxlRUkCWJ/SR1yUNyQR0J5Ir/9nkFtWKvecB6LfsrH6A44zJvJNCm
Nk0c8jL8UfA4x8Zh6zOJ0iO91WKbbLbY9zpzQScQV7J3tp0bNilA5qN5S+jjkyTahVIcxN7RNpw0
oeJVG5Kv0e4hAItkcqoi06QWmlW4sdc5rFcFYteMpo0TB2aPGmCL78PEMpWy1jyAGPoe75DpBBFP
dItHK4GHKhLrd7J6OM/zrC2kSF98H7MTUZBSkCO3+0qvT9P/0a5flf9cjYHrpBg8QkVElxBNEZD1
BB7q5ZNC4OE9IvnK2W0+7QG7RAyL91Lj9HIHo09Z2N2Jq+qojiqiTunocfMrOkKopVwMUZexp9BX
3V7yzZNOmmLga5+nU5Hn+wnG5PfisWyr3rMdrl8S2Ja9g1CPuUqLS6BL+2hpVKWrz2eJ6J/p82Sj
ZAJWvalULD3rX6IjWyEMeerCaWggVZ7eYq5/6iKEWmZPnFU8vTqqlGUwctdDwI0xrbT0jAgHApxd
QTnKrlQe6wy+3yttV0DNUh0GH160XKhCbICJmcrDqPM/dNO1xpwqfYS7sipe4oQi8pv3q/aFks+3
PbTfhMnrFpqW7OUyIPWYH+pDfY7nCIwpFHLPYN4QcZKWuI6LKaeim6Ep/TjNlGOis5R/qeqXIlyB
B9xQZKcbcJ4xFoKvNobi4gmYmfY4UWgC3Dwx2JKJhnNJnRVAYsQDNkAvT0k9wkmCueZ6iIks5oT9
4CNu+IMU6oFpILxpAcZuxx4ktVZms/CIh1eAd8l3Sqn1yigPXxvJRYF+AAPqlBbAlCENf8TstBOG
6OC6FJCI1B0gt7PW0PjOR6L0kkSWN4bLVUEWxuPUraLYfyyCsdpBYoi9NFO1JaQMIZ5hh8I66Mkj
JNjZup8sQ4K89BedaI1zS9Y+gMYplKyNvtEiaMDn9nmdfhlsCKSVOgPZji2XN6r+t2HzTVD/w4ci
Xp5nquhZN3lPJ6gWVYX3dTACpmM8hwfF0UdSzqIgF1ZelkuSh9xHCQO3+ex4lr+lQHEySVuoq+Ki
G3wG6ZrLV/UBkg/cXaPy7/vsC1JmT4R0bIjm6n1pncBxp/aSUyTHay6CRIh4cIKN1x3EUWadOEzg
G5VAXHEfJqCjkLsN/d0dGjopuxmMJeXEGvbc/cm3q/YI7hC4/E8VJGx0Wk8tRV1YnDb1M6O8NMOs
8vb0GWs/8P3ffo9UGYtITLHFURS9ZCS9UPA1wMkc/+EpFTEaRYDw6KwAIgH2kF8HlchEAecfmOKC
hrI8ELYSOaw3F2U=
`protect end_protected
