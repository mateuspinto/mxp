XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��(�?�?�G��)KM��3�i�����+CBr��Njv���13�A ՑK�A�:�i�-�j֋_j�&88���3 ��|� �ĖV��n�Z[��1p�\4z��I�߷f>+�O�=�[�|���[������o	��Q$ʁ���+8J���= 2uPf��m��=���G�q�"����f  ?�l��xK����-�8O�M��O�W�L��F�9 �E8v�]�V��B�aP�S�yz;m���]���f���r�=���`;߲�&Y�l�z�����<
Na�����R��~�1,�M����쾛P�[I���adT�w�a�\9�� ��:U��C�h��M�z>%S�n�����g��K�P�!ж�����<vy���7P��E�۵�m�]�	7,�ɴ��A�47�v�Q�OLL��6 �{&��Q��3[�ɿ��^����Ğ�daSO���d(p�~��e��V�q�2I��x�@�ϔ�.8vʫ�un�`�6�!^8ҌSE��e&ᑴ�P��~��v����0y<���=Ck%'����|(rtc��v�ұ�m������C�i�}T^
�bP,SPY��WE�t.���k{3���|�����/���[5�jO��-hEOO|����^Nը�8�����6ظ��n�����o,e3�V�u�)[��b��5��c�ֹ���� �`�y�������ab8۪i�(����-���¡��/�a���ko�K>�Y =��\W�tXlxVHYEB     400     190Q���R9�)k ����Ю�~�z�/��:�R��0C���g�O�7Ԉ*���E�fx����Q2�ؕ把�z8�%���U_����@&P�<5��M�c��YV��V$����ø	���0Ɠ�ؖ��!�	�͐�(t��]�V���5�0�T�������j|.�R��bY��8k��;�'�����E���_��?��AKh�V9` ?݉:�N27��F���<r�S�u���;����^�Qp=X��ۦ��ް�`�^��k
�kw'�Kf"t�r���%���v�t�g;��*X;�a�-��Rh��,5�k�i�Ð5����DK�x9Iq�reG��=�[�I���5����HKK�_�	���&v����Dd��Ȕ&���XlxVHYEB     400     140�hh�}�9s[ԝ�S-�"�E52��Vi(��f<R֗�L�\��y`����Y��q����q��퀷H�[���b�w|�Dkum�Ŕ%`��T��*\�:����O9���|�i&��Dmi�	4��3�r��	�j��˽�Ag�x�c�u�PK(+"ٕC����7N���}������"+�=2�	���߯#թ��f��ĥ"ge��(����`p���7~��!����N�ԉZG���"�<�5s��5�}ɒ��%sR�G	V���ȓ\ �4A>P�e�8K���Lud� ��{y�(�e-|ۻ1ZL�į�XlxVHYEB     400     130�[�Xgp�ܛ�iwqC�ܗ!z}D�J�X��m�d�6z��q��z���a�r�6}N�c�8�*7Y�DV��<.�o<J���A^$[�p�U	Xs���%��L���q�Vy&����D�󤋥�i���y����歮�
�ε~�$��sƑL��d6L:����4��F��[8v�o�����]�u?�[�ݪ����-f��U�	�̔��1�ˣ��MDؠ�M��g#Ҵ�:�ƥ��)8M�O�+�[� ����� �Ѣ���v����� �U�IA�tÚ	�pԨN|Ǆ\[�Q�w���	3yXlxVHYEB     232     110�g!�Ǎ���cD���ALK���1��)^�1��������N�n�TS����7���޽Pn�Ӕ{r/.��+F&�/!l-��g&��MS ���J��HH�KVnFX�xp�y���H�i#�>�}��"���b9�Tg��"OoU����Q�ޑ�����������k/���FR�ض8��5nխ��뾇 |{��V]�L�F�( 2�<E3�$��^Cb�����?���P�M\��{�h
�za���0�� j�d��a����X