XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����2���_���J��L�S�[���K�~n`��؃M�x��ا�c�4�4����O������#������T�.��^�L���h�JO8�\9!+�0�S�ܔ�:3�b=��s��;���jÄQDפ�|��::xk;���)�F+����$�l��h��	���z=/fKC�5�3�4S!0�	,���ǹb�*H��ۍd�d���}���-�'d; P�]I=��;���4��%v��-��0��t[�fN��O��h���#l<x �Z7Yij*[�
�*չ�H�Nl�v�s��F����?��A\�"jY�U�<��Z�T��Qv�E����@���FI��)�䙹�d������ܸ���n����j�]�4��+N�Jrc�D���(#@<&z�Ɂwަ�d�w%������qj=��CV�$M���Ҧp4�+��������Ƿ�.~�
�+B�=V4f>����2tG,B�I&�����.@Xj"�q�N���+�|Shz�/���Ѕ�N�Xg�>ys�xT&g׆W��+	��Ɠq��Q�kP0&�$J �.����q���:������*�B�:(����v�Is�܋�4c���Ȁ6��Ktس�
>�a����^����}�-()���~}C���tܪ.{}x��몡Xm���m�W���{��c_M z븋����Q=�'����9=�F�iz����4k�$P�m�\�J�)�`�: ڠr.<���>_$5�Q8�,C�;6?�͙[���L6%(�	S�XlxVHYEB     400     1b0\���� ��F�)SkK�iB観�_cQ�*�k�`z�o����hW���R�<^։�G�	��Y(ǳ��4�33��R!���12L% �A�w��'��V��� V H�oh:`@${��Q
ՄEj����v��4S������y%8DWKt�9��._��T P�f��kj%ǚFGg˚���2N}Rc$bM��j�V�}��v5@J�M7hY��C��������r�@���-�B:$�陴|~ҳ��wM
���-�p�"��8GU�p6��Q�ng�cA� ��u%�z�>����f�-�E��1��.4Kȫ|��yI�Cx�=�k��Ʒ�Z�l�BH��qxO��N��#<�#5�c�n�,SHH�����Q�	�07��#$]�Z�}\E��?�c���%�Ź��]Ԣ:"D$5i����/)R�7]^��XlxVHYEB     400     1b0|�O!6��x2��y�S���2̡}��V�Y8��?A��6�>v��F��ð����`��c�{�D�Y.noX�q.&ʋ�����bI��L�0��A}6Y������I>���y��}Ϸ�eV#vPF����,#��"�p�� �T���+'-��$��e%V�pB@�iwu~�!Y�P<�
8zy��F�r�>��v�`Ol�5>}N%v�e��w�����<��6I��ŵ�%�6:����ҔQ���y�_؜>�E�ĦR��߹�23�x|��M��Q+��1tS�2�iњ[Y._����i��7NF�b���C5�_)]�:0�|���c-�f�����lNѿ���e�hwb��8,x�cf�Ep{&M�����*1M��h�n.G�xgD��Pg�DM
��V��7�k���WI1����UEV��XlxVHYEB     400     130 B�Il��[.t`v�-�]�
����>]��G�^ȏ���e�FuP�"��*�54�oMC���&O��8�=�9���B�?��_��*�!���?EʼދL�6E�2���O�����lo�׾_L�a�7��@V/k�%�S@v�״�y��CU�����o�,-r5/�����FL���<5�7XP�UG��6�CNKV�ܙ�S4M�/���!�-�$����w}~ĴE������q8cft�	�R�Wê�����w*o���Ι��}��bP��b���`��4�-zN���uk�K�� �5��{rFF�͂XlxVHYEB     400     1900�����H?g4�GB�ðnc�`����W�8Wi2��Ȋ7�k��*����Fd�Q8�ф/^#K�:�k��w����N�8Ԑ?�H/y��L�v�XY�MBpl1 ���3�Zϰ['w5'8#�՚V�!�S��7ɫ����swVޕ1���$��'�n���ThZ�y�������p$iE��	º�G���˩���(;�lh�ǫ2'uIܺ�5`nS�Ϣ�k�)r� 2y �<;�7}'��b�Q�؜lP��V�Q�&�rһ6��#��V���#IA:��#��#�S�N�{��]�j��a�r��2�&�� �7��-����� Q�AdԘ�΅pc�ހ��.���A�ѩ�5�zw�N�E��Gϙu��,6�c�ԣ��9�����B�lh�&.�!\�<?��XlxVHYEB     400     160Ⱥy_��e�9L��pG��:|~��a�֙;c�׉��_���Y����Q��6���S���#�M��p�l�:��ټԥv�X��aF���S���[�<X ���Q��n(��׌sX�j+�F���G����5���G�s4� N�`vX3Pߗ����W�*3Ѫ�������$l���^Ɛۀ&$��J�).�Lt�9@��6��#�M<���Ң�B%2�	��o8z�Ƀ�B�!=�_��o@�p���ѰF3��D~�£�^�6������T������&�C�ig�۠:��o�M$�}�a0�kbB&6t�N|}<�q~v����һ����u����_�ꯞXlxVHYEB     400     1b0fI \��N�#�T�?�z���� ��x���9�  v7��*ԙ�����Z}e���/[����\�0*j���1J�^��谭R�J���1$ǚ?x��{z��i�&JL���`VSi�L]���Je�Y��V���N1ɦI0zv�������Di�ռ��3|e:1CC�9M�'׶�e8�e��'��q���1O�OeB�P�Ŷ���rVܯL����[�^�6x�A�� �^kW�MvY~�oL���v��w�.���<�T���s�{���9Rq��sX�As:݁�GM!��h�[Y�7$A��h=VQB�G�7g�p!�RUt�ڧ��JO�������ñb*�씦��u�E�����(�
#��`��t�[�5���[^��
�_N3�/ ǚ���J2!G15��l�R}TVǎ��0�-�.h_���XlxVHYEB     400     160�J�]�)"!���L`z"cV��6E�9�4Z��]�RS �������A�֖.a],��)_�[<C�Y^�;�{@k�Ĉ�v^n=�e��mT�ϋ6#�6,���9T�3�w�~;��X���4?;]3�E��;��� �+��E�U�7P�`ĩ�}BEp�����X�?y���B��b�j��dXDD�aԣ;ؽ5�4I���!�/�t� 0,�NJ���J�ԟ����y����c�q���rc�=���d���Cc%�b(����(���!M7#]vg�䅚8���SB'�34)R��fI�c�-�jj:��cq�h�z̶b�œ�� �LJF*�S���s�R[�ZM�ڸNЃ�;XlxVHYEB     400     120 ���t��F�ED㥗�a}�ǹjВ��\�/s�������_=�W����Ǵ��i���xO	:'���tCG���m�>1��|7�BV��FӐ=9"^6z0ۚ<<cƚ���X����>�m��Hw&~fԱc�V�\���թNr"BL�s����f6%�J��s���#%��Y������̶�O�`U0^P¶��ޗT�>�����Ǖ�XnՇU��y�չ����:b2�8M��,q6�b ����[{<S�H���Υ�g������EXlxVHYEB     400     190 xd��� ��3�����������T��Lis���/P=W6p�����yS��έ��h	���y����Ek�����Ke��P�]4�i��4��,�g� �x�t�"������T|Ã��^�|K�<�a	��1��R�zMBu�b&��1r"��[w���Dٜ��f5��S�����5O�}�dUU��W	�ANC��h�)Og�Ng�%�T��o�E¤�Y�v3��Y8ݸ�2���9�)Wڟ��sPusn�������!ͅf1����`9ϓ΀xU,Ã�|9��B��&o}�H����<�_RpeB+j�Ŷ28��'۽��6��O�ɹf��)���(���s{ǻ�q���g^�����N :����)�!n|�=o3���z��$�Lu,!e"�rI9XlxVHYEB     400     140r����UƉ߲�o�F��Đ��W#ÿ&�#�2�� �ލ>n�ڢu�Vt�Ś�	ps��CJ2P��8����s�8������ח� ��a���4'i\`a`��R}Fq���=����=D4x�fR�cV���D���%r�F�'5y;���L�ȧ2�m�u��f����*f�����������n������k�mʻi�q�M����WnSL,4�[)Q�vs���7��2�AXVF:v[��n�M�]jcA[2n��ҧaK��8�����|]��Y����p:`Ccn[f]��1*�D:��F�nc�XlxVHYEB     400     160y.a�ѵ��{�$pI%{7�@�Fxz���=�L�GpoJ�UU����M�e�(H^��/c�s��LT\�bl����{����vl	�w�"��õ3}D�
N׹;����?�����g=n�]�W$�`�g�py���˜�p������+����6_��|�%���;kO;���Y�A���8�5>�仰�����CnDyqF�2pj�^j�m�6��t��g�wS�u��Y
y����#8A�����a*��:ac	�h�@�+�Z�a��P�Ub����B��^��#M��FcuҬ�$���ڐ�<#ڇ�v>�)K!�Ð����h&�� >f�&��RG�FL?-:R��XlxVHYEB     21a     100&��פ�!W��SbY\[c������Cfl��}Il���	 	/�0�9��&Q0f9g��oA��{-~O�Ť�NL3�N�0ͧ1A� }�R@����G�8��-�-=��;���k
Sve,f��6z����@K��ˈX��@��$�z�v�ς;������'y;X*��yƔ@e�@}q��!�D��B�wA�VM�mA����c�o@�j���k��)ө3���%�_�ŧrv���j!��#^�ϳ�'�-�0�>[�"