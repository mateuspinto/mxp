`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
CMvlIrnwiurQTLrBi7pGvZOyzeq2DzA4cCL85pRrYs6CMkHwzhs4PB5m1Z7C8DulS0CtDih1LOjm
Iz4kap0fIL/DnRPuDZlAWgwZaCmh4L8SzQIwGONiRzBDv8tTTGofG/hpOnxrWiAzTJgU4fexfS7D
312ja+RNq6Va1ioUq1LHJ1dLz2KDMWOHW6Mk/m46tYx9nvyvOcGHyEChzSEy7pD2EpIBeYod7MFt
nSXJ7/m2yp5+Xz1hcw3WCJqf9ch0AYQQHwV2qR6VUAu7RQ9Vykk4x3Zt0a7LCiHOcY9qPizWGjin
9fOc5VL8SK/CH8e+krwdIDVlgdLr6abBR6PR3Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="GStfj0tY9ulZ9dYcu8aaDWh+6+5NXxBA5DgeHqkQP8k="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13504)
`protect data_block
4vefgYHDtl10k8c1GhrHPamXXNltZt40SeD96JKEXJ9KzEyRIGPmNtLNhZ6v6VzWWOSUqeLnYAYQ
cTfp76FyghTASKjoX+ZYoXo48UnPWqMRhCQGNK6T5GeddARgcLDRRKge8ByfcLvifOd8Oi+27Kx6
5PUjgLedWXZx8LQsRCS+mn6WSrTk9FZ6nf5o/BlKfv2xQTdUQWbk862iY4ZyjYfLEsOIR7K/ZnkR
eVvW1p3/CN60iTC/rtRvebhIXaLvs5vt4KPJmP+TWnRucDy612mCXnUbnFkz7mwwXYtLbZpvmQwC
wYXzXd/4OmnEWVeuSHVerAEidZpTTlU3qcfzzk6ADZCkRDqSQfmp37nb8YKja46UGJhv7ing4DKo
h1dFC8qtz15J7TTDfM4utzYCB6YC0P4pwASDuNmkTKSp7xH0APTk/gllz2ZkilMBP5qYIuIbwgGX
fks9fLswUU6jtjRQ4VpTqp+uEa8v7sA7F2loehBBr2VxjvEPhONNU+sHSPYrI4d4MuAqXD21s+6q
dd9wEDPKeV5s8fe3kTyVyuaZlRQtWgmNaZNOu2HztVF1j2ca4c//igDd+12sD4u6W9f/xqJ/G3sx
CL8t7Te4YE8JLmYv5/YB+n81dHFEX0DS5mpnzheND8GCiW+HO4mREIR7kDLRgt76Khy5Nz92SGfR
NtplvHHATztept3RvNiAmK1EpsfvwDmD0NYR4dou0vXGs7dqt5OkG9l3DsgtrTJjuvGJygickVCJ
SbsK8YOLYqaeF38nyLT1OO3IK3orgSlGlj7b3Dtx+Pbh3G6DRSalEU3C+nohSmRxnzD0pfvPYBgL
rRXqSMBtOYiINgXpoLk/Ifj1jnZa1hg2CCBG9ltSyl24bGc59/V6oTDeq0OMJM4HvE8thWeKP+LL
8NQT+tcr5VL0f+AhlV5wzxiO7s8lZ2CNN0qoykZ2mS3WeyNAtYj1IYUyA1rMAs68+//9s6VlkZgP
H5otDH7fSay6yfSVb2VV5bSyXU8nnnRPOQq8mnPnrSc/Oux24VIuO4eRGdPJ+ZlJ/a7nmUO762eh
jl4c000DDNiQ6z6HrPB3COvLyGbRy5GwWPu66Jm0Lj0uaSISUxhqMxEWYkfwg7xwEmj1IBoHxW2g
Kuj/W189kRvk1eS/tpWfy6RVdK9c9zG/hCg5xzz2zN6cTNNuHYip1EjE0JgQwjH0tv2Ivpb5tmUP
LqYrQol9gmKDwLFlZ+eklkYYECXVJbdMWxnZIUNu6bO/nM84zKD1jFaPwYH/SBqKHAKesa+Rt8X0
0p8bSarhI/vW0ve91QJrwSZHeDcsMzySb71LvqH3yO1ecqHbyxJUliMJOdQG8dEEchoRvdUTA9tv
uMRlbGH+GyubrNznXEaNtRK2PTy5ybr7+5/NNKasxFPYi0zlMIioNMa4RIRzQ1V3PIx8OH9oHEVW
jIgObcbNlY0sVnCFdB6kRKVfLCxeGCCWGZJcqrv39jje6L7XgdR4UZH9FEPx6xhxvo688PKp+ou3
ZqDGN5q+h5SdxPuCTZ3OAcIQ8+QibO8QyJGYt6KQl4A4bpBakurJnZl/ul4JA1l4N0ik/mvKzvcZ
phjvAfVvmyWXcU5UwZ/Mt/vJZ61D9tXPYklUA42FzUlfhRBRqbwBTWaOlablLpMkRWRuSkQEUZN/
BCTnqbTVLGQo8VYpVqzIA/3iUSsoasMVh9VHZrzkqwe1lPkUIm7VBfR2AmEdOkDO3K6YBvaU/h2q
jDgccMf0yxslm6pwu73LCN3+Srg+eDFXsbaaS4TnKnA+gSpfE2w0y6vPbtjfWGuGOc+ty6NUVJ53
MvS1Xe/Ib9qLpl/RtZogjhfZ0VXl3J98vj9z0IWgBAy1PWGGRN2RRBvRCzhu6N5rPu0j3+QL8iow
Mu6iVV7ECSagw3J7oX+kBY2/vtjWpq9nob2HGHgHsZioK6qp1Uo7KCP9y/8TzZ4vpX7vLZH6/3UP
GOF7qKMzcwL4SICjSLJmbL5fbQMoCxxkEny4BSS5ihZF1bj5zLp/zRmS9mnKM8tL0QCwuq6kpKeY
peg459fB1nt/wyzFu9K772MuUn2seazlxaozNUaYVtKKuL08A/qNmMRDehNkGRQX60a7VQOzMyS7
POHDMKkDXOHMZWhu9tzDzcgjt1ffzsvfzbnDBV6FcAvsK3xxyKSouMGDh9t+LBdVCxkFtjBZjLPQ
iYZs+o3Z7JvrSVlGZv5zFtul3y6OCHJtSARVxFvrRvGC9KySEJh54GuFFyHnmWt2gMVrA5y5YNtC
5O4UD/PRPUvuqzr9ctWeAraddn1FQQBZXX9OqSOQUMCjE3u1hrx9VpEHR4jyNHNBE/dbwzQyRA/y
7NrcDSmOhJTK1PPxIqGy9kEsZDe0974sJUnOB4TvSwI0SGmBYVGHSlwdF3BM9IZ73BgFZExKvBkO
S4KGohsqZB0eP+mZP5sQ4LkP5sPZLDpNjf/Z9fm1TCehxQU5b8G6RxBCfQ8AJHL9R5GvHOC1XaMI
Do9d1MSpuAKgSHP/gwunK9Y/k+zHu2l2iZfgzfHJQA5H7KFnK//qeIVPdhsdXHUgzr/h3LzwKfpH
c9D9uV4G6YeTFcN6pArRhEcAwN0EyQ8JCF91vnjJW3Ibmf7l3m1cH/z8+4e8RA3WbZ/5eoT1+n+y
rf/3hlaU5PvuRy7ujqZ7V09ggx5VXkvOOFHZh1591uPXQyro2S0vF+5ba2GSt70PgLbzhM74Dsyl
dzIffYLSAB7/QQJ45KswhsEe8aT3uD5adHkbkYSJDxDXC77ZGRRV9osxGbX5Q3XxTFrCzuQ6RsXb
gDuM7mMzS2E1Al7W999cS6ulh7KoNu+nr1uzlNx8KoT9ZUG7ItJFBTR7ALlIBLQ0uo25fjsRwRcE
3s/2r0CbY+E85TFv9miVYlsbTDIzS1b0mnQWx8d7s8bKVaF0K6Msiam0T6lirl1kjDxFL6IMTKMe
7Rf5H1504J6XkJhbThQeoofUg0ATWMnpW1XpJ4KL8CTEDSb2IKcS5ZlBjzlJA9Lx9CX3f2W56qpi
DwSWgZWDKHsPONIO+DHUa6ne5BPy5XuRjlkJAQUo+MPCKaC+yOUKkGLJsjbTWmYoRYryaqK+QM7a
hrMnrCVoWBaaK8ZLAevmkb+39kmlyS1fdGfsia2W5RBd8zp8M2rsxA12C0GRcEeU3TgyF1uZ9mFb
ilFxMcpG1FBHqQh4ZzvgJ2fo4u2zuYNrs8GbWqE94/SMhW4Doo5DSRR4gj8tUq+eyaDxofgFZKoR
ATudsqNRyldVIcGfmoOZssQjl7cHj9PpX230RaGR1Pc1hq8iFri4NNrPek/ecd93AU0JAyJrH2xc
bWJMNfyqQ+WYhe00FZpLBjIrcd2de/SiMwhFAwwaXZsUiMckmd52+O+TJzeR2V/AVo8hkhw4W8g5
TNUR7cEE+wwnSWt8ukSFyTV8CTW5kT8pf/FwPGeOTf0DZEVIb0Q3OS04H0LiA/Mmbgn6ZI8AxPQq
Du+ZTLi3uc5vvYL3OO1wi1a+vNDVbPFTxstTU5b4+znCAgtkbE/Wu6T1FfTq6ff477ojMc+Pt/qy
mHvfArJiCebrZeZjeH971a/D7O+TXZgVaG242LwOCTyX9xzQfIsRT5mkeLTqIr9xb82U7D+AYGvF
jiMsWH34oOlWSaQrIO/csJ78L0FcvRc5wg49ui5HiopK8JfAaAGTI9dGs+hNtfUSiGkFm9qbWQok
PZLAbbi0dX7A1S6UcvmScxTcEN9vFLeWfTf0RUJX9z4j8+JR4ZNhNIzZi9Ok5tW39l5iQf4uf3bX
ttX4NM1EpiLPbIKAED+utWmtMO8fNCa1jbc4Cki7XwDKyvpwtG29iyNrmd+84vgmaIvwbjFrEPXp
7WQK8byIQ4lwiPcBTVeU9rBveq0wDa6qDbLmh0thWjSmvOqzuXmsb3L4ruEMta60LqNUfTnVVeki
vdQG/kSnSOtowP2kxf6CPtkLaHEGmyJzBX7e5rxJe+XmhWNhKnY2z/u6DHMOEHu7MKN3Vqd7uEnO
xJQlLRgeFvL5Ky4UgESGEgYP2PY+hzvJKWDO9wKOoqjLcr4CaGDuJaBbFxN50bCb0UuEOiFE/9k5
WQiErwo0ebLESchp4b3X83WxtQpppGwFa19NCvfiyl+IrtdjHnho79xO6J0rn1BSiuPPF4dh8iPc
n4Nl0SFwD/UazZy+7bL2+k29gLMdmote9Z/qMZiaV/aLZ/qNmgUXjk1VKn/HwRlhbmcBF8WGlcNe
ou8+caO/JWiPPY/vystqiwNPGKto3m8YjMWhUthtd4hehH5z/J7TZKKd8g+VXJZTZMHag+v2D/mO
sb+JO1R4XcQD+CnBBKNsaBSAIfR43GUQrN4GaE3JFvWqzgsiXch13bl9IYTr/4RR5KQWqNdntE7m
HXG0i3P2RiG8cwO8ouAcIsqsQMc2n1MDnNidF3WItT75Aeh0bOTL3iX7U1hkCMYuCFWoneL4Uini
DoQ5MnBJ9Yyh3XBWNcTT9x7V4MYOIBM6imYsEMO5nvQsIrphS5i+1OjMzM768E+kG1mWVZ44pNFh
wPX5PiGhg1AYI0YtcHpQAL6wOf8+qLFISbhw3t5JksMgqyCjI+DkpP2y5HkyNt+hIqQbFdecsmYw
89rrVNazKtwncMycgP2TN/M/gaSI43zsvRSTKjLfRGKrE5qhGyDjWK4W1WlZIY4zwWHAzoCKR7Mc
cBkQyplQHw/EujS/ij4OqIMV6B0lge1Vi5UsWr7MaSdgdS5+vhVGEhibEB5UP2lwzBEnfa1AhKRz
M6BHorf7Rf/zSJKcyD82O/nA8M+HViZakIJl5nnEopA7q9B1dDOmV2zmk9ln71Uzk8lrp2aU5yiu
2SBoF0KLUqAuK7ZK+Xj3WKThk1V/nbkjXs9kiieyTHfADUNBg8rhR/KYIy+YGXDa3YJ1Q/s0N6pC
CD1umbtmZkIgiQ5NSED5fxOOK+PAI3xET9HTTmaZ34p0vUGmE4FtaAsf6zuxONmSLWPeVuYyepCH
XVWfZS9S1wl8f+2ROH3qbcvBl9ip0C5HoU+7Q2YrLt2WrZyYB0HO/O9RaZ0uaTBiTnn3hgRQnViq
Gh+1ArV4zjQnA2QTMRlQQ2O3iqypb6ZlFvaOpypnvffrq0bCc1TFePIBFQ1Ye6P7ic3GDzwpf40z
TxscYkCcB6woXUr8r6n4emuDlTi1JNd75A9son5/HsD2/3pEs5QvuHHYkILuW99IZ9fbHlIzetp6
/1jX3JAYRf7yEneXsYKZJI7hYaYKkq0q+ESOGRTZKD+2tLvM3C+Mp6SnHNTpD4h7F1i8hzJpxHHw
aKnQICh+/NlGtSAGa+gajueluHPeKK6PubZPAvS4b2CB2p/tIsu3Evb9WB7MdqfbuP7FjxKZVlXx
epwfPvW2BpnNSd6EINPODlMJu2fT6Bz55tg1YBfYsiFvrUIBl4EcvUbVx2IcPrxTZvmtKm6wmxdE
qXQZnh+QQKO8RrAksBGL4d6vphAH5dfZlq6pvHOUH48ZIBIdVqJ1/55GmBhI4QNQSTeJ5uDO0tfs
avxzMZGvqA5tYuANCL0eCESX96baWXmn5uqy1jVKq6EqrfTPBV4IumH78uGXlRq8MG3aQ6L5OzhM
yq0QQ7huSfCNZznl9JYvMA0bEoo/KI0tDPkyc4eCo5JjuaJMuwFitP+9o+GiAK3PCgpfR5DtRjmR
jlHXdzbET2Y/DVFB9WC1ftC5xW+JCtmO21zB1UUWUYrtUkn7T42OB1INBXwkxUeKTgoPGts4d+c5
V+TknIusgmu/6BkRg1hysar2EsXvVFYcSDIuUA4dV8zUkJ8u1+zQobwPEOTWahgLQXk2/MddMil0
1PEjHbdnopgHo/FYPSVTm8oEQwTzc9HAAMd7RkoNw8dtV7U9V3in2H8SlckC0Ile3Ubj99LBL2EW
q1MPQVvBMBXLSeqQeGARA5O4AgytkpUyJZgTndbWRqlYAWsRPoQJjPZ9cUYak9zKL0IwynWGlWlN
aOyXHXJSuflsBWLPQFWTClEnZcqBuuGGgKm7cIL0vqsULQ9Tn8JgZjGe15yTbInMTNUaa9LTtOtr
lzyPD3h2NzLmjy4Xz2zA2BvEJlfHoJ3iFK8lJzjwNB6MX1Ta94MKD5lu5uF+4Bok61zriWEOiKPf
6aGhCoZ6+kwI68fFlxVnJz+4+Y4L3yn8SRfMBzIyRj3tuMUr9FgCwJgRgF8Q382TcXA/fuoffAHe
l1yp4nZ36GqzpD0ZoX80pbDTwFaEx1wt0cQd368qzS5aWG2txksN2lwDUqygDUUWpRFCmo/bvQQ0
31ZFVXeAA4og6wabT2NwQChA7TqL+PzJJ+Ccyx/z3+UgXjqx1IV5Rb613iSqgdZLBq9+U+1gNAD9
pg0QtT/SGax6pGqP2QKdBx0+ATgrZs4w44H1VS4Ao/wj7wZaWN46k+4CKGlJXAoygpM4c9ZsMBZV
uPwEUo18g6GjT+2noTCSCKSqMP0GYLhq6uxMVJiNm6GrdYVnlnBqHMTXPqYoFnUrEUx36glR/eNq
grh4jmVJV657jM1E1RZIzcZFyJNKf1iaIUyInlbEhWEliPjTt4PGk4SYDnJnc+PHNBMw0pN++Hvk
MXNW7HSRXxpmAXJv8GfWZewgcpRZHHP1/AWIpf1MtURLDonlolpYnjk1BwnmVcDCxwqH3X1iWwbU
vr7IT645oE3VIuxv0qiRKOPXWC6101jTLqlcwG1MoGAU6jVGYSKo6fhfte33KiDYBBn6X6FsJJhN
OHO/6jNMY24+2sQeXvdOtDfkWlMxB44mYeFZ+Pnbon8ZOiYBF6BIo2HShlnXfmz1PS3s23AesvWM
P6pa/lnPD4CJQPXQYSsij4mvC+zAUDEKNgl6+SY/gSNq29JmNs+yt9+rvV2igqYfO+O/HYUPCbEC
Om7BD/HPXYwtNxUaVHNFLOt4cf19DKOQ6UlKFPZKGI/df67C5eHh1qM7JJ+pwlmOTsdokg+EJLOz
5QkXA7t1f5S2U0ikUDA9H81VOfT/5pnjikpUkuUuEmj2lkSnDMou9shf8JDS/JSSWB29R7xaQfit
RPC6zdxlEi0KPW4vQEfgKsF2J/ebYs5bsuAqemySJxJHiQWx0wVePz6lWYnsfX9WUTS7izX372Uq
+M49T1IrfchyxyWZNS8dC6NeoRmjtP1VinKciuKWrD3nuN8hl3O2rUK3BVR7BMOi0uppk7MJnsz5
zwwwIj3z/cfWaF28FicGbYLvhtnFa5vI4mbhE+82PgPF7dDqZ9o8bGM1K1t2K7U1WitCl0lr/Hvv
s4E7hCPu2s+bbI+tXGU9g7z3DttenTwq5VQCXPmV21iRzNWgo455KKRtNHRzGoiSTn6cXvWAhIxh
3dP4X3TDbzx8vWLtJRFbnyBT4oZ5VO2/6ZQOHL4ef7lYReid5p2VdTTRXF5cxwxxzUU65zJ/HNzf
tL6viZKF85ecsPyhgZZWOhXFQU1deb7IG9qITh9qTrewxD/NyYL+zOruwxIoUPGtiCEWGGS1BZc3
VE32KJ/dPovL4HCatRFhH2FqkE5/6Q7ojAVz5FMGP/whZtFIz+Gai6OfsXBNRKHrbn7g1QWm7Fmx
V1n4f6WPeAMchMmlNzm8GTVNcHQ/p1sxSook62R9nEoVlCYq9Zc+zu62JF+GFJ0k50gq8GB2McQI
YaKJjR5aln0GHTp7Zg7cRBGaVFCCqpxHZG/53kPLx3OBiDKu0KunQpSjPErnFq0pdXlE3fPNObnW
rqudMPvZE0paALfVZVIx2b0Z0hxmS4MX9LJSdrT0WWW6nCd+UPUp36WWGui3IWn29jbLw5C/UZbm
QGea+X2roGYXoYfHfgznZti/RESMtK+arc4QQTIW8NH0UIpZHgNZOfO71i9AEqh9pJoZOg+mcjP+
FEM+laMXm0yaBeqzjj4bWGjWFob6/WD+29XWaz8a6VTGYaoXfmBCOD7nDuH0ffpCDduXKyJiZaba
eDYpZ6wqu+kdAHfpbsKUsi5WtAThGlGB1mgKhrwDtVJ9PjKfSn95mQsMoUciDy6CQ3dmtPHS9Pf8
HgJ4Rf3lmwUctfJRfb0PpKvRgfZ7huqA0NMfSRCYuRGBuLBXFQBAwgGgID0EKRL/UYsjBh8XVwl0
UkPLnDmzBRW+DLbCvOEIU80hL/jTA5B3aq/bOuHHsSPf1xvHd37iZFO/XJl6X1BBd8P4rp3vez4l
OI6GN8qUpmHtAV1WfsIbGpYlkDVuUbS6buhatsRO3baLPOFajQ7M0gBu236nX3yr2TrtaHfZk02A
fmqeVyvbxrFtvD7A1ygR03dYpnIlDBIkuSvjsTtxFbkGrca5Ya8Q5kJD7Hq6B8OcF6C1kEnGPoKA
P9ltTiLWkwy6USLH9cT34vPqBxcD839aiG9Zj6kOyPPUs/iQkv8d60yZ198FMAk0bSo4raEr91vs
nlfj3oWiRqIVdLGzS3TYhrz0CL8xH5KiEWc+2mMx4tGu3D+fydzQvYtHuFY0fW6GveqmuKjDs9Af
xhfHM3iVvQBh3e4dm1xDJBU04tUoeKAWOFnRXF75zz/Ow8DEzU1j+KMDnrUk6N1rJwTSZ811Irwh
NQSpMOGnH5x2IQdsdyiaoGuDUhJRSvEL7lE3pLOdrSWMoV+k+RhdjnkVX0i5VtDcjvo6RS/yJpEt
+Bf/YK0ZZRYU7G1GBuaj5ZSvXEiwSzBYDRxS2ZWoGAQ1qMvrRSD8XZbBbsZGrE5xvwvmYFI0WXUg
Tcw9CTDJkA52cW+g62QNDNlK4jT90Fqc76KMnG1+Zlpw33PlTb0fza/aRvwAsDP9Z12oPZ6ZpkPy
dUpTjLH5pEmSGkxGOHQk7WG1oL0SvRgHU6ySKiRKSpRl+nvu3/KYyQEHUrXBY1rfshS8i0afSPOp
eOUdV/Gze8nqAu8A0Iwe0YvGGzYmn59/j7358cHsbDtBXILgqzw8OjqkZ3UX/mBVz1iCJXffNDLg
WoI+GTQZe1OAIoC0UoEU94tHPGPH/obM6M32/EIjFNJ7mpzwmJ20DAO8NlX+jeCWOHO3wM2z+x2g
hY0cSbLNYFG1WlvfRtghdC2M1JrZzBFf2MgHG97qgpQxSwerzydlS6II4jEhI+B0VKDc/3/Ltwbz
64Blth6nK3HzC0SuiKsq+7Da6dU2zMddG7oF8JIfuHEHqwP7vPJlmcPJahga5DcZ6hi5xH7EjvoF
hi+hCXC6F7wN+8H/L5D7xxPdbhxh73OC7cHYaAVNtLl6AocdD+YM5bkC/Ph6Vi1XdJw1AJfxRrO7
zLuxBSmh51BKtSTEk9ynVT5a6IlizyyX+XxUsdLon9uxwF0ttxLODdNTi5y434bduTJSab4LTRCu
NLpMtiz0RDe0P4uG3fYCbaVrby2fuBCzVpX8RG+bwTF0+qXP3ZD+GxlliPjaOMruDBEMamCf3g4m
H2lHfiAGjuG7dwMsEqDv+eWryCn2cI5Mr3fCNUgi6SoUSy0FLW+56NkCYx7yb268bxcapqRTpzBr
SSQf4MaQXkF/rf0d9MlRr3Z9GEq0mDhjZnAUYGytxAm7SUq1ibW8ykpvHckSbH9Q9byuGyNmC0I9
CrdyHWuKvtYoHLIbB3dB5fTUYoJi9mLIBzqTmTIk3ImcNSZn7q3kbT3myfwlN9RN8mba//6zc3I5
0iJnGtjfaM79FqWTZT0Hg3P2T5JlVq0QanIYB/51n1yQn3CCwA/imAfuJgc5ujqEO91NmoCuZpL8
TqHtEZcEp52C+QKZp3eQJx4La9w4Moj07W6KNMPOvTc0ORLrB448hfOXM++L7NGPy1h3IKjWejl0
zr8m5m0hSL6MNYz990vON2zqCoVZFhWCGYZVhG8lABjrJdAmawhrCxeX8amv7cQu48FCC0lNyTtd
dFlKrQUSW7ShZttDfqP6F+CFcqFzuiCU5HziH+NmdyROyHYb4Dr4jaEcJkhoQ792LWx8TwzEU1VW
X/ddk2dwoLkQmjyrsgyjP2K2pGotzeWKzDMPQ5nwEADYRZRH+2MtrZPEsZWe92EhKllEtTTQGv6e
WEBnOvRD6eRcKJp9PeRdcKPDXJ1STPe0CVDZNZs+QRJOMGLQ2MKXsPz+ynav279Ou/N0e084LDvh
3U8lxLyxtK0Y1p22C0WGGwjISlCiAbado8X75EZKXxIfdCfrhEnTYaqFNHoWZZBMaRuVANsrVKxH
Tpo6uszohopNZf+BPkxRxJsxuFhRXjMRTIosJRr3BT7+f1qjrLB0bPNiNyG4Q9e0XDMJd05IE4FR
5jHpzu7sx3wFWH6MuRqbDj92MAg0X7grXbvcNTTnObZaXjWd8kp1tT1jtRNIQYl74vQ8y5hVns1l
IZ9D3o7hWj8/UNeyASCRCeMeJFK57tHOxCKRsP7il2uMHeaRrzW2htrjy0Iaaf4gxshR2salpAWy
MYDj4asqnSx6kscY7k+JYWwLpDY6ksHBwMZRp8UoNDtf0SyyeI1UIslbgZeo7vlIrup93o2jqA3Z
8D4pGmd8xVHsD9u3w/RunYi8zkR5j9DXP1/9L9M64p1+Lw/r5aGeHETU0IjCD3h+wI0mb1tUfXYV
1WKXRgv3pT+wkC/xz4+nDd6k9idNL6qABqv0wPim94bzERGGcPVg+/ZtcY1nQznXhD6NLgw4Bdzy
HxJFoBCt/BHwwvTGiIGfCwBc3t7KN6C7V9+uBJM+4OjKCEyUioPdIkhdVW1mzGb43SEiOP1bQgru
UPfSIu9KDB4LaQ0UEVaYTSQAWYlLJ+wujKPG9/FbdB7RwjqEaYJCKoHrptabH1FiB9jEy1eZCpWv
I+9A+E/Nm44tqo/oyyEpHJqSx2zDabPFoimx6NjYj3eRmWww3iywCyqtYHjSJwsLdj/eyO5UD2q8
pQbP7669wkTgLc+ovTtUXh7S6Yw4MUIzDXKCeNkC/02sJywOcUrBEcitoSU2L5zbEz6LVViXwR44
aOQKZqWujxyL34nFgB810f1xh3r+/6Fnn61Onhez1lDNrjo9jb1J39jXFNEI3p5sztSiiFMjyqef
F4Y0bUzWK4QDCvs68DYZysXxDVgnM7hQH7aWVwngOyh2Z3LXs2ycVdyJZvNszEiZaZIdxBJtz4Eg
uxWJQnai4q0gvCW/T8gOlNyVOQaqfE+w4irL+4hUn8ArIFN6yBbXqhxMv3vDao+uji+ZSl1Z5jvr
wJmF3wZ9YyZXG344kAC4u8RGE0GpU/nTaJrcaAVoON9QoY1rNuqmlsAzetZ4DoNwL4kSth26WzP0
Nyll0TU3vSbCtfLKLg1JGXx4UwB6eJDiMt5S4aAIDM002R7QAonKhjiOf+stfMF0hfXbKzh15Zii
Vdg8NjNaq6t+8HUZtuHBqWLig0Y1mAoX6GWFt5p4dO+ZHKeCcpIVCie/zu/qF3sTaoluXAs+1aEm
xSST1FJbNxrCRTFbTtaSZKs7jrIIrgFizpITy5JMK1CH3XoGghwJ2EvGnRco8vCLEOCKE2XYr0Xd
vYphrO/pUu0DrzDl0Gcrpi2m9K8ICt/bfjWLpc/9IGMBzJ3EZAHbDxedt+eOV9z3HtHYLCOllwBu
c8ibYuAWkYL28pai8MfWiWXc1t3SXx/ecVg1rHG8ukT6cmi3jbXn7e4f7MFPfLXe0h4SfBC0n8Sc
MrnuYL4VYuzAEsgB0PqPuDPLZeAxZ0bB8k2GTEq8ZC+yt5U0jujUEMHjkWII+bMdKj0uSvAp3gFp
xD/mlDn3CpldtRe75gRPrYbTjyaqVvrnh9Sx5JIUGntpRpqloi6H4vyz7NH2hhHIMdz1cy+hvxE+
JXFae+L8azdXigmj57IHSEej4C3jr1UfalPqbfo5w3ahBg+lvLslr+C515pfgvFWe1tRIEcbPQSj
vqSbLfM3eLPD4mirv32is8dVfsbi22ix8/VmIBZFHJ0NtuMxLNc/M+YzCKwW5wEldroe5+ygue4t
mBZPdL1lEb7tPRs/5Pu7tSisdhmPphYkLbzlKtL9X7ihJZgKsUbnA477WXmDTJv454Sn8H/uGPcE
assn4bmdCqestqatabNtGAmP2jKwPul5rHLTGq7jEgEPZm06xlYHRMnc4STJzF6Lv4Zvnuk8YlAn
zJaFrwQkIlT+5yk5LVltngr2m0rSDuWzmNyo9DrX6eC+NBtM6keeq0kFqf0idh5KglYx6BctpFWt
JxZ+woDtMn1YT3wuzjuezkbeD5hlfQbqDS+SEPuNWaY8UCTc6bGa6/WIWAsIDCMbt3io8gPPnDBX
o4US7kfvLB9evEIlCwIRCwvWof99wAHp9Fy41PVN/h37UXUmbCsDtdd8jx6NMLEATjBfpTMaesNb
EM7tXTDcGv1LeNROXY3NOjEQggv7v2+QRsAqJBSs5aOBa8pAtrzof+wP472ptX9F8rEFK5HLA0Xs
G6KO+p2UH9sHFIm+A493J1Nb9aLLJ7WeN9iGyXxbNeygSTDKpqY6lp3Uc5CHVHHrRPe/ZIkHa8zW
XXNZfEgphTVczKMD3wa+1rWw4rEjR1vq6HTdIBSugRKQmlBky1RsNYM6rCU5C/2uMsWwGprqdNn2
VcFTDRI6pPf6ofz4OMMbhLEIn2b3heEzg9RTtH4VuCfjQwRSXyLpXjWcSSQOnQq3FPOQ4pbrnNhZ
56ubSTamhNl953JC4eCgXKCylT5TwBjz8oDmlcjfHgOPHhZbQpk4BXvLv1SSyscmHr9GuRV/d+Ja
WSgo4pMjL/zia/I3LUWUtb4o6HopIgR/xRGDsH2ZbRUrE7gkRfMPOyzUJ6liNRc5xnG8KCABisq+
X2IKrLFQglVlhLGi8zl+PgpWcUnZwV4kN/Y1KqLFJvK0WQRRDMj+J0AWnIpJFgELF5qpUS7lwuiz
kFm4N9oAokgvMmXpxDejUCJ+El8q3LVzQRmS28VlM6Y339kBhUibienWIlZYBVXbGxxiJfvJzOgL
diq74E6V/gqeI6lrwZddJZVybIZ8Mb5jz9JqUhYMRYWFxKcnRROSI3API3lylnmmpr+rmpwN1wS3
26diZbolenLm0KvVBHsYUkhD4v2vf7DwMm7vlXcZsj7KqAK3bq1f9HYei9FgPpJcWFYp04iAPbPL
J3geESoX8/17Ws2Xeg1JIHeCO827GKymc/J7bwx8iV/6ORgtpU5OxVeULMskHjpz5dV0pRjbdfQe
EwQLMq5IxWAgMxcwPcbxfO+AhDbgVNwgcCIPyZHrGn5chGpjzsa/+QOmosXsciJ4oxRmbqjxbYuw
g2jwYJRrcPHEqn780ubcVcgldTMcW9QNswuxhkOlB6pP7iFa37gMyjLQrO+V9h2XZgWvByj6lCl2
dIYfsmvP+tS5mGnW/uy2DnqrFqNb41c4L8KbdUCqKB2ml2rEjLSDIukq8dwMhnvXFiNW9vtPlGFm
5VI99Cn/ivE8WGMG7OUX7fm7Hc3b2xLu1fkt7UwhQbhxKRrPl79FqRkIqTHhjf7NIvFYeZVyDtGR
IGnen4q2jHCvquTiTinovODUbGicbZ9bZYsiQNRjxUPLzWR2diFEkP+OfMHFcxvKRqHEs6n4rWuw
OGvXqtf62HxPswl0KkQAxwNCh3hAwGd1NlOgWMor5q1JMRnTNovRUId1hYGBZ6aI8vR/R7C4+wBO
jzZFHETc5j8lj8jO0RCUIoPAU6BG9WM/akdkBj45It768LvCy494dkHiVHZZcoaU5WeNX0dR+Ebn
scoi6i5sJJ32aGs+Ynjo0k3+F85CR3zQjaQhfALpHdBywnT6WjSd/XECLHhSOWndiEeMMjH3pT8P
b7LQk39b3igD0bqcHyyKrcjRzkQDiHFTlG6HyzYm01h8YGzouSHZuXodNJnIBF9hDX/WNvN/v4Nn
5MwrKMiy/ZcR/PhA5k66DdsE2U0M3/go1JGtdic+OCR/384icHliMjjgG3sS6nV/KH6sIdiSp1c3
ckJqriGY+gJ8978Tqree8DcPbf9xEGEaPsURSxzPhtA7xVeWuegZ46M+dKD7PQra65vVAstrcQ5J
Ql6a2qfxdct3xI/4lRd2AwfBsT+bNHpWvc6cYaelAxOoR58Fc43U2pDj4RcVUX/JZZm6GjfyFpIK
XYMgSfNMlcY8PZyWTwUwYK9XlLE+0oBesu6W6gCT08fvXkQKBP3SA5Jbv6GneolRP17Y78f0YwlZ
5N3/qJDwxDV3orSi2IPV7lkGt9WfB3utQM4I8JFR6/1nqOYeiM28ox0WBpJhSuuCE9nxlicyTTiu
HnTWPz4dU00wG7libDqfCf7EnXHNiVCJtrhFtF4rZvQkDfa+zvPGDV22+4dWCj9pIRKGvf9ysCjj
RIjS5J3OqOKGjr7lap0B3AC0gjRjXLtKStlTjUCMuHIbskRENu6aT958Zt/koGseTiCcwxWo2Gqs
dkP8/I6Mnq16V27oC7xtyWnjEy6ZnULiA0cZiKwnT5p/wJMyw4nE6nXN0QVKLLcWVGfTRSa7ReMl
xoIwekrQr6L4TJE+/sCT3b4MkIVkIwBd1bfiYEYprLbldSyTPnybFc/AIHs70fZyxlLZMBaLXMmc
m+NZQ3kTvOSthue5hZfusqfckGUbgSUKdfoP8X/bwzAP3y8x8yeqmdtAddd0uwxcLyp495YucSDw
fBu5QYLHHM53wiKGxhotrh+7yBTsIkMd6mksJJC/BAtyCzp2ns3s3IkyFy4fV2gElWtwUjPYlJ5K
9TkboLbiyr5Rbcit0n7gWRYCtF+Ex7bIy9P/W9Eh/wGMl1m9xVLHWmklJgVVSs5idEqhycLTI+RH
M11F2rZrePuZT7zptZU/r6VLMK8ZAmq6axlstmtqnPVwg2ucV4Z0eZ+75YwFzpuRrgrjLyOsiq/D
mLm26Amq04V2RwRo6CjZRP3PgRmIxWt4Xx5uuME181KfR77GXTE9UeCDSEgV3c9NfbfSSV4+8+JV
/loBtWDOCPE6MnRdRAth5K4uakgUDqktRuev5PV4pSEObBKpYbgMrk1o0PFMFHgakagG8yBVJbx1
HPN/TT/tPBYSWBtxIUT8szanjJT3+Hi4gruVQ+EsVQyPJhRXWBq4su3t3PUSvmxenSGMCRA5PDY/
dVYuo0u+tiDi9D2Ve/vlmSAU4NHiLcj4F0NBcvCo4ZMsm+i4XS+OzKBTZo9t65nJxOLGXhCScOnY
5gyzGmrHYEwyLAFQwWD2kP6vFWpWn4vXkkhvc67FMssTvL2YwMwqBHiasidA+8PBvXwTwmGj+Yb0
DPg9X5wLxpcM4HJY94WMSxiRQPGTZ3g/xQhdtozNgt/eKEw8KWZleaaBIJLgJo1kc44t4tptqBcr
yC26eSnzsgfy22Sqdr7J2IYlt/yakcHkFtcLoV/MOaTgTZLOr8vS62dNad1jy3RTL3+M3I7AiKL0
Rsio0lorY+9iLQA1fQPWm5J7G98fKK9a5cyQ/cMGgSxrRG3hx4/c5dBJ1sI6G7F5+1zv7kFxY+Es
prj0YTOotfK9VkdHyY54aIlNMaElRL1f3G/5vTzTgItwdFVoeGfAQvrvEOPYX37IhcstNpluC2qe
IN4ksKOKZV/Ar3ex2ThLjVsrJfpteqcUIomREHVeqX7VpwO7y6R5b/C4Tnzisz6ATxZoDZ/WnIuN
pNU6ZZKTIdQA2Z2q9+mJ/PYsjzJYlB7T5Ogj2biUKwZ9yyki1kCqfTjA/hwqsV+zav3dVBZZiAyy
tZR00sez/RzGNtAOekkt7VJWEg/5d/Pvr/5xbMfbygs/ocTFSfKGq6IdCaer7QwZtIW/Tdo6h2b4
p3XeTJ1AzxWvA5RzlrJE8OZidcDYGttMSVOIN5uRZauVV3Jsy20TgJ4TdekKGQ8aWzyeXIuHnjvk
I3xt+xcYQQ6sNkF31PHaBDXVJVNp+rHGB7p5ivk/TBdRhH4+WyAqJw0q6juLnaM8hOMVfiKO1SJg
4whDWhoXse6NOcoTT5G0K0YhHo4eaZHUgT+WunteqRCdKxvCYW+Qm+BRoVMcG1bweNIqSgfrnXuS
ZGpIBvF07OnwS+2aiKnerTGgS8OZrQoktF1xA0BBAJpIvBDvxqbf23H5W3BosZ+rUcggXhK+2NPs
VtIruBq+A0otoNVUSF/9aCE7IFWz2I+Sw/zcNm27FKfNDlFpfp1vQ1gaUBojrRZH4PvOzNyqHQsB
jpmMuhms+wHlNAAKCPQxn6cFKUMo5wcmWz9aLqFIEy9z+UvjpSKHa20DlpwpZReRid9Ga8OrEqsA
Kc6uBWh3EkHXRWMxaGgLK8Y/gCOw+W6afLswSrTQ+CThJMPJZtV5vPE+VmdKtphamuBrLMuzpNeZ
ZMA2shF+3XW0KE9ncogpCw+MYNaqhDvhL6qGXnDFcm2E8NDwAHV2augD9sFa8yujoe2vnY1QJKDO
lfNIkceK3DUgfyBoXL16QEFZifIcYo/63wzgBdId2hnLgvpd0JRulQJ88klulE9SJeQv8WFK/58/
EcftpttCR98Lslqohb+Ef1Fx8Q9rtTm64rrNty1c3XCFvOn/6HBfSgJi0CxEzwpf8n1peqWmGy2C
Tgm0Sal748R91UpO+15TTGLKTQSlwuVuv438CzNlh7EIq352i6jBT7H4GzrycecoQr4ZYIK9K9G/
T2bsqY6Ct4YlTW17QgMFImAIyYE04uZyyrXBhzcSDsDsACeA217k+EOmqQDR2j6TnBgbprht2ECu
gGpiA+Bi7VsVTrdLb9AgNXx4ae8TUla7+qQ5UNz1N4ABf5ht9q6lb93kkEFZ1BJOrstsin0Tv0XS
b31ml6le9A7x8FSITnwm/WYI9l7Q0w37q5wctqSS2BKFG4sWltb7do1cWvw4Cmf7eb5M0GNJLs6H
qM9HDeXD0jEf6F28Ff8yB+vOJYhrtIS133pJq1w+NjoCy3BfRVYIp9fy7vEt9b6pYIYZTBJGwZUg
24UMvG1wRi8IWxKzWE7HXKnSmryy3xky57cutWsURGneQSb8wA3A2l8nM/Dw3gxdRoUMznfvalB1
hdjKbbd+t1YppK+5tQQz8HuKyCkjTerym3p6bTWfA/2k2dmXG31L/kOBKkuxecccDb/5Jri7Gh7Z
L0KPLgSiTgCdrvNY6z1fsp/AP0/9lhpbBikURZKI0LdNBFKPBEDbH2IP/wq1xLMyFC78sO1jac/a
feGS0pgi5Uo0xAGCjZrnWavOHDv4Tm6S4cfXN0ihyNkNH/Ni+2k/JsrIMoFvuYZqt77QCwKFaRjB
Quzd+086qaKrnAuitvf+diy2V7THgxxJRybbKirJAwxOait8/brmoFbQ2zvp2vqbuioVanqY+NQP
CAPGhz/bHDAFQWuyOG7RzBHIqGIugEuqB/1bXoagAwrQId5or7uB8fuB2AS14JR8R6qQJYBaIpo/
edeVyxUfRu9iwSaB6XWn0F9iW2qjcZYCGcsJr3eSLJoCY5e0I0B+2PAdGcqqJgRTY9rCLKUG434z
l1JCBEF0GZCuvDvhURWmL+VFxciVcWg1ErHxLfjNQeUFIN9dIZMTE+iNo/B1/LMCVlydjWdcuQY8
TpR1JJetKrzl133x+BnCyw69mgzBnLp1kKLNpPyLhHOnuXpRkqra3fOmJEKwPhGx8xbGkpAvhoA/
FGiTFP9BgGYOzOBBgSnmsMFOTkXhmgFKHYnTFCLikZqr09mfSW+frn2MB1q1V9rI6emfgBhiAyn1
8z+Pk/9z263icX1Y8Lc61Tm7r4QOUJZfd6sqjFJf/RBa+uEQFZhyCOjRkJybz8PcW2vFeuAFeltD
ylzg7YbSen3z94CO55gamP8EI6kC95jRCPaX/GXlQ0OlN2Hry/CFnSJRO93a/LcAIVuKic3wQGc8
su8RFZbRQWiYbHZd2QAX2dQEnOYDgg3OSLHfvSEO2clY8nqKbxsXx4jjcosSWVPYqCV5xoORW3Y5
+Xy9u6LhHlHWhLaXNOlxyLewS6HWJcWm6in3EedQJY0rdTwz/MpFlpUgc0UBHWFN4Oq7AX7pV7HH
6wXDATT5wgjiSUTeoBG9u0A8T8lNvt/BnBFMlPKdDKqK5XHlzLDsURMlj38U4ct9rCRIeQ==
`protect end_protected
