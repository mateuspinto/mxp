`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
Xzj7MrTjs8QKYV8xJsOnleI7fDhbyWtkGEqBYP4ZVLcCyWkOg9VTU8xx9UOQX1KbnN1K2cI6LyHD
dzX3P6DBGXLhU0jGAlpdD8a1C9gdPQy/hKMFy4sNCgrGLx0IC/YwF2gPvydsbY9DvkBTZNWN4+gd
XMSQ+gO6EZxdbO/EFCPneyz1pgKtLH8zW3khrrEdl1lioLHiWPJf1J8p1p2ScMLwPc8PvHNU9SLM
+NNpOrWelqk7QwGtcxUVI53KV3jOQUgbx0Jt2Cxgk0X4cQ1er3rtFCPYVcFozc/CDs5LAFrb7t81
xgwjMSZDDvXqVO5+fXfOIoNaNP9Q0uMj0Ffc3g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="DK4mUho0SfoX71gLKb8PU0LLoQUsAnTrCdRSxQeKzxg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12720)
`protect data_block
KMndyvohNOIlUXgKxAqW1onavVEcEN89HSI5ZMxtvwuwDLzV7NWJ58QVpa54wBEukJXf1GvTpVf+
w9Ah9vkDIOVScIwzKQBSe3AuVaBUxNGA2f/ghtgGIODc1nBiCqx7+0qzy4LyKpqBmlCBUC14Wxp8
7PbnYZlhf891CGIX/8DNHxIS0fs9meeFNWsBEoUrIBuaQynj149IWLyJyfTMwR0+3L9nmquWFhwf
CXtfjjtFOug6HzP0zIy3kdfJUv8v8ab85KmcJOkrp8TKnqhh2IUdqoW+hRakdBhsly2aSaLWPElr
9rRshlCRv2r0/vkxsaGH9HDtwgdJzwwgBStaknNH3JJHp2BQLPKUaDNA4+s6WPggAd8KRC9t9aId
gEYO5eEWo1E7XhiunAyQV/M0OvqJEiPU6c/8PPame/GsvTtKiUz3Tbh7J0HSkQbfm61WYMDYv9nV
hDXIiNmrIQnCKf+jY9ruAsYLPlWWwHyneTBEbq+mV0jVLSPgxAOhn2bOIwKKKztBuJA5VenmbiQF
yiWeuWfbHSRF8stkzKw9JaHjz2xPd5x8uxSQY+J0FzFSczIAcJ5hqkkKV8I3ln3NssZeYqOnyMDM
uSfzXJrtpkCJrXFjyovdhkq7Lb58hWYApdntASpFtgWn8/R19womtLC7Xsx2TuON2dLny21EgIkO
M4SZv+W1Mus2+5td75tlkZR5u66DAOv3WvFwTQFhZdF8Zkl9YIREDfW3wAOlve5EARFQ85rFDlVh
hziRnOnYSyO+emngFZFQGudrseGq5tT4s1vfnKR14xlyvAyvndrtHBReI3zSjAjGBDgciC5frMFb
53Z8Jw7Ncv7cWNogBJ0AJ3u45TgSKUKzaKi0Tt6YH3fLxtzeYfsmhESvelkS7h4W/jAsCrSB6jTW
vWFHgXAQZqabUV2m1npZGub02IFIF4Mdi/yvZpp3GXT60CtHA1einClcW+rapv7KMYfkcLiiR2x5
30oRYJNvT3VSXm+9qh93IfZzanLMstGIXpilHpJboTNRIrJCza8yLat6RCHbM390v6mqWDhhjiHw
uX2B2RArg/Lqrn5D0e8Ha3pnMXf43VmKkHts0G1ELh31P4CDdqxt7AdrYRBe2ENA1Dvo1BJYhDFF
lL/yhRijvUyfr8SIGZqK0gf0+LgjS8gcCFUK1ntyjYfAeMN/fDcYsafczEin59TBdYSi+nW6MRwj
mh8ujw8+a6e8s4lEVx8fcSiuAxPJlh6FD1zPE58zUVVbYWJBp0wwF2U0aAsmMLOQpNK9RUhH46dx
J6oFwoTW/ALBIjfqmgv57tT0KUfxEizM/TypB8qNvUP4uZy7rgo3G1em8l4OS1lMDv3G+qjfomAx
yCrOw8hsXBpqrHb+g4RvRg2RaIr29Kw1QaVrHbrfCYlePEcNgg9eB9MeSAVWeByWWM4q1fB72VFK
55UsBv0swVZG2Sf9MV1wmyeTvhJwUwZAN8cyqrzwxn30N25+uB91t/G4s3bIbyi+EFQHCmHMiBSV
RtNcGM4NvvJg5K59f5il5o82rt/s/rEqwJMJZ7MST8wrUUArRLtfhaf5e/EU33sKUEKlSTxaIWBy
1S7u6MvpfUGi72upDIYLM/KmMuy+Y6K/q0f491wBKEL6uNq4hlC9MGADpjAhzwtUhrnbUp9yoBn9
OpZb806TpsjjTs/Rg30FKFnLX7oeot1uSTbg5pM+s8Fx4K5kfexKbY3K9Z5gIaE/jz/zrznxCZKI
wkD8RWHTaOHJoBnTJ2mmTYZJLjjTs/ExwCX2wzb6A1uPeh4OxS2iHBDOFahNFfSAESQPaIiD+cVF
cFCRU3f7C+D6M7vtIcB8uJgELCmynbY+zqBOTpwNGBI5n9xdE89qOe6qwE60zhE51OWw52TXM2p/
T51t5BNldD5p6knHZNX/0/ydHQbpmARBAwerxh4WfS83L6ifrelxBaaH2CLCA9NcCUH1LWao/f1F
PHmM3aUO0/PPa6Z5GAdPyV4D9BxGT5hFQ3QeA4YRD0/v5uk6IKMnm009ZSoerDdtgvodbPVtyRif
LaXKNICBQ4jG2vuEkEkeCC7n5L2xjPFvtyFtIGxr4ChLN9nMPh5AQv+JEMsXSf3DQwpgfmJBJseZ
8R3pge7AO91nm8iHljpTLczVXClVxXFLajmw7enPn/SZajCJ04Ua+XxLha1xYyijN7w07hgX9Vm0
vV5FaJo7OevTH3RPtF1Sm7q5HIofXL31I/EiqWeq1jhJZKTSuPjnwCXadCo8ntoYKZOojKap0qt+
CrQG+VdVR2vb13wCXGD6AMH076UipSnrTOMlwW0eiroKLPUsJr3mCGGaPuotUpj2lK7zVzl//AwR
ZYcZPHalfafMq6ZXjNsLXYnA0oakPU0T76yzP/QxA3SHbB9QGlq2F53ak+bxBwP+H30GuIUYnCpM
XFvAnW0FDa4QgBcNotgegA0dk5RycjV/JWaAn/lNPYugbH+j3fEdPyzwGbHjdnsEPJ2jh7UvdVtv
XOA4v8v9fqFg+pbhocoko+FyNYtdrF34oP7D4mroz9jr9syDVzbjS0dRzrD8vm3z0PdyiMJWLXQm
RGw4ccbq2IXFuWUiNNF7/sLm5SaOu9twmjVpvvjC9n/6IMYKs+iFeX53bxKGZ4deViw3yU76hOkq
PW0DzTJrNMMR7k4wseJ2+TVdFChSrVwII7ax/KDgdE2TaGvlM9SmOY8VtQE475JbrilancluQxSA
O7w8N88XjpFRAIoTtfNd3IbAmzVkiCfDVFNvXaXD6h676IXXluKQqkiCFy7wp9mNKn3Zzz18oRrB
HWWw1RUo9f9OUfWf9ZL3o+mv+VAoLL+RcXpQecKUJ1ZcLeXaWZNIYh5FHMa1GiLvTo2vSHgcPUNQ
UZrzYO3uXoPD34JnnQSpxA53iDY8pQBrHfsgsj1UhGtPdYveX/qPywDlkIAhiDvtQujxeEPHEgUA
B/Mc4LFy6WEYDYbLPM6DlDiQTO/FVKf916GgRyHj+rbI79FyFyVhzrwFU+lJtYEnmUOc58SqZbG8
aQwzIwtQSJPzm6ZlB/sBDfN7Tfx3UT9O7LO2xVpBpSADXvrzTzKDGTpW9l+rIH1oUxLL5GLTxWdE
Hyrw1Xr6OfUmoLDpcQGDGYtWIj8+5pwbD99JYhxd9NDwdGzhYmZOJPkMGiXzlXEiOZGGdK94Nvk7
/75m231wnCuf5viwyGyLb8IP7LtM4AwIvuINU8lvJjsRbKVFoODVmxjt+d/Wv0tguZ6VYmtVkoi4
fnmlyIEDGDxxoRmToo5AYHNLG4aVvT4Id/pjUuH3V2oQxBp4vmnJGOJjcUPsRnDtEUHvDe/Nj4mB
wOzLlv14dYtIh5gs4M9NzBtCY7XyyeMUZvQZiMy3WFWXCeRuSgfObX7BUDyjED91RT1wMOltUHZ/
FcFJQv0mtkCgNzHjgbJ4k2zjydq6kIKKkCV8p+qFQOn9Y8hOZy/LGC5Qj4eSCrjPR+eYgEWbu85K
zGfV4Jkw1STKyr0Ev/O10qTOFU3PGowlWi6kTBNJiIX/baeumJbKUbTuWfuW4C2jPYeia6elsy9t
kZ77NHV2CnEeZWzsThYNyGX2DS+kW/YG4uAHbWySceOkGYroh9ICP3goSUWQns3upSxTxczPrSeC
HAy1dlBqLuukeb7Y4GBk26tAPgz+PxIUDQVqOkhBulTYNe1c1WICzEtuKZNWMYUCYEV11MsLVLsd
stdQg0XVWgNTW/hcwKR+i6cqtBzy+OGMjPqw7Ebz6Tla5NZKA8n6JlIcKbfANS6KsGc2AjGLBwtN
mUXuzdCir8as0SjkkqpVSB6GHPALpjnkTVAuPZ210EBHmoHZTVUPAZSw3y6IKenCBnPO3ca/fT+Q
vZGZRnsW920r5ATvzbUYrT/D4R/siuKM3mF7ozgop7/5K8lVrH3eK2HuqXSQWSYyK97wO2CbhE5L
M7Nnr8oYYoJaz/nEgioL2ksUM+SiYvro1BvRZsxKY9YzMbUqFzebhLdgP7x6Ox7ESbcT0WiIEL8W
M0C1ZrymEumxN3QIQ77OGzwvyVz7cyj5oIPn15Mgd6IfuzgByBzrnEqwZ2bcK5Lx6qf8Y3vdR/oz
wLpwZZDDSPqnXALz9KJMYa4QIGrDy7OgbilVfutHF/0ZXfF/tyA1qTRbZ/QmQKVBjVBnro6SvwpI
Uls0M7TuKK09YyImkzC2Ec0rk/8ZyErH3h6cqOzsNG2LsRgbyG1lAU3OO52TmXUK9cAuzP7ieLHG
H0dhn0wradkjj/m23JaoAUELclyzG/cmDDh431YdSThPzvMLnTg970hu1znz4MaeTQBO1d/VYUIv
LJ7vBSR1TLzouBNJrtexuAonzhMUiw5Bjuu6mBqIQImxpJybDaQzPvXnwOouU0rFPcmc2+7Lro8n
3rJlDYiBgyYbE9yedGF+ghPmM3LSonHiEmOciNWl8X1wzAw48wBsP7bbPPA8WL2SNKwoO8uqh+Lm
K8uFvn198hKwj+pmNNCqTUstykhBuSH85wEX1lfQNmOTBzNkDS7k7UlXv0QgSTbRSbFLwl/QXLZg
JKXM4CTzDAnw8albayflfBwRWn6kRJZlXsNQUcLAfWcVVPmYCC+d90stD1O2c9icLR5Dml6rrw9z
N0fm6hOgq8l8QyF0yY+PvTJvhelhq5E4DKTWvP2DpvbPpfVNwamqNYxs0rtHjq9b12K5UDi+/lDB
HZVOK3FGehL8+oMuhn/64MJmipCLlawBgbKV4P9ReH04+YFld+y3VsCw62mRXdwA4Cov8sBULiP1
6IQyaVALwO+rByU1WlixaWdJIEQLCO6GzYUr+7+C1WCCOG/AA23+VsS1hwRzpBJZ59jaAukj5/4z
dqYtiNIDJYwM6Xp5FEcDoVShsHoBxfpCidQmMxSvNAzFm33nx+OvwLtpPBzykbTiC4g0129m4fcU
DXofXuM7169RJJf/jG9PP1AlzrtvsW1RvuFH1Xql2rxekXLRbhpljT8UC0r9wacP82e29Grfx/lw
xF5DPABqe1Vm57Ab81J3mvM7Y/ZNziFHlqQS3Ado0qc9opXluT8QoioihoED8YxU+4UIOThYMQC9
pz/F9YMwn/HZRWl1gW1XpylIzFfW5K/hQwV3xQd7nXK7b+fBmOXiJe00JcBBJINzUIyZiZssXeI5
MEN1m1qPaWVUr0F+0l+sfp38ktIKpaGeFch9wKPstaiC+/DDH7uVDJ8NU0pteD6+7ZvDhq+SXDvK
qRyYzKqDaa7Y1+wPVw3pxkRJG95n1bQo0HIxVGkVcS3XPLVFnB6JNh0vi7hzRsi6nxzs1lRngnrO
mS96GFb4SYljIacC9JftIfRN/FXC6KLkk1nbJb9ZgqxDSzBYajOmp6fMBjxT19v77Q+j5vPQegXC
gfiYPWld2auJ+DigQvS/7jewyMpyiGTBUxAJKPPTrB4SfExKXbomJWnpx3MjffnfB4S4XunCP5dA
3hea2JbjZUVjarDEXrenc+epEK5gKKDClHWg3u7JwyHlnaNvJuO6xp+hwMFOL2foGTj7AcNneCq9
6EiReogvOpOac+qXvi5e8qb44NTCHLgz0HNIyF5Hk+YMvMLMcqdSm/6Fe+5SbEx8b6Ko+vCR3nbP
lxLOtGR7Mnb0lDAmht+xSAFgZW+sM8mbSTnI1pF4KihK7W2GaFqFdEJ7ECYSZqrS3KtViqO4sZJy
vlo1GRN9mnuD0ka5kFcCjV0NMJ9YDFHkEH/Fgfo6ZAooDps0QcODp9IeWoiavBMmj6d/eHkPXvhm
DSPbMcyfvmACuONdCayp45GQh1ffqZHHWfVA0ZhHr3DOsGsByZ3R193aj3rbO3IkdOdRPva6dwiJ
MeC9gMKcu/W88GkM7yTXF9T/ZU9UPilQcvM12LTz026p/4C/srB0DZQO3K8/J8mlHyRpK2i6cCos
HNPhSSL1uHoHJOTwLFh/tP1kMZXUfNeyCDTS6h7RCwl7e0lW6pahiioUqdC6pQtG+XqaQiaq+dOK
lMDuhaFWVyrgQ3pcSdOiQBuc2JCb8IXSsDUFstx+JWV2WE4K9lo5mF7H3Xx1tkrZC+gQ4J/6UtTc
zXreOD2twYYrHmyM8dJ9pzJ1B/lkL0D2HH/BS6D/Bp1xwBSbn4bmXxErElw00ur/iy11rmYUPXWE
uFYFKop18Hdpo4RClzkfkq8cJ8nn+6+TaXCbNfvbPm4lbRUMr92KNfmauzjwwXUpdK6EhElrGxo7
dJpyXx5rueEYCc+DwU2Y+bG/Cki3s4OktILEIViuThssEYWe9a/kOsjT4Muje4oiwL/3GnLj7lFe
BJJTOi3XBPP5FOapIpqaN0mjwDIXCSfokB2IYybDSPaORVp4VyxgG8QBdKeMPIX1qcjbr0vOqcLl
dTyK3VUR27xZRlpsxfmKOMLZlqHBHzu5a9nzaznmHslv3s9X8LVVKzDjc2656b3hMnz8dJYtgAiq
evPRVW8YyXmrsYTajAvfczH0K/rfFivWwQMI9lArvv1R4EPP9yVpj2D5NAg2IjbbGKBtToNmMWmv
SgOB4YROECg+Qj3IaNNowIXSG+aV88k7wO1m+uyRDEx+dDutxLu0C/iPHC1hdrHNQdeiO/o7posL
Oy5uGA8ar2tiXQr1cnBYEUM6QmemD66dXSfpxPzeTvvAQnqY0vjfsQO0ppMlpMw1SlBX5U8P35Gr
/qA3+PFcmpgw9yR4bXK9PekU48CIfOzOhqJQYigf26aCErjfyYvXrO/w5YnnPppdUY4W3/tusxqw
RE9widNdNbejt5BBfwQ4/DSQi7kiDceB0OjtN0KRQBIRzUoyJY/YUOR7drx9NjS+rdmdlGEZB0My
v3N4nHYa4INVXi1SCF0mQfJGcJOCS/n0YlTBsxPIdXJiyulZCHgnyCYwFtg7TrxVbQl5JrLpIczB
CALgjjXj9zzc63n9hwssnrOYOUMqvhHGladLV83K6y7TSHgirSmpFbUaY/TsomI9l/yIu1d0qK25
9mVO8MAWNwm6I2d53nFPm9UmXamnE1kEgOrP1N4rPrcf8Rk9sfA4rk/76K9svhmrVS0dZnEBX+Sa
FS4BYOexhMYSwDWNxYz9ZMe7qVMBLYV7PEpeNTn5YYYreK8Lrbltm4rhysVkzm/pNZ0crufcthFm
p3wjgjwHiF2HKwUhVvuXkkg4Xt+TE+EM32e8vnjtzh19zieoopLvUpNx1secA0f3KdkGCQnK3+xb
GsgzB2Wvmz9LM6uBJsWcA47E4V3alN81K96np/+pXr1CoP1RedE68AORA9I+xZ8jbwFVnjK8tAjo
iJ9hIfJRIqUmkM+lN17NL0EtujMAIkXEveYtcenf+nVLpK0hKsA4162pgPgMkFMs6Js1p0Oqy501
Kf9asqgTza3vjH1uP97UyiqFPF/fAx/jCZ3PCdDa7kqq8Fsz8bY7bfH/23nDAi66INO5vQLmshRH
vkoB0ihDmCYOqbTldW0iU1VzUPm1Inx418R8VMTx6JGWfmz668inMWkIapUhRAAd0bkYDM+ebGb1
BzDBjAVKMXp6Mccx/g6EfvnI2/UjGK22xPW6ye1sd67OWikTIWDQeJXdUsGi1mJNJe50wLJtX1tv
0SvFWq2SYqpN5fOwvWzWB9QTSFucbtW6rPEAW5kLDHu4zJVemITr46K8H1D1bv2OU8xRwVJbgFb3
L98okNaWWhBjOlZe+9Z+Uz1qB2h1+n2jUPFEjztYrzvl8yiJqjQ0b6bR7noILzdKTtSxRrjk3VNd
WaKPt7MxFHiU+Tq7gSUddjRcXKqI35d4E1tCsxAvkQTpZikHVt2PdHDxLbdgTleK/rWeRYkszhuZ
hrFa6TKndq+Ty2TUwYCt0jMQniu8UgWjl41hPWYkKWBDZBT4XMZA+hKV7KQz9+QZMYiRgVNWD5+p
HDyTdvTFuEOdJeiRjUHnGp+61HBs3w+OFVvdziZhx9Kcxq2iwbkbUPI3rZwUbKDVqN7i08ONjk5l
iGyHrc4cYHH9OM3LcaHZkh4Eg+3d0gIg+ISkRvc+FV1fUYWEd2WctsVLbmD7s4JNGxBAwEAO0xb9
ZOIEcfgp12nR22eWLZJeo4cLg6o8mOvWLiZtCUP529+UyvfrpPyTESBD0yryjqd1u2iewXjLlSK3
GNel0TbTtU29qQ7uPwiiVGKLAW39BUT2DJ9uPh77Zgock1Ha8HFnw5bJkDa235ZD27xZ4nNKCWwa
uD1FDgm7GIxPmR8Esrz8uDra+TDYxpQdYlkPqaka8gEfglNMu3cnkOjQbrH0DHzWYsnzlS1kfqM/
o67RjMuYQ7PmwYnzZZ3LgzxIogviYsxE1GJDUGsBEvtrioYIjo3mVBOc8CaOIqouVGDzxHjtpLl3
eGH2TAPk+w5ldcKqcm4SO5MsAj374hZAsETwCjPrN4ShcCt/WVgSObIFWzX4etJDXIihLu+tlXG+
FWhz21aDHlTMGqHDkLYWrD7JCtdOZuXigVZdnLq1AHZU6odyK1R/bZMaO1norEMaBKhQwzpHp5qE
fY2YKOouLOaLXgvr4I17m0FKjhup7r9k5NtjXQDxc33WGbzO5BVhXGguyCbdA1oOa++u3pzcHl/t
nmOskhBAVTXDaoqfEQF6GITkAB9Wse3RxxDKvuLCqcSXoA/Wyn7z8AAG1YNCItbtgxQwF/kbnX7F
HU5Zi9GAqhqg0mJFl9t/q7jBZiO2X2xSRkvem/tPQb3IFREw2EWHMFNWfNO6ACIwHeYxEgGtKA1X
3zFNtOCaUZSasQR5aPV7odhRwwbmfh/R1Jji6n+l0vdm31h+iYdCXulvUnfMZKDfNvmAPqAJSrz6
49cFVP4Z26BIEmscTlvARfMn9GgFG3RU4RM+ZQRTVnFi55ZkgRq0jzGsu4COD2uKauKgDNnTyMcs
0qJ9QLST8umHv83qt9p2GzqfScwDGhzCoJe9UCB7KV9lThiWSM+bkTsvQXPyzqhCV3GdLOHtYern
vbsDCkp6XMfP5mBz8NfSLd7ZHw4XL8BkDqMg6XdZ2f6uRblF7ZduwQ3ye+ghLJhnrq1pnPqMvCXs
8yiOqhi5diLOE+KFUTrUTUqtjY4ZB4Hwsn4AN4bS7FHYbVzIPlk8PE3Kh+oJfn+ULb/993BgnOmm
KHG/BhoexsiVscTPL1jRUwXeFR1C4bwY7o2GYpGl7x34zSmu6iUhZ+I0rWH49zff+ix9pQdSQHSm
SUbvyS56JoyJ7+4+Lnr3Cpvi5xIGiq0PsAvFCebSuVtFvfaZFguabW/ZJyu0qlvgF5zwXx5OP/yS
GjgnBEOH4MG0V4J/18HAt3mj+qjM/CUAqwGmj3FjDBe5CipqGdrv6SjHqcZaa8HKe8wlgAYE4eIc
dxpunxJgaXBONne24vmRoTmvjD7TljGsMlt2X5YiALgo2AlxcWx2ioobxStyjncPnsGVRJeBWyff
pMtEB3xsfkwSb33qyFtFtUfG4+wyxFa2nPSf8NIAkyScvu6z30WQ4UKl5WDtPhZ8XEmxaOhgDaxG
3K0FFotK86B00loldJVJJwIrFuVdTi5OYSbWKD/uRppnetgbaqQIS264C4QD8MV9u7+hOvI/BjOd
BwHVMSxz8QDJG/kcgCG6eKdr1S/0JEjp51evtyBxwWI/APqOxX/mohBQA0onlqFZiQv2DqlV9+33
lFjOYX9+Bz8aSGl9wqkimvbBWyBzNYEvypunu0Nl0hA+TH5YdNjmuqpZ27/C8EqmgFKoQbXwXW8O
TsSjQc5nKTmTrbxo/hh1YTHv+zYqZyTSlG3Mj8WQF3pwCMQJ0sojL3850A3QkTbk53vzxYNSdeuF
HY7KdJNVK5j25FZ8YMEMIQmmu/cfY28cMa4HDlVPpr3MrNMI0RBCi47eXGIVvXHaMNDCPv+h6NoM
k/CDYvCB88Jmgu+xb3PgAqyy4+aAk6yBicA9RKoSlayjk6D0UM4CrCANnDKUN86XCd6lsp+F9fcI
zwMXBazm9LWx7Q0xLyJ1v1bybtwMFHY8uTnI/CLEVj3PzKJcr4u+PcgAOfc30ew/4N0GnjcskA+3
AdeqFVDaL9FNfofuh+7L8rh5r3CcEgwzYpDQnwS8yMkdW25No1A95QTCmHIpjEfjjDaHahhlOrDg
Fz+S2c14pITFcury2yYXLKFTYnK04AM/w6Wy1Scy9rsuA6bV3CfYBA2rp6AEsGYk6WgRtP0p2lUL
RzzpWeQQVWLaBmGwCOY7cHnrAx84kESQrWWqxhCurZOX9BOl6xJgJY7K/F7zruwLQtf8Vhu9sUgH
FgR/ElW2T1g7I28N2iB3DYjktpNfrHdWt8yKrf+S1Eg3d8pFeyMG0/ZKSzsfubn+H0GWjVG4MXo3
Tme0IfOrIxC4BmAvJuz6zrwabP/N08erC6/QDDHwScfFS5kx5YWX0r9XBfVgzj7X9wDK1c4Cj1sn
2YSD8Ycbg9BSqjM9omKcHBZKoBkVKRWaYCbWc8qVU9u1I6sceFehCtE7eZ1ArYOvRD5suwBZVeo8
dvCcp3EdqYabr6BrkPOPASRZRe2OPfIfz7y3p8ipUzCdUR6v9lobt7tZlRRH2Dm/OWs+ydJmDPjc
xyfn297BOGrHodqlY+5n2If0CuGTJasyCHtaAbXM//hr8OKSXkDG6C02jc5V/E2IduXxTJKjnOhT
CE/Q9Mg26OtKXM5M1ufshkmxuKIjGFKE/GM1GymDvddm1H9iPV2RA5KxLQMrqBACR5RvuuC/mUtS
+ymIQySJO0gLqZLnvPMEm+fgQ3M0hTXtczpDrtZkDpnrbAC0vQNAdn+DY+elBcKAmyWUdmLu6Qq4
3rO/Puwys/biIeUH1eSbV3SXWIPidSGAPRB5Y5rgxyqo/Vf5eQX4otHw5a667o4e+i1CaTIdnC0k
8BGAmdBsAMzrTIh+4DlQkr6g0ge7tLy/jEjNqcd+EBU+N5ogZ3OC6ImGLf8/TjO2DFOcpV8U2rc0
3Z3NIBmCpdkdQLgX0NnbeD4FSwB3R1Q91+niEtMP/HoVDHukSzeBx/tVpE2xpTXVfCbfh3+2p1uI
f/oOewBJDbcDb5ymsskdJSXXC7rfSvZ0sifGTxAqNXl+fV03CONqNNNRbyOpsjw9rrZBuB81IcoC
JzbpO55yhdtAf314opNGz+i5sIAnSds9LmWeJ/wL0JlMnC6LxXjAz7FV3OqbwcMqifmuFvmYflYN
d3RCDAiye7F34ilYfyej6D+fOG0tDydg0Iq6pGzELsoPOpD9T+Ik1Iyhm8S8kZY9zF5OBfaeKluN
GKJb+YALKO+JhZyL/TI9Ct9ri+OBLSm2DH4JAR5/hp2ZOtrBhZfjDvQuWx8PFxFGrTY/DpSyPou+
hmwJ9H+OXQp6lsndaiAInxvrUPtHDjHeLUr+xOYNNvxge9dTmxp1fdwxM4fq8xFOuNLM85TBZJEW
7BaN6VceSII3w4zBR8fGSgG17qwheF5w/JRMJLXl/hw/K2RDFNTtlpVLxwTkjWFV4Y4wxAheGJEX
+CCxlznWOAdJ9R4/nRqQqOsBxjsnexQOLpmG0tm8qoHapu2YvafMWL+XOA2s4SYHxjmyaBt0moC0
eK1cKBAz4rMBqg6t0+Opi6l/KFWFkt0WEUuK416NrtTW4WxpeK638PiXGlgXaHSS+OCg6lJUmizd
Xkq1wPSjYNVJ+yPxgw8ZfSrVayazoNK+ISZErLJ9yKZvKvIV6mKkOt97A1CJ7J/lX3VGbiwXM+0l
FlASk9W/es8jJHGY3+ZNnZbxkNmLNPn7N1F7cJ3xwD3oNnruI+IkqT7qGLaToI/AKFgiYbgglJSd
7ItDSe27nuoiFoOD8uFbigr9N7X0tLQKnRRnwCtcd4qwXbUS7eJbxt38R8nOW5yG34T3yqWQ88TQ
cdwdpuv0ROeCxW8f3rs1iN4Fe2KPCAE7yfgcvM2jFTpu3KUV0DIpC3rq0bIk77mw6J9VVADuhllS
bM4TEnJthXgFzRKWoY/hvzwrrHSdbIg2L9jnwVtehJ//Zfz/mtGAC03tZ9mmzOV+I3C4iE7/gkBM
NiQnIohQBtMfPKkw/XukXEmzfPRrPbuMlsd6IAtc1Lz0cq73+FG5BRwF/ZshN8YkIrAj8HZamo86
lhWVfE0+WQDUyVVp8nfzzJfY7TO90NfXuOJ2ZI9zOgKu4tNf4aqOiFo7Tiawj5iAIYhkZWxsl9oK
/iCWzAqtZZCfADiZuYbCwME+l2XKniVumo8tYzYTjfTa/VfzxRxChc278p/ChwAetHOOLadM5cQ+
zm/IxHXz89sTHcaEZgpOn//As9EgP7dtPwLdiFjpaLy4lI8D4+OnXi3kGhAMb3XLS4xA6om6eIrK
UHWe1+zjngRXHA1UliDc2sOKNvcPN8ldm2amYEm5qcO9GtXjRKI0beP2S0AdviWMTz+AI8v+kdbC
lR5d//2SotBsI6AEcASuU1UVejKH1rXpNecS8c+Jtog9iVG9dD0ab/efAl0lwMcJnO+10eM6bZx5
aJoP/gzRrct61JQGG7KiyeveU354YkixlbACys+JjLfOzrkeWVX6FrKrEaxIXjzUUO5xIsIRiMbz
zzppOvIwA1yOHaOoLi3HdB2DDnOTW+SpxSeq9X+2NFJnflKePgq7bBQJ78o59J8OqsDZ+ecic5DF
psfc/F6GGwRVgTg/mEfLq5BdfOBdAFMNCnca5+6AEQooifKg3uXfCDImUaZ/q8stz+zdl4thUXtC
i1ywwXoBAg0NbA7Kji5BaO0UjX3ZafKNn3om7Av2n3yx5A3DJM8uzNQwFmMGE4zvaKJogHgtjjgH
+BXakS5E2OHPLMjTtRKjN2N/KmyBUHPc5mNeW17Yn3R7XvOb4HPYfwI1SGdFOgdGJrTDnJAqqpoq
ixFK7HZT9V8af5lrUBXLMfV5koGnj7WflL+YmoIV2KWTmXr6dC2YTgBxRkHqq5C9/77RAj2EsK+2
n79eAR+ydzKI916QoeGsgwmPNA7fqyf5vKbhgQWgz7UdU1WIQsBXQoR4aXXZSYQq2EY2kQwVd2Oi
l/cQ5UmE5soz93S1FKdEDWyMw+5GMJh5Oc7//uuvs3l9KLiMvzehQnOi1qltTguP2qJMAv3a1eZF
8Ta7PlPa6bnZgFuTH5oc7ONMCW9H3a/AXxmL5vD6Ar2CfL4UzFBTUbBfAyqzEHW5XUlMyrGQ4icZ
uJIsV8q2g/hMeRc8oNT0mwo1FfcaPWPH908JTh19Db7+Fk+CCfHaEH0zeQjBR+hExvykbuaJlZqR
Hf02+roA+Hnds87j4mWJ+cQRNLX9tLjxjTPvVDxhr0K44R6QKz3h48LHL9HwfGcSk49VNwwJfY6M
x90Musngc1nEW+VWSFrAAMs6CYTB2OZ/4oziW+w4CnV6FhbmAteMxyApOBlHbu+EbrWtyPrvaExO
E/moKXD+SHixBc7mllUJ2+m+7E7dZkmzlR+T+sTSr6SYgbupRO4KWy1OEA8ZzmkpynyJAm2ycx4F
ptEKpJzdAA4cY034X8vQiSqqme+oEhlD994G6ksFCBhBziQHu3EMkUxWT31w3m8MLUVFettVXdI7
/2U4QxWp7/YC6LqGdexDDS4TGxsv2ZPA1jJyVDZPelkVuaTqy2dcu3GnmfONtQuvrQ+D36EX4fk9
J0iGb+DTk3o5GCaquQYjKs0UvXXaOsDu8WrCUaqUAcbkPeEW5Sy4Xp2Abay7R7sR6cKJXfmtz2cp
GvWSpkinOfCinwqLCWkkWmQ19RUhf3Fiz8usOfv/7Z5JBbpMyIdr4pfQNEsyv7OaXCNQPUT8weOY
hOXBHgG0/dlp02tgoJJANb+HfKQj1nl8O+4plww5X/ZV498Bk4yfEcDl37fh56TzNUGfN4weWcLJ
p7t75VoTPNcssSQUdwJmrRx6nkOWHs4kbgZyc0iFx74T1O8UYfLeHRm33DU8tuaBL90bOXXXPdUx
1hQoYdpRL1qjsp6sdOBaEVvMp1ui8bYY3wrsntSNy6Rnwd4nGILPauO2B4IUr/Z9jbHWvuz0osHY
Aktb94d9wdsdlM8fW92tIIVy0S18RC1IMKQVGtcZtrez4WwD21LacXcN1fr/ARTUDMVQlsQfnF4g
sQuiiBu6x+qg4N9q7oUzGPjaU82QFUB1aVWAlSrX+Lp5bhuR2TPPfy9CE0naTFQyv3FXbFqwDhM2
3hkvk0vo0wNjjzAF+fEuHCO0oODqY77Gq7LXvvO5Xa0jRu7EntfFcJGhAVeHuI/Jq9N/RUOt+VUA
uqJgYqpJykbaVxh69S6BJERRYkovjP1cttj5sYouvTheXSvY5IMZ0fSlPYBctb1kfAZyUVy536zR
vKzQWTIcgusxMVe4IL5zZVZ0udZw/hC/42qwDXCJa4RS+gaZRkp8UngKLF6pZ4qou15spcB3DW9U
7BJhw2jflmMullBAH/f5++1Z6GTGXd5lVZtbpCU28ra/Hf2B1yJ0MNGuagbFlO8GDzcTUzn5D2OK
7YJqrAW9CZetFK9N5jVsj+6vscQBYUsv/uPFpnr4cKXD3x2FQbf8FQRVK/CRzTnigHUOfic0IYaG
nUHJnGmaLETkgYz3MDmBoS2GejH6LDI2Zlhc2sxuL0/Mq2OlVvmrTZLnHGje+ibqIyN/f+a3h5Qn
GA3XuY5zk7651Vy3QQndfRvv0lRNQUt3zfQWuIxs+N3bElfWYrhTfJm6E8QhIvxl+6Rp18M3ZvU0
BrqYu/7CFO5t6LVNuFBQeA6feyGgux6Jvq1v2Ax0VDoMGodgZKyod5bYLgEJJwKi0YID+6QMrVzw
M9OCFmCjYQznlT8NTQHsqvilgvhy0lRZI4CKlX1+pqALptArv2XJa98DcxjJY8w97F5k8T5riuyt
lG5SFV/jmDZvYu14WrmKZb6oL0eRc6YHMtYQMzxmC561BH65r4Tg+DCSxho06+C3t3QXai0C2ZkH
SbcvPyxGrXo2prhLxIUI6wYFvQ1ek3vcziufOLh0mWcRbUgqfDIvLkX6bodBOw78M2NX4ZYdbdC/
vBaU2jvNCJWHC8saV+hWe4FbLhwMcJjMPEFQVpjiUzxcFVHqtVd3jO6dmY5EU6w0xGzC8FCPV223
sVGQOaOtyhBWDsFiUBEkhUf6Nsvi9c+5R7pOW7w0RAE14VS5De4EPy8JMngjDKwrYx4wJxmXweJG
GtD+yzvNmBol5vY99PzjLFVkkd5FYeSEtYF5nwqIWpEkEN+frx29408oMqwwf3Q2EpYej+BKJa7c
OVeSCtQUuAoJgll/26xhxX7O/y2UhH1tR872cfvGFOm+lvR1rfNLWfnEBI0px8EaxEqxUGf+dXo1
EkfvAAj/vAkkODP4FYe2+lGEjvxJQROcOCmh6IkV8nWov3v/oLEiHk/A/Gwn8EGjRvGoIWoLbA26
byZpwCQLBKvvu29cKyLu1F1QJZRA25C6h/eR7UIaUe3lwFAM0hOrSyENMg8/ggoODGENw/C9G3/h
acfzdo5iohQu85xmF7VwYr/gNHoNvqM55fKHqiLFGMnTxCEbkjOl9FBn90/SU6HsaS7m1aGJrK+N
V2YfOzaso+J/hDR20sEDtDoIeRntNiytvgN6c9Xfg8Kx9TfmpixTVxmMte7nOwsfd1AskfsxYgrH
ateYLxBAmXpSMWirzYli61AbYkf6zAL4pFfFNQELR+aleADyXkb4/dB4kKs5JDSjfI/P1mViCw+Y
piEjPBrl6e3r0wjUvKrEl5vl2dAOssq5K1As8YP+XQ/1IL0whMnPZB7UxIBDneJm03snkNe3lsWE
w7Q1m8KQRvPLZavF1POWXZlW2TFMho59omQGzPXY/DIhR9/GJ/krGSKBCsu/KoUKVgkLv4Y1yK8E
JtSUIoAEEFsnF0TvpV3SwTT16xQjVpJlfjHrpgmPUQagCjnC0084ofJ6HPVlplpyfbgOQUS9KHau
aMVvXNRtmHGl6JHCbDEKbpxLq79VQUzdLcWuCFSiHQ44BUOIbYFF6kHAsmx8iKKDp+9lIGjw3Ynm
qeBM0tZXq2Emg8iUzslxTW5zKZk2iMM7Fye1GUZnXSWiPHzLAqyUG14XGZgUcC0Hg9TrGFVtRG3a
XC0sfNRV4RAp2bJjW9A53paXH2fuendMNllJ0FIiRn7PCiScrmw4maewdt6GuJOrQhkJwHONpCmQ
qjs5AXGhDVqM2Q/MBjfGn31odk9PfH4GKVnzeiK2pjbxkG8SHR2qGqA9FGmMbnbug5d/lKevC6Q6
xYvKKQdASmKzjjelzvjMItUY9LMYegMFvQouGCmKyHKg+5Qaq6Y5gDAYw207PusZhbqZBCYhMZLS
1DgEPyAzyB6GpuDKpNMpQx5VOdubk1GBQF39Z1QPAnUWXkeHtiDjDoDXgddUeQl13xqJ21W40weX
lSZJKwVfhi02wzt3yJ+s/t2DWIjmYzp05MXG2VON3eVg4WRujmQIakOHVr+wWLo1Bj28K9rOr42F
5R8ees58U4y/oFu36xoXCQlxiXhVeaq5k99TFPm2RMEJEYcWRQ4+b1rplq4+uNitI4D5seJGwCEE
I8lgu/aEWr30jwI7ODywcyxJWFg7J5opTarQhKSQzkRTZHvtvwwAa2+tTT+N10qjVrcYcZ3NRh7k
5VvVq1lHW/lj4I0TNmagN/guC+gpe/I5lMuYTzB7OOrU7CtoYLL1QSgk05ZERfQ/M6XYhK/YnSGh
ZifVV9EGzHDNrmHhySS+wyJrEuDf+C4hhjSa+if9/FRVTiub2inGZzUbEcxswx6d1uYeSDcYGPnQ
AhPH6z7pt3KefytikygsD29Wi/qj6jeYc4XN9DVaJo81Dkp0T9oM85kQhu+B+WtZ5updqFbWtCoo
hoWAJNGnhVKE+K2Lr+VfXs91AU4CrV3QLLBuNHZu48VpZCGLbykvB/W49VRG4L2T98Rdcg1uQeph
wiVybveZq4mMH7OUYmYFuTIcndlNt0JGvfyhedWpV1rzyLeJ3PcBfWWnvSLNtyzxjsxMMIPmnuHF
tHEcaMpXHJj2
`protect end_protected
