XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����O9W~���_��݂ġ�Ӹ�i2�|�4�Ʀ9�+���e�ώM6��E�!Z��D=>�KVk��ge�L�ia}Z���.��y�_��0J_OQb8<%��[\��	����T3!M�Pd�D�Kvp�\��{����3���IF?'{� d����v{�|U��N��2޶L����2�Ѣ���{��
�� 48jb� �r�#n#DuθN�L���7�|�"��tP��d��\[�$��g В��F��Ow:�AFȁ���5:_
�����H��Im<�V6M��$D��V�aH�IP����V�����%��7�]h����2�1�I��Z�3v�h�;�qK�*���̊��6��x�p6�\�tԙ�gC
[��f�.ƻp���B�V��#�C ��U�������X&@Q޴�˄�C=�
(V�<2(׭�ƈx5�����1@�ߧ>�i-��T2בx�hU��������cZ��G�!���4*��K
��{h��b���,�DYJ�>�#�ݜ�J�>�|Y�g�����t͚�>aU��B�";���\�L�B���l�j���_<���U��'U~6`���0ct��ʦ���k×i�_u��B�K{��G��#$^g�d+x�q�ʣo\Y���������~p$B�D���6*�'�y�W�&������n�s�����b����}8�#t��l���aa��E�|��#|L�lu���a��������V�1"�38L3��Vʩ��J��׏aXlxVHYEB     400     1d0V!&�쀲|6Ylmw��uJ�̓J�-)ř�AJ�m�a�h(�V?~|�5��k�0��a+a^��TSk�Q_��+h��G�;�ۣmfo���jt���^�F-Bs:�� ���@�ނ ��>n؍�9?'���%���29�9�����؍���O5켮K���޵%��m�[���s�m5V:U0�i�� \��d�ęQwq��*�[�D�zzd��<g`�{o~@�y:S9�;I�u���G��׊�O���}�*VQ����˴�v/]� |vhe,��믂x~2&�]�!�Ē�����{�]J�rS@亖���{���ua�dPp�%~���^]��2S�#�� S{�J�>�hV�Q�U�꜁����U&:��YO*�Xs
8@<�v6c��bv6u��=C"4�N{�=��\#�}�3[�k���7@�y��c�5sQ�ǣO�Df�llݫ�r��VXlxVHYEB     400     180#��2o�^�h@�-�wh�9�G�y�Z?�|�YvQ��.�g �ՒPr��:z)-?��͇�HZ�������Z)y��x�?��[�=Tw�θ�OUQ�����S��7������6��  q�|mJ7o#!D�c�ݴ����-O��u��PAv�Y����-	i �(ra��,�^��Mn<Y�F���^� �l�G����t�0Uu��^N�kBnG�UB��*���f�-ԟ̗�����ڰV���24�,�G���Ct��P�x¾��H�$�Ϋ\��&'C�K]ܡ�����	�/ڻP�g1z��}������"a�?{�ڽqX��x�2~/HMHT:Ɇ�!닇�W|�u�(tBC��+��K�XlxVHYEB     400     140
��HJ�������p��DA%}�m=f���<ЬeI����� ��;�M��@��R����+��n��~8� �ȵ��L'Z�֘p�U�<!N�y ��K��|:N���s�����[�����?���-�"�Lr�K��|F|Mb�����X$A��VT �=�$��'��@{��)�pO��pQ<N# f�͔Z��WzE���N��7C��ؚsg�p`+Kd�6U����*3��3~&���V�n�tR6�O��5�a��D�_D//J�W��1����!�%:�$���7 ��n�mqX�)7�����ao�XlxVHYEB     400     110�eȯ�8T�@���Xϓz�},��6��(�Q�M��W,�P>}�NH������p����w����kٳ6�ʌ8�˦cp+!���L-_:��XG�r�AXm���Ϫ2�?=��"=�U԰����n{.L$�v�<�σA���/�M���MT��<��V�Ә��0\,?�C������vu�^�_���]���_���p �fC@w��n��G������ p� ޞ�}7���e?W���L�,�p�'�O�{�Ǹ��81H(u�����XlxVHYEB     400     130�R������̢�?ᾣ��0܋�s|D"����x6��g�O�Y�sOS�q�xB����j=V�R��I�Qi��wn���O-�m������b��4���\^~]���d��y1�}N،d}�%!��'�@�� l�C��Bߩ��d�ŗ�?��{�oqRĔ�.��d�;��f�y�R��^z� ~�\����/gU��5	X�ɒ�S��g8l��F�'̴��d�vh�Ywyl��5��I��������=��4{�Ρl<�D%�m�*V=��8��I,��;	t���ڲfuXlxVHYEB     400     150d��$��v��cBa���]���`�V���7(ۿԕ��~��\�}����Y���חdn����˗m�0�;"З�����?�{�0�_�Ԡ�g�.[Z��ϱ��?!�P}IU�<%�/Y�%f"��%���Q��͓�t��ԟ�Cf՞U\"���o��DM�ӥ�}��fk=���HR�~u����+��{i3��79��[#��v�#�zw]�u���Ua$�ĵ�G��G]�<��ZK+ESo#�pD�)�'�������dH�h��;��;N<�.�v��'�0���#�%�3Z_�?v6�����a���5�ί����D����p�Ng�Ŝ�'�1�oXlxVHYEB     400     100�/��_���2+*��K������?�o�,B����f�N��Dx����%7O�M��$��M���sT�o��n��i����3T)Y�!�51xu��B���Q�J�����ĸ�������s������\e*"�����f@Du�`�K��'��?ۚ�˗�ięC�T��Y��42��,�WfO&j�Y�a[K��=�-��엹�B����;�� �nT��܉ٲ"�B�wb`�
��=÷؇�%rXlxVHYEB     400     1c0fF\��Ƅ���a(�������a�&�+��i�R�Y�g\��΁����X�~�%2[X��!Em"dZ�L�wY�f��ӊ��M��@Z���Ƣ�~ࢻ9kn�����$�P����o?	'��#����l)vK�qL��FO��gt��������T�[�	à������5�ͼ�w�?�(d��ǔ�P]�ܓ�?^�!(��tD�6JN 1]�U�� �Q�����Oܔ����_����c�K�?a<�ၘoH����9M)-�*fU��>���~�i�b� "1Geg���E(�R�D���=8�K����̳V��F��ʗ�S������� �Ë~z������~@��D�;:�`*"�kH_��խ���~�K�F��k�����z��ج�*=�)����si��xH��f��I.U-�O�PG�\0�p��P�D|�O����:qXlxVHYEB     400     140�Z��"w-�+ ĳLo��	�%I}��D��Q,�uv�P�7���UΏRrü�Z���`7������Aܷt��n��_Q��rl�S���\�Z���d�"������'6Ձ�4����џ+��@�y00��s�L�A�����ي�u�eNDG;o��3�^�������Mv�L)y��b��8B�H�9�K,P��;ƨ�S��y3~Y�[m���-R��@ɭ��j���ZM���
����d�@���UM����*�k�T:[V2�^��Z�x�L�oi#��$�%�g��_.Xˣ�J$m��Y��1�a]^f{����xz���YCXlxVHYEB     400     1a0ӱ��������.�˂*]�m���$V:,8s��Ǖ��/�~ob�k�e48���s>W4��j����ٜ�����n�xlܕ�C���?tٞ��/����K\�iV�c������V ���Y�=��2 ��Ɗ�:���� �>o�	_7Mٞ9�����r����i�5mN�Xm�l?$R�E_�]�x����C�!}:(m�w4���~/q:��#�ᐫi�K8��j�Z~!X�6l�aqw����<=䳫�zh�k��tO�
�~��� � T�"-$�rD�h�\�v>��W�[��f5^S������:��-��_5#��=�q1����a��jS�����NH�/8�h6�e;2����ƺE��� �=�T���\cK���8$���6���������U���{
�P�XlxVHYEB     400     190��`�c�*�����'Ey� �)��WE���B�:	�5��{�@"1���0�Z���+�Y��RhA���<�-�;���^3�솆�b]I�*߰Gx�R����9W��>�H���O�}�������΁1��[�
%��2�XZ��`ޕ�?�r���3dVU�MSN76KB!0�L�V�d��%�V�r��� {������,����l(^��������nzA�A���Nk+[4F��'����/��+�8S@t��H.z�������~*="�r?��r#F���H�����@�1zY�H�A��	>�W0�a�=ߋa�uZ9�J�%���s��O UP I��Vnp�H��m�$w �t؄�t��<�Q��������c���lXlxVHYEB     400     1f0�ϑ#�l2SR���5QD�(��@��A�YP-3HFvy�'\��o�U�|M�C5�~�4#w�9#n�Kql6[U-��x	_y`�yf�i�?�*�H�����ˡ�6tP�-����f֜8��q��w޷JHMl�㌀�=�\ڲ��?��b����,�ίllu�u�7�� B����1\�N�!���e����T�H��ؓ'9v�2'n��/sJ�cQ �Щ�j�FU��=��1˭߹\���͐gG_�*��oՀ_O����5�/��sH��%r��1���􍏄HJNϋ��͒�F��n�e���F�o/g�)��r�J�^i�V��
���E��`/Β�3����> ;Cak;<mh�����%�~B��%�o4wևXʉs;�U�v�[�We]�= ͚<��Y���]?��r~�� �j�����s�a��w���,��]�������r���Kt�����1�2��F�����r��
����*�N�VXlxVHYEB     400     170v������c�-,�^ �M{��&d�0�XL��DG��"���U���z/>�f��Y�kI��j�!��0�r�z���-���[�� ��H��)��t��spl&�&�ǣ����{����ܸىh��EG��~m�� 9�4�,�?�4�N��4��L�'�Q��b[!Y^(L{#~^�2��^����Q�l"3��y���Ɣ+�-�I��P� ��?�O"ݢ���Z�*� �#�@��3�,�P�
�n������oMU�`�� �vn'}xl���"%);uN�M�l]x��Z"tDU�>6�ڸ�(n �&���]�U��j.�\?�X&��d.?�1vL��/�с��X-vE(��Y���#XlxVHYEB     400     190�F-�*Wգ���G�9&i���^h}ܦ{�U�G5�`
�� �7�Ve�lO�sxց�#��Α���I���pi²z�j���Ȃ�rfJ����>�W����5zI��-[ჩs���Y��[+q�3'��y�\�����Pl4�O4�c�Nˎ>r��x�R�5��{�]Bk�AtK�*�F�9凜걇M�g&p����]4�j�M�_Ƽ�6.�<�C��,�yn(�:���ړ�m�Fq����\ �P�{w8��xu��U�ɼ�ur�ܭ��������:!�߰~Yg���=�}"���!�|q��RI���>�_�b@V�� ����}E&��əъ�q�đG��Q*R��"ץ�m!�i@������/�*hE��>�)���K�ydE��tX�~�� �XlxVHYEB     1fd      d0i�%���$#@i![�B��g��`�<�垫��3�W6�N��!B[�4�T���ʣ���iK)aOqBe�)X��T]��Q�&��#V���綈J��L�T#�m�~��R�tN����5$�$v� ��O=�#+V������)s"���/N�*'6⋣��
�����W�­��צ�c¿�+���FK�.ї�o���%f��o���Ӟi�Q%�u�