`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4384)
`protect data_block
0USWSUGxovGsyBJteYpEoZb542gXkWpt5GlWJKm80hs+qaoZKaGMnc05oRoIeBueZLndxMwKplHP
LWXPXLo86ogxg2ADifOhP8JvGr1KhebQhesyE4/XG4/wj7F9p7uPyLexvCvKu/gU2obtjkwvQ4WO
bdKuxtWLJInlni0MueCUl06Ns126aPnwwwJFwt2ECYt6SagK8gGLlVmBHe5fbfTvx3g8/tK+2mpn
tUCaNJQ1nibVckVpINYQVXn3/n47B1Skxlb7fMdXZ6R7E/UO0HhsbU1y0llqmwtT+HehOLwY9n8X
bBSHAebnl7Z2BmqVOZ6k0iL5WSehBtD+1ZSaD5vZExiP+YUiQYdAXPpSr/aGEhVoElPTRrVdBP9V
JRO7yePpf7PuBfTXcw/uoflbPiGQtqP5N5b0B5TFx5XoR0FFEfVEDufrhr5YFSTtrKrcNKyYubqP
hlIGo0M+iWgYQi5SH/7C20x1i+N9Gp6xuhnFSg/mzoypCTgySky1ZsRTQPTZ2QZkatXyglZbnjOv
YoiUdElWXXRE4/BK5ZStqeJRurYoy+3ylGvRfN/r7dXzDi7CcHSeYmYkJ3mMlPfImwPrgs0UOAA9
kaeSlumkb8QWh/hBotJ0ZTKZtqd6U/GDcalp8DpJ3X1YsmHPm3X4t7toaqOhR9vkKvtipvWdcNtu
DynlFLJk+wrNgV0jLiKRkPu0k5xQKezQNHs2WJiAZs4rezfaiiJd3TTqWgJ7y7mPzauM/a0u2nt3
qdsq5hPHYxoLv9UqOFNjHZ29JU28Lke+IN3eeKpKBc7sOcBrtF2wQ8c/oLw0F6QbLlMe87ZQ115d
O78pItJXAUIW4RhSkbbQCsP2zGPxLAsMZyYv0YlQ9QY6iQeKhNshRHY4qKKFp/xGXbpbPCVWIU20
8lwBFCYIAgBntxy50DPl4cbdfWbi+s+Nrtq8hD9755579T4Jflim8YCp+/U4aKqmkZxIR82BBKBP
dsPGs7TX1SArnuI5c2G0vIm6KVdlDgD22Oot8szLsA9l1HFmfbWfCBeevEeJT3OVUNbpDdWFe9e2
U2x9lhd9tx9bRRUCB+Bwt++6T1PY8VScei5MwWXQFqxKvi3HYg5rp0oxWScFnbRXQ632RZcLRv4i
7utkK1e2vhd2HzGjD9SnlB9zz0fV7q+hn2oSPFNI7pPUufHS7kWgA8imQh79uM3BPWGZ4cCLkmG+
YdphU+mDUPKzuA435S2IPAwoP9KgiPHyH69XoqqG65n+w1DWDDVYq6uenx7XiDbpJ7M0OtWDxAcp
2/eOMQU4AC1V6B5Q5rNtThn8qsU/YLQYfppOGpR4K6WUM2hN6EcEqRG1xLlmqId1htWYGmiz1+fm
gx7fEt3nPzzPT5o0yA2QHmLh1X5wrmuHDiZ+EJ3RXbAbAVaRm0kP+ifTpXSoukX8f8Oku4L5ZVnK
EcRpizS7PlC7wtz3IZ742caL3y9gIls/g4SEkQzeDAgnxMvNKvpeYKIUcCzNlhvoCGPqMzktf4Hj
fXEL1Ohb+jEtEw3K5Ngmmy8pHPdL4xC6VJdvjXBDCdD2p6hNOKtB9+uY+ZXdHMbl0D3ZxBizJB5C
o755kYF0UprLaNi50CGjYxq4bal8V9dYz/JTkYP2xuYYDAiQnmyoApQJf/jIdU0GJ2Pv7mQQMJRU
1oszNbwGe9EZCKfyqaiFF/9WkPV5KpjhElFx1jA/KnqVvwMGS0SsYet70yvL+xnz1n8vThwnL82Z
jw1PJ+JtAEVxH46wpZV2x440ebo3c0XrsIlwvp0K06DXqoLVdu8gsg21DY2H6GTW0VZ2LXG/hcJP
kagkhgmFzEHjSGJ7g/BzAWGq9fkyO0180DB8SiFZuSELgP1uxawGFJXyGJ9SY7ArAVWUQy9vH9xF
B/KhVWEPli+u+fCzzumS2N1o6rEdb3RqvqIyjfvFnKIXwj25n0IUZ9w8umTKzyHhK2INa7zm6Mgq
LfmU8G4ub9zT3bZBJdL8Q70Zo9l9I+tJaz4qNXGsa2VQvojhRLaqTQQmWu1Z2KAdkfyZyA7LNkMC
A+TNYOQ2WGczdePQtwMgsW2jJItW9Ia8u4guZrPyp0gaTu422VIsDmdWo5f7FlJao/jjLUG5IZk5
D1LwJMBg8YQ6FH6OgfDATgdAWLRaO9ftlB5Q0Fbuv6Aan+Ua+xnq6wOGYOttNyLBmVz56oKarAPx
nDJfK/C6cWTgh5vXtc537XzoG/YLHG65WKuK+mkA0ExRqipJmafxRD/1K3CfwtGD5n5t9TNanbKs
v50yhjfZ6ErM+tQBkU4462fIB+H5RHeT5RioUxAfuQg6OCvcD07CHkDeFfiK1oQKtMA3Bi4/Tonx
o+DSOyc4Uf/VmroFLlZAjK4JWVPfAxTnm2j73iE61CduhYoDVRgzO7u2CD1/U4BlahNo1pcXV7qj
rhnmSNYBkDzjcAnFRsqXNvKLEc5JN3Dk368cllUB41MZ+2sz29b7ZCilPLx7L3K3QsAgSDpnOR3n
PUV9Gv94usNw+zoKMrR3kmWwFw9Sy8LcTh559BKMvEXMVpyydiBlDFJhgWX+7f9SZNyOLYShjG1b
TWal+NG/4kq6yzXZbSysO4rdpJATIJX5T9tth7eFX6tEXcMl7Z1IGR0bsdfGsqDWcthuKeuF3d6z
GDVK83Kk+kVQHsSnl+IkXCwx0hRx9ZXPa4pGIjbhTaGFUYDj6yolTvfZwzWckdU6FqYI/ofyhxFs
/+jx2YbbYqgbxaUfoVrjrOl2yr0b79947N3UWrryrv1Eab1VNAds2huALdfakAmzPNWsmpKkH35Q
z+6E0QdvWX1D47ft9iuAJ07PohhX+ZJweqQNL6wTs/FZqiEN/iaU+UAuPLma3hINqtcDdcjMvDbZ
SndiqLJgVl7XaN0j2DfOuFsvhXvAf+W+Nv0Gc7kG9VC6GaJtg2r3PYUqG0yukI68GRDxvpIR2L+r
jIomQAHvqO7hL8YZPitKb91R3SK/2vdbdMhNErIRJtBe+Iei0b7rLND2bonkthXS6RREX3IpJS8W
34+sAnSzXgDVLQD5frH6kruBjyUndBhJkvf8DtjAZmVpfItZz+NLvAlZSB7JTRQrAFcU1A1iAzxf
/5iLakHQtgbdDWiPeR+9rDyfiAFiC6S/vGMafmIN1Z0dw5mJL5sJSDDZYBi3lyfR7MyRyYKgYIjQ
lBCEtQ+YOJiLXw2yXFjOE36vSQmTMvEE0S94iDdMTIgeqQYf025Y3O8cdmdZ604Y/H0m649cfAyZ
2gMGEZEk/5yQZ/fbc1r3+o42ad3AJetlg15QoGO4Ms3kTsidROSkqF/eLu0BWvBpwRGw1xn65K7S
++BeUh3IYm6Wjgp/3jcS/KjHXTT0SO1l80JFos/+UIpxtgRWnDFQghmSUBvBMHfHbrdMf4x5GAo3
q451ZgWT/Hrf23zLpZUvCMBGJMUPTowOAdbPAxpMHNviw7rjc2X8hZSwdimepJLVIiE02efjOHN2
5IpgJU444hAkDn2I/4ZRIMiPEzru0szqgYGZDYSI/61+WZcFUQyBjFgjpOJRC3d56mQo2Z4mchsT
pfdWLEo1Lv6DIhijh/jj9G2x5oqvOz9LKZv7O31zGqH9w8oo7Jevnri7m9MJu08kZm9czYKLTTqY
iNOpdgoWcLbbjFuuSfPwMV2njuAwnoQNAOumGj7xeeKQVWQTTSsrFfQgDRsLBgIC1MgLG5qNlJ1u
d16v+p5eTQKWg9YbuRnBS4Ev7e9PNziNMs98qVg7b8LWW59Uhzjo7Gm2MTFTpAOrVU6VFVkSULUQ
wl0wT2yGpgd5dyZiga/AY7PfIpaReBj8mIWJxjk20bomivJfZdooG9TtGwJHAQRjITIJq+jDYo4u
EEe5qCY7vffcBXtljmenTcdqHtlaoefx/zgWnCHL3uKwBZxylvJOekzMSV2A7hLblcV2vOFDMkAt
vrq5BNnlJjr3h/fYxyv+bF/0aharCfQ5hfxksPEjcL4HXB769DMMnTlseKNVOVUqCoAxwS7rATwY
4UkdfAjDgXAgNmINuGPmGNPjJ1WoyusbVKZ2mLvvxgJZTI2J+922tgdTAW6dxtCktnr5TvUbvioo
JOS1UZtVqvQvUiOK6BZP93HBakh7sqo1jgZLsYhS1PbZfglhjbG6nMHqT+FbAq2hAKrT2Iwzh0Jt
kDsYkll/TBvIhdQt9J61TQsry7b6nbCQX/2QH3lS8iBEvPEUdcDIHnJbsK9udKd3jS/aERXdKFQp
uEBGxC63xkdXvdHB49wEFBEFsDMER5mtbwSwwjvyHckxe8C2cPoMewilhLovWi69J3loz35P3PZD
fPEC75Q9NWcTBlp/YZ3q014S4rrSeH13pABS4U2oqSb3kYMJ8NbfHjmC+ZlRGscARtWNLMRQK1Ix
MQr9Ob3S7WGQvfjBlubHNf3K20ZxrXS3jsCS/lVYSZz7CvEQGCgjOk7ge/7p21+OPRlwyBZQX200
veRoaXI2Wf1l4UVQEOfNTz1gwZSkXpPT08yCfKT6V+7OwhA+K+EQK4OO4BFhFW4DOUXtGOWHrYZE
kjExPIPbmqSDqeNLLTMRpUaU+wMpbG0YZdtwzNRPMaF8LfWZ1JXCQ00K67AwUahtRMVN5S+AMLSq
GkxBob3cnwc9QXR/6KMpYBJOAsx1bQ+4ICCH5W1qCieRfr/FHi0YQjBTmoTcQtRIBAz8W5Z5ArTF
eVpzlW0/j9VJWYXz7jaO4qqKCqBft8/1cMrb/6+dnDZVV6aixh4XEF5BLi3rSBkTAgmuVf2s9etK
TuOH4Vp2ayWXaosZxjqaXLNTTWdZlhRJdov2PwrGBTXRgz73ceMy+BgHRG3/CNtVxwTIAQyvF1n9
QYqLWK/z3JUM9DK1dkB5m926DWZg29eAJoA+RZjXNek8xi91q+Qo+g6P9C1/nqw0sqN6IZnLdKOC
DHzTY4T7XbwICS4RBRqPTNmXZqS2PdA4SoZ1kEbi+tPBCfsw9b2pP1dgt1N7X5gje/3Ldk3ydkSH
8ouslvgWsJFIy0fYELnfwB316b7Q5ZcJRTzWf72a0wC28UBl6qTOJ7x79CBbumspfB5NIesZazUW
jNipGYOTIDzrcauwkZFtCDcKFRhn2b/JceNmK34EX4HJk5aA026tzuyA5Ac4VfTX6uD/HWS6cKfb
5wfNPCK0b+z0H3LCmf4RZGe46wUVJGp+jYzPYbpylfcfy7eZOBU0MjmpeTg2ICmYoI9yWDbG1/Fm
k6TGfLhkpqd+uv+u2UEZwtisdEVsqPa2CGjLzvLFe5mFUHk7f6bVg8/uCjBke5S7aA6fR+6XzI5J
TKqzaNt9TmneCVy1/spwLp2k+EwqA7GsXe7XUyWRuwLtbvG94wgEgq4PJdfirtKTONWXWUILPm+V
VJtFWG0qp/oi+/d3ZGSyC9MSZw56AFG+qACGmB83gHV9m8ijjFZiG9fqEchJLTvdnHp4L5G5TOfp
wY4PuC/fWpXC9I8qAWmJ1mknntOvX6Y7BBA01Ivuf6RQtKS7ycmcHblMtNIV7GN66RrMbf8lPssP
SWTkCyGYfCx1orhUPkPJrpY6l+Ru6hNBEU9uDUU96mS78n2oWTcaCm0Ur04HYHgovlmJU4Ri+uUd
HrwkL6+QrzLTxW3aWW57t4+Qbk7dUa4nThvIcKQPzj3Pfk21EiKXlImsJqNNeP6R1N3wr5Hugreb
c64q6hYkQizDXy8btB/6R6mPd0cQgjUsihV7CGBMjAErhzZoSI5WyvxG6OhD289LqXmra+JqhTSw
Sq6nsAa3+nJMwV/t/f4ds8S70J1iDi9nx8xRAYOJQfUXhooskjS7grBctW5X7Y9T10egiw==
`protect end_protected
