��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���!V�!��f�%��5EJ�Q� 5f��n�8�+o�)e�w�Y�@�{��Qo~�㌞���:!�~+$���"�Pu��5_*�0�#�F�g�=rk ��7A��PSL6�x�4+�����w&�9gl�����!��-0*ǷY����6U"�����[7��!kF�(q?��$����F�O���48�p1E^�j��ᮅT��Z
�ls'��S��k��i�+�Ǳ }W���CSW��$���ׄ�E[���Ơ�Z�����8�x���N���$xv��*�3 �`�+rT6�+p�!����%{���)�����N[
ݑ<_� Pqo8U��|�j��AQK��h�����A'�����g�_~Ukn� D��BC�/����e�"�DЁ]p���nf:6b��,J���K���X�L1�u����q���8|�����& 3���t+�S�c�l�V���2a���Ծ�;ս�E6��A�M�4[K_4/
��g� ��y���'��Q���D5�JbX�h��A�E}�ё�@8�-.�q��X��
�lX��1�g����t7� vO��5鳧�r�)%/	������u[L�|N4&�J� ����Z�5��@��QI`�$��p��_�M�N|��:ζQ�@��
̀'K��I��{�5,d�(��1��ԽU��wבrfZ̭_ᓊz��X1{���QyzZ�n�W��Ў��̐��v��WHP�HJ��Γ� ��*��PE�(Zy�b���)�5`��F`����I.S n��y#��y��G�00�˭��X_�(�,V)7'��K�9:4��mh^7��fc�Q��i��06ˌ0�A���|��kA��x�RJ�y��+B���M���]�-�JvC)���eA1;P`��b���);Wf��o@.�bз�S��C�޾g�Db'�#��9&�z3 ,D�d����
;a��+��]R����K��h��+����#�?_0'�握��PH��ͪ7����s,4�_qUD!��DP����:[�¡�ASc���sz�TB�4E�%|c �ڷY�T�-1�ӧ�̛�E �0�bP��T�@�\3,>Ox�3��X0:��@�[��ґ,	��Q��7�p#�%���K�`�����(�ˤ�T����#!�-��]�V��ik]����%��x;�-�Aۜ����;�<"�~|5�R��I����s^^�F!$:J�G�W��Sڮ���v�Mۣ1�x±��4""l� ǽ�"��l���3ja�=�-�SEz$D�|P-]tl蝄DL�o�\ΘtL>*�uȞ��,#&P�~��mK�8@MI���{d�<�y�!����,ĒYEu�]�t�	����X���Բ~|GJ��_���[���y�<N�Ƀ�b����e�����+�I�����~N,{Z�m���e��u�D��i��ޫ�pPyͯ����yߑKP`-��>@��a<8�|D�cF�qh���M�O�bG�������{�+LV� �`�6EtóMf�
�����@���7ҋހ�aVⰵA�x��a�%Y�e��j����=ćVo�.{-��L����F�L��'��0��o<N~����D�^��ε�a�^mK�\;А�3}���Z���R��D��c?�ԁ�F��3.-ÒG` ���%�1�=�͟�$
���ƺ�����BsKf#��̋�E4̼/Y^
�f��M���L|o��[�W6#�lBa#F�&�f�&+(�C��6�����U;T` l�NN�Ы��/ów8�; �uSi�)3G���Uǋ�`�v�������h/>˭(���m�M�F�g�d�\>�D�A�Bi�e���F��h؋�����4+�p*�t�ׯ�H��E��bd3��ty{c�@!���}��y<���]`Bլ4 0qe� t��.���$<Ʋ1�*un����fw7&�`+�I4"a�7&�� ��و��u���?f�-�qL[����ҵ�?��SDN7O�C��'���'������;�W��-T-�T��*R`���{j�ETY���A��)8��X��8'8s��=5vy�Myjz�,:�)D�����.�A@7yԍ)���Z!��a�����������P�^��m��?�0J���7�"M���'7��V�$��}��6$ߏ�AD�~|6`��j�AD��	9��AQ�ŸK���?�q�V&��\D��>�<���S�2:nſ����~˂dд����tn?éܟ"�6P�����#��18�i�.�����<cq( X����(�Ka�����"ĢIޚ��uh��]88Iըm0��2�3���(���h)�~��G�������Дv��y-C���Ls��X��G�pi�W��%��C��ul����Y����ݎ>����)]��)�-�"jН��KS��&����i]ؗ�/K�X0�ޕ�
����K񴇈e|鶐Ra��5������W���I!�|bb�ϸKz�U�xR����8�uq��1�t���lXy%�	�ĥj����9��%�_B {3S�T�Z�>�V��IsZ`����&
�si����'kl?2��[�S�>	�Ѯj��c4���[">�
~v@s���4�� ��2�V;�PZ1�7s:�v�x�L-ˠ]v�˞f�0T��n�����4�l����{,��WO<�d&n� GnI�]�zo��nY��0�@�����c�5�i}����聺nv��k��xSz���6њ�Q ��cf�ƟG� _H?*D�L�^By�|& w�׭��J�r^�z�{ɧr��p�9���b��GW�[�H���X��,��:8hxqi�0��!p��-Q�O)�ߔ��>�3���Zw��׺H% �?c�œ�v��L�Z�Д��
õ�9;��S�J���h\=�Vܼ�?F��
f�HMs�hѤ��ðL���k�`���ܥ�WJ�} L���G��VfJ<�̍$� ��Օ��k�h���W%'�f���<l(l�;{V!qB�Jߗ��q"�J��N��)�~�M��㾩h�I(,r��؏�%*ބ�YYA��}� ��&G��5�r]G�M�qS���J=i�F��<�:�(nH�|N7����\3`)Vv4�:�(%��kWY@#��|�*�K�r��7���H�#��S��*�Ep%���:�B�K�XF�=65�.�~����i�e��n>��p��z˻��!���2�ƉՕ�Pԝ�8�S�7��%յ�T��Ģխj_D��y8:R�=��9�!R:���D�C��J�o${$b�AA�3���J
Y�i^Ӯ�̤c��#�8bݶ�8���=�������3���J0	�9#�?�=$��~�249����X�'w��u�B�E�f2yr�~#{�i󚫧+:�T��u'�A���a�>0M��?�.�� ?"NK�wz�#�����H]���#����4!f"�J��?ЇR,�>(b�ǋk̈���lB>�O��^4����M&��$��Q�,G�R�w'�x�F.���|�ַJ�n�0ǪlY}3�A��"g�	��nt�gC�g81���\4-)�(|u��J/�s7K���nd�r'f����]4:��V�J5V��2y��,w?�1��@���M�-��] ��@�M������/"#o�I�[�!O�'2����[l �GD����>���Jw��Ug9X#��o�Ӛ�4�u,�;x%�n�����X����v�܆��0��{�N��=��ː���������C1֠7��/+*|�c��7^]���+E����#�i�ƫZvh� �@��4���-b ���!�ۭ��4ؓ�9[�/�� L̆bq0��w�MjB�3+2I�3�x��8�F��<���:U�`�U�k�)�TT��ݢ�1^l5 r�E�M����\�JCU
��=��re���xH���Ҥ��+���	�,dw
��o:�ϝƫ�s��T�8[� ����� ��^v�2�> ��#d�o�q�1��q^N$����>M�Tu�j���-�r�1$�9ak+�K��&�LƏb�J$�[iO��/)�|7�/*��q����X�f�x���Ħ�;M�^�ݗmR�����3l�����D��x��E����m^Ћgvx1'���?���`�E�&(Z��ϕ=��$+Ƨ�E�Z�k���B�K��CbD�%�}El��Z#֥K;�eإka[�&�O�QbY�������X�;�PʨT��c�At
ܯ��4�dg�{9=N�Z����7]BR������y��b�<��(�w�����:K�A�N5v/��ꇚH��ԃF��I��a^eaXV��ؚ�F2C��d�����UA�q'2*;l3�C6u�R ���H}$�(~!x��6��6\ �����&X��X�&<cZ-�
n ��oN�Oo������.{�#qz{�L-��eN��K���>S��C�.�<�#�'7�G1Z��^8���>�(�K�o�JP���+�2�%0i�ng=�&��߳KG2NN&ܟ���.�B�e�"�B �#�IPn�Yc��O�+���{�W�wYgnO]�!&�wy���ﺺ ���:���a�2�(	��)ss�cp�cY��C�����p	��{�<���ٲP q%�w۞ YCn����I5������ �������Fl�w�y0	�2 ^�o�Xˮ���Ի|[gY������Iq�ґ�eY�d�q�U�OE&�ƶ �KT��3w�l��*��*��ݜ�(��w �X�V�Y6����Y���Ӌ�+��y4E�$ܖ�C�f@
�H����~�ifƵ'�J�����?�/[�����x���3��Ƌ� ����uԎzf&�Ҡ)��y>�D�c���ƳU�>beKX��/�,p|`���d];��8GԬ~�5���.�m����mM�p4��/�]�����$N^�͝fXP-1W�,�|U�;}��Hly�3	5i�o
%ODf��U�czu�ߦ�F����ZCn!��Ʈ�TJ:Ċ��A-E�:P��@~O	�f݊sڇ\���LX1���:��3�j_�]���$v�5,̹;�c�G�~��8f�5�@���Us�x��J��A�/8'!_+޿|�"W�ڊ�O\�j�t�ؠ��� �Y;踽P���}r��A[l���6,|CZ��o�d��"���9��b�"vò�c�ݝ��#?�*��P��z�A��La�(|�^�e�S��w"녺��~��x.X�.(8n��*Qƅ��
6��dytL��C�p�S�j�,O@O�D�Hyu���h5GjHM�!�u���ߒBi�C��ֺu���nd�����1��U�bwd,������.��$;�����nB��f�N���Za�E@'���r.ڊ�8�z�(��a����v�H���y�ݻ_j���t��:�+M��G��UL����Aln�HP�鬄�<�p��lX�C�zY
@�,a��.#t��p,i�P��!����i�Kˑ��Ii���I`r�4��l�S�}_��y����w�xw�@V毖z�X�c6��9��i�6"�0��L�Q�|������{��p��d�����=K����� 4@�3�h�9����؀�/��?_x��L���kl(���a��҈,�N27�߲�%M���\�X�Z�x
�B�#�rت�o�P)��[ Z��vyl��N �q:J����sU��}4��&#EA!7P�t�F�JCl2�y,T�	���E~�I4CE�jC�V���r�,q�ep�EryR \/�rt��i ��V,@��+��M ;y�"�&�&HN
 �����j�(9�̌�w�@u�}G�ie�<g��pb%"���A����� ��)��X���Hwp���>'1}0���3��28d��Y��q�u�*���j��yG��\��Q��K�V��}J=�o�0����*o�� ���&*i=���/�����Ԝ ��V��d�N�]��et�1}s�����Y�ӞKM{qS!�Վ|]i]���g�/�j�I-*̳�lXXkL�e��L�ޤį�8�+:�[C��5OB�VkzA?* �/��>�K<}V��8���ܣK� Bb���!���l|lh���b� �ŕ棡}���G�g��&����an�٠M�l��dD��]���]� & �Y��X��S�F`���8��w�y�s�E�C�� �����MeL��&ݐ��퐍�}�%&U��b�E�j�H6������[�(0>~�>?٣<�u�����7�U1F�w*��8U=����O��W�U�����i�����KP-�p8�	�3]�:�!�+�<��n��a�*9>q�9���o��Z� VM��8jK�����@4��7d.G�rHT�tP�K�����^ܡ�l�`�C̾��5V9�aM�p�+4K �ol��Eٝ��������������w|w�ti]��3 �ץ�+Oz �1ɴ@��T�4�mAT@��|v<'�Rj����CP0uƼ�ӏ�O�_vh�R}�<��E`�dI]�4�Ӏ��� s��EwG^4,�K-u��$Nf��g,韪��O���u�l~��d~Rj�.����g��:`��L�-�}�P`�7e�2?����e� 4P`Z�R���*�N�3#e�f�}���Л�}<C������f��kY�S�r��1I;�&���N5�� �qL�
����}����2}g-���3@���Y9<����ʪ�7B�E��3r�R��ȸ�"XbW����2 # S�'�BNX,%S��1\�ը��d�S�E����̢}=�]z��F�m�ҁ!G��B��H=1��Ę��v�#z�D����~;c��u�to�=:ۥG�������X�sV�����g�D�K��.=l�D2A�݉��-qV��h%���uKC�tAۥSy��/p֬���ϻ�2�Ƅ�D��D�!zg��Q�"�y�ũBC�O��~����x|N"Rw4݂�9��=�H .I�`�ٕ@	�b�����UO�;ս��ԺU��Y����C���oc��5*�ŗ��&;{���� qD1�����++���4R�1},%���%>o/��KZ���OH&�ž�$������ˈt&�9�o)&a�����4�.y�pD�+]@�;B��!��7
�0y��6B�2�<d�ymɽ�`��E�bo���T�������K�zsd��ѮW��#�"u�X��:a?;�� �����z��2BMmZ�^W���\�� �8ƎV3u��"��z>-���m0��y��o��尲�������0p���Ͳ����!�3�e�z��F�� ͭ��a�:�d���Y��p2��z�b��H�������14�4�}g�+��,���z�g�%��IC1�8�\fχ�����tIR�������K��?=�$�Doi�}��[�8!?�i娌�:"
���(�B��:z鎶5ha���f��g~f���[@�#��^�l�g
@�SUh�k��[d��H���]�D������!��py��)�,��%�)���(��1�����`-��v�^Kk
kK��,�R�,����!웟М5�1
d6�CC˦],W*����4'I=�� l��� [9��X���B����k�����#1]��dA��Wamj��➗{H���~�b̮������V�\��h��mǂ��
�X�pB��Y�4�a��^���v��J�h�v�z�1,�У`P ��X��?K���1+��B�~�w;�5��/twK_W�ʵ����lDVVjycBJ�0��@Лu�U7��V�4I ��7�]@�ٓ�>��a�ɏt�MN	l��gcê`�����BI��";EX YߡO��qLגd��yRïr���J�6^-4���#r��y�r�\��!a�:V��S�&24$��`QO*é|��+�?9��\� @m�0|�����\���?h�W?���x�A,�N��ڐ-�D}�������ꉦ�3ya��i���N}WDW�98��l����༆E%K�^��Cnzُ��i��=l%�m�;]U�@���&���uZ�������������"��A�̀�%��'M��1I-��j�	��L`�þ�A�Ҽu�L��i%��!�OP��$Ӆ�h�ƪ,���&�"�c���(�w��3�H������?�_%��Ϟwp�	�c�J�<��eq���۟y�m���
��o���.�pk��ӣ�$�#�P#�H�#A�_��L� _?Z�3�͡���]��x|u<\OS-�����sw���8�!��*a�[7����H$�XrfH�.9���B������.[<&��a@��,�?�;�m	~ ���=+�u8�1W��&����ㄞ�b����Zk�O�V��)�Y_�ic����+	8��Q���9�-�V���LvI����iP�"@�<l���r�ޟ��v�UM�F�PcY����B�l��3[v�E�£e���w����I������'R���+I��qҝ�~�����w�*/Fu�^�S)ib94=��������a=���_�7�@���%�o�+ר�ҭa�����%�p�ɕ��p���wn!~h�y����K�s3���ع�f]5{��ߺf�V?x�
��<=��G�C��q�h=��t(T��Z9G"������,�h�f_^\��1�"�t��͑=��2ā6�.`��z��9Z�o�a��yЈ��lW1,D;q��l���	�����J�������}�-w�䡩H����O��ж^��5��t�7����{�i]�z�b^T%6���T�&,k�����bX�şC��Ϳ�!z/{�nׯ�^���%ũ^7~�C	a�#�^�r���x��N�m·��u�w4+d�Ѥ�>�� �<��/�D��U��rBLo��W�ނ����sشe��.��Q^q��6co�4��T\}#������z~��"~��v֓`��u^�ŲN&�}W�X�>��M5�_>�X�t�SXF�&�����O:#���C��~�㬚�8Oᱧ.��M��^7��>,�#7�(#�H�-����4�j�N��wO�x�8
�3���[�Љ+H��2�`�����Gk��BfZ����:�`�5u�Iͨ�����O�C��82�=�vgȨ.+P��:���������ڲ�G�l�
j�G����I��T��o����oY}pt������a���I�v����6-���c��ƻ��/�!y[K�E1�^�+e���P?��)�R��*E��x`�B��dMQ����)t�n����,n&��C��[9���3Q�bL�wq9U&{������M.q�k�
 $��P�=t�bC_x�湮=��U��$�筙t�5bBYG�I��p2Z��9�hOG�E�Q���2w:��H^��݌��F]��4��!m4��Ȟ��0qb��%��#*�A����K�*4��s=��?�S� �.�����-���N;P�-�*�w �k��g���0����a�� �G�Bh~V�?]Q%:e��q%�ã�N�$քX��=��r���vQ�����y�zg�G��S����{OFj�3EN�h}��lp����C��Ԉ<�ZR�̣�r�����m�f�	�˙ h垝�  bIK�]=\S��di�P�����	T[`��-��}Gj}�KM$��-��S�(M��[_��iƁѢ|D�n�У�[�i������#�H=]��pÅ�mُ���+fL8+kR��v�=7N%��^�秄��F�pG%s�lZsH�{��i$v4,��M/x͕��j�EOE�ȧ��7�p�o������a0��@��/��pv��jp�uc8�]�Gc��"l�(`fIf������h �'�8�
�WXJU �^�5� ���*j�֗��Y���\�͑Dَ
X�\{[Sj�G�),P���}!:�r:��l�g��$��H�ب�[�u�C7tۏ�oEDZ�j����
 �h�M�W��y�z��y�V��������<��bR,��dK�ǯN��omW� �}��Ƙʓ��}I�ܲ�J��5�.����jt�L��1
;��l��t�
�Q��� (zuW�q�
��ΰ%�wͨ��93�ǻ'����s������E|�>C�W�d#�˘�hdynJ�c�-�ϡCU
�OR�#x֠�
+g?�@(s��d�|<��:��n �ݩ"|������B�ȝ� �K�����L2��B� ��i1��t��U� 2,�b�. I���h��A��-%�*ZM��^(띎�A�Ӵ4bHI%6��u�d�C@^S�#��$WU;�E��9����y[����"����8�J��-M�T���^��(G�^�՗�ŕ�Qa\gn���86��֖ԍ�>���0���*��0]�\�����<��H��.'"#�l�z��n>xM�=�7�7��:Iͻ4��O��F�m؇�p�;��'����{Q��>v�Z�*�3ơ�w�@XeA�׭���B��&��n�ť,�h8P���c�L�E��k�	��WR�޶옴 b��%��������t�6w̿��N�8��m l}\�q�E*���k��B�<���z�/C[�&		���GA�^`a��� �����x��Š�q�����.ON��i۷��gm}�wwh��9IЇ��#��M�j���A|{]$�izV�v�`�L$|�p,C�.�FP�{����4�P�M��|�3!\�&�rk�u��I�_����q��0L�6��8�O�n�j���N�4����㳨�u�O%��K��OYL��џ�D�KaX��?o�Z n�N�XP��@�;�q�;3C��{7�AG�wz�7�)��+i��6�h��I�����>P�
i��al#F��e�GB-��9ٕ�ޝ�\5�X�Fڕ��#:�Hk
����G�o�N�9c�7�ҁ�Z�Xl�b��z�[�Y`����nUWS�/l��������T�n+���
[ks�}�j0�`����N��d�T�{�-)K�FC$:�ଔ�~���EokZ'>�MkZ-{,��f����e;����峾�ʼ;�L�p�sZ�I0Lȏscq�}��ET(v�
tO�g�m�PES�������#���2���*�L�k5���R�{�CLei�s���V��0 _�4^�ph�xf1��8�؃�$<��:L^�z
�y�����4Ƥ��%����p�.�E�0��~��iR�fl����@/�%�&������c$����ѫ��GMv%����B4�	�b)U3g��h�0�?�����rZ���-�<���o���pvd븩ݩ����^�J���u.��u��%���)):��gp
�J	I|1��#��'9���:}��\��g4�� ��QOx�d����g��{�.�o��~A!1g�A��̻�U�Ŏ���v`�,R����|�Q�MH�W�L���U�{{)�:`���w���5��
4��e�T�E%���dWĵ�ܷ_�����.���X��]ʾc�Գ>a'��B�g�Hs�~ŵ.��]��.2����p��ژQ�5��iA����M�TX�1��*P?�t�R�	�ܡ�T�D��NdQ>G�*�f�����(��Ed�Ǐ_Tg	oj�s������a�0(�E\�y	���H�1x�X_�yif\L�Q#Vw<WGa#:��H7o��,B��P&�\r SQ�҉B�bu��T^�:pR�*�<m+���R�i�x�����ϰ�e�����碃H�Dv�#.���RڍC��$�i��[�F�3�l���M)���s��ክ�#5�Z���Fx����&�U���;�c�-[�xY���3&S �KnŽ�qU��x�dbCf�x��շ��Χ1L<O��U���;���l�Ek�����B��}���t��;��$Ə���V�M�)S��\�-;�]���(?�ͩh
��;�<���3@�0�NC*7{��V���ן�	�]�:�z�"����Kb`yT=��g�F �Ց�O��5�p�b�Q@��
�W$cvf7�{��u�_��hN���a�!O}����Q��\�i�X��dM�Ё߄E�V������w��c���%�Nt�#��}u�#�%������Cf�*J`��+q#H��K� ��վ� ��>�Q,�)-�Qs���� ��9��aa�����5p�Z^���tbL�fV�o�c����:��d8�e�|�Z�	���0-e]菊&q>�j+j���@�!��L ��&�_z��'�����O�Cf�~׽kUS3�����P�5�m8��l˵�R��C�%U}=t�ߒ����Ų54$ґ����;N)+ [J���]��R���o:nUp-Z�m�Ґ�������I�O`N�L�c��t�]�#�;����f���|��exAs�%^^V�S,�����O�S��4�c����'oZ+gק�.(�8I����gThǅkD�+'��_7��:[�����J��jӐ��]�+fb�^5�C�8��p�qATq�������l#�R�)� ��>3*<���bR��~�?/J����y�7�y����֘@1E�]&6J��t��j���.�^P��*?�l&��me�S�P*�{�\#��`�3�AB��_q-TVR>��!S�Y��f�&��~�Sm�Yz����Q�"�=+g�
=a�x�:-�TURw�!EM�0��X���}n0��*�W�ע�ia���b�UZ(iܴY~G���$��g<=�b.Ʌ�	'�gt����t�2���^'�#8�!��PА�?&¾v��	��u(g��LR�:m�ۆP��3�Y;��y�pϽC�*,W�l�ɔ�h�#����>7�7Z�M�J�|��135���&��D������^�U�F5mo�`��?=�kn���)�S=�,�m����� �8R-q����?@�a
ĕHހX�G�N�f=�yFS*AGƺu��(�6����$(8�����(��)E1wl�#�f���%7��0C��y?������}v��wRu��JY�]�^��Ƃ��y�M�l���q�F�H��V��lC9*H��1 Ԝr��9���U��#�O9�gEn^�)D1��Ϧ���1U���?��28�N�{�5��)LOO����vYb1��_Ɗe����ft,<bb|�oNi���XjE+]O�3�.Z`�>�˓�$�)��(�|!MB��m/~l*�n@����p�	 F��i���r,Zl���s��G���!n<ٿC[��-��ʆcVkp��Ә &��`V�����v��6������FV3�v,�Eя�����sWÌV�8��0�/�������,��Qj�� n]!�>�1����mZk`�.����� y.�Z����OpE�^Z�	�d�کBE�ulR��8��#]W@�;[�x�hN��G�����qێ�^eRO���*5V;���q2���Å�F��a�fp�B?�~?n=�:�����.ِ'����:^T�E�lB�Ǌ�aY}�Oyc��J�Dڐ�%w4�~���Q�E@���W��E��A���#d�L�^t��'�fSKw'H����
��n�5�X�032�����D���x|��bV��=�f��s�v1%�hDA��GF���=�!qJ�(K+�1��־���"I�ꔊ��s%s_�n;��3�p>��W~�R�������n��"$�^���*V��	�$:�h�:����L��Z�������F�;f�Hv�.鹀!�dE8�M�~�N=�E>�OG��6Yʍ!��m�?}�Pt��I}�7��{$<2S��X`�q�
�Ӛ�n_��͝��ETӹ�,;�`��$�9�G�����_��Mc�n#L T�wM:P��C�wt�LקJ.�`j6-�]���.���Q�����V��,�D�<i"�ـ��*�v
 � ��t@��vђ��}�f�5��*i�ZMMe����a�#7*���8W�/?,��=嗬�8$��T�d|����/����g֚�fFo���+4B��������`�?��Y/
�f8��^|n՝_ؗi�."N϶����#<�]&mr��+�LxR�h�j~��K��VjD��$�HQ$ ������д�ġ���,���(����ú���4VZ�-���&�����i��X�ٓՌ�1ӂ�X�������,@�������H ���Bt�vf�<� ��	%w^'kز�T۷kpp��t�L�H
>㇮�F(#�y��(�pCf#�;�;n䔫�%��N��@}o)/b[�'-�g`�KV���K�ն׆�Ϲ� ���)�":j�x}g\�M[�lQ��7�Ä���$�ޥx��,|�����jC�榱�К~�����
t5)�+T<@�a"?��<!Ә{V]m﹋V�/� �>���c�e���[�Zq��y�4�t�K�G˟ �ۊ���(\⌾��[��v1��&�돢8*���0d�IЕ�3I�y�,P��˝��>>�M�h1�qܒ��%>/j�r{U�p�a�K�}߁�e�-�6�mD��ޢ��q�2w��P�34ܑ�J��0���j�1������F�9i@~e4<(�bp�����Q�*좼yw�ɣ�Uu��N���j�@ �n�����W��)X��t��W,�/��j����a�B�E3v~"�c}E����	6�[$�⸥��D�{�����_"����KE�g�\-��(��H��;=(��8E��HO�P,]SQ��,���y�ni���C�fI��hZ,w�xq�(����ɼ����Sn�����>��WVN�/�:L�*p�qX�Z�qB��u����`W�Jג��Lk`˦]g �:P�/L�C*�$Vk/uT8���?3��d�e�5�Y�*f�u`�z��3~�|�xlA'~�lC�R������J��t�-���i�ha�K�*�c��-zC��L].���k¥��-)�F�2&��f�&�:����u���јP|�;Z�Q 8D�Lwz�+� 뜄��+�{&a��i�̝mt+���cgmq������r\��ᦘ�����"�C�m�0�|��w��a�g�����o� D+����B�Y{��6�_��۫��đ� AM�3�G-�v�=�Yh��c?���[u��B��;ذd ��FE˽�P���[N�:c��P�Hp�p��I�9�t����rY�&[��i����(r�Iv���䧹^�<�l}n}�>{��K�9���߄p��Pi�sJ�!u����5�}��Q�b 
�w��S�b�\vV�vȂ�����Q+��P�4��)�k�<	�C��	�hfr6��s(A��7� /'^%�FGY��?Ť�;E6RuRj�8���9�ҝ�ko���D�]�P{�Ž�W?N�U�7{��'<GKU��A���u�or��F�Ň��w��L9���%$CZ�û�3t�{"�Z�0����M9�1�{��'�D���k�E��}�X�3�i��|rj�x��G�lO���e�CЊ����/?��)hw��7�#���2<���b9�EC�QƔ��m%��1��4M�NzR������yJ����[l�����c�έ]Ё����D5&L�4� v3�:�6�
5��t�Ũ���d夷�JZ��}gXTGH/�l�,��?�#I��ւ�2���u��+{.��8$a*@a����r��	8�*��+D_ķ�y����X|���x⋔��5Mr��B�K.�m:6���I�UH
�.]%xE�c=Fv{���w�M�hV'���^�2�P����}"�Y��1�$�����]�>m+��u�9S��K1�g.�	��2�~�ذ���WX��K)���gJWT� g�����Ԃ	�lV��M��z��De�T ��q�;���� ����Ϻ-|�P�F3�����k��ĺ��� ԛ��p!r�_wsx\%É࿤j�c
.ϫ�<���G��+��B��"N,�M�f�`�tP��N�[M�)C��������g%��u�ݴ
����N����>�%W�m��._,~MM�iq�.T�"��0Kx��M)�� :�������� �E�����Cj��6�ь�&��'wf�ټ�'@��6>�9�y����c�?s�WQm�5~��MLh����<�7WU#_P�=���ϙ��A�q#��E�8?!�Xk�� ɴ���pX��0�$Q����u���w�|㌸Nd���o���k����_�u�L���C��MlN��=��5<l�t|���ϖY ����d�x��"(¾��b�ߒ?�
#��	ţ,���a��t������+�^�����5�]%v�_���(F�b$�&�V����}l	����������`��%� �C��Գ�sn�1tQ�Q��r�����;������,PG֜�O���upO�*��q�)�q�b�!��� �%K�̤C��g���]ez��kf����xK~S5ˈA�6����u����C����8��������cDt'gx:��ü]��.�3a����n���[�0���U�1v�|Q205���/:w8Z�%<l:�T4^�Ε��E�6�fH	��'Of�>!��G��0�����'%�]�e������K���% �����g��P�*7��'շ�A\J�3
Ci�,sTC���gA�H߶�ж��z5��&b/M3� ��7-Ho��9�a���5���<�򌵤�Y�-pS&<�<�i�FU��-5�G�8#ӌ��/U��	x��A�F��#9���Gz4\}|�G�a*��xr��Ziqk�[��Ƌ����q�%�t{496�j�>/�]��f��b���
!o�Ǆ�z�݀��W��H'��ja����!��&5�<�҅m����q���%�ͮ������Mi��ڹX^d�XD���B,��.N�����Ktk�N�__
�p�T�M�c����s~�����.��GgX<��*zA�Df�W���e*o�d�ͩ/���@e��l��9�pӫـ�0�*7��įÇ�k���L��T�g+V@�'� ����G�Ť���j���W+ҹw:
�R�%�;�=�d[�&�������)�q��:�V�ʑ