`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
dYoOmr4Rlja4N4r2UIDD906Ruycb6YjZpabTrnRmuVhUC1nUwvciJNyBzQqHNvZGSD3ofqcUWmyd
9nE/WxmvfN5Mx3kl6pJ/fyZCcMSDk7iyImwiic6QX9YhMRsYoT/gh9qRngwBodadprkTPhCq18i4
Tpy4tZnOXBklndzgEwJp3AXhMHd21pvkX8h1J4Gi6OUMc036ZLBmtIqwxSFUDT8cRmGmQlHJHRdz
pyZH/KEKLAn+9STbMtr2KV782VRF8hH+WaG+T3XMf0D9+FGwEv7G1nGkGxEaOTVNsZUVp8jDCyIv
4atwAPrCl+VBYwzPx/O1jmhx3RLaILLp5FOyxA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="Fb7KGtzGUnj8Bm7WzIq4taLfgTLWJpetT8T5u5f+WzA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
zsug8ZjSkHg7k/v1ncIyowAMaTjzIfDMcO+OwdRhh+B8g+jOI9ymtmILg+WB4GKUGZzKgyzIJw2V
MyKHjGwcVh/0k66glF0h1UrxwA8wnBjRqtzBbeJxwS91BpLwQn3dfnmavtyLAfbiao1So4dRfpWs
J+UeOGbnMe3aEziUWUqbErlaBz7YXN4406LUfjq+QDyFYivShe7YTGHNPq+3qHqoqB5lxDSQoAtF
/CMbEtvmdiaiBLTEnPIXCeqnFUcnEsmO+IGunAZAsdvKr4SjoPGw9LYEGHuWwfqE7Id08TYTJvVt
AO/E2OlDPC5Fmu4zI2OCoLdueR4qScbh2n0ehWjDkxlQuAxER2CPP7pfU4ni8G6cSLEARN/+ERVd
7JHaO2RHzRlkS1Mii++htOoWIANYFRnSyeivPd8GX3yJJG0J06O7KrZ0VyFWLCHNxQBFX6eGE3h1
HHEHAQBVJRluwaxTp3mbNRvpL9mlaL/iDfelE7nCXW45mtBwAcC/PMN7OnFN2JSFW6Ew0VSL3hQH
9jPFGb89c32kmVxSzp6sJvdNOSbZrUJmgEjvcHquEmpoAjrdWNYguQjY0Y64TTq/rsr74lJUGtdo
zwu7xDwn0RD4AUg2qbvEsMV8QWP+i9Uy7zAv6XAWAtpwDH6ql7lP9dSRf95wsnu/5sMAvvSSLGGj
TMG3hVrtQfGY6YdYDrrOAfZSIV9s0bQEWXr0Q+fUjkIDPWR3JSnNrEntvU+xUbkY1kea3ipvsOBK
HSNrvi21Yi40ohHFkf1yq38Q/K3vfPt0Faq88yga5HmgzEa/aczrxnXz4VRomhbLlv54strLNDIi
4gYG706BOvI+JwGFIZiBRb0KXIw/omVx+TjdZ6CAS5x9zpEGPzOkehtVWzw+SCLyKGrnLQLCn0O6
TVIjlqKMCcismzEf0dVZGrHjG7qYgkx0ClKxvuVuSw/ovmiw15lcV+zDQskq7OSxkoeCeBGgAdnK
slrBPYC55TUpGLxtGwEoa/jkmZymXTdh8EY2p9p5/yfLqpXlrrX/69THxqoIUdV1W+yRq9ifib2/
KbBeFb0Mwy1j6U9zpkp+yVBlg7pFESuV7N7CSIXwk9aaeYQZthbR7zZhZMM+UMj89U8Iv140Ui8p
fQ1okGZEakVJEZjOZzliCY3yHq6mgAijORlIsrKZNOfXDZx9acMMRMrBLV+wYUJV9wGH9s1vJIpb
yoaem4+CrGOOs02TtP1092bKbIoNIfOabV6ilxu7GXKAjrTn2I5ghoz7e85fBGRnjieVvQtvUxD1
5OVVkPCkWN1sq2t9TEDzJrrBQxzbDvTp+ItNLgVM1FsdyIsCsh81un63TCxcVuOBwwdOBwdoUhWZ
htBGauJt1avPLBu3bTdpoEfB1y95ZsYRHAJIId2pzBLF89XZv1wuqppGXY4HSU1fpHBKUKoYvKTA
e10Jfuu1Lg4QmXASgh5KT32OGPG+O2nhq0kdp/EjB5NYJOBCXQhvl8tHOSEowlHycXbjj2E3oDa2
qxKGU+xbYUoddFitoSb4sgpfFw6thejPzetBLgi22SRSpCRs4h8D84iXuXPEbIUhoevwB0OpQnaf
cRP3jBkg76rMfNkhjNgdN5OZveA5w63xkYi+mMO/gCC9fwkgHxsKYEjkuDpk8mTl5kxXNRywVFvq
6WxlLxPQ6hvaZKBLT2E3PiJ4Y8x0tvUZXXZ2iq0gQZwJlhBB2GA+1lFuUDu7pgbbSkIC1n6DvahJ
K0CxfzcLpJvzmi5fi0q/qXEQaZ2U6nFrpl5/GqGDttKcpRp/ZPu4M66DiJKZTTAQdtf47gqpz6hX
iAzx4Zm5weS8i5D/OsAsRMjHztul+l746b+XZQoOWprLGm31/diDbKc9CXmikwLuOoyE9DjwMnTv
phEhNJowoqVGBFAZpaLzZrL+NfrG2ZBsA5EyQcwpgSNRXt7lW9Gxxvlv1KskdhxtQum6BEwKYYWz
fBZjZ6BAYyeqtQpVWp4Qd3tgZIjjJP4bh6TjuQlTa+XRssCXwspDpryyte4eazjeKT9OR2dqqBB/
y2WBstWkhowqZp6eOsntm+a5ChIKOekHmpjKTnYtw3KqZh3wWRSfhY/iiUzi
`protect end_protected
