XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��,�X�����0���Bd�K����?no�#��%u~�TB����r�G7������؏ǀ�/Q+��i�B���4\`�6�-)���_j`���b��	|�����t��5l���啇�I4������!-ڣ4/L�*��m \���Qq�`їC�x��(�U��g2u_�;��W
O�����g���8�}��БĪ�@�#0>v�\��R
��V���x("1�@/�� ������S^Ɇ�(�HA]ķ��ˮzک���'��P�I�N�M� �zŭ�jLe����F��i^x_0/��)W��6��7t�]3�AAdL�C�m���q�%��֣�vV��Zw#����r�Z�c΅'\s�����M�V���6z	?�쏉��d�غ(��L��Qh�P�I��5㤀d��ˋ�gif�!r&�۟WI�-�n���"�w0�G6&sn\O�@�=ku8P�ȋ�b����Y>��:��i�ܠtR^��nO�ھo��c��B���[
�$�=w:��	����
-�U�(&�A�۹����yr��X�]���2Fc����fE���/�Lg"��|^&=��)���+G��}���\�#:�fzA��{ ���&�1�A;Z��%?�ݟ��̶:��@"�c����J�^P�] \R\悾��|��<G��O�r��t��@7��(��K4D��RA���_��v���A^ 2\I���^7#�"#*��u(���8�NH�o�������Ue�<Y��DXlxVHYEB     400     190xRq�+4�_��ْr���R�G�Sq�n
�r��X][~�xm�>�yg�h�s<R_��x��-&)򢁁à�n���i�$�A�>�Jy9�'�x�3�̣0��`�զi����s�A��w�h���=��b��g�lh�n6I<E"�@�M�pmƉ�]*Nn�;�������2�pob&U`6���0�Yc?y�l�
�R�
���()*h�N�����^qIs��l���֡6=�*�I{�Az�B'Q��-^Wag	x�Um����x�ysw����<�&����d�ۇv��"v_�ܹ|[��S�����;I��Ƕ��Q�֑��*�46���x(Q�a���1�F�NM��7��Dt5)�&�,!��"�زov����
ػJݝ�_D XlxVHYEB      3f      50]u'������Ew�Q�B9L�Z758�FG��_{^X���K��Lڢ�r���N�ȏw!~[���r��p��"�M