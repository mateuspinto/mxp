XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��GX�\�a�\�t�|�+��h
����tG}R�L��1�'�aSD{w�v���wl�z��50��/�3hȬq�r�����?� $���ڏ��L�	K�MX� t�-Ro��F��i�iǳ}:�]}�RDi[�[�	"�'F4,/�	�:_~�����>a���P���T#ʁnU�Ώ�=��xI��J]��6�;�AZ�=�+�������`2�<�	��>I]��(�ovv�Q˨8'
�}�9�8�g���1�QҘv�qA��1��ٳ{�;.*����-)K� ���˰���ʓzܱ��S���'J4`7O&��r�=��4!�,���w'ii�@�y|�.��H���)��3�~����I��қ����dd��Tp�Ɓ~�>T���t\�(Ƚ��s��M��p��w�� �e�g��_
s�#Ӑ[�,mۆleݐ�}7�}�b������S*�6
h��JP��a���p���;�Ir9��1R�,,fB��5 ��q�-�Χ\�e��f��(dB�/?,E�]��Kv,o������6U�_��2g��Y�����QX�bl*�Џ�%�r�MI���ǢM�{>.+t��#����FB,��hd�V�RnU�ǉ7b+~�����Ͳ�A�FE@O�j���+�I席�r��ނ��F��H���BxwH3��?ʦX���Y?�N�:�P��O�'���)�tm��`�&;I���׸w��ۉ86�g�3���X]�����ʄu/����{�{���^x�/��%<}��Q��XlxVHYEB     400     190T_#�AzB��F`Re�چ��*Ov	2Q���p�]Uy _U�R^�ں��ng���+t�T�6�M��EH%k[p:H&#�󘇶U3uE�M\��'6��U-B�z�g��d�bb���TUWv�/����yB���Ԟ+��:�.P>W��W1㈳�*�5������MY�~|�i��������!�	� �P�������b��۷�c�<5I�T7""S�-2eD�&���E��ғ�w��������?�_n��\����p*-���u´�I@=�_���.�w@n��	�����{J�ǋ��ק1sL�u%��Xw ��} ds�<:}v��Fi2��AR<�]�����WF_E���h6&܌���B.��z���t�S�Ϣw�ҔJL�Y���I�$XlxVHYEB      3f      50E�o�����4�~գr
'���]�J̩z��5$�1N���Eܟ@pz�}<�����޳}S�v ��
�/��Pz�(�