XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����7���X�[��M�Ђ�-���3��W8���^*�ܶ-�T*d+7�AQ��!ݙ^���w�G���Hk�*e)���Vz���P�F�z���p��6?U�²{l0�J�F�����(�fo���/g��7q�|g��s�F �@u�#K)�i�����a�Z}?K*���r��)��0�!�K�F@'��%����n)�ǭ5:`cdؗD�_����1ٶ �R����x@�ʖUh��{1gj�'��������MIM��=:1����.s5!\�Һ��C�!�#�/dĳ.��ͭ�G���dT0f~ff�νK���=a@�rU>��o�'J���6H��O�+�aU��cY���Jn5�I(3ʀ��?���,I�L��y�E�]��P�&�zib�4��K��+�VLE_=oƼak�RM%�����[wK�ґ=���t��}����b�f&6��Z�zK	~Є]Ƚ�~��b���;(�?�E�a�c�
fWCB��L�;X��1���?�(��q�4ӭ�XϤ�)f��5����]�������;�#B�T��XZ�8�)�`����8L='�Մ4 ����}���I�'EMۤ%��pS�Ifz�4�}�5�I�1�3��4Y��X&M�E�Y��D��kC�˗Dڱ�#+]"3���:1v��$�� ֯�@�"���$�A�����LD���ڰ����&\�U�ێ�m�F_�W<��t���f-�(�/�f2�=,n�Q03N���t��XlxVHYEB     400     190�Zn��� Ӏ�E�h�)x�h�mKߔsh�rd��'��޿>�U݋���h���f+-cd�+��(֋i5�N_�w2����<�����K;����MG�+.�m��ۚİ��LTKR�(%*<�m���s�S4�.�/��� ��)B�h%J���נ,�����Ғ/y��5��\��{�;�N�Om�������(�a�%�%sHbqE vk�}@��e,�_�u/�����~9��<��j��(S�6B��^0�Җ�(R��Y�SI����e�{)כ�F*_���V��!n�a���;beF7����T3��)�S
ݦ�~�;�BP���\����T}g����.���N��c����	0�5ެQ�B��������P�+9ȥ7�H�XlxVHYEB     400     140��wup���V�u%��`X�O���PJ���������M�F�3.<����*L(3����覾Klz7�}3f���������j0�4�q�m>��8�FP֔�~��=B(������Z��k��~N>���3q�F�_X*�����ʟ����f4<�����(�ʢ�ѱb�����!L�7Ά�5�G���ԍ������t�y�m.� ��0�|�1�C��9�'�~���kN3c�����C�����(`*o!��V�E���/�5�q�S�Sb�0���D�����i�>���C�g`+1we���ԉ�La���^�n�XlxVHYEB     400     170+ՃQN_��)d���0�3��[�M���J�\��2��!'�ҿ�$ٖ�>�ۛ�%�^�[VM ����ƌ�e����E��U˚�����T���G�HQ�f7M%�8��t�ۣa0��5r]��J����`�4bۂ�Mxv¦�Y� ��EJ.4P��~��4g����ND����϶��Ķ��	�zʻ�t�2�o�R�]t���T��A�D��P�+�pIx��GN�-�l�ї�Z{L+�7�V&:�
��~*�IV��T������x�Ơ�eV���!+?�B`�Y7��Qq�İ���]):���o���I)�\���\<F��#��.hyb��/H���e=�c��d�F�	�7������_ޯ�XlxVHYEB     400     130�UJ��+ǠN�#�d?S;����9]�+e�@N���~��9�/߫��!��8bEd�YT<��t�t0�� %4u���o��%�d�N������f[�e���a l����Ds���� g�����jt'��n����Q4�l�������j�Bӗ��wg�}\__R��灦�����kǭ9�b��uh��]�g��~_4�����~� ڼ��m: �����x�h�!}4��z�-�(�h�&�b�8�錐�2�4�?:!d.3���G*����cb�U��ڴ��[s5!���!U�V/V�XlxVHYEB     400      d0�Z�/j7���zvʆ�4��'�t�T%�)ս�7Ȏ�z�uU��O��h��ɤ���9\q;X�B�7�uˢ=��Kg��ŝ�H&)~I��
Ӣ�������[ڌ[���l=��Z���{����C;�}.���&�0BM�@�J��b�'�yc��%�\`~~�Xi��9�W�T&��4��L��e~�]���y_�J��әXlxVHYEB     400     130ܜ��3�|
���m����%9�DцZ����K����,>�d=�E�^�D�Tko׌H5&�:J`�/��˒$�nl��P^V�v�臗�\L�%�&�4r�Db{|��x�~������\s'y���)Γ�'��\��z��OF���Ep�
��PS���όP�}v9Xeo�)�*�8~j�DY�����xp����]nR���Q����R!4�����|<�I��v4|iJ�T�/�&�a�^�aNl��?��e�ม���;�8�g����Ff+�*Z?ٵ-5.�m��#>��!�XlxVHYEB     400      e0>�[E�+K~��,� �xS@��`���;��غȪH<qY8Ckf?�yg��8�p���$�Z���8�̵�D��D�����ݩh~,P��I휶�>ϊ��p�u���V��xbeKH�(�[�ޑ\��m1���黥�έ��	�L?��݇dG7U!���P~!����%K�@���+-�$x��M�yA�@NnN�(f���-�PUM1a�V��XlxVHYEB     400     140tkr>�'�ex�28W�O���t1vP,;0���%��B+���A���c*UG�ŲZƄ���݅��Tz�%�*��ᯪ^̼��mw��CL��j7gw='��Y,/����Qm���y�|���@K,��~��ϬH;
/t�o�?��R5k�ԭ̚�1��J����s�w?�8��<W�[�K� ���(9��g���{���ZӋ�GG��/`\Q�|�Aԧp����6�3�iN�G�s�6��]�n���o���3V�e�0�lb�b ��8�cRQ�ik,����
Aw�ڳ'��V��p���UT܄�@EXlxVHYEB     400     180�x��Q��J\ r�ɭ��<E��(;\�u�콌QU��u%��B���p�S���9��
�
�.�!R&��|^��ꨢ��%^ ��ۺ��_��,�pt�O4�([1���y.�ٴj�c Lkhz�K�_�]x�Jm#y{�*�@]	������?}d���pN�[e9�$f����9���6HG�T���B�.:�{�A����g�φV郗���;ͫ({�����ѡ�/=�fA-@�+ �i�f������Yk>����da��5F��W��L=%P#�:�1w�-�4�aH��������@���W�$^������E�D�����x	���|x�����5y�o���p_
�	Yh�?��Zh�V�>����w��4�nj�YXlxVHYEB     400     150��2���΅�c|��&����V9�L�����8���;��_�׿�uY��PJ�Io'a7ˍ�f�e�1�͢(�Z�8���� �\�n�wC᪃�~d��%4q�%kS�J�|�yK��h	R���y r���p�Ii���ݐu6Ӌ�sq4��?�8��X�@>��N��xi� �m�C��\���9*�Ɏ_FC#��~����c��KX){=#�\�*`ݲrs��+( ��-�2d;ƍ���Ȅ�NnQ3�AѭҌ["�B��Iu���g�[Lw�U�iY��;_K2b:Y�c�����n?\ЧÇC�r�Z��A�����4�XlxVHYEB     400     160jWXV�.�[����K����������'����%���(%�'.j�D �fT`�LX�E~��,����vt.��U�7T��ȧ��L5��Ʊ7<LM5)�݊�0��d`�Ӂo��[a�MQ�-%�kZR���d����v�����5\E5��;;���s�P���_2R3�Z��3X���M4�'����=����u/F�d�['�"i�i�Áe}�z`�~o����Ѭ.���Y`��AfهV�q���'J�8����t�
��B�����`�Ƣ��[ş�ؘ��ۤ���W���&�G�e�f�+�h���BL��9q]��
O|��0'����;�x�>����LpqX�زXlxVHYEB     400     130Л��`U��;ƻr3�D>�C
�����n�R��Uz��Ҹ�>wۜ�w�6�}<'G�eB�Oi��YӰos騢��д�(�0[7��}�1zJ������ca�����U�"��y�d�4��[��I�3 �ɣbsߙ��/ʕb�����)W�[��,A����Sl����t��J�Ko�wo��=�"�D��)e<���Ɩ�^���@��ؕQl�9Ұ;:�H]v�k�2�"��'^���s�6g0��헉�{�b��/{�����x��sڏv7G<�A��}I#�	�NԖ��XlxVHYEB     400     140U"�o��F0Gt��5���nQ�H����3�I=�Ǩw3��K�"�<U���ڙAM�TK�?tq���U���
Gp�K��kͰE?���&�G �KxD��3��w���F�"�IRr��H�'31K����z�-�7�"� �kջa����	�%c�����p�NUȪ��8W�HL��At��iY�7�����f��!�u��*&#<���:�?�M�ʔ�׫�����4oqC�	8ο/���p��czG�(��8���0I��� ��o��[�#oʔ���!��e�o��{(����=��\
�`u��n&c`�XlxVHYEB     400     1a0U�U��V�N�FA�S�0���s�h��
T`:��#2*!�i�=y���'�߸�w�u���KU@i��7������{�[=O� D�L�,�Ȣ�iG�6nt)O�{̿��>��2纅�3r�S\���v��{o7,���#N�zܱ�d�To���Sg'K"H�d�n98T�#�΅.����۾��FE�&I]|�n�D�Z.=�9��6�n\��}�<>���g�À'i���|���8\��[E���vL]qK�Q�b�RM�*�WJB�	��+AF�^��M{��O�n��]��
�I%x�:��}�Qٶ�
��Qx\�c����)X�CX��Zf�J�}^~0(�N�kK�n�����3�%�2��hW1�`U�#�MP�&"�.����s�B�8~��*}� �e����MQ�XlxVHYEB     400     120���|��Z�p��.�&�$�ǡ��w�:�q���26P���d��bt���A��(�1(] �<��q<�+B����;[v�؜�	�e:%b�ܹ�A����D�α�L ���JLh�.Α�4G�T�>{p�H`[�>k:t�5��sG�ȕQ�Z�`�����t�5��V���t��c�`�g����O���˂P�u&M��ƞ�
��d���ȥ�[ׇSkʁ������������� ,jU.6c�EN~�d�sqч����BC~�k���f�+>a�XlxVHYEB     400     180t��J/t���I���qOq�R����2@�N�s�K�;�g��Dp��%	as�����ĩ(**]Bōվ��a���������+��j��0\� ��qV���گ�K#������/�u.&�������ԁ�Rh�e���K��f��,֤Č-�8�G��;�|�[{1�ǉ�j\3�d�Hb���[��q#VzI���t���G	|@F��|���E\**��Z�J[�4*�)���/�jX����?���k���2;م(������@,�����#�s�e�Γ�\�b�~Qm�O?� A�ff���I�~:<�c�}Ɂ-gցB���}[�>����D�ΰo)���S-5�h�5���������)h��V�
A���<�N�M<r�m<Ƥ��XlxVHYEB     400     160BJ� A7�!�GGaq?��<c�f�(�������3�zÐ�a�E�\ޏc<��̃R}�&��d6��E�~�7�A�&��$@�{P�y��+"ګ�uч(�5�����/R��t��$�<1H|d߇ʥ(,�#�E*�%�9v����ko�x�uu�Aأ��/4^�r}rB%!x��KkzP��~��n�:��i�Ƒ!-��53��� �*^�=K�G���rD�����y�wk�� տ�vE���m3$��l:D������<�<-�S�q^�NZ��V�����W��	�xZ|��ޅ����s��֓\VWF����k�0�pK�VANHB�^��5=ȧч�J�XlxVHYEB     400     1b05�7�ron����Sb
�^#�l2��>=zc]��^�&�X�:�8c 7�\��EГ?J�{�x��&�X;�l�`E���� -!Oˑ�4{��1����Ƙ��%��F�俏E�?h�g���kLÂ���DT��O:��M�1ؗ��zw0/ы�[�X����5����fBɐd� 9|�ԅn�����U�S꣕�O����d"Lj�A�O�}�1�����%�/t�IW(w}�v��ⓣ�������$K�_u�h��TJ�C�Jk&�6ɼ��5/��A�DA����!�<�J"�'����i��寉��AŎ`e�q��\)�֕���R��o	�m�>5t7 �0D�X��8Zy��,C�Ev�8D���H{� �2#��(�M�X��c��`�\!��OQEk������k��롼#�?XlxVHYEB     400     160�d��
��Nl܀�>T�ه���G3Հ*��<e��$�j8&=���S+���i��K�V�6��2�a�ˈ�vnRL~��f�l&�*,	�o�M`��M�,X3�J;[*w`�{$$CE"�J+��v	W(���Þ����?N�x�#��۪��UK���l�iLO<ҟԅ�j_/jǆE�OSI9�8kNݽMU����+ؖa{$m��w��H�C�pO\H�D��]K��m^0_������?�6xV�n�/�lm&clq_��au�7��������&��<�k�\a��.�|�i޵��0Ƅ�P������ŖlSN0	.�S���jyݣO�03��:�XlxVHYEB     400     130��	�p�W�?п���_'��ɣ����;W�Z;�׼[��ܝ>?=��mT������upa*F���uK �[`|�2������\�1�fte*�o{r�A�U�S�ߝQv�<�ZYy����p�z�S�:�|ﻪ+���w��9k�[���#�ǎ+�nV�\�U�X�c<I�\���A���u��KI�^`>8YU"�#���,��B�D)���4$;3���a&F�*`c�����z�cF�֟g1���6n���e���*@�e��A$�BI� 
Ѥ>j&��� {��8@�B��߾�XlxVHYEB     400     140�n�75.�r��9�ZaW��#�O�<����|�	�@����Hv������O�K�F�/�6k�X���4�l�Ah��8�7�P����r��>}5��y�PS,[�wGtlz���.�!R@�"�#�)�-I�Z�������4�U���h�&��Ȃ���_�쵋�=M3�ª�]8d���w�;Ԡ�-�]���]��u�$��+��ϦE�[0|FJI��[q���q��:�����C1�<��G%�1���_O�0�U�� ?�
ѿֻ����[^�I2޹�ՠ¶�Z�h2���F��O��� �*vц�XlxVHYEB     400     130�� �xvI���YQ\Tz^a6�W��l#4.G��M�-�=O1T�D��m����9ֈ�������[�_ҏĥl�|�)aZC5X\gJ���@'y-�!^��$�b��N�Ս��`D�#��	��)��}�b��F��`߱�/�=&C�-;D�4��������gݕZ�p�&�fZ��5y,ߵN��
IiH��hEk�a�)���C���!��������H��'=>K�����5�R��W�1+ɤ��o�,E7����տp��Ȓa��1�Jq>���ꢾ�g�a�;	�ڂ�
��8WXlxVHYEB     400     140}ʬ��2��kC�dkK�XK����D��~'��T�?��T�sE���c��t>�ݧ��,ʪ� b�n_�D��c�:�5�;	��?	V"h#=lیB6�=u���F�� ���)!�lLV�ӗ�,_a)��0�>���BI��v.��ak���dD�p[���Ř�^ےE�]�,zj*���8�%s�J��
��5;���Op�  ��B@�p�h�O��P�p���B�R{�\/� �*�)��c��̦&;�K��E�XU@��7"=3��RNn���;N[��팓�����/��Ȧ6XlxVHYEB     400      d0�`���670`hJ����C�b��-a�5�K�!��h��{�x��$-Cj*�#Hc�4T�'.�,؞�������#()�R�q�Kk�F�%��i�dp��] Ǉ��3T�H!���HL�;&�s@n�mlIdx����6٧ �7&�?}j��s̖U�Z����\5 �O�XD�����-u�����}<ug��U�K#�MSgXlxVHYEB     247      b02�Щ�q�u��6��Pl6�ǚ}������"�2�k�D�\(���c^d������k�XͶ�:��7ʑȅi5c:$�I`��hUk{<��E�i�(8Wm^z%S�JUWZ�����@�����xNq�jv�3��.�!�hT����9�L�6��:��U:;D������q�Da��