XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��P���M�@��Jçd���5���a1&�Q�����|(k;Zׁ�������0�p��Os�BL����!�Ą4�uڶ�D���Kn'�.�O����$�"4���5z�J<[v�)w��\AR��Cڭ��sr���8�b�b1֥�z*!�
� E�gs�_�����#�;�;���Q�����x�ӯ�P�%���z��D�r5_��|��Ç�� w~���L���32�%�Z T���Y ���k�̣�G	�7v����U.��w��
.T�<3��+w�p����J� �][���Rg��v���㥞H�|H�M�����"���ZA�������Dj�Gh]bCt8����ZH`A��a�ar�Z�	���.6Du�:�h�*�)�=kPK��:��:m��~/l�F��[�|�-����y��t��*HD)Q�&7����֜�Y�*����ʝA�I���Uo���㢱 �v��a[�4a��� \I�����4�<�>[l�621�ce?}��5���aq��s� ������ �c��ƽ�x�q��kY��a�I|��Xz|���W�ɫ�m��0a���n�C�Aj��w�"i�0==�����q�9ԎJ����K���R��.�ԛ�G$�?C�j�Z�2ܶ�=]��s�e�sl'6W����ik24��C�jH��ۓD�y���A��Dk��2K���-�9Y�e�>��W�I�&���s��l�Xo����Pd�@nt6?�$�"A�XlxVHYEB     400     1e0�*���J9k��Y	�����%E.!�_:�K��H�:WK1[��^�yyp�t)��!�E�Rm*��S	m8���JD��P�Dzb�)�08I�Kh|�Zw#V?⌽��/�~7K4���T'�
��^���;#�<\> c�'���'C
�-�胼�q��f�"�p9:1c�SN:Jp� P���U	�?���_�� 6���s��yP��Pfm��2���$��!~lV�|׆���#i��s��M�z��l��y�H����-oQ����1	d39�Y@�q�_D�r�م!�0KvYƪe����*uk�	E%�$;��u��K`��a�Κ�/������a��06�w�N���O�<0‴������se%���sb�F�g�a�x���M/��=��6%ϔ{U1��C�ѧU��G��I�	��\K�V>��m\�-fr禝��N9�S�:9�n,��=I=Ӎ}��~ᓿXlxVHYEB     213      b0k2 �k�m'H�r#�@4����^��m�}���t��H,��Vͤ�XGcj��= ��+
;�X��~a�|j3U�j�zke
J��.���Dy�v�v8ꕆP.���1g�}fnN�z�g
 3QOrv�ژv�:�|O�K�1[ 2��.z����Y�7Q���:+~����8��