XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����>�0)1(Om��pL	���LS�:|��Z��X��Ktnm+�6�=)����S��IGD6+Ot����Y�QE���I_�bt! ْ�$�ȯ��>�m��BP��{(;]Ʒ	�%@'����y��,����2���a�c�8ɑ��J�k#3�oj'�D�!��H��@ �(!�"Sؔ�7�qh��Љ�-M��H)�]yW�J���h���$��֕�:�[��fe@'|sw���D��C��Ƌ�����B�zf��J����
�P!�܌�OP-k��_���叨%��Dq�Q�Bސ ��'`�z����@UhU|`p��t�s���)z��
��w Ma9�׋�ϙ_�V��u9)g�+���̶���j����C�B���q�v$�o�o?��� PC��0��R-[H�*�vc��S��wϲ��{��{	FR�xР���e\��5AK�
dE�N�O�#N�����o�I~�0ߧ��7��f���9�7���� g��(�`�qZ�R��y:���v�MW�8 G�(P'����Rn��
�\@OE�e �����rw�"#J6
��`۷��ﱎ$k*��u5m�c�?�z�����ך��c{�+��կדġ�u�A�`jq�̘=���3�ԗ�,>9aͱ����B�O�خZ����)��i���]�H΋튿6v����a��sy�W�ޅ���ǸS|+���4m�H�����i��$���f�������> CN�P��O�����d���x��u�шqƬ�XlxVHYEB     400     150��M動�x_/�j�t=���������X�,]�x*rJU�v��+��|x(��}�W���{�'���}���ڋhQ���/��KҐ`�(�����h�$�"���p'������W8��5�5��� �QB��x��{mErʙʹ��{���}��gTt�[y������;���-H�1��qY�����)^�s���]��,�<�P.'�x��e��|�}�9[C�F��UЛ�_��1��,���.�p�р/^lM���slE�<�G�=�L(��y�'͎�l҅��
7�� ��OA�<�J!��4���g�8�{7 3���&��(��i�XlxVHYEB     400     170�?x���N�MI{Q�#�rd'�Q�!
��a4
,3uK�X���]������:Hu|Q\��mN���r�P#R���ĕ�JEJ~	&��,�+pv�e�fr�|�ќv���"�C�B�ʥ��x]^�E��_~>B��!['����l�h:�APK��9� )`?W�ЧP�֊����[�^Df���p���H9j�-�"h�q3d�^�߳����0�?������_���g'G�Z��b5�"�06>�O�Ն�9�5��ǃ��a�(;��[q��ɰvd,b��C��`4�Gu�f���$�HN�OΞ�ˇ�ы�k��K��`$=R�����ʙD+9���4o�N�Ut*^K�x�p��!�J#XlxVHYEB     400     130�	���9���b����<A�.<t��>��a��aЍ���,>�ox��{�桕~xjJfd�ٻ��:<=�[����Ϋ���ۡك_����Ncښmeb\��*�0����Ǥ�I��Z�Ў����R#�JA�a��Bԯ�5�Ben1�?w-{�w�Y��v�-?&.��n��oHj���Z���mVy�Wې�/
�CK��ˢcTb���Q���[�s�"�y�z�w��V�������Πx�������;SF�p\�|`��)�)ş��APV֨�W���ڊ��Ģ��;�G�XlxVHYEB     400     100�Z��%іe�!���
ڞK���ܕŷ����*kG�����y
(���H=��l�0�:1U�y GMSTV�愰��5�Q���`Ykr����q��?x�8z����˛��2THֹ��M	�ߝ��$U`����z�W�Z�Bގ�'֕>�R5��z�V!C\-:S��7���ѫ�O_+�����vȄ�&��9c<c��"j60��~���$��[G�B���ئ3�]����F,
�����gfYUXlxVHYEB     400      e0le���M���M�"E����=4Z�m�����oL�×�t@t��5�,{V�~�^��9u�Ԁگ���F+g�=z!�����hgYAz����"0j���Y˯���Z@�nN94x4��%y�.Q7T� ��1����@��T
�R�d1E�o�E���F�\����b��(�~�$tM^����W���eRs��&ȩYb�����R�rC*����b�؊ҝ�v_wXlxVHYEB     400      d0�8uma��Yc�2߁���넞p8��5���Ķ�|}9']�>����
�?߱���!x�p� D�x�o�eG� �^�ž�X������':�:H9����&k-c#�����M�s[{�v}̌ov1�\���̀�����SzT%�3ԑ�&-��?Z��:���+���#]4e*�_C����|L:��>>T�����XlxVHYEB     400     120��� ��&��U�z��ϊ�T�2 Q��� ���djv"��l?UK���g-Xv
l�s�Y�"�\))W��z��~ap��p֒�WU�_U���k�5�<���� ���ge�h1]�91���xX i�M��齩m�e!~����=72��j$BI�]�D2��<Z�=2W��54�=�ר�����Ǫ���;ɣ�����������c��ͬ>O���0�-0T��7p�Dt�q"� ;)�2�����·�v�Oc�z�J;B�����.��B�K�Q���v-|�XlxVHYEB     400     180�i������A&��EC����ѯ'����ݍ��V+*[%������r%��+��H��w���c��LJ��+kw[��S�Ifc����]��N&������d�-_X��}��-e	gm�B�����x�C,7�������{��\CE�����v"�?+�f�B��ڣ�$A��Ȭ3�a�#�p��G�v���H�Ǿ�q�$|�լq�#j�5�ة�+0s������-�T�e�~D���[L��w�RG�!���|g��c����R��,ŗ�zr�� ��[_��Py�[{ go���H]�>B�W��q̈́��p�p�&�ۇ-d*���۹�}$D�IP����Z.�P�OTu��&da�T����J#R��XlxVHYEB     400     140]W	D9	�W^r�W?�bz��4��TA$�>������#���>.	���������M�^f���=R�铤$�&��V�+�uH=ε��I f�KSp���&V��FY��!��
�r��C���3��;'�(:1����쭊�1�fvmʬU�V����Ȩ��B��~�);0�!�I3l�<����QC�!����B
�p�t�D�����Ɖ�~��$Ty���'
��P|�e��eW�:D�~�S;+P�,w�0Ҧh,��������j�C�h��p���E{��O~�<4�����>	��,����y ��T���Qj}*���b XlxVHYEB     400     170V�3Ib��9�m�Y+s6�:�2��n�j�k��ER/���C�#-��c�xE}>�3�)lt'bN��*����v	+o3j�<�hWJ}SWK')���͋����#�T�ayR?��`k@�о!�k	?��+U�{���
}�tV�@�'��5l�`�=�徆T�7�.f�c}�ݳH �Zna)5c��-�=����57��(92QJh����ԝ���=C�"X<��NBL)�B���
y$#�G涭��F���R&mk14;a�6K��@ˇF��7���q���WLv>�Ф�V��HՋ�<
�D!�~���7������I�;����:�BNd��U�y�+��1's�`!d��YĖ���*D�XlxVHYEB     170      d0" <ռ�hIO���ݕ���LZ�H��r䳏�9|��n͌L��@�G��v�G���p����p�H5+^��X����_�ِ�.�d��[�Hr4n3��"���(`��e�!1dҁ���S���t-p��
H��bc�9�5;{�a�=�3Q�<� (c������ *�ؔzp�$���Y���(�����ubH��ݷW����0