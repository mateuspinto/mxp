XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ʆ$���A}'k�-��*�&�~3 l�#�jz
"�Y��D���|6��H�`�3�j J�m�W+\����W�Z S��+�9�o��t���j��
��cT�y"�"�ٹ=�v-�u4&Ɣ;��z��A�)�D���:/��9:��N|��?\3�p*�-ɋ����o�G�'�;/Iti��a2�]�U=bam,1$st�7�#ޗ��'� g����E���$$u��P�l�1�o�"��B�65>��7k����A�A���Ԙb�~�!?�w�.�7�"`)S�FS2��凢M��f��?*n{�i��#�ST"�v�1�J$�\.B�\�[�n�1�ފ��}����'�J=O��B轢"�Ј	�����h�\�#T�.�������H���� ��V�[j{d9����L]2���\f�^w���K�� ̈́� z�ȹ��~����q��56� <A;�&�[�t�_��ɂδ�t�]���+[�HH�����)X�͓j�B����%x����2Z\��tzb�f0��N��Ɍ[����{�l�d�b�=�\��EەT�F�ܔ^|˒~�&�|<����t$�E��nG��7X�D^�I�O+Hޙ?�w��*�u_�Z
���Q`��p2����o��,�1�H������rw�e�b�@�6ɴug�S���]{�GB���O�sw$	���|�0u��;��������l���G�O�M��� ��Hϟy]��Uj����z]"7=c�*�U�Hwd�i���vf)�h]���XlxVHYEB     400     1d0��9u�=�rT��&�DF�^U]`�9"�H�Z��������Z��R�V��0��O�t2b��0�����OoCZ\k��@�_�%'�C	�g�0,T���]���kf��4l9K�2���]¢{8��U�p(����4�V֐~���(��@c$����y� |L"3��6���ѭ�����_�$]������Q3��(CQ�Wg��En謘O�T���m?���]`!yOA��lN��@�c�Y�7��O��8��x��s��:Ä�9��,;<��I��SHW+�� >bvXy_�� V����+��
�0�"&%d���E�U���֌4vDd7�`1��94���z�I��8�.`��=p��/+B:ڸ�+w�A���N��	S;,~��ս+z�}�]��**���-ͳ1>ļ�������c�m�[�xN|ӄ����9�Q�<و��Ҳ���XlxVHYEB     400     140J��[�����;�6�I�^�����^(���-��:(���Њ�ߝ՘	��� #�!k�J�s�H���� mƎ��G8넄���ڝp���F�S,�0�C�7`@1FAc��0JēYz�:b�j�oqv���϶�#k��m�H1�^�b��ϓ��ی]񛽵�;SXE�����!��F����}��!��"o�b��]�{��iBe�~��R(����g7�SrX�2�E���v��Nڤ-^����b�s�:������g?\;1hu��R����2��V�S��i*���/�8�� �@�M�ȑjAV�̻XlxVHYEB     400     170�s",|�
��x]�p(�Hh���6���3���aF�Ƴ4�1����2��C9ZhW�V��N�_
<�ѺX���H|*M���𞪪�&���/��a�y4/�ON�2;�Ẽ��`V2ʥ�����M\�H��lT��!K����z�y�z*IBР�W�TO��WF�Q�:,o��tf��n���^#��ʙht��8#<S����e�$���x��eR�8;�fꂔ��ֵ.����ޅ��,�YQq�|;�)Y�b���S���*���g���K�G�28C��!�K�D�Jh7��P��1�h���B��	5����M��3���kC]�\n7�APLR���(q���f~K���9m�XlxVHYEB     400     140@f��<Ֆb��7)�<�g�G�Ɩ��!gß��$HAw�R:LEw;�%\�H����)�JD�?��#�V!��xS�RU�YoV�5��*-zcv�ߦ|1X�N'��.��j���-ǌ]η'�Ec�G7μR���_L��|m��-�����&��**0���=�rMK�y���\���	���]CC���KIE�[�{~����zW�*�V<f�����+&��?�X�>al�u`?��p�H�%�%W�a�M9� 9c$��RL�E;k�zѧL�W\�*M��L&>��+3��q%(C
d3���jXlxVHYEB     400     110�f2J�����ӓ�
J`���͋�{�Ī�.O�Z<Zr'T�>���Y���\���N�`2�Ezv:<�~��s������4���4�l���8�c�©�g�7{KZ�-	o���i7��]x89���`�[ȃ�&���5l�cp�Ro���4Q��5�|����ٗ>M[�qu��q�>J=�WF����DG+�/��[�0}T*uT{�0����#��
�Ӕ`ư{��TO����W�����%Ƃ����_��g����Y�r�˭�a,km�XlxVHYEB     400     120**F�$�J���]���ǅ�٬?@MI�Δ^ZIlR�����o=�R�_ex�֧���(֮�xy��$�$�n�~\`�%�t��H��c)��(#��Px��������	��Ǝ����%;[�_D~>1���'��'x����& t҂��w�/`�J����~׎u�_�� C^�n��oV�ǚAh$U���m?��'ۯZ��2.��L9��8t� K���+��7��;枯s�X#���[�e������H��o��4ًu������u[�XlxVHYEB     400     140{o7=�7��l�Y�\���x�N+�mG��{Y㮜rb4��-W˰aU����Rp<���h�|3��>�k�NZ��@t�ҳ��� ������Z �CK������˘��'bd�Pj#��M+w@�_Þ�&#�*�
.	��Ձ,(���P�}֓E�T1�����1��,�A�te
\�,y�StHV95�����{����3�ː�*�����̑����%��wk��6�'��:늕�+�*rF�e�� �{x<l�
Fdf�#�/gN&�%ء���?b΀�4�<�xw�]�k�6������
�p[4�N��B�,>lXlxVHYEB     400     150$�
��t�E��*<*2̾tW]�PoW+�(��߶�ҟ�b������Ȕi�pWw����0܎�}6���{�С�N�SP,�J<��[\$���SЙ�����Z� ޻�h��
��t����T7���-���t�oW��ٶ�BZ%/�ž�>�Ά��+v ���yZP��Vai[���Z7g~�T�,k��ZÍ텹�����8�U|�$J��3�Ok�R��ϭ1��D�n�M�#\rzFͤ�8�nUd=W�pݺE��
���  ��t�ŏY¥�c~ϐ��֦s��,�P��{H�cq���qqR8�@��%^y��r�VY�(r�����]��~$�6T���XlxVHYEB     400     140;<�l��'����~!A�v`���(..�G��į�7lS'~Xβ-��,a+��Y�s��c6�����
�꠱���$5�O@t��wu�L���������a4;;�^e�!��ɘ4���6��^���U�3���QK��+��,�6q6q�����"	}�T�ˌo�Lxo8q��{������],y�!+vU"���U!�889���yr�>��ZJ%�i#��}]�ٟ�\y�ߏ�'�0�o��sN�kÚ���`��@ ��	\��"���ɍ�X��܉m�5m�W����3�w�gF��}<�_�����+[Nu�wXlxVHYEB     400     100����K�\R��^n��;�R��L�A�Wg_�w�������Anm��暨X ���BVi�e��y8J�X����j(G�����w�L����g�6(���Gk���.�`'32^�O��f�>� :�or�8�`D���S��8'f� �d����9� ��*<�5@ 2<�"f�i���������D�O�`��#�7X�h��e��`�=Z@���ƀ�[���!�}ݮ�c����m?`a3ޭM}6Ǒ�XlxVHYEB     400      e0�$""�N�0�{���v�ɝ��%�u-��&+�tӑ���P��k�亹��0'�|!Žv%��2�����1)녋 ��U,��	���l�5L����ޠ�ѾV�O2qm��l��]�T�^g�����]ic�B;�|ׇ"���g �w1D$���=�a5F�0��D��g�	�g�|���h�ꇣcZ�4o�����,=]Y\���e���.lXlxVHYEB     400      e0{���Ų��`M�Q��g� z�jh�,��N�����m@j�]��ʱ~�Y�`x�f�𹺌d~dj���3�F��M�պ����H�pߒ�d:�� 
�
?n�6�^�!5�4\=����i���0��@>�"�( �f01�9X�=i5[��y�PdD�!��*������%�{�p~��eG�g/?y�ת_���Cg�:k9�Υ���G���Vkx��� 9v�?4AXlxVHYEB     400      e0:�C���2؀�Q��L_GD�0�~���A�r��}t����e���e�b�����X���7�t�V8j��F�K%E@�%�Z�̍��{�fiHC���gb�Ĺ�-Y���`�Q|-��m��5,��ƻ:���fּ���R{m�U�d���-�A�ڑ	�%�0�Oc��A+��3�s�	o��?��V`s�{j%Td�ܷ��u�j�VH�0�������b��EXlxVHYEB     400      e0W�R\\J����a�v�c�%h��\h�)�en�W�:2d��_�7$@G8�܉����#�T���s��7K�n4�;�@�_�MX�ɮ+���8v�8���凙��=]S���$9� �vV�A�-��s��: ��VI�-���rp卌jn="�������U;͚� �O��	�tVy��4��Q�W	�� �<ޕ��>|�"ڰ��v#@�["��$W�46��XlxVHYEB     400      e0l�O�#*!��y�Ю����@t�6�I���#�4�U�=X�|d�?$���/Ω�j��|�g�cX�� 4�'�?���g�P$v^����2�Û?6�#Y����/�V8T�
�8����@x9��S5Y�<F�v���� k�9Ѝ�옔�?kI������i ���o_qM�x�� a��*��a�:<09<�k�Mu*(zP���6��Dv9C+Ұk���dXlxVHYEB     400      e0}�"���X6Z5�e�˕�58@*w@d�T�K�L��9���"${����MԴ�ѧi���;��T���n���|G�f-�M�mi�]����<x@���R���x����<�L���r�9hv��m6,�kT5J�J��2~��[e
Gۓ�dK�H��)ܔ�=��yZ��W�t���N��2���L^Ai�^"~˛̝����)'7�,Md����,0�XlxVHYEB     400     1c0��pn+��U+\�lcF*hVa����edPbj8�,����Y�:�eӜ.��F9�M���~6f?�
팖{�)1�w_�n�r����<x.�2��=���*;��PX���e��:�}�I�ߞ�8n̑s��`��ܐ2�-�/Ft��~���9��u8�ө_���C
i& 2�؎Øb�A�cS�6'$j?ēW��U`�Q�v��pH%eKh�'MfzS����+��&�[Y������� 8Ч*��j5�o2��eq�EN�#�e~q�h.#�Yۉ=�$Z/H�ݠ1!cdvGݦ�pQn}4o��fk��ހ��%3�Պ���h:V�|��kw��mw3�O�/��2�Czs
�Mi�1߲��{�Hȋ�kE#����(IvY9�Fͥa.`�DG΁�ķ��QqJ�O�i�$�R�Mz�0o~LK��q�5y�CY?XlxVHYEB     400     130�T��@��:�S�<��%�pA�:��ű�=�<���b��r��e%����"�F��G�ڝ��.�Y��@���ވN�;x1���U���GҪ.�<�zN����Acz$��wj�¨ꯀ�C�	��Y��8K�Y���������`N^��?��Iz
m��lQ��;�ϰj�I6�+֜J�B�w�58��3����a��\��#�`�C�kE8�3Z�rgm�:��T*v���O��!���ޛ��g�N�h" �+����%]fkǰ_@�w�꣞�OƟN��i�~1,)�j�XlxVHYEB     400     1005Ӂ���L�k�k,��AHx�[|��A����^\���3851�\*��|���;!-�P���
+'%����-ė�8 �3�l:����V�Aҙ�~z7�՛V	o������o��'.���u��&j����)��WeĢ�W�[��YW(Y��^��C^��υ�7T�:8����Pc�\&$����~��yO�ƛ����'�n�ͭ�T��n��+�X)�g�(a���ct	E��Ȗ�	�y�l�XSAZm#�<��@,XlxVHYEB     400      f0ώ��s'Q������·|^Y�ˍ"qN�P�U�PtO�4D�Ab]�v�K���~����ʧ\2*�topP0�z�T1�;^�s�_O�,$�~�Q|�������G���M����1��}��x�=�d�g-��}2Op�Eg�k���(�2y(�EF�֓�zE�/qC��~�V��z��c0ɹ���ye�G����ѓ
�V����TkǾ��&��5ξXlxVHYEB     400     140��.e$iɬ=��%-0^k�������e�2���#�x�x����wz��^׌U�Y�(��IK�m���HX�n����jj<�<��[�K
%t/�P���]]��
['���ؠ����Ļ�Da��$����x+���ێ��l�@d���j��׉��1+�2�v@�����6�ǁ�Z�] �(3Y7e�ɵ�L ��>��O\X�!����!��.r|��2�h�3w;��#�k�.�k�8�5UMe�I)Jz�����Lfg�향P�.��{d����F���ڄ_�%�}Ĥ�Ǣ��bi�.��GOa�TXlxVHYEB     400     150;1�+��߽��߼�R2��������Yy�y���](nMҗ��Տ߻g��h�L�F�qX�?�c}�[b�~�ߠS�~�LL���g�96ݚ �~J�7XK���w�������߂e����$ms81en7�-p����Y�$!{���*SX��;�\��Pnp#�RF���U'U�h�h�3���m�h�d�t��R˩7�2KөiL�pfZ��3�|�'�I���TE���ǔ6j�4y;���W�����8��c�UF4C�$�ͩ�#��r�e�"�MjǦB��,��������Q����_}㫐&R#灣2D;��c*�H~�+�!XlxVHYEB     400     170G�2�y��@��S1B`$ E�5`��M�T3{����Is��׻��~�D,ȏpr��}lQ߿<���05,�g�+-�(�����Y��a��Ǧ��!-�JP뮦[W�&*�y1���O�:��}�@AC�k����]�Z����:��&���+!��7ʸi�U�4	�J�����y��Z]žʐ�����H�OoC�[�{+�u_�6zı�=��4�����C������������_ogt�mo����	J쿲f��au�X�b|��z��Oz&� ߖ��U�jV
C"}*3������RV�.6y�Yu�ϾT<7�	�U�[�@)�/~gP
�Ə�!WoB�� �eē�"���n%^�k�HIOXlxVHYEB     400     160�kZ�;�-'6eHD��?r�n�N�r�4��P�1z9��?���I�FBU��:,�X6!x�S7F�h)���#j�MD�����X�S�(�V�bp��>±#H��c%��?��O�d|��Dc C�.�P��υ5g&]�5!�C[�#=p$C^k�1+�d�n곫k�^n�<\��!�yY��9:j�(���ܴu���k��1s�5rX���¬̠����F���+��~DC^�D�������l�H�+P饖����ݰ7�e�dة��BLe  BMKS,��	�ӌ��4ˮG��=5>�������lhp��O�?���A�d�`�����k�&��ٺ����2�"�_��4��XlxVHYEB     400     180��ќ �-�>��:Z�����u9�,�b7�e���P�CkU\}�ޚ%4f����rWm"��������y��e�c)�4y%����`[��5�<��<�V!	�ݯ�X7S~���I2
��oGF�@�c5�![�C�-��Z�Ȅ 0��%Q�	�ZͺW�_S%8�%a�,!C	���K���y9�IGnb�X�y*�:�5�j4N2�F�,x�D�F��v�oVM���n��%���Q��f+[-Ldb�9+>��[]/ؖ��B1��җ#F����,?>��%#h����g�04���m�a�`F�h�zU�,�|��	��UO)��s��d�o߸j` *\�1i��p E>�C(f�|��RW��#t�;�1$�#4�6
�h�CXlxVHYEB     400     100oxU{%^?SXvPGzKGaW�� h>�]��i����:U���fZ���8�g�<;��B���g��ϲί��?��׺r�o{�ƫJhz��>50;@+ض�g0&�Щ9b1��\��/��& tt�)S�Z<�di4������;e�23���I@D�]�?��1�d� �B���;FD;���Z���c�)/¡',YL �f?� و�J��ȫ#F�KU��+�8�'9�:���fZ�ENz$��0��rj�B��>O����Q%�����XlxVHYEB     400     160ߠ�(�@SZ�PReӛ���!��ŴI���\��c6,�@�6~��0~�9ܕO.��D�*L,Lfggs�)�m���T `�>!ÙJݏ@�.4�7%R��Q5�8�e]�.n��&�-G����<��<�7O	��� B$�/!�O���d�R�<��V��\^S������b��{��ܝ�t���Y������+Td*��Y�w?ɡi�Wo������ޙ�/�V���*�:d��|g7��r*���:�}�J#���C�~؉f�Q ��;ik�	#A&��lq���C(�c�[�����y"ͼ?<q�㾰�;H�tS�=1r�:}�]���&5�>Y5 �?����iф�0:��]�ɾ�XHk�.WĔXlxVHYEB     400     160+�}D˶�!��W������r(���������@Hxh�#���>�A>��~�+�n���B��B#��c�=߮��x��ر�g擾/��RC��*���T�k"�6+3�G�
&���?���1�ٷU����y�S�J˝gT��O���d�C\�XÓ*�&jLn�(�
|X0~�C��n�j��VW_{.����eI�^���s\9QJ�A����C�Аv�MS�x�%
���Sj�8I�w��*��������O=������w���<�Чn��l�=+�Ky�����o�X�ƥ���o �{�J�ȫS$g���{0���qE4Q�o���ņ�[XlxVHYEB     400     140��H����>�)B�j�SXl���r���>д&\��J�y/����[缑�Tq=����(T��Z�q���ASfđX�`N�#!Js��x��b3��5��Ƙ��6�p n}i�N4p�`��]��M��d��J���?/{�4�J8Lw5TE��A�O�'s�to���@8� 6;w�����ip�N[y�~��� >[,"����c|1݁�i�n9��X���#0ɷe�o�H���>�}�8�_yU�f���%�g�e�UM��0'��ɒi���a%��9h [���Ŗq�B���1&��Bq���0�E�Da�8�لmU,XlxVHYEB     400     180)!(5���,I破�?3l��-	�r"��C����:9�;�a����q
l����O�,�����c0Aڴ9"����|:��"1n�x#lD����1�6���/L��L���uzw4�VH�䢍EpX�Ʈ\�؟��ʗ]��ɸ�L�[Έ���rߡ3�7�WM	���e�$��s3(<TͿ���$�mnl�;�㭈��S>��t��%u
�_2��`��'����NO(X����� p�x�2�v)��k�2(N���5���h((j�Û^��aTYk8��0���+d�,uZ�uA���<-�w�ɷ�H���U������[
��$D-j�����0<��+M�F��<����[܀���_�׼!�&�\w��(�lx8r��M�N�j�k;XlxVHYEB     400     140��]ߒ����C/N���y�f���'Iu@�0\�Ib�d�^���*F�����9MbD!>S�%�m�iLagn�O������7���g�C��pVc��- O:R��y��@HIM:zk2�Dq���*�eD�$a�}p�R-�j�h�gӮ�O�X\V���˪H�����h�S�?� �*|*.8�d\p�/�߯���S�ڴ�������E�D���g�,�s�ۚ��]#.Or7?�]��p�s��9�{;�/:��RlRGD�lle5%@�~��F�-&xI̘��_�U|�\)�d��˄6��`�Eϲ���h�Xh�XlxVHYEB     400     140g��6=�4�]J0�yh>r�ќ!;�9yp���~�򚻤pH��ӽ4x#�WL��.�ө�ز�]/Q�U��Rn�v�f�Y8�E�w�|&�B-�/2�+Zg+nIW�d.q%;�K<�vԽ���8�Ű�j�ǒ𨑫Ģh&U�+�vھ�'�R �5u��U���,�y�zF�&��+�s�y� #�Fh���=a�#s|����-ӫ�!���f�� ҕ�c!zJ���v��J�B�������r8����\���UN8r�i{���5��!���q��&j~�nK��ѣ�9bW|G���ȏܝ���1��XlxVHYEB     400     130M�9��v6�Y¢�N���\*x�;��UR= �!�GfZ���ΗYydqo���>S���y$(}����������^0$g�u�s�+��"M%5wSe�����IM�:�#?wo5�o����3Mjb���S�.;^v�n�P���I�d��2L�a+��>��r�$�O�j�5��<z-O����2R�v��G�p���0,�a5��T��4h�&�]4/D)�0rs/gzL�?̍�թ�p�ժ/�?:��.�r��x�ʤ���4ew^����Y	�}�ĎG�WϮ�F�����XlxVHYEB     400     170s�[�`^���΁0�{DDF\���W��`�̼_��1�+X�و�>�.�����\eg�kF�$�9Ys)���Ϡ���@�1���6g��"&���8=�������j�_.��<��X�1$݈G0�I��s5sc�/�z�A�AZ�Ƨ��0�'!������2J-n��� �*w~l*&��s*�<Qn�x p���P���bWw:�z��X�+뭰��Ҁ7�d���椤��fE�X��;I
�6c��������B�-�Di���w�"��-���Z��~�8���_]�e�m���5�N�0�Mn9h�0h��;��q��ҨJ�m��<�l�Qmw9�եi�n��ӿ��[9�m�x�
7 �btl�XlxVHYEB     400     170�C��j^XJ<��x��<ӑ�DlJ�q�@C��uSD�z�Em���2Mß]If&�R��ȉ����0M��ݖsoQk�����^��A�Ga�"]�`~��mjj+��b����x��G0�d���@_d@�~r�X��\F>��u�����w=�����!�L����>��9ʘ4f`gv�X��%�'IL�[[��j��I�3�	��-�eC s�� �ȭ[ˑ0[��'����fm�n*6�4_�:�D&:�`�����jf���L�KU FApw"������)6�D�Ÿ�� �*v���`�DqR��؎��+���|�#K��B�����RP���cO�G�/�CT&����j���}�;<jXXlxVHYEB     400     190MW���~mIB:���<A�떣�Ęz����W���3	��_�A|"��* ��Lt���Յ�\�O�.fZ�!cc-8hI&��=���j�}WMA�� u�����t��,�B�j�����0�p,�U�	���N<'����\v�M�܃V��W�3�}�� 5��2���. ���RW�i}��O��j|�rM:�Q6�	[J/ �o�"��ذ6�>0�+�kN�2(\�e#���B
ù��`D��	9�mf�:�I�R=X�(��ɟ�" .���o�W��F{���<�������VV_F�R�gj�4��������D<,�y�Dr�alDt#3-��K-�'V¥��o��.���R#�ie�=���=Кȼ��ۋU������XlxVHYEB     400     150�P%��.�B�|W/�P��`L��ۜ.Jk�9�Xuw����_�[���~a6��B�yt���<d������Y#�������$9Z��/=�mp��:XP�E��~����t�=U
jw\�e��������Q�5��� ϒ�
��P)����-b��,3�،O������ǜ_ü;V���9��UM2B�"�#S���O�O��L�wع����V����: x����L0Kٵ����E��m�>X�wNz��,١T�EG���ȼ�b���!�������F ��*�(C�-����mS�C�%�8��ю$s�Sbf�)/�XlxVHYEB     400     150W#�˂�_x��~U�7/[���B� ������N��C��,��KpC�k�Q,�>}����3G��PE�K�����M����#��P������	奠�AM�W��ю�`����8Sb�CyFv�Ѹޱ�	Zo[��q�w̼�k �ŋ]�Ş�笌]wQ��2�i)q�f�@	��_�\��L����B�Gm3��F�z��h2_h�h���0�\p�;5�g�W�c��Lha��A�M��9�uZ�}[~��2����R쾓��H�mK��*'�4��	�AD��)�f�Y?�F��"ZI��;@�s��:��K�l�0m���_7�(-�HzXlxVHYEB     400     160MP���;y>>dv?��������`D�3����opb�&��AS�e�NԿ�V�E�y�P�y�zq�Ӭ���c�k��� ;x,����j4�?������ˑ��O���<R�;�v���\2� ��s��x�S*�d��u���H%u9��}�����0&�?����rIq�K����_�ƪ�nG���P���ɵrW`.� _B}Po�i�e�jX�搼ժ͌ �7���c7��h|��s��+R��E?�;@��������؆r!���C�pb
+y��3iâ1������n3�+z��\Q���a�\�eWcP#�ė�+�{�����N�bu�3$>gF����zc�:�XlxVHYEB     400     140'���_��S���}v:���|l#(��K4��6K�f���il���Nq�j��R�d���n+oZؘp��l��JZ' vA��؇�ȩI�Ir2�KoP�a	�|��@�s�Ih��y[u�,�7����M�:�yՈ��ʷ�C�H�䰗>���0;O���H6����`L�͆ ��Y��rn)f�׃�l۷\��ZSSr�݄��)f|��.��v��	���:|��-°&�"BC	�.��CF9jΣU��N��~��cE1�E���F�')�AR�Q����=# �w]��~����z��>�x���O	��" \�kXlxVHYEB     400     170��w:�X�����%�_�y�\x?���}��[���Aa6��Ī_�D���#iQ�]Md5-�4��?`�EY.mB�#!	�S��p@���\򼅃z�~�v"��u�#�"y:ǲ��8O���n(�o����Xy��Ÿ�칧n����
 V�meNQ�b���pN� �S�B�.�����.�'��뿑�R���F%�Ȳ�������#�l��Xu�O�Ym9BK	�E�~�_�^� ��d�P\[f�b�����.�p	���G�^ti��+>n똸{�?e�xhT���o�u�K�a>p��f{/Cyk�h�s|�=�]4����Qb,�@������gהR�Ğ��0i��i����S=t�XlxVHYEB     400     150vd�����I^8N&�J�#���Y<���rq���$h���7�G�egx�溝/ ?�ТI�/�&�3<H������p��t���?,�ї'-w�u62p8���0s�i���|��(,4�ԟ�i�&+�u��}�����-�J��b�y:��u�-��־���^+��
K'�M���a����m<�p�W��DޥF�\Y�l��/nhX�A�G6��^}m���>���"�7+P�8eJlǁ�|\_��ݝ�]'V=)�F�AR�dR�#�X��U�����8w!�ߖE�M��=țݮu��;����Eܜ[�X[O���^�$o�٥��YrXlxVHYEB     400     110��F K�J�$*��^��.�n2�wW��ͨ�����rs�bPj�ī�|�71��Ԥ2�aIo�.�q$��.$���	�����\b[ELz����(d�&kjd�j.�;�f�:��@�[�D�����_|��x7�=�$��ϋ��Ѧ,n�>} �6�_���<��r�c�)n��+����9����P���RR �N�����ׄ(~��,|M�S鋺�Wj��O�s�����������}O,OD1�Iå�N	�ڀt��Nf瀑���^�0��XlxVHYEB     400     150���s�2S��(e'��UH�o�}x��R�i�~�`_�ڗ���O�P���:s��d�i�(��}��Ma�{vϘ)��T.i�6�_ň�����ć6o<,2��#��zW|��l��N�Q$���\��Aj�KmÊ�	X+�e�@���R��B�^����"ܻ�#��m�.>wx�/70��y)s����t��fa)d��`t�+�<|J+rT¤&�D�(�����X#T���.Qϲb�IW������Y���d\B"�z�(�,� �1m�\1+\-m�Ι��}�T#���v�zf�@��7�刡d�vly@���ڹ5���
�|��طXlxVHYEB     400     1a0�"K�_��+)�?3Ǹ�	��17�����q����x�0�Yl�l��j�����o3}"bwj~ܟu�[�����J!5�R9��z�|n�2��o{��u2�'����P��w�C(���	���ba�}m���cY�����fԩ��(�Gĵ��8�Elc���0��z���O冀p�@��IDV�P�(D겠F�%�R���Ad�]95�9�NxA��
'z�I�D���(S�6k�%޸E;�A�Qs���2ah���Q�� r�П%ě����r�f������r��!i��{�������'�C����&�P8��<OPW
�>�'��7��p��#	��Ps�T��3,n��xH�`-oGt���"A��$�~@Q�3^²'��;;�ѱ0���5�%�i���pXlxVHYEB     400     130��wR��޾

B��;��B��fΝRe+��c�;����Se��2�M��1u,�L�3]Ϯ��~.Y9Vh@�.{i�"T�07Y��,N��	2=d;5�Ց�
�mJ\�;�ܫ��T�8����nl�W��o���ԡ�#ib���b�ut����>�:d��c��!w+�{��uV���Hܫ����k����d�'���Њ1�?߼��L9��<��N���O&عl`ĵ�n2��pa}��	��b�
�΋}35X�N�ν$:��}��b4�wM��b��g��Ů�˥ˊ�9,DXlxVHYEB     400     120B��A� +���N[1o�%�o(�o/q�F~w�?xjď,W�z����m��kZ�`qVX�?_�� �L
���G��B��}���m&c�fa�w��<<ʃ�[c�d^���W�ͬ�E���X#��s���qr�����f�����lԌ�������v,e�0����:`���1�1Rϯ��
.���N�,z��Rf���5tB�(H�~���2Zh;��5��B�z���0U��m
i���3��zp}�װ� �f�`�K���[��o��M�F��V6�h��XlxVHYEB     400     170_�����x��� t���szk/_�y�G�Ǻ�i:g<��!�*�s7ܒN���<vbÿ���^�N�~��jjV.$�4���V����ip1!�����| ��Y\g�0{p��b�kx�0��me�~p�H*�+�FN)�G�����d����֡h�/��7��B=&~C�A"���ԟk���T^R*F-�G8=�8���^��W0���=��iM�w%�|�u�����o��������kO�n ��j��B"��O� ���ߤ���J�>������WAQn)O���R��ԶQc�F��>L4Y��c��9y8~��	�)���m�s"*67Av�2?�6��r����G��sy�c�XlxVHYEB     400     160�3.��1ۆ�C�O�^���XN���@�b�!��yR�/W��f��P�0ş6��(��хM%(2��QU�8�O�G���ً�(�mB��h��y��/����sj&��$"�29�{�JR������ֹ�P��k�b�Y�%�����mA	�ӹl�_1νʹ�4�f�x�J=���x �MQUTZ�NOfR;؉h�й�&�lK�F���<��/o�@���}~d���r��EO�Gp3l	ia��hH
{=*�%�,���/��ݡ�E�W���6���ޕ!� �]ȃ
���c���}�:E&Ku�dBa�ﴟ��u��f/�V�<�c��]��^�9i(��Qv8���e�F�4�XlxVHYEB     206      e0u^��4{@���T�\��0c�M�e@u�����:F��lw�|�B�'��y�R��G�>	��M�s8_�rK��,�tN�ke��6P����r'	����O:P��pܓ8����O���,{3Z$=[Eݾ@��I��<.�+���b�w�a�)IWdȞ�zB.X}U�w�1$lZ���!��;�F���x��L̟0{�I�zu*F�@�W�ew��M�_����OW�