`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
K3B6Jo4RtReNN66yjHx/LX6IUcH+N/hSEXgh3EdTlkP0DBEmVRNBdextc1jxAkhqn1o8Rj66qFcY
BxYa4lFAXAsDWLm6WfvrfEaQWzqR7XhztSTAIZ3tDNNnWqfhnH6kA8lhzc75f4pl0GxVW+4dA9Kx
KO2NViV74/t30kAVmRmGTHGjRVWBxcdLIdmIAfRqVDTobqaGoGsLiKZY3lne43JXImkt5LPhMJMu
7HH0l0zLha9XoJ4J9M5KGeZi54UPhBlK2UlrvH/ZlaBHqDBfbwtcIi8yVHY/R076D7FtXCwxy8+K
lW3RBbsPphyQu9KujXiG7SQvNOVY9GSF/j/ACA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="7U0v77SBgzhRYYMeg3Z3m7MbdGflyb2GMiyHlVM5B6Q="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14864)
`protect data_block
Fc7CftjaXQTK4jOhjGI/IYySx0gcodbyUtsLUOLx2F4Tv6077xLOCPYIyHXvoZjGbyZ0zSvUTBRX
nrAdI0EQLSZVQWErnO1YxtYo0lQCGAJKCjnBKwMO69vDmuvmLTio8cYRrONb5dgO3Fwwk2A8lt/b
tKACtx5gbPQtHavl+/VTIPI7p/QCTM9A2sQDlM/CJCHqk1XYFvW96ABXy2/ucGdH2u1UZcMpPUC4
ri/APw3w34cErvoY8aJwu34PPQtnBfIb+JkkT8Sd8VgN0wD0qbK7EiuffMK1g3ui3rFvLnGvh+wf
3xYmBgF6Qn1PyswYEY3bPg8uZGQ/PpUDzzo5/PYgG0+NM4g+VBz6JjF+Lz0RGyz1hDP5Wkv37+fQ
kq2hrDSEdhVoagUxDMzATE80+J6LuB5n1+/OHvaqzw88jxBzBn8KU+KU/IHG73C05xN6EopeexSM
G+rWwV25QTwc+nHN8VOK3LKXerZCXq5bJl6zxqc0b1n6eGhjkE4a2Cn+JhZphKW9vaFTzR5k9cK/
uQhDIeG84VYnMgtRXdVZPN+04M5PUXtzgCiXoOmf6BB730n96gflBXLW2BP0Igst6UlE0nC8YJ9T
THA0tft0TW9Rn7KuDiS0eUAdlvPIXFemWPT/9yI9ieVnTe+Fof5I/YG4CBH+aMjnAp7LLORkbMsm
AGHlhtbUXV58/DGTJPLD4efgSHLKhTEPfMQfZknI0m5nY0veZbkUI9VIicX9ml3zJ2yRgihcCXq7
6qQYNEAqLsvbkpcgSayxfu4acIty8qIBzriUDWsntbOxL4Wuo9Qf40iK8gL4EbG/E8GxbZqLDdNz
Uopp1IUZIVz1OMq0D3yC3VLpgCcFDxrzxM32wBB8efa+OHKw5H2bKu+mDP2BTesLz0ojdv2X6x1r
pFHAomfeolQwGIzlDQV4HNvdixDu3wcsim1vQ87GwI5vcvsVC9bF3nfDlcJXRjWaAJXuZFS5YG5u
GTaRZPAAiS1Sy+xEh3qjM3MGpk60Iu5aU7X0MTPkP5mPq1OIaj+8XYbJpWut9NpfGHgyb3j4Yk5G
l7a259f6d63aecG+ad2GVgLnl92JNldZ5lAu2nPWNef/vnGMabUx4WgvbThK40D7f2FbVWdU32R1
Od8Bq6IVYWNlQritgAqsz5Rle8fPXaxKI7RbZrdQ4Ywq2uLqEhjxiveNuzuCBY16pTa/H507bZvt
AHdco4RT3mMzrAwB2z79vxWvG23oNASDb4Nc23i5kYqcdQlFSQSgQlrQ6erw/Xjy/njcv9uY30Hv
TVJuhHno7D5sS/ko8WJ7sy64Rz8HK1hN9bw3yEeVUeQAmxP2Wk8pMVj3QxgY0IY6463Mz8sbtWg3
djXoS4ZgHczPjvHVdeMgsC2B8UqpF4qcgXZyfhZZf7jHr2FOLZXng8xTDDl/3bYRkM7u0L5d+tjP
32sjrKYRG5Lc7tW25pP0ruNR52wkSGIOAbfInS7+FpIXYDSDYumWAiSJcVNMXKJh0tmGe/wdoNhR
x1bsOnZEWGTDBw+ojVjvI3e+0jW8htEi2bKRQixof0kVa53RYT4Qgl/YRk/tuYSppEsfHgj/Yv/M
WbHIprHGVzU0ixm1UejOUBxrX6hhbWMhJ6ca0CVhJEfPNtvF5nE5QkjGGyLqFKXYnpws9StpVu0t
HsvJ5wSeCnllv4/91+ShsD8GMSII5YNl0ZC0XIpD2hcWqmRks7I1DtOk4/4Ha4lLgBkjhlT9RhBF
xdLxEEh/ETpMsV2jyy3NHfLobFMwTQmW3FKEJ09i4D0db4vEssWTiCp/iDYoQyRhr3MjJsIBPo7u
n9zFlIKynM0syyJqGvOCK6eHcJORwgl3/7Qkq6FNr1kVrkwraRr+HNt7vceTP6Bf0P7bMpl9nSrq
Q5pobFX449KgzxpMoNLX6Cci1gZW/I8Nd+bI9ERvVdMQsCYuXtbOw8WnbcaHaRAujs4G/WatwpeF
ctm0jt6krfz3J5cSPnXdC7q6471HD7+/2uqSsB0y1KESaJHYNs4oyvd6J4SCp8/7xpd96+dCB5ha
PJZzVgPK1qwPwZtTkUWe7ux62E1mSddwClFKJvf6XftE8xhGj2vvMvbGlxoeDLA+XJ/l60plW32D
hZMndkzKkrN9ikVhmGtLW/TWRm/xLLnhY2PmhjMJi6YN1n6Ymp6xNJMyi6+vaWEe00IsgO04nEJx
LkU/pT03d+IetGU445sWvzgQbEBR99/UoRQPmlsXdS2+of9sS3ZLSm/UbSA9g8X2rfb8rVaKGWnu
Ss96ZA8tbswkB5iig0fDpMS/A8RbYloS4RKmCxKqb6O1T7dU4QyrbJdkrcqXKwZV4vIU/AIQCv9L
8wnpYOIgVRQ+qZBnMknVlg9bYJo6GX0HRcfU20Dv1cwQqaByj4Oh+Nfb4oZwJmNV2bJyZlLivjN7
apyzXF7iROr/vLiOEkofhNsxG4I2iqzCUxPU5ZNPUb2Ffmc3wtbJnCsgZGL1r035/5m/YGp9/u0R
lurSeXFHBG58KVUjxHJsvcyh7pOYimFWX6xbNlgAk9t2GEQKdzNGFYucdHyQPBjJwnOt9+SB6Ofh
mpcG1KibMUt1PLGMwhPgeUwbIxucNHGbiXRNMVRN2vVR+ZYkeG/6vQ/Z7fQ+/zjI66CsQGXGgx3v
VrTs9V918D6mQlmryK8poUaiKKru7lt1q0BORYgJdlkKhY03WBMwPgjv0XJAwCXnNFERAzBgbHMr
H7JiaAAeM8HkUc830qrIwaMmX6cLx43leGdNKWQMCj56obKVqOtn/TKcqN3JVAOgUfXSNuePjrUb
aFRNJtUxzQai70eKqe9ghuCkHG++6yvpFG41a3c84lYLUC8tNR/lSIWcrEWpsn0hsFhDtsmZWIUO
OMOIaf35y9VM5UfshngwqSugoUL0y4+kagyrwQjuRark0MIo0GfcMPGEIKZgphKm1iP47q4CtIHH
BGB8ta+R/e83Mbk/4BTzHH+ngY6WKXf4//yB/V+ElFg6U3QA4kDXEcLaq8EZg2q+Nz+CLJGc5glE
6IegyO6+m+9pcKyMTSYBc+vD9FLyKA2o9qZcIwPBvebT4ajGsOMxdMOWxuNrcckVKhr77DQUEv1h
mMdeJwQCZgrwpa0PaIQYAm3VXXCllhN4YYgF4HtHgk/MKmWvj6YqcwVITzWokoU7f2Q/tz2kWQ1z
bxcbxI+6OuC3URcMNQzQhL40N/HL6rD5eoOauTSXNVFqB3de6Yj1dwRi61T2IxibFh1gpHlGIwEx
z0ccSa4oucc5AxGlTsPpMVenNm7NEtgM5rlzcEwJ2nDMBhcyIULQnQKDNVaCXh9Z784m/vJb5dFV
Uh6+YQubWwcOPzcO2Wfars05HR461Dyh4oWYTwGUSA0anQA3GdlzJXEvg7lFopAf7B/ezUrKGA1F
XHopEVo+5hX8Ae03cK1/AQC3vycZkrpS3eIUVBXPLgQ1neK6Fh64L4T+CDm5nbb5AjESu7bM4yOL
OWA/vMS0NiiKfw5Ebr2mDrFoMlwkrcQ0xATfTkuVGjFmPG8D1EXsWLYmTY6UruPou36Myh7aURIj
fNrBDTUHvtalH1A/zwyfMIJlGFpXaGZMU8Oj/q3DPinyl+4qTCVqC4bJIrDWUdTwAnqlZSna++vC
7rd2DfJVUIvkqsl3nOEpyC6ZGgaAO4GLamybRMzrCVZQ6NefULloFdAPPzKmeqyKt9RZ0AWv+EOq
9KaFaR1JnyCyy+MneyMn9Do4J6hL7uLylmVOOU4ahVOfjFP6X+klRa0SxamtQCvDez9MEEhcznSq
Xtjy3BfTysgFYtR3SuUpRxMb3MKLlmXhqIRD//BLmU+niVqjbe9V5c9bX0PofVuJzmIQHmnzA5VT
90dENF5h/NhGz7Dd7fGfGXkXJUHyA/CG06FIZCKu7ug5p/IDb/0xaU9k4kFRVDiUYh9AxQJZqG50
f6tTI9L8UkokvrhAS44mY7T1f5r+M5mFANsTyzh/wS00BH5zN/yF7VUfiAH6LmFZ8k61eBW6j9iM
cnyy+GBiU3yDTqtYGABriNet91IMlKo+FJYANvqe1AhZ5hzmXACB6cNiBV75pGjn85WW8qFcjr8z
ibWyhE1IGwOHMh6CfYumXgB/H2zLyOwESVUDJvavTcxaLmSUUUn/o0csOBrcpV5nxc+QaGRUjQJH
QrUGylZ5q1lfK1YOFUCKsevQwNaD0rQAy8/JMVpZhU1Uah4p1th+vsm0yEag9uiHO3sRDEiadLUx
BkWs6AomXGRQ9Qz5mwytTB9QR4a5v+NO5F+7RbBReg1IeogwElfDkMe/xHxm2MQ4Wfh/dJL794bQ
yu87ghGy0eOnMeq1AwP9Iu7srH7FRG6vYHIjFtTzq3pPkwHdid9RPbtrND8sqjMlQwGJbB+aIiVt
75NanSZyIa/ZVCUGi+tEHR0n8puIsArlNupowjWxxXqEwrht3gXyDfK6HStssmJkSeUrGVOMziHe
2knjD9FXVpnzDKeWjKzJ4aHYBZ0EAlQiWqVRCrLiU+yi6l77DarCapJ4riVDdxNXySHKamWwgwu+
oNi4MP3qWZBHin2kJYp7w3Vyta8N5+mu51q/1nmW+L7zD1MDfJKS5TXNo4M8vW4TduIjJLNPXIql
QpNxI+wSRYOEfhhMggnwgsAGLrAPachIbi4oyQotqKC9aEKVuRuUNUlEgPgLsPBh/T/I5tP5JFIL
wZiSJnfBbiUrdWmSB3/4A5G2YY1n+neUr9wpXj+OE2DGUUkjHxCCPc3vj7HYQTIZQYu6TjYfZ9A0
7gtv6vBVTKXANmrYzVWvoCGlD5y3vRlDsysf+bPiLqxruItoyDenxt3J2f83b1OpYR1PuLdXsl2W
HRJuhP2SoL0m4ySTY2MJ+5oZNFfDhD10nCM/YlgJKwK9B0q2P6VVHZus1d2lXnoAmEaj8nKVmWR+
wo1Ups2Z/7BAGowyvt52xtFPl9SsWZ3iYcErjaqhtDuhblRi5chds0wDzTlhdQPzxKovoKS+0iys
SPycY7QK7lq4/G8PxpwsiZFpcxyKnLOx+DMHCxf5c58O4ZB+sZ5PdU398IrvPxcK6OChS7bePDJS
eJJ2/GMS+qk0epoNBi41fxymKxy9PJuI3mfUmYNux3NrcqiMUMtcKzwkTFfL3jX6BYBPDL54tu6a
JeUDISYFppriY8iNA1eOWgKzBiDi7VE2MZUfxUUKxNN+JBk9bBK7jWXvGGqAlqsULLlvePdP+ofM
j2syT7pWpG31ahkh+ZfGTAgfJhXIGh0ljNlypMJs2WAVjwbZ+wEDMVoK7AbnN4JzvR32jfKeCh0H
579pxQ+C9MTng0Y6OHYFn/Rizfefoa2/rJfjc7YW1tXOIeo7Y8jHmFxKqGYBNrE6n+ofXRiQu1NG
rBxqa0DUmz+l8aX39wQP/Xy68J+eB9n4t2vEA5J7byC7708ie2NRUtE2lVEfGVD9+QIcXY4Sp4xs
2fn0eYJ4StMYqXmc9BDrfmHsUWhxeIKA3IHhe8IbK0oGJ45Xl4RLPEUxS2LLz0Wp8MnLPNqwTNIE
yJyqd9nGde5T4HkXD3In+DKyxaMDNMY25U/EXCiSSgsj2qdNnaGpsFTlkCLqQKpQZf2FAthnKe4J
Vdj0bC5C1Jzw+biYUtrqiHPk9oToYe2vzXXJzGVEUoh3Vsgn0a7lMrEATD9uZd+1lSDl66hYdbpX
PHdP/mJ4BuKUZQY+BoIkQNFalspIARvW9efHZoJiYmgd+RGYM66kdqpIBuUnM0tGRehlWKd18CZ3
/PdxRMRppWvJQLnRI/bxmcEjM6vY6cOFZYUGW8/OCstEJU5gQ5Psaez3s1Y2pkfjmVjvD7XN0dvm
dc2f2dGVKqmG4SrsCUNSpKqEACqAuO3PaR6zIY12g5Y+Pvx0yyoMJrG9A77OFdaFyxOOO7xAKD+R
mdfWb4IFhz8j/a5szXeejgXcqDVlp7jAFtQhcy31UPRvhnMaJRoHJvGNLESbuCuPEdD2SS2q/0g3
I2wEWaWWUVa3FIT7o6pX/GP/fViXNfWVpM3UWMBeXq3yyQz1hfRvcN+VlRzLFuiiDkPNVfzGyMX3
8vlLSM8A9i96b33UndWDhk/DxuBXwIBNFt5d1huNftaf34H8FD7/CJAqjn4AJX9pi/3V8uTJbG0P
MthtwT/5e4HM+/KPc+JwO2l1wOCEDCg5ijL4xfJ5yji720FjPskbXa9nfRQa8AnFozwtsCWMNJaA
iBvWOMxO78mBHoZmWrGlxiBi9/CHNp9Oh8G16hZKNQdFDSYvzd12ThiLm818TgFyHGNxgK7949ri
VrwNxB3nUXH678RHH7MhUWal7d5Rbx+ytuuc8TI7AUU7aEVP6krVrWDn00NvRsYvXKWMeI0+Ij1e
p0TMEwl7VfDSdAjHk38LPGY/AlrMZ4ttpW31TVNq0BQocCZS0OxYeZ2X0lVla0+6VojTWRwqKlv5
zKeWW4BgJcMbkcsOMcjih7kfXAxR08BKd77TXGbfizKnYg4HfrUbpjXIaJMbum76Fh0NNVC/zT2F
Bwmr0HjYvBMySt/R4jzbUHWB1BKbc4VWMRFM1rCIneBsikHHpmlW9vN96nr09iHr2PeF+pm9/8Ax
r+D7ozkR1gvc/qw/KDhNBjSs6VSrmXW1BabrHFjd78RqE0XwUmtbi3qOGIj5RrJM07rqgmPoIO5K
u/o49gan62yH488s4d7ljw1S/YKQsJMMlKssuN3pnjFSJcwgNKmc8W6TwIfArevO7TUdlLY1bl+f
Q1LbXds36bUiQkHTuRByoOOpmpF7RBUENEA8/77qWBJFMkIN/dLbifNMOTBa1CIkb2O6KiCGsgw7
coxHG2MKHG/2JdhwYbEKs5SHUVp9jPB+3FXrMn41uRF/wQqKMfVsP3xN9Qp9+yiEuXtrwSwGz1T9
KK2tH1SrYRhKCz1U0igvdRufk4I2WDV+HHbLokJ2C7mbfAHlSlMQP9wTLeNLIUxfEwjP6ly5jLxS
yW+U7cwEBZJNwvACQKEdsSkOySiD16YKAXY3zzWn5ZN8+e/mRK0qZSQHtYgZFFyRtuC4IRD4ypYw
2x8NWREXPJs4Iso6WdYuWhjVYpDBZ8nSv4Ej6eymckZ9fsgQrQPTRPUhl+Wd02jbq4rtfvAN40lr
DG7G8so2lgmm9TFTp72FV2T50jB1hA+1vkGGjKFyfzobF3MpuON9tQNsvDrmjisiBWwjWlIO1IML
cCaJZd8CfHMgLZuXT65lV5G4Z5XcYc6oX01HI2e3Q3O8jW0aD9iLJoYUmGfvieoAyRvg1iEUEBgz
7fjmSnhPr46XyLpb0h25+V2RkEpikRZC6uwHdmXr9Q4hJGdCQ4i+u/BJrFV6fDwwT2a4i5JW1GE5
ywH48dPqNnBd4TlkDl3Ec5kPj/Hcj65MkIveHMD517mTWa21hTqGrZSbtM1IYPyy1IyuZlSU/BTm
aQgzChwLjXWCcifj3+mjlIIpFbZlgCoN8UM8h5jfd1ff3yZT6YtlXQYV2G3k344uRGxC9Ime3F0a
yS6Al92PFH6/CPQsm3CVVvIHcEPaH3raRhcR6t5QcU6CMkRKrQBKYUuARAZwGX+k51sUgDGtjeTu
WRuhcfYE2pHOyS93Gr2AaUigUz6MOcOB3tJaL/7nzWd2KSBrSrIVfxdTeS4SiLuZLj+rx2IMKsJR
qGq82ysVZqG6w40mKLoMSoa1G8CdMDl8iZvRQGmMJjun4DRukHPdJdrBvNwkBLjmimtRJG7j9Klr
XcKzcXmtn7Jjh/XsZjADhZ/5FAAaMiifuGT1bl+jCwfkGPLhzj9fF7kD8VYWvM1zD9VRvIhJaYdl
Botkfx69xoJYRxkgBNtoZcOEUgeHJxfcibM4PtteybKHalm9ADBBYPuF80PswwXw68IiYXr1IkoO
VIkjv49d9DmYjlqyhzkqEt/tGgCGr/sYP82x1ehCK1wAj7poCf9OcuZcFyb8NcuIS3wwaP7gMD4U
3YNYsENy7Yd4vTzcDLTJNBT7YAbgTr+WnmGTMF/mH46KT+yoB8jDeppjr76k+hiih3xBK2VLPnHI
HKnJJ4biIzopSHt19axULnDePo12wa5q6vNcNW1WchFdJAGUz2R9Z+IOqYUh3jDEybio/Jcf7Ib6
FNkklChX4zf+1NiDQb1zrbGXZuwQ+hHw/XE1EU5e9BEzINr/f+d1GZhJptEgeeU4qPLN8Z8PJ0kE
p64A30XFHji4pTwNUvh/10HgWtvPKxNWJTrJ+iZsv0+5WUJGDOGiCnr2vJ7j1E3viX5LlKjigIMw
Vgz9CpskpdkrdExAKiLqS8uO0SXW8LTKP3iOgTWWNhlio6Eumnxdr5JJizthAvpu+Obp7wJHsoGw
Z1i2ecB5EIxVoPMH2CXvpHQvKrOXzQsWmtdI9ACZXvllAPqPB9VSmbV2c3MkUKKVs6HrwOs+6QJd
ng3565K0VTCbghnvHEnqzw9bruNW/lyrtrieyfPSK3TofP/F75HQ6WTFlzSt7/W/KVTibIChqTes
mGE95BEowZR2rxEFuLPzO9MviWlsNdCFqGgNfO4uKnjvpbL31fUL9cyC6Eh0gGMav9KDS+aRE/3o
uQJUXK7TzCqCKFfRDq5SvA1+/cakjO6c/FrbmwyKNqZdGaxyFDm2TAHPD9ZTi9cq2RT29r5Yh5Jf
O2OmqTL3NBoqxxKPiQEv4+YZRTDROLUGf5ZBpBLf7oU53djOfLgJa6U1+zLSzfYkxFeK++rxdvCN
m67CSd3qWfoHUzvbDNoFhqGkdeVWrY9KcB8ID1YbnLaE+Q7Fhw09Pmbn1pV5Y6RhuWM1jz+jNIky
vpWkGEPE9H/b7ymnrWHkuycYjybfae76ezc97gOk6ZEaAImzosQFzNUAFS2ja8B1lfcAcjvOLJip
quQLaHJ59dCB7Mgb4KCXGU8RIEcXtjJ0dR8b4M+LJq2otQSvBevem7vIDTlWsDBZnCX4zUXeK8zo
ki/vXfliX/r4YIl4Aro9ox1hvAqL7G6noUjXYcT8mhjd+cxbTL6bMTPiTU1ON9X3nAmIJDVLsW2m
RwlzNNrj6MMoJKM7EJmN79iQC+57ae9uuQGyuN4+k+x4pXrnfSn8L847B87axxVsRHWp3tmVZJ1c
YSAp9uGmOvYKphWwjkkCySJO2pEMyumwk1GuSs09J8wr2qU2Oz9V/ys51UNbh9Bt6XyLECcdSoiL
Bi0O8sQiY4jK1AYAoq8j4rDsDHt02lb0McNIDLaq/YN30Xb2VHljJMfd315dSzemMqGbM/EHHIQX
gDYmaVTP4r+z09cSBT45TGS4S8nJVKWnT0NNZhc7BLDMUfd4KozvwncAIOYjK7dSFkq9y4K0H3KY
bWsJLigaYPb/Fh9bkNFihVojf1KN5XwIejGpTQJoU8tsSLlAC49Th2T1hEoBCT7mE8xmpYqumhTP
Rgy3XStacg9K2DNAZfFfZ+QppyhQDI6Cj8ogxH8gHQrRAZe03PzedKHZO6C06aOZBoAiLkNKhApS
z8PccueNwtmSeP6c20NqzUN3dTqSVq7887GIqjDcMd+Magsmb6SqlaiR9B0TzQVYdAr7w/8GMyI+
Vi/Pf5Ss+o8dpBIibO5G5yYRF1LCZ07pzQx/TxmQHNSHMlTPtX7GDnAqnMMnmuS8+pehrO7S+5qW
m67neoD+r0Tzgz7Ap7TvNtK1HhOWnFOBXGdm7VrfSm7p2v1njd+bzXX/68R2q4pIkBdRFdBclzL2
MFQgfs3XMd3lxXgyYfGaIklz1IPLehJ3KZJKlCzheKZD7H6V1wBfwXZykH4xshfrTFuT03gQ2uLP
0xfEVLzku1TAA1fLOLHuBGdsTrzmeghoZfKLL2hhxZjY9AzhP9hX4MiIR5R349oHR6L+j6iGPFuH
iJ/i+oHaRIz2fBSWoq0H47mj6lzDFPS0NTjrReo0TiNnPODUv+vJLR3JL8wCF6Op/vMF7dTiUBly
AC5yfosX0WYKR2wOXGpn8MmlwHWG1TsDNEQu5ZaG6WuDnJB22RZf+8/3UGrnTCUeMreitm5YFhJY
ceqtTC4mfAI57WcYAkZoQfxC21ukyYVUEKr6ivCtWIv679boUojeOmKYXLAWO/44fuvN4TYM+1Ej
K6UxZF3Gz5OCPd28NnmbNP3pn77mzoNiMN/4YOVERqbd8NJYTGUSzQplNhtk40paNsTp+JRLhC9Z
PWQgqMByoZy7My0RPos29CU31DU5Km/Y51BFSXggJ17ji54VQy5One2aXUxQToDkfvEtRKkYGYma
s7uueHh9ykweeP6ZhRQ8g65S+h6S6IcJOxgtHKovRfpJSXSV8qRnjHlf6W/i9LtbtAF5Yo2Z/1S7
v5T2yDzIPrEIYGF54r0l5TLYvNmAclx+tgMuSB1Zv6DbRzRGOBOMhddUEKmEb1xc7L0FZDThJk84
/+ZXiZ48mewiarQmKIUPsQTAnWnlva3oIyPkjlrrlbjKq21Bn+D73yn+vGA1vMSbZ/LvRrgxyjKj
Z6jO0Y1KH5LkLCoqJJly6f9MJ1fqn4JX6xG2OTvN5D2Eajp+pCE9zl+8SuvKHXuLMNzve2DWvORd
gkZO5asR+omX2hWoiTuYTzuSLOsRSlKCyWkyg8z1b2FQ6VzsUhOpw/VhuCPBBGy9ULWkkPSdAO8M
a7KaEvAVldfqH/SHEqlwp8LrZSEJ8if24fUDLi/Z7YAjq7CsSzo7FxIFaWhQdtfXcAIDicjCr61m
UaZhgW9NBX9RJAeWVHNL3x6ejE1BE5oT5vB/Ac8mEcQv82jBOmvEuBBfUEnvm3K+6uD7Xbbvr6iv
sjJfYduWvhbHBpY17UrH+5l+e8NB14X7QxJ++9YozGnQin43r9rrtxcA54FT88qs4fLTwWYyD0Df
ih+jP97YdhdgoAIsVKw4/0tpkU1gwUV5hOOGSWCzaynFkRvsZz6bHypbn148ryElUQn0KKH0a5pm
MaozKjPlqWlR+x7ieRbRteMpP0Zrqbp/sxdwvyv0l5bEBwjnG4C6MaiMBTyxmTsm7b0jbtIP8mR1
gAdBsWvFL5j/lWa7Snm3IO3BSHgpXXzMpjGH5mQKzmwfgNGf+DFWdR/9/GQ2KYRmTL35zovajKHC
IIaxoNQG4+E5UXSugxLnXJ2cfj9wNboIoCQDb7shuSZAjTomUIm2N8avifU74f+o9QJUdY53JXal
AzzrKiLo+6AoizGIDE4+hd76hjTbcsYuD8yzprNnZ+5qlnLDL6h2Cz882sx3eZu2vKAsfh4rEy2v
DX4CZJ+UgK1vdj3Mn3RKNbKFpjxft44gqKVcUtmEGHy4qgfu/eJ4BHxFWAyJcMklfuIZw3FfyAEe
t13iZdwtiLbdl98N5yaQ1Eln15Uu8yYRmZd4cVXxhrzYrWov9EJP8PW0cFqiEYzpnNLatKymUroi
WYGSquxFoxiRXsOj9lznjhsR+kk5AR8Ga3qu8rAb3JEEAeRx0+B6kufPiA2FHomN6qVlFLc1BjeI
RKDTPaOoywsfi6GOWRPjwsHR8IBYFlzLIuPlwyj4QEyxc+CeouLAtq5wFAXXaKiu+E7clDTbbtp/
R3Ptrtg3en7g2oQzx1PeCP/+rZe5CZ03dfmN/D4Lv5s+nm+McJkrZW0BUoJvYBXoNSj6eseSQ9Bn
lNas00/MSShMYU/uQlhcjou+ceq7lP6H+CPPqygd2VeNajEOB9dsfDmCzf4IHtKqUjbWLUouSvyI
HZrlsR42YwaGoVeDK+W3mtbS7vOd3QvvwtI+5uC+iSM+DXLLd4qmQkoGEUblRy2MwF0khYwpEyuW
8F1iZJMg9WRyT8eRr1szdcFeHE9R+syBjts3yGDyq4vTxFQUwfKGjcNf1Kfnppaguq3BmMOlXPf9
3XgRTi5kyr75BL/2CwVbmLheuX38Z2enNT7tDx1zYcg0gIuKkQOamQng0R+OK8mHiaLTKqWhFnrk
xKZEoT7iB01HJpXX6NUM+rIt176rWyI1NSxOY+4VdgYTsVIPyADaPUdKr/RDVtoIAEsbHYRB6Eo5
kxvB+S8lEl4FYpCTpby45ap0HvZhD182O1tZiI198VOYysviAkl3g87fFFBz4X9czAWslsJr0ZJU
hJxS3EhI+9y6b2F/uXHGJuVE+J9NuRJmZg6naHTcjPxOh1yDR/lwfK+bE/ySRnG/IkSG362VSFoB
xWoQ6UHjI9SaAuX5Ei34KaFDOaMT6JY3phEPyTHcg4wOY0fTJyQZ+8ojsY3WQbD+B9ZObPjyK/og
zUP9jKM+UhmLosiFc3R7qS/F1zIq5bEwseuWfmq5bt6MOanAehSgHu9tUT/NJVg3jsRZnhES2AJ6
g5W/h/Tvbft5r2XFIFU6SXLs6QvJQEj4i6MOX+8FG3bDval63f02QfRnEJ24o1LhLLkRaBxuAPkG
jqJIeWygG+OmPod7jZvT8KMcyxYudApPfFo2GKbv3Ja9i6AmrDI+ncZn9SlkJ72VLa27zizg7e8F
x7uC9meL0mpcmHF4sQmBprh7EQUNB8Koor3ys1gM4ameHjcmOV6jzCKoUVkT9fxX7RDliQOYLL/X
+pJbrZYACKEdbHoHJOU9OgVqsHv1EIOUv7hIo5BsaNGQSyjy/umTLJOzGdyQ0YKVJJIXJqlaHcA9
woydydAOVv2Jlclf77BBObcozy44yuFaORUjs8I6hMqCmV4HEzY7S+dDnJ6oe6LNkdecEkOY52Fu
NyHmvlRSJkl+39Xn1Ih5sdfveygUQVlyS4T9+Q61uv2DMP4qcyrNUKtS8RM1VE7BM4cZdgr7Sooy
m+3TBu28nQKs9AMFrrQW0CcglamrjFD84tPcrPOxyPBjDVFGxcs47UxVYzvuB+y9t4tqbd5QtbNH
oP18b01sp65vJMRW96B/7eQaHah0EaaFhXuLWpFjYYCNlnPISltiamIR/o6ZT73mzzN0Q0ekIQNj
TdM27zfAasGinX/0hBVnlJ95Z4WQQcBL7z1w8FyFwGenDEfIaSv3xtpSdSHucSWXjawcM6HoJ7Xs
V8450Z/x6qtO+GEn3zySA875FMhOvoB19Tf4llltR6OTl3XNvUeMJkIbHj4GA0ER9vlwWL+P5+UY
XVjpy0Y8EuvmfY8GMrRKiFidJpDWgBUXbyCWGlMxa2tzjnzNgMrhfNJTKEAfPt+IeA2AfhQRw3W3
Mcc2pd8nC6h6/M9zdNbXFOe8QbbptMTLa5JVmFZdY4m0kJRyJA94G5d8HM7udBy0mSrdWXGDV2tp
kEd0YESh1czJ4ecxP98ibCTL95kOwFGHiR0rU0NP12f+/6ftSEz0j4dXt5PWolRKaBL0l9MyqJXA
lfrPfBAciNvKEns++7AFyN2uNKlREsGalSaZa6B38eINBu9oIzvu/wSQ5eM5ZLaVRX8y1DG4dix3
zpl15EWvwBACJFfw/9kgXpnWTN+8z8+DHakGQ/6nPsWe36qttna4YzNbjmge2CpzRsBzq/Yr1vwY
mbWMR26nmiVAYbn5zE8fBq+QbGXEBr5LecvqOTdjKNu6cIvf+eUhj2EbgLVg7bChP+wuKv83yfd7
178TGqw+fcQ6E0YJDEKvgsD/FJ9oFHKNkpWdD6JamaNt+2m/lM06WSu5jyIRRZJmG6pp7GDkrAQl
aYKez6hw3i5Qf6gLr3YDYEqyhzYcZgZBtl0v2FVRVpd5CizJnVqrNfLkvQJRbJU3SNGbgFqrOSTN
ma7zsKH27nX3P8U4I9Km1E7YFK871KHXkh4mLgwLkeoCwZGnHiqs0jsDVTcWty6GH41LwUVoho25
s2Csz/RRHzgK+vYHzrGQiW/FxufXXEMYKvapKX2SlhOr4fgbVqce/zVeZEIstSsPzvvAhJnIzHzS
Yndw4HDDwxOErRM6om0v+tjdCppZ3DIz0wCHw+1m3dnzxOja5DA1r+brS9p7F3GTGU8sZY9AGnwp
PQ3ua79AUObhYv7+szc2VZo0QXwfTlXgFuyjBy0EjedFpvyLSziOu9K6Z5seIiXVqOptoiWpdtXL
wDKnggzUa1yn9O5LkjxvdSVHBDx1et/3js7TTP4FxhbX712UoDCQI4TZluy5aO2bGo408Q9V+ymh
p8hzHZnqvqytI13g+y0gMyy2kpDHU+yGAqXkzn1iLS76pa+JoeIuCILB8ptABsHk5DSSZhvQqt6A
7aVzLmEBWm1IRvmJwaBwtPffr0tmD2ozoZ4nunOKGPiW2JxEEtrVQiVhsR50xaRBBWrJ1Z+RZqZZ
K3K9h1uBXdK4oOlW7nQ+6NzR98e2nwne43VCWJquL2nNXurehRFy6Hs/jGiNZtoOj9z6+ay4d78/
Okv5VWWFpBI8t7NllElh1uqSbmRh31Nx4wjFHBS3PYy8pkv4bxGGtl7+PYNPwhFetT+7odIEYmdc
k5TGRYnLqzC7fPi2j8RuImKIcxtdyvFkLhWyPE9pfEpqRkLirnhX2IexSHVYfN9Cqi7M96Euxsk7
lO9ScHZ5ywOXoVPhE+9wPCe9ZfYVLOYOd6uTEJXdtQsRgfIcvv9QhOgpK/TzQoi5DmecunvmlAEq
4LKo2JwMmGfO/PPYtTeefHT6qCgt3GgC8k1PH5TSyVKYPdNHTIT1UyUMnam2udLRjTDRRHRWgbzF
4xGXYXXmzfUnWvDqNkiQJfQMvt/hDgDvyzkxSl0tbaJi0RfMGO8iX0i4RraFHUrW5hs2HVEoZfs3
9obmU5cdodSc0X3v+ndWCuYFeJt8MQWWacirqdI40eQF8/YfcWIBZl2yjloGHaZ6CKDVyiWNDmSk
x4MsBIb7bTZuMxI/hCz/AeYC43GrbEwlNTMQ9ba3zFnrPLUUJWJnuHA+hoNkOdGl4rIwY8qmYdaq
+C39/Rs8Csk10J2htGJlGCyoEqrzsR3sBuArWR5TdK+KKhcspA0heVY+nMTf1E1bsZi3ySdqqyC7
MiZGPAAJuOP2td1fcNpq09HCqGTUHkgm1J7d2QAC2IX32gkZUqvpOjqwVmbil1JnkgtHU++QPRBd
MIZ4mw3Qb3Q7/goQcPYaIvA0yR8rURzf3zz7V1AiUVPGcgs+lCGNC2MjJ2jq7tRWoYZvD7k18EIC
ViB7v4bobd1mDpHJyq7L0lOXGQ9oPb4ttlVKo/FuCXcRmw2x1zCbR872rGN0Cxlw/5s40Eh3gdNm
ZyQ/Y6oXsQaMuHJ17tjitS8DVY196saVwjsacslZHn3iblaunR6hCsD2+nMZZv0YP5VOBk4ffPgh
tUsmiZdK58HowTQ9yEvxLzPutQ1DjPSMnv5+KwdPVgU+zxEb4ZXxW1/kqI1Di6XeweMUCK4zadFK
J7sJHQw+YMpIee6aNLIE9jIBahlmscXjGnkdGCzkPzd0rpciHM20wYHKrdwsMbuZKYso6I8k+z7O
fazI1RiktIzPogZWi0dI++cVCgWYSgpG2sOHA/oP7JU4nhPhFyXLXK2WmsLeOVaPWleaw7yRROUu
e506YhiJm6je/4xob+UIlh3Eb32EtZbOMODsxMlTJR9yjiHiWb/T3EGv0sG2YJ15mG7AHEyjKDoS
/Pt6P7q516fnxeStfRzRM0KYFua64qlVnMJo+BR/M5cvLaeZCB8oEL/Qt8N6AIZgRgU/C4FVid0/
aP0qf4EYlecTzLMS6pDXjuDd2qpBWx72jUvYGf95zSPNn2oL09hSruUQ0NfPfatgM5GgTTtcwkro
paeSwUqbxQRXqS7wo89aFi+BJnRLf5rO8Jr7zDpK8avalSATxIjCacHcEILneKd1pBGVlmOzfMLb
MCzgbppSrr04DruiufQU6kpQXK7eJtkdMqb5cYc5LN7kmnQqBIdzmTu8n8xlMHdc63mIeOQonC5h
Ro758dAYqv3UH6odz2m5v7mqOEoXKCgOX2RWvr4tyUQxNbFHzsBA+eOS/rJyh/v1O8fH/Iatub8/
+NYhCvOazBUvU+FUHa0Zuae/UbHikVbsJRVFYVS3Wd3xZcBZxQ9EF5yI+oCDsCIYtjDCNxHu3k9e
BlI5LXl/cPhfJJxBhR3wRkdUBab3vG5B5AhG4yhxMMhpTM0r6DlkvqMvWuweqz7acfZ8HXHvZ2yV
WQ9XJLFgdyyb41ryuGjxDtGqU8rDkT5AmsdR5zzX4JadfWutEN5EZCGaFiv5VguThCDOjfNm+nWA
9YnknPD1PCAE9U3EL/T5e/Yvz/BEP/mxnAhao6h+SKwfjVFL6lPIHmIBChPeLKuHVmjrwA+Dis2R
XXSpQxfyYCNiFvOuAzx29ER8owQru0TbRG7ay/2mwhhlJU2Ei2m6lf1noTTeScI7/BRzcAqbEbOU
/u+nUsXULZhsCAb5uD3DWG0fSPdspG+2DVK0q1/kcnNyVmSdKFgMUMQtM3rKIMDlyBDpAMypD6HY
YDnIMeajIfmP852Tb/6enzSxbs502JLkNDly1d95Ys0dUA+Xnr3Cfu9RzmtEB776x5w/ZhlVQQ/m
79R7uv1SoCVWvGX3Mpw2ApbBwKYVbTLZqgvLl4cFAzezgIn+Wns+Am5y3FMSV4L/cgDCJKYQX38p
Y17KnKzNQ8pK9j2zWUY4vlo7JTnT66+wnv7AwGOlAtn+5IVOJquPXJ8xbHCMaGPdnLOSVybZ7f8D
0LRmMPD43ZvEd4arhoPaMcx7LbxBhvsjKsHaABNkdYejDqPDwltqZJwMxDKdVrowdKWwLqZgGU+c
VcfrK8+MNXXAtNGsnWDZkl0rbOJdSO6yTK9ajRyLkcEeE42tdO+sD60Gx9lYbAFgbgewJgPvuNG9
Mkpav9aMmYUE4ZVz0HnVTeaV3YyNlJe9JDNRm6ZqnFhaXHErl5FLO7UYqrK90oXK3JiN/DeN+1fn
Q4qzgVjwQ3cEK1xeIy8NXGx6oZZsRwk/z9CS1hyg4pxWyxQn/zFgszOatZXbWdMrEBCeGsOedkwc
QsccAxHJNtPjsnsQ7SxoNTAyk8tGA956OclC2zC2I2A5UiSBFHCaGGDexAxu08rmOqnDa1vwFMLv
FxITPJzz2F6SIanaUx6v0DVtLdxvQbndKP7+FZnefdY3vgRmkhhEz4ExoeFodnrsAf23JaQ1cdXf
xFkyNjF01K3eeShY2Q03HrEASQJdRsKkrxgrt/MlxGlH7jfmKcLinGUtjHAOI++pviD7FIOdai5g
4dHGWJf+2p8Ylt3fd7fmsiH52JnMGj8WlnSYzMItCD4SlM6+Lf8ezx3MluR1sPzswm4McJWcMe0d
F7PqIwOBXqPtWgiFmhS/iB+5yil/c1DILX2iXtRD53MM40jSuKbLZggnFy3w9wgRMo6gfvLbMLrc
ppHnSamq480cAH8ua/PU3yLq3aKNfVkwA9FB+QklzzSq4ibZMQWRY6aUnHggbVISTAy5M3+9p8wM
trebvt5YLlHgKlU4Wa3qeY9sDnxr6sVwpX4eMyHaZRHfk6Rab4R76IsKM2Ce+LHHf9C0X9xvom5t
ZQ/gnu+K4ZH7jJKNyOj9KLKskQE7IZP13oQs2+0V5Bt8M68kKP86sWbWsexUJJbKSGgXtolm+/yR
eIHXQhUQ2d7zxNdvekp71JAtIACf6CAbQXVIzGIMPxW+tsFIas5Rl4qXbIyRyiAc5Magt3YuBqQA
HgjhgxlDJZzTRimPvvzgjd7acfpo638LYDF66nFpfZGADy1a5yXpb4/1aNImccyr/VaBOPKO6vup
w3RNHwLUwqKtNeVr295QxAGU2L/3n4Z1wiugTUxavA4R6YkOETLVwRqHFDRsJhTrAo5j/Nsmupfg
UkFJXImgd6k0udu0Mv3wIU52uP+4AOwO/fKRcL7FjMYnOVFnbu+RxYNTSjLNObaixREE51AQ7OJ+
trkv8DhECJLmkDLx8pA+W2ZJzidZfHiLl3SWCC0b/ATS6f9IqhpmfRkuAhBJMtN+QQZPiJTCq1IE
iArSHAsTyxXiYjJkVqxelXOOFCXr1p24BMc1whniTvlLQFkokgG1Z2Cd17LO67TNm/ufgVWL2L/w
KFOV4kU79Vfgp083R2ePLbb3wba0IvfTtKAvuGIJVRJ65fiinSdXmOekLvYrgGcUMNszIqYKtHeL
XxmWqcyOynt8viordRE705CuXxjOq8Mb4QL5ly0ircoRso1UvdQ9b3yhGOowPCZXSXFYSXfMCZxp
mnWhPSYLOxZnvC+Ylz4bhMxxAx5dM5UR0ptU/e9TGJAzpr7pyGMVsoQNeBLRWgSvCNIniJRtCMBc
M1Jr4zjlCsn18dfxaDO7K/TLY2tK/ncagdWtZ6w3yAAeAVN5GqULRu64vNIC/zuJM3PEs0KRUzu7
1Uv0t3F+YrLGHzyEw1muvgMCMg7aQqckZ8CRMv1djAHW2NZDP1ag8ajaSgc++cwC22tolkw8XjpH
EQzW9k58RuC4ZFNSB4dhA8XyEcuE5sPP7P5wjbFOh1cgH/AXgOFahs4pbb1yKFvu2Ij9EqcAYGSM
Vxv1q+tsBgzOPD3QBmvlQWCPBC1DL4rkV3Bfmum/khcvsG6vkzQr4zi6Xi+9WispAN6wh6gKZdgk
j8KbxoAfPzxQDnM3TH8m6iUFVhM5OpTFn4wj6jGFDi+qFa//jKMJuU9qeaoBetL9QEAgsdAlPLNA
3M19xIN5kdPH/S/tKvH+vsPWCqjqO50kSPqavc+r5azEzOFwvwua5ZjjdhcT54NdAPgB64TIROTo
kFGwk+h6T8gaxPaTO0ynGdPHqdlb86Eq48/LY622B/IMVgPubUdU0wlzi3N7PWGkGZ6pdFx+Vncb
Jo3RtKcmJrRcAQ5C9/fIOjv6JIZFiKksvYE+f242ROfG6a5TlG8CaW+5fyEfJXyzgJdr1zky2TYV
Sos/96XSMhgkol2MYtaq3ev/njdDgu0gTVnX3qY18Dgzw4kjjAYcUYH2lJWsZ32z5q1HDQpDuFdc
NTqH5jH/Vn287dj5s8RoiPejAqfQ0Fkas79D9ipkcp4O0MnMiAbaJeoIbbksGkahUQ8ghNKCw7ew
sSE2JfPHJXalt05Vv4TtFyYnpGrmdrDaPjeLu6lBRj4xuehLMKlmRWUcPgcMXmVNgRrvCASMonDC
6R2uQ+9xFXPA5B7bUjSBAwky/zkUw/Ze0oA9PuGI6Q8aRQtb+IMjLwZne4Ua6uLh6GhZ+4d/W6uS
vYt4GuV4sAgk8rhq2tjQ7fXT70PaB9DqWhAo0ZDvCXsXWRAiOSjRqMFQlkWr4MXso+MOIsJIbUoM
yzB7Kzm/H+zcwghuZc8XkyfGwvfQ889bFlrWyzkWUM6Acb0FPP2JwWOM+B9fZrzMk2vNoyr3nJ+O
eyUxQVtJJX12dnY5vzRVxD2h45z/WTGMtRp0gL3PShjFWFzsvsa7gA5WiYt4D4xyhoBVMrj3EMGH
ZcIEHRcKyqy6hirxcr2v6LoX0HMe4l40+AUEcJYvHTgdMFZmcGgx1DN2yQN3Hlrqp4yEiyNBFg5m
PI03nL8MV7T8rbmwaOI9OlTLm+H/IVRJbZBAadIRmG7UNadsUZes4bTpa/bTwYajtJaKms3c2bsH
YNpAQIOETh5Dc6Y7eIUrLa8Iw3l27jTY5c10Zoj8W63PhnncUL0wED3HTY0PAd90lLVXau028hmp
8TSx75uIWVRysmIR1s8GL6glcs3ik0PzDYld9vpn9uQnqi7A7FIwwl7B5Hq178HyO9c9iIv4RCRN
g3/3iBxrgYEr//z1kz936a6AVHN8h9wwiZM9iOCeV77/yN10FcO0kgelyo8xz9yDd+31U3lxG9RK
09fuoU4WJN/o13+6i6kAXuyF+4GuE9H4lMbnJ+nreKY8QF/AX8ykwOUF+sIZGMQxuZRipe2A4/V1
w+NRsngAhrtZo6U55YGDTT9LxYLfK2KHVCN0ZnhY2+rQFsmizzIb2zsAapQ=
`protect end_protected
