`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3664)
`protect data_block
xZ5RbF0ebqfYavDfLYiO7DJ2vJw2qR2HHEq73BGfsJPiAaVexgZhgtwwYkkNo+XAeV0kP2FN/WI4
G+xCnZWLnlmcPwq1Zsr0X5s+GT7jR+mp+CRvXhDfQV3snK6ENlFQKfwMSqKtFvl46+7yl10YGCx/
OME2qxcI4w4xrijnHt84EQEuLHq8u49yLgeHhjktf3FyicGCAmjt5B0wZ3NMCDC/AeFZDJZ4xWvO
R4DTxQEcqGYARRYzI0ZkMKjUveOlT1vvyEW96oWH/BUQaNpRzni2LEo3fDkbc4xLv/96pxTMrALq
fZYdQMmX9MgTmiaHsl/GihW2ncH6tmlXibqpIvkkrIYL6lN36JDgZ6BEc4jvWPm77mDxRQhLs7I5
L153j0n8dXwzRG9AwMu80A+FIZYsLSmJ7P0jPyASjuUVRmj96H74B8qBk6K+HL/nAEjPThx5KOWE
ZrsP1SsMLsiGJJFG2nNyk3dbf6GB7toi5eR/6DQpFRUUAX2maLCX4je4PdrTLJlEkhoxzQ4aJaRo
NEu6HKasWQHXTzdUz6lgOQkpayxA64FblEOKMcSsxbFL/6MSgeuwrhui7ridZECdiMbIAF/pS5Aw
39Duou5erbryB/hD64FZlJe/nApKdEnS+vGm1tkCo7fuNOmENEvw+B4dq2MS8nPvGGV3fECKTHgz
82PNAEMEv/xcq/h4lcfFxjNupHD6koC1uNJ6RtOPXk4Rk8GoskEteumAa6jQf46plPX3BvGcqvLW
SMcb/eoATrdDZKHrGGU29iYOLprXca3DcKMisFbOztqUHKYnzX3h75nsnPwlPj/rs+DZdeiScKWa
0euFk1CanN9/fHefuc18f2kyzZqRDVrcMobVwo5Tun75Z23HboT4j2jr3aKDOVtSX+c0CzYuX1Jz
H0ptfPnYUavq30MKnDxQgLFIR8zNXaBQA1UH+B0hZVsEn1vU3bdmbMqL3xxSv52UR6A0zzPBkNBg
YBnmIXtkj2C3dr9aMrOBou/2MPQ+qzC91Z8quNG9yVQsH08vFo7Zi4/tUZLm9MT3JvbqIVOdgsAE
vJ19Ed7bG7WoLzLxAqAEnfFweaYM0Yrkp7/wZWHJD1TP/FW7vWNWN7lFnVo6Pjh5QoJIKN/FAhQd
ysVK8nA9sLDs7WmteWHNnKrOuBoWSUOvS3Q5G3Ap4LAR1RBSKO6W4bSOcnd2KsS0q1arMkKRwhqw
RTD7kPf3BfIRRp3Qd5/OyOQSOf6ehabxWGReBWCNRFdJveS4k2T7A1rFGJ8IgfrwGf5i1qQ5kvQK
qycT4OcH1LaH8tsbh/VFfY7b9rQdXMEFQtKYMZbMwpW+cDdMaHBImTMvtKlkdQQR9f9GojByQDth
/gutM634oGdmDERYG8MRhmyE2RgzMJd4PqdRSygx6EhADg0I9pRqNy/FbNnVZJm5awccbux4qGV0
IAo4aWhAkJTjIYPXjiSykWxb47N+3vCmA26nxIsfTux284Nitge6KCHrUhvn5PG3kls85HVsO2A6
W1BBWNvG6DlOg6UzmvWYFeSd4EIRl6RdXS7CNZCKXbNSeZUt8c2i+Rqf5Cy2mS5yuvN4QZxCajLC
MndQLBSOgc97yY9gTSvFeLq8XHMfRiBevDqeUZRIj+bt3UlHyl5Ivpx6Lx8sI+RkBoQ+hy8VTYLW
rHmzpeQK91xW9aBXddYfH3/48MS+2+Xju9wehRDdI4nSKs6oI+sVtmwUeTz+khrxFjqlfgk1bW2U
2aSTqs78qjFklnk7Q0ZEGRbffg7JPwO+TpzgvhWTe6t8svMi6ymYJqZUVuC9LsPKZfo9hByBBn11
JzS3L87UYPb7BBmRQbPQU3pa388UUmlcshFKIlZIQ+s0pL7Zn2I2V51C4QHIpt4zgHMRxBkTwIiU
bE2j541Dlm9iM1jZJbGlo5btiNk5Y5flaHSby5jtQwnVqhWOzZmQF1VQVsrmVjxmYv2e3Tt0t/tK
eedCw3qQIjH405jY8RIA6Hl3UpTeGxX2n57IfRl1aulKGwAVY2Vqd3C/K4MuN4O1sp5VxrWh7qjm
5ZOjZto2oWBuebsN17x8cu1ARo9FFG111cfhKM/RVvdJ83+wDdZ2bSLYERRBWG2pJi1YdhKRCZkV
bZePvW2vJGrxJsjjLHKUP9oxgDTVQEU1GxQwJYCZe6Op6xB+JUpKlZJ8eLJCJ4X5LdtlVz+BAufz
l4v9eEIl68f9wYsULg/8nd61Ywsuhw39bX2AHLIcTZWiomTwbA9xHcAgPlizo4XWat9Thnjtpjsj
MM5HMbAAYt0oByuJITYyqCHTI81tGCUogNE3NStdLkw+9cUE8FPrM/oGNMuuIrLu0Qh6U+iTVkef
z5546vvMZRMg9FSVpQE6gWwOHG6ElTLDgDJLEbz64WHe37dCFdOo8gGVLgJzxCdmETW4rk/DudpZ
IXYlpdqbWd2wquMrkVgpeAo6BKrVRJes75PXLHTqByLhl6WfZ8ZARZloB21z79IJUJhK4YSAnvif
ZrPDrK4/wTJ0dvjcY0U4dnsRxD9v/fuMOTtU9TK+qhZmIEerIbnhmzIEcPN/XG1LeRLaMHXLBDrO
4FdW4mUDldUzIcIMswguo8VMYFCBiRe7fDfd2px+VQYRpEY85KnQYCBbzD+IjG8JRrzFCkYlZI1O
+tgTzBrp25b6foxAXn6Vu6dxCUTqgzsJN8RAWKNDWW7t0sAlm/ZYg0wjykKOBaV2mxijt3PkwxMI
hasLIJorBjonrM7i1oe5t2M/Rj3Dlpr6SIt0s65JHmSMwyS7yDKuu8f3bfyeY9uONYneYsVTIg5t
iCR3vhxxqCRz/jRIsWVcOzQVZMUn5Jm6S0Yvfm/pj3zcEThUX/4W3WgzAz/lsz/3E9Jf7HGgn8+6
SUXN27GjnT6BO53vpfeq325gAMDQC7eF3nEX2DyilfkD8faBDieMyFKqH7Ulj2MeK4RrAOFWGRoc
1jJZn0fyVYLMOJt9uWKqIg/c9JgT8n5EdVqYt30hrcaH+6qSN2lYduovgACiNGETZKl5wP6Hl524
yEQiDlP9qhsI54cKp2YfpaK8VjJSvh+KfsCDHSMhq74FjylBavRJp9wAUbE1CNI14VW72gkCFhCg
U71YoIuEdKi/j1Ipb6Z1ZxO4gaIwdzHIBjITpScKNi1ciTrFVaxCvsNBzMnUgSTN15knXKHSpWKU
pF5+Sdde8rarw5zpIe6rMPkXL0xuD+q+2N/CzfqMPW2PzAphwYlk3Z+4iS0w2udEvBPAmd73dVOC
H9XFXhoeIq0pHudXyFcpZnaO8Btl55ugERwVxMkktNLaJKd6WVqyL1ZJ4cE1NEiQLZpksAI19C7X
SIywwOLJboIfl1k2qh5XdYm1C+lqT8YAXOlSC6tfysQGUYx9QoIgLF780HMucoeRHxoEcNCMuvos
3nZXOwQFvz8IktW1dAdLzCa14NIZJT3ABsxFeRRbTlBxMYA5apnUuaKvzATthSHBaM7fK8KMRpl1
6l9Vl8cGr8rXAS5lujRv3p8IRBUKxeRjEudMWYsAPyZ6Q8aIk329+KEVJcdkgZhTW3tXRHJSDLLc
SMHCBTVp5vUz7HGmt6lCKGaL++GU4OTVB1NKmz3V86oHiUAdw8bbvuilQ1RKpn2LUshDOxNCazyJ
A0KwUwzQ47WOQmJG+zblmMYR+1qVl8P0A303mAcakvdTuOr82FqQX7GEpDFFHquUsRSdZNBUl5xr
mTmWSBNuSnUjKvndtuVMx2LsAP4ABo0kN7CpP1Dux7sjlLM7drWGkREbkCKm2yCdqp0gwO5J5URB
1c2XLq1ZC/lNZAdpDXILCXNz8QKIrqa7FRFH5XfDwN53TyhGMRdQvtkGpR4H01f1h1Cb4mKK3ryO
hXP2wdVEhjRpEgDNMT8WBoOxIybzp7ljyFxjegJ0sCFooi5dzaN0SkZrNLvYKRre73YONsi5mu3D
tiKRWeun2riHnFVeKlTKG09jpZodopiHem60+Jhcnb47KIBNbZA8kdRHrrf+sSbvuMJ4LqwhvFHE
oHJBeHqF0OK0K5VD7BL31wHrZczZh59P+GyvT/ODJ1zDMNYWZVOlQvz7lAs3e3WEyQVYWgNZfRgl
YKXIMI+xD/YsaAEmTJVODa3C/uFt4qx6rVKEDQX1Pi68jhbK6zNz1vRUQTiFwx4A1HwEo9vxQnD/
APAlV5owkwu9lFW1Cfst1gLDex+jOjFI07a0M3gHCjOOGQTAlz/+0oGzGkcxLPxWknsl9yT3/1S8
IoLMIpwcDRcQm//VtVgW6GnxS3UBJAnWdTENiduZbDGgs3nBcDDO0XS7++/UD8hCHoNX2RQ2ABxz
C1NoXZJXnCg7LTAUqrbZlRZvFT9W95CDcCALc7c4fchNIm6iZuEP/31IpYQQ188e4t8HEgQ0X4CC
0iTbT2PJ4uEEleJzl2kTV0kEo5oU/jikYNoY3WpoKH/MHPLsHakxRQ4Syl/cF0de5ImSsmfzZxGq
nMrBaBogCvWzu3Vk3qcAMZdGiUqfsNvYayMqhfLMaTwdjIBnddSPzLjlc7DVJtt/JeuTshOZIZy2
oIClzgEjooYfIDO5EWRmrXmEpYjDAwYwiku3npiGty3ArYdyjQCF+3YkYglmYlJrFpXEBMCzAkBV
649Sc/jIlypDdiUFXz47o6ZHtwg7C4DwRtwmcuIC56E/wqzvda1KKQDEJxa+HOLDKL1m5nirJA7C
gxWG7A6Hh9G2EekzD52Ls9UUbnmNdz9G5f0vkjHVHDN9va+raMfAtx+s5Kqp1qapiVsqpG305Scf
7R+OhYtF5IDUVfEcHr0hCqwRzOrnRw1b4RVuI5VE/sQGRZA01hfQgs9LmSvJSDVfXzcs9SJgb4+T
Uvjjzse9nTXg8bU5EQ3+kQ==
`protect end_protected
