��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l����Z@w?�=;���:D�~B�~[��X&hd!�͆���G�e����g����TMk�E�6P��!,N:�7g V��ڳ�ѐ(�g�7�)^*-n���8�>�re�Z-��aQ�l�	f�Ȏ3d�U����O���Y��Qj�2C?��J��A��n��p��� @��}��X�,&%�)��1�8��'d�����J��+�3T~;8�G�g�T�i���sB8�ƚ�5u�lW�C��G��e�
Ӻn�h<�85�>J3L�d�=���qc�s�:��UY*!�ZeF�N���7�GVerr�\�_��(V��F`���"�l�� �1�����&���xD���;�ADo���*���H>�<��� ʌ�X���4_fu��dz���˪�=(�MO��ɖa}拿�/Ye)��]�G+��VQƴ�+� �+��[` v�jvU���;a�t�c��s#%d	}���j٘Ly!l��e��Dcc�����������GG�p��iP�~ݝ����/���&�{�Χ���t?�:�YI����U�� @���Q�)-����OPb�)�5�'��$S��_c|�GT�\?�X�˖|6XK�m#�L�zz�c1t�|��F>(&����ߐ^阢B��`��m�BSEUWNt�d���p�%�e�4y�
2�/���������}~���Rq�A�`-�C��E�.�X����"�4��鷕j�R��/.[�R��I��� �x�Ȱ�h9�C]������2P�r�4*l+�N�S� �ȋ8�� 0 \�H�6�5�var���E"*�X\��*�a
�}�yH��]Y:�BH
0��vRG�i:!$el�;.�i�Up.>��C���qT�A�&ÿ|��qŦWisZ�`� �ڧ^�	q��#���H'D��5�,��vu�%��.8A�d��2���ͫ`8�Y^��p��U/�Q{;�m�\�"��8f<4��,��Aޣ���ĥ�eF/PG���.�B��6��b^ǜ��XWXb%��qT�>>��P�*$eŃ�e�э&
:|�=Hw�#��FG�M�h��1�8G�$D��FVy~U�
��0v��"�~ZC��w�Ղ`�5� j��UD�$Q��K%t�a{!���;��d��T�{�ө������V*y`,=�D�ȍ��0�1���ƿcD�,���y��τ��a<b��|�n7~�B�L�M`ñ��Tn�������9DwG��%����,���!V?�eS�@�g��r-����L�s��
8�~��3��~�e������"u�&1���b����8��da��~a��])�)w�5�Ц�Yx:w��$�+��)�`g�<���P���Q�]����%n��|�������Ԏ���d|5���2�E�ؚmO��4�1���N�B���U�~�nX}�v��<�C-�c�ͯ�s�3��y}F��8�'����u;�p��6p�$���g���� `71`V��޷����'^T*�%͗a�g�)�j���x^9%ٓ=ʠG�����Nk��v��iT���S9#H�t��59���7��)}�y�A	W�	��5��a{�r.��_����g��|1�Fۨn+����G
�|m2��Yqt��k �@{�GY��cE��9���ii��c;��n�~mFă���2��2���u��aL�l�����Ѩ�Mj�Ϫ�ǧ0+�?��RthҤ�76���	�y�e�4�+�����jJ��*�Ǌ&���6:�����~i�f�zs�2ƨ�r�2�ڋ�'�����aPK��������CV�U
Eϙ+р��{�0��ۧWь3�����a�el�A��d��В"�_�5e�NW%Y|^����y��}a�.����%�J#���3J#����B_`����s�GW3h�^������
,B�b(�n���mVe��@v�J�j���\艼�"+�U�<e_Y	UL��GFޏ�l�,�ϖZ�D��w����a�8�$��D#�����]��+n��e�Nܩ"E(ar���g�a��gz�~jU����t/Փ���l����L���Ա�������!W�fb_����HD�'��n/��\	�8���7�8��\�su[01�Ԉ��M�Ju����HX�%���LF�{��'&�Sɝs�EQ�a��!#[R5�PZ���,n�C��@oΧI����C��:�h���
��v|yД��g�\��\�^a����d��'��e1�EE��\f��MqE��#�mɀ>-�Ǭ�������I��E�S��ѲlY��h���¶��Ɖ�e�����H,����E!]�J�ƋS8���8a�� ��͆Q�(���J I��W(�*��3�2W�x�58N�*�=�Jb���^����OxJ6,���Ev~h'�#�d`��?����G����9����l6������6�l/G�����ix�cL���'"l�ua��k�T��֊ׯ�$:�Ba����-��ǺX���eN[P׮_S��XZ�~��xu�{Wh~�s�����ݺ�t�/����ki��hrM^������/Ф��\��&PbZSp%�*'��5�\_I�Jz�A�3HҵP� �]�o�x��%��(��E΂�L ���2���X�Jl�����0��co�����e��.�
ԗVS�]������k�8+x^wM�����
��?^����`������G:i�  ���r.6�3�3�`w�J����}ht��bX�0,d�>7Q�����`\��!���0�Wpv���M5�ToQ�a+��7��WxPQzy=� �� ��-𾡪+���\g�[l�=ճ�㮐�v$ׂ��w�5�LѠ����2�Y��~��C��_�_q'L���e�sw�I	����R�|(��A�a���mͰŷ�it3dl���8�w��텵���C�-�!����'�x�����j�
�����,�[�D	�+I5x@p��Ed_rE$}�S|o��zHV����
�r�@��9=C"<[�=�A/X<N��N��`�-���	<V��=i�0T�Dg���m��G�-M��i�8��'|��sv��^!w�>=$��A4�Ӻ$�Ac2��4���nCﲞ���]j��u��T��G�������On�Q3�y�:*�q�Tln���##h{�������F�E5ɢ�6����`�j�� uK	�8L�؎k�aܜoh��ʃX�������нr}5�Uz�s��R�M���EO?��s69�h�Z��}��=���?�'+��-18m�����o��M>���w��^�B��ޅ��
$u�����]\6[�[��Q��H���/���\]�7���M��߹�
w3�mx��;���V�f��@�F��9��{i��3
6��Y_{���x�h{����\L�����+���Ij{u+��p@bM��p��-��ftA�7�!"F̷��^j�	�?��D��$9>QC�[���1�Go3�k?a$A���I�y��l���m/%H0a9���ҝS���dQ��+:r#:�!NK%*��4t�a�,�*:��j��Թ�tj��B�� ��"�� ���Ѹ��ި�8K��e�l��p V����n� i�{�+�(i�����������m�oF˄�@a���74��2xH_���RZ� ��AA����l�����.|3r߷v���F�ʜbP&�̖�y^�R]XѸ'�=�TIT�Bo�nT��\ʲ���p9O����r^��	V슦��!�JN��)q�~p#�3�F�֕�U⋺9C�/�I�X9��ش���QY �b��v�H�^|���n5�&�3�Ǔ���~��������/��$���n^ u�ڽw��ޠ/�&�V�Ȳ���~`1QF�P�:u�É�-�KXM�e��@z/N �=�pXH�b��_dB���|�;��8��x#��8� w�5��ŹcR)�0��?�.�(�t��z���qF�l]^�br�O�G~�x�@r'a�]���ڡl7��>��00�Z�Tj{H�*E��'=��k��W���&:� ���iޣL3�O��b��V�C7{���� 9!�	���T9P�u]!��u
�'��������
�V�0W���@��ď3��>lVM1�}�2�R-���x�(~�S3��f�C
�Q>�%r��H ��Q!|ă��fS>͔�	uV@a�ܔi���(F�)��,��	9y�	A|��2y���%���+F�	�W'��1\�,�w�*Eƥ�ȕS퐦�n�Z�Ԉ��; �O�z�&�Uc�R�_��
B�n/,�|O��#�
Q�ix��2�����);��4�^+]矕2� ��LG��/Y���=�ʪ�M���ɒ[�+�n���A��J����ſ՚JS�b��6��-��0�o�S��v�}���r��Ÿj�r��T��
ԔQ��m/���,�|�·���u���Q�c��_�@��5P:1�=�qL�E���ι�Gcvu�e@F?h�}�">|j�2tr/���[m��?�]���ܤ8�݃�s���~��TP�Qk�䚋�9�e�^y-���" ���'B2"��x�@Te��s)��p������΢��f�����0&��f�^B�As��7E���u���q��ԃ ���hJF�H:GYQ(&?E#v��
�6�i|RRI�����=�9NH;�9!��\u��l?M�J�<Tp���9;���Lcq-��In�)M�� Ut�����t�,�;>���w8.���}�����q�j;G�RY`y���u�=5梈l��~w�5�H��%�e�i��"�1�%���*6��@46j9���c�3���꽕4��z���+HdǨ�w�MN��u�mv�A�O�(J�AS�tQ	%o�O�
Ȋ�+,Se���	��)~Z¢�{|�?�oj��#S�"� Bx8z���7� �{� sG�	��ԨC*ÏJ�

�h��M��b�A�Uow��pӆ���1SW�	�-,�����g���B��ݒ^:�59+.�z�4�ʗޅ��j:�_��~zp<�0��P.��	�hR��2$d��S��YӃ70vo����&-p�����ە�`�Շ�x$+�-mW��(���g�t�t��O���c@�ʪ���s
!H�({�;�����v/��'�{�`�wK���h��� 6�q�ўT���věZ���ym�����4h�����!i�1���o`O��Io"�� ��_�Q3`��J"�p>��~e�pK"���3b(�$3�S9����M|=��*�����3��py�(�������P(	5��1x[�%�����_rx��;�������h������t�/J���A�6�<"�ֻ�,>�YQT��Ȟ�{�����R�q�?b3��k��Ǘ�ส��-��nT�T	��u`˼���<�ƥtc}؈k�y�T�*��#P����ݞ�p� �P,Hw�T ,ߊ�2}O���U�P)��ݫ:���I^�Ju�Q�Ea'���Y�"���܉�TU��;T;��B��)C:���Z$J�w��A�p	/��s�"�ܞ�%@/12oF.cm�/wn)_(��4�;W��\�4f4�GxcX�)������LX�SWLj�Y�D�xˆ��/�Ő
���}&e�7h�r�z��gΡH#�Q	�����.:�4�˥��f�n�B������{l'I���V�q�5�?�<47f�b
K�[,>BҾ ^Q�%s�-w��k��Y��ٗ��ߍE�f��x Wt�oɃ���ڮ7f�V�b��Z���zB��F�%�Q&�҂�W]���5Q��y�wvP<�Sb�~<DJ��1�d�_��������y+ �'���*6+�B&�x,<��d��O��G�H��㝳�4������o45�������Ϙ���R&¯�vL�a����k��g��%�u�}V��%��,aS��j�>t�g;6<k$������.R�5 ˟�1������:�@Ga�؎�K�ڙrb{p��CF͘x�ք7>-e�њ�Ψ��"$�,��4�����<IG k2=U��6 ��G�(�h�����B�;��"�ΆȐ���:%��Ѥ���tPip#jn[ָ�\r�d�)��-�쇈����$���ٰrUR ���>N�IKd�JIO�R���M#�jџE�V�����1ʞהRv�¦ ��#(�m��Æ�>k��Z����|�.�\�hW�7'ܸ���񨉚�&bGpMvC,����I��2�$�W��!JB5���� c+�q+������	?���o�k�D�-�Ĺ5ʂ|\����P�����&���[���R��2T$úS0z�C��R�����@M���.\�(��d	5xhc�e'�׽����K4����P,$.��|�ޯ.�4�����yTq�߭O�
�.�:�}/���B�+��&���������w��8�W*'2ᑴ�4E������"�Guo�ѕ��a���Ubvo�C$���珤�2qU��YΑ�2�?/'b��f_�t|�x��~��xoܴ`�&��@D�׼�=�s�������1,��&���.bVz����/����'0I�Hん�L��W\���
�&f'���ۭU���?T�6܃�����JsrY;�vAH
I�F��V�(���w��A��m�`/iv�;��g�x��?���xP�)	�	fۚ5�Ή�{Pґ�u�	�Mt�޾�"��I0�{|#�XRNN�s��3��fNWS�ץ��\��| �e���]rn�h�8w�q�j�3�#Z����席�#�T�B㒖0�A���E��5��r|�+��r�����-�TC��q�ߕ
�'S��'��c����@��h>�"����y�;�S�V�)aJ���rk}��x
L\GK�>��� ���.���������@j��J��!��B,�mJ'f�Y?ƕ�2	A+������.DO�
e+��x.9p��Ύ��6�g����Cd�TfWE(#d�ǜ����m�<A�3�u?v�9����(<���Ju�\S���Xց{����s=l>X7X .êM�>��"`�.O���~��g{�G��Rޯ�l���_Ubx�rqx�JҠWs���p��L�p���>��ei���"�;����u}N7��o9b�x�m��y�Ե�]�M�e�>:�E�e�9o��򂑪ܪW	�5U������h�#_VK��oJAdҔD�G�'L&��w��ԫ��_��1}i�	���������Iw�9��5&��A<r )l�q{�a���6!�WML�Ns�ɐ QB�'Z��k����mk%���N�-f