`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
sl4jcNVqRWNkOWybbtGTS0ybVRmAQ3bbQnCTLFF/qcfAloTKWUKyHKJDWfxWpHYUuN17pQLM61Vk
qxHV6Jk73k7nZSraAYzvw+rBNHdy2GhnfbYOD7hYSuvHE+h+bxBgoIdmQZq+yOR0ats02eTCZB1Z
xhw45Grk5luIDm0GnuJFDyNBvgioqZdaYfWxUnsytIVCyv+VdLMK5HhkutQmT7yB4L79e1Afhr4D
2XQNUjZqntZCppRGnwyCdQ+6lDBsPKFJ2aLvvguWNylNcDeS/bG87i3LyzRHfO0IgDzI4VzYDsEr
AzlEz7BA/HOvWN04BXDQbU5yOX36XN//S/jBZA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="px4SVAHRJGzAWyb7RnSNcT6tkIG1deoH8uqRj9O6VjY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5488)
`protect data_block
bEnU9WMj1t5GG55AI8rSpE2oVXWg5wRthss0AzOCgN4wFU2BqQmkzxD54NfVog4x0Zp5wtDXgY51
wJrslrbK4UK8k+T+ATW6hvckeZ2YUXO0ok48BOOgW7HHd+ERhnVg1C5ETpdBVugybi2nOPwqGJVP
+JprJtDtIUY+x/b1S3JcKMyHWBsUh0zH49CL7vFUi3pXzqny7O6ecFfVvlkpPl96Wm6AIngMhGDB
wGiABUaERsAuoK2fzwTit9eH1xScFFgYZ79PFRtomDDiuls42xUFHBlNEd+M9apNR6gJnuJMK2xo
pvtObiiNz2VV52QNppUVjaRkkr3HpX/l/415nn9+AQMOAwrn0XIhBfAEsBQnAX66OjJ6xgy3FaAg
1bDOYiMF2i214+8WFGaWQZdXgMlxIbjdZWqWBjvIJORNNfvA67wzC/Jhf2zo3tm8zSScfpzSmGpP
rMz6K1ne2UiKgC0mhPl0cE6ZqhNiCbHKnnYoQimFZPQtO4db2gj147fvrtnsqZEXWdboMUDmMqBH
AeToSWNGd3sxLGYCXmP2s9ByF+6eRs9cwpwFtaHK8HlWdiNvmxCBM1Y/2rnYFpEwEv1trUxfAoTY
ZXzXRlhKObgnnBueUZiuSPX2eBG6jQMAthUpi2dcHKKbzkF9GGvqpYnU+SIfAa7pFheYvThGEs/Q
/pVPjlSzfHCrsme9GomwQVsk0Var256+XyWoKiF0l7/3SfkZGaBucEVYTzXmyyxzbRrmoYL5M6VE
RxksfKusaOlqborgSUStV9fa2rraOkze0Ky1nTMof/Ju+nm+/vuUlM4WlJJ61+cDnUzxmoQT7wRB
Sxl28G0aAs+yCd+bERvlkcd72ghmYsVcOE5AsLik+eunRnTpFNm7x4VRgs+BYQ57PP1n3hGWs9ng
tqI3/T+Z4pG4wrdb+dQipM4GggVmwvugdGfG7rfX4oLPoHvUi279ACkYH8hbxJC76iBDkPj/OhIN
veoMU/Ik4oKfW/Flu+wS64n1loasNEuxAUayyZWonvbfTFu4bHCqRsVUflfL3s7tpxGadmH/39tl
fiPxZLWcvlMSwbSJeA0CEOEwFuUNE3/EIc6c+jVX7UyJJdrRjzRCOx6SaLfIQHusXxohS9FKV0nJ
bVrM31HmrTsnw0PEIxaRM6oJEXHLkUdtlbjIKoyZ13dZZi2c9DIpZ6gIQLNd4RouuiKuBBgRc13o
Wl9WKWtbW7VOJTG6nviwetJusKt1aL3VK4bH515xEIlixeAZ2qUXBXGGng+hcOWrftd2AI654erN
f6iniWkYKvoPJIA0/GtTVAR9xaw+uwSVT4baIkSZPaSUHrkWehfmohsNzHvBXiWXcI4SE7XYC3gh
3Mw18RVum2Y7teQCmMAGlguijkYm08YPSM1uI9vQuivF1tkGB5eHo31JpJ+vAfMgLC+g4MU/z9SH
4ayq3bMQadg/R+/cd8awyMuU41Z2e/CSYybII6R1lVMBJoET6zOrO8QVyMzhmZ/3FTxkd2enxo/c
SkTso8zOhT1fuwlLbiE54rb06Q0AgkTyX4UfI2+9U8kQE8urJnkFByDAkVRUv9Teuv9Fki06za4T
YwM9ivVC8omc3syQn50DrVPfeSV+wKdHYTGyGUYTnGoHznDUWEWuhCH7Kg7H6r3Kwrnmg6sSVi1l
Vz+i5xvvPezUit7AphC1u9lsDoyWwZ3IhG9nttGL6QM/OZSSMjAYHudoPa5WohEsYyZAMoyNl/Z5
FGxDjF3IvVBrgWHSXGPQD593UlUK0mxtkyc0BfMhlg/xl8QVyw4qF73KN8giF66hwE37F/W56dZw
8Bn+M4YGrq3cupGygV6xdO6HkGOYtlioXyKE01J3Qh2x2fsKEwxTdZBt3FNDgWa2429b+0c1q78j
VLgY/8Sf/2fJPz9AgHS32jH8CdxiMYwwpaCzTkhZPiXZP3k4n00vHJPyz/G2lGEUkiEw3dbV7qaZ
xyqsDmiqGPmbYfWBqbQ5HkUqL5uPsc5Gkaff3gkfCHUKpNPiICm0rHOC6Q0jSIt/8Yx5cp//nxUX
/n/8xr44OhXpiNVa5FqXT/PTNNMbXJq5IRrET0p7PzqMuI13IB4zIzzV2HVbvamFB7P3+YlNxDdl
FTpiHbPFNgas/ub9yb44mmKfJfv83XoD79qRnw/kWgAo8ihpnEY7J8ONbiiXYIzqVoZSGoG1SvG+
SW6ZSQdZFVsQAhHIorLc+eayweqUVJYewod4skspygS198wZZQlD8H/1pyV9BpNjjnlr+rAFeiA1
3UVU1m/fLfidEyfGGc6f9kqE97LUfoM75gAECRXnU/O7orBY8GI2CdaKhXUti0uQhJLlQcx56j9s
4te+FpKYao2CJHQlGL4pzhEkhZ9WW2/733p4mZKuRlXSGq2CAsXpsbLRTob6EsdYsJ+Eps7vOV4a
N4KIPWS1uAZ+DFhIi0/AurWxrDDNr1wnKOOQV+oP99E+OTeYjB513aFsNjkmXNvTpE1VJS6Jl/NQ
me8GdAsKLntzMeXC7GBIEONmGfrRJfNsmnrjyZGwaT+Rf9FaKjkHe/XiPDCEexOEVIK4fiqEya48
oQsEPofar0vnuLIm8WLDRXzILjPCnmWNfDUta5lp+obYXlaELNzelgfZ3vonCJaQNVsjDVMaxMCN
be/YpYQ4jPVc9GrA0aIOr3N9KhDmrxFEcJ7bi/5oRJiegpjLyqoXsyF67qBdT7ZRF+u5fQJbo3wT
GFft2NXuqARGp4vUytFMgRIk5sGxhKZNEx3s+mag9BXy/vGqH8/PyIXbKM6L7JJyh1ntPrcBlVtm
LYu8LjPQ4STKnyi5o0w/OIm3+5ckVe1WGsG54h53ANJlu/nzkSQ0KsLy4q9Yzx9OoO2ctMxP1tiX
rQeg0U9IJBKNvfmBvDnrDdM8o3pyyFaZTl1siT0RrW/q6mZ3ia8v3jcH7T9ju+oXEMi/6vvDQsH5
X0a1yP9lmQQPBQbo9AaR5UATcQh0q6yUCTR/HHwkBvC/nrJDZ55vzKr+7QdmqnXUfKu9YDufB/SQ
5GwQSFniHrxXyrWpuPwX7cOWBbILpTbR5aJnUSYxhdw6MluDYqbwE3bUla/DTB5ywWyz7DFa4tRR
FfrncAbszrSqJL940f7nnfHlBgYs4PrHIJkM3TaTwPWyGiEdlxlRBvkv7eC28hYIEKn0YpWWodn9
h4tOHII/ldcISnHezRH+fhsUJ6DeGDl0tmMsvvUAR/bDukceqoMii9mjHAuu/X3/fzVgxkbQNXMi
fBMgUv9pc6EfoRl+PuLlKfqHTea2bUx7+i7pApVO/29MXCOELwD+fqYaNuNKqUUs8EeHOlhD49/R
46+bXMkLB/QvoD0abSRcJT84e+5OFAC6D4t3NVIjaniRhYHW/nmMglNDDpT9nXSmndmg2hkctgGw
IsHmE3RmJKh/owvZRoGkmOSd0hd4B4D+YY2/NI6MRSvOfRfIMLE3MoxwiQ8V/9wvvnYwLGrFm0mD
bGGVyc9+ZEI1zh+Zgy/Pyf+Rn9NIo6VndnMUjqgAY8YibltBEl3ol5wWovYkwcys2jIj0JD4rpgc
1qzUClF6Jjg1Wa5/J2ALjczXWvN+EfnOA5p1OTcq+b1OYl8RcgG+CgPOhzDI9qMvI86mnG5TGyKk
Evvewsii/oMysOoumT+wlOPWa/3D58T4z0S/WZfpJddZA62ukU80yOcXuhKhMNf8Z6/St1qFTJrR
vDszzK2iAvcaMOaWlV1n4F7MKZ5fx1a2mMGdOx95iktW8wRnHUKCkVDTJ0pdwH7G+qFv6LFOSGtR
H2YccsIFv75PFt/wta9qn4c0ixXbzMZ8Puz9pfHal+tuazimbniEZACAkIbGk0y4tIdVwlcCmVTg
upLQ4XSD7KlvOtnjFwP0I8IJ1YsuQf661wXo5fTyuRSXlBKw351IHpaYMrRKqnobZmJO2xtuV5NJ
YF3rkwAZy923LkZpm2TRPBlJ6OoWt8CMLJZQvxpFUIcBvnDjLmCzxYCTeTO5QX1G1YOE8QeDhG5R
YB4pW2outyRY3skMP9kUUbk5ucvFWS/u+yERByzzadl/6mP4osWXfueuh7kfZCdtq8SKSVltRgsP
ifyn73FrK9BeP5DStC5E7pCEmSHlmVPiDon9ZHWQ+XX0gMb4mNZDki9CCMn530O9B0im4NNzA9PQ
BXWfiBGsXiQwkKwbkeT0rccJwjdl2cLQQxTRFPqrsR+kheVvFArG0gATYMU5pQQgvL6UAUMpuG/E
WOZrS2k/6uUEANJmXseOEnJxNm7Msj9tF8FsQDnp4jl06A6Z4fnsBX2OOCDkkcHKey4ty3G14wZM
mNSbhEOTFkD9A+usPjAWxRp9GV0tA4/PG4ge7KMP0IsbFIrv4zMMtCNmhnv6OgOsKVWdEQlEgipJ
Rpm158rC3aC0oO6rt7oBsb5Qye8qM9HvaWXd8H1SyD50Kwbp6NzPGJA/GWRLOLMXOLQO8sZEY3MY
6DKj0+2M8yp08nrrTT49259d1syDldNa6aJvO+xJieSRkjWUN+w3YP7oa/lwpalTQV0gjtlQDtTv
vwLhnXbrLquhA8sc2Dsu4ZqannG5gBxRMXkCxrkvkGhA1vZPHlp5VzMUImU6wxtCDN+B5NDbVJrq
xyWILEXuS0bYBw6lBo3q27zwvOySay5HhUb+WLZLlWoWhiem+KhAyux+CQbgvR9vJsYUc+zcxJET
d9NmJ2MK2KK0gxtXqSncLLh4Y9QL/RFuiMzBjQkZyM0Mxa841MAJrE+zPKCayyXHSN6dOcDMLEDx
MVRqFEv69EURtMqYlvg5HjmDTTt9qZX4O3+WQ2Kq+SrolHE78NFtieW76Ux7c5AB3xv+QXTLMTYb
UegdbkFmnuVVW1k98r8T4RHZCcVW/KYDq1buLh3HcBoxXP84MH/dFz72f175ViFx5LWRqDUUF9FK
fv553H3OhXiIUos6exDapWE+BWCPfSWZu45XQR4SmdxKNYFqNW48kdaCOnLBU2QbPFd6v9wIpEvq
TXNs9JIdSYNsrgU9hRC6Ja9tojoVXCQ4u7GlqWq4HsufB06V7yK/sofs9bxuDBXOcmzwVAFtoE7I
E0eDj84ttdDTGT9xzxpcBWg/Ixkvc776rqD0GlwNInb+maRWQ7VJUhlGZzH5Hum0iyeTtyLjFtXK
m/RD1HdpBON0ytJECroFrcQCyUbv/tTSn93EEd+Eh4NFdlKP+lmGI62cidEU9dcMDFX3a972tjC7
yvK8IHd5B96Bpspk5K8z7EmDUif15FaBSCqdvA0layMk9J01YI90nPVOZjiznygSiZ1lN0Z3t8cn
T5ACD8t0NdycQiqvbdv+yex5qqr/Q7o9ZzTnQ+D1QpAWw9rfgHHd5B75jiyMSQy3lAu1wPwA099W
UmbsPf5+bi2ybPYN/hFYcsX5MvVtkjK6Y9HPLeqSKin55rAh3bF/9o49tk7SBZ4d60PpYNkSxnFP
jDnlh9PE1ZnS4oH8Q2iBCxDq8GxX9WY4yux0/u/9vioaOoYvHy+29ln44K9+9fF8zvMR5+m7TQ6t
Qi/WYI5l6KUfT3ucYAGfxNAtr0sERmH5GV+afuhrS/qXhuBicraVhzEq2RswgQwA4tf9ievLaYv/
Dlmfj53VXEUIHIuRc1LG5qdQdgih7xAVyQmB9FrDaKPhwWAKvbvz++DBefyX9t4TLvReY4Ac7Q9Y
yXykBXKNiewYsb9pnyRPLpj2X/nKXA/58E72RAaq1Omawr+1LB8SVnshPbgiZb/kmA2r5hrYLvgy
3ECR5ZoySBK1yAIi8HiMN9+sfL3CurayxWaXip4yue6P3p2/beWAG8FBN+HVa0+9V8/4EOmzK1Eb
Tj9Khtv+NU4ao2ENsFVufgkfEtMfCxVIAKimVbDGd/Em0uuXfORrigJ7kjKxMQ4+w+Gbv/2Zsz9w
Ul5dFwwKqAi5UPWb8H5sWodxCFJiuOFI5HLnSvJVXWRMoM5859xAhvDiigvHBufMWrl4LGQO1TSt
Y8MQVJLabYuw/OeA3WFG6rmVGvViDz7EFigkICECvZOEajl/uo3gfC+p4jEPh9iOYDv4/O/5MGwT
47rVSJ/3pm1W/qQlKFC5yIDXIRb/BBeSIfCESlvKPtlJIas0OKinlkAYnkAR7cOMrofVMZBCTidx
KQGiTgdKFKHS9wpitSnVnQpZJ+r4nYqzHZ0BaIiF6Hs7pFf8cCu7R33EW3ivFv+Buc2FP2kCX8BJ
soOnwV5S9Av8CTo1eANozldzXx5vBuU+5TEtR1Zecs0Ziz8dekL3DcRIy60u9SVXSu01PiTheS3O
FTf7YomPRJwo1x2J7YuYyRij5nOWg2AymaYkYU6kyc9kvDm7B5q4n8F/xyIpNiDnCPjadofI0fQ8
iyq0CtYztvSzwMODiVKQE+pJJ05snZ7+fU9AqrgfngbxX+yJni5bxLLQVvctfOVTse59QnpzEj64
FA+PXIg8TLPymFDCfSHqdeRzNMUXNxb/dR0/dhwi0fSITSkNt7rawmrkp5T3LuOFAJOYQJlCptb8
sRUBoD1oPStt5cHUcLlZpLiHt1ZnO97dUVNwcGeOH3dBpORpA+XHcY2oXId4KewVdfrFdals84NQ
ppRtOEQ9OWVqGhG8UyXxjGaf0wv54luILuqgrVEQrav3dIBBhqczcnmN4Etpkqe2zHkjyUTCf5xx
UtYZsOySSWkdA9fN8HBrmjLYgVz+pfrJrsAj873jVeTCKJgtS3gImyVYt/OCq/HeH2nbK7teichX
TNCYlQSVo+qM1YuRdIw7VsYr+O0jqVa1+vhadObrAQqgzWT43J8CxKGGn56Bf0ubuZ8+/Lp4WgXc
StnIdBBytO/T2YX+hfzetj2dTuAEQn1bbqqqr/3Ai+wW+HYisQ0/oeeq4rm2KxZUARy9fEtflC/o
kVfOHy323Nv7t12lZWGNNq+8mfAWF2eq13WyjYoa7BAfrDF8JWUKc+OpGm9hOfcmSZDonI3SGKDD
TD6229Cp+QZXeY7qFX/nFhK+brHwl8dXVjlhbm6Z6lFY7Ppq/Vsvn5LHjvqGPhx4Yiy1/vzFZCAU
8zEwhiR2yUJT9dg3rT2EWgryhu+mLPc/Q8jQPWRIBlFEVa2Z5qle9uUkpPemb7KANRjhzKdRJLVi
9QePe0Y+pLY1d8qXFoDugUFoKs7galulwxuHmLmHAMEkfQW4quSIC5Jkdua8N/5naCkH/K37FamP
8sIxgt+4Zvdx4QysbNFSvI1nTSD/KF0hpgiBsGqRrecKI9U5kG1Ik+GFOK58NlNhhi5GqF+PdJMP
GU/kKdMK7/WzieswTECoXA==
`protect end_protected
