��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���C�F�.���GI�����U�YZ�|��G�j�d).�_V!ZEe|�;�ػ�&I���O^��9я;����	S��뗌�C?eQ�(�&{��_�7*���A
*����pRE��r��v��_ ��1���eW�e�痷�PY<n�r�-�6\��9F%�������v����q�`6¨�В���dϤ�����frw���`�SB5*�̄�`:�\]���,A0֭R�L��uK�^	A�o���3i�>��Yn��6&���L����jX����]���7sa���Fo3�y8��(p*ψ�1tP�[؏�֤��nW�[���9I?hY������j�`O/�?ç�$�x�5=l<���[.�y��V��W��9<���(`ߧ���u��Mo���pM~��a���l^"��	ֵ��NȤ6¼dZ,>�N�����ۑ����3������1#ˠ�@�F�}��.�o5�'�>����@�
�c�K�r��/��yw����iZ���>G�`,��dK�U���6oN:�֡�E����8��X��؋����b+jn`=~iy���p��^����z�
Z�Ӑ3Q�9��4'a�=p��mT`͕�5����F^9�<�&W��G���cp�������f�8�9N��"����I��ҁ�3bR�½d�ܝVیl>� v��� �	�lh��H��2Eyzx���A�B2W,AF��O��xp%;̞�Ԥ��$B��7��N4�]l��V"�쫸��L";J'�S G
�F�9���d�]M��{�iH���q��j�j� �,��]�r�!72�Iت�jg.ons�ė�F	��_�C8[���j-���A
����,r�G9�࿗J@s;Q#�I�$*��?E�at�A���.��rns����}w*rV�<�6L��e�AS���c�5Q�����X5Z��{�t�*w��j��{�%m�*�<P�.��u�>]8�J@E]�4W�s��a�v�f_�<)���T���$�n���ҬnCS=f0��jnN_ߨ�^ }Q��8N@\$X�f�U�3D��\R$�fFV���ڎtP_��Owݣށ�a�A�����g�`}��$�X�p��k���-���K�ӱ�%G3���p���zASiz0�	���[��S�<��Ù'�3������k��Z��%J5mn_U #��:3�
x�'Ko�<��ݲ�Z�V�Ѡ�Ǔs
'1��|�.�s�q��Ir�Ҋb�-os��_6��-3�l�ݮbg�},��m�h��&�N�]�7�˖��5R��!���4C:6|�7�^�\4_ЩoY�Cca�NU�j4�[�HB/*�b#����ð���k&-MA�ݣcE�|�ĩ�l��|��3#�d�o����+Ŀ$ΎȭL�̐�I2����wi���Bo�=*.8M����W�Q���)�����d6���|zj ǳX���#��pH����ܪ�q�rl'�q�(儙Ȱ�	-�r��105ī���.��E��]t�)X���vI�\'�Ǡ
���c�Va���u{
��N�?����%_���[��r��S���P
%�C4���#�Fʁ�w��L:�� ���!��~�I��@��w��<�MK�t�j�a(eV>���',�%��;��������9'�����t�Ʒ�.�A�_�Ύ[�1��NZI���@�YL���O� Y�l��3�!��m_9mn�����THBh3{+��?jHƥ<0��c>��G೮�>v!�Nu���D(~��E�k"���0`�`����}ؓr���xB�H"��Ҹ��~Gx���'�wD�~�ly�a(�<��TȘ#�)��3P�6Z�,�����
�;+��sj�֕�J^sG�����C�s8B�m�®y�<�e9�hP'2tt���kS��[��;�Ȑ�h���r)��x�؅Y����`����GYލx9����ښ�C)�-�?�����Ows
}�Sw�N���6�ӵؒ����Y�4$�fE��[4�.�L�����E)�QRB�~��Lb�qU�p��k40F[��5!���l�A�_%����мޥ�Fdss�.�G�R%˕�4X
י��bߤ^���<����+څͥ�Rm7j��J�u>��HLf)w�w��8��.�(��ȤK'�������7_LץY����A��NLk ��kM.��Jw���W9�5�U��*t�iH�_R��CT��"Q���^��4P��R]oi�tV�"Z��h6�b�>HXK��4P� 0��>�VYd�;9�u��j��ܺK���x)�9���H	��xr��*� ��n�0��RJ�s`ܗ��'��;`��n?��f����}�#�C��2��	���g���ƛ^KvLLm!�6�mS�1J�t���gq���ͅ�L�Mژ�eI!&��3K���R�H�0��:����U��C�"�;��T.���qg,�8q��K˿"`�0�!�A�Ki���[�*^5�茖ͪ@�&Q������I�3�@�;PI�f�DB�a��Y�L �h��2>��,Jp]�0������'u�8���+�o���F�F�����k�j>tν�d1�t�B~�'=��
�G�0�K�Erj��٭��X4��b����3W��*.�("a�a:g�%Ȋ�
}|7��Z'Uy�L�I V'5HԴK�o�.K8Q~< ��m噾������G���r��t�؉��ܦ���tG�������'>�C7�Au����A����"�߄}q�i	!�fKWEI�^���������%��e�h�������q��.�O8|������	\��п!���3��Uɑz��\ �鏜F6�x(�nx2)I����3oW��������NS{e�pF�C}"XA� �'^M�'�c1���� ����t�G<f�^r������Z��I��[��m���~�I�����߳{܉�H���$�k�l���~�Hf�w��8�"ęI�k+���%�G���A��hu/�&A~Lbd*q3��;5c�Er��K��c�VP���WF��@){��u�PW�e�����q)gG�Sn�!&���5(|�ѿ�?����^~��V�
��ϛv" > ,)3�����n�>w����y��^b��Y��܌���&���w��xǦk�
k��M�H��*��0�6Mo�:V���W�N��Ŷ��Ӹ"���E�=�C��� d@B���ܼ���2�F�8��P��d}İ�b/_�C���u�ǹ0:���P�u=N�ug��3ǳ��L��#qʵ[s�.�@%����5d�R~	�Rٓ5����K�<}����HDK$�cUL���%�nO�>Ь�@�'�B�b�$��vB9"D���,f89��N�d"�N��賧�#�f�Z]lO��bJ'9������1j-K�Nܹ�ܻ�� ������=��w�&t�I�������D�^��7�J.�1ԃ��o#
�h]������S��	~�V�G��n?����/EN�����2��!K���6o+]JY;�yA�-Pа�(U��)����8/·�mU<����ⲑk2�����햼�H6]Rpے� ��N����2�o����N�+���k����gc�x����/k��>��/���y����=��)	K�:��y��@ˇ�I��=��l��M���Ը~��#sɲ86
�%M��|+j9-����T��p�؏T�>��������-~��U.hOo3�QN�s8V��u�$�Xw����c-&44�0�����W�cF?���rY�D����k��j�`�ܜ>�01�J|�C1��FY��7R&k/=�)��S�w������u{uff���oճ�3�-�����d~�>��<��R��N?f's��xn��I��rf8�!�}V1��V��li��Y�I|�@��/�O�]@Z����ЦPJ>'�9#���]���CR��G)����d��e����_ ��̭N�+�lRr�Pڂ�ZJ�SRl w�"E/�`������\2+#ܓ��(��ĩu�>�y6�fmH�٘��J
���ο��w�0�.1D?L��[G��	�yH��.ME
x�A�*y�'��/����4����$q���u�iva�����]�h��LXe���F�R��&����N��c�/e��a����	ん0&#�����ʻ0��@^߁|�,�7][}��4�*}ϑ��sz���q��^w,���	9���#�x4��".2����|W7�g���h�H��gкԻA�����sN����3dx�˳_��ZT?��3\O�F��t���7��zօ��LÞ�|�/�*�B��Y�Ԫ���̷��-v�nF�1t�������qJ����NK��}�ρ�Oޞq�ld�Y*�^`e�/|畈$��	ɒW�3���;�\S�ȧ2�gB�n\�4�بn�D���.�a~��$�*��7��21���$-���A��wÜ���Y�o��u{����
�w/5���~V3��#���̬B��.�ᄭn0GC��0�kz���ʷ7��Ѩg�:�A����2h�Ŀs@A�Id���
�����l�>�ˊfPa�@ZU�g(~�Du+f]xӬ�s�iY��H���uU��.uJ��زLZR@7@C\����2�0�MK4"t�"b�{gwՍ�^�Jp`"6Y��jv5��{�ͩ��E��E��@k�����m��N
5��:3����O��)���3���E��j�6A���aæu
g�$٨�֨���B��~�>����i�CX1�Me�n�c��,���,�ʕ�nF<�t굲㸃?R���m�>vn$v9����и���l�A��ؓ��A��E���B�"q�����p��c��)��ƙ�4$�[r��*�6���&��m��9@������� 3gȟ03�9�D�D����x����� kĬ�?������B*Oj��Q�Bڎg�F��Њ�`�H�M�2a��5��p�+QS H+��/3^c95Sd�)PvB�D89�Zv{/4p�w��pǶ+᤹G��;�M5vta=0������f��(�aQ=�a�犪ť����+��[�+3_�
F��&��,Hze����l� ���_���kR��Z���d�v����hڂɎ���H��Y4�})�-����fvһ� ���x����w��<Ō��Y�H4�L�\�2S�����0
�!��m�,0ܱ��ٳ�ǝ�ƛ�NL����?�;��4��\��_P�=��dٸ�FY�qd@������3�T1\�ēݽ�7z[Z3�5'�Pa��7N�J��-\*�Z� v�D���k&��H��S=P��������Xm��#�k�����=2��u{���o��_�c�g�D�[����Ezg(�

l�kc�Dt���?���A4��(�}��e�4�Ȥ���0�Fb�;����6���2��V��'�-BP�UԤ�`�2�+��a�|�ƾ�&�w��B�\8�FGC�*�`@�l�M,Vv^�Ɋ�q��qk�_lsՕ"���=o�r!�� �����Pe�Lq?�Fg:�jd�g��i�����R���k���T$"T57�C�Tj�|�*�_7U��	`3߄�e�QǗS��:��o�`��>�O\�����2�T��T-�(7 N�r��j<;���!zT݋4�~�	����<��~�ӳ�ݞ�a��f��[�4��Z&��7ڰ��3��b�?s�����Pv�Dɭ>@>h��F�j�`�.��vg�y�t�b1���Y �L7���9tn����|>�A�а�u$
;h
�\����ke VJ\ O*Š�9"nr��
���8�o���gi�jpo�����3���	�;�}C�5��5hw>*�B!6�N],w�9O����qu�_�����D��g%�.���C�)�~�^%h/���Z����N���9/"�/�V5����G�5���j:>cd�`KO��\���!���j�����)�ZvQ� ��j�F,@�r�	)�:��-���Z�����Xm�TZ���1]�K�J�E��J�R[J����U-�';��@��� ��f��F-�ƨf�5<�kw"PEd�:�$�7}��+b9H�k���y�m��)U�/�~BD��γ�v-u�>":��\�#���2㨸��@%�Xő�jC��e\�|fQ(ᭇ�֮� �#j AG�8�a;�ZUL#!�M@�Ⱦд�ܳT���g콫V�p2��f�I��ߢ��c  ��\P�,��ɯJF>�EO-A�d551䁒v��7/�Gz��o�m?,�]�^�����
ko4������H"V�]+v��Vvy�I-i�|%�9U�f����N�+��3�Ӱ�)���d�%�[��������l�c�jk��8P��(y��F~�0��.'��YxIc�'������'WW���*pr�'4(P�Jv,a���L@<8����?���$#�H�o�}KP�$����>
�V�/Kv�:���*�[�&����y^��"D�/�YL�;�+@��Cj#%�-@щ�'�t��s����ε����2- ����qJr�fW��h
r�1�K� �Y� �(�4�����qh�KQ��*���="�8%O����h������xC&lG)�Gm
:k��Կ*�C f�_�a�6�tӱ�C��;q�@#�1�J���b/�zx���A�9�w����[pu����r�o_�����?���W��f��4Nub�{1*י���io�f���Ӯ�Z�!b�Iji��D}I�XCT1�
.:t>ڿ�09֮@�;���� �����`
� �,BDC�Nф�.]ҙSY�I�mf���QXo+�q&�TX��A|�Bv����>��"�.E�|*
}�7�,����E /�/�%�FXė����&��ql3��d��g�݌��݃gl*�R���|�G���]�$����m�}�����a�����@�m+t归�e��z��T���d�0tG�ŲH;�#^JI��/;�0�AjH�T�w�wJ�Al�)!5)�KCS�Favm�qo�c#8!�X�� ���vT��w������������饐�A_��*ld�8ԁ�!�7Kk��9����8��� =�}Ba-�_u2����1��o�R��ȕ�В>�����sЮ%��f7ʔu<^{�H��0`*�6��q�c��R�N%�������3���V���u�vH�K�swR��j  ��=�[ꂠ��P:�S����e�##.���3�r���e��.T`�*#E�$�\y��	�*��)����� �"��� �w�� d_�6<�Rs@�ghvǚ��}O���@�S�r�G��GxF*�|k��cp�ʃ|����w�K���MaR�;���M��>o�;N��9�m����͈�M�4�`(��;i�O���p�`�4��M������Q�����&'�,�s���N%*Ra$��^��e�m5��x?��(���v�R�Bh]�2�x��CO0si�'�u1����7��(��L1e���QL �_��sKOY)���� �o�A	P��x�%V	���h�k�HԎ-r�w��%�9�>T�?#��~uU1�?�RF]�����0���,:;�W�ó���:�������J�r�5�傔6���ƤO�צ;JM�C�n摣%��PC^�eZ|��ɯ釁�Jsхoj�����J�j����ᠨ�}���bf.n����J�����a�W&�7�7-*y-����,�x���̽ �"
�#A��CE��+.�K���KK�Uú��:�wm�yX4��r�;YI�·�R�$���p��[��8T�** ����b:%`�I���9anrӛ1�UC��(�aW�ɻ��R��ϑ�2b�9%��d�ӶG�
��2B`F�E�d�̵L��P�gGG�=[��Ӻ����LG�?�fTdJ{��75{����a>�y4O���(c8i�)�y��K1?.,�����FS\��G0띋�i���Zp��
�<k��h�L^�r�-�}v���o�ٚ�b�Y藇�]@̢�3�M�~TsU3nAF��\���2D��|���Z���_<��n�?ݢ�[y;��v�;dBy��~��Q�w��H�\���'��9N���HM4���f�2gt�K5��{��3`g�4pnW�k)�O���
�y�t���P��bI!ENlY	�ä:����܆C%�����3�=��{D=3�ڏKs� 2��i�����t>;x�1ޜXSx�P�X`�0�B؀+��m�Ͼ
)���v�؞�}���G}-D9]�ʡ6'������85h<@s/�qV�k�R$z@���҆�q�bq�"J�k.�����y���_����  ��_BBZmЇ\��
	p{����#���P0���$�+Gx�XGmQs�.�x	-�������jEc_��,a\�E���a�Td��aj�m��W��Ha�O��C�O9otNЛ(�-$��^�g��ά�:�a<��HN��Bs~�yBq� �XeFe�S�&�n#��e�R��HF�|Blr~Βy�����Qw���`A\��c�O� C��m��Ɗ ��c5���O}��|����մ��7�r�4���=F�<uA��u)�+T�ct@�,�+N�Yu֥�k< v��-[Z���jE�4�>/�N�4��$���� �)�����{~E��¹-�>u��߭7x�!�,��Ó��0�X�φs~�`����d�aD��Y��"k�@�\�7t"�>r�`1��^�߶�']R�䌝Q���N�q�"i�d�,�9�ֻ���O�b�X�tf�&��ꍋ3���g�N��*�V96K�
s��yv�5cѿ/�<�v����ȵ9`C���3Q$p�7���s�Faa9�� Z�m� ��(�g;�/ԝMּi�f�W�l�Р��+���:5sj�G�D[�!F����W#�� �' �s��W3�ņ�}�&� @Y���+.`�K���C���r螋���6YX^��_e]�GX���kW�Z���>�g��P����������>�$z��t�RM@��x��|�kaW�E���a��	=r�4�����6I*��:$QhE����EK�U%pk�3X�Ѣa���b7*.}�p����͛S����և��4�\��vzW��14�'��+JV�`�K��h��\����0���{ A>h�Ź���FՎ��Ic?�8��9��f��DS
�d�;�d$���a�O-��A���ˤY��a �����J}�G���בq]��V��7���j?Mi���_���)J���>B��j�M�st%u&�_y��+����t���p�)���>�
�a�0�F`vQ9'���>�٠���%*P��:	H�(������!(s�"��Q�H��⧢���n���L#�"�-4���\.����YDl���� =��$�J)&���όR�T���'|@ce�`2h�1{�� �4��
S�Ncپ�1Z���M�6K��Z����>g5�"彻r"JBՎ_�)�&ox�N�O�X� I�'6��c^րt����#��H��{ԕ�:�G]yP��Z`���%���H��RO�p.� �f��4�������JO�z�a:�~k����d�<�O"I��	��*����� �ޙON�c���s�u��{�Öi�%n=c�:dN�T6����U��ؖ� ��jP}���W��]��,:�Z2��R�������5�+�*����T6���6f
cm+4�\#s�p8�%h��}�����R�6ӵ�[EO���0��f�?2�)?�V(͝�v���Ⱥ�����(ΧAx@����cS<����oL՗0����:*�s�O^���U�TŦء��fG���O�`�Y�jzK�R5��WbF����H�6=�ѩ�]�.<�7/Iٹ����3���^�%�������Ia�M0Xr��w���rb�>�v���.����ޕ����=k>*z�'�����zNn��{�2Y;�>1�T�a*9�(����ȩ���ȗ=�b��LfTN~	�ą ��]�����{R�Hu�<n!|t�ⶳW�בb<h��Q�C@x.�%��1��#�Vmܦ����C��i�tqQ�I�NU��$S��)�C=��}��9��F�Q���K!�CR;��J	�Z\[9��'��E�r���ي�ȕ��C�7�H��NV���^mCa�S�	��J#����mzI�"K��Yc�O�?����O3�q��>Th�IuM�p7��JՏ(�R�hQiVS+�;�7�oLٟ��LQai��k���/�L-�t�ց�l����č��ɑ_�A��E�X��ÿIp�I��i�~�:���Eo+=�� ~]�"&۠l��`C��ոfV$����2e�C|���O�Y�U��@œDz�Mٗo�/s��p�⧶�>;X<�?��|ez���B�����8d��|K�2�%9�e��bfM8��y��,kr���K/�`nF"(!��V�[�c&�E��[��8�P��V�Z�62����Q�}��,��L緇IEv5����Moj�e�W��Cf�Y6���G���騉�jn-GX�{)Q����e�U=^��yN�v��L*Z���Q�A��z�����T�^�t�Z"��'�6Q��I£��=�k\���l�����:���봟�#ʯ��t����B��9ac��6��V�1�Pr���T�㤥u0žW���Uw�_\bJ�mL�2 ��t^y�g�l:��-"C��BE�g�R�ơ�w��'�Pb�}y��w&�UnN߿��&��mt�].8�'u��y�7��V�Zj�C�9�p*3�u���{Ys!���4^��ʼ����5��,)���i��X��Fϩ�p���c��ޙz!�e�;�8w���'��gW���l`x�����#a�W'c�%ET����tS���aFl�d(�A?f���N	�Cpc8���R9�@Q�L���8s��?���җ�>��K�'�7M��>��ѵ��Ƭy��7H!N�����<��X,�����_vn��T&犨R��K��# +�k �j���;�c��ަ��Mn|
c�.�1�Y�C����-M=�3jC 6Ƿ�V������Ļ����By@����!ԥ���u)�N��ޖWnK*���"��n�-HL����/�,�lF ��:�7��Q��'b@��S�k�V�)#z�q{�*J����~������ۃ<���]�]�<܄!3h� 5T�;l�J�|���$�u�/ɛ�c֌�a�v���ױ��Wk����6S(����牲�I�@T݀���^��F~u���z+q��7>ége4	�!��JxĈ<H
��ï3��i���žQ�!��p��f��+9�L�N�	��\T�+����2AG˹���%9�ɲӮ���%��'ZB+��G�Io�r��Ҧ	*��4db���@���.S�B��Z2~���pl3dn|i���(���ec�ќ�SZ4�n�8�y�C����Q �v$���d֡i�}��p{Z+cs�:�.�x�%K��߆��H�Qϕ����+��ɖ�K f��%��J��sK30��
��	ۇzy���9$�t���c�Yu���xa��n 3O} 8�e��	���q.܄��_�lzi��c�T������}�?R��˩������A���%��-�r�L��E5���HHu�甬�ޮ���|H Fh�l��1��z���m��X�/a&v��]���N�L�FOL���k8~4������\u;�/��[�BE`�gk��_�����;�R����� ����a�Q����t#��HϤ��A��7ս}ڐ��V.kG�
�ߨ��5����F�WW�L!0��{���O �Thaʹ�ZJk:;���IP�o��3;Q��6��L;�M��M�#S�,J]�M�8��K�_� �X��G����_;�m�k��<����������Ə:d��P���IX·�;7��I����̔���S����z1�����&L�������s�W�+̔�k��*a����ӑ�H�WeU���HV<�G"Eb�B��ÝD�7X�݄&���o����IZC�+XB��
ǜZ�:�u`�' =��O��OamMӐ*�j��`&0�Գ�+�9NيK%{K�.gO�s Cw��yf��`+d��^���=o]*����k&@�EQ��^ϳ�t���Q�|'<'�2��F�>X^_K�i���T�g@��T{J��i�s�H�����H��+h���o7JJ`nR�B�=@��X�����!M�T.��a�Ce\��pa�xuM9X����82�j�kb���3�mq+s�i����E�;��e�f��׈��ϋ]2��y~~�wK�M_"7)�Ɔ-d��Tg<��6��''C��7�JL�g�����uk��Ҹ��1���F�ճeM�螌6wf����$��+�%K��d\�����a��J!��WasLc�J��$�^1�֡1��F���쬿�����6_kd���{�'>$6O�^Fv�	�M��)���3���NG�8�?Q��[�A��t�(��=jԤhiz�h��Ə�������^�.[�)��@�.�]��7�����i�S�t<Y���$�?��%|��X�t�rxE�/�چ7�XoB�mG_mł�[Z��K�øj�Љ�`�Xi>�;Py-�)���ɐ=�;�'o�~��U��i�<��+�]"I�t��5O�9HރK��!��r������� ��d�6�A/*Ts�ѺF�v��l�#5��bE����#����88aI��0k�)�o��nQ��M?K$�i��L�ġ����m�_E#�P=L�-��?�fS��&�5}+N ���NT���(� �������{�Y��h�VQ��)E�fe{��wC�o�-�M.E�z�ʄ��V*x�_�>�O���(�C�@LRd� P@(�;Fs��E�pŠw��y����!�$������0�z�m������@�S�}�*I���6�o6��*���I0EZ�Y��3�PO
��4�;T3a�R�f��z�EIi{�:uq(��p�2�u�Ș�D	���)��b�`�>��/Yo��A�<r_�!�<p~���:n������94���s�%�*�TUn+�
ٶߔ�lu��+g�_�{��C�%�p���1|�{��S【/���K��U��[�|Ú�t������NЈyD����`d��G�V9����Ϻ�ȝ�XUV��׌����G�f6"�K2����-��(�:��e��R�h��Πs�q�L=��o�zo[Uu��ėើ8��@F搜�������������-v6�_[�]{A�1^�:�24{V��n��y�F���������v�;�b'	D�a!.�*��o���3�Ȥ���kr����U[D'��իB��з��7(z%8�?fr��%'C[�%�V�
tE��4�6O��C���r��Sq���e��\넣�<P$�^kR�u��&Oe�;	���V��h=�>K��R��b(�P��Y�Ϊ�̙�����{<�����A�_;<���g� +С����uF4M��4��IΟ�@�������bZ�U�@oTu�(��?tM#�9*�����R�z��d�����R!P�'�o�p"��'��'�֜������!�9����TZ<�pL�3`�I�u�,R�zݵC,dYr
���=	��h�
�S*�̗�G�[�,�l�I�GW�.@AJ�d�������F��^�eZ�,!����X�n��u�i�2���T�Ѹ���,J�+���G���]B�Ѡ�ʦͽ�����h�}����`�H�DN���"p�J�HQ4� �� {~$���ˆ]A�Sw�����s;��T�C��i *� �u�6U�o׃���8&�s���^�v�^;8��>5r<qު�Q�8�q!�a�̞�����5{�VM̥k0�6�Ŏ�So�8em�w=���Y�F��qHҔޫ���y��=N�]�S$b�,�d�#��۠��O-)+Q�������6�=/��`M�p;^��ׄ���\����Yj��0�����m�s��&�i�	��d��YT"l��5�X��h`6�a0�yP.�Ah��9Zj�bq�W�Z	T�[��"��IU-�8�*�pЙ�S��\��
�OwD��a�N"��^	cP%�X�lJ.'�=�>�p:�u!	���vg���WFaמ�����Z�yy%����LR+ҝ�܎�3��D���͜���e�x��b����2z��� ��^|�[�Q�z�E���|K��?<�a�Z["�3I��
F���M������s��ܟ~\D���P�n����0�,�{�G�ւ����N4��c�L����Ό�]�~�E���3n�p^��~Ǟ6��ȕ���v+�9U?J�Sl��]_�YV�[`w_	���@�4�1�����UkQ�܄�}���Jk�柷h�����*G}��]��~y�f��3�	�y��$��ݩ�v��of�vdO�}vcJ-�l~���M|g=~8��ل�O�Z��"��`oNq�E��!�}����
���i���(	��r�)ٴ5<c����RU����޻�Im�c��cXҷ(�0b.k�4�7Z������Eui��AS�9������E��4X�z�n�lPv!t��D��+r�zN¸��\�M���m�v�m��`�w�a�;�� �d5�,�ό�4��N��[�Ѩ�U���\�?(E(�
�s�4�K\`����[�;�t�(0�Q������2��b8��O��j��C�]�Ph��)X�vp �a���F����߄&�g�nU��m��ⴞ�`�^`�`�<Ý;Y!�?V��0��`�g�Wk}�V4�I�� M�
�]0+Վ��81�����:$��w�A�rgK��9I�!�P��L���Ɠ3���2�X����9��� �	�k�Th"�슟C��K���Wd�x�����=�u���nɨ�4DA�󼦏�͖8��R���3u��j;2��>J�|!`,y���l[����?����_F �ړ�A���kBJ���5p�<�Et������93��?_<��;�$qVw]"���PG(���Fo����a���k?�Z�N�ߚ�\���l���c�t���QG�#�ݚ�'����UT�6[��6�>c��m8�Z�I������vɊ��%�����B�m��&� ���b��o�nR��/�y�D��G�	##�H�=�zIy��Q0��W��ą���9P~��t,��jOp����M��>a8�\:R��
�0��8���9P�iOݗ��((h��,/�<�DI��o�#E,�_/�R�Fy��� I������P�I�F���/�'bT����I.ʜS�$g7��A���C�%�cz �h�2=6��@c+sƱ��q4�gp׌���E'!��v�N�ջ��|�z��<	i�n~�k?<������[btPe��B��)�'L������ ��X<��,���9��׹Kg�Z����2�t&�Z�>��~�^�h�ӮK��Dt�R3w>fR*K��VX�%�!�矯���i���n`|_s7qȹ�-�Ω�E�����'�b�'�[?�~.lmuN��T�5k�Z���L������,Wn�:;Є�nT��\y@��(��7���5&�XXH��fO���*Պ�^Ѵ������\_b��lɪ�&���P3\������>��juN�-�v�,t�h�G�#��S�t��e.�G��˫r��L��$�)��4/3,O�S��]����x5h�������]G*�P�SͷJmI\�M��������@��#��-(��;�j����vϟ cf�o��ɠ����3���n�e�fV��dX���"fk��Xh#�P�t�d*���w���#���y0M~� ~��^��4ͅ*�^���&K��ބ��\��򜍭�٢��޽?S���r�߮�����C_yRrt�Z5�K�*FS����R�q�egxѓ���gߩ*w~Tv#�A��n� @����Y��W�Dc��C��0 � X��i�9RmwǠ%�N��EV�+�6.b�s����
q��;ݘ�z�܊�@�_��fa���s��H_�����Yp�DU�7{6s	�����X�m,���}�P�x��i�7,?3<��4ށ�HGf5f�l�~m(a�?#��nxP�����,ݗ��l���*l���Z�)/���0���"u�! <Ѳ�Io���o��O�蜅Oǃقs���^�/��S!�N̏�֮��x��:�U�KB�����nW����2ڻ�өk,���b�]6����	X=�ѳ<BP��p]��� ��K��nA�������h��h��T,M�V�QD���gl�^Z�2����s7�T���g����㴪�֚-�	9&�X?�n��I�A�0�U�
��������p -������r��ȕ���`��s�0�u4�%l��cEN!��|�$4�ygDN����I@���������$�j�-AJ���zo�񼥠9��NSm=(�:44f��w���*�I \b������!v�i�mc0e�ּ�4�iG��=l����Ox���c�M�2`o�Y0A�F���w����t�jD`�Wu�.{�T��!P��'�gVՒ#�PjT��IG:��5�o}��3ʗ���wt��^���q�BA��&kl@���wA�����(����D�5Ŭ �p;��T�y+Mҟ�!�NҒ���M.�G�:�1���x��?{��