��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���V���hS���kAk!�����tB���g�s��9w��qY!h���D��_�$r��*��aE�T՛6&
yv�J0i�/Y&���^#�(ۄY��3�QԜ�Z�$�w����U2Z߱�������I���\��S�����L�/�l�
hx$�,�64F3x��֒�}���a}+͘\,0qĜh*$n]͹Г~#Biג�
k�*��bs�`Y�c�(a��m矦���"��>B�t���z�cZ<3WkJ�F�+n�	�Z����'P���;+"��:+h(\"��[�h3��a���Ok*Y^Wky�3��(R����;r�)H�z��o5ǚ�}0���^G��ҡ�اk@mba�g���֮*��2���x"�o��v�<�mɌSt�bPlC�P���L�X���9~��̊�n��ʴ�|Rŗ_�j�iI K_ĖQp��pC�����ֆN�P�G���b�rc$B"c�֬�b!d�����u<O�y"�Q�H��4��E�[�9A�XY�M�?�T˳h�ېL*U��E�gPO��e�}�&d1 ��zQd�������s c�}.?@�BM���b�
3�3�T�dw�(k>�AHC��
²��5QE	���敱�&߅�.%^j����g���Ocd��I���*�a�q�Q�W)z��.\�^�ng�hc�|�GM<���y�C5~[��)7�O[�`v��=#a�y�����$,2-Ṷ��G�I_c%N�S�HE��/vxu����<�[��E����-!�����6���@P>F��)}:����3bZ�����ֹ��]9�#§����MZ��&��(�I	�&���ߣ�0���'�l��9�\}�1��v� ������S"RV�6 ���I���?c�Ȗ�n�3)�W�}3��v.��ï��t�����7n�	or1$~�BL����i�A�m�M~���N�Bo�{ui a4�C�+cP�e�%\@8��Rش�������+A/�5(�?�w|�?(M���E��h�TA'��r=��,�,�	�,+�4��v�l�fK%�F$_����GS6����"���p�w����,A���~]�*&�gkj:fx|�$ta���V#dfs�����?�J#�Il]���+~�4�^���A��_���Ez�{9�E�KX�W���d�G���}��(bqb��Ƞ�1u��ϴ�3�a�ȟ0=ƽ5z��q��%B�\$`�J���<]ݍ]~?uT��OB��a C�O_H���\�ʑX��&�������:!t�Gy�оɔΤ9��&8�WU�b��>��T�p��UC��6�^��Xҗ|~�Y*���5ًx�":v��E��3��ٟHS9��Q�&pb�y۔=P
�L�����d;��熎A����"�����骑�7� rƀw-�L�8����1G���~�6��ܛ�10�c뺟C��=��s��x�g��Awi�H�a.u3{Qt]�:�15;����F�Z���H���֞�c�/'i1 $V�D��P.LB�ʍ#��ӕ�$�dm�s<���~oU�+��/1Ӥf�O��l�ۼ�6���5�65xa�����*�¹?>��D��[4.�e���^m���{vJL�{�lr��,8�]X��/�	��Kl��^�O�i��CMϾ?�VN���-���d$ͅV�OS��-���C����茷�]�_�/^�a�V�@w�kpYʪ����Gd�j�u�SkK�O�`�ț:rox�s&o#��܏!:�4&��q�ԋ�҃�Ԛ�&��t$��ڼU�	O���u)��BT.�y��-F�+k�xİ�7��:�l�n	�{��TKo�*��wo~�h�O�k�i�t]�CnWǧ��S�x��SiշA���,e�ĉ�ע�m��b�{H���-YA0��6,�^���z�`��߅/�`f[=W�����b<<S��֌J�@���	zun�eo5�w�J�:|�|(k�[����#�%�PFZ	Z�vE0`4�!ȻSNh
�T~!:>v���*�;x
��G���M��#l �U��9�S�eOt+��ڄ�e����Z��k���wH)<v�|CLf�W�Jŝ����r<e��!��0��e������vY]���}�5E��e2�t�`�v+h5�B�$ Ɠ	��]9�CӅ_�蘈�e�R"�e���q��o�N�����wM���5�#�#[�����zq���k�ЍJZ$ؘ+o�!�������:	�.#�olR�����XKY��Yz�4��a�c��w��K2D��ys���<�B��*�p乇�J�_�+ �(�$�U����:�zAq~�:�V�x�4����k�ӵ �U�;�k�k!����,oR����UJ+
�v���刁�̷"v|��G� P�д�'Z�R��'��ݣ3V�M���@A����d�y4��JGI��a]!�;��9=@�k��W �Yq�C�� �[`{~[��͑"������Nk/A�#OH����g��W�x!
�O��㪼'U������]o�,�a�.��g�f�l�T:QH-}������,��~}�����G;��)q��ڟ�������X��afr��(%�����>���A��B���yw?�'^l���������HR�B{���盦*��X J��?���_�3#D;ۧ���h�KEM�Py|g��ѠzA�rw����!e���0V}y�#�w��GC�ؑ�ǁm�Y��$�I�2<Hb��`z	.�d �͛����cTg� ��j�eW���b���%�|� �ܣ��@��]uczQ��,ɂ�L����a�j*n�̤���7$���hU������������H����.+��A8ͳ�`Qi@!#3R����;E��C�]Hc����)m�	Έq�CJx�g�T"k�c|2[<T�NF������b���i���C�� �T���Vj��3։�=勍�|�ޥO�?89Pb��=~�\/�Z��a��d>�F�W�9l�M�O�f��ҟ�^Lh��89��F��n��7C%��ٛ�6!��9�!�DF��tJ��XG�j�;MF�@�(M�����ǎ=皠͍(o�;�+&�W�q
(��ȳ�DXR?WZ7O���~�]�J̯�:,��Wt�̸���:U���2$mv���8ȕ�U�<�5]�-3uI�(⁙��{h�*"�\Rh�<�r�Mq�?av]��P�J�	�s�6Ǐۋ*m}�IK+};�>j���Vt�V?}'0f6N�:e����T��1���&�ُ����iq7��G�*�e\�,��3�U �����9�>a�R�A���r�E@�ʏߑs'm� �BE)�Ov��c���%ܖ�~��xd	n��{��͟�v�U+�#*�4u�K��"�1PQ{1!AsW��丹N��^oנ]���Y�%>�L�C�	o�Ple�gf�>q5x ErHhZ���XD�������F,ڶ��%3�q1\-A3{��k�ū�u	g��x�Z�P�]���Ӥ�P�<4� �I[�]��&=]��(B�U�m��nxf��Ũ��o;
ȡ�	��:Q{`�Mu1�]\c��(z�Z,���_�(��
6��$����Ie[�0?����6��NB n�=Dqaxf���?]��`�Q�m�D��ғ�0��"HbXM�������w)u��ў��j�^#�{�̄jlk�V��\_(j�H��"k�3�/���Ìw668��s�x=as�x$�)�68��=.3^8�</G��BT2 ~e����([�D)�v�=b�[h��D�oY�&F%8t�qb_o"��N��� ���	� ��\��/|I�Z𾶞&>tM��_�*�ә ��P
c�^���j��M����B.˓�H$Z�do:Nm̠����[��2`qf�����Hqb�c}��|�K��[����i�����|
K�/i.~��a4�X��"ǂ��n:��n�-�!�,'D�C�!����zO�£	��&�'��?��]
�l���
��V����Ź=.E�e��vJ.*q���_�=�:[���<��԰����'� %�Ϣt�����"��mõ�dA���~�nD��d f
e���
���{
i�QX�t�[�L@�;��쨗j�8{�#���D���\Q4G4�@Hd����ң1���H:�T̯�x����2��������\Q�� ���}r�f�w�Obm�V��#k�o~Z�^��ܐ�{=�,����f�e_�C�ǹ�J�`,7ߘX<�֦��8�����˸�q�t9
���+��t�E��R�j(u�$C�c�̙DKk��9����`�%!���d�t�ފf���'V��yI���S���494�ۅD��0{�\�h�Q��H����I$T��	�����໺ w]�#Y]��X�	�B�I���_6G���ݺ�:7��j ����gD
��'J(R�QM�O{U�'7�k��~�XUf-}y+U�n���}W`��'孂��ٛ���	�|Ō�k���}[y�1 c�P���ق��*��~)���A)�Ԥ�}x�/��SY�9l��k�q��:�;8
̀�Kkm��;��YR
]h��0ы�3�bn@��;[@�)ۛ��v����Q�L�u��>ڎu�����U{P�Z3��b������-�ۙ*�ߓ\~���A��g ����5����x�F�ǆ��v�۪���d�J�<���֎e��n�܌��>iX�xA?p#�n1����u�r�k~US,b̢���C��ݑxy��JM�5�JZ�0"Ց��3�}�c�I�}<!b���iw�~����8��!�mI�e-Z�V�f������Iy@�е��i�@�H�g�G�Z����5�,iɩ�J�Va$*�e'��Ư�\�{*W�t�DvEϋ�b��������-�xBF�����pM�\�,�_.c�E��0�Ĥ��)Y�����-�2��3�0SW�*d)��U_�8� �6��޷��,E�t��]����yV!�9��p>9���X*�Դ�u��_��gt���f	�ֽ����D������֧4b~O}�,J�h��1G:L^)��̩G������V��c?�����D#��/$`�s�gjXx���n�U Ϣ��'�M]}pbk�&O%�Jǆ���C�&-h{����O���Ig�O���	L ���ȸ�5��0��N��Dmj7�����-_�0���BpYBu�F�aܙ�]sPc�%�%������N�i���;O������{�6�;g�zD�1v�����*�A*T7c#$�Yr� �9#�V�
W���m����{��ZP��x�����D�.C޻>�5ʹ�(ɟF!��ƺ��m){�ͩO��اې�9��2[K��8�;�CFZ�аM�ǈvCr6�?UOXʛ���vrt;�j���yi�}	�k��K��g�+�ܚ&h�M:v���J�sT{Д5tJ�&��� �4�9�#��W'���sCf�hK�[�}�!������%�[�*&����r"@6��A;eJBͦ�]�ޮ�y����^�����V ��<w\�� h��p���j�4E�U��}�\s�[��ءQ�#���ѹ�6����2�g��yR`�:��\�Hs���oT�2f�.̘�0	sXR�jP���%7)P��oʣ����/�2x�'�ZƎ�z��ݳϷ�fW	l<��\eS;���A[����?����{L�y�H?ޕ��{� � T��@�ǂcO�\in헕׎��H�x�r�1G_0r�5��%�y�����%x�ɪ���*����&e���o^��О��%���8_B��Pա����J���ZQ�@a�?�ޠ{%�g��<_���n���<!	��T9��Q�vֹ���,���"R@]�"�S�V��L"��=�4�3,��?/ LWl_ע����t0IՉ|0�ji��G���Ḙ9��gL��A.���(c��V��-�$�רog<&q���q�i�@9��{����@�X�SZK��6S�4��z�"놛����k����]���fy�������o�  ��8gE�.����7�6i0`����4�W�8����o�=��늂b�JX$eΨ ��ʴ�aH;}��c��
���3RB9��
����2��0���vSS�gN���b�ϿO�%w��oy��c���\*?�[�e�~(Fk���r��:@ �i����C<�A�q~�c�{���-�5����;�	��L�b�<ej����l�K���e�G�{���4j�6�-!����}0���4��Km֢+���#�,�w��Х�H�B8�б�{5�B���v�6��o9{�םLG�윗�l��S���P@lw;�d$�ɒ�M1��v�(����!����4���\1��Xn=��#�5� 1�B�s� �RX��給�5�}�ŚF��UW�t���jI�H=n��/){��O:'^�?�͚"/�nG9���6����A|���Z��N4j���@g'�ϒ|��v�A����&GQ�Dm�o��j����|�-��NB{	ՙ���⻇�Td�L9c�qΰ��Wt�i7��yϽ��$�7kQ9\�c�a��^m~����W#��3�w���'��Fe���bpʛ�Di��*�A}!CRb5lY���iK�9����Q��޳�U������C0l���#6��5޷�svU���?V`U�y��y��"Ŏ�vc�ap���<*���_�\�<�� �1@�P;��9k�(�C��� ���np �ue��u�CU%���0%E�.�]��`%�j��wG�s�UN�H~K_�`�اvJ{[3 �'�I#G�&Om!lC����h���*J��C}�u�e��n��i��