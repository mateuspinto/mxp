`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
cWRCia867n9foA451nYwHkg0/2/o/mxgAs2BSmDmV2dxLysMKtl900+1KlYkO4prhmfuAOXo/SoC
OSlmDh7U0IvaPCSx/DQpFZiPb8llMijSCCw/Nc49vU3HbDAKzF8uQTIuY0liC1cZ/2b0S4PQTDI7
dz3fdeAGhPVijBFJLYd4H1MVzCsUqvGVLp34bWXoJmbbneB3ssg+wcJunpS5oMloDGO1zY0Bmw2s
0dBbNUMD466M1eRQrzFqJ75i/V4ifyNv56ZyETcGRX9KOBteZY8ukKqJ/j76GxIPItwe8IYuhW4V
jA771kQUcZrGlZVZYc5id+krrKQiR1362WQ3CY0CBrQqqynmHaO9rwUuf6S5oVAJYD1xEwfVArYZ
F/1hMoZSD6Qws0TdYM7TGfpnkbYhnS2bHuRpHOMhwjNTpRCr1d2Lkao7AiWgZa52i3Kv7gi13/6B
x97qaY4eoMKGbg0Xz4yFNwT0nWbpXjsk/oUSIjVjWJtjudbbgmYeFhpDTtRQs7ArOMIK4iOqA0EG
W5jyXkS8z6bArIRCvdCBEDs7oc543M4q9IkckvfG+F7Vz8TwSXCfQm4XonXXM5mOILWMIVeg11Or
ypVqCRfmQvGoTwhKPrynEU/fzm7lh9I9n4e1eWCNSb+TBwfHElwtQxlUY9s45ErdMoBRluw7i1vb
aidTLbhS7IguvTMY45Zv8+rXkzXpuvQwth0qYfkEU3A7Qaw0q90THjR+kDLJ2dSesAkcQgdO0FTG
53JLeShWOtuLN3lFrCzQJIx1bMz6aGv4+hRZA4j64GIgWkyAUwoooNtow3irytkNzCCkOTznAxyT
GV5lPqPrdo3sH+cpX7rCx3qOm8KdoRekmo5+KPPgjQdsv2LAh6UEyOMF2jak2MyIAIczqX/sghyp
aTq8UUiVTtgxmltErH+xueKCQn7IcC3wXsHDh6PuGz78xvmVsxHxmDwUeNv0h0EPKM1JJc8AVPKn
4CFyuT7yGJa+2borW+8zeTC0LZpgrofZ1I/jEeHc3UXlD/GLF3Hz7PVlowy6rdiNDDsxtOjohrbu
xef4U1z/pMzY55zOuBUSKbkznX1fUhtHgAfcPQvc1DKsZPKrckVFxJEwMTcJ6rp76Mg5KQZvphtB
GyDJP5j2yal8ZW//WmPmOfvZvAPBliXmNfScVf4hQE3ow3hha1CWMzmcCZRsTRzDOmeP0OK3CfV+
LuAK+Fr9B3yTNBi61gruvay6jqPN+bFoK0JhbqFXm0duqT/8OO1BbDZhH+6duGkNtc8euUQlp3Sa
xL73W0UdGsnkSnmXkCb/pcDeoNEYflS9bBuMBFQuipgR3wEK0UZrXcDHHcex6NfKEXoUX/g5uzhb
+jBWGV7eyUitZuI0znzKXJD6YDYM1OV+tHJ9f8Y2eLXSD7cjc8HArQ4WqqSL+8XFwOFVK0i0C1zB
jlzRz5Pf2IUElssnPzAvKxC9V7HceeV8lkc9Af5nOKAnz0RRRfcXKOfb1cDH/qDI2akbGe6Iwz43
sS4Y46RgKqmAaQkfffudBI7GP34gaIx+V5T0ksoX7gj3vkgw5WSHY5HOnrQi/ssChiJoDvynVnGh
MnLgjZjcjVrCKsiBq3KLiNC25OxV7A+yYot7pEN2vaCyDFVEochsuCnbGqC012K7zrwxv51bnbVd
3TUlldPfy0W/GoBropS/75zsgbHNk2EcK5PCeAbllot81Yr+vU4dGmXsbm7mr7AV6DH9C6xH8cfs
PKxKxZCFXWZlXAZ5QaKJ/LG10l9X3qfoZeN6AQXzXqGFLyBOzlKaGQ4YFO5RyvH7uotRUF0OLX63
IKASjjLaVwdEWHYD26z/sz/Lx1KHuCpsGH7/NpAei49m6QpxhsHw0qnDOMQs7SJ+JRc7K/tFw9lp
Cp1AHF+bxaH4s7jxNhKtuEpfRscMhsIxGbKgRUcwGuL7AutCa/HiZRpUS5lYZsOWDupliFIHsA1I
DwiTUxn1aMizzagB07YgTt8dyH7wllTX9ac4nmbWTnSmvAQg8rQXVOr14Q1DsYhlB36y36bo+1db
DGkBJ3ZbKzZY+wCiGqYa6y6/W2rtVAK6hgG9P2FlMlWwjrPGoT1UEByT6SlgD40cd315f6cRXIl4
7mWzfTA28btkIIuC7TY3JEscZ50aR4qH5TH9NARl6vy1OIqhZ3PcGetxDOwHZ2o6u0JkQs5nkQwq
Jp/jWe3eMpuickmnPNOtrr1gka24nEbIWQkJAAgdhhRKJgsEdZHmgoLUk3T2oo3/HxD9nscV+BRo
mAvWqBKTi7CC03aernrPDoTJAKrhNgJucjXKyQsoVIrZKYeZco09mzl0ighs/a7518NHVZtSIF6M
9mhiQv+LUWwowKKZNzQK2zK7oA8I1AF9IqCMR9mHbi4PP4L7A1dfSdtYCWnz5y7fuKXzeWthPQ8+
PEWYUAeK8IyRNZxg6+zeRZpXuZ7NHNRZx+WF1/rzdiP6GwDNd9IdMXeJg4xTfMQcioBK2Cm5rdSn
9/+4cEE1u0JGUV7Be22HtVS9Qmp/t7lMtnKi76Q7daRp4ERB/4aFSKfLmMKggFXawcrj2Os+p+jC
SpeEEFGHQk9yR0Uh5mDOc/0gta0MLJVa+UwuAQPJ/KWPmMXEygXTgjNPdvFQy+Fpuv8ZXSfSF9bR
LyXDb0N8+ccrmu1BlGs8hNxv9quD5EuX+j2tnKOMg1j9POU/CV49PlPz3CpdwJcOKZKvkBLUMNXH
m68ZWzukBT6BtHBRh34qd+vX+OujrhhvYHxI0w/B0eU0/c0dqzovJTfvk3AAsTz7t04+HTRfp3FY
blBfeU+gg3sWHpofP7glYjc7RlDWBomsxC+QJbRkx4dClUlY29rkM46bUs/3Fs+XCurw/53wY1Bn
E4IAVFN2huIv8MdoqGcPmwIiqci9LjxZ8XR867rJgBMuK4fk8twpDfFX1ge8tsgpSD1hZY5K299m
J+ip0XcIA/UJRWLGncbIDT5rQ9NH/k/1kdKTgutdNoKcMFCCDbzBOoGNoHIMVa5jj/VDxrHxF12Z
2K/sI9W9eV6AjwDz+lYkbPz3jdOtf6P4gF8B5EnXgC1lxXt2F0LRovBuBhq2bOwHA28gD/8+X/cW
B8+OKlQqcZh/AjdsuiLOSvNcsiUAfQpHiPhYWrLHw0jB73kmdZYgTEdY6E2sTwyWKcAmZGHD98W5
z0wA8v92AzeZEtuS19Cbq4gZB9SmOEacc/kfkEdDGWSYknsLVkXEEWJn9Az51m6o4A18fNDzpSOy
CwvaX0A3gEuqHwrfCAN7UaSrrcDz9xa38hwY1X2Tkto/LPheju48UhkqBHx9wzs22+vg+Uw9Tv9f
1QwlxS9luLodWdR0AmOLVbKN7n3A4imnyQDN6Yg2BTfSFN3c4/p/nzTolO/VJ0lDyNhpmke1yoPL
betzWHfFJPFkr+YNXoexYj0xacCXthhgea3Q/MzYjv/y17Fxs+8Wbs/efqlFO2+k/W3bdemusUHw
cPh4FEQmz761DOe2jLHHV40FLAAyEb4wisahK1GPsCSkVVumcyT2bhFtU0luqMipzetpPHgPwMW/
A/shjRBSoENLveT73ZmfGdxz2ed+BzFlzeP+RppPNrTyrnknd9OUGkBeQfvIs4LyFpZwA9XJIsXs
BnZcZQPkw27/RIu0IsF1825aADqc8tUSUeoUGDJnnFk/oXk+oyKoZ/g+lwsJ+Nu3K0MCmKyOYwXd
WDf7ygyP5lQ8TUQBhvN4l01dpxC4VuaLD7KbUIJ+WpSjrynJEYhnT7NA0BteElNhQFow9FniZ0tW
5Ns/oUmLMTMCFpz/EwMYI2MQD4AT+fTzQhLlelvwK2R7qIL5wGIjdd8o1BoGvyW3S4q09N6t3q1U
g3ybcQaw9JibedYweOdN3uVThO9uPx1nRPBXnaXgzPWlFCxDocx35ET4THtB01ZsRjeuFbbpyuzw
VU2UBNXPKrwBQQVbXfcF693jiLDFW/CnJEROqlZ7jyk2pS31FOgL+yiJS9h3icMCbUQkJ5OThqDr
A1wmp+twsDb/xNIbo+RC2sJOOQXx4WqTMtq6KvAwsNUQb5BuQSRt30v+jMx89gOPWATTqrhT6uq5
ZY/b13urlKqFTVsmXOdL3epPYfVQmT0CGL1bOLsH3+B5G6qLI6uSFXT5lSgqxcbwAi8cZG4gBW7i
/PZ9/iTjfZcY4G3CK7iDNf/ZgleeDTgvwSzNHXpuborShI7JxwoICyTsDXUli741H7Dl+WcRO4Lx
c6T75rk1PMf8m5WKq9fcahdXRHUlJVV3xVBKC9TdOiMWbjzIYa+w4vtZa+JzxXxLZTq5t1MEarK0
ZVFmeL9y2a6fPbftoe2B2+p4iFB3fm48bogyTC2GDtJJP0dZLi/3mgDgItmsSplc/LWvoLda0awo
fQRsBJqdB37TZ5NVIvYB784U4MCn0/3JRfe3LpRueuqoh494je3T1NmgnOqsCgucfrBLRjWkBRnY
0DCNJfBeEHkycHd5ghq+dCtTIn1MQXQa9ebJj3nUIHQ7YOpUgHKiXVHhupajAlisLYm13dBqRQr0
OYj41iHris9vXnV2631SfzY5zJGBm6WkAcgPVGAr3QKSh0mU2TVxfgFUnFn+Mwqhf55wsRcyBZUO
8cFcuR+kQAF/Yz/u24AdWQTix4BLrIloNGDLc4HA60hZIJmSaXwW4OxP3hwwxYfZiJ2W/c/nlq22
KAkai+lk8YTS9XG6DbV7hF/EypGakSeMDsWBVLSTZxEALaPmDrtzA+u7NJmsai41cvZ+C4hU5bbw
jpk1ZtfGQaxhwOEBUIRVaGHRZ3H33D7VT5CRE+xaK5/0hjsuhyB125MOH1GineXu+iGzIbvRrwcq
uAQ/acFQDLtxe92hsm/7TQ/XLGYdDlTNx0W6Z1RNjEWDC8MPDizqpCxmOmUwsiWZdR60Acm/FdC+
przNLfPZNl0aKRr/W9UJcB8Gl6J90cFfKe/kLgggjEerNhJRpmPI8KWKWttJpHy6cP4tRCZISXZR
r+xYfRM+d7Yr7+Qi/ejWt8Zpf1waU9O/k9v5cW34n5TuN9fmSQoGbwEWHL66FRpY/FgQYD9WweHu
nEsPUcMgoUQ4jNTvRsIC06/h+R1FyMesM7BMJQFk2etQV9ujHDxjXA3HUSZxNEAswN5qlXFYaZt/
Ugh0uc3VE/vJ/C7Gf1FS3ry2BE/vZnWd0I2sS1+RcCwXJyFR08fby9DbRZUtJf9nTtgpmBnpcWbc
S1+mQtr4zrBBW2DidTGsnSUWmvhYb/02v8tmBQVDfOgB9emHA8GJ5eO4TaNlPF7VKrpAJfhdY9nz
GZZ2BXf1908tRQximqclRj5+ocpbgGrCzojz5AS2vh61dmqh1Jz/S72XEAy0loA84Agk/N0ipzHm
Jf5Nh4PW6XmLRM86vFJSZK4UR3DZUg8Tj31yGukFbRS5Eb1HorslaEOKMVFbUegyrjlFtsvL34gN
08wekquZxFvj+UrTWhvwquRdiNbiuVGJeEliJgVK6FM0XpuBN6TAqtPvzqV09Z58PC8lc8cvdE9I
3qUG9VWM12YPzjtubhA5FhcivvdsMNaWuEewE6Vp1uQGSvbYy5ItcoFty6Bf1faa8VFIu/Mm9L9W
UqigygjYmw5HVR6aMLGN7Rcm2QHxbWachLfdNBBEseZ4YODoG5jKQxkmjiOo7cuICNSXldhVFJHD
HJAeNtRkePs2y6fgnjB9gHJQC2svUMsVdeMuEOugCkAwBuVggirSNG1SNmmrzBbkbgOLoq2Rwynb
kUHSPNIvg9mFYCHH2vqN3ADggwaTXifGdZ6XhaBYNngiIqmCTcb/ysczDWyIwTRcj0LMmohBPPkj
e9wfCgxkwnQYlf/lmHQheI1obDq+u8RW9jaWzCFkUxLN8DmV2n+rbFCW3zcDl65DMlbDWVpBgibe
uR0y4jlDDgUCk0V49dQI9EcduFW2lhvsd4yGP2QvCmD/adWJXZ6R5ptaUWvQwwRkBpiPiXE+0M+R
gHlWEIjiI+dTrL5XwhCWoynxpQ/l8LUtfXh5uY0tKpZ4/cZwuDlKDkekUNWj+5PBsjOn3a5xly3r
L/18FWdjlcIRqcWN9Kixpa5+gpf7FqPA4rowurRXmV2EOjHdxHcb3Nn5oOuoMRZHiy3DqXePdKJE
BPIw6CDAIUxQLNHBQMJVppdhkeHQoARms7Z4Lz/lQQ8hTpHdsh/AIJe/J45tI1uo+GOzP2hYqAW6
ou7m+ppktVEEU69d1BJpi5dTUiAkqJ06WLHiF3liWgTBiCSaJqAbG4SS2hmNrihWpmN5WOVtktIa
/t0+uzvF3RVgHSGQUde9YsYuNNOcjCPVR+qXftkMUNpMXtNeag53kwu75PTu58Lh48lFHenGfEuM
4+4IIKBrxzMcn1vCVRpwyUjOao0eyCXT7/Vu0JoUw/jqepT/oJu+xxvBA4Cg1B7lPe7ENw/p1iGe
EiUIuZhLnD/2N6qm+VvGLEilhI5azgcvosne18eeucNeAUYX1ounJ2WfMepWUYhji250e7YMMK88
SrbBmo2fvHQqunQ47ApEAKyVlA60AhnY70E04rnf+NpeW7/qgp+qTWwA9Ny5AZt0HXHgKotAfjzc
eHBiNRmNA54vYO76Q6HgPxcnsY5B9T/0R7pgJNtzTyK6OIT53WojxY2gAkUjxBbrscUtoMHNqbXI
Abm8Eb9FOjDZzbRro4sbkxSQQOaibgymfH8XFUDupV5l9g3dLiioWHlX6bdNHSoD3Mms1liDJvHY
laBVJbzaIXbn7yJioVgIxT8+HC3pEJnl8iP5UoB2FenltxRX81UTcEe303SP0hKKYMnb7LYUzQnh
mXL30x+QSL9okUA0tQhgwVAgTToSKwASYvOlCX1eR8HxeXGb6JTqG5CCG7s3ykz4zJPbD77kXbWt
WdosL2QIA3NYJNnmu83qUOoGAELsdzr3EDKERzYMAL53QuPk3Y+O9nmx06AEqC+/mKgEkLpQg6kJ
C9GLkyYojQUqQ96NWHbIFJKPmOi5Fo9j27hvDWye7Ct9ti/S2xy0qrGskHxk/u6Fz9OTo/NR6AQX
+eyDOCCqkFj1c5OvFTCKv5gK/pfCY1fX03dbQkNXx/UE6uh3d29cDNJtmmf5Itjc627fWTpPQOk/
MA2oaTiq02OR3UpDC2OGWBRzNmwwG45SS9aP0W7WTkUdwUaEvwzButAgiTT9sioyCtZpkCWy4zua
p49vKW1DeobfiPoSZHIAOQKX6axPPlN30n51tl8GXW/Yl3TM6UWNhjHBdJ2VVWqKVfPHPxDO1iss
qMFUca97JRos2LfSLnwMqOOru3PXB4amGHFEpTfbXsT+1v3wcU0gSZIBvWsJw/s5F4mfdFgMyFZY
FsAXDwyOH5Yzv6o1RksqVCwHogo1ZEbKr/cVIocCtQZpnk3pTw8bs9lQehQEm6tCU4Uv7gLk/oGD
0a3/RUnpfHBCQzGm6B/lYXFZTci0U4tacbwAeI9h5yW4YOWdEaCVB6Nsv67VN/ZSrBJW3iCGRDuW
zREavu0MWHRhdgt61+/7joOt9G1+UZ4qZ9wnPh2WQmJ9m/06vru3nIj1+juqNtQqttVJV78Hdh98
1Yka+ZWn8qvzZhUha2jdMFuyZdhBvs6xYd76U60vY6rP3TqJY9wMFgEM4/Edyzdevwn2DaiFTZ7W
9ao/dAmO5KJZHihQpfO23kK6xSljQ/mYvIEP+hF6HjcaUxds4tUvs8L+3OpYPDerPyH/TKkzDG9m
2xblQsRVxzUuftn5V+mpTFZjrrxr0fMiBArke7Gqal7BQ3Lt34fsjpscP/s9vlLpe3squNh6u+0v
8JFeoQeDnwgypqY5Rp0xcLz9pbpwY9szFjMlMMIiPNKwzUDBFrFL6Jewawv4dm5cx2rWNCnhSg15
aARySqKthvOvtaq3XM5RH2eub3RqsIApZ6pP3fBj1l2XP3ro3kD6l1sBX5DQ3qXBPaw3isCEPz54
3oj+wF5w6dbXrXcp8mbh17QiO79vzi/fvJzTd4aZnreGiQKQ9B8oQjbxjbW0BKaPfOu6wkX+sgbO
4oe69Mc8MIgWekcP3Ziw3sMtz0/37kVmrMutbEkaeXyIu/WfGP6CjmuXz0FkOmBN2zeCqWF6xfll
vOfJpTf8aypHfPiEn6REUfKdY3d3qg/39D3ps+pSATHWuNmueAtI5quHyOEzSt0C13YhunkIsCEH
zeggQ8QehBVqSiR16oNRk+thjo92AfthC032l6ijXAuTSGGVb1982NYKAmBAUTZSqVi2UWuX1APD
/cCfk9ytLCFyarC4OjxdKahXUCITLdQUSv0Rw5briY8KSRb628RrHytIi+kJcKbDh2xNfWkRaS8v
QAKcQRdEXx8QYuazB7CYBYBS7KArHNi6smyfdV5rvghK3991l0lILgXsfLPXbVcY2bzqIB55Shyw
a2aWr24jFYxjlfKlEDW9sCcrt057Y0e11i/hVoWRBsio68TctVntldzCF8N25r1uKeRO7AfDJeos
ux7MfbQqmT1WBBlofArPkg==
`protect end_protected
