XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���FNpj�ڱ���^a�̶�$gY���2v�j��%�ݷ1�T��nz]*j�I֢��t��z9Uɡ��>��{<o�Y>]�i��^8�ɒ
gH�Z|�Nq��(���+�3���%󩻯]bȥI}�C�x��=�_P�
V-!	�?	&�A����T'�EJ�
FI����p����<4Ю�(��W�Ⱥ l;mt ��~���µ4��ވ�R�Y!>��+R���a�d7\��'��ю��Λ�	�@\y�=|��`�G�r7$������*F~6�Af�՗�?�!����	}��j@(1�7R�@yr��ӵ7CBT���ψñ��$(��F?����^�]�9�ܘ���+4�{�/>�V��r����q���<_4�q]Yq@*�աr������t�(:N�`�%� ����s�֊O��A��}�Q��.y�@�L�V93|`��3Z7-�����=^�p�`!�w���G�z v�ڭ,�U�:�%#���^]���S������t��8���(���!R7���[�H.i���	>jҾ������8�@~D�_N�E�}�nmvkN?+ �+(�n�o�}�)V.�/��]׸���c� )S5���-����u�a��/v�X���~y�����Ῐ2`6�G�aK2�*�>I���3��r�9{*��#Mc�e�lk��!�l��}��q�X<fP��߻yfvv�����h;C�ȍa��(���3�,��� � ��3��gR�EQXlxVHYEB     400     1e0��k�g���1@��S����,K��'[$9��e߱4�����Ee�0'�-ku|�x2��ݣ��O�/Rf�<���V����!7�Xz�S�C˾�Μ�sF0�UZ#=)W�I10ƶ����B�=x-�����uE� �#̸S�5��5��:NSD0^�rM�ݶ돴�2׊>����O_ p�^�������7EM��2���yAb~�6K�"����=���Ru���7��1��5IT� ]�Xp��1Wd ���(��t����D��q�k�-\��֠����[��Y��@.u�s�|���M��4m�$��t�$�><d��t��;�d��C�d���H̠��;�4W��W�1֡h�7_��1	u�(S	�Z5�1wĤ�1�6�_�¶�e!G�&��
I]�{���#Ŕ�&�&�`*d���*��S�n����^��nk���8��P���'�KhEg�?(E��&XlxVHYEB     400     130��f�(�{��;� Y0\���"u����9�#y鲵�i(h��P/\|.�Fg��� 穥����O!ժ��Y6�3j��5�in��
&���j�
�a��B=R:M|Z�-� �'���8�������*����O�Qx�G5���h��Ĺ�����8^��0I���u���:)7*;Q-8���܌�翀�LX�B�@[(A� Jh�=o�1�[��%LǺ׸y�	fV�e�-U�xzu�����g����y��"�B�*%j+�����f�T^�'�kF�-	q���RWA��o�|�/ X�XlxVHYEB     400      e0m�D%�y�4�v�M�K��Ae[�QT�p!�������s���Y���`E7Í�;=�����M��`��ʡXz���&�C��&�̑�8�evܶ��0��Oh��Cr� �Vħ:�rC)B�vw�nS"uS��� Mgǈ��<"�c���㌶x����l�?1&|`�'(pt�g�a�£�c\=/��nOudS"j%�x@{�צɂ,Ղ6�\\��~; V�uoXlxVHYEB     400      d0�)f�D�a�Ͱ
C3�L�ҍ��'2��.X�:v�%I���?��YL�NI,`>�L_.���2`:��ܥ+��-��i���͢;Z��+Y|2�Z����{s���0���F
��E\M�e�V����ĳ�8l&s.ͩw
b	o�͗�d$[*O����a�@�&�L/ZvM\ϖ_Y�B�7�;�� D�E`����_�XlxVHYEB     400      d0����d��e��}/'�h6 SA$����[���06މsu�-n
n��u����
�҅��<ΖUIWv��Ӆ�?�S�˶����{�V����r��9îq$k���X�yt�Ơw)�w�$:�n)_d�a��Z�y���wx��~.��&����m`b�V�j<�Y�`�i���/�9��9{m9#aGh���:� �$�a���觯��J�XlxVHYEB     400      e0�Z3-�����5�{ w�OQ��a�M1}�������r�D��|�d(�D&ϻϠ����ٯ���t;񀋮"5�;�/��"�j�T�5Jh��pEq��dq���x��>M��]�������������ܥ��~:���.9k����Kl��KΧh=�D�=W�X��fQ�r�Z�䀣�X_i�M�e;;,�E��rLƏ�}��X�L��?XlxVHYEB     400     140���jWw���4�>��9Vk7�?|�!����Ɨ&鈀�D譌�"�.	9��w��T��G��9\L�3�Ԃ� }蹒p7�4�a�2zM�1�M��C���Js�a�`boҲ3���SZB���_��L��5k�K�l��^kgk �Zb�G���	1pb�"Y�h�s�vk� �;³�̒<��5I�1,����V��\������;+N�������`��&��|��D|��ES�����.�q�j+#�=�֩���B*c��Ϧ��h��8���h�U��$��� �j�����;dEXlxVHYEB     400      c0~��*�A�&��vk_.zsW�pu���4o+��_�2�e�djn�sK=�`$��jF���'ӄE��wg����|�.�a&Wz#�H=h��d�@�.��
P 놎�I�$�a�wN�a����.E���?2n�cӌtÖ]�{��GX&ʝ|벣?3$+���[�F.� 8עP>�jY�P��,<;oVF6XlxVHYEB     400     200�$�T}���,��c�S�����$��Y�;��;��I�V����O ڍ���-s��DC���&�|���c�*���#��-4��YJES���������D�v��	e/X@�������/�ې�<��6��k4��nc�k�,�����[P?�gq/�'����o�XmoZ�N� }�1Q��2ih`��qE������|�]�A��E��>��
� :!ګ�)���lK�'�y�/��9�݄z�Z��@q����=����ذQ�ꆢѥ����M�M�����oҰ3Ku�ă�\��TՁ����K��)�r�N���p�?�_}�vP؀m��Y�G)xH��K��	 <�����:�\HJ����Df��%��oA&���&�,�)��0{��� +:��Sp��A5�])?��A�����z���, �����X�Ĥ��z�o	�	�P�D�h`����:n����1K�<
B�|=�+�B�_�!��/�p������OXlxVHYEB     400     100�!���0!����Z0�l�f����`@�����~��sL������N��~��� �2�<�"{�E-l�8�������h�oe2QroG���C����滪ٴ���/�m��Jݬ�y#��J�?�h�t� �P����D��/95�6L�	��U9��6&#HY�a�L,H�D� *��g��z��LC��``���NY�VT�n⿥.��s_�e����N��o��q�C�b�>����wy;�^�����+�B�XlxVHYEB     400     110gZ�5g>��ŀ�B��.*���S���ނ�	��;�z�b�!R畭a�%��.�E0���3y��_r=����-���㠦G��̱aL�	���ܽ5q`��S
"!!?������LQC���ō~��t�?�ǓT��ބ(���J�1�;	���S���-BD.�����,����]z
T�h�����Zӂ�����3*��l�q�6��-2o�a���?�*��݁�ىer�vm���K\��`�9��\��4g�����˒^ٖ�4)�0�Vk��XlxVHYEB     400     1a0D�
��JjU׋��8~b�`�D������ڡW�[��'䨖�Ѣ|¼�� < �X�����,�h��-;WŁ���7�	��~[��'�{��E��EE�\+�cL��M�{��I��δ��w���H�`��s����⩀�De�>I�H~��*�S�{B�c���H��H����5����IT�xN�h�j/�v��e)�y�sx��s;��g�J�c�z��v��E�5$�A)�J@��ܠ�ou�C��\�MEY��LԴ�>V����-�gR�%�LL�++�a@;>�@[ ܼ�O�;b
ʲ�lr3�d��c�Hr9=�r9q���
�Iժ�Y�}���
8L�On�zĦK1=?�)�/A��L�^Er�mE�=��x©X�(�iNK��m���'*罬�XlxVHYEB     400     130�������(�7#8g�M�u���\���6��QT�v�l
k1����i��.u����i�_�a*����<)H_���Ȩ˓�6^;��|�5'I�.ͅ�MW}�6���+�]��i��*��H+A��Q8�5�0]�B^�RC���'��&��0N�|K ����������"������N���꩚H JJ�(~����T���-e�t\�!��,R�Ѕ��WM�&��,��E�N��^�	��>���5�����O#��u��V�%i��z�)~��Q����&�V%�@�h�2�d��q-�o�XlxVHYEB     400     120|��Я�q�t�+Ua8����U�8')Wx���J�i!6F�ƄݒT��q|��0��
�ӈ��мp�<�n,�"���Z�U���<qշ���S+]��x����4�z��lcIau���gR�>���a�l�n�bZ1{����#�dhE~T�%�Pm�.��>Z�e1�j��u��Qe�Z�*�W��"P�T�2/t�$���Ւ�Ņ�_�Z%S���X�L�!`��<���1�h����7��H��#A��؄���A����A���a�_F3;,ﶞ����_j�d�y�Q�XlxVHYEB     400     110�IA����0����C�m����U4nu/��ض�r�WW%b����@�s蓦+�+�ݚ�.mk�#4|B�;�ˠA2XY�7����%����o��t��kt;П�~z>y���*_}9�4��2��d���p��3�V֮Ջ	�1"m#gȖ�:Ob�"�����-W�3=�5�A^���-�)�鵇��Ei�\1�  �	��-�M>���̭���3k�l[A��O�/��"ep�P�ٕzJ�	�MK�2���*��,�  ���XlxVHYEB     400     110��Y���}PV���ǚ�>�X�v��"Ѩ1u��G��nD\=�V�/6_LM,���#y�����ԷI�Щ��*��4�~7������Q�?�����B��UZ��ZO� �ʐ!�
�c�M�����Że��`Uƭ@O^��N$�f: g�|�9���ş-�:l$J�,�Ds��'�B��κu��p�>���c- U�\�t8�h2$H��9LmI�a���SRI�D���{!ܫN�6��>�~�#�b��Ӭ,������6����Q�<�4XlxVHYEB     400     100J��,'��K`��;�QN��Q�-بB�s��_��xp`�>���|�/ߊN�FU�!�f֜fG���
�Z��k�{�s�"��|��Dj�[�cQIt�݉�b���td�ߑ$n������q��<[kI3}��5dnl_P��oЁ�]��&F���ܲ7�UB��mդO�����o��k��i��_tD�Ma�$i6���j���i��@{#�L~iؿ���e:���%l���Y�?g�J)�8b�o��>������
XlxVHYEB     400      d0�O�u4�� "~��&�:u��BQ�Ļ��q3DE@�������S�:)��c�ùn�>hLͮ� �C�yG�����)���GA��
�AQ^�`K]K���Z�nп��m�~1Hb��q�,)�@�DNfB��;
�_�hČ���ڪ���ѺM����p4�e5�����x;X��x�H����p%S�U�p��lECMs��xXlxVHYEB     400      c0��P�c��1�
��s)�����"�C�W�R4��M�F|�T�h2r��$NŕP�u�*kX��0��/�$��Q��ԭ0Gn+Nh�ݍ(EU}��{�l���3�1/�5�u�	���y���>�����K�d=nC���%���s��{�B-��DiZ^���y<[LM�h�Z��.1�S�vd0:5�6XlxVHYEB     400     100`�ܣ�сۉ3cv�'�>�L:�h�^���+~��U��+w}� *�� �&K�������o�x�*dB�A���	���#�[Ǟ�r�`=�+�V���
d{-e��9@�o$}/�M%�=7h1@�����4gR���7�&�{�*�()&�W⬞Hhv;e�N�I�8ϧP>��&}h��s�.� ��<�RL��#2��%|�p��6��Z� �qrX�D�yP6����Z��w��|ou& ��뵦�XlxVHYEB     400     170���Q�r�}�x���!:�^�s���᷿H<%"BM#�_�l�C�ҡ��9���lp�x,fR�%��1����������;i�ѝ:��\a�p��p�Vm� 1ʇ��QWQXE�RHkn��d�8��o�[��}ո����:�5���6'�}�N���jH4S�`UXz�F����� �-E� b���HR����J��(h���ݿ�)�`RW`)�!eں�P}-	��s��zA��E>7I�-^:���]���'<Bu�� ��B���r���&xv�hӳ7I%�A����Q�������(I�=�a_Gf���<f��Tj����$�r���P�	��a���  yiiĢ�"�vuTGg��i��H�XlxVHYEB     400     140�X�F[7���Z'���:l�m0�ضv�)%d��Sc�3����c�� yX��N�n���ݜ�˅��E4�^׵r���4K�U���8��A�,�J�t0�4��������]^�r�Α4K��?ToI�
rL��bk��,O��Y���I�N�P2O�!i�z��Z
E�G��C����uq�C����br-�ΨUH(��[�1��C� ���p#�\�}�V���	/���H�ICq�㖩��B�N��tb���(����o���2�Q�풷%�:]�Iw�B�7^ϲ� <��B!���z�@Q�8�h�N���XlxVHYEB     400     100�W�9(�GkDe�g�,��Y%�������%`�}��;�H RH/'�e����7J*,a��XP�O���j�p�_���Of����Ƞ,zլ\�����Az� ���������h��"_�&c���^�����{;���m�Jڲ~Ҝ��Pee���3�e	E�-g�~~���Ts(�-�2�Tx?N�5�@�4,��k��僎���y̩���j�=�����(}tf_of���"�l+<uXlxVHYEB     400     130*l�CKF�3 ���O'>�N��O����G������G+�V!�Ć��/�ӗ�o�B�r��W0�l�<J�r����MR)���WK��dAOEq�0����'�?�%{�@ V��fk�bt�;�*B)Ϟ��i�3z�U!���!e��l�M�e_��\���$M��MUh�t1�s3���C��/�VJ��"�!w\�@�#4�Ba�m^�\h
vɴ����${�h|�E�\�[�sF����
Jo������#QZ˹N�N�{�o���)\5>W��^�<i�}L�f{IK������O��;XlxVHYEB     400     170al�7�$d�˟�%=mP&�\I?<R$爢%1CW��Eӏ�$��7�:��y�f��񏀩���#���0 ��7!�;F%�D��p�NC��n�Eɪ=��΅�rs9�����ڃ{d&:~Jr >��ҩ�Q�#<���7*݂qǎ�m'Y��s-U�a�������K��U�{7fЊ(���7�iH��i�k�����Vv,�=��:�!�gӹ��������Ufr%r��?��T����m��'Y#���i��{��h�ˎ�89��
�@��9��������S�,���G= f�*ߕ���K�ы�Q��g
��`�ئ�&��Q���o�5{�u����F`�����,P��#�	��y�����BXlxVHYEB     400     120�S(�6�>|Rk�[y�O��3�� ��AN�,p�4�O^*�-�ߴ&!��uy�l����#%��An4D�?�5	�eM����C%%$	�GlB�SN󀨍��D�c��_!���
�K�"�Ӵl�k(c��F_��b��t�.GZ���&i&vI���'�QT#�Xp�y3����Q��I��NB�䪠^�t���2JHfC��s�1A��^�*Q��DL��mO0��^��.I�t꺃DK��i�7��z@�O
�l���I?�"�+�X^h ʰb+�֑ƙ���T�OXlxVHYEB     400      c0Rt��_94l��i�ժ�fT~%�x��O�РV�t$t��u�)��Z0U������/m	��w�����D� {���y�
=n��0�SQX��O�9�ñ9��!�+���1L	vi|�TW"/]\�2�ס�c��H����P>T�
����#�S�t"�4���P�t*��������V��θZ=J�3,��XlxVHYEB     400     110�s��e��hP3]@g@�śڒ�($�,
��k9���iB}�����]�<!��; (�t���Y�S��:�w��F7ƺN��B̎���@<�+��aN ���!Dp���n�"�(��yHsӺ�_�q�e�fH��P ����`�}t�x�Q�S�YT��M9r� ����*���c���qm�l�R�����5ҽ|yz�hU��2�o��b�܌a�Lx"V������?ʰ���&��G5�z�,��������&�M� �XlxVHYEB     400     120 ���ǡ�޶�
�v������rp�ڢ�ȳSA_`�!�����/�J�"��b2���w\�ش}�S�-F�ؽp��Yءi.FEiԳvE��ߓ��y@<J��%�����	c�/\��A�y����5�!R=c���������V�k"��C� f\M�B���'��,����Y�#�$�ϭ�37�Xǧ��{Enos;�Y��� 4a��%��Ͷ�i�8�l����Z�WO.�8I�׺��2i���8� �b>�d�ᠾF.��$i*UY_b�� ��XlxVHYEB     400      c0辰BAQ�-��L�%I��.X���::K�7x�yJg?�,�5�����3�����Lc�0p�וlkhS,�=ʌ�[����B��C�@R\R~���X�0�Z������I9�����?��6�/�H$XیW?��
��V���#���m��H����c!? £8���W�T{E,=��=T"��<�$��lҪ�l XlxVHYEB     400     1208���\��w��d���n%dO����y5Hk���� �y���Y�����M��ox�&�E��;��1�f�trF��U�ڻ�]�腩'D����� �J 1����զ��d��q���bC�D�%u��O��p�e�/�H49Y�<ŵ�d�i��;�&A5^��3/��pⲰڙ?& (w�ꛒ0���Hs�_+{=l}'J�U>����0=�a^U�/���q��.+	��p�壺h~�9+ư�?�&�C2aTIx�K�h�A���(C3�#q���'+@xd�ۏ=�XlxVHYEB     400     110�u�9�Y�vYԈ��LR���
��������_Z�+G:o��'e!v���"wm
��_&i�(������RI�<���ΰ��Vf�y-�H!��I�FpM�<�����D��$��I�sխ[��\l��r#h�-p�Y����9��xhfts�)
y�3��L���S�X&��(��(mx��	>B��2Klp�R���{ܞ���sa�EzakY��H�������aw�'�"?�k�����^m�G���4`�U��sXlxVHYEB     400      90]J�<��>����d�#0�C-?�m�OeG8%���R����7x(W�t�/e��ރb(���кM�ĭV&���ܜ���ܷd��ɶ�t�h���Ў����A���O���l{�,�h�HE���ݲmL[�GC���=+r��e�XlxVHYEB     400      f0�~F��w�I�~DH��
��襪&�~��fy	L\�#^��t��¯돀�� ?	�I�9�Ӎm6��A��;�T���x}�Ґv��B#߳�D��`��������@���u���A��G�W��*ĉ��� J�	�-����W:S�B,m�y�P�����9M�9L�\%���ax�z�2-.��Z��|gZ������҈���Fk]��e,���^�$�<*�>_�y6:���_Wۢ&��m0M��XlxVHYEB     400     110h))��3�hId�f���#��ЖR��m5�[(�:�r���ŞqY���FH�d1���sN՚˻F"����Ϸ_�sc��Ĩ�"����Rw�8>ii}�}2Q�����W�	�B�:�4[Y+c�Ҡ�9��c��1i>��1gb](�� �q7Ð�]L�bTȣN]	���m�r[��C[pD�xsE�8��hׁ���(���{��$x�R�d<u�?ߟp����/[��l���/��b�B��bh�s)�į�h�ÄT�ݿT��I�N�JXlxVHYEB     400     110VD�5�W#�2yq:���_wnM
1BuVչsz[No;���Cmi�Qݬ��!r��.}}�¶���"�S!n���4�ΆX@��"d�`��~]}4���^�%>%䃕�R�;,G㒒�G����=�Q� G������6f���4A@�T�AJU�3/�TuϦ�͠�Ir��b���k�^^ w�ߺ �G�f�]A���$pY��,���[h�"�4 e��P�b��v(�%^�$�>�.�8����ˆv��J ,$�ߙ����p��'W�a�mq��XlxVHYEB     400      f0��m)yf50�p�oSLTdV���k��C�u!��ϛ�I�ǵ���)�IyZ�bЧ��� �,���>����F���o���s��X�f�x��Dd�K=�8�I��rD�[G�­?�Q'+7��M���1����1[��I5���G�G�PT�i�,w���Jo�1� Q;ݩ��Y���#�_a�f znrm4[t+�7�C �kxO����d�d���gA}���K&g�yiXlxVHYEB     400     130�-S82���/���rw�O��}\����,��՚�[(����%[� kn�����f	y�Q�Z�r§�����}-�ouV�*�݂�-:VC�U������N}��BTx���p�b�-�����L����)�
����Y4�	�,�݉�ݍӖ�KD:����"��� ��7���<�őΕ��:-�β��Q�����9e�^*��3�����/E��g1��1����No���ᾣ6���G_������\EJ�#V0����ͦZZ���eG�,�\�Sũ��XlxVHYEB     400     100�D�I�=���ݫ����U�NeV��d�ʉ��4�y>���TL�_R�Y��A��х��%�o۟S�{�A�1굌��|2A#/Ξ�\r�د�E��,z8wSs\,"g�Xx����T	�+�.{�e�Kg�g�_C��OԩރK��mW�U�n[�X-�x�NfE
�H��;�/F��|�Lɤ����ʰ.E�רX`�"w�
lT�|�=&�iw�e�k�AV��@���K1rdJ�l%�f���b���!`=r˸XlxVHYEB     400     120��z����t���q}�:E��=!�[�uhc}�¡�G��FƧ��ı.Qh꺚�Ξ��ҞϏ܎ߺf� ���W&���j�*<C4�Dt��v�+O�\���LW�V�ea��\�r��Kp��M0�6ˀ/�Ij�I2�8|���'�5f�,����kuw&\�%����po+���'�Ğ�u�)���L�p�$����<���YI�JZ�|�� �S�L@G�
��QX&��ۜ��ۨ��ά��H��X̓��A<�:�wU���8�P�gZ�Y6m	����;�XlxVHYEB     400     100���T�G!\"��=�W���=G�ga�+�x��G��re���/A3|���`��6�Q~���� �7MS3Ťt�u��k8}D�l��ri"O_e/��
��PQ�����gnP$��K�}��ֹ��?r���{I��"l�U${Qܝ���ؠ/w��sR�~��_h���S͹V�E@��t���6��E�(�[��w�[vQ9z,���;����܄}�|1��b`�;�}��rS-5��	1$ĀM~�XlxVHYEB     400     130�;[�L$��y�����ӿ���Y֞n��n�;[_fń��.|H�o;h�\!������<C_9k�Y\͋��?��j�H� 7L%�T�փ�D�e���ou�`)���*����N !>��&��k�A��DRfA�:���-P��S>�Lfot���^�0J���b@�Z=���+8ܯ�>fop!���ض���`XyJ����W�Ն$.��g7�˛��B-�~xc�(Yì�*�l��+>5�y�8���EZ,�j}�k)Q.� �9/����q!,��FxR���	��2�L����
N1�����/�$iXlxVHYEB     400      f0��r�
�Ė��77���"�P�NmA�}�B%��D��զ�&ub����=���nO�L�������1�|cA1a���s���%��wT���~\�X,�1��ξ�21Q/~�@U,&PP����沀"^�����Y/���p~g�P�7�w�.��pz�ǖb,�E͛��/Dg�4i���O&�ץ�%F�2D����2��A�4\���
������><�8��?W
�M��<���XlxVHYEB     400     190n+V3�4i������\�3��ٜ5�P|U�t��vW��&Or� ���:dz���3���Ű����4<l�~��������װy�K�HC�;�=�Ӻ4�7�!eR�(�zr�:G���N	�F��Bk��-��#���?|S�R��i��&S��M����G~���_�\�	�U��b���wਛ\p�jQ�`�=E<vS�������M!���p=��*=�i�C\��P�8����V�@Ʊ��l�Zd��T��/�u�Jf���uqP�:��Ę��� UR!!��,�F⯠J}i�C$�O� p=��\�1�����Ӛ�s�,2�l�[��W���}�E?���roܔQeeJ��֤����^bsq�����6e&� tX���6�L_('e��f�\H����d��XlxVHYEB     400     120�� �\�Ƕ�V�l��L��tD�34��:��<��E�@0�0�G�Ǣ��.�Frˎ��[�ql�Fx:
��X˘����N$* �����U��^^`\�����0�`��d�P���o$�j]�<"��2�D:Lv�h���$�_	� �{4� ٬�r�Y\ DMt��s��^(����J�}���˻La�L��HO��tb⛋(7�3G�[{�9�>i;vԜ%RȠUTF8���R���.�w���t���n�G�9%e�8я�(����3;�յ�=9��'r�XlxVHYEB     400      d0g���	Nw��]k��%y���|B�K=~P[�=��"5<�}A���\o�Ԇ(n����^͈�I����M��S���2S¸���z�5��`�e�NA�D����� ��j�GֽH/��!1��Iܰ�����E@O�G3w�À��9L��g�,���<����By �^��P�fH=}xj'��.Jxe�e���£���h� sE�XlxVHYEB     400      f0
�
/PP��r����W��8���0��ްX�ߧS� Ãl�ar�Ș;�s4�Sl�$oЏ�M�ɛ�#�b�yJ_N�+�5=^u�r{~���P��6��i��� ����-��91*q)_��;i{G�Z�a������iӎ��JC"a`xğ�zX��R�N#]�>�"�%B ��2���%p�)c�}��(�}��(-!�q�:p��d"���D����j��/P��$h�F���V�͝��XlxVHYEB     400     120A�l:�*�.t�L@i���M�ޅ�|B��VtJJ�O���$��
�H�bm,��܄����ȯ*�f�=\A8c��rx,4�'6&���sx'�X�Q���x�w�uW��P5E�^��n>2�`��=�ۨv����	@�ãE�7��Lb?�p�þu�#6~�'>:~-@��7�>�����_�v�>3`]�Z�:��y�r֑8:����M�n�ޕN�tE����ٛ0�����S���;C�$|�h�h<�Ri�?�N�ry^F�8;�' Ԋv�]95R���S��XlxVHYEB     400     160dy����HŁ��|�݉>�o2���S1�<�D��V�:G��˩-���jM���=�m�Z,j�U��%捛�0�ol����gNc���"�HBO�#�ǶQ�\�O5_c�R�4������A��I�0��{T7��	Sj׸2'�OTs�2����!*�PIɇ)�t�į��*�8�����O;��O�w����e�'�)oc�k�n��(��ݗ~�͋ʖ�'q���0�7��?h�"�a�:�B*�DAB��;Ogy��}��3~���Y���c\��_�>�!
�d1�R�F��IU�}���-�EUbz
����[�m��m��ѥ �|��ƭU���XlxVHYEB     400     160�ŤX�wcZ�����lS;�uZ����O�la+*�SpZ����XR��8�h����֖��%X�=��������@�|�q�z=P.P��Z
Y#�RD7��_��}j�V�g�m��U������T�7Yf�ݡ�zeT�jT�|^Q��[~�O�t��y]�:�H��改a��Y*ָx�X�� hr�k��A��vK\f����J\��g�������w�����/���]:$fYst���x���됚Z��SW39jUҏ �v:)��h��i�g�u��g�)Z�%�ȍ����m��׷G�x�ՌF7]����(���( ���&�=��u'�
��S���յ
�8{�i�ySXlxVHYEB     400     130�,x��bR��4�d����䀒��Q��&��b�⊌��P釕��=��jΫ�����u�`�Tn��#�� �0jވCw�7d����vB���4�\U��{���T��Ea�8�/�$)�+!�5�H���RƿxD�f[6�bU|ti�|�ϚE��}�j�iς�ц�ӻ{��o�V!iR9�Y���ݟR���h��#��FLJ
�2��5�C���I"�dKl~gp>x��~m��������s
��!�fx�	q^a����H�h��#�b��˹fi{�8���WH�n$
.~�U\L�>+o��}�1��SXlxVHYEB     400     180Ab2��<j�qT݀�q�mu�ֺ��OF�:��P������p~�N��=䤺qb��a4��Go�O���T\avI�d��KUȫS�M�"�WI��p�Z��KF�ĉ�`,�ɀ����Ҹ��o���as��s�1�t'	�9kl��ίBG
�QM�#�FM�����Ƈt`��C��YU���jL�G�'�Wr5���p������N|o�T�!�"M��_��͚+_$���Z�R�2��;yLG��v�?�����=9b:�ˉj�%z�4��JV�Nm��x2OM����h��9����_b�R�BYl#_��R^y2����!�o?l��P�Lk�,ð��RR���3]_��r2�&߮�JZ�K.��_.�H�n� K��XlxVHYEB     400     190	�<#k�;��}]�R�;���N�?3&���e�o���B�ƪ�vR��duz�Z��Dz��;��!���ǃ���D>���i:���^�}�YW1���:6�7c��Z@5�$Y.�݉���!M���+��f�s�fП��I�=���Ǟ�Y���i��싛E2�f���1�����k�XD�fG�R�&OBO��<p8`F�\�����74�$��4=o�����]J�o�N�����sŁp��4�>*U�!&7�Q�g/��E'Q���;�)ς�Y�#�ɸ��m�,��\WQ�{�f�������"z)-guٯu=���_�.��1�9l�T���
E�߽-�fa������=����2u����������s�MV7�}G����VP����zXlxVHYEB     400     130�޸�(�`^A s\��h4MPٸ�������@	 �v�1	�{�'hX�I֧0��OϑXF �B+|a��:�H1Ս���B��F�q\r{��Ij��Y���$��H�4�&�z>������h�bQ�(����\?bJċ��Z.g���ccs2�|QTK޸O�N��P$
0��)�biW>ic�ZC�wM���1�SUN2#�jZ�͛b��\��eR��;��.��8�|�q�?�hێ�[3Pw�ڃ���Pҋtʁz"��\�����:s��a��"8��w�;?��.t*�*�$s�XS�Q�XlxVHYEB     400     110\�/u�p�zN�ܕL��JP��=pz���@z-��Bu�vs�u�:���ϝ&s��#�u�}8s�=�};k�!&u���
��MֿWf�_������,��)��*�n��B?�f@}G�ڪ�9��1�2�M���Ө��Neߩ�*g�OqJ��<[���HT:��*~�6k�T`�ߍ�}��2�O��&Q��|��ʹ��Cxb���fI�'돣x�g ����f.�p�h:@��b�;^$+LŁ$x��k� �vf	�6�e����cl.)A='��XlxVHYEB     400     100!S�2�;��~�~� Y�H��d��&T���9� ��z�Q��R��A�6�Ub��I�1U|��zC���o����
��d~+R�%q�+�S������'ϵ*��fO�D�m%��p��4ƅκ��Pu?��`�!���M������ѓ��tw��q���R���8�|-��x�mk�;GM� !�,� �d�6�U�ژ�{���>q�T��­�t7�ĳ�����u�I@��{,���Y��u#9��ѼF�\qYc"D1NXlxVHYEB     400      d0������h�v.ш�s�Q�
}J��W��Q�-e9�ZP��5yU8�gd��aj�b^���#�3@����7���q,� �|{I����fT�0<�9#�>A��l�a��'�kz���:1� ��ɢn}��fd�Jn����1�:9c�WR���G������9���7;k�zF@�5�%!m�Bq���F}� ����X���1&�ľ
���d�XlxVHYEB     400     150]��jk�]�>�X�9e?����m�[	�D�5~�h����"1�y�M��Dņec]'f��������}'7l��sLu���OЊ��f+�pI���(�F��Գ��l#3v�4��7'�vq�C��b���	�~Y@��[T�\��E��oqO��7�����"�z>L��_�U��r�$>k?�4���ˠ�j�.���P���җr��+���w?��Ѻ���*���$��l@8��{C�=�l	fAM��>9�0�߬@��8�,C��)��uH�P�ޞ��3��נ�ȥ,�E�ɔ�A�.�@�����rm�5N}�Fɛ;~=��M�� �mXlxVHYEB     400     120�|sͺ�y�2��e4�Y4�ul!�6c�^���r�����ܨ����.=p��瀻�^Vԣ1�>�Ϙ�9�b���%����6�gQ�ed�4�Xk�����T�˴�yv���/��t:k�hr�n�����n��AZ��pP H룛U�#B��;��8C>�*�"����t�_&jpr��2���O����VCB��h�װ�#�O�0��Ϙ�S��:��)�Ǩ�R��]�8C\���;�|�MC�Xh������*�d���|�\�L��*g��T9oᶣ��,A?�6��XlxVHYEB     400     160�q�X⌸��3x�*�d� �ll,Ы	��,����7�R��g�����!��hB�GcL`ǎ����-�72��� 	��͏'���( z��-o;�ǅ�)�.���a��+ 7kw�H�+��z"��k�X2�/��*�3���X��h���|rb�#�{�>�&���ANI�i�jJ�=�w��������,���ё����>�w5RM����o���2q7-�D��!է���&+��w�9�RZJל������l��,R)��QD��Ԉ���l�������#>��,3�;BJ|�4�Zsʚ��2S��V�'9�j/�U�ȗ�OF|�v��1L9]$�xow^=�TB�/�6��)�XlxVHYEB     400     100���"�^�K�F4�|�c��F,m����q�`(�H��Y�����;-]o�|��m+���߿|t�	��� .p����ֵtB�$���gi9B�)��ډ���_8�l�:��L(_{��N���������ZV��S�(����ָqHR�@��]���(�f���j�U�5��9ګ��]�{s�s�}L�
>�d5$��'��J�oR�@���|��<Q�`)y�e�zNR�cN�P���R�6i[�e���XlxVHYEB     400     120P�Y�mV�#�W�+�$ynΎ��!��I�p����C}"@3A�����ov�L�9�v +���8�A��X�;Lx����[�tP���HI��sʬ��j@�9����2.�m���I���{w��p������g��Tk�98<
�!�-_�����N�@��\3"52����AЕ�Gӹ{[���48��d
pB�v ��T>�̵��D�5���1�a�ܐU������������R0�G��M����Ø�*ſ"�6K4wG������Ч��XlxVHYEB     400     120(~�c��P�>r;���~�=4��:����M,��E�� �)1�>����<�p��� �D/h��ۄ�����;+q�H�#dNQ}*{� 9��D��z�����3$]�i�u`=���^SxԙE��J?���e�,�s/}i*�H��V�e�v�X^�Fȕ_���<
�󨝵|�ί`�����l~��sx�(�T��H4j�c�ߌ��,��.)�ՂRF<�W�ݵf!I�5G)�����T����Bߡ��V�o�0!�a�}R#K��Ү�	����DJ����:X�O��Q$XlxVHYEB     400      f05���6V����v|��]h�I0�Z� 9M?�}Y�g�*Z�_�b&��lCcA����FzB�{f�2�|o�mw"�W$3�B	� ��~�!����ˎ�Ԛ�r0��ѐ�=�]�����3(PU���>F��{�^�������X�pcJ����T������BO"*���c�E+_��`��<���F���_X���z��7(�t��e6B���>{F4�=�NI��\s�W�o�}����DXlxVHYEB     400     160JY�l��A�̀�'D�^of��$0^�^M��6��S��Gp�}�8�q�޺xV�bm��t�C��U��bh��_�n����"�䀟KZ��� -Ľ���Q{�n��A BB�t�3���8���
���1�ͬӱ�'Rަ&���ܒ�#y�(�dQf��<�������;G����e6}�ձ��FG���;Gb�V��C�+v=��+л����+zs���.њajc~=�Z���p�;�H�����dW���_Q}��}�6QHf��^o~|��~��o������F�"E�:h����B��LIk@(�
G[YD�v�;��{�!��dP�)'9#��yW��-�sAXlxVHYEB     400      90�j'l`Ƞ�I�K<�����������/~5��tGfY�����ZI���F���Dac�w�dחYn5Ʒ���#;�R���)�-T.��˓lr(�;h�yȐ+=��ضA-^+$I��O
::���#I�j7l�,-���C&���XlxVHYEB     400     1407�<�����ʸ^��H�����0F������y�R|��� /[i=�A_��,��A]�j�������o(J_ĭG�I�4p��ب���ٶ�t<��+���w=�7iȣ�a����,~V�g�@c������ �����Uvg��v�-�����U��5�j@����`�������v�}6툩�,oa�(a�����}
�mv��-��$�����^�_&�|)��2M)��a`� �ȼ1`t�C��O0vUtӫV)b��b�Rhun#!�iچn�#Nɜŝ�2��@3���⬱eD� �]XlxVHYEB     400     100��8j�p^pzQ�c�{�d��f��gj	ɬ�3�_���-,!�LD�(}�sU��y_�X]W3��������g�L��#���0Gq§�Y�� �t��x�ڔ��W�˃����i~�J��XL���wX�k���Y��4	��U֢�l�<UcPd��Aj���a���я���Oj����Du���>��&�5E���ݺ�*�m���K���O-��v��.�5�W�aG<E��WW��+?w�lB�/���6XlxVHYEB     400     100z\0Y[�x� ȷc�,��/�V�%mL��u���z�+#Z���8�o��dI}?�z�ǎq��>Z���{zĂK�1�-FСX�Gj�ZPR�6!�֨�&�r�gn7�A�2��jN���'��l �-��ykj�6�J�����p���bK�X�uxy���Ė0�� �	��4��ӱi:-qc�_Xn�c���ՒKE��^R���Y�}��OL�Gs�(��R�3�J3d����9��Z�����m3XlxVHYEB     400     1100����Lz��O������O��� XJ�i �3N���ǆ��1���)`姞_�8��lj�����~R�8��_�f�eZX�o�&�e����p!��Pgq9ƈ��n�
W,����52�M��AXQo��\�s�+6\
�	S5W&�>�߱�B�3�R�^t�d�jʮ2k`�o�,x�*��~��够/�58m�5�L#0����%h�Eu�wu��5��Q�҇2ASSG��nl[����[�v�����>���O�NP���=&�XlxVHYEB     400     120��gAV@�L���PMx$|[	���0�Fw#і2uϚ�A2��󫢽�����`TחZ���v2 ���~70,��O7zޗ#��zvi�p�����~�����]�x`��}Z%]�X�p=[1u4���y7�Q�Ffon=�j�|�%�4,���6�c�]�~!�G���"JA��Nh���J�ԫ
Y��5�L8��� gD������$6�a9���o-�H@�m��	�.��y
"�L۠��w�P͡3���Sҍ����[�_��y�0�·�d�1�
@o�aY�R:2XlxVHYEB     400     110�ǁ@�̔�5�Ԛn{H�7���Z�����b���5����+⬝��#~f�]:TJ� N�ܠ��Yl$�P�퐀o{Yb9�(��]ǕN����o]�.����J���qo�;!���6=&-�C�Y��Ǚp1-e�58����
��\��uAHϣ�q���sZ���ǡ����!�g\n���I����r��]�D/)yHr$x�y}����1���>��ں �l��Er"�A�'���Z�h������:��(���k<���R� e��_��(XlxVHYEB     400      f0������ɖ�#��Đ��;���i-�����;�'�d��#Ξ#�-"n�����\�<Z���Ů~�r��=k>�P�]�@H ^�ئ�/��(%Xu���z��n�M7@V�WF�����ക����.���Mٜ۬wt.��G�����g��R=I�wήޖFtK���yKLQU*��O��s�z�*��xV��Ln%���D��i��or��IuI���SzA�~�T�9"XlxVHYEB     400     190y{���#g��\W�e�7�Y��
�A��Fd��5s�?6�������!
��>��P�ܪU������!���ު��VS��]�R1�Ȓ�ɂ�v�D�c0$�i8�ñg�D� ���#m���1��0#F��O0�Ą�	́+�:�_zR�*�l`������<j����+|t�jR��E-UE��R]3@�n
�רt=�p�sd�M�F�ى�!�d��3���Ů+`�A���w�c�ް�68��T���c��T�	�g�=*bWՇ�i#��<l�۲;�QH�����P ��zJ���kkL2d\���#�t~Z��f�r����c�N�h�n�PC�X �՞��՚��w�H;ך�#q}rM~�ᱧ�y�4��)�XlxVHYEB     400     190xU	��D�[�k
���T����M��\�4�����x�rx,��n�4|SA��*���a�JO�G��K�,�W�g#�AU]�Y�>�q����z_�L�\��ls�i�ߓLaW�������P<(���s������^&��q�yYJ��U�F%{�x�JLo����r��_��̂!����避��/���˜ȩ��_����e����3�5i��ܻ��� y*(, ��rp�����H�Ĝ�d|N�|�|�_���$�w��!�b�kP�dc�8r̉�ѿ2��6�����A��nB}e;�;�6��A�C��?ֶxy�2D��i�O2

��jsJ Ȫ�4���9 ���H��lw?@���ڒ���$����tFH����@si֢x2�J�a XlxVHYEB     400     100�l��[LI��SL�[.C]����^wȌ�~��A݈a��i������f"b� �+�9'}����*e)�Z�24S��:��Z+�<�1���8
jm:mC�x�W�ۧ�l��ŗ��uWS"��6�����u�A�«�gȩt�j�a��c�v�7�����Q�0�@S�O!�,*g�+W]�q纅���0z��x,G�����7�r_�B��Q���ї���Xq�?o6@UF���G�@�/��&���h������hXlxVHYEB     400     120ۢ'���@s@oNY���ʢ�dx	!X�x�L)����ِc{m�1��B�u2I�r]� �trYð��g��$jb��M�������T	<ְ�lYLHG�����6>�T$3���lF� vƚ׆q�z`5t9�d�Vi!�_*'�:ʬ�}ݫ�z�G�͌gS��XB��r����R*��Tl�`�e�[ >%� �t���A�����䍽�+���~ߖn=]��ݞ�����y��2���WKP�����g����'=`M�[�ʼ)l�ʗ���yc�2`XlxVHYEB     400     120�b!�y�p��p�çpt��yͣ����69�m��	��C~���̑Gg��[�g�o�n��xi�I��`j¦@뼞ѡ'��=7�g��(��4��m�U@�5�}TH�-��89I=͚)d�3V��]tT2�Iq���zz�Y��y2��M��ݎ4t&섈���!�ss}@��ؙ?I^Sf���bW�A���,����f���s�)��C'A�	�m�,����t�0�YN��z.,��V�sB�x%�4��y`��4zWM�f�#Xò�0�D��xx�z_�XlxVHYEB     400     1a0]�oF*9�Cs��x�z��5��%��Ϻ;�[�w�g�T��S=�����$�2�V"L�WcϺ�C=�s��M.M؏��KقC0�X�\�[��:���WD�Ɍ�a�D��CsN#BacL33k�L+��)�C�9R������<��۸�6J��s/��I@�I����Ծ�y%?2��ц*�2/�-�f�a���VD�$6�����I	MYS��w�j�!��@��H��q��iC/��OߺY7�����r�/���RT�΅�.ې���)��e����|�O�G?��A?��0���_��(�uRMg����W���Xx�za�살�Z���mFt����\Y����s'l��;���V�j�{}n݀*�	Q�1��������du�"A`)�XlxVHYEB     400     130�F�;%Űh ��A̠��r�p�df�s�e'���\0�$\�0b�,�-��!�b��2�>\��Ƌ��l\��麔@�@�ٚbYE])3�oDd=)���ʞ�Ԍi������"%�u|��i���oC��J�S���I��a���
��X�֟Ѱ��$���-����+�l��Qp]��^�4�מ����6oL.#�Gt�J���j���q��~1���)�]�ټ9�e�ω��	r�g\jNn�	�<�,��B�])���:S$��P� ������kţ9�&�4��FXlxVHYEB     400     1901(W�YG�N莳�g۫~��L���]D������ޅ�s��f�H��Q��$C�-	4���aZ�xS� +}����B��a�Ԣ�MUgR�>�ud�<�B7�ԅz�5���i���@��=��"w�o6��H,���Q�CedH+v�p�~|!PI�F�z�UL��/G��S�K�o� �6�q�BZf�������b�����D�VwT��NS�5�*lC3�v�����>,&ȿ�剙yhdT�j3����mLp
�؞�I�3��ZĮNw�IRI���{U��k��P�gu��>�-��3^�ӓbk>�0�q�C6gpO������
��ݞ�Li/��4D:��T݉lT�i1F�?�N5�D`��9J���g} v�T�ۦ3KXlxVHYEB     400     170Z����7��4���Be�;H����U���W���p�t�6�RէE�k����cL�Wv��(����b�S=�F�-�Id�x�g*Me���$��Gjc�J�������e��%�>��8D�A�+ϧj�pH�z�n�hE��Q���H��5Ob������Q`�$�7³�Rl�Ad|��)��Ny���@F�0z���˩���A9ZD�����Ԑ�b�ہ�Dg3���,X�m��
��=����a�z�"�.��f�g�}b���|��� �Q]�A� �AV����X攲ځf�upS�dVE���(=O �ZKԒɚ���� ��VKꤶ���a��tݏM���/��5&�����]_�, XlxVHYEB     400     100�6�`V�m�X��������Tܙk�Ĺ5;:���}�4�m�<��չd��+�VF��߳�\lҕe�ԟ#]�d��)���1��>���6�����P�kj���Y��ؾȼ��Sҏ���^�%��|z���r�Le�Ѱ�Q̪~ ��b=>��b,�E��y�����e��Xө������g�m��m+����V�\��ײQ�h�x��ꑾ�<�#�)c�c����e������\�C�XlxVHYEB     400      c0��l$W�+m�U ���%�� J��*�� � ����-$o��ʈ�,�b�V���[W��*����S%W�զ�+Kra �Gǌ��\�0�v�Y�3/� ��FmG��YD%}���4���²��b<����������ڦo$�b�yG�a^a~�B��OH��Z��ku���띓�g$%m<�XlxVHYEB     400     150��%q�xC���?�T
��H�����&��,]�s�I��+�mr�'Ϣa����,�������r9ge�V*��*�8���)���j��:ҠG�����8�c��X�*�qr^ςzܖ��:m�K�͎���,Y�w��R��4\�k�m�\�U������-�_͑�.hT�u��	r9
����i:w:��������W��ec��~�~��t� �|���2��64�,�sa%dEJ��}j���X��������}�J׷.X2�Y�P���v�V����2=��Au�*����g!��!��0��~�����HvvY���'�s&m����&[u-XlxVHYEB     400     160(,�Z}'J���P]�n���(b�N����Qem	bT����fQj���m
@M,��Jx�x�w���Z1��)��J8�8��'������f�{�s֯�:�������_�j���'�s��#���U�e�	��Q�5%��x�R�A�n!������0=��b�UU���ҎB��J�6C�q�� w-���O3���������Fu�o���r�Bō]iu�>��i�6'�=X�i��o2��u�������3P]!�k�KmA�@N]g!��UfSfK�V+))G�7��r��9�)R�����H�����'�6�2!���MGa�//�*r\�T��J\_�;��XlxVHYEB     400     130X)��k�hV��ם�����rҍ [l�G�ڠ�{���m�=%䰣�
ξ��l6��� ��6��Ύ�����c���%.{Q�W�`��҅ɭO	5}�^�㜐���P� ��|���<z���`���@�a�q�Ӈ@�b*x#б�e��F�X%An��������X��4H�������Ѯ���J�r��]���藸.��T:H(�pO��B����a� x7�.3�կ��O��|���/���]/&��{{�M�F���G�����"PJ�>��������!������I���-�E�Q��m,�XlxVHYEB     400     110g��S���!�Q��V\<B��n�UL(�K�L�	�:�I�876��A����Փ�H�!jF?ޗ���U9�`�)���MP tXh�E�	��>��h�r�*�#V��m(��"�PQ���a�u��xD]��My������?��c@�ǋ��9[�6�y�ܼ�OE�6�8ɢ�5k�����P}x�:�ՎdG���4�> �Ѭ�	Ɗ�[�w#F ��?��L��;DPə?�4D��B���ָ8�z&N��Z�R�
Cf�����tXlxVHYEB     400     120`gY+�n[�UͲ=! �?��C!�)'x�E�/p3��mc�J7��1��"g/�����C�!�)VǑS��a($�;��.(��~��ƶ�7���!�ze�RJhU~�6
��沞�R�k�QH��I&�M/����Z�P�b�"�()��h~ٵ�!4�WM���J��1�>/h�l|%���(���DnM�j�Yj��s��叄�&�kJ�c�H�e�:}-޳X6M�����Rk4^�=�*���SP��m�I3��>P[�vR�Y�j��;)�Bd]��m��a���XlxVHYEB     400      e0�A�OS�>o��m����=�ʲ-���r��<G��$^0݉���.͕,�D�	l���/9�  �W���Q�J-R(乩�Cw]W�TG�^�XA��%	}��ކ��nDa<�y"�ƴ������]VՖ�L��<�.�d���(�g��Jo~���ت���zk�tv��,#�fl8VKJkG6p�}"N����|�y�(�IBe���$�\;21E�o�'!�XlxVHYEB     400     120������B0E]�.ֳN���Tnõ8?\��T+6���gU5�	����fG�ix��=����:����8��x���E'm���j��;kgg����㉘��w�Za�eD�k�6��w:{�v�������T����"��;K��$�����gHoҥ��T&�>oih�!�֋C{�N۸�}l�A+ p�29�ρ����Gaw��]z��B`������Ǌk��A=3�]��{6*,�:���u�K���!�2��UN�!Y��u	ػ�֥!A�"��"ihat�ި�XlxVHYEB     400     120���힢|��뵶��aLT�	��.��%����v}�a( �O�5݃.�W���#;��0tR���!�ȝἳN����=������.4#f������p�J.��A��;�WpY�U����MR�|pa�x��ԏ^���Yّ~3C��=��CU�R^+���Ύ��Lv�ʽ�ߐ/����!3��N%�3�s��~��ߏ��|��wjl462�,S���BOЈ#�p)��e�9�l:��p����W�7����.��ưj�J.�Z �`6��h��,Y 	�i���AZemXlxVHYEB     400     110����۟��W�ʦ�WO5�e�eR�k�;~���������_�h���B	{U���g%��$��ǦQI�P���t��u�*���I����.��uXJA�GQ�q`�U�w�+���#�q�pLÕP���̯�Dk`D*���ؿ�)WM�`SY��G�f=���s(-��{*�6?>���'GJ��M8AZ �LG)Q�J���<���we;�����V�K4�8�+="�r|���ThkA}8��J�Z 6 I]� i���ϡ�V�#��XlxVHYEB     400     150i��|I>b�UE�}��5�y l��{�_�)Aj@�����%_����k:Xp��2Ԭx�"�8��̹�������LI���9"�n���d�x�ډ��L�e�dP9�N#�H
>t�W-��Ae��x�8��x�ӈL��NW�-���R��˵>̎��܌魓
<�͖����AZ�vi�*�ԡ!Hњ���:���Ú�[4蕯Q��?��6Ԯx�A��{�O�X3Q:��C�i%@c:a�e\�0><� T��	��ǜ�142��\К���L��$��*R�|��$����5�8%�B^��?ۋ��){���25�Y�.��ro�߅XlxVHYEB     400     180�S������a7ċ����O�a 0���A�y ����5<�� ��?h-:(����oj�i?-׆
*�U##&Ʈ#h�8q��p`�� �Ԯ���ʅ����;�ʥ��-������J��:̭BC+��U��h��/��\A�,g���FF;6K�Bv>&���B���+�-���n�Q�dp��fO�}q���і��2�^6"�p���r��l�=��Z�f
6�?)Փ�^�@y�����/'��d.��i1'�5����Įe��bZa�f����1�rw�E"�$�@� �#s�E����L�%����m��x�t��}׷ո�(~U/����H��T�J��pq���}_}��pф�Mb�/�!��f���Xә��xXlxVHYEB     400      f0[#��k}���i��*�A�cK��?��9�wg)a�reWP�-z�0�P��/2j�X+���\^����r���b�]�Ǻ�|.}�[�^�3��I�ٴ�.+��r�n�y#��p� 	ە7�ke�(K~߃��?D��`�'%���&w,.����>[�'Ϝ�'߿'.��A|��X��br,��aە�V�3�?����5B,z��f-�԰V���v#�����+<@�y�l�u|m-�]g��XlxVHYEB      eb      80lM�'�([IGCiA,a��M Ù�w1��>u�WY��=�
��=H7jt	n�ə�+!��70��ؤ�?��|�?�U�P������*l��`���L��O�Z^���';{�49���� ���