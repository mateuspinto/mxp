`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3088)
`protect data_block
DVMmkTuMD+LGXg+HN1m9p/1r/lBn3hF2eJt/dlay2pMh1SUjkqRiVdZLme7EVTaIjgiW5GMBXIDp
9tsu2bT1tvFUlf8spyJRZkFjz48PhH0KjaoQeOavTZ6nxz25CZCJQzu0e9iJRoW7Jqm4OqVcSBp3
v05+eiZGw/dzskdOHUMPN3V2FG5Lg4allJvlVe7bjEulQ8wHaovKByLWpiP+ho4652n3hou2G0EQ
P3IM/aSInjlNEwyMsEVna6WvF0IY4Vy9C7XeZeRyabDctyzbHVhRuVZFZzM4PQTt7bv9ScYTJRSR
PTERSD/8luZy8Iuy7X4irrMvPflb10lYw3zUPmHkP+0TGLjhscO+Gnuz0CSKZo2UJ7Yb201RkO8L
+/EWx89ZuGZOMgEoMWO2cUw/G6BWI83iMM5ZWMDwMIjAP+Zfzb5Jw60eV4pUCjqr9/Q2zsPPr44b
mSWzzu7/wkrMwr4ldXupiSLMkThGLXdGUy0nx7OcM4ZPENVxFXThkdB1RgLKBHra2/VQvTpRdw6F
yi3K/MBq9Dw61g/R61XByjtDcHqRvGLC38tKs3LvmZMTw1Xjc2fTXyQ298K5wK4TxDWHP2CcdKsZ
wEC+7GS08lgg6urEVv+51+1nxOg6M0x7KGHkiTa9taHc/Exh0VE53hxyD9++HPSC45t4TBMwBqs9
5KOMHrpf1p96Z5kSObbFYczHbEp4c75+6xUkBf+eZnh2X7zslvEe8zhB56K5ntxKebMf7mRsVCW5
vs99bbA0dJQEP6YkLjIrXcSjIaQyUAtw2+P33rdQmbmuYFLU8EpT7CoINwluK8fxeXWjlubLZUnI
PVckFw53QsJjKmrHfxLzJaqPRlQ2ELQJllXPGA0Tf4bYwt9OyQplFTsCzsg33Z6X1IWjH/ba7B1Z
ioPVV+x2wiFvEZPfOSHt3s24BHFp3o8syIUZlaklbC3G+RoVMRIbpz7d96Zt6Qungjulr8jNVuik
T8jMZeJGVgWgEp5JnK9wiYMZZAMvS6bWPjkidmmNfnYplMZci9UHsSUFTGSbzsr3pXyGarZMWtAs
6YVEarCx1Tv7Dy1O4v8iA1lHZj7eslI1iq/Lw2ExB8ELBz3IjJUmTfapMLif+LgJPkXGdG80PFrs
18LfuNR05oYO2JBwNk5NayNd3cisyrcYKmKtWTUdnzF9XDZyUq5ogOy8npIMi6m0r2puLnU6wdH4
T35uuyGOjvEPAZWLwgdtK3PLQ3NHkBk7GbTO/zeAK2Kti3RTQn+SyeqPj4y0WAk9XJFv/Y4b67YI
aLuQuBQp7PGLANMVqQgEWNGnGNfJ8RTFLH11RzopiA5Y16UQn4Q5107KFlx5SB0B+89E+CPVE8XW
8ZhiycacBcmANzyJkktyFmPm3kiiiN303fHNBJoo2xj9Ab9dkZjWc7Zusi9CyAy+a4xEwi3ddKTc
FvjepOzmbOD8bkJNnGIhUit0pXEeWvh13oLyZBgFFFK32s5LVALuycbPfrVsIDMpZvNqDoERA29L
1cjymP5jl8QHSG5JOnmL1PC8+p3hKjtBnTbrQO/9rsywBuH1Bd9YyWKBMQG1vjWMtOsAphYOXjTt
Hq9EXNRhcL3s2Ol2q+PRdJh28IZ3M+o++dzHA1317adB+SXg5R/6hq/n5FEjN5NnyHRYMx1K/8lP
bZTQk9yTsEif4Q4SOVuRJvMbrgf320eoHYRfiCpVRDeUxW8I6Cg05k8olQsFClcoOr8HlLZvFkHG
+CiWnN7HPMgI+0aOjI4ZO9M6AjlTyPKVoHtH58NGE0jJ/9Wf7Xrr/c1RPT3i9ZF3uTb2e/g9vKTY
SDNQp5GKigrRBSJr9BNOPelBlMjAECcfHuc6r+Xxhf9GbLif0sAo8Ks8Kjgm+MHMgv3Ae5t59Aua
bU4C1DthPg8mrgcfH14NqBB7qxYtp9c7UX94Wnv8l1DprL6ko8rrbJ9t8eauC0Sz1mUHHrD1F3Cx
TLhvnaCfjhsCqv5zGA9vY2SlAMXDnKJyQZs/FszwDeRLZzMweiCGZX7K9JessHnnuOA+efSTIrIN
ifH3lFZ5RaYvt+zOyjJ3JytTcUbCPaS931c54ZSjpAmaiSOvDM+tCRh4opl+Vz8+toIhvcSIu+/f
6s7/alzhkVnYpv2sDas0OBy6pn3t0MJMAQNKOeJdAeprd5/BWDFfWwXSod3qJvJ3E0TnrLJlgeh8
MpDOfjjrBZA2yj1YeI2+yyHmbZN461WhSE4VgQVWh4cpGgkkkBtPav3rXemLPYalnP+RILlq89E6
od7ABqMGIJjrzYrRd1fAqywCZn/dZ7O2Dc6PQN/YZQ7JaYPapSZdG1BxilfBLb6xy6JDdMf8pKbN
7o2JnRHK8uGiMbfOkqssSPZ8BB9yZ6bk+mioaSHynHZmmpfQCh0cO9/eEaSvrfouuyhUsSpBeV+4
GNWD5L02QO9TkdYlg6xm6HZXv95wdHnjrXP04ATHssfYELH2CM34/igoOEw+wm0Ks9VHLFcDeuhJ
t3YXAm1EAkDlbXIkzP39cnUEy7m9qqgZl4CzS/gn3fH1f+3XE6/qNs3ewyp2N9LaXoBxmR5BMCuC
3sc73GzZh6LbgRXpJ0zAUGCMVaBGgFI/XafUQ2FeWhXXLijQqzasri/qAPEhEaTunwiINKvI1Drx
0JghNzg3zwfptiHpBpStPbPY2Fv23TSAiSTJxePlgIvi3H/mSLkgm736Ij0b4WY7BW1Dp5i5CmoS
nqWiOlyHeWgy4fjIUZw42JYRmyHeq1mnH3rvBsgvTQ3A3uzf/rffiQSM/JISLdELKf/mNxo9pgm8
dLFhMnAQ4k86OG1qiUoPfory2ZnW6xGFr3yrkj8jbDyC6x4uq/DUxjxa16feX9nUB+uBiIGz1uKE
QzsiOCKxw6JeLgUznWG0wzFr7YwInZJK1UbKvvuoep8vs9RIkjB83ON4ukajrlR9pxEg3pIqz9xp
uuuDQrykeASr6qhp15TlwH5PWOTB9aEvHZ5RwSNHdHEl2A4TSFnNUGYKgUVer1TE0gc0N0fVwP9J
bdekjL8USTAAS6LCZ0S/A+4cfLntsbSoGjinuyv94pDCXTvf5YS1N6FA2GAbEmk3ZEzAFQkKTQ2e
73vn0co4ZLsjpdX39x8lAIp+01kh0ch1G7BsBKA2OiDW9+/yB9aGkp4IOEuzjuk1RvH3HI3Fjonp
Z/1AafsJ2TpjYIr5+alRKpDw/t/PLHuyfSqhABo4l3ZwSGRWYydLscRgNpphqs1h3/FBgxgpysGa
ZyYu3xM3lC1zqSAFWozSh2tOscJaWxduU0PlMFS0t/M3TVNeDzDlPCg9kLC+8PKWndkss8j/CYpz
rCVQgSLgESaqcR9HlObqK696L6vEpSOCTfdmWxL0UJ5Gh0+/grzeXmHrDp9voKluEphEY5XOwVYy
wkbR/rfZLF8oe3FUe44WEWiCaCfZVdLrcRrKqj1+kE9lHytL3JE+tbT7KKR6jiJQsI/tJpfWFc44
o6nZUiWH6ArEIGhQ4dErU0jT4nbCtO1ib7YdYtnbybz4Bgwrk8urzmNq7jJsl3GCh//7C8ka7xXZ
8lGwn5BilG8P9L/b/r/V0IAvFDuIoXnt+Lkzz8FeMEl1LAO/QfoGLfo5rbFMthrqyT5GL0ZgtBM0
gp6BH6Im7Cy2XA9fsF/hwi7PII5Uw/d0AL5kT67WyrV01ld+MW3xtdTYb1kbu7CoikHgCaW3/NfF
nwIV635T5RMlpkARxnZzEUbD+Vj8DHIsz5yqwHdsVGWzQueN1Geb7xMlfaPGEPKedJJxrvNKDsf3
jfGh5gCCr1avhRGKiz7fMe+Nw1hTXs3MhAVxM2/GcqSso2vM0UUqDHebYxpiph/1cRmChmamDc2g
swBGeyOIHqGYi3boZEiwK8+11DS0bna7/fsMsXFMGV+oVk8DX5em7fhRhm2j5wpYc2BPMbzBe1zD
OCGGNYwWWlfeSLlcBck+v/P7clUVirhLfpDpu1fw6ErV+FwjwftdOrl6ecPYNsLRQJzu3AN0EUsw
JkRG6n1UWQkSH/tqoXPMrfLK+MaySX4cETNr3SlxfZ6C5cDXH9PdWNsHKA6apHoRNMctMYoxcdLT
yfixSZbvLJyU3A==
`protect end_protected
