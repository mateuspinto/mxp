XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���0(����OmD<uQ�qq\+Ty�q?�!S�L�F2RȽ�ǘ]�&�p,�e��i��f3��쉬T�Eyu9V���@;=}���d����FС��
��[I"m����@;�~�bcn1�`ק�3�&᾵�V�������>��WT5��3�d�!�l���[�䑼�n�x�q�KQ����X3��O<v��{�����1���p�f�R���z4�'�Xҋ�Tl�W3��t�G�;c���[ݭ�_����ʩeY���8��i�� $v]��P�I`(w+-G|��ҧ#������*N'4�/t9=I�׀R;�)V{���L �fh�����H�P���k�l1�m?�����(%![�fT�g��~Kic��m�0�ȝA2�9_��[@1�>sK��F%/-��۪���B�`K�!���>�t��;#.����tA�0�Y�q��aE��̇��oM,�-�}�GۛV	�_��|\ٻ��(��Đ�P�a�"���7M��������!�e���/����OG��˒��&Z��h�ʗH�;c4*v�O����8C���Jy*%�ԝ�+Ij�Y�f{��J�>�?���x��8
�9�MF�|<F2ioQ�*�:�pN.����	��Q�}���EV̔��փ�\��V,d/��/�m*�@�u� ��ٔ��>�w���̶ҋ�y*B'�%���:��K*i�"��\�[>h&EF#u�m,�����#6�šc@�U��|��B໥i(m\�PQ�~->XlxVHYEB     400     1b0z2+��	}��oȍ	ik�� ��N'�=z�ګ�M��Я���A�-�Xh�0j(���	̌�e@���b1x#Fj]�#j�E֟�FNO��x�^-N�0x�@�g�1�8���AH��Ԛ���Ya6x��5�ϯxy�\JoPG���\J/Z	�0D�v��rz�k돛��t>�� K'��|�Tp�3A�0=M�2M��U�-�
VE��<���|�i�ac�u�9:q��ѳ�Z�N+7�75\�e�;�Ů<hϳ�R.�(��:�_�&�$yF�k����Xn<9��9��N����)�L�
"C~�LEe��nj�)2$-�R�0�ꌶ0q�x��a����rO#qfq�\sئ�l�ߙ���8PbX|��m�g*}N�s��-x��
��(�9�;7!ܳ��{�5�0�O��v���IPj1"�`lo�XlxVHYEB     400     130��mtzI�%�bF'd�:1���2��'��tS{�������mǨ��]
@��G���nf0؇�fq�]��g�x�!�9b�����<��Z|��P-�x��i�v]��9%�X���>���|[9x����W�5{*���}k���2d�	~�^�Pf�9-,[�l �����H"^ƛ���EӺKj�/`g�_8���`�kYTL)#[|�y�ofO�մ���",$rr�)����,uDi��`1BrW9��C֒P�w�n���e�?q��(�;���v}�4��<�!a����gp�X>kgXlxVHYEB     400     120k@Ed� �~�w�]���Rpȶ�?T�u��;��"����_��6�g�V��SW\��ҫ�<��4�sbG^���z�׀mG�G�(Fw���6}u�}���[�3�0���)ykc�o��s�����DH��yɮ��X��{��$c��o*��(i���3Q�4���"ԩ�����SPwe��w��v,�y<��,өkoL��cV�z���N��&�	���9���.Kٝ���O����Ӡ,5)z���3�GhO��Z�I��p�ށ��L����ws�A,���p�XlxVHYEB     400     1708d?�3`>W���kS럴�S�TC@Ɠ�g����xK%ZaI��ѝ1̧DI�/�8P��'�>�������(�9�Dz.a�rق�V)R<ʸ����Zn�*�'�" �/���͗b��=c��f��D���L��{���0f��H�D�A!� :��ᖤ)���%����A�hq���\�N����n����Wk�	�m�V����-c��,SP��ƛ.4'.�t����'���ٲA� :����0���oUB< �ʌ`eZ�~ )]����G���k�x>= .!�>��dE]���Jk�����M|��A�C\��u���cHE����ʝ	�1������u��J�A��5<&���XlxVHYEB     400     1c0B�|q��S��iI��Ȏ�����9c�8*��)���=��g����~��ƍi!e|`�N<��8^Ks�X|`)I9Ѫ��kc�QdG�!a��"h�m�T�F[������Wf�$�`f{	#XH��vTos�|{���P�
�LKH�`��=|����b�<�e�����������v�`��k���Hy�T�p\͐��g��C���7u� PƦ
���%)�����y���C{��/ D�{ed-E���>~b4��HfP]8�P�����\u��G�e�n����?t��;^��}�r�i�i*4^m�3Ƙ ��30���n��X��FC\f��\S
 ���cpP�<S!�p��ڝ�,��Y��H9S��o*P���JP��&�E�6jP�����w�?�g�zU\���������e4aJ\��vs�Ob>�\��^NML=��(}?�U(;�~XlxVHYEB     400     170�7l�ˮ;��Bh�S���KsM���ZhjWz����.��q���	��U����Q��	����Q�lsq��4P.?��O���Y�a3���T�M�
���=Ҽ�y�|U|�&xI̤(�"s���ՇA�2_H���m��\Ṱ��衆���Z����G5�q���:&����jǣ�_H����2jA�kz"q���僄!	��b�bwY��\��� W�d�A�dZ>΀�G��e���J���.�$�IU+�/�ys���:y_�!� զ;<�>ދ�h#I�����1����s�r�n�����YG)�l�l�����R��������ݔ ��>�C�~( ��N�XlxVHYEB      5a      50^8��4 ��C&#Ն�N�A����O'���x�!��ݻ+jvM�n�1�n�Va��R!���>���Ъϝ�a��2,���f