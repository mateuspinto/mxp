XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����-��egj��y6ֆ�ې{H��D�=Q�Q��ϻb1az#.|V�Q�[�]��<5�@����XL�G���m"1��\�:�
0�ϑwi�g�����!��'�,<���|nn� <Ãe�ҿZ=|ֳw_պ�(	�}�x��CU#?�)Z�2�@i���B�'�
�X���o��y�&s���h���J�w^>�Y�B������שׁ�dyv���"���$�u~����:������{f���mל����7�dv�^WǨ^�@d�\�F����%C5Ez~6���iI͘��$��"#�]�q����>�;����L"�c���z7sH���F�sI�� ����ת֜iKii�����Y��,�r��VI��)��{P���4|�CWp�/\�� ��
+�x�A��x�]�A�Ǥ�j:��d�h��ǯZŢ=��}���е��p��1ͬ�����H�͸��1=Y�����F]��� \t0�:������^Ĥس�ᕒܬS駲s��\"=ck���\!%���W��پZ��M��mo����y�Sxy#�C_�[�ۧ.it�"kz�������ޱCw����s1x�}$4"��B[�g��ݤ
j����Jy
�q�2aC��qs���C����T��/����O)�����'z;dx�`��d�/������ꮪ>S��^��Zye.@����S�N���gg�WH�j�	�ϲ�����$�b����7�a���]l�%lXlxVHYEB     400     190��w���@Oyc��v�����
��Ql��(3k�����Y���4&k���0�F�<D��1��-O���~��xKA�-'=#%����SP����:��Z��6a��b(�;*E�p�G���ք'������.�E�U�u��A�䞿;@>��Őc�Q����:�@@Z� IK�"8�u�5*�Dn<��BU����A�þ�z" ��2U���6��'heoM �#,ܻ�D ~BHMZ	^�3�Ǳj��)p��r8��ېN(Y�}n��,��03�N�MW8�?��ʓ��@h�(�Z�]�?q��%z�@�83'� �..�F��_�2�`!�2,��՞��.i�"��~�\(V�be�\"� lǂ�LΦƭ�o�La�]+Ƌ�W��JӾVXlxVHYEB     400     1f0��:�q�unf��@�s]7�k̇�rHS�i@ɇ3�����l��?�"�
B�B��fk;�;�D��z�ܹV���	H���Z	EN�3�b�EUc�^h.�?/)���TJ�;����F�Յ!�)븦���.�vp�CX/�gb+�=�mu[dblh��`�}��:-��(�7j����O:>h�q�ޠx��V��>��2�q7��� �´��X�
�ˏfϧ��z	���c�PPA�uO8���]j�ƶr|�
	�B�5���p�Sh�-ȎxA{��p�Zf,�0�}���N�ŗ���kfWɣǋ�0��ckO))s�������Xx6�c&�����ʦ�@Z�%w��EO�� ��Ij4�X���.���K:jߴ,D�o�~�=T�S<E�:�X]ܕ �u���b��Dm-�̢��f\��-�.C@)ϯ4�%��p�{ʢr���A|ᖹ�gԜ���d�d|� ��m"RH,^yt$!�XlxVHYEB     400     200���h�ôh�#�J���m_??A��;0#���O�$R��Cn�\x��N]kŋ���_+#����@~[_��
af�<�!v�)�;o��޶�/G�� ��Jûj5D�����@0n|���;A��G-*?6�tB-�#��U���b(�;��g�� e��yܽ�}�2@�f�5��㎼ee`�Ix������-���,ܽ�/�(?<�AIfG�#�ـ��A/�ao W�,^q�Zħ���Q3��5Ú��X�nk�yI�<@ȷ1����z�.�*�����iT}�7���T��I��ww�w���2��h��)[�U��s6�������M�/L�/l*3�uP��)n�;)�-]��\�O&��ant�7�#m?M�}�v�fV��O0Ϭ�eE�%�QS	_d(p��w��=�Ү�ځ���0�Q%MA���3u��w!|�`�߷�/��b8�<�w�����坙|�x����A7L����UYS��q���0�P�cCn��XlxVHYEB     197      f0�!�y�f����?���bBn
3T5ſ3%3��gͶ�l\Q&:�i~7�v>����c�_���%riD��eB/t63r�>5����#7�4x�6=�} �\`�	tY�`�[1��7ZѢW�P�1&!�����d�-F�]4�M8ûSԤ�^~�d�dE�pD���:&����N.��y�nˏS�4L���ѽ_)j�&7 U��l��T�8=I�T�$�OZ��@��_X�`���<t�