`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17984)
`protect data_block
ZM4KErOaarPgXeBHapbR4+T4IrHl7KSChmqX5Mbs/FfyLCEvTYZX62rCpAjdIW0CSd6BbdUlW0jC
RM1OXnxXXZsO/8nPDF6tdUx1bciDdd+9IW0ImKL1fXJ1teGJh9LqxUURkhIwpUradHCWIo5/zeYA
CGhKxgX/ZSocUhESRNCfeXlyoRw5rAR+IYVskA0NhpItQQVHnxBmhrTxeHacaOlxvzwZeaHxbAH/
36+KIqA77fgf92lP6y9bR++dpqiyAEbA2CtMQ4djygPETPPK8Fv/NA+LPHlzEB+V0NMIQnEF9uoO
J2609qLNN+TdYX+WNwC+8A50VxtdUciwLdjOeDSbNnBqViaVIYeFubuzYjq3AZwBAH6AaB4a21tb
OplQGdvfAbZnsOGVcvfQB9Uf9G4CblwUKyGm7GKckt13UZsQaTrjPj45N7TCP2h0BgRp08HT5OB6
HWzYEOw7IKNNw0XDpT4sTlBm3aB5vx1z2lEIPoiCzbowbrIAiwyNr6tafSfclMZDyjq9izvm1MFG
vuPCzC37ifXPGnP+EiCwpW3KkwCPCP0tMF5qPYnzIisF3CzyZxW3s/qwNjwDqc8csQWcKcHY3mhD
fGF5rJCgfEIYcpf8MLXv/ckrOpPtM+edsUxemOEUe/PjaSzEw51w3buqYcVKWA7toVftBSdJtO+I
93mLKhSss8TbPeFnv4q8x481kiRs02K3WKFV2BsteUKgzEnUxxLsVIm3baOKiXNgH+9hI7tiOj0b
RxOfBht0KezJTb4iocAWv+FdhcqtutZpghL4UXoQV8f6Fcf9BcbpvlGVfEMgkEK4qQvwXsrrv6hU
lbaG4vQvlkdkenudQyORb04Fn5HPsC0N/hKh1648WfOUreLIsWXAOinqm9aULzl4DtSScUUEduHr
nGiUXdXYd8QaFPjW6mOTJ6cq/BW2ky9GwBFfp/bmnXvnFWD4WePdGEzbnykJu49gjL086fC9uxS+
3grdx4fliG+ru9JpNZ1AGzVrrQ+l8RcTzHehihBuCn8uwGbjEKBDQ6AWe1ofAshv25fpmHM7Xk+/
ctBOKDJAt1Crz5T835HPAt9bP1ZixrD8MPS9MRo3Y6sxuhkn+WCtMqh2f/UBc+v3Gkd3jZVIL3RO
QjgFP5bzVeDrxTPM75TFedTHMOFJNM5HGj22ENEQwq5PNZ/F0jqmLEE5M6FSlj0XNVPJpfbiLB6C
GGxTIAU/TEFx7DdpsIynrpUcM+nk52Q8Bd1CrHIqFp4Z0UgsWhx4DjBIpZg05xbq6TspJmtZdolV
M1GqqpU6+tP0nFSe3v0uINNzUy0T1LOwFquwlQxsrhfTGJvioGM5JfiM2HEx9Xvjsf64igVpacOT
HCaQ6OZTZR1LYtgAU4yteO9nqVkaQzn7TONsam4H8lyAWIm/SkLSBAbfuqgtQQLQXQ49BzUiTEJP
NPp8kJVkvqiGqsfz6nKKBDgISQRfzGMyPFeeUU4MQVvjA0M+IDN+LJFo6hGbn6ZSxF0a5XV43Tdl
AQo8FAXMXCudS8fFeVzO0xIIYHVgGMXfMGg1bQKAh6G3iXLKBzrdK8NP9jfji7agmvyGZ8MaTXmp
/yR3o+V5Dcs8+Cl1g2XHh7pvRtcnE2WJEP4kzrsiRQvzXAtdIGMYyVL6/ms4mkJmzcgLhg79rzxN
BtOMnVOV/woKGn5umw7j0Baq4UcnphWVQf+ExIPpuyMtesWV4RoSiVQgoparcOPTCRTiPPZpiWuK
KwPGWLZ+FSzquyRqG9vYb17TuIQHKioWOjY/qjTA4wk1bpj44U7+yZ8iuIlVBy/lanktHI2Fp8To
I8Ekrb56/FuKj3MaWsgKz09qV15lQaJeludJK9HK955I4UkvaZ4kMwIr14MAU3F4LiJM/m/J0Tuu
BxpJXxMhf5cLtz1YBeusE1gr6PDwmFoWjbA+RtFYIQrtrXmS6c5r0obL+9snlMDw77e0T4Scbf37
BolDTbq4a2SggaIRgw9KsLnAn3I+yM6ODSl/784Zc7C8WF2FTIkAGpyr+X3xfZhwpHbZVVOF1KVA
BbMPWm/YLYKrn6BrNQnGOHZFA4xu+g996WLQBHE0aPKYpclFuQuXnMH9h83rjSoh8th/W0x4XRek
/UL253eUvp+5JFBJINmqjSQ6+OVjdEQIslEk9+92sxaLjnJ/jPfspVOR8wwlCjb6krqmARPgmOhN
+ffd1jXYXMGh9Io/A8EKCTc6o1FJXs/6PNWPB2CV+W6IXU/eEkdoVRR7Wm8e3CmzYAv4L7nELzAO
c+k94BILdujS5W9Zlr04x+7x+VK03wvNLM8VHRsrQR6cWvWEMSoUGZr8aN0wz3e1zSjsuzwmmwlH
c34ugoLqWU8FRU0GtfRHrerm9yG9yQ/BsEMGJItLQY7/DDNV247vxeb3IIU2tp3mmhWG7F/Adzgv
EIrBgNB79JbPCp/9II4ad4nSfOMQrYNeMRcjPASHr5/BhNQJlNXpxZJE3WNG7VsmKLQWEKS5XdQT
17iqV0ta5PAU3AsMy1Axqn9rjjTPppGPbl+G/2N67IzFx7Si5erCmTJQPLH1iJ8H7VNF99vPAYx+
dvz20f2jU+xjHZeDJs/mTxNKsFAfHfduzB/sjiM08RNlSQPom8b7//jDttKpX4sZmi09TWJtTT3w
95F9oYabsGp/6mQ2K/O9+SlpEk3zG0nt6GKgrJ7T23VWtv2TUh4/FUerxvxHG5lDvw65Glbyfczq
w5cwXdOdMdraAQs+JCjYRsvDUlJPihSeQaby3yGT73CQwPsT3LCCbNJhzIIwss5b9Q7/PUjbKX3j
ICHd2vG2vCs1i7YICGicnlMPzvGq8y0YQLm1HTMvXkoUwKKV8ke1F4FrmL0uwUT9e4WamiI8OZY/
m+n5h3ldVYm93jdYhYVVx94SiOFvrx0pACSi3OfRcpJEdT1tvNa0OMctDFb+hlebJvefaFZjOH6/
vT9f6y1uKUbH0bim+XlLL07N2DgAPpBFiC3gtsbD0naSISoKye6A0FsbnGWPo2U5DTfxwqBGHe8i
aBBDHbDpZ5zdY0o+g0Hvp77bpYCDG4rNfUJqbuYG4n24X9zC5feM8yhMAzc28gojLNwsfx3WuRZ1
w65Jwix7Rgqt1kM7Dbg3SPNxGWZgT1kYJQTcUt6++vBKhzG47YaQHt3E7S9p9PebWFzwK0ol7k8W
8FIeX6HRORhvsJdPgQEykFOiGV+EGs/myfXoXroDCqdXQxW/7Dygo2D5A9vRO00aMqFa4AyEvBSH
FwXyTU7FlvYLLa20I3WHQdpeRPwsPX0X8ZvgzIQucqOHoJbKqwwB5Pnpxw3jrx8hTprNM/hFOGKJ
kVsMVakXcXO+ChZ79xXLEeAzM7yfQ6kmKP7RJHe+HKl32n/ycz3GwSZg7gOLUkcl9cF+4hl6fMt2
Mo5Hc4WBfD/DBsj/xfq0LXNup7BxzgZ4vjwrQZphwy1nVUp6G4lx/AHpY34PL3ERSf1K/41/EHJd
KlXa2NZZbbVOlBMSUTfWYDJnbgZU04jvyPgeK+YvV5JntimRLRiudtB5zMBXynstINi5h3WLlkMt
QWYJe6itOKTfbOoBlCDaeiRRFjqhhaBeob2qG3L+7zA1/BNPL4knhw0J83H5bQ+yZ5KMLQIiBoWy
5+Ucgc4z8lQWxWXWknAckGdb+T7ovQq1tPodYFhFlB7Y+XJeck7Kmn3Knb0Hmt6strHEL9JLEvh8
GBiuiii4yPo74jxF8nx97Mu9lAeXTJgYedvyTBmQV5Z+rbk3qKLcKUnRv02FMRi+HVvh9QcrZVDJ
BI8dXbDDHV3M7LYm0ss6QA9W1G8ptnkNDtPyADqeVzkiNKKHsj6hG0EC+TlrYB4lSbAYXdFc0mah
gJJLS0J77Y/QnYPFbuPk9DNuoiZmMSYHwH7E+kauvO9G40MCpe1Alp3SWb1SNrJsa+TFlXausYKb
xamdmGLhTrsJIL5ABHI58+5lRD4vQWXT4PISXxpm+cb7eEuVp/U9QwkP/0UjWkHoAO3Qjt2RX/nQ
+EmAqyMrYvlQco1K66A0MWBbDFb69JfLIYJ0DCXpzaHAmzWkS+Tl/CW10gsrgMfpB2bb/+109SSx
WRdpqxz4de4/iW2UnwssQVevG5uuwQLya0Zw5VEV9ZQXV6P1MzvOlh2Idldh9PRNgPmfwgZCqgjq
ANdGAKhfgeJaYSHhrx4WoFHzCvA8ufmizy8KHZfz28ENvK8GoHN1m32eLbMROj09Y98uRSDD4NzT
pBkILPVWHbnCYV+acT6kuBumu9nsYA7xmCYP+2wZ0zh6lOrQZhvKmE+By9ftyBXBCTbRiyYvYr/Y
ax9MswroOMVx80g51Kca1wB2+mbZkMlAbaRMWujQtW18Oy5E5/1T141pC323SwXSwYYyUtGkVMHL
P4tQAuJ2gYsCsw7Bs6HdNwqeqgr4NzAY1vKjR93e+AWM08/CXY4+KlO+a/ZSyRgL3d48Entl/RgA
/O4BS9i6PiC5TrVSa+utWZMkIS3VnBylQIhz9lPBT0tbhLbdsc9qxMTMjo323b3JIBCtB/wXEals
MiX8fT281mBNqvZOFPw9WIDmAXtAFyPI/27fQnLZtZ5Nc5hrXUAa1XxjVBe68atBX6YxRoHmQ3YM
2vb9/3pC4fioIZQ2qvbmeDyNsqhwMLLHB84J1rroqFUevgcrWjrxKXwSXKKA5LOoX4WT3yWYsj5+
xo3PAldExW/qHpvblmN+Bqzoz5zF8+wR14qY+KIobGRs2m6WUids1YMG8Cegp0KXwhYJKgP31IAF
Eb0ViGnS+SywwDNhGhiPcEYSms7OzbPEmaoHXfWBLX78oAGLQ3+yJTfVin6PuqKMH++T1H/ngQ1G
s7FdL2J0+eRz2JJXfRpuk1L+xp9IQT+pyzfnFcUqgpxKkRz4cOWFoGtEfPA2277UB7NZe03zgim+
SU17H57Ys/MU6bIhj3BmhcvvRUkQsDSZl+A/C9FUevMZKMAgc18avADUmb2xpKfxo/6QpvMukXjB
v1U03vgTjLcYgUX3WrQ6bY5XIgv9XfKHKvpEKBxCQqZJXJHJpgx7YZeWdqJLpbFMiF0UDtT3HM82
zMZQOwk1otqU8sfsVn2/7nuw8XvNBdOEn7rbxOMScAvFmOOAHh6O86WGm3oESWnvpCiw/mBzdF0k
yN3ucQdeMeDTuyAjG1HzOSnblKNv9d8wsOSZBEqV1YCO16R4bGh+3itrLpsx3cCRBQqRB89OERrR
FTRi+3SoYn9fofYk9ga5Jf7QEwTXAjAMTwhDLDcmBRyefiv/iZJOgW00aido86GZmJOSbHdVSDbM
8wgseAOck8rv7rEo0t0o0CCmV8361+AHquLcei4UIqdiN8XsBQkS82zwZ6Wvpjk+4F7EMOEKp8no
C7R81cieKMXUdCq+9y/2RpnyeFRSb47CrC/OzkCd/d5qGZABFULK7364NytOQReF0UejCn2ziSAZ
EFTth26c3dkwdkRytWDOYNop0aY/gN1X8/NWzu9NJsfqlKdsTfSFQzlSPLnhtpjmKisHkN6XkXu8
qgmQwz4UrcvkXysppk0qzrlRkdhlp4FuPBfJvG4YGDDY/1hYn73pIlm0NMA+qdkmza4k0XYj9Q2q
RV5uJaRGQH+eIob6SjLq5E79Yc1bE2psYjvc81EXtkzFRhSF3oQlZ69o2c1WdspXqTFeYgY+icrW
r8ywdeIklM3uk3f/A3V61Q8CX7kMwiWkcPZvok9mfmoJBdIx8+j4b98g3OwwbEhF8ggK2gEoIS+E
0Q8yx+73dfrukjwARDo7qwoWMOfYltGyqhcxuW3P1RITaTy5Fm1EG0coVlRl6BiSutpLjy5am2ia
D/52Y2XW7HhKRytjNJf/zoXPUFLgKiyoRHWmJgWz0C9fNg8RFHvNYnXLjKCAVtMP3lvoAkUsps8a
2UWoaoE9SGWWAX7yAsV0nh9NBsq2vUX4emo3z+cq7VP8eR35mGG3THkXom25hZfNNAh8kX3VaGEE
QSf45S0hPBokGrVbxaG16wpbQobSVf7GHXikCimCHPnhmqkvnAbBzfOOIFEHgDp+Wps5BsGEeO+i
KoErpJQB6jqpXsXOtACEd4LoX8GjGNeVZMpdGnBkR3Eqt5umiiOOcGdwWSR8BNG+VIhaFdeAj6Dl
+CxJWoKEsfATay7bJrxyLDKWhDfy4c7a9WCWJ4w33U3wLTM4a8OcgZDfWVseGrDsOpKJOmm/MyPG
qwnPcSoybv0bf9y7qF2QJi35ew0UgloPWHMGZNjOGzBezb3PHdH6nM3DxfTl7ZRMWmD6aEiQPU38
RW1PIS9eUoLwh7z7BwSEtlgwiSKrMj2IO7uk1/x5+var0LuxJF3u4hGA9MGGGJ2321jjpi5XFtUO
5LbTddEUllgu74G0X9hSDFjE4ax/GF4x8UvDnRhD8F1y2djMgRU/ltTAEKRnsDtr+qv/jhAO/yZq
62U8Pf02aYPJR+77oYhWoHN4A+biw/zCpSfBnoMBsAdEoyCWUEXk/hlasSPaolSiau/LmTIe/5ZD
zd6CFCEN7iaRhAW0WSGHINa2nBsagJ93X8jJkPhuagUensOTHVsgDXTJrw2lSxgnww9ve8HqdQij
RKyQnqCTd19cYtr3VQ8b2gV+jG/Wm1PYtBvaWSt+afLyxTUm9AMW/ngMSfFFUdvX3OP7RSzzaWfw
4b6PyOIzoR3NXzygm1XPriwO5LiGZoAs08AdOI6FD5YO/3awZ/5JZ2FkY7WRjz/5pHrrTKUzz2uZ
Px96VhKsSxiEWAXj+SqJHDW2T6/IMgKsOkuQPHNyl9aIaDjUrsXr5HXw3minloKJjoAF51lpf/CN
kYTZlQ+mdUj8DieDGRghV6iczIjNA+VJ7kEBDtewOt3f4rt/dPnknEpv9hnN3xXNUHJDRzgk3DMV
xELnAXZjZYWemKNJ+Yw5ClfRXflZPQldDUyio07b3qaUTsUKJHBnY5DkBoSDaHKX+YrPyEeTBkdH
YUJGnA4Dpq890PkI6c76DbTo2fAz2qF88ExzgNsck6BNhnc+cXTNgWlWSdiDbsjRzcXG8zaqh9a0
B/KhrN2XRF4D2QqA7nlbMyEhvQ/mJlVh/oBkicpJGlsQu9l5eaEq/jLURZqGb3w7JXIRmIu0jMZ1
DVrROzxWF5LZWyaMYyefctACvh2X2/aBh/WG1dSzvEOS16HGgdMTWTQqLMQHXzW8liL+dcn3KmZ7
74062pS41tcaXdbyg6p8MsPseOKq47c7kuDPD1PT7eK9X1hs4ouCGRdk+YS2itiT6JZCJBExVvHL
hJRLvyI1hFzrh6ZqwD9rJAyjeON/xcu51RQZzJbjSQUaPzK6gKjqXjkUwxbWeNIlritdSQ15Dc5d
feTJYrDxD3YNSrTASYxbl0cBJGaN69Pr7KHMFQcoOczBxfRSDCSLXeSIKgXn730HceUca4Gfalhu
EfzioBfBC7J/rYl9UykPKpENSufh/yqc4rHa5eeTfJ5zJdV9ZdHzvDwTMP6eOeSxqCdWsmgloA/x
j2lbQyAgBEIsGVNqUCcf2KAbGKOT5unc1hUdK1zLyHdoTM1PVeGW/IMbV7p0SoeyuqrCrX5MKyNN
dJm0rn10Yu3w2kYmFdS5brkFfxRpfK2R3Jrfr2xYVdKEe4mq8r2Ecbz9h0Nyd1/l8iTNcM1rQ0qU
HBOCNKTeSUvmtYKo3mN7P4WTJapN+sboO02hOXeZmUzD17DRqYwpKvO02x1WGFhz1aMIgXID96ci
HfAJmnJ7cZy3KfhgNWIDv5jSeXjQiDIDOjsrwmhc6QSFGvoT+gg50mY2SMZ+DomQzmn+7j2QLPWm
K2NUMLLNIaAz9EH/0Jo/6YD4JVLLdP2BGQ6baAz8f4WvyP8hY0gctmCE8fGGx5Z5EixM0/rsSuWn
iIyWlvjbwULVjmAVr1slsbaP4ZhjXVVG8haabzGE5UAMJGPzyUDmR8cLBnrWNvCkQky4aOIt0WY6
CpDjTywCAhmRJYwi+FqX96zCHxCFZIS1MtamB0ZFuAgEYxyQ2tGvyK/DQVyH44llhc+5zMvRAADp
tK+8K1zmIqZ42Wy4uPAQ5b6IdWEPYbdoEVPYx4zbqgwQ3P5g+ZJCYEq/nAra3Hv6LTdYBssokxIy
J3Cv7TtxsP3PBZqLfu00QiGAdO5ua75dWR1q920EWpTaEbExX+RSGWwKJ5Qio6qYQkabUrCCI0J5
59HMLLfeqpDJhzAbwjpLkbOu8Qro3X2zH3KQQYceYLhNF95bHWdlsLvao8+omfLBlMZXY4DJx617
lCjocrxlLoWqavFGcwf17yM8CjhAzaNgu7nNMeIGP1nzpQbtp2pYyg/b7r+/KkDMJ8tIf1kXLs6g
Sfv08ZJbtlvIYxiwE0fspjVuoN6CpDGDWgI+XvRxYwWlQOD6/djc2QIdEGqbdmZNEChuByvWmjgi
9tBRBrx0et3qUKksRe017/ykpHIp7gk+RKLyRoHSz3Mh2NJr4SC9ls3cso8pGj+zPVMXkOLg0qW+
LrjJ/zDqwLipDHtspnH1XdYQD7RpXsL+5eH6BbaW8Mp7/crHkl1pOP1U/ewjbSUcWLlrRjs+kEQH
g4lTNNmul9KM3TYdYLWNZx0T6qdRUIPPCnVUoLJGNZ3rjPMlL2R4lMfJBzp4sK4/vNuOeohQdEDO
cwGwu14RhQVtso5oeKbbnoeUO9fB+S70kEkQ4VG9Njz25bnopVzls3s3mmTU2TpY6pM2DvKzO9r0
ymQqotZJrRC8m90LfQ1ca547mACGfZTpE1Lcs2D+i97T6xa5uk5BMS5duAfl8Wzpd4jf4LLEd0oZ
lQoAje34RbmwpvFigw2G7qESIgoFPQFDiP/1wZJHr82GqSwwe90eYQfJkp5XzlLvIEvsWWte7+n2
kG84/W5i5gAk7lK8SCaY0k6UV0KpoRdlyWU6iRXGyXMJze9IlOMb7X5IRYCDBuKPrDWstXtkZbNp
5YSqDYZd4kMHlo9wJcEF3dLTE8dBR9q+nl0BkDqjo4VHIN5rVx/GBD96JvcUJzWF0d9idjgNUNsO
dOt0Mu/YKk/jYJ0R1jV+RakAAhjXHarFx1XLe6/wPqTC55PLaJeJMMzl702D2pRVh9ppGsVjgONu
oW3qaVHPg4DnCIL1dxvn4XzDa+mB3WbcKQRrX2Hdn+iZY2iL0E496BkBVkSV2w3H1sp0RzzhlOi8
O2+mQVjf5t7OxxVwzUi6ZWwygsMeCLGgi3KVLMsNFc6wWOA+uHl2LeQwhfhwrgFtZkzoWLGKfCl6
hmQkhJjE7Ws2rJi7A8mR2ELQO2ifrkphEZbSj5Tz1XlYZGgW0KeWl0KQmKCqwaTxKkB9NLRIhf7j
f1OpAa/uuKluawXnfXaHMIEwV7v6GS4mwxOeSJTYed8Hn+JoqfpZE25/KOHwA87fwriIcw8OyH4Z
PPBlOtTQSvGmeB856AKzpO63Hdu3XnglvMWPabO4JtXiRo8U1nQEYeLpj8SPnQE8w4VHs2IFZpxe
3qhMLahkRnWCWDpxYG2jgMEFdUVQam8AdHL8YdfUrUzdHe5pChLui6kfEoC3lLNnUy3LisEeJ2tv
m/yGlb699Mn6WUdlQBFxV9xhkEu0f9wj1F6/crKpWK0fgntw40Wq73eOSsay2+LXdHsPSWxQV+Gw
APcv92QexAvWvWrFBaEqbGLoTTMlxWYSexRgZDqu/F8kEm6oidLDe43Bkv5dmoJZxlWuCOQLh+Et
oc5foOBQB3LonylfPvqqaTrcrnBgA5XFvGFYBsuG5tYXOa3YqXQIr2WvoSJYNWdeDMU0SV0yuw7T
yxf2q7vnjqT9OAKSzKaNJp+JpdPM6SpsP+MeQeM2Ar6jrj+41Y1LP3dcs7PDm9LWMv8Lg/aKJC4x
kAp0vVYFOiCZeR98m/mpxrm82HLzkh1BtHkrRuYCWKGwEBdXKYsIzGOM7Ic/a2KkFEVBBjfa7+ZI
bzeeE3q6Vq8XkPj6B7uNpTUHL4RjlOsnXa/GMA2Y8fDiU7Mw1WZJnvt5msiVhzEGeh4tgjRzTbaY
kzWNUzJHQXWuGfE2I63fiV7iTFEfnlnBvEKjrp9/5l99d2QbLv7PmiKN9eanAUW8NLXkhNOrSSfN
gPKzYtqMavS6eaS37uwl+5bRnYdfqYrZbEviiEalKIU302u01PUgRKMQQ4RSzpwSwX13QKlK4D3N
kkfiGn+ajoy2FcgSsQTmEvq+1BPbrBmdMAy2OzHD6bbG2kyGr45bFCoKwg1wbHdfFaOlRmlyp9ZV
kJ/u6/SxzD7IskgT14aloY3twJzzYS9+2x873OHuQf0ZSVgoQaAEbxt6ziS4xfqPz5Fhki6hSeOM
n+JL6dOalxFwcvTAW9C7ycKldRZfnumRSopzjSVhb7a8LRexQUejZgd0JJLdNeLEXYwG2Dos8UsF
Rcy2iEzwwEKNTSnMZ45yutL49NZOIGfbvsLAtL53OyEeJrdyfakN+gKKKThWIVCisIOdwz9EKLtv
3TbHoABzfYGUDOj93VlvKgN0XKn8fATwfq5S8MFfStot1AAHWgkZhBcKYSHy0hihsEK0HiFNNO4D
o6ISTG6gtmmhE2eRE4oYwUvDr32c5taIRo/J9YDcJcy8VwNx/XfbFkavuo/MmT5sqcXBc2ZB+pDE
MMH5V8bICN7OziJWGeLIMA0PkTLgTvngL48raxvh1k0cvNuU09Yc9r11AvXzJzdynfhnNNOqmunH
+6ophpblvMK7Bmuf6BP7k5Erg4vUWXfHzA24n5x3wQj6qBZ4+hHUAXCo97hu8p6qrcVmNFDy3ZWs
pFg5Evrp84qnVHhP2j9w5Ol8leHJToik9a+G5HaFLdw6MqDjPa8yAwSP8siDekCPeeLxPwpzrBgG
v2bk8x/B6sWfqDUGOCYEwg6osmv7UJMjQ8aOeHRU+wS7ipTglScz+Kmj1QSVA0+CUNGrpYBfiJUH
EW7WIkLT+BZgTjfW6kkQtsSuH9FQOOTy/Pg8kDUNLJofPbnZT0qNSMk9aOZ4WEW1pMdsPdBmEM5f
V/rVQ4tP406toG2nD1EQ/0AucPMpkTXrRT4QDGrCz14Ep1S2oh1qzwEyQFoD3HNv2YANVg9n+bJ/
C7Flwe66W9K829nuKPANgIAgr42Zgoo/lwWHfyu6xfFfooNUMC4/hVi9sVx4JkrXU3vNWJBE5mmN
GCCIvqEpT0zb0zVIyXQ4HGeTCNh6ujQMgHS9G4EiC04K+E5aOW1ewKNf5NsuKcotGM8DOxrjArKq
LqIOZtk2RBhzz+zf3AKa48CYQWMiQh9klUIM/GRcYwWl2v6zzaUqxyfNwOhdUdHnHSy2s1SO6boV
LN0VYOPqQaXSNEsftdOuiZBQoqLL/x/cmpJPdpFuR2ARGmxo6vwmjNIcBqdeZyZOA8tIPs+iwxII
lfLsfmQKW3MmkpoPEordYRXdXigjsLoWd/1zznCeOnc/ddt7SysHDy1qNTkgL4kWAgNb4ophQ494
r8JtxwU6vvCTqXBVp7A+BhM89HHHwSvdIFRbdUXt8oigepL8dkwDUYXln5RAmwPx89XTWswmyTuE
d3NRS7reVimxZf0ZN9P99FrAb6c+fWe/CJ1I3foMQe5aWsJdZ5Y6MpwfemRcvPTxz+aivtYpKYvt
cWVD89+6jTX9yfo+cgO6gA7cTcmwuhax4QC8yiTzCMuXgDbPmze1z3tvXbrpG+6qJYuRNqlqj8oM
rqRuOlKy3wf3CskVSWGU4Y+CuM8N2ht+nC33EBvj67sD8IfcjUoBRYkJFYreSTPGGkISaiyYdOLR
n1XaxCMPLh+UDRmMlM2lG0InrJpxvG4BQGaY+ldb+ZhkoE+oBaY4BecqxRedy0+mnlSl3KzwO5yH
XvQG+mXnHd71RIfwFnObiTQGC3WP9Ys3+503ig+WVO2q2NnGt2EFin8jSZ0msqqfSknTDG32XoSU
5e2b68Cc9yc3pWeN0mYFp8JEO9eFz1N5GFeBNAoyDL3/nY80RrOzhuYHRMVp1U9GMpcb1LsKRIfE
aObR8icK2NInNKHJiXqT8dG6S4WlbNoQ6UBMgqFOJfn9Ic3TJs/FwXkQe6SqSi9Iz6ylDZNTzEuS
tbF+FH25Mtrjqwq4EYqOEfiVMQIDhpJlUEYK06mVgRbXcVzCSka1hoKpcVst9cMMtWgoLkTA1Kk+
jnRu0eXFZkJ5Mr7/TfGIzM00R1JNLKToMw6CxjULpSLnrItDUzM7BidE1hTdrz0IrqjlFpr5s86b
uaKEjVpoGDEfvIzcYxT8Hf/MvdJNtvDieSD3YFR2uVQCEti1ZgBSsHQ35Q9SHPUUvO4RxgeiYxxG
+VqlYqqJ+t8zTqlOlKkcAw7j6RrF0b9HOkLrVkQnXYSW0U06NbmK9Z0R4PsuCWaN+l7uDfsmomBa
e1UmJ9cZJtqY7YKFHOJ73ROomDfQhbwXDrT7mo/NIzZZ7etfpKkwsxpNoCshsZtZowIU2DRNRGR+
tQ6t4rqrUa5cm60ILY8hiBnma7OhYtyF2zSzXp20Hie51KVNBaI5/RFZe1xCcWBRGji29N1CK4eJ
0kfu3997C1Mcs2cINrOxKWvGP6Vqbd5sdJPgYlJR+C/+CjtDDeV3xnRhuNQbZFXme+0IiJ3orlL1
8UMCnRPrF9ziTdg0kCKEQvId0W2Po2wFCde0p1TqX8GHIohrWuoaZ7urIKTdcuLHPbbVRwrVz/WO
U+ykQYmQg3OLZWPP7CGujV67vvNkdzoga7q7rfPO6JbSgXjx6jVzCdZB/Bc6DNVRxkjXWbfnBmpo
CZEPpLtLSHPSMQw8d0MrxJOl7bs7U2g59WPDQo0YCVkNyCHUG6j5A1sYtHvITQGu36uXJdgbq7e5
Rnfqke6UsDXHOw4NoCI1ianiV1BN45HyRF57NFl331i/NaW2UlgEJEVq/JqNMDqnsiM/cht2f7cX
Ky9MKun8Y/d7UIDmkk/53WdhyZMr8I/j63QPLnCVrnMWq8BpHLzAIj8WDxkSBlCP4lQLtRMhLmbN
LMv7M5dH/Rq4L36WaJ7twB095KDVrlMZVATj+uFmtcM0Yr0aFi6b4U4JweJEbPdpBEnR/WBZdG04
FmIHGjuLWPJJKMkgXifDMBcaijlTQUXu4sROeGIZ0n7p+Uv8/qZzVTZzYWetXdsd73Nzi+gj3oR9
YZCsqusUl29mBGTjqV+c4cF2ryJ7tVqRYfP68l+qrqBkqPCqnQvvpSGYR1n9Li7uTystat3TSaNY
NHEk9kZJ733NmpBjw85Dr1Gbm3KMlMlDVLfzDCWP0BKdt81M2Wd+/7ebsHSdgkxtOrxT+4e3CiVU
8ZAI1ePWSwAE0Jwd8pDaF05lJQ01Rf7E3XdftnwjUd1US2w1jfmfFYks9yx+hFPBySEwnITLj6aE
qKNzw4aLsB3vlBGvalBfIeRToSBccJzeVG04/XPBTL0wFdzvJxNAANoubmWFxSy/drVlXoGvJSJm
vMdGBNIwuYgdgeiQCv2TR6VRO+OPRpX0y41OV1U9PtffHbp1tsN4kmBh9TXc165em9mJIBjpjXzP
BpeKCUCTIsl6x4sRLa3BBDmARcSdVPyxns6Z3Utr3hcYjtf3nninE7QIqKK+iJDeKYSJKdI76MIs
3OLRyLxVJp8m6/7riPpEkFALDlSX7QDlLyK9nKWF1ZM3kwAb3qk2Y54v9zMN2DPL9ip7QpPn1yg1
L5hpUKdU2JgLvP0NYpgv8XuRURm2ifY1qNOT1LhihI3SH3vAYegiOyJt9cEbd5+wC/6yu+3Rw9Rh
yMF0GpLeOny1j+drVEV/Ap5eM8jgXPuoxVaqkCRGuL9KEEkRaPn4F+CyrncPA2SE7Tn/cLybL2Zr
TkbqlQNb1Yf34anVgjl5IsIchcCSuegh9LP8+gB1Hwn/cwoZt4m8S0f8Hs1K36+6rxTq2k2WTkwU
xdVJ/HZ94Foyu2F4jUjSzxN8rij40VMLOcwCQ7qTv/uwrylj5ubRhPtnBuxSzDn483i+XP66l0w8
4yr9T4DgVfPkK46nVsGWBKzGcuOvBQKW548+ODANF4wXLOUAM5ioew8cr9pQp8NlEbfMsesSwG2W
FzlYZINyJEPa56Pt2e91/wFOYG9JdNipzpDj9Pf/VdDMYq/ukeKwbZD7SmJQeC9mf/+H37vBFoqx
MfwWGIESMFyNMNrKN6NCEpu2lkMaJDMTFLkfywczjQNAFxFtcNarKQmWuGmBw9/Lf2uZb2fRLZny
5R04YKqW5FbNkD5QxRyvbBZIpTbA3PW30qmAgae5Sy3nBggW/e9U24i3SA3PfVKpbvmy2HlS6Q4n
hvz2+5NXbFAHe4iQ7ttGSAcAZo1/nR4kirmKebZQwwqXzF+Xzs8YUPPeLm6TE0Lh1NS807EN56Cc
VmeWd7vuBoIWknahbcbCjn1k6fRJqU3fn4kE/q5r7zabCwsIyKJ5ss9sxW7yScVVmZlssI1ycI6g
+aKDW6PD1K6aBuxIeNy09SAthHJARoOBFSF81mzfaKlgx7Ca/xC4Ay+xtJ3pm5RvfZzSdEOqR0aK
MBGRixLobbqp+0SBXhPjnH5N4ssh4ieHfukTt5cJII8OHtNYJkOnGesGJmheNAJfhwEP5z7USc8Y
j5PIG8GLtonT0+H5RXcndbHD7JK3N17zLldN4QeRI9XXfBrSqm8YzIf7L/bq+5Jl1jys/bz7VZi5
2t/LeBM8QnxQAuHpYrbqooFSW5TwOMDqtiZmbeRVOiUfy50n+8dVQczVLdrLILJV/Zw+f+8gwPIP
2MkX9L/CLwfue1z8tZBDI7ozq/e5f+OV0Cv9n4VP6WuX+RM8dYTXeHxMKRxcE4OMU1igDyMfJKkN
8c2WWJHnMQ5dBbNBcNSnAWnP29AK3Qc87gKgyp8UFPTna3a7OUwr/4m6Ro1zouKLR1ixuLiuoULd
JcAzxbNIWgXjLmFgaBmPICxLnwqD76ZXMgPZbNTRAWfHLjR08OUkE+9URg7J44yC5P+W2X5hOrrm
nhLSd8QqRO80DziVOvWwmV/b5SdiHZGmuNx7CoJK04xVyIbzs34GIMDXQjMx2+l5Hp42qJq8AYV7
eeL+X2HI50fxFeuIrgO2F9Xi7/6FrXyG8rHjB9yh99DbMJOmgltY3mQDLzOna5tqK2A6lhWsS1Nm
+KUz25fKqtNJ0n0qP7VPAiq4kqddpTbJ6JlLzX9SqCkrxALuMVmx1MX1I1pF1JaZOAmtWWjwBUFY
/fn0wgc7qo6cy89OEylXjwKPJalB1EhZhCwqVsSU6gf0yRVW3DNkDNdoiMOlbXLg4C24X3hEmbfr
GgtgzrUSxztDTSpTnkCGELu6LwfR/ETfu7wU3pIn2gc7KbyW1/Huie/lEQrHUrhXsguHoZDQkFWx
2Sc3eSBAdUCymG/akH5aSo2h24cIHYWHE7B3TesptjqwdWLtPtNlYkicu72A4D43V6OdFboE7APZ
uR0+EUepOm55JXQIIDSx1dFZHeWFJdFwclOegCowEYuOmTT7t/scHTtYoDw5M8t8JjT9NgrrqJ+i
WpkHrbbjKxe52jMFN0+BcSX4HKJmjFuqsrDdmh978z1AHliBqaB/8VDCSUQthXbulD4SpynJn+e5
//kBsHUClJPSxIE8FLdXSaDnaD8icxHI7n3uRxSVVEPTWv3vXr0MJ/BhxnYvZdsJYDpmxWyiFme1
dfFrU/ydxn+OJiPqJv/JpKlhQlvtmQBVsxsg+eQEnvkPz5draCyYmCtDB6a5UbyYD5z3mBD41QOC
B6XTHDZq7lPBTIWxPl4khrFLs+9mh1Gr8Or2UIbN+gClEzsawzts/b3a6S4XQJ6PxjKslIFCW5Yl
GXiNFCxNQiGrfAhZXxOAv3k6eSE+8sYPDkl/qdxAE5rYQ67bH3g7RuQMPn7H8Ky7GB7llgSRWZYe
x4BdUfDbWdOBdkVIJh8mszl5nWwTueoZHlG18nVhWFWWzHQAiZ0Wtq/M91Xrc2ZyVIy0/82mNvNn
n6zHYcy+X5yVVy/1enjWkK2S3RFvaNyuPY7t3mf0iDDf/CarY/fnK/3QhtYDfZCZX2T/GqDDlAto
v+weOY956ylXo3eFNxQmfUMJV57nrC0AQASZzcHClDJU48DbpT1jDo0KMJ1AgVAJcvDSxeAKtTpW
XQ5cgDK1KEuGIKO/Ws9VareW22moHXWtSgK0GWplhoBvWVKPsmg7/4jtfgTMeafJk6bisargoq82
UaKHmNID8l69aVkQeBkVwnXbk1MmIQBshRUI1n7z3ITI0emYktlqxxXhrcGt+L4lCfDzXwvAydDh
gIhJHJ7JCupZKFImmK2csoOJekHMJ8stLNh7hlGdpCgFkTF6hi5jEe6bagYm8f7pAsLw/6WQdyZj
XRIbFdf+fdVGXYEZqsoFkrPn6m5LPx+WSPmVMWBN5QIQuHC6h1XTwDaYcjv0RqExIBbUa0ksWF84
08/eVgMs8GqVnYC53blZZKp/dVgrE/oZnk81qurIRnozJLZmJr7+/vBqs54uAyYUxTk120BXKsr6
d91uwS5gkW93iD0oNzdOY+MT9RVNbMyAysL29ODyB+kAJp+SpegTj8pj97ecQWO4wQoFqPgfZ+DM
apb1umo3uGTAUrrF3RPcV1NQMrxfivIisHM5G3s6jAIKESrF4FxCU5Fe21+RSD+fmOsS7hp+tcTf
+5R6y4iitVjSx+5Dbho8HJe0PbANt6Y0BcK65NNJ/v7yweM9DjK3u1Zk3EGf7D6erI3POpZzfTqP
NhWSCEH4JaQQX1Utlw+6GhwpjpAGRZEYsFqM7iKDvr/7D9KWIsMsQU0AC6Ij5h37UHK6HVH6Bjh8
VDpnyZHcm2TbCL7Hi9mkAF5WEv7chrySkQfen4PojHgf1QIUrX20Utd9emQrmuEgsayeTpFLgc0L
SgIRvcqoWCulmsgqfV2dK36ptQgtt+kqcJz5zp9FUN2xUTFWw0qB9amV4qijeS82ubiR9f1Y8HJW
nVznIDavIMAYLYO4yMv1PlFf5+T90VMZ5seu7PLmUI7Jw8Z17yATLm/33T0jC1BFLczaNXZzNuoo
0C7s70ofjkfWXd0mix3xOCQ8sqxo/3Ahexk1YZamubVh9J0yZQMCcTmyviUuSpSCkbUjSyY8XnsV
qqkQEOtpNndt2lo2sD+ZnZDobksurQZdgXfQDHOgePGIBcQO3wsv0YK6XpsaLAxlZ29x5FZhhUxj
wkKNA2DQk2KcYMbJaFdLVNYmSEPo+oS3+9IeAEGCCvD9CqEKJHhmgMGYVtF0KhUDLjcKHXnw3WeT
dY+5aiXL3GEiUiC9I79Bo4W0crL8/n1/D4gPsNW5nTc86MrohQf0pgBCNnSabOOLFSChV4n7N3bY
56kzSXJOVuUMvUMbTrJLioTtsS76T4Rq8zoydTGqI909v22lCMJ72UzEnlzqAYiPeAK9NcnK6O7j
MCkqtzXSGnlZHIO31ZmYj0RgAh66Jn8aCVyWnDpynRvvqCdfrfH3FKF/WEeIrxrMBGjsYKLWvrPe
zZfViChBtbdTKJX+hAFzHZS01R+cuK4F1wA29ixWsxaQDeWcp+bsyI/+KlP6w599lU22D7KW4MPg
9V+K+yOedaWgVadQfabqMV3Qd9QpEU1E+PIZ+GWRS7ml9Wa2uH7RoKMmSbwqeID9s4jNz1UHtVVE
tq7dvtFHtNTYiTrOvVNn6qj/VSFKlwjXYPPcyKHfQ2AmViiWwSwTdCsQRjhSvPWPtT6TfGWCy0GX
s5G8UXxvRik5+n+SCXk52zIGMpiunX94F+fOOj5wa6xxPbZXt444SHYLMs/nBPEYxBkVJo+TsZat
awSRupiEn3/1mLdIEO3oE7rXrWXR9XkB8r3gonIdYFR5cg8mmv0Is017NLwT2NvgTn3W+22K6HoU
tqrWWVuItcFqCP9qLu8Y+4mN2pPSj6MEAN9jpBnfVMIc6TQF1G0pAL4mi4He/chRtZspmYR2vBNl
MumutJP8+C+fRrqvhqXqW6LwyDpG2YvQvi/ZPtfShmeFFjVrQOJn7tVTrJvvzLcyAcI0irfZAjjY
TcxfwQxX5Ou3kDin3xpesyMxqnNtXsejSYqNBpQGk+Fr5N7nluB+5Vdikbfpi3dKex87dqpPu5OH
Dj2BtovobpwAtbDlJuNhpQFclJAJhcdvOuCLqW/pvM1Eign5HsZrU4dUHt4B92kunSA6D6NhN19T
jtxTO0dLzesfQy3MIsTcLAySdKJyRcbOVGZsPHmjWY+B2t1Iv9sPnjbXn7D/YfDdSbDfxZC3XsMU
f7GzL/SMIryAidfVnuxtNCgb4qzXsbkgG1XllMqCizfq3v29O8TaXXesMrPHBZTjvgFgRi5q+iGd
R/XUZ/PA6V44eI2DpmcGH3hT6KGQ9JjbYUi/ZN/4wxRNek16rmHy4cC7UTLkZnr0mKqCkX2nXyeI
ma/c2FDjzkoaseO4Zcuha3bNFTu3kezvI2KZnjbwd64DTZesqa3c/ShZe4NbpUIpk05NDOPGI+6h
rn/uw9qW7/1RL0xDMw5ebUw0+DCTxFJSTdQAIyN64VeN5/LKJcbWsgtu7zB6gFlnD87ODoW20aTG
cyitaQh8k7KHqfr4ygRgcbe9wlstJ6WnPqbdsGoXL8lDoI8sE1z2HqBZ78B2QoJfCF6hzsL1pLJs
HJ+uhhgvFeoLvAKFaUAKbN5lLJCn967cToaibETpIubyBJAfaO4u2pzu5466bofyeh/QvgVe0r41
7w72GJsO7OqXQ65bpyG7SzEd+avyJJ+gMXLIS5SbMByXnQWrbyDD5wRrWP5vSpCQ/z2dVpHgfT/9
PJS/URKTsYqYHfgedLoJUOs5nLqYAt/TPGakGr83Unjis59ZX0xzhjU9Z8n029RPWfmSgSgRdmv8
/5aO7Gv2a/InePM6yzwmGb4etTxToaaRx1Z+dr3NclEJR73Nkg8ETRk9YOAQXwcHhAdo6rhZ3MNb
ZCcRtnifzQrdr/cNXvt5uTU4lfcaJcrC0abvzt7caEz8loIiaDuctyy4wcRDI5U/IhBxM2rPoLwd
0GKD5tPfqAUqBEGBu/LMEvzKXILAoo/+KieKYem2gn4Vrq5J6K1RJDkWPhN156bnPEglRtpOx2Iz
Wn/PxzNxoThNRbNLfh6x9UP5pF8Xvf6SLBHwsllmsj9ebzxRyhnzztbgHHslH/eeATs528fcL/nD
y9KQ1Qi/8lar4O4JGehgBQgx5Acj+Ml/qUA61Hri9KTGB8wD22aeQGwi9a71HlyCvXKhhE+aJY1H
ccW+TJZVYjYDFrdd4x+lQI6/WoMfkqGCIR/mWr89l6eYay6ikWtyrXO4C5ps08dYxoLHn2M+0+DP
aQrMcw2ZQzC+QKbrCoIR1P77VFPju+rZmGKp7/Ars981elqBdP8UEbcVwNv9XSwgr6sqsbiuFQw9
c/2m+r493Z5B0Qjl0Hltu71G9A+zSxoT1wTK4yksCdG5J67pvqUwx6nMVxEnS/aa86LO4rrz8btY
wbqWrC3OW1ua7zKCjKQuqK6Tyc/EsSCm82CL1Vo9kYJeU6kcPY0ycqfg3GvtLDt+5tVjMewFNws+
H53ps3jMaV4kBO3mqQYaN9kg4bHGg+2JbsZxGxMdTrN8QmJZ8vHbggyBfOKQE6MYHWNlWIcjEjBk
djddLxe2XrVtNWxABGGhS51bWpaphW1lW8QrWU29jHg0VUlwBZPB9BBCa0VwsLAHAIvxy2D5vXLB
Fb/F5DuI6G40thn3nyR5wGIe4fCRx5Wa3fI82w24bZ5rBhB99qFhjrtX89ZMrRIMV8NV4q8HTqs2
6ezToqtccIdvn9dRrYZW8G2gc/LiPLDk4TYWtZ3KLu5+vv+X9GoVScx2oE3YUDsQiq9WhTH7m7gC
5kjwgcKndhaTwI/ykTV/eoe0z6lYnIsE5xwkjv2mUIcnRads6hJPl8huVqgwRw5E5wReqE8O2YSt
OG5/5gBJ4zy1HTBJpb7tF6zi8dWz34ux8Nq97asYW3kLPHRC4q6jfn9/BYwx5QtKzp67ac1jQiCl
QvgEvge4SRKzFe79RQvA8je1U2KVqaNH8aGHJwtRTxjtLI3IcYTeAf4nsf0CeWyWXJSf+GVA0BY/
USncAF04bSr8KLaV09/KsaFs4JTG7spzAbwhnezEh83gc0Tl868hnDc8WbnrEob7m3Z90RxNJ8yj
tdwgZkJ6rYEMbfTq60OHBMWwZJaofMFQyX5SkY1W1Ni+yNcmXOA0pf7JEW8gkI0h7aDYEtPQy6ki
1vfP6mlHusNUXj3c2fUxmszQWUhzADeuJfdn7HIXFxg0Q1idWaCg1KpYP4ltp2ZgBX2vLNe6vYwr
4WQXfRZEy2g+Bh9qyD8WF5rDnIm3DTQthPVQczRaYvilZp9Y01QoSMmisIqdm/yBgPn+61MPfeYW
jeNFINpXGO443u419zIcDRDjN+cb3yZHqJyNMrW1Evhhng4eB+KF0uOl9jRp5HvIfjrgyJeTFtBd
kuyR+ctY7ULlCqtsgEgnoJUuXM+cDh23LMWTGYC6Q7/eyygudi862pfqkqA5PwNndCqqqATCn4hP
vqlbb1aM+j3oggUApuICWmwAWk8H+tZGy9sb/boP6V8VNq/ccjlMLa9Vqolb1UGv3SaX9a3LdJDr
Dxovdy7zjzXrdnH/F65C4P9fXCg7Diplh6sn3+seZG/BCJuWKHJ6iBCrYMSrAo4bZjMkMTi7FaOP
kAA+hsvesxZsXtT+xN6YC5X3ZA5moFR1zE104ylkIszkN//84r3B/XzqO7tWMSZNM8S0lm/0L5d0
8h+1nSXPQRuGZaxle0Kzqtlm+w3e9T+gYVlmz7/4DVX/lgns6a5Riw4H7PxTKysE7lJVJ20LqU2A
crHdoMlp76E+vmtOScMXB+nQor97981H2X6h+/Uoq8vE0p8XrX9lTeLZZaihGRMSvScmhw4JCjrw
Z7b8rP5MltbWRhloozk60RkKLKMp9OxEJyJklNHyi+DwbpT5mk/PRUhXu9kitOqq92s7YNGbFYRS
zwb/cAgSEFBpz2fsXAbByHpDqBCQMZKkdyRKn6+I4fRktJvJttHU1QC1qV4n1J4sjKoU1T+8AJ1R
cfJq+Nq4CYzGjzEu/HyGmBoFpAEwa2irPmm3Xxs/u9leSJVAQbplRjC6/13ZRgO2v0rU1fOyNJ9e
j5ZZb93nPbXqM1lDWfpYXyQcuN+QCg5TCYpXDLt+xsw0ZiOILJ6jz4ZiKIdRCY5eP4IQTRDkOzMn
gufFBG2QcbAVLpkjOUNFH0AHXWm+vPsuU/iLvBWZ5kAt5Eq0y7GOxKDOqQjTg3ZNq9cUqsnqTrwf
i48vn1p5kHnLc9yDOC7+fgiD281TEnjdJQ3qSf6+aVh33Osup1GLVY5VUGlVJ+B6AjGK/OpMIK11
Ftfa8Ddo2jhQ0Cst9hr4vNdM+ARhOOpVhF+Loll66nMv4MKag4AgMI9cjVmcngpSHIRQsVsvUo1H
EEdFkE4AvqLZesAJ7nQ/zqfaz/BVEZQZJBQf175WXdfxOact9rsqdJ92N488WTQv517scFcMYVJB
dQUQWNPkaKS5UIRtg7PRkzcZt1Oumh4aVqrcRVw3XAjgsZIBYBbbROW3nHYrIfpotVwczqx2r0RD
v7eLkDTHH9E48KNC7Wn3ZYPTmEI0SsEwCkc+n9mD37LBb/vItfiQNjrJ9jmCvIgYryGtvvGLsx38
yRFx57qPGWlXuO4rH4Wh2hCCmvwBZ7TlmSx7/X7pVk1CbzPGxW/TmeR+wRuMdOnPRSatqpUvDTH8
Wa5yhXJfZeDzirg3emYcsCWsfsJOpzf6cROh5UUdqcCKDcv+3fkTJrUx8FZeKjqNq/Mp1cfhNx6u
0eIuFwVLsktWdvY2gPgNvvrn/DZXxoDEHVJ3qu3l98/X7pSdnBVbAFRSkXCtkY4dS86A2hKGiLSx
OCmlHI8bsBNBa8xJAZ8AE76ri7s7l+XmyzupStrveHoLBt9i09/bb4ww35IeZBbaKJOWU5NI+Fy6
Jqbg9NslaZwBs0BlbbU24fNVnYbvHBhkDjiufVRpw6WQn+0BoyZlLUzZR7C79la2hgiWUH4LATFM
G/shLkmgPR1NBfyYtH64iVw/RynqAwKKSUka+4U9Wxr7ivx2cLb7fz32cyRiov7TYIuHVyKDINAQ
UhpXmnhNojz5gde4jxABQarXSf9r5eozKpKSlCje9NEJpRe7yI2Qf6wwOmjIIrXvHMpdpxiY2Ufe
3oUPkt7Nvor9CBDuoJwpe1wudqf+n068oRwQYDTE4+UznoyDEBWUeauqUlrpi5lDNiYleYzePGie
SxnPOG366WFGCXDAKDGAKKy0BLKXB0SL/L+NJO8VyL2jJfTQXaMqrhpVF8d1qEUYptkVwq0eiwCf
YTNjsaCNpx7T0xOUApfkDuh/I9B82KxLUzEPkl4aBsfXuu245ryAZAj7Ah9+QkmiaEuIdRtnHv7w
Dm/6y6XXeNqtZHwXnrMa7QRMyTjfnLvW/iF56etg2P9OBWd9WX8C973SZH+qRnuczzFNZd7FePez
HdbazYiLPIg3oNMFCTcI8McyFQ+ForfxcWbIbznyG1URBEHd1FXOCuaZzGK1LldIKHkEh3nK26oC
dFUC+nlNyVVMDDB8pDoHfgejrrlOzKKcfllKaNHsz/dGMltCXkcS4a0r5GtqR86WKs+UUmv596pP
Db8/gdw7IX86wyf4Hz4P80lLX9Jf86mZpJLaEjVlNPxWV8CI6LABkd3Bpq49e7BQvVb3YD0j8JX+
Dbk/yaAHSa3l8OKLY4pdTPSElccuL/JExnr2n3OuWJBEeWVH/2LuZzGa3+I6USmWCZymDFa6zKwB
fFaWXvjfyyjHxiwyxBnDNJngSbrqxGI7+QdzH6l2d9CHTYpm8/rQo8kpU70Wd05D1Pjr3tKBBR3O
HiTlR1i2hwIEdWA343jhGtrAT5ia+cR+jRmq7CwwleHBLmKmWxk8h7SDJmgTZst0qRGGTp6iVmU+
NBOEl7q6bml0tn06u2DD7oen0CBTC8cPCOj+q66JD3ZD1mUuJjwX47SJsyxOffb9LjDfikVd/zQz
BsI+n/Xb+Xv0onRcV8EsPmRpfhclaT1LhS9eRe7m3VUzBx2Do0t9DMb9PqfnT5VeTIOF9bGUtCqw
jpo4U6tRbM+Y8Eprk4iojQ3/JNEYugAH3y3otLfSvJ5nj6yQfcg891aNAJBo7W5PF5brhVxF3cOT
SBZ89oOQgimnOYKUbJMi7B2ffd7b7P1WdeHkb9/3xQ+4BYw42/Y9duU8Tb8VSc/1s5+MeUwEp5hT
uyO1F+FO2KU2mX8aCcTLvqYrOkgWw5/KGoL1o/9+QCZsEpmAkPuz+KX3H65fTLLi0/QB3dxDr9lD
E3qlK+e9cecUi9emQd6ebQxyCK6SXZAFQtSOE6DMOUZDnMAN2ZRED4mN8KV9zCBcG9EmvG6lwGyk
GLvP/9lsTCd1YjT3wpz7V6OiUXzKSQidnJpV1+pkEl3Xd1ieSMWqHR/LyHNYQ4578Z1v/LXfR2Gp
a8N0yG3g7cmJ5X4YA6B8sGbksO+cq4OvISadF+cBqIygkoQokhcH2GbxKXKSpQatRoLnCKaFfx9f
3HPtsQijp/GbsKCGy64Ew5UWnTpMiFb24ABMOspyEnoMnV1ayBqJH6rry3BqqzOcalo81/qKrseV
49EFe7XwrQALcQRh0rwl1H3LpKKMVDbfdG6du6b6te1xXJ4J46m331vKJ8J8XPLGyo3RBjjH0oy5
Vn8cfWnv2Zu3dkGQqWbZoh6LopLjefM7+x0Cz+PAdNdYiAMWhtbkWMg+mTUm6hXWS3t0yG8MW5cc
a8XSGlyH+cnDbpONWx/4MRDjMxjsCj+sOWITXRbqGUs1JofwmXGC+SktU0yazNQ/4zvM+x9/R0wB
7A21B9rNeyVDF8PhOmWwKdvCMq8vtuQquzQma9J0wDLZqjOFsCY+zGrEZC+4R6ascHKSy8WRgV4K
rYQy8Dst/vfXTyGTpL+D3QGwRxLBtXKYvA+hdZQ=
`protect end_protected
