XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��%��)���X|�������[<����'E�6���4���dp��(�R;| |@)��k�m�
������W@����*��a�v��������̍�
��M]�B��ˢ�-�����X? 	�+� (���y�y��#{{�@��Ѭq�7[�塿}�=���2Տ�ՌDg�.��Il
�M�NR�o�l�˿��6�!�jD5@F#TfE��8Z'�V���HL>Sm�/\�Q��@�x⼰˚I<}�9D��:��a��O�rw�Jy:�5��4�<h\���Z��&���Q�B��*,�+	8� �q�/XLY��Í��޿�0RKs/̔^ɺȄh��y��P?I��QSL�+ޟd���cX�>h 8W|�GE��S�w�F���1�.&���.L��lȴb�s�1`�v,t�w�sU���;�K�#��y���x�R����%�	ţ-�t�}�(F|���e+�p�Oj6Z3��{c��K�/��	���T�dܷ�}�⊀M�N�։Â��0w*�`q;��@��WR]*T80�����*�3%��H��Et�s�ZN�ϥ�+��)t�95�|S#3�D��U��;��Ͻ��R�������
a�x񤿛����U29tfJg"��,��V�Y��Gz��3"�i��4���!�&��>�;DO���ߖ51�X-D��&�@)e
���[��;9�AL'jd?�>`ҏ!�YS�%&�B6A6ؖY��Mhߧ?u�@C	�Gr!�e3�XlxVHYEB     400     1b0��$�%C<B�(�u�����*�h3m�EN�55�6����W�MB9?���jb��Lɯܪ�Q.��z_�s�
raa�i�Lv��TU��+�c��S
4gn��q��OJ։c;	�+�?rџ���	`�� �K�����U�#o@M.1p ~w�[��W��E(a������Tl,��ɰN�X v���k�_�!~����zlevG�E��bL�ry��Q'�ŢկY�9:�Oi�PL�������@��_�X�	3W)a��b<�o��*�5�9u�q�=9�{$G��X{>إK�b�� ;��!��a0��T���:ļ��]�4��<`���B]Z(��7o�;�ZAt�X��OR����>�h,g}�F��Z���J`V����dn�X���r�9F���EJ�#Ex� �N���+�Z���V��y TG�	<鮊�XlxVHYEB     400     130� "Tb�2��i�78~n�D,�8��k;���q��=*����jT�X��C�3�7���K��{u��rՆ��/�L�8Y5)�K�
T�p����$���������0��s:�i�����9>}����D��8Dҏ�~�7�^�jb�!SvYfsMh�2�hS6z�F�U��A������=0�P\����S-��ʯ%>֓�4�`����F{�ߖX9�#U ��۫�j֦#$�`]1�o,���	�$���\��zN��J���8.f��I�b���k�����Ѳ�޹�����$Vq�XlxVHYEB     400     120N�n�>^�!Q��$i�YY;9s+��\����'M��L.r�d�#3�Q��?��4Tl!�׶_��WK�_�2@�$��'��p���=K�ȿ@]%j� > ������)$�������0���<����Y��O0�C�/?�83aP���y�İ����~N�`}C��|���_��:e0E1Q�+$'}��jI��Im;��� "�;B'ǝ�)�<�"�
�:�'yj��ʓM��jC&|��z\o:v�)\�����u��T�����]Č�T˙<O�,0XlxVHYEB     400     170�o9���@���;Ʋ"���жf��4��4钮;2>l\�Gե��Z��ݝ�Ǯ��kqQ�ै��%e��}vw�^2�8kG�v����5�4�����AP%i�Qvf��K��^"s$8p�*AI�^�B�����2
�o3pNf��3�̫H� �X�wP�v ඕ۝�Jq�/q�r��Qh�U
�)�����	�ܗ�/m(��"�D(5��.���%w��:��q��P(_�Y�R�~��ؑ �"4S�I��A���0R�Q't��?6}�]4�I�V؉���ЌBn�E��u��Gf_���?u�~��E�?\�;>$%DF�+\=������$/����v�T�d߉r�l3�XlxVHYEB     400     1c04h��4���r���Aqv�ٿ����nfS� ��\J�O�G�0(ZknwpII����*U`��9�.��tRt���G�C��&��f\\�����s��{��ĭK��ƺ@ժ�:6���ʚ�D=CvURT�*��:��U��P�x1fсvRIt����LƳ�[e��i/>���[���+H��|���˸��O��!}���[��+ېs1&� ��i`5�2�Ix�r�|KT��+�c�������D�rjH�{��}���(T�~����ى��tӐ��VLe�!{{�Ak�	T�#a�`����,��5Y�(.:]m�Y��<f	�ѕAq.��&�{|�/-@q~R�,����©�Z`�}�Nu겁�@5@�$����"$�zX���JZ�@l��;pW;B|ۉ�4���P�XlxVHYEB     400     170��������ɩ�5]����y
����i�s.6��e�F�W�-�/':��3�T���ʦto���Gs뤙a(=�(�V�;��&M���dl.4#(o" �'��[�
�)ﳵ����:�����Wc��DC���/��Dj���$*��Oa1|��.kp���t[P����~���b8}����$ݵX%�٬E���h"L�f�DO���H:6�%��wr�3!�I���R_q]��[*/A�Պ��>acs)�[��
������o\�79=�5�gg3��F����ޙ~�L�Ν�O�i�.<���gs�{y�hlG��9�ˋ�n�Jg�[lb��%w:���/��-��@��俟^ qXlxVHYEB      5a      50(����E�x4�UM���rr�Lj��q�Y�/G�ǲ9�B�s�j���(7LH�L���T���j��M7�����?���