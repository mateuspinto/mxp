`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 100176)
`protect data_block
lWky/TQvyArhc3XxfAFCibqAdpOQzvtzR+O7LygatkXd14AeWaIEeba5eMXArOjGVw/mEie9mB+U
kPGlQg1/GIkCObUr+LBSeeF1Jn49ojfUDza+tQdM2EeQ+Co+JyweoDtfJ5fIwuJV0YE9NecUVwNm
gt/GPNAjp2vpQNWsxPy5MEuXw33/imy9JQ9nNeonI/gKkq+El6pZnZ4lQElOfhpXaDIa8vpNsaXG
iTCqHt6XT6vom3kvnW9i+heoX+QIOLfCOU5StqjP1mFbrJxvEzbY4dK6AxS21tECTcpvK4CU0qe5
DsK7SV5qUKzeJRyg7c97cq2xUmR8++WY6tJPHhcSagzpCzt0JJBAmeHbveduKtVWCeDH4BH20Hp/
Py/up+rO2BqWMfRNvEISlSLy9jQikZwUq9gfH6QIiUKbTWJXxCa59dlNhpV6TEG7tsnS92LgBOHq
qJmVpvZJfw2fXBYF85KoVv2IgCscqavBEtdx07PIofI82AIWjbpxS92w7j5nooXuBm5AOnGXHshn
XJgBdeNaXde5UEjxpRbjJ7BbrL36SORr2kmMchiWlM+ie90rXwGda0ekkm8HcBUKx5KA9vWZtawn
7NUWmJydBoiUknsfS7P4HDy+ZwB6kXxgWJGYBniUEdM76SIpYiBmA2Snhd3k0Yo2J62khEZpbjVs
w0SN8ivJjo8lCv4QhXg1AixCeNVDtyhJZOaHLplEue4GLUYI2LrbZRlBAKZ1nNwWURGeFwCiKBk1
OLyLG9TgC6VckeBdwokb4bFrGrbXgXY96tKPYtImZMlyxMydIcUuyY3+6cVp9md7tFNFTAYq1N3s
A1lJDwYqV/Z4/J3p1k72P/y6D6DJV21H9Rib11k+0meVfRfKLNLqGioYdJoVq/jxsYDIp6t7vVrC
ABcTXvpsz9ELSETUiIOx5naXApx2PyD0hw5n5NgWkRRDgvafAxWZzimzhRxFUwyk2s0AsaNcHBFF
+E7hJfptKCXQAyUxYAptnzwWxZsB+dwXcFyhALXStFvMknd24lSz3Sln75+OgKNLslBLazcjAG2y
uMQf6ebJ+KLT04fl+rIBpvF6vm9c3r6vUT4N6R9bT8HRDuwgy7IHVSn1P0M3PRfO+RciymIemUSv
/QtNEla2BnXD/rXD7sDOm+7eegEMVXbNCH9noZlTkVkJpecZfwzb2ciHdi4CljWB5syz/eDmVSmv
vlCeL91/6oOiVobI/z4moXQUaGZY7ZXxIGpecxv8aYFJEYStPtEsMh9bWvFdhxOu/juqbdhYcnXY
1UN8GgZKb9FCTgnxkIEKMfxRjpxBGN/tfZTSsa1SA61jvFtAqhTBZABKj50sgS7a8JUipoJaRUxM
M2FAPNx+A3H8DYhk/UARdgzmJ3UR2Y/l0/75GZU+oiHnGwYYIfPU3ZdxcqeeXWLA/lDmnP2xDDep
SehI0uCEHoZybSutAHDck1upgg1G3Gfgg0XwPGjB2yljgMQmswfoKawLGpyyobS/5RjvPXlq35Oo
KmSK8YLsRNS06NIVkKlivnOBL9Fqq+pjHnXalVnQJXM37mguiT7M2ctXkIiAYxCXolWS2o89Bxtk
88V5XMRSVU3DENo5hXLpbrr4DJZVwZPXuv4v1N6ql3Lnmrl0+jjhRKIyO3gFLsmSbrGXEBWP+dl8
U/UxXwxrKyK/RSsclMfKIog4jDD0IWf+rnc+e9WML9hPfsmj5PEIUZHqb5IsR3D3U/mvmgpewEse
3+A2te44uZveBtNzwM7Tq8ST/LaOgpkmKXL4f6j0kJ3awjRj9ir3qbqcGHfDp6GI9wxRsYVPnyOB
QYHAKdPhAShuOtkhZtcnJ2gSPyd6RTohuod3+mpLz7OmWStLU7mv+rn6UWx241xduUaE2ByvyQPy
zqN7yuh+SJgwqv3y5KqW8wDEenJH0818YbJUzwVWn9eVdFU8kjIKqoVLPCAUn3bDaOv/RyRiJMDL
vHahmZdX4oDaHPuUPzcaeLzu+qyKV3JidOJcf19LvV2/PCAy7Ol/kdFbnFNh7BcgB4cfZSmyJHXX
Gxkfj7vWBzJOt3VcYumAfw58GSmB9vquYcsQ78dSlYiz7GRfOTrgaY80edZMTZ5WkrSesH4axwyy
Chgk7HRPAGwCzwkmTvcoA8gLtfwZbRXF9TEsuTKZ6H/qTTM/2QymWsQZlNb6afsU2ceLZkC62NjS
jeaCNmRhAlGbGBPJ4Sb3XakQzAGDTS+cuHspFah0zEViIbjBLeUhIapEC+YDinye5hmOzZ56ESPA
MraPlUazCiaEwhOOilx6XA7X5YtqiSjqbiFb8uvgmZaK83OKpflrh0mtvWPUfawPv378Dy18Vxyg
Tba2a8sYBVEHOAQmp9iRTv+tm3OvAh8GUvZorZu6re2GO31DPRK5DXReKqUVsFltll+v+NmDknNW
v9bZs3077I+64wzCvgm2fCyHD1ZkP+rtajZOjt3UMuJfI6wEpF2Y5xQXFqlIlC6tGmPn0RS6z6ed
Bvbn5sbp4IB9iFKuWtKonN/9VJ1L3EoB7+IXYBHM9MnKo3jkU7Gc1P0K+PiniJiIhmiecKJP1LpH
uGpqrj2VRqG2Skw70aB8Nk+jtw6uVK3rqhO5kFcoFyWeWpom2IJzdbTyujZVmQQazA1lIZG4UyCl
VHlLmTDPepKzzesge7n+l6lmfR0gvUlrKSToKYw1D9t0zDAxCHJUVVEz63w1F/iTJX3MluOUBEKy
WwlSt2k268MhPkOB4zbvgP61HYGsXdE87g8qjtPeJY8snR8Qr9aI5i8vOR3jpXLm5qHqV7GO7exE
JPRE165n57nh/bP0GuMF21aaorwYfVyb345qKpcevkoAO9OoaQm5lpKOKVHp/XaxSY/hMTisVGiC
WSlwA5SXIpKOoubtcpFlcYshxRSrgmC5Ab7LikJnajq5r1hOmbGLdH7zjxvUbTZGL0yYOPnScABo
sWxmurMOTbcTzsDLZ7KTF5Oku+o/NA/EhiqLOgr9Ueenq+B5gfzWYpHyrncMJSOIJkehMCRpIvUP
mUuEzHwMJGFTXjwrsjRK+XqwaWV21ZQ7RBgAiCEpPJQkdvHbVSKrLqxIcQDJmLz6f6PScVQHmIMe
pG0dlhiqCMhZlCLwI0wPFajEXLK8v2OobITyFzmoIL6Ce+/RzWrqHkK8hTQUbWcyRwT3q4q1gh+z
yRBJSgyJnCilQn/eRvy38J3yTtzdNidcTVtzOMQmryhInQvCvNgJxi0ltMka7O3NXY7DpYVdgKbN
9rdRu0BgOvDwF5XjqdFdT75/A8nA2G5vjTxoVwV1GFyslqIEhSv+nhCgJy2xaBZ27PoWrNvGmDcb
eni5civRsjw3AA+i4kWF/ETmesFls2u3vRVC2CBdKpQaLwwC6jlqYVB7FVk1SiL8ZYaX8VKuXram
UDU3gNZsodV3EXEfZukUOzgTp7deWrjkc5S/jINg4CBf2oHqiCvZ6u5x77OZQ9DHFTbUbBypMWpE
2g/D/yUa3uHzmT4ZMqQhiNIKL3+Dkpcdqce4/y5+uWcRL/kOTWL6UrOZrDdu/HKca/Kl9T6RTPPk
sn009JocsW6ezAS748sEUyw+ABOxQQbqPeJb6cdYhe2nmO+uK2H4068LJltqc6wIYCbTdLWpEyA7
9WY/lPXPKAYFzwwe7mcIaKHTLAcTCR1qtqvHXP4KqZJsIrCnCpzTjZQfB/JAMZOA0zyK4q7ax6D3
9IXrGhPM0ddtrgOgkM/aG7ucYOyQ/Rxdf7yAmt3GDHRB86luViUtvJLFMGyz6uAjscDbe+vYo5yR
k7NmokBfJKtfjjzOn4x4s2xl9JMXWMQjRk6C04PPa97sI5ER0D4NaGxMZUQM5UjnoSuxEsb3Tazs
fslpgs/GovQCOjW2ZxytrNYCRDPsr/ocMng0rvRf3LIiqExeM441vwgBzn5WDwLD81MbSyWuKz5v
lPzeAL0GKA0bL01QBze4zRpvpvnDBWkR4xjmvuhVVN9WLCKfYjsG7XumcbDi59qYyITXaztUgpVD
ZunhaqF9eaVLC3i3xqcB6zXkt7+T4bVtHGIGexkRfpmaQOlju7ZSTJ9z0qXGaWLCZ99qlvZlMe4g
N924YittNYhXAHOt/I5ooat/LW6NF8/3MiajeSBykHfH6NlYHwdi5xygWMh4WemHGCycxX72ESSc
z1wwhbvmJrk/821ltF2FG8Q4KclrcpuFFt7RPtQPUJsN91V+YA90z6gro8zWMz1TMn47o51pSvDc
QNNKHkdR1PSAJKsIKhCz4EXRbB7+0pVGTPaE4bRFhA01HGyFsG1AB/ub0TX+iktNgngabXzIYoFu
iSk+Hc0wRuH9tzFe1EbK7FdG/vdicHqpt2Pv1JbM9RO4Bbi/8U825rnnB8teQk6A/J4VxiZRvb3O
IsAhrgtiusFBLjn774aX+D/HHI/DsJP2I7cDVUQvAfomBX+RPAIYKTXozm6/ZqLU6Mfl9LwoG+VD
QVFnqW/S6Ww9EEqJbEcT3gdvfujhdBQlvZ/zty4EYINGD1O+XXlAtFFeKhbpmrtFQUeod3xDsq6Q
iFhXtq4jlMlD3D2zJT13q+vWPm77vgHSMu8Vf9aOOvCjDKmmoHPizLjxUyPitQZsj5E2dJKOBdLw
UaKsWF8KzMc0WX5B2OSEdmpbEs+Hs6hhIsOn9MuWTQnpQvwCEq4reaqruCpYoxPcMquOkNIXTt+o
Zjacy307zXHMjkYH8b37UEgWmURsgF+pEg+2UVw21IWcemUFipbveppe+k1Gc9uESE55XPgwYss6
17unrrwQoElNvzYYU17mKJWmjUGpo3tM9C/h8o7IMfnZe0Sbj9jRvZRO8XNDnqtax/JkgSay8Qw0
PKuWhp7BCOYMb2YUIZ1nMX+k6NHaip1ezq/5ljoH1bebcWQfPCYTdFzumTrl6wh+G/CDr7z8XLs6
WwwQZ85M++rU/n5RZHNm5/9duoxEn70w1zzoYdYhvV03Dm/d3v/5sW5jc6xZncxfZ5BKiiikM9Ol
QJHbpUwu/HuqwVLkE2cKXUFJQ3vIrj2g+DF/5G6PIhUBJLFnk9wHT1YZa4OK5IlfDNB4AxljsJTI
PM5SqRV4zTEhrRruYp+xz7/sWr82ICVNKfCbCk5DSdV8UGUBO6qQ2zsi5Wu69enldgUpGcHgxEas
Kr4CDcbfqvRi9JRqmm0A5SpVXSbGRaFNX2r/wJdoh2V35aR3WQDtTv35sEfIdLqpyDQkF7IXCkFe
B/wXOWOKtz5cnemhqDciVl98oZ635MA2lp4L+SPKHLqag72Dkl5TlsWH8dbpeYcsnuQw/Y08YRcN
YvfeEeiTySAEM/YTL8UKJ9FarQsm7WSTSWU4MsBn0vk77OKtJ6Lxdz5cg5OEqqZWDMunQ5D0NKfU
oBDYvl8yU48vpwZEdI47RgSItOcUkVazMZ32v+9aCFMpnMdgIW1yqTeSmJe3hWVr6i8yXMrjtUrb
uisNn1vhetX2RNYk1Gns9Qm0d4oLyhaLo82ch4c+nHp3MjyH8M7T/2W7aFGPkzO/rn36Fl7Beqh3
xLq/BdaobIUEP3RYfeFf4PVtutQGY28gK/LPtDAarzsP/oVfXEn8rAJtMNzrl1eKBQadxpguGYhY
M9wSM6nTw6/qDyzgf9UTSKM/3JWCtMjYeb6lLDKA3fA/MCOB8jL02PpAevN294MOKBDr9o08KTPz
U/A6vGLJCVmNOIrQuzY06slgRgaO4A2SegIZ79e4usRKsEqCmyqiaEHORzCJj+mn9smS+rQYhSj4
uxO4mGyzO429weI5lHn9E3e9t6JUDH5n4u/D26J8SPXS8xeqjH7282rxdsxwSEmtcuO/vyZavF8d
q+zQNB8H6n768URXJt0rx92NpRqAJLLQUXlHaAQf+fi82d+CUBazmH7jBASkPYvkHhong/JfoxdI
teomXmRnRqf5ERzEf+ogh4uJkYjJEsYddHIoBqVXdk0GjB6FTwSY07+J/JODp8HV1kxR1phjhPqI
80MfxMkt/L8R4F1iAo/P+/hHjtnLl1rhgHzvlV0klXy/+H0tzIld3nnxDqWzOHYpm9PHl8STsgwL
TP75SzBfnh/5ew0hcJ3X7j1vRHnxPcZQBwmeMYBvshQDBLuTSZ17I5HtiGe1M5tqaZLg2Nref9pS
Bascp4GxSkPfVZh/th02BLQoK2V47J+yKsYtwk82VRRMIbdLeMrrSf/q4EBW4qTq0RNU/r8NOBXv
tgADe0zsxe2Rx4WLPku1mrKulakpfIqmNrD5v+SwizOjElgMwezsOxu91IjQ19fK/9UbBsvvSfa8
K+L067u+Nt4BFRIfqVhBr5l5DLW4HjPVrpmL98MK9C/HUZij0751rs8cid9kUUAHM2snf6oSR355
+LIWncthYAIa+YtkoWqefjzjGVbNDeALU470ax185ihmbXBqtAT9iamy8sHh/drAtZwx2zuncJnS
ysDxAiE/pkVitAjBTvrHk9wuYAekPZJzNl/V6yipxfL9cMBVhmuvaVOw9g3IBpDQZ7tloAc+VONP
ntqEGcGkhYyQ7Zp+VPxAMrAJqc8T/KnTENqedxMdNpUCVtb9r6N8T6kkqbpvJKw5meplQU0yMRci
DE37KYOWVmGzYAuRD4iEmzqURBXXxdJo4Spz4C3NxEOiOLVQu/EG8VN/nmmu59xPyGgegsh/2q9H
lZ22alIzrCeScAX3dBW0RtKXoXePfuFdN0xXn/b2lh2InS52aq0f8pY0N7PDSYwVG8SVaEF9gs6e
jRG5Bg8D4T7ZYlejrNnKRIfvpc+3ZBnQH3RNvdPuiD+TyDO7CWTBR5xpjlBfZU/02zYZEYkypK3B
IrgeRj4Dlimky7jOkO21ra7KrLub9eZ6iUaJeJC2FYoxxAd2nfDG1TyJWr5jQ8JTiZ2yw3URrmlX
bfMPR8rkqjWZvECl3xHA6hiGndo24hUoJtZdGhLUg0A3X/xBat0syYyfD89CJsXfpfDGPI7K1MLe
iLJ2eAJ+2yRhf5s0ZVVuHPIaI2nTP5ZE8t0IeXs/Z/znqj0S8djxB05dC8EWCiMqMGkLlbMljD4R
/On/yr+vWNVyD2bxyFotiYKy4G6FXiWTC8cfR505j9x9ReHj75CqpWIpTZ94vmAA+7gZsdhupCNX
QJ9CWDccDXS+f6ZY1/iBTULzKW8jV/34V+9aaNxn7Gv5DpASNj7ZDiMLbsz5O/zI2q1vQ2I/qfnx
Vp3mgv7dNrwCWXWCBrm3/IeIWlPrLFxFRhiwufrqTYUkCTLh2XzclSLDEdN0+DllyMr6NaVAY339
eT1D/2FnOigmTfQeu7rIWp/3p7nPRHbc3Ba8nXy54aYupBMypJxQ94mp2BBGXPVcxMylTovNEnRS
TcLz/4t9gVAPgVyaT/G0jbFpCTlCu8vtPQ1xMVSd0Sy/edrSVTx5SIzC4pECUuP9OtXCD+uhGY2m
IdcR7mo0eC2+hyN6BjHHlu7tMvjrqJa6yg3aooQXedst8k7g+Rg5nfNPsxZtdh99/n3QQhC28T/6
Jm0lUdL66YfLgc2BPz6MQ2inEHcnqTgBSCnntrDw50xlCOIeiCHusYtFjyowhvO9w4RKrDnQ/B2Q
EHjvXK+9fh7ePQ5YgcGo7+Hgr/c8v9lXRexaghedOFcUdAqUq7JQX7zv5XrXkB8pLbfRhxYZUrNx
ZoZYo+/1cv1NJCQgq2roHctAU4Hb0WMao84Uml9jrJslvPJYC1uN0mbS7WgDGp87IHNVyosxYiUZ
yaPvkQxmNIofCc1O8vHauaJMGIXn1zaHRof3FgkN4olDN9nL8ThPdBC9jL+zx33Pt3svyfXkcDRY
s5OhEizvUHgNFEpChcOBtqWq285yjlmXk0fcegfr1DV10WfkpzdmYerURpkjnJViTDHQ49jCJOE6
gt69Zri8TX5usqgcweUDOzApbpGyW3pemkk3CV1ZY5oTLLJbBSPlyS5oqEUNYK6O0dmIPGNOqGdn
URo+WY8BocKDphIx+sHEWnSLCRptSn2g/u+2VXXdXS4LQJbLsLPksUfGj+xsQpdSsGUPdJdI+VwB
SbZw9ceyCwIyen3p/GrOzhCFXhxVah3FjvCKnKENb3LgvUmR7/TY91ysOXARpcXYHeiAHxrxZY4g
RP3lFCxL4EsvcMwOKh6bm9/Iezkvu8K+xAgRWt6E+6khsMSrOfOb2wrWrjRXukuo3DvSpMoUHTOl
NtJ51J9dJj9rTbuShaXrlWvGn8tta3yiEW6HoxXlERy5aYTEGdH10ylPppmpjeM2wC9VgBydUCBX
8WXnixLHdL6UPn/yr/fr5RoR4/7mWYgDGyLqC1pO4/DUEOx3KomltlucxGolXoQgDxt63g1MjgBv
Sshm573casuihgOxbyfLTsKBkspjdQLjgLgceHhk+1SBDAYa6IVN9RBtVfp7scymuBOM0+bdGOPB
E7u/ZyoPgTBebNipb3JBGkxN4dNztTNbFZLMaocRpCpTOA9RpIWlB/TkKn8/JyXvqoVsBKkvscIx
8FciPNwJ+CIbNtK+K4bVUOk4S63pqvDPoYIbsM3el/waZ3FjaawMGvc1mccQWujriRToycfCn88H
jmZ3jxqibSaJR6Vz20Hj3M24Sqr0YsGiT0rn6DX2aFPnEnyOQywdxlctA5+w0vhdDOBbD+6UgOzP
/Nv+exzeq0PhMGanfRSiF1FpNZzcO6KFGbSeVHIY4co/gU4I9CftdHckXe8b+wRIeRoCLwRz7+wE
y3VotW7ohVUaNd27+8LmDsUnMhAJuBxXXY+J3dBkV/p42XWy3o7AprZ7Ph8Mh9sitmLD10OhQ2mf
Uo5ehc66snLXR3XAhuNQrRZ9sJPZ3CJhGF6Xo3drk0pbRd+QA9GMtIoZm4nKrTpxyJ6NaDOlfldZ
5ZhqO8i5b1c4EJmY4ojeInTlW79UEcYECTnpdvh/nga9bwV+VedxobLEAPeXBcBzEFCrN27Ror09
m1F32imOtUj366lfXK34EZ9NhT7QXXAJg774qp74X/82ID0ypEl20DfmQNiXoZ7mrGKXPYiCHB8+
v3Gek+LVGiJ5mkgkedjPNJn9BNCm0QVtZ6Gfo7ed2kcRgYIecOkZG4Ar3HuhfY8YVM9iatgXfgKJ
YnZEYPZ3Qo6GwvsW3B5Ma3vffNeFSGGnTDwcZ4HO58medJ8T1aH6yw/2hk+LcWgPDuW+tklZ2+69
A4FyGHstvr+IjW8B0cC0Ko0OW+uuySSjNlmO8MB4AZ1kLiUYUhLdUnSsSM4TJRx5jNHN1OcO8D19
tMe/5gpJOAYVnQ79BDq3Fm2Nops3ACu/fRNu0M7yPYe5WgVhbZNnBLudRu65oR1y2eQtMhzwmJx3
YXzX/egtIwlzmPLbEAYmgNQFvhJitsD09pornk16ovroUv88kh7KhdNRvaYLMnQCxM6HQn3pkccC
f1lPaiHXmqpJtRuReoYHOxVKFK4hedeRf34uIH6xZN9fXPgCm46IpDwlhQHDsVaTkO6zugpSIqGL
7Rf6C2ogFer5xt6tsv0eL1Alyk+afBHFFAp0M5MEOI5ERL3zeQzcESIi8HjeD6C0dAHKEE3382Q4
ecEGLPFYHK5gMfeQtzeG/qKCF+rtwUXzy0gp/B2im7waUGUVSbN7URN4dCtVAjiehcFWPydnOrLv
A/ZmzM0jayg8iryNCEnX5p3zV4QcMQNnQsREK3KvKWFQt0j9176JImKL41G3scPOA7dUC5GadGsn
AU2m1V/dl+oxKZ/W15h1nAjFpTWnQbIOwzlB5JAtH5GmPUoBOAn8t3/gub6v6w82SvIwJVYIQo9V
n4KnBy9zKCgTyR6sAN/DPMV143L+ok0vuO8pLGvYHfy+UnfSuVXOQ4jOzeXZJFcN3pnSRuLxiK6j
j+5D9G3xyOoo6np1UA8BXsedwll8wU0E47aS1Yd5U64cNMcxPLCLZbwWKEekz03Fj0l0dQNHCF7v
n9osY79KIct4ZN8AawfmthlSJgASg2qL68f6jYmI093+5SrKQDtlzYacSpkzDp5MNKLwT0b+y1Qf
4Xes2Fu4svujy1XqILKLRcJ+2BO+CqNkb1HAaPXR1Ju68f67B7qig1qZnHJkkkyEKP2r0OtUrQoF
7x0TIIt/VbZFVeOKcRISXsmx4aK5h6o4jUaXT6hJGiHoUmTDOnRNYhHvTB/W/Q9EMOVn2tEeQnN7
kSK2TF/9+kf73+f80FW6Ax8+xuXh9DPe+BgH8Hgl9kwhmdSEKbV8IBj8303Yz4vlBkAtrOyX1+lv
WuqbthWMMs26NVcjTNMX5JR1haiVlXw6I3HBYqp3iOzvzigfPfa/gjwrBTtA+LXNPJFoN5q6sQ2R
gA2pWELmYD7WEGTX8doxZC7RMPP97k3icCdUgRm09SYW9QiCWPF7LC03q3QbPyoIgreqA9kGxhZV
lRc1zAwPwTapKIsNPHj/LMTzJ14n/r+367W04auuSqCOCeqodXuBmeEcoisgVKJVsk4vfnMDAMMX
maz5CKySrTFmo3RsnGc0ZVVTVV7BG53TkOthALc0kRly8QH8zc2vBSU0tiE4LLbf46P8ms16wvy+
hoVNht1S8g9Em+i1mlpu6aaEHLkK2fQd4KMGc8oPuWZA7VevyPrO9l3Hlhm8vRqioSo6H5bvrpI7
w3UIeq2sh2rwZM0zyU/+kazChpBO633bcwgAGJmoCIx4AV3WE5M3AvDnLB4CJLjbiVVrRCGeZ+/q
c2DvUecEAZxd5sootwHfAnRrLFPgcySKg3aXk6JUJ+RCH5c6aOkld0IXm6bKma/p8rHuw/oCykqt
jvk0itOF63utnzibe8levSw1Vl3Shr6mnm9utHJTeMn/HNKJH6f5/wxbapdoqrL3XOeRbv3cNAtI
6n9E6e5LuO6e6lPW8JrqtSHcFkD+thqBpGctNGRDdIFZRRVesKdhgFetud9NBnVf1D2j7aSynEfG
aEnwSNMn8O1NN1NaYZcNvNuEOgkcJ5BzcG0njz2wr3cjLo6JJ57VlBLi2492X2Q4JfAwM0PBc3We
RFujc19Ot1kV5diY2sjS10WjvIcn5MHzbQz6SIJB1W1MNwVf+VnM6E2oYKKuFDRScfd2Fz6YlZ19
MltRUQUmRQxDPMtjW3Js7yCgyQFqPCoEHk7H+53Je8QsmXgQzV76V0Rq5COIgve1CMmLR1+Wc0c/
Xxt6ftyon+ld0yWkFZ4r65xncS5UeHzMQcV0M6rCQ94CXOK7UfiQI6OlOjjIBczRD7vuAIRo9nKE
HftDj0Xfg2Al+ZdG4k4oUfrz2jPufvg3aqtChpYBPyoK359/aTf/loa6nvMqjc6ZkhnGQ1NwGhxf
8UcuGviLbC+qgXHfWFdq4fkST/2MIEN3Ic/kHQj86pXpZspRpZOP7roaQ3Tf3tYA6XZhnYsg9M8x
bNFJOc8cB6sJnus/e3Bvncei1rKGHCAQKTh0LREwsJIFcCN2Z7vo+KhfyZYiy0bnYvCLrPhdNZ7m
oarGgl2wBT7kysTXsMz6JGqBq8wgHugHvatvgthsZt8vEyHqJfpkGflDsyFmu6JJE8m6z+riNqJR
QA+boZ+Q/tOVqjeP6TG4pnsPCBeM6IBlhiAgKiDBt49OkIGDfKfmC878XXwmzzWhJKtUs5eED9uS
Vf+bxIcmcWFQGtlrK4M8SgXzxsMRVVOLaxPaUSBDgLt/2YtHf0oko4mLzGgofxO6tzxtz0l0L4gS
MG+1XNi9rIHCg61N2nEDAYn+nG10GmvZeubVNlINkuaMmtxHnlK8aLqNzigZybzntZjXd3CGEMre
wIRT1ea2MGkoznbVQDm9+lTmIJmHH9t4kEAt28BZ13KgyAh8snS9hGlOo21sPqvmrVvgudPbH2+l
WfqkieONLzFW03hqhiMyHYqlYdgXH12Pfh2KlhuGUZnqbMcVYyrLZKvkSQNiAMDAK/fBWyD7Z21s
qwXHEyoDESkh9R2ICxEv1Jx9UGxOuvOmiQepjgZchvyizbNRXOWsjkVpNd43ZuP5chZWM06t1am5
fFBEEZoxGCUUZlHRvKM+ZaseqYECWwJgev4HF19kOnsi4ESQwDZPwfibXO/ERUDnBH2PvQRigPW2
Vp3AQymISlIn3rI3yqMIk71sN5E1nnjk8Cnif1CxH4wvAgaCQPS8YTu14B5/NUjYS/IjSJILbLFH
TchULuJd7RBXjsNfR1tYtWI4KtZxsdG2SGYZvVT8AnvY3nPl8BzPP39rmrpF1ytn60wRsIg2LDgy
3gEtFELz6cLu+XAkK8bYcvvqR+OmpaNkYyR99/Cob9zW+VdhxuWDTt0YOiVqpsfTkA5shw4cj/nv
U7onTy6+B9E5VztsMxArclJYBP0TrLwOVr2Yx3QssyRJ1cJGtjvmeX9Obd9dnmmHqRf4XiLiT+2I
i/OoPpCHdYiSeqQyw+7QXTsuXwqsi7AO+V0vmwK5joMHdXd17g6enm32pcznTxKOJtivJhGNZDbO
H56qYhfW4kVxeAKqKQC6wEI/EoLvF7Vp1Po4BrYaCajZxNVV0QyhezndHJhHbijmTRssWKhBQuPR
OJP+Arl59Q4ROlJa7JEdZQErHIFFJ+cbJP9+LHFIfxZtNF6E15kNFKgQmlGtbiMX5d29abIX9Peb
ILz4Lka+w55G5kPMv/XsLXI7gG3numvWJE6EVh+ZDeFfaPGz4o2N+Ix6K7pvOX9N2rchEBpUUiaJ
d2WjW2UlTZ4pSkNb0Ak9AN4JWjGeANwwdUEOxY7Up76E40MQGluFRWuqfkJ0Vic/fuffwZ0N4bm1
DUsAnGPK9C66QgiUKkGzqjE2+EAhwnw2TafGGOHT8n6RsMrigWRKNoE/kEGSngd5kE9FuM2VQ2Mx
tqOloI/3cbY31trLexzFYEaUA0qmUzX3ZKfCRxoa1KwLw11e90zVddVx2KPeAttyCFUcsO+QuBgY
5kGK8APeN1jgne89PGNTELtLqC6btan3HDtwcNdV8E1MF+mE91MdzZ7Jt+c3I8R/VG8v0pTLXKFh
DzOYuynxsvsQS/rQmrQgFKmo5u7xds1xHeG2PjUS/tsidM3rFl+L6zLFw/bl2GiuErBD0yeIpf1h
QMts0FGWPbaIWRoQCfOuDTxYn9FMMKVh75OjQSbnWDcIWi0klvTF6NrbtNPOrO517Lboz/XnLP8l
4IWhTKW4eQHog8kCDtsWbFeqa5guMEyip7ETeUS6FjdmQ2bTK7+ESCzpzumjlfO8xoN5NfjKRkoc
DguaG9HMVOTTbs2lLcyI//H87kCgTm6F1j/VPKXSoLejx3xakRJYWP2qgu9Y8lRIjqPyck3A6/wT
b8WIxMBsEC0xeJxy2JN/cbR32ZowAv+JbZpKx8aRFsVOYcHrBY0tulEk2ayc3Rba9drtO2Y3Bfe9
DrnkP+ocJie+N0tBkcFpEjbH8OineN1ynEiRaJU1/vRqTG7i+GcuXHgmo8QuC+xHvp08KmNwZ3Cz
a6CMvSCF4NalHCI61lrl6BJbtOQ4ttsJWAXEEl2mh3LdGq/bA38AP/+5kNgrMKL2ZVsnr2kTcXT1
B7TpZIxlx/3TYA1o52//jImym7cOJaHwFFeNC58VfOuPYJ7Kjy+1RoLIllED3nnVtU8px3wXm7+h
yQfJBq+4tU8npw3TS+PK5IFdSgyImuzIjalEt3TetBKadpw2ecmCgf6B+3aZk1b4kaVb6lpU+OsC
N1sI0c6TK+N5UgkFV5wBBOdKfwcO4B33Jy75e1VjsuHwxb8kgbUKouBHgJOYyajBfhBjipeSGu9H
bu7C9qK/Ni65vfXtKsu5213nILThqVXS+EBCVQR1ZxA4CadQBxAROaJzuvtwhYlcBqbWK1Ur6d/p
2DO50y4WyWIvHV4KHoxLM0lGTtGqjl462kH3HEEkggavezBqANKxImK5NPz0FSxSAGx4YRo6GInn
aYfkXp7jUGWuXKgZRFHq8w0eZ5gvGpj/shrQzs06gV4hGk70M8DD2QI/WJHKo1Lqh6VuBztY+PKw
wdYX7p4bMfkOvf5+QVDnWCeBYND3oK5mCbeEo8tB3yqxpdmzphOasm/g/BFoRzSFEJULRR7ri4FP
bqrVsNnVWxq9gTB61vSZZoqbvTzFiWOXUQQCsiAhEMRWutF3d7bq3s1D8Db40pWSzLHeu1Qifne8
spmeO0wCLzn0mxrHj4xXCdwpokVlAt/Ul1kOEDK5i4zK4b+hocHd7GhZMRPuznXQE2Gpn+3pIH3E
KBv3jK4l7qgHCn4+J75lhsaSAAggHeH3LrsqyL4uRXOcrxXbxNE1N4JtsbzL3g1+Kiz4VUnQOskW
fnyqk+21tmUMnooQo5eZP8S4Sbk/LJdgZ7kzgWLD+DtPGdnHyqnbA4aX/8rrQVN/pSmEHhy46yIl
pongHcfJQe/ze4awVu7J5vxak7Tiny+hZLiByj22RQwL9IhoqjJAEcED3q39Jtg/2SEndV6uhAQ5
sKTGQHTr1hQL3L2uQy99MB3T1zANE/CHuqbTtPBQb7BHT8Ii5LGaLc4BU2/g0/kqJttDJmvUlcEg
9VycwVCNN+bvmyeYN503rOw4fi4fh12DZLHthFZFmt2YCjHnBtVeqECn7JHt2O03in2R5DWpUeqI
aUk/Q2Ky9NkBTPAwCD7FND6svl4fKECHN43lYLewsNqAmshkJtIBmtILCL0+OdlaZmfc9AbKIkqz
c3o5XF6sjij5c2oC0lLnP+hr4AbtdA3KkHCRQp+OmouX2NNtk/1Lye2ToGP71q7LQpSezbqlbSmD
/HQtjkK+LaaRHwZ0k5qG21wEwtMXr4Wpj5NAxeiPojAH1QpKi0yifuPtIDDlqiaZ3krg5K/E4tXO
IBO2xcO+oPXhRK3qnd63uYIMFiq4vz3z728sb8j55VZYJJUtphL5vucB35D0/qg+j70Mp6Vq4D3w
WTrX8FX0AO2AJlu1OvpnfZ6WiM/IjCvqU9HLTXL5GJfMVm46nffHrFdKZ7bl32Q0aexuHine/LuR
VVEx2NJQDN0bveNJRcmMY7O3F5lDUejPTuv0VzyhDyREu+R5Xs+YjzHJtx67ttWyfO/h1QlVN82F
tyhupKQSwKAyzYZEUGkPPue6Y61lCaKQquoO7TqDMRM+DIP6ENl2ryaiC+v4OIGVOHoSJ0OhWvoi
mOmjIS9YuNJH5Sgk+S7014QpCvqwU2vp+P83mgTroNwj3A5/lqhdnjDbsmdusScWvQy32M8JZumK
/879N7K0Yr46i8l6c4/N6ACr6hVq0RH49ny9M29Vfs/3hyQbjGdicSu/PdXlT0+9lKV0VQUG05vr
BCzQ4rEdNgGQdzH/V7eoWewcTovUHFGaJC8gS8YEVURuyrdcJQCR2FMd/PylgincDS2Qw7WvOHeY
ggMKNFSvgNesbaR6CGyEWSXoHloaiO+BZJpcoCUpkqzuCZXP0LsXiaFU2qf7OXL9ICeblGHbPwNY
vwoH2X5CPRIXm94GZ8hAbWOBRLw+Y9gI1pPGZPuWR9KXJF4r42A4AanywUL6Ze0eHdFXhjIw+UHd
VnJKm1iuf8Nx/bvA3zdQcVKRwcDFaNb6BgHtqGokB7PRARX1eULlzgaEoJrR2BgUKZu5MFpXIxDL
dUl2a3/VeS7jvtgCLYryCpSzrCJAFEtxfPQNN4O5y48ILWDauUF8MnD0IjlxhVKphZtjpECfHcmy
hGmLHxstM/rdedyT7G5cfxNwnYz1PdZXTn+prLJvwoqOfml3bJhcPmE5hSpuQlwRChlLVGaXRHkZ
Z3VF4S3Vh8oVbQWSWYlrry9axuaHmmmC3rK01JtJ4zYOueD3Gw8es33kJQGwa7YyzSBDAKsSEcdH
sj7Xr67M2Fbz22Fw9GVH7TxJ1wjvoQiiQOrJMRtJBYotfNQ+50hwmV0A3l/7zT1oz8NDajdtadFh
j6bHl+1OKx7KnzbFVTXI95zqbOgABIUCYzLjxrS7qSlSwq8rBYgP1j8LQq+XdwdA+84fT+7TUmH7
kZMKaSi3D2DxuIQ0G4V6wEtGRP8958PRtIrG3G5am4Hj2ztJdcxHyLErJBKoQ3MxvYqYzweMod+j
trrrJzycJrb28Q5hFZEr5uxKaE/83ut58qFJ6xJeXIAwjV9fJhdFT9B3QauVxWOBsM7ZbRAwwE0a
Q7XGqZWmr/afdmAnktdyeuMdMJZyPPoR6eXcL9g39Y+kZZDMoX1kbsRYawp3rB466zbDy3/UzwF/
UFZo0oD3aeTPrIi6lRoS1ABcWZRL0EowZD/ZiM00aMM7Uf+cfznxgjuaN1TCENCyEODGOtJAExuj
cjMrQPDRAwtwrIC0/SF7GiGVArm/NqhTO0Exv++CwQ9RioO4DNkPkrkrAFUup2mcQMX9+f2eAkIQ
zYQo42oX5Z+c730yTcpZEBqwAcRW6MDcR5D95NN/84YSbqpSfZxnZo5YOwhxc7Qr9U9aI6scePuL
c9ikxN+eTmRETurRKjKFG1Bb2crPxJyUPBm/PQlmRA4DsyNfiHPttgoLeHtwf99ibFTZw1foiHL4
xFfpLpaSOBW8cJa1vexTfeXP/36VgfVnLPUwk3AGSaR1FqfazF67k+bCC1gsATPZ3XlmnDJfrYZW
M/37n9+Kvb/7jHEDpv0Qvu+A1ZDDUzZuMqJK+LhKGmB9DNlxfEKGsCYyBJeHH1ZxU6BpeZPewxmL
H0eXY8+t2Ew4LIMtBQsPRWMi9pBiShb2I4x0bWd5I1aLgl4nv/udzA5zQPuqgCN8OhCVyALna+zT
glxP+D0aEqU1w5LZwWGBroqGSwa9bxV2j8BeXXKIQNjVoDpPM1kzEdNqrObKSI2s+L891Is6IJUl
anjLw03OFvTxKcbkp3X1ZLDzv6Lg7H4PNGsongKr0qd3NiBaJ7V31rLNSWcMoD9el1qEr0HFPn52
njwxTGu7Ej77E0cTpHjwSWE5gT6hharUVtcIe0DP58G5sWYl8GZWYoegfsNiDXoQ8558EwNEVgT8
jOpBbBiWxP2lHAyK4ZRJ5Q41maQx8scRsYXSGo+csj0xgHb6NoHSaOLSL/kMj/FEoOfgssl6YVe8
DE1/GHOOo9pMZIW2yRctEtMlIy3umztqZfOOJXmQyu1uEo7ovnHDxWTUQuCOwLVyToTtdGe4L3Fc
A7QZU1Ya4ibIYYVHgVqXg9Cux/rb9mA+RVTmg63AmEtPrt9zI3E6yipJkvjSpru8z0r5hJUDLB5H
v0mt00kUq/yh8lrvEVT5zDkhKBThfJjRemgdTtMkSXh6kmLmEsBmkg6Vjkn3GHzKHFoEcAw+/Rvn
n48oFvknwYck1qlXeScwNuVG2U/B/45/3JszNk7GBti7oggxD62pTQsPpjTgPBiyOzG8+jixVPco
NjmXGyiw68vYERQiB+Xyjg2gVfU8fU3ovuJDV+MAGAyre4ps6ospo9+OAATsfx/Q8qbQB0kWEhGU
Hsl33Ufq55ZupF9K3stHqR4emG7OdILz1wEYmh6S6EWMdbHnFb4+qvNC/E6OUnBD493m+ygyiv2E
TE0+NvyaA/djh0U+R6sMF3hcRT7YTcp3sl96beKz0GFEyUT0YWv3Yp/toQ2RUzXWqsIagGyPu7Ab
mVyht+BQ40l+9tQ6c+WXqIKuE3tvDJAOXTTVtX7O3jsGZAaJ0trXilSvhuO/CTvpbji3iVyWBp15
0gDg5Vw4x2jsSNkavz+eZxDHtFm8i5z+jJSEmD1YEsTQu9V9cRZHiSRgMkL0ywgWXHGsWhlktE5s
JNl+5ESucd7zmoUAFXfStZvgHSvdjAc9C+1TyXuuJmbpUONgfdQNYzA6mAvIGvw6JPFSTqEe4jVj
hyEF37MfVIEQGuQl/MP4AAdA/5vVxXXk9zzk4Yf708UPfwc3mzakV2q3NhT0qA8V0M6NZLT0nLhO
0+r0HihQC83uxqsgo2f0MbHV+Q8m08B+neLZ4Wudp+X6pSvTTl+DsfHJXOvGyh0WClnW9r3Z4n56
YXcbNQkOLp6DgVdIVhqCWDVtjI9uIM7KgmKPsiRP5MbMmw77+9gDdrjr3gj0yA95WPr5F9PiFAGF
nkfTiPLovb29JjiDv3sTEHDEZiph2SpsmczYYF4tOdfYOM966Wkgv6fOeE5hVLbNgc+cOqST0GLp
49eDaE75Asj9yeP5POKA2/FQXY3uksnggSNpckksthZzKitQN8JMpcucFCG8puVIvBgYIocDfm/t
EyYDb8te5FFPG0Svbh1JUZQXHPZTYnQFY+BMARhWqFD2+IeZJeyBN9D3atrQOsKz0/77LDoZCBYP
r43vGa4/zr43M6Wx5nYZA7NYuYj03PW7MhjBbz2+8kmH8UGNDeweEcyuRAndyfrAFgxP3ItSIWU/
mVDmeoqfhWcMYVnu4ZVe06tYIhQ2VEnkxpJ0VPT6x2u+ah7IFMuBRiIHHYdT/K92W5/vqndsZvIl
qs9KdkkPpzD6UeQV5By6erUnSbZGXuY6TRB4e/vIacwzbsEO3nxJabTgKmCPhv3z6IwNmcs/n4FN
Mb1K8xp7A9H0pejW13Wb0TCIk2VAkJJLIdfyVpf/B8Ane6Qg80A13DkkZlZBo1dznRP5n8uRJlG1
8OhcQg2A1uK3EL21fY1j+UtPk5i+e2q1YlEuhUrCWnEyO+oBMaSAW2/IswQyq4gRYTP2Sx7wCdiU
llBc9lsZHWkSNK9mqHQsxuo5RRelAo6x87qCtCQQlLwnf+YEFNihKHI/ZNDsru6S7VhvZtfKEykE
74Iz8tkt6whpgoxcWZ0KMgijXn5DjQsB/qYetjcN1GIJxFXuUzyImXBRz4UDDHuy7gavyeTeZOah
MfLJ7fLZm5AA8lGOQVdetg2Sc4onTSNZ32aQz7+AfKrmUX+y/o1iZqpPhej0iAakrwmH6wkpFvxY
eZWejfduV+JFfEBOVo6iw64WBTcZZBeGp8O+pErvvOOw9GqcQmQoPGT9yA1NriV3GYe+IpgIVOuX
2EaR2bZ9LQeOMOIoDPwka4DZ6RbecmdSGZaK8J6xaJeF4MADLkUR0B6yGpuh0bv954pPpXl9oLBh
2VNDBiX1T08Nu4wi6+C87JHzFjqfERY4D2clcYFBD+Ys4eto48KX4YNgqw8f+6Px/wYOzec3LWpi
h3kAZ2j5pYOqOGdXPPt5RH95bfeXYNSRqzjxO5e0jRYAcPua1g+CH69puM1PtAyoAb8SRQ28lhpc
JevNT63QWiknRyb+cVUjquWHUthk/e+hjWCoVrd58XXBROBAWA3aEz22SKoOYgb1k6UQT1evGCPj
Qy71sLFKFS/QqBv1n0laLfkQ8r3QQh0BKXZKJtWud2bk6yz0joizDq+RaovFUSyajaTqq9fJlXpd
V9K34SUZ8aue/yF5LzTimVzx0n/20yAx0cgz5oyNHPA/Sb8px4vQl8Te5Pm5PNWOvexR9CGSuE1K
mbwcDa2ElBPhch4LhrVe9XMn2h5b1tzivmZQS3AZ+ZGOprtnskks+WHmVhPV+YuKwxvwREnKxxiO
TbPbtDCiRX+qLFCIyZZoJsymTkkJ4OVGrgd9kjUoWYvwy1nwFpLpb6vOYfCKpmVkvRI3X9l31WAh
1CG+CFsk9uuNeMuOi3Jw9SmCQCI3pS3DRemxeDFEZl9ydsHq4gQr4JCZERfVQSmYWLKtH9/WGVA8
2wDOu788eUPQGmEXtJe0kVSPUI+bnFQMJhfOAKK/HGwraGAHdHC/HAWN81Mn+UkUARFAu215o6Tp
VgFuKafvLmsuTrxfwm5HJ3vfuzUHZZa8I/UvE9WqQufUyRcsx/gyiVy5yeX07rUmgLqLQA6aF6sU
Y+P5N+yBCwV/6Mc7mtpeQ0bbddo+piyTZvIWSHxU2M3p7VkTXsCqsEBz9aCEhsln2zL/4vvmsy+n
Gn51JEhvYHQlK9EssKPkdnUhG2BjlW0qyiyzoD3UnCfCQlBZe6RnhvsZ3HohOgelp7ki2x8ELcwV
0bMx7hAt5MfKEBaSXzNhSr+kJN7D1ai88pVDXPQ6ZOFA9P76mvKdXbIkLSjtHSJaeDMmhrdGc3RP
zKnSABW/feHmvtA2krBRguZYka6L4krU8koyGhQtoAW4ct41TxdQwoMufKFCpbebuiyGBUmshNM9
zlkaqNRxGs58n9X1g6XEWVnBK59FX7JKU7gdAvWgK/lh+S+ZhWo6ARBXJNICR/pgLyIzAuOWPdyh
l4ivgpT19oQQlm7OzCK3gxfgHnOdQVWrwN538tL25GoJDLKHyfLJM/iBPfQm7to44dp0QABOttcZ
Eg1tayC8vjgnplBYfsx2zaqRCZbpqcKo0ITHPYNzICgtWk5+wsigwaujameZVS8X/AhpbWeZbleG
Plory8LoEH/OMXXQu83q0rC5yBNp6kpohcUo/DeHC11uC227pO1nreOM+BT2Jp1ffoCjwsThFVPx
QI55mI1QG9bWMXk50mcXvpNnbCE9ZpcUOuq5dpzy3mwNukBV4ZcxG1B0XBrkJAKJl1lydTE7Kfse
BlZ8GZoA/Swv0aZqw9QWBNQW0HSouzImM7H5DTyMMMV30OXwfDtiuQ9K8Rp3OpQomo36s/YcabCF
XLU1tV0ma0PWh3P/OQbwRcEZoFLcSR7sFLvYoDggxVpQkTWMPdEGFE5EXFH2Ionb0VONq4JAVYKP
YOBH0HzReuWw1LvDZWI17sttMCLhs2QYd5yLUAcHIzSWbqhVd/JCUvk21S8NhGeQgT4HzO5CX4en
AGSSxGz5TwdUnXsajUYS43z+nJYXoH2zpEECy9H2dMrMc8prM1f+2xRiCKC6XOiAx+KSzoWxhuc0
keoTGvGRuOrPXR3ix3TclpYB8Z7ORj7UqxcKB5le+Sliqcy3OKQlDE00SzepAF2UxfH5C1889VcV
LzYB5miqGwiPxXOOuYonl1qEklBVG3qAqwc4LqOxZGHbha0SW4xZroEAJzDNK7DgQwfvekF59eRZ
fE8PLaP+zLGiVQEyRbZ/JYnyxXQdmT5hFu+WzSrNODg0Bvjs3GcfDOiNNQxnC2n2hu2Xe1SfH9t3
c3fS2GyHRR7xEBB5hu+RH64heeAnV1+AoRe2cOgitQUJVJQr6Ohh43JcuItZsFs6Cx+O9tZS8hMC
yNDRXvqlVSUUqr/JGEe36GMmo0Sm73IM4nSW9q79KD5caw6qft+Y+mb0kZfXn60ul93Dz8UqAjNX
luxu9XR7/9TgXAx91MSk14TkCNve29BQCKHhm/StKnqTBZY07D7Y1SmoVM2ncjVbuDxvVDtBwShS
9RoZ9ajD/BNYOHHi6bq6vSuzDaoszSQOVPyJ54l47G3+PsMDhIcOqYdifm9CW7xaN1c7eCXA46g7
PhcjQXXb/WgEsv2WF16SQqiP7NmS62pKbj5p4oAjHMHmsmXtGhUQTMMA0awMEveeUWdsg4Mun5Xg
j1LO5Xpz2SQggz08tQOORVhoob7ii2dpQQWYqTJH20GStsffVUSFEIBECGgPmXIEOLe/teRLyoQS
IntO0qWL4vzxgS4AbaGUXpgCc6EbjtjqQzwYpar0JEj8MGMfYKail5U8wv66jjpUMmva2BrWGsid
B2b8pNq9Z+3/QNIXlDMw8F+GC/lb7GgMG2Xq9bdGreijgpYEOk7A0iYATA9jINZ9vtp5zK9rPB7O
Sm/lCq0Ssi9ib33FenNgneYiwuYvhg5T+4RMZQ+QjeavGGXv2Vj51s+TnzO/ypF2RoHghGmGwlUW
Ltq1SJZBO0bzxUaXqOzRPnIDpwj3e6nVkChMjFy73EsomtVsbQRykRDE1C7mjDg0srilKLJZB9K9
ex7LgQCyBLvXGEBUd4WxdP9UAgEw6YfrgAufUxY8hdl5Tt1szMtNtekeorQUX58PMKyKQXG1/8hI
7AyuqwoBfSzBuCBaLoSiqbPQ9bnBEAu51pf5O+xlwwe3P12PsQp2gq0IU498GDfObTLHS7DSBGVA
nC46INxjJpx8iql487QaQ/pqsNjrRX5HwaWUS797Ww8MNY/w0rsuudBgCHZguAmUCuTGhYQSUh14
UcjFsukk1eru+C9qoLECA7p8TQBwdwL/O8ZicKoux1jHtGuHmm/zPX01KjmlCSmI/Wxh6fq3zo5F
n3QeUhJyUikzmQYG49yMF50pbh7l7LYi8V25YZpvhrLDfrE++xv4caVa/g7VEI4Zu5TdmDTHZXuo
1CCgkzCrHnKU2TaA1wZ3srQ44RmKgCZRSRo4noNRQK87IgqWM5ko4/zwsa7GAQx+25DPOrD0h+le
qekokmOs/sQRqrd9/hitov22N1qR4t843+A3by2Cc3B6U814v/JhRA1f9as3sLQpvCvpum74d9if
P15I4R1r3Yo3+1F25urMT6VrwTBgLj57S2BjjK+Q6thkKsRN4urOIN26XvSEH++henb9oIVhz9M7
Npls9dz6DGoSxW2/WUwiO/XEjs+apX0K19bK8wrvz1SkQ2oIjWewa9GF4kIpGMcMKx/Q47aBMame
/hAaogGa3TjApBz8Q3hCZAMY6sArAARi8gcOpblGWM+/5AL/GDnFVCwcm16we6re3i1fX3BDRb0W
Ko25jGhkF7aemA4FOG6izm39YElzsLH5vggN4qijyUF0hrAUV+jI3P4v1Cvl3lYIXooJW5lBnYVP
LzMMuDAK89mUk7TbGKoH6Nj5JvB2Sb14u1d26LseqrifYzT8Y+/Kz6mb280AqW1+PTsHMIUOPTgN
FV4eYj4BA0CYNtKCrBygf182xUrzcnAEwtpQa1H5W1LBo7pjGRjgbMhwY2vlG9GizLIyQGsC//wN
4ktBopAi1+MPhbgapVXKTqUy6mgxAz9mK4sLaMAk164+fZLFAx9Tq7HeeBDX6L9aDHdXdbszdS6J
V82tlfm7Z99HHqUFEmDFDfgDEK6X8xDa8NY4IZhc1jIEU48VJMnHSYqHY2FqG1g7TF8Vr3fA3Vv0
RoGocUnJrBpN4bNrB2roZhL1m2kz/LWBXR96FQeJFLQJxgD2VITEnrUwmhqadijvYY5bSoVky8ri
niaGJmnp7xldTl881l6s3LpdkoeopGgB5KrSd/eszpsE6nvm1trNL39je3Npcpfz1KR+gYHx0uWW
p/MEuyPzQicUziDzpHTv3tTkZIlwcnZYvBLccqgNAhdjV664KPwrkQznan0FTM4Q7VqrEbuKXVyF
MBrN23GZ8hGeII2PiDyeJYSBXKeLzEg3TBKEdkXPrjhFYrHGgad/aipU/dARwwPFUFohgOnSRpPR
DtZQ/EzebGjdepmReRg9f9jROmhmtNkMh58RD2hQFwb3j3Zxy1soQ2RvX5c4YZvvzV7q5NzXAo+1
v3w0WxNjvpJ1QvRxhhUAiDU1G18WW+mZ3JDD2qZZCusvnhL/+9MJvF8TkwBbnG63z1Ee+QHSYHKo
FWQw1MxafixGuctEKgCFODyvv210mGpvxKgyQuYR3jjfAqgQ0xjfrbQdNPBsR9hBD7+k66EydKNN
gAdZ0EBySAT0zS9xwgOFtvVF/6bUJNiuqdJj7VCfWx2gUaopVFoXHb0yEbUnMPAi0cqFN30QfROQ
pwC7vbcILeGfEJpWmDpMj06KnRFnQG5YBQTTwc8uF4Vut0D2G3iBFLMjMQc5K2WAEBWUosMwlBO7
UCPnwRLciRxQ7R9AsFYpfbcYfX4b5/J6HESboxU4YJwfezU9M8QpeZQCY/UddFuObAvgSWzx/W3W
iaepWfDUFVDhY8euAIv5keIcVDkT2pZnAJND9ZqJQh0yNW0bZvq9HkxjhjD3B3v3KBNHKosmYP2/
UUdkCvhtnVdiljt9yu1x87WBMe3IozTq59kWKSO87YSC+uRjm5F2xwsi6dUYFJ286qkwfmIlwDdI
iBHh/g7/+rYGcZMHDwzCJ+8UysIpInw5SfZdZ5Q3NW7ELmSs35bnbyJ+pEj4Klf0pPDlMYHShzE2
yZISon35CUh2kpZlE7uA7wAhDeqpCn0Fsm1X694ZTcBvNYy2Y6876kLpMCmJT9DAhKA80+QK5WFE
lgi6Gy8qLOIq4S1azwyLibhZOM+u3VusauzPW4ue9eXEUBORPTmSi/+nSN2teHGkYrwAasSVR5HP
GOsTpqMSqlr8kSbcZyrswmLCCw5lB/VsowaMd+Hp8FHHYrbTvyYsGgjiYIKvrw2ZGqbhNJtQauIk
Ra6T4GiZb2+c4ypLJk3hb1+0NTLqwNwdCH+AochoPbb+jrKa4JSU8NcSHJ/TMq7CIznnCQS015y/
BC57iUxtvlXeV5xZV3XXGdeJraeOP6U0KIA911Kgj9d0BD6Dkg2me1DZo/hYA6qG1+6uen8RNlZ2
V0wqe1YpX9ilsO2MyukL3+pr7zsb7vAqSWkMGwD4Qp0GKksZTi3W0px7BI34uCk1JKOjaUE5+hEs
Qq2LrBNyyxLtcoLlqA7vQa7mvULS2ZNj7xSEjp4LW1gu3OMbi5XtZYJx/s+BvQmQ/mXOrypzpKBq
bB+VhjdrPM+qzvYYHld/oHX8zGPO8uvnuDYoZMToPb++Kgs2YIz8P0LOt6/rp/0Gr3tx7cFgCR9V
9XFFoKotrIPN7wv+VZfeP7dTb0UQFT0Mj7HYGgsgpBn7L0uhcNeemqQXoAMMB2ljjS31RCmmbOXE
ghc8/Hc8Du7/KFa1xdI0pn3BvQ+KUF8znUrwJiNBhE3wA74KWp0X/IHUbSPIUH2IVJoHvHwHXf3U
lOBjxY7owOPQGY95j5oKFmt8GXzLyj9DYVYhntGAKjwlQQ9ObToMtUJycVG/P6aU5giBdWV8Hrx3
x61kBEbz1Fqe2ldFAXcmqboHzcuvIfTmWqwRK8UmaLGYprWfXW0cODt+JSK1UEFYhON94nOkpvu5
uREgCWSs7PXUhw9asNVWO1hhb+80AvMzSbLLL7376wJHsO/93lGsQT9ThJepKuX2yv/goRhZqKga
QXVS0cIzkwPCbO7lDF3d2HenGWC3VnsVzAza80XPYLIS1bMxyaaiAsYhzDtcnUg2iJpkdhK4XvS5
wjRi3yOgW+obl9axVwaU830IelKklpUSrWYXpNMYdbs5WA5mq2Z5HN4vpuLvfwUoaQTroF4wKwg0
t6p6Ri+Gp6yADlM0IOsx5nFEp05tS6auFe0JSsrJUI1i3B4vQlt991QPfMLL6juxHMnqU7UG4V50
FOaiEPyhlRGFPK13ySV5zTr4XzemrcJA9P+VmBqyit9r6rbS+kW5fpfRNhqUteeuIvbgqKR2V1Og
GX/yk5+Z/FcRNyqD6m6RvRWf/QOXhEQLAsMBvl4RS/p0W2UJRdCz06JdD9Ow8k3LyY3JucS2SHeS
woe4mwPuwBi+iyclpfRGVJ9SpTBM4HtBGF9CerzV5MifDMK1HyYgqQgg2vfpIZviX//KioNED+4U
05LV+EGM/Zj45UQYH7q2O3aF5XgNNzbOrnAIgxsy2DzLPtEDtgDDbJrtgaBjg4OQZjbadHQDE3UW
vBBi/sWWjdfH676mBjHWCLowoigSobv7LEiFddxqlfPgLU19scbTxmuV4uAUDKLdgxvS5PGdIxjg
k4A9PchJbQga07k5YDucD3u0bkzE94/vhDkAAvkOQdptVvTMW1erSzG4DaWmCnaWBIHq48ROFTPA
I63wopr51ymbW5YxspOQKz+pUhfMeLChPzwKVULP6y1LXtfe48H0F39YzST/ytTwrNjmMsxS4mUo
np4qUv9z6IUc7/Exz4rgtKkuHshWfPbGENh81oPdSTKmx4wX05Iu2Hbgbr5LzrDzlB9B1qmZQNMN
4QElf6ZGXqy9bM+YY9zBF3KQqv2rSmC9QLfKnuRHAisV583nr7PaWAhKFUTPcSNdT5eWHzwvkAXC
dH2efpTBM3HcEvwUHkiip0/4PjHzHfFS2Bf5roF7HE/aenrP+MGBSn7neKRUhwo4HqYlNn9A2xQf
q1SrmY6ibIiFDgiLQvdHZvNUe/PR8Ei5Q1nw1Xe+AX1jPzP7EAo6etaw5vLzjlxTLCgUgTPU5ObJ
U95L2SZgN4Mlz6KZD+ZaZiJJVc1esWonOJlcquz0eo/+Bpoi9fVm9+th3I2ve1f9g8H7EqSn6fx0
Tt435SmH59Qp561/vR5GzhSgMquY3wfaEnA5ACCZRyuuVBEU3s9M2jeCIRi6kqCw2VAXWIT/fOJF
6DQvxKEwlGyLS2FsU67iQXQpsZAaCDRYb0XKMy2mEr3Ev7PsQLegfWKpb/meKIEgiWWtIbvD9jGT
Z9Zo7/kE4JYE3JZOzCLLgjWRZBkWQhDf9LtEnkOPEh3qE2q00uPbGyd4G3GGdxE+7H1vRIf/D3ma
6pIZSUuRqFiADg3+1woLFUMmKlYhGD0w6I+ygcICJfnq8PCwYF1A9ECOs9FB5KY52E7/dw/w3ieS
gBcEd5keSRth/a2suIN9vxjTe+cBrYx9Ti/KQVmJjDNZ8JULiR2YQlXNKKZERINec5/jIfhGu90s
MGefKM/r/dT7aF+xymoNU11hlUU7aL+UMNVRu3GiIHJGDPn8kLkFkIu+HTrtKSo5qZcgTdCajKPq
jcmSZiaD9RIKvsTTUQ+CECOl40TU/igboZLVfdEck0MGh/ZaaX8+2uEvjlHP2/MP8CCZWNEjXS+/
mmw5T6K9g4oefwO3Ab6WtcCtboCclBPFld+CrDEV+3fBhpqa+JC877G8vLfuj9UrWpK0DyR/sbV1
pllDuBi6xz+MVNOEUPoUMHSFvxBQXgkOMz9iFyaSFf4lWn5YiC9beI0CH4zKqbsAqZqTR4afN1ck
7SqI9Xklm2aHWzK1ZCH444NZiPWFXrQ0nZ8DhxrRXkI/S7J2ypjTTBwTp0jMgenMrRmY2ou/JurA
3efumRWC8jWF787y0Jh1h3VSTfS6PbgPuivSGPsB4sWyyOWr1AzlNamctU5gSxgZfc55aB7xAEm+
QBLClHTMs66G8/OGPv+KRPA/zEzLoRRpGSeqAUf+a85MySAP65s2Ll0ek+HIvKt7htuwpRdoy46e
41ONH7v2lBRayikCZwk49uL0JcemRilKfyodWQA9qe0pqgXaLrnsb03IRnDPEEtVY6leoDm/fznE
1PF7tYFXDMKR87v/xnCVI/Lhag3O0/mb7kkT88E2VJ5BjVVRjIHQEj297SXbTKeiGtx7xc8UKv7y
d04Q8SL6es4RQDS6e1JjllDWffNBaGleDJEU4CUlUziL4tEUE2IsWlzdBkQsJy3X7oOAW7hI8Oq/
Dn793g44/KsgthvGse9p5XTPT+W1JrBXxqPBS85iyRmSLAw1Tsgv5q1dADrg0RxVeT3HwxyyFJHT
17I3kcF6PrrqVQi7TQ0ITAu2vaxxK4dEZP8pRqNTDzkfPVMe6hZZBYeMR3sDGP6vJKnJ/qcxumVM
eR6Ih5r8REgn0bYv6Ce4M9+UF32A+qi/GTGPwvo8B4aVgVtJeuvQRlMeltS3ljEG2ROEXlmBiqQ9
JlYCQpDI+dlDm7unpdW3C6R/CZhJUrNoMWJKFtxJxIk/8uvEBZjWOQGqa5sGY4s1zU/eNJgDW0F4
z/NyzBI6yE68eb90h43F7D2hn42grexHyuiGqnbyzK0GOR/pkZtEZSAIkW+gYJ5jmHAoLIP8POgN
xiVgbofngsgDaI2Xu/f64hr8wb0NDAZPxdT174WvMwmBcTk9PbKo/2SCPOkvbPTRNkrVu7OCZCTF
QpoT9Vd0Xiu0bSTbOtgplgbyskLjtvGJ6yeiNn+aukU23MQN9r/auFRo4bWswyKthnq3lKHYFhe5
vkAOx/7cDSPWTGad7Knd498LvhDD/wUMVkGHigb+Popw6NrgCNx5brxRVJP/7+Cs/Z2EF6gG0dNN
TVRuNzxtVOp2MYqOMrm6zUMsp0W40WCKL1usB0mcYdiRoFhOBJBp7sImozN1SyghcNE0k/xxHu2a
hVvzbUSqk2gNDedar++a2VrevuaeaevfHQza9kuvtg24R+siVpyRLDs4Z1VZMqFMs1OhzPJF7xkj
JPQ6xF+o7a68mCZ90hIxeEMPp4nrYoQWQM7YGDCUiEibdCIviMmF+V8kwR5qlhSyYrQ8kw+12daD
mr9kXXIYY7OL8zU84bR/RdNTkMfDHTquykMWMUGgNTQXhrP5ilH1aLrLwGL9/s0adUX5XXWc9Zi4
g3VTu8ah76FgcoBL5n86x26neAdAL0UeUSRXxXV7ImZ9ZXw5cyn+AJEJQTYC4QD5EB5LWOa4mUMZ
HSEn70tvU73MtMtGRNK7Lg+Cd7onsQVXsRfYRUhElLYa9tnJi+Zgtu5rJRg9nWRqEQ0LcETSkZbO
AWkIOp9lcFZs0uYMinYnUrKe1AP1wMT19mdDYolN9MV/sM/IjVV119+CRxdkyj92JAfTC0/kQvq4
l/n7paIiQtEgjDGjCtUnFZll3mmoluy/g8gmtR6AUzmHB+CEF/AxXKXFJLJLEE2NOcToVOLfHS63
cKchqSottoQjSWW6oTM5ieMOOURZ6Cd7JNox1dHQHBA7+ruHv5xNviXjW+qm3Xz4avZnfIXN3n4d
Tp7hQ1sRxH/de7p8wzv3b6tYnI00b8nCsL3AIqkOTVSs6+ECsYGMOIyDEwDw4SJILnjJQWwQ1X9G
lPg3I3bO2bM99IrpLaFcemwnbuZ6NwitUAtRFDPB7Pb9AJKEUAxNmMLeB8D0RQ3NXs1es4rxXJEB
pQo+hmQklucpyN+Q86DMafJARFH13QPgCE7kIz29vQK50dT6yCMqIRlr9pwlkMzkUUKHv71CDGas
eFg4h0nelRET6zoRGoo0t0Hz0VUM2P82NJ6OlkjmQ4FOSD89z0R4oQP9LzcSAJ5MuPkXmkMktzK5
PCYIwXjm1brl5OL7k2e3FBGgZQY+ocQTVDhTX3kIKHiV4+SDuNHyW+xK6LjEOmObFi3tr84FJrwn
Bf+cssr2FF1hoMrGxov4oljJ9lYX87J0DLG39J9QmkvZaNnnqBd5zRHuDOkkn7qUknR2d/4w7Far
PqrbdDN96BYDhibAP+LMmm6nhEzSjcIr9yQI7kIglBG778mT4QCEcsVYs+cg3v+56DFSygmbohF4
2b/mHts8D78FBT0jq+o0NpWfdGywmEYdy/gDQ6MbQKwUBk25ZrTjdLxz62YaqSqbEr9X2zW0lvhL
Rb9RUDnJgoKkwznXxPg4BNAg13pd3E5gmJ6/DblW5dlQ6CEWMQ4zXaRkpf/rtdMf2x7xai2qDCVM
G+Z/BuJDFxvblStchhLremYNSt/Gz8fy2oP/qDS2LE2gjU/N2/INeXHe1jxqplgnJrMoNdAKqrOZ
btUVGhEi8SIfHYRA0bxP5t5rSuh6X3niM/Xt9+ukE+yVJsdy/KatW9ocaj6IeybAxV8xDvx8iANh
b88YrnnQNZbbeHOdKhzpXQGc//QzgVU52gFgYtHk9sfjB8dWu+umgN8B9ufOL67VOLMHdnw+ZKrI
rJmqFzzlD9qoXaBDZX3LMPdInoRknkc7pyLsueJZcCpYBqA/yWW1mFk65o9IRnhR1ABO5mUE1ZxW
Gk3iqcdlfZg8JLr6LHyS/kal9aQLS+0CmVtxWMW1YcEciyS7kuxn4ILtq5x9baHFLyFJcRj3m7rc
A+DnsWTnb6I8OsWteJWPk5Ypoio2SOZsFRCt00WMzS/q83iIaT1qwVSvOzwEG+vRdJKO+lUSahP6
ugsZ4MiED+3MNXovVBkaLlfd8SrhrRwd2bFqgRVtUOC/l9qmvccaDWJ0qOVLQ7UBZxxA/uKiwGZ2
v2NeRWc+kLUcTP/nMr408PYVJvz26v7BPMPYwjVSZA+AfazUElp/LGndIYFI7QlVWnjpsriRUNjZ
e+S4qy30HX3TOzSr8NyX9W8KyExrJBCP1Cx2/KDnm9h3Fj5z23CrqEL6UXgks7ttvNUah1Gt/Dx0
hIDEhUKeeJAsV13CoWGE8cxTKnViDdE8fZ5lbcMw/Lv8E9YSmnVGqkZSaBT1R2vN4RaB1kE/rgK3
HI/00ostc3tM0rruSErKPrH3fALkljSGRsBJeRAGUjDbv+bybS9DxDSCcvgvNP5m2xx+374MFblC
8rVEg1Mi4bj/mYk4kycTblWxPwh1YcrI0MyU7THZIZ1JX/KF3L3UtS/+qBakfPLotqKvBwIic/du
D+gkn3xL9Le8VOgAsHpsaf8dz510FDOD9M0t16Dxhg0L6eT6is0eKSz774FiLPwUY0eDDWlp9vFv
4+dbkB1u/QuGATrZzSnxreIY/HeamEPxs+BztegZWmvysWFZSGonGhdiSoC41+oHysj/Nc1R15L5
EiJ6ApvjHnOj+T1H2l+oghNY1vqcrbPLVErtanD1wXDVNP4KOQsecdRtwIuTMEA6FXyXHY9Se2WE
+nWDhJr42+PX9qHxlSK4tzDKvbEjuAUuXz2dMTKytri/NY2l3F7412DP1U/Us2lqs+BrD9Oo38te
Rcucm9YBOl3TIhOYu+bgMMJ+pmdpJ5OUOun/Gd8Pecz30lfKfG8+G7ateF6DXvwMtVb5vw5+sWsj
H4uDDsUQ6Nk4S4CUIqX43yGNOPH8yTA01W7jK8U4UHFjuX3PDCNnGvm28CG9DYxayDUwVxopOVUZ
TgtLcBRuRIVfIjram9tMVPphdbVQEnqQjgdTZx8fNOtKcT5w9/1aB4yqVh7rjeTpYqY52vHPwoD2
E+nfCMbzArs76I1RduXzawwBjtZYcdDOiYBvsBOynPIMqNcG0vv/FPrKvlxFyZZDyCcZwkXFDvcv
YcCnpk7z6tu6JqI4xHVbNG0ze8LjO2jB9rNLHMl8o97Gh8cCVpopT/bvN1ILMVV8K4PbenSTzfHG
lJm+fRPIDrZxf3Byh7N/tiAxctGHpz9aetV85X9HbYvsPibXV/AP1Yil40DcnJ3JEDykwdNb9cEO
SKKdiM8/dJFHn6PwpiynKUrSoEI6bJgivgfzRfpUkn/MMwMiphZOHrHHNVDwhrd9Qv/qwKMCXhx/
DmAYAGpXRo4MW9M/8B7Z7/DRzegWTR0tw2YXuTWEeTqcnDYwAAGLrPxmY3kJrFKvwmAlEjBInjjL
QfnxmmFbDZJ4M51aBi0sEDY12ZCQIwsfQB36fWPtu9AfHJ2tsahsnzKpe7UjgdMsHfGpJyFirViJ
lxa3D3DI/7tqCcLNZ65JMSN2DEpCSFhoMQcfgwrxvzdotd+r9ls5AoHQD2ofKACQHKxzYlVdjPPK
lj1I2qZRkYoD+W/+7fTKzaDr+IE4Q0QSOfMhIj3phA7EzFzq/SpyV5m4uTi/HTL80q9UJYm3cjVN
j2tUkuLLo2YGXe8iXJi8rdwNeMV3Cn/Lm0RsAluwUuyEofdD9i62IRPidIzLwnwTAw5qXU3KnhAZ
4KonEVsp2RGkJ3plVnY+WDJxpbwTsIwMzXo0x65UhUGSmCOVmbzBf4Wy2enUtpYQIf13OFmfe7jx
SUiDnHUi2FFab2S1r0092ZgCOSEwiafEEt5a7GOHLIG5kr5Uex1ltK7Pg4bjkOJJv7OY/P65wbMh
8EkZp0y9ldwYgj7LgZI2gY37XBPJ5870H6UOQ66wvrDYKqNE+y6GZtzLSSdkoEtSZtjgaFjvMuaJ
URw1lBYxTNfwZmdldzpUEGZtq438+eUagNoNUFpJiKneBDtTNT0h7RaRDQwqRBK0Cd3ePl/ksi1W
GQaaOehVVQMmbY+a9nvZ0CbC3fbJ30tq65NTVBuXV43xAIbx0KBzJLmeYJPOgKqzL3QB7LVIRfG7
va1INRCPXAgvcaBWfFm6SvwPvDF14RFyPPhH12Bu9s9Gmc1HcUmWUFH8FkRf/pX70mor85JyXaQM
aR3l+b4EsuCv3fxaSL7i/5Uu3XFIAZLsG1xzaU2X+2RPOXLvj4b9L+THP7ebPUtYpzY0U9/KOccP
dDeVyxcvUeURAi0V6z1Uy6kwgqRlPJrCqPa2DbmZumh+PoOxS+1wf2Z31XnaiA0d2j8iSvCbCsPt
M1qVPHPhml25lWCIPDjoJdbF09IuTh8q3LWLcd/pnYGL6zQI1GXTA5LIEwytWLDVhJb2bL8wVW8a
EvPAibA81ysK1d2P96pcyStv11udrL3AeNjH6DzeYjtXVdTasGSm20E4MtxJMah7ose7gsJ+QA9i
QAPblc6qlGu6HwjSO0RoWfJ4HbYuNU83SRC9Lapn5JkfWWyGT6NmDk1S1FJn98A6JK2gGsyy+Ugv
T5D+xjl2LwjEDaekMFZXezBssHZeVzgPLplJd86HnCcfw6SeHLLomUvAlBXno4PIZz1qUhKhQnPY
GocnNM3+AS1V6z2yh5txSC08Mcb7S9GotXQG4EkaE+eEmUN5U16zR6vynV+jk50jIrnn8UWv6oiv
JrU0gvs04y4tmx+/2jpIJDYxa0GMHImR9YJ6cmIxBd6mFMRju9cj5IcqN7oMRn6lxcIPaHh4XPmv
eTj2nr43BGItg82WR+hCQncIJvguPE59EN0TomoZVx9aUiFI7dDrlRe12UH4Pi1WZi22oWDA04BJ
r1HwnR3HVu9iIRky5KR/wDBTG0bHgwg5Ly9PRDIaQWDKDHENGp1BWyhsDWItfQzvVhWQVHU5D/RK
LlY0+WmjN0zrJa/MQDMiX/enslyPaxvLt+jwHAe8PW5guzMVvPydW7rJBa8K1j/4Ge9d0kRQC2JR
JaJCRZXy9u8+62Ym9mqN0qrQNj7gF6VL+ejsbg/FUmo5N2wHewedNeLP2My9DBuCBMX2b0JQwoYl
MgHjRivDF2wpiU8FyZr2tDR3Hbr+K9Eb8m7MOWS1OJrqX2TI2pi4B7Jw1evnTc555Frxq57RuOFq
sQtiW8GCatpOLOz7ElSOuYBKG4ISbWavEiNz8GUKKUpMTxZzDJw+WhlbARyVqj3bRZCSv6+kFxsO
WDFYUuhHsfJkEb61glkVA4IC1YYhCtuzhKZZp2oq6e9T4vH1sRwFgPgfcJCfMvHE3GE0fhLi1Gkq
T2ghvgCd1LzuvnT4BlPJyviLN2oXvUlUOZzGbc820ivLBD71fY45wKtnZXZUi/athAhtkjuuWfGM
zqWGGOWZfImIUVkTeSXmMKy+PmbpVTC6Ik2NNRO5AAy48vTSaIH/0iptvyRzLkrw04HfSgld/WTc
ACuZB/RhFOev86tF3e2aUUpGAahFDcsC1ZVU/seXB9tmEPeyrseEMPFRS5BxRf638UooSkOWqcp7
hvdD9QQPp007j2de2o127CCubJiDOAGc+N5TocpDGrWhAIavKkZKvrqYjO6CbvWTcLQSNRKNCmpu
E7nOKjdCoaj+9VMlPdW9qgT1+pXyphwI0k6fdvApUN7Tb9KkTJy9Io8vqpzQWb/4zHy6zG7zv8qq
N/cnI9dCQMSMqzj5wq0Q+RsGDCwoEdoozAGElzyn6FsSiSOXvQwKQkKUkS7BrZo8qCcgPPRccHcJ
vm4+AixFohKOQT2AFaEgylErrSmnp7wkCeAEQk+dR7cFPZ71n6kzfl4c0ZRgpNPZZ++VWj3oGbpa
y2BXG+4q70xZMuR5CqMjuGQ7XumR1NvTHrNALmKmzQFCu4BJlAisazeKF8jMgcfDJC7QFigu43gs
I73NNwIVmqI5biVZgvC3OQg5vFoR2Xsh5gd+H/os/GeVmuwVHaK4kupHb/4SkZ8wfWWeLDbjtoBn
ULGnlKoITij0SQlu/3y7ZOENl6PGuQzX1L62h2y06oZuHz72lvNNCE9mtbemvazn2cY4X0Rsgwrm
jo3Z0z5+ETXokD5ydTObbEfF/M85pRFrvg4HytTeJy8X6vS5l3zmHAna/w2ORviGyES+Y4wMSHPr
YEAUDV6xHHIJwfIj1DpX/dzUBUVLL9mLleqbeICpgfvH/iP6jInJa6/1tUU5jHCxfXOEJqe9vLpj
/4odNtjMKeKk1AlxHAHFmau53h73Um6eTBZ6crkloC1bW4Pp/wx3cnD2bG5GHtdJpiJcoHQ52II9
gTUkftnll1eSMgj31afTDLut+iZBMhhGvco3Kqe2FBk+sk+nIGbWK5J2lmM7N+84nZafc65dlAId
r+iPHP5Go+t0Nk+rkjoQNbfEg7e2DULQUz7eJlZvhxOtnhnxN1LepxExLIrzGTbPY+GC4+2gSslj
Nv3UrTpWWFtx/okE2t8YDkTcWKQtI4/yCxa/cNejhEIOgvCycFN96kkLvSRS+HTJ87WRGhVXblmT
HmA490+vSZDuKBgIfO9qJyTDctq+xEjtJ98IQO8aIhkO00XA0txJ7K1LmxLsEPb9mmpHC+Cq87Og
0Bl2plPG3qcB2/oAw87otpV7ol95ix6ffYweRtBGkhSMnf8fIIAc5lZ0V+EGXVhvht7fQ+0mT3Hd
vdcRbwTts+V8dH+a3Hfxi24emvdMRRKMywlmyJpQf36sO/xFOal9ctFDNhsJXlPZxNuDc/RRUU0k
LiSQuqy1WY19FOSBHJK6XowTzd/IN/lIcERJk1n0xh5t+n305V7ZzJHiv2VOSNdBiu46XpK0w/rO
bsWN0F76IF9KvpSQmu3XsgVk2P00iLt06xrWtFRH4Hmtk9+PCRelkEF75a6defuvzb4HxNSewgl6
CG+rqZCrlwgTQXFabaqk71ykfsvhcCgsU2Lt1Suc4ZBFd52jPB+AeO++AVUIkm1h8Mzm4NmUvW4m
ElOhD7DaZAA+KJE+z4lv3WpfMhelFMSV8lSZ8xaIaosQimcKHmZc3tV+2pz+5eH2pJPk32j6W2Mt
jGUff8NvmMIvndBzn+B/Lzxi6qgHU16jSFhy8X/6zUrtofcG4Fw74lO1EvhYivRbWn91qrSY0snx
JXMmV/ndLoXeJ1zht2lis6sbPo27e6Kn3+QwNc40UrNngVjjjI+mhB+mc3mvAZVJih+2moSvvO8p
xs931OvW27uniLzgrcBfKQrGMTlcOY5OxzJ3InDo0RBgWFFMQbXBKxfwJ7iJh8o9jB2ssDuZFKrg
ptRpvL3VoffAmlwmmWlH/RgH4Es3jigqSVyKob1mAROWWGMcNwqQfDXb2TSNcrTF1hB+o9NMjUBb
hBIq5Q4TO/uIj9RdUE1R47bWqNnMBP2tALl5rCPVYeeOtNmL9YzmmbJFOXY19nYFY8ZLFXya1vXr
mjSKgkE3VH7ZnZ9w1Pq9UoUWFjVSKX0/ff0kpOJX8pQS+eJjB3KENUet+YPzApWrCN1kpmklPRBQ
28DUPT6aKHHOy7tP2C7eGTFLktCXTTOkqjtlVDl53R0jelCYMjHvHeLqgHSnvVRLhVtB+j+yUve1
Btapd7RgavljU5nloblQQINvNEgC/x1KPohtXMQbnR9eJSqjwSxgPyeH2uEFovYMB7SViTcX3Lu6
wfPE3NZf2oEn0uCBDr3jQHRvGYRwWM5zuJKD76iNwh4wrxpXu1YW2mwzxHgS9nhNFPI0vBBZK8S3
yoJAGMuHWLT1pJXFl1MEKCJi1Fm8WPQi0+tpzHlkguJ/WQg3SvTV+GxIcjZjhJ6tcGjAjZ85Pp86
KDfKHm5KyAEBv22mwgPufdseFIrL8DGCKGY9vljw8gf4o3J7Htk0mYPROR61UrxfNb4YPzniqjlw
bTN62RV1GzGQJH0eafMMTacLpRqxp2jLkcQMGhVZbIjwIcnIEJLUudjdC8f1FEBJkU8YJ2JjAAm2
h8oXTzS+1fD0cTA5imhfqwBojfRNnFkZaCSemJfM7GCzi03JqrTIE66+yj6CETXorzcn5LpgZOnn
Hu57KGUs7leAeXR5Pjd6Dt3Q2yt3skRnXZcwHgZpcADlWJieHfwRezr5K5hfITS66q9OCgUOgaFY
tf2O287BN2p1Y7zFUBiIQJrR3SO/iTOi6cNuFOJYi/6xX6fp+60YBuLSeCa38U0go92RCjpiiQlE
TLOVFtOHt+BSp+i0dO20Y7M1R54bJJcLrZwZfEHO6whcFlct0JEfE45V7Ys7ZVJAtikL4n5YCc67
HomFEm/IKcd/5frYherdF+aWf2IUtTC60Uzxz1YJgYqStjDZZjwz2XNJg2Pkx187ITmbYuaPkIVH
dJd6FN3X919yhf+rkwuItdd3H7sKl9SZdv9mICQpZEse+juGJ+BtEBFQJWICxtQEAIjsR/vICxnR
jz61tIJPbt4IaQZLMCstL5xnxfgud1n7N/vIc1TUOWZvvEcD6q2LvXk/o/ikOXIPNpgJYFB8kffv
Q5/piaDaxwQupiugFK9szYh6O3sy3xROJ2HTLK91Rbof7+DID5Ve01bQYTrAnfbxq2oKyA2dzug+
23yE1tcYMAVvhS8vRQD38waFExXdenM/3Cu+fna5m6IEymrgwOVhf4igu+wVY9Tr+WFrwcsv5pQU
5UELhYJuzE8z2HEw0AYuGkmVs89oTRonxrMxqNw5c8uxRp7dQrz6h3gqElq6o42i4RnK1PBeTO1j
hap9t5x10Usk8OGhm0vvqsgvT8GjeC/JVvSxfJ3/oshGUWlWUC33ruKeQe1msBEp7++90juTYsR2
pjovHfs5M65aFBxyqfeX3fpW84ZgYXsqitmoYyomPAAa0hCnqauHDq+DleKtC4mQ3Mf7ge4Wtm7+
TW+c4TUJp694m8/TItAiGdqXoI296ZhqPb2FbVytjB6gWJjCJ+VisXtsgxtSWCQnO+dscgYmk0Bu
0NEJoixqi81+oURQROF9jJ8qfqbQOO1Ot5DzcIhhxJysdm5Z4/gz8Fucj2K6diUJRFDAGNwvPA89
I9pu59E1cMmH+YqJFNJzQJjelIt0L5b2sFCaK9lwfJlp3RAXph+pcuCyGO9SrwCgKR5STJjpX2tA
h4qJZ3XMXgupqtajtYVt1CRL+aHb6tQg8BPPF+/QkP4wqK3yvUPaFtEffXyO1pvQofnMQo6HCwZ7
QucduMol3H23RfEKwZaPekLEb5uo2OTripURRDzLOb7lwKZcay8sHZq37ZaACaOhLyl4CYxaaBSp
PBefAw1jLL5+OUp7iDvrpe7epyPmJtynAVE2vXa3wHVRsRkNDDDJH8QMRj9W6xvYyJkwe2eB0jgw
wpEOyko+KbIphgleeG3JHcDdSMyxUF63pf5pmnwQp8VhlELHqkzRLYQHIvqq/FZe1krYoTgm3MC0
zbRkpAtNI1vbeYTeSUq7ukJagKC6OmLYmosa1d2QK0auZV9ul001KBzLUKss0sunqEPBAzGHVibU
lUbeL6pJm+mccgYpuVdQHsDV3Sw0RU+ADxZlFmg9RknKkdPz1ZG+/S/jF964YzVyDOqHIgtqEYva
DXfifzgAsuOSjhEvSeydVTimBZivnxgtbnRBuAB0cyzEOjuuj9KEjxLn2ne3JSWH7YWQi1DhMYls
3xwXWMyXXBUbhMa9PubBF9VWBeWHm5Iv6B7pthQsELGyxd7JBDH2uAaodPPHyQm1OOcbTKmBO0yP
yrvajzloL1AlSLEbcxVj9qIkd4YY2CHqEVY1kntpFc6Su9R1v2cHIfDq8Qhj6dWG5TKGqFbZ4aeP
fm87cETdGT11qxf7RHvnL4oTgcuxXYtKPZmYvIwsS476Ykg1T2SkiZepSYPTk/kn95gkbjxvwRgn
/gVX0WVMz1bwfE4rIpVP+/lp1rXkNfpxgHmZf6UTjEQsGwf6mLutIUOPP7G3AVv3Xyx0zFdT57ZM
G/bxvM3I1Gwc31aNrS6cxx6iUVe0rNSDT9mgX0sJblSTHDE1nDer0Op+SZNvHKpqF8U4aS+8F1kH
xHW+7YnBMyBihzfT62iSnOoxKX2qQ1AZ7I6vnYfmG0cwuNcPhbDBm5EwWxPHf/oBKeMnvgXCeRQA
e499wqPxvS6WcHKno/q+WFKTH2jSGiT93TKBXm/1GMr+p0TVCBlxi5YvI/c9/V7tuIwAxtP4sJLj
jQDMiVWj8NGk8nHwEkwE/jnh5Ge4ZLS8SRy6xJETJB+Nig4HyoZcCm5R+T1VaT5zjTw9mu3G3eJa
7ICo9CC9YtzfedKgwx8UNz/D0zzL6l5TLuKtDRPfxw6qG5K8euDH7+LfWQf2Pt1hpk01gKp2YWy7
4G4s/JGpjyf8ajB/vtvExTe7OUhkDPaKOBKYj6oHtD9FDsNCrAxmyWVahM4/1jmuNl4fr7/HWpqi
T4G6VoldSnu5eMpFDlBitbvteSv0Xs6lsIL0OfgiezuzhDsTov30Cc4D+slL5/bwREGcbXKVqrHA
I36p1rzHGwLiQ6G7CNXiVVzOs/s5wtsqupgr1SYXEUm8qHL3Y+HEAzgZ01t7HqOFNLxcwkpqlsPH
reWwcDwo9c7yMhwPqFSOFoxYtWocacG9ZxNPvZcISTeCRZkOSMWqu2a8dlTW0yO1LDHiR9WTK2Sc
sUjSkK1GL2OeldALhrI90kQmPokjECcPyf6JspF50vn1CWu1Nm47ZeW7V4ynqCGJovm/vAet96EM
GiLqoN5kgwts5pW3GmNXoxq1dABNDB/s/lsForThPeO8mA5IURXq50F8ynBrVHRNPxXJScr/6beU
waOqoMB2CqO53R6HML1OFo9kRjrwojLDUmobPMIbrS+2Ns8oOwuquN7z18ObDsSDOCxLygfS8/WF
FflqrLHGba0KuNbxP4dEy+wHV1NggoZC1B6NxrEhYfpDRlmy8WPz9JL+H3Ku3ta5nrm0xe5+fT9q
80gY2OFuxJuB5if5Fl5fBLdZ29/8Baj++yDom1/zlYuTeN8NXo6WBc+GMa4i51DsFjuzz2+BZ+2O
Nn+OKFFh8/RiePxw2OBWdhvS9lH0WkSTEV8L9SI5dZoLxGSySQPVpczW1wn04hU2fXf6sM+/a9nk
L5o9E/IpimQRyUPYlkosvtYeG4zdjxXds0VTWkoCnAzy/vsBfuDW7YGeKIT0gmjZA8mMZC3sJYyI
F3wgYr1QpxDDl/q4cz8ZI/qI9K5PrLqQINqwOkB4F8N/LhuJLlk5vq1PHSc5TPZYbtLuhMsTF0Br
dQRSwfFJVg4fYdpdayd+CtMqorKnE9GAsM1myNXkg+r9oIjPK3XUS2e19UfNlZjZIKS+Oshh4h+5
gUSRnQIVY5OroJMGRkocZrYDJXTyjdGTt4joqs8cEZdbPBQpzAeecV/Ne6Dmbfr1nTnf7lAA8uPF
0nM1q/uOj/2yHdjMgh+tWMpgQEBwZfXyoyOXov51XPfgiQ24VBu6GxCG2b9DD4BXudjzvxlmH7Bn
QXMqYV5NhUd+4fEkxK28LWiaMRSloHzXqDy7pz8fTr2a3G1zeSv5pw0IIasCdsXN/8kF2PW8PZLj
dAfsXEZ+9j7nKYkO39nKv/QMBhzrv5sDXQqnGwa4UIencb7Hk0giur0EHtzZstaTwMwD2j89jnnN
u11XDqPZ++6JvcvRzChJXFAGSi6Yd4NJsf85OzJi4+0qNZuNsJFZZkfUZsMdyHQ45JNOvSWxFsgm
r6vvoLwCfXhEWgp8tyh1vDgdGPxWca9Vmyd2JntZ24/Mzk1KQ//DgqkoQBzQPNEJEODWuUlcp6pd
+Wvt0znvNzzmXvh6W7FS/MBQGTETaCTrrzCRdMYKt0htOnOdZBY2MYcDAI6UGdTifS2q+dUGCAYg
WHX3x/AUujwAp8+FELDdp9S3lPtgV2PypMknZ7MAbSOnXKz6SwE7rIG4vCZHre92LOZmRbXZdSrJ
0QyMe2Po4ATrT5DWaTAFjCWiMWjZDjV66UShwXVWXNOzht8nC5lMMaZhxBqsLjYIv45w3O6EWa2L
CVpFnou/jpw4dBtJxEAdLbIp0NYBp2QedqPbiEoU6DraqxL/zTcgCXMHAAQg+QWhzWiI+TciIUKM
NU5xkcAlAQyas8Q79/dtyAGGKZi+Pjr6QW/0M619c8lED4XbDRb+Me/xxreKgmkYGC+2VrjfhADh
kqQ9r4oLhVkh2jnXbrdifSASaFRqcTghQTIxt9Hn5gcEMXhGX+x5ajJFaH6rD1ZEJE4Wvl738Ppy
Y7NqdJ3Bc9vx1PylIJRcYY24J58jlh1BfwAmhFIFeLq0HL5LA9Stg6IeV7QcVV2b2TdRR3PgA5z0
8VMubDRUUs8H340GI6xm6mKCumo3SLmbLaZbwWdHcb0ER665UevfHB+ge013eVy0vKktpiJg637E
+hy27Sp0MWDcvxs1kNH4QQ64PbsUJIUDF3I4PvvjhsDHH5OQZ9zaMjHsBwL9aFyBgD79tLo5kmyL
Mi3hwD5dn2zel3nEznTyJzWVL9EDpA8BLuw4N/CUZNSmP1enT08uC6izA+xb7McEmejgXPWYETDl
HytCMg572ITzRv2NGQhqmuApgDz9G6N4tpl74s4X9jW4N7ssVeu50pJc/OD5cvG4H9Q/GcGJ1GGg
rAfBxxxSMj7MNaxVBrVWPx90JcmDySUy1ztmtgvEVYwzIWfrVD4ZcmWIzDZzKhFoyMJqzQIr8Olu
wHcZRsZSSqItMUNHY5YFwY0EmeuvREg/WPabv8hBgWo4oV5b5P8dtWqyea1UL5zxOLRWnHuzV7PG
wDhfIfLMfbGmTypKhijMkyxf9jSoGemA8NDHdHmTv+buWTPJwO8m56AwWrxfeXLYtNgybkvlFla7
iFMstY6ktp5NrpCssXO7R7KUuSTz++ybpw85XBTWU2HMHvnvDCw7hD49CHwWVnR0kDhwCZ75nAk/
G+GUVmypSJgm93X8HutAhrNP/42TElC/Zpj7NYBVObgmwPU1mBc7mE/Rt1GC8D5dl+MQ0BpTEqBx
bATkA4egWeyMZNJcOY3GdtrrZgahvrbNex4h3WPjccw3+3gOhfSGxP/HbutuCQsBO6YIgeciYERf
GagrMoUHY6XSBWyW6zFTSPxowWGLZwI0ax6sGP/m8MX/e+DiTUqCS4cPAhoof9HUREL9+ew6eJni
Evz3UL0chjjeATGqLTm/aZ+qeICT7/9KZldJgH5reiBP+Zll5PDTZr9hww1Uw0kOitn+DhJSfAwA
m2NswF/6FvS9sq/V1r62XDp6J/SZJ57k3aBMh8UwMLM9SZlNkPSzOcdX51iw81tPc7JX6m4LzVHm
k3UXgCSyGr/RpnO2BjQHfhIgmkQTOcRSWcjgEzODKvwMlajNrzb8bbUMXOzIhrYGgGe4IJGTryNo
3sMYPmvG8JUYve1w4Am/4DRDiERVGDsEOOP8k+lK+vgLOzqkUNQfSx46zjtpmP2lelc3FTj6EJE7
FfDhoSrdYObr9gyXoMKIv06pPll2XZLu9niwjfWt8OYSN7bOp4U+D55zqVh33F6GPhCYugOlzKg9
idm6RDkzbFlwmk3g6BFE90euXIVNUOm85Tz6HYYvzgTxyiEPpq/3eLqxR7XJhcsVCnesGzInb238
oleJThJ5H0Oeb2uSSJLt/vXGyfYEr17peKc+3NDF7vq6eB0/zYhKfkwol0LxtU7WPcrb0iuoqf0k
AOQv8mz3WV/FrZi8X6vWxj9cInk4N807subM1sXGWccxiPWqg3PeDykjKYcvLMoolbrub7rSZrZw
j6J771okNTKvDGUsm+5er+QX/noWqkpJlNMYZFEGedhfjY0pKPVxi+kj+CtCPG+xUDRFS9ZrLxM3
vJCQCknqSZ4SCgG3gwJgPAwKVZjmtkjphyaV2riZL7mPZYr7DODeoV4LukcWi8zk3NEwLiJbz96T
LQUTJXDM+lu9qHwSU3eOWvFugpfC0WXmv/V9eWTiID0/NfFoK7WO4U8iaMUCS+YZw6DA+ssRvlSu
hT50Hj4k3fdYMARdG1IPkgSFfx0hnAF5y6zkfe8FUe0R5vgjEtja/U7Uu6hFaaXVSDHi2Ip509lp
2FGKlXancQMqAtGBOxoTHfPzbuvmDrHV3NjX8xlCouTsn0YyXbhnIel68TgnMaJj9ZsYronW+y2s
JTBszTvxdOr/SJPewO4tMISMfdkVGk3FD52YSiEnBa6LhVgWzm7mkSFOGhdX6LQHzvHTxp08YeEN
gUZa+8shBXaXBWDMFy2wZUppBya/gdd/WsETj+LxwhKOFOPkFB75TmDmgiYDOHhS9iKuz+0FREp4
iwW3PA9QyWg3pNj+VpigunSJW/XzZGMGG31/1BB8jvtIYCXXDf8vZLPV1p70NymAM32Q1NtfFTZV
oM1htNgtt22JvIeyeJA3Nwzfl1RaWBUhqvYlyNSfXSdxY5e+mX6e9laEoR2RC/yWn9tn3AOtZtTy
t+eHp5FiOA313JiQ/8V931FFJbHpOb1NlU+A2QnMaTZnpYtZQhaDG1uNGN736cYL9Ay90TLlcv9P
U79FtyStq1nMAvdD40ZW+8yFqCbvpcd8SPN0Ut+ZGkv7PFYaGytOkb+LADop3tQcs2YoltoKLPRI
hBVRJ7AkMwBIa4gQgUzj5BM3dLHNo0zY4ExXkECnlZvfgjbEfoqphZk6YVlmz2wh5zJz2wL2746R
4QSYLFggJCy1ZO0PUXuIMUSHdPjyQU5vzQ8RI63GCVgEJw7fxGMhVAlj4LDmbnJumgnzdSAcS6YK
NLLTQ7a3lIp5shvMowP8uaRIwgdWn00cRuovsZ/Iz8+5bGtFsYhs0cqXKXk/9QdDRXh9YHh8hX6u
xx+JMUK2YzjJTNSAnomfobiXj6q5DuZm7iXF+w0txPozMhrzNRaQ5sSkPfGNxqYNeHmIG+rl3WV0
iVCfE0cH5IgVi6TV+12e871nUV4QEYulYsauqWJZuGJ49HrZtqakZI3Qwy4oIslMJC5po0hj9xet
pMDtqDjFHDoBahHgw1B9sSpOcCA41UEVNKXMJaiVmZRm5u3mTNDdVENF+HYxAqj0aGgX2rWkJe9f
DmCBKShL9Gqdw8b05VLzFTt8zzBD+xK8sqaAUknIu3AorE9raeRBy2XQEWJDVQ2DOcvz6dB9eB0p
GzAiXswKk4sf93s0VhKIVd5ZiLh+xeGqFnqPq2ZkDizLwDA68OfMAx6jmI/KfgzxBKnbBnrQwd7s
HuNN0LG5QuGzY0SBD2F8kDTDtJ3n2/cttJDnPhmq2zJL+xUrgXcepI3NQBrXEu9n5LBCdq1m8vln
dPYw+zELuFjwnWQpheu9c8oYCm0mhGt6EmxksWs8+C5gvQJJqbKhLT6fKbVtWkHYeBwAxBR9Ny68
QHc+uTHKd5UEpPoEAoo+MQwavVTII8jyuF8DdPcclHkAmsZYCz09XhxzBqYXswPdpI+reer+wFOq
N9rFZ003y+faWaK5LK5LNcd1mhOtw4KuBQH9muJNiURtFg568VruwgmjNGrL+Oxwo8M0I0EBA9hT
+Z5oVe7HMMog573vi3n4Ty2n1yQB/Fk/fb+k8/NEasF9CPXPsrVIUu4E+M8UwQkLJs8QCneoLpG8
ZCQ4eVoXS57KvdQCWJGlH9Rb5vLE7yxWjkblBVl6fElasC+uI5r1EKoO9NvUBxSdW+mnAHzdya0Y
B2oJGMbLMP2wnJZIc64ZKDkwaUkjysKymWBv864Gc65nNvDqjo7lz/C50MxC0QLzlyMhrDqvZTlj
jb1lXF8VKK54wJW3Cyc5KEzTdXeckXwKWloVfbR4iow0xixMlHgBJtEdco40cJonvEtaebi2gzqb
+u1qNQjPaHgaHHoF3HRmSl1V6gPNpTMqcPOAiSdEkw0yKaedKZ4oUGKdrSHJK4Y5noFFGTHv14l1
KB5ct6SBd2ORb56z226Niupywuy9Co6t6l7msBJ/Yj9PTc4HlVclzl66joFzTJzzm1GHVwGifPO5
0ORlMv3pM6q81TPLEaz+KZ9PNXQVkH02hFUyEXplCHdzi5rVJqaNFKNnOR86n+hbzJ6iD7HN3ezF
HTk2errGQTIcSxcXY8HQQXzv8KrY2j7DsAl7W8rNLiAydOs6DRUkSJamZnrx7Kt9Fy6ixxesFsJG
I/KdOwliXvwHp085Xw1WScxO3PsfEwHXcnrDX+QP0BaN/GsxiEqtWtuGh6mv5CeqjeBVLHvTxCIT
qt2Ee5l2fqmToVjK45iX3RcxKwkNSzrjWtU3DNq25nX3K8IMbWoOKNUKlC8Lblv4P5c+jUS4roV6
CFUGYgoiBT9oM6WbjpVpUKwfNgZa3exa81PiN2wHqQGLDmR8kSQzgfTjLRd+FZeAZcMSo0abI+eG
7Bow4jl9xhvfluy25qlcHD6Eyfsy9vPTcc0PYsSQmJAxOyokkRCGFKjIecBldrBi9GYNMiVX1VmC
Oo/lAXqUQWjVyVvxQYRxmuORAu7MJKyKnnTtN/MOQJlRV6/OvpQ16h5lNavivJ+k93rtyN21D2qR
FGy97TLbcImKdUEg7PboASziJCPbKl7d64YeXMiYnmDdVTaIv6XKaT/eOhKtx7hvfvx+7Ku+vyWa
ptiSt3F4LCanxk/32CvfDcHnGNv+YQ0krwdS/zgR1r7IG7uCprQWWtkVrKFcuoCW8m7txQBtBesw
CKuUDvhce3gOfg+isqYBl2r18/wzTxU5O330SqMZfaUuJ2n6FRIn5Td8N2GQsLrjaM513yoQkBU0
Dtlg0b2CZ5EaUK9EPAgdq4nQCO5Y8fCYJvM1+vw0vxh06WYKmjpSE7kGXan3pCPo4sOsGin1D9/5
E8G9yOQjEg2D+KhfZlK7DjPBz5ZxWMLcebsztfLFR5OOSRBUpbymuHNdeQpwGBTLPUPGdURFGg8R
Tf+ASe0pUd7ESzOyD693uNfeOkqdAw26K0p0Ol2L5Mu+ue4Vr+L1jQ4aqdjPINK+tlNSWz0R/6g8
XOOydflW8VnR1oVaa8Q5Gsoal0LHfp0spYptQBjt2Qaa3s3Seww8pxEmBalMuWQvfEQgfBw+n9vB
zpAjX0kgFsGify3lxFJv36XZqky1qiMeGTaU4WUPNG96YN6TNNENW94QOuEpzuS39zpCNtPxARaY
gCdRTm8D92rBVN9b0tf94Zvp6OaQM3OdGI8Be6iT7ApAHnPpYdBFnLI2Ngf80CMXSHyk8XB4nd58
C31prlXSuh9Ue1Z6je2MpQmpD1TSLUopNUlMI9au1CUVyx3oXedcPyfeEVfFTJtGytjtZ2ljlfq7
srowu2UXRWJWTSPR6KwtKTdOm1oTT0GMiCZMKTGl25bPRGRl4AOvfv0tfKumGUHfwfAWYELlVU7T
bWGUWOPCmGq6sWDMXCgfP0ZcgaTkqWkFPAE0fniL1twpeSWFy7tDmqXhGAraBdoDL+Ir3NT057j/
KYOMQIwLuvhSjD4GyFBhg8vVwB0S/sK75wMYi2I91g30XboZrhRGfwgfMEO+P9kKnZWsJX9qPMry
Z+iJtHAx7t4ME2i39LMIFdYVLK265lODMxXuhEoACgq4eEdutHrl6Jdh2Ux/DQeSmIrA4psTShq+
nehAxDRJRnQnz0D62i99Eq5PIBmZpTQIHk/3PI2h/3MpiWWPDmCff+gSKGR+IOO2UYyYPTtiSmnc
lfoEcC+CUWNT4jlfoHxoB4SGV8aiPulFrE/NOt5dFS1ai6ZyNry/KoCYNjvcMhcwcISYgr+6Px9i
DpDFa3FtJK3/Jh/hm6v1zwIN+f6AkHI8OVuFGY9GBxp5SWPHaUzxCjC3nSYCSD/KsKjBcxuopCM2
KRBvxgWOyVHPEHOM+P6k3MgKuCEvlfdayVlrX93DrzpfuJJq/0LXX3c13xH97+oHMaGu05v+z33S
24owgkCuCS/RwaJFhPebtIlSAr1fLzVRmiqaEWY5pG6wRQj4L+BeQ/FWqU+LNp+1lha4VYqSV9jr
NPGUkjC2eTo0rjQZAIb03WV6lU3ghxF1Yc4a3+v+zsO3rahWcm/wUbrGYW31GZkpouRYhQY8HfTd
uXAUtQfjTHGazuF3Gbc0vI3Zzih9sPctKU4TXv5kera67x2R4HtligYxTxKmmAz9Zs0qUWsWdsXd
lJLajP2yZSh7jMarKSvL/NuCMSa07oaUHQCeezcR3OsCj/GkikFtS9NUOjt4YnN4ffcxXIOIj/Yw
H4UHMMjMcULmSt0zl75H+giwFJ1W302eakb+lhu2arwtTWafVWF+WmYQqSX3ou825hv5oaZlfvyp
TVFigsEYjmKBGZA4EivI8NAHhZw0bHbbXxBCnP3bQSYHkrWUa8FHlrPeIgJ+8fkz9BJeblDBLEoy
zX0DIHYQtippCH0qvzQPR0i+f4ZhiTe8ut5xtLEEUD4XGyRZ1x2O7E+eClAG4o8FhJuaqHysGPD6
fJoNc+PWuc8abj5yu/24Uyi6U2PIxWUbjfJlJBrkHm5FORTxVrmqvGHso7HI1YpDN06i0/uaM+Lp
vAtRrdLc3sGZ0Wto1S5faukg7wCvovQhYpzy6yum0zjw9aMfNZMkHYgON+QYO4fPSZQv91+sPsB9
YK6rIt+msN/26h26aJAf14gOYscaTSzg6A7WZWKqPqW9/a0YzbBJhga3U+c56GgkFXP92oraSQwv
adb4CKEzykB9pupEznBsqQ3p3HZkcmrI6gwtxtt+Pcy6D8qwfmhCSHzAgCYfQnAHKf/AL4PDJEHi
a13G82zwSDwJeTpln7Su2R0CBpzqtYqaX9rjAlq6vkgBJ2g1xHGdK7u4v2Gd8nvaGYDNe54jBPjy
eyMuo7ARoLuOjFv/wuDgOvkTLWE+VcghGMAH1k/IjoMi2POBj7VqhA5WIXsWG0bNwNT+0HaHHtNv
DUktgviwaz2ZDHiiZEL/1oV00cY1qj6SqmOBslUppON26Wi7hfIEyM7K/tjZgFxdlD+EZo3SIi7F
AjZHEGyt9HL00/CWseaDnzqcLjPSh8xznT6eBndL26L6MmSfXEEsx4GN5YwwehgM6ed8NvoOyFbf
JUja1a/kcBLRXMSzKgWtbLSrslCpGKMKUkzcHNre1ivFx21jzrpMT0aBgh25zZexLUvd0JuUAzZ8
YH36Xq5A8QZpoAwaKovNOz69BdUtmJcWkLsexjZl7dHvpV75DF/r7qkJNMUATvX7v/OBT9VbUHSK
GKRuraFndLCslDZZXI7UG4Hn+NfEc0s9s85e3Az7AzVSRYzkHsHKbL3sU7TLaeVnES8nFoABlPh1
z5m2hGkg5DlVmxPG0Q4fzRcLrvb2LdhnvlYd3MM30FtH/uvnQ4ag6+yjnl+w7EgrhOUq3sEIjK2e
hM+nl7ttY1fpL0j7xJs3YXX0biSluKsY2wLBH3VdNbo9TJnvvVAoYSlVh7vOkp6SQomjm78O5eDK
VkDmCDrpAlgyHajKhY/DhqsVntd0CaKGinEniSbQHUXgFhbl2xdAbrC+ZqckrzVwgvCl/h6pplnj
zMGwGqG7Gw/Qen6IqDCHBg9yEKb/CJqFdkx4RwRKUjRw9I6dn6MMw4H4Juc+wMUmmogaquX+nkNo
/S4qiCCDGXTM84uiL0CXNUyGlo63QrelNgWoyEIxM+5RkOfv9aoFzWm6ka+HyVfkxn08e56EqLG5
CpZ9dV8bT2a8Ve62a43iVmVdKZAG7wR/CPMZ11o6vzPDki9zjNoPr87lPcfsv9hbFvVDO8Mm+/bI
aS06CZgkXWcOFbfQEPr/GFn8THcQJ8V75LMK80ppKLEb7U/Qn+SWjwTpllx1RoHAr1cyyDLWUVUj
8xVAzBZf8UKJ8YMzh9gGwRHfITO8v81XM+R1WoVl4cAJSkdcZQmv9/dvtYB4Xy5puT8ZvuxeDa7j
WSUCjogcQGvebL2da59DSVHI0Hj4xx9I7D4H/nGEOnzDvrI9r5e+x16oOLr2ayY+1jBIgtIljubC
Ypppyy0ZWrb4QaKU5O+VPYn3T4JiqyLAuItObN+u0nEsuTTDnh+HrnVfWdlx4g82Loap+30B7WLd
G3Hbyj5KHgoTvg/BZionlvHaIzrMvXAnl12ZqDXbvVaTPLN7qs1TTd43BenMlltY++4/Qr+dt9r/
OwwkchwvMS+L/PDlxqUK0avB+vgAwzKRzA/T6SYsdbYy2X+sNfgzo+jvg8swQBzyMs08qUd5UbyJ
0ZvirWjm3zmVgiC0F7LUHc8qqMPPN6QotDCjc2Vop5pe6Xk80s7qCkl6bnMV2LvPCkr3XQNuuX1C
gfda/tcF6q7MmFkSjfz1jhSAfRBEAXEa106JhqZh+9g1ELchzMqWLKjZmRRM7knXGKedIuERrhUs
8Ixku1QlDoTwdS8u7CwjyO4TvM/O2VYb7PELujMuyrTYFjkI77ftsseWbJeQAcv4ZwmGbCscd9ei
hkQyWV0/hRPtA9l9j95eied3hpiXh2f7TQFqdC1gRoO/8ZfCAFIYwoG6q7UYEa6NJSzH271s1CL6
EOrEzCWYlaXRp2xGygNq0uB95gpnjPbK9bQJKyrq7b4v3Hrk2l+6IFSqSBB5ubnWPtf539JACXiy
AVncU9EF99orsb+RnX4S0P56puRCanlddIjDDp5KE49oCutBIQLtAcGRd9F2lVyTTBP56+yeiiJo
vtjUTul7bbKS2IYqEGxWy7XRiyb+mhAkbbMsCOsUvs5DgvonmBzM5PQUkPaj6z+XaVXukiREpEmH
1YkSor209wpFifHDDT93xeORLIQRx5Rd3IF1C9TiyO3y7iUqtsvTuWv/MmOpM6YGz98ulmCP9Z9s
GZ+7qwZyptQm0agu15kdLaiic8IfDxVOnadRsBz0JmqHkolTucoxvZ//SymIawkbUhyUdbxaTFiT
XQNIUxEKJG813AOG2nTJsRGIweHzHdcwFduyYwWnYLjejiLQOqh6UgwyFZeCqjyRXJkdYEKY6F7b
/SHSXs/OhIt7gMrQqzUbLFuYI/3trMa73p3dFBl4sfNWeqbTTFad+oOZlPuVoX0IgcUOhqgNHXKw
pd++3rt5PGCGz2KBpl8WwCsghOqWaIORf/Yk3GVStel9x8yyavPpmiFtlcQEfO+Eyx9ex1ofkhil
K3gLdN7NE6eBdsu0mKMB4wyTssVO3HusBwVJh70+gS/smj8txJCOb42ee9CrqBkfpOYaC3qSFR6P
j2wqzmcToiXGNmclexkzuoHI86WQ/X1LqZsqhwyl+H9MS3qSva2UH7BvmvbQcaxNDddGRAl3K2m5
/nppcXNDmxc2mJg5iRuos0ejmYw8ijU6Tpb2q+iHWpo0vuuJP37NIW90SKyl3lWdHKwzTrfeT7TB
GLBp+n1dWRwEO/isjwJDUHLexASS4hkaNlQzzEPCLluU+57paChlHQAzj+EIznQMRVP4htAi32bq
dI55tMFCXzVzDh1SZ4oaF8zInGk5JToiLODBmDeTbdeii+rU1EBYGthG85Wc+9Q1hi1g+oADbX5h
dEglztxL/QRKI0gP4kGQ7t/PDFWyYhTdcIaxOlzcGjYgXwaSmgII5L1NzR16MXTWF5eKgocvva3z
keBYPwZraGLV8dS3cfZqD1iHaXUGSZ5YZhIWkKRtlXW1MJVB1BiNt9eKP7i6zOdsPr5Ay2sEmlfF
bKDnFKIZnm2/TiK3unufmjMdvRpyiLknGzsSHeaqK7JRuBHw83lpvGh5CuP7JHUlMbxThiUAQdPe
ipj6byYi9uy8LMAUxnafOXb+LBpkAR7kr4wEbfLGxdar9ZfoIVw/k14EjsM+neFqdHNCIwlmBqVm
+3/TYPaNT27TCA5AGttxjt43rsacpFIvTqJkcfnWq8eVTvsFC9aqLIe21HjewUVFdHAx+Sfb4mea
1aNVlsiR5R67c7aFbgtOMry45k9DYrR7sW4cp0VhJ9LLlLhdkqZC7T87L79S+t/3Ar2B2ktjKwRJ
Kk/XyfGbAXBhWuLt9Blyk55SQHI0zg3FYkoHFf6Ltl+cBBj9JD8gic8A+kfyBb0JcvCSJws0xDE6
lPUIr8u1vMSmh/DN0eWb5VqtHqv00arjedu7cqIcfDdQkGyIXtmtNlkBOmVEvfF1xg9m42ApUCB7
SKmApxMnS/7gQryytGbjPcHXJLcLwvTzoyuX+dstTkD+AoKfwHO4kMcPzQm9xa/3O/VwJswd0Gj6
GquKNhdMIoQQPXHOD5C3xRYA1OdJrM+1nbwGJyMnu4aatdGlsdox1WteT8ecxaGvwX9sfAs7bsoJ
XMLEWjlvPHIDPlOt+ysqrOuV2UUiBkLFanhyiWapx0Wt52o9NVW4gHh66Rv/N3lD9PjYiUbYXTl7
elApX25BAdnqLfQxFu6dNzGNCO+Ec9uwgLD9yT49tnMLMH3aHB4xvsSLbHdPCdUfMcm+Bpn9+y/q
/8K5C/I021lgEZtOSyfBjmFWwy2kvFz8MftY5hLSB7qX0kA8iA6Y/7aIpIz3T3Cp1Lk8nm7HsJ0Z
sKVsWvfR/X+cfYxX3zsyKWsrTVgapuyB65N4cKqoo5PGnKcf0S7AH944vHCZ3YQTx58HuFq239sS
+BeEqzen2JHLO6RbprP9Hzacu5+JlWt/UqOE2ZTW2xXQePCL8n6yYckQZNRLl7S/QyE9Dxx5oIS5
ug8UI73AvVi8y3iRW29zf69R0a9sEColRyzq535gaWaAtRvqeqmmq4GXn2dO6ARe+a+XSwHwtBgk
+x9ykZ+2vqYtPVJoCWtaUvfoj3ByB4/tKwtEIVuPuJICNJ0xzZruwsCHa5BxBaCBDFunGHj8BGIS
raMgXg1yaNSeOPlm+PEc7Dbmc2DvlXkvqhLuwjUhzSy2Txm4xx9MrB7oS1QNWmn40eIvfcyvQFSt
b+kHpYsX3Pi0YSmxANxKdctJteuITtet+oRsdhoCa+7yWVNAzXp+dNFnL9hx5VOWF10vBzuOtVeh
4j9K3acnJRKcGznWcfcd+xrfVb9QZ0x+qIV4LMA8FCRUWfSNAYL/4PmCOnmt0MGdeTLx2SWtxEvJ
4uIZKS117tM6lEKyoejjfOSc5F57F3Lgb/gKVKD8YCqCjZmtzHH4un/pRAF2VO7Dg6bDSd2pW5EK
7iGi1pzUtYINRcn2ChyEdznvgCmSoW8qqGgH8YjaQsLgBwp/iuJgt0Gvc1rWoqnhQptgY2Uw97Fc
JpO6CQ81zdhE2vqH+UDpwR6N3gk1dgIbR5nkyzX/i5iobTJayrOdbGGpcSlBp6OE51YApKhGsRQQ
0Rze/GssE1bB5TCOGBBmOnWSzXECDpZcIc3voKbHwybyYaFJZl4YJ60AVeFNDQTvaMjM18ow+vbC
sEA/w3m25I4SHdOVsAAGkN39r1pw8p4+N/m0tMBuEBmgt6oEYa8YHD/MPO2jPKL9HelDLuP6ey0A
PKSXqNyMOvBivvmwxMftWo3J2MzK+YKkAwBOmd8Vg7cetSgou7UgxLAa1B4QGlmu1bSQ270NNeMW
+FudpUYpy/eBJ/GLkGJxKJ0ofahQBC7xXRoCrINagLkXb05+jAC8a+AkGgzdL9t81RuZV1GlR8hE
jkouVuSvLLkMHQO7KO1RNIb+cDB4XH4zC/hVB3icep7ER4eiMAYultdbA6ovdgY942/7hBs3suGh
7sMECpWWXoAU7rOFhOfK4zvi6cL6DTk35jyIaNUpwhF6AHX/GtEqGTKzSa/sJJRvcWxMW3q22z9h
oWVYRdUk+EtsQ9G76T1Xcku2aB8qltdl5buW4mvv/yZdfTmno82563+ekUq1PbhZwXdzkIv8Vq7Y
xh/i3zIrE5oh62x198rxCLosiYzth7sdjnqAbsYvMAJ0bPpZUuvys/h7KQsjqIxOtGLV+G8w6c7q
nM41XthsBJ8lll+ImIm1e5lng1PAOiEMlkg1uwULZCpM8djWKPdZHiJwkZzFrpACr90NBJT3IV4+
0TFSQoI74f3XdKJWPyom/6pJmsOXKrsyrgPBY6+JgZXzAPhGngWxKl06JVucbvExP/RUrWaXbpym
Y4UD4JPRRhWFHBHSSybV5WUS8bXF2utumXrBw0XvvnEIPe+bt5cRKT600P0yXT8/cZNzgScCQUHL
vMWr0jXHrw5UN4EJ+9seEtD6XPR++t7knSg1Zbhw3YSiYiZEnlQziKTD8+XvrT4W6kmwbHeh5qss
KbrV91V/2Ud+NBASPjH1yQshyILbLbs8yChBd/sxGLCHgftT2dEqOKgWHTKc8dZdXquaqI1szwg/
ogms2hfzcuAHji68lV1RzuXvzniGHodlphvVFtDRUHloj9jgy7Z75U/tyEq13/PyFFmHRLZd6vq0
NkqV0Ki+9K9X6jLB4ekgrVZHATYrTMsxS1gGgwVTndoT2uGAWortFi23uxFeNDSoIYIO/zJVSxUu
GujL7eD4ul2HBOAXYG17+xXP4dgds5HtN5/998mZWiYEAOVTXwiFkiC+O+I6+qRkw4gAbXSElrw5
bwRicicd38bl1nYZ0Av8hWJ9Jmlg4xGDUv2MUq7aCeTgvjeMWcz8r2wA019lv2sKMCBM8+bn0p3+
Wg5KNcUXUI8sYqFFHfxuIAOMTjb/8W1krGEO24vyjeb865yIflXIKW0b1xu5z+YqU8kztMx9uV+G
z4KIVEZyTVvAKY7MJg/X1z38W2O5xMlJUfWzWHGH7ULo+g7B7D7gUDcfzeXrMwTC5FDD/Gkikmsq
JtOi+kxy8I/0mUAtkFh2scxMOK5FtJ4zNT1lufjARojZ8+A+JsztC7DRvewwr3d4tUKznre831mt
zA16NV62DexlUD+V7qQd+u6vlV0KS+HE+rRnzA5AwE6ngDQVoqYKV3Ts7RCmkOmj1Ed6r830jR8Z
R37beOrmqXW/YcAV9jbR44lSipAT+8rvcvUwpCV4D84ut3TT0vbOQi7YfVHJBWofo5ZgBNE+jBYu
IOQ9QZtdg1JOkrQEnCmqXDQvgDfyhPqX3XgqYzEdiFV6Zcy5QB7mVAy/nOH7rRpyUl3r0cG294cv
kRy6Ag8cWo4vne/IAIE6VFSPOBmaCK7y0WK/Oz/hWNsyOIQRQzkbIKTOoLBfxT+UHttZHwOgvCJj
r88eift7yLVrdeC6VfDHX/D4bv8zGadCr6Gf0ayrmSTKjiyo4AKNotQLFtUwKLXpaonT3w/cxVMa
BMpX0FrLcbQhZtSXV6GvXaJP6E9gDakO7gmDw4cJYIIdOip5uJpkwjEcLlwcKtb4DD41lmMYfjdj
IGlD9GAthO89U605kjRpnvYlCTJRK6uCifkXiXEuVOVMV1x/+vL/PZw32i2h4ftsDDoIktAvBabs
Q4K1qygHIEk8toq4UDnd70el28yyYE+qvN/SjYcmMcxXHqpwQfIaI5JsSmNh+ZIbpvrpG1nSy8jO
JRuydOuTFVKE6h+4d1qMVVeRvOe9LJQ8sA0tjgHXLGGsZSgU/a+/ysAVNFt9cqUjH5N5PwpQX0Xp
hjrQzwULhsc4gs/4x/xKNUpu11Ki6NQ9KxnSVAUeXhv3lIuKjcGh7Zvo35Y4I6fiXLemtAvPiDLe
eqwYcUiyj08zkWNoE/z1QpiIHYzoX7wTImujhBexCY9qTweEOl7PUCdsXyr34obJxvMhvZJ3qNwH
BNVUm9UtszQN3YdQr1uD//+VPBmox9f4J7ZE1DL8+RFBFX5LlCF5P4ekiTQ9KbtFxn2bnTEShdLH
4PP5OLNdNA9SnjqmKiD82vHDXhBjJhA5AfdRfQ1hVoLNVtBdbquIgsTN+LIyVfUCizi6EydVuUS5
6dlDtEckX5T2QPH6hHHaRwMbXoy52Wm7nRJK3Y4BooJPtxX4LnlNKPrzZ8IFkysK6Rl4WuwmBIWn
KEJEFoEe2L0DW2SfjwKvNjQhFLT0SwlMyCOJw3xLqvEomKpytLRBiHwtH5hHh5K6d3xh9AAXUpa7
Uczg2b3tGK7uHrNnZqz04t+hpWxR2FGJZZ83I2I0MPjI0atd8CJYpehYGh5YqsT9dwWHiC86IBS1
mPEIPGHPALrN7N8GRLWC3+KlEf8TSggtKPrYmC8Qr49tHn6vO5njpLLM8MAfPwMS9hX/JP9cuxiy
4MobXYVT65xUEkV3eUVP2hYRIh+dQsmE20Nh0hhLYJrVm0htxDQnakMVnTVUtKUgUsKpJZ+DXlik
hLmqaTb8Vy+DIk4TrgxrfR1VY/znxw9iT0kEe9hZsgF+IQxUME7XcbkLF8V4SKnHEA9VuUYUD2Dv
RDR/GfsUvo3fUEJOGPrfffM0dE4Mf/tDIRg0NlYd0BY1k6L2qOEBeqN7dfrXWtEMLDryd5JPwu58
htTTeMhXSxXflZSKVbSDBUlRPDM71v3zEy5VHwj/0Lc2wrf1Rj4AKQDDIb0WOsAoWe71MmAxXpyO
nKXjYMu6HgkZIIDHvwaSjyQbuRNqBkDiE/uKV+cX6Ncc8rZb8J6zBet2FAmr9jnB3pcIXteWQ0i8
PT4kNC0N4rDUekxTu9sDAlGo+guVk44hMj+sbeggKmNk62UY+R2kiKlZa7yujOee6/FX6+5EWNVw
vJM5fFUS8BoNjNzxgH58KZvdPMPC5IOn/fVnGlx2LABeXxukgP0CulX3ngvW2ONYd6HCbFcCzk9S
2/XEytqkpKCRz8vo/l2GUHcx/AKOl9Zk7p/1kK5Kc9y/7b+RQnWqLR3y8Zw7EevlMEB1RbWJJvB2
GFul54zFeDNgz/BQJ4KzeYi/houKCErU2h9H7nzGDOYllzxUNB4dXO15ecuc1LEpW+F1fOU/erQl
uM7YwWcKnLVdb7H8Xzqq6rP6D44KsWY3gNq+PIbdhvRwgBgQYvqmxOLBwQbMagHnZcha4HVEMy1Z
att/5mjtvO677l0yWRbPPjh1eASGTxC8BHJsQLcuGOneSH2ZqRSZK4hGG6U2BI42TFWdu2JsdLcX
eEocoOzpHUtR05r3jx8/nviHwixZqt1kCSuFLqx7CIEuNB4lM9el6B2/LpIR3/Bih3XWMcG/twj6
085wHrZQ7cxgXl8+TwSr9u0T3K2Vf5u9M59KQdRv+ypoNrMshFha5n6I9Lj/RYQvcb9LiSUsfF6e
mR4sSO/VFPcJmBvyPHGI4j1Ne+xgWT3RNo9jQKkEhZ0xPTeSMaTuuhA7FRC7B2rqNvOWexe4Vqqe
0vtsfLVPcbEGdpw1IOvDa4vnNLB+vnIcsxVYNcMYGuitOdnodFI3LHxM3m+anSIXuA3EvIJZbM8h
l9EV6hv+A3HVQpgcRROsKPqGmw/9xtvppRT3jHPnIJhAGzsrzz0YkeCuSBuQaR7Mn2JZE9TvF/fW
0hKDy40f/C8FZ/AzLHXggBs4RyDFKp4ut/gTdlnjbGqLAr2gXLuZprEt9Dz4/wO4aUcAQxAgC28u
WZBnPjxSTS8AJN5wcNX+96KvBXzBAAJtU3m8qBwJHgVJT4G4Z91em3DMdg62GfOugsGF1Ql0MW6T
RDuq0aK9VBlkiWwdmXPN8Pn3EhQQOBLcNYnifaNFooumtpuIuVTr78Mba5U3eKeJ7mky+gNMde45
kmRNq6XsoLzP4O/3zoSSjewRnD8RmM7n/BdONh4vrnwFjag8SVFdLxsk6yt3pIcMwl7TDmAWavrN
TfjSXK+KNqxS6q2psWVw/fPRMM7M1smVQkEG7GKcBz5EKIT42kBo64O5GL5plvqazgPzctLGLxiU
jyihsJer4q+up+lCRRSUGcsSI2DFrcXcSNCNI7aSDvLkwUwkdbloYdU4kOuPxdZG5PO4kga/pEgt
eteCSzHDRG7CUf1GU8rgo0eb9j8XxOo6AQM8zhlQoezO+LHyO8a9D+8jzDVl3qDHInrp1sIKKC8m
f0feqHpycnk6IvGksTv6Yha3mNssejmrHG0Rp+6eYU9A82hsEe/LRpK1Mfw6a2SFXtNHl5lSSFUR
5mOa8SnxGzxpYU2zhtG5/DrQEyA3SWAunqjlZ0yN19qnbeAL6apUjDJcjDZ9HvmnxoOSyBrf/bGa
/wTQD1E208sxlfO+U+qpKwt+sGp7va4v2fmsEJe2U0/zQtjcaYphRGE1oM+oWkMECnuKgACqJYn8
priIJ0gCJJ9qx7AvltP8flJCNDc0POTcm5Ql8BtLRX0BxoBMknw4xIbQLCV8h3iImmGsduHWyJab
NnMj4QToubWrQJ4Mc2M9ZGMI0NVeDhgUQ/UzhDOlCghHpnRmdksNZ9lpdBXYaJRVTtG5G/VgQeqt
dV+929Om3PudFWkaHiNGoerwyauQqx0IwUhsB4Oolj3i0GmDxxxsCyIqHpyPAgt2TTUvcsKdmSG6
io6vGJ+r53yL+HfOKyOmR8ZAUL6GqCrl0q3+cx7AVS5SN+OPRp2zRkZ4mvZq0ACob9NbHeB2iIIW
WrFBKx8++03rmhiSFWBqehjJBIsFEdAHWtv//uAeQpbYk/hnZpaj++gu3w9wBk89YBsASqHpXSWF
W0Mw7iaEXkln6do2+dq61TcMA7vKOh+SsoTRAyj94/2C2b/MZb61+mMx+pdf739W1D9VgGBwMptD
ID/JtzJvkG7d1+dAMCFS9yki5tucSmjHHmZrk+0qfxG65WdfUQ6DzDkDColl8CGcKxfFGIDw8fC2
XJo/OPTJ3xyI9bBofoF42XMBH+T/E9oB8mL/A02ySYqzQQ3Fhh08wCRlzZ0bUJrNEeHg8z1mUfoL
s1PpDl5H3nFg4Z24wQTV7AzMNjHkQA6RinLvsvFBoUO4ZGLaOB/qXdAsN1rj9eKaJbz39jqkYD/3
4eF4LPySmZBPvzwhrBc8bwFGqHpph2H++Tn5BeT2vQ8XvF9uL6195b0SBiUlVGi6vvnbnDXSAwxy
/kHf4DAvw6SeSQaUwzpRnJCb2/WG/+b2IkeUv9mxePwJQeUm2Mogu6mwRXAVOBjIJ1D6drzrM+Jw
2Awi8G0tehlt4X6nsk3ShLVNkoldULz9g1uKYpCxLYwcy1NB0be/WI9j+Fg3lxCSxFrRoOTz+rT2
uk1Ng6BeUVt5OaNBQHoVBDEipQ5XYKKYSKG6Vhxtp1BhuLTOcoU2sv0O1Oj0gZg9smMxhDP/YV6F
4hWrJ8AFZ5xH3qanpVB81+Q81AyVmz3S0Je610VgEeMtAyK7E6VXOl0vAB0NJwK/Lp9HF4Cb1Av1
7vPJXAzddXRrDdlxhPeahzGZA/CeUj363PyYO+vWvs3ucUNoSm+q4Xej6/Hj3gZ+hWAVpyKdeyBt
RMSztw009CvJcTBXWK5qP9rn7YJ3XhxSsp29bxcexk85tWgCiQRttToKQbZssEjXA9CynFCXB7wd
19jyJkPprafz0pCLzrSu6V54s7ebLpeZu1QMoXlEBL87RpC4r1p8cCR3quo6nSu7W4H9k9kKvDLx
tBYmxfWpweW8oD5AgHVaLiWRV09TcM1D5svvfpxrFQEcV0BIuBvSAsGGSCswx9klk2SDljJG5DeD
d8f8i79wRjV/LHCfpdGEGEyCh7MQCGTkkc6AONVww/2WBguw/MFYhHIEiB6sTsAncfLPolbd/nBC
ITsARHdm5A+LsKcda/Lh61VwwYK2U+yGsJNlmfz+Zerc4C8VWHH2TfHjL+ZT8YuP/dTMSjHaxlP8
U3DDEfYO+iVZfjXQE4YYD4LQuDObjH68pW0VYz5koeF4WBI5EStR1ZMkZzfE1ti8yGnCvfahuo68
zTf5KOBIpzigev/OR/pwPCR4Doe7H3914j5QgrD7J7BGzQH3HUJN4C2L0ZOs8OUSemv21jpqGqSM
ZFAIp4DRdTNF7d0Be90P5bluCiCBX3P5vcucaF3cM8VG+feTGte0SMP6RhePSXqEHoIlsPbhGQQt
vR77OPwN7FdnwYq0CiwbdjJqpgD5nivhm0ALLjhwTgFUA6hwZHiVHtlXQpL+6sLKPmmaO98XNrQu
NO0jbrYc6EhnNrD+z9JAPMeS8QZEUU525NrjeiTBAWAqBFAQQvNF9EGRs5kyLrfG11dpRI+uOmKJ
m1Sar/+IKKeSIAmuFTgySZvs08BiCfMBSd1laBEhE7BM4bqcH8MRCd2Ym5wiEa4hqwQdD7pXwrtK
6V0ulcMrNzD4eJNyViFSmMQrqo6DiMhDsccHR5oDGcoQSaP6c3vHhD0jAeAs7ihkc2rhTdfuioag
waXO8VHG4J2WqPv9xMBLo+oKUgNwrVZNzFYmvITvXd+0M37oAtS4meLFYBAhBBqjCkSX2uNdof1L
XOLMpOaX3kkarSfSNcQsKWBna2mA1Lpb9IxFW4s05fq2DjoshaUPdTL4Ax7y5NDBDVhuKDuqljpt
aajJ9CgD72dWQ91uBsY0fo7fYWn5yX4nbjQ6G3yFIjDdxzVXsuAzQUPpDrH4blh3zZzVm0P70wum
J3/sZMNsJc6kL/jtz/mvSQnoIwwSBL9MrQ8wzjXlybW7OQSgBm5d2mVRrsFCdNqKMALx3iFJ8bmL
ZmAGunR1ckoSv54dr0Zyf7Kd4JkDBEQY7ZveBhZconlKRGOmpStl9KKqvWDxOpR5x+0j1HwnYQA8
H0XXlz3UYC5HlkKMyqKTLsGV1IavhZuK6/9AqaVMJKzi0NerQtYaGESOUpA6wthurXA/yD5b+GBl
oLDa7AR0iscp+Gms8yTUIUrFHkWejXPUPktR3SGfKN/Mts0rVI41oLO6XnHMTeN7Uk6weyAiSr0P
7HKWk/fMdCdbOYYbkq+0gp3nDBtku9UR4Ca6A3JOD/RZ4kw06/jCQyKdzeOtGfDSFM1MFTfiZ2a6
6wO+LgC7NTYh8+j0jsbNNJ7PhOFSpzZOOsWTa76EA52bATwHnJfKo429Zm5ZO48x7GnAuFmbucBp
KRW6Q8Q9iwBZkYQiLALWiVxMagcVFrI/YwrBJ1rtxuMqOp5n2BQ0gqBcSz75GQnrEP5nJ2RfmvZD
+trQUxaEyqf8eeHnadoUOWnj7vFvaYCAWOPuRHSorFjBLnCK8v3QpzXF7K7ICjr06SPJG/e5BsUO
9C5M14fl2cghA2rgBS/ftuUUg6C3ORc3OqP95OK3q35D51YGlFTl9bxqpV1/OPQVa8SzMW2BdrGA
Ef/ajve3e/ZFiX6JdrrCaA6XmcfVglJdPNHIP03pSz+cR73/l03z5jL5jErQLX/QVbjiVFJpSTj2
GrCIFQDNnxFkq/Rzcdpmvb6bxqENuJAWeuCnK1luX4ekHW6d0Xoy+ulLFbOzdmNEWmUs+0KcnPGF
GxFkR27dBUgt2sQMHkld/+s6AHbrWmKDJZHRJ5GGF4drDfzbA1M8+mAel97umrMGeqCwwW/B1Tza
SxT1rcXeNn7ZEdspoJ/DusnaZ/eByGvnWMp8CY2PBq20bWe0vftnt/CcBxtFLRz5z+dDInzSf+7k
O5Wp4vowMvqVW697HRY6YHhZRr42UKQ4DSSuBpKgE9eh7JOqxa7jVjREFMQiWgKK+errUqB3cepS
6JWyzdeixaf/9o5Emqtg0KP4syuxOfx0YUO63qKjLnO/KiBf5+xWbGLR96V7gfigk/teE+ireeqN
SbsDZK6qpqMI9Wtqk+zoHFdUb0pCr0xESDGjGYQkv7UijUyaAaoP3YaZRLlrPjFJJ+IQzYt1/O1r
kSe75bS0QpVHYqK8rd3+sFX7uaj5BMQ2ENcmEaxiKNNvV+iwFJLvgKbr9pbnMowOuMRTlIbClKrL
fiA6scDVziX9t2xP4RY1rqvYx3KtYi1mVcM8rgYIvuGenU5YeQdbyjuJ1skZEt9TDLwClKErInx5
J+zh3lHRj72xlwoHgIVkD1IW6hxjA9BV8B4pDMBERE+GowZziA+p/7YTH69PnwYUnkfuHFjGdTCm
9sosq2dYLpFDHP5h3GuAhWmn3EcJOFiYV+5xXtBgOYfcMxYW7CoBjRenYL0kp9XIW25miAAE1wFp
jchxoyT0orTQ8i6FuRRpN1Bt84CQck+Xzafi3mSE+lsUT1q1Em0rnLfqRCwC3jMimUPBx3oRiNZO
JDe+Fx2JY9pS+qtQr0CjYwcgJPPHclOadcRD2jystdCGhichuNK6CYIlZ4I2irvgEnxKbrYCnK5/
y/O0J5AfYhpYRben+7JzM9PzbQ4ePRiNURE2FV3ZZVh5A2q9yNeynNVjSmN71a/CAmwZmQqtEgY+
GDDppFpXa/3emDg9HH8apG4BY4V08TFSrkBi3xy1s/0/GgNS02XCPKHTmronCwCBPtrt7D/AaOq6
VHxG2AJIZgtlThLUSR+YK7mm4jFZij1t9uPXtcvB13ys9fQlF/Ek/lmD35dGEqlBJk83ISR38OZv
q+5VNRx28gomdZrmcygXC8pVaR+jnygr6RQo4r3Max5JzHQb8iJFdbxXdOSI0RVQDz6UoTTX9P/0
eTiX354Zmkaarx7Aa/4zTQACUmovdO6zl4xLL6HBLSYTolNt13HQjadvEQH2G55xwEUgWzzzw21l
MHF3Hr5l4bVkIOOwD0YcwkEXrO4jbfmI62BxnhCGwNk6KhKijVkDn53GtuJu0nFkaVWZqtSqZBJQ
Ced7sWsiiZeq1vGcWUM+yFXYX5SK79hMq4dEWrJp1us/G8/ZlmgmViPIWgcysx/yfwdJwgmO2nDN
cMxMm374bXFf1vU/Lb1myMrJz1Ib2kpYb+6BZ69BvjAtLhcFHHNkbZhX7a6kyePjqu4dcvT6DOtv
lWNMoLqAeVBhyXs6Yxj5ofn44FwrLZlKsENJ+7tvQ/2NYaiCMYhLSNB33rCXk+ao0aAr7iT/wxf2
6kBcKmB98D8vGNujYwvBOP39hBTSpnVw3Egmnryq5Hc25t/i1BZY5+JgbHjQJYXqdOAlXmgiSIvQ
wwDqJwsL1DFM6getvlxTyedPIcE4TCJH8vusugz9TqhUFE++kovYUi+f87nUseUcI7DCPbghqS7M
B8/71ueyp39KKuKfrO2+h49iRGhbcFJ24FGDle8PcaQ3HXdoqm0OuagXg0CDPvir6J5CeIE+5NgP
Ga6iz5jrWW34qig0kqyTh5Uj1ozA4uWURy6qNlWcqLXv9f7MPm7pqevyAlZhH9gS4mk88fF58vbz
C5JqXTv5HSG6CeVSDN/231VdVAqx8H209OpBK1bG8krd7tNYPozxDSu1jYpE+PIsjAvsEoVS1hg2
sRP+xjlIBUfCXaUutegRKA4MJcNt1LdcWWDwgQ3XBhHnewXiwU/KszU/CEl4kX5d8eZrH2AtVNjx
ZoOejn+uQJz7W5pJsYeHx4QSO9EDy9V7a9UwJD2bQbYSfRzYF5CP7Xw1W+sBquUntN8tGWGkbL98
v09QmN/CM3vRzmJYdwE4PPLKpQ2A7mG3VDUi5mZwkiq60PCrnC8emf7Kn12+YoToSNPNWT4DPEU7
YVcAO6TKB0LyBhueGMExEdqKl+6oNkwumHfWGjoFegZGu6YjHu8VZ41AJ1UcIZbIuCPpkqhtm+F+
XccHg9IVRJL/0dvBR1BcnyhiM335WLF/7QuMmAci1d8ox1PgcG+TMch7IDxEhA1ZvbSVhLc9ooCw
ThZ0m0rtQgawBfBD9HaTmkpILOwBJO85OHRS49RZUKr0eacCQ3aGWkEaTv5JSu8UIPre86QyLYdT
eNvIMemeM6aaYE9ajhmOjqrzUEVYyWHEtmqN5gmRGjaBcPXbqofdgV1CtjZcj7WSO/K4sazisdsQ
OJHSVyDSB+EE8Ox68Ny1lj0k88nbc4OL1pESziYWjmlG3BERwwq1LW2gCcz0IGShD5GSqp/3o2h1
EvJPvfGLAx9XNLlO9pHQDQThDfI5C298xHFaQ3JpA8xbRaBtnWbBeJArA0PYlVke0rApW4MBBDaK
TFMkFuwALcC4EuMXg2FjkUR9w+UoUvB3fGOYTwYQzz3ZmWNTZncclPMitegBY6/Je5bMf3lhaTPU
EE1GYqbxhJES3DCuYNBdd+KdUOPVrKppbedRme4Lhxg0TUEVwFz6i0MoxiWecM8Uv/7Romlt4/G4
p6CzyB7kvE9c7rgveNVWyziTQzpecZBlTc79IS3D2UusGbuIHjqWzHVWgxaIIZXhoxHSQneDik9p
P78/3Wvp6f8PeGqiXDGwhsT2CPj90j1ZdaX9O70q1gHPjaIpsGsAv9MUtgpX3GkZR8GX29Z6O1F1
KlHWxlIpJYdHPjEjdVAbBA5QZOxW6hqxAO8Op9Az5NhEbyoblydLXjCCdAAVdiih8HWNNXuQyUxU
thQ72hlJBfWWHcemO99fxGXYwMcHenu0NrMoI+kzvYu8SOtCbLXwquKO4TLs31B01FdXP3jgtTYX
H1wx7ZS2xb/f1tg7IGFZGGLsMXQRmZN/JIszgfaWXex+zhlR8KppCEXwbZmydM6cdHrDsz8qL1AF
D4YekV113QGhIQ9Ik1PaXFo8gZEpmkzlGyVeXyVp782s/I/Lil35nGgGNfSxgdFzWkxM29Q2numK
gimcv3q+7crIg7WglR1Dal2czEj4yTNTJyWdbkkOVqevsr9whpzBd/qseXOXkweKe75B1+wKLogE
kSQHfJ6TSVmcm8jsFejY0oj/YaDpNCBNIeJYB0h9dGKUBSJBOF0fmu7rojPQk23hGa3rC0sictaj
2ohDLHirtim76OR05ahUkqytb9RUn/On8Ne87a7MYITU3uaBTSHM1a3zdlo6hGX9gdJ4RvAftXIU
coxslSvmUgNcvD3CAtlt6MkY3PlKJlZ5JS/JcA1LfKKcTezoK2aG2eovZYjqpv4A0/Ap/ly9nHz8
1MLkM0yaWp1CR66zkmnGiXEzQG1aiiHciLzaKIsGrjbKNl4qAfhrN+MU13jBqn5XlPAmLy++lARx
NihCLKsc6fJT9SP/UpFyv6eDqCSOS/x8VZwBfeb6DQLCVEuiH9cAzw76XcvCvxouU4oFDDF7zSOS
KKiRDAWsJ3W1zcDjMnTu3umuVsK++qAe1BKj/+m71qf4dCVxhb4c2rFERUV21fQ/0Gn4rv4t48T0
Hc+TfOmE2i5jM1++hfgHUzADFXiCkuXMhnTMln7jRA9tzyvvSuFGUVCCsSYnlfXSptujMLSX+Qx9
EgFFyeTL3l3HLsVszGDy4cUSxuEGfhf0dl8hsdP+uZmKsRuk5/oMRkcyLhZW2DbZxHp0NcAmFgr4
YBAlwSaNNsARe5vxCLcJXlxOWHXW6qWATmipU7E4BZ7lSagUHQlcaAlDB7RMB7FgJ/A5V6d3rNlx
SoM9tmnqhBBHQ/T5FD0RFSPo1n5KAU3U9HgBYA50F3CGlXn43plebv5UNGpeAwbDCkJQrh1jnq6i
iM2S/VUGEfGXwrBHndZfd7qvPu5wQ3+zDT+rIJaaohq0B0bVw3nAXO7NegWq2THOdQKU3YtXon0L
V8SEAWglc7GYS5S7Gw8JkKwsgF/OONxCVEBdDjOqC1PEKJjzcZUdjql7VJkYhcCFjjMqrR128adr
BlO6ZUyksYCwxrRqvSO6zlKJaQwnuCycJIwpGZoI6k40yvSpJDrKBI455oT3/Kwh6RAODEB3mVpF
xf//+nxLlN7CvoX3QIS/JoPHOSLHwUAib1LRJAUh7fz9QPbKiqdF5ywc68piPZnJDIeZNTfaISnb
LQ5aM/coAysfBLQAwO7Gc98xgS7Js1FoqRAjC8/YnAT+d+NNMScLZUWcUBco21FaYE3I6OzkrL8v
7QRoQar1VNYho57uQ3Z00sDUDk1q2W6gg2SAEnoHJf4nQc8/0hWBkyshRm7gR8K8Osot9LovKmNV
vuh9df7QeHOeQn9SmykKAUSA66U3BtTIqrFocBEREy++h63E277+5TKjQLY5vs1FFEkHPxhYZpr2
j/yR4AgAi/Am7snvqefSFtpxFHMl918bK7psH5Hm9Rk0BSYFRQWvK+WTW6oGIW1RBOnhY2Gv/pMK
epKMKeQnEVGCQxE8e+J3SJt6IaqESd5K5XwwmCEiZWB/y1lbjy/STqJDlZAdwy0qydIb6vHF2zdR
rnBEK5jBqt9zGYyy+ubXLQEoO+2oC9aDJB+FTEmUmQEfS0kuPyZcqMI013/+NFSW//fq9gzChIqz
Cv7GvKplUOS5d8PXV9Hh/PHaSBMmMLtj0TYuMWKWz31Lm7jAmSv0t88f9jxrDtCWpnpYtYpbpVd4
px3oV9Fvbzh7LFbq4xOpG4mfbWtPsjDKJf9Jc9miw3rs3V7q7TbC7gsGPYIJvHS01JSVznNtTcN8
y/rWCvBVNwiH42aYvq5R+/LorrhLcWvLy0vpfd4Qg2m2hnMrWQTbAcBrjxKxC5O47C9vDVg6vVRp
IfQRncZQ+wBiCXMk4ULohyQDToa36SASBd0p7gl3XdfHmgXjn5Fr8K7L5Kazyn+VtSCtpXVXtqSs
VWFqZhGmaRnf3zrgNGuEKSX/oSbqbQuVZLAH1Au1/wH2hf6yYdlv79DHVYH4gaeHcwvOiTSoNTyb
K8C3DSuWyRCABElMSmErRMY4qBak/0qLsKimsiisPYKOl8MV8H8pzmQrQS4S2eBBJrAxQENyKXed
6IHyi9cm9s7RfifAelFweUgBmcOfMOLFtCoUwXrY7U94RCU/A5B70yEvVfOPOa26XjYK3R3Hc3Qg
Dy4ZcWZr1dMp6Uw6tFEiygaSDndn8D+kYU5pMsE5yA4NqVT+FU9qgwM2PLkbi0wYWZr7VcQbEKpo
LxBcuslx78zhUWooi76vjiDfP9sqwTiZbojvjze7XzmNcXdjjkce3ZPKjqcU9PcKoq84kMiiDIGR
yQUK56R+rhEM2ufJAJN367S6bKZmGpAbSehpTxZeFovAbKK4cQoR07mcgwmmequv1C6WzkkJHpCO
kk7c5Fj3VaQqp1oszfITQy9rrJ6j5KVJN66+uOiS1kcX5KGwiLtHAbHd6HlMlPA5gd7vc1xt6DY3
byc4RujcSfAe3vXnJHiZSi/nW7iN1I1XAuN7iyv0SL6M1QY4YuqHfApBLQ3eW8ejGsnsAuABhk52
O+RK+h4VxvK73TbrxXvhmI+9rXXJuJrJcYz+DTpLn3hr3Im44BIr7Qm+glZEqAxXXI80tXYvcu8W
I11iU+7vOET2oDEKSMUS4Gqfb1xcSY1J/atMwIuB08B0DZEiQfQ3X8deBXobaqKOIeCPkAktJeOk
to6FcNSnBgKnH40/RlU8xFTxmN4BpQi0yrN/vwZA4knKsKbTHRQah5rP8sGEPr6DOLS88d5GrCta
FQokfiGEwCUIVFaTAS+mgbNLcarNCJUUgX9vnWww7zAhraEJT2yeMG7KagFAff6uJhkHloGnnv90
ZkORwQiMPONP94mJ7D4QURkaII4QiFCUBC6lpobbtCRvkXcDK/uWIHu9E0P4m8fZr+hLMBlfeIll
NtVL/oCGNT6fN0O3/eOF3lBs9YRa7bzCibcw/QMn4EwkqOWyXoZ0pSktsT5A6ORDjaX5VnCKvB2R
Qa1IkZUdd/Ilmh7+uNg/AXUzXiuxzE8eEe2pq4GUcgA29yadvuqDY0tY5u9Vsy/JkTDt9/Z7PT0N
sDkFCMZTCxl8ubQxwOJaUB/zli25cddilb1LKwUpziyKa0f8agPvsrUF2OLZZ1K4G7xly32f+qjC
7quvcAnl3At+QTP+IqEVLqLNUwwcHs4zTja5ZG5GfmO0dlbs7vLgDT3AjPcpjN/wi74OlweFs9er
XoaabK7hfAdzH1OEN+iSI2DsIHGYXn8qIxab7T9g2BCsy7Nj9sJ3xzPfeSLlpbLgPvB3dTry6bi+
2YGmiD7Rt/YbBgJFtPFhRlGZjFHLkDSMOGQe/ZL/ORdIKYVx7Cf9j81BVUoapIPytVsiiOby4a8k
CkUGIsn+dyEkIm6yhubvuJJsIjyKcdjaDIc+gzQu5UHfwUaENUIwKplc6zJR4BFmecHo1THHIKeV
/FtLqiG5iO4sOfJz11jCrHJd8Oe3ovu38XXIXnWE2Ih/M/ckwkH9+IxzKrqKwfjRVrgkkJCllFuX
qWoXyGVPwH2LN6K/Q+1d7BXrMHCz05oOyYqXARwR0e+n4mwY2E7A+oEyPof6lXVzxbJYI8+dINXC
L5s86Vq46Am03l1Hs7LHXtVDqwqUgcGyzLFU+FcrXgqA+ojgDnbTErrBgt3kLw1L0wW9cNTOJJ7R
wq6omEY6QsYR5bMYaW2o629a04KJLzvdEf9HJjS6fmDt/nauzS4SWVqoOgki3j4HN4QK8JMJr4Bv
XLhQlZFpy9oAxexBWk2A2NVXfx/MwXoI4xfQaCa+Jzq2/4bwcrgY4waeieEbw9q6H1ROX9qqUy3o
v/ZJ23Unt0vLVlA6vLRsRbNNV4mrtp73KKP8iuIpBlsidtJsR15R0cnlVROWTaS2VxiApKEHUf0e
9Rl1xhRl0pvc+GZ6lO3ZX3qFrz4v+Z7ToP3co1vR0E5/aaE0cGbameOWDSMyJ0PX/nsnYuA6mgWf
k4fiKIBeiMnrTpHPbg3wnNGVkEXTBit4UyUGpWUECo43QvRTTQu3wRIjlIN3jaFxAYmEh/Jnu/fu
+F//XosVkP6G4Kqe2lIUckI5pT58+bACUlxsg8nWSqMMygu3aAH7BEweIbFowOPuiP0namPRgmhp
Vd1Abegto4c4NvjemCFdC72CKS6VBssYC1rbaK5z0kvEqBIGu5j0J/5uP2TRHWJ/GIMWGUXTY7Yp
RaBNV1TvzNwhz5Y3KytXvmdE3bUb0pTOXYyTWXkQXsZ69VxaDBVNk8Oz+sKG4MqJOuL6zF50KHNW
Xuzzf108vmcidLlYqE4oZzx5CfGPwMepLb7joPQZXPuSWkN7w8PBwvzp71wwnvKCyuyBgrwxpIGG
mI1zgb1mbINLooeUfpTYDvbfU2gnfq53uBJ5q5C+MM++Lye2rIYMcj3OJzABu9CBMS1a5iRvRfc2
QV+6kaMnIW04098JGA/MkTSFOGienH1+bSLfIrmob1AsGKvdBRn7qXmzW8ODvdvZ2qvQdWPvtXvI
Tie9PZFzPfFCFB5ea5aTkyXff2G+yVFki0LrthQADyuR7/AnCVavxmZH/IMIzHu98S7sjRu1im2D
QK2bBDkRchKkDdVrcrFsOD1kPm0cHVKjlVbSwR7AYzArZ38MkkWR88tWbGNctlfBYRCP9wnOnW4O
IMJkVnJkDIYvgyKZR7P/NrSOgmNwCRI7IpgfQf33pbZhtufp+z2jqAmA4Z9zJT5ymTMo4Nz1BRHN
M7tJlXHhCYxNj7PJClxMXSkIFBLYfJFTh0P3j+qbiAIsLlMko1vsXVJc9A4LKZ0cCl4fM6pAufXH
1Dafpg7llXF0bYQ/iR328NfRc5S3xkbT6VOwNUpgLkS03+Gy1ND5dkZUNzA4aplYSzoluzJtEGpz
aKJlg8tobed/yHySuMZwcUhEEXoRPWANF7GCUCAmZXdMO03vy72gz70tRt3i3xSGIPSWcmWDimT4
74SESREKFWnchArBRDukdlARJr8TcS1kU9gXMvpN9TEhsyrG0mN+ooMjJL1Jf8iI6hDles/o3UPG
hKh9PyjUnQamh2nFoYmroXulEJnVUbdrC3wVoKvsYHD/9g3S/31wNnJoSwBlLInpFYtsj6GyS/Xi
N47E+Y4XizWsNXY0BQv8/GvgyosXbPRqGy/d6teC2fjR5dUwN1sKsxPiEavd3RiZ6nwJFZ1dzTWB
d7v/yHFexLxU9BuzBTNUXSSdt1crjpyqRgOhJAcItfjeEz5QPRb7Ey66KeAhQU98n3fVDQdxF2vz
Vk2YfcYTeXC49Qm71vLgFRAHL6+aK1DldUo4yyLRrenuqWzTtvw7Jh+X6WKsZAbwy/+9j2hvCv4v
wKjHM3Tippx10fzPJaMSJ/1bB2ETqYMby2BZETDcwwCGMtOYEGrCD7+2giwx4LvsoO3dcKOyH6V0
yf2ARLwunzf25q+MQlUlpAhKM+0+8rhdPpQbzrNjUdYlI2P/V/vG5Jz8t4P6MA2f/KB+2klZKLNI
txxagpHMCAL+miqoFvB4EjzZDF8e+awpx6M2mpLyLyse/5CroGQcWuIDr4U3/7+pS9SAY/xVs29u
TfPiLch4QLuKn+oxiEBSSBL+dx0nMT8moONOrJg/2rO8WFvosoetavR8rC22ikDm82z+I7LhmciS
qAyhRMxfeURyHyGBhNcYnNyhOOTjnXNuNtTS6ROQRNAZEA9ZlbjL/Y27BkeHcVGmKanwVG2sohM2
cB5KHnXmc1O6hp6uWmv6NoJrmgKNSjg5Y3+1j3E9IdS++Jazd6CWQyu3rpwatWQ4OzmVnaku6Wyi
+VnAJVH47BsWA6fJGe2yvtFkZe2U8F4IKeoa9dYw+PNSk2zcixydyr3JNER3+9ilkHB5eoV7mFE3
Y9rUpRFOI2z1p7JPL1ywazUUWLkMPyZcfLHOkNjp0AzS2XdAiVnQy8tQPt8B6qYe/A6JMwFvFVIU
P7ZrEeW/yHsGTOjkAnWJEekBzabWkwmpcgdg0RBMUi+vJ/x2YVoAlEZqSspacSk9QqlS65TlW/XX
ZTlPNfXQ1TA+gQ8AVjI7I7T8DfOG41q3V5CafpCBEl9MklvcF37KSJFwO+ntJLRQMULqWi/Q1vJ1
uExMtUBMn8Z1YAhk6ouK5lk7txiElfE84VVcLMKzI70A/iZGZwHISRXfn7x3s8pX9bt1a++syEQ/
rSpyW6hWavvqQe/64Vu8QW6z1RD22IQWgM5QV3nmiBHXZKMrz+NOZJMyGDi9qM4RyhQFUwyvpIgn
2FkMnnepSmbEp0s4FEwATMeW22MEiQNEdSRsgYxzGEqgjA6OzJl0j2qS6AJdOoEG+tBUlVTHOH9v
w2nTtoxX8RlajHLt5KKPvxfv4ou3l+RRZpr1r2jWasy+xlVnbz/IP/M9lEpzM/o95C4hD4UQ5pWS
KQOq+K6PhP9YKt5Mc/oA4Aum9yc/3BrV6ib2nXbp2UFUBZRBSPxXzZRnArdkw87Va3M7Zct5zehl
5YU8l6UwGKN8b91h9jsJrQakPWVjMCashEHBmPTYG2wpWl47Xd9AG/gFgnUSef9dRiYVw2MibruT
tFlCdv2PNqxdpsEwuJ7tGK1nrsBQ0CsQ7Z/ALkQJCgxUzY7YdBzjjt2e040kfvADS6WSrAKFbkcc
oniWe26U+HKG78ZKf2iv6pj7tLV1kb5IPGhNd46aaUL2bRRDLMD22GG35S8pAqTnBBLr3ci76aY4
vVeikr6N5dpHzfR5q3nzL0ylJ97ZyVk9gPjSvHa8TsgajH9eZFuM8NAC0e1Jwmh0z8Ybq299S7JA
CNljCATF7yXQcBvtyR0VzPXNUstpTv3qhGvLde47TBIkL0p+6MUgePXN0tfjreWjpyfWaG9Iyv9o
B7cFF2aSPLoNdm/KMOOrNhbGnsVyutPHfAF0/vO6mWwGix7uYKRp7hRXUhV+t41aQDR/hoc+uhqW
VcXaFvNt3eAhw2Dgo2yAi9la79WMBbLCyaoCbc45sl5XSClSn6DZVxALFVgRuENOgVmlo0hL2xOp
KFknH4MrF+xjafDTI1fnSEjzaq1Tgtly3cw3z5VgZHSguQmR6JIyNhwTL00wRE3umMryFHNjwO5c
8pK0UJoDe6QG/mwsKdrlgkSSDrHrfe9ZFx4R+CfJSy6SJr7KwbUvVisr5cnDZIOMLTWHCujFpNtY
yYxqJxMHcbMFATNiZEzfwBs06m3V//jw7Y5BUA7FzztwBtJ7/Nr5QkdFYhkkIULSFrH4UyRtn7b7
YLLMUVFAlXfmAcTL932/TnGX16O3wf59kHfzrTMk/8AevXtoLC8x8DUqoR33wTA/FLmP41rEwITG
HccOnl21XrNtQJNCUGBVHuiDOPHMzlnj7mKOgOAtkblh8qB1U6r9TXpbGwS4fVnqK1P5GCKU9zh0
EdEpBxYKOUkrkP38eQtzOSf7FeggkiO8Fj0CKHp2fl+gCOhJP74UYPxsCw/m4IoZoHqcfQJCft9J
f4Hk83wLo8TYNiOmTi0U6yVhveqR5zvJmhwfe3VZi0QPzd4V5JvGvw4KKfgB2mO9qZ7KheEluVj+
j9+JTMdF9OyhJRFJ7TgxwIac3KkC2qzF/Im5N3A4MR0vYk966kfkRIlQQf7RC8delBOV26cAVdlM
uxqkEykXgapgK4ITgqxxpZE+H1P08DaMMjs/0jXbp3sMOFhTECD3olajjKrFSr/w/FdBs8ZAE9bJ
SeMYc61XaPh9z4Ki7Pi88jXwSOf1hS9LcrTMe0W1x2aPr0qxdqKZ4WvVmHZlf923x6N/3v3K7jKj
rFKMzxEHPLAo1Y/h360llKVlTX8s/vpC44GoDQtHUdhKqn/MkZzGZuUlWMjiaytdG5IlQVIZD+8q
3yj0liXh4Wmcf96ASN1/ofwoTNuQAtq70eXgtQWB6lSYWdsnSgjn3R1P99W9QPMbfBev9vJif57I
XVmUUIqm2WK1FpphwqraGRkMVeJlRPInRVKhhL9SGCR0X2adSjvfLiKLcnx+HaAkUFH7iHKhvABc
FuxYGXO2wyl8toQxI4+dHCtS7NdvrlvzDYCawMS9C0/5zNchjhXjEBSAfor0vYZUo9y120ratIL+
YiShD4H+GNztXFCMcySl3oBYZPSt/BzdckplieTwgdt4B7QkbaUxYD9YE/veBj1tp83E07Zx0rWe
kyKAmSmpBIY9JGpndDn4c9i0WCsCOD2VftQsbKevela35yYz72/RlRbg/BTbnqZ+cBAE84kdQ2a6
uWfr20nc7TMdArTakzdknWANmnV4vOijnM2pmnq6+z9BNuYThQFjoTu4j17X0gwrUnzgxI0KWcaN
YhsRxJ9oWRZ70ITZru7GGYzSsfIhqSM7C/rdwhJLOwaz/uI+z1cNjLYRnUEuJT8mh3atkDuki9Ml
BTupvWybxvr4sr1q/VdzD+q8LMOvc4ynU9ebPMf9VenhrZ5M20qHEn6kV5b2mNEINZYstu/BaDZa
mDzcEuDoS9qxh7FOcThNWKoJRCkHPThwvsjjOb0AKVM7YK5XxJCjDa9knIxLab6ZOIdUvacyEW1h
E3acMnof3c2ogiXLl/p/affzHx2gHfSR7QuQaexHpOFLzICIVhEk7SQzaU1zkxd2tpyJT3ddf/jS
uIkWZqK7k7JhnSs4XgeORNUWvHG5sQwDD7gJLZucrnQbuCwSpC9LV+tTlkStZr/A2ArPUpQ2ALXx
CPEZDj22rZxDlIS5lMrSz/V9IyUIPa0KKr5DGiAjskvUs6F61kvs68ZN6/JtPMTwaFEfvDaiEKtq
W+WGM0iAtAO6zTGOex94G7k8m3A9oBtidwvo4yr+XQZN7izrO8yP3dpO4k5sgmk9OOT/9K1VNyHJ
dPZubSxvO+DFdJ8TYGLXwHVsFUTGbWIvhZbjM3abo+T5cwTyr8zJRvLJyJbBP/9gv8IqbjnrGLK2
6JUaQP10LCggBrQCbN9L0MhDrq8qf/kUYWlKHMxIChKfkfxg0cXwe+Uktn7l8+Nm/QUo/BSMjxkr
61fUZJWOeXBB/ga6Mb80mqx4PC0Aql7mwZ472aFwc+/ctfqPxtAI2VMcnD1oO0q4yYYIsXa2TwTN
SBNsT3jYaImugpDPIE958uKS1/FhypRvDb0//HpR918aRrs9bRqf+Wyb2HK0PsLB+dw2aZiIrZsA
Ba/955/DfkD6U6SmfaRxcgaap3GDXMtsNXsOw5vaLVeGo+xOIJxOqPm6cIMnrBnnZuBZeMObS7is
+6FgftvfPG72WhFyGBiPjwmWjOXpLv9uaUdhzIf53Yr93mHqyLcvp/JVES0xbKNWxluf3Brh0Oln
u1WktCUfnCDJxJnLDs6yCzKc3A+QZjkAcY+YeYeO+y9rwbF3SbNq3k8b6qYNhhd6Oi5TYt4O55D4
bEXIVK7YbD6Xi8lqCItKRAv89DSU2DPNX7vlSwE/F3nLV/5otK7vxN+zkZ9jf3zYF0VsBPnDvYxf
JBPgL4fVoFHQehgnghr7SC6stNDlP1j1nXAeyq3A4zzBXuhx+ABjSgaiHwTjdCNW0MysMAmEmicK
1Btf5YdH83+CuvzUKnZHZ352ZpWedr6i5k3lfJ4cmCm3A2Ii1aFEEdlaN/pD2RfThGwXT5ldXStn
ybmcZQYAh786bqWiggoX8B+yrncSlGh2TJh9LxFFbp8sc9AgVS9qi8vh7MOBGK4zCocm+DFMQQfF
greFProNvr4mRbiPXDh2zHn63Hzycmc1G2l0IP0fzYStlD842q2ZLq4o5/M4C+msIRLZfyKOGebL
/72SjnI7I0hc+veJSxyVBumSRS6YSzHAsdmdODIQTEWYCnU8329MbkqswgSsXqER5Hh7B5sZQvml
93lWGsqPrCBSvHrtnwBFReMfOS4tIs4sHwOgiMW3+OY1F0X3POrMwN4RuYAWQ+3x80/ZhhLaOU12
RG/C9UfaNDZvjXK/5tYsuKZvb39CP/MgiEcNkwoOL5QdxXsNuV6ZlTMigp8cYvU5N4XI3TdK6y7G
/Ah52gHluzDiQ2xm9ZhKnou9gaX1XxeErcvax+W9AVBIDfL5ubpjUtxEfneyLU3cEtApIbwUTiWn
aCkE1MztWa3K25iR5A77fiZLu9aNA40ZbrBpRqczzmwe4fYHRmMVIvyDFgokJjvUFui0gaFlcWf3
DcGUHtrlSNe8kyLp6nPoJnMX3w6i8gn1lx2iGza0ELvhEb4AyuUzdLKkPYx07yPE2zLdoOKdJEZn
KBUKLgv5QPRs4GS5dSsLGbCBiXa0eFBMdZ2j/hXPedlFCJXSNDlTH5admXVJAt5kOYvl4G19ngZe
M8kFB1tqieVGzf4AjD5KRhyctPP+xC+VvGqSmnmZTa38kQGWSpWuDKTlzBbL/4gitg8079IJEOaY
vkI6E8y2Xxf6i62uBWpb0fxvjiLA2+bf3bOkY1+tM4BNDcy+jXX8+mKex3LDEgDiSldZEOAU1Ely
A/pYMzHZvzzlInE61TfyfWhG8gmJrwOHjHooU6FrwpwCiFnjARHqpy5DcBXvAAh8pZkJ5/oQQ+bT
vbZbUohN1jyZVuA1j8P1/d4WcNyzL0L73LJr6oPJjbD1s1VJht7eS4LY9u5j1jj2Ugu/cw/DCeCF
ZPTxSblVrSid3r/bGB+5gJEioMidlrJpwPJjcdfsMHbsmRzQfWIPSucqg+HJSJYsaJr/owvSox5W
GdipCyLDqY24RNcxdM5oR4177thviDnmOGLy+YWYo5unFDKGYjtq9FeizKrTOXYcXqxTNYRgSYBU
dTiT9HU+uShJ9xczwEHN8JkyEJfaLM4OPZe42aTkbwXDU9Fchxu830Isy9Chsh7dX4sWsNKuLCXr
gy4oPabxNJFHC5dUdE77/XxomjNtC4NXKO8KAT1PVkgPHbefRe32846Gto35SOBRYufx5Kn+6d8m
VmaYk0drRkBty+LSBo7gafdC4GqbDUuGjKlxof/eKLIwfLKdsWuKMtqMNgdHTznHZpjZXV4NdMi4
a0q/ByEClD+Sf+fuinz78AUOX8lBlOBW187oLniHG0mYGEKIg3W5aNxixwAXh0xlHqdn4ICx58SW
3H9gcW73+WvPEW44GNDa7gSNxj0Sf7cb646rSe49FD8sQoPJz2NR7KNr4p3qF13z7jH9GkxuuIfv
TLzmguQ++n61tS97c5gQ2XkHUpV2JPazjvTxaSGUam3qRhfHZ09yzq82euDWyZuT0+aD+qVedq5n
VYEGvEQGN4wKLxGRDrc9B2ajUQGr/JZRecwn0ZwCcq3YypwkFVLB49w8fHzmEpgFVMINCPEMGCK0
ylkrsgE7Kl1dyIkaG39ikJsBglS7wca6CQv4Ckahk9uO+IRy2F8hqLxrG29DBTDtA1eRmw6ws8Jg
L8byholMbhGJDlAC2mDnwczfU8x13USuWtYfc1LsArAb0gVnV7gTm6H1RL6qaAN8E2IhJF8OjQTK
CPgvgTjeJSFJ6IyZRqZ3dEeM0aRMnstFbC22cD32jsO8X+q1k/p+pjC2GXVu/TiQERqUs5jV2gzQ
4S1aXQewmo8tQY0FBN2ssyC7IJyQYUjZOE6cYC++PkX1rHYulQj1bHKsoiY8ZxgxZu8kY6/TLRdJ
HGQYM3X1iu1K4p+UNT3tWnffukR/dM46bj3C32DtpsFcjjroG5r38xJ5GpSO7SzmV7PxlQ3oPvGz
GU6LiISxQZxpIlNbBnUhoVI59ftHVbtfVp2gHKBvgmLF6+v1tobZSTSaYO9ZNJBJHwPY+i02mFGT
jwVrJgQQOei6h+baYp2/uNRhfU09MRXxN5b/EhiqkL2IPawvOjc8F8xgyVLfEqIVXOpNm9DSrrOa
Hh50gUKT2nWYqySsdNRRwQUB5sJNNZvdKqsS+1EZHAPfquGqAD/Zhrt1UiEScxSD3E9cpDa/xUwo
IdgMZ/WYARBBzb2n1ZtqD8A/Uu5R8bhOqTI9SvfM9uNmK39N7RjIOthpH3phuPiBCv+bP/CWkppK
BfuNokHX6hcakLTerFiTo5cWR2WHf8BcDhMDdJsn66rwpOtK4us7mzMA5DRU7RW/kGRYtdDO9rNY
6YkM6ZJm6IAmr3gX6mEPg2u6zsDVdIor43sltf2udkyCTCiFIlPHSTJWgVdVQyQGWF7uJkOSCH5q
pwrKAN1ZNaRJRIbKh2ALb8szE1Dn2MBEBxAdRLtbSm8Y/m5lp0hWuOKFHgqLqhzHHSNyhlYmKVBu
pP+raZdoEmJ4EtmubP/GMtJh/DXNZKbuRnA8RVPeHYnqtGpBoi3f0PWhTEPHTzcgQy69vW9HPxMm
CVpcctgOCm/YcsRxbYhdRgLcsaaP9m6fOVpelPcTqnxK3uQdrmM6epzx5EUEt2MFiB2WI5XxDeWa
5Lj4Q4/uY1Cblv+xG/yj9uMo2MiuCIWl7piNYKMJPHANASpWi20bydSbLQvjmFsPFAIzKX7jO16H
Uu5JEwsApKeUDDTl+ajTjHxJVEBj5qj++S7OuaTiO/GEgyP2iZia8TT2lMrEP8Lf/qn6AGGuT1rC
ETFcba3hJmUMSCRxb9KNolriQ3HVOnkIaAVOoEszYtL8HsXeFTvmE0jD3GUvHXeVw4+b4/Pp0O0s
t9MmOgi0O/ss++igjZ07mr/z5C7edrX8SsoSZAQEV3u1vuBzNQVO5Mb0wJXoLZGdpjFP+aa8F4hu
UaduS9+RU8buZBhb94gVDJf6osNvglsAKsrcc7nZRN0xdKdLdDQ2Jzd7gIlAHF/zqS+WRewKAHxd
ZknYuSpN5jfYF7WJFzyTXx+N50hr+Az+KJQWkh/ieTPUx0MIVHpxZA8wmzy8+ckkwU6n1ClOTIk9
qq5225WpMmj0iZrVsZSUvDotpQwiEMTOHST7+6WqeMLlrnBXwBNddF4w3YVoWdO5hfj89Bag1A6Q
VdmKaSkkwiC2NDhsCJHTGZbsJGeCqIJJekRjzfpgpF5yEyxER1UvKi93KT9XJpe2C6svCsWPTtso
5IDTO3Iwxgq4vwrAAM2rfQhtiL+MbGQ4YbVUVwBZaxQpr0/DSq3nQOD+iNyak15VoIlCBLZcd6jn
S5HirYMY37v/W5USbxAtw/SiwSmKiePjyxSHJywpSKiKXJU9Ip+wEOu1Ml0UolzQmCe+UYh/Fzsr
Ihmb7hiMKxy5HenClazlGOCjHDVkEfuvBCSJn6vrQwzFvTrR9oc1GB2lwtHzP0UnVkbq6edz3pzg
5PmJy4ne8NDt/49NGVSX+VdlmW9tNC9zkp/dbzt2ObplVKkuqUgFnkdAyX0yL8OjFv0+y05qG70l
KmzeGAtlYq+6gsV1r3v39wHcRtT0Rpyo/HZ7TnqIf+TqTozPkFEGkJcRqT63w2tfp0cNLGtDFIdt
gIvL/hIr6wu8ZdWYgdm6HO/EW/ottqf5T5s5SO6UnuJeut4GBL0GxlZ3iqXR8ztsJP67E5odJwwL
TNluf071386uXYK8EWezKpucZz2ZJq/c4BbiTW/ntSWZZX1IDYWQ6tgxgvje2Ggg3Czxz/0DPdde
/eaXgfAPy/tb/izZ0XntqJSlEcQfaS0e7HUS1DGokza0IFvJp4x4sTsveO6Tk1BDdvawxaSmRiIB
hA4nZy6v+dlZv+gnJuC6LE8fwpydfaG4T1+nBR2MwwEK1s2bGUpCsIJBnae7XjjdFy67c/s0qdqs
lWWRNtySPOUi692B2o0W9bMlJjYP2phD5/5k+m+QSXodUiSLLwcy2ex7agWlcDkNJj+vzVxfB/Tp
Wny/kCnRbTKWYwXXXYOvKc5xNO53sw0odk5cNTDYOyNcC73s0YPeyWYdLXHZUSfp78rLpnChPSCA
nOQWOk3Dt3kB5pyHhhzOpljMwGU/tS5qrrju/97ALtZzBtNEA/B1WDpx3p1vOhXjfMUN8MQUIDQp
tL7++uYExW1c4iWkyDa9OuNAiIIW/jnL/Tb/6kA6PEqciCGU/R+gJOyb9kyitWe4CPpMr3yEbmpf
BNCqvS6Htzsq39SaqKyvqwVtC9xiYQouS68oTVcwyF+4abbnjDr8OxPYGjlf65rb0j7636YQRhC4
tiUDLPQMTSqvTsgy8xY4k7JiZBO0AdRjthz/jIqE0E7noYiWd/sJmsUHD3wfWwFOAWRIQEB7YKhh
Jcpnpgtwe66C+a5B/X6tCNdYBwx0wCgtJqitahByrHVPHMNmPMDGPl0T30jyTp/euGp4INvJMwBi
n0ACP3b73xhDHu8F70x/y/Mof2/AQtykFHMu/40NQxl4yk3QotLkl8UFam7t2/iEPvEbeof6m0g3
obsLODMKYGSFLKNeUezODOsCn788PYh+UuOE1kjpbuprXCatKZzsxIBdG/uyUVfAU14IH80nKYTm
B72w3tGaQDpftREr8mXwARMEAnDV8PGic+T9E3nCPPHWyMGJg3vN68zcHgEpHIojSuHRTYd74ZMT
mwDlkouUosuD5bt31K5b0rO26voo5cj3/Y7rjKWLaKgTa6t2etCovYxChT8BHcXii0y8EzZGETEJ
97K/UsJtkrXwktkiB0BWLFDbrw7zqcAHDopeMVK8QxMxgtzX7AcskhRfkBJ5dtKyWL91MBAZxCJh
4BELPjqaOpjgbiI5/Dg4WZnbGmJ5rGi+yK+WAzvFzaB2hxemL+49nalhZIuAkU8S137HEpV5e3qw
eHFgrkRsOtFc2UG6etT8gg3lUMkal8O2dLINhak7faoKpw/J6/tL3PQ4rHPNmtIkGxEc7UOoWiLr
45nm0PdN4Pk5KPiDbX/O28M2EtYuLnUGsrg5VEeRws2PlymW2DJFJiQGme8c+xOVaDhIGlMpOzWw
lrGa/Pf3EMnMTPllirQ0BRaCuWuLeLV1MVCz+kwV9YolorZF+U5CbA0PEQUOe/So461zVYLeq/7H
cD3VNyNidTHy0yqHBLWhIHCW2SbZWVYsLa3elNJeIHxrurUh3DID1wUZkZHREggH6U9J4Zx4ECB/
VaQjgS3xjA4lppVnfnwibbQGqE+w6WNb/HGIS0FxHlQiftdt9VzfKTXhHR+knwAsbwd5/O+/it/w
ilrVv1uqAx+8/QlEU6LgZTAWQIKB8k2rCHx68aQtlcs58h4WzM17k/FPx89SK1PDs1bL4HhXT/Ub
L+RrXf4Ki4DvnCY9ocw8PG8iDDDPHhtLVNwBSor/TfElWWVWEx1GQntJhcDvCet3LRaQIIzKm8TF
aSsGsuHhJ5PiKUL1Vem9C0N5B5hpgB5t0S0x/m67XonQJ9MiuIWi+rq5Sl2sFpY2VpP7ybnj2l/V
IOUie0abjinng2AeSH/VZLZrQxcfxWuFQAYhte0rCglS8uZ0FNYqfhAHg9MYTgLM1/BToOuK7ROD
sJhQkGfs0oJosbLXFkwN9KgBzDReXXI8b7Hi2ld9gUwTiHUZnJE6PmV/hm0F2TTw7s3Q4HH6/xtw
ZlsiImxtJCnFqGhgPQROvUxHIycfMCSPB2ubiHR/m4x6XMA6CD8ER5WgGMYF1PdYVpgaCO0tzGoT
r8z2bSJjaUeizRwv0DfZ2b03PIAVQJe6WvW5wo2Ls2U/xVZsXnJSA2OTKV2quWqDWUAgU1rSoj++
LW9/COuZqdmeZzSe0hrXlFZLRs+jqg8HMqfdDQcNzYhr36w94sp9wINX/YZ39mkC2A6epzABOYNG
hxsuYd8ld4QFpz6G1qEZOYmdMMXrYCxzCZEfhGBb050J9usMk1VSpl2sPzbjWxBPJ4oXQjdbsUKz
BZzp45O89MEGKOL95b5rbRPKxAnXJT8vm8omOvRaj+0IGOSA3c86MtMikLSCwpTUK0V+trZNDsF8
jbDw0p4JzDZt1o+GcZ8TYoMXSlPSlAJ4JkEbikLMv1swiXGm0ZR2c5z8Zpw/T28tc6T18rgpqA06
pGAZaU7ZVVuJLldq+Ylcq4NLXkf/8Eyr8SBoLE211G8jeHaNSDkuAjBqIVrXvbsRiHX6R5fQawKr
y0IwB7gh4e1yDbBUuEj4qgTWl/bZdD6drijPmmeNTR6dL9KhCVVepJBTX/YDzFEIZmlgAMB0G/K2
KEZU65yIwpM/W6CrF+xQjNKtVEUAkLUlhiedNc64sLlK9v+gvNW5w1NyGy6tmPrm1mam1Q1kn5R/
7egVlrGt091mZI0P80zUb3CfWptGEtTFBZhi3323FzXkvlQd/LpI3c+LyszsMHiSrgqjidLWrvOb
xEiclpQ4QalaVcHXFBrLX7XLwnroqVWgFdg0toNCXF9SX6Lqy6aPRYugUkeTWpA1AA0msLZQpsnI
n+ak5WQ0q/CuwWyknM086lcg0dkitj4Bt4mfKfl/5tb/MvMoXftlEBCydZ3SgyjD7yNkHD8jQ4Ix
2smlTmfcAtmBQQuwgA36h1nIwi859/OmjofI8ghI787nZUsePI9TgsRh76yG013Ikaun4jX4WAuq
+NTxI03D9dVbATX5SEVUxzxDKxcFmFQi8wlVNfviQ+raICoTZXZEcpGMy4fob/Fj4NBZHWYGbNa5
OV3rqck+qqvroaneAg/kP6RDPkcdcT/zrU7hcGBdBvA6lhbpxDw01V7Rx/GurllHtL5K9hCE1JrJ
GMJOY7xWHY+SZUE9AGrIcRg5QBsPWA0V7kfujG+IF2baJ+8uDZS96AARepx/5BRcxYoqvA4nJcyI
FKKJdZATuhCKCN6vo84ekXR+nUATTPFraIkoH5QeJblOPkBbnV7Beh+YZrhn7z+iGS5Ke3tO0r47
/WStBM1OD7rvldNRoYFrKvv+xt9tki8H+3xO4y/ypi89N82eXRkHcjiCh81ErE5fpzG0H2Yi6bvx
yqCF7BKMd2taipSlm+3Ib0U5EGvxVTSANFi99aiErnP5ZRqXbET8tdazLxncjizQh0CJFC3nhEmg
xoQ+rEcI1T8VOs30aPD1DS6lloU62DVL0IcESdDKP7XO1BE6vBCnDPty+0BH7xi0XNSv33+/8lck
jgQ7vjnhWom8sF9KKD65XwGvKNqDQ7GMkR+SM59voEn9HvbPsTRzBtOOtU4CX7fXfQGW06pZ1hPN
mTg9IunRdpCAh51szpUQIeUgH7iWyl9QEcuD9L/CpmGJLskxPeo3r51WRYb2P+D2mfHBuNV5Y0Br
htxc3w16iM8PybbnpLC2cDQu4AaRFBhObqarnZ8J0vTU7h8NvZOTJftPXPJZDBsM0GhqeGYylyje
L38cypBw6KZER5jbWX6vWZKtCuA0ODy1cFO0bMGH9LfZYraN0xhGy705V/iQRs45ZGQ72njvxrtu
rFysJUm15LHnU0M+eJXOP+gAzFPqn2wQD3VNpLuSpXmzAQwPV9to/yXhCiV2KDsqpg7JFrWfBPtr
69TrlvBU3b6lRUrLCaoScjJoJPMhiicfE3Lf2j24kQYLcE93bvLu5rdiVcdD5dWxALT/PTJQTpP1
JgBbVDhfMuUvSvl0z+XAKnqnTt1hMckvDIJ0bhYnfaIihs9rGGzPzP9b3twJM4Zxh1hRSXEyXIwI
1+2sTMBw55uvjmJyqB+CvIQ5hcmzCw4CPkfwYZt66jjiCLNxflovM+R0i755E9+QcIQyX3lbID91
amTABzZHR3tMOhFDffS8+uzEJargHY1JKuP0U+JbIlj8BRm4Uojx3enUMLzwqM2vhrbVtbWwsu+N
ZgnCma8P377Vpa0chCdFEuOjEtQz0sLa1egRrTECYd7+oZX1+/GiygvCMPff4CPVDys5W+Z/ZWNQ
8rtyKmkkhvrzxf8193RGwoetfhyWzXrRPI75DJDTG/zXuNCcinBSoBdQ8QBi631M5D2Di89ltL2F
BwvN44RzNsmYSzkVpCqy4w19H4VCiuoUiK2HkzOrnzLRTF9cZhcASnAMsTG/VPXIacxH/ATF1453
+TMkL1Zu5Cw+ibof8aXQhGWTjluPep6mHhMyyrC14Mx69R8JWhF9412rZYOC4OvUMHIL41Lsnl17
XbSDiW+82/glYlGjZRnKyzImKZKhPShzxZgAzqRC2kFsR9dvGkMi/82ckIdotiN3IdUyGxP49MES
XnGNz2pVdwW7XNXQat8gi9fSJjUEbOs0CD4FFtsbkRmv5Od4OewYEFmyyNiPOmWA20/iwiMhCbki
dZUcCzzfL5bc0ck7lnCGLsgfcGnWNzglUty328NU67F3k4d79MQZFTgcofBRQff3GApgxLZZaKRR
0Mip1f9QEK0VW+Vfsccjgng2VIJhdQ4NB8tC5dZksicZgfWBYhX3Gh8miCqlnsfQooe3aNOMhrao
OIRx7wA8CZIduPw1+2kbyPGWnn/jASidcr02w/HAGktaPlk+4un14tIFVZEFEP8ZIdqxbeuvHitT
nye4do819+XfQejqAlRjYccN8pMONU63qZFbAqDp2RTxUMEcOBwqveKt7H+W3E4K9CYW8L0HoFJO
llxZoWWRBVkMiFT1TwZiyiCb6iyB6ZATW8NqPx5PF0mjX1zB4MPDF1TdBYzXTdj5ZW4/aYFiEN7X
sN0v1vCWu+784J9jraa6/7o52aZE7lR0CrosAOx0wyUlQDw0MzAZbjuqCwDY7w1VnFWOQqgaS3RP
lBiOAstcCKiUeFlvMp06aHPr6Zd8ljxqs9zeiagk/27V3eip7X0zHhfLTO7r/gB58xLjsRkIxkvY
7Ge6fpN+WGdEBmUyn2Oo0Fm1kqmrM6ix/hLdyqzet9qpwQnRl0ku0opAoKaFnLcMOBqdC6KmnkCZ
h6yFSWgF0SdOJB3YC1g26KvoXmKwim22OUfWw8xBYBt/aVUJTjkLV8rDLp61QdcJZ3mY+ZOOGlPD
OHci5UDzUitwva8V8oEh03VVqHIIQFySemN2rfdYR4k8xZ2uM8ehP7uDW+qXDrvVD3QlQFtTvctG
ZtF0XhCkvdgNRRoZlMmFYn4p/V3+T7Def9DwcGukzTw97/bG60e6nRBTWFNhTDqkmW8E5Ni+sUcg
Y1qdTP9VozspysA0nH0oAQ/e1v13cp0lJXkmRuWaEmwZYMbYEyV6NQrjH83DI5wYg1skWfAF35/O
Ig7ffwAFJX4mrqJX3xEE91E+hyTeKHbz4fRlbkZ8wXf25xHSaCsX58eUr7Bj97a9XJbwmBhu6oQS
fG5+81weFb41JhUhJGGo58ocj0ZV/X30RL1yDB8JpWiM4lR69UZzZPmdbB9iwSdgcoAoW43bn3wd
dzoDhJPbdDap88EHtyfJ69UzVOCdGnV9+KynN5+2LbNWfzBWb6iT7DTqXrR3owzY1dbg9sbJ/qZc
KV/pQTLbal8ROAKOXvSg/myff57Fcroz7ATvv4A7wIPyimxV3X4NsrJWd+FDIcY7oJPG3ROn6irF
PgxE0Q1Rytkm+1Zej6t8r5P2cOaWQyOacj8dSeX1o9yCAoIzVGvgKTgVqWR0UAlLRPQ1KdA4ICLb
Kkxuvt3VAshZiSBHdGHStXVNR/ZJgS4/33BGkupOSQtI1ZNRxuljnbxa9iz4QupSXv9k0zmLWEs4
G2pcZ70IOpVjjkfR6jIRTKJuwB/IoZYy2hUFFJtgRoDvMLAaMPZdUtfKr3ysFgCxVyKw9AHZ3vVi
2P9ShBL+Nh4ApkShoDM+Xv8FDFF68lImLJ9FyDkAaOo1YWTql5NfFC2cObGOxH7Ni9hv4XfJHaHA
IBb0dhB1gEzE7X+fJax8aijRditd5uBY5P8Liz1KkLY1UEe7DAxzLNxxFk3+SqBE9VcDSAjRfPVU
uALZK3JJviEK2IyEMz6Sp1cJ++4onOtoxHNTfuHc2gm7fpyiwwc+k9L6/yrAKaC3UrJDA81et85V
x2/XdX5b+au7fR04h+cEbkkv9kA0At3OLUrfFv+3FkgzGlrfCqsZg83m8Y/UOkRD9fUD0PrKMNx6
djP1Fs8VqBrCM0RrHRF2ShP6ohZYOItgaRO/WfAsw+bxHAjyhn27HT4LYZ6wSbi6ZyqGk5BbelAk
uRNjw2zPjWGAkU04uvA0riO0H/J/wqdc56cD35qWetquhy5sUoQdpNLKz+aw4jDcxHNyY4fAlsJB
tPEyqFReqpBZVAj/EgYStmXYu1b7kZ/mX4o1G2j47oqb19p7t+rtkYvpATZmE5iAPgPuKSnrZqre
5yiQJE0XWMOE0VWoxCoqCP0Z1St5d6YthybG3BEKpXJ640NUYRQ3NfYx5SoS2mNbSPZ4CMPqZ9sZ
UMdV1lxOiBVnfGlsrbuoUplM5uFg5leNnl0PgfB7Oh+4ytLjAOzlB868cMaiEQXhh7iJHZSjjkNc
Cg6dWMY45jUx0Eg7IE7MPHRuj0kTlMK3yvZ4MN3XmyoFvQAFXUQifmvOYtVHyHCWY+6JM3tThg9W
xmGWKfJpTXA6kaBL9Q0wmrRpe3E9oFJ4KtZiPL2bQZD/GrxogYN1MwGm5jeEavKclgR9Bp1/W+ll
rAbowVNdOoOolbDDgEpjfYzuY9gGZdDHExND3ygHIAo7W022CttGZ9lqc6UOZMof8+8qvTZegot6
7B0VOBpJq17E3wJqWLCw5L1KJOjr/t0uXmCQfEHuPcVnXEKPQOwGyI1Oa0PnJ8sqMxcS1eGOTfWd
vmNeUpQOpV1aU07L77TnrIQ8mNpBR54y7vUUg9UKaNkGRR6wAIsPRr8cd3V094aCl69Y909f6k0P
CzW1Ee9fb39od23NjThNWfk/Gj2x33oQROKyCYULUR3sZfMWTuRNxkfM7TMhgkW1m49ddMga7Tep
3P2XX4YPh6iTqXV3nWKV+XXc2q8rCBDwTVYIkWfBmeTI/WKJ/xvtAfkF1ECZmgLGIiIwjcly+7jO
JfUerBLILcZGfsLecVDuP+LIktS9JkhVNeC5RNgmlDlUO91Z6Wg7uhVHxRbkVtBIJSBk7Pv5Vmmz
4d4wKTCmdu7o+a4KdnHPmGdZdfPybDFyFLufICzmUGMxweB5XIdFtAs/AVlL3I/s+FPAXEbqqDil
riXfdcdGOYxsmzMD18BUCrRMWisNOlwkRZ5JowYAAYZFX/GgTBEduz+9onX2uPN2w9INXLWhKTwI
JHxzH4sI6fJm3dnR3ShTt5pJHeK2eMDUMVGbrBS9aFW2EKZ4z8J8nzqSvHBAktujY8YAQg4DyQ0K
EWhlHH9gElLmaTkFiVxFkzVSubJZr9ecAby0a2U4ZwBKWFDizNgIcLdW2mFzqTJ0irQJAiw8m+dm
SHvRnPMkJ+xf3VTVsRxQNOhsQXjFwrt/NqQH+rQeEM0Gu/sqppAjNWbRGKE6pD7AinF/Ivzh80pU
AzAxyBnrOSrxfndUG9Kg+geRdmXZ7zqYjPsDiIE5qwM8epdqeWVU0L6WYAGGDbPJ8PKyIRXipFbI
buf7K0p1cNhUXOvxeBBdl3jCx2t9qARWKl/cdEeGzjD6mdXN3nmwDc51MLmmP8NJngp3jP2gsuyN
w4lrRhSPVnudPIwX8KroApe11HGbkbIxzE8v2sgv8BF9YyGuiF67e2WBDCrdDrsxnwBFhVTngFLL
mqA59XsK7ydkAoDhw5EuX1RanduSIapObAFxKimDYshME3gH8PFDXfVgOVL12Al9Zb7in13BlOTW
hlNPRr6OKk5mmHhqaKSiofS1REDkCtmryW9+Db47PgoMfV5HdSkEvUK2nLX/ntOmtG3XOIWKNDY6
cpIPEh9V2SMyEca6BAmMfwU3HrEaAYIKHhSHKza7ZsHOLo09fju+fcX79EKGaC1WgHY7Oo3UMRmT
7A3noVxt8jUs+X9svL06npsZ0qywMbNhTCcDS60gHlZDqsVIF25b7sl8w0DLE3/NvqmaRIZkpKMd
Op9VNNJSiy0Mo+e5c42iDhG19hKH2OeJfyicNJABelozvuxhcBDOIbkaaaqOF/2T5hLimWfdqvsD
zJZc9lxPWGl8CqW3VwbqY1I3m+dMPtzUF2/CiMZf7w79wLwxUsMH4nY5F6N9qgxpgY4DdEz/GHQI
mW12o4bOKYBdCZ9w4i8UrzNmueDbM0QVEM3vygUhlEEgNt21LNtYcspFpNSetMtIMhnR8TdhC4GC
gb4dUzTOJodz5ZEh3Sx0WajL2TMqTnQf6bxhhlhisARPEiqgZQtbWhNcUZYsLx4V773SvHo4z73I
VyRCPDATBqvkAqX+AS2/eHhMXFyI29Bj9q/pG+6gB81IwnBlzacT9WFNkONbKSyoSjd7quE2heMP
G6seoCG6MwMaLxQ7hfAfbJcNW7v5Zqm459xj88VZuQMQ14ztnTr2tPBBlk7Enitjddgl4MoXdN+2
b5wFdSmVpla4K0JsRTiNx3iawrlhw0pXM8SHoB3mLERrpNOGAqapHtv1VbHeJ462XmlkR/btTopV
RagA3g5OTtj/7jceLbDdSq1WoWWFq2BG6rKksa84mWIk7WWy/rusMyQ5LaU13upb/ECOxJBmfrrD
Hp3nS88PWiqsuv2nvJf9Mo5KDAsGiD8Edz3M3MPzrSx+TCToTeLG61Cs9bESfEBuNQm/XxVQsV5M
XPcsxnZoASZyqqp8LnlJejcbqiuV1aIcyrKVsbpsMw7fH3Q0gZO9SWGwGTRieHr8ll4u4Q1iFQcw
6ppM3H9AbWhjB440B2/CpYGo5L/1LMchXwmjx7vIqHCN/UUCgXbSzkXISvUZVIIpvELz4G3QvxTT
8lq4dI3KDFkob4C7Jom6nShxe8AANw1SNQpVgCMMa0UNvb+hTRscXjV+pFsHMbBxNzckmaFzvWDc
2F/lIJJb7jd6FBU4ltL1LClxLMLHFMXC/8zg0zVegnma8NTfNzcA3eifNVkiMVGnL4DLxQn1kZOi
JDQcyOI3Xe0cZ/Bkk+5F31eYhVi7LKeFoW/UNyMLw3yXj9Gi/3zE7T/UX53iD39OmxaZfZdA0xjX
Zx9aZp/NXDe+L3OJ4jufsMdFTAOO8WeW7rPEsf/VwA+xEYa8uM4CN91zDVuoxmAqMqpwDm2apOgL
Sz3SfwQWc2/v35XyC8VpQEQfgpSamW7uv7OfdpPgISgyXKa5zE4pWxmEJMni2wbK6SlRal164qgH
E5IsyAftzngV1BlXjQ61y6dA6cFsijjt66kjTibj1bh0xUSNNWbKkT9g0l/IzJ82UQyD2x/LWhRi
GNTdAuElwmH3/qcdK+zc1YU7oZGRbLI1nF4mCcRMecDgi4W7pthhhUkhGYQapdwB+g7oPN0T4agL
AOobfo9tOOrFOXz9nzRe7y7z9h63dokyV7eyxj4xZauBnIBMcnGoad3snJwcDmcqI/XkmFzA8+sM
C0n85YCMlO4pIPPivOcNJF0g4apRqV/g3HD2f1xdWk12sYCkv/AKSXfydM4zIKhzZq8t4rzm/st/
Jw+C+Wx8MJoUWyYgR7w91bLGuM6Cq2h4qLup4e9s3e3l+b1fe3QXmP2QeP590fccte1LREHi8jT4
wxIzy/Rh6peTBx7iv+sdzAQbYfsc4Gxg3rjfud9h4c4bkOqGT1ZBCvuK7QT+hwpUrfMXIqFwx7BP
DJkafs5Ms+K9dIpkEdC6jppDZO+Bm8pXC7+NoR31meOzRvIThkXTzqP9yctMWnEFOFSCeEBTfFDZ
LFsWdqUHqgFtqdO9pRViOU6fu0b1kod3I8yvmnX8pQKUfpCgh/AZL4lPVSFCknjI0mpUDBu/RDL+
OdDXEmuMCbNyzwpTEy02AOn9cQsWXq2VVJFwyecGtaqpmQ8igyLtXycYj7ELbjjma5bhF4eZljVQ
6Uj/0KHz2c80Qyc7BrTGG5DimJuF04NJvVVc5M70zTFxT8eHzQy5EvCVX4fOrqw7yeaVGS9QHzUT
9eKBI/ZNpM4yVHULY2t4Okez89QfX5thPhxgB0BdOxj+i4L1J5BTwZM2H7/gjFW97hvVIdaD9BsS
ruWBh1OOwtyLIfP2zkBk5cc/5YLUBJr85RKGIUUF8tFk3xxHN2pVn20NdzAzUgA+Euu0TN/xoGVp
M7bua2Bu+70gCBPiTsFXDF5OGq829gwqx9eIuZlxGKIgyGXMHNN7B+GoOdOt5gzbzrQgtyL97xcS
rZZltK3ICRvsc/ozZpySyBongSgE5VoP1gzsp/0xf7eeaxI5QFDqm6teFO2s3z7grvdmb0zlkK+u
kBWW6zNJyPQhNpv2ziW5uOOkLskRCh4yG1H57yuUHXlZBhBIG3R9geJBzVvlAZ2x4lh5NGYYVZMG
TxTaHyBjZ7w4oca8P5BeYr1hg7g29uo9dHIcUbVjvGXMFJfEdlDJ8ziT08zJXDWX+0AP+f6+BLVz
05L2nLGZ1O+utWSenj+1qhVVajR7sTuJCFA+24ONGnHHpw60x5o0+0DXXeQ3vDSiGEZwzMVLA1Zl
Iax9eUGtIM+V0iYIxx/zJLUUjWVOWzvlgTcl93FXoLd0lrTepPaShVcbPVl9g00PrJwenXbdZ3Ak
3zzkY1CkaaZRnlLMiTW2yZz9YIXjrAKieTIn2OWwzwj1y2N1YZff5+DNrxXI3GTqxpRgnpy2W28A
XugGhcJZ3TRDhSSQAjZgGipve44AwSu8KcQz6eAktgQOe5gFEWqn3OPD0wP8MYdt+zuFnwW40m0A
XDK665Xlw+/WsM3Zoz8qjqaSvCl4POx/WfhtQF7hID2efNm2ZtaFLO0lNcHX/g7ONaucul7PR5J2
Rg6g4iYNq3ovRtKrpNninBLDTQ0I0isS9w0Roj6Y7ItmbB7JURulcU94wzI3GJsgBFOHdQqohqWn
Hg443Joqf4aTvsnPMl9Ngojg+EESM0UGaEpf0PXg3/VEOHTyF14JS78URCJ9XiEIs9M2+bHcv+Al
peERv/EDVxedpy93r4uKZTs5nHoGpxFM5BJxDNDXjp4bcy9NttLYIxyU5h+OOL/hDl+4WrJenBnX
2XsRIwh9kDFSbzx+qPv5mwciCKe+O4S5IStv5CRaVMRyPRMaXsx/qyEimrHODWmDzqKio6SE4GuF
p5u4BpvPivBsu7jvu0qQgdSNEZ/0I0vsZLWE4l1H7tIzmfG3woTZuK2E5eClYSzkY/0IppJI3mSN
ty3uFncoZDwqo52THPRvvZpKe67o6UPPDPrQmVECHoHcyCiPDx9WYdPiZPt6rR3B1MfVmkVh+CUt
G53HxRKYlbIViLyGjlIGiONX8SZr4RybRz6zqmImBWTDYB1JmUIgXLqJaXJMRHJaj+bEZJ+IebdG
uikwpSR6d05NYTZGFXK6QQrX3DRk5ppDAV5xKq/6JP8IhBmeiE4fxipRNTT0wHrOFrDVDn3VmHQ0
zIS80c4QjeNhcBd7LFsCdUT5LNb4wynD40Ux9bibNWKBvvHqQ8/ovG1edpmVf/XQ+NPvT94/Zt42
8slSCSV8aXv3JSk7MAOln038+GEzVhi1ve0OM/ax6dBVxUePF9l2gXuVe9XRCDIjQnLmAz3mlO4F
SidUR7v2ynhpTBmdgFpbjkSqasbi0PrhfONbn+Ehk6MigG4ukS6cF70zkVf/CB4BwP2e2Dtisfa5
n0ZRiJDvb8TMALepmaTK3XNBr5es3eLzZIvJykf2PH1FbnQFV83xA+kqv39sh4p1AHO7htjSkaKP
V3iB49fS/leLCS1ItMUMZkD5PpDBQiBY98Xl3YVsma7AeJFtFe2TwbpIjtsdiFR4b8Ta4tg5b3Wi
a2lysnRd0dFpDmWid6Rw9r+Icmnb4fRJFvwr/x88yUrCZD4p7BnszIMQ+K34RGvck3wi3T8wDAm7
zz8kG37joqlORF8jy6YT3QN1Q+PLWru4nYb0npoAppCG706GzCuy7Ob+N/3TMBwo8ffhZzpY+e/8
/U2QkCFbCeGHsh+xQ4sqq8ZzajtCsTjJYiq0GSu6pONDfqX48WQJZZY5srT89erdhj32v8THc5Gg
1Q3lE5PQ4u3kYOot1ZsrNuIXvmKpEkf7RVnlfYB0qoq7sfUQlUHUOyP5GpftsQ6fjJc8pxUs5O18
JBP992mA9XjLHysfO6q686lzGHCTDk6nxXsGS+9vWaM1bINWkK7ms7pKbNJ+v9c68l/T8fsN3vrU
jQLPQmG7Xz2PhAZcRFhNf8mXiYqZXjU3SQkxboN03WliVabiJLto6FGSHnlefn0GWox5TtTd0q9T
WTLju88nyB61zx2qyxIxSiJ+KR2lFX27zdDFH00e1B9usxJWuTdrp4dTVNp+RV0Muh2VCnnxASxh
QikQAAqqYTA1CcNVEO6hnJRumVXzQpA4QUKViNn2OEF0ejfuUTs/zUmnbw8b47dE3NDTHLMk6xGo
Ag6M49GEuu5Sm+cKWgKBXOnzj+Dn8FKnXqbDFgCPSnxYkt0MO0DeIgQodpxJ2pSW5cRlgdXGxT/v
NDFQNMX0kKjibe6qr7NlO2ksIlsS6XX6ccue/qOMPZXFf44L1hz4mOsH9wfdcNA9eEn8JV44E79d
AZPTBMpn8Ds+kcuIvN9TyGjwkH9oK4ETfTKA71NCDV/6LglrIig5IR93C+QwU/r2z+yYhKL1PuBd
rgsdnQ/QbIW0E27LDj/bp4CCf7aHVzhU0ybN537XY2dRi7GtYbxZ9JpZJHLBBJQdDghzKZjUD/gi
IsFqR7fubdhMIif/CSe//8jOqrSITzzSjjqo51Fy5Sjn7wO9YK/5KAYdam5qvAX0mLRnvZbwPWq3
kPxtQGcLkNrIuyWaNmVG/XR+EkAnXdGKdhU+VEdnb6HzQXOBBVsXyIDVfui7IbZsGkrIQasprETt
wmtIF7MoLONbZ81HjP6WNeYPsfyFoS9lMdFaBvkMc9yoT9tjvMOFCFmnDB3f+8yWhEfR8H+ggyUF
EtqBJKtq2GoRcvGqwlh19TmHIQKFTaL3HQTXo0twiu+cDvJwXFb6wE1enayUpUTiD35bAxOB60yM
rAomke7gTfezjo8psjZhcxCJ397vQlKCDrwi/up4yo6nehkYBF0PPXZY8tIRPneZ+6wBdAHPzUWb
q+TqLJ8OQYonD6UgX8KoDPGd2HbZGKaHi+f5GZrWp9p0TU62RFcONl+TYO9AAHpSoQWa4UQLTAzQ
33o0Hvu+SeVydpGe6UrRdYNENWDZmvxYgnayRZBP/t4FOcMVT6H9UZA9t+d7s8zfatyuk0ohR6oX
hbLdurZ/jvrmDtD2SXtDdxPUDE8Y5sVo40RQlxwRCluZtOkOHQMRyr1P2byOxsGJPoid5pJCAxvZ
mqGNafUT9uz+G5eG4LbsYKX75JykAnzVP4Y5NMIHnh5bwfjXbxK6kY331Wp+aFD+RFhpGZLYMCW3
jrQC8Q5rJ+49duwx42iL0/BrJw3ZRR0lle92zG3HwACO+glvePexedeUcaklJh6KRFUg+8lwGGO6
kHQRBm4gE1T/N++VH7Q1K2oqmrkK/TpXko5JNPuE23KIBlVyroxG0m/b08fVnL7zwAU+j/YL/MCN
UJFoQfHB28HWzs2YvYE/s5Vkac4bVL/GL/2sVrmsRk4GhqOk1cufFPi5jNYOn5cK2cXeJig3PVfm
AEVrhCzhkzqn3HxkkrbvdOWmOsB7CTiCIXh7qeGBVQMBk4ZPntgFzcVaxgBPuv4C/DQAPdz4HuYu
Pewnxe3f/pg5IDkpwDB+GaVCPKxhl8Fzd1GAYCKaGEwcAhBkRErlvG/BsUIjNr4ogWoFPmVc+rQ0
gPI7MWh9uRWwc9Dt8el9AUD37nzy4c/BGHhFMFZRch5b+0FnmE+Bu2MwP7q7vbtBnjX/7vF0atMB
H7AxN2aOcKRAA+j0UtHTwpSdFdjG57KNrY8WqG6CZK5n876QBuBXwnBcMEIYBM4EdlNTKnaI1yQr
OEf63LvP+PljO9ECaUViykl/+tOsr2ldvnQ2buisS+rhK1qq/m+DNMYTtUHqrX+XzPNXvb84P1H/
hGy03jE8WMKv3g7AouOhvE7whu0lZkVCiagKgRLbyfH8YOQ41sO7sCGVO0SQmTJJepJ7mBoNB94q
61Beyypmu54G2CKn928xaJuCawPtlesLjjPq5pYfI057Lv3sAC75kPI0KX5E6SpE8LWrJve2dUvI
UcGGSdzdcBpuA206dL0xTx8cAsCwvbl51P3O+1CQkYTYEN6xu4nlKuxfiXHHjM8qWZqdrnzS6vuD
ruFdgRtpdLU48ipcw6P/YmP1Vr6eQu7Xl7DH3LGbBZYB6Kus1G6KY8NHzUmDyytqPL5hJYpRLBZa
hwfCzcJSkbmLStV8ENaq1gPixaQA/iAzGmhXkZE+x0ZY7Mo/dNCPTe3bvuS2bzYslHKvS5S/dLCC
jxI2IBRDjBQP15KpH0NcXUHJVEcOVp8IYLN9sQmskLYGnEihPAcO+/GW3CfgLKgQK9mNfvDUpXLz
t9OUsECmM10sRPzGs1du+JRUgikwJTz9MmuDFEGVFbvAdoMlKrlOLsjetKekmBsDx2rcvIFNaMy2
Mq9RFnOiAYzq901noIm5HNfg50QQhue5lrNKUGpFjiu5ASiypaXAqXvnJMfMrX1K/eGeeis6mTou
4rAQR7WnH7QZZ1Kl/e3iLiD1JAWPhA/7/VPf/14mk77R4r/KQ0TnX/+nhpGlgRVx61xa01LbSurn
fFpnZNxh0xlU3jbNXCnStxubzDlyilSrkL25BdavYTWlco3qhPuIud78cJtYnVVzznp50oDhFsdv
2+OSmmb/qFM4Y4etDLzFG9GKOw0+8j9728eZ37o1AmZ2UpMMaHxY5psZsmvXWw3klJxDFjiDlZFs
7GQrTQcZEy83N/uvOozasLTwI0z4BrNQogd4n3YHaeOifSKYPT8rAeTkW2vbxwlrP5TG5r41Uwhj
tuKkbLFhZeAa2K8Pk6dLQHLKxNKHtLm1Sg9LXmuZLuZssHh60Ww7/ZuqfowMLNen3/xvA1wHz4hp
TGdeVzvs1WNssv2IZeo9bxRgbds+PeI2PKQtAyzmfbzHKCu/rFRa2f0kN/EYJXD5Lfkv1otxIMzB
wpi67NSUdwX7Q45CzuYbYdqv5jduEwzo4nFtLWrsjSmcH41nBrQCOtgCEjbbFiy3kR+dO/Q5+pqp
Xhu489qjz8DSUMqMc4FuYpSKbN7g/b3WH7vTB/12fy/sHQNZJRu/ST4sOh9zQoywz8k1WwQPpth/
Fhrq8odxaRvh3NK0GI/679jXq52+qQzXAb6GxuvyZrCx8Ob+8NP+6nIaeeIiO4nRAufUdIsXg007
bs3Kmpeld8RluS3ZizZgIurifrVR8rfc2F6Jh5lzN+K8D6icm/8yE+Nx1nsLBtjRReFV1r9/pNHG
OnnliYRgctW9B1CFYoAwjLsqTYU21iv16kt/qQJpTKs0WR0DxSpcxfjBiiIUTcdaWrH4wYiV8YB5
2AXu6ivn9XS37y/JV5TgRI4hfKxmEb4WG+pXyDKZDeeCPX5bs6PbZvIYuUnMjtkGDaiuTnEgKh1g
h19XaIz2Pp6r7zTPjor21Dfmn2zAfKAGoDeHytLnHe+dI2qtz1V2Q3I2u42brJR3k4pHprgq5l+n
OGrH6QXM+11Pydv8dAVJxxrk8D0t0nKsHY87tCzbIdDELyLcMjcEBgbTYLNWdTAQngmjBLu5eZMU
xQh4Sr6i8V6tLERcyixdIq/utGtfkidMkJDqeAXm+IJtiKD628VOuPNI23YGTp0fhZRiaRTS5NPA
7QXOkDt8uppRrKa7MpThbFLyXvzhJ8tku+JySzvhwYY+YWzSb5sTpWvmNrVCHlJMoc22npE3F9Kc
Eqd2p4yc6lcTZT6ugOzamWD5Z6iyx13cBsp0wzsF5l9TkL7qrcxpoTry3Y7U/1+Y2nnv2Bg6ezl6
mXRg9a3J0iKXtB6fOwQ6S5vm+31j//5ut11dxdFCItQfiuVg8/us0bPBTKwBqUd5woxrGmiUrn3K
uZbSV641EmuJ+7AVjjEB1/b8PA/lomw+OwKdVr/wYdvXH9NQGfQK9RTfLlxU1mlLeGHZ4J9/zbWg
VCo8xi3YPmhP7Ul5xxHdZWZVE6i0aQE6hlDE9T3zkmm+4U1kq/UQmCutusjnNR2Ziz9+y/jL1gxl
IbyJXus9IOjMF8zBBdZ2fqUfoPipQv5f2qoTfnD1f9gadT0MZ6MTqOCNWrOr85l2l/euCDe4EEJt
hYJKfFIIRQEKsUB8ns3bdl+7VYj+Qu9+vi6DPvPdmZ7z9qeu0zIqJ1VVUJxq6KpG2Codh5TM4HIl
fV0PAZ5iwn59VEGQbMYxqNPIjMkJOScFqGrZ5tTRgXwiTkpJzmM2j/DSJ9gU64DZTRiYImz8G08R
Ten98IkulZxOncim+KWDOnPzbktUKIA9rEdNBEikWA8QZr/UMCHoPmOG+T+yF/TQZdaxBcLNszHo
gOvKrHxh8gIT9wyaWV+IphkBkuU6SL7gA+BZ/2gwNiJqevymRkmWpVlgTBRhMeFpNdTmPyRbPR/c
DzsWPhlMWIi3MNiOFA1o3+c3fZarOwmvGcYwOKLSdj7Bl4JHvfIqngCcx1TbmcDlNJQ74zkZnFh5
XPZdDEUD4MF8C6bOqZCeMmxw5ka4ZTyg/K/BVGM8rlUW07rlVoUSqJAJKaAY6nSSuFnfwHP/sStF
f2z7enmWiygkEOkDiu0ElQ5mzoK70O2ciSyt5tmn0Mu2iT/6EUwe3rMYZmgFPRnCWXXf6SPD3f/o
bOMCqqVakVkydYZZFaLimIZTuC1qgza5lnFf1Lp8HWTd6EJ0B8PR25akfXaUxhSKunwbJlK2LyE1
rPvBJ+LDAC62pcMdXUODgIf5Wae4mTbORSwbVY9TbjVuUZyf3plKuTLNid/lYm26Zh6WCoqr3kQw
BYGgbrhzGro/tGxZg5wpL24sAc5u16YwJaWq9xpcBYdHIW5J/0NnmtSxl37ru3mevGMeRZ5v1UfU
nTLB6RYHh2ylWazWpvEjObRSSKCNcR+L7tSTX2L9jz84jsES0X7B3vPQLhQNSgQcZ1p50H0lTgz8
eSoIM0MOEzjlmg6snGI4c60P966ljMIS9esa2BXNagz+J41ui72EMpzOiXHLnWQ/hKxe63FsJrOc
q9Y6fuGFEQwajA+nc7g+xaXcwCr0BxbxlDiNYMLnt0z47AJvpNwAYKvmIy8Lc3QvGr5Et4wvJ3in
CcK5ThiuvdAbsetbZMEDNAlFfOF9mon3G53OhMgxbPHccnwF/yH6+JYAaBAejt/Qzx0r/tvWjkmw
VdP99KUi2UIbxkc02i5jlOxE/og5S7+QCThYdZm/gDdN6pnNiWIjwY5fpkVDQmf0KDDR6cfLfMZ8
d0tCnu2GbSYSjOIvG5fzyConI8FcxZfySP5+lagdD6+lq+E0p7A25Nf/EINM6aAA4Ak5dm8vNbuk
JysQz4tnK0E5FAccr6txcHNtTwUXz753HTI9/6VgJAYFyjavkL4+eaZMYwrUVqlWPt28ro8iel5E
YnzmA7FvLtr9t/MxlxN4mgiqyNqOhwobhEt/O6OFWFc09Bd8GK8R22YRQ60lWnFbMh/zKH8EZRkm
3I4k39TtWOjSNKUD5Vzp1rDhQAG71ImflZwVseUmoTY8NKpWMaLhDpdHedIWGtU1ss4mKy7jPRTd
+PxasMPM26auq3kYVpzMjeZz5O9SC1b4FsntQQdZCz+gk9GeCP4FM2iiNNCke2ZmqVTYuO0fOOcf
reF+xe3+0zEXzDbRgVcMmX+aptE2iHHSzKvp8Gorz0vVnZqmn3EWqa+zFlvFH7pPOwOzhLmjZn2i
FTbomcP32twt/lbl3rUv3JGdqe6u/jG5b6mCGlrcYS2OHXIouS1UyN8+LnpKnPV+WxaYmQ9aPt54
6UxoF3sKXlXpBeveJr1Di1nFEdJW1MFSSMPKGxWHQvdDiI0y2nBmgyW7f99SXYPG1Lp6G/pL9d12
ePnLPpndaDuPGBTUBtlpI8cG3b9WJeU8RlpaHc+n+HXnrykFzatRhzMXf95cRu8kbeGqOA0VX8hU
V1+whGh/mQv7IFhhs+FBSgRFk7rNBG9okodJipOQXviv/r3q95ik3d7DLqJhJ3twdEkGwDU5hBaZ
mvJP8jkAKEKXcz6Rj084lkvNOvvI1Sohnh1JrpsX16zL7+HUx5TwWU4+IZwjBYFqbDNI4huG1DXT
l9buDR5KB+tH3pq6Ekdmva9SRreMfTnto+/oR809/mbhWHWhOczw4gyWZyE2dWxA+LN03dYDtA2j
hIMgadhvbTvYKE/1kyEdqTrPtrmLf2+hIWgEZTDF+qmRaR6gNm+vXl22U2NyL+RwCSdL2s1ZQV3u
RMJ1JnzomjGgCSFywWIn1q62OhlZ55aiDaAQc8qsP+GwsS2LUkMok2MjWEvexuPHPnL8pFRYvZyv
qBdMWrkLQkU0vqJIcwLESB7wwHdSF/sASvaodmDuNMmrhhm1uWbKidpMR9Pemhr7c3ufX74F71bO
/LEF8GBol0Op+vWtrV2TD5J8rISDJlJJAXl6tEYQrdJhbeOhxhHmjGcSWxVe2e9nmgoH8YWhqLhz
gLxc7b6n3dKFtPBHYLqFk4JNMXgUysVvHoYWzG3wCERd4/aztI4HgjzUkyop1XEDtgbSesxAQPPS
o0Yi0MrjMLeB21Nabp4eo15/zvS2WVH2ffxggLn17xh/5TVKU2TTD0K/y5a3b9czfxJUwyRjQA8S
sovNdq0DgAJsMwLte/yj5gGTW0FxOGc918UEkuVPa1eRhiJqqh+e7t35H9h9Oa3Pqpg58mgj8+jK
RCD6Jtj73d3a81QWBG9HDyw5pZMW6X/EXSHN5xGI3Raz1pTq96A+hgORsWKglhGazIendnYYBCdt
NeVXqryJgcDofOH76YL9L5V0aoMFyhDMheYZFa1Kn3ItjfViriSngCwmbckqRhL9PdH9VEkPvLJI
QztlqtrsaCGvt5d88Rnn4p7SI1w1onSugh5ebGhrIgY8DTxKfpwl8FJ79HhHKpguJNH6qo7viRDn
Qxrszp7BN3M1ZQvMCSAd+mVELsou/AcnuF6+1L00Tipq9GnAah/LNgHoBkKTfMOtu/3NSo+rS5ZI
m5IyAeEGxj5F+hvBBgfjcyqy9bw9jyufs7GtAc2JTNL5r/RglmJK9zX5iuXo0sXWRfH6/Gbh5C//
4c0/LNVCmyjUiDv4GG/xd1iGsdsaQvkgMw2kPXicvoSm6utcoDUxkB8wRaTjIYE23OKvZF9mEMnf
QDtKLFo5T7aLQoC9xQdFO4VxcLOmCog5izgAyg95dRbnU3FGfIkPVmFz04LqiH5RxX8m6BCByb+z
ac6+GG83NDFTVEGb91HKae1v3ZY5X4qwLKeHg3BNQkFPI7bDN2zIOzfUemO89LcU5P7NZEgfKb7w
BSolFW8mvKJdBEAnr44/dldmx7CswFzs0ier+ZCR9S9xHXtyYmpRcC0AemZwFOYIJuWNaciVL6C/
mVORkcxBq1hGW7e5TI/ALkLcFE5wHnlsxXxjsHRZplpZejegvxSD3V9Zj9qtgFcInBYml3FaOy4A
pPnCNSfXzIftNN0cqaYeezLpFC2PsoZB0eY2vTetvGWs8k6cOQkiLwt7VO0Lt1uhrpVosk9J5qUj
Is3QpvToEwdPj+npAouAnto4Vds8W47/3VCMiPKWTXg8ekiJKkfASWLsApoh4dZdrzeExua1Z7Ai
mqLUv5H5ktc8kH2/vXZGhW4v584Ck7mIOLoJUpyhPQU8fc1Fpi6KXGT2Yg+PP/1GDHtXDq/5lEgN
HsUOic+wD+jjrTnF+sxhV+xg6NHXAvaslM6DAFz3g+wGbJPSAk0X+CkU8md1j3KiYzrPVEoZoLaK
Gj4HLmDZ7lcYbHM2DtithmkfGT32r2xo8T0NALwCnaF06hxK6Jj7v1VBn+xUU+36qLXjOxpbI+yj
yqEASc3VSxTXE1N7ypcvRvir0aTVnEmqyaADhW5dAdeBn5evPIiulZN47Q6GER4nuNjaTDIprqwf
HfaQoEPJZ0hE/7sLmmv0DKRQt7ljXAU3ZjPEeS3HCPTcpmsTiGa4zr0DEiND360J8PxlswCP47Pd
UqhBGEvM1hwdExeakiADqmUeXUoiX6za+OvLMagP7ECFcDmiuAKZ60KiixeNoHOFUsg1FZFNVfBQ
7g320ueXLc9X5oPFeVrBhxvCYg7nH1vxi45F8VhTqIpfLJy6i5ry/SzyFb8voiHwnR6OyP423mW1
/ZyjujX4W7i5LobF5ZQHDqgTVw+z+wc6pG/xbzaYKrfFPmJNZDVbLgSuYVl2lDYpS4APpkNu8ArM
FH7xl2bllZWBuKRV6Tdnp4nHCewF6xUXgoE2BTJqplUJ4L6FYov4wJ8MKmq4VsmVNsAALVULMCR0
1TY132q9plH306bbPVLHsFeUw4kQaHW4Cjh1hPEB6ZoZDv1xZ/fB9kK+xC/7CRk6heEizbBxb/ir
dAZG4KWi3mC/5XkqIJA1frV20B7LxrK1JziuxdgkmcA7qqEhCkSH6sG+SDPqfZUiMyq29dYMCiNS
wLXBq9lCKoGP1vurfyXjwXPEocZUdB8Naans2GuNJe8At/SSINacAWi/Mb370Jk0sgij8i4If1/n
+u/FgqCooJLUzWVB6oDNqu2cpuwrLFaVgP589XaK9XiQbkrGXG3fzBdnx0j3v2NS+ZMT96cY5234
uac6y4prXgNP/2o9kbACHGK69VjxynchaEQvY5bLk+5tROLzhmTF87OcZwyGkKhRDD8PACr2xh0K
0ss+Gjkgxa4hinYhpUdPKaa1uEzqSMN4HDGpkJERsp1shxIe4GjwKZ9xwcbRO/JB79bUPY+lw/Ym
Q9fn7Blx4KQ5Ou4dp4M7vhwUyARZNVZe5d6Wj9XFZ/UIsDcjqUxXGNKy+YtCCakmg2/TPT4cqGwh
5u8WklgHHa8JaoJs+BrT2Ajh6WB69SJaMpTmpZjIuvfyiQ3mpMPD6/uulapadmlBpU8DmYpJXvjf
Wu9YPGiLRVd6peGjWhXQgcCAJX87xu0UPMdm8pDE6o7kIpaOjwnBc2H7z1sokvsLdWxEjXFVaFc1
qYA8qMQncVhVfRPkhIJ7yyR2qP+o/9WKQMnEYwlVbf5iRO17Q71K4Wo0pl+j2jjrLXS8S9U123MT
iGdDq/1OceZMO0/+RgchttjfB7mpHZXCf7iZW8icM3fesRaggAJTum2HcJQVxWkfagQ74yNXAP2A
R/pDPzwIo5vfLPoGigs6yPo8uEVksj0azJqkSSpIl/hxUao8bWQc29aOgrgm7cRVi/SKApPTvZ7X
5LIwUlgQpYMhkDeZ6a8ThpJkFXq16mNagLuITTxYgGTt9ICzIhQIYcvLDtGscgOzTjFugg+SiH5b
xeIc4VvVi4MGAL1b7XUymcoavdWa7MjBYeGEqiNCdquwiRM4oUaNtt8lAJhjvVdgO6L/L83DNBic
Nj9vOC1JJeynuTlwVsCcUbdoB91lL+RPZT37gvy6cLuY9iDj6ciSNxiW3V/n8mLgkwa36W2TLsVA
PJPwga8w47GddRgIqQ7bn1WRTRJPCgRd++Yz6ythWe3Bz0qLlfwonNLmkVdF8h7jkZx88za+vHFd
F+HT0IOjerChZS02BG5b3+H+7oDGPqoFCUz22Dpxad7aok9RHz9i7hMRQBuhuuMsqd5SQhTat/hI
TBmGb1XWW8SeovBz++0aG+WEsG5W7OCcZsAOSEtlKbN69tyxj1jCmhLlXPSxcMG+4JeJNQTFEXXg
jpDrOXJlfiTrMMeQglNP1LL/uxsdZJIBpx0fjgaWHIeAIgNfavhMGNm0nVwsMw+tWCrVqEKwkcyU
HtpxxoENxpfs9bYHuiUki+YgmsUt3KBcmS87M5zScqkmwYGR0BPFmlvRhdz5sS+LbwgU7rKPpfn2
fRL323DTPa4pM+3mssDUSS76KxXH2r84HO40bnahLPVPCTdLbwSPT1ddlh++do/EDKELs+sVULhr
Dldz78wQvamKCAAHPwtcJjxNvkmP+Mjct+MFlpubmVRcaHCQSyMkwtir45wDffnLK6Pi3L89Ju3o
O5+y1N4sPVI5pWMYwngIBIPrF5jivi6XYDv8M7MUuaZLsW4bdLADGN3smcwnQXA6ggghDgdfbbvX
dKn5kT0Ve67vnCeBOYpNoGC42VvvNEPlluHXtSA3vFTjO/6kAmzRFFN6p+ZONeiLN5eJ7lt9WxTz
3uZdfc/k6OHo7ipR8IZdYnWGEMghdImxiERbk0ZNYD3TAzIjR8otMXnHzpsYY3ADRfJPzHjYP3H2
ZxTKko6eEEFLEG9WT0K+0pUxIeRYjFtc1xiITqX3okLUnw1h9w1rV/3y8014eKGFRm82mFgKShOG
rjIJ4LiUgZckT7NmtOt7FvwwIpsTfXFqHMKWP0zB2sa4UnjLdeYDo9dfnDf119BNPikITVc1G1+f
zo60NwqGjofjMm1GVgWzkmaBYxrHk1TlMVHQoSve0L182NRicdMYAhfy0C9H6HSPEpVeGnXpACNe
y0eL8nMst2rZOYotEW1/GUexHhBAaKrGr5w/RMkzr7J90+/TMjVi7y9vYQrGAOdXSy4+PxZ/URQO
Sf2HKD01cUavhQuc2bwYiiIsqU8fyrovyeoltejZymjNlpfo1MsrNkyObGrbBBuv3JJnSe7Esn3q
oPn04Y9doMqszxr/CfzA369AEWu4dit9zM1omJtFiN9ZbL72tL/KeUFZvLsPIFwL/blwvC0aLdf9
Wwg9bHkb7wlUhwweKqsXpAMcF/T+2eLheQu3N26ACz7Tb0td6iGnKESLIpDu/UkHgg1/eM4zBrZI
NLRXxvgXL4m7lIll/HzZtpP79sPRpc4krRrEYfMKYeR0gW1WJuZoQVIJEWUMmCJjY4T4SxPqKW7k
QG59fMSqcis1lObshd7hu0M9tuR+4JO4I6dLJP5SIAXO0kxooaUmaLjvbVb3beZU0iT9Wb8uJEcW
GaY1dSfxPc/BOJTtNg2wZkcvyLrlPIz8Aeu7tpVvF1cnZLOU2qhptGAB/JyFxMfQU7xdYIZI9sXF
K3lviZQhrT6WDKN4QBEvbSGi199RaThxa7Zpa94qBpE6ocUQN64YFBDtQunmGWlYVl/vzL3a4K3S
lO4cmlHGoypR53smSKjI8G4UrVt+N53fJlhsz8aea95XEip1AqeBiQmO8+fU5JkFlRMWOZYBwPQC
WvEWmVrCKfdMG2phiTc2sTD4ZyGDzxELauQ4LEXWYnOpeA+Jx6d2b934xMIMn82gS73mmjlCNDrr
OX+D2WOquAwt5lC8vb9LgvYICFT1+9LS2MDe0Rm+reQhkb0TJvyjX26opGVWC12ImqpFar/4ghk9
9POCz73jnWCi802farz9YoaubF0dMmxEUbV+UpG4RdkQziKoD4NjaHOAPWAXF7DKLm16LkDgC30O
2KgW+Wc9D7ijM6fT1ZNilB9jyKaFDsrpOgtg5peuzF9fCR+snBOuUq3QUlYWvb5T5dh/m0hiBKgt
rC39nLsoRrHqvxeijg6b8dYczdpPUYT0ZHW/oJE8Duc8YpBLDiJDMzmHaUme3aRSXQF6pNT1Szuo
NtLQV/P9toBIASgEXMXh1Pg54VLrI0JwDmTkQSuTwT3n8LS1JuZfmUWfgmS8RENEQ43KGOHlGmFh
gK3BB47eufG9IfyAnmrxts+7moxZ8z6sioEIY1nomp5/py49d7ZvbkderbxP+Lxhyn5Qi1Bo3it2
Q+/zMmrA4yJF9mDckkT7elMVMfGeKGNWLFAXguTUCj4h7NqZfNMwfQyOlxe3YtN7Es7HqU7C+S+2
KdcZqZfPhc64QADl8P3mnEvReWrdYgizS1CeXJ0Ofa1+lzrfTSw0iYplPOu9kCMjptTYo0LRNacq
826DXHA/vZIrX2eIyuOMqHDarpQDM5zYjDWqeMVWV1kgxprwDm0tPcrf/dIKu+fVAMDWFD7wrj5G
UmyAxhQ1Ui7X9FMQ5qbBYIa7DLzOZG7fSyuZKOnVEVklQ9zyDpNbS9854mmv1zUVVWXkbUJIdA43
uh81WY4ARDLA1O+3Z3QZiEYMdOT+0dd1vGGu+Ct5Uuy+UwNw94Egjfw20UadTzq9163mBSTYdd1B
+b2PfbIhgxE/opZ3QZoDtye0VgTa5NhttNZw2B6ggfDHgEkPh5Hxm0+DI+a0QMOyO2Nr5D1aKa/H
opDKqveMg7raPUYqGPhc8MiTxkUzWZC2w9ARZ/MiKV4nBVvMCUAqU1UcJ9BtAlRBzjO3qmYD75Cl
sodOQvY/vmsnl2g42EL+okJmwWjk1B13un372NI5PV4mewwaUvty9VZlGcau29g1874rB4qkKUPc
PvKLXWhUknLqQq03kylGUy/au+WXy3oQIwtjZ0G9lAkpT/TlnSYoqVAgPl3BP4f6BVUi4RkpoCB6
s/RkDi0qnk6zhJKbNKpWpuYbVkJbMhUsbNpvavBJWWeVeZ5GyUEcerLnACp4UmZ5f4GYCdy8CzLo
ytDa2+GJvlj+NnaWPZMtDVHsrHUfkRawVaASf3CQ77b5/aRqp6IvfX2j7zUXqbk50J/CjTtucIs0
+DqArLqrkUodDeFyX2GERoDCWiyydvoqhDbeUXcA/uqxQkPcscNqZQ9fLK2d8HqRBLsRwJPp/83U
ZNy1k0CYFolx4vYDGwr9f/iLiI1iDph4UQKiD8nmKWaOSBIaUQr+nAYw1tbkyZuKTS/XfxL19nq9
ymOQOyyy3M/MCvUmE9Zve5LmqvReu1ynOdxGMT043o8YVQfTiw3ub8a4j8BOjWlONiekANIveAxd
siK4xuofCnAfjqI0K3zBdvC3pgI0KxIVlLvkyqHNVSssZM8oaFYADqW8vPc7kYcdSPKGkmxwCTK6
f45wl8NiNbJaETDKgYndSaCrCUYylkH+lUDcNXf+smAH7oqgbdDYJ014w3V5OjIokKR/DAArTpqp
8eWXdPIKgdoQhG1anAwftw9e7pI73+YgBiIw4b+mOxpUaY9/JeQkSyTE+7IZUF7IRRmfqR33/D7y
S3NPyNQ2aSvelO85GLAYMZ+2vUBLuval3jsYTXBRM7ItxeEtxCJWLmUVCMI5aEopB227Z2Yr5r+Z
MGggge/evQ3hPPrThfi6q//IGNBu1TUBUt0U633QZGKD2Ox9JJ5bwBU4nOiQAFDpoLESlqajmBfo
Wuld8/SPTWO862Vseh3Dx0c/R1kr8FqfYXFoO7j+3HOUpk2KpLR3k8II7HMtEx3hDlC9hC2d1nOl
uvNSryxQsmyRNpuEYehXpGTvyLPKS9Cr5oDrEUm9M3UFDjPEvAX9YO0tjUy0c07rh7z1En+vGp0J
jxMxhgRn5RBYEOJXQzzVC4/5CgkvRP2LiIZatU7JVMmL0PrZtb3UFtyILdzT4ZbNX1oM2FtJC44e
FQLwGtH6gUyjs1e2/8uV2tttC30Eo3FGLDmfJSwij4i/44rNFDq5+lKLzSbZgpmIgFtZwc0kOJN3
YlsMIcMhmJKRI6fs/XYne5yoNAPtQSGWLbbgfN41xpoxXHxiAdfoCmyDvJhKVU1ZyDNL9meO56ov
5wKBC9EDKNYPE4DKQx0UJNAnaggdI51YmYzPXLQ1Uf8Oz2ou5bgToAAfLCNaL4qmx/j9uThnStiJ
4DLAvQ1xmUJ3gv654A1bKlzwF3haz4nHmC5HgwkbezKVIay/KrXk44uzV8R5gjzkV4uq1LJPYhTr
KXONOtxjckK0cbnAYRKL9rb+cpjP4Ia9sqLb6jdCVKjq9cYzYxNBnAFIOExW1NOjwzeCKvS5o/nk
blISfLukbWUSulCivaK8M8q8CfTxV95Ey1+WGhjha00uM74HNkEF4VpLAYLHx3ifEZ1gf1ku06RG
I6l2nEQnyGOTUCiBh4CctpEsFQgeskuvlA2LejLvpXP8oY+eZmbMY5Q6hJ52N46QC1ijILcQ9I4C
sY5PS35594pG10fZ4rE+02HeS2mVsWrKU6co9lZUrxG0CnpF5OskniVr4WZ9U6CEmGtiUS890yW+
AiCPlZwEGY5RG7rfmd+VNUpGtueK57PVUj8s4QzspM1aFBq5vlybBfqpDwfxGVP4DkT1dguyhL46
l2rZtabZANuktvYbw5vUjhbmYvpIETyYHLB55+E4jzFXS3rmtoBB/8ITA3pAEup209vSTZjHPufM
n7B8EhYn3+eF1do/JdsmViguXPF0TlPTWbexcxe0SkiWALauo6MUzdFcq0OF5G90Opr2F8z7TS/b
Oly0ZV9cACAjljOjEqcp7MdJBb8Bub1Yasv16OBXFXZ4PZTU5r5RV/3qY/Cbzh3VQAdC7EsgiHS4
NX2/nPUPP6iHMRQMe8k0yWW6k4BHxUCL4RlHEWCgwpH/U2NQ2kh1TN5lPiUD1WzVUooPIQaRcdwi
fcchuW/XJmhuHjVY5gsjCkprk2/fymbQEy7gZBoKAKV59fyN7y1N1J8jA/m5FpttuJzHNUSmfEFk
hnz6Cd/nO6JhA7AkktP2fsGih0vr6dAqqCet38T7HtFaYaEvT7BpNUZmzgd6sraPT0sveHTZRfnF
Z6gVkqMLthwP7HTaonYzZy44UI/9uMKxi4ikn1pJLNeTU03JxAzWtroxjkuklPhmy4kyJwTuYOuG
mjWlvc8GjYa7NBpjRRCp9tC0M8bhUApP93DT3YGHdh0l0PKBF4LBwFILk6lMjxOGD33sR5D4PKy0
695e44ozweCgO7I/+K2I+7t+IHoMKPOtWmse64VADbLLMKhwquW2rj5LXYE2NrzTDJSK+NJJ8M0/
FKoXCL2W8yzvfHyywJ75ZFIAAV6cnKDqf9h/3qH/zSDmaTIHpZpRCQInFabcaS4O/8TKibNIUtA7
1LOrBq+SUvVYG9hFo0e2e+Wg/heRiXMr7PrwZHlVZHH/3b3q6bubp72ht8NZ00FEGAiNXbDkwViD
y8W8ymGeETGnGwYCuY+o+0ocCitmsP3B0bxpPLVVxtZqBTVvniRUMZyraiYwAlfmScwe02Su5qjT
Z+MHiiNy5MRBd1Wp3EsfIRidZaRP6EnFQ1+1ERI/6GhAgtACjmukz9sGvThk7SHtb5vj8Xvu5FUI
aDdWPnBiNVVZ4RvAg5PIiPx9LLxM4kq8e100VfKMIcejbrAmMRnCUW/oaeP0jkRb1XVJbklVCuPC
1QyPI3c3BMGQ5umjDW10jvs+p/ytGaNTnVtuIxNO5YK9IzyloxC2QAMDOCXYVk+qm5y9ddI9OAhT
Gkb9FuFdU1JGvhr8E2sz7P+ecv1U2rfxm6gNbtWJr6l31v7xOUyyE6SzW9+pTNLoZBmsB0+66qUA
7CbQDbb21b/dUkhGMFez3leD8GIQv5Nkt0Fo7hY2kK/7D9QgiOrMlRJVeK5PoWBOZmS5moL1frU1
Rthp87pfZ/jAdhwGIKKTLGHMnYGfYBLjlzG8GJSxxrvpegfW0gliqrx/9spyB3TF8nlW+gJmVAzr
bgLiz6/osy0T2Rk+FhM1URkVj/HAT5Lvwf5QdGRMTRiLXcgu1G7ZXUb0Kb403IF6kDmfgZPfRRBD
yUVCawHSfL2mhfZtAFpFY0LlVdSe1pqyRw96qkBMKNpChEGxTpvEmU6+HBlvFtS4pJXtOjLJiUVi
kSyjEYTM/NmXwxkxFhalCAY778MdQNL85gjaYo4mT+k1iX6OvaruKFWNEH3VQoWKMtYDHSid7P6Q
lvi4DZ0LBlpU9x74rr7ydgaBFZgJkHwJouXE3ogCRGTmhS2ysZJND0PZgei7U33LRW82wn8DsDOr
+mpcgO/AkFi6KleSHJm22b24H+spmTpqgPl8ECDUMIoE+LjrncH0G1NcMdIdsrjKP8UdaFhvFVYe
AxeOtmVqfE63bQ5nhNJWK6T5SKY5E7pZejQzaFhVLbcuzupmCg/J5VfEGZiAbyT2SEt7BrRdwCUY
lvCodJ07dMSEmBnfDsplFBL2iIg+4qGWIJw4D/26DcqpADLHtC1PadZjNQYbOLJS5Fn07hPV0Gj5
qz1KRq5Pt05aftm2ZQYH4V7K9YPCAIxyKC8ZJgIHdImuoYex324vxIsyw7aGdKSH/vzZ0tB2gNf/
DuOBlv/Nc5xfjMurKAKUvyJ8RCwr6Io/6T6nu/SiLteYA0hRc3cnSMGZYkdAhisl1ED63XG6CYuc
NB2tnPpMvTYyc92Zb4or0JMNsQGAnmWqcYnKhess17oT9/XFMcuKEw9e76otpxRQfMy35MbL+uLK
tUlMzhsUyjiVSESFM6/QeWCbj/5mgGXcCYRf/Yq2XOB5EPCs/NhP81XLaZCCVkTcqUNE1Rrmw8U0
EYGjdIevuN7JNZ+h2NGqro1Q1zevYfy3wemkCnaZR3N71NuTykqBidclWRmEYZd2VVCPFoelmWas
DVMVRVIs5KAb5Y0LMkwGC2de3AUNCbVncGp15wjoumsipU9D9bAiLt5LAbUPEnbZSvDhzlH079mu
w/z/k977tvRWJb2T7APja6ThRxQ61z0RsaxGfnskzauyd0chqZTrfCa47JhRz4FutOxtyVJGQQM3
eNcvvTCydqMwvN7vQaVemmnlRmmOr3I/dUYhRMI8wkzs/oG1ok/nFvkGwcpATUsrzZKCymmTh+6x
xY6T2YQfHGhIONbGGxDjBiJ2HIf1Tx1PPFiVvvFb4dTgZOCfaZ3j+BYslsxwP0OwWHakrBNlPITz
RrMyBoaSv+GVYflMEl0LP2di92TTiuiA0nbkP5BN2SvaweIBhVjmC8E5vea/t0ByZnkwskMiupXq
BSPvYzU/CU6wtqRh/bX82mWjpMRPfIXZl8udafDO1HXMDJlltC8dxuS7CcRMZXCzT7BlaY93cqfT
3mwbvwvbv4McMHbrSwRg4ov2fc9lmZ5y4+ZwWCcd9m2QIQ2B86EzspHGmuG7ukohJgx1WWkSlzS6
z+GEQktXn1GOsav1Wk78wjLoVEjAbojqvKK57ZxchdUcqzotfYp+dtKd1Mc2qV4HVihXGnTVVfmX
vw7m5QnYzCiwzWBWgwDevgNpkvdk6QhF4b+0morddQP5e0exY447U4CreTQTK4db55bun8SzgGkr
Cl5eCiAxSunBk2xy2GWWvMkZaKb3h6dhzb5H3IrNzL2f5CdnMWDeyxyQ8shQ48ocJg34QQTuwIWx
ZpH2KL7i2mo+RSdPkxYNlXBi7AZztka7rtrFUrn5660+mZFXwU0GagprZdmnXnO0KfSu8G4gpWVP
H/TNIW/Ib5kbgH+81Uj8SeMbrCXFcrW2eCSrLSW0ulHQscq/Kgq+6EvSnFdRZ/pbPLh+hsl+1aHN
q6Ce/82gy2y/CkHrHmpaNjkUYiXxmp5uesGFAIyj/bBpXAR2iABmUDB1QReeXN5rx5r6mOnVMwPS
EnDQ42oQHWTYkMmmNiElLzGEEurheraVrnVeSASWA1SHjbtVlWzvEH7rlSTnas6IMpNBXCta4I/+
igVnd4QIJPAFmhuHkx3bGPbwdth8uuArk/QrU3RkB2u8uV/hWBbLGuaC4bOg2rQITY55Z5qR1FGQ
WmA1QOm4iW51mHtbmBGnVmhj4MxpL74Vf9fINTO8dJAwVUmDK5eZu2SY5yH/4v+Frw10f+VrpOuU
6EtNT/6+nsJDX4Z5nVgIaAxYR/nWa6MA1lWxJZdwDHaMM1DaUtD5exvYeL9lXKV2xDOI8e9c0qM2
2X3NavNdWVKWzEpEa86mz5SSZXemam3lkGczm+zdai+mvqqB/6KDpFRfyPYL1iN+YrLHNU7o2zNn
bpX4WFsUG8f8JtMgvMbu41EHbar0H0PujHWID4yorKPUF96W1nAJAHEo8mn2e/oXxDHiIB0T033j
0Lz3tr8wEa5cXKpYz/QZBX76y5GGXpm+CA9K/S70bK9JbkBJgkFFXWraOVQUTeWCBAg1YnqgPscj
meEliv9mVe1XJQXV6qqjT2nIG0FvICoDEu3OH+T4y60HNgGavkx4pJLm63/ILhLqx5awGmL/ElL4
5URnTdRBWeV2tiol9CMxZ1E6sLEGx80QkYHW38Cqm15XDQNeWFzBd/0QijL54E+LRBb3v1igHhQO
fUucqEvUgwQFN4Mp7jqaPHS9QmSeGGGbKwmIhef7/OQLBEVf34NIM4hCDiwQNhHzGeAOBeXdiPtI
OZVJJCXUrXkEfiOKo3FM4NyCfcTSsgENdhwWe72msWa2rybJb/m/uCQCZWO3K01ZkLwD7IDWjQLB
io1CvrQRah15Rni9s/yJfYr2TEDzWUHSuaaP1tL4SMjuRz4+DEo3l3UO8nsQXxWH/iPIcUQD4Zn8
LGfH89h30ZtA0u4Paeg1zzg8iTxbRXVqeH40pPQU72r4nX7ukKPaQ1mHybUkCZ+tAwjWCCVYBf6g
QM4EPO3N3XcYYunZuV2OsrOhYhHFkCWTwXJHFOM+OsUGqVXIdb+oMriFzKBN9IJHNdk2QSZ07Tgq
XClP20NAxVDtcNWCPMOjqfUmlFmjD8HVQrKcxzMGdxTSBze4sMLFmK7tP6QcpIrBk4Hq00ke2m2r
o3DRWblr4qSKKbkHsBRDCsp59+Fnhzk3/ARClegem4G1kPjIB/qNebgOdNy4wMTf8nAkUmSMDlV3
RapoBOosj9BG2FS4U59eBA4+0VCiqpJ8qJ6MK59Ftdifa3ncSbARCOADW7ojg4E1qirnEYEURvR2
AngTIXJI3bR1ImxR048ApZvif08clh5hLXTb7MWDJ/AxoyFPSJGk+R3f24+l5Ql1E9xZ3BHV0Ns0
LR9ZxIGTHhKvplcWkJYobnbdvqyrphiEqZ1GE32fc3W71cUN5wmtB97LX/2Ie7ACSnRjtYxB6Pdl
gja6sE4zPoi3Fc0SH4T4OJu07rFb2F729JF4NZDeMTMEjSYRkOdPbPijNhCBaoQWl6po7AEiFtkM
58yS8QLyHxJf+5mpJidZx9p/tOVIo+umz18iE+j+8zuVHh9mCib1AcUs51fT1V1dnePiIRxiykqo
1p5ZhFPsQyHQWZXtY0V2on3+ApKfFqSc3ppZdgqWqBHxOTai66aUhIPBGkMcJm3lRPQAYdj78032
9a7GrC6JLEglkKL2veS6S30e9itEi3E9TjyR1QuYYy0923sQS0Qx5ZrHCpawZaWvdqFvUD9vv9lR
eesmNGY4tPklGBc/tk8VJ744c9KSKUsCwEKsgX+5OYt/XBWtK+u7xWzTMWxRgRKmapWPDcuVvTqE
ayI12thl/SnZqpvrFrz8SjRXE+TUE0MoWLVRYRexmLFWWleL2TXCjYacz7pI8PVm65gbPM8fDptw
H6qy1ShxXZrw9AJlUNDAQyOys6YHMPLULPV1emyII/5w2RhncTBauCV3dKuKKQEzZ3ySsq9FXTm6
6QYuMgJz+Zfyw9OfbewQ7NBK28pQj7mGNaQzWUKnhi3EYtQDykjOe0kX7jX27enFVJtnRNgCtUQV
r8uTXg5jDniF+e9Z9h0Hd9eRiy9cBXmkS44Jui0eC/V/dixG8pYxBzHK0imuLEa6Dxc0vUIf9TqP
8KIrWl3v0pSbLxw3GxhLOinTiefT5DgmldaKnTX+k/rNRQpVR0VK/gQjr4esbzGkXz0gB/N09RF+
NsdF+OWgrDPX9ALloO5mUtriFawlW4ZmnyAX/Ei7xX/azzDoByKYnlMWOBTG1LK5+L+i9Ncb8r+u
671fUV2kUQtEpd56tqPr4IcRe30TmmWoGjGZuwwDzvlrzCe4Fy0yVlwvu9Mc87Rd81M/9hlMVhLx
fhfSCBz9y+7p+nGGgv7bQsMvj/gKmnUL/3pF7eaEeCcZwhwavs7Tz4Wl5U9eKVu+ZgEudBanHwQN
GGvzBwYEVnjaVkhsUFiagQcxWSIweeHX3Sm+8RCzwYIBbvfJOKT80b4zMYw1SPpWwPlNwD/fKkY5
ppRr3b5UpzUfuD2rCu23JzB+hIr5Tx7cMJNA77XPJQrIjnqucSnVpTfCJri8cgORwSTkQiFGwJle
ds40Tmzg9wlrG19jMn6i6F5elYXoX/HYLQAgWmrZ6+FQR8TkXyPOWMXBxgKRP9TUVTh7+LA1KhWv
MPauATNf3foyaa4zfFDUoCkiwjJX+i3IqZRnNm1JgNmhjgu7PcaocfOf+RLEUPD6QG59RHhFVq3/
g0Ur/Ud4lQGIT5Alxl6XAYpOkWhcWYtEQqGjbQR2Xb8dvpoNMee6aluX6Wq5XY4tH3R59pLcF5ME
MTb3nNWcVgqlOVojGTw5HjSPXztsx2oXQIpQPz5ZzCA8dIjZ3G+7aJhdTNqF4ON1k2/ccHEeQmsD
PJQqIR0Ug0ZASa/1lMXiwF478g+JYqWbI7qFZmRRl7In8n15KsF548cUoxW1ddaif+AyQ/JXwE78
cxQNG8Q/kKBNYHniqv3uL9PyuFA9TxfflHUEpn919GMyMAEpyIqq+ZP0H8wdUaWO8rcP5RA7JVEU
OQ8mECTPliY6CyqmjUwYGm/W7QEF+BlQoFf/KeTAl8mj1gXbIdPCm3FjXfelzyK6QkvRqS/0X+mj
BZGsvm9NRFcajfTHI28QPC0vjx2a71v+SEWDzlAGPcOKkDCYolRG4UcnAjjXCIBTxaZ5FvFjarEx
SZqYb5oIA6FR93S+9XIQda/o8fER2TFYzbtwUmEJtmGGftZHzIh/R75Luitsot0i7NqKFOlwYqg4
z2fLWsDdO53EN4QONF4MJYcM2lMJmci7jCa4QD7dvPmqZ7HWDwc8KYbz5VA4A4WGI0KPStaTDZjx
IH3lWyYtu0bfZeGoTZyNU9e9AKauGzF8IZL3D1oSBF8dV9bzQyys35F3N/zG9VD7JgCisYJsFDEN
MlNA5la9Ek0NmS0tIdmRbRnDkNe+YZtOc5uVhmhUi1+2SZTcUwvXdWfeH7UatJDvsByhlbS9aI5h
d1X6oRT+RsTz9R80E2qc3Tb8/GrScbresKNy4nTVokjJPForqc/j6OK1vg1Q3Cw+KMz48MzIbZac
5UT2vsGKr1VqPKjkRj6OrOP3IQEKPqRq8Zv2poXHfFFiUC9frhirp/uq/Fi9OpTnRinwwikMkbIM
vgXd11T5cEfpfyBtjh68vb7qf1Zo23XNgWRxe9d8VHP6EHRdHdublsCU3YI3z2qdwo5aKXy1S+O+
lQCBJJb+XgwAChrbPeNyuKxyelQEibWUJ5g5p3FMc8+HrL8G0RYbYvhbTtcdWUObMYxJutfHjGRf
lT4WeKLc/+40AZEt18c5bTyyW1FNfJ3Q8tAzmC2e/6Zt0pSlkKmMWvtFmnVEZL/PhGlRumDgxf+4
Ybl3CN2hps9z8dt2AJ/pTHcbbZrXtpGhXqjp5GH38ORVHBiFUi0Ngm1cX21S1aalXgkX635lVaTi
iJVBN71zo/TxtZztuhtkpf1wRrQiHYaA2/7+TnlJoiokt46PqGVUtCBcz8zSZt/ycueTjx9H0sr+
+YBQPmTZ/xCZD1x6Jp3uvL8wl68dgiRNpV367EsxxqPK5qXyNP6y8P5cu33EbIW6dxc+45U/6D2O
kb46JeFTY9tHY6SoqlO3VRimmPhVFK1MPRzJeZCWND/IL7X8JtteZGFO5VTDyWdmWwP2JhYNc9Wy
HQF0T3vA31QZ4VL24h9Pr6OWbSE//1/4TzoIL32FDYydW2ktN+cVzcZWCWriwsKur8BFW99Pat08
QbaUN8mVCPe0zYkWJ5pEIFxx2ta4Jl1QMcs/YbBeeRFMVLJqXIwWXlLAsHwXTOMhToo6v9FBCqSN
afUnPDcB2GqjHR52bbyIuo0o2H2W/KgV5v0ncbVtBCfezH4ZsTDurGv9WHJU1UqmKkMO4BfJcY69
27IZ4pBnxG3LaYVVyPz8wh600nQBnlZfvFkJkSYIlIKwThBcO3FhvLSjKqkPUDlBC+IPASw9Vkeb
jaWnZTcReRZyfoKbhQdvzbHUEWEoxJ6W/JFSvshyXv1QnytlcfocKIRYS9ICw5+UjB9nteZexblz
1Q5iQ2+O55vB3jQHI+SMhj26Z3AZa5PYbLdTPa1MfWc5IxwENInuApZVyqy/npUjbCCIkQwJVeKQ
94/acFDfHskjQk0aBDe0wklVblmoXZmkgyr+Zi9RN3+N19ckynIIMjKfXj1eGCeGWSX+8EuXDpoF
q9pnyWfFMMDkc/LbUEtZI8x44DWtR/a5/RrG1pLdmyLvPLDc/5iAhOUg5tFfFb1ZbIqDds1HwZdy
38Wo6gb9pmu3k6a4vEGbwlQRiiMXOaPPxORPDW3sWUfhW8qO7TZkrlr0LRpabgzMP1/O7EPRt69o
WGNu8cUFoSjep31l/R6+Q2jQi+14kKdmkFOVGFjuy16U4n1SE4DNEcnj30PQ6uu1rXoXIKDDz78i
q3f4cTunBuoh6cr2sY/BFk6lrPxCvRXvpnSaWl8QLxZXrGt7dTmSedji/v7JBbOf0zjqqKgzy+vj
AJn+gmE6YsO0aHYESRjqoy9bp683stANAVK3/6YyftZ9TqwNexdJIJ8V59GHibQLnbC1OeKBexbm
cfjGi1mO0tyz5da9HVdGIxI/XSVFJEx2FX/ohQmdkxrSe9I26Oj3+e32hhK3CYh2SWQhMGTS5L/0
ZowO41OVmsw5S/Q5et61dcs8Lku58tBbW+4uhOGn6LZNt0k+uWSwCfyPRM32g3nPBY+NCOPMUuoL
YqqnfTZ2y/pKCtVFeYrnYa6dwLW+XVwtbSScEwM3h5u0joWULj67Vi4xKmNmIdBo+iETbORJ4PZm
wH95IbLqsLWsaQzk/Pfi5CUrDEy9YU/PHECTBKPo8rMQg/H1xlAN9sJW2H9n5N9gQWr6VrrEprEt
4ipRPOnfViRw1caW6ucDTijlHFU9S2sRBIJN4X1JU/DGxqo46cYfRKhDp71KbB5kHd0FpFBzj81I
0AcanocBhLAh9bnNXvSNvMy4tLblM3vd3Lt5CZwsdSfXq55egZ/A5ixbysT//V+vPRzpOhYyzUa9
D2n6trgpEPI3cSA3RupT5Unz9lzNg4eA1ZQi29H5ZAgw4VlHCPpP1UK5tD3nfwIO/aZT1bV5aSxP
LNjdzQB3R/NIV6vHJsGggc6mX1IAuICYseKkWKBsmNCdWzH4tDtArRdjbMS0wLDFxoa/2UDeSIe5
wmJCr/SUslqVvHmCknuEs7hiy0psKGxWpI9QPH2y2XjewFP2hQj1TmM0A+tUlViafx7P9tNFXJ2X
3wNBJS0j1Wxdk2BuQotKH4cBMnfAMEqKpSJlfGTU/HLYN41NpvFn6xgZYkrf2eAHMlOmWcBK6akB
5wlIQMjEhCjuhh83h8pGkBVhX0Dp3PjMAg5yipWO/QeBvNQ6/21/qVc8ZoUitTCFvcdgwGJuipxY
k2WY504VutK96+gCmU6ka7ZqLmluFb2PI1rt8QB9TPi7miwLsKQhHCf6pTaJsvYiPI1QVvOu8bqw
i51tR+cTTI4eTBtUihOr1MDdxTpZcsi4+k2uIv3QhLIOCV2JWKAJqXM28FF+rlsii0foLsUo4CtP
ujAprChcYCONuwvX71wuRNPjN9EUds+KtW7OR7flmldSYsSApMpXRlaTvgZCRMy7nfZy0bg/Ej8R
azJ2T+JE0RM9Nb2FEWSiR0wkI3FQL81NtZGxdLUzLYfEk/AkUZer6BaKxQlob+31Hkxru+SeAlZy
bqU0t/6uHqAtkD8Paw3WdLRRB0lfuXJIO4z/E+NYH1W2GRUhJdQXoRrk2QXAF9tDCUMCwjZ/pJkn
bRQ0W/jzkxb3JV2INLyHpWpWOjBVNl4lSsvFy/8A7Xf6AWMLvNxV959BvIPP79vs8YquFgnbf6/q
oT6YF8WligA1mHGSm9Z0/ToXRRwpVohpF31g/rGA92c4HqI4jJfRp/cUjbTkCTdRdC7a70PTX4ue
huEWRGDkXr2aT/YSoe9QJgDqOECM2xq7vxm5XVjVefTaNRFM+WLv012NBL1i93pFDAr9oESRYMSN
nl4SI2KUYXBX/s6LUDaJu1Saztgwi7Vr8fKoMmH9/6+RLZ0ElVY9hbNFQuucJ5Eeyu3Mk2jvWxvb
RvWYI74H55EMYxH1Wle9itgRDuRoBsF5gby5hDc5YQxDoJ+1slE9PO+tKzooBpLI9FDWUwJSn3mk
bdGOscMkJaN176lZ92HOhsAfsrY3cAdMF4nYCUhGfR7gkkXX8f0wU2WnYEnYwWhxl/l5tSqo2Pqm
otIpMZmBgQldGyItXAm3HfW9jK8rffgVBGrbDgUQbShkyyT08vco7HDaRi+uFM/igtBwkbgs3y0U
L2GyxzArrqz93SGZ2eMrsROuzJnyYIV+GR5quO+6/rf+S+4lt0wBwcJWq7OsX08/sHP2wCTKejgr
nXF1R81ARYCVfOlX7mzWwghIFGrR/jyJa26ZWyqHtOSQmG661e0rvShzv7ZcNJtaNRNNkCjkn9Tv
Jtiw6CmSrC5vGdoIHMlOlYp5a/euJ9KANo/yRWGjnDBRKfbY6zaAQc8NccV5d/1Q3AN3yZzY5JZd
4121oiiBIKtre8FFr984RwS9rXEptd19/ryhjzI2vL/jF4KJvuJfDGZQS96qkMleZCbBeVRI50rT
yU6ZtcBGvlc6l4zSUVmJWIaASAbWFiNU6rbcVyfpfj4ChvxBkNhq/ppq9ZitouCCm10c1Y5Z8918
wpfezLQuz1iZfuy1O68jkmAE8q4fqOGVKrhAobwkXdFvJpU9TDm/GsBfG6WijACcwbpmCQAC5w0t
BHYMjqS/SoosmUo4v0AyAwxA7BVZA0NAsl60uGJT8bS/mGcagvDN9GPoTidhmBKPTzFO5S37O9Qx
JEbKxP/FpGqhmx2e/zm/QayXfI1ScER+/Svxjr6vvAGB1Grcj4UU/u/XMIdHvzlZ0A/9r/eB8Xkl
aQZvp9G2s/L//sdfDxhmP+oYfx5U1UlEEU3pyjDLdktEnMfKzKAdCGjipP2cW1fNuyfrVZfIA8MY
oVMOsQerTbgNUWTLO+Qt4tl+DjUBgb6YeyMq9q2sOF9X+USRUBMM3RV+gMHfvozZljrG62Qmn82E
KQQF5NvVI215mfwviPg6f2kA250d8H+miZzfx6/doxHEWAUeOijTecU3OIbvAqd/XYEf4A5A0ziN
jkeDGjr0v1SkJClSLVxKZP23CdCfQVDXegpCR1KWq4wh/CdGVaCxim61qMwDW/tUT75KNevrGcxZ
bkYYj3ccdMNnBChpxPvn9ZQJ40Cn/9HRqDOXFEwi1rHfVSoDWvLX6u9voFWVFrXjPmrbTiNVRvOa
agKkoAXM+wEBUKdJebR/Sc5uyCuJLD8wkUeZa16qDSt/ZWpVmHUACVWGPj3zF/EJ3B1VIgSLJHx8
kvHESZfrki3K4s6wbG1gAExBtGreXOFMTqIgZwnfZ7bAzElJTrabx926KuKkZZcBPUZ6VBSojO44
wu5kdJMIRvybdx3qo0LhX2feYvU8dnGoY8CDfLUGwBnspLN4mSDjaVp1obS9cuY1OS8vtuZ07b7Q
8vh1uOIA1zKIm+jQsywYXU/5bcZisyhXKS6WkkMr4KpbcBm3M90Pepw6mRqT2pF6SuWD+gEAHO7U
0kZXRnHJq+5hZGLcOYTVyMLPtk3ZcdeWRnivlT7qGPwgXyPiFaDjHriLo2PS+WcHVd6oWyR+lkfg
ajbJe+9mXGZU788gcDKHaIo8/QKLKqu9wc5CDeJzxlIE4P3vb4azfqrUdFd2RrqtNX0vzVqJtkn5
93ja6SPZ9UCVtEf3akecyP8AK7fHGTIw/miS4+dpJO626ZUad7v8S8zw4++db5HpBy6EGtNGZn/X
tToVoXKWvSwn2Oa/6nW3HBA21sTD41E1GG2xpcubNLI1eDwhY7a/ta5Gd7bWLVM4erP/Fg6e8csN
ShPBQ5Ar+hNP2VZy0CdIHxSfTyIN00QY9MZ7w7jp7x6ITjXcc4VKrUJsNIS9yC9MrdVEbL9jymHG
jdtEgN9kiRFSE3y/z7wibk1O58DDjo6+WFDzVJoD40/9XLakuSPbmlB0hBrNCpKsyRDo47VNP+ny
L3O4nr7b8ktg9ar2cw1HZeMRmdZuqUK5nQf+h/YuuaXzxIfHnILAVBUEZWGOoXNMuxNlSOmk2DPi
mYvpvJ6yq/fY1bsg7+pYyLwUAoiUt1Qy5jq6xosaxXecJ5h8CWXsdHQjlXkcPqdwdccTfVZ4iEJq
wCIKFyfxukF5Flvcyzy6VSs0Ocuo6CYVV658aGmH4Fqzym3q0+8Sb/VjcvPhOI3JehawAfkyziQC
q9r/8NGeTn0HDbfulL85WVtiybnG4yGcnUE5tByuq8bja1wTk0WpVeUj0DPvb4yW5jPG8hgRAyxg
cMtCpFsmhKSC81mvXap//IzxLZI+7d992IomzmFslNjIb81EiweLXWsUTzmCR3sHeCoBDoSbVvDL
ZeWSYaBFPEF3WGf4x2fOWkJgnxMLSpOF1SS9x0qSOewzdxW+XnplS58GWJlwpyubU3n+rv1ouL6c
pUJXWYRAp9KLLamoK03ULaT2y+hRQTD2pLtSGAX6hpHGw6ZMbrdBrX4AbtlZ1gA2kE0Igq2Q3Ui0
fJ7VZ9Sr9xwq5B4hjRgWrkhwxFQ66JDRubzFj+puGzNC/skK30QUxViOGzZJWS4kZ0ouGtO4AIbV
oV5PxV9Vk9lNt1alwGwtlk28KHp4Z2nQM1zd+Y7sd27Cj5wMsmWp/aGEWlCxtm3sGHdf642mC4zS
UlyEkI5e1aOxnIlLfPzeAF66D+dTXx5e2h6NvCII+HC8CWNWPA8DesRlUgWVphVco7aFieBWWXit
fJo3JLT4OMhyIPoiYbTRthtsgrpyTjfzZHlubSt3dgmY4rpLlx7MhBXDJDE82G4xtWh/5JlTWLli
6YzHgVpTctXsPBwGlRATIOU61cpwR7uTDo/mP/5599xPnBcpzaAXDSUa1tGZ9IrTqsaKez+URBWX
WvMAPybvtxiHnQCx9C8NmbGgNuSvNRy5tiZJFf+1qDbVoFHVb8dIk5kFZytFTID7gYiT5UwdqAUL
OC1yX6u7Vv7dlrVJbfiQiSsxB73BTYbLBEunvBxxBr70aZq8Z0182ag1xK36Thdvc2v1Pizpjs5j
OLuqBkHCSH9kAuxgy/Kgwk4gafeIBj/T01OBjzr1U/MPLgABaGpP6WsxFt5cMTJUC69tVA06Y1Sl
EQvT6wMtdDURHzW+MHP5AcRBtuB1qutl2+9LaO4FOdg4N7ds4kTMWV8i4bTXnvNQGxrA3XSJ9gkb
puQAfuYuX+2i9qzrK7kGcoIZlaGciC/QNgbue4ifB45cSJHY6LtUvk5j9+g2lJjopejRGSZRND/k
DjwiX6Jowaq5PVT2n1Ha+9iX6tDs2a8amXlp8hB+oCzcZvHYjeqYdwuyBARw7Cd98RU/4XgnC8J6
pA1MfCc913FS+PS96fZ4P82R9qwDQpuC9Fl+lspx3udc4jwG2W2gNGc0BIO+7Od0exfzwbgF//NY
8C3ZPm2ahnuSVsyI/ttmwe1AUxQd1FXzLPrCf4STMsdoH9TJbujZbUKR06XwqoPf5IC8e1lDpJOf
xWlT/bCliXFLNmrmWh8xeg9vZoe8CCNgIoVutrpAnL+r9QkopBk6+3Jm6Kvfni2w2PAegaLSJsMJ
DjD5E8lFpOhPuO9fHZ21Xn8jkrpTT8GM9ymBXUMyhCWI77V+d8VN5muZev5nn5/R9BBTofGHszqG
GIkk9iq43DfG7UckCFqTbOk3jyDvPN8B4KGVK9zwHDSh345h6Tseg2Y3qn1Q8y+PSMYOtgGyc/EQ
8XjSWM8pWdQEkkuV4rAhqClfsUrb0uuTRulRe21FpanXWoosSSypAVktpRzOeEPnixzSw3qWo6dJ
BJ3ibC6+6r4UZ9PQlJEYZC6CGLQt2ehVWeiDvYZtw0hdaZH77FXnnURaRG1agNqBwwcTtESeP3YG
py/p/ZN42KdtxdGl3WqoeW4LrOZCrYzzXz6t34WxAE2c5iAftiAKs9zVkpPmoaXLEyL1q+/xjlAv
VZv1Par9SXsILzmLi2MOnxqPBdBRml9ebTqEwqDJzU+TfKjU/PwLHpJRC9Zu+b4Y6J/3UIk2byWj
qEvbPCKjOZe1vnW+EMlBwJhJhKKZv21chqnmQbqXqvmI9ZXkxF5tsezJ2wHo7rBdmWU/y3cEW7CD
XuOZj1QAJFC1xpCQan/7965KKhBSRTAXqQhfrzfCHaxP709TP/S4YaGCW0PhX1SrO6Gy8kPmsLfR
a8g/J7zVDVqbY8TKcVBJPeJDMWlVcrPLtzwrw4qrYRyN1d3x+agCGFmxMPcQqEpgY13K/tX1A8jS
cka5xIXdVBZZ3UT6bjZVhsDwW0S+mXAaP3Wn3d3ToqCkTwDojrULVMHUXv/LD0nYhFlWxFIDNXYA
USK2e7k3KCS4hZFq0F2PbWcg91lb4ZdYqELLw8c1r1pg58+7OBhaDVhvrX+WbQOmkXGyTmeR7K7+
V0RkdHhj7IS7qcWZtpFWyx1ODRQNL6QIbVmneb3JahFQCvn7bfOgvVMKAQmUPXX4XVZd2QBHyCsk
GbwC9sC4c2ihNmgGKY6ncBYu/hHxwZCtZDAKG5+d2nWnA9LaBMnauUaGtkxXkuFdrgJJdw2wcTVm
AwH86EGlcVXWDTogE4XGEpFo4k69tnAKXjcU8DOhr/OMZi8ntj0r/eVYRUZte6AAxFndoxfG0ZHa
Ii3IElDnIZ0qsPdfMpCEq4pcTu42m78dcjWEZvfpXzjd1LBYtjpkHp+0NHAMAie82JHthMrVz+6C
2peOppn35Ff/zNKrnwh5ERQJWx6s7p+DGzgVtJU8h+4WmyWMXAaJn38CgyhO/zEPyQF6Uk7/YLKC
AT4EleWyYk1BuIaBkK3Lu4Ozm5iovTraM9wsKGpF6lpAa2kIweT9pYKzhzaPglh3J/A8NOHoRNe3
H9sreNhwPtlV2mWRafKfv5csZ9sUE3VFAbsui62mHFBmhTNXNeVdG5LOjlucb1QIO5GEt0pHQNgu
3mqEX0CuGp4jLbP3uuoP0nTFllLOnVJbarbZq3gNtMsl3WolT78WDzX/vlbbGSRDnHjH3jWtH46d
Fd3RWVQ0SO0preuafTCWqLxnYnHlzN1bbhtcHh7me6+5GR4dygXJ8ZJwDRBaDr5bxyCMJhSe18pB
4JJc7OJv4lgdH05fy5k1wrRJrL8WaAbXYI6dK1gi/NjIDKhdhxaOW6KTHovmrC2TTcHHKQNtIO/V
RqMzoiSqvxz+pu3c1X7i0c9+bNFF7/Moc2fiTHnFhhQvh8MMbwPRbMFPbYwKIr9obMLswJnb0Oeq
gEBg9OdOIc0XSkydG80fPQu+S9G2UwWIYkdfn+pF2RZeklog1azA3a9dN3RzRj54+Jvc6Mf2O3KT
fHDvE+UKEeGyzMpgfzW18UJRCYkcweXVa8pWOVTSbWUtIa4h9xFy4mi9313BlaMsYzNHlw33cXY/
usNcxqjcTJlk8cBfhJB91xr5dq2AHA8z+BZuQV9IfkCwZJldqlO6HnsEB2RxavoBQeUWqymzV2oC
oGnXaZDDvE2a/IlpGkVDF9Rm++7zxNxKh5ic92Ml3PnYpPBc0qxPEecB75yuHJmnxNRPN+IVVRkl
+gcAcr5ub+k+bgy1K9vnFVDkXlYNWVHKhbTkk6/HPRerBJi93VE7l0hsscH5HBgJpllanNGQB1tx
bBDLl+8MlSLPrLxVAfzDLd91XTc/4wuAdmxWJ8Olm1JfIRlBoIc/59XueUj+/GoSJa2fvUvvLSYM
WCnniQhOGDR0/2Jr6Zr3XhWUu6aSCHHGzlAe5h4Vd/l7gLfXn+sspSzzwbNaIIa0KCNRuadtsgl+
3i3iiyP0RzND+lL+vZbCFOCowxLa9jGIKdjwg+jtyO/AMo6DoYM0iiSYctCHFY45JFlMdxZskVvc
fzln5FrPK6haVYTNMypNALqgMOYmRWnEltGHcF8QVzfUKeEUrv/GMybtU/OCx27zU/2O88SgJVue
oHtSAAJUFKyANaK2H3srpgVFNN4TjAOaAP2TGw23Y1FtQODXG6SdhipVIAhHKGA3IMYGBbLpAsPQ
FEYwawLSzuHgHEsd09HxVb7UyEWIqJpqQf6MFytj4hF+BF1OOW3F0lH0nVQN9NqyM9KgEvwNZNWY
baPHfKbx5rKklGC6zMruvKCUCiovcobu3o0wp7GXIjVDYEQonifbA+AuYXvE5bjH4H00UrBv5G6G
EZja1pCRehZ2DdlAFgn09Q5PoT/q9XnGLxj257mh2jRf/umEbNmP+TngYyZ8fxUmAtfiObtmkjn5
gKrVbuvn+hr0FwwVMK+GIj0hosvloKCgAdw7cuhOvrYqyBFKEJcjBWeg9M1VMBKrLR6K811+vj2N
XD0r/JT240ghAlSZQbOrDIivlxRepCwOJMZxPT0shaJpowAlPdmbpuY80BLEr49coc6AaNO4Ce3v
yt4YQCwUe1Rk+kxvhLQ0b/Om81p4WrmOZAceSKWFRWdzzZy57nOaEkYn1cSF69wZJU8Qoka7Nzwo
Oy4Yw5DIyT8BvzGxAaFu+Voj/Jul44EGNZxnfUY+5ARkuwUKasIdruffDUXZnku8ddN5XY5zSZnp
aotBWHTWrZcs3ZLs6sALRGgS0MbCTNcLMa58Kb+pJgpZWHRXfhgDsXpP2AfY5o4gmh/NwTFXumxP
JAdVwycb0kAA5wBzbWGpE1AlNkqTrv8JL10FfIl9UFU2/xse1pKXHxcavp5A2v0ZQY4riNWbdwC4
Qjuf6iAN6oQt+ZwCyYI7HhO9AgQYNKpfb+uLldudnWn+MbjcM5MjM/qZb57nfjAuCwNzgYQ0CSvV
YvBLsGI23WFH0cI0DaDIn30BlDA7DBIU6rxEphyICzsJm6424JHNAMXMwnGu/1+fcHF7iwpIp0vw
iehLpdnwqjtvVn85ktBjljNYAkARxYAr+3VliV6M7vHFZ7nVfONkizIW4Rhiw9FtFGzxnpAmoW1D
5BswB86SjkOym0nEK40dkz1Z6oo7D8u8ZEuE7chT35Nl0RuQAfPnttOmhPwuT5i4ho3VBdNfb9TM
djMyRCCNqViER1WbizZjJ9Bw2pVun+1vuZSwkey+gq1f6wh5evVEwSSKpL+dXGjrCZz5y0mbbl3T
KdgERDNEai2Ex9vxbiyV1w2UqWFnXpLEzsbezdxRn0uI2mqBFu5MY+Gmkok/OE+Y50h1+f83VSB9
/QcnQy6MlfSA6lDLXoSHF5D/xovFtPZWfv9WJx/azDzfWf6KnDi1jN/eldw1Sv+imXJncL/udcrA
zsevCfpZqdMg5gIROeMe0P8i5ge6vVnlyzctEYR2F8LY5R33w+rpFx1dDe9UqHBPEHI5VLUX5+ct
izDTykRZxikNNrsQZw61iga++HtEQIFjyicDUlYWpLv+GHetUuINApfKwnvGu7w7eJgIQQ4T8Vd+
TqAebppWLkljM6+AqV6mzrudN/4EY4iKjoqfk6pKuFtZ6pkHhxKBlkXJ407iqaM4FNFuI0Vo4iaz
Vwesc9rcET4riNBsYdPtKiWI9auON+OpSdkUZxrO/UtBaKMZfEDgKuf0FfZk9dotWepnb+mMVRYU
vYVTO3oiNbqL67Q5TDBSA8+TWrjXnYdAc5Pibk2i3qYEElIPktGeVfjKaKz4UU3SamKCkFlL0qcy
T6DbnK8va0YL6IepzG42rbFmk8p44JOVNeiKIvwrtCg6WlWIfE0EcDdxA2L96GdY76q+ASjuCHP6
KMrB1ME1GJBU8Per6mdK9v2Qh+RCtJjR6gQbtCSukmJNhhDxc6/4+8+7W0t9bPAwccB1b6DheFJx
BrZpDpP5PJ9gKFTAe3qskyQnMvAhxjBPC9wr9VwjHhMLvyuB8YghNSWN2Pxh3apk6//TSB2zPgLG
reN8/2+BKoYiNxSELmbptU34Ao6cGjddAhvL9N3W5vx81BfYcz3f93vy0D9SbOHDb9+5GWQ2DEIi
I6fYGzCJjybAUlHIkxkuzfJXY3b15uPEesdCcC3igEj/I0Oh6BVnxf5Swsw5LEM13PJRPvy7ejHe
vbPfmK6zELoS2UV4AzmyfygsFBoBM2DEqD1wuDWw+gtU4fnMq97ePm/xuYy45xkrb91UHYGnD3wJ
sxAISyQ1G1s41IsdKwoP7CHUoU2jc1s3DtxnWdtBsk8BEzYEtZimq8Chi0EhCwSCIQ3sZvsa0a+8
oHOG15PeMqUxyh96fRlp4nkBdblqCQSqDPi5VTBqX9KbGPGG5489LbqM6pWtY1janIE2Om8HpK+Z
Kk1QxdQXuvbfFAUdRJZXd0DHIXT/VyjftyO1j+1Qh2BNS+6GAUzp6MiK57HrE75WxUjYHPKVCwAO
G0lDYOf9W2Aco1kCMFFhaYdl6edXKSYDTBUbc95XojczMxq7Kvdmd8bTRiqPMKLcvzLtWNYFw3aR
+ROxMxhjUU1dIzeSSIONZV+koR5jrH72LH+Mil2c1BJgzFlZvfpOhuib0LdB4GeS1oSxL5fc08uB
4JrgNpKtXsdk61ZXX4kP3IuZJdU/8+b4Z3VuHCA/lfdp7QJVrOlciXVQ8xqNMG1VVWVWkvaaEah4
JeRqH9Pz4kvMH+z46XMpeSO7690S4ZtfCYkcNKrWYtG7iaBPF7hQPSS/DJ/e8OVPnpO+mb+UUR60
aM5/BxyCNo8vZQIIX6TWovf0kt/EO5ucJBbUpBriHF3lLc6HBDOoSFohf1Zwl/anzXqCBEAln32A
DzQj35NVveKdra8prqSt7PKWLxKcv2UPRcQSwav4BGC/UFTh/t2zW50bcgwQxZge++1ExAXCKLnE
O05t8EEP5NRFm9t5dn/XUS+akee6yCaYm7KwblsKvyhqbzIHdteeeZshceFMmCqKc6NulCnD50Bs
8v+eQl+ivUt7U1pAbRCPL6CC/HaWvPDzCod/4ZfD8D517Majl+/CvrgfCEyphJCH4ZmbWaOjbT7n
r9Ar+skQLOOVjd+P266A+oWpsgAl0DdlV66QGZecZXyG75oqRLdpsOBKjXbSt635734mphRLTysY
7uGVXlkre2lmQFO5Yl8EeYI8MTTSQqwcelmFZfHS+OFSpqOwUJlLLW/kkZkGrsreL281KoEgzjcK
mlDuTF8ahAkQZuZl1nXwawYe8Z3tYrgJoxJQTmsadueJ8Gm7vMwSvbwyE2b04VoOmMeZDpdgodeK
xHLs8HjoTJH+/QqT6cPLuZB9rtjee/sb/ot1Caq5JGlPmGW1Tkis9mIwV8Si7flfoAWvPK7uMBNf
ma16zePZVzpHIzTTF0Qz5xpCorhG61t9g3P+BeaovsmZ4l2fL4itEpyOwZC8glfWV8OksMW5Bo4Y
+HzI29qieA761ei4PwI1hFnL5YdkbYuU4w6lOU3NjiuLpu5o6eMSuwjtRn4rhhQ2CBIhuC9vKo+F
CZA6PN4g1UNA87eYXa7DbetLcyRxP7hMkdmBEWx/ePQudD5X/h+j6MWFt8rJ96qhxv/MBZlnN7IR
wmx6+mhmdlKEoR6I3+vRjXD5bAg4yNLtn2yi+PAXcf7zYIZll+GLXD5/n+etYyrxeACAk+SYfPls
+C8nI9xA39x4MERZ57Srp6tYiDB3Nd/FsZPvdh9tcGf4LX1+t0uJKiDfrNsl2wa8AwiAkhd+FS9d
lVncYm60XJo/FqLbnZ4UI54shYwGyvkKIBgxCGtXJ85sMK/FFS9cEYg7XuIej+kIYgqZMLa4wgsb
+LgMpuUpqKNHOg2/D4SXWYPzpjzIY0j/aoaTtZLYoXg3hpte8NF3qqqR4uUZSE0zm9UDbjgyx92l
dLoTrDCYiO/Iw6O+4Jgv6oYesnMpGBsdhlmpzfyDmtHH0/VX8H4qeNgf0s9V60CD8bQBHcBX520P
dotXihtXwa/cP6us0Nsr7SxRFteCztoBU11mq54E2207nhJqOdrcmWtWbJtWk0IjYxNxtcI+GJz+
XGNmh1Czh4JgHtqjW5BcEVCvoaBpOel82q8ETbnb5OxawU4ykuQsyFV8ISTn76tCwVb09opzzzx8
wdO8k71XK/shrACbcFuCpo6z5EyaSH0hXLzhZW8QmL6oFx5ZsQa6pGjyKfq189xcbjMW4Z2HWu8i
uE9JlIVRJEvzgpfBNgVU+PbG66yCexv9FfYnLvyWmdQhVP9BfjyYxRLYsBOo3IOww2ELi30ourKw
Zhx3+XYr/WfTOWkRn0sbpz27jUZy4ldOGbjkp+heVoxhEkOx+VVEIojBKbUNcDrQdtzLlKhLA8wj
qeyOJUfJ7/vyIbzUihQatRiekDXaiOIVp+X6LvlXKdu36ii+LBx6hcYj18u86pO+st+O9Gzb921F
6M+Amke9kkjrQZqgX27jJbmOE6hR9+Pz04+DltDVHUNrcnse1wpqT6OLsNZgZKZe7cyF84Q0bVLh
Q76YwyxAZvK1rRrVCuEHFjs5AGtOUOjkZd/LJT9umvTut8+lZtQRIihzaBFoSb4lAMe7OTSRyA+F
CU53FvWI/TaZ1G7WigR1an84ZF/mpraJxtsnj3rKV6gbiI35yfnIpKaY4hTrzrni4KrCjGgwA98R
w0GX3grlgZhDZztrHvXUbukNx3cL1+a/Uk6y36PRQGT+mCze0BLuln+ZSGleIl1KVacjqBW+AIaV
kM2BWXSSvBaBQ40AqXR7+wXo0lxJ2/TldL9uC221hUiHJOx65oU/JrES42NfdtZkN0Fr7FixvBW/
QWnolJWzvN7NouaLR8hEerBUNovH74jITQiONzGAEooSPTY4dmkY0FZmJm8I/McC/z5a/PCJ9zP+
mMR2Jem6IQkSrt/iamEPIta3Q45KU4M4eOP+o9WqtroV3Og0AJXz8rXu7HShyRkZ4R4S/u7jkfZ4
SAyuEhg7kFcn9irNBzEsLFjFKHrEAhDiwJ5AzhxBRpBNuyWM1yk1sV+9oavJyEM4X4gqcOVXMepB
w19/qnOabCr0BwbA8YsXIuS5WoW7CnVl3znrl1dn3vDKj0wLbrEz6ZgkmBWxcnBLyacQUaMLU6Le
rwgaVXh6QU9IZKTz6A2idhNcpKXlFOZvQPFeliGnWpl2ouWcphzRlDHMYM5IbFTxJZlpzqtXzVCq
//OedcZJ7t5MEf1Ej4uWRjxXuhBV4Xy5X0zh+soyuKJs2CxZphnVadBA93e9rTOFNlsvlJyQ3EaO
qviNSJjkj/MnPR/bnHyn1t8JxQM8obuNoiqTraI6wmAdNPIkR1dg/ElI7IeaIdXPYoEHzrWk5AZ5
VjesL4WSam668g/ooVCycYnvgP86LjgI8hVypVivX7/HD8B3/rs04w8cLnP+Bo4jEd5KYF0A12lo
2OTgWydopovv8M6xPfVNbVa5UIl9xZc1XDVSPdIpQDRnk+3++uaY2m60dhI7mPtV13A6XbaaDSTR
jTneRjnelUQMJbfL97Yeb42CUCBna9A9rWksuyJgNC36UhTyyG1oG9jfcnSuE+8ncE9qCTQVWwbT
2AJJtscP13oeQGedynlMcP1J0Ir7cRpJcGLK8vVVDxxJfjooKM4nXfk+49AVvGChSKwt1kgsWAUc
//JJ/T5jAfDtWiWaObXUnxhjsYf5+DrFs7PjHJSdqDAeAGyuPQNWftubW9jjfokhi+yjtSRBBavY
ZYPPwq4I2dl8k6yQHkEnHVp0JdZnCTuENkiG2vi/c6p9VLaj34+OdQ2j0u/c8ueL1YUtgGc9oYy0
Zvy1DvS9Bym3IsRQ57PTPXoXgyRTRbCt7+NeWyQJh2GMmGZgR4YWYHQQTkTkSZ8YG1mwVj+Heb2W
Cj4Hboa1W9zkDfTuOFvGohrrLF20hQoHUt2i3fXcB3QWInhl4lrkFFJzpJgDGY1f6+QSzWQeJ7T5
/NQxmwkRBspOhh1Keigc7m3cjdMQhMB5bsI5qlhdLAYeKr6Jj4rwRjafG3mONjLjJDiLdPNHftHT
lSlDUpStVaRTuyown8WMwsk8pC8ng66+bdCaMf3d1uG+IKsooEn6wd1v4JtuhGz45hB39Q/B3+63
XAEsal3vXtdn+jfqC4nrgqGwz7uo9KFCz5eYWPJSTYzgQhp0f+lBChvSqjavlvuYxLIBz54tMKj3
u0nPd/xAaZ3n3MKAT8cIprkDHUKzdheOjZ/ue7LtEtbjoXiuUSZjh2nIE9nDafqTeDT2nJMmikKy
pVzVygKRL5WZKSDpHAubyX9qJEdw8SkhomFT/UoJNks7wjbrlPuMWv7IqRvGd7Oya9acSGDIxq3z
Q84oIgyDBF1Kf2woKBRNmR7ilr2fDo8/kssOtBomhS7A2sA154kvU5g5AN92qPDm5wp/1szH17oh
syFu6XYZUDqk/bXm1FE7/VQf5RZCr76/H/L4l/aFPq5k7PBku0D/nrqcSjP9pW47ns/R/mfQhlZw
pvEFMMoBsOqDa7LwG/3jLA8mcCfGxQX1M64kjeTGJ/1CPW59ydd8TH+U6ybdPUim4LoVWTS+QDPa
9ye0Rn1Usu0S01XYcdjzcjj4bC9G1o7PAflodZYijVvFz8JIRZpAMvFmO7yN5MsfJT8sBsLjP9ZI
YJQ4BTzQfAGjVnKos0SXhtMJYj5+c6EDd7/fK2WQAkEKF7nOm80L29TZv2ow8ANpcaZwKHoHsjcn
B9FIRpBBSg/lrnB1CZhHicP673PjEQUXbkiizFOdU0COCjXxhCd2xGik+JiY2I04e1a/IKq/6yLF
wSbPqcKy5Ysnc4aBskbW4jfQeRU23L/7e0lSBCCINUFgca8AFgqEe9EsCwqMiaceIjIUbyjPJzOh
ptYNbjnkO9ZH4vV8HxejKmPPoAm9OCGaBLSNVLUHUWWu2Rt74RNLO0Z6GHfpI+9HgibmS1lHzMsH
PydL7hqBTPu5SFC5Lu2/MzjMxxg5xNSJuISqX5MOItM5PJqGQv9CKKdwRctkupT1VjqC6g/f/A52
vmnUNWYmCLHsKZm3wGRYNDr1B9Q9YMtrx9KEJFUoT/iqAwyOZRisMswsJ5LzoYAze9afR3TsxWVQ
RPCTlHp7kwgRF6hwbLKsm3mx54SQ12XXFjvaOmqL/dYcU/wGpq3ZmIiiBOP/kxlEXseuQxDFzo19
l+D6raLA/qbldFTFbAPwAjOQFKMTRzAM7KFJs0d0/gByJ2HqpshiviZa4kwKao+tRVLnX1n+3Du9
Rn74OKIVRhZlGHv4UND5Jg9xZfAcir9GvZzirRHK83hmtZmXsBQySB7hlkIdgyM7QaVdPz3RLJ9A
MrjknAkV4CljRWGx9nZTLxGCSBBv1oaI5i4ihgYFdtwT3OdEIKh+4D7sLJGAR55mUwOoojNe1UwI
ZrsypLuLk5IbfBoChlGr77PE5PVXGlrM3YrRgcgwHi8NV4hNYjgSXd/0AEbf+cWUvWj5HuRmHSfO
z5EZoXGKCqJqWFVn1TZfh9rW8SHr01d8ms8vLaKBknaJ6fCK+otLVLyNZ1TNW7Q2wUqwfT6bP+CS
mVSv2RCX2sGvmpuhAFXdBz/yOedxxpvJH766vouN9whL7IWyo9igK9a7bgtN71O5sE5fZueiw8rd
YIAt/tQJ+MFQehk3831YVahsUi4fdE/9t3gs2e5ZJ4//M8VvWSe4KrG2Lp3vj1XUk0a6TS5ucprf
L+RW/ilTU+AySfU03RcJSSV36qpfNmJ7mNa4nCfgKHC2E3cNf8JvS7LXUppsxQyh/0LNoLUjcmAX
2gUgOWRU3GpPwXnQ1DYGvujH+Q8bcBKPNPxl2gVTk2h5FiixaIXX4txm/Scgp8R9q4TQMG5/sbq7
wDZakMMuWtkvT6dxt1tpf5uGgoYpfRVPLuwdJO2Ob7aUeidBZ5PKE5onAxhxlRYJBlThzXTNyM0k
K/TNGuEo5VkK1LZCfXxnwDp5GXdQqgVDinJFivgsXoPgvm74nu3U5EixmH3PzaCxxYM5A2ZqGKjt
0PHPFSQoPhelTk8xWfxFZ7V3ZcCjy6pvzL2sy25jyVW3Pku+DpP/NIMuo+7UW13AbqHD2f7L/IFy
l9zMP1972hDMkisI5rrBltxN2DdCqIRoU682CPmPqFxRRizHGpdnAa4TXEy5x7zNh/Bird5N9d7T
iQebhaqmtYTEIHhTQnaY/NF8muV0jv7689bLijbQ7dxd2Y0vjEXeSQrDsuzJosEp53Sgo/hdBOtH
jhvcMHMtDdhNlXFFIGWjnHaU0d+HykbsK3i6XUGeop0YryIIgyAAhLgfGiuOnBpuYl7fgsPdJk+V
031LdWXkupEYXnhbjQWLA47IB1A8JKI5/cfN3C5KBDO6JECXstGHkzo1edzPw81df3lZxCF+Sb+N
wUkwogRZ3+rvRulS7LprVvYlphTvXvXGNaBD37pxv9uRYb6XE0wFkrqSyk8DpT4xYQ24KkzU28Nd
nu/Zul23628l1S1mj8swAN/z8DrcbLbxPqJANvzoTl3x7uJcOWn/OcViz6lL7oKQIaPvOHUBQAd7
vvA3bO4YBrB4LTaeiKesPTxCdV7tJzu3hLb39DFo/7o4pNdvoZdqFZ7T+/7/WPBoeI8wPIFijEgV
916pCYHYjhqZ9QM0q/IBtOm6okjFbv4T1v9jUcWXxg7/YKsXANHXC0kLrhITCZHOSsslia1r1KG4
BFl8HYkjg5sexcsCP+WDT7rEa63nZvrbuT6PI/MUQtarGVXqCGH3W7gXp4IDnu4Yru7s7PUyh7++
kftNCBVaWT6m010689mHolpFZfE7TIJmtS7oMPlWO8sK6VTPwkoluiQgI0iP0nsS+huxJ3qHx0UH
Y+8ii/pY7IRDDNVC9SEZsCSq8okEX2uUqdjkiSzyLJAIMEBWDIOhMvpYgGkZ3n8ctApsQpi/QvOs
mC/VkLxEKYt+LOdersqDeTrKSY9ymkku4ukLM/RKhwu31FoTBOUP/esLqSXZXe3Fefij5iE7RQoN
s4hAoW/ScWPXCUtTsjvYtaYRMHbPeRV9smJdTBxtoTcwrFXzUp9u6oBADVi2QfYkpM4y891y1CNm
tDSFXl+zhCYqyCQDfXErj7p2gf5NtFKiiM6FLvXjNq9PBn1XDXk2nLjSY1rEAB5l8HNSDW97IShh
TcazphuISKIHtXMmQrJ9/d1SZsnd52oFPaJU35Er+m2iv3dwIbm93DvPatimfv+SXyjYTGjRxtQt
I9wipt6bZY6Km1w/IElteQsVtQJtNse37CrjoMx5ZmiZtkpkYOztWEFqmOdUqy2ayfi9EkWFzZWk
lF+aoaQIOYUP47kNQY02cCR2l1CMASMV2W4tgLK1LOmACAeD2nXo28cMFudCtOg9QgdxUUrw/Udn
uANwZXDaWXfezr16aVxbKEsKL1KiSEKfNrevaN0bfBwEVe9nX0JBHGZKk95/h2oO1B752E0EO+uF
WZOakCMG1m1iiTy8rKvLDndXgbbI3uKNQajAWV/miLkwpC0LPR/vl8jSoqZC/maVKbr69I5UgetB
d2DgPzWjViNyPHbUybkl2E+272dgxIJ7w/KSEugR5Jv5o6axqshsrqLq9B2XpiSK1Grvgc8L12Di
N/13ZTiT3cfvaAMrjuxKfgdGsAcZfOUeaKXXeQ5rm5kqSYIUt/VS9xw9SwEhtjW6DX5NjLykmfv7
7NdQRxtq4zRtJoOm6is3vWetAhWgr9+67n4WAtuVk+Wb/SysEajZDAfL2b+AloqkaLuzHKdwrZIN
fXkyg+04/5ecVHod8XDDP1woEPBqAVfu0kCxlCt9hWy4xD6Q4o9n0nPoBq6Qfh28m/nlBBjtBZoU
uKPo3bSqi7mJZLsQmvnzhvoWPvjhJ9mR8upI4yjQ0Kk/QQO/kLxNbIJ51JL4fxG2KkvdobTJESj3
0rdbB+WSku+IKmf7tpZoggFVOhY1BudpFl+MqEDcTHjOYusjIrNcfnuUTkatPg+NFYUKJUEaqDqh
tSvyXEmUV5X9mlmzRcRF+qJL3k5bWpt4jsWwNmSiDDYgsqPoLlPnCn1YGWAtkQNe0iaIJygHu7dr
RY+CJq0iHWDFgXA7XAyVdIjEpaIPQnl4yJa89Cwshx9igzqela033I5N49L8jCPZGpGHqG7+riS6
DvzQk8jUoteyfKOYKhEhxe/p08rx8MJxJJT6QnaTZwfrYApoCLcjoS5Nb2WfePkjJ7WGaDhyGAML
0J5xxNkJNMUtWE0MxrzBZc18aQnx8TIibwMqzDoK9KNmwd8fQglj95cvCgatMyKPigIJPoiAzYj2
T/Z0vvNKW66Nha0NKelwW6aCrHkJhCKy9i0vTi5xQFr7RafoZheA/zcVSFqlQZ/kPUcjzTj0gJ8r
rImQhxigyd6V4Jr1z4o2s/zxUz/EorAgqqkTu5jkJlwkbS/rR4Q8qeMHLQSHLrCLdMtZ+hg155Co
g3hisJx1rl486LWkA3dJvDGADH4IJUQV7QVkUdwn8XNLp3WcsBTbMamCjo/XlZWVEv2tZ2kB+4SS
KDFUFluLv0W/Gg8TySKw2UbFnvvlI0Q9MvRQaFJj+4jEuD317xXjlAusZNlKWgBIREXKnCGsZVkW
Lc4n/nYHgZ2ox14fuA889TQFsrn74lUewdakoAv9B80fyMR6hiG7VGOIw/dALQTubpMze+XlZtT+
/upj+JZvTAC3VqRejmeWu7ak+7zTADQx6NIfOQWXTZ4Ot3WdvFT0+bDUvlfhNQXGMgchb8ta6QsZ
0bpB5XjXk2n9jTlNDIg6xK94osHZmTJy94OrQ/iD1pxQgwLwcbr5035etkjRTOW5atxP6GPYb0Wl
fydy6g8KZG7VJ4xxCoI6pePiSj01B7LQ//BETou0MvkIjgBeuuzdDLvvbYV0t71/KRsqZ4VOg4P3
ljv+i/owUaLB438zDxIpfSx31tw8LJw61809po7SaSmk/jEdpTMholgwzwrOx6Hmc6mQDUIqA+r8
K70+1767T4oWdK7b+dX/Ru0mBmRs7tfa8xsvsNvNxkBEq70INfe6qPv04/QDgw5v7s4YCwORcwru
7irnEhYtT/VICT6QM6OATP0kpn5Tnm3tWLF9y22/SBLOqwU3fWmK7/HJcsrDclXZK7mPBGmCZyNh
AHcOcdBUcO8skHjkB6s3PlF37FaiJ3cUZmUudHjl5Ica5IhxLqB4BXNRhrxzithE76mF8zQ3fcg6
Qvmp7y2BlfwJ9n6wqzFfB/LIXG3pjTSygL9Nkc9gcjITNhcVxdu4bkwl5TfEKp/+lwSIIUmXwpy1
zGfWwGD34L3ENok34Ka2ASNleDeX9++JLaEMNpYVLKmupPibbuqNu7WSo8uKBvcuL5h9ogT5p6pD
fjs7WsalaaX1kPVTZQGyL/adQaSfNgFa5+OydgJTD39h2Z4NTyB6sS6SukhR84TaZYg4uopLgBF0
IhPjGDZ9fcOlOfTxn9XlyvRRtdpejA85gw1sSZSNMkQUxPYxH+YJo2ZNExnhWvNj9S6cidDL68zA
DxD5QJOnpUP2LFmqKWIAGno0byyqyD28U36s+dJle/8rr7jftB08OmgyN7brLIW2gVp60YvAQoLA
rs1Enk1NVKZCMLudFxhyXtSxk2pY8/4lcoTdNgQTQoO3FW35wYRxRMqtiv4jUtLSFLRg5E3mM3zc
EOpSwizGMiCLPw+IB52d9/10nf7R8PXHwIr1HrMyV9HreQlaLSnmjcIRg5YPJMCr9o9USOllzbe3
HxQ4Qvc5G3SMisgOQ2iPnmazN2CUwBWLqS4dg52orZA11Y/M8IqlCY+PEhFSGEIZ1s/0hxk7W/A7
omT4EbgKz04HwtDloQ3b2aBLrnEvYxBffH95UpcYKR5hYrED0eehqEO/SZ4PsQ7eZUHZiIgqPZQX
5hx7Z9HlagqCtOq95nSt1rLtPfEbLR3E/ETplpL7G6X/rgqrO/NLId/qWRCU2Vh+OIBrZKwRhEly
UROpNcXjR9ew0CA/EIMZ2c9JxEmdh/m1UaT1Av71D3SjmaRGgnr+r4DrL0eOeFl1fbO1iGIq9VGj
ElNgzL7NhnoD0eNgDv1WGNyBqRZiKBYu74QR4dG1iJ49PmJ7a/VnnLPUVOtLNZBVVke+4a4wp+ST
JQDbLLMd3hRBk40YTZoC1rTIKAKSuEv68wGA8edQUYn1Se7OWvU5B2k3rIlCyiW74KND1SC0OTvE
awMjQF4cljs9OlZsp3+RGpoVc9rMWGZ5OUrkGzIfu4m8TmRSq4qs1mIUZ7/Hw2GExD2Bux+KU4k/
QetyNm5Atxn7IS2Y007Tub3Acz6rD50EmFq7wKkTOK4k1P0xnxCNPKVQ+olQt24fyk/uhY/XbidH
x9VNRa02wOskouRJbib9jAjDBOOgM4uVYyJN3Sf9JpvTSLmYkOfXAoM/Rl5UtrhU6CSk3/tUEejt
8eqfuqkxU8gze43ju9nRxI09TtHwHK5fEcqOf7Eepw6qY3yEgfpB3LZFcsswBWvB2pGfd46qmozo
k5Aqn9NOxc+TqHVufAqUfsHb9JhPiM7GHLBN/KupBk+3OEC83U44zf09BIWla0lrLRiM7TEHSzpY
0dnftB3YIs93eKHRhzvBwnEJG/oF5VN/GVFefXK1T9Ic+mm/XrUx2cWYjIESBXbKvx9d/zKDWh/R
rbwN1z5Ota/1E3NtSCXB7yixOL8LLbEZkrN/y0GEoWNo887yy/4rxg8X/oOsv3jKlPx+VbAYUBH9
ihyfh2/YeWgaGWgYYVzVPGy6lqcGvY2tNeMlE942oCsX4uoptDfUu3PJ27OiDDyjF+iHKRhPlVDk
Ks5uAjjKhT4dis3VwCPy5q7ghbA4fFGW3CyAMqyZI4TI458DrNmo0AM0XC/f/aRJ2J+uSA9K3Nj3
e/PhJfCyss53paiOjz/Oi5NYlC02pGbSrfopYsoW4JXZZwLn5arz0OD9FGHFqw7Zk7tX5iFe3aKw
FThHrUQsiCcmIAvKgweaXqEK1YbYYIs6YW6UBYbH4RzOQX8dNL02v30BSOv0sff+huXIsoS+9VcN
oTacTx4NoQ77RJjhUo9dM5OK7/oL6HurXsPUzGXVmuyjCTAYkqu8SU00ogi3zm3+joTzUkPKZ8FW
VogVbrTLhYPXE49FD8pJG1+BZWkx3IdTL7SkpBdtw+M1rKl0WipAKaTe0RsJefym9SnF6muRBzAT
Eyh6GzS/uvjPb75sYYkVqrLTBrLCVtgzuKxIWQqclb6XLR1dT188CGwAld2x4nD9TuORVRL8GXUq
nJRsc2814aq7nsUb69Gv5nEMGrz01veWP0rTVNB5i634qkDQ91D9PTPP0elDNTiwgbdZ98sakv0J
jY2IPcVvHmhJlPuK0W8cUKIHW5ulBRnfmQu6TmyQyS6D3PfhQH9u7+2km4YIsPrMUjpA25R9uHaE
sCwSJCUR9EDaGKqN8YSTS947ATcztbKlpBddclXnux/WcjymzREikGsSdF1nVIQUgMHP7kUr1Zdd
XNlW/eh9TxbNLcrZktE8tAT7O1s6BzRl7zS7v29MZiACx3QaZZ4ab83CeWNlqsIZ0mttyDyLeTAC
bYGf4acqwlg/yeKwKYkqtB54F2mTm5I8HOTn7kK6zPjWFl4y9LuhpcRvAEeJEYX8POVbgqaoh6Oa
7VQTulbIDboXd5CyIIf0Bd8UMW34o73CumV5ad9Z8I74qI+pe9JATAtYVRtvylpIj1rOPxTeYMWq
gGABC7VI/PkP1zxrDXrNoZ/0YM8CbEcb0p7bflhnvtFayri0fAnDAYKYhwPNTHnfqWvpqj05RGzz
aZ/3VZJ/mfrs52U3Nj9Tzi2ssgXF5xo9oXS44iBYXpqYsqO+OVZdNXluYx+HDCUw70pofj0x2OT4
m3V7AIBDkApyndffEUpIGhZP476RTOBtheRqXhlVbrWC8AE1mJ76hPhXmJ8ZuPr0leLnzc12i7Z6
8V7clmifxvNQ6bwmiJqiMMPkGTu483Arx5Rpdv68oZ74++P/Z2tuGAuo0EwX5jE02iZOdQedgA0p
wh9ZiR1RBBkpDOeTMcMRPO4ZGluZEfmlXfQCj8NXuZh/ezkWny7Xz7F1Y44o7jxsbynosOBsMi3R
KqOgzhBMFcUVhFFi5W8Rwq24JZGLwIJfGZOef77DdAMwT5G+n0yzZw9k4ka8SgShoxfVglPMLAtr
Tiku21M0HsbSTNXt6E0n+QaO/pE8u5jhxptNSnGykXYSKVHCbHYJiSWNS+biUqxsqlsIDIzGnlCr
CdetxuJV0i3xyG+N0U6LkF+0zr5tgfWOgJwXaFFSYnqQ6vq/I7Kwfco23zJgh97Yb63+c4fOhZM1
9fL0B3UL7GAMDqyGOxz+tMOdY8Puxd2qQvmsyd4HvCRJwZ0bnYfDW5fM6IwytjzwRLr35o/K76L9
uYoBHnPlT/U3FLoYQNZ0v3dYj2paZfCsgaMpxRzOPT3NL2TBKxVcUChR4Frt7zNlAwov1j+SeGek
2Qv/nSncPYXH69bUlC6Pnrfy0j6rpGtxOxn4S6YRthn+wn+OjncSUwlWrO+nVeYFS2gQEgFtQkYW
sPV/umuZBSwHODHa/0T/rw1fH19dUYbW9iIMlfmFdtTgWD00Yt9qbDgwS4Fh0A0qY5vhcxCJhw4s
kISxQ0R/Cf+QO7hVo8Zhexnx2P74wdN0WQZu1SV1ug18vTogddzTVjI4InFAdJdYen2vFH0d8vSz
HjjR8bnYc6dMJmMvxkeqx2fU1mSDzVHR2f+5t5l7+9Si5Aa+MBp9nHFW3CWVQcTJtdxMmXR0TMeo
tCdbHFByu3qbpz5xFkl+z3KMhUKQ2zhSLBNa+Vpf12zTjyJUJ4iR7Xo9Za4qIXirBusm5VrHQ13u
ahqx87QYb0ulcHxmdrh8i/rpfanzLsjhbe3t7nS/aBocc/cCRL1ExSASfyf3eyxHWxaYCniAWy4W
84LIyYE0boRyePOce0meeJ4g+aA/gA+0/E8+vdd9X4gb8mJz0MgTKhdvFYPZ2JjVe88c3O/z2A9P
t0ws5FoWNhA6UIeo/GissNO3tcurs/2T1QPa7nB8CYd1btu/sNVcIPCufppHirsd/NRqC0wJUxVF
xEmq7WWGvKfIKGtEfYJ7BaSlUDc/rwAT+tuoyRJMl7dNDGefnwNyqjgRYlFOlVTiQm8WcIMOnphE
pfTzoaQlEUbf3TVUOKRO12GK/UAx5BcQC1OrmvAJB/A3Jx7vilzcRhAkMAT/r3XEDsf9shzjCYYE
wBITZnkSuVKeyshlmm/sv0VckUlwJQjbpbMnau9ufw9ig0ZpqvremYb4OvTg1iqqWV3QmijQPyHq
TvcaxGuJfX0AMRwfMSO1GhRxVODD/EocQoSN03xoYDSC42wOdeuM/rCta/t8ZTj7OwKUToomJcI9
yv44Hq/p8sx2mhj4UB51nSLqVp7A3SgdjLXhwe3YTY9QRzy/FcuijorYGbzKDbGAe0RXmWrRYb+E
+EdpG5ZcILQ9BSEfNX/cxPFJLaSN45/FGjO56b9V2KX7Hi+4JINvpJd5ECoTUJ9v48oxM4OsYaSw
MmiZUXhJwJX9p7sLIh0fsWQd9J0vPJKMurC1JWxHnYd2Mx0XIuFEcLzjj6TFfowDy/K4TgOk3ikg
zCXO7gqcWWueBxJnuSIMDlNyjqQcjDLmgZpSrxPhdgNnthPg4v8nOockNct3h42yFTft33E6/c61
rEW40jK8W04a45ox6jhNrISdEUbH7jFywwYajkgMGjx1BsseES5WBbL/O+xi7SEVF1DKS09o/imb
n6xjp/rZvRIrwURGWOObOJIsUfSy1CfyMZcJfXKWxlL1ynUcq5wM8oWQsSw1vBCN1XHCjBd+QovI
N80tsEj+kJZfvoCNCiZh0YX6S7Q2M8goXfVNrZowUox+WLEw4l0fYVpfOOmKC1bE695vTLWvoYYp
IStxZTRLPBBbpJnYryQ4wdJFXq9VpcqDKkDlk/fXatFj2w1hU1L0SZeBDeKSlwaMUiTkGzWlw2s/
u7sYjGk70nF5aqNrZ5akEEimRDH043pjOCuhEFp9QAOqoprwngfKNyLcfS/TTBhIddsEYaZsxtxm
r3CkeC391M9be1fAJV4CIe1V2p+GPZjHJB3dFYrOKQswC0Irk6MUZHf+Wqoa6cXPGcg1T6zJeW/u
PXELXV02HE8IDxqqlCOl4rYuWPj5Prf2LAuTx0hcbbrWNFxIZSqs+EXmNzd9xLRRwELuoEnYIDf1
5QJ1x6bZ7ai6gp1D1mMSht6Qildfc5/yJnW2g2IUC+PeJKdCMwTGJqjJaR7pkU97XZnLXwkFxMIR
hXZDeU4aZ04+bpN5zWSzkY3p5s4hOb3T6xg+
`protect end_protected
