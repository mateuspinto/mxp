`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
qubI6o6XTbclxQJy01edKsq9kVhVjmu1w+z0Fv7kl50m3Rku559TrxOVagucHdQYBgh0StFf8fIy
sqyecWkMaN6DYrbH5CkPbhz216qsSaj2E5lhwpErTUBnB+YEoO09PWWOIyUgOBuR9oBQmkjfmBS7
QJUhtV7WnqHHcltPQaC+WCItrGwg7nLJ0WIy91AJq2XCdu/wCK27Q5//73hhoQB2hqwmxFeYe42W
bMBCDZwokMXW1q8N9zNOp+pTirJ9FM47a/sbuG7mbhK/VVpcnKA2ztYjHdjKtCnxXPrxBWpGJ0XV
j/6YIaEfmmKoGqVaCbKPr6629rmqRl8HYuKLyQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="paia/dsck3hglMrtg91Q83JyIFboIyScwDTnSz2p6rU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 68736)
`protect data_block
fZi2H6xAdOkiKWnt/nf0sAfuOjpgKRXdxJUWd4C6/lKdMucCy4CBmABjlWiCchixwydVYLOyqrfK
9rKCs0qYZdBd1Xz6KXxxKr7zRLu3imxUdqA4q0WmZfX6gqrADslC4nmRG1Nwq7R+eOiRZuo1cQS5
N32A2aiAWivyaiMlSHOPs3AYEr3HHn6Wufct9KFLkm0s+atiiNXYiZU+d/iKVk8DNSCXppDa7CJW
IgBbyQsGZotgfUK7pe9j7pvzEHJzSJM5SoVlcnsVbsujiHhz79YA48ZqczKfRmoKUl66rZB3/qlC
3j9Wc8t3iXsXkeGdnqPCtQ8n/RAxkJ8xqtE28GrFF5QE5Uea0SJEqhZrkhTsh9iCNWE5ZPCpe+f9
G/7yQoDk/lx1kKj4flymlS89jJy2fWPcLcbDAi5SwpM0kUVcmlz7zUnL60SVe380pyNA/NHIa9hH
EY7ZCJ0cAfGA+owgud05bWtoMYtLDdqDnwniQED75XVomA/hnovY+dMZR8PfvjXDHkLAtjqOPZts
/ji9yZIuTHBgbKbT1PqJ7V5y1XZ3tCFm8csqY4tngC4wG0BBWkNQeFZY7scR+xb/j5VjFdE/3m6x
MTQqgBsmMaHNiO7gJ3+uQ7PSLV5bdHAwK+j81d4C/gQ8xGqbltZjT7Qu8TT3xsOieYhcKX+A4EIJ
dNxX647EW4D+vJsh3+18piGhCPb4uoo2cimr0pHmvFAZbKVyceVXQOqxlX2DmK2EmTS5li64+gM0
Zsxkzac6cCfPGDyIgDTcIX18quvlmcEu0dXbGQlpEmvnF4ntNodlq3YKpmFcAmA4+E7R9dTMUspC
FvPsaNValYl6JNUQg1hrCIiFunOsv6BWDOgh8U4qscju7Inu8V/IgzNnvwQWjSlaxHnmXlXdPDbr
Dh16Q8/6XuHNC05WWtVn/V40SJoBwS2RUkb93Szmf8GWOJVOx1JPHKwbBlXMSEkPSRf6gnMuo5yN
4uszRIJgzVQQMF5CvDfytUcVYPyuTPhojvkHSJKqVd4DHb3BQBo814g1Gwt1cNgmxZ0dUWplPIvx
1XPLmkeL5Xp5m9t6kbrdxddRpAybU2MKDTmTvqs6K911/nX+6lJ75YsmyKomRcZcAPdl+IpA7EqN
8D53Vp0ACjKGyHgKzvbzjbjA5sM56JcgfdEooD53+EuuvG8oGXJH5BoS58lJqjLCMpzbirJHCLr5
EOvUC2dJzL9QqPbqhfN8rsiB8Mja5YPI8LOfYdH3tbTSoVNlrLgltepR5PrayqAZvxCysprfv7Zx
hBr2tzvYyQK4lr8vJIQuZ3F+MQGKNz1r2nmilK/aIkihVJ1PQTorDsQYrUrwm1WrcBCOL+xrfuCj
MXljiPKS3xuRIXspO0E7LlXwkSa+OB+zp4lyTVlnjnihnf+8DPSZoAxew2LApWE5BX4SC/PNsOHq
mBffHFTOBUrjBJfW5YYQNp/FuuGzPpJ2OozeNCNrtlUnql2/jI3Eyq0pnKAbY7pEu5hJY8LEDghP
UMdzZcA7S2c/m4wY3/1ISeVcRIAGisuj6ddiOtova2HvmqFGJTF46f4UTdKL/Fh8YdzN+d5IjS5s
BXJeTNllqmT/EPS0nv4SoN60xVdFdhUTO25AhW10HBH6k4ewaD7nTeB91N5MQjnBpOU5kKYfRgaN
P1iksvBr3cKQiPYQeb0xyvOqg4JPW/wpIR5/stTZVuTOM3WR1Ma9oCs4Unm8puU559YAasPLi9GL
K7QZJVID/7bcZ2xIEEQfOJfo18zGLmcWH+NS/mOEb4y46vygKN4aM40GXaBRPGJzO5L7YeH7oDs5
4XRvvH4ZOpyG240ear6/BGkv4947VyhnnNqSxto9PJBlSYEa280cSyea+vJPMguqz+SNNNXjXldW
QrR01WaSg1hiiD0B415eoFzwn0M2/Qwvrn50MGWujbU5UNI9XbqQ6jPAmrjwTFqqsF6k/GFUCgyw
2TS0mKfNZqVhYSH5+hxRP3LvSirM7GDT3Cnnmql+YttOFGE73ccrVC5Fvz4Qi1Y8vWvuACP4BrPY
TCS44aD2UgBYPiQV1yaqIfnUrpHDu22xGzjiVeWuLCkj+ZeNPADUd7ZEXy3Mw2/nrjJ5/aapgLDo
FnHnqnQ0wS5E6wB6c58f9TLDfPsE4cc89nQDUGaW2FRyPpKt063cLAbvthKjDojR+d+3iGkwBaM0
BVvQjJqP0hQj14SlT4ANw4ej0Kv9RVpS5ELzofGt6JjZaYkKYk+AZgsXy0JIQmnNLytNsHc4nlWl
fZI+GJbtyxBqsiHs7NS0Bv/XAUcPtHEuuS2GZm6DABTcPSKBtRxPeZze/M+/4nJaYPNWNlaUesgi
J+Cgqg1vMX14/X2hh2jfkjJYZhq0M0PrgBRRq6PyadH0xZQnWm84kxTodcCxc2kLY1BkS5lMkZKo
xkaZhT4m9MiPBTM29SPmSHKCdNs4X4yfro5h0MHM7dQ+VJLhmGwGRcoa+unRpnxTeb2r8ZcKC0Wy
kWBG6noILLKbTSUnVTMXhS+S0FbWEUuS9i1MwqucYrbkAS0FnOfsdAptM0Cu+ccvKp0p/xQYCmq1
a+nkmN+M1oPvd/1otBVrtYuPorNYErF03hdB6Ns32dUeOddV9R7Yn6+XHGvVAYBhxbtxZ6MBNWh6
k+V3DQNK4iY69fnWxAuwguR/ign+N9Lqh3kloASx/71ql0vctg2RNZ6Bu2gJr38MG81ig+TnjK4u
zIUghj8q8BkA2xOpPPOzXRPdR1puzVdIJyk5SZVSUslSkaS7Lc7Ojhr8mu9rgiEa75oVfOmypgGP
DwlWlD4PmV2+TOh3xmz6O+JYZzN3m5h9irTUBuP9xAvChEzcqbS1lZppn8kD4PshNKuX/DJj6g1H
lTNEQI3mMXdFIbt0oglip3zkEaQaHlTaNtdYYp+LJpdxoOrdmVL0gh/exLJ06ivpZ3txxsJ91xRR
wHkIg69tGaxtX4o4VNd255vrU7J0J5ovQOYk7fSGhTtO9nQsnQyvfrzOyHb8V1pmoorhf9mPJ4S3
4rxWHdJq9aD78HhoCNehdgZ99ZV66VexDbxZStlPi0XNGi/ZCU8xwmhhQFabRYgmiA2nSDkfD86P
PDU/OWSjHlS8dqSsxlT4/fcFJcvtFw/Cr36GBN4B6nwX9QmcDLyVKHawpjfTfmDGJanGXCIDuAD6
toqzl1RJnKB4K+bBxuVYuQSx5DKd2pMPTo3qSMDuOhEWznDmP9n6duPwU4u/lRLhLFplPGgyYdU4
fFQ4cYaDesvAiz+3I16PIGkpgKb61YgrJcjDey8VMZDwGrAqHVCirKMN9hsm3qFUTRi/K3pOx5VF
lYblPodHpbxGNIQQKhScsKvuwsb61qY9vKJ/Qz+BWJRXnw+vwNPyvUyy9xxa3PV/ASe3WhGHlJw4
4umPu8gGQBpJugTSS70P0P9B5ijmeVAwz7D0ljTMC27q7z0UAMjKqASfFSXt27nc7TvWM2336E2t
SY8gDFuYXwhIHuJSZPGAnzapCpXSJL66If8+yLCELkZWglzEr9AQf6iZeGeA6fD7M5IQY+FbFtqI
rzgmkvGoG/DxBK0vj8D6hyNHRr9fZ1Ve0/E3DG5mvoR5bZmiiwKt7FG8hkXbJJ/t3uFcXTnzlTX0
rFbJwrCE8ml9nqqs2k2piCc6LEXhXBJTb3YEniSgNPMjwf2ARi1vOJlqrj0/5hHWuApk3Y4qjviE
LKPLZVarBpj5HUrY83LkNFKOjs/ugvtl6Fha+c63IbSjhaQwXZU7Ary10BGlSH8Qs5Skpgf9dbC+
QhQtICEhCpxbqakAN2EpXjeh7wTBNJ4hbSiDgRGo8z5PPUN/8n0H1TmMZH6aAQ9rYvS6SFlEqdxj
DPKmONBQEDUgoRECprLQrgNkZ4iBewSND6zbTidQ0bqqSpLNYl+LL+dpQwFsxi1xR69/iS4NoR2I
+Acun1WY15ABPQIdQ+M3iNoK5VNM/e0S2VgJAe+H30gzAwx1kYqtR/aWmgNyMq+0R2fG+HP4zXsZ
3wWfwiRzeQJG0ghR+jb8ZRvJyy1C9tnYajHQWwO3iXp1Sx2EiEOQzCwPwhlw51QkvFJesS8c3G/a
81hfOyC4kRFVgU5R69AXA5I8JVFELKHWkgPcAWHHl+YDsqw9XUjB+K/KXYGkKRj0ePEQK7wo4XGW
o/y2KNBJsrVrlUwpy+Ywas6cOKsxIwVx1bnKzKLA+PUbW7EGyH7PqOGMSxvZ6NP6bV5iSBXfkhbO
GQqjAkTHC5CVU904wFtVviKgApMr7ck5zhridojkVqr1rIn3/sQaSbTlyGRmwMZiKj5H0hCxvaIU
FezM6xBJscOcAxLG4e18fIX5qEUTdZ/YH42MkINbvjbn3apRErqgolvk2yznexahcr06OFABLQzI
q2apVbfDw5WU47WP1QdtdQg014H5kO5PwnHlVvaTnQki34A9AQlaup9qiU8FQHpBCv4Go3qLYBXs
eu53Mhj+BTAKcufy8+uYq5F15wlcx/lRl+DY5OMNiq+CBu4r5VddKIgeXnTdVBIF5yJWDXvxVs2L
ORmIpFbFtAz3QvQlIlxmxA+aczTLIZZobheU7Ab+wX8GBMux2Zu3Obm2gpK4ef7dZQZMvdedciyH
gZgLOqnSOgtg6hw2R8kHB+wbKS6dPtRtTSe8a/qNlMNxiq5tec7/x1P83drWPt5Ehd0vhJ7zQQ/M
D+R4LRmJbuuPIelw11ou4ExjR+HD+U6J/iJnW4rx1Bq5p5Kk8ntH6TqcUYFlplSfgFgkWHRNR+nB
ioP3UXJmrsYgF2roQ2+qMijLMk2oLkiTIa7mHdurnRM2ndezzBTFRErOUZpyFsJHaOCIxTWbQCHj
Q75R4yGix9bNMdPFmogy9pFewvXjU7ns7klEeiYSMxjrWXfY/zgn4nM+4RBXvdxyOOff+qDcJNCX
FEf/KRW427MUeo1FXvoWkxeGIdo9nzt5vJCnhDPJPKEA4x0XL43zoSUZEt9L1vlL8fEYIcxxipxY
jwPLQBvgaT3GgLwUcDzObB+BGOBk+q0I2oRSZ+HcEunLKFAECX8eaRq5zxN/h2WvlpUDjxbYM13c
MGpkWbIAYMg5AehvmoEVeSjOR9RHkI0jmqXgMW89OwQR+5E2NG0i2HwFauRHek6U15Ex8IDoToLk
kON882HxdIVgZuZ5tswXOgGEhlb7sk4YXMaERkcyvCGpAhLv/nS2IVgUkdbvsAzM0/uH7zOJztnS
979omd6NCh9MGc9+1SWmve6yiil64YQpA0nWFFEZ+Lm6502NL9d+x6Vk9TJzJXDRU5MJL+tnI00V
M14AdYaSB9KbxarczOop9yTg8AiGmfsnp8fgFgzS4vOkAbUrz2OBTYogXMdizNn6hGtY6CpvldMv
v+zyzXHYFE+r5PxJ4EnmJ6OG+jiXUL627ci+0WTTq3WsbrkR7tLM4KQt/7oqW7tEPgm5VzouUoSQ
qEPBN3+YvSIUiY6819hqcElvuRy2MiudJZyKMVIkhEJvd1zb2FA+IsIeBC+nXRa7nPPBAF2zW4s1
Lzh3vX+Wwvz95EDS27/UNohFUxiuXNCN0sd5aWsVlrIpREoW+OMsSh46kHqS2dJ+vsD7cQAuIxYj
ypVydxxHgGntI/Z6UK7y3ArDneygfMjFKXcmUQHwMhWdTjYH5XtBlXDXk+ohjTfZgP4hziJAKUu6
ebSUrE3HL3ZQsM91cPKv/QdwKQYuY83/uuhLsU66Gmut94l5N92qy2+B8lqx5Wg1fNpv6wQZFMAg
PmBRAWLfLz0aObCAmEunQjNmTyZQyrwax6Ls/UnXnSAvFIy+v7c5xhx0dFxOufzi03f4alNoT/Eo
eypiDWU3crxmvnsLdT2WznAR2uepJAjpxtFVZsllaWOpjnjfOeDTNdrrw9S+BopTxlpFt6NxkcJ7
gNX4ntYm7PPwbyFszNQu1Aq6YXj5iLv8xGezJuPiKIZprcvXgApJvhLGVEQPfBbT/EWDQMHibF2n
6EQjsejqZi4DvigB8Noso1gZ41Pvkmuj7FCQgvS3W9kqPBvp0n0mBW16sWOVp+fe1HgR6PCiS/M7
O8uUruf46mSLxLuXJNK+dJMaMs8B22cgilByxPd3vK0g6BkQ4r5pkB0NN8lg4R5kWSF9CAM9HzWA
IxFsx20lN3/e/K2oB7naRmd+H0UrHKBKPNrRqTMrN6UJn61fhwWUq1/VR000CHXnJVz6ine25tib
Itp7MyombtEIZ6NXtrESygHx5UfuKDqYBdWnpLe0jmxhHCOkg7HbH1n75FnQKpaXZTzuExRVgPNl
gSvgfcVEFM2p2ne+N06Y512fFGOT738PLWu7OA0GvGLxBy9SyvBB1tHcgw5MTTx00HWlZ0azd2Ax
UBffJbp/Wn2bKpzzs3BGSwtDrUlXW/NaK60f2aQmv0oyf1gJZ7vkSjCW/r8l7g2sKnbisCuwI3/I
wZPeg5GO0nA8L5pgL6mkqLXfaK6qa42v4jNw4qcnUhgFHBgioDxdvKZVoemvMc/mT2qGzP28m7Yq
QY0aUQpI9oa994ScgSpVeVAcE3hLY2Nm+NkieSDFpB4Q8bsNU6VClMrMZJ0rjlmMsL72lwQ4g5Pz
vhakPyIZuL/RkHMRdB1npG3xa9omBXgnvTKoiHj9dolkIN7UoXSLOiwHq1yh+06W3SC15GNS4qKp
TkPi2qonx7Xt8K4UAXDRj/yFnuO4ZZ1hp1nmFQ6kvfDKG4m36Lk8FEJFYFZRTPkcYkzLnMmYgk34
3xflplxwBym01hedxmErH+4Vd1+gf7bKgFIedtdz1bvz+h8GYE37b4kZ8TXBt9391ZT+Nm/WCZT3
HyA7PNewEqC67rSwIUOk5CZmD/a7SWLLOI8jwJBudUqvZ/qwbjtNZx4lCExv6c3GP0+MLUEpI6uz
OcBBYzqbaGLf80ZouExl3p3JISouA5iFKi9UvDxNDHclPi7Vtghn7Fjj7+hSTmIXGaV0MC0nUjxc
HGx+WtYE7stoX2xumwhaDncXMoCkP5+GQ1F1FLRnzJz1IWMAz6aeDztT7S5czJVnhPzOGLHMsxve
07CXFv6RdK2chYHcSXNFMKloCrpsw6uR0jHY5/fWbi89YPWsuKDLj2Pt7VQ0mcPX1+qe0kw60lY+
p+pPF1VWVvojKvkXZjxNJy/a9NcJTj+vo6CcCDwGdJh1+Rbsez+u0CmgdcOKXEbyE6wc1R9IOvkx
H3K1FEKbds79ybM5++ZCoPp9jUg9sAJlzobV2R+Vv/wgKfF7ral7I7tb5bFVpKTVwUrWBhH0tPmq
/t+aftlPF+QB5/bjGs5G42C5uRuxLxI2doOHqemvo1NVPIYIRXsVUd+vodcjZ6fcpuFEChFK2zLr
yASIe4ruXi/7KgXova6zb7DoQD6KlOUmyugOvKnGFWXc60jq+qbUsL2EfFH1sBoEBUnX09nMEUYE
7CPSH7eAn1SEdKmREjOehp1VtPhF05UMFeL/uhaZ5gRd3yyfN8sQyeDKJO2fdKaqc/t45WBpXY5z
KOQdQ96e7EhOpsdKdscHRRxqimDv/NxKEXc6y/QEoMZVcWA4MZTwK9XmcIN03sDgk8NYyb898G7f
Rujl5dWVGbyihWDN64/0GNv/9u4r/HIOrumpi8b0JY2rtaHXP3SufPuCO7QulNnT05el24wPt86o
RtUQie+CvTgPY2engNV76b3bRY9SMKaz0G4FMDxQn2biPBsJrDyH9pzgTLT5PuAJuyX9YuHYnPyJ
hd17pMDO/1AXfr6WJn35Wu6dT1PgNsXCkrgn+UFDTLkziso78mDYzqGDQ7h3Sehiv9OeeP+NtmXK
/Iqzeykt0AvMcPNQJekV+xTwKmu0477qMijoS1dNCxafrPd3jUwhyx1wLBlNc/kCR5+dotFa7oB8
Z2eZfMZQTTGoArtRAl++P07Ea+K9q1VF7snPxpgM4lHbNEgtcfL2NG4Nk9sco2wvwlxbMH8AESOh
RLuY3TFJTsmtoJGl94vvUy2aQ57LPGRTkJAxbOKZ8lmLT/pctFbR29SOBMzNVCm0yMWpMMkImHTw
2hzsMMuQTy2tcEWECgHM/IHcloPO2Iew7JLi0EnMf7e7OHgEgZY0AI4rY8QKPsV2axQPDrTnH1NA
zQiCLlGT3o7Elwd7r0K8eDnUPavAcrywmsUoPg/MeEq9gJsipITL1Mkr71eGFLu91zT+bRIn1pbV
+dPs4o9Km20oA7n0EofqgmyvoIUbOjWOdtdCfh7T8W4jQFR2t9QAaqdmMhyQoaVl8mJ9B9RUlWaw
Sa0AgN4sV/d1FjBVS8x5povwurGA5tgtrT0TnWSpxx7MB2RnVQcFkDm/Rj7LtGc6odahtZq1E+fk
R8cCHFMVZg2qjnxM/RCzvUSmng2PQAZjYUvC1Rw0qok/juG9vtz/pS1KL94Mks+Iby78+mco4b6I
j4swm78+5YScNfX56Qcso1M1gxud5aoDKObUOKNiYQ5PYbOP33Syg1xmB3I+zBUFxDqf+oqAfbUj
LByqhfqmgA2sqafSm3CRQqiFmVdWsROwBEllp9aVECSspbVH8wtbhiVheqRgZuZFSPup13sPI7Za
vmiLkF+pzcoVoBWJLmtKDsUo1MpV/TihodKA63HMe7smp1WPJjFmiVuPyzK1CHp0by88x9KjzF/d
tF39hnoZI71sxdz650SdtHuPsx43Lnk9MkmLJzd0S1Qh40V2Ne2N1uZaVZW/I+q4aWZBX9OSTwSG
SyTh3Gljt81Bh9pGUKDBmcYHgGBMK1WktbC/JcNQIbv2ylTjF7uC2Bqg55Uil7d3gDW97AzX6FsB
1uQ/xUQqIpjR03WFOnLmkNL8iVz+2Bjuufk3rEiF6HTq4EwKgmy4dW2pj7JB7n2HjLIkYT7m5Hr5
wrisPSHrqPX13hvLtk4snCdNC92Ke5cKbKaa8osZUUWbhUZU1BDitgxyiC948E3PzlsJXBpaSdOz
ZEllaYF0k0U72Q546vdif7/dqJiWgw3UA0NZxBpzJBFSwMFLUO2Z3wrvEohQ96utdDTjRvAdk50j
uO7MDpltlSyREeb5F0ZpX7teGzX0YPMiuu6eBso2nfWoD5IAvkk6tbOA876yU1RLAZ0jvcEMBVRd
2ASU/+w+KK7f2CihTo6/C9EZ734iik76ymlwiArxU1d6rZgxdyeZ9gDa10mn6BHzXaRQREdGZe9Z
fi846/YuY8NaLdygdEC/kRPsnqD1scGKYqW0XHv2Zx38MEn8AfJSD+/lVSSwidKBGQ7LTF+6Fr8q
gJGHHw7X8Fzw12ZTPARtrRgvchuv9CxDvZh4kzsalUBQE6ZbBvdAEEMjgdN4GHWBTx6/NTYLB0I5
vhvAsLojXUjEsFobJDqifH/wO3RJUg+yh2DMmVkx2cGIcw5SF8Y7r9Q64kH1w+H3d9r1uOwSTF+T
6A5RheHofB8/VcCu4krbC/fqkuZ4qYcNS7FZOYrLzbp+LfeKhai9whlDiD/nt/BDoMWYPnqGS95k
rI7HDj0G80cz61wqg8E13PresOxOpR+yhh4yCDxGdkInSyqGK7/NkOtIHQQZhmmyC7nl09M1fW6K
zIB6CsV03CryJu4Ezv2FS7ArOc74MkIsw2VxlvU18wi4YH9k1SO8HydKq2hfp/MGf0UFjsWBFczx
5MCTKrYdrUpaLrZxnkcjFx193m7fnh0jV9gud44yhTY4xBarSE16LqK8fizD67TqZBsPnd7jtus1
s9vHE2kO09i1DtTlfiEiHeM9uLBv5IC+9RbF3SZV/Q4OrCbW01VAlbN8ud/hjqDT5SZOZ1rx0JCq
ZBS511QwOCR8QcY6wwk7+JLuGW2Zt2mJodqyTtJMiKbkkaR9yOhIwCF1M7hqnWhy8LDYrx24vdj/
pD56UgeefkyOiY/xziN7cTtwTedRUOxEI4wSkSkbvLuHWrONa0irPIHgSo7kgWLuyBV6yuOfvc9I
eZwd1gaXcbcf7lNP2I+3Y//uB+1YjjrdqzQ0wEv8U3LkO4MGZUfKM9/0iIxVHBIG5ssVlyu4zoTc
bsFTkcomcqwM+INykbrGz80/xPfY9eJR8b9B2BeUL4RNBVuycleqac3yYY9FPYxe1hXWssSg+k5U
mqCIuZFGbiKEsS3APiVJFBdE5qbeTyAm/uWJN4sVM+hmzfdc64c7OpIaaJIrLwUNy/Y02tRHA9fj
uR0iZ0/r7MDy7LDzJvwkQwyKc2Rmlgnh2bva47OzmkaZqgSzlbMFHYVplC5kwuAg6Xh1NqifMr3B
hcNlVMSNyqR6YlOqF3LALSvJYaY257q1ihi6jUe36j6z7OmG30l/HcdQxMnsvGrfjwA0K9MhjX/8
fF9NxnRAnNKBXmC8DkiQne60TrMErzzUbu83Iy0mbqXB4qiOfMnklkAcLQeFSZYhPl+yQKcl+N2s
G/KJ4cm4jfOA4zYKVblyVr6++9f6sYyzp0OB1wowg9juUkqm4J1g9DhL6Dn7hyoHbVvrFJQCajpk
MH7gHi4fmIte+eeZgJUXKQh2bF2gzf5Co3LwLoYnNKKWSuWTmbLK6Zzzys2otyUL1nRy7b6YiA5C
r7VusRzXywsR2gvBTe3EqqwPMl9NathZrQs21jKrOn5OOCE94bLKVWI8Prji0HURdQTbcRn3lEwj
REX93MGJD5SKLGHBLtQd+2hOcrRufzIZB4TjGxKhuceoqtIhw3pG+6TOJ8snltwtx/993sWvWFnt
oj63Cy62QwCoWESQ7cW/EHPCDS+NEyI/uikloWm0PM5lK8xFYSXh/q2ccubDnQV2K5fD5PqFQcg+
TPM4DprMvTyfrlSFUp9MdxFRytnNghd6MQ4a7Ix0BeIRqS3JBQ2WDfvC1yf7YVWJTcAM2ai7hbeF
+GwkFkyUtnDKWXneDfYWKuZ5p8larU/M/LhwiQbdrn0EWnTbRT2lltLMcxJKvnhGY2clkwcL5ksJ
IvRtXw+ZPrY1qSFpDSHWYm8uaFJmbqG1n4Q1ymUuLVxEZlwVgglKtdVc+9ssBAUKfYvcSwrzEfP6
LwRM+8RzCZwY0D2WKTJbgKzUVX5szCD6tsbRrs2UKia601VTPaQwucW9Av4a6k0Eq896miwZt1mQ
ofM7dUe/2FmE1pGoBlSOztfyQ5CVEUVxY2KJbUPUTtoIqROuQ6qoqfUr9tjExLyK4QEJ/4PdDCI6
YI/5LFHHvS0TveZCcRRUc83tIIqWXdyPE2w3ChRLPGxz+dRJ3Rt7sSylbKDQRBQFbL5r+Ss35Mus
wTpe/9uDHWrY6PaAGTA+hlPtksjaoFoPjD+zozA4Fyok3aKiMr87HmX7eTWkxPTGMVkMoIyy31pU
LtR3Q3v06LFAU7FqpcmHDDp8G278mD5iXbbIII67HrogFGD59P9xxtv6GrWuENWgzRZKD220FY4f
h971HA+xdc22v/WkTTPXYDdsonkk6qlg1cMz9CEa0rvW3zLnshhFYt3O1dU0Dkg6yiW2gQCtM9qN
qiCju+pmE82Shz1ApqGRdXBU+ZSJETgqey01Ds1mYnR73xfekWIADBl1lm64hHk9wbA12JLN/MFX
rs6y9TirFtaUAO47uhQ4BCI2j/ONW9p4grFzRTGiT8EnvWyOL7Z2shayHu7UyomnG+2wNIVfxTzN
grc9PjLqEWWP1OpOX+/dhc/SKUhR1B8msDFpxEoRnyz8VT/7gi92NkupjB1txW23PyM/uDn+NlGX
fBJx8Tx/FHXjhRzzmqO+Z7wfBA9Q6jndkUmYmmsTJ3ApYnYak5BkhlVu8UzrDkTgbVOc0zkMA+e0
oF3UJhAEahV5y7b9BrMqInbPnxYqmkWZAe64c0QiGk6TjmvZ1Qn3Hvt7Rr2sb6ssYHgQXeVqsDwJ
iPn7LFCQUFnI+lracKs7lP6f6o157f2zITuCIxdO0KSNGt/C78/nGabQRhHNJfOzIKeq+Oucr0F4
vIeQ8Yxkwrm6PjlS05vvXdg8MdisQz56SkDWbER3uprtBAXuSoYojHWqghsMyw45nAcAbmSYn9zl
pPvKx4mEHe0jpakOixyDN0br8MyAGbbIzwwxdSwxdFlrqNUXHj3YdWrzTp/87AVIGrmUmSt0ntr8
a3RlxSH19Ho6s7kBU17bdAExU+6yXiAXSysH4MxeaZCpT15mcSGp0oIW5JCiAHnhz4UPL2BIErF1
5R6BAAAYkBfhhr8xMLqwb8hwV1H1yYhIpL28QuqGEVy5AiGtKUIAIfL7OmW7TNdHZ+APt5xlw0we
cPGRrV99qr7ZtGRDcoGIQ2iYy2qlMdlyG+1U1n2hU+nkMJfWXcvsLYhHHLb4mRvKinGbnBYRaKGD
bkSNm1D0085wV6fhJTrGvdTIh2j+H8cPGUflDPcgFzciFe9RebfIlOigF6sM2IniV5W4vXCjX+cy
LhziFTmHJE0eRVbcrEQSuc2FQcFq+2sN8KeeqAXcEFCV6qKZGr2tsQDOs4+W4Dv8/tdt28cXdr7P
rbklbt75rb7SQ5QBRQaPp9R4cbk67hbP3cy1KA/pfInnhLSTR1S1E842DsLJh2nkEMBZLUYBguGu
7TRHH4b6xgnTSKtc2VbyWoIR5Na6odfxU1Q9ZsoMAOwJyLR5X5uXxrk7597VL1PZWiXM8/VbTxXS
//Degt3GG64RP7MUON2JKrvoU749su7gU6Y7VmXLRh482RtCniUEr4hRcngv0hUD5Z6hrOTFLsZm
6j8Jb33Vw2yZ32KiWFSmZjdSFjOEMSumStc3QwCQhGXkVbrCYZF48XFT3E/DgTvv2+C0Jvf2Nd6m
qDYivhy/FkDDng0dFDgJlovCtD/x/ft7d+sjLTdZaB531RzFmWb68do9nDxLpjSUOV4taxW+JpTJ
0MfCgvgWkrzysCE3bB2r0hZ7OVVws9Fs7Ht2lVjQq32g8Yk2mIVE8vEiXt59L+miu6y5In02/u/h
e73HYpC42nsZB4MBuO5YVmoH7YQB48c4RQsVTPz+MS6CznYc+ceu3LNpOdFphmMEP/P0O70LVrFr
Y+FYP/awkijenssmU92mwJBzDa689G8MeDYsjq0TRBtsartllYqUim5N8F6bUZ0lr8ejiUe7h5Lv
8KHKy2slAdmchlP7V+xEnFO32q5C6dTg8UO8vUFslzzMNbyuTyjWQXJVyXXbh9xo9pKZTjoyEJev
SXEKXCSaxgFaJr49dc9q6CSULMwRdn2Mb5aw6rjOptLY4DV7vtH79bCluMnTU8s56oVu+jl+Y2g+
iS8afXXFd2oQfOjC6+/9sXtc7l253RsGDqNQV1gdBmKxlli7YN/OTIp0bDv9KG0r0CwqaZlxUmqz
RtFQAeXlPvkMS4nK9yv6XSbsBLZ+3PpJ+guSHZl7JDiJUTEV89gbJZ2nw9dl3Ivt8f5j4kSIK9pM
R4ZCCZVMqUEbgEhMs6Vh3xA61MvvzfEgMjLRIfGe3BjmSNa6Ln6jZs2iSbvPi9qQyHTNxCR4fdyo
6u0uSn/0f6m/7nw4Lk4UXsjz/XRs1/nbxVNNs6aSpT10JgeagXcwQsoipRcoPFok4VlQOrROiWyA
Iq3/poBZLQzHRlR9/1toMm10NozQAF+/2Cqht0kYbd00wwWh3YxdNgPuoDlDUxRO7qHNvmn+aGAE
00gTN6iywNpCbYJbQl/DNAwmhU6+OyVi+WPBY/Z+nLiPesUFpde8SrbZLMqIfJ3M0B6TwMN+aGyS
UOoR15eaLn8oyg8O6WsK2NQa7+UIDoYuwmx3bpUlIFRZXWMwcjKpT77XCc9yle9xKqLNRoC+JZIs
mMkQy6TMPTqsPCpp2lZR0/vxg/uKp6ES9HZxhh5H0ktVvaVM1Xwtk4E+MGJzcB7oJA6NIrg8iMwb
gY1ZpkjaTYPdaj8FqmnPMS2mQbQhi0oyU6QKg/vSA/eTxICIxwSjnp8YkS7LhNCBNDS8nUCa8hmc
bzObLN6hFoy3fpT4OWza6AbDpYqoryuAfK1HBfnQWeJORXXXear7qe8cEup9nDaKS4loUoDkGn14
28L7w/6oAEyX4XlzRnc4+SIvMwBCyICL7BG0D5KUIPTkLwvpIuzMlhmf8OE47YrXwxrbOQDR+KWc
9ELF5/9zEG3Wiz8AZfGJgJVCPGl69YQG0WAe0fZ48EUhr1/f8KSvo4d0vswsKWaDwjwjNoa9q5L9
M3fZRMJukp5RWQm4wKDMjfMNsBUS2UCfH5ZNCXC7zXaCkObtclcSSN1UbI/sJstdAOYmd+HHwUZ9
V0YwdBNrEEruYA9Sf8VIoL2WZ4EO0GkeJF8V5cGJCyCalx4//ZJgKRc2FUDlCRhASjRim3Pbncr9
j1IQO7O6DjN2NM18HZm8A1cqWnQRf5cFSR1zSHiMakZt1Rgbqk9zo5ouJLYP+Ad6jJx+1+889MyZ
RG57RLwHxxBJEuPNHz6XSaHgdGYleixXu0upC55y2n+EwZfdKCgse2k0mQnPSIU5/1AUA/XTzO0f
ZUIYuCt2DdyCB8Zwik5aKC3tsI9enLZZ/NRDZ/ibnQt9tBGM9D9SzAtMrdGT4prGywfb3GdIJprE
xUiaXVKucZrZCAflaByUn9Zli8EmA3eG/jzzolnt7hukDwTyO2aS3rFOrIeJrRRCRtQ1HvEf0AHs
GjbV3uqGOMzRu35WILCijIgojjNveiYfrosNSIBU1sau4FYVFdEIXpl/0zwKbmb+7777q7KlcskE
2KryA/Yopv+NnwLEH4GRN+eb3ryhOZH23sp9qbuzIXnAs6hG/ziYSxXzCWBqfb5lC/Tbc9ruhZtd
mxjZ2XVKmR4bWJFpaz+8JimWN8KuGzfyJykhaT68wrOJsBj2N+7CLQTuojbQIeb2L/EZCFPzPoka
0LMfxSVIxQMR/npUcb3RfbzRWAA6lss0eqXtYZBaQeNv6x3A5mxppMYSID2QqLm6y9hNufLlQkfu
SliHxPTJP904kyBt+uMVgFlX6J8gjuc+ZAyOCWMnt/UBLP8nkOH/Wt7gWv+t8GQclLEL3P16SrFt
LGg0WYYPVmTLPQJe7ELIBCFX/mNKMxR0l7FLWsu8Sb1zPla6pTAlsc5odg7Rk6WowNxdvX/xEVAR
mQqIwZgYCXTOuqUA6h4xdPFwXXr3as7vebrbk0WqKwjtRt5TjhcFqYrfLYekUyQCnSb/maqhhO+l
Ge4maDNdp5uuiiCblU0tzT0o3aJhKtu7pgCySAS761LUKurzlwpstTeAg9IR9JAufFw7UsopZ6y7
8OzZwwmCxegKpNrquFUF7iC9s8bmePuXlQD/PBuEEhrpfduP57VG+CAV85cCT7/U2/UJymT4ldoT
oPOWU4lzNzzUXPeW8Blfh6yeuAq2TiiFgpjdrkEXLpZKDDKZDQcONd9vkFEdtXU8gDJA2GyC1ZLw
kXO+4XrjXkIjotpSoTjYWaPJb7za5j1aExw1R7rk5G6nNQD1T8ANSnA4I/FiewxI1c8D+sHuWraU
40s/7reYLzOAbInfZ1DyG4qS3DCQZxcfkrTBjCUp2+ZkOiLeauyrLx4Jx+i3EEuJIn5Fr2NKhYCC
/yakS9ucaUOdtLM3pTNGbxMt2gVWuSOF2CLNnCQoSZDs9UDDYFqnXMff8g0E0/wJtfEHJgKgOE/G
64iKrLwXWK9QkmtVXWAuvMiurMJ3JEaitC6F68Zc6VCZr9AHZCLblhjMqmbEWcBqKJE55lDc4FF5
1sIfm0x/pWJIFJlA/zEGAac3JwsC/9X/eROS0t95bM7vqVnpJcXDInKzyPExCAFCeRswpa0Ojeao
a1O09ddMNkf/B0CYOPCzpHOTOxOmgygxurdoa7jW2qvvkCMOAvk173VPnIXMNyf+IY1wKXp0j+kC
XSM0176QcSkeJjTrKfDqwl8sxrNJ5uW0hwWRdKni83MrZqxFVbnYfJI6Yd3oBlMxEuLv6iHz8nK6
bp40iZdWEgDWu0v61gkh4OthNbY5kEaQCKZ/UNuxggWneD3wgeyNsNkpP89xn9v+eSVmOD92P2Bn
3bA03nH8QnI1vjW4bL/85TRnDFi4EL8Sv+XMWabDLKCJV21k9TjyN/r/9uxVKiGLc7kilPWwWnOo
grAYT0mUn+9HkqPSd4zbNlmjW4sJ9Ccc+MjQ7TyIyDBqCT/LAjCPG2iZrbyetJI5KsyQ12uWgnUP
baN+emS/LuOWXYkjt3yEJ5iJkv5LEBpGUVYt9Jdo4QFjJXOQilYxSRFBZiTXvXlXYcuNU6vTKErS
Eqr5jOIKtiv0KS3Qe0d6NJK2TnMd5kr3npXfT5oJK8yjWRrM69MXaJUyn2J3uRCIro5RAjlR9kT7
1owgCg1kYAKPjbGDwc/66Pe/WmkOMF568gzzHFazSjioJdNKqv7UPDjlHHSDh9ywJo9ozwARBxd9
VH449iSXQ3rEHV8PVJPnCwistUQnu0QhDPJ9czuxHHTnQeF3CkBi9sUMCdVi7cgOc1bzXX7sgbXJ
MpDBtb3WwuqmRNCe1fXXThJnVulCMumc0nYmO88qrG0nMKexrYMOJMIwuWmQKsGli8t/zinjso47
WOhvFPp41vpcGqKzv5LFMiMighP8CSex9napanNejfNRuV/setvnsU06GQ0Zd7qx/nA1yPaU8v6F
8rqSgoN8xv6JeHEJHN/fgxuS3NBZqCIuohVoFWbWYan3w5LTpVsj3yQJQaupBJp2R9BMJS19UIJ9
y1iyz/K/H0KOlf3JK6e00LDkq2ZN3XASQLtmsxwRlolnPr5Q5yCxlMHahm8Cn5OcgyQhaGnx5Nl4
+eyAdVy8X3qi5FMpfwgjLzQ8hvBdgDomrHsOgFbq4DEsiuChhGV3/FRGgT7Ee1EEV/mFjUk21Jkh
MSCNt0ZTLPfnvSwzg6LpfFLrjQqOaf9cPhRFKB1JEMLNVppU+AfT6pygZUkGFvs0KMi7L81sDpNR
pjDyr3x5zkgiZVRxnnUEBnW3z3uy8G/IidoPU0DHdFCM8uiEN40wFKcgbwKXkzBq6KwxqPd2gjT3
XXSGZ4N+boUYVrHCvq9egwj1mYpKpsTeJC52rYOiWVXZnY4f9JelV3Tg1bAEHkJ9KchGpWtpgWuD
LZXafb/BN5YPBhXHyZS8XbZnKk0HpuTwO0bxjEBGhCVF6ICYaWo1gam3SjJ2o4sr7Ko0n89aeKPL
x+MF392Q/2tAsBCF9KnZhFlvZ/GoqQoI2hy2yFkWkv4MJRGzJzRAoZjPVj4GYKp0OSDCCd2bRjpm
rdU68JHImmpItQ7wVignICs/pBlQnAogxRRRc/cWf8b1K0Ps9s855e1X6tG0Rjmd867hyVXrNbqT
4iXQ9/t9M3BMYtBLBiU61C30bkbnTRyNEYRNEQQ3tkVDneQs3n/UCAwIGO/eKROqKUNnUOzc5fOP
0j6KN4y+051mFT5h6y2AL8V3HzXjfPBxd7/kl562agVJ+KjzKmLFzCm4TmZSDd+H/wK2kMIarFzA
M+WKdSfI/HZG6zjcJKWGJCuzeHIXBrNbjr7IIPLk7JkPH+DaUZ2afqa5PwcxHT98D7W+Rr10Oitr
DOvF7mKeKUI/AIPUiPS+2Ijn07NnbjP4WMbwgmr8jpK2Qy7lhEb8Y8SSxVc4BgPtILPQ8xs2KzO/
f0vQA3JicnVOJET+c/9YKIlEA7uCGe0ne5gaw3iQs6RUki5CGEZEd8qVsxahbML0AOfS1R2iEVo4
MHIop2e3lEzgheKvAcwYSAVw+wNpS09rwPgdFPppCN9kcrNDjUpeHmX1vLtYkznb47wvhtzs5l7o
eCpbVgoZ/uDwVHFF7fIdB4Nrld5njDJ/8+lDNEV8fM5FrlTxdrpvLAGGCUim1jpJemtSAWEmSNMU
P9jhcm3VYxaLnz3nHYBtl8dt8zMBaPXakuhfKyrJLDT8kbyoLn13s8BRed6I67VrnjBEWBYvMYs4
B/wAimQovehe/wChUWQcyrdrBI3Z5l5MLwlFHgvm4As8EnR2EGoavJwYaLej/ENcCxhXzS5nHE/d
L+GDa7Ewh80BA7eGMUS2P2zYc7Xq641I4X1Us4AJN9eCdImfuhS3LN6K4F/ROxGoinSihtIQa88w
jqM/R58gI7rzd6kw82FxuEH3SL20xOq8K9C7/MplZ7ddMdtc18iMVmwymUsxtQsSL5Ml2pdKrbJy
Crd8emr1/0IlY3Yp5BNxtT1ma/E3zLWdj5yPxifdN+ECjKjEEw3J76WsZWWyOKkZhs9TE1I46QUw
TQprp+sf1kZZdgnP3L+X/1HKE2KCBrFuvpbE7SmKFW7ZgfBLf2BF8oyku06NYGwxfcKmBD6L6CpP
hJQGG4libiPZq//nXNx8knEcNn4F9f1s548IycCRWdtAmHAbQ2X8eBbsUUuSansuSZamv+OyRD71
ZJl3to3ZtYAQPCKdMGyi9d7oVFtARsAWHxvDddZf20TY9SQ+mO5ch9UaAIuHW2tuRUnyTSReSzyO
8uvv5j5CUAhmYdeB6htHRd+ndTRhOo7vzbGzUi/yrQF42+qg/cjq3NSL2yCCEATxHTWCoi37bOdf
JNPvmlJHVyI7img3K3bDThXUpwh/mRQSi7q5neM1KaGdC6Cf3hSx6BXyjoER1miONhFsaM2G9nsp
Ektqi1glD1Aesf+UDutSrnh+G1bnXJ9S4nSnSuICTCa9hRtP+TEnTYrY2ES/hyCU/TtxgYBiwLDB
Arpx+XQPiTrmcFHkycfiMKuSooj1pOiIb0UyZOf7a476I0pRwFVhAJGlOxBKuNvVZPtFeTB1SSYP
6lNtLvDGVAINpQlPCL+9n49p2LOPYVBNYqiNpWNbH4B/MYN/NhqAPSIq/f0dDe3cxA7SlFuEtaug
BFu7KNykJtADfAZODESXGLpArSJVv1IJk8mIF57ONu5oqMzZ+Zl+SqxQ8uV90kWVHuKQBz2of6sU
9R5xR35LvT4zaIN21ue7PFaHczYiraU+Mn99bGnEJ55HeB0Fr3y9ecKMKdRPT22Ygc3OBs7K3aU2
nYwc7v9q9B0/rDzR6XN8gOd9NGxfhLtm7F5b8DdwnoIMymnSFwszS01mhhi4Fq7s8oyvfbKbbBJb
E04nEB8IqnNy9ce91ukd47+tR4RjNG50H+aZpuo1hNjjaZM1lMtr3jHMQ5AyXgFPZS3ynNvuhoxw
0ZCxhsVMr44zenCZNVGC4TkWeFguPO5IimSjNugpIUaTCYyLm7qc8jqsOYJBoa6e0YVZCHv+giD7
Ea3V+E5fq7THBXbk933BRwFPLhbtzc8HoCflNXaEGX5iJatrVd4ck36GaUc9jQbcO2R6TVpCqImK
tNb34GwymJhCH3RkLk8KQFuSUT+kV44Os1/ABeRD9qVqKpnhSjnKvb3+jRxl3eav1cbq28oKPVTA
Ta9/F1gIqWJscXCEU2kGMHQUa1fhmg+uvAtZO4jKp7dMXU9jqkj/MS35N4849kWeSseurn6uCbgU
MMs+rSy0/ne0zwTGmFj2iBNpMM4K1pbAINTuNNFsanLrQg15RVMYBcdXq914thAz+cugt43cHyuj
vGL/qS4gNEU1k2v7Bydv8q8l9WlIIc5QwH/Fc7bPMwZD0chMsnSJUh6grDZsk8wlgRP0UqysdVcY
70HFAHan/QSJUQ+QXmeu/+ryiFxMsgvbEIwF/KZfpw4YPDVqYEmhznpDUEFDrE2AE1eatpfh519s
IWy02r22pPCczlOnVUDSdP9MnZ/+V7orsyWdCuNJ7QoqMIPYa5hczKwHOw/Ll89xdCnZ2nC6+Ddx
XebFyUwRqks5ii3zqy6/QYMSCzdo7Gy2tgFpNBDUhBIrTMWPdC7vSux9iiAujzgAzknanS59LtCU
Bwr0StZzQHxAvP+0CNqbz1Ra9i88qbU6yu55viKTxTajrW8uYzzAnE5DHdx6onx/09EUXfxGU3/n
untf87Wg8Ds5r9czGppH1ro3X//N1IBHrHgK35TYFayDf+7zz26Oje1TvK8leMTxJpIHUtcaoDOG
w6jQNJUq5AOrwA5DxcCLHrg248TlWJRB9keHgdhK7uLW4hEEaSHi7uwZ29qmi51eseZ002Ymm/18
+aT3Y9qsqKrQ0RF99F3KbjaUmFaIsollDLWnezuvI+5gkmBTE3vBx+xVmFlQ9s2OITIwoG9n09bs
PLDQnP24Sxw+bpGRl5Hq+B7PH9AESmybVbD/zwxJ/z6/FR8o7U5vqXwVNeIXy85EqV4gVugpCqrv
6IwBEK3f+hkXY8Q9g6wOyjReYKDJ3hEitU1PJI5l5uj9PHOYJ8zmuGxPqj9fO2h15weOeO5USTtI
0nzzVQywMXLVXNKw1whlLCBboDYN08UG0PnmcyF7YCAgeocEZzJIYeEfdK/YkrL4efWaaFGH6sd2
nHkXLRxjQFhj/Qx1g54tbzLXpLdMe6stuxZc3nIbKkXsje4WgzvdhGb4s7LSXt5FVgsBGt+P2j4P
54NrcIZCHC+tyqp9KUQM8p5iMewyPOqgSvVK1D3zPA5G3PjB57cMEts81XkG26urVNwQC5jsQ8xb
MzMsAvR/TXSH/dgSvZjB/aa1ItViV9XWXTmtSEv51LVscWerICc+yGuIuq2N0JZy4LZ8dU2oOhA8
C9WToGKixjGBG5aVMo/lsXkj3pdIXiAu1NmkMcxLr7NetsKvVtOIRqgo/Vb03OMmJaWFjk6ZiSFM
AeJsEU6+5xR9lIClg5kBCneWnvfTW0z8wboFeoPUBS5BSoSqdU0TZ8w3m12RGN0P46WEz1XxjdWf
EZ+ZyZI87Grk6V6ARcXfRnC25rTlCwOwptda5NKs5+jLdkKYptwoAyE7fFxpbowAYUF73A1NVjJT
OL0VZx5XNwYIwvFpI4OgQgWjpRHKqjyRlEyynIVVcFbgt2ElB82d1VXSyyM6k2aVcccybHzAowYx
KrtSeSDsim71lkjUSywZpecnXRuOWaqsnQnGt7oXamGXb7R6GX/DMAUVi1nNpFU136B7Lzo2wQcn
TjgCx0CUtkc6q+HGvfdvlnmIeCfFFJSy8yJZmDmixfdt9DsHZFpsMj9x5nHBipuvQ93t4C+nruyj
3jaUtEqx+HRS9Hgx3vr9UrH1vLLTARwPMlwjO91330nX+b/jTr8EE1CbZN1vETrsnv+W0hyWM0d6
PKkEJobHSodIo6qHSzVBvKElOu1A9J5kgJXMM84JRz8624dS+RtZnMCGyYWNngIx6Uo9NawFmJG2
592qokodL3JR+omf35nRieWw/jeshNx96OnWf0PBWfmidwwx9ejTRakk1kIMPB3vDgEr7jXxWu/v
VhgEV2Twdp13L9g/ElJZxdoS8r9LTTlcmQimy/736ML92n6sKOhS4wy+nCj9zPthaKXdi5PcIlyz
6aV+2zkPCg1cVehaXQciN38b5PU7ay6Teq//xSk0POgJzbjalQXSH4leM9Xy+kSTJvscxnYmvl5T
dorhZR8uG3ypRmpJD1Bby0dFg7DSsGDP8rz+Wni6uRMrOn2ry1jo340DPqmFbKxwTsw64msJdGqe
MGdIi/QtURska6FowQkCF/bf2L8NSolCDFvBGZAWPwu1F72pcSXvAPnxVs1IXTQuaFT8C79aj+c0
8J72NkRC3PLeS49t0vhW0arujBfDCH+NT6L6NInEwOe3v61TAUsvxxnq6RPZfDwRkYcRbqX509uJ
EyKDQdIc2Hyikj4pCkB4ypMAg7IjLxrhqYEHkYDOzJm7mFe2GlBmSuIi3Oaw6hfR0+enLbnEy2kP
3LYTGSKjLbvi+WkWMuPFVXkvWyLixolYseZq3engVEZubEfvmd1N72QIA6apE4pmDCsKJRZzoWZ5
yH+LzunSGBxznh+C7wmgVl1cBrxCKUZHD9ynpOpeTZd6/oYlFXeVQncIp5KKGu9cYPzVxvQ+eHvN
rQ4yqEtkBdcEPi0BZUJ77lHiMVuyc4nw8A0BG6o73EGT2X48K3GFXBMBK+PsDfGT/V3HjA3hA73i
/1HXidonlaNesdz2O2QT2jnDy+zybQE95hdguo2+bqL7ZOcRNEK9Tlqnogzpbd+iXD6wRSi9x+/P
tHefraSed9E15DnINQN0PAOd2TZZ/+4qiCLgcf87/x64ldlubZYovdAq45CAozc+9Oyumg4/Vtw1
dgQpM6TeXMH66MlUvLc/Llyhu7DsEudRAb+sjjEQZ1PvbeEPpIVa5AXtNGZD121y28ZwIlN8v58a
4299sdLIeInBIljyckcYj+FaGdCXEgSZKEt+JRMGxhD5OQSiVX8DyrTHtGjbSYK6KZFqHvvDr0Cn
WRnYLq6n57860pGYkkPKryf5wXFnlQZrNYxFi0B6wJx1SqW4qOZtzwTFxo2jKdQm9OqEmEwAH1O8
EBQXqBJzQU++4aKjmXSozk6zTjpEaBTtNcVujxSmJwEaL/L0mGMjXXjtVQ4qJtz5eGk3kbTSMF08
Eu+oBPANSlf7GFlJRy/dXlrDVrwfyiRVKLK7NGyljLVDrEpT6wUoKH0uombqbCHwivtjHj+lFOP2
icXbmN2W8vg2ohebaaEM6AKpZcAI/RdcgMEIrZr94cU4ybms6ZRjdHoba5+vKLqvDzNlJ9vVd+MQ
lnORirhpsvGaiXN/0mbFJ6iR5AJT70IMTHL0VWwuttw/llV7RDXiOp52CQzvoKe11Gqz+qTc4ZJJ
g5QaISM+PGqpkuR41WuLDT9YOeLyGmgkBIM3gEEUKfyjt17+p39KlND50GhpcwUyQQ8EgPDllp40
06hx63Dt6yVRmY7jmAfV5VMplsnBciH99cPB5WTPSKQhuEsd5TBRUUCaQ1EMLandug2Qa4QA7EM3
jjT1HTNwdep0alePkULlP6k4WQDGmquu6bpN4J6VSQlnkQO6wne05yXAh5WBRx2aYhW08T7x+GTq
XwbIFeZ8BwfOoNNYZkt6PzBhxQZY+DhVH0dUXKdkHgfzFmowNFJQRCMFLZ2hk70Fo17v75WtmPkm
qJE8/pq4RchcGAfEzapv9STA4Fx0EqHS6rvG/FmqJrODBqzsbtUKb384D2uX1HZPRBzW8GZ/hjvZ
4Ychru5DPyjTEXxlGlAJ2adfTn2HC2xArvdLF60ZDu27aGPNLffVmQuc+hSXZ2tCeKoILJPOLt9b
dJawDezT1lZwD6zyqBYT+B1nijDwqefh7zfILXwfE0wFYzskExIyykSK8ymlffAsi4mxt+lJ66R+
PjemSOkT6oioXbNwDYZp2CsoPWx3q2jE95WYa8r8nr5SRzlD6BSlVP3qz7eSVYRBMPmT8m+WF0Nw
XlOnaMbde8xjkdyk6Cu85MktUOjY1YqQYp5wwmtHQjuLSiAD5fXbbaz0tr+9t5TteRfiFp/JzBII
XjL0xpzbKpi9RNEtrRIY0WXmXU7Qv1iM5EWTZpPFynWin+RS/mMPyd724biI+QPd/0ZoboZqzrWN
VRnbx1Y/Ye4uo2GrE4htjTnKbmxkZD2cVWV14ZPj/eeK+R/I+ZKag+vGGTUnozQa1z/5YD2m2o9w
LBYOe7H9OFOrLYBEMdWnrp6+Li2ATExcxcDZypa+lLONyJGnjK/MveF00Bg22kzTttZbuOgIKQhm
i92FI6L6MJRR8ZEpTv/3aeBpBfchKIC/AwWv/SfhS/R04KjnIXSK94JxfOLcLvsgz5rENrjfGIx7
wfpo1QWuP46x8pwoh03y5EgAu1a8jOxWcjWSA5o4C+U26mJrOXxW6dXvgzssrki1HxEC/Av3nn+U
SLM69gjA9OP+dVk6JRMVr489mHR25UITiMOQzX2UTsgBYV7xxDyCVthgS6sif2S6elrxpLoLKZgG
ED2SHuNtu4VtJnf177N1w8F3gm2YAqsQLnmdh/swqX/bqsKhOvra02mVNooomQH3nV9SaUl2zDWf
kKzOlopbMC9NrXaiuyx0T9jpRHOiwL+drJHif4YMyMLEkFlfxn0lPPYitVpMxjhWOH/G+agS1rdw
EuDAaqTiZKil6kW+iyw/uIy4UqL63INtPIR4QtI3tzAbfmvKUdP+GIgZa6hoTJOlKGH1j0ISkHKU
CAjYCO+Fdt2qFgo4L7wf8eaiWJy9hTnjiwBCg9nxk4I43h04HJNL2chhNb+2+wFN+goPs8ahEA1s
5Gg565QFI4dGlsPBO8t+vGqU1TRA9a9jLQfckkekz6HRRAH2xsabLHrL/lIujr7vokvyaXn4cPdq
4ysP+enxrK3q22m4kKHg+LUXgcQymYT0ZctDxtGSUNADyUDlcvZmTpJdNYm+hhVm3l8Ov4Q4N7C+
lfv3/tsgcUNvn50nH/oz818v3XldqeKp2XSXIPaFlPj0QbbnuedRUFQWIHhsbqgJx56Bb+mBUDzq
7N7MIEitn2X4x09Vttw1152esaImIbk66R4KqoWZROb39XQIoCl2UPGP/Eq1O9+kVSRRCTLwnoxl
B9G76W2HphAoyEIXWGyBzPNA5FuOtojsJd7zP0e5VXkaK7VFkCPlmrg/ZS1d35LK0JtBO4XAnBT8
VKUi137uv4fOeWHHO9VXKnkCU8HnxRyZJVr3T69Y6krqWRsbIVzJL4wsxITxX/0KH46i7xh+EFrp
OKirAwhsWZNWHMZx4XcjTYOg1jDJukhWoX2t7TPHwrJrr5BGJM1e6dZ3cRD6C4YrpXC0DrMJYQWT
U5Nn2++mZyjHCqWl5O1J9bMX8SxSvH2VLpzPDOplf+mDSdBUdD7ImZNMum8S+h9GoLkr42gcb1q6
HuHJRqjew62jGeYBfuZCqRFMer3YH6GjEJiOaQr9mYEOMYOMU6mDkPRqPWyM9LbvUXhVHsaZnTmX
KtNJrQeVRcC2Eue+7tppPfpoihi3PvUFpgrSrN2cOTayPzWryJWn8C+amxAgkFZ6rg86GUbhtxmb
b/qP38vfuEhOv+t4+dfS+4NpvyNSkiz3yFWst9ZAwTEWVkJyR0al9HetLCL3JsiyRjrkkZMYLE4X
1qOC5MVeH7uV6iN6HH7otC8oIEbLh/6VB3UuLjgBGrUk4SO+IyTnKAn0FTr/Z9pAs+k2UF//lTIL
/a2Oohj5APba+S14KS1hGUj0a/4XMFwroieU4HVlRGCAqbbkQ+7z9Gp8GkzuvNHvmH5nybnUViHv
FXUYD1Q+Hn54whqREdZvBFSq9WTn59XEjUo+CJmj/BnegjBp42oixKApMNviJywvPPAcu4rjOgMe
5F2ji7uFI172EP1C8rcZ5vyoM+ZJQNvNavPiuPhZbH0j/oYXX+pwNbgr7yzsiWHu1T/SUzO/45t9
XW3RXc8QNA07Fe93TJGXbMEx8IX4/WhbwGgerO7b+9291r5JEDNLA8R4n1YiSiCZKharKXHFDsh8
ovNTazIcgQ2CJg7QLUSMGqMev39Odnd/b7ln96atYOfmb/aad4sX6pv6+VnOBVWaJuFaa95Ie2Hb
vlzXAPnPqky8T59MGGjeyOfx+g6LFE1ebZIjd4ldjtlH2E3WJpepgwlHBx/oVwIg6b5hTWrv9LqA
635aqoOE2WuaIzE5Bax8lvYCjjC3AftKo6qVJpbcuMgrpgAVXlLDrirFNBodCzaySLrWYSL8HuSt
fbux+Q/wajt/qmq5EEIzx74HON7IowHSMa6A1falfAQ4CrTrqLNVDiMvkkgPTeEi9GU+9elBJ3Kq
znnspFTViFE7ESmdF6sGQLqToFUH7YMG9sTl8OVDdKiEP1IXB5vma4RWfW17kyHTkxutvEVvFTak
PEqKBBzXgbabVy7qLluM4zGiaMaoQ5GU6ewohUefdxebXpUDMFyxQs4IBu1bm83PpUbW6c7RPzsC
zfQTuJHp0ZFnPDW/NJDHA89zEbmxCENYRNEkZw3CVsSj6ppZmqRD6rNOiyilDG2wXI9sDP80lIHG
Z9DKC2YWYAdKM0JU9FJLcyDyvHrYg+BaSDlC58QWjJaE8tRHg/jQYMbGgkZAyiHTSBJ4JbuLzC52
cnsE9yShw/x8Zz48GQt8DKuTGI3L8Ip6m4VGSn9Y8aiwEXdqrjyMw2awNSEUrmGCug496WqPFUCR
QymttfCbNtB/UT8zQ1AN958XJR/tX6Wg6sKFrNlSiSnUZ8+AMN56SLqgcGJboEUyKSb+fogy8bCe
i3aLEEi2u4Phbf+6/aT8kJUva2CyVesVgEBL+xdAesAmEQgnZAuxHU87zQbXHMnhzRSVw1GZQLlj
j0OHk2+Wpc6Kl6ko1C7yEMM9VKE9YB3KI9uSF5bmGhrQi5CLNw0CfaBT97QZDPCWWMe6nYTtI5W2
1gyDDE5Wny3YU3BgpsxRLbYbJgBkBPaPpyUuXO1lgcIm231FOlywGZ2hC5pqr2lZaHJiqntbpU7S
0eVUVwCbA47Ht48LIs3lSY4tV0da9yWD+p7WwEUKwK1RdVKKNDLlUPetdRz5kaLM0qCnnxKWhRJr
Vy84qys0xCBjMj92oyC4Stz/gMb1fedyPKTzBlfXQ8iqtL7L5HfqeaLK7QXGEkoObj2Jaxmyuj81
YsnI2jZk93FHNRF57yuUy1j6bfVPqA4OAlm/CS4qF5rS4wafNXgY7x7kTGRaZ/wiShZlaUgUppZy
KGDsaXB3O/zVL4XOiHFcSAoIg6ApIVmWgTkosKHYHwf0FNgvvJ8WL0Uv+p1ahK8ZVe2wFtgm3Kg2
EGEOzQl5QYqFB6rhqRAZ9XdbKY5RdxHssnyiMC/0tz6ORsQtzgp2cYiKTcLAGN1WF/3TWpskWkhT
ce2kbpklzBgzLGhF2U+Exgpb9GXOEZWB55fHMo5B8cGfTuXvecU83/4A8GbuCQJSmukCwO+jZ5X2
8lP4T9tJ+QQVRrY5YTESiQjt0Sl6NeM6ZJ3+Nr0ff0OPLx43cAZH4TkDooiF4mfOqQ0AX9i0W4wI
5+B2LpTORi0rZATbVu/t1Ow68CirrGggwDJ9hZ6sasxrHVqMb7zjXKuhzg212PmDWic2Msvfuhtf
8WN+UPnrAzYr/JXGtPs3Sgag6Yf+G1FHzY6blRqDDSP2Ivjv2rWRUcSlO/iOjfV5DNHGqpcxFFPe
o7Ee8sZ+6uet6FfTtGseTPFxMyDMmohGSaDvvL6PSg5xuY17SAord2bQU+tNs/+S1vjHKZHB+a7C
i/QsFg4ZTYKv5dCp0dVYIJmO2+kBSWUhZKUMhQBFYoP26RHjokEqX1OlMabJhbeSWmFYrE43Nc5o
a1O4njQs0rH6xTz+aG5GMpD2somFk0Jtkn8PJak0NlVBzw8crd6odivWZC1OwwZACaVVqSyM/vUJ
zm9WUr8c5e8nQJpH5OQW7Mx7NhtD07A+6tQTDIAEQGJkjFiraYw6gzMLNza09ChAiL+1OQFoh19N
xLBi3RW+Cvs6/j0pX8B1K3nm8DTLu/rndfyykcGU+JAGPEM0MbxVLq11Ml7UoJa53ZOg6Vm1FnrU
wlK9WwFrCRTcQ60iZ2ZmWKjjDKoaYG6bMT6sHaJb3uClPaJPn4ELqujWNvHP3aOZcFlGDYVx/U7r
967qHWGdo1e4NPHvuX6Agbx+MslXrnT9GC/txgaSMQg4nEXNfiH0moZC51cd+BSQtlucZhY4+MsG
GWCfnldJ9YybsTdgE0MdIbWozs0QHehpsMaAcigIt0vrkGfRhQw3Ya4kKyaT8HQ9zM955jvrmuU0
03y4m9naWOQmcEfDG5EZa0CNAKQxFK8eo8wvx0ZE5FCCoulE7pB/1wu+FlpZxF8vHjpZCWRU7ovN
MigVrEfs7LnaPaqGI5o2EVzqacyiXN5uk1abQqj4yP/vpJt7n0gTWdLHLfhgNt5oFLZ+gag4kI9B
gFkhPvbKSvzgITqSBFvyk9Y+bRGNHaCM3k1rf3mjdt37l1MGEqFq2aMIi6zNjONh/GgDRdQLtyCn
68P3xqQVm3FyZ8TwtQlibSisn7TrQjWR8AXgpMSZCBbqMIJPYgK6fx2bGUNsDpSA9asnuWc6beC4
2Gi4AJ7uVw5oDmez4wU0xmqSmrmY9JFtHi3BzlCLFn/j7wZOW9VVjfgu/8QGmMG649aCcc3EcdYF
cKNZ92HOEdui+WfikFBpuVAeftUWn3ry8LXMcD7xIHFPXMu7osyX1VbP9Zdr2JO5r6zQL94000Lv
OnokQfI5l/kD7IneR0HcPfqZ8w7s+cdM/Pc+mWcYEBqclyyVL5zIzV/xM2smhrmhdHVxjh/klOjQ
gwyvHXKNgJiQOwY9KS++XmHXl5qaCbcpRltBedoIaHZq6Vrhk69BANc4RkOrMKWnt2Ca0NuQWceH
5jidNOMGNCmGw3E2ToxgJDiYJFY0YC8Bu3RUXvCr0RCaeZMOXuVlpfpqesGJG/Gq1KzH/Vq8JAdC
WrBZV322XRz8j4xPkY5pQZGHibSDVuRq2JxOOn+41j3vtnQzDSbKI8tfNkudUzPkZN52PvoxtwkB
iPgeYySMHi/IVvAZI+49z9trbcsgjBFqEkbS3RVRhUlV4lyUQnOdOD1zlaRC1Nt/aWzIOleUpbjj
YRk3EjfnMjovSKl/YaMEKI9HVerRl6ZRBNZWBif8R7ysFWOsKYtovDJhpCVItYKC6EKgJhsvgFwe
pR0olxHDRBH7qgCpBHHeP7L0+wW26MF0gko2JjiZjRjhqfExqV/WHRBQBjROR6H+fVqS4fnQykmh
Yreo/jNQWV7QiwQr/YHigmhYPq3/BoDrRWKGpacqQIgE/Pu/HG+nhhpa840aq1AlaUnbXdRex+ww
DR6miKnM4ourUOl+Pkk7mQs9fBGsNYpOYjQiFiCo3IV+2ALjyWUZSOcEaZ2So4XExKyYQKC7SGJj
jep39dqB7O0/6bifeCR1LMDp0hz4B8ePJosO+45GLgJ/0kIbtfxvEU95wXx+oTKDnJkmv+LHrHSo
59DppyLcX1gR6tNAf01g5VSpjymLN3NvtnvowiE5aLExSV6vnRtsTidrMsVYolinQSxtpMwwCF34
GAau53gF8j4KqXnoaAWQOsd0MIfohHLVhfexfQbMixzcIisVYDMNrbVQ8NM2a/+7iojwaEcR6js1
yRsdHUxjtfuksqHr7fz/cXofaxhM09bWg4nSok9BYXB/rNLQNg1iBkiqSoSNXliEh1Lgbb3GoMEO
sU6lPouohovR72aGEF+tVY04T4GuE9EUc7pUbtY6N0N/VbG1HNvprt31Wyn56OdqB53jYHkJJBic
wWErYKNJKm17EX0XJfNAdgMl2T0qJ8MwKapavbq6Qx9xikrQjnOKQ/3dK4zQyDd1kkiA2psL3X8L
5Vp6Y2ebmdJBh7+tZiyPMXAV/Z5K0inFrNsM7sQnyzDDz7mXGsytzPGATxHppJRhnmdEcjvHhoRz
OPgHxCIOi6Z+gVtpV6d4DznLbAOivp3TGuItaIPaMqwOKD2WPZW1D/zo5w0KiBgfxj2cci/P0S2t
A7cTg0QljsO/z/vI7lWVhPthJqdVFQUe2p9ShmmHnTzx+GMdHzA0hAgXbdjjeTZCIizX+u6fGiKA
yOtCQW7eEPyLEhAf3wV4WoGdE2AMXcGIReaZ9RoxpuKkVnaNLmyf0ahAR21MHRT3b9OQ7nYy+Aa1
Be+kfDKchljvxpKHcIRTayxSursm8+Oa3hF4E2Shcm0dOvTxpUFwIxDFfoZYmPRZWdCBb7LDnDek
aB0BiUW6oWJ9mGbl1/rPr9DWYRRCZMnZcyOtEx0lAsZ7PLvG6VlmYFuCb04CZZINzlcAOKfMc9J9
1ve5r7kUBJR73B82Dfq8tbBVYwCzdF1VKjZprUzQVUPtW8t7vaPz9LQu9Vgm8xNVRxfqBcwyN6sT
aZeBPjSr6KnRTOju9qkwzzdmLFjrk49clgoxYYFQE1J0Jor939pV7GJw8pHSU7PX8AKufnKIUHJh
GSpGQD3kJwh50twhG8tGnUe67oNwg38CXdG8HorE5hv3dDEkt99vrHMeeyQDcX0BYdFjTCzUnbhC
2B8IPfTlbCkEBX1mt2064PbLC9KThYtQgIUmRJz4U+xe05nVpSySDVGmd+0Hf/KG/K6VOkTzC3td
IKIRGHuvZAxOWGsZ6Z5gn0h+S5KNSYjNIY4SdGfd6vR9lF2ezQNCH+dfEudlF4Gmb9GVLx2F+/aW
fCZzI7gmMD1yKKJR4lcmyyQb2ce7W6EcZGyjNAQoi4S2TmQPYjSOHXiaD/TZRjqWA6wlu+DL9Ux5
UXDCXFNR+YjnOBXVNWC+Jbhr5aKJ0Rbc/dAlS7pSAUtpJ3hBTL1Pm47+9HqL08gem+s7MHkT5YTt
mVkhNrSwuEuE5rxfpcnpt5ZC4db5X5xjCQSYYGEOjsYLwPWkYGMwRVPPFdxinuLHapvgA8YP4TuZ
tg2htzEAnd5dLB/g8Sq8/4v7p6wDt1HowGzZuDHdWiDbodvnpctuB4xsXt4ziuybJ25+jdb389rF
w8FhwHpKWhCUgMuGZI2KalpY7QkT0GkeNQLT9jv4Mmk3wVyUWxso89dBfYaZ9KC2Vg6dtzuDG4RV
AGp1nuyVkvt77RLg7L1cv2LCEF4uLGa+xz7MRqV6QcefjF+KFrVUqQRZLtT3/n0LvrI1SVHEP4gP
74ZYruKLGmmjDdg82aONd0ThzAXFYRbYKUu2Dpr0mQn9pIn6Efp7oSh2WQSWResElvPyYoaIzQXh
MTds6Y51D+I1yo0Z2O0DnIIqMRzQYw0twXGi/mAdo6uoPYHAuh7gU86lU12cWtfkA9iL2gCR6Mkv
v4K/ovQQWoP5St8DvxYg/osgCd5gOkeVckyTytYt+hxw/IcrZX8ukGLzzEcIaXcK0Y7abbUb2BqH
tUmWnTXdEy5wYpycxqS1ycUES7kmyufBTqw5USzJxCmqcgdI8GBMeq4j7wO3qb2JlOjARojpVnCr
g/3oq4zvZL4AmT1vHintkJu9wvRg6KZ94Ihv/G/oyGIiACDIYXCFdeb2UF5vrM5OV5EmdO7qNujx
iAaKVLB5ZuzTgnzMWufqD+JGeGDhFA9BVIJr72jWxCVwzvX3KOXSzu+7qpKMjkRyZq7Cn2mUQy9f
eiQN2rM5daVoN01FYenUtz2WAnfd2/9Hb4nkMsrFRcx7CyXm16zu6LsWTO7lz0LSfPrT4d2rWOBy
njPbVejaz9cuo3UNVMovF8gPzWkcasWaoetcmoICgoKHz4qo3w3mR6nCiBuDMCHyJmTFr6FPGAKv
9764MjrDhTPoIKZ/dmDdgNL+LMAtFYHC0ME64MXwzkdwUz6eINNDZ4lerZFPDbpmYnQgWQfFpJKc
6BWpFd0MCp4PFa/H4BeAl709YmKgaTVelOmTgb/sWJQKnbRgPKN9s+ZQvwE3JaVKupVscX7rkGkk
fEBERgjXtEDWaEws11M6f4nuQ2L0k9GpQMgOiVknDiz7bXGat6OGtbLRxxCzQMVV0AzKZGUNk55U
ic/tyY8QNb5Ck460XYUFUyf6Jal4FzGYt/sO033DSvFb11m1AJzVbgA17k/1BpXMACgrpBY/FH+1
KQ9UOYUbJZeNPPWd59cdrv5MZVUO+MWM7aJk5eoKWzHcbZ88TOaqtmG2Ho/MH0YMO9mWg9LPv8RY
VZ/Y+xH4JMvqEfpoPqB7ijlA/W0jt86oBvnXYSddQHwxquTlqHSBtANdyCHDMgalrhVVW+jKa/i6
Fx+QTLZzCsqsSFgS/FlhX4hY2rNH2kEh7to1o4qGTkIUyPjySHCy3yw/1knF5QkImZKQWj1X3i3e
qs3y9OacBuds3bW1Ai/hocI05KcROguXklEcbCHr2Hd+t8mOEyiZnK4lSSZtYlFu23ctvp9jO5oF
Dj2GQqt5yiDyM8+DL53pgoJ4ghDkbyYGnDYs7mM83U3qbMFWL96zDUf1kfYXFaFy6lYnvygUlVFJ
aenSBvK5jBZMNwlnoxiO/BzFAAAgxP5uWWjCAW1PdvlmTzJLMS7EOt7+mZVRTliNa5mlrbrDoC61
nlauktIYtyZnHUI9mq+t0ilqb5DvoD+n1rkHCTLcudGRGy0K7biKef2ZwGgJ+f276chmDraCowSB
yyxA3zMmLCTudKh2iSYu2XAFAI31cltSKJOwiDLjQ2koXzfqbeKAAAbKBALqPM2T32fcFV8UyGWN
4tdXhrG+fq7R/8a3VoNHrN0xedEPB13bqZj7CF8elsKEHrlesXoOLEv0M/hmeqNCqRQCLdXWtZqf
jIzKKqFrO3Xm/7GI+czEJRumpZy46j56vLtfJXondotdP8n8SQnEuVn8OslrrHtkenhG8269tDs/
/8/kGfhaeLofvzu2epfq74YDDJJCiViAHSHqPonABcOmUcaSvi9Np4LozhgpAGo3vlKVS1bYI+iY
H6sMFTAnHQKNsLSGGWB0dNht7RlPNefw/sb6mfWnQ8TmbK8QarHjsZKglxO0ZRA6xeXhla0MyZTk
hbbi2FE3k+WhOBVtmh0JKCU2HH623v6rdGNHYNSC3NIAlBngx1N6lRkqpAFb93sx8KK+5Jhw8HPa
aP1+ufAYb+9A7W5iVeQ24KOt4T8kXKYqyBQ97fEbpqHTlDRKUID53ygtCRbF5PAYMXCOSYD2LJDj
lxfWHRUzq9ZbXQQxp6u4qy/9IFa67Ha4RwKDfAP06phlH1Nk2CdZKPjiSs0mvXrGVIDXFaB9RqZu
rs53kgnUVYE0Fkmo6VUsXvlI9zdl6ncaRu7UvCT82SMJaBW0Rak62beLwGoOo1itZNsF+U+zao3k
edUegP/7+5m5rmgHdqg04KF3fcFSfJZoSDg8L6DDdtX2cRHz56g8nPFwlkQma87kOfZfkCDQ2+xi
ddHfuxMxFIIFwg6uO7LOXUnnIWr0Fog6cendzSZMQ4O0kVj+RzqI0YY/mnmF8jNAdhPAdKcR8zhD
8XYeL3pCrnbLXsz3an4O8/gDFl+7KcE4SBJTx54uq5ZFA5BvDOA5mY9iJlWpl4ScEX2IFT07vCPd
stu8YX1EcULNJW6W8DF0dvyjm83oHRNtbf21THkKBfjQTYCdpzDoXZrEhpU58V4QCJWfyARJ2oeH
tCq5l103YhMfwu3l1tBmh+9RrdQGhhU2EZSplfxrL0ZUXSNFAotqJo3cSbURDhL/H9n4T2SVPBB+
qpA625tIHD+Fm/XNfCRNunBCU4qlo2AzblQfyBFscFUXwetDAtkMngJ7DdGdYK0PCrZoQMYcudHr
sENRkJOgSUiQIhsHT7TPSd0LpIwA1sUOx1+ntjPvM2rEO8NrY8wVXNLEwkXnRZEco13qMIqJXNBN
E8p26EjD9HUxzqn/i3p5AGhf86ciW7hsFh0MXLvLOdr4SvA8IiEQsu0HnioQ/jURYkSE5Y0HNT3j
MvNpqXsx8H5u7kqwkKqfMmpXwEeYJfuezZr1pZrEuDczXxrh+foEBhTzzcbwFQJQn0l5s5F1aNAv
BAQk4YVZSoAqiwdpA7vvrzQyDlLUvtAg9ulY52IzzARz/t/sd7cXlGmmYXNgINHWMo/WngeedeB9
7F1f5i2nOoqwoiDQPOu3ndWJMdktgbyakKc37AxW4+ezZZZOoRggrDCqqAcynhXXGy8amw03nXcu
f3lOaZWy1WQOZzMOZIMyud/ilCY2zWeOxAURoUqa+ufAvUKbgF+6jgv8/TFuCZhm5DNVlU/TraKB
6IioiKgEu8tFhBkZaOLN5t1n43LX0ABUz3oyYvnrfD1UI5ED2MthuZnYnb1HaQvW37iljPl3Je+r
qA94a3q7wCDvKQlNMaLVpLOsELr0rF5nNZp0lGb5kbbq/3gPqcde4LrAXklwBpHyQAWRgd5RyRKr
u3yQmJx0bviX3LJ8UZlGOHVAm15NPZLiXmf2o5N8m3+GzBvgbiluPCvW9gWPYErOut+Kwe7XNf+l
MX+norbc71zH7KLij829sw49Vk9qPY3NvVc2bPODWfKgOvjVuuNYk5NWUdSgvtM5G7zka2HHmAmJ
rwJMTlJp3GKxsGpI9V5Lw1ijw8pSZtZgvPjvSRPv1+yNQ+ZsxI6EoI28K7OArTzzMYd30BoCIwCe
vfTk723GJHNZkKDQdKrekcLDEIkvgHWCq8jPLamzyLzQ2Cs2jRf94+qhT+5OInsGLLUHiltiFpEO
+W6W71os3yQDMDWpWG5yxT5cllfe2lCsxe0ms81iLsyYxy18cTB9j/68jvu9poL8b1gwcEY213QK
vu1w6v0DQhN1egCHS4jS3FxIWBVjsHypgzPvBrI4GL21jQ1g7IE+QHv7+LdHaLAF8AJjVCCZiVj9
4gpdMRKg+B04v+2E1sES3KhN4IW+ExthDhI35LacRJHZByhMETd0mh7xYU79JJWCkCWF0wBgZDDp
VitkqHv642vezzuc7TVtIhYQRgX2/YXySWWLv9sXLaO1Y9+S5huEUa+CfxAxk5NKkjWu31FppxQb
2Y7E4biWeSDJ5LReMmZKqSq93Yl9beIzxJz+kjn6ARe+tlww5ZiKe/Bc0fDsT+xj7knWU6kGz0tj
yQ6HbfmMDFKEaXX7j8uJea1YMjMThe9ZyBNDRd0OFefwJJVLmeC2RmeaHJ45/RyD25jEKjZUzfmK
AGKahbnunRAqDeYHzAYsbhq6S6zvvzH41WmPIH5RgkpX2Nox+flMXyWgYVs7qNBbVug5nEuiJKrN
J/zCsjHrOrXuQiWOS+tD/azdG0nm+t+COriFP0Wl6C9sb11n283+L6FTyyFt2fmIJeLNIGqlwnaQ
GgcqAC/CNAu7r4bDxEDGZ8cHqX9uxVC49T3P0Z47xXL064OOT+TqpVfRVfrll2dccV8Qrfs10Pao
4wnGtbS4vYh6CBW3kl6PkzS0ThXS4HbT9pl6zcnEzHQLsyy+wbZIcyx4pdphoFDn0m0cjqZmVi/n
FfKrH+Em/4j6uY8a0oHBYetTIQKfW4ezDvwXfPlbii3Morw4vyh4sbnIXX04xrwo7DLEyXfTMgIW
SomCPFTRhslb1TjrDFG3CDi00SwmFWMLT+CYfvMZ4op7n9ub3FXPnLO1ncIBJaVWqqMLPQu99cGL
EyyUsVavhewIgbQAatXpvAv8XobHRyMN6O/6pDwQ0Az2i3k0k+RjF9kyMtq/Sur0moWx8mxLpHgH
d7/kDavLHAPvYqZCsy8brZnlRAoJZohSS4LsaF+KTVjq+86kNgA+6nUs6AcCnIPDX11oWXBa0VAA
SodAj5j/smyosSGuegPXCI2rVP6C+QD+twlx4Z9G5XI4hBIjNBZtx55ETMhyXzI/AGtS81mE2oi/
fUawq0tk7y4VqC63wTeX/C4YW3gEjItxG3QtiIB60+TL/+z6eR5nQQHsrwS4Z4hdsZm961tLM8y/
j7ovE7GhRgJL8SKAIo5dec2/cfWnrPpqnFmjAS1HdTfrMkRU01AlVY13ZWjjk67Ii3alaDjH0lhH
sWlAKLOCf41Vx4+jTQQj3DB61/2vC32OoG3CZ9Cf3Fvn+YH7OJ/zjjs7oqZ7jGrvaxbJxIojWINe
QGBM1yTsdvQwhH4NuNXJZkHuMXHjUa3pnlBVU+MZU1j2MiEQp1i5ujJbMqApCuDkUaVLhcgvTriX
0JBrG3YGv5AJMDFOI+chzfYYTlP1zSkC7J4pXtUW0JoaEBAlPQGj3Fhgo62NK9ppieQeuLyrEu1Q
BDMvY1/7nrrmXAngZFyE9UMn6+xabDR4nzkFXHmvOIYMat3k77+nUJUCLrPO0xtI0mWd3oPulr7n
nIezj0ubpNMQhyQtOkKDa4NfGZ9XzQUvoCLgRDO9LzeoZh27QaqThWzNiPMmSLi6jWPPxeScbN2G
hlsG9ZOgwY/IRmiPKGHYcbnTyLLYrhcudZca8vaJ6R/vfbmMIWALBd7w0Lzzn7lpR0uWwFJ9Srkf
13RX1BBpkd+3C+AAkMjDO+l0AmuSN6cZRjhXam24pIrKRV65tnVhSlDAJ5Vmowdb9oDA27DuQVGW
r8x/B7WvoZvpKjo1S9kAQ9bRyUpwj5FlpQg1w8gGbnEvjsYKyJECNRanfSa6onSaE9PssaJHDVcy
q39tqElAlUdQ/zP0IBG5KduqLYpMf82kQplpis9RQLJoO0fm1o9lu6tUPJwqlnhPQG40n3pAAOVO
U+I7EYzUUky6Dj73S9v9IfuhXR4qgwJBteLjQ3mr/h/AMN8iVw33O6ATwyQQvBH9FQ6tlwRkCG6o
xF/s6c7usBYHNJEn0D5TEc4zeI6G5e/urQhm2OoyofVt5E9QjsJlx+o3JGuaNui3IMBosk0rdAIE
7/K42q5AZTvu1En6dA5Pbcb2EyVRtnPjgBuAIyrqippmc1c4rwIhxoRaBB0wPCFu2XSD47DdoEQM
hccr2hKQn0WT1rsG4BeBfZ2+xNtxTGXmrohqpKNN3NvDxbdrPrmyQXrWXgpmeZXSCF6ODqBgp29E
A3glGE6RaebbLkJyyY51A/Rkz3NL3uBu7l0hG1E6HblGNvVkPkWl/iD/2VrjsVdXyR4YdKSahje1
ZdnIb4MDI8OKGzKMGcfb1vNazGbzuf83QsiPmk+6hRVsWNgdgwhlilkE1o06sst7NWksa37jecgQ
iBN6+EQEVattfdz01P6sRe6/N3V6uylA8aMAyMukZT9x6CRt1Nhi/KWrDHXYM/pEgpsA0z6ALtG2
59ao4U2yZxVb0kfALyPocxHNcSqpTBp6GKu+Hf/dPzqXcq9/LnSOCzeEk8SSI6ifZ5IXzo8O/TnE
Ds+EnkftaTwMd6n/1UyzN2uzuF1Tr5nq2/NcXUyyUhEFuKDYetk1/a8Jq5P0XYXyDcPFaLx2UqCt
1C77iKrotW8Nqhp+3Vu2CsK4eqvK3yvAsy6x8f5/MRat5zV5DWm8viEUVndRE3ZMK8RJwWPNqvtf
wOIGmuWvgGxfYLz9ADQr/V7ZzsjkmGhO3wUUDnjrkdFs8RxqweHgC2UPV3MP+37NlaHA02M9Na7H
TVcks+Jo7pq7H8b30XZIhkVNQ8hPas1gb1vcPKgL7YWX+jmf2DDmLhcn3a4KAFpmIBAj56abnjaW
HFD9OyfPVGMRHwFF2YzjTbdg0txWAdvcK9bLiXs/QaJFB7T0pmXCDaUzutUzUhYWNRqxt20f5W3i
sFsivnh+THrz9D6Fptep1kiG7lFlnTftazX65pQA82mJ2upcoqOMNAOKfaA+15RuGUnDbl++hjPD
84Z85n/KyTFCN8FutZPXVQyFF2ll0t+ctEkd55dWtP7R6ERvIptpLKmw4MEt5iwJqLafPc6cevas
K04UrBylyyDASzNTldHPtcEXp7XO8RDfH9hpkJcOrtE9bd/8j2b6n5bOnXa6saYlSe2CzhZF0gtq
cAl8u8ZYPVVUcg2yJz/yTJRud1HF8ZQ/LWMELnLLnUGrCyhBMl4mGTZD9VdDXQV+Vh6Np16hYumN
KiwwBVulm6e07heIEhOHtWxXzdakSZKCOyKceP7KVY9u3E8RTqgg4WdsgOFDt55uzdQ5Hx2zsP/5
rSb2IXcNVAP9Qpg5fT5YcMbU3xJjQNclGxzx2FmbVgnMIfwX7accO2ZDmU9sNJ09TtGOsG0bkki6
r02KoFoOlNnzuFngVbNdUQ/hAVAnV+YAjm13AXkBfLlgGwkQFU/SbtkgChluMYGjjSubVpvSYemW
eI0yh44hL7sJePiz3l0COFNOQmfJCM+s6wcPpNUUpf163Ph+6GkSZHGzS3RPiK/oTQaFn88EMoZ9
gHbV0d57g8X8iwi8XiNI5qqBwN5mRwhcxIj/dSZh0c4wLboDwYcd7Gb3ROqJ0vV3kTHxwDuY7sSP
/4NoJqjRVX8tRDgOdlBpTBwl3wAxPzkSOrwQPhM8BM9MVX1dCIjll0Kd5kJsg3dyhK5zLYNqViIV
2fX7L4yJ+KN+pZxPPTSV7oGQBLQFBXb0ZrebL2zID8Xa7qD+Rk9FmJxwUdkcPU132OafhEntBo41
tWJPPmwPs/LqB6NodSqx0RUVZvOiclLZGTHxzreh4nmk2VEY51T1hldBmX3hL7trND6PTx9SsDVG
NjAlRCQdBuQdtu/xKTu48gPqkctzasynDvSmJWqDa4T+QaoDa2itmPZ2wcgHprIMg6vo6pwRdBEV
WflXqMDjOKqiYJLk/QxKo3WMM9mUBNbkIZqta+XqVE/LTXw276Ycjo6g6Snjuc1cxgdOU+qSk/5R
Z+G/2wP3Cr2W/AYC2RGGJxRTTO1iHOVkfeCAf5Rvg4YzO4wsoEuXBE5LDhTIvUjHXoEFAMiNGIVl
BZZA+F42T18Jw5AFH+G1ShfNuMeQO8X8lWGKYJd1vr6tMYqMG9SFlr2G0NwrPdUBHam8Ymz8vZj6
PoM9xVggo3E3Uvrdv99W6oPBFwUG+k2LBfSfXQf/OZyXDbvN0RDHHIxW+3j9HI2Bh3YuWxkH3kkl
4wmx3di8gL44xv6zURcN9Bta6iIt1NIcSXMjYmaIOGJpjVyNoErkSA8tCht43kIeoyYUuGECgAR2
TsawYAzyMyN+wTnT9D+y6jWWAcfSOIXzfw3fYSNLYfEu0u7MtnprKS8n1a8UShfM7O/ZBxOaNtkb
VIHSrDlg7G6UAZjTu1wA3AHIhwNa30elOFBzfW37ooscBEYQW4RVbgtRLwuXZsypMKx0AdWi6ZM2
UHKxsN2ci6QExg6Z68DZpPdYMd5U1G6AeilD67q4SH5lUpKcnZQ7RGfCFWzGZ7PY7IXXkodGTgEb
wPIf51hrQzRVsV7g+b4ixJ1wiGlGyZAM+GR6Cdeg/qyumn76B5uDAIR+I9pzapFNP49XQ1UIR5fh
JuKoB2UiG0X90f4N0jPP2+aSmuRpFDqfdgKEfgwc9GeJSzVVpKnNirsxxAls84/SDj6U6lLIfQOJ
kKRPP3/gJK+Y2hPGS2TCY9vD9JAzYUmph2BCwjODT9xqleowlNir8iRqLEZYIxBuSfdIQCjqz/7T
5ccr4e7Ej8C5hu5WvCcyqVp7XxLBQdXA2sZUXt9jrYQWNkHvPXKOwqf0Ou7LgZ5Gw/2Am9Vv0Tmk
goQNTJKa+SfX0AM8e6ggYGjyFJ4TpGZlG4djl/km4LoLxCcixdM0yLP7XJHmT2M5YuZeXpZeKD2N
77STRt1+Tcyd8aTjo1lEFBuqV9piOZ8q0cMEdNYbsBg6s8PUuRAoqXWu3uHIeNUD8UD6uMgPRSHD
nF5+dO+iHIH1rnClRFzugbTuv2ydA9P2Ga5fbROKajzb9FOPUsF54+yTRcd5N/g9rjUaMZXj1xko
T6HbksaOgaC3O4jlMmypN40gUQyPkABrvPVQWy656pxwtp2LtDb4NSoXHjFD8vUT+PDETfuBNl6D
gRid1KTc0QHJ3oF6zbZmyKL25IZTvHbV/DjaJDABfHLpmUTWoQk5TGrTTfNZeeAWzKUf6duUx12H
qAVPYyzojYFS1AgCRyNbHsgb4eG3Mb0D2iO8ZKlpNuSa34Zn0O3RLTvamWwJi1xSn3MoKLGwJM7q
J/RN9CUeRCJWBKmTxMCgFxU1nrgrNZwZAdXrmNe62E9CaaIwuK03mBC/lIzKa86s0MsuteylycCl
z+IB/Xba2ZuTLCIz0y8/VW1cad/CHygq/crNRa7UGNLfMnYh0bywBvZ4tVGtMhQjxPOsun9/mYfF
Jla3P+mrMBCnNud1k1ESuZSW3ug3AlyN7pkqv8casaLJ3UFIETCVNiwMDUmD0dU30RraLcvLLmEn
xWy5qOOFYM8/aqofIdZvwBQ5ofEHAxAI9CdI8DE3OLDtPcCEwdc7fT3Ium8K6ZJiTKGlVf+BdVVj
FnfsSIHb3r+i/m2sDTBinZiopXTahVC7UZyLk5xk+rqhg77MsYaLKe0jzkKP5iWz38FlhCuURqcN
n22wwXC5Pgl1pA1vO65QTJXUuzhk77OtOZ0w8gk3JS2lR41r6ksnWdC7r5oF54JHV84LATCvAGoY
ZFLAWNktu/vYBdXE7D67d2sAGKlIY4Y6PuFysgic2NZhIjvOgO9JsFHcDtq+FFkhsrBZjAC5ewmj
Uub4fSATeeIYZ4Ia8ljQIC/2vCkfIOjzvHM9cHGZJ4SQ8Ny54VguqPE6Aj164+RjvNzPw2jf3W5t
QhLox48sMtCoRRIgf8JkymDiDxEaoSZi150WC7tWSTDs5h1ZTAvRTE3VDnuav21sDRfdfI6IpGTS
wWJaO5lFJKKE4SJdwiD5ksnVCGWBewm6SNioSgVlZsBFGAvS2iHw5woLNGLOLKk5CzrFN8tusDWs
ehOFRAvzg8RzRsBj4N5RESRYXUnNvd3MgNyFxbQ6yoMkHTca96l37n6FI87uX/vDwZjG98mj/qWo
556GppCvxWpQtrPFOKZETHFk4dnIthxpTW3Qh7k5MrdkGCOtg+KSeOGc5azDsGEGOdGzK/1BX/en
BwuXuRSW9XRqM/dUUM7YPnpIsyLyjDdwpQBpFNeBd/CGA2XKdD7dsE86cb6Ak2jBeApotLh9bUJA
pub5nsHIMrLFH91C8wuteU/qf+rjfIy6TdCyUgy1csGZiemRc2TC/h7z3bMLUCE7DvdZglmCWHdq
UieRUJFoHPsrrdNARScvc/T12RT2J0kXuQIiKREP8OfUJvBX8MifvMVMnBbmiSaAzQD4oDY6LTeh
n1VMVFY3yXyBN/F/NE0SwobOuHSU8YBD869xPzBnLM0u1UUt+2i4cLAXui454oT48kk3L64UdLre
1r6ds3foAE1bLucnVPuwzq1UgdmeIqbJF5RQrcqhy9ZEWXo1oSpCAFmFbzRWA6mLqPOlTaSF7nGf
CHgbJqGsxAwWX/NlN4iaCuNJrOLtbFAAK0eRzkeVQmXc5PtfDQyv1xhqNtxXNpRmnls4gLSO1Oxz
LexmarHLnrxBsQK0ZrrOkT83DTsqn6TLlDPFXQKtU4E/v476l93eBtQKMzOWgC9QpCHaGIUP9s4c
DefXJUMNl78x9Ys9GyONgFqFfNxAZvdMFjbsrn39jbTfgLt6GEDU+d49N5bMspCU29Ck/RKH2ZbB
7jxlQlzYrh1t7NBvgY7A09Mz1QGr1/vyxtWTEBKOzsXnsPrvh+buTAGrSEglCKCJzDlDHr2nal7g
fNnVK11GmfUHboA3BlU56iSEzRr/ZKR6rg5CIRT//ShB5eOqdthhPy7CvERgjKjYVBV2PK04IBvZ
hV3qq5PIGs5enwbHseCYglhG9MFfUpg2JZoq0DQXZIAErSnSdUJz2JizODjpIG3J43tmxFiX6fKk
maKChJDAwOGGwK+cX+x4fiY8hJX3NME+4QL0YFl2JwE0Vec0Edpp39f2NeHg+izmI8fnZMnxl4ky
epRwvS2A3HwAmYLQqJbm6LSPxDh/pa5aM56JDyYsKimSSG6DnkdrHsQM1Lj3NltXKmkhIn9kmrPS
54hvAsOL553EVXtWge7nUDZQ3pCFdc0WI8NwTn4GaOHFrcCnYCWK7OYFsd/ozCGeV3+EaJcZQHiA
CJgBspgDtEAJ1pFNWDe+THA/2J78jpNpwsJU4/B5YDqg3GEleIS9atKz2OG23OtcmH+qCn9WRJTF
uWZaQoNM061px5uszvkfq7oo2E9DDveXGMl8iBaLx1PRv96TsY0CqRciLGacmuaKVIFUAbSDU3YP
FiPdfHmU73aMhx2taYNllW1mCK3MsKuNfL7orn9O0TrRvcDFnSQn/JkKIV6kzU4xQ+WFVCndCxbB
Hs5bxBcyv92dPHWxWGlOvvVrCk8nOPLn7Ik59NLXLZcvXAUnLYZ85bX+qjJUydW+hZ2AkuyaGuj3
hd35OJnm5jBpIORgE+3Fk/yWMLbkmD1gEKuDpTqvOs6lw+rwDzw6iuAwsSEp0PXbxIB1nz8QGiwk
Jev3FaEOHCEfyBrXNI17L1GEHMhOXgZYKoCKfEPbTvlgQ9rvSHvPaS903xyM/J9BMraqM1kjRD38
xGcK2sJH74C8rRA57DuVrPhRvkXK7NRu+uNZDBEJVQDn7bAJF5h6SaQgtC7icoPmBiR0jdZ17GR6
uVhI/KtmwSk41hzqShaGntMqWX7aONwOlj45Dj8G5DHEvFYt4CVjfI7+30CWU6MEl0LonQIN+H2G
QGtVeYhAKLcdgr//YS720hswX2E8jUEQb8dAcOWRe/WnSWAmLcsNqvus3VO3GJBRU3SVn9drBwM0
W11aOFJkXdLRo+/zi3ASVgJ21qDOKxVqMnl6vyW9g9Qa3O4QZcfvZGQlfw5i8lsoxq7bk0cTwJLo
xjkO3wH6LMaWFNXTnJuvfIinRqW8gql0qmIWgU5beMyZ7dLel/5zfIhYaUHtuFdhtF/mxjhDbgOZ
vyixZHK9YPedIogJC/wXfGrsc5g2IjhGxqHf6Ib6OwEDtbWfBeTUaou/BICpfodA4pGrrpbajS9K
WtXmgw3oL2ZU6TFU6cMGUy4h6oAz9nRjVq8OLN1KTZjEtkyIj+/9OmF8nE0nfHdNHB2oo+o1EL78
b+hDIRi+vUz2FpGN/xcCkrbcmyegrhNo9mR9pYddV4UayXnfEIzSjS1w2zck0rv4Rm9IaBpK8LfD
MNB46DG7poVLnhowJUhSb+O53KfghjoR2O292YqnTPbXq1/HObkNOlww5S5zJHe0mLku2HsQ+Uzn
/PndrMa6bJCqFdWDcB9BwarzB/NV6nU5KLfLH7biP5UNRnVLqolZxyyBAv8WVDhcgbb/CgGb5CwF
Sc/kpRKIoKQc6uqMpowsf4/9ESB/P7zNRE+io8Cs3CyAEfnY5O/8nkYfFIycc3tFT9PyuDY5F8y3
Kqrzmepa2LuvIcd59PnCZE0jgEBuob0gUjMGtagAGIwfgrcMGzEeRFlCiClBX5zx9jzK1IUm/7NX
T+RPuKIQldtM6W3cYoG85q9dAUTR92myFcbmPMBKZob9fzNfMiF5d0lYpsrz4zYqjXUMuyL3rxl/
qSG/HvtptJmeq1IX5RGIXL/3Jp8Q7tY6BFEBLiHX7veOcDghmk7c2s6dvZZK5HUksTRFMV81Iubi
NLv92Qy9HhLa1dgr/5Qwv22UJq/ctRMfUs6J1EhYUlkGGw2orDTe4lf00s7pfIaVCDFMfOX5cdNk
/oKR3o+rQD5SFPUoSDof4EDn1lP2G0qsOZdRM3YwzshnAEwF/lrCRkzlJ/qsicg0bVm01+WsWu1Z
Xq9RKfu6Q86N0FsVOjxDwYKVQbGRZ62lRVQ+/jOimDvcU9ZLTTgP7PeOvl7lKnunjinFWaisgJZe
KL4OMqCa0ZI16nbp0eKAMXT88Ukx8myEaxy4Eht86+yNYR3JXO6mDEiaNO3a8gEBAT2AOP27VD3e
D2OTQckfqi6cxldQ842AllJIKuBJdLdv0L6yS5p4jwiCf+Keho9s/SzlV8sj0yGfZiV/g2dH0BK/
092/rNJJYyAlh+b0MiwrOY5TTvUSwtcoZUfSZW0FuiCuv7vf1jteQBDDs2FF6Mo+wG2HEuQQeCKR
dULWtix1Bw4GW19La3z2kXRlNksXlV3IuiwLvBzzFN9AIOTzluTmzAhxX6rmgg+6TO3RYt/5ntYX
CkqiXWlPOBnE31JwmuDXqiGjerLmUa22Q5Rna5cX5mwqOfolLQbUoh/t+qb9xb4t5uR6jqflWtbu
HA0LCAL6qlIPltcjfe4ucGt/AkfgEEKH1m5g4mELHtUZXhbrmP+yXJZksg2osJplymIBV7EfUwOL
8Uf2lRjY9AyWgBtjlV2BNhuZVZVwmWDEr/smANB7MNMdTkbupXY8rrZndShGOTGf+zzB9Mjzy0vU
sZwYEuJsvF3oLBylix8yFHkpAZE5BAaTYGuBRswv6ek9CwkD3sgqUO+2MnTqjP/sFu8zkLxOZYFB
L8JixR5PFDHhXFhICRetWZPPuFzMRTMIx8H4NIGXL7egNquVs+kvcQXiQcdm91T4NoQbX4TKlaMT
OazzWh9+GEmBFlDm3rdtB1ogDIaMLaqrTDgh6uvoeg4FXIMfS7ObmJJwV+Iz17eQtxCWOcD9hjxt
RJkC58TCEYURNctXMqU0TUe9bK22wdgeNgbzomMqLBFAHYRqHuS+VUgp+Gpzhp05cUYiUaAE5V0Z
MwoSJ1vBvfdzvwW3k4NyNajKxjzzeN+WUXrKQD7yGNUlcY1OZdrS9eYV3X0djkrTjMnUIxV+GA55
ArtEJKGeA8ENeBSWponNLEr2rHJBsIsDlxj9t9rF59y3oayJBAjaurFtGDg2MC0hylDEDuncU0He
aXshyI1QvHmwxVypAIPMbvHaazqrv13S+8vb/asjwdhnugug3AAda9kR2evGg854ggOhJa94l7xC
rsBhzbPqekQ/7pkX6qnJADIlogMBiH4rtG2yw/xaIdwRT8o6C0jEVe+8uYDNlV9tDi18gLEflZ9D
UCIZlmV71el4dntepD+Q+kVco2dR+E3Z+Qd1Zdw4ZUX0jJgLOOKquspkeHQXiZqbYJhOm8mWs1Ac
XVw9qrdpoqATSTiyNwelBU454RPTZlEzi5GBehVs04Qv1F+4hzibdd7O4ZeoSyR2PVnLE9+NPQ2k
R3w+FNqf8A9wzGTS0VWEgXoNS2bdfotvs/zFrvKb9/ZnmpcemQxq1XclVeW5IKKWyCqusVDTG0aX
DNHk8yWme2OxZq9+tvzB5VOUjFhdM1629Oyt3Y0xf2LmLI4y5RD3IuPi94DsrWSF/SXHUs927Oxu
f7glnrYOArCD9jd1rWSu+K3GISfoIk6hYjks9hZEcvhvHl/Q9G8ff00WjfrRZV66YNFLCK/IDRZf
Z5M8y7S6Q1Fmb0RMNt/ITInTwca+SVWFz797Tm/OMlwlG73pU1cvpBL8r49J0ynA4WRARiP72qV1
Yz/hMwGvHBBz7Hq5bwDXNjO4x0NCHMBgACvwICzJbB/JVLxXpDMicK8HV/ZLgNlUfkPWxHJOjlBq
8UHftNBFX6XOmZrCXXDi2ev+uSX4yLa0DciSwhzdjl7k/ciYoqDSoSz6fWFbKVIL15y+MdgMlAEq
qurr1QaRcBN60rGZcI1L9BJAb4hbUcIb97Cke9n9ulzdLokahZKcZOe8OEzcNkRRddZPGoIGjdY7
llTi6I0EyYOAOKKZ/gL1Ktd5K/0htaRq3j564YHg47Q4LjqPMhUhVNcrt2kSvnHabLYI53kVZ1qq
Mu+ouSuW/HxDwe+z7TWLA/kIcwYNkyru780zWww1sZkMu1zTlKDkyv7GrDS69zNbsrgacBjqhHJ7
mD//hjCCIBvdLrKY/Vpjmbk5W1XeCHgIkBzMLu03oEJNFWXY5xt7qSN8ULNCefWApgGdQPYs8xjL
A1pEpvsEm52U5dqdm/HVfsZ7Tl/JZgeXy2SZtY+HyWz9c2WZerr+vQSSrNasdPVEa19DarOn71u8
LOMgzKVFw7w+M9Eu1fZanBiYJEunXVQFYK/Hw3KLOZr996nh+ze0FoW3mj6KJNL8enmbrsA00P47
VUHwKE1xW6I1zdqZ8870ZSd/Q3PLTHiGrPxUs6qYwEslRbJd9vu2fMMR1Xjgg9lqXh/cvw76Z+QV
uw4nvY2tqW+ff+rjPjxoeEp6vLQ+yrkUnTHQUyGbl4KmiOLmTNe7quFMI5Og7B0HnQlMFHDI/04w
cuQxqjkJ8rZMCIVxHNBPTjIZV5c4b9bF6ybILWYsTMzYkxa47Bh6ZP3WnBSDuVT/hmJMyyis4MHs
h61T/U3ONJhdHPVnbNeYXWVKVeKDBIdNg5Om8krbHOGZim4ef4YhV+eC9Tujwa9mC4rq8NQtf9at
T8De+kKI+mQgmD0/Qp2H1DUiUp6ox9hfmX8NV33lFNFDGz30Y3F6CEFlrrmElwbEKQ6WcQwKbZxJ
XQwOISzhWSqpNaoC45N3of7nEruGV4vzqLQJxmjdZhLgo6ArIfbLHQQ0K6Y42dTrOG4abdvpQy7s
cUI6dhsLTsY5LbS+PBREPCNj1Uv8qAb7olbafKT6r90E6PTLLJF0LbYn4PEZOz1dIbHhuGeDlkER
nT4o2kBTZNf9FBSBgJUi+b/IjANRNniIO/pld07TNi81AVM3Kgy1JGfjjBzLnhQx3daiMs/BQwwb
8/Sh0M5FtXy2NA+KUjxugE45O9oAWlZpg/jaojlOVTIvVFfFr2cU41IVl2lXNSVZVZWv7hVl60k8
b+xTO99/Lt+Zo7roUUr9dbhI43myLknXkAJTkT8LiBZvxVaAHR+F7hp5HY6mYoNGEUMgoaAxFoM2
p0wFWcypBT7C+5qR+zrBTCvF4IF1XghgDtS4PhWtx+xVvT1q6nG5IQvEQrt2jkCNktc4KpKBpWBN
L7iL0e7dvCTl5+Io62bg2dhwFM8B2XnYX8PkGHYR9L4AK9FF9PtYKCF/trpvQ4lyLm3ftnZB4JJF
naOhATpiNwAu4T8brJsVMWN54fHmgztfMnOl80/Xw7l1whsnRVwpI9kUiBO3rTL0rYSd9dM3i7Pm
KGZ4CO2uWp3kE5ukZefINr3WbhXaWvLnl7FVPZCs4aQmMfRYYpaRQaSA5S/4RzbAayeSRk5yweHJ
HS9MGZGC64f5FwYbgM90qD9aVqVFe0lTwVYzXLUUrWVWdVlnaN88CjeiSyfE9vbM5Gfz6IugsHfu
Fquh+2i9VxcF3uDMluF41o//n1KHFXGp83FVeV67uHBV5Iqg/jygwdvqEUhLt7VAu8g2RwFtNFdY
f1O/0jiAZYNvblF9vaegMAR0D5fyPEmC5GbHYd+n5X0u/v0w8d/VUPRhCWH3FVRtHRDowmJz+UQl
Zjmm1RM+W8Ie8v2x9k0wNefkBDwFa7XINrFeBqQnRrrnFxLC6QIf6xJjazA60L6Ai54gdQGayJDl
k3445ndqZCckay6iccLnNxtrUkVq3t5MFQ5gQwXpwxze23bEv2F8bqhHH9PdRZRyJRIE2qNVG0Dn
wnj105i9v+GboJd+VYqqWc6kME/TW/MnHjYyhp1VGAIfZO9OxNEe9tp159jW0jtE33dyaVF2WE5H
VpJ2xxv1j1qYWeYvP4DzkDS1UoIl8Av5eTlytoSNIUSrMRkLw7G0tAQATTtNbxeroBrCIIP232Wl
PbFF1CrXFbxKGOahpDfYqRekbatRxSTBWUHbMrmCzqbp/Yu0aik2hw/tr9RWOKHj+0Rue6HFDCxC
VuOmEFxAHjhyMe1BoOnt9EqYR28+PAjnkXJ/6wp3bsy1rg7n+lDZeGr6mPL3jfAoDtfvFOMddr4r
mDLt6gM6qB7/dCVRzONYMPOnQ5/rGxah5PFHLFUXblK//PmUwUw0y9NY2ZPzEWHMEf+yiKLovEWh
cwf9IVy1oI0/Cwec+JE5uJtZun7tJAvSm2ZraINhfTifa0+jz3JSub0D7EDepiUn6TTN9BH7jbJO
UOPNvGW3gyKze4/c8UW+slvuyMMLt5ntYSEbD7MFE4P5GxNAKuGqHP3uCj9L9lMigxtYbAYC8A03
g+wrdHd9UjJqEj5JmTEAuUM9akk0KBElQ9X+89GWGRVf7T6NG0sbXVWMwpzJwfvonNiZ0c1r7Lyz
KpOntcHEU4DGpLHKTe3rElvgttTNmdasGKJ/VHbGUxqhG1EjntrakLfU0JGMDA97Irk0XrUgpfzO
/e0RR3g6Qs/o9quEBRVJTNGClmA9Z+JsQ53UPzdfM6tc9EWvKSRIUR4/jlSsuh5xnR3mS+Mgy2VN
HoQk5YkEnF5JXn9h1UOyo3LreMlKTGh9cE9Nd4UNwK7NRhyAzS2NCl1VY3eCcZhLro1ngcD/X1Y8
XYmdldOV23t3HT0IV1AigY6d+LCsMYCoL2G48vpG7BQCEi/+3/o7X8QmLDcwIfKROQ3r/hbl+gxQ
98pwjz9pyzSIhl5kKTwFfqv8xzR/e7cXOqubhEnzFAa9xxxDZ5avVqg2gmdWHbc6S/Xi4aslDmYK
LsQt2ZGtGOXq4N0A4bikzI5pWpgS7X6fP7Jv3la3O9DW5JMCGhzGPrvEiZxCvveZxrXH5hemUivJ
dR3TRlNYbZvCCLBrE8hjQN79kdJD1WCfmDu7w8B+MfV8f1NnhL2Vj5/uHzgh+TpMyJEwqpBX7Sww
P3mdv4CAIey4f++WiFz/sKn0SjkJ1qIfaiLQyBR/1dZMkBzrSrE2sujTE1kFH2/g4iP+Iyz1Zb1f
CZ1dbgY13YYf/Qi7dl+5mDF/tiZfWu+LeMR0jpjE2ZzwLc4sgjJCYgq0xatBi4bZM8kr5rP4ljhm
s/SbQoIoP1xQOTDv2NlBq9RkiEKsWJgn7l8Cjt7WH4ui94uUrcdO7AgjbqXWWesMcxZnhEGD9Z9y
KsbQkPx0+NgXmkDr0TVDo32sjwj6xBHeeHRmA7/hFblfEhFDD56EPlq6zQsekTm0XpqwvhYhx9Cy
OFeqFm1wlQA6nBsEWOZ+nrvm/j5jXNNpCjaukFnyLYFoUNSRLbPqfHOBFoF/rqNvlgb543gAWsb2
V5xfhj8HPIBNwmjcjwhmmC1vst4zEqBeJeV7ctcTZSfhS6h7XdD6N/IR1zFO8w7djjjSfH0QNTRg
OnN11Df7B+k0hI/p0/jfv2YmiovUgocRwKHg+k//Mld4HvD25+Yme06t9dDFbY8APLlRGD3HyqVW
NeKoRp4fkrK2evIDcOB0mQUy06IzJ4H7v/n8gEiUl25oaDQWnKl8oiKtQb863/G9A7WRyvfBPUQJ
yK8wzE3OREYNCfKm75BfqlJYf3OW1BtPdNtfIzwCl3av6jrFKo7UW5teJQ8ptjoZASBi8OUtaB/n
Lw/Z822YO7NHUmzpksDU7MJiKeCVw8PXpdG6xCfnQx111pnXL00luPLEGYvCL36mIA1sTe3NYVzs
IAeClYgg5I3UGF2P5MOC32uIsTYNXrZLEHqDIBi2E9KbYGE23psCi5cuVKz5WX9KC/xigOw3sMu5
z71sI8aiSibbVGltLp33LmTknEWbaRt/QESMlFtEUM2rVlLiqN9cobY4OA85pYOK04OzVsqFvuQp
0/udCy3raiMUbdsM5cJnpachbyRTg4GlynMz6fKCfX0y8SVBLBJ1I8euJoDcV9dJSYQAKQhRf9Jc
HbMZyurRYPP8HaVhP8A/lSMYwqhiwoNs/9JCULo98kVX9gWkjNPLg11SUm1LdDZPAEtUAIxDtU8x
06JV+t75+Q6R7sNsfTcztblM+bMGLNMF05lG2DG4jRg6nbvwam5F9GNVQuhspSWpHdygENIR8z0t
97uttG4FbHLVUguRZ1xUO+0clBQeipnjGlVZXZDOk2cR1M8A2YWa3no9kggmxlJ+gDhf3FYKqjww
qS4R1Gai6buhHqglgX7KUtM9k/n7e6emUlpemVW3lflBP+PkY9Kdv3YE6Rkg9M3h1Hqs/hMba4XC
AjM57IkwMUNWKSS2lOvRDZ3dHTUrnwqJ9LIDj3jkkjh9urINdXqSYC74xerHaVUt9R4p5mdupJjG
g3H6rJ18mzHm9Z872GxBUtvennpg/LIg9OOPzq51MSVFIrxsvJ5cwwjqSRYjRj5YHPMnyi9sKjYZ
PPF7mnsAqtLmn5o9O9clmjORky0EJFSglva47fzvpdIhdSi1gVO7YJK0nqYla6hMnyvYP4sgRFDa
d2aNELOqh3dRijSXP872+CIouKlCtjKjHgmvRrWWsvC/5haSVCD0E0XpBuG41pZlLqO8VZI2nw0K
jzTlP83KD0eNnsbxOV1XGUgiCOhsbxR2pPUAcD/4fmdozixYTA1SiZbZ9OTVTJDbC2h8rfJZT6Mg
isypjTi6OPjz/vX00rPmp54KJoHIMqzlSaiul4+SYYPmUNXcdXatsa5mdimByCMNlbf9bxuecoYe
t2d8Ab1QImCEGC3Q4Tnzvj9D+K2Fk4+F9ICsbwDLadRZutyWqfaIKuiVrwa+JAl9Yh9mE619sHQ4
wbfMf7VWDR881Y591fQsQ8CPBTzZe98f25FKmKVWsi/dVAzniN183v8nDgiDHQXvSqBrDFs4Ipiw
mXu2ApW6YaY/FrB8NJpeIqmaMew0380je885sfP5RvoYEVGsa27A63qd+6IF6Q/ftNLmrUQmL8gd
/SLqIuXYJOIRdOmvWCvoxoTovxzPF69DYJJhHGsyRB6RQkUHtrqpuMN5/I3cu9qaX1sm3B3esi0R
Y80cQO4Rk0LwlB6gwTTLXibXYpt6IxT0e47SkdB26d/cmM5h+tGJomS6+sB1eWxziAKMGm2kvowF
taHviTIYaP6k84ZczZuNv5JzWoHFgY7uWQUNC1qNgePFTzuhK62FelabwtL7Q/AIEk4ojMEVom0A
ttdt+hAj2e1XeLhIZFtzln2nEjBpZ8+bRopUix5PvG9ApDyAPzH6ugR1BTm3goq9PPUw7Mnm1Xq6
81gU7K2fuVxDxfe4aCJ5VsSiXX8n2cIOkTKhK/Jy/MkQt2xoRli9iRSU/OYRoq1CjE61uTTpkOv/
9YbaCf+Y+EcNCCCWRXTJcFAUjMpQVlIrNAhIXtabeDBW2S9rWpSBPmpD3k/zy5573QS6u9GoQfpC
K7hoPgq1j10kIjZogcyBZYhDoHR4GOriBxpzlBM8HXqtWlNSszxtqCISta39sC4mGULgEt0+8Tv3
6Pd/WPaez0YaNpclBAaeIveRDN+jc+F8ooMN3mh91XfMpAaGfbVQ0c0FXMOUTb3mYfDkxiAKRX9S
RSNd9ouqAfoGxH5tu8IjKLNsxNz8KiU9ra3zF8+UnyhoGQREBaD7FTxg8pHWsILkHDdh+MOdsSbv
oC8VPDGar6BQpyPOPoAxamlP+6KHD8TX7NiIUwIxc/L+YhOL2LiHRAIyVdDUgTBvUfws3r3N/fkG
k6abcMrE50jEppULsSGZKpkYkO8tXyKPiVwI21qltcbNuwi8o9NutENw5uQADQYQW4yJQmgsq77p
ILgPZLIL5KvI7dWT3K/vT38KJOcJWeu7pkCz1/+atrpK6OTivqSsT+1QHUWVjTC/c3c/+wzqY8vu
uxtWhxbCMGzCcZio4oTEqaTCpStCJ0ySm7oVfizMaqihmoJi4ZmbuGkzBfqonirxGCoBJXmDGtx4
zpzInYwhCYGjA07jsJy4DJT58HE973G++00EiQkG2akFo/G3/FE7/O1DeqOvjOgEmaeB3RlwsIHL
8szCi5mrtMy0wV14YmvqEOYJA2AZ75CjG///E+pMWb2dYKMNOMc5/llsTeHJieIzhARAEdabqN15
NHARz25Cs+mhqbYxH7sttx9zqVgyuILfMpt+g2/lbpCkKtodtN4yjz36exS8JokW6yDy7GkPpC3T
E5TF3VKhFceXcc/EVZtWk6aPM4p9IidwUwVFfxvPTG1lMIqS1nj3DOO0ClGqHlz4KKGP8x65UEz8
zgViCgr59h9HDw33howgzhorVtHUnsEkjRB7B6goIcQpQp/NfqzjuD9mPusCbO92ITIOy7HcZnWL
QCVH/RUJ6JSn/Ekh1i7RQhldstCQNYor0XoewlW9Nhu7cpx1O9k3LGbCL9S/aq1+Sd7SaIDBLuXk
1dg2LG4x0Tca/u56uUovdq4PD3d3dNT3RnquPoP/gME43cvcKklSS64or3hyoBq+GCAY57yEReUz
sKKzEqPa7yGwUtz0X569C/hyokcFftZtuc52D5a5WLCx4yi7L9NLGDrwOju5gmH5tDNjiynF28aE
tsS2MTifAeF4Y3tQapiQBznqrguinzlvBS9dsIBhNta2ThRIvGWNqMs+WeabglE1nLgLXRK8hY3t
YMOi8Wo8VIjpqtBt9T8u+3xCLG4/a8gSG5vjjbqH1cOfOPlsZIuY+SaiCWIFijAXzKV4bKJdc3gq
Zc8H3EanR+XaCuX3yCAAqDknA+1dTUKuElkuFyXpo+IRXVGIxlfkBOZ3Ws9ceNRZbYUK7j6HK0Rc
6i4r5nD85K+e+IoTbPKOKaHGLI1bEYbKPld3Wu2PWSZ0Ngc8QEX9DSujkpE7xNVjAJnyRutos67v
2Hxg7ZqU4E9K2FK3/RpMO6b2fCwYDRKLohgdhZJ9+NbBu7YA595Wrub5YAPN6FISVZzcVIA4QdiM
UjmmTbFM5OV0Oq4SYUjFvBnGp5azpMtOrhdkR2c9Tbt+PspYQKyog7hD2kWAWRBzazMrKhAIAYrQ
TfEHNTeujUkAOivn6zo14DH0Vb7eBfaLqRpGbdMv68kslSyf0yI2LjoShbAovVOkylvScKIe9dSz
5oQYh0mXRB0KR+uc3Szamu7lFyItR/KUE/Sy27Ae9JEm50SARoJG56968vfDzVMYyxF56kTiCfL9
32Z+ipbMTO+0BzEeH+C8VbVy0p2imaweI1XNZeOmBPJB5a8R1v0mvnyeHvp3A9wPA5ccj5+7s5qK
3uHdJ4HZCiMNoJQdUksoX8Uu332bUfiNw2C7fJTgqLFXvqNxGMRJ/gI8exjLMmsi+qzmS9Z47YnD
whfo9GQ4yukGpA2CgYDBqvwkkMUgPiGeGtyvVep5FYySScSt5D/FAfdMIFNqJroBtOaX+XwAZM4p
DuN7Ue1LsylIwV8gTxi6HuanXKkUZ+Bbgd6aCPUfFWGoltGJA2DqiyB+mJMCXyl+894rV7VvWyRH
tfhiWe37Jxp+csFtwHKAIqWZijQYHG2Z9KIJxBCckXvNc+I9MtkYBrlyk7n9XzVyP8TZpchklkmk
uS6Gy4W6SQ/IEpdHIixs6uZx14Lv64291YknxogqMS7ujI32tvFXg3zrwzyXcXGTFaDtxtU5JVtZ
Am9vYVEh7gLZ9t738rlq/eavYK+GJCPgh8lc6u4dJK1YSHy9WkMoPvIe/vEaGcfN0G+cWxZweO/d
XaL2Dg5RpoVJmMQ7txGOJdBCtw1A1TRU9Tgr1dNpDs6f4hjufC6mwus0xOYjvCkSvBU8Gf4BFafK
f9glQ8He45Tz3Xg482DrEH4hCdmJBiPB87zYX87XtZOG3Kd6f6TtuhKclxa/7PCsUQ0STFx8uWxI
K4d6w1Q5CY7LTve6VAUkPZ+djKkS7+6XqNoYDvDDYWDPYz4GBULB7fXJsSnWBPxeSbf1LnrdeK2x
dmCJHK4LcgH76xL19XDmzYCjFYWhTVdEcACH5qKOrmXvjIwWlj4jh1Q1hnmw9lHN2SRWjh4RWB2E
tgdlVZIEwaYhVwmbVBIpHPNMUHhKZALRCjgJviZcca0RU7aVOwNfoRLUQy51qfLaEiFCYxoBQQ2V
Vr5pWkv0p/vQvniu54Ecfi00EYTLz0GbEojx6AOt404hV+aMWbNuguAoLB//hth75zJ9sxzx2vJI
HBan5qjYkNWOF3upAeUUZzDdgRyODUL2jSByXatRreHnSbWorMT26sGKIVaRrPs9bpoam013OEZ3
VXN3cMCim0CdFSLfjp8rq8B6P5UrBK8sf5T7NtOBzxusKKKXaFs+77gOKg4K8jL/n9G4Ir42869w
x6cQZP3DwrSuLgSHH8sejY75mokqRUb6UkyeKEMA589HDUYa+CI0N2fmzkb7nVJTKV8Pwq3PL20l
rjxK+Ado+OBDECU10ZkSBhePq0RqkxMtmQwgArfCZHhLadG27FUachUYnO8K5+n7aAYW6BEPJjhO
9ozaoX5qy7j7LSeCdWiblpwKZ52wEl3M57+X8eYMwNwg3V2o+4IRmpq9MIIUIyk23sFIICoGc/Kq
g1iXHITI0zEIOsDjqEfSrj/C+l29BYyf+BK7YXd4EqSa5O/19KijOd+nhCsnpbT8yXNrh6RE7236
jbXShpzbW1U1YJp+gSLfFRHKqnUZ1P+GM2u+cruaCrEHg74u3H/+U+CwhTyotD86oaZ97OlZFsaJ
UfUFswBhsJqGanegso6rKPn3FuFJIYmUUfNiBhgG7LdefeAhDsCrDw9tfftsGzAkoIxQYjsfCjZp
UaIql5nPfMjTfbBl0w1+wy064lsNiSdCEQI2oqOOR1drW+RKk/EVSvK6cdZJ3tWBng+YVQcvMy3X
kJ4YfqX8zRdn8TDYjcfxcKkoYEfpa8dE4Sb78jGaZ4W4Ob2ZXvSbGSEGj90L1rFe/RUXSR7TGX1p
POPzWR6fnw2hwwKRmq64zhyIAkIzINCz844EP5AOg2I3tgqEKkKXLrcD0cuxRMnS2RXh5aWzgnKT
Bdt90YOo63eKIOv7Y3Ma62D+XtYcarat14il5sxgUNQMoU2O1Saz1BKg1fxSFhabF5C1bQCgWIxa
OtyuNe+lKuJu7WBeLGGi02AoUqbyeccbt71k0oQVDs65cJg4V0+kEiMSoQPnRefs1aFD48DoTnzJ
aIQpDGilTBCNmiznfisKqNLuUjtPxcAp9gvjPIknFYgH2GRmjsdh6VJe2DMz/emoNWp5GczZlPYS
LfNT33qEYI0xTaM76gqz4VvoNmoop2eTrfe0p27ji/sGFSpmUvILo5+GA7AdkNlqzJYvovitVXzE
s+YNefCsUcUV4sxWccM9pYaRLIZ28xgslLubCz+999CbPT+C1y85PFl6shF7s8znYQmgiCltiEqH
RHBmHSfs/vO8PRhpZS7+bVuKSzcygeLjCvsbn/06TM23OIQXgutNnZQuHyvvoqRwMnHrfim4VmLD
UtiwZlKUHLMMNC5Mbn4owDZSkx3QWvkihCYrrFk6v6gp6JlQzUaK9HEF7on8WW3WsCRgtjFSRV4I
MxfurSavXIImksDZ1VmUSARgWueacloGCybMUAu6GVfQP43vDUNhPdF3vZmgQme61wiXeDx1e5jK
8HLUqLAi3G6sEnta3qVth/KB7lPLErZhBG08p7Q9QCAPz3qMI0oefQaMXVDFgONWenm1BnJn+euq
QQ3jPjo6m4on08fheHwp9sdSSc3nrK7aIM2PSUBhxM1u0GpNLslMx1DX7YZyJL54WbXHoyjnzZ/M
Ym5K2vQ93f5cwX6PIfpuhRhk/iaTUszl3zDzgJXPplzpQcNCSX0nHhN/o3RwHBX7i2jHRimwzngO
ecxYzZmDmS+bIM7bryOvfAIjdlCzeLMVhzFzXps4keTsLuvNr0+JveuK+HlA5zYpP8ueJBDBGQ0l
xAHplACXIlvMHHTU2ygbkNKtsNSMNirAUbkTONDDdxEGyoYOmsHgkoLcEvs+kYClC1wPe4x4A0I2
Xq2+if8vOCzllUA815WIGzeppntKRxOdPWZQ/j1SKFI2Be8R/aON+5RE3E/5epiW50aOdWpaFgBM
hFvxmww5vGcODU3nwoAdV9PcUi1VAZIbUgom7KdLpV8nLrqJQ0Q5V49ooyDql37e/F312oHTJEeQ
ibUqGIlqgKVFFunJ8dulTrQwVK4X8W7F1X8hG1L+vAUOvop51jOgVvbejZ8c9qWJJKBpvUGE18y4
q/pkGhBSYoPXPf6PlRvkdtJ0UuY7ADLFGvgVm00mKAKEsR6XYo/QbTmZWqTtc9LLKFNojlNZNkW1
u3/Bbt9GcT2lbxUhrB2xQwcQDH/J1W1lxwtcPMOeGzcK/hyefm3D0RB+88HcWfFpu6sdFDB4XmUd
D4jltPF3al51rn95tsML4nuWANRSQuRVIOM104OlhPJoNEq1NzUHiSY9n3PIScIjoBQoKGKyDM17
COwOpjhTROHS7OWoxUGjy3AGkxNmCi4VvtePf0VKFpSTpV8Pr9W+QVqK939yIBLEg7yRb7e0vi1T
7Srh5H83n5eu/mB+lE4BauLXD2d4luHgrocWOA2GM7f8NHSuoJ4D7zNM/ubG4GTkQB0bvlcKx4FB
qpFowdrUXJXbotfYf21Dz5nTE4CZGOwJlG6IznYqtCeHuUlBixhS6vUuTOUBTZaz3C5T6079eo+C
SyHAZwYJ/BVxdQQimsMSbalSuXSTnWHuM+cX70GwsbQ3ouz2C1OJpzg1IuGZKwzyWSk50VRZ64I4
ZxnUO/6TIk2s9WAtfTi+t//Fk222CeltTbLPQ3tz3toa/E553/ArsC115fWYRwHSNKZi0PwrHcjM
xuI02pFgEjs0/cv5h6O5IAw515VPcJUo0Qw0uBBEH+fAJbkDatg46n/muxNzP1Qo3EbSruNMIKiZ
Mti+ZsljYAq7EUYsKBmne4nhHcRJd8UXy9uZq5lZKNBNDGaQBlRvTXf5KuqNGgc9W7dnH8YOcGT2
a4osd11TSmoNhifIUmhqsszsn41XIDwKK/CqDLbK6X8o9joBScn/mSXsanovCfFFBu2ut75v4HT2
zfRopQ3bHCDlmVWc7eIbrj1cP9+mWi2or0cBZ2BYhUc/ohUKTej660WFrycMrHGcD0UklTbuaRXr
KA5C5M2yOd5bZ13xi852iYVPplckJnNZ3aDsXOBQ7jKIs6qYcppTaPNPjQJxXuMasnLImoBKaULb
yJ3sZC1CiKEc7S218sFW32GmmbMGilRXNaOxuZs48IC7++j8r0AdqLnJF2gfu/t6J1UhwPDAD/MS
i/KCno1rnGnEvOFDSYAp57TeWDvXmOujrTr6QlZnCrVeCbdntrWWqwVDxuyj2HF5OjZOMYe50E3G
356fNeIwKPPl53YObOSlZn5T+rtYqYMrQQIdH1iq4LsoUNdYBs0uEkmy8JeaK11obntTE8KeWwkQ
dWaqLIx3J2hSIQDUm97jg7h6x96iW2PH+OoIUKkDPAND3ghzpOH32oZ0oKqyawqGelq+PzuLNAHT
vZEKjh72DPgNknJAWEtv1NckE9EL3GbrK8Q0lgKoNlNGt3/FTL/KebBalAlkv/2mT9YQaL2t5GWB
+qW8oV+ZNGDUi/7aSobM/gLnAAl/22JGtc4ttCjl59bG4soXYxGvq7NddrXpaQpQ5gNaRjSPN+gm
6ySIAH/pIR13eSqJ00gYR/x5yM0M7xqTuhSlMkulksgE36N1SRyixgOWlVgq9IOBkzmxxzAD6dgA
+RPTZNWi31pDxKza/+0J+a2/XBewgDKDBn5BVR3VC2eECLlnRD1ME2vE4BfTOdIedy06sItRdYMp
QwMjN9Pb0OACaUF8ZG1kPVi1/vfHymNxpluUmXpKOFsI/yY+8PwE/kJ3ZMSGYYQY7Pj1EQF+Qa1W
GnX8kUO+RkFAOnnYV4N0ffHl4YThrm2xiwZZ79q5BG5SywofRM7eziPXaEDfpb831E7rzquR5jKj
NByHTdijs2YZJTA0ijUJXWOkGsR7fzcvg1cGk7ZPuuNmzA8OAdMegrMZ3ecf6FNIuWjYOXRH8MsN
te2rG+fUNtXDQq7/tlYte7wf5X43+yOkPNIuwEQn64KJmUZXbvwy3z8EsPZ3rn3NwRj7zKvBUSad
rKgU69e/im6Q3lenU8HPN0N0jvqPU6iAfYOcX8EYNmD3USquAlo2uZAB0+U6MezwJ3/scVraztNu
9fbG2r3MNZpDgFo3rbPUXe6DASUlfGUT/FrDObJHoa5lpi2LX2hk4aPWVWTvbgUlRRJUEeX+f0At
W0v9i45IBXB6ekJbuKfDRPqRSpoElz8BrrfXWF8YZA/frwVtxKx9TY+2+aeDnebo/dC1AyqulNKb
ZZbmpIWF9ZA5ZHXdUJVSRVEoc9p7lR1lcL7lgGMG8bBEQjtHDG62Akjq4y6ImiEghCmDLk72bu95
XkKs0ZHp1hUAVEWzpg0OhPUKXj66qvL6AHV2f7M2Mg+VSrQG1bYb24qQK6Y433JSCXBtUUhlTcmP
XFILcnbrDZZ6kg6LUs+k5CjGjPOtmgNMBwsNX2QAfbGfmYaJ/1VT0QQ6yJoABSHb2gzqwwl5RrPv
BDF/cgQ0JQbu4SPHCKUqUrTSPPiA+a0noQwIp9HmfzO6//2ecy/TdevLeJzKBRdj2fa2d8QtRVcj
tYEbOapzh0p4zVnsX/0KZ7YgzN2fpRRqRmJ8om4gTc5BHtvC2cnAkB3q/D7a5ImHrLzkg5JMMveT
btdj3m1KxHjxJGp8U8i9LASKQPndGsZlGAAWEM5/bo7D1FNXCrBLdVSg6p/YEfRjqEsPccI35NIU
ZJwm7sJwOFdTqmFrni3nQOM/2gf7uNP9ouC5A5N+DkYSqggMbmbV1+1NppBV9sMlJNy7bvCJJGTm
9GBUbtdU5t02foxFlLg6Jzjo/443lT8aq5F7WriswCyRbSNbMSIvlz3bIA/r9chCV2KuruCvsGPx
1VoipxNqgGlWqa5BrieD/lx/ZshVm0dq41V0rE17DMR58ipbKvm9dBhH7eAiQsp5S/MOp60wQ5m4
AzGzPQgpVOsbfFHin2n16N13G0WflYoKdJZpvHyjmtMTbwI5G30fjkP+u0c/oO35KqCdJFCXZrzI
56T8N4w4RjHifUONkCITNHoms8YM6DefGZhDPrK27EP9jYdb8Mq29GJcA/dQCBpOGVt8mr5wd9L5
9J7vAf3D5SvN86AiAWbxZw/gxIc5uBIjf8sEiOSlfCGygKiZaJxPfr1NR/aYpecm/Ew6vyLUT05o
zUEIbBnPa9xBzv0YODcWNGos8mHLs6c9QDyfI9tnym/6UGI8OW9gwdDrSCqf+wACgd77kbqA/7To
Sp/CrVBZJ4K9IVJHUbntlOSd57rvWNTqoOOXinOuwmSp8QfAt5IOjO9ercV/oJqBd10M1jgQV+Gm
a/qaBH1BNUubHnwr/FCOtk0QYUHOdvAfgd/lIoT0I8Qd8zOZjVs6sVmCpzBQ0TO/hlzjSjR7Rbjc
gGF3gN2YluJFxjiBn9YJ+wyGC1Tk0fZPCB/XUraZdZSBTWgnM+c8iySa7oN9MMZ8mOwcWMGslc8A
KSMKQQ63f6f+bOqpjaHcVjr8qyKGCmwdrAPGccx8/QWjo0AkuOf2Ikx60J2He/Qm1NjE2S+nqNo1
HMX/OBWNk1vPgx9fmvQzBJPKg24knSi7c2dkwzJ3LxgX2sDcXtUtSiLgGtokHnUq7JyzYOC3+nWk
s9ZC+yeDUB+SHGCFMEvsq6A9N0D0SQ//ESVxEJenAWpsdhu84ZaIN7tqqD4Hgo0QIGkB7OU4Rt4S
FQ4QUs99pkgDQHE6t4uTPRTQP5rG7BTXNJbzz6vrdpTPs0Lah6nuy/tr1+2U9Smt89nZLmFYtdlc
mp14Fgyta89xEFfCzo93U5unK8jCrB4MDwJZvRO6+7RIbQT7NB5c5z5OloXlkLWxO9k9BlvBAEsp
oQIrfqTj0aJRJuQJe676Z+0sYB1/2YNQAhZEQeiBnz2bEL11SlG0yzRZZWjDrS2AIExgnnnGXE6Q
ZxESj+9idewGuwRQuNqVizD69xg9JNjG2P5N1MPpzijCQGhG6mzgBe6ulaH+xxZ9FuV/yxlgPaKF
8Copd/yLMmqjZCw0xJzLZUIwohCJkDRzZrMtPHqiBIw4+SqS98w6x14Dg9vqiIQVPFmnqBQZkGnw
2tRn/c45YjcP+mX5rDeQQ76D83g5gwQ9fFLcjsSiKr1gUSOgc2LvBlBmSg2GJxH1m3MdDVjDU7gS
f8ckzxCtHeRGKq44gFunRA9sk2cficBnbmJ0KTin6pMAjWNqgCnd43yvilRSaUlAyAaxM82o5dXI
79ZX/mG8aiHnT00vcBXbWISsNu+m8V2QW5l7Z56J1PndrNB0jwGbn6Dy5VodE4yRhG9zj4qUX2zS
lJAB3cReqkCJynMYd3pMtJ9/sZ6s6eMlXLanSk7r5jEAl24q8dQFT8sQeB6DflNufLeRprRJBtoL
A7RqiTyrDCXtsovZm9x2IRksaIiXtmUYKaJujhUUmv2uR+x+2s9ltmKmYKjhBYndj2dZqpJAL3Bx
+F9wsMtObV/6rnICOzDAG5CkP/jx6hjGwnXo1J/rLNZxuMtewcAYIDqrHB4Cv0l2qzGy3vkrlWRz
OpUzYtd45X9zFxAHOddWNxJ/rT3Qxo8KY1yznNFxOvOYrbfv1+Xo02NTBvjYJEgQkwJvGTOnNSLj
cztXH4BwOTco/naOcwk+0MNP04l3zQqW9aDh94PBJ62E4o9pYqGCQ7L8RVG/r+ZGI8jnDODyDkom
aDch19qQXYmdRw+g6m8gVSQODRSfzMoFm/MTVLB7OJIfHFRwziHC5RGcML65z8pCNqyGqCVvxcGG
sfyi3rvLrj6xVt9DrT+taPMCtQpgz3WQRVhDHvRtEFRQQQWwXL21be61h66E2kSDqvibjPZzFuol
8gE5VnngGZHnd5DTf9W57RzyYm9P0kXXv6cxAKYQxj8AZJTx+BQE2Gn3YMGqS5s8RpzAJ7tdGcHj
c4ROadGSW1wMiD6hcYUXJj/QMNtjgtw2De0O5TfdNlCTy7/wiKVYDwaHvEPT/nt3AyrRFQKihy6G
3Soxkxnw1cNF7Me+io91zZ9RXKAnEi4q8mey2Ddq0fBCFm+SEaEqiRNMJi0LVHk2TJ/we+Cxx3Dn
MvPQqnY8lINoJ3MI2HQzENHNxZcj7oSZQg5cauFc3eud21sgRr+MrjR9aldr8sIpetfyebwLM/K6
AAdN51gXjHTgABZHl5A4CauaBgQvgj11Ytv6HXl20e3Eob+i1uGtGBjFieev9kx0iX/U2aS8L3ub
r5zhGIIkG2saLHyPmcEYl5r/1zDmrA+CkBebr0arsiMCo4OTe/RucGRFBMfhs+/TfZf5ZXD+jfSg
w2LJrCYjZYBYizL7XB1Xbb0qV3bJXAYVUcgjwi6cAJ50ua7sRJ/vLFNzjeb+puuXpZcaXZDze+Bg
zx+o7b2wNLAxPghAqLcytmoFp3uVTEHP3eNPG14BRHcTddT2b9ys3uZhl+CMZ+vJ6kclJv8kXtMb
l6WZHxeWw5yMVPaCRHGbtKENzhQ7czaTSARGNN0+3eXzwMTzSj7J7M8tJmiJX/ruHI1CueVNAjDa
EHlcqKL23xxVc3uBmfp2i3H2IWmBfb5b1TvMQSV9n2pPLM8k6wyQ725n786Zj0YlgXW7MK69UCI6
awF9z6WyfcV7UPflwO9nyy6I3nKeKMUkPzLWQ8gbqH0k+U3LFmBehmR+zFawzridVbIlpuhfhViO
9IVmUNnwk1eXm7BMn/kQrdXxS6xABgf/kqFVTZ47IPZEY5Z+WjfhI9wP++4YpqBlqp3GoXvu/2Td
t4Dj6walRcWhbD9eH+eZ9V3QJ8fyn3I2kx1O6+Dts3uluQCMZMDkC+WET70M50FuRjgwGsnBzuj9
Wg23Ve5tHD6aZbqnTDgbpa0oMGebdX0lwUMkZisU7TR02Ax7Q2l6fByOZMDWJuBas+UBElfacxVI
VD7HvXwc9tZ4vJsVec5ABfVmHqgFJO3SdyXC8rD89OieWqiC6HK+uRhznlF85INZLjpjZiRWCIlk
PZanzfF/Z20NOgBHcm2eUpea+/0qj+1rHP+mq+agzn6ruDgJyKuOGApFyrxewRN2pcODd5zn0rTI
2mZHmkZOSgwiTCpKKBuYyI5OCU7XD56gijdduNLoJAVGln9vDm8/Bl9XB5ps/qAPC8qmh2qe4PP/
D8odXh5CRekUEZJHwZhmD3By3TZOgo6nDklksrxMstj1ptJcTBonMY2GCVhWhPs0rUieBb6PU/GH
NwpAqXvVYTdIsZTyNaJDQ5Px23D4cOQaMnK5ak4G9FsA9efqdwcuuVNqUZ2k+zEr7sXFsK99H4YI
ZFfM1ZVGfVwThwhFk8XC9ZsXsh++npVma5uKncKD4kudCb0j7D+TiHulQHP2VZlDU8NDmUUJXJ8F
/LPMqPB2e7Ji0iaF010umdzVhvsD27yDUE4uoSporUKHsEHvpbRKWFfS+QXAvhWY4NQ3lcH1QD4/
1WzyQrA3q+jFPrVD8EiVCOhI51Obd8U++2axZopENvKtSmg5oSzgKLfxlyFV/XWphKPLvlQlboMY
+I0l0XXQhqE10GzQtCvTMhqG8v/YCA58dTld19CFZsmO14LpuAg24SAxj2r6prXXkhoef3iYxkuG
yraeP1B9YMRLa3QT/GqelMXz0C/yEE9C79UaY0LZ9+Ns4V1qjTpzHmkbVx6Yd7lMhUCu8DWucjeB
ovqC1+S05d4VsrTaPiZETHnF2U+qUS4M4xAFkxPG8ocP2uf25j+5aMxH3cQ+MBQrglrqDIueuySj
yKfnW2lukB8dsY6YAV2pFp6mwG3ki3urs4PYvZtp0DSqsCP1LvcSIxuVo5zZ+gcfnXk2LMh4Z89a
cnJsnaVgG6qRG+M1xkSTnlBXOffZ+O26t4m2zVOo0fq0GzvWcO0TBRi4jE3jZsoCQEYSXPb7oJnY
2twd+r81wywbWkYvX5JGJ9idIHbp+EgX8Q8yTHsCFlkt+b/xapNeeYyHWwN6o/6dNIqwH6OSoW2R
rbBZuAZGVPXJbsoWnqhIRm9WyG7KVuKUYkIqjJmMKFTqNaawsjQ5m5LgwWS83CPGATBr+bwrC38z
KvCeROBmp9tsCm61jxXq6syzaWb2UDC9VZxCtfbd3aWTIeUVa2ROIa8xUFmx6MVBEVniGOwso4Gn
HmkO5biIeiQs9mGFr97bJmuMO02azjKN6qPtemVWMQW9azuvmo+6ShY5rbqIFQvuwZpB98YpNejo
NweFw2OiMfi4sJ+Md5iCPVuCbirKdS6pliy24MnHuYlCYd9KtUKVsNOeLgNSlIDU813hF1GLJUZA
C5IVlZ/WoBW69TSI1vizMPABQe3ZPd0KEL9n1i8ezfksLcZHK/41qWDDC7VyWG315Fx1/vVtxEXn
uezT9Ir9AMu0U91kDdMhPIwymHkkB78EfZpCapQE5mCj/ztgXix4Py8WsWdbXKX1g/2uh0AJ7cZh
Zj9Xd7B0mBjeoXXumVQ0yYl5JXQKK/gxetiLtBQdWYNA0DXvfqLqBINzy4hL2DJCaXqFPrL9gDU0
Ixb2APLOhVC1eB3bZ1RGOsa2v3Cw1MbK5BckBB8OCpfGBaUuRJbdp71NTQ2sEH1IAnix1vKintJ+
EAB6tnzPdvLzgGEHxZq27e3MowFTaKcOwWEWfA5IK13XWe1DUZgsb8tIkT71osoATEnO2zqBgPV0
pK1IAxtuPvUg51zFoSxCtptIne9DRBF4z8RzNnnzQVSop8c0wU4ctkKRJ4lCV82t4kd8Edl8lt4s
zVeA3yhC08DbYgqUIUScLkyWl73/cGibNHx4fmEzD3OcxIWQmMD3Ptppnz+npnb0L/ojCjFbEkAZ
w47Zph+p1l3FIny/M+kmuZMvNwoLONxfg3yOunNFZ2GfSzIX9qazNheQfjUApatjstMEDLO45gdU
uYHERmKRrmVR5tpQJTTQ6DDUlOd0fzfUef6qh4Z1xocOVU8ZlQthy6cKHzaABIRdnLnBqdoclABi
oJk3n218ZwfoFLSBkgL69XE2N/ggkwc7Lw9ccHJdcaibdKqIBdnQV6s3AFQbYwsX5IJj/ltdlpYl
SQePUNKScxTg1T30MRE3eeOpfJB6llGXoe8CG3GSar/GKmu+ZoLKmI1Axj67RkODH9pYaAb+B0aQ
7H3V2JuM/Y8sbqKpeRXo6we60MZz9LhEERtg0b5HHXTavTnH0l++ek7mTYhzNn2okN9ODs03Z3xD
WVdvKLA1kNa1UN3a8ufeXdwiQB1TPqnfK+6uyQWtpWIUJyM3bEgMYAFIQQAQmyE9rcCq7BDonTS4
OWsgr5pR3DxjQTqVKLk00TGE0m+76Y73c4YeZzk1yk8SheXBj5TlhXIzHMQYz7/JjB+6V3KxpUud
+zVeKgo3G4Zww7LhKJUhYEKHu4OtjKAqi6y4Tk9dDeg0P8tGhoSMiNc68KL7p6IPxmqLYuEDs/Ia
pzsstln6C8XCRrQ8yE+YwZxch7pB+Az+pDnLOcCRUARpMrrdhZThk13/Jcm2oxqvEcYCJ6LCFpAH
mcZvUHBKKmshxp/PSsIZb7DA+YbxhwdCcCjhpOUWcK7uBbXTPkfASKTRZCgSn4grtkEkcHt53J5n
Qrk7gPYf3eOAbqtNws0kxi2c2u/vejAlZebbs/a8ckTn4Yc3a5ejiTFPqLi29acimK4eK19En3PZ
ASIrL0pE5b1DEcaSuR8DN84iQ4+2D/nU6zeInYKmXKjF8rxbkLhQXmP0jS8KD4KsnfYvSXYxkawk
0fGq/8sZdre2ni7Yr64zH5FLLiEZ686yUGj4apbYOE5LfzH04lijArqSnHKe9Qw3JAKvnMypokWX
Yuet2VD3IhE0iRbRz0UuhAutdjFq8Qe9skyuUpQdr9sxQuatAZWCaeWFRNU6T6Sc5VSWz/VUINXx
SA6P34nnpMFgTzEydRGlbHLmKXfNHjPg7hOMwxbZ8zDlz//7iED28pq8ZjIYKqk/ni8hZlRtAEoE
4Vh5TKU4+LmsDqt/Z43xgLT3FCJ3aIi5DP4nja2pFjkqPLFjyZvhX2jDN91HQaSvyMS1QfIHwuTu
lW2spNUghz0OPdd8KTSmh8v9r8Y/bIBqfDwsS1UDSXmhl/xptouikriTb3nzmp/HJSkGBogjMCUn
SqeQI5zoMEWxmgD2sgQWjPPlcZ0IRehSM+iiKpiisTRLmQ0Y8MziD0VCrnOLLREk5/bvixijfFA/
mHNjbjrAGG6Rx+GfsxhczyrXeNZChDp3uiRrVSSgIJYmwUpxWfMH9J97JqVfVVdVeXk6miabmGMx
dHculNZmwvXf2AQ71KV+mJFyBlU/NdJAhBIjrLwAHILsjq8tjkJRzWLRVaf6zD9AcreVYc1hkkCG
wu9ZJuNyLX7hPN+Qs9nEsw3yp7rSVBR6xOv4/M3dcY1U5tBjk62wpovP4IrB7Es1JK4RQHwSjqlm
ZKncSCMWhGDm6Bm874oOTNS1py3i56g8Eosc8Gxqp19eBHna/RClVdgKlYIMuV1gqVU6ycgVM1Bo
HjPgQrRTggiAk3Gm0Mc2Pn/r62AQfnCl3ZSo96BG15symoWpNtlhfsA10909i1BIUsAWnVvVh68w
wh/BqOk+97uGbU69UEJ7zle0gekjsy9312G1fhir28h5Gt+0pjtlY7jcwLpRVPrTHXe4YxXHjqQu
UPJg+5AQWt13sFTv36mb6m76P9tJjGHbYaQBX/oUbCG0+7LN3XWM0jEP5RYBzLLXBtAB35xW2vWl
5EFVaJCMM/3+md6uZTB0iG+8aeL1K45vzt3ZV4GNCb74TKe1ahlgFqR01LrNg2jD/oc1Ze6lyc+P
S1lv6i8RQLjgkQXxyE9x2TqMiEAKCipI1u0ulDyTSzbh8355WIVdOW5QMWEvCRnEp2dFCn9JP19L
zV5zkp12v+RUif3F6J2FZrS0bHSTsN9ZvISHdWcscM5L24MwjkiIowZB/ZNCUeDSxvIH4a/zxc/j
O+0PbAXtNF9sMZcW5DLbqs0VIJ6rluSo2X+8Yq+bnH9M3ZrM6Q5gcqWU0BpANflKeWO3MfWWk+l3
w8iC/3OYxYLZiQE5PNpoBMA5rrSCITmNsBx5rqqzLY3/BwTiU+3aNsnkXyacUhV57vzQRMf7IwRC
3g4+F7xW1vzaVuL6nlbMWg4dW5nT31jGJ88GOL0hi/ytQaduQallmdrWJRzgdAlyEb3bv9puEGPs
gaCrYSI58DvdBdHbp5ckEVLGO2tIC/7SprzFmW97YKtkr72euZjX5vYsAD/JIJLeSsrLxEc7Jm5k
kOUAGFYYoXOoO3rHYf2Sad0/Kl0HQQQIChF5mTYa0KEwsaPQpimRbaGxW+0GCLfn6y08enRS4nk/
cMkcpM7WqI+OK74+lO83vwWXsdYVfIEXM33nv6vGYPRp2M54FbkAyAT46hIbgMtqhrBJ6QSSHoG0
ecRr1Ue9ScRKFRhLQyCySBdoyey1N/+8+3cuSznE0OjY4aShRYaw8Ovm4LoJ/MuMNs01gdOCleM/
+bU5PbaQFF8/IE+sXO7s1J3GU5JcqGUqMrjVmR6OGWHOG2WvtUFMNa3imDmoH9JbwAc3EAzQVKZ1
flmmTrURzPDrf/3MiSLb2085uZYJBw4Y4bqvt+OxcBpMJNx0L0OgTZpC4r8kDYh0rZfaC04bys3v
sZrdt6PcA3cX9+u3YjRkNQ+XW/cOYcbvoVmRB5aeZVCGkyWkOn8rdD5cWABRz4o3GnAfubjX8xji
xTIRY+rwPj+F3bHkOEAUEe7zr1BT3ST5yn9b48UaUEnjAwyW8vGr6xnoD5xlK3ShNuTFE85efhVl
wTSRHnAk9fNKbNwu0ubNFI1Sun2v4vYEtw7xBrH2RVhc8YGQBymZ0y/jqXixXa2PGx2YN4rAO3p8
av8paOAg7cUQJlPS7DpSc+LiJaFsFNH3fIv2vvca9L+apOVhWrMxFWysj4mVkfwnOZ9e8qMGhcej
wAyAUqYhro13+n1zYJy2T7D36VyT04AACkuFIG6XqLQw6jJenxgrTPx0mKQK2B2r5sLmj5j+D3b2
7u/FuXqeSnVWMJh86HAmQh+IhdTjsynBMnFu7e4AUxjb9qtdeIq+HXMj5kbiT+k+areqHOqwYmMV
nZC+UPn9TlcDU0iTFYMBLmLPi7BHV9n8zR+a7deGN1RAzoqz5mjR+0JWSKUs9i6AGUMzzKv3h7gU
c1dv5hm7pIsBl7+WCAYObGiioIDbGUMUg7QkvvayHt0lFnSaCZXEdSsI2KKJJIs97DtBtIIbcIBN
ZKpS1xNPFtOBOHWpxZ5Zg2zmP/Rr08rc0TVCYTCMp7ongw3t+HyQUlirom0eQQjlD+0UDvz1YVdH
F8Pf8DeSX/xQDUc+Ray+2Yj0ra1IDKov2LFd65QTY77PCnjOi4Uuekb/yB6e1Desdl62njxiBpdV
vcz+HLVZuZ7KwTEvlMbiz4p80oSV6/JJe5Jigx+D/TLNQSWEkCF0Emc7GnoBOnFte11iDuE9v9Vc
z78+IDot9nGD8Secm7sIgEf/I/n0chyOwKhn6NFlLKncRCq63+fnTIzSPKCY8hn7f5Idia+IjtbL
x4MTqVL5olk3c2oS0r46tlUt995j++WZCkvHTHlTWdZLwfhJs5Ut2SB2dbfAFGo+TpqGPediR75z
wISywPXsnvhhEjM1RhUPMQn6naVfHtli91tGXfVgdxUg8eOl0k5wKZGdBdf+4GcEPdOTlLIJhl8H
L+voGAgel7y6D6g0Oi/tEKvqbNBFvCsWl8Ca0JaWGCk90JxjjVU7rSXsYeJKDXjVed5AV/t+bzKZ
QcPPJGoQiwyqnOnz8EialyIJn+opfwouH90Q+nJ+ZKMKyYL1McQyESgxB9LUmBSdChJKKIIubrXo
CKruvOHFJtGIjA4nF4cJvTiaDjJmWfkIRSIiauAehQ5IMaUC0qMITVqLc5ZycWzCamTC8WtjxM15
oYYVhMkhnCej4mU8PYvtY+64DYxz7ZNYnrVtTE9bTYF64r/YVuJ5pLI1pDmJsJ74qB8JdgoyQcQ1
8z9EkcXfd1OnNNn15UbffS5ZdMOPK9umku+fI0BHtvJxGvO7GxSWSLvoNjTi6J7TT/CB4QvcprFS
Ax+0hOQIT1i0JVpgOiY+PJNxvJoLi1X5TLVppxcCXpsSxSZqBVAZD8gZKGvfvLpiqrfJMh9jyB5h
lUD9veH9TUXr8sb/tHTJ8biQ4Md2S+T8PqlNdYwAZVTil9qvzZALzenOfp1iQvWlyVyY+29N1+ib
J9Chouh0NaJlPKNKzv9aZARcGXSGD3PHd1iQHdTTigsZlspdXdbNQGog34i1ulwWT0KjajcU0nU+
4v2j53Fsm9a6aXZ8BjFs9k6k7sm3gKukMBgT3rIbNV3DunMfoDt2SS+XdcVLaT2ldKS3GZzAnopR
WQraxdLlpGj7WVhiS49SzpXHMLF7Cct6FtOPb7BsLu1XOinciD0S2R403n0b82t5YRcNN5YWbhaf
f5pbVnB6HY6yUGkigu1UBexyrnvziZ1bUGzCuFzoHX+SRutcfTQm4BvbMK8EGCFcct+PmLo1j5IN
kx5jut7gWZCNj8u0OunKcoPzbiGp7Xzxs0KRPMKW+UG4sYjdkgB9jKU8eXW66xYjQCdqeGtQj1gp
mQPs5GPj12Hl+KoVonlvmge2SIQODsRVqzGY9Xvg0IMZJd1+jbBK2If+InB25kmsFGfcCGgf5+F6
GLHj+5Y8Emtrnpp9L/vHp4LfeXCjc/ajfe8WHmyxNma+HeBDT72RpbEo5ymIXH1rOBSrzCPoQup6
JEAvxpzIUhNgTUmmrDobOcA1QH1SkZTg6BtsKBxmzDrXgFbhQKiYdydzKMpFRpDndbiYw7UWIPRs
WQtixbQ7SnkPJjn2Qfh4VDvCq1geSeKB5V8cq93JfdKuZN7XULHKl2eY9jWl1mxJ4tpFjBYTomrT
XHjtdsHWYXGg1oFIiX4dJOhFdJi924X5jSJNdNrRdORMWqozR23uMxotY9O3cI7fA50q3CamnSfm
FguxCBCXoW2+67uMCPVV1XqpBX6MQQlVGpqGd1Wz5xyCY/OnIynH3BeyX5nEjvNusZWD8yUYpKaH
3J6WMAEmRpxY5Zt6lU2dc215EAgugSA36Ac8RbevYTq6XaAFF7kfH+i+ZZpBtVg92dY4CiY19LG0
6GSbq3XjWhVa4/V69sbCEolfC+UOjrfiwuUJ32dPOHbFadAde2eeSqjXttKbYxtL6DI3XJFM6SFo
DQd7Bg2uCq5ts184SXiltHWxDPu/WpMsyibnV9ylNW3uL7XRbgGIt6DMx/guRpTbJ11YUnQORsVp
DrOgewFnBhPe75jiWAZ2Wsc+6YFibGJ1fjBd/dgNrgWGAOYujL/NwyVO/uU5U8s6wrutkfZaMy6T
W8mRCuQF0OsF/aYKJU1CgRhHwxBY15S4WtG/qg2u/bY9nmdtrRq3K56dnWZTtndUw3MgrQEh3bNx
KWc2j3T2xu59uVOgMID3rnTc6PHQYcG4NQa6szdrh27EH7q57loBpRB1hcBTayMjQjzfIqy0/qeT
HJ+MTGhacJv4GpHT+8RhQmtvF2EkDdBarMps7Swuvij/qX3bR9tku/o1XkeB8004gXGdK+wBs7Fm
bnCKVg7e1wTNAR/h85vpibY6ACYOqfdy+UC5IV0KnkzjQVpsS3QBVBZPz3tv3LASeRwjpB23kXXu
JjqNPnQDymkipm/x80S/L8D4Xr+JSJiQn4y8Rc1vMpznAoCbB25jhraL8VJUgTs0c+JhtpRb3SOH
4raR93HiwYcfzo1QQB+UO5kUEj4bAUd/vBa0ZGD4m+D1dbZnWy2TTkzzrSpM/O2hq9rh5BKKCORq
DPETytaZodw1/sN2as+uMq/ezhBUW0qy6ebp4An1kM+SVb9BAeBFoOahbArlo+xjmhsl5LypMwwi
oGlgy60EvUGTrCUD1pql8OcXGVmEXzP+Mj45abSjlM9R1oHgrD28WrxWC2Egbp95qOouZ1AGnjBi
EL/KXk6/7BvTYQzFV0i6Hk3UuetIBtxQOmxjaHx2At8QAANOnW3teK8svdcDuge6ek65gae+d1q9
0UBWQHflyXqv9P4+l1MEKhiW4ql2oXnOBJqwK/YAttFt1wK/Cp3slOf0/gjkslsazDIcRvF6FNeq
xxLDZZblAWa1H41b99HOvZHkX+uGCpdxx9DJ9JTPD71nwZytFZoXKn1N0hqMGcxqodIrWI3LVNJv
KC2sHa7iYpbdBaU3KDgFUnnDVf0OHfz37Hq9H2r7IvcIMXxCySXW8RZQCxenBT3IQMEdAJNJTF0q
6PLxDnb1BvMejSEalraEbUmzm8764KCCxNMM1YGyvhKXjW8nMnrc/F1nWQIp6xJKTh/HClGha8Zt
iJZ3f2Xe98iLHtKXkh8s32FEOH/yP7icOjxKxwgH0IyhAAgDBldexuc+vv97d+9XvKhCAh140wrM
uy9D3vF7IutqMwClEi3k5vEir4vs5/chZBWF1ejDBNCxQCPoGcddIA98VZXW0TkbLyIpRPEIkobZ
khYaMzWu4gO7++HnMKwIjwXDEwKWsJM8A6vGG3Rp/A1iwRj8sdtnZS6J/eLPVXRE+Bll9kKewnLE
QQfoYGtAl+Sb2UTEREUWWgN7HNTfCaHHFyPjRiZJ4UASv9jzV5DRaAGbc1FCc46BSLkUJCdUJrRA
DaJY6H/sIRxEJpgqn2xlciOG5l+TEwug2RQRL2wsiLRucipiCfi8qoDLAuDpDZKjmQNMpaiksZGN
ozZOCZtKzGqNFhZhc12tMnlXxg9dK0SM7CEf132ZC8WKwOPk4PcZxzKMKlBGszjsUC2ZPtjfHe6R
FGhLHZdLvwfMUxlCjn+AMd0xv53h8ABmuPNJ4tn+UabTTh3I09sd4L5bFly9lLZrvbdCOjz9Dj1n
LxJ+k4ZeE26jKbZQQX5bdaKGPs836guBb5b7NjKnXyjMXO3JI7PmDGkLXmH7qeiY4Yf2St2fL39i
K2/t8tOc5fytrjLEpy8yeqLX5mo7AKy9pVPNfAcKAIuT42DYnjqnpPDqIM8haK2fECZu9BvyEVZB
QpOlFSEh/CPUdYy65x5ywh92b5BFUd2Fo4DQKLAhYBxJhbi/MSiLRmeJZfNEyz2Wk2v9B8q6lijS
W4//3mQeBbWTmZ/381jPqhx838/o1Xu5OgTsfLmUNivOtOpZR/4E5yi/QiL3bzvqhOOeXMXxCzrP
W5CHJwRbCfbpMPsfBlaNR++F9ZbyTr0OfjHDNhjvd5ySPkoMQowYuajWIH2638tkV0sY/VGayFfY
v4wLUgy8A/x5+mz7SCYWFJBU4ufMv3D79QqRPYXuaQMUTjAf6Z9+RXbaJX1ac8O3jCtMqoQVx6E1
Re/qieHUcxR/TVFdnw3eFtnjNJHNk3M2L0VdRHwkBSYWLzpMonM8BmrpcKpTcN1AsbZADuROhPQr
cBSevf6m9uLeQD5AycvoP2h58BBSIMa2Ic/tb2UZ2KnF27+BirQ5ANlbt5dZwIecp+HsOUWqarjE
/BvhcuP7EVz+h4d/VGhAUr1oOSivPqJdPAns0JzTAFdHxdJocGJc1OtIO2VkHD/9FCNu6a5+p2Ah
RySK/mauCYCF5C75GxVwEaygAQeNgXBl0XTEyhuQu8kjw4CFzhrqTqwP3xfXYv5979EKsZZ1tZw0
gYZIT4AbjQHTZxyfbxa/7+QrbW1TupfkIi60m/JI8JwppXn9GAaJJ1LTuS58y98onJYDpQvyAu8e
BzqIJvaT/0dHq1bDEhFrURwCvtwW2cuPE7qa8YKiLJcAjrnsCiaR/g0LKu8dANVZRxDwFp2KlzY1
RKP6+ddp7YIX/N5U72rS96OOqtBx4QKpsxYT4SISP21q/ExmQk17n+0Lj4SQHcXCDzdjSdzQ4lzN
gqB0bmjVzvdosvjpg7EcV8Xdv68ifUQLZsUBBs9gizkjdg20oQwStxKij/DV1vuOodvWGgEQXIvr
Pcvlyt4HU9d8B2OMp6hKomo/NOMv0+IO3sUd7w3jBEwli4odp8R5z+PTas4fQlojmAEuW4zFCAkC
VDWtdBqhtzpy9xvzN8rBOEYdCrCYsLhJMA2VPQxS7jasPtnlwpXfrYtPGOEsf9sExdyqs8mnlgMT
r48y5uM5Y1dwfQCuxqakMRVreXDs2b3i6n4DEK7+c74Z4xYRUCIJoRHoOgWWsDHGRWnLnuqMwVQQ
YYQwX1od2ciNSSWPG0AmMsBRRwB4NO9VD+h0i34WCb0mTP5HfVnLqVLhOCwwMuLaa+M/BE9w2lNP
ApgvoDIj8mfMlVZWfAsJS5LbSADC2BgsEJBmOXVaSQ6qAF5IlxKLboQZtriEjYhpWjcKKi+2VGyj
gtKxHs5Cu5f6JZe0mg0X7/DS4Ksaa9uhrbml/3Tqa42dJIWNB9wLCInkNz7YXCDr4cZx3T4X8JTQ
189jHm4FfuhzonO+W1TdFS4nzQ6VhYbo2PJEz60zM5hofJHMgFKXicW+at/r4IuYtMV0ffn0797G
+EyzqFl+nOJqmscwbIGHCBNGw0Pa2LVZLM6vd+1eOp7XirZbzL5bUT6g/EJ/6gA1xIskqQMC3c7X
WL3aqOzH4LY28mESatrJZre6G34xdH6a60jhRTcGAfVzUYoeNwhyH9buAIVbdgBLjWgNG1IkR+A8
Q/WG6H4r6pGuBrM009b+CSzJyHXkA1cn8mtOprv1ZjeSoEavaBxJRLrEo7G2bWhRgtF5koc4zN38
KhARlFy0zBZ6wwbVSkZNoAvD+9BCj3R6sY7huRQX7R/u2TCXYJgMpnAtwQg1X0mGRubljC1G3B3d
YbzgqfB46ih06QemgMeqDkGtgzk6Tz0kjtgBnaPA/UhWmvEJMXz+PO4KZEKcXliHiQtlyEdXqiHQ
NNF2HKqfrTRRfmssSAmn2qmIgFNq9SfBZ1axOOAOAl57hywiiN27/6sDR5CGi9bq+Po7w6JNXIeS
vBM9WvwOuY7imqoGieq7YLNTqh8ruolk8pLxp96GZcPgsbTyaRR0fc3CQQehrkbdMs5DnYgeNCiF
gMGbbyrg1+ElkDjZmixQenv0v7/quHMPdfs8/GMpu9DEP0KNyZq8MMUQhIqa/qNOJRnOz6l2E/B3
50YF/t0gT7S9P4bmcNpvJwywM6t3PWFf95+jmCqrje8bq3y2vrISE1324xX35mYX5v++w49PUvgr
kA0DImXQB0HJhlGygrmP7c16ToGUTkQGEmQ10SM9jjGHleUfSpHxG7LIa4d4XbJDVA8WogI5gMvt
1cYk0FPLzNh5bnhyGqfLJCTeydvTR7Gzv3pk19XmsIDC8oez31UTJPuG/9qCka6feCRpStouNvOX
bMrOCRJPyl8Vl9fQdqCm63ZwrI4VHwyfYQlkIWmaHBRlZTFpwvNbYwPZWP+LTrsNeUOJZrgYFJnL
Y0+VvQPo9BVgWDXKeyIcUQiMIeQmT1vrF0VjuGSMl/IuVshTmas0OrU8gwWi834zGI+ujSjlgtLo
Lg0JFwA6yFQiXEVQXrNTNQjK7FSX249uPJVFSCsJ7d1uqBhBsGVjNivaxpgt52kbdPZ0pJ1dnFMi
bKo4qLuUd7X0XvBnrSGlIefAeAlphM3bRs/hWufG985qXmqGv/DRSrajSyZlrdCr97TKs4u4s72j
gEf14qP1NTYjrcuWtacd+TwAuNZe91+ryk3VGXirlTB6Qycuy764kF3/OPspSnM6Jcp9AGvJUr3k
XPOhRhs8BGuJ2umwGtv1887B9S3KoHao0uy3Aq3ywu3OjFsdLTYSqPc3J1FsviH084dtDsQuy/jF
TL9+nG2vXGBggKCfnshBYhH/u5d44eWoNmt4RFzN9GDwWxFVGX3QPO6JelGoTBcJT8sYBQXacn1I
gYRcmKpLBGskrovwx3/uROkoRPWEMDhDpfjhHT4bujj1VPYicuaAp0QwU+i5flwphaqstqAwm62L
qFQzxa4/MGeBpV98VIypL659QyBYwSKi2GCPdsY872LxZaPKNbb3KoCNT6h7mdvAHdCHPuSuBK7Q
h3YNQQEx6RSmxNeRdg69Mk9vP8yVsdHkfhO7Ey5UOxnyJXZCt44TbQgZeo+S4tofjiEAb5qen7RC
yq6w2UCpAYP72GlikD5y5xchAFh+z+VTWzv21Ne2Lf3X0Uj2XeL5PgLqQytAnj+LHwAILVmK6BHG
7riR2VwpR+gR9+YyKJOJXP6GPmg5j4G+Zjfj6GTrbmfx2cp3wVuUtsVbTnhGFdDBWNFokxTZEcSR
tDVI3OD5jTlZV+566gd0WxJSjiXV26CWDuwHDPx25SD/tX4WCpJWRHNli3X1RpHsi07psPgfa8aY
8j82+MmSNHZU6641/W3672l2xKl+1O5S9u9FIf/LoEC+aau9TTlltWmsBD5ZyTSF6zCsBO2AhdS5
nD/QxmwIFugSCb0z23mXaMt0tw//vLIaGx+1Dzss6si/7v7MWv0K5y5WWJd8kGkyfpUtwTotGxLL
G3fAHsOMAz8iRvzYpPJsT32N4ayNeKgMAFW/Loauguz1Am7fuA75CPePveDyk8wB1CKJ87AeApGD
Hke7awYzqmTGk0nKDOX6WmA2TldYphFUmPs0aJWeo0Q3tojQP6femHyK75PC6PgbUK6bvnGaINiE
5GJl/yodD7Xhomcqroew0KedKGHr4/EtqaOpVyIli0ItzsVY/MWLHTuGwWYFkyp5YMkCT/c6I7zf
XcFEmUWuEY3zp0u3LQfK/Q7HwO6dtmGHpuaqU2PfTsZrWtL9ltekZ72ATIkLfqYLLrw5FdsQyrBa
VDGSr57Gi0xtbN1eXsq0o5EFeW0h332U8vqAQZ34bwFT5tUpY317RW0oCPPkoJfKPw2tqpTnu4Cl
6fIlIXDkhRf7eNXhVrG1TVyLbO4u3UQ5shBeFJqCxZq9xVA/SxJYTAYqKTfzY+Y3YGE2ZpIi9K2V
tS4XWzM4IgWRCWrJ5thAArdojYhEfcYb7tmd8t7doF1RZOPeAo2t49BxikCACROJTEjdC3qjBST3
VgTUxnek8IFOWm4brPv41niYuvxxLiOHASFirxeHDvv0BIaId//bbNN27p3WwXWrgVG18RNVZ1Xn
tf3h1RDGvt3OwWRi79hPb0ykqyNSn83RaJDH+uPMpDVDCwugl8+VJlwsBpwOud9pPFDNqmPkBiaO
YPMhzrTqE54WriA+i69X9ljzfa5PRfZupt095jPijsD5fMB6FbN0DmJ7oWVqbbQoDuSXpOiKfJNF
XqGVX/8BdnuGJp0AVu6DI0foaAyURHxQ8sz97z7j0MQ+1RBrSMdpK/o4EPXkHXH/TeWJ12RrGO0G
ad2hddh1+6RjKrcx0r06kPqwx4xVi6ikjSf8kqKugoBPEciBIn/5QrkjoGXgMCBc4ttFk7pBD4KR
3DHaQ3b0JRsYjs9tqnvlYmKBuuhDxiThGupQVz7Wlk71NLRQ3b+J3nFQEG98UQ1Q1y5zXMjC+uhm
E45juUosGrj8W+EPeoBWdaTw/1FAsFtYAzuTQVuVmP53+5Tp0jYGoj7+pKIajIF7/IgdZWkswAgs
fGV9AQ66Y4owZ3qQoM7PFdi88aPtxX9QxKYEYsRKdUrkcCDbSYw0fNBkJPCIhv98nkjhHZDryG06
rf26WEFWQXVFfw/wu+I9oEdWvk5l11Fq/kV7LP/3v4XdZPpIgASc0qolnca8E608wBgs+MjA0HF2
gW8DdNGkqY7bVLra4d2Z3arWF8tt6D2I/uFJMBvWzSZ79kwTB6svrSXDzXZ7XdhQ7RsQamM8Yo1N
j/Lflf7FdVEfYYtMij1luaWBY3zsho7ODn5Ve6C2wP9XGZH8QYIehERTIFgSL7I15dU/S+wLY2Ua
bSt2iZxUp+H5bkj7iXiXPCnbsICVTF5sI4DDCMVtRdHqvTJxNtL6k5Swh5J9zkNAM4WPKkdao3Zv
WYWoR+SbjrVzI0qZmbnnZPyKAvFU3xirJPp5rbhjFD5oYUFcNurk5JKKc8gRe13aCF880TP9uuG+
9JXERUxSGnXHMRog6HfK/0EcMx9R8pK89etBlm9a9DHLrL998XisGvKBRyphJ1f0I/DOdRcAhPcZ
BU5CR+RK1ELenJ3Sk9tn+6fger6gZLAKQWVl2bDNEe5Kz2IJJ+kuxzvy37/9Tu0EkmzMZustiUwS
BHJDkT90yhk/wWaOKsiZpoEifXxRmI99uCpm5NcHZEGv1cdwtlelWBdtMet26gjBjlZCmiOirctg
vt/euoBPA3pPxMislTg+YRMWR4kSBKpDGQOn7OYxVHMHVFnRCagx37Q6NEahAp/r197zlIJEcda2
v96fqeKl5ElwEr6NhH1C5qE3Hu0x8mglmw9lGuA6r5xxDHmYJPY8EK1a/+eryKbbsrp4rCcnPiX2
G2X5bRsvg5EIlD9E3HEChe1h9v0g8NEcpvleC8wEEN45LHmnd+QuMZ0qHNBYTF8Ss+qoloo6fyIC
xezuQT30cVIeNa4HNGMiytwEz2+rIGGMRFQm9Bns3OJ2Hhy3KtUCnp/bUEvrgYAOSFsFo8DGnW0w
WRgurI58InZytXheCGxqM7QZ9rM6r52yzfaM4LGkk4sAa08suXxeXLEQ2zK5biV3KQ4D5yTmUZbe
jbersPhcHh6lOXszDrJ+nf7UH259iX89mT1SlJE07WLP/UCduWCeEfEAjQKQAr/cTTS7AgjtblxK
fjxi6PgPvKt2HBc3GOGFJZ8ZQeC34cwgNzYxOTU82D5Vh0eQj3UzXd6nyUnNgwDqhXk6QWNl0he5
9wuro01hXcpLT0ZARjLT3EevEpqgx5giS1HmT3r2lxqc0fC3wjv6eZDOQlmmDEpMTFUp0f+wYIr1
fWzvNUHTV/puSMatc3883PfLYQtgIgiIEeBXLdXOgki6M2CnbLJZYPR830IVu4mv+R5kh8ro2kW3
9fFqiRUWffdOqmlW7Vm61O9BidefjF52FT6YU+Y8A7KuPH5Y5cSft0qJG+o+PwPE4NFhtnirU577
8ZqkK9YcN3ID7i6hMfU2zWzbS+6EKwNKyZZBngdE2VmhWSGxP5Xfu77tjdvVt2I2Kwr0xk5tdNdV
XPFzM6ADWyzou/MjHbQcZJzJ1OQJRY80H2Um7WMUXerCsTBQ6tg+BYDkfS/dfhWPYPvTrx6jtVz/
GKzkPX8lqtIFQvoUn1lG+sooELcvWVdW48hIfXyWNVcJ4O8EGOtjoFuXqtu5IAgpLhHKRNDluBK2
vkYvqYgrDcEgcQ1rSGmJFy+o1NPQrx2xAYsRG7T/rcCLwDZ+YOONkA9/YVzO0DMyZOuojTD4gxV5
3M33nyOVvxVQmi8uu2fnIF/bNw6j910XEh1c3Iy5zULbtS4PfNgh3ixL5vdTLyB3//wdyDYcIjhK
Tw54HC/EXJhbVFEEiLgZR+x8rLtfm/w9v8uR+Z0loE2qgFuLud0Go+l4/Mk6udgWT5Dl/nLPPlYp
NH4wPcpb1ZHifbb9cHURlP9VdjKXD+LP4ktZ38RfmYkJflYrSWZiTqByrbs7W38T/4E/nSggE1Q3
yeZYbHIS1pKvcvRj6kVt13cokoIu17VTvtFp+y2NMmyxnV5Lv/J+OH6oNI90XLfFggIBlr2BoiWw
CgUig36NG0Sg2zrqnLh7wrPBmtxgObqtRx4XdFJWYSKxb9HLIQylkvzU3Jv712ZqL5oToOeF3p1g
8S0L79TwEiFByIDwMC2uQRI4ZhqwpnKqVH2XueC/hn+4/pr09RNBl8661wpwy2F5IKPq1k229lCx
CUGQ0UiCMlmnL1EUGec0wJmateg9ffwh81cITUpvGaOUZMDY/iPj4UpBN2XcFxJp7knC5BP7ElwT
o9Sg+efz96zHI6fqFKf6wCk5XCHT9LfKVyKDp5xxBEQSxpIk4hR2pm6frvb/GNwF3Td1TuAe2JYp
9Y+JCpZexYSL8/favmp71CegTvZUeo/XZ66O4p3gu79VwiXlSYdSr3oEfRhY6gofTd7qHOoqBlny
frI+pWPIdAyY2dGCpDZpzRVpVIT/kWqi9KaVHGNOyy4EaNsUSFWpHv0CMEg1bGlhXJggFfkHZeTD
SoyU1Ww0D9YNKswCYS7IayXGGuFnL6sA7qDvpgBaK2XebXhzO2ssQd2mHQRvrlFxecZvMUQjBLTv
y6dIN9zjHXtq3EHn00neiFhJ94X/+rUBpVq8qJBjXOilcC3yw5pnfq07bWvrpqAiOgp7m/PHaKeo
GlNL5TpFOEqwd/aCNzb16VxaHMjofrgb/nHVOfkY59BbnKl8r6GXSu49P8qmhR4yDebLeJyEf46H
tw5Of9fmeVbz2EMMo2L6BBwaIzXFmD3DF2z7m7V//woJxui20cW9+qsfWUDBLW82/Mg6j8m2Qtmr
SSguqALpvQwIKeyYrF6YHsC6Tig0r6BJcGsrErr8/sWhNZLEDiQJ1tUhc+UirQsob36GhhjeMhSV
EoCwOvmLKq919RNbBA0GEzzwgVPKil0WJ68EdeqV8za/4xJzhZSxnNApwIweU1G+1bFwnvAS3nEz
0Ma3KKQ5LVG0rEvxCyjpBTEKinmZCx4k6zfefrEnnwveO45hv4SCHYW5ZGWL5UFiQlJcEE2izFZo
TXnW5CgGzy1mbxxl+BLof4gC25NSCziH0ix9C66VQKqPPxBTF2Kdf2V8U6h/VFSywoLJtrge0vTB
1wjwN+3qXMGtRNQWmOtMmatmq71G3dcyBa5gdYzaNUgNFpss1BztZ3KKR4tBCfT7gApUTxUxt5Cw
nlNFbzPxcyfqOu6s7dHySIyd3OKSb/zoygLzTJ+VYYNugthwQiOUYJsTer66QNSMmui7mf3xLG4H
E5jMd8ycM617vegYZjgKGXcCqVwelnUoIUJPbsa8cZga3Y2ULYvsDftRfrASI7Wzz4wGgRSk3LeG
oJs2bv/69A5BrH42kjw03TTzNeUmIdwHdbe1TPP2SkyI1s41/5zD88d96NLdZSysGR7NNpOEh1HJ
7XswhGhrpbXK/snOdrCiHPALKKGpcc/W7Y5UHIrCA9/GOfCJDLX0+OOhM6NukATh4bPlpFPENmIx
yegZnSmvJkeL84/3h8dUXz+pqd91oEZoLM0MlmarPQGx2M0uinKxZWpOBtoKdm3Naq7/AERE2Sv3
PgKo0WinSDNZU89ltd3uAnRMGELnoaE4UbtXUXQe2O6tvSwJ3ezacRb9PVEsRxRMR3eJbKei8cQt
i7tweSAhBWQKLFztQkMgAGzQTLZ9xAAu7nX3EQLCWp0Jg1FX2hW0pxwUYNO5/SULFurcVJhXCR3Z
mDa4ArxGEAEDPZ8dapFDhQwYhxM4ku4YoJG6TeYNGUe2w1AN+QpTAOYlwLsIawzGHushyuAbP6A+
wGoN2EZSrMOPigqyV8+hCGEfTF6zXNoN/mX7QgwllIL+MGsrMjCbsw45OdvMMYkORgIxBw/PN559
9CxZxZxTEN46awOkhC7PnPDOb185ISw2B8yuz4vL5wUWtU1ntZmY89hiSPuNcMTExN8Mtdf9jhUe
oVa23pCcqSmRMABj376h7cKpD0+JKVAIuhGPslhZ+I05qVHlMqCCVXfOi8S+jbcSwtLu4HVPWeXk
1wIZOjmT9sa/3ecGfCLPOOD1+TqENWMzhs7zQ9kUvbJrHHLy70FW8T7a110M1mO3tJALpPx2tMKJ
qQrcl7c22LO9UGhRskDyn0nRw6oHj1/OklfwZbKIs1rBdH5m/h4J9ONTgmoRtr5MKyKju0UuSxva
Rzivu801wrDHfoAbwkSAKYOuRtIkmYqB1IY8eCM7b1MBU8i+Hp4X/24XoyOhfwPSzGT1N7tS1wI4
83jmlgwrXsSs7tejWIvGu/cbWDy1OJOcXzNldWzAJHsrtcgQ4Y/PzRiHtWhdlPNsQ2/YB4sET57a
T0ukQ6n/sEjEKWzgM0K5Iqx5Sig6HUAu5Cq36rQIJF/6VkVxZdFoj/hz1r+2UCpC0Ud+QMs0Ze5I
MdJSmfPYx7SuYcGqvPMhbcSdU1yNA4XTh/3eFHfF3XhrdhkPhgnX8QuXWdXq97aI4nrP44R4JGec
GE1/AalH6pq7jl3IJ+Wb3YZcmdQmfNLAH9YqwNAtiUg6a0nhUgXLizGnUVvXE378Bywz7oeLGHKj
YKQBYi0XoesZhKOaTsAMSS7ggUfqFLwiMkv/qrv2O5Ca+an2Pvr18QJsEIRoUMp2PQzKWrapCLZE
XJf3JQdtJ9Fzloa1v68eu61dmgIU9v7fc6MpZVbgYbXiJb3yP5EOxijXSYwewc5VlVYiy4tS31Zw
81cetnYkkuprzwGZhxfzeQHQ7VFWIz8CWq3TqAYNZOHYqrNUeyJaD7+FQGxTvnHqDRP5A8A0QRpO
0l2WzLxaFzoUaPcoEJeTY38M1OMCi5fSB3up9LYwdmulyYOYsti5NxVPD0vw4HfStlzpcQrFeHQR
dqYsynZHJx9gQHEeF5RGSidH/HTWPTRYtRjH/qgHJImD8MLxjDufwFz/9IO0kgxafbycg1aNZaG6
/AxGvmbrOGtC7jn60h33n4VLSqt4QdYx4CGLgsiFVrhCrYQdAlDKW+qG250yzUw5XAka7y7Mx4KT
hcG1gm0bBsyrBSh8Z0Y3ElL/9FBh38XRKA3svg7o/N7jQYH6N+8YBNk+3SI2JUZtYbKuz8NaegzN
8MuJLtnGYeuJwGiuKjikVnSTC69XT4yqTeAiPwju3WWpF6r1zxYHygXiSDsiR5uq7bMfJ8va2Anu
Fj09MZuyUvl2UlYujGpnuiWQsNWTysmo4fTQLeKTKaBTH5gVqo0pUDsCNfEnnU41Mw9BoZ9KUFZJ
uzfAHz2DBwkQ+MWF+4T/Xmhx1DsGlSJKjd2X1lnj/AeqIi08lPBEP2ovjaJvBRWuTmCm/++jqGmx
eEWRFbtsFEnOFx3cefrFsa5KuOA4vDO75KwdXPC7BrlkG8/Tvk79xTEHzgpT8qQVBrW6HYLT3zrd
D5V1WNyg/+PvqQwQ1Jr55kkBejyOkBlKcPDSOW7SFURwBO8Z9Sfj2TxYf9KbN6y58WSqxSfcgpYt
OFZVWknuNuhWMjYWWGHJmPAu287X4PNIxQvMua/kfhn2ExhHQ/AtoQXaTQXyo0PF1PGknUJ4K32g
TyXuLhSMQF4RO96K0PkRTKRM7SNNrvdanN0FQtCHpIABYNU7om2SLZVFCx7rrQ6ID2XQnxv+ZYAY
1K3Cgv7Yk8DLWtfDztkEbchbcM64cyaHj2E9sDJB4QcNGpikVP/XmtuwIMo+utF//R6HAJp4+Wn6
K38YAsSWuDs6wpn+QcvNC6+E9a5qjG99hhp62kUCnSKWDHrEsArfb9bkb6j4R+dQb5jNmAtqNIxh
/cvKzVjg6+leLU6tW/6xZOR/48WQUyGel7SAbZxCqPZlGDn/HGsmSt42atSibg4DnYPRAMJbJ2Ol
vNZ7rPx46NoiO0F8WchP2cCQAtKllGdxtB3wBROrXJBqZvcUHT9nzNYuvY7QZMLjjuDrpfELKGRP
tptz/bGi4FP7fZGftLBJd6EYSMS6lp6QWiZwuiuFpjuGoZRYjZgIFRUcvkdlfXaDEcG7Xjo6gujw
h169WA6KS1caWSa1j3fTbkvLTS7y5krzvLo4EkmqLYWyXuxgHSwUR8y96PVXXU8uCtukoEtZvPd5
WmoUnYbMpATjugCBZO7nnaZXTKCvqIo7cVQWO2jjdly2enC2BiN2qzgm0OuSlhJL6sTCWZZMfJIb
CsbitNr4UEJwNIx5F8t+URrxGkjEpKHSSTR4P8KtidneWT5z2/Lq9jjKXyrrhvBri2H1OqcSE5ul
mHOrt6zfgNmXh+20HAQtQFj1FEDku7J4U40e1lFtXnarEGIQUsJrYJiRiSdcuD6Ml0hG3a5JfTZw
u8guDO/VP0OfQASb9k4EMiy0HArKvMoY8wHfF+x3t6MK9nHwDrNICkikn3oWkZJr6uIFCLGtAkY8
AdLZLd53qn3X4B+4BBtFDxNHHTvuTvfg3SctMQbFh8gYQsQaBgsJVGL0MUU2Avr6VMpXtqoN79y9
cHamJKmhVHSh/VOelqwci5YSbxmZepS0rUtL7/V3ICMM2DRPQu2SZQ3IRMckdTrBBws+Hl5JAQD2
iskmpQl3iKlVz5sXO0VmPpr+710eIjxdGEzB0MStrsz+RtAs0BaV/D37QgRQ9K1d6yXpS1yIJOJn
H30sFwEF3MO/yJXJ1RSqZwGQpYgziWzci64X/0N+PXTyYJEL5+WCg8hK5qUh5nCNAro90lLutvti
CxGXQKJMb8SCBctOOD/kNkcYuQbqPkK5F3VIDsC7ctlkk/bLc+fxj6bPxREEiHYN/TAK4HlZHBvm
7T9VhvuS12qbaYmr+HubUb6X2X8a9bzfyIxPmwj2ruHxTz88HXm+Zhp6jt5br9k+rhYPqTh3IV3+
RAAeNJGL/W+UKjemPlCjLGMg+IUF1EF12eLObmfXtvmzVl0HMh60CFkwwgZtfRANNqiUn5+it4TV
22dD0zAJj4p/JAtynygmigAPMq9i77eZO0tNEBAr66r1GbwCgzWESTODgqIT1smt5BukVXrpQUwV
/ljnu+MEVQO/FNKq4epAEwFiidmNdvPOtlOTf5Tqbm0yVUdZphTp3wUv+x6cFHQA4yyv68C0uLlJ
Ir/uXJwifw/5UDmfFndsppNEuwVQMx8CpWqa4R2Cvsg/LYDcKIz6x729jYY9M9rg3q+ClJEVd2Bm
Qmr2zMitIEo1iUef2bF/q0kBqidB6U/RP4W5RjoeNB8eKYFx7QdMa9sOKsACHj3e7Y+gG6SDU8oV
HIbVJiYOkvTZUPqahQvqOS0BODK7DKxrFiYa4jMakgJo1g78deEJJtZkiqGTIt0oMZMWF+yUHImG
vX3HLES7Ym2OJcgjYJ3htbcEdxOS7f6mMuT1OHcncTWznAfP0qfMmPMgxvpXfNzXdavFPyNeUXgL
hr+VaDdqDk6zLYSqIt8Axy0OTZ+Spv4Cnl3d5RY7XdqVN3PigzpnK4Pw1QUC0IEuARzmJ1HWvWy/
0vsWOCK2Zh2AC7YJ3PKXL6xraCM5BWD9wEHlIxLgI6D5IpR6ypUI0TYlEgBO8z78seLyx7kMtf7V
eLzu8xQ+eOzY71z2OGyt/9bpDTCiSR4qJMcM7ZBcVujAtJV7bmYptCtUR+F7PSAsJLNHVFKTtCvv
uTMeocPl5IK3tPVax7SZVsG65hljZEEdc6VuF0Wnk4xYOsF6V/u7fVk6zYqaLS15DOunF+92AMV4
dQmZtEQr4qGehms16Swd35WmplXSY7addsRueg5576Y/cklSuo9F5pzQQVdo7ZBZlqjfy0S1weRa
GIKX6z99TxvLRS+xwEe5l7a2M/TFkFB2wFfw601D2tIMtBLSN8+uPRmQCYJQM55HRfbepJlXobU0
9vW7Tw5+ysjlBQDK59JWMWAwVjmfZHcGBaYy6kYZNzfGCAmPrr8iEuCB8spXNXwhwkGWs33Z9MuO
lLEBADvUWmzZcz8SM2JqD4nDv5Mq0k/jn/1A+QzHlgipKZodJBSvWqOcgHWpCX68xQG8qWHcVzlW
UOhL1nRUfReo8USDa52vjYfQ4C20FWiRIwzPALiLmG+r5DVzLrr2Ek0oquIbPUJ/xOEuQS11W6tU
pWBiY6o4M9ijjkb9XkC3+jPVfdYZENylD8ckP7KezyTWhbWh5FNCdVZWa8lB0/PCgwOkPbvV6lHP
smbRWqda+5JlyJX9Fkm963ZvCP2xQi3MEU2bRpOc5MczCi+6P7DaKmSS1lh9HSjRheMczdGf702f
ZcUMwKQtKODS9vw9dqo1MNArX4S6XAU3jn90JUhPsYEeWbtq1ODfdA+W4370dxefYg7BxANBoWsg
FPwBRQAHLrbX4j5AJf2vvPNU4/+2eemzbW0bL+zcUBAKkZiCnR5dKdq0drOYoafS98EcCMNBPscP
JAQk/XrrYSVuy5nq5quUYfhdFXCE0FuKLN8ARjeY39R4RpBBqffVkK9+6yW+FPawF8AX/50GM9HB
EplTx31XZO5Ckts4QljRxN+yC3bz13HndAzA5MOCgkkzR9bIpEDPxufbtJv4k+UTUNuU3uCDwRcG
7tdGDd4ZRIc3MOuto/t0HwXtYmoOHRC7qZbhvVnuAwL0btXkJ85EPGWRWK6A5gfI2ubYFhCVcMhM
JSW83Mkk9BSTNndSr3zEVLK2CIuKHmXxlE4HMwPQun4JGeQlAjjOTLMWQAmZhxLl0fh5BGyqNjG/
KRb3t8zDUJGh47VP5ebxubFnQrsDad1au4GNvHB21mhtZRIhVeiknKqfHCfS/ozWY4A9kGV7ddBC
311AMdwRfBxzNemQ3kw1lXoloqt/jOkdcU7Cd9Q8QLacJGEOWx+pfEYSdz/r/4NhJutJz4mWC9x4
odyOzF/SW/Cgk7L8hOlXlFiuDLkLnICm+OeY2/p1egFQlpTgWRd+cc5LUXban6PHvlAVdQlfHy/N
hfQEubvwB9nXtO9t65BHmEfuj4HjR1nDdBnA+PcRAohaDh1mAyhMWg0yvwfjUjajmMQPKFc5n/e7
bEvQHexNX+RLjMOZs3J/OnE90rK4D9BYQhVaAqNV303XkwuVeBpbtrorPwQXJWXlbM3cjwizdCnI
16cT+BaR+e31NERft9mfGLJ9inIfxEqlP5XuZn3A9gNPam2qQ/y1iK151LHIUeoF4iwhcF+CaaOw
QezM3jWo2KthZVWdVZtZFfUjTM3tdCZjwFe0esRAAS5sxxl/ClqYpgqBaPWSRsIIbNivMO/V3Dh/
dh6IQOu4LsjgwdDgztxyzMWWGNUb1I+SYf3g8BOg7qV/ChILwE6rPMpX3YT4fVlK8hcI9Pk6Tgn/
xTE6jANVGWhVAZR0Hyi+GMM8fcoJVHqgHTCE5XR/SRJX2I3Zi3OiBHbkEzaElhGcTCxwu94xwy+o
wY1/tqmZ27f5DNmiFf1JadjumLiPQOdiIGKJTTEJK0emU8o3f4F28myCoBUVRqlfr9UyLYzGVao6
yysTN8meTWEa91DnoWsoWS/DmmJO1trPi+Q7NtsvUnRJxUgX5ILfhmBRftucTN8AKyMPWAj3al9a
98HOYQPS01MMWZ+bhgagYiXlMlNCA5Tk9+UHp3ChLr0SvrDXcSgh3+K4lOVj7FnFPuSqDVHrY01K
FSydYjESx7A8SG5BO5yUPExPjyf+AJ9f4HJJtJS7e/rDFUO3VWMM9KJ07xk7w853hIyC1VEhSf3e
vKSAgtllKOkQvaM5o/HIPR3mOfmz9Y2vpgHFGnxQcOdWsX4qwI0iqzwyBdGEME2UTrOs0uwYZ48Z
IPyc7YrSR+H3wC3G6pqkzvY0eLPpwPMVXL6YJ7+Zg2ekVgJx1UMLOxc7ZvUDNd4F9lKWtxz6YVUS
M6iJ/SCyWDksb6lfJEouHynJHiY+f0WDM9bmII2bgqIg2r5/3mANaAhe87laCr4fKEgu0sEwMJwQ
Ng5O+1tJ+0KTKgt3VraeFN1NKGRiX35Gilcd2uGVleT2CUNKWUYSZqMoPXU0Vwvy75DT8QIKLRP1
2Wo38kBcdeiBeMKZa1FGUGJC5Krp/0869TFE6Dd81eZIxnHv/acJPRe101Gw10DtQ2MKCTMYwmJL
emqzgrdRMD07e3RFkUCMnsF6XndwVX3v+1pWD2EIJMZYR+YRuz/VgXsceZp3Av+xogUdsAOyUvDS
k+BoROK/Eocq6RqVcg1+PzforUSYJxx4/6YpGKqHI1CcLkecsUR7OYM+aVmcm7jbRzVeks55JuhG
mqnddbed6mk18EetuGSMKURyRMESLz8oQoHyOsy6ZKSXWyfJ7XidiiVjvmT/ssiyO/DHcmKrMU0l
rvmbX7AIRn1FRhDwUlhuSbk+1qeBC1nmx7h88JnfDx4rE0YPdYA4yLaZb68KGXeiBKo26p7oEOUz
lNNY13xb5KWYrywnixQ//pOxU3lm3qdm4V2jdT/Lf3KsIrGCOn9eW/u3SQz3sz5YVkasUhDmeC7S
e30urtJrKdRKKnsZYIZYro/c1GSlP4criBJXaCf3m9uUB6vM8IK40KalE51Br54AmaCV0xCY1AAK
dAHfx7X3CKYk8zokx4GJRL0W6pmurfJWVCNXIHlGPfUbcwjq/NYy3gmsJDIKm3Vx96V/Yk6u6N7l
h1uQrztwo6ujom5chE/K6Eg4AIvkmImmgpnCnsb5WxNnlzTwg4xujNs3ZcPk/jZ8KR62AOUs7qTF
TY8PcvM4yUk+pyJvxuZupnuoe5c0h3Hd58SsTmIyQfPRiw1VMyxv3dXzriv0u7EYI4LDSzmzRSSa
z1PKib9bQBKF3wHvcNyQWVd6tKeiOVWFaW1vRbzyPJwBx8UUmIW6cEDJUakaA6pi952656sxCkhU
QIQbR2QvxSh73d0gtjLzdKLHcyZBPU/9KaTGMWXS2Y7T5tmp5W/okV+t/EYsTUx6eB24n5F1JOm7
cK/7PGlV6mGWziCbWYdmBioqTHwM7S4N5Dj2IQ58mdzuKKaq09jQlWCw7B1w0QttoVmF9Yoy2QAz
q5mZTuHzLpOuCZIjAdXEOwRmOcJ2kB9L8G+TaWScVyRiUYiX6MYNBWjxj6ocveGUVfLtb3XBlvK8
gu6FVvmzRBTOrnZumclaHxTh6/Q/Z0OSwGvVQJLZd+r6ZwgELRrtShR/ay8UjFTxO+XSVya4tJ2A
vZQVKZzGAL2HSv+jtlQoQjU2ugC8hQgUGAsAE7sr5eDQYCdeDB0Oc9IYp03E3vnzNba6FpG16cmH
BP09eYZ6NSvvOHdDyxiB39F0O3CwrgpMM2Tc9b+Ytid0a+ZSvlSIRv1g2LD+viRJUIwnGGlHCqE9
Dp8pLode59rH8fyLIy8ZpDzcM4xxxz3K61nLksE38wXKh1rZQROTlnvdBz9ZmXBcwNqc5cA+ZpZH
kaxfMD/17KNoz0q2MGy2geHzL5f7pqKpPwbgdgj7ZCVVsFODz11UeZnb2EodWah/fhE4LSSu7KjA
527ZT7jwaQyVlNIpfxdkISeiHd48edrx0F3RrLj5hAfxMqDibuMEW/YMdySac51hWbStO9tZCjrT
YcqXX8N34A0/SI5aMJumURTgnXXPhoJe2wJoUCJfZCxpdsAXk3sAPCuBxmf98lHHIWMb3mgjamBc
eOSzZp0siFKRnd4YnU9cDanGdQchqF2QaytpgMGrOorx4zijnopIbdFpnI5VxCEXjp28DS7yVu+r
X4c9jmLWwgUbSoH2aRho11iK3Nha7gkJdcl7gy59lF0b/ubaq1mp0/ejtKYw0mt2zfGSurXOPwd0
O6g6YnsOcG8NrjZtUnCIdeDX3uh6VtAqIQwCM0Q3cVT/RMLCYqb5356PkenQjQIUpwAwKnIIjxLJ
QzOcxsxJBDedMLHnRyLMgEfubMUuKAHNE2Fd7d9ZwrQBC3HnHfaAB0NbZ71US7PW3UWPDc2zXcq0
60shuhsICaW/Mvt6iRZzpVh7f2o7APqRxbER5IIIN4b2jlLgNyDKaEklNSYOIfd64EmrtcSxkSwz
qVk4SaXD/xVPEyV4Te3OizLJpXNjlmndfO8IFopma7AKXoO2cttZUke07s/4jedM/P+vvMhRea31
Y9gCQhrgw6/sy3aVuRpmQs8pQAY/kxnqp+9wfLn9EqPSuU/ReiRqIAkPLf+eOhGMUTxrYMv6lAEX
4JrjUQqDO62/URsNDwcXPcHJsSFhAL02Wrs5nXJ6uvnORjN/I2q0nd/TVS3blOTaTYZEBPwqQx14
meeH5VNV+viWsmJfnAr2+XJQLt5KnvaRJxctEVrVAgkFcowVmjxUMZiiTpxbUuLBOfXNjIDGcZ3O
bYgAHaZsarInolnFFQglVdYuttcZJw7eKTfNmZcTT6kECnkGVrnLfb6f6xDQvtSkE6aZj4tat4TZ
Th7x2pRVBKx9LmcFRZ07y8Hz07CBmvxx7OOnVuZMKoMe7K7Rxqn6Z2kJne9ZWoBlqasKuu0Xf7ZY
t471LE1y73SJIv38U9wiF1nmf/p3tNJ5Cr4/aNC/WVq+fR43iz7nIULCxESvPfI2n/ZcIYw/DskA
suZzFkoPDSLG6di0ZwyruqKNZ4h/dGVEuQ7hxfL201bM8yv4G0FPmpuZYmgFzhA1nJ74NDe6zRvk
YedNGsjyBSDjXKOKwkcAgsP1DkNd1w6RcWvicZAC7vbcaeq2weKsBffaWg2MsBlDYG5hYhEJmd5H
yFHihzKxk+UsyaihFJPHkWGxFWHVuUPqW1+1xacGv9/DKPay8xMraR0HKouCuM90ot5vaN/aUXDy
v6qnVgadC+2W/f+1Xgd27XRk/ZLCxO9uWVfWeupA20eecK68Wv44C1/4UyoFJhlX8O7RbcbntWV/
0wYf+JE/VyfZmzA/aPKM4FfqwlVBYefWGMNrVqA0Kkr9CwyuhLDefGGeBOJ5lJT1oQ2ZKL2Q8Z1W
crwemgV56p9OhAhMjtoJMlw/F2hJnXeNJn0azWszR5gyD14sFEaVUzliik+hejKh5hmQoXuIFqTw
x0DFF6UoNbjqiz3occAW8MXXv6bDEjBw8IEjtnJn0Y48L/nugrqpxf6qKLgX7Xh+vX+lgJkwBVXb
cQO7wjtkt1g4rYZjRMFMmiSHRpz3+/9KuR0WFg7KFo0Dj7CLUAjaLQrGJ4LQExvU/u8/UKh13HJ1
z4udeqAtoRy+4RGUAsy49SWnDnVLBFpRZuLE6SZvgyeQJFrcXo9zvkhuWHst1q+KDNLq9Dn/H+GX
1X8H+fiLtg/u+I+ru7PxroC+wiidqNLGd4e0yp/UFp3D0k+IZya/uek67ZthNn2p8zTt89noRUc8
5K8/kNsI/f/F8SkKyqiVMj+oM7i66jiFi5zaChN+jiz0XlqysCjjSWYj/5UREnO9dT6m4cFWNMdi
lxvrGXdulz5UmAjNupQrwIIwZlc5WHxD21ETysOpMPE4GqqM4i+E+XMfnz5/F5yYhEmhaJtwsVxb
9U7MpP7c0t/Gw8QYUx9zaCjzULFy5R4/CSWs1yC6Eihl/TxFgib645fJUwu5+YTDXz9bBb4oaFQc
KQRqY6loI5P6qGAdbBpxxp0UvryrBDr8n3znpPwTbzr3PQf2dT3v3qW/25ISetpxuYFP1zwZ4a/1
jTF99mWCTHpkCF2emF2ehV7m928McBMSAqqmhonjKN98yIPvWFT5RgoxZkKClBwoAUQWXNAeFqPb
QEePvIqR4pDeAQl2wwKC56EOjEWTwU//6mTdbBEllPdV00DQXl+1fG37ovdUcAWvwwUUuIIfhzQy
LAGAtUX0z7QyliClXLrFOdu6npCkgpuEot4csAfn/7j2bXExOsPcc0fOl6tWqfKVz6/GmUy/WkDK
qLJSTeA05j0GxhGEgy0nGOlO0p7KkWThurVoDhbH72mOqBjIWcEskq6TVoyDnMM2DRUdVITDcxPU
Ke1JGG4a+2WjlFUXgzO9VG78WAUCnvO07L2EfteG0gyMK7u/0tUIllZde3mXrMtYHjlC5jcIgglG
jzuHcPRJlABSBdYw3Z1ej2TgzQ8zSsjz7M8hk3uCeL1CyaO3khjD4KajX3EVlvpY76DVTDQSiPyY
CHHBpVWlKsWCuKKMTp6zgsU4NHY14T4UOZBnUvIW/WziOY1kn4mqKZJ+sjzLvHrAVXkctBL826gF
XRYSiat8x4OhqJFuT620gKQVuQu4dKDf4b4QTRpd0TT0+pu3bUUBJNBg+XIspSVuW9FRnKP3up30
U17LZ/aPtbFyudIHeINN3BzZUHWYxht99rpgsZX+vpsv/Rm4El4pcB9N91KZzvd27DjWbqYLdkD1
2024xFDsyluPmD0EnKQnJM/OXikhfPOL2FcUiEUcqvWylkTkmlAbekrM3nFrPjMqicb2PFrIFxTf
kblV15tV3Xivtfq/h1E4+BHcoElEmaWy8xbdGEY7B3T1rys8F1nL3b8Y/nlWaCXnjkpINMMILdYj
dX1MMLP2CvBrUy5angBD38w/8eBcF0lveEoO1kHyxlkCTPCz6T5P1MbLh8D2P1lvnmCMtKrrnxx+
jjtlJ9tJdHKeuc05bB+Iq/pdsBmVztABfhqVwk0F7i7E7/zHad7SAK5wXt8UF58wXZpdZzWYi3Pg
O721TZXeBFBRmklPGOyxSGZtCFz5T9Hp9x9nexo/ppb3A0u5MqD/L/GHztsNB44wk2qNkhPxlaaP
lfsO9KZVrgTxAY8Fo8XPLp2oCNw1qxhfGpbiJBiZn/f57heL7i/0LdcH3DH0n7ZY+6HrSrXLZ/a/
E5hAfcH0gUCXT2oVB/mg/aRPE5pn+rA4+fN397032HQ1YjGt7JJ/QW+dV7FMBC/2DLWcW1B0ZPbT
mT2JCA/ae6UyHq6c2ROjOJS7VXryTIs2+SC1OLDMQAajDbnb+Pwq6kSPNiCBpuHhx/X13p5HQHXN
oEfh0b2dRs5AOmhSTXIXjCjdhVHHIvOrlLGt8v0dzIy4e90a2FFlge/aHw11LGkkwtJgvae8+uUt
ljc/dfJ8D8UkfJhNs5+Cp1Mt/Z/lXRrl/09tE+p4EeUYc9p13YRMECwHP+jtPp9jc26E68a17q9H
scfgCB712H76E9V/j6MdE2XtjUyCfrhH8rNDPYZyt/VPTBbSaXnqqKrD2I6MMFxDepiRFNYZGrnG
SDrcgVVW1rpxNTjNJGoLM2tyDZZtx/ndZKtJcMDyCKutGuHIW5T3/+Ai48HLutvgLQEhjd+T/yvo
yQPXBNb7wqkJXmG1TwE3zgcAV8e3N92vcs9sog0VkXofpyGj9c22TbYwZx3m6psLIcfs440nUF1M
0B71ATTO0sREEDNoI478RUthltEOPERyOaDvivLjXkO5wHk5q+srgH8tbU2LYYlBT42yzRDL7qNc
pI7QPR/711JCTOVCt7CMg5pkWoJX/c+xjFYauVPV6foLY0BNXNPCXLjQmTmK389umkMFX+AvcFfR
U5aRtHib/j4OU7sRPU5vNa5vK+AnqJTysdqjziRVmaJv4kHop8l0zM4wpWeH2ZKr5tXlkOrHwtij
3zobCUvlpCCRu1nwW6Ns4szJDX6mAddeYlUEICtG48FsTa4U/v04uy9SpoXKoWwox1mNgRA36KAl
BeVYvq4AvFvOUHnbeQGqMJ+5lSCSIpIctA1GkCLMtnKK2iIhltzi210mMkSSImk73xNQzSj5/w/0
lWXFMnWdrWawNdPbrIjoh3VeQWoskchfK7EiM1QujWqmTKWy21bp9ntiseeWPd3nmP6SIm6nTJQr
//H+Wq0+6CR9p77BDfukW7Sjqjv9Ut7LzmNmRFQc3cLvcexEbTxR5fzrs7CECmwdrXndXoatgE2x
1WVi3eUwk3AxVfFERFQ2JN2igsT2NxZC4+J+mgiYrxrkY4+NAqZfaLIK2VWqQh0Cwwj1sbhXztcn
G0tpWELqsWmJzrY5j4h84V5r7u9mCtdsyfvAoVs89gLH6rKK2L+cvKVC4xX0tDsS0TCayGNIp33f
mmE0u8Hc8Ypnnjkkx2f1RRoxEjkBwxB0Dbry6P13/+zP54k+Q0fKTONn+Y1RPAFM5xj53ITrKRJr
t0Kc7vm6Gz83Nxsb0D8Zn1+V0GVRn1glno+HC6zU5MUE81ZKzVya9QXexF0+FpIgN9m3G5qa0A1I
mtJvVipZOytTEU9+hqJ/L6k3eSlRpvtLasTntBBYggPJXzcHi7iaJG4EhvfYSq3zorQYW4UZGCq7
Wvb7O7d2TbqtT/IpW3BwL2fYVO2Bd3RcGRKxhGnNsQoljc9w8jfF05MzqVAKfNuLLV2FqecyS7eP
igz5qy/L1V5vMC7EOJ/YbUzlLvG2zi3NCoEdzhMI1PezpI5ZCfebbAZDNChbHa5O8q6tu3VPbIc6
eaNd6N0G6rgk9bAbQuadXIO6qWADPlY3x7Mc6skNsiUmDgb3rUmdXNLGkPua0Y3M+Z9evyMapKLf
O9Id1+Fb+AJsqYFJ0J2eMzluRK4IlSmATYPZO9HfHmezonDF884cTt7Icpe6daxO3OJJlDRYYRwP
8zm6FB/yEuVe8tGKivHYWO21xyoUvPfbzeLZiuAsDy/X0TKNPA3gGE6uGAbBpLnkufvc1n7j4YUS
Lpugpl+sUcSKAORxCWTPlrZHQQEQ/7P0gQx5j2GAYyRZv9Vvwhaila457YY+Cj3AeOcH+287z5yw
09t85Ta7MZDppdaoMFaNhQCndZytdo9STbm1hCEcr6yOd5V/189/QGENLaKWhBUZcqV1McgBoI56
mY0U8R4CE9txHKOEcULBcoinNEuj0KnD5lhujc1ai7l9r/ni4xuBQW3ge/cp47D1JPs5kIU3DRfM
bgWuDinZha4wc0LHi23QQkTKWPZgR95t8579IwlGH3RafxBpclZnHYPQt5yKBoOBY27kUPB/Rbua
Zy2Cphr9RbQdkTnjmHXjnKv9VkhYvIA5vE0iJn/a3b4g/QxL3wiIhkfU4xMlWCcpO163GWFCTJ1J
V4PZAQXju+ZUSWqOVyeH1aMgsXkKDvknA3Wh1Z2zm/J+E9toRwJpuUp7XHfzmMcPESk/QS2yLHQ7
odQMk+9vYgfOWvQyIxJepvPJw2QiY/hDueFRPyHGqQJMMbYw/lHLm99g1AvlGGsOx6jiPdEwlvsp
dVD+e1+HZYqkEcvwYfEQ4B0ezqwHji3A9sgH3+InoRI/OMxAnobQXF3SS9raX7kFemsrj6yRu7Qq
W+XvHPcTD71HAwYjaH6AiICLC8xVPlXWOazSOQPls5/2QE/Qz2rtzkGoybARL8rn9EcllGY3/y3c
f4O1vg3NVyiDK1EeEvo/f/ayqfrmX/qFYC3c556bdye05V2a47e8C+Q1hfZdlCkn5OxA0d1lDFXg
BMHmetCnCKi7HhNFSzcJnCK+TUKyCVe6bv74sN4bao8ZE3O9iEWCadVEsq2ZnMDX32lR
`protect end_protected
