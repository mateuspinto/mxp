`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
Cg/pwEZvIs1Bd+woV9992pAt1kcdFnVOm5bCyMU4cnASd6YpWiXikHzC4TV5xqkj1Wic1CdQH4NR
cR3oEAyPClJfEXiKGb49cuq/0dmf/gXYHN05+MYpCNQt1YSYyymrr/xNsZqLv4CsrXsPFthwMG8p
e7G+5OANCjxpZOuoapFvGUqT63syiA5s1pSBkX8Vhx5rehOXQvszYRHDaYrDPkYAlRk6osmkSFYh
aZ6jR4GYuzh/OKWfxIJarIW0PYETEZPRlZtZEKk1Nzr6mnTt1eBIdxRD9Ge1lgSwLZolEy3u56hb
ZHA52oXSSjM4hfmBrUwyeuimOxkURUexMxGeJQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="8BSozYmhE5moPXFhG4/lkk2TUiGn3LLij+7eX/C1mgM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2368)
`protect data_block
fI+416ZdBRboRM7kj2Ws8AMvUFKHpLiCc2pZUenVhyswlem0Fil3DzE5rlxojt4cHsRic0HCfEBq
d4GeO0vQVs6AiH81Q2vwUC1k5h0osAH3c0oXjQ5ERJQIt8Ov0yvNMfpsMcL7Zr8A+we79q/qZtF4
P/HZCu0nLYalbTcoqnNzFDK6xSybXJJA0xiUlSZXwVLqYHV585a+oXnuyqEOaQ9m9bnGMejHyqwX
0JMhtdzqCBJ2jcyOHy07vX91Ohk74XeD63wjAcvjYW3Jta7RE50b2+uDMxQXuRzc8AaVhMpfcwC6
js7nO35yZFgNt/ikALvLJ5IRkZBt1oUQ1KaKjRt4tk2O/5djk+xR7SPZkNnUCcwuRGg05WjDB3CG
PZ3v+USYXENQlzeS8FuqblQLRUsRO/rfJFRgULPVsTIVAmwozcjsASVItV770dN7OsFv2ecDVFom
cBiGA5AaDh1AXqt5DHuObxhwTb3LTbNNLgtq1wkvRWdh2aP56E9wpMf6prYDmZElSaRRwn15cxki
eRlra0IMtcyLytocxFm7bAaClqnps+WqygSDLzJezMpCByhFUTGB6f6DrORaAoEhlT85J0rhxbjq
jf95dYbBGl+CgB3BJXGPpQPGbAnqqSOYjZNVg/NieAJ5jKm8VcBqIEhP8bNva3EKKjnlq6SLH180
hG0dWlBfiuIhrrNe7mpxR8zALOo+rAH34JbLpnwO0kfeqE4lFBVL+8rlVfY8tGA3ty3e/s2vIDah
DaD7iym7j+/u5r9dGCu/gOnVpDkgX4iD/Ba2M6pxl4amCaZWwLvooTlbaMD2kCQGokTDaEeGMyid
QsqfYFDbs/3XAkhK8IM7iUPbiW+UeTjgUxIuN9NEhGe8kcJl/Tv8tV9dQl8dPVBEU1CWzadY6csu
dGZTnC8B7RAxTMzMUdg3FRg7EZ8rHe4C9985WU7ctkByCpLCfPZQ0/PsbMaYiHxOdS2PGPp3fGCX
tRu6Kk1EjfaytvIP+d4K/lZmgLwWKJnubSRlsQwhxwkBnEgMt6k7n4yEKio8dVnf+zKNbfGpRRXC
qBUb8Ss75TloWAmn16QgTBcw3nw47vgeFAH3k6MM1PHIIbBkOUpIneajySrIcG6jipzIWkA3fpS8
XPgOhaKXOqssTW9Mk/HIUmKGUdLCtaR0286oEpSGGHroreJh+2j2SkSJit/4y9/3Oh2fnFbAAbmD
1lpc8J9noA8qkn3BnuwVwxanc0CZMUS9Uzlb6glL7M5L0N/zB47L4vxy6VuhdJMpMm89WTE7I3Md
0FTtCzVvCeUj3d84AJ2k+l+vb5zpv4dhYHI5DFJVN3UUmNXrTbAUWIBrl6XYOfW+3M42hjEmS8A7
tkB+qzEUxIb3rTQQnM1azAdEpJ1zSy5Pre6MU69xT3C5FqHD5HvuUp7XqmiVRhT3t3jfl/4CraIX
TQ//eGB3JptEUWhONbzb4Un2SNEra4zmEMDoV83v6I8NOq3nX4Xesgnj26Kg53i0XTNsbQuZRzOi
Klt7GEUwc3A6+K/dXdfqZF4VAhsX2zf3dTA4UZHAWER09JSqsg3EY1xwrmVpAl7nx5FMgSPEQuRM
NLG/yTrk7YiLMVDMEheGjbVaW+0mBb9UD0IRB51FqWN4Xh32F4/riZsAGO8wQMMUUpUqJ8FVNdEm
6PFU6G52mefJOHKuGwwfspQNAXzYUxc18GSfbzjtqMzUtXYo/yB8up3QAB7CGkLVj0sFVzZz6Gjy
EFlgaP7u5wppRAX3ZEY8xe7N6pXqzNfQhf6BTxvUzkZlyT4C/NE990+06QkUzuwAG9vYwiGw+64t
McCgzBeeuvwXQRpstXw7ncYt1qSNVrOTMz7r3KEc1vaKGdACG7Fi63gGVOY4hMCwpMx1MeSW4DMo
puaPDxQS7utmjlJiE7fYeW/ij3r6iJ0uqdUDHG/67NU59aet3RPvNeDq1VSK7jL3a04gc906Ln8c
dnC+ozzrTtdtYOKq16x3S7ur6cAI0gyquhc1inZt2aKNdwEUT/UskYwx/ExO6B1XDV355qiMiqI5
hpj0ms+cCMdhBrKu7lGdCkck5j4hZKaD7aGQE/B4VJSldBcV2igukt2L8dP1CUZPd55Q5tLPtFsm
7h9s8lYBD4xt3Bdwyr6neVsjW6clGl/LLOsE2FW30ZQtZ6Cjf6pDjkuPsbpsx8hVV/1nwFXn0Y2u
abcedhjodn/TeFowDiPFRKQuh0PfnwTNvkwOBVSLLGWEKcQsp1D8j5dFzuBhHfHvpefClvXK5pPn
zqjpJ42Ih6b93wRXUhP2uECr/OL5Ty17T/LnpiccmHclzsUUaxfVVG3StdFupKPxVbWPS5wtgc6E
5LPVuY+tlS6d2EmPHC6lCCVhJmkdplaeBxMD4IN6+mhogzJYA7AN2D32fJ3b8snluaxjxES8TKjw
UYqvnKdCj9b/2U7Z0dk0PyN74w/oDp+dqzHfhlpEtnifc6j8LBO9Vu/2nZqo8HkdO3fEUfb4gWm8
F425XhzCSYXp6RCHpw9Guzb5kZJp07tWuV0Wzjf96S7w5Phhd4i4THIBmSJn8Ci/22Ae8ybeitxa
hwtcgciLuHCGmMgamZWNJwipiNPqrQOtOft6os/IxpYZjRW8TITyynCI+M6aI64wKcOecrGsJHp9
SsxQlycJLmGzO536xxIGoqDEhxdW2gGoP9ah3T9GRc09R5QUKdCwU8iO+TWfG6Gdm83f1OnXSnsM
IYS9wnfdWgO+cx9eUUQ52/nQx1D2JYVEedSQf4WZBUcnOFTOvFt25PCh6A5ZH1BvzXga98OfyuD+
c4MzD3XlLT+jxdLTA7V2VBEDJO55BWBUMzRWl3I3wUzZH/pkJkWBkT+llVx/TkVnLanhpVqWjjk+
AcjR8gmFe+RxlwbQRI5BNPc4o4t6612339nrQp0KiEnd/bgeLx35bJo1H+jyYn+1xVwkvgmEG2nz
bX5qKZ8ZibnPTExkr9UTbOD9Q4NM+qqRjl9p6I9nsDRyM6jBnOTOEwS5HK/GVfZXijwA4esQ8Mob
V84TLQ5YPdNBFm/izjKPO11S1188i5Kz3lKybzRGhYXrDnDe3QwQ/WsLL3FLEFBIppJpX5ktYfXV
brTsWKp/GgGK00juvwxOXk/9gCU/w/aCjKS0t9eU2w==
`protect end_protected
