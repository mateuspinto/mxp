`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3488)
`protect data_block
OoRjyePSHw0ZoCNBE7vXvK2oG6uwMSg5Gx4hO1UD4pEj15cqQuBeYECY2psW3ChjeBcUhhuZvaTY
oT4qstJjoiLHp4a6hgH3m7CYsP/qV1yGd2b2bgcDf1tYI0iCYbLY5Qawwz/W22YEzGJEUIk4rXgc
5snLvZedL3n05YzUpJJfqer9b9NZ/9YwNrwH9RYJ1Zw99nWVw7buRENl35kE0evelnBk0fwdNEQN
wxuxIPGmFM8XtjMhB1vMdyjWi7w3J6mr8wxOHU8Wei2pJ4zp5mlngN0aRklQs/bEumBH2eMMu6hW
dJ0PXJm2wEVv0SbNeGxPYfv2SCYj2cY7IY8mxmIb+0Ek6EQEttFFrAWaFhQbcpjb6IlHP/KUurAs
WsaT5cU4bwFbKZlZxKSAmmen1Fc2ToR8HoTAwKlfdSiwS9jfiWrQC5+7fQu97LRAfCTDnWZMio2E
RScKE5HJr299OsEOhA4VOszo5RP+VdGswkvIHMinpQQSwkNLz8GfHKIlg8q93wn9y8AOIZjZsDBa
hP82r2fXVJ+9XjZ3RPOznDCMHcDDZnD009PCY/SpmLlCt1o00jUR56HELom+6AhCJsEu3xvTMSpk
m5ziH//0E3xoXb3PwABq4SrMz9dmuMGqbBmTMeKbUFb5z6skWLKtNQtJZjlgh/MDOFwkml55euxC
JRrflEqwCOeodRQIfRb5RAt2vA2A4CxotiEesOMvc+BEGtxoLWAwN/YPfEm98+qMLr8s5m0WBqxt
/t7nsGtrU/acQFODfs2Rf/3en6ilx7KcyXe6s28KUqzAL6ZCiH8OYPmrcDVteMJ/Oo34Dj4zyFZ1
2nRZ4Jjp55gB0hxmCCNJEA893TJyhKSFTw0PQXWgaopuL7bnkW05kEeI50IwKsNX4sSURnpAbA3Q
m2Pb/mJaOST3FpaquD4QQqRZmv1sZVKqSktJLcpKu940B8dBn4mDjHfIFpKq6hK8LBqan9vtlN6B
IrbASqyNgstVFECWj5oF+IInoGZaICCTX2+7Gbf6EF3aJU6YjmztRWd/Yf/hycs6OiwFBfdwyjtP
ZqN5CHFnfvDHJ6KhtaYtN7GoXNroB6pKrE2pIJShQI7vj54DtBT30q4+Y9FTJE0AruAdAHL1+zWy
t1eFvAB4K2+XeB1qKRXrDbhJDb65bwSDHes+8qZMjiHmJXmZCEMUZ1u1kVfi03rz+kaoHconocgv
r5ef+3rZo8BspGnQ36mAdfyE4eAKJBjqf8MzRA5J+18xgDgI1umkAxm4Zv76Bq7NZaPsjzFoKFGz
MgqJ8OZgzmGD/yk+oxgBNuehkUq+mIwq+6UuRUL+RitpJmy4cbPwR871g02ZufbaeJieeIyae2Dq
VuGcO6vnYFbey+Ma5E6E9vgKm+UqdOdRJLSc6WIu8t2csLDLh3hInkhBWL7w8QcNFUsJeIdPJ5XO
RNdL9bMppSdj4TK3H1HD6kEHLKkgLPnpViWD77VFlZkobp4OgB1SDMhYeZlXaVqDrYPOEzcVboFM
SbPcKuLwEEpg58pLv2qNGvFi4aN6cZORjXOy3Eg/pMku2aPEBkQXBv0pYLm54D4Jp4ErcMWYJY+K
lueqry9ajYt385Dc0kjMcFcEL4hJJELMWHVwu9wzsT4X2jq7pOTjC0GFesT1YsGoxBvK3VieurzT
H2L5YBKTNEHmHY66YgmxCm3+rxUk8/1W/dh85n0x+73EwS1swsavEsuOHYRv3rttcwKsl393DDY2
Yw2L3j7+LrrJWL89o6FYk8OVuDDNVxMW6/lByLrDBJVF5/f++L2tb+BrYWZlcfWTwKjihbZOIIQc
SRa5eT4w0lSNCA+qAqq4oXm0V511IMjL2vGJnq5ylPTuAfwlDxYk9rFXhEcEJjLyjVNVeDTsPvF8
6EFmfucqfS9QMeQGEFvxZPh6dP3odU0+Jld+f6xAfZeUrti3pM0eanuUHspwEzyENO5kIehLQ2Ri
M6f4/ym/ohu0xgqdRiqlnUu5D+VcDcACOiEvDZ8Ntcvl8FvXri/SezUIK6dtz+/bJ7F6PSIhwqOT
COrFHYI6Xm6fcOHtGY23BOLgLg3ZG9zUaB7iQpgwvo0Pcj3FM077a4/dLWDZM59GQk41ujgIcqmJ
KUEsBPdlaOmPwzEdGEX9W25TY4fdmpaN/ImX0OTwsLHAoR1J/SZlSQJZAu+H5pMHVw77E1B+LXLj
gmkbxZfbxmnCmPnpZ3wsMpEmosCs7+R2yfRDO5mDXW30gSTAWREJ7aOhmRza9W2Yl7WINQB+4cJy
c3BqKI6HYD0LV4czM1YWW7F+dimtTwFiXaIDVSNmumiGUdca412x8tTpHFaTsNfb/CGlK2jxter7
ZJs/PeVwQ7NKi8xSjW4G0MBxyydCpvHTINVxvlHrtRCu6q7qufru0VFFXkxcgUQUv5rQAjmGlpZm
jTQkTLC2UkBc+w43gB2eFtGWM0asuKpdWsZMIWCm1Y0807n7iJVoi0A23rToun5LH0ZhEoHjMUIX
yGFYyoZzYMuj2rmy6fajihwwUbQA5QESfEw8vNO79pyyXVae8q89lqgSp/vM3AS0f/55xvrOb3yO
pN0cT+mQ/DD8nSjozmjEdoCnPQ+xj4p0HeMadmtzG9LiNNata3V3AxKFfdNJ+vsJBnVlv8YCSZyp
BY5KkxR1k0gxGtBjDVbztUxjCr8V1sdoeS6HBou12UwIvC7UN2tL1K5m7Excofw8olQE9YiaGoML
IiGGXIdx34d43+Yh0Bo+VXlso4pRy/aSiRtKL/FxJCet78gtxpQuxoCcbpXP8iofULLoNB8hhPMz
bMzvSyvdcQ17gRR5esGn6bFhDV9gvbAfM3TU3ipOzpdC4vSzdZo+nwfKclDstOEqAMne35v8Dy2U
XzUd62EOq6ET1UIUwM/J/i2hQaDiZrALSPhdvJgYV8/cAA8J6dOTQ6jkOFuu2nwYYn4N+Ot7Y/vt
rkwGVSyddyMxuFKvuT7JBDbC95HThXL6crbYYnK0L31VPl6g3pCDzq7po+CQJTr1mMQheM5N0KD9
kclum01Y9kLGrXYW9O1HBuWDz6BBFM3VmMmE8ONAzIawV5xhWm0eqVApQ6/+mGWvkHHY8GYE3t++
nWaSN2e0qOnda4zxrs8XVAReVcOkr8MWB+KCkeRm3XzJO4EunhcdwcI4FJqC93HWL5fTqnmg6e8A
LvqY8/GJV0Q6hcsUPdCdOQCZ7zk7RxhhXNC0fteNl9ajeQTMWjvaOS1l7KOh37vuD/IJMaynyC8d
Er+fynpHIpCThcT+y0su5MJ+vgk+DEr+tsrihqSKXqmflfwDxkPDC124tVRz67NjyfYd8mjW1xAT
0xxmw4DlgTAwNwp90/rPrsXzV4ey9uwFtpAeuO/XiRbdQX9eEvm+YpH350rP2dMixEfm8tDWsSg4
P43053f56Dnb2tutFPg1Ll1/yLHvz2PHIsMCQLZNhBrUAzDaMMY15gWnq9xchnc64g6NylAl2y0F
5wXrnJUrjTJ5BeRrm/Vl4G3pDk5SOF9UnD+uOlgIwooYJ1Rxa0LNwo20eoxn5kwxLExK8r83kGih
jO3uuxYwTgqE09+Dmx5l+jmHxGMnST9XDObx1p962afqqaEsV+0pvSSwhbPJQ+G/0ea0ZlF5ZxLF
3WTAZZuRjYqUBr80oOkwt11fdhcv5c942uVWxDzz31rB+Vxc36bmAsEtocvKpGoWFFeo+h+GJ6j6
EmcogrQeVBxO/pxILhakPhyjlJEbR6ERoV44iGkjfaHdyVDnDXfm00mdHbF+e7wjeNYYEjKZrhC0
P69raNlmKCWNpOrqHP1qPkgBMcncnCnH9Y5sKfDxGUfo58DI41SboYtMIOdydwkP8aMifBTPbtT7
6X7EXVLjehT7+xa5D/vZe6+KYKqxbHOQEct3JEWbiMP91WDVrwdBQfVdOSWXelEvTPlVhEnFr86W
ktVYqZgHHU+26p9tqz3dIN9fB80n7vdBHilZYGqPGnOHHnWBAdQhUfyUWe5I7tR1pkzw+WuLOCZm
L9KrP19o++MHGyOS0hhFX0Goe1o1e2kMFwrq/EShf1BqaEBU0WU9+HjyAZLy6AWKmImF/efBa4UU
kk87F1ZZSn/kIHrO7mOv8V2VbwKqB1+iQLWoerIhsho/B+LxQJF7qQp7Akdk4OSUE9ipDAORv1zr
ktFBMpEHaMuFfY3Xx3Fnkbs9Ry1hpXyBeCAEsB2FplugOhWLrkSQU0dED43Bn6mrqTrXYcFo7epW
ap61lql/7UhnYQn0tJ9PU11uq1l6VHNu/yJsV2prS7Jh4bZjwNOduEmu9knpJ5E6Q2WT05f8sofq
DMbLlejroid7u8oZoglGF9hK1NluhBN7hrHUvwB6qTwzNMFm1+BLlBsf9zzyMBQox/pqGA4nO/c7
GLoZVH3+4EzW69fjiusHfZPSUrFTw1T9oIWTPC/fCMyLBIb410tnhPQoR6nKKFRVlhWC6uXOnmSy
EInlvbGO2Evxt2C+1/BdQJOTwkoJp+aUz37Rs1bu9Cii7RyYkSzoUDpc1VluYNbUCmZJioNreCE7
gNtLtBvtdNZ0sZmwxIhv6G8UvwELXNIVgSrZasgY6fJfTvLnGdtvESFMDLCqhsLJ3fYd8ix6pFsw
3NVt+ShNX9RVfX4=
`protect end_protected
