`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
lh80UAEZuWkA9hUkyl7K9Bo6+wf1XfXLytGUHygizlcRRqJJDUnelCmTpyQoZKEDd4Wax2jX6/ec
MBQUHUuHGlYZA+O2CIJC5zXWXxogluM44fT0JwJMFDHGakbbPFkS8Yzhub9aZOfxqJKb9AAI1gKp
Cx7cDQE9tauyoSYHiBi3e5xSBZFIW5mtyQWlKf1LXv6imABLNRJaSUOLNOYzKF5e3qi+QNxnuuWD
ZfGLSJeTyYG0auayoWD2hBIn0r2ENViUYvnibfU6mVHBa+vIICuKC9z1tLT+Xo7RzLLwx811ypKu
m/qT2YPnbuj83J2Yi09OeqtEvOxQGSj6eC4ikw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="mI6YLBbWPod3CAIdxBoedOoejgwwamseAIw7U2zpgDg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 94592)
`protect data_block
af6DLRl8rs9mlwqWPbXLqmifnDgWuFKNoqxSQkilBmKESiFttuYgMyw3pho2vO7FUS0EPngBg+BG
r6r8k+u0N5/QtZtdCHhR/bsFFEZ6NF1ERXDXnSslclMDPF2rhZPDH3r47lQTeuQVXkjABKLZujmv
lfmcym68C9cwdZ/gvfLAJUphVmmYL6csEIoIBa5otcSVy8AiiFKGu/XLvgLJhoPboAGwzKZKXTmY
GD3V9zLYg19bUPV2KygJLS805c33JotUCj5AHrxs16rUoCcPz8kL4sf1gHh9Tyf+ZommL9XUr+jS
mu+vA5u+KrV7Ej1DVpho3FtrhREDGLswE26hzXRxOMAYrgXrpQhohw+/9eME03SCVyP4TNXsVdk1
Qa9ADEslNHMEmMwtFjyhtnyE9d3Bdp4rNW6CrGOfr485JsC7CZLqR3b8EQOdmEKEsTPe9Kx67aqa
w+pWDOl8FvqjtZaILlvI3oSoqkCcQXuOmBQT3Wu04+n+hhmUehwrNDPpIuFkU2OUunI36aAwOk/U
knlwNDBaGWDUWlNfVdwFYSWMPxvutAY2Y9jrufl+Y1tRkIFUMGFUCbfn73AxahTHo3TZFPZLDN5x
QgSkqEvRuEfGFqrsQa/c/vTpJ2bEuDX8fRIxvMjHH+F/1xaoddKyxk4C0KBuQm/JCxmOH2fn7PYT
tDecGQNF4N0aTzyEResZPQmTdXRM4+6g9jUiCNMICpvPBn5QHzwc7yx7GyKDk0B7dLIrj2cpf34K
j+pjptVa+fH5PvSS++fLMtkXHGJk3cxuu3z2iRljmE4agD+D+YG1WLMxztGUP6k/LhYeH9zJqZCM
3Mk638fYIbC8cBgcccflHImOqFtYa28cZoezZ2pTWLfnVvXa5YuGiCdV7WVq0NZUQNikmOoEXsMX
bDDYdDwRp3mM3rknzvx9vnHNFzfou3kVzjKBMCzISPjKkm50RSI+u+9FfLZZOmx4h27JhFxaX9U0
fMOWxPlxSWbCLLSRR2ujivp1kaPDE88mBHvO/RIUoNdz6LmhXBfKRD48sXZ5rnveaHHt3Apk/cBu
R7u4xKR4ywaPjEnToybbOibBZ1FlH8gl5p2mZRuGW1y9RbDOAOqxNBF6HfJv9XKrJ0sBvBnpxuC+
JXBBsBvTQjHMZrKZVWgEsUki14nv4RFbqkG52JV0yYtgOkpbqK20V3UOwTDh+yopEzj4sKRRg9FZ
1ILh+uvE3V+4QSKKJdjAk7++xZsJAR+8YMmG8YZF8QRj4VNWW3uf37tgo7A+bx6VhWVahCyio2nn
BPktCE1f6QocWv8JO7ykII24wAfHOgpygaj+zPn0+LCWhL5dV8N6FSGQRlANZq+T0uBtAcEK2ss1
vdRrjrOJW4SPyVyUdLROxtUG2Frruq/kfUQc4QU43ia1rrnO6HkUDjBHK+hxpJkBgM0pssHrIYh0
B5fSYqm8ERiPXcvMQPLwgogIEFgN3qiJoDayUMX8aeUcQeNwxE2cfyOfF7T/hTtQXol0pJReIz2Z
oMoBPlhcWTJiwJPWsgUQ7edlsHE7zNGsi1iPY8nntg54T0dNhNGlE4k9FVKVGFAWqln4O7JrCr87
gTC8ryFWcqQmOnfj31HBR4WU8SKT9N/T3wbH8+8tM9RhN0ffII/mKF0LshecpV4EiWJAEYXdcmHB
TDvg6plsRpdPSzg9/fZ5om3dDNQCVEI3xWGtuBQumo22sSZ2V4qEJmdixQxGeRxSVZ8BFy05v16F
QTa6OiVAcsn5s5HOt10YtNP2agzUIOuvuqVViHPLxpIrm49NHi6zUeAXuJ8Bwd7N5JyaJeLYvN0E
itVgI9xQCQhknsANznZiUE5a8FsubFZ/41ZYyVPPYwSBTvZ2D5c8QATa1CNI854u7Ss+HDag8/KQ
ejJ38U5K/J319MNREo2wRZzV30+6LGE4HFs3W2kyZjtu+4PC6kQJG9Fk1HThBvSWNzbFUyRIfzjK
pWSaYK86xv0tbWcfAKQ/rETSJ0JbNuv2rBwesVd7VDAwJ4obHk0ppNf2zmzV4F1P0+XLTeeZcGJu
gu8qzpLZMaT3mRL4vFXxk07hAD2/73FOwU2L6DN+kKdkbWntBfmIORoBcoaWl98FUv8s4/sSQyMb
ccBwUiLJSn35ADfSWlhvN8zaZEL/qU3eIGPOBngOJNVcfczcEs8oF3BmuW9Afvdd0EgCZfpK4Ytd
06Al8PFYNe3d8OApyZYDRodUlersIpLQ+0EDEyBbfCsGCiXKTGxypgxR6Ofkhw/jZkM1OKyxIsNR
/s5Qhntw8XeAnP+aIby3W4Up+JlJNGxhcagSLH5ZMuYOkvq7C9f0PLgBbSpQOyKAIBOw5DzK7q5w
DgrpHwOcb/Jcxz70TALl9ZL12QQ3uxE5axlBVsqGQviZpgwPNxJCxecIYDxat4zO4y0PGW9DpKYb
NtnpMX1V/msGY0hMEIPInfJNoYo2gQNCp+Rj+mGZDNSMUXxyu0PDmHdP3Luo9Odq1hoVOS+SPgz1
KcRMwSWIrQ8PdQdT36sGRXCMzD6Wra47Rl+xtpsboG9Bg7VpsvVJVWdCUNyFD8NpFPRxLvW9bbKp
ZeR8uc1+Cle7jtwFerCoVo9BsSHHFOQ+1B5brA2+0KMN9wk72f1i+cZwaa3oATHzxlC0EEYJpjfQ
ohC75UG8O4zxK46V/Iyne/TJh45pGZNIw3VsrDINZcjyNW6SgP/TAmpRCjaocWY9It+x9SpJ6W4E
PosD2Q7FlY8yLb0tHwbahPTjtp/uv/0iXZ06ob64/JChsnKSTsuynfiEYzwSniCnJt6UM77oTYFd
qxyLd9gWsYVcnL2vRElghA5AqzcwtleyJwnE8R4YxhHAd5TwOZVIibe7BuBNWdRdK4vy4I9M/4wR
eVhI0FLqyLZjRA4pg8yvyxmb4FxIHi1d1ovvghBLrDjKJuOjtKmtrYO+U1SPzKvQRTeDibjbnnWi
gdnb3wkuQTOpfzVmJd/Y/5e0GLRftV0aGVVinkFuHh9ssId2ZFD+MsfGSs9X6xaLYyarfzY+55Y0
LsSbLZRMiS6mt0oM59brAqBNHDDwZPkRZvmK1rIbacFBteMs+E3dsBirXp9/3KRRHPIrHBbLuGgd
Nz+sL1lRKbvO1wOkjGbym1mJsENJ6ZMoOcgf9NBTjZS10uhLqkUCReEzTHcIXp1wTyoPqg1lBiF8
3U2caySRM8ZR0oQlgPXhVQ0JAyHy2AzDzFUAHMC+FAtnnZScD3sDLAT0lhn6TUi93o4tYMv369Hg
3Tl8p1jrN3lzUET2SxXNw8cWiAkUBtVplehhgbSAVSFRxkMEVmQnCmyu5dnwTjYlgE1zFxnUd0V/
plf3Oq5+GDUQgaL8ONAQ86qkvcWTj9jsVR6j/gpShkQwLYJ8vEaHO6I9iLU1miOpJ5HOJXL0Ek5i
aXVZqhIedIKXOWNXfW3f4TeMo6A5QiZxEGdNEkwAJIKEZqE6+3JZW6DEy2tDXCrPhBVAxODdaVcI
LsEXC3vQjmDKW2yPstEBDIxikMoY+CCfELTE4VBOkhPNS3i9Pj/EDwvjSxcgGtJ1zSk3S3Fr+XCs
CFafYAr5+ZFKnfNBAAVENDAEF7Sh3CT9vpI81P/i7EjPpoHTrzxw+3F5rJ3+PVqap/2e5vvxg5A7
ytHC3IoSvJeJQlkqCvAn8PW/QG3hhJZ8KxbEjBiCIPCuNXONxC8c2cfOLG8btefPo7Us2P0dDJ99
TvNjIhiwIxwlExY77Qxg+INwxMn59Dy4WZHGMSn9E9CJWQ1EHc+BvxXMe8aC6EJ8WKLidYHD6RwY
TuT7DOL9DUvRv6uSJTTZ5lecT4bumU3i7aljlL6MGBt69PE+qatigAVDbTGTPs6JD9EGD0vNdi/w
Go2rfefVPxHDSMLKQYO/4zgKQiy21kzYLygIkvUFv3chPHovtNL9OiygbfkQ5bLCrT8RIh6r9Yee
ECBUeZ6swQiqFwOOza5z//EMNLCPv+qzDu6Gz2yM5HG6MRTZlbvV4UWKh2hDyYvs64dwxCwEAF6b
NxWLVa5enDzzv4wMehCjL94LU0YEZ/vbuFSQAeRpiD3sl80gXl+AtQQ2WHxXh68PErZnUUIXazxY
7za8WgyPMBct3b9qs0jf4f1CqySWQjMi4AgO+tgkTtoTEo6tT0ABDrABnRlNKhjpj9RRB40/MKlR
5rOoYm1cYNgaxHC1qzdhctBkjyWXBWgmnmq4gWHMOUYJzLg/605MB2NmBvzqtwWnJ7I7tOdhr41Q
sLi15eqbIk/bNeHpfixPajVvUj9KvcTU41skUbQ1rlc+CDIehgkIEH7ZVUkKWNepNwzYGv6Ruc4d
M9fqms8B/AjVamiCg/J+8qXrNzPSIbc6XfIgMN18qfYaX7R2zl6aTs5db1wFxbUopJWnBWStFlOq
W1GjDem2yPQPcB+p3M6zKCzHUFsrTZDDLJ1vFsTzoMPtRvBxXbG21s0U/X0t8TlMiK5hBkReMZUA
zeYehqrj/rENrsTNTTeiSSdqnagUA8aEabWllHN4lEV648m0o3kNCfaO/+yJVXUwwBUp1nPPY/vt
sHf/OulnxyjAvf2Z1pw7MkPTZQNEmAg/MazTtdtviXKIRGjUve6uA+DuN8LXCynHQIXlnKqw4RQ4
a/cG9D11zOsEXQeRMpV8U6JFEe95hDOk4fR6ShExX6wNBq7dfXUBhwZ3S4qGREt7jmOjCtNkMnP8
2JIikGbWrUc7iBRDwWUbQEhUxRQxBDt950IBGNHNb/kVQd3/BmT5Y+POrxCinFWdMHDNC8bDz6LM
+EPCzE+Qss2iJT6DhkybIandVGzsGnsZhL6VhQU4IlEBwW7q+pqyxD/0NpW3nh/vNDV+YCxasJEQ
IymOqumqllqYoxJmDseIQkzMA3APUCSZ18XT0jfaGPYEmowQRwFOletLKGqkDCf5jL0ncBcbRwdI
ca8Y0jhLGxCboS/HhilnrlikFuAXn2rbCs6Q5kTOZvOSw8iWpVOxJDtI+n2K0m4oADm55CbFE0h3
4iKSwj07wr6WGatIpNcnwDhBu6qaFB86HnwoBHoz/xPtqt3BvhA2MDIARDHhLjzRMugfPkrYD9xr
A/x9uDf/t2K7RvTUkKQAe5Drm+Pr+mvbLWd2yE5nDsN8+viRwq8iApWXCLrmlhEHR778XddhysFT
3fE6Ff5777tSPOBGE5g3VF+etSamY6pm300SeCRP6OZGwhATsk6wtVbFAetTNibGIK3AHvyvgU5w
Bx4QXRQAou5XkWvrFtXZahv9NxcG1HaGuyij4IzmLNdDjhgB505Y7hwwmjonL9f0JpGsLkPCo+hb
q9yGh+DU9v8jsspuQSHDR++lsHPGXsk9CorWWl92Y/3e0Xr+7CoKZAQ1Tqvh537PbY3ZX1orOY0i
tKGIcTsl/DnkWKlX/uiT4j8iFCQUlO2GVQP6kBmw9hnIrIxh7rQC2SgoKQyEDubORklRPJ8fbkWx
BinpCWtGZGP1O1KsawpfyEXOWU/L+q6hCXwFa4H1J7DyzXiTXTqugwItoTdEqlGA/yfwIVi28+vh
E78O/6PYMkkVoRHrTsoRy6RjJ7tCpMz4tu9UA/o0mSqNFKW8f5cYVae3uxG6H9IZvqAmWKjkIfKJ
bA4zEK9+FhHNRP9s1NChJWBnSjL/3HzRSQfLePAsQMuv4Cm8MtA4+66TPFawZoWpUgYbQyHa0/jA
e/9dGdxVDCpWP2T9ejak8DC43Fq2mSE36td7HSf0yFas9dyGwXznJGv3bDg/Qx1oyimyjs2EvgJg
OlaSoKzzdj7cFgMLsT4Jg/hIlo7fPH74WAtmP5D4ATgFadQkrhlpa0V5RFH69zVHX13otrPjnT3n
dt6zkHPfef60+pW4Zvgkm2sjdRw5qCRFcq8sf8l64DlPbY6WHEKtZhfI3KpgnsBWJh52Edj8MtQR
8ZuO+aryI9IevJ+qqqewH0+yGV3FLvxSAdThrW4OQrCTNN27R0PU0AAOnwgItDwWeeqZbCIY5u2D
SvBprzX0e47B0bO6DIQmLF30SO+dCo0y8FNRVIfN2fMN8uhzGFo0kX6tDm+ywwQw2vXbwSlLedtD
x3CfOZ8NK4MWAQ6wqsPPDkSrE12TH1fV4T30SBoEEU9a5X1/evmB0A/KR+/7mlj53aXlZdS2OslE
Iz0eb+AYCLb1W8qLl2vm4vYVUX3/MUw2sWRQ972kb0+8yVC2PTrVmx+davWaZp/eLMqNrJZ3bw0o
6Wr+rU72iTPFmZAZfHN4ITNfoq6bFgSDkjuw/Rsso3LqJlJfWrLsntTWRgBBEZXY6SMaHnYWD/SA
LcPjL6ni75XwuzrOQuRYVpCj7Jjkzxd097agYFBPwwDlRlkgxNlnOV8sTBpmX2pcZT1UUM+wCIHA
ltm/0T/xRSorMHc2c0Ox4lw/anbo7bOtXaBM8ty+qMbNmzBVCcyEgr2Ux5FYWWGwTPqFOhN01ZqN
neHOWEp0nH9zufzXq6XteOA47leHmm5fUjJBH76oVqYWBWNZakorzEsENxG88noTA3X9C60XlneQ
ZQhu/tyvyEgRC7eWbSsNACcSH8wfYKy/cCNAJbrf/WvZBpVr80kRlnuDLWA0tFP2NUCd4Rjolvpv
10ar64kaTjuQKSOua/Vdp0Mg2WgSZPmJ/AZDIey/q2t1VVWwjLfjQD0wKj3kaKs1+TpsHGckwIgx
+dJKlgnEi/0DPqNMH2gSVIuw2gn3jbYexiRwvrGg72p/GiwKqqG7E3pzdLc/V58L9Zi6u4HSJeql
uxIUZy+5Gsn83TeUsDW/92vj3Mln2SM162qL+71phzFfpTPl4JrA51ipvkDUt+WFCc/jQQgrJlIH
WvOFYazAycdYuPiamAOaPZwe8EagZwEPDVfEbB5zeLf8SJ/o3ujFBvSOjUkcV4XgkbBD7F25wGgt
0dPbp5Wbi/ongDEbqqls6kCbZSaCjc1KsgHPDHxVHj49+PLR99dGeI0Q64MHJhSxgxozyGzPvjkf
W1zP5DJJrIj5/0qLSQmNwk0hrEsneCaQ69oEkR/yo4hwZy6R3O7+vZmk7ypOM1DSsG+2fGAvVsEE
ziImufyGRqTSS3RXgsPdcKCKAUiJbuwfEDAEJIS21dlzysX8e2wyI68J2x4Qblz9cV/G/fKiqaPS
cKbpdL1fNW/JrehzJ5LRYRutGtmYE8f7xcdIe14I2P0SCYRjrusB1wZwhTaWSW6hIzw205Y1yyvl
++xW/UpW9aJhMCWfqN2ScHcaBneGSPSqWCG/1wCq4VUNWOFPlRMo13jbFxT0kBcoucCdsqkBwXaR
ZF+wgbZlw5OGe6dFX0YLi2VEUQPpDToul9f/yAWuXNvBJFH+71lZwchTItZXZVldel7YZfiaBwvr
YXVm7MuJgVHGnV/0oj3Y0xxaeAW78eizLgxtB++k/i6hbNpKQdshwr7RmZU66qPELSoWcWZ7syoa
vPH50gZOuMscHvP8QwWuZTFFHpB+W+S3ueWKY0igcdV22SQLgF7MM48XnnTUpaIZUGhRxqSrn/jY
z23aGIxSdj0KgLNh00wAY7JW0NrX95Q32q2MNKQ94yUFAbO7SiPY2Er422ns+b+MBQjcqpOK3YPm
tuPNTcLOQ+2wMi8dFY01je/gUtk7nXLleMODiMfZVEVpAqYUMGECgmtUzPQ+l5QSOQ8l9ZIUt1Zv
VyeXyHz+GVsdf16nHqVkNBzWn0dzA9wjPFkymrVLqp3r5B1Y4OyJVTBU0RYLeYdDotnsBUUKp2uW
LiwJm/pJt9+qcW6vO/t787n+9MrFsyeNcRHDKNst10Rk7obP2oMfPoZ+EnjvettGfpDB7oYwJgHu
GvwsDBTdyomKcPQVZrNXsWzmbwD8zocC/rF6MU/IjSz9xc3nDSGivOnl5KDAETlOggf9wG7M1acT
Rx69L5Xa3vjJUC/FparHMj7X2YLcVJff3BkU2EImGCCvSjbx+Lbh7A8kE+/4xCYT9En6fZ5oM7yd
s/NzpgSGgahAhU+vW2sjJQmfVHtEhHyJeSt0L25zlfyVyCxe0E5nVMat+mlxTmocWnZntYTemRxy
O87Baxh6cUbliHXUIqYjuZ5joy2CESomgnj47+9YYZ+PzhEbP1WVaNZre7P3IDzQWF1HOVKYc4Wk
7l+XNihiRHECCsAnIveffTflbF2XiKbAHEjY+1kRJjvk0/arXvSIPwleuWVSSglgeHDw97ZeXInq
UjcBszU5dsLfugWcojfBU5uLSrGDNpbxf7y1OIRWwJhSryQliXM/O0iPzb56o4+rzaE+qv/AyQkn
nw0qcUFw1oF+aEKro5RP+HPXmzfiqEtiyt5lYV1SD7ylW7LJxWZomaOa/tBI88xcoMjWD7G+acOM
vejYpEMBFOoWICJ7B9Gg974vJNCDwf7WvoQF480uqs6ARTfboFBDzSQH3JJLc12SO/GfMFwitQZ9
zoQfJg1SRvk/fUmAon0YcqeiszqvvDZ5xulFrVao2KWEEvzH+U8u8CgW6JjShamxz4h9NqZOuGWq
Q7qVJxY0G6pi4p7UlbUFeDEHJcsJWRHS0a32tEUv6j154fKfKrGixD1B2cdY8re1MgpyM3JFtOs/
/G2NU2WYV/UaWnGASH+7ynV1VE0NBsLgg0OGxCuRfR3q7Xsr/4S9Orr38t+mWhFwjIJcbizS0jUp
3wao+QEB+QXSacWVd3kUZpCX7oEy8s+iHmMhL4GQV/uRra+q1RVmW+gaaZoIALZJUbS4khAzfogI
F2kcDhf6ofyX2V9xb/RpUA0G+BI6t0mxbS5FvGlb6izojWpMvecgzRYtE7hcxdMEtiebyTAhC1Ju
vnJQq/wQ0DoHkc2To9GhdwDOD1ZFP92OC+CY4QH+r5EtAmf8pmmu0aSwlSsv91gZeV+79o+9ZKRV
8+Utr63LDnWsSSNJAcVGGjU/375E2ilO5jcb8kLDhx9Nkv+wyMXVoHrFCFki7HwWvDVVQI684qbX
D6m6eAubQ3M+cC7sdHB3MSU+9ISnLHilEDmFkonJ09Ak4XD7+aOIMMxF18xXaoarYUbFHf1yTw64
lWpCCizvyGrfJeBAK20/MOelnjyJmfrgXSGyJkfsuWR2zYskqTiaz5YBcaOQTVas9m0mCAh4jqWf
l9pf2nqsbstQmpyqDuLjq6wTsnv/ATUUw0WjIq//cZeW6TAn4umjQL25LYWJhaF5dqN087m2QO+p
cXoS01kMv/5/bR6NBD2Z+y6//gJJt3eefhf3nVdfLgGPJ2v2UoA7yILmLMhFR8Mvd4X/k7Tksxks
PYOOalBCurTdOoG9J7Y7xg0U2bn3X2Edxw83kfdXZtWAFxgZrqeYu24hQZLq+a+HAK+qbk6b60wt
y25oR7gJp2Z0xUo0dEc4K4SxfulJpCG5oCen7DbwMiIlquHKVPDV9A8A8GhmBJ0Ufb3TtWqHqT9/
poX1HcJhz396T9dKeBdUTk2UYlcyXwmbInm35CiyrOXofJb1PsmMoqzvVWJoM5tKEX/WmW2Zzffp
Y9iFf5naf1Jirny+KAt+ZgYVfBWuJDxxXmysKikbnGV1vTr0wqAh1f570QbJGn1lim+W1SaXDq3z
SuNTPWJDsYx5K6QoIMog0Zk4lv3b0sAXDV0ipPNSy+f0InRHhlMSFj7oBks4hjW9EITCCN6sPvNe
ym8V6+IKHfiIVMbyQUdFDN6GLznLdMEJL0gukCC0gYJVo0R5DN8umHzZuWstfmdDUZvYsHvBusyA
Jia5RV6MJgSmE2TvKGX2qrnzLb0E1Ka3yTB15ddYYjaNupOABKnBo0irP5br6QaDjpSaF2YVMPX/
oBBB3PeOd/SevRl+NZFq1wNPAAaSdCtXymvM0zylpctwmUSlcdn65XTuY0Zi339RjxxcqV88QZ5C
GGNzdf6ODfNhCZ6nqHuUf9BKBisgUgsy9kGAzlmCpMSFi7I75cctqU5ArYhgAR1GbutRaLF0NP/s
POuC3LeCo/73/OVvLhSazi8Q9OhuTRqg6x8PjypKHHPAkHN9vC2P9TVRFOb4UvYMT4xnTaiswPKr
ejvaXKpfCLfQvXoDpQQNkzT5Rg1pM96JhtnGNbMcFiXKkogDslxGOJ/yy8uaBqyYFqRL5TW4w2XC
/e34RRd+2KSnL3G3vEGbFJlsB7KSrZmE3ylCgnesu0BCawpXpZxyiDrajtHBssz1cZvxaDTe0OL4
2b/vWPw8s4/iDphd7HBwlng760zSE2lxHb1J67deL8KOAV+kz7jFtSbsHddUx4f1O1XC0tnAvuJD
jyzMh+ngir48eEqYfNdTphkoNwhNGzqopJL3b/2mAlRNQfxBAOfkedO49Wb7cNqRsmrcCbTWdQLa
OPzdO7fdyH33ucqQPYHVo1oYopr6dJGhnlzIP6M/BJ408ZEhbLGWnv+nDJDL32ilHIx0X/+PtrK1
ZlO9kQ9JCPftKGnnrJf5+yKxE0nXO6I5yct0ZvLSdqn1UR9p0eJjlGeqVxgLBjAafhRDSRQe12u6
gmQF2XOuhtX34u5dYJ2p4YwMTcvr33Bf6l19k5CX6im7D632HqcixU7evsKrhw8Lj9tzAzWtdK73
5FaGF51Nc2onUovbCJGT3MHz5DcMRaQFASARG61YXt5EWY5scybC+TnwR+IajJm9MscsRUFBdCEh
L8YVbtj+Xwp6Fp7IVHsLCu5r8AZqdiKvyEC5iKDIyWIJUmLQZyHXefjsQI+His66HkctppNqFH63
8t3UT3JgM2xhHsrS8kzEIlvN2FCSaljfQZBANmzYju5/xboroG27G7WoOcoIqvqyWxQeFv3R5URb
g9Y7ZdlQM81st8908Vd63brH0Ie2lcNjrJ6Fdxem3D50Qsoq5H3hxVJFtt8cD4wzBKubnhU1v/DD
Q8M1XAQyycNHFpB0j4Z6y49A65pBcb8+khLelpMXzDZs5XBm8UE8CLSEkURjIqasT4kkk3eXbifa
meHOGOfRDgisViiRYEOtB1FxNLeZ6LF9cS0QCyW5fG0UwObwpY4clZde8Yjfz8kNq/OkLesmR4df
ZqHrR0o8kGPbZO5mgQD29Hx2CSCS97xp3ytUZQoMTC3jsaw3OMbD5MiKqL1qGLbrdtFvWzMKO7p2
VVWZXWSMgXRQqEM9UktKV3CncJIhoUehKNeK+VX8kxeRaz74nMmPnCjHteEWQ+X/AaD8zUsgt5jv
PnAAfLDI01MNx5371E+B+sxmqoKMhbxw+RwoZw+3yPDnFqCrm6GZGV88OC38IUlE9cPsSdzwrwcG
+qgVvZyPqg2NXgO5JyMQpBPsM/YKY97zXhTZyjhkm0+uiiWEhDT5UjZsdBUvQGr0Bl5msa579nmN
4GQsgu751e6qKTBIH7Sok6Hkt7mUscyedrwoQjymUmaJ4las8L/2tZhARNOF68K3ZrYQxXd7qxl0
S4k7TBp/lRw191mjy4cCJpL+b3b+TNxe6RD7uPhPaG4DLCOmAXzKy3IZCVlqM98UU60v51x7kAqV
+ii0NsGrmmzYhfn7fVAbp39OUqtO8nuqvnx5Cy3+miwSycMSlLJJfROnCvc/SnxojGtUcvg91xx7
B4JsWg3WfsWcoHvDLG/SB3Rb9VBkwjEA7Am2p5FltGy/8u8VvQk9T5QWaSroLNAN36Wb3zuIhiVZ
MnDsjxfZqanp/0t7TRJ88dy3ikSTWqk/7oMutFFqA9rQDFReA0EHMR4S96ovQS6J8ich0y9yv9J3
uOXWOalQn8GRfMimapEpIDyTeuJfIdUBg5mlu+mqdTtY1J2V/L5u3puQHkDVv+5D2bsj0TXfCJZ0
eLpvnemYo/xZ6Cgbwwbj7LizEJIWG5KrPUnFLZVpPwH9xvOZLvf6/6Lkhzmxuu+PzNI1XHZ9gx/I
MK33jlv3Xn+0jPdCO6aXiKidQp9yubukWEtyRaN4iOOboRilzQ3ssGwndsPVXJPITbVBQdbmGWX0
ekJn0iFCMWbm1AK0gpCcvb/Vtt1nWiSbnO3huzdNj/pdRvGuMvoP924mkt8a38/TYFNAgWR2nGV6
TUqE/FT76EQwfGyfJDRWelLM+I0ycr5TlJfa8wSZczbgCPOdTSvYca3ngyF8s0R4/e22Ksb+U0Ht
5zT5f5ucyUjU6dUzMGXcpZPK5JUlxh9kMUOpmT12oPwNSjsnFGFq9eCs5Q0t/p1RRfT3u81Zt1ov
1/PukXDWaJeGyY4bwxyjEWiGhRE89wuZHv0/msNYgoNdJeQJag3VcOqgmcrVNnZpQep1ctf8p83l
Et0+QcxuQ2H0KCY6mVjG6H4Y+bMyf2MMMHZKBgq584tSdvEJ9FBYykrsO38Ng3nkkVmPR8GinsI6
rOg9+cU8FMDGk3//N249ceRwJq/denN0gEcfSBaqeJxNLKWGlr9wpCZxdiHmEL7VVr48UtLGsoxL
rjOVGDL0Z/tIcUa/X0pwodXOsEpce8wLudq/w26RAaG3TUwGeZoogJqHSiwuwEzy/t2eorn47sW7
+THfTywmoRH1oHcAYfauRrqXOMgedKZA/xXNVvNvDruuZuuNXxtupgnLFekOxiGLeBgEEh2puHTS
ObrSIHERhaUM/4PQn6qPFE65Lo4Y8bjVC9eTlCaB450bikgjNG7Pz/Mc6EGKy0qkCxO6QEWGHTDN
2OMDOBhpVJi1uRfRTDnM+LhRO7rNXCxEj6bEDsARtFvmdBXjslV+pCmYpYM+ynLwG2/Ldtqf6kJC
eBZ8YIFxZFv1sT0aYBJgQl5AiGBOVjWMwCbViXugD9phlKoLTnWk+Yu0h6KIx0oAY2PTvRRac9bl
/dsFI4FD0k+aJdO2eevYMOoDD4Au5yqkNeApYcIHnIx3UpfPrvIv8k+tHzvy+nRbP+ObMtrVAA5Y
ky9m+hu9D8AjDCILxtHzANV20GSnkU/VomI02TncPQiIFPfhk/2dpF70+Mc2aAZl9oSmEATurfBz
JqPMi78Vtx8vq9C6E/RgxhLaPtVdrN+qkvza14f1GDORd2PLZ/zyS1vNGKvqhz1eYplJSONfe1bX
A7umBmvY6pg6h1aL6gZiwZU4rRE7SVhbXpdmkcZhg3JZwl7IFK3dKr3m0OVm6yeJnt01zxLvPipv
xZcrFuJMWm3KiiryIABEpbDf/jxPicq2wXRYi9OW8DDZR03bj4lkqN2mCScDbUQW70XYFrAAdU11
CK8aLJvtLnme3cvk7x+SXfTgYDVIRULepS0a4xQLbq19VQm1YMHzcytJ5OJqaXpnFUn442yL0x6c
yAAdV11X2ZXJCvKB9k9sS857GbvrqfbEPCDriLsUAjQ33M5RtMzxlY9NByWSv12tYMisenR8lT0o
FSy3huve5AFaUOXcry0al5432kz61W4D4M+wjNNPNdm4fyIFOAtCWv13VlvHZi+W8274CFC+QWes
SVfJj3KQL5Y/bkK+JXzJOKBjvvhMiazjdpRbEvWMjLM3n+D8caor9vZ9vs+oe9Vsr2ljLBtcgj8T
IJVRrN6JqrqC7cIHIV7DiQeRBkK1K3SOfWggOW2NIcnzZ7oUQMFjD52dUP+X+0EgEbLkRDiHVCG6
6kNEemeHdo0qOqca9krEHobpTgmNB0O1gbuE1WuZAj+TKKQakpJZPq2VJc97Nf7rPLeI6DM7lqYr
591u6YqaXtKy/hGoiiRSZaYNqXscgvjM3ZNY9qofQFTLxGVsj5BScomxXKb//4W9apbhs75XWut4
UNNQHjhc8sp1UKiWxIAdDJVParOm6KdUEcBZgSm880y63cpferszTXeo2pvORes1VOHXLV+ip7Fo
qOX4f9V7CyMMSxtKjR+H99vClUWHhOcL2yf2WFaL+2vLJ2gv5GORVNZEZfvGr7GQ3l3Co3D4fGSx
dq0lWu77OsEPXkCiotEvG/J8u7yD64K/jMbZIuThSIkXB0eZjHYRf11Q+3ka3WMnovtLddEEc7rX
N4WqW30bpFFK3dgWtnOWXcvpeqk2EkObOY2Muz9M9qo2Wb/sHeLOTb67T6Nt4o3P9Xg5lfe2E2qu
rTe0sl5+4x2rr60YYxPaYb6kyxfTlWmKz+kVzuGeeblkL33BiNqTa8Pkk7qKSpCANvt7GvAxxYBJ
JvPmvltjHHjZBCcGQ+R1TtaJ4mQgvNylcANk6DeCNjNyRrB6Rf03n41nKuT7xg1y++mc2aSbX4DN
ZlVPVYkXzZKJ8olNawre5MuoGa++vcEGETEWy1PBFbkTJl9Pil/EE6MIpg7a1jIGtawyh8U9chHw
2awVM69e9R4nb+rqT3UPa1drZGMQRHiRrr/vTnXWwzFLm7GzCM/i/G/gH9TT1Ow/cTUb1tVVmJe1
EDdpAXlEYSL3FX7I65D3llRrKCVoDt3iiUrvSOMiIzLPtwud0bE+B4MNK+poGlGQ4zoZVomqevq1
g5Bygyeojy0gKyoXDX6cC8QgVzP+Dq8Pr5GgCPrJCyiwfObP4vYglfPS9cJQlH/Un8THpfj4TKQ2
1ykCNizlsIepSf3VDJBMBkSanr84enhiah8TvQKh3pDfE2zs/4nqaAdw0WSSzcPUqojeimRz6hQO
TltjUTFjyuKB3YJ9bUpN3w9b9jDGgyBRIMa/jX9cC6a2Sr6Le1a45mxNczFRUSrvQK4vp9xsZYpZ
DVOqvg8qRVvuOb2oZgeXU4OIryk2DuydxLUJO8GGuzanz52iSwzXXQB7k7C0rVIZyY3MQPMPTBtF
IBouaRjbxt2SB0eMFCec8waGYzAesrcAK6fzN/NBrp+soPtY0ZIeZQnWz5FJh+/6e2K8fLWTXX2U
C1yKvHShcN7P9yM5upZyFtlzBib+TF9AdWWi6YHxubcNF6I/Lc6IVJdoy1KW8RoDK7Skjo5+sG52
jt8Q4oxBwEBoKfxaBOUoG3AEuPwo5f72fMRzpdBdLSBfyuErFlkoUiEM7g5Yj2PYv0Feua+vK5uO
Ed++xNZR4E3Sxr/ZE+Z8aJh+0+ydGx9M+pqWvIgH6IeihfHsaEdrBtAGpiHH7BycS9101H3YMkKQ
k2v3gl4ccGkq45lvc+2Hmbz1o4/22WA+P05u8+a+Hs+knlQ3aseK4XLXgI2BMnv0hD617jjb6Ns2
Szx9FfoeJtkCMCEgfqo35eLF92M35fQt7hhDYhxX/tCZipGElMRY92TLO4nTRw6rtDuFYrQMuIxq
sYXn/BcUYqdjIkWx6j8L2K8DKolXRx4B9WF0VssaRqWFDj9dllQzqWod9R8fpPJ4TrKLdAzG27gD
KAzXwkdkcqQxxlZrtNT7YOT/hVJXKEswRE9I4nT9KAuArI5Ix8rnRuv8NO7FtyQZ4bmQjsRA9vVT
7lMh+guB5UJO7q5kqQB9u75WFEnbcACGlxAzSX1owdKHunwcpyCl/9wLy+wyHAV/nBhdJ/C186Es
qo6Nkri1nvzC+smBqInK0Q4Cs8zLjEejo7hy0Z+nnCIwUo1+GOSg5SEqGMYPkzWKhZ6MtoLLnQtc
AdUe5A5lkS7DIxJ884a5P7AgWtB0xea4KrRbAY0uYSq8TBIgc4lkGNsdrAdCuX29k5KOQCxPBQLQ
NLM3cd29qqkxrD+S3YuJBLFFUrKiqQSUl5BF6J1oTU44xfufl6imiEPcryxlTvJA+E7JsU+crecZ
kdu077+WdVtjp6QgD9V2/DH5tf5yZR6xZuRJ04+xTJBXEvyG7zFE3hTYHqZjSBGI4zqRzmRm0uSs
XGLpWByK1Cnl/7K09tjjgrf+/UsYzSR1PwO7S98vQd9EwOKKV6We93+QzZ7e0bd+u12j/NGusJKU
l+r4kimylbyvVFx1vnnEcWvlaNS0LLNVaN7kxceOyhBrULYL5Z4+TsT0aLlP5sdRuTvo7UEIX5Vz
zExRR+85hWZgArb7QgqahAHcdo8/yW/Q2tWyd4XfcEGku8yQOMTafiEWRIHxrsFUcC65KT5e/2Ck
VIDk8TU1h1QDABo6XsmoUKsyyuByuFX0D4cL5PcRARrPyGFvGfMFl5aatLPLBhYzKGsMyDfdIlLW
BZZ03VpnUJjNfW6bAwXONKQZE9c9fQE9dNIGpyT5v4kUAF1Kskz+DxNfbozbrwTEnBduU7T1gg1t
s7/tGtcgD8PEd52K2vG/5g6+WUROFgc7fbybmwn0HrpOSMrRvLjO1gTZBGLkR6a+czeBQgpcIbHM
4gmnR2dik/j+hWC4KzPITOYuX2PmREBkup8ofh9xurxqIEuBV6FpKwwPbQXtdzEKuXW1RZ5L9JaJ
t/CnxuKOh6nWAsKl4fn3Oj1mt8fhl6e2KRo/5NTGJ+mEl1uBCTlCJwlC+ndxLFZg2aY5lqhNRBQR
kNlpuWdUa0tXwUk/4tijrkVbe+Qhi+Y2BJVYQOWy9NvMItubR0kdjDu92MqKnuXk04QCbLlE8Obs
gwwdeQfPV7shIebRbChloQcuzhQ8QIu339lam8ONPW4dOnz8h5NTBIeiklN56uCQV68qvwr/N6eI
s9nWXa44PjRyouD+BM99SMxBE9RlmYK7GuUosyF6u13rcABeGz+XrCQRzfs6+87MwAc81JeTVeO4
O0QJhntftBMrRcim9eNW5bjU79qfW9l8Ven70DUPb7i5EUtv1cxxtRjbfAHEcESUO9dCaGKAIGUf
cx0+uGppxhXftRKC4ynrGieoup2tcpWZxJqIf+y+UVeWz3KajD2D+A9304snPPaIfmJwSTjig76b
n3cLWZ483Q/47XXeesNsc4I8If8NvcreG/QVh6RlBTvuK4etssVdesRwOwPYoS7PinXjXZ81LNyJ
bRnQCbyi5LyaBKMvllqBMHhWugECfewKnRZ/ASXYoJYbBZgcKT6/JVtHaEFYH53Z750XFk/TWG5G
0gNGAzeijJ7vu9HUaDijaerCxJNCbm6kjvLYzp2Uwr8w92RwV8Hdsm4ykNPeXafZ8NoiM+DsOo2z
MPimO5ODVYZbqoMjdg9+466M0wkDueLfVR5dF9/fOAe6gJt7yRGIk/EjU47dLBhPVEfD/hw2XOWC
pB6UWpWG1toIAVusgL/P4FnRu3AE0icudNaWM7CPS2RcxUL087ROa7gMQJ8zq1zHfpHVCRK8Djgk
Ii3NYWc8DVVKNLcc1wRXaaKnfaJDXAOuBAkWDvJkxh8E2TtEtHhpYDojaBAbhuJARrzM8XpveVjY
9VBcyMD4rl3DXPLYxMXpw5eL7zzy93BAMgMJKqqzVDcEnuFdpqvf+m8Sdl9cm54gEZu2Jg9g1QLV
aWoz1y0piSyOFYGQKWuBBvMsXYAPe8Fs18jW4/A7XeHqQITwOOUk5ctgDT5BtJSPVhieDx6zbOoW
ACTkLF2NZQ/GSOkvBE/XDuCa58qnNJIQIOyTRkuqDqi/0CbX407d1v6XiHA5+JD7q8QfE7H9zGNl
P/t5RkflKoTeqrTDJ5ni8xp0g2mna2M5RgmQ+nmhmVfAy399A5qy4xSbhzMdJCnJZ/s5r5wUMc3v
IelDWI6iKxkCMFelz8whA082mJRiNN79Bgr7PUqxZvxNZttMik1IZCwmZOGAyzVK3gKzK+wNZRS2
GhuqluEcKI1iZMdTuXyYw4JHX32FdptVRGC8eer10MfM9pFHMZZwjZyRx9WyklqvJGYZ1TxJignx
M9JrLr3r9BbMoKggjgrgqqJK7ezbIrZeGoWtfhxAVFk8bnzBApBM4Lfr0Cy6aEbL+zGmY69VRLYt
lWrGlb6l/rWuUH8bSqKMgymfXvRlJNGj9k9z6QmwOQuLus9Nqln+YwrJ+chP5onvlJL22pOm+ty7
Jv9W/Kbxk1r99y4ZWa8cOk92PGpBRhsTWBgM9/E+C0QSHbWLn7tqjdDtwpxJ72L5/uiMDfMJlXvo
QEkhWaduNMFWVXakG6sVjiiVEvQPP+c72f3e5Q/ws+y27zxEwWLrmVPRitXeHUFQOfIDMjPXvoiw
aSLnUnBoSTHdPgXXTI/2SY3BHP1ahBKfALVW+nub2mXzb5bXpOOI9UDZjVPLi9ymSygFJYD2IbXy
RQxDHIZjhqYhHCpA2eb6w3bsw8TW5SJeH4u0kjG8Gw00eVf0IM0Um3+C9XRaT9ONVmP2GHVrZSNS
AfXHRdXKLT+JyJ6h4hGbzwSvPCpLIsU5GnY4LJdO1A77I7KDeNKpgJFuulsTPDyyEiD7KXajA2Cj
EFwQDxFDLZjAXWcAay/2xr4QVtv1SOmNUILBYI/TCUAPr5IbomQsgdvxAtHoK0mf8O5nIV0/3vII
lbbVeiZVoTRb/nJPpdHdI1sjxkesCXEDO7UHkznSFgRRToaUoXly0iPy5G/+03CkjJXdAvc4LBen
nC6Mgbn76nQVDD9R8uLufswbT0GrkOQOvToqnwJueKj9NfeHB24s6OWHd02rp1iI//VWEcwqkhmo
Ue5pDlq05Ox1hUFwhT4On+HkWn5d0zEPIXcTZoV3FBHkaSbKLKPBAHKdc0Sgut34cb4rEqoxT5rt
0ndLPP/Mt75EP6OnppVXBy+yH0E36WAfj3q8llSwV+7+K0Is0SoofCuI6U5xRICeirwVHubh7Fpq
xhgy4cGVw2DOAegf7rhxrqyk7z+Q7mpQCi/p21fEkTwit8Qq3cEzCrDgjBCdpKszIUpPCjCE6ICA
7VX4TBNxWBc7eI6rBlsygTjUiw56WngGqoq8QTUzaMDwBZmmNlA6jW3RXy+MWPI7hc6K2HLVcvPP
95CJChzwoAGG1NpRZ8c0MKM0jYJBGa7kch/+TTeD8HF7IDK088Gw8SuwHLVHqhNQWox7XrR/maB3
05YtiZa1ZWG6T/eK8oboxzNlEVrdns9kfEGob3MQth8kkXGsoesmEm9e/lYBMsnKCDkDgcWC0yLc
ZrU9b07bvRdC+btAWbFl/HucGd8YOvJyvm81mufhshWCd7j9LHHpDBycOKCE35iSv6wuiQrNEvG3
n4+QKCOxLCVHYFaLYLWahkait2AVYdqCaLJhcbB3IlHViYSb0eFHuO4RSdL7BFFqUdq7WYsOId+A
pXAl58frZx40pJmr+9AP5v44yTULLjAdjF2iaojpCFJY8NcdnLOa4isIncUawyB7KkrmlN0N0ONc
S18HuppbTIAgr94HPhOGma41N5DCq+Wd3LJG7OeuvWNoLBm/kteMkl+MMNDD4L+SVl7SO+C6Hi3N
VfOoXNYg2Y5xZdzAotb2aNxF/0gwC2kTY5hfGaMgibq5C4GW7aQj8BmH6x2bexivWHXJSl2ymtDY
hYV7HWT4uzghpO4Yr4YW2v9PatocATw2tDdw0/wRENhj1qoQGQ0ebhqcJWfUnUpY8KnSFdiVzeQx
rRLd3zjgkALjhrnHiGk/2pgsaIbVQFbn2qRlVuD3zTojZwjsGMwGjS8psV28/IvtId8Ekt6YZCnS
cGjKUBiG+SeH1ErgUejL9bjvKuu3I995UwEK+f2gfK/mlyaVjtowSBmNX4a0jh2cSfwHght1zUxR
fTOF1Kynab8kUvPV/7t0jY0FQR/Ohcui20Dg1nUUY4oULkQmricNQZTVyJGzuwRiOsw5XsA2BEsr
g/IFqF1YJYADZ1Nwt3j8KZ/RPUgArMRzqcTKpX4FxxsHllWdhOTDJuwotx+bupSC+isJRnkReUbs
e7Fsqf6EUgOf3J1Ps1rlhVAb6LxnLG/C+HbTo6WVzyOvTF0Qj+No89lKv2x/MghfvocA65ZeTLZ1
GfD44qaMmGlqulXWJ2nbyrQ352wNPKXpLEDxHcfdcJvHJMa+kWAaVFSthUbOg9nNHNor3QV+0bTm
wY2kiso3z+3/ag02xYLPJJOoZGpfR36xMut/dPFZE5xSC6V09bsTfQqUD5QwOjC27uVqEK8+IuVq
RoX45IQanA7wZiSb19467qSONUBNLcuFV4xW0qieTyaOlelpq6v5NcBAvEjhJdy7B8NKxbU8XN57
DkAwngy23opxV0nOH21A98FEFxPMGShCATG9FjasQ39sd3BHR126MFkMSpMYHJ2TBdqrYXUNtezh
q7PyaCNJIgwZ5xbM00KCTPgLY8R9RvBR+xrkIeuTpwqnUORS9unneAPlKTfG8h6qfcAP7N0jkG4v
wMe/rC9OJxeRboVXLOZjUoo2gOWkq4ohpyA03Rofo5ZyNqNjrUhMlOqvFtym5LorrBSOIL948ws9
B1gurKzXWAr3WsboXF9EJnGNjXuK0WauOwYBvx254wVd/Km1Yr1dvG8oG0RxrToGVWCUm+SiE/Vi
+3mGjindoijene1nWamHBHAhCKbMhR2kzj0uhKoWA0V3CWNXTSLZL8byPs1ttd1+q7BYsPO8e1tv
dl/VKXXMTzr5LjsHRxLHCpvA7Fi8Qgco2kLH99agTChcDD+RkQWKeFI3VrRzfLcsZkogCKbMOnbZ
jtc6vKjL569Yd7YcHGI41rg2EXlKT02IDAVbqPGEoMOWNHKoFE7Bylo6i6G+vfKw5r84CP3hXeur
MqPxJbqlSgLpHToi8SlZ6FHxyuJimjfpNWqt9ImSS4jNIgsDtoQMIf26jCTlNELovDBSp0qgd5Vu
pYTccqI2UcVtaQTWXojWxcdyzn4Ls5qKitWw0ypVEHRgU5pJx4wD6Q4QaIxjCrH0O2vC7QeRWvSh
/1hFIdEGbJB7yMIDenEKuTqCDOaQ7umM2UBROh5uHvj25cLu8sXIwYYvBXUixQ1zQQLup2VGjeXZ
dFBMtSjvxwFQcLckQHRFGwcKCoF33VaKFIk5w033+71sP0sjTsrZ5H4Tcf7VZCXplVgFKtkKEHbD
WVGJBBr5GGYf/vesnc+Ujj/+j4Dv7vivuK0rfooKWY1/sohfTcdvLn3XMhpGNrRYXD0X+52upOWp
L/Q5GoVhY2ERNaGQg4yDRoiuA/bkqOVPx6fKrGHkIWLCyceMRe+QcDT6N8oA6vAj2JjEU/JB7+4R
JxGXgkYFQYqMThGqYDhgR4o2Zn6FEWt7k5KG6vBegXxLXaWbjzjqBgUGezMIqZ9qipUn6on8TGeF
49Rvt8sYWhYG8kDgVISumUu/DnWt/MjjZVbC9i8Nf4Lbuv5OgDCCVMhmCg4Il85xFffgcCfvUQvG
wo04Ui1O5lOPZ0paOMpc3br40YeuJXTrTmN9pR1lkq+NydaPcE+idAqY76qytu6eKhpxTWTFtrqO
SsdmxbrXAHzvekJGG09voG2pyM/mc6g/p6/zjQE1PHv6j0OSb4/4qt/lKGHK8BdKUOFX2eO2L8DW
8kTn44pfQg0+IvbppA//LOI5dy4VWpbCuu0tQdV6OjNxkIv7jf5pAEoXDwor5bQlMND0aVgnn1a7
UbIVbf/Sb+oYh/sxCf1Ztgmv3Hh6YZ+PILhJ69NMiw5oKu0KeVX8ifMfLQpgdc5vjh2vV830ntWh
Lt7k+Ftm2/DPqfYIX5kkE0Hc00/EXCSzuqEjWGwq8n9ypwcUMcusz0qpNIhLJXGfDqTbvHuD8FRd
bS9q7xVaQ9ILtBkLimbzdIM9qwC8fcnvK1mrGpgAhDfB+ia3IdVebp0ztCx7HX+4e5ypokuY0pLk
Bo991nKbiSStNb0gBkVNTU6LGzTrqJG1339l2xbzu9TzVXXrTMrM9C4UIbvAIdllKuJvo7mMy7ES
S4IAYzEStXiSrkR0EOlapyE6Op0+GtnvsDS266BIvSxyuaQJSoNPpdSUpdeClZKxGWVouSOxuO5o
GpSpx7tkiwP1dKcpZ7MI865GtcHScdsE5H+SwIWNd4toz+43a/T5T8IVjrqDTxUzpQWkYImzuVTE
inuj/rLRbSEiL/uDwpxbQUKNdOn5aIG6bxOcBL0r+LLnWVDMP3M+IVhjXn+bGwzX4HhjlwnVkT75
mxfa19+vyzHeQKccXoR0XiZ9QQ/mhEA3bnd2hsqucTyJIulCvL9K3mUaxTvl+uCP1RGD3udiMZ/o
BtO4cittHabbfBr4xga0gUlEzTsocHvPSQg6YaoimDHkuhaRC0DgLAMMzoIG/HcKb67HmlfmSzoP
q5kmVb4A8tZAX8jqaHLzszYq3prY+TKO5OA524S3ToE/HHZ/rtkyjq/SLPzIg8HlBWrmGFSr/N8x
IQPHEYajVUKlfWanZkubs/0WOiFRUguH1V/UmgCAZQv1qNdhCEkv6EM8rHwyX47m8EspVpYOwnqv
jUqBnISgBdrJvA6fX/TGiySTV8YmtOeAZ137perv+ACthPR+UqRump+EGOBzxtey7igG8wxzArE+
A2qH/h+9NLxe0w5ivmyuM1ToGyIhiEhAdCUrF5SdPks2/NEGJT6UYVz/VwQvs7edoNUUBM2jyiD0
gVlx8r9E/APiey0hQ+B+ixKocs3NVvqHFe1zOke/hR0OVwabhRVFeM275djjlAU3cqL/7tJxL9xS
KESEVXWpAme2ZCHahlzPAVgStAhC2u9yDVfAxAzaT88/dsRAc9bZkvqNSh7J16Xq6uLkWWFlMQ1S
F3pnH+yn1/rPrflMiM4HnH+jxP1idqQgAxjrZwtaU8cxTABsiJiJQY/4tRjHV8+ANfRS18gJUpzs
yhjxBOOdXYfItoryi1411kgFirg1DACfxRXrxLGcrfqMAyjXAczXDWBzsME+PVQFFnaag7karrN1
uctwFInRjCGOxI+wXiBG1nu0YPqKu1P29P6VJoWmMMplNxvbkechJdK17/c4CukvlpiMwdrVftG8
E898dlasDMXBPAnB8h69EKAS8zXDSlwDzkw76ZwWj+x8+06T16sZohPAnkGMpsmFiXi4Vi8HGGbd
yerkyHaMvzhR7N9JEPspdmoWWeBkuRnlM1j3Q+LrB5slq2zFTXmz6hcNZQw0k1PXdtvORGOLh87U
0HD3cKdIt9DYPZUEyo17W1KmNOrk6diu3+9l4UgrFoEamT3/6Y2vCVhYexe9v5bwHP7nwT1M3CRW
xvlHOIbgNl3EMhOLZzzeow5qvdvmhReJVcxd2AGbKYrtKL4uL1VFxHBRazi8YKu13N6bNY7c8lIW
RljfZIV8XbR1b42l9X6dKJ3PcUHpz9YLbivvFj8G215qxgVOXUBQv0ej3xp9VCFo5NPtPnTUPrKR
2ljJ4h8bpP1pOBkKL8YB9Pp7v8ArUFoJ/B/nrITqphfda8fV+ftNZtxD1kTriFHWL/uli1qyiP4U
N1rsJv/tfHHbSeYv3lxFEdEoXSmFZNL/rXbzG2HSHUqUSqYuihl9JUt7hWWYbo7QCK4820W0Vz6F
BXGHb9pO9IZL9hP1vEbSAuISkYyv5h11DCgSxd4PMw2ETu6NgsGFJKAg2fsmPWLzuNS+WLNzmID3
vf/JjmTg1SFBChwF51NmB9cN2wAHZPFl0lCXvPppDNov4pcyM6w6JCCWuAyh0ZmrM9g8TlBwV2Fl
wh290STVsBnq3mtzGs0MKT6y6AwkGXKBuUqeWoNPqnPECPNBdExUnxaGOXkCttJekbCaCfc82cHd
TEnTEW5C20be5q3D/LOqSBX3vcaMDTDhM5oK/g2OMuvQYKIpOJmxPQCBq1rJ7fvEqbgq4R1CnrGD
hTqgrUaYQydk3uid4cDjx2PYYh7BiJxZDBXEn8FKoL0ZUwybdjUhnt/gIYhzE9bPWAunPHWMlQk+
hGOmPJi0gzWLkkRpn4JKBYXeuJYv2wnPRrcnFQX+j6XmbNyY7ykUS3upkSPf9196S8/xKWgxg2a/
7fFhGnkgp+xTVwjj2KKQSAjyqglbrrQOVCh0OF2bbeyHec/3IJkjtIlIXl4a9n6MqNoM3ZKfJx00
cbS6ujRj/EmkXIhieRnWFihM4A3PZ3ncFg37Vf2rkJW4PZSOkYkV3JZURGMz9B21wniXWxEKg1jC
f9+E2yDxjtqa4z62i0X/9u0GbHMLvQeXqLzZRuF6UvnUYDCa60I0x/syGLYW3xHBIZPTRokjrErB
ERibD58OoDU2WjwPSaANwN4UHTO2LT6mGghzp9XoqzleikAykN+Tz+9/RIyE6AIwcPnI9PCJjf5P
Adpp+pk/Ft0BEeDbWCdySLP+gVg0f2IfowFlOTi8FrAaFh9ElOApjp8yImX05DUKz/jNVqW4pdMl
upGypYzMIXkAeQytQUo6tVOwAmMj00shM+5H7pqgOzgEqdBo+zXBsBeT6LiTSyZFqB1B/9ut+6tJ
6BeGA6EvxfVpA2klYvTaNYKbB0fHFcbg9D2v+HZZ+zWH5yMSyqMN1BG68ExG6KQ8yWv+XmIuja0P
SzAcqv+ho4rq3MUlgeNI7ZufX5uaXII9Pu8ZF+962Jb1A+jJ4nZE/MQuUJi6O/lu8P8ieWMyMmtT
t2cp+ktAw2widMRBYKgtncGNe/QD8hAOUrFVVHXTEjnnLXQ8029utVn4ujNJiKJyZ+lrlhVGkGRV
xusnlc32rpwAW8wf3n4Lt8Us8AXOICOrffOMTBQRHhgPjaYWDblp6vzpg+1UT6zu1kvDvQKIJTO9
lPIw7EPnAfESDXlTS4XAPmSmhtceJEwsh4vb9VomrEIu8//95Wev5zym1EtPgIrzoz3PhRZowLO8
C7JYpKSe/MBQMnDSq8Kfuh4qWrdIaKgsuyiRpdNdYAPVj+fB3F2y+Wuv7hjxxjpbBxdNfIlIDfpb
92bM9Hm+dj7PjwQiiiXKZe5FVC7U3mK1w2UYrUucg/zbrcWyVQSZYLeFvDYsPD7syio2uA8Rdv2R
E/2VgKBGuBGejkstIXE0e8+TxEFjAkdM1ZdB/tO8ZFpmbNkUUvgPoCG2OOi6wlcgy33xeiQVW9mL
u4oK8EP3J4wpKUxQFnpL4XFaL2cZIiGApmSGVJZeMXeNhg7Yi6/f8u/BzNQbpA8OKXI18NqsxHwN
Ibbt6l0SarvSeBZ/o7EhwVKWsNLaaWcl8yQn9y8V3gTn6uuTbQ35fPH0etM1zbVocwXs1xavx0Ds
I1Yd8BPECxcRjT8NR2kheL9NwLPQcqvaYoa5TZUqNgb2Hv+692D9dxoKFi3Zdn8JDS+SpajEOBb3
K0AXiM6tnHfQkusnC2PgXxwMg6l424TaMihXAbhRrfr21Dm/JS28Rwa3zJuFuP8GNXx0viMplHZq
9F+/e+6u5dncX8XenL/08PhDlsha3JBH1Lvwy716TFrIr82RwR9Y5Q27SdH2OHvH16jW2tRx93OE
TQ03X+LjHJAQhtLlN5b/Fh/ZpiR8BixCDDbauBsBrMtzmWVG6k24xOc/0tzgy0i+hlzaOVKJzYBu
pQtCL7TT4cwO/svedXgOqu0XEkSjl/TM4ueBtabmD/S6CU08s5B7ROl3zjOj8guNozyoy7mrRNv9
uN2IH1+e5kJIRBd9KcRzrNwesHSOK5rg2cqMZ5p3ab1tfS2qyvD7+rMDcZBtNxEXl9Ez+rfRFgDl
d/+lpodCksu5seb9Mqa11nBKfA3FVqNCKuTO9JLZ3EM88nF3XXd266GAtR1w2xlhDESphwwLDVdv
OpqFapANWIpFa2IuJdwv5J5zDYW9kN2ZvpkIU9q60oDCM5bWJzL17gp7dfWCy7UrkQAHcOkCjlCR
v9upxnju6l+FeQppKPH+unNHqW/EC4LADLeej8nYUCoWOSc2H8bNkpnOf6cfxGC6BdMuo3dl+aeX
kfW1hObvrpYfklMKvdNlwXG/T3FDruvJF6lEnFQ2oSZPCodGgTcZm/YHd+mXAMTZd/154XrZk6J4
n0rR70pbqEbw3I/4rX35tsUWrHCOFAp7gLjwZ4nmoH6xtSIn/WRvyYuRocQWGIPJOg3KCBBloh1N
ZjpM66TDVC6v11VkY1fbptPoPOR2qE8u1dXMK4imCQnGJmT/qI3RRrKToU8tGqb6JMktQkwHJ4im
JZoTe7pBFIV1xDgJJNj8Bn/Nz8oIjBaFAZ02l+QJKahDw+u6k8veOezcHyaDb9Vrh7CJaphcDW1O
ErMXkxK0d0/IVqrMXu+ZeT8yUW105NHBxW6W4KOwDMYZ8VUPZd/vgn1H1Hy8eOlt6a6W2KaDvG4r
hObe82V4BIrrE29xHubEi0iEM4q7b4Pk5izgLwydjB3RE4bPK4df3mQ+jCh3gB+OKi9sT8tJkv9T
9iwBmMNXPEdHdNuXFQKT4mdZkBFyOkO4pQ1iSaWTyaaetbfsEpXQEunnjobLjyDvZP9hpqcvLg9w
GobrkJzLkE1Z/ICq8bcpFiptJdma8W+rlVcV8WvEkxyFGlNKnJ13oLYBlEStuy7QHR7WgxDH8Zvq
cdGcQ5tTdg+diEF30IP6NrS74DNnYsHwrLPFI9J2lXliffOL/acHF8BaLLcsDhMI/KYVZ05bNp95
HwvRr3Feno5MWwR3q15YCybMUux8vp0MhMIQpUFoWo1jCIZrf4FGzzdRhSzaMkHwmzZsZDSxMCme
ILiSSGKOvUJkFRUbv1KCgy5FvQtxIosu/euQK0Qx7boWlKWEhaaAeNimMMCSWoinSyLx6axoJyry
d9+kkFSGqwiiALLd7Rcepx+ySonU6P3jXgBbgViT45FYoFqtq91cUXxR24l7nszfdHe4Ne3BTopQ
DR/nz8T2W2zcw4lS9XtYKwB8jm7L7qRvX/HHApB5qe+4ldXzYT0DTAmPO3RD8Lug9NwOx2HYI2xF
XobcllTmLAiWfGVydED3J6So5J+X+veFnw0uwrTZ66KxU6L8EbuoLtUVNlMaWBvwzgEi0jmbXaa8
BDuOZ00+d0XtUpb5/VZds3qlQuEsgAo59I7amhh7A2KOkTguBNGnNv2HVfSHfaar8sqSIGcOU032
ooMRlRfz78Z/p6hTG88vMWE7nO8a9Fde7sKtqNMinWqoak3b+JY8tZlKFtOieHL5XRXjryBr0moJ
gVDQKPDgOtQMoBZKoHGBGMYLGJ49C8UeDPjk+Z5HRXUV3P5ruLJCwAZSkG11m8V47qddnBUsbyYh
R1qf5RC1k8rsClXxq0e/d+aN1QPN3tDx1dCrdBLTjijRJ4YGY151GnACUdPrKcZMn4MwUi4klUdE
Bs6XVHB58H+NPVgFBOQGsYLxIEKgsuYcdDC6US+mtTYk8V2Bddw3bIeCxmoqFUxM2JECdr0j/XKw
0R63gpZC6atTiQaho2GBLKHDeL61Ox7x2VjiYA7FSfn6UH+wUw69s4MWTbGxc+C0Axs53o66OcWx
YBvsdbY5dbYUhUttw4h0eqsvc9XLzEUKUOWaSPXbDsWnV/XX35msVVlePJpcubgagpmK7PRfe0jS
+ANmc1a3Ij6JvywZavKDD8Ivnf2PBz8Tc5WlohU/3YSkLy9vg6rih0ki8gFFZtmWNUgqajWFxcWb
xQWXDrMGw1X2yVrgzJFMyqhFNvJu7AUyxulo2h9p5Z0cpXbKCQuOzZFPKq538RBx3eaadcm5ISPs
7u4A4sBMIUbKnzOGdh/sq9IB9Hkr6mmCV7QxTcZGzUXV3Drlqm5LArsXk/OK0ry7Jd82T5HfiAg4
ctItnv20MZhfJIGTvjkpAheuiNVtnomVKfNAnVJYmKCvGHdBrcN0YO/O9aLtMy+c7guYskuyrP6o
STBAteCRjWWp9EZlL/k8SjZHS7Ar8yv1zY/7TmsmfkmTAWe+VA+sGkYpwZPklqZSb5KTm571IwSv
njeFfOYxB49xUJgj8idugJCd9shulADrlCHS4xjGNHC9xPw5nFgO0LC50q9+L4v3v2mEQDAU79VA
vkzmGFJsfXywSjmz8fvt1wzm1ozix1dzJKXIf2ESBIRD5FAC40JKPpX0xTvcGx6iRrZaHBMd7mbz
fT+56ZzTlUw8GFbgn4rvTq7RbVhcOmb2RNEh/O/VuOBAbdq3PTjDuJ1CJ0XZPcT6r8A4YJhcPFkY
AwPkWDXMwIpIIvGm3NNq4eXm/pPkB7qwp79lNMY3WORmLnNrhmUlcp0VaRNbnV+y+miILbwiOYXz
Qzxhr5IqE83WrKpg79pTocS5MqRepS6gNDXdPqmtKx8DbbgwO4GCG+IDmVEIP2Exw1ENLgvaPcvX
FmVFi58fGhem4RDi4Y/XOj/8KTXCa+32NxPX2EHW1+oBx/sXvGUJFR+4sbyYG24hebMx8iFkjAz2
DOJUoVGh07yDuR5nz8kMJK9stz5jjCuDZ4HeZ4kMK62oX+HoR5JmI+JEfvT3axhRKr7Ojx3GiZpI
ZppkoNCNE4ClDH/4xbBBNxvwRJjx1fLJ9W8EmNSOr5PMzpsuckXpGab/hiAd6GvCz9RH3X/RAMkA
oScQ+apjPGIckBMJi9dY4YSh1XxguTIx0zFPfbcc/qj+eal2s16ceCA3p1GQl/fPGNgzxGFrwCdC
hX7b5PCZSDlXFHt8b7kDM/9qLX+vKA3U3/TYhJwqmWw7SucnkIq5zvcWb2Ys2oD/m5mcFRR1cwEl
hZtnj9ZaZTIt06A9qRSrooeoiWHW0k4cMLEuJjQoioXm3HXNJL2VCRLrgR/J6RLsiTDLpbtT8dOS
U+/7/Z1Ee/x3tBpsR+7iVJKJ8YXD5dGyX6gwWZBBJ9JnZDneCMZpl3p+kENnEEPyWRb8wDceWQfM
zL0a19qYs6IfL9kg3OnGEfbPW+59MyUTNUEKymBw8lCgp9UwFBLEXBDEAauTsdJnUkqv9ORpDxv7
34iTSUCsnqKMlXzLCICioYi5QQePnKc4KMvS0sUkGnHo/2M0ad29kNXI/dyvBQRplqriBU0vAub3
X0K0bFsTKusRN3Dh0DPCsktVJbfQKkfs8MBFT65Owv1wG75ZlEYN27vctHNwSe4OYcgRuPcLOY1U
QuQIYqw0l6a88YgMtvqNO0SZ40KGGYAUpg75kI70mCJtSD6nVqkSYxCm9S+dqrrVkz2F9wFtTWPi
8ec6jjXHdUolyVjS6+w+cj+23uU8j9rNvEazS+vSAPkrV5dz2KO3MJsj/6rG6rzdGdbfUmgWcx8o
oHBN9Ie0DdWHSNw/iKZjiFuiZ21Ty5kZChIFxK9rHBJ3Kf+cA3ITOmWtZgKAd0ixgcAfvD24p943
SsghT6WiojUxtttLclJFnORIT5BP7BjrXBF8Y2X2sNP7A6x1rd8OWGlDVTEXe1gYE5lTPJEJUClg
n8eS8hVKwFBHtZ+lw+Tv/WDUVB3AusFYSacOmHuj6xDvykS4MsZXfJJAdt8xi1AwGYylE3IHH6ZR
nrYirKGRRa/FdGYi81euXk4HJGRrsY89ae+pZnPy0YIQBIOwJDAWoyl2P+paAkcrPcIfUSa20XNn
T21r2WRXlS4e85SCaRrgHzMVFMuJBduXSt/MHHGS/9jR+S2u7WHvApuj2wpK64lPSaafs80cWHd1
iTRbnYc4KwCLrRDxn3gTgSFZF5c9VfvmBOvfTgBOmNGlXJwgZvLhuC4vKrawmLg2f4Jl31KtGNJI
6jBzS/OW6cnXBwvm759A2THP5fXDtfth2M87v4BOIYysAHLgVR67tlIjMOMOB0AU4FaDkIA8gbaK
cshXCNNJyE/t7uEMT1dKdiygR0Po+Ot1uf0/E2B57oQnG8d/i1S0ac7HbMyJYbJFncaWU5pzHkNl
9uHBdhRS1bl/pyHRukQoA0EviTi18CWaWhUi4jabQxyb5XxcnGmgn44jGCB2+e7+dYR4SGtgQmSw
5CtP6fqPxV5etHhgYhzBl4KsCn9uXDMyFY+3IzY76fp2h3QLLUJbGj/EBuht8h9CX/AuVeBQ73D8
xCzuUj5oXmL/1ohfmikCurMNiFqjbczcQ9/aLO1jycTdnaLIN3Eu1MEDEjRoaauN0TZELw4O1zBB
FHJOxAXirG/noDMPxqH67xBhc7DQRDgb2sOUQBrbHyTABWpRyq3HaGLeW6L5pa14RlLeJzdhOJ5x
Gc8913oXt7TcIHVdx7MPvpkceX6Z8AsuoB5rMp0KuME4OTfCHN6sR0HPkRBI4/yrkK7zxp8QIZvX
752Sh+4mk+Fg7bfL9v2nVIw5vkD5fNvYrT6JSVWI7ZA4az8eF/7TMY8OIM4SxygFPpiuQwfF0aFC
lD/owpi1RK/NT2NtNnAix+HL6bEudpVIHu5y0mnqnVar7d/w+NvFv1GGoeO48DetAYCgot+MJjju
on0X61mbOFSp1uSe1kaME+SQ3gdCvA+I/xD8UEBd+6t9ObILxRtp/+AzIS5XtbNtORScHF4A9YIn
ZL5tWxUuh1xnAnYbjF3VsJw+ZkUpTmDOAXh2Ol+MV6QCmJGDLLAFTZOTIl6Yaxr5SLE1kvVNnBCh
WeC8BD9ks3d0QcDfJN26M1Uf9MpXJ62Z4/sy6qWIdBZSL+fn5Lr0/OaRuPjcW7Rkr7QaAw3EWdh2
JkLusaSpgNTNkGwiY4QTpxqDh1Luimh9B1EkGmvUfOwyjj8F5brCHBeUOcDPaM6avpcdvq/Gq/nK
VfyPlWWmF15LN47DNlhBu66YRFSWTVCs2ExOajFRLW6av5PUwBMVo4hFkZ4hT2u5wR0GjRl1HZgJ
k6/ccb9nYFVFaNUrmHbVtdnnGe25be96BwFUs/ypo+z1Iu6pHghG2Samh29GHOOlPsT7Lw2pzMZS
om5MQUkyOUGuISUNe17ZPRfdjKjip0HMMvicSmrCGAWvZZGo5I8hONaM5zhvOQGdgJKRpZqAV3+G
E6bqCnH1psYEo5CKx1MTfJSMTba0Ibigb1sEO8jsOlX6xQioeb4bz2RVXFTxmXULALCxJJJjFEzW
Qze1hBVbeafSs1zXRgSe9oDVReADpf72ZknzpM6cjBCTgv9Jb9PwLN7JbrbWHcO8XrHKHxfMKQvQ
v+z43S1PrVXuc2P64EVn6F0c8hsaAI1rXFo3gbFhRBqtOKmkloA7H9XD0sAQmj1UIiXrOA3ZpJ2R
tb5RrHoTKTV7EBnyWZJzB6BJHYjwT1LRArmG5stkHA5vecOt4RjyzcXWpe07pds33ryIFNAO8n3B
QGexfIAY6l63h8G9JXvRKJ1ZV9D77e1UAi9IZ3/Udnkqmxi4Q3Qoho62wBMMu0xWAglMbWHYUtbA
ongN89Q8wTxmaoe3osYoAoVaNkQJ/wTa+aGz6MSQEpy9WZ1/oKZE5wtx2TrntBspKns4/evcZnCj
KwZJzDnP6JDYMvw77r6ehaudFlQF2uqKsjXxm+wM8hHRghSAPx1/TMcUHXrpzt1TyHXFtYn8yo22
CwV2e8BR0ZWKjTHwCat32LEWQRNco6nsSgCpAlfxyt3Evuf9L/ZqRw40rraW0ZRteuA6XTUU3lIC
1045B0FZ+0UjGryDujWhtqOEfr5B++GmRIoKJTXASp1t46cOUDXe5ZeiPxJvBquemn5XBMEr4FL6
b7+1acE1VcxS63NLu5rLWtFtPMoC5MK9FT86fsdCCTtCKGirox4jPXdfy1BlPpsFEKgA4xE3uxXw
U1gaO42tDBbPGavEqDRk6QHPEnu5kJTc8w99CEfcZ1KYDg+n+e6g1EBqdVh4MjgRPxF5EMZcF9tF
QNlhoxYnif5n4OyUhi69k7gGL/ozlJXjmAJaSMayzLMoEOBdcnU62Rg6YVfNORlmW9J9r/d9iEzZ
JDiYOKhP0KIxjIe+UkidPJIJBN/trvTxdFNesdXajZvDKCDklVW87lHkuhw5jPE8BOQwRQRR2QZT
uUPxx7bc2saQGuOVtUCN8IKR3vf2nltJh/Hw+MjTarEQHtPCy1Y5WJhx9dZf/1iVS+NfWpjbP6k9
5XouEwLEkDa0bnCPkbGTnlnvxL6KFOqP2EefAvZxJF1Epl2UVyDqW9H82Hlv8a8F7bYVkjhkLzFY
YkzfBhyBUWqfh9Dut3gFfDOxuDg9kzrlnbh0rZWuQoNaLcvbXNDA0T6ACOPX/XT06RscfowNoyDe
uNnhb3/nrH/jGOol65xt4kBCeif2VYoEcZIYZMnQ6dAwTd6cw5WOarQXeM5Ivbq8Y9Gk8DYZ4FxD
1LOKFQeJ66HXD/6BqGFZm2Hd/fHaRzWj2D0UvqhS/yS6N+osKS+0RprAhiPwhNM7D9zC0Ys0Wy0m
JE8VAF1bgBCKp/J+pW1zYaDFC8AU8EVkVyCQfC5SaDADHOuZbrwqasczzYtG3eHiVnvV/gG+ryXM
KsHR1ZkJOMrpvxEfwXoWtuByIh3l4THkEGQrdRFwdrsceOlBK1lZB5DvUo0xhSIcFBf4Xw4ZBJFV
yamIVN9MdsB9S386lNRG+0wHHuzz+1bWw+c3ELG+NIyKb/OAgtaDJDf0e5dRT6rHW4TVWOIQgjqj
AfZ4iH0jzw6awL5dzPtbB1es3l+9cG8J5i+OCQU4dkmEmbvPnSR1cTwNUF/nhv9LQQMOq3S4aHoN
0+U4/UiInyr1gzg8+n1FM+HnxmpjzVSJYO8OYs+deKOJQniJEvS4jMujwzPt5tdqM+P0esmqMWMt
ufmz7x8GMSrc1GWDBo/mYJzpvihqhPnNm7UrPxv2RfD3YdKtvj56v8bCtpJ0x6RjMmQ5Q+55+ODn
hThPQjzu+U3l0hHI+/RtPgfk6mbujLD0TfIgcSIqTY/KLEn9tQXriioxNLImqNtpPF9IZQpilXo/
U4fE5vbVzDEXhY5NLXQYNx6zGHrFNFIiFX0+Dd00ZSdUUwNJIVHiZsoQdr8zR08RSy63AanATASu
RcjdftRrxPHKspEFS0StYEFPNqPBGSu5J6LcFnmcGsIhzFuAGgbGXtcYdyEASooILj/SQvs/ZvV/
AKUCBt9tJGXem9tyZDGEHTgAygxaJHhyVKk6MgTpV172PTfEer9hg01uZRBjtqKvdBWNgKa1Y6mW
w7uea4qBPRjdLP6t9BYYK7qSc+5a/pBgTjuA/D5m6HrcIAUz/rK5vMLAonSOnIKcDTO6f3OFT/0J
+W9tWzCbxpEbcr5Fjx9iTdr4tiOhCTVAw4ZGibtk3RaOCFLgt5XNgMrBjJMWHlcNvnTk2+k3yNdd
N1l6l27e9POU9MtaXex3xI32hvYEyZR7JkMVhIPDL0U9t2LOD1g/JNpCbZFnrwxk530V8ZTHhcix
YLlNBTe/kL/VsEtWwVnXms4qme/Pw7SPrBbnSmPBbWOiYpdMhmVcMAF2GaDZamwDs2lMUtAAx73M
tt6RjRnyy9MmdHJpbmh10eEz826/6qi4aWvgZ0yTKsQLD5V9dz2Jq9urlelC8zhPRm2j7HUKPdRH
uYWD+ZMi5ZUcxvDXT0tuE80fcd+pxxJPcQ2K9wLnbd198t90Zp+cOVNZwE5nISEb/VR8UGCkIPnI
/dIQljTtEuqkHFdTL/WwIRXkINSVLcLx/pqSKitFHLUI8yUWTLvhvi7eVbN7bf8crsznIODkRqua
LsbfAZcN7olfaoH8wRE1RtP/c+c+oxBiq8a9BO3fYG1jDmLAD2/NqqcEYIkB3zJ7zt8wJXrGqHfN
DjNqBJnE0MLrE3ox7d5oLwrz257Z30Llf1ve3Rczt/slvVSywfN3Oyz4bN3zsYphqxu5pTYJtRrn
SucDDHh7+k28h6oPoiJTyZ9V6VDgqUITPBA6kGbBkwnpQB0BR9AilADKL2pwOsskWUXGSBCfrVP+
RjD4tjhivrsD3txqPABfnlGNy2AfC7XqpR2O3S81vtBYMGNmBK1QgmscwRcUupM7wpP196LOqPuP
f81YVqVvklnIHx0IkVbW6PRe0Q8X6kKlw72W2ReWlZnZU/YsEvTCZhR9kJobOzXc1PiUiQSMcTc/
PXvq+eF0E1xDuI5K8fS9Vbfn28boKfT+86S3V++IPX45ai93DGvu7Psu7Xi9tD7nenZqXQNhuadH
y7tXHOyOBftwfcVfFSMJgKGJ+ggD8Ud+BueCTi4FMqFqrvtB5iAzyeFu8ihEPiYS5Lpdu+j2QHCk
NpMzFkCuoihXLEn3xRYoqd3Fgjg/c4QP7J6KC7PCt5s6FVTjH5cBh+JNEd/sMdvleBxFiidI7pT0
Mcbz1FmqYah/51m8h1aXlnRCp1jHfDZ/sgQ3ZakEWd+Q9vS5EXgPC6uU46XDBSoLz3FvAqgCplXh
5I7MYoHF+Om5fsVM9tKRnWdoP+T1CfWBr8zV0P9wvMbZ7TspCtlR0DACEZmDf/ieUE958kpmy00N
O7yPO+yhcPPwNq8HxiDNQXM7soUybu0bzWv/vVqTI5djzmViQcNDeEjz6O7Yhmq5LyRHaDuYsRl1
6GeSZtbo4p4TM+WOC6Usiq2zfhCsWOFcbRvaWGPbosXBIsaaic+9Hsav+tjeLajMcbWUxjJhDZHv
1eQYvKVoGcwbQgI0ZmI93pT33M9cVxw8RP0xl0LxaJSn7RIkY1uike1dcq1brGlF5LgbYFXORcAP
Dx7Waep1lgl50Lk1fRu5n2e4HhclYZ5mycSgN06SmoMxSOwcDHo7BFRqo2IIyau0ewJf0YJMjOz0
2QEh6fy3G3gvC7fwnhCkDk616J6p6FbT7UNCH7z7KydgzgS2HIPZ38ZMRWr8q9o52Z3/eT0Bc61v
PWySV/smTLcH/GJ3dhVhSdB1rXsQ517y7Tlhbs38CHoSywpU8aXUhyVCXGqjZFLICOKDP2zThh9A
Gdh4POm2Zmqg6jTXqUsjUBDdDWGdATx0esbMHzoDM0NJLrWv8FzQj8MiwoIbCjAwPKiasuLWUqWj
5gmFD49AXMrbS84/Ba3gVnizYfAXrr91hzji+Krwt4VC1+tUFh8WqBSCffuHqW0UdEXLgkcp/WJV
NVW/9Rz+hMEEPKCkfYussHhKg4G7MVXLbo/biN3zLAVaIB+5xM8FbDXEw/RMF/fJpC1aYTzZGoJX
7oW93JPwBzEUEyPfOM5f6CzS1uu1TbURkW/qRbYuQT7Tg6gSmi9vhBwphoABepCAB5f4zDlcwTmy
UwrNOSJwBAhM1Vm13Fy6PDsFBtkw8HFMAM7onTIqfWGuAVONTbvDVVGhF/ELe/pBIMooLht8qoCL
8N9OOWor3iu4bmFmKiRrskNmaZZqvtYSV3ON9bjtG+NMrHd4+yRkEzzqfY+c6YdWaKHIpkhhD/Ao
f8+nojiN/VqQitfgwPRHr/n6Be2Bj0DDNfdKehGON1SaD3d2FRnJ7Wu5rN+OUvnAO8ccR+4mv2p8
L4ljyXxM74kTNIrEZ3PxH4PIkCV1oO+WqRqsMkpC94OMC6bgOZ7pgtd1uWJd4FIhyjogbUy0xKBn
AesTD0wkLgbj5IfEn6+6E5OapS28Pn6ENaMQRaVaGXL2iy4abWLFfiSwLX4+MIpOKfT0ZrmZ4pCY
0egnT81rW10Gp5a3UH8VyARQS98f9wuWtL+QACn70pA2TONb99fp/AvQT2cDqXZx6UP1W15soocf
nn6Bx+wsGx8CjetTkfKrPgExcrIN25CPCN4KzGmq4f9MvCG5Y2D0TFz5sUmWJ6KcfPMYRT+qYyUS
5MQ5WOrwcicC5M0gRFklL1JGbgJQ2HKuEMPoWlaDQw8AJRvITY1MFhWZUYu2uV6NKIJbZVHNLO34
SeaotW1zUY69v16StmjNuiyZa8NHxnwhrJs1q6KH8kN/26ILXA1JoJpd4Ow7QzzcNc8FLrlFULv3
X6r6nB5PVFfhs6mtm1YejEmFiCXoDeyOhg0MsWlDacy/xLmAcFtg9qXeTClmP8XHggnZhgotMFG4
+vyzs2NSzMkccY35skEXdMOpwJrRGUnwOBjk83/gTZpwFJILd4vkzABck/tZowS05wS2BPdEAEOW
nLvOBV0NiFyBjf5EF79JdU+GTsgBX3jZPXm5i1J1DVbmynh8fR3ZNQh+a+kZC58snKl4VcPuqetj
h8yPZ25dTMxwoLS0ANK1EC0K9nxNc4PWwn9fDgvZTCjm76screu5go7mj7CaHfpCRhT7+h46bPfS
w9pgUmb4IyDsr07UhVVZqzamqCVgOHwS/u1K4BXfG+YVkgfy1Wco92zeKl2TU9LLHVpY/ziKKWNT
fLxHrzNPQ04awcZzedxCe0Gyh7cDIH3xHvmGzYa0ql8MZHWTlBjwm875sgGbDqyJVOETU3XNxWRp
HmpJewJ05bPbrmMzE0MdKu/q1b1S2uGNmZXZcWJE/C1RSNPU39n+qcQhvvgRLqNyjZJPVQzn/bw4
rjTjSREQlZ4TG+4FL+RuNTxz3vHsnMh5e6FaPWRpl5GDnU6MxlbaVb2b70HSeDnOYYEycOJncSs9
KYo9beWXfZfXmTL7BXdD3tDFOBoT4eK8wW+w2g1dnVszp825rC+TWMmaygRxjo373a6XDPgQjb0S
KegvxoiUrbhxyIeumrWH3Pu8SOT5KDAOYZ4rLDDyJ9PjHgYdvuIKHQnjQZYMBTNb97WAZrar8RQY
xjKE+ShMuD16d4LkYm4n9cWz8TCDveWmicp2n2ZvXNScfq3jiqg4Y739igPiOsnFb96t2P95GBRM
DdezIik6fBa9ZIGjJoKWhj6nYrFtJG/Z9ilxpWs4AQaPzavHWtn7aMpPrStT3ZfniMea0koEPQvR
1gGzZNPIRleUxaLLypBwbBn+Ay1yqFhgm/4vsExnedjPPhKWVLYCke4OoYJ2woPTzQpihjEAZTZ/
HY+F6CnHDuNSRfcmhYhgJfsot1rWb4Z/bxEIOyCQnz0BLCM3arhex7AGg/t0GbPt427C2Bad0M5W
yTOyIxkSphR9IsW4htbdmQe9YA79ts5Fy+yAyKyKbz/RGeoZOL/1Dq6prLn9Cl3Q9NFuXVxRcnbv
VSMZcfHs0yfJWsShYUR4P/2dyZe+vlj9egEvl17otmRzCNsDV6Ep/ItwKk1vP05hWnB6BGB/czRq
DZPktBluXXywvzjZam0vKyattiTESnfW2UV7cy954jJRdo1jUhESX844oE0MQje2Lp/dRd4Vru4b
o0XiQlKdmc6Ivbsk7BqxF+OhoDIFDXa2MG5yQSsN25ldL5HjnqvjfQuyxaTXkY6OM2gDligftHW/
inUuSk5Zt93rMqvGS9WwdUQPecN5Rwbg8AuFW3MymE4rNp8OctQpcBqzXHtr6MGZp81hQnitZoCn
3i7JyV3mhQtjFN+TG+qaOc2FluwssIqY2wbh/tpHRJdDuXDLWeD0dW/ZiFO6IOBouci8x1Ln9rof
04fGxeDX4bJbRi5F3Y+w649qty9SxpSQrHyxoP42syvQjxa6tlAaEhh4Qguj7cutVahqHdEjZ8d/
4XqvDub6G40GvPatlpI/XBApwze6Q8yKYPk7P3O6lMCHPXipamhBWnthwwgeqcLbSIwkHnMBorI6
IdDeDIxDaNXNyu9MJFwR9FWWNVCTNkiBKGiSCjHPWPL80l2kZRyU0WGfSlQsjGAOV5zqZAla4hCh
KfSNGvYjNvdSfs2qcEMnEoX6W7WpLsygLm6pJjSUQQy/raVqXz65XeG7c2eil26xGPKOX9KOir/L
BjloqDRcBHhpF++MvJZUVhBPTa0jwU6BHLAIVrIDGmumxCub4xTh0Q6gwe0aZSkhpwia9yTR3rTg
NQpQRa4R1DFr/KhojzPp9EpRHXkaTlaGKr7/2FSjr85MkXu79ArsinM80MBy39HXdhX6NNnbcSws
oPpcdZomr4K7HkhF8+OhPG5S+obQqLVuFFq2+4Gu2Ce07DTKAYzN5UXg06m4E2UyxVsKMnZsm3Ae
cErcVLxVbOl7ZfXjkmYdOCRJrS03YQKMRt5JkzCMEiz8MBjRPZp7eqpn3AM2yaS+Dox2s0u4WQ2s
v+PANl1XJ8mX10C6g+d5DHwC88GbbzKfRLF6idWOCwI0tZFSdtPYQp4NLIWPzpF0SOHH7azG6OIa
YlB+d6sI3Dbjo8064nvUsVrMIFekO45ik1+X5uU7MxEar36jtqhkI2jFYPCfzQF80RpMikvYV9eN
MZFirbKF+dqhErKlsb0qRqduhADY0lOh1uUAW7ParY0bw84p8KNYi7ZserFMK+vSqqGYoFp2Xe0u
cG/9nP7hEROQqWDdcV7fRGNbTCw6pvcdjBldG9ZMDk6VPElZQn7huwvtHHV2NM5lwKG6x08HUdvv
is3XAs+s/rfvjNE8AN7QzGmv1bWnDcp8v6f9yCEDxa2aQV/C14A30LfVhdr8UuhdpKIBeCZduiul
M3hQxNnTpEIq6PG8WPt3sLmtaHMA7uAqZQg8drQJ8ykmGz2FSH44Nw5bnMdzVpZ/xT46D8ec8I47
rxhtBafWgu4p/hLLN8SQij7JtQDMy0Ns7hVS97acSMnfqUEWBZrC1l1rOzQ4kMlHQ3xZ/Jxxvq2J
O7P/isJs4Qir327jYof9Qrwb3m4f9h3Pf2H49Rtn3NnD+WuvLFF3owdAML7CsFnKwv8cTRXxj9zf
pVEavPwTfyBvarssJe9UmYQDqN6cBTj+NZog9ByGs6xsfWN9V/R8UerXwB3v+QgE+bghzmyykPFV
WTwFyQBUhR1YpwUD+zseXVWXvaNxYZII95JkVyu03yAquQgNMLQugZNzLuG25NjQQDUvBmo97tAT
JJE3imVLvUx0KYGkKyNCiF7T+7nbl21i0opy4XvTkfG8+lUF6B8/Xis5mrdkDHhB+qoOGNlYhgZb
yHCdCKyOiANtI1Pb/EbJ6eVqKRONAx4iIp6O7sHpLLof+OaGk1cauXwUSr6awqYxjaDsFqtDC7cN
lSks7gdfV/AUjyaRMcylko8dK0Ig7KSQFdwdPKazZ900u8v0h3yA9rejASzB0kmYBvGQjX0nbVG3
5oONwKlvDEPPaxDmGWpWEHQp50FczONYjMTYchXE1mE4pfAfZVyOvpbF7H5KrZz0dCwBP4Q3Hf3I
mXNNjw/fjEuX3Gu7SPuemRFCLMk9JRFw90iG/mUcSlDKNa8XQrQAFcKusk48zMxPUUQeohATje0p
QX/NQrO2BfZmAOxwwMIWTAlbC5Uo3A6QggTmttJbxL/nL73SALQGay9ovs+ANQgg1wsMX2Vf/Sus
VzKdzlq7NyN1tGLkVgC9F1KCTcnLSNSHNntVaf9qPc1dv2eYvkVLpnzN8Cgh/rUScmGz2qAZZE5H
jfYhr5+zbL+HxijPfdGQn6agEVTmQXlavd8ht9TCN1j8GJgXjKgdcwrV0dlNQ5EYOPHajIlSV8Jl
IJ+2ud1GJNtPaDt1ej0oYyzesVue0FNXJ0/ZC7PT8lBS4wHf4aQOxkN2gcFWNuw7pVg1YoF7j/7C
l11mhKhES4AKUs+u3cqjCkR1aNwmWx7ym1jT90A8g+Of640VYbQHypKjFtwfG3StYJjkw2DlB1Tl
aC6YfEK0XBkVKvRL3tk6qnmh6eTs+F+eYtUNtTVWlikJO8RVv4m8jw2zy5GhULosFgIjMMGyAr5i
gQht4ieVYgYJdFPp7wNGpLevz8ZsFXe3dFd5GqLfshcFtxpOWJT788uXL5Ri3rrUREwz91DVAk2O
EvlT9w073VOIzNYuOJgm8SYhCrxA2KSKpblWu3l/xd8S0hFwrboTHOEffHoZzEAN6ttTPtp1nr6H
OfDLwBkWaLCTpZHilJjxF4Nx7jDG4TM3vleHINPNaGZm+QRWwW0I4OWMTu88plem0mWYmYrhawzU
pn7QRt6uDb5XXyS7d68GjLbbaI5qPre4fTP/GaFsVB0tEUUhvNNjsbNhO4wLgkMirfMUOo2KHFnE
7gAUGh9c5GEDN71eWINpbfmAN2fVeLn0gkpPzDfZlgkk1vMvfagWVqVlZ3f4BBHccZkcp1nuVDdx
tOoWa88MWzHlKfGL4tuxVF3tbAoKnmee8sZ9ERNxp8GzDJfGiSb7kG46FK40Y1DG+1+UQDmypNXF
6qEEibBjZfmYsKXtaAgrilKanI7AkT/WxRpbJXR2N4I42vGLTbcscgiv9NiU29nbycDCa+BJtIz/
YfCovqnpEn4qmnUYlM91jQZsp5tvt3+oI6iMWGgH00aDkqlALwOigq56IMLVqdR2rIdKisubm5OI
iEDa+EelsgNqkIB2TQPRUeat7khi7Me8DjWQKE2/4/r2S9bbclBDBZuUd4gcc1Aw0fKZF9kc7LNe
QmwmsOFhLG6xFcCwcrTS9IxqfuUKGm1991WVxJACAOhZZxwWDG4RyJPo0zhGjD5Ydsh2/1psmr+a
eq9rXEdNPi8ZlTZz1m4WtgiEcHf3Wb7fxuM2Qv/nW9cGpdh9vSKuALQCayW3QzpInAaEVShNC6WF
Zi4NF37+YE8hld/17E14hfhMN7KXUwEsXpkwzOKzsSvYYTD+aZxWjggsPv4do6OxzACIL57Igw3y
4znsBfNivgeg0VygRIUpoETTZMZ5L5zxHf/QhFdjw0Q/FcqsCrLWZbGD84tdnmVmG78rv0DXcm95
FqkEOxpCdS5042y0nMNO1l2XBGckzKL6ZFoBLFTGzmg6BRsegq2Cpdn5m7n/HlCiwZihSXewu7h5
0ovHiQ9ZncywH5hhdt3Y/MpdBXsPvnH0UhlClyDyk+BTu2nSCoPwWZnOnmZJDiPktNEDdv8ALwt2
ZhlqkoiBw39oFJA+TqdX81+ALvVE7QpEXkBVtcw4ro44rldU4VVIKXmVspAAXG0FuWlW5qpNhzWD
p0q5Dp0dLzlIZpqpgFwelc+7U7nTuljAwi1sjUriDFACYl1ITCQ0HoqjwR7EtEoywDSfqGgMiPwk
I8K8m3GRHiw+m9IbpAfZ/xtyDt7PeXL0hl2USPqFsho3kvaxvwq21kGU2oTPivVoIt2S5t/scUDo
a5PSl9huqVsDIzjCzjam3DJff6GliHnZxcBkiq2ja8AcDKm6VpHn/ew9WyETLQZq7GLMHwbUEVqU
uhzEqDpAiM9arGZvhp19u0A4AXpOAG+kaMLNXz7L8uN3odYN2yLk6jyAdhsdsHrTpVP64aPYTTtz
CgLNsLdisRaVOk/wh23MdrYjK5XYwO02KvZmqAqL9H5SDC9ADPgE5oOdDzJDHJ3GiPwC1xRHb9+m
PPYO/aNpQpMW4Y7Y8scY5t1GC32v903zG06Y0OO9Xsg25vCCVm7nCQ2Gc3NmtIMF7szuNHtqFyV6
XHMNsv3grgz5aJYsE4P96NnAMz9Qv1eSoer2Gsy18KTTbxPVBvGPrn7v/AHWuveKK2AgD7X0/pqz
AtvrRhyiAfpl9OIcU+eyxdAEbZj6ubi5uNpN4A7pDpFaW7zFq3XmU29W/z94K7CPA9+1JHXmzF2P
DdCsnMZNq9rpVrZVX5H72z0ZECTH9Hsh8NMZ4ifwKpe4dRT2ZrGVbJPccy1EhUoIg4loCwocRVCY
YJh19i5iLNpLW5uuzfkBkwqYYRsRsfDvoSeGGPCFZMUYdXSzvktGsVhtK8wLtjy35vH1gfzfS4I/
npcRMGKrjAacVt4iXcK9jn1JGC2LXagZ40pq7T7olLqCC8EzI2TJlUhnvB7w7LKlCG65wu6umhmL
2Kt0BGcU9XyEHugrTC/P6jrt0XVd0w1JPqgIydPrWyA13ar3ey/vV1iva1fcqrvdv998l3lJyuHa
neXgraYrxyXgaToF6jRc0BR1Uu+mobufsAS4tfYpuLO88AUtuec5vl+oDEsqIgjmf90pOnJgMUvJ
hzbKDxb/71bW1/jzQMr18l4dd6ht9gR3iqHVyVrKQfldGrMh8Do0nkt8NFtodlF4685WpfjMA2Jz
OwauHq0eQDRjDHPMNlANstXnMfDwREXJW5N6F9ZH4gsBON9Uy2rZx8K24NkxCONzGLkny+09GFi0
jD2EPpqkZvq3oSl2XOZg8qiTpEeM/oVwuJ6TMFyu81f3Fd6lj3ZVG9s6AjwFvtWD32D6ur0g+h58
WcZWbM/7GuYSqObwYLk1rJzZOu/u/QTYI6k2smh9NLRac9BMW3v/PPK5NqjtSO4yONl/BSPp/bLM
r5yjwz9GYKlOwXDUd7sd9ffY1kaZsj6zxwuUI2eIzmSk92WZV79lsS3mUxJH+K/b6AHEz03rp6UI
r48TtwMWEBTSR5E0g5+Kbs4wWIuG0dUv+foVXRzW+CwEn0x6TSyy/NvRGEAd+xwuOgJoQhVXATvH
+ej+olEwNcAwY+XS5HC2xGOZf2r92fafMCLyHvJ+FVE6+AJCPTRlqfJa4HODAJFhFEcG7s3fBAnx
LayuOBh8Enw+wfe63Bhe8xhQzgjXTAuNmZnrmvTc8LmC4FSLDWdhMOq3zKkdSbGv4f7lVvKE8GLj
JOVI2G+cT+pL6UNTjzW8+NgRFr8mXT3DUH7IiMXRO9y5ZMdcl+qdcF4WqU9bYLAZVTIPGgLF4lY/
NJTVWDr5gWDl15+u7pBflZ14iQqXGqa1RYZT1POhdwvsLwyhF4YMnLbrlJ8hAS5O1n9AXZcRho4k
DT4glH7Ooym88/DAY8Sa/d5OGb1dFcYQY5Dk5vjrxMZhuHzq1N66OCOt5LUnqK1A9RkLQG9vbbGj
0nvDjI7rziEVltturcHoPc5kzbV98oRckc3FGbkOcXFcF8sgod1nUe1u89AkMKe0jxdW2voJ7gCV
Hls57KziWvsmkbPqogIm4XIUN2e8MFod3rndSiPfABiuUP//k7KOo3MWUDl5ytHaInM/TDktx9wP
kfzl2Ym9xq+r530J7QPp3Yq/R7Ms1yJlV5DpS9OYKaY7/T5lQamJ+1rviMHWAeyS2R5oWXPCoGY2
6MHl1bR71/69ukj7tOBSlBpAmy6pbYilH2m37fjgy2i2W9nQxz37xJyb8ZeVKaTzhBx/gFzY7M+g
TsWUa+t2wRZ29xFsNH+FE5U9b2Qzu5EAHhR9RGU21nBKX3mvIarJN3l2ezN87+wpZDDNZalzHaDn
YQeGjqEPgsNeo6sjoH7XqkOL2GU794eohGeLQmEPDy4XSIgwN7/2fFsp94HIu0ptCsLlJh0uM/9J
Xh1CKvEJxjFMZILA9FZ3t+AUgGtw6LR5bZBWPTSSCFNDM6YHyKuBUmpKrwTDwKjO+/NFyHKMuF0s
CvupvSsbeBFpq6H0zGgALLluesm72RmHhO7DiuoLbQaInRSSU1DEmk6KLKk8xr8SU8YoG8uuPhs5
EpDm+VonzRYMUmQMXxMc2PDE5Yr5Sxt2UT2JAb2HpWV5Mvxo4iHV3wX95456RdNZMVIcFiFImv2S
wO6R28kLx5uW4PQEfj5mCEZFjiLIoremMWjiku6Nbwrt+N/AUB3MPMdy1WhdrDUfqDDAGaNzhJxj
lXHg2/9ox8Ag+191uNz4jjtKx+oy282tR4EJFxtmGkodsX7KRaeVNnj0DSRhOuWXO4d7Gc8jOSfo
BZVYKZ3sz4KzkjRHUMYQOinohulDq/XrZWd3H8nI6tXXq9Xf2oFCO9wywtEfHxqPxsQeVYiV+3kt
+b6WMuUD+Etk0X2bfrSjASuWsf8foYUBUoNRinPNDxOXvJ0TXiq/HRU0lWm6LetFEm9Cwz60FpBJ
iGxuQG8MP+Q4a9UvJQo07KjrS8/h0qdIcbDyGEnmUUrT5JBpac3/Lx0Dy7keKVNSTQ1Rh/gKEXEd
1z7em+nh0sY4FB8I/WgYArccPP4XPAz97X6wAbae0ATGvFuhBBytTzdc5DdU5SpXsrEnaBpGVaz5
fX4uMbwxa105jSYUSIvvFfEirssRLurY6CgCezRBjcqGr9Vzyd356LFD5isGEkhYaF9FnUVaUwzO
fAqV9qBrWiAz2j103IHbIO4Er/mk6ygEU+J4dGFCp07WTYc8KzPvHmVbqMsCiawoeI3V96aIpFYZ
AoRfSDQUJLL5d0tealrD4vNs6q/2EUtSpjjlDSi9zBYxToJEU4UEkfMRwyG1oXtD9Q19wjzImGoF
/dNpc8DqLoTn1e4A0PoOz8oAS5zUdn85fjAXs5DctDDyMb/U1/wEZMvZSCwVw2eZE0dCXWauzO+A
A243kMCG556TsiAKx0aCJS265+/VLwvppcUtmELioP6DtpIhYFQkhbr694NPD4k4pyomDFreJd7T
UGOBDzONliCmXgJgFEWF6A4T25MuXKgjIwgfzLslPITWv/e0HEgkOuCgonjpD3EIVZSzsASESPVh
zTSBT03IimNoriVnkf0+GqKdpXcxc888ac9GDFMXO+dUNR6BSs684ZoztCmmHn3o/vTBn7qZVP9z
m7soQdnnB0J7lJExZW/ZpIxB63k2BK4fYkWGWkKCyuSA1RW72oHwLidNY5FJd98MAcfPY+nxQioW
nxw8NqrU0rWsJFPyI0p80t3qxqjvB2Cbg2PC4xtrDwuA7g31T3LWJC8SdnNM7UNTY/TOP6Njzno/
wB/DQvWNSazCIu7efpukeJFPMIkakFttwOiRmtl4b4d4bjEIyFYuPsJByOKTpp0jw/5uOh8jCLOG
s5gkivBLDG0Uge3JUrfT3ec95Q3vFHJGm8cetgnZ0Llbs2xZs2tDFc4fB104F7z9TxfZgRMP1QCk
mKKmL2CJrt12YdvoVi7YLYwVqOQe89kFVI/HFNQgfiHZnNEw57ZzdkLmcl4t54e65kjuomtobSPZ
lmuu4Ea+ANx1zGiM3ZJIRVMQGF7Ov38CmlG1a4dqjn2AQ3dtTRvCQoIDIHORhFEt4/mrLdRfTxx2
vUD6e+axeIf9Lc/wIv0NPg6DtcvEkJ6Hc1rnM20TaVoEEghKB8lRUS78Wq2g6AnG/lBaxB2ofNvB
vfwZU4QmF/BRZPlF1vAnlb4nvJ9a5MBeoEya5K2MyQhdXndI6fTe4xV5RQzErZyLtu/QPVMHfPG1
j11qyFbIeJrlVOc3nAh7XaIjcv4eF+oYF61MV+b5mBU0Tj/9thwe1vY3zhQnP02qrYzLtxoYciib
8ZQB+7RD3bNKCYvi853i6iKEGATCIi12/QxR3RSUtsdyldm8EXUcxCDASDtsnb9RJQQlRTYhPcIL
2TxEdjNz/5eX2vaiqOaHzTfBJQs/dS0bLoJCT3NL0tCobjuFakFGUj7NhStPHVCmZApNdCW8pZiz
y6qyD0qf6x8Jo94kgxyMfsuZFdVrXtgeKrvsdUlH7jPYkZbfMU7gTPBNHiZOOseS3FRctQMi6MMn
1vEbBMDtqi2bwJBZ0xtNl9+/KzZbCpKH1UESFjn7IELLXrN5x/kk07Lk1WGtRShvCniWb64KKuA6
lnDitiBXhVyygw3KQ84ChUWeoyl60iLimcBXr6Xo4cnukMs9yZP+msgz2A84ktvA2VZFFppwwmk7
Ry/6VcbF4GbKhEqqlNzFfxp6lGajkup6jTiK5kaet0uzy8ZacIAZJrUc6ku/Ue/frbM3e3tTzJiD
tffz9LGQ8NZGzsd3j7yjZUNhCQIAi5rLWhuXTpfnGLm3/Jh4n0rh721EvFD9Hl77CmVtPCdaoVUL
pAdr/So0fckYw8Fwh5Lo8Ngt/pPs5K85QtYicgF2ihlhxRVk8+3HSfdO68vdIJLFTpmij9b4os6y
kETXjO4oVXWvmVdZB30l2ij4OQEF0jIGoXIG+wU15rhozbMOnj64QDY9Lo07wYt1MRNk8cpOWpeo
wsKYYzoe8+QxACPSi5/pJ4OPX/zK43fxh8bisw3Pidgb1lvksoDpEJRmwcDzQyq5l0hRVKO+KsMb
Ve2LjJ5040d+0O4R1+wPdL23FZOMivUabMtnUeRCiLE18NZCQWrPqO1xPITB7c33ldkypFn8r9yx
AhtlRWC2XU0tM7XS4S9y2W9PzGtL0yT9X4MPeeF8eChnkUDNheuez82BOmixlPkS6vD6+IeO9mfl
B1jCvpMwWq7vIoGTqwW6gsHFZCy0ABX7mFFq2jXn4/1pD3mp5I9Pbc+ePQa/g+bDP+WJUmVnJedF
ocuMu5jtBqvO6zZbrkwn3YPfE8BBMsi5/20T9megyqaAmIpDqiNy2N7M3R0ewxyBvoEXHUa693cQ
nYS8TP2aVdo5B66yhNxglyP8jftulU5Eosmqz/jdMFr7Drpok/mZaJt5p1qhucIm8X9W0l7kVxoh
g1vXo58XlmnH7EiCeNm4KgXFE2g73dn4p6hCLFd0j9fvs0ujl57JFQABUFvyxC5fST3P/QjxfbwJ
P52od8JfaaNIszDCb25v1uCZr85minZT/k41L5Z+Uru+Xw/Y0qm8WvQjGpVQjc/77Av/O6DzAkhY
m8UHzD0bLySQdtH0HCO5Dm9Wsi4SKX0Ap06bopwQ33xR2/e5O9+QOy1ghWVqcBqqho5XH2egx1Hu
xWq4y2hbWkrMLNTZeodMXNGrZdi1SmVTwfFLarmWQpIU98TCtt06vTPt6o918wmiJR2sKukMDVlw
5AnWxJ42Uy4+n7j/4W/Dfe9iB6yAtx+qKMKxTkJfUL11R3uOOO+CCO33f+zejNX4VNqj97wQ7VuG
kEN1ICp640tMA98fxGqJo7Wo/wUIm5NENZxtD0c7uIqiLnGZnxnpIvQ3UcMBHJS+YrTQugRC+uVm
zNhb5B/1h6L3iQJxrfPNhxr76pv4X6LyIDOljqmxRF+Ahq4QqpL8DfHbx2AOqtliuNDYNwrf3gNl
DfWE/Q3ijEt4cmbRSd/etlAulKmbynhYsp1w79jOnyUnUh4ZFhUZDkXcQS/d/4XgPki3k10qB8W+
JLhgruHwebbd2tq+zOV3FxWlT2LKhNalAPA17gydMKOs/4Cj3qlsQha40EeTRyp3eeqKsL6mgq57
+7wxHW0pQ19lCyEAVaTiJmyRE9NK5R+Z5Xo7fU8Pw+5kXcGf7GZmjDQybUv5POq/m29s61yhv6hA
G6HW5cmxA3f92RCvCwXXqGX9pzWL7ibrr6lsIKqaAWUBrRoh4FrFhO0yE9BPrTbl0u7NRyoDPeyj
HhbR4aWWWXXO+ytttEK+F7MRJ3UcUj6XWNQNcYzg6U5idcJMzhmaSkGgTXlqL56qFF+y3NVjgdYW
j46h+hVUKhvKa5ywFTThPAuPkMEDQKcbk00GYVplLzhO6mVFfkGzgDcek34wYGX/8p9uEIrPFGtg
pZLB7nm1MjXZDcYpV/hBb0YkqgD3+ugrNAzgdU+AxC3C3sT+s/sKGyjxKERCyWpDdp9YVXXEYIp5
EzTegNe+JKuNhdF5Bl/dhJWbW2S45WH9xP2yZC17r/yI1dHk5/wAt+OaIOMWKit6F5k6DigfeEZ6
o9+uewSZ+WaiPywWnUVKKKzQ9DqO/V/61s3EahPyYILBH7EnwU8bxYiUUXl7n7V1Xq5i8LwLvEmJ
+qGu0Q79BG4yC/8VnhRnl5JQosBKyk02vBJX0PpAkEn01zr/aLqM1yg4Cm6dtTj7PcFwlwdS8dKd
KS3pk96SWmxPNabtul+4GzBx0HESA8MjncWrj+SCgLP7HSV+pTo3xA7GX5nd9Wyo8SUKo1nqCIJk
9QmlXjrXhwTDvV6N4xmjvuNC5yJrT+uRMDj1O8GryiKRIodk4oyngGjfUC59GdcBkw51BCiKmtsw
pO/aVsHKuh2/wuUKq6OHNPo2fu1LiPvaQ7HX1XSlieQCJeUM0jkNMVIKzEpy2LHwXhvovUUrYdbJ
dSqlgWqWjrxBgUpyH37cBwIO4evYcNwNsz7xKy9+h71sq2K8vyO3W2viOYZYtnI7sNSYLObFHKJH
UDfQHCEf3IxmcjHHqJots2yyBeFkbvbzzhPouhzzDwZowed7NJJJvXee2aEzEXn75ov56YV1T9x8
XWjrGyEZUtTQ405tXsgBZ/Rc5lv6itTif6c/gys9hMO2ND6jlm8IUfBJUgYjNRSs6D90sklyslq2
P1HSJ8in5Qip9DQ1ONaCphDjZ9sP7i+OMe3+ytALcVwzKFqoIazXxfIzWclLpWrXLums6idlhmS1
XbXpL8kakIzoIP89oSofTlxT+rRcBwtOZaDz2JuCeVKReEvx+8wOUnBYVPHRxVXMRBD+6KAh4NWr
xoYv164gyrIi858N0XJcKyT76n0UNBhVcMvQKEBUn0lvO1Glb36sYePL9mLeVBpM5PUG7Lw6jr2t
e2LyPGQC2+ls9kbznh3OXA20hRvqOVKk2Pjj6sQujt0LuTQji0nU5BjzN0tT4Kpa9RbxbM6B4E25
OwJj9na4PnZcV6fIpn8SC5GMTza1tRRFJuqO6BwqXqnlzAJnWJCMLZaNOsk9kkzCpFX0DaXpQ5yj
+yhNIAmSjwhgpBLrMRlQCI9vGtbWScGIXmXrwOACxFOoTI8xL+J0kWFh4Lt8lnxg02Jb2R1QU8zx
HC5dh/RAT/A+ttRH7JFkZHykQvZNmfWFZ4SEkmMh8BpXYPy+PVjE0+2jmfdeVlaYlMUdDMnlzb5h
FSb6/LZY767lck0Ak3QGi7YCWlhlWEUbrQnt1Pd5cuk7FYP71RBbNUTT0JxOFQiFqDWJXxGnbI6r
MGH2zN6ZDkwgZoeW6qFfGZEg+oyvi9UN0UemkIJVwW6z7il2d537nT66xG+X2kp31UtaL7ag3w92
z6aHDITsGEBEj6MR/p1/Pd78t8xTC8qB1Y629/42JAPa0sCz2PVWRmQ+WY9rDHvpwugM52P+vBiK
lvo5L/wjqSjqRFCR75vhbygYQlj1RZtIrxCglwl18kq9znjoNWP2EPGJp/pkquSVqeu391+M6LQl
+N8igSItMYH9KKb1mF97TtFnzjnRxM3e0+Rty4x3Lb8puIOIWDkn13AJLkq+wsYgkoT8SK9QfTuB
gTY5K2kykDS3hljMYU0RVJs/sEu6VH7maAcua4AeOdE4e2G5ZVH9Ndc6jBff9LZJXrLPD5FPd9dl
W4OOLI/xDu0puO6/utsiq4MYxu/Ka7d2AZ63y4NQka7QRQlWvPHGAlGMEtZTiErgp1s1UQ+oQ4wH
/OBg85WBYQXsJiylvz72qxliKNdwxDqt5kpbQVgvCnMNkZGb3U54gB6NUlrQchYa1+BGR06xcW++
VbnXC9mJ22RZ8EroYMT/sKcmQcIlnL49oK2vXB7NRZWQ2Q0rr/VHfNjcsgf7qmL/LwU4GeHv7g8J
1bnhk9i/eLkUC0eWc2GCzZl4mObw0DVVrAfqjqQuk0HNENznbGA2lqet3w1XJYo4suYvC2SY6Vd7
pTBF5CyEICG4J/MKclF6q6UGt16bW1eyLGgw7TT8M3oAtXxl0hE8/T1ofEfzcuWtaO/yeFOII65Z
ZPCxflAJqtimiIT5bZygIHQg0A4N3sGbHz8oSkdeB3uT8KHcgXj0kAGjahJgaKRKQVSz2IMkzzro
V9oMiJhJzkkaU2wECYC6Dc0GNroYg1IlCa7c8/xbS07/IEIiTCV7ldqVKmxAEKX4uruJn6YRxvPs
nFv3z671tI5gkwA6SGT2rD3t2CLwyohA50+lvcO1hA9/7TGnfF/iRtFtEw1ELd1gCmgGgO9N7dHA
AKBpCVBevvdYirt9gKbHNiGScNMHzu5IZftw1eU0EU/W5BXhDca2klBVOzX65otiEAhZJNO536gU
f5T0Li5yRPK2c3TL/YTKyMnlnrE0KFWclThYyquVcATsPskXmQ0wWnBHDpYe8XGF+xmJxv98hotn
vvXmTpa1PlyTKnI6cq5AkSI07MIGoPsLgdJHo2p8W+okjDXnC6AZorOY9LcuckES2Uw9Fkl/W4rb
X51FDImMfdOu/Fnnc5Uahs9KyurhKS+COwHiiZcArz0h0/vWnGl9iv0zJK6OY4lgc6rtV2YeqDcz
dxBWy55PUT4IHTHga/uPN1ROgf1u0kNCD9Ebl4dkQLGBREe47eLgJq4s6Zs4gJRRUrydz60v2ynM
eNlS0z6lK5toyT93y4JumrkLP6Qp7btvRGvRu++zs5+FjmC/J0lniFU9S69WVT36zzgUWkb82xXA
eQzbvlCS8nz11PF5nrIpzON2+OO2v4fS1nnZLNQmEHYkPVNsSBARGONXRfikswzhR7ko2cM599rZ
EDsFFvjsPCfmxDXzrmuDeMEr/+b1Pu63mO0Py3NpH7m/qhtEZ2H61AFTECDvO5YxMcMxxmRMfHpc
TpJBlY/1RRP205jzse1oF4UzlrhBcOcY2Fb1aglRAwvFXFiXnnErbvxlJ4xr53oTa0lRrI9ai909
t+mEorPhefLxYCB7f9YBqC16ufCoamZQ63I809mn5KLlQpX3sYIxc48OTaGOOYqB+G3vIkkimvKy
9surXkbbUyEYTuDhi/RRde0+0LBsWE7eD8pPgX8AmjMqOPSTW5a9jjacmhal9YbXF37UW5TI2jtA
ijdjlYuNJYwCA5S5tjjYM/AKY7pP+KCNHbvUjLoP6mJJLxqdlJ/EV2XEfXOX+XD2uZsLrAWWbqCS
BV106rbHG7UjE7w/GtOIRX1QXBronGgKhNIJXtdPZ2JdLukOv95zhr634vCGEgAxDX9qmwHS4ftG
a8i8tbdT3eRD9TK3ulNvsMZywVsJr5tRGtzDc8CxEpgar6u8F7u/XtJ1TaCXpStBYF8DatlzWAOk
M6GwZYllgYyJnCC8dKW/597oUAZ+gC3l++xR4mfhLesdG+vIShe4ifj5zE02e2Y4AJZzqrR9W6K8
KJWoBmIZAH9qPZTcE9Y/0ZHUKzvQ29n4rtjtBKCEaD5zHpqkjR3Ok9hYJCin3+yQcxlQtDDgvRqM
wPFOvwtTOJSZOAMsOS3dTfvQpXbdThSC/t46QhWLafv7pSwVMaloXdeIOPShtAEACie+lq/TCLB7
BDFPu6ZR1txSynxzfw1EruPf42bqWR6b7l+m1TjmptoX3pOg/YmhYGayauqPZ96puZlU/qWpb8Ro
7woM8ZdgfJzjtI+dzr+wO01mtb/2S2xmkHGUSlRcWBhA2fN61oxhKFjcNh54R6agC+5EpA8DcaPX
MpEx11OC2JCmiDNRrAmTUmr/A+7Gf6e5Ob7n+xF4v3Vg2CeN3MdqU9ofkz3RN3dNfBceKWlTlTQ1
NWuGIysNyYzHb0yeh701ee8vaVIWNHq+Omot8EeyoanjsJq6i53cyoYbxgBTEE97g65dMb4hZ/bu
isZIIDjKGH7TB82VM2X4njHtJ8gUGOs8Ot52ROfG51eG+gV9uHB9zmNEaKwAPaNhj4UOA/nOuzVX
XssKm/rrQVYvWDvgd+PP10acy6P6nm9NhJehW8gJJaGNMbFLAejIr87Hu16Nd5F/UHqhqcHedfIG
KuE0QHjdGLiiUUvjWOR3qUt2eDfb/eJhJ6/lmQUqGijGqqnuCwQN+8vhfsNKcVOpd5rzb+gB7Sq3
Vn6rUyxZ5CeZMHm0Kr/ng6EbRjk6AX1wG0yS22wPUUHkOBoErbvVCZ+uLspH+ayGtTuojG/Msvla
3SGYfXG9ra2izQv4aPxiROoUQFlapioViL+f30a6sSQ5Ipnev6RDT24EE9dLT1pfqW2lRgk+QLsX
eTwxEaYGetiBYW638aP7hO0cTL7CBxc0F6fvHtTL/eXOPpr+vHei8wVxa40pwdQcJqUCr3QinAnD
l7Ep+5C2EEw4NlSNpq1q6fmY7qmfsVbqWVVDSWxWtml5aS/AlsImWLbk7b5ngSg05wkuMn//7oTI
2nd/XaYJqE5WNHL0uCC/gaDrtOvkojYJpFkIdLZkSDgDyoB405t13C1iCArDOVs3OPUmX8PZFVOe
wEevY6CNh132sN639JQrzCXyqeuxdmDk/UqRtC/mEMepaYv594g/biDEGjI18sICKillmLQQXbaC
e5Uyme8/o4N6jCojD1XpTfWfGnnOlsEVJwOYO35YzPxD+BKhiMmUy/+Szxl3l9a23UXB7GoMf6vd
eYbmOpP3UPdOIY0WTrtcgeZ/d+ut5FKs46u4A626xdLBqZISB9C9Vol+gECvqd46bMKxe59B5GXv
xLcF+2p3Fd64AOuSwjAKSIJIeoe88fMwZr5rkW7f4kp1clrhxKBmk57qOih6FIToebBZcupx5+Mr
tbMYZt38rH8uuGY0XA1cH2teE81toiQ9hgdSvdkdu8jYT8/gZxd0Odf/RYfANPPeuEc6V1HK9/+9
p/MbcIh+XhoLmV3kqciitJzOjfu3IoLA+hFN5kPtYsXfikwR3H5NXVMb1Lr9+Jc9kkH8dsoQduui
ZGewRIs/G8U+IUO8WWwwdatgswg2FlVStoRN970nECWsRYVFfhEz8i4AASnHczobxLRbhwbKN4+k
AYs1am5rDynFiBIZspRPpevw7ODMsc10+bC6AWL0H56nzu/sQ0BbK2V9qLl2n1SzDP8WKibtprr+
00tQkcdhSjzJfcnXyHWcfrG3YTqM5tpWuyP0GuCoj0t15itq5Lafx5o6aRfLSkk56coIZk9eEaXf
1pxrpy5p2bVWlP2ERdYn+15stPzc+VkVdr37JXt95C+s0jInok6cAeG/4oVtsZ7sLAym76KvVHK+
IBLNReKqp5ZrhnXOfYdkTgRZk78s/nkJpjrWuHd4lO1Sy/I0z86zc6b70DUtF8iRB9CCATM4Fhbk
Mf/94T/m8cTwHi2A3D/bDb9j+fESsWcw9/DO6BpeQ/Nwn/Ea/GTe19jWZ922T7wMrYOZV4d17tEe
k1KQs3ih3l6fVUnJAp+9Qr4IFMAGcMemSdqTxSHa2sB5V8/wpQ6B+oV/ndZ0rNynStZ+9wDxTkG5
DSRLtyQw7vCLq4FvWeyl3uDDs2J0D0I3kpxtxTni4KTkHl+52ga+e5RTG5TRWqmobvNYCGM+CdYQ
/UeskQdndM7BoCW+R0SSglUpMmnUBcd4jLFJBTwIxItT6GOjypmF2T36RJMsho60iwgMYBTZWobS
f1XGMPfTkNAy+m0I3hd3kT5pni8nJqHjvQmJz/VLuLQkidWUlDRguuRoQQ/acf+GRhbmx5wNa3iz
VIznvvI06VO1wIr0/LS2r/mzXVa/v4LvEXlK+7mvO9zNoGzX9aSPvvbpsu4/s7O/9CKUxl7DsYjS
+ThsnLVlYTSXcuKPkSig0GFb/kDBuiKhksrtBDIfjhlcOM8WGPC3kZ6Dajo1O5lUFFhx9Q9mV1RD
nW/xukSbWjIWd5KEp/KUsocC/43N9YRGQ6jHlEXWhy1Swm8W3NCTHJZlA431t5wkl7hz5HVHmscQ
i7zDzwLSeOCk0Iol6WjF/E+iuyD3vcXtu2PLCNuvk/T6mFQrSv7w2amWmCSSLjK2rKgqJnv+j5ZM
i0Tbd0QfBXxzBqcv1WFwknbRibFp4mAjWsa3KxK4eM7oxLqqoHpK96nlF8JbTShdvrFHc5PsChjs
KrHCI2PmoSediWObxwWRykemhhnXYuM8ij62ma/6MK0DyqhmAHBE/Af4ZttqY4WOX991i/bW123R
1U99cqnfeFYi75PsarxEC2sxwcwbfCGc01G2eyn9co4WoaXHy1Uh132UosQDjMv+BP02qCoXn1v4
8B5tvwJ3RYe4TRFdQLsLVwHY5P+1EOvGNoCxeotG65egRPhq16I1ZMJX3MW4uzWMFDdUtFVDuQp4
DVzEK4uorarKtw0e+DR0oN+FzrcSH/r/S3aX4Uu3BhNmPA9N8sBMJexj4e5mPIiYNyEYrxBfQ26t
rsWXKMkr9mPavLvDTiVp0XAsASKkNJAMCj+VbkLd08QpqjcmalQ7za0wMq4pNOfopXNniAxxbvHG
ZZ9bni4/EZONiPSx4uT9es13ZIw8HWSHJJSwdSQq7F3HtJb1CVuxhYHVQzGtfx/usDb+sERtmoQQ
FYCx3c5BH+ACC7p61FIlSyg7GPQVPwagz2r7oOVOM1+aJqqvF/rXN+oVfHI8RrM0Q+X2cC8XExUn
k/fIZpNZJ2R/jUdut9hTsFbstR2JshRATFmfuWYoriuN66N+FFnloIo6MZqa0hlCbAcsvMQ2iGI9
MJQH7REpp4qr6e/+crJBqPEiCCF1aru0hNuNkLnBiKkKGACIpzyqJT0gZo8p/DR94rzr/JNjMytw
vgyY/k2Zrn5Id4rT25FS3WHUj0kZC2ouX3y9z8AUu4X2Hi1ejcCDb3wI6ePKq7Yf1C5zzOzJv6cy
sh3v3Mb19O6VJ6GKD6lf3p39TpbFs9rfQFbFcSlIaTjmxKQexCbUJ/P0UlGZRJw2BK3nXoQeUnq0
vvNgXwT5qyBPT+uFnZRsZ6e4CALDZ1sF5eIRk1Ewigw4zaFmCCP5FcO7t3LDryrSQKoqMp9LwGrk
ZZ9g+FzFYxp/ZEIAS1iSkTVROGMrPoCygi0vFgb6l3ivQcmqmk+DDBcFvZ82MSRYT568X6fMro1j
WZJEwcZ1RkNJFUzBcVWprdf5L5muknSIEcywUyW1kI9BIgUfS+5nfHytcG3ZErSuno8kTaOwlX6G
SS/XzNXMoSR0dIVQFa4oy2mFMU60hDz7HFl3NbPVBsQFuEVDsXkjlMmfE+9dpmlcee7DCR3i2E0w
zCElrEcFvkBvmfEu04PoqY5+0DRf0q+QgeBld4z5yT7x00RIpiYrFrBGNLNPJ1OhlDFPaWvNXuY3
+7LGMkr5s3HOabePInMCIcfY1Y7QcKcU/SSgutBlQrhD3A3OuxYw5klpglWxvRVRe8w//01C9XdW
Uy/ykxtD7iD+3YzFwcD0h0V05oiyibjCE7q5hQ0tibtOpSvgclfUhLbsPgVCtMB5IQsNNx1TC56m
VyKlMZZ3BAUVYntPw8An4RLp8Wvz57zLCgwW1wd7ktW4nFmJ89gJzFlL2tVhZgNjqbN9eU6QGmto
N8uv36XJp8KyJ/P4Gzvdelk49QAtCV/Uiel3LnFpL3KSDw2prRtmWxMBxuDrqVwFUfkbqs2hGkF6
OPkvn0poxDWIRyaHewFK30f7/WRVRIYgtf3ffqPNcDK+swl7g8L4tNGK+cQSzs8NQnxe9TfHSdmo
MccAl2YuqGkkLRs/Xy62yftSL+ZM1s/ecpQ0lZzP7DDG5kmDyDUUXjodDnSDqJZcMTvmkfo6s7Rn
wVB6DHksa86Jwigev76IR7JVpJ30qRcXkSauO4dTFBO/ZcQe1+fWaiQAwzPlMIko092o6m7N5RKQ
j20wQedwwMw+D6P90dmXdZfGm8G4Gcu/6m06wRDMH7MhOJtRwj7wEW8IRljlfXDOW/3knFWnQXF0
EOGLJF3HsynHF6+UFlQH91IPNFd2CqZpFCfF52eHtnAcZocJFLdMxVuhi5frAXg4vnoeUO0ixOBs
Ha+tojrmtQMWBha2PA1pFF8xi8CaMB+W7m5XjPHykI6Wcu5esGVAvRL+i/4d06gEryEpRcL+y8bX
ZCsaoT5Ds16JxScF+troYWfd6tROZ54NUuNvLwAymRLLknl1yeUIl+31VrOlp9xI2MdkXszEUXVz
afAqWlhZQeEj+m4neSkVar3vyFG3qvUu+aUtutr1QLXtSWvNU/95iq5FS+lKBdR9iHy5CpIRvnX7
/UkwwGDwfOX917KEnPsElDOsi3v043ykMeN+mvwwYp5a8om5JiE57tsqYAMCWnjw11mfbKA9YYw5
kKHGYZiyb66y2yARxCI9EZvhyKF215z3fOxw/ZPLbIV/zvZ9wNGkjfIUqER4YgrzTqRPDQjwiyEX
Zpp1L7vEPvUQ6+PHXwRp0cMiAj42DeSZDQCuYr40xSCIrsJRsImPccFg6CfU1K4Jjqlk4e5vBVQL
KiD0q/XyG/H4BZGzDJ4lxLAstEWQ/Bt1HEpNc/dHNG7u0V83KIpiKHTXiY+603QoclnFNaNFHC9g
+QpKciogJdifBX4tyY21I29g+e5UNkVdH4KvubNZisHHn1FJ/s/amSAVEyOp5p8fmxf1q44/TvH8
d6GFIjMI1ZcJs6OWkC2d9PyZF5ZIg4hvuVakYhACMWbJSo7y8vjvv+CoP9dv0A4hBtfO96cJMbor
xFiJ4bGJOXByWWaB3Hk5LdCpkiMRWesH0FU8lAhjhgrhJ7WkxzidUIgh+PKVxFv8N/WBHRVIxYM0
H64Z859aox1Hc6sEFimZfDE0W6ZAQPIeXLO22fmyqHIt1STDOzO1yu5Zv6tsUT+bWvE3cLgqNkKf
jVOYcMz3OgCDw7bozWlB27azDGKzWucWZA2VNKaxogH9n9hEBbrXBfPd/T96yymGq0eTkncfhUR4
DOpBg6YdxGeuIw8bUp2cxzlg0ey10Wf2+RqDPlT3g83t1Zw5aXIj5AqtkpIx+xvc5k1ub/oo/scn
vBEgyBmRpCv6OtN/g9UC5mZytMNaC0PG+DAqnZiW5iI1O1zG9+W1LxcoReKPl/0cBh5kRTpg95Gp
tCrVvQ2mFgnTpgWGw3Dz4hIZpkqiZMT5jo6b48kRGptGxdcDx7L/0WJ1OHvBusUtLYKVFZiNkwT0
Ecp04iXvx5YJ/tdVIjeNVp6n/ZRGzXQ3K/+1HsYksm8ZFZGb2L+taTx6FwSEIghL4PvFJUAbJh28
s17wMvhn41fY8ULK+n9/FodxOL6p6678HqANhwex7jTp3Fm8XpEotP1VkPpv5trN7vqmLLZXMjjy
4xaZbSjqy6gKimOm6CzQKhtffbV+famwaHVjj7d1U79PPASNJxqlL0IGe5VTWVeikl88apPC6V9h
9a2Sn29hf2exxaulbdtbd0Iz2oM72kGKUn41LpmJKYm+DwcY88dbEaCRM6VDdQNU2u4w+zcQSku+
vxbrabRGfVc5DKrk+2fmRqGclbElO2eM2ug8YHpFpoWARaZ6dmKpq+tqP85aBF+AE2SbMRPsg1wU
UcxASC0kmZ1jZqiJjPG+5Ov9dJ/1/7M/PAO6AVSch5PirVvnFTUiGiHXnkG5KziXEpvNFM1GYKZC
Ibf5LFFK4qaJ0KOV/WfsLpgc9uzygJVZ/920QgXcEUu6pL1GlELSFIYUbUsYfrBTD1CD/AyT5FhC
E0DZDEKCIdPLkCb0N99YjPHUq0LTAb2y1uwhgtv4Z/qIUPFNTc//CNfeJ18+jtwxc+7vcTWwvX/P
lM5JmvYlc0K7pVW7GxJScHsS52tKfng0PF8PaulLsuE1FFFFEIODUC31j7uc+gpdqxr07OavV2Y8
ASme4229G71Nx2ocKJtpGw4ifzQMpuJB56/kXuN6EA3uz1OXeNsiwkmW2/5QMyt28u40VBKKO7nT
e0ecZLZ/hzC0tZPxLeVMLEKHPA0meqNWHHquXJn0NNmmfEtu4FOGC3PtMaiXDhpPddinZ+NLkcf8
TOUPWdWVrPKGP7ALVHAxhjlGAocnGILag2/syZPe7GodbYHC/06rHZ3hnKKInIIkUskobi6FkCY9
uEuz4Li9+aLStzKR0jBCaKNMQpmJHGpIKN1pA7GIqa156Lwk7NyiNaG4rGQV7367AeukfKgR1oV5
FlDEySFuOU5R+n6lOpOOguTdPZ1aFBFdWJ562V9Rma1/C4SEhz1tmGn2mheSYHd+9cs7yF7RVAiG
O/uLgJRcwUeIqsNQh+B0Lmssr8OYKY97ndkqdCxpRUJb9bYjCuKciplyeyNNuPXqInp/4iH4g7WE
8RKcLbk/3wPrzi9jWWpdiZcGl+cpZnf2mE7OUAcg3SIYdODKJFmImPovVFEwErNRd3eXqxv797Of
7mQ4w5z/Iv/CYWSlZBo3AUxcm3WNSzJ/YvcVP0t7aCF2oMYR8YKVFESbYEZA4ymr4OQ7vcyZot9X
7sDZBCNTKWW2NOjrNkdRULkiSr2Y+Zg7ofdmykKD3plf/qA6BpQp9HwVlKK9TVrOCPAjKxMz3nkt
0Hj1qgt/xkZ63lnqG7f0a3mbWXWJVRJWt7yn0modkevNnSnW83DU/AFsVe/1lCEaSGBeUEp3oXex
7qKboZkkH0XwrC0F0qVJhVfYmXNkobMsvatk97g2PTKZTeHT0fIVAX3caWSjopz9zMZEdx4pjjxQ
4fmODIPSmMWSewmb2C5qjW7SIYP4tc9T5Xg3sNpU2itWaeFZs+8wLkRZrwC+mRCzRLV+evvcMum/
j409+OJah708UtxvHjDgDde5V52eXMeqnhDFdSV4nQxZ0hBOsRx7xMwqtkZDWhkAEUCef9tgk1WQ
Y5Uj3y7TaJtpeq8hqdNPH4AjDrXDui2egTbYkX6r3RzaJSpUUuKjrn7opuNCU629vOhn0gGJQh/L
V+wS16S8X7WlcSz+1kz9OEjqa2M4lU5RqbJhDLpDmdOfevf7fj16Oo86aOOiaikGqeRkm309nTRe
aJRLGY2OMy+4u91fsa6OmUHWOcjl6ehvCoC/OIejNwlPlupmGaHpLXa80Pey0JPWBIYahHE6dSYX
BJuTZkE0Sy7uiVO3Hv0jzcHkdliyoS+3dOqC9ZjiZ8oNTf9zD6723vGMqS3drzBfWnMvZ1xf12FB
vRL5wDBSRWpPGr24dq+KHnY0KKdYXhcm5WUVbWm31vNgifIFeyHhUq0QCWzoGY+/bPEJntj/jMsY
AhsovK8lUIPccNGh6fyWyke0IUG0p4mrlxxNp5pkjC9uQyMS8o/XI9Tyn4sjwsUV3oK9McXm/kAW
MQUbKVgNw6k+Nrq5V7/Ec9W345T8YSaJ7pXU+jrJ+WCAxyW+zpUUioveJYrypldO1f+ek8iM6m94
VJ5bnjQjEggQvDjnEs3K1KqM1q/ThMWJiGdyKCjYX2CQ+MH56BxoDiOeuIvyVl0sAMpvNbkpO4NU
+LKxAUyUAfGupfeW7Pex8MH5Xx7BErmjOErohNPRzx6tmNMvft0/AxlvIWaHQdwhr9NdxMsHLKQj
V8zOLh5EKLkHcwZRKTyHC9J0Z368ULjaPksvlcJUOpzMaJTTFqjbEps9ou1mboWTRlUBnTFxNhJ+
GkgJIJ6U9kjCaTeaa6Yn7wnQFQCr1+8ho8HQTSUGdwitBGck3P6DQS18zAyvuK6An/62lGeDfX17
m5DVRzp3KowH2PMF+LWcExxLU+obqcZFvZHN1NbjFFaPZZEzbLLIXkA25jj4405pgurVi7LaExe3
S2oqRJrnzqHEk4nAoI/5fn2ibmshn7uT+JPtAKsiHchRNtAIKVGu6XdVyofCNxM8sN3gWmuV1O+z
sMKDtAmGlT9qEU4Lqsf+S+asCfELoPP0Q78ReiCCb1amPaDwy94ro+PURah3p3oOVtGR1vlW6hkk
1vw8ePdFLshlA3yLgSHD/Sgg9prDO1dZUVioAx/gHb7HErCUxVfuZ0GOw03RWNoARKDZeN9ySH52
Cej5umhNnM57AVgfa70q8JCfVVv/0XVxCARhz1URmlrqQKuKOA02p4yiAIwkwWCRjq42V5yM7BKj
GZjbyepk4odGLi27nq19ESu5FTXdSudS3S7TGklXYTbRbvd02fkZIcBzemmUzPv+610SZHH5t+GA
YQRcKTXjNotgbulozV7gypoPM36OBiRjU/cJnWin+am+ME2RZGJQHzKzCqS3PdszMnHEsPeWC02a
AotOhGMVzofQFsiLJAPj1C2U/xP2qS/qa4MMq+TWJC0xE8Z/aVHMz5MQAVZ9dNatBti1qLVXHdKX
d/7kxwRW+6JRpSGAXTLwgveS6imm/a/0K0SeTw4Aa0iRgKY7HnwqPxsTYz/bDS5amNYEK3THhpI9
UctMkK9xdTX4d8wgw/T5KJAwSPxzVVdxU79i7Fllbgjoqv3HvAUnNGfacjIZQO7rLyAzRT/ME5VS
4R0PaEONySLs7GnbuIGFkkaOk0XurUdqr6rJV7Q4h+ymuFDMyNgmzEJNyK/JRtQ1wb8qbucuhRSw
Swe6zjrsdzcz1KyOr16R93jDuAIMesrFgROOkHd3uRhSDVfHG36jyQ7HyUKyvecSX3PvnMCT76an
SGGJ4T4+6hWdc8Ah096aaZCPN44Ncw78LRud6AVF4qLLpfkRDdU0gkybrkkrN5+BL0Ax3KOgqsUR
aMxV8oU2rdsuhxPed69x2afZJ1n4dP43BtjsSQDYze8JGNchpU6X3/2oeuiip+OUFflDbpp0i0rI
ONKvWvGg2X+u6H8CtmMCqbfCx9m8MylDCzyBDXqOSW/GG8RavIqzZHYRy7wynkthNm3ZQPY+uJ+H
xjJrbCK07AeZ7PdcsQjKrCvmvPmlk1AQF8He8ytRtizAPOLdDFaQZNTNZrbotwfjfTGkyLp83j+F
XGs/Nm+pRvVSOimfv6cfyrWGWVebO+cHlGx/aSDCDzn1WpdHF6581EFJLJySM/5OyfiovjKpBqWa
a27sdTzVhrrzo8gTnq4R0E+twn0QKnEmK7Hb97ezuA+shgjjcwlOvn6AIMZdpXsEn+DEsg9yQbaL
7gEy5qSIwbkLxWNN/1GHBd/mIhTxE0yVtunhg96CYQLjlXoUKKJPpn23hYibNyIfqsJU2xTz/NGg
MY5t9xjkGKrexXwNSclFpKHjdQ+tSs68dPOxNZU+zw3BosUVte+ED46DZ/rAcayFpPCcjhtN61DQ
oPHJ1mSpadzw1OKKURuvUla7t2e18BOMu/B6qLzcmw13GZHpeqayV5wm0M84HVSFLCQ7Wl8zkkER
5C36KJQPlj6WwtOZdf6OZg8HW7vyFgBh8FdlefFLL0sSpuqzC31jQGYXETPsTT5vb9h0UPfDOsKp
xL+J4+z4Qo+dI61KgJY7bJpEsrYr3ahcu66xTL8qUY0j75m9nHs9Di1cO3Q6b6MD5MbebQ2jze0y
zVhyiyLfl+9Z8Qeu1DusFgCTetErcXgMHvAPXR5sp/QfcL6FUbd5oXpOFCeQFxrouYV/+/7pTmXE
Nu+5mjGTg91LcVa3Zi7pBrc6Y2/+0fEJaEe9IgEE2EHNa9Gol6ki9UDToPW0w5NRDNHtX1dv8ECe
SmjoyXiOr/DK29yeV9Nl6N216+J9ECgnLiSIZpdBAIlIKWKi+MCnk3aZcZyqNX2HLVCcbShIM7c8
pVIENJfjNT14vor5ELaNpSa7Xz4Gn1adhHzpqVTEWuSAd1RbcaKUfbd197nbKUrNZvlESsq2Jmvs
2cM8bvYG3pPZmvy2rJ2sqZ7uDqO40Ckf6AAAdlDdVa1qkoMzVEdSLgpSRdzZLrYFkAvkZc1xamEc
abWDAGPB9+W+injJ8hmC8EBVCH57mbvaY8o5TF0LYiU7ANR8675zo5j3Ndf7O5uLSUHjcRsJGKFf
sXiGTQMGwZDpWjQ3Lu4N+9cS/NpUYGJlMmrnLZbm/4hVjovnXFaO69pVaUHCKuzZjeTxnHoAC1Vb
9kOhZ2a6R+7y2r+3GgnisAj6LG2Fh1aWJRRkbIzXSxBfRzXPmkjn4JyLaZ2TF9jF9QRJwYCKFPKD
r4jprkd51aOQSNWzbPyr76d3vQubviWd2p339gZupPjrw01KBVQlbuBpl7Qkg6PJK1E6lychy/77
dIP8KMcEPR8Fgt+OzplDxF3n0jbc6e4enHHf8w8CZ1EEJ69kiiYkuqvVkndCPyTbakLMahtbIECQ
u0k+x7QSxcSsLWWRHQw6+5T15vbU8tzF20e5uhbuKGfi9FVfKjVLUSkthP3Etn3kQhGz5sudeFuR
utvJuXMMr9F61QU+NhIbB3VsPJ0NXLxKXyRm+qPi4EOBh8akxw2bzhs9rprN8YTq2knK6X2vLLMW
vf3GdN2HRBhvI1YFP8QG4pX4t9qjIO/Huk41L7rB3fPMuxA0not8XA93rvoq/6qiH5Z2EsLyyQ4r
Tf55DdRT0Tea5MR9LW+w6X7khTafnhQZrCwZ9bx9+UNQJ3xr9GWmn+5E/gKV+tRBq6tOYJdMNhe7
/Pk3SVDYijl909HNW2sPJFvRBczI7d+yOPyA65hpyiavIySGwtNjYS7hXKtpuAG42ESvx8LlG9mB
uCCGeXBz6jpEs3uSsQHXFJCTa+kagr+Xs1Npyhlpi+yWGGiNOVda5pzqHfum3D6hq7gPwFx2015S
5rltI0wt7n86xnoQbK3fmlc+ixOW54/QBd1D/0odlFI1x6BcAwYPJ4YoclOSDM2tNnH11shnyPK9
i0FMWpDyhLVgJDlYBWb37zFSfPQk0l2hpO2ceFQk8B6tVvV8zhH5ExXseJH1uoAuX3Mw1EG84GT2
27OW3a7WK1DvwntpSprU4ARQ0kXlUlMorCEtE6BVIFoJjbn1I9gRKsYKHqOxiEEw+1VzgCwn/1im
vDu6rRSdKc49zjleKv3ic5CNYyhfz7VRblOdmmdoIx3WjsgP+rZnUJ3/T9WL9FfjbJtHWoxa1Scx
RCkmdy4RynXQk1sv3hmGRhCezEs04QKvLKm6TxgDE+3lUgK5RM2No8H620UOWtK6QNUmFMQmO/ie
Pl06HQ3But8P9IL+U3k52nUJAynvCTpE6qEKLkC7v/o118dGbnYuz7+AltB4EIZ70AjZZTgihtGz
o0N3X3tWmqFJoO4Urt8XMBZWdP16czBsrZY4vNtZsGQ/mYRM2Gb5sPUiXJEIcKJCL8lfEaMMFJho
HYkz+FfARMmBWdQKepOyHzTKp8mYCDduizh1AElfxVrWeyiHdklGYxnrHLGETUqNcudeaFQ1lPAe
YhnCgIpmlkMtZxyArXnBlSpO0G1DEJHGuWe896/A+AU4XDzw6jsq3+94HhwVav/jQbey5F/4xm+L
siio8bGr/7qLo26iBh+vW8aofBRwqXyDg6ekU63+Xi0saQovmCSHUpTHv61my37+o967uaE190kc
veeH8pwFWF4ddCBE1OPJlxGwRR942Uvv8PV4CY6VjEm//IYlgdNtq1Re78Hbc1C5n5u6/b4xdMwU
lXn9Ia5jET38+OZU5m3c03DXyKvg9CQdh6oL/bqrsd/wEEX+II5Nh6QpM+6U3dN/CVNlC0Q93N0f
U+XOq6xnwjoQYQ0RZyVg1HP++I46cCObYUAs23qelEo7hBldzMrV9kSCQdD+YkMR9Sr3C8sk2d9d
k1J2OEFjWI+xRx8jCx63q2LiZ0SK3T3az8SxH/lT2WpmTVBuBYLEH6Vcdh86FEZQ8LMvNPM2b/Ix
AG2Id0dq3tc3MQpwlfMzxUtzEquOVv8umaTg+aYq9tq3xxWDx9wRjlMxoiQhXhqXtnLj9x8U75VT
SuDhNx2VuRPcbZXQ4efTPZajD6Y3RNnhPBpS/zZbpbrED/Bui9qgRts0wPbXYRBI8LmXY2lmR9aI
0PmxR5nXO7rGyOwVbw/PHlZGBQxjAGX/m3U/MHocRnDekAHlMmvwbigZ5DjUo3oRnOC9S+IQ9j7n
xSxB3I+XLg4UQutc4MvFWVGZwkpDDmISAcf8bO4YsDNKefx4e2CpQKReoacPgHiEcHxRmm4H6KD0
QNaKhVQq1cPqRyXOKTkLY5APIuMTqlEVwkeFGPX9jHOR+3kj4j644G+76dO/yViiEyimfAGzKF4t
jUrCAoI3f1F4YVyI5yrUdPGIYjAPVOkMv4+RwqW+pW0YXZzblbmqQ3WHXOP26HOWO3CuJrY2eFpt
vUMCXFA5nJGVbXk491B5THwQKbG+cSycs+V0W/SxnlcLVaBMUDHeDttvuXKe/4BVXnA6c4ciUez0
Ussys2CuZNKbUcjfy7rO8PJKcFQTBQPW9dLDzAOvjV2RCEBo2jd1kQftBKArpj90PgJ7d00Eaitl
xfy3jc9/ypClTFH/rBvBcaIdHv8DjHbjQrtqrbkQTCFykDZxVrsbubo+Ka3Jdd4B0SJtZzekvt6s
H/F27nvZjzdwS/A8dR9GoWf2YYCxA8wrPYLIySmH/x8I17ZEZ4LxS2uTAverqk7L/hHMWpyMf/1B
mn/SrKLWbm/CSZOV6bo6jxMMkF3uvrSt2r3SHISvHoJkn3rPjRGp0oeySVHVCE2P32FcP0XSR82q
ygfzyahvngwzljCU8FAoDfpv9hEdK/DjpFrL24sH6jTZmvDSFmOnWt46VEu9gk5rq30qdZyfxIIJ
eQYO5qma29aC0x9iei0ad8iyYefuYt/xvwHCGib53/xOO9lhT+qCiIbi++dp1okUjxpFfWnDe/5t
Rv0IqGK4OS9Tpye4qqbwQnXptkFQ3v9j/1EA5HAaH5iW8ks90rctg5scYn/SPJDBMQXjRER4kkHX
rtyz/JQzRkvsobf3yEYHDmmPa4Wp7/D/LxCtFHlys8cZP3TqgALxiVkQxCnCPyqo3OfXp+591dfb
nyJTWsUJO/T8Rg3HXoT5p4SSS+i0N1OAmV7ZlsskfT35nHVH3RB60RM7Wvw3yM+ry+XyfII/MraO
e6hOpJXnyuFnJet/iXiOU3fsqOPExjXbGht5kNqBwf22aA1u+Z+z2d0BBp5L6eGKzCAlZNJO8XpJ
QS7yCxq4IOah8EVpcXzt725NGn7/7g7cRDNAhb5GPGi3hY5s2qhW79klz+WDukxLTbyiSEux8Og4
659gXh47N7brq48BcrXvRp5rs1ILK6XroRkVO59tdNjy2cg44cCGzU8JnOFtMa5VPOM5FtJNwVeA
TqXEZ9sBHR+pfpJtzIyR/Uo1QBxxxSRFic9oem1jJ+2uJeyvRRGyTIKYjsKoo85opgviGwcoe6Bz
YxMuCmDqEa2TJLnmUsD9TA9HY4KlO0tEIxXsLen3rVcOJqykKCiyeq0cFQz5FIFi3m8zE9NI7Le6
/AnB5N7Upx7O3vpFAtH3lKmlWPO4CgoCW3gM8kH7KCGQy3A5s6QtMagrCo0x9vBFHfIxR2BcnZ8o
RjMY87dj5Mmtgd3R7NvpWeh7/DYNbJ+hXr50kMnI/ZlVG8zUEXDU4IR8jrE8HFWjG3hqF1T6Uo5E
XYUk5T6Pwv9ONEzLW5TyFDqXRt1BsG+ruOCnfye3fwDuWIYriiuwPC/WRrAVG17UXu9OEd9N6lfg
RKvFi+aiTAROU0Eci7I3FSRikLUpDLbVyf89+e/7fSuSIZEFZURvXciRgKXViaf0888D5EgKQIgp
WvugsOPwx1ufSuZpxMYuoMdKKYfVQvsHG51Rr2ytm0tfU5JmkX40U+qhBdKx6sep6458oYRnKw6s
XyiqrHPVkAvWAOjdC2T0OsjM9vS1vtIbaKRGXTFHfvqdH2/adwlaRmcJsni+4fR3rR7VktjvTnuH
OleyMnn00tXicJ0S9arcrgDtLwKbuswU1sehXlZ2OfmS52PUX/a9+QrPDA6r2yjdyEDbMWt/K0t2
fZi4XjTnk76VMjMdyH63QvXDNq5P5BZWm6ofV+7xMh9xRiSPl/ilGCnhVqb8J+fL86xASW2f1zZz
ZhV8uJ5Yz3ycOnE+E1oMzG4NozeaOzjcth7nPxbBU6hNa4FfSIaiNxIk8jmGKUAJjS39saqHonsD
PbzcD015W/padN1LIN3sT272WdXqe5OTiOV0Rrowd5K6gpr53ckSxj8gD7MbW83pAsPCILAXQWaL
ZHpOH86qviQxMol01k+HxUOVCbHteq+eItWqrSDL1M32u34bNEr6NwlNW22kXjC/LeUEpqun3Gs8
suOwnJoRkBKx+3WJbRZ6p311XGrWtBm+ArdzS/We7rKILDb2jjgwNmjwx2/YIsN+nVn8ctKVONT0
NayMs3YBX7IVnx+UxKzieQ9bANC+a0oYXAM6jjww6FBmDWyKm8VOenfeKyGl42pXzzNdGzKsU4NJ
4V1Iin00Kx0oVbKsjVzWeOXl5zMVIJvqZ64IrpWB8z447HK3HTxgma9hkeCllxVGU6WSLg9k3ayg
c4zoFxpp3z6wgKi2ja7tPzDh8nz2YEiEH1sjtBdSaOxwBHJMRJFIsR4JhiSDlDhulvVIFA+yxHM8
l511ZZoRocYzQMAvdZ33Tn4z0DdUaN+RYwH2s0LjCnukM3uGoLtNTQ7r8meRmfGUbs+6Vd4uNkqQ
F2KbMO6EYE61ijdw6pvwdesbZvRAGhfEKYRAOi7ZiPc//0ZO1w4HWK6OrnC/8RcJjEygPEUAn4sT
EKDWdsjbzxA4HOlSdrN7eAle9owpEE3dsDOle9367R3x7E/41LQAeDL0T2ZzYJ0+MHyIFKWNQxUV
c5Ug0ruJuWh4TMf8VdK8imcqTWUuUVpZjUSI2MBK9uF5pNrcnPfJ+GrD5YqmpDN++o7oiQhRBhoq
+qTG4TEZYmv2rfJq80NLlZ8iinbwvIBlvXmKFmWphwgdWoPp+YOVV7yJ8Vzb92D9+HCgkT4Lf5RV
Ui+7/JQ8tAMhJ8rwJHZwZ349UrmyvHR8nZSvXQuT/bd42dhRzCTgYnoyIVPW6PFS7w2S15nJVIZW
XW+iJ6VCPuVz4l9x6u27x19ma5/3rqCb4zDYL2BHnZLfaD466xtH94wqzkxqS++cu8O89n+6GCON
Rd1ZWttGAnRLM4HcUw4GupqIVS8OqFG7cMI52Qem380fSpWh4ESo0KJ8wHvoXf2iYlnMcAIvKnpf
eSQIZkpccX459Oc5sC/zilvScF5kEwYS/kV1Cm0eZ4GhRVjq6mba9hE2lzSqaboQj99RIUqSTCa7
D/OfdGd4iAoRs6PZ5331tmhPCPqxJeRjc5SGBqSiL6aIxhimEMlc+yiR2sb2vJIFI5mlLC2Fjwhd
m9S0lT30xOYU4NlQnH3532Cwu7vz8+tLkmwiQBpJyHFTCRHebVWsLc858GGl/xJFHOj4TU0dEWHt
sCTxNs78tvUsRzOelIz0MW28AKmQT7vvKTjKr/t2Aqal5+1YwftQWDhOsD2r1DJo+XcEMJTDAnzf
5/u/L+k5selg5mYYDOtKUKq3mFDfYeYFovXC95bQ+mldRlYnlIGbP/VavnpcQBBivlr9pFInvjeG
mS9SIWa0wxny32Mx4HW12dSrTodcM9m5bHcXy2egD9QFWj9XLwZ6dW6ouGwaiKflsTj1IEV+6JvA
UG4VPOXCjhlFL66BjsnDO8t4nR5q7lTRr/sHV8TJdJYjiCTRHtDFV59ujexBU1z+jAIAtSdwfQPS
tUtBJoF5KWYW0OYwmscSbVlLP2OPCZnhnLPDs5JX3YSaO909T9LFe/4gOVFRAGcMagGkuXqCZnWU
81ZGGUs5nejZfbcTy2QsDWdc8IdWQay4SyG/2gKiTHjj4CukIWX3LFqL2Jfif/uzMABzoYCNuUOZ
1EbINRGi873mzdWqtR93R/7aMpXwgz9ljltm3ZiTAngDKPyQW1LYu+frVEx9hzeGIkvxBNnhWmUo
D6Dt+f18ZoxtxuykFT0Nin5eOnLuo+ivujSqQ8hKSJmNnLRpNPAdmJxhqzvSA+lNDX3oNkCG/Y46
Dun3Np1Y3WiCVvkvVzFYXkMqBB8EItaBM052JiYR6jYaczBMiuoxj+YqPkWf9+7vqH3SpXsb6lCQ
JVD5XJ4XpCvQUAywB/BO2ZKJlxzE/etYmzbRy0ZBjHEpPFEnh3f0DOx2qJpbvmmXHnqenZwluNod
kmONhy+LJlAkQQxADWGHzX7oU/MFGfzBCKuV9sD+2Is5oYaILtipblm+UHyveSfr8SmSob4ggsix
/Fh9qHk0OeQzG9trIdgRwyVW2iemGAOfSmasJSkL0+K3Mn+5kdoszK8ZDYiQSYnPylmgcMWAV+yk
gQ7mewdqZZSWJC4U1AN+S++Q6+UJ5585s3Sxk+9zPNkP5EhlCGOpNy+QcUFxXgDz4VFfH5MGRYj7
8puEIyMmRenTUHM9DJvWsfmXl1fnktWWJ1lBofNx4k0r5tKgdN0Zv6voi5784cqRYQBhzRQXpf13
N+DO/i8mHz5+v1x7vEHiK/sQE45VhHa+ASAWx2Ppedm5yak/ymO24eh5WONHTE+NFy9BQmcnfshB
A/0j++/IzI5uRV4KYGEW4tHrGDl1xtsweebK/7Ccz6qwTHnNeQGIIrABJFHAxo7oQgIKVrBl4tSQ
5WrOLFIYVd7YmZcpsA2OefnjRxxCMNasbbY+hNrqW7VJld/oHFRPlhbHk+7c5e+NzUjS3UwWhALM
3OohZ8DTe6HVRCgTNoY14h79chTbgcCXHu2C1GlMzbyRTqVPeAY0lFJw7K8+KrbTAQ4mmNmpeTGz
pW9Wpc94TYcZ+Z6aqtrXbP+LYAc1tTPHnm9ygpYhRkvIW2MiyttCCGzhTma8+gp5zuCKvm9g8acF
1rybwyMRZ7jQvUBn2E4AlB6ORKy4LMu162n2ooNOzirMoHxbqTxtv9+vOuznskOHEvp8OWZ0Dly2
vKtI1Z2VHvGG9nPpf3m5X7n7pvdFPPZdO4anEnNJKmQQYnPYXQycS0XWeUE4oJCZdRV2qWM/Hkfd
g6E6j7bhDZRKhbH7eQSM2N2Hyav4lHlhWeABnjgBEQICCxYf/PK4KVWTdSU0CcDvtXA+3RsroexB
V4QWYFiBMTjU30Vf8JDoc+mvYHMtewCCedy3KaYr0Xr5SS9gdhqS/I7/1zkI+dCmJ6sGi2TPY8Wh
PqbHuaBlq6nVN30Wq8aUhrdMNkOI6jzqjOD8TRZypPBBHEPSTNLsVf/jmCBVjNGvpGvzosopFwS4
v3DmHxqIuiIeMbbuc2ilEVnGuZGStOVAujbKc+vIqL5QYHCsrK3LYMPM3iz34K6JFb2L8/HSD76O
ouZp4UF6fJRhYKNVRMpsZq5qGfZgODwehqdim3+2l++Qwe31HwvM1PfXmgDFWluPUPKuVBPp3CS9
ghvadgjCvG2wCu7UWnqaCxoQa6/G5BfMiVjerldKdfhx7f13QC006WdWwF/JafCa6coD59VM6cgn
smIf5gDlx318w6n7n16s9S86rYIQs8LvHeN2yR5XNUCdJWVxHFYqW7AsTeGVZa1DQ7G/ZetplP4V
dva9WkrKLaIU3L1xrve6T/5uY65aNZYuE6qaOVm3hAUn1vCgwg9cyGUGPo9tr8GRaXf4XAhA0Uvr
LTAqYOIw+6BJ+OaIobxD79n6OiuZY3tS2YWL4GJIrcz7h9tw9yr5OTMWjme8cSxZ93mLYjaSOINK
9Eeynuc3kPcAMQkZJb5h8+fl0c4s9xttBxHXDWRPyWMdR8cK4GC046ZIPYptqR5RLvcvRdDck0JY
2M/jZtOQ1UHVqUKAg4pJ/3UM11EY0fxZ56TWVfC5EWMS90vIuKZlcxMpoag9rSRAvhpjEsBr7qNe
izeCUDvuUga2B3OQuBmauRX5McdsiYkzp/6UdW427AK8kTG8GIFYynU3YS2U+jOFeE1wdJnqTNZ8
fvalGhaMi7l7SVWMDLOZ1Fc07CtB9zsfrlhEWXY6aP6X1da/QEs+GXWwrhdifwO08AQ7Wqg0HzYv
d76TnfYcuNyvnB4JwNoXduYWgnWNdtCajTAPtU88TX+wwc/0yFXSBWwXcgdj6ww4xpejt7QApjhR
s7fzUlt9oAL29kP3RZPHWq8IetgV4+z5war7Ur/dfkFF4rqFJywbDF3F0x02ArVERVO+6SPlrgQH
C5XI6cu0C2TTHFnYGfwZJIXTJ67C7zVW9zLGX/HTphVSMP9P9lx8bB4A5hBZi9gKiFpj3UQyMzkz
sYEYaYs8oW+uDZMUS6pEdahYk3T3LjVC+7+QanYg2GQPIWfY2EV+/7SboJf7I63jO4+F1WjjgHTZ
GsUQ9cTJbeiJt4MWhsPAvrVbNxsq0vxhFgnRHQTGuEYaa76+4S8CXMvtrT3XZBBQVOSZiDT2ZUTB
TH+3FjJIwRbalEZleQnV1RAWLLuoPcj4kPxEyM++FqZY6Oe9/eDE2sfBHgw/P3qsxNIRtXcojcVc
837eyGYqeGNKfx6SkiH3gQcGun3sV+ECvsN0GrU1fDoYvpNByjNkuCfALml3riwQuMymYtbWpaVE
BpBsXwTKuUWY1fCemvd+LzLNd5vmVG9eCECh0jnQs8wE59QZFjplIYxJX8+gqZ8afCPko9L0XjH+
49zL5w4wjzcOD9r27PnvmJx0uNcElRMUgPCPS1tVGmhOMdkI6hIMavNOkvGCtn4IswY4wf8PK3ua
2i3MCxuF74xqaQPDH6PQNKzjxTN0pU+wthXD3iluzL7ePu1CfNVbRb8EFsBVwN9PotPpqEv6MtlS
fvy38x/j3eBSHaV+n9A9IroNvXFGiyI6BHEOfk9BnLydaQZt3GGcOSYEutm9oIEDmBrZoI23Rzjt
FxRdcBTJEScXNdh6jKJfkxzefn+7rh4V/r1+mpreNLUHAJzhGH2Tifk7gIftYEe+qOCuVL18/Yy4
3lQkwbFyV1l6iKQIx3NI9KZ08A9Au4nE6kFjnN2kyaL/WNwToWDMRqAlNMnLfBtaOEXEMxZ94RZB
TU/earIRGIlG339n+Ui8t/fDDtBXuWCSoselby923zByV1oT7Ys2s4lDMozVdqzwxKFi2q3ONUMj
ps/BO09IwyLgbPXCkt47gjDX2rePnt8TuoDuaPcnR13JkRxdHk99erTTuEESwU8Mz5XljfkDqwE0
gvvRQyibvLJ1dpmo58Cx5a3QwQfka2PtJUMcCd4lId/NZZhuexcD53LBXVYM70M7A+F1EWSKtMqn
m8mF+yIJxtLHVPm/5s4OsUplHV1LK87Tve2ijXpPKL+mHF0AFpFLJzDHMsgi89tts6QiVHZ8tYoZ
fxe02rUI8eVxAKBWwCrXolsOt4orpF1VWZT807W/QD8zz8t/NEBLflaMA6K+FjGF8e29wexR7mNk
eXXdH/FMTCR/laT+riG4GoL/oNdWV8AQjC5bnlnKygbtKvIZP/P7OCSQZiMlSkbwAIBLdI5LtXkm
Kq0qtXhlJDm2HRuMIsSzyqS2ciJXPReWt63Zz8YGUeShyzFZDwnvwQQEVuWk0mpxWL9EP6oQ1o4D
tQoenWEqxTDOnUlWvfLB5jioB5q/k1xG2L5fjgvv9WTWYSyc0GMQp3HBEakfcHGrgffxr0YubA4l
WvGMobYpCN32XAAhDPacLmpNE971kpAxp1iAhShIfpOkAPIiV0fmBkEsNMpjp7GrHcTM37dr+iPr
Rh2URYKM6NRVenRyZQ0Z4eG1BR4ogw8G8BO2i8wPZRDNv/v7jvBgyRAMUpNs4PGtU/3zN1sFkln6
9nVuzcEXp8O5WnMmaxaQg/yc0KwPrcLpG++w2nZqojlTQ4gtSsPEt9BO1jQdWPpmgTdpBPX3WS2G
eFJAibV30vCW+ZEX1Fc5b5TNScT5z9nNxnV0ome0zUWQbBYZ2RpRwINGEGzDpF26dz2dD1UCyNXs
/q5VR7Y8zA+m/HyNk6r43gQs0d3MDGUsgu7AomH0tZWbUUWXx1ZZgVoljIPofvKYHSgZjA5bCEgk
HA3DyuYwYvlaHu92rNUDd5SNJlALgPGA9lLIBGdLzRNbEFA8lWHICr9svcAbOmM9P60xRtqBbYzQ
LWMjpFr4uZliMmFQXlbKZbQbLIRw2CliSDG5arNgUH8Zm4OtN1ikljlXLVL7nUyuLjp/7KNFdUoh
W7CLgVEy7v9X7fYDt7y9a8CpaA3TX82cf5VsgT4MkGSh7QgwACuVjFX8zudZ9Qbfjy5TVdAqdK7y
LWOR7fbtMkoo7QFCLFq+QO4t09PIr8SaZWIeeNcXDUOERTUAo0gAJeEXFrSav9ETFYAD/CJAoZWu
c/ZS/nl1Mi8Z3K7SrNYEiPNJyXTA9TW53TCrlG0Ab9AvYrMNugko076g2VHoIuhsGx37rpB85rab
OFMI1PoCsJO/44LXe4fv05gJmcPJBNnkU44A3eKdkH2U7l2j3bjf+YUKEOMiAunphEDcsXoqokEw
CeGqSh6tFmbXQuLtqX1f3RkmuXNsCovc/ispUpG/l+nDK/FjTBFveGwqyKzQ9T/vLiUwSGYrgurT
+nbkPSNNjVLzLhZi9+n/f4B/O9fbEWXq9DY6enR1MFNjoeJCDeiu7s69gnJV433PIH357Ltj2BHr
GpYLPKioU0D0ksl6fVxcWuzM5X5/4IwvwKV2RZJb9qqC7jdFg/NudB36/5wbZh6lzakVPMH5bt8E
7nKTK9PUeUADiTM+oTLsUordmgBcd7TMuJT79dMguAAS71RujRI4OlwsCXqY/xet/0vULeJunY3J
+s9DY2D2g7U+5Kl8/uOjc0z+9OeUznG/fukZrSm3WMDimJEusTEBJLG31jc5UpsaUxQn3jDE07Ie
D0hHaz1QdP87zyR8z3UMItFBVqzhQF0njHaLiN0rP03ByEu4pd1RqV40cEcArCXK2D/K7xPmf9Kw
gOsR0x0bxcixIDw7CfsVtpZJ8jVJxxJf1jtkI1KvUm30gNh1HdM+Mvb6pQPkW4u1+0GzqGk9FSNJ
BmmtCuzJP6z1szGyFDEjS72zLNdLoMDGt1rU47N2CIWP4CmZnHhKJ0IUbE1L56oNcmGq/qHH4OYz
qoaLvN/hYAGeVz8i8Z/t98xsCDkpTKtVCh0FvUW7flh3anU5iLP5EdujNsjDK5thO64qImeC1Gxy
GX1YzLtVLml2zUU3ZqQze/Z9hKtaiV4YgHJGjKCF3DOjb8p9rME4ywSmrIB62AWrq5tBWikAN3Kk
80ICB9Rf7Vnc7mX5rNqqLVMbJMFvoIB8i84svLA0jdd3JGu/WxaSS2bNu1Q99NTZ/ljC5LbkNFS9
OsALREM36GUSaHQnT1scD1jfsn7D7j19RyJYU0DshlqBd220UciVpFPPCjIFVxtcZV/gAA4gN9cW
VCu0OxxvKGWTD8wEWWCeQTbS8pp0/BLloMgurX5DfDMJdFhrISLB6lP8frU3MUsw1BO3uTc/dQni
zt0zXEyiViRphMAtyZwrfgukH7pMD02F6dvtl6MM+KUGtczX5/hucD9ULzOTMEecvnnErRsuzeef
lqitmGZlagpbVRjpNt3aEYap+9RBvzAfc5dN5BqFnFkc0rfoZOqvfP2AyGEw9mT/uYRkR9Y2lPDF
0EXLMGOc2eVnIzGAWZAdlX2a9mzG+muy5kjJ/pcgxPHyT3wr15MPOGrSE6wChJM9mCJ44wei+pO6
E1W/F3me8g7XofZT1Ccrc4JPlblSq7Ean8Sp8l823NhpA1B1PCl/4zgfd7GbnMQxgkaLNnNbIqF0
KszpVviMotZdDW/fFX7Ez+TgruEl5E2aYcyzE5aFtxmeXOwopMhdHPpRNhy3u7pzX8+aAUpHYPKZ
4vJkP9JkxJ375mAEzggpW71H+rk0IG24tgn8BWLB1I8H/EOwQI+dMUSNlm/jIegHFVO/n4SIzBqJ
NLtBfasm7ndwgb0Sfpxf/9AeJ8jDxvZr0UK3U+8CPVfipeJOTwmzmRG+GhkK/GewebNn7CDXLewA
jhqsfU84ywRBovqlf9ayMMEel0LPySD12tgeLuOMRb+TsBP7h6dFfvoHqgqVhYM5RhTTPAgUjdiR
WbuT4WcIuegw9SN0OUr18HSxIYlyWz+EBZtNle6iwfTETD+Rm7s6IWUr/BWRqalLQHyrUxNrxzmL
Y3XZBOSyoSlOZp0mrrzIyD1xcXlW53NWwFl9JHYI5DSpLz3WrbUQLGYqf9RVaNdv1auNODAThUmz
6RdJkDvOeNmD5V8tJVVcnDYwP8n5L6AJOSXmQ9ck6rIdU4/gF5985KVcLJwODVC1s+jrobatLijd
SS/uWhY03a0czcrF09M+xZW5IuOOwIaylXFFyca6U+Daz2B2XXQwmwLY1piSjmFLj0f4LRM6pH+g
zmjdXgmAVr6djeqG+vhwheTwQbkTCdumENTkdkXDTCOwwDHv/yDPxH08ZLuYCdSRDp01+CcHQ2re
OlBKUCK9z4i257tTeHs0Zk3WmZ7cTl5Nv7oHZhM/kMy6G6l7rH8ZjFMBefZ+XM2EQ2xGsnQ2tpaP
dqDHAKxKmhWMXml+9J0V7rJCpup2ZUaDSJqlfB+cSpwsAWmGEMsvw7g2iShb6UuCDItgdPSFaKB0
OWMLyA0Ei3Sfke3WnoE+4Yv65Klmek44xPMpQqqC+iH/9t7IOpyWmU1xBTRWJ1AIEk7liwtQ4arY
6zc0IoEEEnNR6JwJfvscj/ILklS8PrjQ3fJMvig2v96Wg7NP+aBdM50rVRln4jG3MdaZ7CwOtKEt
eZax2uPYSOgp8WAy/IKDR3jgpn5+2fFf/aQW+ZPTpMow6SRxnIT/gbwsExsWWoePU4+gwm2xOtrr
mkpK5BmiNEfYOMW9H0wBMQxPHV1kiybwL089gCAseuavExhLf3fXgodiwuNaU85V/MtbW8KZVyoW
yuygQSINiLG2HytpJb6+BEk8F6f3TnFjXMnrsPq8sfnr4+jpLjfuHEx3dJBr9gZg8lpUMX86fWjq
hdkovmDClLk8TMIFe4VEPRv+9CtPZ/Ac4yBXbgfhaTmUqzAmrY0RhWOOyan6Dh8c4EozzxnVnSAg
BctC98ZOP5xgvt1+1kI2M3hdk/uxNyw8LAz17Yim5M1BChu/sCKwIXLohHji78yBALvVq1QSjpTZ
e1qm0QjiyVIlRt+fK3JYMiayppWWXtkDJ76zLgGwzYPjNafOgQ1Z9Bp7G1i+yOE/aJULoiypPXwj
zbdqzLlwe5oVhgwwnC0sJcIjiW6dNmyhKJP42ZR6obtZAxQbnsvAOurGRCHm4QpDvixqPWMlM47s
4r7L/K5P6zvvjz9nnWiCbMnEPGg7XO6V0cjMb181WPKIS0EqOq5tS5PITEz+2jMbr3WAkNLHP6kf
yvq68FniDGYcF8orOe+8oec4xC3OAm9NgCisyiRaIAuICxGad0yEUw+jGa8M1e/xu1jEz8zjbXEa
qABgheVMtYUf7wxJOzTsi65ChUP1ItxgPL04iTIa+QpdGYkICX1OoKSUybgbSebSVqJN7Jw/hYD1
7a5qvUKwyvqrx/fvIgC0jSXLq3dmQkBJGHaRheUHUOPBX+33y4NwIinwfPeQsLPVwIqE38sJ/sir
vU9+GRxOhKpeaDHR04/GAj1OGqZDzG02/MIiYdr5RqeQAjHADH4MCqaTc+pNwRFU8/Pqms7xHZ9F
WMCtZLM2pszJTHrw0lpoS0VUYPklGuwhThUM+SM6rcE3h6EZWRU0DkJ6ysWG2f7ik4wRO8QFvmev
PJ+A0xKmgQJfjHK8I+C1iGC44nH8Yebr9P8xDubwM0VJ+TXabyXtEB24TetBoj+Bq/KBlKbPbRXS
gqHTEr9kvFqZYSoOngyGiGy1ECqUQA9cmTx0qDh+w7/aWK/vDkqvOyhMUvEyGGvFIYMjduliR/7O
XMDoff5EhTGdsFsFXVfm2pH6ByZMSQZCl3lPnBwe5kZ/HVyHOfyzMU89DwlraK4J2kHDh95v1hyt
zX+Qg4jK8iZ4+MP5uy8MKPqT2aqSl4OAJbCa8+k9CcOb0aN3lDlcXJPkmK+/nuuqCKsTLC1G8yQt
F92xzMJL22t3mH3siURdblHslgiZKpMWTYI1BOCQt2nSUzQl2X+O/5f9mhcgnuRX3ZZPYiS5CHz8
pg+vFWuucQGrqEQo4smLqRvIw/CTBcujCnOcDtDvNM66DBau2wdDjK4tJZh74QrL4m5PLfkdq1hl
+Y5SQO+gxar4W5iRwKcDU+uk2QBgENCTaL6l+Lg6cvjYC+WhllqK9ivopnuY5t5lxEl2AURzXyYd
SUJkd4hWoSYUHQmH00HE90XKjM19Pp7yRBwNPcBP0A30P5jj8PISGdFE4f3dfsq6F8UhyLUh8Snd
UZtdBud0eCgGGqYfWBucChrLCe/vb+TbNFtBflr3XA3pSWkDD4UATTo0It8oOt6qtquk63wsQ6gy
Ioch2qIvXWeWqiD0Zea/cepW+uvImzB2WilXFOZGt+ma7LDMfop6uuPC5T7Gv4Mjr+uWCUMRR45Z
zcRjfKsOLCXKV70iPZ2ZomVHZRrR2fw68jMpJlNueV2C/Ckh06PgWDzWB02b5UxF9+aA9/w+8fRP
0UrmmRxDscRljhD8b80dB+aHARui0hFZsLthYg8r3f6FT3P8ekwg/tQB5sqPfF78qRe9jCBs5rWX
QFL14og2uZqHqLFAeDDsj8G8tuX6n9P20+QGJWJ4x2z0G/Ug6rB2eEQVbuQKqrmK7UuGvaisa/N1
2KVzaEaiNziMCCW30kVHhJvh7ANuk6yFkr/yTir9aFdFcq5n6M8lasltXY1nlmxn7f2PMJu/9u5x
Iqu5T8goWlKK1fBslAatXEpD1XTVHNUwZbTQK/BUXDWrIQmz5DUu4FJKn7R2SlEguh2DfJNUPm7T
IeNMPe+EAyKiKzLXbUfsBPI3z2A3PpQRDxLLFLicNQou8ju3g3Ou9SCg5oY3BSj26UOD+a+lUSg6
5xYfcTmbhj7ytF6JAtKMUAtuhx15/2s5uqSMoUh/aFaLNwL7JOTcu//DV9LaKZC/wi6DSfypTjyq
GCaMBnmivVZVvQHMPIfmL4bphz4lJEIyDJhytuIM8TDetphLVctyhZB2pZesy0I8N4HgBrNa5Bud
zuTCducrIoVlUF7NYADRjmWiufsZzLyNrbSo2uQNobLMD0vFrkLQcntMjAXEZnhuMAAZtCgQ/l+N
Wnx29XIfT8iucgY8DyEg/X0DpaRFgGA9vAb+wpdQOHPY7N/6Hi4kws3w9F0oOUrgtGOkwKLa9P1E
CR1tFBXTslcX+XYJ/GxwAuA9DVOvcpKQBUuYUxZBc8+ZthUnV/9WG/94cFxcgaoqrvND/A18hF/A
N6OIrSUKCJoV+cRJGwdZhF78EbPSk8tRXfVoGcdpko0qky1AT3TifQtOG7jY4VReRIwrTEOgdYFT
bvXzdnndBnNEGC22An+UlwjcrWOmH8tbUfmXh+x7cmR17SWmJnMXWKHdrzPHcKok9HDnLSiRMwMB
NMCkSGpKiOoKGJ8WP7G8TmbmuuK2TRdZ0qma5VdKQCHvQcvTEeQi6BTxCBU6XTBVbTyRjPHf3UP/
c/EjYufTV+G4iOuyiLcu0BVV65FD6/V/CpAwba4WmL0r3yBS6FjgFWPR137QRJ+FmTH/3qeMtcg1
RrUBqIvOhFt1wK4QxTHN4kmeVlAWtEd1XqbCgfzCsa7mDboJalhg0poKm037qEl26H9D1onlCjSs
BMGCANWWKgf6+mmVPeYeHAi4qCUF9UHvYBEGjLU5eJwmfF9BM8Q3QX0UgZyyEVSrhoDb58cbnoU2
9c7E+lcbMmCsN2ehL/DhQYovaAq1MdGRUR2ra5GgDcqkcDJYRUzv4MIKgJqq0bhYP4ZyGcEMtuyN
HfHRj1b6YPsjinufEtRi8ZnKmhNFrtJQiUX4Ix2qo+PVg663bh/3jxb8Vbua4f1rvIfY7gthj9/l
143yZCSl5/iYvwRYXVapwlY9Y2LlxSVtzP8BVpNyms6RPgC9DP7ZgQiVnHjhm2uSZ3HjslDvC4NG
MMHLX12l2mBq5lFAKrAXq24FxYMu2nM8cpvvWfIlL6tIiCaTvJgqiNhxIK64KrHRq3L+9wJELSEp
0nYjzHMCRieTXOt9ohYUMpzkGZqdVUcvXYiC5DH+0eJmnF+mRTiFUw2ri32lb2x1HHyyE13o0pam
YU1Ym41y2mcncGQkihgk3EuTfuANDOfZcE98V2+fsFkGL3AsFi6V76SlEUg9UQ5UAUefTJEi9PvZ
wuLZ1L3UY/ISGIYiE3YEB2yrQXp7leG1BouoHl8sr8paAhxTCq3/hcEzLkykyVNFxtT4c2XyRx0t
cE0LHkHQHFwhr5onPtpvPkGTmp/WIToUZCpM9tT3SZm31xKD14wDZwR+1NtU+lxMGZr/yZ7NaT9O
1CWVzVBuS/zH8QwsMmWdpW5psA98mzQ7kxqTzRJNeTz0YhgIkFHcwYGkXy9yLhOLgy4G+KoTkfh8
4ZqMUB+KzbpWF15gt6O6MSrZdMT52srib9gQHLLMRRM+kwYOep4mhbkvD+A63HDA9s9ksWjnA6op
GRqFiF0LkEjM2TyQkKC7lItLtpCcNZVKft6n0xdEi5xPazx+/VOTzTN1jSG23uTmfcmyzGkjDvwX
AKIklu66g76ULX3VjPDyIZNKUiAzTX2WabTzquqLTMFakgqNYUsTmEskscs53rAiHL442sD8TFA1
zTnpBDrCntbaZsd84KM5Mtf6/swpLsBqWyKTVvz8qPIYr0C375KLntM3ZMQGSCxMElQ6HbOTlVjN
PyaGCPZzT0rJcXONeTS3AfWYGVqJ7EndAG52AwfR7XIPkVw9gdvNOoiq+zXNC7vrJ8sQzymttK6h
iNrJgyVOUmRQof2zQIhjMalcqZePo/yXxbQt72YggdYspILRf1Sel01cxk3XBEe2v5RPWCgNRcg3
T/gwwpRGsYhbe1QpvTHLbVY+WwiI8W3CyWNFZOu0AWYJY+t9236vyUzy2hbua/odV0IzK6as5g3o
vmjlCLKfdQ/RVBEgEjuFP4SX0VVer0usyMOE+LvrhFH9S1HrbiwvKaQR/u7uRKUOI8rJC1PueCu5
WNTmASV+RVeBiFHD90yzf9JVCbHf2VlXffqo4XzcCTDvS05rEbqPgQHnDxuH8PaeS7PigbW7U9z/
bdANjsKoZwjwYkC6gOX41vDQWJREiX/cI0inomwaABZWzT5Xq35akxaX3WbWeOMVgz9S8kiJaX0p
0nwtBPkOTARON5zhYuMW+UqRbOKhlW0vnrmhwbEZjQcwKadPsYc+cahsR4kB4Jvxt/HAx7lrZ38X
D70DBq/TFmqeRqhEtLQ6qAdRBg3dfUg8g8Wh9hUKwUmQRMk/Lt8WQKlvCPfGs0Bk4EHjFJTDRm/+
nCQfR3JgxBEMeP3w1QHgnAwqhogBFl1TMpm28t1VRpRw7kbnDZ7J1U0t3vKDpefXCrbTd6HDba42
LWCNEaGhaGdxhkDYXwUH3gtnIJpxEiTKZEkbAsbXSVdKrf1ESwCCxxmCcGZvhRySeOdmyfjj3vLt
7ZJtCZyuJ+scMzRXNiglaY9UoGTC3YjixosJRE0b9Xn3KgREBvCzLjFZEPQiEIU/8TXl7f2RafBP
0jSn9Ypuou0GoHXRmBn9OGGScaypYN3GVBWCbNO+yNmSxTALL3o2teWjxalu+XOIkjPGylxuT2Kk
O0CHeLQ0J5u19FjSdUS9thYFYMVPItAems4jjUcWvvbbg4VHbqA5SrA4EML8IaUlL03l7WzsDvb8
Ic9MfQPnZHOmNy0V2Ww0myvmOUSCLwff2DiD3Pwz51EW3FANjSvvFMK5jxjOFX0xMGk46PdNWl9X
JZC0e/Ejbfvpqk12R5DXphOEVixmviEyc9Su5ODtaTneHgDkdcpXa6Q4gsVW/24U81+CukdRwHQ1
ITunzPoZnj1Un0rsTC7caMpK3GEhqu2/Lnsl5cFeyC0UKzmDk5EytQkyirtZIXKYmeAINzDDldxo
lX089R/wDZ22fxDad0YIevPZjzfHZuPgOeaJjlzeVhAkzwCkluPhYaUuu85RfEbGwzGX+HZfZnkU
57oPHTBitRdC650g8wfOqplSHl/Rf8vhEJ3F0fJ4CbGMPP3CdjzfqzfgCrSamtlE4F3m2ZtScqmq
MCrZscvIcvZxiWlb4R1eFyJe5823qUOJ9cvxS1YBNyW+KuYABo4q/O9+DkWvRFi16/SQi4gl+dGF
6nN2vlspWBE3IA57hfkqyRnrMeFfbo7FXoZeyr7FHSbOnxFLZ88geSZkrVFU6BKXE6muqTJ5Mdvi
P35USsf/+4IOtWIOyxlKuibpE8VJ/PLIwsOLh2WTY8OLTzIJJquWA1rLD3jDUIJJW40XoFy7rII+
3B4Nxp4rRKuyYdx09j8BIU98Q9K1ycXfVfgDSGaBJn9nrlo6LCytMmyv8JLiLujqgQzsnbmZLT3Z
WqSJfU1PwXv38BoAbeQviifXvL/Z0CH90rAhsUL6Xfa8HMaMW3AcOzDDGktsv1xyfjM4P38eXoF3
/heka3XUW1+etQWv4eIZiEyc8QKx3Ztp0PokJNxsqlqGOX08JwskGZEoQlul/JH2d9qvu14ISg0W
QctPohKVcolqIjdxi0ZKHWKL69qzm0UqP3ewSNyyX/m5JyKDU3aDqnx0nGmMQqU3ugegx7lOESWt
QOy0hiC/ek11mKXPcgv+Qazr9a9yJ1pcMbev7q7y+4/q1DOBYqyIHndrwML3IGlilkakay0EDGe0
/HMMYXVi/qicrf7Li7wXyMa/JQDsr+1ge5BnFkdHfOVH+ktTmpLLrpm8O6zwVGmRM2718fLUM2s1
9XFEkaSj2DRIudcpPA5Rcl0d4QRVjc3eX32vqqWpItH3vpwWUlPsDcJxp5lR8lFs+9KO3hfOdZ2h
qIKPAt/4hVDKWQvz3kVHaVWLmupWcqFCegVJJxH/oAyOm7dQoU/byzAIMTIGWhgb5hh1TxxVsgBb
y+KYa3SyVan0iJFkkhSYhBtlGIqMdYnwlxlFeoD55GL8krrFVNdQpNnfLzWXY2O/djv3ySIFLtfi
4rU38mcnMVals66WOfeukishwR+6AU3JKhsKtJPTF1X5oIXeSYVQ1C+U2I7l4fUZSgTkWeyLW+xU
Ftqk/Bp72CyciwPu0bX1WzHNIV0FER8iOveYuLCVOgoRxSiuEPaIqRDFRsZQ06Sr+bY/RU4YePob
E8NpjHA4/n18Gi+rjT0oAeO+JB7U888mkpiSL9revBVs6KRW1QNjZfeBx0941uGL94Y4ItbXwwPV
JgBbaXIyCgMwMl8qNCfk7Z+enDrffX6C+umXKeF/DY0PVvQP1ZtovMIe7ljRuzrgsiYX+DLspvsg
buctkc9yIPmAFOX3vjJk5N1kgbRxkzBIrmJto6Z0X7V44fWuTwg/tcxPSeT5gvF5ABU9Bhh665Ln
Bsoeahrknobucgo/KBo7Bb+Vp0Fes74crmwHv3ZSqQYCofx+PcmhmQo59DzCQfJwb38bTvAc1afj
0lxtYaVb8fCx/K+5r10fIZWXMHhYJrIPRKNgpI1psDyJU5DSntbeYcKKIOs5uV0DlK0AejnRj1VR
rOAybV73ias9Ht4Oqostlz7SuuVezpxrbxD63t+X18X2SWTOCtY7uXlEP2Z08ME1uS78LHOc9oFO
9c1hnCnjegXqnJCupbUMpjSs6EKAkJuBuC8YVijrQGFmD4Es2pi+M0uW3WWFO1aIybafWz5FpO6P
E18+ekD7KEtFcCacrj0fi1fohsIoCvNV8r2EQlRUSRdJuO+c+PEF2ue0ojo7PJp8VV9IFz8zffi1
BG+apVpI5ycQMaAEO0PD3INJryqwLuIwgz6Jtt3nXKxDprlkhXtGB5NRPqwL/9QO/orEpmTvftxi
rHzx6GEesbaKeCs7OQUFOqVQEOHVYss7OPcFCpy3qJb7mKqiJiigXoQhchsqeuGi1z+0zvoiA+Rj
t/vCU7x33l98JWPXZE7H4bwB1bxh4rx5XFr8zGrkWHgzhVVTVCCyEggK27u0nDSvNRYcQcaTIuuS
MFuUXYfflF2DngAhOsLhBxWfSIZo8RnRm7GlJdgswNQyKi9I0zUs5dfanI2fdfZyJB6J0ndlvHHi
SecqDVaso/ZMJSgtAT7FHm29gz0XXLj6HEf2Tzgz9CqwRsTeL7olMQ0Au1Pv514OH3WRc/ClReog
0i+iSSwXlK0VCcA6nTcGHtzjYxJiVw/dlfjgb42vhlyf+8/4h2kyWkZFk01v4TRGiqlE2ewpzB1z
Kq84oI9GPccG/RiWMQXAO1xFlrhgzOntQDQ+sdNbMB2IM4cLyntA9GL9+ZzOhODPzOYvw9PrgBib
nlGbWKM86ApYqRmlZnQFPF+SxKCP7hQylBUN86GeJRL444tqAmg8cfPOxb4+hn1IMQtT9AHE3oaz
zEBBCG8uY+hX4b5v+iFtZENQ1e/LEkCs0VPnIybWdlC2ond64dlZyuHtlO+PbMd1O/82NUAYx8Jt
OXaCLVrONRTHjk+SSzRgRO04pmtTatPa7MojbyW9d/xkBwnVpi8c1tCJ2DABoVFSeL0slOS6OSuY
3HguOD9/o1MHywsoPer4jmAlY2d0TSGkgXRIjLxvxlf2lJ1m1zZGzwkDCSKsRO3OaWJmvs8r5pRx
NA/KjWKFJI4DpRa0CmknvtqGx8YrJ5m9wC+E60k2GGcDSlsDkF86mRZFkkha1CJL5lx1nDIAovPT
xjQ6yJqiZRjuBRiLuLc5/SsjzZHvlKtasC5qwIq3bWihbc8h9rkJ9p0nRDUPxRlpRbwtevr3uNBM
s3gdlcCVf/w0oCJgjxhQ9AJpSAQZdAoRUSlgMnQgrLvkMah4yM0uF4qsWEa07fkjWaIAFLMtpJBK
nhmdqp+AbAMB3apSUUP0c/nr7Iv23f1uxQ97rVfddWSf7mseJnXMiVOOS13/PXoDeNCGo9XcywIe
EWvn8DNeVD+/vZ/9BdVtdga2d5YI7RrqqCtUVuAH+2/bMfp+j57DV2hcVA0UBBcI/oDHXa6SV+nd
OYMznkJi3Quz/RWzzuoV/7sbfv9T2MBA9h2Imzx6ZB3ZZG88/N9n+m2BCJuRcqbq+8msWhuZPAfD
spYhEE47gldEaPZsV0jE7v5o4Tzs3P1CgnPkJJF+GYhrEn7d+14sPCEeaGMWmCQFO+AKyv91Z4nX
JA8plVUpI1rIzgg48cyCeez5BOu1H7LY4UqXLZJU/GhgYLv1S2IXQrldDIkORvLlTzmpgwQnRDjP
/TWu3DCj+c4cMvUV0qK5TpROUuVVvpzKkZQW2mG6WCveK9t9GtV0pA7iKwSsIcz/PWyRoYDQnM79
yty9xwp6RFu4JSdaNrMgxUirPHkpPrGUK4OSsg8hBY3VQz1z8eVmilcoSJT/695KghvzAuUln3KN
+ebtAxMfMTWAXlj7JrIlZDPB8dYclqFNNHIwmtNFmzkZUPhkYiAKnw+Ksu6QiPU9d76+roNkEKc7
l+lDz5Hi6H904uJ6lY5Q5vHXbFL7gExxyA2r7c8QRRTYC25D9/boOUOSg/uncgoXUw8UeQLs7cvl
UOvVA1F9j5zLj5av5nLkQmD2hP4hQIGfOa8KDjf+ZvDQJEiO7g+4aGUZgprj/VqvloTRW3cOgFAL
qErEm77jYwFNSv6w1sCVjEY0RRrhe5GAq0wK6qm6cpAq1hX6mTxz80SPjzSCNIrGRDvXpIF25rRW
VDK8Zrz/5LlFvbckmDSKjA13lvYfZa0XvfElAZ40JdNl0XtS6oMOXKb0w46X041WfqKxPrE+GGY9
Gdu++W+rqNOT7WgcFC+jykqPHbW3PjiCvdyWAtE4sc9O2bV41GQgzAjgOnQSou+6jnLZYSlnSYpv
3b68o4JNC3aWbsnbf19FbJ5aGgYyG7WZ4P5uTyDmFRmaDPCbdTsVJ1LqLZW4Srg2wKUrv8xLcOe+
cXemKdePaCLxlmF15Iap2z1fEeaRzy5rsNMgzv4SCaPbXK34IHe4bqdxItXA4PrgVyMztlCXuqo/
Qk0nCwmVaGsbOtDGbTwXLG92oqz3E35B/XXkG9F872AgeQdjhEyPmx4e+h2P2NokiDa01TfFlnPQ
P1ljenxW38BGt27A6biEH4+xUgzzdd6LMYkCSvoO4NQ6ThzXt1iJb5GismlEKC2Is30MrI26wcXR
JtqqWMMl0N52uvWNbjn+XDBTBsOtxNl3gzNuyhBB/uGHqdsuju5+m0EEwUfFduKPLBejZKwFFJvV
zIhA1RKhPHimxiOpok5zyp5iGUvAAt9fOG5fl1H8HBC6t5Hn69QSMn05Zte8RBDBOMWaqd0s1G0x
mMZZA/+/XtNwro2zb9o+cznh7KxYLnQOol8LpW+ddlVSwKtPprHKu24NduX5CTW7Cv7sANoDEZVw
Xvyyca9ncwCh3weYM9Avx5PV5Mdrs1seokBqSmmS1GQVhd7S6B5GxHAg688uKJJzYhF0A/PrXF8f
IoFdqPYgkGJfGAli7mVF3O9aeMM3VYvKM+fEHV2qCq4yXWE+TovH0EHvVfyTiesEEsZI18Js28Yr
9r6ltyDhrs7dcPuKQnASQv79pVkStnmlRvhdRogBMP1TZETeo1blpyCBV9Gw5OmjycfMJxReezzv
Cut9mKqs4O3mR/OWXm7IYFz5GZsFJxExm1mtJEHqmH1DhBAUB8UMKpE1ZvWE/9cEFOB2a1IuScsB
Io1LUJuAhoq+Zq3Y78t7ygO3ZjqCjfjp+vRm5bHkKtbkv479/88Ovl/BkHqVqbjzrPk8LPFKhCSa
nkM2JLO1n8yhZDISQX0OCtMdItkpSAPd85FHfz2559KUyueITlrLvkTENK7f9WL1uKYFXucTvtN5
daQRFAdqXmbESvH8w8kUwZvA3jsOPP20MbInENvoPs7URDfEJo5pCN8HMc6HBuCf4cO2lMdvKOrg
Oee699UjlO1srfGYn+V1Xjx7R0gJoZ+Mz3pTSgD5NVYcjfj4EQNUusTpTv5k5Fl6qiMauAGLk2ka
m7qm/aZX7MwjqW2gPLf7QyxPLbBUsYHwtIexzGs3tJwV7S21LDH7sO2noLCFrXigZmAkQsTg9/rl
ZsIAqNIcpNsc5z4MREp+DAkHsrLURwz7NsSbG9R0paVLOgPy/vxSASmfH8+Btj7EdbtrgruiizEN
a68trPjvWo8jN/kJTCyo9kqq8Cn72qH1bdMrzTcsN0fvZD0+pdemvSMUZ80MDPJ9RfzRxzJNFMIU
KxghZV9Zz/JSxYlJn5ubqMYg/lP/glXIozsqCOL1WrYK79uHQdzKsL8AhM9y1I67yTqP+D/MXujk
iRPMbPfQV2U4CAal9LxeBe+/TUuT/v5VbSL/u3JuZ8zluCj+tRfWsUYGePCSxzdoSByC1AntD3wN
GzE8jdd9RBujyv1R4iFrIzce8s2vUmWkIpfnMP6gIXk9nM9nocnAm2SBBEb3zVDY5kWe7mYGMRCm
ojWVIHeMy2tXUFlfR5DW1vK72CYRGgTGQBgXRuQq59gpCiTpA+a9h0HJO7llcuqGRyFeyovJnAGq
OhyRbo5fJkLX6tvWn211PwBqBQIk/tX3G1jt4ImbtU5w8HJMbINe57nSrzBTzK47NEnh4BzEZerU
i+kay7o2HvcvSi7nks6cFYbATCjLdmuFQJisIEqOvQN90hPZfNQoyx8SSGGeVPpxlz1imTlHL83e
MBcSHribK7lx1myJAMP4yh+x80cSb1vIRbHEAqSFLsswbZ1SNd7OH5WNAyccUSXJVAnlQUOEOvPC
D4tmCWykHqK43xA3Eb+jFzhTopumgeMHsy2WV7dz1Ec52zOaI4ojCutPg+Scc7BDKi1SXZtEeRFZ
+pqeqSSfANP2Ph8bivC7asG0K2W14Ma69ve0QVi3eYYT3tH8SjGJIyaj/wfWuH7oUMJUW8hn/Tl0
weODPYEm3SZtWq6AgCObDxNyZjY0U7H4QTPRy8hKPgenESKfZJIiC1qH7SU2lWzT6IZfKHVU2yYI
J5a4w6ugQkCbqktzQh80sYyYlkTvPDGyCEVVqcRWhlDLQFMOxLp9J/KsrXXnroVw/ZxV7Mnmpwau
6ui4NTt5QRCnNfoZKK7f6z49cGE0FYjA4F1ni4rOyC5ZdITFQE+V05fQi2KcdjeimgomFFERsKhA
rNBnh3fgl3237P9dSy3BzAt5Qk47YJqxErjz7MZ7ZMYqVNvW7iue56Q7/xBLJY6/Mw9exta5IZWP
tUOcSyyND1ay26L84JSVO8+O2pyKlRT0GHsE4eQJEt/bD8xkVhMu9P3Cqpl8ooA1HZG49L/BHGXc
UV3AkZUowExNpPcRrX4PmpcsqCP+hXzb5C1zgbhskz+n9jTw4e9Mnevq8GXFzMzovGtT/oBtnWzk
pMsOhNeUE6pQg6JekcGbQTYFI/Zqjdjtr6Kn+zSoffP+6kGJoAwIoK/iaUvjNBvF7euL16V/nDS7
REZ0x+rjC/sTw5U5BXYDCB/KVp7t5zTflBUA8bGFHp5wvvAUAB58Ppd5d1dFhaZ3se1OHfFOr038
+HioAejlE/KcuiPz9bh6eXYCG0G+lBm3oz8BrQad3hisfj5QnVZnTzHUu1nC9CMpn8KMu+YJfSwv
VS2dKzHscgc+G82Og7sDmYDpGLFKAKRBlAg9JA6IpaqBiIMcY0ke5/LCoyEAdLQE2NHswtPIOfon
3xn+UO+EgaMYpopcSRU/O9Rpct6SVQN4c6Qvshh+tG7JALVncr31/LnbsP9hqGvjNk6r4qcj0141
D8mrgdVEas6dmfBNbpiYW1UFFynzczkl8/UvalckBwrEjvP/kHjSTmOLT62eGtH1K4GU5PTrpZ66
NKl5Zj10RtWYoLlDAifg6RlWbcExysrTgiUjKKV49VQ/ww62AVCXBkmeMQG2ipnGHVFi6HLNBnV3
qlFD9Rnl8tC5GD6CFINGSj14XnLXRMxtaM33DQjBS+4lRyQ29N3c5N/CXdgLtNq+MPCe+jXWCtoW
kXAFV3t1J/pbxC8b1mlSfMOt6RVn6IGgXk0cSLkIH7vBUZN+lbTlrWI3lM8E558UYNunjBZqTzOI
FSsyD2tlKhG8tUsC35RR/qLIvBeDqB9mULxRUcYaUmeZmX5gmWA43AMH7ZebaSzoGcVDPS4xuLxN
TP5QHYDP83Hqhvsj2iDlwRGT6pFWjj6MXU58TMngHJUjpRpUXh6vQPJq6U9ZdN165LZN4YCn9D9C
I1x8ROcWb1m+2CtE44GH/w+fm4ggm+5rEE9MQs5fPF4vJQ2lO6RhvTER4xDQFrNrrrIrXN6Ld4eS
OIyQ7hfOWagtjHcrSY51NXYPU/5cxbxmFmD+0XQzUBeG/+fcQQyTsonS0igpYway5N1VLiaboqou
oXdat8eqWsCkccCmyX62ezJxbsKZLvnt3NK8jYJZ25uCgAVoAgg8C0ySazrKeW1mm2WTZWpxKl7j
O26nOtTnuTrffFfHwUhaowX09ePDMhPuFcVxO/PcroLxIivM0ua2/Lr5COYJXIUI0rqMYCMGyAYs
TFOUfVYsF/4dz1CI1g3s8/mAHtK/QPmH+Fogv5wXkontFbou/M/ljEXU/Z720Gbn+N2py3AVD8RG
VPZDlGS5OJF0a1qimHa/TFS10t1LxaRyq0fSQ89A0mT8kLPYBQWbHof15jJOq9NcHWRHtHrM0NZC
fDoeIIGy22mXgneepPvRxZRv7CUpzmggd8zQV5S0Ys3mcNQwGXapnsFdbEHublmZamunZmCikggx
8R0IAbp/Uyn2CwXy+gFnoEcCw54BAPs3dOJSZVx1rR29Vam9q8bP7PpsnSTNkSuCrZHUKlljio9R
lqH5ZG7L+trygCElceT+4FlajHvMQGcxUgL+GpZYyK2rRHXNSqrUEYi5qAbx8FoWOlFm/6AExlk9
GqVsWUo+/gV0zozE0DrVYybOkQ7lIzbvaXo5V7teUWSzZx11R6layT8kXNDZDCKo7HUeKDn4Isv1
5xKlNyTmfU71oLvR1AJY9xxSe07qhdku5fFyZVGhPjG56khDcOLqxv6lpZkppVhN+hgYAvqP+SNM
67M1PGhJpgImwiM3Nl5m0ax8s2UXQ0jY60lqvkWkMVlksjFVSWaJIMIuDKxOgd3zwTAbz9gR+9eX
7Nw/cqHMb1xCGV7l3qvRgCmNLr/NdwqvCkwccDX1W0iIE/c4T86yj2nDT3cOZ/9F2DZL32jLhYHW
GvUlZoNCzdcJ5cDorlfWifoLDfOAAyC792Oa32sd/RkRYR62puufiA6yRq/wcVIOGW1OkCwqUqNU
Fhnn9l5IDcaL2dYyfuGh3mfGZMmtlAI1yZR9i7Ige74sG3YClRpoiobAhJr+gnU/T3sjWmgK5WnH
dl+oZIcIH2xXRXjm20Qq0e9EH7uopsyLUWokhjIE5qoHNVbfIGzDLihFiCwm8Knd0u/UMG7HWwK2
rv1z7dpK1Iie/o5ddIekr1hPRKMnaAKsFdSmOuxHLzmdpu/VJdyqt4g7gY3i8mCUHJYY1x+XF5oJ
7BZGjeLkpAOtHPWqBhvk+u3J5vZ59fLv7Hr2m6JdHvw/7s1GgYjpVhhqwedkpIknpi7Ke6eWsTku
GtBj9cUukPYiLA6K+brJgHT3xyLzqOcfWNSQqmrhboNDZQSf7vj+4k6E+5MzmE/BeBhcqlfcbbGa
x27sdiT/1gBvam6ocjG4GBc/3WyHa+RdxGsTt7Tzwr4p1xwwYFLkpwoEss6wvReclU+2ZXD8BSfa
DUZpfXyFDgkMQeSwoRFlCOQuIH/nhBmsWyWRiKy/oFTOLHHxK0jWtC4qs++ZMkj9HLflDb3v8nk5
MtwPvAlXRGhzL8Vk+gpxl9EbsG65VELm4b3O0/oKpIV7XQapxwGIyUQ4c5OeRPuSCdCjvlAxnE23
911m3hSdGI6DlXArK4O7o1INuA0/hYrHzhUfZGsvRX4L8cJdlBz+DgZMltjpEM6XoLZWRGYaH8se
UsEUapeAk1t312pb6qMnTIzPPVtmv8qeMRHpfkkEmopbvSObpkH5BI1KSmWwGXhpeYZ4GGhDjBVA
LsFqVe9mzmKEydRdhLqh4LGA7LKW7dKN44zQ2I7cEUtPnZNs/q+pFfnguua54yoA0TKCyKG72DR4
MFqn4TJXOCVHiPhu1iUraPlgq/BEgeIIKmswTAVmAq3oS9Wg/HJht+RwkAtxWdnU37iV+VxvVm2h
aQWgsFydRsgKCtsVvCAc/BVjU9paqvy9boOPD1j7gKPWiSIf+NSvvKFXAmj6pkH+fMfKOtC5M7gV
cgHh4zMClFK+i+uES9m+d9ccZW9/L3gq7/w6pJCub26BJIKr6GlKpoCDHJ1+8EWxODUtsZZjCAQS
l8GjrPAcXs/HfqWfvQ3zd7UVQyTiR8fuaCpZ4wsIbzbeJ9mpKJX9SQiB9IJNlHY/SVw4KaWS7sdr
JqmfQyBYFQWRp/GCZqkp7wwIgr6g4mX1aUQKg1OhcXZre0MpYPvUWuw1vEq1hn9ePkdp5ihAnFx7
guex6T+of38z/UN2C7RewMDSnz6zSffFysvdr3BUB4HVjw2Dd86tOs2Ez3PvCO0Pcg9g1G2v9HQC
C6fI4KEB71EaGrZtAXIf/DAsmpPIntJfba4J3bW9SXR2uuyw1L/6ys/l92+jkdJMZQ1ElAz1dmZ3
sA4MxnhPXsQfZFDYg94eQDT6LVlVeZDvuiV+DQoyDZtYpG2IIUb70NhJmswq2P+7f6c4UFfwxzSN
GQMexNxkoMxROHX5AYSbVsj0Uwew4uHjS3SBnXR5aoLHheqn20EQnrBI6B1+ldUSOvR0pQ4HUmNg
G4gZPGIgtiluqdqtwU+7ojCV9GRpzhXjMhntLM16xS0yQJvif2Xx5Ck+pMgVRUHnyq7fIcL6VBlX
AIqCOhQXytdV2DYlo6lmjWT1zrFHyX+a2ZBbiPyou4EMrGrkfTwTM9aIp/MOy35+4UEd4c0HHIhg
wmfUn1ZoEOwi5uzqlcgWVd56tOwo95RErpdTJWkp3Ka1APyfeWA+Omi3xH63UPB0BF4iMWMD7ulS
fK6t5CpV36D1NlJ9T7DVN0XMkgTbyCn5m8uOktvWtoxORE9jyBDvG37S6ted3kncVB5X4Y2pm7Pa
AbtJdyr9EmfR6RSTEoHt/A3oNDiyihO+NwNq7BToAkcnaDG9owLSn4jBkp16ZJ/ztGEyoO9Uc2sb
gUA9QgMYEQsN858e0KU4KEFdwnmNqCqzyZBBH+V9tmF9hT/JjYm4z0Aujb+dAVjRHhVUIc38WMnz
je4kZRNzYckK+rgtSA8mRDH4NI81HZBk9W7Lh93Yby550NbM2QYoqqTy/WzwPoKXLF7Ri9Bdj8lV
c2+jjSfhcL+QiLRJZoBSMEOLszgb8buyAE+BRqQMgOhje+Vx9Aiz4V2yHWj2o7ta1dXLraGM1uJY
f5Mc8lstNYC72aL/K/J5gK7yPXS/neCaGe2ucJKm4JN+ryoZTIvVu2CA9mfxLeVaXuzBAy2BaYY2
/nT+6Q76cyvqBYJK7+H1Affhc5q7cuaRcI0GTVGtdbZ2YdEUB2mi69XGycCqx2l4FTL+hnu11jKV
mmVTsA35Cb8138dWFQGUKlsAEyh2GOzDAk9higfrWBHW/hRXiF+9HU7+5V8BN8/IAPG+BnNwGg42
po/cqUVURlLOdVwufR3Ifcp875uq7tqG+gtKX6xAjlXyVELDXW17k1Hd5jUUV0jYO4DesNpAh1R5
0m3EVgsoGr6mhoxqPYzQnUggq4fKXQXZ7ZLRQypSvnUHKSQjVMqB7T8LBM0kLLgNeZ+wYw7QI7Zy
9SiEJKjaFLBurFZR5bA5IGgVCmCq6rDKtHKWhAT7CSkK+YPlFUqVkpc3fNg0xS+b4fd4M7uQFptu
AYy27NUlg18H7rN/s6AlIt14jBemwKfCmbTTfM2Dc4LHeb8xawA2LhpaZ/LSMyTV5UsrY3Tt6Zre
VyFnHQPMi751XH16q7q2xk5QSY9xk9YuD/3+5uJLvPJZSJy0FOmFHJrSnb0JtsZlMRB7A4yKg3s0
L2pV9ab4jYNw10HjGqePBHBaZ6klYtLl5kv7T+dq2E+fk2YO2GX4stOqUouXwj8r2FVgcBsAH2Is
JrtsJpKZ6qN+9XMQWbX1z5oEBJE2IOXbPcLLC1rIuJGbMFf6GhpuUx5Nd6/j9NZOXX57bjSfwk5y
toyj9WygsFQIXpZV9ITCyBdC6A2J69liod2QTmW11UdvyxZOBx7xpI2xo7Lc2BKw/D5tqQ/ZkfWp
CngpsdMj6lr3TU0p8nguQp8VcYUbRjrgpRK+4DvxjwsvfapOhX7s7W8stt6q7rOfMmPFRXSUegM9
0eysHlq9JTGDCbHgiTwX7ZzOMEhfteDTxfOgCBtz52q2vo9Zpu2xOus6SqU7Cabsy46vyg1bZJoh
nFFrDu2j6ICvzPXjS5Z5S/8EPrj/IkeOKKXRx8NV/s+T11uvUf/j/lTuydNqWRLUAof31ZbY2ivA
cptTFAAaxFYJOSGepXE06WlaqzO/9sokdLj7bvOryIJfMQce2RKSmFBP6+Fe+30usA4bWPkkmJv5
xD47O7AYawZNpSPSDbpaG9DZ/16n+3wl7TMDLTdoqTdZzawer+FoFwCp8oxjcyCjQ8KIxr7gjDpd
e9ExN1i7se2xTsZGOU0+9/cnz7r9bmdc0dL93aXANU6UeJjN4MZK2nXEzIcst4id9JbCFqwm9K6d
eR4VJ7I2scXYWwgKFaMWhSQGAFma3nCt73BFzcqYTvNCmx1+81zFPu4MUjuFG1G/NTjITAGDGHQY
UlczAhifqUf72L1syJMqPCPW4ih8bzEUe99ksV8Xe4tdUpDV+4rqgDGXEleQDdQyQTEAD4le8EJj
PIHTJk8SgqjYLthZn55hTGamFPnNgxPhDHcFW9Kltsn+s3jkYennF0RxqIt7XHM82A2Eh18Wz8Jh
o6oDbfvT1mrS7aH1THBL+SBJsttQRBRrXi6QnhWmu2NwXDkSO7mUtz9+9dMHXBAscgjI2tZgtE8G
3paU+xplTJrl84upL/uXUepMaUicVLPR2IeUaOfkO+MmnGttc2xeojUpeNc/vCkdnWjsM2Fsmsu/
NAzxh4AFr8uWrcs497vXefHDqS6Cix3o5AqLNsXXwXS/U69lPrpX+nXymnp+pKb7o83VxQPvzrxM
JdarQk99dHV3ADrLa384oKpmYtLC0VUEautOWOJ94DHQGBfUDFxwuUu/MWnKGo2CegRDqHEp4uDv
iAEdVIuto6kmXJn2VXmix7fVJabpEU7/5l8RgGuVoGJPbh3d5HFKdW8akdvwMCxMk+NtpTmhwbq5
jWs2WJl4bGCKmkVBqGLD/8x7LItgqySeRYJNKumq1oe/A/YWiwaByOBuYXOEDTU+Z5o5m/51WJnN
jkd9QGQ7YGABu8gOOj8I9GVRhQjtrE2NDyVMKeoi/bvoG7QXD6QDUong+ipeurGDGOGILMYkg4za
PUxgbwZClOTzj6j+K9vDA9t8SdHRWU0cugsHlB3PrYEAEvWGSK4fP0lRFR0H12MVqz+37Rx2+qdg
Rq2HEey2GDvVg5AV+NJ+Aph6YjVYfr6xwLvvjJmKR0xr2CAOBxwJtPo4DxvtwJn6mas7SNCZ+sly
KIuvCIGBExykyXwhs/1ywweNwEicfCSKHSe2Qnc/vS1qlM19ZCuACYFlArbbMM948Y+BY+MsY8SK
MVolyxQcscui+f4cAz82sMz1WKtt8Wazk58SbEiUrOJp6+NNFQKS/GRK1KtPe8NOV4XYJhP5fzWn
jiF+t92p8zWrmVZANgyzI4lyaYl8xCNWF2QXUNimaN+Wn/r/tWIyX5iSzKJO7BO5y6ylj0Td3u2N
GojZMek7ndDnTJecrqR2GR4MvXXUZyhdAxVKdHjyps+IjjeRXaBf+JSphAfz9AEDbh8xWSO+zy1s
yrmeYQO95bzl5kPyfKNYRz2+DYSyFLo/KFqoJOJIeZJDN1Tvu1ji8u9WipRO6PSrR9rXjLLwtIHl
XScilBLHmwlc+v5XEh/EcY+3Obr0nPVaFHpYYpuaRgHieELN44SQi2MJZzt0hVuMaKx/xkDUD4I1
vLG+ofgrJe1JUEK6NyqNZH1iDGd7EREKgVRjoESW50ZkaAqbp+/XichJZ15+gb/IX5mOdsCeXemL
Kuv0oIVQGAdDiFBm5AhZFCEA+EdIoTIzV3k+9VAJwYQkt7FVFcadn22JCZQEf9VZ9aad1mHEg21J
7rOAHguaiewNL1/FIB5kPbAxaTvp5UntUIpivjBk09jSl4rTFkSskEE3rqqoiO5fXymJUTn3b2UX
wtdugN1IA0pLXsFaTgFMNcBQ7jHZMy1XgZPJH7S/LRmYpZEbLVGRardMLTkhMzCGzzheD8d3ACH/
ShZOex1Z/i1arBqIZoLPlWYFF6A6sPa2XHpBr3PYANqqsvquFZUpNqoWmtWZRSWzbYVC+/JbKgs4
8WZpfaBnzd23XB7karY1irG7m3m3DEpLgozZ/79lWEaZQQDcdk79NGJgmFyukHnCUq4FgoWMz5aX
Q9N3mQHLOUbH7Q/QabjkgZLJTTYIGwkGkULifJqlgsuxLnGd5/6EjzSJIwAex02xZNmn9Eq0F2b/
1KFpHUopwgT7qz3vNZlbuQtndx6bU4tGAEs0+Mz3mljWNM1bX8BAVGAUF7mF/dUOxCRDB3229WVo
BhRxLXQkRKxUYHV20TBsu1kIr8+kW7bIad5FxzBJMIH29r9ATlDzCLmmpMa2+HvbljNfkBlc1c60
FXO2Qlusa74yClnGToNnOniyU1m09K4/W8Tek3JL3M0P+MDsMP+AOLY+/90QkbCtz/oRklPwDjSe
1AMtYtKHhegD0882H/j5mKvb465QIK6Z828Hy5SNJuSsT5Dy8HJC/znd8QIif4vKD83Soz+YBX+w
FMXCnwGBZv0tlNgu7/DxJVEECsEdNeQnTVj/M8dHFqAuShYsJOqkltNhVA5er5yfyRg1pt6aHmq4
5kjWn4lFf/DbJdeWSHiqEfZZVq1GTit3Dl16aYPUsvsVXdJxe4ACKIyqPCTBBWTfh/hX5IAZBcF1
rts+SbUD/5NYG871fozOAeYdV5UjpozA4whJgEThjgbql8mY6qfgBqH/OxoN/sQFJ3/SSt2b8JHl
bNGwyqh0/05i9Ap+U1HEiTu7LzYkWNKg07TwUDqs79x7mibpjZ0hlVhUu5Bi3R0JzPWCs41MDBC4
E4lN8+8oqi6kocIdnXxUSgkfvmqAEpKGNg+NsR/xo1kdRH3z5kQ92Lx6qydNU+a/qbpwl0LCQdZb
PsJoJTFTdu6nT3mTQ98N1Elqsyxb8KlZm0CKfs/2Ws4tf+HW86CGk/7rrX77sndKhcp4OOcHuVty
oaFgQ+FYY4PCdX/7THlLFv1KN6nroIfAt1WE8dCvWjY4YPggmLXkAFNCmcZOVheYO/bDiGNYC6iH
oB+SojCGYLmoBRFj+3rLSW25XSCvMCZGDGKHPohDAGyEnDcewozYmTaqQHF7Zz7m3rApAMItQa3E
3WwDE2X0ILfxzh1u8h2Dcg7ckeURs8xOZCBAqX6S3D9PrW07nyNLvtMbkavhYj2p0fzA7+lQLueA
x9k+7YnF8qxM6jU7wAthLqXnk2VKFqZQInghzBcqdXtFvtpIVILnELtwCI1c9Ap9psBlzCJAnRvU
Iz2uuAy6IVOjmoOpTrr38e5pm4WiGq8vb2Ihrou2DJ9/2n7tmrW0prYicbuAfqTNjGuG/khaR/oT
wVeoomPqHmmdfLYdzu9BDKohnCWO9wsReKkMLd9aWD5CCBpzYckpUgoak2bI4KaaOFqc6859KaQU
j+kSLSzOh+O7uIFzEi/Nc17zLXR5OpiNwjc9g0V98UaVZb5EZyDFBsHd1lGpaiFYJkfM7dacQGm+
unMWtqyXQYKLgHn3GVWQwLo72yEClx6F/2uuYEOnql5DIIZKW3TpLCGNjzgJJnqw47wodydimS9A
QumpCY4Q4gvKTQF3+6Spd2pZSM730hQsX4rK63hu1o2ks/ZT1UP3PHxbecETnTU3JvNZUB4MLef0
mh7OaG/gRb+3tZSj7vrCUO0Qynb6rdobgTRiaEmwLxJluYEK5x/nmvkInfvUpqg7uyGPp0qu+PD5
0blH58ZSkOGsrlHNuRafST7aXMhrAfnl6/5Zjg6ymzRtT5+cnTsvdXd4FdP/S9vxibF2RpJkgk3n
456GT4WchU8qA/hUFJub/qYPt9Ngim2/n67Lo1KCTZaxWFYWRczlTleYKv5k1gIFI0MdgUlu6Hmx
lT0AogjcQNo4sTVnnSAtHc8xkicjiKkcoaft2gkq4zmuo+4geHiLMRRI1JZMyBBG3XT4UXJLycZ+
4qW5CoqAzJRm5+6Nq5ONIY3id0Rmo6MwE1knXtIvv4Z9DVM2rb4sExHZAOGXXNsfQ3MGigd7FJH6
p0vNStaGKy3juyCg3zMnvhjCkQWJrKhoBS6vzWSnUMuYE3qSI3UbhHwqwK61nAuvd78XEQvZFeyC
IsDtHuFFYSyaPjmmbH2Hz8N4SUCsomRmh0gi3MtkmP2qqsAzxyFcXYcBQ8DPQLh0qjwNsqLGqFPU
xST8D9VB/28wb0thl4RaHnqCYbYKzl4Jt+yij8pADiWDyM11u5++QUe0jjrOuvId8/RAQ2PUAfXC
W5DAvCpy4Z7SsT9o72Y3+glAAAH/yT1Fo1Yz6gZTmHzE1cFFLESWnQSdyV59/+F1egrAiC+xlqCj
bjf3FnVAFBNBVujq/jU+zSRPF9AP+Fz/hd+1OhyfKIfBFO0DwucjwwJts2NnxWO2eNbLguF65WQ4
qacnI/Y7Z97O8A7d6FlKQ3+kkhX/55Ju7sAZcjVJ6R/3jf2bZx9t2gL+lYkUZGILb4Z/GMVlf5RR
WqfXQhg/52GelbsQY2lh9hFVFYRLaN2ODWmvh5gd4mVGj48eXOP0lXsuKGB57HDktS4s8cgFzGAM
FKOXoqcCQozaqa7zBB5MqguKElal43bGmEHUx3TaKGRMP+/tlSrjtzUPa5v7P4Y6kvDnx5c7F7fZ
Mwv2qgWYePWdpNjB2uIp4CVo6iywGyURwDhne7tUNl24AWkZn8G0zmeRig0Vg5fSRKAbQ7i7xTBo
3fRcjXEQHtSjsY2y2fEwDh5q/fXBCMNL5um4clfgaVU6UN3g9kOFnu3EA3AVKwmfQ1xBNZJdsMxQ
i/g0jWKpZcjPYvdTLTgfOPxpA915zh/pf5uHd14WUIeUzZwBZ7KdQoRaSCzEqZY5BtMwmguxJOjv
Fi7LajmcwTJvYurNb6sVulkyQnncja9jx93CXJZH2gbuTQdMNYufL5LMa0SRs6vSfvWnZ1O2INKk
o9oQPGUj1WNVzj9EYSCY+QVXUq6T7bnNAOn7iYGTRVsSHci1qYxw0MCmZstL4RSFmH297F2imEY6
YYWCWSyS2rGRK2VK5j6tyDMVO3F5JZOD/DeEag3S/h2Hse4FcA6XSMDMI/J1C/b2Qh9DUAY1CD4y
WOufHDd6QmD453QJGUo6UsnNAu1XuAVo/LjwKHHA2P/bdTb4oZ4IBnD4AuqBjhFrhqmbhlfAoPgS
5EpSegJbUL3FaaQxwASMz+erdemoLZWhMbRhS7uMu2o7bIH3zz3gKR9DMWaHBo1ulvr1498pp+Yb
vFD/+GqTcm461W+96qSzQDN51z6f0tNL09p8jKMmWGH59MHuKGgo0o45s0bMOO5J3FTR85o474s8
toMQ74QUSg1+heyC0EzmNVMIrnUZ4lFAZHxOb+kpw4numPYjO9GI0pAr18DDjfSilMnhzx2jAlNE
3GSpPdUJN0cMmAT7iISDqf7D9ZmgFXTCeFvWGl01LLfykdPdgsUCiCyAdM+Ns+rHaL2y/guKP4pH
K+D4B2PmwuR+y4aypTVML7g6rt9SUQ2uyiqUx82HZbCIHQtGLZALgb2yMZexJnDEg1mLea4UbFQA
hrQOhthpoG9KldBzGyiQ6Gstb16BsQl5iar6AziBdzNimKEtKoVaE8SSj0vRBgQpxtKp5DVmL/LD
LW0+ObBXJE8CrAAEJ5l0itc80qv9ncR0333rCStwjPk4jKBuerUT2Q50Dk+JxMbh12uPjc1as1wg
pjJtIfEw+7Fco/q+s0F72Agne/MSn0lZSslbzcB7jQlOzUu6islvRmzxKQL9FzrxoFXn2KPHNToS
VTXnWvqAoFb8eQAoO0WFtCdQ1p0cpsMKbgr4m+RWBkkxzN2NuoHUOO04vU+iTzCckdHD9caQc/I9
0XoIQoSra9Bpf26PCkMGqaRjr7kHefGHIQ1Rn5a7ImoV/0dUNmg+HYup+Q4dD3f6D/F5UTZ1HCdb
lI4V7CzUIwXiTiK1dX4b34hZGZd2HbJZlVYGwXxrTqx2SqqodZx7nldiBmuP5ydjtw/eY4NgYHqH
q4IB9kDlec+DhQ/qCKoICBHPkw2N0/kbPniLvpRLdw/BJjYYdfZ5xBM7quu7j6krmilGSxGodTCd
ubhWA9dMckk+KYSRvkTVsjb87bGBTkvr6LqbzAgcy45q5ONU7RFJrosUxzBLt9vOpjNtcC0WZA7D
8laGKt5rGWdOwKSosK65mSf//0p5Fxb0EvXrF9UjhAu6I8DiZ2ZHyJUHvPjG4F2vBSVCql3eDW7o
LpNQuUb45qXDo2gz7V3/dqpF76mTNafnI/s20ea9IJZ9W1UhVMmIIIb+ZkBureai8R47pGY/JOIk
ZMHP9HPY30RsMap3PeiBJfoMWVuhpTYZDP7WsmLwrE+AnR+n8dRx9p2t3cgWwpSVkpK6TrUj8Xm4
qFMmnHfJpdgcTuILCXe173NO4HnrGR8t3bPnbk8KMEAbsRCHWJd9vzHizYq2yXRIr7dq0WmoL09i
6p0S5u9O3kwvVRVQLyHccr2VtU1jV9a5fndp5G5GZTxrr0E6LD9kyt1SnkkpuxbKhLYA3OWw217g
nak4bMtIaYmcdzCsK/A2S8AwRGiLFr2/YXehhA692MGtfclmojgMjFAFXDH14SuUurxxmye0bE2X
GJ8AxxVLd4CzfqUCZIfDuJGai1N8MweIV1h7PD+RYQwfIf+QYfkbgoR4aC30rY+6S8vHChPbzwEk
dYdjdAagTuQtZHHrS+5EkZR/6jYN0U0HZZ2PSWsbgXk1IL43Og5YNB6bDxSPkoL48xpqsLUV84vp
tfO/FdnzYaRp+ZBiGiVItGJix3I2qAnXbmge6dYO7WUTzQO4hNygY0+2JxfRXg0PiJu6mkWW8Fuf
mB4aRFWbpGIRgZxYP2DLnLbDambST9ebfEDFR3BFcfoLySCkmQ7a9vHj95F0QMVRGjkGb10bhZYG
ZvYCw1aBwFF0FndU3h/TDMGnlbKUVZsLM+BY8B3XNP/61av9lwxxOImkq/f8RDLC77TJJBlqN28i
3HZ6VJCTAXJF5DjdOO58IxQ3V//V0DvWgj2Qe4ALPnsqvS3HQCbhtaExI520YY2mLq0GbgxSumnZ
V/x4HxfONeomSAtMsilAXEHftd4AcH1Z0vA0lV+xCjpJfEc8Skh4YgrctjLns+2jwZo9DCznHgl7
kVhIi6fOeLGUY14mBoh39rzD8j5hZ9jgijVCXKLW6xMvFBp8e5Rmmoh3ZkW4+y4kWimGieJIpgR7
JixgnBnJal+vJFgG2/U+VhFoZVSPuv1qgA3Oeq1G48zwaWIRuvv2av886aB6/ynHxEbDNyU+iMvV
fPi398wGax69VIDzDWkGR1dr1visW1Q5Ez+dDSCZbYtMTeYeT7ei++CThLmxs4cQZu/OY/oDG/Ef
Jyt8b2KcKrsQrt16pqPcjjw3ezKObbRmR4g89n5s+PUmthRXHLteJfoC3Py+TL1TIL45dxHrTWU9
mo4T0ujUJRNiutMERQRSA5Bn00NoS+Z6noBsZ3RnuPCZKpm1XHYWhnjfL9/olraTYEtj+2wdJ2nJ
OuuT3qvJWcGtSvo6ZHRgCTt7u7pbmi3xk3wVVBVtrOrG2x75VpPzj1p8JFLS1lLRBuUOjxdFubmW
cJae6W0hEeAjFVZ9XtanP2OvNdWp7DQZlvIrCAH9FRcntOIXK/aTxb7ZWGp1BFiwcyxZWHivEF2F
nKdMg2mW/N1VaAIV78AXc5NJycqKxVzec0YwzDbjPvAo6kCe6uRqHSoy182RzDPrbR9T0loRuCQm
oQMxpNdl0iCURdDVO1msM94vMSUiKo9MmGXb49BjXQVpEmXsZ71t3vHmh+Fo+08Xfnw5dYwMKRE0
cZ9maP8GuxtWxPW1brdL5yiAmiX5rrY7EKct/gsPbfW6CNYBcvBdBotzjRsdEIZi4HtL6MvYfoyk
mF790NqOBJHu9yTUkUkVGRJKFm+rOow2Wwu3lCrmkyVRxkB+7VWbWsvVq3f9yYW7qCY9K6R/4LAX
6KxtnHCzwkGn3zWIi1Y9B54X9yvM96mYomPs+l5ZfAkBefrdvDzpowhM4IelRb/ogPMOzq1NLy2h
g4kWHaof+eVsNC2f86ZRm8Vgv7CB+Sj5Fld7FYNskCB16Z9XYdpsBv3bwvaBJSds3TY7EwiNhQAR
0FZtBod+yQNB6uV9TE/Cwjps90Wd5czMaDfdtrDzp0BujQXOFLvr6WCLpv4rUV04Ad14u5WVpa3y
IQ+G76x7Nt0JpMIrJTsXoJK/XIXnz/62BS+aqLu5hWQo3Eb+gOAQwuWdVx01Pgv0tZKioqok/A08
43u/kAUR8713IZt/pUlnFXHgIYMsAhPfq1ecRQ/G/USe41jeB+8qZBX38lKSrCOrTag/FuECcJHu
u61K0DpzeiR+NgMKdouKD+y+BG5Rf/u9GKAmsBElcuM/FAEwGVd7Zpwfk4dwlTXCq894Q9TJMorF
tq5O26S8yanaKUU3nUmoSDmkDx8ikXcQAVfYfgKXr/pJ3YgMSCAtsbFpiwYVUChaW/zYKbR3eHpP
jXaQXxnBTsHfuMaXBCKJgwmKIiCm05+PF2b1UfhW4k2MOsc2FT36AihZBfEuHCvZyIYOY+mGvDnH
xm4+Hx8RMLIrm4jYL9J/iGNnDA4iA7P4MNU3U0MXfKWaEAES/QKsG9q4eLPEAAxsKZNORF6wxLsf
PK09/Aa2xaksDF6qgQ/eq80e7jAmsVljxmTkAHJDrWj7K8qAYadDIVC9cVWPDZWx8s6MptlUMOBo
VclehS5VMPVveccdN2ZfFkf2IDPl5Xa7OBqJOoPyYNiJS5TMQUx/e8vs6f8m3R93dg5gcsCMSXdW
MO3UxE59biggzu6j9TIRdhnA4Gsmlbd/MrDwHXfJL3WzGhJfe9c9XVDnIDG1LX3lQqDnz65lZ0yr
Jhhd1BD2JqbceWIF0zrdGBDNz1GHjbeOfCF5mJOooo4wStW4MOIKbWZ1TWeY8kjoLpALDDXOEIpZ
+bBSzXSHUTF1VAMKZMMFXWiQz8iozVWRui3CbPkHo/Iup1pzX1FExJKjtb58Ty0WIExZAuoM/mOx
qqmxEGoiP8x1bvFO5LAiat43hRPFbcjQt99PkAkRrY1H6yUB4bQ2vxqT67xyCaUGOjYZ+p34DSG2
GBNjrQHJpR/GS/frE+I83a2GLNd5ICnJZL5rSLNi5I39rm2iu8g9A8KKUxhQHCRe0AcRX/4q+9PB
trQA8T+QmONJThRykQz9EAb1foR+xSYeXaUjJBcHR42xDJO4bUnssXTmyQvIXX+IXFcu5gba6pXU
twdR9GUMQA/bjPdpnCyqSK3k43by5GVujJNb0ebNoJ5FotgnS+Tnffel4rEwAJAA6A9z8sCszexb
f7Zmp/qA9bhyW6BzOZSdnxIi6UE3Gr03FIxaW7wUiIrSDrkNyQu2QQQyPQOkq/H8eZ2YY5CjwaV2
MzfawEnW5DvipLDUxBk7nDwh84fE+JpBOERJpvwnn/9/ZtVhQ7ULJ9649+41a7aqToZDOcs1sea+
hT85aP10vqZi9DKBmCeEaS9p4i+AeIfNDmS3HrWTSqkBQy3FpYwqkiWVzGooyBYTfpxo9OTq/Lqr
WNZOvBHQIHS0l+ptmWkBFx60ofuTGqSSTtGYwqHYFdOcc6AmWzJ+9qtSgevNdtuJkJxkdubqOWJ0
jlIWPSAqGjpkZ0AbRa545S2xoCMwrMldahGHg5lf76N9/7PD04N8JNOTZsGiyAp+UmBV9D7dD15F
+0eBAqQp918mSnne1nS/B+pJmytaZ2RJdO7qOvKaMGo6mRqYYIcr2YSG9npquyQlEF9ct2yTsli2
Oj9RLrx10vHJAFKxW6BkgLf6lry1SfG/sGaJTzeW1MC16ARw/yNOUg3cKpm77eE6a40L9NBwjLD3
exMSRVY3Ej3i+WdZ7u2VL+8UTbyXaNUiHCDHjCG7QTrDsAipWxa5U8X12mjzWXPD7x7be/sbfYxA
VdlSmPH+F6d4dnhzGuGz/tuzIH/ivCK46cajDk54apwpqyLVjho1IEtahjLbyil8WDZh+WslsEWb
csu1DfGciFbcf/nNLR1tAoYtWJe+LHGDbfZkQl1PQfr9h6LMcsd9p8i6PTJElSwUusCaGFfS5vO9
kINAHl3CqRl8wCdvlORCXqVuttDj/IT4/87jvpUDq5kSevt/9aKIt9iNrRim1Up0XS+nTSzLyC+3
vhuo+h8Vip1GQCrfUZM2rxeMw/F7BbekH/NOV7bCnzOOxiHaimCarFsoSkraJyRjZOr3/FUBJITO
oQlCGLymDgYi026apjce8YQAxo+zjDAf9V4L//VC6yLMV/wS2NLsuXJj9EKXoN6ghpO1GBu98ott
ayE8uiUkc4OclT3Fdrg6G9uOuLdeCr5tNuAxg+9C1LXbeOohnn1meQ6cRCk2nCdPQyDQMhW5NKvx
fFk+L8k61GpzaSJMGCh5kwK93LGw659huqAc5qUYoLD4rmQojbMyyXUcNQ0F+yTgsLIw77L+mgW7
oamJIiqXv4uZ4ZBGkf0zHgdyibIDlzpnZ/+T9Cs9fkakwKOKZsFgC7kDJa3M/OX84FYC2ftUFCdI
STAZlyHmx4IoN0eqjbtYMY45lIpFdx/7NBfmsZz9uUUKeFkls05EjX8q7zY2d+2dLx31AOK1IZTs
+7djdA4gILRgUDXTdL1m0/8VGS+OXDrD/VdKtwjrUpU8piWtBR3HNF7d+eus6XiYfa/Ro9bDa6Fq
mpscIY6EK/udDcgt19lN8E+tBDtAH0PtEp1KpMV2ZbD5xO58e6sTI6Gz89d4D6lC7o0cRBTh8uau
t2KPZfZj60vAw7l9ZZ7wHS8+Y6vivnIe+1PJq6IBLvEjyWrJixyqrHRZiDhzNmGEiQ/ojYFavr0p
ghrN+xqZeDbT1pEtXPL8hTGZwtrw18bu+8oKAzsk3Of7iMh9dqTatAZ/1Mjnl5+5d/QWjQTccT2m
9dt1jAQJ576Q4yr92nCjNbqZCWesq8Wldqy0/8MCSJUCBQeH2dSDoLsegCpdIfYFfMvsnz5Uxnvu
BnjyjjaMIX+quaFvqS9HM2nYpfo1nClw5/mG9G5bvTWqpXpx8tPcFe/PahNKTczMPqr7Q2fyvY8b
6AKNQ6BjVlmb3XTbr1xA3j99PreS+h+Vvwkv3PwvO5o5ZEzSoGDZLPWczjNmmz/Pgu1aNo9IYEKz
+9I6j5qk9FQdOcGTugFRXmgDcg+Eh18aVCkG4VEyijEN60fjv+tW34CblnAxOtFx3qsgfFQ2voTG
oyuArO/UqPR7jMT6ICG+Kioi3Cv+9da8MC8NkDEEi5xVly3Y/qG1I9QqipowJWwKC/RvTolqgEne
LHBws/tNq3dywyafsahb5kJgf5dpXxYYcr6spQpi1K38lmmoUwiADYeVyfmKR5UoaJZtjBao6Pni
6CRT5p+6OsV7T0GjQAgqZVaAkkv/1v1q9SslyiRbvRVJhYaziuiTroUS+k6ovba3BhH9d+w4S329
oGcBrItd4ZoxhFwYl4E8aX8DHRmuQlM4aYjHBQ6H7o/IIfoSv7NWV/Vet0QmGpCxtujuvtLs047z
tZs4OgQ3uBwMyZ61PlD5S20PF3+aLCctIQ5OGbM7UOD8qtEGHQo7HklcNh7UwC1alL7+P+a2O+DN
KLhAK1O38zYOq+zg7/4jobSDlSaLn+WUIj5fSU90NhV7yFKLFFN4HWKTqBqJthrS4fRezJp3PlRf
QQOH9e5b3LUCZniWEeVzIgprO7QdtpCIFic8eio+QWfdS2XjZdJmKx142s2NNX8jne1hPkmp6tr3
tpV+c+uTiaKNN8UBjYHi7L88Tn5HXn6nv/d3zcRdCCmpAFvQ7YOB4dfQuzzOgtPAG6on67UfDMr1
/bClez9cdADgX2X7K1u1yVxJsXuFmNg2bAoz8+Ooy4JJltuB/66YtMkfekZF0P0/2oseLtrxKnfZ
uo/7VgEiZn71i+BPFgHfM7S7YDxbxisWPGHqZfnLeWxsqGCZ1XYMln46m3NA+KEWGU6D1pFh4Jzw
sUcpH/5HEShqw21dhXio6vhoy4v7OEtNPNfdEm7CmZ2BLvmTjehmAaVq5zn02V6FrfnZBFeuT7mp
rcgXz+TyQ0cq1PPMYJg8RQqZMM6YC2cXyB6d1fmDH/P5yMLE3XAdNopmAPPq9hI1K227erMjJhzI
/6QlXiNs9Jz+HNufAhEnTzkaUxK+lejr/w407+VpacR0v3b+End0uU1X0AIjm1B9svrIGNZ4CtzO
Z5ineFYsSjOAifl4Fq8E7v/AKqOh/isNh8SfPoPyMU784m0ToyVz9kSQez0VyTD3bzuVnfM/kBsV
MQTTbwqPipFqIm+jk3wnDwdykYYFgk73WPuYNcUkQ68PuJhBb4qkiGK6n6o6sp/nX07a/E76LxKA
WcGOA0KEXbkVnd7XPe3IljoSGYwHt5sxRIw3sxXWDy3To/VQYhirMGVbVLOTUvTD2GZnRptc39NL
Cj3Cd3skn+Hd7pf85683JepIb00HHUO4O7lPms+UkR6zMyyWBCM9X9Bm2p10pGjjBiRj3JedRC4G
Vuj+dRO/HVEp6fA+vzAEZUqf1oMURrrsc6Ji7QMLQ4NX+LhC3JvDiOlWBbs/R4B9dH/z/XMsoRkV
rT+6eUw2XF0tx/iM2cG2hqvjXazP1p9THnNA4u44imk5S0UY9EfGObK+71YdPDrG4Tmi/fsa6Mtj
/yy4RBsVC7tqWWmpiHVpDu4kwkX+fOaHXOi83KfRR4W7s8IS4OeRImOlTOpc9ULH6n4ldG+KEHkJ
gk8KMMBaBYIvTMBu8beZmJYdygvr6hb9Z6iAYEGPHwwzfwsOOnm8WsEDVucCRlxMrHzgKCgiE6AM
o5LOsrnwQihhU/HALPN4KQYeKZySQvFp1qkk1J1ELur97h6opMAWR8z8xjG1nQrrB2fsaIq02sAR
Wfc7GjH29eC/06CunAEj4XLLXhkdV2rRHznwm8LpUDubZtiW40W3mPgCB4DmXl0ubNEG5bOyDwvz
/pPARyrBzKzNVI7sarURHENZtRnB9zMlubqmc1NfwQItzEFK8lKAXy6W5/MYlLQr/HAsgcOnBu/D
YtmKzDdjfIyTxRKZ1j/ksf+48NBSXTz6JMS8rTzatT8huAWjIPLzUnnXwUnI++IANhXZ9bVChwq1
P20Sv38WyAsh5z1Rhwyxea9bg1+7RP6H0dMmKUI1s4AmbKY+9snBX2Qtr4CpU0+p1kaibQ3z2Rsp
pOzjXuGRpD5tLoggQlEE4SaeTaU3gO9Jq3sHQyJrKOjct/IYHgan1bWacZMaILjxbfruwP5idEcm
JQQkwXBbX5K65SyBCPBP5RDnCGb07blSs+499PJAy/L/2MBGhp6m/C6yRJ2GL9rpKl5su9U+f1zF
eOzfOiC0SDfzLevC7kModQjKAYxivMrAaV8YyeK8IsaQcKXqUzZBVTW0SX64s8pfymyHVJCbxw8h
MIyDx34buK3yUwUSQ6Ldajz+WhErL6b4Yg+QJmj6igzrgmEQWSUDqGeojLqsADlrLLW5MM1hEp0R
9sqja/Wjy0Z8R7KjFYpG6INeDua4e0J0xoFFuHpR49k0oz1m1CPI1/xLBuScpMTHLk3C8dHU3vmm
x3L/L1cJYGkHPmlwXpVZ/xR3MOJnEWIBEjDmP043wPRtzWu3KsNQwIYLcEEwjbw2u8J0zj2VDGdQ
G20FqeLMQpkKFRcBfkgc90Wwj0mdjnX0C6kTDh5ta9Q/drY36vAiNC/SWtLNKH+gOR/cHqV5vtpP
2cnRPOuJqSCt+PrCYIS+G7C802DHZ8JkgGKrQ5W71bV96yE+r0Zs4Ve3NxGBQ/4/dkj0qqRxiMqm
vgz4q9ZOAHVpb9GxO8ZqDVoQL8kV4K7vKvlcKfSwSQfG5XAeV0Ikrc50z7S67oHNqiBcqGxswI6k
gp4VZ6xkmVJNEUvxAI3sVlXH3qEHM8bgtIlw3lH8aqHi0XAs5/tTsVY29HKRTxFapaKTf2kMqXPr
2GVeJrqQn2AUENh7XksmP7zVOkVf29VFcWW7GJeJwciUPkMgyoNbin+rThCvmPMADWguhx0Wer7c
m0HpuGTvJzG2ZvFYbjG2BCsZwddf08xDp9FDNIZ78bUV0HX0xk3xToy1IqFoYUNwNs4I5nZ8Fs4x
VXoRILUeN2R9OtnUCIfvCbFuO9AHEyPbwqgaJrGNIEDUy9hgjeNDURRd1+ObFfCU3PbmOQ8CFXYX
bpL5ueWsFxxjIvz0WVaJkJ6PpnbIlSxK7+vZ7K8dP6OeWKM2DYJzoNUAMWYKDzG9kOcZ2zkKF1Jl
h0qfiyZUF+sThDHibhdkPHG7tKHSSz38prZ/nK75QssCWPXoM5yhMg/U8n5h6VGFHLRtADDHg66q
G8q+b+D3J/YhJqLiX5joCgKRLjBWnYL2eqEmd5Qw21PvpVwfOqKQDCVhkz9ARiA5vmVC6BjTDod/
vJ9Q5xtbFfgU6YlhVj/QpwJv0jbALHhTxDikfN1Mcq2eKwEULUUoax0e4sZ6KzbrydaUZc7hiI4b
vdbsN8ke3La3V6OYN1ePcGAg3zA2y+IzDgKy3bh+Ou9bOc2b2UkPcmEDp3sEJnYKOdBEta+ztkjf
cML/J8zmU6YQN5mc86NLU+K6EiRPsNEYwYn/oK6t8xaWWCjKDXQ1zSqFT04p5GUzuGQYeo4Uxbk+
djVWWUnuZBQKquMmA6Q60Hg82AvncShWGrgiAQadrAOLwVGwPg2RhfoQbpr0wWs+R5oM+51oUD3J
K08fCMhPZ7pteKBNy9JDo5bmuIBFe2+Nb34+/Auh81zCwCYi1K0P/dDEqYtB2sn8p2t75RfjNk8/
PxnlBcJ7EhND2UKWTCx9xQHo67Uzj/htlziy8h+uH3ZP2C/LQu2ZMmTJxFE3W0aKJM3B8HIRu6KX
MThy85x/8v1xmmP3joW2KqYyDfdQXnSpKyvZBx1JXpdMW8gLfC84B7f9y22rLLAA89/UXd7HA8xt
cqhfqO2jyvGC0WmEX2xlTd1TY86XEyV+kEkqK6HRXg2L29XEV4rwrJi714eXlHUfB0+YBnWZXalA
fVupjJLpvUGctWynXDlLsgr129d7Ue1dXdrLVtv8pQH7VCLEV/pMwDdr9b5NiceDnorkJnLSrqth
pXNWG5PlPG9N6jhTI6BaH6I+YLeA/ADJ1RFQASPsmQENbHLO4TWZ+8HosvkUuyBID8Yd2JMtAZYx
uv/KTURi628jvWQArnkkCInv5bW5VbV6n6lPbuhkAp3Yb0JtgLMXWBFxKLO8OtOSjIzv0EWbkgFQ
uYq/QKgar7TWsa8zcNyk16W2ANY1M3YM9QLbOnvVa9YoXIDj2a2pNEB8HXd4N61FYvt3fOZ8mDlq
sRGAg9Muhtx6rXA45drjkXpcY4dyCpEAsJTYpKW72aZw5IDGmHgpLQV+mY5dBujxKXlkUesMX7WZ
BNP4kE+k90teywJ/cKtz/xUXR04HqW374AdqBHor1mzHT9EuleduePsHCO+42GHQiG5YHu7jKTGm
devy77fCnixS0aNCwwjuqQRCw6U+1GfKNfdAMbp3NTiv7QzQNnctctVH66QRGnnfaZoMJxPK5Wos
TIH/zaPRZS+BomrnnWXZkQXi+mnVRPNCR2Z0YzEkKAWF5maAYiVIluUBFHHRtrasFdCWP7tGJ7bk
9BFfzk0qrhFocGk3gkxWlGQlNb1c7GQ0XxHdwSp4SISlfL8HBcm6Y+SR++bVpUyhiFZzV17Ec7nC
nSZIB8B8kS/UHEVoISuzKQ0j95SndmYv50gDXPrPFtoVG2KY0Y9N1dfwHkvF29h0te6ystG6BCCI
g5xdD6UK2zfxotrnSp2KFMAK/cRZhyaM80kcP7bho6jrzOECjtk9w6vzJ0gDPbpFg89wOfMeCw6z
dl0AExlYqgM2quot+/vp8OSV6z490JrfsZTupGvIBPg4I1rwsVNdsEm+4+Vvfb/Q1+BQtc1ZSh5k
c9WWwkG3/v+rIjTlHihchDvORf8Hz2I7JWGEdK0F9Qx+l1yoZoupI74fEIUZqlisymi7CcgzB28J
M1nfhJG2+MHu51/ni8POZAHU4UEaZVXb+qqe9zzMM3xo+hKFXbuKcVNltghkn9UwnDRp1xHE+4PX
LlxcDG8erNbYF0gdNnqMFi5Si6CjCJFQ0wCHGHqTbH7WajNJiwgZ0sWP5nzmQH274sKkqHL7cjgr
aVXtqOvGqofwAHPj0xnewR0SCirl0lRuLAWREpnJN1tGlZV/J+TDffkpFcxbNEbhTiYq1btJdNmC
CjZ2Be89Yu0UtsnjJc6fH/sRCPRWUTWWl40w495EunDj+mA0IKLxrQigjQHHtEdPlPQZkbSCnywZ
K/yp6jf78ayspa7zoOFjCnv4FDTsJgLbt6up3BORcQzh4ollT4aPWPFqOhcJPk/YhVJdx6VcNciN
Wt8r0udKQZvBw3xbj6mN/4my8fbYBnbsedyDV8xLXEnI4+aHQCGJbMF3I+DT7S+2l4bWDd4aI1Jo
BRUsAeZqoHxXJk8cCCV9aSWJ2qE4a3VrrQN2GVQbubHJ2Hc/RlWwHdsCviPE/QWNLoiOU/2cpQvc
2wtdu+LwBFJ2mtM9763VKyCN8drjgJl20OjUq/RnpJJZD6ubZLNHrJx6xD/v7Teb4JTmF7ad4As4
RtvgdYQLVmOcwAhrJLa9RgQxL8ivaHr4Ff/BLAjVC9/emx6/FwnyId5DTuUpZLW6113dRYsxBArP
SvARlP7VVKmShRNKQbkhFT8biOfR6UomowKXr+uVrZO/z5qoGv7NiHprWoa8NcPG+R9f/z7UrNOM
0w+dYhENiZC0IxpN4Ijz0WnxEQLMDQNouacR88c2RRwb71BOogZM83ZHOswWXcJQARKL17F281/k
0icCgx7epw3kaphloiHcmWa/f7PwonbswOxdP0OmIxcm8ZC0+5slJcpBCeIZVoMHMTVbeO1ywpP+
EQWHa29wP/KkX4FBI93oeYWjt1pqANU+T9OZGgsAeNkscr4HrJSmzTIYfX3SkShP99yE3CCVpE0W
V4rLFESHbJ4NBj1stDM06wXFYkoHOsf1fw9GofDsNXWHIrytCnjnBiTfvfpo4Yfscsv9NbU48Yt/
658RAIDAWsjpNl2GBiOUqwZiJRVGNXIXpaJdBPQzL2fE5FHuL095k6vP0pf8FbDTsNCz3Pg1zNlc
vY1HumYUTO2mYpo9+FdbgBQVk/pXbNr4Y9xWKRZ6oO9NlhNPgfBRArzuZ4TWD+ms2s3ZFq6ur8ry
pNe2ZUtKdaq40Bm4GZzIWmOgcarUFvm3xR8fIF4GTu2bAV+7jCb4gnntbyIsNWomB919bBf9JNYV
O7yNF0/wp2n1Nis2MHhT03bVlS6nzlLzc3ah+i4pZ1pL274GGqopN44tyEK2u+pKFQsO2NuZopLO
wiLA/8qqL8PA4BINnWzKR+qV6H/7rcIy7t56vYYQURFadNevifz6MB3ayfmFUYUYQ758CRYDPNyA
kEaDYH4nCfY9OClycPHJoZxi3kwozl0iy0ewA5naELA/NgL9KhhfGXXXgIs58OJ60iw3JxVJzjL1
5kxcPaz8EMPJjwY0Nt+ye71ZBj0AEa9OOubx2euIyR04OrEmJWFb8JdII+M0m/cl7Nis0O6zzKGW
2smQnK6olRh16A1YsC31mXSnJKXarGGT5HRPBsAID0pV56RMzSYaHf2gDy3IyrnyYdxh1z7JlQ4k
iPPH/K5JETclNoQZDvfWOK6mOHbPFbWiSpzl4kyHtJc1he5htue4RwZrPOX1vAFndVQI/2mf9XJT
U69XnMOGA6HStVARrEJIk2lm+tgDYafJWQoVvMt5kNTFo2aPqZUixLJKxtgOPxRyeA1O2/dn1grN
3s/cQHS+wiV1dOZNikAqkxW3ytbBz6p3nOQvUab6ga+HKA0YeT/zkRFTh2VT3pwN7KSL4FdKTpqs
YAkkhi5u6jhOyfa456ddaskA68CDEBYPkJV1mYr/TeYcXdJx6HTdaqgwkiFrLu0GoxYftdPiVEE+
DnuOK6n27zqMFHmtgYZHqGq8NtwPSaHmgGYUjyLugknkDKuoSN9ydVzgvNzW3823yqVxgzEn1etf
xpHxtp3nx0XTHdxFLVilQm/AVa3wwvPt5qVXKt6i+m/BCN/CI4x5sx52QU0GcM+xBQ/vDt4te0oz
0wTicDS1T1Cpm5fZ3OjkijClkhlecOQJ+ZwUyo8Yk6lUXF9xFplCgzBmFPW690Gma6R0o0T83q2d
7TMjL+BE5iFJSlBCVoX/brf3AbbwHD8vETHzzwZIqiwBo0P1eWpWMhB2BYG9Km3AxZCzp5lOcVFW
SOcWEyn/c6B1xIa8qBvhWswtdEUnPV5pUubTOjXLeQ8CcThfMTP1EQxvRwzczAbxd0AWRh/NOVNU
yLNi2bgtTEtW9yU7Mnx77VY7G/il6YTcT/0YE80gfY1vDCLtERsCw77vDx/BZmdNi6Iylo1LFq8i
kMcURFMtOPMn+csZuX7YP7/ipTjEZrtMk24RY3W46+jYWs7JQV1/4s0ftOIidh1nqb7lp0/0BViE
SrtCCC6ZiEZ2Gb5+SsWip43F/ObI75W+38Dsc8wWgT0U6G+qmvMdjKtCGQbg2mlPuc1FGiH/QB/a
FAUQ9IPHmMfV1ffV5iApmaQR63B5KOLyWDGviyScU0e5iqepuCzo9bj8slYdIPwiDzr9nYSjBi3u
zheBj8d1CgleMKVA+VlCecdZ/plk5W9ikhJWT24G2MjV3ALrs9Xgfkab556pz/qxQetdBScydGJp
b9rAuNmN9JwyaKMCa/0VaoDEsJ1B5VXtJQfT4HaKS5EmI1rLlt0+zgsSZw4i1UxFoFRJWYAEAKSf
H+SYu/Y3NLEwEEzrSM8Z1UFCLR2o/FchLerUkAgOerT64ND5bGPxSX9bRETNvq/i9iHm3AyU/nQ6
6g/rwd3R6Jlh6RBBw0aIlRAQ3NEVWvOD72M3YYLbarG7pXtn2eSYyDTiW6PU63GXOljZTPzG3l9l
BN8k/mJ0mlT5mvsIvXtKu/v2etmD7KuCeCNlDsWiOLUZ3GMmLhEmJacLRbpCT29sMmLAWjFrADMv
bo7j7m++QstbmsVaZohcqSc/6BAQsZdggW1SzHW/NWKYO4NDW3EhcII90XGMl5Q14am/yMNIltXM
AG94XKXmp96veZx8ty6srb+FSAHRaPkDD5qeqsg4iBQdb9tNf0cTlSuJB9bA3VlweUpEJEYb/I4l
YTz58YJcWFp0ht3N5eJmQ92VCbm5e8uEe78FJi9/saRuqELSldzePeaAknwTLwRT0BD0VcQOPgaH
tXXDVF4vCCjkn1EK97vQSVTYiZekovZKe01eCrF6YdLCvPNv3B/eSTt95cofLxNOY9pYtu8Bn/bh
1a3pjTESepZJENhGwJFIdSP9fD4X+62lg0sVgUtnytjH+BPayFA0+9CUWm06WzJujwAba1ebW6fF
MtuUFT97Us6zdK4Rv7AKt53UHWs6lvE8SXsAfcdKs20w9Q22ST6CxfVn/a5Hm/JdrPh+4f+VwZb3
WQtG2yrbQ11k1zUppTgaNT5v1wN7bmwAhX665VYw7yUVvXqlRqiVp63iU6s0dKEFkr5MSSDFJbRK
rjh2+O09nNL5jg65h5VPtE7+Rx/s/PN5J6ciEjuM4A9n3C7WvHjR5h9tplvL/ri8EIN2LbP8x+oB
qKqaaXiA1bOHeJAa4kuXKr+SPLg0twsbhyjvOY7gpmT904juWDB4yypZKDlnLw398Q5BooEgDh5F
AAzQQXUijmaX9+6DvUjUq7wJLPHY11xDiPnLtxumvtH7RNZB68oLzDOX6sIfj4eVl9Lw9nEqqakp
LSuHXFUaynAFBmsmBJ6wx3KEHjgA7UF41TmEVuOU0ImAWwfZUc69Uf0rRKRED8ZaD72nnZLVxNSj
ui4oCYdydkhEJd4IKJtBYQTbAFLTWXqFl9g3HTEWwsu1bboRd58DtQeAEZpCfqjCEa81h/7xSWzq
RI6vaXO86RLjNmD8B9VY3/BjyDqUm/xZtaVCGL39ndwiYGcVXVrR95aZzMbMAQpKuBftJDkF22wP
vBcxBKsd4htzO5Oj6qj1YYQLZ3//2EzMZsxbCBHvNtggAh9TsbHJDRT61JcKoWRi4Bv0KVfJ2ecW
EvF+hFvtvcSlmKcCXdwxHdDTMAliw8ZEb2TyU4Fm/EjjvdlUoaNlx8tIMj3X7GrR99F/Jmw5IMOH
YKXN1G95Nqttat1SsWLGghe6ogwJiGC2Oo0yrGl+OT06HIlR1hsNsfwYhq1mx2ZSkm7OAk2xV3eZ
SOdpBd91E9Sd8atAf9IhA0gW/mOlbPkoUpgzZw0IaWNYDMQUQN+KNOUhotGVmvNjl5Tg5PHvEOjk
vn8pgCE+NWOGpy3rTmQJd+s0nFj3q+6AEVre8q2bl51q28+OL32ZrBstMZUIHkzoxf+jGOdwxwnc
naHNspR+/LspH7TNUP/u3gLrOE83tGk6uAT44jYBpPWnCj3QE64EUIZjfxglHSMU8eUoNR1QMGX5
6JpiFvVmBhuxz3qaoMI2bIs61hK3a7qc3AOBm9V358HNh1xbL5NlBm0kzHd8aF4PnDtWPeG9KVnW
x8XJ8TM0AqEqc3CCAPqoSjdO9KuBWsenQdtIVTvdRjl3j4L8c/Hvr0fsI9TR4lSlM02YgW0UL179
dEpAej5VEGsAai260ndB5F89aymtggcKC1SM2mKDdfoepzYO70kV1bKI5GnjcfUy4IlFbPhuzkOC
XJItQfnyR/6emluncIhLFROs//E8T9ND5Y/srkVauIU7l3Ll3JyqPfBcUlWVir0XQHDOBeyYFhqC
Hiwd7G7j3OSKP03YmT2YnwF6hDoUXwHAdUVq+xsU30prh8bjLJ/xAco+dEWN5FSYebGAyuhYllY+
ugMJTnRKeU/di3rfVoFmzHC5n/nL0e8N8Vq4IXw4fdszq8KOmwxgnfqupN34/fqfVWeG3XvxJgWB
fyMGkrMgQBi8ArI93iN49DG8oHgVqytJ/Y0nZUE2XMGAraIDuRJt58SSiMWAImd3BRwc2274ixeF
esHGK1G3Wwwrev845VTkbq54+C2hsD2LU6pHORDikNmThHQicm4ICENaVHBYF14SA0iAWV47V6CG
IcFxsHy/2qxj4vTbmczvcO31SIiI8wajIXSO7Ey6E31zpWlTPRJT48DsN1q6PHKVblmzaala3CT1
OqetnmVkwP+9xQrGAK+2WO4OQBrQ1FU2jaJ5HhGAGtiULuf0/ajT06DTCLfMfS3lWSvW5QiEmbp9
k2uWfm6uafsbTkSfS6wsMl1UKE59T2xy6BOXFeOTX1TcAipspTL5KjIBugyiZj9Uo2q8L/6TzBcW
SI71oFAcQdpmdJLOM1rU+tQCpuhd9jpyUvz2bwcEVJw0J7hHU4sCBR3UQvOZwlJxBsUIq3Dm7udT
DudZwQxZG/A1q1AkDeX/4iv/csDkrbgjskiaqjNWziFtAcIJ810A+TmujkzUO1z0iPj8xE0swrU4
5HVJ0SgpbruhXUeCUEqSFOyDpcR2B7s0BCcqEDaJdV3nbequTZ9g1n4X+Ld9gOmaPy0eewjigS8o
wHUzvgXN5Av2UIFnq6xr0rdu84HZjuXQ1P1Gw4kTxrHXMb/0B6ZUPm4eBmMogK8U1Os0Pr7+wh3l
u0Vz35XGkKfdRIeSZkBzQ/NHjBzqXdiKbYNQwYomFWIwANOs7AWcKdnmDhQ0xcmQPWqE4wBL6qYJ
4h+xs5MUy2TlnbApQNGHpjl2HrKQ0YmbMWPB6qentZ3RtwJG/ZBLYH4ZD7nK0lq+oXZzUERS043a
b36a4G5QqpjkpW4yHg4VFsCrSfm0oCYVJYZflozlcDEOVZcVivwYIwr83XJ4VnfzIazrsV6cfWdS
xsRR/5c+HeVBglrxL4s3LeyICiS56a9LH2JbXKqwVGc7yER+darNYI27AORR7wNTu12/Z2QpEKrI
uVKLtp9cfC3D574kqzjti8veSpe+v9+G/+I32Mp6bVEYUMkNFy5UK11CFoWmiVBSoilWbYRfeHQZ
SFUE/07YJ4pgDQAn+eXlv+kgksFTycBmzYgPWztyST8Ee7/jNWDXhyRnZDFdd81w7lWzOcY6ShEt
iUNEXYA7XepXqKhMLssG4NYtibXAcS+y14gMugt/2oOPZWtY8RHUQpQJq6QHIKGMLnMkQxAOl6Kl
JowiElcukBcHzRqh18s1BaUUE9f4Fdpnuiy179MwUmobfwxdOKJy2QbzJx/WhB6iijP+zJ8FcWYt
UcQkzFJn8l1nlnNyowoNE53ts5ekujgHWSdHU4P0g9v0jMEiugWII0jalhor3M3/JI1MATBJayYG
TMKmMxZy26r94BdBaqzdpIU0cgobkGjnSazXgtzBTV6PTg57nXqHEuwDz/oxgZoYeM2ORS1hiA7B
+qbLMxsL7ZctlxR2HvpYuSfAhX8Gt1Ynh6PkWNWSokc5zoCgT2xlrKZKgUYX0WpFWhqVBDcD6AN2
QmEQFofjPK+eKhdCoSCwZ/PIVLW8Iq+njegcxcqCuOAWvMpYsXEAvC+mBWb+zLV+A4MlEUEW9ZMl
wpvuaQ/HlEC0eUagHLbL1pLgSaFgyyqmT+aWTD4N0y8V6XnYIT/2HspLd6zTp1HRuc13rCxFl7W1
BfASBbSV23JQ0aFt8ovC6bx3iq+4QKD88bs3PPXgtDYR0PCtylleKl+MSlljwdPXTSh1r4puv8iQ
jUAqZvBPBXhQ8NRto54HtUFRsYpd3W1R9p8HLh4O+Zuwt4Z0Ec//u8u0wjXt97D8wfgE2uxj0QXb
g6e18pw7AXFOZ6gX6gVUh5jLSs4ByDUdoTDC9sc1o5lcWAq7Ccpy+LwW7oD3Z8w8y34klC3NwKXX
9q62O8ZyA7jfjlaz7VnhhOOyxYQAdTmgcduJGetuK2N8tJACRI8hXU4z4Wu6kCUteC12fVzAuouX
0YrzVGfmnHbjl2P09JcP6zLj2eDQYbzi/DDSUUyHysTzFACs9sPAy6fMnENjswrOhSIz4PbXJEg3
dXjCCdWPXxYSQJf6qPQVswfaAveC54ZOlj1YFQcjHU2i+xDLzJjJkovt0EmOk61gMcwAFIqa84Do
5LU9GdVznNsuIAux5Ha98MSGUsqBPCu8OI2biOWL6fbtc+Go7XuUYC1pXd7TyoTMGuGg9YsvtDVZ
J7LctHiOUzR1aotSL1dBWWr24tOjIvq85OYpaNcsG62K/7DIfxMhUZTj1T0ccbkfRTg2SihiZ5Cb
lIim+0mNsR5E2ZVxwIKRgByLjkP26JbBcXpoSeVnt8Trl3HNMCCddTXjbDegDP1JA7X7Xx8VrOxO
EMc8iL44Kj4JiLarYtkrHg34RqBzUUJCrkEDp/E3BI4MXCb2lnhRkvvljppfuoUnRdSg/HPUiY7w
uEJFIduzL7rQpn1v1aZyXRA7LheqTkPFILrXB1TiqTuvyBiLWoRQ/cUpVcJWvtID/vTy3Ea4E5TA
esJU7VJ/RNPTVGiwp809Yyhmj5Cagxlt5ReojBVURamSvbllpQ5tlKnAg9vE01SBkViiyLhsOrzT
k9fWg96iwHD1E/ukql0N0Hqk93oZq7Lynv+oDrYyQPvsBT5JEQE9gTL2Jda4wumJoA0Ml9u1pWZn
VezYTH2WD6jdWvYqhno1pa3RRtcLBnzrIpC86Cu+KsAeLXdbeuwIvh0o2+4coRsYWzLCoFCC9evF
mePj+YXLsav4d1aJX2GU7SMO2GcdYQ+8HSvK+YuM9xRc97lOCsWakJahtI3NV2SeyPC9bh+xDUCR
nFCy+AI9JgarG1GAPaOvRVTc84F5emeik3mzR9qHAImJSl35Ju2K1wj51X3CLpNvkNLmR/QiC2sB
4u1l5M86eDs1O6jQZvyJDfse5Pr/K5vnBij7jiRDaig3Q2Mt9WrnOU4D6BIrzQ4vRUzWrpmdPjFK
NMy+H07RuwZXpV2auKvPSI56LJVP6q2LG5wfr17EkVEUzEY+N6INx9Qyxdc2R7vhwvgbCleDQ0+f
vfMKJUs7etSoGqNPtZTW87VpcY7WRPKBbagqy0WxuW8Pw4Zhm+OmLsftYS+FXZc6JPvG202pfDnX
cWFXiokuvpj222owQi0fLi3CyE8MD+FWaJUGVpDWCVJQOYUZmievJXBNYPy6llcwH2Aw7VK30eyn
a7/uky7n4uTAQfnmDlBtvguziXuHuSzRDYhNq5sZzEBFV5/OAlKGRkM7UTKed1+gyHo052lRKvBF
WK+Cu4kHSSp48xU8bQcXOgCQo9BRBRJCY9kf5rMW/Bz+tOCAp9MXxrcx+E9nzQ5av/02ica1mpgx
O8wKBJGvhrSp5bbUeRIgGkaTdL9AdDNSSHXp3oVT6A7RQaJ30ojQWr065ostw9eJjm9eDR4INtTd
6Idoogz1T1Qogup5oHnahRK2njwox0KYcKfxw/WHPAm+/NVG8NJYWIygt7IH1QLTmtfoMeJWBuzX
7z/t819ozahP5eYtHo6G6YDyHECtUyWCGgwuylpBCwuTkpcSENAa57eqg0znANiebmqq4+0uU74C
uSMAZWRyC1xI7ZWMQGoNSxLuhVlcBKyjWBI2IAgUQkGany2yhyVYFA6exledhyfZcUKS3VJ0vDfJ
e3RSoCio/SLvO3V16Bo6e77p7/A+GfHADsjBvmXFqlt6OkSW+/C+ovzkRbkC6bxbKekBgguSwTED
bZ+yRTn8D7HUt5duy1da3+t0DQemAMSqHObK1njqkBFPBhaYE6LhXaCwf++NYyJeIWieor3RFobM
eh0vOCTcN10mY8TpPWrM3wgBmVEyAmGZZS2BDExdQEO/DKBzyHMqasrEUuUmPUZtkkHlrsMCzH+M
wo3QQSaShiNv9mj3JeecuylO+RrCt8ZDCBJWMWm0H3+G7T0tQTxVVEEvM6PYsd+Ny8KqNXl4kMke
WsSw5XrstLX6sd2frNp/yTRa/9pHbbWp5hWTFxNgOHBMHN3lNBEaOKacf1vebCPcRf0+Lt/kOj6H
9K9ckw8Jud6HDJFI4CoeWobfmW8HwzHW9fQz/yXfNwmAc48Vc67/7oyHb7za9flSlKOBQMK3mB17
xLz/rjqX+dwuRLzT5GuBlcAu4cEZycyRMoLVyeS5yzAwVCE+yaCcvznEvNHn34ZxmA3GikddmSkM
za2oxtMw46bRSAODq4JsDDxX1K4Xv7xz3/mdLNDw4DviF65oFMC2682SDARt+ImDejGSe/TLzfnI
yv6E27tjAVgwDdNNDbSSr05gK9QcgBL8yq3PHwYtq1QZhqjQKcBPgaLSpdCRNsCtGP9ODbToBpAr
9u3s+QcYNg6zx+l3MAkfI14cKwRXu2uAAo9Ftozn5w1xJO0WewMd50bSq6gtKWT81AzlmsSdZXqL
XLZJVp5pAISA/rvCkUl2o50099jiSsO8UdaT531dTiw5+0Bsy03cXp2WG6N4CCHdCPaGuMC/B20x
FzxyBsHh3gjp6vKwrS+Mt7EfzCePGWlDQfLsg5n52bjrL4aDyTvTwM1WNpWzOq9UmkdTCg2GR+cB
hm2syBgulH2bX7a7us2w8TyRNozTwOdNhigvDFf4ScS1ju+zZmZUIZQye0l47STQLTuMkhlrvdZL
LRmASkxwS54q59E2PRlTOJ2+JUTLxt0rBk4s84sZH1bHQRmZ6AVnK7WSieiQW5G58TRkDC4pg8+6
No6KmtGFJDElxvOi8KlNKdyKDi4PBXOPUZccY4geF3TxKuMXtG111vvFV+axheANHjUAZjWbDupX
Rr9K/brhx+sHY1A/8vTwu3UjuUSAUd1je/BhaJZXKroxTuEKMiD3HoEtHQKUDL4ZkTUBVMnTR3eg
Il6iEyxeV+KZNJ723hMw4NHO1gvIkV4aQ0M1IE5rWuUYQifk5kEvYvNB/SCwbzhknk6fnUtVJDGV
GCFrMa7egSw+GUdk/63h2Ud8wy5bIfvpQWwfUThpU9l+X9/nsKyF7eBTL19KVFM0ydWP6UJk+vAc
q3bZi3SbNyRnpSxTK3w+QuMGCGGiSWXu8FEUARgddkKVsDi9gpDAB8NKFFzfGV/byRFrW1KgqFcA
nHQL7RpDdOJSzHqglbSz2gdy9NyU0Paf6ldUiAtzA/SoHdm2nD0T2VQ4OOsNyH5fmdUGcKFn5/sN
10d82ZdfuM3ssN1bTM4Gy9d/7KgGviTD7DBHOiB8oTZ3SDLLypfvcSLs5DQm/h3/lU86YnYiONls
C41lQNLjz+CG+YskOE4WT7DTy0tLbFwU19sSB9easS+BFL7UMSEeW24S4ccX3vXMwY0mf1nmcTxK
mTab+o85MdblyORAd5fjswWxsDmBOaO76sCpyRC/RFtXo0PLOQso5Tr8zAiQKVSSThQQBz8O0NMv
DIKvhMXETOI6Ni6TentggLBW1Bf+IyHVDbyt/pULwGj+DINg4mL9lj9uTtPh1vaNuHmIVTE4X1qM
R6h/g9Zq0YQ5+H4XTZJtsKnpg9Eo+n3DUE4GiSC5XZ+NczKEcFtCEZ2VNKyxu29mjGviXsTs1Urb
/yx6gUqsCopvYfhL9OESOXdhmdN8UEaIN2ibo6W5K9UcWx0urrWSKyGi7ow5jlceiilw89jz9UNI
Jd8i4RUEVz1lygOyXOF7TtCRP0AVSkUUGXvf8mLxKNwI9luJ6YblkT9Mpkm/eDwH0ov7w5sl9WFp
a2z6Qr5eEQKyIvpn+n14P4/TdonXHdeTHVMA0IBytAKA+osPVrAbjMZUKo15qPhOLQPWdiJPboZv
WgwcxbbC5rI8Fx6f7G9Eyd3qOAaDttvmf86ox15CBtDnlT1mzjWMDO5/aZrIZYAKFpH+cGhyySOS
n/o9WojOQSWrq208Cx6i0Z4MeDbbhURoZYA62h9KmT7HRi6oDj3KdMuaUcxRYqRJTXz6EbUFGf8x
DAoeWjqqJN74aj1lTMPKbObPXi9V2JJiK/K01xHU+XAqHu1/3MLc+rT6gfVU5XsGpo75vjn2C4lz
WA7fEyb8eZqNAsX/DeUPEeC1FPUQLIhPGEHk/lwHDWUjMamRarmjsUGjALzu5PVT0RMjkmKh867o
AkxEiLz1tzRvJrUarvtlHS3NCUO07ZsYb/Bonl+tFKSd0Ry6uV/RP4mnWdJyrMKtOb3xJbeOIZLP
xf2l4f15g5HnGk+lynvXh+0fqkVpccRFBv/LOcUWMbdG4fqJpmLe8XlAvK0Q9LZ2UDvZfMJTJFoL
sFnNN0ZO2Q0wNoldkx8uG3atK489ACFRl2b2dvaEvAKG1F3ReK3anego4ZaxGcBv4ki/1gMB5DkV
6rUgviYhH6CIbrAaamZgYXqnU9IIxbuhvwzDrmAqCRYUfipWYkuraZtYMG7fYSid3JqJCcljFFam
BTxwzRcCgKhlnjhK+82mbkov2UfssjEMzllGqDh9q9zb8kY8OQks+4/1R+Ktlnq6m6uDJluAtBr/
O1ycgnnbcEg02qlaW2nqmdN+ZwrZxI5Vz//4wDPGqWKNqiYy0982B4OMWUJXsS0i7AJOFJOzY+54
iD1goCTwZVQBru7qEwoXqfNS/iySwFr1wTp4MCT0cGUfHA7WNmSvbsOO/BRAlvcR0rv6fGrwYkxF
vgqcDlmn76wvuTujFAKKazu+34iB7ux5JRfZItfy+V0oJ6Q+eGoSMMvEnRqAoT8sR9zs84UukV7x
L2xBo4COPInW5ZHR60YXhxbDn15zdzFnCc4rafMRl4LWEd0zN4/gYVI+0Sam3S1npLxG967rRw58
mkYq9xcpy5fkYZ+v4PB6ejomkf6e/LYDTOe0dadGTyo4O8WYIwmWCSbNEtxfHQUoI84eT1EMRjc9
gYJTvrDaflrUO9POCY9Z2Bo3Xfl+mjCnMnhQeDSOD1/1BFaxMPAa0k2KywjxolYHQRlzCQVUBfyd
yWxyWlcyn4ub0bTaJnMj3ANDQRDMHUPxO2Zb/Wi8y6mES1kmaAaH0xAZ6DLu3YKNYwCBJWM8y/fQ
NAVsVR7wi3pNyvHdUg/ynq+/ipDAsWTLlGGNE36jqFvgt+g3HKcnXd84IDAxPARBMWMu3zrxuy6A
u4YoPauRZU86UVOiBVs9y1ahskaYqzPIxct4fx2rKzBUQiV3GWqb8vZetQv9dfRDE5QpJy4Hd5wa
noUWeKPYzonQ9CaDkbxgCTO7jTzcFFAdceVPBZYxfA6ebKfRWRITvgOeuzkWMMTVTbGRSEQqfHj9
otRIjSLDWYqBlcD4o/TQF9uRa5P2AmltZU0rbCqMPBHxnXv+K1auxJVQYB1uAsTK2FAtWfg1Ec66
k7tG+44QgQ0SJTQkmglPKxvNMh7GP103jOs/mwUb8N9/zV+KKn2U/GqBW+aPrjh7SaSSELaeZcuW
fNEbPadHmvhWvT4/Nw3uPdQIkQSASUNyb77ZFOAsu/wO/64wJUAqfTpAEhnDNni20ajJiTRbirvF
ItsegTA8PUFrffD3xqIWFIfO/9imyEgJhZVfdOD+VA1uEfaPDhvP92drcIJxrqL/f+2CpoxIBa1D
n1oia7iFhXPrG2BTtPvTcWJiNB2c8Oo4Dtl4ITaO1C5nbzWK8Y2LBTWKfE4sTemilPlgO9vgXO7o
hzvplcMgqhBfssmOgAGaN5d+kGyAtFzYkETP8rjWQ5ZDMgoS9m5i+dXwEIwxsAVN1qbo6RD3eTKZ
qC/pdxKki0RzNND/h+OTw+x+jccHoA6w88kVjAK9wszmuG23vj/E7u4iPvRkC5s16sbAHtjOny5G
EzhZJNyMkxSWjIkUTel9QmWxcn57bwN4KGetABhXCLNYaZD/zSmVC/35+TcL0fRlw2MwMGt4am46
ejGN2vI4MAtfiBM+Ml9LO5aJ7dQQeNQ0BkWeQ3bERkI4TAf/dDC1KQqziUeFCTvMJxCxUDR+dEDO
bhFBBRCirCk8TdaF7R/HjMaS5H5pWDTYTye9qt0ijHyOCLFiO6C4pHvGIkTVmTJlqweNeXSoF5Hu
h8Ik4S9MBgrky0i8gipIG1lOYezSH1KDq9f8cxcOhNw1C9lXNxnNSNTv1eYDzB2LBa+DVXGThn4f
pfIVeS7DUzhDr3jX5WGR5EVKw+ZFhYGuQ6psq/1JOdUnXpN+9X/v/H+karlaUk/AgYRTeHdomL/c
F92RRRrubNO450XITEOAsI3zfMrWvH8uMUgSAx6AYZ0+ToLIqvTJ2kzPVw13o4A/cofisUm+54Ob
7rifRn36h6ESGW9euf4czAQZ0RFgY1AU9qYEcu9pLQ8i1Wa/9uispfKEjtw96nGjSA0zusxDbJmw
rU2l7Tydm6ZHPfxX2lMYNAdYLpnwlQj6Bj34My5MxzaXoDoNpxcJdad+HZ3C32W+zKjOVXboKkw2
vrSRvwLFfOepzq3URdTldfigelWV2fF5j2jbV3poDx0aezoTAAzfvMC6bE7Arb3t0exRFvITDai0
ZEp48HQoCEU9vx53ukPTEJqWkRwzLOYHdN8u3uQ4kEkb2pXWIPvUHJW94aTqFh+bmTZg77v6Kbe+
WnA2SWx0oLl0/czjTORfuZradJnVuDjEERo9xLjcOcu13820CoRaFhjZiFEDELtb+Q48FV7igQia
2A3rNKjsidqAUZxkvAWCrIKiPKSF+wKgYpDeYADgThvUmZT6wfSbTJosztZywIbnGENrC0hfUqSJ
tSBHLRJWNKbgpms6qd34GCvbXt4nmp3BuFS+ARkCfWbuFWly+TrHnr43mEVzmIrOrroYGFhMu2j1
dluW24DsUJuUAjZvNsY9ZXNclRYKFYS8QUnJg2Ski4ShzdtpMtGDF09Zet1pL3BWgcpL/6EynOTz
HNSGWXhwt60q84wsV+VpVPZTVB8afN5Yj65S0wZLG72RuTB7NWPgH0CosiaPyRZfEV5b3QBFEgC/
W7n94yA1I/StTS2K8IFjHxp1Y216NL0UGSRzQC750K/HJm88hOmJMUpW0W1zOq+JhYLmvPNRwE5c
gJgZKa8hkazgyMf6lmT6FMGVkWjrDtG3bA3ZRp6n9KbYPUHJfZqfuF8Yv0UKlRGxrkdKA6AMIg9i
mFKyraH3OFgQgJ97+pravi+fcIfyjLgZ5EpsaYkerRcVRpnoPlRtHSS1VkuRU7I2r56phHg5t0Rp
vH6GgOTk70xdRQaq6AK1N1HZkUa/5hrKcuKKrFmx8Fp2y++qXzPiXVwmflkoGolez0pOyHaE6Ae7
/Cvkb1lmRg6615OSlsO3CEnIRkj3a9xJXuJn/lKwwYxSE4nUkxbEnzgPZLqCEXLWA0/DsyLTfwmi
mK0ed2YEQ+ZDSV/m/RCiz9ldoOLlo6Qsejmkzi0OVT72bHW/s+ga2KoNh9mDGjnQyX0X9TXu9uus
Rt0+PhazAnxXbWDueFoQJ6XgViHhnQLOmQpbBCfbuA7wi4t+ZOUjmrJelhpc2FQyNZEnfsPNieSS
MmEhn79eQtA7erQpFebK4FjzmKo38XZEiUUBUj8exlEgBOOLaDX6DIXb0cn5KgX9lMnLhFy9n/R3
NLi+ddgOF4q/sltu/bqeRr9a6tkC2rrpHHAl7FeuyoX42OhM7tKwr5kITkWXS3/kyaJrj62TUlKS
9D9PxfIV1Z71KjSVUg3kmvlt6fiOcInbnHLJRE7MzpmDcKA4bO0xuAOICltb+MxD8VBYjoUTzN/W
b0WlUP0H7CG0R82ummnc2N9e2LBtZ0Z/tEWIg2vbPl0ormkq7KDHUPjawDsDw1hcE0qFGNICymCV
ZalnZKfYVV2KzDZ4vYgwpiOyEpCD6qNyVbWw4W2T0KsTvLqzQ7WZ4TP8VlveBQLb1UQIQ8puF2L0
lj55HLfb2BKxSnyOvwYr36+e16/VBLFEZ4xQPN2m4Tn2pA5uxb7CW2+TLZ4qoGEI//HoVUCR13eN
3KpUq/IDpYzhwz5RnpU88o/ivofYGmbYzAGw1GzD3AyzZ3qD5MyOLYKyYX/df3StoGcFzZSEsok6
CPawIQKtopGxPGTHlQ5EwVUBauTwl/zlkWLjd8xhdr4AsjJt2DB46nPebnTgs6DRQis4cYBDCeC8
Pk33ewIGUKYrWh8mAFLEkfezN/g7DK2qu60PjbM3rdd6AmTn+5VtIt7a34eyFyVVufh+xBORgbJw
5xzUupmUuYmHLScRU1r5fPKWArbQPEIsyFqchFI7Qx3sBQQe3VKDFUinJBBsTrr/XZyTPZg+oXcV
Bs33VrNEgczNs6Gd5xcjLrOXB0CQNR2dZ7rdhR6Y2LdArnvuD76WXQ61elkiaTpF4uX/USVBevXR
60+P6IOgx9WBrmrgdhgE8k4ej85lMAAZHtVoaihVHAYgwPqoVp4HgRlgnl3B5zvQQDeRxKOuKtzx
g+3vxAJ7V13lzm75l2Xq3k3HqDt22ejpbMH9Dh97xVn7cgQp1s1LRHHtM+VajrRS3EmIMUn2z1Oj
0KeylvMjD4lYvyDfd7UppIABhTJBeQNnG5gtchc7gRZRX7TUfEbDr8FhP4Vv826VOREL67RXN2S0
P8vPuL+tV7rO/QKaRHKPvEF/kfEit0WHBmGJDpiWt3wtmnOaR/JNl5ZYtUB4IBRbJr44clrhAWHu
0A0GMrqD1LwBH+fYQwlsV4vE6Pguf+5IP78mVCkDBP/I1OufrYfGa0wLQilFCoJWFIdENqaoxBh/
foQWLZcbbLVRSHcM+F/EIoFQAmjhH5VGImRznT6PTNBbrGmWa1nBcHkkqHZmDfAnAdIPE07Rn3oN
AzEMf8MUOaFe8t87rCP74zXCdcqLGXUVIqhVmNklTnH7RnoUMefpv+4U5CPwPmQ7jPfym58CZ8jT
yIjV8ClmNiigfl3uPtkz2KtgcCsNHG4kHVfnYrYpaC8N9SIkPt2lZtvYIYrrR8rs8F/FO8FYiJzn
r+JiY5sfuGc9jmMup42GWHUgBfIPxkmxT7SYrt171/eom+1ZcI9SdFgS0Z9DDukSfng4TDex8Q2i
oi2N08gJGSj7eJWlF7iaPzZ9C1NAxWJM1c0roGgkMG+vcweuo5QwR6xSLeN+ktuZG/zPio7jnHgZ
/9m3K3/yICRVRhqWgXWzir0JXPx6tsOPKMuxfvKc94FMnZMJyD+8n5Dmr+ShmjX8Sm74ZJNn3+nq
QT/h7na8ViWaPZ8V4A4FnGtqoYnM74S+oGTXQby5N46OSHLuiksI5YerxZL/2QWUNtvjH+1wHyuO
Dvopj4/aey1rrx8MM0oVYRXbrYg4A+px6DmTolu9P6Ijd6tWNuUKKLaVW0MDw/3ENkg5Gs1lsU0p
+6DohZVtk6y7V2NerjG4TOe8j4ulE7Yh73yMH6hvlmRaGn6vcrGjhdFmQsqJZztoJEYzvoaxzTfV
Cjk8u/1W6oEdG/f1M+cABA5PXTfY4iIrDdbkjhMrEGYnLqc0hJjOIXs4Qzit23Ru7Ak9Bwh7lTsh
aAlLwEcWnqJv7BSl23pn+O1BDZpiNnBmjtuiQSMr3AOHYHIM2/cBkxH6WkiAGp/hiiqlMFN6h9UE
Ns1Anoc81bqTFI6NKHse8aPfXzFfHYbshPpKLDA8yM9H5UUa1i6dPqVKPUxsAV7MmEKxO+bILPji
00aQbiRy10PGJshJG7UTtgRAkkb0XT2/R5CXStDrkZ+VvA2pn3yhuusNX4mHM7mLOD/bQ92KQx4W
0SqLGyc4y3SsBaJngvup8L+N2Rl+X0a5tN0mClqJX+RmoSqEP8si2kPDMa0eboyuLoC+yqYhoRR4
hRjxU6Gml7juoGo/TK9c5BZHAdYb4ogeOFvOl3ujA6JcXT1MvgK6N88Ote15g2IyzRddUnZMbpk5
QRssUzRzGuFppvIXr+E+0NKORIIsbX5mkdoAesWD8IVqr/1c30zLv24+C8ESbAAim+x0JgkJ6Uq1
oB51kQJQla9aOSFZDT2BVViCpi7cv8U/0SLsfn9JZDI35PN/qgcXtdKkogaHV2zYVA8NheQmcMyO
UqlzofisrVl5PcpwhhUQMM4PZahFETIq1khZWHN0C4Ss/AI84N5ddQgr9zhGNxeMGfwcqGlmQGTm
wlXmwaD8I/ucXy1/FIKzkrUwuh1Wgma1sLAC1YNHVvZU0iBMUHULCfB/mlBv1FWRFEKct0Eaq6IT
vvouYaFKgpI/0sYwhh5LFmVnaBQdi9vNsk3g7LI/QxzwLCr2xFu6WBGv0mOa3YYrllyotEX32dfW
5lqXmHAtzmyixhqtfANoO2oz9GJIuqiL6Vb5IIO7OI7rbwK8HzPs3gojnb86bZ4wrLrPSG6F+Fyd
G3RINEsSWqNEreyJO6tNNjBJ11Pk7G5AJE7EulBQ2jGQTutwQxlnJU56PtqC0ff7zcQcYdrnhS5K
XwYh94xRYNrYXihMtd8SXcxjyq7NeGlqmx1klTT5189yUhKouYeVS3bD1sU0vE6TuwQSJrSgOUll
5eh6v1ox2biQ8+yWqw5iFbiN8vJcgY5UxxB1oBOzLuG9HIOeEE9WWPYGhqkam+jOTQmiX3kBGgpz
q2mbmrCa7PgqCjySCTGniVhOahKzDUPAJ89zXMhwuDuJQ0ICv3opY18dKAc7DEN4i8dO+k0RJP3Y
YGjW+MDxpstR/pRXM0NXccLvPfwkDxiAwunY7TB90d+5/upVs2QKDoge5gDHcG1GbJqqhz8chc9F
8/L5644Vw5F83DINiFcEa4jKkBtXQPHb1g82b3/7onNpnviPsWvdnW14cRA/8abF+hkKLdSKnigk
0YTXnZvm4fGjfIQ17y1+Kc1ZjrOKUmFDPoxv94jW/8aLBs2tcmlZGEPN+Kztv7AJgUqb50K/lJG/
hCBrDEKMw30euiBNIxbJhOf6DNKYNbX4E4PBjF5fjEILzC5d/uFmMIdjWxoPWvxXnnoqJVV60OUR
lxzjs9Jecwjgii53TTooXn36otdW2jTgJ03dxdyXGqDBETlJlKdKgjMDbOMApYK6R9L/B5e5nzhw
M05mctWHyNwegFzxMtclGfV2Wr4JaXbETBsRTlPdwTDxLsemEvsYXxhf36T5Uv96MrrBeqjdy+bh
G9vNT5PTTJIxd7JqOcbf2Tj4clhroiNQObYtGg6+HNJ/BV68corakHtVukgZujNHqzUE3KBFF8XS
/vkpAOFmC/oybZaz81xhAD6o83j4zMVQMCE4ARbnSWKI68IquHzDe2pxwJrRq1Klb7kZcADdk8AR
38jGdXhnYuKkKf4+31AKP8jcn0NgQHuUdRoUpzV78kxl6mfNMos/Fl73hsHIk0MsoWSLRDbJH6A9
k1vrQoHYrExC7dJrSInC3mAb9xlJXxAgtGqCSaN4qRi5C0hIRFh39d6nkTwo86GKL6WjdEJsgsLi
BcDP4Ikux7SEywyewEALfGUbc3kzuHFEImoLR0eT1wpdMcHPVtDmSA3+z44bZCNQllyCFOEgqfwG
zrTqnphiR2MrCKAkSDgqckUtBDf8CHkdk7N8x3S6+1fPOFjakZ9Qe8SW3kvDup2SWBA0aVtFEFOo
Hq60jFmuKlHPGB5b52wmp2uLLSWp8NIZy5hKkf25Z50ZbQUVhDNIUsYkT3AqWvRh/e0zvFawRnyY
Igsw/bC6uJejJ0spJzpMsoLzVglmNCWtCc0tpYSYQRRysas5+IZaMJhgnp/7ilW3MTXrdY/RywuR
2pkC5U9ORafnOytYgokmdT7SC1zZvwuzKKVfsrdHdwDzOoDarHkXbE3kWictK/RHMw/AD4Ye9LlO
5bg4a8AHXbn4hNT+UzeWwuzGQnKd4pmWHiAF+imA2g/QtXPkVThfXPTmQ6o6uy8WFX1+oofhXwd7
n5MxOPBjBGQ7Jm1MTzub8rMOMo76ZBgb3nPTU650vzFUANa9POgyWM6c3t14eAgAmc/0CK5UX0ye
9OJDdnULma4of4djDgyz8WzpKFPIFaXkhgsN7WEricNwoUV6h35Cbg/m9/yos6ahZPNM4e0GR071
Mj3A4wu+f4PXbgRYse8/XnlfMDKOm/pkXO14JwhszIUG+ZndZ9XJkZyM8yntsssXRq9Q5w5D8vnN
Xmqmkn6tPjXJvnRzZWyVn4o0nqreX7Yrd0daLfrbKNhLdPD1RdP32AB7JEVxdgCOM7bIn+Uv5hHH
DjwxjDye/c14AS2fqke2+EhLl/Hi8mw7aeqm5g5ZPl8Hiyp8/oyiqCLJrRwFqOygN7C75txgZHHZ
XQwEcnH4T9XkxWsBtOfkebjpDCREYjUCDxQGx9XqqHDLBe3mHzNGlcy9RNtveTKetLUrrM/g9FpU
cgLXlgr56PdBv6x03ZO5VNtbtBx4xSi1EovxoTg/oBU55kGAQACYG5zleLDti5CRLiUUW1DfxW0o
5Ww64wzNEtiqb5k8nCzU3Wzfi1IUZGh/0Hl7nIozuiDpEZmk+xz5LzSoy7PirzVsU3lQb8Lxt0IH
uFKaC1JUAwP2IA6muuz+Rsx0ql3Wy5pNfEEDvO3Cz2QDtIVrW9dyFtgVvh+MCrSaagjxQQCZye+k
TFPfz5b9NqjWTOPt7/c4L00YrlXvL1jQP8onV0mzSRsBGQDtj7Celx8k8sNCNy5nrqMwFxx374ja
IxY29ytvgEtuBSJ8RSBEz/hOTPR5yffZU6Gqcm1KdaDasuz3PKKZhf/ORu6TY6LR9HCv+KFAgu0h
4erL/6+cmKEkLSEMmLiy4DJq1UcGJMtwFiDh5LfUTi+YBJ15SU26cIEueozZPXyOpThHxynH7kYb
pvOnhMuTOFp2YPYltAfqhHn/7aUy2zGIjThgq5msKIIbJXinl/lmIYYLhUePmy7ZlWbFNWfTZxEo
JTDif8VG8CT2+XMXNs21um4r7qXLj4yBPSpmM1rYBlKAnGHpcNnFl+gBHG8c5nb/0KRl+Nvkd8zz
4+qPyVFIVB+LF6TDD9UZKCqM39wXsdaIqqN8lKVc/DjZ+NgiBwNxgwQiLSks9EqxycPpL9VU9g5v
GtPjMAaDd3FxHbNySXPsTyAF4FLIcM9TJNB1FAneQuU6oomO3oeNlg5sLBE3e5blSIgAZpIUtuJm
pJhIERzqs+xjz5tro+N0nDRSNJ/QhkxvkPxog3oc8GxiQBEqKF6n/G/XcR+h49unovc2bC/hnS5X
HowK7rxnDxEM0lOdB4D0G2+UGHCo28WGP/OuE+ZrIR9BBU2zPck7GvxgZ1x2KF+E5L7ZP9jQ5aWv
80aM0noApWT4ZvjAeAqH5rp2gJPvjTha8UajOkMQ+dB9Tse6FAFEyT/MlrHACd5qcqQXZ95B0Etc
HkHKuGtDTo2Nh7bdmzOCpEJGM44oHZpRoI1UeI+1tvv1CrBjbVLNrGcN2PsjpTQG39mVsjL6KlYu
RiXlSVNrTGaaJG4vphevMPtigp1SFqd6iuv+S6spQD6hya1TpzsduZvrTr43T+LehT1k5CC2xnqe
nBLiZ1JFVzES+iUs9mtYo7rfmyb21QnWiSB9xG8=
`protect end_protected
