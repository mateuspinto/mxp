`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11136)
`protect data_block
N1sTHS3Mz8XGSWBxGWi8gnXRXNX65qK6Gjf8/XRHLHNhl59+WbjLBkHztaQLDIbDvrhSu13iwJFU
D2lN1g8x3XsDxOfP1dsMAxa8BT781wM+ECBA7nlgqLbP5kM0v8SY3sQkpY7rzAe6tVLQV79XA8cZ
MEJpyN59xc0p5tyJydd0SMLwDDSdT9dWQQ2CfTyot0ogiEPW3B1tzAScQmx934Eq7SSDHha5Qr1v
gUpnrvwxVWMnGsUuUPMSw1kNCGBzNnxNl03ANiOyofmxegNtyXQ+/+sZq7BJ2SB6c50JmBNsCjtV
1np0G2wzpl/5QFh19wNEXqkBkrmQjjO9pyTDMvSx4C9OiOkwtP+m5zLkX+U1RkXtT/MVyITsZOt5
Hex5RPp5nuA8Qar0cvoESMtyQ6t71v6ehQEf6UBxpEt3XVIQxWORY/Qh7FFeazpYGW35vJHS4jW6
F9x7blZIgH+hnnwFrZ/xT/tkrhF4z+9yz04CgfR/F2qkpLXaJuOhXCFI0qqQwgx60Icrzl/Ks8vK
UP91WPHVWHW8cXKMHwWwDFl+Joiuf4Q5jFezU9B1g+BBTgEhK/SNen0OKjwguS/npUO3Pry5Djp+
Xu0NFMjuxUkTpLjII4r/i2Fu3AFKn0vUPFs3mOhQp4jmS4Zs9ggbQ+mNc7V3OkgWLj9zluvsYAg2
WK2ANnzSPgxX+qHEvIigrWR8TgdQIP9B7Ya6qllcbbovwqBDXKE8k7LEp32Yt83j7rEYCDH0aP7v
1WacJIOpV8JGp3b18lkcEM28ekgqqeq5jo7ujHIyOnBR3vyW18IK/owJ00XSvDaov8WEpCLFnnE1
8ASJq9RIshSFk7zzjvHp5yimESbZtT6wfurMynJFAHwC2KNAlyVcpm5082FHHVcqupWOh3s3wrJT
xIakDePQaw4B/IyJT7QO4ju+E0N9zstkyLrQ9hsm7reu9y0VV5rM+EEnqtLXyBfcyOymzoSYN+o+
1M8+nS43tVIOMdOOsSgKBX6VvcgTb7hpmeIqiFjS/x+CQ163RPVHGxyj/3y38B1sLDvNl9uWAwnZ
kGAzn7BIIBtUX035KDflyG/WF1pYQDEWdPeV8ndRwfBO5Tr0eaTJZPRZZ1RDR5RJKJMRw8Qe8ET7
BZNHtE59PEXpLW0+AUXDBfcwWaV1X9jtPCu3iDHqvjCvicc4vpkpCwSJVcGnvS6NlhgO3hcqwBIX
lhRdHishfzotjssuNfhQGsI5QsQ0N7Yrl2TGwbPSi71cBBWbhecdfJfYVgHdRb3OCxx2EhpyNEiD
JCIWxiE2ojWogFzUKXLs7aMsmdLET34tUvkEgQ1rs75dzQr2irxTJiLCigYuHx/yAZ6bIoRUY+S/
VmexV2iJeNNrcHBPr6kBxQq3AEfXVR44wWFck+c8ZZCd00WSox056Rz/4JLzIEYoPLXD3GURxbz8
OPYInesjkm/NlGiPQ0k8o1Z0wYdsnLxR0ln8c7ESgNowjaPk+FhIINmXGFGPb3s5r/x26O5zukLf
07ZZuWwaKtQyW9wWFOZaSVOwmLgdWXHPnqAJFwM9kI6UGPnB5hrSybLv42tz/9ru+KSlEjDRN7wf
kPaOgZDjwjvtaEcvXHZFYdhZglhfH/V9zXvk43TcSr3PjpxqmY4auV4ykIkGB3KC51mevESGEcKi
RI1HuzYoTsXnc45rKGx9MnrPK4r1KMVa/WBkkVazUq/ABpokJZZoho99294VlYdPxIxpJdSZf8KV
Vt94m6V1wSUgsOprTuhwU0mswb0nwzRaZCK1ImFvn7Iprjoic+a///3Bi3OaM7Cr27UaY3xGAaFD
iMzH2pFxNZu5BlulVfThLZFrBovT1FE6juZhQ27S07AGM+8sC0/c1moue5JhqmHLNLrtbXIBQsKg
aRM9SyWbb9+T0Oo5U5uOGfqWgdoUmynJXLy/NxPQnVbH3eBe+YQtGnnGINz+hL2k45RViagNKuZB
Off+/ALwBECuHODuJImQgF5WHbbCDonhaWVCAuHYLpatCSSXI55e27Mqo37jBtGsFZriv92L/CSA
rUmX9t2DWK905N3v/2U3AfsRHB+uOl6lAIHBiYWe0MdDuO94AIraxMwWiVZw6I+Whe2wAd2WNq7e
0358DwOvtlj3qm8smivFlkDZSc2J/vRchQK5NIBzYQZ2dQ2BwE8NytZQqC5fRFx68R3lcE2lXhaj
26rXMMsSd+9dTFHrEIV4XFAtbp6+CpDYbcLdDqzgMGGp5atXkjpQHDJNgS/MEOQWBuEfwnxjpWzK
CFydZzmZ9sXEMHjx27ypa2SzYU+Dnmgqv3hpGHa8M/KquEX8DaJQZiNVxt+x+jygCABs5JVD6voD
qx3oRxOAQ5nYmhDusag3fpy5flkGU3c4l7GXCGx/B1aKyrdilzhqA0dtxOsVtHI9ki+pGoT8Kgwz
uJ+/zdilKU8Xr5b0sIUVC4g+LhIUsjmPxPGFqSxVE0g0XoZdhmUXLNF+kIdM1w4BgCMlT1odsa+G
DRkYA3uNP0XNtgGYXpwpUZ4TihMdvJWoEMLMcxDl4YcsOmTJ//1yLUEdnXCImYGTfpakLzoeGc0k
g7vF47wxzMLxFGywd8ihvz3obq1H/JkuzGI1539suQXzL7W9qQ8VCPmN6b6DmkkxTHwATL5OuvU1
eE9d2X15KPE+c4Ko1/ijp9hOEePxSzNrteOce13ra5nmyb2LNoYfcZH7icQdB1TYSy1ZFQYOCe1b
WB4lsHBJXWaLo4UmUaI0qpUsd8IVzOgz2FIVFYPMTPqqyn72TDNqsptsNcNy6ItwFVV3U+soUbha
/gEMjLTRVbLwwRk3GGC8nQQtfQe7BITLmWpk3w0V8LHdh9Wv+whKMZUcXLapa71W1RpiCjk6zBXB
uouX+HzulEqDlZNvWJiMNNiNBhex12Tb40At9e+vtUhiEkmVj0CFyjHIcOBsURj5nEiZ2w9V4k+4
BObpmB+pxKMg+aNchhnsn4uWiQKpinkPtHzJWG+Ead7eokCnu7WRDavRoEbkqAxBaxaRLwxoA2Oo
44C+OT2CkpjzmtjQwu74zp0JLvKZwIQejKhaIoE1xkfOWIKkR2hH8W/PG25bPedXYiZGM9ppmFku
cRt8KROWAdWlcmfXbCh3bYjUtFNMViREv57MFutZ5vyQmiRgf1ihRKq3wX/VEDzkrR9cEVe7TAuu
JegcefyTPpT/S0pOAjQHqxXSsVfOB0dcAgOFuyiF2rkoy3KjrWxXEXuEIN+W6u/cLlL3F3Z6+IDu
fE8pFlXshTM6AW68eQf1YcQxvVGcdbr8DAx/G3Nre8TtFHWuXmXyIGF0PJ7Q5MUc4WEhpPPE9UrL
hYdjbCPHWBl60JaoFBB0vh5cofZM3qHls9q5pSmak6u54rFFsDpJ0vziSDogVbv54TnMLHDeEahT
3VPiSBT+Yq2DyGXeYsO4/C0NMFre6AX++92Tap9pGJbE63JZnh+3DlQdDCZKcE3kqq+MajLzXFBb
oPvWQfPCtlPSItGyYMGJ3/Ezo7vd0XP5xYhncKid1YKpwHLHghGmBqtOAakw47CYmLUVzgsafH6H
uZLWRhiIku+nt2YOn2bpf2avQ9mJ1KAtfEw/6GOjdzuzTb2MwBq1l2kP1nAuPP6Dos8hmXwmyNXG
NSfrzNKyy/g5BFQdh0sH6MVzeBIZ+yhjNMhBJ4PjBV+DXrUWsAp4F7um6INAERbIQoKCcyBjqijn
Thz2faC3b6gyYQXIE2DFwn9Me42/yILFIr8haca9rrOCBMrkh+QpiEE8rs6RjcKN0gvEiwSbnk0a
AJlxr7h+TfO8+vVk9INB2CL+vf5gS/jyZMZsjEGDURGgXhyzVxbq62WkQwyHfFamBJAJPjLA4SB6
JdDnvt/Ip4L+RoMwlKhk+sBBSsfMXWz5tQc3ZkCAKFPghsYvujI5bY3MRVxa7xJkEKAdA/2xafA6
oapJUQFkl2fGAZQhAzXG1xUIFzxiPMyxe2No7colpyysBwfOrDGG79pAODBxJkmtXdj0IPsAEzPF
x9cnetNrqjDSsv2THkYdsymfwAbE5H8KgTvL9jsnHzW79hEVYTa2VS1WPEzjZR/3mQdE1+j3PYlZ
lebA4m1Sxrquw4lsGc67c04n68AZBlvny1C74dRe8q8dgKjxo5BVN5VvHVJCAclhxLB2Y6VqtyOE
jecqvJSKK6ESAmBdbhk93maG5VlWADFOMf8Eo9a07t/SAo6/qBiVMAvNH/kjmyTlVe6X1VCO1+zX
WM3hFup3MikH4d5u5yyq6Z3GOlf3AZpVIkGLTpvGp4ARURlXjYQ/h4FAMHd/MDx/4TomTMDY+gkA
F+XCW3S7UARG6FL7C4RMUdoHXyKckqTCpGMQGglEQEiYL9yCXJEYsxas/Xr9GZ1z9xBN7KLjk3Vl
Xa58pTTTvgfiIIEQabJoQn4nlikUyvjIG1J8ZYGrmRf0oM65laWHuBfOmL8qocV8IqkPTdcJcm5R
FvBSDpTiI5KzReqCFALmTNzTVg9Y28pZhIe32iYTiuaiaT/2qvRonqNU42ltGTt6dOZPVHWECF3Q
AGzLaYwUyB2kZUAN87M84YQ/XspANvDzZxZKHT/dg4yqUnn1YEF9+y+qsDyKIwGsM52slyOPQ+my
r473kzGliIhQwZjannMgLlNIWSxJSiO/SS8ZJ5Oa/hLRAaPgD1mRja2l3iMoqULD+WOzikUHHB5y
EbdoXnh8g6WU+0xTwmGg2jmX1PGQEV6eyNImi7SEP+GlHJydWAru/sS94GiG0smwA4naVX/RV81b
s+WkeLmkgfLNPXN07c8qjLYYC+LYVR8LBQhWl7pZOJCJWUk6/ZEttD7/uOr+PmrzjhXHZnUELekj
Gd89q9N/i+jtYSpjqhvajzl/nVAdo6w466A2Aqnp/wrRdWDChxAUlKpB2eWuEgSUvrKUZhR81Tu8
HAHYqkTnxPvUq3cpHyIBpOpJy2lmFFAI6hC8vKkpYEoYMaqtBft32sS2KLr/cyJrnCSzg2q7Dxd9
scD2bEraTEd/B49XS07+zkqVa5lNHyFGGr/qKb2lV1ZzH8Nv+tDuUOXQg0hb82g0K1B4FJLnWfU1
yM7pFsJCNrr7YfJ1YP/C1IY+/x2Oz0ao9n/cS0gAINzBja/PsdIcP5xVwPoYt+cIsnDE97PdkBT9
ys434n/13hokpsbs7d6w1l8oLCq+bJ36QQik+ygC4CXin2FwFRdfFMxPy8CviGn1tC4qLOm43m3D
AfvekBkFJ7hbeBfbh27IY7PxYv2o4nZnGvuQBQU1CNxS2ZsvPmRUfC4N39sr1pk85B2cf5O61FM3
tjBxRRbkHYk+EQFwgi503T/o4NrpWcsCcPTahKWJDlbD5u1DFTKfgO2IwbVhauyiifjWDK/dheRA
eUEAhWKCx1CnIvJk/emdW84bbiTGQHSFlOFnAl5HnBnjMyIDVWQJ2pIey9Q5IaCBghBi9h7oeH3h
jYTM+9/lyRYw5Ai0h8Zf55zQJ58fAvv4tHldw2LkiCV4yK541MS90FjD5da/5jlaFmlyUgLvUv6F
5pshgntKEy4RW6x34RBTilkB/phDLGJwpe9jJMuWp/BwyC3F+i6Ntt3atyCc4egcAIBOwKlPw1uF
w73nXs3Z65BUMnxG24ta1JeGCkBlIw04rz5WXGoMZ9Sht71eTCqWD3CsPzJFfG9dzOD3HskSfA/P
oCKLpQ+U5mlwk3EMaTiwRGZdQMeJylJwMNjTtDHkKryyqlBwC5GPp3knvQXgf0RvLIlvWF1Zh6hU
8PxBFxX2QwMI89bz2btPNzVvvkGtxJq63753rinjRbq2SRskl17KgKvac8UXPKzYbzpseKBSqeVP
wNFti7SfzeU8SjLvKpcjfCMsXS6VjK1V9gUJeRNXACWJPjLAW5Rly2Qp059xCYqbH4SAp4vjc94/
mhNY8fj+P4DwIMh/VAkve0qr9yFvB6aJBpON26rCWk1BRjywhh5vIJgWywsdffVDHy4smX5Fun+z
R4VbcvD8ueBpvPaOWkABPuRo4Fdcc69xP7X8/u09asYxR03tYnex/+TozA6wFZaUejsR3iozQ05h
E1rYTKuthdv//XQQUe5mBLhAYAKuSdDNZUpEaGUS3xfVsYrklR1Rt4/dLw6wtuGI8FUmWuj85s7h
gt38+nFrxJZjcMQzk6SMdzW4KGx0KOFDoB3ovR/Z5iVrV/mogsmN+P1SQGbTLvzDgaEkSLRJosTL
zToKA27C2DAsp5Ft1a/mftDUb3ZC2dAbz1Dtpdy6M3rwUh+c6ltZV2mmMdNVVGMuRWIsXY2x/np9
+YsqBZTnfHJ5JZhTvagsYga0bWX1nqX6L3IfaBFoCNaLMiNcNtPUljRtmXnbV9qyidKwFuaPnmGo
yVlwqwhmuf+Jkb7+kJtJrgvPetXyGCbjPg/8gWSw05Knk0rpwUdPFEFDortGwV5FAB1g1ENOyyJD
kfCtmIsJmr4qpY0a4jhoavC0xHBeHC/aRAi5R5D64tIv1vNcf5oXTYyuwqcfyFS8psTnHGs8UAnU
tdMh3d1cEf69DQldHRqgyxdO8mu67dj39+qUcRAXsYPwVpDpPds1EAZOqjOZKjdLvpHjAeGnDGbY
UlCWVy+XwXGTKdl9oO8AjLHZAYuOv3N2yDArJUsRLLjlNu7Vj+IEMfsaAy8TkY/GYh4DHdlwxrCP
8Zs7uko/gJQ8au340AIDyqVw4T/acG6A/uH+WaniptHkDKy45pkAuAtq8Qt0YDkslt67SfTeWRHB
roXcTLeHXMPhuT31R/dP+9Fb6eKr8SWNh5ZphjBJ707CFcJoiqPGSpWd27i4hpySAZOPmeJFJE49
t43mb4JppmJN4Vj2xnRtBgAV6zTxyj+qiLO12VovVvaJflzAkSaOYLDcTlMoQ74EwqLuSQwv9yLI
1pptBfB1a7d9Gmx8RHEeMils4WS/ea+Sv8KhIAOjGPHFrs14yF8lgQ1RMuiO3oATM4dKT76OOAHu
J+A69kHVMnIWHjmgobs2Dksv4irnR2jrsEMjEDh9oG4abRHrVqJrADzhrPqLKK2HUmDlHPts0IVD
z/aHJCEiyajHllaUW5argcMHILkoJnSY47cOXdat16VNnIRRVt8h+wPNOjT/8xX9dyrPNODRBFXE
VAp/U5pKsqC84R76FayYeA2H4imAMWipt+HzMs/DrQ2q2zZpLuDZqdtmJGdIjnx3r9+iprFErR+2
VTqLokS37qh8aUK1f/uoDLtphW7wlxBaQEXwKvQ8YAc+3tDlFscQrPq5Gqq+jrIIk33Q1gwmfAH5
aRwg/PnAqXSVrla+ejPnRVdmB7T7PRM/ubDrotmVWOMzB+X/NDOzKD9uBGNbgBEP7NC/f8hcda2p
2Br5iKmZrUHMd1age+GeeGGoK7G4qTnINJdcx2ezim1XVFVUgEXQhqAFZBfoocDDOPvPS0xzPoHj
OI2A1Q6zU5B2t0x+VUuogF/xWc1jFBJPRgoZXBJyQR4eRGt/rytkAagztf+lgQxlqh2+dLJb7Dwb
+oyXN8fgfIUQ6RLYDG6k0TR62QaecL9fkJYjGDNvD/wm1L2cGWzw6uFFt86WV2Zeo5KxfZwbGsKN
+uE/tcDGaI9G9qBlyrmMF3yEJGKPQEPqfMM1VG9tb4ssxiVKPPFQOXz6ddkPvG5zdId4pql/BdtB
6fGxwy0jzrEe5/1+21aHkqzzMQFXIFtLC1gzsRwEbpgfd1q5PZbDTJ+IrkBcKbvYNvtFpCpbzmua
/jy+PzI/qjfDm6/zrVfH0BmY7xccsoCTkxyZJVS57doburdOR1uUihYdeNViKE25pPCZpIRA1ayq
wttXswMbcY8vXFVcKDhUQhDhHT2DnL3jW/Impc1ONv87Qc+1v7fLbzKHg2KqlB7asfGuX5XYNM+D
u2Y5kRmOlJ9WKrxhybnpTE7hr1vuAb8XsF7C2FVWylOg4/BmbOgyhdorE8AA2o86Akc4eS95DI40
ElViiDNWJoL1U096JpW3hMqSXmq9IG77q7uU5tX2D5P76cafZM0YIpu17veyZ8NKZmz8GE4KDHBq
UapJZwO45SW1HBxTfMjmiwrIpkXXPnhwNQUsEa9lDZB8AN4fZAWF0iAn0LErTxoimtu5kpU+lPe8
ClQXVRNOBgQq5OsEKjh3Mrha7JMoPpfdPGAayIWEOsxB6oysfrHE8xoBv0wanDu8u2gEn+6s+rU/
72K98TeIagViQMqETjyhPzXaVgG47wNs3KHha7tj3LEUHe1KBCGfHIqLSGyuvlqweDIp/RdpG2xO
AhzKkH4fc99iQ9m/c6nOauDqpl9lfHp48wVDl9A6hMb2Gf8Oc2ohj4r6+vThwjGCD78URzUs6u2Z
LpVARo+2hhI202keJyT6pTs1ZP3S6SNJOKaNw33CsbrD/sNKEkDRjg3vJOdvhJP23f7RWn3tZkZL
biWOR4F/jNXDM3UJ9DX6NbdC9jgouj7zfoRP7qpRW+9ahOsT9drBFtRTs+hewETe5g0Xo83A0Hfb
OyVtr8v51N2oi/AG9ocL2dBifaEeNbU3QPJ60s4167Qvr7NdOvqnXU6JB8inhxqVRs2RAEyQXPyp
y+jgonZHjPW841RbY8YHMDda7ZXoBYjV/DQiB0lAKM73LsbzXDTtawVB6yPGWVYyO4pZDSjXrPvd
KWh7pQxy7jb9gIMUSv69c4AUvfLHcDzHpQg+cekERjXgdxW7fKmmqPzFFiLsg5foQhoFYJWyaFvy
cd5zVICwCzz+ckJ8ScqHXQsuZDVcoxfKG1sJO4nhfrJ3yf6sjRj/uZB2ZPbEOrREmY/lNjYdESWI
IrQExKlkwskHuldZca0UfiHNlT8xGtbXRxmrDS7rlGRckycX69o0u8YI6je+IwxMIaJjsynx7LKL
o+MlEUDGIbcW1p4Dft9ojKkSQ47BsrqEuyGIEYpdxZBet9L6khq1pb1NgdkbVpDULcqM6iKphJ+6
ZHzeuPsNJbggkKrPyt9v6/tJEaQcFtqpbRbNLT5Hl6I7jBMmQOhEj8JgcRatYicsVW3CtGOY9+Yt
oE9dKHN0DDAF1+scmbo/K1nGkCr2+PdgTffmMPrVGjs+QWYFBPg5/kcHZQXku7HARcDCp4vJ2SNq
jDamHPWim9x/K3qdLsEizZ2PDGBgx91KQMx1OH1Ygzd1Ua7rOJ66ISyOWPTtI3vaGRB8f0mEDII0
JPqmB/PTSmzmkJJ5WnbX4gAx7XbkwatxSk86U7Dy8Y1UROC5g46mUveSxMEhtKjY5YBDVRiY0Vop
sWiQKRRC718byJQsgTQM1GIQ6EAQKynXcKZFsn1kgBDwig4OiK4teKnKL1L5e17CAQ+hCBKTfqck
rSdtGcXP9eumr24LyIyTDh3mtB2bVugQ4qDPPtk2BnyqiNWpR58UyfSiJHCsE31gJcSINYujUu/d
XlIScLfpAVRBXr7cB1e3epOItdUdgg7lYdb7kEhZZtnme9BA7YIM7aXYdweqVXV4/CoCO3NIhCQz
xO4Wp8rmlWX69AbHYv6RR3DYSsKYeTh97heK54rr25MiXZCatkn4KmYuWs3FoFwff4pWs7Nrcc2a
uHdQIjwvbeMNYWJ2HjfVLIiu93kvEgAtFY3/y9vDSXxDJ2vfTFNtVugr27rVJS7l8+9zIiJ/oIt9
FeAbMHfPED9fYkCmMadFxSkkgNh40IJ6Oz/Kp+SyNZXnKAlaWSiupGAxNch4A2/xH0wPOnxQxhdC
tmkKUJxfBIzG2ZKDOSisV9Ehr5eYKuDSU8pIvQIkfE8CzgjOCYKQaVRjnvYKqqLGwH2VYK536CyN
68TbEXG19f7Nf1CpyvDcJG+uNORUsN89P0Nlt0sYk46iGYprwCvj0mw9RAysGfN/sgLrQ9r9slvr
P8M1mePQ88D0fOsKXNOL2ZJQmjwKbw4fn6rphwRGqWBWG65yFD8TOEGFhCyfAGMHNurVUsuc0AZi
gGdOa7HE1IeWS6BH8IkaHhN3DoRaTnlIoOtfGHvXPV4IMO2iXjIJwRpUJug52dfOQ57FYgyPKbuS
8P8rxSg2aBVp7nUxHt3wraSrpAA8A4SMXWWhfJTVXm0rR2j3H4k2Y2F/CSZkBDn7Bk/7E1oXJ88u
7MTGfdgMZ6I8cazZlgrpS0zeXQIU/y9H/WLzsbwo+A8JgYLBuTKYrcxd4+0TVMStf/Obo2NUU0Zo
Rx6ln5BtnW6yiPMv6uq9Hgt+rcMzXTJXb6m9OeDseFQva3gYl6IitQ/6Kq1zuN/2EPiYj5sbxX+B
2ZnfMPTU2FpYwXhEUXaBL0ZMWt9M59jXouSpbRdTEB9i+1YN8nkQwEPphPOsWh896elzDuL/Y0hm
fSGzQlm+vZ96Bz3i42I/Grpa0GHIrMAwKys1sJyedwKPfLBrcG+ezT8Hvb+D1M/tBk0lRiRA46I1
TqSqyUdIEkrXTTuMp9RgkAmyMfZkfw4KPYb+hy8RnQpwXsNzCApETjblMNT0Y1fi9lLk5673ciIu
5AlwhRDcmsXnYEOWhLRhBXbIlK5z1moOxe+r1jVz77xD+qrnfwTmMYFUP5wr3XTUbZ0vva5xvnfL
bjh9JjharSAP+FNlw6c0Ef3o1FzD9JD2glc9IHQioXK4jze2M4y3bnndLugYGiyeKMSRZ0tLvgt6
IbG84+Z90wmGiIoF9ef8ETGucC2/ylQD3tdqLzBoevRvyzH6llISxmO/lqQYGWOCAo2V6K2ermB5
yYmAK5j2+MCr+F8qrjpSJbtFziqsUzBszRaEVCAcWFjaZHqOpXi2XUGYdJbxLQl5bSdYumpgt2tW
m8H5laHdp4Gs8HUZIe7z6Ys9vmt4c+5GxlVxy5T25NqtvFU62N0YHRJL4cKhqXuqjTwbYioEAd0X
OPiKKXLN/6PGSKtN30r9MG2+oBOVe7w+jJJraEWOKU/q7E8vZWwN4Ro78gveGFQiWoYZg9zak9we
I3vveoKZ6EPZll7gyP0VEV3b9caIMHzJ68GXEmhYLvdAi7RFk3rHCbqbLmc5jDKpFlvV9Cj0dbcN
tcB0c+lebP9umGNgoj7iwiggKITYJOjAJCcP7eekfqjhzPlhsATc6M80ro9lJtQrzssZZNtxehxe
XnYRwtHOGrd7XwWG/iYiWb807481i4oA9KRVACblt0EaiqxuMXm2QKfT6uOq0v18RYHi2H27ntAr
Whg7uqzj06dEx9GP1iltm/zggdJdW29klsyifW/RxNp9EJhqwylFfk6M2Gx4XPTHiUjPxF57g639
AfbY55J6J+zhoj8deGmPAf5RzBes0h1fIDUhj1Z2ZM7u9ujaTwGx/B8f+s5+Yrn4hUN0notDmDSj
oD38Z2i96/7/ZfNVkGSTbQrc0zahNNEfDehkOMfYJvKhyTLq4MpKbAnNly2O+WldxG7J/XWKJ8t2
xW0GaOQ0jLqSJuQaNYOgVMNhtvhy+t73SEddqRFqBAmSipVfAF/8ClmjEk5yrGePrsP4NyR75PQH
WFbTWJmLjFWXNjqKe5489fGvfvPjct1CgFm/Ya5O/h2+9QfpD07HH1C3Lix0KyQflHLKOKDIkE0c
Lm2iO3oPpPKYZEvYLwrOP7Mk0qi+w5xoqWEnG46cYyuFhyIL1CPYale/vs7UCNNz1o3bi4LlbVvR
OKe1IKGneL5ON9/bfPIGOeRqT//+a4YuMg/4M0QKo4opZo0q4XV+iu2P9sM/OTvvP1lLRcL3Cnn5
je7EIq4eTW6aMKvXBkZxKkvd9uwXUjXtvla/MML+JNzkZqBVS3uORy/Bi69nNTrZBWITCb+NM4nd
OIMhVNfdC0dYof0GPyUig34fmW/6cdchzrouqSXB8XvTEPle/whDMtbMXs+K72UAqmO5+z7xsVZN
+D07CDUXrZaJAj09GXee/q4QTtmBTWakq0pI0zZIHMJEYLmoANrJks6dllqZMpt+xfqvzo/ZmgEU
GPj+YqolC+f3MTsDlcL9/QQwuHZrMo2r3CZNQT6bj108FGbPJPvsXRM+UFV7Go4/9EQxO3QOxzbI
qY3/vKXpGnKsGX0VVAR29n5EQ7GmmGcZNoy3Lh5kVe3EqjcLpdi0xxWJL+XlsluGENTUEcGPza9R
fzRLyFeFgwfxyhmBFjcbjLBXlPYcmv5U+QGun38hNvlQMql67GQQbCrzotFy58InW73RvMNFLkq7
4Qlucp7Ho9WFk49chVIRi/ckz4xHm5SyGV5oNpw/1mx1X/jKUnsRGx3Q1grpWcB8i3Y7XiThj/gU
bmGc9qTiCnZBNha79bm3f/1kcbbsNj1hz3gZ85PACOxQ/3LF992zQAgjHR8HahJCEJplAeLMvBCi
GVi0jpkWsoLZXpNm97mqf20f8v8U+jrTdv7nXYmS42guFawzNNLmZ+8iG6E7nXMG2a9dAM4m5+XG
mqUVz643cNIVr7x/30y42oJNt3uV1Sh+pDq5DtMegroGV0tlNXxzYWARCnz8dZAkGiOZ+KFzzGEo
EjnaC5I8PrxbJr8sqJWiuy+PBIS8FWkFM9FK8K35iuCCnfoj3imUD9sEiIHLUNi6VM/zUXP/JsdT
vtClWmbcW5Tut5MskFOGwxJylryahAaDaWdbmtXJnbSdToKD/a3SSKx52n9YEJxzbSPUZNMJx5kL
gY9RjfR7arYw2y2QzpjqojDJVuO3kKg8muboeuh1lPxvhQntk2abdgv8FoHRU6PpStfsm9x6dmZB
hD1HLQbNCrZCMfyiOlbkeslMIE5C53WXxZfRICAEIiWYtlbO7/liW7hy6Q3O9agZM+c9XK+dU7N2
bMuLjv4T035mY/D6vyI9BcAxW5lZMEOzT2jf9mjvNAr5MRM7mPv5uu5gxei1nuP9xevnEtMo8OOF
QmhoyEVeHP2dLsNJPEoSrF4Db9PCijfaT6D+i7dwtwxjViMILkbSt7NSKaE2PwJ60CLmlbZeRqvW
y58RqEc75+lqe9pV34BqgUjD2yK2ymv0od14XMZa892WqvP15qeyQbcORtH/u58l3I323GCuAJsd
HUDvpl5G7fpEddJaTfYVUDcEPGPGxAwQJ+s5qxBMrdOMGhDB9POZ5u6eUhupEq00mK1utrecnSKJ
goVDW+8x1AKBAG8MnFu5qZILEubWrOeYxZqVmiGe3vE/K1tTWDdNuGlkwz4+z7UdB7tR5FfM62xs
X+OEC5nYF6c69x7donuCG2amUDMCPqq6CdN45gLA7BwIiucnupHoj661eoihN6yHY+6SXnXVF5bl
vionSYlSjZVsAxHcScXshumKi68yqiuYqFkRNHkqLLm72Q4oS4YAp5YL76QddFs1ILRepOVaJW20
3cw5Zjz9iMc7o+W7GFadDjXZ2IM/hcVm7obrTXgXEbG3lROH1/ysTtJNLaf20M/HJMaCOjp9sOpj
DVyzdZ4dDbz/JXYoEq7ulvDaY8tB7KqhzxqpJEMhdjNpCpJnnNZ8Ez+OVU+kJSQfU+mujn/xhz7P
hxqb6VNoQKkVua2Y0JJBAJzNegWC5SQquv84Sv0t64o9are1Cduzwca3/Bg6VxCYQNJQqK9CV/1f
u/9o4v8ejHBUF0gBD00amzwfQUsNMVe2o5gvFhH6eU93NddJ3TtdwB2axw6tvsNRWJgtlS1QtNGf
ek4B9E91PE7XkgFk2Nt53IhrilMRxMQgaDvsAHSjWQBUk8Cn6vwQ539/Rl/SP3sYE6wV1JvxMA/D
OU+jnOwYocwF7IXk7cyKm4nWN1r6f29azrSjDoTDTyw80ncY2K7dZ4+pLEiuyJGlrpGTu6PeZTBI
NwDzefS70cdR2SS8QVQKkKniOZAhCGxetsj3NDEzkMPDUeO4KqnWM/8WD1mDNpU2tso9GpvJT5fz
seTYU/y5Hj1Wldm2hKiSSnNNWfieGmd0ZPzuqRSh4vaHlnkehvRARvej+f9H1dh+qTbG62f1n5lO
akML8sgtbzrM3zX0CPNysxIMA1FgQTFEQX8dvitjxE+6VAkBgT+cyqSoxrCUvbTDCbhqYZN0tBrj
0gE+/7fy16Oi8/L3BC/nDFXSX7O9DSJrTPp+Gf29+QsuSOnUX5x3OxOKijh37ZNxghpzD506BP6V
0QqBKlu9hOcKlz9LO41oOTML6EEymcRNjV/M+Wil0JwCVgZhIw343YDAc1mbejmdQujnBqQZD7zj
HCBdSyfudWOcjmSNTunomP3Yt7xQARbSy/T6cdK3L42FU9Qu/VTSRU4KFatjjwQsMOyflCzrRjED
UgS6TDUfkItoySbKLTYRm66Ux/YYVyYb2wLEEJZzC3WpfLSmyfWr8Iz8+kclGkM1DpuiqqI/OPo6
LZkwbnpwaFdKNYNHRzGxbcQ7F55nkZM4dmFKiXNnhpgQjCTc/A9tqxWU7iQAtbrqaW6GcG/60Hue
m/3gaMMoxNWoCctOTCJVoeyyP/RqtS/vtFVVmOynEnZiOzhkzUFt5trqsyhCpIoZmjGFYTGG3b61
zM4+KAj7DxBGKZPSSo8ocWwNJmNZMZB/A/nxjmPLOnc28CGg2hjqUjvsA3MiYsno6O3HLzIh5YEH
n0JbF/B6DGuu6JXyohqT4M5m1ugbhKwvuSuuSLMGpk4r39ZYGs1YGOoDC75nIPjYk5337gxY0uuN
B+oirhCDeWOCRiaZzTv4UZmJmD4+enSn5xXsF3c+vGreZh65TR0GHO3wB9PbFnfFEpTgJHY0t3oi
qBR4MeQSVuvitDIKPyN7QT/2sTBTwdTcqivZL811BIVmVTej1MjPgwH7xXzYG1h6Rl42/DU9v+NU
jz0z+DmSc40MIAwkw2DHorjAVy7YHPg4weyEQ4VlVVaiCCpuXNtsDixy6A3VNvUWv0pe3zihPYOk
lsGwfpeiRJ5hDE1P2LpPellVbnLl
`protect end_protected
