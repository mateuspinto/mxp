��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��О�C�?���'G��p�q��R{�ZWn�`�ޗ2=o.��:ͼ���ZX�N�)�^�V�9��,�!�� W��ƥ'2����q�L%Ţ5�MS�NA���Bc;x%pC4���H'�(���@Z<�+w��M��0=��{��#�66��d�E���Q?kp��ǡO��;
��D"�ޝ�[ޥ� �>�B�,8M�Z�WxՆ}]�[�w�e�X���JѬ��6sJ�K�L���*��Z�����[�yE�ӡ���k���п:�/�_�G@����2�h)Pr1��XP�SB�Q�k�XlմH^�1_9Z��G�W`�6xΞ��rc��X���ٜV�n�g�N��f�<$C�
�jP���
)V'O/>��^�j�w���ޒ�ԏϵ�p��}gu�x����������Xp|#ټ�7+��9&���-���u����bVسmϒ��D']�\pk��C��iT,��أ��30����]�TaR;Į�>�|��o<�B�v��2�n/�P[/0QL�>�@�6���j��d"��H���ǌ��L?AOY��ڌ�j��6	���c.�ݳ���"�&��^���W�5�ċ�ti�0����K:X�݆�=%��ݴ�k�lgT,Z�hz�'��H�|���j�݇�l�C�oz;��^���I�9E
=Js�Y⯭�'��2zP#��"b�_s�����2�7������3Ϭ!G:�����Si;�ȣ�A�pE�ɶ�J i0�Ğ��֧Q\�@�S���%R 
�vg� ���hL�#7w�9�z�o�Ua���k��k����85�=�}&���CMd~;�+i���i�r�A`��g��>1�@���*P��V�i:� ��;�bHR[�u:541���F��x�7�q��#��t��abgn�ūY�4�qch|6�.r� �Չ�FkM�*��Z򨹎�i��nC���`N/���Q�٤�\��{�]N�����G���`�SN����Õ�(C(?��<�W���0/zU������R�\D�*�����.y�2�f��\w/CVP]���~�<jk�,�u�A��,�(����^�&�RO?�.�%��F����"=�U�ȱš�s�� ��s�&67�T�=�@
>�Lk��j8��x�G�(R-���XkJ*���Y(�����
��#V�Y�3���h���Д����
W�Y�H-��K�]SMf�p{���z ��*�@h�QU�����OUm�dJ{7���}L�"���K�&^
�df�X���](#��|Q��L㝗����]�2��ٻ��)K�[�kI�=(��*=u1��W���>!a�����]钣[B���!DҔ�$-�v�I��V��v��y�ݕ�����d�ܨ�5��m���߄�~9�	;�bp�M2���\�k�RS����?�x�^��dM�Yj�4�Yj�^�����r.�����Ȫ^?�A�}�����8mGllF��ʬB�A^ܾ�&y�`�|m�ʿ�X|44�]�m�Aή����a�;�\��-��4�Oԟs;�SDv2c|�b��g�bR���%���s/T4�dL��j��؈��d,N*?x�����]l)���xm�}d�}�G1s�уv����ʔ�~�	�n��PSFx��&D�+E�S����i!/*��3�������d�����U2C�/�Fh���م��/�\X���!G�;� ���L��x�b̬"2���*l�u�S �I�X�����L��p)ܑ�깞႑ށ�2=�5q�"�f����Tv��[DsI����馱�!��-U�W4�^�gG��G���hի��S0��ߖg�I�!U���`���`��������($�� ���S8 dJǊZ��ӕ�e����l�����'��.�U���֦�z[����f�!�(!� نh㶍9q )�[�������2&�R`
����cx��]'�^���l�,���~��<7yCB�k�-�u:S(�k1���HD*��*�3�AJ��me�<�h���3kc�X�����,+��	���˩���@�:/�bZ��w<�j�32�h�4���e��R2��ǒ|U��V~�r0���>���2ྂ	�V�5��uZ�<:;�	�#�p���{�ۡ=2cr�7��h6�uG<��ڑo�>q�n8i��F#�J�"���c0[�u\3J�q-?����S�!l��#A�7Y?�HD��)�`~�l5=��XQS���(�.-V���K���G��Sj�� H�/��i�N�e3i��g���մ_�����8�Pn�䡓�>� �ohR�=�j�{Z���Im�v"d��R(l�\���T�����+V@Gi�X
�:�(+W��w��J.��ٌ�l��c7�"�#I�{�%���l�MKɂp��X=s��ᴉ\W�C&��ձn��W�|9r�f{A/�^ĉ�780��L�k���@1�w�t�������Nfy'�Ix��M�YZ���Ӛ�چi���Y���,�X���.�Hxz�a�H� Iّ,P�ꑝ�V��BvFW�N���f3��%>�"����h	 v�A�c�b�W"�8�&� <��1��)-R��I@�?.���e��/l�}e�_�f�f?�����^u������H���r�x�T���K8i�ܥ��V^lo�x�3�����ՙ��/$��H��e��?D�2�Q�]��?�1);�:g:�#��!����X���$4
S\��S^W#h�����`� �\ʭM����*����B )C���}� `F�c��l8����b�O���:�1$!�Y�����˳��z9죾�,2ѼFV�9~΋E8��h��22���G�v�2�&ޝ��0H����-{r��h�� M�)��ȻD��h�����*[�֊0��;�l���"��� T��u�!{A�A��־0�pi��o�v�1L�w�#��((�R� +�3��mB�����J�3�ch`�q�/L���*)nC��V�w�G�����J]����tAf��l�8ɵ�����ղ�� ��!���;׻h��1�蔅hnX&Ԣ�
Af�s��e�ő�1�q4s���$~���h�	TN�r�kC���<�\��eP�f��7��y�OT	P��I�Uc�ؓQ���[]}x�ϡP<섣�@̃��xD|�1\(�a�EBA睭W@�*�p��Si_:l5nH�v��@Nn��H�`n��]_�_+�u 9��4�/���s3Sq#E�Yݰ���\�j�G}�����ܗo
�F��c
�2��������:���{�~��%q����4���T��\��O�a 5��9�����=�6X~���[ex��2��p��U��6H���]}p�_M<%�cS��" ��}��CK2�tM�*(P��
F�����Vc�j�˖ò.0� ���Ȯ>'�*2)���Tn�+�Z�C��΂��!�ͼ�Zb���XbM֨�H)���������9�@
u"S@����{2��0hP��������ɝχ]���Re1SyF).B<�=��qf��֕���t`h��'�n��D�LuUI*���i�eJv���)}��������Yq�S�oJ�J �u��)���c?M��"fQ>�'�Oh���T�*���:.�r���B<$|Pu<�"r�x�ד��3|ar��鳠���YȦ�o�@.n؈����Q��z�J�5�3>rm����p�+��թ�\��s`2��,�zL���2��iB�Z�1��*�t����l��р��}ԫç3��@��w Qk��j��!R�q�b�b��PM!��^}���p�_P���+*�C��ʝGx��-������̂�9x��?�P��4�%;I��j����T�IS����+�3w�`f"�����������,�,��4�7\��Ud~,{�OզE�s�b��Jteze�R�q6?2Knɦ��߲����Iu�1+b�;S!��_��S�UI[_Ȕ�Ԣl@~TB��+���	���D38k� Gnzl_$����f�DJ����7��/X���ɲf~�����V�u!cK����N
��S�'$?^�A��_o�@��CQ��l��*�P"���і5g�=ʐ�|�����f\� ��4�����L�@��*HM+"3D�ݮR"�|���`��0�$�|��4�T�}�	 G�~G��]U����)rn�C�w��>7g���ǤP4�FѾ�����J{Z�5w)Y7F� }��A���m����=^��þ�u���'���(��Ė��6���Eº��rL��=��e<*���:xH��0+��z�5f��+{h���	���*��J䚫 �|'ὁ�6�������婧�����IT��2?*�~1>��'��G�	j�U�rI��?�י�����ѹc��͜#��~N��o�l��7A�ᆇ�-��`Zc������Sz`<����55�f]�}�=�j�j!�:A�����p�H��sti���47括0c#+��ݰ���e��$�Ag^RS���z��-s-�<�샲dwC�����3�@�\��z]Pzf�F�o�n�j4���ڰXIwj�
��d5T��ĉ�]���Y�g���Z�&��� o�ܩ>���WLzĻ�jA�o�(��D?~�����Fi�E/B�^�!
j���p*�;o0Gbw����%�a �=���$�%���)�s�>#����?�\[ﯹ������k"�� ��!�)váU�م��f�l���'Mbp���%2V��_ie��H�\w�w���L�!��`1��܇V�"� ����A��-���,%)��:�g_vU�z��3�2��v.8�҉g����4؊�j%"���%� ˉ�����Dv�vi�h��g;S��8��Fk�9��D1�␊_V]��v�|��W����أ6��-ۏ�� ��v����K�	Ņ�z�}$Xh&:�d�d����3B}�p�`a8]�*ʓ��onFFM}�����tPxK�ڑpp�P��fH�Ez>K�
�����-9�j4��Tr;h0�;N�~e7��3D>)1�З=�@��*�8����<��OP�5p,����h!�X1�T E��v��n���&�4BU.,lAr����s��������\ĶC>X_������䑤�U�
)B|�L�����ܐ"z�x(�0M|��ќU���&��+X[tS��9�O�1��E�?Hd�tO�5��c	L�ӓ��Ё.�m��H��;�n�t�4�4+|uxV�$���B������c
�'�)��o�D�wqʰ�ReAe9�[�67���X���mz��|����[�-���Q��(%���1��*|�.�*檛+�JRJ�����+�WY%�!���`��`�J\_��"ib~"�Ov�#�|�/6�ޤ��"v-��~�h�hjhH�S�;�vi9>�f��szN����J�~���I5~�RD���`�Ə��Z�F$�3��:���. �ENTi
�+Q.ṳN�c-�z�ħ
��N��yg���Ӱ��q�U�jG�*f3P���=�G�Z=+]�x�t>m9H��q߯��첹v`%�/:�+���2����+�S�;��(*U��I~J�m/���Rl��G�ޥ��C�;���������|˶���i��e��v�Ciaa�9c۪���w?-�T���_�ܵ��~�׽�>*�`�wGyM|��.�?mEG�1�$�;��ɱLvf����K,�� Ճ��L��v�h�J�� �p`�B������dX�4�KA��C��ɹ������+z�j��AԞ�u!���>M�ts �l6+�	����<�(Vt����y�>��_��)�S��p9h�ⓑ��f��R4Ν^�V$t��Q�U�ځW=\	�7�c������gɑ�9�|�tz�֨�NrA�ݍB�[�.}cӍ7%���\1�A� ��]��Mt����)��'&CĤ�!'4B�$��?,�!	���#����~oOfa(�
 �H�Ӥe���2��_��q�$�W�uZ6^I<9��x¼y�>��A��Q~T�^-x^4K�����q�r�� jj�z Y"0�Ĝ?�/,Ce
�PHWO>���-J��ْ,�R�9.��7���e���*���_M�Z3R�R��?uyz�%Q�a:,�ү��֨LC�A9��k���u�i� ��b��^��I�cg͛g��.���QV���x:Ė������"?�N���ޘ@���o��