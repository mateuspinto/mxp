`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
GHdkgJ4gW5/Zja5CXPucJfHh24RyRMgsy/sNB6URZ7CEFnWCfeKKHJLUvGA3mDYDy+VSBMyiJWTV
bEX82vy+qJ7gDEYQ6yh9Y31CvF5xFTVfC1JW7o5WsQqI4LEhJ2dpSdRHQ1UaIa2pJsUwWODrzQ3p
xCnCNbVbX1CS3kx9oIUhRpZ6RjeX13kHPVuLMR+G9orKum/uljy4AxDTA1fnTv2Fmig45M7bzipG
p15cXF1N5pmW2qBBgBdFQQ9hZZlxIbPYUA9FdYlCXJCLJMjRGKRRsjZlqty7ZstAM+r4XNw9Snq0
13lGSkFP7Bk3sd3Cuuj/EkvbndXYcqFOsRXu0g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="ib81SCXA/rvKbSiHN07ySniDYUoyjmEKVZ9F2xRO85E="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3872)
`protect data_block
Qblqi+pkloKefyqycA69PnrePu+oIfQIV8DcXJGqPZ86poL8si0yZf3FsTQK9GAR8PFeP13UnfZg
AA7pLKdzN0AB9CMElrESUTCekjtNlOdmruIs6+fy/WWlSduAFpyTFoNJmOq5h1L31ByPBuQJAIhc
AJu7QS/jVBbnxYAQCais3haMGcmppcV8bXGw1vngoDb5B6gdUjDDkQG/GFm2IAFkTYWwH8n4by6J
Os3l9V3KLXb+iv4OhIeWcR15mGX0PlEffNIHP5e4rEz8z/dkRNgAORT47vqpjWnoTr7KcpIO6xBn
1kcAGls+gQh/81s1bin88ntfL9J+LEDnz6warcOzmrkAb4Qkq47QT9ytD+Eg13Cfd+eZxMT3R7qo
bJ8pxxE9gALD5Oeqk79F6+Z912kATu8bQk6A3PByPzhf4lPUhEu+38zguVc+JrV3awG11svu8REO
otfhvQLP9d1S5wbsUyjjZdr3+K/h6H0pdeaYMxmTWaE7m1b5or8b6No4wz3ZrTmxD7F0JlfB9o6N
uMFLvC2Ia9TloAMQjsUK+QkMNN5pNc9JD2E4k2DckrL+2sofW347CfiWvnu4c7rF4qWp6vot2Uz1
uP79mCK0JZpBAtVTVNyHihGfU7AHyP4arpAfbH0E4DvgACzMFHfaZmtd5/NTX0/mlV5+3NQw3mxK
Lnwq565TgmzejFZfxSeK7uAXZwjgCUGvmBR6kV1ZjZ0nh8LMDG2Epbf933KMyaMGSogrJZVUoefa
noSs0aJopPTtf3FNnEawZ/0U6Moai2mfOEiRjBJxxS3wYRb8/0geWWcIwtOib75LGbfMlICKh/z1
1rddyLYTvm6MVsVbBmwp75e4sIi3rKP686VexAqH1Mu0OD3PfwL+8UTKe/KWAE1efL5zVt+n+LT3
TjeeKBfxoV1jHfnzfai6GPc7cvvtAFxWwqcu9K4jUOqEbNO2Tb8sqW3KnN6SUkjt+qbfdvo4BsEX
PNXedJ3ji4hmmVnQFC2E1ru1k1yyoQ6F5MSlGgCgtU0qwNNLLngk9xjsu2qHJsxr5DDqkkk4fbKt
7fy7/jeKx5ir0e0c0fHdjHWiJVovIMzcWzgF7uzkVlSIoC8a2/2+jwEjtCdORc9IfJUXXPBM2MIK
6LfC//KcyxcHAX9cguXSXMDoOoXXKQ4kO7NxtgImw+v7DKBJiu444yYB5yHmXACFNAVV2UHeO6IX
HakJE5ph0HCAhyvcaEpXAaG361L4fXqtu+S7A7ut8vqxyuIlEj2rkTOIbtt0nHlcLuXwDAQZ9UlV
b5snY3G0gwH3vMDG7zcjB1DuIKdz9EZPAB8mXO4W9gyqRshAjLL4MAu6llj07D31RM075HFAMjxQ
aH4w7L1Je6suop6imVillhnK2oZK74DP0zs8artDy+LCP6rd6syjWgzGVDtZhmesyL9RfmWFtocp
Gfpi7zuS/WB/W1ncI7Roq5mQDWZpafYu+Ij5DS3ihguWmBHyKuzYCseFYzSRlR3ApvuF+Fz1vTFQ
V2vtduUP94QKRsFbxXJrlVnz9DRzOzujqRtETIS4t0TZF3ZfQhVJtiyM1Dcxrh17E0UDitQ7DUEG
Ss9RxV8mVZ/v24iWT78+FLGqUe2Yfr7vZVNUT3bKLPZUGPfC2JKH74UXw6NJ2+HREEdcWwJ671Sp
9BgJAPMYaVFwOy3t+M3prC8YlWWil97r36d8dnUDUHTyozTnTqJNGxNSOLuntspDZP40BbHvsiNq
u7vLWd1+4WKjfrruEkbgqe/mggt+x2S39hMVPNji0rY5CBr9cDAM+rOET7RB0PfKUY0bGFn3ZDaO
WVy3G+8pYbVGxqSnPPxuBe1G6gzQ9aedc7SXCcAyryajxo5WFNAsZ4A+3gRBZ+lr2gQZUZ7JIIW6
vngycMNaEt+9mx4xO2N/yIcAomH2uW66YiU0ekcCESkDH31oocP1b3GlP30UfeA4MjGqbUKtBNe4
cW+UAixJF1cMnBFQ7OGC3fnwfoSz84tQO81hAAW+1xhmLg+39h+i6nGVQXqITyO06ZISrAKrnDvu
xQYu6ARoejHPqqtyWcuLl18LwuLHCtkYTsSCVIdOGSRGJnwVhb97D8PpJYZV0g7WSlA9sFcx1+1s
UMpbUAYxX+dJTrpYd8FFiOMH9ho3wrpGodLaADgw4kJ+vDAaqmTFk44kbqp/kyuXSupcE1MiW3Cq
PVqA/M4X8/QJZle735MKCsgsp6mbkOtON+i2MwCE2fbW3P2A70kZFN/FWi+0T5hIm3dr8zVrKwf8
lXHv7zpxwg9tG6yw58Rj4sCuSdPkqxL1ig4lIBJFZOpD9srrggKxLx9Apz4RJhYRjF2wroKS7tgP
iVhGcXfHHrCgFTBgffh1F3fF5ilUly99qi8DhZtKXB+bN4G1NHo35y9TykfUHGiS7uWjrODaoRyI
TcpTSt19snSjyenVkBNzHqVy+XW/TCfDfPPQI9dhlF6533rFyyc3rhzX+AEkjP5qHp0sYUjc9CLY
oAgcvEcWWuYi/lHfqntQMIGfy3MvovTfUbxY97LCZvSWDsdk9If4m+VfGRdi7+NDs3Qtl62XgXG2
MdrN3MY5n99eUcerzxpOyL7xuTmZotHsaTqupWz5SqNtRe3pTNVB7h16H8TqS/wStewxRnVCUhcD
1V9AIRBhWDKQPlZAv9FqEkHKm/dsty+yEcE5apNX5NM4fn096DS88L+O805FqOkfthjHdA/nanW+
kW8ag6NAv5uVXROkkrJRNJ4ksEU5EWTTQ26XnTYwXHzRGBL7/Exn4CDeHVEN6MegsVnJUDCi8Fxa
xkiD//P6aECKu11GiseimL4JXCgzjaCyzBLO8FQKDxdItqZ7iuqG6p1MvI/t9I7pwz03J9CxV+Xp
F3TRqREbkCY6kZhlcDN5cy9i4tN/ZE0dcmO+EbWQ/fVDRRRE8baQKf6jStSfXM0oICl8SqerTuCU
iGmq/AYIVl7w/3yl5EXzvWB2GuSmH878BNAxLUa6zIo9Be4GDG0Fzs4F01v0ew3Z0xe9TYYl8ixp
wRiTDLcAEi2O1IIBRCTaIIxIShg2ywI+1mqk/jeIEJmqGNe24jXIZ3DFoYwt1koDgfxZOC7GqeAS
vhLW9s313Mnfiq+DWneQEd0VfnezHz0zrUT8D56Q5Rn/89mHZNoS0ZF+cyw0z9JTSE94K18uevRq
49pWQrik3ZuOh8p4nzbQE1+GO8wHIPqv+WFY//ZKkCruxHs9pFrz2wyZxhkt0TYM6SMBt8YN8BiH
SoQz1jIaHVrFUpgloinwb8L7dCZVt8NMb0ISL123hVpRCm8ZCroSo+VNYIHwr/z8R6OWUpTzN+CG
rJ6FhCjJFn/ep+IVvU2IvWBFjZKzm3maDSycvVJjB/eNQGllF4H1ZnRMQwPFZYRCw7bYGV94QgY4
7CbpKNqOEHIP9D2D6xkhEY/X6DRK5yaCiHCDQGhnzyBd+6yNrx01QDGx7mQBGEiMNi67e/DJVzj5
SzzFUkOx4R/MCWsfPUkivdHupb9AMJgn839NKn6MIXTeWIx9PENkJGw4hHetpfkOZXfIhETv6HnA
0rAhXKEvrKlR+YkBGZjzA3ggJb7I+6CQYbZNiS6IxQCLd3z5HqsqEyJywFRJJ7hnCIU/oxxa+7Ex
g/Ugc7QWlMlxhVFx9MNWfA1LS73Nyf6luYzNUFO/5nzcMEA9IspTRt9At2vf6Jc4c/z97XLvzkQs
eNdaPhECA7Q6PaVwHpbismMVPUdkK/92jo2yfobYyAEV5kT3zat5XKIBHcJIQW0SSwLliHqfwf7p
vaeTkjsdmwQwmdm398p2EfZqORya2xg+M5nPHkFz47tng4V6hw17wblfo/9tn3/k0od2CJpchiyr
R0bo9Nv6FXxQTXDqFaxcY2jJEG+NAHzf37FKPolsCvYtivCE0yt6MPqOI4ymtVmWiNrd6mEZTtqH
/zUrE1V4qEEE9793sWId+jLJGkq4YktFPUpbfy9LTWbrWtsBaOoFrVGrUrm9mSs71sgDpX2hdQzD
xDpavzT/xwNwXBLS7Z3pTNWdkqyLPErxVFCUHNPI5cWhme+gHMhYKOnE11JWJ76dpPD3Os8V0k0F
RELSeuvdYamkVPuUryrxGFkNYG62ZX9xzBprnqtaVKacgttS/wQD4qnJ7bMnOmJHeODoMKDugc3X
dRVNz2hgIK7Z3ItxepSQwX9PSJ6b/bPIGfo1XXut++FN75mxq2SlkH4m1/QBUE0lm1xcmT0+rT+i
1FNymkyRSDLCFefMQmcBhrUGUz6/1FL6WjMTiPUfSdjNk8kz09E9ocEjXhTnoKp+H4lUTr+vEXIZ
xFuTw+AwDVsWJ8m0CC6YVAwOn7dB51Bj3LgtLx5k6/yBNGaTniXZGPiEousBLhf08l8GZczzZ0wX
QFO8vMT8Z8aKW7ZK+49L0gYFjkSl0Fojh9jYS5o7ZZt/h5k6qnChp/oUVmuL4rFz2tZL2rOv2BOE
PUvuoTZbXCwtxPNIzDdiiihhaMiH2xPio01brkk2j3YT9kmM5Pruork00rKXGOOK9o9MrMAgew6O
Tkq3VAvYiHuJseHF2Gnc025QBoFPK+L48U4Sfkb6Y3uDNVkxbrgGC5Gpafi+UcWrfArOEb3qP+5r
g37xZPmG+ihhuWLS07pECLILo2Yih901OzaAzY+n+/jHR9k490SReEIyMkOkCNNG8T4GcAEVcohx
+hUkxEZ+Db2eNyRTr2nA9KDDsYC7g30/3n/3jgP6LxmHA5NbBAtLmZjh0PbGDeGnY7/OdxLjzbct
JoVDCwscRSmoj/ZKWJ8BhgCW+TvZfnyoK5/sElwhf9gpk5iWj5btiUKJEJqn8B91GqkkALHFrnJ9
2C0wzvculX9A39jZy+g/WI7pWTxZO89lmvmqdnkGFtZ7ClVu86zm/F/DTfROBeriZ9dUW/Kmixwe
4zlJ8hWvnLA9fGcAAqqp1dN27ChiDF82+MTjn2U7lTLTJyyVWjIJj7ng23AaI/SGfV3SYJ5Cbu04
Ldi2+wEYtSwh8b9AQ2bp6S95Ma1F56gKyJr8MHtMv493/VqxSKzDPL9xK3AQgmd1CpIWSgw3i8YW
xccAVZRJNCvb+8uWy7HYQmf43AeBJdPq5ZLM+hNAVOs9rWJVKF9NfAqxK1diFaTmXa9VMAg=
`protect end_protected
