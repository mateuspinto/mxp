XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��@��
��ݶ����݊�C�Wʔ�!��[*�A�����i�a�4�������?_�J�9����f�b�P���>���f��f����H��T0ڹhW�������"��&���ZQ#���y�w���E��q��pP���
��dr&��'~7x�ʋ�V�}VLG+����)5֎��"aQ�S�&��@b��1vQ�����ľu��%&���M���̃�NxC,�8H��e��L�� f�0�d���,�2�T �[�0B*�1 ���l�ۡᕼ7�lWН����z��� ��9�wdmR�?ٴaK�l+#�Ǯ�,���Z�R�d��E��42N�隯y>��v�n�+0OQY`~a~��\y%���=��!��8�/GR���[�	��a�h��:;��d�jd��G�cs��|�������uRg������掔�Giw�H�U`9�����6�D�A�W6�Ǫ)�B'z�Jַ�^<�6<݂P!���%�$q���pa�qCX��{�[
���� �ᜀH�R&�����$�@�+�~i�"wO�f�MON���+�[��, ^�?��K��%�������V�kVE�@����8���QI��)�xZu��� 'm3����d��zi���xx�l�{���F��S�}X@Vs���>'��~ь��ߕ�p8Π�ݱ9Q��i�_I=�E��Ce�Љ�$�~�]��/��h�,�@�g��N��PՒ��R7��V0� Jb",�Q���[ԀOXlxVHYEB     400     1c0_��ig��4t�ʸŘ�B�	<��b���s�ؤ
.:l<���B���ӳԿ�[o��$�$������P��k�A��U�a6�:2ֻ-��%�U8ӭ��āu�Ck?)9��ZEr�B`;=�3�#OU�"[4}�?u�%��j����m�V����˝l&�C��=�'�F��	8Ȓ�����O�r���m���rAӈఫ[=
�]\��)r1�M!vmb]��Ėc^6�O��vKb��S]�f�{���>�f�6��,l���+"g��B�0W���Y� cb#s�H����G�����"��o� ��䎾䮥\��35��-�Ϣ=�,��=d���^�,s�J&<�jƚ
h�c=�q��3���%Т��nR�q��s(�_d��1̊)�Q����H�ZUo ���>됌f 
�U�Yt7.~�e�A�+d��� -������RcXlxVHYEB     400     150�;.Xe����>GA�O�.�g�&�\C*�У��aOof�F�����Y����7��	�+�4�9�_�Q)�K��S9󦷄݊���r�ر��1ͭ���Jӕv��1XHgT>�_D���8�"8���V�x"�.��f�����Q�{�)X?��dXc�)A�ר�2��t$�db�W����Y�T��q?���m��bCcU+*�4��B��|�ɶ��@�z���]����@p)h��V�� ��a/��Im
��Jӳ�!s�T��}�xh�>�ۅ7�OQ��C�c\��
^ sN)BO}w�ӝ�T����<	U>����rXlxVHYEB     400     130�{;.Vݺ�J�Av`uA�x��BH?�[_�H�q�U�'�~(\T~IƶݴN�/�,Ǔ���=�ڝ�a.�ƮB^C�݇��=n�� ސQ!�b�KĶX�-�U���lCk�T����ș�)�̿�h#SA�k�\��\@K�\x�`�V����ʹM�.B�FB��M.��R�TmP��SZ��$��x���������d�M����ŗ����ߦ\i^泟
�oI�Ѱ��Q�ʯ)@�P���R�r���CF�=U!���Cq��x�o�� h��lk>9��0��r��\���a�pXlxVHYEB     400     160n�k� �_a�Nc�O5o�<�9+�0�����W-�(�­���­c#y�0zLu$%cɘ�;EF���t���5	�M>c�|�}����Ff<w�{�.į\�,�C��9�E/�`!�j�_�*�T��Pf��P$���n.���J1���,��t5/)I�)�~TI��ND��]�Hu�=�ELoymiA}u� �)]��1�yMϗ��+А�?��&
�(UL	L?mcհ��e�_me�F��ʨ�C<�����-�z�<,grG
�ܲpa����]�k��F��׈�f��!��FqZ�1]��'<"��b!�n�Y�vjb/Eƿ����2���XlxVHYEB     400     1e0�y��r�~O%l� a��*�9u�YrSׯT��%y")$l����O�-�:?��mN�mh��\E/����J��OБ��\���{4����nc��qX��E;�h�9@(����Y��p���x+�v�A�H���b�h�F���p�t��z-z_�B��٢���o�RD�� �zD6�Ö�-��\(����*�~���W�<��]�'�+T<d���OZ�?�h�G��˃v�6)`S&�6�ٱ�Մ W��-�+B
q/�m�&*Uꦦ �'i���EI$���� �`g�4�g1'�KL[^M�9QQgd�8�Ϟ���u 쓹�j���?� �[K���� u�O�̺4a^����$�Y�&w�D@بt����@�+jn"�̭I�QUG~!��1��8Y�Ē,�I�Z�����7��5�"
);r8�C^����{��j�j�������r���4��� �����y%ʥ���xk��XlxVHYEB     400      f0>!q���j��y��:&70��;�\+�wmO� �@�0:[Ұ \c��'~�̅'M����DIn.vr���w'�"n�j�niA&�����S�g�D+H;8����w�$��r�h}P�|���TV4S�Z��1����o���������4��$�S��ԋ_7�y$N��1qb]C������|-�j��d�G	h��M�/e��@�:0��"��#�D
p�^����hXlxVHYEB     400     150`�>�?q���R�!�{�D������X�׷��+�T�#^#���+�Ÿ��g�uM�����Ղ�1W���WV�.��z�}��� >�2fdl������w�I.�I����cV7�ق��J�B��0�l5�.�z�2�Q�e^��� Wr�g�00��t�-�r�&��j��G/m��C�|��d$؜�>�279�'��� a�A�0E�4���&�}iw�-�)w��`@�����g��A�w���w|H�naI]Y�O��֒N��n\��Tɝ�6s/�|��#�Z���No ����	/�~!ǧ�̔�� �Up�i���I�U��Z�yb�XlxVHYEB     400     170�"�^�K@)/�1/UWR܅܉{z��p�� |`���!>���zI�'e��oR��b;�4���,%u�mԪ�T�?-���7)ј�踎�
V��dr�=��ſ����@*C9
b߉��jL��'忷��=5z$����Y�D��̱�n���q^�N��ōs�څ��!u�D5��J�R^_�~���M%�t�^�vv����u��c1���K��^��>���4�g�Q[� p��J%>k�z W	jT��A������O��W��]����Y���ߘuq��E��Dc�ps=l8¥���Vй#���F�tP��'�ݑ�>s1XiI�zӫ-��0��'�<�^��XV*�N	:�V���0��-�XlxVHYEB     400     160�������f&������Y2�k��S�.'J�l��*����-�#�+�@_�#O��⠷rfUX���%���KN,�����>x���t�˼*H��(<�C�N����ܘa��,}��n��9(���P�����?N��q�y��!�̇b���������336d����5�(K�X��*�i�yً�޾���Aة��C�l9Z�a��@�:]���e^�	8�T��-��Nhk�K6vV@�@/M�[,PGnm6ϰj�M�L�+.�j���	�8���lm���"lo�>�,e�RHo;�y8��ϋ��BY��kR����(�g��EHe^����G.��a� �����h�C�PXlxVHYEB     400     180�x�{�eps0:������b�9�ﯬI`cMy$��M���>H 1.�6��7��ϧo�x����ڶ���[Y���u��O�8���jC��3t��%�\̓�� ͮ���9��j�蘻�{ĸ���{v�?�1�Y���SF�n�\�Y�	i)��
�6�sN����d-�b��ދ�p9����.�
I1L]�i1So=��ȃB|Ԙ,�?�|�5U�<r������p�W�����u/��Y;b.�Ͱ��;��
��K���j��l"�A�?[F3/����/f�Й�AP��X�W �<Ju�zL���gv�$�����L.?����N��dLj�=������#�Dv��_��뱧�,ɖh����}����˚XlxVHYEB     369     180	���i��haJ����gC1� �B��_�r�Dp;��q�|w۱��%�l�k7fˉI�P/."ox��J�/��XxK�"0�"N!X�E�����1��u�Ds����+�B�S�`��&аq˚���RH��	�1Ώ�����y8�(&�#२����1�:�c-���1��=�;<z�~b��J�>S� '���e�c_��������~��j:����y���v�Ĵ�ŵ��E6G�#���=��#�ww4Z����L,�ֳۻ��"����ŭ��^3��ոÎ i�SVM�;mڱu\t�8��:��>gqOlzd�~��:�#2�t��#��z�(���RY.�d�wI�����\��'_ͧ�d�����=�ڿk�'�Jխ�:e?�Y 