XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����1���/��|o�:��ޗ /p���N6�=�*�t)n���7p_o�!P�P!��f��.��������2�*j��A0jS�Ir��嫠�Y0/���=D@�j�o��*�l4��ə
��!p?9ѓ�7�aF��5h���9 �"�_�6 ��"1~�_���?� �6}�r�ڥ�?x-wa4x��L�J'�(sai�����`�jݮ��b�Ğ�I,׹���Ƀ����5߅���腛����S�M��j��gE��d�����R������9Ue!).�[��%af���B~qx���~ē3���Uo��Bh`��AF8?�~���DG���[���/K4���\������Xݳ+�D+o�5���*�0�J�{��T���Ǘ�[C�`C�%��ݼI���~Ut8rz��7�_OM__8�*+�`�|��k�/���jHi��)��*��0�����۫n�6���!��w�)��
\	^���\%���t_�0S���h����ݑi�d��R]�eXw /5Gǝ�?w�y֓�=���G�9�e]�qA��x����.��V���ɭ��=��]e�����wޥ.e�l�#�_By�o�(���l��u�^nUͷ�'�Oqb�<|��6� �o�ڻ\��$q�t��
�೦P!�vB#~-�O&���f�(����il
+I-�z�B�n����pW��Ko����-յ�zƜ����Ŧ}!���K)����F;Ro��O�ջ	2XlxVHYEB     400     1a0�k��U���?����!d�ބ۔�5!WD�}S�+�j7c=�˟�5k�3V=u�����x������揰`(�J��lp<0Ut��
��x�,U�a����_Ҙ�e���b��i��J�z���P1���[�kv���O��r�Բ����vs
j�n+�@�:ɛ	q�m~�ݰ���^ZH�AФ�`bi>K~,�L�q\�ߑ%zf7IoߗE���3d��D�o_�A��V��JG�#���E�gs	�,�
�6$Vc�>�ݚ�b�`���$ ��{����rM1�oʞ4i��կ��~�Tآ(�6�X�s���e�1��[_r��y��^���,�g��1�b�Ci���Cci��g5$��cL/�b�7>i��9i6�&ݗ���`�w^\>m�XlxVHYEB     400     150y���23�O1�8	��4L-��K����2a2�q�_��� �w�I�/D�$Ե8Y)T�������sWV�՗�2�+@�'�̣�aT�V��\Ǌ�ƔC7�=D�����������r3�J[4
�M0@d���]��zY+��5K��i�۳?�T��q{����}{�]�������?��!H��,�OK�P�<��#[�LB�F0�ޅvH���D����/���kDK�m�D��L�Y����`���](�Wh��N��T����p:a���"��U�(��L����!v���;��ۏW)��o\l���,��h��j,�)$Qh�D~��[XlxVHYEB     400     1900u���t�����h�w R0=IV�Ռ�^�&�ez�����|s�4��q<y:G�8�Lf$�/x�������!���/򇨵	x�Γc
3uF��$��Y)l��ꔽ� ��x�����mbK���D[^�������m�{�����R�1�?��]�{}��$G�G��o����u`H_���;���`����0j�1�w\����)|_h���¬����S��T�'�1�V�E+RY�>-cO}I�i���ܹ�]m�^<7Tbp�W��b�Y(��>�H-y����~Ѽ�56c�X��_�,������������ś
�%��� E�tiQ�w y#���N�nv��!���i�E{�K�{-�7
Wc���� ݱq)�QD0���|.�F]�n� n��\��XlxVHYEB     400      f0��bM�M��[��*�8An�_����Hɗ���� ����2�Ѐ{���=��?�@�*=9���>��B8�*���?r�j|w�;���4�?`���rx�9E� �.\�	���pѠ�*�;Xue���o(8�l���C���EW#XM��&��C'�SC�1��õBz���<1ܘ䭘,���� -��t����C������A�y������}��k]��`�S����P��,�XlxVHYEB     400     120?�6<��t#�n��p=ͷ�����AMՍ%�8q��#��SvB�B_R@���[���Kd�4 ��,E��b����� ,�QC�F��w��#=*�҉
l������a���#	_Pv"��3ī'�_O�F�*e;�|~-u�X[�,��(�+kݬ�w9%3�9�Zb��p����w�X�n(�k6Я���W�`� C�����Cy�^vL��٠�tψ���z=�=5��ry�,S�D��ǂ�=�C��ʁj�l��T������g�ի~���XlxVHYEB     400     150|äݢ+�Ҩ;�{���Pm�%/��	�,�\�x,�45+�c"h����AQB��MG|��2�"�o����<�_Lb{m!#4%ha��r�Ų>X����D��8r���/h��xD[���^��4~M��Lv��w�n�D�cc�hM�`-Ä��G2$E��o���g:��'�i,��z_�4������-\�P��߇.95�l_SM����p������!�U��=�

RX�@7?\/ж��_�'ՙDr�[�zN����z�Id�c���?qt�,�;g�f�됼я�qY����,�|��|��"��0�.=���6��a?�XlxVHYEB      f3      70�U������8a<����^A��%<��2�m,�IJe��|��a2�Y���5+џ�Q(��+�\�!���Dڛd�.B&�b��C'�#}���j	����HBD�(O��yu�4�