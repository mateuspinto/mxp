XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���-5���A�竤Yϓ�c!�z��K�tH���t���B��\�jӳbǧ��"k }��$yl䯫)F߷l��x}6#P8E�����@�O��;�"B՜��01�q`�x#eT^X7]Y��G��U{x���8����( ��~�S�W�[�B=��d��^2g&yY�5�O�JҤ���Zv�O�Y�A�-[�hc0�L����9̇o{�?9Ir��=GQ(����b-8�C/W����3J���~�ғ�JX�%���h��s@���@+�7��-��KN��8�-�J�R�"�o�>E��n��y���"��&2�%��\A@�e�.����`k^�×(�'�4MA2����R����$˾�k�z+p�'�Wz���-��.:Z&��EIW���-�	�g��mV��ƛ|LZZ�~6���eC�����"~"KlH�#*��e�A��d�e��:6K��u= n���%����{�|�oBP_��$��ɹى��-����K��S��G#԰�y�^w�3�ȹ�pi�r�4��%.F\�
���&�t� �����U��p�w��t%��t/D��yxѽu<�j=��Z:�t'���@㩐gS�Ӱ����o����D��õ�9ű�'�BR��B{�?�`� ��sNn�˵"J��q�����`�#1L�Zq����1��.$���!T���:��0F���d �B 4}��ר;3Ì�����1Z����F��c�U�x�|����e���j����obEB�3XlxVHYEB     400     1a0��������)�TS.{2~��w�I�0���/l
6~����B'7��_.��Ok�Z�̛QR�xT t(�٣7cC��*A�� ���%��8�<`/�k����W&��kZ$��rc
ce��|�o0���%�""}|D�N�HU�$(u�b!tB��!��ҵ��ӿ.��X��@w�&��>����:��G�]ϐ�x
�� W�ķ.�T��f�������.���.Bvw�*�ݷ�����ɚ�/u�)�#,5�0����ӕ��ﻂq�@�\qU��
����#��LQI���e�s����M#њ/����p�W�p��nq_�M�����y&as���1�ښ���S�*�	���N�/Gb�L�*\\F�EԦ���\�'�0���7���N6$(�Q�8y�,i$�V�c��XlxVHYEB     400     1b0z:i���6��N���r(yО"V|<�<��F_�f���`��6�$����/r	>��U�t�Hg�IhGH3��F��M�1�s���j��5�q[YTil|��u+�#e�i%L���r�[��Ψ�����z��5�BF����(�s*��)���\u���2h��
�9b$���8Y(��st?Y�r?��N^����F�ZFĩ��/Pw��I����촹7:?�/���Jf�W�kc�d6E��G��y�t�Gέ�kվpGn���8%�CiNm]ifG�"�0�Q�]��K;����DB�}�eĺ:7�|kPzK|*�E�����M˲u��wZ���A�pel�5��Z-�a��Ғ�I�� �a�ZLx*��s���qs7u��z"-��O!
���dP~�E7ClhrC\���Al���J��`���}�KKXlxVHYEB     3f5     130�/�=�H�$�|���3������FZ/��L؝����=]QDN����<�~Z�v���$���V���5DJC�jᙧ��qꔅ�9�=��@3���I��n�҈AٲB�H���>=z�8&��ݠ�z>�Fr.���g��΢fo��O��ݢVE�MHσ����q�f'���hT�:Z����3AC����L&�3�e|olx8�2لR��{�:����[�]F���������_מs����-�;�I�=;^{�2p����`sK�"��ZN#����w�m5�S�'�O���