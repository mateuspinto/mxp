��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l�����ǎf�@�}͚�|ET��xW�(����2u�y_�XdN�2��`�&76����7�1���?��s�:��;�R>^WΓ��%0��})��6�3'�A�pv���b&�*%�r�{�����C���M���5��w�T���a��Cr;_�,;�W�Z�ӈw!*��T��*'���!L0��ܠ��&ШQ ������譵�qQ��.h��d����a�	k���>Tc���l%�p���/���p�C�^��� �~��	���4��h���D����SI틣��r�\��#����L�S]<U�;�
��0: ��O]���iVyX�ar��t�g�䢾����?��5��٨�2 ����V�R����
�T,���\��]���K�9�?�I��	�V�v.S��B`k��L�6�g;}ke2��������bU���pR��u�ԥe�+��cD�rl����^!zx��*�c�l�֪|�}x[� S$%Fx�(f*k/F�ϼ}wɜ�	���` �Q����\�%������u��T��j+M]�#������>�Z-Q��g �kx%��^鏛o��᣹�Y����4�\(Q��֪�W�q�mV����3ן������<\\�ޘ֝ڔ-ׇG�NI
��)��v&p��/���H�MO�7Ӌ"���5D���c?�W[�AI�7�>���V�m)L �j����W�lڼm{�����TD��X	˩s�-�Ϲ�,4Pk��bn��$eQ��m���s�\G���a��i�9u6�=D��F9��G�+- �H}H�/��6ju ���H�1�@�(����تx�l���݋�.y�1�=���n�BMbG*���6f��W?UOe9�]>�`:1� 
<w�_�a�Ta�$՝��f�2�BX'�O��_N֢dO�Ō��kC�����iE�|�uO+�N<DQ`���P:�59oG��[��+uYO���ku,�u��M�ОV��ٰ_� ��G�����^0*��o�:q���
zIJ%~�Xܖ��K�v���*/Q!�<���ag�0�k�<�}U�S�ӊ�ru� ��kG�[���x7cZi�U��Uw��6�{�\���NV��UH��F�I��+d�u��`��Y�,�쩰���惵:���@v��ͯ�'��s��:�����T+�v�5��v9��%(҈���wKD�f�`ol��k^(��� �xD"��ЀQ{<@����f��w��k|f���F��Q��/�����F�f~�A�OYA0�3|��y������c����S��lg��U�'�V�;��T!���r�q�$�������$����6�D�T�4����/*ҺRԶ7a�,,Y��{[:{��akB����!z�O�ujXY����	��q��s��o��s��"sA��E�~��]������lĊh�#�Dx�iS5�Y���t��X�j!�z���Z�����?/���d��2�` �!z3��F7�"hT���B-fW��s�����5�-=�}��օe�_�Y2��zQdY�5\��/��?N2|��IA��zi�t�f������D�3��@e�E�Ɠ�)Íf�DT�x��̉ݓ��v*!v ĬJ�B�V�&�x,����0�[Z�	�`鈁#�:R��o�(�K���n1�n�HM�cc3��w�B�@�!sU%��8���#���@�~Ш��;�r����A��L���2�r��Z|C�зM6�mu��ͻ������s���#f$��c�>T?%�^�^�ɘ>9 ��+j�h�o�&�Y��Q���le6�q�[�A�w���ٌ2��dP��Y���������:!����F���W:�2��O �c� ��c��i�-��  ش�2q��#^�v��ؗ������z���*���R�r8�E��u����y����'tbn@�%�d��Ø��D�����=��.o�?m�z(�	)�b�<-�N��k����ؾVbmR^h�3�'P4�B%)�dŘ��W� �M�l�9)�4D"|�v
,��M�g:�5`�Z��r ����U��Dƫ������r$�� ��h������.�%�	�l�@���G`y�pΧ�pH��cJJQd 4*pk��,��:������`��Un!q,�CRտ�\JRi�S'��΍����A©j~��ö.<7&ϗ��\Ź�T��C���sC�v��4GC�QҡȪ7�����q��3y����-I ��D��J�
S��w�V��m�w��|��s7��d��p8��s���5yf�?�C�m�&��}K�x�=��*�:s8�&�EУ3�W����{�����Ԗ�$�g8.a��g%k�U���R;>���κ�ҟ�M�G�cuK�]}P�j�U��ZIN�	��7���ɦ��~ Tpe~n2^|3 -��i�:I�E8H?7�@߄��P�!4��pv�o��x�;:�b�_���Hlk+�	���[)�c�:�|�qP�[��cY�Zp�2=�@A@N{�!*1-leH�Pj1�=�7$� �f���+�.v�U�瞙��TrRV�,3��C��N��[0Pf0Ы=���L��m��dOa�7��k�L�x.1��hs��[f������?*��������ިs�I��BvyY.�ҽ�H�;�r�W��^:
���������>:��V�n���}�0�kgt#W|R ���t�����G��%�֧��0^p/a%|�.�0L�����#x��NrVi�MG�)I�>aI��%�����.`�l]��5L���M�F[��w�wZ����U�-2~_��ϒ�W϶�,���HY�̑����Do���)����N~2���q�HV��/�ОU񍂪\�C�'�	��m��*��D;i����w�� k�$��(��N�}�X68}������N�棏*X�P�ѭ7�a٬DᏭ�/l�������B���k�i��v�#��ѾFJK��İ��i�����#J�v�?$�����$$��7`��JD�l�t *��CD��>nulu0M�c��a��<d��/u��QGltd��k��n��>��u���c{k�0s�S�5���a]��X�Vn���"�*�_���EΧm`J������5�M&��{=���/��dD5d��mğ���m� �����x��m#2�wZy{E�E\�S��r)X=��
�����-1�0���1���<��#CY���l�i�%���A��84���M�m���V��������/U�%��K��@(�϶���V�:lkݖ�ZhW �����b��QIt5�`�֔rC�˨B� 6�
�@�t&#[q.���m�M}2�^Z)I!��)<���ql��H0v�Wn!�)DYJ����Cv%:�m�r^�C�0Z���YU�
��{ZP65OA@9w��v�bh� "N.�3����7�O IiJ���Y��3>r�y��#��l�� �x��jj��Ev.W�k ��{'Z���\a�E3ս��)�Y
���� ���zK\���X	�,mI��/N�VjA������Վo���p�G�(��uDVHX�l�Ɩ N�/�i,�&�w�m�p��z6���Oڳmbr�Kh�_j�V��)i���F	��7���z\̨8F<.�p���<�/Mj��:[�J��Zb����y�AaZrR/\��<�ޓ��L�e\l���䷽��k���U`��|Y�˔���
��,� ��]Af������b㡤7��Ř>��j��SZ&�'�֮w�~��������.��V����~Ў��� n� ���Ai�q>wLH��X&^�A˳7	�}�*l�O ��@��Re���|�ʁ���w�����S�04y�b��*���O����6���.c���F�&�+d�y����G����%���;��	 .��	��"C�=Էf`���!�Η�di�����hE�vo�bK0�h��IRcss{���1#|݁�I�O�z^�Y�4�B�Eسغ�&�9������_�k{�c�>@����O���](U�u=S�o������5�.^vX"x׺\^�-������[�5S��>K�oR�_����vX?b	hRXۮF|����<���:��0�����I#���I�-��0������lAq�js���4V�����=��� . r?�l�D=`T�@cХ$��0�p4N�M6�ǑՌ,W�l7����{�ݚN+�r����� �;T���:�	�^�q<%<$�.��7{�ZGhT�$ƕ�<-Զ�ܭG��R���YJ�Ȟ��`QP�G��/^����Ƭ4�����Ze�z<�<T,Z�x
n�C����B�,��󉋿��c	`h��[���.�����s^�L��@�k����k���Jo�=x[ʟ���-��0r��@�>"ԣ2�G�b_8>��@��Eh�u�0�d0�&g����o ���Yڲ��H�T�Z练%V+�nn"E�eq�e�6��"��'�V��=�2�I�J2멉���ⁱ@HE�y�n#��z�s���)���X����a�wd-�^l��W�jɴ�u]�d�{����ua�˕in�h�2>L���t'J�`	h��f� ���`��'8�8q�g�s|�G�?E	�		
zo��>T�$�iO�^F�O������	�(��%�v��q�2�i� �.�K]����3�&�t�4>���$P�俧�R�m܍�$���6���������a�N-AdI'mA�oXQ �):?g/bZ��y��9�����p��L4z`� 8\y� �O���O�-r.f�ݮ>Tu��rCuXn|bIP���2�f�L�[�<�VSt}�N
اS���Ԩ�3�s�82���xU[�.ľE�v�+'BT�2hVG+ؓ7�Č�ɸp9�pr�M���J�����H-�c��߀xcHU+b��]A����G�KHA��}��VO��g�� DB	��/Jx�{��q�6��k����o>�U����U:t#�H�cQ��)��2�NPިm� D�C�(
��k	w���>R���d���ACJ�۟����O0���_ElPL[�g|��(z"#D����ct�E�h�X�4��K2�s�<.?��$��0������<�5�&�l!>vp��5��L�|��@by����vX���OY_�Ţ���v_w�"������c9� ���v����Y.9�3K��Œ�,weS����R-�<����
�K�}��W�ox��j�������h;�L�i�p�X@_[Zi$I%�}�l�W��uL_w(��������?�R��y�V��"�m饐mWӝ9R����>�����'��E�������4�*l�:m�O"&i8ze��y=k,ת�`��v�����68�S_V�~=8�z{'>��o:�֭T�ׯw�I�ֲ��YGt�9��e���4��B"Ҟ�8
0~C_�p]��]H����]���"(F�V2u��df>�A��N�\�a�Q����4��	��	��ɏ��wt-�C
�)#�k�ʢ�nx(s������=J�Bj����[����>(�;�� Z��C��-�����2E`$�3�Ǥ���y�˕)����¸a��Y9V͝3�#��Q&�DX�����p[eg;��c��
/�D�rP@a���PA��,3��f��G�:\\�z�Pc;7��=h��p{:$V�)}S8{v�<����,�U�hb�p*@9��L�|*�6=9e�"tp)�v%�y8O���@��ѷ8� v9��$��J�_�j���c�-���J=�h��ߵ��{^�r� �[���]6.�9�?�X��EЙ�c�芋^;�a(�q�����Ɂ����_(��:*���o�W�a�e�<���B�j��h6*����lud1(����}�j�7\dcj��B�͘�6�weSx��M�	��$.�Uރeq�y��X�I�-v��c��t��� ������Hˍ2�a�D��Y��kc;����*y�m�6�_�Ϫ���i��5���jv_�e$7�;y	�U�P�DX��d����s��$��_$M�MF���ɧJ���?Є_$qYY��zj�\��҇���ݠ����dHZ�a��ܝ=�����{Rh��$�aAYW�k�P��&�~Zsw?�52�n��z<�h =�l.�li��C�
���|'h�m��l$����V҇�yBH������(�dI�8���?7۸]�<
���Y��v���i�9�%����cJ�*M`�D%<~�Y
�K"
���з�N7�}�,�P�%��E1��J#d�ୖ�c�+�u� �WѱI�� z\>��nt�g>vh��/�~6�<f�#b�!�2��zma���Iu��2-����m>�9!~���8B��5V'O"���gr5�f��@�6����G�J�T�N��>y{���D��f_�B'��^c[i��֍��9��,4)�ퟟ� ��x�y�I�^�.{Ȏ�`�~ɓ���ܫ��T�3�,ܠ ��{�(��;>+�� ���e�5�g�B� @`��6�D|]6^C��A{sWn�}��c�y�g����@�Μ�,�/qN�*-vܰc.�:�E4Ets�W�*�B]I=#b��k�?��*�P��1�cV�h�<��n�pEQKg���w�6˗�
7p����GDdX���j�ը%=��˃�t�2+Tҿ!G�j@�����c)[l32uV)[��,:2�X*�� ���:n
���<��2[�?~ߡb:�����V��	��$ˇ�w,�o+pO`)&�-�Ų�s3r�
<�T���	x�:�~�)XY�?+�X��O�*ZRf�x����v��#R(-&��6�Q���ii����[����ɹU�G	�4�%ew*�x���4G�x�6�;�q"�U1t���Ӣ���9 ���L���
V�ѥ	X _b/�f$�'�k@=xM����Ͱ9�E���b����S�8,��R�t�>��FV!3�\x�Q��6�&���D	��t�s���دT�b����ѯaVB��(�J��m(#��]��ٓ���"�f�D/��f���x��VۅLZ�^:[bxIH̨��ހ�0Y���P�pP[�-����G(~|�U�V"�3+���O��	Ԙ�f��Z�\��tAJ���Bꙧ�G2�h���S3�B�}�J�V�ju��g�<�R�Clߩ�w�7�c=�u篌�v�_�����t�:��)�O���O̜&�;	 ���^��m�3��HTp�o�g���ӷL��5*�7<ʋ&���U�*���.�&���C�JBmà_�0#V�,�)�`R�38���f]$� ������}2Įwaw�@��$J�讽p�^��LDpw4�n�N�֞Q�^y$�θZ����%<�����a��Wp}�`�i0�C� ���ˀsGj���>h�mZ����!K �|�uMqc��2πR�(�"#�l�f_C� �,@�k�5���T�ە�h{�i@���u4�C��p-]�V~� ��vyi�J�h�������d��������@�}I��x��Y�̗<G�����L����w�Gz��l�����K��m��J"����!|O����`���AB���4��l���#��+ W#���W�\6o�}ɪ�J��?���L랗X�g�O@m���XJ��!����\H���t��������[&�!�^�:t �/���� ��7B�x�������c+V� �8V�Gu H��	UWl[�R&�꤈ j����.@I[��qX��û�c�;��T��=�(xjg-�}��xf����%�T�9��]6�#P._:o�)��Y{���U��m��ORF�����"T7o�롗?��Y�k�c)��]8��4C5CL��B˱x�� 5�������C��6L`C`�U�D��=~O~Q�d��I�>�Sb�͂ںOy�lݿ去_S|����Z�a:������T
{���qSo?^]��7h+�K�b�RQ�l4���7<�O�����3�SD�kuEsxю3��:e�>FFM�'}d&�;<I~a�ߪ�f[���S"�I����`����<D�c��bo2�?w�͢Ac�gL�x��=s�Q��(�4�U�z�;�I��VvJ+��YǤ�{�eEZ�G�>eOVY�Q<������U��#��|�cY�3g=�i{ZC+����bq8��BMO�:;����q�5x�I=J��#�^TiF�[��	�9��dI�/˵p��-^.d4����c���ԑlaa 6���?C�k�̪��g���%4H1�������J��q~0��ʾbmY�5��
I���
���.tRK&�������};.��EV�ᦝ¤��ST[�D�C��
O�#�����ѝ������p��%&����4$���#:h�Re8�*�m
+�_$RO���[��U,���T� ���C����Af���S5�_S*~���`�=�{�B��p�M�(�]Y�E$QD���z�2"p��^�EP��L�Y?��H���r���h��N����}�ʧ��I%�M����"Jq�O���<�N"���?G��{��z?���TRֆ���=R�I�ӿ�A�������ڳ���O�*�������2^�!��碒��5rƮ���GV���B�(o�l�R�+j�$1Hp�٫4���M�ķ{o��N/��k���La��o�[�G��䗛ߎѤP?.p�+���#��Z�]t�@w?�d^�2����L�풐m�dki���
Q-vh�Q�bP�AM�/`��W���]��թV݆ ��ߍA��:u�(y�Q���@ ����sJC^ןu~��y<�0��p��d4�-L}q���>�%�2��_X������1�P���@�!�W�
	�f]���xBBCq�2�0��R[e��yW��"��G[l>�&"��}v�K�譯R2Q
�8�p~�@���]U�����-Q�"�8�HK͔^Բ-�S���I���Rq/dh��Q��.����u\.ZO*^+<��%t 
��{�oQNo���v�벃^9b�a�Z8}���t�ݮ=�|N!�k��˧e�ա��׫f�|�08�����Q<c\���+ڃb�F��i�<��XQ��0 �3���j��w�im��{D�����2y�,x-_A_a�j�Q���H5��v#�=n����!҈0q��uQp&�\U��L��Z�[��(�.�a���=��,SA�J�hŭYo�2�Y����><�����7�=�����%��{_�|^���~�5�fj��
SG��{Y��H�ڼ���!�ś��[r�и�V{o�d;s��_���N��6 ���k.���E���YTّ�z3�l`��t�d1o^_�`�Gy����D�dyf�p� g�hyvܕ�~b��֚��y9�����ed� ��+�Hs����D�	�,�^���z`�������4��Ŵ�+�/�KZt����A+�J9ro�$H�$���Ӏ�"v�sztk*�=K�m"99����0r{U"���!2^��e�<�~�%5{7�~w$=⢧#~*��k:�zE�'��C�V5���g��O�Fת\0%�M���H�}�����a��
���Y�˵Ǐ�J�f�b�k��:؋��r�fK'a��l^n�#o?����
 V�t[L�
����TV�Yv�F:��9N%�����W�E���[p��չY	�N10�r�B�hh&�p�sچ����-�&Q�H.��1��jy%���\�q�W��@h�.k�~���u�Ӌ�[z��MO�h��+����ၳ���W��	8�x�X`��3��e⫙!���4�����J�
U�(wFs)#� �%[J�@`��{�
{|*<ͣ˄�3�dhřTu5��сlU��	� ���W���1b���Ou�^4a��l��V���B�@�E�}�:F���rd��H���T:�R�б����HH�v���_�sS�H�?��x@ǜ�ay��/P�]�R(]���+������V.+�S�S���'S[<r�	׶�k/ϑA9������h���B��.��b{��`�0~����6�"�vT#RO� k��Y�l�d��f[*��N�h��{�i+ێ����}�W���V� �g�!�
�����PSN�U�9�Zo�4��W��v���k�a���9٬Pz@%]l�W���b�%�7�0HDn� �q���^�ie�cn} %�L�@Tc���N�G�@`�e��zsP�`6��q5yhY�GT}gLg�g�]�l��Ԇ#㥻�].)��?ᇽ{���� qqbg �Ux���<;��E:-C��RQx�u#"��[F:���8�< �#Z�2�����H�w.E�r��k|��׬O�ԥz�w�r�C��o�DuE�^9�n�C�?�%�BC�U4��YܝgG�g!ߢ~���$Z��z����KѺ�9Ҁ3� �(2��C݇�O��˫
����v�ׂ<�D�M���
�Vvr;B�oʇ�-1ݬ��.R���]K�b\_�.����Ȩ�R�~�̷8��Ǡ���_M��;�_kF	��^���'ۀ���j��;7�$8mR8��,w��	����E��Kc���_pٯ53�3x=�����H]�^�+��A�J���l*o��������j���׈��M�r�Ѡe}����s+�.�]l)뺪���=���Ru�q�$vw/�p~��,چ)"	J�-���Ia/��;�1C��S����qĬi�}�-�/����Q���<R�!��I�S������=Ϳ��z����蔯yݷ�����y�����@z*��9�b�*R�2������j�*�n��wx�,G�;�g%][;��UA�ư�'�JÎ�b�Gv�6��ڢ�������Ւ��ւ0&�~�b��H?
�*pە+�p���뤚R<�Z�ɝΑLWn ���6)�)捛T7�u�!�.pQj3��� ����Ѯ�Gc��N��(9�ʲ��O�e�� \9��`�
l�-U1w�|y2�N|cΗ��=p���1$����3s!k�����hTt*;���{A�`q�p�����"�T�{��F�^^�yn���w�)���`G�4oo�K鞟B��ڢ���(�#8=�9�BJ$�S�@ܝ,"U������ �ށ�E0���_�����+���}�34��PL���!�D��/!��*������\��D���ںm%���J���y�"������_� ��]=Z�=C��vUy-։�4WJūo̟rVĶ�Q�NZ"!���L�Ǐ��Q5%L2�Y����L�k��k�7N�Ҭ��}�N�I6�/��=�1i���$w7�m�s0��I���S@���*��gO�����v3Ξ��d��