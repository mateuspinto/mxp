`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 50720)
`protect data_block
xzspY9Sk/DaSxt5jYlWzSujEYqfLeJ2DYuHNbLB9uszfy7obhmLAhmLY+FQeNvQrJCWUQHZDJl4r
pa7+o0zU8asWNqcq1CsBdxyEkfPuyrq+UF6HwUL9kDye3Im0D5NYLgkVRSXZ8fJxclP+Q/HoMAgr
6OJHVnrRuwzQFl6cm2Kxs9eWk4J+U2h7k+UMIJgo75T9I/aiB2uEiuhefn+l98riN0dTlqnVbiWV
tIwaY8Js/78h5h4sotV3at/xodl6rrBdVZNoD3eMoCYgTW+22rUR3wHnH/ta3R/XVHjHhVjRY83V
24N1uIDYPZjuYNYtRYWaK9uGkWwUiUMzWGDxXSt26x3oBAyaitVwkVfGX1RM30Jg86IFZ4ZvMk51
HgeAD82oA8s4B8VZyc2Y/RnvKwBKET5/mgNeYK5mQhWwKlIyuiC0N5ILKjVcyh/25NPf+tz4+XYk
2/Fu6nrVPYFlaX++VCpHwrT9hi+mBZNnyyyAsHb1pW5lBha/jaVNfe2KoFpVaXNetYJFJ4WcRaPQ
Qai0rEbp2LjGUk+UxOHWuEmcJt7Vp//Q4wU7tV1enVk5AZM7PPEa5dXrjXq/CkDqmuLv6G2UEkPV
79JmHKoFTMsA6tHtskmTOERVpfGjspz7QFRu9t7pGMifZV+x0VSaXGzlHM4x8iH/oi5JRc4wvmZN
MqBmP/VIvIwT7zgSHJiR8PuS6Byi+q0dUUNwDmeHMwtcjy1OhmgnznlwahEOwWOV1K+OXhSkjVje
Oqd2/s7/ZGS6pCr6ohBIHao7jxBsHZjgwXQWyeqvpgCTlFOU2oSE2qMZAwjCASfsKtI1NECVhfQD
ggifHccCZV6Jlli9D4yuZnPBlBELZuiFfH37puUmHi5CyZcsVBZOkHW6dINo/0VX1LIAnh0SuU3g
poekX78BJKMNJbvmr7W5jnzSeF4DJoMLzly++BDt062vv2FuVlYrJDsPx/brn6jypM0kMkgzzHIT
YTFT7J6MKHcbO99sBwNDNEKaA9HnK6fXoHHIGTpCRYJPNytG1buitJt+Tvb7RKKndud3W98c0TCF
rhdm2YcvzSQFv0HbkiD71USR4glCPtupeqW1Zh10CKTsssHULxtW8414n1e/M8NVRJF++YHVzfFn
75ziETvUweLwzH3c/E7IVm83bOCpOpsPE7GtPEku5kFRk1Ikgg/bG3XHBaC/g0sjsom6tyKj4f1n
t9y1uf2Y+WxrZHAeBUuuTigoSY76IaXCtpN5N2wVjoUjkP7KptJbNVWe9mnC6nzGbwkANEbP6S5a
MjPW+Rqt5rORNLqQDR5qjaDY3adFyvsc948oPL6wQBFA8Pxsk6i/OYZ7/RM+wrH1F3eklTKI6WOy
vCUrlohOpES6odpLccoC0AlJIS8BX8aReQlQMCdl6Wj110ibgB1bnwcccHYW9wEzrn25mvPeW+FJ
xf0i6djRxjSokhxoeBLqKwA1bu+qQvFxrtsjGczt+6g/8IAkEjQklT0xvkp6qlBinb7KgGz5HsrH
ixEIr/Dt3WbtHOOzZNxO+fvrjhLmsZCKqq0le0k2IqcWSOeJKYtEapQ4xo1ZALzfEeB/zVhA3Nh0
XdkZlea/l+smugVylFsm5+7m60uyqHHQQ2gcDZgLOt9GhPar8kT/SkB4DdDTPnty8CvvzkjDhx3F
c5jWLj3JlM/DrDuRXNpeLOYnnZs4DUoX2u5l5KvQYaANyHn08afnZgNK4unj1sKH0BUcKWgbvqnE
Gx9vMdf2VcxdjLTJpTKVpHmpi7M2YzDrOiTHzeJaESYB8Qbq9D1gwQBFpgm/mDeyw1+mJPeWGw1p
mObtGrl+a/ab0Rm2u0VWYilojJeBD/zZvJgYNyolDsIiaExsLL5MFZyNNP+rBL09kItp7y/FbMi+
25pPLioj/vZ9KrLXrVTsEvbAQfLyVQf7CCZT/eNq81a2joxz+7fXhOcLiiQGe892EV+0NFpXl4VG
6T43oVxBDh5jF/MwJcqSaQNzOf2gvWdT+7f5QmFRog5qz3xGZYxZeMG/ElxtqVGpSxwm3cVSnI01
q9tG1bd+2BHIsIkt/1TF20hYBZ//u4ebQpUByVReBbjBmtcRohqrl3UTUVvH6bERLej5HdvY0YK7
FgQixIljSDQNOgSFl7HpI7Im02bFxy6jVYlmuQE1Wy9kMpwHFBSEhedBsIa9Q4PkMRyIdHl3q0wm
HZa1AS00DuoqRgUiPatBY2rt2VxtPPIEUr3lTYCfONGtn/qcRZdObegGeJGPPT15BOYbRHIelweD
J/UvIvVJDBheqBi+Bz0miAFIdj61QzVL5ou96nq0KT9bFCmJOj7hb0xXSpVUxcJHynLVx3xNyCo5
ie2fvtNOz+Vqx6zKE0nBqRG/dgzmf85bSSsSpBqlU1fOOjaykTz+aup5F9Whn57e5uagK4Ktt02F
zVb078r+07277w0mU97+gg7dyia0EoYE/30JK+JKD4ORe70r/NJV9oGzEu6d+W/mexZ7vtUD26Vs
snA17S7Xs0zwEfRMIAIOo8LdCTxikioYVMX8xO20oPmlFP7PS3R1MbqkDWi/tCNnL4fGUia1TLDu
aYODPnaqxhbxsbajXN+FaCsBpudUs+OlXuWwA0A4KX+h6dZKVQWOFKoxyo1AeXysAo3+yuGJBrie
mWlLOf3LmVtDsS9gMZZY6+vv/bJ8iVBsiJ0gX9FbfmcfjgGv0EOL9du9BHO6PNmt6I8cXCxcmxLj
K6/v8iR8NCVZgNSvMdYQK3QgQcD9s2heyJGz5eyeiVp45AeEOn7j9LB+wVouhG5cb0CYRURpYcXz
Lym3tKClaYrZrTLD2zF8laJo/Bld1OqhZ9W3zs9FdYjWGfMht69mMEUpmwLN+qogkY3hYIIoXAdM
cD6B7cegSnUtqf977jMg/MxznRfCo8Bw7AnAre+ePdDt38m83981w1dCQJ51lDSwf2pOgLyrvOXy
GoASrlvwlH3ACO6ZZ4joNR1YdHopPJ+7TDtuNHRswDu6SucsZPU/XKtjZrcEVJpwD+Lx9msxBcmD
y2lsJKMqWxCRJlXGkM6XQFCSSltRJTSRmBLIekGTFESJMFO1Vxhed4sXCizVccXYR8jp6hacxKhk
kop9NT56TwTgdtIwt9ls8jjfMO8sL+YGfuqPQxZMlXPiY7gvjuBqmQkk48bFcTExAGpyO1AF1kOq
MK651lBrzIVozv9uK7FMCoexx8ZzcZuIluPPArd3H6Q5YjFYr6ESp0Yh3Mi7q2JGnupDlHoMc0bE
Es4G3bT/EBZZKoptZEJzG8l8jUNjsIu4MPQlAjhbTglz8/xSBr5GpJCrziD8JcELwC2N9U8WbV/p
YQsNqf+WYswV8A/Rc5lN3F/+kPuSh17My1IegTf0OreIUv/943SOhVsPTk32LiaEHHeDTmQQZJDO
mZhL7YvozcKlTIrYnsKyIVvLs6DZCpb29Og6KooR6vVoqr5kxG9LKf7JFcgg/fxT6fxWKSQFvtWQ
QbNfM7iwxwCyqY2wvv8GdqJLKZJHUB8TPxh5lntuOPZ5Qq4Nw2h3QYr5HnDOR5ZaXeMp8BadjWl6
GxdugmwkDOSAzWdOtcQ3fwBgZXioK2R1WA50UdYzKnf27WKgrl9rlz32CRuAlz5IbtsDoJs4rVrH
QVR9xDGxLfaI+jZBIzJ44+FmDoJUe3pDnyIVCypw/LDnVef5Luf7rjVy1go2NbtEcWr/V0/oCpZs
M17lFKub4HhcDtZzzKPKQmst/abVBq8prCYc4jvaVgW3wlLGrySRndgvV5Wtuyif9KmJJVaNI5HR
yRQbBxqb/msRzvZlbHunoUEYcHPkXvZKdOhoeR44sgdtlsvyH2wOjsEwbequUK6PYAjleZaTnd+u
CqUMfT//9WnT2m1tHW8gWluOyYvhrv0lIMHjWMV6d5hUYnebVUGTJVnqA8F09ItapfmxfoASerUG
hktQIXCNa0c0QuIVRf1V7arBKrHalBbVrvmlSyh4ZsOHF/Jc3sYeMKtVWWzTuV9C7FyAw/tSoQ01
Op3nFUIEmrIxLQWWY7/4HM4/1j/54d8/vbePS4H/9jXPTzzfDCc3LN4oPqvGLCNlozFY3rmSQgko
jFkKxWswjcQ2yWndWkg/xCKkeR9hyCbzxOqQW7DJXd/OzvKqv4ENy9+CRQLw4+5bFeqBdpQ084U6
KaimI4JS9ID3TDqbdrmCAsgG9p5taOlP725fc9XPntEpJb6VRDa/u7YW6as5Iax94fglOCyrZvs+
udPCUzVDmkBmIS6JaNI7RMBMBtLyK4Z1JBPQ0mmUCZEbX2aC1LNP5srzJUkBd/omROR5MUmfrzWJ
AfexUgAchYMzKQ92IvMJxualtKaPWDo75SH4KzeQMhOw2KyMhAkpBL4yPW7/Y7ZOXWOgRFp5ZIT5
474cuKXlsOyfQE0tOr9mRdIIDSUK4kn6tQsGlcd0Em3tcxKByCe0rGPaKLn0kTcWif8jmJ3fTJxs
BQQJ9LgTCVTKEs3dCCRMwDG2WZ/KNaP5I88bHzWRb7G27HfgstUeB5FnLnl7n6cOm2j1ohgmrWHS
OT+3EH643u23Ma7K626eK+mVjMgWBH+zPZ5xlYNMqTMrqkc+0EmXyJlIWVFkm+Uzv6xtimTsKc8M
jeh4P87R5jUvwrWWzI8qKjr+3GigKkQTf729+3pUKW1fVU4iz7Z7WeXimvMSPNZc3J3QLzG4chp7
MGXg/D0KIpY4J7CcVVIRjpdIFZUss2cBT7wPpo9u+MIy0sG1aM6s+WyiMhvQp2stntJCVttDMrMY
ojzkQaC+91Df0U20IbOxw1pboYTdYsgljAKA8zPgIGyeSb75bxfNpCJGopfJ3633DW+dCfyrL2fC
OBkEUNd07hpOIkY7Bdlfw8tGaX6ECypj1VUzucjfQELsGei9l86mYLPs+9z5BFXvOfB7IgTRTdNc
+Jl08Ruf1noZsJ36vPEWPwTx91o+OEIk7puS8qdFZXPUqby/n8tbIjghHm5AWfeq4TJnqaFQK77A
U3KYhoAJOJhMZD6GqJ/gwRQ4IoylBMiaFm/6NbEwEWLn02Dy0aXVfclJScGZS/nHz+T7GwKc3+eA
5B45dP9Y0dFcC7X7FD0rdy1XOo+5ROWMutBytRj33lbHQB8km7VLqnmEB9JDcxvobf1X1xQEGCLg
CDd0Gn64/uMgNYDTSwZMTLJ0ZYfVTGa+G+4A1DCzQkhcjEoyBl0nSCZ3vNJJpru1enBYS24LkZvL
MyOu5spUZXU3Qvu20IK/eXYKGJkm2qCYVreKAbr3cjNJmHvt2WItKPuUHLR8+ixmP0o5QnqwnAaE
RgXvccDoh9BLfulVOyvZzOsCkuxNUn4D989QfQpGllCIezbU4iX3DJfj/y4ISBIj0eJsP77YZscI
edwroG4tehhBMxShfrbR/Hp9cH+l35fL7s32XLqoCX3j5C1WWkHep9ZsUAs02k4DiDz3hyU45G6h
nqioT0RWM4eNluu/zOCp5LONBMz7Ht+p37s68+Cqq+N2PSIqfgQhfAFM3/B2o2x5vAWv5fUesQjX
5SUF2SYUFXAqwQBoeV9dvkjBNmBEwekMJezdQOTKAQcVcYjep1oWvgFutLGT1ap3LmFxwv4+n68Y
9KBZaRhy2inES1Sy5f/CmkbLkOEDVpMY9VTAW8/9H391mFCWcUw7Tvhnhd1eaKrz3bru4OxSGwVB
1RuhUOayEvGnRCP6R0AoaiyxpB43ONtjwJFb6YUKfe7Vu5U4x+5RwfvPr5mLdrQJzZsiV1FJ/q3Y
bgOu63xWi75TNjlshN1bbOHt3JHLrRtw2603H7XttMpuMvPt3+p0CCX6E4y4DSc4Fvjyro6eq6YA
mDD97KhWs6U0tA7E+MSXy3rvBE/hmZflTjpGQKQPaLNzhnqC3mKGMDWreL6KUaC1KUG9vUqR4d3S
NVL98/WcTP5zrWpGN5u/LkwPBl24uKxuw9H4MN00nZ3SXus8M8MJuLbIRGBjWR1xE2AuwkMEDw81
2cbPsOgdoalqYMnvKZSdP7j1NHn4D1fQgfjZ3tSbuc/mbBLOTXUjxLT5jsdL4kbVTwJmcnHmNImK
jcmCfs8+Z6IFBlPkeG2fm6TPQ5U2F0EQsjuj0+EQo7cPV8XxztK3XI1h9hXtWIIyroPqpFsyFHSU
maDwNe1FZLNH6FBknrd99Y+48uhAKRmq+O/IQPDO1HSHXjrWMvTN2pBZ3xxKthrrvGUZoBTE617m
W79OCeKF3qq5PvDxT1a7MePAILmNzsliPp9sTmYOTdwFzI72wBY7XX4xRO9KTpqNUOKONK7Btx07
DCYcDwY9157Z5eRV8WHiP3sblcWJ7L1Y0bo7VIoZCZEt2zKnrCt9Wjb4dPzlxb0HQcZuFAg/IdTZ
SiXrgNXP5UB9TL191Zh/ICtPDK8U5ZMA15ER3wy7qjt2jJAjexlg9sWYkk1kcGjUyjX/oNfZzpFI
XxtHkZs+qpGLaLjUbJjH6e0oLFoQACcIVZA+XjfOF3y3ONP1PLs5/wS/f8MkDAxi1er9M8v9vPZk
t470tK0qpZNDtjQ5y0OY6t2ktJmUtvKZOoLpKd2uFLcYlfX3a6m8HmgrLw3e0Le7IGuvdRe5iVIK
BRqMNU14p5YWaDScxGISAwdcHqKEa37Xbkeog5FVfEd3xfmrVEbl/zm+niy0OelawUgJTye2ilaD
9owrIWlRj9HFOqAmssLcBZA5x8IeqSp98dQfDr4ZbTLfnatgNNjpL+olhgJHCl1b8Mf+40lGB0/T
YIK7a6DMi8tdBj8fEM0ciEAZ0fKfvKypl2mHV5mRA3rVWuwiiEj28VtrOQKufh7TWqwqd/6PYv4y
P+xbfds79Dqbmu3bx6wolaoyIQOKrAt+Mp/HDXIb/iRHZmetITAGjZ+exAFfN1NBoqHkO9mfOxSq
Y9erKZX4xmVkMogLYn0SCMkIxaqhEMjGts7t5ZxTa2JGiQtA8ZQQBL1aOS08OfSPKT5atielUgzi
mn9nTDSeGqKP3PdSRtTl7bEB2fw06sBfsANW831ajHZGFTdNOXOpo8HEmx0B4YjMm24wJ7K3dWsi
cS11jU6BtbRhTxLEAfAuHjKc6lIy3CveX1R1dySiT+VL1k2wnQBTWf9t0oZB6NlTXX3RbUYkJ/GJ
QG3eee4LkYUttO08lkvCKaVOZNa4dPSKL5rl3BnIL05MscnDPqWTZVYE6IB3Ua2THwD2mvGZ9Eps
gXK4s6XrZjypuJvs2ytM0t00NN5ftNb+R2YaS7QpwvhixA5gqWMjSJLlE6gS8dLa2hW8SWuzzg8S
mHaeSuuvws5le9zK1CqeWQy/TKYrWhmX7Qh+Rt5EXWvnF5Oa39hO6ktQUiQL77r0/zbOkqo6iV6s
pm2twAndTRt8lUe/Nu8nQ+ktSMMSukNCSk9MiRUaXiCr6WIR9o35pZicHh4vC1FsHcbOgyZxQdql
XBsIr7gxPFAQDwRGSN69cSuAITJHWT1PJkE22w/0WDSU+6eW3/vugOx70aeQ/u1pjeXczc9TKBLG
UdZkr13CYTIf8HwyvDSrBfBvvinaIOXVFUxfY7oEIogu+kovbgh/pG4H0H3CMBclKCwkd2lQjAcT
sgMAp/VlmswPot5WIKJPwy/HYZ1y/aspv+rVeG47rZSvMYvxerNy7tiT/CZfvs9D16gc8colw7bJ
28hZldApo7TwWmvL2zYOJq5MTY5EiktxkEpwHgbQS6l/T3Rdt7EIuQ/zOhCVA/bwqQcG0AqG8bnA
KKFoaqxvWmlplM41awXVgyO9vIgfTsB+4EfGcfnjkEuVFuwy1AMC5gQnGxCL7AhE/1bLl3Mh2cpo
4ozO/mACuJBSfiAhqHBcsV33Ap6PI3HtXg508AMT1jyJAMyQ9m0jfPmd8J0GPONYXtwOh/N3rQVe
jZaBHmH3T3cWioRR56TaNRLI0W0ADzz7d148g7qk8yvkQBUubvI00BSMThnQIdzvEayeBkt69ltm
wboWLUdoW0u6BAZ+7ykNuzcr8YYnSa5aVMR2U0nlHMJpsnTMooOm7+sIhTa2U4Wchgh5Vv62AjY/
s6DZ5cH2X9K8SbmGji8/PrBFv2kYYXl28p3iCvihogQfmutE+nw17N6mnYWG3IdM+BGglYEo9JRi
cXS9WIr5ODtAEfsEhCQD9yx7lUx3SC9pKiNeNNKj11v3WLFT38ejs1RVHkITYvn85UhvDWtkzxGE
nSzefd2wktRhkY67ML58A+Cy+enf0R7IuVPyy9zR7OCBQN07MmDTE9DF9NBLZQBPaV2c+X0WgoZF
qyGAaPhEMBb63qUk5qPs1m8JwgnvHUExGQbC6RKbIysalN/dX9xz8LQU2EbAplcpTFQ2Tcs5AxNQ
HH2zVS1Razx2WhPSg6a83MjHXMq1vpZyhtV0Do8Cmhiz0uaYDlaMPLKwctkN3zLIp5NBtr92eNYB
muOvp/LEu9n7KIN4ZX+agV0aY20WdK4uRQ51Pnxnm4gimFc06lOiGRxha8pboGnZAO7kAz0n/Zdl
YG78DgXvH8dpDUPpOa/ehwhgINjYOx9LliMPxwnfP2E5GFoSworat2EGN1+6BY8+gE8WAUS5Prks
RosaXjHsMDwGFbmAN8HA4W1alJNE6FJR7dYvXCu6A7xQ4eYx+0JrSWFkfutj9ta1ESw/wjI7Mupn
vCgxJlNEtDAiYriiG0COwbzmE1IH6iXiCjXeerh/PQ2Gi/+0DIjGx5K7b+YeXSR/ik0iWXS+oBOb
zwWIj15uQB8eKegqbI4Qz6PBV9/lTo7YRogjoSZg/jgCSk5OjMq7Y1HC4QyHSTwJj2tjBVozZEWv
Lp5NsHTI0bCgUwJzuMASPDpqgpaU6BGo/iywIlVSjcVUhdgF9DO81MW6Usm5MvixpyBmtOARJmmV
WvuMAv9oGT7/LiirNaCmiOyQSKh1JcKpcxoj+Tr5Tes3q0fMf31a0VVjgxN9Z9J7FSpeKG839bTI
oTCih5dsMfihYGT/7aNU7s0F3ssnz0F9IpbyEKGYhc7+g1PTGLL+FPDC3UDCV3JJZ+flvCFnyy8W
7S+b3KccUrSOUP88/cyFHtS2WRb+JXfKgJ18GyYlI4WQg4Lt3Y621JrnThXT9jgMlHcZIaFYVbyT
WQ++DeVsPhHJipsfLsAbFzKKqX88q9SD865US88ctmeUBzwN7hDuL9Io9ZHdGFQOkMdZpiT7IXA4
ZfFQp3GLR2uIIl+MbUJFC9U4w2Rqybo9ZHuopF7q5ZkRBPNUH/ASWaSsJ4v4GtMzFoimlaFWYYxS
HUZjchIwH0gREvAIfW1kyiDYU8Df1LMxWbviPiB855fRaDQBFcQ4kb7dsZhss30xIYPr+JqHC9Dd
iEmj8pIRl3kzn9hH9cYEoCg5ShKhD2TIXRjtH/FC1EKMG0prMzQdGt1vnvqP5q/p7r46Iyz6m8B+
HSI8ipbUTsV2JngtwLKUNG8lBbTe5ZaqddIy1pRRdApBTbBb+vVznfNVDmdZyv6uCf8QV4mLCaHb
96CNdRddYd2fUsXmE/MV6cr4vTFcSEEFOqMpjZy2TXN419y7ipHsVTQuN9JaiUbn1deP6Lw9w9l4
bveppv+cri1EJdUmLwcB3ztwJiZwSLJSghBXfQkP6dmcYfeVhkHcVX+G+WGx+7yynutEicHEcNbO
lXJ//kt7M2OmvwI4oJ2uH/OUtxBI/BohMwQpLT8z+xE3YWZNE0feC23rIax5xNyLLBRAtVRDxuv1
6K4GDfy9y3Kt4k6ezY1/1q7/g4AbSEa8p4huNyHjPjgV2uYM0p6zaxYh0YSwZDj6nxAmTZ3RtJng
jz5Tu2PDcMvwmilnywP2vJg6X8AX6U28TkkAxnaH2eYWQKbfHcPIEynow88V3X1Ap6+U6vOuZFRP
WjvSZS3Gb71t6Cr8zrHtD1fsFHxA2hanHGCR10hjTffcsJ7zj3AdPx7ARmMQhXDO1ADgt7EG4Z/+
3eDbpxAT43ZYsZhY3btKOnSTnWKmfeAdjFY4zCqJnqAELCcjBOiz4SZEhKIK1BkkYSq/xsYa5k35
jcpiWIP19/bE484EabIvDQKBMHQemWrU3wX8wi9efF5hxsBYqxvonZtCwACVFnxqEyXL6zdEj1bV
9lOqXywkC4ALRdJmdNhRxjjk8L5WOFJoNtdGuTNGvMB8YmhUuT+Kt+unl/uvk4QTokjp5ffXFWAH
ljmTl2AgYcksVVKuR8TQNTMLiPCHzRqBjDdAwlSFwZWxZj0UkklUQfPOo0e9eB5moVhlklyjts0k
dzu+UvxJlzH95PwGa50TbSTUKObpE6birA/3pIoyN/kO1LGl/lAK70vfrfhwE+5pqPzBamM/riQO
dEC2Yim/AAq6JIKergwuBPPMV5kYmufQ7mO6x+Em6/+1bR03sPT10ovGfzzyqYGhHWJc357pCEgZ
xbrHSpYIkN91p6BR1FXrkjPUl/9hZdEj+X0icb9yiqG5HbMC6eBBXHUbFf6zc9dfS+ji26wKeIJs
SRHkECQbmqv9vEtzhWExpbE1hiDG5Qt9SowVFcjskVJH9p6Cvc0fcHXSQOJ9zO1Li54jozN+nxbX
QQ9KUSsDkOYKKwFQUhcxOcLaYSS2vD0az7nbYSmHJlECwmJIMdeR1eW/wJNIXJNzu0ybIBdps+Ed
ZW/WNvkv5CAM3WOuebTW3KdvLcPlP9l2ySTq6v9bKH994YTuvvzqgtRMhs4NknRfo8Ou20q558JS
+sBRpByIMfuPuO3LCqNmNuR1frxg36A7hCl3U6J3Ymhg2HRoerWUr2uGqJ6zH4Gh80a5vMXm9/wA
WPUPr7U/efD/BP7yHN72sxom7ku31ew8T/3s7WwYE8BGZ/0krMrSKc5WuTU1fCANu0K4DcLg7KLG
5/7egf43jsJuJ91dNLYTdcu9ZSD/TnAlwXZootT4eWdnrPOAh/qAzqIe4aWSr8SbElofG5VRONGu
Qu2/gKLZJocJpdtLJ3hcxMLtCf4b6YMytnMsN4HsiGj9FHQmc0JKNFlkFyfUVNTzB/Hg7CmD37In
RqhXvz9ccDZyUGEZ0Y9cnSzD+u79JTh09z6FdS7xl5rQY1hXQAAA+s+XJVhKzAynA8ZC3O5QzLUE
Z0nNdFqZtThLmbKvgMfxO7FrXpS4HjsvohKh/jWYez+RCQOb+ZDhnrjjDPOCcZ7S+F02qCDVRgzP
84OtD/+3HT8jq+Sdl6HuHC+xThxfOkBBvKLs5VgvAWXStG/ePW39jwzuqFcxOjuJowmwjXZNiPCp
WY7xQht/VFKuWlN0W8xtjQ4t0aDXdKGQhy2wypnr6mKcN+TZEUDcIfU6/SxWLy3jNuOp81IVxnjS
YyEzYzm+a9+jworYHBFrmvb0PQMtRGlByWpb2nyjb4/z/vtV0pMcPTDqQuHVbkPxvAEbr2jybdG9
ViKh1HiEkbJZb87LNyb+Wil//Hph3r0aJip8ULjxvC6LeQpxjqi0D6kgjfFvegoOBte91ZKF6GBw
I2uikUj/b35lyGQUA9KtE3mtbSFQ9Uy1BMkcqEzhOpDz6zo57SUNDtky+tu5/Tdusb+ICX1U3gP0
5gu4pB4dRBlB2+XeRR2UyCYb0vAr7vX2yftLKIva3QGHyHih4bb1wmADcd/YJPir3A6pgOjOJJXU
OApDrLmwggD3krC3wMevOhLetMhvaF8bkAMyp0BHlwG9Ih5eXBBPB9BIzTCMQqP6FxisQcmcZpyF
h0CressyglWaTIi8pX+JUROjpQfq+0ImkxqC7VNTcK38PrpPyphzpI46R2EJUhMWSfSBxj+G12Qt
ZMDC/iFZazNaq2e6mpz6bZk8xLzHrhcktVIQvuUC/nBIkhHHLJLtDldnTZuale+Xv3/6j1ka+hAw
jEYrzhBWXQiM9/Mfs4AdiASCT4NGjHNlgp1Hzlg8qvW6OaR4zHCq6OQnEhifgi6e2zmokY/PeKqD
8IwkP+L6iqeYzBorMIVBgYY42j6Icd2iQ0bCHzMTyFtBlurXEHWxCWz3mhB9NoYPctst+/nPEQ2d
nb1q9WB+TJmHojanh+Py41i5627nA648oOXYAzxokBiGueHjTjMxdYY9TFLftQo2MCqxPeUrZarL
gafkfbwSFHNRIWdK1srGW0RhTH9E2/bNu26e3PpcDhc0vr2I17sv9+SZZ4f62smQWctO/p1zAMf6
CVVbjhPTh87NnpWHyrM8m6eJOm6p+eHXTzE1BBVMU99jcUHd/Fib7bB86RdXD/73S4dWGiibyGL/
1emVVvKwMm5stpo/GGuP4SG3q4ZFGeT26IIU6fRbQQxeHzGptEiEDM2B9EV+Pt/9S386JTF0WFi1
ONi9S/rT2HgT9Hl/CFREFnzObkGgfEKT93NN5TDva4mcNGb/9mXl2AisRj/g8rZ3otchWaaq9wgQ
QzjJcaGo9Hv0J72FS3WAgwttVC4yXu9IGSmMovfq1l74pm5JHlHUHEZ9xJEQ69Ke2Wu7JyHnPb10
nQABo2X50S0HVx7Ox5wCAOT6ROfpl5jAUakFVbs+uuNNw34/WEu1gR986BrExwhkxI6KplDnnN11
4K0CX0gPPV0fAA0AFWiCnzfJfKtC5rczD25W+gPTTIK7vUtuMoDC5BLx/PhTWYAr2DpyzdNho/Ge
Qp16v8pfbvfNBH65WViPeVKnsrdEVJwEyFy2OcgFxm47cQyRL/mrHDWYv5KJPaRqdq610p8YZUVb
pyELJranqhzMPHE37FI8w7neic5xCemyqYFSIIHTZS4YOoaou+RTVa71ZYjmp9MAnecn5SVYBZwT
Lr1w7h2kS9hzIiqx+wQmhXjIgL/lX6CXunNJxhVM8uvu/N/vJGjiAC2Gdp2rXjm1fAPUiSJfBO1Z
RMKQqDe7SX2oLvmZkVKYT9mAKk/Z8ZRGwMuFcvaDfJFqUtDVCgPIWA86aqur06fRA0n9FuSqHdbG
6T/+S9SmKtxVDsAFkZwWqeCVHgI8OXZ6eH5qyzhnISuBDh74M1SEZ3JqPsWUxjVo4wwzv8eFljRa
/yqmcSOsOqdqGo+ItKFWplmdg2OE7+yLGfyegjuzZFC/86FMbEFviIlLrRC4TWo+x3JKPqR5J1RZ
bt4oxTeOo5Fnnad6EQhvpPzBlRfmKtcyE4pq2zv2BNmmBR2zTbWl4AY3QWjF2OSDyODjKcwGT12G
/DSscKPEDZXPc+QTx38ISJqNCQU2X8DgzgugroI0zSd8dA61o3ujQuKVx05gflDHizdA1TByzfQu
ItUM/6F1y/yJVutEawb93+WULikGQS/+VFaO2kwwqDRwuqs3B4MIvs3fmmeGttiC+9hw1n3iwvgA
ArJTurf4JTIJB12sSCRzZwqz5QJmsRrmCDXpK2vH9Yya3+OCzQa4aswi5CuhT3ILHSAU7pMclrnm
OTsm7qI5L9WycPHbz1sCiW2NPN0lbIbta8Nt74Qj+Wb1OVKoqVUi9d3KoBB7/Ci+TF5EXaGGCVe/
opCTHGAC8wLnpemd+LVsETwy/PvvWQfp3xKSYsZDIKhywsX2ADPlRcFK58PJlIc0iwjquDi+HpFm
yRRelWHO2bA1p6UaiqC/jdxasaJz6DbypONeQ7/gYy13nZLJ1UK3zP1B2qg3SelKjFCwTbUBmzHe
lAcJYFnTnFyNDCSCCWiJvlN7Dwe2S0JFJl6e6FipgGvOCDy8cgJaE4HDB5+38aVZbjbJC/VNiYKA
1q9c/bT1RFkXEe2wjKOrhWWGwSYFyig3j/JstCVUoyFJekLYwD6MxVIwIR0oV5Cj+Z4Veq6/zWzq
RUkBHVZ7CcnhHPHoVVsCpknP08Pm1hcFedrU7csMvi2TBdhdww1XoG4uo4FgTfDTMZhW7RjpgEbk
gag73mIosvkE2CXBc2okqCVJvqJXsTAR6G2OGl8SAVvi4xHScaTl+kCt3Bm7OA2utPRxf0K6svod
XRUIUEpDnzOq7gUzUJ6XHWd1XPSlXhURRKuXOeXh7iby1Ke77yFGKX2m42VTBVtKsohW4YsvUDDR
W6IsFYxrCuJzV+HR05Leyyw8+qiYuBabXtRnzJVKiV9TK0ySyuyJv6LZJ7PBaq9g27Igp2aVnjTO
UZzmLp+YE33kyaMvzz3srJyICarLQOiJi826e90hPJLH2rAMRGsvAlpSaK9Ls2xGyykXDsw32L0v
pgekDF12L4rSa+ND2dKAyhp6JrWX+ovbwEL5tRCrTEo7Z24Np7tYy7xviIGUCFyVnFn5R4XJ8xwM
J0AGQ7gp973VytWArtipPEWlmLGRyy+t+Fnii5aUD2uwzxykKL9xayW4jaS8MKuCr5LcGU0z79sn
iqyzScNMs3MCjmYVj4lrBDb/URWPIz3ox7hQaGy9YeHR+CPGyF0Im7KFD4lTimcAURBP8yrP9DCh
ZsRD802/NNR2N1YVtK8rjjoEpQ00KU9LXx1u1fZVA65xGrHW/FvcieSjwCThUrCSNFJfJvLaq+kU
nFTO68EwH0svzNGXKITWyYnLJt+wLB8PfC3Z049hY5SZJtWrChG/tS1bBHjzLqC3XxqWbxuDugb8
Cs68unnsv85Y6xbSvlCK8AHxXhlMvhttnmQEC1zkL07qmAkVd1ZQpPvg2YPsDA8fqBz49isRW6qR
ptaMfoYBrJXbKllof//wODVjS3UDzJAHxgsKffjRbFbl8N9tBH5WHkTlWVz1zvH64VnALyEfCH2B
4/KhjInLG7/iQjVXto4vdgrknYZiOaEnmG/47PG002vobINFDA7XSYV/4/29eIKc/Su87bCL027B
TL7UGrGTsfld4IVHVAHDcHfRUymmCTcgszPO2+GN6ISvQJehl/PG6jkMGgufqOB7SKcvg+yyVLgm
+fZSwOsNjuy7l1mFuGV7V5Xi4RBgzsrAPcWY+Yt1J5Rd8yBBrA2ya4QQlY63iY31jThVaTUnLA9M
nP95Eo5xD2aENBp5AiYv6spoN84lrtThzKI9ELRAerwrFSGsZYH4L14X12eEw9Q6IXXJoa0iQUkp
GAwM2eSOOtI1H3meDFUnR3qc0J6UIGFnR0i8yJldE2zS3AxbGXxCTuVfENB6pZisQakJdTwfi066
TUieLBX25D79mmqCAutP/I6Ytakey9Mj6oRYkW+WPW9Glt1giwYixARmTYuH8Oel28YsnS33SeMH
zrgDIM+uIjvh2/okD7MmVuZ6MITypj1MkkVm3nXoKl6QRprMWK8GSN3yPAdtfu0CXm/8YZPwELwo
Jo0s6YnIBP4zGBKx1m6QRwTT2zYhp+KyBO3ORMrZcvLg7S/XcesEwG7YCdET3iL0+VLTkxhd94WG
MjSHPcmIyY1HgrGc1ZtZKNPrFrjRAti7xMkBADe6RChoZGqjHY5duT/pZfLOUsAn8UsFqI+nG4A/
YRNsKsu/7C9nVjO3LSkAcyUfwU5yktvdFaf8GV0OTL/1N502VzwgkBy2cNVmaCdoJVPwfS/L0ums
9dVFUgq3LgxoZbXV7myWV3lpg6Aihj0CrM4jgrlcgAfifaLMpIJTP6VkL4aHjjyhj+TqFg5tIWGp
/s268lfV1DXT3pkLCfeQ5NXgumptEhVgZRz6mp7LGXSQwBvtC+0Oh96bF+s3VPkFgFPMuD+5kscr
PMEklAs7Z6YJQpNx7BKomutMiz3MQpCEbWsmK5B6B1xmbogQoFT3Az2Tj2RyknyW/8c4CirMMntH
kup5rB5aqpwYxaMn/4x3SF7bbURnX/9DVegFQCThETIMF7cJanC0BF3rH5fNC97geo+5+CDIAKZz
G2oMjo13ST+ypqPOD+ajizvNhtYeQfxYyUAXLMEJBpljA9CMg/cgC9jAe2tfDWOB/BvHWj3itaB/
fv0LZFAruK9I/smVhJrzfh7MhsOMb6Mk/bxfpYHZY44Il3BqlMu1cToj0A3/ovT0arQ2eSxeTwrO
OpcHS8cY0ldUCaWj5quZdOiaYrmD+LoPsGZLt0W73npGwHNZYx1TdChgw4kmiYFMgap3hrDY4skp
pVA0AzUA/m4bAmViEobj6ZS0McK9tjwNu+4eOopTCM2ohO+TKokKjx0eBoIf71Nna+Fr26lWZSCi
2Smg/fa7yV1FGHXm4kZyn1CwSUYZX5kRNxrVsyygh/xCF/qv1qIZz3W88MwF8ldDlzT0dzcT0F4e
Lb8I6hnxSrl25qRCZo/Lqcs0Kflk8FjxxyxLYw3B7nU8ZSiWcpzg83se9DYgPwHfRu3dTid33xhX
240ZmdWf9YL1ZlMOJ0krCz9cIB/OohWVEbbTCBlH9MSkavFkpsc/ldX2+NDDXt0lB/9uFTeYgtZu
VEmTv/v/2Q/BLOiiKVvt9vZVTzA5MLM8CgjBjGTzN80KeF8r4JNC+73cV+PVaFrvtTR/i0mxsIeU
RxKQxxUZiz3dmWG498hlJypsEB0VBrqcW2G+N6hVrHe4b2YyPEOismBnB1plktPq56xcb5PTE9Zt
GcVQSldjxekJPb1gnL+Iddb02DaafxGoZjCtWY0ihAM2+zfLNewxw4u7qD168efcG0420OkwNLco
nSJS6lvvke564rTrxTZU6Ac48MdgxlkXV+1SS4CHrI9GXx6cRU9CH2W+D2UoJ2KprGAKAnzb0hCr
CNvpZcjVtXganbHEKbFAdMGXyBdD+1LCm8vTfb6EbjXUUcD6cyI4M+A9+TYZk33KpZm/0UXufGZ4
bz78SUpmH7a0a1JDY19i+PMIqzFl0oujwnQ79JR3z3KAwjLdxq+OcbjBvPFYgeDNoHkzCD4Jhx/V
w9hv1JRbOsD17BTZr9wxCt+dkIt9iuTxPONrODTn8/T/u0C35MJPW+HzxjONTp3pRmFL4B5SA+dw
ht09KZs91SMTCMH7iAxhKUpJRsVRdsb2Pg9UUzKqJyxS3ymca8MnF+kNU5dzpM81Bh8ziXhs6bs5
bPx4wbMbdrZELNBVd2Y6Z08oz2EfSo2bVM7bWWPh4x3dIRbrb25STERjqRR0pZ7K83EgZjafWYjP
WzqDMM7aW7xyDLVfzdIxTft11ym4BXwhY12Zhae20Usg5h4EIoHOVATc7x9rnFl56Aeb+wmwuyUp
wjLgyV8rBvoE7yeFVgFnJMWEU3AOrIviHPBcwRMcimidWSRt5E9dl7FjxnRt0oKMg3QJqtT9mycX
bIeW4gsXJOpH8VMygfWM/VnLrbvX8SoAmZcdKX/JR19Cv4w1l2atXXifnaRAL8bWW8ETnfDteEmi
/YKn7Qq0t/HNFE1gL/raxEab+BDP6zqoy7QZrrKyv26lDqnwcpXLi45ct4tm5aCxb2RAoRWsyoAC
n9WDkMx/5b0rGWOQwTBozxjuXv2Tt8Coyq7eFKLEug2nAR44MzW+3bwbJwb5TNTv3oP5BOv7rm43
aNCKJjH9cxOYY1+WCC5bnge8leYwcm2HV4IKXQsfXDfM4GgtrFCjhpRo3H1xb8ZFqS0BUvbKs1DY
6/99yhAVUTVX3mgWSdUPzh2bVOjtLByrpIKEv+Mn/7arQQxGhX7XUXlFWHdD6ExNKXnpYpSbU6I/
+SRd2FA2UWj/ua//oR0wTNppj1dni8132Qchwxknwc6JgeKgMNViuzrd3dT6RIdJi745RITj2FFw
rL8UobKd804b/vgMcGxUq2IfMT+kG1x+2BwIYvt0/Cy24AIEqtC2n18dcvCsap26wPgbyYInOWtK
6UZe41Bgd8euRK2omoe+FpQSaYkRcxhmgDIkR7TSUxbtMFtsAo1jar1etI0NHZQrOtaC0hRnAahH
QbmtO4AjTYkGJpLFNLQcGra5Xm8YqlbX1vBtLjISJVuEWusmIbqkJEOhiJuzxGEs0vyhPTHUvd75
CIa0SxKSiDDHpdmx1mDNMZF75hOsURYUgemg7tRkiSVmrt8EozcjfJv6HwkTz9bQsyMuLkfBh1Ol
SmRWvfxu6t3/IvVULT8JI56sialcLT23cKoPDReOzel5jLt/OxMP30hAUHyHc0o1MSqoFnBiPQ9T
pykTxtHpRtftGnPFRAxOXpEP/2K1UtyxkCChDwFDMWXJiKtmp+1r87qyOm5rBTRPzeAFCjg4QO7s
oow//s0zalYphDA4Adyj20CwR5KCkSriUj5pZItZteKIyfyqCGlTxB33g33IMibJHM3y+Sg3b6I/
QMa3v2I5/DY5G6DOQDX9ztNsVWFUZ3H/VkmKeG0YmYs7BUqwZ58vfalF3Mp3Y5MSjGizKdBJ919i
9kJIZxGHZEggMOgpmmKRJXDXiK0lTv8XkJtvgyM3JWO6kuAm077JbqHPmVPYrvXitQU5K0vseqvv
re+wfEGVClva65wLapwuZbOQU35mKZ0j2taAoYcZ24G+RzBLJ9Oa2HTCtyMoQaJJtkaakFDWh1bF
01nnalINYh0oc1O5U206EGUe4jbVgU9nUoQboIYgLDQxU5bdsfAevE9fVeltLPvsTmBm7xdgx4nm
HbLNZVCatQdH0eRDZwk/yRRFc8BoADJqzJq51ckCTIWEk7fUIJVC344SNoXRIjeEZhKlY2WhkIA2
yqBG8GgPnOC21lgIDY0kQndJm3IBysaJXZjzhkzFELj+zQDhJsKfjDkp8yWc06Q7Pg8g6utZbB71
EhYvPx7aHJKfSox0gCxgCOl4gmd/Xk2J7rKyYTCvSLy/BSUfRocB7ekOZuoQGrrh53zNaU4JDjqU
t4pU6EpThFznqWs30He70OVk2yIPnuEnAl0ZTXoaqHMQvBFDERM8SL2NVelEudXVR0Dbsa+slS6l
1S7+5ziweqzcx5Io/Yq1irDjJAzJ0HPJAxIwF2/CQG8Mhx9XtP7dQ138Y91dTOe4BO2BxuflWTsP
KXGcJxU5mH0dWYiQ3kzM1tRA/x4dndVdnzcKJA9rf2Pc+on/VvpSmr8BN8GbtqzP4nmeWxbfIQPx
UqdMZbUB3tEyNBf45XxffOWzSMDP6VSoVUXsoEacE5j25QtlIvgqSKPV8NpE0WTePxS5uD5dJsxM
H30qH1wHr8OoXyR5mttPsR0kOdhHXz/Xmru37A+O80rxtHVXa5Kvcpt7/CTnjeL+5h46EikkK0ve
2QrZBwVcvMM4rsTHthXxbxwLl1xsqjVtrD6Pf0Ru8E3ZKIOGpXFOo62FXgFJaP8Tt6z4KmU2Zlxa
ST0QCbvrH/E+D7R1wyIT/nIR7ZgfteYpBFFeVKmhdfKciajS3Il/8mkZg7+sHyGgeavIwayvGOkX
2zo0v6zuvAZvj4ofILuQf6qcF7p4hMa5J/lJ9wKrYICsDptIYcBvVltzKBNRGsiQXu6dFomDKw0K
I9jKfJOAlKCR5zyMw5Q5MBJkv2iXSHBaP6TUM3FhsFz7l6L4L47LWYq22QN6NmkOuTdSQ9AX54pI
okgLmstTwtm02aXWrintd/Ntg+d6G/p2sgR8U0ETPH/WwraBvFOHcApCVp6D6dTDmz76PqYcu6Cn
5SrAqRfSk98HmeWomQZqHe0Ian9ywtsUQV2SFoL2J9ZKXcgH7OKA6g6BqFbx1BxZn3kOysIB3J3I
O1TRUXWiVYPHlugjwPi40QtHoySLgTfI+wqCzepfOLgfCIyWdSzwWHZ82Cx4UrMyLaX3WJR5cNva
kGms0BZw3oc24ytUSiFJg3itlOjR3LVDfUZ9FIbO2oKWHXEVHhehy71NauZCc9u95rWEeGkiuxdX
jgvGxxdKc1jiNcubuBHWF0BOhaLo658g0tlRH4Ta+owvbCV1FpJt1mZGAhP6SpSA4wRIsdpw44zv
3KbSounJACN1sC85b38N6rDP1g/DSb9MUaSrWgYQilqGQUr9YB7lUOvb2YBB1FEpeuHye+YHWAIQ
tMHj+c80kIK5VDFKrJpfOCGJNIVaQ40NaYg9cP2CuLEKQzqLSKVj1CCmhPpyFnnO8BZbMAq/SrMq
ilr9Pqdebfxg28QvyNxjSUt1JEuQgFOQeYXt9An5Jnn1wiXl0NAc/althMRUJO29ZZxaTwki3o7n
UWFJwMEc2aCPLlMLRgzXKqD/EXodaBzD3KxUAR1xifLdzLDmMlB+c3ntIZ4A2WgEUohpTNt7mrME
j9Holku8Eorgf/pOpnL4ayYdEPfd41wjnUPZK6Q5zCGfgQY2RtwTmmO9iSaGVxLiAP378yL3AkUN
MN99PxCuRjorKsi2cEr+YjFX9RO+Of6VAVSeHAcHujCZO4l3FSxj8vKfMgjetHZkZyQ+onlERfgG
r4oqld67098IS3hZDYBsd2eaE9nBR7LbpNkSlNiSy2XYveI83SWb0MzWwePTCMxxrT86l2X8F6PU
lV3vb8JDAGWUP0yGkzOeqdfdxP+Mtw7CJRz2Mxn/vGw26HLxKYNXalQycyY+RmMr08ZpiHJzSmdT
oPXDIpYFbJ7FNE8msYjCgwasDp+N8/mURYmeOtpLOTw/SdzZU/f7Zuv5OW60zRiPihH1UWgA0lbJ
7MStNOYqF5raXU62HVRA/IE2Hj0kAlJUL87wOV18p0yYhvBIf+ueTXJmkTex9BRizz7KYSjHVIUt
m66iYe4TuCP8ptBLKqFQ4Nmf3YvKU4QyrfTjgKn+uwtCppg3uaVCG2aQ5cSv2y7gca77O7PON6GS
xixo6rpE0R/+qQN293dX/0LrszFksSgaq/3+DX/i//3vqXx+NNfQnd4NK4l0Yqo8tOGZpgW0KyO4
xd6jF+6AMM9mwLM412XdUJ6EkcZ+ExUAU+/uxKdYEhbP8Ijlxp1UX2kDBzinWDn45CqMigr4bX0J
R13Amcrtn5vfEt6fppY2NENXfaxArA5SPQoZIZZxmmnKoC9rkO7xn4Ft5CVsGgxHvFwBx0tWjMnK
BnxsafAreYYpuz2CoqC/uIxAk9KstrgAlFzfV+9wpJHZhCDYRRtZejP7cFXwRsT27DL2KyPHAAYi
NVGWNy3SXAkNKlwzUp5dXq65dvWTugCWx0tcGvf4ZTulm0Ly57jYPDWVIBoweSIURHDilhyaXX7o
uI+pjfNUzvqzcHGhyBN7RXL/J4MhIKEWtyuEHOpMZI7VH0XAwPIcQk93aA4+oziPUVWZAFNalk0Y
W1eyS+Fge1WAiy0h2lqE6nshsA70qJuJ2cS7FLOfI8+d2vMDdBAU3XEMA0vMNubySf2eW1hvYJLf
XzQ4xma/6YWix0f08NQa05YP9y+0IN4Xnod2ZGlTuWzYuSzxYQJWJ43N5Bv6g+6NX+xOlZVRBEfJ
hF9QFQf7pU9c47oapVadlCMlvFUHYtyaFd35wGUeLzB51y3BWL4bmWbtPeo1J/nplphd0FHoU2oW
MYy0KAvdgKErr3BKLKtJTAPLgdv0KI8qs/+Lejv10pQVbIiA0fYf9fHk3AViCRrG4z0VDsIguqZe
/7cGm/HgzmIPeRwzCYlF2Vj0KS4UX4fhhoBbdtCP5/93ZhEB/fAX8/cebdLdkiaXUnlV5gED27uK
eonA7jl6UQrDT0TdUrj6UxpXJwSb1NxTKW/QQf7slnQFHK4MJqufNHxQXJ2Nbid6Vo/XVDGMgyMt
PynsKdNEgzKd25zqFj0vz6rUbqqfmBrK5Y3Pn/efsdH+w0eN5gVePK7jqDOVGyAxp8vVXN3ZvG4o
WHCAGBvNgkg7Tw1HA4pO5gz1ooqK5sBqZLmzfLuU2bvGVuh/J+69nRld0SJxLqnldJBdI7RQ3LVZ
WdDNxOawSAN1Iv/KWobGHBwGCqV6D3sPcMavn3Rnkb9qZL9h6lVnpbGnmkzmuTFKqWzJkJ5QGyu9
P/nqhDrwNsnmIYBKNDoeSlEKJxzO1nBjUYxJXTiyzmH/2tUnkwF+ZlqAkHtBqp6LrwDihJtNDkC0
OEbaglxhP+dXB4fK3Xrd4QOV/ecFyG9mAYOXmhbGH70evj/u5Zk58e5QbNf02LgtcYY25xaBSIaa
avkOwrsxG5/PhJ5uSF3H/f96yR7oBD6Nlo7FyAuBEirQATRdANivVE9V2/se+c5L2PqfD+VbmAfh
34PW/YGffLr60K2fFM0DRhE9Cjd/z71DFU7g5MQOeVVdhHcA5b3KBSf01cNOr579gOabKu5XLvqQ
eLUiV+dDGCmp9JV9zEFoA2eCEpubMTPXUqjweBhiGNZe1aPLuVVKTThHwOToEvgITdqFZg3nRBmj
gaoF+rjQL0VeXDZFw5+Sryal0mUg7F6Y50MINUTqx8U0JrXS41FVH3/OyeMgFSeQazjzOVi4bAl1
lm2hA9wWr3U8H1K5dImLNwA13ICN4QtbI9TRHOVaDQ8zLH4kt/5x7hg1bDqU7Hg8gGoD84LnkQvV
s1RcT9g2XYghYgsIPkmi20zkChWSL8JQp1xmDkaPvqAXLv5e+wc6wuyTIXaTMVZhS3Aus/Vy8tBN
bXMXri75uEXlbslHQBGLUf9nqqCsl6ommgyE7AJc/MXeODfpYcHcnfKYJCKD50nD0bTDGzAfgkGx
1NZ7Wbd2LgasKqDm4kC9e1jcfChPHdjsjJbrIKJPqqs1LzMGIZ8v3+/bFF3lDN+lIlc3L7f49iBU
+JavuScIQjP/YDGAMqjDDkDazwMc4nxuXhagGm8RjLwIiUMAwdM01zx/psVsbqXTzK5LqGJlY/WZ
zrZ8ATjKD53YkwiZ1SQDOKJJx7rcOG9BOsa0Yj4i3w8r1Dk9vQGfwqOnLjadDpZte2cVWNVEhB70
K7bPQ6Ucx25Ea7bdxJQu5+8AOlCI3T74vsrTC+n0heRSwGkXGmXBgdCYAJWd4KVVuqyk3X2a17vJ
7HWodUbDcxDnJL9Rs/7WW1VBRRatj9EUrox1oKCgxE9UNOedHVra/XhRpsFammzT7oac2p+t8tXK
kSJkWZ4cZPM5Xa5e7h4EVJ+m3M9M5mZFfN1PLioo6xQQy5JXqawnStxj53gigBFSjCx91CnKplZX
hxxGriorPXmJtzXSunv+1R21JDheoSH329Q3n0zeG3EeE6JTb6bNV1H0evQyj1R+3M4F6vC3K18W
9lFa8SiVvoL/Xh5ng10TOV9NXm6wKmFBRTmmEQ7g7SmBei7HoqsnYmkdNOSHIVGHJ7PDFOIFs/iU
BtUGpfiBW1qn3CysJyriubT4DX6Of+0bSzNH+uj5FEGmikAkvRxqMLLl2e00P0zW9cDuea6soznw
5Ei6lBi22lW3Hgp1zn5xsdMeSOV/7nVKrB3tAFxb9gmT2bpk8yESBSUOWp3E9oeU3nbIU/ttvX89
7nkQgVUXxvqH4lqDOTmvKiu4B6XuEFyja9yS3qRvZyWiPLKEMJV19IllOIiy5kB0/xNDIZOfJHUy
iDNyU5LRXUWCe5bQnsc3JvZr2aZxCh6mp6tSwyuvfn0vqabK/SUjrqLe8Hs7kxvTZyck7CUhy2y7
Gb1n1g2kbgDIZhf+Nt6+MjYupYpGYgeV92bBmjtIdJh6j/CAN61Fp0TnP/5nnIWN0LXpM4Vn3vKa
OZOD8lNmzZiUcd2yBTWZNuD7tu6/mKs6Yozbn/QOcrAjhOZUsb8FxNnyC9jqy3XUdVqlcd6yaBAv
+ufrygsKmUGEk6Glj55nYLB2DR741Zy2FbF3fKN2EnQ6RVM909QWX8NEMaESG4f66v8Cz+r4okRl
bSWH06Yv1pkuBTQvW4TDU8XI6ToRdWs06tIE3TooSgMSSVhpZKEK6wDZ1GE/YovLFgs/83Pb98Nw
LgxLMkyRNcxvO0XJsvCs01WK3nhS/qckOrDG0hKqXKo/h8/9G7saCh7f7KVNI4Mi5tq6GdwBKK8m
5EYwhC2Df4d4TYfjkNZXZ+r8JZ1NBO/Dzbh0oa56ujCMuOZyLHCwPsg0FOFb+JZvfjeZYMCY1u6L
XLkzAqAGfrwWR8+ZpUArK0KDcjpfODimbY85dPGq6wq/Ykn4oh656I5JxOBdpOwI1669X4N0wPDA
OQkc6vTxMar0TzF5AGq1jo+N+x1RZfBwskKJsxyNoCkTi4TCp7rhxbt16Cq07OLqghwJFvs5cB48
Qlrom/uJfIo8/IjhFqijxgJ5bP7DcxQKNLvazPhBVbDJrmisXp3+PStyveI1Zu1w03DyB1Yajh0v
JIysZJlup/kBxRJbvWfJE25apu9BW0F6OHRWgQKrm2Z79sANFt/UsG30t7IBvKZUWA3XAzpQW3gX
wSdZKLVMqTfWhe+hTRk0FIBnATEL1QeuAdaUlyENOqKs9SSLYpuByVo7Fbi9T4UQROePRumwKpBu
iJqRYCpIScn3ZNgfWiCVbx8Gwg8/ZOtoXUSFqHuTzk4PjwjbX90lcHerCMc06IswSqCqGxRptws3
R2tE/G8HdG+I4GMVXsJ/uDUb/yDkKVYCtTiN7BWoS0KwXH28nlvLIAqZ9WYjHcqSbzBx4CS8aqjW
ZxJcsdA3pZ1+5NEwEbnMHVZARezwHruYAKT9HDFHiDMbPB5J1ArcQdfMYITbkQdKd8lilblf74dF
F2Pg3XWTakwWZiKeMyaU9cozwjy2ZjfT2HsP5wyXwsQLV2IdrDiKroKQ23dinfBD6TAlDQTIVVd6
5dg6j4UeL1I7e8Nw8FM2M/Z8zlv4s54paGA06awl6cP+BGiyfFE/S2DxL3RUPwBLvwDFjGSFq1Hc
6iryA9YFduc3pbmbf0/wgx/HDpX4hWy+1Bm7soqEQG6KfOYrsTYI0/T5Wbj/t6Z1c9Uf08JgmODR
rqulxOlM8z8DDOH5/nuzieejigvQmYcEPTm4xC7axgRjwkrK07n2Q++N0wROpBay4ldUS+jCcQcd
Q50raPRZPXGd31kwBSn3x8GOOTDh1EIND7XJYbxPqaoSbAbvmZTHw8sDtMwkssNsoM1e5Sa5N/lp
r0514QDPSSLl2lZUOm5TE1u5M+61uVDq/WpzCL1NTqf3l10dlLDUYuxvWVxfvu3/eGfdDwGwrcDd
skQO01a5rDTEXQQCzfxh1zJdKgqdiOLN9EWo3ow5i7e9wgdVxeS3SlZicyKSi+G7wPHbqmfGM3ta
fTwwHT4Cvx68oOawkUrOUofsdwejaDE1rupwR84Ex8LIw4QGLABodl+/VZ7Rip4Cu1/F0/t19zR3
cCI7tQP7aNh7novWdlA5yCUoftvY6X4qhg3JC8QRlju65m+rPFKuZ+gx/pYeT6cfmKbZ/JtccZvd
RNp86EuDsVGjoGgD/2CZbt/RotkE8IBDq4nMLv1rFD1Bsz4bacfR4ZOk1j1iu6JNDM159n6HUfc4
6ClwQ8Y7pvndBCsMecRXYrTwS8uxS9IguE8PuX00ecoW3iyssVxWjyxz2wH5v5RWJmPYk2h/eUwg
JymPr9MuIFJ9/q6i2EhiL21iFC+s6WfCpXhU+BLrRLsFRuYWEVTo9WjA0Qyqxq3KwvrKEfKTNla5
ue98nbXaF4XLW2I1ddafeWlee9myveAskt/Ds7DGcIRlZJUdi/21+sJRgIeRiMwfUn5ExFwncg2O
kD6Ku7E1hkHbdpby19LBIkT3+o5SJXt6GgcaMYVK5yf2qD8sc0GnR14kkqgUEYqKAH2Q/Ylaxmqy
dW2wr8siJR6lObGAVB9eofvSSwrXo9Z+6gQRWOxOMCe/Po/vbdtooAKcY1aqqRw2BY2U8Yt7oJPB
JJ/Ws8iPdBRZRo3IJ9D+Zm8EljwueBz5HYTQEfvwElBJ9EQF1EOD0ihMZw9AojgpJSbkZknoTl7I
ZiMvh9k56xC2kmR9unnpD9bh3RPkfSU/xIvWtztxtx5wLQyC5uyfO2BWqcn/Z+orzSVOeqrR0YCg
lsqOjQYSdSLyqCkmPRK8x/QKTVjLPHrJvMv159XOcKGCka2xDauH2OqAJOQcNFcbnpB9RBQ5Jicf
yv5TJrYaKuTEg33p4zjnJGtMje4zucSjek+5/NPqXlokUr+Bdr2/+0qQx8l0WmJNtdXC+e8zODRF
EzimSSOdFIFuRJX9f8XY1UUOq/lAUBovcSeT62JH1bBAMaXQrNXnIygMD84FDepyIYGTsZ/ozRMU
iQ/aN9ymuxCvKU9vQm9rvvIdmXLzNg8N6y6LO/ruuWxePJ7s3xgErC1O6fAf7IEel2dhauzyVTtI
RVrbYC3DGOiAVyPACdglwD+THoEcvw6WnSXdzwH/N6SK/uFSkNkwLs2ESGnC1MhtOkg5Lt3dWdPN
F3qgqD0iLoGaou4KJHTG5pYZorpWRz1iJarg+QvobMlAqy3mVgI3U8aXkKmCek+HDM19aopULTi5
M7zw3JLrlWRNs8CaQYa0LpbBtKXJ9bbWgxhulQbPG7UbvuN8bYEpriD/6HTzuQvRA+nefNXT9M3R
GNz0UPt4pNY6AU3taaBcE5vZFR+0kcPp423C07wIm2E16NJdurUUEVncI7wWt35AnWrWH0mAbxdk
OnTn2ui7aaKfSxCm+9ZI43R9hYJj2veiXIr5UFpuopd2Mtycy900Qn/UWSvrUb6DvYi3LEu2VYSM
G2beS8MN0WjANAnHi4meA3Hq39c3HaUGa3jB/2tZIfGh0CvT4qygppnELBjkrJoJM7fH/vGu2iHW
X+AryEr0pxLeeiGwVnRAxDPjztGKr6XeZw+nP2ZuVSp4WCD7vpoAdcRlvC++h/pCmkykOZ9glyJ7
prmp6q9EP+StzrJQNipIRQ0SavgGsrAM2kFqEQABOl6nIldsyFapQgzhlDuJZsXceg6uxzPJ/FIL
8dYpHjHjKidF/QVr2P25+1gDb/NBY1FbFuQzvnOqG+4owFvxD0crHGMxNymI1xyBkMaHgEP55ElH
wUF5z5lc+PVzC0OX1mZTL1JsXKQiNpqssw9yYNLNpAlU2kafN/h61CVd0JLrbFTxX1VWHV0dT0LB
Fm2lpTYW7eet35Ti7qw030SFBZy9hDie2Y9Ooa93LDiWAhp8gxRsPjPFPWMrpXzgrrdnRje/VMHp
F2zanOojdgVPUhwPwKrItnZTBFd/nTsjHVPbalBoixzlKtQs3xwbeWY8YbN1TnJWzur3+fhzCgnt
lWshzadero2Et67X361xBL0ELfyIQ9grVQZ+pQX+twD0p4j9g4N9vo6iOkyRdNjC6oglgwlZaSiH
cCS59mbMq3gTJCiAwM8Bx5S5KAYoNI787Hs1JYwZkJSUIOhO5xiIKg0z3yp7uyi0ecvKgvuV9m/u
P2bQXNAK6DCtqY2C6cfrApfvp4HogxFg3b0RRK5j6EmilZyIKTYRkBPWMWm06abiRr90adqPNvpx
VT7hX2woFxGwqN4XnLfH1INpcgofAR0BFd44+ZOZ+3H9UtXFmSecjp953eYrz3pkSjCqc0iDllX7
b+euH4Pym57y/wKwqCgSFnC5ImYdlOr7gi1ykpYcMvYY7oCJ1+uwP/wywCdFzvqXSnTJt461HquH
70nYJOVZCGVP/gl+0c4qESG6QIbmdkwsLVBRE/LFCXxEDnjZ7ie84TnHhbA4R+oWvWK7Uyx3l2Ki
1z4pffd11yZZhGGXVNZn4auxVYmhiszq3NnQWtqU/irO+yETI1igl8xD8ys+sPI2I+8afCnwL4pZ
r2irKwAaOELvpWEI9YGfv1hD785gruqRSpJ3zy8OWuYE1EHUlxzrSU9kIVTP0JHQEPND0u93RQFo
Czux5NBQyXIUXl90esbBlvRQeE7XG2wOX7JAOYXeP2uF/aGW4PRsv9jitxnGUfQdqCN77lxWWn2d
9JufLe5T0wTHpCyNA/bmtuDkfoWDCCvPuMa3FqWIoZg4NhUScmwKf5PHZCRB+sz8oab3d9zMQtiS
tS/+AoxVjYfC9KSQWvDUs8yJQKW9yacyBQ9/ITn67FaBP97jLKRO3ZJHwUK0I0ZUvQP/FH5MpN6E
mqxumarCd/2JFOKMdHK1tpRAcGIytIrK6VJGDHBfWYd+yqAt/4Hd4daN8MlTNRSlX78LfcpqyN5a
69hddHfoWfRHFFoMmXm5BOErkmaHz0wJGzIippWfhvRf0wawdn6PVBG2ZdaH9aZW+GFLHQywA/jx
SNUqbk9GKnJdWGeiXnXMfxnDanOw68UuO+22J+xROo85auXddj2z82IJjA6WisnnpFAuEBuAil1Y
dgw0hOyRQl34+QK+3DRKw9XvrEs/iYOfuXq0OGXRrqiErI8tc4NHzoaLJnof7AsMvb4A6m/sq04X
vqr5gppnMZLFuDeLy7BNrCxQfurEIF4C54yJySd+kZiHcqRKVcRGqNQ4xMI92I5hOBdAs3MwYIH0
Mag/jUZBVwt5MGNieIjvPMTgFuWEJEp7PdeWZI19dZwnNeKTYonXeLP6/cdoXloi7zzl8khI/XZq
r3tAGFZmhV3x/FmiYP4ZH/XBa5jOmbBVE2vJXMtngWUP+ofe8fwPpNgJg0FyKgzDtFL7q1BisOq2
GrpBFHT+Cu5ffbunCxuKouSYrz8KHkAZeKUwX2E+467FqekD3esLRYLPrOirGjFdOoPhK9b02f66
fgustnivUU4+EPsBGAVkHd95iicwVbZK5sp8Bvc8cha7IjrhtRp6ZwcMFkdme4gkF20wwlShdB3M
8yU+llr91rzhQ8Pa+A+vIF2YHJ3nAAKnOzWWlXf7EOfuRkSF5I/PxQc3XOuBY+PDdfVyzqH8Q5By
qrPuYCgVsmG7w14hxuzcO0IE8Ak35jDwgo7tvO8Ta0C+ZXgcFVvTR0SClE36hWOTJc5M8Jbm40H6
xoT/E9Ydaq2zUY/NCn37ssC+Dz1+DK6injZs3PdRSKVHKRxbrOJmOPDAnm4ick6yu+oZd8qP6eQX
IL9/ZpTJHfSstpGjcO/pCqJNr19ycYQOYjGCWm9bvpP8TpW7Xlk5RtiRs1kbTzh3HYgp9G/dZCnr
EQLuroV1mRZrVSF9vX26SPHeQFr6l6eleaSQvlUyEFbZxCEgN01GpG8flg1c+06xA6VYboo8mNts
fSRRhxszJda0HQ39iKSoK47qk+oz1wrwt2qH+/ymYeyEz8N//VUK3VB+k9z54M2cdKRF3eIsqGfC
T7v5ZgyKhxTJrxaPFukMoTW5gU6DMKLugbL0T+uKsoUfzoBvAYHrIf71SS1tGTXMuCyt/wfPftBU
Jn5NN7sPv2HMcC2S3fGfDin+Bynt0E0erNkg+NoRt4Das/emSYx+tZvThbTExZS6hqAOJZIDZzDa
ShJBeduA2yp8ARjT1JGzRruWYWxGsQeknjkHQ8tJr4Z9kv746LOKgt1Ms9j7NKIVlx6Q+VqsgM6r
+o+KE1Gjx6dGmOTC70FYn7TpBY58QTVyoHDIrC0zjX5YTudF+k4YhO8uhL7chv6dXamWGHMGwdCi
Wi8E61jOUdPFxZLAn/3Wke7P28gHS2xnvu/FRzGgrQdqsjDJaymbDlii0m6Gf0041t0IDVI4TUHT
W4dcyYXMrr7BN4wjpTdHaN1FXNgyz+Gg043qoCtPU5LQiKePHMHOeLwV061crdVtUiO0J+t4ga+Y
ZpBErHBbprIJiGUfk+OTyfT3JapFSuqkpbByspXlzE5wmXBFNnfry6zZuWjuW/0KEkyFOPPlQsKL
wI/ekrcxcH5FIxOTo+YW2jQBqrGYQXg6fd0PfWH88QSDitNzHBBKHHyibX1zw7zL1ztzhD81mIBS
q0nN8tRnO37U4142H22rInIltc6La0JiK+DZEIties6Tva9Tn98a3ANihHKxy8Ns4gTIyH2VLGbt
kCdUTW7WENT1FmIiHrghIl451R5udiJjn/WsNsEWZo0hKfcdD454hMYChRx6JZhO8HL49M/r/+Ns
mmtHCkTCuKcB+BPtpke5+VWoSTZ5IoK+N2bL7frWoilyurzmbMWqfeL5Kx6qOGemXIVCCF2hbVlk
d44ypXx/N1+isa5FzIf3MP3IayVTS2py45MXmagzLC3YQHQBXsUEhX1TYxyhjwuBaIwPgFW8wlMe
3z8w1kex2JfB9uNwza6M+jKi9bOpoRTwkUSHeBeInxk3a21HSGTVUqZpV9Z0DKEPowMRpi4iOUpA
hjf8gQb4Dti0JtqVwtQ5h4FkASblLX7qswfGTKlcxQ1czAh3La1QYVE2ucg5NJ7rACA4BWwFc3uC
/E0ybMHkMN1iliD+2uVCIN0hLBWQzJw1JQOcQtSUc4lR8oIUbRXtkVu8ZmfPC7ZsugN0GKxAeDYb
4cp/zopf7D6zfKj8pDCC7/8mbtF8hqS3Rkv4VmoKm3nnEVHbt/fM97iYw0UQXdghpYC9AFrXd7xg
8OcRpGlf7ejUklLqCdMSN1SxfdknVtQUN98cloHq/XJ4fspqmcGTc13fSvi79uZsc2qxI1PdrX8U
dlAUvgdOowpx6sKZVkTNIPMREtutAoe6HragPDxlnnFNPdtA18NuwGIlwstklYiceszLzIik2rTq
HtHnUf8KhH3eFJHxmLfi76Tzl8tBLJFLcPR4q8h8nKvPZmj2M4m/Uk4zK7ewWdUo7JV4jU76mDrb
8BB6qfnAJ02yYA1kzm5c1S+pPROlZP8RbJlao82PyzIQUkAmnyRN+KKIwECmSlqAxc/R9GnwhByl
qNPNuDEH0JBg9eFEY2TGXg5AbhgQPl2tx/IUj67qiLVybz5GQEEZttJyX/WYjZiIQTnigsBadJJb
e7/OugHbnpFoyZLm9xXaQsYT9Q4zeUOE45ZtPdSayOq3ckIDO9Nnl9AImEtm6nwhQwVPf/KORFsy
TSBs34yqqkxHbSxjToxbAxpuT0WsyHHdpKe7kM9QDDYFRP8mKfzhkrgpFNLppMvel2sHaf77CZ9c
3NfDg8swWO7d+lcyWrTjDs2cn4ZR0S7NN3GGyT0jH6JSQdAcoUNnT2UWJB3tyVV8daxkAtghKn12
xTeZBuFaM7Eg358anVCvFM+nzjd3LTt+nTLB0p4LwnAeN3oQp1eIrhOfAmNXPliT3N7iLkAOjO0C
umeomqc/i4LSMNmsZdtyxXJTTu9agD2kI5aX57/tNiPMCMY0ozZJj7D6fgAaYCs2mWuQJV6mL4M5
1me6+mr6KGdGot3XTfq6kZ/sLOvlczF1Nyl/aT9rvYr+GGjcPn9mZoSM6ftU7qVPjQwNqsrkMoj5
gdhqF7ggrnHoxGmRT+n852xEOq/b0Y4CzmzkHLs3GuofOnhr+DhosYuDrinlPD1QE2v0V+inlnB9
bKO0p2NJmElZGEtgq9eJ/4jDhWzXjdz/OOYh1ni7jwpJKcw9BLDd1R01n8MvwIxeQihGameG50lc
t1hhMMhEBvV+SxYJ0Vi/98PviIxSvFt/xyW7POXQV0eUqI7heX6PEyccaOxgec8ySVNPjNZMCK36
12wViBHdbzafq+118aFuMUU8yQyYt3CTHe15STR+XxNokL8hGe288YDbGzA2g36Cv+G47olL//zj
E/XReyY3XWKNScNCOcU7ZW2ta/Wf64iC7Nlc4L813OLHui88YCf7Yz1DsiMx3N75igOmU4yDmfdM
6+1vm/vJcChPPBe1jeLSlF8BDFntDkO+4/MW4eyH19TJsCQA90m+R48TUy8qJOgHz2TWnbULBGFK
gqdOjGiTQW+z/Vdi5sfZB5EP8N8c3/UL4c74a1WhdqizOUyxPLBwo0Gih8EHzPuIrTONl9ptvi24
D7l+O4ray6TDH3V3stC3kNkwc1Rae9AFyoDoo+Fwr66OH5dmdLjAcS9bsV6KTLyM8Vsql5i1duxM
JrGBXmMcINQpGNYduMsrF9y2vuQKjeRA759sX4Z8DnFUOa0eztY3jzLKLTm79KUEO7o4oNw61aC5
Y1pyo+mDMMwusHUIFNYb3NXNM3tPgIIGNwj2a6XaajQC/RC4AgsZN5dTFl6SJhjmfybXpiG634Zp
+o/N2l2WhcWQrqIy4zMExn69Chv8uZh1eF4SNdG8QAcco0zzyK08OeO+gezVlCbVs0F6ruZshVrC
rFO45/uSAUMx7QGUCd0GPlTkDK/jdJbs+cItLWlNqG4Vp7Jw/awnD+XxVmQVzk2fCCXalSHzR8kj
7g9n6FASxKnAF0VOJP9+xnnlntIg7o3LqyNnziV7YJncRZIrL1YgVH/voMl1lUnJDVDa7W1H1U23
2HjhX4dqwFmqlpsoHiUZpWSR2owxYRE0gxUW8Q1yE9ma+mMDAk1f33+9/zN0GcUKkpeqfQZ0Vfyr
7jBrcNSLHE9oXrGNWqpEjpVq5XTgfl0MlHlTbLlq2sm5h4B5LG1j8gQniImBZFX5CQ7k2RcwsmUP
Sh59tB2/fwdZZkAckzgCsfdsEtY+LrRBBMU4mDqfDYye4JVVclIammAdJerULHSAFcG/oW4Dllaf
IHBu3wOGKq0yVWigBUa9WrwZhOrW1dN5/RQO3eOtrVig1MHbaW5Z3RArohs+7Fym7+tU37IlMyOx
MHcLNcf4OJqxBr3B2wrCz2TyxtshiRxCujsF6L89Tz3CBgacOKHDs7IsQrbkp1hcW3NPdY5+Q/xk
TcMZ7JCqdxN7CZtPuRSsm0ANLqkWd8dyVASEQiVFfnc1KUTNM8x/ygQc/Yq4GJQ1WiDSRInS5mM4
iE16eKW+Tn/6X5ttFMr03Zg5BzxGwNO+Hu9XFDQ2nZFM6pEP5Re+1YOcTWTsgDLNwd/GlSiOYEPJ
Cimt541KYrs2nTkY3qLhX8+7UTPfU1ni2D09d7RsdciQQIW3x6lW2OT0Bauc+8EWdUFboTTGjjD2
dDdl0vIcx+O5cCbhd/Cj1ZI/srddDjNhGwRGMVoV/N5+NSDYr50wQt+MBI5a3bI+WFPmp//jBygE
eLwzb67DRgDBaSumG22YiVg9zbN+hto+JxaMYc8PB5dX0CMNWfqW2PjoAXiVinn1aa4XIuB/TIah
UepUhvNzt2eDsNpRMmEeqwGcZ3L1AUUrWXs4zSpNc9UaMk7Y28bhLLzYrakZrt0uiWI8bwxqh5Co
6idvhb1XtR00VPFAOVn9p/qgcS6u2UtWdwm7nNnUfTmHVRL645p0hAq7dQShDW0f4QLIlio15A6L
pXoCepIEc/Q56aiBCdhdjl7iTyGESOin+np+oLsCIxFyi5iLjvD4zbte5Qvzz8d0fL6TKoMMI2At
TRCECjvae2ROAzocvNRKjRRGBS7rzymBQzA+C5FXaJuWVmaQXHiHqRE2CR2aceDcNCXrMNk0wO4/
vIcrxEQMDdKO9XM4meUuiqeJ5lRLAJb6JOoBSRKcx4jm/rZVqPdSIvG5thrq3gkwp7KA9xtEzTFg
Y9HowKAyjRgL1gg+aT/WIJsvWPlURPMlSlZU6rKKnavuYVYMq/1q1QFmSgWLeWRbiE3r0MAqJVJ3
emOAUPeqIGPST/3HVqaJPRRqrOdROgdNMvwy0Mgv1Pmh7Ldwgz+LE4hcdxP2GX4uh9iyirC90DEe
sjejeaq2oxNJaYdhxJY8E/uYCW5E4znTxLHwuNetlQO1jubFDZC7BAd+MVSJdquuhA3VUxdeTLA2
X0l5bQx9UV2QHPpvh417fCJXj3GdIKkR+fu7NgkPBsyJS9BE0UogDl5z9tvEvhUdc8muQDg+G8XE
3zjwIiHub1dKdYQ8vX12653utFsOCZpeFcNK0MgDyLC1SS2/SJP/7ZDnqceWtw1/eyLg0Xr8NBRD
VBpaHMCTb7dR/Sh4pjbiQXhp39lXxFdC6Cdp2jm0o94bn5iBK38iPvxxAeq1btKRG5eF6XEYaVTX
TzwIAj376dqBbS1zLCspwssN5TTb6TtZsSsL/3i8sgDIEyKHpta57OgbWTunkjhu33+QrDPtYcYt
upp+wYVbP4v5mWGzAbzuaRGzKjjdI7DWdX38XEYq7AWzSx3CMiKjofBGCx+fFgO6UVVbTRiKElRj
NZ36YmmHF8E4Ra5dzEsurj8BYq9NGFTthucBFwZmEDKX7TR2ycC9n7Tie7vwhb2/l4xQCfaANhx9
0Xd/9KyYKujEVuKn4XGm6byhOvjJKC6OD3pCrd9UJSYMrRGMZz7S0WdTrGkFSdsxpMO90xXMhs0A
8xBADRN1LbrLmndRPXRPbKNQhHX0rOeZGhclgNp9fbNE+bF+NNVePaa1q+8rNN7T8kumqMHooTSN
l6/VdFR40AslNtGOws2YSAFHekIKxfond6wHI3L2g6SARiyDrECKr+c8smMg2xCmc5XOQikZp6Gf
FYxbFTy2NbR/gVfFwDKcy97wFbfPlK/TvkIOWa5Hvwp4a8LZmHhpWp7s2WUEXn4cmmBx1tQsB8vh
HRsMDVVMTqdhaTzxGMXZB8C3yJqQeJKTb/m2tZMwXpZR6RwTkt1d9eUmXZS1vv31Erq5szrwu8Ud
29J+pPCWEHT6h9diNHT5jUCOhMu9/Aq/2PCkj4bCoIH+KJrkIV2GfjNx9GJOuRU9qLAuLjc8iM6c
U/xkYfKq13V9sq5+CLEVHFru/UvLo/NGbF1AA1BRlBM2JEf+cxsQw8N7kujHf+JMnY6gTTRWHV65
SawmUqeil/cgrn1LjoM4B+F2WMFtEgx0mFc7UEsSUTS+iHhZklcp2zPRHYWpKJamatt7u4fRKTIB
DBifBY4yO9OdkU7U7fkuZwTLiNF726FMwhc3sXU02xy9RdKYWNj0heK3UmzmvqgCDqm3g3EDGOwY
lJnGjtplq8IcDecAkCgC9c8Yzd330JAWDkTLMZHuzLHxDJD5FXrPRouQ/6QGnX9gebkuYD9WP2un
A7jkMqUGUPvHRN7hkD3JqD56pocIeD2EYfXTiHmLsl5bR07HAlJP/a+upBz5uMI4MZ5VtoqR7iiT
TbIS09FOS3nMHhqYOAMHhB2nNeYbNvL4jV+bDofxUQ86lxaeccw1qMrdaYY1MeLSAbql+QsrKYPD
v8+9579bhKCgr6Uny6Wu6CMajZeuVi6ftv6fDdvOGED44jB0JMKgmvdDPUgmdvPdwi8OzSfjUef/
J9PBo//+E4RyxhJ7guO4nHK65KSnyp7ahUgDfdcxhuZHqKxzdHo8ZNzVv2hbvLyArtkY9OGg+MHR
IllrYLhmXz06TLGIT1JU4fnvTluHvWU9tK6++sCTmoRk25ZCQI3gIvBIGVLYrwfqYeUcNtAXXPsh
wJfqFsUKHpqZMrFO/7MVks6YLI3/ylHbZ6xR+sPOrfmbUtHfiEfGvcdCwRXkhuNUfRdtZpN7B9Wz
KvdhTKoD21OLeGnRSzMtljr4R8W6igRsbO1jI5TEayIdMKyAFptBNX0zVuF/JMgu3uztp2pkNfrc
gCDewqhndrbu9BFed6iLPPXptjNy1kM8UEWMSfP/BLLkJmypcY6gKGV5m1NzCjdEpqcRoMRIbe69
PSshzHyJ5+TOahP4A+NuhufVrL2PKc6QS6tp+/7B2Gls2RiaRBHM7Tsxk2aiHqbdXEmDWjaoG3KM
lPWMjJXwssvFIW0BAm7DAnU9phzHnyWxB9rTco4qjkSJ4hu2IMN3F6v9zsX3F4jxQgHX6RAqjzI8
C13X3JLlho6VmKiPXz11RzJChjFAXV7OIhk4pZMDmfOWEYPo+g1z+c2cZNiZLEnB5sFsI64Ay34A
NoANifCFRbQedHIyQ3ZL1EyMnngQzT4mNXjPEazC/G7noNXvKPR3Pwt8KaRetV9+OdPpvXFdDu1w
85Tvm7SLhQuESaL6F38sWVbFCSUKN6K2drvMULK1AMtXSYVACEA27qgm7eb+lw6tZ5jdejEE9BF4
sp4yRaq1e0hMg+FIFVXJTVcboqmdpBaoEIZvksauHgoFSr8DpSePikPQHGZUC94RbySR8NqcRoYz
f+GNgyfSJ/ulswX8Rclumfu/FBls3YE7eupTNlrvUwas3am4cURY8p6Pium6PnWIfH9G9ZhXT1v8
zYmxKheDF4KoaXnOKHU2VfUA+gYXtCZM17R2a98cO67bnS6MWo+T1jTlIYxXbIfJpQYNDOUxDk3s
75w/X2+1q8g9PKvBedQ0+GZ/GHt3i9iFX0TExymfCkM4X8F1GR5uS9KEJffe08j6FOWGXwGTGBg0
JA7hC7+pOb3KIpr4OI30x+VUHyTS6P9DnFnecGd5ni6JDyLmlWaevE9uAtlPljKFASHQ8s98mGIe
5+QKkmiV8UpXNaPFru6qPZ4rGVyNOWKMc2RnJQP2omDdbQ4FOeSbF+7xj6XA4HTb+mYP3BwFnktp
780sDrZtB/+7ERX8/YprQp08McpLN61qiPiXLLYdfX8cSjTLtt/8bmjvEwRuqJyUogQ3NLdlfcci
QXh45EG89NiWrkCT3ouY7AZyelT/1jRX209adMrfklBd/drZmSIRgYe+Tr5Zatn/3EHsFBw9XLty
N60IfvkBeNvwEsNwfh9gvcWAcFLeba+ZLdTjxSbwCvQf7sQqlmbuKEPypo+6Nwg0Wf6XE/YT3egQ
AOHUTQA7RnRUzw+3URo5FzfpAPFhbtQIgrR5yy4Rkg9vu1u9NjRp90IG2LFUOvkEV3GsuuOWFCol
8TyMftq05KeeRBfuUQh0Du+tkgY3jjHTenSYsD673K5uAHWXbSJgY/0Sp/gTCj7pB1YT36/NDkui
MaMloRxxB2aIRXF2T+Ks5S9l4WahLwDlKWfmMhObXAmgVgBsdy6HK9k3VREf8K45K9IJsnNfEgvw
rYiu0HxjWBWK21iSMVuFPzaLje47iLInhdJXhJgFjFw9CKKT053YTy+86c7klgQm5CCFxSsbEWQX
qVaHcW/QJpJtBvMGYl7OcafEgcoOtQo46ALOZD/wcB7e4OalyplJyvBLuaTXc1LHEsWnGfY+aa7G
9Ov5OMgEMx8VotfMg53NeS8+zCaEI7XiQs/YXrEKQjtP20AcBUccDHs0DF149FK+HYxqKAIRjDkR
JwNssH/wrXOxcIqneY/YyI+eXjQkwRZhezsSvkbHGTVofN42QLHC/i4FIt/1R9sIwYO0oT1cp7Or
RlryBUy8/ZbTD/g7VIOMACCP21u0QPqSKxdKteR52eyZgkFLxxA0KwmDZs4Gp5QrlSIOHBr4dfZ4
PcqNMEvBwkBXqHueSIiyImKjaOUPUGP74zpO7xYpbiENjrsDJiQTMRv2F17QqAZMuUBmwh2BtZDL
pGKaev0L4CsBNc9Yz0Q1ZfjOgqPA/LbgGcflIeSOtsKHvUywxz+Lkyn/y7V714b9EZYaGVRmjpId
6pxYoAB/DQFiIgzvO3oZnAjgQ6r1f4cMNgnTSz6yhS+MioUY9IWL1IK1nM2b/A/lBS+42Yt8YvFW
iLU5OLC5bkIZH5tBCPDjqPok02Ne7+1nWcAouopSE75+ygSBS/KGYnj2LWBnlo1Oex9HaFRv30tf
56mi9esL07EkKCS7+WcC5I63V5mzA0fya1o0ZR/xpf+U5Q884cBdtEA1f8tiwJ3brRxV2LT6K8N8
z71S8pfNIdp5pLB6MTQfN4eKbDeUxrw/J0r/CwwKLGny1/Y2rtaOSrX5TcC0cyJL8cAD50RhOuPi
jE5VR7/7wAJQwm1QYcq6GWQ4Vy0x0NRpx5CppTGZ0RUAYS6D2VFgRqJRiQK/unvCDDOC/k1q1udZ
ESVmYxRLMzYtggIvKwCciJ+m3eslPN1nbEjPPBBpHKWGGSOfts+62ro12wQU0Ht5yHFHVohLfLl3
x87gggfmLonPUtruiBL7MDrPcjMGeoCHB99K+b98n8oTz9TpdYtx6j+sHPEG662/WD2PNCNUBa0g
qv60SSRhtwfi0clUJU5jnF5qPq3qw1r3yW3cGXzmicWK4HfTDy/l4uTkxEMaYgrcwjzJMSIgOiBW
Mrg+n9zopW3ozoM6m2coQnbT2YgIy5uKqFYHrVddCdR+a4SXcJtUjMiv0m6peqkhLu4Zr0HTdiQQ
Uz9IfuDTjqjmR81vGO1fpKTk62zsZQapKxW7F9h7rlckq8fpt2Jno1HyMRRC+3oGcuBkwaOsJt48
qOz4IgWQRJr9StAi4DsNsgASZ1kwDqyMVPLTuVVdcYZEg3XRg1i/liIEQ5HDMIDoagxPQoH0/n7K
xFYmk3+g8vzOQLdzyMMfBnU/PxnAuYe61P5oMrj837GI2D+93vKViujmRbfQttQr2i9Z7ArEL+LH
WH8xzC7WgTeQ/sqsWKwS2cfCieZ7XlyTeArKjEDsKhg5sT+wr3yBDkhdKMnWnf1y0xJuGLktuzeA
y5oqjfebL74bmUw79OSpS3BdqiTxgeq1GurcZjVM861n7UU14cKQg9yKGwibuNFjaE1+sx+L8pD6
NXfx/4jXYWAWg7veL6iJwbyCVqblE9es5vwfNEpQrKynOSoQy4/KaU0VdLxhqRyxtTMEJ+U8ROkH
qJs3lAgRzZYmGncrdcIYgLP9kctAmOsZQ1eHop6pa/Hn3qSJzNFYx66h0JS81XBw40KGGL43W7/B
lmn3gcvsmfZ3uxO1WobIYfQVTo/FHVbZjXGrezgxVH8/MLPKue8nxBjPmYBV8cI/ZFOCh4ySSPpJ
Yj1bOI2hCe2gzfnf+0H1l6UvIz6lYjO1zkeGrH71gSqYNsutpUJA0ZgKTg8gKEMiYOzlgplSbXHj
Wbm3s68GaVZozKM32ONH3Mr+/kOh0A2BGbkOhy14hipOoflydA4MqIuDJ58IkwbOt0WItKRpn8RS
t06Smj32P/0Tk7iSXq5OzuhWecZihJG3P3XKCzw/BT8+XwegEQQB3rCpVGJiwsmZn1wHCaJhv3Mf
2H79b8+CKDTvTHuCULXekB6RIKP/+qFbVpr5i+UJNBU+vGgenpEH7ULfELroePXNyoOVi0/9Ugv+
f5cEgOGadqc7fOcyryEEvwXkY6AQ3LW2t+Lk7c0Uyaaat8PM+OvDzifYd6H4BTeN/1GxyKzuKGTH
rKBfQpxcpusHpRRbcRmeDFRvA2zlqm0vQ8Ew/x4mKhXdXZcWyCzwu4zsn4JRPCS1tuMWtoQtOofx
0dAdei8JBzXOW93qxmodbFiww6111dS6lVKphQrguoVyQKxmWTIMMb3wbdRNgjkP+/t54ZmhUk8L
gNU76IOHTJVgCfoosCidYLlK5/IofFs9kLlYQobuvYKntDGOcMNsiyokCnImCehwEpbj+ZkG7lYE
UbFcbXvQ0nsw204ozkPywWg3jbKRavFTuUsv96GTv6lOHCWOoJstOLUsEtJyB05GWR7qsLOy03K2
zazusHvzAqbsIkuvLYCBoXG3POGKGGCkKvRKMnNnzQbBAYVbTao/f4R9E3iG253HXz+Q9jqnaQNr
J63d/hpwMXZKP+N0vqgfvxg951sf0KaULwB4mKMtYkzobqnsRg+mK1XyUC+cHFwe3LrEukAKkitl
xw9nQBYns4AsbXCcDx03i5dzQ3yw8G/HdGe7looMy8fOqbbl0LXfoqu4RfAmodzgcJzeywWhIUUJ
AtgdD9UWYoQWKLwX8/KkjPRfjE3QTb7F7ql0D84rgKlkycoUg/zrt4r5N12j0Yksc/tqtBrITE2U
f61nFTOGKHzwQjrREtGrb1vtBgl119PhcigZd533IwT898Vr0fBDMWKKDHniyf1Dn5NdFldvzHHz
sy3OkymTYOLeQ9KsjMgkC6uOVXeofjQJvh+Bdpgoe7ulaCTS1GUWRVh4E6JaiMfJiHaW9G5KlWQA
ZJNBj0tJPXtQPgJDmrc0pxomq8XFaJf19jRJ1IgF/pNTGWe1/TPY+9rcfOPk1HuZYfR2pAtuyE1k
p5UtyIQxYuoWKbZRGgjgX+QaXW6asnAt6+9HMQGmbsF469w7ghIr9pfBk17/Ywf3JJhppbgzSMSR
rjzvevEBeDRw40tAmR+IBOcThamEELOf3Nwlg0tPuUe4P8LG67UycQHbwvkv3dh5IGf9vRW9s/X1
2lYhshBZmGkGVuciq+mZud6GZm+sBs9bLVA0I/XaQfefW0xiWdnGqS14ARiCn46oHOiJuhjIYtVl
13Pbn/T8N+3h4ioQAd81pPl+mrRVwnp/HTw2IUefkYuc+mIswa2RCMIOx9/NPAyg4DXmEmP0C6ow
MQDKOM1ocS4mc4UjuQ932sA9F8KGaCEdm/95wQbAhkK4osuPMk4JARpDnR5Ub3bp3x3fHq//Y4jn
ciUEWCycRB5t/63vyQAi4+e6psEEZasMUg1A9/iFgpRHo/Wt9t5pqSe/Qri70EUBJGQuJ15v0nG6
hwGT0ZH7CP4kmr5bU/3WDRqXbZ7NJXXE+sQfNZAKhgsFDnKl8pzZrV8Rk4FgisA1aCIIrk7ZkLkL
dfwyZ6gqS//1Nm1OAPB/L9cl6FjzvT4JbdZdA59rbQxD09oTcVGp5MfTzn1Lfpl4oHlkH0JUCiI7
vEz08Hpq8DHb6ofXw/DVMRFILg+0zWF7QQU8S4unuOJnJog7k+7Z+D+aOXfLLXv0KpOTqvPwaGoO
Tw777cQpK5VXsaXWaOtDeDbqTsFWTiqykQXHlHFejLyImK6Z8Gh4R7hT5qM4HpLuxbSZGB0OhymY
FMRAPtEc34/+6gREWMIeSe/Rfwlm2u9sIgkRdMTFMCC5i8fU2FCRejDoEXPU/vivUC41WCzM1ypn
rmSvzAY9NsOTTWZbJeyBkHP2JvsTdueYRLlJfTIWrbkErONivIbaHVg6PIN/yf3MhguXNCvGLc2I
gWRRULSWclFE9G/aGKD0NDGE03VLNd8RoFEcvC0XPrlRisVAcuE3nbhOfytPFGTNtiTP2iFv1aVh
pKFGE8kU/aJeuzh5LnZsChRJxHe9TT0lj+q7IRtxUyP9UoWx1UKDHnKceqOLaneXNm/PL3I1vEe+
VgXVYRPV0DeODMiDSJGaZtW0Y/9bfi7DGbX+wy2QhgwjOODP+FdbvQW1vMOSM8dn2XAV9gAcdn43
WKLu6EnCVfLGNt5Qsb8fKSS8dCa5AQEdwMklTaWVPaZzHATd7vGJA5kB0aVMU6pcvU8sdIeEAoEm
94HZkWtNy0JjgkNQ6MWKetF+WCXZXfh+YTI310cSx0JTfbg9g7988WFrWmc/8erS37azawoGfKF6
IcvtI5KYNy2SlYDtgnpnJz10ulMZDqH+ZblAbnM5ef0MzJU0XCTLE7PIDX+X/9t2Xy4flPyPsXTM
ZcSxp5TAwukEBHl9ssH/H/PBdla7yyuXsMaU7IB9+ZH3MYIWameeMK8NLojGKz350ehiA+Z/zJgJ
OTsLFLwKJ8BC7ghbKt+/pjT1WBdSwg+TG/OxOep1yvYVAWfp59TNtiemr3r/3YWltjEqHR6t+v6X
N5J6HToX8ND3t6hF1W8La7P5Y1EzoRajJntdjAeCmTfFb9fAEBj8QFdCZJ1NeJOQZ4gxnSulboQy
wbQr0ytwo8DYrNx5X/zIm9sUxwctaq89+GyMrDNhLuBuHpEPKyzVZgu3tN3yo9lcecmR2VApBc5q
MUM962I/K8LAvmNZ/61aI5en1yzu52SQlsaCVKfA7Am1rQ7hU3qLZQA4B+WztWzcD2kW9xxIHaAK
LXFyHF9RrluLkm1szyEcrdyylLgYMKOZAur3kAh00oq4M/YL3Lh/82QXYtqDO7pXuoRFNjpK57Lc
NkQT91EFCT19Sj12DjvjFclHdDPqe7xN/WSkvGkp4UBFkTdjrL+MO8jObx3Ja/YbVcf0oYpH5wWn
7Eic5PRD6iERkkw8sm4v8RCu/dqoHmWNcUVx4rMaKuW1YzLJh0rFQ0dNBNS3XHT3im8DAG00oU6B
xYWussgd2/9hamLn7XZ9bLfStjJomeL5gspZxvkvfDpC5GT+ZbOrasifM2P8FoakFoAPJHvJX7pR
LxoAA7WK7eaZpMMWSd8ehzxru6bOW1O4YbiRvSnRkoZmuX+6UkpZNYnBCJTpmW5ys2Fc3DmPcaLN
WBDu2t1ZgYG+xrFzFDilQo/0H6lQpRs6pbW6oqtspPnQEvlh9b4fb+Vwu05Q7xou+8b7xkG6JTGn
CceELfjTkcvN6eLLU80dnl/3slDP6zqWWY5X7sYG2DZOHoUYdkSIwWl3VeYcnrU54nw9SZki+ipK
eEQKLC6qmYMFhGFGAdDWFBiEkpAI7cuA/9TuWnt7kxXh/W5y+kV7tveDpGo2KTyB3TPEYC7MdL5s
H5nPEVOj/bPoWZWMxXzAAyXDjCXr8781XbCcNoRjWR9C2qczgJkT9qQGYXI2qg9wSwFyUptblDyl
3wdpUZremUqvKZkLlxcbcwobVhJBm0pJOGzH+HuL5AcS08i2wNVE8CvnVNilk3nQgm/DwqgC4oKO
qhl7enKGcJPLiYoUmqEL/Gh1PdUDezFtv86mjQR6/9PIR3PIU+zSfEaq4nK7zn1TARIqnH56SCZu
lSEJsEEiXpipoLZFSerD1RhRJf+7sYUOpg/I0jkSMuDas4fwSOAl5EQAMQLZ/9M5aoiVD58dJqTY
RA2WbubvjmMiut9QWxHWgfNQ2T3V1MX3I1XVce38CYAVXhT2qHp3M2spJuWWCEO398s//7XwwIYS
zZlqGWBt/RJn6/s0C2aX1VY8Trai0a+1SgFQ5MkFG9fPmq0fmgqqDOmKkqrhOceNwLG7+dKQ/POS
gE6K0AnTxFJHuFhilaGnm4EbogbCj1rS9ly4IlDeDDTKXy/jofiwXCtSM8CG6GW2hqC/zVWMgWo7
lUf1z1HXXNFbu+ppWLk2/k2xFrWpKvdnZkNtd1YxAHC/NTmiOXfqs8FskOuFbZVDNyNppIbSLu9t
7eGU0Si922rLB1HY4hhUye1VOhLIMARu1mNYglwwHDcb/3OyLf4IA8OL8EJmrp4vBdcG9wjmFsId
sPnYqh4stL46xqr2hJ66J0NNhIbhgfuIOUe+TS3XHLVGE/85bzVCvxabLDPGmmWiGiktr72K/Mjm
wDePk+NEwEUliZCJHjAZ57pr5wvPw9tyrxqAciJN8pV4eWZl5Cqyd0x9YAqmCFDM7L7ZNS65IA6n
gR80KvjytOkhw9IF2TUpLiYUay6OuoqjR9deUH9LIF0jJ8qhL44NajrQe+iC1s7/eusyhO56rv1I
CNaYTPRF8Z44P5FA1fFGekbTQC1+x3WqSwL9aB+Yn4kjWf/7mNyVBf7naFja47HRfJrqzUBqvZYc
I6LOEEiK4XtL4lIuEYuwkXXawTBen2XoUsOhuwVyu5o3+VHzMJ3cMhH0kOKwO+1hfIw85rNNgQYF
vuNxaVPfN+N+kvwo5wTSQk1gcR+RcXTsiCKmXewkUKQkiDNIzO9qYsD95zl1EHHAwrpcktY7akqu
B6LrXyxobHQxnAieWYq34OLq4p4faq0ReiGLZabuu33YW0m82R9KXx4B2dWgLqN1XnJLV6Jtad7Z
xF3xz+tAMPSGNFwcPK841UdtjOe+BZh5gdwe9MEHj0kHhCvr1gAtZgcUZ7OqWK7RDgJk0A36D5nP
nH5a81YZyZyfM5fS2UD7VWrveEO2t5m539kEMsw2LbUNtxKSzBXVGLqAgKf6+6LKDipsbLj8QwjH
NOm1z6t4W/p+s73D0j8/tptncJ/w2m6rVbZ0c2jhBXUw5QTgG1EYjQYwURidlu6w2MAqTeDdZFHm
GnuTc2rbmBkL4xEUHJ6yvAd9xRM/JzIclOi56p9vMKC8tAbTNTjlplcRT+n/umaNfseOu6YFzSWf
AXC03cOqFJC6Zy72ywOI4kVoxeL0v7W1jKtXwP+fZJj5l8/WvpUQnJE+PLTEQrTe+4bTbGelBr3I
zIkcGhLgVY7+xWYTs+9FmnsWeD4wEENiWofd4ndwo5HhNZAwZFqT+AqQek1KuyncQW1fr22vsayu
DbFYnteztxjjzNXYdXpNlOGXJd4K0mE4HCjSo8DqSD95WoHdc7ABaAZU1mEmuGd6o9uc9Pab7cBz
vGcuQyKsHcQTP+GyQmM81X032HkXUAR8X2jYhNOD+YulNeHuW2/buJnQmXBg/c4u7K3SzvIM24Ih
EGyLb+xmr02WjzgVutEUpO/YZ5IwMyRZjE+ISeNWt44KhCkNDucnVKH/b1ZyVi8LbKXEHOpCDNrD
VFH1hFdLXLPZVxmIE4Gv5aFa1W2muyqb1DgAX5Ic/CqB0AP+bjK9S+FmyUTzamKUKME0vlV9YUx1
AYl6abV/DxCtbS+RMewtRqOqFdEhQXaFZB/bt1dEU3oz+vqdj9RRrG8SisXK9Dw3EdDtoA7FwtKl
uGBQN2Xmo8n95evpk3qe9SfvxS3FFKByap3dcryuax0jiovsoK1QTF1SvbTo3SweJafrsBAxyf+B
oXz7/Z16l3OUy/IqqTFbucxKAgqDEJdz5ykF4ec0QKdafqBzY9r/nVaR3RPKR/up6jMu0IpqoxOA
TcOsZWHrzr+Daul5AtbXlxcNcOmNi0I2MuqBkSpEZfulLZGeXtoU+GBRAJlwLZuLfxfl2vxKWgBk
PjbvbanqxZuSnwg/kvbX3yG60r2fxeIPMcOxzQOn6ufY65Aqlt2sQHYVglNkf8Yt9Dl2HUU/J+Dn
VZ+NIraXoEl34OetX0ftJL0eVJJyjrFmHpY8uZkCSKqjSeFhAxuxzYJS+i5W8LZZQla+q4y3CL4U
g/M2YB0IvlBjhHJxGAT89+lE59xx5WhRGenc68ar4VOUsmfiMiU7TnOorUS9VtPvCK5rRZFXSC3O
gRbz7gKiwnjlusVXEFv9aJq/6zhvTOHuL7cqLQE3O04r4XbgUzj1yWrjOz56kCSibllpkcWs6e5v
6gkxqKsp4u1UMDaGxCj378IPZOq2Lh2X52rfH2OTC8UBx8vWSt3EqRWml4t9V3DdoDAn7Q3JbLAa
mPevwfVDGtXKblJ+FayXoSJcC3usYdwNdHarCCZ/lgDB0XDmHOP1vFI9WN2HNAliepLxwxkeU0lC
gmP9HKdSUjlpGylZ3rBIBp+iQjY3pfu3M/5z37E8TzEi1eawXfDuNAocpUO6cZOvmyHR75zXvyAc
hj3gzfKaQEnmZV+xl7sWng0NXstPmbjwzKASWdQxDCvIZcgR3gTnBXoJzWXXUdyPz5oK8EHv186G
e3ANn/NyOzkTuUl+ZIKtgEcVW45VtBEtS28ngDf29KzFPvJxAMAlEWibCjr87xIzombRUBRTelDA
n/yxCHR5fvO0vugBONnuhT7naNpNB6gFxRmUxkJuVi4en4u2/6m+IAcazmzrc6Vjzdw+XaqJlWmB
ljQ6yfVjFzOGIyn8VQ8wK2d/FPVonGBH0Yy+zWylmYIxx5m/FgxGB+Xks95J9Rgcqehf/QBGtzaK
F4SW8vCkJJyumm0uS3aXwwGqdxXx2wo73fzFuJD8eQNt33s7L8Zl0pDwUkmlNsFckYsmQQKMt/E4
cmhe8CH+uTStPpcUlPphgoyg4pEPQwq4DbXcIl5zY5YP7CUa3Q5lzrqldeo39c22qGoOEFof2SVO
9TaMBAb3rGGHR+4kJDoyIqUB+P4RMe1yYXbLANCEQemNPMyEWa7gZK7Pg7lVK48otpR4sNrKpiDr
aUPaCsyUNdFP/DcARhIaYUsONzTJ8ocrm3+raDTr/RObZvWOCVz5a8womDdFJuJQbkHIKBz48jOf
mEyC7YJ+HY4bHzf8J+qLwDLZhuB/X5ZdwjlaEQC8GSxpiK50Pwt3tL/x32efaaFT2BrwheYnS8Ek
Zh/yJp6GakSxQaLcGQSRhedtsg0RD83Othg5AuXMYJHDRZu8E5PnremcCyh7q8zGEFjw1ruReT9K
/a9dWWttN+XviPI/Yx2EAlsyyXu9aEdmPESXZf5Yzm6rh+Nqa4wpQg36fpyYlhP8VUgi0uabI99W
tyU5OKVLx4yx+gf4bNOe8nQGCT5inO7bJ7NEPTMSZqq2r5FrbZ3TPNhCXiI7wpjRkbpxozzNMISI
LV1acgyW+CrDCSSEoNHK4rqQZ+QSfr3wYoZ8UROsDtIq09Uc0I3rWRl70B9tscjfSHI7tY6956or
PLBfNHWz5gBbFM9UOjIKolfbMplBrldXvRW4QD68qmk5rKc5v3OHhDcceUY/NfedQzAk6CffljHe
Ihw9cr89qglhx73AQVB5hRLmjbwcCgEFxe7wMmswHzXen+Yr8CduND57RDg3/LdnPj9Q4k9iGdli
1z1VKmEiN/6omv7c5ohvt6Y9r1cg9kDeHilKyL2LJDh8j6AIQoADXMNei3F5DAw2wL9lg4S0lOqn
LPYxQC+W6WlP8Vue4ZqlDF6y1zRQujMrN9HlGZcE55HSrqKhU/Wn5+1baq9BcenmQL8DWnbjKYPq
WYAGeu8HJwfHzdCePuRK9Oc8enOpmlmTzWfu3jXWD88CE+PiFadKoD75YBaV4C26VuNDBFHVe2yS
dP2WKGdv7FSOZsR+kylyNwRphCReSPaPqBn9kjTZHxmf8BXawfDerkatwJyAuVuar1L45/dJD3UB
Tpo9fogbq+ffufGogA7LLKKu8/IK2xLWnVeyYnptMI9gbEwIoLb5K3FIHXBzWzvKzdncc3u13Udt
GlXzkvNeKcSD30oRq35AuCNo/tnxCjIpnTMGHWSJmhcdW0kviWapeJOkUpLt8TKqo/nqjIGfPVaL
g3GljTl/ZxN6ilTHAukdF8eihlhCi2Rw7B4PbSbDv0Gzzsa+m5ZdAJlKwSw72Yaebk+ZVGIjjrXs
VYf/p9bRkCLwn7dTGUXOWsRy5sXSuwTzByWnzgsml/j1lOb0737yRVPD/J6GZ4X7aZZ9dB/wZpRN
tinF4Abt2N/njaUeJLxtsL8l3t+Xn6KRE7JGuOjAxMnQ1CPCMNHu4qlD7AD0GqHozoejpIthblSM
UQcdAkERY1y9ED51uWGviDjc3rZhpIIJ9BjrVBz4gLZfs6mjXLW78K3Ve8DHgro0OoKHWNkYyreV
dFEG/VJw4SqDoO1SLdbc/00JFMP0f0LAxiaMWLuYvW0GGYob3NafHbGIMKum4saZwRrZyAokrgLD
/UpHX8v84cO0+U8gsdEGN6of6pktPCDoktpKrmQecxouXQbqX4YprDb9txNzIMOw2YP9aeLKSeB2
uY7jg16V3L15RY8/4EpBGFOqlg7dzAi+S34ieCf7SKLVz7JSY7Tf19s8KZl+I5b3S/297oeqJ+3I
sQFgO0xgesu+1MyAEcvEmRNeaRndJfY3sa8Wli81nbzGjgQvovk+YwO0x/CXvZ+nVA++Q+dVDvqx
cYjJIYHq0L6mFFBxEQ/BZXwDS7wrnXqWU53Tk3AgBl0Y0l+36MkGH7Un3fWFL3REbiDocc64rVe/
/VrdBoyKsFdLviJis0+FV3qT2tvXxf8Poj+I/uK/fPzGvTAry+jKK40sBtTbozG609lLddGp4GMl
fvkljZivaBqnei4bl4ASJROVWUfqJeBFu72LvqNlAsnIrP8WP/hFiJ9874E7CRLWsFVvwuUUVovo
knthUhikMymKbf24DAehdDkRAO3uhMdsORpCfO/SHLKgnRkpwu58ouncmTKV84pbW5/SNXRJPs3m
hzzbRqzUWnj2NC7CYJGecYvxjNYKiGNqjZfJecz28trSLqj5VcwD40IajNUE4iMR1RDDCT2y/FrE
OD3KD7w4tETrbIZJTPxM06yMwwKvRBGYlI7ZAlvpTP9TWjK18OgN+0nFb0UZ5twTicSSMaWWaq1d
jJprus/XAfOiEA/xAWP15aOJpp2sq1TcyS/lUDK3Xrc3pe1ToMYMD9/vw5CxM6antZwmytiWUdSe
TgjbcNaI6hfEuJhpBCBTOueOpGQWLv8S1lQloV/EEMDHKk4NiGvgUYvSOojEzkaAb/xQTdgnJEYU
P3E9hv1SqNQe4KpWvbIUCP0fGsptU3k3T8htVK12R1xyJw26izQCENUw70fIWxKHk0H66/I2GRjY
b7J+XVkksx8eSTkkYd+T11n02fcWz0CNv42LsT/MTd/YevnWFfxF77oG0/InDwAauKrPPTtudcS1
lPGW1xzTZird9urvrlDhQYduWiATMYPBK0EIdsiwQOl44wqF43ZoRhU329Icvo51SlPU+2v99itR
o2t8Z43ZwUG/8vJu40ZxEm7UYbaZHDMgZGaXblW6FYK3/vNcJOKa4RzPPc6eaxXxnWTYxnzc1sgm
VcnNu0GCqX9GciV7OdAVVgwChMVvewXcmoFNN6HZhanDRfkIvzJARduwCdYVqKV5UTNKhmIc/zd/
cjjJG6UqdJqKyIPUEQp7gOf/UlIiJtxJEw9gBu6NF7dZmGnefQ9m3Cye2LoR/GlZFHShqg7IOa64
0uaJ96iwHI9eK/JZ6Dz/DY2TkJclVSRfSabX9x3ez5VEolSaVm2mV0ACIsmFl5ojNOSCMnL4ITzL
5hdB9iOEvqLS+Fn0gwfKSkxKzezi2i6XgPCJU9kJDh8FvHL4vPYdGUF7NffGxJNukzvlcskaS8pz
WcI6ucaWOTJczHKV+B1l7S97RrIfpD+ibQRhtKROBQkrVrqsZcp9X4ffDTc+YgoRDdnQYbWbEbwP
pcAFeNQeoODesmcN8A03QnT+BQeuxLB0fArDavd+lV1hHdhK2mbWoqP/Yj37bcs409K70zDwyhdU
ETkyFyShvKp5LJwRjaUDBQNV8JGqxPLS5DinK+cB6MENu5jCcTPVG6h9+bwZYT09D2QpCRX7OFLE
4FFNO38bL4be/nhzRZq5/7Mx68MVPBJwe3/5q6IucDnPVxtkvAdBWn6+vB/pcGM+ZglkFx1uve5t
3Z7pkIxhClXnhMgoHtyYSMC79Y2rVZ7pKUkpaXySwJlq+zQ/22AyWOow/GAUYl8J3b33wqFNCxfU
JSSqzYsT/EoRiXiOyRoG7xw4QrFlNd/as22zMX4pYf/SBYzC3yVcyI7+/qNJ7qxvJRB0EJz5ynnJ
XSwS+Ad+4RiG5FVhayXJCzzKxI1JUlsktKptfEOcxqJxyWaDjM1BMoIPb5kUZStwRNUH5IBOXaYx
AvFVnPukGfNmyLwAPHMmPOe0IrV+fY7onyypWofyBSQ4fKD+x+fTQoUyfMLLKqbSg0VDIO3rzO3l
T1FTguh05wtJyFMlDVD+w1iKNoD7+qfr+8GPI8jEZpwzBTHqqGZiiNRtMHV+0trV1vZ8QVs2o6L0
poEi1xXQirwXmjviLo5DECaI61N2f2K7zsQLRXwi7iqP6FyaygznGxiRLvurjZebSG0/xBgYuA4D
7moRtFZjJuTEMbj62ch0DbD+t6WYyoMeoGyI0uP8JXvFiFSa/guf+MvszXi/FRIzC9+8N54qXUyh
vXmeVmRsj/HTDSYr8WiYsWpGTpmvdBYtNz6zIeqEQ+qsyE5dYuKUmIat2ELt101bjWCluehSefi7
VRnVWu51CBMbQYf2vDc/5nRUXVsEEhKC8Z1a7l8nIFHHDX9wwyEm/igP92A+1qAlP/Czoxxtcyyz
vzqlXM/5Zp+Z2GrTJOxMPIXbofAwnCwZayzLB+l1wc0sD7MzIudy2C9pzrwI1nIgwj5VOiuCrys2
mkI5rj/mXhGNWefzW6R4/1qrbUYg7lcy2Gjr4x0zrE+d491GzRJAnsCBFD2lUe5FNVTyZi2EY65w
5xaI8ffwQGJPX+EUkrOjLm+jAKvs8t9uPZWkJHYsYdP1WT9juIxXlhPDLmXqaohiogmXKM4EVIcG
EpL2NwIyfU8eFM1U6t8/YWb39BS8Q6RHYZQwdMcAJgRnRT0eGbyXIAHwOGtR9NyE8gbpKCSlY1ZL
7sm94Amg1hGyNGXczppyYnjaVuufxbb0qjDnFtRHyuejBHrK05r2RzPpmaqkfC+03hQoOiVnV4+L
pZHexAzdP51xpNelQMxyKBaCvaOeGzxepLX2ZUTIYmUjbQOhKIB5bX2BEr9ViHOrb3DML3ffjl/O
MzIQNUbAXKiOCdX7g8FRAVBZjIrxQ7Y8WplGatVWFAhwNfVK3DBNd3apVNSJr07geO0I6aUtDnzi
N3kLqFkNZ53vVLMgPjWlI3k+CMJ/8AZh6j3PdVPTqdL5+RpPOUowREc8jxqoxwDaiUCABxN5On4Z
hbaM2axyavrLoUNQ7ICRl85b1ZB4+Ep6BX46eXl/lbKP3I7iFmNaZiBOvxHWjMwYNDqjup265isN
oseW1XgglZT/QiUnt0Rc2bjBZD1E7peGPaa8kEbztBAzC0IYHgUD4TjzeDB9kSMy0bfi6To04/MY
wX9qb6VaZX777B5fqZXRRN8615mrBr0OSnzfLoT+VDbav0tL6urH7zABgiODC6U3j/PrWpYCuaBm
wCPoT0XCmJ9fx4gN7qGFLkKAF7U9eolcROir7QqcxGnvB2RPwLSKkGoHPDXUXRRSy+RrzkBYXKxU
ydhTrg3ptjXkBF6YgZtm6yLkP+UsAcL78fa/uZPS7XY6ux0QtYJRVda34gngYLTI4z5Yo3C25GIW
5vg0Lbl3crECv0XE7HH4rmjYodTIbvBNt2FWL+TOAfiuwV2kQTbUlMbQFhE4X8ZtrtrVIZrhrhBM
zt+8BQqmgLT1yLJompInobE9AYA5Bs4sL19QArRwHrmUtkqCPT3U+nvwdwHS0Lk7fjduhS53oZIo
n+CpUPcWWeBvrq0pdLDFJvcCFIuT+6QrHT1MVFaCM4C/QxsBu8dkxkKAkjsdaM3WQnjjwtqDvUpc
F5B8Q/D/joLID50KmtUJhtoHr2tSnzLQcx8phR99QNjPcKRRcO86OaGjwqHdZ8g2fpTx5Vi1LCZU
rptP+vbl+79UFSIHm3xX2s6tAywLEWlM+yCCjdlZSeviyiMKw7L65OvhUGDxkkhEwmSIyGqGDHjy
/ImPXzuEs5/PkzRvn3vShJM97nwM4GWhiLiyuB58hHBiEbGcms4aMwSPk4WhSR5pKFDE5Io7satz
VdfHU/1AY7WLLQPE1oprOPGmeXV3avzzlB6x6/X+axhtTfwB/beDXS8uyi2D4lQgqp9cHsQP+ZUf
ncblanYnRVfQb1gIo6Zasso/ET6kQWAJ/SKUbbbW8vhwpOPV1JOtxmHvS4z0UJu/perprUdBpPWe
5DFKI8nnKfJcLy/KQDPyO4m9BNxKYiz9oT3c3Q96JsO2UR2gkx5xqg+PHCgbadFT7a7h3Nb9IB5r
TTDSe47CKzDH1YDEihwTxqb34jCGcXc878sSXVzT+rsokqqUbz4ZnPeDPrS6vVEmvcKURcP5CibV
PDgO7HxzSF9aQU4HiFTED1RPwvdpuqjElNcuKGKHRs+ykC+a43LDc9nU1V3eBKHVu1S9oOJTC3ZA
sGhm7ZCDfl+h1alc/oHIiI9K9o9uxJAIFzi+jxXeU3a5UIEYZLfHe1SoZRNO4eRUmgGRUejpseMR
njMFOB1mMzNfS4uYM4w8YotB3Zic7FPz1SA+a4ia+9LW47Nk/Br6hAuT0Y2y/A5G/DG5Tv0WB6Vb
iABSA52OOvRqddC11laY5HK8nlk4OJMcIxSXa91sttNAP6PM4+ZTgjClCJ2KGMPh1T32VlOZM3MA
TJnZXR4g2CHIEg+TuHdg+oC/s05JqJr1FJ/ab0cmWSpVNzX9wGgPWhg+A4FXKqLlJxtbaJkcUGOk
hWhFTNBWkmJbFHashj1my2Hh3Hc7Al3gHPBu/7j6fW/hmqkVEFSVs4uhyDKzwgkXtpIvCwHu98zr
7o8+KZaaC/jSeGLHsPKZs4K8fUj+Rnri2vNsAVd9Kxoia7mWqcwGCxDpmX2EWjg2JsiCAvdBty6f
Xs/a6n5EqWMiSTA8dtYn4ApQGD1ixBA3RBmSodLj3oUY1Bsqw2mPE0+46Jeds2G2Me6WW0vS2UTf
OPf2Z7LHxVre4GkmoGqA2KepZILEPprUQ3CWPmcLyGWjjKoYBnSPm0YB/Q9ISuHcUcpkBV+rRkZb
/0T68orHR/vu3dzgnxZr/eLFCKSPF+S+C3q+dlscDnE9fkWNGLT1yb1Jb0CPYXirY+twvIWfZsSv
8xtNdnWrlIiileLZl5Lhb1ChNNONlLsyQGmBku4IjX2X6cT923THtEqEHDHZiP9FJO8czSq3ZUzV
SITT6UfuQN/7edqNoABW64L61wTq3NC5EehyvENn20nWusJ1uMXDxoB4qagLhgeRuPUnmhx6s+dm
yMz23d1uJ7YFUoJzqwlxmw4M+KCOBQHRUofbPINSJHL786k8srTSbGZSA4wJlhLFl8vEZK0CaHmd
7B010uSocNMx2sf9ePMtNXjghzZMwjF1nfwnj5HVWJaoHr9OL0YS2hJLtn+76Ku1iwmn5H/TvVIc
kZTUhy6rXBL8UK6a9UJWzUibBdOrzNZVgFflQXdmjQj9nqqJARt13RcM5TgjnfWjdFcMncz0dG5c
ZI8uT9QUMztC2mbjOiuDYc9EDlvfeWDd8sf9QGgCUHdyT9uVipR1iSJymCrA4Sb0CAwdfqFNOwx4
HyfHZX+dB/pk/osslIqwaHuTWiB747kuOvlXP76aBARKXYPv4JOikuak3uPsNZbZfmQc49ZwJw0j
7zpUf6KqnXvDO6L0ePDL8l0adfD75AcWiHzVIAh7t4FYpoav1BZfhn6CV32I/K9M3fhpE+PxGXgI
47IMuDEGdKJ8xYtW/d0HNrMVzSouxL7s8AiTYHBUpunmIMFgF+nS4n8uZBpMQ8BcizYJ5p2+Izah
2e/MBwU6OA26Ge9f9/gW//xhnPG1DiuC2hnS7e3tYARJw9P3sDprv/uu7bf5kEoes1qQ1cE5/6wu
Eqrb0vDtpHHlY8sQbrQwdZj1hmzQeIQbm0Bswcna5ik484OC+hcZFvtQJ0Jxvh9cFzDoy4ODBqiO
+NxCsxabj8SDGmba0S2EVSLrjXt1U7CEplxD4JAl7t4YoenJhCcv1DEm6bJo5QiRv3sjHOtvziNY
7rXNaBB6CX8B0u8kuA9nQff72MwGqDEAqVdE+oxm/waHBl9Y5CxGC3TrgU7LWC78QDpcxPVglNtk
DNz9NP7RTq1sjO5X0Ye2xgxpObzhsmfeUSGR3r4txg+G8j/o9dzb1EmlkUvdWH90AjrQ7WoTQiJj
//YQaKm0tsY7yHnrk/MugrrfwGRwIlyOKASH7P2fBRbDA/6t9WklMA1njTMkeBx9fjPVy4l3WRT5
8e1zJxrJEw5oVRWBkV4Bi4ZSBZ743TgQPBRVaiW5++DtDumfmRxaBZb+5rIez0GtVKdlnC2SdlPt
Ys0Z6BaivHPEl2AhHA+kBqKg+noZ1cQ/1/GWsBwQQU/aqtIiU7/bmHdni4AV5j2NxY78XuZRGRyy
GZdSiC6nyNh966AG7uY9r53KQyPf9+G1728IYRnJIzRU4qgBLMrKeRIpdTjXiGVu/mIEir1u1me1
QFDd3qQ+QLO1tgcEWeA6J/yVnbSeX4r1yPMzRy/NHXWepdrEXyqs0BNXUjSJm1Qtq+5l7H5zk9hz
iWdybKtYyGzMyHVse6xBHvqpo5+9ARznZbYVmNidxIptsUS0TLPbK/LcRv/aDgXjjmO7aRO0KcOl
Lf4ekFsCfzGRblBdQX7/PjbgMyk5ypXbFtvd19ol3FTbSoTnZyD/Qd/9ewI+pKBY/xIhzmeJQIlV
PmGPCnmf7hIokTA3hrNzOROZ22Sd85ht18pIW9adIVAZDriU7l7dFWGIN2vUTXIWWi/rHlwLzXma
lzFyculVsArrSFLMh1QqQwJwz7le37AEPt2fHXvXbG5w3MWudAcUdZuAn6O56Q0uxDknf0QCiMKd
fbcAtaZyv7On/1ZrmchSKqWRchvzOpebUccUjWIXvOC01e5qswPzmsPZ7Co7WsB5OuH3AYZ102li
i3wZuyw3i2pd1tgonq6G7M3jpaeV+TOxVgOi17Jh2dsT8e63WVRTNaX10AO57rUoHoDgBW0F16QB
59XdD2QuWqehOEQQ9Le/OWtNwZcmLuYBJACja5dLpiWTc48zCYjVxp9JV7g02L2gSEnjxwZB2Spe
4a/JSCUFUXaYIRzPVFEstFzmGrnHzl2Q+LauzprBVjZS0o8/7XxwCQAYBT2jQmQeZdsAx+bXuya4
eEjmIu5IrRd+e3Ipoxnyr5NuvsaR4ndDQ5Si0k2FXIz/coNwTmEtvVoM5XEooNBY+NCInWbgEjXk
v1Q11O6mq/hhgHOEOW3zj5BUU423AJODrF8BxwQdDvX6hB//fPmFe9QQHehVh49R6cJ4zGyFeZ75
tOjX9kICueYAmIHerzDMr9+p8RSb6aRj8Yj6MMl1wJqcIEvj4xyyjwQPN+n5pW5RMB0qQI9LtSkx
DBkOP6dJKuk6Dmd1YNZk4CN8eGS6gewqbKEpH2zegIzzvNxRauI9Sm4K3PzcYR6+uVo6lWDJlvMF
6vvVsCh7RlTsIDFQjU6qbj0yJIu7B0M4fjrMu8p9OKLjtxqHZb2/ZdYqCP7OJiccqV8TOiSLD2Al
WOm0cfbhxv9KMNPv6AXGW3Q79rMdPLRo+xyUTfVdeSxkqLdMSE0nr9wnWpLEy98YlmsQ2ynYInN+
KLhY6vYwpESCsmAb+6gd1tdZvOM2hSONBP5Vkt/sB7AJbkv8Zvt4//WIUwqCSRBAAPUXuw1sQn9i
Ig+Tvz6TZTE3uDaaJk9aazqRpFEZYQfKCHa2iIMHy7BYBlNR0E3oMnc8EL5YCKiAfjr3Rh3qnzMS
Q7B7jtCBLF6srp4urPxsajeiI4D4X2fpUhq5RI1IJFJY1klyOH4ECkOoum/WCk6BHjEDNv1AZATh
u0G7IeIpj0bNshCHD9bbsq9hAdiGTN0pEmwfVgmctkcTvui/CSSkJUohBwude5/3jwUC+LM4djWt
8iWhFdAG3l+bD0PgE3eUM4VQUKm+TmcU3ixSsFl39cmHJRIyOCiSJhPKjzBAf5DPvptppjVhWfDs
tXy15E/PHoMl0dGPtleyT+rTcOfYFDN5KSXf0d2K9NI5krCltfcSEu3NL4WnXRoM59v167+/VWTL
8amPFarpwQDbq2YQJkHhn9cr9mHAEM8YmUJ+tJVWW+M4wOE9NQ8g7BD1QYtsKwVQCRYXXxgthzZr
p/DwqHAycX1O4cui3dR8xrE+X9rXVnHvug+EQZkeKjbnR50rOujKBw3pIEhlCjlPzOWxNi/OWynS
7oGsgHcCfbxOjNmPrxakNxhhMcchX6LcGKBeHUjS4gVDaxOkZ78h5lA/SzLGa2FdUq9jofFcrDPw
R0Kbhe8/7YXw41pqCxBFVYu6PK+skZ6tAm0GlzNO6qnJGpCJJBG80ljzB3dJ4LYEQlIUe8gqEoVi
+ylBqNcBNlWxyhbmU2Y/CmWzuSBf6I84LF8OPFtPDCKy4tPtU+Sj8/9KVeFbFtN4jnm2BmMp625o
eJoYQZOtKyy2gC4jnLk4rKRpn8Wow3Q8jgbdjViRIz55U+owo9EPdRCXgbhxPMnGSkxu1VcWbVue
S+0ia9sKMB4ROWeRaaR1FcV+F5xdslSxRdOyReXkRd+KEOP27FsqvlqW/hq03Z8JDKTHicNj+77j
Ix964WP4C4vlBfmopyxv86U+WejpJZ1FytaL/pJhzU0VMmvmH1UyCc97kg0lWfCT4u7jqarJNGlE
RKlAGjjgU69XG7wbNeLJjQgYNDuSqX1RIaxuPNvPLR8INhiMJvlptB7U8z2EGiIVnc30ufC+SQ/6
f1uxxAkPkbco/FLBisGFEkZMd2fEVq5GecOPwgcXzmlX7x0VdY0wZmDlYO6urO5sv1M8mHOGhRuy
IlrZ+dYzXAx2AZOTgkhS9+8rzkcpisAre9O7tPnbArcF+LARmerxfZS6dkbNYM2hlSgm5R69FC8J
I0PqxuiHGntpPE/ATDEqbAaH7xse+/Uc2HNjVCD6hL02v8zidLykcPrvoPlyT4hjf6DNaoqnNigN
nLSIs0BfV8TQ3pngLGBp9eVSthcD4JWEjAht2d9z/bZoIzRud+lml6pqUj8fC8tnrMEPQzlpi0I5
1875QZbCZd78JvpjSY/ne9Bb8RA4UY/fHcTE8HMYF9UPwLdfnozOgbPEuaOVONmROXq232Jqka0u
C5Bw/DDQmkHVaWVDfc+wz2QUQ6kTTwOS920i29BxVdT7iPsiSSwvI6xgBZfF46NGA4weqGB2nOp4
zr1+f7AtItme86q0m5/S1u2M5U2TNW4W9hqSXrpGxZAs/U40CLJ+UuVVARn60G5GwppfTrfr0Mh+
rLM9mTd6ghXrMRQBZQAb/rJ5rOJYTeQYlmFFU3OtFV8aPDqhQjDNDYwReszhTcDmBCJ02vUeyq9m
Yknz4uTW65W4n8DiRR7do923YjFjb0FnvBk9dXG2K7Rd09ZB/69A36RKXhaF11sl1XZdzpefyoX3
QBi56mo8rAQpHLZ2r9Qhxl/I0ifPpzhKomL+RzqN8vgpt/23rqrVcIdNEgYxMSlOxgZmB6pXqmgQ
4vK1jsLQJe8hgrOh+Z74GsBNAz+uujiKCd7zjSrneZhHEnJjTX+1EQFxILo0C2doWkyCSoDYdfPe
doHbvyGHhAFUnczPDf5rkaMsNGUujqvjQc7jVept3iIavkfaXdMGQIM4gav+5T1G45U0TLPSQmkK
fNHv5Egk0DZSOJkGBg7lzRVGdACDXLykck77+i1L9pv9TZZYUISgE6u/HH7e8CWylsB1ifdUeZfw
DcV5m5znaY133GUfxdNswLOKNzcza7lwRj1b+2vIISFmWRYiGKsW6ToKyxHKREr97nOkyLQqS4Dy
P0xEgVSJHtaCIE0YHZPPoXBz77SdkqpRCSL5pm1DI0Ut2xPNEcC4Ng49TdhfisCUBq5KUZuBX5ZR
YACROkjryD/by6h5GX7kEDkRr1pBwTDz2bMTj+NzeMcqfRNI7d1FXIr3lc7bXlh/w4s3y+mCIhve
LkJTihb/mTlN75yvvbnL8Qgr8tbmyTc2jZVaWi88SB5e7Rmbc7TcogBdjHjGf7yk5E3qJQz/Tn8u
+tUD0xueSqXZZQwvEgKaU0hsAc6qt52jP+nZkVzZ8VUAhy6SUO7ZzoVgNzoNzko90nS5gq4UhO8Z
O8SgiW2nbSqnzGQPhSItCgCOkk8e6WYCDDWx30bjyyPOD9p4gUgVGMfLIwQ2Bnf8YLn69fCj6ibw
4uZYflXwM+JeJ1PEhC5Lo85VjP/IOg6+WQtb89oGCdDi/ilONgsGQMcdyBIjdY6Xst5CtSOD6tkE
vHpciYKPpro/O2hvNWfUnOWFNu2KhKkdKmqSt5YgQv9y4D198F3ElIFJRvDBdK5WmWDe4wZFc9EO
N4CtkZ5bGbi6EQwcqTKX3z53menGUvE8ldO97vafOh4gu4+EShanxlN6QUSGMOmhfuKNhrZHEGTj
lCmanarRej0/OUAelbwv3qqvciPXiPcDOBQ+TA1MlQ4SoyIQKrJLVpAhg6cHfOCvFhMwkTCP1Wcq
Rx5pF1aU/j19Bf11F+74beHDnaTkiJ+XI1tGK785fiwxZUYaLE+UjpQ0c/Aw1bivWP/O1DUk3w5x
jDlwpsjexFS4nq1WXzuL/WGe2L8B/TVKEJyyumrnGqPzvFAaq4NIs03qiot+hqmg5wBRNPzaF48F
xTb4rp7P67soLgjQIn2Porzqe0XfRs/01Ltx+8uX6EtdraNqayfQQg8+n8zCVgv8rgc9hvvL9NUO
G7b0Xw8vJtv4tAWI3JHu6ZZUGVaeo3r53utmigvbrlDlOoYpbu8xOCPFVQq/BXQ5RgdZnvLGYRgJ
/NgtfOLkiq7urXVDboD9VXEJR7kVK503c0JoyxJyF6Dhftp5CPwVYZZ/ChlGiLwQQ07g/EpLxlUO
hOTH+xAnlFstSlwBJrSxVx8KmBLT8Tst71vy7hN/F9F575/fEsngeh31D4DnoIAwSAQb52OumOWe
pIQIaZzj9YnaEjp3ql9nNEM8sF+xw5eWFrdh4kOaJ0tIVILtnhVI+H7HZJ8yH7dJQUM33aY1hoOK
6Nbm9ratnH+PlSfM8pgwt/7uEqE89PuJFH3GfKIhOlyiWjqQeeK291p3QZ7CFCGg1pR1XqOWfUbx
cip5UezOvYQ39eN2AvWBup+f4EtT0d9HJqu+1AZDe1XFz+I/EvPkly6D70eyGpEHESTHuPrraGzP
WMqB6KToW15oXPQIa+vapxIyZI9qJN+h7EcOft6rmdljhwbVhuZSniiYO4ygoewabHaq9xIQAKIn
G7+oTYh6e+BO5VKhrfyE9KCyGLAE8ND4UNk/UboKw/9xnJgtBqXDFwf+PRmY5RglNGsGy9GNQ+p1
8sUNhkEEDb6JoCmMwJrc8WHxIF5fwdtrq+iuuYIxdP2IvUcJF6iv++WOBP1NX40fQrp1ONplbnnQ
mFAOepNHMq/oUMGe4MDWmuzKdCN22ZEJdRkAUFTFoJV4M/x9rnyGDZ6uiY64FnfLVWdrqstR6IQC
7Ip7Z6BHjjqHQD/4YRQcE3HnT1xZYRunVA6IVk1S058I6kJkqRloAprg43V+3cdaf+LoRw8gysx+
EMkKwJBB6eyGKu5z1rW+n5lrdYsAeRbBR17lun0zKoVamKZdaJhSoutG5zn3w0VLCeMgOwvGEE8q
Bd6q7Xl2pxdwEuVlIMBJ5FZc0Y9HQsnmogQ4YZ17k2rDAKSigt1E+1vc28j7WakI6pS3TPk8FkoJ
Jjc+jYEWGj4IUwusSDDt4K1y4j3/Xo6MnqvfLNK3y+daJlEX+dm2KQlh5EwNVJ5n6eHIzaqWimGO
svq8K/oVbjmrVITRz0Ez2m3M+6nVbPostIHDAKMNQA82qBh3exKMFYFN6Fqzfa21d4ZFnGekvU9A
j0nFHJx6MyLr94kKoASdj1tjyUIY+9FHpMEnRyGByQZfYHOpc5+WV1iLiX05n0B8/Z175jptxnWg
7kEh3kuE5Zj2yZ7OgaFKI4PWdpQdswyEhFAPJi4ByDoXteBUIWXSvAPdDPP2YiWiXsptXXRm3Wdz
I8GFoNA1a7Ob+gIiolDGMCi0sLnp1u4NelPcHM7G6pSVG+HCw2KtoYgbLVG5URnawkpHtRU4Rq5n
D2gkHJZiAQVXyCtDAN5NAyfFSwsRyIYW9FP1/lb85s7vOhKtZnWSs9fMLJ2jNP6RubPssS8cvlqQ
gUZ0JyTsueXsl4yo1XpZ7lhDyOZdpHnvr3D6IQU3tQLnzi6bIURV0yKC3AUNX6VC/xMtfhaKNsQK
GmjMAoZ32BdEi4WQyonA6DHjYJ1fJew+5tZbw1peRcpB175luWgLuBJ7uuPKkbMUns+IYeWSqhD9
Uj/6HH14ECZY/MN6mKE8qFFOD0SsoWdHHDwpIODnyWQd0ltYw1UBaC7l+bnzztYKWPNkRaGNk0hr
mBmmHXsNbSlvoAKUXcoVzjz6lAd4XgeHX/fB1Pf+lo/CQHY16yaIclDVS+CiiNr24iEa6doYJNFn
HKEPhJucDgUhueR3FD4Tu7DNd5Z+hKmTJXCABxmTCCiIWjfMq2fae6WHqXyIqvKAJt0ne2Xf4bn0
I9JxZM9DFu7IKkFGypfpkgcy0PkhZzfW45PgU8CJgcz8ODo4Gf59BlsfvoeDVt0HitzhEgnsQ+Bn
9qKgz5x+eIhFGdkHfd2Mo1MlJBV6pTqFEEunsI2YaRYMA9oBBzkXuExExYaQuWISvhJSnQdH2UMv
cJPGo1bJhzcPTj1RSbEb84ALkl4qg2wxDlxtGu3d0OgrGRiAfeRh0pMWD0dG+5Am3oPNiNuZpWLS
MZe2bYP6xEzVO12pkGnRyu65avSJ1ORHQntJbO3s1zjKwhP18sVU0kxS6TzOGk6MzSG/Wmnf0fKj
e5bQ4oUTr2mAMF4qo+i923YLYSMuTQKbWzdXfqt1U+CG/TbaJZgCzMIE/u740ZNEmjnxiidUJkI6
YgTYVQdUx9kDHLsptWyKxUDqlGXxHe2gQ7kBZe2h8yfLoISTLH1Sd9rHjonPEj7AEweE3aUnLdNR
6CP5loiQMmi5cnwiGHnQxhJD8xbNUKsJ1u3xIf8uJs8zQZ2Y2i06V4+1Y5cWaP52XSwQ+oINHERo
L/okK+W219Z4vradFEYOjFDvW/IIJjOZ684jkQ5QN6AQv81vpKNzlVlowfaA8QaTRPVR8cx37RMq
FrH8M1+GfpAEHIMF+FXCrZCen1wfzXj2olfBIZ/NPS44nFrkmBSuAhRNhDGlxa6hm88u1QWPu1En
mh1CIeGaxqbnZAGpWOX/PtAH4DqEnvCTG0Ycciu5Q18JotJcOfZqf72DjwP87PwITZx44mSxMPKk
2zZ4HBX76f48tigyA6x7ECt6EpFRok9n6aJwktsTYipadSo1Dp+xrMKPzmyd+TxHsGa/0SVxoEix
O1shqv9Wsuep92SFMF1YjosGxLL3wz1Ze7KHsIGf/a3i61ruMoXhZOpKUBbZlyJX6fMV2JjFXSk3
8ajRBB1W2CPOJJz1p1h722ZlaxknXxnQ+rToDzZuVnYQELIZLMoFWO+T2DsgqArA9ge9qKmvdrqC
un6LayGKUzKZQrKavB/e3zLSQLNoaWc/mCL/rXScfMLXWnhJCS2n+rCUEoFdaHaPjhImcBAsvVrV
65wc/X/VpP/vmd7jv7Tf/vz5pUQ+Ce0q4D2jHILWGCi1lvqO0/xzwuepuhiqL+VL9j/ZALHJ2avH
RExVf/RV39JFy1qmI6RtLhD3B65SgqGLaXJosxx72bVO5h4+h2IhLad0b/VM6LvXpPrJqMaEY5I6
3zCfhOtFyciROEAE7SezeC1mLJtBuWg1Kg8NRQU4zdIokeyOoGKhRscZ/iAaTVEkZtxEUJ84QhYg
BSEB4+HF+jwWsemA6EZDPS5C5DbEQPe8/I00JzL1BjJI0tk+qXlkVZKp9wdrEb6SP/ERo/bg+JZd
NCWTTLslTYqUkyR5NRin1PbnQZA/gFOs9LddIbUkJlOkNEGj+u96Y5md4gPcLjaLviyySUmTO99u
eXFbxjSIsmVk3eyi2FBRKjjal9Ro+frsYVs4gd68no7jptsj1sbE/zdKBHR9bsXK834C6M2/onYC
zGWG9z0Mdx20CEhtThwfZSnU7sVahKLFvZ3RvZ+hXkRVDKyr9iFDwLU/e+ALCyZf85XcHeHCWyhh
+gUUYKmmRvONX0Ry8oBAXTlX5Kbjzanpf8DP8WYGs0qzDOsuM0wEnHuITJfSVKE5L72mHFiIUyCT
Reaiq0kAJoY/QjRxDVolcUd+K/ADUx6+gc3AsTp6loLmdgnhDwvcnQr26erpzEnCRONKnqNb7Qz7
9BjTSM1lJXr4efklelcnQKEr0xAOLe7pIi77H7qNod6pMzdlaolPK7hYamzqmKzhwt2nJPxyTGa3
dyCVuiKiZzB+xd3zDV/Q8SJpdE+vccluA3GbnXya3hZq2WmyVnx4qIHq4+1a9wnhJNVg7ya7p6Im
tzwQDdLoQap0FGDNbFrQLxY80CN+AAbN9SyvCgEOADtg7+/BTUsyyhq+u+yU8tvrclg91TkuEOM3
4QfdcxUloDij3eJZFJvBvIEybcjXs4zAKnduU+w0Kq32Ij+Ii+V/LQmIvWBp2vRmh+1sJlZlUVyZ
KM1PZ96chQiP2NQlOOkQNt9wLeDoaQRPedTZMhcx97Fe5pQAwXXKfEvrRMr5gFLc2C0AzOivDH8B
v4CgYs17xyVjx0dayhiTg9vufNnCNJ7bTAQxboXq4EJ/6NuE6uZ1PQSzl8NRfR7OIyIPR8JuO4dd
h/gbamqnQqLTvBnckidBVWDSOOufAYBGG8F1j6A8Iy2HwqEjir+NB3WUV8M7PM6qjQ6mGDwsz+mo
b3qHAH3tS0VbPEpwVfCJ8mWItkqhdxWcA93vD11XzNq5T3vyU/SzM0gLcoiV33MK5TFsMvXGuN05
rJ5Lh5KlPQrBaqHcER9RBNlmcGN+FKRHnQD32qd/mv5vt0IMWJvLgUjkW8ROCClueIDxCqXzufjn
IszrsaGSq66kpOq2/uu8DJYb91tP9sadxe/4t0IDcrjwPS6PrUNUrmE2uSJYvCWgeVeVISMUqV3q
FUjyjJ3TjeNX9SiV3JaIlqS/3u3PYMgiiI1pPnLLRx3Q/I0s8rxdJbZCjSHOBW4f6psZzS0KpEKh
OedX51N9LwlTIA8GLjAjmfSAVnmu2CTQy0tfukgfwM3vMvUGP90htx7lY5+U2hhsPQCftkdhiyVg
9JORdzhlq2powYWTs8gAzNC2yz/duQ4Lg8qTaL45Ex8POJxPXtM52cWHLBTYOihOFW7jRhSb5tUV
2z12VWa7gpu0uPEMnmfPJ+t72o0/PYCjfCsMWX+xP3jqqglKwwTbReL0KSB+adfxoYhDJ6IETUGA
pF9nC9azFz+Jsyh8foniG9ZbqkmeWENnb4GacW1NFZ6GB6M+HQh1+ZywRkd+dJ8yahB1+73nhf9H
ik+GtnZpb1gjHEt5W603dM6n8ZkrF1ELu4JoJ1xbaTfIm2A1/OjDVWlUNFkkh3oH00myTEpZKQx7
XDsLvUfiNtKwk2xJuhMPViacsC5MPhR0W8DS8cmz7TUAv4iIpX2S7FfmQtyG00sd2v5RauogbD/x
FHeCmsDxlzPM4ro4c1u26+FBJGFhFDIKaiWog729o2BPZ9sJcWhigHuLmO5FQ2U4YRebqWaaCTQ8
WivRlLXDaUt2p2EFefQY1hUpZacznliY5NAdBw+W/8l4uYfNSkpTFd17mJC5jaEN6Ip9kVz2I+/C
QI9qVHDRyhAMblFIxCC1/nyqS+Ie9zR5GoJWkwb0HCb5KsG9tfnTWqsfwhwnfh99ROBP5zNaRtVo
JiXAWdvofTvc1wD7YYUQD5K/BtlyQfxeilzpgDP6YNh/XuKysxbQvPo4ygnI3kc7BiDErykJa40p
4oLUuR+ohpRuyS0DaxLXcFdu9p89dk3MyEQNGIrRkLJuObxEtKN+Pwld+rLadILpsl0pwpMNwjNA
gFHUN//XZH0dB7RevguiSEPGLKWdOG7dG5id3PG9tQyacsweGVL9vJ2cdnevaq19cSsDGl4cXHsy
0Kc/TBdVLGriUh5LQ+i7vhQvY3Nej6xXR612tiZM5bVZdGTkEjgEsXlin427ywPFhugNvqFatSiE
j/JLYC4CdjARE/C404A6wtgJtGQ7k1S4LexQHSiqDsVBZ8bW/j3XOvEeT3R6KXOTWDKGasErAm9N
BC5MnViEtQ7VPX/ebM9B0kRpqs0jbyYZG/cYcM0ixhqe/NmE9c12WIiYSqOvV7Iej5bVCftTyC+d
B55oRbLhPwQ7idjfkMd90ecpjn94B69HGcj5AjzZ8nzOADvMV0dVPwhDD0LkCIXMCRPxQ46aePmb
4lkEy0MsNjHUNChs7V83q9UuzLAGLs0rIr6TdaVZDe0oxVCC2edsotpA6uDgcXBCflKoL8pLi8Ra
9ol8eMSysRS9YJ3DHiP67R9SZ/feq1fjZWPqg7o7wjy/qmTjgGBU3twmbIcOQAmNg2x8Ei9s8c46
jsUd54NhSjiFhLrzlPiN+IxQ3DRkbv90GxwNWvE3px6XyxzunKqV1b+aivTuTJ+QpQOKpfpGog7W
U22CGSKMjbQt4HyClPfYwszljuB7LcVHpfReA0bO5MGMqcHWavuoRx0EgKYDPHCTiRnDT3dzL0nk
n4opCsnsySpUDTStJ0otCA78sjlBv3YsUdcWM+/ou7NzLjArBgdENCBIsPsGAn1AycIjoMDfLNVg
2S+AfJ/a2GvTotmkqQkMqDttqEH0BlnpWqzvAo1dFlJKVP6rEZga5UPyNOhZcoevvddBm3ocsI4K
zMd41zEtSSix0O6Pflm/W66ou6SnAGte7CDaT/l8GF0o3YkqdCJnKLP+HAlC90qaz0t/s3CUoAJE
B6J6olm94zOfEVcLxWiCK9BQ+xGpewS2XkIJd910o8EcpG5iTKpLpdq9FSD3YCzfNru/y0Qlg+dW
bKWAXXZROc3yYDhSvIwO93bynV8OyyaaLpAAydOtcYtEbZOwoAIA/DRkhdCTiFYBDmR+fD7CK064
e4wwog3MldKgwwQ4XPVVxcbHkHxfhdoZtFtTsFqNInr8h0htt0Am1ugkIaQNZvYdxrTryMk4ww9J
VtmqPLf8C/0jiR6v5ccPnxornNFj6DR5/Azble6FxwnKKPGvzf3ZMTipsh4qNGaBSaOGmEDPyzwA
UFUz/3jsxjQp2XvBEPmf1rbh30l8B9VnGVxkwlJ2ZN+oImFy3A2zI93wbjQCQw+VubalM5vidnwB
1j/5gMKDfF6m6eLlalOJYKwROnOoJlUyW2iMbzU9wA8N94e7f2ngKs2sxMUHWy5Bd/WO4M31H+CQ
MSjngminXooTQ8MxpRHA+KQ4GuxKF2c7hlui6GEe02K1u5Edn5FobqYwdOVRCtSH0aXRWQCWfpET
85lFmBJfoQg3pmLjVQZUwiAz8A0DBsXcpGnv/IhsZZOtQQwetHiIVAFtYV+Z/eq+ldG0SmLHYLn/
ZoevnJzpbqwhMHe20DcFwbXuNfW5a/R8MaaPMXLBR4U4dJsVdMh68ors3tUVzeS3+gZvCMfV7r3+
lsSC4TM4ziDUNfaIYQSoNCwFa347YaLq4+GizSkF03SP44pX//JEG5O+FsN6HtydoSJrnJ4Eqi8S
qSfjPX3bj1GGS064y7VcdidfKhqzWwTdBEp2UmB0aLwu42V4XcbTGEZh7TmVXfSDKsgZ8x1D7709
QAha3ryKqB98Bxovxcd4BceBL29+nts8ihrn5icYyQkg8bM0G/Ud4Bq1UyNUTN+YOgSwsTuaTTRB
Od/CeXjwtOUBFAPGqJW4/hVSjue1gGjwkGS7UOcxVR5EA0Z1iBso23vPm967n3aqa/YSwiIHdnyF
JHwAc0KUcCS7ss+gLW+yNZnoQ6kZy43PWHfB5ekHOM9zQ8as+wzqyOL2eYLz3/y+yX8mp8aKhkDy
KAmONqtI0JBzxU47Lod3aMB1fuLWxSTmhMs2nKyrG4Wwt+te+t01PM/T72ay64IhvBWSdrUiqnoB
pxTl81agxWpsLYafLN7bXWWuuZ3ZwM2xysywUfqevN2bKxskO764ZLkhFnKltiKvTt27QhgSsTYu
+1KIM7Y0sw5F1VQc0TE5s64Ikz8olgIAbu5cfA/pjBTtHmpNHFjsmkqJi8BfaDvqCs99AWoDImk4
SeFrdE4h2wTN2nozMVIo8UcxkA0FqQCXMoLFU6iASXWVjwJGvNVSnurGvXnI2Y0egT8su826TgH9
hHp2A2iPEjV9GlVyV53UFPg28tLaGQYpiRrgPB5XXCXN/xPCrI9VD6UtgyeskWBEnjMtpndWAkBC
Tyg9fAiHdsLAm979T8tA2z3rO0YkeOMurrocuv4nLA7PoI40cGTQ5u0JKpc6W9Kj+8dOF5XeTGk2
EfP0fr7kF5Q32kK0eope0f5rVIrcwBpI6SlADdd+SFpoLnG4Uop9sMZcAiZgTOXsNnUvpndAHLAs
0qAI+jtW7/KeW5x6R7+QAeA7yPBAiGTIxCpPOwql2fZpqAqSzTB+TrmV1M3q2/SHB45geYyDZHjB
PhBbzVHgFDj0Mo2xPrXK64cbyMlLRjGNgzBqgixFqajLC9hK9rKzcmtdD4dcnStNoDUTy48yCCyr
zRbohLzGZLKrMx1AB3fhN1qK1jWw5sZf5vsBMdjO4UAgQzU6Mw3M7eQFwdLEfuqKW0cTjc69hzbO
mk86QYA5OyZjwOZeD2VSgvThaF+OJuMOz8bWrd3v0Yk+XlCCWhmhKDMbaV4hw/TVKDihwj+oknYL
uSPG/BPkpgBs+l5whrJKpIOPTVlkylxTua7IHEJyNqrHSbRR8y6/No+LXD2s23FbgaWUVVsqiS9b
RCJvI+4l+z5CdWzS7ZAzxFLpJ3LCCsCs8X9uRsmXlDRBGKRlQXFvv2xOHwRwykBb152z1EVPwiQQ
be7fVg4KBBGWz3mHNzogRc1gKzC/DlKkXAinkCNeujvRQBvbTbTVi0HeWRHIJy6zWXAkdiNKpjik
cMKSLTW+t4FCgFZLOv7PQSS2jmkGlgr3OdzzO1s6G1tDIxmcR97rsPaGjCHZ8DiNz/xYdaFy2/Fw
Qtj3QTGLIydAuYRoiA1tbe63eAPBlNrteazCFym34LoXTRoLEQBMJ5qIFutZYMqCLIXDW9oMjaXj
kzYyolwJF6T1pK80OoGlEECKXsjKg8lEFWxz6kRVSIfMQeI99ar938tT22+8ogU9ctfSnSg1GcHw
LPVntd90UyLmPwVv/gFZsFfVmSBXt10FcWK5W++a6kS6XScyvbuZrbSspOU8uqU7+ODQ9MuzJ6ey
xEBwJYHSLTHb/xyQe/GN4DIipFxnvv9kv1irZDLn3KxrfTW7Keeh4h97dbZcncLnSG3XGYDH3y1j
aa5N4rtF2KhwpbO9grH9wFY7CuMrG/8zqKPWwlHRtyWeozUjp4LERDa5XsUIzmoXZWVcPOjDdlgG
xupsaeOqvOu730KhkN2MuCwapGg0I4IUpZhUcZcYwxT0NRtfz5NxVqSFWBDpV0X8WfjeVWndTEQ2
bbR1aNyk4nHIXcv+beX/6Q3V4uIhMhXSCEOSo/fOavdmhUk1cLPHNOJ2HxmMUCAijZuuRDq262gF
jZxcKgUwszWc1+doklMybjZL6QZ4ZcE1iN8fQSyUCW4MKlt5VJtSy4Xt4/rBnbj7bZhuvTf0VsY9
qBoTRxJHrKzrOXKk41BB7PRJcaX0yx/HxMMDH5eXw3YCHrSMfKi4zPmSmvriv5byulMUgeb+KNYs
V+j7+iaJuucp0f6BdNeKTjxMGbsak+igkd6v2qe95Lb/nWZ8fVTNy3OxjbkJbCT8HEAkiQKfSLiv
ptxuzmSi7O4Y4dfPJQhXkNec8SBhMxAE738j87z0PFiMxwyQuhHmdpcQqlVha7ElN31PXQeMvlyX
6X2wAbyT13LLDJoAzpFhigUekDz0BXNd8/gdfTDUTMPGJzbwuSkoyZXsXfjHJSgennq7oHAZeqhE
pcqNxEFVpLbbKeKw9XCnqSHzuXPcxtwwGyd0AlgQIyQ5WmoEgs5HhiYkQ169m/fvCbuttXzktUbk
w1akRODy8U/7zuLv7aESkop6OL25TWLd4Klut+oT60B2Ti2FkExrRbs4RPE4f80u9b4RYblDtQp1
kmeqYCcPBWJd0lkM/lnUtFCn/JN0lv+mKQaahRbCkYvJI9Qq2xFznGTvbba2YWsrVv17U1q81b89
u4nrAufj+lPfNWLFS0BmWqKnR7rXBEWEAX+kgzKlIXjLhi9GnoRq7U4n/vqQ2Xh5wSa+tyD7OLZG
qFxGzRXP0diYOm2UkcZAD38lXi3hrWQPmW0X0QUAVAtLVTDj2yB/1Dm/+CTbEJYdLcIcDvHmluzt
f8+067CdsDfPxp9PyIQql9sIpzbdLeBoAxiZkFrUjcKUPYJFUYfjRcLYNWuIKb6093duUnekcbB+
tlpc6JPSPukWIFkobvZzTaqHZXbTfV75oBznM0h9sUThPJif402OCJrgRamhfeHXO+zqjXecEFV6
uPLy3XpXiLUQ5aGWqOTnexkTRcNyz3KsYTEVSDH96S2srymKYFyxFt4XOu2KKjMURYA4O/+la1N4
P/fw3prf9zAJUCn3eOTc31vT3m0FgIcEmQlpEX8vupFChILCUmxsN6geqv4LYBjku0RJo9HDcowA
sRmPeBju+M1i8aaaIvQ7utCYJ3AohoLtlTWw+vqE9DdICw9B7X8azvme29LAVV+TXoB4k62TOvB9
kVNc1vJIjyv8glMUu7quXnNsaJfvTZOyEuAqtSKixdVsGl1iKAYhBLDxDPI29Xq5+PsKV8duDebx
qQ+mIslIYVWBdoSim+R1cUB1FApbotRepYGtoui2AOZkDnGQTg7rPWPdrqJFuQFVCST1jYTwFl66
W7dJ6LKNHlmHqyOLx1p0X8NH1BmWRxpYeVBiM7nM+ceeCzNszWupP+Ck5FObM24y/BMMD1DEF+rk
76g/THvLaWSe3aHkSRDD71VI02+oU+cFcY4LwOgBa7QUyFDlaOF/6MREcrlJnTnCVG9REn/GPST4
hmqwTqM4yQiWCViyAHHeyp0SakaN/aWMUd9Loi7u0z09xjbvZAJiTFVQNEWtXSywBq5Je7OdMFvC
rMEup9tkEUCSPDEfjBwooSlCitFQyQdGfXxbQqBIDshe0Ualu/SHMc8II/oQFMy1pGekCRtakC2S
ZNu60qy5ANwM0+jXv8N47GaH+0caM0SzwIiq2VjYKRfoQHsIXbSvQcWgV3FBSNs=
`protect end_protected
