XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����{�Qk�T��Vkk��5Ǩ2�ǛGGa�q}���Lf�f�J�(��';���p� �����9�����V��]g:�L,E�鄽��h����v��}#�Iy�:ؑ<:d�%<���3'��7��� �T��@���OY�Ky���uo��R/
9/z_E5�7����ϙ:X���d/X��e)E���#��mS�!k��׃�Qj>�s�N{��tU
_g�FJ9��P	���%��W�T���ak�u��+N�x���QT��l�H��Y���YUҵd�hb(��Ƨ��#����0�,ţ����YքoO������
�3|�A� �b,��$�1��9)�pA�ZLS�=���+�j��x6��[E�h�\��N>#ο^4l��kM-!i��~��#|fd|�RZ��s��P*,6V_��#���=S��sJ�6䆘d�t�ӥF��e�9�R��|��������kD7�ȋ7Hg�r��s�BΗ6Z�}2
�TW�y;Xm����nf�&+�&C�;��0���erm�O�G��4�G(	q�)�w�E�_s-��ǅ,����<yDA��$�.�7@�F5�?9���ԤĿ=t`��d#H�2?�b��ǭ����$qC�\_k���ed����~���N�Q)� �"����k��ߟ�_����M�uR+X.c��Hf]m�4����ϖ»u7�t8CB�E>t���0n?�[@F��|�P��V�޿�&�-��f����w�]/m
�B��*��7�h
��y��LXlxVHYEB     400     1c0�b=t=Hr��mv#Z�C��#y�B���s�SOӘ�7��8T��x��G�M�$H�,�p#�PYc����a��_��Vy4��5>s|�ړ}�?F3V�s�*��ߡE���̨��y/��ݥ_��W=��֌�t�.��O�P%��|�M�����(c��׳5�S>��2��W����{ؖ�����#o2&�N�L��Q�bE��3�z��X}��8;"���U�a
�Ǌ�f1D�'�&O�nPJ�=���bV��S��G��JT������Y%z +���_F��iA�������
�����U��Zʳ��\!�^�X*|A�㧹�D�π�Mm���M�0zb�b/2T^5�_��y7
�<�|��(Ϛ�[}�,e�I��V����j`(�����ŃT�Fxᣴ5u���cF8��y3����ھO�d@(�&��8��NXlxVHYEB     400     150��Qsw��M�%���K�,q�m>EB��n#���uБ�Kj��OOzh7޳��AM�x1���40c�Ly� �������i4��}�޶���֌���l1��(2�
����à�w`�B�
#�g�M��p�(�ں�a
�'b`9>* 0�q��y��8g�����A�b�9y�gN��!a�QC\��D��\'��VV�5)�B�q0M���R�������'�ʑ�:N8��sSQ���y�mI�~��.�kȓ\��������{���zH��;Pi�V� n�o�`㰯��)$�4Y�apN�
ɒ���(����)��XlxVHYEB     400     130�&���w�L���8�����Q��4�BD��x���V4�XΐnMi��G-|"Ff���8Y3{��L%����`C-}$��-��:�W�&�PT`x��_���(��B���_'#E|���P#\�dn�H'��y��sE��#%R��F$�P�e񏣅��i-�����d�j���wfg����u��
|hTd�U�t�E.�tG!�(���ԵH�e4�y8��vߞ��;�9�#�?��m?e�̵WLǓ;W�bǏUG�R)&�C�U�d�M��}�XC��M/��@ʼ��]�?�T4�筋fT13Q�XlxVHYEB     400     160���Z�^{�7(�P�����'0O�m�,�{�#bz�ہ̷�� �X�Bv�j� ��n�;��$�C(���C��K���eLgEI0{��7Oo��M��0��kr�q����yF(����"��}�{pY�^\3�+|����0n�,�el�A<�A�RAr3`�%A>H ���	O�K�q+��?��eg��;_}�ov�f����)LН�ѝr����D��sp�T5ׅ����a���A.bd���z�8�M����c������'�<��Š��#��w~�J+��d�)�`���R���/�V4��Fpp{C{�,=�\X���b����f��ڻ��%�@�*i>�Γ�v�XlxVHYEB     400     1e0��f_ñiJB�P�hdwYդ��H��^y�D�G�����kB�v��㜨����Xpb�*�Ӳr��:����v�����"*Z�G��(��Fb�h��0��3�K9b �1��?iҏMS�)�r�K��py���?*ߢ����;.*w��x�E��\�G!�i!	|��p�$�ģ��״�e@�ދ�oj'���~'rW�
[Ç�e&C�Z���v1oq�]�ч�A�3��3�p{J�ϵڦ9GL�7V5 �&���6i��Wl/K���w�p�0�����Ϩ�BPz_�.�q�(g;)_�P� _Ԥaϸk�x#��P_��<R��l���=lEF�NJzG��AN��>]��@��TCvÂ�{O��n+�F�@��Z7��Mo�(̥;H9�u�Tvr�t�է����˦	MD�	�@�T\���~s1���;�0v'XQb��_愳���6�'��B��*H�XlxVHYEB     400      f0�u��Ezd���VVu����YPc�J���D[E�yW�b=~_dݣ ��l��#��Zŉ���b�{���1b��Q�0ɞ���@]�sx<���v�=�{ʰ�A��͎箞�"��7؃�j�f�l�f+�����F����	�JYh=�%t���٧Ҿi����xr�q�\�l 
��m���O:��v��R���9�ƨj7����LI��Vu�^xT�8�a�����t�� XlxVHYEB     400     150O��:�o.��e����h��"x�3�#����V���1ѯ#7����z�A�v�������A�:������s%�4K���9��z��VE�
����Y���u@��|�s��A6�WKV�P!��ώ��������?���tt�����;�lA���mMH!�R�Ǫ�#s�wL����$��f�ޖ�������Q�ʘ�Li?��YIw`��������f�hk{m^E g���L�ʧ�"6�qrC���; -��g�
Ҝ���ШPdGpݞvpܬ{��Ԗ~��/�Ϣ���v1|�K�/G\��&�B�XlxVHYEB     400     170V��f�I��'O<9�h$�
`́�}p�>��M�	�Z�i|��X�FUV���#���4+��'��iwRؗ��b`nr1:������9��!���)<���a��_��$U���T������s�Hp�����q�u~��G��;LS����rA���t{=T� O��, �J��4�i���!��7s$��^N"Q�md�%\Ķ�&1D�}�~��{F��Y�~&�e�\��St��A!���5�vJ��U`�З��Ɉd��0v5.^ֆע�����U������_�p�f������kRY�k���ӭ�MO���e��h��=~)5����]< ����@��T}9��z�η ��B�<���l��Tq"'��XlxVHYEB     400     160�Oi��K[a�Dydz{ߩ�&�6��c�c�u�M@7�Xg�3�2����a\��j]	�??�~��n�ї]�X!��x=����`�iE�>�d"X��B���x�&9�lv�A� 4ţXӲ1�5O�dj���@耵l���I43->f�O*}��vѪLO�ɱ�*%N�=�SZCJ�Z+�mcF���-j"�%D�.�0'��\�8�!�x� ��3�*M�A�q��v�h�(�#m}%�{�6�h��e~̴>����8CY�")���-� F�%T�e�%k�<D��|`�G~X�v����6���PШOh�qBj	k� �~�N�9?�ʸ�����w��Jbq?�ٵmU�XlxVHYEB     400     180���&MG���֋���[޿.7�U�7x�H4�n�Ӈ��w���ę��
���))ѻ-�2|b�l|=��ag��Q�L=CrKg9�D7�:y8B%��'ĭ92͋2�G��9B��z!?����"��L_��y���Pi��t�ۜ/H�-��2�E*d^�xv�p^RP<Ř7�L�vGȄ5��Ӧc_�N��������jʨw}|���ia�)�S��>A�p��a����y�Wa�~�Q�7}x}l�u�F��w��T�"U-�E-ySL�z�'ٵɞ��nz��]�w�fL�tJx:
n)d��)���{�'��/���N�����J����˳���%A�2G�(�[N�1��f��p(�6ITb�XlxVHYEB     369     180&�7S�i#8θ�V!_k��zGF���� �� u��Ɏ�>������H�z�8�Q�NggR�\XC�@,�K��,Q��6FdO	1�ץ�`�����{��&�����JKAg�>��pP��A�?>��s! PT�����fL^�i*'^�+��8�~mN�H�0ȵЀ|�~��%ZPζf7���Cc�C��o��M��a�r}fo�^B�8��@apɇ��m�A��+4B|.�&��Hd����f�f9��)V�Ѝ�1G�l���M��Y���a���R%����=��6�d�%�&k(��,4�����Fa����\ÂfP����4+K����]�llmj�%<T�اb���W��&�ym�%��3���5r��Ѣ