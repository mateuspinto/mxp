��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���)�{t6������i��u̒T>��")Q"&(�$���#?U�
��C���P�Z�̝����1�<;�"�c�׫GH�
���o�k�'��d|U����
��X�\�1�f��}��N��_Qg, ����L���!�_�1l�*��>Z�2��3Ru"��&�|�����Z�.MA	�	�>��,{��Ӱ�s�u��B�T|cOw�	ת�����~7�%oY>� ��Κj�Ku��+	jhu��ȵ7� ��	����g��9񲛎�l�Y����"9�4��M�-�����X�r��P �s�O��U��=���ar ��=�pJw�WE�Zc�`�DR�u�#��"HE����T׊Ki�G)x�����Φ�vЀ;��b�Rn�bKOX�p��EY��b�1�؋�ᨘ1�l��\��w�J7ī�%�m�=qA05DI��{]m�*r��#}T)s`t��wb,�2�a�8�>L=D�<8y���^�tsU\	m��7��1�A����4\l���@a�ܡ"��}�D�6�O`V��� ,�����$��!x\J}� =�;�<D���/K�]O.�~������-@T��V��P���Iu@t�ݾ����b+��%�'�OF��i���J{q���]�n�U�!�y��G|���{��C0�g��f�����Y &�h���PA���?�@�Q��:�v���[�;��C����7���Z��y�2�im�tO)d�O�����$ '(�w���&���Ȭ�AZ}������Mwr�;��ts������.�Xī��X�B�<ɯ�e���R�V���^�p8�圀��,�e�-m����3+yz�F�\U��S�G	Y�-��q�EH�,8Q����_�M_O�Ǥ	��5"A�f1{��P�Jb�&XW/t�f������M���9X-��g��s���*��F��_����IETS�}��Q�n+N�)�kA�{�����K�E(��7>;h�"5�:��|�^e�=wP�AI�����ؾ�ת���|@Jp	�_�j�DJ�D3���i?yRi��PFc*AД{� �tCx ͥA�)���:��\�|w��)>\�C��/�Lw}���u��V����˟��6!5M�(��'��ۢ#�l>Q��&5[n���B��w(N��*��z��{�-�s*J�őh�&����t�g_f�+k���Z��^ S�O�1oM2����X�����9��ɫ�1c�m���K���"۷*hv�{�տ�tT�Xcz>KB!���TG�au�������8Q��G�\�װ脴��R�@LG3_(�g:}\x�ڧ��x��r�Ε���ūe��`�e�Z�ȵB���!����������~�O//��vrWn���\�9r��6i���^q�����I��T�$[���8�"��8�Ba��p�M�3����wzM��z|8b�kG��h@1��n����"y���D��A�!��3�v��8Z�?seѣ�!���D2,sИ��At@͈�ݘ���S`��ڃEHl�����/��h��w����7����%��v���-���#�P�4��v�	��o �<���;�Dn���f�Hǡ���-l�1��9_��h�_HU�b�AFT�vm���_�q����MY�6a���,��	g�8"�E65ׅ��d8� E��oc�O!��iY�A���_"e��e=,�K>����Ml����a~{{�-��9���τ�Q�w�T����c���~wH�^k6���G�<A���6t�(/����r�L,�
�b%߲Uy�	!z�=IH}>�ި0%C��*6|ih���s�%�g�s��<��yS̙���يu�+6;{��i;r�� ��[nD��$ۋ5F����&�,�܈����[���;�G��,� dU�a��H5MnލN'�etry��+R��-�����D�=
ԑ8������hw�k:�J�DU�=����r�"  �4�b�'�8�l��e
y[t������l�R0<�"���9_#=�F�RoV�?�R�^�͢.%*Tv���f1FjK�M��ů:�V�|{�s�S�h6�[�~���R�<ާ��&�	�	U⫹3@��E�è��N�	ƾ���;NBA-$�5�)��e��y������S�!���B��ɷ�`��,��
���p��x��Z���G���Სm��=2k���F�B�H�t����_�Md-��X�	Aς$֪��p#�˱�P����m��ѺBPN����R���,6��e��b��g�`f<�TY7���M�{ ����I�y���J��ӣ�y�<�{i$=��J��j�>��j�Y� ���E� �+����i�;��3G��T�i����@93�?�v��C�n����f��)�^6����O5��6���oL(�oN'��� ���hek�u-8�Έ�cG	��$���9J����Zx�>��� .���W� &���/���¸�X%(#ümK�[C��8�A(���F�~�0y���l��P4���}�G�ڿ1�(E�낂� W���#�Yo��U�ysѻ�R��0�p.�+G�5�F.�I�Cb�.�5p3I��ߍ� K,�o~$��&.�����]u��s�Y�ɻP�>v5�)�u&�{z�]���gw��s�2L�{����C.N�}�v�-��7�N��!�C�&,���wդo;!xW$@�#��$���
 x���"��ݾ�<Kײ�E��3�0b3*ܡ������Md�L�w�7T�l�&*���&tLƭs�Kl�܍޾�>�;�� ���@͢d
��|Æl��۹sɨ�Y�D�N��O���c/#�u��%$R�R��B�u�<oMm3���g���'o��>�Na�i��`�i;�֥��9%�޺��Y�^V�P`�����b#��;�0�H�����;X��$O��*B�FS`��ig�j:AA��GCz��<軽N�#+�ߵ���4\<8-p�%� ��A��-�!���w�!��F.-"H>vS2i�6_E���q��Cq����֐���Q�D�n��)5pgV �P$I)�*Ԙ�8ލ�Y��d�߸�@�p]��(��2m-�/BK�c�8>�/�1��\� �X�
(�e�r��0��t�������`r�]$�bjbXV�W�ӄl��Ȉ2B��܂i���:a�2:����K����Dy����~������xT�A���>H�Q�d�/��N)fy�$}������:�<V7�E-��� �*�Iw����\�Z���RE������=_N�2�X���Why��]�\�I��	�����{�v�'@�H���7��HIۭ�f�*��F�?�r��e��o�^�c��.����4,H]�8S��M�\������E��n�VP{�nD�}����(���G@�?C�\��^�9��O�e���z�X�:��^�6kZ�3~,=��C�_,D��ޘ_4B�b���U�f�а�uV�e�
��r�Ȕ�_���'�˞~%��Q i�����pnP����f�Բf�\F�_X)�(���7�='�T˵���1:V�j4�_Ī�Q'�ŷ*�(���7_a|�HB�r���*Z)^l��ǀ����Q�T1#�4��Ci4������K@��`H:����R�' cB�M����)���R��C�Lc��N��Y����ph�Pq_�B@����D:�����^��Qy\�#㬿C�Y�;)�@�%�V�:�������`�~�Ù-Ȯc���W�J+�y��$�F�k����H7[a���x�>��[t��5�Ju �1�=BF9�� DsKt�gk�Lil:���v�X�ø��.�\@��c�-�&ʅ�4�Sa5�"XtK�ۤP��6��d�Xf@�0�닯:B`:�*0)�r�P-�4!�n3�n+u����%E��߁B5��:��-N�\0ۼ����K�����ȼ΂o�$�12��Y�^f�����������ڽ�ٓ_�/��׽�����zo�F�Rt���H9�/Y�GĄ]��|$��"�Jݳe��TrCF
Ա����*��A��+�|�<�Y������3��qÛ��P.�s~sD%�bێ���B]6� �zl��(�L���}4�E�҅���O��'��Jī��,�r���?�G�.��ڧ�b>����T��k^�
	V��Yz�#^`*�F6w�8�mUHO���sm��3��8}!��q���isg�Q x����Z���F<#ֳ,/,k�7r Ͼ��I�-�Eay���f�X9��g.�5Yj<�I���ܼ�	��?7e�����J?ui#��̖d�lN!��"���mR]g�20;���
c�0��|�ۑ����|H%��9\7[ɼ���$f�ت �>��vNG���<�L�l/jc�(�����}�3���m�a�6�0D�Q�.cd�_`��z֞n��*��"��?OB�u]�`]�Ds�~F��)*�;�Ms����m���Mx H��d�S_~������@K6}Z&6�Nލ~�L�mԎ�v�e�͸A�摹��>�
m(טs��v���1�X|v5j�᠐ii��G7ji�A��4�\�q,@��8�ѱq��E���ϑ#4(��� }9d�ԧSO^/�A��E�����ڞ�	��WӦ�����c���m@�:��T7܇z&�M�:��v�}��M5r���/Q�vX�L(�;����(Ⴤ��|ԝ��K�c�����q���RL�7��5��`3����mt��^�!˺�$+��`e@ѝp��K]��J�T��a�ʥ��ˢ��%b�_?�UN�d���<b�.G������k�y\��PW0%Ud)�|�=j\��]kE��(�7��;��,�Ծ�/�db�7��o8�.�//�����J ��Vh�d��;�T��T�C�����^-�1�Er���;���+��_"�>1�L�%&�/�ﹺ����?��m7�rM/� ֒�领�� s��~wث!eYE�n%��?�o���ЪH��5�|���+�5�8%�� ����ꕱqL�
���}J;�+�m���$hvYL��\�פ]��+�H@	:�C
�c��8=�ߪA��'��Ń�^S�l>�P�hP�d�m�F9� ��޷�5�K� �M�2�ȱ�V��Z۞Z�I���k�������X��'먪J���mv������9 ,�u���o2vo������
I��l��!�}�{���nׯ�.>
�L�œ\�x��`g��!iy��h�! �~�_�beeڮ�7-?�&���"b/X�kӻ^s�=Mٟ�(��ܛ�_Z�����"�p�y�ң�O��7{5>j�VX ��oo��
g㟫+��L�Sn��=����q�6}��c;���E_i���[��r��� m�Ӑv.S�P&���8��j����H�;�5ʇ�X�T����\$}F�>W��� 6yw��	���%�u�9K�Y�85���J���0b熁��&^`�Ķ,�(�&�^ӭl(&��>oj�b�۳KO�<?�����A.�,orK��`a�p�;����&x�<���3��g�v"�y�6�&J�(Nu�A��D���w=v�VJ~����ȟx��������W�"/]e��=�u�8��!�,�LV�S=e~'-����:j3�/_B,�[G�]�ʱ/��D�p��s*C� yyV*ڀ�Y8 ��`_�D���.f�;�C�I[�}a���ğ-nʶ̢;q-��u̼�OGn��Ed�,J�����~$�;�Ǒ^
����\Z������/��7�5���2Y����o0�x�v�JqS����~�I��6s�?�Q�0�|L��'=?����H�܁��vuz��I��:3[�N��s�"J<�j[U��?�����'�����H�K �BC�-���j�����{������=�@����+�
v	N�� �y���a}��g��>H��g���U��ċ�<�2�{O���Y3!|Z��X��c�:v�~�F���7�9���x�R�eg?K�=L���W�l��Q/�_�W���<G�J�r�4�<�z�����X�k���4?aP\7C��Ej���Hd��F�,�G:dFJT#�MM�:��߾����#�à,���҉���~�x2w2,����!�:��[�Q��M��>�d�%%O[�����~s���K?'r���2b�t��)q0&���d�@�s0s?���&(J����XrV�M�N�L��֛�h�fY�D�H��\w�mY[���۲��[��5G��҃P�L�i���_%�Ec׍�u�o�£vM/���m8�{�z���M�P&P���KoYi7����8Zs�B8b���	)�1���M��ģ�I1�M����Mb�I�c4������au�j��p]N>H>8[�}��;v������Ӏ���(�ŝ�L�M}� �H�AQ�c���ϥ��.��/p�����������*"�����Rf5��qB�Ԡ���3ha :P�unq�W~�k�<�p��=����s�jw�Q�@V��t���#��V�?�p���W+�#U\=���Ƃ���� ٢O�Mջ��W1LE�ډD	X��Z������b-�����~���!B�6;$=3h2��
N=u�o*\1��gKW������Y��u���Y���5�^�V�h�՟��i�t\0J��Խ����ۍW���R�d?m���[硋��]K!���s�=(i� �3��4���,> ��D_�s���wB���gd�,b��'�
d6w?����Q�bX�L����� D�Ur6lԖC�dG�D ��W���9OBu��6�$JzǞ�s�3�� W��x�%^����&�Ai���CD�)��
O��X��<�Xrt�FkY�c�1d9:ހY�%�|�������ڻK�K3  �W��>�@J1ˋZ���X[Fk���x���+ᡜ�X��s�U����(A���1��lœ�l���e&�]�"�Jk��
�o� ֊ϫ��b��D��V׾��Ҽ�*�R�K��rr��C���{<ҊbA�.���q"���~';ޖa�ߤ!�b9��D�͋�'�Ug�\O��AI��l�}Sa��1T�����r��rҞ�~�o#]+;��]�JL|��껮<ql�o�A3Ym��t�����Hc�j�ì�1�:�����c�O�m��2Uʕl߻��H1�i¼�z�$�q�C�v�{3��aѯ#��EE�Gi �p:�+Nr�����h�)��ɵC8U�c�E7�?k�l ��1�'}��5��(/2[t��4�q���5aD;�d�X��E��h��VɕCH]���-w���ª�Ra�Z$�¬d�C� �c1a�s���q�]�
��0iu��\�+eZ�*ʚ�/?R�AI�g��Ғ=��M�<Z�&��	0-���I렉�>b/6`�?R e��ݦh@e$X��x/��?j�7a�,@ q��۹��#��E;�6�m�BZBN�āa G�]�g8J��[r�!��!`�Y�br��);���M�i`cp�K����10&|Ɯd�سHH�y��zŪ���s����c�W�OU�].�Fm���gk��ƴ��@�=0����]-�ot��������ɪ��f���V z��3���K��2 �:=`��Q(���F�&���?8e�y�u�B��;�l^1�%�.�$nM������pM7jz���n�$����C&l��wg�d�� s�U�*�3vF{��6m�b��� ��G��([DW�h�~�i��T���5�E8�����Y�KE��A�ݯ%�"���/��bǝ@��
7���[���v]]�B䦌i�y��^
�:[��LtP��K8~��׬ٗ��М3�C݂-CY�5�!L��H>+�Xzk�a��T-{֗0�����M���|�8E�p6���e�{Mn.�9
�U)������`h(���$B�N��8Q�O&�ln����Z9p�yQa�$��Q
ԃ,�6ط\Mk��԰As��ϚFRǉ�V	�����1�ԟ�wqp3���1}2s6����	��` X��\�����y?Z��8�+��Sm�R�,� <�h��o��w��\�Z��DQ�2^�ݚ���j���8���	H7�7LI�:n��g�jDU�dF�,%�+yp۰ȕ�D_]1��cf�i�US�)�./��;N,czX���8�_�Y��"��3��E�+힓��+rsh�Ä�.|�:3�0�bN}�Ӓ�`���$�kɄ������O�)j�U�|��K��TJė���Ƚ��U����.*}�gA���0�}�lNb�	��2�¬�(���لC�(\�6&�;���4Bu��8:tV���+��f%�	%z���n�=�7��p��2"�m����t�ٿ.��(�A�b4��1�#�0g�� 톚��J�Ԣ��AOL�t��w��Z<��i���O��N��>�S��������C�F���F؄�T�8��䝎�f�Q�t�rƽD����m��J?Ka�ힸ��1I6��:�P�W��"!��CD����S~��b|�cKEr@�%XeK��"��l��*�E��N�	�ث�mM�x�m˅go�L�.A�o�n2Ը[b��K��F����q�O�τl�/'�"WǤ��P��q��mnP��2V2@�Xk�/1��ʫk) �߹��&�m����ڡ��i��yU'�7��TI�?4��y?jzʋ��O^b��4���Գ�sV�u�?��F~��IŘ�68[���ޠq��̓#����[9�j�Vgo~�SԠ���C��e��d֫큖���)�Qb�C%-�����)Q���v	���Y�9��Z�mxw���^�0�p���e�p�4,��_3Eri�By�#��"_�j��3�ʎ+�w���1�<jI��I��O������R�8K��::�JN�V�AѴiZ֐ד��x.�U���U���� ���<Z(/�{���$q.Ѻ�Z�!�~h���0<��� � �����+��B���9M�T�ʮ��."��4Q���A
a�� �z��
R)]�����W��������
`�����[�bp]��C#��&a�vct�U��0# �E8��|c$r��H��M��Z�۴k��5˓I͈�I�9��-�� ����DvV����!x��5g=��.GZ�҇(f���3�����qE�*J|h�"���y7W2�{���҆�*���f�{�
�`���uA@�920���u-��r�F+�`����wgJ�o����"fW���$�8�	��g�K�̪�
}��%Iմ���ׅ�֣tY����,[��o�yʒ��6���@?"A�Cu�6���qo.���K� N�����J�Z����C��QBNzFA)��m��ƑZ'g����f��Q�x��M��yh���(��S�CZz`�g��+k.�.�����.M%�N��m���]`O�>Ӱ\:�Z�+9��9!�� �"��`A�y��ń�<~"����n�.�)YA��yiY�t� �360D�[�M�#X��[��ř�86�'-���VHfM+�75�ͯ�����W���>��_�=�W
K�j,1L{67�j�?݃V�l}��.Ѿ���s��pp?Ө�+��G��:�Qe����Ze�4_���>QX�M���M���v����G�<���bk4I8�v�dû�X��=��[c��{
S-D,e�e`�}2k8c\��q:>c����Q�މk�[�s��8\D�R,��v�#�_8U��<�O�E,�����%�����n2yxv��VG�&�|9l8&��¿�& ��u��!��|z��>>'�WF����І������+�`6��V;_�J��M",f:�B�!_�J��s:�B�&�
s�.�.�>
���=����±/з͖�d��n�L֍\��)��䒭%��"��di丹��o��J�J�u����,���z���tW�z�E�?R��Gl��nv�+�I��A-PU�Zm��8�F.=��Q�1b�]�Y�QAi���$X+����)��I^����y}l�6�dj��6�8���I�����ѭ�V̗�F���=h�j��r��H6i�#,�m����G�c�>�MDA�5Gi��9���wC'a�%-��m\��Z���� [8�F䷝�!l��}]D�@0A���S�7��E����̒t¦'6��q���ü���`��J����h(����ĝd5(�����<�������.6�����݈1�H�j��{`=�����R8�H{vw���]��=�]=^��l���r0�O�9k��WR�f�G�XX�u�=,�����Q:p�a�,�[���"��tn��������\:Wbݖ�v��e6�/ޝ�������s+6D�ё��oँܤ �kv`���đ�>���j3��f�m�j'7.�*���z�]�~�􉟍� �+<|�#Y���ɤ;���L��_�u�@�/��z�VY0���½�����O����l��u6���`����ٶ��t�Y�kO�7����tƌ��)i�\x��
��t_gW���]jT���2/A�x��t�d�Q`jJS�E��я���,�=��*.p�u�E3R#�y��K�+�R���ޕS������8T�'���iΑ��@�T'8�a�&�;V�D�Z��u�m��@?+�u���Jw�R���J��/��!
#�U~���*���X͢�x�G��(P�vMA�/�{��5�쨃�K<RcDƽT!���K��l#�r�R����i�L�n]�M8D	�/)c����	Z	�����X�� ;#V8ݯ>���O���P&��L�@J;��장��P���+(\�KY�Y��͟����7�d��,�N�Z��)����zl�DQ�"�uA�P0f��w��v����`'�޴��w�42_p���O����i_
�ļL�(�E�R#� ��A�xܸ	����|����GVw�C>jFθr�_�4�}%A�rq�����z��5��6$�8����E��B@嫪�]���N[����H@�8�gE�5'VD����z���3dd�,��9TE�������;��0�����r�0��A�N̔�T�`~H,捋�����>X�h�5�*���y�J�R���ː$�!@{�h�̧���	g�o��Ob_j~�N�"�5Z�w�>p겳��f�p�\tV����\g~H.���UW�ӷΖ��w�ʈ�qgտ�5K�!��?��B�)@ۛT '�L���;�e���a��Y��d�~C��f|��qg� tDd���/gW9����"|l7S�w��Y�,�?�3���cE�f���,���C��.ت@^�}�Y�n�䭺'(rz���s]H�t1��8$�o���j��C�)0�f^XD�B�WL��T�|\�*8D�!Eq�������b���>�jh��Y�� Nj��9�)��;��tXd��ɪ`��S�& -�F�&���3OâF"?�)'������>�����n��&���o�[l�3wS� �ք
�����HṲBG{=J��-$��P�)~۸/����K�{��t����ll��7��G���׿:�sU�ļ��.�(x�B�tJ�I��")��1k*��K��4gv�� �+h�b�|��ͪȫr��Q� K��o�Mݔ(��-�	 `�ui}uFM����F"�Vd���F��������"3^ƹ�T�K�ޙ�uN�w!�N: ��f��W�_��N�I:���U��6�%�:�gS�7Q�8�x��Ή@睱D��ؚy���)�m�vN�Qμ8>e�d��&�v�0_��Nm�֋\���W���L?�&��{W�F�yЉ��p��߬�ệVϧ@ߵ&<��f�����Θ)��5��x��b�9S,<d<&@�Krx5��}�\�M´dǫ��K�f�=������ʖ�r�=-[�K;3M�R릝+`Ѳ�$YS�f-Y���d�J���ѿy���n��a����K��jY�z���E͎Fh�R'�L�
���N�-���96}..��?���hO�^��k����	�%.����_����$�~Sf׶!d&U	�FƤ��R�	:+�;���I�HٳpS�*�V��R�=9�^}����Ο���x��x��7Y��͔ħ~}�ֱ�9yS�� ��C�� p�"ѳ����Q�ش`j�K��b�l�p�j_��w����G�&���v��iiNBp�V1�ǟ���6����'"Iv�.�q�5�3�8Y��c��2�~p�}����+������".qk��I �}p$#��w�����o+��`=l�Rd8{��Q�=�n�G��f�����*�r8�0�@�e="+����ŏ�FYXR�?��)NCba2��d]{���'�����)J��ޚ
��`{I��<'�5�-4@���h��O�YN����0y2b��y5{�z���V�rik�l��_Yr�b��#l�s���
( ��#.)b�j���]l����DT������E!c>��x�]2�p��(T�n�T��]����N+ޗOF��ۂ+-����*�F����A�n�h&�3W3'˞�v��=�]��ā��R�/�ِ,��ݺ]e��3럿�kj4F�X�R�B|�1h�-�1��^�w�Ԃ�?35�P��๛_��N�kq���}�������)N�=y;>�2FO�ؚH�L%�<w�#8O�U��㍚zb ��t+����8� 8��,ΔC��C'�g�D��]D�`�ș��n�P���%�O�M�&�3���<܇&�d�X�S�O�!��[�tr[�+�����#�
6i�Yu?j�ԝR�� 0�
CdՂ�S�4��\4�~xP`���]��AH�8�s����^��`�\Z�\v#�\�p��+:�&�����u�s���Xx�l��Z;�E2���^\�l:���.P�����р����9m`oVe�;��'��RF�6�9��9�b��i�t�_�,A�"����O~�d��\�6����j����& *�������fdԜ\���I�V^t��!�ƕ���W���l��a�A��gxy�"/��2�֚�K{6�ĳ���v�j&E<(N�0�d�]K�ύ��h���'�����ݾ���������'���s�ڙU[��O��#k\�N��>%�7�C��]�A.�	�s�/z*��Q
����X��ɉ��>n��Y�o�|��������5:	�'�Q)����>"n�=�ߐXO�M�.�aA�6��Opq�AH���g ��u8��] _^��ڤG�Өoa�$��z\�j�%>��AM���n&{q.F���l��Xܘޘ��`)
�5\��EEr߮��� ��lL�aG�q V)�V�����;*R���v����rYٟ�/���ON�mʍ��
O�?>mo�#P˪�� �f���,)mJG,��]�τ(֌×��7��Z~Mi��a��)2p���~�x��dd����}uZʲ������zo�_!N@<�2���Q��,����?���V1�{}�ؽe�1��0bn�V
w�	&݊$9����(��z�X2��f�s��g�xؖ�e:�m�����1>h�ػh��䮾(�*ߝ2h��5����J��^�:ST��>Ďb~�Vw�,q؝Z;��$��������ew��;�D�bu�u�N�*�
m1�US���*���S"�B=�h�`#%��M���/_��}03�x�M�����i�ɫlW��,h��E�Q���:� J�(>����H7P�Kn��Sbz��dw���#SJu�?�n��_����,����.�5��Z�̥��g
����!}��J����H�;>�i/���<��u�s"&������v"���/���1j:�7RJN!@(��������cy1�5fI�or��6%C8�dm%��)Pf�0�ⰶMVI�3ψ�F�2�FwFN�T�_ě���GYE����b�ը~R̸�F47�\��(zS���d~����hR� ̓0}��a�N�8CGms�r(��g,��H�Rc�'TcX̄0�[wH�ȸ������ۂsW�#���A��Tz.c�d���m�Λ�s;��$������E#�Zr''�/�зʆ�p�"2B	�p���#�(�I�v[�	��]�e�־<o#����v������{�0�w�(d��5M��*���ls�;�޹���ž{�/����˞gԟ�t���[|��%m0�U_��+N� ��	׬�²��k�AE�W��q�Y1v�L���Gf!]x7e�DO~=~n\�D�a��:�Uͽjd �*\m�P�jT�;�3���6���ەC�����xdssdwa6u�V!�?�"��V���h"/~ieV
�S<�k�^��S�Т�dЙ��l�����T�a��֧b`����<�2Y�D�k!5�����L2,wG�h4�׭+�/�A3>6�}F|\Ja��.���ETE����.���
������&˦HJ��� J$��(g��Gr��wWk�e�Lv��]O�"A�2_������`y��A]�YBzӊ����N���W���)s^�ٟcd*�JH<��ȼ�����W���f_;1���^�]9��1�� #Oev@��,�?Du�2���|�/�M ��J=��<�'��7�ll7�;���X��y��c	VKՓ�?�^ز��������-6�lٺ#���t����K��I��O A�u�9���=8�X��]?�R������)ob��ܘ{ ���V������� Tv��$�$��y%��s(q\	`�p���v�[��aj�](�w�Eb��
�C>8��ThsMC�ڋ��R���dfM/$�<���y6�
�`sGXQ�ۆܨ������+h��)$�h�����.d�-�W�^�e��L�q��b����nh']z���[Jj��X˔* �6I�Ϡ������ ���&g�0e�\������4FmAZ�K?��,�usܦp-Ğg�K��;�R���t� �����1h=Al6�<3� E�m8��I�yD3�)�7�3��'�C�²�F~N<��c޳H��/�!���U�%;B`��CО� wM��KU�}A����~֮ j�8��̨e��ԣý��u�e3ٯ+�{ԏ+c�hk���?��������x�=E`�?)�&<	<+Ȇk�F�}����|)+&���q�$� u(j�R\����Y�Gq���(>#*�����c�9��8��d�^���%�:��"���E��m���^@��5��L��4zD"��#��o���J�$�����;ɲ3����b\�5�t�6({����6�[�����f�t]��5�u�1����	v���޽�D����PswC����aG���*+�EjT�G}~�2w�o���d����4J�D�1�'�1��tOb��ƫw��Aw�.7�۱@�֪���܆�&���y�Q����hW��F�+�K�z�$�:�x��C/m��|�T;�󸚅RA���,��T2<����8ĭ�R$@�Fى��W�*.�}OnB5YHk�Ozz1v�j��o���ѷ	=U�y5$�k6l��=�]Ȏ���c�`ͼ�rɣ��@���;�Gg鷪�����;���_�ڡq�8! �Z���񩓁�ZB	�w
W�L���T� �)�KV�R��g��{on�crv?���i�m���}��x�.�M����t��3C�X���I(݄����醶{,�����*���S��%L������[Xo���w�bF;�\fÇ�d�-�O�˰=B8U�j��/�dS����L�h���������yG�ޗ�h�S��Iu	�mb)B)�����@8lh�3ӌ8�j�8M�2��M �vr"x����N��S��^����U��cf+h�e�
�[��o�@'�/ �,�%����!�_{��8��$��茶M�j?���/--!�9^��lL9b��Zt$��DˈH۝U �,_{�O�y	�K��M��/�Ū=�Z��`��.�"n���qj���R���A��[YEU�P�9�B�Q�C�V�����u��8%���Hh�2Qg�f⧸�E��U9z���7���ʈ�����ğ�\A�q�k���
U�y������(���}�+���4^�h$K���UM%Pl���WH�P�����aʍ��LeƠ�����7���*ߝ®��[���@|�1�3�x|:�@wN���6�H�"	v�(<0{fA;��B�׍llI��QG�	4��Ius�DL�-���S���H��~%���'AZ�yGiT�p��S��J�a�7�]K�s��"{e���`��Y8�z���Zu��;����诨ICj������J����� �,��l.f~lB�s)-m\�᠙90��ǥ	l��}��z��F��c���+�������?M��Y�9Nr�@�E�M�D��t�Z�&���T�J�h|�/y�4�V���&S.�m���@$m�G)�s�F����7�6|����j$�f���0����ԝ��_n?�s|fZi!w�2����(9�9��<ʯHXO*�QSD�]�pJ�;���
%i��=��\���f��r�	}�-�u�=j�{��<�_�L`$����G��h�v����Q�����z�%���HI�O�㸚�	~Y? g��dQו�>�����[g�M!�A6��!�.i�P�N���:�$NZ��d�US. �E��i�#8�{"]}1�7H<*�Gc$��Rܩ&Ni��V@��_���B+~,k��^���e%v�ʺw��K? oI� �ݟd�{d��f���7<P�d�*�E��q�rS �?G��l�,�c6��<Q�{Zy��N=u�/w~��DEi�m�O:E�L�=J?k�%F�i|�%����D�䀲�bq�3�Q���� ���X$���h���r`�'-��r���? �r�'h_�ۦ�k�szl��a�ƣ&�u���L[k����\N��Jnf��Kj.�T%Z��=��x���{i'�CL�}O��!���2���S�?(�s�SQ�f����Q>��9�Ӱ�*̣���z�������:7�E�Y�\�\�|p�۳�:;�-�������R~A;�\~cPf�����`5?	�MÆӁ���B��E2���W�Ⱥ_iF�Y x�x�zq4��-2}���~a# ~�r&@|�']���O�����c�S�]��󎕠�#�c�3^f?|�e\�� �#v�d��Z�H]1mÊ����чKl�7X�Xx��?g�?�4��)�r��k}�J�c �˥�{w�a�M��H�|����@|{�b��%��+��I�5[��^��� S7Q[_?��t� g�v��y,t���|l�GG�q�f�0�n�uf����w�������^r�ؘ�]M���,Tò�\^>>N�9pg8�5���I_죣*xs���D0�,��ϟ�\;�����35�ё執ne�d��Ce�S�'
aʗ
��w;>�c4��~�%\&����0��q,a�/Ȫ:�'�@�EV~jt�$>��F5��TB���bZ̾ޛ���=���IJ-���w������x73	Rۣ벀���%}d]�S����%��s�� ���׀�.jif��7q�`\&PV-���'[�#�A��N���!�&|^�	��a�j4�[��~��7{<L\QܜL���GsH�u,�1Y��O��I�l��8�ֿL��(�$&��ȵ�t�̋.�)�RL=�o��~�����B(ͧ�Jۡ�Y&��eh��=6�ï��V�5$QT�F�W<5�-���1G�l������U¨�PQ�<��:}9�\7�UҠ=�[\	�t8�I@���	JC2�3xS��X ��g.Ő77`5��Iۭo�k��U��E���R���]�jN���t�p{q ��Ri=��3��Ҥ�n��?��r1G�@jb��5�֪y%���������8V�ibR��r����|�FP� �7pd����*�&���x����+��/@W��������5V����F�OE\����̨���*�0ں����.;���P���Дx��;�%ꐚH���gX�<xN5+�fl���o�ߤV#T�<���ˎ���W|�����@�~�쾪��T���'/0#�2C�	A��\)������B3�.P�ro���
��������e�h#���E�ή�
M[j �OiY��V�7.����ϽW��<0a>�tZ\�Р� NM�ؿ�����GM}���:g�Sޭj�Ny�m׎/ѱ5r#����;v�A[zAh�~z�N��/_XG.>�����3��#�M��;Sc��g��4k�7�����X!�g%�X���N��Nt�Y�E`ib$n�.�Sso\��1e	�K����v�HM������f]���1m�[���S�y�q�y1��ohg�+����v�l�H�C�Ҽ��3XUd�+I ��q���8�ޗ0}7�W3h���E/߶oFǄ��y�9�d�}u��'���0� �)�r0|۩�D�d�-�G�$=�T&\��T�N{�����=��"���π�fv2�=��L���O���y4�_Dݗ�E!��d��u��g��N� ���C!�������
�'�;�t�dd�U�oǍ.VM�;�)Q��w�H�
��r;,�� �yY�R�~Lt���4�����[���٨R7�W��,�kՓ37���jT�?b�<��<{����.�b�;e�V>�ML�x���9a0 ^�G�,A�����vb� �f�T�*�=ě
&���� a�K�Sxʍ�'���H����v'����j�q7L��w�ʭ$��Y��',��z����^K&e��\��e��P��uM�{��+���* �}X���p��7������Z���+S�%"Yw��O��,�<�{W	�E��Z��b�a3-���ؿ����p����?��x����?#&o<z��L��,+0v�ۅ-��*bZ��h�+�s^{&=�D,�xNH�������!��ڇr.k����Q��sF�$���:ʿ�&��c�����$"@���W�75G+s�>��woU!'b.��n�����(��P������ BvEZx��`���o�2uz�M{=����i�d
��WZ������:���Rð{�D	��Qrv/�O�;����1W�ձ�x�:a�dX;p�2V�,Ej�D�g����uW&[�hT}�B�gwq���μq~w���\Տt�jz�a�s#�Ӵ\�ų�~��D���*��x�Ux�P����TA=_�hww%��q���/b�m�d���+���כ������8x�W@ L��������װ��q��M���ת#�!���ZV{��r?�s#6��QǲڎA��(:���j]����%G8Zχ&��1�}W�����:���5T�Υ� ��}�n���!�}ci����#9�:�����(F�K8��0�PҘ��&��=D�BUe��qW��x����2���ۿs#O]iI��m��	�e:@Z͚@����x+�4 ��I���H �j{_"��4���{~;�7t����x���@�Vg�W)�d�M�1�YK��k�T��$��\K��8O=���6l�z�}l�H �4x����}d�h�/��g����}5;u��#�С�I�H,�W�7��K���.�׻=v��6�e�t�*&F��s�04S^t��	�5&U%�(
#���AV�XAHc4_��lǾe��dENc�	���g�������{n���H}���FyZ`�GŅ����\TO��
t����}8�F4��ؔM!�=���aS3����E�1^�A㔤�s���#�e@�f�2	sI�e��D�l�	�(�>U[���Q��bU��L����R\�a����5�O9�/p�xIki��hH�] �	�= ���.�ztdq1v����;�&�L��t���Y��Vy� k���{�яz�l�j��7���'5n�{`{��Ì��A�|����?���I�v���Ax��̡x�ۙ�O0>�f�4G���ԙ����6����cC�E���Af~�U���b�-��UTf�s�Al��V�F1�xь]K����|�x=���vĶ2�,�^gմ��[�g`�	�Q����v�3���J3��]mO�Xړ7OB�@�mZt��,Z���	=���[;ȝ"����u��a�F$_c��P�Z�k�(M�"�,�lἹ�Q�KJ �k	މh13=�\���u ���h9�� Uo�`�4��R�2f^�Ԧ�{K�z��~�ru�Ʈu���Q/lKj�]�9/�7fͽˆ)���5�v��3�)���d#����ʙ3C���r�6F	0��H��0X�:���(L�Ã6�;��s��b��ib��ڙ��T9łȅ�K\��i�O��)}���t��|Kl rTzϓw�I����.���B݀�ZGQ��6Aӳ�=9�>u�!�Cјh/�YX}��Y���yv-&]�B�u~aJh��q���p!���N�d��� �#qh��韝;�VX�G�5}jOq\`-��y�3�ܫ��@i���(U��I����h��x�J�t@��L��O�`&�����m�T��=(�	���	��]��KDF�����%��	��]v�}���r`C���G	�Y�&��l��[d~����r[.�a-�R��C̷�m�O%nG�	�Q�}y���Mf��������{tx��쮰f8��v]�������p���Ƌ��e7al㐷�T���XJNc���yB �'�4o�H�rax��Ra3�7��fN�9RAV2:0�2a�ťӋ8�^��|�vi|U�O,�|d/���-t��D ���V�9FD ����܎���&�R�^GK�_��5 Bis':8�(��8J�]��<SF�c"Gu{���Kݸ�1� O+Pæ?��Lש���C�ڶ#��H/
C�2�����֗A���Fݶ	�4#zh�=�����?r�8�(ĳ����h:�5�,������(�oQL�`���W�%��A�D�#A�udO��7,���Jט�-��&�nD����*]����^M�����)�F�X�C!�D���,�p�G��H���t�P'�ұ,��Y�����R��e�`��p�!�Ƅ)�Ή[��L�l��|?�w����eL�:�{Gþ�`@��Y�|����#�0��~� �,�ZH��!
�����ZM���Upʸ\����{`�:|&�7�)���V�u���g�H����A��0bo�;�E
��͌�#V��j�f������ۂ�w���w��X��i��[���Y�1Kr����՞t��&�"���.VC^MF[Տ<��1�Q�Ic�۵��~�'F���܇�]Giת- E;�:s��@�~z}��^
�Q��X��Y�4�0^�]tr���2V׍�w��[C��Y�5d�'�G!�y��� 	��gH2=9O�����§&:Mw¹���qāk ��i|8BL���H�;��Y0TT����X�������^T��"��{1E0341�r�;�n�j��VT�47\ r��$���bd����6 
AHؾѫ�N�ixJ�NH=�$�9��� �`q�@3�͙�G���Yh��MUt�Y8SyDza[��%�6�����]��a�f��8���Q��AI7:1�a<�8z9x�J!p��L�SLd9d�XV8�����͔�)�,��6ӎ���F�M�C���b�H�LZ��,3m�	��V�!��=��Օh�IA���/մ^���c����U�.܉ft�pȅ���w��ޮ��1�9nQVF9fL}�Ai��r=VΚiuo#����$ M�R|~t4Ee�����#@]��.�*Wm5S�\���X-�a��78Ӆ]��	�0\�'�_��b��Vo���a���,s�E�d#ϟR�i|��3Z\�gѳ��Z�H��2}-��D��8��"��9�����-I�������}j�
�{ٿB��&�޲����n8d�^��?�#g����X�m��ZD�-�{����/��bӀD܈f�BI�8B�UIwz�=��;5f���`���r�c,ַ�ˎX*28Ģ\-�Z�R�K�tYҝ�z���]s�+8x��0\�\đ-���I l��b���1d]X��Os��b|�~3��H�D�7];�ݑQ\�2����J]�Q��W�g92����ǽ9:�T��1b��tl)l�;1�UP�/�(�=A��u�	�8d�{��po��B+Y�;ګҧmSS�A�0����?��j>��O��x�;�e��\w���)�1�bs!�1�BsXA83]bE\��[�Ƈ�.18Tc��Ȋ�}#P�o��&մAx���Ҁ�����BX�HY�j_ee��xϾ�B���M�T��*��pH![c�j#h��i��G�������S��^�L8�n��ӭ�3�f�;�Mf��P��>/Eb���U)�P�#���#O*�^���l#m����*C�)�ѱĦJ�̺�h�(�d��qdj��i	�C��\�g��O�Y��KS�� $��to��9G��\�B�\�'P�$F�C�>I���ࢲ��#՝�4�+�C�1.���i��9��֜��r|�5ŷ�7{?���p����(�������2��Ìq~%Jc;MKT�(�G�mUk�0�H��Fz�� ��c�J4�J~��ZX�Os����g�cG���ruM���['��y?���9O�|vJޙ^'�Q�ɺ@�3#իC��Ys g	�?�����(�u�Wz�S4lIgi^2�@W��JO�g���i{���^a�8�bg�xǨ'�\Y`��-Q=R�׊Y���k�u���a�w}�ΈL���U��q���.2�DD�_�N�^�t��)fH3�s�@	������i�\��N��N~���,�E�s'�0k��ɨ�}��^���H�?o�߿���
�tMm�Zs󰏈P~����ԏ8SU�ݓ��G��[�׮N���֨�{Y���Gep;K�V}�&?ki�HOӡ�G(�3���.6����~�Sb�'��ٵ]����� ��5[W|���ۨ�.᩶�85v��_��A�?�y��8��nD)����8�
�8^�����S�n�����<�����zY�սY�4 �L����9&s\_>1F���Wϼ��a�k:Mm����	P���:
f������^+��� �u��V�QB���K��l�M{-�Ԩ�Jdz)ě��U^���`�.s�����m���(}9�w�t�h�^
�g�����Ho�L2����שC�)]4iE�dlp6�xV�J8�t{���sW�� )��t��Q+�(�_%����>�'��吵�&s�d�T,^%$�����p}9���#�C ̩�!�8H։�w3:�rf �A�ؕ�U���s�k5�����T��O�-��-��JC4��MI�j�gs ��oLkԨ��/�W�LWLR�-s�_��� �ըd8�i�-=NFF�"��&���x�Ί���/�y8|�V�zb,TD��v�̹��1ʴNCە�R�j�/���ϝ��P�t�S�wc�;�W̕��!��f�[���3T0�_z�"���9wMV#��?�KrV�adB'�*�Pi_*@��:9S��,�!%���xF���ݞ�ȁ�?�΃��t����{.	��.�d�_������>�I� 3�]�5�v	�p~��|=�����xH"����f��0�9�������e��xM��|��ʋ�x O�H�'W�ѷ�*�����9�J��N�?C~5����o�����.1;� Q�U<N��,Ը'���(�����+x�,��H:�(�!���eO���O��z���r�����?2�L��T����˷���ڬ�w��w���ĮU�n��R�x�����lۛ���oi>b���ݕ��E1�S�Ÿy�����I?���qKЪr�uw� ��i�/���6�8,�Nz����# �����r�w�F�F�w�+����x{��$�K�����L�����W=ot�e��9��+Hc�0O`;�4k�V�\�_+�k �)����+���╂��QA�_�vP�m�s��7�L��VV�3~
��/7��x	�y]�\~K�}��s���T�D�r5���5�b�~��5=�s�����4g�?e�1o ~�k|lׅ�d:�Ay��h�3`���H�4�%S��`�2hb ��+D4�2���x��<=��<z�G>Q���PO�#�]�jtp�s׉��v��Y?�~q��g�0�W�#�66E����?���ڪ ��/�B��_��Jg��p��=##
#}��r��s���7�+�I��M��������z�1���'�K�n59[���B@��U�=d5X���o��-.�!�<(���Y_�f��ެ|nut��.2�5�`���I�#N5�#�U�xܯ�Ў��d�	���0_�T���g��3�����)��Yi��&Q�)��s���&-���92�I�i3��:�4{�u�(���`�!"�>�v0G�_�>������-	�ٹ&Gg���J?~\)ۮ��b��$r�.�1?`X�^�غ���B�UY�ˬ�
�6����~�X��{X��㫛�("��(�g�c�S �F�ЮqX���ܪ�i|�9�wN&���-��j�0��{�R���Wѧ��V�#�}!��b�?��ڐ�����C\8��zg���fP��`�Pa���}�(`H�X��јB_�I���8ۙ�-���������.ۥX�ǰz�B�I#(�b��L���nyǘ���W�=�sK��v��n+�@暈n��ʆ��rn���:KU6�I�~�]���~�׭><x�Y����\��w�P��p���hQ<gS�|���z/���1���e�oGpD�^�x��[)9���>���2�J�ޥ�OQ7iG"���I&+��?��X\���hZd:��Ѥ�@�q�q��s��7]�ܝ�`��t���L�?���MZrM[��ν�ӫ��pm���"]�z�lD���tq��@v��?��C�q�����tE�mc���(C�'������+�A+�S���0�2Cc1F�� �$���!|T^3ʀV�Zi�ҁl^t�Jb��c�מ�[ŗ&_|��x��vbAkl�s������"_�����ԬDF��܅��Z�"-}C_��8i#����s䀡��Y��.b9pX���G_�6����ܡ8x�r�u/%s�ߦ���Q?c�BD�0��#C{ox��Ȁ&Ǔ���Φ�rH�ͯk{+�����h�A��B+H8�-G�讆�y{!�:G/N�VG����{[<���.�f�X ��n�]�W�S[|ʯ��9��X�_Lm	g�S	�H+@�Wz~rZ^�K��.A��iy�F�;Kj6��Dф@�J��I8�&>?Nۼ�k�&ܵ��x@�.���A5<���ؽ��0���j�/�  �{�<0'ď����[�-g�Vc�&�P��V(�89_��b���%��`[	-���I����9�������Ĩ��x`�U��!9�$���Io��&�䅇�*�Z8��Њ�*����q��#�QU�z�H#rR��s��,U7 ��)�:��#`/�1�����s�c�S�ywՕu�h��'����V�F�a�7D�(?f�{H7mY��@k��L��寲��*J�:9�^k䉊b:�]z�4l:g����YJ^�=B�놌�^�:*y����ss*�n���GNqo~}G�t���S���U�E���zw6hı�a��� ʲt������/�8�̡���Ԣ��bˍ�\�o��|��_#��?�����j�w�:m�����!��Ohus��ZG9�5�Ksz��r=Y��PUu�1�b���Լ��Lm�)��{�>�(�u�B����I� S��^��,�n�K�Rk���x!ڹ�mqφ.o�Α]�_&�G�_r��|���1Bh���ȑĹW���3���K��G�����`�`-�� ��;��,c�:5�̦���x��Wl���� �� ��mi�����p��Bu&�wO>�0��Է������gV��f���FFU�)����y��st�Pi�� �N(��t�= B��ص�0,�o��T��k�����BI�c��cK�D��8���:�e]�r=L��_1b��9��U�~�L��z�$��x�H�P2�h���e���h�Y{ԎvIStۜ�@��5,T��S.Zf�@���u$!ˡ0���9nEE:]���34j��H�Sف;~�ф��԰)�T���(���t1_:+�p��u�
�8�wC
�,��C��F�O�C!�%�ΣD� A��@��ٓ����$��֦I�-V}�CM�s]�q�G<JSf�����h$~X�޳��R\~sz��RVʅ���U#���(�k��
��4�QVM��Y�x��s�[3��C��&0�D�ڐxH����h�|*>�Z��W=z�( � <�׾Q�|*�j���y���~���5m(V<�#Qa�ԫ�?�װ��s�kp��/*>+�X��\۬��WS9����n�?����[�,�3"��w��C~��v&u|P~B�R	�zh�h&�v)7< ��z��}!y�H��E�ẻ� C³�����Y�N�X���c�*�[��ݐG��iȂDL�0��@��/P,ƛ���_��\��9�����V�t�~��U{�Ӽ<���~}�7�U�(çQ�NL��CD�\��M�� jCI��_�I�hM[ƻ�W�wW�a	���4���(�̓@�G��h����-�K���<RX��7I��-�����
�aɛB���?�}!�Ʌ[Tw��ר�^�3%�=�4����a�����Lc`�Z�9����{Y�����B�"��W>��W	�Ի
��>�