`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
MotMrfVaHvfPhPCBZPRW2Vp7/sn45TAq1NJd/HSb9eBeBkuGixtKwTbiAQk2mS4GwPbvYppZeKgV
bQTCNBAL1TXHzGFJvb+WR6ZRs0VZdxhntHzqR6rBxwdiJw4uj7ybYuXP1yQEeq25c1ZYI29ILrmx
WdqNX/2NUPpdOBnICE5PNoEbp/esAIO2T6VnnhswAOerapuSA/9EiybepavGk3oADnzOJCzJtKmI
88EGuDXfS9HtUxM7Zd528pfMM8AmKjM4sHVJBqw6ZPxvcd+Z6/FM1Vv+QJ2MhnPy9g92yVkLwmGX
P+KaCgM4yS4t5Py0KG9VaUCG15scsPvIJObFBQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="FU1L9FRs/Osyeis6/39QAxGD+zDK1kJFys3bwoMN70s="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6288)
`protect data_block
3THTx/qKh0GvbSLmw23XYXdlDciBGyePLDYL/a/jcxZ37uVYpDUwWyR4MmDWAM3tvfFM0/mQ6Auw
iuR7/5557+LIKw79VDNqZWEuccgcHCDgdyx8TP4Jwo5SEjEATfjN/3WAexVb2J49Zc3sqJxshgmB
K4wlnxKaQUz99hn07330/Z4baLDMCa1ESl+746xchKhOv0AeTF6p41nz76dwtzjKO1eRz/Hs+zds
z4pMEAycpniEJnvpIcVr/Hp0v8JeLkCnTf6RXoN6DrvYu23w+G5mGj1qFsr6y+xvsCxg1iZCKLAT
wKB3Qs1R34LckX8dhGPBtb+7X1UjBPlCTR152fuoqCE0WJeoiDnoQRaQqoi8q0Jm5Fi8fypoRBOG
xuUL3Za3yHRe9YRIt5VrpDnV3iAXUfS7ifhbjhc4J9W8ZYvqLlDN374TW2n489WDgSPRyyfyqYXf
MXICXUtHr2SYR64zUwhMX7K+KNep6O0MIuyQSDYAP+mm/nx2LnLZTmWHjs3zP/rkdIAHahAeCcft
a//FzoJLzb2gKHARWHkZ+NsaFUQj3Yi5wSz6zOUD3Bz+d29evUwTS8qV+bHMtZv6SNvQdhjyAgIn
Q61mAkqxwcr/TxRWgQ2NDio2uxffBn3HwsPFqhS9Npy02wJIernDJumwSRvwEh3s1OOZd9raWwNP
MlFpGA+Oxr++A/mgKhKx9R5ICbpWQ9tQ4EOZxoMn9ctYbslKa6bHC1gCbkPnZKr5p7L4OnNhfww7
v42gg99ctrG/m3wrqXRjlrvUss/n3Frng/KzcOlk8CsoDuXMAa00e13d7KbSgWi4evGW8fUWzLdo
eyYxW9yA5WQu231rrPGadIhgf1ruUT72P3+GPenKirX/5W00ttvo94R7y9/WyBWp/o2wVd22xJ7M
WJwYGdMjDrvGdYMPABLta4p6Sa1quyP28EU88ng2OeDmvfNHadj7uurKTQg2QgbbYMEUQmtTzDVd
HZ7VfBBdE1p2vpRWwlxeuGSeoKa4aTNNsAMEOMLuZ61xzbvASly4XkcaxKUkFRhdHKlsmJdf4tkB
499bAOV904G4EqNjYvTw+dhgiMv7/87qWvtL1J7uhZvLlAelUBr1TcKBPULrDe7FW4kX8VyndoyH
+xnL8dYcjOiB/KaE2JgQmN6czdxk8mirGky63t6bcaue8QlYkKoECfgvofinxvzeH1wwdlDAzIWM
ikH1LjoMDiAQEr0EJvXfnfqxGsX/mMyNYyAEV0VA44PbctiZzogY6oTTghCSYWfnlLe3VzS8JERo
LkYxUzsxe9otOM/QF4p0n4SAThvNuY2X5bcKbPFmLMni2X0LybzUEeANakcshHpEiTgPL8HV+WEo
CfVzJOrT+p+SHVP71rrgvQVLNQs4Xi3IxNYpgcdDAsWEvLCdUTnjbtVhuyDSfeJ1EtpmtfTcSVoQ
IhJhZvrkyWioq5qoPUWv7Vk65PwvHj3CPu+9W3rQSxL0kTK5jLzSWtbcGjAgJ/fKhb31YHkBRkWi
HoGpv2rGoRgxVhnV1GoIAew00h7ypeRKEx/ytc0Jwb4dKx4wDKicJO18KCM2Smn0kK9aDUpFQaxP
hgh5z6wwiZghtWkhciUUDPxGrV1YwOOMsK2hgyvgF0bAFenEbPdCt2aOOzqdFR+SvLkrWfoFF0Tw
0FnsxRmUZ52cO6k7Qs8cLUBo+4uu8QWisOeR2AzekS7dHWNpvvbBYxJL1pUxD0FvFHpGolLbIu6u
J8P06KfVwvhJhkzoWgwAETNT0kysqVM3QARQC/4E6+20y7GlfozVqmWV0XKHVgowYRblqqn8qsOW
ZlNJvqlCmNl2t4P9E0R/AIhoz3ngtKUTI/JNpqATihDC+yYZY1Qlsm0JAnLL5xxRi2sdbqmRhvwN
UaQ80ph95aglnFYgn8g/mM7JEvVp9sHsrgA/i9U8sLdHTYpcluu173ksjntqLV1dyR8uZbdh8J1P
evAErS156Q2s2YKbkAYwooz0PFbi4qPvYMDvzW0w2Fy++q8LkU/XF1iAEpt3MpEy/PnQodUwTwhK
Ci25roJKsSf4zi4sN9M3OPt/J3/o75sMrEh++10alv8A81cYcw9Q9+RxFB+1e2L0tynl5UkdcDxo
HJPww1oimekABu6fXBDnlZ6aLEuNgQWPbMFebPL0tnH7SXamQCXayjMXYQ0ENt1Gu///SFNjqa61
fo/tcUv7p/5okyKw+hWgQwsRcFiaZvMuQfOz6dbQq8MzrUclqnHXpAZ2vrHPBTjhNNpM1bNFjq0o
9hpOFglEDlG6UvQscfujmrnSnhaIllWx7Rw9qWSIYtENsqTG8vpwAZKvcwcfsDYJiSEpfXxI92+4
3bH59K67h1rOc5DD2VTCPKjNza9xERBDhMhj4bUdA/VfoRRSWnwJseRoG4zWXEewidPEwcAOKAbF
09CPMOKlhB2TymiU1OOOeIl5v+aepZOY+SVk4mqJMgp+mURSQ/4i49a5U9h4OWEO14MxLsBGD8Qx
43wuElqBW5PlwAAtTLemCdUog0uvsKXhbgZHlttgxvYEwDGU6uRt/OFEak9rNmtIbms0ZoD9Zw+J
DQYu3mS44oOcMG7ZaHVnd9y5Ibd8el0X1yWcgHk16zBdbes+eSUGQPDNv2osF00hD922P+5hBolp
7xei4UbW2QKkXgEfWunVTiiBK3/w9RRhUOli5Mnol6ltYpRDpre26LbJvtIAlHi/ZaYwl71TGoXN
+RXQPdho9J0G2EKfFq3cUtyZ+axOQEcONTT/gm69hvnMJLUXSNGiJzF9jCdW0f+5kxkkMtVGu3LK
Vi5CyfVn+OMT+pQjRoIpwTUHetSfVgVtJ4Muh9qBwPnGR8PzJg+ymrsjQAGfciQmSLGdpgTQKQ64
jGhYUFSGasrHQ0Os6fLPFeDa/VHwv2F1QoPKzUiBn0SI6HV2fuadxGlyTm4GKvO3i5ZKzxkIsBA/
GOYWm2HvsFf/oCpg9vzl1zF+m/aBNdaFkGRELUm6X2lT118+DzwkmLZABv+2aCVCzKO+hArW7g4k
8Z7OIPJ7EvXso6RIwCRAkVFNxn8sa2yZcDJVht85aopNsmDa1hRANSsNjvMRGRvmDjM1hcFSOw60
codADu81LrAMDd8+IF9VhPLN8elPW17WXs/Pqcgsm4LPrkwPm09Jfy8oBIsyzyvzghd0QHpp06QP
5kn6QCsI+/pe10mmJCGkgw0ZPUiwkKkSzKSUkV2qtG55Rhbhyi8TUtqAT1JUG0KGhP2cFRR6rXw2
FXXh0QwBcbaaNOl6JRCZ5N6EY0JdiA+GC6uSudKURWWerCfGE4GVO7Ej7Dlohvhws3gn/Fvr5q2b
80Vb8dXUoL3xUVR2Gab8jXVdIBp7vP72KhUwT6SGSH9oAuhmKWezqmfag6uIHkGrxZEkFips60pX
bKz1eo9uOllWv/LSBjccxwrrNGQ1ifY1ih/Z36NrH6mnhTiNhXbVV+4Vdth0CF60p9qDXhsMeh4H
UPGcVtXCv0wGVmCFudKlyEWCd83qIH5fNnQZI69+gz2jVYDPmgEl1XSj6nspoX9oxiY+sohUs1Jt
TTNsH8koFOD4u8RTlf6yINHYq+WhpzEgJD7Kz+jSrOBo7yHXSMhp/GiaFLohtNslyfVQ1S1P7UKN
Z9DW7ojcEwQNKtXR2mZFIQRdFGj8Ay1ZZHRaPp7pn8i2d5588jBSfm0tQJL4bDoayn+Uc/W6yHej
MR1W8a70pt2dVbc8O6ewJvDX1w32Rojd4fKLDCVC3cajMm0IPilk4VBeCrM9RFgQw2aN6pE46Jk6
bKG2SLIE9opr07A335AEMXVq5U3r/2USZPCbN0Py0YFYouvzcfN76a3SkuLJ79P7dCnoUoK3IxRq
f0f2i6QQhtx7gWbcKEFwEJnSrTqh7YoGTwBCT4j9RLx8/VsZu+S/wb/LI9k2ENOs5CSc/ypAoHRw
/CrQkBbeatzTYMuH7QFr4sj96nb1fqq1iUd2I9Ka9Tgla6HPAjd5NFRAlhXvnqhlL0fgt6E/VG9c
ttZlLLudubQOuaNXO7ySv06i5Ul4SAB8vRuaDhtEypb2Bo9weC3fBZLbsJSKfdfdBKlqpmxbFJhl
JPj6j4SkqcFS6z9rBUZb2K3NHpwXaeTpdMBwGE7+XRGJWCKj/wT9FPaKCtOLRIQSBzlL0fM00/Lq
eBpfxLszHVXVcfssT6wItlkBhOvR3g6pAqZ4rkSYd6iY2OYe9eAmByvH8j+Gx+DUKY/2gUtKdWfl
pE9bPFDX/WwNebDhYCUAsa2/rhxZ6ueQ/GPdo+ZponApJG4Iu8cp1LmzZeKtlI5vhlfPHwvWQHC3
dr4pAJCGPlqCRrsqHP18cEM456dQrn5ug9Fn9G1X3bCOz0bsV3/wx/AlLvIrH7tLD7jgshDtQf2e
1Yzfk1Udj8ISsS5bRHq7C84q/c1+NxJAi0YnYiSvYmkl46LKy6BH3285TP0xjOBRv+YLrVniiQp/
r+4tvvg+Qt+YVMmKrzzea7wytsqrlaEWu1sQi9ciYLHJ+obBmhmlTwylv2ShRoM0+Fp4i56ZweSh
QBAMwUXb9kfvmw7q3XWsId+s3TrUf1li2hBsdIDdUacVYyR8mrslud3lZfI5r1J38T2EnntzQ2S/
yIkVLZJe5DhxCVEkcl7xlI3s/3/DwcmMcT2iOMNRqunbS76RQ/FkSrD63MqJrSZgJfbQRxWUX+Lc
tux27vL7u3KWFajC6KcsAYzLNYfv90OQAghWbZ8gCDiLZg84/5MJeAVdiW33TfPYmyZrH2pAtB93
gnDDOqi0NhWd3daicO1GAvjNF1moZyERCFC6n1BcolqtqSptHyr27DmSk7Db2bWorpqLjLrm19z/
J+fJmjt4R0WbYil+MqCPDfho2oE78kZ5JO9AjO9icxPeLOfIbI5/0usJRvxSDQjHPelJe8CUqOl4
gpZnA9qUgBW1N3ObQSbq/fOEXIVNRnDQSMCD7Xut8caU1FSpTc9d8r3k7hyxpxZYZiIec4vIkOEK
QJTQAhziyCdvTF3cZfpS/Xce3t5lwd6cbl5i5mdx5DjQNaKUmE0n+m904NCsdjvTSy15yv/ut25s
88HFljIMS+Ut+CRWa6Fx9X+86ZTki+4r2vrtwfcfzj2f+YpHFEm4PPyziVEuAmc/MN7VE74HkfTF
181YLAC2lpOlCyPRRxe/m5mY2bFdmyRGU0lTQkH0lT+s0Gdppv3PCDfwHywZavumYwczZ8Ofg7eX
niTkCf4vH5+Cnr7mNGTbBqRTU3Ln1mISFT3foj1+qTWnjbzvRFwZ5pFv9jxHLSDhVYWVgkvRHCPy
tiycQTMneKOkxhWzx9hUIX0W9+BzrP5xH9Wo1gh7dmXl+qmEY3quJ8mWtmDfKk4LvNmAq4P/LcAS
2yUKXl/Itl1mlwZQQGLrGULY9qryLLKqERwOMsBD7gFFwomjXBq+3IKoHE0CJ4yMjARtl81htZD6
3MUUbNdhagZy/aoFu77c4MoQNl9S6KPt3Jz6SUz9wiDNc8GzFybwMb7kKwRcWbAWJlzSOzn8Ti7C
vKLl9JmSZFRFT/3ouzoPeRfxQqPCqjjrezqcYjcMPcwb704zYLW8Ex1Hpny9SJ0CFfuekXKvg8Km
5kAN5mggRrZhs6roKtwnn5QTZsqwVz9CdoH73TpIbvoXAFG8LZnC/HQNf2iC+Uua0qxGAQUKrk4J
RhgZabx19audvxWfS7pFHqLkk88IuoW5shD1Ga8HiaGThGVNvw98gF7BWpz0NnCocQFNs2h8qJQw
nMV5pdfmnEGw1sJjSLQISRz2dszqdlUQLw++shchlr178V44lC6xBy6P/yb3uP2eL1ki9qZ59s6p
mOF3We7c+FzgUJomH9Hfs63lJe1DObKtPHsY/g2D+xh+ZJcYjFP0HkAyYRzQZ7rpD+yWDMsht0Iw
v+bILL+P1Ur9u4/CUbOc7ua3I33yM6ZKGGRA2P2/+ni6KdoW0ExAI9n/NG6pF00dVOjE1b+3ye+Q
KgfdINjJGKhOf514sckRbTv+4iaocn2upBvl+RXK/l2e3Dnkqetf6AdyLto/Rk1OJpayoPsqAU2N
HORcr0eX4GJpvv+VU6ghFE52gxDe67XlAcxiJoz2M7Z9SM+lE7mjg9PjqvAGJw56cnsYx5FLtmp8
t59HrehfDOSd/gRYE//kEMstsXz6aKZZPVer/Mbvgq3Ky47nyIImPapeKFDRIv/JNvhy6o+Ci0nt
iIodMkmj49foeGnRBuF8g10lSxEqHj80XO6hRHiiqf0E1Wk2OIzcfhpAwhmGEsKV5Wyq2c/Du9dS
rVUYEv4j9E+IEdZcL/aiIDWCARr3n39X5PGO/xQnOcy/r8kxutuE9LyDO2yhamZr2YtrztHaHU/z
U7jlWwzCou2vqKjj8YTmP601Du49Q9A9Me32tth90lUtUXJpxK4LevO/l4cxnPFvyp8Xm6whTnmY
HT2EspfWYq+EmVbDkVgupp0/rvU0jRNNv6XtSmVsRFkeqXWgIIlderQJfaEoZk6EsFJybUbIxKUl
ilY/IoCvNoNOlpEKdCL/BTFV+60ofE/MOdZ3/PcDiNcAW1DGJzckK3JYcwaLv4yawJnvZ2ByggxD
GJ9uq30tp17v5eshHEtMigUDWUm3r4VFJ8J00J5OynGJN930Lz9f99x4lrkkqrmj+E32YsQsp5VN
6MIC/p/qC9FqCsY05sbZoyAJkbfLBIasxIcUr6LemRspQYHGPuJiIsdMGueejgM2c+BcwhjNRSnr
jRfv0/3x8zPOB7xRvbDmC5Z3SRtWAAtb46lBYAYS6ma2yKjzdEPJndPAs9+oXD8+KiwzbpJSnNZm
/0lJPuISSsBS6w608AF4HEydyVrmnCSOTCbcke1cMQZJq9JXsuUBJNeyjz2PcOZFjm1sp1Uh2N9Q
6iwXlsu3QFrfB1EGOtEfX1cxJimIMI9Y5ry6A3lbDZ/qZUuAYR1duW5gb6l00hQKJybgeG4achAW
LeWiu7r+Cd64D3I21V5gk9/ClfaCW4+65+28+EntBFklIcBsYCfyagjFa4Jp6N2/uFJmmkMn7m3B
cROPWYX+KGO+jtzn3F25UNspWhyg0Vea+WbASA8UAshBfhcT10EorBfqLgTdXONBo30lLFD/QQWj
LjLSezZUSiE4m3iJBrCLymcKOGCv2w2Mrs3H2UlFPN+hNKT7+eexQ7r5FeWqBVVbx1DXTe6RPPtd
uo1TKMZjiR10Ze0laFhFucxKB/AHtQGwPmhPMQ9UxqnTlBQW3zCAZWQA7tUvh8TmwUrrBIQheYYq
lLsoChUcBfcRXOZQdDX/lKl7v7/SWOI9BCI+so0SdxGAtn1SPG6OFuhl8L7qrH00B6OJSO+Na2C5
Ly22KpYXe2gzuCmdGNYKNS2rNCTfw7dZPNiD61WxT3eRYCQn5nFWMpqR9IKVI1mlZqFrqUWN1Eej
sUMufJ5CCmeeTnpgp9lLMJ4+rFkDjweWCMk7cEK4Ak6TlcnW3urzD063wnw7Kk617i6Vhu4Pvoq2
kC0L2dWs5FfKiFfXeCAdK4GVdnvY3Jbisaa5ibxCi7U+xfTzguQyG7uz6CPIKIiT7rYm/8gxja8c
0pEafZvTm2FUoQ7TKGUTZ8mZpeoo+cKp5sT21HTmsNa3jJiFTTwfVdc7+siG4S2ff3EUH+F2FK9T
lqwCDro6DqaC1r/0YWcGCONJJ83MBKTkl/FLjJjhbVtiEaFicrp5Pq730aJie1WlgmWiaoUj6zlf
UnkH2EbDvOVL6PHuGoA3UdelyGdPEdBzr8rkI0mZo5CKW9sGOaPjwe191uffeiIwFaJ3LMqzTerI
p2DBR4u744E8mrWJZ08jf4YBl2ULf/e4Uz10MK8DVdMbLlH1yEjHMmas1U5FFnbZUV/AXChspNfz
oVn3lK9EPSCq3XRsqQq4mR6hnbDgZc9ik4cVozti6QJVWrNuokY6ukrJQd1ZMW5vERebfxOUJGKo
wUj5ah8Exsch40kajB26jj+6LEhIrzeeKPa9HlbmP/6QNIvQQDHaDk16+m8Unag8k07rXTUVVSha
apIlNR4gxiauWXInT8CkQ08pSPgNrHVkqR8Td/8mBaCdZsZFqC1M/eNnlo7vukOPIvLA7v5T6bbF
chynfa7EV/cEjFVzRhnJZM4HJoGyz7KRmnd0RSJ7r/6c9w4IFWe4fWWhwdYWNwub0ZqrwJ4t3efV
utyPrW/bVIS8taYp7zBBapzVRRy2eWEPhdFr7mn2vD1V1TKwEvgQ5WurddL2iQh3urJ8im03uMjJ
j92qTFJEOWeGEhnNtMs0dYjrJA+PIJMULUwh3RBGpvBNZ6KBZ4s2yCzaBgc4/9roaQRStiWNwPaU
ICRo4PsvVQcWyX5Q3ZkTX58w
`protect end_protected
