XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��U�[�@��P�yf��[)�4����q�cD����j��O!�#£�)h�]�j�3%��5ST�{�L訋���׊����Z^[����ة��̾����ў�Ǡ�}]� �8i�8�e g��{��F2n�Ȁ�,$�I�u�q����|3�'>0Tm�D�z#f�%�s$��DT�Bt^Fި!]8Z|��aL��hK�	�S���ʙ���/*O���k��
��E/��Hs~
��!Bo�q'&6)�ۭƊ���G1��/���T\�P�<����,�M5�1�4�ǧ����  �쀞��"U��V_���H�����4Itp�oպ�$��@���w��f�TO����� 1�
r1�;D�=�"^?T���:/A���V�J��L�_�d�ڽ��X�|�!��+��h{�
M6�8�(1k^�J��*ǅ�DO�o��5X,`���"�6H�r�Z�f��z ���
l��T�hpyY����ԡO�Y��a;̒�꣥(�	�f��5/aȒ�ruQ}��7�|��O3�mp �B��:��/c���()8�KL�F�E�D$�t+�7(%��Tl�'�ތ�����9�2$e��6�L�l��T�6��[�i�\�Vu�6 do��!#�e����*chY�x�TZ�n�WA���C�f�G��G��h��n���@��,3�����PVx�����_��g������֮�)��{�׏�# z�G| <��-�o��of,i E����}�l�+N�����&���c�>@XlxVHYEB     400     1b07D8�I��u��1�ђN��������E�l��dj�Rx�:����d.!��y���k�n@�X<��7�~~ ���8��a�ہv4�!t�ףR�T�[��g�����Mj�ྶ?�M�(�vC�Mᚋd��As����R;��6ESd�+���O�-�����s]b��_:/~,+���L I�
i���A)�2�ѧ�pg&���L��9	;��\�q2f=������f�7�楳6sSY��&>��Q��w��>tn�9��W��ȣ)�c�V�C���a���TH`�sU�جPR���o� _/��\\̂ٷ618hZȨ�Nk�к�Z3�Ŧ��Ȅ��)���I&ʾ�\��l�4U�\���9�h�L���j�B2eetk���"�p=�<��$���"W�v��A���Eu�p�XlxVHYEB     400     160cI>JV��L^-������xle�m���i� {���w����*O��5��<Ҩ\�#�ܾs�R���ی�A��I��-`T&N�eo��AmS����.�<�fۭ���3[������Y5�K��Wr��d��ٗ�������z�	_��$��x���g����OKD��B�^"�nδ*hb�M����gӟ�b�9�Y����S*���J#�ER�i�)-�F��c�HG��W�� �	-2��� v��yP���ѭ�alP�W��slu(�-L�ƻ�PM��D8��'��q�EU3&]9���5���ی45, �����:!e�X�:�	Nܢ����K�U(�$��$s�XlxVHYEB     400     110���;I~��7��U��ڃ�{��:xA%������ȅtn3������AZM���>� \pq�������ם��.��7�8��rqTG�oʘx�z�4e6.�r�=�W�31��06��Ŀ?M;]��^m��H�*
v2��C4p��g�iF���,4mC�r!P��|����������|�|��JD�*�;9�̟�{�����z�MO�8�ւd*��{$_�9W���*[�P�ql=Ȓ�W"T�Qv�gܵ�>O�p���>[0XlxVHYEB      42      50"�W������QU��H}���X���e���ؗlG�U`
�5(8��+���X�p��,��saNu�?p��W�g