`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
tCwhFNcS8nNgCo70iYPpGgq7mBbHLkbBOmAk6/Kzoq1alxUHbZEeD8AiWIg0ruiQGAO3R0lAoKr+
C4RXczQBm7xfq05PscTyxs7pXhihPNEsqI2C80hzoHpSmWmgSEGTAHrGz29g6QZBRG6J0dOpN9b3
nISUW6dE1/R7fPCWDYQX0s44zayrT8QCAqdctlizLKSVabhu+UsMC0Up/yydJiDTkNWJAQ6EJAxS
qNAARBecphrEdUqHtcbOlR7k6fSo8AzJSfGGNnDaosttlVSBwDOMQ7eZLr07kPwDK+DsF9y2atwp
GdSCinaay9OG95lRrAsQpjrx3lotoFTHM8OffA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="gx/6ZsiZwD1MG8LgadEF/bdjHl07JZDRnLhKrJLqxDQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3520)
`protect data_block
f12Wn6bBt/ljF0JZMtqy9KLXxOr0STbpU8ue2Xugh/SvQRNcWyLg7kPMgPxiWp43R0SDfyqiigVt
uqxqi2vqAaNRQjGpssww3Vki6fmCnPp2SMfKV92y6efv8Cgr9GKhydyw32btxZqApQfHF0X9I3vZ
CTclA8onCBRmXIznCf+GOAx0js3/5/qCRxiEgrOVAToCFWGloe67LYKNlwxVgLoCh8fQUT4zEPZf
4m+IkomXtOChst8C/jQ/noG+N8Vdpp3sBLceq4byGdTSDLlFXzbz0p72M0FpPPWw7eEHc30QxrlR
Y2zl/JXrmdKTnAEDZhql+E0skp0xPXPhPoYmS3P/eVR3oDg0NL+Fj/YE2cAexEAxIKNOS/j6MvBM
63rnToaAu14/z7dtUzm+gYHUEvuAMOnWm92X/abQDFUsjcEpwrFgTgFEIJCTPcvXgSEOKK6NYWXI
v+e7D+oOvc+/RASVMXsITHcKWcp7mfmtgf4g2yIIlXXLN3Mcl7W4Z72WMBmpntb+MQXwC6NssKyS
ksgw0nVK4SVnTC0dbrtSLJZv8vRo7yEWuM7Axa+jt4Q0WM01aiOXQuSjTLazWtyiJLrGTzzn1X2U
X4kUf/p1Q4/DGK2lhGOpWdF8poeVBl/tZCfE2fT+aujUdY3INvRra+czSCuQxZmaqNkoEub3XVgS
zWi0GFuCI8ldEXfJDLgvAPVtqUrUA6i1D9uhn7fiLHstxFZrYci0t1dHIfeC+uOTiLRTYKQgUUdw
XHnx6Tv4ov1PLMUYpW3mgy8AbnECMdBylHewORBx4tN51DRm63yYSGcijJquiPYfVKbK/Ht0nDGu
wsHil8lZ6+eR/zhXp9YOY9w4n+JHSckweLYlzzq8NJo+/ghp+jh0QnfenrgsullsotJhpuONMDNc
yA91REw7CliIytJn4HiYIGLk24BUR5D7eqi/mlDdpqLR0scSWpqx0qeB0HZhbiK54BAMTgFqy/m9
rB7yxPiemIAfOsyqNtqYgXDQkQh7XL3yN4aAr5F6iek8wF99Mwu1GFviAPzMAD38JNbVoMTffGsx
xFsoUQYbkfOqMOD1pX4U6EEMLw8TtsHvMC8iHLpY/5w3j+G+gF2GnYSRab+I2E22Dv9m9otpHHgZ
zSJ1LZDKyXP/RsbQD6OezcilWugmBmMqUPo7WxUGxPWFb5YYgkT1H7AaH0n25SL6hv3yfoaIjBOo
VkqZaEH0qODHoR10SiKfA7/oaDPaNd4100MJqn3Ig2f8Vht5Rln9hMxzNYE+hPoNSRy7Kck40XMp
Gqs32MG7stYdErE98CJCy69IJr70XxkwVLzRxfqd/TMt7sbdwrfzSE3ROtv7LBuvE6i5wj4szaOZ
BsH59dV2MLyI1ZUTCaSmILfF86PUci+6ZCGJg6DOJkz86cpjqf7yIfwvYMx16yzjVN2iQA5R9oYO
15rAGLA5ttTGY2J8XDT/yShhgbvG5k0NH9/aHoYbLqAxw6nDC/Z6I1eCMDocGEoAifRrnWtW7/wc
S0/H6QL+lTLUOOhbw+iaH+AQo7UjyOr/96EdxoFPM7sgFvy9v6S+WKOS+Q5LpRhWObiAwmPQ5odV
gqdOMECO1SXEabnOySQj+vv8nqJXLRnAdVPJou0XnOq2prJ9hTnNVhTD/vvySMe/VjMRIcXCeUva
9PI8Xpybzq5U1k+XgmU9abVYmD9lW+FcxCSZfFVjtHwkF3Xp4uRLCNot7jWVAX/pOwj8liUIkRbf
xnAQ6LfjAKgttLK+xZFLb4kqjNdPNyGholFhporlURWZC/i0IMOv5aOMwPjD0pUVyEaWl//mp4ip
eU2GrOP+SsoO5cfz94hs8K5SgJG6JR0+WijDM9Yw2yenyj/v/peQv74VlSAjazU8J8nrN0s0VIdz
b7PQoYorL5T+TfHnxsYvVk40r/G40bifj78NGVkxa+GoToQms8Z3CYf//yDSpoCWeKJwrkhlFIwv
DqZGWIGjtjR4giGeAVIsc+PgzPJJ9Jv2EM5gSVVnk6E06UREYkE9OO6nlGdpInwFlijkVmj1l9TX
+gqwYrRrsrYohckVbOryuxJplUn/snigqzIJ6lfjlMmfFmW9WyCMufIucwVvP31CzLpDzd1X+CUH
VSypXMaAcz8gZdO+c97MaFR5lhC4UUWHDn5j+yyNH95FPMYvZmxcT02OLKx4ccVra5kuoXiMkpPi
EQjp5qHUag9so28vXPXOm36DdFVPTZ9VwjGJpRHkL2dEO+NGvsLOeKcP+KRHtgrWdmC7PsQ7Jbw0
DwT9HZdmvcHjLtNv5QdhiQsOkD2FTJRb9Hrc+m8DwpyJiCnA2wi6TfeXK/02KSeJWCZmXWaDDWyL
F5k6sC9pWiyBp9d/I6J9GijFzU2jPjOpa2b9UbhPbqCOQ4tdqAO5SnEQ8b/54he+BtmBLc7G+t5y
58P7FUlzXbu+yPtFTY+oaLf5l0ocyMzYMOerwO0/6h0amqRf0VGqJlQ5oA3L8ehqKlXy3Y3s00wS
/gJvwxMNLN6olH4eOh2U+jDfm5U1piYpfE/0hKH2Tiudn1Vfw0PnFk2SguMrkXGdfa/ySAlqACq0
pTLvDNX3JARgkbanofs1hRutTCduDdFAk0Ogm+3SlxVd/fUJcP8Gi598or50ZDYbRZNVY7oCnj/2
6cixI/B0F36/qU4G+EQYamypUlOBAEiq9nFVxLaBlAQyoT1mdHSh6ze4sbexdspWCD19eAZ5jCMK
kINQXPpODPDsm77RZ0CwFN9JjIj0Io2NhsdsZiyEv8UYGvDKesH8yxonEi15t0TMvkZuAR1t94Tn
fm23l8/QmT6fHb3/6zN4gdP0kOwFZ5KM0XqVUr3BUh0ymg1vd8RnCiSpzdazBX7Sou0+9xXtR+zS
J6JZHhYM/WDsDDDw0y6NAzD7T4vp5DoEZK9RcqpDF9DesH8ig+mhYplnBaKNTwcajluYiNm1i/Fd
Y/8lKr86o3CA4GEngwaPn7YtFy1D034jiNerKdfBUx3rkThaOqb+nP4pXp8rntd/XWpDvH9O32ox
EHfgALjP4998CXwHVAyeZsX1sEA7m9LAUk28qqdD8v7uPbXd3QzHD++Qcb6hNk1sAfOxYprGoD+8
9/Ad6Miv0B6/rrPq3gUesw2NmHe3142tc2WLBUAMBSVPjR/UfxkCe5gdLpppcGX20/uPpQJWZQEv
9i4SY9fz9vrSd+gTEYcb+pqAUgYTVDV/1x0RPYS2cPgBITatrKB9qL572mrNJIu3neyXJeUioz6W
j9OTrEabmopR9ZEMph/V7ATjHEmABnfqHc/4p+hiJMgi/iGHcEiSr2ZtVBWhjuI2TtKX70ODIjOX
4j4XPpx5ryCsvTJ9HPuVHFmEC/WvFnlM4DlBFEI8Zm+jr5y0qQpviS7ZGvzJJw0ZmslaBzoCAOXa
IlRzLB+WLPdTZyl0XZTvpM4cYCCWMhqFrgAp+KmIoZlBUN8ib6i8oiwUJSEL9gepD25fzIA2NqVG
J8PDATVbVW6TA26tRJ7na0ZikLC7EmPxacVWqCLmwGyqF7iAAHKVa1MUBMa+WDnETfJ0xpJ+eZov
nxyIYbsdBuRX4uj4kul3rCZBPbZbXExJd1++aR+fkLiX+DlilrTI4C1UKEATl6c6ZnTE/X9ubmLm
uz7E+X9WwyLSYVu0QqYkRkhmbF6DNjyigAtvc0F/rjzn2aDeir5fyVCAwN2g/fabuwZAV4riTdWZ
FNvOzapA8hWysyVzBLy4Pg7QFEs0EYEJW8ntUWTPQSL9xGN85kcXcSXr0aWPE2J4QX4D1IiaVe08
BcAjJl0jidYPvD2ks73OCX3aMPzBGLZK6uSsaep50zxEvbEZQjZz/VRZYZSHMi4opqX0mB55VNh4
5fedfWzsvto0k72nIPSwiNJd+29XA/vavz1Ep6ou2SDsULyDMIMK8y7mz7Sj9Zb1W6VSWbvnG0zl
W9kHWtYO8WHRhbZh8Fn+Um1LYaAyssWC5fWcYKGX0vMk2e2bk09zT6SA+hc34dhv/iG2FahzaHjF
JMkrpV3gb8vo6irYzXBkJoAgXoe6DIKg9Cvod4qTy5/Yc4b0P0BG74sufCdgy4xOb0KNmfLmD4fL
8BYoY16tPNPT6vpvqziISP8LDEwLkM4SB7/SrJMZmngQN0OvlQ+LCG+Haf1oZ/t2BtZnpbribjon
Djjw5pZzqybUtFcjjxUKN0Nb/e58iOU05ebzWSCgXSpWKxRy/efLoZdNFmzKGP/T4ld7kreRZgMG
4Ci/5d3imyxquwNetmQu4i4xztrdnR8wR98vaJSphI9Nd8BXAd/abMStqLqUTgmJVhLKFJc01OnH
4FN4SOHsHnbqS2xQEhFHKsGxHlQyaYMRMh3dWg7kpvJGZ5Ozr62PY6RLKL07wWAnXz7riblA7ONh
2XVYnBSTeNJTT0PRObYrmOzwtabz3zzYIJkJqyy73F9c3UgTWejUZoyKHaQFcHyMa7ktxTj6/bcc
owsSm1LLrHh3eIFofny/JQFgc08hhoDjH4HBmTc+YHbequVAY6QvSkEm3GQ6UIvd1jOEfEvGW4ho
lmfSYygAnVfYhb/sDRW0oy5p2oWDbN/F69R4kuuhNDwN9pXhAeaWBQJyR/xyA3ZbOneq2JRsmwQV
zh860TJk+IyndqWR5PU9ju4THbUDjxcJq1lhsTPLOf6OEpTcZ+AMFLmORA==
`protect end_protected
