`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17984)
`protect data_block
85WqWAyW8JaHMWMkpeaAIfsS0tPN8YH0R7OD9xntrZsqBRUwp5QftwJ76Zr0bFWtL0zAQ1gtNc6B
NgKQt/vK5IP6b/8+7CHCrASINR/080iNW9AKoZbDZ/hWok1Ggj9rwW8s7QwLf+ToEixwHRkcj9du
DA8huKS7vRcVqkfjBmhPNbklrljFxe7yQH/EFF3Ye7OX4B6le/+eRJDHjoRCFVE7QWgVPPSj8dbS
muLpw+2/xSYBXDin7OzaACCmXZT4Hs04iU1gxuQ1QiL53JmeoNBOx7a+LTbvnM+S1n0Pf6wMd0B2
2JY8q6CYpwaYwpuz/53+uc9+Fa9mcx+JkJJckkZ4CpsUySyGRdAE+gwoK/dg7Eq95f3zjz/8XG7j
u5pysRMPH8yyp4idxBtzuD5IbAp+G8b3kGuDdQPVx4sMrp2juYpUg7bU/QZBWZm7+hsXPP3SObbk
cBE/HCjtbLNzADo/pdyWCZ9DdXho/xiA447IfloefFkLeaMkqYyzv9uDzyCQnCW1IkF+TthiTkY5
hd/44J54Etsn+oqj1KntM7gGBQx1v0S+GuDYSOtQemKvFYTCoBay2RcUtMc4rS/dzTkHNUpKEB4W
NmikgoszUHWqVXeQYjfVwxxStCkW8qJGgihOnHLu8hIKc2c5oD0s3s0rF+MBGV4MNRrpSBQgYTJo
1IV0fPJVxVtRh02/PC+A49c6JjRuVCcUKZ+TBRlIVAeTKRl3g+Z3ZdeFl/j5S25kx+50Fv5lzd44
UcALM65pa4P77q7/oGBPVnVIySx6Jlt5x70wsiqGb2koubZw5o1BgzWdiMBlzM6Xnc6KnfUYWAUt
YndB7wa9DBqDjaCWdxshiUII47yHI3Y2YV5u2DPwH1UkHbzZ52A1erQq96BE3c8JaWJLHfghwUsA
TDxCmTPjwdy62+puX1T3W8Aw8F4ejpBrzwSOZzVO6zztO2HGzw9ST8e7JIR7H6MnRbbN77C5uhBq
LhhmwcpyHNYBlEK6nDEXpp8a3gPVbC1D/a1t6FpM5GZ7qcexf51b3OWiCVpz3tEnb+f9d/E7Eoij
mdVmwFkMABJWUCZAEbQ0cUMv6Fd0ypcymOK/eGlxhuMHnsHx9LnQLpet3s+2MchHyIq67oVhZccu
+TDT9XxE+NVokAwlmi7Q4gui26HAdtMOqoMEY4uDukcTbI2qxfOCtZivXIhwR0RqZE6BcjbEnWvK
Zm8nzp7P7KCKRctaJQHv/aC8N2ljA2cv/8wHstOizWla7w/40ZfigjnrEhzxE0CRK8XQUpNrzvpH
/93aHxaRq++UUHt7kgqElLJI7IcujPUsyNJo8RbioueJzb86Du5Ej6eL9TlhTI2eLu3nLb/Dm2oB
v9LUNjQ7W4H67DWjMSk4Z7K3zp0K3HphRZXe6UavgBOmhhJoX7kXpFroGD0HZrMCHXV65uf9UWt7
Cwoya94k2/1ldG92DVpTYhUfd5xrH0f4MCuTLKxQzmCxmsXl9aW458/Lqka0nbMgVngp7/ztu8Iy
8/XTYPGIP1LkoHgEJy1a38fM3GQXjBfeKL431DpiAki1eSDN350KhojSh3NdfJxy30+htKWwnoAV
NBkgpuuUKQiTndJQD0OqtsRKgYxGxxtJhYA07fr/9jovQSNLU+x0bEkzEaKdcZc2nz3VwUR/k/Ye
W+rMr1pFyNmBbqYrHjWxVtQYigI1wN0QMYyFjcv1w4d8b4+jIt9LUUXZgtx5lIKh/1GKWNc+DZ3o
+4BsMkpDAodHvBgvi9m/0I/KybuixWXySbvD5Qgl/DVCckako1nJNqeTLvzI81G/ZDavAkzS7YZ4
ZZS+mhGscK4F4YWVHcm3kiM9Tmxb/+Q0mx1H4CeDzOU1rqtuIB9qQTBHSZr7LODJHyS8kj3sqeVf
WfIW2NHmzOh71dNuRmYN8AEuCfAx96Nvjqr5LSGCaGY0lBXUZVUNrxrCIVBx2QbkUj1LbSoGsdMr
Omvr585qSlCfu58BunQd1rbA1JVMkxD5NuslHEiacpQCRTAibZmHMZbNvraAO/zdZV+NWsRAzwzF
KgegNfUmZKMsTDmAPkOFmQTZChkOP/b3iKBfsHvJuSWvVa6bHhmdwfMMyzWvmCHmKSQAuLisKEi+
SQW92GxgP7qT15+FVUgkzM/TscQFE/qNQVzrPU5E3rERwni+pNcmwNvHXsfDb72sVkR2DN3/ZWUA
sNq/rWcOZ/HQPSnZjKX9MGp2P0x7F3u3Ct6P5blgb+14b7rnBFIiWozlwkFFCXVAG+6d6pV581Ku
zRGfF/oaLx2XYq5aesZVQeZj5OYgLiMSUzHde5+k4eDS00PSZDEOZN4+4669Wmi3iFc1hEjWzcq8
xSOeAbixbugccy2Cc9gHtOfJ0XHFj1uqyT4UeDdusS0BGFPqpBYm6Jj8RkZDiDFTmH+qrLICaECX
2nuLP4I8hGRzKKBZa93riHX3iL4Xi0KW94+SmPIDuDbvetVYP8V4m29sFY9QgO6q5HhyyEPAqpWB
pv0J38mXeL2/l9E73E+M9BbQalyXY3Tbsa75YFI+ccxPn1To9IhuM9F4q+MJLTGAJPsSiJudmNMJ
9CfRv+ruJGbslg8n8ff2pdzDdmmlDNE6Li6ATrUt/9TatFyyI10a6G7TyyrhzdWhuQo5C+7uEBvW
z+1EpLH45JUraX8sVGlsRH2JCv+2UoxlHkwOauUT/sERjtfFTFfnqgfECqWxyxtCzbk7gkWWaV3W
8asFbZYgLLAObtmcwvnKDRg7CbOL30znyqwcc9+e3jD7n+zr/OvZEQYKorHpM6GUt1SMZKw2kY/I
xJF5buYU2/JO8hYlfzCf0q7eHBZwui8dyYXcJn7nrqvnd4xabRQrAFUsnz2UuQawjiF1CtZxbYY3
0M7PAXxUK9EVKfet1b7DJj5CgADpuPB0BYdYCjHHVvA60wGFI/YQCe676nDq4nX8l6QypJDpBdWq
UuxXgQfgkZgMKnILGpuPxewCoMFd4joMfWDpbMemeXx511jDXMUzWXm4Hfn8cyXVFdFF5KDfPyiX
uymMw2eOrUfF2FyNQFfJGAxO549l3LmjKk5eiOnoLtwMCBd4a3MQ7t3tqG0eq6ukXdXog9JKMXHU
b2BXGK2ObcYK4DhA8X/ulOshSvPKaozKYZGxxVbkdawehtw1mlCzcHKHG44971cGQU7tXTXVrjuH
GdRzn+4E9Qhfpw1rP0lv5g9GeTl/visc12LDutlzn06+xZDGtpEJlIuuQiEHynzvoNhWkqDGrKbw
DAB5tknXXgMArSosXr9zIrtmm6TwjOX+Dq2W/ANBtt9wGeG8px/79xlGhMg5lKs7aCLGsm39puME
6R44ARwIY/ofowRC8ZBYbuOv6/7iV+MB/p+cqo0UyWGqRjBZaej4rCFs+C7S/+CjKu/GTied1j1T
9wJSioV8fExmm3Y1Bp7zvMKtmzECdDgYXVi2VeXNlWYItAD0vBtFBB5cr0Qq2WhK/4zP63pxTmQo
jISWyZqpspzRz08BtLcwaJn8lmVnTenJ7yup32UuJsMqna2aAHs6kVMc1DjgkVGi/xjWkPPUSObS
g+U/NFKUCi+x9kYkP3fa7IQ9XaerRKlsUbw09O3i1ySKJuHG1zdzbbxBWIcI8P7Be/3o0l519UlE
DzE8np6xx1a9+i+MXleX5k/QlNzAS5UCsC/ogM0mtpvayclfJeJRfVQeDMNszt9nBy0cdi4hmivj
n1f7nQSR3IXFnFwGTx9f2R8RNOl7WYyAGbIr5GsKDvIvV3WLdw7fgfxthXINkEc2+RFDubhgTHzS
RWkhxBgVs0344mQfYPpeeKGFkhFSHm1brPDBGM9YL822UHjKvbm3myUMfYaFsrKULtFA5cz85S8E
E+RrTcgNZoVr3lLUhvDbdxZk79LcybvjRKrl1LOgo/79pg/sXvgD3N9I+X12nkwnE9ufF0czl1Lo
7wZds6m3mt5mJnVcVgvekqOrHM+nt65CpgWvCYSs/MTXBDOrWZQ+Puo0PuptcJ9n2+3XvO1LWgT+
OZ6hwf9gqw4iW1UHx/OTRRVt4q9fqJE38pUaxdhatdSZBQCSNuWmpgIRDv0wu7cN9vaJhgWOoz31
rmPG6uH5xRUhKK+TVVHMQ1jv2MmIgj+K1Fw0at+gUbN7HXnINaGVQuWkvBYA5kPtndMUafv7EUq9
DXLqldn3yn4rVCv4jiuXTRd2IS5/+6tBC+r171eLCT09kxY+SRPP12v0MJ/6Ex9cgRM+j1qHIBMI
C2DFp1wMZkEUKFStMgkU+GXnYFfCkxP8RPaEaTlShbcPJ/fznXhOqK8QqacZbAMhiNQA98v0eNdp
fr90OgEL0aufff7QFOXzYt/HOvOcBdfCyqC64r0oyzFTWhuMzHav8eaU1tyzeQ3+PUNT6nxyXUZ2
TtaI9Zsojaws9TKVx1+0+LEwGzpmPlmcYGhTloaAgRkU/ZbrpwDgbeExePhxYk1lqBPmFizeNDht
msQ0aVFCPkQsvqNxbce95KqsvNN95LLBL+VPT3ux0MzTos4vJD2LwzzDQiozvrC1iWcXRFebXHJZ
LukhYDKP0W5ROvlQ1F+ipIqGEMxYi9klZnOEEsN0qpQ/fDjzSSFw+ifwSEK7RC2/0+de7rv5T9p1
S7/Q6R2Rb5/a3NmKmdx1ZuU2lakDCcT1UUs+BqEftdQNhiT/KW6c+K6IIk9buZjHSWwvdc3+UXFr
aiKTthFgRBDef2rKMFemzxHvHnVQy1CdR/TBfKkwOGI/MXzBZ3627JgYaEA98kChc83a5xZIdpRC
4TyN7CU7TzsNHu+j50/QLj7cS965obrduGbXtw/T3bmOzCp6lXWHU4XJwWN+T+igaMs6EdMJU1/3
Ctwkd0SnmmXEnTYa8Bt/bmKP1FF2KovQBLZZ2gBlUJWhicJyGPZNIFe2xZ4nvavuW3Ib1HxLbQRT
7S2kDWC5ZtZlteQxkR/pHr8lQPtqzLpD5ZoD7Q4U0BHQdqp8kDY+bV45FOnuynLAq1BcCbAZ46QY
srRmeRTVIO6YNkLO079qZUfA2qVhNbeTMvfBA9Qjz4w1A2JqsEoXvp35wolMPK70N0mz6F6OQBg3
V4u1KDBCpHz1LZy4yEg7CCheIw9lpXr2Uw8RVAqSBpba12L8/Lnu1sq2ZKXnGnkxTWi8sQDnzmYz
zZvz2qGkOrEDkJRlCIOgsV/SKD7TnDzajYCv3oudCbRg63HNEipjfYB5UA7art5TobQVp4yZ5tbp
d9BFamE6cVlzJ+beolfqINDWtY4fD2pP9GRI7K0+zaMjIXuYZ0crMeaCCSIAvTSle+lR31fJGPFI
mlUfgEwjIMlyCikVeQ6BqInvxJnAJiMCmtGqbiVqJ1VN83MrPKm+xMITUy51qQ9si+U8wUVqmZfm
wKK4tv4Wbnj5fJLlxb8F1jXnPq0aOJpTO5zkxUmRpWzzl8yFP2ldcejsdDpe4ORBGvj+Wj0d+Jje
Q/qbIS74Hs6qZgYYpg832xsJ5VjEBLJNRba/LUytDOBSdX2w6wueL4Zlk4W41k+FivJoqiE3eOfK
gp+MCMs8mc9uL6Aw/v/FrFplPjpx4bCI2q0F9eALLgO0+tL+8FsB6C+gpjZmKxrlJKHB3embE/ZZ
K6Eguxk3cpTkCLUGio2IGfy3PSdRdGVkGwhFtX+OvFScEUrlzUCkKvj/UH0gPhHYIUSZ/Bm8Wa/S
B/Y+Yg6/ZTOdnp+zq2jlvSLlxo9VPzemV5+lCbXZH1R7vTz/A13npe1yW2RTE4E06PV2jR9KPHOo
lz9I26ZyEhOOJUT/i7+hlEpoJMT1qA2TNZMuLedAJGgo+ZyxqrnerZzXOu2xm2g/APAm99WYh0lB
HUtFZFgvyJ//5CJC8Y+3V6T5AgtaUdMZ6Icfx3OY/w/A21GYgSzK95D1vz87LxtgkRPxN/qXZMlp
VkgXGH0nPl981UBnH6oloFVxqbuZnUG8J/rvXiWVY5CogMwAOnReECN0PbqRWn2Y+BWDvC6qh30K
XND4CE2Mn1Tz1UuFoDKvqe0p5ulko5/uDj5cbf8cClf0Dox3TEYbtX6cjwVR1brqRmmyeHB79+N7
bt6qNCoUwUvzy7fTLJVG6NEMirdsOkHfKvsp9EoyGmRV5NrddJmO+Vdc9aVyBTr8jos5crwlXdlI
fQYktiO+tipSJmwJVsmPEoM1el7MTC3ZTNaeF40eWOPDOPcX1Zsg46bb1leWyd7Rb47fV7/aMXQ+
Cb9GJPaLqF395P/RsLplx1jXmTFkd1xY5URJRUWMK2LNYP7Zm1Z91cacpNCD55VKjeLmgUJilODR
Q0//uz3/EchYikC3Ry692zVYwD2QAXq4dawxh0cX+GWj57oyewD+8SBoUTA7aP8v0t36HOu0aQcG
irCgCWhxIghqu7LD+q0Pe7JQ4SsR2VAP5B3roPEHAS7UeprEXcatkMR5WeCVN831L60XDFPmoCOa
KHG7XI0xFobIksY/e/7JbBSLWRboE0WvpEgxLkTfSgwkL1tJ/Gaa9xGSklbCefwmKv2nCKH6FlmO
gfdfsAKMy9eMfjvHiQKupSYMJtziL9+TlGKzSb4VPnh3NBJ3+VHjW5Syahxs36FXs+k9ZGDgb6KI
8WFDfjqDLWxSnbNHewYJDOOt2yo+nvLndPhTcicQ0ZGUbVccAk8g4yJiYyF9pqiWDjdg928QMlFy
SA2wBC7LBcdHvA8n44yGBSdZKuiVPnREnbZxLRu0YAVEvAfn/uAGtCuTrFNoDsvEh/srlYUGmDJE
et0iMlgzURdqoGJT4n6F3ug2/luTmzcelhy1SK11WXJ9yBYT1qKdAY8FxwQg4NFwxEhy57ShIhkt
SOnylG/nHtvqeLBq0AawjpVeOjjMerL1zKN+Kj3itA83wFhkKqtimb5gMCBjQ1AW/i2v2d2kney7
D/7NLTPAeH5aXAf3H1+/d9BIVQht7WvU30J8Avh4MzLnj4+D9yp12cuEfr9X3RIV8yztTVaYIkG9
dlYFMzPyhBAbAJ75QGNSdgl2rTG9DtNsC5Uv0R6c0LEJxdNA07mhG3P+pz1teaykM7hb/T5mYTIK
moqWkM0HEZNy4VYlaWMskz2Jvlf9V22Ri1NSeCAHGZuRYhDu0HHEObdPgojolpMnlqlS9vAvGsiT
VuQNx49kaVrcx18Qnxo/JfX3X5blzlDBMdVAWRcYX08v4Jq2nNz/EJfhOJExwGGGLfMPsWbZGzJQ
qQ6SMxaxL3dmNntoYFhch5Tt6RiR038AhJlljJemUIUd5XoM/iwE3C3S67XI8JCXndEFhwG0RcZw
/O/PmOCWbmY839PVkx32sHdwyWbFhjIGETnq/B6/lslnSQHpCIDXn3rkIF6z6UYUVe42pX6hokm3
poqL/3TdXorSHhIrlYEPp5DQ3i4rGC/+pauo3X8eOHCB8BTfVIGzYpRfxGkhB81pV+woiWrqxF/t
9I+Vll7KEV+/PjzhoaQbacznbUX4vbAVTkjFsHqjM+7FQNVm1om7iGdTv7Lbxkh3s57jAuzK4wto
Th6xzaSC+SHNJ1ORMSjaf7olYcFK/3VAvpSylsLTIGqKT5G74YFZv17+kZGy4CizzqQqGKfawyCy
yb0gPO26SdLoeI0fBgTeDQqAxm/7dYx/aWtYYZEslDOuCswGs+JN/imfv1GOJkG+zeiDu70xSwnu
3J1bN8s1pik+FB3ZIws8E6X2XkB8kxEd2Lz0kMD2uG1PnaPn6cfpJy7vG9OZ6lmoRWNQW8gc/Wew
H7Bny0HhR54v+TsqFk8hJdwq6zJ59NVWshh/fRG7FRtEqvViTVE5fa2tOuj6McO3ii7A2xJV6WXr
MRzt8CBJNmbUulnC87VETn79pgC/Kz7/y7bBQjf9Q3LOGizZSFknuN9JyLn3pdSZ9fCv1kdT4BNI
vXoomb/+vvHxcgck7x4PCiXGaz8nCgYjnMRncnR+r23mUWyrkCvcuTDg4xQhjIFl80OBuJ7/xy5q
1lL9vBRteZyCXA/KCqvEv/ert9gSsXrZ7TEkyQp2624Tf6Rvv0fWarO5AyFRUGwBEBl6GTy1HHrV
mQXVW1l7HHSQHQp/V6enHKT0L3XrW1ETnq0xY6R8LazJ8+57LlSZvdP8HFdEIQKWNyMPTlXejwy5
4iSChyeN7wzOxK3lzbXC4MKykL8CXFmXwVA24H0ajxXKO98WYPR43cAUesCBu0xPhk7C7Q240dNw
VQAdGqOqnWgb7z+zuc3S/WUSRopY4/xpF7/5IOrOpLduAjFmZ/thZm3WlG1w6RfN5E4dtvH5CJp5
veWgnXcshcqUGb4NfrbBpfvuPEvXNNnUfVh3IBCcGWgkmVNcr4udLrkaX80MEVnoz0Mzln1t20vT
pWnu6rIDpL3GhPIxOZ32JnNkgQYHU8w4FYDAeVaTXz742JTIrPqk18H4/IWLjQm+VSDXVIjOCbDU
RymfdgQCfVNi/eUZ1wOKwuDMmgpRtZmCsz1mIcwlA+nYLHsMdzeUZLuajDFJwd63qml5pPgb6ybo
qVkWP0gQ8wfxLq7aDcjsL3s72V+DbgTiSu1WP+iX/wfPNGBVYMgY6rd8MQRGbaSTUj9iV+fgDLGi
bWHfYvQM+jWbqz9NXoAghmwyvLpIKXU7vCROjpQJRkyRGuUTUwCRvzHPCQaysad/1PRn5V8JV4iP
tCk6LjVKn78vhhlM0XEmLvRbFbK/rFdStEBg20rXHRlFn+4jQzKTlhoxnVN34d4y8FkKeRjRwcqw
DFD4S5NNQfQQuiCoWF3hP+WFp2iiYArn1ix2Vgud0mXfgnZRuYB1d9qABCwq/R5NRIT1WMH8qK1T
VocSGvtQtaq6hlfCphgoOuMILDfDsi9/uTYf53tsKnbD+dXQ93PfwKt/PWeCU1niMLEmuIowSlhW
GDFsh8jp9Wc7N7d85PqJ/RBF3sve6rHs5KmvMzlWxU6M22zxpxUADcKP3CN39aFI/+DLsiu1+S8P
4SrYWCTHaxr9Q/QVhesxk+gNbdAqO8Xj7tCxa9r9xBsAGIZiJiD0v5Go3WVNkDlmCQOhwMMUaTkD
yuf9IX22d1UEgiwRCmjnCKQQWxr0VlqDwPjVrY26IrJ/rsFUeCMCLHTRSjLEE6GlklSi2ssGSUfw
R3z0Atpre8Z023q9bxe9ENi3oeH/yAq1k9FZ/oI+t4BMJcx82VvBVhWazaDl2VJprhnVHsKKvJBg
j0R8eaF9dqJvq1t5wwyB9Nb/tV2iTFCFKEdsp0rSuEZIsmwphqoyOcWf5Qr+WPFbgpx7LHh9b2NJ
0T5NIGHY60cSs9ZAy+ZQGAoX7pVGF6zDtvSUzf2jVIs2bNSF+4B6cNlmJ1mOl2k/a3gDxPXWtDV5
A5SRfgemieee56abdFkyC6PgxZbknh1HBxEqxZdzlrW7twuh70watnd9lQvtOpTFaFS4n3YM+llR
CR5v1UVxYncJFhv4ItoboY597XVSKLTO2ayajF6pUtzmFbIV8xe0sUuYf7pJM9kQOMQQ5oWhhqg3
ERj4fLZsmYHQgenlefMNlanDf+8az6ugN1SrCIczKkzBnikk26MGKh7d+a7SSinMY95ktCOzAq4L
mxYFa9B5tLmrlI2YBLY8KAXC2e4El8X66K9U1mMZIx26VoE/nwpuPV/obIeWZZ7LGIiwnhjkyCEc
3r9eJrPsaOf9ox8+GJA6GSI/7nlsgs0cXNi53NJVZlXSEv/ld736GhVTBXvomXnB6kcQkW4UOHXf
2+8c3t63WYbifTHWS5XpJNCkUd9pJSahTFQ7lhqdn7tTFClTZaSJjYkWfegRG2xbx0yY37aRkqxs
tk6mdWIOrP0Qkd6Hd0bdhGsGrMQ5J2WD3OO7LrV/MAA4ZAnivqE0/cxmDRhMcU+t4Ei48Ipecu5L
YKLaDjADMNHDLBohGtYI3InByIwO8aiNXYtzmxFc8+BUuUKcC5GnSC3NanNtr3a7912JKVH+CPOV
AxoKnZljt6600QguvVqrFPj5xI8g8cEyHv0RrZHfdJGC2du6dlNTfNcwjdeikgpryEqm6Z/eZ6i4
BM4bh+u0/S3lnUvNmpeS3tv4v5/ozTXIo1EyVsRWnerrzywdFBK/zGwI8nQ9fcno5BwY3r9Di8SO
4mo1EwwLdtlMOvLzlkzeWeI8Pz9NEQRr/agE4CvEzWaf+LNc6xSBHQA0P+26igD/g6ptlpMjS6NM
ouEB+chI72pOvh4MQAPtmodBbQFUU5Hsn1qVIvhS/R2yU7ZWE+2BxfPFC4jHxJqVEbEoS68ATs1O
UtWrs6zheVICZLrNc04zxlN5HMkY8mzKY+4ea2USV9OpCl8y/PizwiDbgu4mVmfMaJkH3j706PLy
XW6aPsmFbLpncWaLF3WVxbTbkhFCHv4snOgs/ynSZeOTpYmqZqsKikXMseUfskp8yIT5Fb6OItQL
+vnMQfdo6Ldx547qcveTBT96OQJmYs3bv2+AqBvUNM9MhKDpP4v5eynKepMMUUBzowleC1wfMJsz
y8mv117WYaSTvvTE4sU5XQPOyHS5Qc22ML65RR6r3ZUme2UHvuHWXAYsYeDD43uBuUGiYf4aqamC
xCJELrmBFVhq5k/CW+RtvEUR6mN9ljmClIh7XPcIfxIOsXoFfU0wUmWe0K+U/KIt1320Tm7ASF76
xTpB0Kzd0o1AqxoXl+f/mbBzwUH9gUuIa70RggLuOyxKutFYzr7rOtzDTpATMHABDvrig/aw8nUt
BQEYRcpAbOODthCL+nkXRzjZ6n2Er3Mu8+/Cd6R+0kpfcw2NGHONOssVEgdgPKd9M/nXJap5RcyS
SFXymzNy9fWVp2ymn8wiCBG2eOBLbC/aZTDpnXpw7htqNO7DntKdPA6yI9adUZwIpjzlshNfjeNa
pWs0CdUryzbWUp2GN9KMx8S1vnoj42C0xd7D2K1y1EGe8oh6Zk2s6ApzUVYMyZ6+L7BO0S6G99I4
zVLjzIEpffJaAaaCEtY2Y8dlqxK6B3Y42xzTv2ub5NbM1NJePb3iQ3Llp1qQ4H4WHzvDwMTXh1qH
/CmJXIpF2AsJMvmhocfsxHM6a13wdKjElY79uubx+bpfZOgqRCfNJm8iFhcbWWRaZ2zNCubZ8UTM
oj9qroi8igFnrPgmnM30/VynNpOzIsraj7uMw1vaakge3lY+lSgY3wUSQVTPdnZO1xNwZIf3Gbh5
rWXZcaAicD9DH6mZ9GnF6DemrgI1KsjFYhmGBylAGMNC18OwNREXraYh6X6TRbrzI9Ca2xiW4dOi
Xm0r6TOd+ePkPosEr/bzJK0O5fs9E3p9HXznQwahpOngDvdXTiv678CbB3p4V6/LqOPRYEiG8Nej
Z6bgTc2Xf/c7JGQFO86/tXAaqkT9ExDROwuaTwHf+5PjqeAqvoP50S8nv7vsy7Do2D9mhM9YP2uj
/4zou6vb9wEXnjTFIe/eOfuAxZqBhUZHNR63uUspSRl7RCE8lA9tG9qiRmi1gtiVE/E7aQZywSWL
+pUbV9xTQaExlyp0qrW7RWO6PeAUyqluUvnkVitfv6BHcgLc8T+IH6Wskzl2sMuhwQo+MaMkadrB
yUsERTE4TKTYt6DgmzF0XlB1EpS74yHA6xkAedymdHb3PRwPX9vXShSL32+wp7mv9WSfZii6Iqg3
ZAxJObwEgdeMfqu5/RKC/4LU2yuxOaFtk/zUA7sEEJsQwJ53/lkA4DghoMcGvjvVlTFHp77/lhDs
JqdIdw/gQI8hPtqZYhyS1LTvl/p44NusKQoWpLZEkODBb4BjeidqDNpYlVnQTzz0Jw5fAUshfkGZ
QbiTbsMONOTE4FbK6D14FdM2P3Ee73xlbjYwjXBg3sLGP+jSzTLlU8P/0PHX+Fmaw3va2nIrpMCZ
OLw26fy/yuBOT8hj8gFU7Is3Vcjv8b7RVvMSi6ZE1Sz+VS6163mr7Xyonyo7zrM8gJXUS7R7sqax
iMfpia8hk6cO+E0YooTJe+Bb3aMlCQd3EbFuS6DOYwBlPTlPtNJRUDqWGBPat6XMDmKIUm9yBltP
EoQPz6gSEWlmm/NsY5KG6iof8TQRxxhNlHyVR2X9TyTjJIs79D6gSxrIakOVWTUiLkRfh45YUyaj
Ztv6Ovl3k0ChsTfxHm4Mn3PCIqUdl1xFxJKPfzYlkfmBPEcs9LigjzlIfQQOlnHofIwViKWmowgB
ohjUXyit8S8Jl61YORlbCrhxdlSOoa9wfa7M5Zo3kpGC9otoFmLTMZhFf/gnvnGnks/XbKss6Ql5
7nSVC7/fdkuLJn0eJdME5mxQMmWAz4vjqEf046Zyy4ein3shMNZWB0jYQ9IrR00zFTtNHLBGPZow
CV8bFvwojn0KHwCMPTDerQ25tCUfsK6fIuUs2b+5oSiAVzkOb8edce/HHzRagDH5udw3LQKk7lk0
NxVyNXNvEdKpyMeuH86Ig4jenbJYlgLV+JkxfWNelV+AWbBHZKLKoOAoYsIylgPyrmsPq9qtBHSu
r/ypIucwG1/ANjnjx6WKuzLtEGxUFLP5c57Ju+M2iVczMD8FtEKq5JZBYrc7iEDyli4cun9PMTFz
U/DSnC1Da0coO8/udlIHi9bevOkGrDJuPiUBCMT5sCc5w4MdEAddzlXXqFwTZI9iTTtVuBeaIixF
9tnjQWcpM1OSO5DJIxR45pamuH1Rns44eYqo7bqeYgHbQSLK0dEQ19pGI9riGovIPVj3M24JvImR
3WChvP5n0nPNXsYlkOOf5IespIoc0OlfZ6k7xaTzt+QhiVCf6jwxEXk7Tti6c1DY+7Ne6WkShq2M
5VkOTRK1fnwZb/pP99PNIYOy1yMQBr+mA4Ig6xcEw+4j/7Cu3cnErH295TlEOwJquKPCVs3L50ew
fWHjilWMkidzl1lUxGJGO+BCT637yQwK2jaMi6MvBDMfpsVJnV1GXZrbb+vifsmpMuwgM3TOu0qI
tzIBR+Ltz1/u+Gykprn8wtPI3RewcEE0u3DMA98NxnmqQvoR9ywPczoMZrH6VW1bk1GIxTmLtJ3+
w8aJEaoLoSENOaBr7IbUfePXn+nXXemlzPtQRks0Tg8RTYmw6XgAj+mvm8j9MnfkdYAmFLofdmgL
NMBYM3Q1V4WUNZvOsBc9iDTNbWGcEG5bYFmYqck/NyO3P/2Jw/SPtbxJAQyVmc7ZFLLQ4qXX4JTi
uhYHEyaCTDGE46qQlVMwcmrD0rnSNn5sSswcHOJJsjyce9HZ8bTtPY32PvqrbtBsk6XnTjDlGK9b
8sR2vsvGyNj4JDlqXJFcpsK4rWeFazh2dBdLmeXkx2oujv+bX5SafkvviHJP0ZPVbw1lZM7woyEP
varpDwobGAqyWTWX5+52DaCfWdfzXQN5O+pQIj0YkT7eghIANGTfDRKoe/FX0b78hgu5exDdmTnb
YBW6GQ5+il0JJhck7ErhM/xi1gr6yr92XMCn6w/iNaYEnnULPMHUX07L/3/0A5ZzEIpMu7B60LBR
LrKcu2VAXbkgVn2UOsjMT3LaskPC5+D3wECSEYmlKRVwr28z74yvcDbiT0LBQBiP2sPZrbjmfRHH
HlojtQ2spew1r16o74RAL7buLljKNh+/JwEEZ9Ts9pWa2Dp5SU0dE3qzO16Rkl2nG/ezD3NEwdmK
BVvFGZC3YMeufxTklT3a5Aa2YXzlG9G38aKGyMHwAEk+gD8DBOIsNCjAYdTLCSaEtRocFCAndjym
nnhGyO/SoTDEjiFFNuFqitz3vSe89mrabD4sBEuL8N6pg34KL2707XkvS+fepbb5uvh6Ph0xC+Bj
Ae6Nl6Y7Pv/ihP+R+AvqqrYGzpylrMejFHtkH0pVXohxGxfDNLJKyZ2n+GdZs3FBSP0HPub+RXeu
KUNOE9ZzBiizWp+SUmFpo3GDsSZTrzBkfMoFGOoD82wzcJq2AYG8yUtxaAb7/nV++z0Ps8JVcylX
T4sSvbWz5p4653WOU7+uQiugXU85P9f+3YebmSWak63EMeWXwVvg8/+rlyXroFE3ASWof2KG7VZX
JL6ZlpxRSfLKadTr1fTlNNDmsJpgecvcrei+1jGInz10w6tVuq8jEom/lSMDfKbgGMLmpBqdb8v8
kjHvoLfOHB4a9ZwXyFpiPSO4HIS6xv00O5USZKueFDHJvSOgwfyXQ+MF1HhIHyI86AbZc+1IoROv
MjXb6Wmm0Fa8mmk/He3yI/KC6PeBGmCGPSTdOFYIsa4Mlr4YS9EQ1X0ORKxinLL/3ayjr6zhYzMx
ELlsTn7gWLeaAz6DRWSwHAnP5JQ37f1u5f8ZilD2eAcCDl0VCTFut6MsMCatnrmvmfoGVAvNBPWw
hE2g3QvpdtGzBrGMZ6zT7439xQYRhjX45I589BeASR8TWNB5u+mMJnP/gBHb8sdwfFt00qdIpYCD
+XsX14j9ws+Q2b9GvLuxnUYL/VoaxUP3y0k2hMGH0EdHwtoY1FUQ2FAjt5w31FvavI4MLTwgHaJz
XBIA7hCBbfyML/mc8WowY4+vGTmyXEAEEwrKgd1LeUHxYM9JMo7u9fYG/0kB+5KTtBCMD6INZMq/
30NdhJEJ4ZQpgDlpp2lXdh8I55M132609cHYvePc/H1fEmvQA1cJgQTJtIufTewMQXP7dmPc9MqC
uJwIIH1VnEbBbANJkOOJjCFJ9XuzHjV5eky6FGXjyJdmXDQU962BhZ69si/AJL80Jwx6n50LU/sb
AmGEbGtCAnssqcTLXOyqpDwYrddoCHVKfSeu1L55ccSlwfBxoXjo1LuRMXyqJwSyadVJHikJ9aWa
ypYcyuEs2rxqS5oMQNMqmVWoXP5tOhwj8mdkZ/Pt2Jwt9pI0r71lBXfTCIA1+ZN4gEdmXmSc+zcq
l/5Zh+yyCGCEvQR1QToDeBt8tG3iivkOee73qdBBP0KfyaxEWrFn/IlMtFPhFsiKbqOLBmMSwVDr
nziCrqK8+yXgSTyumSfpkjFj6glAJBCred91NailZAZdsIJL9OWOfqfp4DQQ0Yd/jtLM9A3G0wlo
UwtPxfxtCvQTg5/8/FWTticMuI5PfuaoLMT6sxOPRHm3mKOVRig5JVyPukBehh8WU1IfHy3ad6gO
sw6WSBSl3ztAh4cBnQmBcU3WcnhVk3wHRXmFCr2SZ7oPnMs9GvHAyUqmig7t8m/FOFNILLXSWUv1
LQXMxEpynyuJ5SZoHVkx1guKrDx9EWZXR1IU4yFil/tDUE8SRZaG84EMZPX1ktTpuejsQRIYAass
q88ckE7PJ7ZrFGHci/6kAyb5zbZ+TuuLYzMACB4XSbFk+QqpNFMQbgqd++Hw0Z1D8vA+neOEE1ao
Db+7ni4Psoauknr4iuLnq0yjlMpU1Xen1AU9xTDP/z5VI9SNzxm5hj0fWaidnQJ4ElT16L4jDuhc
OLwJe39+nXG+bBpOka83ix5Gn/NIphXkOAKws+GqW75nuInP1ru5ChNMHQeiHAntbLLfsphpJEs+
cSqXz2JDRe/zL1t3Orpi5Jhl1r30C5eBo+4AgYHJ9D8ROOzi+5OZlTK819jeka9Oo2KjPYbogxWQ
XwTai+12zj1jONU0/lQkYeWiFd50ScXN5unAzONT71BWHzJiwoFfXlXWDYl3sUGJIkiMB/Iea/K3
GIMQ93NhCY9yh3/WtS9ghqctKMurfVfBe1vrTJmmacw00B2MRExHcJTIG+nfjv6hLPJWAyPLfL4o
VMI2/fHsL97piuML65zne44vGmgHrD9eIKi4pEQMb2u1SouS1TBvN/iS5eC680A0mPU/T+KJJaZy
ffakcsFTOOToKWSf4anw6yFW50ZBgC186FU6LeGT70ITwIgbS/xXF3r+qj8/6ggWEtm6Qv3g9zzy
VImDac0e1U6DGQAdlu/1qd0lKoqOXg9cM9Xk74d3Q5qTK1bBHwQRzioa0R/ZFb0mNgSmgH7u1HAM
/6bMjGxKUmAFcYhka95L2AB0HQ1vR7LkTbVG4/oG8djg8lPg1OVkq/ZF/0kVmIav+3/JSV9YkGeV
mOJcMPH2eJra3/OKdr0mE/UsmKRnjTJrc5AWwJ6FUyg7hRhgzZuRxEWaGCOPAPmZIiq7bG5RiU+7
7Dlhbe+9/poaWlyqL1fFEMl7jRrtoFBA9QtNwJMqoiZgDtmDfSK19mxI/t37OSSfzJ/f+HKzK3w4
1fZL4QFiki6XN58GJLgVowezJhCHz3Bv4fk6d6HCUaGzYYwTGbywbjVgZDc7hgRicbY4x09b1Sss
woQ557/keC6xzyno8UgpqEXzDj335QJNMW7eepk7AihzDop91L4blNPRMyeHHcJUsCaayIFgNy27
iF2b2KeLxmEuMaThcIdltFMRCfO6Q9AcWmniPW8Qxl6FRJC2kGPkrOJOE791znEgVzaTo1y309aL
T5d6M9oXY8CGonISiMCgbiwQhgUhR7pvNYfqXQFyHkc53m6oe6iPPlvaSoAo5A+6xQ6Z3AzwABz3
/CxZ5QIL5HLnPtNcz/HS7rQEtsjEhEVrKUVh55BzoqerJG4+kTHlA2rd8OOIVF836+v7yAN0Xk9m
+imyWiebUJ7/EbZv8JBEHdyznVcTKbY6TDI5DDjFZq/bFugLWQF0Dlgza+z+AsRXltWH7u0MHQuS
XokhNNwEnEa9kQIl2ia6aPKKyC9tRmQIiAsUYzy2qZwOJnRhvPL5rXnSn4Pp/ZFhfIe6GDSRylLs
SZtQWeE1vhY1T517EmiimracRPhpjoKYIJM/o+l5IB7hdN2cl+KKmR1CkVVIBZOGuiMSg5zFe9T7
0OYczqlACsxSlmO5ZAYulwVNwyOJ30W11IMrbQFsCLKjPN3PKJ7e9+IFK64src5VCGoSpV4HSuZP
rqJ/fGkPN0rbinN/gSVv8plaHeKTk1friiGsBc+eMUrbHopnSovQ2CNqVg6R47ovJYcO1gKi7w1p
1M3SYPzaI6Y4gKUsHaKYo3PIDmegiAMI29uyAwuEQZn9sljVonDjKzQHpFlfy5DDyN8e9LGN8jT1
y+HH6J6UztfLmnAl7ptlyOV5Rd+6uDUur2al4amFOmqtMtEybkcCKgZVJyfaoGtXDCggEjCKLqox
zNhH/0AFpCWE47+WI8h8ubQT94rhp4GZcXqlDhlcdP3WkaPwJoMuttlvnKW6kD5yFFrYj1XSdxVY
t1/jfiA42V0cWl62q3+3+5rwg3XvKwhttqStQtqUadfVWuOg6qjQArmfzvvdupVXWCZEOKZfcn2F
sjd6MjhScxp4wKV6xtV+9jitGGzpZSdcO5uk7h53zS9Kd5zR8JB0gdHi5Jsn9NMZYYADoYt2Detm
V5cNaJ3DRxYLWicyohZ9f/VpZetTLrLajKxzPb/PwfNKVoTSpjkgTZ3i88ZG5oCF7ghthOFVRKTt
a18E4kel+yMHS3iabWelgODSRCiQxfGV2Y+wdoSlzs8iAi0dRIPNOCcZ3yovms9Wpu5/Rl5VHk58
oVNgyZutYDIMI0smZhW+1XyMypwXQTJZyIVYISmm7j8X+qX2Nrq4QJwgCHDItUPOYKR1BCv49Sey
9/fxez6jUR3bH2gEqy/NNDqRKrQ2QLigESKeCpAuTRbUdpYjDLqyt/qVjamMNbFURRxOdBlU23rL
ktJ5Od1tvA8zmdqPIDQt/VBvjg1bDv8yrw3sOQVLfw1cg0qUfjflFgp2GcSJZ7QkVccWD/xq3gCA
f1w6lbaKDp9UQP7ZeyevzlOlwVZuPQQDCaesr3fs1ajM8fQgxDrBEo8HHfutF5eu9glbPbF46SZ+
N1MvBTGuHI+Vv81IhYvcvKJtsYrSQ0RPrdf2eW0wH/Nt1ilMaoC38K6aVj97tAdqILmQbef6KHA3
MIjB5909D73VZQWkvx0HqLmZ1UOXP6cH6vysbeqtPAhJTzTY6TPWy5kDxETr2CjDHGAOgCkeZeSZ
He0AWqUDFVmtmstKLB8mr94tzvjEOclcaG64LMy5M12ifyCUejcJsgXlF0EUPwQ5rHBWGHpSpILU
kIFbyj5WxellYPMWulEM9lOcVtbKGAcYX5813PDkgscNLcjFb2RGWkf62MTqW++GIZT/4Mlkbh+u
jPxLT6ltDkiSWgjBnX8pyJ6mtaUEsYuYzsLH9qKEfSuII7koxhaP9PZjFU7B+eR62mTm2B74+k5J
ZoBhPzy9R0uhQh725AAABGKGjwTFTpGdy+4nBd1ui9Cdzb0Vw4qwEGJUEPXmhFPcf7Niae3P8/rD
G+HLYpXGNxecro9mIvgVnisSM7t63qR8Wm017dfkRPWYiGS3tF64oxcS9grNlEIpD9cSHUyssvwC
Gs2cOAV3zFXmHkBZnp7aCIf2mzNjdx7jK1ebQp16Ygqs0pze9cnV8dvwH2vk8iTq3PYyY3rRCAQh
X8MCSqtCv4HbcLwIjJdKQpJR/BAc/2nd5kxnBaFEvQ7M21r9hpqPolctBOtDU3WIsz++PFndVM/w
f1CyfmatHlf4mz58abWUcNGWGDb4BtigG51yMjCIFpG2YH5+uio59/pGG9ZceRCn1Y7B1djyEgPR
6RKNZc8+BJCvMkxMWWXOjj592B5jFIo+3pCXrp6xf5X6K9Ud02roP8G3JwXXmm/vULTyyBlc0pKk
LhJtjSpUMKshFc6zyEZjRXFOIDA56CKQArl1d3Sbm6FAoOieT2PacSVzco5fJmIMdNc9KKJm+z4R
E6KMkzxoFp7/jfAGERlSbI/ii5GVq+pE3TCEKTHU+O8GAC+yICWajR4t7lRXd72L5N7tQgPGyYb/
GsefEbaJvO0WzPkCQe4WjqAH4lCPvmOb6ddEFRSiGDmZ76wIujinxjrSXzgCs9ZaCqTqw1C+/e3J
MqZd+4pWenszVLbd3oGBGr1tsvZAOHkeZfX2xEldv/+Eq3R5Ropy+noaAhvGl8vscbCCr7iTKQXs
BaVwREsXv1xZZTZCXcGGsDK9GmuavO/NMN0RqQAQVuz+bSHm9ALT85xDhBvOIizLeAkyshSyaWk1
+a8GQscCqDpzp9WvYw1jfZZTI6D05h+81cq43BIqRZfT41tPYSs3d0G3ikF0Rr1YtlcsTryEEHPR
hH7ap6XYW4wV7aKJ33x5ogTUFRJnQjnWDi//Ic3u9LGfASghxJVdoFQn+8DpC/+1ebweiiys7BgW
45nwfLZzjVuW2DkEc1siB8flij84kE+oYYfKByuW1boYeTokl24hskyjDAo68nHM+PhQypSs5kGR
gYSVnAaZQAo2oA551iMnb4BfwngNNra8LToAty16bCEzviP4LFKarEBsndPFrsqWBLhQa9fclFfZ
U6vV3UwoaKJFkps+xa4rw2YPJmOEo1QN0TTX7b9pYI9SujAbWcs3QG01M498pNv39rPjEfQAp7ps
eA1DnxKLMblQDizQwJdDznxhFkx5cNAeNX4t2AyXaGoaHmdU5Lw4kSjsFcBXuJStKbBOEHTCrito
t7RtRpVL1uoZI1NS5SnUNAqiU866HS+/fAM/kRrIFVL+bZit6OOeEI12cMNvPVBO8erlSuZLEwIL
Ye6NiQ/gxzdABFSl2CdI+99lunLg/kTEnM0oK2OnQSKO9wYBHgq4ZQSQIIFKq1M4Ex5aNGkftWkV
aiGAbrQnhBCA085Pjo5+jx88Wc7+eCisbAjLAq1iGg8aSfzZ62+P/9NcYuGzIGqeC9tIBvNQcv/N
0k+9zRkG06NwTx5HcnaYP83X4klJFi2Mn2l4z6Mgpw1qrengx5VMMUpolWuS/EbtnZdAyEwzZYnB
/7rDPKsBgbaRmpfXFzu6rHWP7BU1fZwZZ2z7fVREtY9nZ33vlnKKTH/bpmLSN2f8qXZGtZ8j4MTa
4z+Ikmy772aOJon/Jgw2Dc5nR0J/PgUS/kGyAMtqyd4f6RginM/ke8vbf2KhShVPW0l9Gc0ncBG8
3VE+hrQ7LZpWL1tGI8VPX1g/CpyZVW+0BICOLr9PehxFBGLYn80vAn75Vk6UxmkNPYAQ4KF4JPwl
/R8YfCx2102k7K9RHBGfFbOubtwrsE35PySwh3AW8wt50VwnmvSBbtHw6Mrd7/u6Xxz4cPmVtrUr
wyhu3ohsrAnElKAV+kYt7wvHjG+tEllBOJZ7vOaHscn4xVTZbCfCRd85EK4TwXc2LawKoqWPQkNJ
64+UD9nm231mjW9uo/DjPj4//KP/6a3y1kOKasPw8YKinayC334El11FaDqQJJ2Uq6/5BOq1MSA1
vvQIsaJ8G1tZ1SGK9dn38AFxzeP3yX7zl8H6bE8cSOuw845zLGWyaSXgF9lPyhi9pzrMn8aNwXZ1
pboa3ZPiGssuIrpShpwsZDMTekko39JgB9QuVAq6+kC7XNtwFRny8jClZZnRSbQqypmNxdT3nnIf
aOGXaocz/q+bVxfiEnqqwuONKOtzvuVrQBDGo8BT5wrvZ7Gfq/6U5J1Q8Rsn5Rsia3w2VC4OHFWy
l5+L0EXEiT0yM5YuIzK+xBzOX1N4z/eZEvB5aQf1iaBoCeo8kWxXB+YSZBW/m99at5SFhSgmaOkL
jGF2nrHTuHzUDyybOBJAZOkKV5QyRL9ZvUuBrjkFgwiHwdyZjYAPigxzI5pAqTfDoUHqbkHjFVT+
vG3Kb7z4ZqqVhTsNKZkFgZmpXYG4/SY4tdXRofQjIjMryR5lTWXMeKMXk64szPUi+fKOWGiE72UU
0u/PrMVz+w4N0fj4CJoIwr8lfQ62GU72d4uej94fzPnVHmeTRn1aGmdyj863hT31ib6crNHggfiE
9flGcw+LETjrRUShtUhPhk/VoxrlzjZvbW3hqCna9FIzGlgnJycyn7wo8Zy4eTLW5tviwekdkmhw
S1IE8ITyQia2y+kK6JaNnrzC6bwX0vIJ5a9kfG6XwIYhapBWJLi3TexKCKjNo4jUNCaBkAGErSgS
lXngNlbD+34YHzv9CFn6it+bki8AlOhd9xbLcp+H5Gu1sa20OY2rAg0k4G5Hp5P9XvWg37jeGl3O
YxHfdEJGX5WFAY6kzk3KYOsWEqBKAqMHPzXVAIwkO9ykEfww1ENaN696skPg5ADcmFBXAqK77wpv
blRqawNCbARHU//gVT+/fCEuEu7m3RRdWjvf7HD2lsFwfmAySFjuhELp5N2BlRh9qj81o5etwvyp
LdIrUFtnuw6K20udmc+aX/rt9VidMfVNk40YBHN9ZzjoBHClgYx4NFuoA+Kd/ID6JvYqD/yKvpmI
h6L7wr+8c9Q+u1XBRzZ8nJUXItFJvxkO0BwQoBwAws8Ca/ChuVV6atA8g9oCS0IUo0HainKkPxXW
plNpV17mc4gmESnqHy4M7d+y2UFJHgudWKovZSHVSCbXl9KJYcnNCEZgi+9JwGw9knknXo7vnclA
BeieHtzfc/lfXIwCCIEHVhcjJeYCWmVsJmh6uz67QI8SU1L/Y5J4RpdVRkDapVzl+sB5AciwH6O1
kjA6a+Z5HAn+hQ+AYRnV0wp2E7q+GWczJNJVlw9v8bdnZCvq8jReiNhi/6alxHUt/bvZoRO4CGFk
4CQ47CkleXDV1MGxtyc51HSn4LOC8dkylzi7Q05yjl7S8zulNjPKud985MPz3CSOj72sQrgaFfHK
RjW9MTFENEe5U8iajStxIoFxFYY27FDREIu4YqEI7Mjz7Mgqt3J6LX2r/7qDuFfQSfkmQHIQ5eyV
tBonmWFXxyD8zSrozSpAws4EyKb7DwizSbqVRwICVivEiIYrbxW0Vb9oBRP2aynlUgQihu4fWRn8
KdCInNOStnklNOCI9qbJQvhULtP0/aAcUxKNfiUS/Qk347Yxx+Nw9u4r+CYRFaV/q5nIOTn8uEZZ
A+qkxcy9C2RI3rlWUX9rkbFbBsOVIAe2E+a7+FwduWZ1XU3eIo4+ddoCA2xEuLOFc1eC194IXPlv
rBnPgT4pqhthlQUi4XEzk8PPRysixsDegGasfEYhVRkM/IBDa5ypBFBrNsAq2qZJpaxsTL4vKyDm
SovplVo9Ytfj1ozB9BtzXZxE1QiXMrcd7G6YzM3rnP/KVglrL5hwMtQ2JpHeD6nzDuc1yBYATGyX
i1hUtvH1M2JX+CE2Gmkc8KuVxedRG2Pyu+nKBVTKyZ2ik/BonoIPvZr73iedWYrJ+gyzi6VCIw8t
ohRqADHy6DfxVeqUKQ2ikGGT/BAHv9ltzqg7bY2mK5vcFdMxQy4/sPvzUH+oS3UMnAM5LsyLs0cB
jPuuVGMMtCc/hFizibRUE42ngy1pUUyzKwnaH/fCm5XpZxjHL9PkSJ0HRc6m2mMcqPpGHjx8c0ll
C1G/m0bN/oUASHt2QTXVs3kLBg74By8bgjecOUtjW43iMcnIq/06364pYDLlkR7yyXi5gLKEs6XH
g4DyuJZQJngkEEnFRDuc6i6swvh5+dJ2qkvzU0SMm7K+9QLlKcp3W2dMC5jKFjB/81d9gWAiGAoP
djoYFVCxm7+O+diUesdKUrNNPlLl6wS9V1UDQqTdTMP8MgqdKv3GYLhImdlZn7nA83I2JDo6l/7O
c7Cb97f1IiOA7GTxjeH0Td8QGmQXdB3jXyWdqi7CLx21urB+L1yBEg07dfyoox/3Awlaww/OIZqE
VnPu91rZCCUjh7g4kUQvx9NowncJi6LbaPNb5hoLV4QdygPlPjwfu44GaKLWtFYHIWHZ8VSnRfqg
0xmmbDgH44BrUB73CcJKJpHWyRihwhfntUPQlTQ5fyrQj6oE3b4BqHXI959QbU/ZZfnkt9H4Envn
eUyI4bNVFOTCc32iiAC4G1+whfZCupXbXslGcnCc/azntMzdBAzeTo5x1cSL3OBfhNWAQxu3xONZ
jduoDnM3B++h8MnBt+nig4Hfwlg2OgBXp0dhFgG982qazlAEfK97OWq9iLZgmlEDkMH7nh9GeRFL
vde68ShGRyc83fUGubWDosa1EhloFV4f+x+a3yYTpTviImvK2lDT4h3r7xGrMRhmxAwwwfFV6mif
VNyws9P6EUL5d/oGX04bCg9WDgXD9grLvpZUjsmBTCbm0AibYNgpoL51T6s6WDj+hioLuipHC+xO
C2+0jSgMaKgLTHCj4GJOAtNg23ovXZk1m2Df9tuVkYC3zo0Hu/kLS/KbOu3KXDzOPJRZS9HKMsGX
53l//Z8zMEbQsY9DtrvKyXWlZtETwe2bFkM/l6dFzZg6u6aaMRyCahK9hhf3SF7QZWbYY6sBxhyE
OFs6xce3PJlLFbnEvS82Tfdh/DDDDvcMRZaN+IOX423icvPkKzyDZkVysPdxA/f3Rfa0t1OmN1e3
Dc2BtyMK2h4YmGE3N9LTZCx8XhCnDj7xAmJM1lky3FgCQLJM2nwNE7lzTS1Z79BAzjpggIS3jVNu
3HjIBHSa4MYTWHqJ2s032EnqsfE30MFHn4NdSmUK2dGWacjikAVbnm8ZpZyYWyECj1TKgAi+uXpX
wLsfXrsXlRavZ7lKhTdHZ7Ns6NDQyM0wPA6GL+wCvk11DA/ACDAikzjKHLsDeTYDXhkeGyZoOwSW
VQ66oR03IudLD8LTBj0BuJwVpi3/Wj9MjYDKApWG3D38gpHQp0WKxZW5C64KSrgi+1cTsOQOHDoN
GJ4OtDYM+bgJdUYFfeo4ZDrRxIJB4F5dgVs1GPUUapOjOEi+nHspghyV1YZl4MoH3vKA7haCtK/E
Rs9PAO82bOso9CFpzFrnj+TJO2N99t2s6zmeAlUSQzjEdZpmOPYbi5jRTr0bvTljZ99vexEfwdVp
IF/1Zjcy3VgJ6n3kXfSbHRoOO4drlmqCoK9+M5KM6q4+Y29eQr6CGzCt+lpOkUFAjCnRPUi58cvV
5HxeXmaYhtNZBXtkPQk3lmPYfNnjxKf853u9PWQ7gr61CjhNL2HfLeYY4yd+9Qf6+wMp+lrBYbH5
EkeiE4oINL1wv2nwSdx8PE02r/zcYaDCb2LPx1H1JzH3L0u792T5jKJlfmC1EiaCbpY36a/ggDmP
MKyC698XYd2x+OukALL+rgCBaDRdAKGd74vN2xqzvloziE0cQRm7W6o/Uvl6dYovRyxWvxde15Hs
EVcCWz8Put3meOop64STy5NZX4sdxG6aejvM1q0=
`protect end_protected
