`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17984)
`protect data_block
0USWSUGxovGsyBJteYpEoWIoafV9OFLI83TxNV1dwXPx22C3akmhPYESpUkJ26ebUJ7tLct96jvJ
0FbQNJDQv2THZw1cbWyLq0ITf2PGs9jqAFub9MYuH3cV1GQwmgzuDG/ieo6GTNmxrJ2iJdweFlMT
sHE1Ao2f7vfivzyAM+rtPlWPL4+zNqzAU/TMf5wJi52Kf5TDfqcCRAiQTr7x0QKQbzAev96BXTJd
7lFdOiRTDBG9XfD9qDyMYdI4zJ87KR3xeT/8AO3JvmbMIVDZSqytehUCnh4xrQD9H8spVuPkFMTc
d1ySWs5bOVrXvOy6976o1JD6kpSDPPoknIP909jIFl2g4tKUM39IPS6unTm6skGC52FNNa/iircl
m36uHTgUmyGxPk7YVG5USPfyL7LQ0BmilQ1al/JB57G4LXv/G+cqHZMwowKmfskeHSMKIjVUiFXQ
NtBrVBPhLLto3hKfd063Fe6thAydCbvhxRx+Hnd+9QU/TC6meg5RKohS6ySfbPnQelIEuVQeS98J
PYdVdKAV5ghBRcY88BtmlBpz3UJRut9GmnNmhI3koeOujUdhJDwQyATUd9HlA+Rk8myRXDyDGPGt
S5IxtfKRqBYxqCesjxTuksOOl8PoBXa/kbgNtjSkZ/tl8LZZCW9S0T9A2ovF14/BSbgXPKhLNaip
+sqdkEe5p3BlkSKXFO/7A551CSNFNfK63Uuv9jJpqsW5r5RPSI+UVm7zbzdJ9M6AvfarKcTXI7wA
j1vt3enFoEf0KEr8or/lAa4MtnYLiYBMNIBOiuHER9DWe3iUeFHohzFaCtmmopFI/irRmgISU6Ar
ATcYjhdqYvsM5O+g5IUKq8VZFBSuCZ6hBXjfzpVnsDoQS9TpYVRcMQlUK55On/faD/bF9dqCUZLU
zNBNn3+A8MqQRUNafGwgHNtm66EZ+6ZNgNTs/mLkO5ZbYouFCuhHwZm5jt4msNsQI03xg7vqS32g
QaxXkSVXhgc+QfXpkpwzUGT/VnZ/aHw/kErhEZx4fleMcoGS0V6GhqRzL1zxVV+4Pq90Vfbr2BN1
+wM1YQ+ttLICdCS6dfoz1r2BabsaUcJnA3TjGpRDIg/lbbWxJkToNvlpknT2cCYIv3NckakXcnkZ
GCxQFqXhQW3+7b6/98zkP0wme89A6GR+wlG1UbFgZVo7GH+0yZ8Y9DP4SFkQCUieOajji8xrUdDP
Nv6zcbjDmAnsR4BRVuo2uJScy7QxcqPuyrqtSVK27zPtL9UxYZa0G6jV8pP3stMK/HsCI/xfm/xi
9g86bVyXpoS68QGqgBm4ZpEEM67jFjU6Kr//bZnM5vAHuXnEqZtFCdO2mRD2ZEmm7Mxmkd2zCtDC
g6ttVz66+NkVY9WCkADmVBt4+/tTU1T0gt0mTTgzeFPdQpquH33J16mYSv2TtvO3mHqVC5iEMYDM
rE5iuIAbj9geVoxo5rU+C7a6YBdk18Z7DUN60mdOtletcAkKBxjFDQnXnVGOWw6q7l8pT7cF/NL9
tQKAfxh+c8zAD+jMFs4UE0s83s6tcRWUDTghgIa8Ht+IqUQtXtwdNjZk6uzQ3tFFUPUSU7+H/wbe
v36MHa/lHcHUpteSQsJD9KT52gO+zg70LT71DDrf5Omu/mylOqYbp2pwgIK+8G54arL62ncKHkOO
cEIFiL5rieKQjAt1dmInmeknwVl1LowTs5e2Xpy+c60if66KmrGhdfGrJk032h0FZG6/ySvEdrd9
2Z0dmbU6HutaeNhsb6dHK3EvXLfaVzKGsgqBIW4/0vdgNjng30jE5d8fOQXHz8Wdr2M+iv2oZ3/b
soMJ5xCLeyGf87Y52THd05uNIonIlaJnN3pseq//+5ftRtDG/g7Y7CVYKPqSZG2w5p28AMTni39j
vE80fK4x+kl/mhzIXqlJH26eJ1SnpvauvFuHP5Dt7cUcSD3tgz09hRVekm+30MClngsEtv4LZPpF
JYNRE8VjOaFu/3UdPFvHWjCS7g3BO1v1sIMCAEGbKNfej1c3S5SCri2WUN+k3Dyc1/3MxzVpEglK
LpmbfiOljbtgRPMt7HUVr66v14lUtW0JvnFFHxIQct+rdGH/to2YZ61r36+M+ky6dyvOkpRWqcH2
3gjMwDNLZ3oiRtk2I/wkUgS1V5bpsVr4GhnLakS7JECIb0hbYUcP/Yk3k+NJeoagp8AmVIUo3qJC
Y3Y2ped5qt3YHSQE+eQwtBA76uyDHqT3LPeZavL5EEf+ACUa0JY5x9MkRQbz/26UyIi1RFHbHVXZ
UYDIveM2MnJWdUO5AvZV02BBucMGjqe5bJg2A2xPU1gS4/x+Rb5AATxSUWe2BwVZwnnuNbl0Mz1W
l9gw1v5KR5Ht1e5k3X35piDIfWEVDXNoHzWnUfGfKIw5OLmOB1BlFkG5A0WUO5z2ha9qammPvFHw
Ga0/kAOJIZqWfnuAosbeZVG2QGrUp7tP90HKbWsUJ+9ykNGROuEZsSdAbSYRhFgQGfwJLxAUc2/b
d/75gx2XeiW6yxHQylwTRGgvvQYFtxOeb9tnLrnhfVbjpmNuC/ckV5J+x6BKKk3CdOwQ38h09ddO
RVoy3Sn5isO0hessvRWPiM+64Vpiki7BNuJUL/XRF4ddntVlymusvRuO1pQ3jC23WfrlS8xP20oe
zHjHXSjVejt58NnN+Sn91KpHvNEef4nMEPRD5L4IzTKDdH2+XdarE5Bmp55Bp5HPZZbTO9QMxVpg
OnyCYqhMHJvWKnkWS6cVnTAYN+UVRlDYF3xFnmIDaJvnd91kPL6tC0pogA2azqeuQ2k80upC76qB
YsSv0wgvDEIhIsAHN5cM4JHcBkJQFPvuBbjH8O34PATUAhiRF+XwUAIETFsIK+3991YCSIQkfYLs
rd81cWS3J3R/uJA5vt4nc3A6p9k3DEebthPE4vwQzrC/LFcwuBD48RPiAXjaE1ffZx5edr+krDri
HqUJzOipJbuZ43Ilqqgkes7oz/pdwiF28bfLI/lcAg1SlZZVzy8UESNBmDbYKQu1C22w0Qdf4SdF
cXeXjyHSsCWiroad5uDGIU/EDUC5Wf8XhYF7V2YsfPh8g54IJgmWUFhBAmQxWUDr1KOiknaYljyb
F4I5O8fUxYmkhFJRuUqNaJvf46SWhdbHACiieq1hcHYdmpb9N+/vZSoPJGzNft+JF0LqAf2lQ3NC
Xrv8tRcJFDtI4FDDOtsLvRSrphtqwrDzYAT1aBGY9uHy2OTDgVmEC1QDTzm3g7pJ2ToHiaVZcY0F
HFTaAYag8YTyaWlVGasXEOn0jwFJh7byMaL0LXecKnwa5w6PifsuGgU5wPFMh+rS62S3UtOgaI3f
pApceQkflja4ts5doXUY8l7FODlftBIW7R/PqdzF0qWxBFDHiRS/pA1o4qXyXrewIDmZuRZJH26d
xjdJtM6Y6S/eSR8ixEa3IBuWAUaN4kn4ZGmKgI5ahGAy048AdxJP2H1gMxztrpG1j1A17me7dmC4
IZIksEoBnJ72B1eKEs8me6eMZ4v21bb887DspnFqp44vEUD+8/GBjQrLpw9xc9yhDvvMahip3nE9
ikx1nDvyiCYCgjVwRgNtoh3a5Im6BCDNF+mHjnZIgHn9ETf/ycXTIYSOSOlcVcox1crnvulxNvuH
p2Kkr2TAIApQP7nVNPD5cmgUyJmqq9HWkKdtFP4oWJihWjw1/dxa22ioNOUjCAoMjziaDSeH+rCZ
CySz0jrHpgF7qFLQZWEhbiMcYUFXfhNHrB7BN1ll8QnylFh87t41op6p9cwYAy8mRwjNTGeaI7J+
qjGWkWcQUMYt1uDE3+MEGmblJebHIXlp5YRyvxJQYs/0VljlACbAicIaA7gavnFCXXba3jvJeUGu
o9Z862tst0CfzI0PqrTNgzyNVdTsZYURUqBcfNCFNAfhHG3LbIWkHglSchpak/A6AhVjsCNYX1W+
x0jalbNJVZ1uY7ftYCso9i9VrBAzy71xYJEMQV0lopia0155uYmGOFbLUnBknpEbS37MBwB2CbnF
6c3dTJnWkXfZUOevibUcdBsiYI7QbtqOWvGCovHTVmk8G49TP2YV0Uewi0bBpJQjZ6uTJLmxTGxm
rEHho6KJq0l3csWU+iwn8dL8AKhGYEc/TsH7nYi10AUfE7RMXIRG7cMwjJoacWCZokU7fu+ljN33
EIDRMPvv0cZ2ju0miWXwcFmHEl6a/luYhNDW42ic4SU5U9z8GB+ObhkX4rNPXTVWwFnPeSAi035m
MFK4zyOFVGkA3AFWGVcTJ5ofkxIOHXnYwYqbJ+ppduk/b0xV/eshl1Dl19yRDkrUI9RDcm/etJyf
uWMPssaACRC33rZKihuF2DGmCioNIMHqem+UyHEVxL7LLkiR7My0CYs9+eNZOeLbKhta34uI8QlK
qoew0XqwwBmHIgCTc6VqvNd5B5O19Gf2SWyAkvlGW6asnZMvgi7D8uEpAKgt5qNQQWKWbC70fXm3
C1i28nstVzxL8lE4oLjWyv7yn6GeLR+l1cF8QyV1sWGtPVt9AJwtJ+jE5sFkdihllnLNNwkDm9Ah
tB3HsqIvuWiLPw86ebm9mGj+hNS+4jt5v2ncB6DeSBc9aX/d43Y7OLwFDnSNB05PW7F96x4pDHlA
LaQna8W7QZNUuobLXAx7sIi+9+qEW/e36Rq2od/ICukq0sCbgqKI4VcIpufXvR38Ct2qKfO3r4t0
31KO2+TtHYapQFOAnB1LuSymomjhKl0VKtXt1qrQckb2PZLPkIOhBDwPSpIVGsKNhReupVkTa1Gl
aaYXqc2mtx6vpugJtxngZUvcdjp8i8Ta4LdvhISa7znhrqTmdGj5W+QbRcv/Ehb7hi9yi5enMlyU
n8QVbUfIxYloO9SvoMdcd+dXWAV2CWHpn46B5Lsw3aAYUmajJCOchmd3e/NU5r0qHmpiCcN2634O
2GzK8fnRuhwlMw3deQe8DE+zl4VPQfxY6csRy/qVmYIiCDVggHKV2ehy81HgjnmwWR3fpEHZAijq
ZxOXZeGCZ9hG5+q5Zm6yVHQZGCD1ZbJpEPmmt8tG487hjpt2/XKrq3zVgrCtYeDQVyAUQwAz2tBp
SawwJcRC65xZZQT8sBya2pRoE2h1kNoenUHVNceuCAxW3FR5HSrru2aQhlhcxaDjz2Ta7bk4ukFM
pe1t6y9bUSq8P9JalCIzcnlD6eOEeeOEFep4n2LWNFpRcQsulmbvCRmp3GDKA2H4TAyYhD5z+k9P
OMN/p9Bal8XRsD+GgFz93trwQ6Kq5lgjCuccvgxOComW0pTDfEiENzaFrZie9blJLA4QS1BdxuqO
iEcomdjK1D55hUY3KjJK6HxGEYgZDrJ+sZNcFLVqO8GvltNQq1706bq+fmBcgN4sN8Qq9iQ02Wrr
F0IbZ9+97tTzlHhKfz5wQr4yABqFT9KBHl/XBnVUJlIOMAIk8b6S55chiN8+2H06T+vJ9YddlWXV
zTUCANZH0OGOc1WD8QBCu4Y+V+WA59b22ln7ZIXlnFZoW4fXeJ9/NXJuUVWatX/ujA9js10W6/09
8fStVLC3TX0yR78WGhZIBWUUJi+fNF4nppYe5smg0pDgfG6bPCOPtXyeptRMltLKpGX+aN9fmNEw
K3DF086/Ujki3PZKpClc3GvKhUITFsUpLjzWK5oGwdSCVMd0b6US58802aDUVHKCHHfLNm8UEhrJ
ZZ4yIizgzDvPRdSnUxpSec8vDQxg83Z66oUv9dRh6Bs6RZY0BsaaPGHkxJztDsx4Etfb6fHH+LYj
IVs0mUtd9WxZhSfqQBm7rJYvSMcs6ltm+AVytr1SdoRisrW4qGsrsR27n7a8X5QvkHuvt74nD+8W
hK+ouq39EasjR3omH0aDBhnZ8Eqq1LT5OdQMRPRK0FYvYpK/yMkW/7iA3zIdcy+auS+H7Nfpy/p7
f9i6RCgNIlVMy3aVKTV5bOa7CQVLtVZO0xHzSnedNAL+0WerR0OcMCbcGjedyDd9F6YxHRGUFkPP
cdcRo+s9MMAp+KBVRSA/ZwNKWOr3kPb5pSsvJEo/tDW+HmjMa5tHVkK1iXlahlFHziYd3wXpphdP
lIfqVDEZK3eCElWMGpOslNGVKofvNxi84pJUJ17ztcij9G2ZCJPd6wOO4FKC/ApGhZwvImfE4tLB
qFV3bID2v0szNBsi84a1zG9dnFltAYvXZ3cRJGwbp89wTjyh1CIwA4YhlAGTy/fyzske7vw5TAK+
2ip7HpTldztVY59o6AG+hFIHlqppErO6Qawy2ODYQclwQ+KV/m8b/MSVbV3YjlKt+c0pEon6P2MW
2RXJaegLOkVPORN1IMnk5MLTW7a9CLTFYe7PGWpdiVg/mxiyBDs1pg351EiiGBhvqYoItQnhvmDW
4iEY/NtKCmzXm+25biFWQEyQIKiqx+zTewjEkWDK/Ub90Iu/b9WauQA/BydDcl5cmAdcCiWfQUDI
6ww67r6Pg0ANWkyV2jtmpSK435BcFkivl/fJt68r82LhelIcXvAEvQHiaMZdyESXb/p3QAwhU9ac
5WkoKZXWZMAtEaKuQzzqJCy3OY9bKniSF7iXRy4x22aslSnD+ccJQHP7s5+wJfj+abJtoL85C0fi
7u0N053MUQuHxlhV1x6MxGyRl+7f0ssgdnrnBJ0JlAs4sTRah2JCd35WvlOHb3sdVCBhEKXvlsHx
Q20P7ag5vF7Qko5riozEA2r8dGfffgBl1yWEvevGA++Wg+ixr8Is66+pzyRgRU5Aj/1UMeZHTdMS
/9hwu+o266pozdpQhuQ3XX+o9UVxTbkhpLlELpW07CGULugjSEh1ucnsTMnpI/JZp39RatqvtvEa
/TuDznp7K8gtJX60QSlsSI/m10B0leaaQy5UKEj8WkAOHHNoUryGvebZ2fZIjT8CujPquOcfGGsz
Sjx845w1eX4X0MOA7wk6uizFaxiZknLG0uCY6rDtXp0Y+yvx1m1QsSej0pgzXRuZxDXvxOMvDPNM
4QnC5KeYbJp7Tz2FR8YavmNDZNJtXFp5gNAUDbjSr2xcjzNCT35FFK6ySV90A6Oa8D80PUw3Asbp
FDAKj82js2JTHuo6n8LtV5MGOV/RWr//jvAGDW0BFrr9LqQv/NxymXC8TnjIG4XH0bbrocPadi4O
ygRK2TcbS0TGaDJxbwHxsLYrMeLPEeRtupRlkcQxHLopJSzwmK30HxdOOZ8G6tpiRJgHDnfZz6rz
Ty2pLx7z2Tnjw07QpUk7d1W4429oo7NzhNil3O83f6/KcNd0o2v3zvXsHVOw0GmtrIfDxQDqJYIJ
fhrN6Q0g4WrR3fy1ZqV4PEUYHtZzoESfyMqsaQDS++C3lNieY/rkZ9mzt3NantksFdxpQ4fIPC42
NygcH60mouo/ff6lbV6dyLP2ZhhfznH/h5zdGkSm6WpUdsiTUmBiGHz6FDAXKSzbPfRfN5Nx34Bv
ZPuwUD/FjJN+4pxuaMC+9i+LtYYUPfeIjxQoIUxnMKU2WBcMsTmNUivPjr+55O/MiQTEzN01iCch
XPXEG787Lp4R9rooFDkfyKXSw74mP2zPp3upJmQ6scDR9Hi3qNzS+SDR5DjRaNsrb8Hua36+7Q+h
qOguyZr0oicaml22Fp5jn95u+lUVlIS+Q/wFFnI9mZxNfN/pt+1MEtixm/iJ6tx/nBsdbVcqAdHc
2tOlRa5/SFcIhGte/SSevznC38or0fddt4T9kKy1DgSyegS5kogLpFgVjkx3Tvr120PqnevP7MKC
/Vtdvf426HhOiJSQ/c+qfYH5FUbeuFe9CR+w6qqibIlOFa1Pt9BG4F6IDkcbqe1AZSYFJlTJy0wY
nj45fcUeXxDf5VTX6RGYnF58wEC5Nl9P/pYufIyGzUs56c7Y5YkIq1otrClMThtEXmCreTisGqYJ
KUQ9Onmzb6QkVWN/T/uZpxoqkB2Xi41k0aQ+V4H4nC0lQvG/TcbRGy2CsIp7Ypl/jczbtqcn9cZm
fkPn852EGeap+Mf7qw9sZ+Sz5udSm7UUHnLxdnkn/w6jSBVxoquCuLONcb+NFuz4pBJynsM7HizI
0dheEpE4OkEnPVqST2Cwk4fcuCyWAp27xZ158+zUd/zxjjKQs8JVMh9b/10oo0I1sZq54rOTSxb8
eKeLKZ4BaGa7a4BuZzvbEikXAHqt+U+UTJ7e85TV3icYJXXCAWwJ3+QxI2H1priz0pP1V4AJiSE/
0Pjxi4yM0bclmTVgRsw+kg1N8vJERMQ/siIQuws0B11Xdb2L8twBpybS8km4agamLKmWsjqQrXUP
0ATdYBd0R3cmfYMAW4X/QiXepzEzsYV1U9HrtrF+IwSpnBRbpTVE+4DP7btuySReblfFkv9ZLS3U
R+ExWUaIWJHecrn/lSMmi9nEM8r8025NSa+pQ0ljfJys5OMJNg/31TyBOum6lBeADEGzWctL8Jmr
tRtzKH4vBMC8mnTwbd7Avy5rHnPIiwhEjjvbOzQ/VlWvncFP60TlODxqMF20P5TDPqj6ZIbI+Qhk
Mc/dovO90/2K5XILzYTNH4blFmUfzZDUq2v16pDoC4rEa5j24at/JLAZs4R7ux8aJ4L8aF1HSGH5
2Fj1vSNJu758S1zpH9s6ZTw3zHrC7nxjSwCNPeDE0m23PkM418CC58NQZBpw3SvfpVZaITzesL5P
Q2Z3Q5Z815kv2myglu+rlveeZlWsoTNQypQCp5CYx+Ykwobwc3gTrUPzRnU/lgvdooypdfdYddHD
45eY8TNpRvuUgKU5PCzN44q6wAfEeI5nMBInPucngjKzFLqsBBtzvNAOZI01SIpp3yOJvpIJy2Ot
swf8IuG2rgvgnL37NH7iJBFUgyEcoHsweJvwT+Oj8kesZhp3RvpkqCMUejMuD1rhQWDVZoCcKtzB
2j8sve52qZOSmGqad0Ffi4tzC6EWCNNEpT4+6Bc6y0qmS09hTo9Chw4wYBlrSHSKP5WIuOZvZ3Ks
2c94g2DKtOt2yqePIDX5NLmtO5jF09sFY/tXAJ/mMi0f0pXNFpchw9h9joU4n868VhSenfbw1Enc
1JTtL+JfZiTCZNVzCbf/rcyHB5qBUFfMLU+/Vs6iykc1K4Oyu8JR2og6yQWPT6Z1Jo7e88GG4FUt
hV/ML+kQlJ2l1Us6iSEY/OamXm7TWdyQm04+aemr0sDDqHRIK9l81CASWX59YtUs9EfAvpmRVdsv
ZD2WzMiZeZM6A03cEYTOENpnFi4Zl/qxZLg4RRuqtHa6GtzdTCbKXcUmqoBSZNEIiRE+kS/U5uZD
mwSNrZKDf0NrF6mEIiP+AFkULiLPvWThai5InuAhJQmNCaej5di9+5EIQ9+FSR5r6UZRJ29jvezE
7xsqlbUFcWI0+N2HVxGWWtBNrjR6UgfptYR2Lkft5w93va7tJvNTf6SEVCZbM12ECDBkg4co8DCY
EBv9oCQHhc0qNqyUfWrU+GC2tXnCAUZk8mQo+UQthEUm93ALvYw0r5X9lwELUJ59in0Q2t0EFecQ
DBI8k/QOtqf1yF74sjeDe6nAQWIE9wVEb8Hn+b9yeha3QfF0Q1Ut47LFt52pfsEmmg/AU3lilD13
4q9CBr8hB9/2gfom2GPxDfKzL8bmKNjiy/2BlDBQVatjSiBpHS2ssajeSZCdQgCjXHVelsqpDFhk
JGum+hQxNzCI6HpECYFqGbDC8c3LDPcEGn+qDIIiooGs+KWpx1KMpIwWdzVAg8SIYD+IytyAPeAI
UvYFIiTZJ2kHkIBtUAGgnF286FvRrGaVn6/wk+5hs9Jzx3CQ23ZkfCg44BFYBpzCtoGxpEhvxTCl
QHQSe/2620TpwPmQHgElkx/2Gw/R7mXHe8dO0VpgM3ibl8ds4R8u8pkUgFD75Ioh/wd3FQ3to1/Z
ADALSYQR9R1wBfcJN2wrM+QiSrWpgNoA8NBKftYvErnfFWeoynTH+AdztgTQS47mrhKT4LBeCzPI
BlLD79Hu0h5K7EKUThJWQpHoCqTyIIMLmqf3w9yDT5jH5EfbjvewXimuwxHC3C/W6ht93otQNnBM
P1gFMwOptAxh3VOi9ktuJ4IYaGHZbSwtJ4x24kRYIkYZLPDwjsah/+/9hcjIgAsKL5VIjQ8REeal
R35TLT3v2QbFoNkF06eT43semI5S2wn2++I2unSrYdcFGpdf5zpVjP8qwFzG01UIjE4m60IMQHt/
LTIJfVli34b/a0+cjhmVfgOVuryfxYW+sVP3AnpMUFbW7XW3m/EDXsxUou1bbr7bhxQsI6UKRdM1
a/Cf4Cv2diJiCxLoUPETnTR0PfTeohyKk+EI47jtHRP4ybOwpVHOqdFQyWll/D0SOWMQbIvfOQJG
rqjOgBKP010fX1UqJPa68By/qpQd52lRV4kym/fP6+duGEd6Zp5t42oy0apeUdMNL65kQe/21gA4
7p0cfVTPyacIa77y0FqkX5qRg6hXGyP3bFn7TVqsGzF+SlcowGq6TyOqZ7Zh4PJi0M4kPuKZZpcs
JbyJ+Y4rsX1HXBoTgRAllcUil6zi40z4kHYqrUgnZZ/v33XDrjGhcX/ELjboXv+hlyxEgFZXReKJ
5NCWOQeDhfm2fsX69+8jRT34SJQlgz5FLl2qXzWDW0fSaPItZNpkpYSm7+jXZWUG3YDt2RJoE/YL
rv//9LMtA1cF4ZdjAt2u1nj7SnESLYTQZx8A6vY1G6i+zDtMjrpuGttb7fwuSML3cMiXtiRhoGBE
VeJqv2zWjTR8PtGDDhGHOiQ7D5RLWkxebCkty06q5rFJ/8nSRo+Isjjj/JYuigLwj1oZA1IulYP/
6nYNJv0tWSNU/78IWueEKrpKbOeDl30bHtEse2KVnFLNEej5TASLqwKsQf8OFn4E86zzhotDUhC9
ClH2AtFNmUC1iLQIFmlWSHueEoJXkisuts2uCXttGJsb8xHiXxpAZpI+hv3nIpcss7pctSo+2Azp
LsmNwuAJvclBKaLMVz8pcuZf3VKtHFWwc1zly0ttCjQzfZyrHHrCzFV4QJtibMsYA+G98KqBqKOL
H6GwMSbO8r8gH6/Yebhu0BzEyTJ1hyVfpPvID6QaGU6n3DsUsZc8+oN6sbAn0/lIwB0xEusiBCrb
IySPKx+6cyM+azhkEfMisgMDfaBefs42ukuD0jy1hCZlxjo3yfa9RbBYsrk9UyFRz0XkIZIgi1h3
BWMMK0gXdQhGEze6elfxOGwrfdQ35XstVkUz7a4GTUDRAXppiR0SqkxIGy6OvZoycBA4zYNh0Qq2
nP3thBf2oNBjluUnB/2yB+b5BlWzNDFues5qKd87GaMHhgwez5bayD0YxJfF4rLpa/ZIZPnWI+z9
KBZGrfET9GUuG7aWQsTradu4b4hkjTFWe5rADjHxYl4ly2Y1spuGfbyysDqoOnRb8wTfR97pUsUs
jR/44Rwr1T/AkOP8nqOw2zibDGtdMCdjAsgVyDzM6w4z7+pWowwiS7wE6UWKmpDR5kx5Wvasy3D+
fn7gMqSUxIo1AZkoj5NFR8at+8ELLLPu3fcq8Lfwk+OxHIHvyzYqeFiuRiGh19byc3Ljsu1y3as8
+OjHBrAWu1C2esjuwSLit1/7YZbc7bq6dqo0tcSIKPNkcvip/Ht92Mo4NeMvibWpOjB13RptcCCr
1vnVVow+/00iTf9wQPAaBgJC8hwVNQwI5nantwizlWN0kGyBLNk9YbB+/uln+0ZK1Yz8x5eiHCRL
JePGQ+GltL+xdZEyhqMA82Qb+tuJpkz6aaq3Wk/o/eQ6uz+dIlK1UEx3J1gDqGbnZnwziC9zHJUL
XD/SX9fXIzoi1BlT+PkjuyGtkNSN00v3Gn+q+87OItXTBmZN6+TQRQMV6tVpP6cTVNX8bRd7uiH7
rdXYtYPvny2vQNSt0QX3x4kRi167B3gWqpW8K7/RFTmM+J6ha6z+6JwwZdhVuEB++vUTYkWd36rO
TPNdDtMf8ReSNNe6Zg5WCUytyPSuZw7jS62NQzqW96Ba79WNA0fV9A3WavVgaAd6conr111iG/40
BYV0EPiuqI8j+a6/WdVW4QnsjjH4rxhN/9niakO8P5/EZnuaMp2S3yQ61//E+dk8TGcFAFls0D8M
LGZ1sviRTG6zU4y/GFF/6Rx60Io4Wx3dsV7zNBphNw5fLMKZ4U9rPmmf69xXIvBkWH46tiQK1i6L
S6csMewXSV/Z/1lHXMO8heMHPjI1jdWD0Q5G7iHz7HRpCmG0q5PyQw8isnNIZx1H9NelLLy1pamu
NdB3lGMFL/7YAM62pJ98/axteS9GJvVvIrVqdlZK0h4OFg44mp5nKFAx5m752MPCQ3JfI1OEQbsp
x8BAKkWKQ3l2FQQhLEkSzzP3NVjpDjygz/UcUbf7ByrPJaqJrIYPD66qljU8ZYztbe64ggs7oRa7
opH/wiOn9EghsjpUJKgsghohXFq4jvKJuZyGkpDPt5kHuQlQuWS7FbMlI1yiH+tXMMB3ImjJc9v7
mhA9Wgeik1Zrb4klP9kCzc0p3gqFzqL1G9IroSVirwOzUGZsgQdz4wfK3edFWWovik7pHHs6Xygk
JlN0CRpzZK8AUbQBQYMTqXmFMdLv28mZOLFT0cnueTTvUtWenariQRRK33xTe74yXxVQd0ch966O
1BJBm8z9AcsjMwR+sne3JVelG5tZ34BbVZnItkN1UK/mYcL4QCZZGY9GZPH/iLLeoXzrHzJZb0mm
20LnEvJocFg0wS2/XDwT2GA2vpdLnB4oGlvNXYG4vZZMvqrz+UGz2SQiLV/sIaSG39yhQtd6Oodn
BXGyvvSKNk3O9DqU3eYsthaj23RSdzhpQ7m3QTkycpcVlIuWceAYHdqSAW0SBlsjL+twR2980sJR
RErQqqU6OddFRG8URYLPMoc1ItbyyROcKptmDx5kK6PqYQKNt9LRDSXdA3eTaZIELMPccONpWRY8
YZGh9os8M12nP3c3V/Gp8CFGrz70yfuOwIkA0lEcBqEMw9GF1l7AqJxTxw9ipRv4AbCRw/I9jea7
ExXiYTF+uX0tZAjgP81Ss3YsCV+yPYdXnML1aL1hqaVuHW/ZLKFRGyPMtL89Ln4XPiZLuhaS9Ek3
xoGHTTSeFVv3o8qhCJxDrYyRF0AKzgiLZRO+h9i/nHaltxd3cev/h0HEyiwaU3HE6zFFk9WVFmEN
8LA1yRben1LcNcIR1NdCo337w7EzzOUJnw58kZzphBYHuFp4bHQ1cWO9H4UuM0E1TVHDQGVnBMUD
0cwPJFfrXRUSmGR+7+oTqbULUD4fgw0Un4kz2eGKAD+FMHD3VF0uFDcFDWjIz7iad3VjMp/gIcIL
eVWAK/WDWFukFKHtHyWOgMLdu7DeAusLliYvoaJvEy/RMe3hwj2Riran5tHjmFN1mKdVRGlQb0Sw
OfaHYiapiBXDbZfjzdn/b2fbfgDl1z8e0vMJR4M8XYE7Yt6lin5YprfslGgP0sjLLDv6PwgtYV95
FlwQlAMYFpNbMorGIAyyC7tGkT3p/QAsCs2G86/VstBTJOztMPlnTD4j/+ruO4963m2sjV27NMZN
C90YqgTRd935vg3uxD0e4WzkIxtkUIp2v+cRUj219nX3Uj+Rr3z2dCrEFQVW4SZveYPBKjm+CiPR
VA11GgIy4b/wQfyUPIsqmTi/zaDgvgVNR3NdKED02ximxcUAZZGo2aM1RdsOoclC7OJhE0tY1fIx
KSWT8M9BPLykCIa0lNU8g8B/WGi0rC8FYNQqceBCMBaczaYAKlm6e7xwT8WFmJDyGz8769y+pV8+
/kKuoIcVnnN83DEbq2EXsgtEVN60qdutR+3usDqJAjf6WOJdx+nSfMTPlh6E9Yox8g0BR2NMznEQ
hsioJ0pSWqGsBxiW3kNo1pfQykSF8JHwijmvVu1nL68ECij3qK6cEtLlSIRW7jIcV2rZ0Kt6jpwJ
aRaGOC80JaLUhU6ms6xrtBD5Bl7RtYcfS0IZ//cQPO0wA//GVeSM13YDvrX03ndWKrdccF0dEG84
YZ218uWjOw0Ry0De85e/CvgEPKpmsY2srtwBp/2tBppfMKNc/Oe86B6KKSMx5ll8iopum6qo4trx
6ffhdLlZMsg8TvxsV3muktR5ZcqZIxySR97ZNRXI1RTzRqYO8OdUbQgYM8X/U7ejqpjMpK16cOY0
zGblU808nmPpQhtfXnJvsa9dWvHJQVbpW6GB5Zc4tr77F3hZIX2aKWe4as3MdXPN2U6U2HXF9Dzt
roJjJOaZYDcg9OOz6nDIlgtEuMQGOmompdghWqaRJGBaiJxqEmLG8zAwZ9aR2/GKSKiMKIH0n0x5
bdgCtSEWmjDDGaEpf2BQYxtCWZcjm+fk5FLJ04ohh7FE0db8jdhk/Hi9u4mj5C2aQA5teftf4LqQ
YlxZnyO3XrOOYMcGFT26qhoQes4Iq5HgLe7OYIK6j56c0w9GmMdV1XdRZ/D7BJBr7W+bjO/Ncas3
R45fZrVhe18uo+ekuZAIkWro19Cf8BTX544ByD+jzp4ERx05BiIT/mxXg1ZZ4tQ2R+91Gj33sBvH
7kVSJ+pERd/PrmJwxoauqLvn5pxSfu9pj+Ca7jcaHBWEDLKcyCFaZpJNYu0uAtLXpHN1J0ItDtRd
ahrbBG9OKdQtKZs0xxFhtJzckBlHTM4hItnuY/C7EOjdzLgTD/sp1KXpKLwI4bguuGIl2D9IfKk+
J48sg9ARrYA1Iqh+ZOxLXz6eDbZ9Elqc5KqDbKacE4GTQJAEIaAa9wBO1uran7GpFpcVuC+WQtue
+HZD8/o8k+EiigAYVUTUH5lEbE8amYW3hcVSob+73nRowuHdML0UhBRqaXBz48Agy+rygz8lk6zc
0C1s32SOIdrKQgbqfGdXr5Jz5teN9A8cnWKYVn6uRdwVEGYrSSFJ0uwiXWnHHcUeHzFsZ0smWFcH
g8qkME+pufVwAR5Ee0hNyk6ro/8S1pDbcV6cFvrE3FYtkRK0nKlAW4080UTKr7mcXcnlEg7rr8ch
WgBiJrsffTpj3Gpdv7hmFhmTymi16poIPvwLDqjVqhl+0SYmnbSMpm1aEz7HmuOx/peekoCYkoMz
IWSE8Jm2zikuYgp/Yv5piKhdKJ/bM7nAsqJuSZg3Vcn43T5LMV8VoNR1O1GQbMy6DjYQBKd5Ou3/
uetB2yGR30Sm5YSnIO35tW4JXEIG74am5y5Osar2XSiQO6WszYlTeub+d1b66nCe5uU5q6zI643C
uaPIZu5YGFIbezMJ52GiaUstn/Gwe2zbO2dCaw63GXdyhxtdQfHdiyVOr0gGLo4Zc+HNgpkn5Nfa
EeQ/NWM2hYgaMnJV5Z2Y17kDRj6if4A1tw2iHj7vyQJp2UwfeRXR004cknLQk0OBVD+7pjJ6fESa
xfmqzIXtEo6smpn/q2gWQq6EEXhwN7TkRHLNi/a/3T+iJt5KuI6lw89OOk7YDYu1NDCDDL1r4vxi
u56UUOlEBEAOsCqqoR/I9rQAKJVoxdPLpGK7CtEIydbk+OL+vNzDoSVuKOgt2A8Is1TszGEaBttj
XHPv+9dXSly6/5InwubVF6PsPm90AeCcQv/vrshRIfWurGQ6OPg4VW4UeOvM7AS3ZaiiTwNPEzMs
ybpbRUUtAOWRUjTS2kTDDQo7flXR3+eqQqqsB4sdfrDJH19Jo8hgCrDODtOU+ghkhm2xb5Y/qAtZ
B5VEB13huXrDl5VNRVjH6ZNIJmeR2t37ga+QgvnndTC2NuUbLAodqd+KMLh0ciWVevCoyrAy03gP
Sju+D0vdk+FVRZYKR+5VRZ6hULyF9S04uzizHlsQCuqe47hf6zWPItmzSwmSeCpw7wmIcpMbScQr
FOmm2Q7PIW0wXmuKwBSyDfQiZfpCbC3GIReTlCpM/xxdx5hfAQq2tDJuWRsJF8liuMZalnBy//u0
G4iWkxWGyILKMVj0UEinS368HiM9azQ0DS4OBoBpDs3rikQiUEQYj+uq/Iq7A20x0t05c2ipgfMf
vOanbUzPBFYXSylD8ccO8/xQGR/kj1iZQadgQ1yfn1tEHheq5AR0/Cn/OIxHVkna0hH7Lqz8Z94y
O1Sluh6XaZHbMc2jkPkwyk5A9xMhOW0ndIjFMLkEEnY+4foqxMk/iuglVXpGBiioovusolxbOcdx
W3YOr3AnusfDgYCYHyCYno7qfV7csLPrwsBsum5MtgVoowqD1p62NI+FBKtagh220Sh93cg9KGyJ
UIDGKwcKlobFcWbCpM0SNrMzXTUnRA0m+L8Q7R18k/biZJZ6ysMv/L4BEyiblbh0he/kU+UwitzZ
jq+DNpzgFy5BMcbbewQUrmVOzofpAxhBcBG+LrT358Pup37KiuijEc63W4JXGdoAI//X3E+sHJ/x
mljOSUfU20UOtfYbAo0i0paLfsnaC6FdxwvBMi8liJhbVzvNgBgBcRdpLV5u9K61vAGrw8g18n3W
5dbcxU1Xk4wGm5xT4THRo3Nb4BVW4Z/h0tMm+6yWXRSPj5skGFBJQmSUHlTsQetQsVZQ6QaNjWHj
M1EotNO8E7vdIDWOEMe2FFjCmAhV5+DzcV9XyPcsZIqqaL7mZd5R0p9VAymuVttBie/kvwcKJLMG
4Pci6JqPSjSz6fIvX8ExmOUShcN8VvmkN+x0yaTHFNOiVf0OQf9Gx1w66bEwXqTkkHU1Uqal5ade
zYwBDibsU5mlT9GmRJg+i3i+lyV4Jt85SdjC8/qEBlehyXk/5TjiylkLhW1jxVK0XAB73lWyaFXw
gmoOWjZtfr9upzKS+WnVMSFRWZtqEVuNq2etRsChS9b4WAersgAstR+7leovMV9UN8e/Aa4DvWdB
exKI/J3/s2KCRn/IDpPpVHBWK/FciWnuOS4bf+68oU3Qgl5Oet7CfHPodUHyh3iCqdy9U9CToymQ
DHdMbP8S13TbH3qsXztioYTKfhQIu//xZisWch/43uAAdz5LcpEsUmjKl+KIh/Zt1AVpHzkPvbYY
DOS9xT4s4c9VVrZbMWRkmXW+dzS6uRt/SYyBM0weigyOUVhYwUSFnFHPb42i3W16hISa18mmqYsY
Wyg/AD23c1Z9a73llBCXlpRxSlPky4Cg59h0PRc77DSO74AqPrpo9CEXfR8eDbHLUiHzoinlRGax
0Vx4CtJHILFAw8iEAJ5xVKNBJV+VaMbJ2f13wx4tmUuMYwcpjxNY2cUUP1SObKbfop397aeSnHG1
QYWzenj2nocFgvg5qNp8boySFgJWnF+JNR1k7vmu6SY0QHnkuRG7Zrq65K5AX9H9bR/uRFPyzpGu
1XK+tvzQPmUUHxMOOorUKVbOprob9nwOMpBTVFh7QzLQg6cN1ROrZ8tOvFDyKgoKcpqukt5MbSgS
0AUtDZrIjMpXEsRUKAiJGFCBEZXaDt56pCnFTu0bzgau4sDFi+AoRaIwM1nizgiVVxr3Fp2Cd4Cq
kfX5/VTkis2+PKzz/Rppoxk0s6eAhnhm158fAfAX5AVm8XbIi/jQgRdb1pe4DYQDkcpx4zsBMugy
QOlBuezGO/zyTFI0tB3uvk6pY7hPQwOx4X08JjBN7bacPDzEzWXuyZGh2X1T1DOOhfD6bP8fD8kE
KYJDmpjaNcdE5582qaPh6NgGkHeWgbByvwRuX8lguozsHUPqqNn5zF5cIqnpJytjX8jJTHCg7bLR
Vf4vRddVxaT+9qBzZLmcqGbQyRrQXQqlj46r9tPF1eQcfpioBox+x31k+bysa4f1zewG/PV4atQf
7Le6XJ1E4Ppy1eShYQKBtH+RdllWjZg5Sa3LK7NStZgka0kaof0z6sNFnKF1XJ4ngzMs90fCaM0z
EZxNycJGqiWATSeaSCmZ3S8EHzIgCIB7GmcWzHDuaxUjGlDzMx8dats2LDBliA58spNbqqBFrrjZ
z7tXF+tzIU522cadYCJgOfY2kwNN+npBzVYh0xz0KDO/mB8oX/L67Q3tVgbx8w3zEp3bC90alam2
8BWLrIlXT7D1SOb5AKiwp9Jx8C9F7uu6CDWxJbapVGYBq5wbbRaKtKKEyC66c9qwfc5gyLI6wPB1
V6TtQk/fJG+G3Ei7rzXyMFeayiG/Z9kmcoIQ/zixf8UcB3wKRBamxlRhlx1IsYWtsrFtuuEZ+fBR
yXuoSNEKZrCBjQPrRWawVGFey031JiIpjocSHtDxmoK4mu2V6UOKtplfzzYidyceq/GNCPeOu4vh
mNrKVVPMYofi+GxyIaKvYr44VZ24pFyV7aYu95tRqTw0PMk3cd5kcsJXPfKdU99g/jmffcZFcjJP
1G9l5FhA9iOGUrRbNxGG4m6fCzmpc5vZhiqxUfjDDZY72+ZU7c7r8lilRwrPxtFTUepRD2TiJIPK
FBQNVmY2dRlAqcFOPcqAFyhZNCaNLi6iJ0ZSsOqjcplFk5PL9wCOHJJ+debKX5suF3zJ5YI/aNbP
5p/3v8M8qCjbs4ceMGN4/GSjbLZ6jDAyXtc5NWle+z+9r9jz442VwmjkAaeIy+qguAO/ggAwqgCB
zAUpj1SAm2K9eNelkoY4rJhO5Jscp5iCE2dOOM4ncxE3oXm3yoHAoUWRvc2okDoz4b/WXmxWHRHK
msIvcMTf0MLwlwoM8CHg5WVSef/ZnwcZLgUsAZ4pRXC31XtWeVkqaERlYeHLVsYoeLTBAMcOjPwe
tu8xTJxjVhcb+ewVuKUlJ6PxrPgCKgU/4JKwzZ4fieC6KndYDJe7J/2nMv30kCLTl1Zw1eqs8ck7
AH7ark1QTinHKN2b0nuwmh9fMnKqnlEBfs2KFNnqOzmU4UYIf5fcT2wWn/xCa7gX27ej5ss/1eUU
7dEzD0Ei8BEwK62xZxHGjLa6ArVUOvn6WaNzvYtpX0hzgOFmEXqUftUWzrC8dD89vDYJrRF6wBRx
WgFiGYCkn0wHSdj6Rroql0X8CL7FnAchfWV8bOemHY6y/t4Hld3haxUKu6gc8uykMX1FDZhPThXd
3SM5CzhAOmSXjfK52wHfKM7/OpY3UUeC94JhQHj7HA7qW6J16KWaCnci65ARiSfiUdc8BH1jQjK/
9b4vn24ipvPqMOO4fqMftWUh6Nd3hIeM1DDjQ17zmpb/XXG1tE1lld161Ytk+0VYygvLIi49SlXY
9qpzj9lZMnlRUVz3LIz5F0FJgbzJRwAaSD9EC+4Isf8aTHeEY/ejxcTDZgyb2g/o399QEO5Pd2Kb
EJsahTkmOu+mfDG/r/PDQ4+Issjzrz+XD5dmqA7GU58IkblMoKGYOOnK5u+GAXWRYIcO2zqLWq4P
end0eMc3bwSR6GMSDlzltXuPyms5aMppGbJ4PwK2Wa8Z4ocoqrKRmW+MDpEo5NjbtoZFX6t3x7u9
T3JvhDF+opQEaYEOd36grkLqJnqwYETdlhB8g1zVns0xa0oOW205JkXmWpxsjYqfK+rU4CkLyZj/
t8T4gzOnncJgPK+XPwrGjO3I3S3AayVxLWvylNjQb725x1w16gflbEGU0GZSPWCGyOlLVMuFO6SG
6lY91IhgpOUX8/RISaVtb7HzHGCZmqAXXBb+1uN5Q2rXkepDhQtzIws0nIf/nvZ3165HeNYrO78P
RmG5bpUYVqUpwGzJenw/Odv3SVVmA3dmYvt5e/fLfJtC44wTyoWLYNrDoUMzSMwpUb8UvPQdTiAu
jXckixnm7OCWaiGgKeHbB7HU2kvrQv5EtmuLfvuR4lyB4ZbNM1ChQmkmznKjR+VMMcRsjfLgrEiM
6m2Duw5EemuR79znas6NU/rdz1jVn4sHeOWSLyaMXDbGu11hbLKVXdXpICpBzj1poECl1YkodZDl
PXOpzBv+8Oj7tcicWjZdLWSi6U025Dm4REc6IXGxdMZ5jWLspLtQaJb/hkw9QQ24vFezPEegbtIm
MtWZhs90EdLF02SmujA/gI+fxUMvk5XcgNqinO2R09xFjD+xz1G4S9Nz1C6/nsbSitR9SyW9sdUf
JwD6FutyKS7gejXn9d6MNlZGtlRNmRz3ZPM+LHkXSDhxp3R8k0O+EtFez0CKoqNU6X+W7zezJmNr
hpXUxjy0WqsFmf7b/ygkifb4zagKpUqVePZXdry5txvTcPzTKv9QhlI+lu8BMuo9vUZSngq/Ve1g
lShO6vU9bP7+sRyL3uBEW+b4/fr26e1dIvdyFGuWqSppWlWrFRbH+TjIQeHKdFSbx4rKfpppbhxv
tI4wgLU8mcyUdnXHk6FjQezQu52MGQqM/TA4VUfCMdztpRtiGEhcKOaYBycKgKhj+F/UG+JKdxaS
N7g/6Anb0hPUNM1GLTfYxNNlLY7KENh3b8yRictOu6CxYJZ3PwBZN6TCgodrkeqA2H1pYE1y7y/7
cb0PT9dWIpgPuO2HNEz8oWWoBiltf++9TyL860y0r87WWXEUT98uZ0j1VQg+2i4cHXZZD0ZfsTW8
lAwP8Ao2qxTMnt1ebw5xRDH2d/251y42XofWdJnAZE0gWsLJQ0505uQtDWsEJrTRo294fyBy241q
CzEYjxqKcN4JDl28+eKpp5kQjhZTdvGJdKWX6X8x9Oz2CVrbnlPYDh7QBFPDcIXDB2zUgDTPqhhI
pM2cHNpPnd1cd6Ki3sgbW9o2eBdQ8uE/TZZg1TRp7csySBaa15IelXDajdtTTeACkhJV8SnjjCjK
ecJExTwLf0WpAECm92+j0PMAyNZkMo/KEEWxkfOsS2cWmMeYvkAJq68naw3q3KsrxqYvMM+uEovw
vQZV0PBFx3YWvtiK9z72Atd29sz37pUWQjVZRJGhPFIb4TJevk7BYsXdYW78Q4xWr4Xmlsksr+q1
pirJAKjgV7XwLM27txIhcRWtu1ySPtrhbu2XPe+zCKh/FCGvgYrR0VGfksAzTgXWmzo+gjooW2Mr
E7gJhzepYAxcuIxQYp9015JbOnhjue8TulWz/SPwFXOfmVU5YrlJ4e1li7MHnWXTcCCoKi7eEL8x
9jbXsF+4OfxU72BM7PV2wXLp+Y/883yM71hysnBIh3yM6+FzdYLtfT3RR7N78PiYdi67Rhe6+b82
fCFcS9aVOMuD0Xiwjs0s/pDWpa81Wv8oDIM53tgJmqpcLPbRc3lv49l1TK/Z5Tu3s7oP7jwO4j2Y
VU4rcKnGECzeySVrzMB1AFegXB3i7nzXo6Q2dko2hj4quZn6GupqwbbYwiBjOUyMBFgnMv6USB1+
qlxPZKJL8w7IcBpuJBRHMIHDN1aumSsF3sX+/s8YvYoPwqytSdIlIyNDKVVm+XxCM+EsP7ncEBjI
UJg8w20eWIUEgTqdcD8vP+SDAStZksc1wINCHI/KBwvKIiDKKmwWXJ7pvkRXzgKDTIFRmbL7Bi6k
+dlRLddxarhWuvXpfHw1mtNNTczA+ZHOgxqouP8X3Ajoe5MOqKAzJ6oG6hxorb8Nx1JjDVZ6/vqz
pB1j7mXQbAGJRfJU5thviV91GkU+KUGdBXYXyZPHDKGR0Y154bhxYjbbWrGFiMSBPy8Dl1zQo75G
HHe7Q9P1NsOh559HAaLd35RD7r/Ie4asu4vqSMHPjQbB2r0RMebuu9njhh6DH9wx+qOjBNBrA3mr
2EaexgN/g9fciY4BAwyekwdPgU9E9NkEUw3FpovOHCAaadTAFT6J4EVh2EFOXhc7d9xReCs7jJXt
+59GtIcrvWdqaf71Mwz4/N0PhWZne0n0EUYbBuh6Lrj3ZyimO6hjIC11xh8kbSHmY9iOagKjJpI9
ipXUoR1aa5d38rAqeePc/1koel/DD0p6jz1HnfBX61qKZIDh3ZQLDMZ4wM+k6kD3ny8duKEmQIU2
ue010H7RjwDNplczsqw2VM0hp3NzYe2WaahYJmiliux0EEG2a+vfvWh2oVJa6t5h3iU1DfTVQVlN
yK95Z3+5Ne/1X2Gq0A4fk3dW9Ejf+GzE+so6oZWPcLSkBDlmk02HVvyb2lAEKqctgVQ46vL6e9KQ
dXu4Se1BBiXrgFctgwHvT7Jilad2csJQcVA7wVwXDapMHiUUmUtvTpr9BR9gWkxuI5oaxQhcFe2f
MdYAhHLJKuUI+boLbEH5Ke1SOVxUW+LB5XOv8pmwgF5oFeObp6hSlW5HKZDMrREAgUM7s90YlOqE
e/joazyBRLSaN4UEZ+Gsq1W3TqW0rdcg7F0uQ0OESqQ0xfRebN9vP/WL3IvvQUMtI6WqXD3L/dwi
qCdXEiLKkZN4H20zxSa1Hyg+8JCu5R1XvIq5eRw5m90038XcnSr8SUEu4lYGSITwYkrY8LW1TNSs
7O9Qbz3n8XgImoeUE/SW97mbUTj9U1HnpTfcUN0eloxOxdsY6My1ZY+PcJfDawUjUHVHvahmZXby
AF77mhzlpGfsudfbPpvs3gFCGZKzpz4V0A7h7QJc28PBLfoihdk5LwvtZDzycQHXhLOHT/SKRkoe
c44KbfAk8ShLveoAsah0snKEYaDAtqxCozntYAmbn43cnbR4OF5b77PV74MJnI5leYzRf8ALWnw6
NuCGwknl/kV7VVR+e7Zsu0eXWwfLfVUL/VIW7EDssIEoahnSTGbDyeYFNvDbz2ugyU92ra27c19H
86ALs6/w48BHXpW/aWWWYgBIAhsWsMP3yDEfwv6m2BHcAWIzr2z6DfqEi5Rmyint9P8X13gscbDP
vUUFYYrMBZu4L+Xh3rxmGUil4z3dxRRjYqxZP0gQron8KLPbwi8f6H4lbzYkjnPGWoFiF6UyIZBG
4EY4gAD64lT1fIWe0Pn7wKHbMF4RsLkl81CbgmNc2hvMipuE9JSCgNFZBl8AAuwlNYAFjein6LqW
esXVTM/7PEyIEHGFPBsguacnjpYhuL4ErtSGm2VHnO9/TFly7O9Vd6C1UT2d5aFfQGAI8RM/QHAf
d6bqv2hf4s/QVkFhX+3M4aKDtiTQpq+TVaD3G9UIhGDFLuYo7rU24jhTOqzBhuIrIG5PACq7CEkD
mj6RmGDUklIe1LuOx+Wnx6o9YiEiC+zpEjz44nyl7ceslfuWrYVZWRi6Hl2Z20fFm/0jL0gIikFf
O8aNOk2dqAaBVnzeBvAeZy6dDiw8ulfW4LnfA/wDJ4mDpJL/ZKObSMVg5bTSAxpLyqy2jiHgCCp9
dupkSsmCKg56SmiVBy/py8/DOyrqXdvdhGh481BncOCsRy3S7CkWyKlx+YO8+zxagzrlE0IsIonU
If+DxguktOElC4dwFAsJjuF6GkybY5+FhwFjje/Yv/9pU79cjQh2huOeNjKUXnaFSRfa52r3Q5KY
iUqsXAMd/WePZq8x85A7jugzIFoOyzaaWH8OEfIj0fqvO9uWYOl0BXmzIa8dNP+o93H4fvWQJFbX
tc7wda+aQjN2Wg2NiUkiIb1wpO7IzdWC1gN7TmYsLkG1aWyd76zJznY1qXRqALLvo79B3IAgGKcV
qMuFm+cyGFMu6Jg+uOlrAgPI+6rP+Qwze9sQUvYwu7ljLwGKm2x8t43+AAyIrxJWP6xR18WunzbV
0AaLmAvvm+7Cj2wsKHsI3CDU1ThGK6B14EmLIZNxj+/jvU4touwB2ViLR7mFA+GFhR0Mify6wQs7
P4mjT91I8RGM5V01SYCulYWvur1YjzRomUzOqASVBX22iMQmj9eqy3MQz/i3M1IfzEkFpPaInFGp
69+cfg/ynqw97TYU961j7SoW75kinpADkSbvIFDqnFkqGcf4taKv6qOT9LQEifwvTxfKAuM2abRH
Nzy2/4ai0mqc6tAnlGu8Zwg1PQtr03I/DfDVcGp0JtFJpyLe/NYEqqDPt5oMHUHb4oH55yoe+Mtr
AJXKujs6MU2MXX6DdouQSb2U6Azld2qVH0sPkmPQi7ZUkMDqXb71ogxsVyNCNxS3yJAIM2TSxyUa
IMhw7r0Dktms3YPGvOgu8qtooydFxBfkhwA72Q87IY7/YB97nsmlZLrE6JNsEU3lE0Fd+ZxHXVyh
PVQhnZPMlycBQRkgIKC/KVGvD/rkxODqGfibI1Gl1bDs+R+KBZwnhCgmbruDHxnwJ13jpyTjDhc0
2pG0jydYI2A+qokhFwFkMoVhBiDQYuaK7INavEI=
`protect end_protected
