`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12016)
`protect data_block
U6MMyH52lPfMyZZceWWSVS7mKIzushR3s3qUut2veAfJObLNU4Ct+wuGbxm2AnGDMS9Z60O6K2n3
/XDrpSh8rO7I25Qp9aigr1pPT1ajLH9ShJruTQl3h3zDta6Ulj+k/FViBzFX28bYdwI5ZMIoy6Ru
dYO0OyN04gitUoeLwOZf/8Nzr8C8etB+Ql5ktnYqNKGUfN2BSaWgskNSp8skeLHn3Pn+X9cAxYF2
t1ICz//lBtBNLzHo59/cCXpowUQam7nrTlYG6Ieii37HLcxWMkdro3G/gt0XrlAattm5+9ginDX3
OgbZoVcWCF1a1x/dXcGRKSiyOMZY7PA9O0mQf61aeV4Zh38KJTjucYkq00ftH8Z8J7xwZq+uK4Pm
5TAdotQfKCb0LQOYNMSnAWjQPk42So2Nzkzrss1xhcYr9ZvL4eQL5OOj2DOvWauGx7pl/q/Y99CA
1UV7k3NoHyGy5ZjuVhaoMHfteD7mWeSZXvlFI9ULl3ESdn4RK8plYQ/MwaczPnloafo72CV5vn2T
zrakn1dPmDAFrm9px8EBOdAMb3ovujNGLgctw5oY5NclututJCPWsTuRrkiPGpeyvbJOSEBrwLih
fMnx+Af98b52iLckH+PhNNSvXwkrbdNnf3rqGHlsGIyVdy3KQ68sOwk29PPai1MFhDX8Vzu27AD7
EqQn6IhOW+OE9qd+zVbxuE7p+8sqf0i//KDezryK6XffDnR6BhFA+4Ebjf6qVfVq6YUhE3l5EIMh
rERzqwH3YTjIjWRB2J9NlzIkJeS+AB39yycm0d/xlhCiD1KbL/JHfVHy/+omE6IEQAgmb08eTFWJ
6WXd4fBzYBraQRMwXfO6xEnmBgW6Hv5w+epKEyiB42kkP8er0wfuwVKNPuHvLZZZblfYWQkWgGZy
u1DUo1EcZar1zhaQ+KOEWufG9TZYTB4CGBIBLXn5j1tvpUm2GAt5hRPmWzmZsB9zBWLnAdMAO54n
LCnGH64t4oqoHGicoJgfhG+cIZIS3kS6Yzvx+JTsHwI4GhzsAWofb6/hAZCOMFiSb7SZ8q0eKtS3
hwFQUIFKXCOUIlF23IoKqQUNPfOWsou9hIVaPiDmdTSxZUkpLrT6rO0C4g7S7saoXgvDCnZulWiA
LkElqYFplPnklFuZeIXMUu2VU0mTgAExK7GYYvtYzgKC8m07MFvVhayVGDG2QxQgDPsXomNGTRoG
mUSJMlp64WfXcpjVwNk5g0CCO40zqcbYzv3NNfeLnVNw1NnojkBauXrFXGhd3ak5lCrZ4Y+kzMIW
XoD//uEnwd6ryyvfl5tBbDziiOm5QZit9PVZrjAtTLBvIEjPggFaww6OU+kg3pc80JzDLvjaDXiT
LesvmpT7H7gaMYMBDaef06DCLMcJ7bj7NwWfkMCJTGWtnsUGOCFnPH7RgKIOMlvhEpc0hHcsv/gE
m8ijTPB2saus/EbGIBrJHt2lMsFluZSSb5rX1+po9+RMNwD40IhdaFZSQ/6QB5vbFJ0ui/PoFg3s
hWwt7iKxDqk5YcCsAKFo2+pqmO6NDTUXdrsprC7oAigfniQOLWCTTHlDLbxhSExwFGOEddUlSXbG
0xwpoJqrPh3CYLiSHs9UcuvJZTKlqClvbnqgs+zwiKUsXfAIKf+LuHC8Y8HigsohUaeeTgT7waKX
YK8nI/boyxr8Cv2Qe4UolMO5BfR3LtwWittC2uxIAMt4Ua8ebDbpyadafXp59A1GbX+lw6eO1otq
szbNml3RoWoV5FNeCw1Oq0hjvUQ3VZwefthbim9Ka4fSAvyUpaqT3BTv1Lo77BWMd9cHmjO9WcIk
PkQxDfKifng0u9S9+dA4yNpcXgN/fpG4jd7+zKHlZ+lFW0upELk99LrSVvzbA/GkuwG4tG2SuD68
LZQkZXR9naS1KkA3o7Db0+nCFi3h8NjTt1x+dYDyNtCXbZyincxCFyV9mzl/5ORzFdVYGjWoyjuC
it96tWcX2pfol5Q4DiKWW1GMC+psaeJrALqTeJOkmY9eMaHS03ZvIJlCAWgReFkMS+w9N0BapZHW
4WpeOBH5HbAqXKdmBj/J9u4A71w+O/y0izfEWrWPr6qyE1t7jc5cFflPO3+tvsQHRJmNAGPjvA0E
cf1qswLUnoa/p2B69zh43BRhUJq/Yrd6NkfF1LYia/WzUZMQW6RcQKaPf08ytSjZM4oIpmxBESRN
r3GJLCGMYcpo+WOTbaRvyFwL9cSUuScXrh9tiQEeJT4kMsPxVl1VG58x6O6J2BbE8MZ+iYI8XCfZ
e6reFDq+Nk/Dv/UXBi0kS3hngbpxzt6/a0rjOBLnQ5s/YftS/lgkqR1GHczp36OkGsaygxCIMlS1
WKWEwIDOv30TYSS/NIbP0HD57YsLSVgH0Ef258SPDLfmPdYaGx0DPhZIg2tYESgGRIraicBjrml7
qu9/6D09XMQtPwh7Pa4fFgzwjtiZtaNlqGOsnmBCdgLWm0XB2gmtlJ20hN2sKWNxRlcxG/Z14BHH
aaTaH9dL9o4pN+XCuSC4QF/5YFOmbpH+/lubo/tEVkSnsLXjuKcmD2BgQt/8qCM+yK9Yo4v3kFzz
KRLTXqNcgEB2k5QaSsxNDmpGYjbBiGaaDn/Qf5XZzIFCjXenlBETdoK3jbAoqlmD5tGCXL1/ABLh
HgypFVG5XFsXWPSQ062tpzJicsNmYhGKzLkZ0YA8KTjARGYUQow2OqtZYWyyc+XvmwL7P76J3naR
6PlvW6ld1hfDJB9hA5ASNCGRYxCnOh8DwPShJBjUf6j0RgGBC56fjkhD3fUrO+qaHZplb+ai/uXy
x4+KcjQCuK+XV9FJbI30pebtCtiKyNno+oyO2PuVFX3RJ48YeOiENyDa3UX7N60CHbvBH7bQoT3f
c1U4WS1DYveyDNMg05QNv177dvb4Z4jA5fv2ahvInxlGyuN/kSYt3+4SItZOMjkUjXH8lWaHR8b+
GGEB40c89qicSYcVBddNIng/+LF6AH7eO3yeisuh0Lm4yLygMzjzgPAZ+21C8a2M16NcBZHs2URX
/owwPkTvNrp2mw8TpAiSHoW0RicDAK2jZnBhLu2Aiu63SvG5LEtsEghdPMla7MS1Xgf42Mt2NkqR
vhXV0wf7+Lsg5wL5N6hq1EdsKnweWlrYmGy92D8aWeQNUNXzyuTDsVZC9xwLnQlu2cNtfvyRkvbk
N3GjK5uL7UHYxBE23tgdarUyjjwwA9+6Ts8Q6yqo/73wWRg9lChTiGlxrm7YMitl2AcItCmNP+3d
uRzRYdzGNqa/Rq5NVCDoa72Cl6sv3WnPwXKtfN3O9WXEIvOkIp6notrYZ8Rduoc8nJOgpmLRdt83
uoHNkcb22BMeWrzR+9dtW6Qu69bN48uEn2b/70PUfKghK9L2PlO09O7JN7pyIQZ9fIQTocig7bFc
iabH6ulPREfisBx6wyCtooG8CtegFif0JNAL3CNaXSLSSMLhYDlNvsfcGcHyJLttLQA5FtRXg0bq
+Nzo4IJu9YR+HR79CCkOkbLpvCzDM+mdfeQIP71SvHK35xcoWIrFgZm7MqR+v8aJsD1OKbn/RRp1
VUx1jdArJzTG/CGuCJRteKvYYN7a8+YMIpSUDfRnprWqQEUpQJqy7Vx9JymA/5SIpOcavxMrRAt9
tJU1CgMWeCKjTmJgNZcXqayCvxAk2muSeSOCbo2pbPs70If/YZhr8HdKduDvIWzzYpjDmIAZJdOF
YABpfSBZJUQwVV3iyzAc2ghXi+ihOE8W6UdBmH1JiNGaXi5q49m/x2NvyPv6s6G+xv/hT/SFLeVo
8AWw/ohaEd5IQ3HiI88CyzUvK7yxFCDQU+lSVyur9PRYWlDDgjZs4prhs/lj9NtPR5el6wrx+yVT
/LnRVgWO0b8y7oSYDgcAugIhJ0PnW8/u9V4CsFa3iL9WuTFaAslcWXzx8SXE+KaEsmwEDHpk6mLu
TTDPcmSPNXfpAj6EfjKxAPlWN5oaOhxtPtTc8fjiOxP6vN1XemRk0SK58/nY6Yvh6yf6A2DrawVj
CfULFUHw00XRwvy3j9VI5V81J1E8mwpRF9CzEFUBxZKwBxJ9ZtstqqzQS3hqDnNhmi/iGkF9MZaU
LKAjiY9GhNL50tDwm5RhgCPO+Xzc+eM2uzFVq8pN/0fVye67G/JiMZshBCRJVYfLDOBrAOi0/n6x
6M/wFiRGWnloO/1npceAvZS/0oneMYD7KSvFw1ET+jEEG3Kz/XCBuAfBmFVaOV4vIoEjEiMLgXPh
6Ww8AtrItiLRWh0G1V9t+0rTEsV3uYtcly2X0AsdMtVZMRXZo78QOV7PNiS3zzhPgngsY9Z+ZCnP
wj04MnIhH0UT+3ZhEGfJe5CZk/AZIRwsZuDRKVKUXa2Da7xxWoyFaShomyVZHvVdtWFjj4trhdh4
70nWZ2caHg24x1aCH5Ou8l9Z8/a3kUv0D7Lq0NT4Y5vihD/wwOPnT5p2+SV1b3CF811UBbd2TGqB
ofo+H3+d1CdXhSVlnFpWanjU1C2Mp8E7Pr6LQEXYSQqfeEEbup7o4dJDCU+ZQw9YOGdKwpjOmV7j
9BLE6TMl06b6w1K5WrObiyseBPBzuZ4EIUC0wtiRK96aQ2xV6KNYDGSFVWCKZrJLUooeVqXT2tLh
+gjQu7eAuuuYUvbf5YkP8xJbJ3sJZARECJ++bDI9jo2cCSPWZ+/PH6bjfKXpwPQuJYew9XBYCbaf
+Lw7F8TnL9X8EySlQW4WQhftBBDMwNe85JxTkxjjmSzkfGTefTk2NUl5pzbB2klaUGsS7XZNPZi5
QKzi11dx0D0GUbxs0Kr70uAZl/4xmF5HrFZRQZYUQoJs4Q39n2r/itj+iURpByhB7z75IJlyBszD
ykkMH8YEMqsfHP0YNl+9ConghoksEu/idf2GNTp/+U58miFI9u4j0fP/Qlg9Cnl8oPouf2nO9bVJ
WXIQi8KGDBmybnW8S4yiDWK2Mu2xuKuL7Fk2ULj5etXUBCTsYpKYy8q7s85LigjAYrBd6EWZbpsY
0/dKwnHhfXQu2EjuOuDh9F6ye1SgJaniojXJ321v98oRj0WKj461pM6mPXUzW+8SLv6YzKR9UGuI
0P8DnAir+pPswQgeG7F2umXYzYQPyCJe45zndJcIo0C2kLf0tGGGgXBcqadV5jjBIGKhEECis7V5
2SegGWUjxRrTiQEfP1OX++8aNSlv9u/FoeaekydxkrKS5/2pBu4MPUxtLVTm+RLifBelxVPGhxC+
3fJgT2sMsPhhumhhhKCMKBW4VpELbjpOQrcjZO4wVDIue7lOhgdCaV0RxXE7jKq273wTIWnTy1sP
8ZRzvvSlnbLdCmMhsiRNHv+3m7MgQSrAqYSjeO+aCyJ0sSwyldwXNz6LG5c+XWBJnERf5Eubkk/E
CQdBvC/jG8jpEeceBt/TPVyRqp+PRYAkJMa4EKbwceh4xIc1i3F1x5UZpY64e3nuDxaVpAPfHn9y
fhZ8x0LpmJ6gq5IrjHoIOGk9sZXirBZ5flwMERIiUWCfxDLodGT5bsTCnFG87v+GJcvY0qpJVxQm
jAgO/Bw2yJ0SJ9bMCLKOsS/jk8OWEgE2U0no8G1kX3YJRoooG2CuRqbx9UAzgTa4c+jhY1VwBhZl
Qu3P2FggcZdYqtA3yllgSTd8DCrkqYHC55h+Wu55SGJQDoeHWuZgAEO5haDKKSDfOZvQN8VAbxcP
2IaoKFoumSm02uUUcjp4PGMNhmSSJnD2SywzcaNRmBf5nUt3/ye4X8y6fY+bFXQpApt6qQAEu/Eh
HcHkw06Y3nY9nvxkG5q6gWNM93yi8DF5B/Z51vz9RM6rHqDs6NSMn+cGXaTDSok3pFQXhY7Y2AoH
jfsAG50iSR9nqrxEdelAGDNCY69yoU82ssp9CjzVHrUbyhagHFKZXC55uymNY7RN545oCmt8rrN5
1NyqAZduLHjegjU75KFCY4hTu6pytA8cXhC6ktCkVKpc/dlt5cLHyShN4LkIAy6V8gy4U12elNXT
KNT9GgSVJjvK4f+N8vQDTydGgu+pLt98hFqAs0l4qu3M50p/4oZEZh83oDvnxEQgiS/1sMUqmBGy
yHvGJcnG7yQfIZoI4kb1rlP0NsLHzhnkF1v79xBeZveV8Pr/EJlfb8rwBwUF35uTOE6oV59NCUDW
AXaupaBGo7qFeURj5iH01pfn3tbzx+MS2h6XGQf9lH9SelIM4qJ5OMCaFXgOfv6sbkICMlsGiz0m
gtxOgywSLIN0ZjcrG1iNdwEG4hf+onQCFvSXsAX0tV6P3LYNnPNWx6UHXZMx31lFyQz+Q2L8ILDe
wrKxLUqxbg8fNMID1+0D5sKBHntQA3l2JmokhkpeBbUAtsXnqGGliDe3046VIS7urp/RmJprd+iw
XxxZQFmkYQMETKIokAMCcVU8ZS2uu35+qRdPyzAE8mtbpAbV4KNkToPAGqh9zmJFz5loa8osAYvj
5njYLzDnVfVYRhWf6a0j1SBP2fxoTU/fD0DyXATavL+U52TZkrayvrH2x1ZA/ehQT7fey+LiNWSD
bOP+vxwdNvY788YLqFcxne/liqUSUR+DMIQ9dxkZE8hgxq16VDwW/vDe2UmGs4TzL7UQuZIBsjfE
RwVTFI9ZTVabHy6t1o7pFMoJwAhIgjKbbe2/ZDIFh79FC9DGCPxreJF0qnUMU7Gll1lJwiv6wi7X
0BiUkmD2x6W5bN1p9/1xGCqP65vAmh7uDS7434KCRc1uU2CDA+OnnAWEiCIDi82kqz8XUOV2Gnwe
k7VWZM2SxZA6CQHQLguVSlYxx6aCXwA5hLOeoXPaiYmb+2CPaO3BI9VAUTifZmivcVvORnvrVe4u
9uaDTDsmeqfvGX0AxqJZ4Za3NRNcNbC/mPv6U9bNN3mq5OQ65xR8Fn0r/Uq2qDDRdwu+CBdgiHQ/
cCD1KE+TT/pn92njVLouLqUZN6Dh33dGybhLbq547WGZ/0djVeOJK98SQRD6Xl7tviBiI4ZMhODi
/F7rt0DW6Y0LZxQOIM5ya3U4pfVYgKsPF7PWkJq2tKH4gq3+uQqt2BSZhoCjMv3a9i/8jK9XDSnD
h4nWZhbGXBxHUmGvxkdROfVP4VJYocLcyfGUQXXTY/4HoHEUI3b8D07fvRzQQBLdlMOMWF4aseMJ
VIMUYIRJDJAB4O1OQrhnagS9JkXZotH0uhjU4PDgrfRo8iqKnnEwFjHlKKlciVa0+AmozCl8snsp
vXroA4fMWKKY/StflFpLMNta6+9doq4Gte35OkvXqRWmGOt69lDDL/Rk1i+Z8VnZ9JW+zg0nuzzO
3MeozSD2dRK2M4FzHukABxg3aKChZw1syusySCQ4yr24m4gmtCOa6PsAgFmDhNvLXFFwHDaX1foQ
D/SgZJsr5oMgZZmwRfRH/PTTAHUZxadYdkLGwvy+eR3RIFegCm8DJ4FPLSH4A2LaCKKYpQ3B3fXR
rcFVjzoSssr4YxhUscREoqoHT45HuiEySVsl1o60O+Tju5K7FZYba9wjiecXipdKM9YVOUFYHEgZ
OdNGEzn4R6wUpDkboTKs8oQMmUWylmPHd0Y/VxxMKMlSg59mby58fxR0zv1n6LLMh5z8ZkLHYqJp
tlXdrokx+Z1suycNWcHtX7qvbdOwAEgrkAYrosf1WEtokZn7yBg6aKUKC2tvvolCoHeGgHwUnQ9L
yqPvPzBGSjDlXwAQYN3yLRM8T6w5fRqSsKwBA0LtriwAZfEt71bxMPDFnroej4iNN5rt8t3gjN8g
Xfmu4RqBP/Aqzc1Vk8rdoFvsnpzIeu6bqykwX13/WjlN7hR/3/txt8m0+cMOnLfSawrvIYMebNQ0
HuDkK4Vr/Oyq4yXMShxlq8zMxWGkcUJZNHE9vag2KjKLUOC05n+ctg0wJRusSBl/9KvzuTDbsv9a
4ENTxlDF+Q9Ecem8dx7wNlOJ43URNfx1Vm9EFkI2iePJMG/OWezq07KeaUvOyl+X5EyuXsPkN1OY
pibaeDWm8f7hL+w4y7ylp6egBklQBPjrb35IY6f+1AdBRIbWyqZeHcIuDqkqlGb01lm7DsRXGK+q
FGRUBQiFi0QvpvZNgzaLoSx+NVuwi5xzfoCj+WOilcQAwJm5ntqupyHGJ1lSE9NJFJqW1f716FsI
tEe5LO3LhEdxoEKbTA5mYOMQX8O49egsr0hm1/SgOE4w/RjVLgMSzw+1mKi6qSJEEimaXOJi3Ayu
vOBox4TeHy2e7bn5qVXofaMOvgNNQBuoHN/VtyH5ntZlSunuFrl9P0erkkgANy3mYGUB0kRfiM9i
xwZSa1XdzxOEo4FLZOYxgsgyrA5Pae3HMYhCNUMBKB7icOkJE0DPBUCWjxeUSm/oHTluO1is3S7g
g6J5ygACUbW92C3zIyGHx25AE5DxLcPkgoYjeTB7cSwy0KUfRE0S3gZY8/vUl1aQMzgtsOehI08e
j/6v5m+eOENDcpk1htUAkS/6itzvNIKCX4s2Z+sNs40pXxzxkQjPWtgxDYsBZHDUDAB2T66S0J7U
/od2t7k3HV95DkF1C9qTgguE1CecnMxfhpIogZDpK382FYMxuI+OIp2gimeTSL3fRLmqWKRbNhGv
b+1jMKgdSXh2cGc3pjMRIo9MUhL/EUfinF9WSVLiBuoB9b+l7jTUYYgFfHdBciHe8JKK+X9QR5S2
ux3jMVuD3M7yR7spgFQYZT3WugnCsMg353Gqc53Rr8fjq3itoLqBUfr7VW+ZDfdNUQRsDmdbgwM9
9JVINo4xoq804roV/UFhanuccsRWYTV1UtgaC6z9kWNGjX4gJfarzPKyggbOfCysVJXtMGUo4/jj
FM6i0bl0Zn6AONzxtC9BDpaztlufKxAPLLtYx85JdiXZY8/S23+ZSOweEMptsNPt9T1X6fk1vze6
PoXf+r9LavEE4ktoTUEwc6SYXUB9nG3a8Vt2jwgnn9BLql/xcLWDvM8g8V3H8eHbDkuq8ZI+Z8K+
oVvpJNfr9DucIeh+bPAcOCpAKK8VSH19tmUO2FqJVakaB7M8i3+ukTIojvQpnt+PxnzkggX1yvKa
0wZ9uhkyKlw8b87vwQRj4Mk6tD3+i+2OsRQFpIlX/kurINyB9vBA17jdqsKxqPI/PNzsB7EGoM+V
81OWuQm4X52Q0jyDflr2oCrQ+xKEktA5M2+31vOcq2UTcTCV/zJrwNPVieyb92g4tVe9RxdvhwQr
SlWpjecv9e0SzaBDgJpNSjT5q8rFaTzUDtsadvpgLIg/VISH/Uk7xUtjbC0UJ/2ULJ4rtDHQxgEX
CeRoPb0i+iOYjSxrhzJFLfTzEFuFamJo6zA5TM4ISs+3j8AG0G9tefDD9+9nLeMAjMvRHWRh6rfe
7jwW3EhIVI6BrNR+J27T6aA3msEDXX90p1uVs+NkPP5blT37g94aV6y3KvdnodeJJcw5Xloe44Dm
zpSXpROgN0d80pZ+kuUGfFmaOAw4HC3BUwKY2hBWk97WZvGRICrABN9dhvvDzvewXVEy3YZML5Xv
PfkyXlfpp4fj4xyY1RUDyMi5QQI0+ZctnOgwog5Uwdcjnfq/NbelqfzG+Bl+MIL7HQ6X/Sfj5sSk
6ERXahrDaG/ywl9gFG5cIxQYkhAoL8ZIadeX8qLpcE1ytG/drbwRfMz297/EXnFTGAQC+gfmD7/w
VQ62xtTw6ZvoUoIwysdO0L2xzq5/f9s1V24AmU13bm6FOc6jTyHYO0Sp8C5yuMVqxDIGlvL2oFt9
ZDjL23ZNVcdbSggCeo16pIrP2UfnJpXJ5Dzz0oIcq6ceb4cYKrTsy8Yoo7HAOurbJf1922X3QoUL
hQMrq34cRNsZkJyf4Bk89hFCsBlW3fGQuFlXa6zG0dv+jisV45Ey1IKKoVmCd/gftj+j5npaG6hE
vqUfARIk19MP3Th2Oy9Gc/Akx7qubcz/CBgJIcHqnnTq72qRV0fOI7v/vUok9+2DlegU7Ti3842f
/zJbCFT2X4iTnZiX+s2uWfLmQjFSIFRbmrR/Kt/EAbqRUx0WcnoScODGY6aiT3Qxg6JR7OL0P4uH
CXZS0NNPdAg4iloDYZLYk9Lpb6stplobwdBCnW7uzBFn6ix7WVDKx6Ue7WR/oESZLTtnE4LcCv3J
f1F/VAdZXUHXDFZdXba/acoG22UL9EPUcNj8fTDCen1YX/nf+d9MK4zNnJ13LPkvmzMrZfdnweHo
oqK7v8W8uHjS2Xv+GDoRWYYYw5XBuC0CKSLLtQadntoc1tfiHqDbbJilbrs4XDeABJdg+6S5NHR2
HESSlAqcTIEsmFwb1AEhDmklDt9LFeC0+u3zAFTp1m9WkL4JdCnufVt7XldexKdcIP8YAHfhjh1k
wwAr5jtbjJSstZTSMnKkQnS439hcBRAntLeg/l6f3CbVbs5ffOG6BJdxYx86L3Xu5ceA5MyBAchI
/hdqORKg3Vu64k8Sz9zX6zrbi2fE96rYadyFV5FmAu2JRnWNqECN6yig05eTncKTLGOe+OaWu5aK
Hip7cezQeNt5zZ9+CdFTwCOjLl68k+/xSCBuyvEpWwJ+oBJnneJ/vRQmRe9kpliAHQUjumK7Rvq4
ysnRxyH3WVFhWFQq42C53UKuw8Utax4ytMtmiYCtPmsQwzIW4N7gOp1d5apsndUpMDXpamkYXKss
gn+zajirUdF3QU0tEXDpsRyHSxRod/e7rreaQyZ1fM7WBHST89/jr/n0BPimS5f/5i+ddmJoFnH1
szjxHnlJLqaLIwxBkGOcDLW96FojZybrz0AB9SZ+32dPFtPFjO69tScID4/Jg8iWD/sLWfeHVOvD
R18Y2lBGpydh2vwIEEV/qmnz9ejuEs54ujd4s0sdEHA/jFbswkVTElhu/1cAKJujSWUmTfLQ+VUa
sKU+s05J194OuNs7jUyBnDyp9ylRbZ0WqDFnNGG4Be8y9AS1v9lr+reKRruKh4IJKoic1BNSAnKI
zOZZI22smLp70MhNn2cAlrZp9AmH2X1dGWwp4ZaDKSRpsm5zXcGpr2Hagbq+Kskte0o+JVhgiBFA
qsEPF/J40r8EFpl5CNO4f6b0q/p6ENBUKxmprX06P8yRebStQoTp4tK8r2kwDrAHWKkkz3njUESq
udcGWA3Ml9OLQuWaVFib8mUcuW/NV3shSBFkLzyuKbKEReKKpL93Q0fYRcHMQA6HcWoxwKRjYN4y
pQ7WMZ+M+qEvXYBJU7uqm9aNqX1sZkLyKDK5xoivqMG161WxHKOZcaijCoHRTXcbjvmfwB7pSC23
vGQoDSdO9S5C4PN6V/BCZyv4uN3k4NfuhViIVDzGeoioceRR92f/v5ObUc8iM25cd0fRn8zqnyhL
jj8kMt+In1HoouPqj3y9E2uLRFEwzlYNngl3klag4g6fNekDRG8YEfJj3F/A/XMUfrN/mnBA+Ii6
WUELk/soTcP3B0KcgKKiAaLQtAJEPlr3LUUctB3xKOCdR+odRRVAQIgHgsYXGcOggUUuTWOxszZr
tBLDtyKNC+LERXQmw54uDUwsGfcTP3kb+3AJu5lvcLg+W0m0T9kxosfhpj33Fhv6GyJQtLyetzfq
/9hIsoGxKu0WcHQTpy132BruF0GNStAHH2P214G7kfpAQvYwR7hIBSM0xnqpqrUI5w/lg2wNrF1H
5fsneHPlK3E0D9i0a46LCt99BT0+Q1XPen8m2StaNtkeErUMMApOhXFdVb/PHTlyj9U3AEVWJAyt
K2O1O8eqbT36PZIRT0241W8tBhVcRy6ZYOKercx7fPPJr5aW0vY0JxwsvL0620Kqy0h8zVjLjZK8
Sc728g5ILI0u1QQbDDdRevtmJphqnvblaPzEYvqZpw8Gj3SXLJeU8TC77HXgZxEgEVypS7ZucQEq
4E3Lo5nEjiXEEYmo5t7XP9ERL5QaiTEHLHpkdyKC+bVNH8LPbgJMeJBbVKzI7OpCgVVbUBMmfzb1
bjQtW9Bx5eJ8kG9IK1lQecTZ2mqrFpiRaN96MBHV17GeKJaD+DoKUZCHfl1rhwhDduJrmGMe5Ujw
MSrOCAIgOA/b4EX/T6D3dTn/XbTrYRgiuxoO/0hn73zm8Vi+7DGSVQF+AEayXMvbhb4YHLXLw4uh
yIi18wBfHBG5rxYPRgSM4XflyxLJgOWg1rgw6xc2UoOjFH5MroEDQ2nrSdE3IbmWgoptd3fgVVOt
7/+O4EH0BSyZ4VZWnmk4untRV/Cy9rK4gQaFu0yvzJH5iBywct9ipoR/2eWZ8azc6YVK4mcsojbR
1G1RW2ig+4D6Km6XebnWPMsPJY+WR9RSVs0R9J0yq3s06lpoTIsRsBfymuRODoD6LneTA4QPxl1y
ACoMeAr/YJ0pjakkPwrnIwbnPvHzOfo8RRv5WuHNzwChHup0HKSeXInELY50piQjjbxyoU3Is2oC
Un4jyYv9cIUxwYFJcvHa7oYw+vUDVJih4Jq14fvJAo/VdClC5/4Vty8YhY9nKNE2GNGe+RRftfE0
UOziVh+adV1p59Wa7DMla3Kv5oO6vx1R7VDhUy+CiS2CFtKVEmt40BAzMBxHL+EFivKsdugj+pNW
bIackMu6RESbEpOPlUlArXp/kXDoaqcUgwH+y5pJk5v71Q1dBqM7r8vTr5EEDU+HrQMdbIpTLPL5
M/MM6vQRbyOePoy+bFI6lkH4t6p0LUhYSEQPYtqLrilZk7GBkVpoE5mayF1situgVONyh8o07jcK
KMQb7OrVBzQF9distEOSP8zG48R0NARaY4Pw6H4NdoNQVDPvQEaCI5/xGCJFsUV/kW4HVjrwoMaM
idg8WLXpPzW4OWXP5hVimIVSYl2aBHNlWak9+/WVqtUiZ3PMsmTrbEouCne2/CJ0Cz7/WWUi3iEn
5mY7aDHjfD4GyB9RGne1UNfH3Lw6V+ltjmCkWGze2fBdhN5YfZWwQ2taxPfwTVG+xsRdg0ACX0ve
uD8Y8bB2dcf7a3Fp/rVb1S9F1Q7mMEWxbQWUyKsc7o34vWaXlQ4hC7avP5guJqdgkiOdcUztSd42
Lsh67H2OpzWAeu1jql5ydq0Gus/lWsPqodB6EC9phvH1QzfKPhvmq8H7KsKRcqxJJGyKP0CXzw5+
exVN39ae8Inrv0mw8s94u4WeIooNKytXZxLG8UleAR9ywJAbmzKIL+ykxlr4jmLaM3pt23o1iuzf
HWtbqLGj9BytJYWPj6lzvqIAEAa0W/ABXbRf1NGOnlbEt0qASGGk/bH2l1grKCyfwCPs+Mw/75cb
kyaA5tB5NWo54QuBhlVmEaR6x2ZrgmiBfywLSrFMnLjGYvBZqbADkAJR48OzD6q/86+Fs0by1+B3
jIcRYHT1skXpUUyw4XPsG9JbFdP73VktlA3fsihfiVhjHt4MMrHdTHtSVDywj+kWrce6tL4rmqdS
k4CfgteCZGaqg7Rqi/2fHvd6ubBqjR0pWAQipbVIPqqt2qc7wrlCVFYMaT9tMhvtb5E7V/bwWc/8
N7UpGQdldIAF2QjcB2+mA5bUtQ1rLPJHRK+7/UNVNjWnHFNU+Zao0S6P5K2xybUb35I7hLP8aIpR
ExPhkuEhWCDFq724ylYNsFWLhhJpkFRcQS9fPwo95Devc//TymJCGEgRstTrGRYedN4JePqJjPiG
OjR2v2OKGAGygRA5a6bsoesjU1+bmvTp6DD7XLJDph+wd6gP9wG5pDgdTKiHqZZZ2bRuog3xvcpW
WUjsQdXX57XdgnMwGUGhzJscdOsmbzfP/57GK0h8Caf6qieW0/jG6o53B9iP1sg6RwCTFIYc/lBl
Pr5LMqdrwPShB9td909H3WvwnfWPnNLbNuUPBFy/5I1uD6yWUb6IPgxSGu3MMN+il+oKbyV4A4We
xuzALe3KsRE6NjGXY9xPSkIr+EWAYdCW2PZ427nnlwbCyFw2kz7Q+cOm+swRDwbEgydNcI04ytJ+
3UdjPEj7Oz85Bsh9qyetwgfwGOy7ZGCqgoI4gmmYPz+YgOsl65yViUf1N6HNG+vhc1R5vOoIPVgk
y/jOk+GIqS4361tu+4dD4Kqh52otir09aal9QGImfMxG1w8j6N3PUQSVM1zgxXtwvC1fxYgp/xKN
bBokj7yrdwRxkaKPdbH+Lzr5+PTqUt8FuuOpSA8X90JHN3nlFAMQI09MD5iI8Bp6dxe3VD0sh3Uw
RNM+o2EQ52DL7lYtREG7grMxkpPbYWHhbgJ173Zu6IW9ySm2fw0v5Vad2DzJOYlVVFXebQaxyHZy
oyvF+CGLHF4pNcqGsFRtH9gX+1eYtYhne9roDdm60H7qq0COFbUZKx6Vd7LjIbNOCq6ss7xXwpzL
5IX3xKlQTtsxiuRZaLvwcddCAykYo631cQ/tRHnoiZ2U0lSkwgZB5rPo81ciAFf564WBAAz96Cw2
6UKYDEzSPJJ+2JdUAVp1pHR5DcnVcWngmra1FKZmuSwKtOMnDTl8hbLryhHL1YkUmyi42hh4rEom
L63Cj9tjFvnnhWfnKDEw0GrJyN5Z6q/7DbagC9gSem8Qnp70EiBPJwAc4RXxaY9hTf8V6aPSixfM
br6c6HSB1NrDBtat6UqOTX5gPlCIrDLY408CqF0LJbM15kKDTSPBFKKk50wbtJhjUJyNFVsX6apv
0Rw555lAedgLjKyjgUW1yK5jGn/71OgnKhoiJL5pHlXqqt+CY1IYHrRM7gJEfHEeCynIRI1aasF8
s/DrWwBOeOatKw1bSLZIo7PKImp5FqyXePqEAL6+4zMjMIfimygs9GJtSnZFeG1aM8xg3ie/KKcV
IiSUQLQ8BQdBVQPtzDN1VE8my4y+8zPKctrSSLfOhlmJtL4QR2MeL9kxUTkgVdUa44W2aaQGaTgc
OMCIp8/R6pehnw7/2vvL15VZF6r4fZdt2kmlrDWlJrsJyMdYou7Tkt5yiiO3hE9n4yAVqZrBrbxm
4C2kj8wiocKlovubBrqoIiY0uMT0cJre3gne+sac2uJZsHHKEoz7jhPh7iGoWDTm0QMzzfiGa5+J
3pkY8LmjM87Nez2qCxl7Y6ILjksKuWZCVtLRCOe2BK4+ldS1Zk32A/pRbwjDRojN5uCj3NDW2mSp
dHEUbVbve1tM4ZicT/S/SF3io57ufoLp7pJZdjZxg5HxiEzPwc8VzdPAhhlHxOHIy+VRdO7rE/NV
O+Di9mhcC7GR7PYUifwNOubkjLThtZCp1ZReId8teAX7mmaLHRX6c0xW1BQ0TIoFUT9v+tpzMtvT
EJ8W8jO6J9f2u78XjD/vg0xpQIAi1DrURDebuhkxj7JuOrdIFzWHwWtXEnf2ZwtXgcG2VysGofn8
3CfTS0Kx3JpDHZ4gwfAlipcfLnWtSNejmG41RVyjcwduOJWfU9ZIlsU+ZHkvpLyZNlITZB+toamy
XEgxSl6hIf3dhznd3GDJ6LAfHnN2REaBflJ5VMahmtxhwhqkGcgF0N6ccDD5Zx6hzEzAJS8CrIXN
S4BivFitxHj45ly8pC3jmWx8QHGEU6RdiL2LAQCQlhEJMp6B0KyhG83gqh5fUJGyh0X2JdKLr0dE
EV3A5nips7rtgKGBHwByGN5YqfRCpM8m4J6LLCf5NJYSTe7fTCpkJ9HrZ+NS35nOpwJU57u+wX4G
VVUEmQhjtlYxi/9VM2uyX/6l3GAH4CvqL05oNh9fO6EdcPoEUa+2dzyW73P6JlIu/eHkj64S+AVo
UX7nKTUv+SJIwbkznGDLDbohJKgpWPxXF/cwkHmgj6daB5wNPc09rHdBnp+AtToimMznKomg3K1U
sgPTHKeLxfHKHB9/xEogA+bchR9zn1Qtc4+8ii47R//R6hMLp0Bkrly0rdt8xi5X1kQmGV1vmXyb
LqU4rCjTAIN+OacL39Z3BOg/ySJBlxh6Y8nFx9YzcHOrOsMCdOjDNsmmyXeIeD1z5xP9poiYYM1E
ZRXrngd2TcSSxxNEaNUYouJGokxDusBtGg/jwBTinyiIs5XPLtXgmiP+NH9wuSkwIsXoEHb5QX6Z
ei7B/oATG0ldYT1m8L9q+DwwOFFisnymEY7Vi0y/2yeGqrTPLIY6pO/rFWrzYQ==
`protect end_protected
