`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
ANXFqPn+0KwTVCmzRaWK2IuO4nsuTG33ywgAPxSBrTt1lIebjCEQTvcwGL3yviD0J377TDJ2M4Sy
hmuo54ayY2PKtWIikQeemORURU6eJez/EENvSb+ZWtBjwBhYvyvmhBcMVBVoOGFbnSozAGSVmsOA
lxHTBB522XSxTkr97ixy2rAgpFBwSTtF61ZwMrv0vdIx5L5HwNJnc/2vIx5VG/uuvOaBGpKY9oCp
jrDHvTIBohfJbUezpjBGlc0IC/zCrPBXjUI+IiMpZRK8p4t/6maVxHhEL45Gcflg/M8weodNEDfc
cbOKGOYyg1T79ni4t/qWy0DDf9vOxX7VFP1t2g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="UxNvcb9ejzC2KRh/imYNOYv/SURicdopuT0Tft0KQvU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4400)
`protect data_block
NMGW/vc5bkDi1xhNinLOKjCCZyNlQFGXMi1vEGEPVjmVZ40pAyz4dGChea6McoxKiowC1CocLfNQ
BnLe7EbSEA8v9X4D9O2DDCJHeMq3MsT2Y/zJc3wzCeS/tW4SaLWYv0Tbp2nT+rJERuFWDVivmXwe
pDt0YCf7fiIC3h0adIe0DcvC6Q/+85WBYrYtXE+PXou2JxgDeG6jLbs/37n6M2T6gzzfsIJMV34Q
cSTdQJMSVOFw2XtLsRFRsWtpM8HfOIiOdb0xJ2Ejo+ZpVQ/u2bqigVym7BZfHk56N7SMFrsNqzHB
X69VWyQ18P7ISlNYTMLVYZ54HTShgqWOErS0zrRByG/wIns0ZtkioKURnSGmiVYgDRb1v+d9xXPn
X/cHprF9ZNyDM73TKuiwsfgOMUNkVwzwxoH9W0znJaQ6ste2Q7S10PuVcpRBY7Nc95CWlkYt8SuG
idR/e70yDe8kJTlOfY9dgtX796Xdu+SnNwM8JPRhw3BE1zAkoEkrcO6zHPtIovjUVgk3rKcjtn9w
xdxr4XijkUdioSBFj25H7k5TGjO+XVq7EvREzlXSvUZ3b6+bovY/kCyFirQ9FK7g8INjyrwVy7vu
nToQQdATqpWaOonYiUyL1cdFbUbz0VmRKQeZyoa/pSY33d7bslo5ZBsUZIdE0IPgevKeWBbIZ3Sk
iSBGRbgSJJj5xojbHfwFID2uOPGivLNUX/4iPC+/cowUJeEi25GOAJhfEec8Hl1/arCVEyeW5JzL
D0Vcr1KR7pnx99sIS8ap0RnX1Hy17MBAWPcjF4Z3vcLW2biQlU2zo07Lb0oVK/5HfL4NnZrB/K2n
Kswnutoqiq2G1HkTvD7+toTSGnV9ju4j/rcjSrmjd5ou0afHgmw8hl7tGx6pES9iomYYDDhHto0q
95WMrsD3ka0kHE8TuYvii3Q/Ae2jUdlFGKJgC5MtmAnhvsvIigsZmHv/mIfERizdJ6zdtyTNGWLb
IAYd4aXukfP+snGEKXDxMEdcw2geWEbdmYoHBK3PvYpTIibohoAzZYRagqXsdUovjJWHAu9IdNh4
+50vyZ0Zos2Ck59KyeQM6QSQtUR4umup/mNZEIzNtYQjFlQej8XYh23Y2NPHZOY/NXdPpzAWp3Fw
Ays4TcbDDFBTMUfmCe+mkFB1Ttq65mIc8JMCOpxpzXVBk+XjB5XnYUtX++GSqDVLQb+LVYuETeKR
jpoOep2r1zzbLPmmRQryOyipoQMjL8IkLCnDcHxClcO9qoj+DprXkL9aBB5eYTrSpohQVpkBIgQG
39GqnWxqgZjuhcYBOrvTgpdd06D2s3RoFnNv81ntghg1h2Bq16adnCCMUZGSnFvxxBDXB0yBcFfk
eFMrsMT7jD+pjjuqo6WIEYaeQeau25AK2g8p6I2ktMK47yFVXTkBWEUHCeO3N3hAgHqEsFZtZpnK
09DR1hgT1Xgx7naIm8G9OY/qHJ6BwDCJKwjkNjK37gJi3j1LogvV1ZLKZfnPcXALrSu98EAoLmEa
vPMzBRF8KrF4M+oXI75eVxjgXA4kfCKirgwNb1LIzapPf3QT+VCK1YsmrYqTgmVdrvkM+3OxO4vY
IihHOObcwH3moZXDROqsiBlMhFH8DKo/hdKyE7v2V1Rs07nyd8nbvHwkja8Aph+rkraEJFwbl7uQ
mDVAfWW0eIjnCtams+mG9U+1TwwMFZQYL+IQkkptLYZDdUusTFCKpO9U/Jv7gq1w57qTH+c86AWE
iMVADZIcNZuncuNJG+EQXazAlWcolU+OEtTtJexnayCFByVveEy+TfLQQwjnJ8zrOnCiNgZM+AqL
Qk03E1crqfSem1HpTN6w3++B1NZhd8SkGo/foizPkPNgyPdX4p+LxG02qWcVoPCUqGJXHC2SZ3kq
6eG8PgEzHRn4DKodPozYoc5UKFBQB6/4cdzywGGwbVP/51wulnrRaPf25CMVjwvGPbxssFt0p+g3
MmJ3olZ7S35PJOHMASVg/UngLxWUFK1h/zgsFxxF09j/6okpgEpNlOIrpzHCZh7YKV2Nxa+nJn5H
gyIZPtBH3+/jjZBkfPvgCp5VvSpxPpLvqlJgqKT6pj1x1z84wKvld/ejby7YbIAXc1Cy+XCyBxuD
nNRvx6Q7ln4IyGBB7WD7CTOUdAzSV/UFc6m9PyDu2j+ualt040Ew2RRNQoGU9aD436vuQ5tw7Yq/
Jm7nnd47x0xYYXQ7Xk3j8JVwdykFHF2ugzlIV5Q55REWdfnhLMUU9wCSeXFitvT94ysU/aq6yH11
amH9T62jsylYUFhmsO7tbNRzFTjbiEjFIBy29YamwnBFmYCrjkzpBW9V4ERgqEEn6J+T1NBmx694
hDo/61ojm6pFpOpgu13nzK9gVEydFd+L8oV/hVq5O21LcBVuejaWpfzDM8RyF1yUFnCfOQHeESkv
t4xArtcp0dODyqv6ybv6yy67x+D0voLvmRtc46wlf27nSoPWBOIpV2ohU7DRT+py/0lwAcdl7ha7
vQZVV6TUuSJhHxJGzFOOd7z2IkQ+KJoYrsPEej+MP60aBL1BHWtwYuXAvi613BHK0bjmu7GxPGzK
Kcf3VqMWaHGSG5oHjo2llFETuEOuzvGFLxOAShPgFbjKtDQ0n9LU9bLFnqq2cjfNne/qbHk8MCsL
MkUjBBfYmPvArYUNy/cUuR3FzLdba9qNFF4/ssJICJgeFGT0XIkTUfPwTNS20Zx5OHIE+UgGGavS
qF82KJtJ4QddHtRNBiNCCXRmqP3sglu2c4jWGzAgCkMx3+Z84CCyJvMc2kX0LDuJ1HoovzJlyoqb
BYXSqzAuZhIJe+hvzRjyYczLSRVq7rOJOhZpigi8Cv7+W80GCAsHn5/qpgOdMx7SlQyLb0YqpJUV
0XNIO4qM8VUnIw+MuN6h/wSv1FlWGFXc6t/phZ2A8qkDoVSkT0jVnUENasdoehzKcaVcO+zYHmiY
oe3G1TmNy3XVIosml65kMGQyRPQDRu3CFgnazlUl6UkA9AMgLEpdPK3X2gnHxNp2SC+4j7Hexspt
lObDw7G64kDMIRRreApzidzr43T7/JIsvvo1DFnQkTJuPw+Mg5qi9c+08yDk36eWSV0io8RZB3ce
1evh18tZlz4a2wOYzbSRFLvz/Iw7Qa4BtMLGSnx9tBNfTqHwcc0CjaLSfFO7l1ShFRe+3ldCaqt5
53iV8Gyrt7D9L29qx/4a4uQPjB0DcvKxKssEn0WyBRPGmJftfxt+FO4NHyq4r4tUcTaeHH1KB1ZK
F5tNzrg+WDn9K51liURa96616vY8k897+LRS+Bx6zbbsLWgxsnPx5NrGq1Vi8czFaOYD9BfuXqUx
g0URjfHJ03TLx8NGNFcUzxSPt351QJ8VFIc1zPtge+1Ue1syS1drVTyjOhWf5kvzYNWAF7jFPMZm
/wgh+IqSb/7rjRzPm8DK9wN8H1DiLsazFcVEIfiptRXMbTNwx57JZJsx9zqIrFOXCKau1UXdx4xP
IK/KUt74YDBAmiW0AJCVdStp5h8c0xnbAplpxbesiAbjDqhblldVcnCK3ajMkw+x1qzwq0J5UKqN
iSAlziwkSwQco+KUiVNAgplaTj6g1fVKFgV6yPeQ4pyRO970RQjy3JAOTpB/8Q9bjThAvIrMzBFG
l4S+Jr5UKsWcLKuDOcTwnr85EOcaCqgcX4OUa+ePO0kM1k2X9d/7LJCH6VLd1ja1iKnOfxc5sw6p
OmwwrM6ntzHxsTQUF4UO2F2+rZpcZC352925UQY7GIN6iS11Ge0Ka0AXwLtFFVeHDvEZMV5OqAIR
YxVxq43eXRCRs5jYhnvD/qcf2dQ6JXM5Adm+pQfOtecufbDjefzcGWvq4SS+3u+OwHgGbIxe6Yfi
sjVaP6Srf1d2lPqt1Ev/uhJpdC1UcF5WEpLJcD3ICLeJY1UuUbeUPc1JKZH/ZTZM8bHnL+NNSeUn
Xj8AbwdE0fpMsilH3MXogh4BmPcyrpP6+kJ/2JqA/INFDzuN0aBecxitJIdwKb66jsaG0JK53TLB
cbh9n554c6qKeB4txMRRBlRZMG+luDJJ+RC7JjG3gI4JGpzpEZcenWaaUmWl9Su/dStJuqWZF4WS
IKkYB6NZ52s6LJAP0ujTakO36c1JKOoEsQv9kDhAqBcLslR/M4nK3XoDYFILXzC4yUEn3/zB6/0T
Q1yTB3/W/v1kwRx8e3fNDk90hFP441z+KNS8k/+9awdJgJEXRf/BrYtozH1UbAvk+So54vNoRCBy
D0MPzTRiorVGsPh1NFKtnVR1tKsQ2v9ryvckZqFf6rxb7c8Jr6QLI8Jl5l83LkoGxqpknDBeSxay
MOScJq+P3f1XNeMCVZbnV0Z2IbnbwGi6kGD+nI7hcXlHmZntVuMEwvZTsS1zjmlWx0g3cRnl5l7c
/JffB/x5YsQvMKs2ukGhX9ZgoEdfv+GF2Lc4R09d7FX0ikfIwFiDPF0exllid1fTZtje+C/zcS6X
2XhiXIZmjVsCHyrag8V+cXSV2s1bZAQ4nrr4/JM7OGY6/upaeIqykRKNzx8fjAzcGuc34WuXySlF
2dlxQ9Iv0siw88b48mqe2KI2tlyJZHV3gJdhjHmfpAgft7NBwxnM6gQkwr2+AL/9db11b6Wo3DMN
BJc3YBj086p58tTBuXRthLDEnYvBo0A/Ip0JGHWSGLCyawIkZ+YnwmP1WZ8rPz+eIBEKJjV18wwd
S7MPgOJbqV9X5plKsq79Yr99YIVY3iNGOhBfXeLuLUeGj5Dwvf5yz4QGiHRM+Jhkx1wWaNkNAycS
ZXkmJG/Xx6cduGmLy15OjNzvF04kSWDYziaDbIKtStzPi+LmivfSEbkIHe28rFjcNNxmIKjzKIhD
rEAgpgoS5rFP4joWtVSgZ6ueZ9BmWJqgu0YNQRMbBEexXy0R+yh0YBzM39vCLsoqs60O468cwMja
zAy5StwtjOjfOVUUewow2IOJqErDEZ7zws5TpZXisy8yImL0Kbcon5nYDYlT+G1xMtvcxzDPaE1T
X9V72Cj6aBj2hRBDeRXEdRDPrEYhCMLokAIRmX5Hryv7AtTzvEulEVSKWJHnV6t67aRwB5ApKbY6
Vd7CWy4khpnVvDxmn+QkBRsYux/j/GefY/NoCN/Uj2WusMTYCr3DNGqgkJ6bN02lbCRiZL3+ybvC
Jv6idDTOno4lzqCDuk8EDP3G4mVMSwKhyJeX8ALTFm/gQyxYt4RSA6M/80IeSRwLJYXjBmShtTvM
jszkIvtx/8XbkjJ5tB8bssq/1VftOAUSw8rLJzpemixX/hjPnmPORqDmr2e1NZPTXGe2pAGJ1pbN
/mfcF83NCa624HB0Rqrwt1SsvNxJlV38VEVwpRlvV1i39fA8wRXhjzYx2PMCCSU2l4/1R4QPAcsh
LaKCh5zyBJywtxK6/IIp5aqrtwsxKAhFBX3+6jTddU98PUUdDk7MEuZMO/V15qU7ZhGxJkPI0xMP
9Y3iHcjCcyetavgHLoTOoPFwN7WAfB4OV4J/IiE1Fxu8RoTe8tWzDNgrovCl9ce1DMOaGJmcu0hd
vAQwT1ugziFQU6P5BBxeHwf20n2i26G5yeOoFRTPs9AgF8XftRwiWxlqe6l32z8BTuxn/4vrpVwu
cVSdJsBLiTSZyB1K3iXMUSRyivt/fsXSXocEU6XDx83RnOglOigWMhHSbVozGUxAhqnPud0qvHra
M5aHoOb7wUGEEB3dFjj5blonK5GjhTvt1WiqZT0v4RrYYEJ0bb6QWgrNcdsKC+B3urb+z1pEHmfx
F/4KLOjbFUpay8nnu/awbknxTJkwS7r+fPe6vlg2MDVqms4/0z+nNTtmO216oBlk/70PDaYdkc6P
y9JxWaXmB3s832o=
`protect end_protected
