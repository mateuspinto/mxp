XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ͫ��'T������%�3.
��������ߛ��L7�+s�W�|� �Ң��O��֌LK��#�.<��'�'�yeP����wm��fC8A�]�r�d:�P���Jh��Ղ���/~f�2Dm)hx�Ǩ|�1���A��A����x:�-�$;��Ȱ��Px�/���QJV]�U����]Zj�|��ź	�"|�Cj����������]	����,iV�֧>���5=(��F>�F�%+>�uz�YK�!��/��6e���:��#Fl��z1.�r��^�} ���V���'H�PT���7
�k�,�O��_��ԣ �&!<\t�G%G�R��� �~vZIf=g��zJ,�$�cJS��~����W�R���o����b�MD����� ��Zlo���q'�m�j0���8KP���d�϶2�;p�ω�L����URR�ґ�~f#����ݗ�*����3�Ư�������w�Ŵ��d��<t2���������`��uݶ7�,��
�hl��p*t�׋�㐸[5XY��$gXk�R.��N���S�G�-��}Cv�.��r4� �Q_9�D���1�Q��[���1ܚ9��zX���J��д�$ﴅ�kD.H�%WY�k�F��;��~4��M�-��d�Pt��p7���M��5�>��8�!eRI���1��uo�;�j���	�whff��V�9.��i�-X}�) �ACd�r8e���<% �^:R��y�]m�>Ԅ`�ԈmH�a4�_�5
�^r4�����́XlxVHYEB     400     190��U5�1�U{�sv3V��6���0_�?��v��F��Y����y��f8ZI���DbF����u��"V@��:�j�L|_�C0�'�N�a�� 9C�i�c��0�g�2���nk��Xk��M^z˱Ͷٴn=��a�kc�e2��`����긥;���I�(�7��&��P�u:4���� �؃a��a�avPkBՙ/9��n�����t�'f�M�8�X�Q����������**��>y�S�����pe�	i�h�[X�^��׸e��}<���x�3IO9��y� �td�]b���L�7�#�d�C�^8���DB|oVz����N�'�}��Z��jD;%��"�v���E��br7.q>Ȥ�#���v��U9�˨�oEJ����&ɘ�t,l<XlxVHYEB     400     1a0
�OA�+[��R�$t,g3"�dߦrZ�tFc��'%W�C٩�}�!�[N��\��h���
��n2RC�2~3��X	�8S���v�l51|��p���H���������^���5 ��>e�+����|����$��7�3 '�y��r�K ���=�ي|�-�f�YI��4\
�"*0�W#ߠA4�M�Ϩy|g���6��"����v�
����\�䔺��0�� �fBg�_^$�+`�D6������P�j��q<��^"�����M�4�!n�/�]��b�2W��B}]У���t�&BDJl�pMa�����������+�S�S��/� :�i6�z2w�h�(�<��~z/]���<.\E��k�WXըƝ\������d�'�ÿ��~k'6�+�QŎ[�A�Ą�OS���m�DXlxVHYEB     400     130~FIp>p���"	4s]�Uj�^����a������ic�p��3����YlE�/NB��*����w��� ��^^��*H �7�|�T���l�@���oK�� Q���sI��&T��R}`�mUٯw��5���Gn�$F��#p�8�%�3�z��tO�fs�~}}zgFˡH�M#֛���R��9���v��W�g�y
�u�������ЁP�d��+�ZN�`-����\v��%2��g�W�A����&����0���ψc8��N3�N�O��Q{k�����h5|��lG�˵�hXlxVHYEB     400     160�`���E�$��Z!t7�R�#2$ݕ����O���BБ� �d(��.�>sÏ���x$-����т
��O|���^���9�%�x�b|�S+��u3����z�;�}P�z��U�ry�g�2.?XQXn����U�w������W���Ţ��}��*�<�7K��*�G�[7[���N_��!�4�VD���ف~$So�vM�V]%?j���J���,�rB�7�&��)�ߵ��A�H����vR��as�%��}+��cD�2h��h-E������0�(�r�1�����+c�oN�o���Ի? �g�N�Q"���]X�����g��w�s5o�n��ȌkRp�XlxVHYEB      3a      40ð��L��D�L:�T�̓gj�>�Y��~j)Q|y��
7~3�Z����$M*��GM;C��w.