`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
SQ918xjt8rec3W+fhLcuo307qz1DfZ/ZCCx3TefNujM/imwnFocgC3tmbbxgib1h0uHAOV6gtjul
jwntAYPzkt4yCy1cxjDrkfvraOk0mzNZU56utD7Mv9dYG5yR7edtdypWTrEL2J7xklKQHIktVmXS
Zukx6Y1AeYP+fycB9hEQT1P5QaDWXh2GYcViSUeQzUjb9/E9gNZu9+9kbjwIOjsVhwWtTM9kErO1
D4v6spjk4bnk7QbR3vvlImdEUrnZ3PC4wHPwShEsYErXc9NYrBerqQeCdkzBs7Yg1/nPV7uHpwCb
Tb9lKlL4TlMQz77m1oT8El1XNQP+Kb+vqfSSew==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="4tLgG6Axc8/2ShMzOebX2+hZONAWLRUjr5IGwaL6v+4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7488)
`protect data_block
YzM6waCWIt881Hdf4m5mIG9j4zFe8eqWxVuWUhmSkOtG6wheQAYd66wGu9vWxfI4fVuQvyKqYNLy
URBVRKyqDI2q0EVznDNxW1HbYdl5N3sA3+qJTze6JEhu/5T+vKi7rrPOgV9ZhXBOqiB/uU/1Irrz
VbKXe2hzAOEHKtbcQonbEffCcgoM3MYVzuLxreF7Lk/G8KMDtj2XtbkaTe3SiVO0kOyXTdRbMZVQ
gi0ajuVa5zxWiYoMWg+2l1SGs05GoLHvZGqh+yBu277EST8flue2P20YjAwnx3LiaNSFjthKsmUv
AWTAW+PKQKlQ2GrPEgjGsUtVhlDNo11U5ZmGMomKqW/ZLxcLszjRWuQ6V3Q8G/W3Ml0+TioUWnOx
bMgBV6tF+qaiUWTUOzhA4bXOFGojojrEFoli3MPOB/yAr6fCXQzu9RkVQ74uGAyyx7AWWAbWyKGr
rcaB164XEuFKqj6T57MTnQOFxJnTm28KqTOpq1HnSHFC4ec9C6GHS8HNKTzYKdpykLJtWOagfah+
BOe5+XQPHlarjtH2T3+l+yoUa8XlVxNjqPBnTfTDJduMVBHTl0ygteGNkoJcUTbEzrdjb+znDL1+
ix7LL1ZzOqypCnCetONPGDdvYENpSOJZaQj+UupV2Srs/Y+QzulbsC8cZv2Zux35CIEaTcqC7R35
Z7ZMCsv9swsrlVHrKEvE2Ilu+/fQ8Oar6FivkUXQ4ZBjFCM4QIaFNOncpphuWzk3dKxgyGxfNCj5
sI08HlAPRBlTAEUX4UQqqhx6kBX1l/t0W4r/yz+GYorNi/1c0upcNEB2me9TLhYSosL4qnXv5NnZ
/Xu0l2BljxOdfUYfxn2F7mVA8NzxRfNduYsta4hW35NdQk8QnYssJjgO/V14vEIeRpomC4kFk8O6
u2LrXHxLD/p3eYG/wZ6emgxm1YfIB69i2e0AI8YI0rmfipqj1Ts6kxzKBcwvSRHssJoScGpre9wt
qa3VEumHS9omh9cgBG1AZFgU5Qnp+IX6ybmcrhbpq5LkD9yWt45+QD4YDdogQhfzoaYm16NwtGoj
J1dnyhFlqNRVLhzo97A0dA4lV9hlwxzRe8Zix2EklCqT3sRTZyVbigk5EVUCTZ/q9CvP41aMpbIQ
6+GDTMqY/kMndgxnRyFjZahSNS2aHfTLsTNF/mJtGYjLm8zCFuwaFUgDzg7pUKY1G6yaolpBKG8D
wT7R/jvxSWdIMx1ESsOjt/qgBtTw5j1HPAO0jW2vehdSaF3JXsFIe9rZrRPX+ZPO70QB7F87QoB7
tiP44rhVtwJYa6qdrjQ9dcHDDiB2p2jIftIPEV1wl1rrQI1YPDgIvtSz6Ashh0sMmlWgAkrPJdOs
6Eu4QPYheuIcmSzeXYSIdAPBGJ4wrxxAWFkIIeBTijjnE3s8PiTT6hqUQuTwARcXyFs4csUOW9dH
TgHt4M7+DJcqymiJjIGTF7u3RCPJCsuoT2B804sbMTCmlnGBcSoGu/jA4R+CY+QuaggpY6cuyNXr
psXNPa7Ypk1u5w8ThweV2WCD8tTpSS/PJiF0ASkPi6V3OBQFx4r0zkx5cWKPiRIfPI8HYHo7Xeld
IPtjuvkdEschpPiBco4EpT1Z/qFqUYmoNot5fMHfmSnXVYaKCM40eDidR+xR46wI37gSmbFRQ2kA
ongMFFf4AB6jhZYVKjzm7MaEPggpI9vqlA+iUEoffbdRQoE9wDmnSRPttbytGm/8akd+q1eNIJrb
5IjQnTj0BSFriJKBYV7vfptF8dIOSOekouPqVjmKwhYh++29viq0B+AJt5i1Sv59hxbaiIF1jMbM
tDKKw0eqjms1rt11ZoTFCcSKkvsoW99AW1dotDl7i5ouCqzcUxS80Pd2tAZW7gefaqUT5ZGlHEJ7
9K1DhBQumY/lATcJO4wcSm5ono74JpsElosbW3+WzrhpCJ8MtTGa42gTGju9knQcu/KK6OhrWC5Q
B9FtIojT8mdc1AlFBYRglqZusLoavfsXSEQFVrHfB/z2JoTqoUU9dGiTfy8WYv0gFC9+z9ie0KZS
QzMPhyIeVwyrbvPML90uVGBMZlInw0c5mmDDN6XBqwyMH3z+8HCe+0j/Gz4WGTFjwEWygV7XASXf
QGO7qevIG75PvnqhUW5X+zBrzqlD+dqcyFAQgcxjXoqxaXHXQyZ0UR/BndTDMWSjNclCoLUCbb5Q
arF1goqnfsNXTNZNkGS6ELgzgRAhLqzaUv85mpFY+zbjNxbQ0PWAHsWqaJxItgvXO2aJ6PiLRodZ
Cten3dhwh3MLd6g9cRmWZjpIfQ8NR2DmqjYUy82FLhCIGslakUVUs7RSbO0uDaaOfIqmm16zMIKt
TJMh34egfmjUtqSLpdlqJUgWKG1iwmbyQfkAPA6PqAjA8RJBgndsJoaWnpH3zqf1/TbI5kcBv7Yy
IRYefp/uchiDuOlxFt5jt+wgGLzA29S9oQYlXp6qikoHVJ9gqc4WfkfH4NbnqBPS1kCD58PDdw3P
+5Ja3Bz0I+njjO5JZBjU9UJNQDbrslVKTb5NMG5zh86IolTJYbHElkX2RjObwZxUkBW+oAos1foA
mV2JM+kgn8EEInK+E73fCJnQ0AdIVPUzPwlN9KR74bE7lR9UDGlHW9AaKE4w0QvmxYIYebUFoxUR
GKDYdU2SuiikJTUCiwvkxrYjoq1O7s907oF9JY6tGdT0ptvJMzLrNl8xuqduest4uzARvf4zvb43
tkknCeI+3aRPtHFvL1yrIsHeHWhMHs/FrLixYuXQ5vFJiCxf1ZvwRi0+Zu3s6A3EwUupWgA0Ds6C
xR6a/320srzTNupE60PL5jWqIwvWCPql/cx2p/W9QYMqQ7q9HFCbLVjysc4Oj4ulZ9bjvMsqpZmj
MP/WQ6x7GjY7HByS1noRReV2ubpKWje4ZBXaH7mukoOrmtLpM0FZ73exroYHZ1P6xBQuSGn2XxhL
kQu6aaftlw1gqYumEHV43kbp2gQfF+/NR7nn+wQ42tSyZhQIZk57IfQI5rpNGg5XpEgFjLOVDtEz
U+Mlp6xSE4T5tW9WwXA5Dc2HZv3DfotqoEtylcpGP63omViJRKhpfUuGDp1L7ky7aPNUuCsR+uzq
ksz53itqVYaCJO9GKMsMd6kExjzJNaPiuxxFt0DzW0BY5/0peBE1J9U1X4GSd8bnIz3ncbqTLNo3
/DMLbqPYL9dzyLADV8xKAtTIIKgTFeUFWNUCKGX+N1WZpe2114Nue0jcsKjR++g3YvfaZibLyt6I
u5nVKh0zLl0ACuKyBWfN+UZ+vQBUPMJgYPCoNR5tIHno/6Sf1YInAUD7mn6soZktg/2BionKQXal
bFLcKXxkHyNwPJ0+PD/kL1HpjGIS31vBxNyWtm5t7hLksgN+3Zhdo+QKzpYAkjubuCvUeCwoJBvm
YEbFTpsJcXxHZUS484xsXx03t0Zh64ynZWm+WujV9f3v3XE2cISOuAMXzMqvL0bAz6WJcDoJ5XjU
CVQ2GFai8om1xWNasw5K/L5i0XoatXuEuDkbTIx8KJrwTVRca0KygO1Nwrge7r4kMSKolqNKWUvP
9Ozn8Cz62mv4oZZRQcOzYiuyk2+sNNNlqtlq4ZGJTJB5iLwRPJrZLCEc+TRtj+XuvSEp4uNPNJDv
Jh9MQvWPePQ700JQHqxQ+aQkb/qq/CF7Ux41g1bwi8Nyk+WFInVqBuDV2Ap3xtT9mOi+tZfwU5iR
9SBrMiHDOwrrrtsnrpFgs3HOccPhH+gWfWBoTDNoYpxXUaNFsNl66bAr1YUrYV1BT2cyg5kfwKEw
IsCBt2oBTNeW4Q0/wG+sS3PunuvO8ozyV0jJVHmuNCv9587s0v6hNif2AFzLz2MjSB3I6Kd4eC3X
wExatMPbnt1ox6OG9YknIs4OxEvdaBx8a9B6CDd/72/ivFDG5D8YcsDwlshZSYXh32PWSs/hdk8t
ZjID64Qo06NRHxzm5Qu9ZCl/WTlK2liUV6a5MFvlbS8sm/0CrTQB59X0nzFd27Aeoe0003qjTwY2
gp507vPz8a23zuqEBvzeu4kafsKv//iTxQHoytiEk/TiFhxX6b5BapzbeOQHH1c0QoZzQ567Nln6
BcakCt7GvA5Op4JyRus5yfxT0HBw43JJf5eZggoykN3y/+yyzAg1F1hQsIH5j3XipSsv+9yBG2Y/
kxtLWkhY2A81F10tpON5HZICMmXCrzOTKNoslnqx5ZbaOW7Au7ugMcFWJFRUMgYEx/kfv30zzoqL
y2cIkkXMJ9lBrgMdZ5t57kTRSMeloZ9LK4/p/1WE03pxd1oNbNF5tEW7hE8IC7+BATen/AoYTdx3
uTzHU/ElxCfWoVhswL9eLKcPjwHUPfbX8zn5khFu/CgrvatmqZSb0ZI0Yt3ZiZ5yfcbbal9WeDvo
z9ehQABZ2h9CfpBzRVFWKBiDHfl2x2SD1G1KlUAOi6l9ykBSv9K9+S6F6SYE9codBOX/Ds/AZDQj
7GVV56xLWyFdM0uEVKyF9WSMQhqihdXO73RP93ReYZX6qJtrSm/d2YuvCCAw//1o1LUsHc+utpqO
nV9MDbEm5COk6VHeUaHuUV3CEs56a40VnD9mk7ahf46+xhBXBbO6xZzQT3DPyCnlbyIuuVO0JNdx
rWizHPAvDF9Gkif1uXzh6i5j35SMC6zdf4pQB9Xh1pUi534oK7IGhgHvgnlYD4V7S01wBuXoZOBS
cYiJ2L/r5Ji7EZ2vN6OYUTDoty9W4yrSHoNKKwha+vZ3v4amrgHGjcWC+gtG+Xr17m0V9IFhg8I8
yffIQsMuZ3mKuzuBaNuvEqqXqVKr6LphF9t8l4nTOvmGSmgTXBPRBtWnTKEDeh2C5FKNq3s0fVzF
08ITUh+BsjFifvCpSm+jvbAp/6vTtBGOyo/k4KRQDOyjFboeyLJlEobzEn8NhUtIuVslf2Dt1ulQ
Two9XoCp5xu5vqf4bytkHhtugzGQTAxTfEHwd1ltBQ/Co9IQ1RxDkQR4Jt49EhVDi4Tjz0mf0sH0
IoZ2S4Wex7CzOlooA/TNVeisNjC0Seikbjg8luS0tSo2KUc184kSkmZS7BNBnPwuhp/vXkJhlPnw
bOCSnhgNhaQBowBIe+1o3BGybFQdnbdtbRFYDzDzqDwoUDZd50lEmkQRrs3YVCqSgw2x3MCBusq9
9gwg5LbFPm2SNOYlsY6UCVzlv7EGC4hydtjgELQm9HoUsgqFOJIq5AZ3xI0RW/Vw8SAQK1AVkHrO
Iym/AEDtIoHOL86u/ATD0t+AqdJAwdbx8uPqFELnxmyjL3XVoEZskN9ZPbxww6AdqO7gHuED4AXX
0KIM7VnlNd7LiJ3SYPUWbp/s9KkDI554meCjPuRobehuJN3VkRIG7zKR3uUUgHo8bkVb6GP8tRxf
pbQ/McFrV04cqez2EMHCAdW1NI6hljutTw3bVftB7mhfpMMiHdTtYB5IXCSgV47d0O6kM8DVcmr+
14DehgC/PhlSj6SGxFwl30VXoYsahT7IThEe638H1ZwVUqtgHfFcz9s7gu4c0Z8NPx3KghRmuwJk
8w9qB68D/7GJVr2FGL+jCSTyudwRTbfNvwPkCLd1Bo5DIUi7llVze16FUjqhiyCOUnalifa2JbGd
5tpOL2U7PETgtWBNQp1DCg2O7kPMZFIY9Qjevfn+B+blQq9plwrm8IEnk4codnjExFnkY8byWcLY
wHQjCTZoIrBwF8N6TfPRCplg/dZ0DwhPNZrtZoT1k716rpltifSpQnGMSSQtfqpJYZQ13ZgJfKAL
PVtH1+dRHnTW8HZrWwG8y4I0oUdwXf/C5lKsNKyxCBHhwATgDPvuf02WCOVI89LscwEu3KyeaycV
keEDSuOmkf6c7mNHS5rRbMcZkNJL0CsDIRKc2ZF7WsORHacgC/EqHJUd2FKSupsGc1JdkHqfYezn
bPa4rT6cC2cyDxOJ3Luw4FyjYhTqhMmlB0jvGqLS/zwFKfOYosLSomd23tLW3EYtoV07XWPglEu9
a9AlNUe1KFbsD/GEaH5GBq+Gwb2XJhzZO/sC7BlljmSamS5kHZt3499XzNoPpAcOvnAreqMyfmRe
YgOkCHWp3XJ0SBHa2V4n4Q2XvPTG7XeaQTEjRgp9Ecdv+FZVm+zWFoCpfOZI13rSLPl3BXcnnjPB
+oSb/K47vNwuMKDXsqu2sIwhtJTBx3mOsmJniX1ELluy7Q66GkVrp1dKtJ4UbI4R9EXsPGFVB3s4
g1BMyh6XWEqPTNHl4ERXeickwh0XAqnKUgylzUVSXnyw0hcuDJcP7sEoTVqoYLB+/R53OfgtJ+9a
b+Ib/TbsMrwINJlv8lY1hJGtrm2kwl1u4GLklZx+D3mNlZMzjI7xC1viUFrGA1wLwm2O+iA/75tw
pSCuE+sV4QwrtF62NDta1KcPYAnfSOi4kfThGorSjrtmi4YH3s4+Bm94x3Zm8A0W2W2JZeu7eUko
j5D6D06vrImf89E4mnIgt7LW/dRds7DvylW6nfl6vrjyioZwKacWleGW0wzvU4LAWwFex9ulA5Q4
VddAD6Zqb7Xvyy8KGJZMUMoULSWk+NDB5spvH31371bhkelqS3RwPwGdArOZ6F1zueYvAwmH/3Mg
v/MocGi6F3ghZ6cxHCCftBCqJ94cGaN+sZc2mXMnrKfZn2i4WzuCFxoGg+T9jkjBkborCSKh2XX8
NvXvZs6g6tbnEtqzE6DGN+x5jDsYtGrJFRhj6FusOqhlPNAAyBggwrFJK7fXW64kdGh7tMHmfIvZ
uoqjNvykK3LPNOp7pkkYO+aXyxODSmSwmiHHocBRaWhl7RHqnYFbJurbxzf2rdHVYlnL3ZbhqykG
uP+WZkwnUin7KpJt32c7pr8Nt7tvfwuJPzZaHRBtUMDhnnua6r1o6dZ+xox/fPm9vOFx9Vu5QiMq
6djLJ//9fQ7GKxI4c4MhmipieLtxsHDb0cYUKNgI2XFNvjnXeaBVJ4Y4QOxQAg/ox+GyapcjPlB/
3GW+NQJekF2qUZ2P4HXZO4/t0KeL+KwU5IJGKBlfn4z9EvDssKqTH9Zu02LTVUEiFiv42QhcX5DF
LoejrSYxN47Xymt0+NGzPyDLkEwYQ2y9L0e5BV+cBATBs3op98kqWcY11zifrBRSmfXfss9cgT+Q
ha1OPvR8W1oitoCw1XFHKL0imStqEffgQ+Gfn4Yp70AWy29aekj0psBiXFEftYz2adhnySiUqWJ/
HQtwgPwSbqpawaPCfBRRS/mnDXLAI7T26T1RwwXSBG9kfLWinYEO87ykEL359yjcTcukuqwmxF+5
lTdeHPUbAxvGcecO6BkvH9OJqXrS0+m6mFcBH5PNmZ1h1vYzMIFXGspnycrXWBVpaOZ8o/xXN4Zn
ZwTJNvcr0M14+wlnuJw5qyP0/hAAJejxBdNITP4mFY2XnwvNHqJEoJsSzKBn2HTzUpmMrMs3Gf/C
eyom5XTmdMlRmLGHekftfNcfjXCiEp0tOhVFxfaAeeJRki82a3s4dt0212i3Zdeh5odplbT15uY0
7mNVqJCTuLsvP5dfQXuamC6oyxNn8isorGYln5RUHisgfv6Ztpje7EI8d15b4hUU/9NOoxBYq2OC
L0jI7ZBYth3YleE4CyS/VQYUMUgp85QMtxgiJ/EFiuPXkhbjFqJ731dJcMlNK7EklmTZD68FIAMD
dWlWdaU93TKPkKdX+q16tFXM6/TSQbVpj1wl++f48MM3dDDgk4GaEW9nuNwTkFDT6K40513xF3TJ
xCrc95pMrPw17q6ob7xicKGUFDb0pX2RmNc+wlsRNtP5rKh2yichY8hnIbJc+WNBv4WT683qbwTF
AuiKmmdP6Sf8K8dD7hbo415f3xHBN+0wQgDC2ZdvIrK2uF5egZ0L23Auv36icW1vHV9jEtasO/Lh
r8RpKg9br9bUdvIoVkDfGYCsVkduZTO5iA0nsmtUGK1qvAhCMos6gw3qK5JN3KqzSt8Q0+nOKJHs
OUiwdZ3GiwvJT2mBidykuWiqwc6ctmojHi+UJ3wFGelAZDOIARNTUyypF+jgWf//dz//xRB6W0XU
Rc+SGvFPHylgX0xyZT4ACe151LKcj8tnYfRwZr8cNdFluUASQMejsUkcThTL1e6ZDVwMmBJfOoWy
ZJ+MtC88bNqy0pNkz0t8oaVrQbO4Iq/FU/Vh0+rm9vWByGGMjzvkjbBSmHz3UwJORq9TA5vnGO9O
8FpkjJyQbGROg/TPzOS2fl7pC/3jEZ/pTpp25XJhGoqPuRBn2yu9qbKbkkdbUOFvXCfMtwDezmPw
Th9rmeSg8Ggk8m0YuyY7cqfAY+ZVfeNG7Z2YunlATQPltyMJhVWqoNFfI9asT12fqbZUlHOc8e8D
nXFGqBpY/GpanRFME5PVPdk/TDKGfITNceM/IB9PDEbt0I1+cI/xKY0mbOjRaljddhIyOzt7Tgvp
wFgnH78hAp9WKEAz7sMeDQrhZFVOWmk4IQWo8MfA2JY7HfW2UShmwoi77+CYEmQrpli70wA8xgYJ
HsCLccY7S6nt2M4+IwqhK0ElqmtqjD8T16M/FlW5oMxOVLOTy3XsURX1wy6wONWfimZnlbUrmT03
3/UaEbGPwxeTXq1u1D5Y1RDHzOV1Ax/bYhzNNsXC67VMqdPo9RA2VKDaxqMMVFaXV5Cn080fqIqe
aQ0JInlQZqFsS1f9/iNQGxOteKbV50PbAEgQUzTtQJK2sOEmZerPoabp3ntCPgI8PC2oWOGiA8Hr
ljNOiMleyAaDhH7GgdUGSajaP7qsskC5uYPstFDDjvsA4IFTq2KXsV3xxeVKRUj8YqzuCxNNEHp2
mH172fuhTlXInz4pnYQXhoOHmpvLHwTWMspo1jf8NmYRHQPNPMSU5e4NZmM4kxgtKN2CknFXs9YB
pbPh9YiMwx52FEZbXe5KZYLLAn+idwOw3/Yug5AzcndURKSYW3Q2mhLbyMYS4Mr43e7gcS1V7qb3
9lqrShvV+wrBJuELVyYZGmfsv7SMPSB93hViCaSaYd5Njtsdcwd1mVJz49nqTstirZjVopvArtkP
vlutmkMMuRMHEV/Dhh0rN/Hy/syv349YESCe6gVAXArAGyj88VUxF9s6QUUffTTTNV+h9Hei/Dww
69/pZMW7gYuZ/UBO2dPhxzSI9VjWS0oA+8fe+OsczYyTkgBZwhNLb930Oi1wCICG7qgZaEvKMi0z
ytLR4dkl2CSx6sG+1HJExMrApWoCXKmyh+nWvhocowNHwHLHXNYb9TAlyqO8F7K8trAGJrbLEiL2
ZcEifRSXEw9Fx3QY1EE+BepFZRf6QTklnCGUbpwV0DWN34lA3XpQCggwFXbJHfwxoFWmhLk/x+IN
D4rtNfuHKg9ez/RwRpdPnNvSPG8vxGWlpM72agj4umM2NQRMn4Hapoz7Jm8IZ79SUzqtNg8qQ3fh
6qO/Rqj2/rBBlWDHL2PV5vJucr+KDIwB+h1/4TKA4s865hujwQTsgmCAG37C2qZRo24gn2y3HVs8
StYQ9ujL+DtejYbeuDcKb1EjPRB6eAjPZm3lNAYVKPclpyQcoLqnLVFvW7+sXsbS0cwC5posk/gj
LaI7IyVY+dP3OUn4MhUVPHSRGTMrcZPIxJmgJToiYlyfeTonW/lVxHodGhbnkjHwezcfd8IYMpmD
dfboS7X/XjWHg7M4rrmhm8VYj8+NS+E1+7TwlnfH6qKeaMPgAXb4QrS16yBfmxRlwPO7JlsI0eHw
NXz/lO672XxQSbW/CLJAqyc3wRdgjH2FPRY4q6WZs8CkZrJ6slhlAl8WrUgrwsbZTQRYDnGilkop
DC0WcYvNAOu7aKfPr1H4QL05oOKOQFz3q2wRQ/xZa5n9ZvxFkxSxxen0NonJ//gaROkEVDch2YeP
17MlnSpwvAvW4QDuXFKO91rs2WcNdP161XroQq9DR24+/5A2LdQh0etLGVXrs6VelfTg0P8y1i5i
8uWI/M8VNjYdZxwxxal4xJhtNiEH
`protect end_protected
