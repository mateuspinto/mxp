XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��c9�d	�b@̻�5nu-���u�]:#��0�B�z�k��l�E��ai��TX���ջ�����ɳ%�}�@z���E�� ſ��,�kߨ��(,���٩���]�h}��4°���
�~�Y��x�[2$����]�}%�M������ ـ?�aETz���P�-�Q�Ў>�c�*�Z�	��Vv���Z�k�LH�Ы���O��5�xAK��H�P��󎳗�r4G��~D��>�*1[P�f8�;> ����
�b�D6�f8���/�qɕ�^~��<8����L���$1�U��_
Tq��SQ^0��w2�8[B�_��|9��H��i�P�)����U<^���l��`��K�C��$��_��������sRg��Ԕ"U�/Y�bZϬ���7s܋C Z�9�E=Ld���tB��~����]��P^�V!�v�zq���?��{�>�/�M'}:��Pz]��V�!��C��;p�־7�r�R�Z�%���Oդ�E��,iU^�z��Xn�"��+B�4��Y9M�P^�������?vp�i�#��8骋�]���\�dX�,~賑�3!w�w����V�5\�5�ԶV�����n�C����%{G�CՇSW�X'4(���~G���>y�������;�,���tlI��f���͕K��yBä�Q��?T[�E��je�;3zS������<MtS�	ŀ�e}1�:��[h��%��9���^�d��zR%�	��J5B;XlxVHYEB     400     1c0B�ػl/T�������/ny���y�c�d��=q�t.O��
�\��s�
] �tU=a�d�c��h������^U�`��C6��;]kX�]��N]9�1�����H�.���&^���{l�WK�\�	w���b��B�q�P��ܝ�I_ݒ�TZk��ڃ�KWg��U�"�M���!d��!�IƗ�� 6=^���/��;�����.����`0SC��5�Iȝ���9��/٨����B�k���?IU3S!]��7�8�k��v�2�gw�6�F�ן�	~tM;ж2@22|)��d93��[�2-��n�����.9 4�;���ƫ����?~��!
ڹ$����L@�C����]:��ܹ�{h�+&Ȗ!�Z�Ԫ#����w��!��������Q�m��M��۲|��N ����+�'O�ţ�#5XlxVHYEB     400     150dh��,�9�ʅP�;��ԕ�'�bV�;�ESJ�����X��Ao�%8�K"[ߎ��#&�Vj`d�8$��4G�R�����{8�ڳ?����mę�Q��R>�Sk��\���'�\�p(�{�׊¾�#8Z�6���|��m掂��G���#�_3������(�kVg�A ���]�u.˞�W���M�ig�N��̰��4�;��YO�O��]�[}��)��ТKΨ-�(��.�X���.��I���dL�M���!��)���n�����S�ϫA\P���Ip}zc�?8B�+�פ�Ԧz�jЦ�Ȕ�(���.G�dk�o-XlxVHYEB     400     130[>E ��w�0�~���NaM[���B4�:�6!�|)!�I}dlfO�z=���G|ˣ
4`?���S��ڿ�`�7,b���7�.t�|Q���j�nڿW���6�վ)�4���D욑�]�,k�$���|��NK2�f�Υ��!3��=���!�Y4�edY���L��1�ω�ˇ~�w��xJ�ߵʰ��e�-r[�7�w���"f_kG�]��e�v���=MALc���W�(1���B�&M"���5*;FL� �*̗���c_)P,��D�,���0��\��<<�U$�XlxVHYEB     400     160.]�w���_ �/��j����.K�{�)��JKGS���t U|s�c�c�1=^t��4(#�����繲�"�"�����@�厜��/�󪵃a5 �}y��v�0y��!Jy�S�������.�LK'��E��a
eGA�@�#K��?����ؓ��i�33T\��^��L#�"'�Sji�N���U�~�}��$9w��<�
�tF�1m�5���$����$�9	#]����I���#
c��:б:��k+�����~�d�U�<�-���&^"20A��_��W��:�4=�誘L�!�k�G(r��2���v
	m�l����e}VUJ����7���*$u�84��XlxVHYEB     400     1e0�=�'I��:�����)��(���`y\-������6��Ĝ�i��x媑v�TQ��dA��齡4͎�v.xS��EOcr�����̊�0�w/gs� ��!��P�0�)� [��=A����[�(�Y׳����V��M��u���t���-���h$_y�iЭV��������U�|�z�f�(Pj�:e7e0à�������sY�(�3�n�f�C�M�ƃ�߭Ї�pĖm�|���M 6pwQo�K0i�q'�+���~�Ұ) l��s@�2	][��p� ��������f��hm���3�D7u=�)�,�\�5+*�_첡 G6+4��W�byT&�h�8��،�3�{���Kۑ ��jY�ᩝ�Il�	413��Sl�XV�ǣzin��2��%��,����/��p
��8mi���%������/˨=&3/��!��i�&Ê�}{S.�H��BPO��[���hXlxVHYEB     400     1008�^�wAq1F˝P���c��F6���D��~T����oU�}b��g�3u��w`�7x��)�B�xq���K�W��o�IX@��0`�2�R�E^�pD�N
�t��!/�+���ڸmW��\�*�#������^new}7��2*nWD%kJo�V0�Z�Z�1�a��E�}o��P���=F� ���:�I�!AK6_�jW�c��1���dv1�8�)��W��)p��X�C�#����M9ө���0F�^"��@H���XlxVHYEB     400     150���-N�/ ��mUv���oaO�-�.]K!�Z��	��m��W���H�5r��I������L�[���ꂖ�g�je�����v4�*�8M
B�?nR��T����Y#}��k8�P/� �f�j��3&#��8�pw>�p�i�_�d�z�~����D/75���"�	_���4�!��]gs��sd���s������]#Piȫ�B��{3��2�u��m'{��}���$;�S������R7_�B��u���!YK{:�t�p3�4G�a`nEL���d�{ט���ށ�b�DN6�1lN��
q�d���u��٬��a0���2XlxVHYEB     400     170|���|5��ڜ;T����g�+Rh
1���,��>2`���7n�#au�jc�sK�g.�fՏ��u�U#C͈O +q��ME/�O0	b�O��E���iQ}�ft�����X�0��0C�ϐ�/K��:f1VG���	�c��;�2�O9��z�Ɣ��z�'Ħ��K_$Z�"�oXq�k"�l���|�j���(�D�����c�pY3�2�i< P��AJ@!��gVG])_o[���3L`��EE��!��>q���I�-cb۴u5?�<4�G����Dl�dh�e���.44u�^1��'G��q�-N�b�Φ9u~Z�fS;�>g>��nܸ���}�=��5�ș�O=�6l���)��+0B����XlxVHYEB     400     160��",��]�D��Ё݇;z�L�,IƯB)�f�F�{:�p��GE7��y	�����fW������S�P���2/�-+>���4^E}��}�n3��=�d�D�FpB3������:5��)hb���G���#��ߴ�8z�������4;{�p�F'�(/�#�k����� G��v�vpb���{+>�H�A�E���jQ�y���SƎdF�ht���g66Hb���(g���Y�����E;a���߱�,Ե�|�eg%5'x�y���+�����r^��S �g܎I�sVKm��V���/
R�4��,�Y5S�׶ғ���d���/L�n@5!����N������XlxVHYEB     400     180�&��Of�C��"��L)E���P&�4�5�"�b�n���]$�{��GQLB=�郐���ݩ���l8��J1��`	��X2�Fr���Mc�\���p�+#5�Ʊ�E2�'��Ƣ20�F`]�)��~}���d7.���t���%k���@|<j>�g�j�n��a	(�'ʓ��e-E_P�+�hs�V�{���R�盛���v�����%f1�h��0���_:���`_}�By���hB����t�<��o-҄^�>ɓp�%���8>��⤕���PA��0FD�L�?��a9(��v��s˲u���1�n�W�Px�o.�#�p����`Ǡ�7GN1��:�r-�/}�Ż�K�$ �7U+@���*"&�m�ٍJ�	�\�*�XlxVHYEB     36f     180t$����VYg�\.<���տ1����F�c�����M�Xi��*yd�㧟�a��[4g�Uy�b6��yB�����xjzU��T�ɺ"S��f�
;|y
*�-/��́�IVL;lw�.{Wd[;7��%p�\r�Z�W��]������̯͛�6�n=�z���}�-v�g�y��܀<���l�2���יME" `����8��H��6iT,�̻ct�mI6����}��~�|`T6�ҿ��~�֓��L/G��{���..�gNJ})�鰁��,@7���s�p��+Ӝr�G�:(�?9�r��O{?����&A A`�.����[v��N��K�Rd�UX�:���������r�'J���QY�¤�tp�3��d