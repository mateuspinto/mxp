`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
6UkOvbzPXuisbXHwjN5RKTfmyh9SkvpZ76V+vVPGobKYUhAd+C1tFXTv+6gSZybxyZKamvucEdxZ
hXu630ex2YtqHEWK32QhkyN1H7r4vqLVmA6dgRVwOPAgjy6+bSO/Ug4CtOaOKVoTUrc8kyAOdC8s
UirrAayKSKKr11XIbbU64Oh/khjwaKgJWrDpEHTtUCNUBbLSO62CkY6c44cw3PGWjoNbxX8/XHQ3
p7iWmnTAjOc2vBu2VU8k7y9+N+MPlJ/gtj22KpON6Sabvopc1zpfl6DVGa2syddyDudEUtNRUW1U
1amquGG0TgeGXWtBMvKeOiuHk2rnWnlMbp4kWqU+yVltukQIYDThcP310PBPVHytSUZh6OrldbGm
DxoVIGlkBMbOuxr57FkLMl9OcBXU8P1uoUviqnwhjtflfssZ53w27F4bG4fPY8fvQ5BHCsFdyFqL
dEf+5P48UXu8rGUdsWzW48Zoi1hf5Nr2CKKb0T8Hteyo49xn2PJU9aMXgxYWag31ecqa4nJAepQM
KrgA9ttIhR/7C9GZB8uB1nvC65q5auCkNW0cJF5GJH3/G5z6br19bQfakPBpBExlyIgolzwjwv0/
jWGulA6rZT9rBnAHP1SokU4rSKTO4Tftmv+or+8ORzPaaGHI+e/HpDPtyivsVqqlk2WxGXUHWx8Z
5ACF1c9tMUKVUp5t5KVKPeVKs60on91gHN/TzwWLB3KcKQKn02YXBF809BUpnoj3KcIH6iZeOB4L
dMDIu4te8I2N5zPQUFFZ/lAcc9kDHAtKDeMzsY0JzPbhdLzZ5h7+Hu40A6VuYgqHmpfMYUYKEpU3
hHKQdrateyECqkqdnm+Dl0jrqkkVLdDte4JM1PC1eyYzb3XC+O7/CJ3QBkMFIQj9Mx6MYHCNIc6e
2v7kV/8KJ61SNIuh/wlnU8Cq/8EvFg3c7RK0etFrcLXFBuBiB0Yt2DDQ6/aCV+dEmNcXZYV7t7Ny
iUKxnufKs56rpFu47lQUuCFa+jCwe5SSXhFtQGy8ZTsfidq6I96PvzeXBySYr6IF4mjXEmQMgpAG
mUr7TMIAxgvvBiXtZUi3Wq10bl8HMwhIpSYSAPCa3iEKBX9P5FoJNgW/B8XbqmKnjpy2V237s0yA
1C2JN7VbmVAUpl0l8Qu47oa6zqUfPNhS9sJzdVT36DS9daJrATVeX9v2TbR7mEWMTICeLVFtXxlL
4OP+EYbiXPSq3Y8A8w56051/1kmeHwcUxntLCxcY09cxVAEjnsKBBQtdaJWeq2Pnn/NSp4jiGrKM
e2LYyxwgNdhpwvDC9+rwP6GFBCMTd5fzZ4lAeQ9HRRTcP7Nba5g2s16y9pK9yw3OgH4LoHl2s9rU
Ftg6o3caS4o9WFMrCi0pgbxeY6gIMpFesSgUgrWnwCo973KQpDIMBrKVpBb8Xo/NBtxiG64GofQe
Sbst+6u2lc3SRqBhItdj5y4s37hK3VdfD79nwms+mwpq7sU4Se9sNkDBT1n4IkK6KNYFH1H95RX9
BbKzhupW7CfZ6JJG8IoukU/jkd13W2sIb3BoBemrVcQOUHyybzwjM4xr+krUfbmSPCyG24iahOMW
aKIxdo1zDBiPmBuyPOoubS4dbXID0HZ3xO1gtLTpn6d0hPr2P7/2/EzEzxnhG9Vym22qejf8Gobk
2E9dXCDHfLuQxliT3vUgKEEfi4VHuTW+bnNCZPRzku5hw6nOU3Ol2nOAF0MVyDJd4ASzkS4W+mBJ
ss/Kvxndm/QIEBgfvnPNWErtpy/fbFzQ7NHL+q5A6/cqg40Q7SiqeqzhUq/0YolqAA4Pz0aPQ2wV
+UQBtCQ1vptpUP9yE7pqZo0Q2VrDzI+wNQD/dFby/yyb2pU/DySbTGyZ68HQrJBLFZpQ9eYJQIIF
weWLKxUVMAvBUn7O2Z17RGcEV9RTJNlNSUy6XM1NHdtr9AVvXusZN0BU/G6XVfXFF3WTNzYyGArG
dGuQOQKyJTWYlyRQP2nODfXuQoOGRkXJ3waJmSCTIIXy2KShUfjZpO63+zpAfj7mHaMnZ7LJbWXR
MsJ2YdE3iaiVHfZBtZCwq+j6kMSSsMfVmSYlAD5nE381ihvIewdbK2r/l1bC+ycdmZ6WZSIHaZNP
xqPFvP/XegLW2REgldenrog98KfclkIvybD5x5SusdUa25qErPK37NHpnLqUY8VqD2kslJO3Ecrk
YYCEmyh1gQXVrPMhJF9W1u1fDtc3yYe9APQbbuR+y+1QI+r/kfQNqZ322j1jfY5OxUbMm0OoMaVv
8QYvKOoy5cEhmJvOIhEqRS8vFaAvP6VHn/dWDPeNXFlp97tp8mnt0tCPBt16o0VEP16KLqBJveLH
sduQ1p9oDoR21SI/CWoN6dVigWw83D2Ddy/XaZ7yNCA1f1lbuHSHzauTMxsYzsDAaZtXOyoKLEpW
gKTIhZbUEugp1NfQUyxG0ex3c7eNCP3d3L8poeADbL3057UYDRvf3lZHLpDPChoqFGlrUuWfRZKg
AeYKmHCyhBEVYAj0xbDiRRJGcGP/QQXrkj3f8KhfGDO3Kvsr54z/Kd3ooOYY1JwF2Oy3DLHN4oQ/
6fX4ApSgSO6PCNoFAbhLNcnL35X736nsuUgSUfnaGzM90OiY2crQ8/uE94odVmeng9XRhWEmMpCS
iYk0BN/U3cX7iYPP10dAv8VvrqLJkSvNYfvaykvBB5/n/6D3jjX6ZWjRcwOld97Mz6jIrI/vctTA
svhL0byzjVQQpqSBUBoWMT7VnaNUyiU+o+meQJ9VaSJ3V5tOYKM1gjYrPKGU2sr8Lp8JBSMwmK24
aX44HhKIKHd81ljTsdFNdp36d4wFyIsZdfO9jhDeYziA7DZzGyIo+72xvT8I/GteWN4jb0/NQemt
0TT2Q743pNSKN/jGdpy0GrqK5/AR8ffBIKDRWyUztHZ32HIo4SmIoyTRmr7HqaAt4FULYg8pUsJ7
zyZLk2NbKDCCVxaTYJUR8cWaRr+JldxLjtqc9TnI3zHaVy7Vj2RhjIvEB2zwwzSItSVfLuNDZzGY
Kp0jr9FS+cvAo7CXeUsdMnyxq4F0nxZyNJB8Jg5zG/kKkk6gN+0rtodERwGlZiLynJvNl5h7uKRx
jmWmymBMJSZrsrw/BnM/pdMdqENFsHYy8/ayR37FTCwhvKR4bnmBA5ZtLxfZduHujSNbw7J2Fkpx
sJtWL+bg73L7iKnWMWWJQkRhPaQLlFzDBimmVPisLYZyyl4iqrJHuVBcLzLtsMc4RY2/IIOBk6PQ
cgDrWjRA28vGFIXIWVi7+IyX2rmnkw1rCzPC5xtZ0o8fagif9qr0hABmdk63pGMLxleH/b/R3JSJ
8gLKNokZsCaf+e+/JdslRgAAKIme/IacDZs6G9BoaO5j4rm3ik5+uF5MKDUYcxegxNJ0CRVixw/v
kKSNU/Yj7gfGooofbapOaaif5QafDVfHxjzPBUwzxmEj29eg9jElCelUj3u2ogy0YJk26b0LtlRm
2SeOVWdcOOnAO25Gr7Pfy8qTOjt8K9/aKfPMKtM184v/qgpzXu2i8hgrT3w6iU+vP9CQWCZP4F/V
MPTv5kLT5k4ZEToUvRHqk564OPAl56cf1j9IGlLdWq4SHeZjKFOOcg/zr2hvgZY1JGa4mtRUf/yU
DRi/TZONLvximzsHvodXGOIIR6zVhAiD2a9xizcNwlg1cnx96SXwCXKS8KQLTrCNmjE6TL5/JJLv
7TfrVolh4t/5vCCsd8I76p5UCiidOsaSy2IsI34+kNgzjc8HcSCvLO8HjPr+a+liTPtUN8G4C6up
ZcD5LNsNgdfcDDt2M42y7a8q9scbqo9NBgVcOd74JF5OZ6uWW62qqS0VOePUXbc0BZa8ywXIIwwU
LptqtLSoqF/D1QhIwNHr4hj+wVPHohl4LHoMJHZWnYct8K9+c/xMHnOmRsB8NUzyK6W3hObb60WS
gOZj5hrDomA0cqvkVJWJB63Z0kvIHt5u7Owau0OpYFzPDhAMKFMW6Gnp9DLQhreymwT/uwdjHQo6
LrO55XbJwKFF3GtiJLSwLG7N8CkVlTlzBuLrKGRPR/AXP8qD5iK4oFJinAoF+l+v7Dx6madPjOfq
wblATlDSf5P7JkBdpjOAyEHdP7cfefyBAv7N7CpA0OKZe4fZBqLSnzupJSvDE9+4qPAejvcb3yUk
9TXka+1LcZETMM67nfWcfUjTjj1hYix0e6pBQ2uCPcJ8pWRwak2w1qfqpAXbO+bIOpXzZhnP1wrC
q28fKbF490v3k/zba3MFWoT+sdBF9peauyKVmbge0/L2XjXnoTm1CrCcKPLSILnaFTh7SnQdBfy0
eLZixzgtRHKJaICNp9M54IC4B3eJzotn/Gts5PiyGkOD3DY7PjOzIPdlg71WDSxw+6sS66ARPWrH
BI3d+YgIDMEm2FFQVlMSJSdKB6P5RkfSFQ/qPhTfsQPE4Xkx8ItkY+1j7sZAV9lHuOanYDFLbZJV
vu8E25NILA5mfQut+etWaMuFO3hfoBNjJgPMDLzthSgfHAQD7wchAiIpCsiGZ3tacY0hH1d6ADZL
HXbDvflNpWE80/UfesWcmRf8a2O2WuVyWtjtb/7QG4hcP6U6BmwKdpTsVQVFRY63PCqOEw4eMFdw
vZEI47DPpq6eUzWEzYdw1f4T037KjqZSrsm14onIPIIVDPUTacytUZfVJU5FCELXzlF3nwjfSilO
dcoKTPtwtaii7pYN8lxdxL6jdzsjl96UWBgEPJ4nVWhr5AbyNImPIoWoLuGjbuZ+uhnGZjbf2GTe
TAElE/Z7XprGJQyOFzTyeVlw/5Yo3uVrHsW24m3cMAn1h2lcf+CNMsixa5ydaWlGOvwf3YbeZFdh
QJQ7ZlH8gDwFn0hx17vhZ+/XWzUIVA/K30bC5jlLGEsYL+BSOGlzICI2NuloZ4vVWOe965G26P2O
Ib24i802hD0indfJoUJho4Gd4r96FeRNB+GUvSRz0L7hx1Xxs4ISs3aI2QWF8HxDHIntFgI6eqZ0
qPkjOXE5ylVoX5q61waVqYbXQ/H3psqQMxP6S16JB+BcGHNM4iW3YOMa2GUL7Se0foFDlKT3GSFY
bQkM+ER5UJ/jScd6P73DkTCKMsUaapv6+RG+DBuZUVhmrvKg7dSvD4x2DhggKDDLClwfGdEkUKf+
+YqhMWe8Oy3yWz8Ap6jbKBKqfL2zAS/GFIsft0ARnmSaZhtDstyMccLJ4gFmeyXuAE3pRRXbde2R
Riw4xutJYcuzz1vtL6U3CkwLPJ9aZpLKCVve3TgYc6+LFwheFEL1FQEVsHRTIfd881cmZwv/l/Vo
6qPAzbNOER37g1H55uu8n5+NWioXZKLkNfjdzT7MXQH+SOiilUcFrGhaCi2J6sZaDCKkC944+E16
OIWatEzg7ufMzIA8zvyehHGjedOntDHeZv5OX7ZS3oipNlOulpRr6uhovWWquCUlrSmF6t/6nkIV
7xRcL5KnR7MONiWzUh6ru+GXvtLCDG3PoMvx3ZxkW7s0k5DumgeH6ZfcHnVPtL/hsiU96dq/R6iq
nP1LZlQgCmJa4K5BU+cmMLUY6QVnWn5sqVDanCs6jq2lbZisfKKMVXD6ufNYhfHA5DsDA4avolfa
7M/FBCB1qAJFTHkLhIpTRm3kD0GPtFvQwCWX/elv6TP0J3DD7vmqezkrT7kNF0MOlvkI+eENyxV+
P99/wbpUpWH31WTxz3no0W5fwZE5hW3aHtohpYDnFy0nB/tUj5Z7Bjdi2RSMswBJ8sP8kZISzvi2
NgX+lkqvkvyM1Iwu9s+ColZvW7mcWHtVNOF2lBZhC+/GpVpicG4e3M2P/8Kh+MKlQLjK7GXpkT3s
0uJKYHOG+Da6TImK3Zgpmhn5222pN2CyUt99qe+0+zg0Iubl9IKJc8POLZ+vrdzRP1MsPNLShHhG
WuqSRheQVMyPMyRyIaCT/PAgLbZ3jf9TFnkG5WOgTenjsoBtQX0Lm4CEpDczUp2vpdZU8IusHXKd
5TrqOcXG4OkAb91ZQlPqRxbljQPmpXcT88+8Z7OAgJhGL1LgaxmSCfIlMDScVQATGlxjZ+PAqmTh
1iCbRBjnx9r71J6W105SjJePyjqzZ5mNvg1Myta0XhFVkfD6BpFnoC/8txP6sq6elo104PDXsoir
WkkOTeFqiNoD2+hV+lO5AAJw6jpTa+xtB4kaDHbyuddelbquulU8RMneKMT/j4zJZeyzEJUBlhiv
qiODJMelkXCMiqhPwOZHjUhk5W3h7pdS+v6YcazzQ9rmNRTb58NuMGMLSjN/Ts7bmwg+CBc0GzQz
FDhbX80zHAYnrnsX8ciS+VEQx9lF63HoJjZAv8xDAefH3cLgBzen0fGXvTy9Nj0QzStO44FN9K/K
+Ju5flOUsJ34soiV2c4CzV1jSDuXv3RW8lwG020okOhrtO5717MavC89kYRBvNGe2XsLrNeV843s
g1rMhLvP7c3ppzLFtvsg7gXk4/Q0mFFVAfG6z6XRRNx8WT+sNBJ6+3ZkZZmGDdBuamO8pg/krGHm
ruTUEa/kkGQ7i8PjMl01SsCdOxsnK6Arc5DR/Hc0JeU6XZSJzTczaVvk3TItS/2aK8RimHbntdPG
TCfC4vuwISA/rflqGl5UfWN23TAzXFMpzYceAuVUQCjzteZAdKKWfICdD2ZtzcqS1mF+YJx7cKMf
MqwPJvxi9Jsof1jb5K1ehD5Woz7RWE6pkKeJ/cNfe5hQj57xNR1+Vk4MW71j9B1D3ZkQ7i0uVpbD
Sbi5AEeTji6wTziaF7GH3rCPWe+GzxPdN+vVzQI6HE3ImVnNjIX5FiJJTopUbr/mVnReNWCcseI1
HR3dAfYruYItdR64iobJ7ZlpKDPC4Kyu0j31TNNt0cyEHjw3+RByYlFwL7AColnjLlYr6rPBXCf7
Mu07xvOS1+ub6feAScJA/czig2MZLbDDGLhzMSZ96TyoB0URKuNfzaElYa4iXDmJ++kNDVzWrEpm
xjSjnYcMg3aHjvnbWmg3D0bDlilGEfQFX/ivy1168cijSXwuzJmdS65zZKtBRq7Kj/m5CnU+IHOQ
GrYxGXRwlTN8bTkRyVJDFxR9ed5uoMSSHOahWcLaAxkQbYowqrskJW/YjUbbFVFJPRJ7khArjFRh
MlRMUfBhSV0oVRxFIySHE4KAcIyi14Wk9si2eAGfSvg/d4H47JdAhYuQF52AGqe3HVmwEUD5AD+4
ylb5B9NTk5kXwtk5u71tfledrxjbjdclCbIKLKsB/qlJGR2/9lE2fTk9DrOcSXt6ihT+kAHVLVnP
unYNRK5NzziMM4mEZhIGX2ZmOAyKX2SaMBbesw7IqNmsAHR4dRnnmpzpnAHVeYTUm+ORUSCoxSY+
RsQsSxehbxwDmbB5CIU0qw3ao7kE4ESK3+WIr0gbw67OkAU5w6ZUamTca1hZPw3+D9/VxQGRlY/C
SRSzDLfL28K2ttTsf/8lSa/isoQYDsuFmi8NqI1HqWhXhv5ZWEc6y0JlofdWIquqcb2cmI1rTUaD
VVjKHddQAM79D0keEwtBfdAy1xLlOYAetbkjfdCrsBdujwXtoj0cgKfm6tDCXZxZPhuQGobB91b6
QcrvPemR9I++YNh8LJOWroVeHAxru6bBqbIiYAzfjbqW17I16+905Cgir7iobYHByeuJvaX1uMCD
ZZGR2/JBxRQEmK/Cb8QVRvXNJ+n9+6YXvqdro/+Mnfi9YvYVmAIhwooytQZDjbbYQAV4cjkxXIkW
oXCv0rXapVggFwjPGD9e0zqN2mGbtaLxtlqkDMOq4K+jDJb/Wf0zLEv2u8MbKuGJPOI+/T3xN7mU
DeiDqN+uWwkZrYbT1pXzqacWcT04Ag4oSnD+2MuR6IYpj7lnxsBruDHiPk4q2BUO5VFPXH8ujd7Y
SrtwVjUXbnkxi1bS0m6AUc+jN/z8cimWuvOvWrIph//EmEs1PR1M/SQlY87mrjhrcYqwBLd/0/la
4djh/556VdFJh/jg8/lGAj9kqPXOc7d+Vpqp1YXtuhr+eYXmW/wiHBjd93jF018hZpG7MFI91zdg
Dds0wVlV3SDtQyoqjsdddfIaC2iSyOq2z0M7/Z15+aS2OTRhAMFX/TyRqOfer+1olJqMwbw1NIf3
WobIva69y4SH5dD42vdZB15e8nvZneDxeVRb8dGzCTm6o9CI/vLJ4SVi6ouZc2c0lDGUa/N1si02
JaBuiyMW/0AR77xiTCfJsARJMIidvLG+EaHbFzrj3i4WD7L0LvaGbZXSDdAGuSzxW5YAVVmftDop
nLsxhUt2q8QtD2F8Mjc3TMLDLcNMvc6rU0yZ9LdDVjHTp88pzlyuTABbhg3R/HAFe4yq1wnPA8ui
M7ZVHFodNMvjifvuzJB+QFfJh/JwKvgW5ht7tNvLAYmgyrku5u0eZEQH2QzrG/4pSjZQb88MzIRN
98XVRf0vrKadBGkCWaXkBfdFSysAwh82L1OEEe/rFYtvxIxdbJ4oIN7vtHoB2/kp1aqfHB6uuFFz
2L12zWDhDhAM6bM6REALjA==
`protect end_protected
