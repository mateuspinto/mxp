`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
j5RuLD5bzDKwgGv6/tNT4KD2ZAgk11MOsIo6nPRqaETJWC6tTIbDMdff5xNoyfblMcLk1Yn+2pb9
53aclAGQRTxOmG4WWiZJ6TRx8xR2W/e6PVNxERd92EqJh4/BQgk1attBL7TSMM5/fbl9Y9KJsyam
78oRpnHi6ST+OxjnMzViI1m9ifVYhLnoH5mMlKzbweOeeEJd3H1lHurR40EvUcRg9gykf/3y0GbB
jfZ96y4mdhuVdS32bbHFTOcxIReA7yIVo7h+xjvw3sa8Z4HLEbF9/BAjImlt5EHnwT+HuAieP+up
A/EsAek41V9KtaKhpBb/WH3Oh2yZFoJW6u7uBg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="KHN1t7BhPons3iBGEYv+pXgj8+c+ZbJHbLrWeKqoeaI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18384)
`protect data_block
sxdmvHvY6IkEC2FgkaK6aUKtExY4GaPujx/U+RklImx6XOMpvdW1/eyjyDXkXHKTwpY+JUtN4jns
/zW4nzFjmmJFydDFx9sFKSEQK0RLBnwoncLdK0kUXYD9H/pr8u2vSXNs315lP/NQEkAvs/Og25oG
lyntrWIPeZGWKOWbhw88BACbnfFJhc3bfqLMWbKK12J8rPpeJ+1I/SPz2R3fPTGANLzG/pL9YZa6
6t3ec6IAp0w85HWOkcTE2OvvG5XqwgHYAlk5Up4fnSuDq5K4LOBEa2NJ8VK3h80Oh3ChfATiGsJ3
l8ISNE3tn5ip3jmC9oj5lZ1nBWA26FtNcUCDNpNf1fuMVw0grRK4bVPOIAHv6J5DRZuioU5/VXUS
COniIkXCVWtCrO4SX+ANrL89o46OLgiBYjoWmuuy0BjClJdtRL9vKIiohzSPKiG/MlED4D8Tm9Q0
U0NDsYXk3IeadfKpab+EaM3xbrNs99ZOyLUDSd6I1NudQ3MEhe+Iu7tbjS7zAzwkAmQGHSKsmTjI
72qolA4Uf0ZcpOF6HwyznGVq4v30Au+K+ovZWx5CEED67hY2vgo8ggp1aBnx6kPy5YWFbi2dsa/8
M9iRKdKk70KBRTeZEp3RiK0YZZ4WDS7wqdehBFh+FZU2ICvGNHItceXQ3OJSwk11+2EF//QU920p
WzqPmCcrX/0j7HQfk/OTAE5VYsMSC/L0nDVmNHno4R+Zjy2/mLHWcr938Iqq0hLevg3dqn8xw7Qo
ARvIqM4LbPKXymr1XZHtL5VQ1Y6NRRisKZXmD4lTPiioYG4CtMGJQR0nPO7cjZW/oh4BDPVF8seI
JcGcGZyFZW+jtp5wVQ1in0PREcQDCeDfVQRpsXLXR38w7MNC8u7iK8PUhYv/qOyuVf2ih6mts8uC
I6KMQ/FFKlR8LwUEFaCdSZrlnTCz9W28m+4fdu2SjFkAZTLSlXq72ww1m8MlyE+SupZATTFgNxoX
EkAN4NOf6Oqp3rasqvJ6MgLJ2GIaX6VRQJwGmyJwf+VX114xg3HL0+dqbwv1P+9faU2RGkl/zOb5
YZkl18M47wVuGReW5ZGiN7hNcrhtuMd3t14wVT9zuE85FjeQOai3CyncyycF96jzHqmWL/u2F4Zx
or6OJ/T5S+9VIrLwRBMkwpeFvx7JZ1jCS1eGDuJlnlUesgxS7vJyTavKzESFCPhEcTHXgjHpOWcA
wWgCrmzKzHoay4af1jT4gA5JlGt3J8xsDjBmUqtZCC7zcBUT8DZgORw0Z8YQncIRfQb5JcntF4WE
0o4bmNOIhnbs5vaHdK47dHs5WTof7JBdmSSuNf6yyWVuI0ev1MN9fDjqRKgDowza5H6qczPv5Gbi
s8YjLuLnaow+IEZzJ7Gje8Qxpem6MCf/zTLQNLGijdA4eVlJjzyhbBGgwsvcVYzklbyvgAcWz+gf
fBiNz/YulNqcaWsHKgZl5NFjiVPJnZD6U8nrsC/7LPDPoGeuBaaxln4A0qEjld/DAonoMMibh6Ht
y3R1gMWYXRxo8uc+aOENrxiGspgxF/cwZoveY251icghGxoycJ5ArcD0qAjPNBWkMod8aSn5Rrag
lOuDx91vTueEs05jhAduGppk9mrkOJDxRkro3uRk5Fb26Qd910acBF2IVZC3Dflg7FIfJsR4x0Ve
e47ejCN2qtwXPHKIhHp7TibmOy425T1Admc/QPGWuU+pZVVfYXnpi8zfJJQH8mkPioC/CNCH2J+J
ICoCGWPPiNm64KsTbWmfSdLWKx07ElepQhBXmL56s4e9cWaJXy2w/sP8lNnRPNnhmV33OLw9PMt2
TBnXaRrQQA+Ao7J0t/uVlK9AKiI/tew35XL27dgcNgCVl21WHMq+79zb1UEKX/p9J3DWJQVHuUKH
2jDnAfpPMZyzrGY2PTPLKl8gOfLb8gjrr2+yEFJTPBdMz/F9qxYvOdsxiWHA92wEjUQfuqpf4Gdz
jVvegwo0aewCcfhbnZGZcQVhKc837WT9ce7PPNkb9G1BSdIDZmb7M+vt6nDln8H7qSX00zn26vUP
nMqc5ucK1oBSpWFyeP7Eyky+gnd6MjxPnh6/bU5SyNZKO1mZo4jkJWOaiv9XxjrTQU5eTfBVQsuw
3T9XnXjPeSuS+ZVBk8xBu47lkkklPjK7y1YvVHbpDNiPn+hQohKUOJOu04kZ5DrL1s3qqxoSBLGL
RKyAYfngT03Gyi+Bv86HSvvva7YBY3vYiIhHvVUCCuvwdHjGYnuYQyqhgAmjlZf7e6cH0wYl4x0M
11Z1/zgdmKASuquxGAXu2JSTF5pDrQTj0JsiBmfGfVPLXgYOW+fhMlLjVxMQ6i3Wt6NjWhuWrADt
CpsD+6QiRLgjI0oZ3gUcgV9BAxQdURNFBg5sz3Kysg3w/AtzrMnj/Su1VcxkpMDmNLQHHTOa45No
j/9waKiSjQvb7dVxlfOYySB4HxYbU/BLvgsB4vQpME754kFx5jRqNMI4tW45ZOXQBiE/HgIA0iw2
JpUITQd/aTbp4I1CK0BgR0NOcEfUomfb7E7I78TLo6mCLaAdrYgOcw9WusM76NzraspwtIBFGthI
Aks6JONZrZHHudzAj9uVvUzCuFGZBjp1DKMGdk66eUgcDXnwA4Nvdua7PyTgcHXb3/wlIglhnLE8
yGyQgQUF0228JfxpFWHqm5TC+jYWVMT97xKN3yM9UM8j+cRkB8ShapH13V3qAK1tc0r5ShJTyZg6
yX271yCmALSYV7R8UTuA24BDxCX0BRWn6S7JOgrV9/0/2UxV/PEimSABYdZsg0Og48/hnVKodeK5
nYDjNCOmP2fg6+g9FP/Sbu2O7pWsRrJ6cBGPmIW0j1y4DUj4oegs2cDfovjenXycRNLNHj31xAFj
QzKurA4hLXzVyg38EpAc+Y6m4kfQP9zJN7YLrsU8Fi715eXlnMv6gtqAODEr8o62kz63SRrW05ZT
THZ5jjP9TZ/PfX/FKKdSzjyYXvgjSzEqc4eaYgO5MdL3r4oh5lCGhC9cUAJeTOxxbCsAP5g8wqFM
3bs0Idd+f0SW89hWpnDvn8ZckurDOgPymJ4Q/MT70U56TYcjF7Bmqni9s+enxDWOBzKYptHJXFWK
zr6hg7MI3ZusSEwK3WkE2q/plrBabNI1igsf3AZso0g/FgY2JxqB0sFEmLkahgxGLQL5/xO/nKcs
2ImDbAWIDqexj8rNaWp6NHGitzp2F6o7qny9Du9eCOVekRVdWCpUXSHEs1KYxwO9ed/uRe2iavz1
8/C5aiQBNUW0FBfCyopXUCD42W1MTQakBoi4aZu8fs+oUtF9Jgy5P3CQ4nFBU9AqAJcN3f8Wcaz7
3suZxkaU7b9N5yRDEOqg1qgOlvWQ+6KpOcTd24jwudT9udBM9MfJfACsOSfGYvBpYj92FibxIpTM
WOLINN04UOWZ2vQqjrOjv9+l14z8v6XVFKGG9SJcgI1Gyq7zXBNOL/dUd2/amXMx6xKlR1wPbTqr
ed1Pw1RS+VeauGT7rXYLxWfZIEms0reK+Kj+xDslT23s3AchS5Aawf/EupKode2D8yi2CpWMiK3x
d9hKRpzbev1roReY347vZRhRVEr0qm6QyL6jr8Fsxc14Q3uFeuC0QwFnjhWapYvfobBB7CKCtWvD
oZVtkjGKeKk9/75qWQflTjFGR2Wln3n0GNC0VJqiuWDAyCTBnlJsRqyvkVfKrGUj06fDjr+aLZa1
X+WSDLL+84mVPF+NEKXwpxQWqbPYaaPHlYlmxhnA00S40U170h619IMPQrkMLMpgEWWexOlySP4N
8dn7D/A4fpKa8mmv87FISpDxk24eZGw95W/rhiA9D9c/1MmcYGi1U1A8bKvi5DZ62g0dMR4vWy0Y
dlIQzeArxMauTj/aAixnBdF9GfX2pgNHUtDsbAIerpR+c2vvxv9f4VISgM/e9RHihZ6OmF2ydp9f
tqqHeZYYn6AYuerTg5IiEzwR4doRg60NOpgDhWTUxNns32RSFDDJHGV6WneYWahQgWvAb3BMado1
sfXcA/s+Q9AV9sE1IVZMbl57xSOVaMgqbBjYbxjGvx9InH15c8OLRuX2slLml4efTaPDo6vKwvXY
XKOINi8mES6R4E+CJgbL9sVPd1n0SVFjZlVKAzKmsV3H5NwwdGpVlT7hcIqpSbzPQOFmp4TpfB+O
OUl+/Xf3gQ4iZc05LV84OEQDTG5mpoIUOKB8FTwMZzy3FN4Mc5UrUdBo58YO/laTgXJ7Rr4FL36s
AbHT/NDoe/KwExJ6GK/ctg9fAA0IgZdUCzgmbTVkVfCH0CLAMS3iUP73XffvtPt5uQkCU4xYBQuE
1ioN1B/XxKItln4mBphGz3M/hkcqK/ehxWhGX1ynCYOFqWF9BeTmTCdhsgt/XKf/P6edmceWzF37
f/JXxeMBFEwyYkohryrY1zIC5t1EgnZYqKel5SvE/fkhbIA+Jr88M3BUSU8hfYsWDSx5BioC89zq
z+MysQ5iq7AVdsETb1KCHOWAtZEi7YYdevcDAFCqxTiIeSX9S1N3xSkxWrJQLojDtS4GkskxqqEO
3/9doSP/E4udpVwbP1icvt2Ga42Ac6+esFQearOWYIJNZXjkgKM00C8jJp3opdgYX6N/y0D9E7hW
61yIFT2UJ27P1BqwGta1dzFhPSkICrb9kUCkz+hMSc3qAnQyEtN8DYd07ql8hkldAAPJVuxy/M9W
v9fQaKiShltYRNsVlgwJHiUW1MJTyG1lQ9E8+go/VzrP9jjiAbCksgTJJ/ppGpMMPzvA+M7xS77r
enkDnM1FfGLpsgxOyQ1+Wr37uf1DzpfC1D1A5wYWFyBB4gU5UUXPeTxs1qnrfBw0WcPqDzKx2/iE
5HcD7JjfbB0HOZeD2dswMZ4+nAfK5f/4i3Rz6e/w0IqJcgn6aEeXVJ6j6eXSh74xuddD/EqDSsWO
LW2FLc9/MPEFycCQopHpW/Bi8Hsl1LAUd0wcAEmj6wnB30zGqTk+zL/OZ3kzL9iIAU4TrdAG2gex
BVIvnn6KHlphGTqwJR6VLxSIPC8uCn+S6hj0fmc0zynsgBgpkjmO/KidaT3QSfn2Vh/ctW5+KgVp
2gCmIAfNjEnHpyutS3TvNoz6jhKgR5oLLDkibrOW/D+RFnD9HNbsNQiQ2ExIAxsh+lohk/bGZ1CL
BoCpat8DnDCXA3rv21byIZPV38XsUAv62DmqVSjgo8f0ZsPB0UXguT0m/qqHdYaylNgCqCiJL8/4
x3YweM/XCNy/DoalDte9APYNm8EYeUMD5IEhfmruagjfwIL/MvBMwZjzPh/mpjyvcFNFQzMV6FZr
8KMwHRTzZtVgjh9koJZROdFHxD8m5O8SeAPhiKZahp6qVAk3YfZ0G8OYnDEHHx+lCgQEhsImLNmE
oxaZFpQw/ag7kmnRdlkJ95s0vwAAeZef6SQAb8y+1FEj1AfzNuYqfl+9THk1FB6hsaRqcDeQ42BH
9oxihnhfkeVhR82GdQmG5YyMCEmzunDakC9yMmhvuajR57ezlzC8mblb/JdWYFFpXh9Wz1pDW5FU
qVI2aj8K6HDG+SyODpy9jUACKchnxRemNP/QX4mSkYaTXvABJhpg56VPlkUqx0d08KLaKnGKIzmb
RMuEAUgnLAzTJOYYNzc9+P/iivZkes+krd+eu1KIpltr4rqoV2QIorxsOfI0oHkvtXUBtKUy/fGn
JRD9C9K2R8UPawQQmp93OnwvUda4udhA325ZJs97aF/w4AR1OoKIXQWZYnOb5sDiHM7M4faMbGRw
/K2UIWaNf3El8Okxwu+M5A0LwFED/QyFk9Ca1kbiqWUC8VHAsrDI67Iz78NLJVmQyoEbaL9h6cCy
c/UQZkWiz9NcRNccSJgSNtqJkrKCxliHvNL7DZxLrrE55eE1cXGeu8S1le0FrJLZ+JeyJiDUSHUH
xhWl19pSGJexbb4csI3Lzct29i2YZSCNFgTYUpHbEL33QCgy9aqT/bMIXy5+X4E6s/gjqmVYPGin
/lTTuMS1wGqbwIUuf9uORm7soX2zNHWgmPBJ3b6003BpWLbbOtq2ChEko3vDc9IqQI+f+75YynBd
DPdJ5ZO9LBiGps0DCbfM9fOsmHMnaUgrvGBJtRvaLc3ocBJKgsM+pxKjeemCKpkcigpwrDwVDAo+
0hrmVfDyLBTG2NYNGG1iKOpyMHwr/9O2w3mtC80pMBqXPB4hM864LlhBlKXjve4jXac7wpx0iJFJ
DntGVJ4kK4j5whY1IcC3E/Er+/nRzZ1LWxt/LKeu5Smc2fvsbjJ7hl62XTDRTOlHSwp7ky9+nIWH
OvELyv9rklpstnuJ0BiMocGHn/Lyh6EYzqxvkfOb45UtziLjHAphs2cHvLKVupcD3NNzty/Dic90
mxbmYWrxxl4tfR+hdAkIWtBl2ivbKzlcCDqFDUUEkk03ZhHsoSlPGyTJk83hqUSQHXfvzgjY4HhP
WrRwXt3TQbt+WIWRUlZdj3cj3OtCSeqSUTZ0McChtXAQiedXFipQWkJTxxOI8oBzrdrQfw1dSTJg
wHaU6fWeL/G4UPVQ+MQlWU56Ao5uQzwXRxhRj6TjjJ1b775DJcShEHX+mmtKpzJZrbFtGpRTd0FX
nBI5MmbrO0Foa5zfEr8tN0+wZzT0dI2r0LXMotbFi5YcKhGKYDu1k58sy5OINTy5buXvbn7RYcMU
cZ2nz7EgBEZfOUrlIp0jrWHij730TFA+oyr9VLgA0i5EpCO46TSo3w6gJibHGojYs9AXok9A0mMz
NDmqbj7n1J5HGWHZ9uD9wnwLZbza8TRC9/nu0NuTmsKaO7AsMWdVBf//2LFv9+AV1trU+9KmsXVH
gXwLtTEARqjJCAf1Ohz2/Q5M/vrSGtXrFivzny8BFZM9XagSbm1eMu4ZxGJRXQCz/Dg7FoCXewTI
CkWt2nPYvATl3JmH2UuXnf6J/jcKc87OyxIF7Wgxq+rJUUGrV04CGpPe++qXhNNC5gghOSEJXsJl
rlvaj8QEWHp69hNvFSYr/2KeTWntGLh4Nm8yRIKSI7amOzfU0DRgGHI+hyMbfmMJ0KiFnL+VYCJN
b28iahDzCqW5dHPsX2zdSeaZG4DkGJd7ZS4UDE7+QxeounMZOPZuLWkX4wfqryVSJBPvifIjiq9O
/AxRUAYUdFTp6y31AnbHta/njEEn6pB88rYYd113tehGjDuFwzTTqX/18O/Tvtuzkl0F/rNClVNU
bhIBH27fVSNnpLaKlCvGFBn1RKzxjoFOqq4IeLqDINa8r0wAzfYtbeVvFI6UOTZ8Y9gvTtAvNReq
rJw1J/sDguH+R9lm0D4xRbsLcSNAm3EMVD2Gfxk3boFwLpUF/G1n8qD60eh96lkLLkCMeb5DdibE
jqpWC9oyO5gtr7UkQrnUz6oIsLHU8dW+RELG6X/XP7iEhjpNV/49Ed+puAQ4h3LOoVkQ1GBnbc7E
+21vHw/FU4NyHJQn/4+OlgjzYKHKdggNPxHJT2MSA9OdaUVzOPjkBqA09jzvFuOuzoQbXUlKt22v
728cfFQeKIlbG/ISXbNK2K+1HcDJmELqeD3cp8xcaUwtDlX12DB71KKlrIW/mrzaQMmwVItwy1Ck
LekOF3XlFV8vMHPmgL6HZ6q8R2zs6pOpNhrr+8KAIaVJGBvA4DDju13cEvqMHuo//UizDDi6XSX5
Xeyj9aq+9/i/S9TCOVUgfFYZa2HcIG2Do3lN7ZN4oGhiQiCav6RqzSUxZBXZhgw7G9kRRX/9YsF5
xRSlQPBOzJTb2w+rLae07p9ai2obBk+nFA62QSY1JqnEFoY088u6gDxS8wco73b6hz/Yt1Pb/cND
Nkg/REOB7SRASwfSgKNxegxpsRKwKcXsQKR8U4TxQENuQ2IE2iJQVOFj3lUDepfeHwsdwSRuJ/il
oBdhD3t2ZRriq3RCXE1G+3hmC4pmwWHBk7uQ7uaz9nUjVjp/3D/621Ms1kmmqYOkWJI3cOpgq8k9
whdN89wgxz5VTFz2rzlGOpbNUYFZD/3+OfVxhZJm6GyGP8iSFIadPxTnLjgo5tdVEZMwlkLKBIUp
XO+LIYvYIYlihyF7B+rdfMQUE/8kQyM/Xdi7OXSS0pEneYls3PZOl3EPH+tlQcsnzVOCBsgTbXt4
w93bFsQZjB945992EtetwbUPDdMS28SOPJcKeZNmm4+ZGRNTVZo5gxmHdAhS93sLQ0xMUfQYbuZv
VszuWJcFa4mf/bnOK/sDM1OR7ZXO8ki9MO3E4G8umUsmMwGdb3biys/wquZi0MtMuJ6Y6zGj4iOi
aytNdJiscBLHPV9z+osV8+4RmWSJoGw3vQSPyn/+4i4AfpFxZCZPuw75Bh3uDCFYsunl02aBbSti
ipByHrAEB3XuzjOFof/TWnGyF4itqkYvC3CP4HBU9YdHc6xbrgJ3fhNsRDM9CYgfktP6jOpK4mVG
vwPHvee0NbOF/3RnH9pZnCSm2PPEd8hkx0oVrROahNO06YKGUt//Ynh6Zxah+WBIyFOB2HBWUdLB
ovNJj/2xG1WkFZvFePlssQWSHKHj8l0W6JMKq5a8U52Bn+26dCXlW9fMuyvNS6VXzbpBW+QuBS+2
q1m9cq6jg5w5xGDeo2voKRqA8tEUJxf3beIVNHsWe6qRDDR3FOYR3Fxs46AbCPiv3j43Gn30VrZh
rjq0Bsp9Exd6SBB46DQmMDzd06jrf/JPI/SSKWGRf39kEqgB+XEtfgSj6U1tsmWTsY5oFy+wisHl
REOCVqFDG1rJha97jOifV2IV8Og2Zxg1B+Vkt8b2RgISrvMMw6+O3bo3KPsNY1461HtlA5H6Lxbu
7pEjMdfDk+WrWZL9EX0wz9MFnXa1L2W/k8HzIsWY/HiVICNTUCEz3g7U8PhVGCbWxb33eE/+dqRY
AuxLWvEjKTF9vNrsXX5d3RYWApreo6yB2tI7G1xZJZkeikdSzctjnzoJDszBi0RvTn68VezNOY1U
DpvavwiTMQOAFFATM/NNh0P/kDoyAPguZEE5DbluiRP4kStea8aRLdCuFvQhWJLivIyJIVIjJKD7
C5MiBsEYowk1lmk+TDZ8jb685AUP6TaKOJQpRp7B3bFtJf6TlcHhsUnrPaRzsckfgWWp1S6p83HA
263gI6T0Pdc9b0YCnyt1oH6ApJ5SzZksri7AeDgQ+HeIgnSvo+rEiRxqs3V/9pLrj760eYHn0p9u
esCelN1vNYnIABOvDzdP1N3G3V2OX41TAIUcD6+cYL9FcUaprmAxPVJ+dJcN5/XHPnwunvZiaNHO
qBy7ijp42KlAW2M1dZJi3aw9u0WBpUx2u3YV2JhGqt4/2aeib0lvuEOTVsJXVxL7lWOT3kNoS8Iz
MRWFTh7nQ7WCZIrsEF8BP6rLTJInBQI7u2LJ2oX0LAQDmzrVV/rlFVhLsVKIQzJHOZH7cQRDMgJR
KC0BaJbRL8InElABe3pvfc4gOen3ar1hENUdK+cGXgOriDzSxjm5UR1YmptkhLywQIAkMR44kRIH
eyYZplBf+Jah/pNNlss2V9IolSnIt8hE5Uqjtl3hosJ5hCCnIjdjhei4yYicdzabHjofOYjDMd2r
uaX0SCuqjzyPhGjauJMBsQksIUM4d77BSX2GSUtjeU39BbPx8m2hYGtKwEuho8ktYB1ACu7bCeuq
WnUM3HRnO+gS2DW5EkJAMxeCUYBzgVsEvR3mNQqH+US9TtNBh7dSmEtXtAG+AdPsLayfPLMqtezl
n5FfmWWGxk0UzwRxX04eBA0CGTVuixhWfcw8IuYsWAqTALc4dIZqq0plpuSnZFUsxdCDn3kqcGpD
VNrhlcEUgQNW3Q09p5br/UKD1P5CWruQhp0c2smx7K0y/FoKWt4cBpDWxCma/Mwqgqm2r68Qok7H
Zg5ft5zA3b/vot/C5lVvqwX+LQLbEySZlOgqgODTYisDOZCxSDCvNEqjJMMwhvOIMhTGLIElv9Ep
dQc6KHkG8aDRJB4tlmf6WWw3cusN7xHygwUWiADmE58p1o8GfxJ+3sXYg2tyE2iqbcgIeADm14y9
AgnvkYQH7FtV6tWBsCZvp2y5hk5oUGTTFUnBz625CdcUCuvt2nriXVL0TiM4zekDT50514WFOGcd
aIxQaEFnPHeNMKq6RBCpX7wjTPDK/BHSD9xLx1AW7ciyLH93fio/paC3Lp6EVInbuXRTmJIs0Mef
wv7+Kr9vv5qtWleyU6IjobWc9BZA7/4UMjJto6BRZzSJXBhtt5fhMnB2PkUl8ojUnFXjhUtWd51s
cbznV8ixvakuIUBDeg0sVq/D4ohVd+xh+eDPuKqCAAcw9F7U7hcNlaGckfgx41dls15ECNJ1Oj41
hIdSYJ13X5MyIxSyF8OzgI2/bkoraWRbFG4rVZx8V3FlBCuQcFB5SLfhmMIQ6PzzIneTiEZui8yP
PI7uomZplqBO6hhpFd3iH8IwhYCRKNx+9DplEabUDKoRXG89lepPCqMW6vM4FdjfIRqbMcIPP9Yh
Xb/MBEbyQ10GAJglmNKCpPu9vzl8zeXjXAahSz7E2R2dAzm3OtLCSn/nEtdIlqzH7f2kv/sPyc9K
p7WupjCozJ83jhhnAYrHCWJ4li4BCsjp9P3I1BYSTK27xnfhZvAhVeFqQXPHLT84c/I/dwBvPaij
CArrlb6lK7qMBG8gEAE34NlGli203SAh/eTIHU0O7E8jQDZRqV/RBPmnOoYQ7L2f3L1fEkOVCm57
524C7FlKzNR1ZYlGrSoOJzvJ7J7EW1fCgBlXxY8jL90HizVdevo9p/INUjJ1nORI78vq2nOwkyNL
rjW7TxufTc+djXlTGJj4POJKPKkklspXQPD0rEn1bw3v9Y7hFhAWGd2RN1/afLT+52SysWnDkHSu
4bQ8oi8QVb1ZzkncotSh6OUrolN3EXrbIatf3PETjDwaPH0XF1N4WF7OKjn9cwUDCtk2D8BhXieU
rdNLT5zLGsw0tbBm0wVjEJpURtnfFKHnLOdqja16yFWCxpQ0UwZyPUfTwWX+ssPe6YwhfJovh1iQ
ZjbLEqC14KqWY55zmt0yt1i6kbUFmqaeyLkUGhKBQzq3S5hmvw+rvbsmc65A252a9KywIa+fIqQa
P2D+/0kWpxmqppMmPHfcFMKqwWtb4i71SqpOIT1ESPZqnaIxiYaSRqA88qL7T/kiGv7313Vrui+h
zbzr+0xGNkCtZ2IvVyVUw224/Jjqr0gPZ68X3ZoZnLzzqnDd74jBMybj/P8bONdwRG5H19+3roA7
zdzFy71WQ1zL6fSGnC5W7HRq9pa56HDogZ78FCW1Q/bA6fq8+OJx/efnFORq9AuX9g8uD3Z4NsiZ
DvUg2464m7N19TXc4XrN0M0GsKjilMTWaIDTLG0G5WXTX4Cp8aQRGSllopybog6Nh7mP4qatxbVR
o8PMGD0anftrNopN6lTGnGrv8acOFf5OzfUpEwAqTegr3uKixuk+W1N/nFTxdRIpQNrObL5CNSLr
7EsihdDX0lx9R/YvVpB+GfymaOCVFhZgORQHO7CDqkFjQewiN2E6ivKN6/duMfScPK9kvGpexv+z
6+nfb+575PVeENHLra+LaG0EEN2U0lcUcqNcNw8FL9HrzRJXRKSZrbo6bePbd/djSnMI948F98sg
z+/9WPk0p/Q1nM9nGmfFoNSWUo62TNu9HdiLdYNYELjHLUisjvger5vbjx3QfChXlAbTtwN92xnv
FL6dJAOIRQRZ4CqGMEyZI19I226pSCR85lZKIjiMtpBlhyoWVIBU0hyOdhSKsA4szI3h0Lyn36d3
bJWgh1lOw0lQddpl604BrXQXVMNP+mT3UDtXl2e2slQfkH3u7iKvYBTyQbhg4UwM7GrJ/cgZYTk7
HgFzSOUeuDYZnYbEKR/UPbZ32zUpsZy+keykO0TcV/dm+I2DQHqPReJB65DJhyCTaZD8y7dbk84k
j95YUncsFpxgHbeOpgjG5o3xYrLaPpbaFESo1bGob+EVNSpAoCyw2VYcNOxhgl7zDvYv1nGw9iD+
DL9yzUJs868j9TQsyOJHQCZm4pNlTfMgHRgO4QQPycgnsmP81T7vfEFTxn4bUaUb7+sVsp3IllIG
UI1i4BlsHfu1j+9/2gJDif12DpSGYMWBOUuM/uSqvzJV1LFeNrOqqj3Zy2mObEyGTb+h703ntzff
If2EzU7Svo/uilYoEu1vV9+VfpzPL1kq8W8miGpNAiNUMDZwS3NKdPio91CRFJiOjcoqF7wSlYMF
P7p3ODC8jo+2Pn+i2U1qjivWKPaj6hfW+WFIatxDxgCa0DpPaM4IO9UAvuNIH7cVtw7WNx6c0C36
USzULFRXSMYU1pVVChqEWRHhwykI83aQKuV1MT8Q3C8UtWFgjT6WFoRvPNgcLFq6U2WihWxBUFso
lAiM4llVpvHaqlGc00NJNfxPS/ZUcM15RJ5S31MBWWXV8z6vsfJRCG0NuWqdt1tO/8sxXRiOSfGx
Frnh59AdewiwcEwRjzP6ZRrEmvR4Cx8oGwq49RmDuEnCfF3ZyPpl9bJR4TNDsVi4uyt7eRK4DNjj
LQ1KFejD3r0mBNtbITDUcYEEgf6HqqAhGXmGkM1/Vjjkz4wSTxziD7yxY82xLSveR0foY8x8vXfe
L43Dz/h1HWhTza+gqcnn1u8fAvOB1WBV/8xn4/rVv+3HS81vPivm19loJXw5FvnlBTABUG4EOKMj
ULlqYaAHWAL1Ge9s5M5mWfoRBl2iKF2QBfHRLeiZoZ9rq9cZ/vq1SS9K7qUP/FqyNZAXIrwS/0u3
syGNid0HwMe6o+R/Nyvcg298TAOcCvsbl1YvKN5DJdY81Ch2TUwtdxHWZHjo8W+NsYT9GvpdBC1o
X+xZDp8zT8TRcq0PTfwt3sVKYHI8macT6Eb0BMMspuCNkhdopgnLxJg0zobLw/Kcq7N9B+XqT1Sq
fNaf7FnsW0mlsYO+vs7ZDQkxdPtnmV8xX7/JDJrmOln9uH3GkbJEblZ4+TeWkZHXI+kVLHzrXGCj
dWR17R/2iJLjN267GBfOwVtPR1zKr1VDUSomGKZWzv3kbwQu1M3vuuxQPq+D8nbdZSEI7rro2AfD
BSDYHT+WbE03b/8v0ccj84Mn0xnvDTTx5Lqk00Hxt1h3gR6dLZMDLoCVhVqgyd1uhb8F1VDn/BXE
pqPxkkBacsCUW3X/wG5Rq3Lsp0y9+RhzWdOUk7qnY1pUJDQWwh3U1dIdbN8+QscCFufkwDhnu52y
MnCSIJqAdPzgJI3rSTCh+x1xb6wWvSynW4aoIRL/mC5DiGZ69uoNQiwYkX6TQCb6EpYGflnm+gpb
YpwbQzSNf8o+dw0Rxd64qOYW1MNB4uWUPxMnBwiheS12CySm3szn+vOHy6+RFhwu+dFykvTuA27A
OFx1TkiBWU35kr11TBheQDsxHxJ3NimeyewT//fdUhoIwpdsL4JsVrtRJwOeGGMAtu2GHNewbIfW
St0jPTtO5HOddnmVoMDGWoK+wjknvNYr7emWCIUdlNCiP7SDO/vYv2tVyNpOTmlu/c0XMNM6ccDw
eplHu5ZEaCnGgy0oXoetlZ4IHWbn9SI+YARl9PjlhHKoV8c45oym74D0O6aAkmIAG9U4VxCXXG8Y
wMlcFGc1rYtKU7JdCeLw84LlgZqFmWr20e7fXu7Ex5P7Od6RdsEcZ/U0ltOQJdMwTC8/MipUZoF+
114WAOaC97t8Wzkyq5DKWBM0fvTRHTPJEpkZN7szMI23lhuk1GTSfNXjBks8tJYh21jMoSfum4YV
otHJB8CbAPvElJ9mr2YGIidxrqbaJsDK55YZXCKViaLOkRfRYxJyj+ujt3a9vgKVU0dThdw8tzTw
VNpMEDXZ3BtVvM9bcywtHecv4fizjtweCWwOAPkFnE1odje7nEd4UFvPdIttKXt0ykE5U2yvRqPo
/yiaT/zCnEecIMlybOiJG7hjKdARxFvucTdJ61Hf8IszNO3Ttjv0QAUST/jhajEeAWUs12MQadga
ahNaDENwjbYpO0GzJ3mnip7wOEdWUVfV7L0J42ed7urrhrwShaKtIrKG8Y1D+PWgREm23vtaz+Ez
q5qrjMUTiDvJw0lqg4pbpaA9vwX951juC7s7fWibi/AvwJLyLlymFwegaIQ48+U2vftORIZrEAtP
DSPgPi3MngKj3wCe6WhaWxILZY+25/MLw90V9tFU88yE0IH6KezYikpZfda5qZ7PUGfmcS3ZDN98
oTYXa2XdiNwB96+tL/zfAUQYcXXhjVL5qvVGJk8yHYSTbvFrvi3STT/AsQWV4gs2Pyzxfe/sHVt9
5BqseU5VTJxWMGP7cBPG4m4hXLd8tfrYgMH3MIFhH9LM9jlTJfc3dHjb4doPo63gxeCUEiHjt6wo
iAnkGGeJhMPEwB/Z7NPkngTw9VeF9Sc2muKf+gGIS8kiAzzBKrnIT9Zuk7vkt2CS4pWF8sP5n5bg
hiysmBycBBqACASlX3Qk/HDM9d5YqCWjlZUTj/tQUiJVLbZ4/f+WIRj44RIbFdUniw6/CI5ChgHA
2vDFpEzNx849IDrSYk3xRg6Ius/3gh9UJ16fsuMIuOGCxqZzduGdIReHFo3V/qLSoWLWtEZ2qMwP
XvFAAGBtI/ml+5q3VdqWdMj0GzwnVna/WRJ50/izw05cdNRdRH4gJ16HIMw9PKm/FyQCX6ICX93N
oTlGCQL531U5vOvqemNzVDR9x7NlVeGeJns80CXXYTS2aEqR59HMrixl67FQdZfsHijbHGva1IOQ
0CLvC+y1Iqb+McEdSGLJ3oaS8XoPhBx38RzUmn+vm7nscUSk/fbvklVVYyp9PzQXHAuCr6Irj58l
jhQm648RKxmrjakGCL2TajZyrG7u6ebBqJkFtX6ZNk9ZMD6YMufSZZaQO9ycABP71d7ACvSJ4/PK
Say6W/9CfvueNm/8wIDaDdx3twghcYldfMzqEZBpO8Xcn4E/OUWlBSSUoCsk76ogw901mu3TIeUi
SbSj9Ofz39VOrnDHjhEJUjZRhNYQ36K/+vj8cZPha2NjV+1ZX5D8dmCXe7FmazfQVPzbnzBQajmA
LpmA7+zV8vXkp3X8/UjCor4OV6imAdZc9LgZGXsKHsAuZzaCJzbG92I00gNlglQSNNjTFJ0OiuQK
fI92bIIyi/yIik6HOMqWtaGafvHWIyuKTbSrcvMMexSqB4+uqNOZlcPogvSXN0DTFkD6r8BtVydb
V2oCNApgWxEnk0RhqCmUkGsWXgxNDLrOAJOHRNhcxvMd2cFw4GzmiCXPAAaQLmyMIOFXV9UxxIHl
+vX0ccqH7KiwzuXCFTaAUsNrQsh+Wm17sr4b1azpVDWBxnLtXxXaLZWo3DE6yD7UpQvwBipp6Lvr
+44ZbSazUHsdktKZpn24Bp4FcG1kf9v1yx2MDrnLLt9GPc/QU2XgHd888CxB+F0gyBEQYdwXar6v
0jr2BFhh+l72icVt5ICE0JAa82MeHtUXAVyAPbFQOROar8lped6L4Cp+SeHNElDob44B7ZEURq0R
IMFlZt6NmFxTPCmfsfURh4n6ij9yP9BxPn/HCQCk3MXDY/8lqzp+erUoGhLycNd1gQeiFgZOswoI
d07JC5uGuYCy2rjyZz33ut4Y5n5NsMfQbeIcuKPpRU6Z2BwsVepwe97d42DMvqOlZYIwgOuKfauM
GjDpkJ64JfbdRxE1k1PMxE7tMq/UycH5l/fyt18Vz9PE5+lvEVthSkEahecVG9r8Wf4oK4ut3PR2
lbh+73Fmj8tgbH1VFvrhUasaBnL/DDx9yKL8BbH0ILMt9gapavhSaggc6RmMrqzWwbOPfSg9dCev
N/K63NgLdStt/fKgku51WKAwKCBHgTne6ymjmqRXluR2v6YfcdvnyXZtL/f/Je+pEVX4lbGZsunN
NmprrPpMNHanJ8wfAwKuHokRQCxpZxjr8R1CzPyf3b6q5iBMRQ/CF8c6ae3SoFHq1+5ue/7aqDk6
3O/O2A8xOsSgMgkiagKfTK5QZhjkUQL7ZokTGAr8+XOUmyX92vdciU4GIf+ejDR0Nv09fZonlGXH
wSUwhSTbOA0brLJ49Q0OgU9Qttfl8N/Sd6Kf+E1Ji2Ky0/GppyOrPLjXxF1PaA6+ri536TVg1fT6
LHqYY2X3KSPYUTcpclJrc7t0HlgkepKIzEbvaIghZxsh122XDmYhZS1ySJqQuOwOLgJqROUVC3k+
LV/ObnMLDAxrmUx7RfAVglJdDqtSQY8WPbjoFC6WPqvkQ+kh0R8Y0ugnlyTzo78RkdrTsphkzKsW
/51h0o255oW9uEwg0sKVyhtM2BOMnBHIkXNDGZ6/Ign12md6fgS1ZSAy8k3Jd5gbyzE+vYGP7ey3
LDptwNY65TtT2RwNUBPIGdQKv6PEJNLX0zA1gP+67ofMOqZBRDPcgi5yL5noIr8/2VDpX8zDjh30
Au6gkV/rMlW63v6z13QXOaYWfHEahdLyIWqSiF7FbM1Qisaq960KstYhdVYfd/irIr8PRRAfjeSE
TX7+NGMHDKIzHnfG41ZxArhAkNFSu+RufUbRBbJn85ojTZoRV3g+DaKbOno+9yRTyr7EhEItQJp/
yAAvSdW695or1RkRQjskOyWe3BwMpslH7WbmwtXqdH5fFLNjzrbtJWe7FHcgOjoxMT7p8GjIrNTr
GGXXO6AgPZ99Z5AfSTBfdP5PL75/vWmk9fYKLP3knGTxncEWCU9elcisytfax7biz7rDj4E8Gwj1
hJDsQJ1e5uZI+KGBHDfnknlexYz/q+JOu6gWT6FYMJDznGpV/PPgLdFechWIzPC5OMs7nVkhpnxs
k0eayqiITvfrE7jD5WHDbaCgP+TN5MWy24UmApWUfBItHQVug6rsBfJgaaUqZ+s8xHyLYQVNH6pT
wviPYPwpFyiaXKWUgzIYeAVajvRX+1nvzniR1DCq4EN/n+gpITg7o+DIbe3JtYXNXBwD+KyyC2au
l/Rl3KCHPHnw/BPck+mXgRVA8aqNTq5IXHm5lVdvYAktx5Hahkj6UWBRFZS1NBaXNh9ve8rLrwA1
kwWwvrCITxcNa/afgTa+FZ0jO0StuHhsSXT+dgyuj4aoqcyScumU5OyCi4cDmtbOFEJPt3c1q88V
28VvSj6RofMJsxhwviQQoEkPqsowr8rBfvhMNHTJ7tHlAJGvkKoxvW5/2TNbY0dKiDMx5Vs1/sCX
kODIwC7rik4YxrnqZksWk7GXaQPW3QZ3Z5wKqHgR34YV5My2JfejFVZYTwuAY5zaVvhQgKCUuMpZ
KjTmtQd1LAyhXyptHqKgFtQVglp6zERTUTtfvsBvkFWxMMUuAHy5GtBDuA+6i3yzCHzjO/+IKZ1g
OEdDvwldB2AEP1lWSK1p4RiLkflbv5UA/kpKVwuSywAMYZiyDtjSHPpdM/bLPNJKGsMY1+9tYL4o
NfJcvIj05lFYWTB1uXJ/nGqWyhJTNh7CHJIGOqjZs/rKO13ccC/lDH6LYrK/1sdLw2hhe2Nvv6kj
PURUZxLENTdMk7MJA5VOBiZJh+ynY+UqbI8jnyEshp5PRjAlRqKlfHS5WwbGY7AHcrZidp/i1eod
goD4DpVIDPb8MV6WqESR8hNFwMPIAPUT829rBkOJiclkHw5lCpdf7HOLhZ85gbL8WjFyJkKvs2nN
wZ0UVau7cIg9V2KtPEThhd4X9Na1qhoExFNrFugl/K7oyUv9OWwsYHLQSJRLavDnesMljY7B+r1X
yQmHD6qkks9wLFVFeiwVezVRDysLiZNCcAq7vJH3fRvn5V4QJz0nqexM5F28O5AqC+0idSX2L3ld
+mPulqbpOLUoeRVMnkdVqPCKANJlJIgfQKRNFcCsvndTAVWsUFmOR6LFeAb00RZA2tPfH9UwSjww
iG9KqZC80R/KCgsaLf1BGC5as00Ui/kstdt/P9c+K8o0NDLwdsURyuBRnD2W1gxK2biRLwVn5SlO
dM6xewD9sURWzbWzcT5SqzZPpQcGtrNVhRzeLtklzgLLMCdx7Lgb/WQBET1I1wZSoJtqX8OdfIEO
mHecvaZ1IukOs9qW34tCu5r7zy+Av3ifKX429UkU3My3DJcFbXy9GuCpUiBiOqDFzFzThHvOAT2X
nIOLP1Y2JRHY1wm0MESQD6oKkPBwMLPf/7gbTF32H7+YsodDnsY1mVugKr+/R9yn76GF/Z8bEOC/
pxbzDmKg+aVvtgiRfhmfAywwhXQbZYWXRCTCW16E712/emvyCdz/+3k+xjMmDMD1i0XEse28qmvk
kXWWEhSsVqoN24y5x4KdYroeV27/0rOcsjN53e2sF3560wzngOg9eaY+OLK1DFiNlsr2iQkBvUwp
9wWIgJAnjraK+QkUbHH5nJ1TgRGsk0CoN8TfFuwqlz0ss7YX4/f+KTV+UHgaQqPM5Sv/xsFOARFK
u2Am7pHUL8MbLdl1jHhPFMOg7epZmC1VXfCLfcFUX64aShazX4VFt/OiiQqp6DIskrKrKF7skNCD
X6qTCb3iFg7FWSXVPxwo7ExOGqFM2y24HhQhYR5mQzqM43vzOUsDAN+D5DI72t+L+C/1bGp5zYz5
Ip0sYoEPuvxJagDG/4jVgc+mU1ncJ0EZ5q8qXkeiTF5br9bDN5OEOrsAzvfI/9RNWXq1wD20Y5IS
g/qPUYF45UeD3EUg/VcX2RV6PKQ9oT1eBUPGTSG0IHeCw2r87494HqH0W+nGXpkhDYoXFYMAzD1g
908kNl1Y4dWRP3Rq+c6PCTiZPV1weslmPYJYSngNfMtt5DW5OTNMdAGXqIy+wPWsHqVvh676I6YX
kTzrGT2aaWzzEeMuqnre1wQcXkH3Bnrf8oK7x4AyBkeP9bVQbORi4lz+EvfOuCY8bFk5tgY3n3tO
bQTzUgW0YScWyQz7+8lioyrdaAXQ+wkpAibeghcTqs3vSI7xEYcNAN3jaPB7SYBqv8OAMwdnN/mV
ABWCjNIOjxA/Rnj5IoyjpE97xK4EFxuvmh5/ZMU3rzKawQtKGdEYnBl2E1YOqSfgBM20bkn4fvnQ
CtDHkyFvmegJJrRHOONJmumUq5yZW9ETRewbtc2oGH38s7qvYyyLv/aDaGw2kB1rEn+LXpYO2GpN
+h5PtFzEp7suosvZIEb/kfD0285ywLQFErEo3FVOYGbxliCp7/LFfiLlputs4jyty3hyvPX+yi0k
X6Gw2Mgm0F/NcT9aknqxMpYX9lPoz1ZqGGNB5nxMOVEZXQ9goC7/e1OCHG4u5DDYT6v/fnTBwmhk
ul/iHfuQujDrbjHPFQUUNpuZr8jltKvqtVUWUi5sAolOiu/NYIvs8qzrRpHtSPSw1N1dq9n7EEhD
j2chYj3gZW4NQ2VLNEP0jLdZVhCQELz2CCbTPlFXS7bpZUowofSZnvv7V2+7QqW/hjlyzbBwiwTC
aMxjQ4KPka3ZpfcNk3XsEpXcF+g21bSgNReRFWoOOVxH2t7p8KFWJbSJYTQuEoZTlNnvClRCVktT
5rQRHpYiryEORcTE32HlJKE+iiQrx2YCtTvxHyYOKhyhJoeV2I+6kQidGr+N5dgTExkBYxN8Ug0H
kbHmu18zd6hSOTEC1Zo8TocI169Hue5Er1kYgBzvYRM/yEg4wyBJDsElTNzICYWieMVT42nyXGp/
9IFrIrhMru0K/XRFoGw6CqVi4ZP3QauLIHb9o7AvnTx/9jDoQT4LayIUug5WPlq7i//t6vzZZU6N
23VIWD2yvF9KyZcKlGe3SQQcZc3ow9U0Vdmbg6/vs586hlsQ4LgvUYotpfcsUJdv5vLz2Z96wtfm
JoDYM/7bOjTgUxchsESqPvNtYzvivy5BJgBk0Cqj6EAAy2lZbZrndXjePriYqM794yeq+Z5Flfp9
kCrKcIMQOvrujhCoutpwSY41wDFSMIdFIZiMIMYctY0ZaoT6/k33hT6QlTOHYRm2GCbTqh+oJ62V
/2SQENJoUzN8ctGyrr+zCYOIsqnANUGe74BC592aVFgGG5qyCy6ayQ7K1XJGrV6m2ws05nOsc+6F
gzPpf50T/OFblnafgR39JWlikupZgq59mVciO0/dICBA/fwVJZx6pkHjBosIOf+C0Z8DONEc+wIf
Lmm548jtYkTjq6Z/u7ewdJpo//fUZlxssudAQsW7XS7Sg9mxsB9BtMmUHJijk6T8UqmAR1B2RBcB
m+mCq1tzLKswkZ3Q9JB2ieY0v/1izSTM0cARJ79Jd6HUDvAE4nXUwwbgTa7a/YtV6j0oMOiNSDKA
EA4ktKkN7waqQ+vzlr/7UNrf/vl9wIMf6pWd4D8R2czR4WR26Gu40Sr8zjzKjXFyYIKvJE1c2wa3
M1wUxKKlOtISUGDzk6TD1tTqPXz5oWiYi1uNa5AyVRefv47HRERVlWG3ft8x26IanzK4u5j7TQl3
+wEeYvVuLZvI5ZnjWKJHm737G4MqTF+W3bHLurq24JujDoktWVgDdDbUY69HWR4lwCIZii0stHix
QsqMjf+KterUJZqUSbTRaQmB4vfkZhT3iCA0Lk+OrRIyn9FLrS25SwNJl5XSEYxDq4F5sm2mUl9J
btQp+p6HWbn5+HciubhwCimrMf6GJUTsLQPPPaaoShab45SKvzod2j5KyObfrvOJhx9nUq81A+1a
H3ADxt1MFZk1C4TxG9N3qbIkBC6graa44+yITrj+RbjunAUHJExz2IArZgY6y+iepCjnX1icOV4f
rBuvu44bwbI3mrZ2PzYLhujd13lwKANLizcsrD9Gh8ucf8Ami97uLQqc8OjeMfawg0WTmzyuNHqG
kWR0CVgYsXSwJHLM+029uHneefvR2Nf1jwZy/n12qcmJMJdM2vkbRTijEevZg+kZVnMym66LHXy2
e+KMglRoETQ0BybJtivKZIDW6trFVa2bEreDiAQzQd1PoAS8QtY4A8Ftl5Of87SMwqiD3SGGT8KJ
qtWRLlI9uap4GEq2W4/QHEm7NySK8kKNzGOxAvmwnxIuTA9UOHvGmHCJosbJhrv3i9S5of5BiKr/
tspwDCv5HnrNblF1kmpLFtfhmRLg5P+syRdv5wmCyowIPgy8jm4jgHBjszpWa0hwHh3r0lBhblFE
1RHAkBIIuUg0ydKBdO1gpElvxstS4Pjrf4r3aSA25fagFGxsTuiXi6QZamSytLy85fIMiwJtPl/E
o/6MjwP6TfOwdxnSACnlxo0z/QJN/NU/6UM98tFJF40zixE9Dn15efh57HqzhhjfVOraI8rRm4XL
5AACraM1LThqx2d0AS+AIpohp0L0VIEHplFNPTjZwpBtunT3tQ6kgX7FSAgS/NDicZDXFb2y+XOT
SW9X+bwrP6+hmIE1bO7hnrJKGShwPloKN7uY790Y5HAYlM880OQkd4eff/fkqNmMRZNmvTXA6Gme
6ByztCh7M8F9mQpvC2cPlfvmQGXvAo3YKOwvI5QtWMGDIWlCKwcT8nnf+GMbmqt08xX5bWkkZNKY
v0AysdhptBUzfmMSmPsY9hTbeuUFqLHhF5ITHgsswvs2uhbqf7F5Sngl2jOb6Gq+PGQp+bq7m90W
gYPmPfhw8iKflR+bQG88ExhqcnMR6lV95IFXqLq6VWtqSujFkO3IcWrDXQzMm4V5opPFO77HRwQb
2lg51t+/hWIrryKT2/VcQhhm5axUSq30SLIrx5ZuWA0Cbw4VL6UNDROrbC247Z5/ljZ8t0VPYnD8
FOlA8UfEZvSGMCzSfnT6y6+Jc/HA9V0N2giVkJMEgxXsGHWcwI/G5KBzMF5Bu05PiUaQbpq1+AFu
BbsQVVybMttPIL78FnIIHbIKMYwAo6It/ff7b6v7569fkMy4eM26MDXChRq1xDAWUe/rvS5ZJOvw
2w6XRLDIeTToOcMVT8uWRB1ZAlxtZA7iF1VCtMhWiWybjFDtGMar83KdbzBOMujZVMqCmiiQrsWc
U2H050FQmfar+mOwrqS17ViMoK6a5xVvkP8lUT7h8Hh2VUejNPp1+Sy3fTgJp/Og25ElCLTd8ssN
ar3qe6K9KfLzsVonjMIxN4HkUSyrHGtt5Z6Y2bP5DBTXnPC3czzzDpZM7sk7bMyggDHKDKnRQ2aR
dBzvtLMZpAzUJ7fIO6wT4iRSHWSFVHEwgXnTltxyA9FxT6GYJMziIKs9LAXIX6ja/cDBJCXHkERl
UTXrLm4huluXz1pib5ymrwUqzwR61bkGOMuV6IRkVrfKWIvpKvQqhkKNgBM7gX722vh1AVbY1NEA
bams6c6SzTRM5qJLR/xhwcISOq9kXmU4YqQjiyX0vrJTORoojTBzK6p+B+CN3waA0qAtQR4NlGSN
bPdhTIZ+pMDVPVhJQfOhMxFhWKCGs7yDwu0daDJ4onr7+6VJUJ20nYU79gUMcO8KHoWnKr+0ht7E
JIdeKbr09yKjksG+P0nQ2PnagvZpmV9+XX7NIQmI99iku/Q9oR0PPj+MXSepYQLHaSn5BsCgreDL
jIu8QsE6IgAHylvURz3kq/5aHHRhYXgx3crpQJNGpdXvZAPze+RWR0ry5FBKcENeeR5BtieLuS6h
2uF2Xt05T6gJbRrxxUeDugPZf5JINUAUJdyeuU/OxH7NTj6ZS8KTOfLPbkCyjNwmQtgzFHtPpqbC
Osq7xEdfuMC6CmRSwLEkBOdjOEULsD/+EqbCVPpG/NdbZtMt9wFpknSukFVaFqz/ld7+CxkxssTN
s+ABCPjXcNt40rjquv2beAXXv27ByiYEXHhO4IDhxnmXlcwX443O7K91fvPP9ov/pLJsBAG1DRPl
ljwxKYa0ceIrm5hRqFdjrwqbb2CXQnU65h3LGtb20zhkmA9FjELigoaXs+lSavgYfghnRc1yUaQC
dEhmXVXZWEXI5vu+JUW6K7pKkvWyCYBOxG6eL5jGAcGzDjMpyXN2idyJMDk28URKW/YgTpukyDx/
fb0y7ZFK3QqYASQxeriNDPqcMpuh2gGfN1XEXEeGOoYhmR191FPvpZeqdqFaWNqQuq0Hll3qZl6g
o57vQaWelnayR4saiMo3alLTNh/aq3KzBuUmJDO76WilQhr2OB20Kcv30bhsDgFj5bfrH35qJm8U
Zh/ZjpJs0Hmewi5Gmg6DTGhfqgaOkf+bkEHNWbCpRkfoWL0zdi6qNsHE9A4EOM7LJv7iIkXCwG5y
mjsf2RU6V9oMrByNCLHfz5kl2VLMV9xXehxnvXD+/RCL6M9jjeq5oqVIiRCwbXkYSSiqc18zTyy/
AdX52FiRfXp3b+05gwUe+KzSwRMib5OKWr03lO0Vwygo4cRJXL5AbleXna5/35X991VViJnrbIN6
HvhO9nJDes3HcpKN2qAXosnEaAyGsN0hng70b8V8Jq5cyhin6B2S1YCaMT0yhfQVTLjD8W2xVQGt
BujqVnOYWYjPmCEjr4Q/oxLkxnvP9qbyuUh41mUo93IBJxTVed32n0L5qcybQGISgW/n7c5ImX9n
ow/KVcuN0wZJTP7epX7FuqY4gDJgGPyoKuWMh3FgkpHvPp3OZq8r9mkuw/I/pTJkcb5taKXtoDz2
AjGrG/tog518cMf8u9bnMn4BHpgPSDUQrE6fRTldCMmrcjW90Rbq6KtkE/wwfxW6+c7yX/KkzdHX
ftH2bE+6xW94Lc6AACX08bT25z7tIcozDKF93guRbL03Jj1JrOB4R+vy+DuRyKP7iMQ00d3UIA6D
BGPMB6T6xIAW3XbAYTBb6hK0xJE82ze6G6srfz0Brx11AWc8Bm3mccIxwHaEafW/HfMzHFdNKBgM
on2T7DPRc9rZZ1OivvQwyC070/Ty9zJR2gNlj7wGYnrvAKynlllxCzRSDwSjIsjMR10Tnks9uG1a
ms9srw6ReqfA5/2KfhbT3NlZ5+xvRHDHjIrtFaVmyiRmHbMvc/n8SV3F+hB/ttvqZGt3DjXG6xJ5
oVb9B3y45fjqq78zJeDwkKiqFwPuSvBeh5znPMUr/6O34qzYFMs2HkwzWwQ0cR0W9UI4aT55SOQR
2r6LmFhVa5E6vxvroAyx4Jm/5ika9Ea9kEVDvkFpRIcoxXbbL2td9dlIPaWnGANMdoiVaiVcvKIH
eVlm21jSRcHJgJvybwuYGifxUAgj4to5q2m9Ycmuzub0qXyk6mEPNaUwoAFhUo2s3ClGVJAq1fot
9l997hpg48pyMi2HuAfXoz3q8kfcNVd1r/071BI+SMeSVNYShSLYXna7hk09aiewqVlZWpUT3FRp
Whfl8Fpb+sHRAnmi6JM99LDbFZEKO9nrkbpMvWSb6uYRaPggLgxKVANmJLFcniiVKUqpF001N8dl
5v6QHNhgOUo3wC72NgcrFJLRFD1sB5EsjVunt8dq7AeAGABhC7NN9ZMo+KE2uVCA+kZTwJ2JBJ7l
8Gg5OIleLqy1XDFb5r8xLWTGQKdBx9a1oprkp8ZNQPfYmxOTl8tAyyc8enw2DM0lUxNps9MfaThw
HBpwcXdxBzhGLIo68hDvpo5OW+w5zzYKuRPJgQwmj8FxygAS6MFBAKMuT7fPqrPHqk/49ugdmRu+
mWdO0UpIMSs7Xo67FyaF+6UqtHL2W1BXQO+SAXVv
`protect end_protected
