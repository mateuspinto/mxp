`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 69072)
`protect data_block
FjufzIFmRiHKcllQAtqGLR92fqkiegrLYdHbE3c836vCC34+qAlT+SeBChFaGD3y1iwQn5FvITJK
vfVktvO6hQcc98SmSUW7UlEeGLojFI90a+1QNdoz+7XYzO5JPNQDg3HkeD/PyvHYMz09ov8+DO4J
4hMX9ZeGbYNVha+FQJT/vKRDwYih7Di7eB0hAm017GX1jG8M1TiUXU/MQKN8SWS+ki0j8Vg2be/g
tp7VHdWVy3zG61maU+8l5YG4TghSxTLXXYcF4L65RlXGfQkDA9j91qBIPCHK3V+MuSgi+FThBAf/
3d2xoBGITdV35IEdOF3XPSaMlcZUQsseiO3131aq0atiws5IUYyxubZe8KDtZZ8t+xf3a0Hk4bZS
Y22SLKyKPuapiiHaNXH5MKy8OJkeHIkswmzFphpxFBw0pA0ATN1tQQyCg/nJRbR6J1omQBUYWQou
LrIOcxZPT3NMd/7Hxh9RXYaPeP/groyPn2bvnsHsWhYN0gF8wHSF09BRGjMrFxOW8eO0p5wT1wBo
ffNhb9nEsdfB/u3l8TJUL8j3ssBSVsQSuVItC57MNcct3ne4J9fw3GDTrnkwKgK2+c+ZioFytTPG
wuIckuhHJoFTj76qt7ZLgoYA5nkkwNfdgVSBQzgexcg1zmK7vBVOi/PhYqzWEjwvDmAKQIMhH9mM
vAdLxTvIGkxWwQlyh/WLVx77Y26+UnX5aHPfDsJDZqteI6dVVi7gMltcRWsgV4HHIgRDe/d09ulU
3G9C3RjsAWiWQgjzH9iR7SaVSouTUAvbg9hCk98QaZVGMTY++cbIH0P+4mq+unFDUaIgaqGoxSQ+
yyOnko2+40mGZ9P1Eh+pmUOH0HIy0eskjpqPcX9ipwmJ6tqYbeHuypqLxLrycVLDEb55FFCYzyVo
SoWrYMY4gJhuS58SncRLlRYURaMGGgeaPbPm9vCe7wCo75KDD/buHFGotocJh1kTJxr9SC3QWy4k
qb259GiEVB1eWbtM9PNGun4novfDI09xSkMw5xtTYXDWKPOVZiaZ2+yX8DciDEJLjAb77zfdrhOq
URO7YKqyjKm4Dy04hrUlN28amYHBRhtiBmEy6i59Nt2fZmWEKRxZS8qm/id6Ax0BoQn0QBYaYdVS
r3h66jHtFzAYFGaXkANnPQ6ma/M9T1xjPO4krUccpmDcKNj164HhwXWX8v13sY7DAe1N7dlDB/ho
3kY7J4Z577iOkHxAf1kDKqz4vo6yo0RlIpBMu29Mn1lR2HUkMbBYcgk01LxiVlJL9QvK7wqUrCJZ
AfUMCwhih35VuP2GXp2xZrCdnO/p9Wdr6XIQwuxncc9JzF8anksxqql/P0MDINMfdRzfe4dPpHMb
xkZ1DFyGs/EWhypAC1w2Q+7zXmkhwyzQ5/iu1AD8kmFdE7vJfzGgC1b1VYzXNoZjKspBbWustG8i
weSAUK96t2BpybRa6SD8oqOtJps218RhZ2vqjg1UHTn2CWFbpnuiCPrWGeP/rj2OYCaJk2M4DHe/
of4RtusId6p7poz87hF6WXsxMYtzym+Gy9cDJ9CQjLnYOAM3JyTQDU6yWeURV2qI+DN4/h5tgx8e
jFrXGHTK+qmLXEoZsIyhb2FYK0w6bvze+Pt4zBMhtRcxkDnrJ9XVyBa02CPv5jokXq3252Qf7vnR
MF7sVwsRBu54LyZX6Ck1v/rJn9DYT6pYVV7kFE1q2ls2dYPp7w/regH89MCFq/mAgsikRxsF0Vpt
5wpUH2gNgO3rbGlQ4L0EnPJhYB1wG9N4zbSv0x2wnkQs+P1ykWVaEqI7HFYfKdvZUaAzPn5t7ZvN
2o3o+4Bkd0+eAwsNuFXCLmo7BUXHIAgj1kKQ1KmCA8HIREbvCtHNgas5VnWo7MpdGf+1E5wcTiVp
a5dss9JmSxm5YB26Z2KVEqh94eSY/5RW23AtP4r0nteM57dLdJYpGZGEIbyS48E/TR9cQueSuFod
k9L6tPhKZMuI8SK1y9NQg4Egk7txoT7LfTeZw4NdeKwsVHqDh9Roh9OUVEKqerVe6m2tooBHS5rJ
18d7SlvVZ1mMKTUVxGioaHzDh+s9f1hlf7t4GZDJdFtQANCjioN4hmr8o9Th8nKyz6N86QOs07Tb
8nGx18fZK21vnNgwiHctKMTEy9VhqKJJB87G4hnW5txcPPW4ZvN4NYeBGp4PLcd2NSZBTDPvTbyI
WJoPsAO6dd7sb1q0O5XDNuRIpfw+S0K4yZoM7WZCPbVXx8764fmN9dkZcZC9DwbSstnqlwkAOxmB
yq0gj2kbv7XWDXzozgnZvA/AR51iwOpLjTwygSysl/eRGZD7+oqONz1ykAbL5CFC/512kT9rc+OU
jaOUamAPqQ0KVoZwRd3AltPetM8Vo6tRBG3Ao+OcgSkksroDJu0RPyu4iCJ4k9CSAjkpF6IirFP3
kj4mo9R/dcqkfFKpxf4y0TPe6k1vv3gtiL8/keYohbfC7Pit+Et3qRjdgfM3qJuvRsXK5+DY4AGY
O3CAXzzbw57oao3hgNFHMx+yIPZHnMWTPcIXompykPiqiObP4hFs1GMnZrWP24BDt6RuFmAVcbFe
DXjqzeM9/zSJyffXdYZJC60CQfEb17JAhq1y2gnCivvWyVcVUz8rnsD4j3xFINYT9XwVpsul+mQ7
ueQ+5kPjHLZVFAphAwU4MNK3YdW8MCBCudSIBUC9iuW+0cZZOYXFPx4WimClS6RX9cvwhi/C1Syt
hYjvGDhiNMCs42UzYcnpnqUqLAuA7qPktO3LlY/gTd+9c/iqBuwEhQcFT0C2gmtFRK3yKlBdFaQQ
/qiiDwIJ9zjJybm1EYZPP1u6+8QnYgMkq2syCGqLYaD8eZ8awiwBx1q0/jzjQckb1XOmQNEQIP//
YYEyGIyLoiAmR8Uy9oiEUCG+SESaNX8BMva2d22j/mlyfPPm4iiGofa6XimAE3oVYTp08Z6Oajkn
fhrr3jaLgtP0m/Ox0QmbPFWq+9G4+HAvZwseRffafY+mzNwM7XXWOIo2Tskym6075a7ENGqACV1K
yJaxPZpyhvlQRMpq8b9bC8GbB3xYCTrdRVAsQJyrvKa3Agr9NF726SDO4bWQJmnrc1Rhg+slRaAH
QfwSKjtwq3wB8ePvIN0/M6221oXK7/dAQDqQz01dCNMA7O1sXrzjWbP/Dl2PnUauEZgK8MXwEgkj
5fqEMqPhu3KEU5O5p1OtOHg2hcjenjn5PoTfmPMfRYVVh4uci6QqcFvMC5Nn7nhif/ITTG6HXQK2
kxXuQOvT9PiHKgxPJVAz7CfKN3E3QMb0lbBpC8bDrkD2U95DbEsfhXm8DaTu2D/WPYDBuzszaIie
1y/BEMjcNjzzwxFd0OgwQMgAuq27csjiCoyGxS/x/ai2ZOFLatsav6mACL4GdzG6pq0y3wzVPaIx
yXMRMQfO3mP2+h+fdMTJgf0NJ8GN/BsrVcBKXbXxagTuDbR9JvwODXFwuLOH9U7gYClAN2s/TlsS
+gMObtRqZMqXhZ9dBJEgm+hQEFde8667hWjuzpF17rvrzDgCceiz227AJ2YxZeNq6Ishjq+JdFlI
K0v9h2wWuajggdJx2QuGcwnIyXBdP4SRPwLDOrXgkbpHtYt5ygfIvYaRu3Woldhx637J6atgVIMX
6lqohg4lREfsqdHtmObCg73KEG9UkAzC9BaW2mXj+6VGKxuOwLIfiU8uIKGxKs0wS0PuQHRD2++C
ZkZKAdkDicUUi8sEbIFeEw4ddhHb8FCph8wGzx2+0ok5dYEtPV3+1SJ71/XDvxdIcONwL5LqFo4A
3T1XhYEzM2qJMYW++3oHBeyhrx+9Pm702bUZiojnONM4c0+NH9CWwa+oZy+5VbcWjfZ1dcZGD/B/
qGtIwzmMP02Y3B1OwbxfQDJArAvI6HD4CKyCFnBAIwrRrhDLPGDHvSO27WdtDoLYnbmHw+Vk+S9j
QbgOqNb1/d/lleh08Iv2/gmMFip/KT/TgIs1Dok/mkviEVxfUp/UwbTr2h74mCQY1jEpImywjiba
+zRMrZhOrypQncXJqORGgZ+u7RIni0vRUg4xnDir+wqMH/C03hMw/nEM4A+9fKB9cwvoEpynOmrQ
JmA+oJxJebUTpdeK0cFtzt1UPdCP0FPQkgkcN0k3ywtYANmZvPIorSp8Y+fZAX3YiVf99aaUWmYh
f4CBGP+4vhM70QvWBSb10I6iKj+Iy2pwFy2MAmsXEcA+PsEKXG4+LtK/ALY3BFFfoYHfrFtZzf3a
9ajlMnbZUfY1ym39WaqIVTduwuyRS4lsBZ5SnkiHTYL8gTU44yWXTVhUC34xVW89sb4vSEhSkt9M
zYblDWPZ/uRyfzPjw4V611O0v2wtnf23vVzQjEXsQW3cz1/k2gfl/BSLub88N6hqHvR+tH9XF9fC
ufyFH3ccGqqYA2DBh+uF0nHtUKp0MmFP9n+enL4tUCLt7ELqoCFJk1y3B8TGTFHduM5YbrDEisD3
4k3mQFdLgvSYTHW8wLaiuN4+7j78HSxcuJMiTCamN4sUvOUz888y5rvB2b6l8+9CzQhawrTPG7TR
FQlA13BLDRXGl/PbXFVR0/NCtL0ZvMoAK1yyO3OACaEhj/o8Ez9bjt563ZTsmqez4hgMIGchEvPY
lFKoCXhS017vMdItkdmqKCyBdxbkaTSaclj9OdxmlldVI1+WKwiqmKVLCjRu8ZAUdIJaOjfnmUFi
UaUKkIoN99FhHc37TzBBLH3WGCvd+6OZ+DTcdTizDkXWPcjOMngH7YMR+8YzrnUo5bAWVV6XSx/G
Db9pwy6wz/0vPyNx2NDFO1T/1UZSF7XhkDNfPPko4EYClF9h2wSA/31TR/ctoK8dhAF1ZVQypnRC
q08Sgyowfj/ogBS9lyTUanvsXQbicDWi67z0m9YUgkpQN8WaoVeHmVF47sMMiDH48YjgijOXFXR8
JohDV8DTp+ZXgKaeWIXfLpLuvykXyUYHFpdMlxGaVcK9Sb7BER3U798c/gpot7WR3j0JvtWUCplM
OKE9LjIu3BtTzNwrZU7PcPleCB50kDGgAmVnAG6OX7hHYjrO78B/TIFtsZddOF6G0RmCFLCQKLX3
4F5X3+9GmdRmmdSU6kx48ZUa3fe5FJauLqTcSbDoc9LyhRERviT1iiDDZq43m1ssDoK9tsF682pe
Wn8Lt16E8h1aaGHEAvwK1vVGKTo0Na2FHEm4gRfWY8Sr03aH5a+oNbBtQOb3+j9pwPydATH25GQh
vb0kervaC0E+Xew141Bb78zRAjeme5dMaGLcKxlwJ0ZCtVSOSWjA38TxWbge05HBdfytUGNZDPwx
KCXDpgmfXU3kEPgm073X8XOVMBIZMrtK6+AESZzOr7Mq+/rZyf0+9d6TmGO3Bdzm3A7fFJUEWcoO
kLrxplYV5Xjf5bC43NRTO/V2AadKSgB8pSI9yul3XtSxLWe6an2oMyYl3vpiaGawvco/N5xEdjgH
KbQlmGowUjU6Q44fcpXkqGtUyX83VGP54AOWle5C8K3CLMCHh78T4DqGo2bZk7Bl3Aigth4gkj+y
h/yLFN12tZu7ZdT4rEeDHCqjBljzjSAcK70zFV1iVFEyCotJyKi/T7l07VVOLHwh4gW+moorgTXD
71lyutXuLs2Vfq7vcGHSGBNgNhqUWESWMXyBpYMv++mSwF5bnQxChnIAtFFd2vv0SsyK0Acu698A
hMKjWWoiAggHVLoBS9BE2LX/pDpoqhY9u0vQDsSYHJYhthhdTyagGxvIDkxk+tUO1wAvmlDoGE77
sWl+OgmxyCphbizXvyBx92wjRvfcQ2buTiAR5Xy+yLNZT7NGmsge5QM1HOLp+xafBaDWG8bwRMCK
l4S31Q0l2AA9gJGTUNG5VAZEYcZ1KbRVmJnyunKsGqwzRH5NCzk+gvBACARW90Vidjz5eQHrebLi
eK/Tg81f2M/nJUrRAM7WrnqHbEuJCBrBmmp+bYi9zPncASa8S6GEWE4wP5+TxBEaf0tZ+e+xvXbb
0kkRop4ChnHxe9zUSrvc8qZko4qao20JnL7tu3SfLdcngTO8rKguJKhpfx85OjHFNG3Oi6zn0Bhc
zoAi/rFzV7VKsq+/eCfMfj4roKgWqCrMgt50pvGPMn+XzEerJHVeKMo13NPJ7SRldtd/ps5Tjb76
C+LIhhYV+saexRdlbJS42NBhigG70YuRMdkRQuWCX8sIS3GZiqGIhBncvxWoecC1x8jvZ/1J5Pf+
W/nULe6gTfEqkzzffF72olYThkGLC/8NGx6pOFFIKYVWF2rH83G1gk7dvnKKa2Cr+bG3TBUbL+Vj
6qZ4wc9y55UnktIX5U51ebqeRivUVe9XoIqBCue0b7EZJoEvpf3nfyiYwzwDdHFERw3w8K8B/faw
YNjFf1kYKGyjIbQjH9fjL7ytUk/TKTHGESXt/8NwWHv2NqWywjs5VPv/LCcRbGPJnsO1b00wYFce
wG4ZS1wit1P4g7VPIiwboQ5xUIXRmeaLIUVL1GS2ZwRzIcaiNC2HkeVzcL6VYNAwPBZudhCW6GBc
9noBDktCNy6KylkEVXO4s8Bv6lHTis1rKS7oaYwC0gdxlsRC0HpKfg/JaT440c1vH+ySXyRs0bNg
NNsP/4eDZrFpePlQ/icBc86KXsQEWtyTovxd2olV1hxTm9oSX7km8wJzUlruAmcpWLQFptOEP82Z
qAkBvhp+48InYlvUxmoVMknEODgcZ/1xoCxbhAzAYuLIjTvb5xSBRxf5mSejMAuGjAwmrO6JpTZe
DYloZZaSqBzFqd3nO24ihmUkyIwM+nvCGbEXRzyCIjoYgsKnzycYLqPQs9mI17DFd6x7ilfmhm8D
hZFv7MXmpSWsRPsh4hOSCdIcqNoMQfONk1z/CXzzPKUlqbHefNLgzIw0S1KS8Gmc58n/hiqz7hEx
dMzdsrSgA66TPe4Bw3b7gWRIjcdms7aIKnyS12jBxZEY3WDqNqxd2/6suzD8DI1beQmWQms0vpVz
RJ7UmwcCT4PtCWKb28atEq4vcRjtJZ6SpuAqshlRzI85oWsc7fqpRnLkvfk7hK2TBzy9ad92UHPU
YLnV4PfJ1s45BUZCPCCp1D8v2t2FE5/tsyfv//YCv6he1kzRiez+Jm4q8ahAMNcenfppP0L1+Fwi
nx6QxJSjeGGouDGOUDyO2eSKgxlJZIZFJyXu7qyDgzMArMtAC29UIRwCX49UnFdYXUdU7JPe2wc2
1RphlL7nqESv1wVHFgxIh6HremxzI4AInlgX/qO1PPKmCt6xeNd0ws1FItseBUx75Mh5CNIU0u7w
pelJviJTvOUX7mAbftZ17TG1AR5+VVQ3fR3H9BAzoo9ShKm+dQH2Alu+RXJDzVzqRFCqVvcOAjr3
6/Qocicqor2h51DtsoTrn6fzL35F7LQQ4b692sfTp9SFQ9HBuqBTMe5ZnAPBwEN0UUwOMo8U0//6
7Ekpf7wNP3sh/cHbsF9/1Wt8L1y4KU9+6qV8mQmrlyR9IgrB3qTCgAQaDerPjgPBO9fDpQd8asDx
MVyzHdiyizGjnM90VmFUaijaydBf1kABEdYNGBASSnIArXO/H//WJawoz/4JbSYNuyx+bLF0BmS3
ue/CJ2+dB70PEeBPt/UUCMUfD+uabrAkDsIgdMWg/9KTqJYSBko1QUkbDKJS5vbzmIJ/MU2DpZyR
b8XOk7PISsmh7oKpUOTozBKP+IPCzehBK82dJBuCLfn7KhmNisJmQMII5no8NFUgAsrcbHyaxuYn
rBNHFvNNpDKRCbio4F53QHcU+QF7/pCTIGdwaG5MfWixMYsoh6JQbbM8kQ7zrIDXvqrGpiFbUgXg
Qt75WV269Eyx09soby//VCOVQ+XgaPwcd6rDq4O0dLx3eg/sCDopY2KcBVo7kA+H7PH/sN3Yx+t0
IIQ6kYkz6hwI/SXlGvdjhGjFa7QM/qaPt04c/Tt3OVeRF+CLLsk8BRjuYzmBet9jWoDh3MkLZypF
5Srpgqtl6ekLz8tt+TVITPwT0tL6EhR3cZuUsJc3KjwAvKX7fxmCcuuI/GhkyVHSSuDwjvkvBciX
iqTsUfAj1rziZ/FdYFg/ARFbH4tnO5nw7tMeMGs78fHIwaEsijNjhGO+sO5EXJq7FXVRjkhyzTse
dNKE6fBStWjuxWDOeAGaLDb5jOhe4C1R7Gf7Zy7RJJgON+BD6K/6n1x1p0uRd9OK5dcG9XQ/NZEw
cTIZ28j7eXD8bwKyyfum4VxNuumFjhZg6VlAXpei2jzxwsA17qPYYl579cVyZxImQmNEMiCkcJID
mwD8FCft4c3DR9OHHRqhQi5K3On/RsSw3UTHvCR68XZivb4Ya2+ddUnngAsDEW+wSx4l2/yayXCm
ZKj6+qULO35lWW4aVVzJv+7DSVDPU4Y8RMp1AwzhSpfFM/+w3y2b+sYXRCgnOJ1s+Xkih1SHzM/n
O+3Pbk3UaXHgldvSA2FYpJuTTlzyVGAK7dpcqek+8BtrsfgRYEGPI6X2s+nWi71SmrHRL6j/4KU/
CWexkswoO5wBW0tisUEEOwZGI2J4xGCiP18qgAlDIjGu18wyuKy3uW8ySFtJv3rPRvc1e9FeHEr3
8vlPIhohBi8rZlr0Rg+fMFA1cUJeSlMSc/JwyuaLaawg7k5QewOOJhWc5ONvVeTpyeL6bu0z23ao
U3H3sRPTThQx34uIPNQzfwZqVDjG15z3dmLLshS23TE0zvaE+b3hljqkNv4aMWJ5/r8x1FUiq7z1
lL2TBspRjapWW//aNj7Gj8u5vtCe+p1OR4DXYbxm8O/Zm+3oaXt5jJNe3VijDz4Q9oCENIXeQExV
ups5ojM8AFQ3JRZUCuRB8EVJbf2ehhWb9yTWVfdWVwJWt/YV61CE0A9LK1BmRuPtZo0ssaDkwOvN
HVfGCVTrkBT5k7BcEB4rufUUheWO4Ggg6lWLumi9Hwc6YxjY2/ivFKXyxApoEft8x4+XXJpxFECk
D9tBq1XJ8G7+/Z4Ab0hOjl5yQxltMwssntqOHPP3CkyxWNZtLGiu5YWk1z3NaMuOgBxpx55iSBRt
jlvXC0xwSCg+gKz+HulfX8zA9tGIlpxbVF8eyKDwjrx5VWyUZFWXVxW1VGRq6Us3gxPTxtBYm/wO
YPwBnxyNaGo3YiXqNtjcF/ExQa2aCxkyWDLnWbOD0hmNOc0JZfQlRKJj/6uvL2viImbHGQJKPTGB
ggqXczOvdWk+na0FSCI0+4ljiE20UcMGE3y+BYqr9Our7f5XCkbBLHp5eKWW3T6wWfzn8rMBXxME
SK2FREM02n2slWuqy8vqWB1AOvWubTSU8coPaMpUA94lRg3PFb0sD+KFwApe26qNPlJZvUNN5+tH
l5WpQt03qqH2Y/4VaWjDwwWuXOdQ/pjmDz9KB52b04HVDK5Ed2WA/Ax9lNXzHpjq5tdwTsGtTpqa
+Q6tTFO66xtgcIBXfH+YpESGj4mXO4bZeyUFN6tYGLfRwTG8OnIVz+hrK5avrxePWs82jhUJxSpU
yDC5OSxLxhDLBUO5r/J+iUD60cbkye+/SDHKl2r/7Sq26/3ruGFWTgteUxflnp62swST0vWPMZMI
b7A6COsiy8MkuUAVb3KPTygN2yIjaho/2i4D/i1qtNC3MV2AEFDCJg4w5WA9/FW/xU8NSPmhxG5R
E/JJPGWFqsjpRAJCRqKzu+v6QBD8dofGIBeCx/OFSm4+cn21ZBomE14t35Wpwm9MAZ24F6lMRsUo
CVZg8O+IeupW0aNNbDmN4NjwY7E1M32Vu8NiLNCUB27Lx855RKDwU5Fl86ckvDe/EEaW6NP3fsII
N8HYEzRR3EHKYKszvfJ2cENulDqB5e9zR+LfPd7dQ9LzUTSlBeTq/4N9gOLi8bDsieCO8RNgeaqc
ltNkU3vVFtFJWy4WkY/t+THFKPxCprno7YvrrUqJgEnrfpMLw5lGerfONxaBpBOUa8Z21WY9lP9v
nef3dHOwTBfu23ZjIiqjcTM+YonEyZnI0hVM7RDgv/U2snQODGYQgUIXRw1RWIZlDMJUPDj5q9RM
YbNEOiuAgNvUBfFdJ/jfh9pQ916UyUnU+IXxb/lD4glquvtXZHLgALPdjZ2G3yn0zc8MrT6XvU34
Oydt1cJ9GnLw0XwG/Q071YpR2Q4FzSSAhsmTHrYyBR6Q03sgmcKAEa9bWeIm8oCCvtn8yAtYPszW
eSp296wKqXQ5B7I/AMkt0tCOrLD6m4OTPiJLT/DNlzk9Ey0GPTJMqs5Ep3nRinecJGQSVOXPemN7
xdz+hqRSv6u3Eh9eSnVTwwS2vSP2czzYrjPl1Uz7u31s84aiNuIwfwEnOrWEDFaVo/ST+xRomKHD
YRbMMc6eN0JGRt4LCznAyGfvKuVvCCW71bMoh+Zw70TPBrIrn2G5kn52kZyEuV8+mqojIeLjBB4/
JFShtNc9OBilo0kEJzXLW07gmmZsGWOeJ9rNgyuqVL2n4SSNVUrsUC3F3rKtG4z3zarNz3TmoeZq
dUWmbYor5z2wB40BIpwE7jjDuh0U1JFD5SlGcyUlIRiCGJpomsdVHD7rt6ek13OiA1obmMME6JPJ
WJIgdZub0HiZK1CTa6fCaL9h8sNMyedq3gZEmUZUvOzN6+J5zjPv2Xiz3iLnYRUBF2jbFHSh3xde
s8nhiukTkZcVQxrP1ydg2FKOfgraI+pmnNsa50+YO0pGNx2Y3SpGq+MTa6wIFayE7i0YS3Zv/Mmv
8k4hCdE5cGkNz3oSKY7mXCSZtssOA295GBtTC5kffgaU9i0X+1lrGZtYIZdWC7FA6fBC4Wo+6M6e
UkDWOTfa4FEnLoMc9ZOmOCybAIObnaOy4R3hP2MK/2OYla+w2Vvm/F2XBYSJ/9+OkwNc3NQy131J
tYpEgTnVdgKWjOP0wkJ0GwmjcFyw8+O9xnaTcwYmPxAaVHc+yP5zJXti21lgbLH30wH7Fvi1wzfp
kkF2gApwD9OoFPTH/gjyFTw2ZXLi6r3d+Si6PuRvPeQGaFL/M928uDu0v8j4GAdiif17FBTdo41L
Pa2ui/iMHGqICrrHUMitLn1YfDw+dplos26wXomg1gngC9zyCMDJaKF+cdMBzCOZ21sB9V/+Yogo
Aq8VB1mpFnKs+Vz9GHdVfFijh9/q6bdzWGaLGT9nO5/AufHEkca2ey2a/kGGbyf4lj9oe1FpSWfM
zlcdZidTvkG+Sfy4SpLj0T68ZCiqw4L0TtS3NDEE8T2BXAZ4K5fBoKZqdHVnahLHgCWmeKXcMZCA
e7vBjo9NOTwJiv9yEN3TfRsQ+tV3vgcf5P43vKviaJX15YTvusuLlWc7TQF94/17UiKFsrK3zM2q
jYvGQbCSYV3EEPhTfmJM2HFmjgGMNMGq9co62RFe3lNt3WCfr3Ed5yTLcJv7t0l2KGEfX9k+oo2s
MErYsJKfHHMZwHyFt7B3SOmwMV57aDoxSK1jbaCM94WbL5lR1+PFGITxkvZiscfB+ibMi8dMR28K
vI9Px8PGRUz6AX2ZR0uKWwZjPX1bjTozV/cNAp5HwESCrLyNo3amh716gyuxIBSbBajPV6PCpWTz
lR3yOamBv4loyrpuDqKJLgKV4K/crjQcW7gw8QJuJ3ptNpUDHbS8X73+pLShnIFsz4d3dKAP8Pqi
J46Dbgf7DhYQ3wmwoQqL1XYkLmUHngvWwtYokry1VH3EDKv+ZUfKsCIvPilUWh87T2sm5X/NS3Lg
h1RFt4ZGO9kRxQqd3A0F9I0PFIhDXuytTN99dzGF0d7vQ+UvsA2LgWXGNZcfaLyomDEwS0FcgY1/
ugXdfREDaLAFeLTM+Aqbgm2VkNZSMPORRb0PMB+1beY30UUo9BS+rGdySsW4Q+4j3WOcHf3yQLuI
8rYi3ZsPg56KTEMuH6KPeo8yTgqVgLa1+EF0j6jYS2HRu46kcMhKaxjrCzZ9KkccRCtPvTklNIwU
wiWp2x8+AT6LdnXSqdOgEdg5p2a/RJhoGlCkOUOhRfDlStBPv72Ayqh7o/e+ZF2DUr61HQn4va2R
UDu/TmmeONWQM0MdV2rwZbpjJNme9V2pw0oI6slNQuqnoV/seAMqhc4jbkeUHv2RYA0m8kuVOqBi
OKFMlXDku2gu8UX1trIYJOxPXtr90LXfGZmBbS6Oniv82U3qcpqTW5rOO2sf8ZRLdf5ZiAFFA4qQ
BnTvEQL/dxKYmTm2ewjMNilzEDJMtyWvvQ1q8HUNzwjwiU87UoO4Xz8v3gheu01e//BUEZ5F6w2L
WGqQXL3HzS4gb4MSqY9Hsitrj1ywDsk8DbRHFktLp8vB/3e6YiXyiY5mFjZtPEzCtGb31Eza2KhS
KVlTi3q29kE2VHtXIZgHAvhc/mgLxDw3fLyUpLcxrl7p6QZQiSByWGHr3ww5DJo2bhmjWTggBL3w
4GgK1vfTfLVg2M1BVNlK+kQlGmjLUyCcs5FV2BDnmIXf8tJriBC/8L7XxJG9UD1A2TbZGOLRkTO4
lDwdYtlA/YocNuJwSqEsh4xVli+l3emE1HdPOxgUlkbnB5okfSiSaxGnL62tAZrIp+Fo9P91dgeQ
iiJOeviG2c8aBC5V+juJx+NXTuXpRC4HzAenWyr+HYHLuluSz1XEaQU51De4FUR1sRHyjue74qgK
S5kF7GJ4g5jayeFsnRSGPHqsk7vb6BFFx34aBuU45mz9CcHOw/ifUOh9mnmVLo8/rJNr1WjVajT5
z5RVabEkEws0eyd2RfFzrx7+Cjy1uhvmE5QMI5NdJquD4XN79Ye9TOFnxUYWvj+Btpg6UOkSKTcG
umZSYgE7aWLnIzRYCG1UUEkp7xC69DAoiHfRWaLRdzchorzg/b2qvjG/9BMyhG3jnHcrVTYmPPJ4
h3BIiVTYQreWysYjbaInnGJuZ79ccRQ2VwghvYgIDoOvpWhk/TBvNc/Wbt7OUIbMFaGs0bkJdA99
ZYUbkUcCTnd6JbiENvwwvgh11333Bepx8Bb25vZjQnpx9vBuD79g+aTdAuvWhEAJfnwn+o6bJFtZ
Yzp/ylVVmHJA5O5W589MzwgSndeaBewuoXdwcPMdRBHAoovps1AtGCAHSG2EnWQyz12g0VMDPMIS
LlwVmKpDcsZc9Zlw1S2iDIz3DyBaC/ZmW8MsNSZVKXjTQFfpX5bp2f+8xd1dzbeizEo0Lv3tpX1r
JJNvMDWCu2/udYeQPIX3Gxigc6P8UTWiShrl+0/qY/fmsZsrCPc9EOrJpLIfFu4xeRwbcSAOuvNU
uQeNBqYHl3RLzEEX7MTNmeE6lZNca8+k6mTjcBoRw0GcG3Kc/tr35CrqAp8jUH3DLiLVo7AKHc5n
2bEKP+RwP8M4Y7C0TP8BgrKB1DfZzk+qaeU+gaYgzz7RioHjdqlK2SEJ0Vc55O011kh0uW3iB3sw
LK72bCnaQzqlv/RniIIFPaP4ta6anpB6gs7m+qlBdOD5ewMWLew1+uwegwu2n/wbrQVB4wKPHNc1
Ub+9E73qJj8budaxOU6lWTRjr+ep6mz+lGsG5IcPBQBp+C0PMPyEb3EyhEfNGZG1D65Flk8Df3HF
4zG6dv1JUVQR8cAAZAi920ggq5RsTP1uDNtcD2eLZkJQnUXh5W/r7JhdR0gCFMEbxT0h5cBGXOpv
vZa/oLxZQvG3DO9WNYJLXAp3hklrO8TGkN4QAXxZ4PVtr5WBRaIObyvpQgWOR03kH+q0aQcLIwAn
yoLSreBL+RzV4WNHSz3jfXvSpOsQv0X02/6MQYXP78DWhbsDZlG+9twEezkbCs/EsQ3vvlF2q/Bx
EGeEbBwZEpJ+dlrYGEofQ8Bg5sREDKHwSlJKcwF7fW/ou0/DdSPj89szlCb5lGfb4VNOSiQCAI8X
IVC4TT4yO6Hg7icqetdOanuV1ghTTX074L31z3ll6YoHn0DaHcBtnfRlyhbyolDpktrpKbFMAgcN
M0uX2WN7m4aKG2RZ86Bifkuy33crQ0LzaSp/Vh05uRd7MCSLia8IHJbqKoB8u0KpcMSYZVmsFbFX
+WhZ7iI9wKd3Skxq7gculPVYCUNZnWSE+ijxBzAeDl26v09qfi4hWSO74ecJ4DqO+zxrx7rg1d8v
PtwO3D8JxbgUM173vlX4TXITL7WNjVCA0Yrqg/Q+Dfj7diTmgcQdIA2kyZWOGLFzDsS6QUPaCYed
lCiB6MAEXWtHdDL0KDjRjwRzOlvx1mGM91ehPBy35MI+aj98azLzf9TaEIwmwGge+VzzzdFymmXA
AS8rf2fCA2SlrqfBnpUcP5Fjy4NSE6/hnCXMuCNH89JBBpkyknhj5+9zZglOvVXCzp89TWX7pelV
Vq8w7bd+lt3XByBzr6DuBkTzIPNkWInuMIY+wUJmVT2AYgPQDBleEnmYSfaeGbHqMOO+vJNo0q57
7fi2EQM73fxgt+8HwbMykfyq+bhJ40bSh168BkCfGV/zRxNqoDp5pcXorFXLk7CRt6yARV3l/HY1
84Y3jdsTbe2W/YDVoMtouq/2gLJ6B/GQmrSsCvqJ4rMW0MWP8ghsiW0Fl82JwHLWRlTely3APOK2
8wjVAW7kK6RI+rilgPKnJnSVmNDrUb5McdCA78NX19oPhtRW1P2tiJGJfkfvwdIDInD7wk+pNm2x
gG9LaGg3FfmOFgJulxehSHZpH0s9Rkl03dnA84G+Pb7rFnxSpVFxt95CZMsqI2VpHqlgm+d6002o
schDf3vzWmlhPHXXv0259cHNPVO1fkLUW65uZBUpvhp0dLp1C5C/Wsq6utePJ71aRfxw9h1HUAMY
/537UCiGwdCrMjWw0SMiuATCvJ3pe0lnN5SNJ0zz//vGfQTtjg/VkRmHoFzWeXNXWsSxzXLuY7Sz
BbYVOywqDqWfQVUcxwvFLAXM/2GShT2vRJQPq0WHUVexEbs093BABM31qMou4zx8R6tcO35jXHL0
dBX1wkO+m1BK7AnPewPhDiOYB2eLuGC2KMPYMl13unbmiKyEebBuISIJtJq4Xgbc2dQgkxSWmyCT
khSjBtAdQig/47TZzsn6sikBsnoMs+cXTL1iIXSMAZ7TgGZnOSHgpZ7MCiQmWsZ5L7kXlUuCVS2L
xPiMRQWZGxrfj4WPMdCMjxCadNnDmjaV+1RZhj00XL0uLPlzbHcd62iu5rSYaWpCDk/amMXBeDAE
q66SJQ5IW7Q0y/K30WIHjMVfqSa24gZNA/cjXUdrjQxj2cZeq8Pe4KuHI1f7iZ3uo5mOIFpgWEmd
NqrkL+ntkURPNeI83xbMVqvhcso3FHBFUGqRNZjgvixxyK/tyC5OMvrMHYPP1vqBwVQ/oU+dAysi
KfCeH7Eb/QzrX8uHSmWrTO/9zV0ExW3N1Kj7kuroG4aPNR6PSp1LPojZse841PIklk//KSJtXmTM
QxiDo+Zrj7EY4pMJ6oAkbg21cgHS/ABTxBSrocxus0aGQPTURk0MLiMo/eKDSS39/qepA/foo7iZ
hDOhUD/ZJMw9b7aD9LI89fakoiQSuUSmJztEoRpberVgvKJ2MEktm7KDBKJh5CTKP7SWBGgc0IsW
46yeUMJ1SOKU0/dCC4A6uX81+qqMuNHR14qVVUQIhBmzaDuHZ9DYmXHz9oW1+U5Yl/I/LeZKHqUt
iu7FHmB2jYzGdQmcoAWZ3VkWRPUFVKRwEIT7YtMPw68gkJhDwIM9eqSJ3UsBZtVJYyf6bb3MS829
7gOFc4PSnwk/k9fPPPSkFiU/G3TAU6INa9A9i997vSkgT+DcxmXgZefGw/n8mpYc9kcurG9Uqyae
EhTxhYdgtYOPujHW+iUeaVRQxIvjMVcH1lPd8jcu2HifmmSXLwmz34SIGPAVaczHtfTiDZs3FEbR
7qANm+wJlkmKyKZW/c3Ow+q7GITSR0nxfPaaLIrwPzsyQIveOse4ie5jyxkkU5dysr/Ul68gD4v4
mVTD5frJCEStYx6I1O3J7Q+bHyPdPhiQIY/aJOQApKt4UcW5EEH/VkY8j3mvT5TPvaLBnhirgeEY
+lAhpOuVq7VKsG+An2xYfScdZat6i4zvmk9bIaFNJi+rYTvJ9emwRgze0M2XFbgVNEurBOpAuXbC
JaVnb5a1RFUreLLfVzrwAbg3fiZLr3jXzO5SYMXvorg15t93q6tVa4dsIeoPq1Z3eU+QPZmBz1gi
FBzpAsVlvY8jVcH4ZCIAgVcCDrfEKmGRULojHOmnA2X0sycNQZFBnpOYr16OqWxnuITLysVvPHgh
1OxfrPnSvCnieE8yBQfdtliXW9eSzy1dcE9CNtAAiRNAxRm93jYdUgPK5vOqJqjGwMSJJuWtNZKH
5cnB5wgPh4bSfi712O8n1v4HYJEzfmT+2sddJU7JUrQ7e8px3N/aeYO218E+WTWAWqE1ss5yBMBC
H6EGd2Zo6yhD3LJbQ4GCWxDhqITCQYeNv4lu65fUtZ8Z9QxHbszmy5dHNbjmxOSDLZ5DbwnkNSiD
p/zwoCGGtIBy7jnNljXvRB4eTjNoYKhIvxhEVXHImXP4uFiAUPjD6F20IjNcOFclVNrpJHyiXchq
5eSufct89HhaH+1UtXuIZibBCudQpd2SEMMYxHGwAPIS5RR+LR9TwyPNF4YCfziCUkG4Uk1IK5TR
AR/uWiDMuvUd1Mh1Y/6Lb77+/8YuzREeiEaoV9DagWrwh/B0trMlMyVFvtJwoJS0AujMrZ/d1l6V
qp4ODwLQMTEDW69UKI4j8Tuc0sOZfiSDLFLz0dSUnB++syH+piLCrsqWtIGDGrvvVgYUWVmACA8a
z09tK4KUwdAlw6wFCginCyQ0/UZ9SLhq4cjcXiM3pD95MGTB+tuYIiKZGdUVZv1kijNrwnRQj/uF
VqXbZwNyj+kN/0OK+f7OM8rIWeDkjnmONJQprNcekvPeSpmTrk8Bu63dj2oUrDr6k8aDMqntejEq
50O6USDSA+SE1/axCXP8nfM96gk/PzVnoSfoTzQUUBYe4Au1rfs/sahCo2fwxvdM22k+l62+r/s4
LLHs5IrO5/WZGfJX6jHfu5SnW3nX9Iyv/6MlsrC0IiOrqGiLOA9laFp8UAQ5royiFmN7m3wX1SWZ
SUIegc8aAxpQOjAgquGZmi0CpI5Lhi9slji3UXufccm7d0Er3nnWMAVdQSVDRnMMj87lwigBCw2O
eywxDiDxJOQh04rNj/+U/z49LlIQpl7/Xr6i1/ZnBFkdu3ytnHs3oW9jmOiEYJ+9WXoWW3Bl3Bac
hnDKBgX6z1nQ0YKTL+rpn1THNGFzT4lGSqVuiZv2E7K3yPv8d+NgdNLRr/cq43X78HrN7s57De38
hiUvB/L28k0vlC2J8BpU67HZfc0XbSU7gKMmKFEptBfo7RIJ9T1g9XKy1HFmRwyxy4NO0au2HqsC
El4de59dM7elDC3dYm7T8Wp8RQfK6WHINNamUmjNS4Ha1PYuO1GAZIFDmUWuseafYyBcu/LJ5t6X
zsFfYgK+3dPtDDwZEcBq5sIzO+m0cWV0rjoQTRKnrp3713SyUUj1XLh/jirypQM9ghe/BIw5u0xd
UIy70jbZo89alYAKLTLo7m4rrcKsxIhuGLKSmXnrbqUq5c/Ww/mpX5JyElLqXlyuTKHCic6gKLev
Wi4tMcItTeI6FJp0fMvv8e6Rz/J6Ru7X6t7tAtepHzcZv0JkhkwGVyU8MQ8bVQlh39U2OxJ5S1Wp
44v21Xks40PedOvUtFCSlK8WNgzkTuQ7Ore8zxVGVGJO3POUmmLpgB67u8MMOAam7pfWgLlLga5B
+HTPRjKQNR+8O9J7xWOWEq0PYz+Y6k2pe8TDnAFdgYud01Y7qziFvB03h5WJHnoDu7RDJWekUVlI
kW5uxovRgHSAZEmkzE84wCDqw96jCwyOJEX/qgOQnZ4VJOGrneAuhkToL/LPV5mpMPoZH8tOFstX
KyS5WBUpIxJNV39TJDlYZXKoNxmXWkrAxc5r+ffaKbNR+3Za844e9JZlm9lnMH4YgEpbkCJdnUeU
r53w0wn0i82nOV5+ETnFAeB5NRcl6jALsEQd3Jhgd6sQCuQeVVWhlGFiafbVrfEFHrnSibLVdAGf
/7Lt4RtjtNL2s87g0JQVQGjfsbnbDy/taFP33Q2au+6kM5jIgH/vuku4Ni3Kg2fe1CiuNLYqyDwa
smQOQZcMeDr/pRVIdm/P2/5wHLgfNP4ct4uA7vMMR/OIJubaTNrp+54tLdu9HwC17h3vMTaKRPDq
NvVutp4it7k/7Z5Vi49ome1aQ2jTZhtS1tIGPbZrTj+eqtiHefGMV1wrq2ougOJppDP4TcEC+ieT
9LcfQKjMH/pptd3IMas3PDauCUrRyBhiEJdqC8WeVOfo43OB9fPvqhf5CJxukW2mtYIOjWTI0qH2
hTDq9KL6P0SdnPQSZc/0vw6Nduf7vqPfiKQfZIyXS8vME9DFYsNfBMhUVLnvbDgcqEOzPX7bxqU6
5nJptbgFgegooPoPt+f/lKvBJa096CSIRLd0BQS+lHHnRUlxkPJxTTliqwddFy0SsMK+EPPRnHXZ
EEMCJ6dQM/ziJLWfgFmUDpu4AzbVg81jm+T9GJRjTQ83h1ecZW9sBhpLvcSC7/Lo+gJyK/WgnxMf
u644OoqMobcmeDq35+RijFu3P7RySHDopQze1L6Mpl6EDYnCgNroa4CcwUDewF8/cDONiqOWdHgN
2wFG/DFursH8RGS/2Q/D7V58UWZW9q2RAUsR27qYeVL0Zzx+9sOVxAevZVbVhHu23vfY/JT0QEch
zjaLSPexQMHrxYzetki42my4LXpxN+k+abotCeeCe+DiXG1p+kby9A6kWb6s3QfGIlJQNOlE4D5F
ZMl18Nn2c60xzSfqAuHGYC3ComZTtj6/mVD4b72ZW3niBUqmVOevNmMBkH5sfOsdQDuwDgANPiqb
fT6FzEWk5bRR7wf1enq+PRm2S4skfaY1yR/S7w0MPU5f+2gmox4BKR33hzXQq5VwrojdeTOJOOg5
ITXxzwqjV56a0sOQCfCOS1PgmrTU0Gq5FHouGGac8q7Vf+38tmEnJwNLLAKsm60Soi9GzvA5l8Q3
+XH7azNTCXPuSICMkuILvpx7HYrf4hTMtZ2l3BmmAhBesdr3BEIvzPK/ylz4Y4j9kUWUf+o51qIn
ZYKKLvvYuJWqAJkttDcPPJMLVM8udCjD1w6nUpuxw6VQcIsr13x+FhDgHkEkNJKigqokE6fD3GjG
B3sYUSMiVIOO7xcARSZqFiOHxUOPMsQ6UJFoHU1L1nq6KsFNn/z0O22uRg9HL2iZQT1RKacJfMXv
MuBMXxpzA7NIJ1fdWnrc1a/o4Z8S0O3yMM3r7vQqUTX+Bv9mAP3MHfv11443fOx9mxiXwFVkI/g8
/9Faw0NBGTboNZiLM5qMT3tlfttTR/v+l6kQ1yh6vBOxlv8DMJuuy3lvuKo2h6hl7teJMo8HxWEs
nRW/trbt7QuRTRTL/Fvq1xzw1dYqD8hPzPZmYpLGp6USuYdziseFVEmzZCZkpCrrp8BSm62pnGuK
cwIqyrFCqxE0tdUVU9TyUb+rOg1LItHNOHt5k1roUzdYNVHGkR6LttrKEokBYhwOczYGpiGcI65u
mhr6PUDRaANF99FiZS0w03AHlSjZxkRopdVe9xCk1xdCRc3UESmxwlSejn6fulLRqv10OWAFuSTv
8hF9c0LUPhxJgwGy0P7MWvd+IOJZMfQW3EdcXRa6uvICcgwzYXg5t9hNzb2tqgV+YGnTZ2x0xcY2
s5FQxQeu13VFft/bs7uOxYFraM6wKaywIsxzYmjnC7sDSe7hrY6Fg5K4XT05lR/0zyZdava+mmJk
P407DTFeuMW15iVK9uUmwfzNDjNlfn+NaZArbLFT/9re+kHxtK8VeXDabN4iIjH+867T7/i/uEox
rOi3hQb6hh1MAJRTRr6ANEb01McjfIp3cvk/Ou/2iuMfLLMEwtncObWKtAtuyiOosCh5Tw3cmg56
qkjhLoLCYhOhCQnoiJTpuOY2ipfmIm2GuRxOtYfUcLWmxAx8CUKlYsOzDral3wGl23OimMnXrNOp
UY90Ol+nycqhD87Z0fF5nY+YoZkOAvVmGX3y2/KaEyxLpcDMH6cJo/gZWkmhINAzX4wQx4v2rZEc
7OL4k4xviSNSWa7leVtJYry/6ZmSrNrnpZguCJNzS05S7qJDGLhiyqvDSi1N8ydlH8TVCIq7MPgZ
qd+InjjLQ6V30+cRHufl7rDUty23UjLJ1JW27y9VIajJL1656l2uqdgzw24XID+zSKj00DjQXE+l
W86NsJRgNTxHVJrwzOpMFcMUbCtLH1K3QxZCDUPJMLBoqXvkdwYQfQ/uMqKq8RG6DFfQ3T8kfTC1
C7dFi2/VSqVX/ZlhOGcFOSLpCnyQzp8oTZ6av/WQdsyfNFpldhcHNVcJLWMP3kTsvSU+ZhlbkvqB
YuWvKx+Kaq3jzYaq9Pp9AuKnCUL6wP1Co/fW0BUBev/zKfwA6DwdXQ/kSZrx4KZdYwUgmIGRLGoO
1LbaAglGykhnm5c8410Cx9HaIMlnVZy6R8TrfIidib6IxxUr7lMzd033sl20Bb4/45CKv3dBo2vP
we47v0DVxXbhOnzaNO66UsJuipYyHAPW5Ry3POZ8avLk9Kt6mz1KxB15wA17lemQhL3jStyqlKVH
i//EP6f72Jax7lfx1idhby+9aQrJLZwk9Qv6W2FanlSb4UrBDgkvhCjJe+NXu/rYCL3pdMBZ1xKW
bgt1W/Wk6/eZ4yPO37G194Ufz3gu9hjnF53fWojdgzcGNd6MN+H959e0ddL30THBLTUUSSVq2RQ2
c3yf0c8FmRcgGciESiqksv5tOMzZSBtWA4Ep+4iTb2kc7WqSX1H8QR6KoQNlCu22ilp9bCCwuclI
UvaTZvh0aCZ7D4ThhV4KBzYtKTzzvbvqv8MxV8cZkrNB+G0Q2NcPV/IHVTX5fcjNrg9vNJoolNYp
0nnTfOB5RubQE7m87uRS9/Ji/fROpAa2x36Fk9Ov26ppogsEud8Xs+wdm0tO4wnAamAU2t/+8Rei
oIWfLZW6JrYzDfV38tEeNMfFkVsFrSZec2Ed5OMnQBi0zbdPWDL5QrKOSz9pD1sViNSOuAEp59+j
/nqSgom+EfYwu2YlsKfqHFiYxsnvJasYiwV06zhQ3iwALaYeLJfziGBuxg0xJqjcjZIU1iG39Fh0
Qo1qeB6IHw6lWrhf6olV5ug3LvNhOtKGDrJiISxfgJDEBCa0GZLOCDJt7xB0Et11s+OxAQLMxlsz
B4T6YDsktlEqZViYilsUi6KL3/7M/wbBoy5GOJJbb65ytixUkk5K88Qc6P27spYpvjyCrSW08czC
ZeXex6KkGKB7uuMDOtkeY3VSrPO7HR2CH8RZMxxHEVbDmyBNjoHLvTusvKG46Qk5EOz76jabsr67
m78zH56aT+cauyGzzt/bamXayO3UhwrePINv3lUN70sIvj1e+rBDvwjPpiz5bMfo+ZtlVMCWV8au
z4Vj3uGXsMFDzDrmeB/+a8HPO4vjYptv7mQN1X5ksobaSGKKjNb9Zmifv8Ku16MI3oQpYUzbXIvW
KNqsJitL81FMVqcdfPKeS5K11Pk9ABEknQ7geOGKVKr8Fti7+ZAEooEiOtfDFhrdGF2Z8qL7GwIz
GxzVHJr1NB1VVZeCRu3fCB/YH1wQntB5dqmdXiwK1dreohzU6OnMjycrt4FhH3npHgYj66Kl7gUz
wNRNq5WeEbQXrsydtwLaD3nnnIi41kFSIUXWdnj/8C4BXzLHypsOKmwsTuGPIeFYSIIyHytMBGDL
JG9/rFvvEK2L7tcY05HAvGZ/guy9SO3/Dt8KLDMneEvSZ/bUUGXUN4RhWjBBxOvhFMW8rcmCkOzF
cjjQNs+Yt+wRsYuIv7sorImPnXbiDEpa8Mdnhm0h6udnR0sLX1kiRFGrrdjs+2FSIgfa+8H6tP2r
fDEt0bayTjn/aFXgWxY1dgVEqP7SDAAs69exnm3InQrUVolCgnGeF4b3I9kzN3ljCazBK+Ov3NVG
zZRzpnP8uKyhexzEYSNMnDynvM9RoJfQ62CaNbePESxir2FCtqjVkcsJFpRSCmljoUGB/gZRE9Qq
cB3M9D7VBYBe9jEIMK0SJMJx1bbLT3WtzQCjWVS7lTOoUWgQ4zeHo7jX1zQCcjh/Wv7cAZ+Sseth
8bzlMFZwC+glFk2SmlQXSxMp5A6huRUwaFxlar9fafd/mCRdPgEzyUPoA5wrvfa6mWBtTX/hbabH
q41a5eZxUuZJX7WfhDNtl9JRoQkGlcnaMpDkSs6oRhdFshYolFLeHTaIkg1cDypFmF0Xtso+p7SO
ZaDga4w2xXmBuoVlnGWLe94lV927n+s+XUZ/F41IsfsbFjPvrGardS6luV+/jEnR3W8skDFVLE27
7lryniHTCw5Vj+hJoST2+6AkkRAATbkXSo6vSxf660yomRvvso7IK6Rzu6kIe0KiDyQXJv0sgRle
iF3MzrbXJmMjBDRPVn0SONzh7ezGruWcISivpIN7cLxDK5AuRct8hKtwENBV1B1MuWmeOYwTR9k+
07gGQeXY/X8qBovXVSD7GkULw2z03j9n9Ns6dsGv2QZa6/BiqtsnuySCxD1Hda+Mp70121d5mHis
/BPECAH8sq8rKWt+NUaxxuAhnZLzviiALQiSJZhzUFMA3Hk5qUAgGe4Y4MXkHpHobw1SzERKyqjH
mWAZ/mDI8B4kZgjdiO59Gc5zvNZ3GAEsnycrJBC41MTh7SZawlsUTr3Wl8pbvIYnkuJNElDdOpnZ
MKPrfTfR3KTVszy4E0fdzeo+wLz1/XTjYFDq1N9AgnpsgXUXZFOzTTTTn+BzApj+OVaGftaloIOc
SDzwjIiwGNi7hQmrUJygkX77G1NKuwbIgR7x6WNDhEXejv+9Wn6fapqycWYa7bcbZnud307uNoul
L5dSdhPWvf+cWeFULIzRKTP4NYRY70WOZ5moiPd2K0i5hTREA1U/vNncYuX3yPJt9GjIQGmWNEyV
UxLfLj8TljT+E6ODRVtO9X19KLzQ6bM/2FJeTmJKSrsgAuvF1ZiH/nb5m0lg8d529zURzQISI7pF
tFR3S2OMKWl5jfTg44UP35VDAbu7eQ2J8XfZMQ27Q04nPNlhy764cK1u0vKAnGhLRdk88urRRokc
bTjq6AgFGf85B3Dyv67g0Bzi2tVmPA86OVF6zglVZWunrKZrzq/ZsJS/H6CxamOmM710iyJmMawq
v45toMpfm9Qh4VYdgjnLTJnMYHfYm69MIVTH8oosODF9Pi1N3BiPJoltTAMXeXLSOT4QglKfUNDI
lkFWAtp4JFvr5faxk9UqegyS/Fh7EGtkyMZrEsvApk09ZISBm+CjCnFlgWl2XEas20UzeBfURb3R
H5bTDRRtDr5lVwEUny5Y1+brwgw2SCXi3yegOtO0O+KLNMqceyB2BJcYuZSHrLm048FQ+Yev/scs
giR7xBow2TAvznNb0d/WoJDoN8wytob2Rxo/y5JP160dmmBPyYlKj7IRXf+D3xGVg5HojhxGqYpT
Voe/0431ImnEUTdYFCJduyorNPrNOtOB5ibx6lb+nbDYoetUnjtZDwvzPWvqmtCG2B5jv1dbFUlp
Mi7sx82gtfH/6xgr9dtGIdWkO701tGMR0QMsr9EojxdoZHvabdkZ85IR3TohCf2FhBJdc4lSRpEk
ClFfFme23v505aAkiaXB+qrgkAghZ5FwGg6HOhT4IdSRKq5zCjjQHTtXDb008oxtdrcd9+8T+6h5
uxPp7/6loWtEcwpn8GnrltqH5oU97pM9nXiJaV9KxwPlrYnEDk3bLK/RQsGWUEuPcb+aOIsNc1DW
lwGUQyQyrd8X17IbJG/bxW3hpMi96E4HZH9q4xYCvCi/eN+c1VxYQCXrs4jMhjlA+ix3ZX8Dq1g7
ZpZ9BpObu6zOHj0IPRv7NtYGXe+wnES1cldKsrCbFexl5C18lTHTITHexxCaTPkWo2pQDQxroQjn
4wmzCgn9fR1LrXwLX5uCFrBIN6W9289QdVX79Piz6tRk6WsLlrwKJF0zxw0RjcobHKcRgIiivEsz
dYL9z9klyfZ+JIAX0f/WTm3uizQZDnKxfyEvfqhSUsZ4lm3wsliH7ZohXI15LzCk4TidF6h6UD2E
8IYyi6P+EhSvlXm8zgujtOtAxYM5NtYg7dPMLiZrs+T4SxsAcNvu72Vs/YK8K+bbzJu2Fa0OYYzh
uMD2WpxJV/47XEKlGw9M1XdVvHmMXHsEBKLIf5LALHxVDYOeE2n5Y+dROGlA+gNyl3gxA2OP019t
oh2JEOr+SdhpAndQlCT7KutnBwBdpUn9Qahvr8dQHxtsQBCFdM1WAv1bfcKNO7f4Otizhnqt5DRV
Ey+qFnDjzBmesLpZkuou6tyJ2IwESPPdZEuUV07E2eFmSz2sDJ4GbDblE5YjYM2wjWOvwkoHcG38
BVwaxZ2AOvPBY4zi6yd9WXgz8ztjVkm5cWOHW6v9TEkgFDjv7HdVgVAzcyvSvDSxneHg69OxLEtV
tT5Wtel6DuCenpgGf7bwRHpoyyJx7IOho3qgF+J2nv8J+Km4jc2z3Uae4CrTep9wO62UGN9XumhB
gCrhbrA5I3RMO0mCcfVARb01ppOjpC2mFx8/qQIunkQne/jY9ijWTgjBRrBmksotWj/JvsYB/yiB
AoETW0LhayroDLfOqc1rhO0FCKXVQpcd+B8tJoYHo/8KKChP3WdK1OO9I5L2mC25s2QG8kArj50W
1H1a8CTgwx+QWH2H2GsQwgf1yoYeq3pdhl4pKgu1FETFoCWuAMktAd2KrUOIpLG97nodcIzT5mh8
T3wAzAEkBEMFt56Nfggbvsnhvblwg10sEdM63u0VnEanxlPwlnU7F6XeAKe0L5oGjeMzN5UDwbrd
bmhTE5GVDb25760gVUEFS8RBTD8uiFx7HkhVVyA9EorB35rjO/0Mvz6iVLGWtzwN3C6CP5RmdaJT
7dSShAWxn2bqh0tvuXZN4ac5FAdscQ9cCnmNFyWd7MMRGzsa92uJEIMXKi31rDS2eau8ihiNa8bY
+VMp9aeSPmfZacr4r0TSosm0DHTh5vW+Rt5/bX76Dezn9YzfseqaXEudDHkBTVMXZNBdxK+7DNAC
pbINV4SHkOf6Nm/FiCL8q/EIy/7wXy8JfL05+62+MuPVB0dKvQtbITe47LQmSnKXJyKP4bVVtcSc
UPv4eb0/WzHOaAFn00XyGguNIkV0KYvJ5V/PWChtZNoFXzSKcBcVG6PBP1pOGgFes+1D1UPSrm/6
8cxO6LIf8ZhilcjCkMZvV6bMvOmEVaPplzy2INVrq8XdcSrs6HsmADQTRi6JHdJKxZsU1Z79eiUK
v/gACexvvQjX9fuGPgBgGwE8/sGNUkkRaaTe7tVgjMXw2SIeEjK8OAfOvtXfWglPg9hcCETfiCZI
jEnYygIpNtdls0mTR+TwobhCr/6nbhO3HOU5+MZLnG9f9Ut1ZS6kTm1hC4FeMDDeYIbi8AZcH8Ad
WuhzvIBNo28KCvnT8b1cG7W0wfI1SsxCBgZVwgGTXx2lSCAf46KPlurZN2tFOJJWwlRBC7gyyeLd
IQXUa8j7HkfBFzByKnRhpoAc9slaOY20ym2kc63oKdYj/yktysaxv7L4m8cbqh+gzv/kP+K8WW4O
af6Kw/IC0XO1XF5kOh9R0AEYLLcKRmtRiHHV2HXf4SfO9b083dSXPGOSe2dYP9pOpObTytm86918
hCCdrANUG9mO0u2BfCQMMLPoCZR6FtaDResAs958VSYitBEi97tppI36+iSFQZ5x8w1dgaDVtGn/
fMyai4VwFL80SpTFswVPM1eFOVP7qJHSZabVpt0x/DG98ZsRw2c0I64b5FV8dxnbCnHM0ogQcY41
yO/b+e20Xwqc6IZN6G6yiltbwyiGgqVAk5M0kkwYVJXT084I3roJw4uk0rQ7cgEYeenVHgd8f4Mp
8p2JijEWNrKpjEo3HXijyMEkUQo36tgYekBIpn7/fgQJnTw6xKDdViPSRRapkuAyVBygEMrqVYPa
JYfOV8lrLxf+7Y/3BBphLyFomhgr46D/0JEwj2AcIoSe1vTkCfUoaeR8PY+IV0+k6oXsohjmorHl
z66IztvYunDvRs7JyqhXL2F1tCE2x4aX7qhMJgxrwH7D9UOPTOO6zO5xWPV+2KzlgDx1pmN4s1G3
BsY35LNtw139Onp1J9zi/F8JnGVtnccOWax2lXqHQRn4+Xwvg/Lh0PvMk7FkfAD0Juz5WY1yRtDb
r+oGp55RMz9HaMthX3kD4g/kj6kT3NZaKPQktwoMwQXpI+Ox/4SanXo513A08f7xGb0nkCgxUBZ2
qyFdensp1udCCNmFKzK8z1EiOJCgwTGsHNSFs5/ntCMJuYG/4fGwBldludl5b8BxLFcinxT5sxoX
jcN7TkJAQN+YCcPQ0p2Uv9AEl4prVzlvqbkobsqz7Gq/WEv4sD2yXec4WsUqBS2EA1hef1r5uTlz
AqKFX3afAVGtyV8eHa0LdBXwyK97YEpWaiDZYriVYR4+AjHSVFcjO0meyz/dvWk7IjJdo56IVWhV
G4e8UseNXO74Eri8cGpH0dqASoS+xyLVqceMODDBrlsXGUzu2OXxzvjeleGaetxn7sBKLqmH8WEA
LzgIcPI9rNLcoJcUfbfukuNoIodVTud96qR8uJd/4qztB9fOZ+1ZD81bLa//bs/SPMg63blOR5Jj
HiuHnjbBJsPZC5vngZxJH8KjhxhjeWm/uYdhJT7OGiV4V0uRs1aznZFH4Sbb5glEOdoafcZXJSG4
Wc+CqoWgrAINaURDgFn7FgUw70ancKlMu9zS10Y+qJDu9Sqt/5JHquurhgD8lco8dk82KmNeLweT
XTQ+2+zm5Dj+38/1DwfewS3ot9ngF+dfT5nq63JGQvKyHe7Krpqwyc7iECBKNmPnQL9mMdTrZIv3
wA0UT1wJm2SWba4IEYCfd5COokJEDEXYJ23QCV8uqPD4/j7tEZBZaTR7MtjXxT4iqX4tJfFsfyHv
XKqCGgnufayomEwMmjvgQVEbhcux3ahqa7J2XAtifSUL4vOGUt4zdWgW3vSCpBSQN6i0n6HFHElC
xFRiapAaNWMPz9bssrJfJKK1t62ZQJIxF0yz1YbDTFaWXjyyzwGpPnq/FURxczx2UeSvSV0Pad+Z
QGjpjFgy4H0+Kdpc7S0UEkxSxYZLhCge5RtS3aC6o5Ok0kZbW4sukhkOrDCm3YTjFlxVGULs+UcM
ucqCKmoOehBSSLSavwZDzb8bBjOAaleZ3wDX+z46iAa8RscWOT9CD2PKuikyzR/JT1fZAb1184QS
PlMuVxmEX8ooAKEXVRaOdsIduUMkSEp87d2gW6VZIduLIo/dnfEchgORTGOygdMRi7p0zBC0Tofm
aB/XOseCY4iWlPllWrgjpa3UFqRAxtFWGPwctXPBMdNRUtjFZJ2/tAXstuSzRnaasJZcZ3tEQNYV
AraP4dMdpYJvGBq6mMEzvxt20pxemvMtsAoY6me+j/KfHrcEZ/BqEbhstEuYqRCUzMbBwV94Jbzo
cIsBwvQctNtAnHGNS4CHDGUGqKkzOuL+bHd7/PtSRlwSFsGMvLh8aoypTh9HBhTxojo7Bl70159g
aNJYtPO38DjqEuvGNiFEiyDHkLEIfVu8NvpnvLn+rR6TKlHeFCy9bKbCpnUn+lyeG4Eh+uK/KjN2
7tlDEPbNvIpjvrwWGeTlkXlkEwn9xYpfkvy5fXbi8EreMXCRKTT2WrrSoUG5FXkNSxc0yHzGWh4X
0jAVLbvJelO/RoIinXqaghyr3mqRmOEWG6tndXbMyMw+MoJ8LtteHeA79ysKCUXh234hcm1RDzNK
0wbq1JvRg9TtDPiHonMuH63mzy8FBVMOtgF42R1HMhjFBUUOojmwAQqcMRyagVCfyaa1psaOmEb+
yYJ4aGil+bCDJSrwe3yKQdxKLYFHyscT1hbYOQ3hf8AXBkrSLHS8OqyBpmJOhOCTHsMZCej8DQt2
Gx2hlznj/aYE24rm9acN0Ed9VgsPf8B4+eKzpJPffTim+YveLzOhpvKn8UEJCyJFqO/FupyfhEp9
/vQoVWa+RyptYxF6PPcD6sQmn7pQwYATRHHbGRpwO6Cjzglm2eQrHtKElcHb9YUSShAJYcGRvonC
pfLOf1eu8gElfzYMkkds5SQGevOHaBMGq0Rre9t3v9f+QKrRqQ165hiQsrJSLKfVUKGzBS8x0xu4
bv1xriFCszlBMK7GjIH/VEPer5a2SEgBFi8NsR6Bj7fa0T4K7U6X5IHZuoanfEUXxkc37dBu+bmn
mXANuhpYb/zqH2hUKNq1x8LIUtHdjYBJLBw5bn13wfW/OgOLHJfjtvOOj8nJWQJ380Jm8r+ED9Lo
nZTg1Kg88fFCt283CzAqyDYWGnTq8ncVCkgpfJwCcUbXJgGD4P2V8WyHe56Av5MzaaTGV99V0lT0
rW64mYKyBEusqFo6i2lJJ5DK+Hku2uF/DmWinUWy7b3YyZsyeH3V8vR/7jlgxpc1y6E24oVRfgWT
f0WpHfNy6eSop/XsS6ltqjnSDiGedK5UDocmcja7UiRv70Bh/AyAyLg8gsfu/YcmSQeIcNKEEWYP
oeorhY1ITPbsWKxNBuBF7o2PyXda0m5aA3NVOW7FWhhzdXE0n4bizzHlPoi7wdBIjkLeozeFKuE0
U97vQ4hWCJdyF6FF+J2Z7kFHp7mnLazjVISlckd74j0uXNIO3EJup67sMOhqZr1MQlDxCNvlcm1b
9mnOzxRQGR9jpX1/ehx/CiWzOuWfG6AN1byUrZ2t7xgNCHpR+Q8kewwQG1ppo2yPknrKaYZsE3B6
WBRVDekGC0i5juUKLWhuMier7xtvuAmaHDFfFSY9KoJUZ3eQGaw2SiA7uXYP8Q4UHhpYN3DGo9fl
6fMhGnTQuEu+GrRWj74+NFnPI3Y4V/eAd3HaGhXr1rQ2HxaD7StbRVaSWsjUlPlo0sviRh6USy0R
zwwrtB4b4kn3X58HZQ+bLJhCWKDmfbtJ9ZcnNm4wSSdGe2MbdXV0RNG57SsGAeT1JGuFjHjVEOTK
n6Hfo9PEPkRQvmBfomCEFJ9aOPIkG/hkMBrObslDD92e8/UcHYMxv4U2bOHP7k/ZIa3yti19N7ra
wWvv3pr1z17WvoxxhMxTREijnseO1BHbT8wxd2KGB7b+Ab57lZFICjktiH62eZgQRY33KQf1GKWz
pzovF7lvrxFrz+cW3aIhGe9oulST26ONWotscoaDMvA5tVD4jszKvqskmcUuj/DeEPSSUCJALg4W
/gc+40J3xA1VwIzpwujxqGklHMAvgpL22l75JYnHP7wLAMugruq32vue6F97UCBy8R8icCl91YMK
MtcJBDJpWLPC1ndneDOCwfvfG0UfbhsbnEvfslffXLpD5yKtKrfOFELMV6oXhoDgKg95y4JJIGFu
kVuimx9SR/FeRR+iPydKgfcX2ABO5Q6atuxWxibFcYJtrB17s4VJ639owM+FZccCx9e/ZPdnu3Ep
n4mlmrGHwhNigE86RIpmcX1xAxAywaW6tqv8I3zEwKQ7MOjtygAN0r0gIZGposIPPOgTTxn6OyWA
34pM+yHFTIF4cUvTASYYeVFJeYeVNVCGnepFOSPmig/gQx3GhdfS8ufqkYFRCpdra9AImOaVSPzs
0p+hpuPRrKsGPH1UeAPxzp0BjJJGYaGkJWWgOtyWjZ0ybqMGe2WUk9Xi4/c6Tq6mUlDK5luUAMc2
pZPZdBnxwKeAchepNdSEdbK3vEXiW3E6cyr+Bj/9AJTBLcO49hEEInMh1sw2ZuAJIaIfMbvhC+WU
ge2UKLTPnM52dlTy3nRuZPkE2O2Nx1SGJOdhwM3wJarU3GD75FbiA8NMW4PwlXb2va0DFFMilBY3
bkwQuS44fasrri1hLv4FeIBaHC9deLvyQuz0s0n+Ypsl0NljOhYAvd5TDvQ/ElWznXiyJPE+rK0u
ohqrdKYwbw4mJIE9S7UcbJn6LGPFp+TrxKQVaGv2++JQQKnpzWQdp9GBCur0BGKLbULfFRRDRsnz
aU1HV/ZQBuNRA5JbPMHko98AdkBFRxYzSt+1VM5dpjkE4NI3Xkce8bTKzUS/h7Z/wnQhmxM99p9T
72U6Ha6R2yLJcrE2Pg1VczbZb9YPJFXOw02KPMnEguaAk1iaimNzBR5oRJXOZniLOqEsfz5WYTF9
18p5WwitjZ9GtGs2prgYkrd3gFFgt1m3Fy/3jj6+6UxG+GHtwgeYjYDrLgNDE45x0R1yInDytJuq
mG0pMH28ukKcIb8ToX5sYGXiXZQK36fMu1G3AGwjVDQTe6hAOThcVTlZwk0CYkQgiuGJ7v1WURhh
zbd/UcEERhReKEJpBK6qB3fQG8opHmoFhyqr0riapmbtW2sAjT5UwiXHQmRT/SeSI97k9Di55geg
GIuIuACp82h3QBLED/UmCrlZOvgdRCVtzX3LU4d3kYdNQmizauK2MUsnd8E0ujGoEMhn+0gWuBOU
/AYQgeciJgj72+OZdcQDi2kYHRqNFG2ceQ4RkCyU11+ekxT1xlQCZ2Z4j4hZsolOHnOiuYO5TCPW
O7Mb0xJipc90yb+4rGjhho0Ajwpgdak0tHcizxv9OCw/c9h0zKp1ZcjbqMtS/ZNNV79mvm1h5Snu
HaM87xXB4Rt/+uJlEJ08X3jUNudkfHOT8RrwoHy6fwu9S33Nr+PmQoi+JzjjnioZAJJLrtMDurNi
sOnAhh1pW52MDgjVgG5K2jEfzJthInXtT+uFzcrQ3KnD+juLfrHCbkoRkiPALXPWZid5LZgvpTJi
jTkbINeBDCCKHuTTvfzS9B55RykxG3R14o44w2hZ9HGeLvmq2IuJ/uu4c0CJGr/1NrdYXL1fCft1
KV9gcx3eVV6imSX/TfE8UPgSjb8xnKGkk+5Poq+AgHTTLPn+DnN05JPjVHKaJh1kMDa67Gp/ccBy
tvqbWY9Yw/HXHh7WapzVMwRKqMIiAHN9IRcty6VemWLg/WHpKeF7LNDY8MpcExCqICjx9e6bJFRX
od5B6JgCm3rvCmGzt5Ayr1VC6/iDrKBmCZDDxOf6fTgOUix6g38eLfw25PdiGeyiGWRGuRxF8f5H
N2Iux1lkE2Dp+hxvcJoCnbSeW25bqKg2YQ80WbBaD2cdGgrRQH1Gyt8SIGryHUIXisuKZkuJlw1T
qLxxt0GXvoNIY8eTbM9YfR3s0lFpXNjy1WLGJu++o1aylD+DLMM98rd4i7pcM8qaVwY1Me7wvLzA
vgbJAOYDQ8sa4SIdkP5oaGnYH89+jeU8SxF7IvedwRb5j/JmyBg25Nz0DnatR65EUWBsoGYN2Iz9
B08eLLckZvYdKws83ya5nUI0237GJnRkxRIJq8VqX9gM7l/+n9R/8W0Pad5q09HcEUrzMWA9j77i
OJDMSytVFL4N7xvnbJ8VLFQ9bRQQYyJ/ADOcNyWFWRO2CDibAb3nFcL1sGg0urfMpzdt7Zk0zV6R
+mO+Epi3EDVAaSsHL2wU2no0aKafiGDdCe/9FMpEYiXegaVMwpmkDwfK9KK+H8F1TtDRTaXnUzOL
AlXCvBSEc0tFgFH2QXx90A7JILzdGnNGPuKfjxSymHh2/UT7eGVq8cLCNv5xXkWPje6HNmXQF/Ma
mKL07Ki/IQ3td0J2C87JQZcHHyUFMMjh/uM9lAjUjlof6PUm7GSuD4mKI6KkxZEyk4PlT5SSoULB
qdYUUgNQTq5FKvSIDzX6EQJqgYZPPhLbnXU9Hs7pHiJafsMo8jn3q1ZIn9tWWsMDGv0Opz02tcmv
U4ea1aJ6hwcGG8QU63Fwuun+yALYlrzOyfPytmGX+tPLJ+M6mmdYOvIdXbZl+Zw+2XT+D5WKkjd8
uYGb011apYHuS3nSRBb+vzgB2vusu35ac0kBQ7AZ4y07XPZax7vginRqzM8uXJz82/JZX+0Obh5W
0IRMk2FB5cwt3ydfYfjQ/X86OGvwxr27V4VZQRUNkHi/t1IZEknWk/7VfLyMWMtB3k1jlOWVO6m0
iV2QxAXNu24u1jzs/I+cNwTcsDEDgXrfg3Ii+n7vOebcux/J4Ms6Dpr01XUutUxNI8epGglZg/Va
T5pm0gOuUPklA+IsBH4ccsOkZ20G2RXD1lXzc8eUI11moHnQ3oYV26XQijIpBxpaygukUs7BihRT
YhilkgFpwLYFvlohr86qMNeMl/wBoClHCqZHiyIHhla7LUSIFkQWsmn8cDybqSKSlHHsElCiiYpk
MCC3gXkgXV832wTZm61tVQviwEQe33/WfrDi3krF+VXO54pq9b5ARe+qwikz7o7kS9aio8RXvshE
DnG6Zo7VTSYprB03lQSW6bOup17d57uIvuu0s1d/np8GZrU2hnOFtWzv+qfPUpD5AUFp0RwxsAKe
F9MsSwYE1y4CZwIw4JlHZIU0RPo8m2Sz2Bkc15MBAY0FpiV89iqqdRZprs3bFWA266yz0NzF+QKs
WIdMvkX8dbyueZU7LxgIOcXdNGxIK3YGsXD+uoZUzIp/cnQEZD9TYfk0lOlSGoA9U0OsmmtdoDJg
lUa2hC3ci92GzYRX18A4WjizpwWyRqacVyuYWGaBDNAeEhx8HehvzaC9QlsRK/jWytENrx5wQ6XK
4V4oEiKB0SOeJVK0AbJKrGsI1wxYnHZIEGy2WOphPPPjHPs4CmIanVeyIC+38qNWUDStixdLe/NM
kn2bTyL51UxOxD8TJlRD6XnXkoqCbtfhxVG4GOPO3XZlx1iufmisHh/18Yfm6Z6uARXpUW9K3gPB
fa+CYRLVv27vdkTG89nnOf/EuxtKlVU0xhPnypkDAP9hfBi/hCe9RXii3OkhBzGkicMVHfEqnKZ7
JSU6y5CGL/OhBQcEY//YkvHwk9AlWawpINNk+gp0CyibqtrbLKjRlKqOo8/lqp4SS1J5OcnnJ+B7
br+DrGSIS2I6TWAXx50JU4CEpN1hVKouuBZt1KtTg8r2yXs2+hUeGMrRv2zgKxuaVZZCaBLMLDis
HuadgHo8YYgP8jdsy9qrHVzuA3S7ykBR14zXDTD6Q24No/eGdD1NQgv4BReeyPmUaQX4fo7IF8RT
kTQyz0mq7B7v+vhmMP3l2eRqqE6AVCOHptCWLlafWu6j3YRDOMyYMgZnEy4eWXfpnfDb/7uGDeub
ns2equlg+rGEhZHqGfh18cxSRvZFMgYXLX8EdvOnWDoRdfL5iNKPsrLLWMlS2vWSyAIQV1qnXUPX
2/QP5MD0T+/0shzhpiMU6Z8BgH/XUNW/FBjYCBE15r+OBeedLxou1mhwqj0vGTOXAhzG5kN5z6r5
A8jN8zEncJLrS+t7LQT91UrcbUbK13QiHh3Iq0cpvXmatNXkSvg0XRg9T9bmGlSYsdRAM/jLHbRY
ZG9vqB0XTuMZCGTXUPi2RgBBd5h+ZSpE1MqUm+OD2mE5qLtF1gkdTH9Fc/niD7yO3lwA0a1is0EQ
XC1AXPqPwRNtI5XCkyBwP5mB2LSZXAWHAJTp7Wx4mz/LMgf5b3WxxtZZr9BVSfl/IEngi3WrvGI/
U02S8FVFL3n0YLicUI4smQ8vPgbaaGTWucUlumf1pqLxrDzrLqGEXzPqiT95u/aU/bx6xcmH+RS0
FB4WfMPve8sxqTdD2FnnixO/8wBojUqe9TuC8JiZTWq7nPGijAQYzIYNh3ddOpm6LpuXMbsqBnNI
2cjQeAqG/+vev/rUSWsHbjomu2UzMx+Zws07v7pGls7OcDJDRVtyk0vXTdSzAGZoAv0JE+YwKLSH
0Ba2uaawtfktSh2TEAT0PXTiWZLfXxP/GAnch2m0cBuQ1mRNddaRUCdXLtqTZNS/82/npD80acDu
Fn5O0wGocGg30ug2J51othiYqLmtJENhHxlWor+U51x1EBazkZi9Nv7Amhe0mgwFxiF0BFZN++Dv
dyeHcdEWOT3/gy8HHHJxOmkj4xnIbGZil9zFDtTRqE7pzu2ZvB28CyW/6NqNUGzyQfLd5+SMXrvL
X9nFCqmXglpf6pLmd+n95yaWNQTjpem34kXxsp7BBzsFlxOTsrlnho+kHgJ7KaFYSislhcbFTntk
r31sZX8IWL7FKVoBLATAhfm0pu2QRMu6D+sUJuSJ/CSVhClFOLFFhDLo+kZBbKdFlz87NMu3UExV
SXO+qkyJQeIxVSQXZqq7NW0ULEXakWxoVlqBHub+eE6gg62KPP/AhjfWHamrykFEYllvnHlO2Yej
jrhMqyBtjAKWfAqY2xCzXo8acG/dlO3M8QLLAg3Rj683f7RDmW1L4MT/fG6j8mQm/mtQ00ceOGyY
qqXIUOZhLq/jagNqpnaTvRfYcJ1yW8sEQJvNsGySpmwdzk0U3BTyoyoN1wruvZE4BVW9G2JFIxgl
jl/LGtObQynFKT2TPwBCJ2Lsp79janxmEeSwbs0SGaf517xqQP93Dq8VnsPeSXuO4EaIW+o1hq0v
F2ZaSlVyJ4cIPEsjdnCWVS43/mNSrawNxOA9Om9e22MJAuBPgOzjp/ZivcgDXZHkb3VTIPjMr0y9
6FL6XnUH4DL2mZjXfHhd4hwDVJXbgKdPNwm5sGj3EtaytwMeG/3+UEDhWn8xFnZnMGfkVT6/9k14
gHESCAftG8g2xVX7wQdmO4SQbhQgKnODSlP/vrHOeavDCnCxJi2jBy6tlx02u2d86wbxxUsccPPE
BlEM2w4/QGmAB29GbBNBTlB/tYtwbVviM87JPk+pMz1jsQ1/amrSTPaklbP59CnomQVylgqkTq2C
BGMEkQg9llSUhtAvRtR7+8ZT9eys5Gd/CeS6IEOTvvFFOGT7w3R+vfapSILxThUnIiqG9HZeTvqp
EjRVNr20wChDx8igf8swmlyzx75nps+XSIgSa9j/jtLeuPWlYS5Z5tbB6YKqsK+4BKPvJ/Gw4rgo
YdmQ9392ViEHEJMGcIk75A+t4cbQpjmrB5LGi/q4XWQxiPh6oxW+mOB9Js1YqYGdZ0ltkyyGdHLR
tWJCzYuMy9fn668CiILKJq6cgCpqw6C4oW6e4ypOOeNEjpwdt7eQ0c9SW1x7kz3o4FMt4/u9gs/A
1m2tuejwC1QQuNJrIgy6fWEgBl3SjkKGGi4FyQgfE9hJDmtPr4Y+wX739sjh2fYRJuPvSvMHzlOk
w2vScRawMhq250YC9u0ItjmFhEMWiX+J7o+gqKHR7vuUvQ9LtQdcETK0QoLHTbhFqSxzSNp+4crH
GhFnL/6pdyJKz+U3TIaMYIVRH/tQCvFocxXam32E3eVA5duUO0J1vr2iVqBmCZ1VXldz87RqiRed
qhj9btZra5sOvwVJTAdQF5Y5xprYnz9gU3sKyc84Ts7m8o4s/WvBjpKofKsJmvkU4g8bFpRLyTY4
bF/JQTtUaNwAL2QimVvj4ZZrgVjG+f8d+VqgVVpn7cXxTkkO4Gz4UkJoe4PhxOU3aG8FnRGLOc5p
9CRwlf1op2TOQu5P+dw+0beA+NcsF6Qys4tW98nqX+WLWSsLeP1Kz6+/tPtuMN7yFr2sPFICjqd2
fFaM3TAMJxUW1RJGESgRhajc8l5TcjIwjdllrNZDpOdmZJdJ6b983X5OGe+2sMkX1bVmjvzF/yIp
5PPq3np4Ktk+bsQ9itp3OAmzBLpSwzxtNt8/NkUUHsTZvdqdqHge239Y5yF+E4YcP8EvdGtz/l+r
Q7ymBAejatfV1eV/w0WvGMWxNE7c/Ur346u4sbe4y/1D9ov0ZOZl/z8+puaee6jLsrg8rdYNx/3g
G7+ySpcsMU/fYayudM7G7y+ykJkqwcIVf18mclFm8rXajbVM8O0hcrdCVUrA30uwOoW7hD+gfcOc
yYHOJ1enPJZUBv7o1v505stOWxkEPlWH9m33Z0RzgicVXevbAS+RpnnOEvunnFnqjXJgY9HyACFq
ivQW+psJOp9XQHcTVupQbguyud47ezn+v3p6Ppz0kLBQkEpwhGzhaTuhZaMcQvYJyKyGE+T5jXXE
ePeUYYvt57P3YGagKA/z31VNqtq3BBi96cJ0TZjtR2XrAjYTWKAVO1+zP2wBXGMxI26hYZEEJDy7
DthdNeWjv+daA6el4UT0Jv1l5aqOPPL4w9JPxXDWepNnsfLZPsvrmeUc6Ab+Fec1QJvDQB1yc3nI
IXbdsRisncu6DpNm+TWNOjdj4O6ODEN5WJQ5E29yIGrrQurgDxR151CTTlXkhjSWGd1e8+GsMJeE
KmpV16g+280aK8NW8h+Jfm+BtgtJnMAiljk4NbrLPz8Xhz2yyWSAyWTar6sudaMDYqfuH4nHusaY
K0oV/wGlAlLiXk+IGuXekaDu/anyUNdMHQbNHZR1/HtMnkw5d2VKsb4VBsJvCGmPxweAdEogrfvv
Q+Nw6AWpdFi3uqieZhKDifcJWTTR91G1O9gZIh8vx+Bxog0bFzsA/xymBPnZWnp20rQvoTbEm1Js
/jNVRPKZnFqfmuVWObn8AQEoM0LMfoLE2UKepQk5hW6ATIIXgilOOf+MXJN27dTmPVEv/5xrtGIe
x3uG7YqdGKoM9RTrACegDXt3HInGoEIYYd2XKMJ6uaeu+pa8dzrJ/HLiqqtA7xRs2pAzUsed8Sus
SlS8Nao0MpNkdCKo/y4fAgl0xar3tUt0GUVHFR7HFGDVHbS3nS+yF7ZmkIHI+ofB97oOf/N2EJ8n
W1tyHoT9xQ9JhM+fM8HmDuB0A/AuWaV8uePWXXSLvS1yypjgE/lM04IBmj9FnNLSj/5kgk/bvKzF
/M3cFcT0BvCyTI5z+J7Zl9fV9gyJiYUyzz8R4LWFowoTi1pLy6FC0gzpgMTLQ8UhAixLOVW8r5mE
QwVvMxam6AdQDOwprVIOii8GJHg0Ca8zDq1MWxwAjX2uVHjlTUWe61p+1FWP82GanJT1LnDTEgFB
FLPN80CNHQ7r44hY5xc9cXBjr34M7DmU8riRTCV1Nn+wIR/sz5/xQOTGl1ep7EiJtiyRsia1WLxt
w+9u9Y3c5P+qHwLAKr3NhGS2dNADc4nI/wlSYGIZ84vAmCHVEZ0PnSx6nF+6aZh5YxbvVertmmtA
5gzrlqWQCQMus8o2tcs3w3m9FW7sVx26kVv4/8NNQRR8LukTetATp5wlqRi1xhL9Y4EY+Gx/12k5
oXymdDosXfI9+qUN4uxDhBYtXMoLws8TYnq5nKqLEynfV0WVgFaX5Y/KDzHJVh4kISvOQb+eg1ZL
ChvqQStertQ5CAP2clUD77K2dPtOc1zqubK5erSxO+c7b9iFGeBvsC6/HVsy9Be0LmM5Id4qFjq5
AaOYe3SRiyrLXjafu2mns9gfH10hRscYQuUaXJic83EYmleIV4QBX/G3WqNO6Qof38XTCQfp32S7
hb1sYh0IoffHSACFZkkB4cSBphNiwTXQNugHtyN6Vfdge5FW0fnVOl9u2uDikXCFOBbuDup/cS85
Bva18orWZkbnypGIzLMW0fMBb3BrAFcRABFgtkBgvOlRX9rXvv19mAYSgX52aSqUh0Xe9fX/hwP8
cZT2/OBfznY48X6/RQcJxnZ0AxzxKKWlcCsD7DpOyDZLRtJq4fxOyBSc8gKmS6ZCcqxIb59c2EjO
UxknOE2ibS20XN9Qnb4rf/rVy+3471EUz8YmTD3D0eONuHFOaPsI25ZxOCkK1be9GPMoyctYnA/x
7qgUZ3CVdW01iabKErujATGEi8gazcn0Iz7DXtAD1XY9k007ntvGqi26UFBIsnrp1RP5KLk6VhbN
z4HvwdKUAf8do3WlW5dl5L7Tt2w5uMKRYhhKVXS3Q5Dc/3bQBJEztSagszSv3lWF8siJf4WfXCqb
mCgYUVaGt3amCeQIKPcH0LV13zTVFzMBAywrXdV0SpZp4m1+VqARFEVe6SHaLUERTfi7G6z8BcaF
hetR0EQRLcfDyEhz5aVDlwx+K/SKvtKUaLiEaWaTOj2Ae9XL6k5MRss/3Iq0hlLU4hsC2h8WNQq7
Zo9sApXOKTxhQ9nnb3R+/AXxnno7HfIkh0RUFw4PEWG0Nx27hFwoNMHGljZwEz869jR4hZGD1wcG
JmepqvU4IoPSX8TQCpjUiBbfvHVg/wqh0yUmqKG0x2X6lZ/EJbdZ3QVbgObrdxptyk1RW9V9JJad
fL/LqE0ibouqKbQdW34xFJlLSbxQBgJjM7RzHFMldlzHDvts26DKZJfsV6Z4iPFOcBV8hiNTMwSg
Iwr3z46gEdClj8Hibll094+xCs+xjvyLHz8cd0k4dN6ZMHziiAxb9S05vSuYA613X5MOo4OEDFbc
bq8NZQ0VM8UZxvYbjVJLZGjfp72np5w4H0CyInd3a5a10kGNMKL8F3E0J4ITOyITBeQ+k1Jj4GB/
wRphCpbyl0AgiU9CLb08By8Jzgcfg/oD/cwYUIrTqvzWqoHAjGz9b5ASK1Hpc7S6MQPBMWwdyr01
eGYIs/i9zWWWgOGrtoq47zcKGigxkJiQqvdZsmJgTJHiEzZ40G6QEJ7B3HP7TYPPHKXDgzgiG03q
oePF4mzBLX5qSQm7Q3r7dyMXcEIqdRqBCPz7uAYJ5YJhtyqhqLcksl+HZE5RestU2QL6/LonUSmf
DErQovHrPeEy8bbhH4hr5QJbNwHZgc8FS9kPUPhvdA8q5GskaPgCwB2IPk8JeB0S+Qs8MCY51QnS
j/8LSdMrO/1DQ7WjHzpSREU8K/y1xefGo7xF4lgHOV1OkJCyWItLzmBDNAJvyn4hEJIR5IAFHHXC
rfLTIJiHskVs36QkMh9PUGnaV9FpfLhdmwf+5fbw2hOwKDLiubLNh42k9mw2JGvD/tZm1OrXNBqm
5cHBfCM1LCTfVd8dqNf8D1K08vLNIpK8YM7qGwQ3yDQtWYKxGmqqS30utMFvx4fr4M2D8dw7J3zz
n7HqhwzaXEv66K2WVicU2BF7Vtxg/ojGYojweUpJgKekNyl5wW3ewi79mhMVsXPK3AEYZEU2qoDk
c+nNB18RpI+H/WALz1qtUKPivpk29czFobhWUmiYNTdmC1CdeV/mwcOJCpzpZMdQ6QyahWx4OnX1
J2J5jBLt8ihhodEWOFRRubXN+eQPLpod3MVqXUEiqTZxd8dVtkNOBL15+V0cq8NIEQRh9fp0EN/K
XIgNZ4s10wRMy5u8mJW75wXRcYzVrknXYobAcvd1tSr5+GobiR4yYBNQk+221wLPOVwmpOq0u3KE
zBZwRRHrQUUbC1/OJF9Gv6nrSh4p0GH5VTARHsZQ07Af38DIyS14ygwqFBggfnST1Yslz+mirywJ
BjJfvktAkAaqCpoWZTQfUi0oNjSSpmBoA/Hfckv8fQW2U4ZVAQ5MCYGvS9k+p4stOAX/SSOS1+WG
kOvq/1ZwslvJhf3i5BtGrnEOyb+5wmShdvysak8QZow9gL458DY13SAqIfpAsfBVPhcWvc9bHt9C
JicEUxgCbJwz5fbOBC33Pd8Zfili9yFrQc6ino/RZ52kdZaC6xBknZ6pUqpuG509W6phz9vJWORv
naVaubRDmp367EXLN/yQU/ljxnMh0QDZAdoL1VTxRFTg4pYMu2TpaVabVL8dDZ/DhKAX714/tXS4
b4IDhSavJWSg8Y+igEjcu3l10B1LaBn7LnFGS9qW+yru3XljRjh+JprmWk/BLPthwUo+6UcFbuEj
lwl0sjnXTeExZ1f1TUvvNa0o17/RKFaqC88IW5JVBgy9xS99WZY6U3wdLix/gnZa9xlfP0qnXlVm
aU/bRCzkiCjiDJ71BMPG3dra33K35TCIVRYm6xkFs0RRX2r1D48G/xYT1s3AxaLY3hXlz97kLijW
+gbwBD2De0ZRHW4zZQdJtNgaFAAEY8EaruqbPDbvNu5gYoESfWqo0ZpLVBu/UMy9kBVXxVjP+Ch7
GyF/Hnx/ddICOs8ehlQRS1ZwQgXpqAlL48qBXcQLOemAInjzsGJvSVnHECUgCASvSRTDJWyz2te7
SuwaDDaIzKbRI7Z7bk4UQFCe1NVpihSV3H9IYLV33/G2iUcPqBGLrjX64+4saADPNe7D/ftVdwqp
XZbeLirgTrqYnieVf1P4qJbMOkG4W6mXhogf0UqKsQo0mQSnSnnFf7l3F2elysI1bCeV3p2Fn2Fb
FNR1ExW/jz50XIc5Cf0d1jSe1VkOTHG/40tQrsaD6jsep/HHhS8PYjJihaisomSGwoy/dXcyv/PG
uUi2FKw7MHCfg2XHMXjoMnxd65ZdG+jgVQOIn+y2QPb2bnQjOjZuwSSsP0kDsXCRP3n7lJlTLHIo
B2OocIFquFoB1rPCrbLi+UkWg3HDtGrp6NFEE8axnOo0taMwterBfSsujvGveiSjN3J1Ddi6y0Rv
ftbSVRjSC6VncC4rwiyJJqTGCfx/bNgnWSxTHy8oBe6ZhZZSgqMH5v0kIgVAik+vJpUIHkB46Bli
8Z/zOjc8rTNpQTTxpXeXkpeP4FxpL1p6ZOxJcAX4G/hxpBN266VomBuNPYejiv0rM/R8Cn5vqdDK
Zg8P/VZ4t67FaefNeBagP2pjQh2unwkc22lkgIXUrxLYrptPuR808TvCy4eDkC3gA/I1Bfz7Dxsc
1FwLTpbrsXp5niaPGw58nX3wZt3Hil4A34EeV3Clt1RzvsyrLbmiLR/LKHUUjg7Bf1C0GKXFD8vh
Y1CYGd4bwN4cc08zzZSbEmEHKwvxeNENEGyi+vLGNxIVMCZa+HBsfy3Njv5yhVX5Zw2XetCae7aP
77nrJi6N4J6Jnv0Jm4knqLaBrJI+WZe/Ns2D5EzrZCvtph2+a3sO012r2fTdRVU6Ps4UEyVn9Yxs
yjwJSkRtfq95ofwRduPkdsFBWjD0Fxzyunra45Yh0tosVYlUTFuYdQsuoYP+8uNtpy3RVIAoQPP1
wSzUOMkWCMb3/dMNWGGyEkVDTsUeuW3jNzmovgtX8QTXL9st50JkuHzYI8A3y+4il+DCDcT6z9bM
5j/S7ldbf7mXzqLgVHPRPgQdwxtlYO2h1vCmJG6sDiP6iCUgJSuW2ST5dWlKOy/YCtu6eXaiMtnb
udM04alyn5+DA1h1y5o8VTPWZJQmGtRV8kTM86o4ye9ec37lNdW8lqBOQu65nST6Ij3m5Ngoea9n
vwyNnTQiYU2JR14WioTsfx8pWZrhizjE5t5pYL2HGLItn7ue/O8f5wZmrCi7xJ4Nu6uivNg/M3B8
Y2XsMzD6aBZEYAH5oIcnrHhxHpolmO0UX3orTQVbM9W6k0VujoTMOHcSRyFwbHyB4nzYneXk9Vvb
XLQM0Vg/EB0/mgStR/zUmEhKR741i75aw85TI9HgbrpaXeNEgTLN+tS75wLd3+QhtaUDHxQ3gwyx
x3OZcBkcIdJ2gRmh1Y1KVHOGZgy7tDn+nxq1N7NtZXBCInKItZw6PY+RfYrvP8UNIA4t4tioUQ7U
oqp2vce5U0ltOzSk5g2eYdlMJXGzC40botGmlq1Xv+rcoVVGJ6WORk4+p8D7RE49QlkV0hd+2v6i
auXbIYyDlb36DLIhwI+6mHOFGJNne6M1xMKG7A71tcBt7xgm8PNGc53FN/uJxwAlSTB0hIQHhcbh
j657VtZZtjZtLl0wDyts78f6b5fZGKumWZ5zezfYZtVynG2/mWM4bJm3smavbrAq0co7uHFfet4O
j31x200llnvHVRjKFajORaBqbBPF5jwgtyiYnviiQnaGawsSWGgk0LCXOOHGYAo0GV6mwN01m+2l
CzjY6hHHEDYU0cMS1IgCO2M0qiq4y/I1tcu52Ya59T/Q9JRcG3TTRTGwU9bW3GS7aQDLrTHshd8e
DITZSuNuzGJtzs3z1c3RijRfGA3BKKc51163Fead5quwD+s+r3Fu2enl1O05ChRAzK69OESxNvn7
+ff4hVn+sd6CGSwyCSvLoPLdDuzG1Qe5Jm9ggrAwTcJYvBLc4X9S27u7u1zjfD0xfxo/lWYkXEdc
of43fMDLy1JGgLX6zKBnH9hICLOJ41xJFwLg5FLMkPuVOkrFh/LlGIHwkbLElmwY8z9X/RZ7rkkh
HOi62mAYvnbdlYDLb7nmFQpZw2KG4AucDGXHH1ETE/1V6jgHmuq5Q3pDNxLb7qfD04ufebd8GMdS
njodrV7KApm52kyklnJ+Gp2RX7q0OYBBxnCPxjWAWqloqLfiCR49GrVhPpN0UztpwTfCWTONcVIq
x/sSPZDzA9Wyr+81bUKKzh/Aar36W73/uyEiafvHXZNYZHuwmsW7NSqkqbhQ9YxyBxXy/MT+hoH/
YyOxXm/W0Htft1UdA+8j3K3ZLDJwbBWbc/s1yKy0FaNW7e7kle7BSUSg+fIrLCU+pVacBPOZ6F11
Q0m90PiuzkpzC6E//DjIwUN6TbC6Gxx7V4GZ3MsMPnYTMBqBVcsnS5vDt+06PNCH5MBuavwgKRGx
Fzyf2VsYXSnduSybMmDKSc8v2fI8Qc+f24IW47AvZx1r5HhJGPkP3tHbgH7IJzV1fRcLWpXw/JEe
ymCIbfkjkuGh3wr4quLreYgLjLGHT/lbl/lduGXGXZnybKo5iwSecEcM7rZo68T/j5ns1twjMDa+
IUeg1EtSre17I0IOCZjoQ6isT2dVRoI8Evhqj+nENvD56GNX3si6rN1XKxGhfJL0D3kvVZh5JFAt
G+A9HZV7A74Y9RlysDnT65wme9IIxOsamOQtZTAzF8EeA/MvAvDlu9O4o+lua4NI8vvOwKnse7zR
ABzBgeFqLOWOcF/peQdp6uLMGL0pR7NdFh3rgDAGMjfqLRsDOHRH5kpifffbQuKWK5WsoInbyTmb
8tYMajRBRqx79WlGiX9/0Fg2gpDOwMt5uoY/5um/a6cCbbNl8OQq4plJ+U/VvIDtaEK1Lmy84cKP
rThBh04mH9fI4cApyZwm4mAk1bmizeKBl++UfbSGl30Sc0KSgnr5ypY0FFIzJzsjLUZKRom0LN60
etJ6kqKNbyIiSacWqhbq6pGTZ0U5qZ2IzjuUhQKxehH5bXJJ9YSEuSja9cvELYM/SaNWeZxUpGkx
BzYDYorL5zCEeBYOx2DAgM/guzV+YNdG2G8RNgjA1BHLvZFiasXggx/pf6yTx2lNDAOTs+bvm9G3
vimJoapzy6LKV0fcrqMVZh4UKgAv7LUf1Pu22Oi0xV5KaX5WIXX50jJ8iRntoaJJAnewHdEXVZhU
MwkJnYcou+uwIBXAhtSaklb1JQm8IZ8t//uyP1kbTkLZK75ko8BWwz3JC4gAzELLsjQgUwuzC7Zf
clPhoVf/81DPQ6um0OO21A6pI3JKgtizt0ua/Rpt39iI9KrZ0ecFKvLn0R0d1ZSWmEnlyZ9/3xPi
M++ZYy43PEp4N38H5ICl1yU47qksI5E7sJbbUU3lk2h1SzoiOQQo/Whbahxz+NOD3QgEk6nFtDZf
C77KEW3U79AyZtkeaU0ZGDMOTBkmzdV+BQJhgsve67FwC7b4ozXGoy7FiW3IBt6Y4XcqIPSjdPd8
RRtagPcdI+JtjQUzZvyx9u7qEaeq8ojKDfHfAMGlK7vDQT9jwJkGRiEjvUAYXnWgsHEnU5oKD6cn
b4x3TFAzIBfwk2ZVpsPuwzWaNt0SA/+adR7HiinrJ0IYbGG337Oc1NsdKdSt4RO0qJ2d0bCmcgGp
Baq8z5rEbLtQnS9j3aOytaygEiq2Nu0Gmrq5warw6NxicDTGHbWxbl6IBMRa3fHU3ZMLJLB0d6UC
04vroMdKiNdCQYKR6K6WsRtmCb9X4XuzcGluI9O9LUoeWrrZE4Npe0wM2JoR3ywQ8fms2OZVVkAy
OafdQW5Vc2Q1rC34z0mGdijzH+3LgZwknHhLjLeErmfvmSFh1MP2n+QxwzvGuWKWxb+fL45DWD9+
u8Ujn4LRwN/ENrby7xs8YsWWA/Aqco7ap6sJQ3rlf59R/qPn3oiNWOjb+OutLb5Uma7bFbquEhST
JgJKjbB5j+UexlzEu+1wTvkqhvS23yvCf9XGWTaXpRVeS4W93JGg/TKjJyJV1Wgonn6Us7l9bjpg
kTjn94mbfx4x4jBJNA0uoP0wJiclWucK5aEhN5xS6h5vjTHee/yNPSsmSL7jeOjtxdV4ONLybz+J
r6u6ZAd/WgH4w9GvEo6CBwC+6u6bFNjEDntburkH7zJPMs22Y+9pQ0fAHaVL43DsUfGVSI/N0vad
1GGrBFnHnyeQcDER6QJJbbJzwm8h4nHcl9SaSiVzQD62ZynMLpAiJbaAJ2vCCEpzzce2Bu9AKlzI
FTfdXjw3Y52SaEQg8N/Ct1TWpF9VBXszagetjEMjk+vg4LylenDF4VFqOry9sOVlu9BuzT5Las+p
+VfGhkWsL4ZOvBPFyIlfnnc3cLQSkVkVJqq9HOFbJiQ9XYXb6AbgZegIwPWybyTcXY19HehvyGwl
Y1aClhRofm/lDQs7QyOxffdOiVLkwRRKHKuqD8oWC1JiQMT+TOjCbnCWH1W/2XjSaxp8Z52xC9qq
Mz8Ch5Xr28P3WUzS6g3gFvToHJT03QfIJvdAoalSibp505aPgtCH8Qy90bz6yjRdpSTYb8UVS8OY
iNg1XkYztgnrc3/h6B3+JR9OhcAKjN6MU0N6oSxDstXEidDoqfBpA3SDQ8vhoyZ2IoQMQIMfJrEy
9BDeI0lBQ7FDURd1FkdLNbMjQd1hdnOL7C+E1m+TFlXICyAKpIXWh68d5JAgPikRi4mwZVGjjFcq
8IZxrHC/PKC+uONH6kSF6VXIhFq0eQLWmPzhXuSoXGnSWXI4YOZEpyY0enN4GaBOW1aDYKbHlEjb
GouReslK5SNLCGHR2XpzzNdUTS5mycQDoU1VLTirzlq1xTvZaBZbY6DrBHqZnngcxTwfgQmR4tzz
mWictIWzNr5zYI1H07DVvO2K/E6jqaQ0Rzd060A7+HPehPpNKsYgUWCsmWwV4eH2rOt/rlnZOnZu
P3dmpAIoPFC0nR7QX0nG9p/9kDkMPkFoQXBbzANS6fskBVAbwJm9hHx/bZWRKMxfXg2oQdtU2c8l
Wa3XYokNyu8gyL0KYtu8KyK/BfQhdyjzxPtZJ8DsPwJyWkFVCjegs18Sy+n3vvsNube8GOCK3Mul
1URL7wNi1bEK1XWxLNczPGGBOEkHzHzNpUdLAl0/hzSsbjiEtCQpWB+UXghSouatDYqxtsrEq+x4
9RMKaeXBc8UjGLDtehWDcl7by1szvxk5P642v3QWlq0AiL0Qcc1DHelVirQQGSDQgQPwfzsXRrVr
I7y7avozof86JO2s9UtJX77gfpaJJU3CZZZQ7F4GeVXtmx+gq0mbc8qN78cKr20DkEWpO7FOu7Y/
Nc4ehqdMKq87TfYoTARgIi/d6COT6M4NoBxHQ9zVig1D5Lp8vvuUpCNgQ8+7xuhZH4d8/jpYsoqf
M8BhxQTKP1XbJ7Javg35XG94TdK+RFLuoQ7TQhPL6OSOf0RSiLtmligpkwQROQx4kegl/UMKmLKF
P8PQOoFvm6zpkWaPKqRue+DZGbOyJMas0vEq71E5SA1BV3/OxKuKgdIMtXNb91qlPgIFGB+YQB3b
LM4R1ZYkPfrPNR0MV3HOyHJ5cvKLCt/gSDOKzw9cP0RdvwkIILfhWUK8xgJ+066hcskLoXVzOsa2
I9B34y5Byf676+fJyBr+dZqSThvIbW8GmwXrVqlbkNa5kRd0stoI1iTGilwci2XOVtswVaLcmQIU
LJ49bei8zvSGmlb9hRSPWugc7HwDc7Z5WpfZZiiCeIe/rSvqXOLfE0DVpv63nHI1uVfUQUcRcjmt
bYTjSqtQhJCH00f2nPVyM82huKLjccbd7UtxKELPEk9Bt5OlfvOMBB3SVK0HfeGbgHCNYNgm7/5V
2m+XmXxbIjKoj1//dMbSZtubejhmmozTLPk9logOW8qoy/GHIvxLQDzdaqf6CrZVVaMtzXJvhbyQ
ZQVaAkTDRp2xJVP23Lhrd+lUy1NXJ73SEn1wu+4Rb1tQ+YDW0ikymeGOdDhOmSjTWAKri1TCQa04
4v8rVioecWAla6xDQ6wjTnMdKcJB3S9siJ4Pya93HSLVm5MlEXsYLXFXsE6z7ecf9OW29KaMaf5l
RnXxv8B78ZRrSGh7+4FnQuLJYDu4E2cTh3oHwJ15D/Nub8SgEIN0IyaSjizpe1DPQrthV9QEGSFk
rbMiAgBDmYnEDbB5wvEb30njhkiKKQMtgt7CtLmF/O2I+5OIDdC1DM7LkmGFtbXzushlj2VYeu9b
5wq4e5GnK3UpJKMoQUNiZXHuHTsPzVgH+3x8pT2ZOWOG3p2RS1KF51Fn0giyYL9UX9FcRbeKnDHE
rIoUuwbXbineQ6xuxE5a2SZcOVA0d/o6zOpUtbRvUtGONAuzdLKYnKonjoSIEw9GG9P+at1qAnl0
lsun/3YzoYzr/8cPqZaJ4ZGaqu5ptZ9aXP7hpdBfZf4s5NZTQjUDRZgbGsQ+hpA4wqAdIaMSRsyW
ChQsTdMnxKFzdAod0zGZ/eQUUci/zaAu8rbu6kqPjOUaJ+Hc3wxEoTb0nRm9cshVk+ZsGwhgHBxm
gBk4jlD5FfRNwgCct2SKcLxiK6omOoM5FXWCn+/I+glvMBbR0q5TfmbXODkezy1kDaHjWoJGjaMz
8cWektNGxD506OTHg9yfiyARE5O7eOkhGOwM5PdQBo+dy5dTgv72gAVw4htk5+/pqhELRJfJXPFM
KgXL+8MfbtIPtu6PkH7OK8nncfaMah67JqavNYA4DfStCJjWrGeE9pkPFuJuT39EIkIJdhIgMPGe
3Ijisz2/kDKqLC7vMCM9AhJV+DFGCm2zEjmBZjqOh8phultyptKA840jbAPEqhrOYW8Ld0MXF6TM
rVLUpE6eID4Hc2IfLEfRbTPfLvuZJsLw8G8oVmQ+2/Clr1doYSbofVA2u7Ly1QnDxeVcXJc6nLO8
V2+K/d7DsgX/3/Pz97RfB7KqKE8G6NdNHexvcQ2hm6WhkqAOrc9pZ5t0+6RxGNhq3UIb7GZbIelF
OVx4aaVcp7LRI906jFckpsxnf0GAVdubLgdfKzoA8TzPuEC7WW3lAm6YLg9jm7BmzW/QbNPMTE7l
TED/qvC1FN7lgpGdDc110Y8osLcpRct4m8LwPvKqyliB8ZCUV0muCaf4NT7N85psbkos9qbt0nX/
W8T7HYdR+abRRnXatthW2JyrfhPbo/zgFI/3Gqme2C4AoIsnKPKkQ7zsyCzaB9pTfplFVQLIJC94
ndVl0pd5255eYIMrYGHE45QsyI6xgSU2b8g3EGWTQNczI/4jBy47dMmro/OzGn7ZCsUMBMhTb54h
EtuS8CFLJ5h9WcThg0qvIew9VxhbRB3CKE/jXWRhhPi7mIuVllHGfnKm7R459Qy0LMJIHY7g63S3
i3k2hjEeJAdjibsV4XIuwO7WPHY2ByCJTt9Y/3ZeIrlBnX9T2nnHOqexwneJ5b+P5pMn/t9GDaF9
0RbZIF1tcgfP08fiDvXYCIP42LgHqTKwt7KpRr7673uXQ2Ukucasf8V0Ujk6Gv1nUSx41g8fJOh6
Bx5UGRwzPwI24gEGv7fQXRx+vcGqSwQEiEK9/x6mpNIwIu60Aqnpt7A1zTMa5PaKfsa+J1UD2hqX
eiNSQ8LMfqsbyBMnd7rbtVo6tMT1mMw624q42BqtWw/G64b2RTr3KV1rrKx7Z4K2uVjH8ipzBldq
/M+mb+o2QneJXRqrqLCOOZgR8zwYeu9xRXhm6UDiP1DtoKx4ns3qIJIXZB1fI9X/8768w9KCT87S
MA3gWX3xAxHweS2rhYrnMDiU4WgdayVS4fUXQJbP2j+dUO2NvTYndM9W7JCOVQLZb9ytbMG8IPNC
d18VT9/e0zwVS0/B4cVOynv1/xKbty5b+Zv9Iw44vLNGi1spnKcOPzrgkcBX0i3Gl/uHijH8Q7wM
1tCggH+YW8LFRW5W1ZY6flw8JtaB4KZvfq0I/sziBBQdxx2g3CSvXa6DurYwuohSl9NW/KECV9tk
AnP8T5TwWpTqg2NW3tYSpQ2z2Geei/VN4luq6l8fezuVQsJdKY3zIpxKUhmo4b6nk4UH6FODsbmf
KhPozAswELaDkMZ9VcZneghiqMnHGGoYxVIfmgFx9C6s6Cg25QIDeyVdzOqMIjEwEeK2QIiE3Pka
UnB+wT4rhe5c8C7CT9pa0nxevS7kyu1Zmo6YrWT9N3r3SF9JbPxsK/YvQPc5MO8tPck8X6yyMY4a
X/+gs8ITCoaezMblBUssuK1VEw2TCuqRj4EvW2Wd+zX+ZNuKcSiN/dHJSGU7lTDPKxxCI+N0mum4
LKCCYJvait3crNyZMT7YCrsUn4y0B9rtJSn1wkBC4/Epq5i4fCJmaKY0qH79qxiCng6sKstwimkb
WiB0s3LZPwURVQTnHNUVm4EBSvMwR2rEm1B9PX81H8G9Xb4+6G2xX0LxXRLhcHJBEP5vQ1Bok27j
w2Nw6Stk0r6HnLs/Hp3Aj8U7yWNjzCo9hxzQDvKiQ3ZDqXeFp7OkttTMh6dXzQkpJ7jgoFD3Py8A
gPga8/FXgHwDjlg2Poany1HHKpkkyEOG5tWUlwc8c8d082QlJQN1gdmVjWI8uAwqXG+EqmCCy8i4
6HwsQl6staogA7YXXhVOYOw9iN5qpzyh2k376cCRmrWW3Xjd1WbG2ptHDNc/kYoZoHwVexbmupvp
7QTRMbvhzQbEDXUexvOw6KG9/hqamyHu4VxDWj+7f+OadFbpgAB4jkUXp2oMQ57gfgM8tRuYt1Pd
vff1PM+M+3ccTb9a9hdbn/WG9OFedjfPVp3D9IJm3tuCETndOLSRFwxU4wcGi1SmLbteOyFZAJ40
S3FP25T010f9YGYtmM8N04m6tLZFQoa8OoI1wjyPB9RTsfYuQavjWaXj32QRFNrvqoQIOiz5xTnM
h07jviivNYfVib8vqsbPua83XpYjtOMJN/cgR4kmMX3/BYhbuKNApaInZLycf3Ccb6tKeGxvBAlc
vFB7rNKOouXZ5sqhxWgE348LYcBAefbMYl/gBhVVuimXDcnRs6MoP81fylEgX7gs/6xGxmJBgnwd
8aHjgsEP+DgP2h+Oao7YMVb8EOUGX+P75254AfHxZ6r3gUec1BvxSamIKMq0ifyetd+15+N4eoIn
pIIRFcP/S5MkrLN9MjhOkL2objZ6yTLSLhAE1kKAOElHl/3VJ0T4OGRAkfW5VCsxPz7W/nUoPqGr
8kBN/FehOQtWOCYoR4DvEgyJOsiecMgV+DU9rFCfgX1hjO1V6D3Tkjd2jTk2Pev5+aQ4RaT5XY8l
VMeNxt4ZVarXsNC6DA/Wsnf06PcTiOibK8zC7ON0+ADSy3HKeUtnOupBTeGzup2RQziB8yMN+GqP
MVnxfss9GlqEjZ5DyJZ1Q9CpnsCKUGpYS3SpoBEBIK5y0DDZ6acvKVDK6ntsgWKsAcyh4f7V1t0+
z/1OyWhtV2u0LN3B5ciCR4mGcciCnbLWooPRPV3JZ7id+i8xYuply7SKsX5NplqZV3Ttgh5gWgt9
7jnjAVyQPijpRCuSGdVwytE75ZHH6s+NbSSF3cVfxhX4QI0av/vO//YdP2kp6FqzHFzwbxOWg5c+
q+3SgjEshfDJLdVpnmZfYmrhSj0qevMbQVBaQAOwCwPDxxvioT8VGIB7F8wSiUTyA7Tby2r5+P52
v23PqiPpu2kGyEjapcZMY2GwmP56SQXqlvmLaB+8Xoinn/LLRBedZq3HBRg9kkc0wRKq/6aMFWto
mpEfpZYYsowavGE3vcIP1BphHLtI14QeZNfV9GTYAQo8VznNqnOwraZs5FUxdJbaaPRtf6lproyH
tQgphXDLdBMnK4NM3OxL6pgDy3joPmVbOPCcgaGAATFBi1A/HOO3RtQjf/g/jEExNrPt3ajkMMa7
SUFerc1yXaDWjGXwNRpvdrlPZ7dR80jLMpLdPfq5kpIp7ttOFes9NlxKSkKWUuXGkP8VN/wY4BKl
4fvYd/wvxqUCZUD4JLOZ+q+Aeyu0x0lJzF6xDtKPFsDtB1uCR5Ri3c/sN/dsfYwSDS8UZVUjycKU
bhNVynBKD75OaDurbtS3E1wAqELMWtBgVwILLS83ovuQop5PznyRt1AYnQuD0QT+sOB/1F09OlYl
17kZue2n/a4VG4BvhGTpLgedeliHE+sydzLSCaWU0+6GJbN5aS6S6qsmekWXUk4arSgGhXgoPDO3
/XJcWULIDiOL5sWsbJoBJ81T20IPN/c7whOkB/7ad9Kj/X7vJyeuUAgw5C++EBbXQklfxWg2sLCW
zcrOvdsYrb671DPl1LPEN9StvAXj1URnHT46RGFRxfUA9RKi1Neu1pZ/eIrnsuPt1HBEQLVMNIqe
VgN9iUA62oSmh8ZuBA36phXypwUiYHhNzVHlnrYMGwKyZajaauAC408KydcUrlwEbMONtKSkYG3h
Kmecu/Jt8keZFf9jjjffiyHbpsIMTeeHZ5JMHbMQPpw5LVoU12V4W+zBiXJiVmOoh/6kv0S8T6ml
bBNfHh9aUSw26EJRE/F1ZUZXBebUi78G5kCHPnb2dFhUTiE24GQbxEOpNB+Rjt1uY8WhrMorpo7J
uRmt2XMSol2LIZE4+BCmSubhLOuBO5Pii8HJ1GpurGli3+tkQfeM8W1XC+blG6xgwQ6227rmQGuK
VomhhCgOt7VpHKq+vEVXqOkXV5BWuZtfraHOYic2/VWvWOaylTFzFCFrzkOaFldaRIIY/Qb+uFKM
WOg6LM0NB0scXflQidu4dwkJHJ5Gv5uoOEPGfDkkeBLtoPvNa3fB8aen53NW6IHbK9l8t9OO2Rqs
buoyUt2sINFmC/grFSRuE58+0AfxsYhAcgifTBGsgVaEQ+tHvVN0dfrZv3DCiV4xn0VUt5W4A+HT
URJpaPJ/Bre+xynOJjndGqp2nkbPvOsKfi3fQxmpif8XkuQ9Vzx34Ihe0Rd0PfACKcRhWKIX+I7J
no0JoN7E9AI32faYKBZNx2fGx7pSGumqhkShOBdD5RoStwqOlVw36ZKVxaPBtRF1rmZFybGapv9w
mQ3qL5fb2oGTP/mYr+5ndsz7Q+7E1JqXi3qwjnn4mK1u3qxNZKsvDcGG64KP3eXBs9zfsvqh+/Ou
GwMJv6HaibmvO2I1AJRRf0HwnD7wI8JfVNVyBWxqpZcPFEwFNciQWRC+jCmyZ7fbJKLxYhggHVTG
XHYmnfSuhvtgzc49zfybhcRgdqQSRZK7wKlWxhuHuPDAphklDMh3om4+xMT1nOrYpK3dPrf5kSnO
yPUN/2MgioABMq5DMstVW4E6A/ZOiBj7WdCn+ey65Ox5z+J/lQEl/88HyiRov+O76H+6q9YIbx7K
d5o1SLTSt4CNm29/sIygoDTRgT/nUzJ6NYENeZ1z+STt0pxvj3xnUcBSXiwLnk3wd5H2/3yY5Hx0
hlYok/aTRiSIawMXMQZNlUgZWVNDS4VSl9OABPHpdW0ViYWzHl7aUd+q9HbrEW2kI7HSzR/Vb82h
9H70CFQhzB6ApYtP4Py28g9JlXSqvoswx/ttudOhEeUN1n66XEVa6FZVSJF08trJnLGE31jKH2eB
+f9/KyhEJp6rvJeh9HLBpw9MaI46+KhJ0j59dEwuumkgxwng3hx+zFVoY14h7mlWbkyYAipIVM/b
8CdR/vShusmz0voNHA/5DJ0RGam9SYsGtxcdNIO2GIhrXXUFX7oYquVKYMqXXECPrtThYSXVU17P
ceEKU32DTOEBkqEM7aj+yBSq/yuTZtNEq+wBlX9dJxdYpI9vGGCNzIOzrVB5dnbuVMPVZqsvh150
NK+gFYNp0sbBedTdt1igyXiC6zbrbQ0M5N+XCCKHEJvJih92jr4BUo8Vy1cAbj4ZFVUK66X8EocZ
Kxw8ZuxfaXteThqep7NqLXioCHYmAfXmT0LK3BQa08Ac3N7bpQc8Hw22qCX1DntrrUxN9EKyFxzN
JfhzahMG7hKUalIQ/ZmJp8Hqak7RHPVoPiMUmhViAmyT8HSxJM933YctelrSysjwNlZKVrToKPyx
v7py4JNdj6V4OEB7Ok5TpXmKFDrLAmfBlmXeWmaSW2FItmevgo2wHzgTacLNFneaUGzPCJZpRFBN
9NzNfURYP6kv1Q8ZgJdHSBsHgfFY8btapbg/IPJ25W9cz/Mww+FmLuxo9tFGvMpTr2ZwfTu7Yjgq
6ppapN9tB8HmgnOYPIUs4YLiEoYm0dLn4ja/j5vC0iad/Feuy1NJ7KDY5VKVFq4eCIxEWPxUIjMO
FaZNM7QAk6KQ/kKjNtPNCnThhRkMQO/fn9xTHUUr0SgJeHpenfOG0y1n1vqOFzzWR3jT7VNKL7Hc
B1kgGFE2T9gSvB8bye4b1q+c51ZnXF0drqN3p8Ppfqu2XtecZB8MQeKwY79x9Vq33V02/BHdf80D
fx0cS1mcdl+9Yx46ggsIjTYnRkD7dMonnsI79SByEheQh1kdbERO27P3ay0GQg/0YSKajTOH0U1d
DutFJIBh+C5lV/KS5rMlya4gii1UGlJh3nAoJ1gjjD08yjxexmHBOCRvUGzgDmHLAJOn7QfB9+8T
rPRHNolOGr9lp1ltS6HsbmFYt3njXhSQ/W15IAMi6JQ245UtNfJEbbkkDoWLIQxtdXVnL3rnd8UF
o/KzY6T1wHcRPg0L23h5wO291ZHPoZXrhqHxtCsoqdlHG++2WiyTTTjUbGF+40l9g+HuLwZVe74P
1/ivqAcraZ0WF9QVVR4PvQC1rg4TiKs1VW8+50TVqneOwyRbIvY4G/VQpcFLTa4QU/yezx7DrR0d
6C66ilbKq09zebMzo+mfx9kyyzwhkNFsqIMMyS5es1ivnfKZJexp3VPfmKtbKVi2rakqhRESLMfk
c5l5uQtXOmFGhAmh1V++QjJ4vhR8WPrIL3Au4QUxWozNyVgmfNFdeM9vfakzOFV9m6KQ1AIVfl+u
t8XNoOqxCKnOwSbaE8MQFFBR4eqc/IINtWLomvAEaDTOLpuWMycExFESXkCVzxIJs/crGpMig2LF
TdLeRLL/8f1sXIrRzjW4S7WtXn5jzZT4jWC55Lf0IkEE95o2rsLcHRX/JxZb2qCXYC7+BqGmysQ9
+1lKEhcQFjrYcwz1hrw133RzdFspuVJsYA/h6NuoFVCBTDc4c/to+Ff6iMi6AnNbmIMAdN55eBTS
0aEJJch+6jIjPXPCMb/FEpGwys17Oe2T965xg3McQ9IRPwInrjfqHOjwi5GzgfmLtL+dTiNocUSN
5OBEx3745KfGqQiBCcJFybZmh3ieKJrRlA3+8EiaeWedkzBfs4nfAM3EQTISi4vDoA7taKEc6NIC
37xhCO6DEDHpP9t/2kPiKD1vN2fT8L8rTq+fL6nOyhAsBTkauuzxWJNjLsgBxEHAJfsd0J+7Rbiq
pZZc5BKqggvRdmlxnaln0RtWCFWPat/mj3+hojVPpwVsPpwCFlOn4O4HvB63SfN4WWOBTjU23EEB
DRxaY+DpZYFq0MBORMuZn1AN6CzqoYG+kfAXKEp8uiyQAEXwS52ddxCmjbJhgSc3G1iz1X+iht2T
S8SFoOFCYcVyeGp/K2+IXoP1N7n2C78sraKhUADksymTU+N/21+IZeonseKx9uITlZdGVoGBmNjS
DL4pvKWzeqHJ19r+2dgbujUWT/YPQILSNNgcqJOeMZlusfRPhFlYyZO4b39H4PXpCDcCEsJDPyB/
sznosHsLO7cpGCwUtgtua9srIimZEQIvkNhSrUVyqndOfX2JZQQij3FLilSRMKbstofj/rNaP+Xl
xC9ikqbWOyR3CHD/UAH/EtliywBcFNg+CcoI86uXSXNaS72+180O6/Ciyg18Px2y0dwKLtFtH54Q
0zdZqbmH3pyjScOEVddfg0CguelVw2lFh/aSsKjylqY+jQ0I1q1EjRI5lhQOlT+VL9SCng811aKL
Y0dlZ0AcPdOpEBKg1/o8QInRlODSf1CKDPfIjAd/uYpGcsxtFvboBdyJAEoS+nB0vwFS4tWw9tn/
m+uDuvOAv3bSzDfgGOvyT3MCUS2ch0oEfxjyX5Xtnop2RZ1V7XpC5tZedq5Imgy4W5P1uKgABTmq
VwZCelZKuukiEVCe43KSx6hodvnhA1/TSYKy4MAHdHbEadyE0uTUjilGsxVt1+2gx1NC0FZkWEHS
97tp7YfI0eSk+RsVVV7DEzaZog8s+EXMpVyrL7O2zQy89c4zYV2ljF0eUk4caSKxZqUJNUU81/kF
1gOZcvHWkmNaNybTr+zqNETfD5Z9L0H3LBdiUu7H4kRo/3Sqjdh89ZVinlvVvKXy2xsWyV134h76
cvJ4VJYLTFXcv8Ao4Q69tubAooNzjzfKn4b8UjpfmoqZncMxKH3aywT7065Aq/3AVv3m+4rYPW9C
Cdjm/lQ/tQxtmVIBM7hXkydng0gFN7u1dq+2SxJ7zXHCc3OYpcvgjonUzTmrDpmjT7X6WXVjxWlc
PhjWKUHx4O/7gn5D37VENT76F03IRXfnEGw8IxzKDIA8PZ5GrsfvtJ190p06mdBylAv/xBgyraPb
ZsRYouqtcL3Fy0z7jiumhjp0BdKBD0mSdVcKOq6ipdMik4NOancvHuMi+eRjHO7giGZfCLnkqQyM
gevtUAvPRQpveFAxmPFzU3MCJVMCiXfMXRhqsIhB//7FLbbOew66v4jydUahktOQCNKUIrbsPLqU
V+/E41we5dVQpZGlwb4lhEIgKWhOxOnfc1Fnh0qxcoNVr+VhP1SObbDi9xBPI3ODdSH3yX8JRHhc
cDj77d4xmGtWtFpCYPFuc9vZlluZlcqdePno2iFGLJWgOavGM4Cj1LSthALle6jnrgPNiKHsR0A8
a+xkw6vCXHtbzVkz/czhEaBG9eLGxMnfPa2KQZBmweH2/tmxMKjgFQulVswkMsAeZsIWg7/AJ8iP
qpmaxZjHUdeqFzct15rJdRgTYcMXxVAP8CkbDlomkrhjHThZz57URESB/3UPRq+mfeznf7MKgISP
pRIZsRj5wIJ7Gfe0AHjopGllQYkE+mv1b8tfbcxW7CsVcK7+M/gMgRRr465IEhQSEfSEnwZPpYIg
Yern83Lj1zOcGgWoLH5/5aSrSvcqcsne5sMdiTp72ZqtARyeLEyEbibqHj35rDedbduZa+JLm35w
hjsVe2DNMNNNXcNfm+eIoje8FX6HX8FdA2EKTmN2odaGctTSp+1DyOYcfk8hFIXTdfT5tRJBauXZ
eyLdMbDy2x17D6SFL9TKpwPK2wzLAUXlldAsMOmGnIwr+1p1x7U8H01prxdTOnvD8GM22IJp8ElM
Q6sT8V6Fr/TjHybQioWEwFv36AHPT9ZEcVMtuNZUH/ZcG0yJl9lT3rOvtNcP+rB53mKjHUC4euT6
hYpG2cLj96ZWRJYaTMASu3EPsyKBpu2RI3B2mz1yYMkHloWUJbHXYcGW10Gw8Co52uSFRYKjPM4Y
ZEH49+uOB+KUwO5vnr53z9h+M60WWBl7iW3eT4cpwi09sfo/7OxH0hVeUCMrsjdf5eD2O7e+9W9p
P0a03jl7jPldJfWoutjst6KNUwHFFKG3mlzpr+wiTNHAdr8ty8r/UXTOxOko/m+WTBREGOBZ+o9R
Lg4QEaGyXPOfHlOKwwi6JaKihzvDg+BwbOecDBKfpcvd8nmkDgPCxs109y1NMjYvM3E5hVKvQPc8
B8MDTI7mp8hG3jVuoqL6+HQP1+IexX66Fl6BbkjkOjU04JKkXSczs6tdJXUQYxGa7+mL7w6jWxcG
I78GcR1i0E4gGhL6VIM2aj54dAbAwl9dlhIES+CB1EhRd/5lqHhJF/Visftm9hKquNf8hNqDn3TV
nF82DELihSSLsASQIgm73YxoIeS7Gu2DsVeUecp4ANVA9wjQSDicQNMQwG3xgToU6Bu01Hg1uZik
jkUMsIKdDwsGgFwdouWnFkKhNZJZQHgWrAFu0Oou+jiAVuWXfWGnezd7kQ7+IpqGchWBzmIbDgZt
UAtHk1Vz2Wpcp8Dr2OWTinc9+M3PL3P4N5+WSvgJ84VB+lTgID+WL7pXUfPMZM3v8qaWSGNhu5ea
OzW5qpP9lT7j2Y7rwRT0D2q7kutoBKNe3zKj73sj75NeIxmAZ94KDOqK8uKanfIRpEVQRJZ7N7sY
nNzmjcZs+fygAT+Cv74jGHzrggUYRRtNInsbmpI74Mbvglg0nuiIPO7pIRZmwPNQvJOeV79oxC5t
l30qGgj5ZwV0CryfyK+KzeOqDiM71jaAZ3V3l5mUqHtOhG4se4ADImHOIjQvA/y1l/i8CXFlu/2E
4xRHSNzxhMp2uwus/2GMzm2V3sX+CjVo54TXKD5+nvA6DvErCN3y6h6CzLAFYL5KHbbgRm6/ICjD
6bWEY/eM048Ilr4tuOzCi/z2wBGIVf7x8xDX4Mhh4NfJcX/w6aKrT428UflzQOExUSWHzPqsdqkb
scTpvGBDBJXqPJ8sJPJtwn3JjnkvtQ/eRpRkOEkL/1zYd8VJawVkCJZHDNcex2FDS45km1dvNAki
fxWmBM5253Kt/WBIO/WX1fT7cmLEGz9V6LJyHWkaCNoo25mbjmqVALpVI/xF7xKBDSRCKWNKAD5l
vOsux2qdlm6cE11B8Y2qPK/cnsLBM3t/gUndYd7XLseBs+0rX9ZLUGaNWOH00pSFDxBcsqiiKDP1
ehGsKzIiOxwsyUrkRHX/eSUDZpHAXIK8KEenjwCelSME0/b166SDwFW7QdGhdanx4KyfYGgLC1am
jgBI7c7jM0adkV59XR1eBE7xoxZrYKEtCXRfQ5aCR7oAXyC96uRK96rcaXG/n/seV7CNY3utXakg
NFYzyBd9ia0RdMT6iY8O2qdQ4lKIATF7wBg5O+z+MOjdjn0X/YiRQM6c/Aw7Ml8eKJ1VITuIrAeC
EgdmAMD6Cv7vhApzA+3bvC95Xwb2e9NXPtQE7VH8LEh+6QFEzkvmlKJzBXbQ99gSwux9bTM3Tx8Z
LaNsnOpX6CEILa7c0o+u7R2+UIowFUAGDIHpxtQ4tkgtHrSNGbXl4sND2dDbvL+ZBZeDDxbIxHFW
j4aHs3aW0nJPE91HUSJPuVcS3+ofR5NLokK8BtCnAB1+GZmGO339IrljoeOxK9n9G6bUBDnK0sfP
QwcWKffs+c+281Kv26NjIDTuzaKrsCDbZ5ym0btmTeDa956qEPzFDYVNbeovC+UTNtw/oePeYOTK
CGWclyzsTV7VDsd+bnnqntpBp01qRHL5NCNcrwhEIzP/LDKmjkx6BZe5IhoOYACkV2lt/h6eAHku
hdBoCjZT/anTZZb1VnNRkH7wkA/ZFVumX9ig0615Pu/zFva/LKla7hzefIAQrx4pwzOgqjOqMoad
vBC/yjDvNvuadasT9LoMRIk+GlxiqyQ1EmpOpRC7VCjat0d/OOb4HIi+dLtabMA+1DUZ+P2e2wM2
KxOp5KKw+NZrCP5SNH9ocptd21wz68knJnYlbhqSqB1fyr4XZ64wEZUc9VPrs2c4/vPhynNxaKdA
OhMPjclQdxysVvsP1m6Eralj7kyhVCOLXHDbMCuJtbF3Bii7AXpxfIW5fV9ELozK23OAZ086Z7+a
OV0PEc3AYDoPCsLmbRc6l/Xd68cv79WD/+ZYub26OP2FH7oAYPUyEeMRo9VO5kYL9+FmB+GBwtXM
VEBUt76e+U5bvu5AVmrZ+oMcjPQ6RbzGi/adPRbcRVUJd915DdMQ557I4UhzobYLUOICmRPTsJOT
ut/F8wF1HOYIlpeppnPy33+7qSB7w5lSsrkaF6XSEgwaUqfHC3ZFVtoCUwvBKWabf0lqylgbJqEa
GOB2KSQnAWG1KNGSwG+auA8TehcTlulHvXfY71v8XY2RW5dPuNokq5HhjTJtmjalRy5FxmIC6lKd
m0VwWhT7LtFtO+Q3rYNrlfFsl8QgmxvM1GeL+97DP4IA+lkAULK7A1rgj5Nu+ZpC5JjribGvhvQN
suNI7qLliFuqp3L/cvDXGNuDkgjirEwS/Cj6j5u4O4woxYuGYfrprat88R2VmY+wB1J2tJ+LBUtT
jNr29rzPwdjWYiYCYVeSij6+w+Nhrf/h1oy8tjtFG/UdlTGOOKcgm5A4xKMiTLS3Jb04HwY0K6jh
ifKN6oGCTUaTJ8tvwlEPehrrLhXVqYyps7W0J6LlPi1sd/fha1gi/GJtocDN0ylMVAkH9YlmFq63
eK2DASVKJsyz1xos07mitIoWLItriHLI1p3GxNMKoBOJnXp6nGrHwXwWCXQv4/H2cDXToxwKSpah
bZ2Yt033WcdUcTifk0zX1ipWbv45ehcs/De+Dr+qukWHMwiQHAEQHXXat03YpTDbMLy4PjuAU6Zm
kvEEvN2LaZdysWilIviaF/53vbsBuotWPHhk7r2rckz+RGJH1TTM4PSRqmiAVLAMPLLdRz87kpG8
ijZ6Shk6PbmaEDDoleuhq0VIQlbNUNQsfV8yqKSh2UV1iAHeAUyn6oY2yo/O4Qu1W98eoVekHbkq
YSgI0HhwItvDGvp0Svyf3BtdeDTq7igMKCjbfIh26YylrF+nfsPiIXQmhmoaR53IInZxA4C258AS
8Wq4shHXxaXG+UCDzyAPLIEFmHMMzNQ+GvAJV6S9INNTr4ul/6XddyA9nRgLAGSXAVmMoeJSISad
GnTlWHhBuTUuiHnLRGs7sgH6wD4wrAYSqpTKa+pzBOGpPBNN5jKNQCUvG8mPS6lPJexb8VJVPSdv
dCa5wxAJDVxWvtW1OrHf2eZxgg48Jgu5/lEVTkdJMYftaBCQhNKADdXv8PWKezi6QaViRS6k1igb
K9j3+T4f1r8URfcgn8Fc6aSYi/Q8xwRWZM3YDjtdvhTE6sBndeDER0X1PO4GBveJC+6LMolrAVOW
H8Vp+4J73hAi4qzPakHmgZc0LfdX4FlR72rCBpX8XbCHIX3end94sgAT6xJXQuWNFOLKSuWPVJAJ
SOaTelQl5NOzhjTLDf6V+OrDlCxU2IdcZF0Y/vKEQMdl4SUPkZL44iZQC5cGvSlIh/1CyfX/iZ8z
ZM/3JFUWPj/ckjP4fQmjtkHwE0hRLZMVH8MJK+aKyFVtRNHqb6SRn92PLjSoyw37COdSaH0/JWF3
Sln2AemPDkS4f5nQ7Ga5Yh1asV16DQof761yFPdf4ha6iXsC6XtpAxD1gaHvtaeWVc2OPtPDyPYZ
R1mfJaw449Gf6V3cqhy0IZPftDfS7X6DWfCntORbi631Hyx6PRRHmBCWJy4KWtHaKKtm1VR/MHcD
AOY4hPJKjm68LUcGbXOCfhCoSaaDwsnHO9v4wSlwNFnr4BnWRwc7VesScOBMEmlzMhxBHZuHll5y
oYPNflyv1f8RAV0zpxv/XACNRhwMRdnaopOfl83iMgHXyh6AQ4aur4xLgZeWJF9BemEVfzpRABTv
b2cbpmxVAryX+zOYWuSitBlc7kByXIiSWiwcy6kHW0pgEzku390sB9vzTG3hyNkh3/klTjqkYl/K
8ZfQfXRo7sUPNCYnWuD9PE+zZvFwdTK58p+6W8xcisTTUzMwZ05iMKzIqkYN8I14q1okQA2mMo7q
/gnnCvXoU9EBnO1Bsf4VYug3vX/0RzJDXlEqe+ObEZJSizSMs7U6KmQcJ0ioyVvrhdVCfEHvTMdW
q2EazLf6UiLOTgWn1FNgX03RJvCjWLixWSGhRkMZ/WEmIg2iAbmT06IRvWb/OAVPKJuWo3LrmvG9
izreh/ITDxwALjOdUbUE+N+72UR+T5Uuz/OF5G8+YTks99qkQbxDUl6U8S924ew4LukMzbcpfd0Z
r86Ia8lZXKCPlDdCB52qma1Flj5/0n/+SemTJYTjFCVgEegldWgEicr+Syj2gV5owqpUT9O4uFGr
27EjJBY4hdmOxGP0R1N3JmNUdXUQNJoaSe0SzNpN9aE4IkxXlyQaNtm7ZB5sLPS3QSBZUjgvLqMm
pC+Zgpf7XGZfaFxVltBIsOQ9OV3O3BvVAejW2Vxhn2eJmwU6rz9nTY0rwNPmoOPOGgcIHJTb+rHZ
pLynlGjP9crBTkFfgdgFtETjzTg1zpcey/L2pB7dBO29uYUsTyy+VS5DzV31iUkaaIFEdEMxRotb
ugvJ/pQSq4vpE8aZTZNhI7HpNj7r7zmBcMCrQhDvEHmkAsbZG077Hs4v59HaZ451lCinl3XWU6By
gXVc5uSWURMTRX9xRSHItIzx6iWrRBNwzXRwC6BYLBdjphnr7VKBLuMaXEE/taZucP+gqg5mIA34
EkEncmR7W+NNG1fqWtAHjfhZjqFkN62h4c/ahUOeE7RoMHHZF2ySWx1f1KOqgAlO3YrvFe6iMQZs
Wjv58DcSv/QXDm5myb+Z8eFL8EJRtGdFzn1poFeRJXIWfOvyP0XhZnBAUseflvYydr5mhe313Zzi
O7Biivfgn3QREMdj1nYSLc5dLe2ygnptuPi6nmgVxyh5sbeED8wqT69itTrInGXtASOepF31UZky
XprETp+tDMqLgPcQTclxaKpiVjOVcjkxRV7LhBnLJTWUwTwKoM/q9xojCOl+EjLyNyRTGqdHOvNF
o+tEGfnPflQoMqAyAUdNAevCmQXuKAzOFefRTN+rxDy45lurAkVtP/xRU3W3uL3Yx93W4oMAa6Bh
AKwRJJvzh8d0nXPyqHckgdbS2I+NSTZlOOhySGPk+FVoTbCSqkAznBLh1lZoHs9hnNk+CMtAis65
gG1Ja81fadoZhu1PTnMA6tFnzdDCKQXj0q8XL0e/Qqa0dyUi8tGlx00D45sFq0EV/6mFWS+5/ouX
ewZzmr2BaTdpLIGlKUs4EE1wT5UzeeDkAJ5GoEg2KRkByc4HmnEIs+1R/aczBhhSPf3AfzfqXsp8
kAod2bzda3nPSBSXQNJpnN1W8jDuGVg5fFWxUSTn6YgTJP7T4geFSdIr9l0BQJ7OkeG+2EwdVFt6
pl/Do14eVOb01A4VjnhFDets+hZ9P/FksBybSp/W/J8vVI/5v6SfaZZC2lcW0gkrF5OBMoOcKqr+
erS5HQNhx/fhFSv5g9Qd3YJ3/TUV4n2wH9/NoVgs4qsqhScXL7NhiBgEPVOLZGtpxfxa8mA3zA1u
nxAVkB9AiXm9/i52/1pjHJ80zUjbzHyDdFHB1hEZ9dXPUT70KskQdOjPRsaUt2N7AgaXe1HHjgUw
l/OfKQjMAUK6hUwfuv0xtK2isGGm498wKJI9u8eF5EggZQ53CwANKN61RuPPJ0/TEHtos7aMz5dw
bGCeTqiUV5A3C7PsD0TbTVlCS/KzsNwojxoW8+Ew3/1BJUtFM2WtGARmJm/aMbguhsvptPtlLYKi
j4n5P6eTzwD/C8LT5HghRixe16YQZySQdWd7Z/B0RF/8gsWKd3T909TBMkjeuG9W79g0IrCwhL01
E16OzbamJBMGKhpQjgVbbjlfxKUCu7S2G3Q1XO6B3gtzjCjBfeZIpPovgtR6xuwSBjCsyx8vxntQ
O+mntymAC8VroUdjGU0O5iU4S5+O5gqzOUO2wqkyqjglIfg9O6ZZiAZRO59mOjAsr3Be7ngLQ8Q3
vSKQfHLHBTkfA/EPNLSvn38ToxCWBq/p38VrNtAoCGrJqEFawwi4ZwDbJDYe484S452mLHrcWS50
BsjgWQ5F24px5gGgB1BR8nEsZRgTR+7zS++wRsNbQOOu6nN89cvsuDopYfGqE22Y6qLrfuP4J2Hs
rJvmtRvIu2VUW5XVYfPX40W88rizvDX9RT2QYR16XvZ+Qu2m4+LIoKr6GsEUVAlvJORUBJx4rIFY
rmLneE5SueAC2O4QTq3ni34TBPDqFMZSigpAOvd3wEHDK/d+se1AIQqN2Wdk3IRM4ETMlqeo0qIZ
0SSFm4JokDT/46lyNWJ5RDfE3xWdGnlfa64PcVB3f5incKbbRjn/rnTppfKvesTFh5VJYAqn/zfb
DlQH6um2F+tTC0vppLbigEJ07so+RQj1fEXOvqzGXoik0kLZ5a/8aTlFtU/fCWg7l8qjHsnlfVCI
emB8DKvsGmafLYuvXGhtU0Jmn+57et7PjYZbXw0VWWnybK3IwAZPmG4CbcuW0+7yhs8p9IGm4rDP
72YWM/WxdvSqaoaHa2YtZx94RwYQC5Q+HKvRBqm4ryYFNEhD5Qopsr5teDpNEl6ZrpvrE7Xms4sz
YlqY8jRALbMCJ0ih0gEKcRAzsBM0FdZ6gp9eJ6EDIOT4WZyzk7hkaw2qtCYg6WThkmOauVHxo6DQ
9eC5U/EQ3WgQmPOvsQRQsf9pyKxMMr08fVxNCPb77tcUuGTJmwLaX9gI6D7K6Cw/NfLraNMSEz2V
9W2bTU6aqAXtSMhsB59OyWXLKDwuoQOjvF6Apua1Qatpley7mb+4+GqVD6YtHXT5DDL0vO570dNA
yPn1ncSdklpP9pPphtJgPCvYpwiWiw3WtypPUuSYTWEoOfp/yOdSaGM0/pL3nGkt32UtdTdBSnSE
/kMYMbVLPZy4wuLzEuJLr++g8udlwoXiC000JgsGOWN4jn6TNAeFKvGJ0L6pE/EoLBpcRMT6SUyg
YhwrR7XmOZC6r4gKbT3Yin1DaHMntH1MeEOXG60hsIE8DPDh1mcWxgzhoor+OewKQ/xSbrT5oPTz
/HgU9bFrgAJ9IUo//4xkMSxdfUoXlfCOYl5sLKX28PgjtXLavnHSbLOJuD11DBHuvX0m1xhphadi
G8G5CgAPu7cOtNHNEnLoJzqwFH6SMCu+B1YLOYzMpj7zkRUPKX2bWZ3E3tz8X8KmOOVeRA5Rwl1u
ccODzBNhU3c2fZl0CIW50f/S0gMN+LXPG4Bc9T0pB6mYpi4dPjz2RKhE2iyM/kUTszdVFUjS7+To
NWzb3ozcuKVgBeBTZzeXNndmMRzfJW5b6bVZjhGGrAgxS8yjI0AVIMJ9vSA027BoBe5Cakp6hWeu
EPby7+SnPlr+WN9SBkmdPH7J7MUyo8V3UOJyMrwP2lwbg4JsxPzzhFCDfm8Ua8M3cedUMZ8jcq36
FrwIWJHQCJxrUleJ1KqKCHFmfVbzWWf5PJmMSekqPXwKTF0yKuEVOsbpiXVq/NHbxyiDYUzVUIgo
yEk8V4eCMu7H9EoV5GUVPDZW3yhp+xPXAwyeuBJWNfNr2CroHLzMQL3skiSWnee0VJvh2rfOcpoQ
rvVB1BdFPTbiS8YBRLfv5SKQvsYfGX/G7ic+U40wpqLCVv6dLTPzF64Oh+xL/irkixVK1LPl+qfE
Fg/AE2iUf/1wrtxi29nV7KEUzAemmHuUV+qj6aReXQso7PJVVyHtvUhOuXMOJu6kWc/OR952I14V
3vGidz3WwgJvlUwarKv8UzWEmnAnKMg3whNZujb26emDqR4q6ILgAZ50aNgRW4V6iSoaDPe8JtiM
8JgnXuon66peaMxb9oNA5scQXOkf3Xo0/1Pey8Lodoa5p4BiJUDHDdhcERoXnm3wM89TYLm8FHZ1
H0Yr2hsrTqWXQT4uC19ZXxTZ/RSIK0qdzD4LI2gCGDPeyZSaLvTHc4bbwj0OLAbkttkZROsKLG4e
dPMlkOqcx44JyPgF/oT3Gtrz0Nuu3bCmfyAyJfHag/0xyHMS8zxSd/5j8pTYVOqwpXkeZHkt+gaS
wUt5XVyv8dhIytjaUYCRz3RU8oXZHbSvGmrsS+fCgt4e5NzfG6jbLEoooonspwgehkNKi3nlYAUd
E+CKNJozE6jajcrs12wmzjvNsi383igS9Ini9q9IPRdLv/sJO3q6nveyj+MDQFg2579WO2JiG31t
iYqjxg1OcZ41GD3CzO+LG61GP0eAt8SmFBNIE6r2IpOcbtE4JmPYi8zdQzARaISKe5TngcD5Qojd
fawcrISAUfJnO55GjphVQQ/tcRrmob5H//DzQb74NNMVX7wrvXjJnQxEw5Ge49CkAhtbrmeSnJ37
u7xAl+k+KRlxR8QFw4Nvv3ZDEwdL4fo+TuWdoeDCpSUbAUICBnlr/6nzczT45rJwCpTUvnbiD9Vt
WKmqnSAVKBPE/9bs135zInZnJvpbq1Dzne5vByIE3kkR7iftUAHxj7QNPst6/J5ZmHnbpU12JlYj
DRjHSzAgvo0pPs6rUxHBkVPYWpgd6YMokXpkZ7LQFY7l03Lu9FMkfbbXBlwGQC/M0vcqK7oId1xI
+UBkFHmChvBPCW+NUKRKAlIjDlTMQ0ZE5eWgk89jDYXTSpD1jq8KHpciEyfoMd7Xr3O2Ua4KbwdM
Yo3eyynrEA+6r2FOIHl+LJzofl00arhUfqlIAhOsTOqEAp7pKzP8jePCDaSiV/p5wOEo6SheEYT9
NJ/aGt41nvkkOnyXn38qciODoKRaRAsFNk3XtYa83y896YFzAL79iLtKuWN77Zog1FpBByNxrLxi
+auYBhOAb3qIU1BCF1I7TlWmO5OxgACAKI46ZJhRZR7QUzdqPmZCelkuiG4RWTTZqg8iw2YSylll
/zhQIJO8FSjeyutefhpaLbNQm1dBL8pCHxiVcxoDQo8aNbV4ZoT7xJaUTERQhCWBoLygHL3o4Hpi
AadA/rj5Syz0rxKitgI152+mQrw9lypD0NbUqhcw1lz+ibC4MGjwNiyAspHahL2Cb+11PGIn3ZEm
PGGFd3UEtbEJEDXfyEI+gH4pSurnPdmQ4uoL0rtb2juej+y4Brf3IEblNBVgdNgcWaEieUVAFs0D
BrQehFA9JOi8Hs+MwNE5tCX3AdR/ZiRWN9DbWaR2hogJsk5O3AKCiKWDc9s1O5uN12XL02u3Tgq0
7CTXwhXLP3B6pUZiXg+g/h1FPp3pYltHycb1YOMFUM4Cgqd9k8nOsD3NZpO2lwOnkk6Fh4Ed7sCf
fwUxOMWHQBwsXwAH2cdi7h/aLp0TydrQxaFdQfwO+cyJGhm7dGuXbvM6jY/8i1PlIje3Nh82gBFl
28HzkaqXoWa6gVn8HMyICMoK5u/tZ6W56LOwaKwrVFrzORXVN2T7SIsJk3bnN0PiZmUesJeap9yt
1MJX1TCVcjNSee7N4rNeli/kUv8Zll5vrPSmWea3rNLaxzyGYcYEADx6t9CR6bSd/KmAq800iflg
u4gRCytIhNqGc2mNvRyZfunDFdutAEI4LvZmKTEvBoMA88Vwa4HUCJTceyDgKWs+VFyzDFmScf2g
kUZD207rCybasSVBH9VNb8+5PyI9chmczXj/oyQ4LXFVxxPmwmOyF8M7BgVuFbz1UrfAzmdPiMic
Wb7RfkhfZ+rHt+jl/jDP0N2r+Lq0c/1P3PKEukJjQ6Ib6mVIhMwqLhO6mo5C1Rps1KsNofZoCEis
B5FNpB6LPSI8lis4bpy6Xm24o4/dF64zGXfGZYY+bTtZOZq6MQGTNmFRgV3B6uv5PqadeR0ydezo
yosyDH6EuXK7Wt0xa5n+8F5z0uxD2Sjr7nVbLWfngsHztb2DIm5ALHCoiWxkgczjZk54fs4V8bZm
O7kx/JgiaTCUfajqKz8K5keagEJqnMmnKwkLJD9SSvctJ6NkzcBSPW8alzM0E/MBevJRRPnZ4cN5
IjOrti7G5bH2W/lOMJGMg1dAtZnWdSKpx+R7Q5DzbENa6wjT6hZhP7yQQJk0s//08HRxqxPnZckd
Cr/y+SrpEgML/Tfn9tv7nrgjV47iYPShlWKOLfqzdlEyvF8fvdictvYk//pEIBXtx4topiidi1uL
/xXxDB6EB7NThG05C+9K3ReIYWf8KMICGib42cvQv4agCAP2IV8swDgHQtaN7wAhxYmlIr/YWouv
Djoh01oNidVvsnbgc0afoo5+3X4JqtnVZ6EkL8gZAr4s7uw4bFAzHXoNae13al8BoD/4YXWGsbMo
PMJ5dFmf06Iskweip8/L68BESDJOCdGSpKBYXGeh2+hjbXvhrOffjm/36Lfz+Q73K04ZfB3WtWCX
XxedWbv13MSeAxYHKeAAPF00dWj9LNgxP/eqO2J4VJDk5NuWG6syvL5Mws2A5zXwZEy6QQsIRin2
5RLILAJ5AVHcgQO+61sGeptEZKwsOtlpwCWgqhJ7G/NUqq6K1Z5/4XKX9BLuX+TCDcCbkJpJEJ1W
2u7usru5VqaNRfCoinsBsRAgSmp8lyImAcoHpsKWVybqgah+P1XHZxaS1T8MXW2Rb4r0O8QuqT52
8Ws4jlIvGokjEZlT25YDxx0lcW8YmLRMzcfFL+POg62o3GlJrzOv/uB683No0Nn74IyTyruA2din
FSQc25d5yd0Czp9hzwJqpuw9/pvTHG4o/NxieS0+V0j6uyJi2CW1Oxm6tZpIQSFz0xDz4ATKbwos
2vSKz1ySAlw/sD4qyqG+NzBfwDNT8lK94Q545svaMfktC/RWdWhvHDsU5nPKHkedVVMteEY2nxEM
FZwGF2BGeFfAcuZ7Nr2DUZxTGPyry0hOAPVcGTghuHT2/MgCxzmEj5q1qjWqxRshPFrv2DwC6CqF
VKmqbcdkjxyYv9SiWYL0krexdABE7IHSBqj2tENemaZQMlSYYpHKq5M3DtxEP9fYe5LuQfgWNVJW
lZ6Spvk+QAFL6FvcFYDwn/gpzBahfVfg3Z0oH++S1YNG5Ccit8pfJ/8L8XpWDZcJcgvnDMb+CZAK
Rain4CZOW0gVZk9ov20wJp1MAdBvUce5hnHE2OdK4wXIoLAeHw44FhYEfdGNALEjljPd4ae0K2uD
+6E5OnfQnktZllDdvDmSufcE3njlq/URVv6k7aaeDhrJH4kVCajhPkSU8vQw72DkVT6kK89UzAW9
sCcvP2zS4Dq7Gm780wSj1QKBTSSpbFx7r33V1ZOrNzXyWr4v9sM3UjhuS2f1GwA+9H1Bq6BqrE3N
7bQeZB3k2mEcCxNkPXX++ezFiJS/SHgIfpejZdfctKpNNkhiXCYZ8ytyF2T/MiaUBfmZ/Ks6eAo3
hoYmjUpM8j/HuteTyOwo5u30Ugl0Rm1IdlEn59+BqndCW/aCcW/YgWrGA8ZIaPKva6IKtkNQtgBt
jjNjSElUetY5d3d1dqhZo7X5suBD+w4KNpbwCxGQI5VE5Fi1C87y/CUAzfkcTqf7l9Zzeqz8VNqM
pH7A8mZwdc5c2fhEc17lh2jcaxq6HGp0fy1v/KJSyTrlxy76bbXutYnsc2zYIRl6gssqYZmRfIsI
0z3HxmiU/oIHGF5eEw9Hsj22T78Op8MsntwzzzshfmxcggWEu7XNAu1t53YKyepfeuny0w7mg8uW
Id+Q84afpqa6gBE1iCUscwUAK1RjcF6nqIEy8gqnNTs1vkqujlQtshf8DJUmDh8wuwWlPoD9figi
x4rdXXdHzLR7ZDrsNPkK3xzZ/0mq1p2NEA6IgBFpzTUDXBtxuvaITLFiGHWUdyhaBVXV8Nyf9RQQ
29UgKVTt1sln43Ey7JvxH1saZpIPaINUq2qjERM4jjX+Nb4CZWAN5O9IflGFEwjsQbDsQnBnX7Je
4YNKT/5/otOrpY9TYMhF3xJc+tfFCfcwh1g7i8RChkPYVQyhlnhvRPhWmmysxIh/IcANKC9NeOt6
3tDg28M2ymzEnlUM18aFGSfVlfj0hRjl2c4X3oCKM8hgVpvG1kfugeBNNZRA81WRndMtyWxknqkO
UoFtyK98pa7yKR/3f8yT5pwVytpI2lOUahpRqCb1NRhBwZ1HSKgeYBiWNFQMzuVMWT4CFF8m192E
eZiYrKeKfDY5/dlTBBmWuGDQEpRR7euhXHSShGgSOOAarzYPNVwYIpOLcCO0HS5xEg5T4/7jnnU0
5XzDZgGnL2bE0kUsEVmoV95W083DUrGEikY7soxODfZc2jqGqr4dlRwxh/XyM5ktqCbTapAmosfa
geTDv3UON+0fc2MOwMRLCIeZfGcxhiAYyn8xlHXRfAViAZIKM9F8AySvCti6AL7uSsb9Pqcde9Wx
umJYCh27UP9wCjt96iI9kHmd+CM5uqLa+VWUk8Womj6jhUhkh0uqyqIGgd2de5jirnqjhYiD4TU9
ouehKVktjhNP7EFzWk5R7uxP8taTi0n3BrhwujliI9Mki7BGVABzQRMX0SoINU6NaIQ8Q5G3hNaz
6gtL5YaBSn0zP9CLMHf/Px7hEWpTLxL+VrD8IdbSkoFESXZnlSrJeFET019um29C7hXn1AKyy3qK
qCcNF4TMsxw9JjMso2mShuI58w4veinv0V2IZ7xFzNQ/1cuk+ZGY4z75Wc1KxZl7BMYa7/Cdygdd
KApuYm1cGf8Qu4W96icsrL0NCq/q071t88UvO/KdSTnsopKzwzieb5DZt2Bd7oAAYIB9WLyj9k7G
9K1D0qQt5iu72F98TrjQzuLnK7I3NA6F6R3ceCEhghWnMs8El+92SSm2gECQXhCUI5A6XVC7Mp2w
B/ml7zH3HQhFjrQ1E+1J/CsKjaD3hFEOKuwM5WEs8F3RqJBGwZrUJhuOJoHMjN2eUCvoohzziP3K
4h4MbPNhoCn68s/kQx2K0k2p9APrZzFXpZLvsiqv+TaOU2L+f0MBVtgBEqSqNZf4uc8P79bxi3ZB
htIAA/gz3bxBgQ4UP8pT8+mIP66m8Fu4XH8U5IiP/qRLGm0/YX2mxqK6X2P9acYimH6ouzzCdcGK
RwBPkamZrG9qKp/Kmut95TOHiDi2eiFjyCS/4/5ZB4+TxfCae/TjPXGV+IV670wugSeH2GK3/SsJ
1/MV2QLkWVRHs1enep2PaciQnz1X+5qHTjcHZpSf2O64A1Tt0hghjzg+TCvgKV6gmbZJjFpu9di7
WioJnLCv2G+b/E8yDYAQZmuvIo5CcLU0jRBQiWWuEwkiuCTmxVKnDE8/jmFFZx5aS57X+2mn7GdZ
UD0u5FTj8zRu0WAXwpc8tFLcanquvUijD5h2R73tcrrnVJzv7ulkyN2O1TsUTzhV1S+wiPlUJywD
HY8TQQLNzxoFWCpRgKsHYf8V2lLfaCP2wPRg04MMwoeu2SNuCKFvi+sEPP3nq4UlvNy0W9V73pCa
c0b3OkdvFTGBeHic6Z02bANhmvBVS3Tjmwlj5sXF7vG4xHeayhUaDaA5YCrd8Vq5lIDLcYmrzMQ+
ZhPLJNlSb2YHIfVSUmMz7djxmMyrb9RjS0oNmcN3aDjG6k0o9qUcaJccNowDXkAcn+lKnk8+Cnhe
ooe/IZX96tQs7rOKU7oeOnplSKm+HWAs0sWvZxSyFC7qTxmNETfnacB7pBQbR4BQpZOGM1Cw20++
NbAEdkTPAB/jyX4q5Wmn4qBhsYUGDAnzERLGoIqBxpQr9UtWU73+AnLOYwDqWRad92tX0yObs7pp
G6sfEDT4mjTZq8NwJxb+V2+3xT/RjYzDilFDgDnR2rvXhv3PTBUVdZy1Vg53yZChrPpBOeEXkSxr
V89ams+j8BXX1lR/iGEESQbj2Ra6ws3+OPQevV4mV4IaRa+TEHz56dAipZq1hF1lHi9vHNMylxRk
qVzIdCm+7X1dlI5ZHWN0VZsSlPcaKWzoGzDMXGy7DLj3QnGaFbM2zlxWu525MlOe8gfRY3B29b2B
xjfWNZLYtRlTXAZRzWwtYu4M6Mgklggb5q5leIJTl6tVtnskrllGxe/83pmBBoiURenMMljA9OBL
ajHUKY6IM50p/6tsYmdFpVONT5wk9klLmGRPKmy9GCICX1XCOPB1yzSwI2gaZSimwCH7r6QzLJss
DRase4Aq/q/hNmJh0KmHieWYB96ypxcq3xTMaIyB2vQGg56A8AOgwF42jsn+vao+qBxuSSPMV09F
WUS6S7ZSXc8OEFNdxHQ/jAw5fUooeMyBq1vYw/s+dfhvq7MSIgCEkHnP1LfRDbLftX2bGp2ExXfF
pecPtgzqPsCmxAJf5NDjienWsqiSD2D+HdOqQqkZzqh4DtDACKog/KQZEeCpeWPEEQO8RI25/V+q
q0KPU5xN5nnBm1QmPBWt7xQECndCWoe0rcMiuayQ0aykxLqgb3FuhlDwwQmNMHDbUqKhvdjG99Qz
30hpTtNrB/FOXciBH5+I7+5N85mpTmCE5IYB8lSaDHfcK0hDN+4kqbgcoBXusm7h2M4Q3bFR+k0k
D0/W7jdTI9q3S19H6zQ50GBAaZFuym4XbvbugOXyI0pBtV8SjrG4q/3z8bRGTAmSRe+dHThw23V7
Op2T7ie02qU8LIXyB3Mf2B/59qehd6LYs6Vp7CIe9nhG3qoB25O+TeXAIMmgVff7nIfTP/T7yT/M
tDeliCN9S22Ib8uWJyDPJuCTQFLw75y5E+L6MfMLaiyTCJvN8mz777SEAcoltoj8chf+ZwIKvHOD
n6+1jvnsMQi49RrZVeOHQQgG9Xf7ryniisfzZqa22rFzBSAigpGj0Fp56/B9RGMGZNxZJOcu0MAe
bkmnH5ioS7mEJ2UxHQGnfQDcwljp5wcNCz6PByyrxhBU/cCoGy9I3PsdUcu4mGwW00CcL08MVV3c
Rxf7yw31rmI4YOMK7hb2EajreCaA+f67ubxp43v05aJiawCiFQ+GnR+s+D2SQi+GgSYqYl4d5O9U
+19wa3ekUzj+uAiSZMDo+YRvdKSGVMy77XA/zZlDYUfvUS8QBvzAVTj+z3UAc6NxR2Kb8JJwPD3I
qFV7H8jdKvwGOSurWFk05vddSWnzcPHq6EnNVQPdtB9Bs57uvJbsVVC9Yb4DWl67CGyE8q68g7um
fFrXHd4izCZz19INuaE7R2lU1HMeGV0c2f2JWrO1TwKV0r5qoDnaSFgrVUWv6PVXvQF1WO/UHYDE
luCrPEzCCYlp0wCbm91YDPeuuDJ1zRcqwi8hdNjpjqUj6a+a3mn8sVYlLLbEJJ0Zz+tA/QJ5FSWA
VbWCCF31NX1IsRs0iQ3mLeA5FmQnMTg6p8bZodyZ1xJF8hD+jhwL9yzhJVMtTQ/7C1u+OWLbG00U
E7JeBxZdlMVGmO7J+qn88SHIZwABQ89H3RsUsrJWhnCd3CvOyMvMf4VD/IHFbhCNZtJ8J+3kKXQR
XQ70K2SpcBosWYJr9c9v3Z2XFsYOyTIi34TzyQLw6XMOiOsLFq+4CfF727QEwJsPJvLyMyaH/vR2
9EfVFH7zo3j9Qc2UxORIR9SKNUfVfnTwgDZEEKSIIfKn89fvT145rDzuFay9LefzIiQ5sJLFfKlB
sxZFsnMoJgqtI2UUlMWZsIr51iQKpIs2KyO1F2nO15uOD+pR+MCagzGgLla6bpxLdFIErBlrPYRL
06eCYCqtBqomDsgSUvz9QExyfsP6Xol/dNyCxdP5DrRUzoPKKLJrSi3XfIaVU+YRoArZjf4n8p4p
dcaed3ugRcj7GLa0Jin7lXXnC2h/+pnBErolyIBDIcoCJ+K9vx4ch9Na2bKqryrRvZvIa9Nj2spA
16XIqI6IiSVXbbt3Ns1/lOmHF0rF+CuopPd9lNyjBDJ/M5CrduZxp1ZaFmeQQukwSJx6IuxzX5W2
6zF0YJthoOE+8wg3qUFb8mcwJGM5xXlafXDyPqSs/P5DpPw8ar5geKIjZm4rtMHTyAGP9N7dzMOe
MepDr7znSVV7OdeXRBvrWHQFEDV2rX58AvaVJR6w7JLf4HUoNBdTl5/Xtsu62zt+4l6lU1/KpSEm
JXkrnSuHDd0akyTnYLzdF8RioP2qsIeuI7sB4+qjBCX5CqUGhmktSoh8fykW+4iIlxIzWqMcFV90
CPayUOksqQ4FQZFzp2WvbYxe5zs4nWoOyhKwp6fST2KVrnx+X5rgrcaJyCjPEtLuvDACzakdrTy/
iEGeqCHneD6GD5+WvGRyTPoct4I76Cs8mTMsZdFtb8XePsnWxvrlH9bGd9rwF9h0KvtK3r+rNqxs
rIjvvKoddGH+XSC40p4dwcBMrEj4Blz1Gv31UFhK1IiqSkqax6EiMxWFeEhl4vrRU/SjStqPuwM5
vnU4cVE6yl627iHOx+oOteF6XgcxQ0eP1DWAyBgZWN5yG4XPoKCytbO7pUCFDp8T9NKArcTKspxL
H8vq+0UVxIPyL8PSKZS2fhHMQhiyPKCVPWShe47Xh3lG6SEjwqkLFLk3uytDhCr//wh92NBHe1nd
pr9dCeXC0Vb4szeIUlA0O0Bjav+qMnFP0R+8XadQlAcLBlPk+O+Me62eF79CPq4krGidkqypCE+n
AKYIT6hQUXeA3ElosuqvxjbzAKslNAL3BQzTpXdtCCD3ryJM4GNzeSNQ89zxox07EZuoBZ3iTHpW
HCMrMw6J6bXgZy8WoNgNZh1Mqo7aBXVlo+j++ro2pePHMqhi+mR/1ujAZJbyiYY76cM0oT/frhxG
z51wSeCAZP89k4te30s7QzUlFCLRWMV5ph9tYhllJFI4WsRZOvSgS9OjuSDfZpx2bsyGPzGXd1XM
QXw3vil7gxF5i6ekE65VB39ns09s4HD32xT788TVCXbCr+Z0frxNf/TavBalmUG6e3mQXLLemIt1
W7ajRaA8T5bYRz4Sy8ZzhGdEgwgWYuaDq7wCm46WP7Sf9OyYDOBNo2wGa/kDI9C412WTbyb1rHd1
bD+udav932BmxX7Bx5oHUENNY4aVz6I4TrIYH0m2E9Aceb7KGK/5ZRDACulB46PwW7lZX5W5cca7
El+SgfK+s31fzjBCI+pqbmK4RPO8CTELnDaLtPhMKTYjfVTMagOHqC+3ABk8A1Ns4FbQX59PpEUc
EMnFXu9wNXFKXN8uTSmcoCRyYhLQCQHCtjvXs6m8k5aY2yqaAf6zWm7kKSFJbvdGoCE0L9MXE48j
SbSUtKtHNXK5a5bMoheuImKEvLirc8IiXXRoOzAJ6g7Re6VvmxyNT8iPu83Fdu0eKtl0kNcZBWeu
Xa2BxtvCCJm9bEdigpe0ON335wyq/D6EsRlzxJ0roxeOX2on8LBPIF6De1+vfDTs+XMqJ9ThcGtm
kW8dJJUjym7ZrdT9sRaTzAXn6gHQ78D4e7ky1kuqxrNQfy8Pt5mD7KyEY6BnLmJabGKMmJJOe+gj
Z91tBHiEE9RooNgn2CFB9BCSadrJE0ikPNSRZJVrQZ0I86NV5XsIRdS2uqqUeLsG+wgzu2JeEnRW
I1/HbJQsdhYpNYgvIYco51uXPUcKogt7UVD1yfV2ZmyS9wjaZMhSPS5i+Fjp6ZBQbBXZyI5ldRwZ
T7zs7v7HQqcOLeXQOk4jJTgN1GZdI4X83z+ivq242+pk4BXU7I4t/i2VUJC9ZdCZWSLbglD0i8W/
3zm2rPduT96N6QHs/hs7ZN10JTicW+lI3WZ7qcvEnwadsqRiZpFZFiTnyBnj3DYvGK0V79FxkLk8
XaGxuvpX8S7d07Nyb46xyS/pdv/BAJwaTdPVMSjRVWtOt6uELDpTjJGsWK4DeXT6MPouh5cioKFu
dxSO9xpzcxxg2b6tFB/5HT3UX3/lyaV4AfJU0POLiHJ3jK66UGJlK2dCfOboWRsp9emJIeHCD6zN
B/c3HqLnKrh7c+RFceun8Cd17KL5nVjH6zsDjY6JrXQfDD6JGbOBrZZEAJuEorjc0exoftmSGsfU
y06RdteIl4iusCgyRKHE0QThqMCJnDvvH1UWMMyL2TP+hmdF/emorHOoUyN8jd7QYZEXJSHID+6j
dc5AGvfIQraJ9M0ye4438zDP+b/sNjPULN+UNug0XXQQ+Pw4xB8RgxutjxsS10LpIpBNWTY3EaGU
aMoZhgJO5QCOd404Qnr7QmFTnYn0YY4tVP/6RThbyE+o7WkcJua36GgOSDdkiRymL8DwS3mzZCLe
ZuGzN/2X5vFPrmI1hKw9kTRUqcMWODkh9QzWlt6m3XxWSA+fFdu8yBs6T2VF4EfuALuq7VQSGnOg
O2h7+S5xFtfQ+ziqXajSD339C4rjsrVjShG+fBz3TalYtC7VHtyvxoxlB2y5/XIC1FcaORCio1oV
RkVtOZx3z6Y2+zFGTDXgyo024xN/2tBXW7XwctXRQcYOUZDpg2aRA29r5XjOm6YnMtv57Wr9pUjS
idf8KD9SZ4WfQdJNMA5EGfGP23I2plrb8c3T8gkvGaZHfw7cKoRYYUFcO0omJOYU/P3TrRgwDvIl
qo5DRx5YeK9WZUe9Hwur8+MB1iAift22+76xT4qpgLhwaDy0qDGiyKrCnpKepbnCLekUlFMmOSAH
bx7GlEraPbORaxGtb0qXGK/QTWCzJ4qTOHY/33obEcQQmY/wI8XIWAUNzXMlEYxLmUb0n72/Yyl2
ubrm9T3FcKHkwRXlVhKo2YxIwIe8VtqXufqJhwszRJRRUHx2s4bMr6EiyEPAlbGucv0kbFokHkpz
q9dlKLEwfmrf6tr9o6PrgRKpflyDX5+3GtxcuU6uB2MECD9gb+q7nyq3rZLy2Gunlklgq87SCFEq
MlebjBpIYTQ8Ba9ZTRTOxz4MPZv784zLB5t7TebIXM1WoOAEEqik4FmECEveqXvaXYCmXz6QXVVX
0zaEzBJPdy8lKgN9XuD0R8RwdDJ85qmelMStFNjq0gYDcWMnT038i2rCklAHc0YC0R+rpaZOt737
/5dobIAIXb1mfmyNi9RDE7kR9DAKN8P+FQjLw+NUmugYpOrqVnR9/Tckpd5tKIvtCRqSoUM7e0kA
qcI3r7JGJ7RAIPG7Q6jGkdgbHLOjwCOgDv6ZjCXfznRKDnxPMOnBsjHtGJeDTsvrbLSHGfJZrPDY
Jho036yACfZB54FwR0L3JJrhIaqCv0W4Nl5pxxp7e74vxHXi5B4a8RbTSLAQMbbVuEvG73GKOUB3
GFzI4Yf4zCQEdiM3jL5nAIy5NnjdxQ67fTlW2bSDY0oT66tv/a8gtKdMzJelOEVLvW49jta6BgvL
afDQf1JeZZqy8QyFoXaD6OuNwgVdHSWT9zZX+DbTU9eMlYSqqOmotg9aUFzwHWE69zs4j4DyYORV
vA+PLLnWu+vjmXeXN+EaMeWSuIW/Ay9lzxgYVbQBiBbw1u3AXTRY4c/QNYQYL8Mc3iQY8jcFHetM
InEM2KRHNz3YaMeeIPJWG/lpql/HPMHXSUVi6rNoCMRULMSKxNIahs1UrRxGuUaYcKqCmBHLL+DM
Ym7yL9LKXU5vw+7r5bmLNXco1eVDTcfkgAjSTJt/pz1L2y45cWbMnSQfL/Qf2eXdS+DtSR4qdBcu
Yc5dFrNGVu+tM2NBb1tgXQ439XdbAsYzcjQmF3YK0Lot+LbnR6MdfiEUid85SmyAy4Bc7nYOD9km
EwyLMlVVcphLp0Ob9X3bHUVvQZxL+KT8jscEXFiWWMhuyBLm04wdsVvgq6lAwJQ4bSuT8eMvKE03
yOCxGdeG4dN/lHBtcc4dG96R6aqoBL6DMpfeCOGsegmNBvb62pyLgHinFnKN40HySaI9MCFIf+Mo
z2IieiF8DFNJDeif7IsW9dILabZfhuCIvuz0Ksn2+1RVyXR/WicYR4wuryNdw9ssEaEfIykmeZ1P
xE6IsZluZ0u8pqsxTuf5dCGxyPu4Q1VtDMpwBOzyck0GkN4Z3qYUB7AmVGlvfk1nUshJ+ILqrukE
8De0mnyC6U8lqbEJ42Fnk50M5ztD0xwc3kl0aTaOClrQfEEI5aAjfw7eY88Q8FzC3ag4k6+OHCYx
RuWkjFwFI5evnVnC/ueNtoa7em4z0j0c8gRVgID9midt83lAUcwaI0jYOpUilHsB27wNisNfzkXv
VTRaWTIQdIAbIDXudMRBbSW6vJlgW/kJycT1EqLETVbXLIphAbt8De334mHBED0QiI/Gwf92NfEL
tV/JvGan+QPlDUXtTQ9XWIZicmYEV0qm1w5+Js2DB3kmXaUR6EphFDRrNGpB2/fI+m5GQjsbM2MG
FD0RVYq/1zZXVDpJMp3vfupoDH6dWQ63921haYrsmOYbP4LRdveZpsqAFY8au+4q9ewy/ef88Li6
SQAJaAkYUxb1G0RDA1R2tRJ4meUPT00hTMJWHwnJZmkBdnIhqfD6lhiL1pgpzeQ7hSG2oN0f0S6Y
BoMq2ax4t6Svjwrulp7uvmgelregPiuDXAE6ETxq27v0P4aRKQkYFewWMphp7ymPTUi4xuug9nHs
J4lLxgZZgAQxu7etkILgq7DP+NohpwHMkuQPFsMqli+PWi+MJo56BSwcPIonr7F+X9szQAp54FC1
g+MsSq3KEjUptWsY0XglhqoJqRcMszzm+5HtlApgntc57fY5o4VWPiZkfgUrG0xAywvtT3gAdnrW
8Pwe2YrK8j0GMFgr7gmEOyUDx5WviOOIIj4zJAe5glCzQkOQUDPJgcTAAMA5ppqpoAb5ZuNTPf3J
T52PjCdyMBa49b0nZ1YUYpFvAese2P35OvqhLa/Q8deajVrYQaMTjAySL5ykweNdT7uBOXRQ8yQf
+8NYQzm3zMxZkBwM2Fkf66mLisU1ruLQkVdnSRP6YxmVOt1/yUrlLgu1pXuiTGp1hfpeYirLUS9g
/FKMAJ5o0yrCvVpoIjwYwdRRrv1ZYEjiqXbReygep9Qp6bsNQEe+nVIFLfWUnuh0k6kB/bfgzIey
NIVCWCw7g36ILkTrBkZ2GrsBe/X3GkUhlIH9omhJmZ/4AuestLeNHjXv3KuXPLwPV6hgLw5Fh15O
CRdItG8Zu2SmOKnENXSdVto9Fq1Y9Xi10xnk+ljUs5guuhbvp69ZSQbv/3YePBDmXlg6NWVBvXKb
MffztV8y3yrcFun6uRC2ilYAg/3jyDe5QzVtwhhrkf4fE1E2N8v3KJLyC5lo0WKfXs+3z3yuYNJW
2LEuil7woknEN4EQeIFAz59hBf1x/cTCXcQuogzYp+vuAXqnv6B/iSGDlCdJwG/7eBOgUsZhwb+Z
4ovkm6qWVxEjbC2A2jGneBfl/9vDmMTuP84+OwEN9TfelvnHzSogoa/bAsH+P8x/1J/WNw1kxs6F
kO3ew03KWYa4Y6u+6VChqZckidz5nic8gGH61d6zaIVFfumX5l8aeJqcQYZ2ZXGJKxA/zXuoG103
xbHlUyQx8wE0FLSUk/qrEr1QXD2RfShJA87kcMjs9m9HnfHk+VVRKyL+Rz8MpcVlH3nFM1b5fiLx
CB9mY5L82kbUlopDNAb21IHPEjaph3keprAhouAQahDlCIt83lWRZPb5Hwz18n7rh0+oatLx58M3
WTzd1pAhCbD80eo8k+JSO3nr4ADVo4Oy0rtOZDsc/H/TGaCQitNrx0HHpLIsxuajDD3FRVXFEcCR
LNTsN2O9yBYr8YLovDKOptIrnU8DciUaDUdrUjle3KbTshJg6yA1vYoBNIVKC8PNlwzLmHOJr/DQ
pyB97fIW8v0AvvS4In3i2etcfN8y2VZpiUy/37kctloBxU8wcq0RyBKkh76rcUdWbiLPCxryCK7v
48XTuaOd60NPZAjBTaD9MAWSQCMQ/UpmVFdMHjn5o6bTNKtKwRHLu/DJDLHAB9fHkV5mnNoBGnY1
TivQ1d9w5fbtDce3rVeKkuxlmZH0vnumrKZfnIb0eXewPprt8cDx74+CAkOGwsMgoNO02+/+9XMa
oulBRpZGNDBhPszp6NguOMBF8S3/wqG4NseohBOH7bgoVRbf07iUQQ6gBPINs65xosPrrgBoHb6V
U3ipgr8mGIO3rl1d1z4hPww8GeNCCJrGB3qPGxDuTfzA98zoonk3VHjF5ZY3BQt315zbZs7GQ6Tr
5ItI9ZArsu7eYh9eV43pcMFVR9UZw/glPA7vLUT+XKjSrODYY/wWznlFtTapQs7++ESvVHVXeg7m
mNx1gxhwn0CXoMAWi24tWHxxkBHo1tpq27/FcdOEqyL4Ro71uota49cecHBYFOHoKjiDbOY3uHfj
yXTuE0nrypCf4R3z6PSDDy3lHQOOqzqC8CK5FrlvSj8QcXvi6hsa38eeRSXy70ES0HcV5cqCP86P
yg683n/yxr8Qg3XxsP19dOmwqicudP13fp0guJeGlatXbBo1qAujSPsFg7PPG6/cSd21MoXgxusB
CA83mLPTrCBcUObWKjNqxll2KvX37HecNuOVVHV4O1pQ/8Hj1klx4C/59sGdokdpcGBJezPi2bwg
r1kHeFDB852cmTlMDT2oyg7g8TG8f25b1uIK1hiJX+Px12Z4Av72O4YGbHYBF6XQCD6kOrNN3nzQ
aEyHy7BQLrdPR6rIZaJ9XPJ/NEAfJZ96Fvc0tzhmDYUzAym9OcMsixbsRJzUStQ/zkC8wMkAz6mH
ZN5Dmg7HJthJ3l6klRo/kQUP6Z39+EYaTgI3whH4feHj0lVi7WPCcBAeu2F9ueNpQjOPEaO0CvnQ
PrSq7TrbzscBual81rZpGqWxRWVL+k0OdRMb2cMPOuV6k3BtorlZUZi6a/qJGiiB4Q8gx2SAnG67
UYZb0ZmlCnwW0EuntACcebk/ItR4Ygx7FoFbmuH071xnmDvF/omOzp7gidmcymkVErn5NGXwK1dk
D5HCVNPqkJFU/txtYfFuirEuAIynOrYLc4heMm0lKQkXvFTQei+oUt7EVohfLicpi9T1eT75/zun
Iudy8dsESU8fzUtYh47/WTm6F/Kxa8fSMZFiXCUV1ojJg8Q7l8llYbP65HlQC0bN+18DvZd64KTC
D0JCQw3sqiYztXYK7Gx5R+r5pRhAnUknUu8QBc1nD31V1p1Jo99UMpa4+zj+JqZiEXagTQEef8w+
j5GQbN6rpKR0neto8bWVEWBcDLQ9k1eVOmbwuUz16OMfv5cDfhqFtRzzp8ImOVmAD3kz2hu8pOCp
E5rTa7+OOIdp5a635ywjAUz504G6SHo6EfrgPkbjP8RUOfZxfQrSaHzE6h2LbsjQ4DN0W9vGLju4
757T7M8Ftb1Jos7TqBnr6aaA+zaD5lzixgCpKEYU51gqcUtG4L5fp/oXXuugutcKPN+6VM7dyycr
v8QFPswjntbuVpOkV9aLdfktKB5E+7aMVoBs9N4ON+griAa2qnLIUGjfiTj7bM3JYZfysWkZN/1S
rQvz+ff6mWFSFzllSxWkdbj0bfU9L7+Hh4+YNRBPpNhPf+ZeCUUlGoFEGtqIre+iuIPZZF7FllL0
hgrgrHz3etO72VOveVUBcx1UopJuK7MJnL+/UwoI8YIRYR5+A5LPvxU5fNoapYmlF+c71arjq7cb
KCJ529pZVVidnSFuyYSQFeppENNMhajrLGLuLyJ7s47De5Cpe/QRsIp4clOhZHGTn3KCuqoHWi/M
MmU+zNDEwOf6eyiR/lZJFdjgzoYSVz3Knic6sQZiqFDfhmBo38hZmcr37JiErCOpF4v4sI1DJyfy
YgnIoiKkyFyyzmcRpmt7GxjgjNlMY5vr0FdU4mzM1cpW0NrLslRDTg44MCwBODNCiL/bssjMtZ7f
f+5Fz5pvHsF59bjwuLP7d3D8+lEh36kVCKnLidqWH9pcVTW7QMXo9xc4CY6pGoLurE99EsC0BXLr
/rIdTEfGSSfQ5AVOvYz9VM7/hQsLpM+C88ImNvMZW+4IjM3ZgL927dn9GI8J3P5WdUAdQDq+LS2Q
TfGxZ98ixkzP67rL1Psr59uMBAnuaSc2VUAWTh7Bz2jwezQ4n1NSWGh/MvLCMem1X5yqfVbfmu5B
kTvzo/WfPHEC4md3u7FvEMsIIMyRII3ICQWs3V8ZHrMpvb993DCeBlk1OT3kYdngXiK+S1FzKk1M
LpZyzKiqTo3KXV6N+TbQEnQ1OjFWF84y/206Dz/8XiPKjk4LQz4Zd9aJ2uR/aUzQxN+NiUYS/G9m
EcoYsQyDsuBViyl8coHNW1OvDPeCjwp3YihAzY7MFrAGuYvLwCSjBxqmrh2pdBgSTNXgkZg/RxU8
w7XkMNFL63MmuVB06KMXlgrFHLSSUaFZBQiVkpyr2aB6RCRo3uERa2ge5obiSI6PQdneYDw+1tcu
mpFSacTNWzjgzWIXOs9wvpJczaawSgDhG0/4dzBJO+AH1/9yYfY0oD3qPWFSmotPHGAI9iySi0Ws
OdJGkTqVrGWdro0OYquhBgXdcnQqgtIixgReAh7H9NE4GGUegI46AAquNIMqveE/D5idKe0GPNAF
ufkuFSA9P3eZDWq4X+1pqU478AhnpWryMREeBzZVFtsnzoTxPr8hDEVL7YSs2nnGC+8X9VndTFs6
kupxINM6HlvFZ+WYtpmREI+RrV7ThV6irwRqVoHz/gc8c6g29gjbnAa1itRuOqesjDCAaIH0hnR7
9jOcmNaARagg/vvZw/ZCnFJWfO4jsKWymaORaQENFgewjpomuoplB1Ss4y0Kxc9ueogshp6Gav81
LVDF+SJ8qS5502Iy+KufRHMNRMc3GZmS1wrc14yLumNkdWNeNuwYih5oX3OzG84/VuEih+q5Hzn1
t7aiVS21DzrH5RQaM29Y6WSh+sk92XfUeZ/sU6GMx42p9NSlJVmWv0sAYTM8aAW9pdJ/oJ4SdmdF
9VVDh/nfVPwLiLzu7tlvrrlFHnJ1uieaEtEfC1k1Wy5qR5+1aF7zCnHasNmwRVY86JN9NjBo6BuS
Yk8A1erkHbuQZBPiP2ljgeD2KbrvrCUQaqJABRq+kPLjMNeCKden/rdBAkfY9qdWLC3F4nQIWzHf
mzlxr+6fYB6JYIgSYdhtn38CcC8fwsDXrEz9qTUoP9Lj1jec9lGZYbLsAHrexWl+PTNmOn1xWXOT
mhUcsKA+i+MSolBvACtEcRDgHoJW64NYSz+Jzdw3tAKbaEvump1FCxcSYcKCRF0NUqB1UmGNQKgI
C8HcMnctDJsNiToX+BN9eEk8cWzh4R3ottaFEABVNOGUHUXsjXIWrvxTK38ZhdlljDxwv5ApuD2N
HSS6LzVMxpT+cu+wF5QkTVSIklc40fKW+m57w+skdzepP1+fLdjkeXrFwpqw+ElozCJLMEMMMkcq
BBjiGS/rCkmDowFQrn2S3Qmg4bAMkCTwSWdobhiZta2CjSZsNbspL7s5T7R07YWWYVm709DfXUAg
GChKqS+fCRyNBU0zpuwFjDViqIWJaKcj6+jZrwqSZkiYhK87u30xZtbgCulUF6dJ3KIgJp2xKpzU
RGtWRpttRtxyBLBD8dg1LpCkIqcpW031xXQez9xIaju0ylBISnl5SHOLceVEK6F84fm8lnW5IeRG
0FpyIrIK2YVUzbhdtWBg5ySZ0D8jkEy39R1u1QjYMDVer+r9dyWJibI+5eKcGNV3FKjA6wsBpEBM
Hzpqd9gvjPkvVuig9MbHIWIszHitqRnVbBRSBK359zfakagNLxTS/GxEtKhzeuegcIGRC6KYxtEs
Ny3DdUv9u4G5C+7aePidj0z0MICI1aPmwVqqHXb1O60EM4VLfv3pIU4I7Mxq7G4cuzJdwKtOLrtQ
coDpc/51AMSNkAByl/8lz96QqpeyLqT33RaiP9N2g1vi0lowp8NH9/iUPf5QRVUf1PducP3SQpVo
KUcLHVgzDaAqqmomUJPGKsjLR2GD03w/Fq4VozgM8ijh8qIxdtiFW2nXK/G2lNemEh8FtWCbU0We
wU1+kVkGp9mYsHMCsKS7rpW/fAhoWu5qrv3WR2YZt5JgF+gtepgKj/4s3wBG7skpkGNltarW19/g
woMQhieoo2Tn0vwpfvobb8L0nw3sgmd9J0MmjMMMOEjfk6+82kQ3NLGpI+bmpihl8z7O6z/L2RkD
uqtL2EdVOm92bCqILv2B4YDPAUyEdKsPA36Uf+UJrVlUMm16qbtbMNWe5IyAonx/rGcngXC8kC2D
ypvgT6Q8Lc5lFTVniFI2B9DeMYfZ/9XRY+gUU4hWqP96QEvqGclalHae19j3YNsL79FgjpULLINk
Hw5v4hNd5wJCzGz2iNkYPy5fEju42D3sBRfbnuU3uQe0o64vLCNfkw9f/cKCA+oLit8es/ZAXP6r
VwE9x1p8tHc9RO64bt975N8t08X3EqkELxmVWahAncYzrFPcVVPsEIcd5jsfONkTzfiUg3zi56/x
iuBLByD+FRfmQBy+Dml/snK7JaEjNgerJ4SvxoPILPGoPYqWasczDvR16igkGvxkuHcBKuTajx4u
nMujV8cY4lVQxsoNBY7uCPVcF9X/9O33vAgQSa0cYswN/sB6XvNW5JomGPMGEf4oNbo51oqH5Vvp
LnxOEqweam96+xlVd1J1bUiaufQRhyZDnI+g4RmmcNH5JMVdtP54rlxXvkLzo/m+zppgD62XMn/h
TlOuPlaXJqrZ424Xd3kzQiDZZuUAmLM57ZeGxZHZUjOT76AOsdtb0zFC0ADOHX7kgV5JgqVgF2YJ
jIf0GnPRAU/d3RjuiozQSv8iCl+oGiz8UhIoODSZyVHpIgJ8YzB3iNtL6cvVZbrJCIrwN5nGTHwZ
7B6YTqJJvCuxwpuXHgAYMAe3fmx96UXfPKIkSaZetJpzN+tQIgeiBQBII+TboiCCVhR14U05gHqI
jfLJTm0w/cJx5wt2KRGnbc2bwACntZsI8IdNhI58Fh8AEt++Mpwj5nZZuk+bIRNLvzUjEATot/pP
GPYJ+7hP0tVv9SuLS93D5Kh89fEQtK19Csjtf9D7jpyxkPEL34FXcW8EH8CzT2VW+wXTFvPxan1V
aQwU8F/r7FgzN0Vd8jZyUH+41X/lZA9MUVOeZFexNUWz9sKwz7eE2lpwXQBB5O4CBzKjfCx7AtvD
obCdDi6KSS4fPVtXRlJ6jY9fDQuLHcFveXDLF2J365YqPkbcCj7p7K1nQdUHz8W/TuTMsDV0kFhS
di898SIEjTUJ6IfsaDSA+IfI+ExiRE7YYjyi1UUAaxyJVoAn00TU/0v0IQ4pYldgCw0dsWjlsGD6
sCv4flz6l99Z5Z2/PDUz0l5QBrBi7xSSzaCY5qzp0XFS/HMxOhIcTeX+yceyo6GqyQi3CEXRrQUv
LRIbhwmHVnHfiTUxQd8w8TTeg3tR3r05oFejc/BuroZllS6G1djcILV0BtR9ersx/4SZGse712fJ
V+cY+X428T4p+UEuomU/HtJ/MRa+lRMqrh5lR4jSsFCfixL40WafjD3fH+qLHxen+uK0wjGCQxYL
0ul2YOFgMMaftbQ3zSNlz4O5xWUt/yZ4CLwSetEjmujpYf2Zjj0UXFgxcxqnlerovagcGjv5k40/
xIZLie1uedyd6Hle/l2DVFrNTHbdABPgnhp1Qp8dEvDdWm1x1+0ge0T23e9/mS9DfqRhs9lW3xYD
LfKMeHJP/IhIT2Ul46euSyD6heroY3Oq5L9K+QbkcclPtb1i+Ym5sAIPFMAQZz30KkGbx7zdjE5L
6OVrR6I9OF2S1UI+5TIh5G81rIhBCI0Nhzz1YLXAm6J73wsqGMcYGM5+YS5OwXDXrsKm3gGMtDZh
DPibQ0YdcSQBhgddRsR7Xl1+cg8oaCgQ1R5EU9JkeL/0OlCaMsuS81X2JOClz3+hVSD6A0/GEPyg
lS2gSsmTI819A+U1H7CfCaGNAZ/36cMVmV459h1twlhabi8j6X/06H4/VjrTUcBJQgStp7rqPy3y
iT1QnlXlblYizu5Ygh2h1yZ0jOXcAN2D6oKB5GD98qwTp4LkphIpKM1AFiXnEkJbBCdLo2y0Fzr4
a5LA1AuHT/Xv1/Mn4bdoTAepdj5cYIWU6QK/FhrBsRrPC63LTGmieZ6lHHL3SdTHYcfhPgEuxNLd
PCp9v0np69VtI+VebdRHWqJv4j6tnZcLSebFjJn+wyI0wlP7BoVnIfzuBPQXm9Bd5YMk/B5zJGOY
RwLNOrnptARNgQ+SCHopyKI/U/NnXOPJ5tcJQNdeIfTntS0IBpdrengdALCHncXEtuHlURUKDIMM
JdEVYHnOcRPOPI5wtJGSG8Iva4t2Opl5Qc+d1vClZ1KR7aN6LLDVwvn4firb1nh/Is5Rgr/FRO1Y
PtqGNXt9emdye5iU+ULqtm0V+kwG+uurD/e5crNQ/V8fvcYIIHCnb04E0z5kSqTiLHclHY3lHaNG
slNV7Le+2If6VGFqZwFNigPDZ1yDdwrtTGyjJUniiHb4DnkK8PH6RaJcC/GxUY7QizqXCA4FuCtP
KItrEnykOg0iQ6x/8lQPUfS0gdXO0bmMgogckL5QDpOOphF5dQxsJobh7E5ApyHBG3raVMGDcYcL
kMwg8Jll9+pXZjUFvTQjDexoLMIKaAy+3xyn1cOzngP8OH8ggsKirejesPahqP2CVjSaSTZtQIv6
sRamsdXWHIhUufFGBBNsPIkIleQkeLnauvM3/17avsqhHWxMlKwK2fiG5+VPumEVUYv88rLRrxGd
CwK1Eu6wExVzbm3qHBO0X1GWMoetyt1/tlZrw3D8aZAWL7UcNnke6SMnD78FOAahztYctHLj3kUT
NWMRi4b4/6PlxmeS1+WTAO8+ubYcpS9BgBazbJSgA0SpUFB8trJjAlOnWu1ZUkIzuM2me/G+rqvC
gbHa/re76PMNQ5d6ffeIoIjflTy9Qqbe6xclyOtGxvEFWLLAhkrZqGy/+G9nptm+Hg68Ms7t2xnK
S5vFOZbXenHUDlRLUi2n0v2vSjASyNwiiQKdSAHIaWta9GPvzNgKbfRIbaGV+6oxP81NqkMap8SG
mofFjy6YC5+3tSi4pQRK+qNEJOItbgl+teXP8Gaaed6Lbf82Br/aysr02Vrz536X6fBbVomNbsHV
atWTpgBUlpyuFd9tZS2whyC/Mb5tv7Pawv2rABdAOl2/AglY1RlVtVNJr7K571xhEsLX6HAyAsAn
Bs6a/lew0OyGJ+h+XwXESmhnfxRyN7v1qTMtryX69ekoD/Y/Pm/Ld1pNzDeFLonuuxEHMneq2h7e
b05Uj0fwwSoAk7QsNhzeRn12PrMoXvlMGHUcx+S5hlUuVxoGcNyoN44joWKqQ9ZVgwRnE4jKLd4W
JLXPkB5CwmOg29uuJHPWIjGzM60eJyxOdOdJKchnBWhHsZVb0HI5Jgv5PCxV4gvWXtCknhvGAiOI
P5ZCYa6vpbaZcTprOrPAeO6634YvQTxU2rk2xg1+iLLbR/mo4/8vMAcHHBFwx7Yb8mtV9hBqKG6a
t7Hxgt56DXcYchGySs/BD87Z9kMhSclOplh4NbiMVrPJY1kwB+FQk1AWDu0+fZZROwYNqpTOpOlV
o3sITbXWvQwKVTVcLyRB0ZsdmYm2zxMC5HukY0NhFwc3DpRgm6FhZhgnxuM+AtByBVxAS8e8aCVk
FSYaLfgpka8eyPcpSWIV5qdl4IX2yJLF9M6DZVIHlv5BQWnMLCkZ+/HNTdWGoKXETBq4BcmgK2Gv
5xWZAkbJ+fe2Co1+QSBPs77XCujtw46TLiXArAHqR3qtK+SVuBr/bCxM/kcW/Cp45wgfYiHHeKMs
RQ4EnFUNxGzfRfwn2cWaYbqDJolzkI/yoGnAy1+15vppAaKQM/hrGLcMqNxYaG36MHr2Q0virBky
ceLSWbNVnQDbFkk75otmAkpCuB/NyMo4TA7FkTkoupOSsmb99+yfcUikZ2p+Ek3Q+7RYkO1IKfqe
XiHxLuTZCeK454DOVMgRnnn6qZOl7ZUA5klIyB8qMMGFY1N07uroNPzNeQPdJdXlw/KCUqgWNOz3
5BSMcyynaMDB50Yu9yrapPoWI2ycVlRP8X3PCwPGVr0a9mKFkjPE33NOEdVe63Nc9KG2FUdhCRtB
7gW0niQ8ncdZjVdI8WFKj22tbge3u9KnhI2OoRQOYEtSBs6+Et+khvj1Ygk+wCSOOXRAxY6lTYEf
QwyaViyvI0M6ZS78yy5luVPPJcx7qttCoe3Zp4UnY0dZ4JpUAnOYOR59ZdDvK6z8/a5LGOQpUwsf
D4t0/Gjsv06AdHzA0My9KoS1Lfxz7HjMUW3QcSxrrqvXnuTMe2VGn4crPuVzfNezzjyB0RWUkQnu
uVu3QYMwYcVUQIgUAEJi8ViCAPqB04yTsyTniWU/IR97q648COZRcngi4lZoBNwkXD2U1JjyXq9F
7m+CdX69GT1Y+hqwCEAsBjzVVorGDGmra3kGlAQE7SEiKgQ/tT3gXtCOIUX8kh4meJ49lc7oHAz3
Femu67CwuZ2jMicMfqkFezp5fH1CcjI5zsl9D/YoNzzYMgWEpVLKa7JOAJwoIHmw/MISIQvxtLdn
ewVVXfL1haBBhU00WyIZ6edEd5L5YM5Umi3In6YGbuOkwvhHEa+9JA8VLB4Ih20DgGKjC41hQVj/
GNlizQ3BnG0X4RCW5safBOAf1b0y+HHLl3Tga/YZk0WWJpAzh99U4o65zPfEwFkwS9L8x39PUDtP
6Uzk1vplbTTxeH9eWnfhrMIYnMG2QjE68uiCD3mab5z/hG8TQ55gWLdLxMHWVk5QgQha9X6E9UZQ
M87pn/L8zg5VenbH8UxSxzPJScsjFdzl6Qjw5/5oKaxtWkQsx4JF5H2U6KX4XYSSP0hp1m79h3s9
f3drQUdKt9DSCET9l4w1W/DrBDGPV2QyzWYPs7i/qydOamjIhaXMej/u8mWQm50hZSybZ4KZmX4B
1eFA6GTwM++DqShWeWrfO16iykCnfwIZdD2W1Jb+PjpycXnveW3Yqth18f84pB96ZdLSCgQYdpht
3PWmAoOnVZ4BZvibPKcS9/KqmoBQAq6IE8qfeUG+AW8YgU1jYxASKamQa25s9OiS2vR07SGvyM87
jDK8Ldcmq9wYo8OI/JKofQS4qyPq2FQH3skzdemr58DjsOYzsUYsjMmFnJwSHKuipKa8byEago1d
mmm9kYqGfkktqNifeeRuvgJvo9r/gHPt8ubaDQq5INquNw/y/o9NG1r+b4ShvWatyWyu1og7Bk/k
6kWxIuP5k2BGdeF6F1IvvWwiTov0xu9OoZGaJj3p3jYHTrWQRoF2kWKICD+1QqAENJjdrlsqdpu8
2IFanxDpXtw/1uGwJosHlDxbpsprRNPmcqBUAE00zahF7sMnhciAwhKfqTwMyRrNxhC2Q92U8W0M
aoCHoe9l5TepcY64rU78t0qSqQ61u+Ygr0TZ77w4HCrAlGI6ZY5Aq3maNWsBMa+30SrnbdgLqe/5
hxu6tWXS6C7wP7SUK/vbFn1/YOH+ERJwd6aN/HBc7qzsxj02GtPRyQqUSxlHR/x5eEhMT4mADbow
N6xlQQD/BEMesOYyTeynNT6Ww5SOfadJnP4XapFeKYRlJ55wNbjdTuw/Sow46xEX55ZA2TDryi+S
sd72SBI92UhX1k8xLz4QxbhRD5FcncbWaZ4wDE/Xn6vgJ7xlaOLZ7BO8X3b3OjanV/IQ0YJmss75
1FStUj2azevCLT+GIRR4Z8oXIzNQ7y+PJ0HVqnnum+77Iz9EamHmoQrmJlU2MxCnC3K7VBIEq5fl
090NdofQB7cZNzqu+yTgFr1V2BksJQsCFgBdQA0NMW0BbMYofZHXnRbHrS84kFK/NzY9D2KzeON6
InaHHQuZkQb4nvfV1BW59E1hfaOVZz3fYE/aibf2SlQFUg5aJWOAZrhWnXGkCUsbC31s17m0msBz
HsCOXX3YWobo1X88mnQkUCZx5Io3+B+MSHiyyDQCB7w/Z9YvIDzOoOO1QCBjnOzqO3E22X7vQT9E
bZ2srBBH2NEHMQv2NbxQ1XPwNz0Vvy74BEUrK49blGWEBt6n/qd49P+vB5XTy4AVgSgT/FU1XmBm
0qoLVmnwxxMuIynzusrDUsLyfE2UBiC+3D+9jMUAQ8Hf+7t+xrSghPUe+NjoClf93EE1mVU/WACR
wWqxNHfdtKmYhtTVhm/Qf5hEMRtph68p+ACk06wpatMB+16s+/tGfN3K75S2ZTijOFdezncWXcTj
IiQYaSlTiKD8WxSTVi/iKl4wcWnOWbQ2aibSjsPvBgj0tmbxSwdc8l+0e5sz2RVTz8L8awXHaq1w
xFHAHNpz4l90oPIEzdkNr6ZIGUenuN7EFeBpzC57h33M+LJjNKyJ+kNYyNs2BXJPCOeKcUEIKZNO
ySkMhLjTm6ifYdMjGFmGHDLyLYy38IknxjyDOsc0A8Z66cgjH3P0kD0q9irQ//tCDFLIZgbCqzTY
ztNayxgA0PCbXR/isNcg/byL6GA8q7d4hHFam5FMhK8CcyVEoIvwO3Tpv+7xALZEo6jCenIOTdQ1
NNh8Feh70dRECXT+bQwghC1ttjFKUi3KHvVtYuWFyJeJ0N7L754MUE0lvrZScGQ4TyobsZFKotEv
ROXwfnth6tTjolj8Gr+UugIdNnAz4IqvCqih1HAiv9+OdJYnkupM5C76PEwTv5IwfHRKoocKodTc
Lf1TeXJvx0KC26KMN/49j2ikKHsrN6c9AGlbHRQZnqHTaolcSr2ipZtVAr1cx3x/aE2Lnc/tYgcA
MIzili9fBPXv2tvutmiXPU7Za4Ry1Y93aZMSFfkcuClPchN7B/UB6fbr07CtTJZXSzMAoY9WonXf
u04mJwSTrFIP1qmQjsFBd6sjN6lb70/go//1JRfyMCTpAV5RaD8E3RNw11+I6w3wV+LUGv93m4cV
ATuZj+JLcR02xA8Tt70W0g90viNgiT6lNzYRrtm7VWZic5ys5eMR7S5AiKjKwZ8PsbnkA8f+wquj
u0BkZVt7AxyMU52E6ii2tozApdot5KY2h3rhw34MueEcoSOiR0MfIomrqriFplWXlTXAFi/keOrB
DGfbD7L/8qONztqmbSoYxPPb+VDfNX7eetwAVxf869It+KNKjlU9LbwgwsnBOppI6lrp192Y5d0+
iFs4m4Ix4fw3Nyir98hf4/OR6W6MpD98MmVwIEci26Tn6wnAuEYTc+XeKooM6GUBipF95KshxyQs
ddDy/06h+J5/QpDCKJj2WUIhuzKZBPw9j27ogfw9OhFfo1hTgBwUg9gNv0WShcb6BAjsnj4jOrID
Pt9p1BCYhBmmrTelNyD6nLjMdytRmLURtjcPpDd3+upmSwT09al58PdvqZ9lNHj8jb5ECwLVbf78
bC4+4W5n8ywmMHPnQWAiMVaxfwTYspfg/9ugbDK/ijcawRRky+KodTwmn7euEA4v9xL4ZdMIV+uu
HcfB3whxIXk3yyksldO1UZ0PXqaCCtfYttAwnNoLeLNHY3rogmykxSnO9gnuSeZh4bDr8aSkGzrR
BUarKcCLJboUZyhGb5fG4yV1f5cdtzf3yUpk0R4X/KZPmYmsN4rqzsu5682zm1YTKHdeQoACx04G
kaXxXdv/9lo8DwJm5QsXBCaT52aF6MFxAAeaJFEbn/5lb3DzWEdZmlQe8OATVoitgRXFc12kZII2
EMW/HAUGhX3T82UikDC+xRWMUP0F+xvgvPIFVRhzlzThPVZwDvkT/v893eKvHy9C8MUO9bz/2eLA
DRRCTYj2cCHSOo1Ay8oikFFWpMGUIRGjO+oRNPF7V2qfjFDjwvg6RQRvvqWev1IBrsOcwmgC1/qD
4udRtwt2zOcPilrGx029MQUjEsFOG59TqCYL15VkHxIXcQ/YZYkubUCirvrAVZYLDjExJ5kXBqW8
lCmCE0Dkwv947XvNeMbEW0KAYSNk0rNl/5+Y4Ae4F/Xxdin/J3sBcINpbZFhdbVp/H5hApg8XwbK
rFMeVrmNLUk/6PXILdsMa1ZPbeXUWD7i+ErTQbPXyZp0eaovOGGdeEzyp7uWR7uWcMOZ4ZMX6nqC
28HC7Cfrl22KdO5He4mBI9g3cnQdTAaPSZtExu0JQUxf0NkcDjPAwB14G9OZhIGPL6drXzT255tg
p1mch6YzncHInKLY+f8zINtXypbqxeo9desGOXDRFwaC4IvhAzTEJsSYk3O2nwkIv+97Ev0Z+Cy5
TTfHY2H92U0Bvnyydvlr4iEBD72oL4NtnQDYzsMJaZsqbeaai7mJjcrWlVOzMr7hLfWivtyDR3Qa
RcigHmvDFsVIpkPBfAuWXWB79w8DE8VqIQLTIMg6M6uJRtXHeeA10BfC5pcGiUtoUOwa7Mjk0Ll8
5DVvfbh4WcP4vEbF3aLyanM05fsz607rNNFz4/jKQKR6rnonF0rIuYgtNBwfgddsJBZNxGovYcAs
ULN/452ZtCcta5Mop6b9oma7M8LLypon2CUNkIHRrcjeQv13mHLTGl7+bXNRzi/VpUmymGXqHrmP
ylQarc5XuImSH2LWQLljuSCriFWlv6gzo2ANBzDA95ZVchv0wwnPmJRib4MrLlR2RvGQDaVTlIZJ
iV1abraBiVhtARBe0ULVcwtY13c3O43RLw0WQNNr9rUSmN+pqKnZsH3bbmPVl+7NgxZJ/GU942hk
GRgYwrtBa0nd8fG4Rb/jGs88tWe8FDqnmurEJ2cP0yyzSwysfHEagJDDMVjYOnKwNy0Wh6vxPFpW
8Q8sT+1txCILxYXntwkuE9JeuHcZPK8FwzuarFZarI8C8icoNCLO5ms4vBG+Bls5QpbQRmE67+ts
tCqVjlDm9D8GeT1Ea7H8DfQyDyG49C88+jbZu0KiiO3hfXBCnioTclI3rFqwGii0Xin9Hs6pqBaK
rQXvO02DeLcZymvvuaqntPQ7u3gx6NokOnospxebYKEgXB7RRICC8gsLRQaWeR00cSOnnVn0FhAU
0sqvtVYbyj5Xmj1HjaVl5y+m9lYO6Ey0VYADckdkUiK0LohSJApts76qxANmpdLxfQ1CzvmP0FEK
auBgl0dmTE/cE9d9kn+vf7bC8viVEkkWiXnYNEKT1D8kNuUOF/hB54+g8iw+nv0/3oRfkC6mnW9u
f24Q/tt6lqTr7lclMvSvsHE6zz9Ks2wlMPQuRgyZbqsoUTqDIV3fRGj5Abl65Ij/IGKZ9HeSOKdd
WmcSxRZLqpXu528p6O4Z0Dps6yE8edLCDWzAyGT3ZQ29/VJgpIj8mw8BdHC3ioG/rl+53p3MBQe/
9KVQ0y/76eJqFpgoxKL5BnFoT1CpptNnH5U1GhhAboOYRfCUHG60dxpZwbVs/6QqBHKN8bk87HuP
9ow0CAQ8KfRW2hTef51ZbBLUKNx05W8XB/NTsjoKpEWVrulm7MxM0sP7BRHys9QnjepKzBlfSKAD
wzK5nhknfojEcDQ89vLP5tHKJkeJHStsnqyFpTB378Omz+7/e+BVUDvrbNpuBbw7LSnSBRidOsfN
TxVtCQ3w0dxi9/DayLc2jshDP4ag4/aSqKsw47REZPhJZ4NlohkeCtVQyx3vEdcj8RdQes4RpUp+
9Dnj/ZdzRZ9Fnb4L4N/dtnfWvSrjxV125M8SC1nWEyM31QiyOqum7OaVa4Fi5OldUmVI1ia3FpzK
lvj23/40RaILIWhmjeGoh4EUYG69c+YakGiJNPqnRBL+aUEndmxmt9RVQwBVbu9xVdvp+MadpC9n
zHz18w3VPGv09K6EX4u+2ed9YXTqVac275xtJsQp17dflD6W6/j/7DbRS5Zr3LfYF4brMiq4qq4o
dArLB7s+QS03TH0NW8s6kurWcLyMtF+V5D05n9gYGJnRgDKMU3i5Q0kH3YfPy4Qz2aIRGJk78phN
Stt6GBmQrLW9MVs19WtHi9EzJ0yaahUsX4MlK9pDQYBSmrQCfquRWkN/FTVghygj9u4M2aEMvaxm
THRP7Kgz289vtcLTuU047LDDQn5nksbSC2zqY9PYhr8N9CBm/MMCOuqtH4O3mR3BPjUSGO0kqC6i
P7l5hKqtCAz5bZou/GNOrv7PA8kRmDtxGa1OYBEHBr/xh9LmPXtMba/4pxp1C0wBpDvyBIKo0y5E
OJNHI/mIBFP/0+Tce77AHt/7axnWSjkM/kJuenu20VtxJ9LRotb2XVvq2FmIPboIKd41sJ5JiGHR
2q9knv8hrUxFRil3h96n1ombtL8RgL6EnRSjWSBfgyaR30MA6ibAHqMyjzH4kkjXLCluX9sFEDGs
Y/E+ek5PH+dIwUfqg1BCiJz9ZxvfaMHxg7lQXE/vh5fyN9kR5CkLnCW9Duj5HwgnwOAZErG6hBfr
AxNeIv+s04J4nXxgaIbSpr3Nb6OIJqISFH8CqJBs5JYs5w4Dz8xeaqr7rHk1H7mmtkuZ2ZkiEb42
M28ZFqNOXSDwLNvw94Pykg+An5+3T8Vp6rQKf0/5wylnuRRKtVC0YxFTpf6iDMQuU8t5qJiYaobL
yydYgk/RIFyOu5rtMe5+uS0T1e5CFjuSbWUmKQlDvH3DFA2s/II+kp6v0FRgCgAxAuNYLo0v012j
MWz3SG5ABg6i5uX10u733eiwg4veo3OjPEKQ/hWBFLPxZhcc3eDPTxaloDqNHNqa4c4ntXs8TKaJ
KGIfO4UE2SCmuROYxMyf8O5yHEZFLiSrNsBGXUsazElpbx5pHOSwMrAQcor7Y61bjyC0VaUe7y2t
5ef94Gx2+sQljB+FmKDp3AWTUCzMFTPJzDYMTvZXJMhKcfqN7yq7UtVMdnXl7BF56Dv2IilrwbTx
0Y5dae5Jjw1sO2GyE/2o48OEbJUaenYbwchvRWCp+DEp8N3NZCV3zoaK3SVvJe9YLgz2IQVWEfq5
86SkMXEV+lNI+sqq0uUaTBugNzEMzripZZHUZU+R4nAdjLcExDzbn+kxIKME
`protect end_protected
