`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3488)
`protect data_block
Gl6NzlCyJcPkOTjtFIFgPH/S4NvvTIBME8q0mk6Zf0K/GWXztJ3heonLKOGMbkEmQlXIOD811j+Y
lyDwmx/KMArGNaED5Iw4anpShibvYwclUDX7GIq+OGCE8iMMC9J5gz9hQBjFFRPay1mRau5mSZRZ
HCvXDhxvMTwZ04W4XjAhUDlmzdr3Dy66gUGF/Nc1F8wWsqPm78/Cq9jchwYsoirfhjW/5A2Ih92u
wF+NruqkaLxvSBZ+OwdX0891FZ8Mg3G2dFCNhncdqwf3tiw9o5cMyIqJlMwCKGljDDBPda84i5lI
WpVxQOzJtSvw1kg3bdxFjVtTuFGSop9DLs5JrhgKq6MrDcDHAywW9Qk6uRbr7YRR5CA+mr0cABFA
FW1NIlciGhe5ZMFnccKTZ7JdioTtFYm9XLihxBRGMLXM5HtW+wTsb26/dRWSc+IZ7RZD7Vf8cAnT
u+ZEU8By036fHOVcA/v4sKb/uKwQM7OEhVE6hhR4O/WrH2e1BmJo2Ra3YOqtdcCXL+izwKnlOZvx
2l1JfStMMLbQHHVp+SfVVObtbTTuBj0xGF+qKFYSiz3EJqSCi+cbwibJR6eUvYhwLPjhQa1n15z2
Iprl4i16UlDoG+jbRqwZcoVP65hWLh1FnS7qHClwS21HnEA30hGl54HHiWGr/rtDRk1N7+8OS9EF
nuvgZ1Ps9gHhyxYuSrzP2rTfDbRvAnYY9aj7eW6aBPJ2e3y7ep61uFQhSvCljmxNDm6aSSO13BkK
0XawJ42QWAuwf89zftqSh0tH2jKbmMIVFEa4UIZpYwfd4qBleJ5KskK/qjuZKySRox9W5PsOd6SU
eUxboAIhCSY7kRVogfwKjE3YWGPF374YvX77jguZX6FZNVw+BG0rfWA6zMYkF13bzy2AhSd4l9j1
MnIEpwpCkATpn+feZiTSSrJgkUDSLGGULyDsmm7+hmHOKi2HPNtkV8p3Csma9lcdDYlMSljpUJth
oFeM8jQ2YbaFKzVqky+GJNDP49C5liQ0ekXj1H7IWpH9m9FCx7rW9BHotTxhnH0wcT7WrBmqz+M3
D7pM6Rrpy9vAnITtLm8y7el0PzDCPoy4fooP9x/mG1ubMT7IFTxsP5IPM2CqDxIK5GBnHb6tOl1U
BjMAOf1jXDiIkkIGOw9oofA/6idEKqBeJqZW9sYf6lYaYrcRow+PW5V3jFm1bMMCZHN1UfLGjROS
1yO0XO1LryavN3jCcD7MVA1RkVsavlbeCvIWJDzn1rr3GJAd+DxPOxF9ofMnwlmeRY2hJ5hhyk+X
D7ohOIl+uRQ4/yq9Zy9kkSkYAfe9Cl4Ll1EytAAZ9tMO3RUA6SNMfmQCSSRyfTw/xJOWayyN1RcE
1FcR60W6+4Bt/GokdgTre2CQnrFW/uz4VArROwtCymd+tWWbUcWwHTxfLIi6CNzIHYuP/HbuSE0N
sV1Us5Svr7Sg03GJ0aMLk0E1p9FnNpP+eakz9nL/LMDHbvvc/4cD25p9WnZvbgpQpZU+AqaR4kWW
th5i0Qx24am8twVzyeAoXlxlyY2ETX7+yDXEAD6rNcgh/dSblJLYsSbLAlu+V8EUGDPkoXcfWakM
vko5xywPWCN+GO7X/yCRKjzUymEaZcm1ESM3hvirzK7mav8xUth1Yoprm53DOsEfzNCyibW60oK2
gZ8BkV3ZNOjN/AuOWaT+TRhXJ0aKgVbXTNJOHz0NIUFtYKcDPo3PtAIoZW/JC5VZw9vDbMTjkLKG
R6VfjLU9i9Rtl7vY6CQZCgXln36HSLrtb0uADRyTBjJelnFLHKSz4G3ANvqLZ33BRfmyV2cYls1B
FDLHtuGy1AKIgPuEMqWudSD6ks0o9taMGPkpx4xQ8Wp9BCcC5UahZa3CQ3LSQeiWmIY0sno1REia
UBnABTUKuESn7tatmHdCutwnin9zM79aUs2RFN0c30LuZXAmd+z6gAWLAoFfDUiKvQBE8gqqbO5W
96183CBsncuMaByC+2FZ7HJEzuTtXXFfThOLd4t2rUCi+9hpvRQYR5q4ftLKIzYJqgbK09xW7Dgu
BtUR+8rV7Y7QZ5IYpFxomGwaU9tyTAcZSyDaO2zCStdqUxDGz7LiVDqiFv33aoz37qXrcudyoYJe
2sT1zieBKTbfQfznQefhhOq6ptKVJNxJfLmge21d/g+Vnqle+xZR08eh6z3pHqh09BQD60Ox4lmX
PwlLXdRBt5ZeWWee+dec4j1hRpY6lAvprhZtFhcYudi6rFWA7soP+9bxxuCDHWxTm1OA0MDXH2hz
UKQk5d+E0fxf/GnytQEjvDbmRn1LQ3PmDACaOQH9kfl39ffYiwLa3qk7cbfKvu0Z06xUuTBngc13
cdQT0r1K10zIpHMnvj/mP5nLYzCddMcFmD5xOzGJRgvohF0UPNrqw78RjQ8nkj6WQG1vdDGz+up+
vDzc6I8Pv+Gw8fDQBchMc7v/hQsDCFucg4XrGkc4dfmOly1bEWfn+2yR/i3CwAuGhRndeYQ5Qw5g
B24RQxx6gGtcXXFZXf2uxQAfCzuvM7dovor2XSSwOOPCFJOV+BHOx9lJA+ELJlsoepEWXsQYPiZe
kPMrRFPYNWYWIiT0FwA+EJIE6pYOEI+QEKvXnjHllNjTvOy+qrwy6FmtK/txFU0nfATIIVOtTcKG
loc2MocTQ9RGzRjh25oiYo/MC0kmrN+amzn9op7BonkUO4kdRfwoAkj0lLZbDSqx5CAbeqQBIycX
cSovlBoCJXdBt+/BldpoSe/NgswZzJUPXEkZHucFqs1JLw/uU86xnTGwM5L7StSRnbTj8dp/Exjo
3hh0Zltel4DlGhlBEbcyBeZvHcJ+Pj5E9z6Mk+XutQRItpo8SP9/UkLpw9Okq9Hpj54519Q1fIn3
QD1TTqtERpW9/kaco/V+oHIy6mEX0gzgYixx9ERfJaDFSEgDwD7HkG/mQUnwanfQ/Z7423g5VeOE
ebmwnH66v9UqyVSXFJj29w4e5dOFYA6tkTLMnij5qxVuP2sN03lw7lNL0zCdU7+4+zQ4+mD3rXBs
kklw60Zrc15eJ9nyLarGXSGGdBGXjBgugMHVeexdPuyjcsnJMRwU8pSzwM4U96bPsVRL8tgaJLbD
cQc+zP0zo1plKZFa8d+sFwMfbsJk6opxFnXipe2yLmGeB2wlXD377KFnbJtPgUQ6jIbHVBYO35ta
vrFpinU5gVijSlaDFI2J6QG5GtviTjUt8Tumf9HKlUd3Q0b86zW/j9ycMK66uw4ANe6dkk910s6g
qG0jPH58m/aTIjYHwrXKvNHza6fapy3E+iCDjhSPPO0G2riKM1OGXc9+utV61MKgG1tnBtRH6oyT
gVdwIQ1GombED8Y0/hFLTzYiQJ5iVDEEWkBOasmZ5MTXpFb13oMfJLkIi0FY6abfe+CTjF27Ut4Q
O/DydCr5pwUeSovp444WYYX5TQt4cpb6BlbICtnULRJf5ueGJ3rPOhQl8O5wkygWlvqjkLAC9C3E
OTiYPQ8vOqvTtN7x+2s4TIfQTY7fUdZJ0CnZ7Yc1LEpfcwtfmz5T5YagVs9Dd0xG1uoTuBSfsw4i
8PKzbMrzl/ONhkN6V7i4FXBg3JqYWkHYu2NOeUf255oB2eJAkodZ/U3cb4Dm1402uyT7le6m9KmG
0Nuy6+S1feewRz2CxQK6ufGzMV7geC+W4kiwPWMGxnrfuWXt74jKKERdDB8RWOcCWbr/L5y1/khn
Oy6d86fUDs0e8li2pAIKqYb9o1GizZf+HNXzjITHaDi+FxK/syWxdxOMJJ2VlIPAaMjzsOEhqABL
w5AFukwWxnlUbF7J623HwCr3nyZ8mHzI/LA3HEcQDh7nLSHatkJQ2X/zs97ygMijMgawcoZHtrvp
UcaaoN+yCYsse3lrV+QPQHG8TCnax0E/Cjm6Q3mazyMWGStD4pu5Nw6GzWRmVbPcrWYwyqxwhvqX
7ZfNAe+QE1ZtxIm627MI9znvjwZ6oRHZt3CUmy+I4a6ZCRvcvlFpglVD4U9O1LhOkl8PIojtx6Wi
n/TZKH2tSiDgvm9MyCgxa6hxFjXkSonGOJ6AAcDOwD2rjuDHd89JYY11DQPtMlkC7y5O3E0NuUcV
Ywr19I4CcofP2Z7iP0sXDXU/w8B96dShPyWpYayax2NSpaMoO05Xr1jJIuEZNUaoj7ryhlzIWo1J
LD4N1fNdnBLEAEyNZmO1nfgug9wA6jD6WzxBHuP1XQ9tI3HZ6zB8A9j+V09oT/jZJiJ1SZX7e+p1
7c4k5qr0XXanvDTdX9KzmTuko2bxI4jo4e6/avtHzIPLV97tjfhwC8E09chsGDRenlTfQLTxn8dY
C86OxjHbbDV9NzND8wq6sDqrgCHtiTkwYT9O3791gf3L+camgBBSlcvJHqxn9tH2pQjOOVR7R/kF
zvDdrl523qrrjbcIvL5oGtt2bSm4Ihonk/jIZ1wiXKR1yccJj5ezy/LNAz2u9e0ZceUTlBKl7eBg
RuEX2cDGhUdHPdFKagesjwDdaelxa5GdBfvo1KovaoGftm/wjr6m7RCHoaFAjm5QQckA8TaPODGH
oZ9r9QNaRcx3IsWBjf/L26I9IAWZWnxugUH3M3ZAYCZSgcGarlG2zji41Pr3bzoxbpdbvrMklSoM
dnou8nKWe4aXiF0=
`protect end_protected
