XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��$ެ����Oȥ�
j��<Z����� �_٠�`&�DB�NX��!ۺ)�*P� �U�4d=�ӣ��6�Lo��C끇������YE�3q�IB�V�!���Zˮ��>����6>�jG
�+�3K<��L�O{��Ȥ�;�l,�+a�9i��hZ7C�7����x$��v�{��p��ɛ�������4�tA3�?)�FƅX����zA�/��DRn��l��_�����w��/�'�Q��TYY�ɦk���}��0�@HM��2 ��N����_�:�]���\hV\9��&d>�R�'�:�|��b��Z�x�����La!�d�؃{���SY
���l��6�ꀫ�ٖ(��.r�}tp���g'm �� ,ڝ\�X5����������yJm�'�ۈ -1���,�B�|�"%��V����m�I��4��XVl��j3`��8ͥ��tvz�x���6�ib���(Z�Y
+��#��۹��dy� ���̐$3�;���F����m4����"�)`-=A�,���k���]1bf�3��V���v�%���'m�x��ac��h]rK��8��x$/,�6oA[;��v�a5�	�j$J���e��"\���;������L��K�mu�Gny̱��X�m�u�Aon���5�< �����.�9��W2��ɣ�k�[�.�J�=�[�ﵟ����Ip���B6@�.�;�]|�-pq.�)�z�u<�<O�^�泤�s�t���0v�⯂�}��VXlxVHYEB     400     1e0Җ��:����^gsP�`��|��X4挦��3�KuY����{�?��k4r·�LH�FEk$T'q8 Im<�
�Z���1u	��.i麋I�X~0^�)���/�w'����Y�髎��Jp,B�"�
��Y
&�	�.3i�B<Z��
*4@ ����M�Z��Z��o;l�{di�
U�xei�j�Z�A6��ؒ�9h���G��� #�\%*��i���Z^��[1�^��w��ć�RB���C;���TsHp��M���;�(�~~���r��˹�*�&���J���U���Qd��R�������Ȥ�~@J������0�tX- BH�u5��x�|��5#�1�[�����;�g���k�3Iͤ0Y�xE_�P����)�_��/�����g�i���y\�1��m� ��U{�l/�~�Lp5��;��ڍqrO�X��ϏP>�7)u4'/�B,_�2e�BXlxVHYEB     400     130$�cV��%v�ij�����S.M7�P9����}D�X]�r{� ص<�w��@)���%�F���+@^�|�g��N����l����J"4N|m�S'S
���ޱ �'xF�R�h\�G�'?�����Ys���*f;{8�-�[�2.5��'/���@�%$3��������[YZ��Aѱ,��]�
7jFBx��J�	��J.�?ӱ�X�]���b���6��p%������w*,�;�V�r��J
;�l�u2�ZэRO�-�����F�����	okQt�Fn��Z����tFniw˙�L�XlxVHYEB     400      e08�N	���zgG� T�)eS)�4?����B߇&�4ҹ�A[�n3Aͯ_ru`m���B����E�!��E�6
���9��.x'����8\�[��	�kg���I����>���	*n�*��pL���eN��j?��[��hbC��x���^r�r����;�����2�2����TL�����Y����Թ�vZ��W;�H���d�;�ϸ8��K-���XlxVHYEB     400      e0���e��ɨ4 ��y�ME��@}���}x祥��zM=!stuO���ޅ}{�!���@�����OD�+nHt�qũ����`����;>8nu�
��"�P1 �:��-�b�C�����Z�H���%�|n�R۞Pɲ��G�la1s�a����bێ�+5,� $
mk1�ab�7)�v}�����1����P��+�@@Q���[�ߗ��%�u����o��r�XlxVHYEB     400      d0��t,�4}+~y�B<l�:.8�V�n� 5-3����OG�y�&�%j�����S�H&���`�RY��Z�ܰ�0^������p��6ʤ��Jq��ˌ�;ȓ�����d͊�Pi�a�S
�C(���J�ik%4`:?��c0ScPf�$�>l�I��1��'��ǐc/7�.����壐Q j�W�7�����������lQ�XlxVHYEB     400      e0Q��4���ay�����D+VU�Zg�\�6̕H��xP�?�Ǫ�Ơ쎪�m�H�W�j�!ĸ�:j�J��Q!�U�$�i�묡_L~�VaK3҃�������&�ks���-ǽ�;W�����[#����Mf�~�<�B�e��(Φ�d���$(�?'9b�V5�G���R���Gn��#�h�Ve]$�u�-����U���Q )Y�@�DIkEk+��rXlxVHYEB     400      e0�@Oy)Z����0S�ܕ���R6�T��������t�ܪ覰-�Co(f^�,c�E ���jy�*�c��j(�ğ{����6c�;ptjK�Mo,Tz������F�23ZT�˗E���_gj �/f��;�";N��o Ӑtc�����"�,�I��t� ?�L�37���'�L`�+�H#����9�}��s3�m7%�@�~�ٯ_��Ϟ�1
���Z!�XlxVHYEB     400      e0 jy(O��k@,����(��[sQ�!dl��xY����f5*�U�v�I�D"�<��SP�� �dRㅿ�sG׍��'}�E�,D-�[욞���o�����\�4=�|��So� �b�r�ŷ�=�>�PlX���O�?0j-&<f�g�� �~��PM�t�fe�4ͽoc-�w��_�a}�?q���:����xٚ�9��++V�ա7�)���1Nh���	�,XlxVHYEB     400     1a0���k�����w['��o:�ٴM[hL�K��%��טKo).��{C#�\\"�ơ��4�v�J����e� ������!n�K� �#��{�U��KI�� �A!/_�kR8�)��c��ıU�Z����W�Ȇ�B�,�� ����0w��ׁ�(����Nc3^���w�'��A�9�8��j�-�s2J��(�l���f�NQ�^#!���qH�=�lEB��	�V���v&.A�x�H��e%�`�{��.0�;3O��3��`�,�S.��+ HC*A��3�ّ���ef#6b���mi����.��9�z�J2Y@���	�����T@O$e��I��s��/1�Z��bt�kc�(i�Z������F���]����2�C65�Ȍ��?��p%B8�ޏQM�XlxVHYEB     400     120����Xh�n�1d�^��X�a:l�E*�14ח�9����[��3�Vih��z.�Ȝ�bU:_r�d�kܣ):)���眠"�l���Z������U(Zi�Q�".�94_��M!r�*yv�����ZI�U��
�A�Ǥ�M���ҟʏ��:�<D�����򤏑o
g~�N�ih�)�)n���ȭ�Y��+��D�cj�q�v�k�!�M��$m���
�SI� �d(��Kf�{Nt�|$��O8z��z7��s���1�=��� 2+i��M�eE�2XlxVHYEB     400     170��I!�(���&���q�&��,s�DƸ/5�~�7��Y�\',g2$:����ěI�"65n�o�O���2;
˚G)_�b��mP�˰kR���Q�����y,�e�q��9ޒ�4�U�i�ۊX�\�� \���Xe�%[�쬞z�%�@��g�{���*b�_C�4P��������Wn,��B�9�s��v��W��䟬�6�t,��[~�F�M�<Y���2�Ψ��D.ө��VS�g����"�*lR1��oW*��4�ڶRVp�;U���e�3��]��CDB�Q؛"��7G�� ��q� ����5�6!�T�1'b=�^t�W�[�Y:�qs4(��[�6���d#`��"���XlxVHYEB     400     130R� �������į��W\m��="Tr��\t9_5#Ħ���y�H��G��d��7�"T�@�Q�n�mɩM�ʎ4�\���-i{ �A\7K��
痲�ΖvgL,�<���Y_����R��&1�i�(� +��'�kۿ���O*)�sj)�V�Y����r�?�ݶ���I�d�~���ś	p +_jHt��hsYm�����+\����VU!�]>cN�D��Q�;��8�� ����D�V,L"_F]Io�ip��6���A	�G�p���2`�g�0�}�b��XlxVHYEB     400     150����+��QEM�[�$�<嘝ՀO�VX�V@!�2����� �L����� O@�o��H��y��_���W����y7iNHh���h�y67��y$a)[��)P\�j[&�dCk�Ŧ׎�+n[��c� A 2[
]5��O(fs���d�?� �e>�Gw&|�"���fZ������.�W<,�ֽ��] ��c�({Cf�����sW�-�N��k`w�ܩGS��A�S7��=kD� �(ؿ�F�>�A���ƇH׼�(=�].�Pe}��7��c2��t�Z8�z�4�����A'����q\}�0g�L��D{G0l��������{XlxVHYEB     400     100���C���W2e	%gm�5�h ,��iZ��=�+�ȅ���R�վ�S�q���<�YT��&3/kq��cΗ �Q��Q���� �����U��������^��V�����!��K5�8�Y^8���9i�������6-�Q�m�I�g:���.#������&K���5���0;Y��{kNSM	�i���9�o'�? ݞ�,�4^���9ͼ��~'�n����ۻ�՘�`=���/�XlxVHYEB     400     140�z�6��Y$mbeA��k�=�(�r��a��(�� ����f��CB�1�����1�lU��Um�K��o9�A�{�~��F�	{DEA_x�@�`;x�hʹ�ِ�qh�I?���q)��O�, ҪU1k�ͣ�e�q`n�}l�6E]Z�HH%,�;�Ǵ�nC�ǧ���#��������,-
�'�5���oe�"[��y�Z-�Q*{~{j�Q;U�GÁ\Zu���-f @0�S�1o��؜�[`� ^D�bqxThVM�M�����^�i��=<��I9�N��F��)��h�,���,��R9ن],���)?�mXlxVHYEB     400     160��~�xҀ�)l>[�)����Q_�Ri�3	��.0�4�"��B�(�Xx��(�c�܂ɰ�m;Q�Σ�`�/'�,��}����'�>�jӇ9Η�=��n3���� ��󂧋��B�@����Vw��uHX��lg���j/+�	`�o7�C�U�����]��|e^���Rot�2�I�s��卂v��-��ٟO��~ڨ ���v]f;��7"+�Mt՚1))��G������\�ӓ>�6�R�K3���؝2z�3��������n9]C���]3��:Hڂ5KS=�"�uPH��LX3�	c��ZP��u|ޜPb�{���=����N�1�c2C=l�>�94+�w&XlxVHYEB     400     120l��{3��p*ka��ˉ:Gg�K�t�ޢ7_�c�_�5���L�]رa�*��8��nj���ڮ�fw%mTϥ�t�O��TV ���O8�@���u9Z��_��MN7�CB�px��hQ����i�8lﲦ�,'?s^#g ��J���/]�Y�-�%��eԆ�-����U8�֫'�g[D�f�\u�=�VoNٸ	T�G��ˌ=��0�O� �1��a
����IMr��2M~�v;���0��c���v���ꊦ�qIց�vX�n�U�aż9�¿J �XlxVHYEB     400     140��Ϙ���R&@q7���`�v]݀d�e�,p�~~��٤SC<C{ސ�J.[L�G�?(4l�c1b���j6����k�迹�^A@뜟R�&�:c�}��q�|�5��:6�ZK������Zu�x��zX��k�������-%�nu��㘹��0D�~%��BP�=����bn'��s�q�@��O6Q���;: �L��40��*���W7�6l�*l�E��2����ߞ����+��v�-bm�{Q_��]��L�g��kH�2��k;iw;6wx:/�w��U:�ns�?Ur������~��mXlxVHYEB     400     130�J�jA��L���U�"޼��U�6���?-+�N@�f��֔"We�s�y�Q8���X�g��S�Qg�����7�����5۫�a�b�Id����N!�f_����=��ʍ<F귌�Y����*�>�$	��D��lPڽ��?����G�����r����Y&�J,O������dr?ctڔ&�=���'M>���'.��6�yM�*�1T���e��1r�����i_g�B���oT�r߽f�BB�q��*��p���tی�i4%nz���j��_�0�B� ~1�v��H��XlxVHYEB     400     150q�1������4��n�r0Ѕ�q.85:�w�����.���>E,יbG�L�?������ΐfq%'��_�[��O�ϙ5hH4t��r�\������(���@�݀��f*��Gں�T.z��������q"�V���t�Y@��1����a�
8t�̚x�n����ݍ���n<_B��0�-/sq�"�}P�$������FH�= |��e��R�G2�GG�$-�{a/�~�y}�˄ǔ�k�k�M-vf̷��z KB�����Du:����\�{��^�������!.@��/�3��u���#�����rA��
���b�]%4X�dH��OI�\XlxVHYEB     400     110=6�.��.|��zR"ԊjN;^xWbL�!s8��B�����N�i���Y�q`�˘ݹ{kK�J9S��EItxF"91������B�I(c�6/�F������5���-ω�FP63��Y�!����O���&��oq2{��e��3��JXQi�@T�ϗoK���ّ��(�ݩ�4ps�V��7�����{I#���δmI�	�RH!������*ʡ,;n4�B(̈́�&��b~$�g���P���(��?:j�#�Z����� �(��`�߅�b1-XlxVHYEB     400     140��ѻ����1���V!�Xn̔L��Yfsɿ4���:0z��7� V���f�ˍ��*Er퉦$�35ε�����O�n� ���\q@(dv�:S��W)!�I\X*�/��/���N1Ucu���)����,Hʒ���0���ʂ	��뉢��˪��5W�j`��ܼ�<��>��6V�a��ڛ�m{����0$RN:�M=����E��,N�U��@÷�VJ󚓬/�[*c������-�_�����	�a� �Yp��L�yt�����vH�w��rS0Bn�t*�Up8^���:���:�����EO�}�σgi�XlxVHYEB     400     160�	ũ7zdp�U�סp'*��G�d&��Ţ9�qnh1==k����1O��p R�L�����l���d}�AU�9pkNOߥ%f�� @'�H��s����ʬPﶾ}�b�V.˕��r���*�����Q�R辆�ʶ4"���8�\�f�ۥۍ����_��pvW.��bA�o��zP%3���LY��˂��u(��L��T�=����k~v[�c�0,W_ˑ��ل�䇽��\�ӻ�N���g�*���&_���"�C����}q��p�t�C�}x�ʠ}�Lq`yވ�!9F�r����b�c�
u�y�{/�/�[d��K�m�
A�w�{`{0�4�XlxVHYEB     400     120A���8�7MkfO� ��񬯧���H.�_�U:=;2y��:!{�ZWL��1����B*j�h|�g��6��=�4U�={^V��^�
0xϮ�)��M����aeaF�t�aZ�Ѱ׈/�����>�	�݅Rn�}�8+��%��e�d(���
�`���O�ɬ>��.�U�C�R=�U�����@@*�n����C���p���"��;�8x�̨�SxJ:H����%k�1*[���y�`F�z�-��ڙ���-�qiB�N�6 )n]�ё���gC�ی�XlxVHYEB     400     140��Ϙ���R&@q7���U��`6��Pԋ+�n������@"��Cd�(����2��h"�1K����	vT��͒#6J�0��P��f!��r�ڨi?���[�p��bC�㗈[i�옥x���D�Ħ�M��j�#���:�L�cP���'Rs>ē���R��',^����^��^g#h���9@��r o���/��]�Z ���-U�gѨ�VM���L���{_^������5S����k�N�D�vn�Q��S9�j'�4������M�*�~�p�*���gw��w[K�C�C�����6iuJ���ѦXlxVHYEB     400     130FN|�Y�?V�#��q���WA5�K���U���9�-�$�-��㪨���BT�Ӷ���gVe �fh܊A���r���y�#E��6��Qr�'E����2a�^�2�qf~�CL�{��ّ�0,�����m�V�u��)���^���48{�����U�_m5�l���Y�P����5�W��{�Ny�n��?W�Bx3d?R�]��;�L ��I5�1=L���:�r���x��&�ځ��e�.�]� $%����{�CͪHܘ�P}j��̄p+J��g�Z��$�I�<Z G�XlxVHYEB     400     150�P�Hȕ�x*���ɉ�[p����'gc�
�]����*ż�v��_q�Y�0������Sn�Ϸ��!a0����[�qN����7D��L�8��dD���i�yq��Lc�ӿ{U�$���/ɕG{d0�h�������L��*�4�$9[H��T��$��$�#'\)QO(���x��n��rO-@۬-Ts����5�~vϮCP ��y�y�1:��Q@�v_��3�*�K�.O����?!�w�	�:� �>'��{&��N�Y T���4<��9C�>�GL�9+fI�rY�ݢ�&}�����yI�x3������(9�@K ��@�\D?XlxVHYEB     400     110��zj|t	t�����ͭ`Ʃ�gf��Q;���X�+ATj��<qnW�R�S�30�|��e����5ޯ�&J������	j��'"��9�zTq
PW:ƈu"�gOȼ5�+Kߧ�!/��0:nU�6Љ��
�Fh��/�Y�T�O<ҟą��3��Ps9u.�b ��L�z�v0�惙1\.��F+n"���K�x�bvq�.&�j�@��ZD�&ȶ�5��-K�~���@l�����'e�[A�<BI|`+ Y.HJ��hОK�`�p�XlxVHYEB     400     140� E3&�X�ֻP�R��-9D&��5@v�[�0Q��t���MNR���LP��pQ���u�w�a�82Qv���=Z�q��J>ƿ��Φ���,n� �C�9��-G��*�֘����ah�c9@��UT�5G~W;ot�Cu~~�dV�#��+��(옞<o�7��@��ŷL�kB�x�|aX���U��q�dC.A���G�������m���̡�;m�aP��ڰ���l��&�k6��j"|4�$`�ؼ�^����} ������sӽŐ)�K���uT���z�GJ���
�24M{Ĭ�㹊�ߘ��+XlxVHYEB     400     160��v�)w`�ܼ�<���L�Q�s�YPP�_o��Ҽ8���&�;��4p��A�}wi�P�r�����	�	4�Du&�XCq��s3�[_���Zq���G�fq<'
&�;]��1�Ң��^7�	�v��T���qa/Q�üz˩m����R�rNʲ�cO�L��"�����M�G񏂢d����X
�[đ݂��w��1�i���̫�2R!�R��;Duh^��S�����[l��4%	�Ў�����aƵJ�1{�`>[G#A��V�#}?��Px6��زU9C���C+"=�;92ae*�י͎r�.���G9櫢V���>Vq�a�%d�_��Md�XlxVHYEB     400     120�W���<�%S%Z�[���D�p�H�{g���P0����h��^��]4�V�4��ȡ��2��UDw�2Ⱑ�+�X�������q򽠱oB�qԴ�I��Z�r���,�>�r�d5Ki�-��m���8�I��J�5H�x�v�L2��%iVzGY{�Q�"�%���g
��� vn/���+�����<�����E@M�����I���?�C��!ƽ����QT��ݺ�鹣r��̮��5hs�?�?z���O	���M4��b�<�6�#��15���3��u�G� �XlxVHYEB     400     140��K�$VJ������(�r�����������c�.�߳<��2]�_���D�l���<wc�G�:9i֓�0�s�M�� ��7�<�Au,�	�EA� ~�U�Nrj�W�'d\wDw�Z�͍�_�}�\.>�	>�f�����|�� )�˵�yĴ��dͰĴ�7��880��+t�9�*��3d��pF,}U��H�X���-�v!����S I#�1U�~	}��>�yb
��|7_��DD���b�n�TA~g����'�տ��^������{����$��~��L�J7C@�%���:��D��Mr؉�+�XlxVHYEB     400     130�J�jA��L���U�"MR�u���Ge
:�$����T�қL�IX����6ɷ��A��d�Xf�@�4^�O��jz�.��;���C�4��s�����z��M��'��-_�(ZRiߝ-i1���ni��h+(<��'fC�8�F�����sx'�����+�}�>~i�4U>Y�����I����Ŀ-�?5ŝc�C ��\��<�^L~�V�9�.6՞��}%6��@z�#�sd� �N.4H�SN���p7f���ŵ�]�Y�������zț32��dl�gw=�²"�a���3��/sXlxVHYEB     400     150'Ǒ�V"����"�֏�L����	np>.񥄅t��2&�!doxK}]��� 5U���&\1@;�\�����\V�.e)|��>�v8�����\g۲ ]��/��Aw�dx���'�(?��{uG`r�(~�د�'�p�R����;�\��<��W�k�ּ�n����) -wg�r��E�K����>=7�0��C�.妼��u� U!pat�F�zg/��{�5nZ�8i���:�<
.������ ���P�����WƈPz�U^S�*�{C�j;kde�0@�++�#�!��915��*f
Q���QD��9��F����w� ��V�Ynf�c�XlxVHYEB     400     120�m�rQ��22�[��ѻ�����˙#��͵�b�)�C�v�!�R��z��6�22u�|
x��jr4?��������JM�0�I�-���E�f���	�Jʪ��lo����|��Siʒ)�*n5�"=����L�N�h�!9z��$�,vyH���Y��p�[�;@�n�Z}./-������k*��^�U�l�\�d���UǏ���G��R��D\�J�?�NؖJ�;�t?9��+��C�5������ >�p�s���:���;�N7�3fcW����/�"vo�XlxVHYEB     400     140�X�u]�m�W?q[;X̯��{��͗[�~�L,Ne�&���A�9Zda�͐�Ov�U8jb{����pJ�n���c�]��8�s3"�W��7^�KT1�{�N�A�n���4B'hDb8��R�P4�	h������VS2yO����.�e�&�[�M�e_,�+��E��
���PQ2����)w.F��Nl�k����f7!Ʉx�T�u��%}y�P�Z���h��������:?��J>��* ?>���?Ty�I
�S�X�'��D��H[69�l���a[i,8k�b�!����_!l�;b���s����a,lb��7��b63w��XlxVHYEB     400     160��W���z�9"��z��o�䩚h���SP�?'��������K���UX6�n��Y���֭�2Yp�O5f�efU���Pφrd�d@�Kn14_�ȟ�D�&���]�2���G(�S�t��б.i\��0>�UG�NT�l1���~�<�D��K�ߥ���\v�^J$��6��;�}T�O<�ZC��G�6_�)Ă�y-���$�B[UMT�2`Sl��A<$Z�KqrNLd�s=��@:�]�mz>�J�JC@{b��O*�P�K͐�.T]�ϼӝt�B
�N���ai��M�J
��	����Q�o�
�̒��<�j<6������)C�-�,E��<�!��i6U(�0�XlxVHYEB     400     120P�w8<r��1[��6��� �� �6�U�NLo�׶�Bo�R���$ӳ�`�sV��h��\���j�9C��lc�����r���'h+�$���P���ݞ1+w���k�)��f*��z)2�=8�a�Rv�U���C�!�I�;�u�
�=l+S���ǿ���6^P��t6��͹���"n�@���Ǉ�>c�:I�yC��K�$S��k+|b�չT�_�����6��%�iB�K+�����S;3�#F3_]�����0ַ���ٔ�������3���"�v�j�iO�Z�"{XlxVHYEB     400     140ڻ�l|s�U8���Ȏʙ߭td_>	_�h�ׂL@�͐��4�D�+�(����[�����#nV�ux)��	t+���AƦ����R���1����Kg�]f���eK)'�#��c�1���}����v��'���͚��<R�^�g�j������z��/Q(��,:>�{-��;��0BbD1�;6�45j�ω�lW���o��Ȥ-g{���ʘ�ǎ]�J��[3y u;��;�+W[o����~��$KL��Y�ω��K��N𱝥������qX�;�LI����ڛ��j�%��k���b��'���`�ؑG��XlxVHYEB     400     130��k��C��Q3<�C��o�(\1h��MK��O���p_j*m-QDs�$#�!�L��ڍXJDǔ�{#=�jX�?!�����ȷN߿j��*Rv̕�p������ݵ2��M+�c�ZyQ�>­�4`���v�J�#�O��,깞>'/�a�9]���6�h�x;p�T�Gt#-af��+�`%ڻR���i��d^�h}�t��)r{�?H���	�`s��X@�ܟ�]G:~$夓q!f�����L�U��$�����V�&݆p�=qz�l����>���ˍ>����XlxVHYEB     400     150s�� �H�GTQ�[3�m�&r�;�+��N�oF4� � ��}/���%1�~�cԢ
��!K�;�!AaM������҂���|(�/�B��i�G�Tª�S�XMM�W/[]���X���sX��̌g����F��+/P��3�_�U�=EӈI�X����G��~Јh�52�{x�y��{@#O�CϨH���8rS?��]�{B��	�fN�o� ![��|b3���5��`����C�L��a|����`4��$�<�'n:�����W�^��p��F�ȉl�� b�/��-���:9OUWO��Zq�C��PKP���(h���dG�o��XlxVHYEB     400     120�ˤ�m���\��4���xOTJ�|E���Æ�7��Χl@^�3�S Q_�Ļz��#jVFiBQ͂�W	�Tf�kW���xnՅd=��e�<��!&,�K2SN�}�)g����n�V8N��M^��n�=�0@�MGba��i�]'����YVeg�|�#�LQ�zFR�����{̉Ab|s
:�
]DSx�Nf:!�ϱ�xLU��
�ಖK���@��ҍ�M(͵��;s�8�(�����˿#�o���I�(��Gu�f�±J��	[��lk�2��=�2
�XlxVHYEB     400     140=�bO?Q0r/&Oz؁�^9�$-q��G���!�^2�+7��ݱ�#��$�ЁN�l��[���Exi�*Rz�����[���`@5}�Ea�ׂhzL��=U0T�k�"#\$��?h�1���Fw�o��Y'�r��g��z�
��"����t^��I�N��r�j��]f[%����}4����Ē������ ��d2�J��3�R"ķ��IT�����X�%�<�����zp�,x���)g�%0^���>�-�Н�0'����u�H��08:��ʰ���V��P-2�����m�̢�y�p@����W'�XlxVHYEB     400     150ƽ��/��Mc��Ȁ���S��b#U�\�,���FA@ *���C!�nϊAw���$���t$B����4) ����<���u��`mk�Aʵ
n!�AnSH��>�Y�Qa&�5� >2U�{KW�������GDI#盆S�	���C�m�k>0)��+���c�ꇒPM�*B?gu�=���*�k�`��,�������C�i�Y�+����X���_ş=��R+�sV��O�O�L�Qt*�U9/C,��8�����2��폗՜e�|�ur��N[l�$�]5�{2*��C� ��b�!�I�*�*�j5�M�"�S󫾴>��7�ͫ���D5�Rr@NXlxVHYEB     400     120���^f��˱W��ik�:水j ʰ��(��I��?�_���Vu����Tn�h@���p~^�!RP���.:�su��ERf���O!�r�0����<���u>e,����W"ca���*A�t}D/V�-�n6UdKP�.���Gn p�{� �&h�[�s���j"N@���k�42-�����{Ş��!�/OZ~;��-�)=�)��	s��2�Y~g��HE���N��T�H
����F���n{�1sWl�����Zn�l�KK�F��l���O��Ӽ.#XlxVHYEB     400     140pφ�{o�"���k�i	(�; ˧����ٮ0;�*�@��
F�.IF�	e����@�ZOxo�$�. u���(*cF�^�/�9���q|gf�N���R
�|�R�T��3�*�"�1i�W�S�9M���)��ϬT+�HRZUhz��a�X�՘j���w���aßr�n\��b�2/%<�*����е"i�T�����A�еZ��vãt|�2%�U�'�������q��5b�U�z�h�qX{���u�,�]5��3݅4)��5iH�SL>�N�hwx"�����W�.�p۰~a,1�ߛ	!�#G�8�[��V��+x
N�@XlxVHYEB     400     130i=3؟G[���`՞t7+B!* �܅�x���u[�>5kҬ+%�'���#.|�����n2�`�cw�Ӧ��e*�;c�7�4=΋������~�a�������%�,��\+��ۍ�m>j`�ץ���}�I&��3Z�!�nh���^������r.Nq����Ĕ��Q��h֍���|��(�ˠ���́�~H��?I.�Nl��'�<��}*���k�TYPE��i�?�B�S����*"g�蛽X��F�2�`���0�V5:]г����:৿# ��0���QXlxVHYEB     400     150dm�y�@�gN�]Rl6B�Xъ���P�{iDp�s<]P֧��f�����5��$�e�/���� 8i���mM���d�N����T3�c���9�6O��p$�M��l�6�)���j��s����byͽ*�o�W4S1�o�j��}���A�(���,���`�X�W��/+۵4~�#�[��N9� N�v�åZQ(�z9��[I�fQ�W��Q��W�\�Z��3�0�H*p��όO0IM�%���h-��1��G��ւ[�K�����_���D�-Q]b,��	g��>�k]��L��5b�ʕa��o��ˮB����C3�sV��)XlxVHYEB     400     100̫p�l�&X{u����f�g�S�1d�\��g�̱������C�l)�ڎ���~~�qR8��^ �1��,��1Ͱ���x�D%�0��iWF��W�mL���5�)��z��k�jÕ<� %���ٲ�9��LT�٤H.3���1�C:h��/H�Ǽ&^(h�IH��< ��w����F����"̪��M�Z��ܐ�N�QA�\���O�j�oz�=�vS��a�9Y�=�j�%����k0���^ޝ���XlxVHYEB     400     140�����ju#��ǛD�/�`�2�0�6	�&B7)bU�@��?��k���	�YD�û����I5,zE6���w�VgH�v�Q�T\`�ۖ���ڢ64PƱ�Q�>i��'YUt�����)�Hl�̆:7�/M3�`�H�=�H��h�^2�Mk�a�b������
����EGA&���Ư�@/�"Ť���6z
���Q�AU�b���WgZX,��0�"��鲷�0.q��D�҄%��a��u�'�Jss��`ڐ��������1|�B�5�y����
`�HE��M�d`
��gg�b�������Aώ����]�[w��XlxVHYEB     400     160��ͽ-�tn��&�jӈ���6(��YIo�H8�r���/I)C ����@A��u�5�M0�؁��� ���иYd���H��P�*Mi"��E�kZ�@0R�mv���S�c^+J�>:R��j ���|�&���ZI3�ɋ��e�S�h��Ձ�@`�����=�K|���ah%������t[(��A�#�L���a"c��%��j#D��w���|�2��k]"�3) %.�P��'F�)q�0� �9��'�L��Ĺ�K�/S�q3��+ĩ�5=��Z ՗h��N��?���|2�x�Uk}׋��rt/���A�K����eޏ�I\���^f��e�XlxVHYEB     400     120>w��L|r,Tg�h�}�6�mQ��d!��!�nG?O�'B��B���<�T(*���SwdI(�N�v�4�{��9}[��%6���=��t��m�ꓗ�|\O�,߇������+>����k\���5��,��XZ؀LDX�gT~
L_i?u!$7e���s�F��2U�F:�s��L��jIOV�O"��7y�"��$���{N��f�E�q"k��5�����\x<��Bleo�[���oJ���,��im�B*A,(���*�l��8���L8�O��9����XlxVHYEB     400     130���ڟj�UF��r����<jW�}�JQm�ϯ�sm2t� �B������� ��.�P��	|�����ϫz�[K�@k�X"���e��.����r\��5�zZ��!�F��,���O���C�P 2��Ip~>� ����ԹcM�
"�+��n���}jMЯS��}�wͯ�� /ff��9���!^�,���
!g���@e;uAa�?�b��1� ���=�󾠯ם�u+sP�lJ]Kf����,���8��:�i�ٸ�6�B�>twJS�ͧ��<���p]�,_�5t�zXlxVHYEB     400     140���.h���NI<��}��cg�ϔ�����13v]�*�^yԁP�K{�yU�����V,w�P�aS5����y4Ȑ�K��ED�o���R��?v2uZw�Lssп5�-�0��~�rT����uc�i%��d6XhX��C��ң����g?�����b�5II�������y��x�^U��k<��)��0����#4�F N���SV��G�G�E��IІ�!����c!Su�ED�!�b{�����)�M�8!(v���(j�:�G>⯝�I��V<���Aף@�5�,�u�uE
�t���S�i9�L��+�\XlxVHYEB     400     160Biq�-[Q�ba������q3!��\��ƅ{\��	��&OAoKa3C��zd��2�y���^v�P��<����%��B���P��6�H�_����r$٥����g��K�`���/�ɒ��P�e��uC���*��<�I��aJC��^z�7&�-dKM	�2,��p$�{�!5��ȅ>�?�	NJ>�[����� z�n~hK�+��H+5 �����hDlqQ���zM���
Pz��s�:�
���|���9��9T�T�j�g�z�"�-����8f�%�h`�s���!����i�G�U��x��7��M���������-�!�cYa�Qp�N�XlxVHYEB     400      e0:g�!}�3?PB��1��L�VI,��Z �v�tm��@��!"t/�f�v�et��	���d�*1���o�.9~*�� ̲�����щץ#�L��U!��]�/X��Pi77X�ˏ�[	�L�Z���fg���2�p9��PA�V��Ͷ�uXI�B�Ȅ�Xײ�Y�Fn��t�ۍ����&E/�\�p�v}�*��g)E�FVz~�2u]CM�[�X�9XlxVHYEB     400     160�`@��g���{W�y@0̟���_�UA��6i4��:*ߙ5�=l� x�d%{x����f��8���<��I^:���RX?�-ZeԤ��~�_�ά�w%��*��s=�V��jx�Pc��SW��� O��&w"'�E;T�a0AOI��ȍ� Q�"�b����̲���{"��怬4���v�)��.�+�q習�#� @���Ir��c�!���B�E�h�׭��4'~9-� �8��l���-|����8�wL�{ێ���/d/�W�$�%L?g��F��i8�g���3)+��P�z�Sr�w)�^�ƿ�L��3��<��!.���Nx51��������Q���XlxVHYEB     400     150*�
�c3��uH59�;����vS鈅�2�δ�c�ݺ X�����xBɿe���D�R~r�}��#���^�tGJ�9�_B������c�M��cyp�/bƃ*�k���� A��Bs�M�N�D�]y��铽b�:->K+Q�Mz�Kwhq���H?��H'.�4�{��Â_�;	\N�g�p�� `��1?w�
L\E	S77��v�7K��z�d̖s�R��\�J����.}>t2MV�@��{��w����F�/63�G�������2/�N�B�4Kw�Z��Ie��:�3h����2�@�W���O����פ�]W��@nE�vRP���XlxVHYEB     400     120��	^���%�Y=?�NK
�ER[Y6�-���G;��/�ɴӺ.c/	.�)�6�þbx�">L562�*-3E`x:�� v:���1��zR�I��D^3HG�8�K��j�U�`X3;�̓��S��B*��Ѕ��@,)i��e�z�P �N�hu�C9F�? ��� ;Θ�衯��ᖐ:�����Xٛ+�%��l[~�sw��������Yu+`i�[yeG�(/V�.@�����!2G���>��Z����}jS���ցi�����%�&j`XlxVHYEB     400     1304���(H�bz�2��z8� ��<5���|�AT���;~Y�r	��;7?1�U�� �-�1��~Z %QQ�I�"��)�SE�o�|���ډQh��9���y0H����=4].BZ��K�Hj�lSM��H����t���#(�z�A;̉�O���U2;-Z�~��_�iz��� �.
��d80+�~��#�v���Z��J(a�Ǯ�$�W$�n#����ȧs�-I}��DƤ(��Cɔ/�>d�J�E�jT���>�'� ��ڟ�`��9v�rN���J��r���k\�W��R
jx�����uXlxVHYEB     400     150��"������S���`g����u�	p��S�i����������D ��TF܂hյ�]����9��Ec�ER_F���?ԜX��fw{�?������`�,�̂dx�w-p8��x�z�m+cZ��O�C �$(�J!K���@ڎ�] ��|8=����G�?jV��㟷xʂ҃>U~��1��[F����.��� p�l�"�s�7�롚��$��:5q?�:[h"�&x�)Ҡ��'�&1����W�4�C��l)�׮yV�&��!�u�ѐhU�z4�_�<�_���BM�1ߟ����:Q�%��Dpb(d&�U�u	�`�,����;��[�b��*|XlxVHYEB     400     160����y�d^�1g`���pU�d��� |���B�t��ݒd�{�7�Pj����Mc���J�o@������ɔ��bNE|�ꦞ{P��� i�i�!��;Ç�YF�{�tFW�&��_�"mǫ��vt\r�z���N>��1�N�H#��d��,��\gZ�!���&�h��u���8ɮO!�� .�����l��0� �2j��ȇ��W�HX����!���S��5Qf��9����]zm������Z�m��_\�n2S�9�kU3�A%���[��+O�O�f�W4$���{�!��iũ� F Y����1�ZX$o7�v�0-��HR_9�k����,��oK�غb��V<yvXlxVHYEB     400      f0�	�H���t���eZP6b�V{�6��oi�'�����eu��N[�1��_��_}T�~9��:��U9�%Σ
��Bz�<U���y�G��TO�T�;�OM��%Q��za�M�bM�ʧn�8�#��fBRx*�{>����#��=a�M�Y״��D;0����%�0x� C���BQZKH�p!�� �����_��
i��(уi�{1��5٦�Hxo~��ώ&� PsK��U�ՍF�D�A�XlxVHYEB     400     140]}<������ ���1�)z�q�ŕ~MaoQP59p[5ZL��֘	�'�J�[2�aW#��ݗf�5òi���AmvX�:�X�lѹզ�^_�;�aa�	����Yʻa�"����r�JFL_����+������֨b49�)0�q ��V�A�٭�6j�+6��}7�ݠ.�Q(�d�*�X�e�ϖ;w�;3��cYο?�Ž��c�pO��b��FvKO��<�䮇h�����n�gmr.�Tm�n]5��0 !m�ϧ�Փj$�@�T�1,�O��)8��څ�`j�`.�w*&d�.gy��RB>��D�sXlxVHYEB     400     120
�6UJ��'Wꔓ��1B2�5.��נ"���Y6X(u���W����N@�!���p��(	D�2����<�����PZ�87�J�l���b(�BH��Z3�l�\mx+���S�ΈθH�o�ILղ�2���k����}����/L�Q����?ڼH�����B�	�-���|��/�͕k\rσ�&AR���!��\��n%K�m��rv��8�0��")�:Hn:jO���/�-��^�<��F6fLQy��o:��m/&��[&�����x,IV�vy���XN�8����pJ��XlxVHYEB     400     130ka$�����P�:48����^�~F�T��e��axI�N:ܞ#G���Q\�sG�\D�6��W�wr�-H��B�Yf9Ҕ�
zz������
5�H�a�k�JZ�N�c�4��xT�@�0{)�N�c��4��e��ĻN���`JG��/��7��m�a��\�]�so�l�+ M}R0���������� �|�*���H	@�����:D~g��saL��C����Ktg��ؘ�8
��z r��~�k�%;��S�l!�hH��R��3�>���"��"y*�p_�d�v�Oǀg�����1XlxVHYEB     400     120h<z@�&��}Q�y�����H4"rɅ�o���M�v�\jAp��O��X6!=z�1�}�����.La9���ι��KB�J�%�6}nca+�<�6��aZ���_�Ě�ˏ|Y��rȦ��F���枔�ș�����[��F���y����!�Z�a��J �͓��kֶgD�j�%_p��Q-��zf�j(@<bC����h��#J�T�['�������e���uFq���_\čyU[�}v�9���H�W�[P$�R��|$����i�ƙ���P~�zuB�?�hXlxVHYEB     21b      f0�S�\J}�~�C����Nv�ԋ'D����/���ְ䮵�e_ �Ӓ��NB� ��%�<��0�?\�9�_Ya�_kkc����_II
���pt��y/�5��D��Ur��\�!�B�u@_�J��!�y���&w��1�F�g���c���2IEw��k�ta��`¸	��W�-`�$��"i����_��	�.�i)VOh��e�.C�2D75���մh=sf��p9�/ ��S�ז�