XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������SP����b��[����F�I���mƴ-�=�{���|�n)1_�0GU�z� ��������p�R.���a[>.o7�z�Y��|�
SfDO�u��/�3⁸u��>:��0,� ��"0ތG�A(����K�Y���c�2�}6@>���\���V�����y=r�aC&����u)9�,��T(��㻣�;�_I�h:>�#�N�w�����VM����S)�x(�r��υ%�f�\��+�5�mB�Kȣ ��UJ6��i�]S�"��GH��"o��ObK����>I�,sY��&��]LAl�R�� ��ۃ�=���a�屄����Ç�y��8%��>��k��� r�h-�����}�J�.���qZ�"dټ���������a��� z1�,����fB�R?ڼ��ɏ$�!I��MӠ�\��&}e�ŢS89�g�5s'dJr�I�?�GR��t�6s�z%Ț���� H�T`����לd�אg�6��Ɔy*\��8X����(oժ[K�����;n�kLD��%�>>��TJ�#��5G�;�A�d*�6O.p��,O�g�$�@%.�ʑp����$ҵ���Q1Z^9���+9��R�˭�r�B��"�4�b;2l����]�,CR���:WiMD�e�{k��'	�K���5�'s$n�"�ܭ}>��'c�Z�q�����`� T`h��o-�A�!�̒��'C9�����H��{M���x	V�.��(,�Q��q{��XlxVHYEB     400     1a0�7�|�J\�C�<qeS��5/�9A8�{�W���!��x'��K &\�"�`=0s&5�:�� ��T���v��XU����X��&i�+��K���ݕOi���k��Q�j>WO)���}�*f��)��5�FS8����P��@�2��	ۘސiY|��Wm���0%��8;����3��2[t*5]V����g\a����'�^�}��'q�n��S$ �U���~�h{���rU����f��6/u��ߖi�UĹ�=����*������W��7�;բ�8ޒ�ɖ�'� ;�����|ݧ�Ȧ(1�`o{!` �%���uv��@*��a��dFbU��c&���ܝ�����0�Vٶ�J��? ��LQ��� ���;���PnF�M�pf/A�c	���'�XlxVHYEB     400      f0�%�1>�Segߣf	�-��~����N1��t;���V�t��m�*�,��-�h��&���אxyP�[۪�6k��Ap_�5��[��D{�]~})�������8�`mo��b�̳X��k�z�e�3���~�g�Qq�+��o ��%2߼�Ž�;l��)��ſ�g���mӄ "�X#���ңIUS�7�� �SH�pne����k��Չ(�1d���t\S�i�2?��~XlxVHYEB     400     180%huH�[B��&'��l���`B7Ex��X�@s����|q��g Bbr���#��5����5,��U����p�ؗ�� :jN��O�FŬ��$�C\�+ScZ�J����?���ݣ-ŋ>[�Ān5A1B���y�	�ڒ<��|���g9��}���SK���zؔ"�Ų��p�&;�l`߃1k�0�e�c��I@sc�듓��N�y��	�1�+��ko����Isf�����s��D���)�7?� ��je��m�I�Ŋ�ɩ�Ʋ��~B�Q^R@ƭ�8'G���������C�=��K'L�j�Ǚ�u�YF�K�:F��"N�=24����P1���~�[Z�>1�����mE'��#p�XlxVHYEB     400     230Va,E�
pP���̠��I�A~��D�U/:`)P�6;��n����L�Vm�h[��'C������g�C��e�:�T^���u�z���#��ʊp7j/��{�
s $�~��
%�	銒6��p�����E9�)�2]�0�9�< pOybYߕ��7a�玗,+��iG��,�k�}���3M�P\�Ux�����p���d<�\ۂ�Ƒ�N�M�C�#a�m K<*즞U�F�)@�w�Tog�ZE_5Y�Ƣfq�C�����@͛�\��
 �	��*�[*!�97��Rp�K�yTn���t�� �"��
�4<����F�s���X���!��r�q_�-/ou�����u�$������+���na�Ӳ�8O�+`�[ɫ�Mu�;�Ov�%&Hr����ق�4��������?͖��F��\�^�o*6ڏI�Ւ�������@��R��8�E{�����ٌPBo
��(��t$F��L:��ge�m,��i��Ea&�J&��	lk��|Y�)�'�ްr��D֮ns�(����`�m��}P袉ss,(8,XlxVHYEB     400     1c0���R� y��U�,����3l����X�>paa��h����_��3�-�Z�-��q��۪���x����m=^";>C�,�-�a�%�D8�[o�r�.���y���β�N:�rV�*?�����"�,��	��G+Y�>�'j����� ����s��/�R��'%{.�bw���^��v�߂*�B�(�@"����(��хSVmQC�+<�Pa��a�h��j��c����2� �R��ݶE&�����?:��*n�Q����9[�^9I��]s>�(>�	O���`�>����Sf� �moFŉ�>p�R�$��_��j	���$�1vY��0hb.��P�n!�I�z�
�����L{���d�&4}�����4 ��_iD�3f��t@�0���*^���l����*D�9�l� �+ �`�t���|Z`'�t���FXlxVHYEB     400     1a0�v�7D�>�VP��Hy�È���h�MM,��sY��+�ګ�,�>ʊ�"c���p���a��^�������S!�	�͘��
�$s\g�����O�F�՝:�'ҿ�7��#���w/\6�����ڽM�G��1ZՑA7���O������q�������G|&3�[�iI��L��a33h�w��R����g�v��<9y�ݦ ��.4Q���|�;�L:m��Q��@�m�|�^��c�u6�@��J�`�^�?bTJ'D�>�~Xx�Д� ���#KFJr���߁Ƚ���7r�gC ��~+����Z�mL��o7�V~I�S�m	e��sp+��?W��&!$H.eH.ǋ�8D�͆���5��9��'+�GNֿ��_!�|�yQM�[����8���6��w��g���C�_��1XlxVHYEB     400     1a0 Q�`&�5���x2�./aH�m��)�LUVҹ$
<�-�t0�mP/N���
�w�c!����N�<��ӆb����y�������
W[2O���m�*F\�C�s}0���������C4���4_��=�21h���u���<2��Ej� ����(S�����,[t��[\�J�w
���W��&�!�U��c�?#c��Jm�l�����5���p9��Ԣ ��֩.�,(;(�`�(�֝��GT� ���L2 ��A�W>�_\��K�љяQ9"�W����@.?-5�J�|n2|
�1�!@v�y8ծC!�������Q��������<O��j��Ҟ@4k{�:2�k���O��@,��Φc�~ߦ�7Ls��(�����������iҐ�{vI隻���:��tXlxVHYEB     400     1b0��Y~q0/4�3Uvk��!(�p�[���n���Z��[ma�������m��7�P�st�z�
�^D��"����DI
^�]��i��� MGLO/��8���K>��A��^�%VFBH`6�{6̋���D�`��/�C �Q��p�W�m��k�Α�O���� �������7@���di���Z��Ga���#�+<�ꪪ���wU�0�u��� �m�8J{0��G���IaAԆ��󕟨��cM���Xd�a�=��OI4,�M �4��=����F����Ch�0M7te�#��@Y2�JE�9�Oj�� k`i8��U��� h9����ǝ;�	ց�"��Ɍ>pEa�F�H�%�p=�XF�V�l��C�!6(+�K*�\k�5�*���qud��v�>}|��:�
��Ã��XlxVHYEB     400     1e0�D׫��,2���( Fs���V=Di�t%<㆟A�C��1}~7�`^>w���ܨ�E�|���S�y�k�Y<0,�kmY�GUs��W|�QZ �3X���%]�nfL�z`Y�s��M�`U�'m�tt"�]����m����3uЊO+E�ŷ�@Q1�cf�B�����352�e�|�e��2u]��NE��P7�$|ƈ����0I�3�(��E1���5X:!q[���������u���S��B2(�=7~��<,��ō�*���������G����)�J�9URJ�sjf&� Z[7��58i}j���> �سV! �F*�Mp�|�������@�je�0�ulW6�͈/ |�ڣ�+E�X�`kgs	�1_��S٦^Wt��Q��A7��-�h� �xdc������&�Dh�P��#yEoL<��f}G����G��ڵ9��1B��e]�Mp,겧?�{�ʥ�z콮XlxVHYEB     400     170�g����
�#���ҝj�>\��ԀA9�j�2�ldGP�l&�����*m��/r�IJ�"3���03(�庐�=��=��YE ���Ѷ1T8���`H�d�3�� �U�b��0��3�5�Qi�Cfyan�'�����SYJW?�Ui��o�Ս��g��K�ws	�duD����`K#�a��|`�����܈:?��ge�y�nA��\���M��%lqA;���Ԡ1哘��*EBV��%Fb'LΙ��>R����� OU��x��M����h��v,yg�I���RM*�B.���!<��w�?l��u8����ا���p�[R>�C���e�7F�*K�Ia�!P���ڀD��d����_K�5~lXlxVHYEB     400     140gG� �$s��~w\����+/W��	y�� �����MO�����Ke;��*�A,��:>������s}����V�p�_S��=H!������ˆآ]���6�B�Q'7-��4ع�5�^�?Q�tw������G�LW�۾�zq����7��8ɍw���b*bs�?�e[��]�oR���5ƺ�}���"!�\^�g>̋c
��:�[�'�j�Ĝ��ҊBI��r�:;%��;ٳ��+=��_�烛�b�5��*��ir�t7j��� W�oV|3gq�aN䉧v����\�fq�v���W�[�
}��L�.E^X�XlxVHYEB     400     140)�)�Hf�,�!����U$Gr���M
ㅼ��`�W#���J�� ��|�fh݋�ŷ��ROxJ�Υ/IK�6��ɨѥul��H�A�L.A�UJL�u�	��IS�Z�njh���눭��'u
X����N�z���t�o�Ը[�E-�9�0�<�M=�H���y�I�e� b����]gp|4r�&�e9G��ґl!z�<���;���ɣrt���m�Fs�M��An(��8n�#�
�N��A �::��@h9@[�C}@��
EzB���@���>bAT�B��SuU�j��rW�:Q���ϗ��<��J�ᗫ��XlxVHYEB     400     180�j��ml(:��aY�����ɞwo|�"�����C��c����_��h�����(�e97�mPw��]�����`\�S��8�L'�9.����N�p(I�8ڢ�&��աv&��p�x~�q�Z�
B�x��?hu��}X��{�5���(�z�Y�H��Fͨ�y���5��V�D�)�=� 5m�O�O�H�������e:ߗ�����\���Y�D���{�_�hڙO{I�yD�#����U��H���h���y�}�MӢt��hX1
�5�$z�n��@V�z�Z��>'e��ån.�^�8�0����N��|�u��	�۟L�1E��)�f�p�H��Rܠ�\ -~�S��E�p��.	^��}��W@zXlxVHYEB     400     180]M�H^�ȩ�<y?˲|A�:��z�BG���}@%b0�k��
��*���iF��-��i��jO	���Y��ݭ�x5q���t�����ϋ(���{����"�7-_5�\�;?�����<C�5�����s+!���5	M��]XG &B�
�����:�S������=#�����h\ʝ�N���K��Y���G�5>�8�ﻪ�d"H�5<\���O����?RF��F��^�;�� ��U�8ơbp��P�E�\���9Ys�{y�E�P��W��E�+�:T�'��:6띠��\�`�_�"s�Ý�8��Œ��'���3(3U��{�Nb�-H�	�e����4���JEI w_�,�"�������l��WcXlxVHYEB     400     180��k$"c୅>#�:���uki�j�A�*NYH�c8U�3]�6���~���K�y�4�:��^|\�����儾���+�f-��฾�J��p�6^q)�t�y���x�@� �Žۄ�(��>io�& y��K�5⭊ =�ۙ��6^٥f����W!���Őw#�{r��=ib��ʭ�X�5� ����I2����19J,:��Wؗ����EGcf��ڙ �5�ZՖQg�! �h#����X�|��cZj�di~ϼ�rOn�W���E�6p�.���]��r��(EX�Fl.�e�b]X��x�Wn����4n$ t+J������s_դV[B�!���'cR��ک&�����/Po����ۺ�/��ظ����2`�l�XlxVHYEB     400     1a0�V����z�6X�Ҿ��mp݀%�pV��u�f�����҉��t~	E�yZH��652B��2���;��x�w���ŋ����}����q����K�����}��h�ª)��g��D4���n;��d�y�k�c��.O��Q�y�p���eQ�ja`���a�]�#TcfM{��ݮar
��0>�= ���Xv�7��͘'�2�K[+�ml褳{����<Ц� 7u���/����[�r���{��� N�=`�ef���=�����]3�5%��DP�����Mg1��Ȅ&��`�=��p��J 2Ʋ��4�D�R�b�S�#4Pu�+����q��Tu�V"(ʡP6�̊C��	���wOA6�w�+M�6s<F�Z��0�����{7l���Z���cV��� �F��z#XlxVHYEB     400     1a0upԛ�eӋj�t��E
v��<�[9�a�_6C5a��Ymu|@҂*�ʷo��>��P�|���h��(���9C;�����(e:�9�%�`�F�2>��4��V�@=�"D�Rw�(漛�&ᶩ�-�I�*�8���>u����tɱ����?Y�B���H@�g��[������E�nwz��U�|���jB�ޞrA������ �S!�jA���ww,�A�������f��� �U�1�c��h~YټL��?��|�ԖϕUQ�vƒ籐����Ě<�����Tx<�΀Ÿ��9A}�t|�^*9¨��a�낵���ǌG�̯ҍ��n!0�~t�(vyЮCN7<�n]BP�N�t-�x$�A?߷�<,������D��@�+cj��Iw[,s����:�.7��XlxVHYEB     22d     110iU�I�~݀9��(���dl����a�)آMt�,]�$d_���J���)2%0H�f}#�?ޝ���T�+���Dz�����M3[mO��g����4g��J�Q�Uv�"�O#̓]^�ߞ��~C\�m6�^�ф�p��?�\o7Ϗ���Q��05�2�@(����fYh_�+aõ|�����khu`������W��#����?�Xa�F��6����N�"��o��Fn�	|yi�-5��H���nK0A���.�t������o