`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 928)
`protect data_block
NhAWXW3MCN0fqvUFkOQuWnFrSCnTEMzsbG+72K1PDm218AAO5C8G1+gpXMuYcvxXut6IEGxpr8cH
8IxgxwNiXMmD3OLZC0e6f+9EXLkIfXWTeMTeZBJARs/hNYbCcdgMlmt2A92ekbigN1cIL0dwwJK0
NfhLG3CnjhAaLS5hy/N3ItqtfhP2BjHdn6tNKkME33xm+UjlxQ1+2h8+RHqDYO33LK2iLqQKYqAY
S8b4ty9f7VEU8iU327jc8vmx+AKWTpe211m2+VB10oDBLuJwoT8owiWnyDWqiAK7bi1DqefYiwaG
9j6awM9FGTBeFgQq++bTNRO6//homyokxZSKNEW6+JkpvcomDUuWvQoB8JOw9kNWGJIjud74ALKd
7aIwOwHbOk5xn5aVdIMAI8o1quYen65Rry+1fhRwZgjEbSLQANbh9l0N1AEptkEmVNqqc3C6MApY
v1bY45xv+/p1zehtAwU8e81ft96ogyIQIQ4xNYbVYGf8b+PIHcyqqjFvaWA7vPBwFaoAHJqONujj
BRroaFRzvGRzUvQ0D/XZeJKb+nagzpm57AX/Wcz75oqjQUf1N6mRuyL7Pywo+Any2f4wplahKY7y
XUj0ZLT5Gm0aZkyYpYCe+c3sey1uXtzjdtlBmxVL3Ig01SvBFjkGwvnEjHaUQfY+Fpyt0qcYgbdK
5mVSzejIUU/n5bY+bPbB7KPGclvV/GeoJj8tdQzTEGqYT42XKgBf7vxDHZyobuN1Wh6FFcX1DaWH
n87DA8eVS/OZGaxDCD5Elg7GgupJjasfNkbNerI3deszaH5RH489jQV7ni/jkYa6QunQqyMh/V6S
MOiVWHAFepghoZFT3rTWVsJ15/C9KB28llsLbQf1Q7LCMmEUBjNR24MLIjvxVfseqWKuX2PyS1Z+
/9HdYIZKAHawD1DwDC5iGBdy0p7FWMdghm4DRx7EPDOt5s/1pB95HBJEBkWl7iMb03vcKItY7E61
KzBWBMWS7lMAA6XQcsE7qifSY23xZsPKxgH5sJqhzwyOk8AuF8OR/UeXlbYn8P81MrmmJDPnZgF5
mA9LMcgELMPcE5e+LJKzB2zd1luJJVmeHKhl4PimoOC2qcMF+qftCnBWMWC5j0gfj8diesWpjxWJ
8NWOCbvdC+63E8EoUn8S0slOYA6nlzFsL19SabHlNBh+semz0zRv+NbF9FbH+yzoGPubS2qzYj7z
TUNFagmP62jLrLqYDOM+GA==
`protect end_protected
