`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
ParDk3yuQW0zX6yNkRDNDI6GkoWgCyVaYrW8ju/HU1BEUzSDgtcNX4nEUQk3hJGdPz8Un/pWIWbC
m4ef9LXQO/NYfe72zyz8Hxw/tgNMy4NH2N98/hVwqabcPX6Kio6YEs2SeDq+d7UcHrdcUlell5Ut
r6120pboEazcmrD5juMPNI2yqb5DPvqa+/jXEDMVHr0pkoj94L9CizkkOd59D3Yqrk0YiQvxCg/v
9bN0s8aAoLVfEGhTO7I3piMf4q+AYrfHwPRGfO8WF8XzM4VVGo2MSPFnseWxac7PtuyUjbpQQBaB
vNPdRyf1ko/Yxsh5ppZ41uCy3c2R7/TBgBjs4g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="vL93OXfiQJYNjIIo4a3bxRb4EyrJP8xkxur/RRG3GT4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14032)
`protect data_block
oX6Nud922cmqEDZUCGG/eXoOZIIgpzM89xTK3QSwwVuuYNRk+jYU3jE/lxrlRNm/2yCGkoIM3Hw0
Y6Rnmv/TKmbu6E+p1yw4mzJVJ2yeHLfa0UMDCdc6gE3M6IMo9iIqvZthhEwhlLVQ8wYEajyQvxdO
dvL+BEyfx3ChghcDjI8uXz937vz8Ljgbz74KrYLXBvX0+kcZrMcirAflahy2pefxs2frcIi/v8D8
S9KD+XcxuerfiLd9CxtS/YAxf1V4u4+0C2frjrNlyAu7jw4961K9c+XtpbnbIAhru/li1JJeqQd0
u/SI2GJVAGSou6tBBlPSCzQYqXGo5/5CGgN68FvafP98LVQ8MSWtUJYZzhuFmqhVAOYt1dDuJ0Me
HQpHwUXZoreYvbip5L6JWE1oIYEvcyARG1PyzRwFDpcQWVA8eQzf8DUgVpvfCqHSiPfhukySLVOh
v3vcuAEYT+yZwFOArJ+DGx+wPBP7GWA7qMbYQtgudBGKp+r4euBjhUp2R9Riw0Uq2NysgOuXtcGv
AGUWYk9Ja5cMtOh7QEPqv+/gq0kfhkVAdAHFpuCt6/1u5EqmE0xQgM5ZRUlJz5s5FuFHt/gWsFyk
RhJql+9k5OAbUgcD/EsdAcsHNymvEDPZFNDT0oQ2+bRj8sMvvVSGdAv9kjap+OCSJbTThtKo+nwg
b2I7mw8pnk0zGz3UG0UZu5Ku9dhBzDiTGwifkrzsder6JjEqJvkwHiluqOtqhqpY0nIgt3bwJZhQ
aJWswVSFeFo5QLwoV2gI7bx+E1SggoNYOMGmCTnYTN2swjqPEKqLxExuF4aX/JqwTPSOLKwb3Q6J
tXLmU6mIUZdYhhp28BM+u30fAXu73BcvxYiZdnZiu+OyeMmQTs1c4hiG4y/E7/WXEX/2q1vzDER7
41ytgcBJ9sQ2NW5OtooxVjy2XwkEhjrh9yMqtTA/JFK9lRwiN7s7wnYfg+XAW6vztwxIXJtyZWws
UHEaQZAE1wJi+Ljldh4LTkMuJjY5AYKMwnR7ZmEvf8E9R7nwmtAlWbtnAKs8pWVCtb0DgswVcKvy
lhxTK+R+neRRUKYdOsPluyVFrFFr1FEh70ZrxOvnYCg6NkT7CUM3sjXZgF/64iYtyeIbZ8h1E1zT
UUhndHP01nmJqcFYxcPxj6dknUhtPV5j7sdeaX5m80W2FQpBfcYtdMj/4Y+QeH7wKLT6aUPguOm+
nhGqlwy+FAyRrp9vFDMBd3lLaTn1xAOwnboFiUO/DXuhzXLWiXkV0nkHgvGsoktLIunJ6nWV2DKl
zG3u7I1qyrJBMtu2pu6/J8bSRVeXHDshzdalGZfVROj2PoBYt7zGiTpNUZD+p8EqU9ehXVD1KMla
8oisn+UADHI7tEgLbga5nF6FqmbaEKHmLTQHlOhiNx+qdk/Q11mhBg5W2jvkotexp+JRM+X9SKzY
0yy1tdxSqp6PkhXETuVnS3uhE9NF5aigaHXfkhpu7gtWIfW/9ptOI22Ew5kI25ZWA4uWH+oeksi4
0M+p1HBsO7AS8aREquhYOyZK649nFLGydwan1KBmVcnTFpNx1puBD5QR4WjzSgXWM6aE82FdZ8+f
jJH6airbHfzoD3Ie+vrXHiplihuQ8c5ZWCuAz+YPoUF+hSDMlsu+mV5lPOPSO4hYzttOuQFSFGna
7B4vPs/ZG8SUdMw35tGWG43HtMHC6ZsStcCd1ObPqeSwO1PLra4vB6MQ6SUnxW4WR/OS4S1YZlM6
vrCObnRRLAgG8gpuYb25gNZe6HXLkCXQTpstjGXWjWkjc+gSQpmnaD3RCmk6EvLKNECye6W1aZcC
gfq/1Li0GBWY40wUUu0NB0ItFW9egiSQ9F+u9yqkAm2lABZ0NARa/4pbSYtSBsWt0aGXzE+88Qv1
IzRA/+jTpP6XS8VAOGEwm7+5yb2ptwrAgN0Bt3+WNgeVhrcYwCvSNWaDtiHnH48M5aDbsiukUbuX
qdAdJ9F15qjjU7YdM1xbZvERoiYJa0d24Twu41Rc0dBO29POR/XeNlm2Uwyqf6DYSpDbhbyJ6S+7
4qoCr+WimMaaW545kxaDcvKNClULaKXTkgL9nBQ4MX2t8EkETsp9+OhxiIDEFJsxpOefA6I8mvQP
KvTICFkBpA6C0ARRNpb6GH7dOKWlL5xJkPDIJ6HSsitamd09+BTG1AX3/8C49nhw7T5L+C6ZGUdy
qAtQGhX1YkhRD7/lo985Ap9GcamC+bt1/ihuQVlKvl748qBE1gkPo66X5uZgDSeEAL6MOBgyARVh
cgz5Sy9hoFVVoYCyz4WwTUj0GWqrbIVFzQoyTVAU5kLup6hMGqcDogihWumDsT4uXWXQVJsvb4e6
uoPgOSXlJvzJtzoEX6g7fuDwVbATL1luu+UUpoHLO61bo+ARRC+BNXpQhGqwsOCA+QtQOMGFLtF1
bc8WOW2go8Bq6giyx2pS1/HaV1EsgyHP1KkMZmM/cGs3AOrDvDdJ/E7re+vTXN5U9yUQlB0VAxfc
laYbdI6mtlBkgEQcdJ1DxGODfbzbOrrcOXmVfyGN6Xyf1mStfHagxWgyt1P9Wo3EOC3xniuS6/Nr
VBfhRV25BxbfZ/XQPuX9pLbHkmQQEpMOPWZKOkrZqEPJGMgV4NLx9zT9x0UmG0fJ4GBvpE78F2gq
eF0A5f1i/BFS1a3fBmlISGWUjFKBZzSk8YG/49JsFUDSQqilmmbigYZIlfnvR8s7UQd99+s8rqT9
XxXVwNBu6AuQdOdOJn0SDJA/kEzkgkmyly/0saeTWX6Y6rXiyXgcoVW9okZvpz5tqj/j4ih54X3r
t4pBTci8uXZAFKO0MY3HV8DB37f88XdDsD6p3zPwsOB2BPM04yFQT1xThpcCPnbUWORBIfhcBvSK
xuzg6K5Ux2+pQZd8ioihP7WpSkbmXlik4dw568ByjwL27Ux8o3RPiLWV53vdZAoeW363Ax8lh3yf
xOj9kmMJCMNjN6BIBVIYuOD54YW6/b85XjanMEiNIG2/uycSspd+uw3S4k04EIqKO/rnJN11+tnW
OaPnc+GtMRSjeCCs/1DFYOhDG7ZuZal8Cfj72YWKX9n4v9d4CzKv2ls3l0Ts9pwQdyF1434LUuqQ
4n+eAt4v+NxxMUnMCrRBkX5K4gUYdLLxKYg/7nqMSZlO3MimUVCUXHWeLvEZK7zXMnjxKsQNbjgE
ttabms7k7OxG3gP0QbP0F3P1xkmghx2WW7oBqgmNWa5PO3ia+3mLWNcLa6AzuQODPZNGovG5Nmmr
ggRMh2pu8AzIihzC1cfoKhGAZM8LYgW6ag+IsoRZYK4FCBn690jaVdfO9hEKbLbTbWpSsBZ9R0bj
KnNayZXbYZKTD7kz13dzQAespsxG+Gu4ZWjJKQdetK4FiikU9xdg5rEO2tcL5tzs1r1SysYnqj7E
Bi9Y/anw/wDBgJYZ0ks0y0/hY7gE2E9wBJjw+nkdwx6pBiOmPoGqvo3MqKVfDa/WzPgPSeSU3SZF
GuBPNlFDCoIIVnalzmYSayPDf3ln7KYoevF51Qdl6ywOpnCbP31gDuugH6rxAqKhWvQvBMic+RjK
8aoDhqQSAqKAIEw3ewS52YJr5RsTSHV4cTd2CL8yFbqG5wU2G27VhcEasmWf8bBxRs1rT4cYDkND
4czT8vPHUh17wDmSrm6B+ZBwFVBRfVKPFzaR/o86KtN3yWmybh14ncyppdZTCm9UxJGTiKtBlBtQ
1GFNz2T+hT34P9SvSkrlDMjwRCIIPr7BhO52cRBDqSpb/RXMMomD9cxBs4bdhOpMGmeF0BDgvA6B
JIpluMw9TrhldBJi/nuX7zHg1v82QVTlkm3QDOr3QcIGKpcYfogrK43AvrXtVgiaD4biqg8OcAC1
M2xfYit6svJpTzPfMrg3/L1k63+AGuMWo283HWtL34Pi5mEGfMCVqlJ/wqYycSlskta8kaMA0iE3
jojnPC0rRLZW8ZHEbEtwjCLyFQrtKFu9jYMVZOq7pCLi3F5Vd1421akkmunaWRxqcZThvWzMGrhd
py1fMRitT/ui/OnVsGtbCw8LXBjGsjcGkkbTlcaFuTUIN+NDilNgIR7lhtUnUcOC6SSmpYSj7wuS
jpA39cd02Pg95ChZu62AT+n1YenG5aNkNTbs4sePIPUoGDVj5eXhH0CdcvogRRCyoZq3TtNGfcnt
57LA3055i2fWhvB8pSAEygfIL3PUC2trhuILWAYg/PgfImYWedDC5B7fyIajmfbvCQOnUtlNY+TX
ll7WfBmYPu4R9AtKCat9/kdiv18odJtQU/ytXJuLfEvcQzq3H+nJmljOMTBeBLrt5/8jNVQUOeAj
wnfEcL8ujZbP0FqDhttoe5ZxrNspmH93EQ0RmakeiuLFCk3UM2kZqaKpWvtLT9KOqofz+BiyS57N
jxnsun5WSPEQJLoyCTVya4Xgf45aNR/2FtTdCuRXXp0noCZGmRW9TOLMozpyAvZBHJik2MLghIXH
oE7o73+AmGmVtY868KmyUj6i5jHKoO4jxMprBuZ0B2vGWCn+TI/zHCdtghgpKeuZinPzAxx8HpfE
pNpPYWO+DBfIdIUUuqZXs6jsvT+VBMRfW+i903egNr7f67/nahFLLDbGira0PUaU7HSd/qn39gVi
PdIvPHw8DHdelXwP87aFq8Y9IACWD7a1HpvGPA2mik3RxcWGV5bS2uig56upOp6LGptkkEJiQ8Ez
KbDLYrIvOlOtlSmJ0efnVIt0KcsiWdxjfoYRLFWgNce6JSXh/JVhWcMURbrqMfxyEhR6/icNw+OX
FAmkPHC6GhkVTUPKzjWVGihg57Ulmw3PDRAgVSYUEyefV0/VN3jh+WAHPd/KLuTJcOW3uoir25RR
Jze5KHql1oZ6NvNBAeaNBJ1C/SAgtQZqDkKO1/2dlC91/4GI7GS8D/TlCOYyleaz0sp1XACZBWq2
PKYyNlTapFmkKQjthtj87BiklTX78kWab5jFoD4o7V6k2bWOl7EnmVFO/K/u4QsPt4kn4I+MCoIq
l2tk7+3UI6R8KrcIJlv6oV86eZZOmNgxF//YjrrowbH2X3qWGewTdG6KCokw18jr7d0lZCr0nWet
Pz7H73Zl+k7/SVcxre4MnTE2dkYQpLyfOtex2893XibPthERHnJUGnnAk80ZRLAJ0f0Pm/UTGEZT
oQ5+C+N7ZKrRfUqcNyDpIO6a+/bqw4bqHFCO3MSJbrpPVuJErMPcT8MI8yEP37TVxSkiXAjZI4fY
0R+srZoLGueq/ACoFvr79Hoh0DruF4TxpQlEZ60qtM+SrntTNw+206873NI9xbhU0oxOuTKv150z
Jo1C4eVQV7N/2e31cYN9lka0WzyH9sx3WbQeIPF7MbXS6MeWARru+KLHdbAsS3IRWMczltUwiY32
x8jBWPNFGLyuf951l07nglQ2Lwm6AEBwGEHALfTNMgj+DQz953jndJzr0YooHidO3SPb1EoplWlE
71DZi72xBOpNs6oqEDo2l8SDKYNtymqBdz0VU5kPShorJwXa9n1QhzP3Z1Mg6a1O/o5iyZTS+elm
n9E8KOvZUvg0nuKYGpKQz6pAF9iUYZ5jGsFHvXwJ5N5s4OgfIGxkczN+6D7Jmc8aSehi3Vo5O5Et
kGvCDvRIwvS/Cr3pvQ/r0n1Rq46K9sBjdJz10VemWIHaqDzoZY9+rgcVg/9g5KytwsebE2HDnq5s
wgTy+rs/DSkNvV/N4ev8BwYxV4xFKy5k8wBks8z55hP3M/Fxc58sy5GogAwqCXCe+U4aCZk8xzrV
kH1YAbTLJwlGHUJEsZx1MRddyLupMWEpI+09WD7w0Z8Gwkt4znqTocfW6ZvvHxyvn6UrRJw3th24
w0m+zqiOLu5pCJiDIS4TVZNdn6EYoEoj2V1bye8CzEQPzegOhf0VMyNHgV4dcP7uhORwoVTmyJOU
AjeeYzrTwiILPDo8zmbsU9aO8WsF/lkrOh0/rbv0m6RUWGAaH0t3rR8OnR+2jOW1bAGCNnKD0xpv
GfdxdSuBo7rhWvEdZy86ZwLGRQ5F/nRmBLQawMCJQXlzblYldhn9uG4xXzyNnhMzzqC9r/PuH9LA
4pnr08RxwkwoaTtz6CZc77t4pDDA1Pk5TJAPVwk/YPy82Z9pxZ1IC0YWzcU7oKUCiArdFhxb6uyC
OPAm+KFSHBjzlVm87fdHtmRyDTmybttCbX+m7dzdYpgj/nXZlR20/aRW6TNPts/IeMhQUESIQoNL
TZjjf1Fqf1vtKIxF/iLA6m8/hs2Hr9nPqjURNCui3Vfn4EZVZE+T0+f7uWYHfIBd4yngnPUcWa/+
LjATK+pO0oaStFfLfS59T4y2AvTddyJCdIRMXCNhdeqXU3FFPBD4fxYYPKPLzGBqNCfmu8LyVL+k
2Js1GrIkVI9UhDjaY4GeC7R71gvgh64cwfrmN9D1EhGO9Kz902lgcPbQUeJtN6GHDpMe2daEEZUx
CYaM0emHxc9YzHnkfY1rQCWlY6vju709d8jfW5gdPUstlJpVkqf6FtzWekLoVRDQtshN8qtVvuqe
EVz0gjBfYu0+jJ+GYRvNJGo5ElUQUtbPAfgevYESpp/ymPbnSWaEccILFYlIWSVbZ6QxidrGln/R
flYWRJ/WMO4YeaEaSHpUAlKptODLoLyTqNMAbz+0+y7mwgWKTMEoZwGaHbY6uNPsb46pUh25v8ZN
6HGKV6khrzw+zq74tG5CQS4OwP/V4GsisPooBRodwU6hK03VupM/fIkbFrbINipzXRzvxqMVZXZK
RbvYYqo+4weiRrKRjSSbAGXb2hQyN2RfO8+vaOaHszAtoXQsvPLFLAZ2Qc8DJ8KkPoVseTeGPaNT
dKTNm5Tp83OGqgTn+CKdral4qsplkrIx1lTRrwyRcVlUupjgKthkPl+0ef2S6Ax2ID0k3qhWnFNq
E0YSpRxV9/hy7i1z0Ko7VGglEEXrEpRBJUFH2krZ2e7cJ5ftviD4jMOpGrMqOgv4s6tU7Owk2wG4
Q3VsprfPEjBActM/WkGCcgRp8q4kBEIq667V6+cgWHjp8NMZzWh/vz6Z9Q4fuOKzOp6K4KQPfpjB
kZaBgJRMJ2Jr68Pz0omsshdA49T7Fcsfc9YsKGFRy3hE6o7NokIu+ODv306RdAT6pJppW/SANE7B
safxL2myehCkXBBAFGdFHhASOYe/z4iyDsKZATNB8kfZD4th6l3CMrn+Iw8E/2wXoRuugl6QHmZJ
Mg71hfm6UO8xeQBAShtul9GrD60XBclZbLjDD4zzqbWL8lccPMCYqUTrNSY4jPuRiPkUjpx/iZEB
XlV3rjD9d7WNVMbRO7eMzH+jmktbZZnBz+C7hWu+2fQRFsBcf/FKR8GgYdQtp69zzgSNJd1Oz8Gi
mvV1gZbs/1+GbqrvqDjtaWYW0eqV1K1WAUynNvck5GFZAeqQzvErhNgjsDCFYcllZ1l8VNpIeH0i
RekgF7QX9EvWvNQ0diPZtfHNz80aZwJmqoJxNylM+2HzXbcu29xjGzyPVc+drz/rQDiFFaPkdtTa
53Q6XF6BLkrqCr8lNrf8KLK1VUwGy9Pt3o1IVVle3LkXbuBGjIKmr+4UacZchvYgJpuSTFbz44mR
Wnzo0Z3zwZ0V6tikhIMy9g06vlYBCgwE3Kvc0CvsUrnNzeInJlVpOosRoowrHqBUIPOCMvZ+OAzL
qDktYREAr65oAwZM38fjmfxHHcOyDeHijseb5TkWM+44r+XReh2a69eeHfvCnW9zIVOw+8OsUIV4
c59sq9aieNZgcRkm1G4+6yfmmV9wxZ+29vi91iAI55wz+VXX555bC17eDrZ6yb9k75kBe/RQV08K
KOT9/NgnmcS+rlSj9Tdhcx65WnGy6B3vtrhB/515xYuPSh8dv8BeshxydnANb7vdLlDG1dfHFYjh
iqBkVX5NStU8MMh62eY6o6yu6oCswYMVpCT+lMRlNL1Gl/eAtE2vdLFY8oJA5GRaYIkzaQ3fz/P3
eAXldusBX4OxYvX3rr7rm9cGcbNRRIzZKbIh7yZAj7Fv77Wwe9DzhCE+mBXNuPMjApDy1L2kW7Mv
mThXrPKvC9PB5mh158juTSW0OlJkZ9UnQ5smi0TVkajiN6VTIPTXnyw6xYve69EIjWx3dACAjJuU
kRezx6wNDRjLN10eYN3fL05jJv1s0Vv7NA55OwKSrvkj/ME+u+EngFDuJPPLugoBzsvh1/f56+qX
6a5y/K2a/6JHp9gUumkjAWEpteppjl7CWaZzIX+pvflBHPNTKeMtZNxd8g4qeCyNVaTCL/mS12kH
crslXnXcNtjhZU5xWqv6RwZL3fCeTc8szNa7j5i7DneYs01fewvgYzDvn0iYr+5FgsA2AFFSm7H4
eI3JoNC4OSvZ5vAiPp8GD+wKHggeSmomgiLxXjmuZ9DTCa8jOAu7hiWQVRcUHzrLfWvoUFF44pTL
+bhbgfArEROdcCm0c6WHSwArOm1ReKvVZAkWnXw0H6EcnYNAcNYxVJS3+jERZiE0b5lKB7fmdIXM
um841qMTHy6XDHQ3vmhaHQk+f4eRMIKL/Ryu+HW4iDWYXmUQNKK5A9J/HVg193Y3GqL/8TQ6B1tL
KPBKNHMJfTiUb09bAshcBxZqXSVIHNBI6kcS6Fx7ZqZv52XOdK/XZMVNPJXEN4v6oLXP1A0fswd3
JFhNtPpGl1eM9EojXfzhyAch4mQ75pGlq1c3JdGEUezcjNb11AhjFDUSXD/2BQYn45eEFJapq9nE
3n6ZaMl99ds5RtmxcKIwO0oNVGV0VVjc6O6eBbkeUMYCnEwK3RDGcftE84zpyqVA8XSYSxTrGJS0
ZszzDDiSQxPvHwQ+Lkr6KzsKqhBn6LvgAwo/l8HpizJILnztPz6OMVxP6VHyncmkbYnuPuYu7Mgr
K2KoPbQ7eLGDmpWU0kkLx9GZL8tVaNds24c6xXTfETAaLCQrPcJZuB9T2XTc1rw/LoFw1jzor5qu
F851j1AO5nLIz5nsrUoY3ugG0AiDG781wyJ4+KQTFvzrsD42xzQeGDTK1mR27O4tXfMA5u683Pb1
Stn4xzEPgzaiXsS7xy/wE63KVbCV46jaLXSxlx9/X6hZvWDDKW1Y7DhxGGsotTizcne3jeJykUXj
JQi43p/utlt4BcAZzs8VfOZRXhECNYJ2AAVQUtF0HrtD8hxayZV6OjCNZ6fE50Ea2luTfZHnXXD9
FKu3Vi85nmqb+QTfbHZN1mES5GgeSHwTM2dQtAhMv2KAYdPHmvEdAjLNOSIWjFLgO/NSGNm2p836
mXT44R9vKNUsJRwJei9enIjPFbcFOFiZogHApghLHMHdi6BAQUA25A8+2Nj1rWGHpNHvQXboJU1d
CLkC+j8KsSCJ+Y5/Zk0gyOFBa8E71kxkrr5ywCx04rCC+XET63ePghIijDD9OmGA+JEfjDXMvGcC
ked0oGNUhNujuavdxzB4GLfZjO/yqAdK5Uadfdl4Xqm2ogreqEtPVgzZ90K1/8NNanuIOnJzplXw
EAPMvkOzvwfE6cyUH/vx15sFG+4rdHXZjUmdOK8HI6MNPTlaYAB/T3NeGRcbrTk1ZNcZ/kkLt7iF
/qMYz3NXbn6RkP9IsyFP0mjFPtVlzM1/E65OODlQIGlUIBtRNYKIS4pTF+KhaobbtV4qSEbtCeCN
35nGpGEUjKVCaqPN1rGAL541Ny3tt7fTxD2qGoZCPDoyFXIKJmGHkDBxktMqDBkKhuC/x2C+1yB6
6bd7W2/f04REQNL3Yewt3c1mpwhj1cuFWtBod2zUU97z2l7NjC59JaLcJWzIeGx8PG/Tdv7Z+F/q
ohlANPfaOLLTH7EuRhAn4FfI1Hwp+2lESoisSFsF3nVWsyo5kQEP8quq3fzr9gEf51OzSCdIkBta
z8TqH+vjH1gnNPh7NbyCwXSPxwC8XoDnKYB9jpA2EiJmQYiwMCwKycNxym1jWzApPKsJT5X/xPIY
qL64QFkR5n0T2hujk1KbTQFpSU1QDiku1ebK3u4NdaKLQmdESnkOacUZsVVBoI6XRSDCTr1deM3T
p3NjOIlPpkpy7woNrjsJNAoh+R9GWm7l7U6ZbVdM3x6xrMpszU5TLv6LtuEGKsQd9wrvf7LITnk0
SeEgHCsZdPwfgxzVeyz9/KAY5VK1RqlBOkJ+7mEe+LIMQ5YtV+ztRrEccrmqjbnXbCNgVK5XTkip
2IGIAq/QdLyU/LL2QVJ8LIlnq+cnwFP9qrhJw0VTOgR5VX0Yyb8CqNPbLtu7ZWoJ/wVjeCqkCDf/
UnL7E1w++DYJDxyFfmvnAGph4ez8ftBXI/X+uPWQkQ8zay799sPAHlXns668wKno5ulf6KhKFoxN
vBzxf4+tiLW1EHmc0ujsMi999UhGVkZZRowmUncaxO+Jd5tV7IHxQrP67I/hw73vhojLwcyP52pX
seF2jpRs7kFOqC+sFQbAO5qblmXHo9s3Kyeuts7IqRTx0YoSV2IpHiD03lXgc2cjJAt3dPNYTjMm
thX1rCXDqCrLsBYekOnkZ29D015wdm8m5MxVkGzGEKwzPvBVnoAVdJoqhzzJx2qYBvIOESR9MmHw
JenKYS5Exk4QMITVcdL1vYE2uPyQ0BuGDG7nrrDlW+6MBfu67jjMeM0Jonrzklj8zIqIj0HYh4/L
lu+9H2qjCUA9kCKNei/uCMQk7iOC4KK7zL34++XT/j+s2AR2yr8ZVGgRN/hnK/DX7c5SHbLMjaIR
zrzGoyPAzcfTCOdUpXsusuMUxZIqQbIe87b+oZ5W9LHEcXUgzfrIulA7lEnOQQHU09k1tWo8t4jG
c/ZNheY/JgKdzklNeYbunNSaQ3gStq1C+8X6IV4TB3Nk2Surc6SD4ijtYs32qtOaHyB4mvYO/3yF
KCRVs9p7uejmSOJBxaLOXKrupBpH32/zfr3GZPBLBmHFzML9jwZV6PnkLnu+p4bdM8LE8Bghmu42
y94xRPoteEFJap73o6PBXENxpxPOwKdxs9rspiZwrNalO5KM9R295uWW+8VhruvL6Yq9fzx4ChXw
nysSp/VFajaGZmz9kml3cHheEMCGxoYWNbLTkwsGWnyuTvPJI7epmvRcAEXvb9a83DvxJUsifSeV
P8MVVFYwTnxn3SxQ9Aze36DqggaxiuIhuqe2MyVY7r3OXOAL73Jqkdohe0o/yvGjmIiQb7EKmZm1
jcq1pIqC6dWN85b89qeFDb+943DgZQzxavr47NvOCVvRDA2rSmNL11BISHsLSN1yx68bo1rGsqjL
K2hcydOkwNixIhs4g8O9xc95CSUFaO8OyYUGaSxkgwoLdK7Cz2/2mRBZyWLYs9WOraxd6zkvVaMw
dsCoYDgq9u9WE2y9uwTCwYobQ4HH1yiTBOxYw6QACtNAA5LTam3S0AWPBTeO/D/lMLXYtRuQqF8x
6wcnVfFfiyAHAdEWWQtuKIqi1bPVH7AOMmM+q3iU9sFAQd8arMHxIrqbBkgVlC4W6403VWnw1i1n
9FagdondIk/bTsjhUeqTct7boOSwwYqjtrPJaNoZjwZ7vW1axZm4o44+ZFhWUqvg7wtJbdKUSqdi
O2oVhPY+iaFB4WZLCoqTbbCn4PPVnh4HYUKP2fdlv/c2Z6Utu7bbdo/fsRtvUt22TmGa3Rj5ZTkI
sLXcOh51Ajv57GhdGC8ik/5m1KS519ml8u3CgM1jyBSRmaPDzZtU8gDq2lorTnOoB+XjI68CEDA4
b7Zf0iivDO2wNh12SceWm2TwZevcHhDPPrsk5IfkuYhUtqXqsKmquvYS4XFccVaqSrnwPJg6tawy
ijGGGCtZaXclsOBmhtN9QmeGoCjzER/ClQ8MdcRa+99ld+dsbeYTBOXerw9KkZaH1km+IUYbcMJS
2p3UKj75lKMnVu6rTXELAcyTjE8snINuRuJBcBoAPP5t3BI/94K51sAeDCqBtpBXR7a4FXrrd7vR
+NJbSVr59wX9hlsHXy5kmAuL4seEV5Lkh51CPy1CfJBQHufIm0SlugaKeSwBiNflcMcFVD9hI+m7
UYSnm70nkxg7+Ffw6ppN8jVZSMyzWcP1HZCbAA1qH3Yulzy3y7vIkvQE30jAUK3HfOsl6cjq48JA
9s8NvZq9W8hJPsG4g4E6UnoK6ZNYB99+NJoQv+H5THo6r/Naeojt6ysJ+4KipMeH+inZHDJu0UBA
ictfVuIVMViUkHPVKUTR0Bg/gVQXbiCSbmzxfJY3W5ioxeOwM3CE3aAq+iBJthCqB/tCz64bhsb9
vfOJVfzRmZEPdlzCSx5Tf8DyCb3xGyiz4oST/2duRraneWBvaj0UE00muRmLAkF4O0DNwDqrU0sZ
slieiVIdugkDbukmMUf1pgSlDjKpJPQopoSE6xM40WB5c7TPxhpGEANu/O+d7iCwjrUnVYaOXlQH
kvcYcD7y2pCPxmKj5Khqbbx+vZH9UoGq3gnYc5rLCVFlqBDh19ZWD+Ty0w5XBCYF0m5D0N7qLNTj
YNjkRsFRJpPZvKMeODaobjD8+j8t3tysZ3Uc5jginRcR3ogUdZC0ZVgvMZr92KsZL8K5bQOsAdWH
Kr8aD8oVKu5ryt1D8ypnmzQY1oT52eGe6DqviHgsdAYKl50b7ktyy/u4qb+yo7GfaY2FIGYwAZct
6CJzqq3zJ3wn5VuDTHXJUmKjnZ03V9Ct1Q0ur5bKuVQ0LJQu25A/8gA6y4F/ve+fuFlD0L3Twbed
sXCAtwAaWGI5eJgo+7I55hzEeN0gwg8zomDLUgZSF4v33VKQUxXGGKPEhoERAUnFqCrYIbfN9U2O
ShiBTE2o/UfIPiciObh0mHYmKvG7Uz3MNxPfN4xKL9gi8pilk4xEtbjRLrx/imLqaEiOX67owxj+
OoHgabvWT2vJSmLTPCYamJ/kFRPVbkDQvrl+Eip/LFCYxCM2mCTFW5Ug4d/xTDtCT40t1dKOh3vW
cC3hqR8kVPsJSBc6eh20ZYcy6ZZ1EIFhqU7QqTmV82IWunkHb1+WNquf5QwQPGQDhQAhem6XUSFl
l5KtNADFqs1x+nQSCtBN0XIDr7HStG2Bj/J6JtDICsrke7pG2cU105tvK1Go47zH+LZsjwteYZn+
vyvLVdmW1Q7e2QBEV8NqW/opP0hICEpX38NENAj9aQstO4MjBeOL+OihemuJ9lcnMQx0J+RI8/5e
5mdffRmFnuu4u+KdIcupw2fzI9CqxQ/UNt6GV8mwrv2q3eXzjbjGa5o3Qfdicmd2v8+vfPLqTFjY
qv1+HwXBu2ulvSz06/pu25dSVQEhEZoIFaIIj+DPBHlUDi3pn6SUNVLeEk2q4gCrzT7S+L5759H/
C4FcUu0O//vSYfxEBMY0PBBP5xSCcjfJzz5fswdQVwFc1uShiP2PNcmQQofAdwNuyqUbUtehEKwd
d5AUHUJxQlMsRFprB5Q2MCIczbXLrgqwQMYz2oI4oZ89O0IhcwPgoJTbdyX8JYGfW4FP/OXXv9p4
RcVt/LPvTIR52rcTN1Piv7UyHiHZflxfoBg7uZJf2j//TyeA1BfW3qUVG8VXAj1oxyj5ab5LtyaZ
m6kJ2U7Z69zn0m+jbVqO3et+8DHNMuLG1Xw2wFK5oJXmHukgySR5JDvpjhlOWdKLMF43OZTXlN7c
QSxcbF0DTEzBnrDn8t149gdberZBYxDK9eaImMJ/pcxnEll+MfZ8znZPSNcfmdRsect0PlbgjNM1
vLPLVq9rj2oIQuO0rph0+jdIHY8UAi1TTZEZFDXv1nfVkX5LlVUFbLfK5WdXzUvXjYI8Yb3eiaOH
OKjuNijkNZ+yIyQxul0C9VMLRbzvs7e6O8jt8teWb3l1XcbJFNceQxCFWvFkpX6DbwHvMouT2MRX
O30mAw6VfsL2TCHfW2z8KcgGFfu+7LIx7eiYiJKcN1McEKL+++ujB7mEaGgyN10fv7FPJXxA3B4E
g4SxilGzmmCdY3l/w5kw/xX4pfORRQxLinET7CFxZR4TX8mRovuClrZynUFEu8roYf17USwiW9Ub
ikQi5yZDIkk9JbMh6BzeFoIvTKgHKeRm8Ed2f0OPzSqVhCjYL5UHgKJE+ABHGyY7oECwn3vaaYUz
xAv1ixFw2UL4f0G2gc04AnTCo71ckxOTKryFtY2G1Y/nWIQ2WQP/QtxOS+Lx/xtCNe2WWatUgFhl
m8DY0DS0XEhFfrOeR6e1/7XyIalpjTtrUCCueINLclYTrWq1kgsu0h7FHaPlINZ7Xa/+1g7B5Ukm
2ET/OtV4xAUxVeUfIWhH6Ryo9rDdcEJ33UK9zrxHVr5CFzSvpnXHnN8zEL8cTjkKnuMWppTWyZLJ
i2FkFUSHuJjcq2ygKopP0pyHJDCnP4yuYDt6/VMTGhs5wbnIM39k0Lji17SEPyTsh0Qfr+9dOPok
lGeWo7ccsHu1glAxE1bItIGTNNw1NNznK7NUN8vVlPwGb0UfdL+JOL2ThCkdHa6aUhJpsWP0g0O+
Ruh/H1dIAAkMxNkh4qflimhjPb4fCclzerIE+GDwl9nO3q/x6VtQ3qkYTekFPzSXmyJVW3zwVBQI
iureabYEv9pZB2QZGnZKwKqlo2dwBwDPq8fpqMBWIP0R3xgV/lrNd1Q827hLoJ6B9uY8SLXHYxcQ
PEEe+1+nhh4g9zIK+hxuMWbqlUPkgzEIbbHnv1u1YtS+F1yeMaoYjh+b8Na+EOjCpQDqZfSCO5ei
Xj/lfCQ0/pWOVZpYQwgvsAz6EmhDdao+d9/cMo9CzPSaScro4ROvTOFHMzytQyzKWk08WvvytOVt
pLt6VSbXgsQkxmMvl9qbWXPnavu/5YoRXI/JRb077TYF3j0wTOH9LPbOk8OzmKbuIEUM0gzgHtwi
qK79LJKs8IejsBvHcxnPfdvhjMhcuRmc5lhjRsJWHFgYZdABRPOS8+foERRO2Wu4v3YJfcIqa/Zx
M3cxQBhy0lUwlBoOkeLFK8uTQ6PMxHlhfr16HdeG+R5b43qQUIjCBUTPE0533nwTJ5nwYS6YtEEA
qJ26djiDwrVxBxHG6ZVWZFWtLng8S6JhtshfyC/YKcSb+dqPTU6Ap4AAGW25xWEZSkK22TItky7p
dHhp09eirXlNnYylqsFQtlqoM5T+j7TMbP+phFVUuW46aIbaoMMzkEhiJSHhFdl9udTDmLESIIZQ
jWoNLBfspfGrLf7gBAgneYMR9kCuzxWtM+qxSSjnoEN/QEu5Ubu8vrPDccdB4WHM9pk8vH086Prp
w2OUcZLiGrRHDHtgTi4w1zIlws0KNUzCEDAYNp3JuO2NQQbYC50CucjTbAZRL/qRbarD2F0MAAKR
qf974FQ/wP5+bttVk/XR89aXr5OwjPjuyLB1SpDQybFuonGOk/46ojHY3ujbqgdHnfMeNJUy8k2V
LR/cSXRejGW3IjML1O4fIWyMHTOA2yg+UMGS+O1d9y+JXA3zgw4VrNDtLDAz8urula8brG2xygkR
7wTsWDofIJ+j3uN00l+anY5YOIbVxJ/dQUxrjxbp3CqOR2+Mkf/a1I9YmcG8l9kVc++vjG9uJlEB
Ed8WjU4tFmINorhHUPIBoBYYz2lnVBBr6NT1dJFNme07aeR6wMb6aJnVGd65qKNRdAFLcXYznMcD
uugMzO9eS8eWOTcUOFt7rsmJ2f019lDX7/hhRGiKRq6A+2L1UQAGWNQbPQTnXZallwJCokSqiHxa
kD3qmGgFQVoEmX0lfdndyoS50szVNz84Q7w2w43lDt39ehHZp/F8nckQ0mfOvw1ZQmQmIKVieRZ7
0rZYKPQPkhXz4p8bROC8sgr2BbMILdlzUiSiacOn/L113IoyBzPRG5YK7vpoCsG2IfAfVVZvsLo0
D4fgNmseMyvyJgmQmUSot0npaUjftGiMlRodV1+nQ5h94NMctrApaV5gxURhhrF859N4SYI4fy+o
GRErYuxtdznMc3y8PrJW2V1bKwokBuh+eql27gROTiDeH3BkqsFFUvl5FPayT0c2MJGu6LS1/k/E
GIh/pYlcezDGVXVpOZMlM0kZp8KeSKNXitt8F/oe1kx7cH8+L9TTrDkzYDzeMPclca42M6EQSS/N
CYDb25fiw6c3JS+9BFLUvz6nuDwqqbaNaacyYlaiPn8xqUv1vF2ejled2s5YLzzcL0eyxTK+WZXW
58J5Cqpnf7necwY/YG4k64DCX0DRiNu4KzT8oKtX99BBs2wy8SZJfzQOWlvF9oIUYg/TZZpWDJoA
wvtOJTEnFNxAglwSE8e7TX8BQWNBJ7oq3TlQm9knHgNhCRG7msx8neBQ90rqCg3AcnRVX+YdH0PU
2bu8DX++UzkiZ34/hjo9mIcrGgCObQW+olX6tOeD9GckloqFsNC2UlMA1acbsrwLt7p39/akp0V9
OXn98F1Gjj/4ojONxxI2p7nlEyQdBKcA7Oj6AoYrlxvTG7g98id1KO1MWuJGBKfN7GDOihScXxMY
VMjg9Zfc+iS3w71g97m5gRzgtu1rrxWe38woS5MUjWSFVpWLsiG+rjmNz1vOqKlyNtOz7ACgqPoq
utsVFL3eQRAYkb/apcE58q4pPbZyiM7+g2hL31Wvqa2sS61GTa37u0EWrdMOIdhgoK968Y4P71LU
lUjnSVx/FIpWMEEVEu3aZ5BqvuY14Aw+gZKgb7l3X+W4K+d+UYPhiezK3RDZLP55vXC05c3wpuJi
gqVttSTzGl/txw8s84A/BQfPun6H23Dz19RbKx7fQDNlhWPFqFRd0xmPaFIIbSCrgGiF+vNmSnpa
QB5E0RFV52UG4D/EWto6quISJhDuTO8NxsxwR59wGaOIJR0ZYNfBgUXrwuJ6w1lwYqrnUU52hs2u
QbTB6HsZa1w0BZeFELLMwbWHxv7tF9byrxw3MbBogWbzIefTTkqcyBzAeE6yiXRzn0A2E2WxE+Ey
Bv7FpTcOGJAxOGR5GpPGK09zUl5es6UKmxDd9L9L4YnatR69ilGqSaEbaH19qyNg7qvQASd9H/zZ
Wlp1YR81z/XqgdkCw2QYOK4N8/Zr6bWymE2uCo/YxX2h2ASM5pC0mkfo6+Ov3vSq7oZNOzRIj71Z
ZUU/hIoWh/ywdt9dKDIjQgbXUW9nKmOtQAn5BmjAoqEwzSDbNkxf8u1sv7WWxIhG8TMDBEmECdlU
6SC07eNttJIkoJVDYiUzP/qFmCt6/gNumEFePdo8oYsC2qbYSzYgX5tNukbDO6CU3d8I1Tfx4qA7
i0fS+dbcZ7C6gpAWsWCjoloIzCjLQYoayqRF9JXY1/7vNzIKFV7pKrh2SVSNqOGajezUL3HaoKdR
Ew1le8y+qFkGibgyBKleUw7+SMcNRy7avbrQv/o5qbHWjeTMxrzhAFMOfrypkVYB9q50IsQF3pcV
JJqqljv4QHX4ux1fIQtuXFK/qDPe2Z1HrCfQnm/sFFGgLpLSjbMGAMhlsOmdelpXKjguyHwRp/7U
x/g9cT5tb5/1g+4DuMXGldg0Y6gO6/HfLRbiJRPYSUbRvaKPRRBlTVOfBRzqKqP85jQqnVrtvOiZ
Hz4e+pczuNVqrgy856VEjMvmh7q9tbTVGBTTCS0foIfQvN1g0tY5aVe+iNJX4AbGbYrUjv0+qjqj
n0xW9mvFSibguUSVIiV8UU8dgJV+FD50bzK0neAJXSBug+95JyNIm0VNOu9j3LEndh+gDq4X5n8D
SNh2dP3RK1plkhAjlMeYPFrxhRvNaluHy1pYzAMup4uFMhenwJA3YLqhyuoJB4/hxve47P5Q2UNi
a80AIPyjgNoG/nOj8dA3e8ziCGJqQqdXIIeQiGJVTEwK8vr/FjtJ+iVp1COQkhsq+SlYBq118KAg
sN4HJEFoXRsOSLPSlk7aKCrQtBuU9wJ/EmniBvCfLCGVIE8bUrkFCSSUOGW1IIplhJpEgoiQUS7+
WFJaXEq1xbdiXH94KZiM5XY0dc0bt3i/0V/I2iGhQ03wX65/0udZ2Opa5FBdsekr1/elF0xeL1a2
X5qkvzbwbtQOja9DgjiJP8kcrEl3upElLu3o8i6N0nho0WjJqJ87UISDIGom5wFOIxXX7v0b2ijG
RUeDWxWa4juOTdH2G2fAEnTSOnsQZLTdyEPI/Oa+jZ/2UrG5Z9qLnEemrDanco71BVzgQw7ii0Mp
JWbf/NixQ0sQglhFQFU8twG3xyAFEYmxZL1Cf6I7kyBsWlszQXqa5wRRRBoSJ4ohyJrj79pGMn0M
0HvVkVceSoslskVfHTDLbN0mqnDYjK5pFjFQvNIdS/CSPj2m3YtW1dhcycBMLa8Q5qyV/zjFtaeI
n+i1t5naGHGY04ZP+g9zCIrvxNhnXkf5DDugCAtxDWOGS45bi1OM2bdOYyimfEqyq+EjvaAbnW0G
D/h/aFeBu9fYLPLI42isopfzocF8cGtCd5Rp527cUdtLuhbud1ErelyTbPvZtaustJ5EgKB6pDcw
cTzusjdsGkYT9tBwVEceZIgqIEhC5q908JbGM804YcLkYq8VdQz8QTQxShrrLd3LWDRW0d95OjhU
IN7+wwxB23Gi8569DSZkzTBlxRnxEY8mRb6FEssMluJMSf3gne17W5uaNd40jsXLViLghHvQ6F5U
FFTqdYYqBKTErnDwHWzet/wKz5ixVbrY+/CllbMzR10PBgfDYL6XAL20IIlL70W0uhFqWmHFuhk+
dbNgPoQ33fQLH79uuSXpkhzn+UA4H5DReh336jnA7x1/9OUGcEQFlICtqIY/fPLYiuG3vD6iaR4s
3CtChsi9GSpznQ==
`protect end_protected
