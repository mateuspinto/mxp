��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��Ь��-p�l9qe�p}����y��L�Xݳ�,du~{�/�mt't��UUe
�"WJ�>��.���as��^�o�r�?�>��{�z0�2|K:������@�����q�����ev���@�e����p��d	���v#�~'w)�U[��P7��nF0eҘ8�^���S��z�m���x�/�����tn�Ud��n���jv��Xv:L�҂�p6��iQE�Y�� ܢ-X�����G�^z��Y��|����]�b��E��/���Bc��@�0�Id�@dQ]� �HA����VT�)Y�.�U���H��6�<�j(������6�Fn��,h�jj���hc����t�VK��iH�}f�ݤ^K>D�ia]?������Yt\l�Χ| d�{*�������RSj���b_�اv�э��R'�b��յn� ��n�
[2��"&���Dtb�n5�C�� jҼ��\��!�:.$�)e��nM^i�;4Te>T��fs/�w�8ܓ�(o��PUHz��uP����$����P
9pE�������)�=���S$ɮg@���LC��W�����y��0:4q�(#P����0ۋ�@�嗧�1�],c�>�)¾'�@A�3N���"�N���Ⱥ�unl�������BV5N��$,�k4ܩ�#���a;�S.�Ns�ܺ�þ�L�-0� 9��;��tZ-?a�Ɋt�젊�%\wE��O�6�%�tf'�H���C�mZ�O�R����΃�;J8�|��i��܎�YT��f��j(Iqa�؎�O̟޺����=8�[PLP@��\�kT#aέ�������(�yE�lj�f�9]�ODJ��\0~P g.=wa�����$O�[�1�L�B"h=�z �*��.��x��r�7�ã�s1�����<�$����#� >`Ce���+�3��#��O�ՀW�"\W�1@�:TH��N�������c��)��J�$S<��#8��4H {;��Da2�~@�5��	;��JZ,�弌@m}o��䱾���NG�5�G~]9���CUAs���v!P�������9D��=D	B�c?��K�8-T�A�s�縴=B�S��j3��YA5.��M�3H>�F�8���ځ�%-�=J
|��{�E�8;����˭j ��S;��z�>9����"�o�F� �G����čي����S}�� s�w]��9x3�%���G�䫙G�s"`��ܧx��*�h�x��`:4�HWîc^�ϰ�pY��2,��nE�x�2���`�#(�-��FQ�/�
[��Y���}��T��)�mDQ��S>V�V��<)V]�C':��a�-=ʦ���Ld/@��g���`c�:����kat3�9���n� {y���t�N1A*aF/�PsU�@�Ԅ�b��䏣�K��e�^{p�(6��'��
`�nnET���bRf�r����J��)6+�����yC���"ư<.�Ь��m�1O��-�=Ӷ�X5��0{�3}X��S��mYja�m?L=���v~W�r�Ct���w#!!�^���C�br���n;���+ɼ�rVti��|�GO��>����!�}_�["z��g��C%�x��g���%d�u��5\��є����
�K���C������i�0��+ǯ?��[�d{2�#=��r���\�D{��@��Y�/˸�ht�_V5��c�ؠ�=��%�o�s�\�=�E͏���+����<
X��x�������2R$ P�6��1�8݌L�#�VC���*��i	L�ՙ��w��vRX��鉸X���FF�d�7xf�$�ccz���>�r���>��Vܻ��L$&(���Ԋ��b��N^�39���g��S���SM��
Cn�UӸ>��K���*�z��>�ެm\p.Y��Q�3�C��=�@��l-9���DwzE�_ʺ"h�Pk�4KiMb�z��tre`H���Ϲ��?p@˪W�{��k��K���a.>�U d�Ƴ�hBH@�:�G��s�d��`�˴\�{�1�b[�� ��Cm��U�[� �2�������3YmA�
�vR��r߇�۞�B?�&�WtUg��������~��}I�>}��wp��D� /��VD	ɳkj�0�$��h��i��K���E��n��S<p���=�M�7�ǌW~aT���U��b�~�Q�8�8�_>�X�������Y���O��(Gm
X1��OJQ ��Ǖ�ȭM��Ud~4����W�3쩃]��g�n�����lPsd���9|fȍ:[��v�)gv�����ݎ�^_��V�G�)@8�whբz[�{�9��� ��v��V�"C!��ei{��I])�7%*���+�N�]��|?VN�7\Mǩl��hYa�c	u��T�;BM={ٿ�C�r���n�����|NLG��S�'��]��)�xsDl��Zw�L�'����N?����5��pC��Z��-�̜~��4p��C���~Bİ�@�5�Jt�F쇌���{�/�;���C[�ḧKL۳�R��2 ;7�-�t����g���F��<D�߰F�����ɞC�(�k�G!��X��F�.ky�<벸,�,��)����Lr�H�,����^��uo9W�q��7=�	��#7apk|�����%>�Nu�<]J��c~o\+S�<;�U�.�?O� }ȂJ�1JR�W3n��B�
"E�)B�S�,"޸���N��)}0�H��ΪD��������:�f53#�Ÿ��X����BL��8�Ú���&[�-7�b�b���ʽ���~�������K]	��Ɂe�%Xeԏ�//��o�t\p!sD�l D��^@�{p#'1gF����b�y��Z5{9��tIj�p~��hC�� *��3Kc���]{=_���M���I�� e�5ʎ;�j��d�2iB�Qnecs���(\��Q�;�~"�Q Q���tF��	����@%���ܻ^$��&`x�WrU��C����,w�p�R�E��?�[pr�Lf�iA�wYS��x��E[�&h��`q{m��d=��`��f{��j��t�YU�ܐ"�7?�ݢq�����B��Y͢l�>I�RNJN��r�m���q0�!��=��̯XZ
7x����b9^Y᳑[bX�<t�}�ϟL����|�t��H�,!O&�H~�İ��Uڐ*̛eWh��S�j0�����B�~�	 ��V�M��'<���a�����4����7�Cd1��"�r�l���Y���y^����y�����ы[$�f�*I���cő`w��6b"�0Ty���l��M�痢�fH��B2N�������󴘙��I�@�o#����}�^@�ϽS�
b�;_wz����-��H�|f�(��9.���.^�CfzgbpOS2v;.��e���`aA:���]�KI8h��-seﯲ.
��$zŧ�^��2��=7лׯU�'�|�/��ւ3`P�9b�{F<��A��U$���sϖ�P�x��n��ҡ��v�|��'��ά�r�!��H%e��H�[=q�hӰT�S�1�����r`�a�����T�h�(�EO�_�V��첆�ݭ��8K#ᔾ�y'1�;W|��wz@)+�yt�a���l�+�T��o���5��T!q ��t`�S(��_)��P!L���x�f�[	�]^�H0ebOq�X���w��Ѭ�F��T{P�6�|��Z����JY���Ϳ&�D	�
9�wu:��W����?0��3����s:�nrӗ��D?���_	�����AEB���.?{!�c.�_��w�bn��_Xf�)�,� �"(E�Ǹ��3T���p`�QpkϿ��D �S�+k(^�,��UH,�k�ٷTϡ�u�l3u��?���q����������^�U�
<��y�ɟ�hg{������ ����ѡݗ�І�鏻�C�}#�0�0� 
/ӱ��q�?����Ys{Ӵ�1
�M�+u&��*�Є�Bzes�Ū�����CBt�Ty�F�!��,�Ɣ���r��'A#l3:7v��k��pwjK�πF���b{~V]�5��\�Mj�bܔ�h 	]�-�x_��"2=��Bq�L픅��jI\=���}�4n�g�q͵a��$ �Ԉ\�vEK�P$u"��5c��Ds�K�o@_��m�x-����;�� \��|$��-{���i"?Υ�t�a��V9�����R>�l�`L��73-xI�4L�k���W~�I-�������a�Mt�e/�O���lJ@��.8�i/�_� )�=�T�^-��͕'b�"Fߙ�ᨋl슎��q�M���&���(�%��v�6���B1*h�%A1@�%���DCݨ���;Ф�A�G4���Tӗń)�������;X��9 ������Is�[���p��i�je��$� k=uW+�hq�3d�+D��h�<�4]&�\�N~��Un`�&k�-s�P����G��CL��}ۭO��ZOk.QF	�Ωf%V1�';~���/^%���wP�q�O���#-�+:�+�$���҅��L�"o�
9��r�p GSN��{"'\��eڐ��Ã�3P��i�dy7�����׵�q�ܳ��I��_�)&D&HT�\����>��o}�1��nR_�S�ʚ�����4W�z���V����l:�-�"�'��ٚ�����<Ͼ�u�����C	i�xz9�����~�lRK�/�j*�*=#����9�����"�5��S���堔�_���\��U�",�,�i(w]�%���0!���}�N����Q뤰Lq��І��5z�w�^��Z"u'q��2�t\)�d�W�%!��*�F��e�F�u��t�F�.�\���[Y�㮇�I�,�'�D!0�W�/��3�޿Ԟh�F�q�w���^���໣F�{�X�ż7&�-���[.E�5�k�0濡�<�s
�9[NJ-&Ţ�;Ƣ%��]�=ٌb��R�xI"G<���S����t+\'$xr����,�����)h�R����ү�J�i��)vA�o��ؾS�;(ho��Pw^��܏ (��JԈ�ʨsFC��s��yP�����-�h�oH�A�n<rY�-wq2��2t��::~��k%L ���g.e����v�Zp�A1`��� �U��K�Q��ǂ�o��P.�����geF]�uN�ćVK?�ϸ�e:N�}GFbn��[:G��;��Y�3.�z
	��o�
K�=B��փ�~=X���tt��ŘS#��[�'��?��*L�k�79ı΅VИ�"����C���o �N�p\��7�eZ�?c��Ae�nR��t��޻�����f2��
N��2s��rg����%6�6�|S��zyN(cus�����������{�Q�߉�����^�y����?�eҶgEy�ev|!ˣ���L,�w����E��z�i^�6�±�y�5�j�D��0�A)a"�g5��+%BF׋�:>�V�+�6����:{�hr�^��p�j^�Pl��I��y��N�M��z2!vO���l:�P�&u�o�wT���B�h"����T�T����K���2���B
��
c"Z��s6؅�̿E�6j~��H��7�����7�/> `:��d8��*�����.,�'��k�[�z���N�'hR_6�c�Th���v6�ڃ��5MR�>"�8�9!q�`U��:�`^� E��3-H�2{:�7r��l�o"�8]*|u�6P�q����Z��?�ssc�����.����y��JH+���2bG�r��N��T�
�{�Z�2����b�w�h���#������°gY��B������1�ne)��7�o���ۣ.�z�����9?�.�X
h(��]qZ~k��
�
�P{�@���m�T����x��Q�cI;��$!�y�:S�ԝ:V*B�2��1;v�bF9�h�ay]��y)��۠��Ī�n���	Ƕw���4/� �Xc1�H1m��L���
�^��91��䘝+�;�ܠ7#���Q����i�N�uG}�$����Mcz����=v�Q�]7��cBL�sc実e#�&�@h���@��ep+���kof,�b~��os��<̳�q�n�I�]�i�p���r	*���� ��_ɐ�E�*�c@~=\G��ݻ���D�(/��![[��͐Ų�Bv�!D�K���vH��z=�7�9u�������J�a��=O%�b�p�f�e�e�2��� �J�/DV��.���&�B�v;���z������ 1]� *
����.��d׵���'N��l&��Gh�;��XdXV�ެ����M/��ܔ�a��c�ҵ�q�F*���+�*N6���)�a7�dHΟ�Z����i^|�Km�)�Sk��̰z��^��.vI����1�Ó�i '��b���om�ă��4���>����*{C��5��������C�
��r�1Ǧ�V����w����*��bn� 31�3'Τ�p�x��Z�׀Ҳ�!��&��r%��4�wᠢI/�z����ZZ���B9b��c�ƄJ7�\Ů�b���$�^^����t'���Lb	(�� q�-l������30|O@�#Ʋ�A1U�z��0YS#�)!_^Gg�^S�S�FEB}o�N��i���gK��㼞�!�J>T�0�jsKk��o�^��;�{!���M&�������r�0{Yw�R=��!���O^�o	�d�CT{�F����?itQZ����J		Ccj|5�Q�f�7N��j��c4��2Q��ek�˾��!��_Q�������"w��v��-ˁc>�o|%r�Q���Ȕ�3������h�cc����։�{���x�2�����*��r3�,l����x���ç���q�w��h���ﾛ\�������Th�7VƔ<|��I}��c��B��Ү+F�Id�};������AÕ�f�T����q(f��ң�h�����)�3��yi����!N����,�b$���m��,I �th����b;+L�>�\�;�=����4�"�Ve�L�+�y����k�x��p��PM9+�^S�J�T[}+�c�Eo�.�n���_��<�K
�uV4
�w"-�Dh�,m��f���IYW _�=��M7Ik�Q��$'\�%�B!}+��Է՟0-煚UŒ7c���A4G.|�P:�ު���Qo���O��kjA�p�J��"\��J����O�rd��έ�O�����|���#��\+)�h呣1SH�K޽�^ݵ~k%s��ŘZ �e���e$R������w��8����L/��m~p�^�����"�H��]��7VR��Iv�H퍌�>�i��|���u�8Sv@�텯~V��y��4_���㷞��6���;ٸ'�Ě/��=�p}�i����غ���TRU��{�P4$ނL}uy[2�d�s�o!O��54� �mE���i19}l})�7f�:��렾��Dt��f��q����i7α&b�b ��s��}-�ڸG�Z�m�]��:��
ȍ�}�a@����MkNj^d&	x�R3%��;q��H��^��&����#���@U	�E\Q�<�߶���G��"������M4�QA���:�&�����m?�he�x;���!c�������l���sGЊ� �O�$�M��H�d��Ň�I���Yӆ��e�^�ޓH�4�	�ۚ��/�u�&��y�b�K�q�-�F�2�^� /Aq2�Ϊ� t��ކ<=լ��P�)a�����VNH���Em���~�:TG�ľ5�uzptp�r�V �ת(&A�.�����ȕ�7'��j�Ð���J�{��V}�6A�U4�{��w��ՁB5-.@a�-k���G�)�!Əs*�l�G(I(Mv��Al-{ �p=Z�>��@o�_Z���i� ��=
��Aس�f°�9��-N��һk������o�R�� �7������A���X�Ԑ'���:�[$i.O��a�K��?e�|��k����}'[3�Y�o?����m�4�#U���P����㭾�������5��H�RF�2֧�+3{�+�'݂@�Y�h���Ŭ��� 2α?���<8�H�ک}_8nPre��M~��Z!�n`/�.��A9l�Kj��O*#��rԾ�e����"2]�u���,"�.�7f�&�`�̓I8}����X�W�ߞ�pO��𬬾�;'_k>{ANc����t8Y?IU1����V�(4Ċ�8�r"x��	��L��Z+46i��0�)Qra��>p��bA[d��Y(@�Q�1�\'m�$E�\Z��xE*�d,��_QSs�zԟW*�	�7��f�%��Kb<ݘ����r�8oT��4׈�����������!@z��%Ae�;?��RW���&�.8���~z9oJ����(غ�z���%���Y�ߎ�\�9�+M������{Ƣ���2h��.`s���ѫ2o�pP�U�M�\w���lbi֥~H�%��I�nA����{݂N߂��E{�Vv�?::�����j_D3������ɏc��#���e	W�A����&׼L�mۅʫ�k���E�p<4����O���ۂ,�ߓSky�F����S�
��I�u)�
ͿG��4�WJ�r�O�:�@ȟK���Af�s�Ԟ}���ɺu2���@���S�$[��;��,�GJ%}	�#I��x��4j����]���d�x�����bܺ+���Em�ք��!�-��+��zV�EZ��8�_�U��i$�fE8ݙ�D�c�lY��)��u7�	���^��X�y��Rg�̓�0&�i�x��퓃���֠xėX(�a�F���)ה���8N�O�g�s��y���}���;��qM��G�Z����0�7�e����M`m ���/
�1�Yk�#��\Պ@�T�T�r:_)�W��|(����v���+x��
I��}1�Bؒ�4Ǳ^��҅^����٩\ӄ��ʨ��]�i%��wy�6\��3_��.,��J,�q݊d�x���:��:���W��b-�jl��e!r���	��D�Yqt�q=��ddڝr�o���Gz��"�i�֯"�nh���Y��)�qB�'��4J����l���� ѿ�A�L�2��!"��_xW��<x,�>x(�,Z2�{�?�{��w�����Y5I^�R$[P�&�SC�{���we7�����}��|N��@^�����
��5�'�1�_WλLv�-���ųB��6J#9`���v����e�����e�J��u��|p��-~D,�^#6'/
&�u%��X���r�\�'�뭧�:�kj��?Kp�,�&��Jν��N�K��gCC�T��$����2�'h���[x�䶺u��Mx(�����6��mV]+�H2��+h��f�:lt�v[7�kG'��'lb�Wq/��X����8Q�T=cx���p�$g�H�^��o�aD�6410�[mS"��ɬ|�`f����;�R>�ڭ;�y�R�2��톿�_�.�mh�L���	U�wb�u}���2f(T�b�f;�[��C��~��/����O�WO� J|`�0,�4��E��8����	ɬ+`$G�;�l��A�nJ�焍�k���a���~�c�e'�'C�x����xHi�Ǧ�'C��O�����8���v�e+�P8��%�6W��C�-�W\��Q�Z͏S06�"�EP��H��'H����~��L��y5��O5A����q����=����u���WKz�=R�����-^���Q�:H����v�2�{� �,J%�roy
�U/�8)�Ԧ�c�N����O�\��S)��k�KU:s�'E��KS���tV'���J
�˓�A��2��_��^}��g^Ĭ�ք�YR�6r��	��j���>v<�Ḱ|9�_)  <,� ���*~j�~-j����D��ԉl�L+Nr�Փ����9��&���I8���f���1�R��u�͛Tex�V����e���ni�ώ�*������s��ʠ>�㧻��Svk�����r��T��os��u5�9�?�.Wd��K��{�24/�#��$�t��Wk����觅���ꁸ5[����nƕ,mo6A�`F�h�7�4�)Qai��gB\�g�6jb��(^jh���y  t��j"�>��ur���G� G"��ʣ���%^���9y���<(��HYZ��^��]���:�D6b��kj!an��� �����3�n+��}�S]Bn/0���]���J�zV
H��6�Մ}��J�yPg��$�Io3�g�:��w�P����9j;�!y���nCգ�����L����M�cp�`)C-�@��Y��u��q �g�W���f�@���KfN,xz%��%�k�I�`S��-T%x���dW*��eO��hA��,�OEz�-�Ɉ����3�`����R�$+|��PTp)��-� ^v���݃�1(���~���^nn=���D�QU�w�.�N�lR�k_a�7�� G<[��rԗ��?i��˚p��}Ϧ��zш���z�����j���*��߼�I�����IAT�t�<�34R��$a8g���K���v�}�%��Q@xӤ
*��=�G��B�%�N�⃁�l$�T߭����Je�(1�6���N%ޏ��6���}f4^p!h�؈�\��|ˎ�[X��B�����n��(���6,_�W��=�����H�.�b6W�s�*���Zַ�?64���(:�`��s��ֶZ�a�+�r��ɶ�v�Wa�K��R��n'�[L@��еl���l�Ϲ�!�f�����-gew|�B�OL엙eK��h~���R���.=Ȝ]�v!�!��ݢ����E�K�5�{�+��Oj���jc�>��x�35��~�t%�T�2�l�-�}��|��B�w9��[�QXDi�Y�B(�Y�6��ՠvb��%C׏���6��ܢe�K�rd'̀�]*GiQC	���\4�"�4�'/ ��ٖ�܀���7k���$N$7[��ğ�bA�=�j�_�&%�麖|�4�j��C�08w.�`^ZZm>9��tn�Hxb���7�ޱ�l^���;�8(���B*%N�֐K�~�6a#��5(�n��Q!�%���.�8�?�R6���\%&P�m��z�a���VC�3v�������n#~zK$}�Q'�0pP���&�@O�I߽E�6�0�i�9�g���k�������X�M2�\��'z�WkW�v�3+g�t2rW�5U|�V9>����_S��}}[�.�n�[�+n�9\���4^my0MR>��2��'�Q�Zi�!3z������"��c��,����t4�-��bӢ�&Ӡ��},l��.�f�=��d��c�8��J�� �C�A���� �1?:�/_���fF�{�'o�*�·�J��(/�{a4W��)�IÏ�S�v�ri2ㆠ�!"�6|��b�����+:�d�/�pFZ�7���N�8�Z/��{˻8�yz�_>Z�B_b����om�.��z��m�BG��1�-�c�:�H�Ya�����=KO�o�����Q+fG��T�;@�<0�/^@Z�^�Ιf?��hۄ��5N�B.��W��v3��/h쵏O�u���s��!6;��_�L�9��6�%Jx~1;������e��9�o���$��:|5�$.x����G	�����N��ɞU{��VB�����:trű�DJ��NrEw��!LO&��U@=y2D����@@_�\���|�48��2�ڡ��O\x=~�s�6���`�����iD ���0�-��-I�e��hST� h����,�g\���-��12*�IHGt���H�{�gibh��8��z^���Q�3�[�x]Q�� �r5�����惀x�8Z������b�V���
v�>B�=)��;��α0��6&;�l��95Q���>��tL��\T�J��E\�1<�7�0�2K]7$Զ�M�P(���m��jS�N��d0&�k�m?ת�7(��F���~ڗz��<�ae��.G�p��s0�=:�ip9����~�#����'1K�%�OZ��VA�'_�Pf���hF\*
���$�!��*K+�:�D+C����^���u����r��r������j��H@�W:��ק�2��;[�}ORi���h�U0<k4��O���'a��%�A+2�Oq�L�������P�qO��9IoA�a��TJ��ߟ�{_���0k�A�+7X�5�V|:Z�P�Kħ��<�A��-�#��US�]��l��Rb�~ K�b��b�\��:&/��?��3?V>�=�t�Gf��m_,�
Z����m�mb�~ikS������O�`��(*���+�sy��G�ff1��~�p��nM�����'3�fz9G�L@G>�M�e� ��&�c$?�9z�?�%OWn;�V	�i����,''�f��Yŕ|R|}�n���7���@|t�J�A��ɞXܠn@�JEw��PZ0�|]�צ�J�d�2C\)��L����V��Aχ��Q$rQ�o�œ��];�<��6Pkx�� a�!}oV�������z%C�/�4��/��� .���i{9�0��MW��R��iB�-7�=�U �l�m�8�O�t��Z^m�Q�"��Ȥ�Y��"�"�}�5�SN�v�zͩ�|17��(l���\��2'����!�T���Pp!�tY���勯������S��7�%�\���1��{�_҄�454n �ɍf:�[QH����/����=UV}��E�K ���6�}Þ�X� ߪ�ԃv�Ñ�sf�+�� �=T{���-�|x�=xtdO�sW�5g�����6�����
P�7�U�G|ƺ�����d��������Y�;�	�X��[��O]����$*�:~�=������p"dg�Q��3ZL>���l^�P3$\k���N�C�mr��&�;B/�z��:��1ao��\�a��i?�A����=ʉZ5}p��6FlQ� S��<T�hn�I�	'Y��u;?��5����!WM1�HN��������;4U���>!�szыy����	U>�؏ڛ��U�Q�v���o�C�@�H=��C�x���Cӛa�$n�����_���R�����Cp��aC��0���v�R9�a��<�	�yȮu�۰eb#"+�MGv�4:A�^tكlx|�"6���^��$�:����3���4V},�'R���[�/���1L��D�e/�8pp>���:���|F_t�jMo��*X���l)�}�ʍO�uW#$�r�g��CQ�*�20~?;�����t��?�Q�v���0��ү���/	+ȡ�_�i�g����g� o�fMWO�r�%����H^Vb��]���]�
ۚ75y	����8X�z��	E_�^?��3U���W4`\���H)��u[����M���+�̫Y��v��(x�9�I��8��"�Ys����"�p�[��l`,eN�Q������v	�u(YC���pUO�^���D�����B޸)r��~�E��+�1�I�%A�0���v[?�(��W����y®b��DgAZ����E5*]*��*Vr(����O��*k,sޝ���h=	�S%xŨ�^N�桑��g�-j*G�?����Q�DsP��#����`s+,eB�a�V�(�����A~��纟���4XW�A!(֨��D�2����%���z��f:&�ó;�
w��t�|-$�6c&����|Q�yڜ��#ߘ-��aqY0U �v���w:�o@;���m�փz��ֿ)���k�ih�@d0V���&M��9�
]@)�+cI^�,/�G�����y�p�������P��(��(M��ʇ_�5����K�=�雠�vd,-�SCj�ir��G�u�b�s����]sQ��� ub�3-M�(����\R��p�c�ZM {��"�6s>Ϗ�_�A?�7����y0�vl�ȥ��d�? �e��A��
<�~����#���1��g$�=�s�ߠ�u}W�2n7R��j"��c�;��3U�M�	�k��
�@�4A�o
�<&}���d�T��N��$�r�&��l����L�9e�(�I+[`u	G\�<������yUK�}*�H:X7Fbn��m�#>��Y�)!�v�s/̰�_ah�\�&5{���&zC��!l=�a�a��m`�G�x}[Kp�c����i?h#��%Ү��)j �U=�ט��Ů V�T�_<�0����\�����͙�xg
��Zi(��<��F���&|��C\��j�'�> �[�\�~cI8�c	vi��l1 �N^���b3:]]�l���b�m\׿�no�2�4��j���R�9�o�'y�����K�0�2�Z'ω�/��L�i�m���Q����ӎ�#J���^�AOٓiW�uC^6i���2�!@���4���R�1n&�bGm`�f>5�:�3��9�k�\�DX���:��D���Rʉ�>�&�s�B^s��,k���/�_���s�g
�䤕��q�ZU����m��Ӱ�-���Z~O�e�]¡�w�W��Y�@aƱ�[��t�ۊ�8r�˜ۑ�^����C��ѷJ�E�����/�	7 2?Cn��_��R���)L�Sԁ����˛	����wN��E�����x�3�'�ȍQ��h39`�7�)rkDCVcp3+�t�H����S�*P���$�w�hK��]g�Y
\-��SxO�(ŗ���<��O ����_�]|if̇
 rF"��C^���/���(4)�p&>��������`���:����+`�<*y�'}[���,�����f͏YV�g�*�6��S��vͣ�;�C��WcҀS<�/�[�(i��%���r#iM1w���m��[�iJ흖"'���d���t8�If��<m�y���$*��w�=�;J�y�"��t���:�exW����x�Ǧ���W/��Z<�h��gу�lzAx?�n���M�/C�Oz̴��)	b��Q��g�*�pm�R�b�"��R��H�Z5ec&}�1R�Ȣ��������IXƘأL�TJm�a4.�����Y�����7&bSu�Բ���f�֛�<p�a��N��\;�(K]&o�#�j��ʅ���?��k�(��}���PAQ�p��O�^�r�O�5~��U��Z����RM#�%��9�H���b����?�(�����+A�D	�ɷ��ӿ����*|���E@�*�,�k�i��e��ox򏉽�H�PN��k�Ůh](0�T��
?63)��kDc����)��q/�k3��~�voF#t{�-D&����_,��n� �-���i�(�s'Y���/�ik�;�1X��x�I�vZ�U��`�SV�G`xn� 6G�Տ�&8l?���m��|:�8u����K��9O�|��t3��3���5K��|*�be�K��_O/�O����y�~��rBLL�w����YU�ݓ�o0����12vO�+HDh����OW�&A�t6������B��Y/ӛ�Z�X.ە��m�M�4�W�t¶g[��������ؘ�r2�] �VLO�_��lغ=q� ��͸��GW��!�W�侇�ȶɳ�=L���Uq;�}�KUixzߨ��AKD9��9����9��t��o$!��%X�P�U����tHf.��ka�5������u0���!B�3�0������W�l�� ��_��N:�o�� �l/#J�6U|uhƐ,t2U�'����Tk@G���������߅g�� �C;:��;H˾�?/�HƔ�U�n.���l�Ng�ov�z9�����nOx��Ր���>�� �n[���l���؉�+�b��H�b�32+Y9�2۴\�AE�h �5����kXd�?|��d�����<�p�zN��>�`?:�/x����n�e��E�A�t�RQm<O�\���V���g��m='���:�wqF������<e5��X�D��/�`dI�_�*3a��Xو��G00Ym��\O?���Q��&�g�o]EF�z��[��]N���^�.��U���^!����N���d1��ya�ࠜ�P}�6&�:E�}���Q�Mw���G_~�0T��*m���e������ �;�3^1��;��	�E3�ɾ��*M�[dJ�ԟ�p�q`���˨Ն��Vg�:#OH=���G]aYTp��7���E -^?�W1�����>S�aR�!Ip :cF�P��m!�K�0�s�O����]���oGh[�}f�BV�t�m����ٓò�l�qU�2V�Gڠ�힚�n�<�-�:�o�Z2⪌�g��E,�랒lZ�����a��&�J)$A%Gx� ~���_�d=�B�xmb���8��_�o%C��e�����9(�]]|�{Za6���=�� ��X�vʑG�ˠ�P�D-��f7ԃ�,�M���~¾c�+�����?�m��f<30뙖�s����U��e�*�Z��uc=���e��	��@�gP�K�7�؞�=̐�
��^���H��l_�,i����;.�Ԉ{���u��	3j1�r0��A��ڇ绕]�yhP�y�?�P�ZGn.!mO���B�O�D�eD*�/�40o����ںO�b�E��L���4��xd� �K��^X�;�e��@/���i8�i���Z�����ےv1����	W�eM��ع��}ư(��ͬ�(��&��}=��iR p���9!�T^3�e�_��y�Op�Kr�������5,�(�L�����d���}�a���͸��\��-����w�� k�<DpȮ�o�8�k��L�v���!��Q�)��X����O�:L=�-
�m�g��|�АY_�Q�F�Q��|��q!�?\�4m�ݪ���x�f�e��g>�"����� `����Ii�W�Al�S�!����Y��5W�Z�����Y�ǂ�!3kuf�c�@񩇓��G�F��|jo�5���4T���Ki��I��j���ǩ?����� ��7�,���`�C�;5�8x����"c��Ա�mJΠ��Yi��*Ơ�h5���ŭ�� ���a/}�W�&!`ך9@�:���6Y��w1�H9cV�ݧ��s�3�����
�^���`0���U����R!K��mğ�\�:����&�$v�a?W�ށ�m=��TY1˺+�x��*ZC�d�4v���uH�6��G�D���E�SwL�aO�FN��Y8�� -=���H�� ��=���z6�� ?*��?-T?��� �%���r�QSe�-�ЦtRV�����O��ۤuo�K�AE �R%��p�
�c�7e���IP�1�V�GW���[��n�.0rr�Rj�6_��¹<L�<����d)�*��W�����o�v�y������47B
�~1��r��K4���,�O��ߚ��d�9Gw�*���=S
<]�3=�EF2���ޱ��;�p�[�C��i���3�fv��rM�B
�`��@I4����Aܯe��ݟ/����`�9ma�>Fy��	|T"ɨ���3NR�6���n��:�#���2PK9�]���mۡ_4��E������^FM(���2%+�{=8�!��;���ӟ�n�0 uzB������f���j�%�f3Jـ�Q	#���k��׵�_{p2̅��w9U�.��E\�P�ܵ�%�R3h���ƨE6�K9�e>��ǎ�j����D��Nf�R�pf��_��i� �2���l���;07���_xA�yDT.��Sh����)��6<���]N��kc.���`��c�vAS�o�b�
yGS3�C:P�J ���p�H��� �Ȥs�	R�t���}Ō��O�������:dJРح0@�[�y����
JoSpHSBB!�UΤ��>n�`�2����ǲ`�� ���Jk!�t