`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74256)
`protect data_block
0USWSUGxovGsyBJteYpEobS8pRuGVCL1d83umn7m+GWqBnT5HWRufLhoHlhvzp+qhM5wdyeG9Iv2
nhpuhHdf8JeKAjbYhi+qNZGPwCpi9ymAGN0YMO5K5413Dd+qXmz+2AGThw3ytTA1WB/0Pq6gqaYW
gi60mI3sxkOT77e0KEC4yM3GhDMyb4KQwfk7Rhh/lNDwG7z53IdngNPfz0whtEwCYYmfo8Ida1WL
UwBR+jQE3PDask6wMMBDZnpCgBDN1Rjd2pUbnmpCbOqbje4sdZMnjva4HH1dXzSGWUblGQ1aMFn9
WK1ctE7wVcYIPh6urvBh2IFjwNpd7HABYAib/G1peLoXjWt0pIuUi7TPr/MXGcvQtESDkXr+MQ8H
vG0by6M7/scS1gdwp6pd0PlfsUkfSZBHL7YzEjkL+PSpEMbrSLW2hCnleSKeHcyqo2laUT+/JnV8
xhofoxV9VIMAjx9rty/qMO06SYYe8gDBLpHwoAAJamoSEYY2x24VmIxIsJFyt0TEhcAlALUrxJWK
mBlleR1PI7R6LGdvyEqiFLcknJwTJZ32eepEKh6wiGeYLa2KQ+doEka4rM18J8MCBuHkH9tXX8Lt
w75oE4N9yLeNdROLBRwGZJpTWGhOMGczPfXQ3/1ioshGsRpzOWxt7SOssJkEL9Evd8vlXjM+dgVr
Ax/Zex6I2SzneG3HyM5DGfkY8YaQy6qhuG0o+bmf4OzZeMEd3muzUeTDsgW603zfvJ9ebmfM4QEt
sNEefVXrzIctesvVdcTSnLfxWazhVOOlPPtw3S/D0snxnfcrKF6NTacsVaQa59Njd3Jk0eEd+MCy
oqIB6s0X3HXRU1azErF2/UdOH43x5c8SjN9MSWS8dg/fMIaRkYJsfdvihcUHVu7GMrdJ8gLfi6KN
GM9zGq4tnc7FP8LVJoWe6xo9Ykou0mnqqh5BOtNvqgvLkmShsk5beAie6skBG7JuyjcX5hsP1c3+
xFG+UdgUChhOJB59Z2NEZtFX0Es/WaaXbaiQZxYzV0q6vkIwV+JzhJnZJDocTRTgYIptFbGGNj9e
w9hcXHDiqpXRVPIkFRzTZvwdJaJSpiZ9Ar9ZROQmGxpDlS134l08h3j0BmRU2oU1VNtRDyjQiLii
ZX2o/NUr3FoUIXXZ5NuMeyadLsNjqM5qmmh2nJEtuiFErRzUK68HiVuDoQ0pOUntT4UUsW4NVvCv
Tsys/XYwuXSygmrieylmcc/9zETVn3xmp7IgJg+eCWf92evJ1qXu+PDMd254ic1coHs8CoCYndPv
WK+QuGSXLvGR172p+0QodF78+Ej3kH4ca0E2+id/RgHqxl+qwENzKwVB29AghiOxnEcV23eZvCN2
jTUUb5Zwtkn8we8TOrU3vIQRA84QndknG+HHYcAIAVNu8nt+FnMmKTY8y/da8jTAHfQy+01rp/s6
G88Qw6hcAi/6TrJx9T0RyA3e1PNt6irMAPw9iPptn81YcqToK39USC1SVhdKoz1OnJJtQiOnCKZV
pI8G48vWIVC1vH6uVNDvV0iptfqEL63+tj/T9KWkWrxrL8cD6Iyqq10ndkATsprKg2pZUiyT/fI7
IntwRido/IMoAfEE5Ay6LBbHe2+ggHnw8XRnroDF5Z22B2ysaenYMoUUPG0EmFt83iTMNK3w/MEe
p6UnwSXADkUo8e/KrrXP1ZaMSReSjfY3BiqBvCnwRKsEq+l52TVF2Eyhfbp4pqdl+oRtScy33QMs
PgNPer4SRAhGkYvo2LzcJrbtZDjKPHCFDjY4N8q5ZWOj2put60HRBg9GMANW66qKOuYVDRCSZCkW
RXbW5YvoJ7KdOvllo6xq3X4+7HmySR7y9mwEfqm3bXnONZZjMLVUh6+Htnz/ABMzxNomf6eoHPud
f3cB8joikO+64vizfsq3m7TXjOdRpqChgr79h3MtkeEZKdb29X5iS3ubrZwwM1v1azhVJPl4l+eK
9Bn00WV/GMOr/p24VeRJeqUD91eyn3RUZv9kY1IkgkbpDu3D0kHBnuDEuASbBWKoceOoglupWPWz
h6fIJLDHct0fJOBCVS1ylw6SMJB3NYMeBj3fcrbpCaKNJfkfYehIJq1QU5h+PBaCiQmjiVTPAFI7
N3GRoJ7LplKrToSzk7EfMNcZNP9viIlHFjOSERSIQEDIVZ6vswDP9aMXj7g9+gKDbDUYqXz6NDXt
rzzcKReW/HLHCzgju8/IzIgxGuuOxUDK5s1IGyYb3rxkRlgvudZLAyuIMrnRCagwAjejnq7T68Ts
/SB0ArbXQI/zBUB5OvmG+4x9zfbbhFsaolBCpG9iS2M3Vf8Dr+wcJIttR1CJsFHu9qextIgov+qJ
C6r7/Ya8LwXY4dTpl4KzLwdQJq5BECgksllGMN/vmPbXQT9v9c3wIFSeSBZL3TVOJ9zK2dg6hA7t
z0fg08eaqncVeGa6CGLblYY2f/Rptcy7thr7haBxldQ0Ya0TUyVYUlLF6P0aMoniWl5m69XFF8+V
OQTErd5oe5+kRrJiEmqW9n+aPEZFswvr1gBvKw03VnrR1i3FjuLIRuEkb2EJHdU9fiClKYXgoz4E
yugmbbz1yYGQZgAOD8P3CGQEuhOACaHwdwp/AJ6zH2bC/RkTLHxQsGXHhZD7PbBHvJPen+cxsgBM
Iah9BDi71oXj50rq5FI+NOPR7FLpXPMFx2FyEn2PeKKquQTdzn/j7Mf0Vz8UGjnsjo52XKkrjNMm
FqkDOPywJuFHm6UD0JSIPwMiFUzyvnc9lh7b5MF/5rq1C7QlHFstsnVU7Af0cbt8zUcFOthqR77B
ZFZKACCZJgqvzJAKW7y3Wg6QBpLTHWFXqya1yYY5WmgbICxCrn0ir8y0xvEVesvOnQTuaMDPHqnm
Pmzn7PhxfKSnXRd+/h6SWNKXldMPjhaqiiAd7IQv29kMB+R1Qu7zY/O9kZe8j1Q6fnrLAG25v2G9
Nqdqyh+XI2KTt95vCLKwu3wxp0i0gDtCHFyUvZgL3f1VKnW4wzGR/CrwOzFTVsfLG8SQaVEPMV4T
Is49j0q8z/rpzfvYvP/UwXoNtjtl92jXSx2+Dj0POhS8HqNi7YVM3cYSdt8Ce+FndnnUdEchqFLs
rlZc/okna4PI3RHzhfJN6G/petvV+QH5AQoCSun6645ewzYEuE4dA3BjCYk89GJn/Pgh2Gip5qoL
ekafwcwjNHcZyMo84q6snKJAxOEHlsntTTUn2Fp+tRyvrvFiRD40YiP0NtoB6x9UffnH5aSZIjET
FZfOZieDE2xyjlvAgSe9dY06NK80jkH8vlKoOPdub4WruoksonSXA5T8TVCCxxlUQrb0L39FyqsH
07Q2mnzMNw48Vn2sB9K7pBXlxzTCdyVKlawh7ND1mXsF34kRz79SFXvTpTO4FUf/ylT3yqdYrJOu
ziGuRBsomDfxLtanLdwA4KlyXXz7u/INDd0A6Pet45Ah1QQ2dzY5dZNd6FTmfCNmfOztxc4w74Su
Gpgsb3XicjBct6G01AWNTuKD2CKYsSudB8FAIjYXNTMN1VSjXIZOka9dxXEdbbuKWDh/oz4bcUyS
AjmhDDO5HfcQnK5RsGx2D2eFaPIvF2G+Utd5bIgtNxO4h55r3iTai3u1YClZ6UlgvUOtfbZ13I0f
bafm18NT4xyBKZgW3LgvTtQqdbgjxsNkUV/8qjlpLb7XRr4iV0oYOdBduAlJ3BNZL1JOl0G9tkkO
ACwd8Sbu+IsOo62wtszUSEW4UE+vw9RObSrS1NIPPFh2cFiUXk0SW8DwpdRibZU0+y3jYuCqyFur
vWbj5EmDgJt1RTm5XOhgrOtIzHw4VUURuNYY9FtCLewqltARaWK5meuv1OFUX2ZM1Yfpld6DSF0I
7JMYIRNDrnp3lm7KVDIYJnPPVcuFRpMZ8g2HB0HolddnnRDDeN1Wac6SulqNbM8r3WE1FQjbXq3F
pYOKL66sMmyUKdrIMnsEgobzpVccE96bN6vwc2VKQpNB3JPqQaYUcZckc0GtDwz/sGJeBBKA76NO
M13JahlpS29Scyt3kychYmfsoP09iQ0PraHB6u3xx8nkN9KMowKqnk4HqlmGMN+G3FNxq8cI/NAB
mO3sGR3cOxKOytgTsqLhqQDfB6DeP4HIHKqIb0O4/Rv429xPxoNzC4oRVJrYwX9H5ngoR5pwGMUw
0VrwpVmtH2w4rVUIezKx8SpySFWLO68MIbSenLDZH+oDawlnQAhBpUC09Aw+BA8IAZAaj9pW/mGC
pDiNyvBjGUsL39rnldXhZRMMB+FchfdKO3xXvYhyRcPd1aOQqOnF96beqYOwgnboIh3+Un5tuF/W
G9y/CdP2sDUA+/xvzYZnZUqR/AYBSIlk8RH7q+CBCxJASCWfOHMVJG4WjtA/27XvfeKiFHUMVpIn
IJi5ZVLN/KDtSxydGq+1Hk649BxckTIg5PL48i9Ez9c+0PUTojkvkcHveQfaE07uZPioJUnCnvu+
JVMSnncLUx3HouAaZL0cYNUKyf93UC9jbvvUcvjHET5MxjgkHqjQrJyJabxyCZ5gop2sa8klUNdR
w0ZQUUrDS80XWCkWpLBLk9ATCXZ8YqiedH7g5MzyiRS4i8rG0bNgsu+8GCQURdEYXNaE0DLBaZ0X
8R01RTd8KGzv0pol+QNF+z+sJ9Xr3OhScjIIx2stnIbxA54Z6lRubH5k4Voui7AbKcIZbN3cRGbh
KnPy9TrPI377q1Kmaf3L5bnLLxto9TJH8RfjDiLvxBC1MaiAOCE8+yBavman8B9WLM1UIAkGliVs
jNasRYRPrq7/8LtEX0ZpOLKAe0+mwuazLO01IMsdN7bvnD8AuRZedxtMgJBynoxKjsC0cX14g/m9
riBJUVj3Tnv9so1vR5d2I5dkIstzzM09mK8n7S22/XV3b9sPq9P6xbNmC/GtTO34hIx6ZMzwwdLL
VFnqnbVYgLgSpeQAiDguaaR6Lto0O32BM2ix0KiGPBGSQwTNtEwqD9ZYfF0uTb6qyO+hAcqNN/7j
fUz2Pl+YfqkJP+lcp+eRBfYigHgpDU1X9UKNLyLD1blacp+qzuk4W3iQDj2cAjlpxJsQkD+3Hxlf
BaCdf4bvFL9YEGc9d85xb7CJv/7o9o4d9DWmUXlHzPON3y4NrmQa9Yipr4Ub7zZpDIrCqp+b+/Xz
iyt41sVMqtSBlWDkVrYCtODLLv9wn5lRKhauE0q84fcN2S1tuZVrAIF2hCWwcIlGnd75Cq4bEhBe
QHpv0GsIwmhYcQoFVS/yTJ/cBke38s25QnElLs8vK3gfB5YajA1i81tFKOMAhXZ2pb18DuKZMSrN
OY/qE2WYreoo+KhEbxgKleSzzTYJkYmfkh83KFjaCSrgI/y/cjXkGxDYRWDr5LKuAKGZAMFMUZgI
YkubZucDglLMLehkK+N9CtHQJf9sUOidJzIJTwaZn3IdW1df2Hw85/GSFSovu6Qp6lwM7je3aLYc
rm3ZkvdbtEOahWBG+A9NlYBkD1qPj5qVqrhcmcSDB9yaFUxSS0Tau09yZkXTagYpgtuJKGxztNOJ
26EJCFTzh0Q7B/uDeg/9Jwr/vCPH2M4wsKqwThfpA3ZDHqUpz5MktqXlXjM8NVlP1IBTYZFZox+7
LTkDGFdmDuG8sa2V85KzbcghoGWfGxq1AYYDLa18BmqDXNM/iB38ZS2iiMiG59ww6HGo5Zx/MsCH
95EoKU8n2cpDx1O2COLS8fKY9WccPGHzSWKVPkI9jWm7MekT4tCK85MFZlkltRyM4/5kC73nC90P
SnZOHY848d0MLhyItILkLL106R4J1aQC7pO2usNCIzhz2JJVQ642Xv6D2uw5bh9QKMreQf3+773n
j80xmbu+v2i+OJ1pEJ8d/H21XjfFmd/Ij3ah2WpxHR5q5yeGSTRYo2BB1A56Q7vsWuYYDrOmxBWj
YLz4Py8U5Of0ZVSjHATxttmFlFpfx4HSA2jKmHFxmUHnlcNKIMuV81X7OyaorSLRGamRlvKVJG7M
3Y/eLay+T3PlIAjtPEqVixpkTF1mrn8lJaRcPxZh0mXewKXEKhZ84ez8R7rG+PBaQAOdkQTatMsV
xhAbP1d11vr7sw6gKnMb7McX79ojj85sQpliViZYBBkroS+lPcx5CAyjZhwESwfXyhdytiYeOuXL
KUKSGSLvsXOASmIlGhgRUn/ew5B/UsKvOczscUxFxHxbjSZV5Oc8sduE/QL2Wr0mMJGpmtzum04l
w0jlnGdoy+f2xKNo66gmDpNAjYyPqjqlkw+fGpiM+RcF8dDzEAgU7dNeLBUO6MIFgZmpgGKhNTOc
vMlfgBbqWxwjMhmkaXex2sBLqFeUrkaZ/UEnoPtiumlpmq6hhtOrwfVqsee//7+03us1sbm1MEWH
EnsRvpsxL7Xbs+pl+VlcY406rrdf5pZbXCzUGcHryPFlzvrZPQquF+l2Id4cNjAnZWnI+RbbH9ZW
j11Y4uSPbJGaXLwCMOQhjrvfuHjF+FcUx7Qh+FGv5U7/WWmQELhHThovAOFM8nruhrE+7FEV8LlF
eXoRKBaR8Z7vPVXSA7jnkaODJbOdy0RZGaJhf8F9vq/ksKpKSY84c5j1j7eoXcMBDLLYnMzZJxPH
MnlFUok9id6qo1WPBZA5Z0auT072GOquKgI3o1PaBZGlhYlXnPB3OqPvWbzsbGJVtc6v25v3Zi9k
B8M1bw8azX/ZgLFk2g/ISNkyn7lmryX/Ovr2VTHnUwMib+o7pqVp06Pw2NHHDlRHCLv08Q1OJhQo
2mchgC6n4FbNEplYgRWqm3zi+KXNSq5pP9Rhy9baH1QAv6siWLiO1SOgzLGdwsg17SrG/wTakDdB
NrZwuoyNdilAsxD45FbgjT4V2Ff/2ucQ5fetuxX3RFm/t6s3rrU6rvwRZHaBG8Qjv+B/TwCCTJCG
kVbR746h8XsrQGlDVdtB4aVKB7rm95dLIioNKr78s7SO6rZUaPR946XcmU/MDeNBYZJSmAD1bEIy
TqcR9dXsqiAT7LYSjVuXRTyWa3xrK8+p/fnhZ1Xh8BvjwRrQmfg2hnzTHqnt2/sZAZG+06HxHZu0
dqPLDr76QrcPGGML8yPz97eEkgUldXNOrh28W1lEI2AGCp7Hv5MzFpYfn4BfSoHSDX5yRWuzVaSK
5R613AG5/VbUZh1EY638O5xmH1B6RpXsAvhCpbVPArMnOBjflOPptLJT7MAQ52AzaG06US5VesMk
MY4rNi6rzn4VHEQIu1eg8YNXQ58jCmo8utIWLtZJUXHXOkJz+ZymuLyVnvIYJTq+H5Jgn0/biLFD
jCxVBkeqkyifiiFBI7zylcosD3X7jjT0VIgXzTwA8Dz07mLY84uScDfWaTfc4T5seCXuKNEg9s1S
529n6qbGPZhDGCT7n8Y4UlXF/I25/BKGcotKGK4zkwvuJ9+oBZIDb/rKmShvMl0/+oFtW6vE0+7z
91kdDVDVdsJr4aIyY5f2dF8Ot8QqtTHaDiHJYfPuAqxuvGajZcT8ES41LSqJblKOiDSUBGs5ACtw
PFFOMMVZuc4n+L7bM7eKs2gO64+Ac+aoXhsJmjlH0DkVUPHOveYUe7Sd3VAQKvpCDLQGv6tJbTxo
djEwdhEETfRooVEyb/aMHHmK0Ljr1do7oOGHQi22ZTkPgSqsgRKzlctcV5AK41Y1+om5Xpvf8mm7
2JIeJUbu3C1B5GefWeAnIMnpDDE5Q4Piy2xDC0S/LbWGVtvM8uNyVLokJNcyDxtTsHYdxNPygTQw
QkKVlNeLszgZMbX32TGxCjHO2GGZ9BqQfnL2lTqMFPGwUzQI63zZxdzAQX4MzoWQOB40xs5/Anbg
wmSwVLWQufMnS+lv7LGWKjfTyHK9XbwDXBfcNEu59I85hfZpWxuVgPh0LNOZJPebTYvI6fBz3CZY
Lkio4ssRzpuVtRPZMyV/h132GBHg6amhG9IDdJHSv+97QWnIdOCWHf24VMbgPXVrflp/9fSHRGSQ
KckZ0kPlbupDjOdkfNQ0G2pF1Eb4YW+WUrPxBceWcyy5aCdRInmWIaKXWc4FzGE6THFq8Y9pCaOq
Gc4LT21YlARvEGnnkkkfJ/Dui5Bn/qpkF7tCqvMAGhk2lZ7o7gUnw6nu0Lf1zcJzrEyJaI0yc0Mf
JpuPwU6/2RUJ5Kag9Ykbxy68mL5aJf0FY7MVVinZXu97gr/43SYtlf5X+YcrsW7XyA1NWd/5Lo1A
1kHsU1SYdPViM12fpx8iSQj+MTBmdsI7jYXvVZkcEqpK8MTywampztfQjfA9auRgBIBoZAqQfhvJ
1iBcn2v+i8JFUe02K6TDic9EovvszPKUDirvyPNt7GvToyFcn7Ds/BRYKI464INCR2kJEHDq6CVt
hMGFcI6rnVKaN/vR1uIBG8aEgrSo3uB51k3lIdWKVZ/u3MoRj/uJfd39Ffn3T+Ew2+l3aucV272J
ggjMMP1acp2Vb11+MzFdpBao9IunU6z2xSW01K+S4hpxBAcE6vSgijttF8amKbd3VD+IPdKCmgfj
rVO0XGjtdR6Wy9kUU0MVkBjQYltu3B1+HoBw0ulcjcycPp09zS9mbt8p676ovOuDeR/eDjLYnfE3
wuT8Ui2shmx1mzeeFSholF1YKTKIYFy/6ZhKRI5ienMh/oE/43RYXt1EBl0fmaSllorre1+RhxnD
+Jl4+JNSoA1NUITReJT5OQ2ykwCRsgU62NQrs0kdhh8V+8t6eOnTCLHUjyc3+41pLKvGy/8fya66
/7rmusaTwt6WS3oNs50zfxQMdXiS/ISJBWwmIz2QO5/o96obB7PfaHn9Tsry7WxRnPRPkAktQhXS
bX+PmkJi4kIY2av4/4gsWeE5lZuqrnoy03BeeuL3JmQPCCIApv+4z7B337m7VfxrIHj7M7IJP1W7
8qMWn1UCNqhTvfNr77nL8SIALShuxqkDmE3jMtAkqa12rYcqG+efKDlUte/B2T7Bw4YYW4KjbbfW
ZR8Q5rOI2Q0QInifFWvqCuPZT9fkdo7fruBbk9EGbYfMiCO+yxHkcXvEhJV/QPxnH47x849C1WbD
5pOZY2qUfN4bfde5IbP2KYKE6xvWQ1TgaZzCc4VVzA79m8Or1SHY8xS52wb/jcyECw6dHBNpoHpy
yqoYHsOnmSwlgcQ+OId6UOdK0sOs9IE6+srrFYRh0MJKLOFnDlJYrSXf21Aj/9myK0x6UNALrpxR
5ibmlpig6Kz+9JZofISEqyjTvWnrHlkswHbzrPo6B6GvV0lFcaqwXhRpueiuAwrpMIS7QkiUV9VC
bZzQXuIGrAXohSiAwocKf2wM46sTE4SFKLh8oGXzQbPdqBRwj55m8vmJWBkcmzo1IkjPEqePAbjC
mQnRHyLka+arMl5hWDrbxrQptZtaXtHvWwgcmeSWslH/p+6dEecX8Or4Z1Ser51gt6j1bK5KhVYc
R0SXksRG12M+2UTRKOQ574JhuAMMSjWZebXMryV5cvfkWghMdAu0OgapSZA0wHnhzQdqOai1W8+F
ZdMr7SwQAog3kslaii7NjxraNkDapAsNDJXxjUuy/DWpA05Pq3hUate+RZvjk3DoJFOcL1n8j/FZ
xGugYpP21g2o3Qo6D1qmEB15haBfSMe+lGS3/XLMpLe3qUpBg0VC2cTU4zVorQzaZZ+xbnlcoPze
skMNJhFPadHh3K1qXWFaxM9m+yI5JjSIzrvnDZflMAk+eIpiuI8x7RuL59dqpESssHosh8lStGWM
V3AaKjvFyRIk3k+gb+kw5XtAKkdHnOuPZKQkLecae0cDJ32OwNiMItyjt2q+DJy+4rIJ7kVMkS1S
EIZM2RwcrXpiq2KuSZdF9ndQ38HtqiLZbkw5Zz5pzU4xNYPqwIRcAnEuW485DiKksgGv3NHbirL3
Wy9Qf93vSUBL9VAgTKZpDs6qw+nytz7Xa2isY+RzDEyzHrjPiisz2GaZlVkqj4GGOV8obRNEDUk8
AenSOpMyv/FkkFHz7hhV/OnX/MChQCSCgdNxWD+KPQxyPuu3q5CZcnWf5qiyweTmdlgSGYtVesij
yUz0euTqj44ckZRuL145XbjT63t9ALWVAruulH1/ksoZNAmwQsT/wMFYT8drBnY+Su90qzpjYryu
QKBkZC/QMV9I4GrXhGbJwvx5/BkyS7PrkhaqY5x48DSbjofUS1Lv45+456qbJuy+1t0JCeqmHvDu
ALZyIjX/OK1gkMKQwfae+u0N2Bgu2r8WTaUUvkutx+PBSSpKuOLnzk0XLTq3CZCyYEAl2wXfrUWK
11PrNbcMcbDDrAQQ/T3fVGhRRPvE6p4HjJjpPwsJzed8wY+tvdrjNHVDSfA8nYhBfv5bbcrd4XbF
QeNQw/mMei0/5EnuXFGCkRKTM4mPIiUt6rTXgtALSyC1KeW5QdqhyBzJguYQ4g6ej9CuTg7R0Hau
YTDDff92u34XSovg8lPcbmovbN7HYpudsWghIliqXyTuY5b4cTZsWPYwDJwEm7m9PbF7nG65qzZh
Bvd8kMzYFbPSJNmbY2XInMcZC/LPT+Yw/ICvF3kMGWCCwPJacGjxRwlxV9XV4f3Gofph29FEjb5l
lYxrhZI6syDHsuNrphj1/ZmBrZg5F+99GgvZDLqjhZTkKxh42c/dKbJbcHHI2hw9NvQcPJpub3/K
XKO0im+2QXgFxou11X6EJLOBXXkzPMlooRjQkWSwUiVttRftJ8uYzE6HWvFz8Mup6/89Lc6CUtP3
zXt6Mgx8N1hD7UeFMldg7ZeYjWswBp8IolABvAjkTJR36QI4pkRZVqCZPKcOGF9kx+lyX697MDHn
AFaVzONmvWokq+AZXozyQL+9027Uo1uAaUYKdRdXFUwqGXiAknycvX+GhsOMAjuA+bHuTus/wgVK
ZSkR6H/ggu83ag5PI2iCDv3J9xDSdH6XxEU0oxCjzBQbYtbZVsH1LEWgKBYKDUuwEijWRxJKUDfW
NxmkADMbMYcToSr0Md3vWtHawRtoUDnNRgy6NpE7FT/x4qZ2s0JL+0XuU9uGH7MD8aR2PQICt9Q8
lDHvxbeTcJ7c6pbvzTQtsjCKlqpasjQztED3obcbG+UTyCc0VdH1bJXMN18rnnUYXzyx6S3L+MCH
AgtW5HU9rGMmPnUQkD3nw3c2TycgSBssDVSl3iIKEsUpRXuKGnTcZvHNEmXQHhNBTKP72+yy4qX6
+pGDaoW9/j4Z/RlvBJ+WxdzBAR64q8tp2VidoU5go5zjCR8VIiDWWoIHqvILP5aRLu9Zu+kpFvs+
hrMzvEm3ARNb14KYXfPNHZgkeLmSEr0TNKEGfDKQqvtFSHcRX4//qQ8lHPHd5VlyzAVacWYHvldv
sswBPFLFkZC7PvMfMccatb7a4eYx3an4OZEWmxs9joZ6rYlIgOwFjbBqBAQ9NsmCf3yYoWvu+soO
S09TUukPsNnkIySvnl9WMbQqoOqi0AVWFLymnTgCcO0d55XFCgvPY2emaUBO2bi8SWBWUB3pq+KQ
Wc1QYi5Q/SvEVhZ+l4/B6xoUYPXq6VZB5XlDhLqVFPr0zHtjmYYUZ38H3BcNwtfQUVrXuWNbK3Z5
4R01iNNl0KQKrKT0+zRn5ptKO7WinVW+VAD7blNV8cpkhwVujlzUIaFr4DhggQf1dwC+wf31Y+1Q
aHCFqiIVu/H0Uf5ouWe2DZSzUQZ52vTqXxh8BE8CB7X4gMVXrWIEgSClLYLlTqcbVeWESLl4z8/z
gB90VMU5crXzotvBu2Ad3mOGL1SO9rlTdK16rKBxJ5mbuwR5evJJJsfuCZJ8Ch7/LgVT8Jj7UMiq
xG/a9RhT39B9V+7B2LHkmDZ0DCEeD9H8Zc6QVCHvo7QZGSIKb2xKIDbyNVVzy2txqry7ZRdLOw7o
CVEckjNa6HKEsQdYOhjh728HVhgD3vPL3nl4YJEFNxHFP6z5SXV8vtw8Pl1rLdhpRnpar51m6hOB
7tsNFrapxXypxoOKDTLCE6VV8Rvg+zvFHTlEkxLXt91bUvrLAJLWtMndKz2dTITZQ8VL4nmyns+f
vapTgNX5Mt5KKC0cNmAS+FmNpwa6nnsFdzCRsIjAZ42d4bReMqZplkK6bpaVikgFBb+1FasYA4b4
u9ychrwr6qiFezrH7IrmXl3//1k58JgNY1B/Z53LLTjhpSrWgRxICzplz/r0XslECYk8tYH5/aG9
NbuiEJHkotIdosbYk+r4I4YS5NR0Sj+y7vAzH+47AHAW7XRozoF7AUK3WhcHB/4y43qXacixajl7
W5l/MCPoNZmYKvIGxJXMbSfOzRlT9soXaPfRs5JzJaLcloiTSZXkv5UQsGSHVfpbHVoElzrcHFr0
Tvx39iPS/DqhkPjCIJRXiGPXcY62XJuG+fNTjPSYKC51uiOygIRmWH4R186HB+L4Y1xH7cb6X70w
G9EVsDnc3TysDVLCiNYFqKjsHwpvZin4e9NU22CiVRQBWXNA65PcV2wxPVtB2JTTg0wF9bu7WKj/
KUayEDDGqRT6vloi3tvUIT1OGwGlA+gj+T7XAh5iJv2m9vztNOEbwvIbVvf9IoN1iNdCT8S/VLYN
7ouL801h+11ARMcYAhhcaNJn23zSqdrNEzMdm0FCSm0F2XpO1fQT4Tgjws/phkPIrV002XCtHNGS
aeCMZqqDkyMuwSa7YymhnJy5qCrEQpHI7H2y1nvJ+f86ByoWO7+1Vyqxj4zoK0cRGyRlvZgL6b72
lkoD/ogAOTxtEN48rPMzcUEuzX5USINGR2WwRjva//UnO32vUapanIgjqY7mNGl2mtKkDUJRd40I
MCX5IivnLOeB/nRL2wUqKb5YvtA3Y9BdtB1gnmv/VGY2S7hzeg2BmMks4LWzPFi9kKd1MO6TdlAq
TUdVeuNjL7D7CvzJ+iczOLML/ICgGhOgRq2ySKvSWiMIF4iGLyG3L811lhjl6aXCFaeFKlFNqMtm
atr5+eNwqh+R/FDa+q+H/VuEFa7+obnIqQmvkBtg6BjfEjk/1lK+DkQ6La/Bx1WT0EVBXNJhb+Vb
S9kPkPr4Xo3mzRhyHzRWpoXsYJC+Gru+0HbVp689q0jm0EhkZqZH3tGk80RI0QCPpaW6nN9AR1yK
2O3NId8dk09RxzgAHVsPE65OI1Wza+GXm4SY44OgJjkjJj8WFo4ZjHKPPS6zYP/4Dg2VhvedKYY6
pmk7Oo7Wq25bDFqzT3oLikFLLUxbuDvEp52e4lEHFWoEi7vzMuAzHHKMdUtlEk8qnDzPtySMBZAo
CHYTColEXv0ZqEkzruF6xu0mn6lhyIIh/qU7PCQANadTcjSYXvCtD9mOk40kiHhFItPD0OG/lDb/
j4joYmWYGi2yduFvC4LShprmmTVqOO8lFeEB+qi8A8pFkkcQWbOGyhg8kiAKaCVZGbfRMnsshzF2
xyuiXq8k2QfhLwGRcfVfJy+lHron0LZR8a89a+s13/zrbQSYXRTe2MUx3kqPHaKpqOFruRbta4zW
1JJaWvXFuPyYxHInxRhJug+Aci859rouNGHw7o83vV007NX5QXC+pkRFEMyG4YF8Wn0/5jCjHSHS
9wJH3V3ZA0zalu/jMrWt2CIlnq1SxkWpaSIK8EKONak67o5gE0Ds0FnWpIPSvfE/jisvqaUJxM8t
SmC8UPDo9GSTlsWvqDWdYqRcVCnVBt8GeHJ0KHQ0ul7OlnzQ69hAJauNzvCXtRxhWSBjvTsb//Wh
RxO8SIkDNmgS+CgwT6h50iATBwC5sJG712o362gLSJ+0XUnUBYH3WmxHamTLuCFaqeMDhGta0YD1
Ux0sMl4SnSubr19UpKNbH8JmmCwbLTsFt4RwF7IiQ8K5tJYEo2zF7EkeP2lETeSIfvBDZg/Dd9N+
qAVPjCQuCGw8scOagw3NminUyML/+SLTNzq/f2e6/jR3us8kFzXvjQcVjFTlOHAzXjB74L322LyF
TynNPzBHKYGXCdSY15ZCsAlTzrRbviEGR2vdr/UmL5hI5nA09rl7m1f9oHbA4z/7kaqPM46XRHFQ
bX2oHwh5DoE50UTdJc7T/2iNySk7TzXQH1JtvOsLPFSeqki3c5RvolKGrmGsKoeEWKDqvAzPPmqr
pAtGVnfcBPD430je0k/3tvNE6zu1Ds8EiKLLG08Mg2FytL949UEZyulLhe5XeQLYQ++H4hG7N5Dy
MhRwA+hyoKOiZhcTTS7oUsWgO6DX53Q3E5YZ9lOmkgbdJXqd0w46VsYDOfI6PfUxWv2McBTavXW0
LJ5pihaS3eOYbNVAkLQ8n11Uee3+RxEkXaF89P+VWezbSvow4xWxTbilb674TjLt3uCMBHLoMTrm
K1WBtyapFd1kv2wl/IIlsH6y3mLTtYtKy03snNIIbx29eshykHb449yVpCy9yCnWPju4gpGcUAB2
G4Drh2p8/oIK0Wrob5WCoce5H1hV8PAMq9zjMajcitJ4fruapgevcm/ApVLRgS85lJSF5Mx4uF4K
PPN+0w8n+MYWyvWZITeoxptS3TbcE0zcGo7wt+QEf45Lq+yFrZ+be5MuQ6B5CfG0507V69CLqhBc
ajmBBPsrewrJoQJkjcjxb7y47otdAXEd4EUyVTuSKqJmYDoZ/Q6s/xsq3MWzDN3XBEVm78dIs6KW
KBTTv6K+uPN+Oe9ob+QyIc/EVSlit/8T8zg2PcXKoCGrl3OnZZZktpjGUW/umw8I1mO/udmkwhQ1
JuLQEuRcBMRPPsmdhFCxrC1mw5pge5RsKLENAWY/Hdz+rldkSbE1tmCp011kKpw0kNMI84Guf/WO
yLAVkXOvuuh+xHfohI4+gBcpCEX0x9Edapx+rRbLPDF/rsitckJydAMUGQGF23ykhYEmEpU7Zhu/
9hU33j4O5pvj5SJMMF24yHzhgRn6/t4u0c/r1C71fl2DZs6msIPvFY9W/PhG0IlcsJoTwc6/uHyt
9nEOMSxwSq9FurMyqAExFcNoEyiASe6zgyNlzPjN+UopitVkFdTT+PAbX7ghcZIJBlIBMVuJT9cc
E0jahbiNNqGomBMwVmLhLtYvaUAELyVLW8TRfPWY5aCkS0Db7DKj3+TRcG73ejBiBCnzBI9MClCY
/ZL+AOF8TMyPp6dOtwtAD1DWiZcXOekK88loVUm3cTv/tVmEiNxkk7VkkFLl42ddvHHogXgNHdVm
+BalfCFLqB5k9+ESWIpGV8XsrjailebBsXJMSOYRyM8lGE+LN+tzt5TnGmg4qWDH9esUfQpk/Hiq
m2S8E2Mkc4LOTxyRUVki112i/ylj+piP7xCmIlpdgJYRH6AGkzE1xH4V5IVJ0kfYqDDtEtANRTXd
FJhZnr0YXzga+LHqqD0BfIsbE4fpIXxfq72EbVY5nAwvEMoD9ls2l8vMOq0IhAbs0gU8ThCOfrba
DqGxxbiH5s4mWcadlpvCgqTwObeE0aqiVEXd8o7N1AqO+Igbo2eVoGmNlAyUlEfOy7IanpiysFtt
KfmDedHhdMwWioOmvr9tT0L920HNGUj2RBruCIsrI4IklRVYWuYhBlsWRH3QySpcRmAWo3EUJW6D
xHrQQLuUAIVFYXwzJ11BMoEEB/J5dsN2zBafP1nfH3/oRrdE9e3rDklAGh9V7jFiXodNqogA3bvV
HM0hZcwX340WfVDln1pAzfHdUF1UtwFS3fQsU8JR9I+qVttkq9tfAGg/yS/ylZQTPg6UtnRlrY77
Ut8XTgOO8EBanQFzIC2kGqgf/g3df1j7xRuLrIebW2etPMgS5cgyTVQxhdKDySZzN3etPPR01ykj
0BiC0yn4OjEF8PsxME1xz2wy8dvqURQyaMGSuDLWFq0uAj96KQkvPtVeBMLs/uDPJPf+yg945gMd
qynwXyqYeh6k4NsizEbJ4w/aqWF3u1fhZR0PrRT/9IptD40T5enLd+aLpZ8BguYUHlDizV/IcFpp
DbzbgAP+A133VTYK/O5FAzVW/3fL+6xMPLOWVs5Mre/10xh6XPH4rHHYhO8QjcOSM+HHnbm9SszJ
UTQNtgQmXPOZ24lTfNVAmEdm+5HqEoRuDsgMLfyiVPR40AK0ppWf5i71YFH76zQieC1XOY1hTIEl
Ju2aS/vE5z8WepiWsdEsUp4MnFjq4oTqc2sWmNgSANIRbXoh/Wy/WRB/MOBGygsJFHk1F4DCRUYN
KTu6CiWvGeYjLyBNHLxM0yeJspw5Bvvg7ZJl1q+mQUdTqsibBk5le8yNTgR7QDFVPW/2UtGLBnlM
KA8pjPA3lLwdHEFWrLQVEBwGQfLJxzeBs9nGblENLxzNhqwxsUugiLa3t3Ohc2ShYnDpcP3R/3zp
Md82N5C6enhY64Goj+ZWXoLjsZ4jBCevPrSntPHgaboZJcJ7KXIsbgv4LIfYEetsmZjUjkQlTjCQ
ytt4ME9+uISbEG4fXRvDwsATIXUFAdB6bkFQcJ4GQAuY+sbmYpRpYi1rBJhUPcT8Xo1A6Bo3e5fb
n+TzoF5mXaQ2GNQoIbbzDRnfTc2gA0y5Nqp7eSYeF8YjTB2Tqc3eQycxrba3F+Vb/G2tFI1uoAJK
BEGD5l/yM7FK5xDXOalvftLfgA+cVrNkGzdi49+fXOZT7xDcTIj2LPp2HMqfFzfA609r26yom9OQ
K+bNsZ/v473v+HWagJktHOrpPGGqoQXQ5Ra5w9E5o7vhg7CIoOb+SG/IGDEMXaovwUbnKMHO9BHj
ZeriCVjr/daMtbmZN2JzQwIxSSur4M980KD2LXb3Xlwfy4jkkORd91Va4yLQmPTFoopZ7x4xOF7e
RhlEQwGSeF17MFubACqqovATDsi9mwbPY6Ca8zcGrx+Fwo8sPFsh4VT2vj/RfH2rDAnlINugkGfI
/KGtShR8r7SzNWjtSfeDWIpsUad97bUwaoSW+c8W1h39PQezLTk6aHP5CEptnTn6M/R28/4bB+K2
prNxFTGzO1MZm8djfIR7f+0c7WACURUwp6U2KJ69Btm2fCWnwE252ejUTUg+mFN44pduebMSf/oR
vwmcfPKaTNdtSLXxDhpse0vFtHQcKlg/PlnyUzQ1Gr/k/+awu81CK+Q9bWcb999pHzxH0o+KM7Jd
e+qW66APLIlgENljHWHVWAt0oAa1FOMF7C5d5aJe7GN+0skgNCkDNZq7yZQCAbs4qZ121SaXHzCi
qO1JrtbySQxC9E14GKL2WjygwgyXqivJWC7rZmrfFJ7UtVjpd6uJqdx5c+7WS85xtBpxNfQ/h9Np
SLgIKAyxmVqMgS0lKMjZ1s1UcltQBvmXMdRxC8N/+A/eLy+gbj9bKL3WvWjt19xDcPIQGvuhEinl
JAYFdn5Oy6PHPp+QU6+1cHidYRInpM1QKUo1fHPMq7fF16W3Wif70+/ytTCHFvCRnDsMY8b37pwU
faPUlp/3nF35daz1fX6VNvWKpndZoFH++ZEPpIBQiC6nuMxZ0HgaHI9A838skSubFIEqwH0A05y9
29t762qa6TLVl9NLTcl+jaBAChEiMYoCe3DDMVTMInEs4pp97fy1/0b1s2XrBQZPLCblDfEtOwrJ
z99Y/c1omlHpG3hz6kJpmkwkuvL/TgpYI4me/lssXTzt/OYLLC7waGkf/tC3YnWX9GTKUepW++zY
DLjwz2VtaKv9wQ8Wmv9lMHp3z5ZGLlQCZLSP69zMkterU2KyQMHZbXpn/Wi2C46zSYUKr8rruZAE
Jr10DLcvHWJGNjfr20BEG2QMiwVgPwG7rK2A31aZey/9A158xmlOh1jvEiFmfJIrrSo7LnM7HPPw
MNbQciaPKguMhpBI4kfHi5FuSLMPG5sHQ5zmLsmTwut62HEPmGiAPPpiv2jxc6RU1NtmC2i44vqf
7qImsAsJ2XHCsY9YVUq6gfq5lgkYQz3AZrRxSw6jKqVCXuZqMXMSqQX01rBngrTFdqCVx/PPmAKx
XVbAmyuCQvANl36vadnEwcKyCwnE6kF0DjQKgVUD4cnBixDlvWw4ITfCassqN+FYxFrqtNDZdhZA
dItga9nOJuQ8PLeBe6O38TOO3Vlz1rfUW/thCa9NAIaDgOn0IaaLGdfiWb5u01XNY0RbVLVc5w/O
DP3/ZLy9B2LUmAPDEZPZ4wbLlmumqGGoz3GD7azBLO6PaB/3jwWS4E/bMaKQi4wu5n/dFpt6HsOA
g21Rly2GomlLzPghE6Nw5jlYtdspTk5Ku/C7YR+QnnAccegg+URcGRJcreMLi8YLkv3UB4MLlFJc
LetAe4CCdmWzQfSd2rnuHEVVBsHpUyraLCrffInJkLnyTMdoYpUjKyKmuRjnXcDGJ9bwuZXKJONk
lPrLCTWZdzoboH4cPHxLHqLMJGvq/gH8LtULn9lJMEhhuGt+gy6ztMMrRykW2u56cD46R3mjERq/
i+8DPxBWtMdc+OKNYxBNLy7cjgd48IC2XNEiiMiKf09quh9eAogr4IHSK8I9t8eR1bvGDDT+Lh2l
p7f2L8MxpngIQJ7AsFHEOX+VIeLp3qCYAEGQAAfnbGOWmcn/XTD7fg2Di5dvPvGLycSgvFOUrR58
Xs5JDIkLqtDCcLYGAiuT0Jhvcq0Y/wv8MwYqG4i8tel848sNddD+dGMy3E1WGYBcahxV8mUIDIVw
MAtlFgT0RrrSqTp1pBuWzSdK8QrD8fxwmmEDzhydItb0Q1QH0skuSrdsMpjWXoNo9r5HHKAiH/Wk
S1gmNHrEpea4F1q2S9mrIia1lD2bSi3wd24gdke3g0LREy38z9AZsFdNri6KLWfhLcj/3P381hcL
6gUyTzwP+lZ6kNGJvh+CNWRfkN0IoY5d3Nz4qZc6YTDsjO9t/GfkdNcfzYG+zgBLYL4IxJLDOzNL
ZssALsMoOtPsiuASNsoRp+cGi74+EZTNhSf38FiNtmE2vT2p1hPoyiYvOBi0F6RJcNsMbQZjQ32k
ZtNuHVEp5HhH9JyPLgqk1W5gp4sB2m0iU0jKVDGhGGXulqRmPevYYCbZpgOOdmQkhvJUOU5672Nl
tQdB/HoMzzWsJUY+tCFIrakHZ8ezTT6OiWZX3IXy3pnziWCpcjsg+U+GAXrQ02vU0eg04oG6zOyc
dDiwqyZcUNhYR1fkDpmv6OKsRDBqOiAZomHLWfC5VX7Wqs/n11huDlNT9wyDIC2pJDQQGgTxyNnf
0Adv/hJn8enPUTi8u+l66vYIFLcGwtGft3CJIyjXbm5+OPU6dgktrk0OxRVbDdyfljKR0YXb9ead
mF87YXgGbPFQ6VybXiTbBVoYULWWVyx4IssoBZ+ghEuMcT52Jw87+gSMbBU3TaTd5aBj6LEAYHCX
Bqzozka4IL9gHjg3QTimDh+EamzLkGSUwynP6Jj5AzKlz45M53/JJJ41DpiUo351u2qd5pk7SRaj
pUdK9lW/O2IeDRK5a2UFRocRyR+fFabIbSDYuK3cqFLFVFXzyzd3aj66Ag/+olVyc2GofiWLkPbq
Q/1GaRkqNYq0N4JtmX5FR1ydzhKev9CUzleFmPcrFCHqZNsH0XDbZTqe1j5dDB2MenN+kiZ/u8/4
+e1aiwKG3nqg9X4kkd2XeCtKY4VItR7OSo03D7zQV/L4+MREmhQ7dKAngSzMv7SCcqm8OrbOsMTy
Fp+2tywwKe9KwnOjdm+JyzUpXoS7waNXk+bqvIA70votw3qBNlMKtW5AshZ5r0biV/WlydLgmz8R
0VrLAizYLt35rd8R8wQUI72MTdOR6ka9JrQibF57gvqfiHGcJZTV9B8Rcszyl+UY3572U/853WuQ
nKPIOn5NEgQ9bamOpkFUB4O8SN6OrvJ9yciG2wCysG/429QV9+/75I9ELUT1aTsHECyxerwVfmwi
Q/Ym0UW4q9RMfWPEDIKqf5ZZzOkpJGhj1QfwzwFU6nuaDDf+mCmiQGV1a3+csBr7bPpdjem9sEub
hqArNeJ3RBTm3NRd7gUfrTb3EPjfgmXOQI+s/p9keV6BFK6HGdQqBqzVbin/4dmc2uu+sWHsiDtH
tto7UpXv9oC1A9nlI6cscitw7RUC6cfCzTafVOvec2EryP/4pC342vftIZXt46mf1T+HmsJh63kL
ihi104Ofp1IyTOMJ42OFQH4N/KhMrv2s6y8966yATjLtV0uwG6jEPivQ+/0AbgWatXNrTsN/Y8TM
3vnvSDmoFl5j43VgfYcUDPX3yH/1/wnfLePJKUQdFruffdJoSIIaAfJOJciS7CiTlLqLdHcbXc6D
v1S5EyL6KcTEf2HZaP5gHLPk6Nvr6yM1KfP75SogzOA75Mfgp77nEbA/Spj48IrQe+AZWR94EyLf
Up/jBUsF7wS29BuSJFDsZJrPCTUv79UOMdAee4UzXXDArBVIACAd9UtS8sAibgYEfuahGdDj5ub6
szTPYyT33xEvhcFy3nHQisYZLYNtflMmQdRZC+hohWTjXvD41tLYGXYO/krEGPRArASg3IhTYgz4
rT8oJpVLpkaSkd2z6P0f/DmAz5JvBVK6DJ1vnqszBIgfuGyXNnuPHXjERCKS8s5PWqCNoTKqVx3b
CeGqnVXvqk5GsUDg3zEZIRbMfs1xhdaTR5sab5eC8c7glAngDDhe5gmPAi/9Kmt7gX+RbUm8UlBU
ZDLs6EwRdvf5MGvlU4+iYB9GZxKdBURB2c4ABeGdQEYcdkdOs22QKvRZnckTF6WvlsnazisnKqAP
4bKzp9XwgJaRiATw1EJFPy9lNDHvrWBrZN9kuwiCALy7PacEefzkttnzvn10/c9OrgXNzYCtZXr6
z2GHyp5t1MQpPCxEt8TZhEBdIUWPD8TxiUw0k+V5YVCkT14xpdf0GT4+Y6/xa3xzQeHIft9oz91I
H5LVxdkXttAtMlAVg0/N6N85YdZ1LG2EmyIrgtBA8eOVsCt0F7M8FJLdZX2/byLEETQEF19Ib1Tk
uLioE2H6B3bZsUmaLiJcE6LwCu4p1ZfXAbSTXO1CVUEUtBdJtCdjnHTxc5v+2Jvw1r7TElfBDFd3
lSooeNGi4HIuQnV8jnFp/0DNi2itN669o3RJMXT96y2oj6BvRrJjQn9l2koW/YBzM56qDBUrVM4Q
GhqHX6TIMbj/1QFYh6f+Rlw6SGu+pAUytXwGJs0Gtl9Al02oaP/LxaJrssqBj+xWQsdf9XNFTxFR
DxoUcKCqU/yCene/cYXtn5AM9dne0ktiTcW1celXhuJd1/4H0N4d/i/yQDcaQrx7v+1lZWaW1l7i
A8xK9nXmxoYgdA/RhwTdNM3joVY1OTGud/Kl/BTypnokE/Bh7bmsBY56YbmxXgGPUPTeRB2VbnZH
YKhTZ6kMWBGkVgQCj4hpBB5Bxu/1RTcFvoV2Z4FwHQM+AmGIgMkiEwzPRTavCbWhubulb01qorMi
32CrdjXEtNkTuMi+esVEStY3e8VMUsCkCcodNrMe/cXepyf4jSD1DH0UOY2xu9Cwaiggg3mIG5a4
bdvdvh6H5/UlVTiSnGG8qO6+B+udqoOzx7tL9g+KTZ6xuCn+j9GcDCjHsR9rLGo8vlCznyIOeu97
NRyk0yiHOo0Ty5ZaIOPEbk3UUn6ThqqA3O4OCbR1iQQPo2KxGIiog4mjNJR1jf+/XD/Wav4o2NTf
h7CjeEol2KU8BNJ62ZXvoVs5chka8gBthWhiP1nJriGXHR8EtHiLACnG3x/Q+kJDwx6I2Ce8vvGw
ezSyNM1QW6CM/x2sgD65ZD1HV+0BVQVfml//PFYFtydqlF3M9V2uDmHRABotKGUFHBovWEkll4pa
zeu8jUi7noNsHnNiR/EiOgiPLtSVhCA7kBxqSd8ZzdXFPGbi/qBM7cnzPZ4SlB8kgeypNqWKxXDv
RT3e1hNaoF86hyXWwuBuGWHNb5NLxfl6N5Emy99FHg9hkrM9SHp1HUBFxcGSAZUTsJPqSRmhmbhL
tQta4EyytS+vfdICzNT7TI+mGimiRkpMB/pZ2xTTAwWRSQu8pxPbvcnPCEnCCUsTCrv+UaIXjiEd
jumKWYFqb6WIRqfjeQY5+M51jMAUxvXRMffTPC/5NokXLOMZbeOP6Cx3+W8hVol/u4zGWBAcl9++
Xb9nvV1e3WMjeMnp63uOikl3lsGtXey0ee+f9CqKzGM+q7DoGj2wMoC0/0baEgvdPmLMFTb4OD2k
joyRbeYPPTiki/XhPgajZ0fJLMFiwo0uFtzW/t9QKkrRvG8JIQIkJnrUwKvleSqz5Aofapx3j2/E
yKQdaXCZJ1qaDoo/7vsFnu6c2U/gFlDNXQJhth2EEj1sv8WV9FQZYLlvZ6/tD9oLmu5p1xdTwcPv
DWvKkH6keWtljVBqz5J7NOLpdty4XxWZYX1PxACDNMm/Uk8SEkYjS+I6XBohRFQYILbqmH8eHOd9
JNNnxRMcDsuj2pDVTgr/KsOQRx8WvfIClcUvnZPVIKleOqmONTXzA4TEVSH7tPPqJ4gf3bS3/7/2
G0QD7ByzoWh6hJezEhtlX97MZhAGZopLX7FTcic7dlDLJFysXESNxEtaJsW65IJE1Ua8B8frm7fC
NLr4oDaybZgTXANAAbiySYICtqnu2rXd2uyMHPstm56X6CRDdZqBsDHsV6HkK5gHMLBzPlq1rYpP
Koz4jUuFjG8VrBcaDPxmcZh/S8qejGkboxI04AE0Fwz7i18Pvqx29OlwuPfE3DE5eJgBn3sjXf97
sLAuc4DsWOOYkAqi0q9UF5jVlpSllBFjUU/8kofLvGCAB6gyPXEBKEQPEYBbuTYqo+5vIz7eJgqp
KGAM1WZ6SnFaA7PNlgbGkBQOLfzoX6kj3HMBY0ohJyvyfeJjtaybuz9wqGdt//YEBZXU2vXURKMM
3LKel3IO4vXgMf1cJtV47sEA6qIsR628a1iPBiAXzDa7YRAnngWQoXZ2S6WlDGEvW5fhjibeh7va
u6CbBm+RsHTSn2/dJsPiKU/0H+/Ludfy0veLqVT8vuzVlQuAnrIm/RpSrKPHi9VzaN7JgaI/XGHF
XLFttj53PE+B/gbfyDyNld3KeNBpTPPRXE4JY1rzxpIVtgV7UFC/Gi2gbak28o3bDHL9C+aL9+xy
Mv2KSaXIy+Vv8iO17MX0a+1yRUdSU6c5XhfMU3KdWf+JtHZOSdeed+0kdmb3qMuEqh3LCEFT92sL
Xo49zvbFWHR/LhHhHipy/FG6Ty1p6ZhXNxjLk6a/kKMWC27NABqHvSWx/LLwQRM8CzEDymz9u4rj
2cm5e2HbQQLard8WiT2zydunFaZBwoN4zoGENQ7Ue56XSTSsK9Y7RJE7MhMIrzLLBcBceIGm3N88
IWSZkxqRaq0BUAVNBrg8TheQ89NNCOT7oEIlN5n3OeV86S2vSYdCDGw7L9D2LmioEZQX6XxDlBPR
ya/CVZllDe22rVyRe0IDo51QAzz9i5BU9+1Aa5FV5s9SXjX/xXyRPJseW03rCAoCwZ38el0fcxmV
9x/D62oy+qiQJViTpkTj5ssx+vzpyig2SAMeuWlSuVbh/t3zSl4r+z3pQ1hFe7eOXyoSFh/psYCO
eiVfDkUWLExpPkEkGl08P4wz1tmSPngl1uabZiumOD3QFOKmJZLjJ2WlIEw8cbcWS3lvf2582fO4
lGIvG1edjonfcuSgXj8/0qAohPv3A72SyB/GsLnTuskCYw1UwkxYp6DxSLL6aS0tcEYuprBApchy
Iw6URH2OSDoOrvLC+WRf2u2aNg0QNNgb+DBRnk9CHqnK/grkeLK4seai7qN/2xVvVRBEOMZ/7EEF
/g0xvCGXlD8XnATBf98QRAB6UUdLa5CNB3pcf9k+nDwKFv60kP0PJ9XmUh/qo3LJcg1F87cJI5Kz
j9w/DNErBcpeK6MUXgoapP4UKJUWvMxavYf5vtnnVugenpVGI5Z4thiCqO9uLyKdeLpRMu2oYtnE
JpRHL7L4Sc+SFEJhDlmD0lVnO0OpqPULgwAXaYf02LP0PFrWK28jESYEZ6sBY+DnSEnYCVYAD3Hr
OCUBCU9Uw3C4pL/khZfamnxBd5gdLzMc6/MER8kgnBCwUnhTxrjNzX9bfvxz7LwZmFkj6nLosjk6
ZQ8bbOuFDOP90pleLvZzLE/Ww1feqafgeAqu7aIcUs0meC2919YU/eHjmC9U/MexwIqAPOhn1lwn
mgAcaqrW49NACDjqVvR1ITcRmEAlCMmERyjE2vKIC1O34HEXUu7U9DpAoZkQw1BgM9pHo8ClovC2
l33cg+SpZAhwh7bOYvMRUhVXwZW65moRlgF5zJ12px1/iAAP1HIwckMtR4pBpzT47zS5IDcVBjfk
eVEW9qbUBs063p0HpGCMMSU2xO7dSRRPvD/Q50cM0Z3shy6cKsR6eKW396Ogz0OTey/EllPAR+7L
A3GXV/chlBh8TZM7mvoTy0unI3RjV0X/1kfxrIsdzqtq5JB7tRXQSm2/yexQ37a2GpSZi+tfvWwo
0syjneN7lFVdgj8Nt/hoz/B5ljbWUZYpSvVIFQq4RfenvQbsokPI2bzEv14y7S87OmqbY4xodvfK
4QFUnKUJY85J25De0YXcQdcRjrLuOnUNXaZgHwMrhH+R4PtfrXxcKvE2waY0wDZ8XpN35ItRoEkO
LxFAQolCPQiDgiSymRxeh2OtO/Sq51KJsekN7UEN2Jn0vg+1MwWPVRpFO85HChktz+5XJQfs+jaN
FPbrkEJmNgNfqx47+8l0A8sM8bhgAj99IFHUOD0jtcBrZU/97TS4j4/y5n7KW7ntzQd8WR5Lkoxi
hud0bc2FqXMcFEhJsrwb+SqY+SPVagk6BzYy7L1hNJqbRooOlrGyDaI5knBYPrC4k38KhILHj7Ze
Yk9E8PwhUevK+awUtlYcs/nEQbaGz7/E5xXnHD18UODs2hliJm5iL0ULEpy8VB61Eg8FIPbAEBlK
ZXqi2I4yRDRj/Cek/6Z131uiS25H7d2Drbt1YRAr+A57AT0Oij6nmfr6BR2FZFCXAqlu9hMrc64/
1HErPYM+Yc5AdmdnvJt3rwMem2miEQiXU8NsOe9B63R21U8frNg7kGEzXdr0cIf8l2YhgqW8o/sL
JfgGVags1dsgIRd1tGjbotr3ZpTqSqrZH5V/Cv3XqpNVb6O5cjKjl3jpuGUu7S2lh4oKEb8T3OQ1
JHrbn5Hgpiiovq89THj74lHCTtXoI9VhWiRybRW+oD3slhdYOHK98wgPMZmVnbxSEVgEL05E2C1e
srZYLNX3o1BzzHC8ZMdhAQnxFbHXVpTKU95GKWNuZnghlbC420Pn5hd1Auj8UWXfy3pFsy+X1SFi
MRcGOYzwBhvoN+/Hdw56O4+maz4NGQ24u5s4TLdZzsV8JxNHITvzn7j4rnaZxbDv6Ig7EmzpHn3S
TALKPVKmlV4MmzVggc2RZJBG5HQT+A+C9Us8IWHBzedeibRO0TOv1RbPNOswhSehPa2BB/CHW6/q
0BbVEErYq17+vrfrDVQ42ovUa3ScXJsfGAT7o9i+q5p+95g728RfgJ0Pni5MIz1LLtMdqiUWsKpD
iNt18tBkWdQwoRm0JiNHTKXs22Rz9xuU+KqRSPYcWBfSgUCNm+OQSfxmMxBedzLd+iwl2l9f+P/A
RQdryEpkK6nBxaxhgf3Nkr4YHMzSeM3K1KguPV6EDprN6ElE0fMRm9jrlikrO3dee1e/LKBzvst/
VwuTyHz9QtavBMIBog2KrsMktG7M3MEHf1xLdMwgTvWi3BylO4/HuzHgNCcuv4j3MffNNlmloEKP
FOpNI0T67CXZqXbBCT8okp3HUUJFOWvO4COvQsbXpRE0qhUU9OZYivM7iKEV7UHmIoqT7wq120VT
mMPjZegZhw7iWXojnUjyasK+d6KCSn617LlT1SCCV1olKNoyKv//C7LCp5T8OON5AlBEmIrvDasN
pSYbnx/gJHxjXwXpYC26QKBPDz6yKDz+ngOhv6HzSGIh49Egm0Kd+cK26BwFr1Swx4ue+Zn6XK8j
kiy30w6Vsla8XHH9+JjZX+dZ6pTAQGngTxie3nwF5fgpJzr6dmFU2N2bLTTsFMgVQTIkFkgTCl+u
H5DpheorioAm5xk2el05BNgEFmMzx4N07eH3NV7bX380SUhRft/jGsC4LY3ux1TaV28ETilRTy8J
e+xBa/K8FWAsL5MkW8CzkHhiQkorJhk3XzTuURDBeKXFuQTDjatbaBzfNN9vI7Sb1XzGyVeRPDqX
CL6ihxfm5xVgqBJqnkGttP5zJZiQZ4m3p7A5v0jqAigO+H0wLtU/0y0+SNN2qjzW54KZ/Fcv6YXK
KSVK6vJ3gSls6L97pU5r2kOeG4NKRokIiFCTYihkyv5n3YVBq2e+HpElH2Vce81069vCT3n/c/JD
sH+35u6kbgUVxzLx9RiAK4HToGDCZYbudbi9qXqJJEC8ITS8LKnA+c99j2/v+qSfKFeOxpMS+ZJz
vTHeWKfWeC7WdKAkwWYmSavYfF09TKsh4Do5nxOtj4TdupaqZN8AExsnKNtw35myGbD/Wpyv6s2C
uOqqkWhVVx5V+enmo/+pf+B7HUBReAjpGuQHuKaGIOMr0EfzFX+nqOQ8P8ZBZcT1GXcaaSsKlytn
kBhVatGjU6Dn3kG8P9lSK1rHPEi/FSM0JABDaVHRhNGy9w+TrFv0zNDbZatwAZGN7tdJ5ISagoYJ
BZHhiLm9xQkpSzPt7v4En1+LINFS882VgK7++9S/LF0l1uEQljTmzv0afEnk8YJqxV7n57hXRZkM
POFN8wy3mHsNvpDt7/OSjBkZMyrqYrPMcoaE+VXHNnJB827by9UXCZhEwrz8mwVlgpGvSX7vGzLp
tCOoIaaCTpmxTmHgGyUi3DvBLly+rb2tMDL9SCZIVGGamk4Ed/FKEK2m+E0+WkG06kkG4VeFyGvY
wrwouoauqhmrJKirKQe4umEuHfaSDUYFkaDUlEeWuEux3cToXsgz/yvQB/ZK/5HWdT4H+e8ZtY26
J7Isa7Nhd/NoAhsZ06eDoW55sRNjIkkHpwJnEBBtxmi05kFlRyiivIBZutEWED41mTIb1ckHmyTp
Vu914EVXl+Urc70MHn2m4JGb/BwUBkelv0DEcf7vnXB/LmYzix1Skxw5HWwkf8W320MKo+jTBJdO
D1fNRdsLlGSQKK7lmxkAesaxXn0/ltWWZKc5Ax0RBG7bG4lptzbbv7IM+xGodOES9aIlcXmm1aNL
2hnssa4PKiHhAS5zkW6s5I7sW71z3yhiBkgY+qzh+tePyocOxZv/AuEdtz3SJ8KOZoG0XAmXaxi9
/5I8Pvf9Uk5SzMV9pIBWwa8teF1OVV/I+jpdpyXtcNeTxQSKRRrdu1bilOW0fL4wUHttmHIBKK9O
kH78tecL58gaSrtiDdeZpHDfwWlU8m5o8B/qoTF0mbciN4llDeqOtLc3dRVVzMBg+yB1IsUSuzzD
hKtzwHl37lLJvyQnvyO0J4giH6dniscZMH4tUM+HROgrqlneC6dmQ9H3YWPZueQdxv+dHKHj0m2d
R+nUhy1/7boeJ73zlaWrfMeg09PbG3sZjs1xuYyiCwu1+iEZmq7seewnangOzezAmHh6Rfaw/ftk
Aq0JwHORSbWbP+Lj1BTElZUaUAin7mt7EXMGFliGrplBz9UTemoJfxZfJmJyRFx9TerR6DgXf+Bh
vyyF3cpUSpCNqe6wCqCOlsG6Lwluy9MAel3FiaYcEtFzk1JC0afigXMUsYBSIXyAU4bT/vro7a7U
tsh4HsyfwJOCF/OA9w6v3FLPZ0kzDFkpPjic/sOwnvMrwA/wbu5g4bHCthhfUX5hx1OJ1IbrrEre
viGpjSn1NdS188YUMZPa+SZsyoWwWoKgWcQv+GF12yzsxYz/dXQvJHzXMK7gCE7w2tnkuHkhixQe
5mGwuAFx9KoMfMSU762zgrURhDtpyscV4wChpycXxC5FoBeaB1+yImJ1SY7y/1L9Y39rz/OKZ0c7
TPvkfRcMNaEiIzPQl9cgqsc5Ys0hoUkA9q7A/S0d1OYyN4QJbChdrQS5bQwEMsGQw0DBrp1PBey8
FdjLr5fKiCc1IDK7DtG4h7PwJs0ElOtnoAid+Nismvi5AJz617BhFk7trIIyvfZr7OKjAGtBz+xh
m5EqvEAJEMnKAPGkcuv1V5/8N4EXSbAO36f9/FAv/pbyOI4PRB4t+DT29Y8SCMbp8+gjuRZFJVrf
Z5B6ta0yqmCl8ThAhV1djpIvobFwfW1r9SsNWg/+ySo9lJJQnz9SWLnqru1NgWupQ8AEFfJoPYyp
MAXjWVLgQ16OFcZ0Po/BBPCgpbyEvUhrLOahekRHybV6GoP1Tg+wwFlWtdGbilJzQtH48JZkwyZK
nnkfydIVKAmqsddLCSLHt84HYZqhFrbkf6aEE7xouef1V2ePZA4v01Ugr+qY6oxCzffptdoXzFvu
O2sv+RWfi49QVFskLBSp7wcHg5XkDMd6+SWkHY33QprimvLOOQTnK9IjM6R/jOq8xnwJJ2xx7O9U
z9Ykf6MwhigIb/Dcbi8pbc9sLCi/YW9+Z+IXv7I1ClcH1qXbysfIt5NanUuDvVoEc4EcagM6oLO1
f5u2uBlvrv14AA02R2A/digaBr2LNE7Voz+eQP+I03b+ZgDf2cMBAZOaiA3zReINQD1jaifBve61
tQBYJzen7RO9wfn4ck5YuhX2zbzRBqo3csAc5YPcOtE9PtGes2ziPrHYKgHY2zpavDf4D90BhXIQ
kOn0QuaWG/ZSLmaZGfRKDZASrtfJ4pjwGxpwTHlyQt4vkozE73SeVyiivi9miRXhUwGZ88t4lad/
2dpM8fBQX9SE8eSYrqz+PrlY1yQ1PArp+ef7DcUMQfrPF+Tei1qYwJfnZFuVA8ySq8w3OVE6Jn9i
xpVXzH+fwNj9nqF7NglfUEBsgKwYEiDtdZSjaWYYrAPawNMwzWu1GLhYOC3TaPW7O09zfU1R5J5i
pJaJdNpkcTmbucycuVpWu91qUlYC85nrQw7Ve9UEJBLQY3eO8ILZbp4XsJQjUUao6VrRlXRoDqeS
m/+BDcCFKLiUsrPzr86ypJVgbBkkM/sshBSKoCJhz1EBod/QSieahMk7ToibWqyL4dVUuixjGECA
g0AjXm5R0YcYkAGLKk0NlqWEXyue06WTv8lGhHYTH0heJv4PhUjEjI7jlRzgeSsLhce5DiGKjarx
acUk5M+hYSxewkpgvQSRAie/8sOclNbN0bhF76lnU5HpW6sOf/v5WY7iKhC+L7Sz3DzvcKpiGPuf
18ndewV4QQjKU2O4Q6A72XkZgWw8jCcPMMEDSw9W4P4G0X0Q2H4LLAq079+oZpqQxivH64XgGUXa
g/XTu1t2gNTIAk4LNheOc/73zUIPzgY9ln4/vBuxKRtEVl1p2VINridiniXTPWbKPLF+HC4O6hSa
j8Ezt/iyXkRgnFiufBmW6iCqM5qYwim2QLHHJafFrKy92/gHwpGvEcmCyXcmwOPXOZOEVbSrohk3
Hai9g2dB8BUp2CQHeTPuD4cvgWLzGSR4FxDmfwPafvba5Oy/DwbvMJo+p6M2wOCAFrK7mo/MKjMP
Yt8INOOPTmgac7j/eFauYGu5DRr+PokrV58V1mIQfHnG+JgE0uZ9Bf9hEYsdCqJIuhVt4UIIf2no
TKbiL/xGWz+EyPuc4YMndQAy5KmRhSH3eFG9B+0h/VXQIMR4cvOcLa/wHrL5KU7jn8hauZQQUMjY
NQZqu/sTMWJIRnkpF8hrk+W/eC6msaJu7G7TMHzyn+fEzJwLZCjzCjVxGthr2l4HlX/M6OYCQORq
ZK6zEha05LFt6d4x7XuvXLnvueWIR9fqyv+p/HJOnHMRaeMtHbx+7DBh9/wFG9iXmfW0sb7KG5T5
HLb53XtyIVcwuPkSqiSr8O+uhswqr7HjZBTKJLeMvUaTKqoSBzgD82eipxkYsRVU2hwdtmxaYwE2
yIepcNhQRpodCBx0LgyQJ3m+Hlk/aIaosobZQmW7DzxMyb7gB4UyIItJVtPNoFYiZjfBQ2Ix2fzO
uLHFbYb02GcF6MvS5gOC3weuOmCaLAwTKBGmmx9K0VfATJdJElooAFsRjtZ5TWgNg6fj3dG8mySl
r8ZaGY6bevliO4+mNvenO2HU2eCoSfcWNzUpmLP5pgwOqfT1h0dJbLyWtzcpv6G7fFO+kLhwyUBd
u8tEw3sSQ3XmZrbY6nqW7Cxm9xT+aa3wlDszxMQG3bPKLby/MeY/VRMdDXzpqaIs4D1f21ntFiIq
611/lzJ0XxVsrPhtXOAf51Imwik0fnA8xVql7MrGCJgQdf0+rdUoG6nbc1lxZpuPeclwqdjIEZRh
C7I4ziEt8+CWBE+zNrC0848DGaFEGmT2P5Gvaq1MPIcsn8VSq2DhW/JF9kWv5AacI2g6avlk8x8f
+j3xouiMaebzBAbYqIDxUJMTa9Dph0pSZZsMlMlrNYQyv7sJdqVNT1D2PVguBMJngXELp8o0rxQH
8rSiMuKS0HNEQUeXaldf8c1qsMB1/Sc/Mw+oiMhsUCppI0ncYv7Z4yPoCcKSWjVxLofI9c/TBOt0
xToMo1qwMnvE/XvH2cvvyu4BvjxV9WvTKZiupnM5tEBcwwpJQyT5YXQglebg3MQbL4SwmzQ9YnCE
rPYK33ZdTfchdVTeQWJgwNCLrwXpW5vOwmx+SjW0hEm4vZ51EM4gcRWijZC6Z3lKw76yGmOlY2e3
cnAaEbOQ8AKu9wun4zzRANPBmqfsbCiGJNePzh1irtLh6bWDCb+xUpHsJYjqTZRnhhbhpCwmtWTz
/dVuWy48pRnU+/xAVzI5dCfRaAwDsncPSSqhHkqlwqHSqeH1DFfKJtiV2oYlLbsrLgPuF7goliu7
jPIZ6AgJ+/83pgoMbHXKNeHor4maZgDfm+nRhD39Wn1SCP52eebOZCLvfty2foTGsOeKy9U4GuQ0
yZ7lmB2y5LFk5Iu/asGqjRrMQD1XfhPFzBWRk3lyO/x7YhmvrF0dOOF3Kul1CQX554z24sLqzoz0
sOFRSr+tm8AzRDlHv1r3EaxxO+DqDV2dxnUGRxJ5CrNhsjap69uMu1kIiy5TJrJM251cbQXr5LJz
PsuNjyGgyn+SRwZBTN8mh/giotx5/RqHisrThvcgxbIVH4Bn9fvgr+GVgmGYFjSMBD1E4pMUszKH
3XOUspqlLVfAvlhAIRrat8z5Y4d5oIKCKjYVtyqN/1jiNmD8gxuaYTumGp1+8OZVU+/F+U4E2PyG
oDo9EkSuxExEZtfJTJm3emBrIJNsEw7XWT/OIvAnykaRqUEE7SREZDEEzA02IOJkDto6KVAjFwFR
IvAy7ot9ORYEcWuzD/lcVO8k96xk/EKHtg5UZnKFs7x1Rt3zK7fEXGijp8SmWJeZMprVK+gZhaSQ
l7dYw5M6AwNvGAaYVCfK0fwUkmpgOK7GWFwTC9CMtYvux50551/jK5UjoeDdoUDBtAAuWug2iscQ
ax09sk/1B7fExRra9+/ljnZMfHW347si/yBgbmyyOPj84SuWgYLNUNTWAbYPAQIiYXTC5yMt5P2u
wmeP8wZbgd9vZ53wsS7qjuvWwzvg3l/XUF7xyK6cuUgUK/aIZBPHIyKBmedrUnx7JjaIsNa2Boht
f2YQc3nwxoOqU4ySC3+srYSyTHpuDPxDbN7Bs0hmaLuYiMvoUVk/zWgZdE++T+gJ8a3Zroi/kJAp
DYRperGKl4S8Q3Enqc0ZqtQrCmWTAm3Qrlk5uxiZMrs4hBKLY6uqsN4KeWvSzGqMNhS/vqXQy8um
7Q5VjVztY+L/RzHBvGq76fVkDJ2hGrFUB9u1eKXDwMgqiyNodHZv3N3q0fysbQERVDjmqvyXksdK
G6z7eUGAwlv7CB1xg8z6aiJ3xL/ufO8raxsNHa8Mi/rylHNEeMBQEwOQefKyvck51aoAkeV8kMyD
WKXgKVJTPNGnejD9/IpvqIQWUDEdygCYYaoLPX6NSIMcbtMIq4MgxgNcCptSBoadgZQsJKEktsGa
uOJkaagVnMW6DjC2nIUhrcJNIt9mFJcpZJktIQMFXJiZyC/3V3YRviQEkQ+feWnk/Qsh+TumY7Ae
J4fxmbKN2aPqD0QblJCbOLIaXKRfKOMKiaqso/cRTWoqXBeHOrHmbLR1E/GDO/AqvoysHdrT9CgI
hXxP+l9lC7s4OCQTjPI/yG//HHaQI9Vqs6Xlz3viRJNBaxule6Y6bbBJV/hq89WJ1ddY7WZMRX9S
464UlJ6vDXlqydnpY5/O4WvU5pQXidf+gAXryFxPp4R1X7SR33mT7MF31Ha8BuhEc3CyfIA3iL20
7p6TSoA7mTsjqZuQN4eosT7DQcuO/+n+tcvcWErfujuF0Pkeo2SgZze2l/rPXREeVW2BOVQ4jmOQ
REPQGvMYVCgERLSVm175a60DhsN0ytnBP1qWwzy2DwqsgvLRw1OX98z0ViAr072x/C/+ifFbVqnh
0e8iZOlzZss+J5IX6oppUllKl6Jf3Tt/68biD3FOYWo48Q3djiJ9S+t7F7W7JcEpxXidMHDPK2pB
GSnKLJbiwaXnk8Zqqp2CBETY+37AhQvkm+amEvZ4t5goI44SDBoPX/sQcLBxNJCyD3eU70o2FrLU
Ecya/qvjRZUffcREH0UssaiHWJpecn8tHDHR4esT1K27ao1ZvHMzFT8d3rPywYskrY1yhZWWGnrj
OHfUGyHrohWHL8BZE127AL1hcD2MMMB358Cae0VMMDMCHeftCBTko6HrVQs+Xi2SEI1fUSBiflAx
f+carvFqoFb54YUbjRrP9y0rOaOCsQcvi1MGPnB9ljdtf18l6TKaW+xfiPQwHE+1dt6TnJOXaptL
bjdvsv3bYybZxPg8MsDOPWPxa+CXNoRJlOV0FItg9GTueTps/SyHB5bylPL+cKE6s5sQ68bAWCC4
c1lGxdrFMiVVcG86VPvKV47l9acyF3qb5porvpsNkIMpdi0x4+Chtv1zX0x5/xvqgl6bTu/aYgPb
YaY6xPDI+B3NzcBiPjXkb1t7BRal64h78hv+O06JD2q0T63s1AMbAnjU7pFxXreRdyX7s5EQYPs7
vrVhFwhWdyiI1bhH7IoTdYTIJ2snqU/xBKwpSSi4wiuGHntbmYtzweRvBfybOtVnmM6MT1OtinTO
12ZjjAUqV2vA5frImZQ3w+zvztACCglZP3/fTXOa9W1p+l0G2CwZNjsjGVhg0GFoOubkvlSJr7Yw
5InBFS/RzT6+MPiYfynjVEFO1ZDprlAV4dQX63T77MxNkCA3Flmw99xSDpc3XcBuWl1BaoKLLPqr
BlkgarJQjeCIydgiyutEXIApdIMW+m6SIzlyxkFXKjR8buQDCQV5uPlH5Oe6Tqa6c13Pjt1Y+z+P
OXBAB0ljuWX+fssz5wmr43BmNo78s1ThndpcdSA3UwJ1SOaAwqF5TvhIbhu8cDHK/XADy0JwB9lA
JC6PD3mcSwhrSz8JwCDZ7YOW+LiWVVXVh0NgHrzp7wfvO6HaZN5g6Ws9fXvaIf6j9Vb2SgTKGFRL
+shMCZIGuq8ulYwvMxJrGH4J2Kt+JHh1aKnANxNdM+CLmrRR+9tUQQbTUicOdNr6SA60p9wnKt0L
vJqy65hYpSqj1eaaqwBdFbKOHZuKNJfvKRESV4KQZnqJiE2fEj2qylHA1AIBEwRIJVxSZrSZPeiW
60qe7tvOcndhg4+5+BPjxZuwPRzNPbsKjJu0mnMwKxaiEVHb7mX5WNMLzZ3rFRACDyTwxwiUFdPa
XmNppyBU4yr/04lLphQi92IW1GJHSI7+YQqGPPM/klFzk0326b3CkekhpQWJwlRTdNvJPxRDd0fi
9Qsjc+yKeECxzZWeV0+jU/CU5tMA1euTeJxxjemCWsuAxQaB3NdeMW+dWdVBbqZx970f02NB8T1B
ZGk3qhDygsD0MNtrfai5KR1c5mgLVZsSr7eQP24HZE8cM68S464jPqqvLJnjAVLskqzqhd4SUlwE
jiwqbkz6ETq0izeeU+W3klEoW5N7W6Fo4Yqi+uYJMGTcDN1Q8p7qSQwQXzXu4fm6fAaxNJ4ATpAC
CtzRgHQ4lgjmq0SmAk6CcY5p7KqEylIf/mArEMMikNOcgn1JcCReFkvKv3bDFdxCAbZmbU9/CXiA
+2uw+eNnW4N2kF1wnBANFxXcF2T3J0Br+V7DpTesL2uxyZ52cpO5N37vXhLQEGbjpozO0PIlhABs
NjxfQGFFyI+QMBmTXmpF5klYOVsOZ/kJ9Lc7i5spKU8ErZvOb67MmM3HWtz2Z7ZcNy8Ahk0IQlpq
0Jlv3pkH7mhs22e3V5pcTrHggYBe2qiSVkj45qUyUSGmlHewtm8JQYt+m/fWMiJIYKInn6mY6qs/
4v5x4VOt1zbKgpyUzo3drM52LDy+trsxap/4lDLyVq7wuNJkLc3C9+LA8NQVe/Gm7j9YzOib0gXJ
Oqn+ykuvVyhp3RQ20JVNfrC5fMIfZsr9gNDpKfj55s6k4TMRkrbNUKW1P9AdDI6XzQ3PUzg70WF9
Wz2lllkJ1WtlG3SzcAupuEb25mlOQX3QEWiFXKq5mmbk6KKOkpGDzbLBnX3zJTEuXz+Ky7bS4tsL
KbCQogSM4p6iCWxoGEU48RE4dX3ux5aOLe1DUEHWgpGrX5mlTcWQ+8aNssBbXcBIC6F3MA+mw2/z
ycxEEC74hvmbGSD53j+51zDpEJYHjx3yTJjcb/46YAbA39Hezrb4PXocQtjaj+X+i8v3Zat2EL22
DXA3VSBW1UjaIQ72utNl81hmfuNgmghqn7rIXecyFPfJ9vIgQ6ZM4Egi/0NqInpfr/M5CSqwzFRE
K1z+AnZhTaIvjgnngsffwkqpDiqs7uTiIum1Ox8UVHq/VDpxnfWNLaXe0kZH9IRVqsy3Ntfgsd1I
sKPhcjXc9Mnqf5BNE/n+wJ/i9RC+xqITrlNfvPs6NuM9RyALw0OlDZkDM9zBbnAqF/emFkNYoutK
XOfIZcYkzLGLHM2R8+zWEne3bN3yBFsfV59f0tgggmrpmgms+zOqqWJW/C64vYhkLFQtUhd0AeaC
DBgik2sOE4seRn95fT1WusRsgmvQjyoY++Gc0cLcJAR81mGxdBOV53RAk71fVBk8Ir5+J8uGJadZ
EW0x4nDbQOMNc8P5cY5gLZuVnaPHCuV0zqGcPG9RsATdxgr9bv+msBMd5MQfM+otM+H1ZQwHx2x9
HnMJ+zs8B/WDDfitwC1ZR1Gt6uTOudAppRgq0AEUtQA0q/kMLGn75PMQ/ajSX/dgtajnjDIXeVYN
ZYWkTAfEMsHDW+GMP6T4nPZIda4TCPomJq+pJw/Uxt8BtFxRE9R2JHyUw5XMklcMxBGUhDezxNMu
lMqTzTKwR8MLgF99JXnndTyu8ikMefATQp0J30jv5096yRqxKZDI9mlppJ3OgIh4nLVwLqId+81E
EyaNkd8qXp8BNRQq9sCXk978RRO1nr5sP7HRF+IyZon44KGE5U0KngX1uCCd1l19fHsauEhgD9Bx
a+mahByTLv2MWLDogsECgPHcKWe9meFClVlX/USgeKShJUkaJspL6VDSOGA9bOdVtk0L2Ch1MAQN
lSZlBxBOuIE/xUwS1EM39eO7NfyTXrvjGiPSFhSGrpEebXamf3h3yjTWgqlnjJFLPPrwfKLwrFp1
JpxKT2S/rKnU/QcZAObkeAguURI3UZXU8owgsHjViXcMIQc3BN/1WLgSn4XFAdfSQaPiBOl2829P
ErmSgtFbMWqodEYTpEAkVXBFPRScDm7Nr9jg40cKTb9iShXQUOBLn9r00DYKCVyeH9md8OIrN5an
goQFJszzZJOuqALVNv0ze/ns4PKr+Snqa9A7eOy8GEUYxg0bNoK9qHQ0/Cri3ku3A6di+oBr/8Bw
X2dsXXzDbfpsThk5cm2J/f97OU+L7ynp2kdPoiYi7uZTFvFTfZnqgoxD+zQ3sX8p+CHZk64wx5Ix
Mgu7BYzLCRewKDtrNvwrbAkfh0/XtjvV0ovD3HDhURxUVH64Gd4Nq6lcfg3dShUTDECAGjQJkpFx
VtXCvkIxFtE5wO3PnKFapqtUdxwyhpFeY2pt/jwsSSPI54NKA2i0q05RwqLlrQ2U+mZhz/lvH6n5
s3KCkCMbkqjHVdOW1PnjG9s8NHXwl4UXfqsrojpWoIxt7khI2ekelSwzIFEw9wEC5HoOWmUPPSfB
0A3y0YJVO3JjVIbwgI59pWClpiN4+SqDH9n6QHt62faHgbRPyfBKWJVs1U4RypMWZjNr8SRk0nX9
0Vpjt8+AE4D8cUBZmqCc7FQhHkOveWFheuX6F/eAYPJLjRnJPyLioECDxoxaBAaaoqv8gyFsAXgb
1CX5gEMq1uJbsNMWIjrzCI7MMqKOA5YDqmCmYpjSC/2SNc/I41Dp5lo/FIdL0USkop3LvFQKg7w+
0H+Npi95i/PiDIrQL5/h9rb8L/faYDT2OtsIvVUqLJcoYjy0k+Pd2oHxk5VJDwzxTTUvVqtqaclF
8qEBTcPXCdmpP2jDo4O9gt4/oST89rXLqzogCRSUaW0H2vk4rvz1/1Whg8WNOh6ChrUzuxvfA3xC
MOqzikD22moV8cZLWORvNRlL7Poht10GfFAlj7sWZ133Y/ePXoDiFqy0EWqnM1iB6/f/MyLCPWpe
1CjjFi0ypjxhWpS8mvGR4FHtUfyEBcq+mj3q6eppx1O8rjPYqyFybwFPtSnf0O1bJek1AsmCu0hh
5TirzbMFmi58O+kxwcqSLEPaZ+0bBPb9NGEWW0KJabdMzFzQNQRaRnjTX1CLlPdhgTR56dU0Ws0S
GTdIj6qsEfXp1EWsbYzLfkVwHt7LDeYQQ+dcy1qnXFDyyhQyIlhAIKEkL+zsGTvb+bd5E66bAIr3
v++TvmjnLf9kR9+cMmUfYMMbQm8pcARds8uHb4CCA81Q0DWhWFJRj6AnWjzf6zuSMpffIEYKXY+1
++ZHRho1f3B2uSeTs6+sG8++UrfGaw6wdr0q5wwQMZEs3SoY8jpoWDIHQbzqm1U/Y6eB031I/dyI
5KNk9iKhv4y9DDbrz86qlMx2CO5oxlf2nfuXzrBl4Thu6Ct96vgJybgHQhGptc6dVOIu+hRX4rim
2uPp+llIgVmvH3jRX6ETO3YNmTo8m0qvltx5TARr95uW5X92zefboOpqzZxsikB6rzypfPHIaQxN
VCCIv6FiV6yrHTmLgIkViwGtH2AN5S8WQN2dAk0IxI2WLEDtJ6S4yF/4x+076rE6oWwoJVswT0u7
Zoh8e9fRt30i1nVCx5FDXihAGcrAaxOGAQljXyZ/259ve+ZPyFyfd2Dks9AJgswYar3xjPRuwMj4
srjh/hgYdPaA8g9K5QtC1SCkB88Tb1ZD8BqXy41w24FRacURyquo5tyBY+ruPQHsPvrSDzhXWlJk
FCi9HSw9RJJ+i4xn9sXH16VQq2KzeZ5AT/WlWf2DdB/QfJKf+wZcJOp9FoQTyJYpw5s/JYhcBr5O
TMRBBLwM0zHneZnaEbRKgVREIPlPj0EBKcbYSJmHatllaI+aCFHso/5mKPMrDiDYEvzpQAzzBO9j
A0GclgfOCslaqYZgUZWa1vDJfLLWLc7C8/VTB/h5ZuqIZXbuzi3LpKmfl4rwFN6VryBiHQ7GKyU/
rro6/bWtjMmdJ/w6fJ5584T1H7qWz7eoPM8gy8PsqKahVNL4canyqpgqyfLYbSKICmFEcCSJxOiO
Bpdov0JehiYwCGRvoTRCoj7OAgKqxiTG3fpRZXe+MtsEmiPkHiBxv8xIGfqpH0GT58lB2EUx9gJh
AGuqiKucRLHZ2p23uB8+kuv1sZyUkNewptzDL4egWBQ+hdoTxCcs5pAfhnTnI32A050o7Z4JPT3W
qGWvKIHxLXCizgEFzfd6lwTkRZ6wb9ii4CHsyaOJ3IjziNBAKETLrG75nTM5h2QNDQmJO/q+D64v
AxKO2XGkUODT3StATx1AUdBATCbAnWGu5TgQXnyprJckEU58BUxdyaCrCu4S/vc+uQQ2P1MYVpqZ
BNfafKe8vPeKhOw/4kPlhS9goUKHcOVqZ+lt93lbd138z71tsHjWMaTNxrJisW4+gFff8vlg/2NN
MjIZMNQL2uUPY89SkeIHicz3edc+Y3blOunURui+xKKCrPA9xO9Zf1PqZM+1XDWB0zDsSHinjl/y
gCZAvYKaHaEvTq1fJlx/nVQ26G2VS3yKA85Swt7bTEAUw6k7sixIiwkACuATzkPiQUjZgCntLY6B
04YF7PQYT8LZ2mYAusQz8FbJ4SYC+rG4oRzlFQbb57on5O+pnL0Ss5E22CLNBz7acyPFf9y+WbYz
KKwquon06Zu+/2w/9N4+RiFGk3hVV6pY2KHbr2KkRf/cP9Gf5LRerw6R2y6rJei3KT1bx6qAk3Dc
cXhp2BDVVh983W3hlFbuXLvRXwwkDIdQAFL7uX9e+2+M7kfLKo8ILU9EGrKabsjFJsEAg1LsKlCt
Qyi7LypR4XkdVs9CIYgu0aQyinA+xyl3aXXvFzthjnvRHUZI6lFl386pq3Cbaw0iG9YMNLFKjb/w
l6IhQGJfV+KzZOjSyxylrqscdXSA+GVMdxuMBI5bWcr6B53lNfhygFaPEAsWVpXB8IcNa+de8eGZ
234jxA5ncSGWsp9kHN14TaCY8AIinI/pPpgj7g9497hxFrAgH6bX92a7rBis+iv/CqYLvz/ARm+h
aCTZvQx3AN9XrFw55P3gpQUYiJtz9pXgpFNQRfdwnj7EaKrBPyqAJw0z52ySIi1beenusBfIkdZK
fKlhK0AZJq2eXAibTyqnBNARuc5jtjGlCqBcSqvHtfzJ/4Klh1J8+1pmymeSIU9Z2oUaAG0Qp+ki
vegmLzk3rfbsZjb3TVOtN16zskbXWidqellv4LUFQk7m32GR0d3Au8zBscnMOkwpNDFBYK7NzY+v
qSsKRL4BcGqI2ZWbRxFOsUXwWmyujdi9z/gezGTwdtGkz78OPdoSSq9IK9pVd3pWtF+ymsaaG71z
ajsZmQqh3wtnv1I5wiijTCvteu/XDZJB26jOOWaNyl5O+g1eURGcF30nz+ubnaoGjfQSdvFrLU41
ZBjkYUgLZXCEQIa61JleTvUUdq2dvD0hV5kOTd3F6I8LV7H7P25gE31pCpeEmaWi58n//tancteg
q9LYZUAGG3iuJDg2Elb84+CCbcij4aRhk1h85RROaFIukbs1A93ACPmePpxxaZYZKNn7iYv8d4jQ
Ilaq+4pJfOdYx+/qH40hlX+SJkK0NBvf5k58oitTcXZSQMSWYiqmdJcuUsYSs1PFG2TI2H2nptEM
+va72mMnByzzvhTvjW57uye5362SIO3ZTSbs+RvN/N44olelxZonxACWddz5iDOdRc+U3Rws+wS7
sjuf6kP2iSFvoP4Ns4rsRI/x+4R6fCXXzkkNSIdzzxderiWsZ/yJLsJW54366nRE52n99866Bn2E
CzXDQ9GEYRmz0e+cbIf274DKB7on/hlJUPZiAPgbJXgq4dhG0Ekt/4NcdyLCqHY1EjOi1W5kSnh3
Ygog8wd/ccFayILntr0PPFkKcElXT2fxPFK73InnK9VU45W0CUFAGqpSAefEvo4PWGuJomi+Nu9c
99YBCqYoRTScBmmFE1avWhoEz62q3vkRpnufiNbtQQq3lKT7WdG+JYcUgRkzYxULYGGVWeRxwl7k
uO5sWvuICSblYx6+RrB6nbxGM/pKYPyWwKVcGYkwBZnFI0HDun35oLrm6UZjNmTq2N4dOOZ1GZTr
thssfU4Kq1StX30nwMhRjhRt1RYLOOkLyn93M79um9FIqv4s4f16C6XdnQVc/1mstSdoupvzM2aY
Fp5tzr3V3gJfyLnzOYoqyGhOcnGT0BgInm9Qr3p4ZGfqR6HEq/7Whky2Msu4XqD3uTTMYVxHAMM7
YvexBs3It25XT8ErTfEQznngztEdx5xsYau8K4FmxLEXN8MJx0SwWIjbrxN7989QSR/VfJBSFiYK
acg6D474hZPAiJMREyzaNiM0a1YmZ296YgeN8uqZpHQiVOWFewcy79H6o7uJ89gJ2L9PX6jMof7A
cA9fjn0CWTZIlqeU/Mu82O1aD1p6iY+F25x0kwrcxVc9iHe0LERLZ6A66Aun6HteljmsX0oxELVL
S1hCcCrof7L+KvI2yZPHJbLy+PNWcoEWOmkrMeCG+5pSlGFZgJBEnntSnO2FeEa2/z+Rh0y5ElSv
oG+5vsC11ObUeglxiTPgORN+QJi9pYse8Q9gc7H3enoRFI8EazXRgFJbBLvBvL5c9ojveh//6FH+
2xif2sNVSQGowQ03e9+URWFR6hMl80ZFvMkMMDZfNTUQoeBD+SPNUJvlYvuVbmZzKiispQnKMSMN
aclWPbJnlIm2AbA074W+0n2TXR4dsfAJN391TeLDe6eet1s29nyguZxPPln1Q4Q+UrPrO+Q/JAhQ
VojmIqBGC3gmCMeDb0U7fcL1qT6l5ELEEmjwCK0VV26N1wQKP5RyuDIPTDta0HXpJ5SYo9OuDv3/
9GU8G3VwPh+uUiHbYlfvcKY/0dIGSKho/76eC9UC5jY9XZtQ06jMX4zgaqXSVk/kOH8/X1kskP4d
d5R9llLt0NnmcyMfdaaV6MMnkGJHjf7s4tJR+LEtJSQ3ZJVX1D2MRVVev6AYeQYZj41HzbIkVkVO
kFMwcQ7jUlPyQTDcBM/Syo/ZuBCZMAXmD3lJ4ZEOYuMc3aI/Mh8//d5Cxn5WxfZ3ufZczCe+R+QX
H22t60GdPqCleP6LHqYi1eR5TKtqdnDwdcxI7dqTd4prD5SI8CxT7KZml3i0PwUrJBnOMY9s4FH1
sZw64WLnHIoQ3e6myg/20Yk7ifoZyxRIswzrNp/48vy3OMC2JuWOSSQr67LxSWZy/zXMt8uSxwtS
oYcq9PQOLnBmHJGCT4z5PD0vFfocpOfiFmakmcj9L+Pkog2s7n2N1j/QRrkgmm38exSFdUqqKtnU
m0QO7bEjzGPRsBPR4ZY8pxqqvyyoAwgkj6ys5va19EoECSrnRDkJnH6EloTBYckAwtrDw3CJXsKH
QeFsxiMFE0OjE6ctK8Rta20gyntLw7tcOsKrSb4hUMRGV2bqQbBtpvbwMN2i8cplTBj1RiuPth+G
kp7WJj7HpZetuW/vb9RtWBgCd6Ls92D/FbJcjiGpUz+jeaUgh2CdmKqEVs5my9ztO2O4I/9kBxk1
F4ppFuyQi0QvSi+HY72NrYqF1RN2vyAN196BLMfaxf9NRxzNs1KWzdsQIKGWFGqiBQm27o+ScPCu
JnlTswkrKbYM87Ly0NmqxwNXUWpZRs4Pt3N9le8Mg3lXDKoNNGax9a5kmOYw2zwKDfN+iZsryG5L
HsD5/VQkk/9o83kZ2ZtczlOs2rjEohXSmwF9kX0zbz/3moiB74JB/fK3oyt+ejUQOj/UtyGiLK9g
LT7vPUR20nnmCtW/2MdtVJ+Ayq6EU7eRr/Apn1RZqd/y5G2OSr91cm0GTORQXuhTFidy1+f6wsOm
nit5JdvBUclzaaJiVmH7CbhGGsSn4e7aKI8szbVAJwHika2siWE6LtBGgBl9AifhC0JCWHeDiEox
v8Y+l97AZJoIB3mM6NHh18gFK/p4PP0QPU5qm2tV6vmFzkGXWXqFnxBTOTPwdjHo//aJiyzDIWB6
SPYHfH6iwu/llfdUaUEpasybyScjfmyq7clTx830u3JbOmlQ+eXcSU+sodz72IqdtDcOc0YKzskJ
xaogJfgWh7bbgUOm3BLGwAbjptf+Inzjn2yLcLXwxkM3v/wC1eoQFDOlHRcETI9cTxZVxzB6sgXr
qWvQDsMnKBWEqsUkI1jt5ZkExjRgRgoc2zw7x3UQP6uc6WJ5Lp5pnA4KrxXyYiDHOzV5Navnzy1R
LQ3iItAQDU2dY0fOwx3yPBdbvUG/LXl0wytMgLF7SwDDgHwoYQv2z4pJvu1yfv5VL4KrvmgN4+fa
OdO0TTabb2BQGq6Bk+ma2Sn1HHa2TntMQ/d9dZjU86Nkdgbp5u1Nfz0mcHrr4UzQ8lZYsyxWTk/F
WxbgPBmD0DIKhZzmzoGPkwhNsn6/HhY/ih66kDbvnnGo/K7ogexs4tA2YvepYPOJoqTI0jG/CiVR
M6yHFvWgiGO/MIghY1lj2bDksMWqNtWRH4YNRSR2B7LP1aI1IGyp4BdnTnYxMmCXGqBc0y5l9gko
mFSsEdraxlt5Gy1vssiufzY3wijBxRwMpI4sHYEBTiBjgRSHXll1q2sTmOm2odOerA/zfpSS/XyN
eO2lDHj1v7i4d9Bxt1sRIxaNKWrn/BvJvl3bvkpJ2bD1BGitFZzs1VsGfWTVKvtWP7neEZM4556Z
+hVtbT1FG3fk9oCX4D+SjBrQRes8pSZI3ezZaBmoanhveHQnyVuZwOnZvWvf3yvvAD80k0aRxgFe
M4viugOf0SSveoVO4vTKN6vYKztUDejoJYLl6gnvoDY8x4gm6Ju3syymRTU6lSuhoRkdFWveV87l
v6IZdBDyfawgIjT4Af7zw8BggFNqpvZbGepWyUPSD/EVnbPqxN0IoFTwpWLhhe4xPykA5c4x4jh1
X4mt9swHH02fY17Lv+lKRe0atrwvJl5FZwfLmPymBXVf0gla6kXwzQnes57rV1CtbZBom1itc1Yj
ps3eJUISfLw+sYFcGXVVJTOjN5q1HwZSrK6a3FOd7LfYgSmcGw3Y07VeP0Wh3Mr/OrBQpAh/7EQf
oiOXxiNJ7BWuDLN1e99aOYIkw65Pf5BCK8ug3AiHBkbnur1sXR+P9TWmGPY1KGjphv2cQ/KXZ1J8
sbHNTXVcE/nX2rnIExRSv08xIr8enQUp+9aPcDzbViBr3pUs4dJvxxJXj7lL2CyZsP7LYGR5oPJv
Zrg1XjQBfFqxX/WITMGn2X7QPXwVuCFV4d2ZNlBWy3VQHwxUgpB+vDjnget9wmS6jYFNlXGEThVT
cpxVbWgZpGnOioZ+TsCi3WjxOm1u4vxP56gtmq2bXZE5wnB4vjF5IoHIhZKxNv9OjyrYhycSgpZb
K56rJwoo3xX7VqkBgnMj8GnH/gERWaW0TJM/aA1nUfATqYZIDSup+gw4c7TDt+Zze/HmfjkdRD+P
INzT8yKmpSDUdnHYs0sJe+oa8s3QVqF5xee84PqODk0Sy2bliJm2ebf30rYOhQXFyfR5EtZfRgCA
HSfDOcOpGTTDJlJMN91hX8qdYI50Q5M2lNmoTOgr1uhYXG8Kyq83PRclUmkvfKPDqBA6sT0oft4i
bgfWXhE3lMW1upiOhVf0a4L/8Su4qfner4k9MrLOBkUVp/v0UQ6GJX1sgHEtRliN0i8bPvqdzeT/
/FC2qW4nxB/rCYBxkryrCtiC/jBtoLX53hEHAj81iU6bV8WDv6sfOVLDRb+Hv/E1eTct1QQZt9ZJ
H9G9bXRfELSOmjGAx2HAXFMwhd6jFY5QuKqWqfXNCLXYFDLkA6O0ovLhZkNYjK1x8Al48eFjR+ge
5HjFSBSF7PsDPzLVgtCf+VeVVihy1uQ+uxhSPYDUQPAU4CyIQifGzt7gi+B6xXJxMa789/V3ZQxk
FrHzk2yHZKmqth4Pmv++aypfxusCDeWxDO75XEg5IQ+vGs7/d6SNzRvJ4oiy9mwj/rbKyn4/71Az
01C7++b7zxCUtSGSCzVqIk8Xf17Umf6VEYjy4RRIpgzUZwna/vTNw8p0axQgm6zKHP2I33GiXDwL
zeYb6HDF/Qp8+2xPR547zNq17BebjQnfIXFLZjvGetlm1dChXMhzJ3emZ2NFAWXrxHvr+uMsfsGN
zCjVlPdfjpRDpm8UOgBy5suS2gRHkBJ1DJx9TuXVseQTJxxgCSwepi9dFS2E5aH1vAH46dSebikC
cPwVUmRKt99NaXw69IhHm1TMdUtB9w1+DNrnKSG8aFlPrkdhfD/MZ0yiLoXrGUF6cN/rVGbHiy4G
+DXVejxZ1TTNnEI7Vj2VXiWIVn3Bbj/Tqs0iKBm9Drp1igW4datTcSLew2+1ZtHOgSoFcUyPwvrh
7vtr22H/KCCUefCumXWcXm+t1C7EA6/lgfmVBs34RtLrG+NnO/k0ppMp+ZNmnz7IHSB212XOEwKL
eDHbVgAi+ipZRBpk8puU9c8d21xug8zwX+DUOhg9nLIQKw4XpOloNfogFTLuQQO00mkKr9NMZTTx
DhA1pRJ3Ua/bUeHSty6oF1/87DEsWnMi2uKYk10fSGTGrUiBh/wUUwMpYBdnzESQMte1j+8s/HvC
NYDUM9AZJuJjN9z21/vS5jqIADuBZW4ZrfOySpTH/EHYxiiYigkl+z/3Qv7U3Lzc5+KY6wuhJSFf
6vND/7I/DpIACMP9ctF+3RzIEB+CNTAc7z4n/TtTdfC0pxvoBVg9NfS2BUcBkGGuEl/rqwSHPm5y
pDl/PzOq6esf9mfKIaw2OJw3gQNyuL0MaSfssJPF7ahk7/S3RqUpUqNX4OuKH+QKT8WOsn1fXGiP
O2fomweH1nN2fJbKr4WpC1ii4QND7vTWp9yF5JsiGlvSkIQodImyMm/KL4Ow9fbsohoKRQ02810H
H8VPMKFzLQcC3sGT7XOH5KH52lXsonoNTvaMUsv4uMOl9TJpKeN9ABt/Z1ZkzG76Q+hOqH1kJhIR
pumnQLQuMiKBsivjtLaAgKYrwojh684zeo+O04Eu6TDDonvcOijacFWsuCtCjWDRpjkHTNxyaY0g
Qdmm7i2Cxdtj1PKOAO1pWCNIOaj8xynmgqs1Y+vbR5Zv03J/+G8lcba7XOfA8DvthD2DDjXkxS3P
JWhZG31BpbNYkNLKWmeTQ+2X4Gns9GJXdfExLjdfMCbQcdS+1RLd9VLI3dGogjBKsXZAE02bBQhK
MlEvDSjl53ZBR0STcc799T0cVww0JIWamTH+050rJKwk5dJlACBx4jEmemBm/19o4DQoQKtgGQeM
voOg8cbyd+qbfGWYXAmhLwBJell9HGhqrMYSNstCTdc7sA3ubXHPsh5jj65OnzD5aD8clD2+x798
mV6pTigyrX/Ah3ddNL7Hq5KgOVXb7Zk59GYdNpQ9UabBFwMLFdJD0WUcDZw41u7A0rFy4/IONkV9
hhL2CfcMHRWODBACnqDJWNmSGWiBLbt+gr9FW+bHz/qZWyqprLAtJbKwdizqmKQb0FLQXLzejvNa
8YtNBVoDxKFZ6PuFaJdlLMiQYBTyE2SqcvzSMr+xKKHfWEy1yeRhrSrGGyWgxiFSBjICEDe58hyZ
EsLGK1ZFPtZ7+Dd6qCICFYkDoZNS4k2XocSzXidt5T431n7vXuQyojqPwuoWsufUM8hsVQdIc4A/
VYcUV/NSAAEFgz9AItyvfiorHtF6j1WudL3K7s8zkhrCeaK9TNb2GPKFTU2wIo9+Pq62r7B0lzAM
FXYYZuxSOxvXoFNMN2g/crHl5YGvawEOidiT0Rpg8qqQiqd+/YVyigJnbHSZgsDjYeyYbVduifW4
xuvCFL5iWRzzrubxdzWQlJB7kTgBKts0f4y4MdAqB9rlfiToXfp1ZoSa1XHswLs1CuSluFpCc0XF
m2fvf/OGA8OXTysIVL6egG21neLqDpoUkeD6U5M/Fy8KK5u49mbjYn38cP/ZfRfpw0ODU6DyzTa0
UYixigJw/Ii3/gPARsxaIW7XpDTqg76jMPPcWwsn+7c4yn1mM5wHzMhqKBnCFyqIjoYK4nJO877r
RQybOUqwyjUMcc48Ni8pQRRW6KWvxqd63mi6IvMBFSc1MiFIgk8N2k/U9nIVIR+hx5AZO7eVeRWd
VhUDXanZp8HeAncdQkylsIiWTWphUrJU88+uvQAY+5quVBsFlsrVDgAfV7v/5GRaEGZEpzBQVVCJ
7z0tvMyC04IkufvS4KUhlJ/NnQlyHJU1qtvF7SE4pwf7gjNLaS/kbwpusON9XrNom1eSeSkVLf6n
xvkyUilp4Wwu9mCfO9X5yWcyhaKtNsY6Jwh+t2eAV21bNLR1YpAgDMYJJZo2s34OM1si9lMPq0dj
Cy0rnqZDbWI9iN2HJjOlG1VP8n1ygGgdP6JhvUbUdLOjYA9b59htoP5VF1SwDlwIn5rGVQyGd2qR
bm1DhVrTCDqpuH9l+Dzdz8jclSL1eHCFap2p8Sn87PPxtQrOHueVI+L75Lwh+0RjX+99pv+xIia/
GEYDUJZky/fUlW2eSslOVTjJf2VwyreosLSTwbvFo0yfm34AwbLaLpEaMpetHYZjPetciKLqTE5c
GV4akAkXbK0U0JO8VE4hNfkkF59B7sfYznaROew0SosjOthByZN6EwL6RjGOFHdtNkmFenNIt4K+
QO0DcNPOklLiaawUb4HcG+uGZsr1U6GYZKrTc3H7lUGeixxg7j2Js60mZVjTH+v8WuYFoDz101aZ
wvHZ/vQQuZl508kZhdK3U5STt3t0u5lMYYhYgor0m0uYZaZyH2lgJuXC98cmCvb0BvFEaLtyP8KA
48GI/2zRhLFlQDeTEuuf6eS/HJyqazQp3mpSGdwlSP7mhgQC4VgKwS6pBhMNfCZ2FceYguijYs1e
8Z5kAAcMEuvFzigTe4h/gN8tgq7OfYUh0i8thyH2HBo1ahFnRl6lsYPtQokIKQKVS7os8F2Hz/3h
YWu4FzdyGA1HVHhX6NFaKYr3ysHjSfRetzaptcmAwmgWzTLhxJqMAuuwEZBiROpC2F9lrNUCwM81
J7NttT8vzvfpBXH+5ZAlGUSuKR6v+m1lWL5PeJgftJb6O/f5IGUVuUCph4Wq2YflIbZT/V4KRBez
jUkjIKFBsD7pKMRPyVb3sodFEXldnOu/Y+bIb3DVX0PvfxevO5wfOj9Ypkd4+3bg6VfzKXu6Wjry
vuisCWp6DMWaqKp56fDi9UbjGMSDYCALovmbqNUnr6ee/MJeLo8ONbvBG+4CARoOiXatxyMdcKeS
goY5fykUTuG9+go+kSZX323DJAQkz9qyhQs2nJ8QcKeX1tqU1WlCl3ydQRYsjZNwP/mCNd0D5Tl8
WIamE5ux7qumNr1OlUi+qF5f6sCq6zXZk1VVzvPLtDIkjLlPJCmOIytn2XwM9pFybfyGqkZxBjGv
vIoVb+um5Vm+iHcXMdkxghQKJzqWaLy5vx6Ay/iaXENf7hys86/A64vAnqwMl3l7b1kYE+DahKvD
EsxFaoYTiHcalR1cz9OST5ZAox1GHu2wdAvwWwb4Id4CAH07AyU8FvfZ5KqFmtnavqgYq25q6usY
6sKgKl71fMFoEVPAtBcReyo7n7k6n6DGN+SeQQg962PPaKzSFW1l30TUB29JGdZ3Tu05FJLxRSfR
/OCXDZjd6NuJvC1U+OIQLW88dhTO/TAlDDamiO/mXiJQxnNQ5tDg7kpnvxQHKxLrPcAxrDdMiOwN
C6F8hM+ugCwtVKOfCbY2npQoM4CK5MkIOJ/2ZzfQmlNqSD4+TIGa/qrMa5JZhLwG0nKsudetYXGm
bOXjHOeFeJyv46nqBLZyJIfYHC/Ec8j2TW9XLAC4CV2IMVcr9QZh0SSqANB3S6305yOhu+h5hsTe
8CoZ9GLsdq4eheVSZ6K4eRqd0BpxkhO7nmCYXBk4KvU3Wt6DTstuZumXDSmAJak0QTIWBwVaSdrh
PnpvWfJ0vKR3J0odL33SzxUN9lLX7NJw1bTlM391EaqCHYev1GYsqEdRcsMNQz9C0yDnYVg/RvGe
mrK1Yv5KUl1SNa+y4GKJXtZ/MTxuUMcIdhFPxEEjaRrLkTfn+JCuXRdWroUhO+52T+aTV2aEmPcV
BRxtR7K1E/p1H3OfL8m7z0jjiFc6dHsOzMaN52kcXJZstHosuIbXisq6yyN7cA6A3s3Qi3WN+AXy
d5hrD40P+Il5wQftXrzroJ2hotRt6BxNzvXuvs/AQ+/YvnjEP5bV7gqWRP3/7VlH4DesIhANXXNO
9EuCsern6oc8XoKt0JxoHIbhNngt0LOUnbHDc6zN9PJNY37VK/8eKiytASsH7B6AlmTbskndVGNI
npPVGdd6olJw804FZvd9gqoLytCqPyPWcgUOwrMjsCHONU79xOAKrNJslBaIWhv1fZBWAg5283kQ
e+VmTVigYWLFDM2XxTrHLFOnqJ+94aPSnsDRQIQrGeEyz140bpYZx+cisiVBz15Awjj/oMGUxtIf
vTyANbwXU+7BjyIJKjhHLcd2AlqPJXZ5bYzutAZhrvY4xELy+cfV/SQTedTcGkon8ouxOfY4+a21
HsAhAr1su572zNgB3P+dKEQ86saL1G15kyV0gOurEKptKR6eelSpRtaaiVhjcp3AD+ghNkWtjDIA
Gtcl2SWEBpXFwXpsNk4MNb/UhXbS65TbUwNG+m44y7tSG1pm9BRdEchH/z1pkjvB9DVTC/s7jxOY
A6Oq8n3LXRDKaBf3+yn83EATdEwjAv2HlcKXzwaSLnNOTqwGOCL0oiV0O+VuWndFCe2VGq8BJfKa
dbgNDaD/l0avqCnThQ1TYDhw7t+6ZHBlbpe6X7wtenuGx7qzcWtwGg2OyHJEBBvndE2qLp8WS0YH
olHF1LbGZjwuQ/JtgojYI5mxmcK3v0vab5g28OAJKJSmlbSq4KmM/M1qWcJrIq4Kzo5J7ON+XJWd
XpaiUTcfttr8uCzKsnGMP8MNRknoR9w9YV3XLA8lvu7vaqLxcec0R2dPV7d53NwYo/z0abOLBIXA
ihvSozLCTjl6PK/A5mh6uoVUPu+p/vraAkXt1nKavW55Bqk+l8cLR0gFJgTtZ3SgaLbzsOUccwJD
OXicvpwc8PyL7dsCvf2na462l2Nvt3XlKr+woSchbQbpSzv+tGuXrDQL5WSFLiQ9PddvDim1p6+2
Qym1wdtFoFC4c+vZRThNt04bUgJHphGZ7Sd9FVIMKxbMpv5A7Ug1EwghBw9EZWT2Nm//hZmukbEz
lDBVVjRZMKzBbouI8rKXQoS4oy9jib3ItZW7Ap+PISZSOMxT2XVeO43C1F7hhZRIRVmo9qmRizd6
FrYNxgeyxm3dINV/vm5qbtJsZx56bRQL4pVqEDlg7rRfi47Xc9IF7iMrHsDknxRXDBQ8Nm6nlMDI
+f5Yzib825gVhOICO35/CKP3jxo5K4s2FHk4+ZJ7zomqwAfI3ljpao0cx/FOBNTvvgudQFbDp5NQ
Mw6RBNRpqMzjftTRu0ytbU4/Isflp8QWaRDJ4EBWCLijvKWp+WcDeC1R0BOe53Fy+xUm4389aGA8
Obv2EUX+w3Le7ajaqK3dNmkik3/PfZ6h5udD+2i58JsWrvvyu5e4aXNwDXDkvKkzJPpjpMa/sBCl
5Rk+vMTQ+g7jtWUnSJcQHFORLHLMrXI/J/h9zx9KUmggSznl2+Kqj8zJkoQ52Lqy3EpSydjGRQ+/
T6GPsSWNS7haF7VyJf7jhIMgTtYn26E2L2IlwTG50jt9zFmvzYLiYM+7P9VEseAdvmsjDpv9ZF6b
1GOe7gm4G1WaCHJydZs0HEPl2CZkU5kXuz5eE7/UFN+UCPeUPKhd4jBJL64p72iRh+qRoNto2Ckt
TzDCBP+QuWgjeGZ3m+qkzILdBuVNN9NzZMXTsd5hzwsO4MMmP/CX+8Acs2KdEVtMKdSQbJEBFfMJ
Cwb0JmwFDCvAbKga2AWTOKDjlSoQl11FnAldnR4I5fC7VuSPX2/V+QWIfo+Ziz9cClfeNCfFI/iD
7+Hxz7Ds9pHZ9ix15OqdXPdLw8ywRIySLetpN95avmpl7DzNzaMH4S9jXyiMfBDs1dkTk7eedSn/
vbfs9HOuEN27uY4WLPvhpPpgmbcOmt/Ks9twkiyUX0AQcdumBFbVQp66OhkAZ/sdDcdOH6zIW0NI
4SK01gRsy9ZqAz0rK9gX9Eo0DKTNBm4pNhq6hQeTJSjksEd+xtACAvs7CunmRgrZrRK8hIaQNOOW
DnDGxAZ+HIH4EQ59m2PPqdHIcaZ3zCXyp58Rr1NVYELZ5aoNEpbUxxZtourMNIqH+tlmQUXuYmvo
OoGdAnvLzL6wYIBzYmOxrq3ATkihOml8LqRZBGdz62+3ULaWDeSmZLBF3NOcariCye6z3Sv3XySj
yG+28QsvhKDm5TN5D3xVVXeByoMVkad1u2ZLBNVAJA7aqVn4GNnHakE71MIOW4pLxVjoPMCq83t6
46GVB0nmVNadeRqzd2PoHrBYT9Wr9tUL1V5SmTadElDeWejY6AFdVt3rhKfThGYXCmzNAdIxoGe8
RjBHtnOkQijBRIIZF2eSfne905LnrJcPKshzeHQ77yXr/3goxQeJrKl/j9ogC7JSiROhX0NBwIsB
KSoXJPoQcPDh1Jo68jtTclsVOlodw7ST93RFymNaN9FcbQY2Gb/wtwwEMnM8zEwEpeZfJvPxqcQF
tVoF2snMtB/1hv+iE6OkHKndVW7yo0G47jgeovslTGho50q64CuTUoteR4O5p0Ery2pISS2kWP/m
R0wMavxqBByfBPPtW/kKe5gHYP7HECWlxU/yFJq7Lyp1rQtRfJ+Hw82sUNGSvaepkEiDoWwWYbry
q8WlWWQh8G/dXteFLGlb8dYNdaOGo2UYQJa4x8S95X4ntKK/xlgAn5lLvvXOvt5P5655k1epV1Wt
kz5mcfyZPh4bn+BtauOZ3hZdqLrjmXM+4vd5gjiphdQOS+xXhI/LNu4ReIyxQFtFH7dWYV/dsEje
4/9c+jS8NZwy4+Coq6ooOws4zDvZ07U/wda99niMrj5PsPtzfYYpRCHTTJVlpZnFE74mG6gRgnvO
MyXSoSqSHhva4ezAP7ucfbMREK1nDzCWctAsuW0/iqrWkPOYH8P0WbFxr0UcpTV71GlzPtBtMV8P
ZbeR2zQohnzKoQrP1EDyZCI/H0AeWhpSyArO66ccnf2MWdvPEKn9FTrXx8mO3Rm9I9IwY8hyumMS
FhSbEXDa1ibBORx0EtDq2PioxCpioZIA/WdTqB7/oltFPFry0EFc0vSo9vxxi5NExGkABrPLxLii
KEpzgqmCVyVceExXmP8Qyl6YqYh4Fr+NchlPpUBwVMSjoy+dEpZ9g7MG37Be1txqMEz8GFrDwCF1
JlkeKuuTNWdMJGnvej0zC4K6kOWjugW69B3jL4Z7kQGeVPJ5TELVyaJRuIOXFvQm8FYWtVAUlWGc
sd4CXDtOy8Ar/D5YAYokWp4GQ4sajzKz2uQMZyzt9iPATt11P/1xfJcqAMU8Q7CWYPCXjszrC2jr
S71yD/LZEKd5Tn7Nr9JL5NcNMc4888Kv+B2iAuXFhCM9P6nrG+uRmVG/dCy+Y+6ASZybZctBEQTO
ji/ujkNLzt1/LoCvhLTx5yrkVSERNHWcjqHK+Hfua+LKs406NgMaZeuxw1PnJnZh6EwrjSSGW5u9
NBqiHPMuA/yl5pp6Z3Igx+nT9vHuLzFphrL6KL2Yu6ZV5rF0QulO3+6OOJTeQUgIfMPbH63eJNsA
9R6th+obJ3ccvxUUAklVBt5uPg8XCQ212Lho4LNTFwZJu2EPMoemjYTMC/FgcCJZC1cTH3kOB045
AeY65rPZTyieI4uBxAClRZL6rGJk43EmK2dFHDCEiaTSPVMLe3x1T/FQl02ST9MCJd1GBto2oKsL
WWrEUMnfDqZkaRwgfqfQS7ASYyM93SroktodSnARKCBTV0dwbVpPEt3/pQiD51FxAPLRWIBdgz5I
IObvGvGS569c5EXHCZOaRbpCkZyjxzVQ4j+I4BxiBfA3h8JIQGnM2LyoGRnaX5nz3H0M++/eAyG/
Q1QfB+HTo8qAojKyWQpyDjJzUuh1Ka3Q8vyCG+VrAU8G4hmFevNgj/9GeUKOEO/Hqy9rdDooTQPi
KZglpaZ6DL4BfTuPPQ17Rq+JCh16zWaOUsgCJ+o6XeUG15GVtGYAd/7nVpXoXsl5AyY6WVQj1N+J
vNsLi5UP26W73wsGZj0+W3tBLlfQAOZyrVJ937WAcBpp0GgLk4LUb3X091XhSe5cIbO2W9+bxnbu
y2alGwbYllcs74q/jq537yT2nxRKK3RnYBD/QKUhr7eMtV8YoLoEXiCE0prQrlSfdiJxMdeprg+o
7ayUrb8qNcryPXY/chUzT0RfKs+umu1pVdddLkR0DbPiwFJlLx2co8/qPVSKP8mbouzqwX+xvE41
T4A+ssMS0Bf9JhbQWwHFajBW+QV3JumuD/+jyYapjnJpDzX7fAlzwTqN633rAG/PLV8Zwx78ybrp
yGVjFBkhsmcNEhutdj9y2S+0bRRxCUc/dEr7sPcZVxQ5oE1RVZTWbFQ1wfUzfGq6UCw3s/Gjk1JQ
H6kd7YuSxAefQ999jwhrX00VyRpdA5ZDcrBTICtjoes0+YvrboQowpkDME0fIemE5rbn/8m51FS4
Msie9Kkr1B9qb9c4CivIFa8L9TPrIl4UctZVXF4sEk5YNnUCCS2hKZ8wg6KunEQfL3Yp1y6S8zgs
gaoSFClEYxGX2PxE5nVUwUQkQipG99emcLmExYlhvzdr4Y/HFRhV9u0VxZ5rM+ZRREMJbsSOTfI8
HXcECtj3D/LnFHqsz098cLNj8tQbBVo4NGK4NAyWaeLk/aOIQEXHXK1+5FxSIKn0+U/abQ3dQnCb
TQ/okYaHdDZJlM59tbcaaU92rbqBYS6qIcAQN9QIH52shzC6xWXgmiR22mUj5nT0A6f/PdFsheAD
FNT+w8dSl7vGK36lBy21Q38AHphSmijPM2cz8j7uA0yL2LGzCV1nHwgqZ66iE8rOj8GGnRKHfgg9
iSccNXEwgmeV5cAR8dwePpJDTZEbtIw8079rChDEgVEGsSLIWUFJfo0ACLwSqKXUolu+7mWJxLq0
PZuBhzSHGeo/PSK+5UrFXkPo5JPXu1QEA5h+EH7aQI6N0GI1ZJSiT5AJTiTo6HXdH1EigPQzXrpA
t4Yqme8MEp6/y+GIrcH2hHZBuzRDluDmjFo9AFGWlqF18DSdcfAsM3ngyLF031+hsTjSW4n5P9kf
dcevtYnLllqM25cQB+WGVkEqJ5xJ5Pc9Q2HRNeZsDJad/efbJFDstCgUI7vIquSggUzyrvV7a50S
CKV5GB64FuZD03JlP6eVzt1XB5L7OXvitd9twhMn5sp81iJGpume1f1SwhrR9cbGyNizwL0PZy2F
4oVzGUKphkj15oZtItRD124XzYQ4FsK+boQlhSbMS6W2T0JqeNa2DldXRPMDoha1aahIF4wKN/C/
wa3lVIJjbQa5Q6KABPaAynE18+BDJMtW4j/7uCV9l76vsuykgikG3lFAeEYZpKtX+S5R9woyfoXr
FnTQKcgnnusTRqh9mNMaTN/HXcIZ9WyBXL/k+igmQBIPJC6YWxZW76g94HZtTk/Q6fffWNeqllMf
DfrF9riFCfm2o+Uv6v9e/5fF8AjMb467Ih/dTk4iYipSeS+BkVy4q1BG39eJv9QriPaCsietyMGd
oyoEJHYM+Ww8b3xHXfSo+keQoRlQXnHuOAYwXbVKv/k/HakMHZ3VW0B0oQkYz9VgsUfq9e2VUHIK
wc/gjGnohHom+z8FL/0YzV6myIcQRtAK0WCATUrlrDxaKOTRRuhiPp72ZStfE7rLssSobCmAZUtt
WA8fisq2OMwqzuBjQMeycx9FFRw4sn+5FslOolLQ8h/dE/Nx1URnFFE4OtQUdJM81gJsrAwW0qPy
OFlLARRC9oplxOaAxtQmzSQTNc4VpPGefZckVHlhNDEk4+9pj7c9zEokAtegq6eNjc7qlTl8imlb
viHtBSgIFzvngObb2HXqY81itvtj5IbtY5C7iwDts+YRs5C8n5zAgFZ0OGw/ByKE4J1ILi0EF1G+
g0e4rqQjRxhP6CBp+dAhuS9uXCAeHPNcCnGxH9TXgiX4JQAA2ujkePbgjpaDZcJ0UGCyH18sCcxE
7iuVqUFBR0QgSq4XC/6PzLwaXQXO/JjTCVO4ZM8GO6kTKctzXjTNFwmWubBvnfslbX/QcksHFsTd
+ehyUGEgM96sAzMUBORhBkcGjcMGQ5uZw1T3DzpWV5ymNSCedzD9FINmKbChV4nVFKys2X8iP9ks
HfdgmCIEQPexnADqlHZrUJqzuQ0mw8m3OW/WY6GqpqMrBu7DRnUekkHs8hflf9XKafghRT4EZyoV
Pfi+jd0aBYYlDx+Y5/G++RpVwf55kYyRMpvwEsn83QEYdCX5n1Lnju+OLILivFsSUOzSfgRkrwoG
gSqTHyEifvFQ6jRY5FMs6HcyLzanXA45r9494rqBLwOg472CLWXhpWJfKheiozruTb/i4DgNY4bo
NzKzKF2xICn4v/KBhV/UqZNNDj2V1aaH6nbkTZGJnFLrniQsZNb5qQY1sKr1kID8Hq+HwsPU5I8s
2HFQMB4Qw2j5MU3xsnTrwbz+Nxqd2GYNV3iO9/6JpBZkmN0CyjwWQbzLH/Th0N3DP/Kwync+EldE
rKpyUcwsel65JDzXUZjYjM1coLPGaEQgzocGslu741JXCSBdmNpox+OqqPMbtMjA52+ShJOsouWA
hURwL9pnP4+qYlayzVSNckmxfZ1bhtZqmY1mpR5IxAgH9DRtg9Djlqv/g9kfX8/mEPDiw2l9+q5A
hNUy2uGJgpmb7iPnF6Nzu3BfyMhVnmM4ZRes48mMyGKpqtKXykB5j4toY1+6mokxd99+PnGOCgjO
GWiAqJCF6aOeQuSby7/igY44yycWenQqGN4QqeEQSmfDTtwI1r+xXeDGup61ROu9KUn0Tvlx3L1H
84xEI9vLzRKPMjQPTIEs2fN5UtfXdi5MBTZZOCbuWD5KnoSfvmiNTxiwyNuUzQJJwRPYq1aatNwx
Fja0gB/JneLvhy6oon5U7SMmuxLOuYow8/4ylhpAyRjhrjbIuJ9UtVJ9LfRao4Pzz9PjQhd/ZNZt
oqbAJokhCkinh0O3Ys8IZ1P3kEpHBlk++VIpRIcPdjgl59xMge7LeXSUWHpeBbr6KBmvm6alwkys
3zZ+vzQff5eTnVd9/tBcStaNI5bX+WTQjQFonJFrc5PbTGk8Ms9MM/JTvZTRr4y/EFAE58XHkfpb
JA1Ekz+o11pXXSCh9hGgGuY6QLYLFNby+up7dAr0+8C740kPiydwm4GS4dv3Mj/aknak6HjIDqOX
DK0HVgAttrpTJgleeZI/hKQcG+upi0efgUSWY0wZmfV8w10qMx7ODMwHN8wEpxOKm/EFrW8IYQMJ
kS1L6JUjpp1yVTlj2t8sjlw0FggQyqHHaC3UAqEyt574aQdB0hDoO7D5P2oVYeSH+i83N9HBivlG
zPDAraFLuzNpKVacOR6dIY+XtmdurzHPoMF2+Vl2egNmVED/uVi1WBgep25pAgGznLl1eWCYOF/+
vmnSM9H/BoMMyBiVk9lJYovIsp8sPPu3XmLu3Rzb7cuLB/6CyJ2p7q0RyjLw2mNafyA6MTOlx5DB
Sx3pwpzw96ObecIKnjddgrp76I8mkdS/y32yRRDs1f95C1nanKUZCFGtOGvmhmAcWEW8ck37m4GM
nh5dN5OpTlwoJEEhjGLAfD/mx9O0rOSXd/p9hymSABqibg+MhL4GrHulo/15/Nhd+bRe1tPaoLsk
sLwCHeIOSGhDCg0lzjzTirg7Z/LWqUGqx9wSc4Y1cXAOxEP832VSHHm+tbE8mi68Szi/k03uxu0j
CGMO50Z953KY7osHlsul3g9dmzqckgcwZd1bzpYblUZKhTs6o8yoGGosMNiTavzZMXp3amBFinGl
UVSsLMGEX4obUVQ9oHDSZ9QqwsMTyaVccT124mQzDlC9zHyMyrRQnz3Fl+1AVaRNaKRfZD6lvEse
VIM8dkbPvDuRn1wI6qzNNNfcqMMqLo3wkEM/hypZPohcm377W/oBiarxnTKTypNi7q3a1av7M/C1
bUdW552UtS8qRIiV3Jt7JINPbztf4di2P09AKdUyu+uiUFFZN+2w+4Vh7jZDJuWYwqmlECs/LgFn
lvKN4zGmtbkohMjledk9IbnpuyeQ787xQsxNj1zwrtA6gIm+c5bPW0EJKrweTjryIztgODPM2R2J
gZzm57UuQgNz82kDGn2Kfw3HFCahdFy/jkbuDyNnih/sfiSLlJJTZuoic962WucIdNSQeHq7UZl4
duIHCWO+oTSpnPqtgn3Wk+OlbNDnIS0x+9WtgNodlqmWlm2Zvi0eTEVNLmQ7puxuqTP+8v3TWJsb
Wccu4fjOjAHh8ddY/5avGcOe1RKh+LV3mtjMkYH5x+s9rOITHDEGNpsOkQLSnn65fZIrs1JgilCK
no++yLG5pAUQ5WzN/z7f3/FTzNvzXMWa3EGEjGYpZ7UdFWfIUh013r/OIg1kEnPyLj7QyVxx7EWO
QItjOTfg/uA680o3RCm+aCp7NiSqfV7r6+UUN6pYR4kr4QsPLyxCv9sh7lcP/N/JVESjLpg3dkmK
lGEkXC4QHisQNesScEexfuo0xnYBApuS5SBI5Umd1Qccc1q05C9Z0jeYAPc1+QrCzaAcw2yvgAC5
nZrJhaVtQPor72mZvWBlrLnPWPnJg0gdHGdjaBy2DSRJAi3WnQ7GMw313fxNiH4WVTS+ZZX9odXm
M2UHvW/BllbTKAY5vgRnURr/OC1VT2moETb53OLAeaEeM0ZvcKy6KfHJiNYjhivHnryY8uJ3IhIy
Hqgh5+rHBw4aJBsPTyv8xw93Clz+FetC1w3KZvdAcXVUWD3b0ZepOPxZ5HtfdG7NPkMha1gYOF5t
nZyE9Bq7/yKhriVDWPZB3KEjyGe4KTpuWFlCq35mpUIrXn4+4uqt3E//9ERnNZCNAsDZ1dvMztyO
KLEB0PkreVbQmIis6TajYELgp7HEeaqlk0DuIes99aMLBXe76xr6/s8kl6BWZ89erRzNQ0ZJ3LaA
9wK/ks9qhWq+TEonn8U6m/jKWT5LdY35iA6sRcrS/Dtr5AC0nVVZb539BsGCwAngEOCNgNJJjV8C
ysMQfTrkuQpt9VAY197WakYp/vLzTt16O5gBehXI+aPYLHCSo5XKH4D1psnoHRtxN1Vx9MbGrliT
TgQJaweddEhTG/AnauDqnIiOwWJzTjzaRdrGwphNe3r+itdKz+vlTmeodUPrEa1qQqSpKCeiXDbv
dkkeZP00q8DbGnDBY7MpUIZBmOEuTc4L5kT4kUVgV8uV1wHDkP1vSjczYjPPfg0RvnT0mOnJzCKp
/QEHmEZAwADsDvcX4RR5BB5dFVgKPNLbg1gDdDXtVco0ldceiDHWi4l8lKpA1CkZijGU+1t42Q+9
vc1MdCvvQMdMzq2suMzCNGJUVe9lqHKml2W6kf4fdOH/8QnT8xYO7vBZg8jlIL9kMl9ZeXJKZeJz
ACfpUkkpuSGNbOTi2JF6GI0xlx3aNGK7ZqrAGX8sZ0zI7/kBHVD2CW4ATZCTkDdPjMyhXkSaBend
AlFRraJ70R+cbwOfkpzSqSzA/s/kC3rslqRq7B7T1OLGqRg7FrA2uhSqfBj7KxKxJA3GqnwIIgJm
ZqkyjA2S9ojvfoyfTBKz6uWkKhPexVgJMRoOJYfFW4RSRfMc/j4bROCZ8uo6wavrxNgNrnohaRA5
LH9r0Dvs30QYBKm82OgGmR5F0w3+ENeU9FuqkujyYzjTbMDwq21IDo05oTTG2gFHLlV3RW844qND
1vu5y69fw8hO3bSRmXvmf+KIPiTWfdRiYe0SFD3pAcl10X6/zOpAr1u9bt4TBJ78izMMBIzhXyof
VWYPKWB0UyttXRjFdUg+lp4xaQpcMYryIllIWms5z++zQPRF8w7f8J5xk/lLpoNT36ISGd+sowjd
a7YNerdVFjcv8d3kyxFA00Ye0UE6pGqbEahJKIJWInFH+Gnyt8y4KHVVLkz2rXEuZFE1WFBV2muA
ByhxXYjVxvZ77L5JJrvlOPnoNqGpFsay3zTFxxAoIWt1joQZyn1xw1uXqWBp3JmLntsuhbmVcWh1
50I70zap4YrcOuyBPpFjuFbz+T0BKloJW2jnH9ljeRTNpE11U0HUTJ7PCFR+bBElN8jmbSeACOUH
7bhDER6wdnl6iL4+hpNygfgNmRuzSacmjTeGOdrIRqC0Lh5f8eDUc/1MWwxZkoHkG0D4yyKW2F8T
DXLhjNnnbYb42ar14wfMuW3CGntQxfUL1qNgnSU+evaA0OJEuH8H5l+4UFUuQ4bWXe80wAAZWhk6
s80Oi/sl5JOdB3ZdiWRFX1zy80PgvjCOLY9QqBRB7++I25qqrtym7I5ydUgghohShBjDVs5oUwlb
6gcGW8kMAHh3Z517l3d/EImQU0HqJV0zH2B8l2q/hefdHgJZsNC9zZTkE/KZpOM5IUmDUWj7cKMy
TuuIXhTM6Y6oTNkx51Szk8gv9QpLNMRCEj3kiPEDnYoNkZFrT2VHv+GGqITqs4XsNCQQYETJGh40
14idBwRC1kgsd5TFgfFMli9Hq85nYJBHpsgBqZGb84wB0jG6L22DWDcsuSt0h4X1uR07hf6oQYpx
/vOspKEEh1mtIwImWeSOTr+DYLTuTwkGXsac+z9Rymof1V7gXlxW6M0O7LIg9yk9prl319IVANKN
b7m/TmFwgDbvUkW099rzL0Oct/nGGXYW/xnTygAMf6yNaRDzM9sBTZMOP29aoui6nYMjMAGHW5b6
AmRfO5lHNUqSqjUzdmtTwyQ9AmnsOUU2b3IMHjwBxMCTk+YLZkPs+QerGJL6vEE+D9QPTh9iNC6y
VWQgiSZz+rXGnDVWo6pHLtlU1UXv+YB07Ssdus/VIGKHhmbd4LsV6d5w0G9pr3thcGCu/bV1DO30
S4P6xx5GyWZh27Sjkad6Ryl+3bgJE8Af+51T9W/GxKDVLfJiVSIqsa7PX5ajR7v4hyBQ1l5CvLEm
0zuEvFgPlXf8S2ErhnE+VD71Ck5PUl5/XSUIpKja71Br/Dd5dHHoIbfOwIFKFWv5ybgvze30AinL
H2UjO7sYCsMRnFIv5LXZI9iQhbEmznSHysbitvbIxCRNVJjTL7FvtuJrS2MYSPQ2vRZCBrv+c7qT
pR5yV/sYLsdb04Qx7b+IHSf1iDE4XMFqWPPzcZy8duSv77gt+90+HVrHkfbfBC6bFh8YRMPIhHie
3H5Q/YetZnRreSfT3zdoRWD06nLn2j2CNRb/1JRApP8qGZRxnoV34Zwsu7AYZrQrqK0foRzLPfdX
tTSBbc6Kc16jAahcZtp6sDKfbBfuv6rx6uHnEC6m3Zm0PJdVtK2ShwDpu/f1FSNWoAnsyLpUSHmY
xQ0b8jp/OKsfZBVtNZmPMZpCnJ5HOdhqpRg3s1aOktGzpG+cH3+0ugj6ZbKALBqOb3DvYbFhlmLM
eUMq/fVs2kZsfuowr3P16GuW7r6WFkN0OiDVgpnnqUgxYSlKyrWRXdHiJfMk383hY9bCbZa4d9sh
yr0q0u79RT8NWy1JLBPQg+6/BcLvCYdxHFR/2keag6/mPh1FdU3Bf/k0T/Lbjo2dakTyqhheg6PA
uQVSndt1ObEcbC6H8796zW497walFQtLPRvGAOvJny0OURpB9kU7eTCEpsa2275N7CB8GytmXBzJ
xnU+vrUk4eRkdtX/TRuJHF5QB9L+AJ48MvbELjeK1+2WbaHNRqHLOFcFckoeUlIpHgUR7xVxWjGf
xcUozffpBj+ifCJCIgYKRTUO8W8/uiP+2s6KYwvr7xClVZr7eDoVcqWqAt1cMVl43eeCcFNQAs1y
f8uqcOC0cuh/ekS9qElgaIGHx8la6HGi56ITv1oGN5X58ZoWq7JUiwJxs3W5bInYNGoReXP8vtPS
Mjw0RpBuAnmMvcT0c1zyke4KnPoMzzHaMYyprt2zuGWlvCGnaDKt8MiizWjXSsBKVlj3izMTKQsa
yJjCSJ9l+sr9VQbjWqMwTRJ/zZCWV6X9hbSUuOYk5IHEoUvVakzPd6i9of/a2yWqBVlVuSDcE82W
jp/HHlNgMA0u/T1GL+ewhpdZ1QiKHZqbWNzpsLNaS5GNLujrQr8u9k+kpx8d3LRzAbUOr2GcZHEj
zS22+8tvA71D/solxX8Q+KUoZjCcZRUa3mcfjckRbj1AiFba+DuBg+3OdpI7W5oCNRb6W1Wn0aCV
KrjFmKxU25nInyhTm386CeezmTOR8tJPX4KoCaiRoYuiG94D4B2bqC54EmHv2/ELd4Stunyjnz/A
NlSiBfYJqnjapbu7+3bVI2JustvWVc3PG5+ZRCAYeFGYM0r22OHcrZi5F+aVDmaIQ1VmdjPYyHxJ
hb8YnYgCe8qKMgBYPOnqNVpdETOomvK1oM/uJ+rjK3KhHnDrnufJmVgTI9xKRIlks6c5rM9YtSX5
cPTx7VKAWQqgjD3kKYIg7cvwyG+xKgslei9uXdAuSRz0TGBui7ClgacDbYEkZ/tN4+vc3SQiQbb2
5EfHoUvqst/qA+99oYyTYuu2s96V/e43Za7ItqBOl9ckrjGlvAVNJCcZK695MCW7PlKe84ii7Vhd
b1ex/7SmaOACrQGSoJqm3xrH7tjsN1Q6rtNikFIjxon0LjxxYTpaLpTBm2l0BUL3ejYD1Gs33+hU
FJvTqjcC+g5uQ8n2zmZ+13iawUu0r3XJ7tuCSvxmkM25V8IXkMzGUCWjTmUKoipjES8SG6JgvL9J
UflkOmc0NqBW2eYJvfBc0s4jX8BRQE9ENnzIaOECnpQBQF2HQ8zQbgSNbwdTp2hqUGwghksPNFxZ
bL2FV0cAKkmlgawQK0sTjgpKYU2m9meBB5tO73UtjypRGRJKFlgJP6KipsDQ+yOHv5eDW/ODH6tU
sY1OLx/gsw9p8q4OjARR8lU2KboRzhu1qj3iGBVOk620lUB6GFkm8UgOSmCNyWnQkt0v+ZmOYmSy
VbFwZpseJn891xKjelITSx8NMT1EYK81mkRqih2lLyUo/tXyzt+jstG9d84UUVgtCEth2dL6dPAk
c6wvYqciEEvtmqs5ISuOUBZ7igwyAxUbWJC/cmZZ3WdxLz7oNIlcuaZueVasTCPxz+fzY/BbbrZa
h4RAsWEQSFEwiuGRDL7IQ8NjbnMnA7o6XwQft9270+YjJ5K+ZCG4JiLAp96wVDnzcPCCI/Eg2BD2
41vh9X0VYt85qWYWli4QUJBSfrNqKPWkweiXMAiPClQhBQoi8LHXaD5FnfoRk1R+THi2HXhrTGM0
uDDtvCYKu3FmZGAHt7GZcAFkakpdN23Dovnqs5YSaljOjSQRR3rG0EHkwddoOmdJoFC2Xu63iaut
kEeQ7+3cGnYKJkeLJgW1Nn2AazsgpyIvLVp2/PWvxC5ir0hRVuBCjeCrgB4e+gAe5S+eAilmHXZI
fhEM8bM+Qf9CUEmgxvlETaoA3Gl9VKYBtOHZnlzrvnKjrLQDHIJ8v4Ojc+vuQrGWXR+7Ftf11+Hi
SMkCn1KXF+dDL1M/WDbRZM4x8XwTatWK7X67GRG42f0s9/mNODV6NGciTnvfzCHEgOjR4eSVFDAO
jr1wDwPCZkkh0Cd8et/ROShPxXUl3osS51eooRB7+9yEAAiA8QuDmebdYDC6kGq5tIJnIHI/KMNH
cODXmaCWkPW5U9AQfkVu8BKsZptiscpOhRM9WpfrudH571tJhZe0Ca/VI6LHvsZ0tr7Oi6tLfJSZ
e4Mm1xRslJ3kKX2DUx6fshZ3Q14apV9ONkk26d2QIJPd3DRb1XZX9CWpllluRIIdUNd+aJ4TaPGh
MgwFMiauT2fQZG0LxkhKNfFrI/s4PvWYjzzZJe/zQ5JBRhtfnOQjkyC/sh7N+YD4OW0t7N8jyJbR
VpRyukX5FYWGMwb1pgfwJLYgZdOxNzkn5SqvTpUt4IlY177fZ1flXyOTjBbD7BllTpX9FSbpfYhR
6iaLUNnFzMKZHHWRqWsPBuK7I/pMdu2Kwqg8YIsxBzGV2CBz/By4ZdtY/mKWZJfh1liryS6ZEQD9
MsbE1Tl39cH3YZQpji84lQRjtMZr6+h0xCrvywQo1F1Z9mvkeaHeM7xv0IPgDgO2vQsX9vuGb0BX
weR5CKro3DmN/p1HguJpz8TBx88y3b3l4gdB0IzzALUeaoB+Rh61Z3BuQ+OJ2JoL880E/C9zJft8
Z59HYgjB7T6AUS+0OKHPDGKBUfepHkGuMF+ezngfCGEiL/36NlJ4WJctHZ4JHTa5mThRjm7DWukC
LkGWZ2jiLcgxmuTHzHMGlzgNKiqH8dvq6COvfhwhBKZ8ccLuHFQRlr11yhiwuVw6Bzs1fMbzoRE+
Pt7o4erCIDCxfOkS2d6ALAGoKBxYumM7mXHDXu2zQPhBSINuafy5gv6xs+pM7Zn1sSIYwqhMhwpD
eAjqlkvzBleobGPMWpajX3XhRZ3Rb7wuSbj07Z4hNlpZuKXWYdjJT0OwiAP7Ez7U+UudEAKLSIK8
Dmi6O1y9gffpqEnIUSmc6lW+aomyJ2SVm8JVe1Zo9hMBstS0iNiQQOV1rYe5rbbnhgxOKqUaHaL2
LcvI8G23v7FaFsJlQDZ8JkUC3OcO95F1SzddLx05Bf5Lkn+UMZkfpbimYCUp6jYPhGtWMz1NNetH
AurxBQEQCYOdPS1xnsRKQRIWAINr+rMKFfw1DQKAijhu2G9N5v9XSE9CwKo0csiXOkMVfZ8hSxoV
NgnO8+JkQmOS0l5JXKp+2/PCNufEgMaiC2S8BlFzVmNUh/EPQ05O8HZbtvK24fB4mWvea2ySkfXh
W+ZYjnqMgiUcxEw1eI8yKl/QM0N+96OCCDAduW/idbFzOPJxBYOFI21eMbKRXf7txpwWtd2ryIQi
Wi2kVtFAeD08488H1IQXncW9Yx0I1iYOwzHk5Zikik17PpHyzfqIlS63ZImahXhPzH/LmZFmZ6q0
x3xOb2OiYflEmw2D3YdlxTDHsgBilzpLksa35vOhGpNTFCMu/zR/UhxbY8QeTmNBcRO/ecObkZYY
e0D/h2R/6KAqZE3aB+ysvOLM/O2fPmgNG/sq+mwGFKJ6+Bgnx9drOtCKktzSlfSCABrFx8LDn++D
yRM2VVqBd1oC6RW/Zz5jtrEMlXYOL6jO0zHhVSuXqM/WiBqTJBtDBCK2ySQK7B1pl+xTS4Mzujse
pBj0IZHIJfz4rI8qUgw+0uX01z5jsyOjJ2bhXtN1E1LtubnAzRQA3/dfRdFPt3g1ghrTF7PSEtoY
koq/9ZSXZxjr8lsD43+sdKmuiop+RXkXbqs33WdQBSRNwvX4jwvXfa4RMWRrYOEGLmz2q50UyVS1
4dFasTpHL4xwhZxRFkxvBN78b1gql14mWwriuRpTVUaUiSVxiLSISB0mM+N3aROIKNup8dJKazXG
NHXRkuZbKuq5TtVmijbkxN0CeWyR/abwH1ib24yJyBMqlCp60HaV7lySI48HBf/U50HJhabpST8B
mW/X+TyDc6DDQK/fRBCtS/BdQdPsprXXWk3BjLT42J2meTxqlQlYRaU2D4PVaoUN2wW7+s/l9pia
L7Md3FN4sknShohtM5K1bpSOUSZMjUzjXph70DYvRwD4bU7pPw0sDtABOzV/9orkkEd0qyRfrhUT
Zyno/HVnhyiqnOFR+glrA8qAgtPDHoqgxW7v0W/CRP69TnYFClXtPtXVD4iYPW16rkysjjnOLSk1
Uxl4OZzqdMv4pqf75xbPw9MyBSOoZk97UI/7ANQ7pVyKqpNN7BC5kPuxKrar8rsjyv8z/Ol8NCQ3
z3S7bLhLTf51FjXIPz9ZNL8wM0aVNQPgnqh3O6KYw+RaT/baIYG15XBG8VfTc+17WTEVx3rog3En
eY7eTGOBlOLevXj8tjXE3w+s1Fi8PxF9SXsPl77CCsfIODwj+JKkqM3m45ZqxAuctGTkpSgmYzTE
AsnA/AcTY4uG4vHL+85ds9dKOFfukGQDidQ1tOmoRb7MoGnP0YDpvnvvVQaRvNZXp8pJpsjpwyBq
1YfzpcIeGqDSjikDuwVxhdjD0fa7pkaJ7ggSZT3v7qboKWqzoAvP0maeL+qTdXiTV3sZiSv9yFie
8GfiXYlRJ/8D3a+V6ouIvS66H8rASYCyWNky8PEpztPtvKgko32S0V7z/8gt9/qsWFMn4EPsKUcW
goTn6bWCWnecz9XCB5K9yq4SItEjmcx88bl0X0CDyLhfw9u/M/9skYuA0P+r7J31sHRw8vKJn/im
RPaknGuAW44m/jRYSsdJgSZg+MGbs9jYIlk95IeMPmmKRSyDLzaXbn2DvftX1yyaKpGbWhqiHi6Q
jLs/zTgo3DNCqipMbH+1pq9EBOx3EgzViemNUNKaoc+/Y2KEBPSyvPUqTgSQqHdHOjJPZAISax8y
YUMP2VAnxDstzbkFJ0f6c9o97d5w3+wA7YhQYtF7vsptgoOBLwVBTZCEQ96pAu72Relf85Vr7kbn
TZpnR0/wCzQ87Ca2wIDUZz9gD1fIvkanlwa2OGwpfGmvCUO7p+2iC69Z7SI8KhGAmhcqHr926+LM
gz71o5naebjjGNfDjNOe9iM9ykqBlqmg4bmRx5R/1ILsCJzXJbVFoU8BlpMF6kw7RX5RN6GAfYJ3
pq1ubvv/OrMUlntpSL6dOoRNjfMdfck8YqPpIjf50d4FeqiyCDygoKthkUWUsbHf4GKCOuhizrTh
omhqr6L/mkcz+zv0ZeRXD0J3jXy/jM90ec3UTKJR3R4BAX3V+H5no7dx2i2x4yPLeNp6PIZbcLIK
D7POK9cfcggEkbkYmmSuO7vGaGMRK1R5sPVeLzOwxZR+/zDVS0ogbFDDsSHfvnxMXUWc3yudVev8
WgDxzIS7UuQ+cBiOBHcirHodEdpH8TAMt8CYo9jKFyK8wv4oCUFuJmR0ue96hWkuKeie3+ivBKVI
9MBHNvmLnuhnHpNH9T3diSbTMkTerMCaSt5zOI9jRJ3QqveiorU3ECUDL+woRNsDzKfMdM/EPAY2
EPjPFeEz6O78z/0M5tfCsjsrULMJP82pgZ2flNiDZyWTcgUxvOPJxiNtCunihmRv/RVIRAPMQ8hg
ClFY2bxdp3GkpwKMwa1T5OvNt9vaJY9fQA0x1mFi3ExaTgobOBZgsaZezXQ4/53xs+qotDlQ8VPC
YbS1ItuJPnD5PphetSnYSVSyp6S/S9831M9tVwlscoDcGK4X1VNZiTmUEeUJdbvqrGKiHTxKvOGJ
E8Yk43thHVcaKiNFVa2NYERlTY3hzqzMfcYGSXN3K0BnXmdO1A9lKzdoZvNsoSX86aRQyFKjtpgh
xv9szjlulhz4Vce75wAbZs6D+5x6SvD1Be/HML6OGpKhjeo7Ngvup/8s9t6V00N4gKQYObC1qAyH
InhrUXTb3sRTw1+mClqmFwpVQuiLug5zJ/4qhQJJn+YlgtD0IsWzk7YUikibKbPlkg9L4gPlZrzZ
Kkb8tEdj7ZWg9+PLqF7oLU58KOSgejaVnlMN9E9Ms6OlAXVaR1QFchNHw0vjAnqk/Nyc1dCFrqiW
M3c+fIcQZM/g4G/bCIOumV9iBA3OL0mqQCyY/Zxgx4/dGr8ilJrDV73hZrBKWsKDGvOpmHX9mea7
1Hk2B27Wc7U0qJXnuY1ynD6WsgQqkpLRLpkNMSY6Zvn+qan+e2mX5zQmTl10PYKKdHvpsnoFM74B
a8Wg493QpIXjiZMeyNw81x6bFUJ/TzXctHXnollD20f9cZP0P3kwQGSPm6A/B/s9hhDiAQa5TiE8
tbDsUF7/AGziOom/VjuCXhGjfChJFN5KP+5Euo121k/fTJPdReyIuQuJYcxBdOCQ0Gsg41nEu0jz
fMRH4P3c7ntl4ZaLr+urluaK600loodGRoY/RRwazwFT20giHnGvTS5Fpx8sq6mhKkxU671AnBMh
w4XdZfhRcDjOM0nwY1T0M4pMcCuG5FFxMU2iiRnkcImdD0BxFqCPUqNnIkidLeseC345dkYk2rje
BPCNRV070aUj4dY//bhw9gYVXS/ecG7uSpsz6jHgrI7X+Y35ZlYEY5auJRO9AKjFYBw/p0qu3sLR
uk0OdAL7yJ5F88AA2ebK94YQZ7ONgOFB6noMeV/RK4/aabBjEK17XbQN5FFcNQso/nXRtJ7+S7Cm
IUEY++CABDcSjNR5YV4hmWqLqf77Lqn2nTEJYr21PSa498JjgMTZ5uqKqEHzXvfFPNgu4+td+1QT
ORvGuxTu9jdRN7bcNOMVYULXwLcmtgUNv4X0LOJjOYeqmCkr7CiqjqfWeUybpKiKPr4SVECIB3Am
+t3W5J7oOBmjF8uEnnTWBiudU3zguiLmkIN5w6lSUVJGzzoX0PzkeHq/tBOF3t2oSGb4neLn9reX
uy6Yz82mFCpYmjuXSLWru+t+nwWPwmfPS0hj2poOrEDFLpw8SfxPphe8LZS0nPqQXHbT7PSodJYT
RAmT4nbWffd0ka8K6HekHEznshuUnWDF8hr/DxUPMkC7KiMXJ8oNynbfvfNiW0fxbOGl9tNzT9mR
S41knMnaaF9cCFAla/vZNRttqo6evT0LTZi1P69Ei4LAXhRhG/1niHQKKsjvgB7+7agbO+3wHV2i
yFYjg5XJvCnNoq0EZYo236C+5/ssR+v35lEPHf+aIKRr8Rigj2IEORzWV2KGHMmTApEz1X8FhV0J
gWW01yXUxBUZ0S9SjN+0NC+O+mwXJq9akzfaqCpJ20NNOZuuiwy/NOl9XhjAyE/ofdpDe5+4bv5z
I/i4CG5Ksal2LD9vVt05q+zLBRQYAaWTWlYoPMmb1TwjC5ckSSCSKCGPpPhwdPKtqDRJ0/0D7OP5
AZsDsOncsnwkglMDukHhiiraRvVSAoqhPQUShVPR5UPaLiKOgeTbd2k/+DA4KeXwHEzjNAKEqd+8
hgA18lu6mMVTiOongNlP0U+Fcqi/vvJcV01EIv1NPhBRqpsxorc68zcZJWfu9RT/BUY4Yok+pqBa
d0ujcod9ssl496Q/U6X9Mmt2mhOUTCzXWzSrmNJaMSZkbVVLnXEEV3g2zKVru265zMrpMsyIm859
0HG+hZ2ZaA0f1OyF9B86c52YuB/uDPWuLC+OLDexpFairHZ8BHf1V/FCSV0zpkoenHEbEsX5YnKC
IgQ6jVCghbesc0DYJREcTc5Ito9XSwzl3TJC4XtZ9AmikhVZMkHytite9KeJeMw4XE8sB9wKadE6
t2DzdDiyS8N6np89TrejIacpVFFWtIdVs+kJB8BqcfaqLpTBycr5YhbR56XfSWVlNw6RCVPoSYaj
ETidmY/8fadgdi21AEgLnD/g9PL1nOjRXYY2ENQRJmEALVNTkJmAcXtmm5inem+j3go4TsOfTfeD
qI0KicnnEIgQPcaUMWrOF3CcORH16y8bvlN85DMWKwjmmM+WMzUpx4GNL7/3RK8m+Uj00VL08Pm1
XRv+1F6MQL2vFwXvmFqkovtaGjwUqIzfm+xWf4aeafB0uXZv0qBvLzObXlgR80eLBzKD4SoMrpQN
z1VcD5cim3r0qZk+9+J4T/i1U8JlaC702aWoMcbipN1B3Km4wjCI+xJ78CZUywdXURcOrb3RyVui
XZAfkeD6LNgXJWNZ6SQXiTG2oNsN4+UdC/wWITaziF4A2iKTlDdK1TPIAc1EWLolX316fTtKUPaW
dSfeL7uzyi5GKw7sdoagqonIyUubp6q5fWP1ZJ4D82sd80twEQ/fl2AwD7LvjBsvtugydscZ3rpq
+rcXneLp79Z7SdLAz17n31RC/0VuP6UrBpAq3TvvW9MbVUKW0d9gUSWv9yJR30NF4pB1pliJP96t
Sxzc56iYIDrtD0Bduck9ULp5gr2mQd9tW7n5xeh5jcJM5EZ/1Mfyaml+OvXOI9KDbMdagdfPvST+
3HitMPK8ZbeK4J6DFSCSzEB6M1aXgFybekt/ITWFGODZYUdowC+c83aMfp9peY2WvtXoVmNCThpv
WuWIYKdBDbJ5wrkY0+cfV9BoqAsw0DAUwmuxTIlKbC2Tr2gBim63b7f0RHFJ/84cYN9k43yybPdS
KYZd+m6S931zM01EbPscE3PgwZ2OBYSg0Nkpxy/NDaSDiGHBXc8EW1ajZOeapCeqz1ohZ3MT+jw+
rthrtgQFUrMFyaR5ktRW/mFJWUusO23NE7L9MBpjCjFtSqV2Y+i+6p6KaJ2iAHdIsqDTk39hlxuV
v86NdY76wLSWf0CAatFhOaZKhI8Na2vmmDnFcl+y1beoXM6LjzHH2GDcDLON/MTshkTxSGy2IFM4
VODET5wMDU6hGhaXt1Rtgn2P5AboTn8VQDhVZvBbBMLGl17zppm3bOxpUaIIBSXLRIkGmbSV6UR/
5JP50OdHFDnQJLViZrmKg/RiCvn+lPWfPt27IQcTWO7AbSdSqHMOiiTuGq4osGk3ZfjSpgF1BVs+
Tb06VxEJiXPjuH+gC7KESYKiWY4b9O/PIxLK9XodJrrWiWkGQlX4O8TtoCCFggQSDjLtIiyQ5/so
e2Em5kW25hkrv9PZuPZ2SsuIZSjaYjIk33LNZpk1tfKzL+Dmdg0d+YxquU/fPeT28CCzklf/iHNF
lnIltnqMGDYA/iC508rix3TarGG54adWUK0ih3VxAoScv2Cql6ca9DeocAyO7V345yt6qY8gv9sG
9R5TiUvGTZVVyzvUOqpKOmwVJdbFgvCGM1MX/e/2F+AWKJMg6FI/djeyY3up27+pQWCKClXqgzvo
su7RS64FjbdbDqj7NUph1VLys4LQkYQXKR4zOzlQRi3xy8VvdiAM+sTRHzG/cU/jEM3K3S3tp2st
0JBXJnkOYG1pbe0SUluSOtP3rvO/ltnNItSSg7e2cUhDmW/lT9IEJxNKSi3DRyZbP2XdH8QKUNNa
Led84P1yTm1ej2XnnH5qmIcjHYq9VviQ4z5TSmMZ6eixDnSgjHtJnT4mxrpqj4jJV+Unzmzw2314
fm6cE0ryjkTnkKCEPookVuqdo2jd2SBzl0DP2m4HDsSuL/YrVnZ9Z0ggcah1ty1zxu3fYTkj70Ce
M7F0Boj7JU1i88RzHJbRPrXnSgO44roXRog5W/+OWhTtdWB4bQT9uFz2d3UhMaOvFwVP9cP2vgk/
QSHHXQBSaHV5XkHr7sIBWsgo55Wg3jKD8aHPEoDX/9hsQXliyEdDZ5ZfHX105zZ+YCUMVELnVx07
XOguXRdbRb6s3aQiimzym+SM2qatJIoF3rkfuZm097oDw0xaTPkhwDS3RCtxPrSKb+z5GPaxqs0e
7paGwML3KoIRN+rdFbjX0UB/B769QYyUbPLECiBDGDlRk3sAaMJDLdkt20PPEfJRcp0aBCK4qYd8
S+9j6oTedrRBkgBSRIlJ/ESIGjrDeQIiA0oKLINRlFFF44/5C2eg3surS8dZn9DTaW6xClnLOcw5
haxxWkpUjUP+pnlYKRdazpxPO55GyUM2E7+VUFDXwrM4H6l0q4nXgbsWkzkS1fkDGTIAOnoi7U6R
JJ5hja8Id9tLFowip3/wJKlxrU9yyhQmhThGzhbj9aLcamt3OtUvpLQwkO5BPQXtSl5y73hBOs/L
aYL6XUzgklnwdYepalX9FCaa6cikQJT1Mi3EYkwjE4h9Ir3g+For+sCkSloPLuUSejQh3klZkR0H
GCwRNFUnSIb7tb1OuZeBUCMWAseMOP5+WCJkw2wTS28N49iQdmxN6y9rh9Ia3KZeyBwPagris268
Ejo0UUb8qAUXrWgaXzcwnKiwWMb6JjroSo7wryf4NhYq7EDZvuqj5hgutZJikw1RzzuL2shxqkH8
4MGP3OhvdH4bagTVNSZshSj5tvVzfzhoMnB1NbMaNK1e2uwfrK0V79PREaZRjFuimc2DWc07U9+j
sE3JVjyuWc65pCfIRdfwr1Uu9gC1ADLKjj4HqlR/NsTNdg7gVbk1s0zqEwaixB2z4hH0rf9m8SUT
SAfQ41LC1B8sHYTkKGAswvXiUYpsS58fbRHDgNU8Po0QO7XrVK0LIci0pIiKuOMQhebx9zpqjLPo
mSrHgoS1hGO1MN7G7dbJr68DemktWQRIoiHYx1psqY859up0kLHL1yYPwd1ZzTAmxNIhGogWiTPZ
dCfegINYPlHC4rSeGv0rrBNsAvmHPb9baFl0hqxdWgqf1bwU458gqvYjgFu+Flef5HqZ3kNRl0nZ
tHyvnBX6ZHbFCf4O3EVHYltVe24LxxHk0dZ5er0FvvXMtXOl6wGFVElTTCLK1znS/sFZ7jPlt8uj
IxK7cUWju5gig4dgCAh1rvjtZaKlRWcRaA//9VtOZj6AjKts83JAsdO6qgxmi1eK+VoJ9MrnxOOi
C6EKg5/M0w+8L/cL24gwW7yzjlCuTxS9P4gwf4XNB2+i0REdD9bxUZP/6VPdxTvuuJFOxPDga8CB
tPApTLJw8vv8yWa5PBhNoF1CYh66rnGosVYmYDk0L/DZo1tDQTlycyCt1zoqM/0rZSKPmIq9f3I+
KxKDXdoyVtvylXnqo7v/RKdKFiEZ4cBKOrX9Jo73oyVR5odiAkZki39qTwSTIDC/B6zj/yGevTW/
6SyRhn/EXnIIPa3GTSwyq8+24P87FpQ/EXAhx8GuJUvjfNd2IS8jYYoQ7EYka/zmhYeNe/nS4sBc
Rfb+E815/m+Po4Z7djC7EHRHM9MQEjgNctC5TIQkGWpk9f5dM3ebCpn7Yd0IYRlzYawxh7JSiRE9
02y2WZ1onPxlavPBWmFv10HM8o5wkcWvMm1SVdRbnsm5UNrak9KyxEfiaKeT9xJRhhR3ntCciIKv
OMRL8Re2NR3o0PfeK3aWhVhoTc/tdG04GKDpfT6346WnyLiNCR2RpiM3gwN49Ba/QnNWCWLtw9xe
HK65CVhXMK5wE0I+twZIosfaOFbROpAxlkET4ngXnM9ZsklIEiSThKgYyJsFCyK7fmfGG4jc7Me9
WJCI9j5OPrJAKKLB/pphN37VyClp4uHkQ0srcrs3VZStLUtP0IVTDPWJtoHvkZkRCmY4QROc/JQA
fyxJz1OnkP/SSeVil+bn5V71J8mzoi60qsSVpYQa/nNSgIBZbeeDuKt4Low6IKBeBIRY/Oppyttb
IafySDklG45McW3Gn5BeqTHHCKvU76dA0JF8tGS/PqLNR48YWb6DYsKu/SLCzOtQxrd8N3EC2NLa
bqEnzmarz2eiLv5OUVAAmqUyzLLz0EesqoqgE3RX2Xx3EcyTbiowVWXMO7i6aTk8nKkl1OjePf6A
yjQ0j/rbnChCqUf9Bc+U8sjs5gHqyBX3OwliI9Popq465TH6czPCrnatLv/y1gHQ9LjcWo3mz0Ih
lAVjZWSsqFfezBbRvfvCA9wo30Gs2CIBbyaXafSCHh7UzHITgFGz/iJjzIjdHnsK8VkCAz3EF3mz
4FbVtorA9qS153bVos4Cs3PE9RBvgtfbaokh+RsCO4AOxz+3BErZUrLKcAfVhUlmzelIdWrSVNwc
jm7tWc8l7MUDh7klnNw6kxavwEyz6KUFbz4Y7BIwDKwl6UEvg8FHPg6AFOaHW+EoRj1aG05DhEMa
T8d18y2NBh45l8JbqQis58fbwgpD4SVT7FyZfx+dt/To5sEeqR1LB8e+M1RdbInscrUyQz2vHIcO
QvSj8xdEPRoDR/y1lpgqHyfjJYD8pkCUL/MI1uqFyjQERQ83kUbnvHMsL4QWZlz1InD8+bJiw2xH
38zIuDfST3hDQ0REUv+qjyQiw2j3U/oQV4I8mz5vwGcH9uVW3LKhbH+ZfHCrg9/lWEWbqll2W+dN
nz/dWR8qi1L5mwrsAga+tnmeuy9nyI56ke9Ek/4bm2+/SMwykp8/qduu7GJa6Flg4AU3xLxKJwUN
ggh1wEa/a/jTqt3gdtCCN3vxU+QwCGirMamKK12denVdiLVUyyV4K0J5jCX3xD25WfHMkL6kOhJC
L93fuW5qOm+g3Hf5PJQbNAmdC2mMIZwWQniOcjNJYYlkLjiXjCInkmIxmucmeM5BalxyGnH8tVzk
yqCHkH4Vhe5szRJpYhKLSpewKVBKBfDJWFP2wPFpcsIoZcfit675eqoiauCh6jIrRA2Tx92sUwTK
Wom8+2rxuSnFci9AIV9LKpmfm7ry63Nxm6V4u32764s/fYJgiQc8Vvgg3znEgubl5Id0bY00tbzE
M8ND4jnoHf/ThvTvw+/6eOUzTrAmDMEHYJdO2FyCI8Vr6w26i4cqDgw2JuIkOok32LECHnq5TrPo
aOVmM3u80d45TLBRMSoLspUUQ6rCVQUVFJ6XrsrOMz9TvLojHBgOo2pXWIdxt5lGtP0IcdPqt+3B
oMLlWXWo31awxT0c98QRf1B2TTKLWl3FAAEdZ3Vx4o9V/krOkfIdjjksL/4pvyke2Ntt5sBPkzll
P+UFbjnf8l8fbFwdGRe8YOqWlpZmC1W9r081nyQPRu8m7Q4adP0Oz+hkZ1iE3WerCB1bW10HV84C
VLiELB7b6pIdDwmT5RsNAYPFknX5Gjnluno7OwYT/NHXSLGnOzfdJIUh9AWXgW3bgjmnk6apqBRz
9lXYjBmQPeADMiLMZ2IXf0jKglB6gmIYpMhyB8f9BOCz9FKcVjsEXdhonRBPsOUPIdekROWW22qW
bcgZ3FRzPTNoczeCkV04XlpCMTbECX6DguCVRj6YEO+YaHL6BmbYe/zBIby9kXynw7qGejjO+9/O
kzm0avmV2R+G0AGipLZKcb/myDK7jRyE0QGCusnSp3bxmfLC93B9vW9eWK55hFgpFm7NP84t/DCs
LwVLzFv/8i+cZjCcMGtcuMemw38nTFzAmtfjQTuhOn9pPYJKWdvHsduFaHMOntIr9fnS5depBQxT
4em9K0Osc4UDWYdKJSRctyk0RU+BDdW7j4EtzT97B4WD4l3ZqJ8uGscl6we5BOlgReAtXYj6ltBr
fWBZ3ij0NIkoCa7zc4W/uadEi2L++GbhJeaisbFWX9xc2QSHC1I9OfwzgNsQ/Nw8XB+ccAqvqcV0
xh+buCdsh+0hrXs0bZBU/uix9n8wbn/FX8ly25RNIiLqWLFzxt+ZKjW1VmU3IAcrWFVhRXpGKLmp
ztZIivynSKzrqaA54vVNzMgdnWCoYFTjLjTVK54OWPcwUQE6EAX+z3dd1PjhAC7uSOU4nEi7B1h1
8JnXJNMkS6pvgLYn+fnwq8egfe00ahjC2EhQqivFqUHVbfBW5BUvN+m5bnUqPc4jFdArzfp8wISE
KH3KUI9ZnSMiTGzanRDNAHGkcvhVjenUjWPsgNmnumgQzv7B69wAxbEQtvR8TGoO38A0sNrO0YiS
G/8pmoFr2FDygQ/0vYQqAc8INh8IioVy9/uv8QD5XB8x+tVijq66XNVJKns5YeRv3t5f9jGQuAQQ
z6tuDIcY3kSLVtZgPiOXYUOcvgZkgqDU4pdEwDvVE3Xx3nK7oMNim1jY+8P9nIJg08aKI3Dr2I6L
8CQ3ig7QFXPtZR/1uFd1/+u31whcvFANy4D5M2eCLR8AQ9SJzFnagSEtedgQpw+5ruANhq4b5N9Q
yAk6J6vVs/apyGQ0hOYTRox6qiDcz0qfiXb2KMCvPos7thBMQILEYmJPvxPp0Ix8b5XP+lHL2udZ
ymQcWjIyIwPw3yyJeMx1Qx63Ll4X15K+FoxeKyQdsa4ZD3PmUmthyfAVMUyBxsb5ZRsHribEpRAP
DvYMSIp02JsMUu2f6KIfDPt+3fyIWWzkSVbjIGqKUvSBgyv6s/aQiEOqHFacePdHF8oybr4cH5fB
l0arz6g6nnq5zJpqQTEC/H1OG+mE2/LT8I6OtZ4UIuqWc5LrqBoPbKGVbU7yzdXLPMQs1jbg6n3T
dKSdSFeWAP1gHhN+OuR8YQNO09hk+Y19a+SBCqYrbR4ZPQJE1krgHbfUmybRf6hhvcCGNj5Nxj5P
DFY57yOCw6W5Yip3VozuIEVWZnerPtvEXr+/Nxe5gu2HKlV/US2768nfJrYVJ6MTU2m2y0yK70ga
n+ta4f3EU5W2crVBnf9FhrSRIaUP8QmLhjAcnxQDW/ulLTTf0wWZgNC7cbbLxqVzrPbw4NnSHIcN
yGBHjrJQVh5oEdleqVRls0udocfxDtpwN23DVi3BELh4WWJ2iAtDtm2KfHo0JlEyYoUvr92yg3su
qGd8dXTGXPiq4DmKaVOfGxY7O7tCJ4DsmjTYjj2NsdQTlDE0pHljd+CTfHRQX0IfSX5PSd7DlG42
U8gEFplf1KQYgNyBtZYMjHXSLVi+W/2zuTeCothdq/9kBDQ9GIFvHvAc9jGBr1VXVoC8BnsRLd/Q
8sUEoYqGXYmArNGX+gzaeTDCEhQwebsn0f5kQFgF8iFNGloV0qFZVf07Ud7okmYnt8arlvSGjRKB
47UNV99u+9+S/ipKZF9sFXC1IxuS+gjMZBCC08+nZQfBz7N8NBNQ9Cgb8PurWQp5JjcJjqgTo3Lp
CCFtwb+G7ca7XGgzPmVpfLak+aZY0iJLiuDHriTZ9uIRd26Ns6jbVasb3bsvbcb+cImxpceWWana
XeD69vGugTYj+Gh1Y7Mg7Dmf/M6gfGg/of+p4pQx0szxM9V1oXZM4xUxhkBpT5+XjJXC2XAhpwkr
BA4+/pyLpj+xVhnB3Aj+U1O5T6Sl2RUaHtQoycDtAlewALDYpOlcUJenudTspaCdhHRMMfKRaN2y
hJSW514wM8tqWKCSwMbaz/1sv2+vOBtnygsP5mWNx9kX8egrKoMUxpKrE/JtY9O4S3377qAI5o8u
PNuYkdRyGEE3hrVT4VGTheqQ1pJWztTeHwycb0PUXRQipgwLLUCizyaS6eie1anZuRibouH2jTG+
xVgekCwdqOyHGZRJ0FrKg/eOLPHwmcYWhnMl7/FOJuH123a2t3cLaQrpPF0i5tgKYMAL1tchGV7q
ZI66zaRfruo2cjUSpD2l6XXpp7TYEnzLv0JK6sexuZ6EB/xb5BVG9hDHqJvCi0viwsRqlgtXxeB7
xuwXMyBPgLu8cYcj5XVNK6qpWrDnt1b+ptGzAgHuVZQOx3pn2QWYb09MpXNa8Ni93sv46smKjyeb
ZXpqCJs1yEmra6dZB2qGVi1fN9x2/rCgEZoRgkcOA06SXA4cI8NujWDgGbaB0ZEa9wMmkQGpr65Q
x2RWZab0OlS6s6OHpqHrXdDFdG78wOWtwWCw+GSih4qGskkiT58Jlybi/nZnOODAW4Db4/y2GMLU
f8p4jou+BI2zFms8ZEdINYwbRWR9Km+QJSgpnMPysceMBeopklwHSECxep8GVBxT2QPv8MCty1Wt
P7zmY4u58mhQyKREPSomF9ZcQD840nPe0W8JlbyxXR8TxQt8wWvwrjNYbGKXxYcOEFLZEoErGyCf
/KouYsny0001edXuZl+K57aPq143l+G9QQtUh5QWqikm8/8PT3aRrV9CWITkKt1K/PgofOPEEz0w
HyEcq2yH25pxbB7q2As6b1sKswMTqiKKcOgbs+TNUpSzAkh5mo4QbQ+G3woVMmJpvbBsDjxszxdu
gStf2JdiyxNgRBG6YbCfFGi9R2zLpn5ASMLFhLt6aXvvvC9+3s96LpOIgBe4d3P+Z6Vc9KTIsh2Z
WeJmYV1Xo9KY4sLwLgU2RYDYqafsp7lxnL6rlyju+AeTIPkufzBPVMiXVeLSdOhwFt0TSxgnqRuL
nuvASi9aYGEVFkoO14AGBd0CKAZ7QAoJmwbuwMuX1meGLZxfST8A3r2GjnM4YEdR+JSfmGM+/bzS
V///1nu80hSyaBRRM1IZzjINPsiia8n0IJJNhrEVV9zAO4INCcT5cz7ttUEJ74ydnSBc+rWkgO8M
PylLE41fOf0nubQZ/SGEW5j33QEHrkT71HUKxQ5ClB5wdB9fZ9JpEtMOuWmZ90cwVczyNF1w63Y4
upooYRqnZdtHxi1ORuxBm2bP6yEo02CskZv8v12hU0/KZF+q1LhoGeJPejjzcPil7aS4NL1dYMj+
2wDVVBtn1Ld5DM9RLRn2raQLwlvDxX2ixzOhxkRbHc0SVa3sSOjkCcq09svbib0IZvaSfx9tA2NH
/c4utNzS7ygyEmlRgPXJ6cPsifxPDwVddbrtbZBpgjqKtK1lBki4rONnDGuV4xswMC8V1Yki8GeH
ZnX+TYYIVFxrIj1ytcIBLkCOHVG5ST9EKJvxHCIfeSg28X8HH8NdPcwoyYBChW8I+myNO9rlLhZz
KrXc8IA9E+fTyVEC+4p16UpAr7us3kNp5aL7jiuNcRoD6cYLwCs0k/Y0GPzJsqSIKnM6sNx0YWWo
VCUVnxOks7d5aZHAONbr48uxeiWdEGIeY2gJ7or9p756pdB1zqp7SQBmrlI8kPqs6PbCbFWrpZhR
/t14BQpv6X3IlxigjwRPq1S2v6M7s2eGyi0B49nmswwCStDceWC2nqNBs/KW0+Y0hhfeSQaarU2M
P+otgknRmL7vpobCKSDK2WjEXQt7XdSoYqmqJ3J9+EtL7seR+dTQDPAo0hank5VQbDpj/Y9ZTlIh
szTzqPGp2k7y3CHgQoK+aR09F3XvbVWt/to9ZXu1bEpTcL479w1ofqfZeVkWxIsvuvI7o0xkYZLV
T1b+GGEhkRbpXx+FfPdWabJGwqrbUtAMb/2uSzmfGF5mEKlK2I+T6YdjdFRCy7nWU8sUuPxd+R0H
8VA7KigAojv/raC82D/r8ugvbLwv33hTlIlza3cuEjm9pBJ01GFsyiQiz/PsiWOZWKwiZ2rQ6m2u
UMuHS9fdzYF7yc8wTDEeMk9YK1k5IJ2kCZduBDuIaMbHGSKAMM1s+NT8jKfYjlgkir3kV2lprZA0
dPkVwyhvjq8hzb4CoTVoVL/CGrOOxFzy0+SBlXbhm9oX/z/h/wQbU0AY2+NA4uwYkxW4UJ6jkPdr
67yU4f+4J4AIXm+IWyp/tbnq2hHfvdyoXKsfZxBozyLE4mCWBSXM8a22Im2ZD7+LQxlGKCvSCKgp
pt4tvxE+zbWjqrot9GBleimdXfK4i8rSriHxWt4G/w/1ahlcWGyC494mMnPeXGvQPOMUbh+vDAud
Bqdd9J5IIDG52CHQ4sTqFs6GmC6o5vkjHr+tXDR2EfE5kIIyarf8r+qdqWMJq2VVMEnUy1UvdM7D
tOoLb62UWCIyfEl664t+QENUxYL9JWHO37TSsyZiPxr0TWQg3u+6CJYCx54aNhv6phIYS8oqDORC
rrEZ95TvEsmzQCjqAcOa7kWCNwl1gKs/rNtshKacSSSfBWDEs5/hgdl+4XfHvPtwhy+PhOF/VDOF
SKoLf+5KZLL+auovEy+VgUjanSmJ4oLr7OGM9JLqna+OSzyuWand6Jy3iCAWFmLAo1hzbWWQojbd
ykWMakDuJiqW9ApGhSd6ZEwP5HQvYV7zhYvM6BSQcghpubhspZHsU3DPi2eiT3ZJo79v2MOug7Ot
iBjYyN8Hnj2XBQqx7nTJrEv6aT7k3rboBZbYSWoWD0E1fQEsKu0zDKgbFXOW05R/cC2PhiAgBuQQ
hRv4KlvE2inKmGZ1+GMtxv+6eyR0sqalhldq+WepLS+oaUyOcYkXnazk1Y4l7r0Z398oZDkeuwqK
NnJt8e4COIB7dlFvg5CzgHZQbwvEQMfNLLOuOaIZ3wyegC2GmoHq85kSEvAZcL3zNnTj2D/OIg9t
dWGkk7JQy+yPRlw4wFbdC7gZbE5xfZm36RLw5OUJl3hhGGwTKJYWvUw/7asAe1ctZlGqsx5IokXp
Hqn84/z953G1dqAipyXGy7cHXudfBP2+6hoHAxjxQgvQgrtn3IE0txJmZG52S/fYWLRz9J4ZEpi8
/iewYV+mFA8E6PzhqGHtivyFrAwqmtAbatBvPe4BoE0BSN8TpDTVexI3P1FfYWu0W7bJ9feM47fb
I0aZTkU3V4un3HAU5NOPdJXFQ2J9yo+BMQrwhA2dc2RfYswhCLqFwrtUJ1xlnkuFp5/SocGsF/JA
HB4w8mC3ECxLgC5lQHx/Ai+qSKdwNz2+K/7Yt+Zf7I1NswJ85DjmmlulfvmfX9RXF/Yj1ynkmmqT
PkvJHc8SdxPShuC0TU+i6uyl6fo4kxVOss3N708nf2PQ8PDK47+LMtD+6s9EfNt72rkzVXryxcr0
s+KclcUyNArIduX680yGU4vYbKTNl2E6T/Kvgnh1Wo548PJ9SeuopPml+sumpgtOhHDOPeamQ3WZ
fnjQExjukwz75ioFMdGca+JB3blJhvGhsDQzW8LFoSC71AYEu9q9BT9OmTjy+KE2WWwANdkUJr39
m/KqXKwbwVPasoxk2Xx7IG7P4XXPg+PeTMyyXXEWdNjD/2WCOKZ/KvMDqd/1g5gQarDK0FPjcVAd
kNybR/C4K/LwZh2qBLQW4Sykz/Ymcdwmx/OSOKVlCrtWVWclcojTkVzwC8wnMB0mEbQdpNwK48M4
sKUqkAeawlkIidmK42Ar+Lz2Vic5CaY/iim4Z9hHT7/g+/MAiw93QTk00MJQrUoW5yO8PNvnax7V
NY+0dIMBnqoen0Xst0YMRcr2W66Wll5TZ+4DeUjoQUGsP/Zt000fMOwwEWcEQSD7anaagSmeKlHO
6wNSIYoRJshTJbBAmZK/XXRGXauei1gIzdo13jtff0Ix59ZH5C8elbEn5yANDVvfUhZB5cbzbIKS
ldVccNxWGJwkKvthS0ghabRgSGZf6G3Z26tEzu4S/KB+t2tOfZNA6yRHzXgyGN+w3lWrZBDLeRkg
eICQEz0L7dNfEb0njeb/jA/4fCDv8OPgaq066TjBQVvQQGK5lxC54u4K3ll5ukJTWi4na1zQEIrT
uZif7zYLzox0oLJJxjUB/wrkhrl5k0apCJtHwPZM7y7q6AsRsi6ocRp03s4TrAbrPvf6BoEHfqG5
COSBvPtpiaGm84MEKd3Q5hAJXa4spWj+YoLvGcG7NnxTvSc8gQGvFPF2lTY+OJVo9Tn3t8uxDRSR
FkSdxMUTdOjtoS+BwLApbDqlSE9FPR8n8QCLVOsHJd+6RfF9vvQHh92awyeAcBlyTQIUTElLWw7K
4WQPEJMAjNQPlimrEhjeMPJINNrVar8nj2OeP8ojVmaQ67hM6LVu9Tm6QB+6fFpnKoM050/aw9KX
nzS4PaUxkLkvVgR67qeEH5z2ptT4F3Bc5eZ02vNYtrJO/8/e3Xe+ygLlP7f4PetOVj349rTxrH15
eCfdNzEqZbviZwIBp9MUnA88tYc6UJW0H5Zufh+QdUkxnwfz7wDjimMEmbgmIQQqWROdju95cRi+
LK3KsLhXvLMqmpWYIOUTbs5hPVmbsTLGcttB4Jtnfh3TGLHjLuk0ve4jBL3sTdymHU1G8+38AxGJ
SPt1Nn2QYkwT11fsMvd/7pLDov/d8c4vUzmFfWv6nhfLncSKdEtWXl6l6fohoFcVb35pqN1XDx6F
JuyEKvRd3R3XJPyRKOm0n0Y0lOTM48xItSXRw6URwY0F3tGwFbiSTAi1+uaH/yTP2vg45K1IwmBL
P2CQeYsz1WQUamHTRHGWJfj2hK64F9eENEuYHiEdvlKqtAdWy4m7a+WwnnFDOizW0V/kdZPqGHBX
H1N34WJlppu1gJ/t05f0vXpi20ylAWuCA7HxthcZa8CQl8CBUtKZ3K4enpd2Gig2iOKzdhNSxACO
V7S4eX37UlDHCq00ksiZlrVG60KnR1WA4sMhiY/hK4Z+7V7lYcBDXcEIMaFzJHyKhGEFL61ABNpI
6AV+AEH5wQ+2gH5/8QJkjQmDsPQaS3u+eXcjBHnkLBrUkyd5L6ZRtK92+6vLLtjCIELkDzX/2Ci1
pEP8ZlgtTBzOo9+HPN6y/NPe2Md+c3xRo9oHgrUmefdrWOXm1InuTU4cOot2klT/HS0YZS7pGw3f
6FF2N0wRLUSuDWjSjLG5UAKq99EOu6b3EfM2oh8QWW1VulZ24xj9nd3nis9i0nKOMswuBRpbovIJ
zkPpf/94U3TLnBQ5J0lHmVSArQByGvM2Cc3uuqcRcyUSEoxIG4T21J+g/QdTivVVAygT2Gws50ib
iU4NGjNH4pVtuSVNIKzpI0DOVRUPqghPbG4YDvuJ/hpUV2KIXnhiGmvZz8Ctf7WL4q2CTryhGw9S
0a7iC3wspt6BnHET0oU9J9u4Yfg3XeOeKaNPOsUWdmvVFO1HvrJHy9A6emGtBxqqOGgnciO2ELTV
sDg8Xn13n9dfV1nNqJDhCr7VfSeeVrBcU+bR4GaqxMmtllgK2tJQzuP5dCvSb8vunSYkYJz876kK
XQBHIPliKQUEoW0hvUcNr7oJsRHWCEgtC60ekL7oIJhTHpN3DzDzPY0R37jbbhPCH8qYruJpRw8w
8kNAMWC791K3WRwR865ePV7bUi0rSI5xvH3P4RAZJlK1q3HC9DjyP+xUJ1CQtV8jOF93r11wXqQW
c4rUJ+hEbfYDtCiU6BrruSSOMvFN5N/1ObHzEiU4zokzoYzsJu97zpKlyNQyxTeDTYsh+nL2UV7o
GBlljo/CghgPYTTl87B+y5YABpd+8z02ONYF3lNjZ/rXbQHuVUsCeDjarc3nQBSrgucEjMZe+uBT
cXLz/vKO486hCIdMf3jNH05oQrrH7NwSNpRdvGL95aP5HwFzNZ1by8TY+Ms9UgBehz7e29ccNdGo
dLBk8Z4Gzk8Oz9IJnYJXjqLSdSkbWjPV2IrW/7+51GV/mHH/MGvXoeIUtmYAPfZs3ZJiZERfrDX4
4x46ImzNmFGOPgIaBQT0E0Ko0ytOHeGcZfbJ0lYZothnY/iks7qY1iNnW/YXvo3YriCK8wBeXABy
ftYuffbyfIWzJpB5oe2g68aYWQCew1LSLQxfxIOHa71HFTZ+2gNQTkjekd55RNVJRFtxCMNAfubn
MIDKw5PTR3IUXDw4LusHwqE0rae1Dd5E1i1UbzS/1oCp+VNcBFThSgBe4wlX8ufGLWuqXZJnnB2a
oUdOdriYEc2vMPk6CcHm80pAMLzOHNLCbx+vtsIzAcPu2bvfIsmds5ZE5IxirH6hGZo+e70UqsEe
7eu4g0JHWJceEzqcuG4ce7aNDVB0jmhLQKjccCMm4EYL7NNhjbiY+AiTbzHkCOabK6pvz6uhdMwh
W40RY/ZQ/li4uZl3XtwwSE96JckCE/kLyN38a7B9xMvOW+6pT4LEd/WGwFaC/vHtcGYm5yG7+Y3J
qeoBf76xk+canIPbNebTcYWel1tVSMeVB6/d3ZiKqLLSyT8hidfzqfcDMvZaepKqImY+LBV3k0Vr
LZMwdArCANgo7DJpuLaljvmnZk9GQJGOWuTCY5HU1qvejbKzgLKaYXz82SOEK/WO8JMdx+1aZh5B
1E29nH8Id+aU4xV4MfOgsXPXjYEy4GZgEmslFLJwhhQPeMN8ESqhDchHwr1tz06FnSbXh9bDVI/H
ahOFfTOyleninQTkBTl0hmD9jS28atS3HVhUk7FaDDuIySGh3k9509DZ7O8KBjtIPCgvZuqqz9pL
g93hpK+5TFlnPlsUYzYJjAvfE7zhtInFa6neQjHNOKFhzLJYoiIB1P2GNv9ixeTo62bq53lCeI3C
y+gx+Fhm52fZBw2pvn4hHBGfSC1xXrgv8lAE6ZiScwPIeQfs+sI4TMdRrQOzSWxUZGWxWpXkNwjx
x5qZ/b78qWcLIVYLvrz5bSIBh5+1R1BCtrZyuFB6IrtviUR8d4q4OsHARfg8Pfw63b5Ug+4EVQM8
joz3ViUPMPmMAs6ZYzLt1JBpjRDDp8tmBXh3/nW9eMWGnbn+9mSeiABXzeoyChR3IZFdWQrcn15z
/u/QihXnnD+GLhKZAnpMTNCljUAvAeqwLibndqRGY6vFhmcyqzKCAfk7HrXOVvKFYd9f9BLSgS2t
zSO/xELwjBSRFn012tvvMPV9aZEfpSMxAWbs+fY1eghX+nO+yZVI9v4QFNiiBbRKVs2+JWX/h7iA
UcdzsD2m5dssq6m1nmE2xYc1sTxdP+NdeV0wpMhm+mFwhAbwulYlQmfMFfKHmkUBbuqgbOuQ47bs
UVRt4Qdv5p+O2qisSxElHlCiRzTnG49xpwZPBCKecE/ZQY+lmx0Wt3R4L2eUuhFEDU/R8pRb34QF
VuSCzlDcIv1SRNCM+d6EDIa2vU8ZD4MuzujNKlKI4sg1bRF54yYL9uBVrEeJRh9azKs1Or5pHtle
wSjUUUtpvy8Vv1adEoEuBNyZHnzz0cQUMjqiB8O63AIz1rDHT4oJu9Nb2dacxNJaDHw8E2WWmCat
NQ3ruEzZn+9cT+E7QcHXhPWimGdPlm29N3SvwT46162C+6moMxCAv/De+BKhPSj+SARHY5na5g/G
wOH9nPhllCOp+OSMg51juFnZw7GJPCkGPbKwOvTCHEYSd/9LK5Rw5DlodbwIAwPN1EGdb/iEfV6Z
/1CQKvmLnj3hF/G57jKAtcHmKxuPyImN3vgdQtOQhZGEujuDTCqG5mqRHvlQkjOAmhAHAbmeKV4T
riTy+jMSHnC8HW7ksdmTJ/xjiGBSgkqLoKzN/eysLZbiXaWnZGzJfwiplXKJUZ/WcvK0RgTz0Wis
XU+gmfGe8GeuXmpS9DtXSdBNdiWzM3jiwzdQSEY7niagUgkzy27MORlROhwOfnayru3RZ7IjXg26
OrxIEfVZO6ze/b2N1v93KnvYUmQ64CUerkN24knkXHDfzjKZZQgquViv6OLKr78VzmYHsKDrja9H
tPunIkk5ow8V5gWMKuivEGv6dHJqROzH71nr0qwhGiPqionk/S+7OsGZlCiqEB9VJmNft8i4SXHv
RpihN5NkdjAaBWR7/BEk/0UobspRXu0TkEmcOv9MRp5LcAA14l4LyNQC+JqVv0bi3cI+im4XQvAt
JNZVA7RmHJfmKkERetX3BHqg+FJ0rBxj0BHZvIhHhrxMBBhX49Ussq1ejEsIfqRCwvaTeUbrOrCG
9vmAuH7xgptxifRx2/7EbIrruhF5UwdnilD6IcmcGX37BNIyGNmvbmHMCkJJObIhNbhMLq+oQSMC
6itmfuufl1+4QoC3lUQqkoERX7iqtXNk7cu81XCwr37bCM86QYGe412bnJqZBiXyaRPwLMmwZ7/Y
+ldTUxy+cBngvELagX0VxsmyiTuKP3oZV8XCgBLB86+/q23p24IB5f2pulsZjrif12Kf6AyX/Rcg
Vu2uRXXdleN+iUSPlbHvVeNA9iUaoPvnGy86B0//+1b7LyCZxU5I+QCh+OCcKe4X1yWTuY1tXR8c
PvhFJgNaPfOfTlGwZtzIKfW154Fc2lsvTbfQb63XM2bEXtiyKDR+R+zzCRe99p2xJ3ae5496XS3a
GlSGF4El/JSY3CLl8xQdsDTQhT4lIsUBRefStuyzXuAgWJQurddofZdTpI/3mMwdfCX/WXrjlJHY
V7CzsU/82f73nZo+8ESq3y27l6OTw8jHpZb3TFydeQ/IhlVOVNBhHkYK53LXdOiXYXnQaZs18cdu
0fHl42gyS1K1/Q8enF1VtyQTBJAFOl5yNboJctw65P+vrmzTWPFU5uKrGl46uoTIhPhlX50Ik/VI
8zBctU/J/dAbc73cX28zFp6B0POJL+IjWFdgPg42qHsLF8f0pcPL0cmqzpvuI4vTZx2YBZiAhdxO
SxwDjq3yOnX4fVBMnEThu9KJ7cXlMnPiryaL7s4irjpb/RfYTdalAR+ZktRekwY2X6G/DUDxtedq
9cUDsrLcj+nM8dp3zD3fMzI+O/AMfHw27GRY2hag2v+MRGTewY7Pqg4YRAUhoXFJ1t++Z1vGQgML
I9wx10p+uVpO84Gf1AMbovrNRPVQmFZzisgOT80Q/OudDBWOTxs/ej5bebBR8nFWRZT0QZEBkG4J
GBWw1lCliO2evo/ETk+wO1EvhgPEuPAkL1T8+GC6zg+rixx0dEtpsUXsPraHlEo5X6L5tmsxfZqR
bye9c3yzLIll1BciplR2et4XqxeVRqxFF+tHOlD/34SqyDQfHY6+5p+QfQBmWoDBORhPegsi6dHY
fDjvBI9toeBasz05ZQ0Dvi87QV8l1LoF2zxT0ig3tXbCXesx9uMWgrnbK4sb4gzdegA/y8Bu3yZn
us5+OGzST1uw+RuwqvixWATFbM05x012Xxd6OAxs3FxMQQFVJT/sHsERBXn9t/U0r+1zRakpsRun
DG4bag8H7UGfGaE23Q5TC+qC8RMZ62MCCzzU/GUy4wR7Bm/i1lVxSdFJZmmfxQt30VogWz3NTNNN
dURDuR3WGwfVUTYs2r/glzky+n61KpvGVsWJksRkxWBWu6bvAB2queX2I34eZtZFaVX5NN32Qt6R
VmJaS/ur6kbRKCuo6zMWr9Rv62bSMbUgDALIewL7Z9CdLBzzYHTCSSaJUgphfeOwANEUg2HSA7Uk
Cw1TJtifTVzFqSuiGjJWZE4C2X8fhuX/bGj3QeReitjIgBAIz7xOgeTfol8HADlwrAoFwY3LHFfd
Z5BCRXFf9kPQcCc2CUZOqJinxkND1ftNtdNwaMzIumqjAnpP2vJ89S6ygVIG3UoLXtEnNq7asnbi
nT76k8HDAX3FvgsGCKbV1cmw6fgHsm1c5ae2GzMfFwlqZJF/+JUZqt/y75MkbU8X/5qLr4MRKRg7
6/zOIaFX3MzaVb6o7x+eS30eYiRdfXF2FHl5Nv35K7dsglCG6QdcT8QIR+2sSz1UJ0AgGUIv1lwz
T5G/XGIlmTrfEPUcUqEdd+flab3k0VTd4ETCn2T7nR+MdbF3ugEVVnfFP+u/vQ5QSxX8R2gZlSDf
Pit/NGdtk1q6QbeFGELpk4hUOIRQRrCVIQLjtShkfgpCtBoZCxPU4RtkEvTMEUYz+4z632H4Y1bw
CxOMLXho0Q7Z4HfUQ0cay4zYdXAqygaaXnA14BWN6caYN+eX8gI6VQpxDp58iTa+UG7Hi172T2gD
LqrVio9piRQVzE3qSPtcjc5Z3BjOmTCweKVDsUUdUeqViKEME2Cx8xpTI05sB3WpAoKBoOvfhL2x
bE/s0sbfUHq7GBeH+UwuHm1a2dMs+d5KvDgLHVvKKInmmxRTP8HNOemlKoCkPuYepE0tiTmc71Dm
9SvI4gFmS/vYeQafRp22SUARt8Cmv5PtSGBdyEKf3Irm7ITZNxnXC8HUk3mCJXgBB7DsV89SQwda
troWQzrxsT++zQFTgO4WZ9csPXKCjqYXaqHNpU06lJDo+eIcKZqntELzfbrlMw0A8LuNd3osN7aV
XyGsvDBpAtxZC6CM69LA8CYdyMqz5wqHQJdzZsxzwSzFEjFI4iitR35REdeplarM94c/+h/i2xWG
EIe/GnpUN1zbNow/vQelsUuEEkiWSRbB6bhEDbjQstmA6OEzQKKvW0WiWXMfDfAHfomSyC9raoh7
+soxUZoczfdTC7CjZnEFyk/o6Rpmz2QWsZOrHHoN8osd/Vhb0uyLCYgSUKj2HPGkLYq1Nd1z0/JM
mbjAq9DMlQAVX2KYHlKdpmJxhq2XUXF9GbNbtul4SKx8zAv292DXgLjyC9+IVCK0JPBKUxwVg0I8
n64ux8CD+lvQXQ+8EhfgTmEX6aBUdOg01u37IcIiU6K3NQlgmsNcdf68+OhFishTDBfIK71kVYmh
ZyLkjH0MPKXaHLfDgoXAaRpQ9P161VbO+zfwAWrJllWRtw5b6oWInNLcOf9D+qyHgHIuiCCyn4Wm
iatGcy8BT+4JDpbQ9cjF2G3nzaRNgxdH7F6aW+X+OnJYdDxWnaXSagK5iRZbzXRGxJdYqgzl/9hP
sjkCYXV+8j4BHJqkqVQ1zcjpdE5lDloK73omfDPZU1cp+jRqGnHr3MqS/zL+u6dNrbQmQLyuZfbd
bnqW7NTspsT252NNX2Wsult/dGO0V+J6N/AcQpRLZfOFdYs9ls3sqozR7jyG4LXcbJ0uxWjVbk3t
g3tXskWilBMdVPk26YUg0yrhTzQpKF3MwfZ5g7WWOPm/txDDlqygpe7n7KdiSFgiJTgqLDHLhzxq
aqrHJCzsL/FZl6q13UQZMxHs2705uJaWJEfY00/klZlVKUhVb3EzIG3/GWR3YLyzBKIeFDZULtGX
STBNqfFrP+1elCCbxqThyhRsr1Y46liUFU+mslJBql5GlffsOQxwM3fJ/kwTNVqsgivsrfym3PfF
WwLdNks/r/W/FP5siJ2eEy/XqOseh1Sdja1JMRCL/ufy9Nq+eG35fqGfcH+ZmpGOAp9GITjybjdW
flmPnl+8qrc/Ae7qOYjclz31sgPeMvtnjwLdj61rv+Z2Op1/BGPfch/nIhem+rIhDIeLlyjH/0Rv
gpV6g0vlU+zea4atxUgcJITKOaIbz9nUzPaCPCO2EirsTZLflOurQlHmRMxdM1g5FJ8Fi1FZe66O
tZNMzrp+9ZWW6e4azpTJEIlhU/9UWTpjLxuNkjLfReJj2+o0HTaNVazKiiILDyUbHAer9iK016mj
uDnk1P9fOvTtrY8DqokVRzhWn4TcE68mpS72f0oeQ1wt7hZqts+0qSbIT9Da+8YxnHLwpktex5zF
Sell7us9CDN1fdYagfztAtLDYAbuQ1xU8qvu2+5mgRBa2s/1NU+aumfJOFNJYLd9upskuxiFCqZc
VHoNS685ROXayRpkQlTLA6HVyBCS7u/fuZSMoSkU2S/6lYigvGO1VtSVlEpXGlfAYTJ5cpsY2Yr8
EPEkCu6S89mUABVqgZ8njguLQZsSN+MF3yXVmgJQJgIjQWFiwLXJelUt95F968NuJsuDl36np0Ga
pYW/wAD3Srs2ifQkTd+Y6tTTkQqDH9BDkBlryUW6ex0UKtFTa0RxqClTtZDfPwYRHpTi5Sn+jT/E
T8CU6CKtyan9A8YSz1gfWw6e7zfAlrnN1lkHpUw6Kcl7oH7xzjmD28EqlOYwLl8SXboFy7z0t9Nv
906mkaE20+slsFhPP5iSi+r8ORphhbSoei1DX2wyvjlTQhegHfh0zP64kQRk+FJroHSQZhFpjApT
gwC2a2N7KaGF5MsuZ46lXhJmxcKj/oPwyQqLGvV0e7qPk3MZwXOWJqN6DqI9/0+HHC6DkHr/extf
LvzonLgPycrCPo+0bQ5Z68VXNZKRksfG+Jzi6WVqQXjutmnxJFKvUXAwzu0OqtT7WGEsJt+iwB7q
vA95qU577CrUQq09mP4iapWhI7pqh0KQ1+HCUMiRb81miKYm8eXmCGz2HBcTpZ9BCKZY+XNuGjet
hrd+BMINe68CIS4eqi8gHqVUjt9kvFlP2T6gsqGFjsBpywIFhs42kHlb0/OpYx6dC9zQwlEefF0O
vAZe14bJqwVO2MW5fvSUCSMNF/PpCHndJ9x3I8eL+9Tu23LO94CX8rV9jxnaTQH4pFvJfTgGGp5N
YL6Y/OG5FPW64yRITGcwLCC3YFxmsTA9Zc7VxHbI12jCoexzpBsWb13lrrh+VSDNJMhOHzzGV4Pv
kqmdIRy3BG1Cu0d644tJLnsL0MmEXBZXxrdiNxGLC4Mgl+FMDyLGwd787Lt5CtQLPkC7mLMWazIm
Hprj0EYI/4SfkwqT9f5WbSVir+6QnB0g5kCAhUCnPsavrLtt6VTzAq2h5Nn9Pe0qTXuwjvtbt27x
zwFS8vc6138jdvlImKHGDSJ2xC8IRBLnJpQ41NVaYS/BXn1rs9CxID0z9rfDEVLsrbzU2fGUUewE
URG3eyu8Ojv9y4ohexIvEce8+6BYlRHQZPQu3ZUaHR65EZdu/2W1+ztR+n3cb+haTDcUvZCTEYQI
jDfubbpfJOY4OGdk01EJuMAR+8mV5mN1d/VFgxeQBX7b+RJAKQ5a5acxeNsLtF1RQNYYvO3ejzJO
s0jveklOHl+pAvMLeG74lps1UFL79l3xbcHL+XFbwYGHTyHHYLuN8YBsZE7jtF3t8X1LijsknH2Q
R9gE/GOJ8pYtj22fIa6a1dhL+OLhiq+UsYL5zXGf7oqd0UDVzkCglJSP0pGDyY9Wl9eS+9MT1zab
YReshqbPGg9BNsmgKqp32TmXyVF1MHiP0ewxJYuu1b/7KwNQO0emXyhhkj3Bh+0SL3wowUd3zlCL
QpofC5OP3NQu5U5NRoyXy6VJ5xxu8oqCP7388gjl38Z0qt2IxI3xdEJMQxBRKmHbqcexBHTNAqMx
N3GJiGkff9Ff/UiSIXV4bkUaErtOiciMO1yY3hZuMZ3mJUZebI9egxWUc6P/RUWUmgRTdNWC7Qm3
/CfP5OyvhSKtBLeIMvQoE/ZJiwvXR0URGIJrB+LMVHbF8QDfCW8w0KNv8qeelwmNKX8rLZUwY9Cm
4roZKfWiTY4xu3HU0qMizGJC6Pw3/tujwrPpARa0RcpjG6WxY/gC8wixaJy7yHD1hny2Omf3tM4/
Cb337zNwY3W1S3mHr8PG/GwJvaoim+kLZYWFz6vK35FAQ17WGw5cQ3aA5c9SpXVEE/EyuXu+zjX8
QuzRCZIugHNlINfpiNkjjcyYBBOJEXJuHTNejpNgzrkYcPbpTOdf8/xWotau9+6UmQtTaWHQSDE2
eVWdchIfNa4TII7Dab6FvQIdMTNsUaD7+eDH/s0j0yS07XP34kZ+gTf4cE1VTcectwKesRNm8FpQ
i0L/gJc6r6MmzQTFlpeweL42A4PMZHftYePGT0A5xmnHI++3lowKUFX2W2VkvfGe07hE8LQAU2sR
XPwJSSyprhea80X4QsQ97sDgxtQS/qmOOuI/zrJr3IzZlnOh+rYuQVwvSemhpkSLZrPzr0AAqUoP
MSHnPSYz9S3b7Wm7ZxnmpHKlvlSIzLTgBfT1hhUUtfQHnwfRhaMPCNMkQFfZoZeOSUw1Nhafb93j
AMrgycC0t9hW1wAw2XtBGaRt2EzrG3ZgMdyHq8T4G4iEGbawf9Eiehrokxr3B2Z8x2UpdIJvZm1q
X015sfvLtjh3nthY2Euln04sjezwvk813IqXgIfebmAsff3hL44H5Zu8GDH+jhtX7SbZ21GneTvb
QGy5EeiLMVdhnBxVoU8/Repe8pvV4vtVWq9tXFmZ5QcglubTUSidLdi0AmNfh9KUT2k08s3aiQVE
fQPeX9Sb8Bcm7ONhByx2Ltq+jrDNH44YzHDbFejXy5JrYGKHTm4SgncTCnISMiLwwXd/4IKUbs+U
sMHhiuvS+N79TAQ6z+PiB+UGOEDy+pCsmj//1ckVQP3pg4hqmbQtB/uis87buZf8o6bqxE4bp5yx
tWbwcAX2zpL00s07diRK5FNiiRDPrjxGMEJQs6wGHKXkp7YFspE+Zf8HhpfQOC2+gG2PRe432zQc
J0imW1MJNyum2uS80iMTJxBjf8WI1wDQAoy/jBnJzC2v44yyNvnHUb1SR0PDGCu28iya5Na341O7
EKcdUkAIU6aMpEow5FvieMRY3BmzaJUdq4ap1LHTNN61hZU4uGKzl3sz/o95pPLnmReTnfsnU/st
RsOG1d1iCjPArHgsRE86YdI8BjE+NQ5SwRKaI1VUO77CzrfLurAPrP14P8kfgir1GqUvdhNrWRX3
zZoXWRan1prr9XTdQQOiGnVpiVbSOfo9pFP+tYB69kMhIUYvpnYQclbXMGdZlbGmIaQtYWVWvD62
8gJG1MHPo0El0cXGQRV4iHVQOixVrwV7kuubchkr/rge3ZRwq2w5IccDSgD/Wsbt/IJXxUV95xnT
Dg1oAf/rP/XXYviC2gnieW6lzqyVm1xAfjwjkDwal4vjSC9P7IEeBTzmRLkCPH9+LWaiNgurc8Yy
iMPvpalFG5IFH8/SnWm66iFpwHYwIPHLuQlNeoYS34RHBjwD0kqyfEMGighZGKp88d5+2S1mySnS
vUFJNyt92AfiZ2NFaZpvqMogP++9Zf/vrLxRj89Kw9dBmdhrZ3GieAfG3h5ERucDOu8kJ8J4CEK7
hPsSLI38FFv61zIhXPNTyLF9p85p1H3D4XDyZplmJcQClSLj3mwMBYyMdeue1wO1jVioOJ0gTBHM
x1ijNQCxqpl+oJeBcatsJY+DDRwJ8K7pMQMULC7Coja50d3U+EdYzae24AKqH1QfM1eZMlfBvnzm
8Srs5T+36Kq8moi4ckPJqfszaserMz4mxBLWWGjkXlESB3dMoyjHxJCqPYARJaYkuLSAlaPuhPPS
qmt5o6im+uCSsa4QhuoJyRkRfTmCK1lWBrf3CNq/NTpl2zOn8AgsI8rN4LBAwLYHj8xl74uPJLGe
+nhtyj4gj0myAtIxEQriMfqcai5QmyfJ8GNAb7mCcT3yxyZTnb2H74OUfg7H3Yew1aAVv0vc/PUD
4K4x9LKFZolGX1sYEFtbPBARhSU6GLO6FMqQRMU4ENNVRCTjN6mgE2UKjjF2RWATo82oaRtqQAg8
6OUtmfTj6PxiFW6fyUaTpfJ3I/6O2vvnxoMSSLoezuyJ/02GkRWwAJPWKFr39Rg7U96CCP5kGsqc
b6vZAIFwdIbZ9F0jZctEw1uf0oNWwv5ce0xkLnvBFv5TCQnUFQQBHjfOINrcHAsl9ndQz3p8QvFQ
wJVQkZZWX0z/t7hBfb/5geEPje6rU7r8W50DE0ZicXd0cAmTlmRsZrysVJPrTY5H0d1UE0BKachZ
rOIZ3WEFHy5XAJlfA2CTzEQdghdkApag6Tx0vWdVGJpzEs9ETKki0lOlFGaXvY9efpMz110xOYhx
ELmangG7C/F5ZXgB7yyLNZQnzj0zQz3oRC9BXyUmfw3mZx9ROAyWox7/+IW5z4Vo1DezSX0vaDei
P8dQxdDkmXr2xsJzAV79qELr0KDiHvsSx+juMI9xl/OdJhzWjRFaH9BNqk6/v91RNUWOrEKiazge
H2OhYouoAWhdeG4pAE/myqPmezusPfKCADirFkdTuPTFz2/xYiCH7JjdtEkoYc6PC2fALf/F+ItE
fIZpXYtwuE4GJLzMmk8hnAM5TJXVdJ/KcAEOCBKuUbU1ZI15H5yAF447Q4iOjoZjy7+2A07jdH07
TjqOXiiwXKQOXijSqLsJhj+EE7obnRtSmY0V4ZX/VY4crNggRJ8pEH9hHHD5thB9EVCnkoyI9g9F
1EYpD3DtOunMeO6SBkop+6GNWaBXY8/G4y9MS/Kg02PE0DNAXhK1vgg9FntKofDTWc+kP7iVQLwQ
1gyw0SBEf0uGe78uiO289ijQNzHTQ9deX8sUfVQuO0NVTsIWgp7RE2B9WAvbZYwRItGFpxnVQhnC
vgE6hCO4WDJS9wrQ2c2+h6jpXiXxs1CtkCuR8lV6bJYhgHP9sMj+43h+CjgnoFwOcc/gNry3rbsR
vdCqKdKMIf1+rzZHkA9jT3cUjcEijhGkANoKG0aXE/+woMnKSyKYYUPbq3JzVorbiD/5ZI3DFtGr
ELp2t2wp5Rb7R3hE35bdLA5zKjBj3JdxtOYl5pXH6RlKOjn5yc0ODhTTcAoaI+mrvBbUmo/Vy6N1
wrdhtT5o9fJoRFQsMgM4fcvwaB8Q/ATyQzNAXMe0AZwTPTQh7i1XVehOHOHwLMt4l2fQzVWiT69B
vttLzkxDJjlpt1y0jgqsEmwu78ltgJfHU3Z+o8E2XPyhFqH26nB97YgKZsoFEZ7duqey1Pqi/vNd
6TU2K0JTxkq16+itg4tTp8NMvZweO0Cd77cKjgrnxLpfXJaNbLIqLCRQIgCCXBgwDj99nqBn7Agu
O9Ai1gPMJmqGFdphbfUz3t8m5cTQcP3gY97qELK8Wu9WbeM6TixSm95r5zt6Udn0ThYCAu1CvlS8
bpKwW7j8JwgvT3knqtQgXxtH+48J4nN6DUWoarMnbOc81XvOmauZhGh1HtKebytNEZPSCMnyYRzV
r3N+fL2gb0o+9hL/MkTz/mIbMO+UholgamFOD7tqKGrhvQxH4NtOE/PAWWZDMINm4GwDtqYGEreR
pcIlRV90hmAfkp66wmwvD5kNSIGFJZpWSCDTztY5y5ix1Jvax/AF6/cOhLJFUdT1Os5Kg3cZaeXl
2p5tg2JoqQPq3K+nKvg/pSaZrsI2ptUQPxGKH3vEETwT9/FnllXLyuXAjMXZHPowIREKN716uWVT
lIk660oQx6PKoOpI+I8bHPrujc97i7Zk/yFNix6blW5pRTKPPcsbrTIvUs3Wws+vSqB8WTAASrQz
aHyvlvxnVS25a+fnLUQsIHesOG//ZneJwsw2GafAxMAaNY9qbUXbzXvby98ptywcHArXnKfdVWTq
a8eJ8D9vo/4cMdA5ICuk3jHH56XKZdeT5RITZvXu7JK0r6lqVaa8RXHqKjktcfNwOhau0MZ2qI6G
iWp00WtwkasER75a1BaNYzw/Fpc/CKqevLk63NDGjUKAxgSrz2M0XkAS5xvHkbkLAlE6c+YCh2Me
KSDbnaL1T+A25DeMwk21aUZGOOF/re0JlWhAJCIQ8x3pqizyZ6Cf5uPBBrqoeM0oniOf6/A/xF4I
jRGk7U5u96hwOWKAjdVN0GSKd4P8sHHaXFmv5fRl8bowaJGiaWIXq4OvkinWcKT2vQsSK5mIY3g6
hskN1Fh8gAwRT/S3DOx+RqhtpDjho5zi/nxSqCUsAVujkQtQfCCjsmYx+Znm5X2frJsqf05uu2fl
Za9oaDpVXG885wdyExQciS8tc+jEJCEurzPG613HHm/0/WgLTmjwkHwnryWfRH1W+SXrSWpcS4rv
qDEVHMfJ/LAKJfazQGHCFxq4hA4EMD6AUozM81N8hD233L5AhStTiUMYyN5qt7n9kVYVP6yVVCdB
Ixi4nQkzWx8znruTlfWC8lWiKoorTCvwZ9xZV7ZI9BigLyElABOFJeMHH7dZuME2KueQtD65Hpgu
vCCh5+OY2Zlz0NximzeuPtu4AGWytPZZVys5OpEbALrooHmknl+i8FEsE7m5Tuft/6/jBHXTEDQU
PaxSlBUfq+xZ1c2XA1JUIpIeeXDJEBieQnIJmLCCuzI62DNwdlFQ0i5RaiUJ5RnA+XX/hK+6YzOu
vxBk6nmMbiEYCtj+jZYJRg68KC3eESSiVrdzYycTdQS4EuZH3ctfKJxvvBFB2exXtj2VJVu7KDss
RvUA9CirCjYv9+ZLihJ6tDUs7VzaYt3/FFWO92mUlVudPuYgTtrkM5hLY0lFvY+hsfBQ6vELXj8X
T99Y7N/AKI7aEqgcx/azGHNHONthGaY6OASr8HIUehbwG18W44h68/Vbe5Zscx+B8blhq2B+1iYw
v7243fY+mkaxRVvQ7yBVz6KetBbekyZnRaPJEVeTXO9X0xdVtf8ncZigXfsNnP//zg2VjpMA0aHQ
sEEg8umsmxV9PC7okq7LAGB42T6VBpQzbS8XqLVWZ24QtzwEv/yXajxm2sZjvnuzL0v9ZFc8xVEC
IwsaPLxqT3QyokZGvnn+WdRgyklMLiG16FRJMptYxNQPtl99+uUwc97jYbLr27ARg1hOMh9jDaV5
zXdTZaIgCkQUnr8hTqtT8t2cfmlx7FOC+0vkTh2AiBgXQ8sXGYO3o7xpTbHKKWuR9akGPeKWwsME
RfVXZAnsFtwPE9/1N+t4igT/S77zcRHVz8SbyzgWWgx2uxlZ/CTd+N0N5pczHmlAxUAJD23cUnGy
DiCMHTFy1CmkCpM2lwrtCooMxaL+igEHAU4P1+EzkHjry+8jsmtfxoUCIPLzcL1Ial5byJTDKW0f
y4m6STunrTvshJQNrR5Yv3cTir/lZFBxaYA3rrKvZo6WoCzvKnJz2EfFYrmXzriq+vRu3+fYOH7E
cOnu+9XwL1oKznikeCKiJJDfDh62c+lIwmo7J8fyjwRxEGDsMYyZWiVpBX5mLrIVYkFWldq99N5p
xELmDyDu+TzejGE2xH3rB0CRQKiX0xZljZX+iVpqQDVXly7AJ1zA/D3Ls82Ky3fZwJMDOGHQ3NDk
oPH6KHvjAcwu7Y9xDZep5fR9fwG3M9TS3nOL1sdnw7amnkYNHLbsAasaO8t+WzwnU0+iBv+0CnSa
A0+Rt83I+lvyBbATFOADXOf7+CO97RoclW3x9DjtZ/9xI+8ibCZGCEN+Wq5WBje62lJjWKQ65KIW
VRyChSiudQgfUXLLX8oTNpyHZ8JEwvfqNpYVG1APxsVlQ+/5ycydc7W5oLnobtBNu1/MB0MUpW54
rhBt7wZ5EgNf86st+hJTj6ESkfZjJaPxmPf0i4127MWUwayEmv1qm9uXeSWyV5LcSB5L/y0V0cxL
+VlXkwVNYjQ7nBpLz5IthV1ghDdQau1kWlsuv57PCY/q0kYN/nzPpFbFO9ac/7ovXYmXC/5MxsJX
JiMGI6jFgaXLVVmhYlRGd2/1UEGysPcnTdUFzLOiQZIv9wSZvQTtS7pmVaFzeqiesHykGmE0tFb/
dLGO0rejLQX/s7LW4m2BTMdvTLD6/4mM/J5M8WW4FTHdKLHVc5TATmpvmyq/hHzb0RTsTrm7R29X
F8565N6ma6VfCBC7VxYNJW+wMXFKNRlJ+Pdj1tU0DYp/H8COgjAFDvTTMA/qcEJTf9jx622EfRyP
fHQ+dBYvAx/KtE5c3ONSyfKH71LNDKYP++fP5GzTZR8MhOPr07nJC9F1Ke8zAuHVWRKf4F7xZFvK
54GJ+48MC2srRyua5WD2x54fGmtz8udXV7K/uPY2vZNCshRTh1WgX9juvD3N0cmbL6tQ8gWt1z8I
eq8yI2WiEZb08erWUjARNXvDV+6KJ37xqiIUwnDeyjcEi8T7CeF+V3Q6K1vmVU5OuxEKwmKXwkoI
kHbAx8xVkRprIPhLGtPTUaMVg7J2Nrd99TNOkCgtArfoUm2gZG0UCdHam2QTkU408G8tHA/4OEOx
r6XMXE2sbbxmw20hPg4sCrZJx4O5d+Jpd+Q6BRUcnpdeUAZmpq37vKH7KWWb3uAL5n8WTphwJPTa
xsO70kvaqqfHuVoPfV5VSUnM/emNwDsWMVXiliYX61imGCuGQy+uUQt5v3VzL3/rZe9VSwDO21BK
Vdeb2WvI3N2DE9CnUzsqDPvDrko3t//W57qAlWBMVmgNrJkUe78x400NEh8b63nkjB67CXrOTv3K
vvGqELXAGpu8ViIQR3PesZBJyCVR1MGA55eZY8c/ckBD1UVcc2OTBannv+1VYs31og97k3GBAt/I
eh0GBn4jnvz3Yk1rQTg0yytF+WwDSCYR289QPITyDqcjT/C1NvFnRM5GxdgCj7UjC8DRQkJPo8kZ
3cw0icV5ToER91I3FBWaTQS0IRO/wRKPDfu7YAykAbSHkCSSphs+3s7SVry/yRG/kUtkL/0swS3R
SGqu5+MUWdiRJPeR5HEhJLxV5jeM/8u7qf3tsPrdKP358LCGEv99R5wzmeWQIbN9sLLExDIksi/B
gR/l8o7lEQtGdBFGscdTSKdybba5csJCE+f/kcaK9P/eNWYB75YaIu2l7zYU/Lisf6n2UbehPu2D
mM1zBggHiu9kGII20BXgsNNBFIIJzsEqtbs3N82JxcU62I3qMf0llR5wHC9OTia0gHdQWdgfohjv
ko0bd6ZQ9pWnkiVM1EUKQj/PGmsD8fY1VA5gYBshpL4+wtCq9C3fNbekATb5Tmk4DgYppnsmJ17N
eh0xNodJS4JM0qGuZHLC9NxjuGEDWWnbja99HK4sQ8Z1zQRIYdz30WWqP/SDpljtnuN5juDuvPte
j1Gg/qtTCjHhFZAQLaSll2LeGYZsHq+gV1EKJEASRm5fMhLsajw7OyAlTqN6LthkcH8aD3DR0GaR
t/JmtrFdq/Czf0u9JbLyNX68h9uyvkYo0QrKBalH5OR9edm1D2yFQsG3mfF1qwWLG4XsZDflGMRf
WI4ROQvempQ3Ux9DL0dhPlaTLbN1RZ2Lx9YdOUksu0AXp6DitUkCJjkWkWR45CrDmk/0IE5082Xp
jJMCfFZqVQf7yNhM2KLOixKPe77lXJoSiWnJ9Ur/qbRNI6ez04q9oZWKK+kmRq0KOPZaQTSZZxF/
iZLDuRilC63Acx/MRMatrb06F/AkyGg1aZBR5JYgcAMnKWpouXejVMFzIcxzKCH9zE9+LmhNuoVr
lub5M92prz+ODuFhxl8bm5ZwinlfanraOD4UGC4Q9ZXQbd0iSDxI7XJqkAQOGIXnE5bBAiUMejSv
8zXz7q8wixi9HlJebkjfcrK50id8EdtTbiof+cQaJUYA+quf7ivIC7DqJ4CWkXEwrfHI4bdH7IPu
rdAxNuBwggY01j1CTxb4DoGVF4Zob1UDrNfa8iWX7j+E/EIeFnKnRYHhLX1kmrxC6UYdNYgynU47
V9KJLdly9wpt1I/nc7bG6NNXxI23p8TF51CTa2Pe7n9D6hQztSBcUYpEMcyAEeDXxeB9XzDZi1H2
ZnZrCzgX2au9LluPnhP7zh5Q6+Nhdfay/ZfoAOdAAR0bkDpxhHLVeJRaZy5iIljhopbWzKVxzCyW
lcMaKeBqjk2ROPd80oVv1XQw4dVK3CMOAoMP2vdI7G+qWcDS4b6OTVwZ7ny56lfiUK3CtTOqnAs3
S8+0rUb4VAsy6F2lGa//3K16MMQxG2flHbw0q77sbJrib1fYNAA2CfeyDYzk31/xB2cBiBQTfiOS
i7FNDirASYMeMhjOPvJC1ig8MAKMd4ed5SL9Pmc1dSZIzEcjBTndlbjmLkKmwk9DucexhE2QCxNj
ry42b/yURCJTo+Q39vFWfaZn/XegwldMAzmuCFXjofAW+nJ/jNQF1w+eHfs6wVLGl3/zeqMWs4ce
7Y6zzK5kggZTFAvlFkM7vm2KXLfdg8l6+bMzEy9vvk+CxMHg3Umja/xiPDdVuEx9us0U+NABEHH4
ol3Xbwebudr2sTn4fiKG181tgTtZG5zIqZ90EKcIZ8hAId91LYCRyzyYJnvcOzcAvJ6Juvl6DGVA
5zNpieljcheiFsTXbKgDZlz5fhwUDJZ9DNOQkLfjohr+1nC8QZtP/7y/m65RNhbvXDoVdJadgNP1
SLkYJDpzCcRQfRZz7o8m9a6StkPvK7QdjfoilbHX4bSTYnOgqj8kg7GrFpz4KCnzBKWd1wUkLIRJ
cCubx6WOXvVo2WTpaJjC/oxYuSgtBIlqQW9Riedgb3DC+49eCwpBuqr10fW38xuHGcYiGIKLk//I
t23yEoWuD2RIGRdBIQZdipmvJ/YpVSjLDiODylBbMVPAsddGkeHFN9W7TWqsPgMvneqDYdcZmVBs
+IeZcwzaaOWz6QJXhmqdW08P52KSJ5xasW20FF0970+RtpVR3C52pVVxbYrYQ3DzKO//87OiQ8RW
7o1K9a1xdcW2y6iyIzt45Tt5eXqZgLqYGMKTUJvhruqP0kKMSEx9U1IwQa5TGalx0+VjopovTZdZ
DNjvH13yzCIEcb0wasO26B+SYhJdgexCzouiBlnd0nhjLrHiFJ2MV7+7/uxtopMBx6Xo6eU2V6JN
Nt2aJlMoHoikZjDZR7c+o50LvrFWSqSzoGcL18ttpKKposbSHYntcyCzehvI+61smGrZzGvSRACL
n5qssVbVyvRcAEWfeHeE8Q3dPVp4kPEFKsP2QyXs4Ks4valBLCZEFBPwiHyOQazlniuEcIfb1Z0s
5a6Tz1RjyDbpnyE8nwuNwFqgMFQiTogeJNegKF27ODZoA4mZRzp1CNdbVJVAzwq1rHMWUIn0Zpub
bM+E5jO/IEas51pslmQv3kFDvgu0I9++t2o898XJphpSarvo2d9wSx1I76U1se+mZkQCPxdbPmTl
4QHhGnF0vN4MRZUcIH2xnNp9m+6CWnMvgOLFDrz1WwPy0G9uUb+is8ToWpKPi88OZn70OlTDBWCZ
kdM5RjiEtV1glMX4LU50NPILM0Hg+CNITMLNDcazWxkgbJBNxyl+lpP9Z0yZxPGRQ48mv/km7XKi
mucLBLO62J/ObWhSRfgJKyXbzrLYe6+N/IBlx17EPrBdAF16ZRx5uflgBLek5Qc/c+uBiecuefEi
kLEV2DgjoZ+jPEfrw3cmtYfCRu8fLeLvXDsRdeSVJ68CrTV/K/LhvUYhyOTvMTheWoz6wTZcptXo
V5DcdirytlNZe/Ik3rNDlBeHASKVMdsLCvXleb4NHUQTvb2FZ3FYXmpfdSRGllNR9WAHOpay7d07
m0D4hqaafy7XhDfg+uO3a64ZpOnx52JoFaOCOW7dT0tOLTxoJL/014B+sYEtRfTGU5yQ63p8WRDo
U26pExbY7A1isqdaVqWt9cTU/HgN92nD9bAadIrXhXtnBlHDerkcS9nJcuR1ip7Vm70KiZ/CZ3F0
814qijT4jYPNxnaihGzpTNe33c6vASp8tpUbV02milHA0Zv36C+FLl7vPtSZX/a7h7OKA0ZpJVmT
tdHyID7sUNji7caew7ojmDHiAKHfNF/nL9GQXCGViZD8QGL75KjU6nXC+RzYDm1UsomlCIpOlclD
IAI0T7N0qKSUJBE10YZ6WeS6QFksmwXhlbsMuUruTkRozBcYTmM0bMe9fE6D5+hX4NxI2eiQwtjh
1oLkJY/4dDRZnfyj1YyBtsPUGnnngq744b22sqIlcGxtNluZXWpn7eNKK8sWpqxwDtLPjuKqDPKK
hAnmbp0J/F8qhakdnZlGoBL/hMaqG7+JcepvbdUy7nsIuyLlyAqqZPTbpD7aG6REhi4uTTDmH9Ma
jtDRjVZQQiVFVpYLXon7++6zAPQk/NfNm/y80/AO4Ez/RfMb+AgAQNhS0FOJtfQeGcjdym73EKLF
WQkQpCKa7AbuVZqSA1MzMPrBWbko0i7g4Kid64Uv/+xMOkOJCjy068bX12VzGKjKO6MimNybjTz8
CIiN8AT/ukYXsFJ+qwCxQDc8aA3V2ZCbYb6fsapSgyLzFr9YE15y0B+Un9A2nfmLPCnNqSt3QXhd
IKi6MK3cWoMHHOG4wnKa0RRRJOyMrIAojDPqaeZXWfsuHFcrdaWjxF4Z/m6kMblv0m+Qoel088uF
amx9Z7cIlzh2g4FmyQKKQw/ibX/RoojmqMCF8U9+5is3fwNdaTlbwesC8NT65lMfr7ixkh6BZDYH
0My9deduaJetIWCRX5OGmlOCQGlRNgsV+tdIBUvsAmcVEDsyMisby5cvz+Tk7L5I3gsLWo0VIcbw
unGyFwY23B+EXQ46d3TtPiNHFLaZ1aaXDQJ8kfLuZdJR8mdrhj4wIM9AS72gBR984vriUOGDWIk8
jW25Ixq43hucalkAk6e0X0EzjKn+d3ZwZpCjLvQbRgf2JHb7FRcaPJ3N4LfScFLdEkQmkiTIdkKY
D2RrRdzxdseGEnonebDgKglGon4Ufd5D8CSQw6bcdklE/eSjqSIPyf0YKE3yrp6Tu608e1CFEvs0
SC8JZ7/y2c/AzmXVmBoHpBdFcDuzYC2PazDUs6tgtUT+2m2amE1diULEeRSZYdOwnKYCA9+NQ5fG
AASlvkKlHohObbkPcwJWqFq4aglKrGPB1V3iX+dzlES4i/PSDHxshP7lAop9byPSOy9ASHZnRqsX
Q7O93NZOuP7TyKNx/gYRLDu/tpFq8qQXKfheSGIEJ/QXQnunvq5s/iiXY1muMU5tWUsid3pFVFeW
IZBw8+OegzrK7rgnZzBr3H/nvvx8DDCFw4+kqGI6ST1fYy735GzaJGtM
`protect end_protected
