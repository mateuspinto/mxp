`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3088)
`protect data_block
+KhFLhd3coUIq6+p3P8BGk4KRaQHn6YXJOziNr8UeSs8r20EKcbbF46TumClR29cY9Iqasf3ckEm
6+TwtHrtlIECXrzKUIB9TPMPkciXfeKtplY1IMISYoIsuHjrQH/pBbLvAWTYv5R5NeIAyet09oNB
Qqw/r3k8CiHTBJnT2Myn7ZUd36BCFHwWMBhnZUtjylu2CphBYv5TkpHaUUROvOD1RSxy7izbTxgn
vrc/y53Y5+69WPgn+wO5bD1EteYKl4qtpSmaMR+hUd7/CuZtZcyRiBhKvWC0TCnCGeBPSmrwg/FT
2n0U06GgWgp9jr/puoAbjSRVSOthi/Z7/AErIKD5dSfHHfxlWzFzuNK+N5uzDSGW2zROCNDG8Epc
vK2dCRhlfe9aZhom4XZJL/Oh9IScnHiuNMQt+NiRiPt5E93QvuY5TEhKkUp9CW+NEc2jKiiVWwgq
LxG8+UP5mncPnmIxTlpbqBzFJ5JxKVX+8rjwbKJGD2qzaFq7BZvsbou/o8iBYwwjBvS6Vtbf6p4z
SorkW0EXWBIBxfjG09J5IBJ8bncL79RNjU1REz07VWWy1dUdpydwBQoiGr1T6AiqEck2G967xiO1
NAZLqE8r6qtKlzauEVBSOhAUQ43ktWxqDEUztIbgldwNGZlfrBUs4KhXrlJg7J+ERJPWhTzdyEHx
VUcwrCBpWOpWtupEnC+cwC9TetXqpRkFMl1yozWIaRtx/3zHhHOezHCeQ4+wkRzko5vD+7bIS8uP
dci74IvDoRHLwa2tcVO3y/3Gm1DA5qnYjVgCg2vuunYnOlMzGb9i9KBfdTvRqOeQ4Zh2k9OEmIxc
crwd05whNdN5B2I3PgsZHwe1+/ufs+42Pv20y5J8bf7qeKmjxLYKTgYTZvoWI/9QMaVzZKicTh3N
m/kqF5hs+rI+3Ryy1TuGmHzlqei0uk6NXqGEiboU8+WiN/fzetpw2KYuc2QKAzKWfgR5hCQodSIz
qgBSvyL3HuLmNNVTqNZXnhHR98/75bDea+nVEt7iMrCNjlstyMfKiSsosTkaV+IqSasr890VOli/
9owmZ6Ube3dXMHd6XD9h/DIJNhZ27xQSnRiYlLto00t3AbzOakNxo2eJHMbluDATk3sx4zzFHM/6
8n4HrUtZrPt4Mh2ujCiZ9TDlpi1abeMwGnLXubIlHWNeL7Z1v76SKyjiMwggCvgCnzDijWsCSIte
U42VroN4P1j7A4MB8v3iQTVF/SGOYHs6kiDmeOtjC99m1Pvdxgpyg1tpPu7QagPjEPlSF45iDBeO
xderObek2kDIQGfCX1ngQ0WgSguXwwbgJYjqbhgAsp/+UXr7+HG5SuVy2HgFYWj35jx/UrqxT6Xl
zKLBQSG6FpWHx6AX+w4pgNKRl+ga0Q4Nv50GHfzHyDwBR29f4a1q0qO33sTAzRnL8xmBmnCXVBoe
032ReYJ2nUNSF285U3m43xBFO3lNr6iZiVcg2vUfdYN6hXqXOsxQHR3cZW5Le8w+sCrvdRoozZ88
DaAXP1EzELXHkdjo1Lrv2O1vN/JeaZeSb/vD2MMxNT5+TgpdfetjiDFHWYmMfJZJrAuF0hePoLQr
IGnIo9hhJOBdSuSmlKCmPEbro+sbrcNU61C8yLZZ463Z7eF5LFQfGGcpFCUGSH2HrIiwSqFDl2Eq
lAfBY4cLjmCPKhnALLRNuRK7X6X25LIugevt/IzFn3y1gfqgwkyTWSQfwK9VEjx/ImvYM4Fi4xh+
ximUiDzsGzPqs53ErxTM1XyAwQ9JDK4O86AgZHEbtepDHRMplNvqcvCauYMbz4aRzPcQXr2IXcIP
HttB9yENpCD/vxduvNvP0WlAVRdUQsfsdt4WS1uvVY+gG/5nDce0lJ3WrOkpQtmZP9AuWCcmNe8o
NQ4V7jQakrD8iPzaOQI78rxydmtAWlX2M9HKMQY53xZAoWCxf6GqfHum2cBNpHKmrLHJTv1F7u29
+TRg/qQfviIAHWf/87TUKhiYm7ra+HWzznVFauGdxwVGlHmIFiWoWTY8GcZUMLRX1KE/UADXIL0E
EhALNYGsW0Ba0jLsDxkNnds48P8DMdZKplHxORLnFzgvhHN24Z1VVsGPAesyehhAQhyRkNGi9CmM
jrymyM1H/plfbagVN9XDVCxz7Rqrnuc5EN7ZhvhGlIx+ftsfv/iiE5b+TeMxy0qBQKR4xWgFLhoE
/OG78cL0B5JTKEGFOmmksjF1KRHywPcjXz1TPXL/3o5q9dtw1cLT3rP7gLf4lOQFsGmF/dwxyc8N
qgPajoCAm5xc34vIaZuz83o3voPdZ6y0EwZrHq6PNjVajPOx72a3uMy6ISxSVZwYfWeYmP5R1FJp
e3BdmTVK64bwR+mZvRh0thaQ+sWAHBa8JWF7HCU3ucg4lGuzgNbxaFqThhEqyQImyd6DfVFXf1hg
+udxTwWSOMVcTRscXdvz2o9fAwvf2KCe9Rr6ZkarirEfUi6BMdc3VLRkicdofJVz8WgWMKTxL96n
dtdBNl2h60ZqIj0X+XNKAT2hs2eDvMzkUpYOOoO/08fg8CtqD2jB6+SlNcE90kt39lcDUL4TcFjr
pQ8v48WsXI+S+MsqZG08hjr6YLqXG2J3hq7UMTbofCdzMXkIBK3XaiyyWHD6uQm6HXsa4m0OH9UI
Y/InenPVT7UVgGTaKn08OndUywAPDgkD+26zVdOo6YJrixReUY64UotvRxO+lc0adbosMZdNFfht
qbTIJ75DEgDJOpcujbxt7jm0mD1lFnDsdfTpPWXDq95HxL9Is7hlIGbBvEDRseoGTMWy7amWL6PX
byPbjSJW73EfOVBLZXOkWykb0dZDRwtVp/cFH3GmksX/qp2WJY5xyKK02dlNRX7nCM7YkvAIOxeK
21osB+rs11oilcRdDTaZ12BGtkd5U+l1LpCljmPdmXWU5CKwam7yyUONYGZvmDtrdLLVc4kTynKO
LZZ5HwU7tmOYri6Ri3+j3LYqTjbB7p8A2ggzq98uAEWrSjGdSqB1JLhQ/tirhqY0jBvsW49F2eek
/aopDPnm6d92iXUc83b8Hfr7/2Nw3WowiXO++YQo3AtKlXZ+JuMPd4vT6pg/zZ33RY1qduAEiVTb
n+Ls64LogT3xUruPkeBTJKs2K+v/NDDlOgx6zPX620qmMs0CIoaX88eJXy+8+EUc0ArMLSxifqrG
6sXqTZChekB4bXLno8H44nvdlmv84hJK1NuRBhhyPLQbTjxdBhNItRE/nrtyhRfHbgeeXuB7orKg
Ge8Hf21j4mh3J/Ul2LKUpsn/pBItZlEqLsFXQqBui7s5NcQrH9aqGEtjtZc0/1Tt3Ch0LdiEm69/
J+81nVQqm17+U+5kTW92o/+0GLjS6U7R1D71PYve/5R7dPBZaunbwrG2GkLJNDbTlC3ZZwdFyOZn
cUlFdEplqo7md7zJn31Wh/l+e2QDXCiKO5TPienCtFUBjlqhTHxnp6sKgw7sSjMMELqMqIMU9TsL
LXzzBkvpp4SYw2cYT6LmMV8rEtEchsvb+Pz8e0FhgiPDyEvZSCoQ42HQ7JRLH67+aRgyauba44Ii
HT512XlHV3hzZrwACMX+YMlsqQ+illNzLnaYLsKzlmGoBKeOyXy+aCF+es8a112dz3Hm/zCVnepJ
TvEQmotrOGJAZ8stxZB00pHQshqhbrxKxJqczDxmV9asRtrPXiUZ0v5znLg7JF02P0CVLM0p2iDi
l/Km5bSZgD9SnstTD/tU2C+4HqwCfQvBk3+EK6jFiRwrXOIetSYOIkA9kNLT8wiueTb8kiQ8aiUE
bYiwvCisQLCusxcADjNv6MRL0TEcW8q8twxZoCQvPHaWIAGoC7w1rv4BH2bIppGUTjQbT4APgrdV
hEJkdjgU0VYfPCttfi5on/MS8d0CorpSWsqod1hfOEh7AEDkhd2p4/49Zesi+IExt15dpIWJLSEH
hWhr48fWtAd1Y0HUZGyrnxA5W+0rgqdEnsMDfu0BYDRznFJMdSj2OHUJz/ptUVXFHVGhKFrNSEI5
aCN54fvYzEgtipTwFF9VUbKFeHAYWaQKVmMdfjxjFeLcpXRcnw/l8DliD7POXVdr29I3Ck4wMV7Y
GNO+SCbsbeEHOg==
`protect end_protected
