��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l�������	���b(�]o��]1����:pƧ�G��{��Q��0��_�T�ƺ�'���N����p#2����O�!��㚭��ks�<mMUH&��2��!w5a$�0�lSn/}q1*�奨�A���X>`4ģ����'s5}i�3 ��4u�(��g��axkA�#�Z�&�i�Y(���D��&6�E����5���3�M
!��h��7��Z%k���!_�W��$~�b�Y*�vK��I�����DLx��Zx�+񐖂�=(J�Nе?�W
2�K��J��4���v���]�{�{�{�����#\�1榫'�WB�DL�w�<	��}( :.�C�g�I9ن~�c���ܔ�$B�/��)�LlL.��9��RSr��;)/����t�^]�e��2�`�k��}C��K�\d5��J�E��D�M��:
��6櫋�v$�����fE&x���?��D�ToAps&���V��cn|	i�.s�d�pq�)��	�5��m�t�ћ�k1�b��"�v���H$ώ4Z8T 4��h\��gg�J I�9���6������R!�2D-��\	��^u+�C�I�֍��t�3����"�/?���?�N���V9���r���AX)�&�	�}n}�#�����.E+���z�m<��S;�/a<q%����J��O�����(� .wt�!�%va�j��~�N���s�ִ��_F��Y��M� @�f�)��בw��0:baWd�s=@V�;���C�<�e��Bs{���_��i_G�)����B�Fs=h5r��~�B�:��!���B@�������)4����y�V�hm�xMU�s�:5�-k�}p�.��#�$2_�s|4^d�ђ�@��i����ȳA����A������]%�r}b�x��|�Є��R���-��:PPk��W���T���; v8���s�?�io���#�.M�)Գ��un�U����j�Ѭ
3����B�c�l����˜�d���QxM ������o,��V��*6Y�2:�k��� �lLxc�M�U��؁	�.'��w0��[[R�zb�}����_�D���� "̣���0��ՑA���w�R�2��OX�̻v�e��C��fv��[J��NNj�^��n�Ql�(�B^�k��
���jxA���Z�����a����Y�p�p�J��O~S#%�󱁃��h�7av
�)��*�Z�K�-��c��\�ss+�j�3�}Ue\�T�J���4#������ө(W�fZ�)�O�Ej:]��n`��(�Z���7�:�up��	͚�S�(�qJ�m��p��UV�.���{i�b
C��X_�q��
tf|�䦖B�q �;UD�L�@P����� ��Y�}-c���K�A0�v�C���@<