XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��! xj�1�Ws�R��f��1H�`L�`����R[\C�WN��Q�>�\i�{Ne=Y'W�a}����\ �vK��n���4#�.Hh��zB�SH��o�$n/�f�#>�r���Cym[M����a��I(BI���o�k
���K%��ѹ��@\3�kL�C� �b��ꦼ�6C�ذ�i"��V��2l�%
_���i"C�-	�D�����0T9[����s��\�"̻K��������hr�g���]�/�K���mbr[�f�?���i:r�������F:�@�п��P�+��;Z\.rʢ�ۉ��ͭ��BB���="U�j�=H����Ҧ�p�*!���2t��%��^�Z���(xс�k��!�o�H�&4 >��3�#�7��O�����J))���z�tv_k��!�rt��S(Z�y�`�y�*��R��W�.���cOV�-���dq��#����(�P?����zI�������Hw�X�?%cᇨ+�֫�TwH��鮅�E;����=m��WFj�%lG��\�?_����J��YU~[775T��E���=���E�Q󈯟_m>�³��2#� �7d�[N��5.�k;�:��a)
�@�b��	*F/�P?�_O��E~N�!aF��e�)t�m�,\����q�A��G)��CR���+�@b��v�Ѯ��uJ%"k+i�(.�<.S����8cV�=D� �{Uz�!c�����ֻc��\#�S�
�	ĕj/���~QXlxVHYEB     400     1c09#U��û"�r�:�L�����>`݉�K��-]�z����*����f�8r+K)�\�h��?C+/�ԅR�KS�Hob�.�A��ՠ��D6h��4����� �6�y:ڭ��l���3��Qb�=�V�c�p�ʎ�dn�b��^YN�h�۶:8�Ub�ɺ�v�g�]/��AZ�ϑ12���d֖����<�ir�՝�[#\༖�q��V���U=�ϗy�Z���pwG��a�7��&-��C�� )��}��L�fVx�=KZ�`�)��	]�X��������H�e�픤�����j��P�>�z�u��|��y��˿ϠA 1��U�2cM~�ӠQz�7�ZC�Y�����j6&Z���,^�N�
9!��\�B�
���j����B���0���3&��D�H�=h�ܤ��U������p���%���ߧ�R)���[�BkXlxVHYEB     400     150�tPُ�Y���D����9��ؖ�8��bLʵ`=V���˫�+`C�7u�	 �����*H{\�ݾ]�� ��A�,�#�_$�;��u�Q]8�ύ\�^�Cp�����2��b�a�݁�E+	��!G8T��Gw^�ƠT_o�5O����&( 8:�H�ƿ�cDoQ��d�H:������ҝk:ܽ�ßu/_��������{�� �8�l�?�!h[��F
-S���j��Z��+k>��&�K�/���ŧ!_'̦��v4�S��@�=�0��g��aU�j�G��WQ<��K�ĊwdQ�¡�#c+�$�jV�%��Mw.���)��t�M��XlxVHYEB     400     130ʙ�O&�b c�A��9x��J���uDl�X!��əf^��
5	�V���<ȽASI?�5����[W�M{���Ǟ Ɂ4��xKG�ܻD,��#�h�ͯaX��p
����C(��(JT���{p��]?��잌�ďQ{b�yO�J8Z[j�/������|u��/�zjC�&���j����3r�T.f�SՖx�����;w"C��g.����H hmݩ����(�7��m��@!�CΙ�/��bb��^u״Ś���*m����b���i���2$"�O�����Z �ґ�\I̡a8�XlxVHYEB     400     160�5��[��P�
`�sm�>Ui�c� ���aB\�Q�.CS���thޥ���N�8>�~h]�L�I�)b���Ӄ��4QxM�f��l�؂o�J>�����tpA@Z����
&c��/��>�}�K!��U(��SˉO��Y5��/~� ^���`3�%��=�=�%�A�g��h��0n
�Y��u��уi\�z�k<F���j���Q�H�����,������&��\�M���1ك���R=__^��*�cl����'Wj����>���Uh)hv��}��>��j����O��p���5�T�4�Q�r��5�3I AIpl�}1Zq�������֙~���XlxVHYEB     400     1e0_K�	�^~&�/$ ��O�{ؿti��o������
�=�܆�q��sɰ��ex �g�F���Mm���,�+0�����*U!W�������mf��K��sF��	a@97�)�IH�5l@�z�F��(J��B��j��"�G�j���,~����e3����8t��795�.d�W� }��� �%E�x[����t��;�*�Y��E�D�3.�Ѡ��������(Ec���꾀N�W	��L�G�&TfY�����x'�_��U�\����ub=����qPՓV�g_#�чH{p��Ԙ��h�?���n�Z���I7�eDTM���� �2�u��ۺʼ��3~��츹#k��|�Q��,ԥ�N�NN�x�=��z����\��B�n�|��Z�	�k��m��7�%���OQ��4�Ŋ��Qц4� �.��r)�Mb��a�� ���]�%��I � @_N �XlxVHYEB     400      f0�4��J��m�
D�dåB�:1�o?�� ���17�[�=>iE�j�q�*gXi;A�@+a����*"چUJ���`��� ���װ�� k^v������f�d��3mo���B�H3m���㤊[�y��)KDH��5|�5=�>ji��Q��Ŭe/s�[��§��Z�Ŧ���c�э�1�.� �e�<}���OK�P��9t�mS����\B;��XlH6�:{����r	�`��G&T�|>XlxVHYEB     400     150^1LK)��6���m�`]�Ben��SW��Q_G�>��t��&E�w�zS��9og/���&���{���#����v���-F�~"�GSFbA��xKR�ڎn�-��TS3�jWr�>��l�Jb{G�lw���SC�+���)���^��Z�=��-�ƞ�%��ٮF��U^��#��Q�>%d�{���P�z�;�-PX����I�fy=~K��լ���,AF	x����J�,Y�;�T~<3���<Tp���(2sE�����`ve�?Nb�=�&L��&M�ʴQ �9��-yWUK����&q>LN��YPC~��7t�st�вEi?��XlxVHYEB     400     1704�6��K]����6�'�t
%y�)8 �i��)+�B�͋xʚ!�'(�qt*c��5-Y�׀l`�/��y�0���h��O>���X��{����t�����I����!İ�S$��$��0�ʌ��d�eH��q^ ^:3x��a��⋨b'/��n��������.v���D�ټ��������څ��-�
��W�v�ٵ:�@=47Pk�g�Hx�G�_�͍?F
���=�$�,��H���d)�gPf��K�/R^?�(��	n}�EJ�qp���q!]ۺ�>,x~^����<�[Cҁ8d;-����>��L<$Ч]� ��e�2���d��c"�\5��xq� �u��.��ba�=�XlxVHYEB     400     160��������	e�
� qk�
��`ȝ����vn��1f���=b:�O8!��[B�B2��:�z���UN�q2j��5�e�وp��b��l��tש`i��֑��tp�TF�ӫr�a�}Z���N��f��z䲒�	�u�\�^e��ϔP��}v|*���+�s�Z�v �@��k#E(���jfʪ��$၀���=W���Y�͜Í~���Xf�Z���'������*��#.�Ռb�����	���;ٵ�d\w3"���N]�`BS���������c'��3��s4�-�ٔ�BRnXc���v�h�aqI��cʜ�!�|gw�ҡ[J�+iDǕFlXlxVHYEB     400     180��BǗ� #��Q%v��7��S<�V�����;��1����T����`���`�>�H���[:�Ч>�p��h��9�.����<6��/�Q�n�yD�©��Y����� ed�}�n�r��X�_tx
�n�놙�����()�`�� _�	0�15����֑ h�Y"�첻��_)N�c	�/��ס�����XCG#@-�}<�y����������J�x�ݣ}N���X���F��	�I��٘㓇�����f�0�Au&��͠��=zo���U�/�؃�{���"q�?���C�	ԍT���9-Xk�s]��٦���%�#W��}"��jX�e�M�4<eü|���\��c���m
Ñ�maZ��XlxVHYEB     369     180\Z��,�g��SDs��FQ1�HyK?-?�2��gm1kL͐������Nl��Wn�O���6��"G7��ff��c��M]*q+k�A��iW��dPx�IQ���uD"�R4:yZ/�Q����T� -���8<�����#�O]�1Y��GI���$3X)t�u��%5[Yk�AE*�<���#���}d�)Km�����#R9t0���q]f��=>�-���X$���Z���7jܐ��M�諶*�O�Z��{-!@��H���F��A����&�t᰿OK7.G̹]��[���-��z��|'��e&\��A�o��� �)g�n��J�;��~E��$܃)6g��-W��=��vM��%q~�T���Vw(�~v5=�