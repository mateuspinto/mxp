`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7472)
`protect data_block
MPlM5fGhHIyuEQF0ZcyI29zils4qq0q/oQCBVLiNpEq7KBd09j9tj/W/0HC2IgoOwQJYlf+jyYDq
sIG6P+toajAs5hvbmvgoQiQjbwiYl6wHWGyOVMw+fL1leJ8Iad+wJUimMfx+NK8AfBUEsDYZ4M6t
7391xhaPgxmEMAb329AYLsXMPLlz/j5L2tdcH54qvQzzKdkf5UYntB+j4v/vJKUAM/mjD1Y/Nv1F
oHsPGPCnQ0kbVt/0AvxkYp2L6AhMtskPh6ukCOmWRoNOaBJi4ze2CqaVO1rFzlNxUbmgqXcIboHr
XaUGdW0aYvOd3BxYijw6O77q7j0SFnblXPjbM+PEkjPi/mlULWWI8noy3HJCv7594XqktDM4vDaF
guZBTb/IbDIOH/PT2nrGol/C2Dlkai3nBL2LKKB6RMUt7QVLVLZeJVOxpUpDsia55D7HJq+JzPE/
qZSsGQUfmBiRJamXUzXRdbnKvnTdYXkYw462hbLhFqW9Ps5utuOAwv2stJWgkHDcGZE10Mn9ubCa
/pRLIiUsa+axsSNk3ec1tSAdH+SQdRpl2MVYy0rWf3uPe7tRYrZjAaaOK6mRhRoADQPXXlL6thix
6gN4BAuM4Mw0jVMqgT+tJsa9YSMwrtORx3bz5mlUEC6VyYIFcFPxjD/OrrC63DTyaWSyc3xwyrsF
TSKtFa9fY6GlPyoobg0kn7M4jo5QdCDRBaBf37EVO7cneleaRtzQtlTLQOOxTvBJz3TK6Rk/b3KS
1TMIaBw4z4ffhC6PhFpVfY1MBcEMbmMwcOLDuPaq0DD3xaNIs6uNVe+PfodDEfxHh4ym35lJbWJ/
TdRJi1xutOPOlCtkT8xEf3UE2N+n5t1TJyYng9Cqve9fGT2aDbD166p0uXNygf8lOzAb9Hx07iwx
DZ8POAdoBIW9QDvfw1Al9J4V8aVsIzkt+1LJwBnOMM1M66vpY+JXfB5Oji7JYuG5xsEy6hCNAdje
fB3htvPF/AuMrHD9NhPjGyRyqlOHHj2YzU2lXX8lB84bIoIbuJAMU9WN1Eg3nZ1rE3RSleeWgLoR
gO2XUV48rraIHqfvIFC4dMbdQm2iEZWchocc9JYQB0OUizk4XBLY4LOCp3vn14hzKYczEsbxeI/I
FwODr3n+EH+EbKQUDUa+gYhBo5QfJVW0FsR5RwHrCDidN2WehLsxf3+uqzdngRipHXD/9x0tKsvs
uqijwYMCgLH6QOQrpG34gqBgb1qQKVVhPaXeJP72UoBtHa55vctNxYA0zYh/tx2BF7IAYyhD1J7R
qkEnIhVH0xWqifD4Gjc4aRjWhgT9cQp1XqUAJDXPkYYt7LgBZw8lvNMy/h13m8By24EqkSVSJotw
Efaceh25kbXRKkmb9Hoqv8umuoJ90gXidMhM5K9ErffbHfrkHedRLo/Tv/Z+ivQf75ytstpjjea7
II6H2EempRrZo/kR64iIt/7/9a7RKOMm+cWISXDDbfd4NfMe7RtmxP8mb8ykTwgFdXpZ0YvEMOop
miXnC7ZQOJWO2e5a6DjOxFbmifdGvqlwMRiAhQE8VJxJ501XmDKndc0MptzgRYnVQbeF/7R4rzBg
GLkA0gVMwp0V7uxEzuT+AHK9oMa3CHcXkIHwtP5pGbbIQHKQpoHZITJFv8NxUw9xBVq3rKmSACaU
qljNwCgHhduYGKSqIFFPFTMSoOgNhpmbUKCrj60e+zGy++TS59IUWEgxCTBsKm7rAEXzdReSUQQ1
rVziivvLrtf3baCSx/j7uDY7hADNYYDpL6lCIRhKr++zg8IdmpYX4HbAwocbmDD8AD3zN8VSz7qu
75p1y4oaU2e211hoQyZCyN354hw9rlGg0guFCukWlXR+l+ZJ24BZTN++wBoG0cYVyE3WKq52WKpq
ggxqjHm+oW4xR6IAmiO7hoc0IKci1OtzeDm/4QwiMvjy9qQytKgGAr9/DCezykpHT0CTtel0um2/
gOBCB/7gDjygAwCaMLpDknc3EOZHsiyC4ifTOJybrxM+6u8o5U2jH9mXbsuUmUEwitcHCuzphX/i
uPnhBtI7eWwmg4hh+ZD4TTzV/AsYXrCfMNDTDaJizor0eObFgd96vW7XoUk3BoPRmUl5WQpj87NQ
7WEy6RmYnhk4hdW6QjXxS5jsDicjU8cjSC2GYMXRImdiOAtGNi9+gOSZubV3XOwXEAHhLqblaaXI
6ElYWLEgY/K9wHDAIkyYXxSAJXDtKFk605ZU5BQPEBqhPwONqTDFRfaYigArpGhEroZFSwGB31GU
mW6AYVOWDI8xvUfeOTxnmWpjAMnHBnvf5xwjptgq7ZZftJi5YJpoR6yyT5emBNMDEncLd4BbPCfv
zZxMqgXz2T5GXthe7vTFalxB2wKB+nRABN2JBXPYJmwkFYpRhhV4z1/nMX2PvAWt+JxCgZjrdNGd
Rv0sx4ZlcZajgPanHPFpJEi45qmERRNMYdTlForaVbcHNqqvamJAZv0cWAzXWl1Ba13Z654CO00P
CWvCKsBDs0yqbueYk5Ion4WeWf0WnP/7zwacK5F59TyAlVoOh+CJ5mOVEBejhcrTTiHHGCYk7nbj
jMT0i2CXg9To9Zze0ZZuoVLB33Tb4uO7ZJom9fOsizK0J1mv5gliT/RbALyyX7a2cyyNkTUJvx1i
TSpAJ09GWGCjz/3yRDdN5kTTCPAEgDbGKK7cQ58B2/UoxlasEcLTPq/BOItRmsCAu35ie48eS5sC
0UOYVuSS8LH3zm/i5THtFkpi2c2jg1CKYpyS/Vc49oXtSnFxLjxGDUACC+l73E4woGCRGkF5/yX/
XJVHtCGkbObSLK0SR8MIUB5WG7qne4kMWK2LJdDz1eDsbr7LnQRZIGpBUo2wJCbuFKURFSzx8qOb
+fGNhKFbFOMMjL7pFv9uVTtaRdjqktMcLE+zApGTl3rOeW/vXlAbwHtuFduDGa+/N+hZZKcqeHXR
Jf0dodIjViLm5aXWx5lFUyazCIWOusRd5LyjUlWvDCFIS8plKWQpw6D3xgOXSifgxfuAbmSGE4B1
LQsMNw0D4ZIOVeKX4/XjNI6vhFGeHCojpbxYQHJXfSLqO/i5B+sFt/LPPFq71jGGa5kTH+pWB29V
wAoyMSKBOhzrQ0LSS5LSpI7n+6cM00XyX1Hu+Ynh5zvPRdB1NiJMt+u9zOt9osFedVuBPVM75QNS
og0McPTM4uEg8zWgaRpdj68nZyQ7is/bqFATyaiFWn+tGwaX/RAVcWI1FuM5syh1ZcISVvbUlSOq
QIPQ+hAZ/W9bwZtbNGHnY1l4SjejCX73Z6i+ZN00y0tSjJ6fpfguUek794i/y34QW84UpbxHabtU
WLrfv1TVlhiC1j+RBkM8enqpH+Wwp9890fXqyGIW/YcmZdYTWjNuOThnW5Ee2j4HKIPgsDHaAwuL
tMn1MGvUoz7RaZ2pegFd61u2NJflz2T5Bhsx2Yeb1T9BehM2Gzs/oMIkLvYhb2+7bhExAEzmnV/j
ugYzg6kz6KcMkg9xjjJ2rGra0Esp3ZBdqHx+IJj/yfVhZ/zxgLkzuDBV8mv9mNFaZp/X7DkSbM1v
ejfcxl8V4JOF67ybFpYvO5cpe61psJybuYPlD2+mWz91ZrljHTUIHdGIgBKalpN6YcUrKSmAaem1
LjDyPwlAUmzg1G22WkOgqhbeElsoBXY6g7kwjvHm5VghJI2DaNbKV3kfpNfQucsNAc/NP81tNhsQ
YMvvkwApbSjjahgiuDfbqUv0mQtdkmec4lA2sGpKaGsFQbp3Uw7N+oQpMFovBfNrY+i/PfHCftza
7QZDR0u0pL31fx3B1aBO4QC+pUglz3g0jxD1Vs9cM6qcKgFovpLAoPH8fwgKa1ExXoq0Tqe/ERiU
uUWni4mS8k4W7MSFur3Rq/RPnRc3sKemq3wWmmUEA+Za2Fe43tkYKwlZBs8D3qp9WAFFp+PSDZHj
GnFJPY9uP0yj1pSB1EESzUc3lHkqBiFH0h+Wk4oCS+fS+6Ns1iSteADy+nE5ejrAmQxnQbwaf76y
zMMMJHLf7LNeXBxA5iIDB1hdC9mvPX8CTOkA/NrHCcd3ohR5QI4ocu1PL/eYd8RGalEkYRJyOaD4
4xIxTG+2Bcp1RcQHMlC63sifQWPO5HBzsiOF6l9rQgAsMwiZy6PbZTjhC5uwmMuc38QrYF72L5rV
rKo9y0oGkeV+gLF0+ZFbqUtdbMfqZTm7flr6Hzc635ZWI3hc6zzurMnPY1pwjzHcrSmcQETo/htR
QLErDigrk+8a7gcLYqe+7/+c21fDT4N+aLsGOqSSH1v+xi9a/MlBZfoWuU9rtw6PfTt6jkaNAwxl
2gdS+XDofrW3YjDZYawk5gSGUFHoh+O+iROIwFpySGwCvVV8lQTJNuygvm5Y9tuFyV9uLmxUQB27
oCJ/7SH+xjXAhp3IRBesRG2aZSZs+V6r9/cOPBah5H6UWMYPrHYkfdDKGqbFOIbZUIeeLzuqFMw6
H1KVruMg1A+M1E9vxoGU2e3oBF4Y6dAH/hqmIqEoBrsvVGnHAq6K6oxJg5rCHFW2YSoaZV9iKOC0
4v3gXEYkPkizDWymfhB9vJE7ftTMJDIc4XxqSy4ySfHL0PErmfEd8mSzdpYSh5AjptgUwPHErIhM
iuigvx2ZvGcRgXeKaQEbpnIRP12woFjr5CrAU34ePFPfaKTAfuCx0mKHKs8h5O1SFkvsMOdZXzYy
AtH6BXqvR6gWd5PLWvRAnoWaN0vZ7t2FkyAHQQncS1h39bmrBpdYE+VamssrBDnXefse+wmgD0Ou
I5ThogHu1n/RM7ukpMeGbNUzYkqb+3mnH7IEkV8olv2i5JYMvY9p6p5ZbXGnm5TIFYWDBduW/92Y
KrU7wlnSxzrkzNRN6KTQpODPhr7muZjHU3J2cjHo2k37f+csJcICJUIk+E0SIbjo+IQ6vN//Um+7
Imj/WybnfxQac5d3FsfE4hC/s4Of2+xndV/qWOGIdoUgYojz+p5+7HOrdftXXnkwwyKELSehzIp4
MKA57tClWxOYbumOCURNM5cPw5/ln2J6YEt5o9j2tujzfqJpBNE3TPr7DYynqrp3SlGfz5xXaGTW
iKRe2XSA3TeJ3qWRsKgHCb3yU8jUFK3cPzya+f7LyhuiWexp95y8yHl1ITnXFxSwTqFwIWTTqIMA
R7FfvujlNdl0Icxd9lBiX540jVp4aTsRYS1Sr7tmVVGPswASQWByT3E3w+Ni9EAXVdtm6YvsO7YZ
6kNeVrippBqgJQL7EV9VHOg1pXKAvHEXNgc6NPyT3yajL35TVHz0p5kJyZ9g8a5vKuJnqxTirSFe
HmhbWVqgvKyxoOB6GPgU4pIOowFxuUxYM+k/7wmVn+gcBxrw7+9drAmjI2D2jOj0edZyUVSC5niK
hCcLLaYhqMdeaW3QbLPwqPrQ05mQqR1YvO75wNM4+hLn6ivQVIm2BNW9buv8+pyYyIWifBu1pjvj
H+r8WtZr7Nr4ij4ILec8d8XOpwuAzLPZCZrpr3spwnHfaCAak1fMYIesFvHxnirkdEIDmdjq1JDe
GTcqYb5J/TI84oKKkyrXBjihiI1dOAwWY8lY9GqE+sgP+6q+6gAjPgo/NX5UZSHdRJ9oNSzUvdnQ
Ar+Q4z2jMX8n5BTzCZaUfL+QA1ev455+KdSrC3zYkHwwa+9NZ3QiDt6I1bW6HiWy33wthNl8OPEd
Mynkc3uQOH3rZzV3vS9lZSfVdC1qONW652eEDGkWdctzdrYhtGM6i5CYKA1GJestGhQ3/s8mWGAL
b6otZ5q7/RB76hHIitmIv5ezFr7H1N5RUizGVXwPiEluFXOncTPOLedb/B+h+nU3vIMYlyYqzHx4
3acvEB21YHV9BrVM9J3OGOmMVxS+nb9WvojOkVJnn5LS51EwQoMYvcma5Up69JfpZtFL5tiaRl2I
QAdCFBvkQlG/DQMdAVYo66gTYGjUMndpHBfhYU6O/G/Hl+qaFZPxWQW+CDBGrmN/KFAZdo3mGsGz
MeDNk7K3WoxGbBTPNV8SoQ06Hmd4n8Uc6Z5q7BfixSdhdm/vz79tz1o37qpM1X9XwYR7lext44TD
HmPN11ZuhnKCT7slH4PDwZKXjCQytY2BjWIfxl6oBaGrYkt09Ql5hXWdsCvcggq8xO4VDyUzyZrL
IFqRvBeKvWv/redMfZewF1232saqAi6zHtZHS4kC1HqkUHCB1XXHqta1lhR8WWMVAN5pUHaASTpH
jCCHKTS3VZWsySU6C9whHnje4QbKw7/yCZc3kAWZDiRJv9KZVJyQoed6/G+tsP+AVf9PR9Tk+dah
zaGvAuBU+Sxz3QOIgV4dvG9GAntzvHHkSuNQeAlhEGXdt/GPnWbiSd5HqMs4X6/a4R+b1di2xhnq
o6+MFKRdToziWzBrvu9BmPAlkS91d6UiqxFNgkauoOo+3c2beM6RMiCH8/aGUqDdZRa4kaBpmdsF
/i7yvHb6CQHriEoMzYSbwtslTQMvjgbZrkq1tPtFZCAE6oPZa47ppaHaJgYzsBVeIhFf7M506lRY
Ry7igtGFAn8R5neAEDWER3w2klnqsOYLC6NiCgUW0zZfQkTs/Y+VTD0QpMwAF20mE6Z6JSfhSGfa
ffBj7C35CZpK+kHAncrjKbq1mRfqVoCq5OOT7XD2dNRxRXCxs7vYDjqg6N/tBqiGfeFa3nLaqJ2D
LAhbXbIMA9ThEGQgsyDLCtNNux24rlXiYllv5avs/AzEOwxDNyv5O+HzeBKP1V8lsCyGuWiBOMaU
W5bQzZFEIdlA7wpi7IhszVrhBHcfgdVShL/PX7OGfaZ+1NXmWdzc6XRuqjRTGY/vk9odBo5+9K+B
vWuahA2oSl+hT338VjLkp39tmUCYYSP/fdGBzfkt20cKTZYZ95/uvRqMeuKQFdupIQ5gNu6+EN63
qMnXoTrcvOAd2cmHmO7172JbrIBwDaBI/3UxOV95ZB8il+CaAumQnrLA35eQTuXA1Qzmc7knfYlK
yEib3xmIp39ev8EbzQvKsVkWEhEn0+i3bBh9o7SknfHsMJxJ22v89TeM41oEWpQCDCe9q2rkmOqx
AR1Y8DdWspBsYMMxuX5mebqYujrOQ7TaHo+LDNe5/CKGMZdhxLDaUrKE9r9gD2CciUG03hqcRwjP
63Xs7JfMWNMMSHD1OIs/+Oot1dS4QIp/P1cNiCzrgXtk3TYby8gDPpZp0Zd+/Vu92KmrTWnIVm/U
Ys+ubskbtt4Bto5dbHrQxADKQCGZCFifbiHwgHrvaPsfoes6GbGsBEyLKC7oTXq6Pi/Mh65BSvOr
PfZHj5B8jK0Xs+N8tMn7q7ebTIsH3oN3wmCL9YlBfE5jSVNl8mFpT6vzE1HOcn9vpjPBsU35CGzi
wYB8DYo+ntMiyGuifMntsSSsS4Ko33Aj+lhPmqG+xjRC84nLIj6NggC7MGXE2zUoRoTuEtTD0aAm
np1Ls26PIc1EbTd+IMZk7GnENEQIdSmUaCp+HfBKA+w5TdDST/43GzwAMSbO31dPAAIyujpl3zwI
Psqj95Tb408PeDb+ElBiEf6y/0liMgsaiE2uUqEzegODBFSxRtScaOoZP3UEqVLti+2izpKqIpVA
Cpmd+khLaX9nYXVBS5azf/1CtFN8aYkyW2Mz4r18ET5Ill4paZH1Pt6FH/7PTZn2LeZOVDCNx5Qt
x2Qx8C4nzvZwJTLmc0MekJfdfeZBBv+VU2++0gNTXnytDE8X+wxff+7lH+H5hTrRqb+xpgwbvzHc
FXZBkTdfbp8IsTNJMDAron/MJZowy2AOvNAoadYTmRvK7mLi7z3+BqVx3PuyXJvtkXWyhxjewBxz
PoVfPChbtGhjvFAUJydHZlvG009cNJdqelHQVrYPQPmYYkGwXIbSTgjpzVoT52b86CN7jAglPuCV
rG+TEF8krhfb0VUq9UhSIdYZrK0hKhZ2mRGEuiX4dD2oWwd9TE6n4P7zIV+4dafx9/iNMJqpvfa+
UKSeFavQkBkwGcCz1oWXIXgD8uKsZizOicNLSJ6AIr9KnyatJKg/dXCNZaMu9tl0MVsSQ8QxoGAB
M2foZYH+yFuiecsqvgk1cp/7f79LS0W1uNqgu9kZdw8QfAOMxrvPm37eUII1Uosg3fbBYfs5pkR+
uaIagNoX/NUb+DtYDVjF50CK99X6V+BxlU+KO2y6Vmn52Ecqp1lapz6v49JUBB7VnBpQvlN5xq+7
K/oTSSW2WTSC10JYpsgg5wmAStiLrpxbN8mXhjIOz9A6yX9IXyhvDTrzfhhKNdb+XRNvpu26tpuI
lNGq0PiZKSsRHtyr8w/O7sRzHQvJJHY2myEF5ukul7X4oKQRk4srf3eJGCsGvUE0ATnTmK9lHQWp
+8zZliw8RhO7BCbN61dQ/3uoQl5YASKBYRWbITbUAHWwvqX1TMtEzTwDgWy6YVAJa2etV8bQ4twf
ocWG+4/+/bz4jfUl+xBjS/LrtAseseB6ctCOhk1Y1iOkANYBwhZiddPi1iRBs697ZXb1rw0qYThr
kKbyCOQthtBqCJ6+/hoQ8EqHJDAn2ypqkyGIqEkaz5S+moVIijBxAFumsRWVhjWURQ46Q+y3+OBR
wWHUS9Su5DQEw/Uk631cS8FVo2SHaVd3v/iRjAlcLcJFkCFcRtxW5EZmq7RKYSaoVSlmkXASxC36
vSC54mQNRfNlhjM6cILqZl1LyoaHH8+yO503Bc1KdDc9swNcQJJujSjYN5btAAaBttGPaQrrzhXl
QTDbwYaGWpJqSlv5X9jmyYSR65p1Hkcw7R3ZcDnI10XG9j7wofBG/GYzgGXlm/v44p0vD7XK0JkK
m+A1ldWvU4eEmvMS+Vkko6LFanFzniXIoW4oPZH0yq8Cc+ItBBn9xUsu/HckO9BOoVMsU9DlK3nn
eMd16LWFSUuN2CeGH+soT+Eb0f+mKnIJ8kIqGew2MCnCKe0wuTWa8ZENbczn6L1inQUJ7ChSaV4j
fPyw7PcwvbTc8zl8LgVeRHtphGn/0omD2pBZeXwHkcrltXewGalbbBBp1Dj19uFnqtWpFUYATy2i
N4zzzgdX06ZZT/C2AN2M88eB6rxV5WfkTyn/LHeucQVtcFgng2OIXtX+3kXfViAkYGRBNmMkMQJo
tiOK4u9mp9oLiG3ZdjCZopYn44PnFBvEpXbwrIpMH8afgXMwjFY2e9O3OtKYSa2m78XMqha0YInx
+UtN3W32CA3b88TfdB47/aGGLNe7jA5Frn7/+GHAhYlcA4b91JSX+L+eIqfOKRlEybpXU35Pu81z
R8U1NDv9fM3+12GvgOuQOOeGp167fjwqYthBrd7tJk6E01WlxTHpPQpNaUgS27zY6zpBsrWtWNDq
U0OY1bO9VDI30IYhgoKw/g6k0EL6YkLE/oPMKeb/n113AC9ZIL3ALOGoXJBJDcpMa2AzWpx8DX+N
YHxKO0yhaBuGgaH4nEgTmFwPlG50ouCZ3fOLAwztfokdoRXgBEwXjJZ+91Ayt/RAyyQQVwv0m2Ly
AMGeQpTlJq7S3nIBW8kn5f48v/gM4GUg8xqO0W21iSEwSCXHHR9/2wDbGKDHQjAwog9M9K39dAzP
qLBvIAu7ge0pb+ppI9xKAXwcrKjG+W3VLdbOplkMqjL4A0Wz3pYS43Kqh2lz1Vj/sXNdemPS2WWg
VBmQrYB3JiZ5l4gTZsG/jiS/LKYxmfukUT68boeNDHedMEsPgLBh5T0LykWorwsf00wEQ2cUg4Vb
gblvD84/Tisd7L1BSoXoaYIhadNHOoWGeDaI66SAx9hSnPRIHuY3hY8+semG1DRkwajGT5oQbx3h
+9GMr9sTrPzzdF41rYipmlaYgvzqprgnfthCIEbd6ysShgWm/DbCp0bgyDfvsa5nBov2x/nOzNb8
FrFd27vTjanzJsaKrXetv9TVM8l5pNFMTVyQFWLHJarzQw4UOS9At1ePlQdJwmwmQPyeI9BEilir
qiKWVtc=
`protect end_protected
