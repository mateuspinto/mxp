`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
iibBTkzgCT9UIsTk684+FZZ2G1SIp7RLQSLZtSXbPNL22knOw2X9ySt8QWDGQFFFUlqp8zmB4YF4
sNhFHeVBjYGjOMkWzOda+5vHOEgk2B1ZXm76Dvswy6RysOp3QmbvVpyZq98wxkAHjRc8bI0zwQLZ
9BHr+NIcwcClhPym7jdlpQy7P9J6yglaxszhRdPd8nx5QEjFfkkE0T1B0mtlDSZnkd3FCpGUiZ7w
YH77bJhHdM/01wJrBwuxsfiwnMIZM3t38q4YE25lYm8ztPLgNQQJXAeAzk/U6FjkC8s41d6bu3ED
J3cK5FsgwAEU1x4x9wvXeE9U/M9vneAHYWyjCWKWFvNkW9VTym9QhuqllwjdgWR2ibAKxEPixVq4
94pMxkUVKKJ+SVmDW4trrrT4hh8sXVWHSYGA1YpneTkBTaMcloh1cy4r7jQbSPgh01nOTGobmhHA
wkekYTkUcmvJ/XbOswx4lsMDp6akSNKt4Wh3pGoivXO3/+HtMvb02s4WZ44ScwEF9YkMLcmyBi1g
Qi7K0FJT7S4dF5ThnJjRHZ2J6icFk3AXl3XkHVkGnINYcpUuatQOeLKGcJhxSBE3wrjhL5/7NNcc
r+yqmfa0zWKlbVfbKH9qHmm87+GlIbgz36+hJbgWrg36tQnCdMVGJfhkZsiLbLy0b054DoSO3bp3
C/IBptPsdz0JHEn20AVW6JPT9KMDHzq4fSUd+TN7mOz+81Ew2oZCD4Tw+5VdXzMffpVOw1BWoNwr
JIjCe6XVaOSRAuPgq51OuCUkYSmsTgoz31H+nzOk7RqtaI9MFXL2VdrHQCLCGLSTuM3JQSDwzUr4
Id6iH6bVVYx8KKQT3HLqZIFRE9bbGFip0bn6CGF7nBCaAyCHpdlEMb0UxSWcDk+Pp8uHdh4Y4T6W
9iK/6xsof4xXETdUcaX4Z0qx2L+J589ig/tPah2/jenrdTLYRVgNIbAR3x5NBaIsIsv1/sJi2BDC
bDMErsy/RcyCSmWSIjThNvudcTv3KkTxLYM2ymQWQJIuwmbjFQlvrvW/jVBts+hy6VLyCicWp7lv
SGK6o1EXTxfRIWOjgowhQ+1/Q8uA0PGE1xegsAAm/9RK5gCJdQfkeipvyiyl434rlgXMUz2N0ztN
QqriQtbrwsi/OuJPtRw7NigjO9YrYNYD4sh3//1eIckB1lRNjP/SuTCQjcWbnSiC8P+FApxw3hiX
CfC17pX9dO2uV7GkzV7euKeBoBaH6xMluKwHY92W3ACjNX5jh1ThO4dSKxlSaud3hEANt21knEvF
GYVxpfRWs1txs2m5zyia0IU2bTY8aMdm6lWE8veDnEy/2Wl5fDHCa+3/XUjT8wP9TRBKW6Td+QyO
KYqvyhRro2x/4MoVfJ6IUFDIY46nwWuBBmsL8eEwDZfewfwYX9F9jDRiNa8W7LfDvmSn/RCltEyH
lT/Y4Y5GqgIFst0jtYYfNKFBe3We7sd7dWiy4pgfs5zp7YwQq5VT5LPDe+Im1jyPwOrzu+ELYXjE
f2lTI4TT0HbL4XDHRA3IU8jgB1fJkJd12maJ49KmuJaCMMjJ/J9m5MaHtBCB91i+35CC5ZKjw3du
YudIRM9lH8Q7PfKxV8KW8BVnIhPj2HQ+ft1RBs9VcIbRJC7kMjZHoc+qP4KC2xvRIRJUQQsRMOMJ
MWK4M1UcUfDcnADrDBkuqidNJtRp96V7s7m3fvjBCpyFTZigH4QWYQQj3M5UeySbVVSV9SvKc+BL
H5A+3+Rx2kN2R0tdz8L+vnBiuEUrj14UJhPro21EwrLh4H5Vvht1Ueq0vfXQborEI6Z+vwhTP8ua
egYW5RXYJRA9+WYWWRxUv9382SkYEkJBMdl1kNNbbbu2qs/yT8Im8jP1qnUPUHoRlE6R/Kqqwr8S
eT9w2S0x8s8yvn4aoErza1XwQL4ol7bqfabJ1UQPmR0g++0yKDUdmlHj/otSCsGyUldHuC75HemJ
DXhqMRJjodmSueQCYuD0ecN6t1clWSs5kpiJRpEtkUDHiPt5DYuKi8OOM550Nk5PHmBtM02uAWCX
snOVWbAgIfNP6OXPr1+FyMwkW0QMszrLKPqJet85PJH0uOJUNA7RbWAmwRAU
`protect end_protected
