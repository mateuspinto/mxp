XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��g)ܿތ�d���l9u������G�bF�?�3�`�M����|ѭ�O���q{2�Ŕ����B��*|��{�s�׳¢��bƙ2Qm�K���� �U/l��q��˱Z2Qf�K�`���[2����K�Km�XUy�h8�1�ͫX��:��Vڞf�V��U��31�BU�U(�C46
d�O� �$V7c��)G{;�)~CZZ�+%�/�a�4-�%~��c�+��H@:@�ˌ��i��������a�7+���r��������'���j���}�]�[Q��������Nҕ�[�����c�O�?�������-J6��C�.�nʚho�)_WaN�� �v5�� ��D�Y��K�B�n!5���^�[����"?Z�A���O����J���[��Q*Hb����#mN�Z���ln��:�s�P�1���>͚L�;�_����Q�C���C�����C�/FNUO��s�P��+�/�r��yMn<-�	��:���h����[c*@	�@�r���'�B�R|shG�8_1�Yjh�a�t�bee��Z"�'�\��5�/=����ZǵGH�%K�~_�p�-BKC������vޒL��� �������!l��0X󦥬��r�F�+7�F.�УO��:�)��G)�h�ަ��c��A�j���ie
�m��g�ᆻ?/��{>��{P<k	.�ѪZ�ߥnF�D喭�N	K�k�}��Px��N��Gvt�9�|��>	XlxVHYEB     400     150b���n|)l��-����� +��]�Q>���|
Xz�*;���X'/H��Ӻ�!/Ly�f��z(�+�a�r|���ET�.)�J)�������F�]n�y~"uz3ArQ��Ⱦ(��fy�h��e�.?�q��M�n�i(/����������~S�^�4�K4U(� �T���=R�?rRvl�,x/70���N���4�-F0M��^�/�#u���
h��\��j-5���4F�M+��a��sv���}>k)��Ay����f��|�?eDG�򔺌z��V�$�h�`��Y�eB����Bl/��"�e
k���N����h�Lj��PP}t9XlxVHYEB     400     170��+1@���k?� >w�ȫ���Q��� F�Z�����=M[	6�- 8����o�H�5���I��n��I�3ͪ��l�'��\dŐ؉�0j=�R�2�	���������9%�{-,�b�R���V� פn�Uo��\Eg=��D���}�I�I�>��c����3p��O+���V�=~�{F	m.Lsg��6�F?XH�z�V�GB��S'#�1x�aD�ѕ���O�M�a2Q�K�i���q�L ���E\��OR��T��w#��2rR�sDs<!�s�51�w�,u������T�@;�٩6�>��bv�9~W���-"�S���F�h
���֫l�xs��0*�x����XlxVHYEB     400     130��k���i�����w�=$���(�噛�M\��y����5(?��0�M�w)]_HM]��D1q���'�4E���2�In�����@�z
W�/[ ՝�HCwc�I�P�?ff]=�V���0�T��I������4�5�sڛ�u^��
��\��Yw`�����b��T4������p��[��%gS�Ґ��&�O��e�*���{/����=�������nx�:����=﹉+-@E�HƮ*%v���xd�9��.�Pg	�2D�����{o3a-XlxVHYEB     400     100��"P۽[2	�s�J�B&��^�*9Å�D��w^��Y�Y�g��8�U����%Ow*>��jW�7o��<~�~p���Gٺr���}�γB|��k눠qT��")�T^M���&^AX�1�F�ު�{	e�[~�J6�aR?hs�6#����R��RLa؛�m25��u�@�+���%�j[���x��o1��kc�pt�/��ų���0x���"���	G��cQ�X̥/�`e�l���˘�����7���XlxVHYEB     400      e0�['��0��i�؂>�JA�.iY��TV"%�-�,��0xc��bm�A ��
�D�R1!iR�oA��D򥹲9�⪑k�i���v���t+X�+����6RL��	�� �*�<�g��@�B�f��@�dgS܁����F&��Y��f}vhhg���(�������Z,C?ѐ�m��3eM	���o�x��d[Dz�!C�G�<�`��`�1	
/-�m�5<D��[H1XlxVHYEB     400      d0-HPx������\��d�V:Gx���'�i��[xq����E���j��?&~�=*��ř���!�����d�TǈU��Z���4`�(-di~[�K�h�nA�����e�C;k��*��ڗ����7,2Y�S��+C}��\Q�]�6��@�]�O�&�p����s�|K�&Z�A�KZvV˜��h����;���"�#��Z㕦XlxVHYEB     400     120������J`���>�e��]�#8�d� bi�K�Fso�B��]���~���t���m�_��7�p�ath���J���@:gZ��I@B���~p%�I�!�8 �{�>U{xy��1:�6,��5�8�7<��\�"8�7r��꜆WA��j.���qBrܨ�/;��i� ^T���dkS58���J>����#���5���m�t���^��4�8k��8�z�`|!Vm~��U�w�]��M9Ǣ���?��j�E\�U�Jhծ}�� ��0�y3{�.&�D�XlxVHYEB     400     180���ò��cp�6�����xv%�c�����(+���o��|:�2´��3��
�ER����{Z�^,�c���tEڄ+�� �el�K�QM��Ck|��1͟{	��3����"��N�(��7����hTk�V��rۜ����b�&��	�	ӣ
rs�=���9����G␄M��˜:�N	��D*��y��U�bJ�A��7���ЛZ��Fd�ju9�c�Ζ��G���9DQ[�������%<�5,���Qz�,ؙ`�x�Y�e'�H]�{I]+�!I��t2j�ry�֨J�w��qx��t\��ٞ�J�vk�}�_*��&�um>@ ������SB�b���!��}�9~�k���R*���<�XlxVHYEB     400     140�|�BRt4��r�^j�R͛B̡��j�&�l*�h��7�^�՞6���� �8b@�H�R�����"H����_;�h���;&7W��9%�����.e'�9��_�{�ψ�lk%��qr��u1��0OڌwꂜkR>��W �k8e\�����;5�|�y����RC���{��A��9��M%�P�($s#�+4��&X�:4�^ 8��M�X���+0�9Fv��X���[vM$n+����e���!���Kp�]q��������%�v����!f��K;�q�{	��#V2��^�
��\f+��.f9��˛XlxVHYEB     400     170 \��ꄠ�hxNo��x��A�P�v�b^u@p�c�@�m?g������	8��2T��<) Ԉ�բ ����Du1O���*�9��ꋒP"�������l�ae*�o@�6k�ܲ�lR��z7�y�9��7}ml���4q���-�7�M��<3�w۷,z���>���	�Y!�كr����e��!�������ЦF��[���+r}Y� ��/����w��F�4��IL�7<y��9n����d�1!�n�/��I��m��R����G_�o�O�m��G�z�y��,BC�����)a.�{�ɝ�������=v�U5ŏ��AeEӨr�$L75�O��K�i52��/��XlxVHYEB     170      d0�1��۫�>���ڇa(A��[�&�@��RI�*ȇ���s���1��4��3�E�<�8���@�m��;�Y%,�f�X)�G��)�lڒ:��U!sU΢�ΑX��_�@�B��2��߮`��D'�P�5UR����p͢�.��u�)���t�w��1]�֎��Ə��i6��VN#�j/��K�N�ѽ������qk