XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���E7�f'M�9���3�f�������j��̑���RbØ�(RT���GE��0���3w�/��K�.Gi"�t�������i�Ũ�����'��~	�*�`�rd݈���F���r�$��=�$��]�Ί�ȅT�	��L���u�S������ >�#��J��ͷ�}���j�?���|t��D4�*�����.O*{_��7~,��/���a��Ȥ2�#�D��0��w%��)l��h�r�Ǵ����If��7N���L��z�B�eU?�W�HL����O��%�@�ZH�r`�>ӴL���2Tv ٿs���~��q��"�&ЪC�?)��~7K��d\9KN��	��Y�9��7u;*�<�G[|�)Ұq���k�q��>ʟ�uS�c��St�c��PT�G��*�o����|��@V���j�H"�������8mz}Y�䐑� ���^�遉�x�R�������?_��3Z�c������ 7�r;+�0l�+!�n��Yl����nK��X�Av�J�2��:O���������9������ �̋g��7X���\��5g1�Y�	��@Pa�%�D_T.c�[��9>���RV�6�� L�r�i�t`6�)�Xu��Ս��J����_]�9�QG��k�&��;�8%W�'����m
Fc,�d���ֶ5�*O��N������b1�zv����7z�?1�W�@�Pz�G���n��]�㽊@��2�Ȗ���/&����/f��$��`�;�"�XlxVHYEB     400     1c0%�D����WؿvO靣�x�@I=��J͑.�Z�R[��U��;��2��x�R�m��J��(cc9�����>h��F��}�S��wwXT�r�hKq�3,�;�A^l�į���]���K�D@��ニ�S��p ���G�C��q+�e��m�&L���(��,~K#����V�;l�ħ�"�Wv�����s���DF�YC!�������°z_�$�+7= �-���7����z(o��{�aŅ%΅B�=�:4�W� -�m�.\�X
��])bz֞]��P��G/�KJ
�ܩt�0{+��s���c���sWE��H!:'Ґ�S01�K\xKW�N�Lar ��R�Nb�/��C�"#p�y�iއ�(+������&�r��j@i�i�摀=� ;���x?�L�5�8Y��Md�r	@|t/[��XlxVHYEB     400     180n�#K���r��S\��
#�o@{P26h�W�8MĠ�4Hm�����t�c�����v�w�ϋ-3��ιF��]05����u?@�!����7�"Z��S���Q��}6�0�,���"���Wq�7��]�j!c�O��~�7����9�E�����.�goʠ��-��g���~;w˽�!�آl���!Y�&>y;��bŕ�Ĉ\�N꿴���|�ow�R���*Vs���(�f!u�H@N�C�8���%�D
���<��9�y�"{���w`]��QQ�.w�5"y�W���	�f�����,��'f��&*T���6���1��u�;.�\^���-[��������E�l�D�̯
���Lq��ƾ��^3-����`XlxVHYEB     400     150y����&I!��2���e�� �Rƾ!v�Iw�_�Jv��d��e�b�h�x�iߏ2�5Xn���e�b1�}d�筓*�쉿���Pme�w��3��f��+Z��B}E�Owsu�p��� ��J$�C�5l�X�H%���;����6w�Z0U�����H�Z��3�e�e_~�Y����_��E��}��]��1]-���]#� ]X���ɕ����%Q����s&�3�g��cM�>;j�V���Y���-�_�Ewd�� ����>N6P��˕z�qt�����d�2�jg�Jy�0u�WrU��b^�(c$� )��XlxVHYEB     400     1b0�n?U5-2��zI�{�v�k8M6��� Ay,��炼�\���<�J��4n��Zq.r�/ ��4�ʠ��2�-�4��=�@�b�"�\���)�Gd4�'P{U �U�� ��F��kuN���mK�=
ȵ)
j���H��{[a�aey�A�F ]��e�4�Q��x+:[��MGHp�g(�Tc���z��vH�[D��Թ����9`���4g���)�q�C�u��=C%���7�^�B����N턅���U�z"ZMաW���73�8q��ޣ��_�:�h9HTR��n(���B���͏�a��fs#P>v?���t܇`xFBIK�������x.
�֦�謎���#�㢫h���%�{�U>�s3�b~�VW���v+�>b�6������9h�2�d����N�S'�t��ςV"�a���`XlxVHYEB     400     100�뵛�F�����N�lA�ba��Q�n�8�b(���)��H��nk�v�|�̱oE�2�Sk�`�-GЏ��E��z͘>}&���hY�a��nWS����(�w����rP���e,�J�c򎷬�B ,�Ʈɳ�vĚ�����%��.�cǎ#���<)L������,�{����o+�c�X?$zq$���i�M���$�{>$G�_�{�m���A�9������t��c�:���n�%�W�k�[f}7�ZL$�XlxVHYEB     400     120Q��i���H�ʫ�s�+DDlf-(N�ۭ���Ŧ��ueO4��������M�L���L{�x�K�uO��yE�(M]����p�N�sH�Z��.԰�@��G�)��}�[�GD�+<�ʫ��e�ͫ��?[nƲD�9�{��!L�!V'}���&.S��(��0�Y��:�x��3�v�gT��f���5��#���	tw՞t�-���@������%�yl��<!U+�$�)��ꤢݥj1�.�t��V҄�08�3́a��U�{���y��pb��w�XlxVHYEB     400     160Ƙ�F�4���|���+*V#��;�թHi���.�3H��B�X��Ǯу��A}���3i7P/�1�X�夨��� �@ͮ�`ދUű��8H6B-��pDJ��'������h���O�}�^��H��f��	��2��(Ȅ�u���k:Q�A]ZO��J�ui��L�4��D���� �����{F�l�^T�Ϸa���kv%�y�?9�3/�7?�B��.�٘���+&W����?`�C�{$Cj*;�~]d.��ȲX]D
��಻� �_;x A��f-�b�&���rVm��̶��S�S����{c�E>D��AK�����Y�\^XlxVHYEB     400     110;6W.�H�ĸvY�K��Vk���S��&:yx�}]����8T�;  <��n+#�E�b4ӗ�H떴{�m�<^�[��k��^�gu����F{��:�j��%VW�1�=tLMe#��*Ry����Nh7hV���o��Fmn"C�!���}�y�D�c4�d�R��6�������!�
��A�(���t�
�>ײ��#}'M����.�k��>@t�ҸH�v^Ѻ�<�+:�R���7�<N9�r"��#ŝ�~胋9��XlxVHYEB     400     100a���?5z��D��!t�N㐿ʝ2Yk�ed9��D�N���3��8�mA�$[.��
(	*���	���=T� ��&p��^�v��@a�*���'C9sd���_��̠Ҟ5��G�w}��q�������gIF�YC�����I�}�cU�t������Vd����M�6+�A�'r�ss޿H�x�;٪I�W��Ł=�L<.Ed��ח�uKs���������E�ܧϝ�K�s]�`ų�s�D��(O��ב4�i��XlxVHYEB     400      d0Gxg�m���k��r��k�sb�h'|R V�H]�.��o��{�	�/�Ƴx�?��z�|s'c���,L��P���\����Z�0�_U���Gݍ�c��	^��`c?@���l�E���X�2���r�
�o7{��}��$A���F��FQ����L'�)}�k|^t�5F�R�˳�VK����c�jKQ�g3ɻ	XlxVHYEB     400      d0�`Y��EKB7��$��F]|F ���ǳ��g�P�l�/>p�+�#����4�a�9-�Y����3u4R~B��E(�1f�?DaR��M���{�>U1$�D���#�����9��D0���[f�(0�,��~�� JkG��\X�x�8�5�H"��V8�K�!��/5.��T\��������V�@�y�Y�TJ���[ۇlb�[XlxVHYEB     400     130U��֌�l��r)���TP��d�c"���̒�������� o��]u�����)�ʷ��|�8�'�G�Sͤ��c��s�p�WX���YJ��9j_�o]�Ǩ47�IM\��.�򤰭�O�ݒ��˥|�晡Rq4$;��Ym!0��8�"�����?������5U�vR��]Wy��es��IRnQ��N�9�s�&*	j��$��'$ղ����Rl8O����J_.7��*�z�|`�-����˞�Q�6���8�i>��	��˵U��p�aXIz�!�m�Z!
D���AJ	�󙦘XlxVHYEB     400     150��gg{�X�>2`�����:�5���&hh�]>-�b���2�e� ���g�V(.o��VH�l5{�Nx/p�MJ����A��)�_#�j F=i��_�$�Z|�/���(9�7d��;�=CpЯ(�h��!��f����>�m��L[$�Cbld˪�o묌�9�K������0���P?MA*�ˀ�۠B�7���� ��`���H!��q��_띏�V��ׂ�5��iU�3��j��<�O
�5���Է�GK�e������a�|H�DlO� o#��W΢������ tm4��EN�z�W#M�>�b>��XlxVHYEB     400     170c��ａ��E�ȧ5[W/�>q6G}0vΧ�6�,b�4~@5���X�c��m$az��B�DG�8��{��y# ��Ώ���b����EfX���aq�?1
q^W��F��@R��ͳ�w��é���a��x���B��Q�)�����͵�*Y4�{%(q�V�CAI����;����u�V��ۗQb�!��^}V��*S+w�>ly��D:�ְ���w<.��>�OPm����8��U�c�H���b}��̵�Ŏ �/��LT�VB�ĝ4_���gH�T2d�
n.��DW���{� ���,�EZ_�v��i3;�C���ڣLHf8�3���'�n2V:,k$H����rf�҅�3Ti�����7XlxVHYEB     400     190nI)�,�����8�E۱@Vh�o)#���qx�q��ih��7��x7��l��M�B��0�����Wtg�43�o;&e�P��b�V�-�8%�Q����\+U.{��Č��Ą��Σ]߲1�ԅh�~(�|p�D@k� �f��Ų�������K<��r�}_��,�B�#-����v�>�4������ۚ��[h5ͻI���/)���T����������^���^�<?&��t�c�A�`tK?�𩰩i��{�^���a
/��<�t��,���
W�O�H�C��I<7�o�KV�??�Ѐ�L���5��&V)݉��A����h�)nbFJp����K��7,��ڀ��g���>�!�o�<�t�����H��,<��D�.�
�"~�m�)|:�h�TPXlxVHYEB     400     180J��pٺ<~�*A"�i��ľv=����8��+�@�������kS�+���yP*Ĉ��4lh �̴�Hq(�_<vRK,
�Cݡ���*K962&����c%�������W��h�(5�?"�L���
����=!^qV�;#���.��O����r2ݑ�S搡Y��9��3�bL��I������9���ءkC��,#:�U���9�y�pqQ�s��)8����8����:˩Gp�G��Kz*@�y;E'���q0�+�	`�:�/��\_����x�l��f?Y9�O����U?��.,R�áXF"�<��]X������
�>WO�-v���7��)pgM�� ������)�b�][h�!wȦ������%XlxVHYEB     400     140��m+sM�!p��
�^�%� �zҝ{�-��{�sI�|����,S��=�a��jJFa�	����S�0a�O�|�+��|��+"�t�W&�ԃ�>1`��>~|�Z.���-(��ڮ,��"��Ĵ>"��6���:��]�T"װ��diQ)*�ut�L��.��r]En�8c��RL���7�Q֋��b7�k<������ہψ��YEF��7k�O3�ݗ�|�}��d3�*ڈ���6�w�a���?J�X�ی#��>8Q�Of1�|��e
�[6��\H�2Eom[���E�L�����XlxVHYEB     400     130EU��|mH'|y�'W�4c}�?�-3�P�ry�5ހ�5el0�˪=c���|-������=����htp	��;rH�,�VЁ�U�u��<G{��x?0�R?���п�6U_��dK)�1E3w	ҍ�RtG�Ns�E�m�F���A^@&���z���G��o  ���:?���(=R�z��x�ԛj]eZ�L
!�퓭�?w�|W�92���h�H��EZ_ߵ���l�#�,�`���7Q�$���Ct���k�H�V�����9�H*��}��q��D���xi�qX'��XlxVHYEB     400     170�c.N�+��F��>��&\, ��R5Jx����1o&=jzak���{��2�c6�yc0�_y�Y��ˈ:܄��{�@��},^C���ۜ�� l$GW�R��>!9��騝=HF�, D໇��Ax�ar:V=Ł�sV���Kt"��p��D�G��,y��&8q�l������,��ro��HX)n��46�%-M�Wbs�9��>��g��Y=-2X��'�d�?��P�&w;�3Jx�H���w��#�K�� ,i���m��k�t����̰zЃRZ[�A]y�a-��~���Y�O[H�G���8&�u�o�r���)�"��0�0]t�{t�M"�56� �$_W+���Q�m+���XlxVHYEB     400     120 ^#\�w.�F�҄n�$�J$0��kJ��c|�W^�n�=��{5��Y3oz4K)p��	z�t�e
�ޖ��Xy�s�oi�[Oi�ǤFU� ��f/ԟT �?��dw���fzU�HDh�� �;����93�N����Xن�]~)A3Z�h���c�[�tO��<n����	"ϭF�Vt�;�e��-�!R�WG�r.�ǚxp>��������l�s��2��tc�IY`�g����-�s���ߤ�ɟAԎ,Pĩ����R���IR���ɞ9�XlxVHYEB     400     130I?܈㈾ t5
%�`��� �����>��1s��W�D�uĭ8C�ܶ]�&\�"*�=FKmH"v`8~E�vTZu�';Uy]5�Dj�uAhy�/7��dv{�Q�[�g2N�0�/�g�4��r�dF����M�#B�"�k�Kݪ���[<��il2$V��2H����"�'�,ڞ�^p}�z�jT���hH}mI�<{BԄ%�/p�!�yK���ƛ|&>T�c��R1���9�S��h&m�1�Bg�BZ~�'~���y%Gr�-�Nde���q�"���֔��h�2Mt�/С�5��J���XlxVHYEB     400     140a��%],��U�l�q��(Kd}8�93�)(�Ъ?����kQ�]g�z.p�����v�%��Jny���~��n��H>�{�"��z�y��51��]_�C,��)������z?�},��8��ҽ�;S^�j�L�T]�����LL�Zň�{�����
�!f���n�T�j�����s�[���N���qq$j\}��B�^-�_�nǶ�p�2���g����H��v<�c��o'�e��_�����P7�>�<�f2�Ȥֲz�!�Rf��on-�0��i�q����s�
h�Qea��!��"�ա�z����ȫXlxVHYEB     400     1a0z��᫇�+B�gpeF�Ǹ��ǃ�g8�R�&�z&k5H-Y�B1�B����¹�U?���H���e(K2f��l�S�)��2/F����/8;��I�T��%�@R��1���aL��[~'�J.`�߅l������A<�e���<L2�ǽ�`C)��z�R�8N$'s�-�)�*I;:�-e
��q�@�F�\�s��f${��D��t{c7B�(<�Y�)At�X�K���C��a0���1�c�m���.�ȿO�Z��Wh]�h�l
�_C��k��|��oa8,ٱ̻��l�uK�丕:����"�a�7�+�?vD���M�PΎ&�ߨ�V�T��NDs@#Ɯ%��_ojr� �s�{	�����O��[ ���gh���(�D�l���u��dE��y6A�p[���B<����%�m��R`�k��0XlxVHYEB     400     180��(��5��4�mJ������������!okn���Z]=��|�5�Yz/E�~�C1Yj���gɨAر㹧a⊌wS��^�uM�lp1$(W�{��4�[�H��yT���vd�2� 媚;��Ij�68t���J�d�%{�����"��a;t^���uw�6?�|�p]fo�DNG�t��K��v�B�#������L�$! ��$�s�^{���L�s���Ы/Ǫ��s���(ZO��.��Af��nM)ְ��M�_D���l}l�Pf��M���?ВIYw_߂��ݬ��*O�O�҂'��Z�i=O��C������%��pK�h��9e�R���E�aN+��NP��v��7��~���
��10��h�M�
,?r�9|0XlxVHYEB     400     170(u��bA�`۬�~oe�����P4��o\��g�X�L�m?s#���°�F��P�;}/��w�^�g�䶭C�lx�� ��z�$V� ��t"_��;��/����A��s�&Q{%~g�g��U����6�C�{���t"xb6n���V��j�yK�$4��4�����z�s �4'k���u��'D�
�lW��΂T���(
��!LO�'���Tx~
w���N'�Y������,�}�i��lvyah��5hF�*�`} �OY�bd��ϋuZy��1�H��Ctc�#$�v4*�䗔"�^��JQ�/"��\S�;��d}�(���Z��<c��;H&�J�P�6�b=��XlxVHYEB     400     1e0vʪ���s���̖̳�������9iB���@L��gk빚0��z��9K�<�=�J�iW�/�V;�HZ�	�ص7�ѡ������ꈓS�UJ�zb3-T�j������\r�+L
GP�J��
W�qmt�_O,q؅g�F}��Ee6{nQ��7Q����m�r���DE8��f�M�R�E��+�or��+�G���1J��~��ö�wmQ͒���-Hl*���'�y:�p�4i�SdV�9
&tSC��4{t]�(�-b��4N�c�59B۠Ycb{�,L֊�+��@�4q-�EU.FrA%w~>|{)b���8;�0��R�뛓����3������\�1E)�y�I�p�S���c�k��(�c�,%�H:b.Y��
B�?��� �G��k�r}{�q�	B'���e���i��a�N.�8��)dƛz�Q�[�\�5J��	��?3�#�Ԇ �ϬO�aF2XlxVHYEB     400     1b0yOj��� K��F��R`�����C �׉��x��؞��(�ܤ�aP��V�.a����,�	�떁��)��}H�8�CF36e�`�],|��<l
�1W9�\r�%��+�	ah@��"�a+=��n�-��=3	q�ZH�82f miv��肣���\�f�q��9K�-�A�A7:<���
t
[���4��92�˾�3��Zq�oNM����Z�����9����ۊ�5�"e�i�Ur�1�+�B�J�޹��]��(��h�hν�C ������ܕ=T#Z�݊��~��O`t������$���������c���Ԛ���\@U���KF���ڬ?�zdDp.%��v�b>�C���
s�T!�I,''�C\�c��$14\Eɔ�g�}����˰�~}0R��x7CXlxVHYEB     400     160!�qӅ����z>��NB�����ͷ^<��,�ϐ2Ua�o��dxe>ݴ~!�F��g
C��;�����\`iBm�Ά�L]��~P��i�$����k2����M�!:E��=�6WE]_2e�P*_O�������a��li���I����,~��-y��t�r���m���%$�om�}$g/a��9H�y��>���b�)^�CUQv
��.i��VČ�j�iX�[~	��%�2�3c-�J��"�īj��m�dX���������|e&�IU�e5:�0s� ,��|7&�u	Q�\���L?h8G���N-�}��^����һӯzD�خ(/;�SS,TS��S�B�XlxVHYEB     400     150�P؅� 2�1�lDx`1��9�Z��ۄq���<�F<k�8�a-�j'p%��i�S�S1�g�\��H� NyI^�΃]�y#���*���!6�L�$ ٤�j�&P!K�9�!��=�|L�t��E=e�������S�q�W��F���P�[���!?�>:�p�ج�������f����ӰaAs���'45CMhD��ʸY(�pO�t����D\x�5#� 1r��ٻ*#9�I��n?Su� ���:w�Q/s@x"`�
5�ۦѥ�@"}?T��W�Os�m1�����,��	����tk��hj� �Bl�;����~۸��6�np�XlxVHYEB     400     1a0D��Z�����[|Z@�r�t�j�P���6�f�.��y~���]uYQ,?2��L�����ak�PN�4U��;#P���EgM��u_�ͣ��"�z�o�/�w��8Ի���G�&ͬn��<���窦V�X�c�P�3Ŕ�\��;إ���c�����&<�Sޟt��Ғ�B���gr���!~�^"�'raBK�v�L�e�-uA�8��
��G5L��`h���Y�� �{r�h|�el�Ȃ#5�YEXT����z4�z:���<��$��
s�Ec�]-(6[���q#t�*�a�d�F����v�*�'y�{F��ul|+˂� �!�t̼����$#]w������O�N]���\�z��A��V��{P�Y���>>�V�7�~�Oy��������$ҲW�#���N�XlxVHYEB     400     150y2�:Uk#ԭ�Y��%I�n��fMH��#J�Y�����x�2T�I��h�wR�>����n��ƨ*��w>�uy�5Ű��S�P��-����B9��ÇAʏ�\�b�.�Q��|�=y"�򈧭�y͵A.�>u�W��~��/)"'=[����5�Zx;n�D��![%9��2$q�	�@�m��
�v�E��H���2�r������w6�����f����c㔾�d�[T�Q�;�)�<��3Cq���q ���ё�x�϶a�Q�"x�i�I!�����l�����G8JN�1|��$� ��CՃ�o$�ʀIGrS��5�XlxVHYEB     400      e06����VYbڰči��:UƑ؄@���,"��0���wKT67=�j�0��^��[L�PB�YG�E�+iv�/�_�:��g��w��q*�~=�B���!��Y��;1����� $�u`n�El5{�]s��b�9b�}R���!_��d+{Іf�4)�x[�w�$>p��Q�l��1����"e%�$��O�fx�q�DP����D�5��=��CO�yC�XlxVHYEB     400      e04�����*p�N���B
��FT��6>����5�	��T���/�K�IӆM��v�	~Wk�!��d��w�:��9�j�;����bHe���b��%��f��4�6����_���\������Rasl���g�w�6,���'W��?�Ce�E;�0zr]�um�D�
�l���<=C�&���� 9�T\gg�وm."���I��J��M>�Hp�`�c|P�%n�)��wvԋ�XlxVHYEB     400      f075��T> �6�7]g�q4�.�X��*���P�#�!y%��2d�����4�&�ÉK�Ճ�3��w��V2ӊ-"��d]q�|O6B0��'ѪI@���6'����#8��Z�%+M�h�`�=֊+q#&�#5�z��^\t曑a�!ģ���F���B:ᨊ"e}�Sԋ��1�0G��cv�M+��۰�'/�:������+�a�2�t��!����Z�uD��SJ\��JB5��XlxVHYEB     400      f07H:�/�C�-� �sT���D�ӼKB�3m���3O7�W���U4u�¢q��sGߣ�����`w�@��A�M_��]lB��YE*���}�&�^j3�~z�(�j��2X��3��c":��FnQ�:r�'���zTYG���/�
��	?ó����8f�#K���;���䫉�w1�<�]�ٯ���W��	>B���n=Ӆ��V����$|H�֒�Qeܺ+������D8��]QXlxVHYEB     400     110^j���7*���ߋ�N:��LK%�_��GX�17��F�&�u��)���%���&��;��p!JW$���4�mZw�)�P<��|�pkm�C�o�H��6H�^FW�D�2��4I.g�qg���A� ڗ� �) B_��%�4�6��l���q~~U�����FIp7TBq��(sj�=�z�������]�p,��L³� �pC
	E��P\�A|�p����S&/�ALqd���u�X���u{YG�T�n��L92�k>{�|�QXlxVHYEB     400     1b0�& ���?�cJ�u,Ce��N"�~�V��;��B��
yڗ��Ϩb�+sa\?���	_��y�]�I�B?���s��%��� ����{��H���
+*β����?L{3�>��,a�GW6K��H������~Z�w���xL���7�����H�䌅%��ԀO��㩴C��č���z|�ȯT�y�N5�@ڡ�J�S��9�=k�E��ș��d'ЋfvEU C��
5x���M�u3lH��Z�2�C�t�5Dy�ɀk����1����m�5F�[	�ŗ�}&��"h��6d��9�geI	�X�eւ����
y}��sS��|���}�H�2Z�H�9�e򘅐DK�^E	��F�h�`e gk�\�,xd��`��~�%~�t�b��$�]M���m�iSI�/��v�C�E�Ns�n���XlxVHYEB     400     1400�=P�Qc�������s��-2=�C�OV\
"I���Z�tF��Tj��YV�J�ťbovH�`�q�Wvͯ��P���5�G�xd�@Vw����q	���\70 �e9Go݇����B���]���O�&8��:9�4�#��5͞���:����l
VDJO��*�����V�DW���Ts�Zϸ�f�mޣ�vn�(yc2x� J;F�	7moa��������L��^/~bm��8>R���a�`(^?�+ZN�]c?�'�.�)#��wB��T�e 	����K$�}��J��(�A��р0��b���.�eXlxVHYEB     400     1608�{�˔rwt�X���؍�uO��\�-%j�n5E��q��2�)�F�Lz�գ�}A��[���>��{�~�nJ����*��	3_&�b���KW6��a/�Ӕ(��{TO'��Ya1�H�.�~b1�<ϟ�zq�N�JX8�&��k#�"����X	cc]�ו��Τ3Z;�~Xs���N����
�p}�45g�d|�W��P)"M�����8_��1�����P�#�V[$��D�x
��vF*$6cDj�i�"0Oe��Yc���1�
J���ˉUfir�97�@C�r�U"0�;��@����R��g&��V�X����.����=��M�OJ6u�uXlxVHYEB     400     140��ΗhW8�\�Ё�v ��;�R��ҡ���8��oC���:0��T��of��"��-��% �B��Pd��f���S�Uj� �WI�U�L׻.y���&�{� %�}�h�d��Q^����6z#�9V݊��͢��Gc݈�ύ��G�ސ^�_S
����ƫ2�������OK�^'�֘o��y���j�˽�(��!Y��ty��$3-� =��}"�Gs=���G�K�����e��V�i��xzߐ5�bI�\�Ay��rj�07�2�|��hM"�&�Q	HM,�v�y[X,��&|!\����F(�%GOXlxVHYEB     400     180dM�<x��z���M:�$��Z��D�F���ʛj���w��bX�^���������*J<+G��3�PH�rIZf�#PqcރZ*��Wvl���8M�u�%f���K�3p���rS���c��^E���]�i0�c�����mؼ���C(/��-��yTd[V�b�t��4Z���~l��SB:����=+\�� ;+ζ?�`X\Ƌ ���Ǧα��d��l�9�9��K�`��k���(if,Z	��� �W%60<RJ��$���oОeov)��iFĀ���=0#~�]�Z���ӯ^g1�fZF,:� X<3PE?��%-���3�a%���V�<��~�#Ca��5Hߓwn!�9uѬ�7ze�]޾XlxVHYEB     400     190:[@�1Ǥ�Zln&��>Om���³���'��*���t�������;<)��+��|���9E�f�<e]�C��KްM�6N�?Cj�42;�\&���������g֊} �C[��My��r�=�*Α�!T����狭��E�����u^1��뫑�
e��1<��H�I��R�yg.��܌C�E$���?vG�)��e�eM���b��n����I��Vr>?.HM���j�����1������v�a�� 0kVB�q����א���2��]��#u7+�d׀��GoJ��oM�n�'��I^+�GO�O�I�$��L]�����W#W$�x��/�&�Ʒ�,�
U��faМ]�	��𑛢��m@G�5W)�z:H�˝��Ƭo��hXlxVHYEB     400     150��|'��ךH���O�S*Z�������t�ٰe4o�L�G�3�-�]GH|���L��]#��y�y>\�@��hD����GeM6���i)����A��Q��L�h�~0gIUu<R'�_7o]��3^�)����[��hw�Ş�>�v^����ů-���* ���.e	Y��3 B(���7͍Q�۝�L�W�����[�G|��iT�PEP,�q�m؋?u�~���6����va���9~�Y^���q���{A�� ��������!C}h[Ή"�6Y��
$	6��wƊ�oI�[U�l�3BA������`����̫�XlxVHYEB     400     1a0R	�$�^i/�=���
ɭ�gbe����&w�k��يۡ�E��Q�y1�횁���:�}JgB�|��n
������3CP "ɪ�~:2�ő����"�Jc���S� �)
�X�``���l�4W̰\W��p���Y���v�$��Ԫ<�U )~�{k���7�˲��H�X�'�չ2*��#r���p�?�f�9�p���?X'T�� �<>�a�
���.h!>/�k�p=��]��]3�/���U~A�hZY�vW�)r�tZ�o"��Zs�>���Egje���v�f.����W69����V����fӘ�x�E�[L��>��F�M� o�}�A4���,��k��B���4�P��_�Yԣ_���Ve����w<�F��!�]�]8 �m�T��aÚzv8��u,oc�oF 7�Ҥ���XlxVHYEB     400      f0(T������|��ސ�Q#�xrَ��r&�3�m�����1�}tİ�E������9|�1����r"��0ߜ@�N�!�4��f���=� C��#�z���`D^@`�?���y��O�h�8�c��1;8L�#��?�j|�AHUm�Y��N�6P��8��dB{\��ҙ���Z�<���%�<��t*T��$L����Lu���k����F�q�mdW���#�K�N1݉�����(�XlxVHYEB     400     100�߃�<Me����!�@����J���8��{9��u@W�Wퟳ��
+ #Ա�أ"�sr |���>ʏq�"-	�+N��ae=w��"J�_I�'���|�xY~n��w��t��:zړӴaZ�1��i��Ag���������1l�\$6$]b��xS��ߔ8�Q�#Y�U�I)Ko�+9��
6�F�Ҋ �q�?t8p����5�j�S�]:���`�W!����2��FL��;�!!r�U�B+�m*;��9XlxVHYEB     400      f0^���V��ӗ7�O�6�?��������$7`P}sW9���ev9�s�at���u�W�O񶐯���U��8Q�<&���OϥZ+�{���$��������r�<�щa7��Ы-�������a �P��2�������ʃ����ؕ��л�ؓ6a����R�x	��B��@>�*#߈~�bɳR���/ŁY�,p���tD'5H���D�~�5k8�z��?�<*�u���V	)|XlxVHYEB     400     120��ʣr�$��6������
~�_"��/zH���\0JS]�a�����U��Ѵ٭��R��=ƴ�ض)0�6����Q�1$`�e����o*r�6c/!�ي�s�+=����Z��c� y	�<U�����b˹ ��A2�G�E����	~��A�f@�g��xc^߰� &.*y;��C!�{v�*2H��:�ޗSk���r�{��eԷ�,͢�<�I�:qW�s#���y����-)��}I( '%��ڗ]#��[�SY��A�^�B��e�g������XlxVHYEB     400      c0����j<�~�m���лpt3aä P��&����ۺ��9���&��D�$ɽ*�0<��h��Nj�B�.����#����.4e%h���lBx�0o�3����q� Kq�>F�t2�d@���L�9���Vѱ.��K�0�j����Ҏ4ܨ�')�,"��m�&�3��R�[ݾ�QT,T�ZOO1�XlxVHYEB     400     150�j�N*F�AӷJ�#lܻb1dh�v����nDx�{�����wA���:Ȕ�7���ڵ�Ru0Do�Y����<��"U͏��n&do�[Չiɚ�\N\(�[�6j���ܮR����s�)������֕ow����i������!<���N䆞�vCu�d߁=�Ig,j���-s�	�(Rv��64�Z&���Ty�E��c~���aeY~/����,}:�zj�}E�KA��]�`�E �24d2�Ko[�rTs��S�V��*�y
2�b�ў���X7�f���`x�%!� /��h�,����ɫJ1�ޝ��񶇡ؾN���H���H ���XlxVHYEB     400     130HX~������(6�E��	x���*���V���.%IǦf���c��1C
�� ��U�M ��W�ќ+	?�"�����b�����${��_����V�V��?m4GM�V�����u:��
���M��GN4_��%���hx�'�B��� up�s����@�uj���N<�� N�i�����u���a��Ƭ����ҹ���{��h~~�Q�%=0�P���.F@?�MjT�ѻ����C�6.р�Bx�T+��)k��	r�����p���O�F�����H9�g�v~� �f	a��t�XlxVHYEB     353     160ژJ�,�mv-���l��\>��h��G���za$�>|����֓L�:�gO��<���//|�o�\/ Q�3���H���nۈ$����;���8çE��h/s�m��O���I���e���!mhnw� `�<���u�	&ي�޻�L�*2�p���[��.����T��Yp�6b~�e�S��Vp�&�_IT7�F�!�m��:�D�����Upւ��d����,^�F�0`�X�T��PZJhS��3�u��i׭t�9���_�D��GՙX��#8w��a�zNai͝�`�ܣ D&���r���|Zg��4c+����g��G�-k�p�է�*�ib-G�