XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����������~f85[�}��9�NKh��#�}�>hZ�`�X�����iU�!J#�H�S�7�LK�G�?�n~H�af���#0.}m�#��0!uA�nTh:漼�$��Ԋ�1�n$�i虜#�AF��W��Y%�����lP����=s��Aq���@��Du�`�� ̄��}��,'�IWi��Gۮ��i`�K����8�Z��c�Wڰ�y�y�N+�c�Zg뉴~�E&��G���a�g��,L���p�.��aR�|�Q$��n�lמ���67UЊ��4�s$U��$���3��u��e�G� �EѤ���t*K��q��>$D�j����Z,�P�:<�%��:��9�"�d9Ĳ  2M�ܿM�puj��).����"KZ�%�`�g7՘��Bw��'.���V�p��٫vR��ٔO��J��Y�
��3��깎�cl_.6�H�������s���0ղ�R6?����M�j��9�\�Pn�G�%�/��QI�^��m�&&�ٷg�S.�l{�"׈��Ŵ��c���A���A�r���OĒpi��I��'f=cg8I��pG�NBK73�&Bk�x#U6���}��Z�V-�[�X�m������(e�#4��<o�f�agW���CmD.ى�h�����L�D?������KN�e|�+ �|��=#�ۘ%�|eW�%�]�('��LT�NX�S\*��+���R:��V�lm����|�%��2᪱�#���V/G)� k�g�$/0?wl��4� XlxVHYEB     400     230.O�=�"Qq#gt�bw:h�d1���x>�`�uX�O�.�����y�[�X�X4N2c�[��+������"c�\9ٹ���c�	X��M��P!�h`�<�'�M��e���E�5�+%U\���5���	�V{���"N]7UX�mxGV�
����(�g�a����&d��ֆ)e�]��)~�g�Ee���;�ds⡗�ݷ#�Q�~0|�t�=i� ��V'��à�dr�;b@s~A�k�w?6�\�~����̪ӫ �6{:H$�Пͼ�P��#�yW_v���,�9BL�}IP!�K� 8��q/<oY��9��m��U�����מk�Q��"�2�_ܳ�ix��ֶX���-B7$�{�N�*f*�++_�/?���^<=-�� �DM�L0M�yN��Cb�?i&�B�c�i���l��x�BB�.<��EkcN'�-�7n��1*��Ֆ��W��p�-�M]����qT{��5cXz�
��dXj��9���ܟ�;�y شw��!�t l2-�N5.  Kmn��>\�GD�!�?�^�gXlxVHYEB     400     1f0�ھ��k����y�m`�N�#�1�����e]:$��kɠ}V���:��^۵A�WXx8:&�w�Ccp���3�{u�Є5�w�E�I��������9SV�K�ʑ"]�/"�]�����l�JOx>�*�����~�r�hVQ�U^�G���c�[	w#��T�3�����d�6/ o������~�]�B3��RK]egB��"$s�?RD��=H��F�\5c��s�'���϶��C��Ɖ����3��ⴞ�$zJ@�u8>�g�9d�->�.�(.�g웱�|`��3r���? �*x$[�<���r 8���=\�%�
8

��9�,���k���2���VN ��O���%O�c[��#6�M���Y�L��トo��±�H����������(AĄ�v�۶��j�$��IHt7W�O.�]M�Ւ9?��l�7S<����
���Q��F�R;}�}!Wp(�}�-JP7
ěJ�KShXlxVHYEB     400     1b0����؊,����(���� �e,(�����L�t��Yۏ��7d!�W���?v` ���.�ί�,N�>��m�_I3�r8z��֦�D\�@�c����\��{i���V���l�Sϗt?�%!�c�-�]'����*Q|/SM�A�ڝ�%Z���l�{���uz���K4
��Ɠ��l������j[�3WKC&�?�
�L�z���ɰ�,N �.�C�ZQ��N*��,�CR�Y��+G<�����-9������|�N�fO��'�������wt�d�z���$�J�.���� ]E��"��4"O��ǼKnh����4K�bc���o�2�>K���MVB���_��^+�Z�b��
r�8Y��p^S��|�q&��A�d2�!>�*]�5����������-���c��z3*�XlxVHYEB     186      b0���1ͳ�P���� Z���xA5W�f��L�N�v��j�~���E�~Q��n�|9w-� ��\��}�tE�Օ�L�acZPڶ�zW褪���q������x�W�a�
�:��ℍx�Ŝ�P�X��)�)Yg2#ѳ��?�MU��ťtb�ȢJt��9��f��2ĸ5��m