��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���L�n�����68ۇ�fa�F. }?DЄ��ٜ{��Hz�(�-�Z��k=��n��R�5���K�:��.	���S�Y(>x�?��6�e�Q>�����ӛ�;�;�3�iE�mDS��wbp&$��wMθG�Qb�
�[8�y;E��B�sr���K��Ċ��st��5��΢uR��4�|���x�.G�F^��y��w�o�f�l�dp�3��@;I�^)Pj]^L��|c�#Gt"|Ж�?���3J�'��c9�����&\� �]=4'����(o�C�Աr런�UfYh�@��3M��
k�e��:|3�אn�	�����s�1B�I�g�p�ÿM ���V���!O���<w���?Н�U���=c����֟փ��3b�_�������1�۟*�{�0_Л�+=R7m��g�Ӱ��|��yL�to���@wh7�u}�A������"x�ʵT)F�I��,�6Go�mWؕT��62������&n9<��xoI�tneF>Wb3��Zf�*I�����=���_��.��QmY�<�!�g�x7ΰ��º.)7�/�.��-�i�������j�2S~��R3w��S〣���<�Č5�ޞ$thK�ΰ�{fC�_�N��&���:���� i��x@�J�=]�E�T�'�Z��4�w�a��q�SA3��y�������Ӫ]mO�^�h�8H�}��;щ��� �m˶�q0(�?1����]K0
p��7�b��j�	?G2x�ڇ��u���u�*��4Ӯ������~d��h��V�s��v��ٔ����|M����R���k�n����u'�g9���}�ĀS��.�by�ہZa)��X��/#��Y��R���kv���|&�}�����Bř��.
�v�8wS��_I�,�0z����*����=��e�M���wT���c�܄('�馬'q�8r42��OZ33!�ԃ벼Q�#;,#?��~٘��6�Ÿ�<9۳g�YK���M��lK��ʙ���V�ՠ �y���;jƤ��e�M~���/��j˼>��ߎ�����s�ª1J����˒g	�5m��BRr�!��~�Չ�z���� )�"&eko�	MS�x�j� �0�����~�U�zɻ���*ϡ���z����;�fR=���,!-�F����'�z�Q˙�޼�=�u�an��m�|,b�����bS�24���[�E8��k\����5�%f��}"xM'��@��]�k�g���ws o��*Dp.)����j��4x��+Kv����;����%8�Gg4Qd���\����J>�,ވ���V�!��W���Ji�P�����W��Ʒ�`�oB`��jO���2������wt�������M���c8���x|EL��wۋ/�~Q톲�1p<���Ǆy�5L~��@8T%�F1��!	�)�H5/\�"`�O=�ԊH����r�>�݃�8_����f]� ��j/�!u��̔�T�{ �f�^�We�@=�1�[(,�@d2�T��n�����H��T��]�v��%����+@§�R
���Z=�	�h�����£�
h�sQ,�<f�>����k�Ƒ�tp����	�a?R��(1��P��&�H�K�����Ŵ�q�@4�	��{�G���|�HC��m��}��v�C8���O��Eu�k�Vy"�*�ׁ�5���"����@�1� �� m*H�6����?z�%�[{pl'��;[i����X��0ѤjQn$vZ��*;ƕ�
�X�_t(�B��7�M�����k�����(l��u������ÿ�x%��{�'N�ʎQ�/2l-���%$6�Ä�:}�)]�O�g�{���V��ʸ�͌��)}̰k��+>�懍� �	�)�=L�����m���_�q��D�+���̅�*�����5Y���w��6��`��YR5?&�&o�8�P����*V���sƖ�F�d��Y�]%!r���~Z��>�0B"�u���M[��.m�H"w�T�a�e0�(���|rn�ߓ�׸k�A9���Z�f�� u��iS��������CJh�:�;O�/�)�.D99��q�+Eϳ�
����K|g���}��E���R��jK>�V=�7l��`���Pt��`Th��ovK��3���$�aJ?�y�hAbr���sXޚ�f�E��b�r^�}s�.�r��Zx���65w�csfj������.�z��q
t�q�D�d'%�Rv�p\�~T��)>���w��;q�\�2��.�um�_<o1��g0�Լ}�$ȶ5�1v�n�݋k����7�fJ��w��k�w�)�q�+4��9��)aְ��EN�����WP��\"6��jtڭ��\>����RO�D3B[|<p-�{^B3�d��:�k�a�?hj�S|=|�y�Gq��]ȇw�4s���:N���u�T`�e�4Y� ����%q!W������n���E�ۍ�˻�w.���_�TX����|{釪k_^��}����������_.�����^�D��U|1�H(n΅�<d��%�3	4'��J��C�ʖ.����PX]#.�L\X%�4{S6�:�+��ei=���D���f���͋Z'��sO��Bno�p*�2�X�䗣����s�6��d���5�"�BԈd����$Ð�v�R�d�+uL"�3ZU�,�2�?�Z$���W-p�V>�j�PV���v��U�PۑEWM�"#rS��?^cO��C|��@���2��';�9�s6pv\z�L���^���	�M'��X���Sǯ��$�ΨlGw�մ���p���+���c��q}-x9��g�1=�|�І���L��E�
V�Ś�������$P�'�x�4~Gɡ�O��W�"#��!P}�@�7y�D����+l̿�9ǝ�Gg�tA�(r�}�Ү9��b��@��z:;Y�����H����H5�	�A�ڢ�%�)��c	�OI51P��GC-�Bȕ�(d9�)m䐺�3Lr�HmvflY�U�I��m�T��%S�>[�/��A�z��"�ܸ�i,G���n�*��+�ц��rc��é�e �ըPl�K@O����ZT�4]ܵT(m�z܏���hy�1�1�WD�7���	�n�g>��P�X���$'��aw�9�4Ƨ�D��E;
�dC8��+G�֒xy��)ٽ� zL��Hn��[�8.Ũm���`<���I�t�ST[|F�qj�����y5~ꔔ~��?@���� g��h�Or�v�׈�L~cuG���5ˁ�����A0Z�;���i��D�A��^�7�Oo�V<��)~�@%ᘏ���:x�o �ڼG%�vjt�����b�{^{���0��]�_�:����\H�gL�(g4$〰��" ��~z��Pj_a'�׹��Kc����f2tyxv;d� �\���9�"�~��LJw�(��G�H?��ҺG��W}ey��Y���(�
Լ�Ԁ�Dףn���jDN:����9���!�To�n�{�Ҩ<b���E;X9�a;��1RT�e�{kJ$�p�i�gY��Ze3V���E�����bA ����������6�'	��3�}~�qX+�C���7�'@ɣd�\Q�|����J����6'/���W Ne�Yۃ�y`��}�M;Y����ۀs7�+̪�l�֯�<>�\s�$F�I��Ѭ�:Q���?��f�/�r_�;N2rw��&�S8?��R�t���خʍ�Y�dU�<׏�e~�h)���]{� t�_�� z��s�)��]�!a`��X0]Gʼa��$�<��i:���~��v�՘fC��eA�rˋ�d	S?>-���0��R��2 f?�����	-�.�e�q�$C�:��@
�yU��ȹ(�b�e���<�(\ĜPi��x���3B�䪺�ʟ��{;0� ���
gU��q�?�9�s �� �ܶW��0�(r8M`���������ax�x��cW���&��H��ս&�V3n� 2�)����F��P�NP��-�F�2���d�:7+����o�Ssf�/��*:��(| �3B!ۊN}Ƨ1d���H{@b��mXbӅ��܋pW���Ķ�D��Q��xa��Ar�Ï9�=��c����7�B��W3�kjݮ�����P,P�V�ҝ8+�꒤�I�x�E���-��C���	��8�L�M�ݞ�7�7_O'�������z��d�M#0�vҰ��*}�)������+Lj�i�Y��1}Y�5���˂�����M�.��[q)DB:����#����c*��A�-Z$�5.�zA�t���E�̥��N�u���Fsh�So,{�H0mM�c#l���I�W!�<��o��ree�M;��Y��_Q}�3S�3�"�$]Y����Zg���#U�T����d�Mu��fS� ��#������r�~��@>��Ez���_��i��9WG�6}a�=J^5�Ly�5E�h�v�<߾V00��a�=�Ւ������/4� l!(:�c#�q;��HߋUB�毥f+
�$���F��?�8���p���' �;�Ϝ���)�HKݸ�,�isN�=�'��I��a~1z�}]��x�֤�&Dqʖ|BS��Z���(��y��*���[�@��f��tf�P�-��I!R�*s��������"���)���q����<���(�����< ���	Qk%���K���7���J�v��o�Xh��`�i)�?���I��j�
CW)~~��1�,M�覺F[�+1l({�>�z���������}����uz߈�.H���]c[?Ix* �U�I�0E��^�p���c,[��M/�^��_eN���j#uK�F��f���G
Gۑ��'3'x�������,�N���Pz!`��~]���^�ܥ�i;�t�5b��H�e� :�e�mҭ����[��&��E��!����h鱽I�Yj���r�����Ϳ�U1���@� �c��FiO	N�[�S����:�x��;�z̍��1��>�ѳt �RX2���C��p
MDq���$)S0��.|Z(0ǆs�u���K8��K����������%��E�?��d�xMdd\��ʼ�6	��Z��"�(�9J`:��Ư嚎�=2<Ff^k��m�?�A�6�w]�1�������b}��}���헯);�)~���Ŋ�5�I���5�i�PU�|�Ws;�����<�g�:ݳ�&�޾
��\�D%�3�@��U���:��h�H��a[9�r���\,��>��pE�O�_�a]  ��uU�8�Pe�>��H���)/�Xd�Q�8��A���俥�w���S�m�������3� ���Z�}�������,��Zi��ն��ˮ�3�[�X����n^ �y�D��qgt��rU��e���WMԴQy��oF�;����@'_;U�^�d~�\X�=���B�g���ђ���xè������| y������,�����&몠���Չf����r�A��+69Eu����2*㼝c�>��;<\���\�� ����2oJ�2fﳸA�1B�W5�99���~��;����k�h�Ē�³�}l���G^��z�B+o>�[��te�u����y\�/p�p`Jvbx��?E��狚��?"١ފ���'��&
jML�M�mP��I�aJ��a�1��"���e���Xۅ��l7��H9���~~iHɏ6�l���}�����ɅE ����0mw朝�����^��fAQ�~�p!��1�9�|%Y����I�z�xP�jh�@.F!UX�NN�P�T��;��%���DI��������]G�7O�"���L�� ç�l�m;_��!p��`U��=�mW�����:�ts8o�woZ���@�&�� +��t��<m�^qִ�<.��f���O�&��i�[�
������Q�t�*S7�^��Z�7�Ǐ�v���&2m�����̈́��3�.2r&����#e�r}�'d�D�L�dƻ�ez1B�l���n0YC:�9�8,�+�[��IPv���J�G7�`0EÈ��A���n�#1��ر3lx�<]��z2�#h�}������l��3h<�Yɜ�Nz�A���O���Dv�)\R6]����1�T[��y�Nʓ��9Z����X���(��q�]�����(Č�����F�K6�x�[����i��8�24.G�x�����[���[FT��ޖ9���m����FR�wf�u�Q�~8�ݤ�Q#E�D��b�Et��.�1�-�C��
�)�aϭ7��f��kmɕ��8MV���4�G#eh�^�����SG�I0;��	P�s#��[��
B�����z�iq��/��=n��3�A���C�[䉊�&� d�>�#z�c���zC���}�7V$7#[�D=hi9ew������� V��+4�}=�pKqVT��öz�&��������7�3q����v�Ȫջ�J��X�BCyBJ�8\+%�'�}��E)���o�N�`e�Sz�f
�m
K���%A���:�����>�/VF��= #�'�3�Z�'��P�����h8���2U�%��:��5���R �bYD�L1�1 �|*�m��ā;��|��a�+<�W6��$�^�'P�d��wJ9���<���Yr��=����ņ���WE4��hԡL\��겊v��f)?��Q��(6A� w���u�VRѫ��xPs���" �l�?�Q&K���ߒs'�@���
�,Y���4`!u������%��3�b�(���{2��O�2�Ǵ��q��I��zd��P�X�y�%����8 zB&���ƫ8�=ͫ@&E��������9�H����� �
�}���R�%.�A�:��v��8�w�x�ߚ]Qu� s�{2{D��/��	��v�X/��E��2�5ך���q'b}��N9�H4𧡯�%=	�O��By�sx
s�Ue,�2n�ҸxŎ]v~��a��C��*XR��?���V�^d�� �V�)���rʚ�y21Ag�P1�=�`ծ<l�L���1��ÅK﷤�(h`�i�D����)�-�=VT���3��!*n=���W��f�j�g�p!Z㓿�׹[�󘽭x��!��;H�}���cĵ7��x+c��Ү�6��ύ��	��x<���o����$C��n�D}��6H�&�t�����i�sl�K��e�J&`�3�D�ݜh�.��qLfe�޳�e��A�tL�S@���n�N�.��2� �p}J�e�sv���c	�r�s�<�����r�O��n��c�hC��4H:��W@2��� b��Y'�'��^�?�Vf��!<��<�dG7��0�
3�ɩ�t�bt�,�8�P�ar	�����L���)F5�b����=��Y�=B$�hi�6�"�I�*�u��<&�p,R��d��`zW�/� ��!y�мv�l���El��*�p�k�]��-J�xb��4,4�o�=��O������͐惒T��
e�:*Z b����h7@���]Cz�;ɞW��CJs!X��~9z��%t�_��ˉ[r=Gٛ�	q�]��#�O�Z*�/����	i��>��򋜶�|���1ǹ��4���hao��3�� ���
=��ٰtg����Ud��
���G��BI�u��><�em�b]_P;ݛ��Eh�5Ǽ��a��>��A4(�����8�Y��Z_��N�cB�tZ��ÂJ�g����C�4��:S~�A:��ג�u=;�,��0П��n��K����̛��[�9͍�/���E儂1�K8����B'���;%�O@�hD����9�Ng��k��-�=�]��9u��j|z ���?��1��֪�����v�G���\�0�^i��ġzݛc��-����c$�[��9���&Z���h���/����NH%gh6�A����!q����T��GR����v��aS'a��L%�a@N^�4V"H�J�i��4�/�Q�Z�9�qj\g��i|JT��� B&��ҔX���>b��{�W����$�!y�p�r�q2���y�N<v>
��f��J�d͒��"����mPߧbl%Y���ג��m�"`+�S�Խ�6e2QJ%�ߝ)<��D��nIБ�avo���qi���%�sQ��~r�b��.$���[Z�`xE2��j�Ҳ�=���߿���e/�=������r�����QSo��y9��Q�/-:��	L�uǗN"=_�14\+(�z���b��/Y���v�����[�@!!�>���2-�}��A�Zr��~��屩��+����Y{!+��D���C�8��X�����xBU����G�$8;�(���%�"c��w��O�sl���6�ګi6dD�����"�H�eϯ�))Ի�'^�����c��(��|���g}^QGgQ?��v � ���_c0
���Ą��%O/�T}��i�?_�Jyb|�v�f�Ao�v��i����	ܣ�M�}�y���獪S��0ڇ�!���g*�� �?�q>1�Q�DӠ��i�'O_kə�L�.�U�a��W�$��閇,m��^�ߠZQ�3����@���4Q�l���0���k�xa�A����<>sg���8o���I��äõ���UEs���~����(����ϗ(��D�����>R%�f���TO���	�h�QL1����BP��h��.=����G#!-I2�[z�(�#�>�������S/���^� 
^�}��mR�0u�x����'u��#IN������=~^胲d�`]��E̴>�o2t[�7��c�
��K
-�-�x��q��$~�J"�@2�
L�˽h�c4L&���qu�GA���.x��lwg�v�01�jGM7�#�7W0�AP*	�:�6��q��;�Pb@����Ƅ2}*/�\��`@�����<0�a���@�X9K�u�l���1�T�����o�D��?�·�Maz�����?K�����e'� �W ��/e1��*��BQ={�'��|�Dt᣷�=)S0�`�M��Ლ���n��K_�1���l^Ž��p�O��~N��e���T\�1��/`�"�����C��j<
!��}��d�
E!W�t,=���$�^ád�	���%�)���U^���ݙm�T�����.֗����P�Wam�0 ŴŶ���'��F�u�Ƶ�^�+�H�5��
�*b3E#�Bv��MJ����,/����{(���ax��>�a@�Vl f:$��J�p��T�Sj������E�7��	� L��f{/U�[!7�:ž�_	:�+��Q�� �+E\a���� 1
��	��uDg�#��k��dy�[����Kj9Ś �3���N�Ry�����aZDk. �k��C�Z�T��������-I�w��Nĩ�B^b�6�l�� F��������LZ��1�2����
����$�Wߞ�C�iYɈ#S���4l����!Q7ʒl��{�{2EnJ.Y���Z	ˬ�7���C��Q���㏒��1���U�t.�M���F`Q����ΜܾӔ\o+�M�3N��ދ�8�]��^����bF�?F�*��Cc˓'K9t#���� 	�h5$)8�g��w,Q="���c7��z��]�,y6N�āsQ�7���3����K�d-�8���@P��/S�o�G��1��X�:m�cw�ۈ崚��u��ro��4#�"�;��o��P�\�q��S�q?f�J�))Nu� �H�B~Of<K1H
��a�UB͇| �[�6�ʭ�c���O:�>!�.>_�J��p��laog`F3��4��?0 �sfU0��
�/Py/v$����tʩʊI������ݬ+*���JE��t��y<V�ϩO�j8u ��ǋ�0T�����-,K�Jk�}5GLZ.
�K�=�en�I������MgҨ�'�B�|��%��0ϧz��X��a�^^�4
S�W�Kl}wWɽ'՜���)2�hb��^�����&�^4f���P�ƞ�""Df�7��*xMU��`�z��^�)�/��%:�@�'��/�����H��"�V?:^�G*$`��5�?(�Q�?O(eC_�<�S�'$W��S,�"'�:�|�fjw�^^9���k��`���	�Ú6�-:�W"?�}��[6dĚO�kG� ���$O�_�X8���WS�C����[�g�QNG������V�5R2�M�����k��ʨĳʫd�{@�%�l�W�d��8rUo�V+6���*ƙ	�M����8V(�_lۧ7f��#T�w���N��x1}�#2*[]f����I�RMZ�L'ZR�(+�A&����wS}h��R1v8C����Yi�`֡�˖��|#�1��m�xʲ�->�
<h`�q�V4�|SNTZ�g��j'��R.�B�#;���`��80�����v �Q�MD�Wr5�dtč�5E�7X��~���f ɱ��gOJ� �����;�0|k�@�`pK�|ٱ���7/�TU'�o�>n�0�_[�P}e�g#2�oi����� .{O8	���1W�H�!����ZG�;�c1�8��g���n԰D���$�g�Z펊op��|EFs�Ņ -88
r�=#����r{_}�8�fr��uYUY���Ql�@�]4����6��zڸ��2��2w ��;��e������Z���+�A[$o����=_�lr�]�������*���N���8�����κC��h��)��ȭ>-���n����jlds	�u��_�U��/|2���z��pO�RRD�V��,k�HH7r�-�!v+D@�v[R�Yjqjq�T���H��1K��|M�#ʇr���/=��U@�HT���"�^=�ז�p`��ѝ��J�<}�"L��Ru-���К������1&�B/����>�.�2�D�*��Kx��	=�Pb�&�I���c�0 C�J��X�i�xNg{��Sf���P����d8�HF].TgO�R���?hͥNUh�A˞V���o��{S������F�6�C��ze�E/S�6�ˮ���{It����=��b�ı�틜m
0ϗ�!@�v\�5�y��)W=Xф�]�<�to�J����r�����+Y�l/��7L��cY������.�n�uP�Ļ�h��;�(���|��kn�f�~�@&�L��q�收9t�=�����c0������E�Q�o�7̆�ր7S��#� ���͘��l� /��
a����G����t]_F�:7��5����6�J��k�N�i�T�4�r(n榝����ku�����8Z�S�t�qp=ϟܳ��t6G�	%�9���?x8��J�#6���-��3y0�#L���ѥ�uzC�l��W�yj��z�;|U"Fu*N�˗'�v �5�6v6�X%2��$���B�#-ܥ��ݷV���7�(���C9#�&�ü�&�s�j�wM�?y4Mg9�������&���_��6���]��E!�AS{DG3�kbWI�"��Z�{���z�^6��� Nh��e�d
���̸�� ��ڝ�W�
�ȻO9r���7�JNFc� ��ac\섩��t��q�������{��M?����):�?�2��%��M��z�v�Օt��4���p���a^IK�u"�b\����+Q"%v�˫ͼi��7�pY�<�g �7��݈A����)�;BHRS����_���@���$�����m�c���>q0���lή mx\S �GM��缏b._tC��-���*��%�"3���҅�*Kx�+Z*���F5�V�Ln����I��S7��ۑ�Sw�tf�ٺ�ʲb�@h�)��|���_98J�;���I;�?ş���t�ܴ7!�r�+22-_7I�R
���a~���������������$�
�J'�{�a���QmN��Jſ���S�Y�T`��f��{�Y�E�4�c"��߮�!q�z`�H�k�c��k�޻۬77����)]�
/B�e�^��A�W]
|�0�/��D�q�Z`F*+9�}�31��X[V��|��
(}��KI��{�t�p�����3��gU��(H��+剪\ND�i���[�U)LR���Fחv����Nm����H!#������gX�󾒂��0��
�QψE4Z���LT.���5��U�ZZ����F�&b�_Ƙ��DW�6u���~_O�I���<�'j�����i�,:D��I��4
���%j��2pw�W �Z@Q`���zd�_����4X�WJԮ>�f7�b�r�`���q���aW�T���������lP�+���=���T�Kg�2��&��o)�L5!Tߕ�uI�bޖO���S��{��͇� �/��6��Z��jF��ǻc�Ӊ	�ǌ�� D˝���f��@���x@�Y,w�A{��z4�cه}��5���0�AĆ�jr-s_��}�/᧟k6�k��E���m���;x�$]��CI�x�r���ר���R�w��*��'p���Q��hq�zOĽ���A�C��4�9_'`���z�z1êi9֖9c��_j��	�z�=ǎ��;��n�N�CTy�⮱���Ͼ�bb���g$�k�&�]�� �+M�*D*
���6�\�ڥr�s����͘��W=�e}�8���Y?YB��J�u�Z�H[½��0g��cf�t���U�غ���H���z���??�|M3.@23�Z�x��]�	!��#2�w_�<Pȋ��A�"�
��^�*�����+3w�np���9A�
�8P3/�$�0�s�+��2���i9�63a�� �����݁���_�5�����1��!�a��<B��4IUu�:����B��-�`mC��v�x-j�'��B�e����Y��뜍�&��C��dv9�����9�}X����,cM��x^e���
�ꂙ��ō��Ӧ/��2�l)�'�Gʹ������$�M����!e�|K����;9HHKpH���o��L��icy���3p[v;hZ�E�X���\��ⴔ���_��t+'4?������j�-��^'�����ѩ�����]7����T}�a���T>��+~Ɍ��(�t���$)c7�"3nAw�i�+0둬D$_��!V�	ū��y�J�T�r\o:��{����u- �F۠�fM��Ud�X����a��G{�[f�G�s���m P�H����uY�IG�xq6�;�ZM�`��䁗�j,w<���Z�˛I�H��UwZi�k�؈��ƃ� ,�)U9�:f�j����O ���AZD�7k�7����*�^���rWy������
]�4K�v4���c�zY�&�hP�3#�Y /b]�:�ǳ�'�`y`���{7�U^
��#�Gn�407$��N禤�I�~r��#\2�UD�D�u�r�ہ[�9�@`/o��9
�S��,M�����7���Z�4Ŋ ����*%���Qao��|� �7�;�5))y������ cme�G5�'�
�DT�zt�Ҕ�}��������}��u�� �VT҈kP�ǙcR*����qJHjȗ-��T/��->�_S��F�sC6r�[!��T$v�v�b��� �"��8���n��[�m�O��q���u8R�dj`C��S�_U+�������Q!u �@������C�S72u2��8m�.�v��5@41���=V�
�I��JL<?B�\�~_��"o��x����gl���c�PGo���p/�A�67�����oȔ؃Dr<�/o����'��q?�&��Oy4þR�j�%��񝟿;�zG��؀�ׁ��_ͫࡇ�.��<������N
{:��Ԡz`$�䳍V��u3)a�n�uhR�kT_����0��غu`Y���TЪ���ڗ��25h�)S�/h�5���V�)�z]8�t�~�F���bRSL?��0�E^���Lr��ߔ������pe���o��=[�N��;% �0�s���|�R[-̳]���t ���>(C+�T]`I�}�T�`����j�T#�{_�9��t�/�v-�h��|R���hy�p(�����p��0'��Ï��R�qa�Di�� a�z�QD�OSߚҕf���̢ \�����tn")3m��}�jU�L��I7׉�D˜�+!�h gT�����ck���3<>���&m��_!�kCo]A���5oVΚ�T0�m���[�fdV�B<�H!VN�0�S7��Z��@��Po:�L��D�9IE�Λ�׭�a����$����z��KTN�VM{���'ql5��T/�(�K�(d�ۖ�x+�2Q|_��]\�S�Q,r���댋��P�w'ˀn�i�94�t��0u�/	"��p��#�N��kͿ�U�%�>�Y/�O�A;�v6�7leCx�`V+k����&I�S�@�D�����#��R���nE��)��ʓ���U��pb�{�f_����	
�e���F$��1#!�<�.�T�(�QC�:�0VW�j�Ė("��ɝs���Y���h�2�U�G���
��y��#��w"���j�.r�dTj��i����I��$��`��")��K.�9H���naZ�j�y#�Bd�^ 8:a�#��逬�p��&$^�*�����[j��40��u��l�*m�Ԃ�n~�=X�C�+D{{鏨�Ӌ/��T֏�¶�W�w��#�W��R4P�1��%v#��{��;D��Ч<mzc��7�s���|���XG�����2˘�W`4U���\z�
�^$�`r��T��� l7dH0~no�����pd	uF�3Ќz!Thͻ��.��M8�o�;;,��:��䶵�Ήؚ�Tԋ�<>�5��]��Du^\��$=9�\i�H���4!	�t��J��"��޾��2��� �h�3S�xN�C�E[�`��e}�q���ԑ_�I������> ��l�3a��D�q��FJA������R&�q����;��hU]M$�:�? 8+��W*_��# ύD�; �WL�W��n?t�d�Fbc�w�ާ(d��P �-e�W. fӽ�Re�'kk���cTw7U��K�s�|��yR�d�{Ϣ���'_qa�X� ӊ�҇&2+�YE96a+�d�3��Y��3i)��P��Cx푇%�
/�5Y���a��"����;\'i�g�W�h���p[Z����c@o�(gir��e�wGH�UU�p`+���{Luw���o����*��Dó].B����z�,���3th�Y*�C�Q ���a�_����[��s�JG�߈v��랢���*��}���V��s�k��	�j����	+����x������O�bNgS{�O�m՜0?���A�[�"?�۞�ͫxo˭���o
J��,)����6B7�9٢�p ��������ۮ!�R�Y_`� �\,۪����V�d1ԉ,�Е±��D�U�ۼ��	�����fM�{�:fLÀ��6�<'N�	hoE$��y��uhaE�b��P��F���(���G��;��e&�&�5���1�<����W����\@M�9.��F�9K�j���!���=���w睺��{�$+��	B�kVف��Ɔ�����~�☩h���s<�
�j�脭�]ht�@[������^�u�!�򵐃OgZ����~��g=�U���@5E�[�F&F�P����Q�����T�.�hf[W����b.a�d��(!z���l�`�8�A�hI�?�w1��
�p-)<0h<��]txno������"���I���.��AJU$&rrS^�*��_kv7�n+ifbBqĉprcP�V0�b�ǒ��D��[쏾O�y�D�M�|��t���n�R���쐀^�:��'�(u�JU1\��<6螙NP)f(��/��Ű��p�%��t�H�P��M�K6�$W<���T��F	+N�08i�$A9���_7ёlc0��vB��~�:p	�f������[�!�>�B��c*F2�����6(����O���K�pO��=�ד�a��5@oN��
J3�p��Jk��2p|-�^sL�#�G7�п+Q�_G��k!�[[e���K���I(k��E���c���l\(2?"I�L6�]�IrY�4�A���dݼ[�J5�+ѳNO�4�;�z��=7DÂ�դ�=&�$���/I�4�b�X���a�|�Ȋw��BSC3�#��X��T�%�hl�x�/��꘳N��W�V��Qx��<Τ�q���0D�v�(�f��Ku��ab��U؞��V	��j	, >�8��.��lf[z�E��Q�H3�np���T0�$r�K'%��<Q{>�F;��)3�a��Gj�rBV��#�̿&�.��q��p��t}b�Х*�l�0�m��A��)w�k��9#Wt,���M!��8D����U�|ī�PS�`L�K
��Ǡ�u�\z��X�F}�ֻ��7!���a��'�|�F�w�N9K�}W!isD��A��%�Ѓr{����
 +Ih!�!���2�V���%o��8��䎪�O�U�N�SC_����"�7N"��Aӕ����6g!Q�1f�'�׫?+��n�}=���ҡ:p#*~9����Gޙd����C��&qE�MO�"�@y`MƫY<O�KZ�ֽv�3��Fz����\cE�|A;{�o;��@�<��������)�X�qY@�#YD�rw�e�&�9.b11g:���%s_�ٰ�� ����+8!L�^@,f�����F��<pQN��C����)�SZ*�ӫ��_��JYw8�]���^��E�(�H����6��]LqX?�lŭ5��8n���S���=��i��#���̟ͳ!Ãu��D�i�ʹ ds�V�����#���@�T!��o-e��D��;ČL%�¹e舥 �T����*��+������	.�YG|�a�M ��J�b��N`GWNR�}	'��*,E�/��$@��*>��C���w�S\�{�U7����z��9����I j���FW;A���M|��I�S���* )��3���҈�Z�`W�CiH�yo���E�Z���#s�Al2w{��~��0B�>%HL��D��j>)���C�ۉh����l�(%�*��B���������	r2wY���m��;�u*_���j���ٳ*��%������'>��