`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10000)
`protect data_block
ACwINrb0iDIGd5yq3Ozb60bdv7hM2AgAJa13fwTxCc+mYrxnUDoHltlOEL1K0p7fDtzTGWFWSFqy
/BwprXjTGOymGzB2quW1k4QIZ0pVi8ZUISJvkBjNYzSP7ln/JB/+jNaKCIf1ZEWlCuqnKj0GLMbg
MQoNhQH12gDyuVNTAFGzZl3JfCX3OPy3oEMkv1UhHDXt5zZhq/mL78YojZNQmZ0yuIA+M8Ln45zx
Hlc5ZJLeQRsihVmO9VkP25JQdrZJ2ZSaaKAaM9pvYk/ZasyNolVGRvEKXG/IB28IusHVDRDNVEk2
iToJ4Od6WQ6QI6rOsb2LMhFniqdlSulUeLqPyeG+6Ltur+xMaYmTnvPkWrlbpu4hrQbCUU45Td6b
t5BbGwNUr4Mi0MALz+hg8Py2ufyzBY43QNUHDL6dnpfSacowDaZXA2/OwpE4pEI5GABaRCj2hVPe
Jxd0aHwyMdR2urgkR6UJPMQ150zlYH14MimKWz/D96ShQOoTXjV6q/mQPoe9HqCSwRbL5UFuRPRg
xyWobhQcLmxR2+ahuk611OMbotJduudHki5FcbnXoN9UuNIbL3LwPumczkjJGgxR/cXrqH5HfsbB
m96Eed9oTlQxXBD4fMoIx+/QWPB27oYvOFYnq4T2/ItrOBUsELzjp4BiQq+8BaFVeoO835QZMuvn
5zXNs+QPMS2R+RXZoJvxwhereJvxsT5sTm4rQ1hvb58ktxz/+anj0jNex1/raADLFBQqjrsfQDkk
B5sW24JG0tTOaIoUDDorPtkBkpV4I1FUgj4rv4tH6pbuPUBytFuhec+2YCwI8M8HMqC7eMw5dgfC
Deaa9MIpQEqHn8c2aELWNX/dfl9BckBOK3BGvNOmg/0YvPafuRBC9ANEEszTzJktdBcGXie/RXDD
FkSiE7MfdjuXtcShALLpOufevnjYu6RrmYViA1gp6/7GtwSvvN3VR/3vNyxE7FSoSzK4MKwqxyjU
ud90YfuV/2HRV7Rx4xn1mSw5bMytt9QMgG4x8vy+GBe+pfo658QF5lloWChHCfMc5I2H+B6/M6dV
Xz2i8jgucr9ET9UCnWb+uX+KjbZlIU7sf1tz+571Tx6OnuglnSEBE6aLbxrcgJcgKOBXbr9C7Eau
vdWG8vi5thx60qJyOQ45siVEpIoL5b8yKw0kJZINd6IbLWDtJwqDxT5wgkf0D7kQq/hym0GM6uOB
X+2dJkHWOc/dbDqZ0J5ptDbOn0uYlhFZRmF8pFeGbUTE+Z36sHTmBBji08uJdgamgFIlCXqbwI/g
t2u0cULs18bk9pyv7kSMAY+YX6KaHkdApUyXLZmI81KSwEbSDlFROVG/92/LVw05SqH8XbF8i056
+ozu+RFiCw7ytt6AoI5netX5SiyBXGs9BlbjBqG/cvJcI6v1jphKXr+drf6YXNz6HiFfLTfSW7PT
E/b0U5O76EtKRHPV/kOU68Y3JVijYN1dhRjNjJAlj6jI6lC0QTo1f+WbDr59fuz2KO55eZyqa/iP
okfHtpGWUroKSuEyKPH9JRjxEhQgCABzckbUXPkhQ4GPToHKwyVuizdAbvtgsjmN0zU4hU/xoh76
RX2FCqiW+hHhGI1DnRQF88XeUsMmu4DwGtbjM5Q18+5NVwdiOHET8pBU7oEFv5vMueLPMzXWgRz+
eAWllAHtQIotKKTp3Yn+Yq/mRqLzLvI/cJG4NF3azH6h0Ghr3mq/b+KckzClkUDPp5f/gvLBEov1
CyPwrB4YaewttU/vNoSUi2R6PwdAWGBeqYD0JHYOp1r2ylB/f3EFhfVBfmT5T+jxXuWWguuobs32
QZtN+e24HehDRDysrGp0FNZO3VoNcXkE7JK+XCngZF5TZMKR5axaXNDDdVrGBZ3wofdptv1Wmim2
EiEPQHPilmbTZ/mHc3uJBQsrCnf8/zc3JlOd1Rv00mX+pWxqzfuIYT2yrGzif8GfYqH+2HSX6axd
jvrXoJh6cnIObnwM2aBCyvBf4ms3crCryGMf434WQoXypP4IhRP+tZmxwOwubgYURadQjH1h3L0l
VYjteGVzCVjNBjMBmd72owGUL0R97N/OO704vCHpFGgns6qryP4JByTr8R8if65ddr3r42AY/QxJ
Jt3uFHi8fLeIMe7ydNzvbmQ94sdq4A+J38sHyVM2OStP3EGf3Jv5fAXEJsONm2pV5rc7sxRJCkPR
w4wxqG4QGOLaqzbLMV8WpP+3D4cS6Ynw4bHhN0zIWtvbH5crfoUZddLxaq7aCZ5728u/4HsyvZTP
ScRpDuPFQ0Fa2HfNpLWHEWFB6PixjFKNUTsL22ZIp0QLGXCzDqdiroxWNDQxgcFQor7AYnOBSjvZ
18hPUU6bkFcML+xYOWM45gVGyoGgO9zRpfyh3qNv7ftq/qH52BI7ARQW76jQNTMfoHjmsYT3nusr
WqSJGsUlhnN3pc5FSrEtbxgFBJNAxQT6/iUjUHNtEAYya4zLbWwYf9L7rxAamGPkaD3DoIzB6UQa
8oNbBDeKtSyLRnr5UAq8GntoA7aRiAlLPczUHTj7GKNlUZK/U9P+tfAV3T7n83Dj6EeeB8iLJr5t
x1Oe3PhoHMHf1C35yw7ZgwiDktBJ9ADerpjeIOKTFDrO7bK6IIgH75rsLX5PdVKv+uEjxq++s9Cm
qrG1fWinoITZLs312dsIHk/k9fefg15c0CYpFZ6TDlPcCgu3UjZvPOR1aJhvUDdTkN1nb7C6cL8R
5REydiiGdUiPokQle3Pe5nwczn0524O4IS8DJiy+DMj45AVBZ/fXXDpHxeYPczEh3o9lDJTetCKd
wYkaH80IbGTqOcCGd57JpDKyirMLMF5iS/Ww74WlMpZV9N2Umhum2QZsGO/qjvx5cUHbA6rsxiEa
u2Y6l02os/3IXiE3eAQUSnMDHdsfNULvzE3bU+coA4JaiHzqzSs39nZ20/3/B3jaP7cSxra53Il6
CrHziLwwBRj0+elRdUJ8HsV7UgB9ROeSfojBg+pcT4JYGMPdmmc7pax7UM2E+NgEPWn/HPAtpTB6
OKo5a8DkxHcZ+iqptJnrjTc1VVBROizORDk2S1LB+KNWQSH+8aiHcWo7/u4VO4eH9o27YdpUGQ7S
wib2c/jks9CXhYKvPqtVK6xD3Bx/lWL4IUteZmhenSEKYBTn4KEt5Kycuoqt7Ute9QkOTkgbzEGG
k9jYO4nQo6xCZdf8FcD8Ttzf7cF1ray0qzzp6DM84I8b9ft71EoWj/qrsfBPjOIc709M23GHb6t5
JseeRWDoMKv2D1yRR79jGuEBQkPOiebciODmaIN56Y/qa89J8zqr54nIJ6nFVGVBGPgBfTYhC9c2
tOjtKrrsJh4/6S4zNXFBLwcsIEERxvW85giSszENGt+LjcYm2sBBp6NkJoXCqbWnENbrQQmGcSVA
L31asbyHhhR0B9XabADwLR4PLmQGyyyRfrKaOavajgCVSYU1lQNjzw5DSm5pyyqk3zpFoAQXI1AL
xs92x27uBXOiHNB/MUg0Mrxu9ySbDZ1BULYvhh8LKlR2h70HqNyq3HXU6X9of+067+QtgqUgF65C
sfLvfzYCvbggciitGOq41G5AEA/c1yqTUCL6W4hNauyhQQ79fj13kBzsYdMMOcw57NcflJuixy3N
Rv9OmmWuOQR0tDkQEoUBEo5OWBmc2WX4jQKEQpRO+aQQEsidIt5CD2NsyeteiX6WNfE7IrMQUpxm
hzOuYU52PwzbIHcGLtPeWDVYXuOSnF09pomQojov6QrXrvjSr9pBr3MLlrsPzOLjlb6HmrcDMsuq
Aoq/krpo1y1yDxazqrVlt7NftudcpQnmE5Wa7BMTh+SvepPOlqUhQyRsPAEgRHfVtUyVIT6Njctu
IHnP/BJ/r9iF/m4zU4Zvve9liYManPwZyKNWDXHSNaPi8Ke1SuRb6LlVLz2DMUPEQy1yQ789D5eN
++sz2EUS5aK2FH6eSBNWlAz83axGSBuis4QRrO5dJnpNfIsaeDWiIUU7Iyg90OcH7arGXpoHBIQc
nfagyR0B8gbz7ij6nWmvdiTKkujLVCAEAlQ/FrU9KuTqHDkEeLX46PUCvVHJURCpawEolvp4vhvE
XWA6zsdio/D6nAXgW/XHdgtK/LyRvZ5OZE6xnmzR3kLxuFdyQnq/pM0xxfwD5Y4d+g15yl/aS/Km
/qa3m1/V0Ps7jodaExhhj6FPV8TZ7hShmUm5fwO3WdaIGjHvwXJb2+BaL6m1s84QT5qTifRjhl6J
+oyhd/ci3zRJfnJFJgIeAgqTxtCMtg6yoNuoc2EJHgNi+gzvQYMAs+q8fp//jh1PfJ1U9tU7k6zV
FCl4oEsve6UnlHR8fUX8OePH5eIE7na5l6FqRyNQktt9LZ6bRcOZV2i/utS8QeAtt8MP9ecmwOEC
XhvT4C1r3UCMu9tdITQHqYZcgOeW2HO7N6MWojdmu5GGZqzqhpi9qkjk6+fSYBzbmx8jrNEt12D8
Oie44zMbbqQP0wmP/gljHHjabCr3SSVhJqrnqxyl2JQDxIjRDcwGa1p6sqWMCGF/E7xNS2p8Jhu3
/NkX4/HK/U5XEEBxqoyOrzEee1X53pDZHUEZhrcETjZpWgHWKq2vxfWUk0RHT/d7mEBYQRJV7iSk
PxvsTrHaQuvt4ixA0cYoFSbEBPdx02rEC8r4kNcnPiuOnEfe7asCRYcVcvspwLrDcBK9zU7dw78p
Phgwzd0wsdCInm9xCWp+N9osO44BIze0s8ZLH4+ODxA0M8tc1eW9YyzlDJcBSje1zDj6BJYC6z5P
JQoy5wErC64ZpQ0/Q76Fu0bmoEun/O5myaWzpLVYWb95fxi4XvKtV+9VUOZcFnVA9wrmESbVcTAw
DXjogFIW1xxwzRTBMPWViPU52VVaYpskln1alcoJ8XuaGfUeax4iVDrlQ8Tcm7OAgSSZmh3QknDU
V1vEgNxnOmTuEZwvqMtFZDaj9bc2tIHfnfGC0FM6p53iM+t0+MI8PguQSLv8nxa7EAKyJ99/V3fY
iXlXm2cqlfg8wzWviCqB3gtw9gE9kMP55TlaoYlYDs+wpk3+x4UXUkVxtWdQmBozmhSC+Tgy+F5p
dpZM/s+aC0exfOlckDpqt7R3DrV8oJOmb8JgKuOhUYI51cjUkbU1KbMXxMBWQWnuowwuWcDVNSF5
KSUpjRT3snRKSyk+bFn+8P+h6N6VWDoHjntYL7xYdOZ/GJxwEMsS39deQADY5sG6swlcc6YX2IML
yjh8frJUlcMOrRYl4ifwR639mEKFrA4q4VnSeQJCRdM+v6doh9q6um/kSegQ9jkacx7uXW9vOBmV
0plJvhvsU3ToYse1kDjjlD2HbxNpOQ+7tv6daN+fBo3eYablU9/Hju+S/8+d1/arS1rHCMYHlI7o
yukOhhmtPzdCZXTo0GrAPoYzFcOFCukuQMlpsokMlUZfPupTN12y9eB22ZmIf9+CfAmmsAcArj5a
RL7MG8rZugImwB82a/M1ulBe7JXxooZh4WgeviN2FCFjl9hqyumd9rjLQxng3VSQ890z2hk17CnA
PqxoPK3dZ5694KZ6D62hCXbtwopPorY7Dr//Xlt9ffllfXiDNRp+5J2YIi3X5PfObm3LdroPhK1v
j8pLWqDzZHMnAqmxH2cpRyilTFhKwahwEKXLwT9SdjHDi38b+QfDUfoeni2tf002OMV6VgyDNM4t
aThWsrPlte+4+5CI2PkmRAsSZukHqJPC+pCwjmRpL/BG/h28dg4oePfO2MtSQi/s3epa1CH4sNWD
I0kvauy85gU9ZVVoVfsFMk500X0Ahj5uX5a/S5LyN42Ld4O9n/RUzoqDHLCs5laycpGnhkJ6p749
8zLZ2q2Q6h6ejdxVQXW5jQyP3CVm9bTQg7Ooyhr0kHYqymkoVrKVHeqzr390VIcwGi/aqVZiMJ4C
9wQvWRSCfSmKeNXsPhOIA8Tblpja2SryMCFoVtnQVP4rai4z49Gr8QUJGHnKljyl9naaz+fW3oWB
duGY1Iznr9IR6OulHKbQkrP4OZ6qG5qp8BMbx1wlSY7qZ3YYF20bnwTxIsCGm4zNCpx2NrqptiOf
0zeu0QM3NQZg9tWuXA2xSpe3Cax5FlPEfBYDaPfFXR6Lq3iNJIRKoYo0NKCjRi+fZ6/U4JBAGXcp
IXVfs+/flLbaj67XubVB4fpqCSTGLWmL3TERExDV33lhDU2cF2cE5ZmJRBCwwQhtCu6Ub6OgNrx+
56VaLFBEFU5mqvIEs6+tYpEURlAruz+bdx5wYGLEWXlNmusacZxGKTbc1LoLkE7EhN2asiBlOwTu
bNmVSiuJFTNtEtRZ2kSLfPLa2OJUZDimazQ7vFPEv24e11zFTUj3qIYWRKbekHWi+ORa84amz7M1
mcIVu5SlnZ2QmxMKdYUWeghm/+yD1OEgltzAgzNDSngE/6h9IIUIBcDTx9WsCFhxxlkx9QVQzaQC
GfdfBYPdKrdJJNQRvZEhEBV2xlEJtZYi1sBPKWnhRGSD9VZMOuWhfw6gcpfUEX2+B24TvBPUQxbB
f+GRo0gJa/erysSBzfVK37wzDKg5HV9vzX0BZrR+cBm8L1sMLdlr8Mb8NRbrMGia3cLmldSmuPB4
JIAEj6LPUou/3ZOr+ZOou/gSj6KrkRx94Uog9WrKoLvUhdq06n596FQ8PU/GmUcRQ6kfflmYXtNF
kDasMOOKDb6cAMWohX8ufAXdCpSXqRSQWCPFeGnkHPKLncwhvk7N844Eb3/RIpn/ensYtGmn4NAE
kFCYFp74GvE6ZJlB0ccmv8A/5i2+hEaNlEWiYyedGdLP7qJAjMib670FG59DFqKHHfM5AAoXHa63
+H4F0N/XjL07xZb0UkRX4NzcrFlCHO0ZClErU5iriqZBgTxrOCAAthGIpjsRxeSH8nwBoPNtIPwO
VdzMoZdZ9+dLpKAj2OVNseYxxjAEpkyFOzbbZCOSUdGAzRcnXPTbQxji+vH4IYposhxD3OyRZa+i
JwLYO/4jrUq54K/7Zdh5cFTgIBoKmaTKqJxDOwEjBtytqGDigjtYBTUfWDdZNcbheQE5bSR6Ulp3
i6O8Z5ZbHsRq4iwyDvk8H6H6amsEhE4D4xoy08IHvOzjw+xrVtjFVMGDp6dTGfunROCYx4cD/Pz9
+lXcAzAsUI2Vxr8r5RAU3D5Db4btRrxWYyhJ6lIl0U0AarMwZKMqfNx9tc51bWrXsshme01GlIsl
NGc2+XIqtgFP5og/Vc34ZJh+39yyHEiru9Rpd1joZ3XHeZEebucvnxWmLxW4GEL53pSn0mSJx2DL
S9bcZ0iXMngJe2l1fTnV1zi5Gt0GETrBOGs5ZKLH8cEEvEJU9jm0VOHn02TQoXB+/GAWVERiJB4/
CFYkqNqNP+Rh331QbIAPHWunc2F8M91x+Qgw+fhHm9qglAG2eQgGSJ4+KXf1o3Af/yTa4/TdzUIx
XU3q+bPC/7n2IcL5/ytgUOx9Qc1R35b7p/A7f29V92fw1kA+gxu/C6zo5njf0oAwK9sEFjl32+Jh
URuiC0ctCZineVtNs+HuC0pqbMur3EbOgCyKhcALBp3uMD/CM3W8jg0BsY3NMHwYIQPHp2yRIdwS
zGhf11yAbUW1vjLj1gzRB7xaa9t6gzdRaxoUvP2HD4yuaxR5CTcmgsxNAg8FgRUDgtUS86THzcBz
pXYxLvtVeLfnMOTap9VaoyzF3yJoj9XHPA5XdHyw69EMGjqldIINA9UChLO1F/nl1HVHP0vrv1Tb
DHkyYsO05dSzP1wzf3tCYD5B4NxIFWqMxDcOf8OPMoFOIypChcQtlQPbHcN9jbmGKgRyyBoWrLQG
cjfSwFHQ2ps8XMMEXevDRDp5J5/H6bHjbtDWL6vno50+LKYpXoPzibMoFUtQv5lBbj4fd0DNvWyH
spFEhxiYTsjHtf+pPV9u8kZ7LWgAWgq/AGDdxhdiWJmING5Rm4aMc/JdJOOywYFVZSOnrABb0dQJ
zdQ2dTUr5Lbn8p9ncPRIrzFScPayDYD8smwJ6igRyw+rW1Ou8X85DtWjP5sxvg9j4uwaHsXNBY5/
bVuLQ/wqP+xcyP6dbvWC12sNjPgFyjkypbSV6M3osm2IJX7bFfpYj1b3GzY7aZkVMnm0sEKXzGaO
M+2og7nICbPadOaaGAxuhuWWonMX2px9j2jXZj/eeddIXVDDqoawlVcRol+IRvGN1R1v7HG2b5Ce
6Q2E++6aVCkzd/FWfqP4d2irHTuvh+PtGDm4W5jmSvHiYyGPxTa6QqodUJKU0zDjhpdpa7FQc42V
1iBg70YhNM3lQk8p0K5kaG7vdWhYLB5skiFCPvaqNuajVfwhRAeDORTATZc7qsnx5Xax5PXXGCWU
fYb3lnhcazS6z7tztYCP8FQ+uqyfUSbmcMJznvwsAjfShcJz+SIe2XYjcXPUbiBMKMcG7Lp0lbxQ
a1yUkFiaA+TAIrYZ6GKMv8YCamd4u+aZ0Nyko6a1w2gUw1E371gUqWwIJ/sNgeSJ9B4SlDudzc7H
DI1CGut1cGNXfNNQqdcRZTzKuryqpLLCRcGmMHbOUxA2EsxMfBl2Ot50toon5J9RktCNt3WWct6l
69eA0EzjryYRp+u/+87+CtD0624bCqIce6EhJFIZyo30wC/Uid8RcXoYPnHFI/WNT0+lPq6dShLn
N8bTxkGr1g8pqRsBTjuxlxKEMFUdO4txpWp2y4wcRQTeZyBDfOLifUl+UpjXuVzGeUFNy0RTSNgM
DH2F7y3C+ARuuETne1pV/oT5Msze/C4mdBtdvYwxbSjq7Xn5CMImOjfN0w+/6hgD2VvQ4wTxDwBn
2toSGEVZVLLgTXQ+Jtz4GgCC8V7IYI6mZ7WuTWBD9ibP/WhFRBo4mEIURM/rbnw85xT7jgq9ykeF
mY06Ss+qCCiNp2rIM39A4QdI+pKhA8GsQQGNdmxe7QMBwCq0GjeflKawzzHaB98BToNVoyxpy/Ib
m7l/FSiCB0DtkvO4Hya4kBk35x3GDA8p2eakQqnq8T2ii4EWwgTKf2ze7nmH/xq4jeqBLON09mTR
0HHFOlEoo9O67hTEd1ZXhJ1TULmiuw8TlL5/zf+GCxVjYKDDEGsZphVULcPiKgUFQGVRaqOKv8sZ
DS7ulVxg73dYQKw2oghdiFqzZGzxSIDa181N/2QLujysaeamclgk5BJV6Gm13wfgnkvHsaXnNIjM
IEMnteeeueAfV51xKxiYr5zLxBAuCvaxvgvTrnUWimbef+KqqQPwjfraqZV3CqbMyFZV3a8f8E3z
15T1JiL61JbiNJF3o9tcTej/ZMX7bRym5dZtFUxU9NI0Zsf94VCJ78olNV471Nm/jbq/DApZsjBN
D+pZ8wDuUO5+TiyPjcw9Gt/NHCLCI6I7MelIPFpdU52la3nzWxXsZFGQtOhMCEEPbSpfTwsMvWjL
v27hXYWzDQqkxoOUdCwnu3abdes7Sq0tJy0e5x0RTZaU63ttSNWx/TtTOomHYxES0IQeQvDw1NFR
qBchmaUOpHws5+Kt5sm3x/eXCHHeFjHboUIIJaRtbvlsO9z9VKbcvl8khH/nPSHLVRqZ4HJcNBr8
HO8xmpo/7NidB20X7WWaj2/OZ0ZovRa5dhHQQbRt0M9fL4oUJ36JZLqPefUDL1oOilFNkdb69vU9
JDk4SW8rFLr2MHW/d/SgMWZb6LfI+njiJcEFILsEAseMgkpX1YJDjSU1u8PeO5qrmo6GwkC5ZY4b
bwC1zGMOHYKP/xluFFY1ta3JxMrk5sCfT/JAXx7gwm1o+837CQOOxVJuUDb7vQ5Od9tgTcHaaoWr
icvIwtppPR2ZattnJAt/SYb084uHJuA+y/re1frvjAq+vWl7Ei8DyRjzJ8zytfvJqyGu8BdQZDDH
UuWcOOBDFYW1MrQzz0fct4VkwVs8y3E0uVMW3deNFkwlOw/mN0fwHAxqfE/wB7xJODCy85O807mi
VVfxTLKOIOBZ2lMxMUFf9zRxWnuOvoNNhBk03lVtKeqWyDan5ABWaBRqqyXAmkDzDPVisqE7MJrr
HEAP111FwIhzwUvng4Wa4sld/nyOuTEtcSRypxPLtwVb2rwUdHpZjoPRT45cK1xQVw39umaWKov/
bpXnBhL0WegYwpjToiMvUxTpdFGFg8xYJ06k+6owXnwE5SNXWY3ilvhSrXDjC51lafPrqDUKXYEv
LN+UcR2b6N3FoesDt6jyF+HFcVjI9D+WN8OT11KRF97dop0eXjIwjAkRPsQaiyYMkX7k/TEOy8I0
iFpT9GbsB5P8UcplFte7WnD8WIxV8Nb5QR1QE1h1JWM8/AE/o5emcYIWMBA4oV63tMjTrsLgJMMH
birYlRkqFaDknyoIz9u6k6Zz++04EB97WxkhMTrsVQ8nYEulzq25tFIzO5nB0fu5aKgGVuSueUJU
4qgyPRaKOyrE3iQDq+W5fvRkXv/EglTUnmlYUipyMQOEoOGV5xABiP4Hqc/W8R+9FQGBR00va2B1
Ppw98rUSe3o8MnlIqah0srI7/9m+/A3898VVX8USo2uATU2vgn3AQeoXdFG+4YAFD4HeASzg3J29
fdJJipRq60BEyL7R72WLXttpF57ywAiJ66BLMS2Q2VOo8x1af6o0xx3PI85z1xrLt91nL8cZO9O8
m6dTOf4PwGlq1MZyXHjx7mfeO7+A9Rxt2ABG7d10usrlAYi1LazxjWGDb6whkq7VbSNVcEY6B5ve
NGxMtSb9BofEFEOVYox2wiOuyo//jSJCJSyT7kxqtlEOQD6ve3agsfaouaPvBJgONTQrjKPaxfoS
2gwYuZBbXVoyRX/mTtXW8+KsU/sYse9sWFjwuDEJCO/DeSJmLz6W5N5vxCjalO1nM/n3v922UGC+
D9L6gsty28X2I/jwPjuW0GABosf3bsnmv1skn97XYnfMO1UObp+uIJOST2pZ1ewUHIog3xWtCqIX
8AjzFlXck+ExUpgs2eoZj3jUCFPmCC3k78tHxf5cHxOGWahZfQN5/nzC7RTUxWo/eGv9LVj/5vOv
RmHpu06doIObi4VyhuiWx+74IRDsWZr3pgUL2+K24AnbKHhuo2da/1Ey29llng0Fjg4H2XHcyyUV
16xymPEAIlXKqX0lENWl/etuvECt0Go9EL+/UVdEuHVA5er9flOWu/yiBRwtcvnFLQeqQgvYZ1o8
TuZecLpqMR7aBgxsPklblmmmG9yfmO7zoK16n667Oxw6Q6UbEKXsHTuFvv2gk/IYZVHfbGTuAhBp
hDeQY4NiHmlo1DSRYkPlqny/NZWJBdCxZ2B75w8NKDkAAln1DldopkafY4iTuUw/8K9KD54xpynn
P/R7E2+BKldIkyXm6VlL3YmbpfKO91el84wX0DJf2wTG1BhlLFyqLwhZl+/MNP2qnmH3EqjI1EGr
sMevLsLGLo6HSFQektEFFyCNK6+ey4/kHOwZiQBv2R4LK3zsMGqj0VyEi59JKg/89KU6HAKRnEut
Wo0TZO+J8GIJr3zJEbkc4mSxOsfiWL1s3sNqsC5ny/CQtyggQEnOYSCIyTLVCy84N1AaVD2LW/9/
9AtIlBnBkHjAwETB6ml5yb1BiDsKvHtlKP0lCWiG7DSgdY0Vjlrcc3LG7Ogy6ihdqKSniquio9JX
iiHtiMBr9S1mZMSjpbSS92VYtTr40gDaDLZYrWKfRfarjv2aosrtGr0yzHHDqqDX7uOgMEY0J9Kw
wXon9hkQSU1dNg7bU/j0HUgaazA4H/GTil0X7k/9AqSVTvFwYfdx2F96OSeBp5oLf88okuAjIrTV
E69jZ5OECS1vjxZdRTQW1hS+PLqYSOBJjdkviFG+/qkBYFXoBZhUhPoDNdaiCO0S8rK/QCeFUijq
En1cRTJFIde10YzXozjfmIcrFt3QE0ft8VO72qOHbbL9Rhlw8PGb6D2LkE951xisbsmvBjdHTSav
WV3EjQoN4HoMfg5diDuyEHjye0Lgum1TYCXLhcrb4UcJzOX7YHrBdoOKafJ+tWs6RtL84T+GSABZ
TKrJLbfnt/ru21qzDrj4t1KtWD/OX2rWzBQmBp3vIc8f9+dUVuiATpMW8ineHGYJ++2PKp+sosbw
AU4/2JN52KItMo1WN+cMrXOQ/MCnLHNYZ9+UHhi6cOd4ZDAgiK6OGe3W0jcEbNBh8UJ3lkkOQ5jk
5oM7byo32xYQykdRvrP4R/5LBSIUwe/d54gwLpUECtPdOma0iqrTsyA+U3a4O28IVi0CNqkh9J2W
pvbNfB5yrJm5Kw7fKCGTE2APjmnSDxzBXHk8DH3wbRDAvy2nRmSE83JKCZAdZDHmMe1tNh+Dda3O
+npQEc2uW0RkNB/dUEhW13BTspb5F8P7pHH8piXnySpHwNhgfZTRWdtDHJPNpRmXCBBIJUaKiUpg
qJuFqbbz/GxjQc13HXLgwY3y0GvEzsWHT6BfQJ0D5pw/ukB4Li7WxZ+jHlIwNeUe0qgYpflnX0+J
sQgLJuqX/Nv3kxdfhpTQ8nKWGeDI/wGHLHcvSOW484WX7JDKKWocKzyPCaiFZbKxVNG4QUTA5A0D
GyWPBa3FkoTxwwoslkF90cGy8XO9dvm0mKt3tbsg9kpMtxss7tZH7/Lf0Hc0S3ISO3TiOEUeBwUx
18klrk3pzOrFNHyuuiABWhs3ivvAzNnORHQaM66YYdxNFiT53Uy/vi7f1mFdxO5px+NXE2q2uux8
szpVS7fsS2R5Peuu4RoDq8XJoSvj5xKO/ucmfaoTQgH+wR/sfNyZht2XqTypKFmc1JvYjWU2T0vU
aDiFYxworXsatob5LGlApbBg8vBWiRBpfR5vSeaVDbQ8j9Jrp5VtozE8uGXp8FQbJ7fclk6ndRhn
Fojhr6Zjofp7OIAx0tBRFCQaPfoOerFOKWH3L1o6AL/xEig93K22aF2iScYexB0nGjo4C35qIfF6
0vJWn8XeVtOto7hQfruPOnuNj3sq71TyaBds26RKzA4TjqXzSsPtdUxGZfSzqnuTXcvCY84Ec9Gz
wyeysYTqbjSRhxtV+TDOc+lh0FJODek38FNTJEEwuc0KXVM1Ut2CacRKXzUHH7EAyltSje8fisWh
WwUSKq8xAWsmK4eBsqSETmRNUn7IUQFVzdVS9gwHMWdpxwmH52b1xwwfiBJxN1/ZtvsQdmeUdYCX
fP1oeODa70Rdg4HAuY2yLWoCwwrSAcqnLwGQn5xfSxfw3ZPyGsmGuOB70s4/YNDkVmXf/2OS9WFR
URrSKBlgJ3kJ09F9EDpSOL42TjTk+GUPP8oi+1jELQn+YuXuk0bK5dmDW9Z7lvWP44yocFWpHgU8
cR9jSEmZAloIDbHmKhUJ7anqX4l0G1mDHg==
`protect end_protected
