`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
m/tQ8xq0KytPPRUVRbARB76iNY00GyopRSgZsh13QG05qVNkkygNorJ5nRnGw71hTIsX3+X2WSnR
vkPlMeWvCXE1I1YPvWv/ZZXkyqEAWmt71x8N5s8bmgI0GULGbFNqo7GT1p2c7I6jXekuxZiC4L21
GoF5ALwlqD3KDKXwZi/NF0MshUp+XL/kjM2llI9u80Ajwi3spqHaLoB2IfquF9ioqRNtb+oJGrbN
iQISzFvtgNl/la3LAoGivF8YFwgMpfVejztxU6yLEAKk95ItcZH8VOeGTkiQeYxQqBhoehdqXYD4
SkUQh49juW4nC52roLGgPpKMMBMfUSg5Q9iaew==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="HilQGzW0u8neqGzdgKMZ8S8GBWSGOkZh2OnqARsc0nY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18688)
`protect data_block
fzhguWZh779ehtmomoELVRcL93eu9hcIvwaghrY75t1+qgxRhLD0FqzxfDPTf3t6fzf8wfADJ+mh
h4uD32zKWb40kG4BtGEsdDYzg0Fp7GKrNKpoTBcQ5WlbkstCJgthwJNvEUwTQOvoQOcUkkTX+mM+
WWbpKOCt1DnmAhdMm1iGNjjM0F+/dFaPyWVllnYafSuJwoCO/6TMaMIBgoWtxtEmJOr+8jE3WMHT
x1v4cuRXIcSucAtpxd5YoyZqlpUlcIq8IKUG7+EPZNXpp97wq2b6Iu8NTjUjLIx6S+iQOfdj6jrE
44PIicZS38gW67vOBLmqM8zWWOXG2IOLEzZx7281qHgDjEvjlgDkKAyqSbJZpI/Dm74cx6rGDQaE
p8zjf4yV4Nqf3a+7vIZh92UZ+mQmQAIh22SnaMiJuLEmD8jPBX+V01bkTidZTTcyPqv40OeGzzh7
/F+txNYAAGTWofgBF0nOzF0g+maGTbMxlUSHzmvT30SL0Ktvz0jEAVlUNA0B96yQTRO2Ku9Kgn8+
hD46xV8OBIOdwUGnAxKUZuKmmd5V6iOUiMy63/xYD6okjzXqRqfkL9tgW/hxoNoBaD4Z+B5glt2a
3vOSQ+IWevDJKKQKBOh8d91p0ZZBGJTXuWNEIHeoJlRlWWjK1NtxKX6IeM6XybIY1F+4bwZfM+3H
BqcEbpOJUJburShsDP4IveylYJBn0lAXCtdZARyhsOML9TcbIDlmkVIkx+KexTMqAfTKzxaS8eHr
qEFvbhY81b1kl9fmcuvFYjsMrlFHEl5w0DEEVCaG6G2ed8nyPnmob5QJ7SkvpzIlSmAGv6OtZlzC
oKFCy17Y95YzoUzCszN+tRhP6vHvkGJlFPugmo2J3INg9jembHVgTd8Wi2Bv8Tgzb+c0OVIHdKgh
JcFP1wsDGTzwp0zFReblvgdlwGK3EAZVHjKY/gwCC6FPcymcxc9GF+E6LBA/dkdAhEDHxQHZ/Bt4
bD2fKXCqJKO9XMMeO7Jwhu6VgQ+oYEx3qxNN0Mjz1KYfpc5zQftgk6uMhinhmQeuDoCmJJ1XvB6a
IuMTSJCLmhBg7EPvyQcEIS6nWnkGPEZ15YahbOQhmhTcDMjwG4/md3RFilNAkoYD0DB18mdKZsf3
Js9XWNu+3yo9SC+/u2RcPWQN5cqbluOuc/mHMrAoNp3c9SyF89xV41Aydt0NRduy8p/PLbxeI1p6
Dtx5VyHFrcDIH5ocZQtJ/8NCEeaWgjXaJm77GZXeMXN1LmCB7jJg17xv6Jfm4hUZJzwOPsT2MexK
4On8DfI+G9RU/HzjbJ+qfQVzffCuuRMtODTYKvNhK97erAqx/7BfA0KdiDuGBS3uj/3Qq1VsY+mK
uiRqj7ya/rPJRdHrkBZeYLBnWBpbvbqiTvP0YFCmx3f5qbNuuBBb4pBLQS79ecMEBdKC8tq5lxmG
iYY4DgCsNyMd3poaNvzLYxNQp8GfP8I23NKRrgOsNuIyP8GiCIXZ/EcGg80KyhOiLjAY2dPRqGYF
2Jl16X4F4rbHz67+4BR66mAK8ZruA0OlWJXvCA41VaxGFkwc0QuLZsBBsENjOT68B1iPspbPpbgB
8Mcn2w6gpLFnBjMXLDdK/e4AClLjb+2GwWIjruoBv/qvkEbfiuJLxDYyO2CFOjhOJMLyUu2RxiTO
icZXWocsKR1uZCIiY1a6dP2HRWqs0wRgOQshh6V0ZoALrmmbMqJh9qERmcd/PV7teNBIpyXur5Ih
knk3N1uHj9ZfXqPA9SJLAiA4bY1ybRqI/1EUPd7bHNJeh0BPgMhf+y85c6rVqG8rYRKf8fG6ZHpO
/7jygGn2rPzwdTvL15kLIbfhN/5a0irPTO8VBz1mZsVJwNE6bDfxVymcJV+AjdnM3Lv4/doWKsrC
n230A9Xj99u0b18dvRdepgM4kRBsAqbwlVxTjIkOGUFJVwV0nbapecMATDpRPYaTO9lL0KfEwZzn
uKwcJX/fhamB+eP/Qk43sHu9AGMo0UDKA7e4NllDlWFB1k8v10qzmWiOFmPwT2mtzFmCPKbmk1Ty
vhDDUd6O9MXHG+V4PFcr1+aWn9whncXRmzm+vL/kaDL11KC44RpVZYkhYQgArXejUUKvWedjHMIk
qHxc+jOdeVWub121XL8mtPQnxWC24JShVpnJxUDpO6SA3SIVg/D9ogljl82OgNyOgKA9kedwm0V5
7IAjsPTExI3gh3uKlADyQuKX6gEqCoIDo7FDNmlyxfJLQ8lUREsp/Hviln1Lz01oIWibEe/sfpC1
3I4YrEpeZlhVTJlee0btLja5BtSgVwyKsPN9Q8kv7IkH8vO/bJFPjHGr7n+AJ1DiO6dTHTr2qJd3
6OV3YvvWGPSkeIDxeHO9aD79RogLrSbgzjkw6AmRRUbt7hxcMdvd1iecK7v2e1hllLNA7WZ1Ex0X
auWWdNAUA61cyaDF2Oe+3T5KyKSPpu2eFzOzovaxL5Ae1oL3rncDYSXvGZU48bH+mKUtdYGIi96T
shuPZXo86drOuSUnCSRtFtRJijeJDoCeUVVQp/Pm/QbXPwPWMTq+lYCIJyrOKPjycDtyaRITU5ac
eBPuG7e4dsgIS/HZtgqCFb0JWMK559IEeG1+u6WGrWl+cDYmrAR0xiSC32TQD377wt7dE1mNsX9N
xG76/msMYvQ5i1I/uhI+uHsNnuAhbCbApfWlLoOYdr1gDa+tQZUDSvEUgaEkj/lbQWdPXAU5cuNS
YYfZ8ntJQFzlN61P+4wZTX/ranjfZI9DqMcih41KyuVoZ4GpQmCBZN3R1YpCeLAjGSoQUpL0Szgq
XPpPL48hOmjGQsL2xQ0vLlYqG0dWKlxTKxUpyVVflww2PNztcgjhA07pmHewWznXob2x+0yztnmI
Z5RPttXFtTuec5aldDxrLFTLf98hqZygDjxN+YMLV0qp1KLE39uI+4okZmpj9oL8PLI/KSrQ5gHk
RA+LegGP/xRx7/jsZ+2Zb/J7RNrv58AWkz6StAzmz1XmM9s4RHPekd06SJadW0vuB9KTGLhauW/q
FoieHe3BF3Gm+niC+DVxhAW6r+h9bo/vCkX2HeWeXFC0HjPVXBi5lQTrAnOCzGqzQYDwmL7lYL9M
IQCntRZEamLedrnB1oTh56G18QvHuhmy8WsPfl8e7gzrzTkwB2OOUp5+O4/nqalBQuCx2v6WpRT6
gaQ/ySVfx9td5thjhpeF1+yX8WfmsIIx1jIOvKsHUaELIG6pmNHYI+4irk1IFzqplfmJ7mg6PJoa
gwYoZFnJpWPFdcyElaRb4UQfwuM6tfiHwn2jjsnGx3AYNpoP8v24oJn1bnjizgb6CSNTTZz/zaZb
lOINQAQfbi/vDNKQ34k6UdDfTkZkzK0mCNYo7XNMTCmOPY4jatbbs2sSxEdNBI/XQM1+iIxubhzv
mHH2HmhCWdnOTTWB3tPe/Qkx8TNLmRsKv3MtbuL1+YSribRXwUeBEy4hnyZ966iUt8xKk5LM0PjV
TCgiB1peA0xSB5u3GdjC1309EAOgzRboWUVEZZiKniZebT4NW/ieNbtWxbIJC+TVRkm9npBULuny
gTv9E8ReGjNKL7CHgK71662sRVXweulkbMs5SVP/oAwyEwiR4gHVUUpepWaBGp+U/eNlq37nuDro
Y6VmsBrD4DzmT+uvOQdSfOB5t+feQ3lkCVcXPj4upuXa9XXN3Myilso/Bq/6hw0G2FHBHNK5wVSt
ionoHEcCmnZCrrrxo6v7sWlC4KmrKocB4eXxHYe9gMxIeyChGnVH0QmmxESdOXjRjKAJ2IFPykcp
TlCyQ8DnSLkdxonvWj2gqjp2RTB9SPZxBmm1CDKbDCh3CjXzYY8uqgNIvuVpB/axFcsputHLQkFC
AQiluDeEI8/bSS7zDbatimz8U4CcoodtNLZxHTk9uFKvNawq09oLsIwXdf/9EW7P3T03/X+YfH3T
HZO6y4v4EpOV3hlxmeKxV8Si+tE/eK9sqmjC6gQEnwerMYKQh4AZkJPl1uDBKxG8/9kb4o4aEoPN
LD8iSSwm9Zxx9VEQZR1CyiYHjT1VBU4jK0kdXDQsYpDokGURDkYLHx0ETYkY+5Urhj9krY0arhWM
oyYYwmK523+zrae0E+J7aKnaaPRVD5c8C3KyB3EiQmSQQ6Kwr3isazIJk2h6+WW6JnHQ8OQJXLYd
AEaxN3qsQfgPVD/JLCcU6FGZWaDv/bMne3zV6zXeyi5ICuRSD4MCXk4WqNdQMp5tktHD/9FVPc1E
2E4Y316kHDRvoM2SeabWKDFEnu5Ua9wxXntvzoPNJFGMRbhqoVgsIw4kDoMPa0wKtoj7tmTBhIrY
0Hk7A2OnHpcIO0T70+YuZonM41ubZkkn3ghJa+jV2A8wqqLX3m58/DWhEW3g/yUyzibKNV0y5Hkv
ZUDw1JSxVM7HYmBN0LI+MgkQBRbbcSme7wemrcCSE0Wurgl+I046hOW/VxwNQK9mDWVmDsXYiqfC
vtOoCTLABbHlegzO0FvZsZMUsnnNtYo2YkNQgHAt1NYfB2e+hZVk+mqvsHQPDZDA9L9ZM2WEhcfg
iyrtDpZRPPS3ovdEJFJuhlA6tv+ObJ3L5ejRnpApVKDrUlCjwLZRxBOh2LU4wvV1AsrCT5gVzvSK
TnhnpQedhVCTIxZssiDyN/jdSIXR1el9ViPPQ1ykA66UZvR6etnLwdIhJi+RB0B/gUEG+nhjmg3Y
2H6/1CSBJkQf2xb3D3e4SUARHP1KhPzWVaI8aGaeJjF8Jer9ErJcYb7rdT/u7qvmHMJ4Cd5FqwyK
G3AsOYMGQBV2I4vnj/ceO+mqnIguc4UDuHg+C7hnyx4ieY2pzjVegL7eD5ag/2VDf0DyDrGsWbM6
7ERUs/70V6cbWMJ967DWri8+E31QyjcCQRNMgsZ3L4KiYM+DnF65tZ0mS+zQrUSXjgxYAg+fLJxi
DeZI+tMtfK/BGxEy6jntIahJdlYpxJeFq2h7AG6NvE1HSZQOoCad3j8DaEVVXz01YjPwAQG00sGz
WVrZjOGv1adIzQmPXiaPjMkRoufQO/VONE0lnPF0uBpLw/Cmoe1AsOM3q3rFBZ2TEaMLI/RytNCO
sspJqH++Hg+4+jnnIfT6vq8c0L3BXnxRlwXEX7gOWIMcm8tf6QcKBJP6r90ZT2H8VkJ5w5l7wwp1
gRh23jvomlWHGmhyjNRgVqp23G5s07jUt3wn+M2TqwzCJ4lNVC5qFmdTSzw01HABMqxIYOFH/b9W
xB4Ymv289FAKsQsCyDQe80c3wMs9f261cS/Z9fdJZOweSdq8syYgVf4QkogIFzLXYmQ5c0VMFSF8
4kTdHygU6+9MkQ1qDcBwwxbAfcTeVWKabdQ/JnSEXsNb5X9tqpgl5TPa4A9s3FLDiQnaU1cnbsDl
Vg8Xxz6XIUsbWyhfM6EwQUrhh6TcPs2IH0dXur7745S7tmMoz9iurepv2tMoUB2hYT6Dh1t0EfVq
GX4cQzwLT8TuCcl0tnsf9PO6AjxwNFsJscNrOfhVLvPUJY1fatq6fcPR28v0wgeWqJrI9xig1SFO
7CTDDNgjExB3bX2QFJNerEKF8nMgKZqVtnjq2uIer0TpchloNZ8L8cT1DNV2st1YotiBNfidT8Ow
J5EzwTlcuiZrSGdLjwl8joYzwS653+LrUnvUJaoaliVZPkXyT7u3GfPIKO/fDKoHST/QKtOznR7F
0P9Hzn9VDsy+xdbiO9B/6uFvR0Bw6I3jn4tpbkduDcpusP5HulwUOvKdRrPtxRq1McEgdxMYmkJP
S6/pJOYiO3ODikVrnvMMxIyhejeFxrNExE0OF9yt/8z80aMmBt7/MfUjX0VuLYh7xDOXOQyuTP1I
B3nUUv8dP8RUDxwjsxK6uxnaMiEx6+LwW8OT4p9FMUSUVXdSqarCjKUy1lcQz5k7A7sFU5z4+Hrw
K0IVkb0JAeX5Nlswi2okOvpW3RDIWON8QFN9hhZsIgbwty31S7TPA6VDAa+xKArWMEJz/ToCB5+h
7Ir4i23ebwCHw+5SQxPD8sRAM0RtnRKVYAo/YtckZtBnnb8WMe64UOHh+t9ju9LIGXqBar/oVni+
1SeSKyDTVV4hO4NiWppW6MaTvYpW3q4g1ym9cL5DliLtfNnwE83T8sTLYBnlcRS0wyhbmJOv6yDL
uAeAcokg47CJ+akG3LNIe9ekQ+IcKQV8TU27q8s3TwH5/U3YMkZYyuUDP9MdsnaCbL9/IAYC0Pry
zcNCHs3i4c/g0yg6dlXxNtIL8Up52dQVWFbtkAgU+Dc0oPldHh5Ec7wvMLn71ZJQ/zH3Ml4lawNe
Bobhz+4dAMTqcM9ubLOkTPokdHU3oeSMeQ3lwTs+5l1rKxmpdMPvRncCGnT0nPprJJrfQrG435uM
gagnjZoUKELmCEldlcu1wfzb7MaPQ6BXlfofQTFxwtuxYcpYsv44i9i0mLfZeqZvA+TufcX3ZY8n
rBdS7X1KMMOv1bB0xUgNDz7hp2AJMYvDlmKJVpPVFIPRCuVj93z8UtTHY+4tL41NlEYvkyLqdlmk
L9s9+PFfzkBPvdeFu1MYa2u9JkhKY6x+qpdA370GkItatwXWijtO+FSoq2dY5/S5FeXtasc/EwEY
wCi7zONUsMsPt81eqcSzDEHuNQLFQUW1WmkJ9ev6stelEbS7BbqiyFgjJW3DcqGeEexXsao/AdGZ
Ny7oHI3C1HuxCHR5eaZO/eNknbqVCW1bjnLf5u7Wbb+HRTE2bu1x23fsgvqMoTU6C/I5tdl+KE0O
JzGTyn13oKptk1Qi3U5ouZ9NKxOtgEIMJUybNHNa/XhJYGJOn2Jubp3KHWfyKmzEjDTNxBP7596F
NPqIT4OYn4CxbiM/5WRpd75eHPbeadUSxyDSS/9htZeEU41jAegK6gg+TQe1SwY0QOfzxboAogqs
JvDYPxNTgInl5GFkFgf8WGbpo5qZbzqOQVAVJBrd6V22WQIEn7MGWF2J/vHgouFkWIfT3jjDx9Xu
BPERRmYqImU1H5Hm4zt8yFPCZChfyO1ymTdaOvmGu6WUPEkUasYz9KU2HpKRRsI8g0sq03QMqpfK
Z2uivgM+kSq7Bqq5ILn4XgPkCUWc9gkDADtrr1spl1BPyM09SsXMPpOGv+flm4yOt/CTBWIrEvB0
Ul1ADmmlWEBWgru4LWhaFbj2ShELQ8/hkczmirV/Y3Rhm0leMtkl+uq7whg+c84YWlH/pvKct6//
0VwyD1ub7WgpY1/nJ1bnwyabOKPMr+vKXb09xXL311HLnXR6aV4PaZ8+i4cVM6SbMOmGf4X5vNHP
tjSMUO5AlqZy8d/MQ8Oiv71Sc9xTbzweCmRfS5QCuSahnLdmLHIIPKA68+53aeJS6jCkcA9riRa5
aM/s7nNgye3Z3WshKaymOBqBQ5Hu8K1tJ8NWg9s7xOApJNk9cJEB/Ma/ZAhBd/Vw7/oj6iSQFzPd
xRz0OvV/WQfirh/8zXPmHLXNC5b3dPknz1FNaA3RVGlwJqZsWfWy3Lk9SnO6Mho1PpDNtLdoJLfD
NKSLOSDWUs+oc62PGID6nKba2eoxvj9d+82ZeU5PeYQw/+9+KEH2tQS8nuuJBXlS2lgGRWD4CDfC
DxPek0YH9u2r5InPA1WSHcerCSCXD0Hd590QRIBv+qbBPmzEfZXv9JZv5ppqDTJOmbPnbNo3z3Hm
y8sEpBKdSYGr/js+FPTigpuDf5eR99QrvlSdpGnPVAw98kEFzyyC7tY4ft7QDY64aMZcGGmEGOv9
tOGFRonMNIU2ql8sL3YRSBabYKRF/GKq40xjvtcxkOEqU3VxtRyxsL5ZqE1mB9M6ioN5NCRPkXRU
tpJNZz62zDln/a5Ab4IL2MSXFsHACGCiU9Ck8t20dFAFCeKpXhXD0WAbr16416sVVtgjMayGxqXT
nvihkkYvjSuppRrZKcnKtSk97oXwIoHrUErY4xsi9+9ewebw4h5vI4uW2jzECci1NtidoSLnL3PV
BtapQvG19brWVPwenTjGyhLlAFDUxFjJIAzVpTn5Tsi5yqjYcqcpemW90M9AaY07/dZAzsCdTWPQ
J7+hQRlToUzLP2jPH6DFgGV2QpP8Ea+ttK3LdskPfxMnphCMcvL0hbwJqlqxA14soSEuxqijFsW9
JepocvfN+B0X8+fWdab+V5xqfcnwZdYnE0yFmGBCj6axiWhjBEozcwF0fH1hRKm4iPp7/XloYJt+
DnTJpCyQXoNVU2pulpjXMd+ahSH9AFWhJ1ye6jp9HKCgU1fg8eibnIwkK2E/45LKkMkpr+8To/D0
XvpDxQIBcjc61F3IQcQoX1xyj0T7oHLw0wRbi7AO+YsiTNY/iFp8JGLGcwnXQpCAgzLNDch1dkDS
AHWm/h1kCveu3kHzl/HeVTfYceebOEWgo/Ve81LLR5H5t1e42nGB1PtlWDU4ncKfdxetwISxYdB7
Q+0sU6/pey7EExcmLEc8nmC/k7hA6LSlfqlBPcxYAhoh6cNYB2m11Y+Zpz3RN3Tio3fD20sitzwj
/12eRq/VmrRw2zTHZMvFVUDxwAA3rk85H0yNlhk+StuV2DWr5vvhZ9vgy7ELy6F7cxKnPSJvD8zm
g5qKRRL2uAHgAjvePRFumGJ6uVQ/aYFC48wPCNoDP2vJPmH9sJrYPcIgOfvPGvn4rN/j1xAI1Qj9
1HdNBWU7kqnohL03KyQqXM/Qq84ReiklQkMC9chNf9OeV55TF/hZ+atQ5i6mCxZ3jm/OQ/qzSDSN
yWnasknWz297qGgWJGU6OmWA5v/naQVIRtmKi8KrYBK2xcBMZWR9xeu1xtMSQKoVW8clc3rBDqpA
vq6hVILVsvpwXlAQov5T15C/9kYDOkOG+dsVe8aS3AAjWApJ6peabHUvtqkb2pbR6OqI+cyMJQDV
opuajIjMtuozCeo4JLHl8RQz7rx/BXLMwczu1gauhWroePu6Tpo5uLc51HCnCfk689/9oh1qAl2X
mZfZyVBBNGgQ8s21uojFlHqAFBc5aBo6gWO/N6pwtPvi7U2ENBLvlWf6XBiCFXnC+O/QMk16qm4J
2aiJrBeYGB9MsQ91JyhYg/EGMakH/sE+Vf6FoOjzl6AtahUHiKOigS9XnooG+45z4Y14dkuBsoEo
IxH1RDQSYt1BN56Ei5UUPZesKICVcWvEK1WhWobllSFnUtvCzR+iXiz6dS6qhhHvy4YMhJPlxre7
rwZvqvUxt7xmN3QXXoMsXmcN+Nvcmsdkifw4FdJRchGgQT0URzmNt4UWXpW7rALPS4TNvXo/JvUI
qT3LKnOyiBRKvQvSArKXenWzlWuBeeF5mtVlFNNX0YQ6yWfiq/S4GaUSEJLanqHS2NRMtqF5oKt3
ZVKNeS51wPPuDboDfyDU2WNt/KJ6cl3fI93XwaY2rt36NzgWGrXQ94THVtiJGnIF6UjC7NRSuIsz
CXTCWsnS9/oREzQ7ig1+67LOkfBml/ZPQQzXAdpeuhB1uwx3RowuOQAVE1LA2eB1gXgiGSbFvfm7
ihCFIKZW3+cHNU2dNJC3hK+sT7TyIm95/N0azYQ8PeIV5628KKzfb3DnX0eUtzAWUBca8IF/Rd8l
1Q5MOkFKtaFo6Zr93L3DfdbT97aZPeb2D+vYPnnxZhjEz0TpbUuoJJaYulhk3fEpnlEbPSDFbiVk
HaWF1Mo5+NBlGHralL/4RY8ioDlVpL72+jPt6N84in7s3+MuGqPIYnuUlSJAddzquj76AXFKnP1p
mm1LE74WI5Vz2Tq+g9CmggYNhXSuuZtRYNIYdPOzTpef/ay1Rj6wx7iUW56MZ6mEAgewbzHU8WWE
osx3bLSTa1GD9V6WsOaGOXCzcFeQ+zY+lwNLsxMy1NtF9Rrqd1FUaWPmHJ3MHy3K1UgGMwuvJ0jp
H82/bVWGWQELJnlMI5//BNSjanl2bTORImmmz3ZPGDdl9dEEOSThWoXu1zdakdmjRrhL9O2KSsu2
ODIPs/OiQROwDTakneKtFxw+S0tFfPujs+rnuKSbUTnYaMYyXWp+hOrun07jUmHlYCBW5YcshLQI
1JHP1E3h+olV5Hmf06z/SYoYLGRK1HF1zc2m36h+PkIxRjAD3j5Ca0YfRE+8GXg4jcMxI9YTQZ83
m353/vy8NHGJ9MqcOCP9E9END1e9g3rsvTGLOnaKq9xVMi62/SuzzDVAjMZZ49coH4y6ffmFsKl6
YPJEUprIhry1uQAxbiQjPk5xedoo1pG48yHnPv0GOonUi/RdOxtVK72NnpJoNrjgvLzR0ztMSqGU
TsficuDPAeLQNjUCP6GtjjmudJaylrCUoPTku8NYlDYfcWWHc3WdCEYSBNk8M8TD8hIpIVRLPOxT
pwwhpzAP86lqY3sDCh8Ks+0FzUgssWOENbmXORL8oXQNtZZ5w0HR7a7LlS/xj/9Hq/bqyC5nGvkU
bxa5Alh0Tk1Tiv8YWSC3PCtgrA3hNYDQLUyt/KhO2O3D7La0Mygrg5ehiSdYv2AIfIx65tPcX/cQ
dxN2UBmjjTYNkjKiG1pIEGe2xcu+TOK8sqZEtz/TKHLlUwVtrlpLXk5ygoJ/h0custBqEBZ3dq/i
jQ7oICif6TD8vYThCvYg7EF1uptwMZHoaDhxIA434ZbQoMTHHgQ5uuqrSZyyRmAqog7zxh2UGEHL
zFHsx4IEGcG5Gh4fIQsNgyVJ1f6l+RMUM1+HYgtjvQ7ks+y1kobyjjpAWJbFqC6DkAAtzCNRzzty
S50yDFDEsg9bgcHOgldVMvZD/kn0HYr/z/WSR+RJBj30tmzJrvF3VUkN9/mk2MW935OEL2SS1xdw
+nTenD6tviJHYnyYQUFpOGIXlKH+eRnj/tQP3K4KY+rAbQk87/cY3lDLCMrSFsWgt5Vj3HUDzCcY
J2ZPO06pKKelNfqKj4U9+E0yi1YmKZQF/qYqG4nNzn+XGD36b1hlE8KjXfSEONdvv7OYJVbBkfGW
tOAFdjGupIzep4CDBU6fWobf1HZXwMpaXVursRFJ6bSGokrq+FWtYfmJNpAFJGIkjowkgFf3OBB8
smLPqFmmycJfmAZ04ClCAzbNpXJwT079dM+Z3gjRJdCc2rPzzFvAcIssm4XubCUfTTsI/tyoXMb1
/63S60+EZtRCY/DHB4X/N/vLapZhEgnbzo7ylQ1r1aRky7a9k7YLQeFa1uhJVy/rkBIty/HvBhkE
V3pwHG5J4qyUTKuCclYi/Wm2BE/pcOA06RXNG9Hskzt5g5kiP1Fsbew2TQauiTn88rK4PWGAdCOc
c9bxcAxedWglPmAF31ys2t4i3IWF6TCYqTBwGzShxuPF9pgZw8IL99KZe2x3tELhCHxj+t1LL/XV
HBX33PBqhbAZWr3Os0LPETb9VeVucDE8hO/yoaDUZxE4jLOnI2/TUFVpiATwaKK//dVzWPptgz7F
JX9ycZDqesCGKg0kWAB4u52zkC/CHoKR9riBvcTaklhtcXAIIBgxJTgns1HIk8OuT3kY9gu9cZ+r
mzpnCb6ApaGyzRIffnewQ23d8Alv/1lBFDbkeQa4QQTgPsHMs7XyzGCxvkwxMf0M9oFw0lmWPlNw
ofkK3YRPcXH9keR3eIAZLByPtbyUKBXuAeRtO9GZd0STMk+DJMzddXoM7N+WSpmoM06vMeXrqTpV
4kDi5cbjkKREfxWykizB3b9YmDe0H9rlY+PAydzcOHH0pV3vDK812nCv4B4yqsP4XBWXR774ZK0H
fcL6idlM+sNNJX9PquuSyZDrj1V3aiwpwpQ/HGfz+NBMrIhzYx2f9jVP/qZuOoUPFCe5LPaE8SqW
gkryLslV56UIxfJZUiFIAjfLAd0I0pOkLvBAbipYZSqjcO+mNGvT+X5DACdoQtVwu94kgn5whO7Y
2GafikFQ3s/83wl7/+l4iVRZFT/XRQZcOqtO5o8w4iUUXh15FHDhE3MwCh8mtEON2ylHcwXas90N
vmz2OjbRvWd1dhD0YZ17aq+R5atKeHnah4UowVcCyXKp1lSyavvJTvH9RaNTVWZ2kXIOUstPEfJr
CxdXEQKrLDKJa8DRiMHyBlnaUAsWhztVmQKqcrKjHQoandBjSXt+yBLahWfx6k0rPvIrV49/uWE8
asLOj0T9W60ktcCsOtOIvcInLMvMwfRpzOBsKCa+4pO0wT9g9P0WCCj7fZ21Y08R0VYI5Kv1s9PT
bg9mP0EeFWWSdmrR107Na6TmM4uXw+DtOljN39bDOUyW++32eDXd7zq7sctZ17RlG2/KBJSRXQfF
SShsgGsFg2PemBS/Wp0GXr5WmdriewVFrs4J3MtNzCJKBvyfJnglaCdNgPmEnJvcGi4PLTlxZ2Ix
YraBpk6QmmztMZkerALbG4epkduTMDqnLY07gwZjSx4gl7NoNisD9AJJGCikR8O/cCwi8DQfTTWD
E/2z5LFK4vdxaCBWpgjW7fa4qW3BSyZCDdmCFC6hXnfNpt0kn56aSwL1zQS+khI7EQQx1ObANkWY
eQjoMCt43jALHC+bKmAyx+JsZV1QK0WIlzZGLP5p8bHraRFTjiiq8IbIrI4E3oFDgVYQ18dNp+Yx
JKEBNg3nIt+43k7YGOYp28BzUzKkqYA1ECT9akeEJmNeL27Z0Kk+/40OUM2jKKKScqRphqdW0wjJ
xOnrmGPwoymz5KdPkgvMOMhgVnjHXTdCmzy4QnVLcYdy0n0MK/Gt52aj4IISppcKXVbK2mMCSOgV
abPOZAZna8egnV2B9DD1ZqW210imcK9+eRjXBKM532TxwMjLw87glIi1vDWwhV4Pzs5uIE9TyLtk
t5I5Hd8vu7BRfpoU0LUZyZZrrfATZNvDlnkoeL12PH0J7FiGuUg4//iC+fucQP01gksvZpHF46K+
9qwHCqLz8DU9omOe/El5vRamKhbumPk6ifRefoPFScG6KSBXJ50lvzCv2BXyja+LE/QDdyH3ZYGa
/1h+V6QuWiKowbtfhgNZ6/tb+s61OtjnyIhxmS64gwORhpkhTqeNuPsKhvV3ng2OImn2GumEzA4s
bUjhYTxPOOF024gBZB+nwYUz2bDIy3GTgCzbhezVisXtcr18JtyZGbzlhunZPRNj6zbbt8eJJ9R/
SOhmN2+VRrOWbqLTKX84BbzJMxfs+1gNxCBr6p3wRRy8FqWIHkQZb3DdUywhyClWYMUW4CUhwApf
8ywRsTt0DAEIjvArolB3rcsK9TWYRbZd7cC14XngUIGamH5kkpWXPWM4RLg9XRiV4VdzA3KCCN55
MYipH+ATCJTeXJvsiZVliSuXak/31eQBvREmze+nbjWptq+rJ16MnndlNLIshoJfrbJwGaTIgA/I
LwvwKaBnafuXomLpcoI8SRH4aOkH2d2PiVFCkWyumVOvPTe+Tm11bZsNCShxXSiudyx2Gpmd3Lmd
aWzZBKxoEJRaFC2RQyf+3dIrCGUm/OOTQGXPjnmJohsQdWQ+EbwaKIDcWn8CtaxdpShkHaiF6zWP
Jita1zZMrXKlliOCijA+KrC2YtsK9pUoOTRmG94CUXJhoJy46VEOk92ibLOxhLwRstqJD3MHBS2k
xC/QVFfsMzP8FCnnRbN6Lwu7i56FLq9r27pOvClY8s4o7Aw7Fa4J90pgNqJSD2tOFcIpl/BXAxmh
67kWff8pXkWdXYwBy6r2TwoRwfzyZvaUZy/ez9hpgU8lOCvKawiT8Y9WRW+HVY4ht1ZHDVBkpLJr
dAA54l4scBDlsAhVlu39ZDgb2lEnSxRf6YIv6+l32Er5LIcr8yuEWwCoLYOTkqoFmBhjv1X+CIac
04a+VE9eG6UQbvBsgoK7HjpcKuMgmTN1kaPQNPk2usZH59BssC5cqjM/2BDQ9gy5Mu9PFBN1JqQI
AUZSOBTQ7HpfEbuDHMDANH0by49AO0/mO6nC022ytKTPYz8a1k9k9aSsSI09K84Y6DxtzV2MHrqP
lo9nFmKcC4hBZRlvzz0c0Xc+1M7p1ups3DPDOVI98mn85ZBDKDW1NSuTjUn7QeSav8dhVFpqo7Ep
Qb9G/Qu1gg9VW4tRSU/UVWztu+dlHNyzL1lBZhB/48TQlnXO2hl8wQqVWvCfqpfodjwczFkShWi4
l7E3NfMqMw1jyyNPIZdE9WHRXEeLrn66R58oLGWZv9OdlTkldLnPyJJKWKPhn1zR14OiL1UhXHmL
+0eB1Hot9hnN7I+hheKqdLfzGnShyGJAnfRyG+W15PjmdUPv7A9oK1LofueuMnCaDJcnmvvo9ZhV
EoifJTyKqHxLuUAwBzRpXUzWMXL5iGyv1mhVKqQymFQOrj5biv5dm2oP3AHzZ60AZ+2Yrpl9JsIS
qQg2/vd05NImfGAjhKcjE17qt6b50AYs+eb+w9qMIuuHHRKJn17prK7bdduRP2OPpsdXff4YD2ZS
nmNGZYd3XF+lsQgT3qdT49b82zDdqcn3Eo+45R7F00VjSjn1C0Pnx7ULSO7/kOgd+HWYjMEGrySr
j4JQd+GNkhb6MoMm1M4FvHo0FjV9+9PYkz9/lWCykl8PD0BCMoO5W2SnSdi2iB0o+jO/8w+Au0/8
n3Vwi+wHpFSuFKnVJ+QFE3fOzzrM+e01+K8EGhXqVJf2kBZXhLPRRsJ50+uHgRd9hJfytP4Pzm5N
hi4C6AZkZ6X3u4m4wgtmOeHXN4OChU8GhWJ1cCD1Ox5mW2v1Xy5ORqdBpI/vfixlZpwJFeztmBte
DIQpjpuDSQ5Td6/VqVzK4XFCPp4btJXB8r0G4W5hYzWGhN1bG2WbtaYSNcQxj6xZMEd1qSavRBN5
M29/HcQfSAUnxlbJ87Eq4fo9pVjva6XU5kvmuwORC8xq2nFVZQh0Zogc7uDdrMVUQrm/5Wz5Cfbi
/AgHKLFVVwzJndnUv5NoCX7OmhdcDVDRVwW0QXvLGnoHs48f8Ksvv8DvFuSurFIRzJmXFm9xOHeA
Na4W/pAYEOqQJDprY8F8hJFt0dc3P5951RNXR3fdG/Vk9U/24V/UIZKwZILg9jy7RWTKNvuhdwaM
UPb+i5wst449N6FmfE5IWpu7T9QlkxpwuNkP0BzRZNR/zS1ZRtMgW3UQTpkjqUYck7izabIzHgcF
f+JTg5PS//hl1AF+Cjqja0cr8mpxNn18pPgNsaFcSRnSNI6xtSM+d1MMvisjZWvIVASwOE5p4D8O
3oJX/UxELocQT9cnLHYeUN+v7wgU7+gj6kDnlsnBtUVyQXxm2+qZYXccA4kHQaiM9t5OS/bnvXuZ
Bw9I+vclU2ZBBPznBsPYK+bb/kDTjP7Qbxk3D8ApKHOf9BH6drcWqUuDQKMCl8Oj176qFRPdStLn
8HKXv3Lw1vCIHFqkyiihH/Y6td3FOkYjUj44zgxCcZINbZ2AoumLtkmbkT1qtZyY43LPtR1Pj8pD
VoIxHXUoyyUQZKm+qIrXTfvZVQMMX/p6D5xkVum7XD+GpHHNSjGnvKHLXTXQfdtrGXXHJFxMLEks
wm8ItWgRKGzhF0htR8acIL61/Um9//D4MqO3e103gW66zuwra4SguOkMLqD5hkjP4UTqLmORqLoB
f2Zu6IBPfFgiwWHBQSIW3V/pP4aUaS0MpzFzvqySL8kqV0iGHeH2oU2hzQQl+bgUbwz1KzPv9Tcx
2AHSY7+Tr1j6I/8SCssLsuG8wZiAJoafvdS/vq/UxYhbyafNaFImsQ5j9pLuv+p3VbkVcMVti50G
uXmcvf51WslK/rY/AG50EP1NEutuNzevMktVMk2eTbeVjTK/zCxi6Q7HC+wSVyQY2abqfuxMLvEw
Igc8tJYFBBMIVqplny2zBFJ9N9I6f8zlwgOSmQ0C+ZkOM2uP0k+HCMSc/Il2okxh2t0FzK3l7pl0
yGCMH0zBnuJpQschu0fecHFuDz8S3V/M7q/nO7wPuRfMbILzIExgqAL+0lISBPluFrkys9ueBsNN
9t3kMCiuSD9Kfv0jyNCkngHc0zUgYVgrYijCi+1Le0HLxhb7PbFlbwgSO9Or/hcLsI6YB6un/oC3
wLz4blxB/6j7FtGUNfPcRIyxv7UrAdghVOowA3zuwoEzmdI9JkMCBh6qIYsb2qv8aA1xqXkeWqBz
R6tA3xD/588IUxgyY5aot7X3pV0ZSwZVdgx95SOKiTJ+Vr1k4uqLf+XmDcHDYwxyoKgs+8krJqtO
WNFFf8ZesADhFj2UYCXwHW3ZcrwGI41lDCuIHcry0FYoqpecDUz6RFVE8N1dLorNBQJgW25xhpRD
MGLGFegPY7ffhu7FyDqg4ke6JlAQsoKnleTGDA/oKIrIu4Q3kjpzzINHdC4hD4f+MlP7XuiO4tvK
953J4Qz4MQIi5w3c3HhaG40QhSqvQGxWNLX9QDqZ+Z3dFUo1lHl21XAe1L7hQIMPaQaKeILEom+Q
x4ZDbIP1TISHPziAgiwj7wLFLvwuNFHHbor4dgzS1qgEL6QG5gAi1woRijYUwwKbLQev6GuVLo7W
XOly+BJtGhRI1NPlFilT5eaU7uukIKT+32vy/OBcFa2+LhYBiz50mQZajNvcbi6dyEzoLEoKeLA9
Xtz87Pvu9VEJ/DwAJxtaqhh0+8ARc+X5ZpS+jnVXA4ONKjSGE8pjUEMw2ex7f300WIwfAWVAZ00E
1iXlJc3Gr4WaLaZkl6DYoCaX4X1FN7xo4vC24TjJR48TQZXiZu27im4qrwjrzMxPqwg5TW7bjzt9
THdlIMx1+N64ABRH7UD6aEUDzKK9VO9pf9nF0eLuK+PLBuGN3ExbUb7C7bdGPHISrQp+BGvuQpcZ
o0uvaXeKBqutPs3ES0p6matis4I7YTzE5SG/tJ/QvpoazIiAM9ZZ/bxgrQJCf2sfOJiWXWeHfRQw
Shxpxj2mFXFyukGxtkOt2HmyH7FMmyjGtCoPKb5VmmRANiY22yuXEIxDDU1mbyLf6za9NxcMF3hd
rBB2zK7ESlM1PKrCZ9uQ/KdZVrcfTOtD+5noHk52okUk5f3M4+UJ/ki9z8Z1XvGF9p2B5qB5wXuH
sT5EqvLbTWFdpEpnHYe+QS76sMVsDUrWhD0WHXbjaWOp2cUR2I3BaqIH4rPzXGli+MPzgTItUHOA
+JYw48jxLPcLndulolwCGmO6+QuTFneeA+xEcp6gtkmvdawA4NC+2FsJZ4mAawYHkESSxUKvEwi5
ZYr617ymx1GrRVqSWfRRm29DDPWq3bYlfbcRLvKcPlaP732wp6ZsknnsowIOTcPlhSGx6Uqvrg3M
xS8ZOqzFX/7knkj/awPhdXho/cXEjsAPUVIr23etEbrBQtWKUTTlfgfaxX/dih4HB4UswAN2/s1w
KdYt1Z5a6uoBEy7MlzMi5+40ZmgtBepBlWQ6iSCPYZE7JwDxgdEvxm8eTj4dqbijx06QA00q7rDz
7251iDuPPjPOClc83+N/QcZzmrQ5esJWaFeb+UMgxM4Xm0jShVrHGpA9FNjI51MWMYxMuWfmzZWc
zLz+C9L8cV/Xv/7RIcPMaLyGMlY6iCMF7fcOTr5xFvRrezvjqVWjCSD8i1Khgpcl7wFizh0eZC+N
3IIdnzFX54//6JGRRtcdojZ9S7InJVOdvCoIhUfkobBKWdzwbqOhRKZ2m8IocDQ6J8wL2ECZLLTw
rxLfyxBsBJJ4Bx5u6cNpnnrJw4eoyFXYr385lSbcN+c8AxOw8O7SviHFHLc14cDK6bxQxE7TCQli
fPUZoezxjb3oMTlR+RmbvCHNH8GJ9i7qemEjXnzL3EdkXD3973PuahhH9/Ne9N6pWbyUWML7rlRM
x10qbGItIra01TdUb56+gsSzDQdj/uq5ozY1sHVRi2uIulTzXoKklETwvmGOiP+JcSEG59kIZi0r
V6HgN/cPioTc0hggqj1cNiKpxYO2IXwOCC/YcO9tisZpXvh78Er3Z0L/Co4GRRtESQ8kdya8z8ia
0jhPERGZaC9Eyk2pfm4sudCypJ3JaovE55g+pnQvcbeSDYOIbrkN4giikV04o79XqYKzx8X6bsTL
KueSubK8gMWQxeY7WR+J5pS6lyhXv9kC0ajt3jynTdI7/WX5AYzYO7WRPTv6vCQcHctxDo1fnhzF
GwPLrcG8IKVkVmaVhlIyRW7Dw9ziIv0c10zpE0DOQJ2xeIAeyiRPecaSEBZ/3Gw/4a799XXnyaJj
bMx7RcP2EF35s+fvdTpj1AFhfGUNNCg6HEp9GO3Oiux2cZ6wBLeApQdfXe06FdMeDNoPHQp2ZP9t
Z2l71mejBCRg/WfzfT+RhbitVRMSaSd/mgjVfFkDG4UnacVQEq4C55GMTjBlheKPMD5Cu9npaQht
h5eff0OS9IjfYPw88KzCX6qUheSZDUvcNm/wtahD7HoEl8v1xmhUpC6CGRhfwBQoPnWEAdYBbQQb
EhKgyJfRvjHXLXV6N5srlqRNMkeG/3s3zWKtD9AqwQhk3UyJKVbmhekr262MC52BY+pw3KddWqbL
DmlwJd9lDeKfp5WH36sOCyRG71TtY1DBJpBMJZ7ku5sZ05C/28MbGdgs9UzuD0/rvCMU35W5m1Q1
N3dYcx37WzFOTM0d7GTqnXWEvLRkuTrrZf9S52vBAwW9ua8lbafY9GAaPACVgDRlHx1A4w+rZMsS
62vmH8KuIEZ1+eQIBREgU0FBDM6sJchxYK5c4eojCp1a7wBxNjndKp7e1tE41EsEjW3bOy/t9xYK
N0QJXLyM34LfrId9p2cMz//87lqWJaDZ3+fRXlN1zSpQqGtvvwmAFu0lnb4+o5UvSJJ9hiHB6rlI
r+XVosGRxkFTkl77pxRpbmiga3giRIySZqiV+H4f6vP6SJNFNNUwlxPhJDdCvQiC/T5BxSE6Ts66
0Mt2O9rVC2/Bq2wgX4PMsqfHPGVNVHHhMlWJGlJOAhD3DxDBG2492Qx+IHchZ631EOcTx17MndlA
1OXSt1xh1OW5hW2cwXHlT1Bkm6tCiX9TILCjdkZWvdWBapOnbmMTa7u7r74g6lL1QPOV4ine0/Hw
X2bhcAjTLvve3Ln47iOvo5WcIMHcPnWKX/ibSWSLKF5630eEhjSiUbGLL4zetUUYzSRfJEBTooE1
ZICeKtjZkBc1B6H4nThBZvAawx71lqlQHIW6dHvR0rL0P0jWfVTGBTLo+r+SBNTCHUNz3AoQ/oBq
DKQH5PnEY2g6dKsqqiJv2k4ePnAku51h8R8SbUY/LntZp+3n6I/t58VYXMc7rhR54McFnrMUvw4H
hIwi7tqXxbz2GvI8PBQeeI7lPi4D1BBtDyqWGODcd0MTSUyyLCrpu41nWR/jftk0uOEd4dElN2xo
pdxdhf+H6+gLdZdflaZUEuiggZuqOf/ArRDqZ7bf0wfNUCOPZ/nywgcIh8BuaCx14+LzKGE9wJBM
8lXlAaJ8rUmOuEnZDamiZlHKJI2GGXEDXgoPvAfapWACVswPmDl0wEA2E/W+BNXmAVEpYNhhtskg
3Eycvs9gtRk6ohh6UPtluQGt7zO/1MH7f77u+R+Yj9dbYFB8GUuGIqOnAm/HCmd2H93o8Fsm1cUQ
vDcjh5j9yAo3egnfALi+tWwX+rCqRV5G3mKNIg9qlgprCO3V9GTSM4Q+ZjoocYAMGbL5UmJnnALI
hD2AYlZo0HWUsqohAGRxlMre4JNvNZp5DxfBj0DWOWIOuyTeH+bsu9pV6XmBNK1yJWHK+Uip52jr
QpEjlCZ2tbOX/yuPv3IbzYpgY05HsoVL2CzNTKVv63RPNLmzh8jetPFJDxQc+sqQShzXIEZKGCge
shZoNHNqQ6aOelgnCankUQgkq+3epn6peabMniBfjBqIUzDqHdPJqjJVQsKlrqbEmNfuvm+7Yhtu
WuQImkAiVEgNWDhtYHBIgmhnBqFlYJ0fvs0PoEG30tEZXwjdqMv0sEA9FAgV7lodA21LRCi03QlY
C3fJaaV7uB/yLOzC9qHTWQppyVXR+iDbToqQAh53CHczFqv3kgcMVogPrOvKcTmqT4qYpJNrD2nI
33YfsDcsz1fnkN27UCZeYa5VnKc6MZztEDIPgyvB1XfpBv+0jd+RR7yAKu4lHUZDoXg2fxTOj225
+OJOrdkg7U0mRkxkZhMNhvGr/liKWX3mcL8Oh4VSYdRTfSCGS6l7uZ+aFA61PEqYn+k6iOAIXVJq
bGqkKp/+CtZ2eLusHdfg0D1S3IW2KuNuJ/sqCg1vY7+N8VR1PZn2Si+2b7r6soAkzoJK4jDZ/enG
q3zcIceLIIphohwwKkM9/5OSeuH09ZnwT3H0MslXJXGmqs5zB89jm7pID725HPvbJBQ9q0pnEN1I
NvOCb/U3v1cFnzApdq7rLQaTZWuwxlIGtrmOdXh9MynEn0xAQxxWf780iWxsT6mw/vQUEBC02VGb
oi274EzHPqFw/4jcID6qSuZ8TGkZUS66+Zt2UcT+DPKZKdJvvBd4W/uoJw5J6PJa4MebRc0jECtt
UTXphqNvddre+5d196ObeHbUVclmt+WEhZ9F2ABrVO/6+yyL8lHyWuU5F5WXM7vVd4u853XSOxEr
ZcjqGjcOWPvkSh70dMt2ywWTPRHX4UlH8V39rJV2g/Vpti9hRPEZrXnS2lDd3hHLnCHJNRQ7C6os
UI65zLJ4XM0U45tGB3rp7XVbF4rTr9D+TwAuIDkFv+RXgWYyr2x7zbJx9RvNzbpSgdw3KfEEtM9d
CAdKZTHeoD/+Y6DU1JCi7ANcOVOBqm8Szyd3fnBLI/h9VyETO9BszGDL50l7y2mUoiTdDdFgnbkd
NoUJQPVg8Fbr/wXjd/DampBvZKKiABlfUDeMJkqLYS+brP1kgbWcS31k+dKylOsmeZoOKWmJF8eV
2/fEaedjPPZfOL8M/Zbsj4L8jKgK4S/3wTvLggsu0FNGHIdQeB/HO4lM89BOJzlLBDzan+8g0piH
DDNWBVmtLlVmSIo3qMgf8CduSEUfWLRFINXaqgzjTFpWBVmuEI+1a1ThTyVFi/FLrbKoT0QPVzjB
ngV7JhmJDXG2YcYzxdyIZNlRNlTdajEDaZQHhohd41Uf6/xHTe9890rIyYTdulK1OXdY4HmDgRph
6J2URMheNOonDkGRaTIzy2FTwP1dqEuwiliuetbEbcF3VeP1KzLlSnPp8uDZFHVGJlz2FFSP8Paw
MrcFTZnJWUqcHmYgmY0HiqKfa7bixoJ2lb4IccFaD5MCq6HFkWcUNdRehUbJEe4Nw2FD5XkZzZnx
umCrHXweF7PM7d8NT2OzthFg7UQnghVLoo/j7rUemk0R6CXGNRdRJyyveJVgT2m8FTI9gLZH49Wa
3UM85SLezt+/sL2phZ3c0np1jSUPltFkpvTDcGKK0H+SUqk+XCyLhwWYT4L+1ZAUULZhs0OsyTIH
tFM5YdNVoth1QK6HNebwRe5GGzZelIqpYxaCfW6rLe7a0N+JIHKG60YFI/hKjkiJIqS5Fo/eSvwo
FcAg9U6Y5iNnF9/BbjIhJMULr+HuyUuVsezqV665ADmNSns8KvJWt7bUqbjN3pYIxUg3zed3UiYM
Hsawg/SiggHMtHevZoGoxzQZXx6Mzfzke7A3WLXAQirWyd6e/dCPnvDgv+ZukIe83H2z6ITdWgHR
upDF0C4xWmhyjQFMZp0re7KiVJoxSCz7zJYlclUofMl9FByugIoYa13AGQ+GJtMo2W0yYqeHG2/5
YMDMarfYa4dk8m1JnB35AY/mhKzhaf7S3UtGi1wAQB2358BEeTiceif+BxuRTsuE9gOJHTZ53kJH
0rpxZF8MrbQ3zl6lRsoTWhXaYdMH28iBbqMUblUCmj0AA128Y/6nuo+CL2MvHAfZ1YLLCjD8o69Z
aPcSuLLOmLawY9iHyRTCDZRM0vQW4e1rtenoa6oD+oVBD38kq3y/nRuVyDXHo5bkvv6SQ8oJ3jtw
1l52YdScJq3Cl1h7tqCms6MHEFqKNyJWtxeazvD5+RYX2PVN+pDAB3Wp0gmaqPSPFXNiV5sxRkN1
hGxnpsUHTiH5qooRRc2clkXh6ihgyosKt4OYyBvicS/w43SEYqbXPaEsiuQA0GuxDA238sozg4UA
wdzYwNuZry4MtDLD94gv/UUOV7ZBfK0xM4Q6FS055VrU1BU3S1+k/lU30Am5vpDBaNJFVDliWWva
VVv7Wvd/l2tOe8JzOSqCzpe+C2jK1qlMElduSom6+k2qJOXvUAfcYsFJud13MMW1/+N+eDhe17EJ
2MjV5L9/K8mhEZb3HY1untSm++u7ih/rGgR1qSkltVOBR0fvXuImS8+jdIxiJvz7QSpC2ApgOCig
U2f/QGXhuQWT3S/8FS5VnoLRT2e9YlhoBZAAGIRF04iqILMTIaggBpVMUh1xfD4PRwckqzlVxWGN
BlEqO4+RKD771kzx6sfOAF5/2pqfSrQmuNsF/oj1OoMCKfVy6BSCd+92ssSo0DOkRXGBO9d0P4WK
ObcvG0sCk8M1FzH2nBdQdA2pyLX+AJV/cKzZNPjPtp7VhDb3Km04iYvvpv+VxAon/+AMljeYuHU3
rq9HPKrPUFaF0r9v/eCN96X+F+rfyGROxePOfYedOngVLS/d1KqnTB4YRwtUZnlL086PjWZfW6nH
hYE9nXqb1NerRlWsMTenA2f/+nx7//RbckqN6HssrOXh0WqzEKUNy4x/a+NfN16R4ZjNDHl+U+Sb
oEYPKiGDTulDSr+lukVvvu3VILoBY2qh+pv50G5jdhR2MEmibzY0Zef7Gf3yKnb7EKNPn6ldCuWU
Wj+/l80sSW685AchPXMyG27pgVl44aYsfadTmOTKB2HEFCkv+4aBbZWzgjJRa62pqu/ZaQCa3+2z
h55dsK+QXBBmVkOxTuAoo2eDq9Wlob+bBLW9o+7kdPMpMmajiOphZOhl+sjUrWWi6tTM/nizJAV3
aWfYVimtiAcICRIyUSuoXQSEbpjhQ3Gc01nqCYvvcCGrC/Zg7pIaPKzbwqUTtZuBDY1J3YJ5IaL3
ZZKFLA8s65tOQJ53lJaVCdluaLw0mjFhiNjH2YQD7/fObtwJq+/xAA6WWSBgoXOec7hk76NbIiY+
uXJQlVCg9gg7exVJKXOIH3Zk4Z6ZwrYVxsuEaJuF1yd8LFeb6u81hS+yRx7LM0iwK4TMbTzeVBXT
3ZAd1uybV571VZetEbmOZ+qy5GO4EwWYEJQg2vzqYpbg/BYwY+83RRHxX6Sx/czKrgV09DpawZU+
XbdzoTF96OKuC1e4s1u7LR7LphOQcm/oYaJfyus/4OjNJwG/GsxOEqDOnzwR1kccf8jNZuYuclNM
pwqtU1dOUhwbFq1fElZyCATh/tAyorbtGGl4m9e724A7Zk1Q8yq7E30H/x3dIFar462iY0XJPFMC
VPDculkVrSsRBtZiVCo6aboKittBUZTQe3YdCN/Fu6oONjTmo2qPT/34MOl7zZQP+/YVRX8ALdHP
mWhvmF2YXxcCGDTIKE/2ND6A3m7IVfz6Rk4XX7HpXfvEjyp+JWfI/6nIgtkONZkwf+/PwFAJbaDK
18aYeuzXtIECnRYmEzGuw5sHqrnW2RWT47/E9n+QOfo6E5Fd5QJuQbkyEus6LFK51+z63Hxyto29
EY+1B4xYEQ20VUCG6Wik8fEoBJN7RGUv+eqpewQ3D7yKYzle57omnde4xb/Xqb65l377cCn3wlc6
uQn/FvxvDipIIH4giFrJ7gER3lwuZB+6XmOIjKfd0+R/4/z4zk3VD67QjAF91fPl6f71yGXHbHKB
+54S5dcfXVu/erJ5E6fJFVL+0IhVwdRjWRpGMPLyzZff5VVAvT7/U0X7fSQp8OK7xL4fnY2K6LzW
eFLsq5L+KTtWBErrINZfcJ22E3jXgVBCDsm969fPQRkKIbKa3HK4yzHrQsfxhVq7+P0YDx5lGVuY
c6mi48SGl96tzglDbwV3PB/x5c3/Y82TC/IfoXlL6qhksSOqfwcGbpZ4zhtQ4R/MfpJZZTbEkrjD
/T6jaM/biWX/W5Ejou6NvwSITr2NJ2IrshYWLBVKov5c+l8sIVjbaZkYnaCQ8RZsND9lk7/JuZNp
PavMtvfAc1MgQagVVe41r3+h968CTRQ1wMC2Xcg+rxja2lkNz/cj42n2MRWwIhWb7qEpTDUHWUXt
3qn4EP63Ofu/XvgzHEj/u3TK2CVW5rZeOAc01o+Qaj2xOGnmRmCgaylG1/k8e3o/BHUM2vuZGMdT
x2vPsFsA5Ebr9lT/H7svTBWR8blliw1l8Cf9CNvztGSh/Z7gr+0q43nt38o+wDVqXtF08VllFGVV
H92Dfl8iFlq32Wmaiox7glEYcw/RvQjEEk5bkq6lK2kSQWZmhw6CuPxcpA9N88CT6LeZYnAf2Trg
WW0QnEpS3G2xoPK86m8Kxw8elVrfn5sEoUnPIcjp4B+StA/zC0UBMdLOVrb4cmlkj5bVjToZltPC
QVGZwkmxIIBlimUDUXBUNcZXmnd219zeFBdOHikx/jzBsZYqkxStiEBEM4ypQSHkATHlrO091zmy
t5nPv0ID9Bak64rkkl5PUW3kEUWNjVjU+hFxN1xxsSMMhMk1WRNob30jtkxJbsxj+ye1XhlnwJNY
1GrkFrACds/ceFYuupv7CSbsBPNGtII0bY00w8IM1DBEmyEA+K/QLAY/qH6yRZS3WFJPyeyLcsbV
x3pmW5UVBu5GQKSehNOoqTgzmgKhQ+Vh4SDfjCeVOLPNFs8l9mo7pKcsas+OWgKqonyUvTDNy8dw
4jYUF5RRtKgEm+xg4h4z/bsdRw8fWfGrfIp2CydoTqcIHcTPtFFLFleKPh6YlzjdimWqQVh9rkZ1
l/tWn6pVAneQsbQ8+6vLAmMcOZ1FewCjHz+RRgaVIUS/Lw3aS7jJ7eaaZP9n/cgpj46z9w/PsTTo
64c9RXWegc9MVictH278vy4ZLLKUJlRoKFfILLfOvlwICsU0ja9EndhgHXBVj5XnjrE8/VuQvsMI
ay5jxuMgRmm43oNMgVoMp0iIBUgN8qlGadEaAuaH+iswKd67FjmRaSLH7Z0ZKpUs9w==
`protect end_protected
