`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9152)
`protect data_block
SUyihkNKvlx0ECrL79FnWsQHfTpVzyDJeh4/XJ/Z4WotbcYAlVhZ2OtUTWDavem5vZAep7VAIIog
2V3iSgBQUzs8cFBstXIVcMJMcf6mkx0g8GAGzgh+ULoaq4BYTgShH75bckMTE5Ia6C4UjSaGawNy
ICqlL+ogkR7oidbd8Jth2SHVmHGF3IDBLgrJbnsvMyUBqVvwTIHz72x1PamaVRFsakFbOv9h25j5
i2WEIOjpL/iowyTSleDHaNsEOx3csrCMVSsb+ynQibTtX5+traV1QDZfa1sGk+beLqpUuFBmCHGt
Zb+3BVeA9OwSzaDG7oHTa5wkRydBJ62Ba2DlJSjWXiTvKQ/Jjct/JFo0waBn4igv0hbQ/PIM0WlP
XA9m7H54O18wSIn+KgTq+A1s+xarxowLohQjJOE0hl1mv03xFyqXNRXBthQfITqCf8I5ApNZMIxZ
ZQGfz+lq7/7ssvIUqyPa5IXDgBUwr2UQzqQAkvl2O4D/5+XoG4S88uND6OK9VKl3Ne+8u0d4TaYO
kKrGcgXS+uRL85EXA7Tk9KMTR6UKuEbK8tmvZDKANqF4rrqdNIxmAu8s9mSCvFqMO9AIS+zSq1c1
AVAsjvzz8LE108mFdCCTcNarLYocoGbBWgbaGHG0lI4GE9coDqOFku3nlCcwMrRxetzA3CNA1/Ye
lI5VlJVllsFk3hn8DHlFNVxiRaPIcoXn0RJeoafsrRrxOpe2bcFLiR5HMhdhu09iVWcKV4ga2CPv
EywElKC/QFQk9Wrsa6qCzD4W8o1mNec2D5QNHvKDzXyuVokRQHM3S7lB5IWBJm20dWwvhCWO8gzY
B4sFocU/KLa39NQOA7s7MIWmSRbsuX3kDr4jVEY0MhY9lvpG5W0KA5qlKGMinAQNZwi0M356bJO9
z3+iI1Z/lLXFFU8zuc84BZ6+HGFXz/Q4weBR1BmMJ23uQkh6JicJcVcZ4DPL1NxQdB1oy7HuXJGh
K6U38QrsEHLr9iVJYZshcy3uGfv4nEyE61dPkSxtft1ZvpMgO8bL8epEKxC5EXf45wWMMcY5riNv
h9vje1O794lY7igi8SxitG4ooz1snm2nfFHOVPBO95ZFmn+9QJtozCwrq+kBJwamKGDorPZYVkMa
SI9sKvriEmDapeuX9jIccHUYITBVVrFBiexWUGWH4fJ9QHk7RYKKAaqzpe4tV7F2q/wX/5FT+FMG
TfTeckIysx/6T/GQKzpiBLA1l0AITv/olaLToQYZxXbHGC7x80K3rFGVQQaPypZFshEiAMqI4HOT
HYEulqerLkbDcAYeVAmi/OSqjHY47FG3SifG3a4v9PFPi9Vm+N9TbZC+crLqsY6RKGCEJVKg0b3c
ds9IM4EXnk4Y+QZHTnhsGRx/m3LMhbP9DsoaKCbEzrqdF40vD4EPk6nZiBNfNtPcikiKTHxTaR6n
2OK3xz/Yo+SONZITxss4uDakaviePSxd6F/ip4Mp+jwXvclzrmc8Wkevm7b9gtqVp1lZEy4qU1Rh
0+GKK3/sNDoGYR2r9okERda42Farnzn5KvS/UTXFavguKcM868T3wGzIXUQF3XT/5uANogttP3Tq
2RthgNZCucdM1mh4EuUtjP4BLzC70R16ZNy0pEDTPO/T5m5ExxtV+xKToYXh2FVOzKZoUrWPy025
qlsMuZZiEXguAnaCPG3XGMq6ek08Ms8vNQywteHiI+sFyLBXfjE1XahghGcdOs0kLEzZuM/EbLMT
JMHLvIi+bai7uLT80apktGHwjFdyYOnne/dF0SQ+jiJoKswQRkMcqKhmb0lcT7yzU1wvVJjKnMki
GJCipxYMRsABL4oDv2OzQxHHNVbLePIdzznGC2DUidIpzDbz+ZD6fAoQyf07zLjk4+V7aqe4AlNG
sSt5qXDUWIGirKLEU+UmF9monFEQEDfQf9PdHSC9N8QhUV2yEvVLRbb9c+V6Z8ETzTHmiP5BfKHt
qPf+fxp/P0JvNNBidiGlsPH25+wV6dFu0pPR0idHA9Mr/Sl1NCxrKGjHMdnTurmBY0eEdj1/fSoK
u37pAug9gLH6eJoYBrOviEnI359wOcqD82S8HGUwkuL4AxtHw2MUjW5NEZPGhxC7SH8WN0hIcbBP
I4qNA9AOwJriDj5FGxDj77yAOISEDof3DFWTqcg67+XWNElqA623cgydemjtNwyBghFypN4W3HwQ
j3W1m0o/hxv/sUfmz/T7jn6SUSPdtfIl2ujoNgpLl4raXEhmmP0X1ZljqdliX42Hk3shtt1vOwcw
h0IpO7SEr1N3GkE5INcJwiLdKBJluutO/hDPfyKkBZ/ZOQtUonAJhM4MdnjTJNq8mGb5d6QH/+ji
hN72C8nDqv1jsuZegS22cE+zRsLRZmAf9lWd6IzsMKXzKPe7p99pgdbdN2UMUEAvtsPEaY2TlHAj
UyD/kLnJ64dGTQyHPxF3a4THRCcEqK/UCOwwubo5w/k1nfsZU82ARGy1XlqAiVa8Vgk2i6iZ2ekj
6FBRpNb6cigRswAlVm0qSRrHNe+v9RQaYbP8ne6DeSCspvjueGHkAV4EMP1OHt4s0KyaoaGsb2lw
k7/CUAT3RUby7e600qyoUZ+juQD+kGMXOmya4xT+V9WsdYAVDogbT+MBbhz2rly+vY2i/SaM1pE9
5FM5ytN65TsOPRi/nX90jKUMhCxU66aiWw08tkriqB+/7p46NTxMH5v83V99wgKAOFND5rMEvCSu
3p0IX+Mr22/QkcFI0c4HRFBO6ZKvEZgDYnQIqbSDJ9wBIe0/01o02l5t7GwgWZY+tsvMXVUUE5v6
zDvorA2R+BuW0itOOmPWqjLxY2IQhsubayibWfc24+T1SAmUokokDeg3+OzIVqoaKNTkZexXwIPu
Dl1HmsjlK6Wkb27c8feVv8yeJeJ87ehbrjc/SmePuPoTy1p/Pth1l0QtV1/raYbWXOmLway6OxV9
uio7NdMtdwrkdDXhYTY2SALAgUNd0lpNFxVot8EwBbrplDsaWpiHOX49VDMoj02CXHCD6a0MyULa
tA/yc+DKbgrO0ag5rY5UyI8YCSq3GuYQ9B6qTpo5brThqDVr/PifUMnB10JWsvTowKNYO7Mwabys
zZmWTK6Nk8CfnOpvuIJnBlMahj9VXZ6bacu+6L3YtWclVEicAoxid2xj40ohNGk62PFBcFAelywC
qBqNz6XctY7Wj6FgRPr9t/bMZ00fUT4dwhhn7DdKzojU9LpwV/QLcT1T+H36rhSsILbdnXJIBXac
xXHV53ParVJGVStrt5QsxwC8hJ/+3HGiRHeKctEb4GqPlam2pwmmht1skkYXmsD/w3EY13iPlQUB
tJE7xtyK6+urGFCsXTK7QYXaudI/GqFNvBGYI65iDOWhyjsjUL7xSwPBrCoWDmwGjheF8IX3kGXc
LxSbcPy2gJZZayj0EHYs8jQI4Bn/oR9nY8tYgnajW3KTLox/w8/SytjMozEV8lUMptCEn+fz+8rf
36UCBVstYZACv081Z0CDMndMnV764No3w2MX9v744UZxn3H1knKbTIhzLdxk0SuAcoC1UFJTdNG/
Tcskkt0R5JloSacVEZ3jj82rrqeC9EGF9e7Q/TppPqMBCrBl+M4u7MHfWb+oOIHKnxzytGcuWKxK
KSFJbdj/PLVVP4h1HoyqIsUl1wZJx8SkxLVel8aOJ17s8VwtmWBQjBMcwD6lUdiLwIQJfVfhxflx
WTWgV4YogOTgK52c0OVGEMQ0Bez3JuROeEhizKKD222G8v2MJZz+hNQ+OjU9Jm/16Osi+uejGNuz
DqaAhaWVUmIlnPI/iTEcCDika/Taz9/GWSRywKhRi1O98kWZIqtv6ntu/O4kopZLd+Ai3EWQlqH0
Y9gqgdCZyQO+KYvKikET1W6m9oRqHHj0BHq3ErovAr0XcnBwnEd3sF87TJWpxXnKLrJLfICZ1m5N
T8Mb45o90RGaj/m/y5yp6h7SRv/6r/NWPEhU8v8f8zwFEAzBDqrsU1mahBn4TTImdLzXi+pkKJs0
fy4QvaJaolA4IhwPn5IoJLuVlHHzhI37vtvbElp6nkVQB+5gp+meyPVYTVr2fCNRRR+1wRzPztqp
XWwcERnIQeUmjT89dleV3gfH6g49R+5mch2Je2l0WzCIIHmfzYLuZe0cpRIZAxFyvGZ/oI/MDSsC
cyukvNTFszve5Wg5r0hyXv1AhzCn8zai9QhHfFcmqTIib89JSvjSL04gij2sLLpuV5JJ3MJNNBSj
a+snAJFMbio8Z+gG1pu7VFZbkxEOZWFGvPO15na9/9HIMT7+H2HelT8jC28DXdwnuiYsN6bQXpR1
yT5g/9os06OoYcZvO9wFIoGOYBl8kt9ugGvdvwJowBpVBVfwvKqSNTZa7wLCC1xK79IHZbisQ1tM
TzPBJRcTaVg23v2w3Sbc4OY1dY4cfwooIkgsNwLkmL4EIVVlytiFTavI+/2dN3HXt/BmhynVQEXx
Nkk8QGHSAnHnJAW2ysFI4PFKqk8AdCUEun/zOt0+CzDGuq2PIzXM0ORo1PnsOa5Ilv3GSwsKlpOK
OdOfZ3MmCKj56KKPuFB2DYZu6rFXW4GzuVQXffYLoAvEi76NFJwjZZNjLiNFnIwG1CLDCNuneHqJ
oZZJNXIIATWEWIKAl5JAQRYd9EO6GF1JanJcLh3311LB4rnCx+OOsksV0pePQqEkcC9HO7DM4Rbk
8Qn5EbmxwoorGaCzdr5P+numlKG7Ruurr/rO4ZNdOslsAEiy7mitw5z9oeyd8gu3gqw+3VN0CVrh
M8XVGDBesKzwJJE7AgRrWtLUu1luPov3jAT0WVGj5iGOdNFlM9LGFbQ4rZNfbVtYAuZimNnlaffd
cBaq0i9GxhknhNVgigDm6Y0eNuZppQG090WE+sn0/+5hoWMdQ6h90aesJ0UlzQSfrV5Xh+X9HXBC
2Rs7mXuBGUtRYX6hLfwwghN2Qw+Nz0UhFhWPaYqJBVj1+QZJNKCn4JmT1eb6nLcgil8f5Rnb6SGO
iBn7V1urw+oOKAiYU+WK9jZ/o05Bfyt9q/Sk/gDS95K3DQ9WdawgQ1xxPx7qItdR9BzNKUHoYoBn
zcG1c8uhhLTn+lcAoBx+/ggDjs48MUF+ybsFSyIvNOa28GHZomBnN/BvOITqfF0N3TaVm4/ItTVd
Zrynw65nfBLdmsCr51R1xFCL9yFhU4w4eNGUeyrDd6Xs2XPqhALVBnO6uMnhuTTIjUZVGcrdLY7g
iElC7afH6710f6QosbZlni/QgS1wpswuenUk0QNl+FIJFwune1vJ+ZZ9VMMFMJ5sUF79GSmrS2Cz
1fn1PRWNmK8H+8CLJ9zSxi2rkd7HtYVkql7YdedOst5dIjIc/1CC+whiZ+XwTSOCR9yvhIj99bsO
ZjXizDwCZ04Qa2Es1n8Gp/Dfmfe7yKk3FAXwbXgGhF8yPcjpTe/r2UNlcHcyTGkSMKFWaqybI/9v
OvBwR8KyEY0ihQkS0Cn5ohChfYdeWcGKQ9E9g5Hw7wo3+ZFXJ5h2Bwd3I0l8LUc2scldholwt4gH
mgp9ZBvXO8OUFL6eJ8gVSgIlNEQfxC4G9p5S2RLNQ1tj8eQKdn5MfSNnIIgXWFJ1MpAjXgHuHUmh
/kJSwZC1roIWofA0HDPpNRJ88UeSeEPRlIjHZqJxuhkSKQyI9oP3JnIeVMj9P/b96A2rg65aSAyi
VYaB1Q4jjlpKrPGkhs3TrJ8ZGxjGQ+VevbYK/WGPmnQs3ZMtYcZzgb+oK9XP+szzfYQCtRi1r2eW
9P8VFvfBNzs4Pus/9xC2xLx01XpEArRzXUu2BBDbTGovNJy1Jr9gbm5a731bl6O7BSnTP1hiEBmf
JN+z4nkEgyO0jFLI2CZ1io4mI0WA0uJS9DwRpbR4lPzS3A4PaQpQr/M+FgYlIhLo8kNqQod5oNFC
c1c2vLOxrSd8fBO1dv45jCTr0BOj+uhwtgD1BkdK+TIwaX1fKaFObE5bTLjPA0gNOUD7WtIzy2CS
kOd1ZiVx+3qBN6XXL0RrVwFvUvsOlkZ6gW53AJrGXXXVEjWCnj5P/FTFORUUZZKUefaa7iLKLLjV
65hJd//PbiAPRL1keKhAkQPMllm7JAu8I+fcHjsMv3HWiy0ToFM1+FZgF7dmBDwiRNLd4opkU/Zu
W4oGhLHFF9BvzPeGc9ks+mazlxEztgyH47q/17gJZL7j9nvk8QOBroX7hQe6icrkSCRf4YzMS5lF
YmpHKSTlE973Xttp4GnK6U75qk5M1B4Gj3Zu/o6tTc4O42Nzs926o7qOUsHCEsIn+btXV/c5iiq/
RGPYgga3MB4sFBGXzZCWol5tEkVLzpHvBdWhi3IXHoaT0QRH/SAk8J4aCelSDsaTXcSS0wlDtr7Z
okJaY8G/DUCKVNPlSKLyHqtnalZJLBO2uheIl7lRUqa3CLigUf1znXnWX5xiB+As2DnlZMvNtKAJ
G4aAzx8hc+Yrw+RJy7ZP8cC8LcKLE7Eki8mMV2dmE/Bjuni8CpkK8rH0pFL4DgxG5CLziN1/9utJ
9MeTUOLfuPXZKNWiUmgJ4/DH6nhR7BCCiShoEEzh6lak9zKF8m3NIXRH//4ncIHQZDBS9hEWTBqr
rYosH3IdsoVF5BDPZD4k8AKBRyGk+xrNWGPWG7lNYCBAgZAW7U7MmxAv0TnOAnMfefPujfRWVZQ7
FY6zAlLuDdxCrdsAn6ARs7iyFac8NZae76Ef4c1hcTotQppYw+Vz7gQu587ejm69WtzAuoujUPer
QTnSI4msKYkPc3Lvjh1AHmM2z25j2QldCSC7Z6s6vnEE0gqCrm6IEdSIyF5Ob5jLwG/PSzdA1z5m
4Y8zNveUgovCyIcX4P5/ZmbHZI7+3uG+8EwMHu9dCMzvWyxw39gEQnKjKzwgW86DdGUUodzfJHWi
7mCpqVgpjDDvv4jhyyk9mdnQrlPKiFSgxNfjWPZyYbX3Oct59IY6y2EVhm7pWA1ql9XC+VRTwPfV
VLX3HF9jOqseWBmg5vpfs8e199n5Jwd/QGPqip8y4VhThCfY0MTeUt8wWGv2lR7SUwDVkzIBzHT6
Isnfzg1VMQcmFCYuWcJZcIQ3xZ41zeRa2S2LUlYImbarVFBloIq2CR0iwmCf6e67x4zB7QGtwen7
oQvmPd+1X56W7tQSUD/Kw/YovhUwv7QAuFynchriDllNEIiDn2Kj548r9XbBS/imwBwnPajkKFqz
oL/evFjgFK8JLE51rj2g+htInLim/Q3G030GlPTxI6sZWKexc2aDoz933qfQlfHD+njvMZ4bqn49
h0RpZSwWJe4xu5E49zOg6kv+YYaIlFAH+E9S3kVtA+3QhdvFeWgNwu2t3n/ZYNfSC6DzA9qxV2VX
Jy16bYTxaJSQjOIqV7HL3+t7X74xhi5ogWvooZGslNajROiv3XHcA/8XERLMFNXP6MhFNARqoHcd
hAW6CmEOGPFsXkvco0/h8pTF+skXvE8OxiBGEee9CEFJN05ot8Wa5TUrXnZRDPhpLPa8HZQi9E1h
Ai0W6pzDx2reqxhn/JdIlTNPQuACGFtJcXFb6NNpvIe0QB7l87dIFcU8lanSMNsQszxuYXFVyw5F
/UQUvrJLezI4cMUjn6baXcYSeCM2g3H6R//Pe8q4q2u7b+2Ej2OhYIK+natxNIUPuYXblxLthKyq
BpcLzyfDOmH9xa6k0pjqEJ/fNAqs8Iv3X7Zos4PVK2++HoqAq2i0LAixV8elrGx4n6MPtPsD7WuW
YwNGeiK4nP2ljwawuK36RiL1B8yXkywPmhrqRcQaUg70GQXZBMyre7yxm5/Fb2XcweaRF6kNu1pa
BHA262wkWtXyvldFnw15jO3r8UEyXQde1iixN4FEF+HwO6Kqp+oMUwsJjTU/zuFl3OAI12YVUDYu
rTIMWdxFqg3X2Jpgmff0UYFtg3+Qo5eZndh462HX2iBVavguVjePp7Q9IizF7EezdorK36N0NQGY
WCL4s/8utpK1wCZEE8FL44uNal9qLJTBbhP3e3whGHKxkvVvbD415JxmqW1J7U1LrKUxjgpssmsi
FEKzp1sEHnjTOFjCCkhurKQDJ5bJYBcna2OP/OkzfW1WZC9eenvepcMvZZ5paqrB6HlgrBA5YuI+
YKdzsvLcHbvkz6mn8DRgvD4+8L/mNSaURnYEPIr8xZB5fhiGdZB1JKPhcoSxujIaQUWJAS3NVF3p
58rjL5GSXnHHp2KZulWJeu+JD0W/exvSRf+11lqpqntpvr9MnMBt6iG5z/GwjLCu4K+GpQQzhJe0
919umbHM+2t8zJZOQDawpQUxJyXF6hTV+E2udf3V3HElpI4YbxjEpfVUwsITeqvhevxVw35jCQa4
04G16Qxv3kRGP3+i4bzSB6L11NlnaRyATvKMrBjog7u5YUA+mWaoLZt/pwbigNVlzTqTQG3TgVh5
TtYhc2v7Sxi0vCZ+XdeffEYmUdBvhlvLJ8ihl1kRCPF3FnvW9v4ZsAyFhe4XlfrMDfyU7ibvthPv
udi72RCBkQ49HyID/0oxcQ3+bOdlkRHlNmDvFqg2oo4QlD4XZiswcnsDQpMrZdW7x+lmmz7SPKGi
gV6A0tsWDR149iBiJRdmPezbfZRjYsQBpHJiBvhGuX3eXl2Bu59BtQ5nIMgb69viv21/VajRlXJa
dIl6IC3hlnSi8eVTSbkf5rA9yqOuKpxCKCXuujHTAcYw1RI8sBVXKYZ3K0rm/eUWNzZojNsd0R1h
iLAK61twpCP5DV1GSeZoG71OPBRWyNYD+wvxZEKiACM78CUpyV8ODyDX3qxnU/VhFXIbUScrh81j
b3Ack4TbN1jXz3KDkDYP6v3vrwAd4y3WoDasK8PQMDmguH+Z9BRflm+Ltx7zjinH82S6yb8c4G5N
xIH72DwnqlhWUo0NLdl6SzdfUOzKqpiDDe3gjCqBQaDypiwoUSbBffoTMkePZUYNQm0sJBRZG5K5
NCbKN3ZuUZRpd3VM2qBiyhh+ra3z1C/NcDBLhqJAtWFLX9wbkHXpJojCYr6i/MKieSIC9HHb94Yi
BEOXgCz0KigeU4vLK3ypSnMXTqW4y6+M+ve8FLG1UZxoVMioml7eViLvdAOJHBaorWC6cXYQMcOr
1XbRmxRLT1/LtSe9G3/gZ078+syHsAJBU724UT1jNv35z2TFp4VuVuvnA/t8VzApCVwWvVWCynNQ
ivSdvNHw7B5y8w1phbbjjXTJ3F0jI9lTq4wJu+gp1Vg7uRI1n0zQSiQAlWA51C0AgD5Yh42pfDlE
GagtQ6D5cDfandaEcey5Q5lJ820gaiVziIPV2QEU9Ro6VApfxwNFPmpXnDc9A7mArBqe5K4Fxuy/
XzACVfoAJJDxPd4o4jOqoVmeRvFAn/8o2NVf1jb9/NjJpx/wcDSdlu4JxGpdRxwGmU8NT+sUmBBK
aU8FaGbWLXFPSXtZav/gw0sSDOUQnFpn2JfXq3Az8jQPKtFsjjA6aUBi3iiTPPGdlZ0ICzC3YGeQ
rkHSsZqbvbdl49mVKftHIVE5gHmk+IqZgBhSPnLhA8sVjHOR/1eVxnYXZ7c+GShZRRIvlKNXmk3p
vKqtaaXkMZ2iYIEtlPRfVaPE1siHcrNRO3fx/tzRr7byt3El/2bO5v15kHwMcqF6v6Rc/OxTX+Hm
OCT06+rTWlEZfKtrjqoz6uZpA2v2mqNqOhFzwizpMEa4eL+pNYUwA27MkOWJeo3gTy0HBZuqRMbp
hrd+oNdUdzRJxFpsesiSmZCTZDYyMSF2wbA64HUstykwold18p9VsrrHUYKPVW7deNlLyZtGL6Qr
xKdgL+9PyjExSk7t8L/JoOJX+MDaD1ryNHnb0UeJKMZd2AuLZmGZKcEiZGJ3PU/A+SWfhAgoqpbw
5lgZ9knnc5+JtW6/B5fORndJWWfXnl0eVcYf9CF1WL3M7T6Jaxxrmj8TnHeyVAu1xF/iizwlWxuR
xsSIMaHiA3hjjwi0VtFT++7wV0jk7tYnV3+PenNb6Hxl+qoxOeqm0DRoKWX+u+RWJJ0rzGiiFZsn
nQDFckysgO1JUZGqgm7mkzHFtsX7BW0NI/VkavN4fEDzqCUQ7J4FJ5lpOSef5xIr5J4nLtpQ8kRc
wswTxbomJ2cNV3D59+BWdJ7LmOLINliAqHHMiLFoViyKZAIoI+DTTDTUYMeeTNfOoffg256q1mkZ
mOlXBH4jQsBBaEQ1xfVvogukBlxJBwezmpSB6XJ8oTh3oRh9zvA5STJvSzIAWOIi3fbR6hoONEjS
fH+5eZCdUoEZzu4FePcTr+4k4SX3Q9bzCycaEzP9s3jYVJCiQQzPofWY1JWomgGr+xv/16JjuJPE
fG2Nn41/fdWsk6lN04EqSNoluTcwbZ9+3zubQo5o43OswMM0r3nozAubGfpdvjBOo5bODaltIXVH
8hlIwl0GzL28v81WcVlENe6orwhG8FfRvj6zxb8i8UGjrKZcNF2KC9igHEAUlkqmPJ+CaZeanWrG
RQVrnxba+TWaZlcz6xzWhwbbalwRSpNsmilNYvZoZZG8ugJLA9tTBMh+wiERgmC9vWOewoW3ooYe
hNg38oj8e8Fo48kJkY9VT7NuqzWXrqGce8iYVPcbeBW3/IqnL9stxrNMeBLJRRvyBno41kl+C6mC
w3PlVxvzaN0V+c3u6yUiQXDt5rpDTD+OeSTaAtzE0TEVg5nBw/1nOKgarkZpyejdqmxpAh7x/Y1+
EXsZhHatf2n1rOOBGWRt3IOP88PyWrziddz/qr+8eJ3/zCvDV5eC7YfjaAxmpYpyAO+W66TvFQCz
Laj9b3j4ZHBXN7/pvjR2/SX0VX5G8x/dyLc/ZNklhcL371jnm3zqWk9vE0es2q7Lu66qBRdep2Xs
BM57/qubGteWXMblMirZL+JSfMAiYKqE004tHIfI2SB6hTYV36g3h0Jzdghcguhd+k8A/ixUD9ot
/JXDaXLFfkD/4+q0mFlfx8QEX2UG7dIBBazIpN8Q2NDJgz7ZMdx0k5fykXyjNbRzFeOkIVv2Jj03
fXkqD6GOaX2+OWTgXb+ptyVAnqkNlAjJcEXKS2E7V2ieMT8v+hXd2F2h7JbFz5f69AFDVo7Elz5p
hBJZzS/Lcc8v5UF9TDHYv4dcAtIvesG8pLB9OSixArrtq6WB/k5GK0ghmRW76GaLHyEAlzbO5pF4
1+zXGpzMWHPon0QgqDoEdx+z9E5pdaLV79EUih28Gcu10fK4EMY8GI3W/WnenWkqTpDJ3AI7k0zy
33KKZ0nsf/D+/zh80ciYuVaYzg4xUF//CZcregaDd7on+yPdN6XDbTCCuuvClG4VtlhTtjybjZvk
AvoiKdSOIdcJvT5iotUcnzUEhaBNZF6fHYCq4ltK6ObQe7XiATRSzewcAKV4QN0HCAtvr/pf/8uw
0t29yeRJRT55jT6wLtcLRvvg3vztggU7OVuOW0whgU0YcyMLHFy3hVEN+VqczKCUKVgQ6ZXHJj0b
MLPaqVHrC4GOY5htfZfMsOXbr3YrZH8ZqKqik0AWR6UU3BoK6qcxfn8O4l+WGU5ePTWhSNo3378Y
9yOaoNGLNNMYqysSzUIxrYyrb5vSXrjnTRNsQNbZcYTpEBvgous2wVUNh9hYp0MqB1uKf4I0MvXH
DhnLf2wRXH/LoAbBkvQOJ3MkBcqfpGfBqt8jHqx6yPPi/Hg/6DHzcBdQqJcCLUCiEp+69ED6oZcQ
waOw2mO5I+6W7yemORQxfNyzHg7cA6VzIqxdfcwfQHaIjmuEuhdiAWVmmPcpWjcCLi6WkmFPghdF
rClPUQguyfKVIcjVLqRhUYiP84xCNyZdXNoYQEENXZrX+bHMu/udBJPUjihpAeZNGx4EAYuPAFoI
iCzoZJdWkebgnjaZUvZ75iLnrC4k6ooXGl1uSLiUfmoXn/PKFWPDY9IUAdce/Hvcpp4bS7UrvKVg
hTAWDjieGlYYHryfZZbA6SEblsk/Wp4q2PlB4WZxgx9SbMVRLeuZjq8LZxTS4cLUql5LFcj5e/oH
5rs2b/KHUDjo6SzeU/mzfckbwQzyEwHAsYB0ETw3Yg+0eLGXMHssUCrarwmjFD7D97o06HW1tlRq
/tVRaW98l6om+g25jA0T+cl6bcB4A+EPsChhHhIkPBAV3Ld4HvmTBdebsaylltFVzqtHHC6qM460
nthpcT0Hh5432LAT+bK8qbDMGndvmG6WhWe1QQlDyUk=
`protect end_protected
