XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� ����כ��Ĺȵʣ�)Ue�;tS��[�.�d �$�2{���l
<.tF"�EO�.�B�G�ڨ�)J�#p$��퉣ZQ�w}���������c���K!߼YwV4�r��_��+���Lʢ�w����bezf��ƒ���5<���s�y�>h�c+wtK��oyA��~.:sX����!3�ɲ�Fe�
��a3�!	��L`Ȉp����Q�����'koѵ�'sִ���(��d�8���2�U:&�v��	�c�f�ȯ�;�@�F�&�wz /bU�*�R�����ZrQi���R}6�Tq��f���?��7�f�&���f�l@��N��a���>��B���,4:v��"+��OH���D���I�W�=4k�'Ͼ'��n~ǀ���*v�6PDAh�@:�K��WϾvT���A��
����4�z��}�5 2��Sp��?3&'A�fTȮ���m�}����h����cJ ��F�Z�~��X����f5�SyU
c�q�a@)��a�������љ���x� �S���|T O�v���UJ[f�M��q.%5��I��ٲ���WJ�w�h�7X�!�Yt��+yW�5�zFt���!� ���ͻuϽ�ԩWE����& vgx���? ə����_4�@]����/l�����ӻ�(�0����G𕝿�{T�-v�=[9o9��T>��ΤU'J�8JA�3K"�2�'��씗U9pLg��G�kw�I
��o�=���ӂ{XlxVHYEB     400     190#گQɤ�$pk�1�	��?(�/�HE�4툁��b+�璱(8�˯:j����^:�'�e��1�?%U)�a�%9�|Z?*��{�q笉N��|}�4���A�E�Z���S����k�C���z��%\h%�|���0��oY�����zէ�e9��<�`��.�}��<:i}�Q��ǰp7���^�%�͹�c���ґJ@�'��J���������C�T��t$�u�yֳ�-DP=,���n�e���©$Lɽ��iW��Y���,���vу�4�����JV�] ��K�cGp,7�H;-�{Jb����h�$>c�/��{�r��)q{i�<��P#� Nm��6�-��Jѡ̬m������:wm*��X�.^�)XlxVHYEB     400     140T��?�wg%|�JK����R�by��}�v����*Hjwy`kT�e��������M�nl�7�t��	x��P[^
����yӅ����3Sm��|
�ja��F<G)�5^����[>�(s��	�ߍd�.v�=*���)2f�U��$�>�ou�c��d�ų���'\���[�p�ԈĿ�O=T�[DS-��f�\M~Bg�G�����刕��l�~���m�y��	1��vV�Go��3�1:��*��qql#�sxHuW`��=�� �ꄺ/)��c�z"�o�<�x�� ���h��'�Z�XlxVHYEB     400     170���� 3�U0�z������>����X��i?������?nsC���4��X{��l���N
�́��҃(H���Cp�IpCd����o؈�TeoasgĊb��Z�h��� ��U�uc��qm�z��� �P�~m�WЃ[0�;Y �V�_?�Q)�ߐ�+��D��Y��@?��!�0�T*{�o7�ݍ?�=\W�08�	�XVA�Hz�Q��H'؆��H��;:V�E�2��g,xrD��й����?��Q&�|!����B��׹�d�$" 1*"�m�Osz�<�Cdv�?��=���zn4C�Q=�Ǌl�c���|E��Я@���K�~O��i�ĳbh�/Y��XlxVHYEB     400     130I	�2��օ��S���M����}"�����ڛ��-�&��� ��-t��Y�+�v&�5)�Z�����U̞�J�~u�&���'�P$��0<7�U[�E�׸6Te��1P]�f�m����o�8o���X.����Ki���:j���xϜ�f���TʳM�J�b��#�wn�������ꑓl~@�'�p���a	���Iε�?~ߙe~��e�1eXl(ݻ�<��!����jPcȇ}ga�b`�����U�v�GB�b����c���K��$X�[�~���r��pA��@!���*�TV�H�%��XlxVHYEB     400      d0qY?~�_:%�{åx"m�se"�Ct��u����@�M�����_ė�QU$��dM���v!~R���t��h���Tx-����߇a�K�% o3���c�I�X�aInC����t���Er�:�u�8v�	��i������Q�+�_��:��Ђ����_Ɗ���3}N�P�G7w�z��]�'8U��'7[����L4Pف��v���ƉXlxVHYEB     400     130V��&����)+�OMIz���NPr��#�3�h���e&wt��ӛ\m�K�7��7A-�Gڍ��xdc@'�� oqi����|����\���Q%�����,x5�Y����/�,���+�T������)�i6�͇ݩx\+|��ѵ�9���lS���s�5���5�p�R�L�*�4?����L�P�"9'UEy�Y�o��T'�3��M]ln��{��s�uB8{T�D�*���*)��mI/ۨS��`�\������"�E ��>Ty	�Mۨ���9&_�?X	K�*���m�XlxVHYEB     400      e0U�\d[���k}s�=M2��[�g}�t��)�#�����0Y�G�xM��4�n]H@(%�tϷV�%.��<Ǿ9�JHE��g�@��ܞ�����@
�g���rPs7ZI�Z!��23Qi5_1PF�}�S�U(�8���80~muM�(47@��~�a2�bH�J�T�Ӧ�gx509��2I\vV��_��,U>�6�O�1�b����s�6��M�ad��0Nu)y�������=XlxVHYEB     400     140J*9� �5���	��nq-�&���b2O3�Ԡ@}/R��|ͫ}�0�����u�G�4rv�_�Wn�%U w0F'/�N�d]&X��%"X��S��S�<ܞ%�>�<*dS�Ժ{���!R�㉝RZK��B4՟F'�*��iy���rz�J�'����EW�:�gJl�[���(d��)���f�{��fm�<D�粲Y�c?a�������[�{�x��H,;��+�G��]�jzǀ�<�Bg�o��dh�3	���Vo���;}wU:�E^鉾V�"d����8�e��t%�s@���F:FU��VJ�ڧ�Pfi%���XlxVHYEB     400     180�4����V�tAT�}uҼ��~� �}wzt��S��|��M���Ṋȃ���<��#��P��[��b��"�O\@��� vs�]�w�hW�.LkS�)�(�
(k3�T׀�7d�W������l���V��c'�f?z3����J �����"��[q�F�9ZK�\����L���]�o2�gm��L���"���2��m`�}��`�)�E���鰐�ϭ:�����c{��w�߲ޗ�t�e�z��	���Q%����}H�v��>�JJ�Id�L���^cB��OI�@�@��U*�ö���D��$�u��-�So��;�h^�{�b�,EX�O���2DS���+�%}`��)����d�-������XlxVHYEB     400     150s$���QΧIn�{ %��z�S�'ζ\�k��F�TAi4�`.�46��5Tg^�) ��(gݻ�|poj���d���%zΥ|���H�m\ ��9z
%.|�J���\�H��(A1�QK�"����Ș�;i��	y@�!I�����=�8Tv�kk\L�wi�nr��lM�j�i���.��~`����{�Y�F��{x�	@B��Ԥ��E�M�]���{�P�$]�y���Jm��*���a��R��g)��;d��`�1����.��6�QC�P�^ |�ϗ]���$	�C�m�Bf��ь����_��[r0�lV�Zm��]c�|YU&t�ڒ,�.S���XlxVHYEB     400     160��S�0�F�YW�ࡺp�-ZN�-�k��W��yQ����>Gi�!�Sw��b�����<��6��1\�=��'�)����w	�Y0�H�9��I�Pvt�9z݉yܳM�5E�"L��B,���B�2��;�}��ڥ�b���f����l����N��@@N\��曑,
�:].Ǌ�Iob¬��&C�!��q(���v%*��R0�����hX4���%S�T�U>nb�S�pB>8�w&W�snK	&c�I#-.	�(E6̪b�\�ݙmp:�3hVg�����9c�8����8�'��?����z%N��P9s���&q�4fw?�[9*u\�f�������H��O��XlxVHYEB     400     130���/AJ����&�Ō��o�m�������Y�f�t0HN\,<4m�iʂXO���������F]f�����"kXcU!���v�������H��=# [uߗ}�ک���w$�P�{n~v���X�5��K��JG`a��[�<����~��N])�,�&�٭	:���&����e�^�v��H��.�2>ُ��o��u˫���4�"�l��n�~���gn���l[��U+�o5z���)y55�x�s=�<z'@��%�X�3���P}�$���Đ
5d��A��o;�U�T\{XlxVHYEB     400     140�V��~���~]9�b>����E�C��pӆ��1����t��O�,)J��V���V�{����#[uBa\�BF��u�n���k�H3N�� ���-��B)W�3��-�Uq�O!�=J�"j����i����^�E%��p9]�0"b�+�I?�~�moE�����];��:C�>ױ)�e�yV�Ry�#D=������	����K�m�k����|����3�^���mD��>M�*G�	]��1cA*S����F�]D�-\�岋R:�W�X':�jKZ����n�@rUJ���+���I,dQlᐱ[�XlxVHYEB     400     1a0��M�{����)����|*�N����^U'����3:�A�V5��B�"���%��9rZ��P���4g�c�\D�{���L���Os���W��ٶI9m�H�zui[�P��3��n�b� ��Ӥ��*���� ⵏQ�e z6��Xth���/{�u�Gg]ڣ�v����ظ��IL���̆�e�6����MΣ_Lgn<d����8�������J�C���%ڜ�8����SZ)S����M�����/6��В%���X҄���c�d�������|{o�y���Ď�*�_�9;]�6.@V��5jm�{�ZC�б�"�=��U*�|�1�䖡$�&�j��0;���C䏾0�NN��j���Fp��(5��@�2�}�y�_�}��S�O�ŀ����~�V�@��Ӭ�XlxVHYEB     400     120���б; �e�ɘ�
(�<�K1�-��!K2�����))��8	0�x˺��2y�U�BG�A�����D��bpƤ�G�u�0��䙖[ha��2¡)��2�9ЪaW(>�l2+�A��9X?�-�V�6����8������u�f�4;��31���$�G9c�FM�fC�Im�}��G!��ąc٩���w�(�<�7�|l�3|� �Y�X��FH�x-d��ж�ְͩ�qa	K$t�o�����e���CB�2�ܴ8"2Y�P{dO�TvMR��XlxVHYEB     400     180�ӻ�^e����VK�<Ȅ����گ��͗��	�3˗+�Z�!���fˡ��=� t;��z���Z��	$��GŬ��p_�$k���yJ���ú�L�S������=*	����,HgLt�A���H�k�x�PG���u˽�E.K->/�}�(n �P!��y�8�|t+��N�^[�%j�k9W\�)�[��fd}h�'�K}��ݭ�b���O�N����'�c2������	�n����ە@`f��y�z2���f i�7�1޻^�-}I����D,{'z�zν9F��1���Iܞ�C���/'=�����&N�c�*������<s��H�tL�G�C ��g��+toXl �hi�}?�(�,��o[iLv��^��8+�@OXlxVHYEB     400     160��1 ��ޕ�S��,u�o���)�9;�[*���Mx�>�m�hCY8���&Ds���\����xQ[����{��=1c@3�����2���f�ٗ�$n@��Ɯ�'D��Y]��c��`V�,{�A����Ue���������zpZ.M���섭��K>�Z��Ӝz9��/��p�!k�Nc,����8'說�n��g	��#��B;p0�@e!Y�{J��K��B�u��sQ����܂�]dP9�(U�����hĢR�f���v��1�A��~�w4��|�k�[�O0�'$})�z8�
gH}ƭ������(�d�����hS���XP)���fC�nʘf�XlxVHYEB     400     1c0P|��C��xk�%����nn��\�w$1M?���kQ�(�)��J��z�8p��U ��������0��������F�yO-��h��@��а����
�0�f�Sy�Vަ0?�@�g{�Hj�/����Pd�7��u���l���54*���+���Bn\�����p�A	:�"��<�%���Mp�$�n�%(ĺ��4��ى��m�U���[^���V ]0�enJ�.�f�Z��~�آk�Bs�Z�X	ܐ_�:ٷ�'W:}��^���7�!�μ�N؜����u>���	�E��N������,r�����-r*j��#c���[�`)>�A6�5�}� �r{����3*Lq�E�4Y�_Dz>E�����2�^�l��όׁK>	�#�v\	�vޤ[��Q��(���Ѩ���<�0�~n�1����|`�3-XlxVHYEB     400     160NDA?���pH'm�Pp{���m�$�V��ĤM����<�*��a@�ME-�HZ���;iH(�C�8c�̽�{��Lt�2� ����ܭ��<0�H����K��u(�K`����1�'�z����Ǐ�@٩��Ȗ/�87�%}H�-��B}ӎʠp���2�_�w��d���1��C(�D���l��ElI����G�-�~�8�LM_XJ��m77-z4@8��\c���V��,��j�2#7ĸ��s����~�$""/4}�0<*}�2cz��

�����ͣS,Y6���u���??�bv�ewl�~�����%�a��jխ9�+��Ov���u&Ѷ�ӝ�ٵ�b�XlxVHYEB     400     130t�l�2�+}��
�'����#U�0�oT�<<��N�<Y"B�q�8���#R�:[(�9&��!r������664'���1.њքrP,�TX����A
�eцs3a��4?�(vr��V�"]�-�+�����J�_af �[Ա�󘣷���P��6(	�d!�ANfz��DĪ!�ѝ04J՗`U�x�r���{���>�Q�rݕ� �R�Y�1��
8"�ı���M�'*~����|>�[:��۪��i3�J�SˑXR�3�wtea�u�$��I�$g	ܛCD��G�x�'��٩���r{!)�\XlxVHYEB     400     130%,� �'Љ_+	�ѱ��;��k|J�U$l�WW�*\\����p=�;
�5:Ib�jMטx���9 �$QfW;c���p�Zs�^9�_�ӌ�ҘN�7z�K�6�ҙ�;���A��Ҵ���vך�'�2lu�5��uZ.Y�5D���1�C4#�IN+�,��7l���r�  �F�:�E�Z��%�ѩ�Ǎ�ńC�R��X�)�p�ό�������5�[Լ�It%-ƈ�������F�@L��eF��T�.�8"��S�ďcW�C�u�]¾�VD�l�՞��C_[����XlxVHYEB     400     130/&�t�D#ʂ鳶<]�k���R����E� �0��g���|1����!�X��+A��^���[��sF�>�`�����¤v:̙��;���K�PUܾ~Yg���UW&ݶ�A]�>�ƛ8_!B/DZ���l�Z��8br�m���fY���0Dwf���|&�;���<�������&Fj�+d�&���A.�S��YP:�u\���Q]�	:�6���p�13'����|��"�	v��bc��U���s;��<��Y���8W5Y�]��NO��Q/wo=Om���k/k������ Hv�d�m,XlxVHYEB     400     140ʉ$������!K[tN��l�M�I�=n�i�B�s�����z��@�L�W�5�%lI��C�f��Ǟ�j�.��ӈM�v)"+�7p+5x�-&�y$�JBI)��g��i�Zj��*A�~�f��g��Zj_Up�X�f+��ֽO����&FQ��6�� �J�WR�X�|q��+�/��W9���Lɕ[BVg��O��Z<L!�@� ���]��B'@x򥝒���@��`�41 JN�S����_n�7�Au�K�/���f��d�\�
:��7��|sB��S,�hP�NM(�a2|��XlxVHYEB     400      d0�`���Ԅ���kG�ߞ*T�*�ћ^e2'��̢W�V4í�����h+�?b���7֛Z44b��s�:�w0k�?u6y4b��#��le�����w0+� ��kkV_ߖ��Y|�@��]���nÛ��g�6�M(�H�^��k������T����i��pٕ��M�����[Q�y�L���-��@3���t܁ �b4\�|�;�XlxVHYEB     248      b0��C�*uyj�����;P��t�ߋ^#���*���{ɲK�N��;F�[�i<7���K���I�}�$Tz�6����_�f��ڄ�(�"�ۡ��d�'�f%qH��L1P���8q�����L'ͳ|�f���L��ߎ���v�o�:SP���=��G>�L��K;є��>Ml徝@�џ