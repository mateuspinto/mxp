`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
Llq2J3rE42EUEzTcq4/+rnEyFFPjWF7m7EYAIIam/K0j7Z16l0T0b8ct//w08G9GK6yUQPRqi7Jw
ljQWnlHh8Wimix8aypX7llhhz8qcOESdDZ2EdFBeOMtjVvuWjBu+OcWoza8YjUjHcvVKw67ckGfO
7ExbGLw+Vlhi1jrky5DBi/eaJxSGa9y2aAzzNY7HGQRissFmx4W4nNOk24u3xzenS1C0ds+V281P
IqG16NC+heUORCdfrQmZiFtHGUEOGe1vQGch5Lcj4GNPk+QmcDuX9o32PqZxQMexC6VibYjIep2A
kIrAYqPep6+VIkBJAS3PWcTQhGrRZo0nAiD+Gg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="H5qbLAXL0eykz3OXO2m68PVgMNHn4TSQlGFEvWQxoaU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9328)
`protect data_block
x36qdRySHGJs82j47UpX0ietJd90mYJVoetH64N0wPCZyTEWm8DE66cE4tg9xWAJWtxmJd3R0HoX
YOk/5jR7VpF7S4TMRDHvZs9e4WYJpecwFdmTgLwQXTKZbA7kq279eF5B4DZrHOx2G4MS/0D8jezv
QY5G0F+jqHM4w0xooKBDqXZINrU/I4yrPVElKf/v5OJiydDRM71Qm46QDRXVqtSdU1rvZrknhJHl
P+104B6qTfItIUomDDX2zlS1XihH0me2kuF/Bj+c6ibCCs5NfrttILHtkA7QWS2HBKYoSlNW9v2Q
lK91DjybtU60bBuTnCYYHFiBjjaS57+r14SdLv2/3iEbu1gDtym3xwNHMj8OuwnutjDW+T81cCQM
cLPviIonqfn5rMRfDl6ANPuyTr/6qxLuglI5d0C1RQbAFkqLmNouKqp1K2N9MjodknbICRcT8Aa4
tie/IiSdWfbrWtQY6FTAY5nnahYLIRDXHaf4Qoqe7MteoGXWFbVYuJwuvfcxfwEDc48uJVqkTeSd
HAiS7ttevgIFYwtZFdQ3IQxBB6kf8SpH81M1/rs9kZB6cLgHlhNoK4+FMlCR25XxG5mYTs7EVkQm
vCsFPu4X5w0k/WeUO5FhV5gtpXq8api/t0uxviU5VOA/YNkgXxr/CwBc3zEU86DNtsIdVIfTXGnT
zuq7zZkAUX1/YAE8wj9W9it42LgUfH3vcEvUdL7oog5iVDR6fmATlyX0s0TFBYNMPAeqQA/yap/2
aSbeHChTQtDquDtJy4wYPCDiJPW5aelwiSxz2qgG1nk/72Pu0v+TQ0XgjBvutDBNC51QcX4U1tbE
KDp7mPZeElEP6gdKqUjqEaqyeyVWNTMIibi7k/3i20qxPNM/XtqVeOnQdoLNjazGSi33KPnExFYJ
R8kwun732cc0osgY1hl+PRqjZXOQVxXXrYKUxv9enDw+JtgDC76FUmjFEcAckifq1qzbQiKCqW1Q
3Nn0wMnmWRt/qUHMPuOShUjYM2c344uLUP2BLVNSu9bAVtQnOSkdRhz/r/C2H11dI9D2SrCPtxuY
gE/CrHaURi36Z861rG1wmWhSJDXcd+eJpewHl5Sv0QNrB83B9s+OnhATtLKoleRJ8vEdun7QzCYR
/V3oZPjslzgiCk8XHQ7Q2tWo/lqrbTTeVTIOfliGY8pOC7B8PmgwXt9p9n+oAAeCfmUqa1qJel2T
G6ILMLUd6bLNiTKxQ7FHlO9iF09VRLKO/Tpze1tXWSK5ng/1p09i8teGjbJ+y56SUU38uLY7o+D4
5y9qoI52K1KIj6SPKtUSFmW5JJa6qbxE5+Uy5J5z5X7dNxU6YyRKIUahW0QPL8Bq9RgO07e35kpl
9gbufK7OlMelyxYk692bjGwkoIu8z4FBjhMeHRS3ZP+v0P4MtjsvrcAm4t15IPwL/KUAcb8Y0n1G
B1TS9lzUcj5gTTyXfnbo54+iSV2lO2JK7GTu12Ypcp39EHn2d7F0xNPOHje98RN8gSd9IlAFXWM3
z8dT08mLz1SCDro+6o++AGdT+3p6Edamc1366+DOh2dBwJ1Ysig3kQHNkFMrPQ/pwUn0KoNFZH/h
Ylj+B1KnlkkUc5a1cTOLmpgpYK4LNLYZxD7ob2dES67qQJ85jEINiGmv+G1GpeFgOyzgZfFvV2eY
LjGFjmTQTGzdMC90J5VKssEi0u0K6jenYFzPCbKNe+JVsyW0NPM6ke1a7ml/UIuRwpczAVsMOsup
OCGjf5gq/DyEExLZduSv4scjOPIUFn/KEblbYIYYfM6wk6UYHFENsRD8LUHU5pv+svuZSbGenOTO
A83y2MV8wz46I81/Ik4HopVOlnDYrfjMW3v4dzWGhlFEftw1ZubNvCZnkHDQJM3tn/dHgegCRpfX
VC1PlaX3X2uDKY4uCPG+TiEYXejm+KXl8VqV/y5z2xxjMMT28SZgzGH/xxglulcxpoV6NLXHy6Hv
10Ed0eRr6LnFIIHD05hllr5sH3jy9I8MsA9N/jp7rLCYQ7OCI3l3qFCa0deIs7ToCpRrp4W5gUZ7
CgJgJ3uIvu2cWMAvKFEyncTJ6Oyn4xU9GoiR/FHrO/M9bWFbHtu7Om2AAOBdcpeoUw3OFthbG3Nw
4Sfu8tBOmbibHNHkhvzcHqiCBe5whzdZAYqqrGKDQH0dDGX0ArIO0PER4hhdZkNWU8Q2DZsJWLYI
qeKR1qsXlLULv9l4bGarzFwLv7VM+/rMF3BYbcGqklRzmhSV+mUDTMDnOiqdeWxilvHnodHWOOqA
qJc2AzQJ5f0pmag2+hs36HGdb0cezbnv4vkxAOcjzVsmFW2PB7igA6Y7Amn5NhcQywcq0vEiBWVO
/ckL+mxHhLqHpid1yrmXNW1qE7jCYH8moBAmdfXWcaAKpX/Yy57uf93SrtsKQs2lvchV3KzjyQ03
Q6IqYOF5R2/bSafOm41SpqdAg4R9GYRr2/9WxVbanOW8STw/Dgnf63uapGZgJ4VVldQA8oCOq8Kp
9Lu+ojUyWxcHOoB+4P59T+jzqQk3z5iwoNlURCicAUHCTIQoZRjpP2VK7zHr7KPqmGIiAGkEQv3a
OscNtcj18whXEU9lLar5bWZqiRK+F7nRl8LY6Ym5hkqBlKBrcYbpIcBai83cO8/8UquQkPk0tb21
YVXSMAJHClUioGb3hi6X3C+9yNcqv8ldDwoNoKoOv0CgvGhwqpkJbnNTj7l2u0bbuLgKDfbeeRYD
7JSBBqcS9+8g0TrA/IfGq+/iUMBv56kfECCqWqPsSYAusi2eR6TxwfqbaH1Qb0U50mkQy1/2LOoG
/KHVAsSS6RcPnZEd38FU+ZTehos0oqagrfKH95SlYNbbRwoZdsGh3a0eAZVQIRhO/8A0iLno01uy
6rOsK/DA+xMg/mS5wsKc9JAoX52qnREVxnZmSgZ7YyN6onFytyoIPUp3H3qpw796r/2IByrZ40tb
FJoXYHycm3v3O6Y09Vwry3R43PgFn9j+FT0C2FZVTSFlb3NcFVqM6jKPLSxapW5S0JMEj9aklvKB
Gucscr/QG++861qTgXuUGWH6SlMvZoT5ERj+aCIz+GHguKnlTLrMhNdBeNg1dUhU5wAQ63S0R+HN
2o5l5iXoOvEsfppF+HtmlPF/2oxTmZ5htMN+bXU5PeK04FGjDLoOqyHyPNW/QLnmLfZ6E6Ubsv/1
PZSRBWUXcQPEmG7V8kLN8aVm7o0we79agczcPlu4YYm4uEvHQuTkZ21QifYPceAZRnGTv5tlPUMt
Nttpzh/HgQN6igvI20wcYhnnEcyqrIuzGtVsY7UfLIeOtJRNosWFRGMBC16Z4blIhSKBRTWb9nd2
Q6sNJO4LX1ZKgTmGQhJCstblP7JjwxtYl7DASHLsEAacyYHWoWL3UCY2a8t8QYTgiQVYpd85MrMK
Ma6DHAOjk9y1wGHqBVifvLOEUOM43q3t18Xg8jnHqBkGGN8ct4ZuLLbejnJ1rmFg3yCIPj+X81az
GhDjKliqpRJA3EpjJAkh0lY0YbxrzFVoUBT0KlFDV778InHhMkTVJbCkrQJDA7OqpmFEfW304SKJ
kUiCO9vjDh6OfbiSQdEQ89UYADwxdYvuLBebr4IBLBA1UToKUZYeHSs7NMUgBZ2+SBhlYJS3KHSO
6rfJBGb9FoFZ3oSvO3+ktuTxgpqwuZfmpP+Dksd4/xRtirN8dSSHofAwDTZy6pbYFP1sM1C7J1Rc
8qww9DWCF/L+H1FuAgz8s7qmmzwxAQW2iwx1sG//nsIJPVyYYJfHDNHuxxSnJiHAfyT5qd3exnWO
/C9ZzSME0LaJ7ECAG3pPqaHxEygoWiUL9uCzuMXW12XYnQCldQbQdTQaXHBdH+xHCGofORRIbltp
9c0PNpacQARNKcixX3w2FSxyfOgL+fOnAUrWnun/Y8x6QN24XWdICjX08V/kNJ4ejEFntzNKJ8F9
vCEFVb5XSiIPy67HyoKt+1FGXqw4b4oQQshFbabyQGKm4SSp43POyl0zzkwGMgyolh/llQFyA0Ek
YMKebFtj1d2BNl8sGGoso8aPOkUizfTOrUxtAHIeeEN50APWxsh4mOpe1CutGstPi6Ez5zHrc4nk
gKAalk8B7WJNGL4bBZyzfZnmSDeSlbm3T9z3CAnO6hHnmvI0YsRDF3879zRtCJpBJ6O2pulNlO2a
PhK8MqBNXFuBlzrdkjXp8bzZUyzEVONk04OyLB6HbglZelV97438adJAfo+SnHaW0HvA+pMRI54H
HzhPAQ4gTeoaIZFIRScppDNYUx/5jAp+OItd/UPzej33WCt7JU60K6uQzNwZRN/lhJiYb9JKE5sR
+XKenrhC+SRQBQ+oj6jGNaIbxjg7jAomKHsh4XeEpuWxa7gbagPjBUn2Kv3HJpo/5k613nplYG3S
/AsuhHtPdAAIuIx0L2ahIixC+JCTr85FC3DxT+ooXpz7341D9M/JSm4tKuE60ylDAzR1x55WlPHA
OUWE3kWMooBJeT9SfKfybxK6iyQCgQ6yyyEorI9Vj27uxCkvkDj5WhQd773M93xL9R93YqDp57Hz
j/2SZlMNGce5D5Wb6PeJGl9y6qERnYQZ3/4opjoSA5G1ezFeoayIewI4fxY0EX4EM152cBhuarww
oJXF2IOtROelDFguydlSBohWonoL9CzmSn2QjRtPtHHUYEq0wFAGehvLLLVFi6+0X7f4LzRnDdWD
Dq1vQC87fK3PsszbHNgyLcrjxPm+UIyAMsz2jSQOUXG1PRWUUSjrrmYdQJ3AOicLw7aqK66hQNSn
AsDDFisYmGhqXFKHgcB4mAcCj+JgctPTJ16fDX6c0oNnhL09j8S/+T1YxQS/0Wa+KUDgQdQm5uRY
bp4TXTdmeys7K8lV8hyCDOMlQEE0Akjl/iRbN+3ArE8AK5Te8HjNd4aGrZ5hU8kVegC6YjIwaU7f
WRI/DLmuI92bRBeDIuIcUxDeHUwnOrhHLlTNuXwjwQnqYMHSAvHxXGmXTFRsiqnpnzkRaKYr0+dZ
FU6KQwreAbS/dHZJR1GERbg7vgKOEVB/okjwLkraYnkQZ4MSixzER+h+ptZVwrtO0dSQuDGdd4yv
5fOE8lk32vfhppMXVR6HkxSzswkOnjrw/T8vz2lbF3GVyrLYChX0StDiDOB4wW/GepWIX58m1V+q
sHpmW7hs21rLhTwTicupZxf9au46yu2aMF6wr9fXsvBVsFWwR0nwcyHiSbZhy7x1v8R7xo+Ju+Jl
sWm9wbdFXGGDkiUx/5ZGYnzgPiDtvhE8k55+I/U5VhrtOKoXNCpLr1q7JxDqJ/cw1A6oNBy/qYbx
T82jqmklzpeGvkV+R2G6p46PRs2MFo95gUkSjD6kI6o6NoyFGUyob0eqBB8sIXusXGNkzRPimVrn
f13pQQ15ByHSMxf/n5HGb394/CFKZ4LKwkkELY0Z5DO11QZLQHzbZZhg4VT8CeV5C8WPQAcTKPvR
3FKBMy8jYqriSSnRNVytu89nqeQ2reBU/b2pQ+MeMrJy/q/AbzVCToxxBEWZBd7nryr/i8+YiZJW
r/wT7qi/Di48CkSmJWar4h/4eCcFuLEACsgUJ8mPnegGI/XD/L0xVpQIZ2U5vs4Wg+DiTEhVQniO
iL2Lao38HadoDuoJZwLVspS5m4z7tdgnWJfhUCL3kJpR7wUWIySMzodBxhnY20KIdW83lNcHeKkr
g6reIyX4APn6zuLqZbPmJ5G84VlI4N++x74UFvsyyh7dQ3vS33h6rWJB2mjR0BrlCFkFTCDZPnvQ
NRTRaSdVhbCQSbdDhc+QjajuaGCXBLlW9hJrSsCUno8Q+vUKARkPaxQWHpEYZ2XbSzpTIcWZojvs
C/Pa8/KBQw2JcyoDLjZx4q/ENO/Z/uLWhI1OAoncLdAZbITjqJES3Z/6CvkvF1N6iivcbXNRsw6A
5NiJgFbapJVzj1oEhMX7zfijHVMF+l88xoUuFBOwp7AlO13+Ca84TBGV0/VwkTsQRN64FYFNa4KA
99h44Q099hdvNr/9et4nEccnmIcpocAv3z0XVoH0CzeWEY+Z9GBwHj+Gq5DtIH4aX55KVemKE7nA
cFgOCSPLpLo8p86vjIsIxgsTk0XSqNgMqBAtmbHLtshjMSnRsZNvExS1Xn375gv7y+fqAvl+0GNW
pCPfCMXKeOSSRESrr0LDgJNeg1HRVF/qnomfr84yLyRy1pyT+Ek5IPoGCUHpcWACRMuoRO2AN/TQ
9UXnqpjN5lCyxvttjF/X3zgkxxm8OlyjgDkzr4dchpdQFHBSJuN4NWKNo7iEHK6MHzdJwgfm/EdH
h2RyGEHL8028gLf6Lz60fBR1x2Pl3jmAKNc8UNt3Aoe1fLlBeIJfWaP9lp7MyJlhOG3eWd0wlwRe
ec2L8aBh910n+qu6gH+TsTsRbusR9lnU/MlWNDhVtlIxnfRsaqjQicjUUd8lswvA0y1IdlsIeoIV
lW0arGnliHZjgScwLmCP8eYbgmEFKZSanFY3BArpF1boLnRffjdYnJs+H/WMbWFedbGWjkrJuGiC
pU0o1aQGvsJ+v4+5DdVHuhCWC5KUpvcthjrlKIvULMRdnMrUJI75BsZqgyAa9KOm0xoKV+0Xp71Q
1CPWkjKqW4SkJgk/xr6lPSJpJiuqlFdi9penz9/Qy0NQSEscYBs3VJ0Fo7zLNT4EJXtSLYqiquJS
Q69AyC8ah1fewpSw6dB+X5x3Qb2OHWI/FSoyTrlsv1NZtIhofSO63A/g7m6tUlaQ++keySqs7C+3
X4bCImg0VYmyusMhO9E6e7uNgrhTdGVrnx9uI17D529uvc8CUurgOpcbbsZQ/S9Jau3HU7hAavPS
Vbs/9rs++zJFe47rdUt55rEm/7jtnx8gUrjplLXyRsSE5OnH+ervhdXbGHame2MrjBwVvQfj1h5L
QjM8mY2h7XF9EcFMf899BzzqD/k38GynnSQjUiVbBUgX9IGwIthkFf6Zmc58lqcJjuQAgjbIX8N/
OUtJuXErok3VLwUoL+ECaSOZvIg8aDnZ2QgRW9AoTyN/I86vFrLsi5k2eAJCQnUp2DvEMTz3fipu
PebS8HPZIx2mkr965N+7h5QY8+AEApssY5w6+WLWkSgaZymw6h3nkWn9ZOI+4XfYm/rzC6GNEX14
652tW6ayxjQA+13R8ZJ8b/cTZjfpN08adM46y2SKeXa+gkq6T7y3iU3B6ZLAf/pjhc/AN1NHcDkP
SnQ08lth2JucdG0b2chXhT6YdVsHJ+/LEjqU5uMm91p/jd/Nt1i4RD/BPIODep85ktOv+V5AR6y5
/7KKe7tFcto4CTFsrGJ5IIw1iMt7HXGkxQo5ft7oM7lNkUDn6fz3XuAwvIEacRS+hLs+d0yXNanF
A8tTdRa0y08kZMeKcbjsS3cDRnxW2gWD0WsfB70gF2dx8VuNLv0fKZNthSaUuC/sI8kJyksp0ELr
eqt7287QdJu6oefSD4bMy7hFukmKYLM4O+pPx2+VOezm0USOOoi4+LXweG/DQ9ajloWHn6zBMP02
Zd5rohET9MhnPtJkXkCOjCTPygCFXftJ+CAA7EmHjNuFCQugL0wPVsB/mtf2YvUqigcht5iw19M0
aDKs16tX6jxGuKsTaIROjKsbNmnHXpyVyEtKSQm5G4KJvumkfBS0/Px8TDc3ik5Uc2CPqZPIH0pz
XuOowCMOoncqDdo05FtiDt5ef0KFMeC57xv2249zYIeFxL5EdnfYdSswyB4LbxDgel0eVXqrd8Yw
5snEbiZ5atlktuaROVFx8pdJsyRo41CWgrCMKD9uj6VD1rDOrT3bgyDqrlFZhgxVEZwCuzxgVLD+
CAC/hj60JQ86/iiDRJhHDNQFnZi5DxoFjaZ0DcwC01IHlLDlod9eiWbKnU0tHYurTZJiztH4oahq
DzKYLWTXlNSilZYdxHgtTQo5cdu991OJ987lwoHX1Vvw6LDGsBuMI4zpbWFDzBJA76HOpdwifcs3
4WV9H7U91nMmbQMHWJwTc7U7FGZ+AfH/RXuU+/mUy/yvQC30uHE6j3cd14HvK9WhEx/sWbw/pGhM
+VWT3R318SQB8aSkKQvIYNzENR9jx13Wv5RnrWAgx59bF+ZvSOQCJLoGG7Rdt4r1Y9riBUv7FOeB
kj0DIu44KBhesMohECNKtc8iKSOX1tsA6/5mT6sAs21zBr5ueKpGxQg1ddcoYxviuDP+qdRm/HV4
FdTe9LCF0/vGeIQC5ovonJFTmmUU4Uha2u760eRqnQf8Id3bqnSgKfU+9+RVuigt8F5iGs/CC1R/
+Z6OdSDzMoz59/lz1aHqIi9bbgKudb/cbG4b1FEvLSn/KV0BoDN6OfZLqmld030RYXOJHOCp1oaQ
q+J6fJ2z+Bh2UlL4dGo+E8igddQGGCh3RfQl6heTqT9r5n1ctbOIa0HhPau+SDVNG4Bh7a/Js7el
x8eR3niqi6cuzujyigF3L5zV7BiJqXYW7vsziyrA9TVpEB/VZVhR1Q8KZ658DIxNocdqXTIp7x87
ZmRUeK/eEsnxJmoeTbW0mGseUU02/a11toBhzSc4HsPqkrcmZIMiRUxrUTKZ1vKDdkMYLGEsAgUn
8WYYzXcUliqFt5/dnHDq1E1fBaH1O1UF+ipcxStVoWuctPRwHJBWV8u0wpZ9+DxCwoD2fEFozi/o
FhdqxpV4h++GoTeglvL7UzOsC4wAC+pOVDfhmjnAMVriH4H6uql3LktaNDM+WwontggTOGwKXMW/
kw8o4FECUAKGdVbRAQOJ+996meRG30ALFI4DOALU8i4JufBWQEZNiL/9xtuO+TVyUAyYeFwbgZTQ
dwkge/wED+YtfGQ9MmHWstKkr5w0rOfTFxbhVhSHl7MyV2VQRveqHn0Y8J7dgIFg/raw4Q6XYSCN
Tt/KBspVrgrj8UUn4xjX5DitIEY6rN43KQulZYoPBsqL34Yx/iriy1bdJJ6Ojm98UR1/Tgj/OvAQ
3f1dhn1GznCU4W7Gr2UKWzN3LFeWzjrAKc4X245rEQvbcjEdk8I+e+9srDevKkgfXd2e74G7e6d+
r8fwNLZycyqHqzGgeXWEeFN18+C5fCxvwEpvsSHj8TNooEEIqo7lmORKCuM0Oxe2wSIJWb5vE+Of
u1vS13z+4CA51ZXTBxpAlyb/LaIvNIpYOFaZSLbHa3av5ADWepiyOOauG7DqX1qIKbzRVAns2WNy
k5wRGYStR3N3AOInD7DM1g9XC9TMMbatzmot3Z3Vn9keFGaPHqoUsxZjkpTy+xs+7iijD1/sls7Z
Um7cZsf6JTLo2qNjmhSffsyRkRGkqT5IKt8syuLxwe55BdwB7QErXAhdQAruMl6Y5J1JVnu/k9mm
hvuV8lppq81yhPQxcwefATz9K+RPEKLaMIE3tm9IWDmqHOOecbIbG0ykkGeVTu5XcI3jHgGVtEUw
h6TqaeK3mlYTV2CEtF0idZd+02WtlRdODGEgQSHOMKgwLJbMOTAtTbhlYjKDmVS2AO0bNIK77Uwr
sojTzkVq/D7MSLHy8VqeBdsN1gpfxaBYcTl2J5zM/EDcvUL4Yk7LRBfu55r6Pyks8L62xSsrjJ51
XMoHTGIAk1MHwm+LTOSTlVAbfbF2wwOW4Y7dpfQDuZaeay7O4wpDJCmoCX+NypUzW+/pHa5FesaV
GmKeBeYU5Y5iKFZz7lGgO9cgeGewqisZ5B6C7UykH/iyshIwQUEK9Q2cIRGGyqMurm02JWmT505C
is7Gan/ibFCK8j7SiJw5EwW0nned11XPEccTYivvOVFsg4mvdlF2K2fGCU+e0lrKYa0Ls5KIE6GA
6Uhz69BYBjL42Y6Ui4a2PyEsq3ckQYyy33m3StgdHE7KtBUYsW/HRNojWZdN5Kuy9+hxH0YgA8mJ
V1SpP7j4fsJVSCnYxkvWm7KWbB2VU9QvxGi/SviCVbPMgL7hXir3k/8krxQaNvmox6M+3UZLGcNU
FsgmMvws93IpyF/jHb3NTSY+IdtJ0C4DBRjFyMzGqh3hVXRIjRCYB+NTJdMLGchPaj21n913+Ppi
rdRs4g+EietvGGBoRg0V3OUd9t9MdLu3vQZiwDwXvs5GCxW7VbdepvTFNDKIXvS8bjmN9TlAHoX9
43L+We1umQIxv4g3wc+4yUw3iwOKUjT9dtGDvSfKPq3xeQyqN8ZVvElnG/8ZKlxUoev1rtefhlup
0xm7sT9h29JPWLJFbtbkOjG/ZUZBzpVfh4lJVq6lcXp3A1lWB4hHhEa7M8s2vmpnOiYe7+djGgjA
67OftU+uhe8THzEUeeoqcUmJ02prqiM0i19VbyxB12PYSfe7y8zEIDVHM+mjt+CHLag5fRLueuii
jQs9oqeL/l4kW35N0I8SP1gXfWgDcxzZTSWfWeEE4rTbgCtJBpbu9VZk/v107wpxD9XzJ6GyR9Tp
p3A0pAtEcCVx//CTjhxlbBRwbVbNaXMuhP839mw8tR424sUs8ksYuO0sGzPSDhax9c4Y+MMB9P6c
co4nmZaKWwL/M7Ao0Swf1QqgsZnOwmHdrSodC2jF9CZqjTwuoxCUgX88uaRN6/05BPvecT6WLAW9
WOMzkqTMs45UnSgCax1ekVrzsDdz9JO4b1GS2gAKmEuevWcH5R3nYmR4iZmOS01b13H0HFPM2r8e
hF2yGyW5eu6dJHwCNePkFLI0fxJod0G9M+rDAdhNNr+KP13zP5oaI1YGRvmGSFw4PpNnYQqYAJXb
fNtG+bC0JQ1sxMnsos+IzfZu/s9HTv+NVwd/stQAv1DxJEYBsG5Wv2FfV6tp3RjBwC1jMqvlUwg4
c/hZR4cCzBXNTcihjrUs3rpiWKc+g7n+1UcH9G0MnlSHbZR1pajIK2P0IyUSYAmvxcgCGEmNjPUh
QoiwLPyuh2OZ4Acvs7u37Ma5QrVz+IsfgdCeDILkf9HL+wUFwmqZnV+26FWRoyR4UKoItA5Y4yuG
2+VPQJZd0/+Ko/wLGjQ8Q4dvPUd3wL1PxntywJES+5aTSaGERnJegmsp5j0oWrKdV41tI37rEBoE
UvT3ke2YpbioEnsYGKqd7NE8mqPJh0bwrq50pALut0w3v68wV9CKIgGU4oKG4fArKrvEwsWdFe8F
IcKU8AC+2vVrniyZlSY8eGZ678zj92RYrncs6Mb1zLyLapWcXhitIcI6uo6qA0AYK28BRjOrM9Sd
cLRRRJsNg5asALfq2dEnnTJxrouFCeOBbFSgo8rIr6DalS6E8BFM1Y6szPbmioJ+m7v+jJdFgXQu
IL5B317Bd3zXZKhyXZBTxYx1GtlNymeNNgwtbbojkEZ6jqjAUWn3Q0wIU5L9kkfc5CxFqCPJSFEQ
gILoZ1v3A/aJHuObf2ZKpRhgKjYe28AzuBZpV08LALzQX/6pSg4XcR2d04U89g1gqJvLLuaCKPiv
rhJ5yb6lpEjh8wplTxRcEjDS93sWDXXP49sKfV8P2DcPnBBldDQRLNx5HHdXpH5y6dLG/zYesnlC
5LdHKLijD9CZyC/mzPA06hUlzbON9syEMQtdxdeARzsTgzYMStALGUcpflDQHWLgzC039hyXSyT+
z6fMfbWtVgROhgmMDCM6B638LR6JzIuZOzpWUgf9OTIq0fmlllaFfcbmC3q1jZenwng5iYlBAXoj
U/7LYmD7QZ/W8FRCiEs9wZ4bLTJ1WNQYsNiGgTwqH5plt8tobF7VEXx9+ECGr0hPETrPG2cuDbpF
7Wd+WJysJjC3YZz6k9eiGc23xobC/UEvtKo4qVCXg+Lyl56tkrrD0frR8dlu5iMsVEyKpZeeWJtp
WWHkQaHavq7kLs0bMZVqlxFzWDVkDHNfyR9Fs1qlcWXjmHOllWVzL0R0lEdWGMETYsuUui7Yzlvl
FQIodR/s4NA/3nWUR2iUvha2EWQzUpaQOP+l1RjVhM/IZN0nn/rFbzLZs33eXG1FuYR85lD/hakR
92ULgoiMauiLk5r2yBIvjpRe2Cnthl4N8KcPWCoqC24HswVpzsQIMZ7HY65J/S3wagC3RBlgIvLL
Ihr7CU9GCrBQ3G/UrAmixWyNS1FzkmurruA5N2sOqA1fbsdNNiFs9ylP1C5O0bgP2x4blNKHKL3l
/HlI3vUq4W3YYO/6l3N/ViuJKTwU6c7Axgzge12AsA2OAcNgVCC1tee7MgjTrXhrkMPpKe13qDJI
0RiUWXRfWj/HNQUudzbEJSPJJptCOY0IK6gLnmRMzmqzNlIkcoWFFHpvAq+t7EXmdmja7N+VkQ0C
svGgFagNDZ7aYWXt0QzjejylZVxMYDVqyFgmJ/kgHmrRJDPsByIhUKCEfZpjlaYybwdIss/+Slbt
2IkLwortxsoMSdn7bG9vi8mFrTw37tBeJCK9v+QEgO5rNU9fMM7V74zWnZ55GK5IFAIarg9u1CoD
PLVVIXczRljO3vODZ9a12AOTt6PP3Yvu/BGv72oVqPqgOVV45w==
`protect end_protected
