��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���!V�!��f�%��5EJ�Q� 5f��n�8�+o�5-���f��8�ߏ"?��a����eͮ��jn�?MX�-eє�
*O^^8�M���lr�0���,�X	5�;�5��;5�k�<�(�ǟ��C6��e�Ϲ�8��eq�f�����7K�s��)wRgc���J���R���vU�l#��o�;�J�9�ទrǞG	�^5��e�B�u���p(�M����I.�c�)�PCB��6լ��]蒾��T՟����G�7Qߗ(*��P�sW-��"��A��aQ:{� DuQ=cx����r.>9L���9>�#����	@�����ڗ]*�	9�nq�}&%{�H�\4��b�s�i�vmVW�(<���ĕü����>4�JʌV�2��2�/R���_S��w��(^�N7Im�<M%ÈX�y[����Z
��z�+����!U���~s�=���@-��r7]�z�����u�#^L��d6c#o�҃��VL��"\�5��$�wcJpN;�T�Á�\�Ø]��>s����l}������#u<<�i\h:����)Ԫ����"��,5��[4a�7������U�<u{�Yexsu���y��<`/Z���o'րk��n?�QD)7�����J���nd3����5)��&�W��V��Ѣ�i�O��H�ݫ�ؒ����TN�'���� ���I�	N�l��ۻY��u[�r�]���.짶�@��Ա��u�Yt�:�������6fbpt���F��&@�{�.��8y\/-�T��:�s��4���8�+�+/%����9~,�}K��۰�wq�l��)������no�E��w�'��� �( Q/]׈�nyP஼��W\��t���LM�U{�nc�7�����]k���%}qktd N�;�7�M�M:��CЉ���=ss���^����n�+L�٦�����A��2q�n�<���?а��9�j4������=�G��Լ$yd:��B�D-^�����`&������]i���S��b�|�N�����@�g��k{���,���ݷ��1���{hc�����]��1p���!3�@{��rE��i|�3R��w�W ��7-���~b�
߫h�)�1�ˉ�Y����`�m����R
�)&��?6�Mz0��M�:cB��8bÙb��=H,�jډ]<�욤�U���yʺ��$#�Z7�-��o�ƀ@!�\I}��������~[us�FZ����h�w�SH���ֱB��a �%B���|�H�+�t^Bq�5�����_gL�#8�#�5�i1m����x+���m�P��s�#o�/���a#P��#7)��x�?ۘ�$���~�k���ԍ}2e9�����Zư+�OD����Xi5�n6b��GzͪH�36�J���^�Vb��g�t���	�e��@�J�4�6��p��g��t>��3�V��K��e���i'f���Σ%�spÎS���`�-ڗd�E'Y#ָ a�R}V��mO`O�9���J^��ȩ�l��}>�64vjS\��iUgۅ?G��</��j/����yK�� '�2�`���}�`��W�{�n��1|Lз���s�*m�P'J��ó����9��Õ9]��ŧ���v��X�r��k�&�<*��~%F�nW� �_=�����c���h[ȣ
�M�ޗ��&e��1��|G֕Lf�\��`p\�t�B�l�Q�i��(��c�D�C����- �Lu���Z�Iݪ�
�pG
jݡ�m*�e�����]]ԅ]����w�۪9H�jU��FS�\�8ap`������<����h���|Tk���4�s�P��C��d{y���h�u��׃X:T�a��r5WJ�ɘ���/���r�
(W��<�U6�	�w���y�6�[�U���A��]f;`d|��q�xC�GzP��W�a�+@tKLB��☶q��������Sct�@Bh�(�}�2�<{�R���=,�k3dV�JT�����:љc�C��1�x�4㓴�ALЩ��0�}3~OX`��`�.¯W�-^�]"v-`�^�����E�vG�J���i��ƄɻiAg$Oa���}��j�Z�0^��
��P�LP��"|��%��k��̕��j�:����ڂ����NM~?�[D=A�*�.�ԭ�迯�`F�G�{E�ަb�����;�j$����v��0m�}��j���^cs��ϐ�QO~S�1Ȧ�R`����+d�	��; 
g�H.ʎ����"ݢ~�"�:�0�f���m>��3K�t���L�aMUrF�����PP��|ë�Bl�uzۊ��U�ι:�@�5��\,/�il��;9�$Pg{���W�T��}�9�ݪ�Hc5X1�3�HA;�V��[��8Keg�w9퓄���bSM\^z>��ĸ@����>�W�,bj��"�z8������5�R�N�t��[O��Y��)�ۤV��A|u����-Nc�Kk��
cgG/F^�,J�.���g��Ylh�s�}��e*��M�-��ǀwl����� �Z;6�-�K��˫<���ML~����1/��b%w�*�q!@��hk���7���������3��!2��5Ze�L*�@:b6�<����'�]�NH����)��r����䛿k��d��M"�j;�wh�'�F�qpŨ^;�V��NH�Oݎ"�|��=�%�ֶ��R-咁����&�:�&�U��0i��E����{ڄ��]�ډ�6�RL�p��)��.NX�٤���M-}𼂫��(/rɔ@/���i�B��0׺�k��K^���A9�O#1�oVJ�yK>}�ś�κ��%�p&�Y�ǜf
���:?H�2_��8}�W��NfN7�g�?�<�,l9�-&+�����M�P��U��J���Wc�e�+O��2�R�D�uk�l�Y��<j�q��,:�gW��:�=�s{xQ�5��k��W�b*'DqR�RS��/�U ~�;U8�$�	"�Ԑ#��PQr�١���1�y�R���{#������[���$;���}�ص߉(2%ev��,�&t��E�*�x"-�%�z�%-���c�K��4�?Xg����19�E����%
~Ek3
���H��
���H.�w�V샒���Pc
���<�h� �r��߹	����R�\B��XI�n���u�g|��i��� ����\�1U	L�̤�K����{�[%��E
�w�i�⪾��� �p��\��zLX OW
hH���9��g��<H9�/T����8l}�n��fS�H�WMV ��?�]�)�R�"]
�ޚ5u��i˖v+�#��ڼ*�bzȘ�����T��P��1i$��G��Ԏ�>�U����o�$v�b���S�%P�:��$�<�17�H���#�VQ=g5��"�k�ćZz�d���X`�.�|wj�a8,e�Ɠ�kv��CO�>�Ǥ�g���2�,:�%�8M��p������{�j��!�+T�l3�� Vo6�T%Xw��Q��V�k2�>@匢��B��ΦS����۲�3On5gT:�j�i2�ىv3�v�W���)�2U%�i3k?�{w�'m�/���ܔZU�(�ED�oO*����G�U1��lѩ;�ו�)j�3�o�����;Cjf�|��8�*� 뼖҃Vi$gH[c�_Vj��OI)ч��fJ!��]c�a�:ʗ�����/@�z��?k0������j�D�|6�FC��$z��.����y�sר�,��fTh����q��_�+��<��2 ���4{0�򛹤3i����S�V���e����&�l� .��%�l����rh��ڃ]&�"�S���HM{�����!�k� A�/�\�)��׌f����4��Z�B�]P�Z������[Y�Tb��r����z�L̋f��w�p�e�~��xW1�m-*�(�PI�`.���Ρ�θ^���E���:�-(.8a.�<)f�����m�~�Czs)h�w�O#O�Q�P���E����I�Qt���9��	��NQ ��aDK��'"4����ɬ��3��q�J�~M��Q���N\�i[�{՗�HFxƠL�wdo�]*��1�K��;�,]���C?�=��8
��,������F� ��>��c�͒0�f0jf��X��A�n[�������{��=����Jgb�끫��Őz;`:j�5/W��'��x*��%��A'Uc$b��_��M⿚G?ɘ�)hÄ'��(�z����c�����OZ��p#d�(&T"b���F��Gl�zo�$M�0g�e�ͩ�[Ae���%��L\�I��p��3���*��b��dΐ
M�8�C'̰js��Gwa /M�)���b�8鱦B�������Ç�	�p�pBؗ�!�m�+��l~���,��N�Jh�-|J�r���߸F��ûm�{B1o������A'O��FH�9T���w4Z�t6X�P���ȼ�ă�ǔ�e)�Ƥ,��R��~�@,�s�S�R�I��,Q��
��SM ��>1ra�����7�9tT�1�\ Bق[H�Y���E���L3Ŧ%�|�?�pÑ[B�ֿ�/wv��u�0,xJ��*�Ǩ�~�w��h��՟��+�E�ݔ�x��}�T���:.H-���]����W���x�5_&"H�y��Nm���8�X�Mՙ*�����)����Z��m���nsb�ᒉ�H!�BJ���}C���z�w���ŻofU����v�nnt�6avL��l(E\K�A�إ@ ��g�5~.���|�΂����	�<���$�1�����0ւ���Ҋ��v�e�_�!a-���4.]lS����Ƈ�c;1� �zJ�B�a�[��f��fw��k�"���z_%�M�h��kGf�NW�}3�Ł�M"�Ւd؍�H�c,\u`ؘ9v��=!^����O7eEo�X⠴ 3ո&�(�����R���m.V����k/�����9��C�����8��^��z�~������2us�;���^�S\�`�ң����?T&%��������!y�c;أ�Gߞ2[�Dt|H:r�LMsHm����T��z���Gݪ>�4L�u���͎Kj��@��-s�͵^�^��2C�g�\��@�A@~�`�Sx�C�T������w�W�F����Z�H6���qm엚�%��(�8��9nr9�d�\o�ȱb�����b$��?K&�fR�����W����߱�>�{7�T�;j.8�~TcS�6���96��je]ם�+�/���ʶ̼�"%+�|Pj��=�+�$�?��VJ�^BN*CL��t�7�`Uą�ܮx��΀)jQ#�����붺R��gP,`%�Aj���~_ dm��5h���$8SQGY��ѐ�^/14%XRw�m��uԢ�j@�= R��l��OB����Ű�1�@�_mЅ"Ġg�q 	�
���ך��H�q3<���>_~��/2�)�0���UebNNI�N�@�]��uH�C�,��4;
;ܓ~��9��\m���r�R�a�'dt䴰	-;�і��Z�Sr��&$b���Q v���B��y}�I�'�x�Eenm�A�@����Da�??���ч�gL�@���ʬ#�?G���~�#��E��"6�'^jw>����c'�cD:~%r<�0K!d �,�[q�PPPT�L�r��!�aX�ORPF�:�_ �����,-T�MZ�;��#��z�(J&/ ��י�ͱ��ʫ*1��)cN����Q5�CD׏��9Љ��B�!%��^��U���DP���h+#����	�l>g�݅r�2#U(����n�����<j�]1s@L�.Đ�Qa.��XW	�<��u:s��\�n�
z�k+tU@`��*�|b�Z�����>�&�V3M���335X�?")t)ϱ˳	��g����nJ-��ŐP뎱t	7T�w������#��`��̫�氒�긇�_K�|��!s�oV�5\��T��RF14W���
�DC~[%�$���0�p0J�rB��#m�u`�0��8�J�U�~�aAM|��[��n�#v�>��5��(N�h�F�sZ����sDS��s�묑�PL����V�c_�幞��oͽ��S��g�*��D��`9�rc� *d2�gx}A�k�����)�Xvso�ź#�ꁏ�JXt�esS14��+��t��	;v�Mk���W�P��Y~�ʃ�!na'�b{�p�@ü^�ݛ�#Ļ�Q�ҿRPC��d�,�TD��9���̹��/B���1�)IU|U�4e։����� ���t��-��>��J:�ۓ����F��0a��y&�A���@"3�MVK�B#���盟�9}cV�:#���� ��W�G`��	�-ڣ�H���*�}$�z,���Y��.��ǵ�Tmx͖�2iN�(T^^�l%������b��C˻YT1��1pEf{�6+������0���|�S�����9ZA���;ӝ���4ip����n[���-�O0�K�At�����WU���EJt�e�� )#�2o�c���	��7�d��w�2����\��o����W�� ����������d?���!<�C��M�}�<QQi`1���D68z�7��\�j�66��i#�W;~��e�m`]^Й��o�h��yB����w�������'�p�W���&K� ��<��˻y}b�f��u:ne�t�:%��G�?���	,g'$Y0�@�Q���n��-�v�5u!��Y.���s򂞝�<��s|��%{����~�p�Y�n����g����v<!����0��W���Տ�����_'�\�Dަ��"�ݑ<�ruX�C�4#fV8�%"T@	�m����[�_�_�9�RP�x�Kc̗C�&�Aﯬ7ɴ?��<Q!�Mu���7�33����[�K�1� ���M^���dr�)=t)7i�r�V(����r��*��u��d���Io��q�[�<u0C��Q0�e�}�L��vۜq�u��K8��P$-
`����J�A�X���y�4�a)Y�R55��2	��n�YCJ}ǐ��rŚ,��;���5�P�3�K�N��q5�.0uc�u��Ԗ�/!���|�?+PG��F�8ܤ ���,S^����T���qt��2&4��x�;Y��/�Pg�Y�N�9Lo�o��L&�����Ή>"a��i\2�T�$��\�[�Y�KF%02�bR��EW�s�(.o�S�$��N�Ľ̷P�P)�;C2�C6�@�nkl	��H4�����f�8ʓ�Ϻ-*$y/���>:j����&�n�]՜�l~#��^�J������Pw����ev�Y�X�`KV�;l$���y/Ξ$YU,+�l%y��4�V�Cl�Uͩ���MIi���[��d-�D��b,�ز=�`�f�ܱ��ua��X�eb�z�P�H$VH�;?_�1�"��V�3���	c�{%�k2_�eFbz>h�{���L�hz|�%���o6R��U��i	���K��JV���H���u?<'o�x����s�agkue�R�-�A�
c��Y��L��8���`Rh��i-&��86��C���q{Y����������c�ڨE_S��Cc��R�K#����� �����W� �-�(�G�E�i^�O�)�#��zd�
ό:[���l<�Q��
�"�5�ş�����ZF�l0��`�sX�wV6rw�����u5g��{/\#
Zu�H�F���^&�>�et�J!����E���}��2L�2��A�l�j9���(��NϵH�@l�4�EDi�`���ѷ "�]��f$��e��ňx<r
�5 � ��=oW��]�� ��)�D1�)�4#�_�Xv�80��f�e��y�Iǟ�d��kR;�|&p�y�`�4�W��f�!ץ�N�����	��J��y�Zڎ�Њ��d> ��y�kVu)�x�xWͦ3�1���=����;s�'�(kڳ�G��8@mk�d����V�	�!8?ÊE�ߖ�Jd;�!]D�\oyq���b� ���"����hR��6j�KҎuv��4�E�I�Y) E T�a� �p�T��2!�H�o#�_Õ ����1����'X���K�G.��F�sJ �Fu��-[Xx8咛4l�b����B?W��ӣ���j>��� {J|~����s���`�#��KV;���Xw���Oz�*��:A���\�S��3:JN��$�G�i2�fu-�0z�����hKZ\�&�tҪ}z�'�Hz\.��=JtH�^F)��W�&A%�v��)Ү\X��>�^R�1*��ڷ�����\���	>�0N�l�T��:/n��)n�����8�U$����ݞ�����E��π0@��K���k�Q����P}P�us�G��=�؉�#(T���>U�0�: ��z9K��6^��	\��/)`!'���՜��}eQ�����dUGrC|.yG��&��rW�a:p�o����v�+=]H���
�UUS"NC�e��UqX����P�͓?�o q1\��\)�-}��1�o����0Z<�&B�¹�G��:Fxx"ܮjNXԦ�T�`2��7C�M���z�7�Ж��!��X���=漨׳�rb�~�	J�W&��<�DyE�>`&g^� ��O�A!�M�L2�
�{3��`�a��=�W���u��$���q�ۓ��]ؑ� ՜l(?1.������wh����J�`|�aF���I���y�	��[��9;0?Z��'-�p-��;J�K�.r����QB��O�_0:�TI��]�V�4���~�o�gRr�2�q:?l��?OzJ��wi�2u��_�!�ijf�,.!�X��vW3�xǟ
��-5���e�`fH��w�Ev��L{&~��-p�3�*�1�^j9�&�ފ	��L�'�%�����񅅍ak�mG�t+����K�W�2v�j�-��A���9x?8�WE%���_$�D�҂�/jf�����0�q�.e�-De�5��y�춣����[��0�H@8(��
�N�"�	��a[c��1�G�L[��eS��M����]�����Is���82*)�X)O�����8���Vҿ�[O]1����0x3V���O*�ܭ&��"Lɻ>6�X`�Tc�޼|zY�U i��?0U\%��W��n��@��"4M5�?,~p:7�w���-{����[��*	�_bv�6I��wS+�A�ϛBX��I��%<��a<D4f�1pg{Ӫ���F���vvliD�gC7YZeg�������s%n���8&�Z�{܌K@�j���->�͑���H�K>�B��&E�0xl��0<V����u3���&���h�:(}�����d������oQ[��;�	X1{�V�n߰ɪ���l�7�b�"4[tscS;���A@�71c-K��:Y.�I��m����(����	�.�$tw�9�����	K��D��i�2�����Mx:���tL2�B���V�~����ީ�3J��5��yQϋ�一u��se�}������1
5��V&�Ć�_������i���<i�*��cJ!���F��?{hm��"���g�K�ڜs���I��AC�� ��ޯai�͊
�L�H`���x?@o�����y�I�g/`�tV�Ax�i� �<���7�)�Q"��0��0���9H��[ަ��0}�����ᥨl�(�P�/1�jc�h�����fzt�ܸA*��c�J_�{A6M��}��Ζ'��;8e�У��m{�Ƿ��`�Q��x�sĭc^�I�2�H�a��V�7;��ɼU]p'o�ݺ^
p�$�>_����uݎ�O���K�(�U��(��I���JtjGY�%� [�g<P��]T��鸛1ڇ��tߍ���ŉ1��g�|s��Y8�l�-Ld�+E����K?����NG�H�?ˣ���6�֛����OR��vMxs_ˤ:j.P�o�bU�і���?�c4~��s�DB�%��Y���y�9v�|����WZ�k���sh���e^��Z�#���ʺ��K�]o�U��7��6y�ՀYdͱ�W�AS1�/�N}��ja	k\9r��v���ݖ�&������S�ė�Ӷ�����S�_1�9~�Hǭ��Y�ӏLK���h���Y��U'��iߕ����z��K+� +�hQRʫ�Е<�Zo��p�����.�o>>�/��u�u��#����'�8�j��3sS�=[�T\:(G��k�;C>���#�z�zA ��Fl��ET�^����� D��umw��b�,���p��5x]攒S��܃BU�Hdحz��`�mP�(�W~?X|�7u[[��DOJ�P��-�;Xu*����� 9*,lUqS������	�b:}�F��6�����7��
�+����'���_�R �W�/������,q�P�Nӡ��Z�N����-_�MXB��!�OLCRC�]����jp&��L�>,��s|0��{;=��-��¯b��V�{'�h��+y�5 ��̎�,�L��7�7��0[��?;ÿ�rK�RlqS�2��45�VAr^�@��eua}����{����9����N�['4�����ׅ�1��M�m���-��hu��5�sX�J���S��b�����0)[2+FX$-0?�ɗ���3�����/��m8� 7N�ܶ��	��6�L�?�[�9�D|��s��#		Q�D*,�r����aR�V�:�	 |��C���*4��<���cE.�8���0�5�B�5�#S���^���_
��Ӌ�BSNw�&�rS�Y:&�J?��$<��H�����N��1wG=�.̇:~!���
[xo��1�u!l�A������F1�9��VYR'?P<���Zj�R�j=M��3J
�!#�F4�*�.��z�3ǭt�Qt� i4�(�!>!��34Vt�GN�+�-�X��˯�^C'�|,�����)0|�.OZ�����(�$��1cO1D7j�Ò=Ǘvtr؜������c!���с]-9h9�B�k����D.�#<A�]����F���HKdT����4RN�kj!^�k̀_������k{ ;xɚ�j�p�<|�@�+��FO���^�\�G�z��/^�]%c�h����Ww�)v�aO�ʑ�nn��<�C٨�~r[��ԍ���-e���	X�é��T�~��C��N�B�ů�Hq��'5-kF		�����H.�7">���6��bN㵌Q%�!�t��@5���� �܋977$-E��&�K���-����t�և�w
ɾ�b���JR���߄M/W��*�5���f�aW��E���4��!^���v�<�@nɶH�~q�&{g�I�r }�A�H�ÙVr�U	*�)O�S�آcPD�l��2
C��w��\�;��4�ݘ��(���>�;z��6pd� ��KttP���:�.ǭ�Dk5��hu@�Dvq(��\��5b�� W�n�龬I?�o����0���<�G����~��cd&M�y�*[��:�z�Y'���v�J��ش�ɡ��')(�����m����#��"��V�"$�Ih;��H����7ȩ�:n�
�!N�6���nl��f��u���F�y��Խ�j���狈�X_i>"������<ܰ�f���mn��$����ѷU+]��.E�+Jf~@2�!B^��� ��m�� � Up�6�#���{��>M#A
�bkRvZ��ۏ#]��M��Z�<i�\M�	���%��C�d���X��D٭����Wg@_�?�/��M4��S�n�o�����<���Ý�o�b !X�;A���b[p��ʸ⍑��n���+���!�,
t}�� f�@�v�L@�s(?����p��'���$�<�dRH?p����}��/��Xw�^2��ݣ�sj&\��%�*X^��V��6Q��@q\�n�0Af��w���<�r�/oz	*�'0X5�b�ک���'�ߋl�!����v��ybTG�Y��D�>�q��qmN=� l�`��0u�t�sw���I�T<M�d��b:�PL��@�邨��{P/��У����q�Ȉ�p��`S��Ụ���j���:x���e�5*k,�r�t#o�i���q �-���ߎ᧸�_?���s�h�~��oɇO�_&<뎔)��F���SOpK�#�W
  G��B�ǡ3�&�����,yEºAD�����ω��|���������\#L�G�X�KI���z�-R7'ug�އ6�	H��^�򤾞�),�u�>�ԹLh�F��W��;Ho���(�i":u��|,�fǭ�� .�񺍅R���"5}v*���ض��Bz��e�0�g���z3ڛ|�(fju#�Q�~~{C�տG���gc\�-�Q��10�����2̰�y#O!l��!���\����
���ǅW��R����F�s��4Kw"���$P��*��n���@Ȧ���F
�c�>��R{�H�Փ\Zq5��zh�aVͪ�:±⣿��x�L��ѧXkj2U�uc��!�G��
X&��+��Ő�$CE�e���=O���E�S��b/aa�h�=H\��\��P�J;�z�a�?���7��Kz�ql��U������U�6HQ91��1 3��������);��k0���ѿ$[p���Jz���$�T�˻�����U�R�&�-�3|s/�%�St]F֥� ��o&��YA��)��,��l�ΙU1%�pN!0���_]��uO(��r�Ѳ�j)i�f�*G�h~}>6ζ��F?شQ�sR!�M��,L�Fv� >?����%f#�h�j����Z4_a����
�g��7?XR��J��F�����/�vL���^��7�~�F���*�"��(BF�A�^\�N2�ldl�s�r(�T+���d
c�7/`ũs���WF-U@K��ҽ�m�[�Te"�E��b��:q�*��� ��	���e�R��t`U��PO��#yWś�ycA��� �7�@z�j�;0L��ù�Lx�q-����i��k�⩀�Uٓ���N�	�G�[yDσb���dxX��|!�a��A�#��A�G,u�y}�6vϩM�D�9�U�x��������.��ٹ�Ip���!����.��r��a��#(�A���V���6�)>.�wdCs�"MO_�3@��n2��i��("�xgWM�TȄ�)�ˊ�nύ���Z�O�+#�'Yf��t�OL�W����[���6L&x����T�OY�ȷ�i2]��t\�Z'�[�g=( ����1��`� �h��p�V��|��g�^�������|�p0D�j����a���[�`�^B���I��b��إw|�e��v��r?^ev ���)L�W��X�e�kɟ���!�|g�m�<��M�Ee���$��_����u���ɋ�o��3X�II��tgd73)l�q���9(꘢�^�����0c��i<��7�A�,��>9��7d��z�fW�����-�j 9X�	��U�gxW	=w�F�P��<g��Iw�wɌ 
����6�S�.�E+JG��w��0,%w;˛84�Ӆ��3�|Ԧd�4�c7��Va�S=%��v'�ϘV�&�ׯg���b���i���w�ac'�'�����bf�>M�kE�Pռح�x/��ظhڧ�0��Rj�@[~��l�R0��� a4�V�;���TcSUV�M%�K����٠\�Z,���Q���P��'i��#e��-W�ŀ��Ա������L*Ⓕ�O���9a޴�V��ˏ�v�'#|Ztv]嚒V�/8P	q��uU��t1Nӝ2ҡ�a�vD
�	k��V�kB%�)�	�1(��Zբz/b��Ŵ�'��;^�-�d���K�����sx�����/Ag+%�,������BqC� ��H+���ɺ o�M����ł�ZC��ƭ�|<���14��.�"�����K��-�Ȩ�.�!��[x��N�쨔��9m��$�ơB�-���,�c��m%���aB��n�Ŷ�}V�XY�W�ꐲ�v�����y�^+��3#��S}(v2�K��w��ƀ�&�y�I�Mֈe�p��B�t�Svi�A��dEvW��o�|�l?�������s�������gO���j�Ԟ��>��r�J��p��!�_�j�&g7'��� $����޶�5��,��$��ֲ�ց&Gwv.�y��d8M����'K�L�S~��,�{n�@�p�0ԉ�Ek�c5��z|J!%J��@`����r��YF��`�Q_SySl�=���Z����2���R�y��#si��zy0Nq�<�c���z�c�$���5��M-�hw�i?��y��:ޫU1�h�r�9�1 Ȯa�'�[Å$�E�8��<�)��5t�������Ew\#����)U��}L9�U�"�����ڌ�)]�Ĝ���گc��AJ:�ډa!l���]^�'ʘV)���6�*ѵ
���ں/;�����प2�Io��]��_Xˤ�������m��h{��Bm/r��m�|�%C�"Ϛ�@+ª��4�h�=nw�b$o��a,�c9���̿�����k����@��K�|[��Hc�Ƿ�����r9_p�"���U��m� ������}۔W��1��O����I�F���hm�M�Y�}\��߱�S�i���ޞ{ٮ�wo~f*�%yŀ5x�k 0@�g$N�מ�F��*S���!��2^��%�3ro���I�KN2Ӣ�J�R-'�&55���_t���D�0/��w~���mSה�E�\N�0���#�^=.�o9�feL��֗�| P*R����#QI�뇅�.�R8`!୊�\��rz�G? j$�z2��`�7 ^��F�G��ٹdy��g�M�jsY�G��L'��?"�D�P)�-j��+�ҭf ��_���2��n4��g!�C�����[�"��H�W�z{���ݡQ�+��5������C����3�����J�}�����#(���aMÎ�NFij΃�SIT�p�C��Ҿ�0cP�&n��pj�8�6�22���X��o��r��m�r�m(���	�3��� ����{,�K�� �6��SS� ��g��l�������n�i�UWZ��K9�����"�"��� �`�-�c<���Ⳋ;
����`�[[�eO����'U(���~��(����r^� ���j,3���<�A�.V<����9����1�%��-���
��(��k㰩>�ζ�:���s�饭���N��+3q�<_>_;��?;o�W���M��`�-�0��m�#4���fLG	X���;�����\�
�''�ȣ} *���ͽ/�U��F�u���0�c�JW�F]����I3��$��}��vt�HT�&9�/�h/��qWn~���.s6D{�a_M�tH��W���=|&�d��%0D�K�s�ޖb��}{t���SK8{� x'E�J��z�Lty�f5�h{Kl_-�� a(S�0��孑؝3�i�Q��	g�,+'���*�*41�L*��W��k�;��\�z����|K5�� Yd�e��?��
���=W�SiK����� [E��ġGsoF5J�.��L�T�?�<H��5hz	S�B@�Tm �.#4G>�WC"�"��������B�j�����HD�^Ir�]�ძP!��W��q�� Q� P���K��w�il������(j��
xOz�.Q������؏�+mز�q��)cWb[����},�ܟ~���%�nk��s�P�l�K�c�| mO��imf�������3kz ���+-�u�;���%��rt��U�NX�����{�g���r���G�Y�!=�7�3��=��)w�������d'ӛ��?�,K��g��:�KK���?�	���ʚ�5#�9d�G�_vP
�-^�P�"|�,b���c�)g��L��A�ţM�v��LzS�
�>�jX�=��Wɯ��$��s�`8��YA��/���/%�$Q�}��̞ɶ�����Y�#�����:�����-(F�/�y(,�ؕ1.]�X`��RWqwNRZ��:� �Y�hU��\��Os�ٟۢ^�n-#�=}��gs�1rw��}������V��:�X�xO��(X �K����P�
����08� "��-�*�#��_����������A�FQq�w�Q)$���(��$�*2�뵷��>ݶ-A�P���C���J���<�ڱ-�rɷh\?_�p2F��;�4�`�F���y����	eD{EKK��j.eo��pr ��W�z	y{���U���&M*�9��elx�D�����D#����4�ݞ�3����(�_}3�2U�5^ʷ�g��
�$��ia���äU�Xt.�]�6��\DN��f�W��J9<�y�l���k-�}ªvx$��g�IpX���AA�-��/��K�g�ư�-��e�K�\b{���CO�
Fy:�h�P�X���E�/S#d��OYP1��Ј�V�!e���U�=-��A�-����ε/9�)a������_��J��ʹ�Ur��0t��������2�e��΃����+%���y�DV�]�����yVs�/:h�|G��S@@��d��(�E��iPh�[u+p��"��Q3�����\̇�]�!�eyG9R�9b�(;a#�$P�u��E�w@sHN����)�yR�C>Hw�`њ���+'��3�e�3q1�ϡ�L$c/Kz�JW��P4D�p e������o���(��=��sM����-T��BF����ȡ�1����ь�E�j�U:��b��H�G��ʱgG0�f]��Ұ^1��>^���zjk��M�����i� XT��2߶ၛP,Y2Q����26'AЍ��>������^��'������s��`�0*��P>%�W?��Ğ�s�:f`%4���2����<a]jX��\ d��:�@��&h����_��KF�[dU9;�A��Q��i-8�
 T�:�E��6�4��t�|فz1�|����<��+U�X�u@�K����n2v�&,f~��3#o�B[Goc¾��gqKw�I��."����x�;n?�v�E�{m�ٲG��$RZo�Cv1꧙��罋����눁G�bd���BmWn�/�ӛ�xO���J;3?|?$Ѵ�������տ�������~<=)�H>l���6!A��w�X��%.U�f[�[;ZL��onY7"�*�6�Rz��h	��=H�Am����,B�)E;�q�h}X�\c�'z|��+C��%�Kd�/��@��c��Y���m�a/���Tk�ZB;3��:	L����؎���F�C�� �q|�A�j��/.-
t�ƮG�쓗��=�~�i6#K�x,��$�6����6�8^�tb��~S-����ٻ��թ$��z�A��_W����?��Rp�XPf�ەz��&�YQ��p��Т����:d,��N{b�%�5)2���Vz��v> ���9[���A�� �8h+��x%̸n���>�A��[��r�Ƽ�NQ���(���&k��8@���}]+�S��%6v��r�,1wI��ώf�H�"�/k0dg^J�~��]�&���\R�Mx�d��*�� �f�8�r#B�5�Z*N�U��r����gjj���"M��=�	7�=�q�#�4�!1�z-�0G��Q�5K$�~e� �{��\���N7���x!�=��Xd4!	9���8E�<�ux�z�r���õzV�
:���������lf$@���N˧�t�+�>�2�q̓LSk�o�z��]�r37Y�J�$H�D�3��UP7�9��u��y���Rs8��� #�gh�-O��������˭�9 ����8��[�ɤ�c��\٬봑���jF���5H8�Eu?!9m�^��y9�iLN�C]t�6i� �/j�ڗ�?�/å9s$#�|�����[)��6ꭊ�5�]#� �m�E؏A����a��,$e���ߛ��$�^�$ J4e(�1�Bv�X��&�Rh�g�l�FR�X���JL��&ޅQ�ro�ب�dZ�z���Kz{bhtK^J9,hw��Hc ���o8b_3���;�kb+Z�T�Zn��L��([?�.CIf�w���*�
Y�ZA
��Y��:�9��ON�/À%�