`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
GZSIT57VbdhZW8bu9tgKtPMEgHkacGevyfg4c8WOYSDyvqrahxYlbdYAikuo/lbRhQkd9megcSMX
vznrBdQfa0jQRjmtryGhvhsqFbNFZIkLRjGKVTbn0OVBj0bNDI810QBzhQ0y1AI4Kw1/NE03jANE
aX3VvoWK7TOIv0PfeI9wxJ/7VPv4MvS8PLmOmHU4Vpn4FQfVu4OzoItzw0Aui0O+hpU+UazfQe5Q
3j9QHJU1UZyhj2XinaHob0bbXTBqtFYZK6RWh0VNgSlRwesePnBKbBfCONDmItc/AYorc+E2XpzK
p54utHoy2FExnzEAKODBSnJijYd3CPMLcYRtvA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="vRCHPD2HZOOlafsmJImLL+MY/tQRQJdsLttiVriTzY4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11808)
`protect data_block
UupeHz4ZUjC62MIQPn9ioGc7WANlpbJ4DQh5VyTitSA5REGxpsxWMKUqV+FterImHvFKZTJ7B2eR
LG+tg3vczCa+4w/8jpl4KicQbc13oHlrx2h3qrL19xNTf2CUzlcS0FJ/d4fmX3g0L1JPKYVnXaFW
38E18qJx1su3LV1qy0b8B6H323sHdqGSHFlATxu54huDWeb4gS5QCVm8pf1F83/fWLwf2cFYFFly
OtbXfsg3IZDTKNfxCobxkZCpjkzA6hhFeuqGV76VS7PoQcBp1JsgqREaUmUD9uOucG9GJ3qf01qP
PgQ4l7c2w6qyZf4rn3dl5Wfiw2JOBnvmFTZAeTf84Z0R19jISHfPZdgu2uJBg9uErmA1vzxnxsFK
Ga7HM1vVVtle9ZHIU3Q4kI2DsuPQpgWt4bbqLPR1Ka8JkMPBhmkXdnsV7STROQ4B1Spoe6P+rmVG
WIBFuszzSBxQw1DYLbZQrK1o1OkcwiLGm7k6s7p99sKH9t0plqZiS4NJHX04D9hhAjINruM8lkmd
p7YXEX8vJCmNmXRis7GA7IQ/QdrfMFK5jafi5lw2sU7FxRwcZj3qpOAgXhupy1iAgjG3QwL+oyaM
HR4PJnzM8CS47heabtVe6zvb5WszH7lZdg5eNZE/dNqIolIpoHggWoNBAyF4mCOL2dbAjFtCtcCe
QDnajN28azTzwqt7GLGUjNqEx+6cghOhyuk7NFrFlNFEIWERbFgcTKjfjhhXqcs9jFelX40DGwzG
wehzDiIwVCGvGFWrAA8o0Hxiplawz4pdvgEZDRMQBsCxMVCEWUBQy4YLcvuqtTvPzY52fAMDgvCM
1qiT+/GeQjsEHBRaO5AVfXzN9sD2ZHjd7lN36zDzvZ2g0bDEjZvk996TFoai7lucklpam3Y0/UDs
Y1kxZpq/cfG/n4I/l+cqm/+Ia+xT/CYhAVlhRozSwasSzY6V+WgqSO3RlFYIIh5Fyf3c88GFiFTy
peWdCSNeJqGstrmmywKfQM0JoENfjWMswaAtrhXoFVUw6E6yljoGfHway34piqu+IhyKPxxIQ7fy
Vn1zJ7Ap37hpHVQjdmlnAsmd9q0p4bGHl7ZJdHfTvzBRS7CI9cXlEp9tRdVja5GFls1/jZnCBBvK
KZ/btFYAdLT4Ptrxi7DBQlk5XxGVHTtkqTInFHdT+GFXw/JqaggbYPwI15DZzxeJ3l0jsOqqH826
taK7jNou8sf+Ox8ovdI88J6VoIWjVLlodGvht5ccngofL6PXf6Bwwc6lA4mt7o0p3S/OnImdVv+K
Uvk1WLtzv/7qtp6l2q7WAo+BD+zkXZEfwfQ6hXsjVLvXTEsXvPt+GU42oQ4iHJcI++mwakOzVm06
KbTRYpxA/hAYQPlVyfDD4jPKuYGOrhMkPNQCakLtIaJ5+/a3/f99x1buq6Dl1r8ryQZYURzU2m+Z
RdWpTXqiJ77djZWGGafxQ9li8ChI/TxEIC3MxxlzADx+8T71/GWUo3H0Gsbw8TVoCiOlIRPms749
iu2MW8KDWV+lKf7d47kpj3rPf2Pr29smU4xX+px/QI0YlPfRbHUhqifs8k7j7+/356SkTAqW90eT
b5j16Q3cDTmcRRR6yjtTM8d8Mr8dYweVGnnfB0O2a99t+zhSilxWnNbOWjmb5xvJ+Tqm9PYDuUNB
vbGrbcKwUBBtICxJkTdRFNAHMJQPoKucYBhs6GgyeY05w/bePNS7yDsqo6JFH2nJjXdk/CzYKo2W
H4ZtDlRVp8QnBksJPu6GET6oUGzu6WhKJaieLt6qc0AiuxErJBJVmq/fhhip7/qOAD5w/jVdZOuJ
O1Fqf8/VUNv7I9OHviC/U7z+GpQ63tkVFpjKwLGznx7bJPizcKNB78PX8ASMdaaB2LqsKbWcaQK4
s9njExd67zC2jEmL4HAuGDmQiFcqKZQ1YAO2iVU43DR2qn8fniaUE3yHLgpcKIznVL2+71kJ5bx9
Ws8BvYic3PJnKWG7HXUafe50v1Mr9Gigv2i6B1ZHwpYfFkWXCyyfZX7Hvh2LijXjOzPGL2Xe//N+
l6XGQec3kRVqxbd6ShtX6JtJLbLK4S7YPHl1g+Lp//tTGFGl6H0mYFdiXXKky6yYGlx3PgDVCySg
1lpXmNVb+KOwp2qCOl435btSwuxCBA2nCrUg94SVbqsHPfItOEyr1xcjHI/v+N4/dUpdmIh3Tlvr
dh08m/1mhs5sTZlMUiwOOzaFknjKUqAwRJWvCFKaBS92IBRmDJOY2DNDj0CSvwqlIibAy+pgPhp/
a+mRMfOmVT8gHZ1HqUd6TwQmaQKsmD/aD/Ln1AzOn4BMBtM5ul3FU/XQ+phQQurN81TloGjFxy8l
5bIKd6668WvBsshnHZzbxHxpjrJSNYQ2t1O77DTUgtKCGZs6rQkCexSpkpjX+x9CHTGYZuB4Sl18
UWuod4cN86AP4rrhZVBEU/cbSwrNkEXxp9m8bUUp6M1TN/A4ST3Yh6Ulx9IiDS/u2jOpjV9ja2Xt
r3fnbW0pZmvBa0DPR6NodOJNeKpc0LDbEI1DEAA9G8in5AAUTvX+LLc+paS2+B8N20dCkHYeFnS2
NTH/Ulm/Jwas/d985/oGzxDmrfbBNJsGm/3+v1wSh0X8A8o8n9zU1oLSmBh6lizPbmfhE7h6c9eb
Bqc4OS9yS+dvAfNHM6CJxivAXcoh9KV+pXM/RG5Ykmqzn8evl7Hh+5YA7e/jjKhhagU2+/JPbCzp
D+hBfUithfr2dZ7Pq0JZkHiMaKHwLh+aoh64hsS7kllc+Fko3MuVzAuVKZb5BnwsSqI/HV1D3AgQ
Y3zlNYVdi67MI+RtQctczPfOg7nIQXRPTcnuUJPKWlwbuMMLh4VGHSy3pFO5efEwvIjX3P9rsCVT
KH0Bj2PpsWlRp/chs1Z0vDY+dzP6zp1rKaYgQba/Xap/QNCbXG9RZrkNEs9eoQypo+1SerMNOuV7
mq+QSHMVaLmz8CqAxMJO5torbHFylDoN51TYZMIMgbWyDbjy0D42tFrx3wFsjUlQ0VmMWFCQ0jvW
leUjtDDHPjYyJWRajn4AZdd0j/16LZEvsoUExVBIH1DDADwiRMpUok78a+bl1MledSmAGuL7kVHm
umPexoE5djjrdgdagdqA6dC0kNuRAUCoWQaVw2ghzc9EI/4sT45wYAVgCI9XX/0NYflLZi6PeVfm
2oOOKmY55bYdZ+OnLA1uSNQhHZxsKDJtHc5UroGltDSvCdWibNu9A9lyj8G/fPpjkPICubhOcpVq
MA/fgHdjDL922qeUIWaOZjEeYD036/4I9MJq4srZ03l3jM7O6aigI83tjYEYj3/IagF7LU/jPIg0
a3UTAoWkZqT4Wnd5c58FUCBBM8s6QHWCMD5mIz/fmAPbV+bwUTdPVz/WfqUGVGe81BVSp+RSvkLf
ZEUJP3LtqNowRz1Bvja+2F7IZUB3DFl5jM1zz91HhJfvZzcs2GJrqFr0vaj8sq+CUGGC2GTkcMrI
/MiJbSY4o5mJeQU+yp25T+nmi85Jay5NpE4rNHnWkT22rUXYI2fFhw6mLdphSzt0sVPoS+bdBlvF
MkCkTtfeQWDCpQBVpv/Ec4zVPyznCp63BADuIiTDQZHYJhK9NolSQurC0L0G7LrzxRPVeobWDoMm
8ILubki8Rj6U9PmAj+nxKRnG+ZVC66QGyWP05xqK3AQX+1erASzyLb/VSZHeojJ4a5T9OdTS7NYW
KTFKrkWjDL+zKcgDiy2+2E05KIRWn2rIG21xKtB1lQbRXXfca9mcR0sAUeRw0uj28O7cqFYe8gms
N+tx4kxazvpB+oJeV/cv2a3UgptQq6TKwRP//NrMuB4ydvQxJb1QVI67muwFDYdZlWtzqj6+cZ8Y
pBzTQgcptLugU7Cch+d34oWZ9zkkW7zlCpkzT+T0Pf4XXWuDsa64nzoz5AsRQfBVYPmH+kS2Wriw
M7thA1mhQTSCrPr1E3u5dXnFlq+RkXSlurjK+t9oBBlyXGeNW1x2oBqqmY8JkvwpzhYNDIDtliIZ
o/dte/nkNbybMHPqe9qhmYCQ9cFUgesYSuEEZhxOvMN9T9WvnjOzHDR3RK14WxC/ScrN6U928SAy
t6tXzhY/ARqhdlAzU/QDO7yldFMrAb4TzxWybbKkp8WTGEUN/7X0yiZDRlJyLh5wZS/FQgPxcvCf
h0FaXGHFUxOj4Fns8XHN6LEBmSTrh/rqtURxS8bOtBmtgH1pF3dLbcaK/oz8jTgHPcxaMN1HBVfY
Te5RcwRfjL3ls6b+dLFKoTgg+2zMW8tmmFO6w7934V86KIUyp7f7hUv1z+J9Bpx3oKl6Uj0TvJfV
SxpJmE6tBLlXalQLfMzMxS1lEvQzgKCer/+1vbtW0J519etZvCW4f/UJ1XkFPsTd0tSAgX9JAjGl
PpGVJ5wGuTK+o4zUxxQHaaPSufvKv3eoTFMYGY/2J9xmccmxHRupv2/X8XC9i7VPe4ij532ahXVs
cWWJb2A4neSIgjKB+V2N2JTLHwkbUcq5dJ5OE6odUVxxiMSmvQ0QJkkd3lACvFhV1Tx6fK7+qbGs
66oLOqidFiiUdPy28WOKLIoYzK/ES1AnPPZSZWjteM6eakpIRqGdN6/xXbBzExD/fnLSI6ZLjAAR
Xly3qdXTIP8Sx331cChym4OMaTHb5AVVPhfMSt5NEoKY+5dp+9J/hjQcrqWz4vjDqBiBz+WyMXf9
o19IXeU4WZtVb183HTrSkCfewchgxpovyvBRl4Hs84qMxG8cyv/7/efFfXn/K4ske3jANRtGrde7
W3mDyXOQsmlPYVeTkGlJfvwsSHstov7/3KTfxO9iKNPMvDjmaeQkOkVGzQG9Kh/poZpanQ/XgiIo
GQKTHajcxtHdsjVUmgAGLcwoR7O8Ma/Hv29O3zGRhR5Hj9PeORrFQPC+oEHD+2feEqwS4XzPI5yd
PCo52m2ImRhqpxYrOLZPVjqcSgREav1urCCA4TLMLgFLaEUvpy38YDwdSj58GIsfvl3jnMsuBF5A
R0DUQiw7s04/RaEgXI9qj4n5aFQ0Vslb4D8W5ob1jkZSF/R5YGaSVBJPJf5gp6TUnc/XgYW4QpZM
3D2ZGjnTWOgbrQ7S1tqcvssSJLTMS+vl67zF86HJX8SMHahKJpOKe0Cg2vdL1noGXRlpTrJiq0z2
9uWoFE8H2iYetPmI+aYVJsUSr4iVvn73ij0pCkFqCCdroVO49UGvavmQh2JkIOzBOsPhs71ZoloA
EE89LxY8gK1HUyk+x2RiUIabFoIM6QPSrhwkNPbmv31yPprfcslWf9sKdA4eMy5tRdTiIIi47kst
3nQFyWNwg/ae7KjPFkO6G5zCt/DR4OSXSSXDPfEGBZy2cOSSCnxrnUJiV+NMkgxJ3W/s1FVrpaHV
ixZqpGk+dPf5hDqB8uQQTW08EN4Rp7cw8zBTrj2lg4aeVdnPaKZVmZWiv9Sr8aBuJO8pnKVZeeXp
rhXppddaQ0cPgXhMrQEdt8SjnuucE8dDJGuyPtHswT5kom8bZbuRBtzo+c0QJR7BvWuW/sarNirY
qgif26OmfIuXJ/UTUTq93DVHP0IJZe85iyjE0cWbrVfGd1IfKqzy479e0bYbTqozq3L/olHB4LAS
o90YN2j3Apj6rlUPsr6FefD8YSOBY6M3k2flLOyQjjzAB+6E1V2F1Zoa7LbZznA0kNisLw1ryaAh
j8TtCW5p0Z4sWyp36cgjiTlXMEiBdTmQnwvXDFuRioXBY7f+NXvcTmubYjq473doxqsKlobgfN28
fim8iFWAOi0kyJZC737KY+g45IxhFWn5BVNP9G37Tg4rNFnffM2espIgr/HMptHBJtDs2za/Q1o+
wahKZg9xoEjiRPDwBHodvPQWI0QJhMryclrCsnZh1lQ2NkL2TE5OSdY2xrCN/Hd6BCTP7A6GRoh6
X3ynu5wIaCZ/ZZqL7ghkjzXzz/qepRmY4LeSfoHpQUPWuoHQCMepaWQoCXGn4GRPfIvdOwJL/Rql
DsvgUZbfVdBgqtibLnlWDmQdCB5m9yWDbhykoAHeCchhVZh2L4VinDb8ZfEQ9ZPyyHTdeUveKf9E
gSVbhpBd6vhrHHhCQAMVo5k1hzcwBlOYnlZishdXq4YkR6WaFD9bs13Cxsoeu4Zm+8FwsoXScrxs
ELR/E4p/AUPIiyrZtZYBWXJDmA9bVv6BILiFs7no58HLwCo/+asU1EU+ByvBPF89bUx0Jabk4V74
nr8ZNcJa5iqWk7Cx59x9JZKMFmImxIK3Czvj5g8135wdEAmk8dHQN4lw931sNvwTk0+GrdBRYSfI
5a2+uzZEakUIAX8uWGyM1MtZHaso4bkch9ZZ69lbmRBEAjPKUyMQqpb1lxXu1wLOYjXSmAP+vQVR
IRTh0NtUf/IbxZPuYKtiyw3Gkz0tTouJbmsHjWeyMAVq0PwgPrgF6Wvv2ZQSUSM6aY3I+Z8jIRnM
Qz1b5QwHlSSSL35sQK+wD2CZqO5c4CraqzZao/6oqdzeA7pWoins1HG+W+0jSMCtG2OCL0lNtBVW
6cWI8j6WV+xrMUi0uMG66uchP7gyrp02bSYnNj2kfrDh3f/jA788mNK+VkO8UDBE925i065M0hnF
zT/VrhDyDtc5mTFQ9KGznGmHeh5rjNq0K5Wp9C8ZakR4sj+IKIbAtvCCdgFxAJ0o446b+VNqv4xg
a/WrKZn+1KDY3V6+SB7HW5y+TomFohcTcfGeyJJX0iqgL18eqpRQ5j8Nsls01BV6tM9Abh+QquL7
RKC648ZqVIAVbxLIrVC20q2p1Jg3dE90SRNg4Iga+2w1a/dsEuK6BjmSk9KKxyZSN4McOlfDzBbS
nM1h5bbTkGDF9gRgn9PaMbjpVMVI9q/bJjM0Po+/fIZpNOo1NUwVx3zRImoJEPGojO0oiLtZxpl2
0zjEh2caBv3ScenKEKEix5eo0ip7pnbhVFR5QL67e9Wb8fLetp9hZ8pZgb6Z4ZY9kf7Ax8k77oqh
YkWbCAdpQD6y2qT+YXaLRy9qKd5F/yV2u/8FXDfGWd62C65xoWSBPhEDrhAjo2I0kvr8bT2kvKpr
3gpBGWNLfKJMdihG9+JSBGkwnqqK0f+05x7rwGFDvNgnqDY8ih8UZP2+ekEd9fOnAOPQnhb1kVTf
Su8QibS8aNKWrpGweurmfle05WB3NCIzZZX4qpQEpM+VIYDQt4p1lrCeJs7/5a183y57whTqwFhx
Qp5/OUGP/nQqWB6TOScIjA11hZ6VAtdbmQ72vpKIa8IVGvZSvaa0o/OMOCuXfc7vINZhvtZEWZpD
MwbhvkyFKVbk2ZtYj6OwAenZEFiAIJjuf36L0DZ5hs0eYp/YeJXGC7za9DUC20v2xu7E+NA23M0j
O8SB4xkRI8R9jFrZNIxC0odBCNE80cQ9E+SyvohkC/zToNJVCqsRhaQRC/Ry1Cn6q4r2/CodKlii
zzIeoRyMSwsOVXfMJWq7Bd0IE/1Fn78lE5LaZNbeNP4oZU6H/5BesdNUpKIu3V0Nd38ai1f4uLHU
jsIFNEplnXNT9n6msZN+30LfugMCHPcf5rthELcb+jaHGFSWXEgaHYxhrv6pTNCoGt5Rfhd54Ooa
g5zTQ6ILgdzQFIBi5GwkeRk7dgLu0wasD3KYFB0hm+fqM8Cutd+AfGnOTPDpbJkTGa92GJoE85vT
2iJZXTAwv3g6hVA7RdOKEURWP9fBIjD9nZyQTRT03hua8mspYz+MXPPwtyWjgDEQZOW9F17PfBcY
VB8joMfFwkdPyHIGiBnRS7j8mu2AfiQwprXmBj51SkoPrQQSR/yWd2O0xyBoHa1I3l8a2gUahUa3
+EDOZXyod4Gobcg8acdbsy1inFOJvBYhq7C9gDSxDv8G1ZFxMqJ+y2y5o/WmR2KyccBxV054m1XA
PIhM9gRggVgylQsZy1e1S6fDLCbw8pJ1M8t/1LsjLpeGvulUz6GofqaaJ6h37x/hOfAanjV2sXoj
Z6OeGVxDPYJRjT97O2JcLj6N8+Fnmc18ejULlcqqA9oum+E0Ra1/E7HMpuZj34H74hX11teerwKs
pFYd7auuiO2GNnFxzx/7F7M1S1rAf8YXrS/EIIPEaFN2tZRenY845pljobpWrKET21YKkcnPEhOk
fBpZE6Sf3DRMxSOyxN/0ijSCidfyhLU+XwDaf1tHqqmA+Cqlc6QOuQX1McUVllomjgNyMWlHQtk+
oNAbd9AYZZzZ7ldBLOijNZ3q4/VbOhaHCNyfTGO+cNXZtVBdvRCfLj2pwQJ3AnhcrsfN3z1Ielnk
Zc5ld+mvS4nYrgU3ckCZ4eVwHYlmYN7xYogWmSV3pfkMGE6/r49k0TTE+NJFNTwrh1zyb3nG9a1d
WWolUmpdCBq6qnz/85hzM8Ot4Rtu6s+vRXJ97vGR3EtvUMuTKXDr5Nu8MpfAg3NALEzAfZPGX3bC
Nj+i1f+lqQm9d87w0xMlAHkLNdD0mbFwLbZTsrO6pVbZsAKfTnY015gaHFKdEAWjsu7z7/WLjLvx
0JSdvoPH+pRLUXqBL83BpEwCCrcrjcalN9iqYcCMNPtu6Dpg+ATe/Y6wRvBOhoxmr9K4gabxRO4Y
aALYN+NNx3QQkBzqeKPi/qgGNWR/02XN+8t6GPyWrpkmECVgK5lGvv75LwXW7x3O1tI+YedtRwDL
ZgAaNqasAkhtOjA2nOARCBldrlh7R1JSf7EEOp+/ip2MZmnDl71D+qJtHy2FjF3Vl+Fa2/tU3OJY
ms4oBIlL01SHDCKve1eOAScsBfWwJFst2yvpdZKHsDoaP7shrvYhXHN4G4bEhXLg5DmIDrF6gKY5
oH0WpbSd3H/weXjhIxSDx9ef/rLiYnXWcRt6SRMd90sU5A0AaDRVapbJq+PxuC7Syhkfe4/wxWOP
UuFvb3JPQ2PKjwvLNLYVI6unVDqpFdjoYxoE8iy8BvxYmGpz+27waCvmF4HmBRgaoqtd6EGP4XRV
22MyepAYry7WsI1Zhgyz3SjLhVrgw7wA/qLB1ihM22eMIzgAcl6aSwVjXVKNJ6/NN6JzSPNwnV06
H1Ag19xHzs+m8uJK+ETTLNVpOu6qDVsB9FyvTwLwTJf8QzeqasVKdW79SoN8xjlzzNmuEWc59pzs
v1RgvcX82ApmmkGUy6aEAAzKsbsf32JbmsxwR4DLNSXQQZXL8tmOIqRWZMnaBfrpkkgHC764bwR/
EUNmWun+Xy0iPb64ZFzKUY7LlXZfQDqzKLkS4exQ7q5PLNSrHcRLnaK8y1fDHM13Y2toGxIoPX/X
Qo7/bSSLl02DJVK1zo36Syt/FJ8wVdjcEZbQsq72DmpFGwxNR/vGEVXzm7zSUYqAoyz9aaPZefhF
RtV0J7HL7J6JL9JxHDTf9saK8MzglfEebF5pPqlDRyYqcTJFdukS4YImVZZ4Zm45j0sKPnIW0FVQ
zHrkkW+0oi1Ch+nvtOSd717tJhSCmJUIv6iUHnyturq6DcPa8KrzhCoOfXfflTe7RGaXQVEE+IHd
J3cBp0+npLR6h9gq4n3Fakatw7AicHgC6G1bedyjnXaZyc+4c6DsvtSATZckY9LygvTIeUJEwdZ8
P4IUbnZ1wk5IHjh6Y0noQlP+Nt+ELk02oq+6UJol87F5j1Ao8sH10xOOjMl3o9Hk7o0etI+X649a
Q4F/euamjAqfnwS4ezXpW7SutNXMOMZ7Tg3fOaof9NCgiN4zrXO2FdybTB2XjSbIKMb0ZdSFE45e
a090RjNHHMkqLFPWa/Dpc2vVCUnLsP0cVk2xll19tLwTZviT/EzG6Ubb/QpHSLUNpWeA2YQb6KKf
uGIesplmZ9de/qdxkcbjhaPtHsu9ACMoQROAMV/a1E2tQ+JGzTABpZ2piHn100J4lgywhuTre2N9
5k50a3EgK4AkytYpcLi8jWJAlN0eL9PoJtJ5/u3+hMZW9ETkIEHNDG7xeh4+/7c/2ZEE7AwMzbGh
t1Ez1kGYDPr2cTPHTtfg95Y9WqI5Mk+VxT2etRR4pGzP5wDq2lUiRtYHBzxneUbvMpha9BKdOa/w
TRnfyd1AjFeyCeLyh5AMLrafurkPPlVIPk3oywBUJrCbd7d6C3UjObIMDjLK3oW0Dsgy1uTxtDIc
LbitKM5XNSwkj5SV3TjJYe6eX1Xt2ubkq4YD78GT2mYjW39b9C4L9kQWSkXyWFjcgKaGzYiKFq6T
PRWKVUpjR3RNcJSACwrIhfeOE6V+gTwATKEhJwJs6hsfjcEjC2IbiZmKGsbwyVo7Cx+FXh/DahNJ
AsY1cxvy/JIuPK2DtBttsdTqKJQWwlxYS3/g/ZaNrUXBwWzbp2rIggG3Jo9S+NHxFCn/uTK/pH41
OcpSBhsknMJkDih4CWpnBfmY6OmzsHFog/TSyecCBpxTNEiWhEYeCmbu2rkSgGu6D+GugdEpCi1l
6pWbFuxicZusQMeXJJccAlsrVXUiaY9o6k+QQ2NWeuex07hatBE08YbPf/rKQb1GKxQ/M1qd8fNX
VwhdoblYxAUHlF4lf4h9TeFob0NiRM25QCBaPXPm0cycOZGPNIyqquG4Vo4Pbz3zg+FOx/oyQxzE
eEejlPz1CyWsViqiHmp3ozkWLUDgLhvzxIT4qPsmwO7WBTDXgWAeOQAjVlxd+iasZhoItUveB6nB
3XQ8aaeU1wnRc00V3P8SZgb+KriEkpDGT6HKoAzkAhfPCEXwEWkR1yUssr40WKduS6E0uGCisvWI
zJ5jidR14E+Bdf5D5tqMl3U2KKuCxOWuotOjV9SQOk33mtKjFj5i8E0i0RUeWjO3SbsiCHB+aBLH
wZwfnoejc6P128X7HlV/HQF6M+WmZrei8w4spHy7ojZBF6ySZeT9hQWVGmWaCDB80v1vXM0QuBqi
Rd+MR7JKE21qLY03ixQkWFluwo2paVIQJWecX1eGVTtdKR1ntydSkZdlSH3cu8zN2HTeNqo4nKFd
c+HIxow54dOjrYvmB3y5tdzzAFMX7QJB+syB6wtz5mqpn/II9aHDS19Hrj8BjgiZiNPmi1gnklcD
FPk9iJUDntHHcS2tfwP6Ki/oy3ttSXZIot+M2X5haSAqiVV2IdICx1V7OICq8LuCaV2+dqK3J2FS
EOC///STb/YmeLGifekG7E/7zGCloe7bnivGsLQJmOCtePqa+I++L/4oQFnfJuZeVWpIf+2mKfAX
63WAqvM8PPAu82Gk+sE00ApTXwBhbogAdi/nKhHatyChEggrLKyrxqhxCgu78uGDuu2/HJclONkx
a6urcF0njTpEEoCp5gPcq6LFi1olIzt5qNoFDo5gz5jMzWAXUrf6Z3RuJ6Faeqc+06VmJLw/LFFi
/0ykVvlJTewWGsIhOX+vkeJXdOVmGbIbWp34JowMTD0waMBAq2f9/xWg6ax7UNK+170JD6cI0WDS
Hn5HgdEBEytwMifexiubygNY6Z0EdZy0dGBSC+SNIhZ/dcq/q+tfXu2+4syH/sfB4KIqRa6YfUh+
ca73znR/nwrGgGKM921HOOuNH5bjVrl5gzmHNMOxApo4wP86pOdDtKCIV39ZVtaPfHGqSQMbj+rl
ChF+O3xmbbAqpD6Ju6rBFrmQoN5f8L0GYwfCJNwaKDoLiCBJsKggQ1HvVjwRVLHgXmvahzi0uzv5
jh4pGquVQ3FNEBL8fGWXBO44Y1DdBv9xC2kJ/tRnu8wjpLQCkfFyyIN2cfc6vw8DMIfw56z3UUcE
3YQn9JROGnAnhN2QleZ7lxl+MQkSaXx4wLd6Vz917MNgSQ5z03t+Ll+3IixrNtxbsnhEMYoANgDO
CxCXjUK/AcjaYBi0hLkmYW2I6ZeNBlF/pfAOZCLWbMxdClSBJHhsFeDok0zHCmkCjtOiPHqXKiIH
NJj9X9bDbe0WHEvqMOD1bsy00IVsvxlb3rDTEot7nvrTwuOQHENNYzDKfxdEYWhZQi6H1ghsSrDl
odQ1QPyTodn9tLC3PtKFd1PvwSdGbnkel2xt2HYQNBcoX+5Z1kA5/KkNsiv+l41Dz8QRbuyUyezc
LtGu2MT4urgu9ZAPVS9zy8/YyNNSOH5j6BarQsTTkHTfKubNJDlyliw6xEH2u2OehfD7Di54c/og
JMw2Vhf3OGmmVz7nP7SUzviXcZ46Ps2JqX4IXxru8V5qq/gEamqt2MDyI3W7DjD6T8WvvPkNAR7E
WvjQEhztah4JkY5pfaWediVzSyp6riV+j5kLOLZG9hGyFWgWRDNxfO4glW7mPqJ9Zl5iInmLJg2k
G9/3l63TsG/l7/29KVUg6Sr4qAiBo1XhNJlYt9HaLhQFnO0yHEZ+rqgCW28UHhgaSjJ5GY20G8gF
UVuPHBtPdXlPZidvdGZPCtq8tKaC69Xn2Xrpp46rnPbSQukmIwPkSacJWhytMDMXsCuOFsLzzjAh
8aqrEdE9908DwR7vVW8UfFwkcQZY3esywFEm4U92uGIf8lCtymefMBe77Otvh7yg5dd9J9cL3z0e
Tztzx3/godNp2W3X6dLIQw+/YgJmrT5E5yrsE9fSjQazp6VzvsNSsbJToXOjmnwKpM/6No6nBeHQ
ZdT5FbiVJFgmaieHMDVevMs+yRQ2lUdni1BHkyb0B14pQid83zEzmUUDpOYiUkSH8unEBgFG/t+N
4oH5sVI6nyDSaS54OMiKA8m7I2sV39H3+fAPFoHCTeMIYaNpTXx4T06TDCaUYwdXTK1zB5EMb5Cq
cRQ/HJasUiGR4R4j56exMy/0Jw50AJw0/SO+Lx9zSqU6XHKWhxiN+zf/6OQVHY1zcNgqWJ/8Mkfw
ti++BqCxEs9YZMnHP/T6sXX/E8fJ8VLeGzICfgmB+M8saF9wUD9hUQJx/iJ4fKy8J49ntMjy11U0
6eyKTzZEDqz79J099iFmeRt/HkFVY8lgMl5ym5PGPdlHt+0+WrHfnklEaHPgnA4TLQKKhzfNzQ5L
43HbEQEl8RuQtShu4lpd8RExtBZiU2aMQLvJkPtraIaDizsKmRqqN0PykARRV1ETZwGlUBfKRikR
qLWxhCnE11MU4vU8V6wHx/8juEQ3lGTtVGUoag4IsX56tSQJ+h6irGIvzIreNjowWrauWIf7Bwdx
njGQ8AxE0GLP1uAWaL1QDxv5N/wYG/7h89UWOukqtvkOur3d2OAfqPblFORzgba08uIItLrqTRVA
wS4kY71BLb7plHaTPMxRg26Gntx9vsa7BaVnIRHL1GuFMTAG+sx3R9hJrO2LFsR/Z2XNzcuCR8FM
Gur983xlLAkkaJSrDMkRp5JuKQvhDa9wX8ySruIfeaHX6BKycJ7eQw6/2jlnGESIfr2b9BzSm+dk
A6fILo3qqyzXbav7bgbyNV3bJ/f9Asm8SguJawSKL+QA5tK1M36qKmTgFeCpx71VPJzWMC4LtZPI
17jkxmKwK649n3P3slJbmQwrJ3C6fWcEk3Ro0dfAfjXBGKY6m7C3juRJwDtwjWcwFm8A/LGXmgXc
80SUwl9iTMOljafnBZw/pmYkjRRT8yH46xX6+VgaLXos0WfmOYodm1TyhhUxutbOgJ5MRLIfyFn2
y9V1B4BusxqxXjkiBx9MRo7FmgB1jJ7p9qQwgNFcZrrh0hoSYvUIBJg6IAxYC6bvbmwb2ssb6Or0
CBGhKDq1/R/108R0U1CG6xuZcZ/lRW0J4rLI2Z38VHhvwk6MKBnRJKwR8kJwvVModEDsadMW1MXh
Bj34ntIhKekncu7UArUP2Z9V5oUclCAgYdL3lTiMLskiNSML4s6NSj6cRFF3BSZsX7PyCba87UXK
LSUArOUPzrfhh/eNRK/IK5162I1yffiZNd4icPCdGUQ9jCO6h+3rOl8FQEB8I2Su+X5+bkx5L2x/
UOyx0KweHzd2Z9lBWFk+vyx7GWq0TE2sa4I8qGfukxhQ1wksUe4Qizn+5yF4zV6RZ8j4QZsI1a5u
gxQn6aYfBOKwtrNLfhsodWlftKCliLs/t8Jpbzrdp9PeWsESCJT2J34Wnw1fPnlcrIC0o/vU9Tib
ppBVuG7R7y+ikTMl/ShAOQTJcB8AvR9oPGlK0etoQWgBC9mkAF9G/xqDHwVR1bQCQHVTmjygJYLD
YNqueF0uTc4xxwYfpGvnXCoYy9Us0jH2mw5mXxyF4rjTd/zDJmqPbFLwq7orkOExMBMbeg2qN42X
rojz9QNsMeLOj3N/EHz19/HMzJ8L1XqZOhD3j4zq5/rOWjB0ZnjwONaMF/ZzkvD82NAt9gCnxVta
zN7BOrrx2l1mNNgPNFCoey07XcmCDVcgGkytJkA7Bh9RiByQl0iK7xMMnxLnMoKfZUr2KPdP4EHs
xApEj3Rw6Kn1bdUTuRFf+pLqDzgRHbukibrK65UpkEP/Re0ErOKDVnZrTX6lyMVpd0rMPXjConal
nw1n5PRBIDMTiAgKliNo/RdEuf9mqwVisz/lW4M7c6DFUnDPacZcPwIDEffnSVqOUsON6gWMmw+x
PIxqtsc/5oLUTfc5oqgKB6iz0RHlirfm707SrkvMSRcpurNfluIAmVbzWx5lVSeyI7P3ymiYlnQ5
VDkwlpziXBUXBEz75eUYaa9iYrSxdwODhfMzMSg05xfQiUOGl7qRqqUbi68n9U32dSu4vlyqoOpi
Q4YWlgl23gkVBfQzCwvH7k56LbhlpBdYEbM4Srr/a3g5n2x1lmLRoHJlKKhxvmOoG8CynzFRYpci
pUz66cELhPW8qn2eqe76wz8Xz+/+DmYLsX/90mNQus+xeJFy41dvaLyLjmvDVSw6FdCd3S6s/5Lr
RHCjNzXi9t7l94t9xvqQtyZuKbaTibotoZRHMZIo0aUh8lMbf/J0S11gRbL9uuVyGU/f14Xa/ghq
JsNladaj4uB4HFPW3OdHBYOuEjXsZamv8mA2I/0g62Jr6n1eNgOruoeiI+Ff0JQkz6QIFAjNPwGd
8Bbw3hUtQUueYGwAGXFfFI/8dL5CNMykqSaAIaq2wekiv0X7wsSzb+GuRQLsG96KLTX3lBYKn6qK
K9hnyTeC+f7p3lTAGgdHhDw7Eg5oVOLr5DMtyR5NUIIV92zJQ9tpRGIzxT/3tR4bOXLkccjrOwR7
VJ3UvAAIlBZcgKRoXLskfT0tcm/XyTbmD1GppShBYUWlQcPhqqx9tFNkP6E4Yr3SD4zriJEpe7Dg
PkCSTsdNCafRKCZNn0iiY7aKxngQ8cR2MpsW9DC87XXLzvrAMDuS9PZZtphyAMMIqbwStNHFt7G8
3Wrgn5cygQAguWwsGaF3pjpP/Ir/Y+W3ZmYHZrKXKF72JVD2xKUSF8u7lO4kLNe4qRKJy7eBbXog
Uuso3rIBbVov4xsBZSBJhIS43guwT03q328euYBayQEDbrxzhD4BD28NE5mGfZskDezL+S/nE+9R
cxpqvWK3OVJZ4/q0Rk1gI7KstZMak3GS7dI3H6Rw/i0Xt7wFvPdRdBgp4QT/3+uYSMCkxO2Wh4J/
0E8W4oovzmMhnhRG0GYtMd+NsCZn4ujsu6MdLIRtGTK2QyVuvQcDS0zdvAHF5dKMCskIvCu0XhiR
3G6VNeZOR6GUDTLTi5G+/8S0OsaMK4uuN5wBWmZloodTTzKz9xWlULz0Vsh4RLrAblXgq4BzBPf7
03KRQ1fAN8ocjPJmeWBKQN1WhqGEB9LBoLuGcP+SYA8v0kr6eqooR4sV86doEmc/9DgasLZavyau
oJH6LlfjK1MgPSJ7NLbOgPCuBksUtVpthr28o5Lt03tEfxx4MXuZSiU36RhFkooNPSq6Nw4rNYBK
NvboURy7Nh/5
`protect end_protected
