`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3840)
`protect data_block
01AwlhEP6Dng5hqX0ucpwQj9kbVZlDr71ah6JB6UQ2WWLz/862LBOfRiF+fxoR77UY6DcaJ6Wb34
dzIGh5UWWTuQUBYWqVxjXyl+Y3dtG2S9+hs9jnkWRaiV0eMne9LqQxXLfGbqiSFmZjythr0PnNhl
YFZAF6lRZdHCedEbySkWY6LTUdUWTp+JibbYGs+JwIZqoOQchYRL92E54J3uryxQVB5dkXOii/Dx
GFIvXFKNMglIQO25X++sYFdGn7EbMZC2SS6iCB7wkdQG6flg0q5RyKIAwn4dNFwnj2M7Kua65Jrw
/R6El+HNJl7VASLF+7wNstiz5VyAJQnbKx7gBvXBhf3HRiYTwevQxvtFwC4yJJJcBNTv25PYPjUF
hAC9tLJxA+1xw114WrIGuaZYOB8So22zGhpm/F9h1Zc90CbMCGxMl+KUIU1BuZn9d+8FON63CjAN
S1tRGkHU5XbPVb6AcIFYRa6/G9A2qnhYV65+3oCxK+TtYiZyh9EdfIVF3lx1d7ajUoc9S62PVDy4
Tq//+OQByEG4p2DrUCrkwFdtlbx9FaGM29VUDfjX0EPN27yKQexsjM6F7tyTejPfVsrPmApEK0JU
e5FibNxtby+aYFOLyx4nZJtJNHGjF7eTPtpJcdt9Pb1bc0l3juqUgABm3LwhiKPCtAVIYDndcCK2
jv+76AXFqz1RXimRWThn2vzTcvgJUlL5e8O21S30OIz3s5tNei+5/J1jr3NmsPu797Cpg6Na9noS
Xhbv6cLmv0oRb9qXy75cvFrshkG0G2RTp3Ocf/RtVJgvGmexP361Liq3VU6JmwtKjkDITbsztddZ
6Ix8T3kk4ugSlVgFLxaxUlZwS2n4dbwNmeQ7+Awr+YeEkcPeo7eL4NIXY9R3QZ1Lb/2W5IspKQxg
yN3JoKSkQE5bv4oThpXHd9Gmr8th+zwjsR+FFcPhGL2yagOr6q1jtWG6VxOUiOo84J+ICNL6tV7e
VvGbNHPDpG/LrnhuyYNkqlcErDdsekw2nPDkqJCBA5s6oGn6ES6FHEtjrmZLHkpfL715hTfvaItH
SH9xpuPp0gwDKB5kk2BAgMx01nOrLuRAWH9t02OtntQuHSjNZ9B5N5B2KYt6o/pMgXbcyChyoJI0
nCv86WH36d4pWx90NUHRaHcE/OhzGBydcCLTrkgmaNrDIEpv6WpNwL0JAMfwI+xGXY0GHjO95Gyt
65soo2Ue/aJHsabTcsf8z1qg4y+DA/1l2FatxXkQpzEDQoPfYeDWDP7Q5RXE+smpVzgIIeQNjE6D
BSTXurkRm44Ond3wI5zTcoI3aZMcfxf+SRB2IlgF5y4hk57Juj4s8kzQpXuRSnECPm/hy8cvM8Fp
q0Qz3iJJxpCZE8X+MaL/hPH45051Hbb/vydufVkUqcpERREnURshp0qPgYp2GvfOO5PnlrUDo1ND
IeNnv7VCtYBlCWBxZqk87HXBMMvjJ6GuUZzkIUjtg1GkBsLZF5J1Qr0Dp6g0SyTE26fLjBSWv9yM
xLt0BJLiid7oF3IaKLrleFV9aOIaGnCMsj7RxUtzdeyGfMsOrT5PbLMt5/NevzJ3OofiFVATDwIY
PFmtD8/tVHFJ1xCvUjF5VQHl/JQ2yHRrMYk9+MTZV6IPH1SsM0EgnO+XOmHj3kVZP3+LqgwRRbO7
1olgy7+g2kkHbeNhuiE3oaRWfcDOqeuRQ9t8nsjd2DstoUqKe9w5xVbHbsYSSzSNTtC2evfyel3L
0dCVc6rJ05Gk46SE4nneag3zrk7+qcu7kj03u/4Vj09Ps1aD5Koo+S1tZAK1eX3SGQQX73GEaLpO
Le8G7B+aOkpiGThLtL4v6S5SuKYAB6EzF+jeBVSBCByr8N9NqJDjY41LypZKqoWvmH0Zr0en6a7X
N0XCa1GnAgMwghRz4TgbtgLY7Um3Y3Y02i+aSPcIys5vKZJQhP6x66i7cYn39P1H7WGLl4Zym8qG
K66xAvz0Pn0NNHtbx1EX1sn805f2kZBaXHQO+2/j/JKoKdpmxolWzpuM8/w9FANyyps81mMZuC3W
QWI1ntK5emK3UWAtm9ZzszNPQvwW098IOBFazENQ/4TaBiPoHFhtAg3WiCqRPE4xFxeCKM+N7Vgq
uaGLg01w1pueNri3GXpZRRmKB82+Pj3sbr4Fu7U9IDaCZBvOqrNmnYnT8csIaH+4VQjLx/bc4OkE
YxVV9ej+aV5jpbYY8PfAmFIZGGfaYfko8nS8684tf2QVjKV5tntprXL+e1Mkc0V7wLKiL29LJ2ed
o+fttsuDap8xAPWmUdZUbsmVm6+SMzCUORa61ngvvXE04CXTRlyJps9b/fki3gb/bGbOmkmxmdLp
pMarGGjvWP/sCxfO5qmpHRwNlCZCcx5KwxtoJhF9Ca2UwHMcl7D1yPFJR0sAwvlkxJih6ioMvxvh
AJyT5JA5oq3dEVl3IfCdmtQ4zJk8nkvLGbZWotVC1ErIhFFdtyFB0AevTv3WLKCvp05B8T+0JXFd
TOWORBrz6Lrm2J2MtssQn2D53VogqF1G9wnyAyaZNHNx3IXUfiqVBU6aFO+jfXA1Y0RgW0iNLS77
0iQW3JhEmoaLxriJQCrhTfSeNUF2sdVLXQToTrlEWwxvC/0AlwWb2sawsrRM3IeOvdFGesDKSJXa
NZIEfrsduDEwvzmVa/EOC0lbTOODF2UHQJE7wDdEUBxIBt+FcbfKiV45S+WBtzAbIIx5NGKSL6EY
Vqfo7Of1a+dQWaY6qwdnRuaqqn3H4vw7G1+zsA30rQLprn2xxeURopdN0nmVLuoYQ+CnupgOEOkE
oG+10corW53hsf8p9un5KpLXW0vXnvXQ42HltGwBFWVxokKt9VLnR2Nf7c4bmCjgJxz5lnRmIox6
2ST8m0J9KekBeyESrUL/T+mk4v8/7C4EFq7D/LJBroq8vfRny0/iFSoqPrGioTtA9FBXlrNrpepl
0WbAyHJ47LGnY6+oPnNo3JoP2bUw3UyB9SablCyeJTtjjN3wP8S8flDUs6keVyrcipVv8UIW21B0
Q3FdqKW4QY7DZ68FB9nflV3YokgMlSclVOU60rzdsmi6rv7s3xRCn9dyGnBcuNFf7jlSnCy1Tld6
BfhWFfg3FfjWqdm8apCR+2ay5BjdXnuYGs99/m+QaPFdWxEjfXX4HK1/J8OXixRco4RGdUBotIC1
QAS1bY9PzbpHMmjE1qGbtz8Z8HETMxpNtvKROF8w5FUcKZ2zE6GtMvfqygP+WFlhWBOHP4lTdQ69
0CYB+85H/nP36InnxFyVeTrCLqUZ7GqFPzCMfpbfHEtrlOC3r2r0jNjvZGBRonTvduB6YSnO5Acs
wafuue2/E3ODtKs3hXoY0wPz5CGRVUemCLyR5SSi2WAEl3KNqF7pV4A440nm0gXZz8kvOHukCspb
ZWRCrazk6MLyFu2JnJ/PWMLxyFcx9GkllTm6/WgMA0WsWIs6MhLpwjlerGeIXCIxYk6eV1lSSuhf
DuHg3VejZHd0MslEkY+4AP3AlzLUkiFHdSmUTkqQrbyryPUY0mCaZMvLrSdbm/a8EWNtTXrQwcPC
+ug92XTSivZxGjAUmArE/Zl0ECxgc3Hn/pLQr6reFJI3iDnzBqoz+dWKyXGXmBaMW0iyspfnEhY+
cw12LoUHmoPY4VNsXofiiHi+5PtOvc35hnOCAUZN4n/Uq2plv+PakBWmvdIPOHm+ZGuWih0cglTm
MxosfBbLep8jzx1iSsP7ly1TL0q39jeTKum0st3TgTuUw09vQX3o+U4asi89uaW6z8YB4pmbK0xo
ZIilAdk28F7XkeU8YdhKrymvhl3nz37HhoIgl9o99JQBHhie0zV8/s0ePfV6rnUy85lHdZUYPBkZ
wi6txJu6g9qIijXM2EcxVyOoaJnwof0g/nayRs/jB+MWyrHa6SGXlM5CzbUQ3UijNmeJkexPweIV
h+iu+JgXVnmWvEwrqYJdkJ7/7GbFx3iCEW+zL046fEpnDCx2LxGzWEXP4EMw/Ar2eup/O8qlg5az
NQrqT0pKXRdVQHM45EbLBaSGeeUZh4wI3lU6IRmbQzor3wC3qFiwpQDUPHwTynIkeBNTwkNKSw1P
wewSGJ+ivffSqxcEbFl1GE7ae/EKcFQn9bhwTQxnSquK4jkCRoozuVvEPSVdE1FBHxxUhFt7pUlk
hMe233903IJYG/A8jdIC3+e7v744TbqRj7EExkXdsZ3mBuKxQcZ/8vM/6WqE1YyqINboWqKSkPr9
qS83lvf6Y0tbBWkYCHFKOC8R9ouyzw2xQnVQd+qe73Elsrd59msB8lo21AEGSpbmtHmfRXyThVKD
a9vmvMJIrNOquOw5hY8Aq3TTG78XHreqmeGDdvhV/MFQ9N3OopW/AwBU28vLASi7/wzfYeRoBguo
6zqjPmdU2t0ZivHWSTSdbQv0xWVo/4WXhucETDOuE8SF1IcnDktvoWWf3dChmWQqY+OzBEPNQTxw
WCf/hLzGQzC7jH9zXp+JrjWbg0qm25lF3br7ucDjrLx3XXppf26liif5bk/D/jtBnHA0qF+w0VRY
8jVQSEEVexCL31/0N7AaOjAE4HHkbWn6G51Z3RmvUgqwFNundUN5+A63Y6+vYxINcELKugg4eaqP
pyjYKgy4yVKFW/naZ4ww0DJKoGoHBDPmPfV/FwM7sdqewJ8agAGWa4FGjZObnpnGUXfK1q1Z1vAJ
Fg3vD1tTCyS2zI1M97C/j8YYYrwqi9j+qUxxC3Mwtyd3Rm7YutoKz4tCJJuU2iKfd7ozTjrmpRrz
lGH5d6t0c1O7lIcGQxzEzpNhUXnPnukpcz6jDCAcTyth0218Fiiv8oF62gq0mlCTl2Wn7hKv+5WQ
dM5IxYfIG+RLq7xsMXV+K3YhWfBQlrMpDe7VWwGGfTEiq91LbNI+G9Ze5wzovtIfS+LSnSay82/0
x//kDfavD/LJr1BhS5icAhRwJ9j3QRZ2ivwQ+qFaBAAjQMOjIENvcy3q7UnrflSQmDAMmyxhRuaY
7kjHuMfO47w/VzsB7PoKqJOwYGm8SFS04II39xurIYJSopy1HC6tpaQVtoLq/XZvbp6fxpPQIJ9H
nGf9fblgHnon4Q2RX8TX79x2F+cy
`protect end_protected
