`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
baF6smnsQ3rdKio/dWb2kRIoVrRhYcC2KOy0heg+KflXPZjYbIHuoFqd4V2m1fEqfvbBmEAlG0yp
CWrJdXFafyTH4ht/jNImtb1+zKYn7Lc/UXFrzPVesvh6NoYpFxIpBiMpMIjblIY/V5qE6eQm2nkz
jBPk1kcpbOEBpv/3jDaU+HNsIr9oezfIRrrn1O+1F3Z+rHt7+pTO/M+CB3te3TKqvqzrV0QWkYqd
GqXUzufh0dmjwZlgtxLimbAIuqwFD2l5vwYcQrERyk0joFMzrYbZYF8PDQFB0mes+qUJkxJ4rD3X
mV/XfUT2naXFghUck25ODUHZxPXWMx3ihQkspg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="0fwFDrSkWLPprffOOkVd8QHvXWw0u4SrYYPM3G1d74k="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
CSNIc4W+ERRCxBi/7W89idDoQiDA29MVaA3puN9wj1aqLkkKuFNCmUw4s0buV+j8E5CB0lZapxMS
OpIwTTFzoxOfwbg+Ye7MEBLLE4Yt3l/uD0CcyjZKMHtxkNz7MLDYD8WHa5EqeJJuP6T5dZQeH8S5
trXJTimzcySObqX9hGAYzV0kBeDCWjK1tqThYNGx0ZrJW3G1InpmYovB6EoYVZV7xCDOfrdQnBY2
1q/actALCgBo0/qSh9NE7qVqpKiHeace6FohaKgkjsvSyMvpDFI/ECrRCx53vmxOy+AkH06CZ+PX
f0nQ9dYqJH7macCNdtCTL/9QHk6j4bkvxmlM77oTpcliBP5MTKy4Om01t/7n/ElBz3Ku7l62m14A
MqRlAT5GRBTsY5Y56LDRWC89PoRuPEdlIud99CHaAAD9Y33CYJpM0Vx/IebzKuioDGhANOah8UHY
3bJNxx66zeEbo4xnfRssqMQJfZkgNgFQjqX0hqCJkI+/nGMAv1ATEY8AQ197vevkeNOecNy/c2EX
zxYJTX6T8tnlcDmX1nrOIzxBbhCvDbZ3DDXqNx1fTIzm5iBCnIRuAVAKSW+NKz1ws+GtEzw0l4o5
dJQifsLKAxDKpuTEaSr7w3ksDBXadz8Ds5aAwgcrLstOtWJSFEwn8uyIF5T14bWlvftvYeYn7IDz
G+gCWbzMGlWCbtsRNvSjbqdyd1/M6flVosG8duuFricBJFcoe9NPyleppmTVM8rzLf7IQDUWqmU7
j+Y5oddty/d5VOjc7DVRlkTugvx8mk+m2I427R3mAH7ZcXlq4TdYFqnJvv1KETLqD+KioQO9j+S4
cS1QIcnUJ6yrBKRrcmbfYVcF8Lyrn/Hwc5vFjvJNWdXfeZnYQtookYIE6eoeMpx/fskHLqetVwY+
e28EQVmxjFy8zXu6eaWyX9m384vEVNNlNGsn3aXs2Yw9NisE4Z2fn1yI1zwEgeohBFJ/gxyFUQG5
1aE29T/zcXbs3fw4UEkwgmSgdFtH3vKKnOvXUQDgsq1sIkes90mDeVqFYPsvGN/0bYSKIW88BdeC
wx/Y89cneGtw+lr3SCv8Ek6bAJUEP9SLkzfw7Rk9oME3DCT6nq4SrvYIzkiEhBapD2E5EAByi5cm
D0XWBAYCxcjDiD78waYmAxzMpXA4RaICFU1DHcRukroEruvBBPUGuN8H6VBPcs4KlXCmjc0vda4o
IRT6uiAq2hjCLwf7jC/j4uvYi/55TNWqWcu88jacZB8jP0OJXIhD7PDa1SxEiAQ2xT8mJP3+hu7G
Y2qNihiJ7gHpSdBlfXwfp5236hg3dqK+VzRzocFSOsXT5nAygBcOlCrXvVimJH7Cf1gogGQ/ZsxY
vkB4am/ESqkTsEBVa/c6jEpjZP4uvsLpM08I1a575kR1kKg669eEg92/BCtpG0y71hxUY+Hwior+
ZyPWLYmY8Vn0Sr8s+12uI5vDziFFciEQamXj58aCzioXh8O67TX5l3qlxOiL/74t3zd8a2/MXS2l
6pZ8Ej6oMZ56BBEfkAnBK23ChHE3V3CI1POulbAnkCPb8sem6Nmu/fSyKUdn9Bs/GUb8xe6K1buZ
l0He7T91lczqHT7OSN+gSWvJwm+php5aMvMuCBgTBvpKD9XxuG0KtWyjKumtoAr6ePW34qkBE53X
IbnGhIJPbn45sKbqTWr4u3HP42BAYGtADHkl8IRj5ERDm+lpTisX5eqBdVQ0wSXNtNGHzLWz1tNb
zvqJMMzEy0DdK+Cu4SheSLqk7tAakFNs6DGeObe4QIQy+wIN6WWXVnmQYbhQUJv+wTHZjUYVfkPk
6jWhoQ++OT8aA735UMtC0CbEqBMeMi2LOsunnfEhws7bnxANR46qU0XHgLinUBPmmkjL2BqTmgEo
onp79SLfcNI0slxFCj4sqjd8zBMeL9Df1dOTkh3adtnI1B9+L8lK3VZ8CEwG5MSEVWHqOBG2W9TZ
x372/ZSq5F/NID4oBNRm07NkG93sPGRWUHkPSwrn4nRbQeTS0A3lh+v6R2Blx2OazN8eMzTOqZmD
avQMm891TItsYSBe5HR8Mx0iLaNfSMwqQYtWfdK6hPD8DlSLwoaWMzl4qI/N
`protect end_protected
