XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��k��M�1+e1�M\b�:҇=m��F��:�k�2gJ���1o@�	�(�i�Tnƚ�^ԏQ8Peu*p�`%� A�MP��zr�6܇OWE�~������rɚe�A�1���e�@�a&ϭ��/S��VZ�n�(.Xè@斖�$�񮗤V"Y�B�?:I�)þ���[��'�7���;���q���_�d�p�m�6.��3�5?�T�sI:���hy�-��_���p)��(�󨅙3�c�5�$NE�E����dE*�o��.L����YKO0o����\r�vN_d���g�ئ���|���m��Z���?�ڙ��wl8�^�Qe��7�m�"�2���i����0�;k8q��5x<@����D��C��"ǚ�����%��U�~Qۗd���eM��h(�h��䩘�O��|6S��z�ԙ��,%ߤ��aQ@)�ø�L���}�N�B�����7c�D�21�p��ZA^���O4��?`,�1���`s��6�"d��J��:�L�����s1��`�L�go�rӓ����(�o�X��a�/:5 ��I� z��i��o��_�}��v�N�96���[���K��f��ks�N�Zپo���gs\����T���ފ�̼fH�W4v�6�U�i���|��G"��ov�ҟ��,e����w�Ҝ�@�d|���S���~�X��p�:��U�e^A�^�R$��E"��E@�-�-Uj���X\`5~r��uz'�����Jv�TѵD���P_ȣ�2`Pl��XlxVHYEB     389     1805Ŵ�}&.k�/���K_���!������ud����\b!O�4�{�4���_N���vtM�	}�@ײ�Qy@�~~�!�5�AKlp睸L4�T�5�j�W�r���#�����1��R��Ji�8�'W~;f�V�X�	I����N�����8ݤf]j�O�S#2��d��DuBJ��H��� ^�'��5��jIC���,e��	;O�n]��=���M2�� ��0Y���� �X
o���/��B��ь^\����`�f���b���֮Sz~��g)�ϓ��E��e�}aM?��+�93sm.�an�!���2��c�+�G�䈵r����EY�]����p���S�d"���w{��bPV�6�̇��}��