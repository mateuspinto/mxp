`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
kbwjvOZM1DDFcqUcHik40ZXDDfFy2u1FlVAnlZeJbhA2LPYpT8mTAZywUlmrOgGiFYzaJnNPq8Ct
dx6Osq6CZ4BMKCzFGrt3iW+rq9hubR91Bsk1i8D5KfL3KmmwNyTbOU8EdVV2z2HL48/LyldG0ClY
itM2Ds/mWkYRV/DbzbLI45ku6JAsD1SZyEK0m0gNDYI2GYmXXzvZWA9XSiHSN54LvUCcp9r+QA6M
t5XA4ZQsRwQC3MLzObGZeC/85H2ZQvoHpl/GJZ3FdiQZmNdU45LlWWsQcukmS3mc1n39WikeoNGz
40nbtwpQWPXnvdtQjbe1IgvToYyY8yEV/Py/Pg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="bBYmPLkC+y/a+15wbNbJh8Ro/pPk9adbNjpC0zw1KQc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12208)
`protect data_block
w1PPKWwUBgVAA01TPBKw358Pf2poqbkO4SOzpwwJKYFUZYv0sUbWi8YgMTEY2FYcJdE8U6Feu6e3
pBjrOp5MXuyqDhmMdBtNy/hqldNMz+uLL0cvQf4VN5oTNjSah0hANDDSobuL0nJzNdnfqmY+q6YV
V7jHOZRVsKCtph9xRZviEfP8vFtmqlOmZ4uy+xnBVGwEfkwIH6KhfASVoGZw12SwPkH34Z2G5kIP
1MxS/0CI6wDYWWPH7g6LfZM/6X+Ndqc1JXOUXYVx2/3KYNStM0NXzvs7c2jr7mZG+QUJAxAwnf+b
mNJcGxpWyPO7NS00Hm7aj4NivKl+r3tQAXfK4pOX8n4hsy/bH++U/ulGqUvrHbaOR19OgX7zMIqP
Jh9ZULnuRPBKEVEAqjnn/tEAehvS9FWUKkDTafWFiowSfTroZNoMNxKr2wKyXaF0Q77+Fy88RmIs
ypxwPVBM62QwbhcpRSAYPIRUM4lyjIQUhZ69tlZbzi8blozMsfAmJgYd4FWDTOerO0B46LMmXzIq
MSGyArEWUdnzAEESx14E4CSnRmpRXyY8BfYShrqioH6n3oGJbGgjYIlf6ce5jBSUB/CQeK8Eazox
wx8I2lxHlUhhv4LIL1ZzGTKLxnz2FWdle2mu/yBYK1gp0ikZnUwn7UIQtg/ux/szqlmHr07RgetM
bDOKf7xT1rSxJwpS8jb+lXB6tHqhdOQ0BWdWaIwSsGU/nImXgfNIPnluw47URpL3jguSu8FCgwKV
2cbUB+lMdI9v7/ZuCHEBrb/wMf8Zyb15MF+oD4vZliz3J+tVMxzOPO0PPQ/IwLSAMQO/ZIrsbyI6
5akEzB5QNQvtAN9URMxaw+68Cgd1+SCXloSvAGjHS8QzQdrnJPg8jBFL85+UNnsJ5QVMKRD1ZsES
zGzo3eWkEEVTvVUTJyRcN9YfzOd1vOX9YL4fV4lMVYu6/0wWQAH/EjnQn2d5RKu090en/xp8gvdp
ldZapdUgKY9BiQcH6BolCxzvjfOsQdDQqAnguTJphdLLA9rRuYz4RV2azfOxP4cjC+FiA7F2fX7l
Nn3TldlO9Ws9yaSkW/bbXcEWseKwYPrbftJ+Cl+zwyravuAbYzngx1j11HV8q9OXnB3PFBGx1gZq
qaP/S9QqlIHhm7QGehcz5TprDVlDJmeFYPuXplfvT3Ihpp4eAzMLT+oBgy3oo1zcHSYPtF+L2d2V
oST/LDbW/KCPih4u96wyQe1AJ3vp6fKqQKWjKyMseOh/cm2bAqDKKqX7jdIcBjkmcA8qccMs2QdV
ut3npGirjm8dhWro/dJ9tXD1kFKlX5zL+BfRCghA6ec3rkhikxVWyZ5RwhMA5/VQ6Jn2UjVnfAWN
zcPEJxeJYpwK+u3c9t1Ku5Z0gXas7pod8yCxlfm5m2wPGruFdCtlfgvlm45SSBruQIyBO14mTPHi
bIk5meEOGUio33WQO/nIQMUmUQJb7qeJfPHBgevHw8cb8Fv2n3djOzC00StDcf9a5YMyIdBsurey
MRXEGKGfmvY8D9ytfi5eTEsEYsvetY0cc+p2DZALDYQ6QN4HGjY3E6lrCek6FMzkPpvDFxghqkeQ
Bbts/tQ/aG+a3DjnM5nfZSX4FeepWs9EmZjA1kLI6nm38Cr2fQckBHypdd9O7jXWAunoFH6Akygc
mVlcuKvmF9mJberfHUX1E9/w/bq6TRwAPB7n/TOtp7+qsfC4CS8266EBAaFzbAIIs30Di+9bAw50
Clw0mQkIfmOV+4PwnbE9aEnfeakA+YxBqiik2NR/WYPBHqCXjgssvpCr3ljGVipSmEvjgiV9J3I9
LfbXOT//wvpESGZ3QZB4GZqUBzf2p02aBGopD9d9Ba8X9/rYzgvkDIzry+CNFpMc63dAeR8bc8sZ
WOP/wdPnq+ZCOi27ItnX6fpOyidt3ZVOHAu5qM/PH2DQ6ITlM+YXUIuqmRuSYov/X4iZxICR4hNT
4r3W78wics+79TkpLF3LnE5+aZWnuLwj3WWSJnrU3/oKQhzUTGLcqB+owmJOUB3u7CPS7llRfo/Y
otpiAqltwmyWXijqlKWHYg+0eValWtQV0n4ESHOZoTnBGPK8S1Aw1w5lakQFqd1iUxwh0Cfyi9D2
l0zWwb/6UQOJg769lqrhfAFLMKQNcOb/HtTBXGYNEBX54NGQAyZh5S547j2WDyb2IcuZRyBziCUg
WNMaV0ORhIE2GrsqdIGUHzrRU6ZoEFBNZHyy2jiy+ILyIldghqXLUMUw+WGzVqbnMYl6M1BWGDfn
my0C7mHH8YcgnfBO3S/Il4kOphM1y8HSeoJTotu5OWA1FW5OssDxg19sYoh3gtVJ5bMGAdoZHoA2
nFX7E+0E5xAJux91HcruzAmI1CkpEjnfyDfOxrKUs3ZZ+8CZmJqhf0o9U4OBTyVLnieoqQDcXkm/
RrCVRMS8H7IXB1LmYPgQDTQLj7GoLGSMFEYpfq+pTes2+Dh6tnvHDV33ubtP2hUz4Gpge5+NfSHl
oIiaXm/13QEIUevfl74nB5n55QenmpZKO1xAGq3nv1pjpy8+sHww1guctGWwx0yrcv/Kw3US8Z7J
kzwRONJYOn/bqVPIB723ww06ddz5MO6ketTrmj1d5Xv7CTbmx/DnWwpyMdjRnbgvQd5mikg5B4WW
qGtVeB4BtSCjYm0vsvFigTpb4UEfDIMZq2YuSuCMNZ7dYoNnUvRL2edR2ZBnSYcqFlJ176LoYIyn
QTS/HUWbFtgUY3ExLlv1Yt02KVxwqEFCBKCdj1dvcUcFXv/hu9swOXeU8EXKJM2DiKX1fSytYxP+
q7XugOkTItJwjYNulXrw4pVDEJkQe0cTY1fgZKM7WO8ObxheA9qfLcS1014zVhBmUsaBztD8pwkK
0RstQgFvouj1kzz/fAwrK/fIhPoKFECGoRxE5ySFs9x6QqB4KsSQNPCI62axSF/I38TsArDksuTB
wY12F0uy2UpbcINBRXiZqj5eX5+5dty0arAVDJbSgz9e49pmbAp0TDKF/dcSuWKerA2955Fj+K9Y
Fgv0jDbpQd8qqGDi/slw7+y98w8D+Bgk/YDKaJQzC2isIhPYagtj68gE3q+aimBjRq9MNAL8AKq6
DECFZSUOpRB3AX4ikTa8Y9/FmOLS/SIawHlHSbOUkWHmluIcxlfZfopOU4ZlIqo5tHfBJR4M85RY
DUViFtj6dJyGrEfZp4BU50hEP4+LCgo5QurfvFcMMLFztp408Nd6Kxkmfca+/YgXe9IQY361A5fM
AfK/HdJzFyy4e4doulX7efd8dKjjrYf52APL4M0WM2URziq0zSF1jAYzEWbc2081TOp3lxYJkFrd
oi9NhVuVLsId/e75xVgoIFdF2ztohTRYC/aPK6Vf9u1YxyrqFfA6C0aKIL1KYln6Y9SUQ31p4uko
v0m0byUgVCSZsaUFbexxieS3U1tc7ruEkevGEm/RbHhBWdZAHWu16P9KbV+ZL0hKPXIpwaUCwpUF
t2GMRVtyhYlrIx5tfaoxCpz0EL8WatGKjwkVQplPIej8LJBc7y6C5j4g6WYSHY1HNqEtxaEUqDMH
UVewQ6yyZcJRqLzo0PoQxhoxl2ypDvJkXs5h+xvDI7irIJ4VUrogwQQVvC+nxjI2e3W8ZadP8PeT
qRWPBajHEAhRfRNDjY12I+Gkzs7l1F1bFsGq7GHXbVNGbLt/1MigxPLGP2Xhp95yK+ympOojZdGt
8AK4olyTV55N31s9cy1pWzdxWZKK0mwPlzwa0f6suBtxORGtlwrncdNvhyFzFppZu7ydOQRfb+O6
iMAxbsf8hB17gvEDhPjCli5251rvT0i7ZVW2xBhNemC0l73BYp2oRdzunnGlUQNH9dIfpee87Le3
Md8VDhC6VU5UQecjMBNlQxtYudH5dQgVI5uKrA3E1dEhpRgMdaPZeEfyBv01T76ZN2hIFE183nL5
crI4ftlqnIBxb3zAhFvj+549GyYdCD91xAahSfNpUVfWkIei0pxuqTdB7OcMuVybDYLCS5sS2iqa
spPrfcR5QVGVgMHJo+BkKriVpQDB+0E364ufQZE/gm2SRCfyZQgpY2W0h1gHRAPBXcOJV9QJcHRR
ewBwJagLI8CGgDkBtsoyZeZfsX70A8H+sUSdSdu6pipeK6fRxMBvV0cbuu2RhkUL4ob87eYc82V2
vW5Xr8MGfHY/xgccRqN7ljwaIvHpTeuuq7Emp+57xPxUuqt3pnkWisON8ozujo7zfR/I28RpT7Qo
RmM1Mg352lvH9ncdqa4Y8WwgY9BtvaXkV5+GjH1r5tkbvZ21fPgJlY/F2KpRCSMGKH8thefVnOJt
euQmzDVaIQslpvR7v9ox0d4F/2IPfBEskEavAERznkmATWe6xJgbBCAGowxigyeOdg61hrAj5gcJ
MPsuWlfJEfLlMranY09ovo8T5NBzWt024j/EonOInyoG6YQCGvaOdMUrT6cMCcX/SPeK7d4Oa9sk
oGupTvUjDRzJiCIJa6OGeM2lDP9+02eRUEbnt+3cc96mmJHhzcW15pf1gFFyl+Bsk20C0rbst3GP
a/wWNziDN/zWk7wrZjFXE9OoEd+GR5MytE9cH1K3Av5wFVKmeSIv2N60PU+rwPRCu3o51BJcia9f
PQG1F5VdPMiQMm401yyTD6BnZw+1U25OVV4BFpamqyKshtZ5SgJZFIWIhahaAKhy4Z1SGnrtO2s6
k7kwqPpX5G028XwZY5yaN6Puc+UA8rdbvYuTzLaVLJ798B4CndSa3eJ85IvvqW+w3pfAwOfoViFm
LpsRCV0IqjVUYvxs6iQX4RX54xB/LIZKsVl3KKDquTLLf4IV7OYdx7iusSi7NdRtyexgrFxBnaeq
rVE+gyHE7XpLjtvHRTH0EBQnqcUA+VoYJtgn4eJJXRrbOGFpj6EDK9ahcE5AP1KwDk/4oBqjImPr
Tr5ewkgqxUf9XTg5qoUQyq5WJrd0Tx3MEKJA1JA05qMnhGdndsA5lo2QFeLGg/pGLaNi2zKZ9CLl
31Ho30HhIbS0D6L+ceUHFDLq2DOrDrckQHxre8RPhZJ5YWEVLmctuHbj+cZsi4KCrjMPUltadBIw
mIFskKQuKisacd6H7EMzXEpv5ZGBoHKNk8+1u5emLTdaPDd4cyDxVdQili7QArGM3w9lOp9YmddY
LTXXuv90d8Rjn6QRt24GEfLV4r+z19q8s+rRjmpedK83GV/AGUWNvKOzsB7bB1415oUKtxeHtMXV
Fwe1SgZkcVeC3OAFnKMYoEDyUrtJpAAsX98o8DsfRKf39RMZBH+2dbQhlgFpLwGnInzZXjcAvp1a
tTyGRgyv4yow9k/XJr+Kv3bsugM6uuk3NDHOXu8SGpXz7XIw/h0Kh/cs/fBzEoeHfDDviOhF5fqW
QfgUpYBhmIVcnPlArq3JhhK82CBcCyVQqHEZ32/dYajWE0cp0W36Z/mv96WC3yHgY55BBcR0IXTg
SCl2aFEmHEzBCWbDKo1o2OHlJuZsmJiFgex29DwlEOacORx04Gs4xOBIpnNN0fvG4oSHYVQ7PkG7
N+rGnISpJqZbY6VccFLal770n4nswl+T1ucBdd4TWNnLNLIE+4Qw8SR4k8I5ddyRd8YNzrdFei0N
t44U4y2FIMEEQaAoDCX2Jxbc9/VYjOahB8/wfLOYbk1k/O4pmfaGo9MElQS+Wnw4hSmM7dZlxNKC
fuyUESqXFv0PcJROIiesx5E/8xjYvDRuPV4AzjSRsCug50EtLoyqumq9EkFM/jKgBF+0LYDyB6zg
u+SwF9U3w67foJofYaQP6rBjiGp2+EWaM5a6UQXkph/9UM+owNr/o1M/MCdES0s+tZBL1G6Bqhlt
SSSoWDqRcH3iKyEAmesjIIbLejTJiLkEls30AkLxgFQdBVvmu1TkMYfGVYKPRoJWio1SsfQnN9+J
7AtuPPKyI1oqOTCmesU2a7RA2D4RTua9QNrUzutxRnKjk3wQYNNuR/yRF+W9Y+2uroMOPynzFPh+
Ft4zfQWsuTEbVYBSZEjvTwA4azGbvmDtI+YbqPPN/q6KDZ6tc7DnAi84saQ8oOAtsy81dYurRygA
+XxrIaNOhggDqcEFuD88vp/i6UcrkiRR7KXE/miSGem4DBhg/qzvSWSLnCP6buSWnig4vhRp85oN
LtZuj2lK2qmC2ljK4hxMQFvEwjseys3w/GIG92bKQfsS76jiMVoeJQkclFSZSo07wCW1Smi63r8i
vobRWCGdrdTLvEWkfEhBJG390dQOecOnsJFOEdlysVkMEsQw0wiZaqKHFQFz505qvdaMYOaOIyay
jQvOlWGy6F98lMiHv3g9f7EkmlYw89dTmwgmK4MdnXIz7CHG5X/i6z80dcZQoX8xuF+YvBU7CuB9
e/qap+qiAVdcxnUnDfi+PpRzRiZ4u811SvlI0hNSL7wYiO5bDtfzhCqZnHQ7JCfi4S6NF0SbNNSJ
0pcuoiGsbjeTpRkOJu+Z5ljgO1X24lGpeK/TvPFSVB4kNHKBqMFDQ7XbqLIAEIlTKvi0mjYG/E7v
t707PJFJ2q4BPoB9SH1nYNAz8E9XHCiZTgHVQaTWKoBdZDd8Y/YvnTfmX8sJtImglXhQEImqYR+1
Nq2xye9qlN52eLsBQLbg8DEXU+ZebumCocQvQkVsW+ByrNnMJpP7u4HqjENAa60emACbwOuIttGa
Wobr1/Bl9ywVzDPtHvHW4m/9Q3KQ6Dre/PCf9ITPYWMAOvggthkEkc7v/Jwgkc2UyPTnoBd2+Y49
s8CsMGcATVVZIxJXiv+OkBSYL0GVj1JvOv1NBQR7Z8FymufJeLmlGgTay5NIAcLfrMTm3pRFv7UM
9iXM1ZmGDddBDZ2fsGOor/woLFN8sFst6JtzJmaM2MaAtP+/9dJU2SI/LGWkRibbnMAekG7jNYGu
1mvzPIh00aVyykm0ntaLOOMg0klg6qM08fMJ099gzIw0mKNh7TgKojvhMUa4jp2GnE7ff3zMllsn
KOmuruNO+ub5XS+lQ9FKT+kfQosEaOm5kb0OKq6Gd1jjzg/xgtRLaSc6WafDz4XdxIcGmHGsNHda
bHno6q/LCEJV/rlVVN6oDwzY8GzzzM7/x2jNqAlzCKokXyMs1mnPAeMFCGsiS2tuXpJs0k2q/9Fw
YXZA52HVS86f/evjzOOTlRJ0e26XjOzz53SOYcbYx5LvTpm+ffFKk0IuCTs49VxRbaim3pj1jA0F
yT8qmdzySGeqylXZxdjmkQEHs38Z7eRFEHbO3vxvbmQ6EKDI/S4y4I3L7mUawGlTZsWIGt87oUdW
IuNCZx5xhwSMpim8WCIJ8IJ5r5xdtmVBDtzLBwQ5XUHzaa23C2vuZciLpc/B8KxerNbl4FUaHMXy
ffebJfDZJcE/9LsaQ/HMi0xGupsURodloMQhs6EoTQsnagu1Kv3KQYN6GcOa2eBOwuH1e+HzYb/m
wkBFM+dm/z9Hsz0klsFiquN31/G+egCVBzrEa9RJMUEx9V5HhtcXIthcx+llZl/kjQ7cZXpFOxf4
jCmUUKngfBCBZHqj+zhWRp1eTDDTLQmQSQ3fvUQvNzU+MdddUVMwWVijsoKFzRtpOEIGW2ZdnpNi
N2pgFfXnfkD0TX01QhdYsR8ikOwpKxAQAbd14eg2KB7wmf+INImbki6ZtD8GIjz+tx48S49Ay8Qi
WZ1eeo3tjhhvBKX12ECqG92l8cI2YaKCiOczYKEy+IV08HS+3scTDZ5ppBPSmgontNKkc0fJ4Jnu
vus2oheecqveaDOr01jEySzX/EkuOnQg9V7N2BfOWJLmVRXu/JWc9uXTcAY6CoXeX5yRWYIKPmuZ
wP3MBXNWe16znLOWBwpILcaN3DK/wtu4lob/RRZvj1Jfp1HdNDv/HgnkUxMSRA7m5rdtNHiPbgAv
JKqpP7rwOS2wONXWnB1Sio7n6g1oGvp/iF8l6QL1miNB7vYNDmRbjg927RNrnIoYO6mnHbZX1RoO
iEvzyy7o42ruCVE0dpnwf7eWm1qdeFDD8KIF7iMerIrNlkZdEw7ZM2II1zYZtnBZMabC43lXVJWx
lwYPUjNT58Dysn/RC4N6x4prTnWwh3qL6RADl16wAJTNzVm7Kj7oQz9aSekE0I0z7Uvu3xt35Nu2
QNpIRP8nTCVVwqMIx73hqf8+dRvrFE6Hzl3IZ2dHmNjx+vi0BUExzzC4JEHArCRUnAfY+DlXC3+u
1XA33Vpl/3WbqAJwUnY5Jawun+Np0tcIsu3Be2MGCf67io+B7u96zjJmADSWJd/v4Bx8A4o/ZiGh
09IMgyT+Kxks7VfVybcJdYDPFHkuEloZc3XiCYXyLJbrHj06bmHmk8/S6MsM8H2FeCdy3L1rCM6o
Bo1nPc/we2VQH+KC7pvAilxf5c8VDMLRSvqOPEfFAJQzTMeVh6KVxMWmtyKxi104hwSk3l8YaDnH
lsRsSJzZpLxkRoojI/QSa3wobxIHy1YMwdQQlbsoBTYBFBBAZnEQmLyMLd2xMnScf5dpGRPYv4SI
LAWd5h23t/ot0oM7tQr/an0T4m8Ngi+eT+Gp9kcXbBgIgCTuU6GoO7Rq8SNEKDkKwrik846+6Z2m
ibtcikP0L703UmEuP9VpvPfbTcg6XrSSP/JIAyB36aIPkSNLxfKiHAo5Yh7Ijz8rm8gXbtPBNzFs
XDVDMKCgnlOhmbXZWKaF4wGiLOWPLwEzYzsin5QFwDlqFe/Ma7ra/hfdqf2X2ghH6dgEK+XDhy00
B34f8v3zZw/qv+BUG15gu6qDYEQBe8z+Tt3AvN7AT9m8U1bdQNbDR79PjtQ1vcSst0bKoYWAQ273
fbAqtY4COuMTIvYaD6GfUIZyqTSyjsASgNjKG7QiTn3mV/ybcrAI8g+3xym7npWFwfUVvF8jqU7p
T9t/yqi8QNPTUA3p5Me/0dsnaaXe2EzRFDc68RvjNJRSSAUTy80D4B8PxVcRkmK6+TF9Ua1loGxv
EOjcir3nzoLUtj+C5Sn0Z/4qtu7NqaC+kpL9RfmaSkjc0fMKpO22owcKZielDJZScHK7s1pX/u1j
5JAjfIwrEqVzD81/owZZNOYzkNk/M+AXnAHLGicc1uB4HLeY9YOxQBNPh1dAMkZqdOCSFB+Lh9sC
WCj0C41nKQHKyjTDolpq10d3kgdViZUVx5PPFFvldnFWwFkJV/0ZYF83PQd+jm7g5hjv9/SCHVCC
4HYoYABNNoloJKDCLyvo1DC14PH630L2ry3V4+Zt53NcWgXyUDld7u2l1H93UxUUG46++qr5DOH7
STxlZJyPDoXQILEz/4l2avtZubZCKnbldPQPVO9Rbqvjjf+Hy1oqWRuG/a2zMIvAWt1N79HnOaaj
l1MRIynATgaCcu9kAdCqM3EKlFRKswC4/SXfnxV7iE7/ssMwerUlwvuJyl9UM4vDU1EJzDg8fJae
BELlMB3Nx2BmX/9vOOUETUnnyOmcjzqreY2ZItE6TKDq2Bj8iWLtoH+t6kCv9zUhJ4g2S4f+6mj1
TpBDcRbK7zOjJZaZ24sE+5+3eqlTmw0QVL0HAkAeA+AaNwCQT2Z1OYWkriNQkVzq6/uMO2A3yVsc
T4Wd8Ft8hc8pCtLgrC8sCrhmBoI+oiuIG7ldtzB8jiOb1npfurrgOghjHigUbIxrdr2q/Fy6lNLR
PhFORVG1zgoMJ0zVYROEUfzDXdrfZHerrDM0c0t+3DGyDR+dXfBmOEQC3OTqGls5XGZ77hzXg3AA
vroGqTjLopx2PW+u4VK95pzrZlnAipeJXCjpStkOU4YrkdE+OsvJ8bpPm8NMnBIga2s33OYxqlTs
0wk5KE/iaYKVNlXzmlXYuucptByfiBhScBgWtwDofNN2q3vUsJ6ugFXcoxOJp738j9hfaqFpMCiQ
1W1iw2lwFOEoCJDmOCdsZz+ZJ7Bvto5JZa7dD5f402ND21reThMUarjIIh69LQBaefQG6OdWE6Dx
9tYixM5sU7O58OvaykYxfBAf76QcPUW02QoKav6Z0AWS0I3p1MGQdDIZg1aiyJhbkbUUrdNmXI4a
2RiFuW0mP2ASRg/1O3leKKu5PhW6NNvm8DVDrQejnwBTUJaAGClhcfD0ZCAZakF9RamTOVlCDIMw
kdERuZ3QtA3or3gh0WC0RwKuS/F3/+VgJ68GZ7NI/k99HDCGChnf8KLG/oUWurfWyku+lVNsAoKf
xgu0lzBCe+56hnJU3hrn324EFw4Zq0hh7PNr4Qcuh7PM/CdBS/picIgWjYFOS2FOiT5E4elIvodG
/owdD9WpPVtttqoBbWNXBgYROjtpgs7na4bUj0ugxq/uMSBBrk+Fd8PWd8cByT6aL9i5NXiS1N3/
SZrhHT/pH62vCtL+vVYv4U4j34o8JfsuMUXwQUVOxTqZgR7poeSmNbt2I2x3wfzAegFU3o57xt0R
1QuDVWqC6wsKfNUxVaIj7mgqDD6eZAsDf/a2EclN66ncKpsDlr+ON20jDugt0z/avbDfNOE9cFUr
afs2UKfkHYpXIW60pqRbxcvxmo8QIsJy2lLsuCdX2rbj2KXlwsZT+J3rKCNeqMDA7yAXrV/XDNMy
VZFzRDO5lg7ljXGTLOeA35jmuCV3ev+l/OxJwKgg1DAreIIjGRVJYqZG4LkIquhonw2DZ5zdF1na
FFt9dgaNwIiFawnUcj3cV6fpi+OVqvjpGbypoGWpsRqtUO4/tGoKKh3Nn0ClHSAGNirPVOjXNHol
wGRXUV5dcDaObIND2YEQrYG6+obnJFt4Kd7aJHNin2J5JivPaEw1KlZo4a0/2lJDs7QjV59ejUKX
OhcfViIuGv7CGFo0bOgMPORp+sFf75CrYfs6YjzN5xqFLrpFjqK0OzY557p6aLiciqlfP7RCCeE4
OKa39PMOGMOQInIWIukTWfDUwylm2TDfH3uLxXyF8ICIEZnnPGjvV2GF623Agq6X9kPyoFDtftVw
7UaGptQIAegxAWdktLzDdwXXKvA4I7r08fYJDEX56a9mDn4ocR9gizZ1oSjznrvPzxL+H3BJ9D06
BTemvxhwtEjXM+LUzely+64SA+yYkhQYLrbfI5kZd5BCMQuQq4YbWah1Dor1sWZplpeUqC1pd+Rb
fZLfgNyVBQZAYzfRExPFVYfht2G2QGZnarEz3UPTEoNmS6/WPkoENAymtuJL8pMSGPH3tJn/JvqU
DX2WUMNKUgvLeYL6Cfyo3bbearVJzzp8cHo7NID0+aipjVrsyYXUb5ppgALHL6GzNXDsox6y9YWP
RcQ/6d1QYnCTvXC8TTuVVqH1a4bWjg2YWAjwRzJ/ccSk9DsjYpUiGyqZAUytTzvdaDoeUtmRqzkT
F3s0+czUq0+eyIlmY9gGZ5JXYONeN04/Prb8p14NT+LFGEETtrmIH2UroPvhWcT33JCjm+jjXKXQ
plCoiaXMrKCtJqi/qm3ZzvTbmcY9Jw5+7Vsex6uQlqgPtA7rEwbeESsQyc3kZAD+/qC7ukNeDOSk
8WRyvzYbLTkaF+2psWJrxXisPeUeVH6Sut3MbzgFV5p+sWJoiDqsei7mU0hzNOQf9rn0GX9ouCUk
eFxOObLHwUA/f1t8xs9MSDjX1AULI7rjx9q2ksGXSA88D6K8ieJXwN1cT//ClByf9JI0P/q+C2t7
hhfI7UkiMwP2R3qyDGUyZYCjb9OPSPMOkAf69yo0SEesmNlpPjF2UYiFiRvA2dntnI9H59PUDXHs
ZwTngi7phhSf6FQJuXhmsfMeWfPjmI2Hfoa2/4tDLCooTRR4BS/L+rVwfNmjmxgXftGcSczgvDuC
aoNGKVvgfe55jh3aUo8A599CAetrzeFZbzGF9f9QbsZ8ZtudxYk49C30iVKw8BGqGDGhW3JhkTfB
iI7Wdhgpap7sIzFmYwE1l2WG+rHxSIMFIv+UGzaitqTRuJtX4yLthNEnkm/XdAJYrdcW987LLE0N
wldeDLM+ablQCO3PbZoRD2+ZKp7bdkj7dSGiplcluA4QJhFRq9VGjLSRU1/BpZ87HQNvkz4Syk3r
Undo3a/sU3qK8swu7vLL0IJ5l2cR5VKBJRk4EJYM0Gz//roI3nngTJ5I8e450boAxXxgv7CODY20
930rTrinL3mlt9XDCCU4BsptRACyR5uyLCXvbHa0JS8NX0P03LekHZTUFUipWx9bItJVVoDwT+6W
j/g26XCJO+TbduTkYAbodpO4vAPh/hTVtYlIOADQPUyDSoRMMvtOn7phUtQS34g+yEbTtevtqTit
Q2QOlYp6rlCaM1xScuAt46ZdZ9qXHF29pFRN9T00uItIq2bmKm6wv0ANVanBJmMx1UOYAX/jLHFl
fNU19y5ZVOt6QgIP7Ox4Ccuoe6RzNatZB0XbdRwLp8fY/YwUvuYsxya78222YAbCpeiHYjDy42Ly
dyAZ5LY3SJwl14fHj6HFLEdVkoAqAE5XYKjWtNexI9j5omNer6OGy8Me6NMU0SzAnAJCotp1odFu
qSqN037b1YMPHNosT0e8se3yFIVedlAvuJipNzUkiLEkVDhMyyir56PbqTi3P3CIT83uKa5su6lm
l8h4AJoN5Yw0U1J6wkS6vnolWoGrf7JFATphuDNNGao2gnD6emezK6MN5DLXIjvHsA25tzWVhZUQ
bMygdbiPHhg0IcLz9a9Q3t+esMzORtbqBqCifZzrz2nO7uPib7Xh+vwW9GftqKDt11pbUvx+Ez0+
+8rWePHZOZHlrDR20DuSy2ODGD5XLnlGr8n+NvL7KeeVDskjPC6NZn0JsZd45dyhLqKgLveLUyhj
ZCDe3Je/FRU3pTGuvOl9UALreJCHKU8eap3UxeiBTWesV4n8qptPL6O13ok3H1jXRRyw0Pon6W+J
wMvOd//tLZdxZiYOmvFeGbQXo0GBbgq0drtOOFeR1CDmKxfIc+dLjiLa1Px2i27Z4hz4cvT/Vojz
n9zzqWEMgAfac8UEP6TzmKmrLZWuMGHOON4DOrKUD5L8WdsD6U5Z/FG1qE31dF4Hssp96YZkZnU+
yMT0Hpij4wXJe8qYh4ycYbAnQh4oMaRcE7meGESoxaTmI1UO4gfDGO8W+SjBxi9G3wsMMTdFSokf
g/CJAxkIYE5ClNuJ6n0UVvn8XTeHsdy8705q8RGKNVv5OG44Py1qEph/l20pdHP1zUDXfl2D/w5n
AyRbSevmLq6t5d4rQVdhULvXtUBo17143jRykOD/zSJLvhrulHk9XaYIT6RVsqHg52HVc4SvqvbR
cPFu+756FCGmOZ1rZg3IZFRCc0JW80XadZz9amBk+6TqFqcSpy0yuaf/eRPNyQa4LG9gd0+IS96N
N6qMfCEC48EGdghkJl/+Q20AD8mDknKuDP4eTP2av4b1/Tmuysme9n3avii6MALDp7/kndZBNR9I
HoC/hfuEBdHeqvp9cWSm1ub/bgoYCd2sOrQFyEz+wnUjlYcdwmgd3OlucGPhc6lGEiHcIt3w7C0U
T0+vJSbpD/pAWOCl+G5rSu57zQkIg05/Zlgyf+N5pLtdApdanMT0eFY5PTMfAIJWkwXZzPaEkQt/
PvCh8mFmAvF8CATf6WKMOAqR+oJy4EXTk6aXAUAHP8dPEoskUmR1XSea0gez6IUDuU7SdKA0mj3a
wcwuH68OQQXCMC9D5agfFF1R7wtoZERjHpsfL/PK66q6G+MycVARou1Q85AUF8Z0Q9HPz5I6Eqqb
6nlkzYcPhv88CKliyrTF7gSRMYqN4qK/vjxuaBUbwKYyLFE4+jqKBZjDQHqos+c1kvfBRKCGRnK2
a2iWx05zU8pOUdxQz5FzyJu+w7N03WFWjSFShpbB8mCftjpfU3YpKuBZ6qKaH6eB7RrLzs1EFPKD
fMloXafWrpPHqUVF2ObNfPoIGqVF3k9nBkAnyTHV1SP3L6w9iMtSxM7R+OLqID/Hdefpv8ByrIRL
HXfy7GTcAP3wFc3C/Wmhs5v0QPxwXN9obZ8bM/9z36ocFixoF1jslx1/W3aHr9BWLleABCv79OtL
CTJWrEz/Ec9Ubqf/PpTMFvoxdimaLq247T8CTy0UIWbWuvpRy0pICJwBatpbvA0Dp8dNfU6GlGfu
8d/gX+6wjlIovqxNx6/f3K6F0vf8y+wazTFgKe979+dgZ6K14fazkIOe8SPCl6xeNCLyJ6DcwbGG
lc8E7iaLC5lqNHOVIMj19lNUjU1rEg++xJi7NzbX2NuF2laG1xuh8PoO+ghvzF+HH8zNtYHgTBdA
osPLlTrncS+aKsveaxr8dobLdKdKS9B3YhX+84kMqAdDUe81NTdovPlZS3EwQp4My5LYvqfjbdJD
NgccEBnw8m/bCmOTAbgDm00+RINfS30hZfMcmmtY5vA0aTUKbZTaPglmNjA7bvKXYYI3Gr9WHbjU
C+Y2c/x+yTgin1Ro1xP93n6qts5+GrpBHL8gR21rBh93kpg01KMZHFNQkPr/oaobNGE7MJL4BQ/M
wFZjLctdMf9TQa9SEqOIXVQJb4ysONE3rnr+YVKyAWYYE8lEV9Bokn1yqaJnLyrqOr72F5eCLCu8
qKryt7vW7GNTb7SJVMATUL+O1FvlxVBRVu891sV6UfOs8DQGIYDAYs6XM3JQ3XLHoFaU2R4cFhcv
nrBDnsr/G85Z5JwVb7+6wcIZv8H/E1vcEEIyUIjwyk/KbcqcTa3/Z1PLf7AUPp+ccDvhbP+iT9Wd
NXPjy9pl71wqyaRqpTQJ3bCMZUcE6k/hsMdsjVUIEszXWa6U8oP1yRrWhlcgtazdyuBsfXFtSIr7
1HyJtJXQnWrs0VahPmuKkQ/PoP4+ZQQMNDar6OdadoUfsqDOpF8KjNaH7cYujDtpoBM6p6oSWb5H
VIlavoAwunsf8oBE+uBYX/DR0OOzA0rc2KICmSO/aw2M3ugUdSw791qFE660X8NDCw/KjWZUeipr
P/OlEKvLe26xM8BAyF2ouf/+JfEZLQsLX/94/gG4SFPgfgLXEqmqL+cTzfrLAWaJBIgcjzDl1YOt
regpVSyhxIBUpyrVV2b5Clmn8BSPGGew6IoLuaHDB0zlaG+DMySzwlrjjtzqlr2M20XYJ6mZkldS
24Dc51p495QdQtE1LRIWSd77jsKwZrAXZpzoCNXAOpcBb9addSuULf2F8/P98pxVp9plQ5CT78D9
HPuk5hwGN6VJ2ID2GqhGPXFZZwQv5+35zO7+rig8ZtTZY4hOJ71Wt272RD3pQvn87zoL4tXXL9PD
tv0+cZNbf/6RTIJR+AqKKdIdoLGC3V+4lJ4SwiyCh2ls9bXxeeZ/meOXRLKaEEhfNZ3vUod1fYQz
hHwtcJq5coFY+8BgE1wx4dVZVPE9XUbhcm27qxrrcjHI7AiTO2SsmVHCrfKsCprwRe+tdCA3Zwvm
pW52/d29rDzTs8GRA3+tdl/VqRC4s18IsfZJJrCRFahqloBgdVi9yGuL8ToJwMaFEgq6hYxJd2eK
UBSqpbyEYsZJWaBCatYdQSBHO5eFGPqFzokEXtoyccriQMMnYn7HfFjkzFdI8+WHgsh/NfmMp3SC
x7/ChD94Uei9x1ldeGoh/8yKi7oDMaqSybAElCf4n6PsMUGib44FEF8SxF4rzPePimwW7Tz3NQtC
8KLk+warJWXKwpr18ZIpuxYM3eidStwuETznLRdg+Sq4CbGdOfxI5ASXsKjyhaiLlfEXhAUVk59g
m4sJKpjdXdTsBtKQVBbe+COTaJgs+wHdlVCASoWBP/4X72QDgTRrYs9BVVYxqHGDwgQkjxZdb7bR
Eb7omNsiE9Amt5klnOqglPPN4sVNcIDG0fHr5z82WYI7BcK7/a/i4pIpC6IT7wPWmjr0FbPCt0Yi
UcKKS3yD0sacazGAN4QozxAJ3GSra5oaiRhhSFqAtggdM/IzitEkfGi9hnUJWVayuKHWwsistGeg
2hVfLc/ldvrIyzTra2YnFJoTjAiaDL94R1PgP72TjqkNKurr8mtLCQJVS+H+GZ1OnGKfPV92LSL2
rWUlz35Xem18Q/M3rk3fNv/kmUfyP9gqEAVYcdg2524YGHLcicfGQgVj72qSJ3MaJS0ioEAykdnV
x7iEqyRc+xqhaS6ttLZOsnCpgnptmKw3MReeX7v0QfZmyeBa9xzHr1Trze8hThdGgaS3n/xIhAPj
FsvZQvNxzDrVyvTycJukugGMwCSOr/I6Ffp08YUW1Z+oczlLyRVd8HMZloUIva4YZqXwa5Hy135u
P5bSYrCArGlGFcL2GRYSxQvR7KtDyA7OIDybdX1G52vdUv5Mueukf09bKXx0Le5Pr4GjVE8fcWfd
qeMaIsLvuP//Gw==
`protect end_protected
