��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���� vU���%�]����d�S�}�� ���G���KZ��JK}����ޓ��R�,�D|Z%ɐ�zGf�T���tjŋ�/�=�e&�=�&�����J���	qą�!��\����~n�o�D��xEQ�VL@0����
�5/^��G%�{�Dx#�?u{pĢ��V��z�Ӟ�\V��{�I.^�����KL����z�&Pʸ�B4�%��?�-��G�v�H��P���kɭ��p���:i8[2|^��q�z ��د�c�o�r�
q��#���6|����+��6�T�0���LѦ�Fl~ma��D+�LN�}���f$[���R�au-�́��|���s��n�o]��D��Ҧ%�q�zW=����������P�6U,A���U	B�6��/"́v͵��w/���a����,�:�ΦL/I�� ��?R�X3�vG+X����*�����FW���+�$|��Z;E��u�ɚ��:�Nj�K���~�v�Y�{�����ከ.��{o���缸����)R�r�	5�˚�ˋc[�v��������3.����;!%�D�Z�Dx�#,1ؒ���|s��\�^�d6�4�xL��� F,,X�.��TMj�OK{��Cn��]P߁?�c1��ڴ�bT\��ӎ��ڍ��{�8ŗu��.�&i%+����ŵ��Շ�Թ�K��-*c�\!��|�_�[ѻ������{���_�ݾ>�ΎR�}�k$�e:Q%�3�j�$�_�O��ƿr�Dz	�+���^C����/�]���l��������s��P��?H��F �*��m{��-:?Q�>���{�hz�;����Ȓ'>~ǁ4�����~zL�,kU����7��7���Λ��ǻ?1t�����u���M��O׽�
��¥�C�]�;W�`��L��U�N-����vO�[�q��a��@�fl1��A�:M�ܫ���������)�|���'$�i.���,�L	7��d2�GP�qa��s��\��	$l6��H���n?���f�[��x~cX�A�����I�ށ�13��W���L�V�e-dϟ�h*��C'��_�9�U���׋����m�.tÓw˫oh���*����O�o>�ј�+�3"�� �=���!���=��K9ҭN:i��%��Aj�]Zj�|ވ�j_$�
""�L�z#��Y<$�����-���֚>*��SՖ#|?䭥�F%S���N��)��ӻ��
�y${���ji��ND��7��c�P�A�j�G��i�k)���@,�%"~Fb�v���[a�6�x�ʲ�4.������3�'�t�-@�j�c&�֗�T��+���HO�V��*��}�5�4|��fj�'����'�)��#
u=������*נ�H#��dGo��w���ر�jwu�=.Ҍm�3��E-ԑ�3��p��o���Spu� $���RGl����� ��K��J�	Z�,�v,��yym\=6�Ŭ����Ƴ���S�<�������kV�^w�+{�����Rf��]dU�K�i�N-w>+�������[AG[����gT󔊮J��(a3ń��U������Ǹ�H�EKZ���y%�]9eo�*��G &��03.s�e�b������~Z�е�
i$��$�{��h6�l��"ڠ�,�n�|����9!i/�w.��[���m��Z[9���S�i5�o��ob��g�N�g�<E�@�J�p�_�/p�����.F�.� ������Vyz�:�����F�wf��ڎ���
��_��|$�ڌ
 ����v�]@G�/-��I�j㨺I��m����G���L�^S�Kl�sv8�1�)t���j<9#U��933��b��A��n�h�|��.�p�Ũ�)M�ek��z�� ?`�8r�\�ԥCo�·N�v8��"}HA>#1EV5��ȍTyi5�=��ZqB>�Q���2���E��^B�Ѭ&J�\�hy��L\�oV� 9u\��"�G�+�(���NB�&.I�Ns���^�]H�\е(��kXO��M�E؞T�'���׼�"������m!1���;��<�C�)y������r.x|�>(a�#��%�z4�8\��åz�e��wB����������-1�obM)p
d8ɓ��x0$`c&po��P�ʑ2 k̫* �ח��J@�3��|5���:އ�Y,�oV�=��Ɔ��?+aQC6z�T������:�(�R��dM�7�mu�rRx�-k牝�-�0����v�o�����!�'� ^��9\?����g����y�K9d��Cnt�[��~47�%��F�Vz�C���@��I.K(�ڼ�{�57��k���u��+����q�
�r��WϚ�t�W�qţ�٘h'��_�8mm�d^�0��n��}��x��\z��B�{(e�����L�HBk=��������l��sL�ag��*2����>�Q���Nt�WG�<?����t��)Y�R"yO��A�f�"c���gw�c�_@<���
ąb�Gۅͱ	:���"J� Տ��S�m� b���,E�����b5�@WW;ׄ/O@5THj���]�Bad��Z��O��,F�8�Qi�U����a�,���j>��$��ss���O�>��v��`դ���5��m��r��^�TK��7��IB� ������
����r�{��ձ������dh�u�:��;���5k��+#����zv��L����{j�9߄*lcp6]�5��x�G�S��I�TZȞ�Tww{=!°��r,3���n3���l�	�����:TR�&\Xx�
�j~��/��
�&�ʾ�㇞ �n'��ՏL��ʿB��b	h֢q����!�5��b�۽�,Y�8��<R;C ��e���q��������	�DF���XM�׻�n����n���x�W;�x���g!��1V�j�vz�q�NAx�(�:�Ѷk�Ѱ\?��f� T��--�;Asp�\r���K�DR�z��uXD���t��x@�ʏR-�:t�&1W��5!����x��-9��zNLE��']<o��dׯ���5�1 ��t]F�G�Vu�PfC�%�>b��a,�6g�#2d+����s��X����4QF���M���I�t�0�5n�$��a���{��>Ty� W��,��Z�JhŒ��fȓ��Js�8��-"�r{!���E�l{xp/�4w�Xf����S�Nɡ�5Ҿޕ^M1�B+���j
��g�������e:��H<x�Y�������qu���~Wu��s�����U]��~W�L�r|�⥑�\�A����`<�۫��퇥����e��;ӨHN�]��JC���ګmZ�MZ���{��TնX
=�Fy�Ȣ[�
���i��>���O�*� ������⊹q]��Nƴ^���'�O�� )�:�1��S�i�v�3�å�e�G��X4�DL�Y:�h����TV�>�a"?ݑၡI�<�vZ<����2.�n�H��5FnXZ�v(d=�l�4� ��Y���Y4{��G��kE����6tH��L5\���1�\s�1 I$����gJ�]�P�3�g-��㧫�:��~L"����WP ��֪h�u���vҙJ��W`lׁC�+���ѣ�����QFf�N�_r��\��j���������j{�#��ke���㐎�����X�9ȶ��/m��t>�_�Rb�<4��.ă}GZ�e1�f�J܆,�*4q��9��ǈ�XKm��� �d��W��x2v>bP�D#�cb�h4�S��(w֔'��{lR��uoK�����Os���oU7R���Z=X��@ۆ.�>;n��� ���A��@��x�<����>_�[^
,"��b�#^0A9�L�� ��"��iqm�������u<��#���*��ƙO����8���W��OY��"_ h�)���0b����.�����ь��q)e3�8L���\M֯	q�mT^�e�S�b�f��,QN��ވh9�O=�H 6#�<�>��j n�O/n�r��5眮�``���%4�7|
�5jb�]n+�y���S��"l5��Ѹ�q�1��R����u��3F�8O�t�&���mZ�[(��@���P��/K��mO�&�
���)'�>����7�TP���gU�٘���ɧf��D���b���FH��1������+n��Mu@�ޏ3��9��W��Cd�=9π!w�YboWZ3��c*��3p���(P؍��e�(ߐ��|��������wZ��i��ǜ��o�\\m����?h
���w�CNY�'s�U�$�^c�?�LfC�ES�fk{�s�l�h~sL�O�;:g��Es���,$�����Z�| �ON�pE�?��,-�hz�5��X7���S��}W{;�Y4�[gw�7`r�{(0�!1Î�z�-�)vM�9�VWۺ~F��s8��.y���焓��4ZE�1k�H�bW������ߚ���s;�<��+��|��Ŕ<���_���94��fj��_�Q�6�4���vH�Qg��Գ=f&�s�O�����<�md���t_%)w��g�4S�0s��	ǸlY��	��c�{5�	�ס+Uٝ��}7Jϊ�\��C�R�J(J	q(�b��`����}��ƞ��r7��� e��!1��o$ps�N8#���8K=h~$}��I�).i��1��d���E�(@9+kb�6N6ւ�~A��bii#�ALd�������,�RP$p�����V�c�n��?f�J�[?ًQ�e��S5Ӊ4���IwN�´���X�+u{Q��S����G�h���?��$�0��Y{��Z�1ܐ�6���h}�Σ���B�{gh;�Lp�"EF?�d�q.:񀔒�\����f�<'س׻��-uaB;�3E�����Z�6��r�>`�yN���.�I޾�=�������#����p�U�<e�?)���[;��{�Ꮶ���U������3���ޱ��~H�`3��Gˠ ��@���Ő����.l���5Q[z;� �OեLD��A�DL|y�����o��I�=]�:�
�7v�=:z?����|�2��)�y��]S3}�4�Yb�������tRϓ�X�G�gC��i���kU�ʕ���1�[��u�]��rǔ��A�ؓ���^�b.�U�_>�cU�>��g�˘���D�����#L��V���q�y��]d^��E$D�@v���i8�$7��D2r�x��Q��QJr���Os�ڄ���Ҵ�Qw����]W�l�A-�J�6��Y�!B�y-\�Q�(������MK�e����X(���@�ӣh�x��Zc��$k�ت5�,�cQ�+��͸�ڜ����*%ݪ�̙O���%[�<��eL��|��&�i�
�z��&�ֿ����_����}KmcTT�v�>Q�񟣖���z2�S�%��?��|�3����'�L���ZD�C��5��4�0p,E�� 5쵹�"&�ym�!M����%l�L`���A�O63��0��T� үf�C:P�71q�L�t6��O�i�nn�_�޳���P// �lD��y��0�3 �@ɜ����E~^�Ǟ�D�k����J�Z�~�a��,�9��?g�i5�P���I�G��Q��	��Uiqo � ��6o�0�ج�ӈ�F���Ma͘�
YK���;����N�e�V� '�D�E	�=?[*�R �kv=(E	F���W������|�����+����A����R曁70i�t6��A_��1ģ��e4��-iw;wЎ��vef��?���[�TL�*M6\����a�59��(^+�k�8^�~���U,Q���Ixdy�`�)��a9��,0?�2���-ɕևU��YЙ�Ԯ��.���{f�jdݔ�*�������R�ƸSs�T�7�������CKp��f8�*�4(	�q!}��H𞏯R����������K}����U_j�>�}*��(�~���'Mb[<ܢ���ʟ�S�Ω�l�(%p��<�nx��1�^Y��\�C����(�p�Zg]�s��*�\���tf�7*���@譙^1V����G�Q c[:��=+��ӛ\��1���R�/��;y�.��|WU�\$ZH�c?�F�4t4����m����/��7��L��ex:�0���Ћ8,'4�U ����@
�c�f��`���"&��G1�c�]������"��,�zE�vFd[>@b��!vk`���B���bI>u�y�S�J7��������]�a�z�M��!�wT=~�`F�'��QXe�U�W	�z�Ns.�o=|�?'Sp�L�|�WZ�Rcd.|o�!��J���a
se��َ��q˱����..U�G
H�ݬ�w��3 5w�E=��XŎ���i���jo
3/)Ï߅̑����8?���x{v?y�����DpE��7��璟�oP�%����*�X���+-����?���Q�BS(���g(����ghX�1n
�H���6G3�v/�n�y�t�5PY�܊��-��3�|�=M�f#(�z��e�ąB�F�s;�bHKG�O�n3I����sa䟜!�Ƴ9b瀝�����\{��5�y=IشN>Y !�f��燝��-�.F�ޑ�: (2K��Z��vnZI�z8�{Hr���X�ϰv�z4_zY�?e/�)�Fw�����V$�����_%tg���g�M\�yb�Q��Sd���$b���]H����.7���<����kI��އ���?CU`�Io"�U�MmZ#o��"+���7<t����>�c$����R�U)�(�YӐ)���$+�K���-��"����BeI����3FV�O+�D��aj�7������S斉���T��#:
v�^|nm��05l�2���[��r����*=Y�O��jv>�:��f��	��p�ξ����3T�x�m��E�:���rsnj7Z�ޟ�5R���桠, �	l�XX%(޴!Ԑҍ-�Xy�~Ж�:G����<�8��Y�ROE�=A����z�(��o��Y��\+�-���3v�m37��\�5�[ϺZ��=r�<W.,���Yò�+�^Ԝ��y��Us�������Z�vy}�L��dWLGuTv�#�BV(�R#�ǐ�~��#}���(߱���;����C���Ɨ	]�Ȃ���|#����;�.W�F�����������R��L_=V�S��,Eh 2�N�LP/�U�5a����eU�ɬN6���w ���B�Q0q�\����㻭�߇�&h�6�)bv�c"�~�<�Н�J���=s�D%�/�ӷfV'#�i���5��M#|���s���G�&ػ�����	���v:�F����*��@h������	���?�ο��eH���ׯ֊����C��Nn�荶Gz�K����^��6�Z�0 �,���i ����I鰠5�{ �]0�o'�3<F8bK�|���n�N
���Ak��fe��V(E\b���}T���|>���Pfg)�d�Wߢ�
���$ft���=l`j�w{d@�Ի�0��:��T�EB�eYa
�V�O����ι���{�J��K���f��5Q�����x2���T0e�l
��I��d��^�6LTf����-z���d�u�92���.{��*n_�Wg�T�C��Y��^t�2i�v˝2�a5�?.��[M��^����!(.���-Ɇ�O���2�G��5Zj9E�ZXbí�nP#�-]�lDf�0�D����o����
k��M��wC�h�h�gm���fΎ�w�4�8ח w?`�Y����9"��r�������e^]�U��g�H4)ȣ����ɓG���
�G��{�!�vE�,����f��@�m$�#XLv�;u���$B\���-_�4��7p������bJ��.�l�H��0�J�K��J�FK��b��y����}�ϣ&b��{�v��.o����,N�I�K�L�9X�<���{��0F�^��9
")�das\��<���r�^b�aWq����rH%-r����{ewL��A-�����(#'�q�+9Ip�>��R|�`o}Otƕ4���Ϙ��/��:�q��F鮂���@5Uz -���Z��Q}�3�ß�/]v$l�}=Yں�	���jmk���d�Ո-�q�����2��� 9cB�ӱa�(��w�>b5��
�c�!}6�d��p����-AN�kKm���ΥX�/sXA���䥲����/u��;T*�����873��ӺB�H�����'����{B�Z�9���s�����c4hS%VR����!6ߘA]a��,M�"��0���=�~0,�9�,��2�3���L)	A��u�!�����ۡh�r�gZ����������ک��������E�dU�r����Po#��0�G9س!�l7��2$�����7XÚՂ;�`}#�¶��n�#�t�/�����,��1�oc�"q�	�S�s�^ځ��!���<��NIl� $߻�]ԫ����nU��Bd![�Q2���7ٓ����u��I�H�\�<f�֐q#¾^���<�R1�������&}EN���0qVA��®�s}X:-2���<r7�i��P槜��"����[������:$ӳ�'ɉ��q5{��61�,���K6�W���s��,�GbkuM�AW��O�|3"1*/���	]KP�JY��,#�8��y������=���_V���OTE��8�� �nU�Pb#�8B�dd�`� W�\#��W]%$�Ԓ�e]�Z��uer��<B�!<�1�B�a �Wx���Ƭ�y��}|���17~��U��q�P|�!���)��4P���wp��j����k�O��p�`�&а�z۳6���{���y>�֏d�,s�c�^�����W����9F��w������lĝ`MWG�7C�?��mp�B�6��`�LTbyt�\���.���4v^��?,��tc��4.e(�
����f݌/Z+d9���W��,tD�����0���{;�)�|EL7	�`J�cyŴ҂��>���a)[���2���w�r������Ț�C\����Q#=�\L_M"Ͳj����U��\�f�y�:-\I�i�u��lX9�tK�=o�O����!%b"+iI��*�Iu,jT�jֱ���U"�J/��:�$�:�%�0�c��B���'
�f��q׊��f�m�l�������9�_�}�r]6F���o��5�Fr8���I�G�u�ћ'���j�5U�=�R��ݭR�����tp��ssZh⸘=���n�Sh��jD����g��m:f���'9��3$̛ճ�'�?��k�i�[X�"��9��w��/��	M�]�L������wQ�!&���h7�L1�k�����Jۏ����+��3`�ް]׆��
�89w:q,�45f/�5$�����2���_˥{�Ii�'r3p�]	��N'˥�/� ��n�Y��RD箥�W���E��ӄu��d���	�Y,�����>�0��#�ѼO��JTSo��ze�X"7���	)�8y�AA�>O��38���+�j>nܐM;�qZ6 jfDLz4���ߊ07x+�hV��|q��ˉe<��J�Z��ö��OS�E��;<\�R/�)9֊T%%��©4�����P+-����}E	��M^�_��Ԫ��7g�fN{w�b��RN��O�ǟV?L�m�A;��<�/
B)ѕ�r�	ǚv���>D' Y�n��.��r��o��ܖ?� �l����-��.r�n&%��	4������pܭK��|�����\�+u7����ZЉ��Y*�>��z��bfc���ݿ.d"�78���0??��f����cX0|����gi���C>�����ႋl�|�Q�I��z���֩K�F�����[�4��N��4j[��,l���	O�c�$s�EQ�Wۣ�ӣ�u�<��S����%�q������T@0�yp��z���E���\zck�����b��X�1[�F��������h��;j��5l-^�Hy�Vq4�R\I�%U��QgU���aX-��\�����f����$
��䅅�)r,�Ou`�,_?d7.�|L���:<�H��P8��K<�iCZ{��uA<x����\fO���ih�E<b"k����u�+%#4�t�6�V>����}p?�)9Ρ	��D!f8�Y�-G�h{��"�[��6�K��RN!"�|_��;a�Ш�����@;�GmXb(��ʍ<E�WW�pX���=�D�P�ٟ��܅��u1ܪ�}p�*�#����v��J�~�� tS��A��rv�vq�D�I�~T`{�J;;�c�b�i�A�Gb�wT�I��wL`D=�C�uӱ����	)䞂Jܺ�36I�=0�-���K��1 ��5��R��&���3���s� jk}?0�b�j����N�:	0H�c��3�h���۰}�u�G;9�7��QzY��k��{zD�[��W���!�`�Rr� �q�8��P�����\V��FM�hoz<w|q�[��L{���N
�����. ���t+
-����Pq|K���ǔ)c\��0lB]�1�I��4=�iJi��O��DA}�x�.�*�J�֥����È_�����s�SV�m��K��b���o6+f�pr�!`���碟���~$��u����Y��_(�
�|�E�(��
��2tFe��]ߌe��K&���H���`}�򱗯�V�_��ey#���d�s���XV���J���iړ|��7��+!��_iFhw;�����{ٺճ<W��.~�;�����ҢZû�Th���[O��2&(,U~1�2e�l)P#�+O�W塌:C�B���֑�]�;���)I��Q��VX�Ѧ?vׄ�"�&��D$���}25��dGO�#VSP;�#�畃�y)�5]Zn/y�����s׊s��3 �:�p�>��M8�����?�i�3��� �1�$�
X��W��o�R�H���%y,�\]���\~�g��β��y�^;�>r6�L6���;��,d�W���^���/�\HLsU��Gf���'����Dj�v���@����͢`Z_%F���܂
�� N'�5
FK�eۀ�P^v���>kq
�@ЕR$�U
�(�^��ۂz�r��GC�����Y�ݑ2���Kj�G����	 �"
�i����RR%��ܜ��<&����3��e�4؈���w��Z���F�x!��l�}@]>8��Y��e�)�7,`�@��|�ч�TX�xymW���C�\���2������ȲT@x�c�yⲢ�-&W��+x�XM�T��Պ(����U��W���'�֨rP!�@���T�1�|=���B�M��	}��uƙ�����]'�rs��0E�9��ㆀ�x����V��%3���XTb��/-���5_գ.�af��2Ѥ3�p{�5sS����bɚ�ȼ�ˍ��)�(ꈫ���$)O�`�TL���]K���D�03�V�N��f�)�u��,ΫP-��1�g�"/}�K2ף����5��%*-@�}$+��Ӏ��������T &Ъ�R:�2Rx�*��Co�>�^Y����Z�Ӹ �كhLֿ�LY��V��q��=rci[�NU�qI7��濑�RQ�� ��w�&�p����'�G�v	��(bɊt��n���F
	�`��.��5�Ќ�d�����ݜ�����C�>�y�D�T�v���82b:W�:Y[z`�����N[4P�<�v�R͝b��6�#�3v�}�rl����s��wܕ�M���~�fF�I���O��9dc`,�^P�9����pe�A@���%�y!![]DP��gl��%�i�\�?�K���Oy4��Z�=�R��a>1�m�"e�Ǡ��#��^ˊf�C"���k?k�|gnJ����܏�@��L�{]#Rxk�� G_�fD�������<�w�n�۪�D��0P�'׊��S����Z�3*Px�IuTn�_� ���r6�u� �Q�^A4^Şs-��?�}��o��O�!�f��-�rM���9I~��E�eԯ*�^h3�Xk[%�1@�R�.��ϸ/��f���p{?l��j:Y�7W��.6 m������ೌ�D�H�����`�\��gE����b��7�$���OIU��x��W����B+ϧ���wꭇ�M�F�ݎx�ႁ?X6;lݾ�kn���� ��rK�����LEs�³EDN�Yz��D�}�|',-�FQWm|()�j g��"g���FKa-1`���uV�\d�k� �&dzs?u���q�=*;XUu�q�gq��)�h�!o��n��l*�aX�7�yPO.#���1������,�˷4��A��0,�C��֭��
�����o �Ż�nS �\����������xRZ�Vֹ�kE����%
!�=���1���h����"\ PMQZ��=S�&2�G�ز�^Vӡ���}�u��Y�2L�5��C�ª�Lnɸʇ��k����D����O��2L z�ó�g��v��LWId�0�{alI�p�2�i�"#������!�xf=�����ŉE�H]�ȡ��F�˞��먆�xң-0e�g��=fkHk��������w�ma�%���F� �\S �r)�e;Q�j[�ls7���F��)�}G*t/K5vwY�1?���v6��7��x_Z���}�7�+�c>9�i%�Tk^�	
l -��=���(P�3��'�_�]BFH¡�v��=?73U��yT�_fN�р�h��w�ž�%Y��W�yԃ�����C�Og��P=���l�4�V�E���	���U�s8��e���R6�ǩ�����@�x�ભ����G�����q��A�"�����	��	�^�-��
��qMy0_4 �5���{V���IH7�NPv���-���^�+���1����m#[��`)���Q|�ZQ�$���"�w��FٖaY��<��*x��ZI`��2�bt ��oI�>���f,uC}��<ie��0�eB6�E��yC���y�ٮ�����!.�U��G�V*��W-�����l�&!�j(|9��2�2��DiU�D�;���˲�2�.Ն}=���J���ŉ����Msj0V��k]�˾/��eE�9��w�|�z����Xbo�nh#��]��H~����}y���j���h)C<z��G� ~�4�:<5�A.�����m��k�U
���=��Y�Uʤ��L�|��z�
�O�]�(+m�5w����Uag,E'6�I�7��
��W�%X���4V�]�� lx$߮���#�D@cQ��ܥ�F�M�J�ƣq(���@.�Z|���@�ʍ���is�)���1�*@G�21�O�Z:4���T��<��p�R����T�����JU:HEv�$ך�U��fQ����:|�~��E7y�u�i��s��aUJ�p����rҶ�t}G�����4Ь�D�=�����3�?;�o�{'d�����R�W�.�.j��%ĝ�T�s�XiưK#k��d����Õ]�1��5�S��r����T�'�gR,,�X�����B�E*�w0'��φ(Lg-]�pa��ǃ�v���˾}�w�]SKwK�Rnk��L��JĆ8���K@*.�1�靊d1 �m0�k�M�ǜ8��͡�؂�׏P�(HTީn��gx^��jЂ&�CqK���<���8g<Mh"��ܿ�g�B{K�a�}ɤ��,�O�,�ɀ���#�8rʬ�M2E�3����F����W���Z�o]sS5^I$U0���/�A<&�\ܲ�~U<�G��g���i��#�O�]r�Ë1�-��κ ���'o�ѱ@ro{�'��yf�D�x���)�b�.2J)�s��!���j�L���y T|��;P��u�htv�o.�͋�%�8bݖZ4'�f��Ǡ0��d�G���G�����ܖ�4�xUN�E��I�i��_��,��hn��sq8�d�9�� � 	���x�Ҧ�ڑr�^� �U4��\j/��c*��TEq5�(�J�R�āCp'鐭7�4|;�;�$��z�jM��|'�%��g��:�T����^[��
X#4���6pv�Db�������l��;���-�m�I�C ��NٹL'X����axH�d[����Z-��� j0[�3!�9eW��l����	�0���8]^��*&*�� a�nlb�8=6%1�i��Ox�W6�4�+aT���t`���M��� _<��ϩ̡�Ρ�]i�¤;�UyY����~Qc��_e�G�8��9S"f�N.�M��(���юT�GM�c0�[�-�^iK�j�����3�ZنP�+w�p�g�B��X�_��y*�-����7����u�����Mdߐ}��}R�%y>��?궧_����~V��7��=	��)T�$��D=RvH�9.��0�zg�Kj��
�G�||�1Z�p��uM�g�ׄF˄|�lZ������Q����G��ڕ�K��r�u�XQ[C�uDa�b}!��7����W�;DD��0j���v˩�ϒ_1�s��[�?b@��lٝ�*���1���U֠ݍ=7���*K�ip�IO�QIZi�k]B���B�MUm��D\Zb'�����>�V��mA�ß��{�lN��l;���q@]����HZ9��m�d���Kt�"u���̈������J�_�J<��5��Bb�|��<`w��Kc��(��R�ج)�������E��3��;S�&�!�cL�>�8n]��?��	�υo���^��5Tj��Ovys�w�ϲ©\�CJ�  �H4ؖ_�`-|�%���+Vwd_*թ�6���.��b�zik��1�p_���2����f��Z��Ő��6(	xk^&S;��Hf�ah���Ii5�J�d�yyp��ftg��fX��S��dlL}��b�`&o�#�pLt���op���������_V6�uh�6�T��c��<9<[�bi��C����.ǋ/K �u�_�(�Í� z���䓽_�L̖Y��c2��5t��'����!û|� ^2'����5���y���ّi�r�y���1�������Χ��TD��14�*�:��(MW�F{�0�T��\�f��z�O�/����I�ݧ�P0�>���r��I!��`J��ߠПm�\���a�d�`| þĀ�/r�K+3�=D�俦}���^J�o;Xs1"���8�ȃ�� �b~.�5\B��[5��s�Y#�!S��O� �^Mņ��`=^�,�w�RO�̶���9�hdBwd�?m�-��g��q�V��8�M�q�N�=�R9��Y�	U����2n�s���bZ_~ߓm��F?��ں���O2~�S����������7����1j�,�FD���R2ƃµ$9`a{n��@m��'%���Z�a�#�J�:�S�1Qt��>�fT��R���/���/o?�-��:����ľ�YAC-=�b;�ņ�I'��o��]r=�| "|ۙ���`����M�	������¨�0D1��\��!j��E�֪�ȁN/�"�	�X���z�l�ls�%��(���Ѧ�f�E�Tl$W��Ĺ/�0u�����%�8z�����#����M}l�?�o�O��K۳�H�,����h�`��i�]��SǄ_VG�J�i�-ɯ�w>�C�>����}̾�嗐������ޢ\�Vp�.�ۺ-6i�q�/�}��:lH����y�K�$*Nc�l9E�e���Dt���
�+4$�Q���@wxIM�@*R]��FsaCNncT�?i��ĥ�����ñ���IWȋbtl�.��_Q�'���OL����)��K� K��MbP�3vƶ�|=*Sw�0�TXa6.�(6}�oz�S�{�6�����Qܶ�0��4���ң�>�Ֆ�����B�.�T���"��v���� �4Б욳	��"ϙU�#a�Er��Wt��r����9%Ar�}���jա�����<5T��"���G��)p�����HG�j�����g1����8޲ಳ��s�t���h#�~���p����3�fv��;{(�>�P�����E��♴P��G�#ݚ���V�$Pu�PD�-@�%�ZA���ji�Ӧ.Ƥ˥��g�r&+x<��*�=#ĥ�� W%㠜�镍N��=��}���v����{_,JEJG��AVp��N�^;�L��"�5������^���S�o9 +K�6��'ȶU]�F8 �v,�	K���؀�-%���adϮp���Gj���Io�0�g1?�+i��\♹R�'f�+o�Ģ.J�3c$�(E~���aĒ�$!eGlk���"C��t-5����7{�R�:oc
%�)ps�H���e� M�E�d�P�]#዁��N�4��P=��q����m��G�(���V�r����v�:t�灚���V"y����>9HXM���Z$�.��C%Ωlh#������������l�e�4N���N����>A�XT��g i�s�OL=%ƿ�B�c8�W���i㉙�/��{��on���s���]O�����
a�g�7̿v�OJ���~T
i��I_l���6��;m��@M��%Ho�4�r �oKOLˈ;�S���e�`6,8�\_3�k"?77�w�ȍ*8�d�T�/v�+�[���ﻗ��Uz�F�M#�L.��w۷��r�l�|��ŕ$�a��]���>e�w���q�H�+A,4����	�����}tiS��7a�Д*�I�U���L��E�U)sz����Nq�Ew��.+K?Z�O7��j�� �yJ�v	��@z�aP���N��=���R��bQ=h� ��
qQ\�|���7�z�$��a]�G�a�o���t�yE��3����+n� �Ua^A���?
{�O�]5���	3Yׅ�-.l �[�Cn��Nr�D�������c�#�%g.���}B�$��mT:uvf|DC�S�M�O��M�c73�\OȄ���AA���U7+��ǃTL���c
�r�/�ж�L1K��I,����c=ԆF�ȿ��.��?!ǩe� ������P�#���]�ޮ����:bf���L�-1lK�?��d���4|K2D���]Ie�= N5���)�snv��Nb$�s�]���Wd�g�\$�!��v�������N�lГR`ȟK��8������h9 ��Y���l��ϑ;G�p'ڻ:�H%���^.:���܊p�W���h��� �����E�fIڔ�p�l�E4M����^�ڵÁ��"��	[Y�%�bx�����^S�$$jS{F9���q�d?frj�St�/黀ڀ��?�%㣜%F:�o�9֪����_����\F��SBZ4�&L��*&Y����,6�j�Qƍ���¨kF��d�_f�)��0pv�j9�+�WA�H�{���}u��.1:=��[����[h+<��|]�gcԧ���(�������N�쁈��ft*X�c�?��%���������_�C��*���,8�W����wa�9n��ތ<�2������鰷Y��J��-#ӗ$e�#�z'줖�o�b�2ʿM�:�.|
FUId�]F㽳 �K@�(l�z#V��i��5l�d&�m��ҕa�BC�X�Țu?������c��>��#	4{bV}�Y>q���΃>����o��'Fw��!�pg�lI�7���Va�!���&s
30X }.ު:�;d��vtq�����L����  ��{+R��R8+�`����u[s�=ڣd��<���PF{����q�L+D��E��,h�I��<�*� @FM�R���
�gJ��Lt�
��9c�H���T��C���=T����ᒙPQ�[��n"
D��P�%���z��{7 Z[k��O�_�m���6@��팴i>�j�9���4E0�ډ���R{̦�w��컅�� �i2����t8�� Ii_��j^5��,�m(���L�~>/I�}$�i��4���䥢Z��\�;����ؕp�z�QO��u?SQ�.�b�W�O����Kv X���r��[�� �[�2��5%_
�kR�d�<]g�p�1c'Ƣ�?-%�k�׮�-|Mn�ȅ�Wu:���xƕ�]C�)�<�fZ������Ih���B��w+G�s/i�2�ҩ0;Da�N��lOU���#��E���f��wΆ:�B���X�҂Cq>B�!
��!���h��?ϛ1�.N�d�o#�#��o�+ u�զ�gǍ�Ոu��<�J�Y�� �n�rC���%D�T$$K'���O��T���"��T.�§ma�+�P34��ũ��by_+�m�;�c�!0]�g4��wi�h�r_Az���o&��M5�@����^��]C��H;Ե׆Z
��KX$.����b�z������צ�׺���z��"^Q��|��O3�J�k��DK����O�޶�&�X��}�$]�<q�|�=q5l���.˧����!�c������Z��Ʋ�=I3��w-�K1W������vTO��Ns;A��D���B��Ĥ����_B�	�ur�+�ی���4h̒�`W@nM���5o|����&�y�FP]ӘSX����87�?�7uЛ=�Υ5��G��Ý�!��O=�M
+�IP&�o���<iz�w˼�����If���1g�[��\:����K��F����g�W�j1���=4*��X�nb�i8�<	�����!&��'�6xHީq��WE[i���QL}����.p-���@:R𸒐Xɞ��%�:�e��W�T[��<�
�2�z�f��@�<«�	��^b�����4]�-�� _�&��H�~b�=�`V��B�j�� ��F����dX^!�b�0�,r��/Ɗ�:�I��:[;��	ZoӐI���y_�,��6���h�)��/d~����D.o���S7��R,�|1!�b,��R��D{��[���2�&BlF�ՇW�Q��㾂��������gKʈ���g�����^��#�xd�{|��Q�d=��@�B��e�W�����ωL$����L��x#�S/���To.�����.�BN�i��� ���S�X�������z&��D]��s����I�;�h����>����$�._�{C�j�}޷�	p�*EN]t�h0x��o�zC�:HWed|��S��0�zg�h����9����:q4�snO��j�Ď����6�鋠%l���^�x<�6�l �;6t�] 0n![����X�ꍺ��5��#E},�Z�x��؜D��s��V�K�8-y`��̂ӭ��Xn� �(f긍d�V���Nf��4��\q���6~fd�y<��R��n�l�m�	���p9����h���*Yn���t�eXN������?@�W��.���f�,�`�1���0e��^0������Fйـs�/0�N�
��uc�$�5"oj�! >�A_���d8��!3�/�o:ze ���2#�U��&Fa��9'OՕZ�	%�a��A�]F.b(�{8;G}���[0�d����v �N{`�]�����s5�~?!E�q��8��b�����͹ޭ'e�`9�S�=��8�NX&u��R2�M,_��Z, �^�G���Dj�)0u]�@͡,�TN��_O���a�E���Bi��˥c'N�)Z�kh����=�Y�T2��R�vp4�}��u�_�#1��%��:h��6�(�~�0���i&x�����Č� �jğ�(�	�D�%��+^��(�*Q���,=>�i�b�$�:��, nj]���~�"�(�"��3DB�]e�:�H�Uv���|4�G9֨�b���+�`�
&�3'E�v$Ձ�[�R�OBv��>�^�#xCM,��ȇʧ�����������%t`P�.�'$�u��.��pg}�C��.��(�Q�����G�i�%-���8R�x��4�*�M�4EU��2y��qN�t�V�$l���RO�ݵ�+�2A���u��m��)�3�𓻕22�b�Q�[� x�m"��i`8��"ڊe����S}�-�Q[��j=�~W���1\W�p'<�p���Ũ���$�M�+��83t�u���.��7u��q��1�A���e�][�(�.�aiI��}�,b�����/�m�M�ɏ�5�r�+
 v������3����5�Jg(%$09^�Vn���L��0��S��6�$sG��p�P%ͥu0!�E��a0�fn%Rc�?�y��J�d����.h"'��R ������ص�j�h�aW�ګ�̊q�DS�>��T�KXϧ��%U�8�u<���� ђ�lШe��d����Ĭ����h����K����*�+4J�ۇ�$.����}?�)�ѡ��sf����+^l'o��ew�:SI3N1��V��GH�e��EMm栚�}�x���ˉ��q��˿	��R�z������&|1�9�Q���7�n�{��X���a��,���d4�I�J��F32�w�,ę_|��D^v�j����[���R�� 2ے�!me�شct��j%�9����Z8ʼ�H��s\�
(;F���O$<vK���b���G�]��ΒI�Rd|�_�R���w/ɦm
�?D,^Q��+�Y�n����� dH�@�T98i&H�.��9��E�����R^�?|��0��]V�"�un���1$�s�I�.0�层g��=h�"��*i��	'b�����4��e�ѧ*�=_�vO��s�\,�Tm�ؿ n�q�"� X9���V<x�s�!<[cg������³���(��`� ��T3��=�)lVc��J�&�I*8%�h�N����;�*�� Z�Ѭ�QA��Mg.^GK�h)G��S���2~ڧ�UҒ�)u�a�c�Qp��4L���á,��.\ݨ0O*�*<qS���G�G,�I�G��6�HЮsQFR�;�bPԉ)�ќE����	`�OR�ok��aӻew��� ��p�޷*��nAU��gf����?T�l�Q<���tf6���_�2W���[=E��)�ǿmM��v?R�TP�}ɢݺܝH���g�e�r�O���J�$vɚe�gi��>R�_s�Q�,Z����k��ew��\�s8��y��$x�[�;P̞l��RbG���72�<�s]'5W�I�
���-p�6;�T5S�*Mgx�]<�oJ��U�[�u����m^ZRO��. 2G5�h�E��e �N6̨�6z^Ҷd���XwͺiDJ;4�9���/��y�C�c������u$8!�R���u�:����}�:�^_��i>\Fj���UՇ$�<�N�̂���	���߱l���|�=��~�$�ɇ8Km3��߫$#=�`IO� ��*kΝn4h���E�S4�!4�O�>��=&&���$�2�){�zY�~�שּQ��P��K1F���0�k��±�(DG��/�=� @Sɡg�P㳻�ɻ����5���6V��%��Ͱz��4�?�&����E�DZ���|y�ǿ��C���| uo���s�G$=���r��jZ\=�t�Y��sF�iє���-��ف�@X��]1�w�b����7gU�r8a/P��i��o���lQ���I,��O�y��uv�Jߦ�G�!�tP��s8�֛J��-�x���B�=C���5�qˍ!�����etY-����k���P�~���j�~Ob�&8�������cm>r2U�����6�:^��&�@��C[w�{Ft=�1d��0=8����KOw��]�Nm���[�Ȫ���Av�{�m��\�rJgO;FF�6B�+]u�=�K�8xD�i��H
+���n�����;޷�����X�����xC
�^l�uD�|�v��ͧ��f��f��isO�FW�#���S���- j�bBb$N��h�J>�e�.Fu�JN#�� Mt!�^��q��C�h�'�}Zx��m^��4Dn��#p X��SX��M��]��x&���\����-����D#�VQ�Ev |�4�x=�4�������F�c	��B��:���I9R�h��#q�8�c�y���!��݊3��.��uYp�ㄢEj�q7]��� +�� �����[�Y;�T�rc�
r}ԤӪ�.��'ۃP�r�C�[.��_#��gJJ���]]�ǰE��pKd`�2(ɜ��>��j�%:�-��3��{ݷ㺻�6oDr�i5*>�m������D��$����i��{U�$JjC6��=��յ�F�i�_�tY���N��⬦��E���52r�O,�6�4���\� ��s�,�H+�G�v����KXL!��������q����^����q��s=��T�@!�b�P�8������Z��IKPH+�5�j'��A���ט+��ה���؊B�ش'@+B�����g��i�pX>�S������3"8���;��ʠ>�!h�q�B:������ ��\�+���jר��#�9�Wx�z?��F�G�?0���#�W����^HCg���#BjҰ-����)���*4k�L�s�������p(sƐ�C��k��.���Ԉ��3���æke�-7�Z.X�s�-�k@���L3�CB���Vnq��
}�i����� �6�J�l��Uz[�'��l�~��[#k'�kA���a�qPz���_˅O���y�A����[i�c�g����^~|��!�y(0���K�����A=��=Kcɼ��@���q x�ź�X/�#�G��m]��X��� Vh
1l3]�X���ڧa\t7t)�ۺ�]q�eU�r���vuo�0�%cS�����0_�|Ҽ��J�a��8�CnŘ��;�](LS��C�HRȭc�BP�~{����gW?z��-����T�t��m���gX������G�)r����1/�>ݡ�2M���X�ڟ��$D��lhӡ6�/|<��<NEӀ�r���Y��5���TϤ����U��Ҍ	��.�
�0�͍��x��Ǻ�Q�X0t�5�C�׭��3^sg�%^&����	���r�[�����a����
���6��m��!�a�`O�H\�~��N6Q��.�H�!e�8	���A�:�+����NuH�J<S׷TG,N��947ʇ7��=�ޫ�^�HH"8�U���z��xdCcyHk�Eʹ��>���Ȉ��S�މ�0����5�[�տ>h��۽'k��|��ĩ�W��Md��Fp�x�4�uC	ʜǘ�+�+]��_^���*�����S���6��PG��D����[i�Yp��A���)pg"���
�PuƗ�'N1�����Pj�xj���u�Z/�vu	0�F]�����%�%��K$A"�ưӟ�Pu�� a�^�X���.PUx�z:�H��j�����M��]2��^��ᤌ����ప0�������I#
��w�,�OʯR��g&�vz������C&���Vϔ��!f
��%=!���|Q:�A.z�bE��zdeZ՗�c]zL׊�p��_�C�$��愋��pl�4��&c4�u?�(����d_?�	��N�k�`�!��bm䪦$��1��I?C�ES�w�H�:R{������؎P���%�!��A�B=�F������wy:����í��Fcr�c��V=�Z��uW���^�W�l�����a�k7]�nĆ���c'M9\S{ض�LH��f�E����_��y�Ǎ�@�/}K���!u�o>��RA�2�ˁ�oL��x�U�%X ��O,�y��`�8�N��_tZ��?u��2�!9�p��;O�C�Q�Ҵ����g�KJ�E`�
��V~���뽝�t�3Z�7�q�����WZ
 ,ҝ�=)����;�+�1Rf�W�w؎�M{�5$Og�i�L踆BqO�����jȰ~����5�� �F/ h�	�j������QӴ��|Q>�d�=� aW�gQ�!Ɠ�$}�z��s�d��jԗ���cz
c~�e��慨Y��mO�6�R��-0�s��K�G\�:bUU�q�#!Ыˬ{����E����Y�9��?�ܱ��y�ʿ�000�ӣ�J�t��x��償%��V����.��a��S��}�	P�q�_@:V\�
~4�o�Ť�.�g]Z�B��=ۥ�s����#V�,�I��l#������KO�p�~�*m�<��I��C���4/٠�LM���#`JYˬ~}�/���I�!�f�|�;� '�v|�_ZE(��a@ qp��� Y:����!.SD*�T�H��Y�f�r��N�^P�l��Zèǝ���]-#	:u��9/АU�qK�F�?�&B0l�L�N�4X�v!
���3��b}�QX�Lk�F��&ˆ���bz��u��~�0��_����FQ��;[�ةcW:�o�j��S�1�Gs[X�k�ț�q���ȅ�n�p�`��9\��	��Ͷ{W-:���Y\���;��i�J�Ҹ��*O��R�nU�h޲Ip��g6�e@lewճuL�NOH���D{,����v?R8�^�1>����
�2��a��l���۫o�EYI\�Y��p2���ϊj�FCu�2���mWA�&@�z"=K�G��5$�Ꙣ��A�{���-e�V����O�ؒ�cm� ����/�Rb�z*�uO�0�6����G��n�5(��V�VCQ"�ir��\�+��Dr	YnL��V��N�a3o�垄�c�j��R���yy� �B\�~��W,B�i�>���-P��INp������ ��i�y�}
� �(��Z�Y5O��\φx��j�VK�]����W�m2?Cgע�Ky\��4A}�lFB]`��,���q!/>�q�WF��sE' ��޺Iu�={+��)�A��$��Ur���՘^z��*�|ی��9���^fĒv�ÍA�U4�����rZOS�cr(���N�(����^[���������:�#�gR��`k���/��|m���0b.���RK�����G	b�r�;�i�w�J��gKA�Q%�l�!��!p�F
���;��6#�~�H7�Np���p��n�
�����^�Q�I�b���@nE�#�t;�2��v�`%FU7-��'���:'	;���N aZx!;�SsmGZ��P��hsbgKT�,�4-��>�mhi�uv/Z�=�'�K�1[Gm5f���B��μ>y4�n��ZZ�d�$�3~�-�s
j��Z���XwD��z
5\��v�6�4[$�uG��^kq5�Қ`��Ͻ�?�BXM��5m�-*�OfUj��0Q�;<����+���/���1
���+�+d�������Jf�*�t�i�k��"Vdh�#t�:q�՛=<�gTY�6/���L�M"���ɾp#;GUw,��H=���3��l\)Ci-���b�A$�A����������j���( ��3>m�