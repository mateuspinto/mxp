`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
imsSDiZyjy65Wi6Cm1XJ7TRGWNw8idu+ynPxKEYdvWTvN5YJWrVKqZelwADo+FQePAnyTTD71vyn
tK28QVUrsVEpdbmqFQEffJZSWnIPG0BT+ukIz8Fm2zlIVQNcUMbDWVMum5kfuqJeIqbbiK8rkR9E
jmDvJPRH1JWjVwNx4HUKoYCcq7gb8voDybOzIr3ZvCQksj5OVSHTQoS9ABNYmjKZc5c8h/0xG5TK
hHw8EQGvqvkYWih992PVP/HCA5BomOsKXcnYxbzrY0qbA0aRFfZjlAqzecsDyGtIuINNZOT4tmsh
wlWlIJXhwQnMCmNUBPZv4yN2dq6J4pARoHI/SQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="zCzvWv4p8iV/svfZPUMnjoM6mcC4OSUb+bGbLqEuDCE="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
ntxJn2XSCsdWJGI7qkcqjfbLAUIaweB0QqFaHudp7zb9qiERvVNxMwqZs3Imo6lP24fJfT3DGM9y
0WJ7qZbi8TFk6Fh5XjYg2msDvrJBPrTp64/EP5K5eL93Gyc/2GRf/wBWbmgUInzp4uO5rd6lVjaY
bp0X5t/CquEMc7WYhi9vIleTrDs2QCDqyTSaMcAGFFPt6nBKq6IlDDg1TBsfCqttjh61x/WP54OJ
NTs2vXfazuwuHT3z3UGgY/C+OSWFH2fr+cvexbMRQldLZ/V1NuffaNShP6EAKkdWpN0pWYX7yRfE
V9oLypV8MNpj1ON+QhN5O/ENdFB7PtC7YuA/NIHwnCOj4NykKeAJL7+cewaQyYRfFShEE0S+cFTb
91V1YRQAxMi6hOcqmHLhp3wvBdI8kBqIBvzpIEa+3OMOiPjZ0tP/HKzr8HqhsZvM8fXnrV3mhtwr
fwqKYsG1ddAQiNL1euaSmxeyCJOw27jIOjQ16M+Gf2NPDk722p6/QrmNrwnNwLPhO7GyOhGCIAV+
aILjjW0Klh2r0SPfYAyQipBG/kEkrxXfxjm+0XFDeDqcljz67+Q2jJD4wjFs6e+nyIACzGRxajP5
CW74krNDx+KRxWJaKdnloY+Qedi5yX56682uu4TB5nQAXhUL0QKnkAGGAl6wQVQl6/gCOGzGQyT6
IrAR+Xk3Txii3nb3SyaV9Lna9BeYb9wQ/MPr7UmUMAm6fKOVKE34fr7/Gd9AP4CfYBo6SgHRL9ci
Xa7ayoin2uVbFLxmE4wT5E5wj3I6b3yYX/AdEoUW73WNULFUQvkR9ZxYJ6IAPWhq3C/Z1Vm5/WUB
0TcLfr8eqG3g7dW9Uu67ta1Bs4ZSTV4i3g7K62mYohbeSzGxDHm+Jog8DZ5ZvjP53Ovt6Kt0ptfW
6SbVlvkAAqlGAllPItuypryl0Yjm447C24SgEOMNLU4uoOWiuzR3CwCqVSyiO7Esxz9TBA6A8nsP
trPprj8Bus0o+zG6kdXUUq9Fx+6BU8kMUxWA/s4AXA48mU+3bwEyo0o1eUpJa4T8/lnA84VeK/kX
IffSbZRMOBZMOsI+C5g6ul83gIV2mC4MgoqyHj1MOTpQhgr80hf7d6kz9aPiNQbw3VU9AKWRBGr+
8JZ1cFvqNJr4fhT+PRLVpvVKm6gjQOUayhMs378TCtFAeGbr6qURtixBDk4hLvdfgYnqr6YmLTY8
cNQ0zSkp0akYfy/JqfwoF0xreOzD/zf75qgZXvbQUF6QHpESX3nIlAj/GgzWejQjEUrj95Z5p1Me
qNA4f4xN4hbNX2njrCrL5gtMiXN9wOY/X45HsWGifE+uSg1Ly43Skc7XY3yGJfm6Ul9hTu9Up+mB
cIXmKhGEwB9sLm1coE+xOamjBI0KpgQWCnijnVmCf11yjP2tFJo/plJ+e6hRWBCRCUb+s4mF0XCn
lRDNlvj6SAX32P6EQQGxzrBOt/kttfFeVGRYTVzzd+s6jdjA0dA1N8kUF3Bw6KSPV8xJlfRHh5E7
zxVcmjgUA6pTAbibjSK/aADYXfoapDzh9CKPglKLSCXkZ553KK536448g/P4e4XzBiNvlYtDVSjY
YGNLQBctR+5SCppQEdYjba6pW7U+sw8rmvtd1lE9lrWr/ws0qF9HUOmAl64skXnYRKO6Ssx+t/jF
oitCrLX/iwfpOchrDfK3xK8pA3lFs+oN/u8L/tiTqaQ8jb2KDZvV/R7l/pZgF/xDhM0PXShN5PMU
3h1+kJh6wlxZl0tRVWRYGgHTUDSipSiCYQ3eNwfEFkFwdikxAzWRGAWiuF+e64cC/jynGw410TFW
iSzkHSShsYFbhOvfa4unnSkY6+Eu7PvaMXfvMm48Y+1bzS2t6drC0+FopSjjhMYA/7yyJ5CqXCC7
cwqHaBvBtQZZbvqnecy1wgzMCKCbeHvAgTvALhUPkTfbufPL67SADLx1CmP87PIB3SyoTbClpoYA
7pionbSi11cpgf5WKU7Jlk10G5Q1GkKSjZDNuSQUJqW+rvY+2juos5sn87UD1p3MbPhEjzbXshmh
fb06v/jn6OvnjgI2H2wBhs+C6JR8ybj59G5bfvD+e27HV06BBkIbQw9QIdnq
`protect end_protected
