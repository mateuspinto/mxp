`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17984)
`protect data_block
0mXvm4FG+Hi9YfXhgExicIu/RRZCF7EM0amFeDVgoIXOUERINLHadQ6OKtBiYdtiy7lOuCoADBRv
3lsLj0fy/YjLILbuTZ30qu7dmijD1kMHCSiWjaKnxe9/FaCvYeJTPMtWiyWO2IDTNgj53b3kp0H5
X0cxH4Xjd2JiZThgMVPvVYkhF9Eos30RQ53LkjuAlLoj7SGbnyBjFVXhv3lNBY1UW+lC4wCVT0kt
G0TvjuQagDtCdChGQ4IEGpQiETUqA2H3nBPPTpchDAIYrjwY/a3sIVzVo6DKYcJjlxwCCyeWqpBB
EQaRqsIp7DvcTpGVsjOpDIQWFpT3zomfv7SQbBdVnie+vU/uN9uYmCvo0aizkicNdEu6V/qw2uNy
nJTXf1vlIRP0lmOCvEW3UUyOVC+S6hJl1iL7pz55LcERhL+SC35tWLqCA+GVOluu3Q3BdsOsdZKt
6g/VPLJC5i5wB2aujJFH+4sWx2qEj0bImmqQT8X2AFZnX2K0+CasXM+VECmGmXGQYBVkPm/psXu/
IXcM+ovs+/oswYJSjXUSU+v+kumbF1JOcN7+QdG6b/GLkEGF9t8+6zMDlfljGPKNS2/glqOKQ3sr
Xkwi0PGZ8QMxmRuqGKuu+JK9ArmCesJN81zHlWrwaR+eLun1PLP8ay5DxG1CLl5U96EfjNt+MKsy
vDreC/y9yG3oXrGOfvXj+DEhMttp3IpeKwUWaXYcSM+lBzJYkJmaecrcSv6HkboJo87ydSSMSQI5
HTzxPz57vsj2gom0Fch5cks7qYKfTuSkiMJcAKLUU+eLJ2XQ0qW1veU5X6CGob/r6TKgBWiiTVV+
cBqvohyWiRVl5e5Xqgx7q3XQ6bjGDKx9oe+9s8FLmBfZihjbbmwLMdt7+T4sHCIhe37Ptfb0iUNl
X3arA9ko1BBc2ZatQmXxdHlwVuSOiTlKHK6IlPHlMyxX2j/ON87Iy6w1l7TKU/eiNJqK2IcFtujo
lXdk/07FsZySRWkrjkXCaDkYsP7A8Yu/CwKz/3VWuZUdigx9gfcyzgd9pmQF+nW13R2Rexwkkqeh
IfQnRWHLAjD6MGv4EyQI0sjAI3kxSgg0aQPf55bbCYoGrpu/EGZUugAF3rwQSsZ5yOzkzsBlPgwG
9gz4ccvk9aew0wRPcNIfJjCgxCGJiUkK8YnSYsMWYFNTXg77PH5nG6Pws1NuQKKuYDu1VF9xtZCW
Y+teIsX9v3T++s1jlcaNqUSD3adqt19O/J8oY/RGKdbtfYahTTi9YY7gwpQR1Hya6mcS3M7nEGnL
iyLkgs9R1cF2HDzIA6PtLFn8LEHAXgwO4MbVn8wqDS1vEifk1+lo88kTTz/ypJFc6EPhnf7TyBtI
XFLSzpYI/ZXIq8CCRFKU6cuehz4YjMoOX7Lgp0YOOjNVolPc3YgHl5EiH2JRHtJHL14jX36+gsUE
F5qdhItemJlOuTgAGR3qGPTubeX7zvGB8NpFUy4LN6yD1vdZlq90EyY9FirsiIt2qotOdX2Du70i
FCrAsRCFS8aPOEAQBQvJUDM4CotOrLxU3yuZjV0IKBKFAAJjh+EYMtQOllYu18vydvGMSWyJzjVk
1vELqfP6sm+uZLsHupghU8a5yC7UbbTbDBzfb2GmIW8n3KdLKonyTZn4oUyGZ8GAiEFndolLQ7vJ
Hy/JNmHydepQarz+9QOGSLBXz3dcFe5LVd1D8mRsR6fcKSyvXf/RgXV801hJdVP7LEEvLY2o8HxN
O8DTyoP0PpFu0rntZuA3kaVTzzyygOz3TNyKq2e6U0Auf1ruI9bUUL+/VC2BwLH3SEzSVOumCRXw
RceGOQF0Lkk57mwfli8y5c0vWj1gbJkkH3iv9KEOhuDkAO0DGl26kdnYkawbxBzVVwqun8ehCE4S
mz1tuzwiw4jlUs5iTIkda/n4FVwfNWo8cpMaoDR3JbX0i/SAG/RcNxykEdp5Yb6EEvCAJfq35eiZ
0NTkdoo0KbI+kZZo/emAfiNxdw+y/LQsowrZGTU2cbhiG3Etru2ZAjmpH9pEX0Es5KHCYeKZHMX/
1LI3egre4vKdcFQzNsx0FxU6H35On8G7iBGN6w8p+nIMTr9/oOVQGTppqOrTQxXQvcoO4m25SWJD
bYAYffURTS6UfdLfLoC/D+UHP3c2BzkKPUv0R4Cucqm4spCHZPlvFwdHn6lRJfiTNm1zOiZKFROD
4/2wShQiUmLjBNL1re7t0hOTRJWBXYlYKtj/zwullFp20Z1T4KMlLAEUhVyTartI28zzpGyaK8OV
NEfRfndFuJ7k1AbRa+SYbbvXvd5tmqyZfHKswkeMvo8PyZOUjcIQVnjnPaJxe0BESxcx4y/7vv2s
JzshHlcSzYZXurbuA0gpLKAPRO59FKJEXg7/POq4qHCU7BCB0TW9ll5Xss3OgVZBfuwbKiBgg541
j4GXtrLg1PgpMxGQLrXYLZ/Ldsbo18MVVjNPy48lNXEY8QmtUgFIknUF6IIMNfUKtVmvzirDo1RM
O3NT2eOMSb4v/N/2+LP3I2Nc0SAt6Vdo3Hun8TpKqNfzPZmPGMYVHNNrcH0z1vJ+ZiylTgoO6qph
/O7/ZPR12jmT/ft0EODNdVVwIWL5VTtnXaYNNsjZcy3YICf7ty5vS4CIFkpL0MvL1aTWjROAtbFw
D0uzb5bW3YeEnRCX4ADfkqy16LaTZOArJPOos+W73a0rUlkG1N0qe85Q1/CGlSmobU1lYRNlvAlM
EWEj9NyhYhDGuyuz01WQI4+19TvfFzGby1aDms2BvHRJuSrb3cQuGztqTSrfOFg6v+EXKjrR7uBl
CKLbZHxFnEM+tiqO+HANf2WBZ6KVVpQuqLTuMbjAH1jW3YCPt7ThZsvJtJ2effkyfsbKB0/Lef0n
8d8/xfLR4PsKa4Fdc0RG7IMlUuYAekKFN6XVXan0acrB7mUh0i6n6LeE3SIo6FegQm+shPaLujpR
QvTfr+i//yrEDECkefOWd11yOhh2+b8jtTq8MDsi3s0nf7IJ89OWtk79I3KAGL8glNNHGVct8J6V
lwKRDblUs2p6zgxLahyT+FmRWmZX3/2CSOGceIVS2uIsLAHHLK1b0oocm3OQeeLr86xzTQ1QFXhJ
36ZKZZjfjByRt6TdLAsQhXqzo4lX7BfhC4klBEcBHjLBn4C+l+uHtXjpjWM5kGJe1usJStdImbEv
D+Vo+/0d3CL4TocPgS3JM4EbebgW8BEU/tyzII2mgV0FQ5GxMX8YQzY66MdpWTgwKF+n7YRNQ6u5
lrQAXDgfsv8g8GsxoDPZkC2z92gNvEIE6+5YxvwiYgmYTOi5nVMaI0LoAGTzWxCa9cYdiTLhJZmr
oMVZrTWLZuspyk8U6ddwORG13YO0bDCqDDBrqYKTe5zTAY0PVfN4xjfcdkY40D98rTMkgbMmB1Ty
19RLNKFpza0VVxbJhMWk18XFjHpFxrueIhgp0EGHD+ufus8wMDtwCexi1ta9y4EdZV+h1iVAU0X5
RJxaD2ALAjxRUl0lVI8NGQiuNF3psAavWdkQBh0Wfb+LPJ1/uzXXDTuFUts5+PKZYFeSXylCgXtN
Upsc3lScFWCF7rPSUZtOn6KWTJgg0LfvzhSkfhQ3CUifixJFIPVOh89Yh3i7uWpn87RrdDvrCMfi
r26fTHAzy7wQ1WV2PA0BeYW88P3HfDYSGZC5fWcxWXvT+s1htDlNDeXjUbYIcMHHD48pgzs7tXWN
HKdagYHlJl/U2wKPK84a9pJYBc8i19SaRrPPvp5W7eBTu8Vby51Tw8RkbMzBSKN4eUxY0vc22lZF
jA1QV6AOfwGcqYWLdEO+/7FI+DoTGllFwGKqjpViXMBdZ8aCuiudAuoLAFwEZmxwcrmtZXSQ9Ecm
jOyVIh6HbJ5yVTnfA000Tkj0cXaTLbhPUbQEKjaUh+pbruPPXa6BOkUU6LMrRJPBlZBA0Nk7IjrZ
N7JRTDsGWFl6Y+hydmuLMd7neexV8VHEF7B3eGKOlEqXf2ur42337Sb2R3ra+kfWRTQTHq/ajoo7
CZJtdSi7mbii1CXEbJcunxo5HZd0F3yAvZ6lFJBjgaNoj9OilNGImqg6s+LQ7JV2ZqryKeiX5y5J
FMS9U4mEtoXjLrtaOQb6n3T+/dzsYmAnav3rlS0a9aeRcgmvANu/BT9NgBd6wlge33iTwc5QZwce
SONY2ASOaPGr3WauwAgWsv9ESncksWyf95bR4E/go/7BRG5QYIzY3QySR8TBqU6pyEzEBD/TSLAL
M5qwy4wkFIRHix4xEzDRIk2/8dTR16ATr2zPar9pbAUC2nPjQDu2vIXJa2K9gBLOmqQHpRAIK5LP
PAX3ETR4JQK2pAUoIVgJb3/3IkUpUsT2ei+/sW4q2JH5dHugIXp5xC0tCDt/OGlNl2JJTTetJNAJ
DcwXZW+ihYOZK0RwNhp3Pl1fwEMK9QZWIAnvf3yBJntHrE7JQojldljTkkD7gNexADjO62PoU9FM
gHd9lLpwo5BBXisaiKvgeB+ItmZIerK/namlx9MIzTjcw+iVTtKBGOMbiDOFVuhOt6Rw6wqQ8lVF
Ve/sJix23Bj4IgzDfgbtX/vpjEL97GsM9eVRpHiZzgI+yLArjGiBN0VMYzhSrmUBpIGz0kmNEgZv
i/F7ueE/pxEbBrJIPV10bI+PMAlAMCVFXmhEIblxc5Gy0eEBsUhIUTXZm2H4SB9Zx/z3lh/BQAKW
MvKpu3DiPyXtqkVZuwGEFjOg9mQuEgvT7Qg2no3DFkrNhfnzpsUbTceWXEwuw+gSuzsP8+5xC49V
gXBIkkdtGPaCV7QgdvS7LYhSfUVbx2t9kqRFTpTeji4AzcrtZwwS9PPvDY00zHk4bpJ78VihHXP/
L9o5Q//Zhss+PU+Ae6fHSyvEaMEgIguC9h/SCqVRANfz7hRQgnL0DHCUDfTEGVaFBrq6H9+JS7ru
2mPRLfXUZBSAB7X5sWs6fhCHSgU43GcBhDhYxFniZfPfbx8xDDamxFu5E5/s04+ZXMxgX6Z8d1jG
o46+5bZ1oMbiPBQVCJ1l0cCldOU2bg9n4elKnhqjA9ufxJTszQF+NwCxmsIBo0m/VhJ53VOoVxV1
EoyzCmjhCnmTYQGGuW67HI9WKmwqEcFM271pvg911ukwtdDVIDAGENGjBgrO93dVikA45PVceFuE
gJa1pQ1lMztKJlgr0NuzkVHuaTkva0/AGzsdJLbKDLVCr5hYuo5qZbrUP3Dh44+GCAC2GQ0NBVPm
/2HPA3MhCE3DfENoirRWRXWUzTkrlUdt4frUyH7UA1GheaNF19Ii/zWmCJsjeohwSpasaQoXG9ij
MHMd7W7gL61PyESY7K4vsP3+HGepy1AQP+nGudhdo7DV8HlaN0aWbJnlbBsFZTcfUETb4drp7fhD
7neAs2Q9JYrR8RSC0VlT2+4JsZwJWTiKpGtl8Ft4bslHYHN2bhDyQh8HyWJ0qrdpjQpFMJriCfFx
ggMrUkMcrixchAc7DukLQjbsvFpYNie+6wq38JDxcMjXS71WMAeB+Bj3/sAJ+3eA9bZzyMcMe/Rt
MSHTpKF9VQiZpsSJUnirAO1MnlzbgewVBjBb/zRm/xHEMAenajNXFcdbP3vyNdcXVirBVyZxRk6Y
zWjv3fsHsPhrytMuyDOGE9RILsw6ZJ7yqAerENhwT3nr4oxwbqXtD9uB3finbR+e3TPcyaRe638O
RJm6rJ6tUVIAz8Irp9QsUV2gpJdQqI4kN77h9/VGzeSGqHsUEOfH7eadEjIEahpXBIxbkxV76gtW
dLLPsWcCXQCxSqZK932EROgtmXmb9hiXIBU2AuiDFkYSdZFtCiDBOZXH7lutWDM0BPEawD3SX5+9
tWF2/O0S1DSouulfpga5E4hGm5dQI5huun1qVZNfHkYq4Nbk6E/Vc12h134P9wx8uQY7lo24EgbE
IymCNIn93NqtZkzxmsWgLOnY9wX5ITp0LgSrhWw3vg/uvk1B9pbIx8nz0M8h/XF9s1oeHiX7WNVR
TbuDWm4ibbWA7EYnVu+EGKyAkVxarhg2FJNM07Xh3/CFXFLNg50fyq7yRaG1NgLBf+pj9bUtMose
sy/FLkRp5d6LuTNJffELd7VWfjWLYmc7JUu/gQHmr0wLnQzKlNhef7aw3l1bwiHTAke44ulY5ysg
aZHQVVT3ZTJmKhtDLWMhfaT5lDP4SbGSmtJwGifAUok/N1/rNiwY9OkVj41sYWGrY6LoS/VsfeGP
GfJEN3liXIp78MrNPdavhK0qsfjbP4n9wAifkqdqcLV+Ajh6/qJ7F5QqYlYbVXhX4vvfQh/73blP
JN8bk4aDu3C9Nl9YW2t+5jW1JiOoXOMRFfzvqMugnOrZmQMDxdUInyx4XvYoD1RUB9kC4t+OSzQl
En3qPe1rpW4BEgD3XEfT/Ip8QbkpKsWcbW6XJr/m32skQquxnL5pvN3Z59b4OlMJTqWMPNjAftpo
QSR10omD3b+ukf0w27NlCU9D2KlihW/Da5AwLb0/4+B9BLDxremdYOjgiFxloWfBGMuzAUkrnYaY
I+islVYjAq0/+iq4zakK4J8k93wdRq6YA2bw1m6gD1woQfq7vZ4CeJP6h5hCMD9WYDIA1LjReqRS
UeQptFcV5LnZDqamYttpOoyVXEa6q9gB3mBdZWtrzKwQhAQu8F0DpsUbDl/tzx7kt1VJXBrPpTzT
V+cDjzJdCrLpTmdanB3asxcZhUG/0UysWzqjLX8/T3Djy0JgdhEKAL9xTV77CcrnUeteK+1KBtEU
A3VUOakT3Zo5IAxeVkmPSa+NTqZrcoZgqfG9OmQLlAe0Wr0XZUH4OLPPQ3epQVfpCo2gpHbCbdj8
d97MTyq+p07/2VWEBEHJ2xSEx0WYPDeyYAoG7odAzJBno+nG6GlhO+Ev+FQPQPC61pwidCwTu6G2
un4rGRxKc/kyFz9V6F/3slfyXuei6cIP5NvWapshO1rHVaRfCfTBoKo6WKjKkcjg452E1uqnmvui
7VzvpSJJP4fHP6JN7UmgOGwsVK/TZDu56DWR7wY0sv43eIRgD2s6KOHT3WuJ28dNUY0Lc2MJTud9
M1eF2s2GVGfWwmreNqp8H/r9vbyi0rccW5XoCUWLxvqB6tIT3hrrU00exjC9uFsJnMBbxbZXxCxz
1gVsQBhp2LZ57WLrdxBX+VOqic8zue/PWwNpAEuQpDMulSRDsGAL2WurtL2kghdxLBJmes/Nbld7
+RU33qFKSaBt23yPM8o/ZmeuGQ89wWFoZFz7XcNwgXbHTwnRt+0k3fNmOuVzI+9H38jU3ngKyAv9
6cXFrDazLgquYq20/Fq96SvcBle5WRHx+x8Vi/y2rlrhv3hSTHhVuNqnudt//DHiRlRNAwXxw+6+
GSBXhXL9xzwxjI58B4eGG90IkuvvQjhdVV0D8f6Gb0DZEHG04sX8XSXzDErmr0nyfZWe4fns0zrv
5kFJl1cL1vE37m0FUr11m+1EwabH6SX2XHhWUZfmUm0YzvJstg03lJp4ET6RcrVkKrMhgN+MP/1p
mI/Bixn2/eSR7MppoU6prGHVOltDesowr2XnUnNkPxaZYJMZwp3mDrTkES+AJtXIXiPseWZkNU1J
+lWnHTADQitd6kY8Jyy4ihajEPI0a4dZRKtMEFsAXR6w/NZE5MbNHGSmJe/kKKrkOlq1C0zbfqJt
GPYlXdgYK8VeQ97kp9YplgD+w/jp2b71Ew8GTFKN4ycc3ccTho5vuJDHVhL3Yj60f5OzfCiouL1y
BYhg1uEiu5hJr4w8dUjF66cQQUkmOfYsdnuDz4c2N8ewjuhvq5EnbKMSYKqTWCUQ144ao8gC2vQo
cq7aw2gPGCRk2chrQ3oEdLOs05XP6+KcpyOc1WXLYoYLK1wsR5MngQjbLbXv0nLPxAiacqxDQL0i
j37Zm4cvBlPOdCN2AzNWl0mLnpUijIG2WA/xA6cmnpUXDYa//TnLUAEKGY6Pnw9Xq4co79CpwCjn
HhNxaWcjDZ+5k7bz/0fsbac03QtzQvzJmumzX8S63YPKOVKFJLDPxAqEClLBVB7VI+wWJ7pY4XGm
eiaU6SOLn56Nf1WKYFydMWzag+w/e8BZU1X++LSRlDyCIIEl7BILKu8P49svOXLEd3Qsq8bjF47j
lxJbhrCaTxo7FEwUo3glzgw5KFdLCN3e7JT985iPfjYANOIVQdW9pj+tD7+Hh37O9MOR7+yDUOGH
hH5pTNi0hFjyjbBxFHcGJKL7y/ReFcXirSODZDHZbtqfRBJUQM9yW34MNRYo8Bkuh7f44UP3XBl9
d4aqMkczjrSgMwEOyz3RD8TTcwJH8qaPbqHkFGtsO8C5opgj+2sWbMlxnTDu3Hi/7ttdVusYzeoO
lei+x1FkYNhX79KOIZrOxWE7WQ+wj4xmg7HGabkctpoPENApWECUjT1khQsfEdoAHKFBL8a2qnJl
PbxNZCLd7NAAhGNeXcgLoXucJ2ir0M7nER4v/98RxnN0dcnNuUrPec5d1b69hQmwmUWBKUKOeKbV
XHLvDxtWGY+0Eu6uTE7YsKegdBj/Qen7Q51nklbV5Jj8AYpFh1IlQe9T5nDxOnYQCEN3oiJFioDS
dbKaBJIvwcRpdRoweYJRH1rQrmwYznGlt0RA/3k3iBIPJNSiAiA4wT0SwFMz1u9PI02zQXxQKW0W
BGLgPPyY2SK3MynAft/fFiAKZd4L8Z+qU14EMHf6BrBoCaBplkrfNF51AAltAlh9xQAGbn9ANYAJ
coC0e19Am1Q/7b18NjQs/XSlOqPHdvzE25iJpNJpeiK7bj/MwhoBd74/wXl930D5fRL5KpocVNYf
O+Ge3sdkECGhCTFpXt227mzGFr0Wevg7T6p6z36SkUfZBYSi/Kffhmbqo90XrWlBTYImlD50O0iM
4SNo0CPbF5D4VDYhDvoEcs8vFc+N1mepChXhyddPVSGH3IEooRcvWY8L2zl8bSSbBdliVbj4qWKP
p4A13w6AoTabsDFZ7U/QqLijNYXLxMRarBGTD0KszClVx/UBsUGHPchKXAQG43z0JBeD7Ni9WJZi
17jnsOJY/xgE92Y+9tBiPERWQpcyJw9MFWDGopFrp0cWOHrJCsz6gtRHjjoGFozyfyDGGeafAM2A
DzNiyv/Ui3eAFpUpiTJiiFsAaMdJKufNtcv318uOuOEw4OtGfkp1DkF4XPWlgkcqa3yNgbZXfwiJ
Es8MyFQnd4NJ/DJwhTvHRwnTl7/AdG5Apse1z4zeDp1c9Fk3N/+z8He11UPwsjuef4NU4omkRPH3
l2lZbIQvsgtRGH5iIhBsqVfuxy6oSfJZGXn5Fjvr6fNkzxtGBZ6HHMg1ShpEUifw1bKSUQiLRA5c
lPfUsvwooVBa3ZwH/WUOCFwNJPPg0SCJHaWq4X7tWwbVmpE97+KzHhzZg6yxX21DNE3VKwK0kruj
4i1JeR44jSel3rIzy74HXuixkIIyJnFNQdRw7UprFbVGYuAOgh4Lk9kQcSzl+UGUztn99o/taceH
PRLBvofY3bUhUT0ZAhlLk5wIIwZClyrllNmczpewAzn+IJfQvyD9F+lDrd4BDG0bpkjf9Q+2brqR
0W3FH12JWtmEUL3OIHTYArSChJjm9vJ9DO0aa+HCB1qoYcP4kmwr9ffr11JSZlbSuk+aAjmotHkM
rCzvfnT0b3WtnoCdI2MXXbmOObmuQgVxXgNinulcYwU6ZDStrqKBZpCWyW/SY2s7fM129YqwfEdK
HkWlVdodN+qzTdtHUzIR9C7T3rQ43b6Evd0JxXDH59odiDMvekaXP4YXv+dlQswV0Y7EjHVA4SQJ
qdgFtuwv1dcNW2Sp12e1HX9oI6fWWHaAIlzBDkv+N6UABrqFeLuOsriVVOR4ONQaA6ZA7pGvG7HV
WpcXtUgn5l6Ex0xCZArRu4B4jeJxWe0ljBskc9iARijc1vtgcPQTGMhoAg8tUiajO2nUXK140d5K
LBe5IkfuQAfTik4FJ1BNJnOJQ+VhVX++tBZTifCVeoInMeR1bqVteI3vvpzJ4PJIpk+imjgTS3WS
m3QoeaxBXEmKiveGZNB+y/tquJ5O1VHLWHAhwqdUU6NAQH58rMjyFSeklfqd0eEGvFh8puGhaEgF
QvCzbF201v2KvlLaGKwE8djtwY/FS9ION17Mrp+LYc9HUH0LeIF3RlKp7Og99V2y9zzq/mczm7FH
/89XEpqLvSB9KWQDtQug3UYRMLgnhXqZI6uux0LF7sDMByWY2UPLLgg3GjDhtaNpmL7uXbup6uge
uQIT8c3A/fEtrAgcRNEr8c654+fvaZINWyQohZsXzYYAMEjEI7ggaaCG0AIxC95b3HbsvRO+moDK
PusWpBD1om1iFgfPtvGNudGFmhFlMvkrkwh9tGzokgnUH9b/9V3ziCq+eQz2hQjuaGlCJ710HZ/m
36/07rTxO223LsWuDsoDIz/iwDKmrlx0n/B8Eyq/5PDHjEH2AmwkcOAh0IzoS4IKGUdKyUDYfDRK
i7Nrwyc0bB6Ikc9vveXZSGAH3VO0dmgUKeXKvdUr+5Wd7N4lH651bYSYqpNq9rsNG/AJKB/o4RWi
KQQHDcoBG3r02z/+npSpimMwNASzKH/dzCLA+5Lho2bkEzAPUUZlFxR93foH7OfAWEeIUJbDa9Ip
rU8rkyFVHL+MitHBZ7qKjbP6GmJAVfgstbklgjdNvrm6+FdxPX3P2N/2WZCM5Z4TvNrbZF/TFiOg
jIvGZJfAD+U0iJ/daBiq6Df6k7eneLpVRsbDhQqGWBBEOkHPfZD9PrFDUY2pAtVVm60Whx0RY3w8
7pN+28UVlDQ4HJixaXluCeNN4wGGNviXXt1WJJwQ38Pl+UHS1Hx5HCqPdh4PHw4QIypY4kfGj9ju
VvCUgHnf4Cf4Cg7tkHOJYg1vrRase57h0ju+GDSsvGZqSwfd4BN1mTUfUvxZUrQ21jlCbVxgUYx4
iWgL6H/ojmoIWAFkN5z4eJl5GTpegSuA3/5e6rJ8Xg6Q4TGc+rHWiecztpJXDwvizb2xrYRa8x5W
wAjOBbouooC2S6EcJzRyFpIDzqz9wN3qbWEJrmrKYB16vrEKmgsPc2RloYoNUSki+V76hDddBTbp
0F5jsoSRRby/4MAhwCgeypbIJuX2pU6V1Y0+thJyOvYsZcP+1n5qjF/OCiRRV3pBkEVOG5nANKWU
tQloXeAYkb+jsYarpRtVwco0d/ygehwLy/5wn4DsTuybC4ESP3FOB7FlmYcWTxNyku83qcLdJG2F
yy+FJuM4MHVfwSyAxd5uY/MNjmzOWiug3dmebh88Br7fDmGQmBC08sFv8QVWpppVyIIT0GMARV5r
vLsUHMraCSqcToZL0kafFly584aTmVBnepJ5b3WNzhYEjLLED7M5gQeGLVL1IYcdmGfe02sSTWqG
Xrpdr8HTSv86DbQzUtC2Xutl6GhLbgA2gjM4eqd+A0mKpOoFfHzvsC5SvNp12tS1222yUcEksg/f
Aw4iZZ/qhA9g6DpOwNV02S4QDfBgVxEtDtMQ3Wj3TRU9LMhUea6uY6gtToFBlbGqexQcqmGHlJig
QGgcu1uF8HiqaOxWxbg0KEGCxkuQM4vnR6klcB/MzlAyxFdD7wwyL5fSdqqsktb4Y9gdE3Olo7Re
J5tqMwl5zUj115uBodMg5gTNWHF//hNcmFbFXxiB8F77C3GQtmwkH9JxUC4t+Px6LIJDjTimdBSN
Z2cIVjSQX/xqBBsRiXU21maiu2cUCnrFcMzrILi/lbef09Y5lGWsDvrAp6IZgcmfOf5iQFpd94Uc
RAzj17PuXTuZLcMtygAV51QXeDHDSag1Ujop0QTyvJvjbYxsnndh6xPhQ8ydk5+hiTJvaVuP6DbC
I3TT30SuPln6m+xOllo+nXwuwUupRjws/j81EQ0wqg1o/uaC6314oY9jcQA7x5+3830OelryKP/B
Xxd/3ytYCUYyAf6G0URpBinFh6xuxYBw43TbSIfxzS27Z3TU+6VNV+1iW+eogI+JUvVyUs2+FpHy
B6JwZlnvsLdHYMDLgkbdtk9JFA+g629fO+Pen4R8xf2CGw+ahiQDPBar0NDMOTxiMEq7uwrq6y4D
aFRGwUzd2B1T3Fs32SCk4IN3LjBfpBv0AXMYdDaxODJvQLKrdP6KrL0VeHh5bnpf0dgdpvADvNEy
fdHcStH+U+rAhn48V4BIN6Adru3Cxwnf/x9yalrRDfX/+KjnwLON3HfmBjTlBFx25Vm2YTx8C072
1iZo/FKfoZHG4gNS/K2mtOp5K94DM11IKLUEYHhQgbpBzdTcHNxn4n4GgRoFA3xQVa8c+vRNobo3
oJ1shJi45G03vHc7zFL7LvaSAfedT+ZYqsC9SpzLgV5aB1x03K590pMeYOpzS50wzX9Af8YvvoE/
MnSpYlLyRB4Ol991c3LQZz36TT3+DSyIbFEmX+bLElS7ZOWks4e0z/br9KV9HM0/5ww0KNpzbdOU
JShbKm82e3sqQgKIRiACoXP3uUZ0ehpKDNiUs4nc7L4viJc9lclAGLY+KAXy982fnnqrXAZXrHX7
6AnHP5+wzb7lbeRbRMEgFJ3ZDRBYAMmFY0WcZIrv3wVNvAgzFC9XkBh2/zYPMLmRwdP9iDxULcu/
5IfH491mwh5+KGS/YutILIYKFwsbGLP8+arlOOjGTv+PF60buLg8Oud9yw1vPRjL0EJ5Gpua7DHY
xPze5TN6fKomqBoBO74qO5DjmbXCFqv8S6MbZ3aTxM//b+4xavK+MnDfOo5eqRW5wSwS8gPkogJb
3g57q0E0mJDfZcYClCcjCl90oPc/aOvBOHts6DMA7cMiHva3EqocXAY/yBgW7E3jN9etnkcdvBt+
gi7ME4+Dm0MMaof1UJjEA8zuD3/gxamsH7c/j67inJaIngRUBjazTTm6X9XTcQyePfn+XJ4HpQFm
4b40WUA1D/8RFUZvfAeQQzgLhz8Go1ZMOvb/YrBaGSWr9o+RTzsRUesBFyhI0KoFG/FZ78kh6zuC
YTyBEgmEjCj2q0mMWMtaxiK1Jx8/ms2O2LaD985iMP9IO3/nGww3gROFXMZO0z2803tEzUJg7W9Q
kT7KAiGaNUVMYpTo3yatMs6ZWuu8+Tq9PQSAecpZ6po0fmqkBSMl0SNfBDl9QOr/S+LMT7IA1ekp
iJnHJQBMJa0xXWQ8HCL5JP2YBGWxjesEn127eIL+iWbwnGS5vg1W3RKBQ8HnRK5wPHcFc4ButaYB
1aXMgWx4VReA+yMAR8ydSVWsZQYiSPWf2P7kB/v1G1a9gNiJXV0iTdNDYCMxDxNErsnswVQ1bOj5
1TGcYFAQU8jNv9cs/aDWs8XDP7DVcMlGvMLY/7ykpH5n/tzC6dnLI9rzvhXbAyX/oa/cbcAK4J3k
0FR8nZQTeFQPEgEv6if9wmI/fJolGF0rpl3n4rH11WJm1KZLypAElD/s5RPMpRUNRe8fkTYLyXH0
i8a5oxs364fkeAis5hcJ5lC0dQWhtqJN5h28MG/pjv7Hi29BbjtwPqx440CJ/DflWheENo1As+Oq
I8zWKwJDmu0gsqWTAgHKTS+Y496+1slN5k0aO8SaL6SZyLypXOLaziXiSmRdiIrXCqTn8sybMuL4
lijifQ7NlXfedwbnQ6NQyrqDFXkxdV9qQZH4VbJqWtlbB93UjKP4b0YNwcP3zTJNa1z9uj4pi7rg
IeLRy6mer+Zp10+Ciue8aEXJfHY7rt9jtfMnKQ2/Jc8eNuUuoDX0DCapks05AVM1iEac6dr3/CWh
WMchUC2g4JJa1ULBcUNcb+kwFLSKF90v6g1peOz+6+kSwKAVPSMGdZ0LlqT+XBM8lPFoGWXygxhP
oU3/evWW928NcYIOlkDMwrhb3I9eCHc8YUdOO4j/deDdHX8DN+GsxJDPWWeYRYxPEffGXnnk+n+g
eYydPBIoWd1M4vOqzPOTKTRDPaFSlY0aL0CzrF05sfhZBd+MZCxu3Y0jbU1u2O993MmldesACsAZ
pXjjgR76KTVb/OkWOV4Cl/+3u5P1MTubL/vuBVHH8mZSIAwUwDXwyOxxA/HMdGxhA3Nes3eIdzLu
mOjdIBZ44tfPK3CX9aLVdJyw9sF+hQ7FA5/+1nlwxLV5aztlbDbMU/dNQMc5hvmXTrmp0vGp+yLJ
eJBF9xr+dufM2r3DS8VjGlGn7FtF3P0DSF8NamCSlIZXSNXFo8x9Ud1rKee2GvqkRgOuy/qDvkfu
jBihNwsrr+XY5GsL3PqfFzmZX0BX4ca30cX4g14aN+hpoJu6jPW8x0QNMAnVIxu+jpqlJh2Sv569
YczYbPUX1mhDhVmnEGzj1vZX0XR8td8pfOOijb0rCLnPIokwL7BAez3N6I4bU4yzIzV/pKvV9D9K
R/7h+tAB7NngYo50usApgSvnbw6v6tFDxfArzlqivFp6BLcKkylXqd2nnDbf8JmcEXSsQVGMhyRX
IJF0n458ocqE7TI+7dYeI+8T7yASQqDoSff27AKNjF7J5F66y6Yicckbata5+zzxo0svFj0uudn/
GPicCLp3TAEa6UDPV9Cdj/sMRVcCwoiK5rYuXaTwnVnhZLfecMJ1qD9OT4hSHnhdFinHSaURJdPP
m3lHMyXRphR649i9bGnKoBK2pKG4I119l75GHIbc1y5Pq86GRacVFJa5zmaDtRNqlg7UEQzkLo7Q
N58LTe91VXjRQ1P6YCMwPSK6VTnWsbxpYam/XAp37wRITgB4bxMNC05Pj26Jh47kzIMsxRCH7ZpR
wnNRToNr/KELbvPub356Un9rnmPnB8H7lcC/gc0go+JJq5CxRU2FB60U3sKDcBVD9jSq5McDQQZa
HXw5uXVbAW8D8eHA8O+/4h4/D32cY1vtiqD3RPDmioJzxEyPq2sWBUrXq96csrCqwEliO1bKDuvw
93BGtbF9M0EL1+3m7BfeaX2JfhP0bjwQky0MdIz0xurFJ77Piikm0f50y84F82dXFbwNtIEuVbpI
eGbLThqfN3PHOdxkILU2Tmg7sYkspf/CQGALpz3F76fP+NCX/Yw8Nu6zoA57RZU4prv/6W7g2i1r
3GJOVuj/FN5ntKRI+k6db9tSWDUfTCkcbU8shby5zodNNVmTmTEi4CQM8UxeUespasu79qjqETRm
u7T2DgZRYFSCDZezcuDEA3Z5LF/gK6bUTP9lHmgaEleABjz7ELVtm5uHQ4UHFBLPwMqIVUTs12de
lhPaAekeMUc0BG5WbTJEwz5XYpSCMT2fdzMKTr8jIkTizHm+TTz84QDxIfcnxQbCIzvj1vr2TxWh
JAgCikl0G7A4lQi4frKudbepA2FWUjXhZYIVfwQeYRyVXGp9X81UtvGwsyS8QVVWd0JaA9/i62FP
aFZio7hgsPUBiTkns0i0xeKN14O/2aEEqlRCYaQEmTiMAKEdoeT7iw25OPk/sopUAQqQpnXcGokI
6chyUTr9eGjpvu8EZdiH3J2LJjbsTP6Trj0AebEVYuFcAVMsyacZ/MTK+7uA5AXCGAO1pvg9OsI8
XO2U8r7Mcej2nWJbeeaRwPjxXanxeQisx8VceX9h728eR9/CilWYSVdvK7HRSkUOrRjnsegTvy3X
+XhrJaQh6hICtjJdBemafh0o5hHwuXY7zf5Vv95K6Xrq+ng5Of3mSkJmjolCg5hG2gmzPiNycl21
U+JPFjRlBaRXiaoZ5p+LZOejsCcbLWUP11foEJkwBmICxoGdtmMne0eRRU6Osmikg/uvonIc73zz
obfCHrrrl2Dcg9IWa1/brcaanH1u+FucjNvw+OdjTT2aK5KEHau53gh47sSPSa/pfebO+lhw1SZt
M1Ev8/d039/ACnHk0L/n4FE3/S2+WnpXtZDt0h6d6dnYES//mWoCCnVDigfVjThaiFfFRPWD68vb
/qQgVhkuL69Qxi0hwEkF+Y67xBgl90aX3M+Vk/uNM5U0t4FjhaYflTIYNQutadzqd7SB/VBLnjpm
VJpd8DCW8Ph31P1OQLgf8DfmjrcLDZ1gqWTHCuExTmMUc/3v7d8WudHTwOKxNqNz1hX/kp2T5E5u
MLMbWxB8+ndm9rtp5nivoX6xmNbydGxHgNm/V0kk20EA7IMwVtemLwh1jdILkq+fc2sCZd+FEPHp
rNMpJFiNv3KuppNUgUuFCIVFbbQh0G4BybD1UYFFWdjcW3TVnJjZF7/CCfF7Y282D7H33gqRpQeR
QXI9ukVnGb9j9eDOPzetJZ7OdR17DzP49P4nFWYhg1GW1TymSTWZc6vbiXyOVZoSuKPYEeuWCazM
GVMxYfSjFPGYgmr8MmqTnjLW3Fwxm7FT+RlM33oqc/qb6Cm1sFilB1XeoG6CJMmWvRBAGinWjgx6
FF/1QuszfRVlRtdIjU5imVsmj34nfDZ4RaUn5AXXyIg6B3R2XsqgDLsc7uzzwa38My0PGzDocaLl
cM0Udgy+Ys7MaCjQ9Ny+1CZAzwipN3QFvspI1R1IV2SgAhFKqX69qqWZvg/v256cWNWzzM7VrJqw
U6uTtVDCwawXn43Abp/JbrfmDNEqMptwgEwYsh/uyBD5tURn8OZsea83K370LWGmEq6jVp8n1J00
EEf8jJDPZp4SIScN3rYj5jfe31Cfatx1KSJG5nHg1os8e9e4ZV2nKeqUkb1KxfoYW+e05cLxTtTx
J/QphYkuSuE6Yl93jp0ouZTb8xIJyJBpt4Gu9lLDCBa/3GBPwn9GNIvRndQYqT4uCs8vFM9ObBB4
06h7QD2FIKfXkN1ko6ShHrtrIke3zaw7M9oH0BphLU5I4YvbPWfItcCBsL2DgRVOQ4sFMAS1xuFx
x32pO3almfqRRS2IV9XgGuBRMFpiHMpHe4aNoqQvokljJxOuhY5IzkAvsHycDGEuge69HMli+Jlo
a8JSSsir55SpXE8TFCvv6VvqzNttqZIQrzObhmOE/NJJCCueNdaUSupRdwJtupceKmFkMMILrnX6
eZ9v+ie4tCytDMEdy0EiaPWzHW5f8dp3q4/KGmug1uiSmfqd76/QWYCIKIMPFjo+7xpKoENp0NUj
Fzfo1GUvhjXaxuUpS+mvMrP6lEM+ZiyMYIqkBrN5gUW6ANt/GlqccmXZK7V7D06nnnIjgDj/KOau
XKsEFgv5yBmoN8qmoSq8nR5/HUcLSXrzvGAvguDYZe+kq/cdMhSSE8c0GCCBfFry4xbWJstxKHrk
KEY+yMCMgnWqfnEgodGnZhXgjpgLhfg4Rqc8HxWgUKHTT6g+2N38eDWaLZeR6SFHdXehu7DGILAD
SiTxwvqfIysnol+Yt+3qwoJeDpEf/N5HxD4+M2OnK/JVPzhE3YUVbLCCNhFHEfzDL4hljozNqSLK
AeVz26Oa4Gu2DmztIoBbf/prcvym6SRZpnuwZAWKhYpthjGr2DfqlMrEeMcLCEhx1PmD8Z9Jd8Kh
ceVQmHk3k7fZb5POTfA+ctuTyWv1Kwh/pMUiuOCa14aUXsL6DMbT1q/Pc3K1rGmwX9p5THPL0Ngr
9DK8WMsQ5//aJgOOY/K3/ByZMP5tGYDbnNtDAOWoUnKzZlXm6CeeNpHimcEPr33juEhbHDUh75A1
+qc3btW20zBJpDWpVt+FZGkvR2UsE2D9bZnjlC4Qcwuh7iS60Zu8WIxhg/2skIMamF4RSRh6bha3
CUAVhhcWOK+/apcAUxE8tqLsTTZ3VJD/8+BEffANkQJG5bKqK9lW/ykIgb0FtN2HbDrUv3W1s9u1
Ax+Ky4WgDmjeDFSlxBvAZ/r1BFmM2qrdpHLOGD/+cw0GD+bglcQ94iq5ulaW/7j5pbWisUiSLFLL
6BjI7Mm5Swc0cmM/Sob+5VUbcpRagmaq7dEQ32ksdbopDEbf2LhWcBs3rIT0voxT6CrVMlxoWt7H
KGncEFDHSYyu/BEa1w/8XCwlvZzk+N8OoDfZDHYofcxTEAnxGe25BFwc8Bzpe0o2XyvaThCz2yRC
yUgIBmnBhPlH2mSu1aT6xs3L/sFT0eq//mXXqSRMxKIHItWB/t3+JcdaWXhFxCXsBlAcFI4zdd8q
O5efYfj/KXgKKk5Zc79zeG2TsGrMwM+P9ds/DGinBT7GxNxruO1ebwb0R6xw7v0JaiHUR66QBNUT
Pu4WGfdoMISeUgqzwHmtJWiEZeXoe2LdA+VWmuf1oxhZ0Zu1AjUjdP2HDhEzEV+cqPQJa9bWTvJK
R+CxSsojGCg6Ss41uEWYrzJav8m7GkZiUHW21J9fvnhefwZAmYvETOPXh/0SfLt8vy+/CAuUWce6
yMtI237Pj6zNm4TOwhqWAWHE+hELQg72qpIufuK3zckrQ87SdOrsvQlsvWqXTZ9IccJjzpIorMZK
Jl1PxpFSd0bdmEIa5daqGDHDK+sbPbslA2ivDxFQtE4/mpOvaslbm2ejfndN3GzvSlTOYYRsERYc
j822HXF5Fd9AS8BCKDS9XKUgziBy9DfUEXe7HsNenDZAQ+EdiNbauWwDSbQlvakmGqHvgBp1v38P
JgHgISXRg4WqG80Sqlt3jLToATaAZXPo0ZkARxubLM4BABIhMqHcY6h4FKemslQwjoHP0YAsiavJ
ule/B1xNbYTeH23rdbmzv0u2PepSnXjb5PAX4LXaw+vPrFXzEBNutnRsmjVbGfcvzGgwX3c4IjXT
BVHX5zruhiSo1NNeV98S9j8CkEFBxjTixSLlXl/JL09DgT+fRc5nVltc4NtE5pgth8a+x4jJ3p84
Sqxqst4RcNEFvuQFxBYJJtSUeRIXyqZLAM95cRjiEvvuXrbSBU5L+wH6rWPYAYwqGRgHne4OrG4Z
xapzc6jXSOjEl7tIGsJ77gcomAOJWw45zO44maYzZYlVc/WehBKFYJX58fjrSJicvyoucuOO33Wj
2BJImq63Ft70b9tuKTPK1z0F0BzINr2S8o1v3p3AvLSjnn0BCv12oVv/W083bL4ozHMVM/Husj9s
PNHUZNXvQazsUmhd+ib445RQqgeiDYuj9evuLbamWsFEmG75d5Dn44x/UI0CE+kMHKgjvuYS/BGo
wx9WwO7aQN6+IQTeQNjBdUEpi5Y6E7lx5ajvk7EbjN2QTayX78v5vrWK/nT4DSgk6ubXQiwU9GzM
PRBE6VUnR00rmSLwTH0eewxM2axVsRGrokObVIsQc3xA3ZFwAmT4ryyhgf1U/w9vfNxcFKrWAMlF
WKyI4WRtjCTqhnhcO8GRF21Te9UCZ9JIlJ10kqj63qx+1GtceHve8mPDwxBkKiZZxRD0Ze9CSmk1
0cIcuz8zWL0LPNd3kNzVq4obBPUydDCYzyCARJw3SUu2uqKeDaebA/acK87C7/hd18FdTmhBFQRp
O9wDZBZs09+SbRu5Zo3C8/yQlMlOeFidZ3IiswdSeXRSgW3W88obFaEkjScXXoCmecCJEFWta2J3
2mJ4AXrasJdsJjlr1FShgNbfibG3I4fkZTlJbNj/t06ApHi960aO8BpDzMUdRt7DW3fJ6LkdQK/y
b+SapN0C/mGwY5Yre9XnkKEUgJq3CS9k2PCtnVCW2hVpuKpHHbuOVtybpR2enCkAilQyyOKvMgAg
8TQUXV3tqGddY7yLTWhlUO4CTVrCvwu4Li4lNSn0A6E8YOiyvNSEHZfwM4kAgHicCWF5hsNNzx3n
Kt6Xaz1IjF7qIbsSzgbS86GAn1Ti4H6kKPpMK+cZ7kb+SpvP0creaH70sntFOUi+ibRGCUCNdZeB
LhrUDPlwRp/1bI4p/Lm49jTgi/H1BFMKml5D1VjfxNiYo8ro7w9HQhDy0SuBXrEFk35DMxvYQTkv
U3AZ/7J78M9FXd9Iv1gjf9mz5swVB7i9iDge/d04FR/U0Bx9pdR/GoBzent/fPUwioX13egZeuma
NKZAuh/fhp2Ecs5JtmGgPPQbE2dFQ65RXBFtZiawwc0lO8i0w2UNENPlE7f58Nu43Pmr8QzmaD+R
s21y9TFjKfZopEmKfh0J2ZCCDecTHHDqaPpuN+5NVaKnR7JcZyh3qnk/8yh64jwPfgoUznEOYpi4
djT1VT4Fno7B4KZZT0F/8RFRFi8PVz2K7KjsbfrbFr+rqzdAUZsUP8roFfOVYvUVBRYkErTih9Mj
xGJOymKk2ZgaPmM0NS2DHuteBc6pD6uwaxqVG/uI6u2UO0BzYgSj/0qo4OnE2VgXqwr3d+iLfNvf
rEkr9MAqcbdA/TIcSB4vLL4s8yNtAlzdYQIG8t/AJ6eV2bZK/jyA/Nt9iVLGR6LN4guo2EO24JVy
YwI9oYkEyfFUnH3MVSElFjBgLAinqlhKTW8OHeOiE4nV+hGybUcSf5OCBS47w0fWV1YIHqvVcwwQ
S6YefRPUN/kxegFYpq70xM1uoCSwXC0Oa7rxMH8nKwcg71/oiDHAd+X61ts1GjFLp1CM6bgP0+lH
eNmZatKO3mocWg7GAc9+qgwqalLcyu2u4fKzkHSZ9ZGnpihoUR+CpdMkAQHASaSMcJQllFvVqxnD
2T/2dt/BaY/lbQS3VeisD4GAevwjNw5SXQz6mQCJwripYSrvytPTQ9h0+GlRZrwUPR/Cf65ec69+
0gx7/NwJdRx2G086DzJOwTNYNHmD+9TU1Jj6ow5JkT3SzhGZ5xWfKEkr8yV6i8OV8XZ1wLBtjzxz
tgB2yT6FjQr3A1b8eUFwjGrsGZQy+Wux/JZizAzJl/fkU7ml+4ZI5AIVMQLvbS7oKpjwAUkyhCnR
wED/3qFOT2q7BIdVydCmhMZZXM3gC8X5cAaYfKmXOzFFbGoxSKQiZtmZoQkSPbIMZluVXTbyCp9Q
KollLNL0R5o1X3vsqkLjjdjxJtf9l2CoHEIbcs1QfhYmtiqhjtWfMxS5kP32Wy9nYqO7hx5dFvef
r8oEfTPZiZb2QHMT+cFZ/iMKHGNpjVPpAUvG7MAVxnPf24yAe7bNYJDdZ2GSkKyl8bLuUzpAxx5o
5MT8+j7XQDZe8NytDYETCRMeRho+6kQLgkuolvf27KIWg5Vfa2KiPVdVRCF0pNFCGuZ6wZ+qbMuG
snMHGU9+EFsmqTMdScEdO9STM6yFi+OS+UjpXjGVBckd7yjuASjovGF1RxAW5U8QahD+krYEcsMT
aoOFALcup7vSHxwF9MAcwS2fnJdHd4/zztu9b0E5N/CpZqCnR/lZCAkgTUe3s7QEfTdlS0Ut0UKT
evjZaDY400nFefVRkceGcUGaqMZYPCauXSE9CcfcKbzV1E2OpkD+jozYI3/5FQAyGzat78AMjaWW
6/4/qXru2NekUcbt8i26f6qCCJILauKc2nG5htP/YHf8mJl4qOs+mtQt6dTVw47HPzoRQhtifFtX
DHyabu0Doe6Y8Svl36kckn6nYw4qERPxpIThQz2rfihWG4+rDBbr+RBVGpik+ifV28L6VaIfmnVs
+UGX0C2RyaAVcokuhQnu1+CnAOf54iPwpKo8DZV/LrdZ9L5xrhI5qElN5lOOe47X+wRhy7eq0gDy
xxUOTtZKiPy9kOPVk8WsLmzzVgsRbC94v3QYHkdvD9w3m1NL+tEZ7H199lMjHMkigooIP2gjlWhL
TqXvggdqI3p6sQTIK2veZ/SAB+FSwGdYsGiSIzzUivtv1prso0RPpiE25shiVYKwi2kJSoVfofIi
5AJtJ3vPytMrM+MgWEtvfgewkFCsyFmOOBCnaEYis4PY1XfX5ifw6RBBhAFMTnWjBPtTr0idjp2D
XUCffWdhThUEC9JrvQ02mXPeOv3Wk3IKdAgDW1TtfI6B2/U0DX0jlzaEDr6a94zylqaBxYQD12bp
vz1UFI3Lrx0Bn9x2w1FQbx8SMit6C6pFy8E62vgJVeprtiVNDEaOP3TEf9MKA3N2cILUytWlR1rK
pagCzX0jjlvFoX53LxV/dYNs6SOzfsq5xKXDX8wB2RqxeV4mMMJcj23UpmUFM+28LKz9MFKTh8n+
3gfoJYiSg6IB4CHuhsyCz5zip/gwhXrYKsVz2lfBX2MS+MlxXLC+tWKDMWy6vtIbbWAl8SMmB4cX
IVwZrvLgW8BKZfSrU2od1NoB8BfkuBPM+Niz5ln7Rf1rDSb3x5f+UBU1m26H5fwj6IQPZ+z//fYX
No0biG8Okds13PMtrG5XqTUdsVyzoBiNfPjWUSK6NDTwHh/anN4RsCFxBEuh/ReCUphC7unFcxug
AphvpHuvcTs5/koqcGReiZw6IthGXiBrCy+N+QsfEXsrtDQ9pGNDiW/TxjXr9PI22G4J/KaZfDJ1
NDz9o1n/8Wwzh4pty0SoM/K8ozPBCcbn61UaUj/zZ7nNekTVR05HF0KLz3PD2F2nIgq0rOSGtvPW
c3z6nJDOXEriZhhHiK8qX2jESJROOz6rvkPMx7GVGmJzxvXg1lxgYaX9Vi84RYyfjzFR40C9dIwc
R2X2EaJFqAmXcUMEn9WD9FWtgMmXPdFfkPJPglbyAX65Noy3HtbPkyAnz+FfQ59i5eTgWDVJHIJZ
sQzc1uHgBeWBqS8P9HXkVs6yI6gyVhdDmkPjM3Uq9riMb8jQsR+iSIquHMQfg8vaSTKdkCtStc5F
PFgnrH6Nz/WKmDn6aDgaJcxe8xpiyRsNU1x+d19wSIpUvDLKFn5W9MacPCml3Ks5wy1xo/Ga/cNZ
F+fkQ7bA2FbQgfLfzVJRCDCsHbxoN/a5vmDQdjS+pEW032Jenha6IjbE4xdbt+DBq5Xj7sTnbn1D
Jcep+ZSB1dyzRKP5cwL1IM8sLF0643ZStYKQ4FBKEjWdC4iT6W4KoStAPdQkjuykqaDiLYq9++F/
Y8bEreJNTHu1AUkBs8UQ5OZi9VWJy9fDxv3kBX4RD4AOidWx5Z7+lrLY3bWxjbj6z4r0zzUmTsUB
bVKsR9sa9kBPU5giHbke8BclSYzXqXD9zFq1M65F/oghxzBPfBdoL/nLQ6T699WDFiHnfQ1enon6
gmaa+nnhgVCJeKrJ+Jv8tCnNvgm5hEYAe+NbRjTCupHd+LaSL1/xGuOC9WzAwD1tdcGvLWchMW9/
zcOxZzOlFvT0hsSqO2A6g2/YreZ67rSt7J76r1kQ91A1vrsjUpPgmGpnTREXKjioNgtd/uts6l/b
XV99RlKTXmxkA2+CWS30dARS2KWrEH41ViGt1aAN4CH3KpBUxudwKYLY6mGaX6u54oFzKQNhN0lF
JPve0bzINmfZY0t6Zobfl0P4Gb1rzseBpaPUpW1FhhjeFoNKz4eGWYyE6tUeuI/c5d/X40FYXKxE
OVO7LvnfWEKLJnMmrOt5WfUcFlhLg8raqNP0HROr2THiOvuVtzMhj/mC2wi7rVlXpQzaMFhCvOrf
gAgQ89CbYw86GLuonEcf9lCAw5YD6Ds16xzRFFHvQzzmTJJ2MA2lQt23/kOm7KDN8a13HgOKhlXe
G7lnXHhrmb8TZxGQ/5cxhLVzrK6sy1WuSBdkDWb3fmSxo+FFt3uyEHuim0Y6EqacBm3wdXpt4z9G
CwmPcoOCVsy+OYH5kQYVrClgEEb2kFpz7gQHfBmqV83QzL9WjTd3ppr88CTKTDESwby5PmhjVnVx
u01u1rHYGUnAgf9e20pcMj5oqIK6dCFEFQhqxMCxpp30XtFca6J0pR3/M8QfnkBO8jJlIlfaYnTA
Rcl8++VSpYJj+uwU++4gnXbpItASSFg2zkjhOuKClhJdU1QKIlnDE5TJkPKoo2EW7Lw13C/BteXT
9v7DR4oJyAqtYeK5RsNhJA1Yyp9cuzXnOGUiHsPuhwUHkUwdTPXocyCDOGKyb80rJTv4F1HfpwrX
uXwYSFQzJTrEjXRtc/iS8rhR2iyw7VH+RJh7tflEZNwzyPYVT0Dt3P3pQJu7qiwQM0MJMrzUhQPz
E/GQLpDwPOwRQQS5wf5S4VvniYFTu+rel+34C7b42ILSr+e1fK+tai1T/Ay+ljgOmlaE9fJ5s9aB
Vfp9AnU1Aip+jjUWsrlkA66YVWEsvDaZSaoBDUwzFfjWxpxCvKQMtCPax9Br74QTKK9xAnLo77zM
tJmS65zR9LnyEYq6L/PI/9f2irUOxL1gUjBIrFk=
`protect end_protected
