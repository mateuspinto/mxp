`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2160)
`protect data_block
22PfpvHNoQqNYioVrmUVzSKAGjZUxFcffNRw/HdXolHZkTDe4RION6ba+SvTtj4Yr6+5AM4i777w
43vqHxsvumRXrvO7lMILHHQ0CUcXaqnEZmrD4W0RoGt6bFR1b6jVRh4UjM5qek9eIQmm5O9/jhev
AlSwTlS7gF6piePI7B88YJwtN6VxBiw7rptUtw2xZC3QfoYTVd8xwnCWRWml+8vtuc/prH2+2VhH
Mn99kzAjZriS7oZRSZZ3/5bnsIkNLAolWSXm1cc/VkULSNVqOlnkMihRfHzY84cEidfnngMkh84z
uL5e5OeiOXWOxE1GaTR5aBPFjY7GXYSs00ueAuz250quY5Hrg4iQHivO8y0bQNcqYA+Xont43yhB
HNztFJkuN83zU1+W3Qgigg5VKqfp8RUBJeHV0MkRq26bLLFMPNz0fofWkOpianaHLWh+QO8wnyzc
ekVPnE9ybdY3Vf3bXA7ydnwTJnSMNWzjWoVtqF2BSvYu7ADkMtAb1puz6lWIGdr9rXFT3j86aRD/
rNv+S+8RpaDX8liTjUD2r2lnmcr06uqxb4vtmOufP+N+Gj9uMKBGgSRysMZY/I2BJT+w0mxErO/Z
pt5FTOp3mM9KHmoK3B03BnNK6Ru75FkUzT1amX/nQtbYcvzYbvl+DEB0NvuPHtqp/F+8q6UT0lIb
1nbOR0q8E58M7juVbBkpSZMIByMgfStjV8MviXDjDAfxS7hPCtcOnkG7XWZ1DrGYgLiK+YVkrJPm
pfsS0TQxAp/jbm1jCrEca9nXLmZXTop+qXe3qY+XVQVTIHm/Xx61IoWq8CQLju7wmI8Cc26Mkwqo
0v16OCuO040pZK4uYdEOHO3oeXGLVYnRWNTdDnGeVkrBu5k7LXxpoVnO9Eu0wSp0Iq9Aao85hgeg
FIfUYnw8XNcJUvIA9Hf06QkRdSRklvkihbqoyzBz3IIh0egXAkFJHvCmrO9bLIXiefwXMQWXXXl2
C4DzVRH1gvNE9J3jEQAUXgbyJ1QhXlQeFdpxx/bAw3N11Klgk0obYHOSWMohB//Z6PacqoPrRgeQ
8wgJ/fIK6X29EzirU27LB5b0Qjayu8qWuA6u8LbGYnMV730bCgv16Oz8fh6jG7cagw0gbuhLeoKY
MXICs3BCj0XK/JL6mag3qjnBKuHr7nkHVfEcR64y7TxfVNZfNaI9JVOH0/dx6iP9RP43/or8MjCE
dVI2cMOCJX3fsGgfuKVYriha2l6XXHPcCV/ToRZt5OvqSt9r5/cRE4Ln/sehFPYTwEvGcbB+qtTS
VbsIr3pDBcjY9M/yBUQPFsbWDLCUENlhr8wzEXkPKSf978hoSOCFeLWdYDEk9NV5Vm7hbSHtjYft
k+VwG4n1HWx7SsVqCzF6BbAyn02g4620laxAz56GIw0l0JaqXEWLyx3X9Th7hbuH4eg2yICe4Eq4
a4BmPi1VMhaySO6ptTeGnZ7ixCxyleYlVxRxZX9uopQU1Jc6rNR3yGyf9FJbq2WVl4Y6k86aQMIR
VSgX/0ktRRQ0TuGzxuWRrlq/NR5TAy/VWC2cZE5q30LYW8qI7owfNIztni2bQuGxzm86uLilHVql
PsxXbbE3qDkNc4LbiWQc5U9aJzifuAc8jwt24Vc7dFa7sVjkXN09W1d0Q9igmVTK3qddtTszbuZN
0NY8j6ctZlUt3yh6Sui4S/r4/CrEcpxMHbxtIucwjlJ+80zjdVYcoksAcNLqSiVBA02AXB5PTB1n
e9pzshcAz1dXr3UL3gcBBAtQCbvTPCI47xeMnRQ6+mYTMLmbTZRdBOMc/0aEaLPdaZ8rtC7i1x4l
teM4XmPS/QZXROZkm+8C+IGQnpYXbPNeVzlsH81KRVxUnhnIqvJ1N65bxqkxgRzkxxGBnxB+70mZ
3HPDVUUdWiQqUQc85yt5QlSrWffrXVpLWIMpv3h7RvaS0v/mmdo5TydnKlpggEfdNUbQBGDHwbsZ
LiVJy7+zJdf3XQzLd2R6srtDQVQT6FqdaTO/LBlgXn4zrPsmX+K9Sf8nHcHCCwa/pF8rW6LVyuMI
NXwBoPdQQMCQZCy9gROSBtbm22vb+cyDvoFYk5PyR8MuHF1byFB9Nwdk/z5Okc3KsOLc/a0/b3/p
imsLvVrbPd6N4ohn8y+rb03EledRGVO3yvcHTHJcnXC+9b7yrHx8Kfd+Zc9ayK2nTOG9PYV8PEXe
0aeyb2ike1wMyZpVZxUwvQr4XUs3EZhCPPwrVP3aPZ/Bstsida6SMjcJCk4Oe1RrFPlh90lGi/oE
lCeOHPrlqeDQm8R+vJvCWZkIWTSImQcRX3gfoGfA0kEOYKJPrv8C1iOgQrvoNdyq3dxZPH5vKzI6
psR1/ZT0dOCtMG5bUClwCkOawQN3WNr0ZTL07psZSsVuCrLr8PDxxHaWJYV2kvwo72dCLFhwm4Dg
vEkHmY4gQf5pwN6HdN0UL18Gk+tzqhJhOcmED5sGBAuhlc+8iWLKZkggtGn2uZRP7a0NAo8TC3Qi
aL4atlWDoXwnLPxHomotPR3B4EIIs0AWj5TXX4e2DfjkBukPaMqKTJ9wXZNtFDk5AcJM8FlzOAdN
GxNh2DOQq8o6UUnGyoy/vTGseIOywYfpSA2MdqzZ++fVQpJUQel6tUAzsYaACehve+Ku97ETQUdv
cdj2OMZhk/U8m8L9zDmDC1ebQH+Gzo5jLkvDGDM3JIJzghOGa7X/kJXbCFJxVuKX1T4Jl7rsvIaT
sgmKbAMGGSDBE0tIoqNDXvwI47KqqBIJIjgcsUBec6U6ORqdH0lc2IIrBdAv+wbveg+j+3PO5TPU
Nau8gjQTDSN+uRxoT9ZFMH65ftdBlma2ooloFqYnV41y0rAF6pyQ94IaYnVqygbzCBuI
`protect end_protected
