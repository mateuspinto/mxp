`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`protect data_block
B8dDmn2TZZcs/o3ORMJyj6l3Sq6JSCPwYTb5psaGmZxF3paw0riEJo+IU1S2E7QERiTSlhMZXGGZ
nSoMRokdi94cysRnSKPfaR1c7q1rMVHbzXaBtZbH56pFd8fMgv0Cv5soywTeCFyHF8sLP2niSfGb
TEKypKoGeLkkJkhaqsyG8aVqNUK5Hb0SC/+61ULlEvGDoClVz0C5QDeFTaO0jie9F0rZCJETVGzj
k4cuKpc+7WaCywmzyXMGphWk9PRJ6mQgYyqXpcp2hKrKVPYaylv/bx7vBpG5Hvas5h1tzvkLIxq5
4HtrRRaJLkkCv/q5pMAbAMdwOgo/TqB4j8DZ9NzpIeMLm5SJaSCnDfNHQnG7Yn0ZiFXJwg07f58j
3KrnbID4vc19yzCseaoHgzy9Wv5vQxWQqu9UBeauoSBXbHUT3ozrW4NXtoxkwO2CsXoNMkMEQhPd
9sHioZ8zF/bUUeKqLAb6QsUetLqbCSqh6HapUbCOnaZSznC7Iim8o/tgMFiB/FEBXPDJh5O90a6o
IEdh5eyTgvmY5z2VK6VLhfhhq+5atcBCGo49Nbcv8UQ+wx4Hsd3F4Tzm+NbxenFQid0Zz5w/owtD
CVMXeOfpy+yvTj4GdkDY5xAcHWfew6zZSH1MYbpIL/TWQ6TUMZBa/6zvsffLnN0S8Kgrha0U1nah
S32o6D+P7f5eHcXIpyvKSXSKcQy/vYYlS8c0IJqny7tWuXxp96QuZGxMYttf1lSIW8xCS3IyBCEA
gQxK5jebzOguVoyWQMmSR7O2c26MYUp8+fS08k5Iw0jBo4a1iv1acCGou8cbr760dZFqNM1GVqX2
1uj+UUn0/EWF8baco6FAi9ZPPAWfx7fCACTuRJFVa3F4rlNRWNvteVhYy/585GufA0xCBx5NOwid
RSjXSt68zXmGwYbOGj47/ApdZC5xqbyu3jmr5H7RRvO4CAYC6b2ANnTqqOYGEBOyOOZAg4QAZd8E
uaBTu6Kgl9WzDicqAvyU5NmvxeK4/aunTFbOzjmsOXSCRDmTl3l5yEfVePvLmSCahBXI6OGlCt/O
aAkYDMXVjo+4+LKx3xEg4C2DtqVnve9TAzVSrVuUe+sLeXGsL9E8H0j7STN0G3w3I7WEuEazmpMH
V20qys/ar+4vgyLCs0/bwM9wQNjZtExGCNFubnKu99gyCblEFhi66ArUXXAyAQROBHm/Nvz9KyC0
R2ohMnbUSaISjnSzobH3jjFf1eX+zLGooAUX+SqhqxBNSmVr1cAhfL//KOgIuMtDA9UxZe2tm6Bd
Zd2pBtBj4tC9LclFPsMt8Mlh4d9n3f1mIwm3SdiyYmH/JGb02fYEbbJMpfOhtDYq40TbUa320kRS
xHs5f4M7RiXOnTKqosFZ3eqKH3kWAZcFOSVR5i9LbKDG4TqMz/6MC/O3HOmUD3hDj24mdQGdN98B
93T08iEJU61hU/zWnLTEtMYsPsJQ4fASztPtTDQT7GIv5Nvmui4dL4wmqMlACYZuJeLeSvxNAF77
9DM3FjI04tfkoVkqm6TB17zI8YvhILiTQGouKalhhtJMYisF6MbogSOhCIpEkvh0JmGxN73voP++
YoRL79coh7DDSY5trJ0f2nsmTSVnIJu2PH3+rASC/zEwc/ACuKQnsCZjIdmd9HPMRzmEkPgo2kLN
bTNCXbKw28YImcS1uW+wUs2c7Fr7Yu6LzNdnS/YtYt145czAU6AZb7HcsxmyX8qOs1c6oOMuqOm1
WMEtPFdZnJtw8kkI/ZNgZei8zmRk99p6KVTMGz4D78G05ED1fBnuXMm7DwrjU68Tb3sYHlblGHws
G76hbGVljHHT9ntj9cjdyfavyZSF+DJYIj5xEpWfeJ4SQFbg824SZkPVNJmzX3T1W1ODWTmj88Rd
X7jd5Rdk/cbaxQ2pnc4YALB780XYjNMIRP6dJpNUWwIy2o58GaFqOHrdfoePN8ipH568aciWHOel
dX0M1KlnEo+qTaOK1qMKwWeBvprwZywp5kpCWtevu16hO6x8e6QLXCmvhOwrVyaXp0Rjdhfy2bRx
ishzTHNBDP7vrCaodJfip8/ZsVSwdMwGz+jttP569HaSxdkFv/fYFDmq3V4b4iLIRwa94zKLRK6d
ZIKen8+SVBx0Hxd+P6mVAU0fe6Hq1jurOUHgLJZvJjXO4938CcNys9S9pdaedu8N/8/nf05K6EKe
FdAJOQeBTNa9cz9tZPJnoF6UJaR2FQ/9MrgoIO62/FBhNTQ/nc2eYLDbQT5mraSitGfP1INhL5Je
ibH39Ruxl9AjAjqWf7O+Zh6bb1rDhdPIKJuJEbw0j70l7fKQedh6vIBc8JlztYOL2otfS+/3zp8e
tvSp97SUOBlO/8YbVorZrsCnYN0ULklB92PY0/cy0zwD1bMzRhWXNfWd299wWko8GlSEGp8YoB4H
uHssXW9EVlqUgOCDdLWUk9tJ+svvPNoHSDovWlIANZaAt/nqmuaJJWfuHtzSSP6h1wSgCZuLeiwT
UyDIocUI68pljiYSczEvD2Ena5i7C1l/JYwsPucFbl3059dwkEkqcdOzxe5o24tqZyaTSdWynf+A
iLJGZULMJP+rnriUUL0RsNeYY/XwxtrlCGj1qEQEiXSf0IYWPTMBBzoNmFA95uUsrcsiW7GZtzzZ
bHK+SiIzE1SJ/Sq1oDcrQmzfcAiMi19xWSNxg/ibRZRAlLGSl6XosntaD3YtzuZO7zdYRDT1v2+n
9sI5I5B1d3pC2Bhl+E3ibr2TxaVrMO1muV4C4Yv6dzZ/QWZB6jE+UAEAXrreLkjr+IMkllPDnGl4
RD52VZZlhkhkQTXRaPsM2KpNRNzMb7U6ujNkPgT9eH8UTEvEohgZZMNPbz32WPx7Hrcx8svZysRr
GN08vof5ZiPKkR4cD3pGrrrsDYT8YW1UZh6uF88UgaR/Tel2peNYKg7x70NGeY+hBZGdTA3+/PIa
swtaujdPftWA2BNf/v9hXLxM+tZqzWSgpH5tToxpp1KuU21ca5ubqCRqbmG2A3W+SUiXuPHCNpA5
tWtI22KxXGRQLpmQ9AGSyX5cXqg1mPtwxZ6maTLHnKrcVMJ5heG8TUYSbRqmdEUyaiTFqzYaNqdU
z+0xSffm5XMZumgS3gk6kZi+O77ajIcugopLsDmPtDwWcyFCzoxDqwKgYFWbqku4udOmPQvAR5U7
MYzZ/6jyGLdG/1MmBSzV9/xRFoBAmoNreHQpeG4NT4q4cDR2SLBOHgIPDCrITteJGSc4jhjtz0rc
pRPYxtmHC2efMe03wmKVgsOll+pwKQ6Wx/oiyb8ndKLdl9NbCtXVhaMO1K11y30VvRTINtu33H6f
aEyZYGI0y9IXtiiIsqvZoJDfU7j1qzkkU6/Rpl2A7Vg2yhMQNMmYfmkXyZ5mLV75kjGcyLil+5wp
9rA5pG9AMBVFFZDZbBwaqtXYKvp5szthpINJ6Gc0hMEr81n+fn3EAHwV8nY9tq7K1NQFvmAivUbJ
vBXsEFz/sbGuHqnTFcnpOdpeZn88oi6mMY2e9c8AFlZ+NLbShWCnUlx5Fa4oUKD8grOfsb8mug+c
bBSfbX0PpPuc4Uujqj4ysT1iZviOrb1FnGt6lz0WILBbZycf72eVcXuPiHwUspOMegayazjwXsDu
AbfnVm0W4KKy/Tx6Od9xs4r8U9hRWmsSCiDQaaDI4AGbteeED1dp2uQZtuGE0OG3klyNpZiPIoy5
WIVyY6+qiO7akOvGlxCT/iwl4PzcYgGzVLNrA9kEVQw8X2g0Ll9IQnWJDskLRjKtHAXK2Q9pNWuk
vIyRXqRDJS7Q44n3CSmrscvqgXD3zQcBQCGhKENfdu0727QBMBM70gDs9xyBMXGmPBq5KK9MN5d7
PXG4p0NHiB9Q45ehMSY2T1VhD60hpKgCeXF/8BTUCTrzlfpXMz6lTeMWQ1HIjzXjC74V4rRew6Fr
SFRa5foFGEAPZai9YZuULQoDud5+0gZs2YnRntH5ZPvM2Kix7nwQ9pFqadJa/jBjQWd42sXAbtLh
yUekIHmT8xu80I8kb2whPK3FYLROqWVqBlGoAI+S39kCPns6PWbj0Flnt1/Rj4qr6S65dzIYZp9C
qXCiEfSqdhCgdq6nzOsoNi7T1uEaTFGxKy7VBYO+xhzGpRgBkjBCpZhF6nyvFxRNS2Hof2cp87OM
LI9w+sD9c9RvODkT1NN4mSXulhNBR9uGvAGuq8hqecVBqyGgVSjuOWbi87VJEmFh0ZgTIHAYbdaY
QVgFW1tssA0BSB8HnHLYHfW6FkSDaSqL83O2Fix8YDohknWYwF63nZ3mseQkb5eqP0wmw7adHGNY
4DPS58ejq7flQMl1D38ZH+wAZ0E5Kmdp3kgEJASpDrDDdm9vJ71cfpnA4GizeyhwBkydwnbtuli5
iDfAOhPE0kQ2D7fw4fWrPg+s2aoc71O4e9dqkbNwJWKj1fiUuZrcqm22DShQS8Xx3fDNNgTxPFJU
2PKfrD5Eb63f1LEtAzq8WlPBcaMniyY+upORKNPpdNaNx9XXa+NpC97vkIb5XQRxqz4yUsxcrNQr
thCu8qT/nBiTVhQHpd4n5TQWIthLh39Zy5/cU7nLVld8lTF59Xe2W+Bj5bTMTWUSDxUeZ7jOfpQ0
JNUsirzS/ZdO/3k4rT1o6TLykWO/DrhhyPZH
`protect end_protected
