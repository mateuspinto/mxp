��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���=�:~�R�Ÿܱ�*�_3���Mb`�5�tp�������K7!�S����B�Co�dT��z�s���2f2��s�m���_ޚd�y�	oQ&@���7�y&= l�y܆l���9���U��"���\�I ylyg|]��6���8]��-�B��<-�9�b��C����]�e�l�/W�ㆩhK�d��3Y�7��R_�#��#B��~�temM�8�����'�C³�v�����{pX>�E�mh���+�q>��]\ ���҈��g��Uf���3J�i��6g����m��3�]i��l���Y��)��3
i3�S�Lg�oy�@���#�yid���W0 &Q�D[�iX��e���;X���?M����\gnW�4�l�AЀ��B�_Є�9O29nY���/�p��M�1G*ye֤���k0>��J����6������鵥e�G���m�?OIh5tQѹzl�wãf0��B��1k$�`S���K�6D��;���2�)��B[[$ov�Q�,L�j�:.R��p�Jf����-�B�k��q]��Mf##�c�]*Ptផ|�����|��p���X�܀-c��X��v�cQ���o�p�`�m҂�es���千��E$�f����]\O�N8^YD���>���{�h`�Շ�CaXp��g$��Uqxq3�<�Ǥ̧�]���K��l\&0.|��D-n�&�O-�H���i�*j]��	%�C4>�T�ڦ��+�둻�5�^ZN�t+F�*�x�HL^C�K�.eEC �y�F�𑽬i�B��-�[E`3E �@�l�c���J��Z�Bک�%�^�sSq?�b�O�>(-�lf�&~������?�N�>^�{���"���5�j�O���o-�y5C�6��xu�7�;a;�;HYإ�B�
���`����qF�n�6,�,ժ$z����A�&<�����˞ ��~�3t
��[�2C6P��e2FTAu�gf�ѡ�B�$/��)�%�S��ߖ��7)���u���ܢ&\?�����!�y����u����d�x�`��6OSV#+�O� �h������sP�â֗c��:x1�T�
���\L\|��G����ɆJw'���U�'�[C�֊Ք�#7{I��q�<��P3�O�lҷY.,���[P
�B$n鄶N�2�]��<�����\�Α~��&����Ĕ�tڻT���<l��%#����ACk}�]��7"���ӷ�à�f��P����}�<� �,�5>�>l;*���c;�vʳ��q���
��Vр(9�x}����AA8���\�*X�F�;B䰑-�"��ۊh���+�m�8Z���)^C���,��	��A�QU��A%E����fli���+g�f�m�����p��}�P��N�C�t��_��W6��he��W��ɕ!���~ Պ`V�x��V�]��1`"V�&//����7.�;EF�4�c���V)��!�����T)�����ߗg�����ea��d�F-�2/�+n�d�c)oN�'1���,@�IZ�����D�fE�0A�NN�cc���I��n�8����7���"��cSl����a�|-�o ���q�͑��Xf���|��Q�+c<�H�օz���M9U�N��}Z���.��>�tD'�=Dw}dX5{��	�22[�>[И�U�~2�<o�
��\4���y̒�c£�%Z��Q��sD|}�F���VF�]�2(�h�x��i��^m������f}��@!��_�c4���%���
�gy�g�!��S�TQI�b����� y�S�:#7�}i*z-���g���O�~�(��:簧E�2t.q�ѓʔ�e�K��k���H�&:|� �k;���Ugt/���e7��S{��j�7���(��������B���72{�ʧp��Q�W���8�u�# +{l��A�e�AW���v�W]����������ge2Ծ1S������6�?�#�$�h�j�J�G�?�m���c�Kn LL�,�[� ]��ˊ�Nd+8��DM�Qw%�ǖU�_^mm;����9VoY{���/�1ϩ>T�yO�(d�����}�E�b��.��~[�?�APF���p���$���X�1W�/���Ss ?����j��7��6rE�z�43��7��Έ1X�).��19:l�jD8���j
F�|5��Gt�;Ƅ=(@���>�(���9C�2��T���T�*��4�_Pvf�nJ	�q�f!���{sAbN�(���5�ˁ�*��T�I/.��U͠���	�s����%t���P�4�m���@	ZD�R�>_�][�#���BX5R��:��U�%hy`�C+Ǔ�}�%5hγT�\l|�x`ƿQ|���^ B��=�d�vܱ����e�������Z�bOA/����1}n�#.7�����h�-@����f�I���).���o��%�]��3�-�B鴬��f��z��˔�7q�!���/��E%Q��W�5�k�+wg���UA�_���-����3���d�[���_I<{��Y;V�v��:�Ƃ�{�������-�o����=~Q�= �l�oCk�I��l?�����@��꺝X�b h��Et�,ͣ�"�xg�o��t"��}��H�<c%�XM�{�Rì\�����ٙ8oW���Ax&�Sbn�>|̗A�ͤiM<�L��J~�G��r^�E�#'�a*����A[eZ]}2K4C�[�+��wK��}��v��i��7��N8`�U�
:/H$�vr����c�c#r ���0���QKp�i/=��@��K��ܗ/���0gLL���3y��x��;�vo3Vl�de�&��������AB�k�Jwb���9��E�$z]Y*��?��GAL-���ANz���7�t����KQP�eڜgD�����(��J��%Փ�[����t��m�Ǚ��	��5�)�o�Ƽ����x��6PA�����(�?Ë�,�U镪12F�[Hz��� o�|�(n��<�M�U���*�\�84��EA�2�q���(N_���n�u/'�j��f���+/Yr���c�͞>k(��Z�;����گ���HOш}����p^�<�K��O��lܲOy �Mh�v&%�_ym��gϔ"u�K�`g�5�� ���mV�i��q܅Ex�B!�)r#��1Mо�D>x�L�<��2�m.�m�X#�Gi�"Ů��{�ҕ�_��W�z�h�XZ�'�t��s�?���}�����_^s$�kӼכ�"�d���\��
S��@�`��y+a���Sz�l?e��f����9
�� ��Ȥ�Cё�k�����]"J8��H�������sǜ�F��ӏ��2>���`$�;昧f���I�Aҽ�A+� Z{6�����
��������tRA��`�Gw3��������<h�M�I1ض]5sB�)v���NO٧"��5r�� !0��gt��ǹ����-��i?�~��5*�� �r��Px `eP��l2���<����y�\c�VS:m����9��ׄ�!����T��6^objcR��M	5v4Ţ�A�^0��0��� ^誃o)� DDq �[ R��h�� �}� !�WE>Xef);&}��l&�˝�bQO��\1�]�V�B>��D�F=�����^k|B�:�� ����������p0`��<���B7�aX��s�O��x4�w&ޅ6��Ml��D�dln�{�7���b��}4(����Zd�]i����� 8����|XY�����1�'x}�l�p<�P@�l�y�.Y����x�s�OM>�N!L�����q��r2E�_?�ї����SП$��h�����t��._ ���O~Ӝ=���{_��֗�mumWP�ʦ��9BW~.�hİ��\]��sM�lV'=L��R��B-v[MXq�/��x�8\N7���.�1Q� -&}�{j4��iL}���[��e�7V	��S�I����?�h��v`4L�����j�����^	�lC!�B �e�j�|%����L�ha��8�1��������c�u��Y��gtz6��*�!h��A�x�R��?�v*�桑8Yu��.���>=��5V*�_m���Xb��ħ��O=wH�8ŀ�������Qe}�!Y=�2��L��r�t�w����M�Ȍdh����ȟ)Y�$�a 1��o����R���6���UN��:
`���ӯPPٕ���ԑ�"��i�Z�e�n'Fl�seT�$>��~� F}):B���eUs�#��H�?7U�\� W<yM�֞���KA/�JU�cV���ƍ�)q��*a��Z����-����Ka"�T��n-u��/�ѥ�6�@+�F]8�5�q���` �.3���j4��0k�W=� ��\~r7f�"a;;JZ)��H>��T�47 ��p|�()��12B*�Ǿ5Ď��*)`r�D��[������Nz�OU�%=�	��]ieH�����Y���e�3?��rA��d���y�9"\6T{�HC
�on�Y%� A�Ɲ;7j�|�4��^M#�V��,ɔ�K"��C��U|6��Jh�`4�1P����`d�����N�3�hs��Kn	����rG1c4f��6.Z�5A���ׂJ�Dm�.���%e9_RmH�eV;Y|�Y��1�����a}�D�ɰ)u
T�k�Jbpޏ�����F��"�k|H(��cƫ:��3'�W�ȭh��U�S������z�������*�3oJ�J\� ŧPX���S9 p��q�0��^�_���=��-�$f����ՎaMt�|��^է.Y��;Ȃ�WGh��d�������o�a�p�cf��S�U�� �7�R�S�Ma[�ۗ����п�NlhZn�=�%�!�Swx�ꪼ��J�xSlSO;��(:w@"��V �A�
��I��yҞ��d�e������_c��<}���"B��ZA����;bC�{DׁN<h���`K�"��H�>��Gl��l���zb"9��i��1�:1C[�����9�eI?�m����^��*�I��$���"�{ML��/ݛ�I\Y��0IlAo�����YV�`g�fpP��{�d��ޒ��`W���yk<��ǘ���Q�|aC��˴�������M�CR�k��ġw��ߩ��hyp�0[F�����l�=q��z����T���o'�ͧ������X��P�
�R>&32=�0,{D�8o�r�WWС�fɠ� pe�K�-�+L?�Z��S{_�>#���%=�0b���=��΢2���^�(�%�F�G��i_F.�756s��(�����fz�Dŧ���}�4��&�t��-�)�%wV�y�:/���޹A��jw0KFZ�4m*�/2�Zfs����a)��m��{$��S���^���r*��@�%қth����Ow�A5h�%�7ԑb��d�zjQ�8�k\���Pױ�g%��-}�A�+�M�}�v�"@Z;{���q3����t�A9џ�$(��!X6���~.o��>1f�M8��9$�a� /�'��/��g�7L�́�BY��jV8K�쌩`�����q�1Z�Q�b�1^?Ƴ�ñQɶ�8�	'׼�M^�Ȃ��롡�\�@'!d�^����I6�#�����`��.����ԃ���Cy^�=��������ܡ$��9Qq��R�*Y��V�5u�o�C�Hp nm��E-�������s�H:�]�.r�`�\[G���
�;��V@�j����k��Q6ܽ�U,/c�v��} � � ���te{6W��kg�M�:cX��p�I��a�fa�����Jg(����<��-)ʚg�c2U������݌���/���fRwB�ku�bWx�������XU	������8 ��g��2�G���!�������b��|׉�?h��l��Qs�X��=����h��_��fO����]B�~0��X�� �^��Zރ %!%��N�ڻ\Ma�mf�H���Vq������J�*��������	y㚚���Pby=�E�)V��t�t������W�I�3)�9�iJ��w
vak����Yy����Q�J�*��XpN�t,~��]դt�,ړ9�)W=ln(�%r��@��5�>%��~�ŭ��oiK1'���5A&jݸ4�������:D�:�����VC�(���)�%ǰLF�	qe��uGx���_O��C6���>1̚Gʰjt�C�