`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
J+YltaX0SneqGBvZQvk60SNZ/agkGIOyL6izVRdSoERsXFLGGVWMzVGMePHx8bnO72XBxx4TRg3G
pXpqle8yuJuBmM6H3GLS8dJnPRvxqhGPTEhays2Yo1Nc4u2Hna9FFhgtT+pAftU6/Swcke3s1DqU
XSbcXsgpxeJMuT4ZGp5bYqZ+lHXsWnKfQxRtivNWQzt5qLmP25b4D3amDBlIBIIIxkymmXDqqykb
+M6TGI4PAXcwBNE/8wrBK2PkZu/wP/AEWsHjkxpXUSzfO0T5w10TBEjzviwhe4O7+B2wcBOzOgyU
S02BxRzoB97qct4yfUXSNfvC0Dhmt0SfY7vBpQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="wFba5QM6W2enYMsaxFSOFaQtQfR7GApN/d7cV+BQTZs="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1120)
`protect data_block
OUB/Mn8j2La0PkLgtMj8/FmKcVpqplAYRjRl2FhXqv4uVDlpuaRWPoJSLm4ijWFNmA0IS7IqErA1
pl1x4lALMQrliJ0ARg3DIaSkHh0ZyfdKcJo0+nap3KQ3LmJMA1hybrvGSDQlZg+avfi1vKbx5WqS
Y+dwmoA9TeKilqsyZcXYDsW/Qz1gGThovBgL03k9wN++qxovR8u6H3TERTXQsH3lTWyav25xe6TY
B7iFySOYsZoRMUSV/3f4DOBihALYBrSZMDUqOSAKPXtTxw1BCFMr2yextQAZ2FJOntkpUpFx5Iyv
GX4G3mJHIHoLyl12sVgEt6hjqOBKyhppLAYlYh9H4lvC4LQd5WqIHWETmpqmUlqEsMlP+gZgbT0E
iL1G/mnHFk/RWgr37/z4y5gKI5qnBy9JI8t3EWGfYkGt650yGG3VKxSNdeSN8X1VcVsIBFjvye7J
1l6frKc1TZRnKn5b3fjGGX0qAPOdO5m/yYgXaGqo1FOxe6WiR3Rfqfk2FmFxQggPUgvzvPsQ2Vay
k/8HxiASghr/w+796QUiDdOHFk2j97bXHf80iDWQfn4LwpGsdyWzYMPkPBQh9tMocC8ODcx1LMFR
TjksG/+Se7Wy9YhIZjrwIDfD6d1QFs/61fhnCiCNBjV2vRgZbHxXYFgjvTLTu+zw2AOgMFpCRL7J
sgTwVjoe9KPOWAK2u+K+6QERGzHxOA4OC8LlzmDzkAv4StWYxxvmqTUj/TIgJ55drqKk883EftHV
OoRQ0cjXYWBQQm1l3kONA39taw2TqAuw//SVW2xstSj/KMvlTnnkz5WFBvkfzuwVU1qt10/tqecu
F3c126nirN9CxlxLBMd3VTWSfjqj8p3+EMHNdd3+MMdHxzKVXNmCf/LocECr9JOoug5Z7PmodVDS
Y0/5JHDcDetT+wpU0MDQxnWMHvXhlGGR780noHWDgF+F/rbMM7Fvri6Ma+R2LDRQHfQvfGldUKk2
trNI5yj9OkjDyRUm90nEVCsoor90JTGh0cpjzjyBaWWSj+Jt2SBka1rrW5f1GBhU2ZXRYuIT7JNb
Y2AQnSUeP4U+r36vaHZRNe8ZS4LvzrXFfBG6Et+DzGXduehIHU2nKmoZqv1iYg/Zyij6voJpZmhI
D0JYZtt+j42kQ4jb/vPhmzqjqHZ65FOko24euezcFjWJB75RwPq5VEV9YlIn3kyt3r4hL50VQGBs
N4H4evVjV3wO8hMMKvEW3GqYktsZKQYuqVUVv0W3+cdcZ7nxOHAuKBqPb2LTZmArlc3qDX/gba8N
/SGUVn2AuTgilH/hYWyXPLNCuzeklbxn8Wtf5aoyFb7eg/rKe01xzq2xn5xEuL9kDOC1o+jpEM1V
y3pM2m4CKpef5zQxn2N0yUn2/RfJnKk1m9s3Il8VfeFeDEPwLT8eixmjqKF3G0PdNcsiWDXQHKx9
sPKMgxVVH4H3RSsT94J/4t0xZEtd9x+2KOfd9Un38tBcKxDQ0w==
`protect end_protected
