`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45824)
`protect data_block
wj661hPIflZG9wLbVJc+d88fXI0UNbRVQzCPbe2ugSwW92r9buW6oxbSP3x8hl532q+6ri7FjaNL
O1tJrmDmtsFmCnTKX7dpTqXN5ADmRQKdKFUDobZYhAOHHngljU3MSAo+Ra1QI6Jteiid7LVgDZp0
vUtC6GqDJ/nlzn0u6kfchx+MxiwltUZhjZkOOM7jJ7efojed9VT4Mcz8qRU8Om849oYFEaGPThoe
gH/TYMCNy0iOQHXLhn6C4gBsKZkOdjV+9zkTzfVGw3irw1BuqX8aiNkyJLvRRFB4xAFtprEl3P5o
mdI+L0hhWqE9zxydgWZOJZCXj7BS+2xlBxBgFimR3sVQ3FHviVO59IDcaItakuMVdiUbsR/oIXEc
zlJlfG630iFrldYNBVYkvEwvxCVmwv7c3+jwbef7n//nbyvYnV69UamAab6d61Im+BpNjRUJzAWv
rObUtDwQF7OPo3Tz6C7HONGw3s8kCgU6YRE0rEBM4RDC3QVyQ1SUs4Pml8pCtObCndBYOIC6/jRE
pwqW5wdLuPUZAmRcU1v+SPPskN62K4JXbMBdVWFepXLkEsBYc42/dSq8htZUkHb4ZqAyTu4EWhHz
/DSx27m8xnqFGAgqWvcL4ofumXzzFIL9UI2PXHuyCp8IFj2xvqRgQQnmoin8q+FSkhN56kyJO9yP
CheZgFleB+Q1rMxs9mDHxKIKS36OaZHlG8zAfOzh6qhFz8hMiTAZY+uTnLyTTFfadVfEKa267WvC
1ZJn9rj9OnKZcxoHuDHCOCbJuopQpWEVbo/VBsENRoXYx1p66f1hPKLXVQVZlr3WX3ueizNhM6Yp
jV73TdyUZoqcXJef7qOKpGsk5eiQoa7sgJr9OsKUR2UpkiaVgtnq3OEAwi4FcNntxqZUD37ai4vz
YpJPOwNejXRB5L4F3ji1xjOTNqTCMB3OTytq/JP/qltUDo+xAssL1ZKJnoPRjpJ9SA4nvTnZn2QM
cAPD/Cf5akwB9pjY3zDq23KUs5hMd6csgKQS42Olk5WVjIUuO4l1t8t8fOzpRy4ay8FFP8YnqThF
D9kqyjVtfx5hlPXX4QnF5nf2T6Dqna58RrMcfqQkoM4Q1CHksiya0BTJV0Etycp/ZXqw8J2tpjmj
yUicazEyrr1kSIaz1ABf/c3ujeDM7oM5NL9zEZEoUQ8FXJnpyezAAT2Y4i65ew80D58sQw9u1vy8
W184ht1wf1CsGUvv4xIL6CE5axZAiXv3dfgOX/THaxttI4+XD74hU8wIqjMZD0LnmHeeCbRJqu8w
XRBbHgQP24rRA7bHid7JQyxfbtnaGOTzZu9QIt//H73djJFOyJm1lHyTyj676OckcZihDNPhawSj
PAW7nBpPw0wXqYHoR05NicwVv7tPmqYrlWIPoLCBODAxAfPeQ5IllzXciFNTvAtE3ZyoAfVE0fLX
97mayTmx2YGw1ZgtAx7SEicNbwc3+Ob4fG7RcHmUos6ZgIUufqmNMcd/GA15RGfkKTh41THYlGMP
ULn5AoxWr6AtlPbk9CYuuyGmGqdgCNhrTrKVgchgCWuwebyjsdtBFwAA6FglBGTUm9azCPfKZKrM
QFAgSoLJLfFOUEaVxSBH1OP1tow0T3rqQQGR+LUIzAdOtfWN/gYqF4IdRxTp8yBIeReLIK0wVk6d
LiSaRqp1tBc9TcBHknw6SyuP2S6JIVEsQbbZra64ttMplcpSp15dooXdjp42h9l9g2eNcXS4O18l
q41qvQgeOX9SZOZ6zKkrbHYg14xoz1gKIWAoSU2/H3xstveCpgH8rDaYWOnzhHLN6VmNj/baytaj
dOTnSOkfPU131leKz+moxBrQw7D+qRjixhcvjC7X1Px8yboMw0Y5c6WDn//AduAo1hmBM6ohfZuJ
SBbM20b+U28CxoU+5BCBBJMYsxa/cGVK3LU16Bq1aPyBU92cA2LQqkS0UWaSqOPrwZBnDYW8CaP+
8ksgOFmFD6x4FbvTlmWWYHPpA79lCji2lcwa5wMrSqHFEMk0FjbkXq2U+6Ev+kcoYwOPH1hftKky
44EBzl8vNYJAeeC+HjmGDpyfKzXLMA/lfDYV03YS4HOJ8ijIlOch1+13RVSYANHJJqa4U1/CDhbO
nKLHL65LeMKR5ahJXDi1GNFqYOlMqbiTdKRJrMI2bYxvr1Ov6MsmooRLqt7GkQo7y+UIOfMBjoUC
CVWNUjnsia0ErbDLHam13YYYeLoO0EgoBOpQco0QTSd8IDv6MVk0a5tQSPk63neD0G1rSM9NTu22
Ijun4JkGTuEWSHK9NxuD52kR2VF5fYpSJPAxb0YJln6HaQSzvLkqqrZ4WELXnZPXXuG2p3kBt4Ic
jiPabWOKC97TRguXwu6khvPk+Y+V5/Y21JlSIN5eYuDTBUTXfEwVNRWAyZ12a18AdkBAap9nxFwH
HEMgcIULP7tTAxuU45l8A8ag7so0RdZkERu7a7R7Ox5WHkuSEoOzoL8cgvS4XSJgsfdgDB9RdBU4
go4GAs1ukI2tbPn4jXDPTmm+vCtsQAozUYEB5Nh1JV3KHbMw71V54IWprVm/dcs9sAfRCGe9usOq
i8pR4wcKfNuWLSUb+cMoMtPLGQpXw73+lJL+/gFjVhYPlwbiiB3aM92JdRM3CwwK/ai4dhRWUiK2
kJrTDWFC1hCwcEDnsMygNStvEDdB3JI+NSV87LOAUrwhtodTk9koJ5VRaupYfS+0QnLk6X5LAYLJ
szeubVaAmsLawgWLuO3Qsr+TMcQ8vf63FhA0ky41IUeIzNvcCiYlJNFFjUkoRsT4AMSqovjbabEi
lHg2MaNTHE79kVRKJDjrz1NL2zv+P0oLmugJHz4AL2SSy5XIImW+S1U5ptgpvcrU2Es+DRBMvh8C
vZt9aTG89gQxoqy3XfZh+rB6DsjyMAZCAEOmL84iJEuZTwbwB3vZxAx8P6tDmglO8rgLnNn2CGhd
pQIqxD+tug/SPkmz2oi2G6UviZWyzeNif9yldFY28DUbnliPMiiaAdQKYqC8T0AzjeZ0O1zP64ES
vz3F9yhUZS3P6r25vLJZTZYJq5yi6evVDbL2XRhf+GjXdBAWKGYcifCaYrI61sKlllruWAb6ZHw9
SMRqHhxYr1Lu6B/bAxeji3XwYaTAMqrY4qE+jpsgFxf0d/EXkdH1UZPDkCNB/ClkkRErPcDmIpID
JdN84U+4+47DUTU61lwqE+JGYiVgqrpbWJCb2rltMpwpLL7sFaryhUDhfsDt9Hy+tu/rPOoKmFXx
8bHPUfxAO4veumzji9rPOdH0Faxq3pJitk14ZmrGu5XsY2VXy0ZLrcaNl7/wA6EI+fmxh6s+8zgv
n6Sv+mfLitgzQXjp0GsNN2E91K//1P31hJLC205p6tESsOHZi9WQ2TdYrWsjGrLDiY5jkYLKO5Me
dxV8mmyT2bw6l4Grae0gb1wDPVMmfuRNdgNHTTr1tg/PPmVPw2pJpCAKR45LKYY8TLMXz3zlxwaM
dB0CA3RDNRyEZFBpZBHbDnXtpie8LE33udIGQIYhNzPG/OVBdJZ9vLnZpwEWQk+F4rRZSFglb5hi
MxNdwBLLjIVIfss/xBThiD/l0kjN/lNj9wunitEN7VVeasVoJ1PgCaaINUkuiDIbsrmHYeGrVMs/
/7YjB3xqdYu3rJsLTpq/N/uw3+dZOkyrMpt6GJUWoAuL13g4USRO1O/abwkDAMUvhBOJMeB+vAkp
Q7HWyarWNzOxeYtR5dEaJ29H5/Bd+Y4OrHwm9+qodQrUu9s6MhOzuEYtio8GcslDL+JacdR9LF/z
Q78Fmu9IiviWawuy06c4jd471JtrRFb7np1xFirkQQgEmkE5sHbYfkMB4ainKkLJyaepvG1Ubz2Z
bKh9FSF7DkSLVqRLbJQzb4Y7JtoqtceGBv+Mjd6/Zu5IKJ1pkGUhSNJVzzjxL95RTCZKJzQA1rr7
J/QsAXK0sqEBTWf71otcu00cs3T5cxthv+2oDJCliRuEW4xJ4L9hCuPaXGmEVqoVNjNapbuaWISz
STaxHKC507pzmnF+utRqjNdrpLwIUaa88cqjAGLzp5z+dprUnp6qrZXmx+hMY5AEfuoEy+hq7BSY
Cb213pHYhrkJBdh6VWz9HoC2suJFszrm12eNppr+hJ8B0Nr3IZUbzzVD1dRbGzPfeYEWXE29p5gp
Gz+cdYA5bS7T8W9XmF2l70d2lbJy8IbC+Rq48JVPFvxDmWWfFBjLfZ+W0AsboLHRLS12/hekzFDd
pOzWpNNR7HdnU0UBW0QK2TaarU5g5xt91mAjWLO0XX/w+cZ5KlSJ1yoq3OIHfB0cNmYj0oWICEwG
d1LrWV142XluWVmcWhkgOPNl/mTbsEWKQ5aWQH1lTbovShPiw4QlmFHzw2X16CsmkyvCgYD+MFIP
60gyIlCusa7Y1F9DPaOc0fxlDuNoV0Xj86Cz4ZHn/WRKwaeKmG2AMgjdudkblVbWkuFtHo/wND1b
a59+QZgfJNDwEWz5PnvsCdNcpaW4eXwnAAG1XuJLyP9P/1nNCQuyg5bfwZAPAO/HsQGYuODBV3DL
A7TFKEizvhg2Cjl9hldDGNvtOaecYV4SlE0JkPHYO2IcomUvTnA2sF5bC5l3W4Vdn2RVb5jfgjEr
PIcqd0VOL2JqgE3AtZ0UwxQbDVa8SEs+tViiV/w0qedzk8/1IPbvpWNMPzyYWlx3xN0E5Pbpp76M
e8+teWo0Jp0VzJKy5D7z1vhS6eKM/wW6LGiwSe1+djPDWtmXlA0JJVyxmLngKzJKj4eqETxgbRfu
QeEq5mmuaDq5yRMBOKfVwKRtCyzrYSdRg87Lgcr6b/97vWTbIsItBzuPSsTpWmKvK42sqLLBdsNi
4kDPTrLhE5Jpqu8KdEaB5XJZZHXb3lpiptlfN2jxC5o5LZfVfjSWNdguJ92NN7FVteAYi7XrHyhr
K03vwD0/uTLJZ/DUBcQVPbyRbW8yraGu/LuSLQU2yLQQ9yeF0dBZ5dfrvUzR/0QozUW6Aa47S+3B
qCiLWzfDjo26D3YiyM3xWvtUDDUVWAikuC0BUUDTEXvcwc3fuoQp9bxBsp6QE66VItHCnYjJpTqI
JnHTv60Rn/6bQTfxLoukErKJzrzIXNQxW0mCTCQKfTE8rj+AELIl7c90O3FvV2a5Gq34drJFHJEM
sKA00c77AO8cAR+sE4xb2woynWOYixJEeoprken5ZGyy7i+kh7z7KxRuxWVdGA6Zz+rgJqijp7IA
xAuGfk8Ud9AWb2r4DYYoP0yRRzSALPU5wiR3sO4AKtctVWR7tcqFrErdJdSPZN2Nh8mUc01X21Mx
Kx2wOidxWgNQiC2v1RyN3wWPdU1zpjbxG24Y2fkiz0/QadzvSP2dq+DJy3TpSAOXJ27NxvHekkA0
GLbIc3Zbo/XaUkyEpTrJpvX3Wi77yHKOeNqNlZMikWlrufH1MRAZ8XTdmfdCPJZ4nJGyw5Zf3Q6q
3b3hbCxvl3TN/iMSzcQK1bFZuZsXfZ0t6B5q0Zdki8nDWwd4EYchGWPkoVJhZyvNnog1qRWCGaTC
rl9oA+3kBHuf0sRji7c9U+VOW+lUjyZMmPsxF762a/1xxqkCcX3MXXVcZ0smvIsIlEkvAGRBdEv2
N0RtNHiM+CQrJh1S7K8ozANVWw2+ckiw4BcQUwauoyFaqBgZzXSPewPuR126fTm86TWv4hfNrKZw
Jz3xLp2ASnrPdOY66DsS5fv8qe7jd1v/3jzqYwVFOsjanDwJGFN0UPn0Smlo2D/ywcTNUX5fZuCk
fFop50d64cXXeQnnKQk8GMnSwrAAR9RpzxPuP1SWYNYbLtYYCqeuuXUIjWY8g7GboJPtxY6ceHP5
i3G5G8DCQHXa8fX++HfBNoDVwkiOW2BkvXimbv2+9Wd/fcLTUdCuGyD4wEHV64IeMKppclemxvd2
n4Xro92XtwPKGTX2siMcW83oiLrb8CrOo/ooJh/65oBjJYL6oYUQ6nK8EUiC1p+UunHIcBRhmN1I
ZJKOeYSt3C5v7vsf+xKRQu09JX56pvTdIeWvuS/WgzIDjVm0VKMJkEMfamYvTNOYyJY19koWjyJF
2xufSPUYO4hbo6qGWk7yu91KrBSmheHE3tSSEjC+75O7Q+J04vYrCCmrdYUQ13JkE/Cq703LuZjY
hKDsi8w5laQD5I1yl4bZOCd8Oiqji1+0eiE2p99Wd3sVdXtAP1a/d9XTWLNwxU+JWqzjBH0W0xwJ
AWQwTiNRYcneJ4uYsuTMAfNVjDgeeMZkEvpW7cqjfhfGwjovH9h6idvjPl2TFB1q+h80Ip/dq2l1
yZW8xT1Xvdcj6wf9WWFxMMTCxd9JM52g66Kh2jayV4CktdB8gawSsm/qghFU+aJlPfSSOG9D4jNa
esfUz6wq7DdlQ19fwJdhGd6wDQnTozZYCqgZfVY5oYerZJDmx1kKRBjJUzaQTEvewczF5Vu1Epet
gUMzNBow1k1wkFoqCy9egi/9EdfzUg9LlFmAEZBTz7SX/Q8Up3iX0jnCDfiHkBxAhwoZY07QaZsX
sQI1d+umIUz9CK7Qsek44c5CWCutQqtHtBJjaGCzy8Y0fPt/0AT0g+AnsOXsn5pg8RWLbX6ND1hc
Yhpoigb+3UYcHj+V2c9TG5tXUa3vJWJQwOl26PIfCg8eBPkOQxi3h5MLBqnDi7nLEXETwqqkThvM
bpHfwlFQVrJlOu8sUXAx4OtPhisHvf3J4c1WKys3hYOJ2uJI/jPtg2+svL55NJv7wYkjty2OHa8T
ZAnYxy4E1Fx1+IFS15eidP5u6rPeGwSp9T7hC3giTtA0owpNZy5d2w+luy0zEcOr+w38Q0wN7k3k
QEQyHiV5SUd7QBe6W4/Xs8cD51CqW8GBhEwpOCNwBN2dwtZGJR27IypvIZUOMIIYqLcL+HthibBb
+FQ9SkZD0q2EGaCNO0JcuiPk5gjJY112LeVhjhe2eobifC5+v4lLd/4ADZ8SJxkx94ZQ+svgphfW
2ALHPmWZGHoBK7jb372m4V2hQv71MkpGnxFgRVe9yKTJn417p2tilBQ5YWpxEpuR0FNwLYpctA+b
WUPVbfpMbna1pcfzOyJrHqXF31cT6i00dXIgu2a85ixcHbouSUM0iLJTuLBWaeam+RU+oGrWXRGj
/n0hSDzolK2D6xjakiDrUkJd3URlkpsG9wnNlpuQBGr84veVdWpgmxpDobHaJJb3zMPtml4/Brlk
5xylPTpyCoUA8/HANOSvdYDIBKy1P5Tmjqm/7agBCP/0qBMA5fWDPzwT568rSJjkIQ4Gw1XSKI6L
pJyFrxsqm1wchTwlBWRctkZzkKrf2jzQ98obW1DeNd0FYa/IPzPaIuF+2E98MIRQ9BqXpOxHTU6F
9swO1kZ07QlAHR+vRfASwsruJoPsAolrROnYJBsfIPVDWhB21QuRirRjmmtAQWK1jA6ESYasq+sM
ZGlaBhLO4y5T0u3KP9XvgUFx0RFhjCof3HCvKfQ9R4aicVGqicvarXRfamjlko2Mcf72embj9sjE
FN4rFlAp42P+qCUl6z/vd57tbkTzg0ooFRgA0wHiXecKhNHKrCwQRmEGrqToldTrMhHCgwZhoj3b
4TOgfIPD9R/rYN24HAI3j7T2Onb8iWbNbXXtIPQFrvuNZBvw13/f0fbM5ZEP/y3P1IihwYy9lHqG
UPep5uSdTk6CIMb6cmzqltbEX8+87uN6fN6Ky+cOFDNkHjuyGdHL8zK7u7yI+Razh3Gng88+IXvM
xmzZdDX55P7Q+qUWGWSuuSzaoJwCbLR684ZsnAb4GUmR6SrdmXF7v+5cEgHPI8XwGeFy7V8D8vS2
A8wLIXKTesrHCgqV6xtRciSOgVqra4h2S6nOxPK3bczWuy5UeDkCOnbVoC4jfj0GicZBuWELkxlj
EtQVoai24gzNIFHqjEBUNWPh1cMKp1RLYzOJcg0J27NpgbRsglCgjnzertwXWRcWNG0faDwwZP6Y
worhK12dtgQV6Nw1y4ztQfljel27Pc3vFDG0lbsG6fedtDg0ISaCM7KtPblqCnB5f0ahiyqu6ZK4
DtjLqlWRFs7TaV8F4KH2HRUoOmVcyEYIOv8v0RNu07MO0BOdSRNBst8nydkHR51blLRWj65lEzBr
ZPWeCMMySLsV2sxPGncUTsJAhIuxn7xfQXmM2YuRWJMeERyWWTgHnglFWLKlNgRytic+xvBDo2rf
Aa1TT0avVePnNGDwL5FjzxuR9TkVpmN5+ehrLr07XSmMu+VD6juT3jNfQIpX/yUTr8OHwxjJpI3z
wZJxoBpJYaxi3Nq5hnGkH2FqfcQOUyzcLUQziugdUK066+ORQUHpob3oVscgUKRnXyZKZnU3Fky4
OeLhUsKtc9iL0Ju/wZnlx2YV+pH5uIxHiaHFGVcm0ad4C7XNGE65AEBRQAun0MnMMHh88PmwT6t8
5DhkBxsr3hKbKL68HbRNk9O+M5gugtvEkbGPARuqC8TEIii5GNWeivyxdx6lspMtxVZbAkLKSgOc
83/RSLoKWwrU7Fy7ibUDwR5eG9d7SOv35sIMhKYzUWe023yLCgKPH5r7a+VUih42oYROspnWU5jV
ljrz56WmQFgu/pJNoSxkZBniDIpx+RsFki2A6PMF+9ZRUPfFazW900tve5nQ03TzTxT9BireZ+6X
9qjt4K9qtinxIfowEbrE60t8RwWsob3DamXTvJDG/kZV/t4lr7DxlyCu8r9Gyms8WKmx3VYhAUNh
r4toopWIncxdPFbS1Gw4DtKLXwjfVCeqyk+UpyYIyp5OjOBxdeGPgwC2TYvQcQ6ngdnJYbeZmO0k
h980TH/oF9NDVnVOqTgX4Jmd3XSJ9MizyfylDN5f8V9US9vapTYrz8merCEK+xhDxF14o/RaAnr6
+bc9tm2UqrTzgKqAiFqqGUXRwzWez3B8FWp0BL0HSVRoZBFWVyhO+Kzot6gXRJYoP855+6CHGxLk
ps+G0InRXfsxHV9xOQPKASsJSRwqkuNHlAR97MmONLmWqRLrWqRF5WVP/kV1qSmqZeGqhOVQmc7p
9CHEqaWgmrEy/3dsVTZlrs1a7rcwFNWlGMjCiTO4fJY5e31mPaTODYu5Bip5VbyR+PgjfOHSN4pY
7+eqdXdHyG1ZlX+4poW/iFWIk070wqSqyUB6jz4JBXbqcU+BScPmJeSJmH5KnOP/mI8oxbfh9Aph
BsDNyJDLn84ww5wJASURrCIHna/KJNC/XSYyml/sIX1Xgpfo5dxBnnd+7NB9wu/Ip3WUy0hJJUEr
sAFjpXINRYAgzKWtOL5Lw/ZMhaaXhvk1Eug43VPzN7MwR1bHxLzQl/z6j9PJvE0mkde0zQjZaT8F
m9fgY5jrvG7g2DxYpS1qRAFG3Th7uAJIPudBzSS1ez9SeUXKyl5Q9OzA+wuHrApYQXJkXiygu8tf
c/gifrsXPZWHjbliIRJErMFLtDLZKx/8L0lyNE3tITr9zWNzcjaXcRhbLEQdSYEglLp4yrhbliK0
4emZqDNMWklJs0YV+jBRfCgMKI8ixdy/YbUzNZAhz5DELtTmofsska3q4Xkm6NA7BTBsCwwrxgPS
m26CeaMkwWdZN9UviBYWN8v+oPu3CYMoQGFFvPnji7oUGU0bTYCyrDPDq2gPL8FKibNFeLUQRwU7
cKRASAN+uxk5T3tZlrq858Yl+acHj2H6Jt2jiinYiIJTs4LMq53trgPy567fX4NolVhQNdJigElt
krsZjRlA924AnuDcItQ4eUCBnOfZ3oT979wruRLyTdZU8QDETxJ94v2TqbFtIT3EKdZRFZEYjELw
Yqz8+gUw5L2u11RLELZS40Vwck1UADYYMP9VHK3YGDCSz10N0JZDGHDD6CTjoC/5aURJYuzH/x3o
hBrhYwsx1BLgpEP++VRkhfjOcqpISV4gIMV/Se2VgHhFIQLvQUywptwzOuJ1Yc8Z4BKVXPiUeyPz
1m9MoTb7yUOETAmUkGOMNhknAkNmoQAg6CWCHKjyhUXlfjeiZ7Fwn1GWyuEi4vsNsKy2SwF4QJfq
tyIrIBhykzTdBjxmdQVufCJMif1vFrwSteYPtl+GVhV5rkDczS3P6+ASpwu/ynAGzv01YwpWzsbV
t6ZJTaUhTLrvlSKSIOUShJg41j4epnNz31TQSF5q2+c+9rfgkfrXFMKYkzOeNprHhQzaWg8ji4QB
9kyEvOg8FQeHQuIKf4Wx7WTLmUtZOVSRv3ck5ZScTjtXPQ5egu4q4O8PoBzcJq+I0hOOerZdBikn
hXsFzTPITfI+z7JvdnImMiryPaBok6KxNDF3udLQuso/WQphNL7UcVGV3r9qoKMFQx05Z4kACoAs
a/yDXdEO4sdkMXGv9RD2W1LTD3LnmycaLLIioRpCiofeUvtAvpzrpMDTaQOKGGJns1/y356R4GCL
QFpBKPf4W4kk/UtjkXieo//56us55bCamc5OdPSCIUZuo2tHKpkykYyq39Z6An5DotRc3EZLwM1K
pLNuTPzlW/FgGflM+PR+gDPb6otN5tay4UDNaBZFckGYsp9o40QBImd46IUrSbjGmDpY8cDFZiJr
0YeDelNYDzXL3yj2HX02RG+AWO48G0H52yns7qZqGVtT4n2XT5qxovlzaKqo+kOgm6Fhh0DOf9VJ
ZSC4ll5SJg+4IC+Ji0ogfsEesoav4dd+V0Z1tV6hZ6AKxukeKprJCcmPFuwfKBYIeNLz4AixtL9X
iN0Qet6+ZU1F9kWYsN4oSUezO4s/AUh2Z6XmyEtKyVoh2+U/mEqNnJl2ZAsADCfNv1xW+8vCL6zI
iMLIYW7XP2rnHiZ5wmvwYQFVWsSvb281ndfIW5csy/4gB3qS87Jz6C8C60vTIVX1E9WEQIZRrtfk
j1U2/+mkvZQQvDhU5i1a+zGt2cGLr3huuj+XzT/DkN/Fzt0gFDTfWOqeS5J8yh+dyV36d1y6al4y
yfk0JyjL5BPPAdHl8F8KmJ7YR+rzioJK9d6nObEER0y6nQhqeaNSF++TrmQmhTu6OqZvWqlEZAw6
Lg9ENR3l0Q4Vt/LMAoqRvi5MH+49Ogxvh0mdUJfWiGmhks4/5TVmmauffnDTcIcDkbB14cYT7QZi
OtnVPfyUGx5rFaJR2eq/OqOIZlfTc6M9s7bWieBiMnyIr6FTLWW4EcDowI3SmjHPnemBDG/83ysK
2+nCgPwsXtftLx81FFZR7olWopUFxCbLxdjyCd11F9oMIBcroLGw08vK4bcmfNWh70AG4E0h/jWm
oKXGGOrcKDBRaSw5Ho1SSveNsRNKaKTov5HqOYidVOdtwRgvyTjNM6x9Qow3gY4qd6WxSyqFzstJ
3Dkz+g00qNXwpjRaZlz+Gx91YUe7gtJOXH86rnNJUks2bZpgDkOjjLMVj2JoJqyhB+4SWVk6BlSv
bYSX/5gR639BAeepO0hH6SLPJU0r8awd3H5TqUQUe2q61V7TR6D9R8XZseTaO8l26w+9Vz2LghrZ
7jLnY+5w1yyVUwslwUONvJC0minQjtnqXrfJhK/EdQ6WlDV60q1fDLyY9X3a3mlUHUJYy6jRMhTF
qCOsvVSvSzgjreyZpFxJ7Yr0sEKlexGNC6XA2bCTL7wWNGCxTNV4lv1kdUVvlshUpjtgXoc5h/F7
+e2wKfbr7U0fGfUlDjgptEybY4lCE+0moqQbgwgW7hUbLij3P6156v/xjeA4hlirjANQG1MUPS92
aDoI4D+3aJOHghP5y6uJvHEeJ8IJw25Mzva+Z+0ixjUYbDjCzEB0cKNQqw6JHUo1LDfRoG3XJydg
xunhZfwhoC5R/0j6YQ5DYyyd9KoBjaKQ69M0o2dJU7n8WiyE/vNKzFlcEdoE54QZv9VcuBCPBHlh
n5lKgjApZTBS3eB9poN2cCM+O/cn2pEefwDl8Sn9Kbnr2BIdlsfVQ7W6dMxMOosYaTtvdjPebkh6
oTyUyT1vCxQ8qSx8YLKNk+owBR//iAXnErC2UnkWVZZHTSmGcRrXpneMLLX/JlnyTnPGRhMRmGR9
iYjTkAhY9A0vuB2noMtTKqJWGqlUPgFnhSrCdaIPX60eGGJA3SG3lAIn8k0xLVMeRgbFjjV2E3s/
GwWeP0WH6KhSDDBfjcJEIxtdGolPny7Clhx3wjURvl/HGif5Fmoh3hm4tkQJYRMWTF1edvJYnAqB
I31F5kYhiav8MSIukr9fTYcdDA7Z7Y8+ROHnOCS0XPYrXyDqJSlJsVaKjUhVOgNxC7FP4rh/qN7g
2PmOrj2i35mE6CAXFT2JpcQc6l3FRZC7n/TVaG9Ge4vbcTDhRdom3BXAl4ntYqlMJvuL3Dey1kTi
xr2fcln61Wn/ebbnAPnKdsvifvm3Y/gonV98nQvS7opeAreIpBVdv/OIEm7myztLS855mfd7VVen
2XFIJEa2hl7vd5DVYptIXFANtbH9HOs/zI6ocvY1GjhPKKkYd15ccHxWq3yEAneqWi0NGs9juWyE
vof5HShfvx17eqONctTxuos50X1s1ZaSMfCSVb3LSkxLw7KXBMvUY0oRPAfOPqC0yr4kIlMYwH1w
Us8gjnu4o8dJ0AMdwK/t0hD4CK/LhWraACzQ7jA16Q2HRxa7N/bcqXNZkKWOMf/waa+PkvG1OPeI
nUeFVhVEh/3nPNFR5ZHi5WFSq8Xf//1FQ8oGk9MLL+FBB/2+PMPURq8mw5dTOCNvu8szdVYUenWy
hXEn+JY3zQ4Oc7AtsMGRvcowiFjbqPx/MD20VFoHJsHtvY2YiTuTdvc1V4Jk0SRl9qbu1aKKwrl0
7H6EfrLAz5P/4GVEvykioW6M3lHnKEKMwyszbXX1gOcPfHzIf9z5WTH5pZcFVyFqYL101D92pB7K
Z54zjl0wz8PxsLo3g8ArS4h4jccKBJADK+PM8bZ2OgncSdRCnDebB4y/YlBDTM7Y0KPgPGaJyGwo
8ShtuWfLGda/gAkbtirPCF1c8G2W2HtBevU/FrUHijbI0SMSv7/kqTOSJbwu5oKADGHJp78gqa/s
5vFdvv3EWoSElsu6m9JhjPHcgWleR8UxqjC0VGmtrDsLFv7UrbWuTGj4I2eQoC0IYzDmdsVeQ6WQ
I44uKL1G/SkYLSn0WQs2hiY5NOl9VY2/D49av22i3+eH/YBQbRYk0leEHW/HFz2TUtnJ4+MtFyWg
lLrD7KgOK5jmi7WPM6XCdEWlcUwHcR0Kz+Fuj5wiFLZcVNR3dg6ur/Mys+vIZJ1BZohcHlf4IApL
kTGKNr5ynkMS1VE/SByJ139H0DMeMmMuyKcovwHkdRnpWXapF2Q1d+XZtORJUT8Ja+hFAgd1oyGT
QqWldqtHlBfVoAgR4AmrmGJP0gl8enbKZoY7KUCY05bHRRWgnWHFWIBJfIMzW5MJBu3ORX/6UQ7G
4gu6dhIWfydbfuO2Zq3x9ZNfsb8TCjjAPS78rIFFuSMM2iKkZ32EUQpOgcFGC1UrOdldg8gW71KD
Bl7bPrFL5aafL9sPtmeccOX+macYm9s+VJeEwwEtV6bvnwU51msbZs6HgO8o7T6etPwAAd+Mq82u
/yD9dwYnxH7qXeBl2J2+gm/uZl5Dw9Byxz2hrmodsD1A0zFSbI17/Oy3X+6ohMXHwuqUUQzHP7gX
iEvjR67w0ie02tH8gq3weyr+A0EES0RXatXhjkiyYH8g+R3ur5j/ODwvzn5nJFJUKm/PsCCJGOfv
N+EtiKXKRtfrxSYiU6sVYkIRA/Wpe42dUfTFOQ69d5uYuumgUuj8yulwxh5mG87eNnhQ2bs0RSUs
wpFrxtkO9Nep/PDs30O//WB+6LBK/TrCUYQ/M4ElI9lBhNY43gO3BcvL+zcmzMhNoNxXapdmsSl9
HkdlaDeAaLK3t4bRuxnA7ZQRfev6kBERhCo+ky5nopZ/AVBuERrMpZpORRQxK1BWGBiqq51LcM/6
VUIfc8WerJFtTQ4cUzMFQDOcW9aplp8I3M38EU8clIRAg1DLPmzxxhzz84jtvhiPDOMhFRjP7ou6
k0vhy5mRqB0XJinj7rAfBb1MmSzc2sieVfcsFuqSRbSMiUn2QGWmXGdznQ6Tnp06ggwtKokxm9Pa
2b45ZxSoBPgrRkaVwY9Mh8aEHLWZDN/9NJCOxLFSN/O76zB/YEakmtN+IHVJsJX3S/Law0T9sx0F
leM0Mh2brBgAKVVMbJuSmMFOoOs1N1wxcRMGcLhTmNNM1D84pfJyUiZpFKv+Yv2PetuORWrYLCG3
LEhR8UebNf5LmdeZz4A/5k+ISnoBITbwrNckRMBqjnLZKb4KpNJiY40yvMMTK9GITNgc+G0Zlb+T
WYi199t1DcsPn4PlgtfL1ZzCgOP01FdqhXgUYA4uUP4DQ8V2MVBiMPAz1rrE7F6hKRhzHh7p0fKC
5PFS9ujTUUMXzhC3232sANHwJgEXX4nmUiFUpLt7gI/FRHHtFdbzQTZKamkTudwfALvyE03DZrcM
AKVCXyiY/UBiankeMZoU3MvYMd4sV6lIu3OHrYjoVKhXM8jkEXSLBMwFbhtznAIqSS9de39FDNvR
yk9zuzADAcaRSafJq62lkychArc0OezP8agInFqALAyBq/ws/XHBwrc9634QgnSYMEDDRpyb+aRP
5OMYCtcEg3jniLdw/UePpahg9mOVRdke9Nn74onQkzT+hSY0TWknjX2K6lxUql5OX3TPOl/mPIAI
5/MOl1zzqjPAcqpClVV2I83lc6HL1VqF3oobGsiRMdlOtcudKcp+8DjCEBSZhxIWJKhLWdBdAKUf
plARv7xa6g6c8EI4dQlDLCFWXoNXbxLhgc1b9pQdNGzk930EkdLKD4GWz4fljdEREhTVII5UNIvh
GbbBLco4g08GcH80knNFoZx/kVrjO1YqM0a0mdWCdx9UVGr0anWE0v0yhcFgG8Fy59DoPm9KOgFR
CHep3S0+sbXlKy25i3/X3kCXciypjXfHdq7KAMNT/PUQNa/tkr42q303thMlDnNKBXo0yd/2N4an
mlXstoPRK52bizMcfmKJerj8vbOJlVcFztkzlRi9D4YGJlO8BfWj1jgZvD2jt21Shg3a7ny1Svmz
JbP95Npk0oKa0QHfPwOVWxC3ydB4hiiadyFSkKmgpJc8FpaLurBCT1aDgcl/EkFWLzldefs4gRmk
URyOK9flk215ndSwdbgfFI1JAa9Aus68GHJfI+LRhp40nqPhKdr9WWwPxC257aAqdr3SXCBLWWAa
DmxZkv0uuEsLp7/82g6Whlt/WCaVst08ZAVpqJjlAExxGc/MW0nl9CWAtGR8X9kmLjNk4kMHWDbK
BCFepsMfqEZq8jSKe+paxTraXE26i9gdGIkFOlnxM5fEoVRMOILI2zt8Oz/uttajHFDKAOgPprSl
MYodskyC8Gb2qC0lOIP1ytWBRZj+X7NeG0508Vo/sMgiw+GWYrT49tTeZK3Ogdt1TOSCPLt4NYx/
PRDzDglHJoqLxcPnmDzL5rWQFUuVBwFt8jUYtlvuADA7YnhQuk0IzP4FwAXLOho7S8kU1hliavdQ
3rPStOOC4KefINEih616lH0dx62JpF2eJToeAFX9wsfRkTScydxN3kUSPQxkS45Av7zFpqvRm8M5
S4p8nNoMsE9/6qrK+Hqvanb1xENuBwyIhqQigwtz5BdRBvBvrp9gM85r35Ac5WZzUAQJtgmniLxo
xHzimoWiPOEtevSRlzhWE0W8bJCq8VswpjFMZ7mduxe+lDi+6A9g4oZCqwGoRQF7az0jsXTu3sDA
NvRY68dcaLXkKb0Iy77W6zFWr9W/J6Jeti9/JI2bVBWNJoJ+2GIwiQHdPzMeh6l3RVaEN34utGkS
bXIMvZeh4CXI4UG/htCIHSSUt0tIUXpQI/ctIrhYpnXwcHS5sncDeocO4GCOPTmmSVjtRsxfy3M7
E4N4z/pXVD2dUy4UM4nVRsBEwm5MQUFC6d25NaIftxIrvz0hW5GMnApf5QWBuUL09bL+882lBamx
6ONLv7It5iZL0GPAb2ViEndVCI4rPjG6sZYxadxB+tiXkahrUC1M8uKB1IMpVsK3ktWlStnBwp0H
qWgLOlOIQj3OmGXAg7PmqSW3CCZMkYqrzTk29GbBZ0q5Xiexxu1YVUob8cimpD8BZ6YdJAxj1vAA
/yLbuD1z0yKXBS2+JCP4Zzn29EfClrZAZ4PmqAV4t8rZzdWBY2jXCD/9wng9E5caDzxAAuKA4uZC
XU+ehNZpUl6n0UfOzUagILMAx1xxQJnbcy5mIVp7dGCIDDzKoV5etHpW31+N+nNLOm9VmSAqYZ+H
YO+TVJNzz+lBJxCJJxFeVX02/7NLW3IQBcf+d0IWehbzgA3lrIAHNTWrSHl8hvHGjGCzB7GyoNGM
1kDmdk/rbuAwvCmCNBwDtgiMAKnE2D1N54Y6x3eyq04bRFCA6vr+JsH/fSfUqTJC6gq0lpd0i423
KaiEIyHJjkESaIwSZrWrs7aKYRjpmG17Cxlyc4/yDdkRpggG/xuxiTB4NwHGC+GZ6m+TAbNgGSU7
BtJUSVVcuyeRKPn5+4VwjcdhzGpwa2PMsT9drOkh6Aifd/vPfjBflnzISMTCipXBdv+v3W6iT6jf
HmXaNP4aaHoypc8DIjG9LgpIeIl8CtOhk0n7QjNtRf3SLWchmm6FnoJIW3d5/Z2gXA1Ztiwfqx/x
W/AbLVJmlWQ7LD/oji3yM31MOtfO3LjHyNjNngj4OGw0GcXxLQYp7vkjqTI+ZOqkxb4vgZl1hp/W
enj8pJj2+xf0eP9PtH96lCEnHG8YQzheqfS4s0cSz71izZ/8PZvHItRfNr7qyh+pTQeewjrJ3hsg
4UMsnN1NWnsoSCMw1NkoE+9XBCvfGUlob9wfw+OlPZoZvEEoUisyaVTIjTPrFrkYNXS+moR71zEd
YGJ+9aFtOiSYESi6vkHYAP57X/0AomexzBcBXw7RsVh7KaLPJ0ldmQq8g2xyt06Vi5ZCrCJg0efp
39r12Rs1Cph6Xr+N/vlw+yrffniRJYU/hEBqHfHJWew6T2QIIIJpL9nStyrC6m3v+YXXGhjgwhwV
3fESSt8DeYFSmr/IvFDdRkofWdKBepVJHhbAP3N70hjZAtnGuuNMMswN5cCmTck0vh4XlXC28bEH
Gjx1XMkReDSM7TqXQZz7e8xfyrq7ialRc22h3Q8ZvFq5WWe+I03vUf/O4B02/q19OgESP0AufFwI
3flTL5Fb6zJDxhZ/ZB3FL6+Q24Odh54gJV9eAMfe/n4nczbWCN/cfbT2DG00KU1n11LPJyqB7+Wg
3WpRfcNNT8C4QvLC7v3EruvyZlemVIpniBumxtfmnUMv53NRzyETxvdjZhan0EM5GqgM6V8gQcth
u4rJwUVWoBLJtR4+v8gAxvku1VJKxULBxr275z8JWDypIivUJtf6bB5LQA+CeBfWxZpBhp9uRh4D
1hFWV2XMq20PXV82MOV9bjYHYLRFLkQJgYnnaEPllcJxdGJQrN3wJLVUxSZoL9Yekf75xYJMyj9M
drf8BxXwZws09PlunYD+HpEd+M5NnxSjlTwY1H//Q2GeNrMHac0B2HZmqJuELfkuJA2UiEZdpFOG
Irx0XA9cQsdKv1vhlYgb//4IdAGGLk7UPkhCnyIBVHa58yS0LmWQ3oFhOqEC2WYafa5/XguUoUtT
sJZdquRk1oeEpgXsCBJNXov9PcwbkwMH43NsNMpi0KhzY6cLhfN3s+iaa2lMi0WWer+KmF1gyn9S
0AiyzR1tMRtySPtSjJ4LlDlnBx2KE6b3eh6XM5FXCOiRUeqrRjHlEHBGVxUIaaf77H/c1SXHVJgD
xwVA8vuvUdwvs20J2DOozLtD4hXIFEqM2Uwt44LU3myiDqlzN2Slh1KE7vkm+nqyE7pUuzh8XT/j
5wQYhJSfRjemlRLe/BGmRXbeavK0yIsZQKV+9pO//JSzxyypxJBd/33UhiNe4BdvTwNkMOqrn0uv
4vvVTTx8ORx4d5bjCbGgSkgAFeSOPNZBrhlpUvA91DKupJVeWV0d49E1+NQI4b22RSkX+rohCVAx
8BTudoh9rfaVIHt6gbqflBXfrvBOasHyhLBvKruY9X1lRmDnB9DwfX9IQ33+zjAmTqyUVUaMWV3W
XcNkzMrptzxT2QnB86UMoa5OJBYZyibdxfAHUCK6Qg8midkuVyvfNRUKtS8X5lEffe134VBMOtY/
WwkiSMX9A3EgQtxI5sSU1EKBjW7ROAV97xcqB4Mre4zrOZwqAV5hPp4GNifWtcviV4ATeQZ87kWk
g5q7EZspAUUFFjubXhHi0f0+C9YoUplno8ZVVc6gC2ccIanViW1BbH0kUiuG+Y0oiB9msLNCrE4o
2ZxDOb3ARXAIzyCQ3AR2X/soYaPwg8J7dc73pElbEz5iSPAVl+LdYQU4tMkRfcXAwfPzyxJvZcdA
73S8x/MnVLy4+M1cn4dncnc9for3BVbQTfH8dXOmRv5RH8d2T754h7d1+1BztNi4bBbyz4m7SF82
Vf4ab8iU/V/rkp4BYtpHs33SXUFF31gy+ytA/Zt93GbJYwUCVDTKXt0fsADdrh89FfI3WUsEYQOK
PITTswFHHh4FctMZWdUVkgdeaA4O0UItjY4nOYVCNCaOKp2qxoMBsZvTGotBxx4V+5kqJkG3UrA8
xLlBXVt7Dc348fyhiVOqQ6to7qzKg4vvAsS5XUZ1R73eYXZZUmxkXAlgDXdFkgJ6m7T+KC3z0zOD
/bxF4Wr9y7EKGlHPi2QD2qcJ7qA+ScMjzCQF9LDmtdS/Q45bfM46RBSBz9eW02Mo5jv4AZGc6m8b
K1p30WIFV40GwUqrk+L8eePx3Y07Nl4lgpTD6KfkzY86Cftq8pxkwjs5qFqF+8Q/pxntWn9q9m7S
cTgaQ1R/DVwivdtdqtq6NPEmEyn/VtLd8m3OCzhDcwcMqUIJB/9c9XGuz1vQDksKRvpAZ5whhXSD
BoHkUMQCD1a/ORw84vGEJTyl2OmgkFpluJtZ4AC/saoJ1xN8LQS/upA+gObx4nvxTujY2/yG+Pvv
YZMZAvdwdMgy/2Y/rDIjpB2LfI0wxabWkrljQrYL4iOfxyagCWLwYc5HwEuNbe9mTF6BNLQ/YP9D
lTzfxAAO4v3+5U+gPYPFt+gGyP2yKUzoo7EovSHuQH0M34WmAGMBfQsN3qHg9JikU2CvjpWGEMnH
3RKlFdKNt+ou1jEn6uvA7cooPQGT2RxqpNIw2siGkHaym4V2Wl5NoerC6QZgTQy/ZN9F9TdXxWnd
DONbFMpK/q5DxlCHZoAy2jsbBJd1An0KBsngdTnTUriR0I8arQBYqQ3qvgVonNJJwmeHd25oeWlb
jlq4B8/tb76fkrKGddUTbvVBjTOZ/uff+pWolNBAzXNZwKgAC++KAHz/BqPnvHTmUcAMwLiqdimn
8WXDb98p299Kh4ADN6XF4kMJbDVmKIDEd7ROiTyC78enUh/dq3SkZCwu4NIoQpggmcSqv/5M78eK
Bu6lAKKwLyYFZ6iEuWHyfdFWzS67uOf2TDwBt44w6Li/WMjmGANPwrmjVFM6CMvNDWTpXRLVIeqj
12KDbz3xmZI7lp7TSqZPaDw1vAMWRN6c5gBvV61Bm1Qxb8x6zkhhQagyXRKQ+gJyo+wmmyC625wz
y4LWPZLPgwa7xrhMILCXowLwYQSEexXZTqCXfp8Ew/bALsjkcKxLJz3lQvr/ue9JIBqfEqZU9Yuf
ceYI1yq8mFbGTSBWhxIY28TpChf32dotT8xay6IMvAZ5/jSYJeevBoQYT9kR7FCRHRbd5AlwLTy2
mTEywg6whcjrkU387QQbcU95dXLMr6h1a0if2s24CBV/4PxCJ593X3g7EXV1M+penluT77OLaRsT
VKaHHtCbtuMEBNqPZNF8rKf0+rNe0x7b1zeMI9EimHfuJiMYVqIjDgaxV97nlGeTgf+r67ItHYwW
Hi6Cp4bucc4NplsSo9yAMI9vYzqyt1RMtmmQm74nmeEpk6NX5InwKe8m4d45KQX7dBCCl4YZ3cNz
W7Wyey5tM8oHslENbzJ+36o1TzwH3r4UWegrATxEVXJSRB45w8vK8eC2C5zFVY2PYxipMxezKXc+
OuxR1Z7DPaa8V+4o/wAuAsu86VlxPJqhCbEkkO55MI0g8HRoQT1/fsRMNmxxtMCzDQBy/3ZN6s2P
+x16SnT/DuL2QV25eUlEuq0acj0IAB03atMuf4uwwQhH9Isw/lR1WE+J0a+vnGsb5KE0Kk8E0/zT
ucj+/hKquGuUl/4OwfqQQmMk3W3u/W+hKu0AiwntA3PSyuCy3QeAn534iorYtalWyYp99a63Xe/L
pU82zczO9hjWhwzjU4GaDjqqKRyJM6B3jYb+DQ7UeTrT5tr/Dj3/cnQt+6VltnbApyJPIw+xQEpT
XXQ9sYHCRjvPCRwvn7n0Qv/pNEJeIPMQIlSR0EAmO7Ryk0MNun/cNQhoW7OwXwCpDUuOun/Jno22
sL4YJPh2JOZFbZkH/hSf93khSrvtA9Lka4LYEIY4deuZfRBF/hNOX91rXKcwcD9TMb1FcP4l7mBA
82iSE1YFhN/vAFJT1yK+Zs7Mts7Gjyl6MSHqgMJCPlSgmnfg7+Z3px19cyWlqkkM0YI8lZDdB/SX
TPCPTMYCs0Zo7WCgCCKj7h+S537WHfNHCYzoN0GTE1e7pjRjBERAL2QyyH7iBsaFt82geUB+iZRK
yIaOM/c4OBjeFbtGSsF455ZJo0qczCj0jzg0B4/vcnu1t4sriHRY9iig1N+PVwp3E47ysOY37vTn
LNX+WwTBHsMLDmaMfVGhJHou6loucnbbb3maMp5vMOEBOKjs91r+0ogfRdYmXsjyxWvg3vZo+Su+
Gc2gSTTLKyshdaa59apq4vSD5UoMgrI/8PYfAFCQEBYO2sx9YPSZbOdqGbkwmPAzaIoEY72TIh8p
02ij8uvcBRVJ+zNeL1pgcJcwbdiF6exKGuY6GzhtPaUDfU9NUdN175GhvZUc9HwpVsWsn000kJiW
p3kln8hPCVNp6myI8JJZXLH10zasRrGfSqD2iKQOx5uXROaXc+VIfZcsZjrqsoBGJNi849BSJHjF
K66tCh/X6NjvjdGhqVeDED6eLOKtDN2PGJ38S8n9TQlhMpszwX37sQHwauMVsY1hQ/bXDNe5nPCM
XCCGR5DB1kku5Gc8/oTOusbHc+yJ0IhUI4xZsaDo3mwSb2kQG+p4kic/am+1WzxclJ1cJQkOTEZv
uDIazDH1B/EI+f38V39IqfbTL6DmA6l8u0QZdcdqvUuuOTMwDW7iVMpMD2Z3CAV0NhMnwe19GPYE
pxF2CysOWe0PWZFHq0/dhJP6oSyrC6k0uUSga5M1ILNKyphD9UY7k6vPMHPU0ipiWYtcv/gfo4v0
sE+duLUTRcY0VvFom4o+mG3wEp276MROKLCWKWyj/iM4O8OjGPGrGnXK3ogqVrhINPCnp0Js8rPr
nlAfZ5xZgRWQfvD1mHeSS64J9iSDN7j3ES1x3PcMvMdXPQ+zwsVE1Xyt+/f9T3WzPXB55UrpR66l
chVBuByAWfyGy7nE+zI/tWJsRrBhsS7SJswe/I4FRu2MxY/FntQDUIZWaY/lcnGlx6v6r+NrkRDW
p6fkS1AJ8QJV+yTAe4Vz2z/zps8awVHzFYagqWqh0fqciq1IJoTvDb6SwCnuwXNz7nlbpQPbVWDm
Bp1kewg/R8J8h1L8CJpr3iNk7HCHQO+vB22pwKIesQqKWjM9Pk3WdiIbJJ1/sL3ITAktA1VOohsw
l4gsUJD3pU/abYUFBpGRwt0O2rf6QJTptTeEooyarMneOTSq8Y7vCslFpHSTL3u+v/V3o6zFIy6m
uZQ/eEBKMkjbylQd6YbumFy2PcsM4D3VNjv+54JG0hELqo/MwDf0GZUomDjyPbLOp9dIxQKCWJQj
6Puo1gWEOr0yQNMMl7IjfxlMPX1jhqXly7yQQiPzQlpdeJODgnaJtcXy8lgNhroWwXcKGFBrSeFN
u0Usj43TtpgQT4ajqvVjTKlrX0Yis/q1JwM6DYVYEMKp2ZnyM9YENKOmxaZwvGRNyUuKRv62vijF
8pSGmtUQZzkn0jL4s4yCpuTawRKkWxa8M2JyVuTwr9bmoKc++sksVv75s2ACBNo8n2q+09nesMB4
81pS6EBEEeFfgMOtUo42ENA/bg+oUaSD2oKmeff3kZbOzLzDNeugDZlyWm0lQ49RS8UhmZ9BhezZ
AUUKMptmA8ou1Du3H2XA0nzDsswtfM5XMYioqUmcfLnKTgRW31364DXi85Lzlswu+9Ub6HUDM+eP
u0GpMOI0ocuA3nNLYB7EF98KwrNrbnpnj3rCsf1puvqt9KiJxnyO6AzcLog7CIlpsFpGk0VUPrIu
VdIAe1snv65cycpA/R2u5OZcCmdFCk51YBnHq5YUNL1PxgW281wR7DIiWQq5GCY6FOiXvtkTJzR/
auuRDm1eJsGSJfOBC7jJGt5/m2rJkBFNCWCLAm5ChSXjBySfLmd9sMfEtUbfsgpqFz6lgz/vi4f6
kA0uBergbw4qD0fK40IISOxrGmc26UQOoNsrV1myC+0ZqY70v/EycpefJ0O/bnzUV4gi0UI0iFQP
2mR2xjaJZGbaNRSnVmN8O4DgMuD5BPmc+mqWgVAqbPYQ9UxagaW98dzxnHqneqNiM1DoRJ/mGZYZ
IMQ6PE8a22kv13YiY5kqhFDZQqOe6Vft9RF79D88L8BlKD8Q+2llzawlIF0nsLqGrtvGPf9AE4TJ
8MIILo8AyDL1omDpmAhEv9bch31dDPflrFeC+2G5Y5U5VC6KML5yAfRXxTr9orKZcAPkbhFQoDZP
LjKxiws8uvA2v5O1wkNBKqtiFiMrcuw3A7qTa42V2oxCEjhQN+WMjK2k78qyXf43Uwipihy0Oc9V
3DsiSedhBLoGQN/LENMwKqwHlBFLFw6N3tqPByB55RZWES//KZ5uoD8sZ18yy0LQsnsH161Hm8Sc
LIhc2jAcpMRacZEyHmi84NdJOe44D1j+8q9+erl02cyVccjFYE6zI8PaalysohlW6HMj48Cg0jtz
WzIzCvjujgz3XV0BKsVkkn0kdhgKhwRyZigJTt5u3KsDk6waSWOMBv0ZDwVNChbgnQMZ3TGmDdrE
jdP4RHNjEErBFHj3JV0s6hjaZ9DAC0KdiqNu65XvDVn+GTpCCReykEW/FOivk3ZyUPI4rU/1W33R
PTHzzkIhs6qTfle3IX/XU3rmT8ik4n8f0q1S0NvyLVi9fWjjloTy7tOUMNNcDsbNkkimCmPtTb+e
ruH/8J6ZjEPp734wc4YP2wVOkwCuEez7DR/kIUNZWkJssTPamAlyxXH5vGfymyoNubswQDtu+1Sh
yPj9/LI3kaRePus7H/dOnanHFPKS4WM8qWWZ7K3Z6sJmWZgO9zZKtyDIcNY4oVsAJmC12bJ+EbtH
C0a07g4L/cSgoA8aCPrSD+WMme2S7RMDUB5D3HKSagcvHsCQQbOqufe4j3FUl7Pdhm/xHlrFgjX8
Oh1G10ZPp/eNF4MAGtcbc+5OCDcKCZxBCLlFT3bYPdklXxP9hCBm70kzYk6JUos+H2XzgM8Cxc/P
zP9zxBrNINIaXJWB4EOlclMcGOeYyL/MjRv2nGUVYxvGdlpHKbsbv03JiYZ+lWoUtV1CocVdqEn+
f9MfNN7lzsWZIEo6b7OUlG6sbhBK/aOfLhXFO78EEGO4ZaO4dxPoRkwmS5vqPal0OF42rAp9tA2/
BK6n1kGq1zcnfjXxlw9N/Lk8W7Mz9Ha0pqSffLzEyrEPz4iZclijGGwPAcQZgOzB03Wdd9yZ36EX
Pz21NNsw07e0D4VCpOS71+2yqag5XlfBHQy5mbm8oljzfucLjg4ZM0mZBS6YcUIbfx148CkYtXju
UI935GsGcTRF/k9wBBdeHMZjkLf8u7GZv5H9w2hnxjPuxunq81lqg3Sramrk8QnKq7BVK2o8drah
A3ZH/IzkW7yKuDzd6BwwYGnJsgFY69h8PAwAPUP5O4E7zckayaSVR1xCyI/7VeTvcFPypWfGCtBC
uZvfzPO1EBvAfqOmIOEAztBNx3AFzhZUfgiJdyPAvu3jv7i9c/dm+pkrlqCNkiT1dEpKA1hfYwAO
D7P0hUVg0xKfeOeI7R5TIfhqClxgxSI14fO28FrsU3b42fEMES2gF0Cu+P5ZjIskPSSGQaVXX4E9
3NLxxsHdYWJmzjpqfs4VBsmdKuFe2kNojOAFo3OkCuN5TYjZkFGvd4qqlkbudGlDep5m7tKbLM8S
0ICtFCKdfwdGif5ND/6XNStZW8WiQXT5waXZy0FYHE2gxRFDHD+vlmmTde+9bu0WKT5fVjZBxff0
HWpMCZqs9wEgeHF7ttqepqKdF0HW7cFEYzm4l0bTUmYm37VwqoNVkKg7QF1g58e50lRk4tz1tAQ0
a7sib2BZRdSgxhiD9ksO8Jtk0JdMNT3lVA+B2LBQXADlxcWj3Fji97dTeDXULvsaeoyEkfdWR6Er
Lo69J6UuiI9YKdMzs9peHREF9FN9UdBUzr9hUgxFaSbiJbudzjjqmVXjbu0Z5nKe5+yuPyqWkKhZ
Ko/FHpJeL+4KkufMUgpr5YJjMvhpp1wM0lpZPRLqKqxFvvnR8/hKLNDL+2ee4z3+iNnVsyzoDmr+
0tTs8h9qZFgXr73l7Yq9RtY3eiDVQW3m7OKSUh6qiOnGNPjFFoMq4URyDoqj4QqBWBc1t9gPeCPl
Xr7S3JJrsmWtbgeyvKHSYAHjgQbf571QWu07hFd9lMyUQHUaZYM+hYgZEExa9KDwzXXwyvlbjk7R
aK55cvm6OgHIC+Xdc/uvyt5XSHCvN+c5nMAI5rCWqttVeombnDf6dIzaadT2Ro4MLbyGzc6wwEYU
McoTLupRrgxhPRB+HyNHn/M9ZM97ljQbiNitzaO5N5Cpd5Ur8A5Zfm1IiuOuZywhJxHMxlM0ANfo
jFENOKcxCoObVT8vv34LCnCIf1xcC17oPl6k9vHTxMPjUevrIqGhka2EJKUD8KAHJo8p5N9bFwSu
DiU0Bs1F55SDOQKQZpoxNj6xRdha0tOkNUiDWGmhxDtP64qT/6Km6TuG11VCDjQMI1IEqMSw0g+q
5UmRkwRcIFRYRR8PjKZGQntDeTD40U01+SZ9TiH03XHfgWZju2lCpej7GcUhOKUynbkAG705Qzu8
z62alGu7kRuZkCPBz1WLFdu0DXnPzurD7RuU0dsnJoHbaxBg/yUvvPhGywOqCB7Y7CQzG0Ormbev
61lSVVEvTGgK6aKT6yA/3zNgVcMqZowA+r+nk6VE9nUQgzTJkuJxfIqm+RcQ+gMd1SSNLvAYHzSW
HrM2nDRU/NJAG/Jtlf5Ut+bsR5NszQr2gR5fngHhcv9GsYG3N5XPbxWupLPvZI6albXB4UTdu6uB
fpQ9OPcoQOXOtwTHqcGaGcKsbylPeczUemYXMygfdIVrB9A4wJpYDL8KIU+/3163Y2Ue7PUW/f2o
Xta+gcrKhNgy2e/VQFu8YXMeuQBgOEFQxxcIMXjswYAV/E9eP3KdNQnKJU9LQ/v4E/n4uvmkcUvz
EJPvoFf/qqHQmppA9XNa0MWVrt0dC/lAmlBWsoe7+/elW9OxKYLPc+3s77xxcOOWATwIFwxdRXqt
W8J6+GJsZWPKIOjbxY2pbNuEcWMtDVnrhbATLjwAyPTV1TIxUi2R0jmQ6Py7P0iedgCcW+j7Vile
vH6OjIxrw6uhY8mmbHuh1ZzEqaMOg5pgSxfblpzmH2D5zPcEy/parRUGAhHCuUjJXq0ACHExoGsX
9RvRKmcLdh4Vy9GifmnQ+PjaxTmaUW/V2O5lm7B/kbrLG+wqeJgYavX7ObDIhfFZSywqKxyj7Gtb
7ZtNRcMOLUuRXzNQSOuCcmXyTLbLMQqnMo2LdwD6J39b2+PBgxLutbMPsCVdlU77bptb8ExmBXDA
SbVRe9CG9alRlG9SjslfVdh/a8U7Fs25/zVSOpvfzmLbL315odvhfoHGeRWReZmqNpucJoeyajIw
SgCbQXFOUqwjVCSa1DmekOPvf9xFZH6xZ4okhU7l5luSBsdYtRbC+gaZTJ79b4S77mHU/kVU8Pr1
urYFuj/RldY/p/BfwsTWwREyoEtdW33WIKnuxvRE4Q8LM+H2iLpXncHzxkPh7I6Ci11eUGJaMRsj
8cZAhpINYMvCMTEPqu5qtPFG3M4XNVje8XzhhSi/2uRyZ1Pk3TnEnWKrkBec60v6AHF09ZTU5+rD
91sDj6p6wATDbGdKq/FYGtff1AQSl2ujkv1r7xHm9rwg4ny4yeNdinAQIF/TlQyg/5pfobRP3Dic
3cp0m0X52XUyFpPP39nec8IFc1x2hxu6oNsrXVL/9A/+hYxv2n2ywO1U7yq4b0KJFmz9BU5tf4D+
FTD/i5X0CYhL9Y3B1++0wb0Zhwt7Hp6rb6Q5YPO5spye9Elag5+za8BptxwbvLGzQg/WD/Z8Oc2A
fFrtNUBiDMtCVefhN4i7vzY3vloTOI6dweynJojGAOmt46bpY1/RmrxvTIwUoYcttbiGXq0CjNKg
EmGjh/1Hvi6YQCEgt9Z2W0uAKig+IMIUsbQ29tixKy2T6IS48DY0lfVRBoFARZvjFartetGosmIg
h6wKhEAKVcoWKopb0xR9ULEVd+h7isFSVdh9lMaz7CTct0wEE7rdbm1j6gEsvlnf3kTpvlZjKmda
9qfVegWx3uPWhMcb4RdoCEFJMa0IHb3XZbeXmhUFqXFjyzQ1dNUl+zKJY1dPrpPvR+5WYi1Qdngy
bw2WDO2VjgpwVnfqdpQgwW8+f2B90KSvjgaTvhLq59GqiXcndv//aCqOA7HJFJYNfUqxcYyVFgDv
RZmR1/Ue8DZejDNjDrl1krKCwMoQNzIpmq/LFDFGDDry4MNBYpU4+uibqhG2zagL6kZdydkq1KIn
G0cuAyO4NiDnEdyvGidb4Zn3bpvYHrMDHhdaxfAKQDfew2intwwUw3BOQZq5wUi9mnlQuf1f4mo+
h92QVV3+Xe540YbX8g0a/hwCsq/wUeoLV9NEKBTL/F28uQzS55eRwVRjvV5vkCKurgCk7Rq2fT9l
6G4MHNQt7f5TlqjqqJqZ9OKeUz0sowg7Ax2mlQ5zX5TG6+qzzF7tce80/QAlpz2yVMcJQ3J5gFA+
6qHvnA3T5Oz9QCK0lpkbVmDHvsClLJkf8mCHypMvrb3brxi8qkPD61Z9pFWMeiEydtVEJDdeu7X+
VGR+cvxwsTruW+eKxQ+NysxhucZbW0FMnPrYA5c3sprHUFtuYWr5b2FZRm/U1HEXZzkGiEUoomjI
TMslBVFQ+dHZ722epYgJ3IFjvQgPgGtCQDDvNhl25Tp3NbUU/f9/8woPOZ6H8UsNuRORq2z8rzkw
X4+tuQnmm4+9KxIbW/BoE572VtsAF6EDQPViDiGNhjECBWuE+k3NzxRDiQN1gM+7lKzyRjwTFnA5
IMnk7v6BZJH/K75YtAcSlIJ6ssEMkIV4yd2U3n8zB3df24oRx2B1aYtH35ACEsLMV7nF8LO64ysf
HZmJLB8VaD1e/zRjyUM/noV6wM/vMLWid6IA5uUH7Zn9JBC2GSijJKKAItZAk/7QdPyfOkJ40jTE
iAVlDEDh8lO0JM/JzWzP3cvyYLhRmGaWRfvfn1+JLNY/xrSaQkPZ7oRuuIQ/XPbnR/6E4qr5AKmw
uj+9DuaixQLIJ3Ax9CTnwC+Aj2z+uWHdKUsUTZbpDjTiv3qJ2e9wRKq61rruSFLYWn4u5l79Thr9
hUFebitBRDXycpOFzR7SA8NFCG/CqQdVGEzlwGSspESczNwrja0EJ6G/wUiA+uqEsGiWEezdiasq
sW53EquUMBe3ooBUcmSp6u2wb8FAk81w5iqhPoW6D+OEQtad/CmfJG4Qd8oT2/Q+S+0Z3JoGQUz1
svqqtKFqFVHFLcYstHUqofbzdwC3/aXdHisBYFarjo+k/AS7CAorWBgnk8aALyTeuWnQhVafT+sA
CTeQfaqcIvyzpgrdvkwBMOBpnI1b6bBcJQu7dorPNxuQobflf43cpiUBjT/D14n/36Pl0hcK7i03
vttwj3cY882FXDBjMUBHVaXj1B961y2xTD/IS5oHBipuKnsZsSfjsfROeK32jPR3mlV3sd6qH3Pf
ObtrB7lJHZsgyhx3AZ719eU4BSehP2+NVHcclXAsiLjtRnF4a2fAS9TzNQtbsTejDBkbENZKPaxs
nQzV3C39oM4O11k1oQBRwzzHDmFzE+y4xV+DfXPx+D1qlOJFflnaLFdgdcW7LaM0WdQZu+8dHF5b
vWmSLzROalLSDHRAUD+7w4W7i0W3ehuLqi82ciIQMoV8KPTiE8C5m4QfplvXpXQUpqkixYTTY1yP
22xNazO9FrA+eA4u857o4KWqn4ETRXrmlUF59TiaQSBJYsO3pc9xALijbluZnzrunHbSI7YHEq1J
XVzVj65AVQIxlExf5K5FjZT9y8loHvaBOlWiTCKsCdNtvRAcI6wi9wrOoDMqWi+DWA1NMP4Hhqry
TNjxUOQ5ip/NbXLrObCFj/0r6Ep7EwdtJt1QBz9kSP80GR/qRlRLoe2UnscsLt0Gj7pdpVXggT1e
XaEn0/56tt63wSAECyc07djqDQPlULruGFF2/5zvUibi1WvESQ5Ad/M78LGKJSeC1iJ26PwLFlUp
0nm3oxyWObS1LLkWyJ9hPsP9Z2G+sXlxy0XITbxmkDMwbSFju8JjxD7FAptXX+yugl4cZZe/0shA
pCXzG/GE9R8cw/yb2lnji85zS+1SZB3w6Vd7Udx6bVyMn8czKTbo0OEnBtQmc5Gd8J3gSSD3cWSx
ttyg2uU7RtkIPbkFRD0lvxFv/jHYAtJZGj14m1ekIViGxmOSy7NoTyYS4oT49N61eB3B9/wrvBa2
wPlB1Wr5YfD3xSyqFoWoNqJyiwaqoVBjyyUa1vkhAeIFcJlnv83fE1dthKIHwuxidwMOeP9gpXd8
V3vdcVutBLOTFT5zAVmur5GqpHfHxjp0bqQM4zd7vujJ3K1E3VdBGlbaH1BpVkvzl4CwhLlOi1JL
PaAIV5BZ3zi/LA3oeplmeZTov2UEn4WNhjiwjcNk6Y7n/kPg971JCPyXgGS/Asuc/BJQfGtRF5WA
viyk1lePBul/SMafCwZax99UTLquz1kqptIlX/dp/KNn25vRoyAE4n+WgZYFztCugeXjMhukeMD0
O21bfFpKABneVhI3X/9ZdUPAIcFKwcZS4MQnAAAm6LfMejYh65F+7FIWp5sAE0ZbOFIkZLBlE5Pm
mJVK4yvHnEXyfOJNjniSix+mm9z9ii+DfjE0PIrEWDUKrQIK7z0sq1fSspzkm08TIv4u2Hjm2J+m
OzbiOwmiT9UkQuTOjQDjgGurhNYorIUv4Nq3kjrm6Rj0t6gmiPZP/hKBPe3alvLGK5WJL/EWrxrG
3K9YnGRjQaxWPpp3/UmuRf9VyZWO04c1JY+SihMUQuJIwLm0T9S7hWZ+QOrqmV+INwN/bY2g22Ab
p355A0sf1s5WUSIHIGI08MTfdrUVz+Qg+AXTcnsinQFgEw8dpIWSYrW15FyxWhIzgcKHIua/9OWA
M0ibNJfUMpTPVb+HsUWnzKU525eCISJiU2x9NELMvlDNp1mLUbwUJO1Rs1BrSpmKfrIDYmgBUli+
Q/ajyb6DLF92piy40/YBOpFnzO3t+ZqfvOuIbziOkvgeNvfFJrusEHkAyvYR58SKkR1FoJbiVrDM
F5svhAq/+VDGYQS+XT+xluUPrkKPsNw+hxkoCSclhZVWxa35jhKSVnKJ56jw/euoMIxCk4Fzp6mg
PJz6R/wtU98U208gnDQexVvgh9MOTL934ljrU3saIOGd+igGfsJvAXHBMypQ6alk7L+c+l12Dyui
DlmvLF3y+rCibFi88AoFt6Y/GTM/KqaunWlvV2YJABiox7Wd849QVcyW2wl+BpjG/py72ySbbCCT
JTbFhxkZG2wSiZT14NYAt1dZG490KBlZEsxAlB+/LoWadFMUNpnOU/RTqSQQFjvm2dgmVE8gmpN4
OOhngHSj0IDWn/Ov2m+KYW0pH+VK3M1RHuf3hogkHf+QthyJPjldW/fC9aV5QYuTylTK+ObADua3
wEG4N2KIZpWo1FuCYroIjlycEgEn6EQ+mekz/wemUiMgtyf5Ie6UqODElmPPY5N5YtLaEdfLziAa
Ri6/Vo6Yu14AhmbuJDiHuTApctN9Qbea0N+txTqtfUv9/ieMtXqu8qJL+AzZAlvjSBnlS5tr/OJF
tbYpaGX16gUj1lT3vRjwdejkfIwvv4DmuFS4ox7ztt5d3WmVJcCrTpxcs0sZjTW/K00oKDuL86rG
evITYZvt0bz7xTeKh4l3UbFSfsRT0Sg4+LyU/e1h1U2zkBCoigC7+3mdOVHoQJPCsuwN7YXIft5b
wMlZ93EbUssLHgnSHJXMlN8QJJdmBBGAiBsgPBDDPg2orcL7Bu+YHUCkv+gMn4I29jpHsT26m/53
tajPlLdwcyBGnE3yEXMPH5a7nPn44iP4x91/L/WdAnkMP8nrgKWbJYETS6oMQiazTH9LSEH1nF+u
WICrQSWLhOCuILiMSQiOH87p7CozDQX2nzw45M9DsCQo3urVyXllKKIj+bXnl3dCZ0q0H9l+2BY3
4GFVBynu/D53eCl5LE+ZauN5wL4uUPHu4fMxTh7wvtU4Axqk2LN2KVWZqw02jTPMS/Pumw3egpOK
cmpZW/Nenxq8OQUk61qbNMRoS9vAhyeVk68KLZSTgcr9OYBEnRZM3NvNw0pBd+HTfPsAwy9Hem/E
yQ45S0YIl/3DhLrGxtNNH2mXOw09qnvvVYJLNIBQhp2i/hNp3gpjfpdoJ6x4+BcU6/2r5dQ062fg
muMR4PFQASx2A41bEKHD8l81oF5D6IZdV5rr9T87DRISjCBmxw8ABkxd1DaNMfG/lUvallbR100e
kLx1vtzBW3pOBxDBtznPXsi1VXgEkLZP75GEWu6HTXmNZncpwVz2Dy8WOhklmeXePx7oLhxCu0EA
Sha1P93chheUmHZZWAulofR6YU3KVD7shL4fcbItPJopY9PkpjGqnjdqn3D3ZuV3xBkuo0T5vSaV
/cfLe7v/h1FbwYV/akF/bblEoNlanVTUfvHSXEwxGXbZDCVuToJ7/HJXiqkCJRt0wZEkD3RVOv7g
lbNDfx2L3NxsHKrbAVAKxx43MNAzZKqioAolpTG0C2dW7mfnq9xiNcBRgY1vI+5sYoMFkv6jNRiB
tkCtr8hhg29Yw3bRORnM8AJJZw2AchLUpA2FX09jLWVMT3fx7I99F/wyc9ItCdCqFpS+GpXiLx79
ctN5u4ewEXWyjdo7GZdBlrADMCFZy4nKrZl+UCP9wutswZSRkv2O+kimtpQ2bYT9Uvr1Y6zQ2LJU
VfzlScx+z/kFf2ZnF/Te+6oohy/3H+p54PNVRrEt0Pn1XUs4l+fNv3OgGuMELhyYLtARgxWthWrp
7G2BPEqqzjzc8eaQKe+i6dhjvmdrCkg+MQBJERw9XsE/rMRRgv3CnuO4imHP13wppjp7t8j1TrC5
VROzqhR7/+V/hAmDOj1VhpG7xUptcFhjwDz6T4U0BMHwWHBJSNUHnkpOSw67MYYITAV1WWzC+HAZ
W78nsprL+EWLSnPsuudHhdKPsnBOrz5WWHmQ27021q59HTAxrFfPJ9kwUoHCayPdoaPraYMzaLbV
+1foyLcGrXwGQ7M1J8W3Sd5MdN4Se9RPQcfr1Mc4rnMZhjx6kmCMHvQD4CzJFPqxbPdCR3PeX8A9
9ri8b0AZCKjAKOOnui8DfUJ7q1sG3ThNDgRy6N5zyPrdYz3TY/rFQhXovEoA/NoNFH5+z1Ynwn4G
j8bpePD2pbYMJWIGys0mUu5WRCYVBqHOAfoOsaSmzAOlj5rqXnEMKTac4ISm4bOw/JByLsnwPt23
GyKD7JD6Lhgb63tB/k/3ZM8zFI4kyeSwQU2l/uD42WQQ7VcFdNxGeicR5ueqzZh27xWTb48OWrD8
/XCdsRWtWEfvENBwPTmZADm1nvjzKh7Tx5RcVJsbqRZJSKRU2x7nNy0A6uZfHKk1jrsVNk3jRTwX
3MPaB//NronI5eXWUrPfbjOEHSZI4GAIbjNg5HV0GXz6MXZj2cGTR40wnGWw6wCBLJlmMRXen2uE
JVl/13TJ4JOvbR8/XRmDeJ8CiTcPyum9GCxkaPtLlK7kI5/YqvvLv1isaeqJ1T0YntY6QanEMF6F
EpwSZS5lhMk/jZfJDxE7mMw6xr5BfdmIzdi0c+8s2MEul2cWDQi5b/34fn6f2HceL1mt5PN9ihc3
9qPmx888KjBuEfQAj3Xm2/AutZde54fYm3k4BxpgDUFnn5TxSaHIjQ72u31CuXrfKWY51ud0kGPW
Aaf4GGHRREY161Ab03Sz+gk1caT/XcbgdhjsFhc5UXz8p58FTZncaSSxX5RYhiIgudTcvodq11hO
qAj1mjWBxHrLNVB7EETuDvU6fmdZDJXzaGdVkLmyGl9eRjuUpAn9t/YNTCv/f4CLcb69sVo57Y2l
nNjJPV9/e+Ly8LLRQPw3nq2hgxrYfcLXb64PkQrWXKM8bLTXPicCo8Jvhg4ny05iXDFmsAuPSYia
MqD1GHQ38qF/yECyHPxP/WtjaDXL5Kva7HBQpmTIjta8yzkrHBu7jU0iaTiVtbemYnKAt2lHwcYZ
ghS/v/P1qGcytFM/y0IsyFPN2jowEu34+8s9Nu9vQnIF5uLPbzrivcUmjS0sIkjxI4t7SVE03W5V
TMKer4O3LBRDYqJmmQ5jVdc2pXDPw0mJijEMgNVS352gRQRdjhmrIT+T6k/gHwiTR2u0GKGZv221
Qvl9iCAcL0YpcaQfOYi5enHiPTCgDWfnsFs8iHTaSq2cWFoCsiQ/xM+hyXsar94OcCisvxMRQ4Ki
LVBz9Z8TwHr0ZM1QhrEU0Srd6RYB+m/KBqOCFYtMBeCMw+3SHnrc9YjVNSK4enqCbA0LOJ6I5JAE
NohMEAxy4/NaU+zRwR+vmW6TlVnAqZTphECF82yfw/vHhuaEUIXBGHrKziv/4Vv/HQLx72d7JxfG
u2/MV7NCJ1Kije3hgVA8xuGPjdoV06J0jxtKteM5lokdZisJ1AKlfTSfzhHqfD7mJjlvWmEXmWO+
/8hb7/hPMjaG010oj56HGo0u/EZ7FwHS6raa8LAsn+xfMwBYDJylFzIJ/iDRgu5sIRH1lYBYpvE0
pAy03iKVTmAocupl8wi5W4ZpgssordzwJIqnZXeZIilwq2bOKFk4qTc5Wq/EEZP3fJItyfLgT8bF
6r4B8LiBCTgDsw7BUVweUzEUE4ZNrocWuyGqsjZkv3h8MCHFjNjAEV60lzYH7JgFsTWEaYoDos3D
NJmZazgGgAsrGOTVINt0yFBcEY/LSZ1I3DGS7SBNyhLrw6incGYe5R4s08NWDmzTT2qJEcoH+5xQ
Xk9ZtYO8SQkVEmJ28IEoL00fdx3LsrdeYF+ecbvzwPEDgZEAzJg1rellzjQ5kO7XOu7KJt+VB6gp
nQvWDPnumopFm8b7KgowryLGlUMiZuXMHrXAfauhN6l6XPt8g6ng5dxWulNsn8FrIjVZDgCbjYQL
hVyEH7JzvAhtq+sAhru8hilYL5SYQldfVsTYlfyv3Jb3Jfr5WtL2FiN2xS2t+Dn6efPyZM3JFINS
d9HezouParylA0vbUX5lycVGtGLojifxDHW+RsWWP8IUPmLct6WsSjjScm52VF9wA8Bh5kTG8gwV
UQKRkA0O1ywXgzuOa91XI8gztudBjEYYSDf40ZXwya1fUdow8QUHraKO68Yq/5LPQwzMtVwObKaV
x0JTk0iMd0fP1PJ8s08eqhek/emlcNQLLhwN3fpyHFLQoaU1Asn3J6MKiL2WZg+RQkhFVrv4dFm/
r2UJZkCq1lXqOZ8MkuPpRJfMgwjvy3tLJW+39jkMhHhP7KYoojRC52q9fLuHdAkoIclpIUMLxnCg
mOe/tWce+/G6eJwSRAxouPcl8frsuKrta+KwO6rYtYqQgtFRbAxrx1yne4OCjqPIUDcXmj81rmQ3
dY2HAAMaP9DDpU6/sHmkLnH88+xCRXexFxkQBtzQrhf/Ghdw9tRj0D1C9VBDTs2JthuJXD+2s/a2
l4tyAa/CABo3Zxd9a7cyrrwUCfeBfpLG8tD2aK0M2gToO+1etsP+2rvnitWCh6SZsR+YLslc+Pdz
ctKEyYuBraozPRcV7BMmGhcrmp8rypjOFulqhAtOLRijVWNSJrGm2vMoKZmougUu/bQUAdhPyfrq
nftel0T+S8BpROkNRpYEfLdH7hSVOW73G9Q5hL7oysRiGHPQOs6PcLGg7Vq5bO6tFwMN0MObZl6E
8PU1O/T0JwF1T7KsqMrxWZqfb5KuLvZEsg8T0pi82itpgeZxetyh/cK7DV13qPOf2IECqPsRj9P3
OSIkcY9hmWpp1fGbkoIbJ/WYkqA10LFai+I1HH8QraamGF7KkFi2+FOLP2mfYIFWQ1wqWFkIEJ3k
iU7uWhfQrHooRRPyw7yVDXanbGs6c4ChAmqwXHoJ6pSaV8lWUTgy9VzLmU53iy+od57sc0cpyHp9
R8Uiw9e4h7xweczqMJd4f4qb99JIoVXZjEbhng4+r0s6T+As3tBuGGNv2TFzgTdmBcz2WDRxuMUB
yj7xhAcqT0cd52PQpLUgJGhrYfPWMTGRj9lYbzYSpsfPYeGeKw9Ve/sDSlaYdG+BpmEhFakaNbem
yW2UaAksF4u5YRQI4WX72NnEcEixyIUV49EJfEY0x47pWap1Iu0EnQXNSQYEdSjYYgn2SpZCKmuu
73N0hYzxjO9VTyAEwy68thTrXRoHa1GTndjwkTSld7zL9/z5fqTcssgf9ZapciRqRhtEgLSRIv6B
gWmd+Xijzdt96rZwcGy5Fk0sVidY0AwjKHxPIe8x/9+7/gGZFxuRHPvTUU526dRn1mH6MYKj2UQ/
vvX1SbiEAGxmgW2utcgKd1wyyObe2xpESoTaywXEaZlrCiaThJ4EKJvrPqa97Q0DpPalXsHJyVvB
hqaJLua94ybX6lCm5IZl/jPjBH58SsHE1h1umrV8bflV4adtjROTVh+yBgcHmDJqQ7dTQ5IeceAR
OVCiwHEs9BAzQv3dsll1J+2j9cLA71gGEFrUzsgvb/WbQWwM7L22mgZQ5ZV9m0uluSsD7fI/czxb
xmJ1D1lfOZgC5VY47a6cs30tr7/HaecIuzvfjMtkOC+0PsRvFvra4SRXgEKRWekVGlRV456a/VRp
vvrWv3AL0cHCAhcxB92/MuSGdbrpl8ASmwpw2vcQVj5IxasoCdxUrFcosXkdMk+tmk8oOw0avN7x
Esg0yBYpJ/RDS1dBXc7IWL4FBWvp7wbM6MP3Jopfk/TFmEY9+/xTDRGDQ2olE/bTkmWnRXYhfM4p
CILqWd/v6oWokYE4Mh6GGSiDyH9tJWbMgPL4f1L37ldHhPi2Ghne0SgKqkO00MYVAGceRYdv6G5J
kSiyFQMow0dlwlph4tyEwDvOhvjerIFieHCntiz7wX/nrVr8lFPkoYU7koxGpEsDWYcc2S3IhI5w
n3ZrPWmAj0j+ghchKXRO1GF5A5jUhyebC4PNeEc1NKFknozpkS7a1m/fwqOi1PnD4YOx/uQd2MvD
0ElsCgFS38QM6zpigUEVNA8lcq42F7Wrkac/xbjLztT310yHKEdf1n6chalHMAJOOmGJyHZl2lbl
CL5oCMgqOnYaflHv6Z4SwEaYheofZ89dWM3pN3CoX9DzdD19Zre4beTCP4yyeDH5lsiuIOpcst4/
6kuUBx6h3Wvc2UZxf+SJ71GkNEBsqqRTBGKM1IKTzR+UTkOwMPFUIYuo2YV7w3gmHI7NkC7MGfzw
3Yl7YTxptW344afbBhP1hSfrEj1Sgr/+DXjy+2xhNA3/LrfsPW7zFbLLBRAlFN53wcThCG+Ft5Am
y4nNEKKmFJ71zeXj49DqIaW9tzVg9muGT1ztmajskgmdo0kpeZrP6UtfNGIHP4F58gKjOf+w3lWU
b1ZR5dNtOj2QzP6GB/ePv4Ak3MmAEmuvp2DeofeNKMT7gi5/m90xerMJhxa5LSxLxa81rtK6p+pD
HPBj7od8bfV/blctTbPz+YY2wQxVthNGtya2of2TeycFia75z4umWoMYU80BiA17dLiHCrwPU50f
9G8XxZNHUR9wxfuyJDBcj/t2cNUa/fOwLP9oi6GlmyzmT7BTIv+EL6fjmHihIPidE4GYxJrtxirz
CN5Sj/t7+v1ohh9mMbtNq5W4oju3Yvm/jBQOKoQdHbAOu76EP1iUh6j8+HpEdmNHztTLquM2ZFaH
umrntSgUJJdEoYCDG2DJ/apEMkfCm7vhWIRaPEO2PzwuJqjIzQtqVSQ9iqOZOh59dLvjxMypp24u
DarBlGRfAaSEpaH/d7f7ZKhNrMUGoP6WQ2aI08eswd9OKnqvm6n10gKdQAG++5EJALj+mDGY+rbC
zrycCkMgqbOWjgGDil4vsDBDLxjsalsLxuCqNgvrwibLcY+GRaecGAnTD9bDUAP5kuhqzAP5yHND
TfFo+JjkZvEsJ19o3vL7mNEJqTspoD2yBIJ1Ff3oTqDwGwx0UiU+Ks2k5+OHJWjTjzgj/8CAWSQ/
AB7hThvj9JUSYX0F9m9mboplvVMVIgQ7LVIpw8Rxv1DJAhHgi/ZhaG5ySGHXIwNZemv68DJ8LJQf
yW/rZeHRKsYyXBu6upEgopjj1hZp/YxsHR7ypy8d8xUJR1nq5IqBDmZeRHdZPjfkOGreZ1WHCa5K
PlUC9LSwtXpyz0KcwlYWk1Hh/+Je2yyMN3kYY5mHR5rI8WEkfty+z9xI2/nWh5MtK6R7CVb1cER/
5/4VepFXU1XI1Im8J1JDqJ92Nsj/AgxQ+wYI6gM2O7Wfddcdp/Zf113E+e9d05m6xlVuZ5OxNU82
P7NxqWO6LYSkHQGjM5pmBxrOpQ1qEFIrU6i27Ee83tSqapEQQuhIi4Yz1Xgwjmkza1D1KDgNsA1a
h19h5mt5Ho3WdYKfwaaHkhMWrujVZW8peId1ZmNQZUbdyR9d2qRtd/E0hCJYaaSv1wMhoqP/yw3D
5i07SaOvR33DOYqvUQ9/VLbFoa+PCDIXHCQ/RL/sfoci5E6g2dwr2AJTfY1rDykM9UZnap9ZsZdn
qNxOEzWSDB0NVVYCxE2UCCarFzc1tzeVzxkRQIVXWoYood7G4IeF/BytLzEDamD4cVMBx+Da/g65
gMHYAUvwNAVYZcz9Md536fM8Bt+lo/nSqxIu+YP9ZCfXZabLyVKeaeXWaPm1ASqei5JPQGxrIP8o
iGfmYEAuLRvSU4PVWOpgAUzHsKetW9Wv0DFKd0of6FIBrYfwI2fckPEHAKCwYCtflMu3bMwUlUdr
v609En9EcQQd3PmMQMdm/X29JP3YSW+buNEfEFde0OEbpM3ntg/AYBIh0DA/0LrsF5xpOJ3dg2aP
cRtqrfto8b8j+mpUXMTDk9RcX76uknDlAJO11zDzC+xQlYkooksug4C1NqEQs3ff9neGJJ8iww8D
m5FYAaXHOvC3eoV2gezY/vMf19HoIsNYiG47fv/H4nLE+k35zhzD2ObqWMKt9b5gODYCmpv61N4U
rxRSfOGU3fyzpX9/GCzHOXuMiqf1lc3wFV0JY65x51z9/G5HnuA5tChx5nmv+AmwFakozbl4u6xP
aztI9QoINwWbQUXlOhkf+k+KT6sVxB6JV+x7zbZNldVLLiSoq0DgYBqNQTUijG4AU2S/8ctX5n16
P/CjH57vufWEifYEJMppw5zhZd1MiEDncKS9ajrh+UUgxlYQrRl3ulBUVFZ7aS8jUQaUzhtRV29k
A2lZHwrLy/QxnqPkYJZZriAW822mJsQnpdJYIbCdwoOSW3CLiPucwEN+T67m40BIqs9rmKluNwjW
EZ6B9MyuEbWPFJPkPEZeks1baHwa88nQyAI15cehY3It9N0x5M/ZRT3S3W/BFnnh+v8EuJ5M5abq
135jOyiDnA8qOJvH8nFDdTnFAs4XpIfT3+KozerwYjzAEXf4a85fKLHtYOscf0m2PfU6EAkdWjKj
/cYeVhAp+jdB4KWOJDqAZsd8V8/Li4He7z2H6N72nqJWL/0oXaJmrdjO2SdLKayOI3aqw7CFR2NP
rBT4L2IkFbrzuHch+eqsvTkDrfym9nHt6a9TjTsDP5PkLXVHRzsViNCpLnKkR4NtHcU7stm9SmOg
sOD82R6VRa7LM4XjZKovMa2IXh21JvJ3hXKGnmSs1QRT2oZvvH5BtQjRu3qqo5yFuMihlCzSWBxj
YnnFak5bZ3JnWAv0d78gMVLBzTvkNn2pvQgTKZvGh0pER+WtfuJ0yY7km7zblcFkLCLjqjAbsE+r
Z3gExCB2JupXIHdrdPoIhtraKLvJJ7jZNf2hJH29Tz03401j7cfn4RW/Fs1ZSICIK7zwZexchq+V
77Y86b/qRjh859rzhbuvu1Wk2xyzsHWYtLJ2r9cpc82Ss/w1dOK+neWGZGxpRygMvKieUYozpA2x
a/JDTmsyNmTN07WcFJY7XcqpKsJVXnV4zDKquCkS0WcH8eDVH3yBio7Q4IA4451Pda7c6Gfz0E01
YpjdUTFWhwh2yTCRMHsZ4OUKk9F0KXqMgR/D/sYdxrQWdr75rYWwVHJQ2DWOAxuQK0yPnqV/s+jj
EjZKgpg6koOiyKzSWRcT7ZbjHs1C4/TWyTZmSu+RH/4Vb9pMjrIX7aFhFFQQmo3YzAi2wFoFz8wb
Es+hQv4KpZ3RBN6icJTh64J9rt9TJatO5vV7rQpwNewxNhpt3oLrNgzXhGJAbJK5IAWw1QHH0jVd
pQzBbyU5HR5ZIdfsI+jZy1eij6pQbDNQ3p9DGynZquqAZ4upMvH40kmR1+cXL9/6KnK1VIwGAfeX
sCmPHeCwx+fO2I3TQiZYz+VdzaaUatPJWQQfpvR/dP/Ug/ISMpSOa9AFBgY7KxeEGBmM2muItkA0
C6p2Sa7AbL1ySnNjPGQX3Y9isi7VJqF9kmqm8zyw6llMz4+Uirtw79sJ446sZNyEd015lEI/RT8o
AsvVkOCvbItjMAjc5KaPGPw8/S0IUqjkgibnd14CB8uEkH+W19GsX4K4XpU/hb/8Nas+ldjXYi1Y
Zx6IiJ0VhCuGjfJawsBETJvH/PNzFfAM94rGarTapNQv8KGP7U9n3ipGF8P+ZfqJc61UNBfZlMKx
ursSE1G2H+GXazAWjwrbhAdUEl2Eye1Ek/TQkHkO0owALsI0Ltt7caC52wVxrDxcnBqPL8O2TzDw
zEPqE3lNCqPQmiSrLacLzDCxzFRh5gPmDis3iDXgYDg6U/a8OJvrgAYBnGoLUO+ZBGcNo4e80WJt
nkXbYT7hmHwMCg75Jjhcfm9mkjTRfP0UbwHBdmlELBSsytC2Xt895jOJd+C1K5etHkX5MlO/jjQ5
EZhTIMgrJqqtXzUYdm2Djz3Kog9oGEgUXsZVF3EepDm9ZFxMQwjgcRw8JfzpBTbiBtKsFCdITFw/
m1bvAKpT7pACq9KihsHzZjCdsJCIviYSNXi8CtkjmrZtQOHh9gZVxzrrLRzHLSu0JSbBesxl+Q5M
59A8pHnfFwnrr30g8tuGQz7s+g8RhX4EkvPCCWLZeQRGICfcOzzyQbTFqjeH3NILmduJ7uIPpJrY
T349NWWeE2gaN1yAskk7Qd6ELeiSDaYnyNnDJpC4U0QtGzQqYqD2I+bQDq4LMskO8M8d4hoCpxpK
O77ZV3LfcSRGLND2no4AdTBqjs9sNaFoZH2YyB/WQqonVt0Pvlmw+17d51ct7HnfgxmBkYvZDwQh
fXaSAR5lX1klXcmeFDAgIDDsY6VG5IAMWsur1/a5vTUxhos5ZIIiCieXvmlVAfm7GHx+e1GjdXZb
km79ZoW+7sEyCnLjCaTBMeG2cHwPoPn0RH8Oio9DlrhtK6d4iZQjvXBJbN2t53zgwddPuuXvFEvC
t2QF9P9jHhzDSslaME9xJj8hiXJXf2f7Z/miU4mkZ4pLa6T1wy0Da76mdoY4+Bl7OLuFNjL0167N
xi2HsylwPGXJtKEy8mupSfQuRcxr6enIloVtJ3ov69YSRcLQkAjgD3fxKMUXhXURw02OTSwk6auo
ITAGbj/5fEY5/0mitppCCjC23p2jy+gCLLqwooIFlyvkEJvBnomP0HrVAX/I9CB0jRLVpDJxKHsV
mYIt1v4WOiY+f6iAvb4EZrtBkOLxPJjUgsvUwJ68o5Hd7lYBaP8KDTkVSULbR+gwieq70q5OHVpB
R/X6HPsKvQ3GWEfOVzemY1bO4D3ULy2yjoJf9jBQtn1+Rb7e990b+pkmQziQRnWgSPEm9QZchbI9
PdEjeBFerHzcMusi8gkGEpQO0Z2PYx3rn07/00PiOJdRg6meJrTUnyvU9pNATaJg7+I6VbJk2ynV
4zgF2JfRS+dSh73IscAmbFB+7dxv+AbO6SPoPKmuzdR3AVKWb4IqNYpWrr9TNrFkweM+2JpmE8uj
bHXx5It0BT32+Vso9DDnVwyxlkyU2drKfEZ9Lwt7bSOOLm2p64e86iDUp9IHIQzI8YIESf3MP3pY
BczU4D+ty5Fw1Yu3fTompAg5GBSKGYjXQNH8oDnlKB5Pnbj6I2njTEJZvd2QEwbk5xc83Bs/dg3u
5uGS3K3on9ez3h7EUfYAybY4PDZ38uAtaVJhv54DBOjVwYdAV4YQMLdy8Qy7Y1EtZap+CuNpQarW
ImFqhP+cO4a5P/oIBD7r7BAiuJ5JWZ7UVbxQ+0J9l7rpYR+Wf0c7NnzQSyhXmrJYt5EhhKhMn5ik
AEaGOiCvqJRFFMH2ZPHmmxrVKHhc+k9ofIHPV/mp67MRjlKzOE2Jd4UJjI1kBPt3tEDsTzq887Gv
Dc49PtXD6lpmIxWo2uYRC99Fm5tt0jU1dt+ze9cesA/CtxvJHRS11EtAddQfApyvE6oFGNGDYYqJ
EnbAPKEtL13eHMAksJjovf2B0x18nhd7u80Ej68rkffgMP5dtTLuP5i4wecWo3WxvMD5Dyl9s47j
6M7yfHRptiWZ/Omh+c3onmC6akFIAPWYmNAxTE3mwbdZWX8uXDyuMcZ6JvwprN5pZLvIdyB3WdR8
YEt8CZZLfZ5cFfIUqDU6E/tyuL/9UpzqMLs/EIgjyPOUcdv7v0iPkqdyFPJaAky/Rwap6G9pZuO2
R96bpnzDM+PdsVFsLT0cDHoa8+jvRXyMP93XJFXg58hyoO5Aqbn4VHQwMiHEDXxZrhtVpGvf4pDR
vvI7GVwUl5gOqXBjb15GIOszBSAlshdXmeibsZRzyAucu3d+NRdUnftogO4aBQrtY1T8ss2/1AeF
yJKulQ1CqwntQ0dOXOzguuAUJ+FsR5HsIllfWC/RAE5o5I7qDk9JTbGik9gfkTuPTb3UOdPylnRM
vQjdijz+L7Wt24f9mHYmUKLQufxzXYxLfaTRqeHwyMS/F8REQhbOGxGJ/AyrHN/cDOt7vgmcNDNH
IHP/8Fy1HyfojsnNH6Dif8EanQgazFTyKrGWXF3qEREVd+SKVd8PrXRGnNUQa22VJp+W9PYsBtti
ujkMGh0V+Cdo1DSbHlyR8Q7BYnJAWDhN2kThIO4OhYrBUB8SEFLNGXcXUJ48y0HmO4wbXMvjqmDM
57OgdxTrEAO8E6fjupUCR7+FbV5E03LlYSoKamVkgj0ICUwlMoDcPXqTd2cuKfErihD0vcevmvvQ
YAiXd+970b6zfJKriwmgPGKJ8DZH1rsDt8WWyAitaIrPOvlbLcV36yN8UER8+y37Mk6QYO7bu5SJ
BaXVR1bYaa9dzOOsu5ef6MsgsLEA4r2e9gyOhL0GL7r3VwWvX/aS53GqAzFUuBzl+vhMout/7DpM
06ZT5fG/+ZRhu4mgq4K0Fhn2+TviiTS+Ex2tRw1GEjTa3+47l2pJo7b2Mm9rxzOVrS4ywBGVhC/e
EDd0rCVMe2RLOyuVOD4RKE2ITqu+yKTfc3byjTOkd87ZV/f9n9fVazvKtdAXvbPMjn8aU6ONslhQ
zhVWLqb3/+AdFZhRqvkvXDYsw/QGgXMfrKsQPUHHFXeaWDQlGWx5y8WPiJazah+Gu9XYm/IwmMOd
oz+ZAGhRfRHKVizNutBbpx43/Kmq4YiiMvvpl7GcTMz7cM0Uuj1ZTNU5729qZy79PPL3hZwROXbt
b5rTu4QjESNM5W4MJXQbea7xrLa3mOiZdM8heFUjRZKApmQqmwn0ApNh81uHTIAySsl9aNceXA8E
QkwmrYaAxZpVhPeborWgGLChnBlpkuqopuwm3yxqtT2Qbxvk51LI98YZoRpLoHFfoJRCzMVd/Mim
kXoSRU4WUEmhbl5SJTPf9PtAlFciLbCVd/HgGItVEO/3SZXaEX3zldTGs8U8bmG9E5ATeroY4W+q
ZWDkWbbbv0ewkg+KtfAHAALCYOOCbLRoLJtB/YlC3qogLWh2K/BruEHLbW+I1pcV6rcSKYnlIbop
mRmAB1Ld35d6B4/ZuJNGNwWJ/izCjWwfw70qsoRvhHkFxzXtWDHaR/5tASNtY9eLYYLBpVnvxQMe
dRZg3UKffDciKOkVcNLSxPbmTFz6fc29lAq7Icat9e/SjuWBy3l0JSOPOG/sr6WDWCMo0VrUxkpR
cOYfeUbmqRQBGSpXSce8aQnGCxzwyJ0BSAJVj0tyOcz7uyVPSMX9J01QbHvyWnK5APN1lf+QkfRC
B+P0I7v9rXHI6adrBn0eHGr3rvXbI0dodAGZBBmEfmo/xeoqfegW+x3WR4rqRH32cnFEV1jDxORh
NkX1e5Ki0V7wHjSbh7m47buHa1ld5dzSv8Zz49e/T934m7AKD0dqPQN3Qy8tRSqv+Z5tbYcTIaOY
JHDqtcMEOjhQ3qFWavRRZMydb/ChrnvVaf6gQMoxm/0PLEZJeGK+mKRh/RudY1PZrIual1Dt2MnF
3P2t6CRS+oU/YjOv5fWFkHV6TbLYpN9+iPa08qXIXPIpDNpeCagryhSKtkix3DERHMZ5FgzN022F
9ggclSMpr0L7tLOXE+INEb3kc9Zub9ZjDuwObjWNIH6LpQoojLfS0rN21CKM54/PcF3g/oUH1uSP
MumjN12HGVECCFhVIHsVn2lGnOG97zTqLWMaAM8xZQeIaMzHD1moxl43s6STexsGAhzFqpXAYf0P
nrqD0FxfC5M54dqyVSfzaLt3EkM+hBDonbfCtB+phIQ0pJDEhhfhOlUrv3uwOGPZyOhkZLK5PN5t
jIgHDsPJB63VU+W0xK7ADU2bvzH+6b3z23AKJ5SWlVhoEsLki44Ndpx0YehZgCKI708RkPHuqI0b
tMV90JWCXd/9PZkZS3tID/Pq+KludO1hQkjuLnnUhNtoQUnPLcgNStMYKzveexOMpTKHs3grbC+J
TQmjPlFIXiXs9INTwLD+eOLiOFYOkFykJC7OnYb6RAPb+mTA0VsjxhU6CTZ80bCvh0Y9NVLVW2XJ
z9nvrrrUM1SfnEFHV9Y0kizkWJboL02VLgV8wcm0s6a1SqEGfsW24i4ExPKyAt1uqDnd+pFoMcSh
mD1yiklRXg58ESFgbq50r78cXcFqf1owc/+sqYRtBd6oWH+yTXHemr5/hf2Qzea95YrjfYO2n6IE
ROwH1dAt0VVNt96yZ04VBLF/Ovbvk8FL2agMiDnhj/2Skze4VlF3hXZpLgaTc3mMKriGr1cxb+z6
VTwwI6sMkfuoK/1/Jlst/4L1Biq7PfsbwrjRvU4G/0FC3vFahc1zgp3F5A4e4db+LhVCz069a/82
YFLZFsPGe0Lh239i0/8aaQsrOxZLKI3vrIXQiwsZ6BHKEbaq531TML9L5yhbMidlmV7UslSoVVBE
inBKcYNX6rP2rFkFnrIt407Z9aTfTwgAs8IzybzqnltalTy65H2pcqk8uG4jEPPC0uPRC90a3mfi
L0k68R93xHtt4WrvVGZ2kWWIWjtXfIFohedI3prHr5+XO11uiVxE6HFS4JhFMleq48oCQ1V5Jk5n
kB3TVUUs20t7l5IvKbxQpz0H+oIDoP3ILguRVphxfJsHW4JG/rwAm9dOf3TTDFqCCxa2SuTa3oqn
74OjVfARAP5WHAEvtQrP3rxJ8Zp9l9kDkMR1drC0EOTjZkUxYImt08dWXQkp1sYZZWqXe+SZ6JxO
KnirBWVbWPvCrm9jCJfk54wRThLYRwhdzMbi+ghVRUsssR6/m2zEg8YYDnqhBhmBaiHUXFgvbwxP
IJnGLYLluTjOZkNvtdZXVJyJhN/+0880ONuU4fyojqpDlnmTowr4nWranECx3pEgayiIlhNfFwuV
e+eVPhY7JgUmaqv6E/Qf0Q58BT8luDn6hZlgZMSJoKpJh3QAVtcex4KK7MNp9cnfLp/saJqp2NPQ
dKJA3LUCs5TQAVnJ3PiEUz2TxmT/zJID65kVTFFkwVNwIYObKKetXKrO/Gpi/1se7LBWoVOYxY2C
mWoH847QAX+8XljhamleF/Ua8hE3am4yT+EOHtpyvr5ittLwPY78kWqBnSIWk3PRg9KGfoiwY66O
+70Fq+z8ujsIESJl2lNWLfyIxzSwd6uIPyooylkBGBQZm/xRRibyms4QhBArWsgrcVoNhotlgeE6
oR19bEEtHqS9L+YHHw95jIvMMF9+H7NtDerF3r8qbz2K54z6T7V+BCgdUCh/WkHCwpYU9xfXZaDZ
eSI9G9JPFHnhGeg/0REhkF+00K1xR75uqUAg4Klj+8XqOBXlFJNsY/zPbPoVarFQwmj/q5wmdQ+R
55ZENGdGRnrWx+vlhU2gBM9AARjuWW2ZoRYVoN6tNMGYqQWKcRpBEsmvJC5QGKdQgEn+t9O+5MZf
4eFADj41/w6Iix01zRGi5DyZpIB9toJ0lB0E49eTHtepjbsQxqHtI6TkMtRN7xPVDOfBAxLmaqL9
1budjwTgUBOuca8Zy+ErDDdYSxQSEB3ICmqMQweVeQqGG6eQeN+v30mFSycLfmD8tS7xI/9XtcDw
tUI3Ku+kmwSvrys87GoUAenvnMNemZog+oPt2I/UPUxWuku1rb2oNBYIRatXUj2chlFx7qljCju5
b940xsNC1FARSIT7G3EoPOOYmYQRwOXlctGYIVE/iDIDcEQ2wyjV66GMW2c/eMxktrIrZx6AljpH
luRkCumvrn/VRsnvzfByyWA2qky5W61mxGyunyBLQfkbQADbyj+kf1TdPjXezJLkPrCdt9PeJvAa
C82JaCcfHye9JdPi1pJ+Jg9/ZzeLT0Isr6ec+ZRWtsfVtgcTKqGf8ZN7HPBUYcKWzj6/MiWpdFET
4R57TAxXnUK4j4oFLhfDPna1Mz8ZMhil/jXsk0KESLfTtCMSYCvz0GUIBIawtU8n/AHRAtqB0JP8
Rms3P9bbi4D95JQ0XHoJ35lLtP8c3uAaSfNFRFqubNZOAuc12uioom7FoYNhmiuqwkYJGfEM6grg
BCV8kmMo1tSnZQWVgDAl/3MQkAhlrsedoQdQBfYf0Z6+8durAis3OZA9SShstyg3yT9ABXoD1I0X
4PGYa0QPujAbePw+bKyE9JK16iu01YRZOl1WU2doi68csdtVt/3NI+ldv84hZKoiwe2d5n2fEtah
tJuUqeqFP1JG05E9//mKA9FW2qEogIu+rc2h91L+2pGHehgXTWeNAgFxlaX+1abFY9sae3SOrlly
GYIPqRw45MHFQ2R3+rhh2haqwC7bIMNBuoopU/1o2ybxe0Dr3oMtfvWemumuGb7foGRNCz+PVPfL
auwbLPZrJi91rS7u7qdQ1Y/kftyBEbRbvLnB3JPeJfdequMRm4LUSadMYgn6NrfAO89+Wx05k4sX
H051J1ferE695T84Cl2rQ3KR8gn5BuBsDPOaLAkASsTcAkEgRUTMBTSsfk8uAKCwT3Bc1DjHe0D8
r7KjOB7QL7IRd6a6s/j/a+orgcF672zjYj+diDqtjzALeHeIXVHUWwBEeL1dO4cQsw/zfzidjU1e
vbz1PQaWvEH8fR4BRAmALIQotYqoG9gxHKfSlE9QKAAfonhN7Dz607lyNwpw2yJGDij96Yfk6TP6
PRn2wyroWpe7PUHJ2mtht5doH9KqL7SGyK1HzSaOwaz2wkdDKNY995/qDPfVbRAdXKLJgiBr59wN
UwFGBdxjMPi5TE0cr0wQr+YzVIAuw9GLfHzL0nGzX0G4XY/Q/SLIFWs9UajbeQ/Ry5ECg2O1W/3x
uCHxfFSVGrCinTk2EwLYOgVObwUkf1CO2K83ou7Z2dNnPtJq3+kgjFRNvm41PhJo0krwBUruUHq6
GHJO3drC3qMeekC8KCT/+u/lLwYe0EZOluSw6vhu3M4w0stXdia32dsC6UhOwM8PzAhYd1FY/zRr
C8gIoSZGWrjeMh7+eBWnGdwNb5z25c1t0uqTvgyoF115et9QnoIgcLb3cKjqNWD7WINEM8vOxOys
L2ZkRwJWCfLWBJRizDy+qCFYGB154XXUWs/8x6pZkd8kGtEqwcX519gjUsYM68hDjY+F3ljshFq8
uItkh61RV2M8Y8g4b6c2HvVms+c3frGaS2WEnpZRCXiuNalmRdAzIPrHE+CbYiDsVowaIYrtnt52
eVYPeICHRQ0BudavvpstLglkPTXVYFolFstsx5z+JmViBZyVavLPkOwrH2zkoPnSdDBW7+mSfyuK
5xURli7GY2s/8m2/TgMXu9Gsayi/+rguWtPYdBMTkUuFi7MHV4GKk9GxhVKkZkMqgjZ8EaLNZ/gA
5/OQOS4/9h3K5X+uwM+IguC2PbJnZht1pzb6rF7TZ+rmRO8wjGpJDUC9moQm+GmRL6nSauz2UKxl
L+nTtMe0bK0PwkOnjWLT3REL8yyqlK4MfpCzjUbxLcsu9Z0ugwO2NeZtY3u19FuegMdD7ckMtYdd
p2KEu6HeKTQREKK1WLiPuptLpNWybpJuMmxVUlD2sZIrIC6hdbjQgl4Yc5kg3/jOCX/sS36xOmrX
No7zxg8D4AIfd50A99jB8cJGhSWV8Dv4IDYU3RqV/4W1Cl8Pst8/0pesXr0noGfefIXfOWi1nLCJ
l5RedwTLNL+OzKxkHzJQDRQcZtXC5/Mvd77XA3/jqWZocauHo/d0JGQaMGJA/8SLXUKicgyl0rkt
E5AMlblg0NPG5EJr0GAl+JXm0Ty0WyeGPYCz5Q6Pbz6jv5eSb6cHnXEz5sYMpyUB4wbWklhka26F
LVBWl8ZD2gX8ccgzqFnkukuQHp8C8mWFsEgmqsqoBVPovSSzFqb1kf4p69ixHkvNL6YPLe4ljZmM
rpTLoFDXgIn5I9/skxI6/vanFcqB7cDZt/bk9Dky1nRdO52ohTuktG10ROMYDZZp2CC8bzNu2wZU
j/VyEqb0DgxDDA3X/830XMdBsmlXGtbvBHR1BXANOl26WIMnsA6E+GayR+ehUv0hQDQEnS0EMvBa
wHKLecaGQLx1joZWPxa5hEhcyd60qzy6+bBp4xyDBKovPrBGp3eW+FgXCPPcJGfFZcc031mOx498
XnK7D1OvVNR2x5lCci80zdjlDDNPfujODcbjjUrTNclTKbBq5b1SD+Q/aR/TlDyPVIKJ1K8KS38f
VdNn+v8eUlK+8TrGC3hvmd2ShIhLs3clwnz/MxH9kvziC188Eeg8nn38aEg3nbvUwVc6sy85QJTi
7sVmIUpv9EinV+L9tp9AP0k3q7GN/fxVnP4x5nOCNZQF2ho0TznvkAJ+FJRSIi2gkBDyPdjQT5qG
6o3dteYSxk2tX+ygI4d/xifMxJ7OCMvjKFFqoPTVeXkY/sKnr3mC0OKKBTjQH9B8nUgpYv9RYPfA
M0qmH80F02wmQEeMUznpx7Ha9XauYm/Uig1c9BGtj9UeBe6GSILCbdV4vzrwOdrAbEv597ZJhWT+
fcWvLzBive/kc3Wgv17BuLgjZA4NUobm/VsZdNTHeBOtV3Ysb/fia0t8neDQ/yeOzdRlLhfbVVbW
Z39eONgWm/YzJayuyUe+WYdi8PWDrYgR8r0hLXa5SBkp95SFnjh86BgJnmnP5ou93E1M9Fuy+vF5
fu7PyqVyM3WX+0lWGOBFVBhNko9hoYOn5HNyUzgSivInXjKVg8u1ZqUDwLoEjhpS0lmPFYxXazgM
oxAq/iYKRqED3OJ9stH1lXZoolFKWTZ6qQj7svPlCTIQFE7RTAmNnHfm7RmRzYYQYrlfu9bFzadd
/Da8YgDIGVf+D7N5V6jtY0sBl4JhLnthm2k8EcphyxBiT3Y9ORiLWdNy9ikjrrfLzbvJo4Pf1ueh
7/E7MGjZ5Y72oGVB/rCD7trDku6GEH8UeUETL5Sj7jD64zklmICohxuG0jCVSgTNNqbQ9Epdfv4Y
8HsveNABDnK5bv627YijT3vBw/Lj7gPzz/dBL2quzXTsdTejlmLKY62w6r6CTJk7tSx6ppzt5zdP
3a6o+ottbUko9rL2CtAXkBTT0DlZo2FTHx9eTlsT5XIpoMSKTCe9ea1sj3uNXuxWXY97JurF0AAX
EaYL6XGWtVNPFmSyH45DvTcphtcVc4FDtB9iv/2uBGvN5zvki9l98yTHpO90UnauPEKsluGzCBve
qQtv0dYLpew4kEB3QngcvE4RMaFj6xLeEtt1L64jLDIe1X74yDJNr/aeoNUEptitveYsGvCzUa3J
Y/RIrkbpSQWJ51jXBTaR7s6rvw+jVrG0TMvsSHgIRH4e/ZRFXL0vUfLqgorqD4UgdpwnIGQEn59c
f63Jmk1ceLOAqsJc6sgK698kC6PWrtqf24aDm9GR5FkCIHoODq99zgamkvQvUFGNonavptvnSvkJ
Cy9UnWkBdyCyQPvpAFHr7oXjmFwqy0kZxgSB1pOzi55LpfgK2WA2sPSSKcAAIkH9npNYtaCgWMj0
t0RxcTjEpJrWlih4H3Z2P8n3lu/An8Lhg0B4kbb6/ChZCyUKLIJr9vo2mBni9s5gPsWxjDKwWzVF
fMVG6CJluLE8ueRarQrK19513akbpMHSVIVZK/OCTBNAvxmeM0atl+hIC8azLk4hm/k706YC/UAK
r0XPl+GaJzpXFodWy5veXf3uUv7QE8pdBGsQ+qkh6XqvwId7sFhui48FeORazL1Fp0dYXRhtKWAY
u8YUyuKZADHvMk5+SecdIDRq5WWRk1KyR+hCjUtT/+ZMjTXQXfYDe6W4tzU/zKkm8svzMdUdWTi0
nPcJWK+y4DkaQ8StPUvhS7B+KWRmsI3MCejfQ3keSUKp3dZtkBs/xZsdlHekHw/wxKAKVMSXihZr
LX7CJF0/p+vUh5JhFdAjukahivzGFGWqwrd892AQGooW1+9GlS8q66rr5YfXIsetAM2FxWIWzOPb
ad11l0aqHJis2RnfkeJp4m7keitevAS3KuBC7SOlVAX5V7mhHqWzpv197lRnQWqsx3UCBR61VsyY
HsVXnLlL1fPiVXZmO9s6cyr+PnA6nBufoZhrUHYlIead2+rRDVoxhLvH8ImlSRm+rmsj2q1e0wS/
zAV5JeUdxOE6VMnLEenlKpCB+ICuHhQwi7cv+m2ThEwXPoPrHGHWxnNufvLV0LLKfC6MQUS7R7b+
KINnfqJHHt316n/ouz7QWbyKwFe5CYa8XcxCC27odbXFuPKzGRayO+MwyRfGIj2rF8N0Im0gpChl
YtHmKAjTVIqzqfDbo+6InMfvVnW97xS3KsWS1DTk2oNrF3xE+FLY3C4GVwQO4re06coagf8anG1I
Z2w6C+D2ISb9SlPhKAJSgAcrCoO+qSaZQ7joYSQPNIXn0+90/huti/2APLO/N/QICgn7EmECXTxX
68s357kC18/BPJ3SdvD5DQ7+CmnufAfrpU19x8d6kVudcpEZBbPJZM4SN3+exTXwD0po5JiJI9U2
/WTBZqkS+JL+nGgtNmUsE5SG9Gb8Q6k3q/wBwwv9m/Q05lkDYW3Cef0zDx8FoycMhPNBmxpx0uhd
AFSBsxLkExuGu8bqzZDsel/EqF4BjEJ8gdNX3Nzyld0abFbYpZRo5RZQbR8uQm12MVs5ZKiPtq+I
WoPJtPHMeq0hmCq4xpa/cof9zgut1950BQqg2owosg/JJ3jg7eIpOJGXVklqOT8Fyoo2eBf7c924
JIjNNwViNOIC1k6q828AinWp9QgfHqPtotiBp8XNleEqvpfQU+41mbfG+TjqmJbsjNBWW9oDhQKr
S18fFtX5qxyLbOcGqd5TJMteb8Utm9+AisgtXSgKUlll6ZMIC9qVHuUrXtdnebVf0cxUKHDLxnTd
XdgEww93hM+8Ri8h97xkKPh2//ypuHTj9SMHX7DrMueInIbKDFRY530d9LD+ljFsy2vl8AYIeTx5
paJARXl4hQXy2Nril/eduukYRSQ9MEUXlvz51Jq+jjL9CEJWZLg8g06P6OwtIlalqx1KRSeAUTCq
ONGYDnNZDsSfO8cGdEELTjZdPCUlfJn24n0XUZPVx/Rc8tqoVzjWF3EGshQOhtwObirgK7rVodHP
+RncOlp9qV3CK7j0waoUwGnjHrXXgtmMKCfx0ayciNPKax5ji+nPkOlfsqpfTORaZ6Zel7gqAA1z
Au0rkgmiXKxFunUaKAFP31t0r9JNlkFOzZxNUQyiBYvKFWwoUwivYSij2W1aXT8VsSYH2LJvM4Np
UQOVDE0Km1gIWdff7MAJEfr0/t1c9gysRHiJ9724qu4tib4dSA6t0RMeaV5JiBwiUzW7QULPBSlo
M93qhXRyxPr8ShpLZ6DVzVYxLDXwga/JCcRREku1gCplRQ5oAklE0BbTPhWKfITRqxFiNox7osA9
AFinRfGMHMAgowcrlnYpXeRKTfNYjkV6bq3Rv6OvX4UGOU5cFlQrso6TmH0+/wlM8l2mgElkdxTl
nCZmYPexQjYCyYFUNYNQAsKd6d4QqXg30p51wyTVQOT2PiewhFq7NXNABP0fx30dDxU7bK75rOWF
O9XuAEdcdOfM8R5ov1mvXt1Wz7hLXpaML7IbwxZTRZkCkme/qG2/RQ71zcpXktveGpjnV9fNxiv/
ChaSufYqojql1PPgokf5rW8HVIVA44jdcz9Cy/QxHY1HXIQuW3UBSUvmq0AzYwDvpxg1MJkCY+TH
oZ62BmsWVV/YiZdWrWFLbMw0sHgKikpALZoXbUa+RL4rpX83717XH7kIVW0HohdyFoyTK/G838An
6w4wggZOgaI/8Ex7kqkH/QiyP3w1/SLLr7Xorv8Pf79zlbd8lb1GR+J+wrt1YZWTGYeu/uq95hof
Hzq+FV0KSAVaT88Q8iuy7A4o7ZPNonKMxCyAyow2PWn6d7tr56kQ1KT7JJpk2LVRCwyL5wfIXcWM
EemOFkRe81uZwmHkSJQOk7uVFGNsmXhEOTL5ifGznXx/yWyGnfzvpNuPiZbm11U24atx1J9P/8OX
u3YwVK6LVuvgWoXlsBF2neSnoP/3sBRsmvrBPT+/u6d4FKbwy9KEHhal2bJVh6BkZ79AqUft4QhG
2UFQutQ7PYmdw4dLJEqmt9kwNcglbi9V+8ifL3p3TmJk+T2GwFf8eIoZ9SkfLSBvMhFoTOWVJVBR
3XRpWYaY+qWxnUyu6U7ENKQR44DruLqhVEDcSoAo1Dx4ntVwLYL6ZGePRsLfT2itOi/3ZEHgXAWb
MA0eqAUcC49k1fcAAj4uIXIO5l4EyeVIxOaKMH9AbvYmZUhHbHenAGEr062oqhX1LQOCN3XHhoQI
bDam2QO1LZwYvrVRZwFSDXiYtx2k557uIZ4ToiB0fWajmvIaVIMRHIYTz2aSNiFeke4M4BmYuX7z
iKhGQi1Yp7qXOmtlEjhLHM/WGxHxDqChAX7jPZyHAH5PFa7aYZBbDntQI/96MFtW7eFQOBJBVdiQ
otxjOo2UcKhRYdYghyjAlK5M+t4kLC5jt+7rGE8493oR1fQheynpCuFbHHtBhEWKsOQDZNCOybIx
3ujrJ/lHs1KH/MtpKPWH2oE0w1xqSpNMi9LwOo64wGujB0KOoLtgGFaDnuZJFuQuWxAo2+071xV3
pvJLJY9a9BtCJlLzo0M7iYrBcjDJ3kWTMm3KuWTV78N6OjDiV7XXpLf3CxhqZwtuhktqLPKtAPmm
mFpUcu1KecsMFmgCjZNdnrd5ciwQ6vDf4fPGk5XM7pU17OYLC90/hzmEdVlYTL+jph4qIh3gxxOl
8EH5d10JvbdjjGzNCnxJzYwTD9ykpflZ9SHargvjur5nOr9z3G2EtESGRALTckJiD5CsT4AqD5rk
/yHAoM0fy2HsGEifrj/t+Ce73oUtEB6ohBKAwX0j2aVVfpZQizRA02IPvFHUbU/5j3xpdDgCnejh
hjKNmFdLyMaAk/ZhGkusuY8c4sAae3Gd3mTtlgSiAiO9Ct4E5F3k2ECGscCawkAY6FS4acXUEN6f
LcZvz4U6sgSbcXq3UQrZ0zws97nJ4NYLxvf1R81r0JuBaYaTdXeDtJkqGDBUTu82Hpn3Sk5ddYvU
cB0SaWUalPC3s/o9a0lbINxcKt8Y5LgtNPxDKfv7RpPKFiB23ABTq7PG0y8i6SXn96fLivBOPM1G
NmWXN3BYqkcDb7mxhDdkS9s/q6fgyS+IpOOSbbaleB74DpciIg49Vxix30WMK30ucvlEhUTW23s8
dW6tbbY6n0WWhXnYFiLauvINSN7RpzxpLQ9SqX1HQaKI35FtcE0rahgih0QcHwf0iIVrRwXv0rIC
qCL/qw5wSnxmbm9kULv6im4SXTqTQgYTjBI0oXZhdzVMpEzQISBgPbgH+qb8iSoNR0+TY77q3/Gh
7ESL/w98LL4qwfhTf8bbx7WDC/KSj4HHmjXnzD7fJgSE8JHRRirdIRno4AKc/rjMLuZ19gfBpVC/
XguuGVm7rvGGvB11t/JB3y6gv7T0k98DvoZp+J76CqHvJQbk1TDWo0CUAEk14zeH+SRJeOTVtVD5
7B5g++M+RuHUKWavGu0hbnBH82aL1WbRvsf7bUUCFE9sEaNKJDpVExiElnBROgDWc34wvWGSRTOd
93EqhtJP+upfuuNk9j3De+Tq9eLHyVLaX08iY71Yv+SHS5x7Ae0uEbzQMtP0Ceb9fHzI01Xm1zsK
hMimSsxQBNdpk+p+wnmi8npltEXWkyFSuV4yYxMRDpxMKiGXgbzJb4NvsEnwnLIXSKC406+I6PQK
Z/fUE0GNSKd1lSkD4h7O4SkgK02VXduyyVPsdCJnVJ+6A2W62SJl810DDlo0kGbuB6Jbzg8Tfyse
WIkamDpDgkrdXvgWyfeuqphL7T6/WdvhnIi1WLoFoL7BUntGW0iCHJCYgfnAdHmSxde6inM/+k8+
qrQMyA7XMN9dFd4l1y0KxXST7iOqCcPLaJC4ngn6Harq2eKyoGkE2LOgvWVZyN4HmSE8K6zJYQnH
v2Ag9rx1Jc+LYq08j4rXJpAa+KGgBtYLfBNkZ7TcKnM457LNaU3boQ3uwRsqx1AYA50G07FZ/sCb
MUr3lBpNSMd+o2N7u+HLiPfdQLf29Zc/gSFOD1ZDMFIBgWPomKbNe8E3zE45vilX9YIfrP+GoHWj
CC91jKLDoVApQpQMTVwLazndJ5ThnL8L62N+GyUml+t/RpwyxShp86oy0NpFsPqu+oymiiLl7sZw
wBc4M8ULT3DtMHN8rB0IEGJd1BCBJpDx3VH7LbyA7goIZGvAqAMymjqDshB5ZOYdAVvTvKqLh3j8
gi9b/zMSMlQ+rdoPOUbZv10YjEkeR3aajJ19iUpTiYHUaoQdh8h5eGu1P2q/dFYL5uPLlwlIII3z
lf3BxMQspKHy7yJtDixe5vforNhHjqj02J5rZXaZQ5W/zdUC+lz0y74ymg7nerFYYuQxifLDi/ER
bJpbA/TmvXh9eOp9WA93By7AguchClbqACJlGvYXy+cS9hsEJ3xBijXDIsu+pnt0SlGhBqAId7DR
nNymDiLXCmAdgqUWQpA3AkFCCCy5KBta1A0syOFoOLXxpOnTuex2g+2u/BjZNA8AsP5NGMj4lEEV
v7bmKLHP7qP/H3D3U9X+SCo6fl9kBaJ8nDS2nJtGqiH1hvRy0zFOkOyeVc6zBHudZzp/Otp24GI7
yO+W48gNJYgAQNzTq48UPWs9nUT5d3KGYXDiZzndrimRtQolPev3UDfst0WaDm4N4M1vXaZeKds1
6dBVaPVEjMmhQGXGAls1+qM1EbUES/WtgAgUG8XsjPwdeS65TZ+vix6Pe2xHrtgrSCigfLH5VhPN
B/LWyJfNRIjANfd1jII4hs5Dxw1j0LYnuj1gQBC339sh2KZORDx3BVmcKwS9UcCrBGpxDTxjLDbn
bq/t6ibjGIv7tAJVW7MfZ0vQWPqMugUBCU3rM9aiR99BIH/UoT5I06XQW1yDNgZbAIsqbgiQ94J9
OJbIlooYcbRUAAYRRRJAB5rPhMs+s2ZTOBq50jgxpEE1iPAfG11NB0KEHko+GZJOpgwU0sWYu4T9
yBzQy6Ie8fq6VINWZkP0tb+e2T3JCKXa7AqRYo4H6gJTKK8iTn+T6MkTpYFScjbL7dQ+TeyTEqAj
+9W1ni34i9kHGJ8wZuaWx/llYAoqv2Vhxo4kkkqnNESPTmJWs1mLQYVzJ7dhJt10W7osU0vhHjZC
OSp3lAaG5KWxfMwseN2A54r4FAnw4CZE7ztiLyYO1TlJ6bC+u/9ahNiJwPkaOacIigHM9K3grHbp
hm2MHGQs6OIs8cw1CSprvf7is2tn1yxsLNXia+89kyB4ctWdmmFE6v2WCstYUkcCGm3e+WpKwduI
iNKJ1jbh4tRwXMK3Jy6h9pzuABqC1MHgEOdxxKWcTnbSc9XB81XM1b/E9ZpEgPyLLTBzenMZ4SiD
ywWYLQFXX6FFM+abLST4p7cmuhLurL53p/Y96XEEpivNlrjRq2lWVJHLPhyNSVpuHozzfTTZ9lp9
rx20oKHMQ4fVLlkaGa/2+6YxHRWymQYDE58YSoI3I1uj87/cdES9AvAnGNy9IqclGYs+dIK/I6uf
zLqxxKvtNsoJ42DIq0WTD1qg9DdUYWQDJpvdYsGGmcoJJcPrMFv87D5Lpm6PRyd8WyYIKX8r7tQl
+/5IRxKV30lGr68AzN6MQBieFFdB2Vk4Ze4TV+E8Z80VUz54bt5gdQXYAEQ5hwaE1dysFT28hPfh
+Kqi6N8DEaMslgj1Tylo5ODfkUfcVwWceqiNv2S8aqZc/sHo6zXZqTBAZHCfKQ82zlyfSHXdl98e
6LuYdGnu3ofstPLOjoW2hs8QRH9WSAKElRS1o2wunWwhQv7lPmpegm1/Ck7uC1pAWbvMJn6oQEpP
a+QggH8uo/jqdT7onDYQXhJJ1/Y8XcL1hTZDIS66GEyVzwmTUl2JtkbkyY4CGU9mDHtx4Ugoy/24
aSAgwDqZhjC2AvLj80GIZSCUmjC/+fR/k67OB8Tj3aXdKwIkI+dGlXKJj+4I4x7Z3wt6+KYuTs2B
jhVWW5gH4I+6upGiDAEgpPMXkxbBRn+SlmfVhh2SYRDMc/r1Peo4t+jzuMRbcJlEbxi8OHvYE7sO
5uexqDbfaFvbGXvSAE569aU3bOVf3o333LTSKTqSJLF6zQ6RkEJWkZFjvj/kAhtQk+GXZ62XN5Rt
wXkx3mtnSTl1HJOm/2LuKi4H2SoSSET9NtRW5pdeIJWrAsaA5s1bkdGVNiFClZhVYx093hvyfET0
PmWUwQi0lzaXrhPXGDqT7+J95GcFmf+pG6q+esmruTQF4xmSibDPgZHmgeFQJn3GyzEHdVA4UjeH
BSJrxHVLdeDfH2LhHzFL8yEfpK21Pxk0sINwrKyFtdJOfYKUYM36O9OZPE3ey5OZpcIKLDW4SRSV
eXZBYlgqBzqRpi+G/dWWGg6WJIfUxieUabWC+mMDFMKaF8PjId+jAu74bJndkROy768ag1q9wY86
PWLXf2c8DyjTv21DNErpgLYhMpGeo6hwlwrLH/tX3E8jkpWZr8+ohETguDQ/c8c9IW2RaYD1FQKI
CK43q+E/02m8n9WTkZpt7Q+2s3X6ISU4L1pcse5ZwyHG/Y+ZlM5AmGjMIpZaPvypNPewEkSf54rq
XODb97R+O5jG5GDPHnUlSo+0WLuSZ86gcCw+GS7F+Izumq9td1zyoZuRkFs+8R74ogbeKfZrBpGi
jHZ4sOZ1/Pa+e31TaLpj57DW3WQAG18TYB3hjrQ7FIdLvc+yzS5UD6By+T9EEZ5dlC1R1TaPYWlm
vIaxxFhexIzm7Y9GgUyB38l/nF7CJgUIuO9sR7KFMdbf0YJodL3lYcrhGOPPpdywAArjP209NBof
4VZxU/VEvlb0+/V0Z5+QFDGVxwTd4DXXRnoSMwFmyJJR/RltZqnX8y7u5rQTMRPYlubDj6EOPBx0
VvovSVxK8SBfbkRera/fsFDxOtnfRv6Fuf0oL2Y2vgr8MReVE74DmWbe+MFgSIkfTG4yPoAsWRW4
eyoq9dWIn+/RDM8zwO1MzTbU/rEdQsXlthNaM5LvT0+E1BtyL+jeMeIbtYxb5wGIU9ZKp4L2xvAM
P54+HcaHb7cZ4aTuARWk4dUGzS+R9ph4h9C5yZaF/0zbL7sG/YiVQzcTeXQltVByccEFokRrWMjf
+BwvN5rQyubrR2UhKPcSxDpp+qQyjFAXTtYuYAvx9CSfHWKFSuT2XobGOXPG/f0QpkbVi8WnZlH2
3GCOKU6Mvd3RwqlOmFEImfoBJvkp6vOuKizFMtsT1nVA8ZPT+NX8BZqbGbKbqMzKwTVWZmoat8IC
zk6LD+/z8uhC2cybr9uqNdtpMzVBHDpyBdz3WO70ZwinOKsvLGiwkUCVBH37ZewbLWx1pjOcChOt
bnmz6+6EDcKJhqWNjNjk1Q6FkPl2fT8GxYhp2FYgyFt0x7dJBwWqPHv+k4ixyp6Shhg7URSVHyhS
lnODndleNQGL2ZYhblz49VYMeBi54iIZF52Gi48OYHydXI+6nypjs/B/2djKvlcQpzm3MtYxBHDw
S71brnUt19XBMFHPVHKMcsqH0180Dh4zEsfEi9j2AsxgvOzl/FW84+kQxBKz9MTu0S1LMga5lftc
VRZw6XxI0CsoL+nlXzhkZmU/zSpzYFe5K4YMuEAtmJvyURn1P6IwGIKGRx9d6i8FKwbWNlbygBfl
ulmsrQf6Pi8pQmjwIT+h1Y4+oH5s9N+pTYxMqpO8/LiC5Ph8y47Puoy2NkQaxLqyQ/M14YKkwHDI
En56qqfe7e/bvl+dXu1KX5YzyYVSXwAOBpgwvuhK54bUQNJzS97fqCAYt/n0DuaMHanTHnRbpTc2
IckxGWCC9L+97M6zThz1cmBzZ54e+/TSaplVvBYtCYvYaHbys3qBToBMtmApiCjSHb766AKka9Q+
QVXfT7aO6XB4xA4iID1BdbkjpNfqrIkNWjJ7YyzTWD93ijx69BWcGTct0g+CrEZXUSNLJoPSFrRc
a/mahcvpVeBAwXUuygtdwjmpKTrBWqK0iaAYNV1rS8hUNexS84Lf7wohxUCw0lAKxRGU7ye3e3+n
j/ZJsKMVCcjOLsz53U+Q4I/xA6jsWsJoaElpBNuu3YFtPlLiToAjfdQQbP95uQMPhbdf44HTuZoW
9xeybhY+EpogXHGyU+/00xp+0W9Zd9PiVS0dUOqyeuhnGROUDjD2zxnO5XDLKm/4Chp8O4pVbUCd
fzRZ/6fsDUQpsogZMkPMfafiicfmZN3Oa6swx7s2+ZG60UIcHogsp+1WKZvtIecZ5/CrxrtzERjW
nVHYsl/o1FcGwWMB14NEgy0WUq8HMuotgzIbB629w2G7iSdVn8n122n25LLyVmLJzHbrA3X6mQx+
dt87JE1hWSlXiJq8EbtG9l2dcGTIkwN3wbL3QhIA4jjdOE7eGoYONBrxBa/pBs8/GHWJqO6v4TIk
94Ll1oH73ehwBziFoJuenHNE0wU4k/VVhre1B8PQexD7nqk+2BkUQjNpMH1sgr57FSkmPN6h+Ulh
rFaC1qKQFvJ4BgbA9Uj1o8fTKC9y2PWN6knXQV5dLZno1v9PWvserXXTwuGnaDRDujInGiWrl2WK
jWQLbUCNOUDOAMU6vx1JHPC1ZoUAkgw9gb+ExsPx3SF8QVumQfJC5/znjYDH0wGrZWsKuXhSAEcl
UR4rGJlIFnl7TT0LUCozwGz9Y4eQ9T2A2WXM7RVIwHfTOqdk7cNvEp681lUOSIV9k5jjvscSsu8Q
V33/h9qan9Yyp+sTkACVeh7g1OMm4QkcjY3ZzK0odb3XbegZGZ8RJ7Dpv90RSlSZKsulCU+fGRAc
4U63yy/1Yc3NRIjCbRR4UULO+eimFKumgcZk185lnPItjuTY6bCOEaW8pYQn7bSLk9WqMJHUWfpM
6jwuznE9LWVZsCqdQ1NGHaLOUt/8PqVm0Mk9XuK+Q3vHrwSgt8Vk1N7vUEvbtShXTJkkgIZDsv8j
A3n/eLa4hIuxMGQPy8XKX7jE1AxLkoYq7iOfzrJnYgISZLETJvjFqcd6/vD44UV5XApfKEK9ZUdX
ZXKrYzvpdVXJObOCDRoNSwVELRivHPzAq6qCWCKnOrj/Qp9n7xsT62nDDf3ZUBeT9VbG9Rk805wp
9CduAYAsQnoA0+QZOz2GJTaPwekWTrEDGxH7LDJsQ2DBRnMHnJhDQc1OKRySPzvajbBENkxJ4Q3l
/bnTCgGVIg2z3CFy9sp8gR5pvkwrc9g3NdK1jKHrRprtGX4cPKKSNDqxH34Y9JOL3V2KgJesSX5q
bSdayYUNzYNIKn2BPeNYAOQBBrm0XyMFduSKY0uelN5ZKDHrkh/ufUjAV08olh230bSuGpqUOBT2
gZGs/1SkE/LI+RMIewUETtqH4VZhUXxn8VO6w1RoLmDqh4Ut+tQoaduHuzP1gT8F68wp/qDARKpG
ue1jnifCETRopE/JcBvz0lzuv5TBukmJoflibWWeRCjTO7U1nqNEZ4YgpbKLh+WjE+wRZjBxrzTb
OD0v6FemF8WG5+IoXvtPuUb58llJB3UxB1Du5EzgqA8/w/KREXpOYY9y+kyjWFXXcl+m/+9Kdb6w
MIgRdX4xLoHALllcI75Grvevse6+jqaWA07bji/bf5TNuEfkDDWb9Cbq5DVO/plzVkyPMQg/xFEJ
CxXjgcfZFQ12Ib7vidMR4UCb51l34hn8/Gt3q4ehlZEQvv0ueOWH4kMnrAGmucIKhdBGspXN7wSu
kekbTRaEPlWSKwK0aU3iQma4q3CHsA5KHTZNkb61wZpy42Lezkv6Q9uHsXq7XPq1LLt7si7hXAs7
i7XhMnAjcoDSQ6jFDZV+9R5CVDMYdBXFXv/F6wLCsN1YxxnGnvIiiM1EmFI28AvDaz4Spw1AAcDL
AEhhvnh3S82loXmEI6d8M8RKD9a/Ako0AA7D3zwrwbi973H+9eOQK/CUjW0tz2QgIGHLumOx8uKq
pRMS9Zqz7yY78uii1rKoR4A1FDETkuOtBMeDtyHJxIzRP34QXPcVdE1fCpJEOZr0ujnOcp7Peeg9
7ua8lzIkBRK/tjkA6jcyWVDZg3JdrBAejCyqqcry0I07TD0+KpHnflEMsqjZc0MzXjHvqt84Kvkh
CPYGrq6EOUdF1Cx7n/7Eeq/FMzvQpUtYuu5sTzM9+tZQf27yNA4kKDZl/YEwsbQ8ZKywG5KLXW79
spfPmbi/PuoEFNava5lU7J+Uy6GGa9NaNqpYUIiTdSN86sSmoKjAoRDd5DbDDvV/aFE9dn1JXH8E
BZn/C8V/bE4zmXFHDaz+6bMhqRBGTe2cYtz6uxINieRHwNL5rs6HwJSxhcgWj8rcrGpFwC3nzirP
AstTfBiq+dx7FV1LHzaciEYa5hxMTISvEqkQ8m3Tw7jX9ZBqkHIMHPDgkj2DzN0zlMxlkkXq/2Qj
lgwlapnL4N5326oHrKjRkzQVziANcYsvH8jiRz8qZLgUO8/Wqd4K1v4nZZZ3n0qvAsExIFzHwAJ5
MKkcZA9x2A96+Q5zuAog+NonabxqRYNTSkuYYVtMfQZDTnGbQb/I6NICDB2+1e2IkAz3T1YHPNm4
LkBF6W45lpo3T78+sEq1w8ahx4JvqPe7nm3Wj20fxIFU9cHWjK4knmdcmULUNBlZ7PPJeXOsnsyo
su40aQIrzHB30m6BKdxwHKWNPN3Ir5RMfPO8tx2JmMUUVN+WPOLhRcPiVyIdA2thEnVf+1ABuN3B
9/TNO0OW2n3PCFFA3DwzDkzMJ6XsPMjTeqJv81xFmfJCRLuOP9fl1t8YXBh89YPaUoH3wQjY3J8j
h6VgiBFK1rSrSME4N2MBPnaSTxx95Clyx9PdjDsXyanp5yWhBNZSmUKwdUjuTtDGHSkptxkQC646
qlqdfKkMXAc0x0aQY0wYIaVaeajHe+SVJyEcLAtbGfLvDW6ETbX5kUceAPIJTejY59Mo9py2EW/x
lH8dz4eGC+LQIxABpOe2RE2GAjV9gtG583ChVY+Wxp6/cR5hrnV2qEFjuK9aOM0MD63wsVV1fU/0
E69X+/4akwkB4kRx63CCCnWmUaHwDpmSjJ/YnpBeilT/a/pzqIsLvRVBxlHX/EDZg4cSjLaU0XxV
LqLWJIwSwzyB4voksYwCg3U0zlavfUAvGayFnXiHBffgiJsGnE47Po2YGsZlr/OCHYDH1jvgdObn
3sMLVXRYW481kFtXEyfzgszEoeWRm5bxyOpg4fsGYJ6+GddBJRMnuH0CSAHEBkxa3rTLMqhY3IwX
8Efuss8p7a9FfmJaFkoF2d+RLir4EsHWIKEl/ea7qyhN+lP9pOXVvtAccdjaYRQaieqMNoC/R6aA
uFrDhVMHpmHx3hgerNhOXGzTV6/7SylhIXxiLItHDrgZkmJom5DJtXIFnejC2XmvOjoW31HeR7kY
y7cxy0Og0CXzgRduD2xTPXVFFR7J7fU1PO6r/LPyexKtTtzCSI1a7gpalx7KvzOKvrnfUtFFagqT
KvSrc0CdDU3B2Y+3YjlBpc5BAu60AQOnOeDvJBNLWSryKNihiG/llwNRsVgnAr6GoiAHCPaqFT+H
48MnsYN8etTn2HuDSlbfweB0m2/jSuYaMSDEYeaxH7lb425SawIetTQWxLFMuSo8UhP43Ef6s+gY
6/dv+FUnwc/o2ARk3hpkDXYC0BQt61tqfKEYJDkkonyQV/ylZZoXJTaioZGcTUuSxhgp3oI=
`protect end_protected
