XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��r�=J�T�i@L�ؤ��8T����+�p�$��(�).d�h���b�zz���/��b���Y[܋o-_�E��(���
�_.`�g���R<3 � ?�IѿR�I�7ql�$̮��d�яY�|]�O���3N;k��
V��l3l�x�����P��ww`�_؁t�_B�����ͻľС�f��z�%
���z��ކ��<\��Нpx��(
B<���Ǔ�x�J��!���O{��J.FO KXiM�'��-ہ�t�Vo&��x�T��\3��b�0� ?�r%7���=�Xy�p�6�@X[ҙw�{f�/!D_��:���P?>�+�ACC1��H��؏�����ơ�b���t�M������Ř�������r�S��}��-�L��`/�����"/�d�X��u�<5s{���&uOu�x�R�ӇC�]{�����.w�'b��;�U%�O�g��-d����?NN�]�٫�Z�ڶ���C���]��prո=e�:,$�Ǚz���f��8�2;\�B������O�)ڊ�͡(�1$Ƣ�;���u�\�F)�I�i38R�e��	el�w%�[���S�3��2��&⌲8H���9�T��So��y��.?�^�ʴrV&0VJ�`rI���<�<x���ԈK�G�`�l���*%�=q&VH�/��8�LKuX�{:�AiҿF�t^Ds�3F}�=��_��2Zd�Ħ	�j�C=������b�I'�,�6XlxVHYEB     400     190`m0�!�)0�`�+t�P���p>�8q6�B��M��
xc����V (9`�j_��k����xY �� Y�ͼ�؀�{9��kx�K�o�*P�Y��-�v��|�(tɁ+�&d'����}V$Xn<
�2\cĎ�����������Ǽ�T��UE4�`�où�&˰\׉�Jl��Ě�H�k��
�&#��ۻ�Ϧ60c���K�ͭ��^~�Fi�c�\ךk%'�`5��%]��7��M9�	�SF�P�c���Z���a�����[�_��;���?�lԘ�E�N�|s��=��j�OQ�#G�}��5�Xy���2UU���N�d��l�wUI�'*sTV9��t"-_��gE�8]�����o'+���X���ǖF��vN�G�p�d�(Hـ�XlxVHYEB     400     150��yl%oY�SPX�mN p\W�$���\u�Ԡ�N���JӿP}d3�?�ҹ�;l�M����A�%�y죉��܎h�L�MJ t��2�Ym�����}m|L��%�d�Q�
qi�|!,���-�٧����Wb9ԃ	�G��������k����f��9�}�a�l6Aą6���������+�%9�;��陔���N�Uec����ndQ�1'U1C�\���fݪ�o(c����İ(
 �J�H�<X$�c�no����k�^���n1_�Z �� �r��v%ze���V}޶R��(���E��;;|�% D���XlxVHYEB     400     140v�y|���8�W��ﯺy��ͳ:�Xג�4>�>�զͥ�����P0E5��x�f�;H;v	ェu�w�ڨ����!�V`�<���ͯ����,�z���XL����e���Z��Ѥ�R9+��/���\�8U�GzZ�a�7 @X8��8��	Q�,�S˵�sL
�#��FS���&�1�6��Nf/�2B2����@��W2HB��u��Wp����k��^��7�M�q6��+�?F<�1�s/?[�]=xWz�w�Ti�7���ՈiD�}�iQ�A��-��1v����{xtH�m���7}���pszd�%�JYZ)w1��XlxVHYEB     400     180�1����0���H�N�_��]��˰�5 eӤV��͸�ի7ֽy���{b)��_�;��Q:�!�ZA/zs�/U�|�ql#�IH�!a�0�����w7�ߙ�0�bEYF�Z�<��S��W<�?�w�7�A�\��5�)�VW��@�$�,���Of����&0,�6c����x������clH�"$Pكc:�2�˕10��\W�b�>&4�|�]�G�6Ҽ=�=���y؟���N
R|�c�����R���F�F40��m���o�:P2mN���^��c���h܀���!�� z�_7����^
��[huM�=����c�nd"u�»�J_ Uр����H�Z
�k��:��gو����+{���
���XlxVHYEB     400      f0y�i�)̀��He���Q�����5�7��!$�p��Pl��=��k?���)��l���āJ��-vwT�bz����l����+#�@[-Ȃu� �+�)Y꽍r�=!�i�"֏�[���%�1x����0'OeV�m��5еd�b��ҋlS �ZQ����e��6����]͝��6go"�7Ĩ�'��_��j��@�Ҟ�SB�4&�c�2��ei_�G�X��|CY��O�	ȹXlxVHYEB     400     150��6��Ąe�o��������'�)>�V��
{����UP�*�C���0U=���_.��2HgjTs��֊����[I��N������/�z>5b���:Hw�R��(R32�rA�zx�@��l;�t�؟I��⩰a>~�/���9!�Io!\[�9�Ƅy�ˍ*���G��i�0's
�h�@x.	3���N,���\@���WϦ�B���ON�x��q%�c2O}�N�8�l_&��A�qK�'�W��6��W���K�_�,�]��%rFx��
�u�KgQ٨����N�{�|����Dw� ���v���³_9�r`	vMm���d�%XlxVHYEB     400     150)zbh�G���0jk��t�INک$��f�k�5*�&*Z����B?��8������z8��#��/�W2D=��N�45�?�OB,qGZ�E�x��`�ѡx��#�s��|J�d�kYR�C�R&V��� K��ڀ0���yX��4G(�E��d�2) ����R�^���<�tb�����k�^"%eW	y��4[~c��7������]��@siSS�'��X����5m�:�=�hZ��-a?�K%>����禎J������`�sv�Δ��*��O�:B�Y5��Жh�c�V}� z�ZJ�������'Anz�	����}��hRDٴ�;N�sXlxVHYEB     400      e0*�y#�a����!=��g���F4�{G;�a��L�������'��������u��;�yy����cα{S�
��_�4��TeYG����#��I�j�Z��Q����o�#��#A���Z��ʓw�1����m�l�x���G[{���"=%���5C�9_8��)��	A��<|���-5���!�O����׌�k��Z��b1�It?�.G��7i"���XlxVHYEB     400     180oe���5���7	� Y����"D	��lX"��jE���o�MJ̠����dOd�I:Geg��g[S[T��鰽�n}5|QC�?Kt���f�`z�����J�U��:�{�����cW��R4H(dSJƅ��՞�3������?V#Q�QBC��ρ�Z/�Q�S�T��MU���"GMG'�
mu����9��1ܝ��!?Tu�L�g����S��'��N1
h����6/��[�;lΔj����;�BK��xl��Ԉ���Y��[�p��.���H'�w�嶿X����{���]ݑǦ|�R��/"��A�PB�����pz�T�j�W�YU����=TZ�����o���)K$I�K��a_�<Y��b.W���G��
:�p�*g�	���b
lXlxVHYEB     2f4     100��5Uզ�K��/u﹬-7�%9�@�ķ߬P�.ip���>LGu�R	m_�?<��<��
<NL��X(L�&-�>+����@��T4N�>��xhd� G�XH�Y�G��GqK��C'���a���f�8ܾ�S����a���"�	V�q��ٱ{
b��EҬ��4W&���?���M��jC�|�
2�4{/�05%W�g] 3ւ�XD�l��:S�"+�AC�U��0#�Y��!��?�_=c=<	�