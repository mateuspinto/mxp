XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��;k[�u����`�׫��]�G�mѧ�5=���v`d0��U�͒9J�������i�fT�C;9����R�-ۗ���	L���G���~�F�E$;^���6����`$����o��K�g^5t��ބK	��:~�-�d��P�W��O+W/L����.�����=ƪ�	{�֥� 7G��Ϗ):��s*�G�Ă1�Gh烾��5�Ŧtրn@�����r�5��?�Ub�-�#�q�m,��h[I��ŗ�[}���k���t�O�ӴDr0��i%L� -��y0���<���4MPl���Z���Ҵ����/ҟ��:��ڰx���U
�(��A��	V��c_�nl=�Sg�E+^���cO�Y"O'W�¼=��ɀ�oEQ�����'��y�A�v����&��&'I*���Z�Vk:=t��,n˼��<�Wђs�iǸf��y�z��ǥv�H�R�8��ಜ)`;�k�w�$���.�g�\o���NbzF���@�5r��c�AV���R��Z ���A�g�u�yu$�NĞt���O�A�Q;�\.|���*��wG����IM��$\�6j��"�J2x�3x����!o�>�̩Xݱ$m����-���T���Rh(2'�~ BQxqY�T^�Z8�N�ƍ�z#���O�!�a��Ԍ����:vSGRf攰��u.�x.�4�4N���cV�!�����ZÕ�!Hm� �ᆥ����3��E�/� �T�C���ֲ���rfs��o���b��#���[�PXlxVHYEB     400     1e0�Z��iE��t�~e,�E��$�r�ڂ�tx�~玂�)2w�S�A{W��G���c�@����&:���$Ǹ��*�
h
-4��1��˄��q-/�Z�����쏙P����f,f38q�UB*^��|c�����$��4��oyCE��9U�^/ I���d�Q��R��Z�sٽ]��/*P���4i�����-EX>j���� ���(��-�Mׯs��<L��3�5��ʹ���T�R��9]l7���{�@*�(]���Ma��{�-�D�oЁ-%qE���xڈPi��/� �161@dSԐim�A�/7�H���������}��4�+)��y|��[Mf�-��fY��.,��c�)u�w����x��lxO��ѳ�TA�慳r6�RdggS!�futBZz/��s�CFW���w��@��y��0��� ����s5�hHgؐZ���ޑN������`/?�^/ ��x�XlxVHYEB     400     160�c���{��a��I 	��b��6��g���TM��s�)#����t����2�ϮC�H��}]�CX�ѵ��0�-�QՋ:_9*���@�#�v��D�dL^B�G`E@��9���m�a���[2����ʸY��(.\��ؔgA�~�mNI"��rp�Ʈ.�,�e_����U�[�E���nva�J^4`|C���C!V���
@�C��Q4�c��[�ئ���̔��k�)��>2�V-I_j-D�V��BMQY3�V@<� �B�n�!���"�1
�m�ӝ%i}��@@.<Hc�=��{9SHlw���G��������@�p��<" )��HA�/Rl	F��,7�v.���XlxVHYEB      50      50!����w_�:{f0ɰ�]L�Bg�L��Z��]�d�<X!֬��d��*݉\j�&K��joOKb-����(7�D�p,�ރ*