`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10640)
`protect data_block
oiAGPgKGBarkt1mwVkPS74eviokV+0uM3D70xS2fv2skcpYVgCtMX4LgY5TTPAPcsfxIhQQXWW6O
e2e4gmSGhBhxHKmU3AzwEgEpfKEa1hGMw9yAp4DCgqCWqX+8kcEM8uEFtPvSaPg+pxW9J7CrVjDP
sZLg2e0SPGOJCQV6BhNeAeLPsY5+UhQeFGyHA/UYuO/6stkIwzBo5gcYs0B0B5K2+vJbrsf+NHmX
Blbnp8tJlQnNBhZzplIp3ufkakTHulTlHSq/KYxYMbq56GREFEr9aDbw4PD3xehVeaYfNuF3cidM
yizWQMwex/jA1cLpTYFJojpBqxNnaFLHTLemQjygeGYYV5SSbulw9vUmW/eONstQ2+IPVMSX9DYH
sUDIqTBfn3OMVzCcA4FMbrpBgjDWl/8PyefpdJcd8molM9COVfDyvaP780zD1Ml7ZiYP8f8xKNYq
61J7kkr32rnFBGtguQuBfZnBZik3VA6i5jGqoazsLaNt+3bqSd0rXXXfxxZUXsdwx2cWF4Tf2+zp
ZfwH2aBPeOH6cBJ6iPvl8WqHf54O8l2Y2r+TRMeTG9KYxkFDXAGaHMfQA/TvpK5C/xw4d0MS8IB5
3wAMiA1XxMh5BZsfwaP9BQBZ1++BTMs4+SS8OUrFuUiqJVTPgnUFi1Tep98cf8C10j0EhXs3se5M
btaIfN7B31A+Mb/49iDtlsqL79Ar9kzRIlZ/V1ZOUUv6eRnBOMQfmD+0EcMpNW37Nrq2o5BG0OBd
IrNCD8HiRnyB2As1vDai1zbMmmZyJBjbI1sZQ+kARp6KBjiZ+ZgLiX5kMfnPHIoQu2yaef1g4ZB/
6YvpuxMuDkvR6TDHq2wcVuhpPoRSHiuw+u4tsqCk/PH5OdpqfsKcIB1hAK55ig5eQtdGvCUJ0yUB
rpIJS4nywcejC9PJBbxVZRtxnHr0ZgRmtEZTKJLBjdB3Ip3Pbyg8iCmryVMYaXk1wq/DBu0gUdDs
+6KG/cynMX3ZhfTAEiknTM+l2UhSVP7v/bvpB8Oi1d32+cTo3DQ0S4BL2weukriWufImRTEXPmRs
/XckfJCowg2Ec11YreyxUVz36s1o7h6haqE03o0qambOMJqTkGz23kzf3BPR9DH+ZDN8rGPBxJ2g
wImGU+h2AA3uilcRq9LHkFhqQtAnDV9+ZhHja6L6+pBb67VnY1Q4Dm9Xv68K9wDq0RC3HfpZMiIv
WETyCqSH62dsAWZUhDrDYgWZA/cLf4LecZ6nVr8fTsm12yNZ3aEAIJ4eh9TdHWY+DOySOMoWlJsD
Ro1Oq3rRQjSRlLEw/Kvjr+RuV794NC3+3ZJrRuBC9U7YSm1bz6hJsXBKPJrU+CPsY27BdgMzR018
ME2iBSYk5Ur1R0PGa8rGTbvklJedqKjGGg7ZRJGoDQCAZUtaJykNzXOYsHvvNZTaA+/6lp0L/yh/
mQ3jWDRYFb5UMjIZliw3w4xxCTmPr4x+C2DoLK9yUFrYDv3q7NkbSQrSXQ1sJd/66lIUVzcth/Ri
UibWtbhiSXsBd0guVjxswR4kDCbOUPGHS36PEEvczI5//m89jmaCU0YqlNNzpwKiOVK4+Rk7bjMF
MT6B1apOJH5brv89nftMT5gig8U6V1KKByIwK1RDwVIMuU6g4B4kJMGX7ZT+PVRH9eHbbhZRSQKy
w6leSAve6qmWJuo8rseOTr0KOipvFOTfPCF+MgpkEhbrXRgKmSN0nSpKRI4eih+lT0HJerXj1lpy
vHovfcD42SN4iI7bUYjz4KYydU9VZRRSDDhTOe2BjDhciZYg+J8Gp80J8ORl+cYXfaVUkPf9gLNU
YIm1jFmsUpe6hynym6+uGGyREQgANloMkyXlwmvD5ykQ0VbSanr67tIC6kCfN9LerC0zARUbop+j
2l/0mbmwWa601wP+NV+XnpV3qqFCghoZ7Mfih4z+NzV99yM9YqD0qIkz3vqJd0P4nqv57oFB4aqr
WvST5ucuXoHjyYljLQ6jK+ngWYn7d3EDBvIIusA0Md8EdxeKRW3SJPEjs+5JITTLvjOfMAHZ9Qso
J+gkaFoNbntl+CTQyveDPV6AUp6GchKcO0edZJqA+DR07h6gD95XKxNhorE9ey4fL/PKQIbfbmDZ
K41jaPYjxK3KP4ZqcuRz8O9PBah+1fiH7kz5NfmT7/WXrQRnLUFT1gNt7BNSwqmJCieHMuLQxLWa
mduzxQWSVFoPmHS5xHcwvMVHM3v1xZyGj5/dRBPPwY+iT4Blh5LQihXilJYGwcctZn/s/LwZunsv
yI/2Z9jvzSU+7KJqKMZbT0CNz5Q9LkF6e+Kc8TfpfpT5Obig+LqvgZuRx7oQ9GXJJNeXKDIR3uvS
oaDtic3A2GMOe39NB/uTRObiWO2YnuAPK2nFk+pIM3gIK0/7PY07KWmfGNvQQqTbKCXeLw1vQtKW
Flcxn9+VqKF1HpQAmNxxLktPaqovb0bx4vx1lQLYY3+X9CS9ZTWPKffU0Ah2uOinITUllCF7TaA4
4d/lnPfJhadQal2mDBPLfXq7f49DeaYXrzHNZvo1BhoW7tWrVUtneS4SBvso/nnKq+8LqbMJrV+X
EdINqYFyyC0Y1hmlAyJAY0GBreQLo4gm3P2zXCj/w8hMcJOCKoQpb2mt982PrRXyccRfBL4pwnsZ
mkCM5BTvdmqgpqME0fcYU9qjIw0nAIa1uOjKalKJzCPTAW40yALzbMvRKNOu5oViYRWF7sNv4eyK
2xo+6/ie3HIaCjB3caIvY2WnLnW+PVuowDcFNYKy9DzBvagNtqIv1Jbo/j0dPLsOJNcR6hHFtGG+
08zhMOAODp/fj6t3AsPL6puVepPur27QcccFUj9uwcNHblF0o0drvgsaUo5zsCgZyVs7iKAO/009
WnpmPVgEzejqQUudjkCYqUOObSl9ivByZVex55oCOSP1DmedTarM5CfsUrIZggqKwxi8bdCQusjT
O0NWL+Yn4HFPUbjYof4GA4IsW/S+czlUWfuaPFb48L2WRWqaNjqF5ne7lCoZYKutQUV6rR8/Nfc5
CP24NEpj771gkQl+m1WBV7LbJNLABnBIlWp4dfwMMkbs3ag5ezzBsnNG3nW6YRGLLP1Ls9NAFxwG
WSjcLG/2NXrejv3UXbq1ktCDa71waC+bDYvlMP71HjaPcTP7+WXkpIVuay42S0mMurmB+g/epDbU
IVMqHzAAo1nQyjrLbDw7sV3lYIWFS+66oenj5d8GPPEBnLAHUzUeGF7S9dl2dfLnRHvmBQgb6jFY
APPDjU4KYet5WAGUltPj2AU3zhGyYky69k7Ce58I9BRRgyqqnSYM1+kM1kV2qpIvXeOC8N+U/Wes
5r1oK25T898wq492Nt+Bi0rWgTV1LQeiVPbyFiUvjb6yx+E/UWlLh6g1drNXAN+hrlw/qj96FNjJ
Lew6xaD4FZQ3egOELFF+F3j0i27DZA9UWpzfpygE7iTT1/JAVzSEi5b11qJPqnzxvzHfROsANz+n
SABagokjaIGAGvPh6rSTnxWXgqHbkVNpOowrmM77IArM21Ey4QGG9mUj53NvAvFmRXy4fjcwDRxo
1o7kC07CL87qS7OeITiputnoebzS6FdmwBohslIHjoG7VtZ+hmMPgTLVuwrAkB6cnsp+R0D9XZ7M
V/2EZO/XgyM+Q0zQ9Vd60JJ3R1zFuwypE82tHYDOxop5rgaEbn6Aw+lt+DfMVZt2xWa1QasmuxlM
/1sbqz7jR/h7IQ05gY/gzRwvD2N9J1vPRKgCx8s+ePxL6FUG4num+3R08JuRdt7L9wfb28KhmSws
fu61ttuGE+AZSDzlPK3CzZ+mKTinl7MQpn9UCcrj9VdAC9Ct7gGaBkQeaKJAe1QBtaIIITPyAZ0y
iJQ1W6CrYbyHYvDCNCnZb9vVrD3i8RwBFQ4OP6w2fmGk2UbfsXuY0yahWYj2oZ6zsafPcnEUmsT+
hPxKGt/0UDrsL76krHpJ806xeCjy/m/biiTDQaIU2O6y86tLwywxfuvnp7LL4U3AfF1WVfFr77EC
/xlH1MgZlFve/jm+lZw6PG2UO/nx4q8JTbAhAY1tLLqyP30nay2rmco2gOQAu+060zuhnzMm16lq
Th5XRf5Ktgno6HRwFiCLTRDu5pBpWvF2g2nKcPuLPZixfHHdudUevq3KaAfPv4nn6SBgRuJ4p7vV
TRfFENynQvOuvTOgTaxdteS1KLq047vwJMdVXrsLLsHuMWKe4NMWyMh49l8xl8t9Bwli/4LUWYTE
sXCs/EjkgHGGfzPpSiALw7k7hcD0Ewds7OGMPT8p5/kxlBzxBlGipaar+wh5iq0bzu2KH+KXKXLu
R5mb3nNbDpoeTtyeqlh0cGSprsFEtsVeuMoGvpr465hZxdaUsovs4EmJCFOz/50J8KjZIgxPvL8G
IPyTPDHT6zEchwKP4+lDfI1MAQSIGDcmVoflYQWSV6nDIH/qfEFp/Es+hvf5HFoE/PBP09gB9CzC
Hxz9EN5KJzYj+AI5zZvCxocUoeMWuwDst3CVmJfaVBjtb76Eb3RmBDW2f10Ve4Sm5WndUPXR/59k
nkUMoA9EuEm7NgRvz8V46VjsWLqApjHaShDIOjK2UAs5ObGFBTguQzbEp4WcmsMYzEGckckDhUGe
+QRXbPQK3nkzm5fRbayou8iPs4RUkGsiFRzvi9yfHjmMILk/WfOf0sn3nDLEqIz+Z1cHFg3RrVPP
wSqCx9LzaCaQbWHAo4Z4FaeQ2Rr4fhzP6EZsmtRGu6lFCljg7rjL8AgS/CPaGB3pfMZ8nKEyw3oQ
5pyVbJZqQ2vTgMAaSRCehlLK5AV6nymgs2ExrFRFdnqP9MqwiAz2MwyHa3L+E9JK1hJiw5VcFZza
qMvODkONEGQ/u57uK/BrNuB4owC0/x/jDEtsXH97e2ojMeoLhIFHNV7qv2DH4ZS9foChLNO1m5oi
J0HhJ93uzN5bkHj2n29HnVVFmGR0oXpmd3FI/wW3Xj1Sf0iLVK0pzWJJuTp0q7UETplwnWn52hJW
w99pOO6Dd34H99k1W8d8nnhdMWnOvfBbZCavn96NmW9AWWyOf1Sy7FUIXf38RA3CiHc0zG55ODFk
miHyOusFpZvcbm6JXIyYHNXoTGCqDGLV6Uj5QGiPUKFlPdlJvDMdBFMJMHiDCvmdyFmaS0AT16AU
Wlb8lS8jepwIWPWhjYSUZN82gbrg9eJfnQzfq+YEqPxRe43rIyAAt9eh4xfvXXJHEanLyI0LzQfX
8Sd4iesG+hKzfHO1S/ODMEfkKYyM6Wo0b1bUDIT13ltX6S2uhbCM9HFuY+HdIb0F3a8RgH1prDKA
quY+C8/Edf8nVFRDpfOOPatBfPKHKWC8EkyC2F88ABfEag8p78PkSAPOchaMEqF8bwiSMhIQzC3i
O3UKApnVuHb/mDYv2PZK0NSBigMWf9GVo6R2Kvff+EwjQk7iYUi53ijX6+qI0NjnngvLJTq6Y57k
96A3qphdWHBauZKrFIPUnv/MyRcCnSURE6OhjM51s22RvdKlu89waA5PJL+rXhpDTu/e4QUAc6AK
VGNF7LwgMcXzJ4JxeM6joeJpzbdlkvADt9V3IG9VQysNMVytnPDyhUtv4UMIjUkvhW5QgE4ULRLP
Tx80S0dSJ4FJRx2l6rJXC8tZT1SXHKX9si2lPyBMhqEyGPv2Qxc3JE0u+lIEMeILj6iyIYS+U3An
7cj7ggajCdjVTRR4y4svmA0OwMtwN1gjMmfvN9ySGpfqYYlM9ST0hXYCka3HwL6+aM1OTYvtbTWa
muMiqBn7rqkqAijZtZqj3aJxKZs2uAiz+NIoEiWsaZ+IMsm/iuRXCK6mckwI0dvbRylQ9YO8MerM
3xB/lNs2k5tzo096MiZeSf/e+uu0/an+QT7Hf+Shfo+a6snXHKC+earzpA/Ds+61koi/9+9qUI3g
AYucP5CwNoxkwPii8cc/FFzCJ4s7uUiONatbWIPJMoxtsXR5Xo8aaVr7XsG7Uvb5xHH9i3m7+1GD
awHpqn7tEFbquH+cTxsrPHwl8mQccbjpdhjVssilUQTRFCey1mdMELPpHSeFvTVyznkGOrpwe2DE
4F3eP9NcxO4i1OuYObfX/cma8O3c4Qpdk71EafjkUJihgHNgSq9afmlrHz/6j1XHbY+/qYCc91oF
EbkssbjCLweF63rlmS+3rKVQu/atwH3cgoNvKCXVFICzC7aPBG/eMG/6yLrwH90z75DRuSHH1/EG
R7YbcLg+wjMWHwpdNW+1uUUyzQ9jsVTIHJi5Nq96T+NqDLFIuc+b4BaHV8IZGIsrxA/QCYLyv0zW
0JmO680kWAszXEJkoEL21TjS8Ow43SXScFfda5OG7hlLxMVymsjnJKTF/Q5mMp+Msn7PBvenmprW
X8JqXm9YwMWI21i8xiR4rgYbQq96oe1QmXcWATIWsQWDleKLDq6Xg+3tE4uZXpbZfR+5UaSR1i7y
Mr65YKMZl5wday2t8BSWwYsufbHv9wbVo71BGHbL7uSRvIh1IJfZMgH8fUDnjSwg2qVz6DXubQzH
Oh5L7AUIGKjmlKCfNiVTouz0MSKzK0nE0LQaQpebmVOs4FP5XXxpqMxxBZlpzuu3QBzZPUWETkV6
f8ZFyEAipodPLofOPz5NoBoSzzz72/1CJfXtwNK6TGUwFAY7pxMp/MwzdZNUGof7IN0/lfsUqFVQ
9kwXniyD/O17rFa1ZHaWadaT8no08tIINGg2ZC+7qquJZhP02ab9P4CAXUGUiaHqCLTr8RcEOdj2
W3wswQvNjNLvyTP2jJOY1gOq19XuhVafFpOZXCwhAE2ZvnT5wmvSte424mRKP0/w8/wbW1rfvecO
WrxRJ4e/DWD62JjEOR2g7Ct1wTa7jstqUdG2AQwwGuNMGiASW4xfmXGkQZ1oa87+DSLrec5WTfIz
9NS/62Iy8M+PYGyfIIdIFRoppE1AqmHy5epcWRTxCaYZ2Y9X+XGJUjPIJFjW+gljLSKDgg7/oB4I
liaTYYTjeClD9sqZ+7UORTVXUv4BKoo4/9t2JgZlruFlYavTlt2Gu25/Q4ThuiyPNgrP6V62Av01
mpp7z6j9nMFr8wx++HwuCcDYSIpn2IeuF7zA62bGmWh8ON3kCAremVeeza2TVa2jfVM6ztlnnWxg
mU91rNaJhsZeFqlLgAs94p4GiA2kdZ7yKwJNWFH4BDSukNLAwZ4DcLakLJmjx3o5Poibt3bYUBwz
x85auA772clwWa7ZyXv/2/Lkoa+XOL+5xbQYFhIfz9oDhptoIDnFZng69IOetQ/u6RenBYPTpafW
pwBYLVzWGGiz1C/MH+MZsJZiWEnrVPRgjhuqhpzhVJm3Fj4h1rKSbHwOdX4qOq69kHovnkhU/upR
eHER+aWhQMMNdbWFsvUL3Uh3UguqelZriR0E/0+1/pqJT6y633+nqrrNKaLhK4ZLoGPXnmb3kkpA
UPQcJODFfSweIw3CGR9w7hMKuGNImVFpOTFjN1khSem1uYmugBwmNAEpISeAnUcMXZt2Ac9tKIxR
BExMEMpWn5cnfWoZqIHgGpIaqG/Wq1zx0051P8eqh08tbx/Rk6dhk/qQaU7ojYl+cX84X5kqI7YV
p+meLnLNoCXdrpdK/mHdJwsbPiVMIBzKefacgH/Xu7aqZjdZo/rNuXtJMeuOlfcUoY+RI/K4aeVL
Cyyn3iI1SNPJHJyhkxZPz7J5W1G0cPs7GKz/gj79IPD17JvMVQEXsN+2YfOuJn0LGhnE7x45CZN0
HO3Tfl1iVD0Fsn1Hw8n7P0q9NtHfarwNugCIMV5ZnEmd7BBrTOkivlR29ZszQ9T7RlOe4A1LFe0L
0HbrvAtrfVFy7rgIYFhhMSgmgDIvqeS3ElpVd1+IngUEP2fPBlZjSbz2Oy0T/eHNb57zUd7PRdkg
IhPMv+o37bgPDIlkKVwGBYcj1V6W5QFG/yt0JYuWd/Ialuf0M7aMhBZ9cj98Jin/gp+4c3D3b/l3
kEhXA/xIlCSot7OPlURMZM7TkLGyUDoaZlCCkPv1NbZJK/YZmWFNPSkYSkzRfyFSAeYd0HzlFQOj
7zXysS7FhjGa/8fpYR3IpRZGfJzdCckZ9D+9TnFOywBSihw/OSQmRDcCadYGdfW6dPsdJ1zB5hbH
4QtpTrfZBa+GbCBwpwksITcOFPiKpJz5KmlnoT8150tcBD+WIuR+E7frNE0jmAjP+sPRsBLCtWAf
4LvVDIoNI/frgRn+0K647PqLd2si5crDncqVQ4cYqNppWhgRc6xplemH7QeSbyC9MIQASdhepr19
nIn9bh7MCA36rOA63ZmZmZfEQ/5wWklf3o8eKP95H4YO20aeT6OBelZqgTvXo0Chtia9p9upO+Xc
WvIP6YU1mkGRgdEvUDuxiOCK47fkkIQwa5EVdUEDzwOkdwz/R3t6GbFpqzoNo+IQegaTufX3HkKb
u+rGha8WWjWEs2AJ3A0MJ7BmLUn/nCGwyGLAb26uiBu++6i5GAr/8FGp9LoU8SQHXMhOyH9cSsRo
QGR++rk8O6Oqn2BFKlXBDacPG3kQhOVn6qVgaIvN7hH4LzNy2zj5jVwVO4kszLKFYma7AiA4YpXI
i8ye3Uwsg+8E4z8QTSn7qw0Mtt5xKzIKHkviBnhiN78nE33nLaLu3q4Nazt+cTpEgzQBnxUo/8Kl
4QXbyxxN4ypMA65rRE2jDB9DVusQEnQU5/HaLy0fdHKOAjTLFQmBwCx5bEKB+fhfptjiL+38mSUM
5QexDBEU78aeDUvwTZcXYfoucuOQsNZgSuEg63KuT8iT9LXCUPntOqsFqtKwYWLdptw9fx6VxiZz
du8fsTnv05tQWe+ztM7+1Dr6AN8BNXfWvZdASOYzDCio6AUZzTYu+UqwDXrJHS7ZFNl6mH/Rh2/R
Ir+h4ow9pxtK75sfYVxb5OPVr6I9FFftvFR5Ubxf/qAMvmNT8PJJFZynHvNaI5z6YfDwtMTjDWAC
E8eUQ+HwOlUQNEceZtAFM+x9nabpaiApumj6zPREVjI3bRhc5lqwkf0+EAYUvkAH1bPv+V4JgOZ1
2yeAEBPIEpAhUbL5T/APIZ66ZM5bmSWUaBQZhL5aUEC18L+abw1CDLBGnoeOSIREdvB79f9oqECc
BAxmt1PCcAHuipijPU9VLg2tYnLgP7dCPQNW091uMAKrAcpff0e4cQHGGf6L7rLS0WHlY72bGSlC
y42dzDvt+7NoxmXqvrLDr8rzGvDRbsVVZSfPzvx3VAncgboRA7Jfe6FPOw/Fn0f4ir5Gw53v16cl
BD/u7IL1VSmycY9UQ0QZXF/JDiP6T7VtpIRCgVW43bG7MxtR1XPoeJ1GqSTmW92+uAObebQsh0Xo
s1TSa8D6dV69ObEBvChFRUK0ZuQGhyubv5n/zr8e6VVs3/mWkzUcBx3eygnCs3RxOn0ys20oCjac
zEPOdR1tKDbsMZUEbiRoQRgTKInhHKU2mZdnZc09Vc1rz+lxSfC0vGKZBNlk6QyTyrTG2ehRdvrU
tUgEOPHPyNKbt8Yj8TLzHWAnP8gYq30qT60FVzdjgU3Z4w/7bEIqfWT+GbYjvRrHbonycLvncNDI
nZVH1gYQSKsNPZOmiZVea7aQPK0pB6OPJPMt/WTiUoeJdkmLEeQXmKFAbMtqgxKq6NeqLGfRylYG
xYRk74bmCJAF4nZmCpNWjRtDqiPpbd3nLO7zew2+kaOwpn4N7x109E/zxb00egy+mJ/zWMKDkLQu
v2bgpgojz6RFyRO0M5NTQKZFPprSUmyaPf4GVh5CjcXItdtl8Y8wi2mBYruN4Sra4ZNB+MkTODN1
RnzG45D5MmVQjtzvuzreeI/oEK9xUQVu+6NNqMd6dx2LGSwBK0FEjljtS44NZOsMY6HVsECOgRlF
iOq2TF0odCEK0yFSM8ZussyexhqEekitYCnG/M+9UDSko2ZjYRksFz3AgZKqiWrJ0gty32gmFH7B
cKcalJwlwIfhrvsfnel8eixr74yH+EKJuzh48/jNGWCs0F0ZT4I3fkSFsZCS131Asw+AA70OT3N8
a4FauyN3UoWE53QxRb1MFQzmPCWfQ3XCGRssXpk6OEdnHiHU/JL2Fhlw7KUqI0ZPxH9TW2XwEkfy
laSGEmSvY5xKz/4qAdB6XCk3fwRXAIy9HiaRXrBV5+fY4J8dxZfL352Pke3C+26v8P3DmBxCwGIp
uR2yIDm7Zjgw+N0HDOkJYaj/LJ5YTcKQZ+gIAtqhEW5TiH5iKN7xvfyy+hfTh2N+GZy0RZcka1EY
rPI1rFHmjeuaQrNA4sxgv+uiO0coVzW3ST8oBYttoDOhKHPwmDsyCHh/S0mPbID9Fy7mG4Eyer7f
MNzahTSLcYD+glICmJPk1YMje0mbon2ymDLvwYkiKLEa+12I/1gM2O3F9JQ3bp4ECo6LLIKJMyV2
V8nxjxF78BJT4XQm2l89phAO+XF/HUkdxbR076yzU08dYQ+Lg6Y5eatD//CmrYkVc3DKy+86uSJl
yIyNqFLiKcVFhO7xsj8R5TJzM/bWxKn40FXVLOxrkAzdjUaIggrEYaaML2POEvMxRTaitHe7Z06w
wJqgQdvvVMf0/tGsOEuy+Dl2BNoZmKMFQBG4YUUnLARRQy86Bd+8bDx7W/sZraAy5fqBXNA6J7wL
Gl0FNMzqTaOpacW7peXn2HRDnIfLUboJAFMFilKgYVn1cGMXIk8e7Thk0XCuhDE3fwQhmJlbTtxY
PDOm4sXok9MbZfjpuDx+EWk9fTyrhOdT8NnSbQhHZvCGXHEkuCN/3908/GYLiUUUcuJWZpqL+412
m3UbZbG0a3fYbX/s8OEjDsadpDI9MCoLrWQQu5U90k2LDaHZ0qeV/SLm66msgJR/TBkVBB1w1Hub
ntQolbw4pD1/2x4Y72MAxnx5H+dY5SJvRmVWpIoR0+hXFh+hq8gTxeuIR/p0sMDjwHaJ4sJ0KR57
HU1WPmF8KTrtbMol+M/zjdO5LHDmuGs3AsONghABVA3EWk5dQEVKV3KpzXQ1QkjwFPNfJp+XNiFM
/Q/UZOJSuQ1yNyXy3rAnHD+ZF2duC87cEnNxxCu4JfOgfA2GIlEO68iWHWv6t6lJ8XUCTnCLJ3mY
bjgfLANwWy5nycTJlhGjbknYNSNVvMKsd0DyIRQYNW+rt7P+6n5zKo2sNeBuxEF2nANJVNwmN4/a
VzhCHb9wvl2r24w1aulwJeMiOyC7/EVhSPBFMOwXsfZuhcV++0UOjS06x2koUwcD1t3O+iSG6m/s
k9yNeQgD2LXTJ+uX+afDrzlGu75GZ2knBZrTLXEcnbb6VQ8DhjMk2bkOA1+Uyria9i24OB2opZtE
se3ffuCWxvxswKhYwmOIESA4XnI59atSTYlRIA4zvcO2tN+tUMBBEITv1zaBnTvk4LgvIoa4ZCUy
vcg1tx4MLOxpVaDWnCip9+lCmtZSinJrnl2fyQ5YCnotC97bRDgi6UVmI7Xv7SJ/lBxvW7RN8GoD
zGbccHga6UwFVBkF59k6lSoewctHyOmG+wcpl+6XANFH7nV0jFf07mfSABfIH144zi7tDCBoMXVl
283eOgkNRjWKS8Xne4tTop0O6MX1SGHJR00UimN2rzJyc+LLYj9KKSPDQWsFTD5YZMlm3XmnJAIT
0eGk5wkXMyLC9jK1bNAD7uKfbGDAoF2HQHeoQvNqF/cSRVva40YEs38t75Kh/v8aMWOaIZ1s6JqT
Av71as3mmg3cfUTujRTRzpUYj2c/G0cd04ydI64EXq1qzs79sXpqc9SH6poKHvY99terYrx7cAUj
gyIHnBlz4ZcwsQU7NaT3d21HMMtp/KrtsUSJE1GG50KdfetTCk5d0fP+5xcKfrWgdneGD6UKpp6A
TTSoLLMZxYzuuyKaiKXQn90/aIZ22ci8L5omnRHqebSMXrLszpfVrDLM52Rd9HbXHW6p98/QxRFs
+9+I2tTSltX16viQ9RukEtQDGvjzZn12Wjodbxn+gazfQ4AC5H38SQCyP0wufVZQ3RZOKuldjK9v
GKVHUakLHyu6SIkxutgQVu+r40p5EQYGjXL8uMicP1lkVctYlvw6Dr2hTZbpim0ic28YzXR0LU3o
1ufL7ekJKX2HeIO5O4+1TnM+fvOzYVAp61mN2oPAl3mNkkywNlu+WGCB+mDZs5QFyPiFK+7OLyYN
3ll6NWgubK12M0JHbYOOZvTT1dGkb73JBo9Jq5WVgDM762WpzPpMKrCyr5B+1eevG0YGFfXlV8QE
dBEXMxnqE2dW8ctNFux27AnA8hmIYyd+1DAxSAY2VReOP3nnMyJkkSmHdrb1uMwyZRbHy3Rv8S2C
3ty2YMoamZMvX7JYlfVgegpW0VEwbNCL94TAnyv/6ycdfttQ4h6adPfaEQsTQ552L11AR8yec3tJ
Y+yW+PoghnuAaTaTjlaaU8UltB2dSj88J4OAD5C9EXL65wUSbQfi9SC5MDkV2gow6LEkQ8rwFZ6Y
JcJ4xgwgeDu2cszKju+SsnysoEkcYWQEGP+aJxZvVd0GkaCeCffnk5tw6mA8fJjbGinq3qhdDwRF
ci7ouOGiDXl+FVtAmaGUMar/2lkhR3Lk06ANl5YDRRn9ZO52XGPnMkay64vxwKsYODuta+A2OA94
Rxrsa9zwVrSdlxhefJLIZOINMcU8sRoOYlQns9c4AiBo8Sio1HwcvJl4A7rG+XBPxephz69gReiI
pfs3KtrT0ZVPg1+iM8BvvOdPW8tzr0s2FQHJ6PzPY+3zymGmS9CtYYywUL5tZez28q0bs2xKInFU
gKtbyMK8WFSXSPmzuzOOEx+n1haEIZpVOLDkQum+GuaCRaFobcoJWtGLPyWelX2DIz3OArhjVrNr
LS2ECRIMz06dZrxvzHxAJWGk0CPEbGfx2iHbPyyWbnV1uIffZmIycbHlri5zluB0CKpiXvCXWD0P
FCQVQlKNJjZBinzlf0Ies3uM9ep+ftd/1yAGaE0tQkVjBWDLSUjrojWf83Lx3gKbZuJbXI+6MaOi
V8Jor5Fi3yJHuR41RaYLLssEwMaymXZbTFZjOMIrSWsl64Uk/8RCtO+GxuWoSZiPxsN6K1sK0LB7
g5mN+RKaT6J+kB6es6yoaiSanwZQnAsHzG0Rqfeb7O4QTaO/3XJHA1bqNLwRUbrzsXJAuQppHsvW
v0qaIBKnJk3w7W5ORpVLY9CCWDBwISGWx1j1o9aoRvb0Uk/SMRxEewknG2SJznbZXqvwXF/y4rr9
cGKiwy7XvjcCtMmK4xvs9L+NKnsMrNlT6KzW2+/z7o9nwdR0gCHd+31QSLSMDU7RYz05z+Sr9Jfl
SUhLKBGQ8uvkaPK+cFSo51W0PBwlVYB77cDtCs63KGTvc9EiyaIajw3uu0wQFfWlTNs91SPEiTDg
BoG528kr3+bQSjl60pPL9xJR50r1c4qEBWfBzYKHw7vLSsgeNUzvQDjqUarf1GXR/cRXzY6evD8F
vYGIkG63ZxFfRyog552SKyoYCurW3C8k+9AkAm6yx03y6n6ACb8RZvLbVfzhvVmxVVJjPzjOdcbz
gWJ6G1El50ND4lI3sUnl+W03d1xHH+PNOoDGx186xjfqVoal++pxbR96ZMAJ7nnLwEz6gkIItcYT
2NtlK7MSHsGJySvyvqyj4NSK2x63R0uZeYSOvI8ZsrMNo8QCcCnuGeaUV2706xpTsGWlGsZ5dcpT
hoh6osU5GZbHZbJ35P9LaOhDvWz/mZ9h8HFVWqdRRQbXhK85bLS/B/n3qDoQ+coHb1XaDYt7V/Aa
WlQR4IZK1ibD+LYAyQHl5rMVDUlhN+obOLaZKTzrNOzfCR+VDcwwBL2vcCXCnRrohIs4NH/kaTQW
4DFc8ViIwTpjp7NRB8K0GxZ1YuD6H4lEPdxS3VYyISOyrJRv7fcV7/XK5nwSltFN1mLhskwr77Cm
H8AmSNkqxeRN7msmg9QHMI1S7ooYJ6HwjUxF7ZWqwMYEV9icFFZSHtF5SU2TwmADmqLfEZc3sqvF
9a9qTodGzdrc5WhBCC3hc88ebLD+a1fRBI2DtadcK8yRK4wjgnNS9tJsep1hxphF6ASQyowWtkYQ
LHrBEXGsYS4ti/9ghUY06NS1BPM2BYF/VPjaXgIBJfEGCO1kVRIHamVT9ZrIlgtAplKQm5G7OOTn
jOZE5S5dfxiUaXk+D9HW3lfSSVS3xaopVPQUg06OGN3gx6dXLoY=
`protect end_protected
