XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����������\�Zg�9�z@�����aҞ��_��~�p��n�dZ��pf�m�a��*s��g䭾��/���:�0V��gZF�Z�FȖw�?�����G�����0�O.O���ۥ����&7���Ef�ק����~.Mb���U-&��6E2�}����d�k"�H�a׉�q�d�7�\ �'M���@	�H�.��`0͝'��� ��埳�=ީf�����i(���!���Ħ�%F�y�|w�����"dPK���٪���^�a�e�>dh'��9���U�o\D�2�ZZ��(if���n���-KW�������?s�v`�Q������g����J��Oė��B��@ c!��������W�2��	Pfn9�
C[�c}(��]cb$/9@r��O�Է�HE����dK��������n�/5��w�!��1���e��,��Qq�m|�y�u�ٷ�ӈj:nC=6^��՚E�WzB'�Qaؔ�����OԪxc��j������	[�B��Qao�F`��Ur���g��&�4�)Q�T~�O����̮���-��� �Z�$���
�����R���K�O�]U�*���#��9k��17)=�Cח�����?t��|�l�e�!�iG�P� �`��TPT����С���RTk�_n���>An���ׂ#�L��R��d\�����;�
xم��M/�C�T�NW��,o�O������[��XlxVHYEB     400     1f0�ض�wuE�s";ޣ<��z�����`o6�2��~�]�0h����X-.,WA�uh.���������k�Q�1 #�ɣ�xA:,�U�2T�;��Sj��>�*�,[x���0�
0���� NR��|ܾ��xJ� n��:��a�^�_F�u�]��JY���;0�&���盭]���io[vX�)L�~J�[��܍ͮ�'%��?rI1�3.m�� ��/0>OosXdg����)p���Q��q*fR:���n�������X�M�ۇ^��Vkč�9)��e�{������b�˳徾ax8��\����&����ÔC����#4G��K�2�+�C-�*u���u<�����ȫ�/�FH��B�&�$�7a��;P��>S��q��q��ؖ��X�K��d'��R�$,T�K��[�w�"D�ڽ�����н��&�N�a>f���u{����'��[��s���	�[R�1Ve��R(K�8�����[XlxVHYEB     400     130d�Э13�o��y�7�+Yk�Ya�q�Xw��)-�}��ذ��lhqۻq�z��Bҵ�!�B�M{�qן�r�K>�ߓU���~j���T�|�$I<㶠��p��-S��)T(��D�<WN�ΐu�7�����bW��9�i(S��Jf�\��s�:8���e�K����'�n�"h1'�����M��!�����!U7u�rMc33��Ⱥ��ɣ���qӌV�yїKRN�o��%�~Y&Y�$y.�]o�I5�T�:���ɼ�������>9Ȉԉ\j��+�4g۫;N�H?���`̈lXlxVHYEB     400     120-�A�M��j �O��l�<~#7�y�s��\b�P1����@���>�>�X�_���݈����'(��%�H�/�l����Lr0"$!�_��y;����3���v9B:F����n 7�N�H7.�V:��-y�u<6�����!�z���qyy'��#τ�7y��}LZ�^�����+���Y1X�x�mt�G�x��O�<���J�o='$�bˠ�2$��3C�V�a]3�9�Pb!�|���4�5`���Hv���4i(�nx=�!Th���\�_�7�=^<kD@�����na��C�8�XlxVHYEB     400     130 �k{Q����۬g�s[�p��<��^ � vح��]�D����o���.��St�ҲYi+c�u�I�3J���͆د�VjsD
;�v����%d�)Z���KO�%�ܢ��2B���[l���,��z�|X����\�P3~6��t�}C�Tm��m�"i�j���bn238G0�hZ��l����I8n��`���&���ռb3]rzY��0�X����̜/XLc�&(�ϫp&� CQ�},΄{�0��Fj�3UL�0�h3��9������*"����f��0^�ޒ	ͥ@�U�.%�PXlxVHYEB     400     140 �u������������� ��P"n�`����|D��R^
r��g��]riP�����s��C��*��M��~��u���RUj�~FU�<0%Cl���5nr���O�`�ںr^��:�h���Q܋�=҅�s�ߔ1��/��v��J0V�n����14!PQ�ҮI� ��s�M`l��_�9p��u\@T�5��jñ�z 
�Va�8&��2� ��0�Y�ä5�)�޶��pw{�������9j��B�9����R�D��;�lϗ#���:Q�b�V6�̃�HtI=B/�p?M��	��U#8^b5rZ{,�&M_N��XlxVHYEB     400     180�U�U�@W-��I"MiXݰ�s��v�B�غ��?\Rcr��٦[�����xf9CA�v�G�V�`<�S����bv*v�΀�V��C-8��!@
1�t�*��}����SK:>��tY�MnQ�Y ~/�Crifj1�P��; ��_�V�f�X�]Ua�;�`p�`�{
o�Vӑ���-\�uY�(8D���:�Jm�Mb�I�տan���u%3�i�������;�'�S$K|n K�>����IE�<�I�o{c,T�ݝ8��c8?D�g�� 
Dy�F��)W;�<�/�*֠4vlW5�� $��J��Inv4�=0w��X�@2���St0�
���s�+�o9�Ts���|S�L
�l[�q��gK(XlxVHYEB     400      f0�{D�Ae.j?�p{�E�%�t���EAW/IGxJ��)yx�ѫ�DFf MwT���?�hdlvT����֥�Id��l��������Y�$�cW��J�)�cԠ�jo��n����{��5�]�Cπc���[h�����'qN��E�2��֍xhp�4g/ޗ�T�6�E�m�i���O��8�m�<O���-O��X�w���^M�k�j�)��Yn��*�6��kn�z� ��?����,i���CXXlxVHYEB     400     150���!� ���x� /��E6�Q��s8D�R�sM$R�����V�ƃ�2��UW�s���=�2
v#Pr>��56���]��FOò�֋��1FVl�_`γ�}�o+�{�`�R�@lɺѢpoY�W.)�?^�UT����VԚ[1ȀRX��F7�������T-j�	ʩɊIF
�'|��:q޾C�WL �y�K�Ѥ�(���3#�$�'[�c(:��G�}���,C^�#�m1�&��d\/o���my�E����FMkS�d���-'���eYn��f \�c��h7B�����U�M}H�_�<%"3��R�q��X�\��,/�9XlxVHYEB      b5      70�9ٽA�{�w�$���2�&��@��QAo{y�V.����䷱����a��"Y_Zx��,��-w\LC��==�����I�������uK��g$)V��7YR