`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4176)
`protect data_block
U5CVgTlMlYpkVYxF/RHASDYBZZL6BK0Nl5VuHZbiCiLvIbG8+50Kh2VCxim41Qb5oS5Drhd7pd4R
rhdRkWGB5/TY875XND5mpzVFnBFNfTfaejJLpw6geHWy5cZw/ENSplv+vgOWVAhajGPeTtmOdlCQ
YQkHclnlH2WqGgsZwbQTd/SZxS+n6MCqeR4W2vOKL033dy4jftUye/cQx9FkI/Rqv8YLIH8dqPhH
Q8xowxe4BIboPUMxFOZaPdPfrOdHZ6hygzsUMTKf2ez4Q6aenv3D3aoqioQdHD779gYKRFdn6ySw
fQTq9yMc4ehdf7P464sBLcFa5hj5cxwxXwiQuLZ0ZOuzIDIgjEkqgCMcDzBeZ17iTds0AJgiPWIB
jdJfndCbF8P2gkBTPlWF9vjpBgHNVG4ZDFe/U2fR0e1CEP7g/dodixZO3NR2BuethquBE8ssQNga
xV76ElX9d38V09TiIbLbihIgdOXQ4bKYmPR0W4Q7nrlv3M6KtkshYOYvJzVYsQnvwuKKKrOVl6ft
ub4YseM0qVaSoMkLw7xfGLNRqZJo1mNUr78KS3kIsCcont26tntSihm5APL0MRaTWYhUJnnoUbne
HbbSHCHGDf/uiwhv/F/o0FfqFkVSCGhqjCQvhC9GZhUofb3riOStQPYbNC0PHIFl1aIsqkxUphjJ
zCXwrEsJ7XYNSIWkeSFuyuf6H45F15EQIeTap304Ew0go/aIf96pjFrtF7I9AwsfRDk+9bMMVEyf
hzQPkuf0Sjg1wcpFZ3fpU6xnkhM9snJ2g4QCimFGa0z1HzTTppb74DUb9kYesodKTR/YxQ46r8jM
wLARbK1zzwYZVLPCrXT/WSYQ/47wXAP34q8xikSqDhtDC2Y4EBTQAU7h0n8Ehc2budxrPpZoiehr
kHV/VlJELhwaV2eSbC/AVQgk5mbatGA87tkr1Ua4Of6a+IjMBsPO8XCzolhk8AW//W8ypXsJzD0n
5oMiBU1asVL2Z10peTvOiDJoCDOsro9y36EJ+dlW2HnLftZccuBroB796wVEKNKxatobiz6cXndG
qY0MNNQtcstPasLweQg2i166JCH7/Tcuuda5WHUf4Agiyh2IIf0PuZV+JJpCEcu+fdx5TRdkmf/4
paZL5s5JBib3o9fQ90lkzPdFf7ppULxSQPoBrBa/09q2UTuUAK6KHixV5aGP/olslbuWombi2DOF
8LXrWqmHkhww4TtVc0oZEH/TX2VroY1Dm5rbqnzYTQaAvpJkJT5g34+a7DZBxXkJOCwCLCi4hqYY
AENNp6BEQsp+MYsSs38cRknipm/VmvhMTsNanngZl0h1nVXFkuU3+gPm6/CfRcs/Tj89ii8kvmQW
vHgSadYWqZBBM2WMSPcEfsz8+4s9MRZTo8DJ0YGRWmuLclIO22V+lcV91iFfozYJscGqNxdTN/6m
wFjfhnHp9ZClaRFXNcj9h/jKujIuaOqete+l0R9ZjGRe8XWye14bN6rfMcyhGRxcNf3Urm9HY/Q9
2M0qPFADF2Q2oAJifjnIerlIVlaGSOH6JpsXmmIcGlBbqnQeKwbA7eafONsiM7gXtKrMyuQ9kMsy
BlAe0bV9e0prlowiC8EydQisQQPtO6IHPPj6pqeyXz5GM87xylOtZy16f71DjCf2zfdI3FB4f5mB
ZP2A3Sdzd9BL3Z3w4ifIgADDPustzwuG3xvK2P7S5IjAk1miyOpPuh2419wyEuYArwtzdPHcR+Gy
mxpVN/FAvRayaQm4Kb79UeMkOkUhI28xkZDAUxY8swXemXaiQOwAVieUiSoqi6Ok1l4+TXZmDCzm
eI8PJuEaH14ZB9Sgq2/h1f36zQN7LTE8c3TVrUqgMINVolRpc6ZsfguDBxRVeFDdpvOH6Ddd0Hg6
v0GwCPIL/4caS4TuJ0+N+psfGu3QMrryfYnnxZtgFiPjGTg4J96tOYSgSBAHUMXDKMwjfyovampJ
e/zJCpCp28s2q2slj1rxGe0dpQwrrqL4a1iNhDqxOSbk8QSXQ5hUt0Eeh7fTJ8QJ821YzUFbbNzm
QvKx96jDXnOZUtOuIrRF0N/RQvKiqiwx0c8T58Bc3O0lSaaBuz9RHGgbdpGsPgfMSE0yeXaJhBVk
HKdq+yb0uIDBHNcpcZDOO/XRRkrdfyEXaAYoIGQhE3OdGWiaJ5vPp6jOYR2Jcl0QCuz3bt82wZL5
DV5eDV1trwqDd2bcMMuQTWqJMS1MMpwUKSxOdCZ2X/QZJwDhh0OsustWyahES9sKKqe6DbNNKwWc
9xw+1kwLhuETkSrEUzcqJHfujByY0iLXxR7EXckkCxiDw8yZ8KofM/NLjIqJkPlnrPh+xwK7f3ym
MgZM2bzy7RXsn345z+Za2Q/ydteAqxveoJWueRC0jNN8Coph9nuoTX+yMF0uDVqbkpaX5fGNUvpi
Da2/CLbqsfHwDhhxWTG3yrz7762rMhOxprU7jfsgQp9lPYtSwnX68+6DtlcqzYVj8/StKpfMowW6
cLK0VWyMCKWmOtRFrKlqdoj2q3I51xEWRuW3mcAzabQJzQ4C9Lb/IraQclL/o27ADX/1VQQeLpph
5+HsUboNsn4vr6z/y+2sMPeu+a2uL1QbbhHmNAohgOZSquCPSjo/4m/jf00l4TYpqjlfXTyy+iZz
OGIT8vj3NhpuAUiA8fx6RychWFW7PNk9Fk7HoW4uT6p9xaSXo/kwUa428dAN/N/3KKwOtsEouzTW
JJZk2+RRVKlJRzgiqImUs1G3c01NslqMuzejC5eImyqgvdPFkJZMnm1qNkXnFUrx3NGgZBU94dnM
Sc92gaKU6uH7qck9p6xfrooWLg7Z1h2UX+nwhPnQqrbwEZGijs80PcAYceMFQqZvhne9C/KZeOhv
6LzY/LGX0bLqK0qXxqVvXQP1lSalyojI9nQMqE3NW+ZpDGsNCRzj9lNERAqBc1+O6Gr+ZrAOMgPu
F5QibpP7oLoBBimA8DupBJSH3c2inXeyJCCKSzbEW78ahyoikF172Y+XEyflL0HmdqIezZjvcUYI
m03VJE2B/FL1pQDVIsZcQ3UvLd0wuULTBIlsjoghCqSAzIGzevke5wSpQRsWp3FpXfRNTnKcIxdT
CEvtR2IGcCz3Y8HEU3ileAdGcpwgP0vhcw2Svtn2QNmDkJWM/xmz4AYh/87UviM9kdAL0ynIgUb8
rTtZzUX6NB6yCg0eokmve9CdZAnrmZ3oqKONQvLdKcqc4iPGFG6ZkCSTDeLliMs2OEXlJpEFD+Dr
4tJYuuLpSBVsytTjQdAecALY6cQNQzkhCaIr51mM2pEY70VIrC0scmx7VzqOiQdttfrLbMK/9s/m
gcv0ka7ZXpXcVIg1Ib2G05/fckRqFThEr5zcte4cPkPOYaoW++0WEyyb3qoVXFHLroQm7AZckywR
PtLNXIk6+ivHZQRrVSEgzs3f3HOTIvnh5OJzil7UW/MDAsf9g0GPEDU+OaU30GhOFl4cNMv3XTCH
04GzIN/nzFQrEF/tP+uWiZy+dXyNBNCk86RcOsDNwKtSnD8xDwJR9nsLuM+QLTaTIy7xCkqWyL4Q
7C8NnenHGxm+QkcsCqKpvtij5J8nm0fmYLkn7eO+XoTY6IYa0ZTFNYW+8GJAf+HzLOYsnOUlPC0P
DUwQj9oPmA5dOyHxUGAARjM8Ip0vUTlPB/hDl4V/RDkuJ6gwzyk1JUd+iOJyML4jif3c2oH0Wqzt
t6wFSQifpWWH+bmJBTuOPWw2ZCoGyuIw8bY0OzEmizt1KIZtXuHXGqsSVxvzaXKGjhMV4vXdw1AE
houd+0qGdZ+UePXoP6vf0u/UOCQEbiHLJ8K9InzrVBNiCn857uzSeoU40iBaczMrlRPUuBYZ+DLe
wvAuliku+ZxhdIdwgLaBmUHleB1OPd2KfwLxawLStvFQPjzab2QvNL0VO0FrxHxXOXD6nMIiagg9
nD1vKNxFSdwYwDu6NT/iqMO5/9GlY/goON8crNW7YQM9KARYJaUt6LLgNKz6Pg2neCe9c0HYYyGk
Fr+ItbBhQC+sO0MjGrQ6HULrGEvnkmJNzRCjOuggnCOna5OGnE/vikXS1RfcbeWlBUbopOi+Lu7H
muVHxfSu7eMs/LP4tt+BcmqekWLwplnq6PsG8IREekUtY4m7+qPiIKM5lJPtAGrTiQyhfceSh1fW
rFW7ZXrqLPrLCJFRyM0ra/2vVZagO7RHDfzbM1S5o/MPlNN1/E/uhviJj+oA6N8o4aVWE0kyiF+/
7aE0TxRKXbRGYujJ1trKWh6hCUwUzljQ8MSvxjEFEgQiSpaaSwwG8jPKAgys+PrF6XQFKCwQGMgd
KZ3dy+G1spYfsLxcu1qrT4lxItLrhzA20YyyqP+PSlLpBrjYlgcdx3HiWdK0tEriKTETeF0hC0aB
Bie+Of0L8FJMGUnfdU2vtfuDxrXzg6D6FoL6lzcELTIRENQH8ZaSIkLJpk+ZUovK5ghZzv4hLXaC
Y3sBul8kE8KfCueOKgQDipdaobAtGQdR8eBPUuOPloumomuT9TAvFZi5SQxzLbC+nAAMB9pCc2Tb
Z7pb6AeIwhHkNqzvKMA8TP6wjppRxxEJGPWt5HDn5Rx5+zI00zlPw7I6kV+EHSq67TcmLkYzxZgl
9raI3Tvyh4ZZvaP8xXImmDtsFvYZu3XDF888jp4dCpWy2t7PCT0ZylrPUmBkdTj9B8+zX+72cg5r
MOsPSWoxD8n+ndI3WHTbrBTgnyNFz62arZXGbLuzT9eDsBkWzBwsR9ONGRb/LPa2hospSMlul8at
9jqDHnEHocAqKEdAd1VF/ga9ZRQYlI2q+DBLIOnQwElEtvvifix6iWHM34Thsl9PK7VVxsfKBx4r
n3PxgScdc4++T735A1/m0mhAPwchkhEP/1leAacdMwGgCTn/p0NF1aCL0bEUxcilb0exD03aoWTg
MHMv/Z9xHV/5lAsH1fFFKg+YN4qvSxHqcHAZcMi/CEerIotSQlGYYn0gYqPDxLhXS8ZlOKBz6KT4
+Sl/1G6KK5FUsCMQ40EErg09t8ma7I/Smk/7qsL8uahmplRLOZzMviXiPPrQxgaZeLb9tVzRUVkM
BVZDd3r70hIwaX6vQtU9cOyTDnMjbT393BGe2kvwamdW929ZakD5NAtI3vj2krGVrwt8jDhesVRJ
852KVicsgRXbcmnAKkKOpLrLugRRppR/IU0CeQY9PBJ42b30K6vXdSVbwbLHKsp3wQ3WsUK//OSP
Snb/dGMm1wNYoqjVlCgayL3GGkHwdTw8uNovl3M65Bfv3j+82YQoNxztPUJnkXlITSKLW8TpuZcJ
q+sOAhVtYUFNM96ZFK9kJ8aZReeXgGMptDvyoYUKBLW67TjQkC4pTX5/mtNti9QoJXMHl2GpvvXc
CInOvl8c17q2whQILqrbnnQ6d1kA+wnEQV4d4cZNL8ubarkLCKLpiSyb4EXrnsfOUUEM7wYgdJ0E
jOraH6tAoThkG5CFcYdc7jI2JUQSQyUP1SwBS1CK+2Cu6WEWaSF/UASag8FwYzWRW54rEzhXTRrC
XfDT9sHhCKfOFrMuSXaO
`protect end_protected
