`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13920)
`protect data_block
pkoG9Uelq+Ny9Bi4J5egQtwb0a8FT83xlJQWwUtJxjbBPg9kaNA7BepTPRvlC2Hy0lYkboWQtxiH
CDhgbL2qD6TnFK3h/fdtyaoY4OIeTXsE7zjYvXixOcrwcB9+m1v+D02PxHbeLZYYeViO32XLLeOJ
GgBoPOwU7pLTlDlq4E42B8+p2WkNmLGVS+gYWuFgpukdn0BCdy79tNxHDEuCG6pEo6IhOsAzip85
0SGEooaSAqJIk2kTqTFC9MfRZK2i0h7c0eMJ4m5VjyyfgcBYN+6qKBiMngkK3f0fFYouJw0srNF5
gSUSnU1MaTVcUNHp9UcUyndG4M6Go61oDzAD+f+yZd+BINJZMMkLIIMgrJ3gNBzq2qy27G8yp9Ay
XpqI3UxF7G74IbG72dsTEDOe25dlmpd6zFaK+9r7bYJCc4GJ2pIjZUlDvyAFImCLrn8uztwJLptY
6MWp21Tz6SNxbWxJ6CCZRuycegJezxCj2gJyYPyftbY07iAXaHVyQkWXJxstV8w4wFpJDSfHM3cj
cNsfCSZrEmE6FY2ybwSVq668Yt12S0DO43aAL3rpR/aF0qsAa01IGH/icB+6VS1zbps5h9wfaFC8
QCnAPY+f+BMCjGHmG++EJd2eR75yin32hRFHgK1ld7+sx5CHKPSBxVVj0j0iccyOXs6atg5XyQXQ
MdBaZDjyBt7lxHAIdrV8EiXrhKvUmiIBRhceKILjBjkTFvJGMM/VL0gIWkWc5APLIadqbaulIMHB
++sgf5GascRrUkbdHkjN5LAvNt+BYZ7H37lQk2b2D+0+PLPf1gLEJoehTmOA56r42zpN5gfyXamB
ooScm+pgoTWXzCHTc1mtaMVeAFhGubTqEiYLQ+TOrWlHyKwvBO/EJuhJNvLyqdYiAMmnFuz12GM/
viKFGMVAQDtNdxta4h4k/yu2gbdwUOaoI0Gb3nTnqdkyjceOE1WCtp/0AEJX8HhuzzBWqFSOdmbT
Y7nF2homB9LtiAaZi3aWmdvFcvG5WeAsQyL7yJ0cWJQgY/Cmrs1WfLO4D48HSboj0aAwMgD3lIAK
h+KNJvbD0/S9gi5oH6fO1fBxfa3hKW7j7m+/DEX3UXHCKBoYAjcchbsCWouYDkRg3YgIv0Oh56PN
oY41mlvgPQO8wAsw0FW8llQDX8EshiVZ8YvWa8qxnpY1c2DbE8s22LCrEayNCBmnZ888oL5f76ca
jA53CEkTCBVsmVvQit5dlGIz3hQF8dhhes9qtXrw5HoIWtODd0A5tVI43eJ3KZLA8zfQZp0cryum
1QFscUs+xA1/Cd6uOyZvSdKAIqaPocCkpoaydZ/K72M551DTPu90EEw8kUypYjnXab1hTuTMq1EU
SuwKBFq611OnSY0Wz5SUyMtSmt1VqYWeju028l7h7KuV3p/6pwJGac6+l6divNiANlrkHwKagPxV
Co60CH281t77WFAjzMzgwUauDSvqB9S4OVIYeveEK1sSwUOu0l1pzuEhsu+xEhumyQUCZqJ7c5tA
s+qOhs2rEN17PNHzu9OQce0toGvtSm9wkWXXSnqUfUCbS7ZG3i1vCSP9o2jqLW7LEvB2C5L9CIoR
5y1UCq15JxHcYETzd6vk0GQUE+UaV6Q+2xOoD5bmN6L24qRWm4LqkSAO0MYEmZFzO/hxuFag1e7J
AFOrMRgiXoQpW7nOG49lDF1KGR+q3GDk6FYMvUcotZ3QK6zwj9kGOkEtd1WJFbmk9wuHfV9bRwRb
2NP6Ut3xyC12xO8b9qckuqZAxv7vUO9KZ1dg5YU0bqLcBjGPsQVs3Wv1alicg3LHdq5wFl4PxBim
h94a+wbhnvSUpb02TBs2P2Mu57pSZRLS4Na5TGjY9tmASU7QaNvqtyfw/k3Azc/2sxhtnI0r8XyZ
yLKs/SgZWbKkmb6yIDOCne1XFKqSlYSi7TOuMQRPLpYZrGENqVNc0JXgLUowjwPvR/FigESIndE5
GXGiWPMXy6d8VYBr4ocOMGRZxR8GEUTE7jwAQG395bbBfhDr6ejvR4U25JIFRMvhhsYuSl8Hr1k+
cF++ReQbVdRxdUHIAIzNV+o/XKRnCSJrwPL/x4j8T6OvKfP1Rm59fsFKGSCn8YjwY4kL62AgWCos
1194F5n+spz/Nzh/yoApWWhVmQckdF9dZhFavX3r7zgJe8uZmtUpUTnkcvR8rMnlkpNhTjIl50Ur
Gd8xrMauSotPD8bGXVqqSDe1DbI0VYNLfMXodHlzLVrE4qEqI7wj9Mx7vofXbMKINo0LH+gzJSi4
eEU3p+3GIyAFLvkom5+7C+Xer9hGMVJSv71+cXvfLxeO6D8+xQsDBarPijlkMs7yEdwIA7UN5Dq8
a8PlEKssf2+Nij9j7VnvsYmc7WEpXi2UDl0C7I+Qt0tqAyNXIOwAXK2MCzg3/d60fceLRkEug507
hYiCUcYJOppnIqv8B0wJdt9kW26OoR3DwJ/JqLtTTyoI2hnb61Otn6C9B1iVnDovnTwq1yh3gaSO
vdMyqtiabYwpD0PDzo0XHSMFFQsoMnH0+sRizI0Raf2Aly8NwX1oQNMxhLy/wqa/BWrhg55LhVw2
fojSclaI6YZK/ddkMsEaaYms2ukuJkU/w0ZbUawwcpsEMwEAvI+oCDU+aOklpjB5qzvQXAattC1h
2qCFOw90kZoVK5xpo0PcLbQ09Tm+gkUklO476LI0HoKTBRucO7w4k/X1x68JPtKpU8nas66QbZhH
vn0DHfFZ1HpsRaKECB6aleu7c9YX+8tQMCyOVqW6Eq4583AajF+IL13ijQqas+CjYohzzPH9UmM6
/BREfSpviTZMvp8c2UOC7d/ngkrkeVYo3ka/KjsbeMHDPU0j2qkOnJ8n5SENO8r5Ii7tao7cdg/i
qvTInNUAZMr/jL3NUY2gvpOPUHbznspTfhB1I67VDEyttBX68GFkUnen5rlKSTwgkGQ423swPE8s
/xc0FpPq+DapJCjC+j9f6sqMsHxKOKa4rkLUOxUOK/brBva2Uy//26YE4MB0X03KKZuQvhes/Ly2
w3jhNWef6VTS57gmpkRIaQ9aB23Fk00osJryEc2Iu4TQD7182Y0i9Rkqy/feM2N8G6NCqTpvF7n0
corL3N3ZtFr8rKUXtASbTy18RNmWNVtkgj+pqVfkG+zcGmby00PxVut3dmx3jyM+OTYb/cgJu/u4
tZwRRSh5LhWYgmbNN5yG2sOAJ89vqy7ep8h62kj131kY1BdydmfsIBVI6u8a8MiRL9tJFigE8TAf
6OK+PNCzf0+3WEU5nsABLAK6OvDiNsnuDEA5r81d+QdVAiDTiEeJDYORZdNckuJ7sUhLU2jvSVK+
5OKrW9sxIevDjBIpSij5w5wu+yGR9iKs6ZNVYLv9R/24WOm0XN7cQ/75UjNUq0JVxlHa6b/qmj4/
6IUdq3ILDT15EyKri4/K+2/HCfncwdyZEKn3iKtr9NzKsKwkXKGUiPyd0gUjCkQ/28EczruSX5dO
LsPU7r9QREnIZuoQ7tgQgKBghMlwb6+mMNvyLXLbE1e90ym/53KTQuBj1wHIWOMgs5KKzeonDASV
yFeXM2Mx5i9JnFxf7Oh2APz11dY0U46ExYL5VZtwKHnyPjzZGGZ7R5VANZ1+uqooS3dwWDv5ufOJ
HHeU1Q6L9mbJ6NOBDQKmfEqkOEE4Jk4WTm1F90Z4uoConzWz4jy05HhqPdMIV3naR10Hm1Xis0xI
+ZXJOLugdELDRfcgdsocFhtoMgzoQbSvOQg4pHTp6wYyGuLnQ5Cy06nQy/4waQSc4RKfPZ6W9Sc9
ORCKLja8bOYajeY01NDxJeVQ9chFb2pROi9y8eJH9qsCLxMhJGgzi4vdbZ0g8U0rCmnGngZ2HDSv
DN67BMFWHyVqsv+BeBWAuEKCavHR3xXRSnSGvMysH0Dnm9OcmmRnTjfJwiUatHPrJsIgnD+zNqUl
gr1e48DB5BQCRFOxQONEkawGlHclVFrQsLyQbwcWJg/Fmr90HerOJ6cHyXU+9l5AXSzAmPjHCY9R
nWPlGrE2QsRzzrncWjhfRpqRcQGKm7mx6RvfTRH1CqrCU0LRsynlMqZvCqUEhxgCgL4q3iAie4tJ
CXZ3vBIvUzMlz1sBbZaTjecvRJxA6EihN41Faa9ugMrs4HdJ0ymGPATqoW7zcDGJq10S4QtXcdZF
2CUQRkz2tuA0uCKi8fYOXW+atko5NsvycKwtdpmM5FZyzL4VAtTid71VTiK6JSsGR5TCicLHdCgk
ESbadkiI21HiNwLzBz5DcxPubXljkpJ+xdFv8AhFNOlL31Um6XIqNf0MuvfU5X9WnXcteovylDRK
KkvkRW05h78nNey1Nhk03GxDqpvlLSDmvAu+qPr49t5z5wYxxXFWOQ7X2k6I8Pmwjy5gf1FwfkDV
xyFHLfCqd/WDKq2rSloCmTZSLl9iKvSN5FzJbdblkT96yZHzJX+J5jWz24FPwTzcahAZXcMY/DWM
t1NYP06cwKcqjRzlM1OArOawptdv1/i1BzC4AeOXAVGdd/L2qm/VuASdg2+ND7+cPuc9jOMYws7I
EdFrk9CGOsxjLUwYZ4dee2pPR3VaXeI5tR9g3y6OOwh+aM1iszD2c72InxB9lpbani+89OBgXd2a
BfZ6o0LU0YfkTUxl3Qqc8OiUFVZnu52FSuBgREtbFzXE6LSR4f6E6wQsXh9DOhb9l4Xb777Qb3gC
yGvVJ8seSNC7uQiF8TEvRqHtb2puCi7qaaCB/OSC41D4/7bsFCcGN66T+R4CxgB6p6BBqemM2Viq
2CzRtyW6HtJuaa6Y3LYFqp1BdCXh0vjK7kQ0w8pd/PS7X4NrylRA0BEmDWoHQS/QOiY8X5hishq6
d5nJgofJd/1Rw69vZn5O79DMpmdeUkD/iWoOyfJ1GWBybusL3H43VIbcARHtHpmJ1BUJVlwLQry2
6G9cPSyh9raTeDz/4KgaHIU41/Sx9ZEhbjtByDgHOEla3CiI/ArQ9mX75cYl//aaDO8bhKe03Cyo
K9ftwANf6HWAqDGSmnwmeYHGgbufPYWvfra6w293ROjJAga1LuTkCz0gudZv/si2plg5pFB5VGm7
4KgpcKGvulp8WpzhnmxVkhAasAwqd3simtegPKAcVTnXAp6FRparg1kG/XhqGcK7ZtfDqZ4YJLtC
+k+ZWw1v90JRqQy7938Jne/arluNgcSs2MO7f72lDCgcWkTmjgxu2yumu7pREpFnZlIv62AET74m
mV0HIKeTEPRu1QYPZsG+p/OciWvkoO0C+kQrvvuv33HJqNO+mfgnt7KYuvlV1o6VKVyFfUYKmg1Z
wt7DSOoqb4u698v9k6TL+WDqgq4qw5mmG/SJS2eTx6muZim9gSLL6bHUfPae+HN8GpOPM9DSSHM4
2V13j3ybwSs5zsm+Tu/2wCXR7CXhGxyYFiYCiJXpfaUFIxWmM+YBNQXgG3WzuPOuQBpnFXTRbrKd
JVrQ8AN4V8xLQG9tbe0luG3CQ2rXRBnPLfyNGes5YXA2bhbeO2Rn64q/bIov3oB4Ayl1Y/EYcum6
KeYgJ5BEk2V3gZqcICc6u2p4uMXGu9QmRyreW2S24EXLd6ARZGaDx7tt03c3HqV3LYDdyWCcYlrk
0twKu+hPLHIvY80o4qpCGhXS3ocoUwdqU+ZkD2Ng94Ja5U9YAQDg3dLaHjVqz2y4/ej+FcNq6Y6d
WRcaa+sS6kA20LhXFW+devpUoL5QpTvZuc3f0QaCUqV/zYS0C8NcAGiJ6JY9toQfRyHZxiWw2mAK
4OtaGebGC2nxOBdRxLN/1CrKGKaj7dXB/iZ8tgFp7lJ5sJO2dj4uluxl+v8ieJtLW0lf09KFEUms
oRsI4q7w/vRi1+1jQK+l79HJssLlgoE9BVl87BLpxM71Ch0+AV3OG9R6I8Eg9nHSMNCELT77E3Kk
k2mBqeqziAS2I4oOPs0MyEGByEbRuuCIasRUVhnPfG2GNzadZwakWBQ+RoGTzLIvKVRBFohqJjf8
JkqNfOGi6M1uDV4aOMLuF2bM4p4YYQjqbQhAfzwBjleuzhLF7FjnTCAXxdRr4Zk3uur8EQmcIMhG
mUHdVCsK6Qd/vnRFVJuVD7d7Uv1dStyJntY3cGKCxWrHaxMVu6VBaZ8GJYnJYEFcFQXk7nNRNKUY
mexTDS3rJrYF64cAVxkHprooxJ3BpfyvG7I5W9hkgitCGfNBXesqSrkhNLEOPP/S8rHrV4tjusQv
0f+vS0dKNUCBe6ycY9MJAUpsOlVaI7eO8K8f0Y3erap04T8UxH1uwNhXCJQES5yebh7X4vljIjaP
dT9JI6irlAH6gwIiGCx5/tw/JRDnboNcI4Ke6Xx8ZeJY6/9Lf1/StWxGXQZ/iD3RcjGLUTm3thuB
8UrDoTdQIg8hMstMSAtPLzqH2eAuTE8Ns57AngoKpw6gJhLGNHJ6mZ686icad/t1w5kIN56bd2I5
0OqOhdeGqHI4kAbmFyVUe1IwjG+EibpfE2Bo+wNmyP0Rq7iWPaMrD4zKHHdj3pX4AYwu7TXtN1zE
snLtnjmTvrkhjYoUVmTA46klY2SOg04+CM5zRvpiFl5hMPmxi+0txzKHPSpRZDu4cCEq3plFLwMg
oMGV3/W2i9Q6ZbvxroLBdTf5giUtVMiVC9qUfotPYIaW/FXOpOF9y+OPFbePnjVR/FhCOR7Oi6cO
o4o0skVkl2Tmi/r1Kp6TBLgVnLQp6tKG+feFjNbW12vSl7Td1JVHIcy3rZ3xeVG0SFcjAD0Kh/Uh
TwrsH+hgJEqE0ebdByjqPsOOC38vGf+gu0usAq3FsCWrRlNbWuGI11amlpHwqKH3cTcV8m+z9WFG
zyCzYzQXFwyH9cm7EHaWpd1Grl9BNh2EsO98oZoIzlwxg47RcpFI/gwGTi6hfh6ol1wRZlczHBwC
GuhhDFXL1ewCnF8ln0Tpsc6O3YXXIK4jyKJPJr0JfS2nbMh7FOeIW61n19fN/1UQAf9MYRBZKuvu
GNhzWlLeOY4/FrJQXP+Sl1lOznBHpfN1WTVb0+TNhseZ4/X57E2QkIEjdf20XUj5an03UZ5MitSI
s2VWUzzHS0LdoD+75muevc+L2xO+CSlK9vL4ASkJ/FRF6CZw+jdv5oyWY2iau5uLhRGGwqO3zs3z
t7Y9j1SsaXRRkyj+WYGa46+7jJWyMMRoTCGZBfDRV8kci0snwgaxbuHhgcYwcWTHK8/laXbKOTHV
2yXRtNZ39LVY9KWMcUV13iDqUC8EVgGEv/QgWirDgiiL/tQAedjPGo3epRSnRvRSCD4liKoZMPEw
nZc6fL3NMHVDZGn5Sdxpn9bnV7+glGC6RlQLhjube1191qahP+lQQj4lgErfjJ0wl+4/UzDBZt52
cJVMpDjYdkBRlbRTMlIHcqjNRjOmY4pSYbfD3RMeINfjRwkCZLKEVQ3KWtgLqC3LyEIWU0QhQfWu
fco/zgl522JjAZBw8JR9yPbG0X35FB0MUgYK5qCLcmVLieitRs9szG6HX+bD6x1/YHtNlFN4Kx2G
GjoE24SWHSSeVccjsBsvZUp/iu9Ejesu7ekyQZSrMqZF++5jRPgcG82HuRoGo3Wa97HD75hmp2ac
vnffONDjiasCqbnDDugQXxfP/1oxBxHUzzB/zBDLGVqev08npAYDR+JuPyQHuxc0tX1VADq5rhJo
KHMTY8JBkSxdO49G/li95UcxojjWEwZpmEjn7rqh9o6L7c4Cf1ik6rMseTo/Avdyribu87vRIvBY
PqEz1iYfV7TWoLWv//LKCgOm9uC5QXbdCp4VkbnLJgWQWrCa5S6MGi9Hqn+RpNf4rpVYnDUvzBOv
SaLtgLaos2zKe1NElvGKt9AyUfMb64LfLBPj+GpY+GWHg/tXiI0oeRDQ3vNUqo1U044Se0IrbKh/
FExGnPVW/JfaLHdaTJx8O7EHWjtkG2rygJcW/himmxG88lJTyxL2T5WwosDdzf4P9FCVA7s6MbNu
3CmnZEhVwv3EZ/6HYR5FA9fRnBLJFhJGvkzyXLlzJeqs+tdJVJWrQsfMrnaR+BWibkaiKhlqLHHD
c/TL2qaCBePXwkNyst7gLimRs7c+oLoUpYg64pP3LOyHlTza1qxZCwNYBpDoL0jAcaWRHygHNJ+c
ryn3g6xy9cTdX3vNgKuLhQnWYImkf2CdPOWbUAuGjrKf5ibGwpf05Y2obiT3G57vD5/IfirEuXrp
z5O7q+qT10I1tLnCpBBNMyijk6JziEzWylzTmEuNGj01XnlbAvAvttrk0CAypC22eINOJB20YMbY
b2Clk/6g+fPSVn8hqoIcwTNOhXny0H4ad67fcXTxbQirAj4hJCeHFH6o4Z2G1w7WdG8+j6XIZLsz
UnJMCYLnyHDDhUKLytaGwBMhQIHwxiMv5N9N0zBtbbEErR855Bf/QIm73XvMuTOmiyaGoz3xec2T
rDGDen3mlS683pBtaTYpxTNqRzmUuPvQoScBpkqlBNNDv1UZxhLxTfmcMBgET4z+VhPIPx0io+c6
0YCslhI6vpSjNZ/5M5EBMkfjwaDMY3JBnzLzcVUhyN2kwh+/1jPhLrHTQqnneh49kc+KFVM8+h8S
fB81WQ5stBXsQvFxvSvPm2MwBx4gbfFRxUF3gti5ETmgq8jYXClbUga2CiSXBBhD6eVfNeGlsDa0
n7G/w4U87FjZ5VNaaW//bKa7f1CAReaGKdFWrLVeST+aq6hQFPoegegUcySfI4nzYvqp/c11k0Bz
3fzqzzXfuY5igHxK4x2VSR76WRidKw5RwUbODK7Q6gr/SrcTZjMFrM2A9w2oAwOm2tiwMxIGKlcX
YaqTrSOPUT4/NMot0DaSYi9htvB8stcj1UemmDHJCGXc1GkK/H2HK//iVGG8i0var7MnMus233cc
9kMaM/1goNovSuxPULq07fYINLfjsYo0IJWKGfcN82tdqvi/D/k5Oa8JXKPLdTz7JfyX6bJa3OWx
6dSXX9VgIe23JYXw6JK5VdNlwNKEkdmtPCuBENB9G9auBVJ7XtYrBFB0i0UpSEthWqsjgCDs3Rwy
jHCnBE3JrrAoCE69RIcewwZnaFk3nPNhn3Sji4MpgEPyNWb0Bf+KhA9IkDJKnToKKPDz98l8ecAh
Z8gpGJ+UA6Pm3Bv04HHg4sRrPz63PV7biyBX9MV6rvZHYmlsp+lT8E1oL23iSZW9nCY1zg/6aoz0
YQ+6nhevT6JkeOpWwWkJREIPFXJ70dyeCQ3D76zxzKwIp1AqeAirKOL5jA6jsgpzZ43+frMqLGk+
1mDJdQEGy7bawGmAhMIEuaE0GuBj1max8VcMBmr20Z0krW4Wfl2WX93TBVrzFKg6+gR7AEWiVnWh
NH0854oZxlK3r0qYSRTCZ5ThlBv5OwJW56evTPKryIUGPGBFBPo02pSkCb/hegQU9PeWAmgbN7Wb
rJ+YyPXwYUuG2uMAbbJhjrEMHhywBBP4VEe4kuCEEMnFRrZ0coYfOZ4VsExPuIdpud/7LO49qS3l
JwIK00JLiCn8EF8XzuD+DuZ7l43Y6sojuh0Nfs1yGzcS3zBrYfcIphddYjJoFP9tDpbMg1fTRQy0
vWhlqoJCgxHDiRt1EHI9HuPVMD/IfBzXKWHCgZdPnyq4YSDOyUaJ9XpnjqYzt6rqaPtTNP7DfW8g
1pszi+TrPxPFqxTpkBbX4NAUk1MU3rQdFy74duYQWVk5rrB6m/nU6uGaRpImRbtq8MiSDjiX+4/x
V5eVn9wWZXR6c/s+FQYvNLGI/NN4jJyAe3bbK0+x/bP9K/vHhFrstP4QfFBJD2iQHfe6Vk/zykCJ
VqfRCw4f8MlvjnlkViOyhu3xiIx9SdfIp3Ml/C/oWGfhSvrLfDTS5VEbGvIoSui3lbFi4qQYVFAd
Z6Zz+bY9Lt4zA+jQ92r/nWJQ3clrYnbtd9amYi5LU0U6ieL+XPqgTBx/9KKPgdCLo+fPKKE2PgeJ
VFqyreQAuMaemT2ERcjIaHUEMu7AO6jO8xMR/LyvRFRpGogk27QavP9KeSVqHapIkqMGb9FxOguQ
1+bdiPX1FixjWYWRy4kmUuESPoaX7iC7fSAu6z/qYahOaWiiZdPjOAC2/znSfBGOfQtHIVWKY8HS
TuMK4IP6DWZt95x80aEZUIqdpsXF/xujlT67aBipnw04Fb5TSH0uEPex2SAgmFZBienan/IlIsGr
O4jxmVwldOxKzIQkVdJZMZGz9NEVkPsn/8OIh7EYP9pEjJy8Al470FD/LgptRFKB+iY0/Axh4Hso
PMX0p1h8AUENdeyRzymVd7tDdG7Pk4IqBIao0WKTX2PLtQ4KKrGZoAFEhVcTIBw2Or7+amI8f3wN
mfTuXh3hMhwuGE4jcLcVn2SkKEP+Xl+J7g8zegEqkJ9CzXC3J8Ff0G25U7XaEsd+QunLwWeSE8Xx
f929NNLXgE4qCd/4iIAZtUKWqcb8ovGTp89en4pR4T037khj5ABZ6C+qNl/X3tKt1dkh+Qot0/r/
nGFlHh/7vKUk27L37Maz2q7Pu35iYHZ+RQKdfbgTjYJd2Ytkbldxfgt+dd9njhIA3sYzUZMZVh2Q
DyC36KijHP2xVB7k6EqezCWQeu8glu8Esav6hRE3AEbTxUEQxvwbqw793R9nu/LT2999GyGzK+W7
GgzXiUvrt25m7xGxLVhcUWrMqzOGUJklQVrgovH739NmBn3+wRcr8AXdbRj0zQpbqWskwNYi2PPU
fcjk5oJqoQoFmbumiMV/y0SxtY2Y/H/ogrAZ8qz8vDRLp9KYovoHgXlZozaxzb0wOC2nX+CHhFWv
NzR2iCtp4TT/w84dX5PyYrdHByRWQQ24IZkNxIqNJRxYPsJhhqML8MwdDSMeuPTpfCJT1dlajTF+
qS5Mgy1z05BbkijedM+hWbU3UbCSBKP8NK05nSvjI0ZlJI6UGpbuRXnm6HrSSvI0h7OGKsatmuId
IRXOnPE+aNO6auduD7ObxQ3a1oB4w3UT9LYMJBPp5PXPML7/nFsauqJbycJ0gOyOsz5azDaKDDVT
1farT/+b9afhlow90d5PmyEkWwtdBbVZ61ctvz3NRLtDikq/RVgJH2kpUl6gosVDFBLIYH1UHiNO
MDVgrHEyMnfBpRUdJ7o6oJN9ZBJirv4Cgkusu2gUiGwkg9bjDX82vfQeCfuDLkBNCumCd6Erv6fB
gkxUxbDnznuXAWxyHC18qwwfgBXPYRtb7Lu6TCUj7lCVwebV2VIslkJdO3LFE4Zoe3mhsKfKmlhl
9um0SWgM0bgd4qozdTO/a9GC2x1W1IJ2RI6+n11jYjQ3ukI0uK+kUjL6JXIp6QGSZbHRwQSRu7On
FiPi5De3/Ovud0DbzFvzdwkv9wn0b7x4pRCm1wuoOq7Un52It4cdieUetQu2r7xtMvg9ldNHyG4E
MjPxJfFnT3nkBnIEdQmLHkFcWJKSeIw6j9ibJ6Lvf+MOUPrnyv9kFv3qhVvrhqjADQvUA5N4ZPZn
/nqsZM4Z/WMwj89bAd9hG5bRw54kb0mqAbMNSgZhELE93jfWDmtDg7XTZNRHlmZpguwIWdJ1mQko
+tCguUwxTBTR6nN378CRnpzHrkAZUf2IYy7wWvUS3mC2LgZrFUxyJ508oVS4+kzQEpyJvnsUDvBh
GZjnVHkaPwPXbH7QUnB2yOY9/pagaHgOvZDIq+6W/w4etvuM6mVVh8UXv5HxQPzTd2kMLXGhH0mc
vgfvoSGYJ6pYp0Hw4zeXCYvfY+OGWxnZV7H96Hu9nnBUsuPIVewLitRaiFXqvCp9FHmqdBf1wrLK
T9Fug6oqwAaxPp9bUSqnO3cNzvO9hMg6Epz2kuKfkCgpVUkFwN1B8poEfetf0viEjImb9R6d3aGb
VCmNxo9rrAj8PzF7sU5n/PlAXsDuFR2T3Jj649nGIEMPY4ZPecMRKIgeQebFKz3PF9MV7Gvi3ZGI
rcA9hB8Mb0R6cBjO7K8LWWdq5iSl7VEZp+cyaqPHN51rOSf2q0EivgtK9dsv8RYUOTrFFergGiYX
44BELrC5k9+peDUBG2p0YYyG3cWPzPI4Rk36lsL31241S4ABvOeQ03zdyYWMvzX+1VLCRBTP3Cvq
YcP8IW1vXrabppNagpIsiC+6RuO7iQalxNS08gvXqsIDpUXowNf648X1D8aL55BHgYne4AJnBkP4
t8kK6NwmHz/MQ4NDyCE78vuTCjGX/konvDdk1sN+9ZqU+mMdfEJM0SyOSMOfDDrugmId6r45BvpO
3XDEtAJGUpWaVfIwpmW7iBWvTfzbxlp6gGnv/4PQdGTXv7vgC1vArELOoAitxfd70QrQofT1fe3J
XXThk1flFq484vT8Db4xQCIdkKf9NtQIAZwZP0Vyao8xdQcFT23juqYmKKyGVMTH4jwtmWPTSY8Q
RaqKirVxtDvmPkU8ZaO+rGpcxluhoO3isA8Gp7lORMjELiElI8ZosLDeM7jXzbucODr6kxfdFfMK
EvXRLO0pk9cA/lKT6MZQ9IQVel9bM029x8HrOFQSBz6nowPGiZrzege/mHasPHJGFqa2OBWuR5NA
IAde39gZ+oGmY+xWylgxR7qqIgvpzT7uXlUavPA0MAfqdd9CvQJbBemFDwzCPwNJIkxhp62Q7Dwg
XV6qAtSeRNW05BbXnnM/q3ojJMsodW7fCTtajyTpvh0SuN1Rdq8ZI0xPMrrvCBB4wFXljglLvp1d
hpX7aYN6BPlLl4roWnP+91uDUhNhnU60ISEuPNpNeL4ehHGqL2jZrde92jDHkBOEC3ftDlOvh5+6
/8T66MeKkOHrQXeUkwW7xVaO3khP3nhKiDE+BeXGPIi1XpIRoLqBWWZRwcgAlrWpnkCtYXxPHLpm
5wW82LDrnl0B2H3v+s9jIFyfICtdRVVs20gVGo46LqehazfcXROEehdvvKYm+ar4PegUtEAQMXfm
YieoPksmKGs2GJAlJE9+JYeQ3C7dxBOcmq9CktELSaAhFQAehah0izd869bymXe5rUPQ+Z5OwXo2
qGyNItVQumc2IAOMcZV+0GwIfYWA+LvE6B4ae+2mD2qSOgAiydMiK/84r9G+AlExeayu6umeHFyk
L3zLhv8rgv2bTaSTM37PXbVEv2g5hguVsulXnKTkjSbX2yH8f1x3X5gRcRMR4zhAGq2+HmYl9nKf
Lwx1SYmVhp6sudJ3ih5yhSQCoBq93kinOVMUqPyd+XvpAfOAdabrRLmwlNTjyPCSbtkb0gkeg9yk
sEPAWiEhnVIiTLjjaq/2VBCQQmnnqivJ1unhWzcgJPb+uo0qgR7gsyCnAD4ZlPCmdUNCyeDdSJRa
u+mNk5ra02NLDJlmCsuS5YBWvzumuRTUBr9MZwAXuUZa57rBeYeaVyoS/8c/Z9+hH8RHqQvkLaMZ
NEEBQXNEPM12oGMVd2mlTlNH364bcU1eeyWY5zoHykZYo4H67rocWIgNgw+PEuLee4M9c5dJOhzU
UoIL71RQ9zNQUh/z9t64L3JF21UC1bvv/Fk4dF3vn4bmT7v20Fc6/ovRlotzQFmLL02k6CKnk99Z
5dyomqBx5WVIMRSOSweMmfy5rgvfOWnJ9riJush1o5ZxDoafhiD0t+7phGVnpqvReSkClVeXbgmr
5Se5726WnarkcTL9ngWep8kDOsdb/HF9/0EgsxYJgQY8Azx5ZX3/NvXlSdVRCFToVvCsXUemGM8m
2y7YizqiPzPE26JnQRJtP+Qehv253rVReNTkvLSp9Qog8hbqYaHSjBKfsN38WZh5zunBf6Zjzy1r
n3wt7wHuV9VevgnZhJF8sVcR6Js3S0sudiEqhDL1WmVY0DnhbkmLv9ndjfcsnsKxlBjAN1OkdgMq
m1Nf1p85C8w3LoGbxRILJ6jlXSr1SeXcxvhNOJBSUwKWYctOb8bnlDmgPbW3820Y7IJSrThxCK4t
uB5EsuMaDRjbZ/UPWVsBZEGduIUlG0NX5uf2ABZ/ZgUaqrVtlSVievoLflPbeMp5eaP4E2tA73DE
zq/8UkWlEb+qVdh5z17L3/oWWh53T9zOIl/mD2uIcciih61UC+OOy5uDM9WrXpVvFa6leP+sj2pm
/PRa6R9hGXPXo613iIWHjMy4rA2rC1IFxWdMG4grV4wbvWbmqGerbjXYvsbiVPdf49ShUU1gT05V
4AxNfZMGGjyGjZ0YFhmR2m1RbuM/HBAfeyaSFMk43RHlousZjX7NxfWYU0HLuUhVDDj3MaUH5ynq
UkBbWRFyCoO4tk4cQ8Kkb010r5C3W6pnQRj2Dq68MGLJRfVrJNZpmXx//a0QZIuwVx0WwegsKEbY
ejGVhBgcUv5CZQ1UJPVhRYVz0vWS/IlPioe+JaEwfPQfB+xAfBJQMoeLQmJSwWeduFbCDrF43dDv
euOGN8tROcZPRWCQm+xZ7wKCPLu2CY7zDUgBDIfEWzgz4lSK9CnV7YskHRRaTHQkrj2PIbxkbcph
CC7RxCUu+clUZAqlrS6xFaO7fzXS8ZLeUIQxjiat0CNEf7G2Df7JKIZdzkbMT9gOGAUzD59r7WV2
i5crOuVrwABCan6Oi/O/fV95uyJzgp+8GV+c7sUJrWG/nXsAK09IpCykHshmJjsyfkRdZBrrdBCH
6g1mnKthvMk9/nWPAfaWGhVJ7enAw0etxnDWzqeZSvLq8nWwUg+h+OtUYfQev0el29Q9Lkr4FsyM
9nD5J5l6cH6wKP7SisUX1BnvIWExRbiQgYe4yqs/jrmVLD3IvbX3CYWN35mKXYC9dS/P4m2Nu9Su
YX5hSokwcffngWxpFlb1AnqOMyaF9CmKfhD4csPiNV3Dul9R/3NT/1ygJ2j8ZkWATcnqfOm2aqjj
MnehuAOaPHPeAcGv+OAB8B7O0rwzJkrnYLRp+qfwCc89dLrp/sV90fyREjrfVhBxqEbWFbgW23VL
BvurLwF6gibBmKMVdUh/Ge+5KS1zL3Kk3lTAzQbltnHZmZmk9mm0EDYDqYxMqsWSAmK4x71xd8YM
bzeVF4CwFAqWUOCZLzWTFpVrnri5xDfmBa3qG/VXyzzXTIy0AQIdByFP1dF0DlLvRqu4a9Svdr63
MwZOZZPLCKVzqaafiy6BHk7BdVxAJHwlh3TqeEPJwpNCeYhIC+YoupL/mg/lvgX/lnlBIzqsYYee
MKncJkIzH+u8jYUtS71BvV1BLd4SuEaq12HqLRTHA3r5IpzKEIF4koqEnA4kFSopDUxL8JdeYzZF
hAyFK4YlGa4MmKBrIujmdz4ol2AlzKfBdmqEC6SHQR7/lN2aSvVTGCO5jG8xX9axKARRAOomhbhf
efMdsgH+2Fchr2i4uVhBOu9ybjIeMWGwImL+rmEzD21A2Y84UmlK7liTwQWcBvTRzr4ohcIXcKrX
UR2yzYWO6yLYkw76jwXzQf//bE7KvjESGxQC++P35oPnRKEpchT0uPwqL5uYOcaJ88CHmeM0aJtz
TbCYXomOhy5DFxgZ6T4YxaMqj6AxxDzDzb70cjpBft1nFwIawjFpUoP5ZCnmEjB+O2G3pf4Pny+R
hg+e5QjNrGs7S5rZUIDNiOnAEJa8nn+W9/jI5rzZFBieO0x0NM0hVOjr8x58D9MX9x/i0m/nAAT6
Aa0GnBZT39/pRnD+F0zD2HnGbJhW/RMl16v7yuC8BjlLHj8CD6xZD+kVa3vWgwuXy3qbtSljFbQN
5HgHbuJoHEJzZ2dp8hsNlDl5GK5Ovtc9sIS2Mc7QX5UlKeW8frhMz0Q/kLswoWveOfvt2Jg2emgW
tf/8p6PulcMsNZLrzib+ZvYMW7M/z04BQCQguB9Dr6zFhG+Hk3b+74XXZiHtd9+twSG0FAk4gt1c
psCHuromlfNeCqH2aBM38Cd38H9vdk6twlLRFV6RG5JiPXPwF/k2uckgmTZ2GlrhXJDOt0h35FKC
c16lwxSPv0LmcBPici0wNiypg2HguWnB/ALs7jUGGNyOQ07rHykZDj7Y5jnqFX3jrei8+MHB1y6L
sF68bq0HEH7pVsvhNdnFTjmt5JBFxrJz9OS10KfrJvQO5mV10yn+Y7Id5BWnUkuoIdiFoas9pryr
EZjQi9MvCY8WvifEN6slWHznmGHSKNg4wJ+f6PXCSjq8W7soa8AmWUhg+UiZTCtEV/fq9J4IuMlR
eWB+Ts9nhotCrLi0hKY4OCbe/uTuE1UV3rrknuRQpGCuiPxXdguYg4hfr+oO2/kYPdAfG0sc5ugK
6XyzsKjMKiKyVJJygED3w3hPpBr9dcDZqXIoh55ys3fuku5IIXdiRj7OID+rp6OG/bKKiKyV2sid
v/cyiHSW74hoJKSpoiF74wnwlIBq4XMlS/aBFnQAJnJ2xB6EhhSPU/BK/7ofPHtYxg+yziJMefXm
kwbxsO+8BYo13aaazq3wJQy/KvH/loCSnaOQ3XmDVwlWWakX9dPisNAfPdco4zSYuPP0psx5ebnH
3D4vMYBxqklLmmx7Nd/aqPakAj6232ctc2lxE9joHmzficGF2TEs0y+y+yTXp61Wvz+NEG+8cUJj
qhDlQBSzhv9sxlg5vkXMmsrPSnkshoDbvJ3qZgwr4rXjBlU2S9+prtc59/FaXx1gvZx9KRADttoT
heGe3pwTHGoz0ugAdaw92lN0T31deTciaWVLLJ1F46EgyzlpCVkQBh+0LbfImloCZDTU1NLy7Smv
W2OMyo2fn0q9JxlB5TybiMTQbfGdBJB2G8Ag7nc39qf+RfxuPcUjDc5dxG+yyVfV1EfOaNJg46qH
xBuYfI98rgoOxs1b7LIyV5Hz4mrbM1j28ymih65Tr8/zKpdQi5K07MC+9ROPpH+LzPjyMG2fexgS
Yc9KI0AnQXtkgmH+Cl6jnileLprcO51+UGtQSwgFrj7MY/xBvuWR9wvRg2vAJukwg2XctieaUpmY
85SYGT4IR+B3kZIB0f2PEsUjqQ/lhwNecCGu2aVV6nJkNIunusezwHgn0URHIXOaVKoxD6hW/k1r
XXEsx/XLVjv4R0KsLHjpmV+UAOdOWQTwendyOnrtlxniRwSj7RrbLjmtzyMm3I//ntKmPqbycOGp
geTRBQeQ23uu62SyDDN4eoRcxbwJd7oZ8xVnOlsPMXyNJDc5CBQwWY7TJ9Ww3Ih2QUzhaYSsKeEX
J/IR6dVHMyKShEycegveNnsaLyk3PZyzofIFmG31F/j1zbXMGOX0UTfY7dhhrdr9Hk9ybh9veTKk
gR8aDlIuU4vzclTb8s4bSQ9kbz0CnaAFSrnWcJ7Xg8bW0CS8DweB0LXb4/XXc8GhGPlaj4R8AIii
tL10hSqkpytTn5Iw7D1m2cS+mHAMOYMNqNRPZg2zWsFVsPa/3PEdzwHdWKLvON/AJoASxJvBiosi
Kicn/7H7KnR76RqpvS/pb5IhnIIk/KrapU1RU4ShRjrNqkbC77vBOzVgxyMFCE/aasN4JLNwmBek
tr+LJ7J5Q67gvktED7hEgyZbr/wQjABitjtHuc6zvHw8Mi1ajO1Z4WLYS7HnTO7KmctgOPOXIjJa
Rzwxk3+7wGIldt+70jpY1UzGTnbLMrH0CTFQbXIc/4uH6clufF8ivN+zKw5ljqU9OM0pvMqUAkfG
3Yai2G7Idb6EolnnJ4wz5eDYwUWB3Pn9bXxk5KFGZlgCXcqRAVZuabgJggQf3UfJEGon21nq7Xal
sEFifPRoI937TGqrx3LckTrRJA/e0QDC3lymjlLrcmNiFhhF4j7ZClBPHF49C0aRmdOAcYXqinNb
IHr1dhLjkUCNMeIKnufiIBeK0kHAYXpv8ahlSbzkgGy9BrA3qBuOaj8iTInfrH1zAakYRtPNaCUV
ByswGRAlrnkfq/a6SKjIBSiGPr3sO4Uh9qVXvfNnmHa1prNUEbbFcNua5gc8FjkGrOHm7Al7rSAf
y408Yce9hK3569DJU8KuWZ6m4/wiD57TOBBn2F0YpXFJuKtd2kXHVVzXuEmwWyPpactbL13Gwlmo
s5d3Y9rKU7HF3bnluphQpnQeFMWibBJbDUNVSVIm4QuCFpIau2Abx9HmMxJCrDQ9InGNHTOGMLnb
Q3tE/4i/bjbt6VfjBQX8P5TVx8Vy3uHYB4o3/zjE299saRgKBTk1bN8BiM2VNeQJHF6NiG6yX0QV
htpahcXAifuvRe1s8qUFyq0OZogIaLAxhnPEjyO/OTDEuJwqO+vUstKlef/9i++fHbWNWmDliM4Y
QsqMH+JSji7lywwwWQaxvG0PxkISB/nLc5nfS/Y3jTml7+qt5sNKm+kJUycqQPr8bg0soZCq3wU8
GdPQNSQs/snOC+jkBt7iSKp0aJaYlStkrsa6E9wDBHtc9qdI7cQ6LNU4mqPt7LjKU7/O7/6R6jD7
r32AoSFXt6oyThF8MkiQ9hMSJ3BlHAo0lyYqZ14hRIZIv09IhBJA5wBXbSUCY5qbmJtwdgbdmBgO
s6o8y7Gg8GhQhyVLfhepfbxC4gUIwP4IjgIxEOaiMm1iO1n0/n9UdsNadUiBw/OVQSP8F0KnG12m
jwBzi9C/2ziLD0J8HLXmXs9uP278VW3jz/+XgUEtcI/R5bT6piPQ2+6aFvfEu+0FWZ75tiMt+syG
vaHb5fsis3XkQJyD
`protect end_protected
