XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���@���C�8
����w�`w��w��hv�7�2,ȹ��+����ׂǟD��'���T�µ�v�B �
��*�6r���=���\���R�K��L[�bb{z�q���l1�B���[^C|rq��DJϬ`�퉚"\�+������b�&C��X�©%%[�de9����wu��DZ����|r���*#7#��~�5�txx*wּ�[�_ܢ]�b�a�c#�4�$��!J��V�����ь[�:�h⋛��G��5k�V�{�X)��)�~$��&�`e�;��_Ա����8�K|T�\Hpv�8�[z�׆�y`Ӡh�po<���KY�r5��a�(�߮�=a���,��ÀK���?�½^���j��b�l�U$�1��)O���k�7���i>.��`���}���s��1�?ES��(_�IK��3�9)j�>��R0��t��(T�7V|��o�`��1�_�1�'�+�����`;��	�%������;*e�5^�����>*�5��b��C�\����˸u�n%�!�Z�w��5s�M6�?)*�F1�D�l%_H����X��<�c%K9�Z��q'vGa��޼�xO/��5N	��m;�Vm�|�s`�O:u��s����c׮�w��ћ :��S�vޕ;þ[�9N������b���/�:M��wAQh#T���X]7��𼄠5sI��0^p��Ȩ����4� SSY�� l<�8G���"�����^&up(���{�XtXlxVHYEB     400     190��Զr����K��o�,��5�8V2��n��iQbh$V�g��D��(�4��f�k���	9���8�4��t9������)u3�$h��xz\ۜ\��c���,�AѠL�5T�B��;@��5dySG�+Ҫ_��8�5�U����Dq�8M�\,�9��V��82\Zhŗ�_�Sc��tܬ����vM���h]�~C�F���*t��q2�_/���"as������.���B��]z��@����ͱ�'�,:�mł�틭�^#s��v���h�������X��	ԥ
K�S:\�d��I�@�>�= ]�8���I3(iq�([���^8�� �~��'i JPDg���� mN��N�v�H�J����`ՠ�W�:�4��l�@t��!�XlxVHYEB      3f      50f2T��&�!�"�hc�4�JH��;Y���p�D>���h���� "Г?va@���Y9s�ly��>J����&Os��U� ��PeN