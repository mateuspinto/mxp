��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���� vU����U�a
��0�j%�+1�X�aJ�t���W
��S̃N!6�lm��F@���u��DA�TuF$;��7s��U��sX��%�09�/� ��͓����w�$k6٪eSY�~�+f���6�p:n]���Y�s��QVY3r�e.uW���lAM�����40��]:��7'�~uؗ��ұҷI���fK]L3�9���k�,DP�<�P�b�{*�5��/��P�?�I�vX��b�|���M�{YJ]q V6H���ptXq��@�g��lu���+�>�s�bQ��-���y��a��w�p��/�r��'D��^X��0r10>=^�o������gQU�̶Q�n�H�
~&��Л�P�]���:����%y��#��G]Fw3w*���_L�1mN���`SA���$�/�?�`�#��@��ր6wW{�V/:���E`��!�����p9�2j���]]�Z{f���.^8��j0Apߙ�B��ǐ4��ׯ��?)�t�l��PL�.foŗ��=�e]~ׯt�����ɈL�;�0/�~�XM���>�%��"_����&�����Ej�{����1p$�q�$��o0�Ss"�ya6���߮6.r1��y.¿>�a�u�� :=��%���C}@ʻ�q�_|�M��hLp�o�(�#���姟��2�,7���H��mCѝ���}�����'�"��{7&�Q���7R+JK����sF�
j!ԗ���%^"��W:
�T�&����8 �Qʷ���#*�M�ˊK:|mƺ�壽n���*������'£05�]�FvM|wt*�%g��B�t�ͣ2ha}�9��!��b����h �x� ճPa��d�|b1-oy���E��h|(�j�Cjz�̅�:��IH��%)��ȗ2lS��G�<V�Q7ӎ��(��C��4�f��@�v�P��ȌU|6ØYTA�@q��(��j�ѩb���.(���%���6ĿN�F��ڈ�^�
��ۇQ������M��Fmb6�}wB��Hr���1^h��45p�A�d�|�,@�� �	�{يIl�=h�bN0nw�B��(��a�.P)��������-�y��M7j�}����e!��O��+��j�z�7�(�}#ZSPR�GQ4y���x�GA�Z*�Cz��ȉUA\*y��oA}[}t��Jf���mS���;�(�rw`���ncy���7�|�7L1��,ےBI.&v~4��!��'M�y���0��|�J^�A��r�3XL��	 ���h�6y�4i4C�1�A+�Sn�v��YzURdOd�n[��P�`��������Uu���h�}}d���C���D����widB����4,&�EmB�!_��g����f]e��صmK��<�>p��Z
�l=�O�Y�"V��%�ER���5ܵ���rc=A�0��q�OvJ�c�]�Z���ǣ' n���`U���� Kr��c-
w��� �1T��d��m�nn����Oq/�ۡC/�Dg���/�L�4��T𐢢��ꔛ���< �(�KS>T5v��i�kPg��`2k���E{q�u�����L@#���_MQPR%�{R:o�gA�IY�VQJ!ϼI��󨃾˱�2�'ͻ��-���n䭗D�-6�קH�Բ1_��zT��4���`�k��b�z��4�(6{�2Z����v����dDÊ�*ɮ�ǃ�Q�8��2�-�kD^�*�;����.<{߯b��ϣ���[�9�;<eu0�3��ғ}"V�2��x%�[,9U�ɭ ������O)�jF�4nUs	���U�?�����r�/R`���L`��[�-�c� 4�8-@�KQ%�|��m��ۆ��b���g��/��Kk�N�0Y"G�,Ch+?�������Q?ޖ~�y��_����n�Ϛи����I�0,c�7{�,K���,�ŋb�aw^B��o�0�'������]��O�蘒l躴&k���)�R�)�,VCU�D[ܳ ���z��	�������^&����\���`����/^�{}k���I
�����N�dc���v�c±q3���z��U�/Zޱ��+Fh��$tz*{e`p�7mrN��[m����k�褎�u*�a�,埰��u��@���\Jy@W]����^�#��v�okU�%��v��&�Q��5ʌO�TqN@�a�9��|�c��T�tO@>�ħ�O36�0��z��9 �*۱�
����\��SN����8�g��xI�6ͩ��P?�"�0N�H:|���q�M~�W/�2��L��O=wkG�
�P�Q�*�.���<=b����s#%�:3l��9EmmAZ_��D,uP�M��&��	̓��T6��GxƮ %��,�HW��h���XReꬼ�&�r���#]5����D'���T��W� �y�9�6v���_�EX�؎p*��v2���i�G��&����4,����̤K���4�aU� �"��(@� ��s"LkH�M��_�*��v�ƀ���K�%b�c���6f�
��}d|?䠗D����n� �h)JzV��?��{���Ϸʢ���En05��ݜ�K�#.U����Fp ?w�* ��ETYH�^��»N#E��~6�m��;�[�J�o=l��H��K�W�E��V^%��M$JF���B���q$�<�Ġ����(j]�&�anG�,G"�Yu&r���@�K|�'�x�Y����j����R��tS��2(��P�\vR ��_x>/�Z�(�%�)��p��L4-���/5�{�P5�ߵN��fR�K5<��{Զ��p����Q���"�y�������ݼ�o+Ӣ��vқ�D����r��;u�� S���:��Q�j]0�ɸ����E�X�7�[�|i�����ek�`��ʓ�m��C�s�"4��´��C��}�7q_J��P�{h�(��!j>�-1� ��W��ޮ>�#qfen��dc�\���2�ͨq�W�^V-ă��!���?�j�Oc=�_�S�[�E���B0�Mϫ+=��!̋Mmc���`er�t��d�:￺@^t��	W���Q��I��W��Jmj��n�a*;��R��Hv���]紝��s%)�\�up��r�rľ��9��1�T�(E��C��@�4�v�2	���N@㘅o��o��Ң��!�D�
3�|Mz��l�@�ǲ���S�����p&S���##��7��5鍚|��R��s9�0�fw��-:�x2����>.�VT�h��]80���pva)g���ء��r��qܒ�o6�����7�.P*O?q/���]�m��)v�2�z���b�JlF������oO�_��t�R#���m�	�]����ߚ+�����V�d��
���Lf"��!�R)�IT	?��?ժ���dy��j�3�ӭ���2��QF�fXJ4>Ņ��F������>� Ef��1���N��b�7�#Z�8�`�@ x���H��;.��;.���k/����~#d�Q�&D��2x�&l"q{U�.X�*�~��.��JL�I;mM�ƸD�kB��6`��UB"K���1��ĒH���`E���:�A � Hm="KevC�;"�����E��M궃MC�$9������Ab����>7���\[�\6�������/�2p�g6v6��P��)���!
Ҧ���<�p><&\TO��bLV�v�n�����"�u%L��H{�w�4/�z�9��~���Dpw�D�0z�$S��I���fz���R�u��m/�%.�Svı�z0iv
�:����/���?���n�Ɖ��.u�ru�C/������ܲC=�^���|����y�~���㖇0���+�ݱN��a��/	8�0��:���j��]�9�֔���P�m�DOK�<�Ч�6:+N:��F�
���E�7D](W���&*u��[X�ul"���;�b�o��\�y^��.`�A�B�P����X1O��%~�3l�3�'ҜܚF��"���c�(����������i�P�kf�"�x�����I��f"���\" �2gf4��G�N��
-���+�Ct�Y3&�6��IvB��|ß�?�!/�C\`�{XQ�'��K���� 
��5�nݸ�+��6h��d0��q+���/:Q�>��A� S�FJ��=U����3�v�"w�m�&:j�WÀ�; ���9��T��}#jOLf2_���׭=;D��PęL�<�����F�Ӱ�ZΏ�$����h����̃�t&�43:��&`�������Zc��S�<�3����(�����
�1�:�(�]\Y�����,	�f�v��,.�ff{@?%�%r.�!�p��ǫ�Qe�&��N��o7d'	p�m�"���XY3!yU9�&��>:2;ը��M�F`[�5嫖w,7 ̆�&������1��D�F�)�P��zb�)��K!�p+�%n�HI��t<ƥ��Y���1��L~w؀_~��3-�n�;��<���|���JÊ�1Fd߮�k���ZK������Ì��!���ˑ����R��3�"|{G���/����.���󃬒��|�묇Gc�i�GwaFU�?�y�S��Am��v6NA����p®�῿�.L. ~��!^���ͨWx5}i5��~SvZ�-j�?��mg�yi�D6����G��.���8[G�� ��)��~����ZEɽ#�-\�&W�m�g����A]�UH��ȕ5����6X
eį'�P��I�8Z�#��{�����������D
�-���)!ā��.$�W��Ɩ�0?��"�5��5�oצ���N��V��x��� ���1�-t�u|��3@�J[jU��7"���pu�1Erԑ
E-G�3Ddʨ�AH�ƚS�u=W���F~W2e�X�&�G7���Ԓ��KA�."#�nʚ���u�=(��L�w��0�[ڗ���`�;v�v�� >j��-���Ѕ�� �E��p6�Qt����<��"�3��e���~*�+�	\�����F�H��PUtԌ1$��ʑ��P��G��Z���ȗ�Oa� B=AfC�t�i�ހ�O���I�����t~�6l�hd�U����.S��NVVV�j�a���:��k�Jwy̍�P�I@lC�J����8�'��	'�����pfwl>��OW��I��F����e�l�҇7 ���n���@����c��?c��G:'[jbٶ7�q#���T��U�Ԯg.����(Cq��NÙk�i�����xŅ?�z���\7#��_̖Z����j�YP�F�gr�}�n(���7c�5C|߅��Nt����V�m�f�~A(&ԭR�Ʈ-�.�E��� ���h�ej�5��'�}X��z�Ux�N�����ܼ8�-��BM�K7����l�VH��L.�F�+ɓ-Y�P���Y(2c²��Ҏ�&���}	�U���R{K��Z�[��b؊��H"�ec��
fkӆ	)��q�[z��Wn�����ơ��`�W'�4����

��ژ�����~�h��V7�0 �ùE�
������ܥj�.z�L�'�zAnaɝ�.�`�#5�Rцm��\!B�0�s(s������6���]w���'2�f�>B��E���.6�.�6Sz˾t��-����Ĝ��Uؼh�N$�?M�m��.k'8����-AxӜ�Bq��dTZ{'���~V�U <�-D��Ø��|�p�F2M�*!Ri�u<Q�̜C����H���Æ��Ø��X��ò0{���~��w����/�g��P?hPx�B��� �O���ؚ �t��n���8��f��1�>g׺֬��k�C ��|$W�Ư�u�O󃫁#�ʇr�[C�?P�g���=��e��� �����4���f�Y>k}�� o��FW��{o�5j
yW��bs���%ߠ Z���;?�3C�<�i?zS6�m�E���EJ�)�����m����Q��t �fB�=}c�{�EV�"���z}_�����֨�zeB %�M�p�ܳ7"���v!+,�+���y�4�U��7����@x{ե�j$�"S d%R,�	J��LwO	��(֣.���dF$/&�g�s�I��c��Z^\����n��%����m�i2�8uE��%k)���x6
Gq���r�w�%9�b��ј��q�*M"h�L]��9����r=�j���l�c����8�aR�y>�)�r�	�� ��ߍ,y��1�e�<A�t�q�{����Q[Э�i��[��px��UU�����-5޳�a�*��Y���Y1.�({�p�����j%�g�/+V�G����5@&I ?��BWP�, ��t��6]��Q������2p'h�P�1gJ/�.o���I��������Q\�^o�CA�D٢@wD*e����C�&m��hmJ�
8"8ý2�x��U�E��8��o�]s�K�P<iB�0�t�w�2���;�|w��Q%���i:�b�iR�8�>c�����Vۺ^��T8�.�c���������어�Nx�R�-�侖��+ZrL1"�7\�T�)��azD>�\� �w&�S�c=\ܱ�FB⧫��\Ҽ:-�{W�Ѡ��Ib������,%Í�,_�WZD�:�1�us�����th�M�%�)z��8�v���S7�	�v�Wsq�݇J�Dg��eW�^�����<z���X	�ao��_Yo�Q﬒%'$�����Ӛ�7<���C\��h�H���:���`|����U"���b��}�ǯ��/�HFl6˾��*N�f2�ݼ��.��)D���;%�!zq�<b��(��<��9�<�d� �g�~��34Ү3Pj*��B��m�%LK�T�����R��O��:������Õ�͕��g��E���	������;r��Z��j/��7Ɵ�����%v��B�E_�l}=��"$����7�q��i&��r���VN@�Z�ǚ�J���:c�r�*�� ��2>�s:�mOu���.��z\�(�ӂw �%������̪l���,dBɦ��4���s\��S�U���e.�w}D�3��J9*T�0;�ߏN������#	�X��ʒ�Ć_.@;�w��?^bp��vɒs�`�|���$7���t.�"��N��#�4���A^T�Qm��d8Z��[k{��\b8㒌���M�G�H��Ӯ�&ʌ4��Y�U��T>X�H%���������^�	��{J���Y�ey�fG���B\�R�=�{&Y��b�N$#R4��*�"Hٟ�'�����N�E�7�wX1��C���wjx���V@&��'(�����C�r$���5��F��8��p��:�O��&�	��"���(։~�o�4�;��A��$�ȩ@(��u3Ib y�,8h�����LC2�	Ի,ɷR��.�s��g0<��	G��C����Jb��V@�jb�|�6��
�t��^�����s�i���R�t��'6�bJ��CY�|���0</�&�|,J�Z�H�D���N�X޶x�g���)����.����y8�9�
G��c���:��A��AN��s�2OZ��N�b,�� ��/�_w�����8����k��R�2(˿L�\V�D�?��F�d7to��Ib$�y�I�zz�rL��w�B��oKz��~�	��x�	�����t}@���PH���-/H���t��SW��+w�v�Z�%Ώ�h ���-��՝��1�%�
N��8���Ds8f͠!�+��p߉V�����x.N�߶ #�y�>��g6{&��3Y��Oܽzf�Šn;�Ld北M8�L�p��?�!�7-�-�c�C��UK��W�0I�&���G�:�^d���
w��ru�郒��?R8�e����\e�JD�jT����7�.�a��ӿR�'A��3
ѻ(G��\U��s�����3"v�l��k�T�p�l������(8H�.��F������[z\���ss�?��>��xG'����.YN�ZdB�ޔ]^&�WO1�[����m?xH��Ƚ��ɋ6Yv�t� U�s�!zE�򛁙�'u �ֆeW��&�Y���{CF��"�_�u/r�X��c}�7����+�R�c��+Z���ͿM���<�A���u$u���J��d���ω��R��ڀ���w#��8'm�H�f�Q�A�oX$\,5��LǼ*fH�Y�KU5��	�O��V�~�T}�qC]���V%w��}�Ê�K(1���_j���L�CL��l���������I=�WĒ��hJD��,�;�_�B�C��!�H�T]�`����S�/ۣ��/[@U�oK�s��+N@2�bw�5R�Cq��&�QZāH�q��EȦt�C��{�o�Z�SB�̗.q
j��Zd��WP��e��(�(�\8 �3}܆<Es�����2�s|r���VUW>�HWr�L2
��K��/�"�* ��^l��8ݦvX��[Oz+����.������D�C@BS-�f!`�Y�n��{iy4�uT!S�����
'�����v]$���Wac�)��2D+2��)�aD
��C���[C�R��ȳ�,�hztн�u��U�x������w��#;��?���h,I`'�NT#����ߛq#�U�w�Y��8��\�eq�
�a貘@s�Г���l��,�ǐC:S#���8D\?��x�'��c���܎[_�;�ⵟZ�#7�L��7������%$b��+5"'B2��:A�Ua�S� ��!=	\۾嗍�'�D��vݸ�V���hÁ�*�'AW^B8`N ĖAɯ���pį����,^���%��1KP��p��s;���i�_S<^��4�map���Î�M��/��;A��ӊ	��Z+FU��g�ᗀ"�z4�T��}�\���4�0�a�g�d�t0�-7�4a��q���M�ɫY�=�YU�����'F�����b��B�e�����|�|�-�RbbҌ��h�#�>�O���a�?�^*����b͡�c������	�Fd�է�4�

�S�>fV���n�A��F�.bCc��1�͓��69�9֫��A��M�I���EӋ���FC��i������S�P����`+cVe9|���ﳔ����l��{��;,�D��4;<�6.����Iu�2�s4�K� N<��.	%�ɚB� ߸��y�E�����>�E�*4F�PB� ��4w!;��z�f(Wq)_|���Z��	��J�AP|`]�/���Q�����|�|���Q���M�8乄���0�l��YO4x��Us7��Ho�3��"��o��U��Jݑ}04��ny�;��[_m�ֶ�Ӊ�##
������&�Nd���\?�����X�݇V��J�wA�%�hVM^�2��w�~� w�J�_b�\�⾿5^���l��?w��&�NG�����{��E����ma�����4�\,����h2��T4p9i
S�m��N`�1���b��(=�C4,���� �)���助R�>�_R��>���Q3沙4���Y.�{0"#S��B��\z����o��?�y�J�N�f��})O�Q14�{�)}QݗJ5�s�3��#��ֺ�p�D7�HKG��Kf��Wh�P<E(&wx�~sl�i�=
����� ��jϏ� h�p� *����e�5��X���޹��%�K�
�%�����[�v�ie�08x���N��%�H���BΡ�� l�P�M�@�7F4ݟ'�QFe�
[(��5h/# �v�}��Y���#����~��1aa' V0Hv�cF��Mڂf;֋xB���f���\�5��\��m�6�?�m{j�A�m�7��&�j���>����<ϡ���Q��.xz�(^��O�b��<A��p����f�Om=��� ���٥ra����e��ag��?bd�n}�L�ԓ�s>1�Yw��I= ����O-��	_�C�$�v��
.���V�[��*��ŋ;>�]l�-�_��@(R�9˩X/�,�S�ޛ��B��s�j��N����V�Y(�J���'�����4DA����-*})�>�(����w덝���Иq�:����%&)t��w��N�����/I M�4���ػ���ԥ��p���@�f�zU��ſ_O09��s͒�M$�5tlOWu�^�ov�b�u�5�ux8;W6����(1-l4�u`���J�������j��tb*vT�f�|K{�d'C�����������px�@�>�>!����eA�@��ii�?(6�.s������.y���'Z�a���Cj9�3�E�%�~�����:myL�Щ�zk�� �7�숶�P~q5[�9� ����<�_0v`B��nE�pM�Z��a֪��ռ+��{�m�W9����2��������Ѻ�E���Zx|���%�٦.6�(
�Џ�
:����*1&�l��D7�YzD�z�Сwo�s���잞�g9B�&8"?:I'
gF$�A��(حMi�\ka=�ɬ-g����QK�:��I Y�yj`�
hx�?�ez�k��%;aj��G�q�XG�<�/T�F.�-�v�ch��{�Tǒ&g
n����l�E����/Y�-t�e�ӴD%B��3�b4ϺwHCl��	X�![���]�A�尵Z��o?s���E�}̻:7��-���{_a�,�l�q�o�Jy�7�=w:�/HQ����p��F�V�ۤ�y�C9� 6%�Z���j�gL.��LJ�Ԋ��"�)Ҧ&�ף�+�I�D� �R�>�%r?�lh}L0���Ňi#L3��Ln	`��#��:�R��k�v��{�1��%n:d	������.���ؙ)І둝�����ѩ�!���C>3u��,fOC�H���V�s��q�-�s��<�n-_�? �� �4���m�"*@qy�e�v@=�Vq�mK\�P�7؟ZK���Ơ�m��k��2�=@G8(�Q�𣉩�w)[EE��c���o-ZLHC�x���=��7�Ph���w���)x��2�ATOyX/�/���X�'�N���v�TO���I��1M}ĶZd�ʟ��1�iB�)T�<���|l�
2
�ة���<F✚uߪ�Fb�l��Db����.:/�g_�����xsr����z��M'qwQb79�ه��,Je�!TQ�$�n(\�]$E�,��tg@��IV�Fc��JO� r�L
:Y�LRsk��n��S��N�U5ހ���.9�q����?��EA��M|���He�(E^f��^��t�v�}�J�/ǅ�E4�b���+l����;p�y��S1���o��RS�Z�l[�K�&����u�6}��iS��(
��>C ��z@�w�1��p=9�7��7V�ޥ��8���P�PI�X���>��ᝦƵb)��,�o�	�ܦO��
���S`��a�S��.5�&���|̦*�:{��a�30n3�R]̼w$9_{2�#����q���C�B� �����N��� �f['DI�C93��G��T�#;��~��I�����{M�k��kL�
��ye�tS{�����M��q�����;����2��z��ͬ��3����[Z4��w��:η����`iK����M���^���!_�����r�u.���ި	�ᵿ�f�ۘ�Tv/�I���AÍ�񡢭Z/�f����\�� e�����ڥ��K;O����rr�cw��wA� MĠ{�&,>�DD�n�-E�<bx�/����"�J���bD�����MKon%>bV�	��v�4P�pR2\�n����ވ
ei�t����B���Θ���l`����|ȦԎ/�� �fToI>�E��O� �c�|سuTFs�ؙ]��+��;�:T���|�-k\���.Ŕ�cʾ�25V�� e�,�Oo��RV�Z]ۃ��M=�x�ϽI�!�K =7Đ�t8"?:8E�����U�P��y$埲��+Dl�O�b����)��e9~�6�s6��=�3f.��%�X��ZwR���e��;��w���!&�	���kF�%�}+~�jGF�z�	u\�M����Qb}�-���8:I�@�d�I:��Ns�RFe5#0����k���?!�N�xy���~5�秼5kG��]�����i�9�L�����A}v�Є�;m,K݁���*�Ɵ0s%����X���Xx[c�ʒ�%�H�R��-ě��}@��k�Β8V;�I����g��
�G���X�0:}�������l�:��n�e�"��U��w�r�s�N ��0l�+��5ƛ�����.��g��z��?�Ai8O�-7�Ҕ�|�L?R��5�C���y&���SW�"b�� ��٭���lo�0܂w�O�,{
H�j�꓆ec����a��R[��CyE�`Ҵ�&���?H8o�b\��f�� ��u���]��\�ѳ)���#���%��������)(�UM`
��רQ��X&�hRI��h?NG��$�0�U�=Y�����{�����Q�x�燮-��?jV�7�
��*b�E������ݫ���� ��{�����(&����4��#S����(ZX�?N����<P-�>X1ͮe(Ѕ�<^�:�������
郢�64��*	���D:�n��1$���#@@�2A�E�*����Po��R\M�L�<}'�Ӓ|�c0���gQG�	�_ǔ(%%����]b��h.�lP���߂�D.@Q�7�<��
�b�}7-�ɴt���6L�p�?i:
(ʹ(�x��@"��`�+���z:������l��L�<d�*��t��Exr�#�ڡL�s4�r`��!pk�C������@1�,��n�-/j�1�|��(J(��6X���R0ٓ��+��1l�~��}0�`@�ӄZS8r0�斄5x�Y��1,2�N;�`$�OQv�F��$8
(�n)Q�� �DQu�Z��Q5`�ȊU�d��G��Z�eϨ��C%ˤ�or!Ro�zX��;埯 ���]�	 �<"X�
��'�߹h��v�����oμ���lI�'��/������u�WC^>���
tE�S�l�c6��������L��q�5Xר0�	<�~W�Z�"V.�d� �_�4·���L�S([B?�[YJ�D�SP����Ǝ��L�1��/�ѫw�1rAgG�{����0ռ9S��Њ��R
�Q�*�8����/ 
�D](9�?���ͺ)0Yz��_Y��u�1yS.����b� ���%�!�����Z��CA}d�KVK?�ф�&��8Z�<x6��Ú�G����?��-��+�����X�J��K�=Y�B/�?A��݁!���`�LU�-2���Ƽu��5�ɵ��ņ5����<B�Y�:;�
���]�f4!@��1nLG2gH��WOK
+�>�VB�T*|�B!NAς�ގ���H�u�k��c��G5� |*�i1�5��~�(MGn��@�vu/��e׻�B���{��}j��!�?%�	D������6 @I�a,F9���"����õ���d�p݇ ���˘�v^� ��it��BڥR��6~�e%�8X�}Ǌ�`�f�Y����h����h�og?D�Ϫ�.�(�����_���5�M��_�~ͷ�B�8�nr�r��tF�2�ݖ��'���^��'<&Ž�{��zc��]�����A9�P�a��ې�q���u��	f[f���9��q���Z;�epQ-�°E�':�u�׏w��9�D(�l���em����V=ї�	�O���O���`4���L^��^�ť+�r����a��L����6����?������MC&3kܶ7Q0TgE�D��s��k�,jedFgC��`x 9Zݭ��5��}H�,12��
]�E��A���@
����;����V�̇����/S����w�kXb�4��F�4a�.��Ɓ���D^(�Y�����2�2U��~j�ţy។�<1A	K�U;�/2��׀�p�>n mT�_-��2[�[�>�ZH:x��Hp֬���u�-K��(;��d��++�e�l�~S+�]b-�t���>GƓ��RO_ГE�{�M��7�;���C��m��2/Q" $l�VR'��Z�d䴀��?�k�%8=G\���!��\�c..~����$�����^�y��`�Y����w��>��_p�lҗ�)�.�,����R$���T��f1�<��"]u��qc	e�H�q��׾Αt�ଁs~���G��9K<a�]	����	�3ͻ9>`�/u\����n�j�����_
��h��qa��k�/��D �?�6.7zp��Ǝ�9��YYI���׏& ����������͆ыR�ǲ���T�$o�Eߎ�q0qOȒ?`	&IR��K��