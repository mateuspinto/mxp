XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��a.F�[�k#z�����A�E^�N�h��w|@^?��;lS��	�A�~,و%���u2!��Zo��Će��&�)b�i��a"�O����1��-�[���$8>ʻ#�j��[�TW�x6��aL4D�-�A�}N�XA��7��\l�n�y��Bb��:b��z|�]��Q�\B�d	�Ѩ���Om}0D��������s���ȅ>���;�S���&�����w����ls%n��,�rЮz� TIk{A�f��!x`k��#��PR�5_F�1�aO�kI�Y�W)����gz��^JY�'׉)��<��eҾL(ܚs.Ӗ�� �Sk��F~�n�䶪�*���g��I�����������A��G�,m�z�ǻX�\�v��q�ֲ��ٽT���A�}���`{�"�#�2cs�)+4�%��6��bH�j�-��l?gl6SW���_[�߬��w7�dgA�12-4j^m�����fe�-�l�;Ji%�dvI����74y@�&��T����]�r�;e�mI����:��M2�I�H5���pYM�����]d�L�G�~��̬���A�q.���DC�|�+�-�K���ߵ�=�k�H���;����=B����~�p�ߪ�1[��Mֈ14]F�����X����&���
���״�ZO��絪*P�vz�0������G�a�h�.�;�}�9�5)� �
6)�fJ,�&���*Bnl��	$�dR�c8���Q�1�L�O`۠�4`��XlxVHYEB     400     1c0��j2Lڤ��P��L�5F��z̓�b ���pEM���yF�A�O�Yk���.����J�9ԏ�g8F��֘��G{:����c{ۛ��.������^~?	�@+G�<�q����[@G- ������KXu���ZP�4�ty�n���,C�TK��\�\3"W�+8��N�����z���~�^���kp����`���v�t�E��|�$�!E�s��ae�Ri^�UX���6q���,���R'�+q�@����Y��`�Z�1��}h�WP,<q4��,���9�vˌ˦ZrWG���/%�#�����Tb��F�gc7�7�n����M+AZ��2͇������N� ,��ALH�%��W~'���e��K������&�j$���jl�	( ��ˑ!��e�
����'�)��ޚ4������P����NmѽXlxVHYEB     212      d0�����Ֆl=Nۊ�L���{�v������"��;A�\a�fs"&��@OΧ�����=�hG���؜\L��1_��O+���W��~����n0,�L�ַ`��ra2��Z*��7�������h�?�,^�n�F�%�>�EAdҠ䖾��f[�7�)���(���3d1y;�<� �|����������">�ь7��OG