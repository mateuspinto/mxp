��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l����$�+g�M4� �����8���{�ck���:I��Á�y���)Z�uhr��;�����N�yJ��g���zIc�ʐT�r�`>c����4��Yz�0��S�S�pHvW	�,4@ �x����T $�p�o�a��,�S��ۡ.�-���:��Jz���a�L8�۫B1I�S�|@��σ
�J �!�9�M�*��;6qq:��3���$e�8�$��~�{�M�&�v����1p��f��*'Ŷ��CX=�1 �Y7�_��G�����ɈhKw=�S@��Vj���!�a�+�)�娊i�����eCt���s ooan�7x6�}��:��)H���M�"�l���z۲��d��+�m��Y���p4���~|�7�m�oL4���P�'csţ�����5̀/�ِ��A���ƍ����iw�r�.�ڈ;�L��↬�D"�l��Ȳ�A2��g�s�V��c{�����S�g~��N�a1P����$�Zy�`��1�ʮk���{#�f��!.xGb�����@!��t����"=�mZ�2��+6%2�� 5KnBf<�j������ϻ�[,d2!�$���[�"���U9�q�b��_���>�dۗ
56���)��|��Gv��Txm���`V�+`4���QǲN�}�+_��/k�s?\?�̋�,@soU�E:}s�Hǀ�'���\B�o��?1HVVe�ω��g�a4�,�@��@��U�ln<��s���:�|�#
��11�����U|��U�e�3�v8Y��Ҥ���4�@��aj&��v\�
{�	�|�p#�̆kee�Ɇ�΁d}pP�n������W�MF�`���U��[�Ax��}ذԖ}E^�])'pd\�1+��ijK�T�u�T����y> y:'̬�p;�XW Ny�AN� �5^�;	J r�k�Ww�L�'����R"�mj�LI�m�q|�&�$���J���ީ�<�#:�х����n��U�kM܄��zV�o>�C���U����$�/&R��Y���G�ض�z-���H4��$��v�t�8D)�ѽ%ѸI�s�.X�<@1Q�w7P�8��]�	=x*��=P���_/^3u� ��m�tI����Uo'o����w%��F�hUe��"t���kQ!xc�j�ʽD:R�s�n�F3۰o��&F�vd�o��W@�������w|�PÕ��;�-�Z;unRN��0RoB��:�c������g�?ų�O��֕u8�u��"a�a������k���|v�n�q��b��*�w龈&��9gj_6�lZ�F2k$�M�Rf*
h���}�1h��$�m�q��+��7�^uC��0ь��=��Ȋ�������dV���AD�����N���*<����3��$<��o��,�y}nʪݚ|�}��}�gin����ז�͏:��eQ���=�?B�WPq9�-:�$-�=�7�XQČ���]=Ψ���Io�Q3�Lf7����u�u8��˥�"_�$t���=��2dwQ��}?�~c�3�Z�Aޅ���S�_?Uf5���;�@�E�[b�}�Ѯ�uI�0����V6��WH�	�U.����L���~U�M�Wא���ů�0i�{�yjS�಍<&7`B��]~�Rg��f+���:����\�v��'�pm�����:�g�k� \�����Β�׊r��	�I#\$m��mF�Hy\7�K ��,�������#W��C�G~׺�_�V]��?7届'�阑0�8�ה`�=�-�g3饳�Q�5D|����Ϛ���A6�z�b�Z��NL׉^�J����:~dxϗ	ù�\"�P~�|�2���S��ӆa��ITQ��qZ���Ls=����{B+M~Cw
%K��j�\c��g8EbV#�6� Դhp�N7yC�H�n �D��;���xq�\p��]�&�	�U��dSc�;���
Y-}�h��trÆ��j�ͲaäVםHj��F�K�1��i�%}�<%v7c�a������:�a�dօg��Y�<1ơ9G$���m{����]/Oq�?lg��S�?�!&{�?[Ո[��G*��"���L4*����w��Õst��Lb|��̹~��h5^��3g��IA����Pu9��G����e۾�D�K�>�GSں���Q_ɶ�d�7ԛ[)	h��\`9B��L��"�ɽC_Ra�v¹G[�^zj��g�ŬǕ��!�� 합������_��Ŧ/���������V�_�D���C.?f�M�[��8N��j�� ��Y1�l�r�c����O U9������ژ�13V��\e$�E����A�	$<>m�M;�9��1���e��)���tNt��k��{N�������nG� oewĉ����gr��tt�3f!���/������-��SR�ηJ#t8?��(�%Qa���� & HM�����Q�6B<sCf�I�{޽b��E���ʁ�L�|�������^mr������=�����"r�ˮ��%��v����=,�l[��?U��r`�R����A�Qm�sٲ��!�cF2%��O�,�)Rs�PV�O�yܻ�RiR�~��o2������$�t�.X��ᶔƷ���h�ʴ���I�z��m)���r��m�D
���A� �]�oh� y$��W/�#��<������~ ޓ��­�Z�:�w/,�Z������~`�[��#�U{\���F�d;:��Ӓ<P�|Z�u�9���ml� [���.�A#�5���^�rwN �)�ф��Rg�⳿ۼ H�N��G=�������
c�۹.T��6�Ǚ�܎Q�2vM�d�^璧�0�9N껠2?n��s������ 2:u���j�XN%h���'���A�ɒ-���\��Ż}tp\�*,��B���%��y�(?��(�c*1��,��/�:DJ2���ܿa{��#n���f�u��pI߬�V&<���֫hp��.^�P�U;\�1��Nհ3���F%\5_,�%���D7Zp6r",�?b�@���?O'�h��0-�|8(��)Q�&-/�Q��#��#<��U��:��O�	�S��t�G����F�=�Y�����1��eޱ|��9Ch�L�o�p���|J�:�[�W�O�kK�WO�a�_�����^��|	���XdS�����ℑ��jQJ�!�n0��_7�)c�2"� ��E<���Y�'�váL�i�g���.D�Vşg��gd^�G��p$�gVxa1�ͦ�)�"]�X����L���|���P:9q[5�M��E�%�{|����7��e&w'��Tn3/x����M�����j�/Ћ�u~��+�����xe�ݱ�> �ZX��k'�����S��H#�S�'`N���Ib�"�֤ѿ?E�z_X;L�]�ӪU�^�Y8Ȣsb2[���`����=�Q�
�b��y����9�A����]"�o��֕'�wJ�(� ^'w
b��	�B���1��꾘i��Ⱥ� r�QWD ^���9\�ov�&���v�7:S�B �^�kF����,K&	�G�2�\F�;o	=��8x6��;@�D��us�ɚz`A�c�K(�!�4�(ɔ�êf�5�IV!�O������p�߾&�]��u%P&#��n�3��	
l�z��M��I�Rz�N��j?{�z��C1�8��ǅ+N�rB��,
èh%��r��ܕ���0���ać��#@�C�.�F�֤�8���7�������l�U�Q�ӗC���7X��'��"xq"�ֽ��f>m=��0Wsc�pW.���[�Ћ�wzۻ��r�i���d$9�)]�1٘pC'"J��J��v��!4/v�"r�t�����<��d���5S�i���.hlN,5�;e��EY�!2��E�p�ql�w��t�	��a��K���mM�'�\	�s.J]���՜��O���a��+�@lU���+D���3n�trȈU|� �݌��$C�l��p��-};�¢�/�>��7W��x�wk[�trwl���֑�i�	2Ku��ʎV��̪6T�h��ՑE��j����=��k~h�p����)b��8e���:���ڢ��M�@`Ni�o���{+��7`�$�>+�?�Lf�E;��?��[��s�{�`�/�<p0y%�L��h��_���Lō ܺ;Q�l���꙾�L���ZRum�dB�C]o�D��W6��2���"M�rCګ�Z�DR��� ��}mՌ��v�T̤�S^�9��н�)�(m��۸�`�&��jh~ђ�^��yY�jX���k�L���E\������gfv����^ϻ�
��@�]�`�m���/5Af��7� �bsG���-��S
��R�`���r`+f1�$xu[�K�j��;A���_rFO*l�	�J���o��!�OA���_/CA����kA~�l
6�,*��9҇���6Ԁ�d��cI�-V��I���*5k������I��7u.>�W�=~����"E���,뢝��g �	�|?�%��#�WR��A$�T���@w� �eV�s�Rn�������H01���۩^*�7N J�q���&�~�s�NbH4ًQ��l�����M�]�;]�b������^\8*պ.�=�dʜI�R.0�޲I��0��X�d^Я@?H�cЕ	*TsUY�x��+�gF V9z�l#�s����M�!�5�e�H�w��}�}�bH䅵���w+��-Rym�x���d6	�OLkx��W�tT���	96�����D��L�s�&��5|�����k|����v͍h�ӆ�p`L2#v�QS)h��af��&��~ki����o[.M�B����v���/@%|-�Ž����TI��A+�	�$�J�mNǝ��{c��b��օ/~5Ks�����ʞO���l?|�c^MT8E�]w[�#	d�[F_�f���G��,`��B�jjD��ˮ6D�۬�0�Cv���u]`�*�p��Q���K0�XH�U��FK�u>P�V�5_=9�2����F���5�ՉyG��4
�E�?'�ղ���EW�C@'X�ݢ쓠�+�p�U_�IĴ|Nص��ul{�;���#���:Vq���5z�-0�]Z�,���@m�P�����e?��<��\��>'!�b��=���3A���¹B%��������hc���Q���X���s:��jV:h����L	��^w5]��Pd����?8��ֿL�9���B]3s���	}y��9^���9���z6D����n�����p^��J�^+���t�V�Zw�&[�Ƞd�F7a`�=��r����`M�� Ck�7 u�|����A�^���D� ܢ���<��Ho+�xJ�������M+����Y�� ��o�(%�	H~�.|��lA+FOe����]���I݂x[���xu�J���$�>�dj�^Z��K�������s�#�u$&4o�K6��?5 jg�C���7�W��ɡw���?��ރ��1�$K<&�/���|!G:�;���A���	]�$��V�#�f��h⣸_��=�s���'��5���e�g����]w�oN��d~�$�n������T�"���x8h���Ȥ��~޷���r�D#;�j(A
�SL��\V�^���}�6�;gO�_҃>�	#��x4�6��Ԁ�C�U�rBG]BixAa�h�"�R��:r��K����	��f�a�e���4��=�i�7bjm�=@�i�Oս�Z��<!"�.��5���~e���"A�(|����v�EJ�.C� b,�
��`�u>��}K����'j�n���
h;9^T��G�Dci��l�.�H9�=ː�d�w�)�;,�i�u��4L�����%U����@S۪��p�I��(�'!���c��s�h��`��m���N^�!:|�V��%�����9�2���M�1]滞�_I3��Zb���^��y��I�9���9{�����c�?;H�y;+u���3�/�(D�xF9��:k����-`g-���p�O��������˅<J��n������Z�^x�
��v��Й7E8H���`�ga2ʠ�7S�1�����ةx�G�pH+ܧ�>	�����O�䅿�z�E��<�8iV_>ϛq̱��F�iy�e�ڑ/��:AeC��`�n9�����J-��8��<�G|�{Gwr	�1�U�P�[<'k:b�O߹�}��֗�=�:��:o4�PgM�1�����nJ�J�7��m��D�m|�����w�v[�u�,&ڕZ��vqQ�������w�Vm��-f8�����n:��鄚�P�&�L;�QT`B1��䮍��:�"�q��S]���03����Sm�jih���eA�k��r�I��#*������:q�T��fKJQuLTg�
=��x*��n;�X����S�i�����a�__گ؀�����*�(Z%�-_����%Q���$�1��+C��y�D8=�$eP��J�����0$6|��4�q]P��z��T�+j���5�X�1Q"�vT�`���E�Z}Xx�([ΤyyuQJ��mr!a�14�+
gt5�gP\��C�bZWף\E>�g������(�Ĳcڮ�0�_Z{\pi�I��٦!�Tɟ����\  m#�TFg��]�n�91�p�]���VnǑē�$�����ƒ�~(0���K%�{�
ͬ2h�b:(�g[W��k#��1��H!`J�y�w{G�dPּ#oo���-����XS"\��'�iI2n��AT��UAv�E���!vS�2\��Y�*��������L_އWIA�B�I"�P���̼����q�^F[�0&�.�H-�^�V�Hq
+
�g�v�����;״��C`�j�i�X����nƻm9�oH��^q7��Kd�f^p�Z%��M�g=y*m��jCȓ��ea�Ft���t>��=g�
����V�������B���������P~z�Wm�XP'#7)�I���ߌ�s��*=�d�B��G� ���}�{�Z@�����^h|�Fi��K"Ž_�����Y��O8Qܣ<�'��l���eނ�0n>�#�c<��~&5��2�|YA҅m�w�,�J���jF6���AB�鸧�����w��+)�����\��%&8?��d�=P�����靡�s)T�A�����J�����Y�Y3��R*�S�X%ҙ�h����Gҍ����+�i?
�&N�\}�{`���6rE>�4P�Rb�O��N��8^�{�"�R������[�(�~��A�]�:3_�n�L�/��dI�nr�	��U����pc�m����ᚙ`�Ӊ�K)�#kp�a".љ%�Ƌi1>8�_��<:��	�h����`��bG=簶�U�=����`��@�[�u�$(��:���o��p��[J��5�)\?\>ƔX�K6`�㿃�>��	^ðG�l�9��S���?�bcS�dJ-�ǀS@
��Yݙ<,*D{һ���
ݛL={S���k��|�@��M�^D���F�z��[�l���z=0�B#�R�P+#	�yPe-���*a[ʂ��6�8��Vb��;���rc�}ྜྷ�����&Gτ�Z�7�^ۅq+PϞo(	���ܥɌ5܈[C`|�|]�b�nP�����9T�#��BkU,z��{���v��ny΅O��2i`��!wf�Ug�:&`D��)��ypcbY�9l��:=�l�q����fW��aKݰ�����Q�ZI|���g�OrNRb)�lU�А>{��|��ן ī	]��|�M-dsǐe��j	6�#��1���xɴi�_�S�L��c����2̡��C�Pہ�L?�L�Ն"��!�EA�kU��Cc�����I�U�L��������V ��;�uJ,%�k����\��p�E�����U���䖻6�G�%G�3t kJ�޺PTZ�:ω� &&���T�գ�.�a|a#�n8��KpGY��+���}2r��Gϲ�W���'��kQ�\	���	V��i�gD���+�M�ZnQG)94bh�:��S2�R��Ջd1��lnh�F��=��s) �*����~
�̷)��U��"K;(VX���9�HJz�*{L������k쭞-��W3���5"`UZ
�����Oe�]�!T3���T����3���4v/��LU�?�槪��W�Ϩg�3ƔC/�rU��	䁶�"��4|�h�����:��op�7&f��g�r�n4Ad���ޯ
Q�$k������
���U8P�6>�������X��G���Bc�ͨF��퓮$Up�z4��͛�������`�F���K��t���� u�ļ�T�7��VY�8SģV�꺋7��J������n��h�F�|-��K�����ܝBK���+_J@�}4o���϶�/!>z��G��$���I�JW�>�y�TE��'��h��lMżh��"�W���C���q֙$�,��V��/�����*�'�艳��Iw�c"���GO 4���
5�y���";f� ��zz���N��A:0�kQL}�~�12%�������k�4U[|��H�}PV� 0;#%)`$�Ee�Z~���S\E̾R�d;%T�!�~��cGD3D�G�8�x��δP�Q�V�'�@�%�qa[p���O���,u�J����â`�yI�C8�f� g!�׭�����]7�d����u�����i7�6{M��tw���#q��wb��͢��lMw0�wl={\0�|������_������t5�K��o6:���]��X��пw�^"��0�+�FsblXY@�3�6��Θ@i����W���0��;6)r�_(i	��ki�6�bd�P�Ѝ����
a����1�[���Tnk��:NޭޑJ���˾��-�
��V����?��+���vБ@h��F��4���}i2��Z����q>~����Cw8�*m�?!v5f�q�l̗�������t_!U�n�,_��r���yvy���:|�"�Ų��o%^�@eU����O��c��Zm�%�a��I��)c�#ѻ%.HfZ��>�n�n��RQ���$�j����pX6��e��� $B6��g��,��Q�(}b�����D���3"1��������O�a��%R����:��ȣ|x�-��g��e���	���A���+����;�:�-H���<��HXa��Y�Jq�������t+�k�E�]z���*�B���{AQ=���]18�{&f�p���C@Ƅ��M޷��F�}��c�3���Z%3�Ǭ�\~S�d���-�w��%�غ#�A"�hս�ٛ�T1����Sg&Bˀ�W�L�*�K[xԀ��ͶQ����1?3��ɬԬ�Э���=]Gd}޶6��5��w�^�>��>T@	�.�Wm�;�HϞ��İ�au�a~��a���0����3��Fo�.z���W`b~d����{SO�u��L��ٞ^Òd>��_��+�$�m��(m�Ŷ~��̸?_?��Ž�D\�j~�@|,ID��*�Si�V�F�������@,X�����0M����΄y y�W���| ���ˊmG����tf��zj���IV���g��V]y]|�O�� ~�f� ��Y{�Ţ(��������"{Ҫ���{Y�F�~�
�?�ɭ��o�k/�E1�(��\_�4I���l�ґ���D��S�VC� .��ѻ4�9��E�N>�Ls�`�����]�43�m�9ʂ��1T4FP���F���p�9��]�-"s�E51�������?(3�\!�EY�l����㭭��8�����8(���@����#vi!Z
)�5U3ˊԬa��M�jZ���h\��8�c�8�sП����"܀�׺�<h� ��
��������	`k''X���Dhp��I�G���ДN��iD<
���[�E�j�T݄Լ:�=l;ak�)�m���Tù�٢=nMkì5[s�d�{ΉIF�ɽ<e��c/WK�(�x�����*@���
@C_ 1����럸|��kyb�bV�=���m�^�B`��	���[���*=�ć�qZ��K�����<�����<����c����M��E[�����43ц��%�.1#}ܰ���)w��ԍ�����]�K�!S����i������n`u0qϏ��2Ʌ7/���|��V\��{d��A��o��G����H�n&�N�&"t}�T�uw���Ǥx�o/�f��Ym&�E���-��%q�܉=<4}�"MTGl����$z�H ���9��M{����6�U+����!�{�V���m�釀�&��iBS�S�yt>����Ф!�:�Tc#�*�t9z7�5�e��d�R
nT�*�}ܫ2��w�X�7�Pi�W�MU��ν3 9���c��߅���i�~�[V"�͏�p�����7��d�!EYuٽ�Lv����xD��)y>VA ��ӷ�F��>��(S��7�B��Vv3�����}����������2T\m�Ż�ᛀ0�ZSq�$�a-�>,��'�(s�`�kH�͏��יD����jo���H�j|���Od�Tp]��B`<{���.~���ء��W��BL���[[�`C�-q/��8�|�&n�N>���B�K�^�e󟂣P���Nɝ�͵����5�b���@�M�hp`�;!�V�#f��@b�!H��8~�<�~���򖣓�EL]��ၭTڇ �4�	
x�U_]��mQ��z��,��g	c�UÐН#��T+bhZ����%��O'}��zQ���>,����踪��\���W�$1"w�M���rr�ҿJ���T��|hHKP9����Zd�������	�شJ֚b^4�)��)����q��/�G,ͧ�C{45�m2��[$iՊ��m��F%�� �O�����h-����	!V����@��0Mz=3O�钇V��pD�T��>��w�çL����iJQJ��������s~4I��b���~;Wl���r]�Т��,�nN�)�{N��f�Guf�ɑ#t�F����q��Npn`N�k��9x�/��>��6�� ��Y��|�0c�#n���t���l3��f �+9��Zl��H�~�]�m<v�_A>Kv{��'�\
~��E?�U��L)/L�{�Z��f�J]���$��`��U����VX7�����ì��2泓@�KS�݄!��u�%�䵟T2��.�y[~��3�:$��F
^�H�j���0���4LK�ђ$ɪ�j�pC�0���_6�ɷ*6�8�0�ѼsY߂0�8�=P����jQڜT;nD�'Yf\%�S@�p�Ȟ�v��2}�6k.�Ӕ&<)��+�e�y<�-�55�!	��+��X�L����i����r
8!���q�<�d_|�~#_�s��0^(�Qi�;N�>u���� G0�^�43���{��?�(�<��n/����\MIk���6̺�:��Ψ���Ύ�u�� M!+������md�uz��f�BPT
Q�~�X�+�����*d{�ǎn���X��-��D6ي#F�(>��/k�Vl�K��ma��2�V�Cu�-�Aku奟՛���q�[
�@�&y�}6ܬY���s,�B2Dci���P���u���:�� 87�kNy�dXEHKe�)l�[G�<�U��+#��=��J��0�]���q��Y� �s|	r.��S@���\1ڭ߃
T4��DH>�h ��P���M4����N{%�jQ�s�B:K�Ϫ�K�VK�*��_�K�O ��<
�4�G@OA�͗o$�ɓ�Fw� W�m���0�
��r	^��i���
te �h}^�N�O�0�_���/E��Q�����/���7�A �I�=?`q�7b����͡"z�8	�ʧ��߷36��~A�=�E�Dn��L[?�QW��5b�;sC��;�}x.�͇�6��Wڃ��N���j��7B�
�ZTv�}�R��l�cUw%d�݉�p-4�q��qզ1�4��lB��[d��]�dJ1Œ7��tk�v��Fp�l��iC����	�y�R슄̉��Cxpy�>)،!	�ߕ��?�X��t�v�?m$b;�99�	hb0�#�~[3�J����Q淎�@�
\�=b��&�:�(����^&��j�8�"򒵻�����(]IY�z�ԫf��2���Xi��A�bp�j�sK7�N˝�6��NҫW�n'·oɯ�4�|.)tQ��W�g��u���n�=7th��m�S�A���`���	�ɵ��xv��+�S���"�J�*��Y���s��!Һ�o�j��Y���3o�}�=���<�g��ȔU.9��(vT8�R�z�j�6����B����-T�ʱ"�{4u ����Ɗ���.�հ$V_ճ�ͣ�~;�xyBDZme�IM�]*�6�8s|��|ϸ����Ӵb"(y%˿WND��䏟��%�]�?U>d���e�$إ �Z��sd1�n0�,�/��78�B��T@=[-7K�zY4�b �V8�f܅O1q��H�adz.�nrOqO4q$(��bG�k�4pM�Ɣ��� �TI+�L9�W����EC'Ʋ�M=C�'��zՊ__:�����쯐�����B�˧(zh1�O�E��;�ۭ������m~���}:}�k_�R�ә�"|V<��"Xْ^�f��+�����<��#!`q��R�~@��i�.I	?�yG[���i��xr���\�џLB�rܔ�m�ު��yr`��뙐����lT�X]�Ok	����Z(��(��ᓼ�;t�AV�~��ϳ����$�����MX@���׬����N�|�H"K��AT�hj�H�;cjP=�~���Ak�"P�a��öp�;���<g����{�(�-9Jw��w!���-�<��l[�B�����m��W�x� �R�qk�/���U�o�G��BJu��9E�PvecY���8�)���VEo+�����wcZt����E[oâIg�h�P nt�~:$��kz���jd]��.JX3I�"S��5���诠;4kƮ��a�I57��2�9�ݧ�$?0���B�&�![�����t_��F_Tȋ���1���k(d��T
��嬑Z�X�|��������c��}�z_e�eŷrŬ��T
Na>֧���q��v���&	���8�"cO=���T���`tϕ6:�Á��ց���P<n�.�X�Dj,�����K�0�W��3g����3,���:�,�G	b�&6*:/��B>��'(Wq�G��h)Eb�BZeI]z<z���q��EmL�
���.�u��6����T�kM�,��&!vc�ܳ��.�B��RP���h��"�Ҩ���*�s�L�1�&=�t<~�|�Nt�,����{EnFm!�y��5�'�j��ƚ��D��t�N����!�	*\ajP=��A^j��P���H����㹞��`!F�j8��ZI�0 �L �'�z�X������b��ӗ���..���6�_��-tm|@��;�Q7?W<��+>��w/G��*��Uy87ev|�=ѩ��sQ�<�YA�Z��=f�r�Ep�dz���g6s]�^+����]����{Ė����Ԟg�C=F<�I��;�
ߛXՓw�wھ��K�p�RJ�B�t��
�ת\V\�1yn�;y��sẈȓ��-Ez�~a�!Qҩ�"˰Wx�c��R�ݪ���Q��3�������e�Yh!d\k~DU���%g���v�F�M���e �K������:S$/���������.�1iNy5��@�Ī.��i[�:)�@m�v��JP��k���&s>Q���ů�+ՌV������Bu��V�Á9�.�1E�k�RP�uAPV�M���}��\Q�u�c�P�Ӕ��!�� B)�#���	��x�iˇ��vE�mFt�*I���Eq��b=u&Iҥ�y�z�&�þ"1I���dQ�UG��4��V6��̀�s4����M7�1���@#lƄ+pRbP'�Z��/���8Y���V_ˎ�&NP���8e���6�g+s����дE:f6	i�1-7�JTa1�Uz�b؊ 6��],d�rD�� O���iL�X���)�a���޹bX{��Ŭ���C>�Vw�j��,���jbt�L���S�3��� �m��FÓ;�t]EX��ﰮ�u�i�[�ɜ�#J�ē,�"UυM�����~��c���ޗ<Ǎ@\�ό�G� T�N���$�p*WL��m�j���¨srb^�Ct����o3�"�W�W��.>���}B��z���q�����E.{Iҡ'��[�-Y�Sa�*;E�^�\cx�N�TL�gOc;������\�~fA����e��tE�8�����~���%��L�ɸOm�3��t���4~��B܁��Zë0�+$��������A��Dm���5�f���^������N�"T@]D����(3/�B�R��4���>�]��}�g���z�~��������Î��ڔ��CC��t�w+�^��
�����v��;�9��:2Τ��(~8�DA�G�M�^��Ӏ�s]���_����o����ׯ\`�Be��^=��	-����tAk���q{k���q�oI>�}�R�
l�uL�+��57��W�7�uի�E����J�yY���Y�<�@�z�y�xvX�HokO�u�L�0R'��[�v�����X����,�[������i%!C�sZ,�S7k�����"{J�S���aأy�Z�ڰ\>���h���|�U��ι_/����䁽���n�o't�;��Q6�
�D�A[|�&#t�[X)�i�o�T<(<�]n!?�E;BR�7�ga��q�y�	]��?a���A����/��VsQc���HF/�+f9��.y�W�@�������zp��g��h����_�~�������OJp�
+�TO��0BW�~���m~B	έ#;�$pD��G��ִx`���4��m-1m���5�q�뎀��� �4�Yva�e����nf�!��<w�B���&�7�tj +�#g'z8X��[��ʰ���W��۸�s�鲩A�\��/�W=v��$b���y��6�⥃K��2�C�'��'O��M�R.�m��VFr���g*6X���&^���Bl6�t��y���   �0Hr�墱�������2h�C�7�E�H���3�O�Mˏ��~�h�,{û��_�_��������!�'���h��¤���1�y꫼P1��ע��,�.��1C���7�,Xԁ�"�(@��.��k9�燩u�g��_�'�$�#���7�{�g���q.9��݆�L����Ef�3a�m�ڽ�2���I�AF��m�2��������1���u�_��-���@�,|c�rq�_�.)H�YzB��	~�$6�,��:V��0�
��'��:���5�L5��RE+�9ir+b��Jm�������o��	��L)�5M��0a+G�a�7D�3��,+����u�oD"��`f��T*��{��w��$�8aڿ���Zm���[���$�'*09���Td����1���� ���������>�PQ�҅xX��Y���b��n|���Ǩ_8`��ک�������"\m�-�^��j�}yS��/;y8��Ppf�/�
_��(��]���N1��]m��,�β��J׆]1�!�B�"�Ԅ��0|���f�^w�Ԟ�S��a�h�ųL���"���ݜ���U�vGq>V~,��o��'ī����&c��q�n@��#_�ڙ���_��	7�\ˍ��/�0�{���sp�/���J[2�T�%ߢ�0+/)4;�b�?�*�7�Eg6~�����#	�^��m�������^�
���(@��2>gD���.��+�i~k�tYF�@R��k����g0��=È�7c�Ju^�5�$gB�JdQL1'r�$�������(�)�]s�PJ|S������������{'����A���b�8��Y�3ԥB\��^�B��Y,��ܔ�X%�`K�c�*6/X��Q��7-�b+�����ʹe��?pm�={fH�=�����T�r=�L����H��_�͵�'��Vy�H�T�R��KCC�e������i2HZ��4�I
W|�c/`�>�T	jMk��2����n>��߸8�[9� q�A�#`�:�~��� 5�s�`ޏ9%ȋ�L�:u��S=Q�<_cA%�iN>D-��GG=y@`����B��dS�LC>�x|����+�LD.�"*=�~nB�g���H�M�y��𝺇/�fE�,z��>��ѓ^��(�H���aɧ�<�5��e�[佴Y`�\����+@<�����h8�2ܟ٨8�:��a5k;�=QT/�N���0b@qfٮ�#�g��A����ު5g�H�������\�/�������8�Sc:3J8��cg����Y�� rNH��F�RXZC��u�[�8��2�`,��z��q�I|��;(A�3_�r��̞��v/�����9������.�nm���6�
=�*Hb�mcfÈ����4Z,����[�]QE����L.R���G��׻�^�ũ/`���A��)�|`�+��.� __��\7yw@��ګԤ:+����Ȏ>JXYof2toS��@���WS40/n�M�������"i��n��Jd�ɪ���6�З�������6"P�a&�i��b+K @]G�X�'���-�.r,
-�D��z�n�����O���z��Bj$�vL�4걢A�7�h�����0F٨�ߓa���2��o��P+�[�������R�x�������U��	��D��(�xnu8U�llJBk��2k�;L��<��Ax=-ey�O�lb�g? #�j�Ʊ��D�s.��".fϬ�j;��'eͭ�cՔ���!]�nU�t��!��ތ�,8����r��'i&c9��.�G�Mm���9�p��{{h��{,~z�H$�� �Na��0�@�|�j��c	Y�����YL->0Wm6|�4�[�s�&��e��j�;�Oi��9\���:�AR21b��S�Ss�5�>m�f���Q`���ln�)�}D��/�V~���ǩ���C-uӾj�5w��\:�J[�����d,� ���x��:~�и���k��9L�,�8��%6-���6�a��9�	�f
Ψ,<��$#���� +/�Q�om!�W��Nk��^{CT/y.C�9��ETҰ��\z� 	g������)��s��9ǆ��a\��i�C<I���`�I�J���w�ü��K��H�`�.j��0xwQ����'�AfA�4;���!��V��>���6�����Qi`�:�g��t�0�rtT��JV�[�l�{ė|���p޽U꺝ԭQ�¡�2��b�8���]L��j��=���0�߱$�����g�;+�����L���I	��ktg'�׻MJ�@��1�QE�v�J��l��ӹ#>��w\�������񫴸�`BIiQ����I{�mF����'�7ubN�o|~�,��������s���@����u>=,G���^x@������R�P(�Z��͓�Wzo��!�A�=�� � �/���X�iL�SJ�F�|l�%�%��0z3���n��
��g��}�kn|X(�{�Ȁ���,������5���n��Pn��I%F�/�Cm���q��+�����<�Kڛ7E(�L(��ߑQ�vj7��pj6��n������d͆y��%�En���e��J��4�%�ٴ"&W�=Z�hC���2����N����~6���Ѧ
� ",��t�����s��w�~�=��&\�y�����D_�t�jw:_��l�v���ė�d�W����t{������ѕ��k�l1��g��9��ς��!�L(�7��x�H� gI7��Co��/�Imha��$�keL�"����5G��wз����i@��#Y� XX����y�}z8�7�B�d�.?b:��7�Vq_�ǫ��̠O�ʾ|�|�Du�\�����"�V"��X��#-p��]m{�΄�����'�87ךA�Xr�J���i����9x�����E�Qb�ܬ3E�N:K��u���K�/WNr!R(�Q����H��B>7Z����t���~��߄�2�umv�/r�K�����BLh,�.����N�1m�+��$�YR��:��r�l��.�M�h����7?�L|#���(!U�&y~,�ey ��<y��mq�)�|Z!�K "�"���Myd��!vE�E*������ec��8���8�#��e�?���A��_زaD�7�5XVf������U�l3���㥪hHy��fpsG���R�������o3��f����k$�)A�Ĳ��p�Wʦy�CP[JAb�3���'a��CH5{�5�c����,u
� ��	9L+��GnES��j0�� ,�$�W#�����bYc����!����%?Q�	��Ϗ��ع�A6/�4����8F6��l�*��(\/�T�A��<�����Y��'\~/}R��B���f�+F$&,�G���x��I1�r�$S^��{��i+��Y|P�=���o
�<�p�I�$��ƺO�6t�n�!E�µd�D�i�m�"��?Y궖94����!����Vކ��s�f�<�v$~o�x�,=�?F�����	�#M#9n��[K�JtBH�*�(/E�c��P�QiP��m���1u�*\4��L���@@n����5�ZI)����uHƫ�����C#>-�:;�7���?��Jp�vq�d3q���*�Q�(搎���H�r� %��$a)p�N[;S.Ґ��u<���.4�Kū�}ڤ62m��\�
�ޒ�J�t�x�%��:uK��-F�C�Z���#u��]�w��7߈B�V�`��+{�6�X>����jdv�_�2p��L�y���L�tc���	��0���TQ��'`e=�හS���+W,}��/��{����Ni���8e��S�Ƀ!�L��\����"w���'-.���&���w�S�?j�ز��L�k��F���w0�b�rn4�r�QZVq��U0K�h��X�o�U;�&�[&*Eni*�A����q�~�Ă�P؄���G񴀦�?�D9����\-�aܒ�����R��*��"i�Q:��;Ȃˈi�hjJș"�B+�U�]x��T�V~u]�[���G1ՖB���xA��e�ݿ�Bf��1��gH��� ���X������ctLg�d�]�?.�:�c�)ˋ���wJ:g�/�Z󊧴(-W.$� �s����v�g0�z+�҇}]��ӳ,��b��RL���ª�L(���[�S����}�*�A��� �K�z��,��;����5I�텷�RѶU�q����H��!����Q޸�����������,�=܎.���7c8>�jU�
Á��=w?�_��%0�%o4���6ݪA����0H�s�>���TB���y�r�:��+��$WW����:�sV8T�p�\'jc P ��L��tB^ϑ��]�lbd��V-�{�R�ú]���zo�6���"Df�^$�Gk�&���p� ���}I(��o	��kM*��u9S���]�Ub	��M��+b5'`���6������W��T?�WnB�7o�MS��C^��ˑ��xޥ�l�2p��:T�J��@�x,�&�L&�+��"L�vl�/d{�yP�P�vC2ć0�ɋ�qi�i��������-��`�f���<��C����-����JM!�[����F��T�k��V"N�'������`���JәΦ�Xl$-����W2O\/<mb�7���u�g��7���$S���_i!兀�iϭ�����<n�T>4�vRԒP��l k��/�U:æ�Z,��P��W{�8�M���OB�I�8m����o�"�-;��$Q�G��t����b4T��|C9���`����R����vh^�>��D�J&�<Wl��sڲm;��N0� �]�7���~�I�&z�eT|���A.&�=`�@{�k�����4H�ケ�4Fp9#X��88RQ&��$�f�����h�:�9�K���	ӭ)Ǿ'�V�D�P"ojU�:� �Xe�R;S�ş3l�t��Di��`Fą�k:�{�o!��*OR��5I�
Q�&���{��b�%cU�*5�v��5��C�Ӽ�Eپ,g�\�ۤ˕�P(g�ا?]\�3z��޾�	����>�ɦJ�'�ϔhh=��1=���~��O��g<���]�a�aAZ[�CF�;ئ���1�!���RIb�����e�FU)�*�zʈ2�	��_|Lف�3gUs�Ȥ4� ���*
���6���%���t)�bZ�E��Ju���5b?Lv�F 5.�Okk��|������\�ǃ���Z�@'�ƞ�x�R���{�cʂ��d�~����G��8�4������\A�.~s�����Sz�:_o�oS' ���n�K!��ul�s�0�^��8k�8��a�N��fP|���0͑uT��I�d��?=�L�ZZi^w �+[Ev������������O�1Й�V��°=��e:�&����3�m���)��]1|s�p�$�ne]c8FH֭�8�+���;�B���2'>�����l�	�~ס�K*m�%-y��oo��<�����5������&>h�v߰��͋����?xS�����/J윑���]emh�d���r'V�O�[��?��!ۦ����~ku,�UbEv����~�qT�`���˗ɒ>��d�+���Ќ,:�����Y�L�պ���?w���T�a��&��ot�T� n��R������ņ*WD��}A������膊��9u2�A�U�/�v��'�2��� �|�]o�JZP ����1B�l�ɍc�B?DǮ/<�&y��|����'UH%t���r��-H#n&�5���'�qjCM���gN��i�1�����hd��\��$gJŤc1����ol��[�(��u�E��z�z�.�I�3`�@������b�&��29�03u���(ة��w�]���G)��l��	�)(���i, �ywʝ���Q^^�?�&'�+n V^��v��7du�Ra��"L!*��z� z�n�r�~X��K/Y��\|���]6�0��G���f'�ǒ3 ���va�;�x
'a�+�c"��� l*��u�3{��ֽ_T�d���7�q�͏�`�?5����=4
����+a��sf��`�!��s4{]�7?��}�n�%~�Z�����@���\-�Y���<���5��@ע��G��,T����C��sA45�X6�x
�ڙ�ܫo��&U�s�0�Pf��E��*%0����s�a�_�sGq�� �	�U��(m��[�ei�r�	����++߲W�+#L�n�&AD���Ae�~�gG���t//aE�&78H5�-]~ρH_��1���,-�6o���"���u;h#�oy��e�^�N�[uV4y�C� ?$<'B���2_Z�f�=�|I�hO����#���#_[�����\����v�D%��Mr3���g�V1������⫋"�\��*����_�+��>���d�9��J���D���. ��>p%�JS�k����A�w���=�OK�b*�����ߔ���#v��ATN�R5�4 ���x+�g�����u8���D"�`��/-?
$�t����Q�

?��k%G6 �'�Q9�:����꭪���|y�%9��Eqo~��=�m�Rp9�@�pB_wSS����ğ��+�C����u����@�� sN�1y��������C�^�4�70�nKnM�ɧ�KW6ҺŚ�w��QI/�~��>��[Q �@����&~J�k�mޙf�ߚ"x.��c]n�`�T*��ER�����v��#��'�D._�7G�a/��=��v_.�2�xU*#��`����l3kr�Y��r�Z��۱�2~uV���7�v�{����Oܽ�݂�ܻ�������P�)s��Jؔ���Ê��)�_��Ѕ��a��!�0_(���7���$0�X#���?��hR�XƂ�:�f�ߛϔ�R��*j��E�ATƍ,ǧp�7�#���}�ljw�p�b����\��:��`r���'���"��u�:eUi�L�}�J�c��qM4ώ�Pq��!؃�0�](1?���S��]
5pA����v*��pԷZ���b~Z �-h.��@�����y�iz�;b��N���bP�7�|��pԯ«}:��v��HI���ߐ�'܆�g;B!{����g7�`�B$f
��`BǮP�D�~�O����#3�R�+�us��9Si�o�ȏ�3�l.��t�7'��<�����V4�U"�h;�������g��q����ryY��5#���m��z��Re|f�
$e�z�͑��֊މ�J�I3�]mNI��xZddJ���l $����cF���]��z:F"��5�bD�&�+����}���֔�޸��kfQ9឴f	�zi���g|�G~5�#����+6�sԒ̰[��
XB���|;𠙴�X�\l�����([�H}����v?<���]}�b)�4P�o�h�{���B�J���K�� Vz��NŅ;�2�3�I�X>rޢc=��/'�πgL�^WF��{ Yc8�ed���-[�w j�J��d�s��;Ҫ	�A3������x(x��a[S��f�~��B5�{��6G�׶1u���!<�\��-��s��_10NS@�����ޅ�4P�N!��B�WFV>�b}�,�C����'�B|S�l�<NA�|x�f�F�8�;����l��pbY�c��-�+Ǫ�[������x�3�?z�:u����L5��(=*�3M��i�������	:I^S�s��Y��>��ˬ���9����@z�͏RJUQ%�l�0�Z.�����
��0׍o�O.����!,�&�M���P�����$6u��6��Z�_��gbK��%V��%�Q�8R�5h:A�7@��E���$�>9���V�d��߻暵l���]тёe�i"��X4��fޚ�/�����n?�)��c����~ *��E�瀆�"L'��h&0t���U����0��9�d]qH�j���԰K��Ng�;�A�G�+ԁ���\[g_����on5Ȁ7����J�>�H]普K��tC�.�jG�Q�f�
��H��� �P�Ӈ#�E� _C����y�A����S0?�\�� lAW�j�&����Ɖ�h�� �����|�3��ړ��m�|w�BX�Z*����4h�|��nt����ͥp�h�-����,|*��t����ͱ|k5ߑ{�vQ۟"8w
L*�jZpo4F��`�M
K�`_��-���,AS٭�mk����Ku ��<O�_p�18� �S���ߘH��ذ֐�N����t6�,��	<v{�4�*�v�*t��9O~��k��]�s��w��0�����r���+������l¸��4�[LG�m��	
�8:)�:����)̘��dþ>�O�.���6�lʜ�@��37�D�GA����&7f�H:Z�g?0:���i����$T��X����
�x,�uB��im����(�$��`�&� ���?T�M�f��N���E)/"�ﱤyz�"�~��U.��dc�o@����_���^���[T��J�,S�s{U�Y� �8�jwѷ,�*@G����h�]�AnA��s՛�~��i��<���:��̑�K��e��\2V���\�f^�5WOʆ�4+������X��rDս�{�r�B��i�n����4����<���b|U�R��[̘.�<�4T��۵�^��k�E�H�c����6���>zxa>0魒AG?)��Dq�I|�V��.��L�������j����t�5�P�G�"����i(B���c][hҶ�Ŀ���q�zV�Q�'8�ce�ٽҳ�e�Q��9ږ�ۂV�ðl��!XE)CG�[�&um��:�1�Ry<H!�7T��J|��@��d�����(B�Q��%�w�.n��i���r:�\��Dk���-ۀ"�@���h.��w��ӊi�����ʵ���U�2.魡 ؀�KT���7ŊeE�<��!�����S#K��/�X�X�VB����Wc����Eļ��+U�p�4�l�T���Q��%.,���ybm�z} &1�$��9���Ű��3�P�}cʛ��*���s�#��ps���hR��ό�˙y�μ,Þ���YL��(�T�{B3?s��0,P����w���,?��!>��"���G�� \`�+]�Ͱw�0�������x# &�|��u_G@ߒA�ZB����Y�3���f��-�����������q�ø�p�V"v�hѫ��1��i+���M�;�*L��~F�g�"�I�i:@#�<��3X2yaV�Ƚ�~o��i��(�5�7/ҫ��ˍ��!�]�8a�����`j���5v�C�	/�y7�!�
�����ԣ����?��M�VyÅ2 ����Y�Oׂ�����k�����p��u͙;c2�,��R�����X���w�{ө�#Ѩ]�x�΍&����a�5F�u��9y�u�/)
�@a6����.�q"�E��p~<��Q��2�(9�3�R��é�09/�Wm�P���Vr2�����Q��������>�i�Ϟ=Y��6#>�����v�H�٥ps�K��h��q�[����=�����6���Nag�8E=�TYJ��CS:dg-Ne�vUo���Ѧ�<�՘N�g$O&�v�7o�\�aK��c\�$�c��=�*�֥�N�]��Z_�Sh�25���9ܼ8L
������w����a�L�������6TSu�{!+iK�*�x�+ C���z�p�9�gl73��B� � A9��Y��#���diŉKq~��+�۾�py]VyYC�M�I`H�^�}(14ID����e�F�,^HV�[^4��Ing�6���s ��6W�wL�!��2�P���N�����TՆ�ִ]����MFw���}�4�������zR\�a������
��*������.9��ʭ`��`q�y��U�+��J����-�O5&�	T6�]���L_!Lr�H` �aW���tlы+�=�-1���>u����1V��3���糽X��M�����%i�AN������7u��Zg�f�de��>8p/��}����|��G���7��m�W��T���,���}yEm l<�N�&��$�y����%���7�bL���~�h��b�;�]ޚ-s�x-��4�p"���+b�Q������?�2:_�˿�v�e�3�nmıfY�+b�~t�ǅ
;��(��� �P�:��P�=ξePoYg��z�ƿ�3o>i�-���$��.�����<K��/��{4v`g�}�\�Z��
9�߂]n�)����7�?K�Q��~d�TR��1�8Cޮ��+�;s�^�A�Z��E:�n���(�])P<���,��}[�b�%Fvۼ0x2v�
$�t��0���g|��`�/�_4�N�-Ĕs�l�%�ᯚ)|Qq�R���+槒
B_���-��R�Gd��J���$=.�����z��Cl�+D�~�h<O�Y�xPL�Wx�(`g��.��%Y���%����ߊ�n(�,�O��9N�����'E]��)�?m!���MF�}�l r3����E��ؗ�C��g!QD���Մߞ���(�i�뾛�`~�@JG{J�=�D�7��^7�	:���FN�bo��Ճ���<�&��E���z���>�ҷ(���n�|{^�z�G�g[/�sն�Oh*j@ȏ��6��Z(����;��q�D�Bҧf�&�Aa�EF3}jm!P�P��q�E쀄�����P*��cH6J�Y�~Mϡ��h��pO�P�Z��|��
���==�h	a�K��jk���~2�F���ȲoI�3��)��`�L�蕲6|����^�H�h��I�g��O�N�;>��L&T>A��FS�R�C�F5(���w,��Z�#ڥ����5�[�mF��i���=}��lR�n�3��9�zN���!H�Ap1��DE�U�pG���U�����a� F��
sz%�X�ǜ#'���,���'Z�N2��'��@bh�g�#7q�����Y^��� *]N�A��	��4<��g��:��OQ ��S�M�h�p�� �W�/��8�K�~r�g��7.n6������la��g������9��)"���p���J�C�D�ʜPloY|Ve�`R�%�wB��u����iI4tC��s5�����I\�3U����$x���ƀV=L����f)he� �(���,c��C������P� ��?�8�8�Pu<��U�^ ���$���w<6�F;�Z!Q�k�>��S�,���ն��L�{� �T�ȴېl��(N�
��,r/}�+QO��4Vf����U͢�ig,���R���D��i6���N]�5刾]�x/��n��f$�Vm�
ʵ�h��<R��&s,RPTX�?�o��@�����+J�{���x\t�'Yg��K�S]��T5�ߊ� <$N�[nΉV���A"-�l�b����3���$mSn��%p�EWB�r	�z�r�Z�#a�J�C6�
���7�۱zD�i/��*�]��~ ����ۏ^^��4.LH�����FnP�Y������.]��F)C����M���a�`����ͺ���0-��`��;�\.�1���# u/�XF۝Ձ��{-!�.�R[\���$���������^)���E1�m�y�o���-y+TN$#]�8����M��Y�e17�=��+?��\��vW[;���b�J&ƯW}b݆�%n-�1jy�?���h������m6��e���t�F���b5�߯Ô��=e� ���ː5���
g�(h^�����S
S��Đ
"�F��Ϣ����}�׸V���(�yΕDi9l��&U�iu}sp�WL��ܑ�j�� bP?�;gyHb�]�J��Iw�/��*��x�1���Ka�i� �D�褧g��vPǍ��<��vx@F)����0��V�߆6o�W�ܠ���Ȃ�� !��]����4٪datW�l1�F̆��p�=�Q	�#�.K�2���[��#mADQm�g�]��해��uF7�����ٽ�<����~�H���׾k�⥑@�6F�ӂ�����
2r�nK�ϩl����PL}O�3!�K�Ǩ2����������>9�*�6�F%&��qI&�#�^M��}G�]�v�I�/�+\o7�o��D�|�{�2qD�X�9ڣ�]�m����f��'����B��4ӕF���C ���"����l��|p^�jz�>��d0��:y�i�C�
k��Oɞ�=YM�WRLa�����C,��x�.'�J/$�U�f�[�?�Gx6���g�,��?�=py�@�m�(�Ձ~����CoZ%��ݚ䡥��o)�s�7��0���;��>V/��}A��g�!�^�;�!�6;�<w��t{��l]d�_�F�W��r����EW�:si�땒2�
�>��-�|�[%��"ͨ��FMG�l����!�߬k`��
��������zʑ�D	��7yv�;%���uT��{�=������8So�	�u��7�wcM�*�cY�=}*
�]q$�<�=��*�4�U��ezxu�X,�壂-^^6es�2�%��s��գ�Y{�Im��AlU2r�p�T�NHmΠ�˼Q`�#����i�պ2�tU��n=�:!�{<��Z�N��n�~�HK�׹��&nr���<��h�j�𙉕~��|W&.�������
�Qnܓ���t���#��8�Z�~ӭk���(oʹ
,^�D/�9��Z�d��$V�X��(��:�Ӡ+r�3���F�TMT�4��&�� �'��f`WK�5�\t�`����Ī���)�5 ����_6�5���ݕ���2�z�O����/CR���g=W�.�(N�1�H�3�H=͑�83��\^��ZT�\�yt�ul�4�?��L����)7m��;���.e'���7\���56�!  �X�����ޞ����//^�h.	�O̪�%���'Y҄�7�ۿʎdQ�����8���|O�U�)�l��4|������, �}|&jp�'����������{ό�CC�!`vu�^�h>�N�n���8QE�c�����E�\M7��M	�	iv����Y�OF���H'�%S]�F?��m�"��6���� Ch�D��^������/�m�����I��,"�o�$�j�S�K�,��}&�`m��Z4ᨘ0��^�u�a`���&C�x���W��\�P�׎.E��nyF]�0y�K�18]�Hh u�,�R)ރ��#h#Hy��X�J{9�1�ed��%�� 3�C%b���_X�t�,.��~�\�g�	��'9v��[ l����d�C���MF���Q���m�
q����,�7�����������/Uf�ɮ����gn���D�=TT9h��߉Td�\lGE�����/d��	+�f�/r��b�|º�V�:;�ӹF�y��F�����$���� �y�c~��:1(3QE�8c�ۡ}�v�����XuC%t�r���wr�M��U���7��.v[��Q߸�Ѣ�_����7�}V�O{�����wԺ����>���U��ZA�XO8��w�L���+�O�}�Ƕ��>z�o�0:5wn�d���P�ҒU{�gA��ۋnFŷ��8u��,��N�}�=�ƐP$�yݝ&��]z!���g*sO˯$T�z����ҳZ��w�9�]��/4��D�|�=�BM^��|���8Æ������[�X�^=׬����q�ت�@���v#�E:�mo��$��NV�f�krOy❭�����Q0���I��Lq����E=�neu^�1(-$��
�i�n�o�Z�
ʹ�m��o�,�ʓ���=���ӂ��J�?�~SV������.u�`�A�0e�	�����A����`�-��ޗ;Ler����<\��/����spȖ��:>�m,�X� J��T�;.v{┈hJ
�3W������i?��oݸ>��t�2��y0(�]Ɣ�O��k��P+����r$��#��8�j�/�\*����m�T=à��g����<$P�~�d��
�J���نcƅ'��5$H��� ����٥� ���%)��D·���(W��=3�-�i�&�q؂3G��\�QX6��Q��n__B�T|��|I3`ܗ$�Gq���*��~yC3v|!	�|���c^1h_��Vų�Ǒ��L+�9g~����@����R�b	�&��H����3|]Z�D��7Nyϡe=�U� ؛�@��O(���0U�Fa�"�/֤z`i�p+��"�]s"&�b5nT��l`,`c2�e��Z:�#��oRE���"�H�.+0�Ys=���(Ǩ5����q��(�S��;'�,L��� ����;k+R32g%��c��%C��B�8�XU�C&ܒy"2{�^7�"�^ ��k�����k�!�YbK�R�f� L�A��/A���<k�΋B��.]QeV��ʇ����a�ȩ}v��� �Qin�K��*�Xa���G�'�8�q:��SW�G��JM���|�n�z�n�����5?�(I]���Ǆ7A٦)�}=�m�.�)��6FlSr���e����@�� I�``qo�ֆz�'�nֹFc��J1ֹ�᫛
�Zj�I�N:f��T&�Z�7M�@��|�I�U�m���+��c��j;���m�f���ob���^�-�/�|��9+E�e�����������hJ��C�p�!�=e�(p�)9*=h��J(�F��z�bD��j! ������	v�VB�K��7�0 *� 1�tS�������Hkz�R���iW\ƀ�Q�F8o��6�Ë��WaL�g�38�BɴV	|$r��4��o�p���	Oi�[�싴7�xߥ2���'4(Zw<�vL�s� 6no�*#C<^+��9�<9H?Zc�7�"T�4	�~,�1���FV��9$h�^�>���w/!ȿ�P<�λk+��aݔqi�-�Ф_��ݕ�/�gO{׹T'B�w�2�
	�:��}R�Ҟ<[Wp:�(5���6�}L�kنݍ/�e.�-=^��-Ʉ9\L��`I� �+/���b�O>�
g���
�s��3UyKU�%~����e�9�1x)�|�y���{��Ƚ%l����Z�]�:��=��0���c7��@��2{��XA4.���6�Ο/Q��#+Gט��,;kԑ5�>x�G����<J�U�銄zB�����u��b��)]�S(�����*R_'�#1�2��%�ۿ�/|�|>���"�/�*fE�V�)Ag�3f�竞
�x�PˈTT��L�~�U'C���Ԛ��x�,_ <���}i�!����y�w��%K���I~Se�6-=��t�(��\h����3X#g�˳c�>BN_kյ�_�.��xfܘZx)���m���X�����`����L� �Q��V���Hm�h���' ��O��g����u��ό�wF��*�s��^W��HT)֦T֨�:А(c���U���ea�XJ ���Yq�=I�ݩ�$(�N4�����.���N���s	�(4\s$�_�nA����L&����)���h7P7��Z����K\2���3��	��;q���đ�Ii�`e��2�b�ͧ��HD��Ч�hzY���"q��٠--6pDɸ�֕%1����. �\cK���E�Җչ�s�y� �!	,T'��W�������4�)NP;�C���wYW_0AɎ%I/sC�Np<��ZI������<R��z�[�®&���D�ၧ�/���C�d�!��֛Z\?���\v"�� !�l��?}o��]�QQp��N�ٴb_����|[i�4^�7��)t�Ϩ�_֐N��S��.�G�_�K��o��o� �s�ٟرW}��h�WՊ��w��J���t�\�B]L����fK"c?[]4�q�֎ɘ����ۀ]]��ġ��^�F=YرDؿ�-��Fa�Y4t�9q7OkUp�k�9�/�+݃�25A��J<.��
�B�ď��#ť�Vo����5#JG0�P��������[�����d7��6B�U&�V��Y�m����5[.>	��i��9a<R7o�a�V���_�:����&|BC�F���L2�"�ݲ�$FN�F����w^s�:�M��fP��+C��')#ؖ��K�E�_�ir� b\g�NTm�>@7;r�+j�JلB��D+�~���W�|2�ǪP$S�o�hf�KK*����zn��K=Et/PO�ɵ�'j����͒oX�7�䐈��i]�ox�ؖx�T޵Z�� �b
�8q�#��o~�'����w��C����7H��s0A48�gϾT��_��3�y$�|��AD��et-�_6�y�,��|IV�tS�P��npM#K�*x�}���hJ�
�9���(��e�\���ɟ��|h���-�1��{���+�>)���Y� ���M���	���<���~�n�0E�Co���#�w���9}����������WL������r<�*���j8^�ff6�ڔ2w'��������̑�Oz��~�=���.���$Y=�㆕X`q��h4�#(A
o�S�+��L#c Y\�ǥ,j�-��$�$3X��eO��l�צqac+,yo���)2ku׶��/���~���O.
.�f���#�?nr��� �6�-��`���� S�V�|#�
�+�Y�nԮ���D�����J����04���f�x ���E���c2�j���;�׭�������[��@��Hry����S/��P.�^��I*��Z��>��_B�����w�kSS��QvӦ��pD�,��ɤ.�g�{>�K
� Q�::GUt$?'��+�%]$�'א9�k۲�!ɛ-ﺗ�d7��n� U�ٴ"�r!7��
�3�ܚ��2H��&�Wc���i��7lD�	�i�'6LG��c�NJ&�����
��๑$H��WƬ� 7^�[-@�����=��-3E�)�Q��� �V1�
+=��>�A�\g�O몵�AQ��������|;� T�9�`)Cmr��[&���j��I�;���;;	DA=�]z�D.��tv�.ؖo~���B�E2�+7���X	�٥gٞe	~	��2��Xu�vV.��r\�~A��
�m�R��Y�~��{��KpM'�wN����@r}j�So�� �F��>x��G�V��G>v��������wrG��P�L/36/�a$L���#���~�=������W:]���B[]�p���X��M5����ٗ�å�"�� �^Tw �!ͺ�ص��"�o":fI握��lQB���e3�n�0�r׼�վ�g�e<�^��/��_��N���L�<( ��FL8���茴z[�e�6�����Z�����fA���x-���0��!��'�Bh���i4���#��5Kw��-?V�n�ӧi�	Z�h�2��*�s���U��i;>��]�MIIR�ʞ*4`ºV=Z��K3�V��M�{D��fj���Ը`�o����k�bm�cS�꡶�U�0H�B�-!?�PHP�	�������"�em����_=��� ���Z����V9�vZɓ�����^{����~VعTv8��F�{�7?@6�n_��[摂2�&�ͺiޡ
�K�#�?��{��,�����#�S�sNb8$������oG.{\P��b8����\���#��R.lL��	�ۊ˕y�S8x����5�������iZ �M�2��-����Jcʨ�i~ �>418kE�`a*�Y2�Db}�$L���G���_W2����^�!"{�qƃ�)Ut:I���خ�M%I��IƜ,�D��㮞�EԼ5���D����gz���@@�c+���'cS�ad�㦒S�iΰ�z&Ǯg�5����k�뜺9$1'hA��Zy��;�Jra��Q��B�XKB�ۉmY�s���%�Z���e�d�,��B�;�?9؝u�;�nh��3N�2�ا��M��J����]Aҷ��3AG�� �O�\�Ҵ�sp�'C���E�p���ld��/?%�����1�r���ŧo�&�$�4��/����R��8ݱK���mĐZ��b�şI]��z���XrXoH8��YD2�7R���K����(�F�1;�b��ҟ�ʃdo)������p���M�˚dPo�<���5��(��*Ȯ�4��(��_��oz�g[r.l{��3�4NJ�n.K��6���%��㾦��Q��t��H��4(�4��Iw���?$7 3������w96M%Α�e�t�n��]�5�$��md}<�d_G����me� ���=y'w�]�H�,��_�C(������`FDF�0��۟]�2�=N�8=�P<�jM{҉���3���C�6f�ꗺ��R��
۪d���6����T�2�Q�d���^��jW�ժ�W�2.��27 �f��G;�)!�q�{M���	.x���R�÷&�����C��+>-�b��hJq�Lĵ61f����;x<\P���}�@���\�ϗGR��4{�I+�����%�Bo��
Fi7�5�t��Ihdb׆*�NT�P��W��CSƞ�)�������f����@�s�(�AD�S����E	��� 1��C��a`��`�%I��mo���'�ik`5���zjƃ*ט�Il�Ǎ�Xf�v������n��ϕdch`�N�6�y\��]em=��vc���b�C��!�D����8���jU�+`�ٷ<4�Ew��e'+�ݝ���$P�~mqi�	�=Y3n/V�rQdJ�e��?��QZ����]��;���W@�s
,���G�|�7���F����g���)�Nх�-�`�j�*a5����7���[]>�ށ���N~��8��]�/iD�'�,�)�	�,�x�#����]��[E=�]����3بA74쨔!�̸�?9g�jl������l�x��g4��l4��>u.� 6
T��*�E��z�S!c3�'�N$���ϕi�tt�����$�6p��Yp�IJ"ON���
w���'�0~�"ي���6ա,q��(1�ȷ��<�Ej�s��݇/1��j:��thO����V�2Dv�n&M�9-��uv�x����855PԶ��!�����tVZ��!��#j�O��7C�=�H��ws�+B$����en	�H;��2�dס��2�e�d%GYK�����Ze�y�G�KռF1�|p��:�3��U��͝�P�.),��K͚&�((f�A1�wm�2_�}�;�D��pmK�`��K�>@��R�l��Ȳ�x�R`���TΊݞ9R�
Lc<������H�]�/�m���,ȗ*����}:�0���S�����-N�>*V@i�i�5,�X��v�S��cXz��*���}R�Q|��8�u�զz"Iw��+�M}��9ZBY���i���;�[�;5� ���V
gQ@~�]������߿��dSIB�0	���R'i��H�Q��yA���@Jd�6޹#�\狓$G5J���Vܓ��A���*�49� #Db��6�g�d-yY~�R�� ���gHn�e�	�TXc��sX�I�s|�2�!�_
MtJUF�����d�4N�����stv����+�<��\>��]a�+��k�X��d������^Q<�\u���#]�����.i�8yo���.S"]+=�G1��(�x���v�F��
�q��볂I�D�$���?'P3����ӑ�܀����D��&�;!�4�+>��C*v����%꥗4�ǣf�DD�jP툾B�V���\�(=T�A�����)��Y��j���w�<'З�|�pq%��Q�]m�Ġ�l1f��� �.�3q�|,Y�p%����t�#��9�o����L�ļj`^�����84�v-��m4��<ejr���B����۞gL裘�
��$[�~x��	؛5���bý�:���#�r���~@��6�qu���:y�H�>?��
�@8�oWfi�݆{�����C�Lv�1Ӹ������+�~B�0"hܱɸ4?wf	���J͜�`���W[2���'�Z�|߈�Y���/��wM��ܭ�)�_U�y���_T�ҜN�� z�;���N��/:�p!?���z9`nu�<���9/b�un��=>�e}��L���D��a7� 8���B8�\
�Z�R��� �?4ݓ:|2["����!6���"�� ��w�����n�ڜe2iM�vc�S6VqcE�u��Ɗ�N�B��sc��F(E�^K��m`lFy��|���S�R�g ��+�#�i@�)�)&�w�+�d��9x/^6���<���H�l'E��i6�Ũ��P��H#[�J���^��z��bxm9Ы��.4ϟ��V)���>��pFT�%��G]02Bh�9kӋ���t�DT����s�&�{���8�/d��tz>?�Y �N�-�c������(������M�i��n-\��v�aw���&mǩВ	���n2����d8�� �c����qD1��������F��gsI0��Э6�m'�x\�.峥ʟs8c�>�4�"{��
Ć�& �γ�`�ן������A�l��T��Hj���"�)��nZr������\�Yp��P\��Lc�Yf�1{1�`+��)�{�*7���++� +�ؔ��5�e��CV�aA>'	�?M�J�V��¡��}���D} ���nç,�V-�Yn�|�����5�8,�m�mӾ;�cI��Te0>5-a���)|lKi�W���- C+�d����.�I1E��!@�'{�Og�6VugA?�gO�Q9�+Pd�6~�uj?雁.|��f �����l�C��`��\�Wն��h�Ѿ]�r�����M�d2:$˅z����I�#��������f�]�L��b����x&�L���	���痿���J��z�0�MiCZܑb�Q�}�P?�FI.ߠC�T�D�+�n���qS����R�Y8�{�9�O���cnW{�`vSXY�jP�)��R���_���~�v{OI˷�w*�t��4:)|�Ŵ��m�i}H� � p�������p���J�͍,�v����6�� 䭀r2���|�3"��L��T�ʭ��>�!N�^d��0T}��&�l��kf�j8hf"�0��$@B��?௕�Z�OD0P�k�~��)��姐���X5ם��j�Q�y������ 	X�֥�L������ƞ����d�J�ˆGɜ\n�Q+=%�����V��Nh�����I�Ģ,ۥDK�ী��3Q%�z|&j-T�ُ����H����c��1�!}�i�E����o8�}K,���*A�^�*�@2.��M���AFVc���!�L�T,P��WR�,��C�`�:aV��8S�	����wq�y�;�1E-�P�Ǩ���-�r�]���=d�T?w'���0��<	�~�%��aì�'��文3�f�}`�m��ˈ� �3�e�
��`���A=�(�c��۽4�Q���'Ɩ����D��M"Ƨ����n�%X[���9|Ӄ[SjZ4xH1F�n�ONq�?+ ��F�x[�����:�`+H�|��nK�H;8���/?�!�r&J�w��_tR:�0��H�V��0N#r#�ƯO��#�Q���ㄍq�c���yLhT"=�/��פ�+���,` �0�Ψ��״{T�|�T�^cJE��2��^�D@��|�HQ��?[�u%X�FP�c?��GK�N�!h�999����%����G_��F��W	��r�/L�-�����t��1<-���Ϳ�9�[��{5�Y�,nV&��g=�pØflF� ;zi")W�PC��,�c��>�R8S��WT�+=��bL����WS�n���"��:J�?����ֹ$��-��D��R�R��ֵ>��F��M��ͷ�k��4�x�g���h���i0�����!O��E���6?�����H�}g���W�~��1ʀ<�X�4J���dO�.:������]� ������3b�u��s9�����L7��ѫ~x�;��u<�8��&z����-�����-3��+8��4���[}+ţ����&�Y�=�ӏ��.���]aBD�[�9��F��|IӦ?R��2x�5U�LO9
�W��2�)�=�ܷ/�*#��cX�m��S)����eLi�m&ɏ�lh�WC[½�8���W�+ܤ�ϒ�c��,���#8����q7B��=�W@�;�x���O�'����-K�E6cI4Q F(;S�w�s{��OS.�fIW�ӡT��l�αXȟLU0��� ��/�}���}�|���T�����v��^�1ױ�WOcɊJ�ohl���#'O�B�V���=I�*C�q+' F��;��ud��JT�bb�,Ǧ�?�Z�s|�]"Kf2SJ�.���
q�|�[$x6���-�<�XjX��� $j�<�Lk�KMw�M���U'6S���{�cX�H�[I@��d���uY���Ԡ�͈�ђH�?_4_RQG��c�+����_�ڢ�	����%�h�`Ċt �ݼ�	k5%�`��~E ���Z�j��t	�Y�ň�U=3ٿDǚ9WQ���3�fIA��X/S�I�$店-2t����"K���T�>C��T��z�������ĳ��_�FV���~K-�|.��[�@�4Nu8����8X4lW�t<w1�ZtՉ��X�W���M�<���%;�w��P�GqK��7����%S��<�Jӆd��Y޴�^Տ=�|&t���d ~H����e��N�)C�ϋ0)��g�s�_���w ��/8��D!��Z~�[�؇��N���e�~��\쐃��ź��F���6���3ְ�{V}$ÆͦC\pD*"Ʀ�hN�"
��c6`�/��"��~��v�G������!;���9 E�������֗�>�ti�U������,���CБ��u���ҡ�gm��"��G_�������8p<��8b�f���G��N�Ma�;�qm~
I\:��WV�-���xt�{*�ȵ�Z�qA6]���g/�~,P�F�E���:�N���ߟh��w0�Aߨ�hB��`�i�5ك@��(/`l$�	�0�����.E�G��������#�������-�X���X��	&J��g�v��}w���jD���5��L 7��.MU!��]6n���L �,_�h8^";��/R����;��~Vd���NoW�h�->:���U0��R�R�;R���Ú�A�i&�����!���L�dR&N��V^���y�/T^$�ծ=.!������QFoU�����3�� =v��i��ȴ��1J��G	0:��}�E��SMB�tW�y�>c��-��p�n�ʐ�[:�r�h�is ��}"v�M�M~k{�t�\0@07�g��e�F�T��X4 �87X���QA�?J��C�ቹ��}!��e��6���� $�B.�k���+v��	BQM���
�B}+_z���
GS�9"�w"a�Ŝ�;���j��w�!6@(���t����7N�[�f�F<� �}�ߐ���
�9����"-�& ��C��4�[��,~FI�_d3�a�M�썈�|/�ڡz��I��^��&�$SQqw��L��9�l�#$ܳ��J���~�ݠ�e��]��t~ʸA7�jR�d�`)F�Z���=���]G�̀�~�A��F��æT?SU�8��b�W.�_>��LM�0Ѥ>�cc�� I�d��񙚷�π���A}V�!le3�S[+)�ŪO���uӌ�xWy5�z�m���<�;������� �����1��I�av)�]&��=���S�&�h��M�l�� ��z2&Y��o0�	���+m~~;=&�x`�YlŊx�I
#ʍ�A ��w�JM��88��/`�`�U�>��'P3���]ū�B� �X�;���CEؿ̲��&Hl�1�[e�{T�C9�l�0o9���♶?o�q�m��˅4<��%�r���&r��L y���\O�1Q^���K�2�U���(�]T]L�|��(leYh��db�m/4?	gkVٚm�kL�8L�%��	UEzK�'!�X��������^�r�4�u�g�gG�7���/��f`��p������C����b�7��'��&x^���K�_mk'!�4H.������b�V���;qT��LhN�=��a��c�S�!������h,iS��AZ��|,^�>��w����n����e��1���*e:0�њ�?�������|����?a�;#O�G&�
����/����ɛH��<Ռ�W�92���W����~�����g��
ᄅ�Q���r�#]�^O̙Q���ya�.�'�d��	#��?3M)	�/KK�S�a�Hő�w��<�����d�yB���	>���7d�"w�;��
�gs"��3>��hO�>"�7i0@�h�ǥ���j"�ɴ���e�lR�;�r����oq���1���e"�IL���C�?�)Ѣgk�$��?:�����i��6��EsWⅰ���{�M���i�(�[Ja��X�2?g�8@�T15�Kc�x|"	�f���{�ג��f��m���c�=ޖ"��= i��?͘�o}]5�e���%�Usp��FD���H:=g�eP|������˸�*D�ܜ�e�
�����f��u[�_?�is<f%|�2�JXXd�N6�'�d:U�������&��q>?�V�T���Y�B=��k�~G��U��g��2o2uK�}��m��tw �@��!���k����mi̲1J��`�ſ85O8�i��XR��,N!�FToX��Q�ٱ��z�Ϸ�U%	lے$�sШ<Uv;\;/��w?��=��u`���	+�����Qw���9��5�'�](1WP���;�$fYB���F�C�7�]{�� �M�e�P���{��d������v~0x�%5yV,�I�O�Zk�M�����&�9�2����Q�Ã�{8c|v������'D-w�Oxe��.h-��9��ۄ�W	Dv�T�y+�N	r�FU*P�g: j����g?�}/�B��oI��h��Ѣ�G�4�ZZZ����I�J�K3p*s_��4�޺�e�\�;��2��_*��ؤ�#r�#�����s�)�á��q�L�ߩ�3D"v`No��`��ұ�鰀e>�)l�e��]����َ�yEnnIx����+�Mu�Ag��4���a9"�ե� #ww�y]n3t
��m5��r�)#K|{]���� x���N؄����;8������tYH�9`Ȉ����̥���m��1�w3\�~*oN�ŋuyQ����Nw^�L��p����aI�H{{�i�n�CI���&9IF���*e�OF�ď"B����6�6�[��˲���1}k�m�.���h�
A7�||A�zjs��T%���ٶ�����H&�-�t�����;9��2^(<�إ���2�Z�����z��nQ&�%��j�G�T��ӭHگ��+S�b��mOʽ�F}���¹"� �)��o#!�Qt�CR\jQ��=l�t�\�oU!z06�Qud^$��ʒ���!�iE�=��F^����{�������	`����5������`*r�nl�u�K��O>���]>iQ�~�OF���Z֚!#EDFB:a)���|���G��!��',J'WX���i��a;��[�?��B��,�m�A0J:/��(aj�wV�&��J���B���!�9r�P<�\��θR�FL�0c��8�|j�.F��/eF�sk�ƪ��%��"3y��GŻW��K{֪i�U-���,0~*���w�v�8�k���T���nx/:Ĵ�y?j����n�oI�Βsz�O�M�=R;��<�N�t��,rS��!-Hn�f���x���L�'�u�ZomM�e������<�7mgTH�U�Ј��s�3 F�K��;\�H#,n�>�cq~�:W�%`��وe91!	̻OI��� �z<���:�.�E묵��H��� �v�ܡ�A
*����5{�>�cS��#��$�h>�=�_���1>R�r�>���슆��]R[h�:�������1�趡XxhO��P�Q�լrY��D��!iI }\dMLu�m?
jbǓ���R�m*Ts�zY��3�Z�W�p��}>=�V�RW����6I,6��=�(����Nhk�@��<�q���쏢<L��>��H�	:�*|yʄ���ʐ�����<�3�2��6��hÀs��j٢h'���o���E�j *�<����~gI���ΡɔɅ��	+���"���$K�t�G�wӋ[��Q�k�^o<�Q,Z��*�ˑk+h��W��ID�-h���f��.�'���)
����?muM5Ţ����".í;�+D�9]U��B�^��ӕ��W.�ۇ?��1�Z�^�j�.5�m3���������MV���۞Z+W�(��9j%|��F}C���o����]5���_�)�����MD�c�:����){������X�w2�p����$�*j��@M�(��{)T��U�9�8�OLq��q���Jw�?̢r�dg�q�Sj�d�w�w��3A;<���Dh�������Z��6J8�'�̿W36�5z�Ȭ�w�^���b�ɑ�$8���V��Y�qE^����A8�_��4Y��c0���D
볣�Pr��IÞ����Qd���U>����a�vw�Y�ш��˔���y�\��;.{����q���avۋ����1J�i����$�����ҧ��w����!�.�ڲ�����m,|nC�}�_��v��_�Rh�7�X�70�+m+�:�+:*~nZ��EvIW`4��5�4j��*�&�4@��w�8c��w��m��k�KŇ�Wl۞�)O���ӗ�(ۜ8A�*�a`�ҟx�=��gh]�b���ˉl�8+�}��+�@)��ў#E�0�*���R�{Aʘk�֋���Y�e^~j)�# b����)�5(����{��ۂ��=��T��h�+�`]7�:��Q�Z~�㩖>��6u�pҡ������A���"����<���Ҭu��9bAu;�����;������X�#و /W��l��|��%��U.W�Y��ڭJ0�-
��þy� �i����wçߥ��Ǐe�1a`~J��	"��tE9hqM�T�ד��+;��P.`�ʕWl"��T�~�֨wY��W��7�4EG��*r���m��4@Z�\P36-���冗�ǯ�b6���H�G�U(w��Hs�>�5�鰷`>�z~ Ѷ賞h�LjŨ���g41�-�{�-��BtN8M(9����?Ugj�T�M?�P����;���*���e��ew��<�_Iۛ��	�$Em����s��lnDw�����a�:��%�pŊ6�u� ��*���V��x1!��?�"��D ���^���.�!�.�@�۝���&�\�&�ߚ^k-Jz�k�W��P�}՜]V= �P���6���C_q5T5�d�Gɒ
��E�wl����=�c��wBܢ}(0��lt(ٻF*�)�	�萚�q0pڗO�ڹu@�S�(�|�@�^�<����C��]�Z@LevÖaM^��UB�qx��\����i���H���ѩ���2�1�E��6�q~��iB��w����A)LD�0�tZ8�iˆ���5��i�I6��;��H�5�z��z�M��VSe[y��A���/]`����=�1eaEw�!�O�)A⎋�`x���k� �!����	eP��H�Ki$ ���Йt��wlE���?��+��T��b.���M��o��F����Q��j)4��;@lM����!YH����{@KM�4reͩ�Ժ�����.�����#�X�~���b�y]����Zn�и�e�t�[�F9H�ܞ!a�R�:�C�qn�2����%�_v���������f��ޏ_9xT�T��QىK�Ve�׽��!k���徭z�R:�� �4d8��+z���C6N��k����|L,,zCe��VϤ����ӡ� ��D��g4�M��hq������WP`�#D{x��0^�����A��� U�H���� �=>"9G�˚��s�Bd�g(n���Ӄ��~�L�A���Uw`��g>ˇj��Y\�zi&k��G+3K�s*���p��*�i��~|��B�+?��}�����փg&|�b���K9��T[)�`=�A���ʃr���J^��e�o�Y� �s%��Y�7������+@^�K� ���:Y����1�o�-����
�N0A;[�cHJ?vy�.P�y/^�a. o�r��cS|zU*����湜�(=���2���?we
��F���AcfMRW�]O��Mq���,J�'s)��2��M�or�DgW٢��x�#���gsjy�_5ڢc�[p�~���D�Խ�OT���ܡ��ƾk&4A2��T�~Af�c�����(F����������J���	S��Ȯ"���}zm�;UR����pF��KΉ�b:Y��K�0���>���Lkg�������K4����=[ q��[!�+��g{�j�X�U��/jZ���_J�n������z���l����^)4Ecb�W D���M=0C�8.A���'T��W	����+����<H=I\4\�9�7�Y�[��
����=-T[7�v��+���%�:0�Է����V��ύ3B�Ǎz>#���[,8�^��#zH4��G�)}+	��`����	9�G.C�ݫ߃n!V.ڼj�nII�c����)��#��-X�^�����U�E��.���{U�H�fC�n(hn �`����o�����.v%��T�P5C2E8��2���ho����LťAu��|�{�3fJ�ƹ'L���,�LU�q�sH.|�)�f��ܰ��})1�����[��B�"��N:��U���S���/��=�L'�4�&�yM ��y� �l��=�S�0eo)5T-�=���F:\�&ބwy��V 2t/����	{8���࿤�b�߃]h]�s�cbg���U�J7���]��˦��$q��&�.�	]��߲�n��n;����!�}�B��Ē}TGU�[Z?Di*�A<g5p(?H]5�˴y�o�K��o�C�ɀ�1���G ��-}��e�}t�_�������g�g�����L�U�H\Њ��J�Wr���K�����w�ӛ[fC<�'A\D�7�F�<���,/{2e����h(���$6���O��9S�����p�R��K�=��Մ��i�� !�K丧%s��+Q�9�XgU��x-���!*-uֻi��6��%�>;Yv�}����N#�f�*�e�T�8!T)�Q%�pTP���dÜ�:�+�Q�2F�0t
MfG��{F5NA��Ri�݂j �hJ���7���<C@̿#�u&�}�0�_ڴ�����.m\⊤�����/@NO"�we��1yb�8����Mf�[�ъ(��
'v������uz��D����Wn�^���ܥ��4g��k�
T����[~F�[��?;[�N��_�[	�H�&� ���8���HwT��`���2�[a����W$�|�h���e�)�
�5��/�H*o����Tͤ^=']檆b�+�0�&�M����V,�v��}��[3Qq^����<(���t�mx^�>[��7��Z=L6��O���*�.Z�����ٲ�򴮐D���i�6jgp�5��~�{�c-�)^� e���,[5�W>w�kӒ�[�D��<����N
��H�SN Hߙh��u �1�7�:[���ri?ى��>��`�����`�5�<�L��,.�v(� ��]r��������� #�v��Q�{��]�q*g�����y�z��4f%���:rI>L�%�-ZZ)�-pV�� �(�q��18g.+���O��ΩHA`�,#�ixM�V���kX����,���`5[�f��^���`E3$�"�f0��0@�v2^c�1�5��Q����DD�ԟ
���<4b�9���K11jX�-�׋�w��N>>!c/1f8����RK@�Ra1��^�{�Z -��ؿ�K��[��uۢ���^W+WFe!�[�JGܫ�����2uo�n�zNd|��E��(N-^�I�"�6�|��14V\[W �6f�IQ4M�W��etxk�^��Ƽ)Vl�:ޖ��h�6�6�+��L��4`�j�Dފ��P��r��q�J���?tϣT]��f��4�!\
�풾��(%a)��T9mRwv"e�h"�avHB�j�XH� 
T�����C.UA�2�-B��ꦤ���M�j��=��&���΢B����@�e�UլZFi�)	��8vOy����fh��妠�����dy�7��[������Z��)NJ
HÃ`�+И'��9�p��b�eS�H�k��tp⨁ڈN��	��_;��?���NKg#٩���*��h�����Ø�4+kz4rKյM�x!p�ʟ�ӊ���TZm�e��moz��8��ڶ.G����+:��1��!K�h�EJkCJ�8s�L��^LQ{�}����̨r��2P3��Z�N�!�6P��_�j[�;�|�9�C�� 5�!���-T��kx�����5����շ�E�kQ�-_�Uǩ���̂$h�}G�q�_�#�W�o^��	��9Xǋ���?�
5����8 ��T�Ո�:U���h��M	K;�j��4����i�ą�4Z�P���yxi�ڳ>̂��H1R�v��E�%�Q9e̚p�jه&�%M�I9=AigK��Fo���6R���[T���I�g��E�V�?j3���%1�y�j�nI`�$4�ئ�T2W��=5K|����[+=Kn�!�$�G���Oc���Cǩl��Ƃ4���$ �yP"Q'���bt�Bi_�6/��Y����G��؂@g��mG��*��'6��ޅ���cXe���d�a,��rt��k�ٟ�5��9�}�(���<G���m��މ����ݡ;S���jA���s8�h���@N*��F��2�'�F/SȮ�]��T	�^J���AK/l���Z$��!���W=W�� �0浹�{�ݥ�~�e�"��0�c�jIB�p��JA��歛�@��R�~Ǌ$$V*oL6��RH�X��l?�* :�{�9u�����˴��1�@�KȮ��
�Q!}c�����{�Z�*>b,�~~��Eo
I[����!nE�ԇn����I�>�5b�I�'.��X�u�CUk[D�gsZb{;ƚ�.��n?v��j/��]n��<& �P8D���g��2�~�˭�{fJ��ˋ��8�'B Lr���ØY9|܆�?�+�2�T6�W�][7M_��1!_"ϙ��`�DFPK���
_2�؅K�	��8ڶ���<��7r-B���d��O�o�!]o�b�;@p�/VWz~�g'��e㼠Ńd��]��y�E@�+��&�Q����5���3=� ~W`�r�b����n*[���L%0�r���2Ў���zE	�>�Lm�5�f�H���y�H��O159r�2y�s�}��=[��7(V>6�Ư�=�B�p6���<����������=�s{T�ܭ��i��fK0dp��,j�a� YNJ�R�	=e�^�g宁'�����������]M\��e�F�q�Ck�~������܎}�׮]�������!E��M ��AK���Ut�,19��!<�f��"34mt�V���D��iMH;x>*+���lDzX��CT2%z���n�n��i<�E?ֹ��/�+=20?��J�-#	����(�`k/�'ܞ��ז���*��$��f�;�d��-���ڳ����]y����E?o?�� >
�!v�V�L �6-���J-Z^�_���P�_c�TVP+sU퇖$���8a�7�-Վ��.� '��C��+x|���u��l�>��졓w۩�c��g��Y�9U�L����Ak�铀*���IK#|���i��I�����ڲ��g��#6�X��]848~�:9��&�����3�p�9�e{��:(��L�_�*����Wahi8��?�I�})����O�\����"Pt�cӭ/,Z���߸]JQ�W_�(_�\�����"���l�2� ,]��lVa���~/����m����h���!V���ŔD4D�r�����n5���i��5 ���	�Z���̇ Q�Sr嶰W*�����2 �X���H�L ��u��-�u�jM--(����=���O�X3;U�&��ЃR������g��>�_��L�S� ��xxoS��g��~w���V-�R_�Re����!M( j��'y�Y2Ǣ�x&��B��@HA�)�ݍ�ki���b�z�"���P�d;I��a�^�����jdb�5�8�ҋ�����WɵH.�k�1����xI���ƞ�"43�����Kmb%rz�6��a�Q�:�h��XEP4�M.�i��uzmjGR�W'yBF�}ݯ�cx'[��W$�Co��B)����*�[[�+Q�>
����3��vp{��|��Y&,�����m�n��Wľ�ЗۆAI�Ѱ�����z!y�!DX|��X�����j��z�o�~Og����\�Q������Aj�s�O�ڿ��"v�M��{��$��T�����Ǥ��#D���
�I�!c��2�e3O�b�-W�b���最OD�C��n� ��\����t��:KМ�)�^���8Gi�}�ذ�Z?��J�)x1y��\�K����ܟ>�w-�Q3��P�pL�j99��q)͢%vy�n6f������k�"<�(��(�.U?�dbŝx��Ȯ�?�L9O���g�Q�;B���=������\U �g�bnK�?X?��Ӹ)Gˣh��ymfPF^r_�P�����a�sB?�ƻ����,������-�n�A�?U��)���0Mm���,���u��M�zi�����a7P�`&�k_e3>�����:qů|�ļS � �&�N:/��^�(KĐ����:n�N�6��:Tb�3�2�͔+3z
��³�~��&.��MĠy�x��s���Q�	kCC�飠7ƿ���d!0h�pbE�5\�R����8'}���cĐ�OJ���$ v1$��-A�_ v�
��b�훕��nFw�����1�q�����"��E���'�����	򌽠��-_�z�(�O���Q)B "��%�1�(���7�wY�O�PƈZ�G�}T�ugbPĞ7^�3m���4	��MX[v�"�q���LO�4?�X���ł���|�X}m"�J@	�Ӯ���#M� ��F�|'X��ƺ�$�&��OS5���d-j]��
|�O�;W �1{��u�Q�-�FÅƅ
q��iT�5�E_	/��,Z	j�ɜ�s���͓:��T��$������ժ��J=L�n�O(q�֟!�O����A!-US��G�E�o1��I�#�l:+�(K�U����������ds����Od>���V7�Rm�Rp�����{�z��n7H) p5���"5���b�?��%E$�`�!���4s�r�NO)�M��$���	d�R~�|�<h�ZU���dM�a����'�%ŧ^0-��/[��Q�8�?�޲� ���[� 	�aK�7#T��`�����/U��H\h���Ox(��S�H�/6����\W �Sy��]��s+R6B�ޗ���*�x��-��"�U��zT{�|9:πl5���L���3rO��_+#l�+�I6�@����3�����#p*į�� |E��SZ��1Ki�*��9�~Ìj�,#�ڷ�"���ǎ�m=��R��׹�	4jh����-���h��n:��\LJ�D<�K�n	.�\5DS�Kk*-�܅�tU3W�`�g��Zi��c,톁BMR�ӛ7L�� ���D���T����ƥP�E��A�'�t�-����Mv[�p���bAr`M]�5�2_u�d�.	S�9	����6� UL��o�Jܼ\Q����)@C\������CQa�G�ǯp��o��CٕH�q
�]0m�t�k#��׊����,��5��>L�����ƒ�~���z��~����lx�Ö0��+�z�$빼���w1�NT5y>�S�W���t���`�gJ��\jN���t�����1�_B ��wc_�sC>�W���(n W��$�T��=�ؾ���S꫌�t��5G��-]�J��;��Q d6�p)��(Bxk�4���5}7U��u�{J����kC�xAx��"�B��'���߈{o���)\|�G�B���e�T����o�a�Đo N�)s�.ݗ�vxԫ�<�v��4iZf ��2`g��c����m�-�8DQ�ͯSa"��5�{z�.o}��2�K�6��1�ق��S�jC�����+���̦0�W&�j���n{񞄠�g��N�u)������RL�o��8��TBK֊����O?#�`U�d��u-48ׇ�Mΐ���pu�ù�妴�`�|��	�U;k��+�k����8��a���n�[�O��K>/�^f��ÿ�[dK��K e��%���9��q�6H�Ν���ij����Щ6z�=�]�|�.�!z�-�?�����A�WډX�=w�Ľ��4�����ӟx^�D5�Jt�1��r<�PK�度q��2Si'��5%F�<����(o��X�v�����0�̿�H�"=�JY>UT�������EH@� �'�I5�"Zǘ��DX��ٱ����Y��)��Um�8�	4�ȸd�dGlZ�I�(J�ኍ��&G�����JΌ}�-c�ZW�=���n_`��=�}&S�W_��5�C^��H�B��v�e�]��-�h��d	?����9~� ���r:���7uޮ����,����4"ޘ6��>�4�C$���쁨�])B�_���UW��4�m��}�]-��	jH�~؄��>	��Ħ��+}�b�~�H斲0���]ތ���~��D����/tǢ���^c.�d�*�p��FG�.w�˝АL�XnY�xgM�}h.p�� 9Cfp ��*�w�B���=}q�����d(�L}%����HS;�BD�b�|�_��H��9W=�Y�
���N2"mU��&�R�+)TS;}r�?&_ٯv�D���	J�i�����H� � "��%�<�d�_b<���F�p���L��CX>���B"�m�����2-��C���=|�`w�&��^U�Y酮�q6/n]�0R��ؚ���T��%lb(b��Z;`j����fIC"�^0�@F���ێ����`,E�*�K��>l�OZ1�}�{�A3�U����i�|��N4�<y):�Ó����=[�30�l��R��2 �Y:����'�Ab�"����s���7��7���r=MM\3��'.i�����h\ڮ��g�1h^�;\ӹN2����`�e����G�����'��f?80[Cj����O$�5�����|Z{KJ�����aX��-w
77��-�k�ꉷ�a�(�[����U�s��}��zk0o��[ٖ����+�p�}�F�ڧ�V��YLP����J� d���E�QX��[��,��~�d�lG�[��T��
1�!��r�F��6���ح�Z�8���V��v��jL29�i�����6Y��7v�E�f��z�A%��hw$�*�8X���?V�v�]�z�^F�DK�*�,I�U(Oo�֮�)����;MM@�f���㖆s��>�����K��\Ԯd K�Ɨ��iA9(�h��ܕ3.����X�- �� 8e,vYX�ÉIMi9�)�z� �%ds��F���G��*`�S����]z�qt�ʷD�SQ�$)�$L�I(�E0W�����]��wnХ�NM�Q��C�����)s��ssU��Ia_�QH.$����O��/J��j���F�Dz@�>T�:����@�(<d��FW��Ǵ�)��2 �p"௚Fvg����|��+�Y��0��h��ZW��Bw��|�Q��~S�_�5�IQ`
�IK8���[Iiq6��,�'WM����³۹��C�h?Գ�&�O�g;�s����vkF�1�S'�#��J\x�:5�y�b�>����5��Av)�@���Q^(��u���?���5U�2_���x���I@k����>�8Ӥ-���b�?2B~����W�D*hW�RN=�s�$;����J����w�y���P��S�9:\=WV���+8qg3�A�I��'�m��bm��]fe[�7j��_Ÿ��n�'0Vz���R�a��h̞���w�<2�0��J��]*9qh������`��%��Oä��͓����ry��S�j����Hw�,�n�9"\�k�*(m��0K~�`��|�ʐR(���Ї]�b��?���d����a������@�bz-�c�)L%8�v��`Bƾ͝��Qb���`q��o�;R�N�A�i��]��`]���f���y&��>���eT����=���a�r���|e��-�B<JU�b��2���Q" >C�*�lm�~~�"a���7�� �m.��1�ԅ��d$�k�oy;�٢`�v�7��@���Y��������Y8K���<��ǔ�*C�������,+�����}<5d�	 ��Z��_J�4����{�Tg���P7�jo"�c�PQ��^;�m'τ�V���_�|n>h��1��֧(&�N._ڍ=���J����{�(�=jz�����ph\����ߺv���,�X�Iv ��ѥ�y �B(n��S�&4,C��9�e�苚���ȱ�Զ"�];+FS�~�(S��,���@�c��+3�Q��9E|��<�s�h��[ⓚ��29|�ZD�K�.�|��Υ���#����5\)��i�e4��DC�ưA-j�ghetuI)��Ӛw��/up���3Q�C"`lzbSo1�=]n��C�S_��ۄ����2�i^@����k������ǣG�t�\���E�]��#���@�:���=�u�X���.7����p3�>�*��`�٘�Y΢cR��ϥ���V6Ƅ������v�j����<D�,9�\��1�4�~@���[IPF�Y���Ljy�IN��_@����Y	�24��b�:����>,���n����C��u�)��jk�F>B=˓ͳ��T������EOv(���X�o�"_.����	X��J���e��y�el���;B�<J�j3�G��Sj��9��ab�B׼�U�F,rY��!��*�p���)�`Win�+&���0���? ���n*Ʈ�'�+r������1X�37�� ��y�?H�E�;"�p��<l9�<N h���*�A�����I��I�O���N4ښ]f����@0	��~`����so�M�}��Ps~�E��8���C������ěUe�1��y��\��g��	(��k�p0�}2��Ϻ^'L�_��\4ǋ�v+>�֐��@[��̍�ѭ���<�J4��t] ��;������.#�>G�yg�E����r��5>�?з閽���B��c6W���Z��g��٥߭�h��������a���Ԙ�!`��`����+��8z�8��c�jD��*p��%�7	��ٝi���I���\���Q�����NN����M���aVl�|7�`�~�Oߥm�$�~�� ���G<杘C�Uz�о O�/�i'
&��[7��X2�b�O"�0�{�>L����9�>t=�?vi��  �S��)��ƀ��s�$���t���psTPm�4����@��4A�58֪��Ԕ.@�[8�I�&����g�F���4Z�w{/k�d��
z�P���h��wW| �kH1��P?r:���D���:$���U���r"X���κc�� W��.hP����H��g�ʮQ����1�=#.��x3��PW5�Z���lQT�{����k5M��������`q�<��i*N���v��Lf��MA�n	d�P\Ғa�r�����d���`^\���=����Bo���E7,�
��E3Q`t4���� ����4�r���ˈNL�`�ܪ�$^	3���f#O���mܿ�3�����4��{W>'�	9�i�����
ώ�g���%�� 3\�8 ���:��Y'��>K����R}�?1����Ql��*o)��a��/
j����ȿ<�O)y�9�nT)����z����M���z*a�d��W�k 863�ڂ���ۿDn N%�ª[�Z(�U���|O������Y��DX%��9���,�]���5H�!.��J��."I�s�:�ZC@\X��?:�ג�)��bn\Ä`z�v��j��D��^.�i�:d���$�.��Æ@���<S��Ω\�vĂ$��`���b\=WX�����`Gh�f������T������׈^���SW�Y��m�?B]'���$9M#�{��wr�\�����u!�,mǷ�F�G2�_(�
 ����nw�Χ��v<�����d_l�����G��v��?����:v	�$���J�32��-v̍3z�tiCZ�f�f�9U���!�[=�Oy��}��9)�K�T����,8Cw�,�b4n��5��^e����=;F ��Z3�\�G�wD�XU���J�
�췭��w�h�b3�a�(X�u�3�[�����x'�L�˽�]��t��U��a���G����|Ic$hk4V/����B%�tz�C9"�?Q���o���*T��tPP3g�(-��B�� >���I|@�&v�G���ܦ*��L@Vj�}����,ŷ�I�^B3p�6T��*`���@#���Ά˴���c����i���z&f��C%���,��d�N��t�N��Sw�m�"lf����R�A�(���^4�\yiv��p�5U
ѷ�&~
�h�c�j����0��TED	���ӂ����'��HR�(��24vh��������6�5��w�3�!z����d���b�T���R<�h�/�k_�j�l�~�hvÎ��!0����B�[,}5�#���J�e�.S��&���~����Ӭ &ٛ�f��qx�{�X��<�L5���B@�����K�&��L�|�2%
�F%`�q�f����ϲ�|>�h7�o��@�j$C��� /\�>
�p���t�r��؝�|�&5}WS��o�\��ʃ��f�W�-l4j�����Բ	��J�������[���yv��{�@���G�;�n�L0���ZxU����/`gu��@���s��uTkzŪ���:&e}gx�������ލ& l����ۏ��N��<^�!��+Ѿ4�n�{a���8 \ώ[�c�/%M{�Mn����	�&����k�ħχY'�v7��-�X-qͰ.��5�$J!�T!�Z��<�+[4ŏ��E�X���"����p�S�-�n�n �Ǚ�_�>��p��Cs<16a���KNm�v�����~��M��/#�;��F���w�4,n�<�����fB���$�����H�zfSO�EN�|��m�@E��B��	��%p�0�S/Ԗ<����;L{AS��V�BG5s�]�דXo�D'B͜K�d;U��n���F��H���vG�3N�B���JE�O6�n՘Ӣw9mW��9����N&��o�Fhp1 A�lNV%b��5�U����-Q��7�PXQ|�s�VG����W�7�|�m�V��U�ӢP���g��rMoɀ��/��TT�n�\u��6����'_���pTM���c|�uÍ.�͒�o86��
/2�i��ȍ�[Gu�����Eş,.2j��oZWy��~��p��q��$X���˿������g�5�t�/gCAc�A�<n���t�ɱx1�'�G�����,���S�G��x1%�0e��^������د$�%T'4-�Hʁ�%3j�� ���s[�M���2��P/.�I��g�ۏZjZ�d���h<��E ,_=�*"J]A6J�ZF؉�i��L�����ճ��4�����+���f�	�ƛ��\`�tj
I�B��4���˶t�Ft8	��,����aR������%4T�n��Eu|�.&��a��>�</�78�F1���>���8ԯ͍���91�H��&1ֆ�f��E���Gn�������<l���]�[u}��R�?�*���xy
�����%s��)�22�ms�`J���IX23�.1�����q�x|J��k}�� 		4�[��B}�S�e�(RV�{ D/F�HP�A*E.ʯq�a|Ǆ���[�+��) ��=4��\Q���3j�XbQIdL��V�`��u۴���&_���r[\�x��Y_�JH�S�vqU^�t5���f�a4m9STߗ-�&�v�w3=������N��C��F�/��E4A���V�C��i�����(�<�r���'�ss8�+C��F����M.��m��˚y��d�N�m,���`�Ӽ3���-�y��0��@�fѨ��5-x:���%d8��(o
>阙�5g�#�#�-�����$�"Uj�ι夸A(�"i�A�쵴c���j?f-!c
���^~�b��wt��Z�;�7�c�����MS�[w�+��!��J�p��,-��!��छ��:�~�f��� �r{Զ��\����F�RBfO�U	\Y���9/5���/�
_:�κ��Py��Bp���0��-��G-eB#s����&����6%��fM8�Z&�67^\gEp.p0aŊe=2t�U'��4T�����ɻ�[�Y�!�����Gw`zK-��6���0�p�-��J&+�
w����<�$	�F)��I0/P�<H�ú����8;˜M�@�I�)�2��ă"d�~I�����TH,���!��@��	�RZX�x�����Q�7qL�1U,.���u@Z;8d�7����W���ao�O�����1	�'e�y�B"��-sz+�cǤtzџY�������nS4%%�7���َ��I
���v�8�X��]|�����@��e��8Ur�����������F�B����.C��;�*�
��+�M�Kſ+��	'�sY����ЃZ�4>�F�o<�M�^�'�����2��(_:� [}��m�` 6S��������=�Ss���3ٵaT�p���W����q`[)�:�C�� ���rc$5m�K⨽�N��r��] X��f8D�J�0M����7	�7����d�޴�����4�G��>@�Od�������'GU�A�k}2�a�|��ޞ�
����3a�����5����j��G��:E����<i���k���@�'@�4�8������3�_�V�P��r��*����
0��b��T�__mKt�9�Ѩ��9/R��/`� I?��Wh+�Q�(���y����/��	�=92����w�q~��'���	��٥�t�
�^�<$D־�N�].�ʴW�bi[��x�����b�i�K4wBQ�<�1�C������{q��0��?�)�Vv��=����4Fl�����6R���v��"�8��}�hHK֭�'0�Ǜ�ݶ�P�@.��&�/�0���'<�+G��23�G�+�I�ǲqx��+��p]*��6/@26�fc���N()�\ XM�<Q�@�$��-�����<hƠ\�"A�A��y��i��q���*��,MC"c��=.n䝣�fkLcf��SF�~905�¨m����˰y���5f��].�#��/��~��4�4mJO�	ƪ��{Eb^vBڴD>j�	��s&�?y�?3�O�v�� ��s]�3����o��'�XY�TV��4uQ@�]My4���e2b'��['In=��k\�ӆ��Z�9D��l�8�:X7�'�t^�� ����xb�?H_�I�X�ax��'��c�S���;Zt9�
Mc�ʚb�..�W|)�f� S^�QJ�������BK�`Ԧ9�/7�c \��*�[fQrÂ��م��?�/�)"�_�[&����q�%���RV6O!YVY��@�"dm�KA��E9�5�d���,i�<W݅8<ehy(��&t�� ����6����(�*�������A�ie�+��ݲP�`�y�%�[;��3��h��QO�RE*�5}�J%��q�.��R/Č�I�T:�Q˙��8�Kzmֈ����SN��W�4Zue]�FcL6�c�_�"
�t�c�'���E��Az��i�	�u�H Eu[
�^~�@b;R'�T������R�����?;�3��5���M�:�3�k��Ώ�i���Ď��*�+*t DU
D�Ŝ�o[
�XJ-�,���9�a�BM�����^��a�4e)~� ��
��>p�d��0�m*X�4M�X{���`�)ѧ<�C`�6b�`�݄9��6���sW���ЍV�����*���]A��-�FXH���E6�)���t�c�2>o�[��S(嗳������y�`b��G����*t���ǯd���sl5���{Ă�z��w�2�.�x�t�|6����
�Pژ_��o{��O�_0T���(�����"u������$
��F�kmKj�іGcZ(��d����%��T+��|{
�Wď�\hP�5&E��t��3��
i���"�NQJ����X�����1�n��Z�7�gɽ��UD�D K@�Y�ٓt���&r!�0���-
WZ�ז�����Ό�xL��P��	�Qd�r����f�*�M��ι��-$VL����Z�E�$�����u�?���aPf�r�4�׬~8^ُ�3�f�5�2��Ԃ�p�Ș\��C�X_��2����y��~<}�="u�z�G)��])ڡ�8"@P�t�)�_�#W� �kg|��w)͟�������p�
!���!B�	�BG[a}��v�=���D��|�<�#B�y�+,5�4�i�ěF�ZI<B6WX.
�����*�>���5��>=rK.�Z��]�J"���B�iBV�s�d��
�����v��Vl������0���ʃ]�"�~�h�z_�ц�ha!�C[tl�&����g����u�k��ϋ���OZԍx�v�-B_ ��|���:��8\Ԋ���(N~�[k� �np�Jm榡��wx�x��x{2��gmbU����LKE=(����]�Tbj:| UrZ3�Y�9�v�~H��t~�z�b]�bY�^��#�^/�O��u-@�WoIP�����[G�&�J=2�ۢ�A��P^�g3�p�b���$�Z�� 쟕��k�z��D#o�T;�6��������շ]Xp�v��yl*Twj��o��6�F����j}���t9�!3F�"RЫ��g+��B��Ӳ�ks��p~��\�8ȱ���#�pL6�=%[��);/&Z��H~83�R���������3���J��l��}ǧ3��saʳх�*V;�n�0QC�;[���I o�����t��Ia��"������u�J����P��Tm��=;:�	@o���9�FR��.�h�TB4�zF�Vl=��莠w*A��Rc��.1 0�3$g��Y-Z:�E&�o���dt�@��b)x=\ͬ�`���g��8�u�7�;��1w��/&"]Ƽd�^&N����Lao��,�Р�v��.Z��P��,��LF`c�ߣS�=?|��%�fگ�Q��Ro�G�t���-�7[{�"�����1;�^t�����?7��~k�gI�+�܀�4�7���=w��ۚ��YH6��-�?���BG�U�����`�]�4J�t�^oa×l����$ي
+_�2����Qs����6��8]�=�d��?�qϮ��Q}#	��Lܨ�$X�m��V�������u��c
/�)���\<�#Y?�.l�ё��O.�@�nP��09'/����Έ����3����D�w��e�g��/��5�kPk*�)�=�C�H[ΆE.,��8���F��`Z�R<]�Ι#���(���*�g9?�ڬ<� k[%0�s$;v�����u��yGjU�,!�msiv#֦_���-a��.Bno�[�~P�{�6Ѻ;!���u!��r �Ӭ��`�=����2��̕�Nݼ��w��PY��
����ܙ�����;���/����a�)��8F��.�v>�(������[`L"Ҏ\`�)�6�ˏ�=� O�o��b[u��RL���Y�f����͕���]�ܫ����c�&����k�;&ќk�͵��<��H�w 9��j��S������bGc? L\J&���8���߱�:*g'����ke�nY_:C���V�_�~0Q�m���b�E}�ۉ�k�7B��*�l׿�{7%�f�WSZ�'����j��LP�-8��U�?��/̓7��wFN���}�ϐ�-�
�YϯD�}��;�؟B�o��!��E��
��n�kz'��UU	�8�s��(J(�;������ɞ喹�V�^S\���u�j�iš�c�
M��ә�3�P�NQ�L:��l���,ƒ�+���U�[�W�#����#[�S���}�:�P�RՊ̓B�>ə���G?���u�$��r�լ�j������Y"�3f���i���'���{�*����h"~H��T�]����*���L�nM��C{�jCk�wtu��!'�o&mt꣍/Ü�j�jW4v���Q�x���Fm��@qR�l"���ϐ�D��q[�S;hw���V�r��ܱ�������F�0�\�#�yevi!��]��!ʳ�H^��*[���H���9ŷ��a^���i�o�O�v����Xx�Y��p��b�N�=���FGtZ�q�w����F�8�T�EOհ#S��M���5"�^Λ�����bѼ��~�`�X��}w��g�É��M7H�Vf�����1пҸ�x���N�k?��� b����`��f�"~s��*z4"җ���w:�����S��a���wo�GD@��z���o�t�P�GH6c$-�HYv�ن�V�hD�j�P�X�!�Q�V����\���յ#�M���Z��%��*T�2:Y�P��ε�?h��h�;���~���=�� g�q�>��:?���1h72 ^&o���|5��窛�6��h��m ���o�Qa\��ĭ[�c+m���,0qO�a�[��i���D��L�����9�+��)�5���Vu(�˱���p��!��b.Ic�F`�5����sd��Ҟk8�ֻ2�-�տᇦV��Y�XQF45���{#g��]E6t�0,��Dƥ����-��;eb&��u��wv�ٷb%&J����cÊoRu�ڏ��k��c�m{�ĬU.Ji]\bK;��f����l�6���OM�R��~}����M�0
�%�����־��*��v�g0y0!5&��G����;A��h`�:<��P�.և*�������f��}��C�Z�ݚ�0
����ﴧ����!ǻ4����6��.e�p�mջ�Mr\D�1��"����<��{k�'�ض?��o2}>����4�t�u饷�힆]k����󟮱&k1H"H}4bF���c8m���vq���g�?������k�RvS�N���S�ߒ;rc)1�Me�����?�n6驿*ff	��Q͗"d~�:���[U�2ִ�r�9�ʰ�n�f"���gl�K�[�!�$o'X|�:�K�%��NG���2qðMFR�>�W�	����pvݮ�������bk�\�3��A�?e�-�Z�H�D<�{%��|B���ؗߴ���k-���׼vB�pR�A^���c^U�ܑ^`2�*��=:�g���Zo[�Dh�1U#�ҿ�eFM�̐���vc�PP�;B��O��eV���;X��JX�	ng<d����!�4�U�"^�z谆���m�\�􂀐��!R�a��Q�^��P�/����}���Sy�#U�����W�?�n�n�=lY���Θ�힞W�
�K�ےa➅��D���j),����^�X���blr(MF���_<3�x@�H*�UN,y�6�Lq�]�Vj@S�ů��7��eA�����R�ְ��vEa�0�\�����T�@H1r0���{W�F 'L�cл�?���-�j�l#B��8��C�� �qzP삉}� ����t��%"X�G�����B��m���"�NO�o-�tk�A����PQ\������S�n����m1�[���F�$6��J�۠�&�0��W�ؐ���U��]PJ N���5�[֌��Q�n�ߞa�b�Q2��N����*{����E���bh
rDZBTœRLPT���A��LV�?O�E�sM�MZ݀�a�����_m����Z��+�k������l-�7���|i�\�E��{p�U'�//(�#]7��>�z��.��+���٢�����6�:�8���zO�4�s���Y�d3!��Ʈ�ZC'$���� 9�/}KRAB)�}'^o��`�x����ܣ��k�R_��4���jOh�F�v�����"��!�yYp'��Sך(g BV�:�r��#�?�����o�D����6������^���u��g���G8TB����4�2��i.j��*5���n�D{r�t�*��y�Cu	޹���^�f�ȝs>��'�c�[6�CÁ����'�K��h1�h��K:�ٱڦn-�h�NT�e�sZ�w���$,�A0�Og%���h�-���e�+����S/7;b�q �<eOV��b&����7	A�O*ZdX����$�I����Aa6?�0��|�	9n�+
��i��0��f�F���	���Ŝq$̈́!'[�_1�
�k�/��eg�m�X�H��.0Y�U�ԾJ��_s:�&��1_f䏟fP�V��N��$�E�{���(�_�9 �ؖ/�Q��@��}V�h���7Eo���-$�����<ZT{D��z�[@B�k<&!:�GOT���
ٺ�d�(�~0X�zu>�W�x�f{)��v4l&&���cP_����h�.��V�ٽ�Ћ���t��π���U�p�+o!]T3��^�%$��m���;R٬j)���t�VU(Bs���~	B	�ye��I���*��Ϗ�����Hg:n�֊tY�.6�5e\A�å�Y����b@���ސW��!�l�pP%"��W�[��^b��W;iT�w�� Si�i�OMs���^��Uu4�������}�C��Y�"W}�~�~�_����	�JP5�y? �knxo�=z��#�$Ǳ��Q@�������������I{Q~}7���J0�O�F��y^�2aѾ�o�c+�:��BH�ҡ��$k����.��V<{��з�����~��1������tE���:C��k�:�rۑz�d�xep�B�����mN9t�Kx	A��r]F��D a�5m�N=2�sk�{�{��L/f�	^�l�/��o� ��լ�5����	B5�����o�����O��^9V�(�2>�d����b��YB$M g�mu���plÓ����I��rx{b��ܸa�6LSYGi� �4���šDp�Y�<�#F�L�k'do���&��h�qYF5]{��=u,�q$ʖW��V�@k�2z��q�$g�4�����Ʌ��/��L%*��Wn�"���ԥtc��-;�m�����]㡴�{+�@r,^��Ș��U@5>	.Y�u�BR,`��y�Jz;��רQfGn�L��Y��w�TI�j��I�g��Q2}�]��.\�`�k��'1���"w[{.0(�V��*����>��h�X��p����׀�E�	�k��[n]���`tB 	ݭW�E���`a_��G"�Z�����;H���N�6Q�٦�����^f�RrJAm�.)��܀�U
?Ȝdb>��;(��������x�=*"�~E	��YN�s�Oz�ƫu�S��.��Z�>�8;D�l��i\}�d,G���{���g*@�N�Ib��]a.��Ȧ����w�2���Ы⇈�d�f�M��sz$o9�k�G�Vg�+5�Ԭ; L}Sj�;�9	��_�@�^F����̳���zjx�.'9X�]���Nq�����FFla� r�n���LsRW^b}.q����Ў��+T6О0w85��v�-��b���j�I-p��s�/��@a�rE�wV0�#��^ژf�����EY<��)�r��Wڂ����^�(!�&.2/�J���(����"�xp��^r���_)_��@i׮��~��ӊ�� �G�m�W���y��ݨ�e�{���Xz-�sbQHS���>�U� �m�8�u-�K��������Y��YgR~O�m3������@B��j��u�WNR彨V���w���[k�z��-���N����,��/&`���|0:i��\�T�ZH�������6���.�֣K]0M�� �Yz��HY7����{�r�d������t�%��)FY�#�-:K���v}!��^���+�7�G�E���;�$:#��f�V2��yh).����f�#r����+0n�#��� �.H�%]���k��SCc���O�_��PV�2��`�lUٙ!����]~����ϭh����u`A��[H�Q�u�����|x������l�.��@0(f��H-O��F��1�^
vz�Ul�>�b�K=J*}NSԴFD����kV�ρ^:����Tp�'�6�u�M�a�<�Y-�`�Z��@򾛆U�@���_�nU�}Ɔ��Ev����u���������G���.�gJ�x-����-V�0?Z��K��o�a3��%i�Nf�f:`����i���������?U��K���!�i�L�E��Y ��^�'�|����=�'
 �V�jw�j�+"���#�	q#��i�P|��?��GoF�.^%�es�A� �}ƙ�wP#"5�XE��#�i�Xb`���$��سX���<(���H9,Q����8#�n@?N��z[���܉���| `�Ϛ�����*
l��/V|l����3�����SU.:��y�7.#,�x��g)"A4~-��G6��#[�C��w��h ��� i_\+�y�Ѿ��,/��������7Ĝ��i�>A ^q�V�'�Yn����](蚭ڤW��ݞ16ܫ�f�5�w�ܔn�LTFMtg��Z�o��S���p�Q2�>�ÁM����,�۹}�%'��ml[6�	�5�NaI��AZ���H�`�u�����7�<_Z��yLm�wY�JY
f���+��l��~z���=]�p�o�(i�>w43=Z�&�Ȍ�=�ҲOp�/X7)��������7����x�X��"r��6�Vbi7��F3���GFB�qL�e���5��MZg����BI�jf���Yb	&1
ܸҵ]zdWX�e\r���	H�+�;��!����s�*IS������N5���)줙�uW�g��W �̗k�}��μ3�y���� DS�>���.|H�]|�6E�]&�>�L1�}~LG�J�����(0�_L��\���O��,�y�gB��rt=�Pmm�0{G}3WYf����@,��P����1�1�ʩ�|��ڡ�*_�/���LA�f��-x���n����j�"�m�m�s��K@���c�(5�U�fZ�/�U}JB�4"�x6�3���M/J�QJ�]e���1�`�Q%�S~�8o��De����d��y4��e[��&��kW t"~)B��K$jmJ�|a����LDq�'8?�*:`�����������d(�n����"� �a��F��w`�I�4�]2�'M���Pgԧ�&0�՟&a���(��0o�ڍ�J8��P��Y?�BԨ`���-���>�Q�f�h� �TÇ�_�\�q�����Ѕ��%q�Z��?v#�h�ǎ�*rU$ÿ�w�šD��e�Q�C˰NT��������q�9�Z���.�o0�Wv>���a�0�_�.J����.�ɂNl�0�i</R�N�f74���������u:@�6�F�UI��(
Sl�:��x��w���*��,4��m�4D�?Uh�gE1�Ԁ����I���c����h�d�'�gx���]A+<�'��*�8�����J���f���+��L:�ju��iI��3��ڐ�ݻf�P��J%��Ѓ�﷤�F���#P(�{����$�2u��8��8̞�9Tn~�ӡ^31��N�
CGa�4��	��x.�pQ/^� �7_2�J�D3]�[�m��AN�S��A��9:.d�bn�4{A�� @!�)Il����m�0dH*��@��X�4�܊�c�:��rv/� }j�B�V/���j�]Q//�+�����QN�MKWGnK���@�	z>���(N��`n�`ߪ�)w#9��]o�TZ�1b��A*v��nwn�
m�u��L@���)ŢU�
Z�0n��M8��S@hs7��߸�&�r�"mp{�%����.JG�H�����@#��4�J��������y��'�I��������ƌ
Y9=a�Zq��i��;��'�\^�����|~��HMㅂ�в���/i���x�,F���N;ZU��tS�:P<g�A5�a���?���}gX�f�]� �k���I��*"�o�]����(*ޘ�ݫ�4���l���Xs���E�J�f+?P�����)5���w��{W��}��*��B��i�@9&_OlN/.T+$�UbMiY����J�;p�O*����Axi��X�5��Os�C��3�J��I0����ix� M��+a�Ҡ�E�S����#�bZ����ʨ��z1Y^�z�r�_b�z'\�u�"��4��ͪ��'�)-l?8�S�j��l�7?Z�T��8V.̤Iń�Wi�ˢ�H�&Т��ҫY���t)E^���<��R �\:�{7F�{y��u�KN�����
ҔA�ſ��_���2�O�{R<>������?q�`����s���O�/�G�杂�E현t�f��q>�S0��j�mT�]��x�J6�����q�4O�JQ$��'\O�Cpؿ0�ޢ�;�Uw>��X�S����E�rf.��0���Ba:�Tn�Kji��J�s�"�Yfx����V;�<F�S�#�ߣ P��8���}F����}�`	�(���a=nԭ��mtS#T�7��kڑ�\��.�X����k�,
���)�Ԝ��;W�1'��5�W|}S��pQpJ9�l���mZfښ+�2X�M(���P��/�H�66��5X6ۧs�?�j��̱��ކb@㿢�����a,6عtm���G/�l)K~o$;U���E�.�O".�U�	_0��Azp'�žqt-(��P�����nK/GtӪl��S���V���	���V��O>Z�1�c&}��\7jl�FΦ�G�ZE��L�D��a>x����j�A��A�>���)�C!����t��9��#�*~��9��$��!54$ I#�wq����Ts��[[��c��6��մ�!Q��:	&�[|e����w���Z��M���3���9�\*�H�Zݏa2j�Æ����7vQ�LLj\|���Q?ۘ�����U&p;)ͺrV֎+/��!��M� �1Y�h����r �1��1�2��xfOY���j-)��4}�u��&T+z)�N�r(�G��
x�wT3v�T�����1N>{9����h�{k���x�ySY�Z���g���PY��]}3�߫u�/�3����N:n����]���~a&%�%��cl{��W>�&�����S�G���b\<���O3� ʑ�J�vC&$O��N����냡N���X/���<DQ{ze*[t/QÛc�#�u�v��Z�G	e��ˈt�Ʃ#�(�C��:X\h�[=�R�	��0}����F���J�]���![�K����Ꟗ-�P	�1y�+����A�Kwy�:;��"@�y���}58;�h�u<p�)h0E���d%_v���8��-�z|ܖ�V[�0�w��g�?y��<ڍ�Q�_�$��L/M�^X~��n����8e����Mu�he7|Y��[���{����gV?~�k_�D���䡳��8XӇͮE��~�\�tOވ�d��Y;���af �z�:F:�_F�ia��C��s��3�w4K�ʫ����u�S3�]� ����%vq�p�v���R�r��+/]�vh�:�t�"	Q���ه���+nA��6|ɤ���c����=u=�;KN�:�cfh!�ؚ_ބ���=N�[j9���.zw��	��_"Y\4�2aEhS_�\�Yr*�%-�\	�7��T�ֱ�u�nr�e� ���/oDBF���Ή���gǪ�D$J<��d�e��F$�de�x�"�f9"{-���m�0�"Z;�X�.�)��1L�_u��V��A�F��[��e���[I�?�������{�=-�8j��q�����ګ�~E*�b��(M��� [����'PI��
q�����G*�
�P����H��F�;��H��$KZ���ؒ</�C���{�Xτ��� !��8����ټL���0���s��p��y�9�˗wY�d�����Ef�H^3��.��k�;�.L�_����/`�=n�37p%�ª��{*@�{�찹}Ep�x��!	�^�΢���]1�.1��V-;�<��}��4�X�3�O���8/p�L	?9FX�p9x��+�k7� �C�IkI�W����7����I_�S�0"g�����]	�ݫ�ϒ�y�.����Ƥ�Q��d$�C�)�8�Ľ�86V���I��[��2�i����0'�r�����xZ�>$��b�ņ��3s�ރ�z��L@d�l��lwuoCK����1���3��8�`��1Ώ�^�
B�nBfđr��W;��������>�������9t�:��=������wȪ d���ѣ�o��(�|���,�	�Hqa��M����T�&��G���@����(S���r숨�K��*�!��h�.�L� KB��S9~�4�$�Kd�ق~hM8�^P��z>�~�����_tGE���-i�W���Y �-���"��"b�9*����p�jh����p! ��f䯫���t����$"�+����hAڒ(�A�n0K���t���&uNH�����c����|�|��|�0���(pXt-
$�Amx�8,k��3�A&:I"W�Ձ�z�M�c�2�D?2G*F�b�1��,��j�;��N�Uw({b+��
��<z<�.�&�L����DB\��P���$P�	����K;�� 3o]��
ކ�gG�u���;�
�����Ƣ�n�+�z��#�e"?O��
�k��;��[�x�Uņl�����՞`^�~���Yg*�rc㪓��ÖdN�w�,��^�w��H�	�'��\W �^�.��:Ei6��'�����1�}ܜ�4�2����"�<&3��E6�FC�gfۜi�N�{��@Me�%';��BxP���X�Jҟ�?���n3q��2.�3�Rm���,�c�7D���O���@ьy�! �!%�ˑ5Y9+���%�ylm]�|'LW�B:�,VD���.�����2�h5߻#���s��^J�֋�`l��)!i�O��Z���A$��⤡���9�};rRsK��&�͢�kg�_��h'i+P��_N�H�g��~I*]m�Bys��cl$jV��!G�(�s:��ds1/oX����)�ڑ�?�8�7�[�&��X����}^�k�}v5Û2���f�	�z��E��1ȦŊ�Z\���H9)�?ӰMWŶ#
0�[(D��o�E�>^�T(>����1���-�%����W^
90�ǜ��@?�C�g�[k�!Q�{]��sD������U ,���m���i9Oڒ��?]ͮ@UG���R_9	��$xe�����c�NJOzw�7���U
�V�mM�N4]]ޮ�W|�++[i�5;�w&��$fފ�{�KϦ��c����3��
N��Э�B.�<�Wۊ\���og����:�l�B�b���X k�r�b�r}(G�:S,��d�R��.�C�uv����"�_��M;KzͳwU����%H��g���]7~Lw�aW�A�6��>eH�Ǳ;���w��%�4x�!��_4�Km�&7��Nx��u�@6��0\ȥ#
띌3��!u�'�(I�h8�KWB}�c�FMy��c��@A��K��W;��SBK�<~��<]9��� �Z�:��ŝ�OX�E�k�%:Ÿ��s�o ���x����6�cY`���~Z��R'��4���'H��N<صT��\B$J�@���;���Y�]�Je���`?�LKSٺ�����Q��6|H�#�:����"�f�7Ƴ��Lm#�{�)���`8�|̓'�bfu�]�on�/O���Կ#{Ջ�+��x�L��Gz���x�yɲōw�������-��Nw:�Q�Q����4[	Ċ���qBڵ��#�,Ȧ�kٱIYh��9;2+�{P?yp���'�򛌶f��m>[EȎ;��8������F�v`6��S��n$Ie��Nij~�,��}�HU�^'�3���y�}^�V��*�Fg�33Y����o�ܸO�Q�,b���W�NM���污�4k�F�*��:��$��z��	a Ĩ��W0N��86�s���LD�#��� ��P^�Os1�z�[�\��)8Mm�����-Z<h������ӡ&��0��`y˸��L����:��F�8:;���o2+�fK�r��*�G<����!7��8��*N�'���D��G�^�!4�b����&p�<��ZO=8�W[���.a갆e}��$�=�.k��/�\�X!Yr�>d�����hIέh�u��נ���.	�@��Q��	�������ަtbzh�`7A
loD�̵�i��+ٞ���զ�*O��Q	
�6j�6�U���O	�����Y0��ǒ���a�&�(v���5ҺCIo�q$���!���1�	%^kn8��7��*#���'�諕x��$�#y5����H�ކ��R����:�so�{N��H�_W�ܒ�K"¤n}*����8	B%� ��a����]�tZ	��(����r�4�)ynk�Ğ{�0�n�4u�B�=����4��).cY��=&��͉~*r|�Ͳ��RS/��iv�>���e�nh����<K�nҼ&��Ƹ6`&s��
7Q �έ�#�2�-˯��wD ON�e��7�Ҕ���u�ߜ=���Y��$�-���4d<����g�#c>��\��`�JM�||��`�9|B�)��?�aޤ/�A#��^j5
j��\
��d#��ʬ�0�������&�*�L��W���>�AS�x�C�&�\�f��A㳘��IGC���-��L��ʝ���}�V�r���gg�R���=p�U���+4�w��	j�ْaD?�9z�\VZ��m���$Tc��H�>+7�״��W˹Π�rEX�N^��`n�f�z&�,������A�w*�P���%�(7��I_��l�us
�rEZzV\�����W�2RR�����{L
���)��癱�=]ȗ�D��
A�d!r+02���S��_<�Zi�ܶ3��������6KeBi�DK���i;m���[�$��9:y-hC��O�=����~�L����,ĵm�|��tBp���X���ndV:�.��A{�"�K�B!���'�ہ�>�n��u(�>������6�W(�k&�D���"?v�ataE"�	� ���-���r���c
���D;}Z�X$���$ǥ2�1ӷs!Ņ�SʱR�c=�-[����6��1�U޿�P�X���x��|F2�È��pY����֞�N��Ԍc�`��S�á���9W�e����AV��n9��P�L=�3�s����K���j�Z,`]�U��U��T�:���2T�u�h(���7~��d�u��5��H���KqgNi����r{�^�VF�5������Ϩ����Ѳ�sG�
%�A�Uf�s��Y��XݹWn����H;E�@���RK�d�ۭ�y٠�fz!���U��ea掾�xA��A����_Z�f�W�ow1��\Q�k����.�5q�톄^?I����Ί�тg�;89�GRw)	�7;;E�6�Зě(�P��'��i��9c�	B�h�!=�������W^��wU���w"Fǎxj�ޅ���Z�]�.Y0����%�\��˞ݲ�Lh�.�;��<3�*ۨ=�?���>?�9ح�m��&e���A�3*bA_3#�^������(��!$���}�Ьg���j��ve:�2�j�`�ܦ!0d)3捑	@;��eC��Ƭ����SI�<5	{Z�t�ʤ�(}���ǜ��!"�����؆rO?��?�x]b��`��c������(S$��Ð*���rD�䁭S�
*o�z����GWAy�Wf��'X���
�tK�nL��|�g�V�s񥲭79�k�\�&sH�n��ir!�M�H[�� #�K��	�/*� ��Y��_��L�#ql���l��N�&���6�v?���.���W��Tj�d� JE?YѠ,L�}��=nd.����%=�7T��KQE��!��HB��q�W�ԀXq&�u�� ��9����-�8U�w��}u���B�����w'$m]&�1��	���Ъ��jq�:bV�W��̰x�����,	J�[ړ6��Xv�F�Ʒ��M�0�O����9ʋq��X+�g�H�)�>�^y�C� �3�*(]���ק'ު��*qQ8��k I���]	GG��|��29�e�sm}���<�'�}I�V$��]�-����'�c��1�Ǹ=I���I����HH��t�G��̕i@�ŷ�I������e�M�"lm�ٝ�T��r�������`�X��ڡv�q6��׻���O�$ "�����<�7)>n�a
�h�O(�C�w��Ǟw*#����)��V>a�ꬃ����񤐺�W��VmqXB�]���TΕ�Ķm5gt���]�츅z��r���}���]�*Ɋ��j?�،P��8��e��6��4��-���,��V�����Fج,
�j1�:��K�Ivo��=�<���}�b��`��#e(O�}��3�V|��E��s~rQ�։`�?��ev�$������S�t<2�j��� �ò��w�VEQ���j뗅W>�=���'7���E~������V��~
����V5jk|v��BΗ/�p�sA"��Gl�W.?lc*�͏�G7hWr���̞���퓁 `\uM\�/R�<�eq�.Ĺ�(�>GR#ҥ�6�h�����`���]\��U��R\&���u��S9����;�!�W8GP7$O�Q��Q�_@o�3ނ���8��~+�D��n�NB��F��M�Qfd"���)�&�1���9�b<�����:om#t�ԗǇ�I��f�s�H�^���;�O����+������$_X}Խ�e_	�*�x&��M�W��4{�ޠS@<|���^=Ӻph�O`��T�o[W$c�� 9o��lkyp�.U�9ƇqL�����4�6���j���2}vu+��=/T��?��pK�����3�c�V�\3d���=�_��������т��=���Sf4"�֔�f���ic���;�#�6�E���v����y�a��*ľ�.��
��B�n>�~�;Et�K�͹暀9ؓ?�g�x�s&
�'�N�I+��6�C��Q�H+-JF�����X������T�}���:<�b�ۃ�5�c��E�O� ��Խo�<9��~�/��C	tE����C٨\�?�^�1+��_&Y}��bB5�H;!��v�3����x�n�@�*�<���Atg��{P�d�9�4�N�{߱��,f�~�D���i��﬇����"�t�>�p򠀰��:�H��P'�0m��1��gW�C����m'����.*�2��m7IU��Jx�
V{�4DKj�7��\<� Hr��D���S�l_�7#X�,] ��e��]��6������;D?oH�]��*��SV�3r�� D� ~N�ZN�u���΍S�[��P��ֲ���آx����[?��(V�X��8�|�,�7 ����U!�ǵd��Q�O��$�^����Mx�(��H��C8��#�S�[2E�GX�0<�1{:S39|��woeϡ�z�r�"s��F�v�̀�p�q����������@����ً���|�4R�⾾{���|��l����0r�^����s_��5z��aJG=Y�\�XR&��E��]���n��<["质��+
��e�	�.V5��'���>���0��MX- �s�rB=��;/�k��oP?�Tǀ{�r���t�����;�LD[��Kz{��W)�b�b����B�{�S먴�B��qLb�X,�9�?��IG\�(�FҎO�9�@4���bBD)i2�0q?;�ob��6�	_��4X���ӵ����&��r�<yh��Y��A��bA��2QȽ��6��Ɖ
�ݯʱS�6��8�f�����sp���\v�n!81�L)��/��`��z��uL�gvc��R��ɵ����n},G������}����|��ql'��6�&����T8��tKqx]L`u�B��x47�݉c �����=E���`u{�h�M6_o�L�x�U{�ē��������*�L��8����ҿ�5c�[<#�	\�?�d6	2b�X�S�XĪ���=q\I^��>C ��Bcw���hj�P(��b��\�h�۽ E~���&� ��q/ F~Bt��Ė�]�H�u,w�y�?��U������>L��<��A6��ɧ�݂���vz=�l2�Ғ협 ^"�A�7���,} 
����<�Y�xD[G<����p$hv/��_�[:�����/��˟
�y��%`�}V�f��u�;r���&��ᠴv�6�w���S۲m�.[P�qԖF��Jk�N
�������3��#C�Lc�
R���
��`��y1�H��FZ�m26�.��䐟/�xF�G�cQ�k6�/���uE���e%�h�_�N��q�����1"��En0bÅ?�}W\A;���8���դ�L	,��6���l#W���sstÈE"��`O�-��F���\R�	c��޷�;2���������g=\�/��[n�5�Wű8Ik��bFL����~�W������5���D%����Ȼ����ra�O�x�TY��*=xt�b��vE���6\���wL�ܮ��䆬U�i��6.�9�:�o�B��4S7���Sٛ�v؊!^]��qƣm�l_���)~������J����Lͣ�0P�5e"����?{.>v�_IU��?!P�cZ��/gm�76U %�u� ���Ds�����Bc�[`a�+)2m�Ph�� a`�wo�\�,�WM�01k��Ƚ�q�1�}��>ͩ��X*ijBS4����ΨM��A�[P�����h2���-��" �q�$����8�OۉR�'�����"�.��z�,�ܵM�`8l�򔭨t�(���%��$�#�.M�g���#�EP����`r������SyS��-q���t�V��Țp8ڻ[I�QNu���!&S�N��wl��lLrgI������j1��:"���!rVx�+��2c��l��j*D�-�x]���ua�YA�Í��xI��D[��d��Dz�r��ޔ����h�~��	x|�6���{=7����R��/xc����Iݠ+=B����"��t�ͨnXڪ<�@��Ί�I�:�(1$W���O ze5fM���x,�T8m�����8�A2� ��>^;�e�`8y�a��b�7���w�"������dԒو���7�DT������$T��7wU����<A��ʨ-H�G�{�EP'�iW5گ��f���0�G�F�C�t~=��Kze<�L]��=����KT��ծޗ6��Jy�4;�7vg����9�V��Tާ9��"�~ԣ,辬��E���i�ju���2D�ߊL���2!�7Us�Tlȋk�:#�f�3�F��]�^M@�O���̱[�D��-���;�B;y!�#�YO�(O4q]�(��j���M]�i%�����SpQS�V�<{DN��g�x��L_@8��F�aǇ9X"��;�����s��.��@����TA^�����,"Z��o��]m�P�]�{��"*Q}=͸p�unp�LS���7a1g2�~��y³&�-Ɉ��`�"Ёy
Hj"i��+���J.�|�h���E�O�;����X6��̴}uBHUG�S�oՍ�ۭ�P��N,#˺��d�`�z.�X�'y%7Mb��@HP�[+%^c��ۇ�[����P���F5��34��y���z�IN,�VpWT�T����B*��4�b/���J.�1��8�N�Ze0��,�WSm%e���4�L5�Z�����}�񌜱�ȩ_Ow��M7dHl)�Y]�#9��� �D8�4#2�:��nP�������S��0$/�����S�R��𷐞k��1�g�5`���xT�h��1����ͨS{!�����<w�\�%Z������{��o�e��42��}�����5�,YgV�=�k�νp����������~ �TW��ϋ3ԭ3���~�G���4{$Q����}�\V�~���4���،(Jw�)�{��Ih��H("B.��P!K���_EJ��c�������f�e�]�.�&��Ia!ڮ �:���@�ʳﳏ���1us���y*��u�uf��5Ul��B6`x'�+��Y��}���D��n���4-ذ�m��L	H�0�����F��[��i�_���۪ݳP	Q�qڡXǣ��(�s�uѠ4i��M�a���TB���
��m���s���%F2M!������c�Xa���A_e�zE1��
��+=�O��ٖH��댡j=w��xbbPˏO�h�LlԚ
?\�uwC:�4�s���	���u$�k�ߗA���҃k�'ɫ|�d˹��v��BS4E�[�ħ��S��ku
�'�ʅ�К؅��;��**{�G�������Lk[�E����'A x��|���E�0�/�v���.u2�^\�ܱҰ����݇��d�GZX�ƴ"���@W�Vv�^��)1����ZqiviF6��P5��5B@E��<��&8R��ߩ�ȍuR>�*2�L�{�V�"�1��޴�
b���}�XNG�	���czƘ�֋����k�k�r(�u���h ��݆�C5���PS�_�8/�0�nLfd'dKݟ��y�F_b0\���曃{՜1x��5�@�o>��m6�{�#v�>׵��^̟E����v�z����-�J�p��#ƫ�(.��}{q�Ǵ�Q�V������9�f�~#j|8�ք`s$U����o�RC��G��k���i���}�vv��5�H@%Q�)V~@;Z�����؝A��f��ΆV�à[��^�!��1\5n�=|��:�6o�C�PG��b�1�.���|�v�)L� X�PΤ�0 �����m��<z�W+�:"O�+.�U� n�ġ�	{S��nރ�&C�`�׽Ï�!�埅Fq��o�4Nj�c��&�G4�A.���9r�ꠀ~�sIc��d�����R�j�L�c�0̼ ���L���#�;��iI�5m�����nȑ��!�هi|�]���W@"O����8ˀ��EW���v��B�� �K|�l6��M%$����)�ՐG����3�i^tn�A��z!�	�����M�k�*�QŦ�(s����"uC4��ݖo���|�~�X����(�-��d�`�-¸-���8��T��rv�:Q���T��~|iI��=��M�)����/���)Hˮ��#���06�#K��"�۵��J���{㢨|'��Ǆױ#IY�^K��j��X$w�H���8�'O:��ǆEiaG�� }
��ms�Zf�;�^^��C,v"��$����`?Sb��-@�ҴB�FJ�(!ҙ쨒4y.�e��$�;�e:)rvqSQ�w���^�����G��~6<�Fd����7�5��+6�+F���D}c̀RK��`�D:V����Ft�7��}�
�q��[��ٻF8�2F���s�`),�aC|e�vN(��F�L�s�V5=�R*Yq��Kc�vpO�ʎzʱ�aW��c��AO�n�厑6;zp"XOYO#b��;+�e�	  Y~<���ˎኟ�ˇ���ԥ`�9�)�nٶ�~�;�4�������*)�J:;�C2�I�/�ߖ� �d�6�B���������w�zL�o�~�L�_f߷a��P�dp�Az.*��^�ҀM���ϜL������Ӕ�#��!����ҵ��;ZV�S@T��S�@:�iwh����jDm��K��c/�I��L$���ӟ���&������Y��oy�;ԑ*��>��9 ��d[>��i�}x� 
�:�5{O7֋��.0�F^�z�Y�Ry���U	�X�����AB�8W��+��M������31g*Cz0q�C� NZB�K����8��{�K�BO��KLX0M]������YU�6/���*�[X�r�pc؄-�v�oK�S�1UF��Ի��!�I�n�;�Q�<��Џ��i<s����1@93�w�(Krο3�J$l1<�b�I���R�E��w�T�m���PdڬV���^��y�֞�Q/�P��c/k��y��8������h?�C����ҭ�clZ6���ŐR66��5���#����@��V$�E�<(�G�0ҡ���]M���u#A���xPzTˡU��S�ٚ��<���]���6�0�4�<O��+�s��{3�q�<� :3�Q{]����������&`6�p�ӫ��@��Q(����iJ���7Wh�*�ld}� D�I��ێ!�y�u�$em���h�����������&5 E@BZ��2Z��u�Ab��_/&��,����A�V�-Z'�M����{��b��+��Fw���L�tA��_�:�s�JB�C���W�i�& f�C����4������/)`��&~��ڋ�^� �`��gE�X��"@��*���[9�r>(f�,�GKT叵�>+7��b,�`{�����ߕ���#ݗ�N��En��FՊT����wHL�� ɵ]lL7ǌ����"���l�_g�S��b"���M4�"g��a�1���2K(���'?��ډ�.>�b���t�,4�|�t���w�y�_G���p~
P�m�?���1��B���<>4�Ҳ��Bxn�� Z��;��"��4�����|N����@l����z%Gx�2���u1�	���٤d]�v���#��5��SN��O@-.�7���\qUX]v�v��0�����0��Y�P��2΃� j�A��f�b2Q�4����A"��:����j�Vv��d��6�F�z��{l���`��A% au&�gؖd��i�,�RF��W��ep�\6}��N�n�zET��2�ρ�>��xy��8���yOrs��~A�MPz��c�΂R-�8��o��XaS6�����̞�� ޥW��YLNCLC�5O0�m�3ڍ?�W��R\��8���7
+���i@�I�W��&L�_��p_�����rM<�٭�݃V������ ���L�а�:���:4+ݙ�!�*y�x}裓\s��N�S#o;bD�Q�~�_���bLD�"7�v�:��w,1?Ýe�w�Çc� }<o�f9���,{��v{/��@��ӊM3f�����O�K�#C��!{4,��.�)�Z}�=D�Y�ƥ2��H��TM#���f��Vs\�D�F�	o����4h��;DWĄT�M`R�� �����4q�P M�X��2ji�}�K1���ݘ �LU�^���m�j7�|E��̅BaD��h/(�bײL���?Ă1������yԧ��H�
3�Η̈�rT�K���@��$ၹ��8�}����ݔ���9%�rd �&.��;��+�T��N�&�`�9S�X�滴|[ê_��{ЈyB-�q�����A���%��ֈ?�H:�H(��E�U�lK�����f~�2��N���`j��=��	��_J�E/����6�o�%p2�k*ySr��Ll��݃�Q7��H�#��|�0�jc�AT�#�S$���^Ji-��vw�G�GH�d�T<�<*�X~Y�- �HԺla�X��x�ʹӘ3Ԇ���3s�x����£�j���=^��՝A�P��("2��F�5���
C���S���4s�+���g�"�(Ä�3Q��Ne!C���DO��4.���Q������ҽ�����g�:��!��]�=�N����B*�_�2H��V�i�_	-q��{�������l,��.!�n�5:iz豘�yR���DU!����T�4����E���E��D-{�a\���&����s3��]�y�>y֝��6
j�RN�Lu�Ϗ���>1A�2��@�b����/�b��h��7��N��ّ^`�uKj�9�J�a.�pI�xqh��_��)����Ց<��,BF�U+-i?p�?w���2v�������K��KM���7p��X(O��Kb.�����.�����W3���λ!��CQ~��_CD67-VI��-��Bn@�U�fM)�7XO�ZB�L�����DI٨�k0��l�29hĄ �d}?��������{N�7/�u�.��2S���/�e���}����.��"����GMaD��e_�Tw@&��?�3Lh��jl�qL7nu�"�)���Ȇm"6F�X�╓J:��Q�l��AE�^�KSb
�2e�[rb$��Q�I��`٩>����_�Q
���FW�<$�u{ۋ7"��'�k��I�"
	z/���S��-��dr�]g�+=3%N}�&����Һg���NW�ż�N_!�L�q�q6�S��Hy���ń.��`�*�Y�����f��qiWÂ��a<�8�
��B^��F�O�~h2��B�l�+U��9:x'�$�$+[�Id$�p�[bS����#����寞�0��{[4t[���I���i�$��c��
�����~bYCp`�_��ׯ��LDs���'����8��0�Z��?K�̩:9k��-3vPj�*+�AN�Б��� ��+�'���X΂��M���T�8?O�W(�ő���B��S���W1fjj���'<i��f�~@�î�**�����3�a�!K�n��^l��5�̓�?Ms��8��|��zs6�I��b0�>��[�O��5y���j�GEy횝&Z�6��֚v(μ�w͍�Xz�fM&��ȿY�� ƪ��͜�C��e����e�3���>bH��ª���KÞ��T��"|���H!ͩ�J��T:��b��s�
S6���Ez q���-j_Z��L�d;X���%�u��?s[ML�X��I�5܉U͂?����<�7W��&�' ����}c%��JH5���z��Ӡ�&�*u*��pP�q�8ǹSq��ˌ��c�ZgƁH�ĜF���ɫ��^�3��5��� 8gKުL��МC���<��������R�+�,5u�W�p*
%N�Ͳ�,'��� )Ow\��x�JHp���B�m
Y<1^���>֔�Rd�%���W�%�Ct�}����tk�H��.ݼ�S�����8G"��������L��.��@]�����n�y�9�s�7-ٛ2r[��E�����$Y�M��<Z.�#����L<yV�ÔFQ�Tb6_�> ��e��+/��O�E����hF��U���%��&˵�Ϊ�jb�2pUh�W��f3���¯�?u�"��T<Fp��k���.`)�g�~�Z#��s�?3㘴י� �e��u�������<C�:���L)�s �ý��q���$*$���,���>����7ߩ�Ϩ�iF�F�ͧ�:�<Gʏ(�cIt���߿���D���W<����E|�w"�^<����DTWo���*/i�р)�d�gƊ4�ߤ����!��)&͒��?�F��@sbm=cgӛ�j�ڳ~�%����~��)�� 7��8O�e��}�&��<%zP�ٙ�f�R@.Aw�̹��j
96�ƭc��$����VBO�2���(��dF���k�+[���5��㍦o����	�h���qW��8���'�`{k�3%�}�0"@���������rl��'�[��
[��J�������B+�gU�ҭ�ܙ�2:yS@d��ݳX��E�NI�����{���$!ƞG���9��g�V�ir,�?Ϯ�ŁK�ᩆ_�e"M�*�}�ɗ�O�����ro ����b��jH�Q� v� �-l�<c`�q
}���=
�<�;G�ܩ�8�g\?L��Ÿ�������TU��s*�ߴ��T�ܭi���}�e���r�s�$���*�k��7��)c�bE_X������1��i�ܥ���Cm��,�r�R�@@�M�c=�t1T�G~����G��kc�55Ҭ��b^��w�<�Čt��!���(�-�\t7
�M8����t���H�ʮ6�_H������d���d/)Ng�S���=*T#l0Zi�e@/-��-}E��$*E�$�1|W��u�'��ޕZ��N��='7�tv�ďe`Z/��k�x�og�w��=���=�?Qj�fT���Kt�O�u��c��`
��ּX���I�0���qa�M��#�����?Ng��b�*&t�#�K�Pd�R��l��FX�-lV��b�H��1��L�jū��#���4��r�=M�Lȝ?��.}�X��|��Y��<b�W��@=PV�������F�E|׺Yc��6#��Tg--�d�5[>�>����kD����\�%ڿ�D�6�WЁ�x���o�{n��O7
>YÀv��O�O}?��GَMB����]��u�AT5'��Wr��8	�a��ns��'�BR�]~ҥ`�-L;.Z�}%�Y����=�m�G�6P@�&���j _sMy�����M�ns�+�0 ��4"���X��������Bqꯕ�S�s�\�	��F�#�z��q6�Y��Ym��`��#r���`�>�`K�0�x�����x�t��u�F��/}e}����D� �7���+�	Q{�6��-<����P�l[sI�D�y��cv�vp�Q�
_��)!YwiEG�"��~S��/gGM��@���ZB�St9ς!��'�٥b6�h��߳�'��G�oġn�|���[k�2u����E�2홭w�N�Y��ȼ�qKH�ţ1f��hD"���p&$e.,�̏r/�3U���VW�-�~O�C����I�f��~�١MK��e�3s-'9�K)K���z�X4���A��GUˁȔ$�bMO�^��'�\���Lv{E�l�EZ��|�o��� :ps�sTr(S�c����M-����/�o=��G�x��(%�V6ra�p��.C�ci�q��d�^L��{R='{�F��8�a]�(�Eb'q�I���5��I:r���W��B6��y��Z嶱���2�J8���KG4�*&����(�o�Q�x=�ʭ��4����cp:�~�e��]���j@4���q������#Kc?�����Q��J�!,fb��G�]�=8�XΩ���M��k����8�E���s*bA��f�@΅ �pX�(=r�c 婾S��ql����E:@�%�4��j�l��:��@%hdc�[^�5	o��,��Ƙ���ݷ�w�����e1��d�jy�ׄ̈́[����D)�N��(���u�h���Y�?�����oT��6��^d���^�$PVꞄ���tPŞ��=$��	���VGAJv��pK<��������K�0P��bN��b�˗�1w���t���F����rLlRf{��pĄ.|�[5��C�Rw���������1Y�k���h:=	�B(���%M/��T��e@Ϭ7� �x�OE -���,�knz_�5�vGt�,X���q3hqs/�uCa�`�f��0�&P1��>���ڑUBr
����˯��3J��'���/�+x[a�FY7_^�a�Y���Xްk2"l��4��z��Mia���z�y��!r�Jsda�����hvn�]�6p�N����9U�9��A���'r.a�R��	�4ۓ\c�!�� 9��<��!�ʳ3���2 �IF �Ri�\uJ��s�o*1��;�K]�z�G��򨰇�I6��D�������A8��Xcc���,���w�2��j&ٳ��:�l��x� R�����ו��V����x��䍦f�+K@�G��3��j�`�f�"b��x��E4I8��H�o�[=#M8�X �����S!��)�Q�8S�8�s5�<�o��n0�ɽ�k�)O��F���YO�qQ�0V�J%	�s�JD���"G��6�u�������!��El3dm��v���C�S�u�Bύ �;��/U"�x����sҀ�ͯ�``�W������p��Px��m��{b>��t���[�^�bv6��C�M�.��k��
��W�M�t�Ƅ2���t�S���E��
�?�}���n~2;�^�'���`�F]�4z�7�&g��K$�h��'ѩP�)9V^T箲�vA�b�E;��Ô�8����ۿ-����"����@�9S���}��Y�������q?�!oO[Sg+:�E�a��@��8	���]���J�E���ƀҦ�/���/��]M�z��D�	JG���(6�/_��]�Z�_6�G��az��g�O����FL�1�\/��'�R�ܸo5�S��%o��[�p�x�������)�[�t����0�oM�N]�2�Y�|l�6*WC̍T���|���6��k���R2�	�G���	lA�{"�3�Vz�mz��F9�J)sͩ���B�5ZdFY�����ᶗ�ҸZ�)���ba&[#���_k��������S�Y��{��p�Y��"���I�_j�~��y����ȥ¨iQ�R�� ���y�y���Z��=�.��H%R����=v	�rhe��.�sX�)-���ɯ�4[�����~��_ۛ;ں�=���g4��8�e=Sr���L!�Dӧhl^����J�B� ��zّ���}IQ#�(���f*H]��4���=��=����s����3�t��V�3!q������3�i��k�b�t�[!.�+������,FV~��3Yp��ܒ`�0H�ˣs� %�W�[Y�E�J��a�{}������=12sT�P%�Osx���G�X^�
�P�;�D����Ĭ0Ҭ���M��B0D	n6���{'��A���R
Sm{I����*��?-�2PC=���̒c�Y�@D�:=rO��<�so��w��y�D+ð|�	T�J�����T%r.��t-ۋR��C�Л<a�|NLC�ue�%k��s`�H�����M�/���i��E1u�&����ɋ+��nu�(�z�^��#��5�pfƹ��5.��!}>�ꜵ5�*B��_�.��hL�;�7������Y;^R�V�!�Fg(LnIK!i�n@#�v!1�͖~�Ք	�>G3#"��R%`y�%&r}5�{���
���^ �+�M��b�[�n�2�1W@W��2��uV�l�l�R��m	j�ݒ�\�_��2xr�\1�X�K�W�f����ОN9@43|.�}|̨) J��.T�˜���)?����+�-���3M�鬴J�����О��0^��q��?�.[�_�+]�Ȳ��Q�/"��)�I�62���CW3Z��ڍ��$Zw��W_if��a�4.k�6�d��Ӳ��,�NZx�6Ş���>+>�7�Dm;Wn&)I~�KSi�� �V��=Ï��;��l�����ߞq�O�4���a�KI�ba"�<M����k~�lp(Ƴ0_�hgkI�pB��*�~���}Ts�Q#R�����e���������d�2�(�e!9�����1�$faHRl�փ{�^u�bbM���#EHV*�N�5 lYڭ!(�@��֟ܺӃ`>����0}3�o����x3��([����i���F:�?�eC��f]Ee�֛^"���o����G�a}R�*��zJ,(��-��Z�M �I�Ǎq� ���N�a�@�f��W���&�3NǺ�2c"=��F�S�#� *B���Ο����@�^׿h�>%� �[�?��Q.����)H��|����\i�$Ŕ���_�=��2�P�i�\I�d�S`-�C��"��� )���S����,wϒ��]�,@�VL����<'θO|�ﯫ*x���E�A�_�F�57�ϥ���E�-��+�MSaS�p���Ytl>�X@+��tR�*0�p��] �H��_���n�gO�c(�UB��1�7�3�EKaD�G��:G�=��@(�C��������\�L'	����%�H<1�~r���2�S���n{A+}�XoI],*2Zx|�A�A���~@�4���\t̚ ����'!?F�ŋ���*f�_���W�40Ԩl��بj�N��$c��FT;�a�H�Ӄ���������Yy^�+a��+?)�z�)Ŵv�"���>����6@�Iu�����
���>��.�2�(��-�p�)O��
K��2��,4� A!T�>ZӲ����	���Nfuuf��k�I<J�%J{����5����#������4В8��y�F�<����W+*����W/��V���f�3�i��u�cQ�&��ǧ��T�a��D��u;*�Cg�-U/r@,�?�ŉ@f�*��u�9_#�h4��+ a/w�_D3����6���Y�ʜiÑ6��aM�+����5-�"K��ٔ�V���y�fa*M�\����|�rs�Z�摿���Ж�#��G����LG�[8�$l�Mk7I�9c��A�U��a�/舁�_���p�7r�T��6;�q/}�G��J#��B��Q'�T^zf�Sk���F��h ��ޢR[���C�����Zi�b�EJ��"�mɽ��������J �i�?u�FX������!l�O��0��/�:��R�;dL�-����(ѱ��w����j\�I#�J9��F��bא_Ｘ��X��%�����Oi���࠾:Zͦ%���R�b�
(ی$��4S�6���VC�e�Gb��%ꤽBQR���	�Z�9�
��(��#��k5[p���e�)�AȜ,���ROz|�T�̓��'?�A��lҟlΙ��HQ��gm<�/�m��ڂ�"��ى�Q~�Y��9���K�D��G�|8����3<�91R�ux���A1N��}���[r���/�HS7E���_��Pj�7��X>y$������y\
#��	��C��[����wZ��{^��k�%��n$0�C]-�N)�NHH~�$:)�[ 9�BbS���sL�\d/�]da�T$(�X����l�w�<��^��؈��+�����CK�3� ��Ò�q;���b`Z*�r��e�� �sb{��i�C�3ō��_��PU�h7���6v΀
U�\��˅�!�	N_����r�]��G�6�-�_��lz�$ya6�Kۿ�i��C��z0��LD���A����_p�K�om�36m�������9Z�C�d�[�G8 �aF�+j<��C�X?̖u��W�	�=��a%TM���e�ݑ���8CV72%>s!-���h*��1�~e���U"��1˒�v}7g"���e��t3�Z^X��<��5�(̼���{�jf��,�J�Ȅi%a�]ac��?��Y�������*X"xyH���]V�$	XK�iN�,GC�Z��'ϱ�Tpt�[ꕢ�W��hk���8�1����v`�@�Ah	�6��T�p`�0$J����vK�yU�-Bb@��@_��[�|���w��n�6����<�@ۏ����=�N���;&D�l@�������Fy�;H�0�����NE���*zjCE9G�<��Zd�߽�Zcۑ���$HZ4�^��a� ��SS�6��,0pl�'��K�)��e��(��;C���j�+\�!��]܂;��Uj�B8� �lG�S cN�3�;�=ۦ9��DL��T9�`�������(
Y�J6T��V�k�n�$�Q�a�� ���ir`ݸ�>��ɦ�����c0���d��`����+���-�
}�cW��0�O6�Eʬ���X�)��ޙ�}9���u��5�)�D"5�v�Kt��eVx8��ɴ�*�c���|H�kJ�M�S����N���	fG�/@zTD�Yժ��{'A�׆�K�B��R�;fQ�ϛT���\f���λ{��������X�bKGg�U�Ҳ�_��	���]3��	,��	��"��9n�����|�?�B[�Z���5�*��ԛ��O�[)��1:�XsR��Z��bB�p���RE�Dţ�����oil�\-��\]�	����f���«l�R��Vi�'����m�3x�۹sۤ>rc�E�6p��{���Jg���dG־�D�!M+�A�*����˸ML<��ޣ7 ��h�ձ+�P���b'����$������kc9X/�J�·��BYZ�5J��H2N�^Ǯ���A\�'���D����8Q�xn�y�$\l�l�+x5t]Q�^��|�7̿��U���`B�{�!I4h�5�H�i�1T@�=�Z{���~#�b��F�E���g	>���ThXLQk=��3��FV>�����C�/��k���eL�c.S��%H|>�e�4m�(���� D�Et�ې��C�����W���c���Yߊ,��x��_�Z띪�	h�SE*�
���7#H�ݲ�,0�71�T*6�x2�)\�b�s�ܮ��쟁k�Io���K_YYp�D�+0@�2T���ba`.�4�7����gDA��c���yߪ��3��^H��6�6Q����A"�Z]�ͳ���&�=�j���>_���a��t������"�]R)�fI�A�1��k�
=�`��!�H����![�_�K������_ov��q��&f�Ky��-��F0U,Tz;���]�����u�[r ;�C����0�M��T[l�[�7�&����x���n���P��b����gs�)��*�X�C�#e���^���~��o�N�E�îX��n\/���K�Ė�<�qڝ��\��0���]A�Eo���]3�%|P�é�
��C�/T�1Ɗ{�1�5�2�eo0�=,LL6��/a@x|��F��㦵�^��yuK�������A�f%Ǐ=B�Zf��7���3��򝵘Q^>K:Y�F�S��wl��	C�B�
�q�@�(��	��m��FZ�Y9��+Y�G`+�H���4P,sk�V�o��	Sw������b3���)�~���󶹪���U��ƲW@o��+n�F
�̳�l��l�\0��#8�}3����:���ĭ�����������J�}ǲ���#�Y�n����}�����<e�d���ʛ孈1�H�Lu�8\��`�(��&�
ϝ������Ut��n�H�]\�ǝ�����)�C�C�^x����f�^R��<���������:��˦��)<�(�H�݊=C��)0$�����u_��aR�#��~�!��A�Q�yjG�U�j��]a��t�@�f�,�hQ8��{k��.}��{i��𓅂����p�� 7�ӓ�V�s��]u�Un�}'�]~���s�(�׏����%�w�/�
��0,�>��t\�=[X=}\ ����ī�YK^�Dc��'��ŕ&��p,�p�P�$�S��Tu�F�H���"dg��,> .�����ð*�i;p3$�>�)g��2|� Y�8�O/V�A}�� �7�`�I�i��$��J�!o�{θv��
ے�=Ns�h��hV��<}]�����rTY��%�����Q�B�6H#>/Ntn	��m��}l\L�0���a�kN��H
�����dc��U�?���i�sK��8bVZ�g��v��	�p炰20S���!�èI2�mS�	I����!2�Y-E�i�Ya����|�H��d��9.�R��Q}{4.��^�uK�tGa�&g�A���\#�O�^�{)(
)�fҪS�ʒk���b߶����A��E{XC������������*��������)�d,��E���t���<�&> ?+TՀpcE/=�È2ĸ7�B�"�����^����8�v�K�-:��-���d��ci?9��G���`�:C{Ec�ս�P߲�����C�*��B�g;sϔ|2�^ާ��k��-롥1�]VЬ��
��ԃ�N�0����T�]��e4�Q*EAz�d'���iQq�镜!��W
�
B|LG�NC� ����X���7A�S�!��� �^�j7���������5�L7e<�hmO4I�5�	g�	���Ѿ��*�|�Ri������\�Fͩ2ϓml
'Qn���Ϛ�;��g�`߂H;������hŹ�3°��Ze��fԃ�$(�����N���&.��H
܀h�=s�������L�������Zn�V��t�'�A�|�j� j�4�X����})N�f�}YM9��<�a3��j�}�̒��._�^b6�/����J�l���v��z@g�.�BZ����*T!������!(�L�G��`L�(L�+��(��p��&�X�����a�����`���ڞX-��z)����q�Y���E�r�~	ķӨlW���ˣ�S���
���WF�A��oF�0tS$���v���ͧ,v�MѢ���l���τc��hT�*r�$�b�Cq�2.�e��	"\q-Za+aRXHݙ� ��j$�y��3:��C���Y��b������.fpO٥"�ԍN9_x_,%+���d��!��~S��.�������������;^ߝ�Ф�X[���W������>>ԕ�~�F��j��'��5��_&���CP���iիz�94�3�����:C�2Z�2�D���4C�c�WaHSo
"6(�l\$\�hprC9�Y*�������Ox=Bx��y/���$��a����!�t��3����L����h���	7��f5���������ú8�k�-�O�K�h\c��%�CU��J	�&��Fo��K��O� ������@3����?O��I^���-�|%Ē�6ug�8�� ϩM#�Y�}�m>�l}�i�dСM���l/�O��J.ūC;�s��1��ct@0�JC>�
X���F#_�A��,)
�Lxi�e���������v<kZJݱ}������X����?b�!DZS�o�F�S�]��+61fQ�Ǘ'�������G�F"�%C�pi��f}.*����C~?��'k~(�R`i�ț�T��tP�ٖ��r�,��1�K`��c�]�Y�$*�#zHDУ-����@[5��˥�(�$���&~���~��|;2@2B��`��u������d1E�^�L�x���t5��i�?z�^r��[��|�:=t8�])tL��b�� b��>�%�Ӻ�D"oN9Dv�O;c�g�W���+���4�u�@#w���P�����B�>���W19�)��� ا��h��=�X�D�o-`e�<�c�8�b"�[D������]��%��N!��iF j�"f�Ex�8�_���q+ر��DX�|�A��k���cU^�;��[F��;48�'�Lv�?V# ��ˍq_0�&̀��{�H�f>.��˖j�����|Y��*A"8��K�@*َ��B&�|,�;�RP���񑧲�����L|'�T��%6��8��*Z�ͅH;��&m>�Հ ׬��u���ܽ��,���<�6J�+
n�ܛ!J+)a��B^,��%�Ʈz)inIÒ#� 8c�*���yq$�7���$�M�H���祈�T�\����+��b����3��%�,Y�}#��?�)����X���}r<�*� ��KT��F,�*x�U �8\I����/��F��d�c�d!�µr�C�5U~�\(��T�p;���b`����2���֪�:Dc�
�q+z�l�F� w��I��e0����5���y!ֿ͈�͌���V�k{��KKj�[�?[u��
��H�b0��*]?~�4����'��@ZM��Ֆ�E���Ę˽�߃3(�!����hF�՝�0�g�N3~9�I�_z2�@�1.��h�+��� ���͵,"�H�@,��ီ����h9GD�P�خ_"���~Lp�O�`o��2����\[���D��Cu�xgE�RІ>B��y�:*X�4��|�cp�ő>���a�9�j29Kɽ��m�d�7�)Hva�>��x.����r�3��>�XЖ�R����!Xq?����L�%G�+�5�[R�4]!'|�d�bW
���;#��ژ|9�0�:�.�+�Ֆ�@�<�ܩo$�(AL��?�i]Z�U@X3��m*惌���۲���
讬� ����~�IZ��`Ƶ�C�����GO�sv�̩
��mxe뎷~=0j>���w�
s��|1�[M��;�/�x��z=�(���$��a�.ߐ2���i )���ݢ*N�yځ�׆]�����-'�eSC O��h4ẕk�����CV}:7�":�`(e.�Z6b.M�$J(�B�7����[o2�<M��x[Yj}��Z1��BD��~���)0��'nq�4���W+oQ?�+O���-�[�s���)W��,	*��J�"�|��z V���h(�P��K~�����pg�O��<�H�����tܫ^�֦J�|-l`���&��9�^S��d<�'�;{@]�#̺P�7+cK��r(��e�+��y�Dk�,~����uӂ�Bk/�0j���M.�,�\�H�V�p_j&W�<���s���|��md�k]�ɭ���-��f7u���h5��2���IU˽r�3�����]O�F*'�Ǯ4Z��f0�����C�E�&� �,+Cp儤�����,��S#�������W�J����B��3���� V�	 :���E;tvl�I/�p;Yt��r �MR:=iI�M嚚�k��Z���`��B���@�2��^��c�Ft��<����:@��F�4M�m�H2��f��
��¸�[f���H�׬q|i�ŪD1�#���
�!gA�N��C#o��/���a%�8 J[Q9y8�<٩|�?�+����\�(8����
�L�v�~f��D�����	 Z���[� �������=h,�Dj��fC
+��g���?�ڌ��48�eGNgѽ�KU6_}�:#R���l����g�=�=u�h0��lA���� �Ϙ���@�ɒ�$��N���Oq/|������P���b��ڵ�c�at�1_njKfG�LO��p]�I��,�	�?+��wx�72#��oB��e݁Z ��ݵ�
�Vv[��:�˷�e���ׁ�.��� ��j�HM��:�N+�pX�[�_�Z�G`ѭ��v|����;?�]�e���,#���`�'-�?;��;�Л���)%�<ȶѼ9r��=�D:�||�ޕ���X��u�r���#���0ϒ��5��pA��+R�L�q�����ŏ����X�b}��+Ǳ�܅���� {�L�.N\�8ɷsU�?���;�^Ů�P�'	LW�!h܉D�*v�Hҫ�l�t-ɹ�����j����Z�'��޺zA�KP����4���i�U��&��L��.�+u��S�:ŝ��b���az�R���V�hw��8FX5!����f��NJ,�
��4+��]���kGN��&*�R��S����L'������. jF w�ڇ�p�2�{�\�ٗ�~�~,;f��IB�5Y�Ӹ��?�%x�.)�w*��&��{��ĕ�s�t2n�z3-4H ��1�zu�ά���L��7 l6*�cYf�y��~o7!� Bu��y��U��N�)�
�V�ÐP'�`Q��w,v
��=KwET���U�3l�4K��,m��YXwY5g"�l���1�V���4i�.3���h���7�o�����i�	�*�U�N����Y
^���}��m{�/����P��ES�\.p'���Z9=��y�4���
r��i��|L؜ǔ,}��Գ�=sݼeJ������3�OY�rB@�#��%�JR��;�,�q5uP�8:e.[p�fR�HM/������ί6���d�k��k��h�v�/8vb����˝��ǀ���#ec鑓Z��΢���%E�1я*u[�5V�	�Fq�������U���%���%@��lQ�Y�$�q�r ��Z��g7XS���nI����	2��ʰn�M���.���Tu�#���C�EoQ\���x�[�!{�i�*���Z��Γ�y�K,�Ҁ6�W�4�s��S����D������+����,.��}��46�Ts�zA��y��hԬIO�@(�9s��&�lU0�80MU�+�^<l������~8[TA��$%Z�f^���BD2�np`p<-SDE��YR�ո�*AnbM�l�L7?5�l�J�S�2���r˺��!'z���Ч6��d�!�M�������z����u�F( �2;�Uܭv}5���J�q���+�r^M���!گJs�y�X�AS���J�@��1g�p����!n[3ƞ�_��*j����Λ`�����x�A���aP���m�����$n�{i"���M�o�� [6��$J�ҁW�ߧ�����N���ȗ5w�Am��&dP����D�q��)�k2�{��F|6�SSrJ�����T���^ƴ�iE>��ή4�v�R��ڎ�����+y����t�_�;�����;���o��?DC�W�	|�0;�VCU���p�-���a �����?Fnv]�m.cd��pK!�)t�0Z�G#���jό���b
�p2�.�ԣes!k�b`_�H�Q��x��Z@6���y&�l��d��9��'*4,4�8���3G}���q>w'�?�i�.�K>j�6Ep)f�K��jg�-�R7��"[�f�]ǇN�f�D����:[�u1�}^�������]?s�^o��}c�l���D�i���
�4ۊufN��>:EV��Y �b��S��a
�~�e�����\5�Z�9 � �DZ>`�Km
.j��t�NȾ��[��36Sj[��
 ���〆#J
�$�'G-�Û���j��M�!f��������k{d��
���D,�!�f`UT�zXđ^vXS����LJ�V��y(_�JO[�s��R�s%�q3"'�Q�Rhc���S}��/��Z����q��(*��ۨn*�`ީhva_����U��E��<��X�~�ډ8��)&S��|�5WB �V��uu�K ��\�I�'�������躀�"Iڹ*D��f����9�H"/���$e����������)V���$벞~�2�
Z�'\l�#\d�:�A	��c�殩��xP�^��K5/,�,�OP�Ӯ�#�� �X�zPũ�*X�t�`��צ�	��OR?�LV�֝����1u�'��o�w�(�C�O��4����la�Jo�ă����ATD��<���f��^,�
��X�j��";p�5�����HRb��[dkt2J� t�IK�I|�A@e�`#?#]?�2h�-�\��^�$���WRMy�Cf�IU5׼��;bk��n�q�&���N��u��7�7�m��ϻ'���*�v?|�T!��q����w0���1v:��ٜ��Nzl!�6��X�?�>}]�v�Y��`%E�K|w}�m���č�?w�<������ �R;��pE�0FU��l\��T֡(�ʳ䷡L�"(��B���8'1�.�����V`�˝��]�&-�1�834^�R���b�I���N�F� v����5�"�4t�[/���M����JZ�G�{4-��8A��㍀-������H�Z��6�ĭƲ�7���BYH�婶���N+?��;������zd�yO�^�е.]80�B�dS,��D�*�{D���ڜ^&�oП"����y&�����"��N�����ޥ��q@ߊq�o8L?�%����0���;Ld��_����;��
�Y5v���+�x|3}��x'����q)���J�X&�۱�!�J�u�".VS�P��:�ӂ(��3g_���,������sOi\��H��A�L��r�U�b���UsՁ�cx�iY���f��w����N���I}9�0�w/����m������^G*�~.ӻH��HotQ��¨��NGd*�ι2ߤ!aO65���jn^%oׁ�t.`G]��>�}̤3�A�Z���zp�ܮEs�V��8Xk�q�η��)�6_�pD�㒌)�#Q�%'o/��g��H�¦{T�h��X�x��G�ӏL@�*E��Rө�.@hJ����{��o=�����d��/�	��c���"���[�Y�r���<�?A<~�QxA5��&"��2R7�uz��9H9���!�w�5$�m4�>�/Sq���r.�ķ.f]+T�l�o)_�/�Xqy���$�$�E�U�Z4)ʽ�f��-,iT��P�U����$!@��A;�����OP��x�pBB�@oDݐ��6�N�(�_J�g'R�������@~/͇��/����#;��Ȃd�H}��^��`���.x�&�n��B0:7�6s\��#j��T�J&�_Ό�o�=�7�?7v��~�ah�F�"J�>�p��D���G(�}.s��_9�a����=T� $-͆��Q��/��Ge>���us��d�+<�S�6x�x�X�tj	9ߎ�ٕ!�w� ���P��U�u���~���/�AR�M�ֶ{�@f TKe��ZAo
/��ӓ�����nKf8Cj}BdxB��j����w�s޿�u�)&C�<l	���G�oNHX����(��3b�78��B�f�ņ!�v���f�*�:>���/�J��@<;J��WK��8(<�ak6��H>T}ꦦ���P��3�x����q�f_��DX+l��Λ}Fc���`�=k,�r�s`��6�ow�t����:.|Z��`)�>�'.��W/"�N4�͊t�V��h�����3�	���5�IQ�ֽ�c%d�8ڈ4��^�k���2텦����M�{��Q�!X9T��g��l�nbv�����	�Z��Wx���n��I��\��)�+�(n��:r���0Q���]�ﱰ����"M6fM/�P��0�x�[k�+29��ہ��JA�Szv�+�N.M&s�f6�5n��	)��e�?7��{�DJ���LX