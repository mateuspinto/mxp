XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���t������N�Q�X������fUh>@�`�$�h��9��
��gaj3�?�Ȗ��uj����mD �ઐh͏/�Gk�<�F���vz�zM��wvP1Gj
�;r�Їo�?�x'Og'O��7���@O����v4�g�G��@u�wr(�l��<d�I�ݬ���'�e���,���oWj��%�IY�]��Gh;����Ɏ=(�3�G��C
ȵ�_%}���n0V�Y�[k��k�&=��Z�s�[�mRՃ�tl��)��1=b3DC�ߠ�ѩ��a�+kN���_}�̫;fU�q���4����ەW�KT�<�_���Z��Pc~ϡ��<�|?(�X�7"`��RL�Z̲R{{���.P"��+�=TL@ׇ�W���bcC�x�50`�X��C�=%J�vή"cl���Q�E�f2\vԤ�zG5�{Gk�-��0_�*���2�&(!v��$�p��;�@��}��z�]�!�d�򧦬�/}�~1���R��F��vQn�SJ����橔1Ou�vC�"���l�g!�AH�R��!;m��w���m��#`Y�� �?�����?/�%�/v�u�?cH/X@\��pmY�}9�&}�&��+V1>]�r�r><�B�YZ>W������~�^�Aq���إ��XG�[5`�̅@w��R��/�<�M���oY�Z��1�/��h�P�q
���u�9�[�f�6ߩ�r��_nA�zp��6���D "8+N�O���O�Q�j�>�Dy��a�Y��8mXlxVHYEB     400     1d0��\N?}�\�ը@Y�$�;�����3��.O'Ef$~�ɪ�0L%(c�)A����&��q���X[ݮ��O6����2���ʫ���\������jTm�bH�.y,�)	��l�(�[fFϳ���E�W���_@#��E"����(��'gG'yȅ�["�Ŵ���"7�x$�q���UJ��P��p��í����DD,tt�p�v&F2;O��͕\ܙ�߰�(�"���<��&���[����i�PD7F�ɠ��9�j�=0._1��ӡYl��syʀ^㾳��t3��k4U��ǔ ��&t���ֽz_ױ������'���7828 ?ªK(����jm��sΨ�7jYϭl\@:Y�a��M��e�c�k)� �j���'dF�G������߰�+�Όٶ��O��Ʀ��Q���5�Z�\���#�类�\.�Jiu��_��t�D��XlxVHYEB     400     170��Q�b����V���ҕ��e&�TEJ'��z�o�{����ڴ�y���%�x+��c1h2@�Cޖ~�	Y���2{��� ��Z�o��9���Jۯ�l���B[��
*��!D�5��Av
�1w�cZ�`�}�������	l)�Ug�nB*Q赸��NK���Ã�[ޏ~�Tk+<���%��p�d�jM�f��f�P0�h����h�f���"N���ڇ*�Dn�6S#�r��e,�e�l�ӝa^na/� "�kj
J��bd�T,�/{�m0!!^*����7���`�G�z�!�3N@;��șLgX�y����v�앖�,LC9]�eg��X����B�P/A���d8p����o ���XlxVHYEB     400     120�Ɂ���$"�2�c��VG��#	"(�����Ҁ��("oG��#ݖ�=�D}����q�����8�c3h{i�Ij�?�$1,4��9W��Z1oA�U�.�(`29����U54���ett6�!u��AD'���@4X;}CeG��ȸ��PL�ψ���U�LΗ��$SBE��� #����,���#�i�Yؽ�4��uw�+$	������+7����G�ˈ��0���6���D�;���(W�VQ]�����i��%.4@�A���ܛ�9��꯷�0(�xJ�'P8XlxVHYEB     400     170~�9�3 'Y��'�U�f�-�����ju�����F�����w��<-U�b�C��*���Ιv���j6N� ���#����>����X�}'pﬦ͔����g��=�lC(�]LG&�HG<�W���^:�fB>��ʞC�
$�X$�c~Ɋ�CPk�.+4����\"�ic� 
�=H5����'�e�O를2kQ��4��ct'��V��ͤmn�\����w/��y�O
O��`���3��*���ѷ��P����V�,*'=�U�����~�վG}*A��g�n	q~$!��Zn��MAZ�������7ZNA*���s|Т�'7_�3���}mnXF`�`�Q�E���S��\�J��u|nz�bXlxVHYEB     400     170ww)��Rot(C{C'������x'�3�A�1��$]k�����<��@ԏ����W2���6�v�n4��nJ`�ߨa�_���)P$�}���q��p؇ꊗtf�!�����T!o+�D^2��U�O������~��Jv�܎@��*Lb(������[j'ze�IF^�c2���Z;�/�,ae�A_���%��m��C�8*I	|H7{��n8�uEq�� ����0�����tL�I�x3q�j�ȺtO}�)<�������f�Um"����v8��7K8M�����,���S�S)�g�#�3*����Z'�
��xv^��yj"ч
vE���x�������H�����>�
�:G����$��XlxVHYEB     400     140N�֠�Qm���1�c,Ə��ؘQ�bj#�y,T&m���X�H�>�"e�>Z���b�v�W�
��u�k��Lc�_�m��hõ���
�jĭ��(�w�p�c��}��=*� �B�0wu�ԻT����^]LB]�j�����M������%�����K�j�i�jI��n9ڷ,f���m; e�s�m���qPo��M���^t�o˴W=1�tQ�Q�^}�Al��o���t��Z�u=�<�����e�&�s,�ON�>�{V0�tӨ5�lELAD������&�Tg5|� ���-X|3	L5}�ں�k�੹�R�D�XlxVHYEB     400     100@�(~���؏]a���͕����Qz��+@�������!�?��[�[S�Т�D�z���}Ӊ����?�I/Ø^��^�&PGYL�?}�D���<�"�,mH-3���k��T���~�m�Y�m(��C�G
+��΀�t4�_�=��b��WfM�~�X[&��^�=���#;!˔�;l�U�������JTq���L�c�>�b-#�b���#N��$�c�y�5��"3hM���a��7�#����d��9�XlxVHYEB     400     170��/����ש�]���Js�z�~��~s���I! ���Ź�&٧�lqI��=i��-Q���m=�6���r�$�{�������^ak@�c�+H3�-�V���9�t�y�ѷFX�pv�l�b;��g�GOL�,k�g2kGs!�2q%�(_��'~��+��
���#͛y���]a;t����6�v��iV�Y��B��f{P�_h�*x�{�ȭ�J5�Y@��OINS".u� �jq�X�!n�hJ ȏ��A��jX�O�GH@��H����<X������*�s���q͋՟��zoȫ��.�b��Y!�fZĐfŊ�[^��BL�c �i̵<������ܠ�_R�0��	�O��XlxVHYEB     400     1b0V2�ۑ���j8��Q�7~��-X��*�cV�wn!4}������n5���O*������\��"�1�e��+;c�Ow��� ���L�R�|�鐯vm�32��ۈ��U����'��i:<X˳.���Z<6��>�"ÙR��A����ϻY�x�N��E�y�Wa��|���P8���Ȗ���Q����I\����FD����F�=�Z�'P�lF
�)��k�h��;�]�r�)|�L9 ��ovr!�a:@G����[-�3~Ǔ
�Bc
��ͷ=�xS{�(G�ݓbA���Q�����h�V@o$�0[�Eᑭ��n+4Ԓ��R������杩�2~�{�hp���G��;����q����SpU���Ӄ�|��MD��/��D)Z��{7�WPO��d"9�d̢��L��͍��t�B-���K:Ӑ�z�X�XlxVHYEB     400     160���贆g���"q����+�IbI�1raЧh۰��h_�Y72��j��⼜��܎��_�tp��R�e���F#���	�Qܗ/
;FL��r����G��f2�ïhɚ �"��τ�Le
��n���@ ;��p�"8�>�1�:�8ϥ�����rc֔����&��BT:��ޜl�ܔ���_o��w9�4H*�`�]�Y�i_�"z��?w��"O���LJ��Ty���ڽ�w�A�W�B�1�R�e��J����k��/�'`�p��MB����V����6�7rR��^��Z�͐5/Rΐ�����Q��������w���67����N�=z��ӜxXlxVHYEB     400     1d0G�K~��͟�|�>�rNB���G���ƺd&a)=_ ʚ�O$ٔ�zqT/D�jr�4��R�ߨW8l�&Cl�;�}�Hw��+��w�Ұ0�`�]O<y��>�>t��݅�?X9Q���pB~��R�Da�� �߀�/�9���
ʷ����%D�h�y�+%�7��,4�O��X"�)9�"}tc[��w�\:�V6P)��g�+��m��s[�-s���k��*�2�P���S��IVE�d~�Y҂5S�b���*_���)B��}�5n��;2O�T�L�'-����;��1��'��'��ʅ(�����p0N����ﳥq?4\�=^��t�2I�i��u$�3�ON��^@'��O���=�+�[Ttcuv��Zf�軹�'����Ȣ�6�7&H!��:'/��u��۷����+��oHX�Y&��6�WM=��t!�U�]M�{����:V~i�7�n�&XlxVHYEB     400     170&�g>i�}®N3�]kxd}9$�L�}xEw-}).��^��ޭ2[3XG7m�U��Cf����>�u*r��@�1jbAd[�_k���)N�OXmϯ(�:Z	ָ�����̉c�C��
�P��
s��L�v�ruU����p!�:�rt�^X@R����ݒ�-�^��V}4�Ou��Ҷ�y|L/���P�A� x������ �@ؾ+O؜���X�*1��,�+�{��
r��ц9�Ҝ�	RW���e���P�w-"��cǈ`c�e�3�*
ǚAfv5�3�PA���y���7y
�{o'�U���6�<ĕS�%��n'�ճTR8OLp8#��w ��ܩ?~C-ܻ�d�l���L�^XlxVHYEB     400     160�q��c���}��}�@��0���
�5���|*K���,	�*��"J�[����4%��-et���/O0%��5H&���,�o�H�m*��i�;�
p��n�`���p�����l`Bkb�\���:v咵2��A8noF�[�85�hKinIC�ϩڠ7vtЯ�d�*!Cstg;���R������Q���[��(� ����gM5�VyM��]�s���4#�y�TR��ytLY�D�(���w"~����ǹ����$���]��G<��	�pω���'�sq�S`��e�Sq[�b�6��FL�s��8F�����g�u��F��%��q�I���4�Ћ���%�4\XlxVHYEB     400     180���'�{ �c��֠�P(m� �,��u�;z`��T�t
�Z�+�R�:l�#2�N�v�k0֝���<f���q��G�9����[$����-�Uh�왃�1ߚ�g�#ac���7Ɵ:��u�iPBv�}}�Xh �ևfT�Q�PG_�p�Qߣ�W,B���ވo�4�V$��𒦰B�Þ��n��#?%�\���N�?�+yП��K1Z,P�{S��O?��P�~��Ľ["!�C3�J]�yD^ܢz��,4ps��U-��]�m39ە��L����"�^��0���9/S�dnwh�ب_��-�1[n3���C����H��Q�s�}|��nي(�É��f�C~�ْ#��5VA�^3����4�ae�A��l{XlxVHYEB     400     130�֐e�?׸�V"�>�Z�������uZ�aFiXQ]�w:oh���E�P��5�p�g˨�K����;�Y���haR��/v��,�GH�}Ա���u��_� zӆmǯLP��n@mG,�)���|TB�� �n5���9����p�~q:�#�e�$�qvG�d��M��/��+����W��l��x�y�\���r����:R��2)����4�.t�����Oi�o��D���\���o��Rm�J��	:;|6MYg���^��d���^�)�q�5��>~����J �o��"���rO.�k�XlxVHYEB     400     160��xc!�a"�)r�|�2��nZ`Ҵ��W�G�a	-�����Mu��F!O:�R$و�Ձ��H�iM���W�����O�ڹX2}l��9�d���n����Fd R�Ny�b�3�@&��_
�y�eP��'e��z:<Q7Y��q�v��;��m��\
D~�1�S6&����I�\���v��ns�
k�y
N�d
-��W�O~��M�/f��K5��
}���
�+��^��>LUi-�Iaњx�c��K�b���3���sڊ��l*�1��D8#2�C��?�}�F.w(D�.#�ٺ���Chg77����E��On0oz�A���GQI���g���NXlxVHYEB     287     130H�l�:}�u�,�1�l�m=I/
w������Ǜ����S\�/M�KT�L��IPB��M3��BeBe��!�����nk̾��h[�>�e��|>��@H�M�l�C�x�P���!�I�����2��{��؄tb��x�)�*v��^>� �'�@��Ӑa�
F�gO����]ykj	8z��1�l�f��V��r'x���t��BK�������P��-L�c!e!��~�K��NU�%� �,���\n i6P�Ҧ�,�#�(\l�jb�3��,�(��=#�U��d;���