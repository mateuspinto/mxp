`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25696)
`protect data_block
d39j+Tb1Ai30idw9nx5Uq4BKsac9/F2QZTO5I7RyXbMT59QmTMlJWX6jVxbbvpi6FO8KC0jKRyNH
/+g8q7CmP2xCyzgGrjMBOfAUdjv0jgns1SwSIzd4bv/sRwRIhG0m79ku55g3CX5DwmqFAgKoIIZ2
MYoxwgS1SomheyC8CIaRWb31gAU0almhVXS9MxmYwkuiIC9x9tZJl3DD+p7a/EwdKnCqnE5GSMyt
cjyxp8loGDYm63zDe5ItDZ3wUEYGNE8r6AFe5lSbfovpUsykAlRYFLSWkAztr8tLt8HXG9c2GfLq
YSD4QJItBy2ta3d7Dqppbab1Q7+XoGpbXIMwA7En7ThhmDyeX7LHqdui02Ccm7Kojc0FOB6DPGJr
Gr3nwD8Njggf1kKwChuga9pd4+++LEyCrs32rsCXLc/ZOxfuKxLQTpk4EFcLoeMQnUXBOxXCRBO/
h5L3eD5n3djkFHPuojKcVy/MlT7igeO0ID19VTcypujbgpiiL8DW8Y3iOn1q/vM5SXxc9Gh4R6LR
thtIqohv1odXz1FxqlWvhmH6GOShsD1cZZvQ1WDuY4runzrogBPYDPabesLSwPvejPpT7897PMnU
w5Y1jaT98W1EXoVUEC3Z0nkf/SZnGX0qS52TVchSShgcUf0aBRwyLLIg/SEm/6g/BrgXob35UaDK
M/hlheHR7QhXjs7Z4d31g1OBSygv5A6CvyA5aDW6bettvS7oWZvWrPitNIoaiIIk7q4zw9PW39yJ
N9Jleciry6qwJmDN+u0KyRLrbdSLAC9tOwLne7/WvdkPgiHcLTByU4jg0mHwHShF8R1cVBbggpqy
SOWjTIbJW7qt0+ImemRPimeNkwAkTYqGrxjta63j+5kHPmZE9R2AniXsDiCJ9UninPBEocsis7o3
g0z2XUP/eIfMFU/O09ghv078jR/0L0+ltShcZfdH/C+FA5Lt9jJR7kSPc5nn5hbaRmUi3AwXy+61
R/SaWgwS+n7TDkp6lQ6exfzmgy2cS1wHlOPGIDzeGOz6gp2QewPbmgdhgbY53aNLG0S8mMUyA8z6
o+bvHhdoVk4RKd5EduPKr2bNi8q7dGkJw4bqcBpuqQ08L7NDAtZE/3D7QfY8vgx608A13r5E9A1s
VKhxHjcr8HZ417sLuEnTgmi6DIAMAHtj2NYv3Fa7t2sX4NKTXXhAsE1mHKLKF56gG4NoKyuiSbNH
keOwyBpqRaCZu/kZk/UldeEvuHtbWi9qs7oMRFhQ3aJR/7WtzmQcfVHWjiIGMorL0+pKdlraVu8T
yrDZyaI32Cn8acETv9Bhoq4p/J4beB12pUXbXZRKouneJPVEguHG8KMlXGGFNO2wnSrtsceVTfVX
5yrnLyuhj+MlxbvdQQIBYWCVM27xrczjTd8ESDuoeO8QWYpOaYVTVqJyHnS9q8ED27pIq6lO3ENA
n+6NwOn1FPFa45M5xo2Bi9RqpraTbKLAIBgWJYkJAXm4Mdn0OHi8mC2VSx8Y9LyFRG72wi9pmJli
Ki4EdYGRRHv4S7Xzm7Hp7wkdvv9TKIjm1MRw4Mtj5ziTawMYo/sDjhR8w+zfsX7TJF1vVTjXtFfM
66TcrSp057OHLMVTRya3nTpIdJ/pD9UIUuANFBrk7PzwYrdqTokBxe7F9S6HTopWI2ro+L+JUu9j
qZinLihB/tKAwQDPcHUqbXx7wEDaYfsjnRnW5u52bkwIdcs/+hZaXcoZsaKBaChEqfX2Tx1AHFVJ
/Y0o2kg22dYAsnWzWaNBj4tcFBSqCv/xe//ZgyTbpmMjwJuOD0qXURyACPbT4SpRxWgixO5F9Gan
FFFcBykE/MeR83pJUSJslAGFQNwtT9EHwYDpbqm9XIXFtjCyPr6fSVMlAzQa9hg7hkmDMmtH76mz
zvODfU7E8TIfhYN4lglP4tDqSmVDqlf9QBUETbepOpPUrvRMxVPTiAhrM2Lj7VLzEeDy91ph1hfp
5cdCMG9uO0JDyZxxanhFPN26MB8s8ZDOtE+4zVA4mBnqiTBt638XOEh3vO3mU7m3e+JWjW57vypR
8WGUqsXozkqt+qIHEfhnnzw2qX1Oi9tqCci7MNA9BRqloIhanPi3ZG9vWcyATVSk0sdMq3RNKOjB
glgwJ/NfpBOtqR0PoXziwBlvzCz2mNtiLLK0ZU4fxISnwqb9G4LD245tCJitaOCElZH010SB1y6K
tdyXaPhWyDkNHujEaJeUwvL/YDv6CUQsbfvadFrH8jYQAs3CLQCXhSpTgLp+gGSF7YEqtbFyDSNH
1givI0GdJlwQHZnUdJu2MzSDAiZe7edmW2iBqXWCMzKrAf929i5DPpJTL6TFSqjOCmcv2F1JQOzh
de4IJc5cN15Ab1GRCGiccMg0lsUazD+JPQdxWsci+RLLtmak9oGZBC8xUXa/7SiSxe1kBqBJ/nM1
6/MfUWT+z2iYYekvdxf5krQ9ZONg6LQ5w/OqKDkOxXYSo3Z6tV+nM+Sqsc8op3MMj0k9H0hXIsro
Jh2yGqbLiQGN4h8CF+28NpsKynptg+35hw0GUpr7hGX3vyqC2yDR0XnsqAq0GoUPMOuDjqavnjVj
0ZMQKqPgEzoPrbUQjG+boD3X1gDSed44ikhPzv0WxWolmkLr2IZBqwx+apOeX54AhX5i3h4U1yxK
wPw+rBjRvKJ7WtXzXiqbU2uzQdRfpHJ3NpgLPDGxM/gnep0GXOvUsWbCIGU9aaU9qa2nuUL0lVLk
DW4GZhyMIyCmQ2lb3KFVsxV7mkvL62yqIjygeHZUmGAy1r+0ys//1VgasovsTPEbN3mVfSOsmPZb
F2BAGTpxZrJ3N85Te+tP129iNu9o84Kx+dE+b4JZ5c0J9cxAcqxTcbCNR6fvvfhgv1/bATI9V+Sf
oUytE0y41CIJzT4pk2KSTijd+C+PEPJm3VhiaQsDGPEp3Uj4ZaXxCVXhHBGw42gc547bT5WWXbz+
rzEsXJ7JaLFxaxSZNi93wkn+tJEXEfadzP2BNnpVM8MS64uZtAigSYx+29F3rRe1MjQqYGxHxv5J
lQ19mXEvJnpGvXk/P4p7//EXZvcIOWn+oygNHadoEwxqRiuDNKPhw0/3BEqgq3B7FPtjaZGRVrIH
jgeV0oNEjnDtDvXITE65u2piF+iXgVdg9zqrmFky0hLUoX7e95B2UOEHAcad+HzK/3rcKqAJCmWZ
e2ZfvMuZrpvSWddTvcbBPc+Txc5d5nTPIShJHGD1Ljk5lvRTQ9F0OvkDRTaxhAa45IlrgbzTMnVw
UV2ekJt3Szdu4OOr4JbgBUHGllJp4ex97ixGPqX3f1BRDBdfQgzOseVIYHnMn7iOg72MdwS/hixp
MxELkV8rdQDfTgCuzeqQ83I6Td0CX1851iXAophsaQgEBFR6nGpaD6LQh7DFhshLqKv8cfhcHuvq
6XJO2qlm4731hdc/+xreOwQkRrAC43s5DcXPAxTvC91LoUkD79CcUGWQk5XsNixtPq56HhuxEcw+
sTgTAWlyU7rbGwvInBtPaXrkpixNPmBntKa8Qi4ObdZRAJh7U6ER69e8RZna3KHVLtjUYV3maYWZ
VTpSAU/wNK7Q8iD0nywsUhhek5VbKGz5J1+Zu9MJVyxb6xCO/EI5+CRjq42AgqeG6U2BNMSRYGct
aOjP5n3cPiRF5TJzDTjWfYvV3xsBEd0kEqEvL07zAi0UYdcN/s/3CInt0luLdr4WssdajiEi0rtc
yUS5EC0Hr8RnR7IN6FM8k1dJf6WEk4PimZPKMYdh8omDGNRYJQpdb2joSZTbfIDb6AloqbHcPkjy
VErgtD7HsjFErmgY090xOI0aUG/VYc9uGjv1kO1wJfAyruFBvZXPpnUbhrcFLX41J31GSo5mf13d
6GM5bJeuwRI4nV9Am9vt5fIWPw6x3iBJA9kbQrAiHIxKevq9BzVdGx2aUCq1UvaFX87p3Zup9WWc
t1wihE04YsraOMRKdvKWbGDpIXZt8SWgzuvvmIhjHko7v2PUXy+92rWDfKgRGWurM+f07iMZEo1N
PD8YdREFKmhi5j3CPyUREEu7+eBWIOaehZXD1H03DBC6k5Fy/jlW1n9lVCO6tE2lNZ0u+W/IlKTZ
Wl13MRCwPWXQruXuOnFGg8Z/WJRtk/c3snNZrevAj2aaYbfPB7tpgvN2NlCiNC3NBqKoiez32D/0
6VXSRCI0em0xDa/DnmnBrOMgMQK8IJnCwbS7iPfBq7a8D1Evt74bH8fstVUXd5OKlv2QwrNgPF7S
QC1M8GUbpJPLOx37oySzLSGzpFrZY53S4ap7sEDdzGEtraCEuIgrzZJRdDc/fv55OFLKpi/3WCCI
DukK74FcWwPn3dHf8WbyZJ3XDAVB0zbf4TFPRpmwdtiSXXcNJ28qWJmZdTcXvXfe3t6VLVEK3kbD
zpkpIWgbPfaQNwHiAquHAi/DsuZO8wqgxDJDz6yRCB4Zw7ZijvO7TChGiVVycLlPnkdWKZQ/tSJg
PD9QJB1JvAuVQU9O40oSochC2kt7SG0XeAU07ZQpRyY6e7ULlVzx+LIuM/qFMKJ/lqwuUeByFrbD
UZS4CB9F2F6N70j55pew9ttuC1ubtZGpMQ4QXGMLxIfMGIRjg4ex96lcJacPUj1OHlMqhaRn/oN5
Q+Hl6xVr8XOcakrxHUD/a3eA3XlilaJBNdGJVXn7l9JPgsICTtfj6tVTrMjylqR95eeHyzwPO96a
7Xffo9i2xks0DQckO2qjT+rg73HMXM2P637K01jwWZ71f7Lj+Ou0isgl9BAbB4so1FEfgVH8046P
Vcco43fXxocseKR0sLmbBqBD3IHDnl3nTdIiRPu5d3qij2Iq2PoCkKdz7qt1mE0ifMAXFbE8CjVv
nm/FUCT/8Picf8xfCyDdxAVt1dcXrAdMZ3DfwhqverTicMVzVksgUcZGpepZ48QuN2Ptrax6uU9/
bIhLc9P3rlQJ6k/tH0FfFxQjJZP9KLYHVgEfu8KHV7OCAZvuFDsEZmi7/7UA9aRp9eY8/3aeWrcb
2yJjTOo3zhg3VY/AYzvqtu3G7K7KxgdazehwgxAMh3U+9cvB/+jxk6iLqhIemt6j5YQPe6fI7WNG
Lm0bXRfRvV0itSd0OqxoG3arWQMlDbiTyCgF6iVs5ormQJycAERm/VCk+VAiW2/6yYkMCt7DGqRp
HyCtkBAakKopPBSirIwt33Dp1swcmdhetUOHIVSeFsdSVSXSi5jsrZXNib4PcmetROJmjeklAY/p
zXnI3tvqfASR07qWj5I0H/7dkrHj43AzWiBizEk+L35zr9+oeRLwIMbdYQho3WDRyxaGK8Bmgz4s
PIUaiawDU7Nrw4jAM4BG9XcGbrJQSKBrWfdy2gIzOuSxZFUn6qUHKEvJW3ITEsrl3dHJjBX2Gi0+
ERWU5Nq6bG8BRKzG30bqgZ1jFhZo74dBtmzE2q5rTLDxtF+MlFvoaFzYeeWMoGjYT8IKgPebtOGD
SBW69Hz6qCEv7mtWrM8AmEk1y+u4sUyAPRtn8OXiJWzjpzeQW0qUOaWGEGlg7CUOkvirZYJ2i7Wl
miNUeqPdIsZ4jaarIwHX8UYoMwIAy8SkM6Zr7cw2DIl/dpOXkNTH0koHY0DeVTUsSZyTfnRPGRuK
Yy8ISpU6qLg27m8IfcpDh5nv//j6BWAfS7+Fho5Unxfdqm1J9Q+XPUOmLE8ozoRMikZfFPoZhT3N
eLm6++ek/feQIXXb2V6CWbVSy+Kq1pX5HhlWCmBixHU5ih2sAai0vm1mOIpt6yJDJiBw7go7WITz
LWjJsY22G0j7hOhpIUhyglj5jnOK9Bo/Nz2WGbsZbPLvYOK0bASf9yMc53QZius5eLeoEqxSips6
4XGwuuXHCqL2YLSuL+Cj5OKS4F/wGrK07Pqv3StpJuhf3M8S6q/lYJeCXnxiAt9IwbX8+jTi9BNz
bunoz/UlFsBj/msIpV68iY6Ra7vXmVMem5qjJp15p728ydHGfVWubab1+c9puB9fV2p1k/wlWtO4
rYlVTrsQYS93sJUEGJvGrGMcabo9rZLUJYFXUl6+64gvYXY02giC1W4cAdL++QOvYk8TaRRMZJif
/A0ow4LCCF6bjtdEjUZBzmKKxAwemTToC39b6QCJ+/fX52rvIQh19XyOO2G4vey9Lln4KhAFmhEq
7aCGZYOjLLzf1CgO4VhJegOzLbZ/+1i/6es8aBTW6iD0Ek+E6uNF3MJNjr59XKlhQSyT9ec7hpZ6
3hEs5+ykyTAFNqEAWCD7UuwklY5fwI/k7S/QsNJm9JBe5fb7MFyDkXAhJPm+byLGLb3sXk4HvjqZ
fFFnmKNBTyO8n1CqPRBLvZWchpwqj7QdqcgPS3w1DQ6l+1lUasyAfI/smSoVA14S2nqMyzsCw91D
7nznlCNGr4yQJcFDwtOSUCZ/IGzKZaFcOgb9g4aI8jqFPjPYsxKMp6cHRNbUqaW+qSEoBhbP0qYB
A3tWR/gFjsNi802027+ikHAUJzeK0buQSRA87njkzOOUCUHv+bUUvlUkbSz03GKm4urE5osrnfvn
bXVUkbHUHarpYwZsmSrYh8HAmm1Mlj7WBcM5f9hBKtq1MoNakxplvZaGhYiCE2pzS92q8zUJkbko
O8Qk+sqy0CHabAouoQ2MTyxOr9HYTTR0qHa9q5fb18NWB4MJnLPcsB3SLcXO2TU9A/yt1n3yCJJ1
bUPcKuwlClFtwJrHga8QjK/1yjhVk3tSR4zVHEsWwnM6Ta65TekU4d/SNCLZbf3pCnuiCtBHjvnT
g85zg5z2k4xU+8cx9+uSDshDibG5NTNELQRDyRMZZq1yHQ2KBFfSA6Id+zNL7IM5/ua0rO18auKj
jI0nKZf7g1iLH+p572dfROc/O+0R7xTht/WNOuQ3HdX5XSqItwQ7zWmSpItqxfYGkP7j/mHlciZ8
PxFHcLIZnUKMVRyJvGzvHIsKQEmy22Ikxa92Ow3FJ+9/rmxN2Rs1lguOrQBTQuaVS5lMV1B9D9Ti
q56VDMlUZ6bpC5FWuic/7X7xLA46VGfTa4LrP38DF4g9UAQv4WTHKN0JfSojWN2y4+mFBUQJkmPC
Q4lipEqBRP66I9IiLfvCp2k2aoC0JrccZVfw7Y7NxLX0Fn4VjTBblFeWm2BIs9DEg7SHUpbrTu+N
QctT9vxvJ6A8ZI8JNTCGczenjWGIdTO2G2mxL+97A0hDIXGtLGoJiLj8M9CWQxHWhfHttcVNjoz5
W8KFKTHMDbGFsbwWMSlYF6gpA8nUkQ8+xHrh194+a9yPmaSSWVCjuunmPVuyhSgNu1V0xlwjqeBT
6I3mulz5mg3E4ZZzvqc+TYcstAmiJpZ+SDxQ0lZZOrPS4bj0yyslDIVRFphCi3Mjn9BwBIbApcbk
sJY0r6DQ0t6AB1XidHbhPuOq79/kiP9DXYTDGAyclnChU6+r6SW5t4FZv6i05wBVX3rnK9G6xsgy
EpO0YYC9cRhS3z6ZcO704d1ZjdqdZCubHulMj948O65AMJ0WSB8/4CW8JPG78IiYP2M721a2hflD
QQ/vlACGKdPoqURJpjf9PZTZPto8D8j7OJAo/VFk72apc6t6L6UTqYyQf8JtxI4JZ/6p4LXTnNxT
RNNXLMcXI1S2H4NQr8qyMUBEswx/wo8ciDFZe0gcTi7BI9uet2jry3E++Vm62hJdRoYtd1GPZQ0K
ME+aavHmScevV1iAYLXOKgQGie7ERYmc1QjpWRmK+VIGhEly1MH8tOJXl4KoBlZQYtjnjWg6TS+b
UppsGCnfECJCXYtEMtJ0uFszLi00HhNV4sqgAEpRen3f0FZP8MG1OXb7ErXw3tUTJnKYeW2kNbIe
+PgVYWd9fOa1wF+LF8pFUXA1MUhvELBN5TId2Gnqm6w+hZIFb13Bt/5mWlojw8NtRdJYqWBRJcda
Q8puB7agHPGJCres5TsRMOGMVYRTenVWYPm2arPwe5xmD+VY+km2rZyVcURVm0wOEw9hKp8Kz2zf
9escncAEt3Sp5iu2AaISUEa/7NU7FRv8zCFNtmhj1pFyyQx9+SqTPxj7UhwEZVZqF2LxLM5TWLar
aFbIw87YdCQVh7XnxJhe4znFO4jnLDb/yKBmLazpYGZb2ZXYLMZrlZpjvhQxM/S4tfTfbt3jMU62
L/g7z4BQpm/rBO1w7sEsswXXD2kHNwE4ip0K2VBIRiatl8lWGT46y6INpAvweCFDDb5jJ3N2S7Go
jIzSMK4KrpWlMfZV/yxUHwpYLx0w5wYuwztI+1XxQQTNoeXeqN1yv1LbyEdsH8/oGlaFHXBpVSa+
5pv1+o4BwJdiglaUNVbstz9Y7kR0FRWXQUuxLbLRy7EiS7Gj5CMGpIHSu+0zVHjO4T7Q6khEAFff
YLK08KqSGjLLEHz9wqfETfsvP4OoXv+Fc5AsBCOzZyz1o94fcv837PXP8c4qQ/s5+T75Y9bYVv2N
LxOFzQYl2fmm4U/9V+oP7O+IM4iFzAJXX76/ZxQ9X80b5WRMZLBWU/WWJNSQhQSjdKXzxtd8Q5UR
1OJyLuNYqg1SKOtONMzn3iOb+KghHVp9NkJSD8NIxCLtzop2pASNC38Pz8s3cCvnoYZphz67KGbP
hBJF58pLUFDnQ5qDbWvve2xPQEg/eZGDS93ZTL0k342GRTD6z1zbqMQw/6Ca4h6h+qhA1GJUdbYj
UZTalp0G1NJtXIdThLQMLoej3RnUDilm8wCo5R9vZH/TaXQ302RslPLM4LFVKDcz3N60lsNv4/K6
akC2Onw4ZEUUZ3aXgaTge8sFGCTKdQ8RFP499GiOZq/4lHUx4vn28n4+JRoYEzmrC7Hb2amUfBcF
JUIX+8shchqSh3JQYdvKPc7cQ60QjyaLPKKWjlbpzUzx6B7Lcr5YiAnjPEUuKAToSeXPeiu2mKxu
jXdlwIC96gnzf76RgTTuZinzwTGaDH7Kapwe30I8BHqn+t6uCCaaju6eQpPy7lynRVGIdp41ETNB
aGGROR4kRX5JA+rUniG5MnTSt/du1AnjopVh66TzvugtKr0R/7M0WSxeJowexsL6UcQ2ATc5vVlv
XtV3xcuZbuTnaTcj1BUvLhnxjG9iy+FH6EM2TirT2fq7VFKiF2Yf3GcE7zGMZhofL1l6SnhgG9XI
VGieesJPixX3qkk9OFhnRerHQH3rv3bfwveHno7943xil8FSc/e5IossLeRNFg+Tp3m0N8pO/fPs
hd7vmtn0WIGAXWjTa1kFi6wSgSx/J/pqD/pevOCx+TbCgv0SvwyCwq34ZVxXUk3beyRSYxrr1v9W
tUDvy1f3GVKlqrxmZfeW+4cOuHkTID+f/bw1mVT+AWjYe161InIlE9QVm4iXAP7Vba6wlze7DwMi
GRCjnAmz7nIKNbxpMZAlLBGb5VsYG2qLnrcxF3rHaqX/5x93a/aHfBSruMMxUpVVd78W7+ug0+r/
wdUS3BB+ElemkxAo74rM5De+ck4SrM505xafoxR/B8+bKdt5Jtq+1/CbSl/MYFjnLi9mSxhL4Kqi
Tds3i+P0QipEgyzKrbYg33CNRxk3f+3AB9jKSL9KtbsuJ8DITc+XfDg+k5fiYLHTfMb9zw/1hY1V
W7eGP1ylgTNS8TP+0zA9Nvv2l6tVko5VcOXVdRTyNXCja73ty2WV3PqI7PMUS3haHGKj4pdJLbrq
sQyWZbcXNeWm3HoLqGKuEbyRv4L4s76LIs1eo6njPrQWaTEUfom6DEoHuamuytPBQ8nHZnQ96xzO
4ku1oFM+pdCtPpZuff2Rug0cm3cP+0VvpEUYJSqT/AzBQzN9YGVQnoVPGia5oEykWfFVggeNoV/8
acTSRLDnIVIeaVgc3tIfAPZmUimhbKQbUyTb3PXmx3Ro2H0TheYD0rBzWETZAnQ8k3UvBW5RGAzR
txE1YMRXjIoqWGFNpixauJd13fiabjEqZ7/mKBXKfTeL6mWkhU7w9nQOwDwmAru+sS4mzGPXzClA
G7akhgW0lIqJwkBpmS/oT3g6IB6paaQcDYhBFH4nb75aJ1fvmSiyFRZOPmPMttZOy8fjP418pys1
5IfnmUeljE+LkiaDjw1DQmitA3AGukMvPBvvevVosx3dYduaApEK1t8dkcKZFJ58Z/YqNJJwJr6X
pd327eLs/xAyitWuYuLpwXQ1WGOtEJuJNHyDQ/7I2KDbbuJkk7JPPrlWHv9KzmmNFQTEYlnBpI+e
140zLa09F7+2sRZsZyKVzrajonxNXvk1I2vttwHZ4YIJBgQG6sFtm6QLfx+29Wpu+6l4pLm+mlw+
GECg1rxDViYAncV0Lim2Q+sugFJHhMeF4nzX6v9zJG6iOFz1IkXmHqVTjx10LuKi/s1fRVFR4Vvu
ffEZPxLjizdNUtr72OYynThaTus2CW9UxmXm8tLD0s6m7L0E3fI2wSUOdEUhpQbKwTDrdjC7FBbr
nGbiDGFLRrt1zAsFZic2gLCQqw06o37p+jR+xhQiYLT9bcJWk4UuPCEIypsNltMLZ0XskMjZuj7I
fZ5rAF5f4Kc1gkQODh7AbOs5MYqVQFYKgTG4OhgRhFzXfmXRjYnU0MU8NjC7l0QcXockuohsU+12
jEPv6FKbaDux6bJMqAWZebhCCPBSJwAZoLo5grl4Zx2fS0H58DrQjZ3l1a1mw76jmyEIn/Eq3cub
Qbewl2WyloUsxE2riJ3WNgjTKmRUp8CQB0eYqLT2zcJJceH/4Huc+wdqImDSHKj8IHxeMiws0Mxk
3+7HVa+JnljW/kE6rKCKnRw3CtlC0a/H/YTGj/ix2usrunVxExqV4KIw3PR6iafdJC3IdJUEHjeP
P3qyCjOEoj61yl3iy4fLwLszWRcUMOw1FXi2b2FhHtJpgger1MOBFkoRRcN6vortysG03mNpVI5D
DEgA6+pDMLWuYuf9Sbee4dNMjcPb8WgCT8jjC5hueWHsU4nMiIWxwyilmW0jrMCyF+KWcpl4KZpj
9zhtRXKNs61+XzrfcTfkTbu7NYrOgrMK1xTjeuizikLWRTYYELhvnXxy9RIcKi2bWdUpOi+8FvfL
p4qmnnuWVhMTdNx7Wx068IGtXTEzWRxR1kalBQsg8cHLv1u7B0dFkCjZEgDBJmF8p8gIVydUiWOA
+bPfPHESWspA7mWSIk40KVHBTptzSHqo7tsnHo0JSXLZGbR1IIsgQpoxiKDjSWeScAlFDLbaV/xK
8TZCWDyfIniMGMzM2hghI9fDjA+So9gIE/uVIH8yruzCk3DZuQ25Lzrk9Tu9R+R9VSMnYWtdn8/G
q1BW2yJ7kbv0og24eo8O0F+SZSWQ7h0sYSkqcrvA/lNN/jIzqAY0tk0wdziLG/qT4EbiVhsTrq2B
9qrkGhBP1qCTkeiIDu7CWDVeTMYnavEJBNvy0rQFLtI2o/5wXuwas7pC6ZSdBsO6S29RIlAYRAoW
z30HHepdp5oy6Fhmrg5Ob4jUkzWEWIzz0baZwXZiNObGmM8Q6j2FqgRUtXd4FfKFUqHellpu+mfZ
DYADPSPLIiDbp1aO/JRmhiqCxY/gxqFoDblpPHL03ehIr0DudUBgKnk5yAfUIegM1vgv2+T9GR01
kH2VVuYrC3YUqAOpY89a9eA7NPzFXm6e4wOKeUAV1JBUr5/5BF7EWKMeObveYzVk/21dBicCN5r5
YUzBJka5qidwb6XEZRq8qh7+2ZhKVH8QwfBE9MK/80bjOdrJnbW+SIYbyEltrfqLAHztCDw1+mul
eOgKJLAY6xtXYUPai+jpPdDwHGIcdgR+51jfcAZEBbqCQ75ZvK1JreEWmoj+piKOZjN6YR8eaJBW
Rsd+zoRziOxk3rXAHANYrLskwI+eOmPS1GAV6E4PJkWv5a3OWqBDbXaUoT5nyBgl/1XNowKOw/CB
SSvc7zQWb7MwmzINieNDgL1CGlaNO5ISXHwfw5o6gdX4PKO4+OUqHpqXkBFGlvCUQ4E/mgQ1e3QN
rez9132vtgtYyLhFU/hHdmKwySiZTPZhWcYy60kPM6QGJChTwjGnQwS/WosujNRyn1+jnbh8FHd/
lS1eVZ26nwsUirQDyURZRnyVFy1yJYYyeeYheVgnKx4vLrPoaT+p5ZEdgog9K/s+XuMQt6aG0rSD
HPld4JzUOK+lVcilOWWDNVLdM2ZfzWMdyiFGSgJLPD+Nx62+bZykyC7bFbss2qePdvyV4Yvu3k/B
5vcBX7JT596AuRJ2bGK8KrcsrDHEp699Q7LVB2uoqR/HvjqaN0Fh0DnxmbHuJKPIuMwAnLdvWMWz
PQtjMU/9OziSg+RG/tbBTjquIrSkz571vMHmAtDqgfwop3q7ZBFThToGuwVB2QsXpgrCmjBMky7R
42HapAOhSVx38jUFJyn/eQJ56rxAzXw5TwwJedSPtmMZF6cbXmOMSuG5BEMvQib9qVsdd4iqdNdh
JqACGSfJwj4yiYQQBrE3FitAMi2Wsrz+opyiUxzh4Br3yZZNqoIjeVaNDBiJwU0k57NuakfddHLJ
kncLqw+tUYaZ39zMRIhEMof2UkMHhorF4RJJQUvCCw0F6T+TDPh/NiIRV8lZPWPR5LbfVFYHo6zJ
zkNXmT8c9r3bap3i9kCMQDC9OmbjFyVKjdrrF25nuUWsZNuFs8jCtsKoRu2xrzAWODEYc8jqGx8z
enKcyiqdJ7UC0fIX7AAZXF2PDnVKq+GAYLxIdH+txp0lfpQuQMkAswPFDO2VFGlcERmARwHiIwIa
PIsPj769LnmBFNWAIS8a69viBXmL4LuKpEJMUv83fQBct/hTD+LywLcrL0X8DbIEBYc3DIEc4k2B
j7T3wsioowhw+kXHyJRJPcVOz92x37Xhy+8vZbBfIWsyHJe7jLS/NZwK682HGnKoH+rVzN4l4o8o
56SND9xCyzk4evoLLknjoexU+aGRURlfQ9yOjq9FsKkGCpmKg9a6MH8/v8kYhbmN3rx4OaJqQJib
CGiOCVXVFTGsUQwuGVDeS3fu3J7P8Gyn8MudG4svVEh/s50jkcpS9iTH3isbOD/loMC7/A3S4QOk
TH3KLUeN8isWwlHVbdMmt3mFmjRuAWPnO4987SWZTrIPPx6v2miL8ZjuoBBbExeW3rwjKO6ynMUq
EyB0ZINz1kS6YaQcdNuOSn8985LGI1aUv/0dNSWc3F1amsTr+uxnaMqRz5VJ/VSY2bz2pvljJui+
8mbsKyq+ZMyauLlvmjG8OK7HFRkdvi+Hm3X2xDfcq+VmPDUnHYgf+abV4w4BD0INe8v72zR7SeTS
HJsBO4qIw3GUKaKdxSHHAJkztLKFzTCRYPGYQrNfp5hwoFE70qFQ8VZp3vtZS9SWydlm7megWXli
8QSNgw4hbvRbzpRzIBpu22L2dH3ZxeEHf1RxHyzZh/3Z3dUdXLByxIjqwJexAjkwDIcp6t3Uyjnf
fwTMSj/Z55ZMXxJWtg0kpyuEtzWq5mmifPC805WWReT5Z47YtqPQX0wnH06LMvviP12ldWAuMnqA
NJEY3ctlyORNj6kyOaUvNfTP13V4hC47k+CpVQBYPO6TEVLoQISwCav8ZaR/QSQw1mC4Jzkco0VB
gBuXu9lyoRuzknijxnRU+nQwpeTNiVHfpQcP10VLiOppqrUo/hGVjyCzSzBLQQWCpykxt9UNGdEk
hD1LrMrOZCxdZaEJooPtLqrY4aG2qfQuKw8i5grLzEUQryU2QjH4IXf89z7yN3nnx5hTo9+t1M+f
iDwDyHUN3CgZ5M57qctlzU8aEC+C1mHt2CjJbrc9dutoOYLbwJSw1i82s0AFIxku2CA6TYKdMyWd
f6UHFlQGpZ9wcVoU0RFKSaINm3jMJmauoTjgchXXdmy8sOOtnGkM6VsNwFjkMWlwENtnMlVBRCrB
JDZkl2kp6j1qijopEr5PliaRKTlkzpzPjCcOQ2E03ciHCmZQ5dmqGPaFiH857/F+gvDrGiTucd3X
W6Z7NYnvsXX3NKHkt4Gm7NSzhy4gcG21gux7WBEQ7n17Yy8/UdmKOHy0P0XoAIvEVxUetSwCy544
aJbQGvYcgP5rxx9dumswmfMllDD/U1s3UZKLQVMb/Ljx1rzBokc2olHAbwVttKczm8safd/inqy2
MHiiyLRtu2OLU3DHOV1vzlw527ZBDWVx03rE8cNpnxnGh2eGGo2/8lp+xRwaNF+yrp949BI54eDm
xViuasqg81AtFyFr5PNk68tGYrTBE43rbTqPtFUrUAaVv0kdMcfK8u8MIAwLmTMjVWGE/vWLUbkB
xt7Ng6T4FTB2TpB3cEoxCn6nc+ujSt9ocBo/ENhxTtHFkCMFOiMjwxSJ5ZmJdKDVrKdOD65+ouRn
E8j/sSkVxIg4yYAEA7xhjBohg0wk1Fc1qG8cEkm4ZiHqiowVYE0OD4GdlMAnXXTcsj8oqjVTg2gm
weY6JISQYmY6oJoOhUVW69Qq+5UlgvffhjYeTnkDNLmnxZIwqctXCIURfsvUZ8XaE0g72HlVnc4B
J4qTFjbfZ+cSI5GnNoaptvv1UiTJgtp2nb2n5zn6ZZs7sVMWBXSjxD0L8Ne7j4Zj3LLvcK/CVlEO
1GPLDeUj7bXjBT6UT+VbYjLROWnWR04ZVTJ4+VcxvnaOjHe6+l3Ksb68tRmooWDUeEzdO8MTpE2e
Ssp3Iwb3X9quNJ+I7FKbb0zaosIha/z4Q0t1vll8gNWEjbZgzy07whcgqyWThDW/zXwmJKTSdlzT
zkJLCiYwaC5iHm5/3u4zjf9WAyvyoX7j4y9D6uB93PFBt7B1dynO5ywVIXP3Z9861t5TKGgyrmQY
Lr/84vsSNtsWtAiRwFU2QH3LdOnp0PE7veHjP5Xekb3HT1IvkGUmLJwU3dRg7argNDzfnRIycwBt
JzZFRqBLSMFgSRhxQCuIQUYkE4turKSW10zkYf3J071L4aRnkvo7fTaQ3sCtKGOLgyTZlq6tBQw3
l2+edtP9GpTY68uf/yGLMpprCSJbUx++qQuM9bv6MHfaVT43yFPQwnnRYuVASzvXGOOQvlNdRA9/
q8SwtpCHy3YafTi6frN9VV976BtyqGRq4BdMA+xF7yW4eoD+j/kCp1579gVAhUv0dA/j/J0KkqiH
WMS1p3isfvW95OGHslPRLoY+f94LVRkFUFcXUOcfs/5y175uz+j/uIk3H6CTHgQRpWNmuNpQyGLY
4XhZIkkMqkw3DS5W2fupMJzwTE5Ad78j84BOr2n5gEzR/cS3kMpqS84g2E0DXN8v7PSCBufnm0Wu
Qh0Xjzw74+E7ue2VvDu0Nf+Vq9ngmXUQl/I0gB1r9/BPb2H3cxDKS8UAQp7mVZPeZKPKvXmo7tUv
S2Ab1RGbZJX7EMI1NKmkSHzb2joBQTsuQSdhUwTCPRTr/2u0JcNHhfKC0NpcQmhOx9+YMkuFXwXi
zEQHTZNKT9lqWOGQHSGjXj+PBAlB9uYOIqbK0egyLZk+a1cCMyuNNpT7B52mJ4QA+UJT67RoX2Sh
SJhNyXnzvDqK6BJO+Dp/5Qnn5Lq9NK2b9x7OVOrF4XCJxNUnhVkw6gwPxN9ChgS25vXdePnl2Pst
EoBWLTybPQ4jjjOoVnMTw1Fr55K4IQX0JMqKRjEuFdPgGFz8cuLIdg5KDl7c3hsVquMcIjaxIq2i
8QuG5czLbupyxxGz3oQDb++U6waM58LlXaaEfq1S5AjZSIkPp7y+ILwnzdo7yb5wLfVOXZ1KBddr
68TtL8x+8me9M12dk3gXtxiBKZJNLw0UnL2apiYKOxCnpuPsQd4oyj2oOy48sUw4Lfp/mm+B67rc
4DEI71Au+nc1AeygY0dqLoyiLxVJYH9hOpTYPFl7P3LVXv+/rmDcvyYWH0S6deF0G/ZSzctdBrGb
l2lp1qPJ8vYNAfhraKSrIhScQ6dacKtNYUiv+mSqPmyxf1PKkBreLTcersJZmm/criw3pAKJ/ink
74FsenZhMN6lT2Za4V2kraJNZC5Ss9EnCRn7k/kB1aDfM0cJ4Gv7z8fvW2r9+mmz7iQemJpCKOWa
mom4FAdq8eJz8yoebYCgKetinP5lXRCf8e3Qse0faewvJDPWAWILrRc1J4HXMB0NKceWLZIufdao
U2+61GHIauKpWPkffQDjy6/h/rlemURfUhgsVYEbW4kpgpcNovkIPYJd/DgbcmkA2ffmHoZSgM9r
rdPb87RNNAts/kVv6RGBJcoSHXtiUfYXZhjPSm3VIksLlDlAo5zdJENIXT7iPSmXFjOaaB320VRW
wflvinDYtu343fvhqrUI4X6XE7Omvtlqxc+gulyU02MwpexeIFZak9ux6awtM4KdEX0fZH+fV0z/
cG/axtIBoc6/pFRfeI4cVpl/lKIJaE9WuyaKIvXUbYOTjPzCy7nMroEcAtYnNHUAPVboIL4PGf2Q
jk7CeC89/3JWCoFgEoiy2s2k7lNFv69XoFZj6zhwXe7Cg4ZMtETX8S0cUtaNSuBFDEEgxdJkxFMf
6CxvbEbYV+ta4KtUct3JpLRduSAtW6iNGajznEuQSf7yhjIOdzUk4pogCx83xwPV4M2TT7cGhFb5
J8qTC3+CllAMHcG1/no8s1jS9mnYo7+IdZgq+bfkvDKcgZnJBgfQoc3UopksmKq7Fq/DOxAKI3Zr
4+TUnK5wmsKTFA7mbC+x18adzNgeKMQyV6yB0a5cMVodIlNQh01nIoiCTb9pjIkAZNcrK0o2X6zv
O3Ph6+nNbnKHCBVu1WSgyl2rw/1s+1Yp5MhZooeL0u3EV0lg4Apj8B46mtqtd/tD4PqN95n8JlzK
pTAmOa/n8xmuiw48E4dP42iktDtmOLOa5ijtGjh/fvZ+uHUGGTSvH9/uM/+oGAE18Oxj9tEXfLmy
tUc/u/Glmq9k/Itf/GtoJWJ6ksiWPJIfXe9hOM3SIzQl3f+rTbFc32833HMFegVrx0qs9X45rV5u
sM9U/3WWtNyxig+q8QQ13+s7V3N+l/dKdauD8OaU1+yFAV2RdY8HaJS5cm2dfEurXkYjkWk+Cza7
xyHEzGgb+3d9/ubqJ3JMsg1cUsiQR/vwDFofGli9Tm0Z1bHLbz91UUhzwpROnrjJ7Db9Ddw9t+OL
kuGtYanGQuG/L3p3jCKKcFtet6fU0PMfQ+dj0r9HhS4WT1Z2sGfFT0n4a6dTNR79WCIa52eROZn3
CWq5QhZ8MagQOrjAXg1D5AEzxHbzaM//QaTXHOi7oeORPa7Ijz7N3Vb88wG32RbZRV1TlWFvcitt
m5HShHrhR0RPqOo+R3OGEdLq8LnYHMLi12aSiv1F3njAv6UpJ0yM3vZsf0JyJQFnglsla4kSDY7V
oVjYEX4olTa5w/lCmooWz6/X+4ArYgQsLWn1GEFyEnnZWJD31tOy08yHrZKSdkgPUV8rZPcQzN2d
f0UP0Wca8UIBq7AbuXGNgSypha1pv/T3naEVwN4qbfFXcf67K6N6p1XMB8NpxKMNM/5VhgAHDVQg
R/t9sx/56ZduJx/eVZdG5+tvlgkcqBpGbJWcmGLGr+VHk3mYea2m99ZQ8u/FyjIpEhsNQejwMU0b
yIiJdvl7nh7UCryAkg9dUYk5193bHB+l5WiDoy2GC+uch9OCGscFBVthxwYVCbHAwoGpV3FlD7X+
pPatjUmicRUNC+4LF+rYO36lNMQ7d4R53MUsAT1RkG06diJQyLGjcOlsPD60Ml9n4IZwXrVcSqcV
i1zOtJDj1K8nbimc2Ij0/5Qm8yucqWKP5AE0S/OdIET1xrcNfhN13YzE4b/V0i/YivMZxvdtz/tA
JjDIyy14U0XNkq+gwZKDQZ9dLuvDz1o1CQFWLoDCf3+U2MuDIqokdYKn++usPYZYhLHnCmBWpGyK
pInYGHAwWEpQ+vacKPwObeO4H1uerXZsTqLy0q8GMtjvUvmJeloenhxxVu7zloie5k/TRRDMI1vx
DK+DycnVLRn8YpRQoW/zPdeGfYfjCX958bQ69WJ0V2bxo0ED+7B83+BBEPnJSz57pO3mD6WVVmK8
WjenTTYi4pnyvQ45tUuOPRL+106qALCELXb2TftJFBm27w+Qb0Owd0STR+RtqK3Scdkhkt39tnSO
kjQ1y0Fz3LS0JvJxmeRg2Xr4G2iJrs4pA7q1XVB3yMcrL10lbR7bjC7ZuSovgnMSuxzNCBBqzlI1
ynJPGjvyGx6F4gUpN0MiWx3INGCSrCUby/udB8OCgPaRkQsgmRiMfkpNYCYvBpiThZtJuZY7f5Ns
HQSAMpBXqbVDDVMuBp+bLYTgxHbhP3t38nquSuf9zvwfpDmjODoUzZowyQx+bgX1PEUGfAAx7dKF
yZUltjOs9rT+mIFKzob3Bo9hXa8ipuo4i2guKTRKvH3UIcbf2TW/8jjykN5T+nQUiTe3Mykh8U9Q
TEANLLOQd/X2SN9w7O/DOVGizm9RPG8gAivIsD6XozS4SmrVwekZxYmPkXG5usRv8ga90mG9kckf
AV86aBuY55YJjLsmAr9i9k7lfafHtyTD+GmGG7dVVVyPjG5eF+y9gOQ/tDfut/P30M6D0K9DGCnm
Ji2b8IpJF2mi81yvAN3/znaJ1e63k83S7sa4Xhxa1vCC4U7X12UdK2rzCFMpHd+M3nIr+j7c6ERz
uwxNqewN99ltnHMvPuHQwO31enhsbPgZ42pwVoN/zMbSVJSoE4uM+HP9bDSYQs8p1ckAhNdAtwfV
gzdaqDUUPpjvHxhpnOOF/IDXGEkFVZQKVpfCSH30vGFwn8TQtrrpxwHy9oKQ5LBv2sg/my7zEdVj
35IYxOI03lMKVfuAlKpt1cAetizpX9dbaiI9UVL5c3LR1UtkN1Z01Vf+NuB6uR4AjOYCD6kLlVjB
K3xwDAZx3bIEg8W+Pc58lW6xk2Yb/S0GU4CcHoXsd6fSuU7ExX0ZFJpaAUzd8ob85BkEB8w8eocr
PCzqyKj/ijoCdpmak9pH0j1hmsXWH+5yKpSRRezvitqIq9b3c/Xvqh/sUGTr06Gq1SRP24TZwmqx
FdVtkbtLBqkP8bPJsx4d1+jwNhv5Yw4RajUPPA4SL6S9ovglgJCd13+SCojlQMxERPMHalsDRCzZ
IMGwpCihIkWFDWwXQ106UkIItBF+KvMcGXRxY2C+Osp3KQdAXLzvUSbjeCmqr79OAKvYgL8zfhuc
DmwQtqWi5r/Mi56vmCKtQFc5c5T+6wWhLm7qS6EhpifqIvChDLBlfrxKp2NVUucYbnZ00ubHvy3d
4zTikt3j0T3dEtP+2AdmASxBT9W5nrvoSj5mF7/oW5wjpQuuvd346k8IzzeVrz38wKSsgunkGZci
gHsHppvSRJeNxwBD932Q5+TPPOisN2IEkN85EIlQk6TlA4ta7nzNf0fiWl80IKQEhj9PZFmxmja2
aeGWgquWpUU/ZdedV0LuBMaSHFyZl3GB/SHwjBMCXvx1idl8MeuUdFakuSOku/e7qrDIBkAiQE+X
poH4MK0hq4Qj6MveK1R9suejYJdpAlTwNt9WndVWB6b+23krxTbZZhw1tcxs1TnlRAEZaL6Xp7nh
78vGOEQIC+k/BuVu4pZ5R2T0789aOHcGgvfxGf3Rw/6sSekieERLaXbH4b2G/zZpoZ+agcRdLgkB
s4Nmlm2kjujwaqyT1DRlbjd6Uuscha86wV8hdFEqmoDWSCEu6LbMRn3M5Gug1UvEOLnWaRueHuXX
8w/2n9iguh2fbayH4/aaWA8UoSTDSSCqtYvU8MIEzRYKyxl5RjccxFEDYdxsrnhsZomVEMcPF32E
4D3inaZP9m4Od9IfrBiiBLwq58mx1jaCve5VKx0lL0qM362no1HA0gNyFFpihCSvDcGtWEDEm/Hq
hHGKONxYd619Nt7lAvH/TMmECpod2CyZ/Wjmjdtyita+Q8sXIagsjuK/O6aLi9xQmoYsKXK83D+T
7JKyad4fSQFwMOD5M92F4LapRsWG0PttxWJ+1ZqKwQMa3+58jUqK2rSZxbqtjQI0lAgNaDaqZeK+
5OJd58ttAl5pjB6oGExnfyKDUhLL6mnY/0nMbrD9gFXvgKZj8oxosUKNSchu2i3SrprUN+6OY5yd
gzVarBfUKPSQb4WsLq7ledFJnKq/H+BfQlIKkYL78Dpky27hFaUrDQNWVGytisctO2jVVXKcxDrg
uSQu26uX3RasUVeKRlXEkv+5nBhd6eSV1OiALb7BqHutnW+QH92cl2NPjusD0wGH0oRbExScznf0
R25IT7hIyv+HAUxYaoIdns4Rxt8D60ZpGjt8qAcGMRTDVCsyDz4x0UgIqTBXfXXMfyeXEcsyK5IF
0OJLz9APy1Kst7AkwT/9ByWm4k8QNN+xVXLPktkNwSHw2DnYxzYuI3jsaUOUzCH33xFzA2z+8urP
C2VpKkkGQYW2kdItFvgg2wSvFrfLrld9OINdDLtGD6Ok0p5az5Gmk1nWPsfC0IWvw0Y27tVJkEsT
KXlPls0G/MMTKS7ge07HYWfq5+eWmY4SYrRqNe5sjPAZK1KH61C+rrwlndKgrA9V3wjnlNjTY/+F
6HhzxXkiKO2nL3Mxf1NBtXOuTCJqWO5G6MMzV92txYP8gk8GpCkj209yCvZNhGUBml9RAXPrfB5T
t7WFFA/cUerNUtGn1LDXXT40wqjL/Hl1vre3i6KrSSSgbS74Vd+OtVDnWBL+5mu9mJoSYa7RVfkD
BZsEM2Wby/rEgXov7CPmD4HHL4aSidGxFibPXO6seY7K2/DoUJfjKix0mbIwSsDM+aA6uF4BIM2W
JAegPvTjboCjyxiab7WSX3js1SHNytP5Yotm0x343f2SCxdTgCe+aOZC43UhwcQf0EmndzYE0sS0
ZaGNmiG3n4DNS20I+BRQ8yvkwrkMmc1t7x4NPL3jbzG4IJCcjcjCSx5kutf/xzxv78sdIBqPAK/K
RrsVHUPHgRPi3ghQvMQ+PmYYPzQlLyytEks8nthmYwMw/Zgddrwq6q+7dLbhP7u0P6gtK3Lla6KG
tXx8MGWRs/oFJn91Haql6ulxRN/jMUHc8WK18oOsHkJP3n/FOn6+/apQZDTgTshd6/upIUxU8Egl
sBgtEMwDlW6i8qAFnrj11uATBsT/KN4QA7EbXfCHKKx+O9jfBtHTqMfku/2nqHruHkTr7KZR1Esq
d8U4XZPy8d4JhOXqWNImGRX+2H2260uJd/3vmmtDSNZOZuV5h+nRHuJpRiPcFhEpSOnH0nIs67FP
1Q2I/yO5J4TQPioByrxe5VObgzwmgMxK15z+QlddwzI/ePZrV4va+n8ZTgkMsnSS83D59rsfIKsT
FAjva/pzjcIEp6m3ZQegWLOsVV8lzti5F9YZOXtsxp0/13erA9KQcrfPYYmpIAya9/zy2dxCAAvF
CJBhc8hDllFMp/ANiLdxnZCkStoxZfqYTl6wF+563RjyPTZ+Xr8vJ8MwYy3kMVUMrbPK1vXGWw4z
rZl7HOTjMPzuOKWeyYqvEW6ov+fduqdZCEpVGPSCmOmwBNU8dDq9wRmRlpyL9wPE2dzZWPf9b1+W
qWcc7Pp7XZJ3lGhWSkv8U6QRMCennxnVuNuQKkcYNIu6TevDB2+B1rzNpP4T6eBfs8Can1ExS5ht
ieO3z0e8wkEGf5mdo/o6N5SZwFBzr96pTg1axmyS5k6q7Bpomv//GtsCHtcf5cWZWE70Ho8azHGS
wNRtVJIJxe/as1tVq8kPrIUmOjqlY1CVGm2RZN4/S9/8nvCToHFE3nvlJ5YrGMqYz9syCJz3y7Ii
zB8PYRf056VajxbdTCaStr0FSgtSdnQjvxM0scpeKLSdSp+Se2VYFgWu1s16X2YWzF+Du14vWM3h
TUIueIkxhkweUDb1f/zW9O10QGPeycrV16d4aeEWX82q19pJ8giacSj9RDHe84OTZdhBbJQ1kllr
ndAj4YxWE1sPb7AN1tuJzBAC4vQUl30xuxFziI6PEE/TDJkH+q5ZYUXI0ExTa6A/BoL1jfQag0S6
PCdyOxgRLkJWTm5aoJDuKBSrv8pgYipzIQWgTH/a2kwB7j7y0pI0P1HdimnRJTsqqAvvkpNZgTv+
arsL/MQ54KF7HYetapheuW4pGzujNYXDAtMNMuz4lro7gqpnbm8qiln/iT9yEOsDSh1KZurqhE0z
YHWpZRKulnXMtNdrjrMoXG7b5uxODh+Z2fIjXQKarX9BNEvyKIAFBRj2zT5hwPL8YpZONGD0j/ER
zxOk44rTdm+YgefuLytdaUcFPY66faxjbGjyGK/wL3N3+yAas4kIFIgr3sRK3K0KD1oYiyo3dbsp
0aoO1dJS4K7kCivl3i2OkOOTWu+MjjavdapF+mJ6TX1ACaA3hO+OkGflh8cAfz2JDpgJdNv21LpL
uhpucKrfh4QiQa0h4bWzEOPn0izc2s7GM7BGGB+cUzdvnU9SFH/yme7nimSjvPEIBv0wWBMlLskh
5XV8Jk8+5az4pavUpGQS8PNINVjoXsQTy2XW/0y6ZbMI7Yf1bfhV2HisySob1qwGPXyIBYDc94vt
S4PbMpn8w3El7lJVtouBQzriYXKVUKXpkkkbmDKYWTkHCXjhKIHRQSFf/ClrrJROvmPsvEkXNysp
2CZCTprudmp+y6XhjlVtVaAZAj5TwqgdoFHmCzMEZSxyAmd1McCPyvVVjcmydrFHRCKzG0dowwjA
Cq1viBn0qfip5bNjsXvDFJ93YXrFKq+2xyvW8Sb/lJRyV5UQXasPTjsP9uNTvJofZ2Y2DC6yrne2
ZLpxokyOGAzAL23xcKbwBS3cM8BWZipnoJlLwaP3CMsBDmVNsbgAFYQqgVUj5euphmdrsvga1ghr
nm29zTfwkQSs3bxQUWw6bV+ls8t3PaZ43kWHzzwS+PdK6fmiEKH9++ckGYWFdWj1tWphwNcTIX+g
Encb3YGyzSH7Wqrsyu77tSKdH8FFvJ0ySUMIzZvvVmKuZ8nMHwp2tl8Ep5JBdISFfp+dNbPs76LE
pGzq1ifcCV3pp0lkFyQUhNJx1vf9SO1M4fr6bMrYPZJqaxj1h6K3jaYMcogYKf1ZinDHk/AWlhgG
a5W1VfnlGxtaDCk7uroRJk2xoNLXWnVqzgz9oOxbIg7mEN+ObTxJ1HUNLok7UF8GBGu43RXOSCx/
R0c6iSIK1RaKp8BsNfnQhEB0uHSSuuQTEsfhNLR5EryJ3u45V0dWfACSPP2LOG3fc7j+8mtvRh/j
zjsj67sItqxtm2yKZty3R2/aBd3v4iRhaCqw/u6VZl9i+W6kFbD7WqcZh2AzSDhAO/wPaVJsOXOM
uXSPtUZrpOlAeyjuzZpoIr3VFKP7S8MtBi+ALFH42ryF8kr6LgB9+8m4xm1FfKvpw8VDgx0d6QzK
fU3PPQ5Q5tv/vdwz8uw5fFAZVaXb3G+WQu2Js6/P6MiWPb8QD8CZHSSwxPOstw/MMECJXxzDePHN
lnYdytReIUhu7x1xpUNRmLO6bjaucv1mYk46Y2Xf5VuGXt/h3J3A/0w6MuRc/aBsDoXcEzzhDgyq
uI5BitZYNijeSRFxxJvwYkjAK/G5Rb3AolScCqzsYeMezmAIue9NrGnoD2c+Z45ty27wemMKrFdv
S3XobfAdMX3mgefdDIhBLxgGk1G0h39w40N1eanvRz/JXTc9HmA+nfqQpxXc4Kp+3Bo5VSTpIkaD
0ANNA+305Y+2g+DLR84YGltQ48bE0+Tsu1nkMPl27NwWA+5nxpzNXDqL3IMOwlUp2JxPVylfJXJ0
0Sl7p62q5I9mATU5Yrscaq1ODRT4qlicL5j3fEjROu+tWXPkgzTqlSdknQ0lEM2Z1NppmKquvteA
8hxH0aFRa+xSgMN0qwJPEwR57F3dMSkyO03eyXiSX67YTD4nVSTskneMNpZ77+Npr8BoXrXQITue
Kd0zVSGeCj49b2g49Tm0f3q1RiXFZ47FjjJEHpo3S8CuDbwCv1E58fMFLKzggYGWeB/d7aiOiXig
RzFrNjsEz3pJIFG7E0n5cLwD5b8PkSuz0UTtx2ScLHhgXDREVKxsO80BFWIxJiXh74cSnRFejBo0
hs25z47PQlV5UGOkMo67enq7JL9vPViEPBU2TEqiNf8ioZiogYEU7QEIqIwzqvXyRZ/3r47ar2TL
MnfeXebBkPqUpyo+44T+GRCBjo8rDoHWRtCu38DFqpXc0MSpybPE9qbcKgKLDxa+Ras6a0Z9TeQj
TXu9dlUCVc0LjFI42WpUhYYfXbjUndkCh4tjWLDyRapni8u8XwwxSvD677iNAbbHgZfegOMHcPzs
CtUwQa9qnYjSGTWNAPsDqUEzrHhE0CJ1AXKtyh/5rFecfmKfQ6z2loSe9NxYfg8Nz5P/ntFKtuWf
Hg+OGFhD9BMiyByqa+hz+sv4lur075jmc/LMRQByD24+g70hFhzwqHOPsTp0VDQnymrc8+XjPn6F
jlAFBO0P9ulJPaRh3NyFWcmal4Qbz0dpbxtKIABwrhFw0VLeyxNKeR527QJ51osBbq6peLRh0rWY
sbJ6l1DwDuUj/Zo5ZawvNCdje7bt4hwNt3zu8qXwISqRPeubp9OUNzlNnfd2a8Tjl6lbXYjsXUQC
aURtw3CnJItUTME9cAICHAe+jcLathVrwK0UwFOau7nUt1ewR/yiJqhAAwuhUmWSZShIYq6sEU/H
miW6Fdob97yZBBOBWeLwyJpNtmwRLkvNZ87Id/2JcHhfeUaIlDWiTpu2rNgCpfoCd5op7cqeHTvZ
4Dzmj8kgGw4e+YUrxJ1qiLuqEm8Rk2xwYUMM4Xag0V8vlKQbjJ9DfEsGuzexBhuuju7xfnxj6NUP
cVKmclLJeqpscmLLK8nsdJ5/gaF66rHnhPmf37mWhs7P3/+y+KqBGqcIUFfXDrJ69ZIU36quF5Oo
3TC03FFNAnqO1jecguO/VIL0fh3Mbwg6baNKQfn12rFVafJKcJQqT2LUWidZWhWS69GiWuEgPx9u
RRPYCCKNu45+8Ah9u1j76cQO8CNUuIK06Dos0qUPJYuq4PWKoXvlRIKdFuSvciotiMqNcUbumxeq
0sbvCKB7Fx6Yl31R0aNji+lD5qnGxwU73YC3QbqT5yCF/GfuT9WkpHd+IHuDIRdpxsSmTIEgpRDU
pd3Q+OgqcwZpoGsiDOUs2JPkZ0XjgmECUY1yUO4lorGH8jDgKbgviKo6LO/qYQyYaBeScJYcxw0g
e4MVanYZX3WCuV8cTfbkjHGCi6xpwXJZC62xv8mrR0hOFQlzb/4tgz8DLuI2yZd+BZzd49jCOTxN
iNIWhSBmJIZZAdGhi/uk7ltwNkOnpqhX7r4CkJeLOHcZmjFmTQzUot4xYe7+iqqImZqcxPWK06eN
5+5vf16OAASFY/6KhrshCGwwkrea2pBtkMP68CY1iof83zacQGzx5Ymcr/Bm4iE5WI2Nz3JkVL/7
uHRJQU3ea6wU2Ptd+KUDSuNDh20HQUrInz/6uVEZoaTZjZDvvO0MQP2T7Di7BtIhJM8ZcR9KO60r
8KeCnrO8GSdaoUoWI1hxpWnDuvqwgjdDrswn3dvhlSVLTVGsehOn9Y3go+N0TxURtRnfcthjAl0R
BAhCRoIJRLB52rIs5Bv96RrSD5mWO3/hEW2gfcxVmM2ROyYK3ngJmUwYz2S+NO7pSARcQCx8G39/
gX0M/gb5JO3R6Tkyk8NDfX9+hipkfaCO+PQnhDQeuxZCVHXXrELnPXX0PsTHYRw/bDdSDCgefyFx
tdWLSr0P8rQWiXbsb/otl+O6F5HvzUrIK9KGxD1ouT+ZJGjp1yPwHYMXVbgZ4AiiCmNUePNoC1Rd
g01ru7z6yTAIIm1yXHn7DKHQnbF6f5KhqsFQKLcFcNScBYU+5LgoVruiXMW9iuJJuIPVTZDvvtNc
yEYXOao2hg1OMxGIz6z3159Fw9811gb4TpL4U0wERUYb9+EvlTzweNhfGiGf1mEOP+7al7tzxe37
P631SaATOUNXqB4/uWpU4Ge0UzMNhpZjJdl17EE+t+YZ2u8REMexe8JwdCjIKsbUYBYfHVA/vWnP
qpqVSfa7OUHvW153ZT0EGbcf8A8A6UxE3kipo6Wjt+IYm3X5yzHJqtpdMgFIp+PAxyoydDkGcI3w
/CwWLXVBJDf9i+4iBjEnZJhgrxUb0b+BwaQjFGde75GkpVt2vsxV1jwQ9FQ6NdDWX2sAnYnWYiPn
vLWKxg1wN0deeCgK/R5hEv2Akgc3C8RUwIp2SzIVxmli5vOKU+KqB4VyYj+9VLluMxCuCucuF6iy
wZbWBV3DBc9yfc+yoPwHjq970Ywh/W+/F7pMBSyIm4oi5hAsIZaUFekQtQH09CRGjTqSWPyELhi7
2g3J09Ybqag0dw0Rmd0lsIG5BmBKG0TruQF42i7e7f53BE/V1iZyy476abq3eqZUGHro5JoYJBYE
LFVDqp0E3BdnqPUxjutMJ2Xy0KZdB/p5F02QxmLaPEH/ITUdp+w7cvhtO9FlTZaS+qt3pirTmPOS
xm6Wsj2Y1Fp+lq5N3tRUvCUXlF3y3gMdKEcs0wmNtDCO3BsA9SQbrJ9UiZxAWZfjV+KJiT3izoQ4
4ye0MWJSIi7L0ALngY/kStyjJYxbch5lYGtFxNivWB+WdEpkLSuTCqClVp7/ujoXAeNGsgSIgtxt
XGVPi4gd/R4mZ5ZP8zRcqbSpvoLmQ5PdDk+hz08W03po3gEMQS1r4lRahs37m+nkP41Dm1QkoW9g
O0nLjrYSdjfq80JnNObc8mblAicw7mQU5gR72z+K4obYzK9NhiKNjRdOm0r9Ec0jKRSZQuQ+WfAW
ta63aT7p8lkArGpRVKyPuJyjRlCr4y87dyYjE1XMph23QfB3XcujzwVxs+CUzqCPZUyc54DS+BEq
tbgHQ02mk0mbHJEBrWLrx1MRFyP7LAKLVYxLO1dCIJqieeT5OzxSKrRAcQX02Q+/n2RAw4OCtm2h
GpM5TOOWAcTDw63Vmtw0F1lD5ivLbEMQTvE1A1+811D9i3xy9SPebqBndYVK7+y2V8z2eo9b/vl+
M4ZWddmjq/9UNcglRVCVBoAayza8a86+zfgSMqFtM5PepVIOzPoV8ZkcSHNYab7M3c7hn63BhH5f
IV/5ynJz1zg4R5H2eJjGlOpw0WuE3AyPNmm5qIN3/fFmfJVxTvr9G4MuvfZBEj11ZedIOSO5EbNc
5dGxlnubouRwhp935n8IaZAnTDJJsHQ6eqaH5cbxeq3iwVmsYKyhyxks9C7qn2R1QwO/4Y6vzc15
kfC30x9tkPikrtPLGB07S43N+Wyr1oAkis/gsIoqsHIpvmaQt9OqM/LLjY7Rdtarr5yc5eDOnt/Y
v+uxVbMBPG5y+JKQ5PwS1+ZNFApKCrKwFqdkNCRZDgBGTKVYZA5xmQslt6mJUnBDEiLAEh5g/R8d
z6v1eQuLIhMpcynV3SuAFiSYXI5atnKhEJBj9t0o/LkpLMp7ZigxirfI8Ar0nAzSFV+Rm16Wawd9
biLC8fOX/eoa+LXJwfh9oTErOaITOtLURChEeGrvh/RPOHuQZyBXEy+/sCjaXIjkPF6KmjKR/pyf
8gFPFJABUBqvQ6N9KYRW0Ye/Rp1mbQIwZWqTnBpnKfrizVSBcRN0F3bvGy0gialpnmFGBtZuNiN7
lcaiVH7tsYnOdqR2yoCum09y+i6PGcNxZsR0g2GlDiQ4INP8IhSJkyzbC9NYdQEuFI6K4aiLZ+bR
fYFlXs8rAX2h22hog4dCbYj4OI2lQaFL4iI9jjtqaXOejPtcJMbDgDpOFFhYgwBMoQtuID9YRxie
SXjxjTFqI3GxhXhDhJmehi8ofDo9+ntK3JHeumTKovbZBixw3kOv2G2HvDHmm8qCK2qfM1Zcp2gh
0ewjZT4TQqN4mTgZln8+T8ZZbOYL/gN8oRtVY+2Q3nsLE7dhfhagh8QO5PlXt+epetxV/9jF9j3m
HvVHMtt5OeHn67ExmVzKPqs/JE6qccdS54X3B/Ibq7906KNyU1zYijQp9dJF3JY1AnefgevVuU9K
ZHcWnp9ixCP/Z0y6ZoqFOuyJP3J5C7llsFm4Qth7xxZbBMMnlgG3rhyci6VqA9nd0sxDfQ2zh+aJ
fI8gxxL1eULKIWrNO/AiMuQXk7E/1ezDnizzwfqm8BAokk4yzv5kQ7cj029kVsNPkwwmS154sVXT
bHh4d/NyTQo7JvmlY5uFbIqWZDEOyFNhi9YzJreOMrVqitrNrKrZFhrVe4+nOhdT0fB5RTWBrCcO
Zzt17r30z5irCfeFhpcOjri7ExZMaXKN6MsoCmkY1oeTXCXC+CZ5PKzJ9Tvh7xWZhS2sBl9rUtGA
Re295FCtOhLO5WkdgYukSEGPcEt8x8sHfgsAi7Nl3YC6T6gzUSDgl1NZB22qPuLUq0RjfpUYvphI
1mMHqcrbR8IzOnungYyIrvdskoASixmFVkD8tvTpmhswDeLKmCf30yW5/075g+sH6N0KGj8d3k6/
XPKBVfdeKtBYa3vMN9rIBawQ/XnRghGHK2Cb97qsjTNQPq+s2RT8/CV/+Y/0tnUp6l0xnD6Sodz4
ynoCuB8usUR+FkI+9scuuJM8LfGmq+lCUOrPwc4qVfoK0zbVf6fFwl6aGZ0fb+2igff0j3fTRsjO
2yWv5zPBaJmhMFNi2+iLwISCS03+OhmbNAjPEk041h33bg5PZ8sVzO3cFk57NWJd8DPKYpS1/EMB
GTRLTKUU3GsF0slfAhl3Vgjr2Imn2WG+6Bi8Z0Pux6STf9m74CYUH+GkYYVNlfxv2TnCePHYzPF5
SuxtWvBkXwfBbzHL2IT3J4PSmqGMcpHNq1I8T5x0oi4CBYVA3nFIfnJFQe3aLgV5Of2wlnQgIxeF
dcWn0vLl+x8mqnzF/yK+VKCkjrD2QCfa5SC6Sl5wLVl7KPHC4OOTh9T4tl3e0IUaagytso6YUl6e
dCUOJXKonqGAhZr3UO3UycdFJp2T/CjRZNFkZI/VZS2AULO8vKpPlLe1JkjVu27VK5spro7HuA15
4OqdgZ6SGd/Q5sdI0qT4jZKWjALFKdLryax2tXWHflXqDU5wuOFnOinCI/hU9o0oXO59iMgs0PkF
8jtXMem5jcble2G4+B/+R5uUMB5XVpPxwrzwkuTmSJY2Sa8E8/NJTR+KW49UCPd++yONLM4jaFT5
gJYV3sZTiHekO/Q3nIneVubpgFYRqfpALjiQ5geGJweqZq0QW3FsH8M2jAN+nMLRv2ixSsSkQdEt
tqX/VaL4nnZos2r4yEbNakh8AWw3ahoHjkUT5my482c2/MLzW36sZrBr0vX6NnRomi6+SkCP0Nda
AAQIERBkT7gAhAThWCXR+S3u2KmEuStamc3o4dcUzp+6qSsXJloCUKI55pzrn6c5M9AUKUXDTZIF
yYROfSySe9jUDUDuqbii/ouzBgIj53oyjyTDNmyVKql5Bsv+BAMQgPwOnv+U9UU3llR6dxVeBlVi
x5WEUgo7P0/7Ql88l2ElWaHcLlEaQmQ85E92KgTxoQjxrKqHf9R6Fmcf6ZFdp2FXGzb7Yjsx0uT0
yJ590dnKXKxhbC7HD4VZCulnaG033wzIN8Qs5Ce32yEXdpoW/pm+GB4mgLucObY5KCYQwjXPQnr3
2S01+ZqZqJvdmM2xi+J1NW391ElLbqUcIBN5y0whTwiJxHwuE1F0JoxxAydRUapIZs+uwKvSo3A2
Mcs7wMn/xyvRU/k4ccCnC9Z29QNwU1pyeNWUBSnld9yIvdiLBIzNZKm1djtJDjVy562GiZSyPs4i
Mc3eloRVRf2zyIXg2ThhSMwpFJZhr+U9Q2GGHY3Vc+e9MiCtf+Hh2wWRdyD9XVatO72VyoX70tih
SXB3sd2G75mvdX7OORhRJM0akrsPgekxBcl6VlsGGmWpK8hY72Ft2hedLcY64cVPlNSDqQZGjWPt
G7LsTgeqS99vTLpi3tN6bmblnSnUYhGmSAvChSU0Q/95tzhVpUxDgDBKkvGbJxazKJCi+b9RDATt
i9RqQtVe5f7MgR+sDrBUT52gHFNrrInOGYPCGwzZUOviEvhdYIhNjKJIRCRfDXOCde/mBOWFFh4E
B8VExd//JyD8EyRE4Y+e6LG6Bz0OhAh4V7ymv07jmiu6GTOiAhUqLoQasbxelgstVmepjrf/3+Gp
gTktJnav4uudKo6ymyr/MuRVcqO0MMVOQnSHvms7y8VFUjB3JSvNamDsnMmO324Yi7EYazc2akrY
z26pGfYclCKkIFOxlaQvW1zuIe+dGdBfXm5Ej+sOJ6ejw9WJADdp38zuWdaiBECrUN/g09G5ljFb
zM2PyDmRaYJIVURuVlcz1YkTU+u7AYnuOjP/ClB4J51z+5zOpfciRyC2KoB45lhQhwXtLNJTCEAn
o78tyNiCO1Wt1L0Bzn44l4LPTqyDh+QBZFEsG5nwN4OdXJVJ1RH1/c/D9AkXV5lGRHH4Qfp3aQnM
CBmXCPEgxej0EX0ti7cv4K8GDSt76vKQhiLdkb3rM/IE7xjFrxNKmw0XG33OwoV6TDlKvhZXquA3
6LhQxian7Zytsf8No+79Bow4SQ1Cat1NdoRnMj5afB05JgKNnIek++lYPXLYNte+ohIejDfNod3E
Z4Z2ufwufiDx3Z8r7bItbHxUZ3wKz0sPmrH9hPwlu7lVZUgbSbjpFOiKUUGyFRe179UuVLF8V5m6
LQ2N1n8u25aMT/2MyN82riZfZQZxkWl/nEl1tg39O3nD0XPq9mxXRXrrNCHnX/AAB+LqTKXpmlUl
mJpjDHLtcM+gRF/W5f7WNndKxxOh0j5zcts7KqkqkPJ/GR0sXLGG1SHTd9yxHHbHKqZn/LfcqZF2
I7xnUJqoStIGZsnOJrgo/LbjeVYN5PkBzUfi2pLvAfRXZqk5PVwTmbBABoNOtiujtsbxU46ODHCe
c+W3MK/dSzkj4Umifzp4Le3wdnBefExQoSArTlo+gKe93/hCV1jb4EHoEECUSNvJFqWCoiRHHjSG
/MUDVYBwtqx8PHlwdCc787sIMV2ZIf5Ga5E4F1cDI3kowNlBPVl8qFJTCAT0Bli5mXvfZGvK9Khk
FjSbkQ0vWwmm7DThWONqDbd9Kwbtp7xvC3RYh162Vs/uuyGpaA+25r90xYXqy21YicSiH+GrC/KE
Qy4IxBHE2MWxlWjqus79raxTwIgvqUgLJfX5zy+LyeH4Xr7k49PfBTeC+vZsNnqML1asCRzVvMxW
AKyu3WD8i2Y64ophuy1gthyAuHFcSzwsmpDV1kPyg0i2fAnydbyD1oEMnvkQmyPVz+6QBYqDLWJu
YrWx9t/v3x0Iaf9oy3LsXfNcmVFtfWUxbYQFibwXRAGcdl7Ul8owSk8nlw+8X2KL4aDbpc3DKtvg
oSGpISWrgTAb1VE8G1BFDV22eDuSMT/ItAubn9Hwqv6l2w7q/coy9MoF3++0qjucq5Tf+kMY0fhe
nv1uqGHFwDtPPx+noXIikK385mAwK2EEE1j4yfwqHBMOKrvqIOJYXh2gffDu5STHc+Ra7wb30Gnf
xykHd84EOaWyZiQz4fY98UyvYPui1O65Di7IeVXnXfKfe5rTToM0kmg3AnfH5dzg/i0E2npxQGGs
D2omwhoq/DAQzeU7sKMYdZRCK5wu+a2AiQ/HAXonPsXXoSn+yR3do+0KdI/hWS5cbg7VbOBRDBUx
wLnnnpekkrTeToIQWrqoOpjhdU8+gUkIEBCPEPAKz6hLhYnpUDA9pin6TsXYN50q0KOW6bh5PYs6
HMK2qWC+zZLjisQD3cPKyV80M2HmSep2s3B8d8T8h2Z1bJVAJV2evlOKqQVaon1D2XuzPQBCLBDE
0QBpFTjlc1PRPub054rwF4k14ApjxSTWOwQigncClLq2fpmTfjpHkudVXhQhZSc3SOsdv/TSCu63
oqV0m1dRwlh+zo6Jvu90e0PfLvE5odGAQrj0vr0gA7F3oRRVw85z4l6oIKC9B6JaYV7aeNihHqY2
uuc0DLgUg51MYLjvOGJy4h0zlwE1bgReRSKBt5bgPmOlODyub5ql/V6goHdhJTgftbI1WnRq1BmD
7be0wrk2+fNYdrZWs7UkPcRqF0uCc67O5cesvN0VgmgUWeMa5vc/Du+Ivy6wriMLGP8wxk6ggGSl
1vnHqThDmoU8v/sASchTB4zRZIRjdNDp/DlP/oTiq3AHXblOJP5zozlmv50LkXrzhdbxkNR9ytja
HRZ1m1RjdRogmEkIz0gvpvJwBPBP9a4j1v6NELCqq+cNckkWB39R++9VR48itVdxcgegqM3JABO4
Cywx0jkbr6QkjDip4wiHy2M4tyfnMT3CtFHXGZRkZaDSJ73vVzaDDl4QyNPBBlndkTRLupJCTuZE
uJHBY7yiblZDzF1BMy9JsLLlTYjFRRve3jAzznnvpGj1oUfpJicreflhFVm2EdLnE8jEZXbnHAvZ
lHkyrs4VcKFS8NT8qUhOf1s+NUm5zUsVFz4wb6vL4yMnO8O56DG8X+1/tGDDWqdHOgnn5oz5RL88
XM2+YlpVO2NLs43E5mS2L61YNbDqZ3I+oArsXZ27rVZxC0Sbf5/8iZ7jsJOVrfCAUe8RrMf51WQe
trEsviEMbIm+meNg60HYiBtv+KTHaIR0x+8zXVMXB6P/Ka3kK1S8XY1xvwIpxg3OEt808FLRSsbS
RsQpXB/zX0eeRtCJrmNL0y2TeEOiapXBSYtU87JvMxT39eDtq76U3IioGN3VZ/mrgceZeV/7pYKd
W+HUEighIq56xy5gCFOfy+XIhm+knQo/axgLbRYCvDCMlxpSU8Rce33wTrVO4vAx8kiFC423IELN
sDITr8mHgcgv2gzb8reBZsxIKB8G4HkN4gCH8gCd9FkZIMwlDE5i+1/TZJsqnVWSGkLckfj+Fi8C
p8DLG3Ly1p+p3CBmXvd01sg7MN7mMrH/JhOD/FBCzmr1G4tokB2u41cFrGoJ4Kpxzi+AWpvaVeiG
o0f8qaoJxZECJFJu37DkJG6bOAGiNFNHJs9dGCd1gWfPnerZ9Z+iaVYBKANP20kF9zhKtsrlE8zn
riei3BuFMCowY6fHe8RVGX+ZQyxEDpmoahUxgH7a+Pv4SSIidvVAedcvkZwAZYpXn0TZO/RA/9hJ
AphxKYTILIvl0/2Zctq7zqkeSEKtTbk9d0uRzWyfISaHFF3wowJ0+1mtKL5klVty7uqVRUhU8cDO
a0FAiEsBcsqUBNwq6SgNVMEOIm2p6zLWsc/UMMYHTLt3DjOICSkYZD73tHmy8i6eJEuh0mmeZLxV
zpGBbhTpXkOCIh+NDReoNFX1EqwpzvsSlELMAGfZvD2UEhi6yMrCwKjZcchZRQKe/ePjnrc57ov2
nvkGG9Pd05DGJuLM/TR34zvn+9RekidZ04nArgKP4Iz9QQIcnapYQe8unerJer1U1Ci+ibvGCuqB
IZU0GJx3nCKHabDiVnBLHsAVEsUhdBNXq2jUrvkV6+XSWkBIk87sYoEpsxl9OKVF2T413M1WLmNx
tvvzJE2HDJKdiCtqiEDCRPoJwOR1YlWdnl4lwt1jq8B5kuFGku0SUss3c8cY8Kwa0WHLqB8tf3hH
UMyfiUMBqgk8ZtUeoGu7Z+Gq5aND2pgZRw3+gjETqt9UcX7/5DwlwO8s7FxMnwa3ntEc/1Oqhaxn
4Ln0j5SHS2AiJhpOcObt7KgOUABscGVNOGQ6VPs6LGoH5TX+q44WdO9Bzjl/Gz5rJgmp4bn583Ui
QD7xgltGLNhESECi6MZF9uF1fcXN6yAwiIT3n21vEt+7uvtmzTGXy1YOCgfFOGethepAjU1AELyC
R2LgxayYzA2APNqN3E0gy48E6plu33UrFePFmamTf5rOM0VAPe1Mcp+lkD5lTjEezRmVKFVaLanB
JYQZH7QyorAoIlLfl+MOVRGpPCpe/K2myDCFgvz0M9YJ0XB3X/CYNGkSG6u3oHhvUoICC8tz+ysT
jSZLeycFSiIYpd9KdDwFBUDH+k8LF0opndNbM1P4WPzrUlbPcO0zk7kU4haO8raAakm896pQLX9w
VAUuohtGILoFE6Rz5ugEScg2t2DLqduxoU+zfWtekEc4Q1BbfrSHvrLcnHqMtVRu10qux5xj1B9o
Aoi2EL5plgjhq7r9N9Fml0BaRFEUxyrhpzAASa1jFE5oukDt0kfuYwOXTui8JDNFDQMtUCXIvr2H
d65pqfEpGcLux2QYTf3hg7STpMLOPHNDyjDg6+BnDyA5pSzFmLQaWTixtoK5wbvyfh0LBBd5jlgM
gtaGdgm3IDPncvXuWtN2rPdzJsEPciM3nfoE5cqZgqE0LPOmOFVzYrWC31LyxSREaGQDPC8N870L
QB4ydQ8ofot8Gy6tlGkc/WNTRTn+zJz35lNTCzSpAcfqFdASXoPyJZ51fUdEgw==
`protect end_protected
