`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
qpyA0WijCXtjo0xVnUu7sDlPt5Jzg1uPL/sta785mYz57etTJd7nREGsKylYFpGqK9dUSDcuLQY0
2TbNQRUYtlQT9fMCzlc7uVbMARyAvHTnm5WGqYbI43fDq9ysz27YwHL7dzJ/cMWWaNf6tA7i9190
zzzlwbuXCnmBhXELwGnPeNJlkA4S9xaRXpqG+7bwhSTa2yUr4K5c2NvtpxJ3ARYSqiDCxg5zqI0R
hCg+ejBqvXfiNax9LQyGTjqsx/6aPSLsnn9a91bvioFh2yt/zTzBA39F4tCX34pKF33LASP8ZJNV
lLfK50x8YAaIqaYNd049JxJG5zD9xXtoyT2uvg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="gxdR9PDc/5qT5r7I2sskUwKpu99mZl5l5i7RXdAmU+Y="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`protect data_block
EXXXIV/u2xcXBWiIjiK648t/ZreHZn67eeDjc0kiJjZehYozEKD5y+e9qag+BRjUmSwObukqpdte
xaZuaEoIQrdFqMI0gEp2Q6rs+5YIgSckzCMY4SLLynM/3ahxWEi8sWDKjClD1zAI720VV2cYclQ7
7hD94AN8yWM34UrvZWORIMmH9iQB5UW4IcHuHwuZ3R6dj7lijsblGaevg93Q/0s55tIR3/cEExcx
yQlWfvN8veWxrlHECTWkI4iWiqvDswFKLSim6WHzaNHZ6vW/ZPRV361sp+WOVjbwxU6PVGTC1vsy
AKztCg5pO7Tj7OaUmjVMDhEB+TI36MgzbsQITnjZbnLqzbImljB2nHb2n8WIZt95XqvrkQrt/tLI
wVbmP+SbRZQGF21rNwoANJLZKjYPfYjv2qULogci0veeB3YMCJBtZqrDjqwPaj4byLhSueZkxHdB
VMSzsYRzp+8+9A+4tEOZfCNjjIa8NfgODhunE4m7QiJH5fgJpehRVKkgFjudFNBCbBjnZq2+cwya
n4QSM5I2r078V2AsREQ5ebpHUavvoI83fv5ZKMOT3dgi/SGwB7LAok+cTGZutPf8l/6bTOso0CEO
O+pn7NjPIfPQb5zMBkMaJnAAPbsL2UqE8ZtaDqy+9aWYXPV8Ex8Dah9afQ2O5Yc9yZvaXUTXksT1
ECpascTVhWUG4GnQbmumMGBGL/9pBtkk9vxf9xCqUyJGY6JczwwrhET7+N5lU02A8XFAijWxoV3R
bStHraTjlT4xcKteBItdjq/9fK8qtbcdgmgIn64D1kDJj7IQJ6kMZXe3OPcbPcI7VBTmNdNQGSRQ
D9x8Q1mFEVFqO80A9wzF4NlA2LulDlEALErdna2ZCFSfOU6/wu/2RQCj40yHPX37YRQ8ZXPEqOED
KuRe7ybhY32MQyL5wc3OhiFizHU1+J3F3LsGNL/GjUe7g7T3Hg0aKqEe9xtSww1ILiayWrv1Sc5v
IMfPLZC5G/pqqF/1hGq9MUIKOmTtCcvCrIhMP/NCJasgqs46ZeA+/S2noOurrbDOcHwvUmP3Idjb
dqlCDUdQ2zWVZWMHto2bqlX9IRfr8LFUbc/s2YFGk6f/kfmEB/+gRkpI9jHPNVW4NUSkNjFCEDpW
husvkKt+JUR7elmyz9hnW/l3pTSH6UywsOC82pG3sc/kfXgf695kgPNScJ7CmyPj1MX9s4jaklM0
Ji+cVy4kwO350lxVLB4jajDAHGvvU79AyEWajoKAAu1QwD0DnyFJrxurp2V2po4rBANJWKlcp/Uw
zdPZVeF00cuHRZ8Poovxwdkb8zwaPlCfopRm/onl4Ys2JI8FqtwosOw4DFxrLamzWDU52oLOWXKM
RFBNctBnrtMwO5ngaNugtFj+ch4SFVC393uXSwHIGIyFFQ2vpQzrekPsThf1j/JjgTMYgTHZ/6gl
RFjYGTe//IWaGxFqlURSk0bnlA+dfWIZeRawLh65KYFj6/kE/KNE8CjU2rAIC1uCw+NcgY5p+TMd
YOR23uTaxWhvJn/EwfzwmEoaqc4p3sF8SlP6gmfFFX8N1BK1cLzztaaJiWgvyIii1xz1zovVh2rS
7kRuZTdXPkM0AU0yUrKV7mP++yg1tsMRmIG4WDjNNfW60woa6V51uFgTsPWhyBzn9Jsn2qbj1G47
hKhaF+aZedrYTYfageY5W91p2xfloLAefR9QYb8HxJK1XaB2tmPcHT3xkuXpB6Hnn2IPWIxm7dBq
jz8BkA75H3PJGJVP52NNeo/HRiqCAregk87QVMOUc/FjmiYDY3tjobifGo5eyN3hA/1TTqIfW0lt
6xYVUAShUCuWmtiZkytaTqaiE5icQqaHfVLZltXjJIT572pFqiNKt0Q1TjzbfvKFFIaNGJCWWVU0
tekCmMMcjwjYCYh2WYjGIaD8LyGqJ0r1+Rc+Tsv7TwF1uUTUVNk6vV4docj4876E50+YoxeNKPFC
jW4gZKOUqlsp2j9GlCrl30OXSsh7qOAXBNa+Ktrn9+ptC0rtk6e5YlxkXMc8DgH6kdvoH4xB98Ut
iixOqKkHcuIfW16eNhsXJg4Gligubzj0V1+g9NKXhd2lH4OnFPdvnWYf1if9WlNof3lYm5ot3Y68
8BZO4LnYgMad5qeGetOs/8+AhzMWRt3MwTK32Mo/Js9Du+CClnIacJU11cA2R9X1IcGPK57UqMTe
C0FBUuyyir//6bqhu2d1ZCRWo+sA9xuibBiQyUKmoUNHIvMt0KMx99+0pmueDGrdPWiJb1nnEVQ8
NP5+Ah9JYqZduy3nxq7RM4qHKwgzt+r1AvvrQ90msNQTa74s10wY2chTnrW4NBH1s95x4A+fARLS
zhsXc6nCV6M2bDF1PQq108jRhNX5XCVYN1nEYPqxdYx8mN82MO68M5ZaabERoIvzfeUZMC45G9zu
DC8aCw7C6M5og7ATDXOuqRwn/8JOps626DhpVov1mOR1FxWi1L3kbo9RnxE1wFd5UAlSfB9j3jXy
B8hdKPhOI6FkgfOw7ultHkfV/Nu8CuzAq4HEy6xQhryO7Cp8vNcV7iNQ9ohUCjGkSPT9B7d4zi0U
HxIUskOlVz2WAcTYgQONnaNhJFN76lSKr5mW+kVDRk/WqiyzQXTfzzCAul5hfmsElS9Lfinx9re0
wDcbg2BX/OHm0hek6BsS/BGOcvkCm+qzMQrqzcJehIti+NvcUOfZ1xiOJnVWPdIkFNBUKxFHZ0vO
13lZsSJkd1p+WANxiGClPeEBE8tkfYsNP51kZEBKSethSO3a8p8Z/1J29KsvUW9JZ1JKFCy5E2Pd
6LOFX0Az96HVaMBGymdNt2b+GYHcXXSaBUtAFHy+4lSRJ2xlU7K8qphM3GShzC/BSrfOSETGd5UG
McStx1fwRj53ZR6hG50PsUR8sIwNyOoEuuATE/dv5VJ5GH9jvD3AizXN4ZfbFDbFGPRrChnD0g97
+KRD8zAiP6RNK1tyBHvhiKeRltNa1BIxtGkSeTd0S0mQIHXyRQHqqcq/cYEbwKCUE/DRWQMT7Ah4
czwdrzij57BQO0N+m9YBL2Fucy8Xm3Bu55sNFVeobhDZjMNfkM3AkXJJFAPEadWUSYvQjrp7xchP
jb3RqrEFmUjcezRn9MdMmJjqwuGhvkkSxymlRVRBkJLFfV441489P5OaqvCZSJlr2+gIDQAccGOq
7n+BrQ1KRLy4kzpoCAGAoQSVmyfG3L2F2+VKrGJBvTRgJynKhJPehDFRIOAEUDVyFRHNcC2cOnSh
JU+dcqeTBwZLyWqq3mbHlirMaJxPLAbM3tNZuVlT6EIyfu51pNmhMjp5J42WIisYQJZ6elrnN8Di
O28z5Ei0b3sDS14daIQ4ou1jVVsAEeGpHs554bUwO3DxlUDwZ9ahvgc03pt39iMX3jSydiJa5XcQ
aPHV53XSCgp+l9TA2Bmsz0VYL0QLKGSGU8kS3bIzueNt+hV6jwmAPRXvKyRHwa8p0+2cK+15eR3T
ZafgpbNCu2GnW9OanTpBjIPBncXuX6eS42hfiP1T0I/CPRIJGQfd7f9S6ca75nc0pF82XgG5lcIE
Jpz5GQZQr4b8Gk3TS/CGnAGSBKYWqxCGit2KEf4mQ1w5tG8hagxRMqBhVH/oedoV5w6XDv5MZ1t2
ze8Qyg8AGQ5WnvcyX8b4Uu8MN4Y3B0xx5MgM+4uPQBQj1rbQUpktQvqPDWq2E9YYK/z/H6m/Qcuh
V7AuAagrtmMEUVRBlP88sejrhRcd52XnJSLQgDLqE9EFslHkKNvBEKxXdFZw7qUQ7qbrPblFyDc1
pZmO6cNu/2AildT7h73jPNCLPi5mNIOKAxNpumnujz1odu7SGlcACLJlky6TfE20g207Qk99aTE5
G7xCH0NUWfEFekCjesRvGXDEdIm0dz/A2I6o+AW2sHr5+vjofAPpLPGr73emEA7W87dOcMV/AJzJ
6r4Dv/xzYpYWZlNasl6Q9Zwu7TQcOK//rvHSv318d2egLmCl7Y6oGZCvlMYFmfFoTawQInpNKl3E
6YJ4KDAvyQUouElEk18ezQvwBXtBio1Fq1qiS59QhL7zO+xyx7LZS3O2eW067j6+KAB6lUp8CiAP
EwKNjyLR4JdudrzTiZs4WRvpDulONmcl+hx0d5J4MIWwzQIDv4HVhCSnmeGgbexJESHIunyMJGwp
GRTjGCLvpJs2Zis4Sxemee3pBTmfqjKmzI1jLaZC4znXmFI9LBh/hNYQGcRPToNC8y04tLJJ9gVO
NqpVSxArPqu2OiTIFe5cTxtxEIGjzCJ9aYKz0GSgYph3SX9E4PdwFEetbPc7eSYJuztyVUEr6SHR
SjxUcVTCcg/H9ueiP/7kLcAIP0coPK4aulFlkXEGJ7Rh+ieEF+8dtTMER7kZc4BvwA51458lKunN
7sM2gzaXMcmd2A61W61Ie/0XZjG1ZDC/NXbHWQ1OIodCeerAbmAxuglouWKjQuw4DXT4mjWndNJT
bIphTns0SaZxZAEfEh6gfn2ghNzTOKBGm/ncjz5BwGcOZZzP8fhUTmmo3J/cL2aRtJm688CnON03
jDn9LaPWgwD0XXbNjzoM2Ouvhm1ksyBZU5raAf9YNxAmThVDqlZb4v3mOZCFGMfzOJveaCI38k96
91doy8M5YcP8DgXavfrzRPpz2WEHcC+o7oxr
`protect end_protected
