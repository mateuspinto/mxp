`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
b6AMGK+56pTs8FCPbWtTGsUaOwUQIOvM/cvEBKSMJmlLXBu+YFm+Oc8H/wgqxf2WfszC8uYzXCQ7
TBBG04oFN79kGjO9ViDs3R2JSV+0ctgs7ORokWm4SGi6ln8S38xihGqKL6NSIdikqBNzWc1DNwUR
K1faRt6gXtTltFxWXRqqG1psmHZttgUDoYeQoYRnsagN+YZpNzcSVTUjDoAlPc51uidTdVhBY0vi
mnwEr8kS+5ZeyXZ9JheKYNBQHFr305e4PMoBkam4e60UAeRujxizBiso0C5y0NjXVL1QE0zEFDxy
qaIATSVA0FlL9xCOebYhF1D3J4StqcfudUojAA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="s8TPRoNY8RPjGngqtep7/M0pJquIVVLqmZUV5F7mVRw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13856)
`protect data_block
SKucDbRyU4qLQS4UScujd1F8cmkoiVXmugEUF6RWb5suY0JT6xNQYLhWmNkdziPY7kDolnGo8kbd
lXz9iZZjQPpX6ZAI86vUiOi/CUCkZa//s845FSeMywpQ/Z/49NpcpUo4nZBBjy/DQU/ggbHwvJuX
AtcDTfuxDT94GJ7VlmaIjX7KPWRoMgV/id6RoSQt/F50380B8/fVVLPUpQHazoRyMb2PDKn1/LsG
EPO0HBYEtj71eCxsKKMGdBlx7hX/xAqdHpdmgg30AE/sUt4FRml+ZR+jZggoEaPvE3hADeCl04GX
ySLaAzCIm0t/p8m5UZHmh9xQmQEgm1akGau7xAJQR8IYg/EEpvZl3wZnk6Teq4TjacxOJNB+0k8p
8e4LkD4Qe4w4FkWxnZqc2p6zoA7U8KFID0zcGNiNEKLf+9sW55h9KIEpkzUvTlUvTcG2ELwRuJIN
2B86RoqhWJe4uwgpwteYgD5jTgFJ+4Cfe8nj1HetrCZQKJxdSSHeYCu3jPbgOAUO7pUg8Ras+IEp
kiSjuQ/u7n3y3luRI1yv7umRebgcQ2GT9DJc9RDxTkJSYViXS6m7V+Wu+1opAF2qfAkYZkUXQ8jr
o52GvMoBLjsL30sL2Ll5ceO2R5ScZhb1v0sv8VCw/BD98qm4dmWR/bLZXpu0TJbwfYgYI4EDXfBY
0kLBtIA8iduDygsZbPxQjudFvAQLdaHqvUX70sIo0dZdS2b0WNewYYIuhWhKBOij/Myu9rxI5hEt
V8hSBPS2mDaGMtH5F6IeES47V9VWMkC0vQFEtZ5RNTAickc/Og7Clf68YlsuRD32mNxVrE8B6dZ/
fyxTaQuUyZ2sS57QDDVtqt+/QkfDaFlNYsliI3JVmqp3Dg02PaS5BqJdmQiErodBAvhF39NAzvum
GIZTLy0FKuBSiaGVIDMKFD9LYilKK9trHMdkbjTGNDC+VGqmj7ovJNwlvHoW7+hYznowVuiKC3eI
+DKtxGFghPahew5zFbHAwCYPoEsqHoToi3t82qvBumBsIBMYbj4fPw5xVLGGfn90CZAEUxsHD/uz
ZbSlcA5uNB/M3ELFkDaUm+ScU112eKYM0wVIPmTkpxQKaWdzJfwiWk2GaPbTCrmoeI8DQhbXglx0
24pWwVyfbfjCD3N4TD94eTf0eSRPXMnQmHCtAvffMlpqjuk+JvbkNq90UZ3Jd0VnMLeM1x4k5arq
gOHWnwUhc8zJuMU8QDM4v9IpNfOk5M1dTMRNNLRL3coPDTcCuKhCIyYWmI7EUP17bR23cIBdZN+2
w41DOqgCZ3catH2MqjV4dFsNPieU3d9/LnslV3BikwybUY73pMz1/yy+182Ln/EOYON3VnhD49QZ
a/OlKcl/ceQRAkWqfkgPmqUj3j+EcZxJ1Jj7j7Mcr1WuZtQK0zH+PK1n5ksxm5WD19KXi02g06d1
ggTPt8WKQSTvReynqc534STyNdnEwDUfYUAwGDZL7EdOTWDv1/MD7Qv7OsbSkhVuKfNTCRSTkFOe
70xeh5Nl0OxWcMeGR6/IrupnMQJgXVL663Dbea6FbPSMZTIL91CQwKgQfk9OqIXItRzlW7nAhvjr
XP+ObQ+izhsvPOrRu2jHYsP6+Ssg537kwC4orlzBtuBlKjBrs84pNNE80DOWhGzZKfKeM2BsPAzZ
VdUKRz6s5vkJKBqrtjV1uufAXEn/uhGU39vRSOK/5LPAdQupOD7LBc2kzMvMTI2/8bbQfPhIPpxV
OEqBo0S7Ni0IqIiL8V2sqITnxyTmFxr2L3/Q5GvNp9TC+leh5I9Mw+ElbmOW++Ve87ZnOPrlPkDw
pmIYO52eyVbIvxEKd/cNItmwtvOfXXYBwgtHwpjSGML8isGLNzxNYP8qh6HMPFDqmXG98OCQMmOO
92rbMO37b6g81GKXz27ME54YxoVi+wOQpjzI6PikF2Opa2afKKtMPgE7TuD6SbdwTXnx5p6YPPJk
qBMDQjM111tsSGs7kJOL02BpFMsUGenCo0lahuUKfY+oziQ2z8epWxxTKyvFA2Nz3l7vg3qTyPmn
z45J5URP/QAAR15F8bg3X8USseQ4jU7zj1CHIWpQFt/7DruN6zyisQycSTSvk5xhYaghAwlW6Q55
fqvkoKmVD4l5sBGTveDytIrdlHRUKX1pc60GTqc6pGqyXck7/8b9L6hdL2qxGfZwVMOs7ISZlD8K
sEkd0WSoJRszF8RWfsWCpBwI7KssWAUyfwgX/jIK48KbC64tW1HrJ5OwGzVx8g52zQzlN3rsor9g
CYw6mC9C8uZFHdFxiVg6WsO9zTLxuZqCajHChzj62Eo4q9ZQv2FbOhKYSwrtgba5O8iiJZO4c4di
7PXR+uLJMywzHwOQ98wvn6ksCG8fsA4bZ1BQs/nrtuNMJbrSgeVOY9g1m5t4m9V55jG5uWETtU4P
SOXk3xMJn4d2j4EOXCBTyKdTqQYIrly86j3Q3X8LHk7kKX6NcGzKD2mYnoq1AooOeZ+vznpt2Vq+
6n+inUbtO1Cb238f+5B7CMWcluziYMd02A70hDJvkEWFyZAVS8VTKpniveBtwSNZ5uWWm+cirBsr
bE+EOSp1m1dHO1mYQXu6kcvSL49rAnmCaaQF8B1GBKUsQYqHTHu1FXehmZEl6m+wP6Ek8x8zfK7T
RbbrjNacQ6uqLX9PNabWMckW4uvbIAZ4LKIXYpLAugR1d8AQJpVEZxcMz5VW1MxOw51EkFerp9Xr
ZR1B2MurzsTFSkogTJ6/tci63zyhCETYc7ZQAhCaE/V8dP0pu12s2T7m4C5JgOdHuhvktKziLPNT
ruXICnMLG6g69D8/xBe5P5mKwAGX12FhTpzlAMfwcTtk/ohGiI9KcaF8az4FkCRlqZTk1WHIsUil
B7523SwbbqJTzjHBO3ZsRY5YrG+PITEymmvOEtVHYzSKPcmrj9peMNBWNAU3OlPM8BMeKD414cql
ivk5ceRApksCQEAYu909//YBEvpa2D6pKeQsqLgrqAAv/6Ofe8ps9OBJ84ya/RgL5PxfoCL4atwl
kuMYLARi1BAJE1fObVarzqsjUbPErmSh2O+KihhNsunFmvvNmoFzWN7OMC5P4ZUDDvfQbxFo9Zui
vJ2aUS06qndAmPi5DhrWudiQgpNgxY/aIR2Y7p0Yho5qmVC08RJzrpipqJ/C/12TWRjWqKwLmGju
tjOG5k7sDq6z4ITXafAPWPoQFRgv5I1NdGY/SEw/4naAEscVyN23Bo5K9+ZhIiQrOi0iibnOTwCN
xA3Li+DEoGZsv/S9j3mSlvVn4fJOgJunMCMZ2+J03mlW2EfaczL3xkdBY/y7K6bDgLJrFYiy2jW+
hs/KhUAvjMkRxTLFHSW+5UbydmXKFOzN4mqPIPRXZ4raY/JCnRbj0aMM17VkVkhZkJW2pDbtHFA4
Id6zCnERODFjV0V07naCQ33SzrFZpg+b2N4Dbzo3By0dJxF3mNH+FsOczUmQZu/urelEeTO/0Xkk
PJiSQsZo6EEZRzPoabe6YJMqyeANVoVgGbgkfTIyhL958Gk4zz2WLcOC81akMVIDTWoSesiGZ1Gt
hyraB6AEBqcqmdHfgdlHhUa+/e7hYhqqlaffzWDUYJjZzwEf8UL6WdYCS+9EiO/Ryu5LTm000wrT
XQ/0sxO4s8K09vT/fRLCVSCCZYFOuIAtCWEaTFVxhgWUoEhMelcMxKasL6YuDoBqdjfQRETjEMk6
kOQOv0alo56M8KACSuHby2F8m7829NUe3cc5hU477t53R4Su/NGHh84qHDlxIs/VuSY1VLrueIr1
dvAwUObMF2a5aso9Dps1Flv1SocH0xprrniFR5CU5XM2Fd3AHtDRPFAQVVl9xxmNzgt89mcoTGEE
fm2Z2s8wnpgzgmUF+HhQhOPNebo/cUif3Wyb5v24ZKHsXhghhj60hqZ6VHb577KTAWOQCMbW8Rlz
Xse1xD8t6YRsykdZc8rJD+nW1UGFQe2uBLtGqKxIt+XI2WpaU86O3hf7k9iZSqLxrF3b9+jPGtrX
bCI27B/YQ5OZh8uUOOPkIanf8QJyPdf5mJaNZ2e4S5MGplKvn2p72KMUSeDBQWbN9KCEl9vDoZ94
0+yYIBcSQFuQ6OeEbsV3cDrX4x4NncXUTpi6qsatTZXM7/OJnAHp4HtLFliJL4LyyMFsRLIFCQZN
hN/Qfk8RilxXI/9ygFeJsIQQA8jSHtjywQRLQBRCIfaQ6VWrhBlKKlNZ8paYTs8OlncdKjmNMqpM
uk7lEwIGtGwoI4CzV0h14HHSguZlSRJ18c+tYGUdqnau64Ocvu8OYq2ta/1lHrAIHjLY7QF9bmKB
cd25t0eyYzt4f1O3vxCnsLzW17nSTX07mTUQJUakyFZ6UwpGdLkIQKhKoY/2Mtcb1mvidAxQwMz+
O3CDPdPZaQXbgvBrlALyQxtWtawaQH7epqHWtzFETFUDJRVoq42aPWfUxxQyaWSfhoVRioLh/bnt
xIBrsHG6INIQlpdL6wJLQXmKfYJ/8HOe+ZcWkoAG6nUCw83ulNBbrMuP6s8wU/oa2esg+x0KInn0
aqsp3SYH31GGl8+AFOzU3HDlIvlVM0OFGCACPAR45m6F1yMuOfgmpfn0wg1iNQ9ZaCDftHQwbtYU
Z2oPierneMMrMiG1nZ3EFs0HXmR7OZVzjqu/vVtt0v2J/ttVDX+TkZVAo4/gGjMHUMfNcxRIeMxw
P4TnDVbQmL/NAM/jqDyxXuKVODkSP8MyURUUcNYo0v7emNqu9YUGD7FsJlO6gioI6azQbAhpEWIS
zpWxWFMpiUTVLJIlhKjd4sXcDSbchmgzZq6CCS61tVnzX0jHxD8YuCV8LngqcMl71b/srUntSrp2
ckZtXKrMsd10dH85YgJGL5X6nVM7Pz7h3qurahN666h4Ewm1o5N8zBk2hjxndnQr5RMfKcfGFxNs
pGF4nW3u4mQbaCe9s0u4ATshJELjl8qKVaoOBC3qYbS8z52xAsjpS5tjNReA29zuTxiS7pxRpem2
f26YNEAUThR1po/dpFF+UYVBkunWCfQBP/yXMWDqXg1DkLSAQsgV/luQFvUTnkCGUOQJsUJmNNYj
ioci2Gmk4MfPcdovSaAK7h6n4sXblraUYUMdCv9Zk2ZpVwYr9QKZA6OYTMSUpbM1GZvjBhRhBgnI
1eChBouzw9ONMvn4BXMHpQo3LNf3CEfTGyL8+Ehj19uzxsTAkSJ6GE8ilRdHw+YwUdNbDiG4LAr1
lgSUkkkegPLURoHjry4x2iGHv6MmuHF0Bhg66R75otdqGZHFFaBwQEdExFe428bi4/6uU6kNFUHm
cHa86NSWYwp/cpIRUuOfEJezVCjc1yP1aDcSfaeWQqxKkEdXubuZAyoc5rvb4Z+7WUTvQK4ibVJJ
xJTEZ+6UazHFrS51dKGbyYRstaaxKhfcZX2JNZqJH7lqF0R1GKe+maJk9YnOWAxhks9v/763tC/C
SYYBTDWxCVogfr3sxCKAANP/Pj4KauhEmGmTD3Ma/QVWpy61iDuTiwnfv0L/sykVYuzKgr78Z+8c
9ZiZdoA89ZKh4IPMY1beJfixnutHCdC0s43JszQPJX3k5jBmXMUQnMBY6y1ucLx40tEYiQkvnmM+
Md8f+hmiE53NtkjBth2JelcKPTwes5gQ8vpqxW0iJXQVMvE8p2EQDWdwqWmQwSwfD9CPB87zagVh
4w1KRjfVAA5Y3O6mEUvI1G+blHgdaqvX3jcpS6E85PlKCEoyABFQpDBPdbTi7J1ZvSAL7MzHZsiL
b5pND+wqJrvwP3ICVQwvsDRhjX/JKUEp0+ryqG7QurwHEJhKC1BYE5USPlUqca5VYPjVaZER7lMh
d4gJ0THukWTp+jMLwWHVQ1nwEnglA/+0kw/qoQ1itSBKaeGE0uqqhCSVD5XLm+1ZzXhul02j4JKG
lj/5p5ttFskiRqd6vcwbk9+5J05XIHIqredMdPNaKHfQ3szrGGbBgBFzauN7tMc4Hb783sJIkAVe
3ZLpX5MiiThd24ewiFJRV0ldDbPGi50U6hwIRe+y0t3cpG0LdcIR/MqKagWyFGcBpMQQezBZnG+J
tD5fRJFI8hIdpARx+J8RvpNJgC6+7N5PgEcge37Hw57e5Lf9LcvyGgloSnYkXzAnLkclh8eIXIpI
Xcd7ys7GUZdhQSrDSE0jtKqDz0fIOODMqb663Cj236ZeF4ZaC8Uo9OM3ALEi7C5XgzeqOJYqbP6J
ldqX7oslz0962iMk/D5gbv0cnWaouI4NAZQTMowvqPqLSXAFo8WhNcQ7c9tgZACjTBnRH2zsPWBB
EbWnM92rWUT1ywNu1hNJVJlVhRKrZqts1Et5Z0MUp+Vh+uii1QobY/hjLcHMDqdJCXPZCaHtyquJ
p7R8Ql4O5p9r8t0dSC+2BQgT704PCoh1i1Ictq1Rw66x2jMop3ijRTJcuS2lXsseQ8yPy27L/1Gp
Q2ZEWnD7AyoNAq2fnaX5d/R5wrhHbm0V6yr7v3dRq8Z+3AvHZ54D3U8qmQUXiJuaYWXgMnxNSDDP
97Mfm41shzXQ5gKhd6NnbMEelOyo3jimXzsJqanvI1ZS54mvSlEw6M22Q0cfM92qQOai5tfypXG8
IN/rMhnqlIO1C63xSN5kCGPJ6/y/uujDX4E6qv/BflMm9TGo5/whHRN6ImYD9HLiEl45lgtIFyDx
ebU5NUzJtxeieeXFd9Evoaa7H4Bt4v1OTakiANbJLLriF9e321bepB0pr7D/2mI3FO4EN/MvfFBM
vfux+N5UyJGc4fvQZQkMpXJPGK0mtP1roFFxWLkpFBg1bsGvCUKI4Ehu44wuJGTqiDR9lKsB3dYW
Uzdj6+3R6pWeXd3Z3MUMKVQR1ouODWAJDxxWHG1n83VPQ1iVSdGA4qQTNCUlsuS63BtQQUbpcR0R
ObQzKBaRS2BkEf8LUuQ+A5eoyG+Kaksrfd7ZtSQMER4+Ox5UhrjFzLmGLx76JHmJzkrUkgiKS9nq
QiXkt3enzFQE2QOZubzfbWUe2sfYBtMezhxdlxyiInYyhV3vdayCrjjzud2RSkgowTsl8eADyXz0
nBd31ogh0pZdjdqw5Ur3ytkeiC9M/hE53UKWYZzNhoKjrT9BnLp5XRe6SrWH6jrvusLL97Iy3pCl
7YIxMymvYcog7b+mEqEyWeGNglVGJ/hTqgd5YdQDAgf4bwEqVyTeuzt84Plwh85qv6TubH59idmq
Ch3NxrAdsDxdGk8HtKhgeKPvLCxTGislLWG83eJH785NRDVHjphd5fm8bLgLiN3mNblTIftcIyBx
UHIJiozNvZrXzV42KV7AOWoqCZDxjkGlA8ll4buInc/Bh7YppD5zKdsw3hugLvWrtGgdA9+N51oq
IrLScPc/u1pCIARO2soQol/c354NtJX2PWiTGEZBG8TSBZjm/LY6R0BbBg3KWTGN9Dn+Tg7bZn4t
+z+H1TEbQ3wplzFg/TF55ihOcksQNwoX6GMPC5VQ4l5KRfZ36s/bFCHDrc08U0vdBs4ysUN+i3Xg
RJ7yc6r9nORRrthEaQPg0d0hW8jgj/AFUKiYVrsPweNMkoEP3yc02P/y1UaeFfHc2P4cfHPhqaUo
Fru013jlgROkNvgbR1JCd7z7vUqU7J5PlvOPDu1qduORKKvuJ609hGVbbmIsL8H82kL+9ssX7nZc
nYOagD3Zx4RZ3glA/ztrq55BvcmQKv2IgV7fblkTYm4PaIv0sZdUmXmt8VDU5t+vbkyshi8OpE+s
yLMl++md8iM3owBJQrEd+zBHEJSBZT6qIJ/XsmGiZGZJPEbc2Qii/Qa707qLQkRfJHLUEnkA1Id9
/ZMB9zb4NrfwBPq/sCCNbOEXWBZGc8xBb8ujbStXn7nbONnkcVxPrZ4gZUPG7IHh4sXF7w1559HY
0blJAN48amXLUDdCleyEFwGGNUtK6v/J7yVTmaKTyA0mj59oDz73XgbColBYl7jl/AE8qY4+ew2r
c7xhfoYsN9LUiU1gn5WI7rl7T1bBPbAgUi7PGc0Zg/RF8ipiEiMiEITPhB/MaDhUB5l11wlyxjq1
2hI+mBbphvG0AH0XEciX5lBJXZwDjjt2won0ff27D93llv8DxtVCzN4pAvJpLJuWTIm/ZTjYYw02
8HMnry9+08mLeJreaVtvkwD2+3w/et0p12hkMv0K+XlGDkvi7nJymQ1to5nqi6zrd5kLq2CKQBO0
kJ3kaiEVpsRyThTPkJ6oNp+pUZyjiHieZ25jh7a3l9xVsc6Gg6a70CMIKisE//UwEc1i7pFRfqLH
u3WzxJQDzQgL5Ot1cGnP/xEUMquuwXPIUjCxlWZHvY1eF3b0OpskW29aOQ3vDo+5unwHBHK9wJq9
txkLSQRZDJEiuBUKEs2wI7FPRm6zp/WCErDM5BHoCxO4PKDz174m12Kf43oJE6RNZkC5Q+f9Lq48
Yn/Bp3/BbqD/NHjvmY5B3bgPNZXyuYqqs0Yf0mZNhrJ26pbCmnEWIDPDkSMSKsYS8UCCF/h2IaWb
BI+kEpUETDVPnEZcYk2SKIMyPeI7FecFa1dPyr6Sb5krEJTQh/7e/orCm4TIrp6xvUR+hxZc2cjo
gp8np2dGg88C8tTwsKmvvZWy03MbOnuD8e29vU2b8eX5rRF6WJvm0519wJqL7jlmiwrJTRcSDotX
MT+XwT9ArNYbOSHUshxTQ/k9gFpNgJUVS0IMV5Ecc22Z6PdY9EIUeKwxneFCxULAmvyXiVY5Et0m
AmtVGAmMogQ4b+mOgfDYllA5fJyIi/j1/Fwj5BTUoTwKC6hSdsE059g3rAm/hx/0QYEOt0ueU2Rq
ruiSVJrP8QpzaoJztFkXF/kZ4+C+j+sP5De87vgdgFmktGhqVhj82IeARn1SjfxD1vVn7lNE04+Y
rH+TnKNI2MjWSsvHdIivBTqZTiHBYfZ/tkLGXEaquUc/ToK9dZXz9xRTO5BcoCTvUyGpf7UdEXwd
qHJ6OJQ5liGAB464F2xnTybASKyCKKp9thxXWe4gbXymUmURweoUOVMQpb0KLLXzEsd6ITKsVMbl
WG021fLnAHQCorpK0wb1hxgco0+QRWpm/GZl15W35BgLI/2wNQTDxz8kwepuE6cTGI3ueyjNkyl7
Rjifj1x6rIqev2hajc9KLanKVFLTU3AG6a/5z+erJyKN2nxxDep8fmXien5r08zSzSo9U/F4pREH
oWZiLy4/cjLokublVZ8ANdQAKxe5mwhFv412cl7xdo+hvjbLXB2nMz0lZIthbUTMQH2w+juo7Ftm
VDnwdG3gDlOT5Z8oSdmPHTUOr1AFTnI1EkeR6y0V4q69NXIacyIZEJCdpGlhNUnZlssn+uRLEai1
ncam7+hU+2496HlGowif3pFjr9d9PhMpF4mQ2rtDJzIf25uS2dLfgbB6jINSCXAF41P9yH++OY60
YtpI6Px/9G21nVJgZdpjYin5qgWjoNcKIFL8XiW343+FxIdkdP8SKNVX3LjTgE9kgGpcOWkt+fzF
iyB4Pde5HGLkDQEb+jyej9MBpjSaXFDf0W0llqyYwks5cMyA+F4I+VzZIEZkQ08Txn5wFZNqIYfw
ENQ8UlO4D6X8O+NWSJ9yCfp1hBN3/oUG4uew3MhlB4zp6iNGXDIzTVMo7jDcOpmpQdj0zhy/MEcI
mxkPsOKqsBxhm9OK6PPiPLeZJCYHAoKAHVZUgRz17UoDf3W7Zchvylw+MAi1me0/VxoVY3Apge8V
Ui0CczSVj/12eQzLS8eRVHXX0Fip1cciVw6c+MTmRKpN1ra79qllnGQZ/bvqUTcV+enQ4B+SgW91
WvWLGBynsy/TOBvjH6VtkonScuGfoc0D0Ie00Jsjr21QIbiyqD35n5iiFGvoGEq8eYo5TTdmzzIa
cdfOv6o8XvFT7XvWZYcz5yHp5sZvdHoHqdjgi1kXXuLZStQm+TDyrIBj9BYCcI+g84Yui31ToJ/g
h/AO6rVq/mrEYTVSlcjFn3jeQa+4opLdRWFssdx97HH4Ax3CfkmQrHpXgnhiKez+N0fOMaVz+8TG
S5f+r9ml+ZnLqczM9hqUQzl8Si0X+OcJwdr3o0ovuXqs9tMpI9QVTyLNbJQpzTiRQlQvUMCHFGu8
NKIQhR5/sPOhnnrniK1e/nHgRwxurDaWVCfcEpRLNtZPR+RhVgZ55qerza386Bo3QBkf95s6RyvH
gGoElLRwZ5XDw/l5sxQv6gk4J54GxrBRa+Z5ZF08SN3/2UaczrEFpgKmVxL46UG4YtHdSOSgFs9L
ONNgzi6dVkY8FEN2ErYllcCz82a4Z+37OqFxMSD/B6SV1nAgxzZgwAT68CX+S/nG6Qyk8R8gZ9f3
WtT12VjfwFNunQklGjQCcLtR/S9QehoiV9xneGlhx7pLTnNRdPABYGbDfK/hwHO2kxHkKv9cMvPe
wjQnYFOoiuUz78CYSC+vySWU1B5HvWZoct3nFK/pGAf9wkNWxBmsvg/I92feUbpaZmeukG2/k0ks
U8b7f2f02iT9kN/3hdnqbhRZPJXQdH8kWfdHzxvnM8fuMIQO5Zz2JB8rNdhuJxFA4xjBh4pp2mfc
yrmmwjM4Ja+ivh/6T1Yy/qe0BcvgDXwhc+NkL6TBWUWvaWo17TWMkxc21uSuyfFDV5K3U2+XgRor
z9H3pTsDfutLUK7NuJYtHuGFiWzKz6sVsIsEv+sbxxHcrUEzMWWIKEs9pDt+7ILaCCzsYwR+IMnX
YgmJ/8Ssb8usimrOlu8sWG1iQJ1HTbVm8k7DWw+wytJr3nqTONB4nTHItudsrFnl9IR1K+I1sD3C
hFy4NZe4Nd9QR40Kd4yZ+9qP0LAgINQBiWkwCyM0ey/MKmBI/ES5kO/NsgMkVxEKRlz4NMG2iFjt
TsP4ievDxf2hpMzERo5vn4WFJQOHOznEfMHeHCnCUJE4B3R7ntty/3aZVV+SoBkANt0b2ZAQm3j/
M8e862vhaJq4Ej3DqB74ncLmnPEziY6Tr9l8OjO18VI/EcDhL6uk7BXMPM48WApWMPbRcFOr9bfi
AhWq6iIba1B6LWXnpddenDuGWHqT0P37UFC8vpqX7dq/cl4Aw8VTi2DTuLj9yaI7OOcHr0Tv5zJ6
wooaHY/tIifjngKgXV0q8qsdz4jtKcQ763CV1WuwCmjtbeEUva6z03m0+YezMRisL8jPvW07g8uF
cGejnGBjZ0nnAp6VaIzDZGm1e3wX15w3xULC4MPwmfXWjyYPvzvgC8i+9JmB5RrH5dmnyt/uFwA6
5d0BjKXtwk612PqTrohy5sXJJQ39fGUYorw02znXRTmPfGVZGLmIWgsTFHhrgvCIQd+DhIuClmaW
6jsOWsWecL9avVnhYb3p//uEc1ZgWaiVnp579dHTTs+RH2Tc5iuckuCLYdG5zvQA/8IxIpvpys9q
CuG+gxPww6lYJqbqtpjM+7MqegIluLfgAuF1c1C5XxYiAvqFH5vogTMXP2fJTZ/vv+T75BiC9kC1
ShkxBBHhKSVq3gfjb8FD+bmILXFrYMSRXLXO7q4AfutqK5YPjTtaDzVBTI8pnsZ9x27XaHnW48J3
KGgP+LndbTR5XoQmxUfUqhE1NeekIT9RtUQI5FR1wxnULn+X9HIB2/589gMaeka6jE7SRprN8hAp
JlHGQOllI+XhZpwdGP4nNT79Lz7uFjXhkalm2rmu9KnFQ2JyTP/VVGWFLI+ePd05HYVNQg1zlqnS
CwGTuDrFgVDp6ONlq4HMWMeLPxcoqt+dvlDMw+3ATco2MrofNrzSK68Pss7pO1ZePuZMAW+kNsrl
+eaYZRwSEd2ItU4l/1v3ryK5qYiyfMXtOViGy2wvSMJW5yqkdQcs2B0invwnvJ8mEmh7GnLcVes0
sp5ADGqiG703FQUb6kG8D50xKE+phz0zGG9UIFzKCCMWBpF3+5+2LQps4y7rh+W2UtD/O9E3TeMC
3MxZWvTDGymAhK6hMzlPtAOWJV40pvphZSKU9yZYPnrQAWm08rpszMDbdRobX/vgdQm5yOgNyaJY
KibrKPeO4iTkTzLMOhzWx4TmVHh3Ec0WuwLGmgbbrP7Dtb2JDqO6lOHU18NKzlKcqYfsCSoZTmjC
uMTRRBtuXtp+Cfo4PJOoRC89cLUpn8UGdrI9Dq4xyZdARgae8xzKX+z1GxWfeKDeC0oOWiI9Cjwx
6SXI8c5ylo8VTkAuPTyhLbkkds3R3C0AxLtluLmJzs5v5WygjuLVOwo37xD1oGWOYAhwQBmYWOsl
IYCwsITm0k6DHmNkhD48KoBG8guDDnQsICWj5qC7820hM5TgePRjzcNXtc8wvigHiTg2nUb5rdvn
AqBf5ynYJyy2U8VEUQIjPN4gZPwh+uZmGOO5E7JGQgoDr2tghMsw4+/boddrMPoLkUFqY6Zgyypk
xdSkP5MdfuYTTJr1Um5wGWAK7OjBELwUMPCACsMYI0W6kQWyX1hzi//ZDG/mfg7jdJk5lLSszTFH
07ruBgu+zgI+M3pnma8W0rNcLHrDqcquASGzqQwdc4VnnBG4GRZX1a+S2zAaUhO3AvgO3EWZDUo2
M5RM1MjnA6zLDz89N95lcYGI8zFPFlRVzQhoxbBEU98FsIMX0il7N25lYFVdqFhc6qdmM5wMPRA9
1cZZIjNy5dZyqFv+8R1JLxOsOzhxsF+iHde9/rOJORBIdDOhUQIQU0w921358ZEXkumCUuDac3sr
jVkIKAPLnC2hhEt21nW9Zb7yOTrrHx5Bwo/ZAQ1pvOR+RqoEAwQVcb2NLbQrHVorYIkilfkLALpz
PAyt4CiJy3DZFwh1+t0nXIZjSx553OntKwjLqcPhqC8LTztCu7OPIQTBIR2IrfJKbRDgc6fohKbI
9XSz28SawSCIBVOeTnVh8a2Q+S8ftYzXoOwydeQFLsC8hW6e8OfTQrhr2GFPNB14VPowmfh608Rx
2kvUrJKRAENBgYtvravK1I3eahns+jh4S5gAbL0uYAAPcKzlE7+mpHcOH1RQN9IjJ5KpKg0FrPxb
m5XqAHSlAy8vOl4yPYEHJkI8urJcrhUHB/nTKoA1djeg7xOV8nJd8u6LHUeevSmIHO8W5jApM8bm
+JrCAc58OnThvV1WQyuI6/jEe2LlzbVoI7zlpYKXXqAP/U0k0WKaHDgc1gEiJw0lb2QKCbVrZgoa
ZQyPWlqmyfMefJ6ywPgOP8tS5xnrlPY/fOftI0323oiP5Rsvyo3BLKEeDD+U8FDkUJ2nTFoM4dUQ
riYWoBLNH2m7W2adnxgFwqboCTdK9T6jX+1YEBEhAOeD8+uFtD595s+IBI8inKzJknOmpciPOenT
Oydeui82E2Ti0PbLJ5wf0f+IH1Ip1V+vhus7OlsHy85b+FTCIEgBj5xr9QniRszuPEvgvkMjhOF0
5cwFt7FSZ18PNzNOP5U/0CJJMPHuM0TEOgY0mNWEHY5rFpLrqHuvlcrjIRnET76ri4efMM5RcCX/
B5iCMPBIHCMrkT9uVGu8WU8yHec+To76+5Cx0WsIoBz+rYf4nT/F7IZXYcgIdJnf0rkXWHGYl75y
ntVBncjtNGkbbBqouiCmEKTcCHoGEaDWxsYHzifv/zXLovxylajjGpkj1gr0yRch/vFVNGNROTY5
2V379+/URJ7BoHSp6VjJtYP6N8jVvguIc1TagYUJuwu2FTzDjK1q5I6k6tR0S1jF+ifsVDMV9kDc
PbnttW+vpKti7/9MLnDbY5WuJxOe/4dhHIMg+2/d+Ddj+XvESt6E9FvS2e86ynbM7icvzwr3prgd
asu+WvgHtEPVP0GWLmCKk8baBDKg+Li6MvBvGLyrDyp95flhMBUgs7w8bOPSpMz6eCAIzWbi/XOy
uLx9DhZQbo4JA1zvIN0yXb12ndqd8Fa/8OWG4W3PNhSWlKAaJqd2BabIF/ZD2MmALwXwBHPsEWCg
srCnybI1TX02MrwogsR8jm2lVmtYcJrajqPGxNV1h6qjmUbHWJdYRW6YYjrIAyZDaZOowczROrpB
UtlNsxQQu0Ajce3QFozZuBm3m3aPZikImNvOtxp5+9S1dLR5Gmieu+Y7lIHiXsunIKzUhzJNgMuw
w94eCTjjlSVZHYVFZe4xxIYCXX2HonRTNIJj1KdZzc4DpDjSDQzGN7GHrjK6Oasto65xBH+JJQWy
AYsKnE288VfTQ3R4iSDF2U65mO+8avrx8GYhRvf0gl1UrY+bzinIiFCOu7/Y6ly9R8ZdxtB+u/7W
zmZKm/xQ+jSYuQ7RJ6ewtTH8cpS4cUM8xyECRqk0EoaWjvWJKB9vrOYexXao88Fn7EGBzPIbbikB
l8IIP7CjAmrtfYQJmluadmQgm1bBM5oQD7FuCk96ISQKNsv/h28SWj0hsYZuLQvr9tXQdH7i116Q
1AJU6SIr5PrYwaL35ppl00SYJAveFD/OkgLHUo4vawMzqmf9N4qdvijiFIIuDVe1mGMT8M2s9Na7
53PVa+j9mJiSyAZKRUmtpDbTCEZ7tMsvlYUCpt6DMXn3wNpy4A7Mp3EP+qgb6+Q3L5E3ar4+7nnc
oqW1ceZgKs4L0f4W5nGCNw+Z5QiN1fJGQmPMBCjcZDAiGWK/Vjp1b6vP2Umr3jwWX4tqpolZtFMY
OB2hh6VbQ9L/MQgi6eVInF7VA/s84AxoPyhlpxNtagZIrpLEcw+arjEEgGlWtd9x8w0RUS2Uw5ti
qvl8//5WuWQyUvPbgk9/diN0ajcVdgL7vb1YeiJrlhMdAAaNbsUv8fiSMAUWi5ybujNAyMfOKpbs
hsmTw5+H0VhscOyCS7eL+Yb1IPhX6SWlAxwXWV/ccuRyU3HWafD2WD4jwfk89W/24M7iva0qOmR2
KEfqXBH990HstRztItQCXIxzqr63faoBj9fPMeqUgLrvAPJhoCoyhEYLwPuOrsfBtQVLcaCb6SeO
o1CIhOxaj2WOQMeTqOq1Q+3qehCNfhMjilfMrqqNVa49veGdnH9zbivp+oD+T/Bjde0smURK7ja2
3ynOTWTns3cbAWI9eQ4x1ttXYb71CkfF12ifAgxZEcJf7qpXyyt1qIj3u5OSrzCZ/c12OFnPf0/c
6/85GkF9NFDAIUfktdWcsQgm8AdOrlH5oqJ9kw4NX9mgo7YbUqLOHEp+Ft11PQCWbrGStM6gzZGA
8nWC50TmYBQTTe2xS+QVOiuDUmXgQp2fI2o4nfQO5sp20ePDTheWMUmd0zPktkbv7UToTY8x08nw
hH/imhJM62ClQKNa2FzOHGA8vqLW1PDs6m4hoNQu4KRo+wu8RDpMzYUwTw1LS5LMYlbM6qeR0G6A
Xcd/C5UIZCiDjBCSX6ON4gWwZg+gYuokgYmXQtxWfL14T2NC7Bfxv7EklUu+9HmKOt9iqzgOkq8H
0+yqcXcVXKtq9Bv/TmvfA4EL3QNQ//wu25ZGD4H9eF0xF9xVnV4LWrkjglF/OFdDpaz0flACo0RR
8B+UaFYBVTOZR0udbBkOAaWN1AzDUjwy3kS+4E8HWme5OCtuiH3asPQeJSP5BQOaRVAQLLWbmV7e
ii5QsxWbUh+32r0y6HBd59j5UWUZhNa/eXQhX5hDvJ1WqTiZfmeRLxE6jxelNKDH0GFQ8g+q3qxb
yAhmWyiXV6pNZ/sjueiS4Uphl6VHW2tKSoiE6JfWSYlMuoOZoZxKbrKshauYpBstx+J54FJj2R6O
1Y9Jt6OCYFWrnP6uKuMuO1Z/yLsffUPiNC8ni4YyIffsa0Pi4srI0jnalLTkzy+hqT9gZ71VKZC0
AMej5BIidxrDDEO/NbFxCDIAGU7FxGxlvF0rWB4f9hkCWesesNQoPcTAAWX4sGU+axxeGP6eaTuC
qAHCrcIbhQuxGOuujFh8Oh6xaVLNzYi/l0YwUxnkclcfgjfmov5kBrtFF/Ey2olLqtcD4cygzngM
EzH0T4m2ght8ONiFs/u0CL9fe8l+0HmPxrP8AilHCmPqgOEiKQs5irAkyWZOrWLUrXjhqWbtHk/8
Ayu6c7Yw7vujkHppyXjnqodzvCU3/PbGrCtMwwtpkrI6CPRG/pqESOccjaBqcRfa8VpTc0R8ROjq
dV6+FEtaXLmuRreY6i7Jp5BaW+u69c2vTt9QGHY46uhdPTSkkZIiUtnvcxs+52DTUDZD7QALR/BV
UofMMiEwDymwJ36NwI+zkkYGabu8Qb9ZHQ7at81HFViGtMzfSbRQXyVswqHWB1OvNfobmsuH3pYE
bHDt4xrZaOcv2EN++aP6xYh9RD4cEGn4hRJBEdBa3RMu5FjehRG7S0zCDbclPuExoMhOdbcEd9aO
Yt8FJsKMNEOWi0pdH6jYT656jHfljKfN86R4SPvxe+/4rFQhbzVd2aSFl52Oaur4bVNp2UGK6q77
tq4SrObOKPfGRJeMIJTPtubzoY9GnvndyYa1cldqT3NF0qx2cWCi6tQaqv6EvC2PVmVISkGJbx+w
qRoX9nmkIpR3p/FK3Jni2Cby9V3UPUJ1Cm0zSJjEVrmZiImL3S9WK45UeC5upZVOUZ95FehR+/0m
Q5NE19+KGiSOlUmKdMQ+yUV4btbXRR/xnkt8orv07/DupShuca8F+zU4Yteza5eXOp+6oB9Nfosd
Ps9rHaY4lCfyGa9gcBdSITcT2/wlf3lfocRAnpMLis9Nb5BPWbtYkdsn0h9YhpLgsmPyn0IAKQKJ
hzHhJM+iID6Hhq2FFkL+kTXZkZXBmyXvk5ubhgJVf4A1kTGuC48NpSP9AZOKCY4YYYyECAbQl8NB
OH9AraFm/QSHqIKse6I7aplNHP5tLbVyIz4HYSCIuaOzQZ8a9/E2h85OYn3e6JVZmeUHFh2V8OBx
o1Z/bHeuXHXk7h9u3XyeE2oKb3YGJpeNUahMJMpOmyEXcK3AlLRg+/jR+YnRgjwCElZGacS8xUsl
GC5ro1rEJPgQvlSJYRGe7rLZe4qY5K2fHLxLwTXC72kvE8OCKXL9KGyzrwrV7+HGjF4HFnPyCUN4
NpjJKtBE+BS3xyWjb+pIP88JRKtQuwqx8Dq4Vl4p07oaHhZGdr8Xfe5dCESQ8I5i2ogUwUtMnXGe
o0+ISQXUSajyJy2hKWcdphqiKeetRGVYMDcZBNhsj36k7hYJq+xETU0GvhY1/z696aKPPzywCUDO
aXAb+RLNCUriPc5j2uVncKyK8A+cn8ppAxi02qHLRDKYSXbWFFnnJh9BmG0+mFyZYt9Q6pbcv10O
iMypHyZwbwEYv8C2ImFJWqpvmbQv+I9A4BbE3EH//19lGv1hotcNsj8dHvxMu08D0moXPykWt/aQ
Hn9Gxe6Fp7LF2dndgRoZby/k8Pz2iIdrx2dVLnBHwOFVDg0NvofN1liqzLaF5NChtHWROROJG8+J
BHWmS+Rc/OmJh2vJ5El9pIVW1jeXuIj7h1iOGUe55th/1BCA+84CtcdRJWFni4zAtrMUS8FjQHrd
vbWLtEqFB+nOHW4LdA60KBrDEjXZ1Wxb2Pu6hNHup9ygTaJvRZONjg4aAkYIfq5Bojcp9W12uQ4H
ExkRrIGXpSEkqpR/JaNjLGzGzt/GvjPl/mq2iKk/C0oGHdwDDaWSz+wLl/j075JBDR9fngSWppP0
8HAvtmM5kzIdKtLmnCclT8VA/Xv2HTJ8J3AgHiMYt7pfWJjrsR6NeLdqSmkxhIyWCpDYm1ovADtc
xrFG+/05URLZrgubV8SBjHqtpmlxLFfpjXvGcumAAf7iQiOnDI7aaQ+hvRkF/qJqTx3aOoqSElcZ
DiUuuZUBJ3RAqB7ubN+VsicoeJNeQvGINYVPsZg9kd73D49qV1Y76zoPkpBz9ZWzOHf4Dbfj+RfV
AgeGnBeOjNIRwgZeg5eNKzp1tROd1xxcg64vcmbqX1tn+cWiP0sd7s7iTOe+ojCq2v9kBXiFOYoc
DjbSZ0UyRwSQ4ZoNGiL9bVQIK+A8pnKchjeaUksWLFJtVNWsZhEtyE+zvXjWpDv8cm20XK7MlwTg
Db0AXdjS8w1zxPmxQk3bNtcOuWuf9VBPg6HiqxHj9v2z/nKj221bH3b7ztVJVGPmPaLvS/xPfeYV
kew9Bg3yXS405tQqNnk22L4PT44k27L1JJU4RGgsQeTvsC33N1+6jvD9TD7eMth9ocbP5beeydxy
AFU13VgHTwS8elOu3FuG4rHdqxAz7p5vqbuQV+K9oKtxR+vThaAT4PnS8tRR8mU9/LtNE5aL5uBA
IlTva/qTVIVX4Vg8qfc2irzgbUBpWE9Gu7qgRiyS5leqIXwasxlXGl69BKvroLtmivtYnPV/Fbh0
Q/QJkjfmyRVJ6X0OyK7F8XQO3+1uYqKaY8yKAE2zswegW64gzjQjoldaUgWIcFTGgK29uSTMPOy2
S/rcLC2RbYFK5qE1xPSqBaIfa43DMgu9YfR9q3/FM1ZfZJcHjn1uslAvTqlZ22i87zmokR0Nz26Z
zHhjAeaACdP/D2vo2EH40duFKtKO3cU/FLoNNpZF3Bda7BSXH1Tv7rXzKZEKVM8S3tfG0AUOETa+
swHBrCA=
`protect end_protected
