`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 69072)
`protect data_block
NS7oQ37INqEm5wSYxoUhuHZVRqYcdYLDTpOgkDtFDgCPul1jSmHaEsMBOnQfisxIiARj7dRx7w/i
Ddmcz9x0UYjhkEOGE1MBJqCycSFlYCOBec9W8ded8AeX/S2YRRPXhGkG/izWE61IFeVOje0Boj6Q
xrzEQuUhF8ZUHWBFK+A2wtdUCHGdYp/MatboUmKGtVpA78XbL72yogm4xQOp/22VrVQo3NMQnylY
Pvi4HMAYb6cX9yM/wW5MwcCrb3TxUL7Lc4c3ZXpQUPRNWH/sC2A4/oTyLM7PfsD/G5h33OC7d/d5
VxjcmupoqwlIU/qUNTx+NSBfQDHbHVEq5JS1a/wgQ43kWcs2oljfdPax1Okfhgho8a9FU7mfdSuB
qtqCLmmFMLNjqkAQJ9GNDPwY8ItnMY23HWSJ+D/9z65/kzb6KWXlJghXDCRgRIbD9JvChD3ajPrn
dC2eKbiwkk64fryDt1jje5tGm+VVGUFyIn5GLaojE+wFCjf774G1Xb3U+Zi+dZQCAao2gBrYXTVo
J/wa9sHHM1itPMZwjFvDBgX3Yw7zMq443tU3VQWZsG9YnsKWTmwvRQyRBUV9sjYhIe9OWOCjzy7z
QZ8lfhzVXdYhiJLLlBcYxOqXdSRVnChDRlNQKHhtwFeogtFCkPtNGuaLciBRLFId/2UkfaDyXCZB
YRVNKQXqmssbx2qLwtD+mggaO4ila9sJ94p5JKveGZovHFvpc7KimWU8qtwcJZiMx7nSdKgb8G67
i5b2zVrcngHIjyeiwZd/ywiKDwALGj/VRdrHZ7e6Kf9elaMw1iCT2+XoUXK4QFn6aDtK9/Tx5ssk
9AnoGmmL4Xc32fpW9csZHf1JAEKtVNDBMjhUj/Tu2s1DulgozWEESsGgJ2dHhR/Ir9x/74PMYvGo
dyNft5m4d/oDPLVE5jCqQ7Dk3AIQk8wIGs+C36Iuxv8OKtBNiMyrMwWe3O/IrUop17qLIM3/EScS
UxOqxr8dp4SzzfOWOLvCrGyADM9J//q5w5oemLZm6w/pU+uzYY+ctSzp4Wlx1jMGdqjoq1U27mKc
5kibXJ6eBaJVQQPa2STKKpe0OKFGOpyTpkaYf2NC/R3nO9FsOjYYRb5n42X4kourky9jJHOkdzo4
t09tr44aK+7lyp4+JMdh2bNSVNjOZXugSnzk2Hx6+bk2nwgP9VGu30ea8+qdmAY5GcKG4lrZClKg
7GvKXQ47WV2hlT1ZlSYUysNzR0ARpwzsgC53tmjqLE3ubatlIdayFJURBu5/ABn6EdluH5Eyw765
pOeWbnbYIwAeynCajGRgvY9oQV2ca3ENyGYgG5BmzB4AmKVQuP/SY7+yBzoQE/B5ViYa8z/EG3WO
5vrtCh2PPEyLjv/gpG6SWC5vfbNSKr6a3aLAZKq9R7qOQ1OWVYpRsmyZtr4/HMF0K8umRIRB9x+e
vLpzQ7L+KA4mvh1OouRMJgPPoAjWm1qpKwebOE3WfChjKFP9jL+HOKdz+2F3/Qf+OjOkjrol3HLD
4nCPZkRrgyZtHDKqTILiyicaceDt+cO9oNwfxNhag2pg/LPaRrGlGfOxJvUSX5HINEHVJTSYaRGr
s5JE6ZCEzeJ9ciOmt7YjlIYaLaaaxIBdWmRF4VMEhV6jey08pYhIbhDLHw/nA184JS3/VBdjsIDU
Y2RsFE4+panxm+UzSoONJdik7bVFva/GybXPXv44iHZX9VofUhHULI83hdyoq5ZKAV/tTlZCsfSJ
YLDrJFqb7g9IIoWUvnw6JcUzjnYOqN3xL94+BSdD949wUSl/MY9S8xeIuJkBvaOP/IXP0NuurRZG
twcPXA8dFXGzhRHVzR7nEsVHmrzyIDmj4405GfiFY16h4LgefahrJzppilf/8CIz0c9BJ6Mmto9P
T12iLNZO3iDDBc8MMnXGFOrj7dvb4lk9glaxMF/nJ/RrjFp0xg6Z/xsZKMxcXoP5KOfRaNXae7bC
dkT56i1v0Xf1qcY/FxaUKaYrMnAPZDGu0XLedP3TJIxl/hKmTr44EPRyHcQCxi+9TnL22c4AaJBz
90Oz+/Zqgvf0YzOKvKEtTCYNiXeu/2KdASBSUAdAdx/1iUYsV3rwfpPzOdmmJElgYhgDpeYArKW0
I7STS62vaInlMwjhzAkWgpXRTdtmuLS+vNLwIAqS6MHjyL3ixrs5Lp4SG8+N0wPRCHjjWuWr0C53
rk0zoU2/j9coO5rts2rKCp8BQmTTqIzyZeT+XMBXg0Z43tUmSZyDE6ysqQqGvocd4gCUHCbLA3am
xLFFy9WfFAvfgKpAcewL3pBaiiu7POvoPjSAwnP2a853gir376FpHeWma5FLJTJp3OqmSPyAQMX2
205hsGHT4vrMDtVvz5g3F0RBRB2MA6UxvCxU48KWjt0S3VgSkel/aDD3w+5a3bi6tdq4GUmqD/dM
lXxYK8vDZ70jejDk8alohe8fsMMwhziY4Yd2OoonJ7jXmU0rp0MMSZ69K2y9OLOWxDP1JQIgiRh0
bgtz6hqnTRheKkJe/thjXAVN1s5180EX666Z0dQK3stWE0C76oMJK9exwQ/YRcVWggH/q8DRMV+M
ntcSe9vANXqDxJW0D50THkwstmuLKXqA7eIdyPpqvER/i+B6t/ETkJ+nAdNyqZPPDyJwZwxsoAQ8
pkg1qVPvw2Il8Yu1DBQeolbvKs1qmBQa9oWET/Y+Ut24j6l5iLrbP3MsFnY2gx+JvkjnfzaRyzMM
D/42zGXeSjY8qzFTg84JOLm6XJmVTB/e9f070DE/tFDbw79rXjWJlz3Zt+pkTAA8heKDCGTwsBsD
ete23zwpfX4flXB/WUjkI1j8rLPFF/eCiio535X5wxm4CRJj0fimKwe4+7MfGi55QyQNV2fI8f20
15yDayxny5rSSF/2wdQUaILCSTTTqOoBnKruBtDNmectkhB9eb88KFFzhPoOgnfIX7OpfbidFJiU
iTludMefVKwua1y+mureFx7LUADJnZQzmWLLpJ6NQLdE1bh0cNkVJ8Wtf418IMkylwfy7pHX/8ss
ga8h733ijDNJcUo+wzUfUM+/HtlCCjo2bXottoejdclzS603D3rr7Qkk/E7J4E4dLXyqBrXjGmQr
wWmy4qaNw5+Wpp65N45XiAe3jnxbFwRARdS0e0NL/5vUcFlbJEULPXdmCe1854du8rB0ACRDM/BL
JFvn4MKb3iJt3CN/GRg95yDKsQE/ZvzYhlUN0MR4oEBu4qXXDz+ptdODY0zbnWfLBAcv6Z0r0voc
zooxcySH3DC+EHF8Dv8bVl2y/hKz2HPaGZZrXSEED9TtmvV+3qpP9zBvp7c/DvZvo3QB10Zb8EUb
SSecGok0DuEBvhqv2Ook8C63t4LCxdPaPeX9IsbNrRnpOKGfRZew3CI7HE4JvhUe01U16+9zlV2O
EnJ5LBeZtlpxsuYIp4YfpvHP300DYGyqE+A5r65MKzwxTds475FVXPY+aDjUrTskGH0EIE+miSI9
Q9fW9A6aU7tg9p25W8vUPxUQBaYk86MlPKggDg11fGEtASmRQ+krMbPcd4MGCOaHnJmnMv9VOy+s
Cyja0J5GEvcpX6QF2M1I8aGffzq3RRraZmDpGCaLzjRahCEPuyCNx0mPDc1t2uu7O92gomvkNZm0
cbdnSdC/I7/sJjN0/G7ZikuF7DHRBKQrrgVpxtxsYyEVGWGKsJsN/ocjgrBqgDAbG6X37e+O1QQ8
FWDfqo9HLZ1g/NebG7+LQmSM+xGVDG5wDcgLpLhvFCjH7+i98xOeuSnsmSvm0/aVwbDfiYBnnHd7
30E9IjeGXw/XCgSHSXt6ptXHFruC6FkvxCzmoYLOr1GVaVK7XGARFY2gEHxY1nQw5XON0oW39BVg
vEhTr36ypFpsUM22Z6iIrpN0yjJwNyHkNh28R+bU77caYcCzMqhmv0zEDTzzSKc0MeSNMhtHi5h8
9rs1K3esNOW4tcrTZrXBEYFwECJn8OeqawKq/w2do2/28t6pp18x/+c4oRWr6L3gBtEfzIVR0EtS
YS/jTLd+3VyUIKvkx4/Tx4/eC0xKKvp1H6WZU3ebDFj2PLj3kyKIbhX++C8TV36xbhTxDWUVgxwm
+KwzZdqU25WKuSxwEWUdq7D5/xQNYqMTmX2BaRETAz+6grYfLfb4csCAoPrzO3tm/22xkBhKXfCY
wHuFdtCGSoj821WqHpG9GeZKQR6OLba51vNaLMGrpUVdu1Cfuy23FD7qetS9rnPTzxijY6lNDVoW
/yh7hZ5sUbCUkukcOEaZ0FfURewXMqljB4hWedQs1YSETfCs3xFkeH4Cd4+ftJRFNHpl3+42/VgO
fcIVoWX2jJAwaB9L01YIl9P/J1NHsi7krFbB1+wJ5RVmxNWxstzigQUt8fkaKHXuGf3E1UIXNqyy
bQZr9JxGZhZdqCEHlX10xo9qryloBRkvebxHSvv7mHEO4k46Yfv1zwCANJ4pdYFrtgGQFE0FhmOT
1AtiqmPxiacG74jqsFrqR0Y2mNdTfg0Je+/hdneO0uvUXD6+a1afKzm3zKv+TVknf/vMa5ABFm+Z
cqeyfIGRc7s7+6Pr2TIcXv+J2s/x9rToZ/asd2GJVKNkblmvyuLQz3/ZVfab+k2CA2wPbcmtU9gh
XeV7wNbKWZqMA/RcYDiHJxHMzMp/2UmS78O732TJrdOz0k2el/vOL6RHd/GcXmyQGNDlGzyHMknl
ZrkqJLZdrX4E/BKgQ9PLm+2L8ltvh0efDcA1RC9LM7LWWAllf7lA03sxj7J1aRhnxIkY+6SGZk3Z
N9kdxbkhYGYUpvBX4GSrtjsgswEl8ULvNAtLPT+sEIr8mDkSnLjGZtcMiob+fYt1TQqs1JhAZ9LX
BMS/iAFtkR6UbgQ6UN9T9uc7gXrHEhOckn3wAlteIxNW2bnWCeCYoFuhNDZKWQ3VLgMOInCAILe8
QvldBqtqeBRtrcz4bDFZwUUnO3l8RhtlpqW//bYiVHGq9StWvEP1WKm9RIghucj8oJVplmfypqFO
ODigWGuXlmH5/tHpiaYG5N/RrOyl56f4Z6YIlHtu5HHcuBJFYMJKHTm+zF4SH9dfziBj5B3YO0xL
HNF7pLVrOjZ3yA0Ca65eTnDB94NURVpjdf+mwE0CwS215kx5/xtcF5r7EP02YidFgztcu9MAygJ1
HoB8gFlBb50X6w2z4LKXzqzX64ESyNHhVE0SWW0FhO35b0wCHk2vjLRAxDxxQoBt97Gs158ssfhA
wmFeDoSCC+WWkDp6z/f+8ZZfbI8dcARhwc1GLQIlpFgGll8EGkqsDqGGYhKBfjHa0U/6VFuw04DZ
KLqX5kklj8kW0oz6ZhFsztg6IBtevIndep3MjfMof2MX5hK7JCSihcoC1M3UzEsDbGLVc2ltSep/
9SsY/neB6uvlZ8cNqvW0mPmTb/OXvixGiH9PYX/HNCLC7g3SYeTnTBHhFsBYmPSS2mEiK06zoztc
SF4/O1Rqj64aPAGnFxpfbjEkzjCUOJg9cRZ6yLd8Fw+Xkmbod+h1euOeIILyUOCQdXT15ufvrYRW
2h/7BaUB7iHcwwic/V2yG/6rudXBeiSsGG17byuW1l4eZHmslBek96/FYpsYpFK9UTRSkE2g79iz
9JaqDFRLsFiXrDwpxXuM187s2cD9MNuU4LPdHk68WGKq29q1jZr9vV155x0EKq7YBHLywJOhDSyj
npU6KDjh6gNfH0b8NsNrUTNRyfZbbUhF3JlhUBFkH+fmzxdhtW00pWrrq1HCZhbNPbeUxb6wWo2U
fAoUgU2vgfYe6wKUfBhswPYrM4jIySdNnvSaAOte4zJxpgaQDr2tbxtQa8UIO/2JlRDm//cAGrr4
J6UW4EzkpsUJBTg+FzPdWUfBdd91BDn76UZRvOYpCvhvRXRvdP7MePmfDrCX8FpTy2yj3sVRBLat
JnxPAes0O9s3mVhAltfkGGftd2n55XXY3+VgED0NHk+EUdxPGSOx0p3oD8diYY1CVb7LQqMzZHFE
Tvj/pIhh1PW8EAIFHCPoFdNefDNdj9F3nQojHoSBNC+hYhJm2DH/NcIqCP1bABmzNxnvovZZCUQV
5OuQArOmzBVPVu/qUviJU6fAwLCVDFECHrd4mGI/TtzkE/wPS2Y/ZINQ+30GvkRfGtUihsh4tpBZ
tTDh5JQLg7En0hN77+UODoGOvFKICqdY2HVXIXnT6p8StwCsps5Vb8X5/103H+DcHoAYO0N3GUbn
gZGQLIqeVyYvxF+1sME2SW+qnPfDlSDVtJAGTTPXvQy7Gro9kbAfj4/I3cIN4vJcVvmDvsqKBTcG
B32my/vYa6Mk6Q8cTqWHWm6iCWrcn+G0cwsw3IJelKNkjWnnRqJnVQmixeFffTrT4lIf+SEF/tnA
Q8Mq45PdqVPI0JIb3nsPVg+iQSIp1KZOOsV5nyZMp0YXm1UKG1OjNf2oVle5yuTJZlU4HePFTgJR
moUr+eBn0WmIT6T+Re0zimKX3K2U8ItsO17iGR4k1auzA5fh0glr4qeOtmTjJNSbGF3OLJJIKS01
/KZL8pBV4LrAp8dDOeYseYGI3GZX8qjgyCpFK1FeXNmqO15mmOP/u9DwZONxGrXd7d3W8w2IVsFF
ExYADz5ALb1Oww5wV3IYr/5h1refQ7+ZB01ZkeYWfRkwxMPx0BU/tOB3IjabTY01nMNA40szMkif
DjpQqXx4YNVuAub6OB0juu/vd1qEtM4gg5VqmYK2miKG9kByorxvgcN62XmSHSZg4MnD378zliPJ
6BdHbTLisRz74Dm7DKA8c6dWQZbhT9WFPrOuyAxsozEGQJLkf68rGZVJV/M6b0IzzAqWGseFbIuV
L3DXeBE4c2A9Eqvf1O/GYDV9bQxTx++GGSz66Vc6O2HGd57l9MLwlKSLSUUyKtGzPILhZkgpHjJ+
bbdrmjoKSimv1g2dcQ8CMOSYLaWU+P6lTxf9cVcCiqjlJmKSzHhbT5u8riZQVlx6gmEvCqguE+EA
7sRykxqPrqV/DXYUb0rbSIXPyF6D1dmT6BYVFGucHiWikpjNdSRxMuZAZGm6MV6Kne9hRWDdy2y6
s7B77eUcKmzhVn1qWkXE5Xz7k10G7HaW5PkhOy/dYtRMMeizke+C2lSyiJLq8MdjIN4k6mDZxraL
R2oNQ2VwHrizKlMx9hEEhNoV4xmsSImediRLujvfEEoBo2F1zL/xpZq7q8H5o+PIKXkstath2Xs7
rFPYdVL78bbuhqL1mjd6Ils8sxjhIaBVo8FRGbIkgJkcJeO1ewmZ+PYt3KDAnuaLqpO0FBwtq/ij
owfr+5S4QdLUJOWBfPxu/K8Nu04YGqcJIqbY6iAUS5mDV0SkohMar8jnsioFTcASX+hZgrJOAoQP
kYdgBvyovNtyCGXJBImpeAqII+7MXIblY8jS9g1zjpS5OVZMHtykmCcLJ6vfL8qN+2s+i7o60vD6
tTx1HC+VzxGZZy7yIJP4DlTcuy//LkdnOFG2x3WL9P4lEGrAjofGjeSNFNF3CFX7forkfBmoI0Fg
zXpQTVLVfoQyienG7SlB9hZKzvk1OwCq3q1wrFjjJ2eShOs7xZKXUq+aj6QKJrQu6L/lFL/mkhGz
sxrpA7LWlWhOKdQpTCx4TyCdtY97sVYEYQscgSq5fQz4r5xWEf2thTDGB8PFP6/3Rm4vWR9feK/z
myKjZGFJSJarJS/Gty1CE4mXhZBL43CU28jPQXGqw9Yu4MzQF/kHgzlBjRP7lmfKCuCvM+p6ahqZ
jfi6HWS7SYFl+uIdQCrrjBil905WLPbh3INbBAbGGsYDyuPchYx8XXfY0J2u/QoR4JXEL0oR71x8
qZ0wqwqKCJXOFaGKreHG4rQvUonyy9KvqJ+4JE+DY6MYXO4NyU2PBYy7Mu1HkFLwinbbWyReqctb
Gqq4XAFPxRpchxKQJ1R+alOzlZTL7qemE0Kyg0bOCkn0t4rXSoTVQXj4ki37JW6xlrZKk0H+2gWb
GuNFIdZoMtinXAqxACJE6Dp9UFc88lnN9O2U83q1oEWZj2BuneuAG2SsY+NiwC2bFg1GRU9B88KL
s2Uhf5BjyNGwGlPhHJ+4OB4F3MNJ0e0cJNdY5pjtAC1kushUV8kJNgnIw7PI0e1D4BA+vUoND4b5
F8USvNhoJf47ssHD12kA8OnWPW8VqSc8JYcxiQzckJVvtXVezZAac31hRztsr6EqzL7QaEi3D7Ib
XkxkWfKuP9wj04RjAwZXIf2D77JRTNJ/jn7ATC7hSFkTVeF/lzdoer3V6sz0NfPo8xuMG6/ktr4c
2oCJ1qmdgDi4o894RXjf6PNfr6nSoQz3Cm/DvGVdLvra3g5G61poHynLohojtWkHiu6nWOBiZyPE
VEmxggX5swbRJ9FhpeS4n0JOatcB/OR4zOipofx5sZRuHRobJRmSooXGJTRsFOTZpG10ByuhUW7h
KNFbA+6S5ut4ItoQqZ+Z54UJRQVeHANlaPtEKh1qItwkvSbEyL9mruYjrQ5bD/UDZzCcuKAtkoUn
jrSz4wwwoM7aNeqKxI0CGIXiATMuRY9z8IMGVVirYddoacjOotjlUAzWztKYqVLyuh3HqXo+wS/x
t6Vxsn18yexVBiwh62GrTsaru13qecT5TxRRj0KXW7ze69uVpa/2qpYMD6EfJidqQ8ner3SQmFAI
S7hRqGbTUj8pF74RDcAMm3AzZtTy1D0Ok/lQo/VfL7xF00oCHhV5OiRwu0Xd2jcuiowN1lsOzATI
pSHswMD00xmiNKHZSfL9IkZYqtLFfMQOOXhf9Bn6rslGPyvWraBXy2Pbj7aEWdQE4q0coCPld2z5
FuHoCknZiIvXkPEGFl1Tlozlfjkid/xe7U+bXbAsgorluirdws37dWKTG0UHHJE/Cm3LwEDOcr69
grI4LHO9ps544v1Qtj9Y3XErxVAclC2Lk6JNFc02ha2sLCLn/HgNX4tb86jJbYZfl2gxzej7Y8hr
waYhf8vseL5EZ52AOXA9ZzxtgEfNGnevboibc5F1V/ubAMycJfvuy/2UiBbs8iNguq6XVGdFmogZ
a3sYjhLoPFwJHWHSBg3dmMKFgjQXGJPAzKruwPN/xfE7y7xGKJRcuweai6Q9YUoqf0x0RpIuvel6
HOHmp/2CVYGfI/ibQnjlTklpVyCXoSbRP7OGynkt2sr1tuvslZK/G4PdhuyymexVXyqB1+Wgh4GV
HbwyQ4V9FXWlAl8pNbpu6mZd1AaLZvzPb4c6Vo1qva2+qI0pm8YKWtW8UFCQ4HyjpbMohbHgGVjR
pvHhZGFt5XJyE6+cI62Pf7kize63xMVUNuYZXB/5eEKrIM3yAFIW39CiBW3s3rsSziRB+fVZnapN
58cVho3gKsjD39iI8i9jL6QKDy1uA2RnjDmVkeT3FTHt3Le5/LbQCr/UZN6Azk4T4V6dpFiJ6Yco
4RKBRhLKDP2nr8o+gW9FrNaErpFj17kHP24GvkcxTy8oelhF+kIwMCj4Mfi90EPC9NusyamFtLKT
hxM8EzyoDmfx/18nvb+z47gjfTy2qL8G0q67Xr8QUh9BI7rHdqIPXfLTyVMU8KJg8/FmN0OuN62B
zek5RAhqzpXbp+KMPPEi6bnM92TuYPjlaYmiraT60/MAayqUu2/D7syIuEaahyZPLG/V5+m1gh3o
Fju5BVlBH8qIZdZu4xNUzA0bBo1gn2NEM6DDwuxDmEUk8kukJd/DW1jBGSjh3qf0hGyP4GCu+ry/
Kr09gH8hhh5uloipYfOxbtAo+xYQkUGVdJTiaGTn2xopjrwRKHxteCjtghUfRnUUV32y9ZZMmdPp
xtYXlY2Motbq0IQoTzMyBWnzYERruS9DF5IwK+fIXr3anCUQNQsKJzvA/pGvEcNJlV6O8Ddx1jNS
By0TcoD65h+T8vAYQWwlWzHrl0+ekQ4DEXpVQ7FXoq4lH2EpiMco38bzIpyA0pIu95JSYPuuO1k9
SZPPorjeukMCBYJxzXAOWT4w9BB7lgW4xxQ8yNS2/JK3aL3JCSPxqJpTWYvLdEFIgjf78Z+bdaV/
Uaglu00uln2vn/+HbHL/5cQf+GcUL2rxKTzJ7HiGsArkR+b05u2u//12Wbx3YOtsR2pX1Jnt43Q+
DlvdSF8Xwf4nDdIv3hSLI3XHSM7Z31R2cx0SiEYTP+qEg0jsOnjxnRW80UsKTD0Ej0jRo0ZrvhuI
n+iSvSNyenOIUv0eXmb9lGHJdae0raSUQqjlDJOyA1+3hgfT99Xi86U7tWm3rTCA8r0B8va39npL
KwLyz6N70FEfchda23FdFu9Rnc4dKkTYC/WIIY2N0+/6gHfW/uXWdJjGRrZiK4JxtNJ8kFn37X5V
ECv82Pvqi32QHv9NxDPz667pLsztMt/C1UeLOLmSofSNVA2ldG/Y3fxeWYOio+bFCi/zMyIylz5T
L5il+0qA+1b5G1aLV0Xq9VC4J/ZZI+HQB9m9W93FciPykU01Jk/qU7Pevvlbhv5qMAX26TMJYPVH
CYajn684gId/Fc0CcLF+cX88MSglGlcpcHQUAaPHVndLh05Ib92pJhT/a0StDGSl/f2QFcK/QeL0
2dGyM+DwoNQ2qtkVL/TMSzO+Jrog+GDIcrEvIjuA/S9v4pIcBBS9L6bgY8riRN0d3KFbUy4bRkT7
foimVPgSmXfyYdawiQo6y4dSfFhNQvag7IaaGRSmbBbZsODDSjwqYvbr5Lb35AVzA23JN5UMt9xg
zhHwpIGA0blJnNJURifTfFdktgdoigFzQiFNw+NsNJrfUV/dhsoo1Y61dVw6pVe8cvJQ8hhTTxXi
bZqLdx2arJiZZK7O2joZSkbUzWlSWygNFp2v+fEXyBUGxDXHNBhS0CcQlxliViZMqxWisldo13G2
1lbqcNJH/2Pcr7yYyJPh5YQ66MyRhd5ByXtyXdKsSKvLO8sFcYHpHSgBygfU9mZ6QD/33D4FMnG7
PxHmoXtRUxZvFMoqyiZ6+hhrGR21flYmxZYzIzKYs+MEyst5cOPovZPTIB1c/XR2y/CXy1Qo7L+o
WyR97UL5Q7FHQoI0PtHY4gasanrOO0/xsG+hAKUImrvHxHVqRK0qb1At86laCb1DWU5CzWST+bNK
TqAt4ToAdG+pjoJ2+Ta1rKwzUVvvCgST9s8m6FKa44BHEfmcseiYJ/87o2RgLY65aLQR6Hu54VMX
4Rzm+GLsuvRIhX/XmHJdv8RK/FnCc6LNoR33TyqkG7x03ty5K4nv9xqA9bFtX6M669GzUryXZyQu
B1VMKnfGVR2Wq7o9eW4WoCImBF7Lv1yJrpsjB7aiHuFBTtt8tOEyl0jzU1bRzDBiEocdoCe7+PPC
Vg76oNf8rkXnH/3wlJPwgLAyzoB+O47Fa2ZML70XR5eqGgVuFfIPDJ1bzV2x1zL00R10kUZSqYIE
N0BWxLTO8B3woxpkMpTSS99Hr0WjGFr0RIxIG1WYtXDw/ZhXQOyuQscP4Ep8Y6jxM7dJdTk/XCK/
EVZecW1X4HrB2ze4cfRS37f+INkj6M4Umx6CqTeQf0fGwGQ7A469mupozZhzUL80CKD4V6FvtCma
qroelEozHx1gTJJVJkez5PXF1EJRIKABhU5CrhrISwNqN/bUE7LCIYpfPgIJ3AGYQvoJS7rvoq6J
zlX7ffZbjUcCGWoXPQ3e9PMCL4j1Z5w6iBPSYMGpYd2kfXlrTv7kumQ+rvDeXJi/Wd2uotJKAiPP
959abK2MpCOC5hDD1PtEUZazZUi2vLAHRHfLT+OUfL62d77Y9a3IHZlnX6UKbefSg0UKIkiwXSFS
P1bY1FWo4zVQT8nZWTTU+hHNiHpNXXLlNFqcP+uDsumVN1yeeuWvXC5QqeWt8AX1BN/Lw0478CEY
zXfBBejSMx/loGaOPF1gGw2ho/KNMhrlmh1/HQG3Qo4Hh5ZRfPU+3VlARVxFMUrrupuWWukCcz1r
bAY4Pp0pWkkcd72fYtx8j96b4+ZfJnsDWfQ+CWdWAOZ4tX8W64C7TWPCy07KlIIyxR45XL3q5bL9
7Pd7wbORN2BwuhiIeJmCcxjO0TSNd+0370x+2gGwhCuTjMKZVY+IF8s4QMFCZg0t0jBX4NLjwf4k
FJtyJCjougyYqSp4PnxlTcLDV2nMoaperuM/Strjbfy2cxO5cpmvE5UEvFTJ+/wnZ+Hqh1gVB9Bm
/nfx0yU8ymV2LHjVhcuVTjIbFkUEAKc1IElUFUnozrhw9keOF6Z2PiqZmESxrRsRYT3VsYZFdM8T
FUR5p06sWDYUbZqv8q/RuhXAR+StqxbrHSgjAYXWtzgbnMiTpXbjYqgC8AFyczffGYa/TWadyilG
rM0zTNyJWFHHbqX6qq7mht48PvQiVCkEiG4GbKEjj0tFVBK36KjQmab9lfQ1/cGGJIU+MhlNjaWF
bVMJyKADYRfZNdbS1tq+uKRMQo82GSS0if8wM3ghpILnouJMvvu3nGCKMCgQAbFjODxXUgue8J0k
CFnO0CwP7+jlOtPSlAL5CRilpwzJ2NY9HgM7gKjwozN3drD1veTMRgBQKKghk73+TRgLqJVq7B/Y
vfCAQhVeCacKerBBwVqE4Lu6/vEdn31j14Uce6Gyo5TlHVjY3Oz9/C3g0NZsP10xYsvUOrDVISwv
X+3muCAOrgPbutGUHNJh6Py/KblYwaNlylc2PSv1nwYH25j8qsoYZRzJkkEyrTh5b0Ygn4QM6cJV
p+flQsKSI3qLp9KIMdqBOXrjRdxmNCBsPjBcoERdu08atTF4bmRo1HJGh7JPf5cxu0aBOhus182A
g94vxyzVXd18jzCGnBkpsrVXlGPBwTNb59jh09CYkk+eE99ACG7GkHivfg8w5mhuVWiWQnx/7f4e
7q6kDKSYbwAOwVxXjyXyfJg+b3PeG4X2gNm+k6YJc5TLsrjrA/4MkOzHOKOaCdeka4VYwBqskpNL
4FxjjmMWB4qopq5wnfKiHUNL/R/XKcOzwsDhCkFwVeKESAahtT6rMIDb8XLGc6T2aShoj089tq4P
KRewkgi15bFtrwf7/DXuQbXF1wbEy2kdQZT89sMV1soh7WrGQJNF6xCrUR1QTVZMhnW1toH8zv6v
Fmh1wb5Jx/+Kj0UnudWnj8xxRmBctNv/+NwUB8h3qPSM3parNZZ0ziPZdxin+t+118FBv5ACyPdS
JWjukotoKmakmz7euTQ0DGNXU7ai5FZ6czO3ejLiOyYmh/JKA17Gglc2ztHRoX46rN3rDFodJ83f
R4WHKqeOG1gRHwtfm+SGKPkJ42UGGlnRlevtywyKX8icDLo/nRHT1/Oz91Eqi9pprxTQrSQUOk2r
ZvYF3oqLoVo73i98e/zy/IhkhwfwimooOXGTH68zS4+2yejrr3cLchGjj/QPgDfGF9G6iMPejGAO
eHZc8U6qnbEdlESFpyPD9ZJryEIIyPOUcb8DGAczuYS97hSJoKCwcd1uWdN47xuWznrzT+JYS1A6
iEWcwf4v4EHcNlDMGLSB3YfR3JoCyhlGbOxEdiYtF4WTyV3kCXK6/H/Ad3dcKVEu0rw6xzWc6N4h
lSWLX400mvq9GJjrce05jXAdN0Byl8NysQbMK3ABKcnpkwTLApe4ReRrHrdzvxE+sWL/MqIt5GcN
TZrwO3hDanQjyuGQDonRwcyCkP8PS59U8etiEbuKOFDlek9GJbYKrPZxxm8RIUU1BctkbocxUL+W
9iMO+IXOFXO06+vNsTSyY08sq8S2pUp6SDMNpfruyFLAZV5JgNGN3y5lEJyps/BC+fur67BvCJPw
a2EL3mE1lNKiYH6Ghd+3AKJk7DWZWRVsdML7SmRxr1oICiRNXOtLOC6S52Y+DLrBESi0q60n8Quo
euP7AiFiE+prDJmn2zDtdxunkDTJIppzDIzyR3XMoiYXilp0L+85DUT9X8xxgBvnmvJR7nCGThod
w9UTEkpr9QUuwbydTKRkXBQqsk8Rz0SvzegGrgNP0e8TJZFH5tqaNx+YReUx327REp730I3lRCqc
tj056muHZprg62qbKMC+GNj6Mbpew7wqDB9WiSqpEVFgm97ODKmyzxULV2CggQoTl2vNDuUNPgOH
abx5aOjSR5zFB/GN93CrNhDagM2vxWoLWxkzLgB2iUlHQC8P0YA3qOU//QuNC7z/e8088dO+tNlO
SS4AUovjnlKQ9VuNgi2FdOEvoBhA9Z6nVhJxunukpB3E9dJV0CwyL61AWf5CZ3oZlrUiOL7oH/u4
NSb0axzXOwzfYy5b4orBcPcWZk1gkd7Kw8FI4WhPSHRPZ2/1ceyk2cT39lY5PvQ5qKjGKqfIF0Ms
jT4QvsHRqxsrc9C8iF0SS/5yai9y6le0GTlqDCGS3/z45wUrrGlnIHym4lX5yeibEJI6CNQfqUpr
E5YzkUAWmXzLQ0WY5eo03Y/NwDZAQZ/5AYcpQugrEsqfQq+0it0xtqeNTy/3meaNgFhxzO+YrcC7
XKuzz2P4ec6R0EsaKaHb3CymCSJ9gH2lz0qau3H7nNCRRDHbxL+AxkLhtub4gkZuTwiqAA7XvON8
joEnG96J7dLOsRmt4J+yFBNCTObW7bYy7a86qK1WcrCpIIunS8cJ7tmZIP5uqqgKRiG/jieNoqv3
YPPXmYr4q9vKld2cXnA2e/EFmhH5onGGqAwF3CamaJXXWlXRxfz0RZe9DXrSAU307QcmeUACjM2I
Hjun9QNtfIctVmu+7lUAgzNnbJYqghWzRx+uSymt23qWOOX86l5xGhbMtZIGxKcCnUCHb3SNKAdN
quaGU9qYu4xF+j68n1LKdw8rlIFEHDyp3ixq/a4zbDGWGRCoJHkAtcZkTg8DsQ4H43FV1QO17gDH
rb/5kFMNuWKFrX/jeH1z80Xe0xTUXICYWkzMTm43o9jzNlvtdJiNVPub/1A9aKeMuetUf5zLILQ7
ES1OJ2whFDsjv/+IjasRXl18HjcnvUAEoZ9HQbVNdyNcBc/0eTUaM36bbDDOuArYAdpcxyQ4W1Xp
aAkBhyiYGXUawSY+PUH4Lt4LROWn8uBLCAoZApy07SMYeHgu1lDv0rjdlf56ldJBsGtqExb+5vS8
1vPYWj9Wp/DUOSAIdLOBC4/gguJwUk4yotqWWaQsDLJprygy7qA55N56H5AZvymVcP6KLEfKTeV1
11BBTaAwWFhwzP1J6U7SASZlAwpXSOFJmp38bgcTYuSQrbAFJzJPHyQB5AnOJ6wQuMXeVU/vw/0P
9W3Z0pCYUy0/PyshQQwS0iZeZ7/DZ7j7pDkF/Ly6NKF2tO0uOt3wB5VM1pG8oj6KeDQTMZGfy+aD
v+UWctzyavTX36kOp2BlYTnfdtepwcFRgQWhbp730ZuwFRAnk4cfeWSLoU5f2TAQlQvie3kqwvXG
8cRbFZc1lxdyj/A0iqwU/wAhV5/ulHwenjtgM82NiU2TpC2RK6crrn5kv3MFaJGe2kLUfk365yy3
jK0LuHpfNJrCKGctvNiy17v+4/TB/tXdm3Fc9mNxgky0mQw1Vj3B6NUxVl5xlHElcjNUns9QX+zn
a1OuPmnRAedit9iVLaH2zgjN/ELUfre7s8mLK3u+ViV6ZOez7ZwytyyiBNIxGBvopb5fvrCfDF07
UpG0pTOvjmtRs+p3HtKWJStG3GPzKjoJRYZZ5FYV2PlE6CuQCQM6NcqwK0iKpZfPO/hFkAGQLbQH
XfFRyX2EU+BXAnyJoGJXLALK3Y1y5eJtc0/mGLsVtDCaJsMcxgsEBiwMf23MbqTvxNqayIHiWpyu
jdIR1ZO1bnxNBtSfl5QBP992bRm2ZwpUMxPoY4sAYhUv7fzOjBWYOXgbKaa7yOE05yRQbia6E12o
GeK84l2avWXdQGp1hzEtorw3YTPhYlm86pfJoPVxQ6qVfU/xyBzGo0gHdqcv5gsM3DCxyKBKiQem
x2V8+ADhu7LUTqK0tFmjaH+eSv94rR+JtC0GXhm9MRbROsL6/WWviqQdj2mxna491JWS+FFZ1v/N
l/ZlTnhrs/ydKq1inXdz4kr7pgW4Fx8aW/MWxifF08ji/D2rxnjMpDK9RIisUi3t3w4Pi0s0WjbS
0IKZuOspzRnoDp/Vz37QFFfzqYLMUUlK6GQGS0fU8QrZgAoyHK02R59FekLxvQX+10sMHa87wBGM
Y1OUeWH6Oj0F3uTQL7FuIXwgPyKfEMw41L3OOx43DauMCVL9vNd6E5CP3qLuohyXSNS0SX7YiQv0
8vN3aQQfdz+PZW0Yzj+NMIm7f7EQEC88k2PsssHWfUHgw/GuMSMNjyYqkw4prvDUeRLmtl5xqPbw
OF/wUJohPNY1tf6YkjeWQXcSxxCY1Vyk+fdcpx0MNV0Bl10dnvPjRqA2DFrKdfVcdIXw89JVbeVp
ijbgT6TAA5SlkZzZQRV76gOwzdYdCM3DTj+km0tlAYdYofFeiLigj6Xgnc0bEWX3nGC5mwsSI1IQ
aBcKfFSXBMcj8Q/gjofCdkqtCs9RbHPPKZ3TDSBHNLb3JkIypI9tEfXo0UrvHBMq/6Ziw0xCPNwv
fM1VxO9fYWIKm+stRD0wVHdQpZd4GcamhK4K7WfyS1QOmYV2eUUfxB+y2Ywi2Rg7p/VPdI6/xaGY
Op2JhdT/D5tIQ0A6SNdG9AD0PBt18iquFFDE4MlPexS2uw7RiUA5YTBC4jiC6DX7NIIHoMSWNYc4
4OU/g1y4eniCCUjtkYO8LG147otn09ZmBwyWNDOnEW3azJLHFw6DkMHjB8MZAF9Ifj2821LK7dDd
9TUZWS5isoB++BN5D3VXm9pS067cez1uuO9wTwjiSjKdZ91flaF9v59ZJArF5i2u1h1ZogbESzOq
XkS7PNr/nUNbaKpPiq7veHpHm6igdC8+7sP9IdqTAUL//TBojhta89SjHNWw6ToifWIsTaveUz2g
COLG99qDVGIDzYn8To7uxkg+SgoF23IfGyDY1XS8D0O22r7RVGpIf/SEmwws4J5nmdpFkQHrE7c0
elibrc6zJgjdWSs0Iw2vZZ3iVCGG2vxDjgi/L+JdZW1K/1GtP9/JreXpg5J2D1booBDUI2P+cLpe
w9La4UbHnTnKFnRq/i7KRG44vRDgpGgzcuXKgCy5fpA87Nsro2GD3wRiz4kFrER239wP1qDqsxb+
uPv+evw/jli+mMjjco/3hX4tgX26sqvl7Wd5sM+agi4GTi3KHXqNrj08YJgh0APd+2LBw5im7me6
7C9GHS7w9un4K2u230UrpcNJHpw+jSt7iadwS/BH0t4nli217+v/ReAnCYP7O5ZqVHjfmgLNtOO7
eT3/z9NZFx2/Wob/+9LvCLqEIpCEhxHmmj9t2e8UcVUYFJpOvmlqIbXPuvL7gyRBXSiE+BjbFQRS
K8HEilrj0rRKNL67ngz+tOplbaWx2GXPHT9vP7rKSDVTiyYqw4OJCDfUOG2/Ft8LKPNIBySikoIr
lWzD+b6XjB+rGuWEKjZ6tUsPW4nP/M2uoLUYWJN/aTkEssUhszNDCz6EYuBhZzzvrmcEmXfykz0A
PlBvj160dt8Y2Vma8xadMCbfEJr677bMvQWtwQedk9uENx4NkjkbJQinYImZzbUNacQm/aDEUs+T
2BkfuBkfFeRPXWGxuxUWlDhJfUqNxeS+Kl8PAC5FQoojvQwR5X459ui263/T5N6w2bryJ/LK10EM
qFmEINNxmR+Lm5AliK4JAYDVNtTCoHsh4AAvDS4koA/k+Lmcdor5se4C6pA93KSWLoQ1f0iUqusD
sF8c10NgZeBgTg/QOji0WEbh8QIvrs2y+xXWR0ZMdgR8ZsIig1+JUKeNkxSUWzmCQUvmKktskTQw
l4dU6zPzd1cOt54mw6V/Bf7U1Jn9wY4xsc2SD5eTjKgglJSgAVIi5UzvFcSkYSzl2XUWLXVdvFYJ
AKVIY/xIWIwdC4ynBukXz2oTgyN/BHlXL29nE2RygdG2FhgW4fwRb/n+GnX6WN+X9nn8fs05AkI6
30Ikr049+840v6FJE4HQADLL+1ri9JtVSAIzlzKF07pAq1jZzqgyUmYPX/z/8BcSBXOY0aglPNQY
Q+1NOIh4FYYRq8yBLSAvdsbIaxmEj51HSZNx2g71jDayGrsUue7zwgcOSuCbxGE+lR/dn2QA8klM
gKHCoB+RY6F/Ufq6GG94T1R94U4Et2p0nooJ8TmolD0JGUetGG4klabBeqELGb89ANKQMKsINZYz
DbsVcgd2hCRfbuNKfLPxm5nJkxD3N6FksW65XwZ3GbtdJleuY2QCqefxy7GlAKGIige1YQa4qXBK
JqcYlK8k/EYMo8/xsvQa94ta70HZIhDUQ11+S5Fl0F3wdHSDtd2RgoR5/5TicYb/U9UkfVGvrYoq
98rgqI44sboFlrIlFsTOUz4MtkdNzHVrFcoKNKdHIisXnMeYeyXWu1ceVqHarmW8JVg/iuiieuN6
iq0qUBuBE6WcmLcEWXDAjDKm3RTmHDPrvD0i9hrfdvAPWXDVG7mGukJbMYXkWk8sl3GSUon8tpw1
kM4Ln8JC24JrDYT7AR1T+se9J8dhOGRN7h5pDfEeM/F7m5wUtJVIsjK9BMx2ZGt2YW8GZlXCHwrc
amebECEoTu8NhQGZF8+DTPs9p/rzikErXwnPeYm9SQ+eb0pelBnPbtPgOvkGUowPljCOX1NpXLvB
SvxvMSCKzIvVzSU1GIf8f6PKY04lZvVmO4TG49yfY9sRAbzcKBq0NWZILiv4iPRNsMKgi/zpJTP/
jd/LWDbfFtI3MiFXucfFqET1y7OafD3d1lW11zpKpu7MNNxmxUZ2BFhuEgT8/IiU9FH7iMY0Hl7q
S9ONvkpMmQkNtqG5RF50yxBfMCdeETyeEO81DTiXsEi/fDjQ5vNNq0Ok0NENW4EXqDNKmCRWp+o5
0mMRYsLiVHaJ/LNlvLj92du9P++lkf9nrhgr7T1Nt4m6OJLURVrMkYzlVQsnvFaTZD5KkZLXvUeQ
VKXMVenP7Mm5CW6e9zCedReWuuG1LsNkN/RWKi/JdZSVbm+z+QAAGuOLa8pzhI+AP08H2qSyF3kZ
RDPkvhyOfzDwaXI9vPnbRGvxc79QsywZzcYkGq0vLz6pRNRI7/Sz65DGP1vADhIn1IckSTuIK7F/
IFYEEQKrcc4JtHNJZSGEgmu49SWgOmV1l9PPYgyqq6L+t75jhTJoyMtZlXLW/iv+A6vTup0g7Tph
jyr+WXLA3HknPA8i3Si1v6NRl6BlLHtKqsMJexKLMRRqnMR3vd8rw6zDuvph+LOuy/G6m8pl4hm/
fzfhG7x1dcGcH7VavCzftq00Psfcs99vZTWOPyLEojpoV7+VaqkWlDyNnuJg2B35YLSvJUdkdwQ0
z+3Cf8RAewEBkrHVuRS4lh4mlTUujehWDKiXwLfy4bolT1w5VH/jzw+hhpFN4w6x3txsxlp5d88E
s0INDNCrzRU4ri/pykvwgU4H59p6aaihPgPJ/n0o3xo5S1LIqoXJmCeqhfsGnUZY/QmOsV1/WuVP
w5qqAPMyAS6Arh/ZhGBW2lLBD03i54+gBfWkbS6fXx9xItIu5OT0+YJfhin2GToZ/XwZyQK+pHBj
oi0DYo5TKg5ZlWbCVsuvvfJW6jnNFnQnxMkw4p0LKPlKLOFviq8hgkoF9wU8lz6f2Is97G8KhH2q
VveE+IbsiKKqVOFStTBAhaM2xyWIWooDrCJsEnhgcMYTKOO8IN1UcdSCovJ6nRDYiPWedtF4YyWf
SecQx6/9FdOxj98nHlDt/ENYN974qDTGro0iDFIcKf094T79yxIPiL4JUT9iKaMgL2qx6W8efnjv
6HJ/ggFgfQcJULpNIHgRyk3ry+EnUFGNPkp8u7T+oe72rkR6SqUQHF/1YK3fX+b3sG33btDhEMNJ
vxavMPnBRiq7NFIDezZn8MQByqcHgE3zImGmckX5F32nKn62Opzx7WBB8U3JIsKrsSSQ672CjM+D
VZjhbwvB0tVj3Loah6zIV52/aj2JyN7+zR47CMLWSBByFazIoFxSLdrm26e3M+RhEKakP5qrvf3/
reuWjOmXVK0Ny2YT6nlHRIyD12RpLYvUOy7aw8NOONCICjeluJp27Zency5swkjK5KlzNHEabJWa
7haoep/QfJZ+MBNXaUCVwswR7PKLt6nyyTqIj7yWv2mqAMHFuSuJ+WQxpyyZ6ctO3VaRhdOjaDdS
RriwQsUR48GWW1nGpSdXwpz2G+BhAtx1OQAzGz6vPPoRQnb/lqEGEBf/jFmmZ7rziXKjcdE/94YI
zZoT4jvoFh0Xnwoj07w1jNyZXLoBztWtO4CREwCJvk/ePOPoM5S3fWNmiPSec6KzKlAq0VRHgF9i
t4Swoy1EF2hh3xZA9H9JxTKdEQwyeFH/2VJ++8nSgStmGTyvUBuyknghWglvWBdrX1lHvaAObVHI
lB96mCwW8rOquhy6W38K+hvGKkNCjOKmOK8cjD6/AFNGPHXqdCWuu6oun7Y7PjwXHGgaiAOWTeJ0
eQ3xhdF9xjTtKPgaRj52C7nNb42klrSZqqXe6ureYrqitcID0WVJQ8IYaXarPqvkc5etgqmkiiQU
EwG96U1vQhiF25ClkSC5xrniS6dWnCDCgNPh01MIkUiey7qyl063XyuIkOcqQKdgsPx5t/ZUV0aY
E4irsPeEHLZJfNJYHHiqfh5zqb0s58DDCOUsJsgifJNkPeueJwhKYJd/2jC6IOZSKvVtQytweygt
mja1q1+e6sf79zoOazySs16Rumr7zHbxNdHAjVKPmeY3dvqX+EZzJ2cLaaQlGnqQSD5aV5q+1mKM
WfX+E2+pQk95+/kVFLGVPYdzYbCuv+SOQOrPz4peMRucCyHtmkNCH/vfHMD1gnQ52Av7nM7xFvQt
cqAaG1o3yAttmNAAvhPRT6i0LX/bMRgI3xRPlf56JZSuBdCgiB0ciAvEsNwhvbY/YPuy+Np1DT9k
r33GomeqQCQZKcjILh/jirXQuYtz2X4DLvoxGsn3rXV+BrmnGW9wqkOQpxtqQHH+ca4xaLhOOAUy
7NdmH/Q3s1XtrwY13gWn50dZs5Lje1xqtX6M0cwuk+ydX8YbvHQzzObj/h3/tbY6zmu5umfaqRkx
dXQegrEJvW/Qltue9aHp4Cez5FDcKNm+CRAsHxBODPULxaKl5UQvLBjiDr+X3nBla3g3Nhj61HeY
taKSTPJfCmRyYLkwGJwzeOXpjEcJMaYFV6s4TbfuBpgHVkmT8/PLc3tGHtkwKV1BpnJYAvwUD98E
t8xyAyZDLcKUR3oA2WiDxXgnkxPyig6LJAFVBR3cgkO5H7fj6N0XLrC1Wjw8G6DMVnODV7+G0fdi
At/2QyY8yI2vbg5JpB7GECM8C+RQwXCv9102t/V+l0Pn18F2sgtu3o3jZ4pyIF8sDsLY4quEaWOa
ZFk+B27JJQFtUO0kSseR+BEgL3+JKGyAkLVbCyFhuPnB7GvDMMM+uTKOV5XHZPqvl3nD3eI779fm
O7aIMFj63AIWkY4d3eZVA60c18FVSZuuAut3YrG9A00H9rRrMjPByPPin+cCWSbSM708YBeQRR1s
zMdYpNEYMUmAe5bWsocClziWBBMyex9KGzCLpMWyX5TKpuBSR15SW1A/hmVoqpo8tm7/UILW7hzg
vws2WdMYgMQ+cezpD5PxkKnArC1dIqQUCWwczeLJ+k3tNjslOf9iKsV1gQ3x8r4KaC7hYKyZK5ks
SNsK/eF+HyHIrxkxhQc7gGYWoASyGr5kRhbIqcrcDuUqY1wmBH7YIEIsyUhYQXM5n2PAKUFn6nCX
et+HiCXChqtLm218IZWgf1X3uQd6MiXUvLqWx7by63pWiig3pdXmwNx1tHboT3D4BnVeIsXoavp/
Q2zKNWi/ddk0Qbc5y5qF4oJEOPzVlbSa4yFiGbDhILLZ7hrUGxgAErfTLN84MiPx1iDWF9X2DsQz
+Eso4QttZ/P8+MloAXHo81Qbsjh2ZYXYKHHh5pWqLGmyt+JlZhK+vnX+jbgOUuLwyB+By3wCXlQk
Czanc3WWe9j2s3UZ5drqCqNI5jhEh3Xdc+kRavGSDctkpqHt7zp7U1BSHwPeMIjakymvQc7xZkoB
uboIqu+ifes/OclJpqS+BnAhtz2ezJb5WvfXT8h+Tb+Eix7+Ui7lWUKVLGNgI9OqzFJrr7rs1CV2
kuqn6fwF0e+hgB8aTn+s1dyqBrWoOAeZo4Ie3u+S3hrFVJr/rDUplZ1m3BdWwUDLtFO8jOGDlMQu
MHqzNVp0aVm1JHdbu0XbHM7FQZv1Q4S4yasdrehdDqTzoEDUdvw/0/pziJ2i4sxD9K59lH4hltFp
zCwSqunF3rT5bTh5LzsNbJJ6GMLlJkF/IKbny+nSaINfNoJ9fUanWaRP6GA/eXfQe6I6DqlgY8Qu
cV4IkfQ0uKiKaM54aGtG16is1+HYQOly6sHbAIjcvVW6W+yV2n4xX9It6AtiVtGSGx3yCH2Lvlra
TEMoktKpIAbt3sOksNMdAmgdqKaMds/bbpJliprgsTnhBpMEnfj0S+r2/3mWqgo8pMSvdFCHVaCq
8GVjT2APvwEt+TUH32Jq8TdP5X5qZnhJzgug9ou6RdHqoMRmD1xd0XRcAIVv7oYhhq34vNIhoGAH
lZQFIzJgchmzVBHROBbDsxOyowFPceRYGgVJY2w7x430wh/S80OzWowZRcaHFBKoNtQ2uLwJFTo/
L92ZxUeLHTpLsjdwZGpF6/xu6mCb1ed1USC2C//u/AN2pYXkZrJJQweATa3LQfjp9DEd0LD43KFg
nncUI/qk0+ho+XYexC9mnnMF7wwVzRcpXcH5SZ234qCK8zL2Izto1dKbp20bf+I68FpAvs5+K53C
TEG+oizgxw0ZZSqTe3ZYH+qvuntSwPRZd/MZxJxHQukMClLiv9yhvqiM6H2xzhTPMoBGkkHWZ5ho
RyVTnWyM0j7Yi1isLjdXZBqNMhox49xLqSv0BBU4NT1bi1EaSMuq4Zvr9oYVZr6/XfY8nVTWV7aG
BrMluAzCG6UEsICMpt/SqbHtcmsWslL7sNWUyUwRtAYzt9wBXxzgJzE4BoLQZIzAvuk91TFjwYq/
ay0dYPk4y42yL3swzKEcZbzEEJSTyHDfwe+RC/eNvX/qeKuM3Hz/BeBte7hdtx9PbcezDKHXZkNb
G8AQ8eRq9Ha1zjN54cGgnEQ2TdPmG9J8Sjc8IF+vDoFV3QTHIg/kOaD9zv0Ktz1leuFX4/AwgIVh
NuWD3qR8MzvFmhU26inU96+kbkvBDAYxk+GdCPLUB0uEgSEk1S6QVJybVL0+RMiqsJqkaHX6mha5
X2Da/tY1RFqTjlEFx2uPqCZoT2gqJy2p95frhN4VClc634lh1X7XNezsqdvjw2PBIm7VZZQGSxa3
VYOhdzx11YixLnY34RaXxEObr0//RP3WKOgZB5tmVO587p0Q9qa/GRvbrHywMig8ZR9apc+JtK/4
E4jn5WcBg9xoyHwYMNt+EJaY8rueRRTf6oRaNsYa3F6UwYPTjXNs3XKFJF3EEEt13vjGQPH7COie
4g3KSzvFabWnkZPJEliKHhiqz7UH4UgUAB1NaG2LCajWOXkoPdmLERi4xQ15AR/eVCi49IasBZid
/9UUZHHr3mDhmnZqRES44j5L5dnqq6i4D/guuiFIKeWZSKJBRun0CZPQEFR+kjy9x1nmNygwQN75
X9jxeZ0nnLTJxR6zHCW30tQGC8Kmdm1p7tJUXMMijuK3o/UcAT4WVqXKzs5bJKs1aMfuUHAKeclp
jBmMow8DEQ0Vwu/XeADj6tg8pnbD+5VOgIza5IoEVV96bz3+0/LIhKheo61wOpbBwv//naOXzhDB
zFh2qbPn4w0fVIRf1gXmmgg9R4VsJL+0e6+2fBfuPJTXtRn0p03uDdLoMxkMEK0je2TrtXWMxLx8
kkTL5rf2wTNShTHJqmye4iOOrRZQdlrJgw6MR0RLjJCdA8xTcEDiiobCI4WRtUiQpGgh3IlTAS7x
i3kMVlwGpZLmLqAqBjGCR4fOguwv8OYZEWvYtqZc/2ULMkwRaTbWgsIis8sEAnXH6SxPCiVlbbww
yyZrmEgVB1YWdE4ouc6CdPjN4Vtr6Zy99BFq7n12JUTt3JXDjFWKCbfWcxcwF27v/yZR1JQTxj27
Kp52AP8YNPD5exw0Pv7c42stRPExVXhhuBO/KUl8OuPf6dplJ5RaXVD7TNTcLiBW5MtosPZ1TEyg
l4QNsYp/7GFMt1VaxzkxHRLMJ9KxXidbdqP3Nz1t/AxzlEAy3KyoysuACbOM6TB1KTQ0k53h4/pq
m2yiae9jZLiXx74eWA9kp8/PZ5AM77NxVej1SxGFAicO31Tc1B/BLOpWhRY+4s2z1e3O6yL+8nvL
gPa+3Vv/+YiZEnm8LcoNA3WF65VVD4WN0aNwty9W5yuMCJDpkVohuSQndBEiTlSPGncmFsVPC+2l
IEou7/FMb+FBLGTkuIMlwQ3f2FwGxYBFdnKTGzh5fxF0qODm69Alz4d6ZP+Xc4A+97eQGOQ3jkL3
4riHkoKc/bIgMm/JX67iNOxpAUwVCOnDvHhPEQRH7zcySeBR67Im08cdOAsiXw7qZPr2MuyD1xhQ
byxemw5cqXse4+PfuT4rzFHdgnhKpdE0d3nBY184nu54LD01CWaxON3ZnldiKSmsGc2FU+F+wdQP
Uv58E4g6ieblbHSSvX0iS52yAQiEUl1x9hWKMJQTGg0qSy/VO+Ol16d5yVNRoA78BnrA5vQtJfzZ
7Me6DnqIxvLgGT/LeptEZiJnSC1KwN/wHzAotgu7P805/zdJlkGv+gPO3zSyhlNJXbDm038KfTza
y6+jSVYI6Ln6mRebhFGkuPVYjHQBZGIB/jOfFyFLpj5gy3v2UaOkKIN89B8Nxvn6Rr5CLDL9UwY6
f2l5Xi2M9LqZhjeg8f/SxC2Db5o6TjAYM8a+vQHeefi62o78oT1WB2jRy1TLefGzWHgkXGQ1h18r
QtFTXYb3HteQmkV7sed2t+MnAOKzh0+/9JvfHRxn6RUYeSfsBSF14nEv2ArChORQSrn2Be6004P1
n7qjUCetNOvOM8rZl5JVIylvYU2BuEZii5VihyluYmgMz8k7bomivl8of6f3vh1qJVyC5ONWTopK
5rtNbk1nV7Ursj4KAluaQXxE+G203d/Pt1wMIzQbM+XStjqABLpPfTerZaDZFA8mEgZCgJqQ3W6a
nhxQzSt+13BVEHcIIf35XhXvhIcrW6HciY1jxxw3iIv+/vJLnty8mCeQml+0r4OhMnwvXvaJfqIQ
lT++c6mlPEmYhN7JWOZboZowQ1AcR21XgKewR9nUNIz83Mc7bkWaEDZYumMysZxmjTRVjoq/x0Aa
zRdfJTDLltdlV/06RPA48fJJlWVn2TIahwtXtM1ffurOVm5F3P4umvlMY+pPsvRsKsmyRH8tpseE
xdvrSOIai0gLjfYMaTH1andhnh50CaMaAH/rmJTicnOweiJp6Vtk9RH8B8xT1+1MFdR6OQaYOlyh
jk+kaWl6vM613RUozFt7r7kKpGpDNfgLZauLta5nbcLuLk1/FRtFBi1OCL+n/mWgcqjVC2WiU8CH
xsOkKhV/0Fv8etIGlexujDvHirTi9ycJ1b+6SO8L6xmJnKdxkOhpnH87EEsT2RWg3PqOzxyYvO62
mG2QTVUkrhhd70vV+k4SXC3DNj+fD2qhm++i5hLYe8moHDDgnXREyAq02Dd12IksvgFPALbkObeP
VgvN7xcanK6ZLYv7RYh4WFcT6sw47XyhzDIEXP6LkTCr3tiX0c9/kAbfbYpL29PqV4EB+2ny70ks
KVkhGv09HOer6VqdPt6AEuEQ5WIfgaqPQZuB6pJ5Pk40ae9xmvXosDeyvl1vkKtGnNyjr8RQ+qEi
Q/mqjvd90JiX3LhCqn2T7rO1E+ojuSm1/TbztWkXfIip5Uqd0ChKPXXT3ZEeXTeH/i1xhrB39fE4
KnAqwugDZl4vo754BbneTPoeTCD0tDbS7L7EyJQZ5nAbff6vZFhjqO8dSjrnUChRDhR2I6wFf3mo
8z16VfviqdMgy1aBoq2woLFHD98aQRD+DB3fl91uMvNu/NgZtUdRh89rb2r+PFr2kRKOEcPWppre
GB/TtSiGsMmBIFhH32v1ddndr/f1rFjll1J2+soRa3lZ2/ljmyNKWVV+qEFHiAnjvYeNVOTgpAqU
l7FXudd0CGIxwvljG2E0Zsw5Td2bYlTWv8GY5+LEu+XxfBTbKwC9wKGw0nkC+Y245W0SG+SZKLTy
yVoQhe9OT0+jOuxz+Qq5FgfKXPyBeTk2l9EQEbOSgb7vlfzBBL0x4x/bAy02jZOxvmjI7VCsF6dY
VvrjdxQeu1BtfCmE7MroiF2XlcXC9yqZbtJKg4RJyZJB0pW8AvTSe9KDO88+xpypZsRP//Y9dmOn
m6KxBp4SaFQeThvDeCLtXdQwQoOS9/xGJ3Fh2IpPP4D6zxLXi3hsL2e8qJzr9V05ycNPw83T/Dhf
4DiZQtNJSL3pD9F330zDVrb88tqzdK8xddG7jT8CgLA8+m2itIZLLMWdnIiTC5okx0gamqE3xbqq
G2PHYZ2+q3QVhUaLCHxF3eXvFBN+1c/SsZXo9g+9n4w8qLLeqCBuD7EWROWac5slYXcTsmmqJeBq
zanWIIFt10BLlcnrfXpXsF/M9RdNFZ/EvPbcbrpzuHXSf1/cW+/d8fE5BOVfZYO/V1tNxXG8qMOr
mMX77e7Klg2dqWMyy2qmfxCDyFxAygGO40neemCFXmmkQFd2QJnoHGaIQQ5ERBkHwa9lH3fD9ljw
C/vm2IYqbIojyY3ka+NxjdFwXR0EdK4FuKlOfMELQfmZLS9mu8NO2nA0s6RW0tT9bWn0kWg1Hx6y
WzjGqmo5tPh1Z/qQAeS+VBtHYvs2APsbfT1R4xLoNB8gK88C+ElZb65CdNuurRA+nu9gPc9wGVAR
vZp6pzwuzgAPnRyfGVW/Jvs8nh+BssYrey3w+dtYZD6c+wurH/4h1VgTP3k7fjqO8w1UwCI6KV9/
xzcMeGTIbJ1YJDSCmUKC3QBOa4mVppbgEo9s9J0jdyCGWwdH75F54cF2RyPf6qP6TlQDD51A4bSR
B5ii1M/XoaQ/Opl5PmpfaNM2m95Nn7qiLF5YCBQK/OEydvR/ioZ6n2552NBUWWcDR9oRUOJkMdZW
z32+SqMpJkE0cu+s8VYk5hkb+El3P1F/7mQO/Zypelb8Ewj3ZFtrQNj6H97BkfxWyqECmCo8FqhW
mvL5p5JGGDQoVdGx+5kNMM6d9rfDNSqkaewjkNlN0YlrwLlboJO/na7cjYilGw9pIiW47zS/UcGh
IGRFhAqqEHPgNSoLvC5MgBjjaAbNTk7FDL3BFoIK1D9KJHRzLyeqrZ89bvkts48VjUohPvib/uMb
OhXKF0smh69vV3vn5NP2JLM+FFCP2ydZUD2FOX72lxMdmwFmqquX5QBriQRBdMWJjU0Pls+UIU1W
Wa66aRpfi9lPewOIoEdbgrPbihchsMWMT/tV9TZsduIWFGoWcPqQCu/y+k0zdAoY/FtWHFHkwO87
Gz1vw3w6zueDaOZQH4zzwSelixzXjAAeZSzxIRGOZ2ndHFTtbZqoPh29pZz2WTetDyOWOcmieD07
F1n/eu5NL24OCpFdHpi+F5cJE2FdKOlOn05C9Gw4aRleWTNT3p9M+2EDqbDwRZtR1ja9ZsocMxlW
sh3fExPL4JMJynNd4i3f2F91SWS/II53PlyqmbU7xIry8lkRiIgHSFH7SZSG7GyEGxMlvWw7Jmbq
KZMgKzJqWYEtmGSvqVGai3Nu3Jq0nMJg24aXT4Na89dqOJO5vzWyQvdeWN0FcStfxzxZAc59U72u
2APOfDeoHMH+z9u5oZbY/I1OqrvEISJEe7Ic5B1fC421FbeEkyWkPlc3PNCNZHuf7s47LtJpjT5V
8vLjn9oylKv+aGcMvWCRUkm5509MY7bbO7QAEZ7quDlLWV4hdnErBPGnxp+Nz7dpvChInHqz4/yd
J3+RlXvzMd7c4+magcXdOAGHYZ5WQh9nwevxTOBy6ic8oQQ6VaYJJhV9LOeI6kwV6UP0R98Lt3hm
lzaGoRjuLn9rPzsjGPuQYSpsvFrHJlTj4/pCYRvl5dzZ8XeTFTQFvE8rPxFv0N/d6ztmlzVE5Wik
8VwGcPccUCtQdwSfLlHPl/xz5AabGvWyiR+W3xQuhod75FsJ57S5YoEbkpoUy/rchh3A+nFTWxIk
KX1HAI39ZkgEJSoqglW0OLZ3r5D6DPjvE6wdVlIfQmJPOrEa9thB/wr0ayAM/90psRCbO3x1ilB7
kt1AA910hfYVzv89VEJOUUaoERmi4MOjwniaQ8Ni3h7up9nzToZC/CeVnDebXbdnwDeArsptteUr
PQMFw0sgQUoyjG2gFKF+RP+9d9k2bw5NJyC7HErdIe2vOjVbLlLaxB0BLEPEUDatD9P0cDipDcL/
Rq4mLQZ1NPf7B5u7Xd/foKGcgyzYhwUanfk+8JxrHCf27utwPnB1CoByW0JnC0YSSE16JjUuSUSm
LKQapOM+214u8yy76nOzh2xOzV66f/gmj4+Ynv142aM0vixpF9HePPJZEdXvzuL/SEEloLBA0U1Q
IS49D9xaxN6Db5Z+38NZ+GL2El+xY+vB1kl9fFuRps3xlxO4ijeOFW3ZQNMjCL5KXVtKOicYFA9v
N2ChT7ADSJ32QIJj9Fe9ABOnL2Gk0p+wqppcjcXlCf+CXv16McZhboAXlzZgna78pkbUImJkyR/2
1OINDHSiMEu2OeU7R8n0DVjO4ybX77VEuuYA6DSBeIEbR418fI9P8aAJbeWyKO6iRlAEkpMVhGAF
q3CFe8su2gsTWe5FHSlrv6gJJSYeY+U40WAjPIuqEgfwRPVmwjCxiKDNdv4Sf5Arrcdhj/HnM/vv
o6sFMOuxpj1e2EGm2prE35HaLcq05hW5/ct54ecTCP8W6QVuPaVbYw24jqKgoipOgKDJahrqvHKV
knRC+r0Q8HX1PfJY2IniudaQQqr5gtoNao9tG8pJiLQgzgKGKJ2wOVOPhNresPzVD40eGjxJ36oa
rv8OPFuYRmuyI2ICTDUIWzEZ8z3vgpz8lk0NRVhi0KdlHmlUA4iwIrzLgdEBieqOKX1YzFjiF7MX
utIJ8FVguCTllwPymha9aYcpfTreS/hEiCQ/YvkriKvDQFv+nJgtLOnD8QNjJ3O/QsSn0HzuQPpp
B6FPSQ5VsmGDClZJQE/tU+q0G5uA5kcUiI7dUTrFpgQtx5fxBer30tfxa7atm3CS3DfIIa071+o3
eyGtELLHckG0wEjLHAzHGr+mbTY1LRfJHEP6MzLdbslzLNPq/FiPxt9cnKsnauvJabMJc5AzKiyj
RpC5Ex4f6UZWNiFy8ISw6KEJD2x4XTu3QMUXXMAGmtqXnpc1AjgzOiZRQGCwX3sY2KkoXSLRdkd4
djLL56Hb5J/2svC2fkPOtV6+HmEy7fwapTwQdGLd1/cvM5MzMXoxsgggtuAI/ErjjqU04cBrwg+R
Iyp5XHFXlEuo89qOLoKbSydbs5wF+/Sdb2fd9LUwXQ2O1myEN1qGEd7wfjbFE4adqW4GFCqBXV9/
KgRhYhqXXJx5TIGjURgT2HG35tRz7D6jGJ+dKpIAPYJJTisyuI04A6FwJZJRmXcEYe9Ow8B4ZdMf
X9151jfl3zorArDWrhyg40M8XJhDteqXhSKfW/1Ekbx9UPCRRriV9JTXz9dIRdXfP73vSYW5YtQ3
ZnsNW/p6Vsar/ft24u1sip6+f6HkpK2AnEiY7nGM00H8+Sp8mQp30pujiUus7F5hDr8rRbFJoVkf
X7uVOIAmLnAfVtwjIvSRj6RTsb7H3waRBpJJ7NbepMfTPEhIs24YAfr/uqYwRyO38qkF/HbbQyA2
Azv1Az94+xdyjR085Ir/j7K5Ul/1R5hLtjMdeChpSo9eUnyytNj8iMse4riEdStR3TekF9P2wBbq
LIQDEnkV3UdV5RoLA36mjC6QUjdbEJ2XVOIrX9xagVJao/JJ0SH9Kah2sg0g+9OfJuLvAQnRqD7m
TRigwYO7NOelVnCgdRZknBUPtAuwUbgIsPLq0aeqSFEgnffYVZj7cURkLbHL6zy57p4IjxQtHdvo
w/GMYDiP2kYQaWVsDh4Uh+4lSHvO+vaUB8/3n4u/85La+XIGnLDvHTdUaQll/Qtv5EIXV+2bbzmO
DjlbSHsZTBBT+2AG1TtjI7rGGv1KV4FoK9WXi+q9QxSJ4zvttTrTagARuUdf1p93bH4E/LRjtdou
FXD5Dwr/Q0Aj2Sv3BupwiwG/uZzPh04T6I8sqcKLsqZQ81Hc0v3E0hANWob+o8rLex52qEhohQFe
9zVIZSoTxyuTybqxdojw9GT88JDMa6kHk3WP4HSik8Ep+inJrC4hWgejPOFAtE5EUWgXC19i1IS7
ocwq662jqbJtnPuRCYGhmk/+8+yk1zlZsnSLsL48atWCoHi0DAiJIQspHuTHJK35JQ0XKHtMHV1A
p09Ms5nRdAQ0rx9T0ybcqakGJZudrbtaeVwdxCADjvbFUwqrGFLnsgcR6RoDG+CAEngmaBxmBLN7
NucqJjBR++wTMvKAIfUw86HFizTpL08aCZmnxryBQueGn2GXGMfJHhlexXTjychFPAvB8oluSk0l
WV3uNGQ3jDTI2yi43CIDl2Ecca6Bgdui0H5FiZgZojwreaNQLdG/saDu/AJvtU2hGqTInoDCUx/c
xoIYEaJlbsd8SG61D+3YnsZwCHntuaUFfWGRRHkrmt7Ida5ML0jiJDlxPU2pxbY8WbHbbuJH78pe
y4kepfRvAH4uDrRGAvIl7wa1Hm8lwC0Lddg4tqHjq0YsR+4f2TIAzk6VInuCcyPQlbe4aa+gMopX
5tikCDgfuHUPi/WKUYhVi7jrWVsTYq32+8caxRa+4Z93r27yhsanOUUNzCHBGHyTvhC9KfI3ILPw
/nZ6J7mAQzkzJwk5B6jwIpKgcnqVQ9VGYZmB2o2m20Qk2b6j9jrBHSsJ+TvIwvUPnZMC3YzEfgR9
KxzXh1B+ffaNLxfrJ/jc+z+Nge6QoICgls1YbQ4IHjfJ8jq3UVbmv18EyzJ9NEYrp0K1piYVkiZs
PVFWzljIL4TB5Y/2T6pfQAv8R/N0625X26srl/h30AypzJX9YHj5OxhdG86GSo27baUqgw6HsRgv
E27JBAS5ZRSa1HTHQ1z1LAIls/6pvO8ZgijUIB8XcoJTZzpyrLb9bs9WannEn+SHAATslXJ6pqmK
VPd9ph3cTOME2qtRQSI9bAgmeWmb/5Hp7c9HUZYmeCxijHWm8pzZlIvcZLt/WPpbC2PJ0guyzjcO
gQ3dKdjkxHy7X4sKZ5EHlAfSovDZJ6vIFUXmOjzPDCOQsqODj9ROcc9GGg2aGnZG5VPYK4hiLTl1
hW9RhMy6MXoCT93tNaN0qMWpqg5YIXiRr99xLs3Hxgbaq51g/CU2gMGUeQ39tM2bk081KTsmto4A
IH65BZdADL75sUC094n8Zv4DRZDtPmSt7MD1By+uMPDTwTKcfZaOvx6eqpdtbOPfc1cKXjhCjrno
4P8CpI19VMlSt1SWtjPzcGqHEK3wS94mL6jdXoJ/fZz9kq3p8Xw32X/QA4RyjVTQww6kKRSlFPbl
XTaV8wCtH3SoCow4WdsalSym1/X3HQQm9UfoorGTI9T4vmJRNKQQHXDNYj9+q78GV71mgz9ShJRV
FBAtOcFm5IthheBzsjURPD/90gmi7IwiReMbqjyP0HeajwCxTyYm9ec2bIOC/t7+V7zTM/nk/r8m
WScMlI6EtG8t9SlD85mphLvJLU9DIqK8tKBAPS1mz7tgUh1NVBr8Z3hOqUH7rsseVe2MHE0KSTy0
vAQ7f3XyuXKJ9rKcRJQH6VHhPQhPkuCRannIzQD33HlwhnskKPijQcFuYDHh53EmRloJ99IHODXT
9qr/GyGczNqWbMnXrFnUVGHTeuWRoE0F5OGDt5ijsGaXOFZzLzhk5kddqXjcFcTu7aitgT9zkFIE
ZFzCpolluxaE9xj6v1F7s/NnO3sZQAguuYn7q3c6PtWIHizSL8VfcognNLqDfFtg4c0a7QU4FUtf
59CbBM0pLKRYiVW+gf/+4cOaQ7mSSZL89l0EjPT4AYSY4asD7/8SpYGc9V8KlSiUx5rKR3lmYmHm
D1kgXuYaEzezIxoPwV/Rsm924uhq+yqE4JphkOCN+rwyEyhPRNSoCJSbjwUtMsvd4O1ovG0BJrB4
cY95ku9cjGAvAAMvQdD3jApwaYNuW2oBdnn6Geli6zmhtOgVVfEql4za5Jx6JlYT/piIPv6jT4Qp
2k9npHTjOFogCA+kO/ZmIC0Dio3kKyT9/deIAgVfKgzrosNBFhFB1ho2aVqeORCevhvHre3AV5Ty
M+tUIOds0ppXh6eaKkk2nSmcO82IZbwhhsAmop+FC1Re54jaW+SVokZexuY399jV85zcyunJxOuY
w9D31LR1s2/XLN4B2OY+wVRTDAR5bVsH6LqZwK7/P8QsUtsoCQAek/5sB5AtmERMEK6H9pueenTH
PIM9j8UDUcWVwFCQdS0Xpzzy6bR0wmT2pD8zYQqZjOPlzIbi5Jyvc41bf3LnEUrIUkuXeUHLybqy
4HCQ4s8nMXwpA/sIMl2juAfitlenTvyVqdIFOxGqVZ801i/dTXMjMQvquYIfmvnD5wGUpAOuO5Fr
XIk3BP8Cs+mCNsh0DNX/CsjASCmZS22ICq6XHQwUKjWuqe8m+YmENBeA2PvloBYpIATm40U0QmJh
QCLFjs2NY70RVIpD4L2jXr8rNGvk+wE9Ju5KPPtfbZPLhfrs6+tOussf7K+MjhzM2lF+77DQRwCP
Iaw2SjbB7ZQNnlERucdKRsoFOrDuYoF9WJvVrfbXXjc5GkofsSU0T6gdurT4P3NwoUc4lVPTeUne
HVYupQk/aC3BJeakWmbGcp+2NXsYP1XdchY1JKhe6psTYu7/W69ZXdnbf6rw4LpP27s2MeK+JPnZ
88Dv32+oML5VMpIIPY+jy2RxNjTwkv/Ghrb+gH+7Xp76WvJxkHZ2bOis3Oqx1Gjo13uG31FHSsKv
67+GR5SOloOBz6Ga32mKtAPe4QUgMtVwROOCjTRBDtIKVGOeuXujSWjnBPOiwJNWanc2fdXHEslT
82VOM/U+73V4a9/G8gSpse5kl4hP6VQuhOSEyOrBMQtEqAfcQMkZlFxIVxJypv1PX6NorDtUhTsc
K9WIlZ0Nu2b+7/ZM5DyQ03DJGHrl0K6653Tb8/qp3FmFTrycyywM+XPUE26erd32MiAE0Y605Mxg
7IKvx088jov+CbjjWAtB50qdORHNGibtET/RIbC/qhv703p8VghlyLbkCJq4XnN8Q+T7Zb3hNsFM
/gos0ardusG5nxzh399W4Lr3DHXvWBtKMxYoEr5gcDh9ryTNQU5BBisf8mnBRhcPkXmvwrmR9zp7
ZS6CV2gmB+V59Qhty2BczvJAAw6LyP/FFRxvW74awDcu+Bkcb+SBrPVbDs3bLTwuHZCToaSGydMy
/N1xjr+e/z39pY2EtjY3Mtk6hVIqmhht94/vhfP2bkDBUPCmX4aq5HBMF5bZwQiZRTyH/GiyW3Dv
u0qDLobbojjbaXNt5Eoz2b3USv3FnNDfNgMmXiOW2wzEgPwM0k2B3DEwYllXcvXND8GQDCTLjreL
PO5+8QexFfYhCtYw3MWsQ8605g2g8nTq3Kq1ASYolH+xEUdX3ApRYU0AVtx+NwxXmhOInNOS9IxR
VCVrNOIi92Jgl9H3Ow7LjQEkN2KfSgbsMWB2pKUtNQY8h860nfcSzVStS8jcy/hNGZAMJsTGlbhL
XhNGdond/EY16j5te0K3JrUmm9UOA+04G+rpcwlQXNfMahk3KFY1vj5TDZLNrPyGEqoWiXltkSMI
AR/q2k1hmNnCUdbar/43Ba/iktYrT82lvpztb7Wbl1th88RwrLwyru8tzYYz0ccHYFAXTPLIUmC+
aMw24C0bdfNCCFOMTJwdaFJE/OUuaJdZ4fmc6FaE2/69nBUp16fD8FFwSjZnU/fR8zGeodPYik9L
igpWfS2uAA65WagTTHaQnQWakFvWVllPc4UPb+7E+4q2xENK+k6Wjdc6saUgVtQm7c8GG+rd23FG
vgaeRPiyZuMtasOL+OLmlprq9YVTs5PV6y1A+BHzQRDtTPttTCNJ3sceXItJP7XS1Iw682wdpaUW
hNhalBfStYgNt3Lo6L/3bYrmYWdiaijj+Z8bHVjaFMbakgxtpp/Z6kt+rCsn8lt9JyU5fQiS+6Tl
ZMAXY5ojbAvfYILYIT1q4HzzTwmF0Bdp70xo+CO/xlyUggjiEekz/vQUu4vhFi3158jSoDuZDoii
//mlPNcew2IO9bQiMRrZXTxArMzVkTayklUmD/bM915EgU+wlaGhVs1YKlOn5pkD3+wQ7750LE62
9Nq65NanHEqXykrQB7c/Ka+UFu0cCaENqyOdn4MmGl+hkkVwpqijU7PYj+44U1hvb//Z8C6nAak6
1du1QdxrDHN8XN0oBsTPgZqRMGgDLU632nttoGZ653+to6rgBXqAbiKgvOtJmVHc1UCwP/ugBqVF
Pdy2uzkAdmp4qmOw8BjFBhy4HHMf5uJcARibIqv78LNI5aznWDShOPpRNTxmR8x99YsxGTSCObOS
4hU902uS21siaEtLS1XZQaIBMjatSHjH65auIjUSHyDZUhZ+25eg80czVSR5N/TZSHRKxyAJ0gxz
0yh6/5RDAKxy3x8i5b/dOHDEYqaC/9uErcFLyQsEt2Hp07VsPtTVxQOQB5HK+C8dIGR2RmoN1Ttw
a1n50WSfVr9xE8crJOoEViimUjgX4SxyBstNyMkkcrHc2h5YSYCYzhREEodRMJDFdvEaU2F6D1Gu
q2ftS7OfIOgGehlfKtcurl6RwKYxD6JAn28IpK7X1WWU0qLUznB56O3/Vx2PgCt6+CAiFknPX7oc
0gK2RiIdmNZ1nE4hTmDRkVfLApguNXsg+3gu+gCmmf6vTG8kiggPqKmRvUiqPK1P+vYXy1d4zBsC
2KGyYGJza5/JgrFuGa9wKLS7PArHMsCYTXvPUZN1R6IXqvht663ybHpI9mrWPztzjbmGqwU9GIU9
V+pWuyMoNKvTv7Tf0m0NBtcweila46ZyAeVRg4VFjAub0s0hBLRWSmezeoLXQ41+Hg2H4dfwSFdC
fYz4s/njpzJfI5QmJjvZaRKunP4GePcotvfXH1ALDv5hEYiQjxC/zvqNK3/EYIQLdW3GpqGF3zXH
7EHMhAzafxwTEcHEgZnKCHbOxW/2tyWxlS7TBNduL4VLbuhMooOSR/q595ozQxD3l7jCA/5MPurT
ev3lD9an6tzTAJ7yF967B2q8xMGCxW5WsWax6PfFtKtEmB/atyrbNrA2DmhWT+TXNZIsWbBFLc2e
tCGnwvFsDyZfsHao3YzuR+kpWo/kDwN8TwUHd3+YU/AyHXNG4Mozn+QArMOPVcVTjdD5KYnfmdkw
fuslToV92fPCR7+w4asQO2Ab78R6PgB3hrshENkBzWk8iRcKQseRw0VBbnSo7QLLAq4mctn06Hhn
5NBsT0S7P6k7iMU2gumtFdqLSU13oHAbthrLfm6/5VBXsEeQxnScx3kWUUz3exd4jzbBK0M3xdAQ
T4/j46lZHlnDkU+Bbg35B7/5etGBd9n4ZedRMJBduiOZpRzjM9mpWESDj/LvchSFaLtJpGSmXnF0
uNLZAmNx8ox4X9qCn/0InJBsTQvkumvA3W55MvkjqoLPC2sTcLKgFy++vnhj0O1XTdm4Od7HaECU
XdqKVx7NV2NmXczhYbkf4JTGa2r+vm9fD5stjnVscV7I0lsAMYLKOSsCDh82nLzn9YRLjaZD12be
g9DY8FIpQSwYcJ59pKrpTqLu+DNPft0DywD8oCC3TJnMuYSuxzx2n8jrFjINO4IEJyrHnS3Ow8d3
dcs+NniIEfgkf4RRqt8YytBkQaH+OhZW+efq5wWld3SeaJpjzVqDH5/m8llaItACtIhNHG2FCCwb
JmAyA3trEHHVyMY9FQ3nqfgR8S1l7li7DC8PqrqUH3Z28jFTBZtHYaXlkCjjHrTpumyPl9YPsTeu
SG17dBcLvtnnyCHQRAoXdSypKPPhOhyZDXP8L2s+rSgnj9+by303EKOGB95Sugv2//V4yH28qfVK
9trF+1gYhv2JfclKAlTiAjlpXPPz1x6sSFqh/tsNrXMPcXbOHH156e3Ukop7XQ0D5O1m6apX/pir
upBrjfWEtg1jJuvxj4cW/TaPXjZbpD4gikksqFxU8lQ4s5KifFUOkCYdg6Wfc7/s+PvB6gp5ymGV
qY+5IG0UeGhtqwv2J4rGj3yN3UtmUGM0V8HKcksRDxwRRHYimpNkO3DaYNzeUWpi7bC69/BpX1AS
yw9GIvJYBpNxYgdCMI5aL/WZlFMTvbm6jptD6ccEKK0y4Fe/VdT+pEkIwChJ0RrHdwlk20oH4HTu
+7ph3oi5QRWLRIh1JUmMPT7eUh6CfDASX7l9A8bGPq7W11Fxz9vnzA1qCgiPhz7NWbbuLL3w14ft
/WcWnvw9BNaj5KcZInPMPMQbqqFLZ8Oe7wL+GbCeT9RAyeDW5AB+AQXesna9QYuI+/J02F7oG1KB
1FZNn+P9/aqUHaLyhyWJih2ATtAjx7QsK2XCpo857hrPeW9/M8euUYuHMlJAxX39vBgUa+y1lG1y
vxniTpOcE8pd3zE6oWhoNtNEicOJLZL0ADEY6Tdu3nVZ9T1Ot5tYAptbmuYRkg5gywpSk4TDJ6Cd
/CYI28yPU1CjKZnsc4S3y8h/FkWQ1Fez/RkfOP+Ga6LL/Mb8SFR9NybrhKHYqOX4KqEFdrw/f6rE
fABdyMecq3Vsc0mS7uULGmDypjkXwbQullf84pRa7ORtmeF9OlK0qbcYIE6rRDVOxsO0Q5V4HT0Q
x11jjVVxSIDJWqzaMMjz5I8Z2akm2teGS5yz89P/UhNIb/CGuxP5JmTVhQ5bdcv/qd9sgaypD96T
Yokik7JKpDzG2NQuEZOjPW2MjVuVzf1wp7upKyBUwEq74gZQpoAOJrKBoCnQyc9j688GgLgYhduA
RPnLuVejmidaESiIgf+XUwwtOJ3OCSeIlXVA3iCCkUn1jvxiVmH0xAmM4gHlzo8L6YgYit7ku+Mh
Rv9c5MkUyBIYrSnmZflX0oJHTZ0dSm3Mynf9zpzpvpO2EcqKoLC1CvQ/D9UeM+GHG2wZyBsZT5yb
2v2S6A6bUSCOK8W17JaMsNgOvhkMM2nop9VPL7qGxG98snS4NNh10lF1JzzBaWonUzh89iyBpZpw
xUIc/kRshBCNEKg6h8KY4OlyWDxQGbFZlUMUJ/nfYv/0supHM+UTN+8G1iFZAzatU8cdbCNX4/TK
WWcZaFkRQKmgpXuis+A2t/fyX8/gSAky1FeJBulZPR1PE1Hb6RH5WCSKx0x+u48MBsZNlNQg1HBq
T5PimDFbIOGBgKci8sPci/LRUanITunjhov0NdgTDeEamKnezbQPXoGD6dVGV7Y7NrMRmfmOR7Sv
nS2IrIW6NnGQBDz+vVLT9xFqzi/u/HaaYaEEVJCum/ebNAP9Qee9Rpra0R/6gpWa8+LyYxnuPPLh
yIV1NHqDW7RleXUbEwLgsP0x2HhC7fyjkYizTZt3Ngvw4T2DIP+SWvFdHwoduOGwwS73T5OoQLLb
uvPZlpzMYfjEmVizU/iR+v6vD9dOc5x58CbpovaZfGZgiUNapbkx9EzF8DmmVKsDcPyHq/jpM9iH
eQ9OHMfvLPUGW4crb5EzuntIBco/I6425UfRWus8b9WOA3nfyUG8ACIdXJO47GyaTxGTn8Ripju0
M3lSpKtKR5XtaMd1OOG3Y68DD8mOjpqIa+8Y1rk9QwD0/hTcuwmeYYz6TEM3XgA66V/dcqcUkaA7
CHkHodEirecWJKPkELLERc70tUP14+LzLwIkXkWfpEMN3bmJadP5rqXUNw3Bm2pk3r/mrq3DAfPN
rua4eRU8vSgBd7ttLz3U4jwLA2rWGQDUiWD+uV3GSg7VUeFI/0fNENxBC7O85IJ3PFPm1zrXDEHl
HPIDt6+mApjjry+NPulWXA0QsyHpUFJzAsiQMlbJ6xom7536P42WqS3k5KcesDUfE14G/p5eU4FO
qRI9JHCyNPqF43h73d6Ex91ocfcnmn2B4tVn7E97XjY0FCQ2wm6ZQkc95rZNXfFpbiUgpfnMScdp
Pm7OpjUPQAaITSTcnIP3dHmpXs1r5G9N31aT5ODjw3hTdIi9XSiKp1p7v4UmRL1lLYE87dUSy5o7
hxrkMATrXsaeg970xzdz1Yh60JShWTyPFbnXh0imgOVHLhVxkO6WZyS9LGuSz8Z5CIP93I/3pi2z
T9OpfSwrnz5UmFLPp5CSqu82C9qXjTa2qSA38PPuTKi/JbcfRthkUauswjazHr5qhv6pOIRJfDzV
5pjQbyDxmmQJF+G+wvrs1U3ISkc4xcWanpPisStojm+jHG8r2VcMJYjV80CKjBxvBeh+05F1T8oB
r2tTy0Sd9L/HF0AQX+isVBVbsk/erBTg6mBiTebIkDZNrmv6NYaD/k45DJvX8TuhLSoHGjtFmHqm
3zAGFqNC06Y40606M1/P7AjdDM44qORMcVYgtGqdaAJm9dKws64QsOdDm5TFThr8wflYOnSIB9Pc
YzH7Qn6QwVO6NMR4wRU8eL64YQVCNGPi1eYsPUKvwOnuKNkEWC2BXVsIDsuKG25q/sU7Z3Yl3Fsp
KTWb9hpMy/DUb/h4pmEk08bzAj4fgHefE381+Ok7G04kw50l1WpPvZ6Zx3bujsoME9ONp2nYDehe
AT0xsfvIrmr7MWOvbg28cOQgAtuXj9jzm7hUM5PMO1CYFPs1PhXpLY+7mkAV7WesqHuBcPC3aPNm
6wyrOfcLRsDQHBSpotwHKbb6dcGNjGKMkYLQa9mxzs4S0wNbc9qi1VF5MD0u72zlE9sM4V/bollq
tdRAhxvL/jx3uY2zvmPK6+BW7K1Uf5qnLb/bsE6FClKhZ5O5APfmz6sKOpODpl5IZkwRJIVDyDV/
QnUs4WAlEMPRs1cAd2yi8jiD7fGqLL6HLcyxBbDsu5ku0ZFveC22hjtLpk8yRQuq1y+r5zFEPu9d
gl3FpI9z3t1H49kf8GbLRW8qy0FW/OoAIzo4tBjqLFn85T/BRaJpjMM8J1WexNDixlIqSSs5o/NE
vpczlKrxkkMuyn5CQYSTAYuOlmUhzvK+kNYEjLgpQdcczgEngd0MECdFqThA3bj7Klwo+au52bja
JZwymrU6RWzhfNKc/wLLgzUJBKLXCeTmVceFZEJE/jjDovTaiQUTeQmWeBIdmK8QMFxryHigxebA
IXNfhTXOYdBJ02we4g93p46o7b9SP7K5sgW2nAQGSBfh/h4E1qVGwz3vtsrpRSzUqXo42l+W1Eud
FUfWJwpJLVtz7g43gjWY4nmcqQaa3nziUHU5Aog2JzlMxxkmiq0sJkyKGcH6CNLvYP3f2SbQRSmK
bcidF1AV+ppj1fE0GPSuAuBuYuXPosAXwZOMXohcJsM42RMTUudDUHiIzr9uZtFXjLp/q04WAOb6
2KWYw/TZHpMjutPRk5sWIlc0zv/afDxYgSE6MiKbiZZo6cpUddWyV/dz9iPNgx87Kez0p1bNTCq4
U2ttAOaL5qTrxscU8Auuhe4UGg4/tL33CNvZVDEb/219arlQn6kAPEpAGlYusaeYTtP3H0QEFGSc
s8e+8IZpUcjT6j3DMgo+7ZdPRhs4TxGUVDN8KQ2Av5x5pHHc9n3/i6Se2kbCl8NALxKNawd9xQpc
SHb2LUkNBbAJibhwHfULKG7bSjZ55hr+MYE4EoC4gJ8w6Q46fPMXz5qwi22N+H8i0tfmLoJAt2MA
p4O+MJoRI18A8WrfOk8XUsR4jUAfzvLitm36Gy87T7yhsxoxhkch/x2f/4CcY5GNwF2R4vesxKT7
Rs83pEuzby9JPCN0Hf0agVYo0v8UPoJUwyK5dhqTtSTX1VMKeIl7wiLqlo+GdlPL398EGue2Gh//
TBnJShqYalpBiopKRMHlHxoP4BsYcZy+MtIJdEO9YiOtCi/0AuugCOuzKXqjCfsoUKWQUdZqBb2Q
aLm8vqboHQeRRORzdXP/dSLoOs4Kqoz8rwOd9zpBpqbu6rMEyT7C6cjSFk85t5PMdzODcpGmZbJL
3RJo3SXEcNjUIqUUYCI/AGx0mjoM3kkbdV4fKXBh8GGXXv9WwUtrxjTbXLNup+pTpzzi1ocbVUxZ
JT2A2QZJtYdwhxa0Iv5ylZ2la0hB2yvMTk2mV5kdJEP0B1ofceAYwaVyUdoFm5AQuhCEkbI1tKMt
SEWedspf4vqnU5eXRHeKzfry/uCAGWJiiKGeiBHo7JSbeKuQp+RSR67ogY6ewgWO6ur91Y++E5jq
KK3eY4m/1aibbjb7LVKyFqJI6Dr+CnSnACHwrw7VOZtkgbxkeeMJhILFTlpryEf5jhwCh6YK4+kx
HFJCRy3HdWNHufWxnMQf8bytmVuPSTj4bUe3HErN62BySdMPiFgXeVKMuqQccWQyWFayHLI1c2Wm
JdL2r3WixlJIRMOLysaf91eJI7xMgLYFkO2wvglonWVVH00vk8HRImBjUbXExIXdUlqPuSS/KyLo
UNeRCMTh524b3cylhdDEupKFf0d08miB+V1hqAFzCyREwGrzM7u4IPuh+pIpDVkI1SxaEtrnAkKp
0HT4Aa4S2/7k9ivcF1U0qckFgrwZsp39xSElCTEOUUz2aBZHan4Pj89tgU2yYHjgfRQwtPiFQf9R
RTZf51RvO1p5ajiigOta+1nSmQoUP2dOwk1FR3TA7FXr7ldFRBOvCgMijO5hMRG+lyGBBp2UEwWG
q4FbHiNUs+lFGpMp1m+rRCkO9JzDpXXIaaKjjzw82gb8UoTaUsXypHJSqnZSxj214wBZmMY37x36
pfyR6ySHT4UxBpaPw137R48/scNix3QdRdmG0VmCRlw/eToftt6vvcbm+bwtSK1XELH+uRp//Ho+
fedkuCF4AYS6eC15A8BZqjWl5QY3ISma6B2KFwpn3IHF0cBZ7l3cjq+3+433sS5c54kSTjBADsZu
9bu1ya0T+kvZVhwsVMVGxtztv9F47NPre3RUDyoUBeQdSfyCP3wFWNLTv37ygTGZaMxuAhKGiHHx
75UcVnqGpWMmTrzv4Pi2kRLRtWOw3+6nSdBavgtJXDxCRMFmAA3pspuo+p1SCYmuqu+udbcw7vwq
cny/WLWAoqzIHhuBHUxXKYg9+Joiwm0wZvr0WPnnYseSeKe644tntrd2WysArpcMR/dqkkzqPwZT
4REdqciePAd6xeEMUe8ktCpYVbGofZtoEK9+/4EmXY/U7Lfa/U5ZTtxqgHeA0T7Hw3wmxvAdJbCB
2Vxu+0rLMYp0sd9cEM++NegydiZ5TEANDkmaAn5Lo4C2zzI14V2TkKBXrdoodpmPtS5qaAAXZzXH
i6Fs/Z071rrur1d9lC4bDtf/3tgNkjzrmzHJTSlYJmg4CkPT0OcZZJY+dHjqPsca0CaNDRhyAMsW
0ilREfDfH9LZmPqa5ipurrZq1pck/wgIB5JO8x0XVswwRVNxF5f6U/yXdP1moNuowhR2792yEu26
YA7POJNFVHBYKGsZ6iLTOAtV20dSwBv1pGjlXYCSOYW47H1XfBZU4kY7YTOj1OBw0Aoz6w/ybZe+
N2085QJC8NuW5OSORQQ82b+BU0kO3YybOwNksav7aVEdR431iPEaGIcBr64ty7ugSCS8E9wCkIo2
7Flp7IHocSGRbvkhRgvin6UM7wqZCWhBxaVNlcsgYdydJc5drRFI3LQCpVUyohE1WGJzjsOpvJyW
Q4Y3OK0w2ZyplwNCOvLdX85uKb+W1MY+SrPMothu5OKWy0uOI1mzTR758Qnns5N2rG1OChIz17Vk
PRC6JB+qqujlzMhuy4eLw4b2xdCYjM57bFCsLxYGu1kQ5vOS+Xlt8q40V7kEc6pAjcyJagfhR0Kd
dETtlxvx+IzRXil9USg18RIYRPGNKWP4q/TcBW4pgH8mbxZllfSkVXs3hnsPU3bGa6BVrPZIh/4o
2dqOWZqG1msWczSpe3MsvB9jsh/UFd4n9tpEouKkSnTxfY7rbDJGRD7WT/UGEYyzylHJ2FleQNmL
dvmOxne7lrwa9sR7UOHMq7IrA0A4PtAImNny30boB/9Tzwgjpo0ud+3xBWZI0/Ui7Nb939GLRVnj
w+u6GTDqIDtb0OcrMO47uQGFmmYSaUKuKAf+P75JdxD3ooPZGszz50dLl+oPu9sTlVIsb/edtpme
piyPammm/SP65NHgDynC0/ZuFCZQ51i5LwC7/TZhHsjR4iL7PCkHDihZnqCq96MWybtIGIEHUOCq
w3qs7Ko8RbiMc8JZHhxeY117JUwnrpI2/0ROtAOXm7m4WeWoY1AquoJl+C4THXl0j+l2kgESn+oD
hF/Q5iW5XdY2BACVShNLkG7m65Brll5jeQ+0++Z/WLNiVnkjEnyB14tao8ueMOH8cET7KohCgs3r
ZXZRgbkSpypm/Bt4jUxXqugUbIUC56TxBUbOpijLqPe6oU9mQd/EcgmtijrZXC0Qjzl9Mh+o0vjm
Fu5b34Untpuo2tKof3snRiYkY1xDnd+4rdv3SRKtX0YnEJA3I6boqWmtexo+97j/Lr1DM0/vWtqV
uo96X5R0SpeYdgJKRt3Zqqp1H20jUnCUzluBwveYkDrAKAJSoqu6tOL4qe7vl5T2/ohjWK341bXN
Nh77xR1zwi/p+vF7G11KylLikk00gPCBvs3SSgwsV+d8VFulP5hd40P2zq8R1rKLF/aIQ3y0mPDA
A50lXfuod8Jwwh87cevmW1JdVg5P2ShOk7t4/N9ER78mY1xZ/KLmZV8+8lo+18TiKlArJp9puXiN
I6j27xtJvSwFKEt/hXIgi7D2BzyLcvIH6slVyJQBRW2vaZp4s2SFxzny4V1tI9Httx53xZi4dgTh
HXugzqM6BVfw7JDUblVdzppCZY0dfamY+IbbjYISwpmGV80OjZ00CCja2wFsciStqs116v6Sm0dn
1boJe6gGyFZQBteUQBYz2jo/y22M4U/BUTrrMQ3yqzWbJKlmNPwlaQjH2+MGIDcBQQeyR1rmA9hV
fK+/doHEN+A/t9U26wgYZg2N7YbGfvxVGCPAIVGz7jLZyAtZtn97e9F2ZboX5JjINOlXN4fylFvN
yq9pDP+Ge3yCF9Ikhb/xEA1KOVNxcBTYkZZX4rfjwU+RVgTUTuym58JIHq/3O3iWeW6ibWXsRMqu
gGa+D8AZh4O/wczZRV7KYwRCLAa7StSDpV/D+PydS1URypjz6+dbminkppXUxdIXJULWfWbOvmTI
Qo8KUE7ihBVqKy04T6t4aThNFeRZ5b4zPGn0duWjIsJNoWZhOqlO1yWlMYvJmk8UmYfwEAEA2vf0
j1Qsf8sSZlgllJkSpquBSFgZl7+pc6bmQBAg4e8SXdEBBx219rogLTW9UjB49ch8W6SLzomLkm2O
wQNxCgu0JFrvaqhxWf5TM0iXm9g0lTYYQMTtqwnUyoKBwkTFKtfT8wJilOnmgceQt9fvuOpTOM22
+MSPu5xYMu1lHedC4qYurVs5laRyGehval0E78Vfo8sQJ6svlQKLl0QRYHVQDaLbtEybjjJ2rPdW
EiBngwudCeaHo5CdH4LCT7KoXcrpkCYABo6OiFQUPG1anjF/AbnINj4olxcH51aZ5tGrhXey2BKY
bIUSusfP9E1qwzdSsYO1CgRDCaSok9FPWdQDXUY4LlYNG3KAZ1t6ROHKJe0002f0WcMPeYpTjr9B
zYUrmV2rBfCJ0/A5w2OsL6KgXozQqivmW0K/FCTacvdV2GCz4SVTHRIcLwVuTX4oQSHlngAZjOv+
M9miJ+ZhPhQQrGyLeztw0v1PsH2pCQUB4+gpVPyDaIUBQ5C6co1kqEUbxVVTBEIxnTl9wjugfG0A
OZ1CPEisKXcX7t7vL47BWzd+hMnjGX3zIyMbXuokpK6U7Tbg7ax+CHVFvfvBXyFikm0KgRIjeKfK
rDmUbZhGzVDlax6t2N732YdhrOCmpFQW/EMK9gIHxaZLxKYJ579bnVloM/9bNlWbBA846QQkxRN+
uSaXrc/P724DOHRnU/RjdhJV6L6PiJXpdoOkZzYocEbY5bp9+pV+70Zu0IA8DsjP/IY9+UBJzZm0
CVmKoPrrx0knSIsARq4kwyCPOppbNF2gprFs44oMX/dababGbnnLoOsazDQmtDoa8ziFddZDI1ge
f0wn2f1Fv40NSEK1wkyGNCfvVZiWr6sk1tHx+CL9yId+ITSVZ4kXOun8wHbjwlqg2Hf1aL8jE5vj
M7xQbQLClwtiKZsTBU6d4girnFT3RObZz/g+hzb5zt1HUm94sVN1QOA0nmrhBhQmxaTDotU+oB/n
OvdsHJBQwPivBjqxefFNK7VQdpQ9jVZjVvr/HgVIM1ITiJXUgqZwGr7tifi0sdX/o8Vd15eUVQtP
HbxdTg6mOGieRzxbu0kQm4gpPlphdDUVGtO+KRFVlPn/8SeZVU3j72H5M4Moun2oC3U6510n8XFJ
78cxilRWcelKJKCNX8qBO8sbRhG0ylXvm6GCGlePT81eq0dksHBikIq/Pa65oq1PC5xveRmyrcAz
GvgakxFB8nvsZplUKvI4sqmCCrf1rOnN6IyqqBWdj35VMFsaY/hO9MTzxKGQlOFuF+rkVDLZitu7
G+1rVSLouUKW2bXmE9g6xYWNp/DxeQxVt17/VmfnX5hwY60htJkwvLyrr7D3rYyCXr5Q2HrIfps6
9kU6YRmU2JwWH2iWnKnw8ishLC9NV9DmVWn6WPfhinMgFEDDcDfhvx2RArZI7+S6DNarGoxoGdiA
0nBI3NzQQbWtaKoKW3DqY2PFtbe3jPQwaDwMoKtWQMV+zKCBXmQjYshSmGQ+BRfFXtIbbPmygP7c
aK/zRhprBuk2ovuqKlb31w5MmIGoYoTG0W2xoK8rWhKrEYKHNgrbmoWQeGvDKz47JDCzwgtgJEq3
LH587DVTzj5XodFeDNExKgc12wwjTk/B6Xi9RhuMpbZ1Dq39ai1sBUKsKTnFykzrIoyFJWmgNRC9
Pwck8n9eoCGv7XzWh7rUxHTn17DxmUNcKtlreqsbz+/28dH9OS91tBCBYudiGthb5puqCNXdQGcF
BmSdBjkHa1twWO3OOqTj/O+BErXwsviT+6NEVztL+f/2iR9r2S1wu7+dHZXFYMJ1JG391ePMxjRr
GdzY2a2tA3WPMIJWbTWkvZQoBmD0OT//bT52ZpzUjrSG8Ibrmfy5u2Jc9bt0Mc7jFTkJRenrcQzz
NCVY8w5tdGL1h2USn6DwhmK19riJa7Be5LeiGy9DMg3vPMNOKm0QC8zFDXPihPM2aqYHjxeA6RLR
TPTcUMoE4xgkIRyEtW+IIUklnbgPSs5nrKJyscCw5f84OTJqKS18lA1gLm0BMTyJtPhqTGfa4RIS
LawIDvYv++8k9D2skLWSEJ7DC8WvSVbXxAN6SQEh0CUjdPHXzLW+KOrl3YFqH6GsYURANzmFjTbh
G/mG92vQ0d5XT1BZOdCJq5nIhKbr6TTNP1eyRkcZWv4A4ZfVUrkipezbvy1vQqqIhTFAXYI92D8n
gTw7igfbX3eRAcDsugnUgi9kBG1+yOm0I/d8FsNZ6PbWgQCTFpbpQIFUTr0CHfFdfD/oj60zWuj8
j8J3EQG8ojFCoPy0YEK0DzSLzB/ghf7oUeRHSqbzQcRL98PEQZJdRLr8me4kHi64ZhwqpcDRLeQ4
tdI2CIOHmj/1kqQfCvlKI5M5bxIFcMhvQ/rZ8mewxj9dzTq+RPXxJbFwcZEL3enKE2YuAfO3NhFP
4gC35AXSIn/zyEa0i8tRVsq3SGnKEunzV3xGsFAlL+ku0tIoxKUg9xzGeHcijP0nE6TI7VTsqf2H
pXW6z7Qe81DNtQWn4mvMYGro1FkRh5vKkgMtUyGk31u4KBGutd7B2UlusS7KjYv2C5MNqoniV0lo
65V2dkNDqIRIN//q1n32n1oVCeoJeMg5PrFb+xiH0TaEwpy2pBAwsGdsuYVMXvgJIQ8B6ZIdo2yc
tK6cvFWQ4LgiN0dAI4rPMI2dwjG5mOIvGXzPi/yCJqt7jmuhqyH1Ysc2yZKBCjG9235LRHew2Ve/
JubYqMMu0OHSb1T8MmX6OXLaZjd0EORjrQ697NqttHbqSromc+p+9EoAbKNQk48cWN71rgTdKLeW
sB3i8GqklKCXQYx6VBFewVGCaisQcG2vYp6lC17T2zD745wHPimBwi+BY/ikQo+WgLvHjZCjSRru
xTC1/38p2kBHXt47L2HcUthtFYx6xQ3QKAfP4szp8+eMzoPBIEPQ1RjJSaqrYDzMXpm9+NCW39/d
FOuMAG/pmhCpeAWKu0EKu1GZpZ5yesfQRgRWU+66KfVPL+UACQ+dSmx4bpfG/vKw0hzrNLRE2Bl0
niOSAPgy9d1ARAwhyHNd+V7El4558mrk0rM8jIQ0ITIDYJZIQJws5zVLktt622a5F0d3pOLMqMhP
cXSkzV6e2izE3+W8RyUAwk3oo1CArG1SXvPYsdkhLmy/pJFT3BcEp5J4HoLONribouOBUN3AHchM
hDL5uu4hBPosyAYkCVZjxY6KpEw03hBxfLKxn2gDKGdMGdBrA73ancNKhrLJz5ZXJT1XOWd5RoEe
7ppvP3Wi/nyEWnyM32/7cL0Qrnt3lcD8dKYH2Op/svyj+oGwQhEfNdTx68+fJw6OhdPbY68uhDUQ
1FEdQyZKFsJHCILnyq+pLQDhWbz4nq9RG9pg6hC/2JUdcjhrPAUu6Gz5Gz+h9s2/XZwcqewdJvyl
ohaqafd7Gv/Mo5AVebx1Q0kCEimO9HgXczgUu7HxPRQCBYW2BMQ1sS6d3Dcz4bFoxjecipCCpvBo
N9zrVm8xYRKYkYTLrzgHJiYwFReDBO8ypsjBwsOcmfJpKjnN1iHu54HuHx379WKbl5+JJ0xZKQsb
YHcmONXM4hfRyhhYGY57vtxxiFonXTkx0mLgXgrvfEYynGEUpGR3D6bSXt3H9M/rBqg+YYrhw7KZ
LqiufmPNCHyl7XEb2nXqskgwVOcPV3lbrBAGSlzhiVFB1ugoLMkuA9KunSLxk8Lljyngz62zEP+f
GqBuBrstyicrHIkuAEf1kcMG2kROFpr45NoOT5nN/YgVUXuMgDUKMmvHooy6PI9YRW9WEVuKgb8P
+naqbKN42WPdj4Ey7ggj+jYoOLSohX8XoTalXTn1rY49XKZ3ceUR5g+JO96PvvA0eOg9mBE7BfXZ
Jue6XclsrU8SSOUJKZTwTxwMjgKGwDkUQ80p4N3YEUzi24j9XNEtJnlutOk/MxQ6icQERqrZSv1g
sxXIwMG5mdJKbPIlB+ItCzGl74ksIUfBUzOK7a5md5eHpV1h1nvScQqbS8ErtuUhyXO0/sOjNHCT
Vn9GhoPEe21phcjjp2Yqr/mtjN9iRDbTr5NJy7c5Pxk0z6y+f3J/AWHt9DwYSSph5gVF3VpIL7HA
K58xexqMqsky3pCsKh6aEhOhXVWIAGGodrMdcJk5xgexERliv5UiLfCCQhhF231LTLVnc59cqi4k
lEs6sXc9pwYOi48hoamLXJP1qRHx4tfrOpyDM9DqmD3ZNsKm0cyTHpJ3Z6rRl6DegsOgI5c0qkj1
i8k358EopB6vbEIilaGmnZtM1DljcUwQJmdOIqBLr3QAsnJbMKV9vOWwq+1lQLQJ721/4yFJPg9M
sHhCpcGwkbi+CqmYG03t6yaWnrKZh+qMlu4+35DPdrqZtb65mxt0G6SC0udKzfjpLeV48bgdkiTr
IBbelMnnbNMiImVYP7CSXG2AgWUZhjy44SH1AsDglffXZH+q8yqyJxvN6s2MYeEJ3DY22J9fIYPi
BqccHG0Vn/buHEMtgXIZPSlbz8krlfCEeCSpT1kl/7RGgGnFUWdS6GfT0GYqEkjn9tqNQYmRnmMN
c+RrXeTh5ETQLN+ZUH7fmbBU+9soCoMiJYZDprznoHT3bW43HLUX3FdroDyAzjf9flQDixEzQyaH
7JUeEmdU0o6lFG7Xjp7fV7xMPZqqUy9ki4HCoaivb7nIvNuSYqX4/vIvaHhY95/MbImzu4R60YqZ
EmILAr8jMY5iIyPwHijMyQ6JtZwsua4u5dcMCM6tpwjKI7aYCabVJ3gB/JcWHKen7mEptpq8i7Cw
x/+LGzHScmqnbrGJzTu9dwUM7Mg7oO6B4cyWkP5bRAje9NdeK9PzMG/PFEWP/ojdtRdqEejYlzxx
lHdO5ZfTHS8VZH5J+CtMAJeOsIg+Ff0RjR0j5q+U1x6twA74/NDd1QQPLX9xtKZ01HjCyGy+C5cR
Uf8ia6DNRSz5jOjyKRtjQeJTv9zvsrYPsEGhhyGU3MhHnrz2/Fut4IZdRkoJAUr4d6AyM6b9TOtv
Q1mUsq81lVuYYZ2Fv+gygdo4uSaE5vH8RwtY55dtrUyvqPOy7R5+7PNQw2FeCcrhXjPGuIj01cyZ
UqFPQ+SzPXb/v8aY6jU/PxWfPvv0oRIGHP5Tr/Xx4xP7f8F7m8zFy2BQ9KTHkI/Xis98WbHjxgEZ
FWZcq6PYLOhRMRZEbU63RF5o9KVrWRpQfdUyck/cIvxINhZ2Hn7URC43eYr9LwbVbyMNfCu0ET02
DyjyC5KMy0x82FcE6jX2pjXARV4UhZ3BhZ9MV3bzFvPFUsFIFtApAoD80+Nf37PxoaJf3JZJD+Fe
LbcyG6H/ezHSRg9du+3xYQJN1LonGg6fbBE7lXDyGRDJ6EPO/vk5ZxjS09IurmsKqBKRtLF6hH4F
V080TK+eL+x6nJjrcOByjeG1Oxt1Xaa9KyyLkmS5Q+iQ8WOcwnQFPJZSxTyLeOuup3KSjBWGGLcL
R37IDid+MzpKeDGjP2B3lJarDRf4ETWui8hqkEdHTuVnArdaTuPPs87w5/jglVtMLwCDi6PL5FT3
RQ45ThF0JMf4myJ2VlzNeXAr0CFOUOuos7hl5Qpj1gyn6bNTXoXeEW2X66u1MPz7eJbr4XMv4Mml
VvkynKflLFOd6GaMr4Puz/S8PNHwU2YgKiDap9s5ZBWP1/sBaNAiKLj2nAy4TzoN9a/V8gVkQ6R8
123CHpCnHPlWVcCnfydqDfz5oZfChv449QeACs6ifuh2QgK8JsyKC7+4o4nkiOo8eI/9XCX1UYZq
GTk6NnmA+9/yhYz65oGpJNOuk/Ab3LcQXS6p+e16LOogusuqLJwBB399o3r/6auMOGwntqGxETAH
aovWtUTBesM8eaP99LhrSrzk+JRJMURzi0vVJ6SszA/dM8/Q8iMRlKpk7hdFqfBRAIbPh6p+0YZS
cNuMDKrwOdYSYGlRGS9+sKiRiENlrOAs20YUJmNqwI6VU2jfnS4t3HsobUOHhMBioy7PtjRdwETD
O+0B6j+mtx7EOM65Ib1WdfKLjrnvwLN43sZGdncTOITvEzRjFbYa1CYGbWYu5h7cx7oGCtrnk1dJ
8bXA0KDj7rkkVDR7QGUsgDYzi7qxhZu3hyYMnrab8MwE4sWh6JU2d4Tlp82p/6hNTuyQLzp/w33i
pTzN9QC6ffQYWDzzrU58N82a8gb00PoQtxVf4I1yDI5SYRBj3VIiDAJUYQD680t3f0yqclfuNz1c
piZI8+Wt47lQs/mnKeHEXAf1UAczggxGRbTv20BhmGLb/xxcX4JW4wBNLN9hl0PjSAbVmKmETwPY
/KlerprLCf3w+E7vJxJIDgVRQDjHj2Lqb1roS6mHpJSXZOw1LKp5oRinUIHm8dcT/87bcCrhr8i7
qBDBS4f4aNG2CzL6nuGP9r2jimaprSSpQUo5q4nHucUF0Hue4bl3bZCma1npXXopQnp5LWq9ao05
DBAFt3FY3968mUQpmrxfBJ/1fEjichmJK1sCQzZvfHw/S59BzXJa5mJjNE9n0cxTYCT0xjwOt8ZL
55nvaOz/d2joiWDS4WHONLL5uF+cQy3tcOuHSKAK+0X7HeO9AAr6e5VsRMGgWmXoHOQ/YoKKi1SU
xnGBowLJJAAVL81dNpf/VsuVkik7+EeU7DtFoaRgQs7sm/l1a8vjcHi10P71OhOkrGPWh0zi7f8e
glcM240n13tMzip8q+cygkMWRZ/VH1XplkURS4dfLh2oVE6lH6/bOZTebsfFlA8WZf7cFRjTjz7F
kwW1vo+YcjAgX0I4PS0AcqzO56LYMMNhC/lnLxqfoAxNPaSxWTwjP/Mhml1VPsmNprKIdndWMD7A
Vf/U2p+XbCq8brxDecMaKINY5ODLZLeD7jRpmpTtKqMMyO3D3/conNbrzrgDDCmdHRTQCCuNoR6w
eXdpEAnwRPJWLlRIXLCdhaHjb5EjUokCgxENemi2NLHvRhsn2kBuD1W/AmROxbqg5chKv+gCc/0w
QFMWPuidg0U2xcL2V6AeDVJDzNzm5G6YMTZS9YQ5D/7P1FE0nIskakmLL3zFQmYoEccyDqBbVM7Y
knCnWFkGIOOSce7M2Zt4ifoJT4FQ4SeLdlf97KH4EnxP9FY+05AW4ioKZJjTr9h4djEhWGFrR8fA
Xa1NTxzoOBVmaNo389Ltamd8k6hF9Tpp3w0TC7MD63LMLthfpa7e/u6XikL9va9cxXiA3A9M1zpT
kPWdDktgYQ0Yq4ikBhsvGtZRJtuH/pKJMHMg5zM1rXOv9HMgD7nIuN8YUoyW741wBAeRt1pz+3/U
EskRSakqYlKfRiL3AkPEsqGj/042iZ4DHnYJyZxLSp1TMKXCduLdmuoMzK8pIepDtzz6ZybZ/ucE
KTv/yWZc815DKWSx8vHPlLJnppohyUDdKdTCTOmRXghMGkprzkrAxAyHcasypbHORvAlIRpWDiA4
hUtTkAlm4yIghnGqtMEXBkc3uvlsd3DBF1OvEz+4N7Fjwj6jPWIeWxAjFQ+GsXixZy0bAE5jz7BZ
xIcwimYw+WpOT4q2PPvX+iUUq+pekefrG3poSTV8U1gm4VlI65YJJY74L8N2YTt5cq+4pL8KDm0K
U3zU9/gbHjUu8Iz5jfd1V2barLEuvU3iaoBupOhlT8hfNr+tVoLSgD7gZUVNKbsswcY39dGJUc8M
HeN7KFtthdPx/v0szp/uCTZ40rokIUYqzRevID2++cyaRkYN2ObKIAZT0z4AG+13DDU3Km+QQGls
oeeRAmageY6IuZm/lTspoP6JNKeXaQntsqRlWud7jW/fcBwNShN4QDon/Wy1cMmf5usb+fDw3pmh
Lr/v3mjgDNHDtCeXuYh3ICh6CdZSqMnqyyR7BH2rLSIx4vUK2sXvlDJ6yDCzSvCce46vtKgMNnQt
TtxRVKnWtW1c7AVUKSSI2jAxZJQdRPfOLwKM4mr+xBG/XswKS8iPWbX3LFwPCyIMDmpMkTm2hTd6
tcmk5ZSOHRR3xpfc5niIaSfeMm8CjYltP728IAheKPzGABH5zFw+zOlvbDYWtoK7PITRrslSxPY7
pJ8wlLaSc7hoJFdZ1//DBTL3p2NckC0CUQt7ZQUsYMfBM5uqM6zYD/f5O4CpptbCdKDc/tEQSEKa
ktCxTrNzLMH7grcMJh+T/xoV6dh5r/3IvdRtRtyJ5wvuiIo2OB2pJpEdNoQct++jazYNpmIrYxz1
RQ17W7R5LqyFmmVPWwk8GybTRGtAQlahpPeYGspIrwkQTA1+BMzH9r14YUIsvnSRr1W88ZIDHBJt
O3sAc4JA3zsjLecUxAnR9uyd3F8yBQABHt/QoFv+hdWC2kakB0UiE6OOT6alJW2knkbBNXGkxsJx
JHcthHytKQXwQc+V0ONas6pLMgulvmgmWUaaKmbAlrL04XPYONyZo+8Ok3EY6s7lKvkLDOg+rHpY
lcxoNeDAREgJg87ydZD5Y16uULg1rKbr17tidVDOnT3aZoqN+hfkHrW8hWTK/0WQHgqRldfuPky4
erSJF8hUyZ2KrRFbLTVbdz2dC46fiJmhEaI4hXX/+Ej39PF3hxMjrg/mq1DBbCxpz0/vXiXk5tkN
qQeWPmLGAOsL/xwhdHdOloVaHoz5+SXt+oVTQJOVxxe6p3Azd27hO9IYzBH8O/9g/WnL6xgyHC9z
XJHHpzCGNKCTutyakZBaboxlw7lu1hV9kixObjYOvz3uAf4d++Gn/l6Y+MjN+ZcLseGibKqrFZv2
Dor5ievLiMrgZqpZxyYPUq4EEjlO6bCM5AgMNik9e7TT6w12+dqvrbmIsoMnX4PL13q1o+66+Z6R
hTWXS29A5bxTQS73AukE5O0sbCOFLdCo2SUGdFbhndbCbZzHav7Ib807TLBCbL/1vWoFjcvDTZbN
Bp2EiDKeYBbbMPZUnYVNK++MXqnxy9Qy13pIObZeqwp+HPB5ng6fwwFP2QNEqeJWXRWT8+HZ7OAG
5AGYF0FjC6deBElKK5MMWgPDeDHgNm4VVokT5EECjGlP1vR/TBzhwTsxkqmPC/dr9Psyzz0KjUEm
cSax2p36J30hII13Czgfvdi8B4hI6qKLtDXWnWIcpgA8B0rWRTREbLFmW3+Q9WCoH+KkY6KEm1C1
/QKuRCJ7YcEXHN8Ke6Avni/4OyB9wCAEis18fAshU/cpeVWGjd9to/FspfvDU4EiaXVye9QrZp/f
0JUYEQXst2hj/MNCyZZdkx9H6fr0zwoYZqBXfVkrhUYnOolRL/GCIg0qf8sSvnf5SGue8eIh7kZp
sUJ5cGzJm5P+52fi2zyEJk6S++TdTZiNJmAKRrFKDwszVGKaPoqWa3P+KruKK9G25cJTY5lmP1+t
JVVSPmZoyd+B7QQ4nDUVTWjUPpMKcc4bbPuezwUfsoOmdiQGCThMTc+R/zgs5a4PLzHvAEaQT1fW
Tweetvb2OcI1rwnvLSLadZA1MoRH2b7nsEe8b76qjkIrD+sHpbQRufRIaDgC/VG9jEyVMDFTlovw
6Q/UWiildRuDONIq/z4BXZ5WbzoI+VzFVs6vftSmbKU/2UO0o0RnlEa2kX+cDcVJwxngQkBOk/sb
qWXX3FweEit/8nKMN2GfD1Ls9drmlUbzL3wTWhR+k+oHwA/qg+GAvq+4TmjU6jC5jjDV1pvND/ec
QDmeOePLNFkmAWQyfxKPU53iuVax3Dp3lRdwG4mo4BaXz4Yx9aUOi0FxXKSBA8MSIKIr/vYEYrrQ
wW3HY1va9qFakeQzBrPI5StcvSq3exkG08DDAngQpuOdNOm0i5UWs58+N/DIlS/6RCSj/KHHejfK
+xaaKCCNeqxuoF5IbQD8FgHV6fHpMIk6zxtogT4H2KK0QGKWxHHxqb3d3zXzT0gv8Gm1W9iHE7kP
Xr4UuJNq6xjatNvCc7tOJvYLXzKB1S7SkzmnBjpZRjwOJHM8goJgK2KSC2bcvhNKMLb3B9+tNo47
NFkACB1XIxPk0AmccCwIpyGvleClN44a+zX5lm72ZI3Yryt0sEhfoqV2ZJaGz6ISh/0vAAiKmq2M
0NP54wKrBnVFqmDkP+kWtdB+Eq+CEa8qu43CVwSHscLlV5vdVp9nF0CO58qbA9CnOOaWoj2wK2O8
/wASzM2lvFQiWkUq4LMZeY5NRWWy+Z4Mmpy/utmZbGskTZGuYMQnHE7GyFybTVWT6pknPtPSkpEg
p9BnlME77/0GFQRakLUi0/yNJRpfrNOovXlGyyiqxmWSd/lQwuR771SOIXvbuAp2DTTOO254TRpr
C1NCJMTAeg1DGEpocwpmnJ/SA5BqYNGaTIunJDVT9bt8jqBcwRw8h+PCBksFPcTtDjPoN91yAcjR
fCnRIyCLrSgk0Es9KRI2x8FEr206bdeuGGvGUOnFbjHsWoeXnv2lfowUQ6S3wx0F1sHel4YNjA8m
ZHwXZKOfYBghnXucUqMB8Jr0V/MS8JZS3WfJu804JkbrUTwTerX70bSVZDYNyA2LBhkOreIVy0HV
tPO8Eecc3eIomMXC9nKvHfs/TI0N8N8ndfJaP3PrxiTcD3vGPEc00aDqh6D3HDIPKWYU6fbyO6pB
n2VvVm4T8QsfUe8/Gwj5fWZ5GAANk6FtoNcQECTq6CI6NuFLFuv+aRxU49h2/hJr+DHWGtLsjt41
8hnwQ5AsqFXFfF1F69WQdzIyBYRy/JzlB/6sa+BeZIymrhMKpz0O9jTdbzsA1J2sqTne/F9s59qe
dEMAhgeyoi4ZZzv1tW0f9Q75kEAnBZUXK6bEfQ7H9zpdIvAaezAz0biRAk0BTGzbQb2uEnBAcsxS
oR9DVWDQr1+Ggzy01WSEulEhhPGJmaJ2a1eZ29eHOSNU2DiOpKTjLlEM19Cx09qgufMO3fID4TNC
ofHiyiELL9fHOV91dlMEztEU0+fJI/78Stazm/aG3g/zMxYuocuaB3ftyVWI9zqWyki5WeuHH8tC
DCAtYGgSy/V4UNm3Q4d5qY+lxod3GbDwTvYaRc7rOz7ffYYQbr6vHG5mY19gLtpTT+LpqdwPeLjB
3WtEqiElWs55HXkuIJslMjLAk7XieSBhS/cqToSxNnalaSn6+evD0p8z9JnxzphxGVhZ2OszhXcH
GHP1KR0HN+if04303bn2JtlVxv1dxwHVCs3R3Ug2bi2Mqoq5H3lM/Htzx+MvVsLGCeEbeuBR0B3u
ISiS4oAveJFNAaO3/Mid4T/YTGvFy66HI0c86US2b+eJ3XSpG0Gq3+zkDULkaaZeTKbZPYBTMb+e
neugUliHD3AkIPwbeMo3opgLugmt666icMqxokWaMknaGRMrq1egGjwCb7fL5Eco2Q/zJMIfrd4R
Y+xYauoLWfD+TekSWEbAG8G1iWcNDne090Gn+F127Iv7s9FttiTw6fTPs7fxWmfkq0Nxw09nxpNM
E1d+F1Hp2ouAnFJj4l3K1fwqKO/+4eEKPP7vtU8Y6gQpfXd7xIIJNm9xohld62iMKQvE0rEOZgAA
PJcASiqsnB38rK+pMI4R/1K4GT+UR4pydHA5jxzY/gfiidhjWnWa0OlbH/TF5J/tPbOBg36A5U57
7Ue2TwGg6ZfoKVPDESbCofG4Qtn4dH0yKXKhoT5NQxp9O7ePSukV+06X5CQgRKVhz9F+V83nMIh9
f8J9U5MfWOj/7aKL0jYl5woEQieOTEajlLeZB7AVc3h98d7FuFUsgnYSWahjOh4bqL4eVEO4/kIw
Iu3cWczl8yMBrzNp8VJ4aYo7Bw0M+K2pcyJyD34OwhlRcS5/XVKo8/OPOobcLQ8qo0MJ1A796DW5
jPNmpZiOfgu5mhBq48euZPDF/jsIYu5zxBZ8OKr2kG+K/8mO+7EklkU6FeAINsyfW0SZHPJGnrnC
BfD/CR3e3s7tB/aJxlRL43uf329Q0tSGNkaZzz8Eo2VDiJMpj4KJVzavxGq2+3JxHaeUbCDTp6tM
ziWm1P1xwvjEQiSszYuZoMUIZ6jrqKiHwL7PrfhljbNci8/5vXTseV2fv7Z7R30Xk8+/mxCH78K7
StaXi/utDQF5X/Z+qi1ubMB1ZYHU+ZXG7ydfKpRu/okmFDw6uwJztyj2IMapPOw66+3GGpO2lutw
yuUk/cGrzUaiSeJpmv7DijE+yqRgPpAsDCP+DVeDQ753+UtwL/W54tF5zs+d6HYP+pK++PH5F44g
KL+xwvnY2E1gBIMTJnErWwOaXUnkwH9JAgQv0DFMzwh/wK/wdWSfFlVMBZocsgtwlEFICF6VXWYu
wcCkpTUnZT/OgY2pCOBRkw0wlAiBqxHk8I94QsZo/1CbhSCmyWNSIBDgEKYaFcnp8kMKcYPk/4ra
d0nUo8I00FflqIidlGQNhfoLBiQYVUDm9NsLrKLDIL64tM4wOx4su564lUdPZI+4gota6fVY2zuN
Zv1WAGF2ZjLfTCNpykZcGj29TtgGH3FXyEMhhhfJFtsAtkSY4i2WnZlAp9UXCZXjgkkpBKjKwcoa
DErqr9jrwELoLzjwbVOxZTnaLI5e67aiJblJSAMizstVg4RLmgUv57UBgOiCNDiKo8pNogFSICUh
cDQEzcGknh+iMEzb9Z+YDhJ12GNb53Ft+EFsY8BpTvIMmpIfFeewsQzBeVtLS/CDiSmEJAvzc0AQ
Y6YCR7GjAd521/ilMwdVKTVqqcnoPd3xAOENHMVP7UbuHKyfez5YiVz8fBQ+f/DZIR7jFiVTcvfp
th9TxGNFHG9Hrjmogz74PNLBJNJ/lxmkImfU0cw22kjMTA+DPkJ8AYJYeSIVm+d0oHwLQ/+7D/94
iFbreBzcUQZc8LPdSCWuc52NfLpJoGvtlUSoh7u3+d2r2LWp6kFzyZxqlPJ6Tt6iWaKrsAXTqzZx
QghIeA2eOQenqG2uIDjJtUviAd+psZFomIQyiiFlYproCcLF+v6hJQnF8H6Oa0UsePiRrZ9YsQMf
O8gDCGzCsRH+zhOtjglWsDJ1iREXjL0UrB51I8/kbeHqvnLUKsnE6zalHoUrhvTWeXcXEhegDxl8
YDHu/dbGVAQw+V8ZIyEntfMC3K0vHfWIJuPS8Bbb3/8Sqm8gb+LPDYRyzUMrqOGaBAss57yFEfmw
rMRqpY78HQHgt/q+Poqay7eiVhb7GG0BHLdHME5Td1WJA1s+IV51KGdgGx9NM83D3BigvU8T4yhb
8Zik0hzJvnwuEILDbcsZTbRuB5lvu5UOzQtS4tAuUYPLWSJC3nuozvnsSojtCHxdsHsbT5W5KNam
P4Av6obt+j7F9Jzxssq9jeEAww+uPH6o3l9gqCT4REH4r9xXkSxuDkya6/oW5l+TvxgM1Z1sOJTK
S5xZ6hcOY5FX2cbPwIKNweuebuEFSLp4XeBkcE8O5ueRROl/iG3GJVuaSd2V1y0cASsgN1tN6x6h
MMQiWl2/ks54yY4sSBlnDthGTct9Dd239O/41L63sMBI9AR14K7BGGteqo8FpxILosjEMRhbj58I
4d5sNS0PbjlK7cmIMxfpDrw+bt/Ygsm26Nnx1KKyAwmwmsjklzkGpMziQxfmB4eF9yPMHRoJoAIS
T4Ytt3ovsN0vN+7wjXwLoop8Jds9PNeVfDvqLJNL8rfx20gIQCHaqhrzVWZ/Fo+Wp6tE3oJJX4N8
BprWjCxqipDWHLu67/Rq1q7ci8QVNegVrlYrNvIdieKTIo/ct1GV86gO2GFMZRC2D+e9Hcts7bIX
DZQXONakexMPJVEKvIe/XWgV+HLU7BJXUNANsJeCnfIOml9TrC61Pwffo+1Iv+Df9cwftSJT+3gE
d17bt/9m/trKZ7CpIZExK0fr6YL2e+uAmFIAAj2Aq6MkDCbc74FtRDY7O/SOb0iIyNZPHqcnl2zs
xutcYrBCBea7Eje30HS8Wjp2MWWaNFETK0gVJCXFJuCXd1qQKS+x9OKGovOHUyI65yYYVwveqTCq
jdJwMVsdQaYsT8ZGp43UdFKtxVBj+q6TLjnWT6aUMRo18WK8BYqa0Ixypq6UZ34mgchHtL/9ofg0
zlsS+utIDOixcaciwg0vJNodObnHCavXVmSReKsRI/vUK5Ylm3I4BOmPxuTVhJiOeiF9M0zrbGgp
RsabF09CbuZrpEVqSRqDqLbFfjA1+Ura6mcomqDV/gce0sOqtSmgXS5mMOrJ0NmUiodt0ffwGTtk
BagMAlu/nLsJaHrA5g+IIa/0tdgWuo6N5f9VyRs7cXZNmTskolPznrhWB7vXLATTr74vOIrgHJ3V
dxDZMnamje6x9uouLK7Xjy1zJMk5Hwuiwgpsyx8cu+NJ4aG7ezQDPZKalok9GAK/AWZZzBJGyaxx
qnciCt5wuDUHx5sz4J0j7pFFSk6df2iirCbJyyu4pKcdsEKDnHY3FhDudRDFjkg+eP8i4cLH64Ml
etaChFfOG/9RKNluDBgf0CN/JiTrLrWywLyquV/MGgY1UUUcqzuYfUk8s0yyeNd2Ir/c/cyRbyyI
lEcHAM/MijKVeg7DswvW97qNG3rJtl/sFWDX4Y8Xpoh8Z2jMrpEn7Zp3WAA/s8qTaWEInkFmILIO
vCsz57eU8UfrJ348+DthgH/hxqCO8emTaoC/zT7qbZRHvNkenjij/aHkIYQ8ZMuKCw+MAwUJ7JRy
LXGu6YN3+f9dmbQzdkyuwLsiYtb1iMBE45yKEX0yCyo+EfOQdtJOe2C9o9NDGmaj402OeHJrwvVQ
kOKR0D8wlhAlbwAhxNVyOXV/tit1FwA3rvmkkrf0hh0cydpxM0r/EZD+SKLpdgrcyAzbGhB0mpqf
6kepmSpZzC5VcmbkiFZDFvVMM3k+yl/Vb8sWj5rRMTSDBLUV7UzYkq3x0yACydlhd/rfg+2Vttdw
KZYb1Pk/NhAy/iAEouvyTRfA0p8F3kiL06lIey6vcG+EtiTs31C3StVQ04KfWf/Fd0dJt/pApS+c
mkhT7mbyjKwbOID1tbcbBNmFuNtB8rZLB4z6MbBj2ZAFEkAevwRT52IN75Lg8E8h1qHIZRJWZ+14
lW79TSeQDfWIvk6J/GWTvg+q+8xFoF8aUYDbEP595hB06mCAkWSXYOL2oJZgTTML5GuRZfwGr17Z
1K6h9dQvxbAJVWnCKmGMAjG3oNKfTC7JszH5qn5IBSqYjhSyqR6HX8K4zFZN6jxJ1oIVyGchLJmN
MhO+Mot/m43XcISsMls1Imkc9TjUlGunNKAf31Cci8ui1RRoE2v9Q3Xzgs8DpOryEsT7gfWiqAIL
SiwK30jnIAdfMynz0F5UO1ak6FmoOCphK2kyIhPcykfQjR988ldZtH5GqJdmqKc3tggx+VP9iNxK
uOLGVONt/fOsvKy5g7p5O8DpFP4cfDxLLhLLh7UzgbDktIjhtcorhbr5QCjAZLjGNm7pQsDiIcjQ
fLLbnWVgzel0Iy8cIOCBONzoXWE4aGvirW2RcVkR740r+Kkx10AJCYLcZdGf96Gq8BjWmxSEFaiT
h8q8dLXG1td2r58dgv6k89p8MJsj0I2MFEsy/+/1zVuAtW5YakR1PazP3PJ7zy1biK8Ob2tH35BJ
LHIn9naiJFmHEJB9jiop/eNfyNfqwM739x1bKjBO4g+pC9zgTUcX4i3bdN4Bq3a05ArhghdV5deT
S9D6ARRAPuu1anWuLRpc4bNImdXMc8NktblNpKTu1y7iNxxuLvdBG/FiluVdWXPbPBo1G/lctafp
h3jLpbFJBMy7Gzdq0VfzTaHkQgL08MBJWMD/hOZ7R2ndTvhksMG77Auag2gvT3uOYRHYHjAt3FWz
GByXjNCHwPpq+JgerLXXIIxq8Mbsy9me2CQdkRx7AhDY9DFL/KQbq4zXqh/kGFkqPPIo9ErNUmLh
tbY7j+WjtrSCBz2h2ru5ylVGj03y6mNDZ10M5MJz7oVHKhOTAt7nEgi+aU7dePTpbqDpbxNnulFY
mnAt62VhSNvLttk0pGpSVAhFaFw1KAMcYoJYVWinq06YkmSl0f3eR3ksj6ubqs4udZmJs8AumzCQ
AzU0S7rX33RVIvlUIBjQKTp93TPptaEirE0CUM2Gd/DUPc7gTkgIx7Om8vXWhcgSeor/jEflBfdp
72XgH1i1KhKQsYwTeZbOqXNWqBMzsCqWkYflnVKw16hl8GrEKaHtjPU8APjPh5IoATwb2X6Ra3vs
h/KQT0mHjnN8QnJCRm2iqXlsKqlqxL5Ew6slWCso09oDAztpwSJ7fXyvFWRnQGUTTd0lkCb13OeF
BKAmjCeMhqyZnTYEQruQ3lHtmyYPfVYEMXEw49uuwcb7sZYG5wLXD8ZxnzTVgoVbtJGPeU8b8Kvq
vEO+aKOVSGPWiTJx1zMTgxeRyATN0TSKNxlZ63EdZB+q9LgdgnAz6l4BzTzAunBXIR1uv5kE/X3u
pOc5DfXIImQZ9gl5KX69hTE63aPaX6yqndhqiVBx82Kcb7HJGHUH6gESvbHUqqXxo7YFDEUuYHSZ
XFcP0f4D1skpO01k3n+tI7FfTlyhi26WrLJv16oDndSoLXImhmQo1MD3/Go1OX40qgNHFUKJfv01
CnM4S9rWfrUxaZQYcBUEjd63YTIlb5nQM4j+SIJtDN/kg85RKRAQA8RI0Cfr/5yM0bvb65mX8Tu5
54HLjPeLWJBufXD9o3Pc2QqkkFb8WMrwHDirEXph6PoSb9Ia3P/Vf27/uWAV+PiX+3FYniCc9adn
LkNnchNyFri3/OP29TBY9xiyUN13ERTJHD3KKFR6fdBXpw+CQk2vBV5HLe615zxZSVQ0bJK4N02D
3Mow+oWMBFfspAhoJG9iOiQpUvBwUqrVUT+kguBIxp0rKc33lUym4ipLxNnvo/wYNBO4KMra64en
76Jhts/NqYR/eDQJJGWS7z16OObZeBnFv2YZSmKW2aIng8Jeh5aqmBKYMIj3Mz3bq/jhvXBvVl+Y
WPJM9foMdZgZxaB3dYM8JnHI+5/vnkZi0+IOqTRe5f/+ZFdhGlAc6135Yx58qvSyDgTwdjUiTMd6
Kn/LT5oZMwvXwrZjcrbTeukrPflrTsxYcwWJ0+c1YjBtjI5Zlmo4JL833v6GPB0dixj5chx2PvKu
9g7UaKrLe2rQ9OX+pC67I4WRgzbdazs7Uq2zE/zfh3t5nhc0x6EElnqWFibowszJkEidq9bwtKiz
9eSvxGdOt26oTYfDbWtXz+L3a6cTSZx77j3xMo4J3wMAiaHsiooIRekJxDlLhmbRR2c7DgJ4UUEv
QUrRkHQYSb7ORTzih3cnIn4nWwVKxwIr1pQUPgJL1kCFOq2hlbchRkNZC0y/uS3ysIr8oAfUkA9Y
XxNJujFosz4D5BDJdxTy69rqcF0hrfWd47q8iKLWP23WJ3ewlO3vGPI/43RtMFgy6/Mf3varSKx5
IP1dvxypQ/1YzL5PWBXJt+bTvJmJoQ5qI2fzORFC7pvf8YFM7XyC8CQHM6eZsdy59dyr3cHUtfy3
PUlhMIbH5maOyk8sjQT/nttgvQMuqvJLXffh91R44+1vz+oSb40v7tgQiT7Yi/0cZWSi1kp/KkVf
7B/V+r9cNh9kKt0Yr0Qs4s4cuuzWgyowjSYvX10Rm/auFfWbTGbQzs1qogjg1dBGfjbO+AsZelI5
vxmB+jI41wwLZULvZT3Mu5qyNY9WVzCv0lxTWNBrkML9+OKu8XDrzezSOCZKa/TENo1hNPioQBZa
Jh9nUE157tWrUPn9Yy8cS+1K55PEKN3s9jQBaEPjtoqbiyDEtgUtQMgjrCHbkrMm2QNdYrsLRoUG
2HPHlsB2bgukOXNeVbjy0rixE8tQ5bOap59T1yYSMuCbJEs+zFH1fQKYCkoH/1EmPFcSfG896ruO
mxkkxq125+Bd+GKYKVBCAC1u0WsppIWH0fwoOYxR04e5Dmudf4XcxfJnCyYgCYO0CskbEYAK4K2g
G7QRM2qqTmicfISxXTX9bQ7xO7S0uMEWQX6gFvNnFGC3XPgeDKaHRTtTW7zOHAncJOos0Q8e//xW
dpS39Ei6jhCzcj38ksvvXgM3o8ZgdNUjasoyMa4IqrmjJOzaUoizFBy0KfTi+rq+uXM2RvKo9koE
kKiqI+V0VCQZxubutpfGmrayU/YeHeVGox16W2dt4wQp3Nk/Hyc2EogTUb9cySMDBtfGY8+0/EpH
PWEN2dmwUg0MJtOmZ9DH317yCSJITk8HeNggrLsvdJb+a6FnKyQtRLWUYnsXz9BHHgO74v+/ZZEY
E6LWcF8QFM3PVMoPX4AgPkNf0/znrZw9bc1I3IYnxMHfJEiaS9LQ1BBskQekswk1R0yHMhzp7iH7
HjvtJfadKUUVm0Au+0ZOLe9TS7Tjt9L5QbjU23apaVIxUcyJgIgN8lsV6AeD6cfFnvvwXz6oAWI5
/cedqHLJWHym3IoEw59jPunUBWs3Ch4HPZ9v6sfKYoLKpqOYnhM8tUcIj0uvnaTJ068EA6pXKhoj
PUhMpgb5Eljds5N6TRIDOZW1InaEOhIKsli6Ls2jv1bOXlWVVisVWF29EP+ljLA8tXYw9+CnO8E4
VDeOQO2/YGNgc/JKOTBzFoZvbtC99uwT/ly1OmddF+X806iKulz7x+l8p/j/cwuZwEaUbN4gSxh6
WiVqJ9dboLnBkGMu9gCKePawl9+izGqUX4/hkpSMFv5sgZZAmZMIFlFNQfMI5Q05nXppNSjW3uer
kWxtRlu2XYlWgfomuXb9/IgnTGvfDniXqwSst1vMhPnmRcJAP84bf0kj9tguh1wdnCsK6RygRBLC
bGxxV2ozUdExYSXnpB+Hw54mm0lNDKRQODr8B4rkbKc1l6FDC0tr7nGlvJKJjyRFHzn5RuKegJTP
dXxvFfwMOXxZ31Qek9mArlGT5CeUCQnccxAMxSLI+m4DdWuY3BDRvn+2etMFGsYCuphLnzjV/e1q
OEutm/mqWUrjF9APEjeDEdIxKqOlhpMOvkVmtf4PTfxkTU0TPfJX7Z2rOQRzG+3eZ9+tfkTp+5Z0
HPH1m4ad+wBaoq2s3ecSQa3hAoorCQR2AKf28gIDISrrIs5DYDuG7xfR+3Nznf+zHL9BSe0zrXaH
H4lYrNAHd+20Za9udND5jfZM4pBN66dLqG2mpwwANsRaAHGgxioaFWluixFiUgF/CmApw4TaU9Xg
9/EY4X27CSEWnw3p1BKID/DSpq2+miuUG72UzH7LFy6HSBITlZpmIdCH1RweHGcu24rg3SFIDeYV
3Ev/9CHlywQ+4P0ldvQDnwKZ6ENEbJf9sQdD3vPO9rUxsryUkeZvGqX30AHQoI5cQR9I05PySrFf
rZVApXvQtz1eEHUwVvKe8f78zdfa0u7dbL37Vqp8a3vPPEYBB2p5AoYMhuiFN1DAKz3AcyRgT9iH
dS4qEDkA7gaI8Fjf+lj+UKTiul4BhzAftzbqM52R1FmwOiHQ/NmZIlqundtIACVh4vo5wZYIj617
dH2OBY/5/5LGZaZH74fdkl0y2Pjz/7ROjpWeQ7fqtEY4A+dp0uEwC5qvSPfKz4h+e/s3ZId9ycwT
XG9dgRZGjRBJbaYRnsW5xwefSMW6QmM/uXLpXQkMhIIhjlK5IFzKj8m0IO4n+Pq1TYiNkZ63h9EU
YgnEQokLfESvJkfwDYO5uaE1RJzDJVCCoX0WTeeLY12y1h1iZ0Nfs02PZ4tUb6XmvD1sYZ8gNX3F
T+YW6W3+6fFMB/U0argG0Ca4FDKPpO5IKwHDAzbU62qVFJRUIuTpyTlz5xdnyZs/CCvk+R+HithR
sSaAgoq8MaiLUcittUmTHxIyhYi2AjFR19rKGS9oIKWqqkpnidOxfQF6EbkhIhlpE+pYEJw99S76
okrpKDRb7bnVp8S//ogPgIaTnfMYeB8LDtBL6KV9ecUEkBEx//yqZ8sOcszmQt+z2jm4iGF/VPac
QWHmcK1N01HV+ad658/byje8li0n08F/qNjy9RIVI4Jk1i+zDzhp7EOvDhU7OmAnSYwIhjNisASC
YSLw2A4pG9zYpKu/0S6BBRvphYqcQlG435E06CDEgfOAIHDX5l9QYa0vZnNOZ03vk+hJ6ja6iorm
3R7xx42qV4tAIWlsgspC+kuMvLcwAqAGCFLxa7QWqMBEiq+G0AO8aU5QWCP34L2SO2nughTG6og2
Jh8bQPXA2mLipCPut4wKQ4OWEYZp3tVxvYYQ67lOfSUzrCSHIdJjyi3OYnAO1tDJ8qcrchw6n/2C
oCYNDdUa0J6UPRv3Lbr0wfZIecDqdxAazpoK8GLATCPU8Pti4KbKad+L+Hc4kVNZPFnd5uSCncv6
evoZxXxcGuEEk0/y4hH5qYv9U37u9eEpecZRQQMlBaQXyuAiaRnZ7jmSXyTgtHcysUd0paamESkZ
Orgd5j1fodIWaiLgzNS1X0svxc7VvIeUmCEJQWKBnzedc8cgcqI7VRi467B6f4ZXt2A5crOjMbBE
84K4wqG4aR5Vd8NXVJf//kXICtaZ+43vtlkpYcOAMnAn88OmphWJZgS3GqkIQaiWt/1CF42zffN3
nlw1cn42i3Qj3i9I1zsaWWLlCNp9Tun178qTVuTPwlfckC0rFQTb2OH/mU2x45FG+URp6gWwVols
MQ2Rn/j3Tjq3v37Yc+rzhBFZGDZHNcOcEebTkKbiYsYucGA17CdZTnZG8iU9uqEzl9z/Wrlm8Q8z
jz7HfjLNI+seWJYS2izwabAY648FsDQJwv9e1oskRcCZlnCvpkpoPvYwJzbI784I4vZGylfMrtQo
63Vao4W0WvJkDBS5byT5jOwOJ3A5jchZOWnlLAihSWLn2TuGuWizPD/WwZGmZEgeF4HvRnAG8KRY
C9pAQaP1F5PVw1IniXqEihBVrZVzvSTON11TetlLq80pkA7jLyrYvtVp0oqxMbl7VAqJEL08/pXx
5PH3UYcdsU5fwsFQVlIB+hnRrv3i5oPFv7j8lofBnAWEP1RvP2mIbFQcew+F3wY6qcNAFpO7hcwA
f3nR/kCsF5V5hCzmsSXg8yqKJsZhs3HR7R9rz4bLa5XYIaMK2WOc9rqErZfaV7kmX4k/JogGFC/M
duwXEEdnTdY5t6eCq7TLaFHaQUifBHH6xKQRjNWLVJItCLno3zcU1u1GhKn/ztLIRdFyZZxGSmXP
ZDtVEEySf/XgINf+HbxhEYZ6SDz/GoaaQh9FxKV4eTMlYUUyUtnEhos4FKNwHEMCCqxxokYug8Mx
/Z99nygiGGWD7Fn9freU+xELvH9skDOoEPdmw9e72T2cFa10WnmcSqGyVfey8TlmRJy0FaJYrqUt
WX73ecnBnypt9qNdlvXDtBvixXZL6AfRZ0MgFMUThrvcMFmMOUgbjzRyvXf1Qo7tihnrcrSnzzAL
xq5cDPODDXM1F8UtfVvNYnsrfRIGH6nD4IbFILXcH18pz0gXIaqzvNiNHYd4zg6RxzhaMGPgDDex
diJkV2ZuxUd7Y8zvVp8yZ9TtSNhgdm+JXOsIGxcn8I2wCFAZ//IsdHDxZ8mKiA/tLcTrWRL3J5gK
6TMxVAC50RQpHh5Gck2i2MftrJPcMKgyHVTeBse8ZEHoZH3EhHQMo6ZZ689ArXW3azl61hmUn2mY
8Im+fjUd8j2saSFAHd4ZoBwmw5zE3lZ12Y8nnzO3TxwOM6oO/k1DgLVIepT6eFpKSptkepdBMceh
92OAqHIBkuABNBSVykyVUKTLmlTlAnZ2+idquG0bBW9gnObdHYBFhvLr4WHPQ34IXZNeq0ughWG9
G0FQ3dvoFmeypboMppy/dpzouJUfGiavlf/jcEnPIZahcjkZ4KaWIKY+TGPgTRR1np+pndmAr5uf
hdwWSZ6sKz64oshBzpsCHWxf1dkR/9/OC+mMSm1r4HaReg81KPCIj2gnS5uiUJPahKuaJmDekzgK
RJ/9I4745RWC87N/JksTAzd+2aQGVb4YfYiSvtlLObzbt5aB3Q+G7x+0NDsStofaQtCxa1H+erQg
WnddlqkYjP+LMUKU+MSrDkYIiDoJzlUqhgwUOJn3o03SjNcTxCFdYyUPkaRlYUVZOOviXS1uoTzO
lOGFpjpRK8IHmHfoXHtV44wfcwe/zBC5lNsqaoEQnP44WX2HHDClGPN5YWuVjcn+0Dqh0BIgFxsW
ZeGBCNM+Ew3Wne1EIsby07c+8bj4EscQ0Mw/lVFlYPr6wuLCi6yM0/1zZ73ZQKlP9Japc+RTwrC8
Bxb1a21umwNf91Ka46tVwXfrAOhTaa3JROmS7NMgW1PngXCnog9gSSmsGlCcD7tQ7dRPTZKt8+jE
6339E5rRJqMNRzLPb59bhnVmAv2t1BWbqkrNPgIa3s4w2+82Lu3eDHdklD2gC3daJ/wp5P2RK2Io
T1HKLxNqmuluMr/jwCjX0SZE6SIMAM5DdVjVIocc2cmKuRX+oXPWap6zl7ofOa0FWzAxkwTgvhGu
5E8DXPvm29kFpe6EGXIM4hueCEIYgzYGDZh3gc92K3PUfgP5gNu2Rs5idUSwg2e3wuFeoCW/bx5m
DVezEacey+jGbI39yn9qdfeQ42cqbg8CTY3MZv/OG4CRCJx05CCkCKqHID4bFbpxgruaJRB3sYtB
BRVJmUTZ0NCy1L1gtyj0B4yYKYQ4oBHvxau37UNk0V8KvyuyrXFZFDewNlNsv/Jk7x8IWrG0Vghf
blGE+NBPc6fhIGa8iCfFyRzHY3itH+ERYt7GlgmRY20PFYZ2fhUB1PzpLweEGG9+GwmwA0dFSUs6
MfycleutZJmf5CWTlkfPin10LLCHQRDvShYARVmrOyUt9TwkZx3b9ZYwskNesLbWvmt6qJcMYGkG
+ubcYIz2kVWtxaz6QuWc9UtT/rEtynzhDpQfhJNpjhmOOgjdLeR/bKLrC46dNdN4m8MSN6B3ALGN
CLuJZyroYsiYqkKnaOsRfMmuI5H+0tDIRs8gLytwCFDWny99NbE0k/q6H40i5nA6l3PG24AIWwmF
EQIpBWyfHFeWh1Ozm3kmUkuu2bUx2WNLoGjeSjQdSr9LHkDXompFFj+8SSgDL930Wwaz/GaRzEpJ
f6+Zf9SbtLnqgSQE2vt6vcY4rwZ/PAiBGaTXOrc/yCbBEThwFyi7RcdzCCd/apSA7J57furARxBa
pqQo/Fe8XFKTXISw7XM8X3bIgFDfdOEGfwqC4WQs78byw0W+jYb+I0vv6fzpD+ioKnpjMPejvFKA
SSNB8k/xPNtrtPc4coXuwcpcw+Clq9MuaL7HxF+ZMdbDwXUCE4XErmCrAGTVMbPSSf1Gg6sQsDjc
v20TEROdWC6MC8QhOpzKUTJi5nD0nMGtv4PharTEUTBRFINR+kEIwkcLtDN4S0LTYeFU7dBJvubW
2gG75+WOkJM5gfjqynSj0UwtoAEwuiWF+rnVLw1aQEHcTDNzoyGl3GnPI1bWw1ST8G2K/sHFZk8D
ytELxDv5BthqmJ3HeA2GFXPbL9bVcS+rf2HJ0Kid1BaVWzHDvquwhpuEPnDwOVQ5xWsy91iKBmgr
ahLfpXp1l6gUiTKcK1splJsk3mHJMCRISX2ikRHU4OXxp5VplsXknXwLf6lvcIu11xte/6t+CcMz
vLJ3X/b42ReH4rbV38OGPkKYktnXapD5oV1YtTLZgNLZQtduS/cdbFqqU83Tz/KWn5c24vzH2D0m
aTRG2vuRTE0WUhXpdKuJjIaYqSHJEyV/SuPlzJ0EVZgWqP30xZ6wpa2wPGgvutlitddv2nlmzs4i
7dgDd2cqWFB3OWI1c0CaJvVAKveI/k0XdF09HQw/kiFiENcOMEoWeyabuH5vEZ9InqGMqTV17BL2
+n0Tgp4619gXcIyDM+AaL4IV2gozhf3doDrewj5DuaRL7v6h4DK4iENJp/OE/sI4NYBV0oQ3xggh
uDyvXdAc/nBpw+cTnmLSQQbf/iL937jMzCqflt9WbM5J7xM4MjPbsFtxttGB6f7l75NhY0cjalwR
DI4ehLyaQcrEnYaRrSaehm9Sw5nCEaLvE3RUO5JzRVfPWcUQ830uBqrdv9PzZUC8JA5mppWf0xRe
4rnBcpsntcURlrZg5K4oaGjjMd5uKekQYGPNcMVq6Hm48Rwoh3QCC/M+LMg9wv4tEaH/+e0H1iq1
I2vzSrjFh/4fSMvvKgYYj/pY1RfVBEU8yGPU7TmIO5DN0WBH2OlX5IWYFOptiRvVlJx6zXbT6kZe
yjqxB+Jd1NlEjEnWA5iTCmzn5SJTX3J6iQNdDRvoV2lUxogAyG96qVYRob+cgyo2O1YBtSG8/xyx
II1rpZKeKUZi2kMsbMe3lPkIrV2Hi7e1NRmwjmNaMsevwStqVEeyzQvEpIea78t5Xxf+XwEZaNsM
MaIs6F2QmfjIZVHxOjk3iIFj/MFnBEX02o0uCjEXHDnYKX/rA7CEzX1CBap+IvJG5QeNBBLG5WtG
3p0+H98MC1hPsRHjMEXLmuf7R3Fm0ipL/htJ2X3XY0Y7nAVbimL+XlQkk3vjAq76XkSE+sz0cdDk
R4cOLcFsLxeWUb8CR1Xo9ewUZ6TKkMkVr2ZohdA9uY/94jr9+UK2IzLCC6mDaE4wlehLcAq2g8+N
CvW407ON+0E4NrSi7icxcspuzoZQSI9zOHZqfMIBiOUMdHIrdQoG3rIGvW8MVvo3tTuB0Yfeg7w3
H/kXmpDgsecmhIAs0R7BboKRWIeC2ZcPzKe7xOVIc7IcWTET6oLA8SouhgvdNKC54t8UJ3YtTIY3
H92XnYG3cILeYj8LHkM+ac8pMGeCII+QHNlLH5NeIoSubBTNeq1y1MJijWDF6sj+8guQ65kwAxI7
+KFHiw0ncwzPzbJ3LwvzJQRXbAtDTHKlLKXma2diz+phhVKSYYbw6LXOro7LAc1uuppKl6dJB+1+
L72GHrcNWtL1PtK27/OUNAfabEqPhm7tIcrzDjVSnSULWVUf8Stsq745x2xPSb7//QbTGhHppEYg
xY/ugbjA3YZnYhnSfI762s6bnz3NCH4mag5BqNZF3kur+jZ/zlari8TurK1Fuh2uMJgJO2gARgH5
CULWIS2svpytnfCtgfAPv4zcyGcViKderc5RIucxdQulTjteoWpKZsALoB/BYlPkMH7CKKjFgd5P
PcLslVCIXoqRm5pvCxWlgkBSpcsqeRt4DFTXT2+C2T3G1MYtPuKuC78pZsX8X8s3cKbxw9ZT5A/s
XCwu9ktxntC4HfGBS0JDX/dKNqPrBPIkcpJNvK7pIqQ7DWz4j2aUc1wJlQIhKSi/wxjJ4vEOGKpS
tG1LgBQuUKFQ64hX0iFv5JXSqvNhzqqVLOQd/21GUKgbfok+YducPyzVv28OmB0Q5jcUypE1pp3F
YOV8PbIrNfIHuP/Yw9N6ZdDRZdtxmJvy9q4n8EjLVz8ow7FeYoTqT3Ic5aUjABZnrYniBz/dXpPM
JvuDf7GnEJgOoUgt5LZR10k/utPRcKfvcAs8oOtvVWYRYDKZDhWICjZ7Mc52jqjlIu+9K+pEcewr
/Dqx/VgiYj9Pzjs85OlKXmuEOaYqFMfSnXerO8BpoAPrczw8LROYI28NynIHhVgDngjKoMd+Fz01
Mt3Soe4iPpyQeHVsNU1z3C6ZK51O+7NMoPd0GxaYLNxJ5jqp2+qrryW//Z+5AYmwuy/0He/ttTmu
hSmgUnFiKzEKy/JLBXA8+ZjbjG1P7qejh/asDxF+7o/9EOvl5H+qSBEyndaldRqBfRAhYHCCuKGu
fOLgeWjnPxq1FARpmV9edPN1bDN+U2KFkfVI1TBZBUgZuv4KJb4GEpBm74UDDnXR6CaTsgDAdVtW
6Suo+4du4C5tEmkow6xliD2dj3gVPEOsoWQI6p7urfQ5/ijz+OGacvd93EiTSU+Kx/7pZ2wt3Q7y
Yg25ovKG8qZHILeX+va10rFSUzymuEmJCjYz51E8vbQi1nji3sdiptZ2/WzJ3zngWSakKuND7ZGB
7sG99BQVixbmlqmVh2mCsSirFlZDtxyQDljXsPBISqyJCSLznmDuro5cO06CfOazp7nmi0nMjV1j
VMJOMqMXNadO8oTWBYZ02m+wd69cGDGjQZ8Jx6W8SpX2+JRcMJS1YC6xu+AzEA9J6+frcr5Db9As
5dUeIhrekpMst7w9N9Eo72opb7/r6PR6e0xoc5sf4u2zQYtlMmLhy8NHIMOcMDGK/273FsD1iNYB
0gMcxxuDWPp7HpHCqlFJaHixF91KtatUGuSggbY7gOLpumWVUknorH1DPMvGuQ3AroBKFUO5SG3f
Fg9J/MWYipyoqzwCLzCdISI+le/Uk3AqwXsnZtpwtHtFxHEplZTvBmUe1DBvI9mWrpZMsqHJvQDJ
bi4xw3yjPATtJtgiRZtvO26xXhyxjwZZ1mw5Nxg81SLzQbCJXKiTMlnECQsJ2ys0i3QU5A/aad6G
GzTRsqY5MgkFpxgfLb1GRjRWJJy/2sjWbR8No7rEqrtsKm4dbzLZTh808pezRLYqUmnKeVQnM25Y
DpIndcsghvz6iHm0jRMthXI0Buo3hyzFiivoAoalZXHFUJNpGHxUZw/BVVX76mHClftX76zgduXX
zZMmSSKQwA7JN+V+3CK1hFr8tlbX0kDzpHLpBai2FRuXwr9UZaZRa/tUhdPZpuG9i1AJt0AWhx0R
qwq+6lAlGifhJ9XRrTwnQN/dvoeGZsnwv+fWGrfPHYZbcthOC6UrpsrO0sUC9ii3ubryqDdqFZYk
lRgJmod/SCPFQvF8xw3DwdhjQTqqxznevzXtSNjTEgnIs26jsXkutGp+T14YGXkztSIJyreaYifP
2uziNZWL1pX50uaDBNF3s+ULjODIafwF5tHwv2fq1+JMcUR8qTBD6/qmuHj36Ch4odlpZzpyM0bo
6F3KsUKi6T6O8+JZGDGQx6jdP+cVrZoDpKlmxc67/cAoaOCY9B2JJFx2lUhS1rmddsdw6pJ/P3ir
oVmd7duyYMzkw/cRfNuWecLuxxh0vhWjgEQ80cOxukPzPf/hztvCuIihvRrQtuKQKW5iTOb046Si
gol0MKK6vsWzlrSyKXiBEiI+JrUes2rUpYWlWmNUYexVwt+FCoqPeiWJdshaASSvkeNSfW3efDjE
g2Aea1inLgCRGUuitYT+/G8/T5F7yyMrDs2YefUWgpExOa8CySUuYEO1QZ9OIPvlOPhEm5qNViEj
Qlhu3lCM27U99ZpEooN93UVHJ8YBivUSW5TkhAQrTvY506tHhkddOVUd+VVDNNB1yvOqARNV1DS/
AQZ/mN1jju+IgiFeBioXJBU/XT+Ueiyw18gwX1gx0BjCYHqtA8RZi9eFAiBKjeFuaOExhyfojzMA
5BXLxWjprDuXsaDkbVsKeDrr7IG3/e2WvLusV1UE/QmsPvrqAI1VqKPL2iKiDLTRt//v3nrMOziW
KMmu9GwbNfO7XjrMNm4nN7mUxKlgxrCajSN/C+N/+hGT78H/eAiIlePBWePEln9wWRf/mwobS1So
pwEilHgPNDmgtyCeAjBgRNLZgnHmRckzDY7Jtjdqk2pSTdGZ3FVkb8d/tqfMXZjgxlje3BGg5X0u
+KVlrjkHbp7TKnfYYZmxfWwYhDK/MPNiFKiHePeoFQVXxzAnufQHEvOjC8JkdCO6LZhgMsFKtx4j
WOwcuxHbsIgfh60NVZiGGFJmXjMdnfnWXgqwzNovVN8+A1wsqHd/lo8HDb4qYO90WbMrvjF8tpBG
AVWiDMYjPT4J/sAoyi21f/b9q+iT9UtTu5df/ktAW0pDAmlA24iQo4naFx50LQGQKOf0HFx+UT6M
Zb6V+HIKGturk3M0tgeOWNODHuwWgDg3cP6gOTwSYX/aCIKnoxzYuk7uffaCu+EFEBF1AmzeWSIE
gBLYN/BIp3MwJES76XqI/wutOBUc8jmb1nIAiyJ0Y7hIetCNc5bZUZvMBHa7U5RJiAcyCXnSdyKk
B5UlF3LXKrQF/lxRhAOvzkyppOr8VdPkRcLB0IOKBwa/zVfSih73WOTMU/xdEkxpnOhKAjYnoaD4
LJ3WVuiVXs09iWwWONx3FknEJ/P8qJP95FwqzzuiaeO08FNBKl/v8S4C07qPrG6fYCuHGnuDw1xF
6kzeQ8KWQMObqjqPRqzem3lhjuZ1zp9uDaK5cLJ2yXJ++QIXbbwRqqspSxFN9VI4ayQhQ6ffog2b
xTfPU9dc+PGPxS+TvJVO5DeAMPbFn4EWiT6tF4vq7ouc9OIGeN+uz8x4xk9HqWAPt9SGl0efkVJ6
R0s97u5HxfcuAq39XZnbLaOutqA0ibhtdDytoppMmA/AhR0NGTmcATSbVGXPEV8TYDHqaohxK5EQ
uZJvlvv6ec2cO2gjR7f3qE7lc6xZQ+CvU7EkeQULWBJetYCMrRjX8c/zvOItifTMvxGeRKp0ZRkI
EtM+3Vko5lzsrASxjur5+VqPBRuRkeq/Wj2cmp77sFKYwx0s29KZD3TeFhYsTiv7/A0+feZr3G76
hJBW27qHXIb2kiojZKZIc3uErzDrzxRBMFpAW0P5xPrUWPRelysHxQqVx0+XuDMTWQVWobVTuojU
VBvGV06R4U+9UKeugqEXBRwMOtiHscyv24VVp6wDUGESHv/c5j6ksLLBKjs9CE68Xu2Am56lERlR
Xt0xMaQ5KtFo5jnFOa7TfTUJBpcTLTPj2J+ahjHjZIXlGomLFhwZdZCK9xnHSnH81oUiIh7QoUuV
7cY7w4lAVFwGSli7BRVodSnO+u5IpWgFPNc+YuFOZKMNJe2LyiKW73RWaikb+WXTRh93BD8bhSY3
vwfHJEIZALDOPglwiYC7yekEq0V9sApn3JSf0shta1a7/NTpRpoIIZM7SCpUdNF4Z4Imq+CdDKKP
EQzI6nV1pwDcL91Wnt+gEpISD6e6PgxgpZqXxU90sFPX+9ohM9OwNcXm+lY/HDxafp8LNa4onFBi
RqHnZIy3KSGeJmB6kDw2G20dkrFINHWuRbqNlwKq8BAPnC/XKJCVqeWiAlAcIbOqFwXlTnSr1Mge
jxQQaEPujI2Je/ms7gUUx8ew7u/4aJSCrAYuzwFxRA2LFq0Qg0sWVP76vnbWpWQY1TQLH2Xq+it2
iVRYo6PHcuGUVVAPmDsLv7UnkGJ/ALFBvrsaTLW31dAQ04hh8qft7huQEF2pXelBsxujjJ+hRAd/
e55eQFVrHdAge9Y5S118rdS3+SumZjxBiuHgXUkrStTw6BrrzxtQCmNSgrbNE4Ks7J7dIeW+vBRK
+AnooYGcFCxZSH5VKON5Ec8Kq73rm0yIIGDH10eCpOpgfvpDwXAFTEMUavP6TNMx3XpJNBEWr3f4
TT21dV1CLL7JIusYxaaFACAO2AqLKUDnRcJZQ6W7hUrj1UTuCWoMLUhedmmnFAgpdTXsTNW3of9I
lwHtZv+UdxjJguqJSgHueKwCrGxAfoiOhrKcIMkWiORyUGtwAr1iJtLuOFg5fZeu9yl6kbkqZIGd
Pou6pHshwzqTY1Hl8mf3gPrceHNu5bRgLx3DCCuMDrrsYDRjZUjuuHpFzgHW2fCivWjaeZSi3HX7
/LDeuBKF1bF601W+iHQdfGve2XMGGl+0qxfwfXj3y8pYk1BPE/yAFdh7PihBpN8APO1fjvAoGz5q
Ev3eeVDHEl0vQhpP2Nw2sLC9P7OkaUw67V0ShvMShcgDU6Lboj+kdDjjTwbeZORUdBH2KVoM602U
m9m6PFaApMisf3Rd9azLUrk+CxP5ME6sm5xmTe+Hw93IUNcmYzNNjLR/NslULYDbhaoP/SuC1A3Z
agv+AviFocffw0J9ixGDhxITnT6YxZ33D/QCHuUw1pNztbgZReSpNNfE7ukAggSngFJDQ6C89Uqz
V4M4kKarsqGCU0IY9AXr7C/3pz/1nJMFjK8xv7tB3leRDL4XDOzVLImKEvuZa3YNmN1thioc8OHG
oEnul5EBAZCHD69cTjHWwyJ2wChwLYDhr/3qommYywTFStrhLSRvxBKWGdNF109cUJZ0eDQOn4VP
xDtcxTpyUDZihXcXQOO55jko6qFx2L+8ybe+CYtljFm8V/WRRw2X9zpfOYKFFOgB3WnNFFrQYm/t
Uw8fkvPGa8yNOdxyi1bPjUNVRrFn9IwRKfB8O73Sl7Ahb/0VOKZR+QBwDu+ihHdLTFLiaHQUqeXy
oJu/3EMJVUTgniD5X+P7MbBCsbIY9+2TSrF3YoLzo9WYcY4Wz4NBvNXPXghyRL1PzSEtz05RNFnn
VpYZRib2UWefnPnkkN3jS0YAYKWqorDd8j+BymWDnFf9Z7MigtNux4ptrL/AibAMjQsFEkHyRkRh
cYDPrD2nHSmPZSO3nkyC8QE/wVFxLk49nkaj0E0OZR5ShROtMOghgMfqGESJ5zX73gcXwFtuQ3IN
r+Un7hKdT90w51d2zTaqiiiUogfMS0rUGHqgLdnv4WSUT1cNaJgQs8EFstwVbzYOr4IKKabeOSJn
fBhb/Lfj2NRL84Mh3iCQEtcNT20snbdQHGOdHALx6op0t43+FsoxkQJsx9WHc531adYHYWWgvlcK
sXCWAChYX4tLvnzl/MVKCxFH+nVk6Lqspc7yeUhgBC48TV8M8NQGsUlazHS0fsf/WDV8u51ndeMc
kCC7IBAJYHRQm66hbMiVAAQArbgG9wfp9CLvELBHSBda3aQbj+pUaSHvaeN3NfuGEzTkETClMVm3
/8Zftr4ZwJb4X5Qh3dgD5I4IMOHDYNCAFvgb3wYKNNWO9k8oncLtInCsoTOEBOlmEC/9JEFrh2v6
+w6Oi3pNIGQvuY8B6uD0+zLNTq3L+AfdzbxJd2IijBOZDd2VgTlQ0ots2nH5aKeTGnLgHajPrs7Q
iZ8DKMJC3gwMwqg2hhILb739qqi0A65uUCvsTDUlSnWTnu/N75yoRUGKEPtWTGLvMYNFGz29Dk7v
PPNjg+NTt+fTkJBVKx9TEwrRwsEMbc+501RfYwmR7qmQm1zZYfN6rI4wWvY2ToiXZ3OgunjoYVMh
ouGKm5xDuDdWGsQUJTjdBbVCat9Dc5PZHreMxosWDFkLjjL+S1BtmCW0mpcpN7TxRgp/o6sPjiG6
e6bVeFcUbYknGUUxaTeCBtbCZtHiZw3bxtkWJZ77ZKsTnI7wemMe/qD30gGHWmahbDXZ9kHG2hJ4
TedqOb8tguYpdg02cZexXzbTCeyYTL9TBjkuSQmijnuxzyE2sQk+i2JYJqDCAPhhn8XSx0eF2Jb0
BcUlcgUUcbYopQzMVS34lVNjJIKryNzNYLz/oMOZnoDrOct8epI7A+mksSzBLWkTf7GMRVCeotcX
7lsndWOst2MDOxqsVpW18bp/JRtxceONuHaUO8QYEkPfGh3T5PkMGi4TvZZpxNbZxXFxXw+p9Xgw
neYogr+1VwGm/XHsei9VcQUhkCc9PxZotSWyU7QawMiJP6HUKSQ4NXizyPyC/UrNqMMwtTeDcjYX
bxKdgIe1n0rpzgSGvijYkhm0V0nDX26obEVpnyQJEbHzOSosWWdgKgEuqt4k6nMW9pKnPE42rEFi
GaR/LWP3JoUHAemEfcPQIY+ClEmchtgxNmbQRpMPubA8byeLcmcAJ08WX7yyVAeZrZjsTDehPQdy
AJ3vRR098M7pWIKWXLdjD+XHp4z28S+AssjIhdU3JlSopx9a7t081JAm54h2ouLyoZeuFdznwxOn
gmwkRy3Dlez3ZP01ZdpehWrkOrUyg3k3eHpcs7f/pZR5FUqfU9ytPCaxPgy7AXuvRHOzC6s1JNKU
E+nXipCayWIRdGkavabDLcLMul+dgIePzB6xogsIt3FElNUuUoc8QhX82KOlk2N3TCLEYmUc7ZNF
/YrfIzMouUIXZTmGXbC9SadgkibkoYd9Y+DTvFQoYRERkex/cbgCWT9eJvK4lLXh8l3bl10grrpy
lvZfFVdHSK1Gy58OyY6u9g2r5+qhsqmgmx5m3KEQB1etlpmkg9Lic+p2aL/YGn1bBBM7IMsgOaSt
t51UTswKhC0/ob+741cCzCCk1ht91b0p/kvZiSTExFbj8NYpNWVq++hEMNvcAjLfiDnuK3M1yQP3
4Bx2JjyiA7/P5xDtKma+WGKke9F1TlchSFEIBA1LL9s3AdwXAQITMo41E//baLn455NTlGcwC0t/
CQniuq4Fa07XH1P0vhrTFIgX62iSEqOrRp1R7CP1KA0wpfJBjOdzvzFLc8bOfkbv0e7yLIaiHtXr
WX7SjsDKC4mc5EGCH7SDme77un1ehtugukT6YktqcSxD9UB/xE42uKt9om9LdZnn12/igro8EKLX
PYCoD5eccy5olH39tZFeazWiIJabeOj/KlQ/AmQCN958D9KszGEmn14fRhNG+atMWuP2hW1tVQAx
OBmV2jfgqJLTL1wN6bd9+fjn0mmuVn9cET4TcK6ysla+HUnHib39TT7Yup5ybuWKNwNK/WyXo/no
ZkA8scDdFZKTe1VUp4fy9aj5HM00Xu67rYV3YSqRcYZJ7J8TIwBkGIX+Cd+7LX6ixFWgabYRKAWY
4hUVQ8RnF1Wguyz63P0Kx5xBG2Qmflz5WxrHOc136Y4HsHrwqDN7UXJkwTv5z6N5ED4+dl6owIxz
LcJUjM3kdaksnj3Hs9wChuvzs8do8Ooi8+qTYnBt4a5hVmOgG9Pxviuv5QDi/uUvNSj6tAHxI+c9
/ELhjUhBRf2vL/DoMR3p0NtL2etGXafsNqsSJN1ww7DqOBrASBCJU+Q9/Y9PQOrQyhBPXVJ/JPVC
/coHGCAmwnNqcNSMgxCnCfmDGDz86tMsw9B7tpBHXoVUCZvJCyOQCPicoEEZgq1+Cj+ywtu+3bPB
PI3FnVTBqu+gg2eoQZgDBwq5/C3bJ0mDx/TbVFXn2G86URUPoezZ40V0N83Dtu/bmkFOGN+uCrhp
fyGADhXNfyczk/8JVIZk7JNamnLxd+HNNoPRFyR0GZ7KaSIV0mFoMztnU5lGI70KO6s1mwMPiJV7
fxmCkti4bOWqKceqXwJRrH4bydRcpaSqOeOfMfSW1sWvtgJWo1Y4fdITVOYTrcdiSaa3h8IJR9Zs
N34whslwpY9WRvgUyOygxcD6n38nwii8VLo3jE4awvPGQJ/pUpSqVaPRS25rmdMUgRe5JKZdRPh0
qDUQJHi4Pyj0u0NDwN1L7HHjjHCVznDUodSu/xQ78fnRuTWylAPyy3u9a6pgXn87z9/hFHBAZD2o
+oc1koOsSxEbqR3V/qmulurUt8i1nOgfqZHizpSu7vEo6SU57dWHy0QnOGJWxg9SgMLhO4Bb6tsD
Cs4I0pT4FSPrGBoa79HCtNB5AU91LBs7FbD8+B+bILJzFtEY8OYT4qmIt6KERj04s6esNJxedwG2
AyIUaZlbL7CNqcOD4tJv5EAJb6gQxWOxtToR4X0CiGOYwx0v186L8Rvw7eO/mttYvn5e82hzHsgJ
pL7QFU4wvC7hIJ+ccS659sWXSF189GZNmD/GRftoOJLCo72OIcp833YCILyuptdnGBEZjDM75jyW
18Db43sqOxSwj/rf9Np11bmKoxbVnDlIpTmeYRsRiPViMaVtQQ+btemRBmS4+F5F8tFA0xSVCZTK
UyoOeigYnQH6s4HrURFrbxPh+rmwpNOyJ1wF9YL2JNGfhHwyjv65eXYba++30rlSPu8EB4Qu+ALd
ny5bYFGrVfnsRwOCFYQMZYnhRlDVmPTq0Ht2M21oc6xTN2GAQJJatMsZWAfgGHMME7iGg7kiQwBf
/2gnDp522dxlAg3VRekuj6//0HG5GjIsa1pSRR4rk0HttfxL8dsOIF/KhKwMnuwDqX8pRkSMlTS9
2VVxM/fxmIitM4vKcVsS9ixW+q+hxQm/vIJ+TRZ/tfkA0KhWW5qZ5c+5KZzMHx/JTSfJQrRPlBOc
spfcdcgm4N9ZYFA7GbgtG9Ya/uRLSP9ruu7K8sv76+NLSG5EYc9GWtkoeFpU0/zfDAvGBjV6Y3ea
kRKLq67o0vzkbkAi1WO4PfDSW+FAWhIgOY01LK/1CpUznIkpRbVwjgZA69LcGYq/YCVTISwfGgHQ
xHVQ9InivOPuIBUSBl+NmjNoF/wLzS/T5I51+b6yuluHrsXRAqjTOTPFEf7DC3R4CqB1M6KJPDhW
ZXQQiaX7izkQMHcmg6FLaajNcmRp4c2ORzNqJKLutKlVGrJCL+ErdU4O3Mycum9GBbqgOO9j9iPu
pttXOX7KL2+ff27Nx/PpzlUA+i+OBKQenDYwVS8ZjPWdBUL9wunR6E1H9MCnmV4MBY7qaJIPxAcQ
uZe78JalOTDdvJQvDZIS7Ss0YxWjpKSc6kD7zTi9eSkXcAr6QJBrXXcDGtSBCwUpI6v+sNT122f5
dtr3RVeorDjABVgTr+AYSa7yyj1Vdz4A7Cuv8fF7cDrfGXGs8LhP8z+AM9NBhA+O71vgx73vqtRb
IPdXUdm4/wjgUIWH0mBNdPzIgRfkhC8Bi+tqww3gn30xJPOrh2m1jSAV5crKuYtIXI1srTIdQ9l/
YUelmb2RhRiGdhEp8D9w4wHC222cxnyXaVHssf5skTSLjEfE9GMoDF2jdJlzgfpmL7P+30k9hhN1
29YGeoaDlW+MW5KRO9GByKKHdJv+tN01KIbbh3aWOD0pRy3dxkYIyJ5EoTdW/pCMpl0PFWl4IQBr
ERmu7YifSQe1+/nlRfxvXYxl2dalO+JgrwfM1C+kRvGNpjcv2oty5nHEKpACc6rpRa2gIMB/99yo
8QDMrKx6XJQRzIziUdpqyojlxPAiLfYk1nSDn5SpD2IDAZAIH8BPTA0Au12buW4YcbQtW9rtWj6s
RCZ/YCr+7aN3MmqL0J23txzRiFmt9/wpMcnftxb9qdyTwWPotL6clSrbf+e0hZk6sJRa5lUlF+W0
ivSgetMF6eW2zTo5P0HGpcFDzI14fj5sOuzxkqe2SEKyHRS+I8Xzj0nA+T55+tZsvwD4Sa+syvYN
V9Xx2cpf8XAelpwQxYvsF3P9pNh/YBVAAFJ3DcgoZ2WG/xpIxgDQxuco7qSJ5/MpgYIrEY2OAhlI
LLS7NVVz2fxbCyHT+myiqf0WtoQXChAEYdY1ub04HVHcHXbRBOqEN+jXUxKNZIzsulxGHWeSRGFv
MdqCef8ilvACQP2WUpbBcBmgVSN39OlSmpvY3Ci6a7dT7+HX1Y1r8iawxupDfwcuXGZ6yxvS5aeN
mJgTWa5EjrQtlZeJeG/ms/5fVGzCX3701b94L5I8rA37NkJC1JajI/KfjTAbVvQcOyAFyTC4rsTE
imZyESwZszh5A0R399PCb7uG5g7ifAV1BlOiyWwbQFq7SABwjqphmtmw457EfC2Hc0H8P9JgLUTx
PFunlc2djOUqdmOyKWOLXQG70+iFBFLYzmaZfSRNoBT7dsFTS85fJhI2z+ICqNTEiwjkW+0HCEp+
YvIiR4EnnnOACb7p5KaN/MGetu80U3rcwiPw9AHSgCH/+7PdeokzYb0iHQs21MYLZmrjkUtU66Yz
nMRQ3RxPBbafgq0CcvWX+3QHoXsTsyRYL5Skle34+IyO22vfxtrdZJEDhBRXFs5qvdu9CL/e2Xab
SpfY/9s50yKBefUrwyh6r8tygNR0gjtPX5I2XK4qU1eA3Zy+wFsTjHqxAZP3qOQ1s2B8CeZR0vif
ldUX53voF387RyqQnONWdUjMzGpqP3H4FEG4Dkshyk6QCYLA4orB6heVbYo6qIF4DzteWWDR1KcO
oHzgfyWI0NkXQsMfhd6P8+UBVlifYg8VdN6BmQlolcdmxQhTBS6uhp35+PJpcxKkuThkb4ygvIr8
hSZ8yWT5QMN1QqU3DnH/XgXEm2bz6RA7hB5Bq+7Za/z4ZOLT8RhaMBeN6sCazsee3TH8iXUWlZ1P
qGjEctTWTzDO1hQRqwEbw5mnOyJLTv1dHmk3JTym5Db4RpcbMVJmotNcIhkJU2bOzCHQpw1vPE0Z
VhrY4tjEg9m1GHQBN9/AWkczIy5K+s0m/JK006v7ZtnzPJLCvUSgHLqzR3V6rfYZe1wPsRQXwhU7
JWC8B613ybzGwx/ASjtp65WGAY5Z4+nYkfMjP5bePY2+nh0qBZoCxsAfm4Rp29JvZoRJrAnm1zmz
RDiHeSZ4AGegBRWGgeBiw32zcnOuWBm60yIEnjMhAei3jxb/rdiAiuWZ2UVPhei8ffsTW4mePcGt
cdJx9L6gDX9ldvFGxf2n0mxULXCH5udBqISE3RmL2WO6UDQxmJvuUdO8lLRQQi1Izx6/ZJt5ecj6
IGZA/oAc5l77FERD18boTQ4AefQMpbSADPMle9TFvVKou5J+vcuCfhWEIvwVZSdsFPv5uJwlz333
89CloggzO/dQwhS5u3C+QTDN2cbexKsNoXtKc8/iWAfkTJUj2VbovoWsL7PR/ErPccc4LO79Hmqj
sgXRGQZL0NXrwjIKyslKA/jAzbk5Ekm19j1WpDMoYKAadwQ1iLBzxvbXGat/hIPb7fnoHqcwRgmS
Qr4zPub84naVTAZjX604nk25QfIzgqleDhIS6fMMDioTQuV5nGR+GJ26ZSImusTNO+w/ve+YtwZk
hN7/7g+GSBMiT5GAkFy6YWEhBIaYj1KYv9dDga8puXna4wj2wDlSkl/hsV/gZPYEoqEjFm7X2TZl
yFbnp8LVFbR0uEcB6J3qxSv++6DFqJRK6XXJHXJWIgZNLSJn5euCb3nIz+ZITq0tRvKEGkfAu4ZX
UFbkv0vLOJg6cUy704GXalvlagB3d4SBcL6aOPZ4Q0EZhOoLeQBWMz0pCkX5ZR2uCSF50PbeK5aE
OTLXUgifZEAmEWN5/GIsHe1G8pG3z9gG+BbHvbY/5WODqgyRNXJ6UVbAg8YZTx56N3vWGKWn46Ie
20yZMQSz932S+Bn9hJD8dsmeWsDiWg5travEkrFQDVQEXk4qfo2tJQhqtd2fBKpUe6Na5kVVbMqN
4qMZA2s574IKMy8MS8rqZs2xD7CpGGuTT1YvNCvRmB3aP+qz4nFA0e949wK8/rj4fVE9hD1V5Z8B
woU1Xk5k1ah5wVDFKXlolVnkyXQvFBOfplM5kX9gaMbiiUVY3va3fT69Dfj76WIw1K7eG5iLgD5g
LXDU/oixoVKtByasbysFV5hyB4krF12qtrquBLqnHoK088mYpbz8slh1XMdPl3ehinpBC8h2THiM
Rhwkja8iIRwZGCDlLbhfSCW5huD/Gr0RdTR1Ip0bvXOyB8N5S2xgsYYB12Zp4DvpkqBg3TxRHIiL
Y+YBv7X2bzuAmHkqbdg5CAJz1mQGtO2V2/vgS4XmWlctfu6jfN++SvZv1E96dMgrF0S0b/3qyuSS
sCxNX1SVC2X5QbNYDzjC50/bX4GbebaaK/bdkUQ3NqeClV+57Im37+Rcim7Zgurc9RrXvKBNRynx
F8IsN3EQ635ciX0W6eFM7uFlAIJWnAdLDB5G8K/8f4R12JbmELKoGPwHokzA2wMvarwIGtEEDB2b
K0EgkzJWh/1BlZHIX5aP+1LFt6PG5X8kN5DMw1+NkOLVh6fuKb9Lw1ihCErOeT3goPw63+zrtm5a
l7RTrlq+/J249di4Eodh7rezojGxCX11RcOlANUaNrv42EiEM2fqtYj/plWlyHODxx53Q/OUmuih
whU+meyLVa1n9V4HpQ5PiY1c/zR/RKMVZksMYXQ3dE52nSB9Mr9hpR3e3PbhmVuOXpTRAdQDRes9
ZP3CJCdQyDwFnljW98kcKydQsRURuPljw/OG0S/52Y5+t1cV6xGSmawcMls9epFI+rvru8xAfmb0
CS9+kHetA/ATQo9ETawXwIG7YU9R/+0azfim9WkwvUGOyylLFT6MpDSjqjcK2Udl5nmJbN6s2/RM
hGRhCHFBBeqFQOrKfq0XX3bvlRuyNtjRVaReWPkSNsehSeodcQno140A+9Kun88ogIW2wuCiCkIk
Nel2Ii/PmUThvI/oh/kQjGptWKJiVeyRiIBOgd+DIqolkjEmRdiE6vdO8Vu533125Kde9VNJTgQb
O1joqbsz+BW4FaOc5487RMdMjYgHZren+o3AgScHQQ3rsr6L2zmIZJuxTaAZojCNJSa4ygc/aFW0
b/Y8sj5EEXvevQrF6Lk2RS2QfkXcBhwN6XfnUHvG77GB0dmuzqa7tFjLOVSvzc7WdNHyGJXwd+3A
MKw13vFIWIVcwzGNz+/NnixIGMVNu/ZXRAIuK8Xa3u2TqSwvpplK75zqyKVpLqCsTQaOA6pIQTnu
1YasDy7QHL21Xj0xlb9NpBWOxbPVbUzU/2pD7m3Tp+vfRzGTwQz5D8jo/L6oXMlU4UfrQqW23ZYd
VMfVhogfEwKi85oxv7k+7Lh8qu05CeWluvRjbqjJXJffUNNX94uK2yrDSRT1+wnU+Oyg78V8TyRY
WqrhvrfP4ihtSSsZET1epVxSYGmK1ZW+0GxM9WsveZo75e95pMAk5LlL5MS7eudG4JRVLPpSSbHs
Cx5crWAE+UrczquGHH8BLYBhOGSgX87Nium0WtZXSgvlSCcAL6q/xNP6zJX+7+IuozlGOvLfjadd
YJp+xnUs63bZ3ZontjTPS9G3XalZi2MuGVPfxocJo2YL3ZYnZ58OTixNZkR7H/EsLWwFtaKYBnxK
6XoxS/WGwTjZH8s2saS19S0IgpLbzBwJVSsBjqgMOYEA0DIziOF9yql5DNI/T9NcQp5gWMZNmDb2
HgjsfK3yQCLaXCI3fnBmIhsAg+ziimLN/bqNPHzCNLNFRyirdw6LUZKVOMbJAzoAgFX1vYHPtHle
tgKfbvryQT2+PfYjA/4eHoJwAjTLQMXhsFfB4hbNOS6THQwWFcWNq0Y1WsqirfiS6Fju4SM+Va4O
uTZgPBtaC6JOOUgDD8DEkpqOF4aTf8sY2d+m0b/fKJI+cotQj/dTjETQgZG2Nac56JYgJOr1tFr2
bPj3F1+N3LRcUEEqDna6lOoVn0ryC2WOELBCWAkCXp8RsLHi8MgEBGcOoAGPVK1OGVsb0VQGw8kC
brnOc0UJ96iq8qpjMK2qbn26k6MVn3OzljBNHuu6VrrsJKZebRoiMDX4+QPPDihNhqc7jGw2fmOz
Kj3Xk0a+LquUGbelC9LFD5Ptm3P5E37B8Z0uI0OZqonSuw/QQf3Ee3AOue5D4GYZlqXtXNyiZpVr
ILlEXr6bfQrFI6nAh1QBXk27DiQIcASWJOWdBqolHKDFws9AizliNdZtj7oo//nsue2kxxWRvYY8
SH2S+Gitenj6TX9vNoVpsL9yTen7l4qj7PkJbzbjbXpcN3DcFB0TtqeIMvF0d7y1JiBOr5VUyJ99
PKyHH0r3YjXFKRV0jRxCVpboNRQ4wCMXjwnXPfalPaRypjCSUlNkHhd/x2uzEpQJNW6/t2eXiluK
Lpd+lh+qaNFB+oXtIK3iBB4DoAYlR7H7VRld5RAoEz3pewYCzCuGKiSVJJg3eWdO76bofjFan5lY
LKtHhbMvtpvI+SgZontrUwT6RPW0p1wWu2K84LwJt3BS2zGVDBUEYAvZ3OAIaoqiJxMIDaaohjvE
WFC3rH/A9FXcrxTEefhUGiB6aj460W4W0wzN0yL83JR/1KPYLTstsiMS5tnq5hphG9zMvf5P+PuB
010Zof2uLz+c32yYe8Vvv27WKs415TxdZmc46PgQDS6tPohfMZkOLg2E246yi/E65wzPNbWOKc8B
lykoKdyFOp55QZxWOLz+MCv1tkbRlSaCchlbnm3DIlw6CtUFZgRYQ4SIXBzxXK19421jUSJuoqUo
csyHfaQfvD9Iw8z6PJtwPmF9IWwwmm3y9ERfgLwHP4ZPH76xsVEZjvUvvKZvvj1PStItJVG76Nxx
th5nhKTni/4KSvkMXxPoRtMCPqPjZDRQqmk6IqfGToF4/57nBxixfQdOTzeCsDNz8EptWmKnyV3u
peKQxivsU46/wMDTV1xYEFlbedxew8sAnrE0Yk/mczK/5Xv7yyFae/q6WqsNhi5wgbuKVF76HW34
kpHS0CdyzIT4cj7JpGdQI9J8u2O3RYmCt8XkX91jEzXlkeLBh61X1vRTZFo9hF20OZg1SvDxu41b
YqQ5/hRE6Y05ufGNnxNftZgWfXnDbIpr5zscy9ILn0l9RUEdFj/M76f7iN9FSRkA7ezkOAINre/N
J9P9oMYhFzohGF6n3k7DaUohuE/7oSVnkUGpK9TJeU0vG0rBjv5t7M8+MNeppcS+1npkpkeAxuvL
dQ1b0ORG/pJWwUViakXFyl40TrXu0h+j8hJJ3ZEnDU9GAg4EPq21uh3IenX0NKtjF+GjMRbwFIw8
UtGbiEEyAJOowFuxRw65RXc6tm8D1mNF6r+UPdp5gU1KgPWDvs+oSlF/0d1dH2fv8uZV4Lq5INQ+
dilg40oJEvlCjS/u3/7N+JULj73uTOlHWVOZmBLGDVYE+Wo0QC1ENKlBdYQFfxFVGozrBvdiStuj
PfhLg2mmE4uzxlypN7NPdMYJUVc9RNAnJZBee3Nj1XulhWl7hOdij72R+4PNx4zPhRFuwomALV+i
3w+JLnDfEYGKPmKDYmRqOeou+b4xw5FYVuLQChYGkQ0/apIZjxUKu/y9rtXT0StJBrOyNLIt5FCf
EJyY6fiPJQQWFvzblcze/bnC7UbCRhIQ9h0JplB5nTUJZIeBe+UU871YU9E5mzNZOurlsTBXR0tM
XxwNdBA2WfvYJj9DZA9JmKwIqwJryfHj8TCfMcWU6Hjd7zCPgdjuVuo9dSfJwKHH655zbgMU91yv
SOdROFcaOw1BqOhSgvzPnXUeXUFVPo9DnDPipL+jIhhWog7XcFXTs6raYkQoAjCVsP17OGmOgDX4
JqaQHKNjuczLUUc6LlxpiJyoCfdjZvn/mxK3ToBMd1/wDo5UFLqBHS0bMZcDIMDX9hVm+4V9EUO4
77MyEuuEx6vWD6XeWbRX1mjxVAG2llLllwQz8SQwXeADX7rOuPLMkUDeNy8RawzMV28zyVumT8su
876v7kOib2FJtnUXuxOGho7NM78fY6dxrR7Kq7YJhAcV1pmrJLh835BHa+zLOZhm+hZlHvGMN15R
n3dmQY6JILENwcTJXELYrLjHpyTSlEYbBXg0JTrplBOo//WPA20KZ37NBuhy68ijU69iZPlJ1Zic
YUO72w0gqhYUbIZuc4GkBbXmMdTw+gGu5l2Y0hmyvOACrhDeONVhekCNBrpjrDf+1UqhdYdK+d+c
Iv+RnEIGiZN0LECCGfL+PCF7U7xg/MAIpN+7k5zZQ75PgDipQxhaUSi1fOuPt0bZI+BH40nj7w8J
QA/oB46GarIVGjsBpajxaWouwMhZWqWX0VejPUh1/gwhxr+CYGtY+8kIpl4tXVQ/6HI4oNUL7tyF
oHuZE6qy5ijC+rRSoBU3CfLggcu2K5MPP7AHwAmozvHcHbIAfUUAAwwPmjJ/afn04qeQdWANOguU
CXfda0jk7XuGkST/DoMrpxHhB4i8EGkrolm4Z5rlOeJXO3abTxJ8ujtUwZDOJp8aVxKFEAz0VUlI
PIT4rjcPHqXC/nLoZHc2bGC15KtCAlaOvezhpY65wZdsyYsszoH4Wcn58lpSVWI7z8Canpx6lqX3
mkvR4B4jHU7kytJRgzwg0RyWQWQinb+5RSvbFoSP0ysQP+n2rvjz0A30n2vyZ53wEAshcGya88yx
IYTQ4o+RHnK+OafSKe8UZGi5SiVmBnkfHEyEjbWC6eGSu8EG16Z5m2uMijotnsX4N+fZZUfK89WU
LDb3M8tcTjL5ooHTMbNs8Ll3GsZz1791a1VOFUWP1EHK1njZtL16yEa4ZQ+PnKqv0bVTZllT8E/u
4koV277GuLc/lg+x+ntkfArNnncMI55TRzFitSe7SjbP73qdrOwYM3FuCFPJ45nW3hxvU5gfqDSl
7Z5l3wv3sykQQkFHMFC+D19RpJLUF+kQSMLfLKrbLYucxtcupYFhjoPdxnR2g1QXbNRx7z988vwE
yWNvQ0PgpxJLiB8WLje80ar8Fh4Ao/cMMP6m4VjWoKHGdCdfIyDkfOPOQYE6JpfQ/J869bDUFKpq
vncwkDvIyPgYNUelqq0s44KXxs9hcN6cWKwbFKkrY0tW+vGrLJf/+LmyoXndx6w0EXr1t0njJVZE
q9DQtPXrkbYh317d4Z9VnncY9t7WNdr7/p7FajD5BgQG7+IN3YGQ1SG8NBpJh6fQHdBJeOe8O1yb
qTWTOT0m+/7BBxPhCN/4EAxTN324HVR0sN2NXWb2/5O9O6tUptkdLliQ3CCoBgCTaure61R3LdyK
UO9+rlA/KVDqvjTsn/PfR8stDTQ4lKmhfAjbzSP8efc/rjybjzeH1P8AmQInOId7oQ095K+pC0pw
2e3HKqewzX7s8BJpAlEBd9tKrHoaWGl70/+xmje58EmT8cyiC17OfsNqefGl1W4HHqm/uVbwn7dW
Llo6z1ebhKoyM4tJSqK4mPdxi0FOPPMK6Pi+LpGF+OiJ+He32FipVS+CXOmspAkxckzYV1h3sKP9
Ijg+3skUecBxpK5i6EnGaixp3B3ixA92uPWHtCfda6COmIecD1zWpppBA+oYloZURXSPMJeb/+gd
F+DbhBFN5/XHFNppF1Y6ZsD0MwBHnTFv7/bY1RUNNWITuPTdpkSb2W9KDIxE7G13ZxsR0wFrxONY
nYmL8yLxrescqWK6EHcZ3AYkxw8H3AqkFF9LD+/JptUN7xJ1ODqLihgd4/Sg+Jyr3tuFOpFM3zxM
RkCSMTPaw7msK7+RfKhdhtV0pX5J/2mbZ+1FsMrS9hfZ87626CGun+s6aqd/LiIXMACLl+UCfTkk
gvVm6qwcqo1ohmTytsN2zH4LLWQ2hbieXYjcmjw+TgFeDtiJukEeBZ/wXxF0dsrjbBiz8byiaH6f
t3ONvAMSrmcBsKQenx+XB/woEUEePuW8UdGl/n+YGo6WBQQpSxr8IuJTbgsTOZ6LWtB54gOWI4V5
hySSNWNGk75che6xiGjCb9PVpnTD6ZoxjW+ywIB/9ZGIIPZlW2LoMzJnQpvhczi/nTKAFK6+YgZc
iLqRFT++Jtnbc/S8DyMgWSY2y6rDmyH0V8ZiRN6x83tZgA2k1avjmeujwtqHS+NyLN+wN4HHUKif
ll9MEAnDmCOU9k9pJPF/8h0LlAxn8XUwfSaGTlmw8putYYrKc5J6aLghw8JFJEqeShjovPMHZn/Z
QBLZL2+hZYxM2T3o626Znb/I7eSQWbzz89y4+9S1GRazjfIHAaGCr8FsocVQlOT1l9fJ4jmQtmFa
z2JgDOqztj4TmR1alr+qZfDFSFr2fgvcYh+5CU3EZhF0xkbIwAdU/hv7v3Z+kZYFjNx7gqw0MOGm
U+GkkTvR/u9rZ/UeDFLxP8AUL5cTFapEo9USP2lDdfYkD8V8CNCwP65Rgz0m2CoeB3sOOuDKlDj/
wiLeVOdE8h6gIMHl2VeqgBYMaL8UM+31+a3qeBOWZYojSKJ26bggpLbndpF2VGjrGrv8Q3YN8Wq8
0b1pu9b1hjLzIEPd74qC8NBjsq/GVZB2DvwiTjdxDjL0p+4WaghMY0XPSOWJaoiF8v+w/EHQWeRV
tutxfnPYiTMeh/Jri5MhsnZZ4PSJSq0/nYlhoe3tzLMEdPx8XL3ALbTzHG5JywdXUThkOrTwbXJb
zuYpAv4HKcwB7cJgjTYkVHBTpfrKLvFgRdygtEDdTVB+m3nlBMLdz9T29o8ddyycUVOQ6V7okAsX
8ph80BgGgYo8vNPcuLZuzzfb06uP3O9fAEQyFVvH0HHgk6iDVSBBTy2+tPpqiuTibl1mATAUdVGy
lAwqZn8yU5GW6h/Vj5GJais7kAJruSL4WYQs7AmVlP4ylobeXzHoRITtUXIvdJoZ5eH0wSA1Bvlv
L7CVSTe7R97CCVFsxjIsOQOlwh0fB71qN9HUoF3mXVH5yeWdhbCD19sXMHyOnqswIQMopu6kwxrI
GlO+2/Vk6/pj3Otcl211YZpkw0GCodXMHWOGy/sSVl9654Dm6P7TL7mPEDlIKaBNxHOsocnq4uRA
Fz6yImT4EHYjibr09oBcZgrRiJL4pUBB5ulMZgfmUm1z2IdlpoHlniwoQ3uAfD7/kVIHaSrx5JBF
J3R+cCRNo9l7SbJ6Uk3jcvpVBWE7GKr/WjLI0wlXQX7PjWOne7gVp0mGYbcV4L87cGebrClWoGuS
3DyyjGdpsWcZM+YH8uaDa3WbFSZ3gR6uHcnB10wt49ptbFJDCtC/1N77mwcM1PJfPDhYABA5h1Vp
HebuxhKKzn+DV7aHizfOzNuMeN/5vITq/Sk7/ZgAnBMlQWfAjGMrPCt9C8xszUDbZd92Fj08jter
sigjUTolswMMBYu8+omJ0UmnUNXw02VeNOQdql4xbeQCZF9x4I16TGKlJNZhlu/96WkLIowy2HSz
/ZjLdgi2SePr7KLTXrS5XaB6csef47g1S4EbDkXcc32VCQBOXvgdgvuZn0tm8I5ZVOGI8yHWvOU/
DenrAklzZDrpASeHZvWTtvpM8tWmrvS8JdoaD/K4/6D3JzE1wAW/h+mSkjzap+smbvLdmtEGsrYT
Wh6kHgd4pP/RwhNaUzU3qB/ziCF7e+RyRnJd4OFN33TkVspZ9gre+SIRCLd7bqAyUmEsmmVgshHk
/HTVfD/4NjmSQYf7Izv2/jIKFS7y4vQfc6V/gVjY46/psM8VJrxmY9DQFtvpKzywiaHM4bHVJUGF
rlEHwJzyOxE0wVq4DQN0S2b2pxebi5y4cDr86cS3C2hqy5it90EnSdzTKoCfsHkMKvLr2tRrHFdb
Tmk1lS3cKx2TpWtluFHxalWT2lqAFjo4Wn65cdDF67xueL07Gk02SObfckPvNDh3kUNmK0uRqW3d
IZEgY7uz1TQ6hRNmNv1t5i5zBCsdXB8lOF8P+TFB11VAYGBleZm+dPYBNWr3d09U/cd0EEOwqcMJ
zUysNQrwiJaDJ5ABklioRM+Mfo7BQFJdA+Lcdxipa/IrLM4a3TGMYIOTI4k9tdMHKUeP7IlPH+vp
3MO/L0HaBb8gH88q4Iq5lhgOPZ+yAuvBro9DPji6zeJWMk/c7leQ2TcouMRXV0RpBMuM0uzfPCdp
/+WGrI76OoX0kB5EeClcqbO7Xk1XlGktFFJv8+3bXHXxd3ZvRDVOarENJ8w8Ckad6P29hR2xYhZ4
nHBxabP9hcq4T00ISfX3z6r4GBKL6JrENdMwufIMISA86VVJgH+NN9Tzav2LI+TByw1kThz45E8H
FgMiXChPbhHBWccj58ICtOwOztpFMtJAbf7mWe4EzV3COOBt8c7UJ+zEe6H246n2T9Kn3tiiCCwM
pKvyx9Trlhhju4TtPqC1KSiHh5ZhqW/hSODHcYk1PmjcQPD5Bc5pCFCB0dTobWP0Zt7ubHUeotLl
dbkWDILkXxSD+OrkBNIWzXJl98ZvDay1HOS7NGESRV+Gr8HAjsU0JHWllrqmd5GCabFkM6WDA6bC
xUwwYQm/xBeA/ZPNSy5dfd3hTKZZVgzENSCOVzvVLgcIKzApK17p9jPLKY1xlFh8Si/LJFUvZIuX
FwmJY0XQQuiiYbSyzfQRpB7AE67n0fbPguqzulfpKFVq/cHKpVsdWT1cMvOO3fDPXjAP01B6Sek7
yYSj1TaUjCrIHhOy9R48tWTEDNXZ9gCBJTWQChX4v0ELocjOBqgPat0qMVnL0H03aPXmDAANt+zN
eaib6elq7ezEne+7lnCm9QvCejItD1nj+GwcNNMGywlKW+HR/MLNnGAsTzw1urSSJA4UffqAdlzL
KMZPOzWoKffwuP0CqnzNNbDaWnDFCharaCjKBVVXj5j+Z53DL+RPfvc2DHenuz1rzDJjTy54eJ0F
Xh4lBc96+UofaoYVtakq98Ta3RdkLWYjFGc3WqwXe8sXkjud1Mrg4/hlRZQjrVAz/jdAIaYX1HyC
pI7GuiXVfmKmqoAeEqFwklmjDJpYpbtoGDMZrCiLevEuxdgIlt1xlTAdzXfdoPRO0zEZNMvXy7gJ
wT8l5AIYTqQY855NoSPEDd+XxdZAM7YVn5BEStGAczH7GPfvGqZtqiien5ZgxMD0/nBsXwz3gfV2
Umje6n5pjPjdIZNrvM+vhZLa7Pul6CqBqt3507XeSlHOnCSQTaArez0XUPONhz5s8WvfIGLH7/1M
5pT2qGEgVgl6n3az6tL6mmX4Bd8D554S+9iHzi2t/3Bdm6r/KgOnVY5S6+pOaA6SLOJ1Db3IF/O4
FZv1/zc6yckrEk0PDV96ic8h0LoAcpKfsolcm1cC7mdLXOeI6eFayy19sXq4orrH18cZXu9Zzd/G
nH8H8jaIAN6KGgm3s/r60CKqqZe18aoDYoaL06l8G57OZTI69NuGj7hguXswLMsdiWpj1j2vtD7I
7gefU5mRUWO+ui32UPafSKNgjl5wwJk+CFZw0JSt/fJxGKVApNDB+eYHuq3Clf6+yy6dbeBdjS5t
bl2CUQEkLzx88x0i1UYvt9zgy7FIMr1OuJeZ6xFoAqlPF59GzP0i3Fe1muQvcMN8YY6/hrSVrcL/
APtFPrG7uvynMejzuSpdG71pAJNKqF0KZs9d4cHjD04D1sH6gLi/aogYhjyf2uVHMfC9u+JrL4cE
tyK79sKIoIpxWry19R3RCmu2nRkWn2fnEMpOixwxETkplVEqWPbUGaXU7oIagvkLqiNPeG1mK4+Y
2WeVLpx2sXbv69sVLZdHKESJ6Ye+HrnKHSQxV1urXkGSJGHUSbrYkKRJtE0K0S8L+dEPloCAs2Y8
SzCJBPICQ3Ogwb5SldFwSuTLt1tXuU9Yvo/33hwS47nqgwMxR8EeTfqUrTUl9GSoaujk081fSqaw
PY+MJkloXKpi+cHqIboSnkb+VzxXTi0h4aN4ckoa3stvrA2KmDf5XZvK9UWNlN92OSWQLIhHRLpv
9WETJgKze9md0mUxikxIWUpMS2c7PVlfUfw3SuguLDBfGLGXDukfny60BnNwj3ZvZLlUIEFZD0vt
wo2JZM4UpEyFWSSm1cd2a9A7j27UQG5hPXK5pPP+yR4d4hRasg1ziyKIvkJP4X/40PT+FIMxcJfn
i1pN8m3ADnBLzG6aC+pnZRH4ODdE+q20+1pOXhp8E7LyGt2YuEbDq6+AB/PSKS7NenUJeDJaGbB+
xgZ1Je1JWkcSuBtj11PCsu8xOp6rDiRxI5TjvVVrBuG+h5ojTVuESm2pHPerlAr40/iUcvr9MCQS
DNvZMhxFYV01I3fsOk5BnambPx5jGWs6P3th/q7Ko/PnLP753VJstAZBZR2PUm9G/0UxHKP5PxLp
eKg7pClyUYFGVVgXLG+kP1hh/pGLcfORvo8GbJwQm/JBWT3DFdRo9zfU7R+SUqJZURJVjruYUUQ3
71v4NS55WCRICVyuPMDz5YMWwJyqLEl34i+wo0UgqiP2QTJZjcqGJPQs4XRy7uaIzO+vsAbUbBvW
xiPzlteB2mR6D4jj7fgUqC+xvWs/9oK4v3th+oXWdn6vYTD/2/BJeD/z3zec6mFKrCbw10nr+FIb
KAJ8hqNVT0dvWMbLPqUw2DlKh62cCA40zQ8TC8nklOhXTOXe75ym5UiPzOMeeTHlvFvzrTdFBfk2
I8mAoSP8ldh3mEow1PGjeV/bdDLvnl3JIH8XSc5vZ/TwQphMN0BrEEvWTyANeX4iVeVCzG8EqOsY
BDBWrQ+XLWZN01rd8itf8s11bBd9IO7DChhIAC7KVq5tzUKl+wUjZ64heX9a4eBg7FR8/1JMpdUv
32QL+ptNha5DKfdmkMCovLgT94BlBf2+VAu36byRo8ntocDZC+32O12cBbUOW2nGbLfYyQ+bD9Q1
Ypqh7sd9rA2g5FqRvqWS5MrQksnskjvHZnpQ3JI3t3vwa7mi5fIS6hZzcw+ujRnjp0D6NapI2uqf
yZUQQnCkqFFSTnb+1TYPnOznX1GGAqPhnLsHvr5Z3GAuWIUOyWU9Of0eR6fqsmqF+EUOpaKxc8KZ
rzIFJ1GBmeTIEIh/BG2JijaIxPzZsgnVzksHWIiP5hkRhwmdMLe/jX46z/YKsipr12ZLxajmh4Ft
0HRQD+GzmsQHTKgY6EY6pfSRqTYjySYhfDOfZjxl27/TtTutU6fpr44G6KXffkjHj7nYBoOX29EF
K388VUFzNhYgcfFh3d0TP7Dw5L0KT031E5WxxAyTAFddKtEUExxSemRhtBRF0G6lAb39B57jocBO
Nf1+Z8jhDnVCq/NPjE8wUGcqrKXYfe65NZAa3bZ9cUrYorSKxlNoa+PQOsVF32eKtIkjzWab8UfJ
N4kZCztwKQpY26R2V9/vybthjP9CJ4xFHxiXzdXc3pC9JbCEd/prmWJb9JiBwNIMA1LWKor+8zAt
0NYj/dGCVDmdsQ5W6ludBIjIKpizXcSw97Y/2TVHEx59jNVxaVpDD7QmRL4B8Nv48rdggxhwAo0P
OdYjs+otJHYzXfpg2iZlbt/iJk7rNUgLI7dFS9rDWxYZaEkESH6qsD9C5PUKe0wO73VWafGn/ZjB
t8IrZc8UfIWAdgxsCAn9kZ6Heral3jP05JZLaw/aw6bdREdeoQ9u9gBC7IRQcYJduV5Ktw3cdhiE
8cDFAYvoGVOJB2sNQsEtK/6Paj26HI0OnCLiR4BLxuf3YHh+bLHyq+3w7tC6ySGSjLjIdGBg9d9L
G0hb1Ef1dY985tB50H1U6RATKaQ/UEdzJN2amxHB0bFlHN/H25TG2kaX23pR4LWI+2LzbQSNg9rX
tNyV0nU3SrMiydveMKwI9I7CdxIZT2IFlmMrXJurOj7jHIrBh3MxUhlP3tYl
`protect end_protected
