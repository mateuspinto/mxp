`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
SqaPmxFjhb12Uh6LXCHQtfjKtmlkBk4hPnLmZDGvyGIepYy1uzw2A9cq+nRiMtggkrifq+YO3S/+
xViIjxL0V6nONRVwzzXfQQFfPusv6ycPM3Yn4ao4MOwGiUlWi7R1pkhGh+breCvqLcJo7Mlyv//b
h3HGMdLylPdvDE5hPastCMStKEcXYnsvbBaGSDkrjiyNcY5u7LDr1EIzDLr6NDV4R4XjxjDxK2W1
jDXm90By4+zscvuyaUUx4DvhiRYaXNVO/zoCU/+eE0QbSXhLx16jbZY0PdcULjiytH9ZsoCJAlPZ
+/F6tzEp2q+88C/d5Yhsy3aAh8lJjp/aG4vK6g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="nnFVeIqCUlQZfoG7tkE9qlXrGyI0Fwn5ly+BvYiG6zU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4400)
`protect data_block
e9rFDomaeNUVfi8S08PRhODZwO0eqRv6teoM6GryHE0XEw2wsvjhEK9U+IgHYEYcKO9PXZi5KDoR
lW4ZWgKaGlPQhmJhExLCuW0hGN5Gyi+DbxwhvLo+fsmEiTiTL9MkJ+t9l0wLjTG+ZXLZh/AY0+Cy
3mqo7UC4El3NeD9un/uRXmAbK1AKQriy4aslWLUhanQHnCP+nP4ZhtFnl+lvVWEC5vhpaGAZ45Kv
xooDv2z1LrXOY6NPIz3WRIgHhBiXxNhNTbVXJiKUaYIw+SpKx+H9axVXw1DXg+FmVTavswjTQjBX
FzqrKTsXVQuvFkOjm4cbXnEY1p9c/FMzkw8w/y7w99GZYqr6+zWLQgeJqhw9djMqDSroY7y0pKiQ
HLtaUQ7jSr5KvAwuXGXi5kPnz1xTkWR8wz6a7eoDvp5sFe1DoiIoOEuIgDV3JQumWotLoCVC7sY0
xobLmX0GED40xxpamYZGeT9q8gMeCRJy5HmVopmeJ7ccGSHmyqyt3xeo9SlL5JfNJ4KM7Y8N4wuC
WNMza+oeIGMn3gKbDILFQuMZ5mAMNWE57JEUtG8go6kyqbI5ebyno34/Qo6XoFkdppyqUbJOsV9V
Kx63/qcDYdIqLaqYLiR60Ev4OGM8NASpHOSKVYA0U5HSn8pq07bS5Ug9gdd26sBt8cIaOeqBO+iy
OWxtNNdkwFuJ/gUXoxDmSNJIMB28sblnj1Vqw8Coz65+RqcCNVBfw4QHBxTLy7QF4AjQafzT33vu
DOGVKiBX6M1qqld+uRWjUC36CF90IHmMFnuPIwM0VSBX1S2jnJAmInJzi+w8RpoIs4pSlYA4ePvI
bR9q+ILFyzS0suy1owoeMkwMViJ+3O1dbtzExT+cJeESi18eL26h1rpBMVJ3NpvpOg0gaUJ/f1U9
O2fZOOAF892hDnnIN8ewhYUoGQjTcu82Daw2iWAv1zUIXx2aOFO4pIi9iHK9HJGlWjAINeAbQkih
bY8Xbm5kVx9CzBWM8nSY+TQkDUZ4nLvtleX036qWUMfrBzZmX/iKX67YdSfhTKqqI1PemPtj5RV/
idQbTcARRoLVVVc4n4fO8fBxCBCJpx1Ztc8Q3tuPAkULeetQuN6El7l8AoyU+SsR2PlwLJj0V7em
QlyJ0v5U9FU/YG9UMUXsGJb8aN3YMFdD6w7M9SGIzwMPAE2+Fq9/cHp7/4XIMgDUP6J9TX2o2bLK
1C7ak9box9g0rCSkOsFSlxXmODrLNc5p0LfhCVSZZSn9B5zNJos1ZaWt8PY+7IEbAzmYDcvKIAOu
swDuKeACoBURUEe067iaRXldqv9A2bDjtcD7t125CaW5Z0kWVNBl4H2pnlfehU1l9MMeK0EEvgWK
rzTs+DzDsAIAHqPLKhX7aJdM+yrVvdrMGYLcnk5Sb4+4d6zLL4zW5e4n1GpdXKdFNmLJAZbByc87
NyOmLjUFdvl4ibuyf/avxeca/f/OHzF1GorfFFGxMB/5awD+FX7wRTYpQ5tN/P2+UrvlqzhwJIhl
b0iv6z3aaqDgjhtbWO1JPDb+rmbZZLpHGuEdwSmlCdFsqTvzwXAIb+Qg4UDP+nHG8b+TikLSlu2O
TbQXzE62LQRSDV3926AVaIBdxvKebFc1upyW1HhlVwfaMbZpmOQDrd1SEOqUMSkei/Hik0IU+ebA
fSnXKIEbVIdKUuktd3CgoD17Rj0ZGatOLTCVi+EJPC60WV3fkKzN2vhWYIkIdJVTn/HkumnOmnsT
RrRdcKrm7Nha4wXPQztxRC0mQMNdAjpAKnrmTAGPzyq7IiTuFhpBP1S9s53OoHbqZ1iF+zhyX/iw
4ZbL9vckyYrk7a+7kUgSjfAkpVTwiI6G0Fj8pa6ezTrruOs3vkYminVWJEsqaSSpj+2WQiIB7cPA
xfq3wWrv8Dkh9/VUN24Tn2wT2GjY3teOYwaXyMwoZH90c12g4ohh9LK1L+cTwk67MtUsLgYpS67/
fj7+Relk3wkW9cDrSLBBlBvwU45lGhZcA1bUemJwZXXMM0IQGW2qSa60rNoZjXHT0FN8N83vkKSF
7U3FzBfbj9hKWpcGfaNXKn9j6Fk6FoM0i4pNofGMdAdR4vTRqhR2nimnrdoHtkpNHLVG6k1+LvZO
E0haqe8VucA/UJWjnTCvcpAUjW8uWtdxZdly17AnVFmOIDDnDdApzuiJ4cTBJuoCrnZyQisSPZH2
u1yed6DgZTHPbNB6W5Hvwxu9VKYnxiWIH5jiT33h3aJ6sXLoPl0uXs/AYNynJBvQ55SUYm+FCx7p
+O8Adi4AN1niDx2MYVc7nIga/EoIAJelPhiL8ZY9x9au71Iio2D5KBov3Adtn9Lcyt79GiUhxFwy
ewQerCFKwYx1A4s9lTuXN+UoMpvYfNrWXK6djmwcWUPtOCKHZuNOGTg8LuHGnNuGygwX268yrXJc
M3olTjQfvYoveK+QVf1paDScD7ulKxPfHxPs2uJy3SbAj8dyFDaRhfD9wTGEfI9pEP1gtC22F32u
QUd1+bxK6dTdjDxPG0/uPqnvJr6k9jfNcod5diGL2bGJCUEfSvBMMMUo74oluvf++b4Sy6MJbOjK
5Cr4/9qaaADEic3XnmpdXWk7nyOoXb9UJ6i+0xwCys1RJx1BJdSnpJ6sj+JiNcek7+UkbjTBvkVT
N5BXY1AMEaIXiSmHXkjX4Zp/vUgzPjNOZv3kMFufjVFaNRqL4dYrhmerNl1Wu1BqlhRHohx+etNA
hNNEIZHqFQy6pqsPvkgkdMdQY2oSozKfoSaqXcxIgzcCYMy6GoAHtYBDCIb42Q1t00eDaG9FFoZn
xeasTRb4/B73UVYtyZFi0hSqk2raJvY7q0FZyI6rdYQLSTmiEYv1b9S352bPTpQbj9rBbE4SmWgk
s+P92J96XUUmhhWYBLx48+BtJ2kSYCwDNn9kjtbC5woorI9kQkgJSeYe12nd46ftgg/AGemNaVIO
Z+xeOB8kRu+dqDHOyZ3OSy6vOSp4sb71qjVMBLjzgec0IMqAkAC+3kpwHs3gixLSah3TJYPmvDlk
VhFOzskZgdRuidoat0dcgULW5fz0mU+9VlOKjb7KYqODZFDq8OlDEbmkzudu65DaBa3h6l2OD/BH
8FYcijxwOpy65EN5HyhmMYsWzRoYW0aQBaIJwG96JdZP48ctpyRBKXRmcUdIH6U5kP/bfqioINsK
Pk2ZmCsOdRN4vXbg/Xieye4COrCKb2/WAQf2Yq2eholPqsY4jvg27+5Sk1UKH83p6S9WiAV0aK0s
b5XLj+adelpV3WEB6kn6x7HhApF5VqTfZoGl7GDVSIi0puo+r9sGtPeqXVzKq6dYlB2mpCRnikak
0oqYNc1m7cEhrJLqv0jMS4+m1gjUerltMZUR5Bj8IYw45nQxOr34mcRQMFsvEG7dA7kvIxPK5kKi
xj77OmVyOB4uOuh6ME5szca9mr0oVzfUV3dnJhMfEaQHZKxkMQaktK9Rog1NHdvL+vSYRVHf6TaN
P6Mna/IF/SMfE4qCTzifLMFm6o6xL1Y2Rx+/uk2CRu5NA2I4NIyZIzySTSnmJNCiGvesN2L+qjhM
rr+BpRYAJwT6Kv2kKwDsS6jJBoPwGB5cSznfiIs/pKZQHdpHg58LD2FvDC93rOkvf8A6FxQZVwCN
MLpoNnbKOpfp9geRslUCNOF/SfMXdY1tJ+NgFNC70z1s9lpOg3/DI8yipajgmtI5A+Qh5Jp06qdy
TAgZV9He5uTX5Y00DHXbftPWs1o+t79cl3h0Oe1zzDHQIsiCSBX1pCiJ5vXCmQ88c0J7LFkbRld7
ekNhwHMIOM2dhKFY8VDq2yFG2u7c00nxZXfUTkq4atC3Jex4aYUIKZ5Dz05b9vT1ERHrltg1opio
kF6VuU+z99QERQjBvu39OtKFzqpSSzo/Ypa7edZFRzXJ7uVDCSFIpQP+5Sv3g71KGX3LlMI5kCOR
ObMG4tAtWV9AKzZ0nBAQI/voBTrfD3VRZ+vKgye46KzbJjwBZWTHBgLTQ/4BXkrkHGeDA1rkLGgf
zsADRDCILmVnW4j5GM+nRrtn7hzTavI174o1TYZZnWFsqV8j8jrFaYNo6eDsFkgqgf4lxgMEa1nZ
4HTTN+2hsT+iK5eMaENJ9M0NIrLPG6TI5PCGjwSL+RgIazQKbhqoadkrP10k65VFXgTPjzDjx4wl
qefwuA5rgikj/cTRDvK2Q5QCeQT1+KZfY/lGxtLq2IiEWSVhKNY6XdF4LTa4sPX+Iivnet6etPIg
YU5oPkrfQCFYHDqVszk82Yrxe6VbX71w7TOvq7gix0RAHfW5GkRmPp+afxcJIADcna9BrT3ynUPX
qi4q1Uh6jIOCNi9A6oPLlp+v+KUKvsZTQbXYbdPZyX/ycHoD+pGJtDC6d+x285lk/9KavveLrdsU
plfLlLL/sLHuo48dG5ByUFUlKRWTU67XQ7kZlOwT9eCXZNuYgwJcmMxwVlpszme5sFWTWxJr4U4a
C4/3bIRCAogSihOPsk3TbSNKVcpAtTvtv1Vin3uDNn3SO/VAI6+QMqCAiRQLIqA8/RSXpAEQ8MhM
L6MlmBdTo+SRjHQWSosBf57p6cDPxJbvL4uynMtR8ipl+jW7GIfBbwLaWOdUQ9OMTr2VvpsCLDec
phA+JlteXCwRzBHfWsQcxd8tYhE8hqso1UJhYOA1aaVp4qW7nnQd5NftolxedOKY64kInqDAjDEN
3BwX/8S4SiYOXMj5GWFSn6FWeaW3cQnwnD4q+gqElb5PV34RtOMT8v/LpEAHlKwtmFroiRDVTOxo
2E+LbOQ55DcyxOjlIHKgy1mcLSwtUCETQ0bCaekvWvq3s9+B29IfHnX5aFvyByYCzkKzzEa6EsXb
GJDhRsxF84p2jMJSFZ15RgNkhizBwQBtkvfQiniVqCd8g9cqd9ZzNxJN9MUFnmF2t5F58m+CbKgD
hIGTmZdH8sDaO18jBQlVBjkLi9+65SeWEEbnYldny7SxI5X7V4rHcjd3+MVNLv5Szp9zoXHSOgbr
89nIjzhBtdrpCzr6i4USYsToOwHOnPwrl+h8TYKAuJx0+Ez23qYew3Ud2mvMN2OuB4D3M/x19O5c
tx8psWtOtWdH1lDQ67Gy6m2BpKOnagbkydvP5yB45NOsjXZNhU0Mzac+1maT4n7ikjnwOi0h3EeH
44LHJOtoi6MOZGCY4zk9lEot0lsK1o1DScHuv/ecn6b6jzZgwYnHjaMmTDrbuRCNrVI01ob92P69
bo6G7n/E0xCwvqWAclE5DpNsRGj5V/taQTJ1MhtACawCp5sycnkRk/piB26POVAO9Nps3L3bT6PZ
+XS/732QyqDQa9+xgP02W9jwA8Bm/tsxhp06UfUOJvl2zzATqdu4wcea/BTXWNihoXYrGFMUaPFd
+kUECrkwiDSt9IbK1ookuXA+6htGUOHx0dwrkoGD+cTSr/8BCFsOtcemBPUIFRHQrRDhRP5BQk4Y
rnTw/KNZF3kyp6qDfGrcgMP9K6lBRlJWZPcyUKx+Zlvdx5uKhXs+eSE+Lh3RShLWhsBovGiNOYjP
UuealegFSK7N2CyjH8xWO96sxxI5QT9ffZHMDqszTef/z15u+C1S/JoTD5DX9p0MlewKwj+BBK1z
oKJxO82C6Uq46M5JEJ2001JkWvkAnE6kTqqsrEXgYO97zFNtBsjVPEUd77GYJw/CcUAzYzDb7+7o
4YiX8r1YBOArn/wJ0ELKjPHBzIldK31VnbSV8jB32P0/E21zjND9wNtliF4h9lLcNehtSfIZBhKd
c4/Dn6AVnkZyMgMLsi0anpaLWz0Oo8b8LA5Lt/T5PapVHx2eLdI/vxqlQpdaOWRXy527+mDHIFob
L3Civ3uf63gQDe4=
`protect end_protected
