`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12176)
`protect data_block
KDYyJ2pCQZCtpXKW3hVJ1YawwIVQMJZrn/PW7zs4Rnhv9JycTaQyWVg3xMovuxLBAGKylT/EYk5y
eP7Bn60iNPMcMPw0KgwqOosQ6mNyLh5FoS4y5J++OEusTFu0Q4+a/FWli8VlhJbq+gCTQydsFbzi
cVqRdyC94vv8aFLwCzcjc8hRKqyIBpTwKpNTRd4sR/AeMGe7idvmuxWvg59js9p0jnZ22oFJ4XCz
iJZ02hAjikfQT5ZuJG8VHZDUVeF06OoLtB5a6I2uaDo8V3ybOnzvu8YWHIKX54dsmgw45ab1/HNm
IWE1aC/K15iiLzlQuhITjIqsgeJEHxNK/in+5fGH4HNty3uUXTxZx50+ELoXKP+vj16+eDLc9JwK
Dg7dmsrmB3+wT2AZV3tHui02/T5EP3bTRZNJy3ECvHFSGY7Mum+ngdQTNdO84fmv//Ni1hlWmA/G
3cblUqJjjZd6uvXf9u2ZktsFXT1WIiS98tUGFOAzjvPmpSALSEzJkzRLpDt9c8ggKNI+9G5mR4aF
h0xIEFReYcXLMsiK0tg/43riy8dxIvwZB9yA97Em0Gw9OT+SZYhreXvFHuGUiOq4/z6hINz45ao1
00yXY/VXh79WnIJ3Xk7qjTX5Nozfni+FatBLTpw4G9Qq5L+BPPkfOurQLTez9rhJr49Yuj0sGthQ
0fXJB3tAfhzthjImt/6DaZDbcDPX2mF9aFV5hTuCcLCRS570obGKcUw0CuY3QEcbFHsrzGXC5mFd
i7CkB/nk3U/MK3QrZ9+ydtm3kY+pdzxiSB0c3CKtyJ7iAujA518NjTEfBXuJ3A0iqhl0neM8IXMd
Z/prhYh7LSyyPi3OPuLduMo4nJrcRlfJiEeCTW1yA5Y1gXdTNF6pRyeDtema8IARD8x+8rE5I7qe
G0MF2V5beoMSJYXpaanrpIqxzNRBHev0i/eIfyK8rM8jldcpOvFJza7xmJv1rF7RjgwNjXaB5ZPy
QwpaR6JiAjSi2allk7a8iK03iLL9hOkTSn5LyYQ7Lq4lKdrVeBqgH9kJN5lFveV6yrwHhskDqJpQ
vLIdzDD4QmGrY8JlCyRt79w7naJUBPpieZJnZhGuCGZCIQOMWsMscMg8uDELVw1js+Vjhl1M3Xxc
IJ+/MuOKO0Y0z5zFFTrHvG2geVYBdkVgY5eSM7npYFVZ9YJ+ALk25hLzcMzc9U7ev7300xdYSR3A
ZO1C6lpGZZOw97HNWty7f6naQ1VaTt33wG6iO+qbzMIeuaoDe4X7CDb3Gzbl9L5Qpyf7swkcZuNC
mtJQIKeVbEZPyA8nQA5OY0Mzeealz9l/CVUq2F4XlLYRvfQ5HEi/JDTruZDbMqlrfE1B+gl4hpEM
iAaR+adV9BqAkzZHEFMjobqCXY1z99bh/4bw4jCj4uzn8vpkTcd6KxB1sUqU4QKBxfqeWYarXSyi
F4dlOBmnqz2l9k7pnsIdS8/woL4DTw4LsnOvnevkThc9Kyrf4ziByLegiBoWurthxP6NZjWd5bQ2
pVX5mIBTS+FynCUpbKCidV7M5XRIPEiZvvaykFGkG6PS1JNV6XO14Q28CDKFNupArYdoa2vKcjQ+
TSw9Gx5XGQK5v/aERpKnLtjY94wb2qlQdehdNSoCiFKWU2PKiCT6/qnc0pw9ZpMXcsas2NVqpOV5
J3GD+NRexS/5FbkA2eqpM8LL/UIvOu1A6W4QuPYx8MLpGwSovPmrS60V+0GEBl0EEeNig1mFA+0D
QIuO8KiHZ8mWmV/b9QJywN4icjRkcHoaLVKQhwQSiIO5Uo/02VEUC3R36eb/E/7NeKrtqc8TYwPB
IvJdeA+kNcRyOhDDEgPsU3Um0FMDYfnNogcGWf6CHnaZcKEPIin55XTnKRZ6lFbNFILf9d/7w5C6
+aywNq3Xfl6xqC5l9VL1956go1Fg5xK1MkB3QPLzwhjUCCqr3PQdQG9fXebBPAHiKJAumZ6XVout
luAVohf5kcPrYJSrK5c4Pme2XVtpOqjugrbldAdwmpysr3xlNVKyme3m6HRXHfLCgSn7Qdu+72EW
m8bpCLTmN3o8fjgYmiFU4kyFYu6q1blgWftXVJitjgVhXOiNaZ4WPy9CsfQnl29VvZByb2jq93h7
iG8n3LuQtrz0S8YPRsMx9NEKdPYEo7SHMEL8399T3Gg9JD2jz2fM8YmD+IoSX9yKaUdp4wrSSMNY
7e8T/tEErBNrnLGAOWdt8EOBkgOnWjZBgoxQpcKXXuvF9N9UQDNPR6AmHkpKmwf4ti+lVKx53lpu
uw/3dmBfp+rNAqVl6YErM7VjnOf77fQKehvcXchAcDiuL9sf9J2QxbUyts11vehlLc59ypPxOvzB
DIs7okbVVJXfzlE7P8lW5SbM+hwVNKurkXd0LR9a5H6cttfjL97qM7tY8Fq4yPImnAZik/XE4bcJ
EzLr2wXqvjrGF36Nfev/m6A6Otar6hSAMzQf/8tye/tDZAZacc60NJE7pAMiyaIoXcCb01YIl+66
0bwV5r1e5t3BAQWa1SR4Ys2+t8SRGIZGld0mV99sYVXaLe4nEx2Jj5Znjqu0N31CnXaXK3e2wWR9
plIBkw52yiOmUCB93G3u/mYEG5NtcX8dPPkCl1/4Tyx0PckSLVJTzlJ5Z1oRATvyRHLcVOYQyryh
CpJm5OMF+Df/1CjmxFhRaSzBFa7BaY8xm96luRBEjLF9FY4gg8O7TaAor/9DxrQTuvboOhJ4Kofz
s7eAHVv3kuPP7rzitMMg/4YYk0WnYNDCOv6tA2883+ue1iBH4xrBN816Jn0Hb21KuiMbBT1PKJ2E
94TGTCitAAU9QIrzQNvG/jCWbKUdsfhEqQmPqMSKxokCJBHxYjOqh0I0fSolh5KWdQ3Uz23GpYu7
VLn65ILkqYSHc2XHPUAo8d1JYVdDssNM5HYvUJArpHkaKOZJYsnfacUrKt2mW7nvCJaQNKnKRqd3
0qWUwDVX3yI7kfm8wIC3A2qJzQ8VesyQKa0dUirf2lWGatqvPMo6WVXjESHkxMylB/hb4i5IsPIJ
1cJs3nn6KwM6MZXuiD1mqHfmYuAxKkZUmJvS69cLj/qrl9RFn/1mB3NVj1uKMw0eNshKLXXHspBo
1PDf1FGdmP/TBhwaVzUnvPSX11PZC7pzmqUgstDf6o53KQeDhF6xQPoxHt8wcUOSYazP+OjkaUcA
BN2thF824WMFkuT9v1fJaI5PfAEZ1j4YW4cB66pAOMZRLXudQtjeaGx7DnM+C4t8AJSYIXdnJLnO
SWyRLTvbBuNjKBu0j/Cg6NdEbAH7ItZ5WMP1vCAm+YdS4S5VbeHNorgJRr9543LcmAZhbv1BnHz0
XFw+jp554zRYL6HS7gBAu7wW8tt6ZjS939iiWxwC95NgRohCdvVwaBuiHWLQFtZIyVpaGueEtWXo
TgVgyvaKJ03zL450ncm/Zv+t4unsBGZE5Ll00W0MzVtt2emnGWR8dY7A+a7EM3VY4/VRrRaVtPYp
5hA2khRPwkVR3Wkl+HbZjLnL1KKjGLhWnhs4a5EXFfTtgdWT88tPQfx2OH9yy03pqQE+ihIpWOhY
Fj03+HgOTh1OHIhw+zGr+AlWlyevunYRz8F+zDpr0AMxZ2XYkcM8PbLtk1NTAp87Tg0P6We2iVsS
RcFABvWQicQbNZpNTM00kTtbsSxmxpM15ZroyFXvLMB5gb1NzQz+aVn8rP8CCotbC3Ye5VZ2fOfC
XOM1G4cR6u9LkLMn81s75p3SBrWe1eZ46PDBA9DlKNXZ2d3E+pMt7zbSqpCo9g1Jc+mDuPCG7qNq
qE5NFE05cs7cOpWxGbtr9Z2HF/0P5R/fv4x2TQ4AOJ6LcWDSKBQY20+vSW7r5Pt0lY384BJZS65Z
fc1jlsFUaCEbHZPWIUOMnBExMxJNNvDMPZMxcaJcOHefOiOlsNRG3VG4GjXg4GDtC0OCsnJMwA0M
Ubd0Xc0tBxRpvS/6sPGLJaRnt7IpO32eUOTZoZagfR9jkoLVmief4XVmTWxh6mKz23J8H1WHEUwU
jO380eMxPlBaAF0vSo+Jo/RhD3nKQipDu1jFBM2DB16F1gZyGeYqtQjloFjZ3Mg8QGwoxJIBAFTB
MFdk/IcsD//U0/TwDqIFETPTjOqIzUXMjwAI/BxXjxsRmZYPieJ0v4tYOc1Hqk+hMrECLPuiCysm
Y37k8Puovx/jUp8y62J6lW386zoYWD3xvCLy3/nY4zBj24TcpnDh2FW+lidVhb3hFepjfzQ0xliV
dhxi+bkmA/ue8ATJ5pwXbYuHDopdJboQf6fr64c1vcIXUKQs5rWTZqHNpjd5A1Eo1dh3r2Weclx/
CzHVAp/k3JN53d0ConVkht2Onl6+T0gVlfK1gB3l229MYwUcswMdTj9BN73D7skyfAUe2IdFB1Iu
8tK994HdJfEGk56/LGeXK23ngzJi8H443aRMu1Hj051ufscb+FAqoTGwHM4DIKvGFGL9UvyAn++W
I9utzMLyVDdImYUNzmX+WD1bOXP9kLiikr94BbdXiVC9MwgBI3sd2TRCvIvAw3N6tAs9HGJU95eT
fnKHrT2vBXVgk2/W0YJF0JHuz7ZrsJMHvIiVHcgJQFLZ3I9PEA2FhMwHBQNP2+ukdIG/0Df0mcHU
WeKR3G48Lm8fCriq32NAUfURFWkAFdfUuOuESRKx8YA3GZwSFLLMHQyTZhtElQVzEeqOdF70f4tu
b/8zFRbo6hj7RF7qjuvBTLGmYKJgNAQ9EA8g3x+qYWflD7GahRIVaUGC+8xpJGdCxvcBDXx0nSk6
xixIM1942GsznqOTulKfRBn7ooUAAkUrdg/xtyi/zVwgpVL8b3PDq9YIjl0f/x6WoVfw6jpdJiDd
LGTfVtLltSzf57oRxUJAn4aQn71ifJyF6tuSW+2fLjYyJifZfLPe2u7CJxVtOk0uikW9ci5yHz5t
S0EZCr9HFvJtV4nkvfBDUsC5OVOadbz3Y68M8N90WEpGTFnVi6No06R9XQfgwaysCIwJi8S2BAGS
H8ctcmb8K8XMkeYZ2Drc+cm5FDYCcfC92fOBrK1ItGQAa4A1DjAt5MTzXFC9X/uz+sflW+svbfs4
5EqnZTDciJyzgTd/aOEEFLLXcC3C857i306eoNBUYVZBDgMWISO9i8UJIkqs3BSXUSLDV9eclrw3
xhqngvmkAD06D4CzLPAfaHiAc3owjMNDwom1JxQ8XGYWXCs4Pt8C89VuRg54g06OOB69akvg+0Qs
rhh3axqFtTIB5WwLeu058zCE3At8MOwF+uBIVwcw8i9anlF/cB7azneCJBNIIN1zvNl9VCiWhclZ
oRcXCHAc8P9euOwz0YlMqfecd3RaER/lrZMaedXayfD5ZTk5TYLinPPG5bgza7RwmtDGooWDJBbG
FpELTjW8EqGa3miPNe9o+NzaonryRJyH7Mt9alac8Qajd+OaQoE0xXeR5AgknZD76WOJxqaev8TI
1F2/TAlbH/0Le9qQt8eH5DK4ekhkVRHtbtHQbSjUDN45gRcbI66hcF1L4+h0TzjXBOh4g1YoBjoU
y0iOM8XTc2HsUgxmQTDMmH/pabhx6sgYK6MOstb0DYAkYz2UTm9wEdERwZXbb0vW2RVrKTe094Hs
Uj7I5eE3uLHz9FDcAvH0uvTHQ3nT4kNZaKDJAUtrDRpv+OBS9qVUnvTTFX0aAco3vYQfhSA4OuYq
ReMswWrQY3lPRapw7PM1vd0T0TLdSvy4R+6JkEj0wFjfULv6XFhjVcSl41D8Ay3x5nTKLuUu89yO
rgT9dSNzFtrxM3+pc/rt6b4paCR9cCnpp5kWsDvMY9YkowTJ+GU4hei92s8zOZAA3cOgoUbUev9F
3HZhf0xqnmfomBkvFExtw2lIOvryC2mT/eOmEUjZ+Hu/XYsBe1kTDJ6Doyil8GdQfA41nsoBQ9EN
/VKGYfsySF5e24ioB0aNNpyFQ//DqXYX3FG0DKIuXNkIikzTeQfovddP0ikSm3eaYSJGizRnD/O6
VNfzcgMMjANucTAjbhZM5bzrwbnocHwi+rhODcA8Em0/ZM6OMEpO/Wn3OjAYgTqhXnmyreTgzaDc
E7rsSQGtE/fuyXF+kZ1jefk+NmJkJSZNzPO5b+uKREh2uSrEC0XVEGS6oyEs99+YnULas40oMTW5
4a9MYMoSCpY9oaxicWLF3W1Qj1XnLZlGiIwSgmoL/RQNWtmrwFvtdBU0giFQZiO04OU1CFb9wXYF
f8C9YCWGzuF4f9rGQ/unZ3vJbV5jWxc/ZVuhvKxTOGOTqjvEMLY/EcKB1+kYtTVDOcNlKi9tWWib
mWUTjBMgceXQLBZJ1IgItrEO3Hwd82K9LWNBPmyEejPXmymZYEn4O/1Bq+p6EzZ1k3C86KMOHiYg
XkQ6k4LD/ebnJ5zbvm4Oy4sMw837kwxAoJQ2mYc0lb6lN8vWNJOA3h9+nHTnj+OrHQzocbDhSbFE
RcCdwaFPoVFstYcH07rhqUiyy8825RO7z+j93tVXPJIedUUlwSVe/kJ0+y99CEB/cummxMGBNyos
0QfGdCF6SACO55QghTt2IZtpYxnCHtNBH2nXQMTR3bDX7sEaA6DhYg4fy2eTjRJ++wZLTKmyCQYB
HYgpu5XIfX5il5jL/zojBwG3o/JbASqe7eTFLkZHRMBwNHi5drzdMIZ+HMSfe+aVTkOv7keIPQEK
8dhkA20pjCwYoWXiWn7f5kY0od/DiLaQ9JdWcEBVLWgz78XoiGFBtfAJIbmRNeGW4ibQeuwrYIhQ
9kvLxVCdGmtUXEybbTE3pbdbNNJaqup009cLnBlVNfb/HxwEAVCxRn0fp0FF8sAsH0EhOj43S3jj
eel+F18LxReRu4azDNteZiY8HUodeCVhjjfS65n8Jiv7OyOar1uJcCX5jCrXyyzvsDyFfWd/FBwa
a6fyeK0+rW/1Yq17hoG6yJOhkLPEhRwCBik17E0bFqKz7EdRdUvdkZ8Tgl2nmsRvMkVZ0SrOMWAM
wgU3aWgZILFsq7Q/p9iKTIpFqaRhGnwAVO/JrxsK00EotyPSDEbjHCQuNJy/hqUvAUEju13DV/Bm
llRsLC2EaDjTagncUlfbGXsbKH+aeZ9aWA6GDYza2BDh3+Dv4L7Fo23eIXo/cIy8K3T6M0FscGPz
xOfVDo7lNqvC080qmW7y/sMjnfXHOPbQ1hPhby5+aC0TxMzqoJpW0HXn0ftSn/LY5PQnDLCyKjMf
SiW/CQq0FXfIY2rcoup5Y1xvMx3/yWbi7ebVVR1nco38JXOIRY7v1jzXl/WERoNSVRqui03F6OIL
do/IHZEAnKQTg/RNE4GRh6PjgY+WXD/JxIvWi4KfrSs4sO+FDA7A2i300Ojpuz0Fs+vOs1xJp0pk
asgaiHP/nd6GfmcEouJiOsprj9khp61vTpaKTEMCRBK3Sc+Hm8TqxpFe4717FsErRlwWUhjph8ii
nkSq+AMgx2D6EUhi+eEwrcPjJOZDw5WKaIkDfk6+tbI46IXcDco2nEtLMSDxd+vT4zLYaCZwHZrN
T02rgADXzpY/9WZXYeAq5Yt2sp2wFIgNo/+Sn4CxYOYxoK9lIsLgCkKDI7F7C+QPpMkMr12kkpXh
idZLIyRKq6xNHwp+EJ7RxK9dUDC+j/PtXZyXa/gGvaO+dv9HScou56te+g51PWmsubAJXpxc8HH/
R90AaAEgWmavky+hphnQ9uAAtFtFRt6E9A7voNo5vLgkMfoUwSxkZt3BYgt8P9PKDonOZTOQWE6/
331IsKWyhI9yYey8hJZiuTwJVrh/lWU78hHKsfVGrkAXlbm26QDaqWYSEdWrslM94tJ/U+TK5uDl
F+Y72/anJOxfO4ftTnmwArsPwAZ+wysZmShZwcX5Bc62Se38tkzOcnJLlOMEBZHNvyooMrrIzECN
AjtPS8vz5qukmWqp8EglXvIKRjMD4JoZAFGCeSqEq86w3tXLf6/XAPlto56v8TBwD6sNd2fr/cVJ
eAoa8DNd+CXDfFxhnBlQXSKtPnXZ1GlWZiJ33J+HxY69g+oRB7hTtMvLhNuk9VYkkkkxipqPXd3/
Be795XMkscQdnDBYbC73+iKZtcnqlawyt5nwp9P+qzslJ2XxRRxyCi1vsqJzbJfT+csszRXuLDdb
iOEcf1vg3JB/pM4HjBXxPOzyW/BjerywG/nkh47p+cuT8Fa1Y2y1A3DZk7b6TMFIUAViCmlz7AYq
U1YaVI1Ya4iNKdwdBWWlcDROF/NUfq2GaiNCiSelkuHYBo29zHZfS/H89F+Ha0Iu+wg3pBAfhTMe
gXGDipHYmSMn4D8D4c7+GHb9vDNC7/V/rzGdJ/dwjxuSWTQDim7c5kL901CNZfFc6elh3/3pAD+Q
BTN929oqL2D9fy06l1DSlA9XJT+V/uAJsmw1eWjwi5DD0qnAWoHyi2YV5e9GEF8xGkZAA/nwM5qF
eup11n8qhmKYBCgAI9d4XS5SbvMDU2D1phWitANRVQ89zyfbGZaPr31wUeK7Ql3eO3RCPQ+qGQ5q
OssBRBdqENKghqxptunDG3QHHlNflZveP0T7qS5TUP7UGi5rbXeLwnqo41rK85wLC0ytnESzA+hK
rO/8qo0SeF66hTZ6WUqNO4GeWOPQIMaV0m339WdMAyzZpQmMDMgOxSBOt3dttgi20ThHmT/gj8aY
ZDFJbR+92V7uxwvPGUNGxplZxfNwuK/l6/FdDZsIQ4fc6h64FkvjjSbVH8OoAFfSqHmaoSo2fpEL
Abu7s7AnZM3ztHUO4nL+JqrCzB1ZIx0AXRGBFwb05xHihInw3bonX1fmmwU39Bs6F2Vc9pzzaXYV
1KCNeMkWPqTDvrRejLTMrZ2oQLaZ8hiI3KZM21s1wl1vtQtvUvEu/gJvTdm/FCKZ4suoKGzhM7Dq
03UnAbbmolcnyaw7f7yqWjE6/H7oH8wxaqs8Wls77QSUtoErpJ4tOwNXjoOr9SRbt65cXP1n6hQg
iVOHSF4eQsXWfp3gC5rwI4iPzn6EAwWOdkUe8/zehUi8MN+ns5BWzBBaXlnPcHSb1kZjBUO6j92J
kh32Hu/zcHDEa1YrtQlYf45WV4jJbMf1UUi4JrBdvHuaTSGLIbGB1urcfpMyQqw97Hrp7PHaWVOZ
jRYwFRo5ZDtI2sp1uhqKlx90IYPVdOy5nhZ+PSOiay2ARPATKRHLFhB6EVNJIohkcA5E3CMkVCYI
5YcFdNquh6jGLISTuGE6xKR7sdX77/0goucdw/4mPK77NCS+tqR9iZeU0P4PTI/9KtwggRh50xuZ
7lX09PvxF0inRBkbutUyuXP/zca7g5ugKURTF6Ink+EBysD/19ci4TM6/JQvJnn8x6mh37TCF/ww
V7YcBsgNQ7I9hS3fcyj9YcTQVBoBv8J4hdILq9toi/3bJm3VAFKbQ+Ht5ZLh26rKtlMcbWXpT6A7
M3yqcnQyGAywAoE6C0EK+F8gpnv9hix9keWDFeV8y5mFJmEtVtFPtZoSo5WV3scsSMB/twTEMZDf
r+pMUvMcOsY9sLZ/Z6nREWkfqf0oy9dOn06+mZF0S3QN+c7/IU41CZKUGPrF3LkmtnWlDbOdGpet
QoU2UsvVLqVKEB17oFdlRVRrI8XXlEq/J2lu4eEYfIFJ3EclmnNOW6Qp81mfVNwfiPAAA5lmVzCz
czYuEDiHK+SZYbCXnc2z/gnmlNL92JHiro4wnyQ7Vff+IfhwsHeg/PkeeGq2el0n0RA1kUkHb4h3
/UygdKyJ3eAO7VqBpkIRlc82orQVibc3B7dkLrEh/b55jHxaL+KQBou5J8NGOIeNEgPKd0L0ly9w
mW2XFPf5wjSVUOZtZc8h+rYIMGM9HrhtnmXRQOF1Quy2QjqYCrAfxL8C2y4Y5WvbTz67/MDuv9pJ
UA2atvkqFHNRkTTEJaIT3ndmzegjJ9049ga3Qj3WpFj7uWtdC/lIkdUtqRi9HkOWz4WG/P0bQLEb
WZr/2cA80rdYqHoGrdhJ9ZAZnWa2RVL/zfvqJwjqy+XRyzRqi0djPj8FVYYQ3amFX3XEMmCRuSiw
6VEijE3BxI3qPxjayjYTN95+akXq0M7FvngVs7iOhxcFB7VOfVO1cZfGQ9KU6QFDgu7Lkc18FxJi
+JGcoxYK6s433TOJ07PSaZYSWfV0p9183OSblP+iZzbkQRUyNPV3j2O9+gGxrI7wt2G3h3I1cPPG
CISxdwfhAmSzNW2esaN9RT3hRJdF5ExhEy2Qe4jZRcoWPH14gS8/vmwJhS6lRwfVBUCynj3kPdsq
Tmud8Fne4Zs9Ix5Tfrzjg7ULFO4O74316dHbY3SuBivu6VkQektSSy0qv6K3/4gA4kcZ18CNiAS6
bCo3B7LdTZSF7Yc6lzNbF3+KeW1XPofAVYDg2leQTWh/ACIU0GCWY+G8nWjvsvOrdUfuVJNK9Gga
dZHxGaMZVGeegaxwirjSjBFyeg8c8hMQ7j1uYjYNQGMEEZ0v5ASKWpsBdp9X/WzG84W61JZduSsb
YNjhrn9qaSXddYgjD1ZP6Q57d9/yEVUf31jHtIhSO2TUOtVdcX0QmxibxG3PrgtEKD+VeNbX4eF0
Sz9lh2B7NPl4WywPLPcJMY0CY/LbEgNOttGVv4eSyV5YPfl5SL01rQFljjjMFwCbPBSPgPOHqs5H
Kif7NvZzkuMlyvRNzMvkD8XU/697VjPMyfLjwMFavBW8gd3/znXbxVv6YHBaG38Z7D9C3dQOlcMA
J4TYxL3pVmpxbsIFLYHunnTq7FU6pF+qpVnwQo4Y1UPBxUvQHkUw/dbALJ2R3jU/qaq35JHjE9Td
q1H31ZB9JkDvplZqzE5hwonpYKRGJCV8s7OsRF+SodAiehtN84dLjv2+XHjURcodL88hTkpljci0
Sq7bqA+k1c791blq9qyfkfwjixDBC2MICEedaRe+EOvA2u9aojwmTWq6sSEWEOdzGidiWyZwdoSi
Nr3v8KUrAupKE0K5lXx6ePazHvC0qM605rwDQe9acq1a7G/cT5iAkGlsZHMlInVEscpd+bFm27OX
0tYndYR8hZw/emR4WfYLndkvqr57tTmOuE4PNcrEr5SK4CGXLkb5uSLXn/y3JKP0x9fOJl5fpRTx
GS/R84OFF11mWFa2y3zT2/WETFN8XBh6Tzx912PV874QPI09DVQGj3zXtz1lZFFDiuhmianrSVON
uALJ92OUMBIbw+xHw7b/NKroF3/1HRCOGfH19iFoyYtiVD2KvfWe9REvQkFALVZh38VH1wcVNSVR
YFpxuADjLatE7WI9k7H6ottKphsfxJl2rbaRya1VSp7OUp6IAmhY4Mq6gRMbxmLL+T2MsI5Kuy7F
KrwoEHRC4DLikkb8nT2s+gWdsHRJ+UhC1X1pctCrSfuGdSgANfRl9jSdtt0dbLZOxqhKGoy0tT5i
47PZqO6IGAwWgwRa+FgEW92LTkSBVtU6hr1TNfY1seElaZtZLhyLhgP+kwQA26DXCsDPdlIIJYqL
ynCgFgOUmUpIlW+MUGEOQVu4NItSmqy+92ty7droaakf59sgMqp5KSDHP+XjXXuenUmeAvU8OmjZ
AJV+jmQfiSzdTRUqMY/rNuNMt0aKp8zEusnVK25ME9iEy3yKQ1OsRGymiBlzMdRQcBdRsdumTtNz
W7LcMQRPZCZ2gAOe8zLyLJ7UAJqqCqG7aUVy5Jt18SFYCvlAxCwuAGbrbyJEVIg5jyHxEx8q87Cs
5Im3p5VXDnAlnNs+/eWI6hjXvSOjGhv03OpL0BGICOzggh+l4pDgxCmSHwAlm+ZYS9zZzLCtcfrK
sJEjTqcCZ/nJN1o0JdxYTO376c8Wt01m/jEMprzMGbzW44J8T/F9v1DkXAm0VKXCJvhPDpuEJZzw
idATiawbuYsPWwoha2v7bZ4w4WpWgDrRSTEE2Vf5RFAKNOOymfDEl4Y6KZSvVMKXerwnJVHRmrmg
WPpJsDcvBRU8MWy4l0gAxeY8KlunTmFSpeHrQGtG+/nEUKFRTCPG7jAnpRk7UUU4V8d0xkvCz1i9
I5aN+nCfLm4bA8Rbg/elsG4t2A9p+9BrZM+fZOYRaLRbpfQPG1cxocxaDjh2tn57yypmYC8LIAmI
ZbpBs7kr+svsY8KNkLi45wQ/Ne+Ndhal79GoMLcH8Jsn96V/cDecbFOozwpGvJ9nsVgpA60xwUhE
6dJW3bhhqJaHURJWRF86mZcGYOMnV/77B4MT2V2e+URb4ZMzCMld33QTbrvYmcpvpeyEgfSfWy/i
s0+GgNBwI2GPbv+TM0Jsv2dKSsWBATX3w6qOYr6UdJudvJcUUBT+bJGcj8ErqWyf+KW2qVoSuRhI
Fdg3MQocaw4IgH1Qars5Wx/yAtmc5R4975G3ORC9QL/o8wpd9TizdEhSt6PlJInXXkaTj6Sk/WJJ
r1ninBAMJ1p4Mouu6lABCIijRPF/6OXRmPMBFWztpfEwW0MQEtPWj/ERyTtgjhpPt4CRn8bAy5G/
jQTdY7stXINuv3a6x3g4MpogoqN2vMpPzDf2TQnI0/9m1r4ACEKMsIQ/UnZikw+obPr6WO/PNiMS
lKoq6b/7/AqPxi3LPpItqmjuqx6WxmbKbDp4r5F2kKjr67MBNryaZFy+SXQkove8ZNORa5Hrc6hu
Wq0ax8ccpf6/QtBrT5h/TZkP9yGetfEERdOSB3X2touEf+sKOdcJhx52UbnlBr7wbSPfPdRMrz8U
j3twXgomYJ3EfyEplLChvjN3zqau5+h2Xyo8FLFUJWpRO2V49SXcNaUevHmNOej80tMvwODk6NzY
NMCdhAMsApenNduhsNTyUk1VDP2nLXCV66TO0mZmAx66AYbiARjM9p96DjHC/3IdjFSMd1orhlbJ
yvtpxRqMuDw2iAHhN6z8MwAYEBvRw3W67wrW9QIA6PCYjtZI/WtLOwsLUushnPBRoRK5w3mkcWnS
fGXxG1T5KO3F9Hq2vf0WIOBN7kvKw/gHxQIVkKmNCLGUY21QS/0haEbBEgySST+l3puH3isAyAJl
VY7Hp3livL/sRnC3ftiKV2mshYW8n203qKaLmivW4wJ+YOwWCLeNuw6Aw9z4KJoBwbn75p2pLp9b
+OpTPvTz/1N5D3oI4MoUpbYgys81Lp404ZNLe0jS3BbSMfq2GgEWcV8t9lbSJPdZSO0XGSmUYs88
6/xcCJzJmjzKM2ZB7mrgoN1oK62virCpJYaAuyJ6elUD7yeK4dwwZFo5YVwV9Je+Ea4P8QqNVWqR
jSXE69QZcGAaGp9yqn83VSYJ/v5Yeq2pCdR0qQ3kpI/4aCFNIouI9IX6OuXxP3Rd2QMziyDqkgzv
YE8AMiBVDXogEr3bd37T0CcgA7VuqfVE1D3v9z/JoxxBzo9l16vH5QH1pYkzOr3Puo8PxBrfyJKE
tkJQapq3CvutbgfL+CI/C3kUVTOG01oGpB33LNcqXaLTGmnaJNLWTcgyikKp+gOwA20yuL5kGWls
n/VbIjSd/wGRx09SsAg8wUZSh01v2ORzC+THGq2pcmCt2QVlTcv/YdDhnXh3FjIuU3B/lK8zsG+B
dvqFh+Q7iWas96gSnbId9xCg6RUhoC0VoQFAIvS7VeuxIstJ4+HffpEN1cyXImWBxeRZ32nbQhDJ
U9PrjP3YYlLEuhrhaoFIKlXwX8F8vxUibB5cDmhDzQhAAauT42dHae8yO0eQ59FV94wYf8QVOfJZ
eRsWH9GjYSNCE11VhtlqgVfCLldkha/D5ADRuJXAwakKq/VsCn+FtsJVvacFJSdGNVdDn6YXVx9b
UAdNjIlO2DF0E2JJKvSgXUiLslbXF1G9f4ebdC+3Mj1z20XG+ILhd3J/kMbNzXbe0LEbkR3g+Ii3
kQxOwtDAvK2lP0lHGMdrGqGmu2zAPTq2zvqrW8+csyHMmLeJtOKH2bdOcYMNVyT2FJgFhAm2h2SD
nhR2WNpkwDUTwEPTh+BVcObQzPLjBtbq+BjPHpfBZMd+VOodR/ePHJ5XWBK3At5QtivfREGtffDg
EEX/TQ7siwFMwtrwCeTTmwnzdQxEdjkyCAoBNayL4IKLNTijYcb6olD1le/nSJ+1nVSWNU2ehIRw
zgwS/vYcLNBVkzUh9gPh6/2qowdxFb+3VSHaya93bsF7Ct3rXlsB97sCJnwHt4oNP2BPEanhjOoZ
upv1lDi7UrkzJl4Wzab4c7BF/vbF/Egsvp1vieM3LZ2M3gZa5fgq0CSTb32CGxPBILx0MQqcMTK9
aQFisxh+SbOsx58pZODdgHINaAZnAAiO42DDXMubKGjtF6bZM9J7pSXGDBDEtP+Z6Se3sHdg3bIR
4Ijo4L1DNmCeJ91ZlTPthtBsaGruEcAoPjnPXGbRXCFjJ0Nb7UgK6EhL89Ev9TJ4G55y6uCK6A3u
UGmLK7eOZz5T9Gyvui1pUoTpiv5YDx2OVj1PPmCJsaLPExgK3pN0HNpNhKt2/9xdZbg2T8vW1YBH
KN9EZgeX+orTJARkKs4y5xn5Un1FldXW9/q5Y7cdr1rcZ3POGvrBev4XPMMdSJTFxQKfa15jOvnE
M1rj/c1yqez7J9JpxMvGak89Iu2jdzg9shC3s7eZEPzQgIaSdwH2rpm4Q+kfkMNc1KT42erSEIZV
zR7ck+BbyTmfSPNslC4TrGFP9y5+Jspa+yrUurnVAYhO4s38UJNdtHPW1ciJKTlF00dhIpNKOm6l
zteAi8YJahRNEcliskED7bHM1rcZhK+L6E6xX9BebLiw5SScjGCxDsiA/6QOjkkEaz7jkPmAQuTs
Y1q0Pfrwj/LOHu4HAjRgsSL5s+ZnCNwsp4CPgK9tUZDOVQfE1gpmHGQhE7QVJwB4yOv75OHDlcpn
w63maP2gdFdnh0ylCXRVb4L10UrmsiAehf+L0eSFgrmxh25BrynyKicnxmnUrSJFsz9QbVNZ0dle
9GGcZ8BUH23cBzZhpGBJF6vOG24iyIR2Oqlk77lNrjQprqjOil/R7nmkLRqYQjJDjdnxMDSHEeMD
7PFsOfWEBxy6NWK6bq3rQOZQfY0FQ/+LqjWgy2+NIvQqdAPJyr02qlS/ZgUE1vWWtNxPeU+bYmOB
LbUKnkHX/dItrBZtqBEf+n05uby4j549iyxcQuuPtVNAIah7q/bmLpMG89xO7knD/uGW6GghYAUc
D93SEO4A4jBQQJXlcl/Sx4SVYBluu7U6p+n/rqHlmMYTdHgH+8cbeG8UHF3C0pXft9ENoSkzObTU
aZvxoO+2X0uaYx7YuvE5DgW4OBK35cWAA70dJkL75Ro4oP9r+3/z3Q+/U143GTIxusCxX8C5eCpQ
Mx8MxaQlika9g39oISRCO9BmkWPexdvye5P9ArRQI/PYLaMIGXMQDfPrQe0q1fomU5ttnTc/0n2p
1h1aeHQaQBSoeRtgWDMAjQrP6VgLW0Yn6ygcQyBvsx1vXWdg9+SBhlM2LEJFymKWRn0CH3Jo99B1
SpitGLO/dw0z1xR09R02aqgMwOQZzo0IAL9TiZ8jURp1alFYq9Skgy+vdbbaCvi64oTKMDxX+I7P
EOLCTy5+BkDPfUdQ0rw9MNQQib//b4llPaCYRQiE/RXxEP+S7GoD2tPcNbQ9H98e2Kd7bMDthvZs
VoWY307oiFRbFUss2+psJW7RFLrmzxx/lJNkF6cvrYIeKT5AuzANo+lhd78LbcYbUpberlcboqB2
f0qSPTVwkV47e1sxrSu6u4tHoL9vmpPQJZR6TPZFBdMrKW1wn9zyyYBhKpsvA7eXHjaqBQj8chZp
i3COBemACZBzEVvLJCV9Q54JZPDsga3i3lUhFu9ylZv5VrafiIxKNvPoBrZ+m0L3PRe6JqFrfxsw
7DYdQ9HVwrPe4/khMxCee7aT+CLpt5/xIW4u7AIkxKmjZ7WK4dGNAIKEN2U20ljZKjc4hBwLLSLG
Q4+Wh7fSvCf9NzR87xLBlFYBrU+0xhkIrr4H7dd534yL0/hiPtfhApaEy+FaDYpoepc4dRjDDedk
bVHr0VfoRxheLym8lroHgYQ/pJUCrjs7G+NlddvddM8F8o1d0LDKQIlqQmDYGxEhFz+cgmyjObh+
xOGysuFnnyc7PCmQpLs5S27Gz0mSISaSWRXL+s3a/hSwgRaEZaGNUlxiRm2g6DQlbRB3tP1/uTfp
9FvlpVwZA1YP424VHAYz3S9opSgIYFnqNYsjnZI3dWHoKjmlLyMg/TF1LtGdC0hZwt8G8chVvVBe
AYUJbLtCZ67torzBVJLDfcY4tLUbTup+z2Yd4hF9Jet1XMg=
`protect end_protected
