`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3664)
`protect data_block
2GcQmZczwdcJOC5nCc5SbvFyT/GdJwKr+MDkULoAu24SxuARarmTCMaD+q45wc+vVfd6JzI83iWU
6cy+jcniCNQtBNJZ3K+JEC7WtBueDGfLKsgheeB6w9RZODcqtm/is994WrUQSCKM1bZ9Wkoo9XjW
TrkAZSyBw8r5Fg8+oqBk6gxG2A7ok5bFyzwtjuVdHkaVX9+MPf6OeUAD2HnK0lS0gedWGt6+7+z9
9WXdK6soS64tzEcN1t8D72Xv9nCD2u/gMHkjXocKkYNDfh8ki0tSd9bLGp+of8X7F3BTbPKWEao5
AbIclrKoVDYqQ9NAE8Tg7p6K0bUwrqJqKk90RIHP1GgIp/O0XjQofCrG0i4YPp5/L8oAnKpOzlly
5N+AZz6n427duuynLuo2mIumq4W82fRv6WyCOk3JGQqUCppbs2pp4PmSlDsFOJy8yka/WLdO+OHn
kXGNeEDAAm2z7dbksXi/A+vnlNaTssWEyPUO0msc18sACl2vbsumjN8aCb5l1ceOi0JaPFnJiqCv
a2ojTzzB9w6ZqbebxbkO6+Cq0PBTf8dDXd+MZO3ISqmHbbSVKc0kr89PoVL4x0Z4VZ0qo+14rHe/
CdHvo9KfMAZzRkYeFmMDlA07/QcLM4pNTyd6UNy4ZZz6k5yQlnjOczOR93huUnGZXjxIubxdE03j
03SWzLFet/hMWUuH+Y0LQvakgfpnRIvFJcRjBu6qbS/iyISKIa5/laq4AlI0xMBTi5WtMf0Jr66u
m2sltxtWhoMm7fQzlK4lq3EK2L0rATt/vKji0hXBnInL2MLD5cEv9ajhCIQ4dBJ5PO5ZNou73+qY
TgTZ3LzVUyzvjfL+WJUH54PKEQfOhjh7LgVIO9LUCR9exWk74jNtEMA+062zcMiiKCOe8mvzkv9C
d5p6Z9SvTtt9B3IzN6uA1Wr1QgB9pCenuRzC39DZJd+5tWWzu+kL3LKY+QNDm520oeyflrgap1kR
9SU1khIbwMkznCIBNdo7m9xQ+6dptgNc6blyPNSdJ0ZE6ivN3cfv5sh11qvGcpwGPv6laFYyfcP+
QVlPCr9qESjr0gzPVkvO9CI+w4mVomGKTPgs2ZduAkv4Z5/5LmsQk1cYdWl75Ci1w94Nc5CGT4a2
YkFCPwuHx2eucokgyzG5WhHZMoxNY5uSaDl3RKhcJxIC3uIUO0MXE71yw2IZSUzRUI7M2ZE3XA+4
yjmR1g3rIx3FAQVFnwipaWVW+tHTbFIPWeh9P59+N3dIdGZ0fg7gegSSoSFHpfpIeCwcNdGAp1qh
a8OQsXgdg7EUBmy0AV1VFcvg3Q5fy/A38ruXZ3IUCawQ6te0VTUqdH+9Zn0taCfhkPnmG7eIMx6c
Lu8W+fhai3w8EwYUJB32+5hN92UfGM/+FzBtztG36UUsoVYKna/vE1QeWj2rkBV2Kc8qbsdOT4kV
CuwW3C9sM09kbHMjPxaDh7yDhCa76Ip8YGA0v5pjbe41n1KvHghFrjuL5Xz19rVoq/6U7MFSuKsc
ENcUGL4DoTb5mgnnk/njsEEz0DI83DpHl4fdKIu0ykrS9B5Tvk7JaGGnzO9vyGpWGJ1YzooeJVlR
JpxedgPZWvcY90V7m6cgThC/OYVECf8v4IrRQdPDgbJqUmMs6N7vTmrREwtFiRg4xcjYT14C4RRi
Yt47/yLqPVRgW5DPnxB/6VukHpCgYASE/cwlZyDVmnd6TUFvH2k1CHR4FfNzLFTJ7VRa41wlS/4P
ntjVoMDPbA1SLNSIOkd0gGY3sC7fCdxoggYboYFOemzAo+IebsQ/8jr5e4qRboQUokiqEIX/JlGw
/wrKtyAEEldqS5RAtyyLsLn5SEa11qjaV6K8xdMxb8fzYg+/S0R/C8qbhROy7L7/4oFk5+qWu9Cd
74/Sm0aaZ5UuqvuNNOH1xI3B5mI15RP2dCk6pg8/2jQ3cZu2si5lkFDB45nXgSS6F9GzhkrCJ3CP
br+dHbFDLwNDIHpzBtfW4sNF9dmELQvNKBaWYL9G59mXDAfeYiTmbjtSu0eTiZ4WN3q1BIONdt51
7R5ORGW1NaefzGRyhBQpuVvSL464o/2foTqM9TOzMaiMqWfO4aeXrv8BzQhaK7teGthtrQmyLqy3
O/1aYfSF/K0KwjEVff634IfpJTyZbBkli04Kh2lSYfgxqGruYfQZnc62fgg5TWUX6gcstg/NPUZV
KiYvOijmiQA9yR3GAjgsCCTzYs5lNeasPxRTnfY2RBqnjynAEJfcKos/GS7ssF/24PV1oFNLG2Ll
z+TDHvUaF/2fG+yAMGw79jXLsYnuDTzdQ/13fjdjGI8imAtHdGmtQfTCpY6NAKZ733qJ28LZyMjM
4EMBtBClmtQ48400xAC9VM8wie9xljxPw/8FmqRb8HSiwc88eSJ5j+6vjXRBvY9ZqnIl9nFZq2CY
sDpLYQmTmsnpFyoyzJn+xZRisMHUfTaeom0x6sPkKbZIW0ln7kt2Lx2HTDngMqkWcFDWj+4zCvHH
SKCbgXbykYcu/VlQaq26GWQTUxyHKcAsbcEQJZJF9YxHjsGQJWtNUkdroa1nTvEU8mT2Cq2khQSe
jCG89AylN7/wd72hdD1ElSh7aggN1Vtn7i/hyurExVzvenoosAgbYMQzyTtQnMHtZU2sI8MSjrWU
rsxkh8OqgzwPgI1tX+9LiTIMo2hT+fEiIbDAI6sLKBe98N+b9TVCX4AJLJ4o2a3henzuNganseWN
opHsBcgc+Rw6ohUbfzhRzICJBU3mdb3gMsEVT7oxPBx2dAsI9AFzjveUOIgDZSNVZRuOBxZpPyBp
PmWMEirXJ/tmbAslrnzRHr1HCDmrm+sU/skl+7wYzi1fFlmgZrgJNCrxYwikAOJxY0HNjRdj8OVh
a/LqF85MewkmDtGCNjZ0rQduzbhZttYm5byfgtr93DsLRQD7rS5xoecfghihpNXWPdKYjAEbtRSA
ViqbUc31ZUv0tlktoOX8b5QZ3ZqU7NoXeJg3v0ML8WHvDB97P9SsfW1imVp6LydQ2mCKCtrN3Io4
BpoEY54UGpC6HKEwVT/fU/GYOx4uAD30FkCbhJ1gidJ2ZyeMyvo+xxWO4YU3vGWmWMjDXDn/e0eU
dDMJyvtZ4VztM6xjLi1BcLMjprxF+zgQBWDz4j00O/x1FyYHI6xSLo3NN5qlVLyoH9j0z4VDFk9h
KD+/3mxqkVuK6DXPqRxTZmBNRjynd4pM1s8M/fb4MLMHsjytcOn+niZNIIKI3Gzj/lqcpX3ziOAa
e+dIWEXanrCDU6rrqOVEtm2u37Ik5Kn7WeHkNz4QGOLibBYR+1lkN6pmaZXYD5c+XcZCDFktxIGy
vmJhLkCINQLGSDYIRPlbFss0lc74dwQwK8sIUUiRMCIlmH6yKeallEh93nDbyYcr6Ng6nMMJvpcx
WdurZHwcPoRDHGPM9y3HHfI32pHPef3vg1PO7RaffpbmF6LKavs/G64Z2fHiQyTEHNDAGU9vMAwu
ZSyJgR0Q/yVqQxvSyxOpsIh1Y/5ELh9Mg0AQKCwz3o4Vi06b3SI1P+YwbBICgznOKO5ynvlg845g
dehcRUZuNdKzXaoHOYgLNX/NsXCtEXaHg/KkUGN+EnsMUkKldBFOxpUILSBsLDcTKMFlpnDYCdE4
y9azKtAn+eSIA0spL38M8kY2zTHBlr4MI8fmyYo3yvIXUQrkOLQq1PySt/kdn6hQw5k8fQ03lCQ5
GyfebuxVm0489pLzfz3aXD40rUionX2KwILuoNwVowdrzevRKvYHT6xOyjhmvQnbddVbzuSNcn8k
Mh6QwmVQVJygL4qivzcXg8vnFJ5z9BztlM+3BAfWEuzo95OX5TndwMltI3YH2hS1VHpTezxdv2as
QVOZkmxMBJOG5O1cfbjVWmpMkU/kYxmfVmoHFVXFtd0hKEzajgiw7lUpZUG4j/NSdl6D282I2eeK
aWRxMsUE2WGdDeuJYC82zcR5E3Gf6X44Xx/ln5yBJKsIrySdxueDDDEI849PkSZANfY6oiw8YB9V
OnD1XAt7J+ANwoPU+8QzXv8XBVHtXKGAgOXPYM1ALlnhsmizdKs/swVe8CZ/JU8qsMpwDLzjrGBX
8eN3hJg6OV84vPHshMHcb0FXob7yIXJkTiDV8fK73mFvq8e1uRGM4axfU0pVxjeolPlBZwzOiVWO
+V2IE8utAwbkNGmi6jpj0bByknKmT3CB/1+56x8tawe7f4zfr2JCnr66HdIkTHFQpHMInt+3W9oE
mOUwmm/7ArWJYHDuqG2FGCgYzeJtbYLnMLpXtCZTxImOHirzkIlBLzhCLEcTAHmTV4zx4txnqSdh
5C2g6ilhcFE2lwCA7/7BMJylB5OQI2JxfFojapDNpYZxSrJUY3TitJXoGZk9UBbwYtLHC3smt718
A1Stup/naWGwn692hnArYF/YuUaIVeHyFy9eICgzqUaJ3jCHZ6zDr1ox1CQtR5WDAcG6fh8aWTOa
VtntvwoVzTmEO1ZHrJYClkBnu15dmA8SeCKQwWNgb2q6XwsMbXPJj749sgGaw90AqTewIs8F3sen
E5Y8CS7rzn6uwHT+DtVhPp2td8cJv3I/3LGi9TS4Q0y8Rjn8lQkiVFN4G+r1AyigtYxLSShTC1go
dcpp0mvNSQrbREN/TAitgqThq1TEEcUjTB6Thv9NJlgw/euvpbj9IiNQv4fyneiwLvinhUW9DVy6
ayTTDs5oX4kkwEb31romg/hgNkAdv2vh1r9oRKm5zS7Q52pC2r9Yd5owDlEH0QToELQ9vgHyjRdJ
4rimERtXLZFcme3921pr1eIgs1w/j+Wks/FnKTwIBO+0BZCTszIXlBwH9QPJ0SzfmK9Er7Or9Puw
Qf+uhMP0wfUrfMFxpb9y0Q==
`protect end_protected
