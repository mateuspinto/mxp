`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3488)
`protect data_block
0USWSUGxovGsyBJteYpEoUYx+W+8OX955reMtwHQKo0oK+uYi/SCvOqjbjZf1cabCguSTFQ0aXB3
/Ovt8NP0yaqpypNPBcwg8s/4z3AebeFuSgEIda/cI2ogZqegaJG2FcwZiw8tABUSKX+zGfSy3m4r
1dVZ+mAb4/rTzUsMmpEk1WPtaCD34ASR2Er6IGLdv7WbJpS3VtpS1CXqM4RVJSCj9ui7l1ql1594
O5VcQMRWRgMsgVD8MYvoVZ+NefnmXGGw4kw1m9Gxg7VaBq2yvQ1garMJiXnLS5KVdEQAirwzYEZ+
Aj0QHKpjLRjIDu/mmv9IolTBDDDDpU9MFejSGuaBQpHMsJ4fCtWNzNbDGFQdfh/IQCKnmw+F+ipd
hDCkaGWiRKC4Ns672o98spUxQKYCrLuICgcg3LrL3pFyB6JIG+MA0iMIM8ZKEWXHahACgFB/krcg
g+hgJnniu0v5y5OF177h4KBdlrPd26s9+SryDuL7XSvyG7EBLGCgVC1fN9BogDBS84gPGQIcbhdk
WV66oibxI7O1QuMjJemN8fhDjxhe6NkM4iMc3ESdPIO4Eu7OxZWWkMRp5tY+Kq2lWHyyTFL1tpIL
wt6ysUyGDIcOTMIm7hz9LPHCDXFy49Dr5y1+nYKStdNHAahC0ZLfiE10G1T7q7Kfd/Y0BAYjJaM/
na1JmKEwhlbey7c4+6HmesYcZ179OHoJovNdag5XxqbzFPzq6i69bmZFGp0Wmntb/YtyF82X3rG4
41JqydaBJdEszA8E1ElrnAGOceUEkEdfh8s5xYNXJIjM/BHEeXMDgWNuDJrm9Giftn4ElOVcE0K8
7aMsIW1jXXE11NN6uM/B6t/8he+XnzSt1lpNizyi+r7GhwDqhOwnHdpBkrFr+6FPdjFauE/Z7vJ1
ygSVtPvlepgBn8RSzS+f36dc9uIlEEvGKNDhFteKCzQK/38R4ksmMZqWh7s3+qP1Tq/OV1BuXayj
T5fz/V4CpyrZIl7DuseOn66RmybgpaiBj58TWyATEuhv3zRF+xB/Lxw/xiORtCIXUEZmVx5+Qga1
0s0kbz5ZrDev1DS54fSHNk/HmzULfSfR2Admw6SjAEn+s8HEuiaoNbDnNCvFZveE9diW0E0BPHPY
qm94ByVGhQa3oJaqdqgyZO11kisD0vbkAngcEFADFD0LjW+Rqr1SpevDLfLebiwHwwnznFZB2Thn
jASU6VJfRZFN87PoJraL2ZXhq1GCRr6eODpDAVrZov33yJQQIHD9dou1UXTPv0eipfemrEspe2cX
BIlhs9zAQMhI1y/HyyVyuN927Mv0RfFshLpsMsfiCk8/AXRFYypTiGU0HloMh/5O30idmJhoVYCV
PYDhGaw/sMhYMJ6WXy3KNnSQoWVPMtTLPpL3+KzKYPVwiHAknixpNdd26All+a73InIwIacJwTaZ
GmdwEC5kTsvziXtcT3HGoC9XLn49tIUQbTkASTrz97+tjSnZt7vQSUYaFhHy2iR0Ft0nl7pcW7/B
91IdhyKrpfHuLpCWzaGfiku0oYsfUjHuHBgA41fNyFMiBPzMfeWsuWbSApZsVU7GM7pB76DHMbi+
AEb+c7oB73/6XmybEeY7GAwZhSRyRQu2Bjo2mTbRLXtWrqV7z/f7lC24njA8maoMw+GGGFiHgsRx
/BBQM5DgemhzgvaQqxq31DePImefAi0YD+7GxcHgBrdOKM5xC4QjibxHRDTl+IZgzgv5ELw9jBjq
u/IQIg6jqQ9OFcdkXscUCf03ZjIUR8zUtzAL7qaJSEH3vZd/3yIXYjz/3IVvn73awoIUflpahOsG
BdkA86kC0shYjImZ683HIxlbiNCKx39jIkqXEQe4uP/aJ2tVartnd6LobMSDWVQeiZJKfdSf+hZP
z/an4fib+fO6VBzTXjQhk8m58LXfVIjraY7PsV4p6vBG/4PcuKvdQGwRsHL5u68TLLO+P8Tj/5Z+
SsEpYaXpA2Q2l3BX6Xlos56nvRRudJQxJJdm9FE/dp6OF7v5scigFfE/eznuZ21OkN1lH31jwbD9
wZLF2UpDql7expMcQk6+FrE+2FQOSBEk+2JRRwqkwCs0xIHWV/YGDeP22WOdiKYWuNoowQV6BXEi
/t58kla1Gh6LgZlmo+z9jddjagiendp0R8cdN1YN/v6tclkkDJKJwS69RnTVlUDet6aspkEmSGG1
RYVtcIJHaF5YA3BHtoatbT9xOrOqm6CUdGC3BJlKjeUrqSEy6F1UYcGj4OopMbYPmdtmmPyOQR5U
QePh61/1CfTR263XkiN0kvZHP8HzBH3jXN1E2Xihr9SKzAtD2Ozz58yHXWt5Gc+UZt6ni+xHpi2n
tfOxlZ5rjx9fSbNzRmAhlyOuAC7Tpp9gnIDBhLMg8bNKDIl3WU1S/bk4DKwzUbpow6uwQyHULBvl
mTki9DIKJnEbg08X+BLovc6/doBnK68Xmm+oaMtqDIxp2yafRiGExhFh3iCvtrgHi7QkLM9Qq8rm
cvVJK6GlSIHg3AtWqBT04e2szfARkS/EKOLdDfz6JEJ4nB2k3NIAWQQfC5lNqQ12WFaW/M6jP0IP
wcUzKgU+cx+oLNTcXfbz7nRKIzlMrgn1M/Jclg5MymEkuzR2EYouyrooNtg0e8MUUu7JqDV3Ty4r
4vfp5bJ5YAGPJccdwz9UDHqUHY3Rm7nbydKjQjUQpzan7LDX8LUti41P03e/KduNRTOKfke/DJK4
Sxm6nFGOAchNRlgHAjJIZUiIPKHgI7yQzPyLXU4O+ikzO1Vo9InPkSwljSbfDyfwRHyPOxz9O9Og
dhs+t4nv6v6amn8WgbqQ8DPdkt0989nACXe9q1tK7cpCk3c70PZmAXZkreBlG/iQmW6LC7DX8ySP
qrSNPa70t3kjTTveEOTLfthFOXl0qW0DDBhHK1Jn6A1BJykMWravIx5f6MIkF2AIVYZoKuoPoLxX
euSdM7CbZkwRqj2iR02dwlqd+GrQFT1JiqWLwd5LX/xeuEkNalrD4+NyOxyHI4cfCu5pRCCFOglX
VeOUncNbumo5dqC6T5vNxOht3kW7+RfcpP/qMapvFXmITMi47Qmnyr3C4j5CWWFvASlA5NCRIrBy
dAvaq4Z9AGnv/OibjLgAAuY+r0KNazfg6BuduBjebp21SKXxAw8vzv3+4r8+O4zez8ohbHyubb3w
hSAOZmW9mA4PnBL2iPPdMBOATyAhAXK9bo+PiczyOyfOYoehVbeGdT+OGhjc2Y5vkBDw2/JrmFhX
1H0hGvfSIWmw+RQTH4I43T0JuzV+hQ1zBcS9G0+kNa1QbWIRiWBnMQyURldFG+wpKY8+NRz7p0BK
Dg/npcKrQqa9DUXnKZanj/Qfdg8Q+rSZMlkclHy/CHqfSua9SZX5pIb3xy0pVrXTW0GsCuVt68c/
Wz0JOdbTgmBhjBTEFlzViCGIjPGCqRXZIR82tqIcTuyFwwIjG/4ztMHdR5DkRSeysgzopNCvlIRE
GpA9UlAeYd120iy28g3CmuDQIfvSu5rkPaa5f5UnjhlAvDM8nW4e5x3bQZKRxneCLqh5ofEnWIHZ
VVdboYbwO/k4bUnWOd3POcNtHRST1MgX8Qswg4BFQ0oy8yo3rXFW5QCCR0FA77KUXPML8sP5AH42
rnXgXcdJArPCmKhYsPCPILncpCyWkhpu8xR5+B8tw0xmdP1cMpoJA8EwMzILZczcVxoGtUZBqUWP
tLWsr+OleJG6xzxQDUndlI0oySfDGQoKe/cs07qZiNINZVtuOBbE1ADua1VieK0AdlfGxaQhCWdN
KehJd/6JVvNN7ETt4lTbqDGV+M1RphGx7eqL0MBRqbrB0qM6cVAoqkSCOiTLZW7uFkHkNeaorzl6
cQh+OdZPu9J7IHkEdGzMY8JjX/XO/qfV2Ga3ewjBlvQvho72ScfssKna5u1y4nGIt9ew/SNSK30e
QirT2BfxqX+UYOA5T8e77TZT/8sPj5Ew/sFHCmef3SfbF7R7vJQJz7MiOaskoGQe7Wzw7uF9EYpV
Fsdtm3EiJbHD1uaICgds80ZP0TWQENmrR9aQiEPYATv3W7NMEvXuPuszaqE18BDCKsRGxOenTtt+
b9Eiq0Pqir6C3anvuweOsh/n1LC2VGg0Os4ArvDhzVzfEaZj/1d4NbA4XNajd2iDvSgQMJxCo2fv
MEqTMk+LcZmSwlKndmRK6uq7NZXxC7ZEXpMNJFLANLIQejk3wqvz0MVi+4ZDTK7mXoBXLbhsnn6J
ArW5ptZlcAcAgGV3R+jqrGWHh1SkazKtRwwLGItUztLnNjKW0p9qdRreogKw/jdFGCQeUEh3HtXD
f3RNZcEJJ8Zcn5MiVSJjSFtExyavItqfQJrS5hBEpzRBMjt/lGqQWEU8OibFM08fkdJNm1lwgEwu
VGj28Vopd/XaK3egZKKPn5ThfOyIH5hhCFpyTJUo/ZOkfTpzrTNuoK1rdYd2BlMat6o/D+82/aq0
CXPRiqHPay5w8dkBFYhmtP6mDN5NrpIkKmi/YjgohBVqTVbi1cRhGGQqJaL0M79qH4xlUOQMxSgs
J2qKw53TZgk/b47wi07J35HcQLqnRXTcG3M11rvI5TJfkV3mxoVi0tgOgyn4oBiIzt0KC+mSuSVX
1IMxy2ChzxsOqlQ=
`protect end_protected
