XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������r�!�:�;�pi��C�p���xY��y�DOY%��F�m��HD'�ҷ{��wȶ*!Ϗ�b����	�껀�<�_)�f�-���q�an��1��0�"^-���S;y�X���(:�5BY�" �m~���J7�߻-�B����(�m�6*�S|~r��W`�g��fH����Q�&q�<���������j��|��ˋ�fD�1�3���Z�=��b�@T�\�A<��,��C�� jM�� �}.�(^����5ii������X�d�l�� �v�]�Ր���m$=20Y�{ե5V1� �q5,�
�Q�kY@_�]>x㮙lTX�+�EA"-^Y&��0θ� �4�.�T�Ss��A2��_��N��zO&I��ˀ�`lj�D%�xG�2e~tQnBέ�Fe��S�^3{P�&/�jJD�T[T�dT�̖���le5#D �j'�!v��8ӓK�eQ��{�i��$�#b��P�>:��H���w�R��[���w3b#�ʗj�������T�1�>�*%����v9{n�����������wS��ol�����YY� b��������*5�%g0��Qb8�s��VSnUc0�1��2��6�H�/Vse����s%�$8��3,s)��� �!�%�t��]��'�W{.>/q	��<$��*�^���(1}t�D�,3�_G-���6ۺXP##�iR�/�؋�0BY��,I��*�մ�F��9���\�-�罿1	��)k�
<�Y4;o>XlxVHYEB     400     220)'��+h����L��Ho�����6\�`�Տ!���k	�@	(Ȝt�@>����"~8K�@-���H,
����"p����W�Ս�w��ڱ=��N�R���CF�0uYD���V-s?�(J$�Y�����y+�ơ�7c������b"�q;�H�Y��/M��%�#��xz�R5*���џ�5�������Ctf���/]�����Y�]r���|�<�OҼ��Z�1�D��WW�U,���R1ɭ�����|�hિ�q<l��z�_��F� I���u��z(W���h)5c�>�z$��5�;1�Z��:��[��U������D_ dl��~Rm3�ځ�}�E��ٚQ�\��#஻�^����%5��T9r��C�O\,�V>�L?M9G�P�ĖĞ�tQ��=���7�<���x�V(M��KQhk��a�N����G��,v�s��">'8YVq��� ѣsQk���A�`gPh���V�D-��8$9�&\0��9��0��`�T�K�&�ǏOyY"�n���b����a�XlxVHYEB     400      d0ep���]���E ����(w���aO�Iq*�� ����V��;ۮ+�� :@��^��6Fs]�r�y�W��p�#4yǈLHj_��_�����˫)t^�j�y-!�_��@�r�R!�c?[P�@�;6w�Zb+�|P�r'��؝q�6����������.�Z���t���DH���@}D�-���1��YR���:-� �� iXlxVHYEB     400      c0r��,Yw~�b��v��o�ۓ[O�NOI��[!�����׌�]�Ӻߞ�twq��O9Y.hh��y��5��#nEl/�wi;����]��l���v�'L�9%b����[8�`X�}�(Tړ<���;�����LŲB�^Ú�{~D�y��� Ѻ�(���	v�OZ p]�pq��RU���WN�5`u��dXlxVHYEB     400      c0c6���ན�ï��ߒd���2;�X����=��B\���c�0�ݗ!(���@`Aj
N �ۇ���`$F�R3�mb��t<�Q����MxW�N�M�m��������7SI��<cN��ZLQ�D���1�R�ݩ��l�g譅u�G��O"����sqվuX+���uNs�ɲ�K�&�XlxVHYEB     400      d0��=oo{�!����@����;g�}٥5����W��5��{UM�o��B?���~���OF}̵	a�>Jo!�G�Rŗ,����0�ж6W�uB̌��8�Kԍ����Q����CCw��#w^��_�gd��ϢB�d���>v����J�k�I�\.��mc[^c�%*V�n��{�c��۴̨��y��'��Y4 P^gZ�Hl>��XlxVHYEB     400      d0,�p쀏��=�_�ɂ��'RPu������(ks���}��|�b\��'�*]{��@��CN$�>D��fx�:
���p�\9��=��Bǡ�EU2���Ⱥ�|1�f�\��Yt�fځ�<
5$��9�=�4�&����~�ڊ��%? �mu� b<J��D
���r�Uv�/=�8���2�����I���}*S��`���2u�<9L#XlxVHYEB     400      d0g�/�z���lq�����Fa�4c�\1��.��� �x�c��j����D���-�؊>8"]����Iw�BC��f��S�Vs �j���]�8}�
����s�0��p��7lM����|J@vt�2��C�`���n�X��(272�>��,/bϟ&U��2M���ַG�H���)�d��{��M#<�Ux��= ϻ�- ��K���zJXlxVHYEB     400     170�	%���܈v�,A�@�%������t�z�o�&�QKl��8V*�JA�K��w52�]��<��ٰ� T{����R��_D1�#g��_���/A:��#��X�m8�
lh�$Uۅ���ԝ�P�O
�$'^`c7��e�~v�ާ�䣧���p8��S�Ɲ���k/+�̖Frl��?I"<o�f�%�.C���2���J#7�q�Cu�����H�,A :e9���}�c\z_���Ix��b��E`�w��E=�u{0ܻ��K�<�����V�H�I�Ο>]��4^*6O#E_"�&c>i��Ml49�����x���\-\�p���
N��wFA|��Y�tM�$lm��Q1u7�Gb�{ XlxVHYEB     400     140K���z�U�&\�+��)����M<!}93����A���$ ���h��q	�+e�w�)�b&Ö�}M2��!���\���,t������)S_	i`��!�^���YC�w���PN��ZD<��`�
�ɨ���(��2��7�J�����#�H�g��N(�9�'�L ��Q�
6 =!���%K'L�4�P)��pn~Q� ӱ�0f��b�~q^��ߨ���<���T���a��ݽi�)�h�x4�H�yR��}AA"'��H�4��s�dVǼ�I�$EQ���6�EI�t��w�e�HЃe�Ϙ�Y ��\��
XlxVHYEB     400      f0��h��Z]���ܲWb`\X�t�i��I+�\��U2��l�|1c4��!r��Hbo%g�nP��Q��Q@HA�.lQ��J3p#C��2�_L�
z�M�,D�m��u��#)<x��\�p�lp�{��O����/6>� P)��m�)j9,+���)��&a�pX�˱�|p՛T�y�Nv�n��%5��,��Z��޸�/ɆՓ�:i|Z@ʃV���Y����sI�K IL�:��B�hz;�s`XlxVHYEB     400     100�<�H��J��ϲfO�&���I ��u�l**�D"�O���ѿ�ο��x��QlR @C~�t�CܶIY�g��u����8�̩(-n�R�ˀAޤ]�f��5ln��S!"�l�X7�T�4v�� ?���=�&�������!�ݖ��Τu���гZ�삢b�� =�����sG�����A��"�&�)��\�q����/���l~l�%:����SD4&c�Lu�T�։����/h�]D����$�P*(�SXlxVHYEB     400     110?M��w0�_s̐�dk᯶�i��u����2��*|�.n��.JZ΂�[Ijͮs�7�N���T��[�3���VSgӛ��#��l��Fvj#Θ�|�Z������ߐov���w��܅�f9���6�j�+k��>��KO�8b�W-��2�Җ�H��{���ݬ># �l<�d���1F�)ı��[nv�T�{5���g&h�4����R�&�����5�m);U�����iq��l� ՘$�aﮱ��sc��|?+�WXlxVHYEB     400     1101¾�S�+;J�>�`��UE��7�Ǩ�#��'�!�@�:B�<��d����V.8}��(��	"tK[i��8�/@;f�.�$kH��\=���أKl���nC1�ȝ'���F-����?�7Cޏ����-@��P���� O�{��c:匿L���!5���,�
�R��s$��3���UʇR��!=6���%tA� �AM�j�#���WYv�Q�#��ܠ�:��B$�وO��湢�^���Ra�Rp8��ߢ���
�C������XlxVHYEB     400     130��g����\��%
ò��(�QB@"S~�g����qoT}qPt�iK��qP�>� IY��k����3�ӡ�Cw��>��,WP{h�dB�Z�?��6��7��M��}���mPf�Q�D�yK�D{P69e�N���_���d#e�2z&	�Rr�J0O0���Z���|1�-�/�`�$B��I]�TƇS����t)�ʙV�|qN���ul)�t_�=��j�e��ơ�|����A�$4t�Z�&V�j0�xJ�;0��>J�Ŕ��h\h�BZsfT�n�|}�"�]q�]���8xyܓ��-��cXlxVHYEB     400     100@�Fk�E���F�*���|\<V��_�2�6cE�1+��	��v���pi���,��-��?�T�1����)Zi�M{��[�/�L�)�9�i�]��W~<��˖tE�c)���5N��hx��Ԩy����`��&3m��RJ�p8S@��{\�&σ�8ly�U��_a���?���v�L���-�E��8���
 �}|w���\�O��ZˮV�b� �}�W��!�n�ټf��Y���)�~*$XlxVHYEB     400     100~=���7^V\4zȃ�4w�:p�mfm����|ؖ�@%' -���M[􋡂˂���r@��aQ=aPJ�L8qS��|6R���/���կ�[�o~gY8m�ޜ0�H��7�+j&�mu�]�{gF^���&D$��+^ݣ��} �go2�������+R�X�u/|@�^Ń�u#E�v�ϗ 1,�^���i�M�]�1��-�	���i��Jqm%�W�����b �=��
Ҏ�����p.P�l������XlxVHYEB     400     100�X_dU����Q3�n�F%���qQ>o(TT�'䇜Zڤ��ׁ�9�8�j��R:'%F�7�=xso�#la�{�sN�XPz��1Ő��jQ���L���_&��o$Xޅܪ�(���w�@�"7	��Jɔ�w|�t>�M�T�����v"�%g6M�>w��#`�\嗮��1�-��mż9�D$O�ϖxV�?1fC?��w<�|�M�&ʂӗ�sg�i(��Eh�L��|<��H��g�)���w�iXlxVHYEB     400     100���pA��8��F ��Z�%u�I�F61�PtK�+�׆./u���}y��L Eȑ���ά~0�`:����fX�����|�C�fڒ���@���eLxKt-�Γ�ːr�L�_Ҁ�K�C��G��f�,#5@'�1!�>��ەW���]ݶ���<�9Vҽ�A�Μ�����wZ���i����=��`�SJI�kS1�b��s��_�8�+�e�1E���@w�Y���}�s�=�ԣ$fB��XlxVHYEB     400     100��e𰰫���Kr�	�G����-؀�|�A&f��x�L�~؜C�؂p�T���C��|�I�e? <>��-`�o�M�j��?��a�/!��$*��7�^��9
g+T�?�8�V��;�^2:v	�t�|mG%k7)��s�����J��W|�����7�!�Wv9}���(�;�%Q�E���)ʘ�px�ь����YvPC�\��:�}�b]N����Lő�k�f�}�P��H|����5BpȞ�U�u��16�F�EXlxVHYEB     400     100�F������Bt�a'tyy��[J����Gk��9�K=��;K=��nɜF>	������Ya�v�a�l,����r!G�ge�$� �Xe2/\�(���Y�����F(�R��9�u�9T(���B��n�}]�e�1EbbCƁ�(ٓY�в��=w�5n;f}�H6�\G��bO
ef���{���ǣjl������pX���N����q��1������Fn�`įI��Y�Y����B�A�J��uXlxVHYEB     400     100g%���cY@�o%�|+�*��O���-͹��C�Z�<:$;��;J�֢�ͦ�u�����^�������02_B|���I-���~�Z˙���|��Ea�>����R7��j|p^ß���>�I�<�g����4qutz\H��Din^���%��E��[������n��%�>���Ֆ~�v��F�f�[Q�͗	�"hE�RUJ�"��'�����h��ʳ!��􍚪�v5s��v]X>?>5�XlxVHYEB     400     100@t�ӝS=EJ�.2���u�oظ�4�г6�͕ w���D���|Z®#5q�h��".�~2�7*�#pKy�ɹ�e�Q!e]���o����`����@��#J�%L��{��M5X\��\�(�����x�� 7��s�4�j�4�F�÷���.$#.�����D��i{z��T{�OV���h�:K�")LdR-���Q�H�f�`u��W��6�$� ���	�|sԾ*���B�A�8�=|s�U�<\α!�^��XlxVHYEB     400     100.!���et�	0(��/qYʾ��Ug�҉�a]�b���� T�HP��e~g�[�~l�Sh�~ճ�Ui�$�=�Q��{b�O��W=�5��
��x�ޤs�	iZ�xZ���0�L�ow�%+��a��3k�<�wGB^�e�ʤv�͚{,=�5Í�*w���"�)x�N�FN�Z��*T{��d�Y��������y��$�`�<�1����e��r��";���v�$���:��A�H�u�9� <�U1XlxVHYEB     400     100�71�ǸY�����y�&C�>��RZ��nw�_w��Ofbi/*Z�_i�؍�g��g5s��	�FI_�F�{�� �� ^�mN�0��1��$@)8�8�/��bb�z�j��)Ð��7D,�~:��J��h������ꃕ3�a�k�}v�;�G��FS�\���auv�1r�#ک�Jd����9��-k�ձg�eM��}�)ﳮ}���h��N��ܚ���3���oQ�i\*ׅ�XlxVHYEB     400     100��#�n�]�jϧ�[�Jv�p)�����S�zN1�Z��L󟺃�c�ġ�.�G�-=ʠ�|��XC��'z|�s\�v�J|o_T�ow��
 <��r�ǡ�	���Ue/� b�߉bR}I� ��k���VR�:��/6D�e�7k���%�6��]�+�A� :��_Beڼ���|	�;]!��:���HW� tȌ%�T�� �D��5�����cy�|!\�Ns<!��@��#f��j�W�;�wЧvB��s�(XlxVHYEB     400     100��|]�[��e0��ZL�u4s�g(�ƺN�}�?W��v�s��$���6Eh�PѦ�*ѹ�}�38^�Y�>Ҕ���E�n'q�Yq��,%ji/d�1�+��,ܶm��n��J���d��e�ؙ�lH����t��":��S�=��tH�~�V��x���:��J�A�9���Z�amυ�'�0�������3�%�|�$�~�!c�P5N{����Q��tRa(#s�<�
�M���`����J�Uꡩ�̸�XlxVHYEB     400     100��}�z�d�z3��'Ax��Ŧ�������� ݜ�	���o��)_�HwG���PA	���-���t�.j��b��և��[}�+	��1����6 �5���@���\JZ_�i:��sHu�m�{N��b��M,���Q���+��&�1��Y���ޱ�c��㖊�FmA�D�2&�����Ԣ�/8���pdEA����o�_�o��9��g����a+�x�0E� ���"�ۻ/�M#`���&�hTXlxVHYEB     400     100�*��G���ɹDe�7^��Q�Q\"M	�Iʶ/K$���,�L����Ef�))$H&�d8�	���$�����v����)#d���D7����S��"%�yc�&UQ�ވ�A�\hyl�O�A�=pߪ� ��K��[z� �z����,�U�^���a^��,���z�:O��:@8Fj��6�fĲ�A]jO&�A��)�'�"lB�8���5Ⴒz��r��0ijD:�=p;臻�M�i-�TXlxVHYEB     400     100r��:���:��ٝ {P�.��{)�ffX!��
�ߌJr#�&��C���o�d���B/P�1�S������˜`��������+����$�� w+k�g�l]3P�Il+��mT��:�0�ւqe�L�HUwkQ�ྤs����};�e<K����SA�Gh�7Ə�(�����
�Ө�W�|���
�g��{��e���I��Y�H��c�lx%��;�4�u�Q�l��3$����61�������^tw
�EXlxVHYEB     400     170�ٓK!m:�vQ�~H��铭�e�5���xX�F�����Ҡ�?tl7'4�	\�].)�M����I�觬���|l:�}w����>������Α}��,�9�R�v��1)�4���!��˃��ģLÇa1�+7R��W�V�cpFɖ����)F*��X�$�o=���;O?�r�5?�oF�g?2�H`�AR����L	����y�S5�H�Ci���2����44D��6�3D�?SbyC�	�f�u�9��@m��'���Y�
�`�\u_x�V��ٗ��%>g�-��Y8p�Ϥ(��F��=5��1�0���[ѰS�E��cT١l�A�fu0d��䜚YVM�b7��F����S0-�w�Xc�XlxVHYEB     400     100W
(����k�l��@�nӍ�x��pN���s@2?�7�o��� G��DTHPr!��_ي��R�"��׹Y6��]EiT�b )�x&U�hѝ���������5<Lx�|&�6䫋2SXs_����Y�R�v�}b�7�+"b�gU� fǪ�a��Y+�Fg���WB��"Tdt�G�>�1?1�o�p�{��Vա��v�^���7�N���b��1�J�D�%ւ9-Q�H0�ŕ�d��3�i�ӳ�����wXlxVHYEB     400      c0�Q�]An����K�8�%K���س��~=�43��!�c9��E[��J�	�&�cZ�	0Faw��ԫ"�e�!�RG�u�X��������Y�Y��u�콚��qҲ;��Z�
>Z�L
��K���L�\�a݂�� �t�^%��@�ui�9uV��Z*��ǳ�wn��3z�Q�z��th4�,x=|xvXlxVHYEB     400      b0o�[�Ë�ur>����2��Z�l�]6g�~N%?	uH��%���t�`�����!���X�d��M������n�M��u�q���6��8�(�9�
.�%��#�����*�gU�q��#�v�����^D��7��펟�R��^��|;�X�I
���<wR�*��&�b>sXlxVHYEB     400      90�l�sk�@���e�)F�<Z����b��˥`n�~�֤��w�rU߾ly���N��d��a���'x)9��������<T��I��j�@uga��A^���TўA�mj��t_�������d��3[R��c�M3y}&XlxVHYEB     400      90�TX��ß�SW��e�?�?o�����<�" �E�UT���]3tMa�cj.Z�Maw�=ʼ0g����Q'8�"ف�>����8]�ʱf����L�����{�(=�Tz�I�MsV��!�	UB��솷[�D���I� �XlxVHYEB     400      90ďD�a���\ׅ�4��űH@�ļt�X�l���V���3�H�0����M�S�l	W2")�o�`�I������c��@h�%�#
�q9F��=��֢,x.K�gK9� e��:&oF� �_q*��˒Y�+��8���ú����$ss�XlxVHYEB     400      90PX�*bNk\FKsm�%$��{����ι�v��3���Ʋ��RP���l4��V�˝k��5Az�E(&���f�k	�᭎��v��?!�J��hy]"��Y� -��v�w�75�NZʀ�:N�Ħ�I	}��?��L�d�uKF֒XlxVHYEB     400      90���^��g���/1U|�����.�`�͢�n[��? ����7�3��z`/ty�mϻ�	�#ux�ZoA�dB Ok{�o��GP����6�Q߉~�Q�s��z�>����B�y% 4����u��uP�<m�\I1��4Y���C�_XlxVHYEB     400      d0��g��1 x��p�4+��~v֫�}���eqp�N�E�~����f�/��P�/#�)#�� �|s?�}�)؍�w�^(�=NL�`�*0P�DQ�;���%�	Od+?3�}�6�]��SF*���-	G��!@�Y}��"s��D�Z�O��tW�`�;Y��NrIV���3�%��p�8��(�����Š�j������XlxVHYEB     400      e0%�=�Q��.d9 ���9ƫ�y.���:�q��<��D�͝W�8t|�ht��"��n �|;��E����]Z��)�|�m��}]PC���n/���r�
�%�l���L,n�8���YO��JϷ� \�il(^?��x�T�eB$I���Pc��9U#bB��|�C�}����+�k��3�%���i���W;%I	c����U_��yf�i�j	���	���~c�Xw}�XlxVHYEB     400     1004CĢ�U��k|��X3o:A�i� ޚ���SC���Ɠ:�!��7<8t%Y��~��
���Hn�%�5WDwa��ݕ�*4�ʕӟQ�o�Lmfj<-F6�N
_a'�g��;p��eC�(�X���2Qf֗:�+s�x�|4�&������ڮ�Fs�m�S@ [���9jh˩X��F�g�՝Z�w���!�������Ը{��4	Aj�
*��=���/�β)�_�L#+R�gǪ���|�#]G��%�3��XlxVHYEB     400     160�E�@M4X�1�*��ٶ��$V�a2�9�BєI�8���Bt��_�C@^虶�(��^�6�ڊ�F\!@B;�ŀ`NO�m�?�hA����/�Q�e�Kԍ �_MI6	����	�"��>;Ʒ/?��M�٬ɧ@KY�����AԚ�iQe^U�3�o��(����ft- ���{4ݙ���~!��Gp�����<����4�P^)���[>'V�A��K+�����G��[=92�������[�C�f߽b������ݘ+��$p�c�Z\�L*o�O���2�l;���@�ᇉ���G����}�6Rϡ��k�O �c�� ���rt(��'cI~Jթa-<�|ZTHXlxVHYEB     400     160������ʴT%����N2�:'�M+sY�����b`������}K㌜NnUlHSA�$��+��0��ð�&���'>k��|�B�і��-|��]���v��޹U��~�Ao��
a����'�+�z���K�T`��L�~�Y�h������+9L���Ml{ytc�~��>yK��CGm�O�!<:/q�C�b�E��3���f�b(�	�����E@El�P蛹d��|L��Q����x�u��c�i��~�8~�k9D'z!I�?��z��Ln��&�kV ڕ'~��F��,v;��.Tį9�l�$6L_�5��m$mq?mi���
�Y���tV���؍p.aXlxVHYEB     400     140��o~x��w�����vp��!���^B8f:n.���x�D�e���ϺO��:@h��E}���5q�^�{�}�c9J��US��2�!�8�5���ԉn�����Q��u]���1�����-`X�g�8^F_e3cwC%4�_.��?�+(��������H��
�iu��l��WԞ�SNÛ"�r�IY0y����%��P�i��ΐ����yw(�m����Z���.�w������T;����c�eO;�B��v�D��T~#Ͷ�'�mIMP+��@�f�`�N�X�'�)��m��~��m���{��:�$��XlxVHYEB     400     170X>۱sʡ�v��=�d�SU��T+���1���j�C��b<Q\���]>T�#[���l�Jo���ސ06qK�7F`ҁWr:�x�Q�\O՝�����:XoO�k?�"�@�eG�NFsdM�e0��*�NՀ<������_�3��H�GX�G~)�Gw� �XnQ��8�47WK&I�V�U	i�(��j��x=un4��6Fp�
�����V�/W���:U����K �cr�2%��y�]*��G)�����Xu�`f�ȼ��\�	�;Fi��d��Ӿ�Y�S�*Q���g���V��{��B�m����QD�|6"De�m>>��v�Sa_�I�bۂ�1f��R��˄���4ǐ7(��i�XlxVHYEB     400     1508�J��-���co������ו���q܏T
X�����M=+,��\��=L
��'��9e=;'!���}�Y�Ix�P�<�j`��jwz���GR����@�O�ԉ*�6��sE^��W����#⺚����!-����N�)�8L
8�_�(��K$xBŒ��>�<vb�LH#��c���DO9:�������%;U!�������P�����A�ʇ|�G��JASk�*���_:��JYY?ueO�hwXٟ�s�KO .��Ȟ㩵E�cT�w�j�X��+̙fݷCӗ/Mz�;��T?Q�2(1��w�t��ּ/�X�N�[XlxVHYEB     400     190ب5��#_�_n:�����.HB?�>���W;���ޮ��Qʘ��
��uTO�|�`�|�tG���n�j2�b�T�b��:�:�%�T�}U'��������kʰ�T�	E�����U���j����"~�vU�Nt��
��YI�U{��.������}�k�
��KyZ��Ηn���3�7�d�I���Jyė��,��IiI�֓�|5�]Ϫ%�����U+��&.:��v���,|]'N�y���:�E���l>� ��p}�({���+� �7%��EC��gP��uFǮ��n(�  �O_9|M=}��I�z�IyR�x�R��]_xW��e��]�^�Q͂U�t���X�#�9̻��AN�<^�.�������C�n���D�B�\���7?��S��e)����9�XlxVHYEB     400     150���H���V �Bs�k@g�Q��7 ��Q��C�p���4���a~n�#��(�̾��6�&4� I	Y���+���m�l��HW���V�$�����S�Kd�ó��*�Q>">��DFk'4��h��e��0k��ĳ�]��8�&=XTе�`l��V<?��@��!ր����U���Y���=G����wk7����)�-��L���)ir���
"$�DI���(�E~�4�0XE��a�1���f+�>~���߅=�/s��T�#e�JQ٢&+�-���	�Z>�Wl)6�L7U
��x��Y�]��yr��� ����Ω˕�d�XlxVHYEB     400     100�*��O9T�@mÑ)x=e��#<.'MU��*I��^G����(�&m�Ο�����'-$�h����Y�6�o�k��}l��ٿH.5��3J��G]�z�\��j�F��7����	�Jgk�?����[���`|r5�������������3>�[�I>�N4��a@�UN�!�M(no�
�f�0��҉�����������6��H4S����
����!]���;wF��o1_�'F����de�A0k�x��0�XlxVHYEB     400     190z�2�W��f}]�] y���e����k�n�,�o�/[�P5�n�m�vl�˓v�����1��o'���|	 ����S�G޷��c����z��0�����E���n�I���C�N1!�%ǽ�����؂~i}҃Tƻ@�M�V����>�,��R����jP�dTJd�ms��x�����7��<���y��z��{����k$������h(���[ltXᜟq������C`@̥Q���:���0�ء�} � ��=��n����S����i@��C���{�����_w�c�%�
���'M�M$���jμ����wK�L3*x� n��[j�4���!��RS�;���t+��eӾr�� �on����_̋���FY�-gK8XlxVHYEB     400     140ŕC?.$����n��-��1�Gp
iM��N�SbKR�X]n.�������t�ő��'׵e4����=�hqQB�����²r2z�q�3!�wr���G�Y38�f��@��;]�7Z�`��ӌ7������'.����_��s�#�4v��������ޤw�Y����*�G3:!KWY�x���%��������2����U�����q���;"X[��*���%>�sm�2�ҏ�Չ9�Fi�(���:Bam�W�:�QU> �ֹ���/�O����x^��C��[�e�u�{�9ʏ�	���N��Q��V�9�8��+�QXlxVHYEB     400     150�%���y�m ��}�r� �!`��{9f!��;i5\D��1(�`L/"1[s��XP4lN	1=˅UQ�'h���}V��S��J_c�sz���r�k�=�ALW�*('�r�Q}+�J?u���H�~.p�3e��r��l������)O>�����+ks���]�.�	\��	�c���Oy
|߁;C��1"��Ҫ\�Z��5@G�w�{�PݍY~��=A�M6MiQ��Ğ�9?c2���uQ�tE�|����O6V�ڧ������/=ք2��҃�5�uu�Ni@� ¡�#�� ����C�G?�_��n}y`I=�#�c�����p��1x/I��(XlxVHYEB     400     110�����u'*��:Ϣ�t`�}`�솵,����$�!�yf�Q�C_��q�u$�/ݺC�dP1~�����U	4�{YBd��zD)�^�w�+'�6�{m� ����b��6��h���̄4���w���d���08��>��k���#q�����P����-�'}�(��0�'����+$ �� I{��u�È�;Q�Q���e�hm2�B�C���E���٬�/�e��qU�~Ý�{~���;�6����Þj��Q�pXlxVHYEB     400     160@Sٮ�J��Vmrt%�����LWԇ��07"�7�f�;Ԥ�S͵�ي0��j�L�L����ty@�~��v�
���V]�:&�M8��ya����^��s&?�Ҡ���?@��]�:����h���㴄D��x�>���-�INqĆ�]����i�&���lX��cv�¼��d��!	���?�� �a��ܫ�'fՕk9o����(�N�e���M��7��D�?~�x�����+&k�\�xm �쏗�i���Kˑ+�C#��� 7>|;�rH����;Z��$q�2�\p�F��9,(���{����2��|� ��M%������M���A}�;߫ő���XlxVHYEB     400     160�g�uZ�y�BM��^�gvV�b��b4H���V�A��H1���M\`�_�:��
f$��C(��;a�i��� ��|l3�܉��s䳥o�e3���Y�٪��2�'��0���Y�78�.��'�;,�5/j�P09ES��.b?�88�_>C���]A��f�jO����d�Y���H/0�>-�b�RyR�glܮE٫�2�X��6�����ϒ���e�)��0e��&G��������>5��Vη�\�%����В�(3��K(^v��6?�Oȉ�t���#��P�����J3�/Q ��%d�.��|�,�1�>��u|�i��XcH���CmY�I���zXlxVHYEB     400     1504.�铛m�Ϩ�s^T�.?�ؔ{�;BQ�ʺ�"ss	߀���P�N��z����Cs�G��h̺g\�62j�yv��sLwrz�r����Sn����JБ8��R9b<p�m�Ý1�#e]Pb
xZ�T�$�m�ĥ���l��}�=O�G�x��W�ue���<C�)��%��+�)�R�:g��p�Zv(��p��<�¦J�]�Je D�XS�Uv&���wj�i�.S��E_�80��Ejr��?!��p�,R׎����� �N�'&�d�F5��%S��b���{8?x�u�c�x��ǩ�V:�:w�C�����`���O<-�ľ��jx7XlxVHYEB     400     150���*\�6@�G���ss�1���;����u�II���=���\�4
����~CS��酘��;�5�mPu�q���l7�Y�"%�4�$����ab�@M�V��$���Փ��o��K�%p�3,ND�2d�QX���ytE�3�9\�i�����O�����9�	$00=~l��NR�*z>#�,ط;���6��P��YoP��Nr�\�ŉwt��"�����"�^7�"�np�c���pq�j��5�kߌS�[y`^
��ձ8�g�>�L���\3�W����h�J���h��$L��^ӓ�U�ݧ��$⑵�^L�Do ,%XlxVHYEB     400      d0P"B埧�����~K��¼z��$����
JjUOx�ȆLլ���XA�<��I�n<��<^0Y�[��-%�֧�m"$*C��mЦ�(+F
���'z� �3��WH^�"����7�HPm�]6����됈>�;֥��2\A)Ἲ{f��d	/���e�G'B*GW����bn��ǵ1͹�X��-qۦ��$]�=l�̀�XlxVHYEB     400      c0Ha;bJ�|@T~H:���vWVp(��%����
l6�5$W �y7QƓ��4Y�$c���Zɻ)�D��}$Tbb
G�~?������l�b."�&<�ٗB��}����������g�ݧ�8K�冠��W�r��0&�8@"��އ�h���
�G´�e�����c]'���L�:���W�&�-�$#��P�PXlxVHYEB     400      c0g��}o�s�cip�am��j����*=�m��%�����$��2�4'"��W8&�s3n��lX&ݱ���,��� Q�mŘpz�n���V�ă�0W��d+m�
EX�����/�V��4�P�[�F3�U�z����'	�T0f�T��΅z���Q��9 ψ.�M��V�V0��i�N���FzXlxVHYEB     400      c0v]my�CO�(�a'w�1�;��|���Q���x�r����.q�2��3'��I (#3T�I5��ʏ*C�D��UՒ.(��t�-@�I�;�-�q�G3m�%y��L:�����r��%�z=l{�u��O4,P��v+���> ����M]��,o�!gX�j�������6�Ô�E�<�$@����|�$��XlxVHYEB     400     100M�|�%��f�K�h��pC�u�.<r��W����r�?�6�5���+<�^�����򾅸�~�Mtx�>���W��K�\�x�9����uB��lW�KBiE�`�s/=	y�#}LǶ�^���Y�6�\������miUp��T7Z�p�L�g�-����يu�\`��Y��ꥦKU��jd5�{1�P�,#8�z���d�Slƀ���2�d`@\^��w���'zYB,Q���k��]�;��R�"9�XlxVHYEB     400      f0ɳ����7��	s#��2D�KR/�Z@N�����-�n���L]�%.?K+����n�AU��Yhgw��p$#a��
yrKZ2���C��!>�@ⶍ��^u_]�I�a�����'�4�ӽ��_g&Hkb���E�x	�:O(ք>�j��ʀ�_����<���^�9���v�I ��O�f��R��{Tݕ� 0]�����H)<�� l\$�$  t�(������8�~�����2��XlxVHYEB     400      f0��qb�@ĸx��Ǭ�U�?��>̺|m`��s�`X���'�
�`�u˃�5��]�"Kx#-��t�:��&	�2 U����C8 ���M�㒪�������Z�xl��@��Uƚ_�8�t�~��!���Y���"@V�<Z��e�����p�6,$��i��GVƔ�\���H�?��,9������(��0�Vwk��]��Vc���g�������2�r1[�h�Ez���b��HeXlxVHYEB     400      f0^\��զ�CuLsqݿ�?-W[sɋ:H�]Z:��慛� �k^~���Y��{|�\���L�JA��x��c�,�����խ)���z��BT�6�o	��x�Hzڔ�v ōV�Y�і
��᭲�@=���������M�aۨ�lâr��Y�5nV�_�Gb��U5�P�\���j"g.b�u���z'6�n	M=W����0p$G������L�E7�\_��ͨ
�,�s&~XlxVHYEB     400      f0��^�����p���Y�@��HҴ`��o�]I���@&���a����I�27�����I��p���`����O_�5�����I�7��_0s	9  ��럟�L�����#fT�#�0��)m��8m�n$2��o��=c�إ}o�?Ɨ���L])�B��m_��sQZӆ�P#�i�:���[Ĩ�[�&��ʃ��Y��	��NT�����	�s\m�[	�}��Z, �����@�c��XlxVHYEB     400      f0X��!���b#*�,,X�+E0��}�'׫
+������栿[֨�z���j��[߬��Z|��s{��~�'Fi+��VZ3�}�0b��7�is��,Dz�fW���9?q
�(�}�{��ݧR D��#�b0������!��$�d�X�T戹���e.�� 6�(d��(�?����cƥT��h0��Pl�赩�C��1w^DY�n4�2e��:���3�m�z�@E�XlxVHYEB     400      e0;��
�g
�������;���i�M�9	�Sm��g-;�mK;������mr�{�68H��o����kD5*?�y�+�}���mZp��	�	�+�'�Z���)�R�s��tc3��	�ރiu��<<&\z�a�Mu�< �@�},$�`>��%����@�����X2���*I�ED�OՓ)Y:	�ĸ�v�[�p������_�3Q Жm:|��+�)���mXlxVHYEB     400      f0����Z����O��r��b�o_�+���I�c��7�E���E5�\�\�_��1�I��d��a�P�h��_Խ�L�I
�p!��*Z���u�f,�_�~�ڵ��3RD������G[��3�3^Q#d�������}AxN{k����DP��}�8�us��w�6ǡ.?�{��&\8��g�"��ZZʵ�C�Z�b8���>�v�P>�y�	C��.�Mx+�$<�����������vz���%�XlxVHYEB     400     150S/&���ڄ]ަjHn[�hkfos�	v��;�i���E����1K��%r|�Wdvl��#:�t��){�BxSeT3�ɭ��azn����~݊~��-�T:��)GV2��F��LdGL;񟓙�s9ڙ�(|��ۑ��Y��3�O�o4v��!fs?����(����k�3�����.�ME���sa����6�|&[� �#N��Y�fGx8�},e�̫�NMNyN�V�4_W��v6*��Pq�^�"�b>#T�z����w3�FS��U��/��������5��=xgTRX�AL)���5��X�l����Q�{%Zp��+�zIga��XlxVHYEB     400     1a0�g$���V�|;����Ƣ�=/ub���k��a��KP=u	�YaZm6	��@�|�6�o�=�R>-Q��M�{'d�3B�/��Ĉ�z�G^��bΟ�v��9���N�pe�YTG���C6�Q����~ڛ!&O�����|�G���~�
&���s��n���1OSnأE��"Q�h3^@k@Y|]���������I�E�x��# (��f�D k��P�Y�}R�V�B���Ƌ��hR^~C� :���T�m�Ad�ZG��>Ҵ���}Y��K�t;�X<�IC��oR$��+�Jk�4�����%�E����< �� "$,Z���� �NAISx#5ɗ��h�2* I�f5r",e�F�N��k���:�ѹ�����J��d�OQ�k��hd��6ۇ򟱧S͞XlxVHYEB     400     150�M�	 �c�۷�,c���(�"��D����3��L����@�f�f]s��?�r�͕���ܲoSY��:�R=�=�R���-�6|Y57���O�+�=We�3�S�m$�p��[�Ԩe��}���B�}����"��`�PPS!r+p_�����j�H���òd r_qC�gS@ȁy٨�d����HA��k(�2��C��b����_��^��f�A�T3h�\S*�]��A��VS�z�
$ҨPRx}M䃚NM���Y���;�M\�$�8���Y
9��.�O��F���u��z7��Ѓmo�eج�� |b�X�ָu:�@{d��XlxVHYEB     227      f0����F���sV:�b��d�;�qtw��H��q�ݲT_�)����� ��}`���E��4�%Ω�75ULaRܔy�4#��׎����d�"]��͟�yT@I�F��Ԓ�O9UM:��dkָ4�3\}�����iM\�&�a��1�4&^���<1�A����q�G�
��C�Cҫ�\)*x
/5�N�;��W��1�����h��^'�H۲�W���,��z����