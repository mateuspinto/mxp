��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���o�*��]�1�Z=����y���<��(�����R���D���qcUT�'桴*�xO��nck��+���/Y뷇�Ė���
:p�=��7��Iw�|��9r��G��i@�A26~kǻJ_�/�iĬ� ��Y~ *��jN���Kdp�[�<G{�Ml�zn,�춣���u�[��kbJ�^�\]{3�6U�qq�g�|b�5�+��yc��@��T��U��h�Ϟ(r�@B"|�Pn�7u��>������&�U~d�w2f+$��=���y2��g���A�v�����n�B����w�vҦ!����[�bc�&[!6�̮�f�"=�ZdoZk� b�����n�3�jC�]i�z���ש��)A�>
��e/��@���ȿO���.�4V�^��ͼ�<�#L�S���奜��@�le�~��nr�S�&���oK����B������s��[(<�U��ֈ$��M��d���1;5:i�_:\H�A��^�����.�Z^����7�cT}���(sR���uRF���n�r_)EL���B�����ݛl�c�[N�?�=�;I}�5�@��*�rB�(W�s�YA��9��ө}��LC��<�J�+�ƾ�}N�2(���;Fv�����߾K6^(��n)<|����ôŠ���u[���ez���i
�Z��1�t�F�l��N��7�Ir�
μ�:`!F�_�`������17�����_�����s�������7i
�v�D#�Q$��ẵB1x%�o2m�`���_����,� �d�JՍ��i[\�'�#��Z�s��X:�ί6�;/�WO��CRLQ:L�<V���dK�G��?^Ů2���J�6V�%yg�ݪ;�0�������s��h7[�,5C�yެ+�Z9��{��A����-��G��u�*Jg`����coV�Y����u��tLd��g����S�D�h��B��f�{��cwY@ACh�᫣�g�񂼫��F��r�鹠��vN���Rip��(�x��3�J��D�ߺ_����H�N�2�h:'S߭�+:�g�y�;��Ę�t�C�)_=����><�غ9����'�I}<<�8��S5L��[q͐�^�lH�(3(���q�7��&�\��)�KGQ���*��򤃧%l|�B���H���$��v���اgnu?)9����A��sUZ[�!A�f?�I�b��j�{�U<VzF4?H��Y�ep󝎓�h~cᔺ�Æ��M���ZBO��d��W*{������F'��_ �N�Fmh[��CК�r�A,��+��U��ǧ���������Ǘ�r,�-������j��x��^p�v�v����2'E���oq$�h6���&��S�Hⷿ�v�U�.U}�n2rT�UXq��̨E�|n�t��$�����f��<��3|R���Ƴ��L�����p��������,x�S�ymf�����0��E]�O�� �l�����C�����<[h��\�8A_��_�J#�ᱭu�~I� ��������x�}�����~����x��З�,Ѵ4��
���O
���	!*8�j,V�F�q�-�U�Y��}��>+�4�#췻&Dm��������_ �f�umҌK����SN� 4��:��Nu��xA!�;A���i��P��?�U��Hݝ@�E��f����?��5?�[��!�����a��Zg���z���dg�� i>�Ұpm�ϴ�� �1�����i5H�=� B` %�q�Q*&��6v�$�뙮EaoL?`�Y��i��9G���mF�ژ����F�����6��Y�?�}�����Qa�]�-�B����k��x'����FV��Sx�8��4��?S?�'#�{����#�J��R��S���SX�@��4C?-'�	YW�f�>�n�tu���'�=hP!W�aiʛ�pL�8^��|�:Aڱ3>��ۄ$��䅓�۲�Z�UN���4�+�H�kD�	��6$��l�LQ-���Jt$w�q_h���%9_G-:�i�UW-��Uxy���xz�bњ4���� �G}�)����Q�;��$alx�C3棧����:�6Ac�W�����Iz�p�?�D5k�W�X���# [�� ����U-�i��9�d��Đq��2썍;t�	�����]�C���%�G�I¢W|���Y��ۻT�&:-��Z�e3�_������89� �b�Y�"�|�Җ�7A8Z��g�Z����&Y���Jм���d�4�J,|^SF�T�0��L:��ZU�82�7:�O��ir�ܧ���0]x��ㄅT�:�|M��%S��y���ܚƖ����uT��~f��;Z~��ǾM}�=��������k�Kq����sKXHz�1���o#�B
@ �OVn����G���e��R�py�I��9�.��j6�f��L�%�����H�`��2-�w��l����X�\���5}\><��A�vI܎@�$qѝ���pvW�2٬!�gU�:���̚xw��p
�<��o���}�4cSU��hB�$0/�g������]����� ��,�{��ame(��ī�"�d��D���U�׎d����q�U���Ґu��!xy��S��4�pJ$�Q�T����R��ą{���W�Z��k&t>�)н���b_c&y�!%D��r�Q0P�fC4����F�k�4��b�uhE���/�Kb�x\�t�Y��"ľ�E��d��8�\U�o���W��3W�$pcC$��^�~��<χL�O��Iw�g���U~���P28��<����E���\g^]H�h��W{�ǧ3������z��J�D���k�XL9����!��t�v�9����O�q8FX�^p�<����a��Ǡ��۪���J`��S�/�)����o�[9l��W�p��(�{��%�ޟ*�o{=��.���<ێ�n��$�+E����iK�%�֋L�RC��8g���P��ES�*�ЏT:ٕ<c�t����+z/go~�?Ǌ�c��Y�Q�v�]��a��̈́�řhD�s��h��FY0��n�M���,*2"�׻'��R2y�����y�y��c���࿚8�xs�D��Dأh['��kȹI�Q��Ɇ�x��O(��!�L����o�u�9W�yi�k�H�����Yp�y����^0C�V��t��'5���RX]f��O����Bȴ����j���J���C�Js�x��1Bk�H���Z��[��-��v����)B�/Y���8��wdN1��ru�T���M�pw�(���lɝv{������0D�[��