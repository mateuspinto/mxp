XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��g�e�c�`�'���˓f|���2i���L{�B��Y�ۉ���Ss)����#�?�s��Y��vU�	k��חFKW������ٯ}�cx!�����'��GUo���͕ͽ���R��c m��>gܒ|/���F���\������F��
�_�SW������3�#�$�r�ܔ�噯I��A���~�vu�Ui�r��#Ӎm}g�9���m����l�����=fw �%��Q�K�����-%*����h/Y=�|��`�ϟQuZ�ێ?�y�?�R3u�����ۭ�]'k�<ϖQ�B���І�%M����NLt�z���&VY����{D �f#�+� ӿ�4����ὓ�;Z0{�	���F�%����з��^x�x��zQ�5��ִ|�ɴ4��ŬPN��D2���Ư­{2��Mby��3`����Q�~=;��0>��<�sK�L�)(���|�&n�]���X�֚�x����2!�W�'_��\�̞�c���P� ֠�}���8�W�ݕi�x���ȂcOf��ٔ
��+����D/?�ﮕ���{�d��ڹ��ܚ��M&~�èE�6��!��a�^k�m�� �<f��R��F�� �P.���+x� ����ι�-ǹ��l��2�KS�J �v
�m��3�c \�6��O�����cT`�j������=�5lz�e�����a.Z0?��\�?ہV��R�G� O��<o�WIossQ/��,�F�M.�ZvVBu�6-��}��/0XlxVHYEB     400     1e0�f����L`*�lX��0N�3��4)5r���K�p�kp�0�.(�r��=M�'����,g��C���,q��Z��E�b�w��V�"@��FL+z��N����2W������^v��&��jHg�Na+q�x���v��;�_H���J�WKa:�Ȑ���A�&�z�\%O�⁰p����Ʀ,,�d��N����7��9B�7>	���R�]�:���c\TQw��o�[*m��&����;����h�Z<3��O*��=5��g �V蠫h4�@6<�L͒�T0���;S|}���hFA���!��a %�me��w,LÉ���U�����O�"e=�0�v˫�h]|qX�a&���b�u�7�:7_�e��7��}�CL̄�(�s[DF�;%P`7�t� ���E����g�_<�^+9���V�~����3zf疨��?�L� f�l�+�[4c�XlxVHYEB     400     140L����r1E�\^�K�xvv�6�[�9�v\G[2Ŋ0�1����z�֑�O��}e�\��m�^�5�zI���D#��v�xt�в���L�c���?�Sh�U�܉&�N��z��ȯ>)�CYO�_$�mG�D4��c:ѵڿk��;�I<����ݭ~!t�!�����[2����U�Qb�HF�epJ=�<�e�v^�WM���b�7����J^0��֒�2�3w�Py���Ǥ3��RA�Ŵ1!���x�~�<�~�]����˳�]��~)��54�3�.=�̜d��[�G�� ��/MA 0�2p�M�I5�4���XlxVHYEB     400     140I�K;�@"��6[0���콢���4�=��?��0��V
L��1d#IFبL ����U���)�~Z��RʀQ�԰h �i�>�`�&R�I��̵�}�JK� ����8�{H�bKfR��y��X_�R���Z���-�����7�]���)�ό�*~���#��Rm���D��L���$W�^�1��[��ke��?L���-ϟ�-�)�^��81D�S-60�=v�r�@0 ���>5I��ט�+�z�" �m������i���v�����=�׶��*d�
f�nZV]���G������)�q$(��L̓��>)n)��VA�XlxVHYEB     400     1a0ۍ.⫭e� MbU^Hm����"���_���0�3�r��@$�.��2�[D�M!�h���F��u)9��^�,¶���u^�Ι���v�h��J59�F�K[lj0?�by�4��r��v�b}��Rqd.X���!1WV~p�T��@�[�D(a��� �ԋk�.�t�'k��r��-~�t�<R��/��;X������[��d��g�e�5({����j*��H�����Z��q���AM@ƥʢ;�����q���h6�wk��|<�,X�37�%�	����2�{�Ĝ\e��ge*s!�bK�حL��n���{���4���;��T�ϲB�*�i��������Q���f�����r+��ǽ3c����S
`!�@<����u�� ��'�^Dk��lZi#ٟXlxVHYEB     400     130A�l�B?���K����Y����HF��"�6��nf����f�I�����RA[8���ei��Q�����H��E_q��wy�^3���Q_�G���M53��5�����/��Fl(L�Dn�M�F93ہ�>U�0z�}�bl���&F�b	�|��X���{q�JD�3�(
.y^���49v�{�:�JL�K��@l�����w��Ja�\z�@9:!^��Y���9�B��*BkH�6
>[��"�BC�3"R�|R�ǐ�{*3Zk�5ʑȢX1I��^�������b���٭ݎ�� PEXlxVHYEB     400     190;�P}��@��	ܠ�^�&��� �1 ���\#�CO�~�<�Sj{������^YP,x2�b�M�\o��E�k�@��L�b&���N��R�i_P�ݞgc�s�2�<$LX�%�Av|%���<G�I��')�)?0�g�w���ە��Zd�?�K�(\���ba�9D�a�K����^	Z��d�:�n��->|�v��o�ט�0cS1պ]�g>�6��B~������u��y��9�L�.!t�U�s�0���k�~O������ L7t�����.��}�h��I(@���%�>gWFLX,��7[��e�����賋U������$�u���={���vF���K�#�$q�[�.��#nM�1x|�G�$\��j&.Z��L4�b6��8�?J����XlxVHYEB     400     160��	�(���{�C[�y2EP�����K��6ʊs`������m|�Z�8ٔ�+��㱴
���@��V�:f�J~��i�͏?�V&S�ĵ�J�;�ꀜs+X�й�		��	鿚:<�Z���4���������A�σ� �b�K�w�T�_�ՊCPc4� �ʴ�Q�n�6���
��a�����+G+�`~�l��U�3�o*B�${i��A���KC�><Y��T^��G��]Q��m�B�V���üw4mZR �q� U���� 8mn�?��1�m��Xl]Uq����'�aY����^^�bx8DRT桘���L��рG�Ù��#<��Q�ȱ��_x�/����r5XlxVHYEB     400     150A�}��o?��H�@���e��>��x3j��"�j�z�x;��� �I��U_M�� ����_�{�-:R̪Y���Ea?�;<�U���Oz�b�a?r'�VA1!	6�ex]MB��jV·���$��>1� 9{6���)��k1;�ra�`�7e�{VF*�H=��|'���Q�
l��p��z�6ڒ�� �*1N�f���qK:Amn��U���V�v���Ȓzu"����zBϨ7j�����'9�-�X��|����[�'���^��Wj�!U�Weei���k���I���q�x� _�c.�!�2�-�2|�0q#ztn�.\ޅY���R�UB�XlxVHYEB     400     1b0��2� ��󔧩���h�ة�2�v�)�[Ӣ��6�i��yE�R�O1BrO��kܵ���еM@>L8���D>�m��RR���LOQ�����	Z���p�WLsA|� ���~��G��š�A���z���+�(ZO	Д����X�b-�@����wϡ!=^�.W'��/uXO$�Q���wL�C��NQ�����y�4�;V�i�߮F��X��ӎ�*�An�{>M�,wգ�Χ� �&&ϊ��?��i{s����ݗ����5�)�`���'"���� �0�D���,��wA!n��ҴP�r�ӮOq�4L	AU�k�p]�_n�a~y����p�=��e�#/�LT���ҋ^3����=�i�rL����Jnj����e��Q	U�9�9�[Y�`)F������ B	����7~�%XlxVHYEB     400     1d0�ٶ?	co�ewM�< �v�q6N��\C����8�ځ|0�\�.��%wA�:s��A�K]V��UjԐ������=^mM��&u�V�CP$�O$�3�k!aIB"<H7Z���RR��Fڀ �z��!Sp����r�<�sH����235j��G��"]$&�)�H��ǋȘ=s���.��%�#<RA�O���`brTe��|3y�gCG;���S�aCTs�;;݃4.~ל��6�b�'ƫh����I��R��ǇkLvh�M؄/Tx2�t'
Ő�K�O��37�h� ]�^�_P2�Q�o1cET���U{S^�o�<C��,�[vW!m�I;���!�i���5�AnX�
�Di���S��b�~��;8�}�jeѭO&�͸D�$����{����>ܽ�/sQ��i��z�G��q{���+oH����10/��-�rd��� X���ٻw�\�ߢgf�Ӧ�~�F�t�^�	�XlxVHYEB     400     160�R�+a�BfHN)�,_�����=�/
,E����a��&p��[�r}J���e1�ɝ"㕰�B�A�qU=$XF[,�(؃\s�x�%S����b�`$��
ѫD̀��a��'j�m�s��d��Q/"g��m��)�&��F&堃�/P �ʦ�ׯ>2f��PQ���b|�t�X��"�]��5��}O}����B�y͡����{i�����X�J/k��h�]��5��\�������Gd�D�a�0�Ήmy2��/9S`��'���A�����KC{��y:�2_Ck�/X��3�7w��(�SFa�����0��D�v'�4͙�2TÉX$�1k�¼;.XlxVHYEB     400     130se�N[�A]��ij�� �S������;~X�:��������)�HDpHr�1��M/�)z:�ET���#2ڣ��>�@.^�rQ[lq0X�>)�����@��KȚ&n��Cz�y�L�&��o�[�I
(�$�߲T��[�๓V�A�	k��x�����\��Q�� �H�f�����$V0H<��~m}��z�3t�%�����۪�dvR�Y�RJW�k�QdJA��C��<Y�}	t��ʯ�=<@F�B*F�@�$axA�TJ
�Z����+�b�c�*�~`�d����LnS�XlxVHYEB     400     180��fs,�IF��6}�)���7��Z�QV
�0q�!�_�aR+Wz�bV �����-(U ��v���-mԝq��uvC�Bo�9� �/��- ܰ>~sx}VQmΚ�ԝ.��t�s�\��>R�5��2�+Q߸�����{+���u6��*MT1E�
+���9MqDc��L�}��9���\�V�[���I'Xf�����5Z/�y�1<�-Qc4sQw�Qߡ�\�0n?i��Y���73����9��/}��W=�G�04e������ON��ۺ&L;����_��m��6���R�Q�T���6�K�g����>HQbf_*)1N�6i�]����a��h��z���Z;ؐ�ķ��R�����8cl9Z�h<�=���ѭXlxVHYEB     400     150X����'�p��A �$�/k���^��)w)x��#���Ղ��v���.LsjVlۡ6�r6fz;6h�F� <�	��(%,Hh��JDyl�tC�󟌋��_°@c�b�*��2���� T�������"
ͅH�L�'��#�F*�88��������
���T)DFL�e��j6�wL�f�B��ʰOwJ�7��n^�0v����糐�ĕy���(K��4(�s��a���7dw�0��V�p��}cكƺӘ:gRU2�Gpc��������+Rh=����xp�l�F�*2w	
�����Q#����4�-XlxVHYEB     400     120�H�!����3��yJ �V���s�88o3}�@��f��ϖY�=�I""�.e�jJ��
?��y"i�˥�����^[+�u���U �"�T �5�%��(2 1��R�X�:6�!��x�,�ߛ���9n$N���G1�yGi����Q8���I�;�h���^���g����w_˓�m�K�5��V��u��z�_w홨�����i��2�kQ�՘��?G/Q��DI����eO��5Ň��ݲ�[ �]g�!#�sN-@�|�Q~,*���4sz2U�XlxVHYEB     400     100F�\�!���e$���O��_����W��u�4N�!b�H:9;��]��@���3T��@��R�����X4�m0;]���펈lx�Ҳz|0�m�ɍ�\d��pZ�f��UIīm�l@��v�e��_n�GGq�����,�p�*b�]�c��tt`$Yb�#�Wm�gU[[	S	ܚ]��E&a��A���Z(L�"�Ymg��ʝ:�[��Gl�G7?T�A��/.Ƚ>�>��)Z�hڵ���XlxVHYEB     400     1a0���
�}~yQ:�=�YF�w˔�d��d� ��*+�{F��ּ�A����H���cEW�G�(˔��AhϦXP�u�������ۥ����['��B�=�L�r�a��4i�]b"'h�ˡ�
UF!��À��#�"b*���	��$�r����u���9��~���1+>�~
���~�֙pH�ȟa��O�m߱��Q��hL���t�֟43}*w.�E4k>e>�*#Tz��**}3/vO���� �K� ���m_u���E�&�k!���M�<����	��&��c���|���G������Y<��쨂�b�/� 0�R١�Q.��Ɵ���2�mM�*ׂ|�y�/o��*W�yc�B��9�$�if̓n��l���E����;��gSh�C�F��`�t������xlF���XlxVHYEB      27      30U/E��(@\��s����^�#s�l��+��16Y�-��x�����