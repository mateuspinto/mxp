`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25184)
`protect data_block
LnMLzjeOA2qpUkbJ/C/BZlFC0pi+fXwYQlydcaSqu1v58LUrBP7M2GdC+gzbLOBJqnczav9d9p+y
1u8rQMDf1ZGMrrlsD0NFQHRx7V1STpa1IXnYa+D+6FVRVjEmrfuQSYjuXipjnioeOOM62yEWsER5
fXFuWzWM31SV1VpThVfxd8Qc2QmmtuzA3qJCKZPMJIlnCHmpZcgX3YfxQkMW9AJwZ4E88VB2NIQw
I89LlNHh22SE6w02sFY8q61B2oJUgjSpCJwIdSEZm7zkgEmcRRD4YgpQcKB4KtLJIBcJeuTyLHZ5
EKcEU0mJRvBtZvblpJ/etqbiQse7R9wfJIyVmdzBMV5uhwKmLJvn+VnpDg3xAOVK6gn2jKL75xu2
tY54nvIyrOWdu24qIYrNT4ex7b0nY3Kjlkh4WpHkLnPt49RvamJ1YmSrC7Lrw2oYOigpMDLrKY0F
0oH/nW2vuxan+LAvXQM6NWYtm/cG76Cjsq1aGw22LYSyVLVayQkNs+iS2KS5P6xO9djBGSmqOAwL
6JCmfDlm0fDwwCUIgrZwcw3ea0NSJfJd8vcY0CaqZj1KuPj7xfqTpKCV0rJcFUZiinQkzN2gZqjd
su3VxvA4TtdReEnEJFVREoUsqZkfhmRZkSJVpj+Q3fp5o1H/0mnGjKXHvwtyEfoXsmH9ysHg9Yd4
Lvupy8QoQUp992JCV8F+MhB5pmwya8PMgU1GcasOv08FouzOYYniYj9xGTXtjTC0IjpL8MVc6k+A
IsqOg9J0w3AERVJnJJMYg7adPMlUXiZ1dY07wXLguLn65QUPtoZ7ap3lz/yFvb7XFsPwgA0vaPFT
VXu7POm8VSzyEHTtOCVkO6MSqiG3h+WmhukCV94Jowd5XL2/ERUcLR44FV50IphzrwECIZGOlGte
hzXpstlp/iDdmfAlp/w+7HVlsmtMxwT5xTj3QTdv2HC5OYVDlMlbJlSjyvEzdn0hP+bmR/aM/e3x
UwwQ6yTBWSbni8tXOmrH8CUzwBQsEBXXF9IE53khTiDXhe2A0UCLFkSrMkR8e07135M/Pto9a6GQ
fSC4IfASYOkElUVwmO6JFaAaXFop5SH+LHQX0qWB/ejauq/hghSObLKqfRYxzr5RXTs2+rMwcj91
IRdcGdlpQM5YRMZuHsjM5W5zo138nbMeI0oAlX3SGjMo5SQoxr3f07fii8VaqtMXVoB5eukmX68O
NCwI9hucBafnh+tFRB0xUIRXcxVp6WQAj5yuR6U/zF32y6KqsM92gAtql9JOQX3rvgIMAhm473cy
mX0hOudTpVfGH0F8pnpRs/X3Kf/mpZj+lZUJQLPhmk6eAngThsXdh9lP1ssKHUqh1CVJpvcSAzfH
m2G5sojXkW0LbqpgzpZftXlU85Q7hp69EjpZJqujU8e1Wnjilt4DMSFwMMhNNU+He66GugRKlB9Y
Q0KPn8g9GLgvvId23tRCwX/w/aqVYZLBllvZOZyCw0x2leCZ3bnirQVTNyO14Jut4QtBj+BaYqh9
Ngxju45mmeRjMCASPLV6gRdCMoWKb2cZarYyt4CNtCjDpwXyX9V9FoRWg1tI0O64jLP3dKAAThaC
47U7z7MGyvn7Q42tnwQho5ahyalv4tHyFhn5JP+VcoeK/a6Hl2g4oyhG2P5kx+epXzJgFH6xzm74
2zJ53W06vSEe2/8fztR2SBa/0C4UNqSr0GGBllp2/JD/ybAh/31qd6ltqBjsp4+gDCU3sHij+lG8
3qO5TMnzgdmQPwadnj30xvxfHATpVke7G5Ck2JtC58uChQCY2xzJV0SMZ1A8ghb4CbnN4cf41hQb
h+vJsyNFdp6SHLvglRFS1gEYDhNPN/YDjGa73raQsEzsoad4M6ooG0/aEekm7Q5sdMjwF1aUydo2
WtFkzGqXHThep00Ym7TymTldzLTwFrT4vE+JMdL+MxJ+xt1SQKHqi9AcolKxdiEXwOQdLlzSK2xH
JEVYLGyDRave559DVMW8C4xGNN9wF2zvV/5I0hn/Y5KBszIhUQhUx31x+/1HkIrie2u+0qcxFc8e
8uoYC59tgrpWQrxkrBs/cCiac9NAE60neBoZO3Sibpwy27qAmvlmQKLA734yrc9Dwf7p6BHYohI9
IP1/dw8vDH5Wo69enS1DD5TpdrwexeycPa2eoNpPkAGLIs/j6Q2W5B4rh2V8bDQVuFnNnE6z9NVO
0uAI2z//kNSBAWZ0MA1Ng+61is6TILYyS15LkHZZxvgt0cCma9J1niz2cFzBnlRmRcibo+RjXIB+
PE8mUjNTRFTqksDlihwrwf46+HS6bUKfEgCqp4Pnwj5IFDfbGqp1naYrVvJr/v/otdYdBbDSVUj7
qHeyXEbXnsZ1s6/PTylws56lbsue1l+BXqV9NzBZi/vidz5uByHF65/3HFOrG6VO/v0uTpJ24JGD
uDK4nWwx1T/xK3jxjwEM9gL+HuDgQgXlVGCHiBmXE9cdrCzkZoL8bHqfK3TtH/HgBFzejH0fxCd/
u47jNJ96YeCU/K38Bu48WWHJyhWlGR2V1CVHCE9vxDuqNSjHRBjq85y92wpj+RuLWbIEVd11Holk
g9CtFt5e8QqSyWIwo4yLEd1dkoiZEq3JbNBmXZEAMfYINaJxtCiVh6/4kwVtsugFBzcdBbtA9z/A
mXl1azTR1kv1iRRdrzUSjieenv9/yZncAEzGBpYTI7FuBH+hKumr4airHQTvsaJNbS8OTgctFM8C
cZ/AAj1ZI35faWYJctj+lG2lpr4OsZqjDOWQpl0hPWEa6lPcvXyRI6plKqNyFObls8GxyCUyhGoX
WtsA0wfFv8rQaGSvbocYiPX3vHM/3ahMRbiuQrqPUcri9gak88Vrhdt+kZZIFWagdV29+W0Dhj0E
CXW1x5Mebzmzn5jZZOALh/cx4SWBxgWjia5rOuECqQZA9Vf5TVl1IkiE+U9ef4ovX7Fgz8Q5dDD+
B2oDQzHfdGj1NLTyuaoXCOXpBjc4rtJcaYcRDlC3g9sgAeHd4dZhZ4Gpz82/nQfY3uzs4pS6E+ZR
frLLCGl2+GgGpMwZuKyfxcAqkr1SNmDOXLRiaitesn6hSfJMxHU/DuzKkojdvOrOj/QGVvqXyhxC
f6N+3ck2MPlbYJbTPorXbaipQpd/VlI5yt3bY+RPy3vZtaGCQsWvQ+itsUhefnps8hVTrerVlLvr
6m1DvsKwpFtKXxP9jqzScfqSOwytgLAZS9etLWGki2WSSGIb46sEgrVJkkcp3xo3XNt0LgXQiGox
21OU/c7DkoOXsdVRLWpEoWEGLw0txFskQg/zaMMiC0IelzgSYVM4lVNJhKkXYpXK1RawMkdJxPr4
ivREXIRxaP9LF0DYsZA/trmb8ZpQb6eyRz7X6hcVZvGqKI5Z/YuEo96QFrvlaqaY2ovHXMmC5ILB
HwRwNNoe0xvpDs1IM6xmqZaUHRW6NX987F7DZnBchOXX+OIkTSiB31iMVd2Ird17JoTQvrFcRKv/
jS9HXYfRnLGvGgJ0fWYD0cEOhE287X2Iia9siJNui1DhRDPVz7OaT4sbO5th+pYToW2E7n7rVW19
T1NOV3PENsGJhHegfZTp36AcOPa7Hd96d7Wt0lovFnNoXf/Qlw8jrD01BexoF0y55h9CZgnR40kp
b7xg+y75gbebxU7awyl+xp5ik4ZW79nEKLHwEITwyKmoJwqcj5/IDTWWvIvnsjCkWxQ4LRtsx/qq
k5aSTZoPpLYmRR4j8blZe8xB37Akl9Wd718SJzKQepmdjkN8Rew7uVRC6WobFuG7ZBVxABjYsXgD
KuT04wXFSSSgflxOVLAGnWu5COJkVLO20lNPfXSs0Na33UaaD47JuAgx5RcZi5tbQr8tVTHjBXnu
S4mWbZ0NcMT7OLZ0Q5yCKYKFmipWSl6T5Vh/kdYiHnapHLGVG/Vkg7DUFWi6CmNSqooDRtT6ytsW
NEjDx+rJ1ycEhUEygH4UEJI2HnPE+8q1cgaZ1OQqZDOd0+INb/m1u80Ekm8txFnEZtVZNbF5AErZ
JdBTVzzh2Q6BX9G7cUuETIpymY9MDxTe59Bl/4+AOk4AWCkQk+aEV5EwhoD5jYfhpZo1XN+RGxAW
xDzfoh/2G1Dh4fsdnzLM6Jxe43EdlVVv+Qf5gKJp0YbVFy9pXlQWH/www/iRlkT/rPnmJKwWpmWZ
nblu6vTGwRGZ3FROT/HoVcSM4LajFvxoJkYDkBPMdhNWYEtf6zmML9nQKKkOQ00VndY2JwSVKXY8
k5W5riHMhTAX9siL91ZCLcIRFa5re8Y03uRPriFh79a7EHBbkvIBXlyBaiwEftyEvy/my1jtlCkP
VHuwO2xHlNJNp+JBYLaYmVXvnYzutD0jKg5GF1qdKyjDETCvMQKUEG/9GsGVoQy9Zo9GouuVvVFy
PvogCbqjKvQFL7RQpyDPx5/19UAxoey8jJgKNMGQs+hM3puFaKarrql54j6Q3w7tFafpnOoUl8bP
bKu9r64YKNErGRrPoyHXWW/7LxK2PgtVsd+7HwSMBDSni7/5vrM9IhGeYqQKO7fELQUNg050ZZxu
kpqqniXZs3Gsr3+YQ2UMUZVHXemxcd0kyC9jLAliVHOeZaxxOpongA7OKHu8dHcU4xiVI90ddvzQ
YacdbANc1fUrBK4MpLkK68VD1lBWqK+9pyvbgXxBmft8IAZOjA33wVbRUSHiId5FbLgGMdi4p+ww
dK5XMvskkJcLLIhCPnb358W8P4KOFPKxBPSBRBfnW/DTvmsg+EIxs57UOBfzqpRyOJdoIXdVZP9/
GnsX1rV26f5dEVQokZL02f2Ps2Tw+AY1i913KIXBBAWL1aPWL6rcW6LrXkQFkUKAQwDAvnMJaWkK
hD7jXpajV/8BWB/qeSH6WC9FQoM/kwrp0kR9W56p2LrP2KUNspbWeAh0fhTnmZdCssZIyGTJZneN
CmjYuTg7TCJkOyC0ZCH8FUWPO5p2Yja1UooCP3TWA9Hlwp94HVpjsncxBSxy7m1saEYUXUlznoHw
zP5NByAwc3Yyg70uMXuubdLxKCoUk9FOo5d4AIkjP4bnMQ4GW1eQ2z89wpc6WbhEbKAyxuaTTfPP
pqHEEsOPvByUWvfx8oacz3w+/xelULGuG0b/bII4UF2qTsZTUtLsCAilaL+O5KAPQ6siRgkA2Kx7
HNlrzjI83Y9jnbjQJfwjwgNZj+R0CxOQAoshhKDQkS5qlcL7JKE6quR5I1GlXtiYmbUgCXMcavHk
AS4WDUD9tVzbOEVur3XCK54w1sgoHM5sUCWzGMz0unZJCarzzf2nbbHhrtcbCSeS2Mg/+20ckB65
b0oJ2iVuY9GFustThVc/EIPhDskKrzph/Sn3bRSI1xm42VhV+HLZLFEKCOvX4mukiFx99rflTJpE
JCDVgfqgj69gME4E/xF7JrxYLr42u/tBSv3F756NnEj3tPA+DxZVzoMgqyclqbhwjl6Dn27Tjm20
BjnGJcHx3saqo2zUzIFula1bzlxKYyexdjR97oo6FeKuVzr/HoeXhxpiDlN1CkeK3oerJt/QdSIq
SIGTUdw1blrEaQzaKU+DtUFzjhQJNiXcSor7okTH/ZcqA4ONEB2lF9EYecBO8Nasql1Qe3/KfKBL
cw7nOQmGWp55MjNLceax1ZLkFsuQNL7fksdnk9ZWVRhE/9LrxF5LhrAOS+5juF+txnnQLFFEGz/C
RYj23yDDaP+PYuzWyz1cipimxyA8bZpzfYB3urKE1Z9xJnWgZLxMbcAaiElnVc5vA59d4Xy1UzzW
ACJ72SH2kqpPKUfnX7kf2gER1ajyJcEbK+X6imvd00uaODzfobMeD0+HKeXZqBgceXqIncgjgHk5
JsgUeARWqKTpyN4Uja0BRTAkHXAn/y60iKWza70ICyDXbI2AmNJobjESYNrAQ0+aCJ7x5A1v2nqH
TC/XO/GwQb3xhv2/JqQSi8IrsARW64Jxales4wgBoRQOMzpRdAGx+RQACi2qjFsHRCqZs++eZbNT
rEmzXiJPfgJP91vzcHXDDK15WrCU2kG1aCRaBCC2gyHaT/+iuvmywGdxDuLnQCTkn2pzFcsWl4mG
m6kSEJks4FMYWbZeqOzFYpKse3yCRGphBZDAuIEwXi/YrHfbFMAlOfRPcV4HWmYvaDzdSr7dR5VB
llbeiPEK06Z6gwQHQlaXPv2ghUwzFFmAktRiMDWTQdm5ordHPKIdPgtOJm1mlfzKAr7tYH2Jf+eV
i3RZPNfb2lOuLtM6avGRii404npdKbce/eseVQ1IkrG7e0StrqJsmNt54IcsDwyzBYbE7XKenbzE
aVf0rG4VKFbBgYOT8olAcxE8Dqd2Kty85uPP7Kw0ClxhA78EOK6NaWh2u+Q7udd3mflJZjF7lcy1
bR+GVbTTUVgsgU9yIGwDc9TYsAKzG1RyY1DVk6zSCp/n5qA/USAS3aIDV1uQtn0EWNnTZMVKy8gR
SVKKn7zpnGeX7rW5GCMk1fa5HDpvLUNpYmvNENGySWfvS5hCzZPEWXpcuw0fKou/2OH27y8NeuHm
HY1bP6NUkzhuAjHj6nJwNlWt4Y5r0sr9CkqBJZdZt1nxZUrGpIfcFMvVPnLOBdUwaSuaCL20UHZh
hJDskDOLKi0myjuqrVyDEs2szxf9bDL1Mnuo1Tywz4Z+3kH9vyhnpKQBMe68HH4evTrx8/aBVI7b
+B+WTJxDReiiFUqIdoQPXl6OJxAGSCoUbG+paIRGHUZmYLG6B4yERbX2lh3/l9eMeDJ4oOruGQm8
dmn0oYcs6QlVa3ZOUyERXH2bWQjZk361yYjrOXhnriyNd5zmsYDlOvdX07OH8iOAtvAtvEiGPVNs
/AG6vFsqeJyFJ9OQ5mn4klral++Iwsb1+5s1LyqRg+i2XNXtbQmZsjr7L4CyCiIxPcotnBWKPSxO
4MiXfRY1z8hg6cYpx+XsSCxLHJ8Qb0zDG9auR0tz86EkHpAsuleXRTyPkzR3oJL7gF4vxAavkkZx
SxbWfwI6mu8i6hxFJwOzhvFHFou6oX/JfK6szie1uS6FADSYPyHSALNLdL92rF0zUlQSoY2GrC4x
6JFC/17khE4WFxFKO+XUrAWvXkqcZpVeVn6HHFWLWoGldZ7FD9OMVQqjJtBJU9qy9HXZ4ERru1XQ
5tqF2LsU1gnNlfVWHcjw+foMJKK8Q6+TYfoEQ9oWWqPedOnK5Kn6alc7pYm76eQgxFKY8KNXaZmP
qaLhEahjkRKRGdDay1clHyXmAakhIWzYLmkK7mFzurzJcUDTEpzw6OopSL4VZdsH8JPg1VyhRo+f
3vj9hpgQK+w2b/ueOVbD2GFM9FtpGYWCsjD8a1ZA+W9jD+emm9Vnl03tW7oTwsgZF+B0XTL28bj6
a6KvgPew2Sjdcf9oODVub3i6x0PciQrR5SFFhsterxME3sX2lBH9gmwe/VTyyBvm8RU1U449sQhs
urTw9zQhgLvEveRDIyDu3D2AxP7e8SEgUnrYoDGxRFeSQ10RjD7FgZYnG/hoIB0PAV4qbb4XsDQQ
W3Kh+DDwTx0tGAIAC/RghxICeOfMOePhVI/Z5q3mPsQAhP0444ZKi3AThzPjP1WOezc0ytiZyzIj
YAn7KLEqRk/GKc57iXf9lJLvOdMiJmrSfSLUEkpnC8GnD1Z+cJubTrMPmW4ZjvYUd4ll05UZ4YR1
514jR0pkeWCGvqhEWPJITbsd/87KJ5XpSPmlmP4UDrueXhiuN448JvA9eRvB5jT31A3lGGkpxfKp
UxYIVqkAUmPRXrVFwdJgaGTZv1EOlbMbTz5XPTnfHjkQH3yTxJu+W/pt1+dz/bI10d455CeBBmrx
ZkQouMO7RoULa07qRv2+ocJP7Cmb0pIaPZlyB6nMeNsz9ElzlkkCBSyiX6nF3bCD85EmkXUGot5k
0w3RDcFgCUnUZbMsAn5ze0r2PNOp3GV5WLn7epdCErpVRbASxH0fArw0rKjDkKyMLggUCtpaOjlj
mDiGWZFhsI8mG1S0hj3GCPjtXry+VQN/CKWv+K5486x8In2q68l6hypXXyk3LANQML+JMYENM4PW
kKdILdk9w06ZHwXYb+aubb/GvggifUPJUkS1JmfDuV5f8nxyaSDEOJ01GWbfnr/Hq/6RnF6C04Ah
MhnSTKEWm8wNYBOMU3Z35iFZM+BUXPDzj+BdBYIyJfHKO7cb8XLLcW15MzM0KqN9/3Dq7h+04Igr
NRtrgwLIJZgNiOYergvUjn4H3Z3yX2TRbA5yRSOl1YZjmVkhzIczD72l5zBqp+zPITAIGHvnzIOl
qNnq2wSj+dO+SeWWiL7EBuEANNeMgMIDepx8xr9RVard8aiAhGWnMAkCaxagdPhS6r3ktSnA+6W7
oABwPNTGY6R4KwgyZTHmqIcq4iDQ4IM+eC9UjDwtI/1hd3fi3iHJ1ZNbZyVh9neVIGxK6HXzgW6i
IUviYw4Zyd6CvF0twr+jjD/bj3EVcPgQLhs2O8r+EpGAi7AX/kAcoQZILvqd13nCg9d2mS5ZSfr1
H/bIDdxUr+lkcPM8m8VGZkNk5dyZUoz3dmkRSZZ9845Iy3fb2rJ9Sc0GGw/ZAEbaqcsDmehjDCC8
eKNePq+yE/qU/G4pmxF16Vm21WZ+Bms7WiQbiLQDzixvsbUEyK1USL0mxK7nP9K+nmopnxNYCrVC
QGGDwgpOpb1yhxHCVvPgRKCKhblQZIQ4Vf/mKe7JA0tB0LUT1Gf4jsYo5StAymdBzL83BOIWQf3j
P4QJa3MwbpkTNl3z0FK9bc2oiSFWZBu7N6XA1xjpo1HJlN4vMjyZQBptkbM5/ndoj9ZTDq3u6JZU
huMXYIvM9IoXPyXW77K+72Jqw1ArzqaFX1+oa0FO93u5BZA3NK/VKjWPtxe1rQ15LrJWaxDiR/Zl
v2ak5oTn5Xw810GluhTQ3D39w1p+5M1z5OUXkhmuv8IHpc+kI8GqQXIgHY+5LnmPxaMQlaJLyBgG
SCEy2PHu4YY8/gxFcvTvNKg8L9rPJ4cjWGATo2RfrzBN7UIbIY7oNF7ULj1bCyA63CnFqXk64Rka
g3idOodsqnnY4xyGrz0Q4+zH72/g0nOTPUZfXpu0KGqUnLf+5HpFeCd2P+Peoxh0yFbfeIsqtfJA
w3lw6bEWswFPMYC4xJz5Mbdioh2k/lHQzoOh0ojJncf17JBe0gh6WbzE22cv0mxg+dTYXoSxivsM
W90UmogZF18p9eXPhp+J0B3WU/RmF+BsW70ivxHggEbYd5ZaZdzcZRkdad2VHIhHYLYiyT2He+yf
hBNA1QyA2fBvn+BBHTcHZFlEjym8UFzymRvgx+Rt6+V0/3rJk91oD4+23dZFcZDHxMI9fRBRcaPr
rQ3qlBWuYZXkmMqMFQ1gCdh4AHdGA8PaQOqThY4It3KiO07gAPpBkH1JkIdqj/riUh3Tkekedffc
vHLwLSrlQAH4yomORaL+I5BjqwFUp6sWDmjbgM+seOWAFzJbxQtbDRy+lUw3k4eFnBIEQs/OqHAz
66WrBiER1K10Y94z3B/3uIyWlojrLhWVYHHf58+29GH34g6ciHDZ0T96d8XGdagmowCThUru0P32
T85EgUj8h+ePgXvlomWNNlIWCRPBgE3PXwS1A+mwMCxE7ksOOG+9mp46CoN2ILoe/dGS15nj5e/E
fdbM730jjrFxaa0a6JEXfXrhOUqmBp1LYgV3dVeSZjhjPRTFjrN+rgciBuOcyu7vUalOBJM1x11V
GqSSiNqylYWiLEeVRjvjInei19c4lZkUqgLHfMmFAisFHRrzn495bJ9u3SKapkrrmfjiKObU2ZDB
jhn/tGfnqsch3kJ/7AV8Br2nh9L67BHkHiCme43O6ayy1jg4hDLNDYdBe+TeadBxD8ubrNdkW/g+
MkNBRhmIUt8tKmIn8B16Fi1sdfdtc65+4kDLGJAHdoPSPMJ/pgLusMwJh24oGhOS5mY1njYsNXpn
3nnISj9NZfYCbKtYBgx0vGRe7MSPGblgawoMOCdtN+kykA6yzO1Ic9wXsbI5qHN+0178TYYVvoHE
Hd4CXcqBI0NvtELp3HKzPHq5P2jb+aYM2PKIGKhkGZv42pHV7mm7FCp8M+9QDTX2lwLsoIYItSh0
j7HuVUHVGRYMuOPQiBjKwnJ1nVK6bM76MD08wTCBABN4byNnCXDL3WXouXFkTwsuj4S5NlBMTqFM
dB0bHrx89TZP4/1Mn3uFqgPPGfq0hIcK+whiiRJaU19Giu/KS1R0QRiB6vqsdQIVadKpTOnD+Mv0
My89PXyNZEIPcvEsnZbWu8xiYzY9xm0vh5rXcRtAg4DrziEOMMkOi1LYmWm7DNtsRXYj+VGv9ih6
GHCZhC/PsmvkVi2wT3vwi2NkALKYJRjYC4TohZ0Q451kGvO4UgZ7N8IwDToZDr5WZh6J/r0lER0R
HBmAO9qwXSOQlkeoVfihm18ywF5qK6enbjsPo5hSpBATYW9qPisvPDVLuwOVrqyjOLLJ76/BNXjo
N1izjrJh7vPKT19geFuFiDaO6TL5m+VGpskRW2PhTBm1ZWCVP7nWclom6B0m5hhvfYcchsdChVP+
VkyjwaZMkBvnQyi4V8CDcRrciXwXrgsYrXHAtPq3y85uG8z8xuEjf+dvNC1Kw0JBOqwvkBA/+ESy
jL6t87fUOtjl3vCFqbYBiLuIT+Zvz5kBBrLX/8UIHplUtYtj/BjYTRy4JZE6k3IMerc6e745Imi4
HsnYbo0aTiCOw+BnU6xlrRA6u8/2ulGXJAwSsPe2Gc935RBoAtmxOhFMczuUJ+4CZuSkJIh9SSCg
Cn0MHFF5zDCfxPjY/CyPh7Qfq5ZWM2I/xrXtKzfz5HlDXmF3RVnTYPXwz1MsE1YwqIA+Vy17GPlI
Ww/GWvPb9DGPcjebZoTuHjv08YfZMck1kd0exp2pyyyRFeIruJu7Ll0lss06DN4Q0Hn0xk6WN8So
zvig7AJ3E+kqS5fbBa5oSBwxxJTl2QDMf31557Gl7wY37NU26jwUghydJJFZHZo00afsMz2VSnaM
TsLOOGwKGu2jRjLcpdTlFvB+OubsFe6LEcLIi6xu5FO+KUjwkMvMkK7TfZ9g/Opcui3lxBAqyp46
CITALk0+EZGZW1uSblDPBRyQJPGNO6u6EI95fhgnVOo1MCiQE6IZ7N8GKugZ6wHsuWc8j69HrXi7
smQ1+vV+1ThmmUaKHScRPjerTP6lQrCAiA6OEZ1e+sy0jMV/d28FFJuuZyRMsef2OlMZN/fo2lcu
ITGMZaEX49Mk/jkKfskqj5FzubEMW98zYG9AP7QPVh8IbjWfWOvl/NixFApUuU7tPmxkbc5sR+Uw
jZM5rtIbNq3fBsc7bH+rgnTDM4oVDpcYkYgfF77LAcDhWRI0j+btkLSD3PixogmPkElDFEJOw1Dq
EVdqHKRWh3lNfvwyxLzQcQiA6YkFjdr1RqoPecADGVtQlHKbrKsGs9tqmuCfvRWk0mKiZWoWPyLW
YTEZf1+lQAn1v2vd2KZ09zDsYc4D+kbkUf2bxG589J7lPWdK+LpzVh7dFVCImVE+PoSJjJsFElNa
VChXKUlv8b1P7Wfh/RSyGAV05NgjM/AzooyuM2fpSDzTV82nLYwvzE3RxEcOgGNIzKJSqph6vFkS
9AgDj9EN8xl+kgIlW+KFiJUYtskLFzLLQIHj5oPgYn3M8ViXB519HIJH8lXEPeFE4M3uB/r6TAjJ
azEqJFh+50MR5zG78O87TzBjChA5JhYF61afuyL6yMXDQEqIfWa2bjS9ureIJ61VKOo51yJ9XrUa
jLKugU9zwhewK0ct/Mbaaqp6GlB1xaM+XDSwRNzFfCWnoHDGPRxE+JfUVg/yzGF92GakDiAG6f5z
p1qr/tM6yMQpIkCM4d5Qjp5aVpo78aOXSwvdxmsNmYnNW0IgVQYMstUKQBO3bSWHngDagWvRg3ha
eFJTWNom/wT8ubRWcnzrzL9neXJ5Pt1mw3pNfVs5w6Hkm/iyfLD7UuC+GLok9MOozxqVDOFv5SV5
wV3c/jQEG6T/krXqYYmKgfULwNs0QJxq2ugD6iTX0oDlR7EQhMT0aoUYxwQ4Y2llAFZ+qz70O8r9
poCi4yz8GK1cJhdDl8hveOb0CVJGPXnWODfBbNHRlfHzTP3/seP4e7VaLhowLOlQOX2jUanO/hwG
J2uUE/KG8ftwPSPpiMHl4QpTdcCO7peWucz9WfuItDkD64LQUHTYW2hpVIWHbOn1jWFg5EST9aSg
zyXiVJ8+rxvyhDBY95WIqcmo989RkWE6lU3wBo6BmaNaSTj3VMkxCYlSskf3V59P84VaGX+B02dG
np2Q8HyZa5R/Ysuacks9JG5uE+mdzSWqXZ+a8ZcH7i0vAdhA5+zTWkVGS7ffAClWsFCSwZVLpaUT
5YmUfZNuqUu27OWItmMWAfllczUqh+L87hzhJ/tWN/R9Tmt4l+yy8MZ/aAH9KqP6Mi/uyUXoLVLg
Cf8b6JQUz59j0DghiRAecrFAt4TbfQd5TIkFSzTk26AeXxyAH/jw9KgoItfmTE1BHCZhvzuPWhVY
cyyk0yG8aXFT5lxzl3S2kZhsuMNIW9/gcLkcFqU/APry3RXGtMFhGWpJQGKRyYP6OPlotVYPvvbX
Uc/2jK5yMIhUMFJ61H8Iekuk9bNOAFUCB++VD+gFADrbDkWRpQNsgGWkCbfNaMMcjvWLAh4NAab6
N+UGe0uwGAdbkix4JGrsG+QulXJVINDtJILUh+g1jfALu6ZpSnqPRWRaQvcVeLKvVkIYoBqkkdfb
hAQz0CufFoKUMNMPJpYiy2ZLBcnBAWNQ8lRZkS44EYbqK72Opb4qSCAzVzHOeG/Le7QTlG7d2Wni
UJJ0XSc3cwHQ2Z4Vbq9u7v9eH6OGYYjKyIlhBf8ZgMY43DQ86iiOb1bmihJ3A/CIUNZbe8Krw5y+
Jh+3NLVGORVX9eUJDnUKaRt0NyibYvXJEFH2WS3UTEoKWB/GHLpLC6bOhN4NtJFoeiCLqmf3BW31
rbuI5SFAZqacecQ4FfGBetsa4gUvsZeEvG9WC4kRq/D2hVioXoReTG4qART65ZcdpvW7foobpRzI
LOsjdXF9sITa0n7jQmp/vSxfKNmri2LLpF1IXxNuu4bQhJIp5Dv54JRQlPAgmLZn/Bs9vy1vsqCo
sIAHLpZ3YZuHuZj+k5XuzPojbuoYhH6DzN1tN3e/KX+4mWX1/XqZPiYhUwIkuKDLe9PmCpHWfQlF
Ktx23p2zsgUAzPwAep31TXjr4i7h9gdVH7Y5+5/HyGxZ3O/AhiRWfE+BWUEDf6QmKbXovfosdhCi
I4nRHCUvsUfOqjsu01eLCn6yk13/dmBt0QYmXyRQ+Ejwu9AE4i3YQcPF/Y4DDPfuNx4m6HA3lBAC
ku8/AFpyJ6twVWHO2oaSla7zLLZDMsy6XMSpqu8qvGQ3jMzpjtAtoEDUey+g437TZV04LTjBUNAY
tg/9uwxnBZ+A35yviKLSSjyivhPtHVAG3ZdeKhLJHVJYQVcOJ0NwNYm/23NzE3UP4XovIOFFmoRj
1gmqKfghnrTq7S+yQGG7c9QibyNtr8l8/d2gLEOcabKJXafGhU4jd0zfOsEteiXMYaDPUGPc4U/n
ybBqgRYKqqVOot+/kRSvHoTALHb9xcYdjxZfZXO+3JzJtA9Wv+yyQZa0+SVHUkL7YBE4mcn8pwBt
d8/zzC41wQpvoDNzlMenUG5QFCFaZhbHNVzYCqp0/MouuJ+sejHa77hiQjU1MtQwXw9nQmRupYJg
EjC1rppwrCghQdo+sQW31tDeGVyxgbow1o5CObIEulbWNK9ZnFMeOc8adO4azYkvkqCqDvpHIvRG
m+IuMeSznZ3A6E35eBLi8G4EfmFOt9dzeoMZh/uWdQ1yvlkOrU/m4VKeD8SlkoL13jNPrWw0MGHI
wbVr+NioeVol++4hmONJyLKukCPxI/XUjZt6dxRBCGAifiMxZ7o/vCnBoFQNHB953JSEA41akwR8
iGqYGk39qD8cOgN1cqaTi8TH4jo1j+2TAU4KgRtid12C5kMpCKTykmfUKeBEVuJh/6zpFvpg6Wdk
3NwyrxOPq0Kgpt1jRqKgBrtTmbjwxtZT3SNMNEhjOc+hH3lALAT+RrphwX47alrnG2b5hq0z8gP+
VZnPmzKDcVeQbOxbxJvgIYjUsKnmIo3lBccU79wIQjHYDvxvrK7VAC7JnmZym3t11iLfRgRpXcpm
QiivwtJuLYxx1kiwUYbYjmIDrdsk0Y/Hpxq5ajFSEgdGZaKzrg3uiFZ0Ef8CUCERC/QVfAPPreAU
tOJuITtOfCvTZPz3ip60vKewS7qrlG2+4glIWGZnSZR3C6Dfb51qePaHFkfqtm4gntpMJj6DuBQo
JReDK4fKA6bGqnuehpnzuce0Seju3v9y6dxbLsGKbwu9VjPthQnFEYdAX5Tbs7jr6fo3UX55IO/G
LkhJv3eLhFBVfTSVbuxUlDMzZt8Pby3j/ACJVbLlQri2yM40jUQ6xdGKP/iniBKp2b51h6ioFVSo
aNjJ6h4crdc+3LJNUOqtC/Omxl28uSoKXl9kOEySwv0ShEWQRPdg3kcEEVgY8A8PWEZRktsoAIDm
jtkZhzSVqzbN5fQ3fDEn5Ijg8xDIduF6KdprN5YuppLq0tdDNGPgD77PaJukLPk3XwlIJ8SEvWe/
iA9ydI4Kt7WGO+llC/i7JgZraKsRt7huJCpYlJyImPBnPO9q0Frgy2/EdU3+Uf3bs2ZE14xsxkSW
a+5OYDv1O96iX7JhVHmzgjVNnF9zRtjAzH0XkYmaVijOiID1weswMg5CyhJCJoVDU6cNHcnIq79A
OB4xYoT0uFqotekgbdg6xTL2brEXr1t+liOXO/57EZ0/JywQGx9A7vsPrduD6JRo4plMW8w7/9K1
0DPuT52R1BEep9V1AgbfAPtEXLKSF+QgoYshk25bs6zgq8KbHJ2/kdri5f3Equz8IWI4z06Kv+AP
npbpqCpoUq9zqBdsGMY/GfJnsRxHsvpvOZuz4rRyP6KqPDE26dtO4oJDWee9s9BQ04/7w2kYhraW
a9u1xHgr65aj/1AlSUDveUaz5AwiyUIcFa5Rhn5STXE7DeNrfeIXtC+dVdqg3NR+U9UzmPAS4auo
XlmGLW598EoBtspwJ6mar9lo9AHF4/7+ct2JZh/GLJG0MDixUz4rNXCbRU+z84XP3PkR82VueO56
Zfec1I8c7WHtwU8VoNTOzBErArepxyEU4qNbYHXaSxCUmqo1MX8DG0KSUplliwR5uqdeJ/TssGWL
qgzfT2uXmpY2jCB78mcOjKPSwNBgIVsxF2vOsTJCZ1KRt407BE2TU3HA5gqE9ndSC1aGF4zrIvZ4
ABS/tMhaZtVMNssucCfqyQuipgVO1/byJ2jIssjI7tao6WO1RsJTAdDNx8k4fuD7tLyVce45oqtL
6NFqfkHDwsbTSVU9wxTiXdHS9pdKo34kitvmt8v4ivLLHtmMqI3jKPQF9I/KG12tZzk6EDhY0GVF
kza1V+3Jh9y/CUEmHs+0kgHx4Ske8bzNo+EY/tGfcJ5HcOwwElewQBfTs0cBPQbY1j6W3646+WAa
v11g/hvA12GBYKtQhSLnRXA57QAnngyWypf/b3FOVEGmtBvKiTD/JSrYGiDrsEZw6C6qF/wMYGIz
vDmrlUCCgpgKE6ZIMNGHNhWmaGlvY+rXHPSVCNSYc9A6e/gOzhxqeqtEX56wF8wWIje0JM3IbBLK
Sujgm/R9uLyof7oj5cS/zIy3ctZSG2bUkWAKiy35o4DEbNB7URLlt2JDy3nYn5bCA8U+uvGSOIi+
f2VML7jo8p2JFlUdP3nBGBrPHQyhvLcJuNB4OFDFnjWB0HU05kf4D8Mp9bus0+nCC7mottbEAi7M
cknId/q03a0QJ/VKloBfR3mtxT1TChLUoja5Ue8JG/ioG9NoxFMD4A+q3HQHLtsKwxRB+KsLon5v
gTIyzjnX84Y5Pz8UlYfx4369foYs+D2RXh59oaxktrk3L0Me9qkaonem8HYC+RJ5YRySqHmrsfNQ
3H5t/I0ERNc5IvoMGFWjRRsTD+ffyUc1YtLT5SiSSi9EqQY6tisdVqHnWQbkYrVbKkAfzzmCeZLn
g33O+vlPB2nenm6J44zHoX5kOi1jDg+yguKFeeW7LmWQUmAeexLqld1OmOD7RTPzaZHM2HL/UX0M
tpEwb60JWrDhfySu0mlCayQk4Ym3SrZ6BsyAcntJf1fD3kl2pCbU0a4v58sYKeU/dhg4yeBW+8QY
QAPEpXbqn2I7hA8MX920EFspjL/Vze7bCNpz6v4mDA55pw7iLl7BOqSvEu6nMqf0JrG+pWExcwL5
5EEPinmNg6cpqWUDTJsDtgeB0wSU09kM7y5TM1Q9I+FYEONc6t2aqayTsLFTGfWRgB8ealMdCZGX
+ZkIrA3rgIy6qiONcxSBz+I8IUl2b+nkAhMKK/NZ12RgXuF01soTVVj6TnvbWEvmAZcksUQuWTN/
wWnZxBXQsvYrfUoYM1FgU0vN84bUQtQaw5D2ZO5czMhxthQo8m3sCMrPlWcLBkjoITQsuq7Xq1U8
FsENnXC0mys4HkDdeKGlNS6QYK0AC/hOoBzCeEYvS8BWpMn8O1xMiKym56p6FPP2jnVnjeuGDzwi
cSMFPZ2jOO5q85xUlELmqAymRCjFKDjKzTaedkLPjDLAAxwhVxtlyoqTojCLHLbYDCJYvPiGgUYv
XqL8ffOsP0y+PmkKidHUuwX7IxUvkfzds/1HG5FHxNw6VPQzFQFK1r6T8aEzBROUv5cESzutwdEv
Gs3BkYwgYMaAiXs5kI0A+oHM0OqMQPulmKVff1VPSNEO1dfLe4dyD670mJPSqWSjuFc7P2PLI8M3
0Oj9uspNVG54p0RvcBm96MuyUEhb2DYvu4s16cZby52hiE3UixUKcImpTOjkFjyqgIAisEYLTePs
nFhg1+XaIZjTOnI1Oswc2ZF7BZ5tNlY3PhW4MlvYb0dTfU43ZsDdf+cZ9xJZaamSrU/3fwjSQwBy
1hKdijhlbuB2fGuX1qTLng+NiT3rN2TvKGKwdomT7DbI7NmkFfv+r/sEY7WGhb0sy/CI2cixBgcu
knO4BPS+nCVO2VznH+pYRPQeZ5h4Z/K5HZSqZkjXkteaKISIb8qPouNpnOjlaMH+RqUwYxXaV06H
PTNa5XDf3frFfswqlKSi3qvrm4MSrWRhXnjOjcYT7lL6D9Xyfz8srE4ONCG6b6ORi4GV2l/OM+2A
ZqB4P8IU6c3XmW6c8zDuP4ZnlUH5BvQqgXYWoJ5JDXtHIus6NZvrCxVtqoqpxmM4XpQB6unTNyL9
oI3ip/zmftSQTItWnnRxQpQ+fuhl+wMnK6E1wOWBMWbxupMHyinRYpuxwSpbTy/8rDlOM3c8l80V
JiPHy1K0uTs9gwtVUhxOhuSdlLogs/dmBLHNTLTEVnnu0WiIDeGkDeJj8pbI3xXLpFe85W8BoO/1
6KIM3JjCFQwZNj6GxwKN9kXRJqGqokFBJpleTJPmM0ja7KxqRTluKJi0aJcQZ8g3IXp86XiTgNZ9
QnAxNxga/BPTP0hpaQ03hnzTvKwOc42p7V0MPkn01T5kEEPgdMWP3hEbVxSGDBDK/9eh+rdSeFCS
jTRzV7ZXJ6mrlypaq5TGi9OaTKJrxMY6VEsioxjQ211TILngjoZQdEsCYp6IlsKFuxQml9Z5hfRE
PzREnv4aI7M3GuU0THEQX5eV8GF10+DQFgSP+00RW2dg/Ie2jBgmcUy+xI+AAA9ziVCwalC8eUrJ
fvEPtaD2Qfc0Cumd5E6Hss6saQ82LPwepXObRYVrB+FwHgOAC7TUBWYQSEwC+EqXrqEiGBl8KlrM
STPd1J27j/ilIOHvlTXlO5WSgqZTf2/ZU58fkCMBpmyNGidKcsfDoIKB3PqwF4yFwY7ncCXyD22V
hsJhrUJyHSz6essuQ3ZooOtYG3TbHN+MYmTKZAj/pxu1GG03s0TtlZ1IusKjq4BMPqfSlDqfyRio
TriHxZ4TgiSo/JlTWREZCgiFhMbz+R6gnEuzfx7xYupdwYdHoOYoml3jgq1o3Pxbf8yCZVQTS6sC
uumpmVHP+nqA5xxk8vjtb8PnbT+QwH0NCN2vzjspEAWbz20GfhFhhC19sSevBwY+urXpMMXoHZSq
u7zdbjSIPg5ZGK94i4t3OX1RhvIzVRR53wESYNYCAA4dmGD+XXaPaVcAiPN6WUw+wx7EUnSqupmX
dSMO8RGgx00ttRZDGHBrSr7cGazY0sKHwAuKDgcre957T0khczY0aAvhLUlNEzIBOFSzRPqLyH2Z
dg4r1246dRZUsbqc9k+/D89pKg8bHqGrv3RZPwbjKu49ZRADe0kVJC9CMd2onSnN5NN3uWCGhtyJ
q0AbP8G1ISo8r01oQeMlIKL/mHMV0HjFWQ8qMKuBJkF5G1IrFVLcghGwOoMjHOdaA69mVAYMzHnV
+CRcwKvCv+ws910aS8TzdC3txxiGQ63dvxqrTi6MCtUvIB7EbVtX16YtFBSPKEKuTUbSvJew+FO7
zl7dCbu4mKQCoPIfvFlqb09YawrNSUb7IeciNPo1/5y1W3JupP+8iEw7eUhNJEBP26q/ht+JgbM1
oPEVyaSMqvUcD/qUWWwi1c+1wR8D6ZB8pT78oPN9dhM2b00tjt0TK1Us/mpwFmdWC4xuOezTYD5R
QUA4xiWftdJExVXmsti27NAXzLWZniHBrp1RiX1zW2n9yYjkyCsUTrzAGtZDg1PJP0a+OofZN2R9
cLjO2iFG48nU6gelde4o/he2CPHhsDfP+uAO/PzozkTzyha+t4K2hFOZrmMQciiBU6xQKULHYrYw
P+CDxJPEl5Epn8L+lJh4eNavE2E/5cPGfyEa1jRXuKPZch9x87MvCaHfqdbCRV1vRn01pc03ci7w
LlI55f+Uva6H43Suu+LrwA2ICnAxBwJehrLOzL286jeUD5ohdCFYxkhLcuumDxuxIq5Ac9KL9iQA
0jXjHFDVijB/yTFEU1dVTft2NgREC6K9xvHtJ3vyjTqNdl+SSVRuzP9l5CFjjMg1hAdni3kU+W2y
/FqK/p+7i1N35ybabealybN1cvjeZ7Ez/YUbcRYM5p5h1yj35bJLqjpCQEpPCI+Cy9DRvnUyUMFS
s9CHIDbSIXOOOWTQArb+BGTBTVTjSy+k8L1W+OTkF2q4LyDWTYaRbMr9+Tbx4yLqiLBjaBrYjQUQ
KF8TNvsfOy4I9z6vF58Q6KjdN+Nd3eHv5tTfbdUzfTtjrWlIze+kUxmn6ziVJQa9qVQ0vh7imNfC
DeLAgxQiUS3O9KmKEOz8lXIjayG8BpqUbX+9tG19aoxMWjnUK+fTL5Y/KFikuNzFmyO80swuEFHl
zkou+zgdU9TdATUTHxGVg8bOlm0U5yRlaEwLZW3gIVeNVLTkvof12O9s67U26RikHexOBp4syOU7
vHPXE4iKF+x1UzIMctfQHlanTS69IGGkrVDnKIxnc0VDft/CWm4NS5AJ3bGI0xZsPXjKxFrwGhRS
joVP2brfWAlbferkuOlHB4BAVVCmihMhh+66VIvgUNP5fQ2SZItSZC+NvJCmQ0l2nnenwm8/oIc1
ZfpXuli4OohXEOvAQzEq9tGiapomLQXQ71FIZF0MW16ojUkGBqph92vs7fhJKZhY8rNM5cvGVwCr
C5pnK8ng20aYClh3D9e+Flqi6FbPNpbFPitUgUO9jKXuXGRL364bBFlocGQhBxcmRIZRFr2NjmHM
AE6qLzyXPqDmDIzd1F65vr4MuEnuehTpANxar0SYoZatnl/PMpCldCjSxPOpZj/fJr5oPDvv5oab
ZEoADfQukbs5TjzMwqt1NK3pdZS9YrtjX/lNS+blObQa6GPRc3ZY/Kykp7Qovv6Ex3r3WSJxAG9o
rXNfHFZ1CTlK4NqCQXdhxnquFBQYZQR/GpS51lUVQGLalP2VdGt1Q0W/ddP5aaee0rOo9bv8VbY0
Iapi+QW47eIauC3TPW+k2LvRPZPLk7/TgL+egfaaxsodh8vy4RIayDBEuPIBbqXbeSUScyJVJj5b
Ao4v/CmPGgvi6/nNRc8D/DzitUT+SE62JPVxu07ruREDrnvhqCYo6k2ji2xc2YQSBbMcusWtpcln
JQz7yHKVPZYGqhGwUuPQcVoPFRa/Ikce3k7RKEME5VN9yGHUgKkIZLKdRofpdTQr48h8qNWiugWU
nxMJTblQCMvHc2+HCsKLuYtOMP0nMUvjkp98OkBqIXBAWJG3TduWerrroLGMocUdQMiGSJqQlpPD
gbo3JhBn6KTlvis5WtsbIY9MvK5GSpQy/8Cp5LaMEjDVKCNEpdlA4m6jmTjqjLTxv/wKrD0EhHDP
V5wJXq4RcgGAom1bqSEvnrDk2w/nImYyttoiB0VTLbPSmA5gWIQzpqwRt9JkPNDy60bux5EKP/Po
FEbE7uJy0XNVGdXbXrg3d8HytjW1tFTLy6FGUwObtCfQhzswaW/avYEFvV7gWPKfNwCIxb9YTIMF
J4lpom/O9IWg011m9bPorvSIJJPrQTokhp07TqKREp9fmfqCUo+Mq0i0z0ZZjceToxSnSvtUa+L7
rTNJl45AW06ppPYHPbT4rjUGAnf8YL9n6wfmeISddIZh+nnLk/zcnLJ/mLzuz4rsab2/Ev5NVqtF
fN/5qsWHLMVXXpndV4o135ytgD9laEqwWpKSMO3PIL0mH/FscYGbas2P0q6ECCwdy4tQLvVG6d5M
vLlraOPvauTXYmJs5KLGt8tJGlOfHoXmjPUnGMHgmRvu/Ktu+y7GP1ECueoHYClFAwz05kDVLf7L
EA8u86cBK7hYwWfDj4HkhH7BwA9pdAayE5h9RUmhj6m7Hmvv0Zi7quAGFwYmMbnyy8p8Tsv9QiOc
9E7U5uAdS4xfELX90kknxCIU9+w5ln//JvJ6Yv+4RY1Exan9PwKb9CY3TlSOPY3ZdVNefh11PxR3
vPktC6t/z/y2NUz3cRU+IXiaG8CaQTo/wItNsRrjBwAVEy2isuv/DaTIecs7u11VDxdtabGs4UVN
tSfFOukpwdCSidE86/B5q+r8a+9eQCGdaTtASg8YL7bA4wlb6axd8uzbmMwBuYKDvs3y70mqRQ+G
rSi/zdyZNwzunP/Ztu0rkqEUxc4b4u+lYmiMpvn5Mize+8C7kNm4TmLHaBhB2L6CG05T0uC8+xs0
MltWjax0K6c1SIBQeYf0sLX3C0bQA6u6J5XGjROBwYDVJZ/n+T/zNmiBUPj/wzkRIln2+HXb2Uaf
Q+0eGeLuHh63lMFgtMp/pW52cFDObkfQJ0yen3MU0s+vzpWvl8a+71Iu2UecIGMHTwgDn2Vkfsas
IVpnGcx7StxOnw1Ps+xQzxeuWvbCIRmQwBZ7Cb5MkgF2+tnrqbtZHF+7iZ7LOzUC57LpbEPiT77A
xhmfzEhKvlZcW2bNAohAycK1ACDLAn2nMJJJllZpUFlWjtt2yI5/W7kp2tiitgHnxUhDee9gRf4b
HwFWGMDdxB4tz0fSs201mkzai75FE8hy7S4IqA59v9AuyV9YK+MFLrfrE6MxXBvn1nQRbZGfXTVK
QrdfP65FEeXJWoysKIzgWq9q1Bz+cqLXbdX+6q0JJqFJfrB36u/Qbwh6OKQLCDUXmPMyYADmMtdY
i0VIC/BCj15ijwkCZSTQ6cepkXpp5TNZ7PxEm61riThGMArs0Kj9EYU8KhyVNa4zzfmobN61lTTU
ucoxe+dOvgt/LNEs96kq1cyBZMKDgGlTWb9XHCFvU8Z+6qALgQjd3H9Z7OnX5qss/7yLCIjeil2k
rVm+8eTd6sJ6DsKdn1QgfBCB9edoTNhGQdja0nlY8zRWsTiaM7Epmrzl+b4X6j3bSvMQxfJyHMdt
C0ziH+8W4Sk42BaHGqwzevc6V5H3uFrj1T3eoGP0hVgDnExgpjZC7WmohgNzmkdUOV4B6OhxrSdx
ZLdjd51Ehd+SVplwIGWUSxw1c9CAcaMNG3Q33RSnhIkFswS/RDe4GN3YRcIfWbBZYnQSQby4iGFO
etLX+OCbb9OjrU1iKmTck70JVC/oYseT7kVgj6U7S1JA93WQgiJYvg1LOYSb/u1yOXj3y2vQWy+1
1m0ucG0HzoAhnCVcnPvdJrB8m54iWHkMIHapyYgDEjcwaBvfjZsOcs+i/zA3sUbYBN0ekNQbm6pQ
+kMOyNqlhZScyIrtp0eunYYbV3NtS8mzyX1uV1rdcVH+EccR0MQO2fxFFG01mJV6W+/45FC/zIFP
CmJicdKC+24xeM+F0A9/j5G9B1UskRq8t3yjvCPZVSbIx9ddZaO8wfi+jpml8LIKuxvCpEdTVvkC
+eWKWl3GTzmxSxXZjk24bGMrRPAyJWiPdO9XeqA+vOnjiTkpkCJkuvETV908ZeFskdH/TOa/CLu1
bD9uPEQohbWNaX7cS49Fs/lixCaa6trxPqVTkkWjJ1T5S6kMJ4VmPlh2cvCrkgXG3xMxRAU7tRVY
OrLnOtz+ktyxz2uac3RYDKxv204VFGshvvQeKB6x1c7rC1f/4mKLoYxxu4g4eduGAU1RWWaNTVnv
QspHsRiT1ChoLdOYg6ig1QSRtebL106hjRZMl3U+ppEh/c/AQ4ZugqkPTHLFKmPM6E3ahA3zRMsT
0lFmOd/pHU+VFAKD8xvwAFhRAdK3QvGw2vdcZQfnlkFhGiJmy/GxiDj8NRvoHAvBDQFLwNcLu9tY
VolFmWxZEiks473UuE39o6s7eHaIR/iBvkhbr5rjtmWKCPeAYpcwRAdq8B9hnBlMzJsH0KGxnitQ
CpRkO1/ygEGjtccYgKN9bH2ctWh397uKJgEGrdX4pRCthdRJYnvMWn/nDW8akgM/SiKA6nfEi1tP
sCX2CvHymjU52p7AEI159vFGqJyrr7DtYAh9Vstb5oY248aVdY0F3Jos4M3OfABnMosx2WXBK5Hd
mN8iOj4VhpQGx8pCCrT55/+qpC6wEjsTQDZ4H8Kvf0OOwPP9hxcs3DbDjXBPDjh6tKQOSxTDG2Yc
ee6/wh3/2ctGWuG1T+nTqNI6/LFIO3IiryQsLUrNQn1lSgpxDDf8K1/VqiLUMAd35pqSF7kePWFD
fBXyVmWd0nbAKccx7vXit3s+K7aMITip0DT9sZU8LrJ4248m4+I5OY7N4NwAv9m7Ezws8rv7146b
dKqtrvQ67u2jIUhUpc0nfWO93/qyUl1W8edMa4zN8Kky33vOfnvSObp2rXwFdpyX9LPk/AGdik/T
UGoKi/biFOc4gnjs3TYWId06oaHfajc31qGWSn377kPi/UDC05LCF0spM9TwI8SgXy+lGe26eq9v
RHqXH1tuALddsAC4eNgWdq2A1JtYpvkJXWfn8PF3rJPaozBCQLSAf1EAjrrJ4Km++hsGYmMEzn4V
AV/q0opHEb8/p5chUSbpnSWzVOiCd6sMGT/t+q+jrGvAq+IzXvP0awcWp7PLzsQJ+5WGLsRovqKC
BScJ5U1kZCG9J/RXKOcJ6THz2ufYa3N/qgkHesi0XNbc9oRLiXFPB+8C+Xp03UB1Ck4up1jkyI+l
v9v4bExs2ADR2hpgpNkANQWUyqeUjJ8hZpj/tSNRcv0FkxN1Zf7Gv4iUNovL+YPLFgh+dN9NQDgt
esJMvU9F8y96wypLxPZUFvZBHtXYXwa3hHXXw2zYjVQHwka+NxjIsUtgIEj2IEPKpKOszXdacrhD
Fr7RNUiUHrE7Oqz2O8wiWuj50lUiZFjtLFSzqZGVRlnlxewXW++sgdQcSUDpaY1J53vqamV5Rk4v
grqy/PNvWkcBqDjkN9RGKYjpBjyiJlRStcEJMKgVq0755+N47yGeI90pd0AyqcraSqTYqF+OypFY
ZUH7MrFO9ULzLNFiXB0SIsxfEAnR2kbA61DYMEO1XrZZKweSCglg6R8BMmSzPv9hWiZNIm2svJX9
uIH4V8QseZHic/G+/MpyBqERTQRfw48Agl0vr1WKQFSusPN/YH+/pOQX1P96LN5Ti5k04uvvd1bW
rGdLETnwu+MgwvG3zEdPQETvK+fbedGOQo504+ppYQ4tt8GhUsNlia4bMJhHNLhStbgZM7yhMvUB
nUKjzbaDSikPs3lKO3wyJCn2NQcbhmnU+MRXURhy9pY2wwOdoefgrAmttcXpM5DytwhkaWXGaSdz
Ukvs0RlrKyOUp3OWq1KqGc/KvolHWawU89CKXWc7rCZL1sodHT/YkhLMDSk3flsvoxfiX91US0C5
rxE4yT4mb5/XxVeDGHQrtrtz7F0fm6BNxGIYDXDrzwkFRBG6CsLE3wvtuEZ+7ITu1dih5phwqvSp
yEHa98FohBgLldAKCKmYBT6QlGPzLcS5ctMofmg0EINcdKlTNg7K9rAL94n5cLLmEWVs60JgZRyS
u5iBMVYjpWX5+OpQ1Op3LuxUuma1Am2xgtkFCDMmJ3gNOB6pnjP9xraDKty5x9Nqs2e4pzWuHixF
82KOVgjdlmOSnocwnFOk4IMIu82ZNAZ59OSemlTjH1NKHLqWUZ4wedqkNlb8mq/AVFSs3xeDCAPf
BY0fFFKCxZcxZkMcliotLyzaAbg88Tb08BR7Qn3y6rLl0e+GsFQmgsgk0UmOuEyLOZuTEUxdY94R
DrDOBuITXhtoWWKzIYombFOnIJ6XiZsLijELKrmJSP5VOvcidj7z6Z/VKT3mOkUeDBiitaZO/uJa
Ww4n6f0Wzb9GMT/T84mC3NgekuwRfXetxOyWJ9h4j+Fyxfz2p5b9wUdPOouGCvddpdEyOx/mRDlb
xJjBkjIOkbDQK7u5Z778iWm3s4Q/krqLqowa8ehM81jy3AqICNNagg27dCNNGr/nCp0Mho0GmV7E
hnPwyskE8MIySJ8aNKakdj45LWML4jX+X0sbPnSPPGsW0tCM0ICp28+oi6mn6UxsA5aCFDlIf9jB
uuLsTZ5C/eh+bATSx3XCbccLK10XCNBc4V0eaqQj01FEs0lBgTVGY1n6PX3VsN/Uhqd2t99V9sk1
6dAHCGmWIIV1uXwevs6/BA/JGZ2jPLq99r6wRnsZw/HQz2MTT6Pd9FgtykwXK/lB5+BCB2KsiAUr
6df04SgLbyoOnAGtmUkYHk4GluXRxB1XoebSaLGA30mkkN4KOML0Owd0l7cEk6s1RSFO6XNaYdMO
kM1oF1hu1FWLExnvYEg+Jo7PG7Czrw9YhT15HaXQZiOcyvG9XZUKdS8J2W3m1P6oW0TKoJpuhg4y
M5+lkCA/nTUPW2Fxr+5clrLLG1sWZ66spRnhyeEA1RF8YRdbTgtXMVl/tihjr9RxQo6BvEdilOZF
xewQ/67HaCE0xxsVCYDCXADAM5Magvhp4QlDQRo4CwGkuNRX/+2+uj1vPwuwYD7xUBgxcuJVYYVP
8MOhqwWij7LTRJxJ8nZy8k7r+gTSexYm/uHRu3Pwgj03cLhoSUb/NJHJw5IbN11SLe09k11SMgZn
0azxjQl+OYvK4hsbkYaRwkJnyK2gZ+6qJH/RhQHVwGXnxUT5WRtbcmBaGujsM0nf+K1VYPAdbHPX
7gsZjcBSlx5hDoIT7fhpkIIjFuMAWx9zEj2gGZ66vR1dew6eo93GcBvuacO8OHtfVJJ+Ov9j7Net
sMun50tG6cSifrwc9afAZTuOKsO7IzoTndP0Hf7Oqs5lTJPlm60qNFcmt5QbDhGjKQ0UN/R90I4U
a1/a9RX5dVQiom0WilzTinDVE8MKJe1fsNd/B+Sn4jLW+N0C7xlD+CRugyS4a8snlSX089/NVp2B
ygUDJPnwp2ZQ6BI9kJ58G9E8SDCo8PQutlGJg8yCy6law55tcPlp7KnpVGmzrWRfzr3/8aesceim
2j0pnDDX3SMsoiQoiNKo2TWh8KwyNnE1ysrU05rOw+0CIQfY9xfV7k6w7fG3Q7QbaLKcEJni1cRt
MtDJ9nyavoQHEtwKEzr+WgrPqy6YrOdApp9vEASDw6ra+lhCFKNORPKo4fgRL5krck/gBDpRIVAA
GnHBZnTfwl3MAuXYz2CMe5BUah08A/kvPQHLA9YVMg7G2TlUeiONu/oK8XfQClUDjkp5U9TcRoqK
p/1ImhWm9k1nihSyny+fOCzfD2ZmGlk31jWGiA80pVGBx6q2H6A67GqaQyO1AUJ9Dcp7VDU62fkd
k2UO4Po81EDTq/0132c5/HkyS44uizl49LD9LEtyRYQTWkXPe7To+/8k13rYlGdHdN7paRsWwVTc
qqcp2Txn5uUnv3IelHikxSghh7+LtHTpTf0zbM5TDlJEdsWuUfZVzCar4ISCSVkJRQ+sW7quTqd/
aWFNMV4poKvGTtmG04XapeEXBdXf5m5NsZUb7SshjcYRcAS3d32O61gsUtiINNQi88GWbA8y6Jg1
j0yuiFjC6oBReSDI1xDSRlLHDB1D1qRHcLL9KyEIq1ZMpuQUjKsXtmNQ0W5HZEZpLksSlPm/WyKA
vCXl5PC979zdbTgh8CCHyDNMvbJpxZ8ST9jXsPWyT8LuC3FpHgVtS+SiS31RFnxlZRFgj09yMANn
HZ6WG4r44LM48zdqU9c+FT5jb+1S+rUysKgb1ewzlIbEeVIyq1flfFO0cZzQmo4XThHbSXiUgErM
jwkYlWFIXDCrQszSS7vDzixz/1B7lxfPTuAoow+KJVPmkVQ8tvZKkTQbd0tzuZD88x5TeUbF/sw7
ix8dSp69UrXo0HoeqG7kyR7Zc3DkJDAlj/ISl7k4zR+lJXIzlzy5rHRwyN+LXz+JwJaIca0heaGz
V7MROMBk2kS/8/MJuFyYa9mtVGM8U+UU/dA7CrsNW2C1P9ObHciax1V4FEgv4YazaULdk5ksp8R6
HWPBLleNsFcPEWd/KceogL+F7/jtjQNpfpRrLS0JkK+MjJNOzGVGc4qufju2n+lPXivQu7/qmRMl
xYP7+Qir1y5ftJs2Zc6yTazjHDj1ZrBiO/4ZEByn2d2ThnMOxO+nv8f5BRHoX3iXbidCt/1yyrlo
rOHnHfu8kL7okH+MFW2++fcrrSclBt9qfqwUM5WZkst7ZZDghbM6vautD3D8WrpIypDqQNSoQPbm
pYIB7cl8vRXKeiTy+EWV7OKKevPBAJWPYclBrrffcV1lhotVKhS3RxC6Ig94Gq82M37ZC8zuAVhC
6xQGTEbMHGj7sYpm+TpCOIRqULc0YEYfsWpLnH3o4Y1h64SPbIeIQG7Kz51rfxlghYSp87G7LhLg
LUBO0M/3EUOUWrHbbOFp2HKnFv2kGnGCBbUIzikxQQjAfab7XDcJVczbpk6JnYSVKIdDPCOvcLL5
QEKy00CvKcrk0VOisnQHTYbRnmhcoB1p0foPBu/nDtMm6HLx6ujhBOaXnFVQo3CuShZGXedxpnV9
jh6uTtEpntzFzy8jG3UO5KR08hA8KDI2YBz9+3az6vFM4E5OvanlWrpFaHKijXK9vmU1+q/W0U1F
F4J0W8BVCDrxA/C5i2iGp/jR//spu/nAxzdq1P0aDT5lPHJjqrD+8EHMtNx1QhILXY11jnCKnM7m
PeRwbbCK2NzCT8C9pVo6MZaQQE04t63cc9GqJ/ul3EYVN8QzX7P4hQ2DmsMsLz4S+l9iJ49mTqtU
T4iqDrdeLQEciAuk2NptmursG0bZxUEnM91XKMfxFw6o7U/tg9xJ7yP0KhM8ENibbgoJBtXMnVc0
/jgWG1h7Dx+VL45AbQyx5wEucX/TB1b1AnfESZv06/etegSqnUxlPE8yo2gBH8Igr+KAE1f5a7qx
B6dUe86DJjQjsn1IQyUze9m9FtuBh57M8ybC/fA42j42GmZFAj+LuD8vcII2SC/qdCgGDYH5HFdB
capaM8gmp57R8JZNlq8SMM3zDGnkDGF2OeM2dEv8Ibv6liV0RNiWIEWRJ14KZAfF/DtHKx9uCtCO
NfAk+K9o4CyI8FomoIPaM3TYzPYKjWQjIMFS1SiVHKfLNGQsIENt7qzmzm6qwVHNw2B6bRLOgW1m
iqb+Yl6m9EU8ybYb2C7lBF1rFCtp1OCLogK1sLzxkCa6rETxdDrf6xG2tRpSNVH765DRsHzRuB3s
q7yiiw2YfjUdxnCUnU8552N35i3TLP7RJ6r8Yzglbbuxx8VurEVdI41+rIKhfreFcvjhqEHPfcRJ
ANAllit8mOxBr2l5ui8q8NmAmob48vbgRpbGEqFlQ1RKkC8gHmI1uS0V1KXqXijhdLjdTkK8lGMH
HO1f9eFX51mxZx+4eOvp1rLl+wLn6dBcyJj/iRxDf/kcZTV2rZB8FT+Bc1xw+YwRINIrZ2r1Oe2T
SjAk0CoBSCLbTINb464AFkhJBFHSlLVnnjVcW++VES2r3a+7XdhwdtKxfgOz3cyKgm9yYmQH1yOg
r0sSTg2TaEOaYeYumsvcIvaS/sF4OvyzlrqP4B0Bl80k3+sUEvPKGhH681V5RKuY20L8JSC57+Bt
auErj4JBM8+ObCs4gV5W4TIVvXbJbTnViVAE8F/6G0V/Wi+/c0IjQGc3T6hu7gK+tvu5P026XxXr
IoLP4C/x7y16KUDxjgHlImOVZg/D6MI1nZ3yqxt399RtE3P8PTxeQPFFq19Uoeo6mGvBWZ8xjyg+
l5PbdyFY+emTaPFU+FUqZpwOY/Sx82s8uWQ+AK+b7ooWQVJVyAFd/xCLc00Yw+DIyvgASz1jyv2T
ezNX6Oy/AYG0gxrutr626AaaB3yjm49K9sdp7RNL4cr1/5OHBttTWSjwwqxEBvcWDYAYBAF06XwZ
j5TvH4MkbQBNdaYQ4n05vnpkaZq7lSY8jryZY0YjZqqlZjtFzuI/2jEP8mf3LMDXa40YePBTW3sN
OzCt+JXjhKzlpz8FS/vqLeysa4gn941ajxAtyM86F3Y1JF2l0a73XK97SA7T+5HXc+Jix88Q1pbH
MjSysfhoSe3sFxTADYOGDIPSEyOwkCIp7nSyXj5aXii1Dcxs3h/HekdiyDL4Y/XIGyvZMUBPr7Q1
ZOrGfG0kCR9jOEHZP60orREPKih1qxqaMNv20Aqs7wn4L4xy50mbZaVoSM33V7iV+kKSwsVcseKJ
tPy3msg7SRcj0XTOez5lMpIAfUTONJy0utRkSRyoA+mzdjzACtCnYh+i8qr3jJRVYnl03jwLzvM2
M/koPOsvBx8efw7Q2QpDCa47EvhrFoGH93RcoJ+OiFVlvm5hLMeKwj4QjnoPzKx8yzBfCuOtjbpK
dCzHbIGaGS0kWKDunUSQdiCa/uUSXcQvy8+gnhuSowCloSaPedsrPqbnZvw+QQaslq6EFjQqzEq9
K2BooGH21mCzhxgoV4h4UItxhYMpIEBOMVjEF7lGQtK+aoDwi2aRUD2/tJv6HJ+g4c70PvG9zd0i
piuaba5OXpRyDRPFP1JVDZ8UL2s9oTpsUAjG9M1fongItD2FoTMTu9HNMuTqV0pQ/+tP/aZ3NIN1
+8LG3QIG2MEJZ9gpsI3qnlgWCbtAtozkWRX1rYgbpGlM5lnDUCyLHmXgTojGEr0wIj2fsXp1+rSM
YRBtXiGzvu7MA4nR6lIMA7oCjPvHXKr4JLPhODlsw2b6iXH4tDSgL0j79Gz0TLXu/VnWQqB1kocn
lc66Xx9a0ZIFoqxoC8aRivEMilAdmvgxTCDXA+FJ99D4pFHk/xnJYYTWbqStZ8r0aBGnezg0+a02
Sdh+PjMmlhKU5EH+XK+rDQM089A+TlnpiWlbECKAPOFRvZJ/L50oeIWZLnwvrCPKYFgl8EHhYMHn
niOrjCBPzAjlwY6NK9nRzRAOeXR3Xn+m1mqCX9TpZOKNzNlCxb3Swtl+FRvQQjY9GEoDcdySk9Ti
2B9btKjz98KnB/o8MmTmeSLKaITxt2ehPRWvd3wymIpRNtaVrVT/rXlpFelVjaDCaOQYqaUTZmmT
7nmlyBnmkcdqjsgJ9kt1I7hO0Cre2mnd4ceTMYtwKSyWSwhXop1h/cMH+dpilsKraRcVKlbsbmNB
U9alSkyEfjnWp81aEbUGUktYSGnVAIXGD6E77qpYX8SjCg1gTs4iPktZvKE9NUVSMlyk52GW9eL8
85xAFrvuWlHiG2MNNySENDraTgaouA2CCqteNYSVJbLkEEmbypAMnNRsXUtCxJpobO2qYVIW2Ky8
zXd39kiBVvUbJHamxUpm6UtAQUOB7gRC9ivUROGOUY0J0Lri40IHEbz2ppwI2Bn9OxHekkD2+v6v
gsbzY8Duxrxz1DHXdznlw0QyulZ8m8SrIOdj6ZpKOMfccfHp2I5s/zlEHHQoOXLpKzVY6b2m3Ga/
ZpmfYGht71f98MPk/PFMJudeK6TQVu8FlL7w+TWCKEPsTAFeok3SI5gAw3mFDa6JukOnzdUshsK2
zaOpQafsmHmqH6puCKrX6gxR4c174LHxoP7BLuFGfhk8JqNh93WjRIryhfATDPu1AdSK3YOMbwvj
4mgl++QN1VMObXaEPyfrRt6oxEmaPR+sIp8J/Tsh414Wma6yD1wt7d7nomwcNaqbRPkiz/ysXEm5
s0Kl2K0UgYxd/BEqQKFdbWTXthX+kvlp2jzgQRcORcNT60FPCmSV0d4FD9Di1S4uYBv5HUunOsiM
r+o5hCKt0bGy7zwyvaXe2EbQ0s5id9XDjlT8NaikKW5ESB/HJWENovpsntoxOy+/oHVu97NYBBfx
te/86vrmPPaUwZNHiuqj8Tt7vSIan06f6uYSp+ji8B22pmtAFZFgWaixS3d+DXfZLm+TntwalBJs
vaL2w/MjQVwhnYyY9QxpJhkX1Pe5Y5+5/Dms6+THXcYas9GYlDeMFVXQmr3HsHILdY7RCXLnh9nb
k3vsUJgkGul1Mkpoo4YSFpt1qFlp/VTDeNq1UswfCX4VgF8/RrL+OBVDGXn3jW4uLwohiYqAAcxb
x5xveExMvuiaE80Abesl1nPl9g0+EY+E8k4SHa8NHPZ3/2TVb2hjUR3lfXjvGVzj43sS47BTH4A/
pQFTKEwohh4rqcHaHiY9Io0wyaxjlSG99KSioeH/sNdbLpr3YqpBAp93NJxW/E30+EMsaMNddIjN
bSK0f254NdbOe/3qvqr2LpQOKADdanidYtEg8MQPLZu1J3lOTLoE0xtKmFsS4pWcUN1CG5T2uCz/
raHMM+FFFDKYiVL4esBSdCQ+6JDTAK1I+Wmt+cNnobFvPP3MacPuCYQ5wgg3De9cCfLtOxJrkK6M
xNkEIKiSZjxtGzRIasydZLepZdlLgiSay6WvycMbDpWkJfxN7LcWP3GFKrLfbhidQdHxVhJHomA/
5HGDZFrU2dZUlFqsnKbTYG0h7oheBoCnHJxOJZ9vbi7nMDNzrVqiRxLDujQ9j2rS9zOpnnjzKyTz
nVvYONb04W44LyV+JmI+pyZx21VAoEayuQB6Z0CRIQmrcE1uHgz9u7vBIBAoV2tozHFzcqmGG6U/
ivXotHGlBwpA1B6XNdjIy61uWetOfZPXjcFCU9fUV7Ydqwwl5wx9b+qJdy4uOYuYYF20Uxjpykif
+BsXzpTtoOyOe9CLxrfnBgO6HSHgwQ16P/qwWlFzIakSsZETGIvEnYAqoxrA13/FO6D4j0T72lT2
WZgL4rc4ByQ+qe9v5DIaFNggwy3ffrcBwrbTqG0EshXtVWSNrJQHkYcMsSVjzUsS7mhTNJX646mL
P3C0hr5SUHzlU6ey/mqpC/ZsC7q5l7AFNpJFGiFG9sCW5RUM6RD9bK1OCRtoQxiOsIMHP6C8Vu90
6iK1dlqDdVB9FAnL5c1cXz1drPEWNdrP9imwLX/0DqcLvxd/m6bHcTY+Ok+IRc+9TAulLBTwaWrz
+a5sZwWxOF6oMDBtgXgnhFWENvQQG1cHR/oxcN2Nzas8/qGbP/NLHaJKtkEBW8Qp9z1Lee3gWgkm
6CxnbBTAv8bDcs4D1yC78Rq/hXrIIUwWcLdpmgdmz0CyBmtWTpyt8+pHkKFQQOl7dll59+D4aFDD
AAhJm3/p8qa8Tii4PR1DsNKNZpULyW5d7RRqajdEtlQnEKmxREhVJ7zYAqk2UG3DaZiqu/seL8Dd
iIpzAgfe1lhhq4HDncp9EPSCPyJX0HqLJkkyCAssRnSYbNa2TFj/ANiMaM0VhBPiTVUqRiHexoBZ
gDKDwELXows8ke9MhLQ9FpmKklypXwXPtoBw61RJb8aGiu4aTAl0psGbk5KUvGg509mzM+Mo2eac
592vFM6YJOiVg5cU1flr8QTvO+ivmW3AvwAZmOzSNJpHee6mzPJS3VEOIJqiBKJ+1Va3STJRQnQr
dDKAdsdAMT1LaXW3lOhU0iYgcbOWIxmZBOoF+kbdFAC14fQz5V9eX8NLl8fV7WVPRckZz+LBKbJp
n/TGT9HT0hnxWtScieiSsH5aPmRf0f/4IYttjA7VgFHlsgdSohfcEcGKv6yGVH153CtGslLI50hp
16E/41XEHmbhpH7Nugta365pV9GYsJ9jUmnVTNjG9w8gxckUX+N9vRjeS4iU+VQV7q2qO0T+0kp0
pwFOUpw0iRmmcsjn+K92VOz7z9oOkl/0InVoQHVPEPfdBglGgWb/QxFCBsRJC8qqWnxNpRPiFSMM
1j9J9aJwTIg3+tfB6bymGp/T7splE/ei7LUrj5j8rbvHEEp0k1+Y3VLlCIb0k3kXjmH7Az9Hw2aw
BilpG1PA45p/9U6I2hYwAAuqbIwkWeEzZKTmY9Vos5UdDLbN8eh9KluqPLVA71Y7XCuvC7vdjnCc
O+axbJFdyByvYb2Y1m6mSys+aHY4aKPCFpDbFuiJbPYPu6AY8hwSNViLDWbtyzMHVuBbdTgoHtGz
3swDjHVJvtjiiDJdruhvfFOabRq25YSl+s5V2iMQ0rNWQ94DKRlJIPoWWzh5iJdM0vPG1QFavDuS
Z3Z9JjCpEp9aAgecDoyUGYOpp1XADRAXurM6L2sKz2SCKAZL8pd4UhM2yYjdi1UXXvsyr29LOz8B
d1BGnEJy+c1LW6yblNE9qtP2yG75By7NLmFzH46y1R3EmOIZ7xFaoJCIE7kpIjIRtUqI3AHx25hI
/bvM5CrdNZw+Nl6EpEYrB33EcpFPBOwegRelzwz84Ow75vvTExjBmo9d4TQlmCwhzrTCVmzmMZm1
kjkemRY4I+0xRlTUxDRYzKvEPqjmTekIEV+3aj+3gXpdSAz9UocBNDNQxnqDWIHNwKsEiTUUcz3Q
YyhLXzb5BLMohVo4sI8LKcnm5YMDqk5uxnyqed5GeZl0LQiFe6GctUvpyhY8JWwEMBmOCkpmF+rw
8+SLIF63+soe2zoPTpf6ozlwznbwY7EBCIV0lUFkyNzTlJSKzoHIX3idVWKMKD3xxoUc37OrRIoE
tHTt7UEjfZ7Q1U++ap+E3RbaFfGfzRVje+em75ceJASMDnZO6bNLJ0LkxHrFzhTACXvV9s7K5QXq
LHPJgqfvVOohLF67nEGfsPgW6V6S2HPyt7cwVtgxcIr8gvw2oT/w5JST64Ca3teqHERY60l1n9R/
K0UNL2zTaYIotISg6P0UJq7fpwl7MIqqqLUMQ3jZwx+/EvlWy3FL5mkCq+QbKeRHvGMYgifQzrBL
kankE1eC3vy1rtToTqWoUG8D2FQj9Gne3s0R0IXq2OwNhLEXwSNbeFJTrViIrDg=
`protect end_protected
