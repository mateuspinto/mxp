��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���:��1.f��k(���zp��'��FL���s���n}ŝl�+6<xޱ�t(�  ��۸э�#��Q���/��Q�}AlM���������-$4�߂�Xpx�����RԷ��p���r8I^͹~��F�C)�bC����R���S;~��׶�q��A�ڋ��؁,٦��:���T��$�Wm���Ջ�m	������<@욉+.�k!7��?jv9���xF�TY�)�M��(����i�2��;V���B~����ߨ����C�����^�߿&�<
���ײ��w���E ��Ӄ�q5=c��`��ڧ�ޘ���aO�%�ӽwC�-��gZ���)���-�Z�~��2e���!A��[�foI �!y���=�s��1����}��ַB�>�
N�D-�����SƗ?����@Fsa�b��#m�fTV4��phix�
>OH�H^ᾅ��3\�,)Jm���Q��`�È e��!��dM�u��D�#aֵ���>~2*D���)w��w7�_�U�`�!T?�+�lĳ߿ۥ����R��w��5�����^�.� ���L�N!��k/U�C��+��Y�8U�L���Ng�@�މ&�r}Z�ޛ��'� ���F�U���I�jq�;2i���5G��/n�]$ �nʮ�אTy����tPl�Q$b7R��yJk`�SO����-}�e.)v8��/�l�O�z�4�SM)�+�]�4#^��A���>�T�M�nS�ݒv߾E�b�c�\�膇�Yhsy��P4U�!s.�~��՚�hB�2�dN�����L���O�0<��
T�C�[p�����a�[?
��x��x�F+a���yR`Y�/�"S�;��,��bTu�@~��E!׺�G�s-��w)�qhW�����)\��<�0��h��
�e9P�P�;	C��()G�#�����\-�n )8�����\$6�r�5��i1��ms�y����s��AC�(�X,"{��r���[���2�|�W�@���)�F9�J�T\[����iV输<r|=��G\Q}�ۦ'8}������X���K��>u�j��?۱|�D}x=����jS�&�t�R�D0��D������eUX	ōS!
tB���B��t=_	a��Ke�e���*���ٳ��q��ㅲ�_Z��F�a���U`�W��:�gL�y�M��:�NL��n�j�/�p��f�wU&��H ^1��S�g��xGY��K�����7��	�|�&9�)���Cc��Qȷ��6�{��~�=����Ϧܓ?�;A��[��"����7�h���P�D�;�j��`Á{���&�i�Pcm0H�Kϐ���ÙՖ��3�'o=��Ex�^莂�˲lu<�|~`�A�?SL�H��v��q�88�)���D��'���� /�,S��+��5�^Lݨ�oI��'���u3�8�����p>���r3nG�9��HwNh�#��*8	b|�l)�(�^�p�@�{�}>���E� y��H��N>[1-ڸ�:�v=\�-������d�4���N���<�@���gP�f�\����ݔ�R9RG�S ��N���y�8)C�.����x��Mȡ�[�u�dKR�)i_�g���JL!�\����b98FKߜ�ܩ?b�i[�c.����V,,��t!����f�y�b���0/"2�8b�����	G�����	�H���X&ut2�����ڣ��BmL��ƪG�����T��O7Vuֵ���) g�2���'�W:���4H���oT���)՝/��@+�<{��\|c,B�������㰸c�ϋ����1���Ř����s+��"�\ Ɋ<A|$U>5=l�m���zX�}˅-Hd^���R��r�\2���~�N��F�,P����UhXϽ2���r��М+�
����#j�P��p����^�M�2�^e
�'Hh��pM���}7�'~�	�H�B��CiG��\|�aϿ���'��,�~�-t߰���|��ʯ�͏|��DP`V}Ou���#�B�vP�Y!�Z^�[_��w2|�s�J�R,v�з����G'zw��<��L,z5ӧJv�i�#)�مY�O6�Q�
�L��N�k:���	�.CփAMSvk������2'q%��1ߑ��H��a]U���
J]}�]��?3���'�-9�#6hN�J�����B'��Du���p��L�;���kQ��r�y�
�!F/�U���gr����\ʱ�3/��r�[6�h�J&���?*�ݞ��=�v�2���,#�&���yW(��m�`�J+o����H��Ju��b�3�|�D�߼
�W�v�(.y�Q�KTau&le8f���KH��=��b� �0���Ѹ����]X��S+c�@BPe	6[GkM%���6�f�N>*OE�2���Ry�5�}@n�Gt�WS'(Ǳ'\�ђ�ho=�Ԯ��>3�;{��LGa�tm��8��O���6�����Cf�F\�%���߫ː���60���u��	BQ��c�)ˊCA� Zp~�2	g6�Ḱk�T["����I産%���굎��̢��/�!��8,eY���D���ǲ�Tj�&�L�碧"��q3������I��p��W,gM�3��7���%;2�@�[˚�_��T��ݹT�8�6�+)Ba�#+�'X����^�%$<�I� ._L6e�B�g�����>"�nY;��Q�L����U�����<��z�`�F��A��x����EB Y�@���S�c�%2�h�qy���qEv�"4�|7�׭b�Ð~�Z�.���Hρv/%�(�@Ӗ	c+jϜLSui᧋?,㩸o�a!���ĺ�5�۱bp�����8>��Z5p�i��u�����w�O�Q���(��r]�������t�Hć��	�aYm޲����^
���,l�l]	V�}�5�>��2�F��Ģ�����lj�瀬jU�9��#�,�( �7�ZPg�An֮���ojS�Q}��w'!N'Gᣀ�f#��
�2��_[!�9�J'�WY�$h41��W������j.d8^e��h��F�����p�S�[����ղ8:;�&9�'S?s���@��i\��RK,����?�%�t�p8�_�n�
@)��y|�il
�R�vMc��� 0!I�N�;,!����g��E����d8T��Oy�� y2*�u�eE��I<��5����Gfzn�>�̻'`�3�S��^r��=W�\Q\3M �e�[��z��낃�gY��s�o��?_���HJ�����U����3��Q�$�^QXea;��.Q8\1�}�؉�ŝKw��\l�w�"-[׍�_+�ô��j}>P����J���u�4�ǔ��Jp]�4�Gٽr��q�qJ��|�M��m�;���o;YCL(%��kKXJ}���Z�M��32{���_�j�b��בc@��Az|NO�M�@?�W�K��SK��x�2�Zk��I��UY&�x��ۏ����-��Nׇ�
�-�O�V���bѥ������>�H�����K��
���lU���p������f��#�1��I2��t��e���6s$�so����.�y�^d6�z,z�8��#�3�z���Ş@�N��*�S�dg�p[�c�1�L�+��f74�Ė��ofk"R���æ��jk$���,s�����\�H�_Mȅ������ ��
5�據%@��1;�U�kdh�ԗC<6K��B��q��%{�,���t��m�L�*H�&F�Mc�%Y�E��"�yi�-�L��l�reN�;���g~i�������"��Q�B��r�z=&qA�B��Su��P��}^��ڍmN ���OfeV�p:�վ��7��O��ߚu;.�Wt��F�"��*̺�O"�2�O-�#ۈ��a�ˢv�=�� �8v}��K��%f�	`�������:'�f�7&���V3-b�����ꯥsn�K�d�pZD�E:����{�gV�Jntz�F3h��U�n�Ъi�`��VL��)s���������i�-k����߄�J�#�Aȧ�8�o��>�F��z�z^��W����\��	���5�,H������rGA��'�L�.��+�7��L��ZבPn����2�be��O�~�ű/m�L`��������A�䏇�G�^߄ʦ8Hq���e��J��Ex7pp2Ỡ�w��Tm="�	US�<Oɜ�Q��^qdsV�CEjy�5t@#ѕԖ!u4/��R|E]��3��._�����Ǚ~�G =��hiF6x+�ݚoԭ�i���V���NG��V8�C 5^$^^ `����p>Z��ո:���#C%ԋ(�WM51;F]�|׬^�d���f��	A=��f}^������A��_�=N�l��wh����5q�#��O�BQ-%�����]vH}�V��3���Hfk$?ұ��C���X4;�lE�>�omA�����So6���
��%`d�f�M�����"�˦�ʳ�hv�K�l�s �jLܶ��A&�'�RM h]fa�<�"fЄQۍaEc�*��>a������Y�� ]}x�-�O��D�x��o�'#TA��qR7DO~���E��S�9u�7;���g�E�G�㳛2Uꊼm���Efv��~ڤ:����t)g�٪~�]�[aA��YT��ΊK���T��_�{�mу���w�M��s�_�w#(/��D����V����jXxM-i@�R<4��p��?��}�2�Ū���U���!?3�|L�J��ɝ8H"�̞�D�N��*��Vs�1�>6>����L�u��j����xܙWɔ�ӑ9"2�\70�Z0h�*�t0�@=NEڊ��#hNc����:��IP%C����@���=ic��Ts�8�Ӧ�D�l�
��(�=�=��S6��������%?X�Xq�)��s���Wc�셿��>��kg`	�[��9�5?8�OP3���M�l�<�ciaO��u?$n,�);��?ױ������"����ն	�/OG(iw�t�˚��M�L'	���TK��|c����v@�����یWwE��t�Qf�	����*r�\�S�o[x����()�,$�Ɏ'�$T���6͌I�����TR��,5-��$ƀ�����(f�[�µ�׭��X@Ck�-G;\��,ǚ�-k� ���|ۏ'c��I� L�6�dhE�U9`+"Oǧ���e���F(h9�$����d�Ƀ&�E[a��V���O��ZE�%�dQ�N���Vb�J��s$����b8�/-������y0�y�0d�Z�/���^�o�Ⱦwq讑u||nS��T�z������Twz���M���S��>Ñ~��!�<C
��5_J1�8���G>������,�2}��/-/T������6|�+(��`n_ش+�AB��#U�S�S�/'-�O:��c�W'P(�+3Á��ͣ�/��J�����p�%��o�\6��?�S����5�y[���q �����o���C�W�$��Wě1S�+lʁKɞ@O��;�n��KMj�@(��c蓣{0T]b���{g�4��ei�ê(Y*(K0wi�B���fS��4��:/ŀDԷ�s�X�n ��O��-��{o�ko����� Y��pOF��Y�2J��F��f����4 &N�>�Ƙ�_#���AǠZ�j�q$���S2����>�e�@w�ڔC�D��)�uK�:�'���2���z�oS�#�
�=i3�ҋ����c;��h��b//ڢ
����޾WB�]����
�v����z	w�#�Ë]�!�oIݣqSm)���xQ}褀�?{S��@M�����x�����S�T_�X�~E�XuZR��n_4��Q���bI��s�<>�x
/L/�BV��S`���(�5�/�h�{<ArK����z��7��G�'��%�\��bv~)u
ֲ�O��ߑ%�t�|��Ω�/�ػe�;V�7pg�3��*�tf�ٟO\jU�����bJ�G����k�t6����,�Y~H��	QZS���o'n��]W��K;Ť�U��෸�!�o���X]F=	�-v�>���T�&���2s�g�g$�xh+H[��'�u�-�ε��D��b�ؘ	�ՊH�.�+M�1(�d*t���J�#��u����4�q�?W��s�������,Wׅ�ˑse6�C�8�u�d �����������S>]��阌�(T�X�����QTi7��A@��qaPl|�!��IX�M���㬚�P�f�6�yA���������ǥ�߷�/c�A���ş(�#�(���l;8\Ww�n�G%�dg��m�i�^>�0��j
:�|iN��?�8Pvi׵�mD�ڦsc��H\m##�J��� eaB(:��X��v\��8����[f�� ���D�Bq���]����~%U�#A�Ue��A����3�Ð/��*UI��7���u���F�+y�d�,�a3]�gWӶ렒��Ú5����Pz�
�ƪ��+�� ۣ0=�8ޑ��pI=j���r��\gӮ���L�Κo�h͆,`$�64��|�g�e�����FR��~vi���c��=|+\�^y#�����멻��׉z�8E���`)G.R��2�,�﬇$@`���Qɰ���Q�"C^!�ͳ��YCp�v����-��#�*zx�j��y�	y�>9�N�OĈ-�T��)�g�l4�b���	oCg�D��f�F��S�YGK�߂��~�;�K-b_t���e��>��R �������+7T��0l)�X�{������pDlC����
��".����~"�Ͼ�M�s���a�����8�s��:x��u�е��9�>I����0L�6�s�/Y*f�؟�f���6PIXEW�+�n�ky��剈o=�~�"х���xb�e���A(s�~�:�N��[��bMeJ8~٠�Ű�.�6�jt�ºΗ��&�0�_E���mXZb�J��e/G��|�s$t�.�ZlϹE���������#gK�k9)����PU�6I�M��8͝a:��!��P��2(@|wB1��Y�U؏z�w�9�e+��C=��a��`b���O����ga�?���G=�F+k�ކ`������k&2�^�V�\�G$�Mؗ�2+d�U��/{8��A�ag��}�L�1P�*�k5��aM�A�w�����'T�'F
���i(Evn�eC��J�#H#=XWt�s���f��B*ǈ��֙GόA\��d�"k�"��v(
��LF �~xv|�IK/��(���$t���a P�	@�)L�/*SqL�I�/I`�x9�WM�{";��SU���(�3J�j|\��i��|��%��R��t�!��
���(]��܁d�}��F���=��x�ɭ²��n����#�To�����>Aݛ��z���Æ�p�Yk�������K����^"�������0o�Im�������^����RV;�����n�,���B8��jl������������~H�$��#"�v�{���ܶg�:���z���C?z�:[_�CR����Ga\Y=�}�p���a���8���_;��-�K"��c�����&����gL�R?3��e͕��`�}�4���X��N��Db/ ��xQ+Q&C�K�3/�nw���/��1'��Kw�<~����m7������0#�9�v,���?��D���=�~TY3]	�6�a�F��Ccr`��H�4�G�f���d�Aı��y�1��9���{���Q��0i"�@�:Utz?�m3L��s�k�����~�&���F ��f�g1�KQ���+
%B4YH ��b=)�Q��L,&I�O�~��y�X���8�(��j�M�q�Ȧ�Y`ϡ��/�;v��'��>R�CL��p���I�z2����#�~:^�r�W-hY7vJ(�tUW��P|�4��P�-� z�4S�bT�wsE�����A��w��ł�����7��փ�ڹ���]����(x�Bb�s��i�:��M��R'���7Ȝ���V�s�̒�saЎѬ��:	fL����	�̒�F��2�[Z�&;Z�qdx�q*ſ��}�|�(�q��2m��6��Ehb?������Ԥ���7
�c�O�ҊC��Z=��$r霐���@�i�|�O�rr��v/i�d$嗦�,�6!�ԣS*TX�%FC�+!*P�%��j�O�����	s[%���?����1��}�X�_e%kl7H`��B"��j^�Ǡ�K�6����<sӺ	*5j�ҏ�]-P����)��uT��oz)/�݅7B�=f�d�|��9�R������ύH�Z�f��līh��l �@��y���)_� ��(p��~Vz��f��}���hi�R�;'��**�5�.�^.�o���R�-O�����_���r�w���Q^ѩ�d1fX&�Al��y5�Ƨx��\���!$�B[�e�]n�ukW+hο���

�]?�F{sR&��w�R쀈9^� ���x���X��]A*�^z��ϴ[���o�b��κn��J��nt��[]��N��n�mn=2���3CK�{��Mgm�@�g	u/��i� l��9	x��v����ꐛk҂
-�o�t����2��[���=�ݺ8�ԭh�t��hz���%����k�����I��SՏJ�U��dY]�MX�� P� �m�׹�cu�Uu��\Y�E��1S"(FZ�U��S���C��� �f�������������Н��&���� ���>��=�8��@�����x`ѩ&��,�e�=A��(~��s8�X��o�2�����-��j��(�WI�k)��c�U��J�h�Hf�=���?����lc�`>c���?��}x�Ȝh}�����Ì#����X`}W�<C�MS�]�����ă��7�lZ+�К��B���A]��	���c��KP�z�( ;{hQv^�3
�^P���F( ��d�wg:��(f,M�|�dLW�o�R�e�S�D��q"��^�`Ճg5BT&�� �5}�-���ty0�ޒ\T���q[���RV��2s �# ^9�%mv�������bo�Szgst
�%p�U;Ap`���I��`	���s<���`�L�Ȯ�V���Q�s����eG:[ٌ��;�"����Ƽg�I���l��S�
K�ia�+J+SJ�k���2)��M�{�g�Ibȝƕ�QZ�o̝��Կ��V?m���s��?C�{9q�_�/Ҩ^u�� 7�!�gݞ�Ҷ�mq���G������=^H�`�k��Ӑ�.��su8�Q<��#"Q��U�^��*Q?
�9/���߄Z5��4 �ᮡ�P���:�/���c���A4�������DS5J.=H`"~�\���b�:77�vE����:��#�I�a)�����*u\�?��H���P1/�VC����1���+��b�����R�p��N�n�b����M�~heP)�����.G_�<�KJ�%ᯖ��\�5����r�8KV���M[���'��)_
	K�����a�Vb��)��
�*��rn�IYq�:�.���ͣNF���H��fUT䛜 �u)��.ܞǐ���%?�Y�j�s��'��k��"�(׻����>���G�������x�����E�B����4�>������b�d��r���G���b�:p��F8��Ty�_�`�+�H�����20'�C�TANz��d�H�C^2`̐wA�G��̈́H Mu�zƄ�������NEC9��:���A������>�ò�eK�lhLX^L���v�}���ES�>��b?���#�'�k������
��r��]�����&�������,�G:$c+Է��6.Cٙo��Vx)�8���mw�}�=�zi���L�_'~�����cy��:S�/ag�;����G��׈�/4q�3��<�ݹt�QA����8���~K>uZV#�S9��@���,C��!�x ��pH�l�8R�DV�6�B�*#� y�A�9��!�$�zQV d�θ=�F��D�b�0���x�I��
�QjM�K����(ޱ�(�������ΓQ�>C/��������a�XА��faR�����GQ7Okg�Oakױrڊ�h�G�m���A<�>���G�-��=K��<Fw�s~/���@�53e��W��3N�)zڝ*'�ώȠk	�!��Mwr�2�	Q7h��h�d�ȣ��e�y��Q���_	����w�bK�HDf�MJ9��%��7(���K�E_,�6l!Х����S�{c��zm��chF7	���]1�'��d�L����JZ㊬�B?G�k6θ�ؙ{M�������]H��G�Sk4!��/��y�k�Kb1��FAs��5+��h��o�����6Nl��Ҧ\�N� k}���hE
��0qGw��cW`�9�.�h���n�ql��f]0�����ޱ6`z�Qϲ/]C*��*a�-Q�W���0#aM���!g�{�?�Sаk+�p%�3;C�|D)X��:v�8��WK)R�A��e;ae�h�����biA�c�����=�2+����B1�_��rBX��ͳ�߀n����Dk�"X��,Z�pfV,�1�5�k�;����B�-
��΍�D�<�p:t#���֗��8�M������̡CeT?�9�xO�Tw���hV~	��~1.q �=s�d�;Yh����VU-��r�����C/㐜�Wx~O>r���Hx̤����o(� ǝ��m {J;�]Q��!���Zf5�4w���~��1�y�M������׍6�!����.��H�K�p;'�����	<_v9�&q#z��n�W�{���l�~�SL�K6%
?\��.(�<�_;@�j$e��a\���vo܈q������t�9@��x�&#�WUꞤ֦��[����Κwn��3ҷT5�f!�{�Ԋ��"v4(u�U҂d���eq��E�s���'o��o}7��ì�J
�n��1��F9�پ���t�[I���P83�]9�Ӟ$�v@�J�9�bMl��*������ҽZ����b�l|�p����O)���O�������eL�e�A !��%,^�_D�%���d ��q�WWig*t���r�G��dUv�f�y���|~��6�twk�Q��˻�؂%�:))��k1(�Qh�Eh�%����`���3� ���1ݣ"��+�w�,�r��HtX��%M�^��u����5B�{���z�jx�؇C����S�>�EG%���`w�ґ?F2G�W�CPD>\T���y�B�l��6�"fr�M�1o1(��wʁ�T�&�t�^�"%0!�I�NS9P|������i����-��A�l��R�Z<��"���{��>j�xb=�:�.��Ί��@��ze���i��P[��U�;Qؙ��r5�5�[U��0U�����B�؆� d�L�dh�X � =�UX��:����J����䫘�rl
"�5�������"**�F%E*;�e��FP�������b
b��?���H����@�'(.7��š��>�X�܅Mm���!$V���W%�ΐ����?�Ģ��AT`�G��3]� ����`nJx���9�&�!��=�=8eπQBU�ϚZ$lx-ֵ���D�aX��!��.c�B�:�������M��E�*�GJ_!����2U�@'�г� ����2��8B!�.�|`�͒�[���p	���FK0/9�H�<��4t��ͼ{|�B;.�+������o����E��A2a,��M�f��J�s�����y����G:#[�8����*��玀ٕ WА7K�جe,毘Ó���yShU"�Ɠ�
�a�+��U���/�G�z]߄+��h_l"��ZM����B��&'�j�	��>>6�z�PO�J����@.|K�$���h����P��6��u�dRo�
�ܣv�f�wz�p�����X�|�^�댢�y9?<�jC����F��kR�l���HYy�0%�b�%wq��K�YQ���1��H:,�P��E�Y�x?Z�Ru�<�߂F�$^���]8Zv�ݗ��y����L���z}��i�A��+�96�����0%�"�m=�a��im9�uj��N�9�N�h~��,Ƶ��(|/���u�X�&n���DF�,1/�z��b��*ue103����;$��ף$�"-W�d&w9@��C����Y� e���@o�Bk���C�����0�>�>8���}m+��
g*q)��B���
D��;%�z7*��vGL���?���ڟ��;��2�9�V�9�x4vqF2��\lO[��J[�~p���Ӷ,�kbT�`�~����3�	b���	AQh����ޡ�����??#<����"{�=n[�Z8�hYϖ��Ȩ��6zLD0�\��ՄLB��y�#�	ފ|su���`:�_�^�!|lӹ�mQ�H=U��؝��y��,ʶu�����3��$�h�~���/B�1i��}����߶$�j�A�[�
2tE�ǫ�י �*�wo��h��"W�F��c)^�"�H$"ꨅ�٢G�4�"y���d5c)�&��[_C�(g������Q{O�附#�V,^�۫t�ƞ{�����Yк�A>�� m%kv5l�:"Z�L��66PXG�x�����`(�Z����ǲ�����O��~�v;_�tv=O�(�g���b���'�]o���3$�~j�Y�Pi&N��/��l]]H���m�b�ǥ�+Kz9�Ac�xp���v�ۺ_*�"��i������6��8i�&L���(@P2D������y��C
k�KJA%e�rΗ�J։_�_���Mv��q\�b�������U�51�G���4
�*ejdD��z$<�OiJ���
n�L��'���O���`tHO,��8�s�x�W?ޢ2�*�e����7#1��O�PsI9�j�E[��Ė�*�0`�<~{L������||�R�Rc���v��>>�6���E����2=�<7�I��f"��^s�,>����(�6��|���U���dV�5�;�=�ģLEm�,�&D�DKv�_�,��eewyW��,T�_�)�u�T�����q�� {ʍױ������z,9���
	�"T���;��ki�dJ��y��f�s&cZw0����J�h_���i��IU3�1)D��Ŕ[�~���Z̰���Um�u`@Cw����b�:*���o�Dw�7��ՂgO>G���R���
��MjY"�6L/�R �����G	tHv�G�P!���_3Է��'�O<��J�|Y�67���v[5Lk����t�QlC��`q��8f���N��6r�I�e�oy�^��9�P��#���f3�a@� ��Tp�V����� 
��`,)Hw.�%��+<�Sĳ��E>�~B��?�|��ۆ<A�MB�GReR�X�����59��[" �� �f�(=�R��Ʉnu+�,m���U�8�x7��y(��Ս�����E��.;����p:���a$c����̾�%-��vz���Y�\e#��]�1۟��*�R&����#�_(�o����G�>Oҡ�DRh-1��Ɉ����BaӠ�J�~���jH����gO��6�5o)��6(<v����h�ʈ;J��V=�ͅ�;�Ys�[�Ě;����\k_P1h�0�ԮU����2UL�d�
�n�H\�-��Զ�z5#E�=�`Q	E[.����c�Ħ��}xC�x$�-^�J2�Gz�T<
��p�ץ~��i�c�*����!���L�X_Ŀ����,�7�������u�����6J�ј��+����|�J��}�MP��k����X"��1aK �'�1�N׼Nn*�T�	E���B便y�I��mM��]0��dM�ZV`�2՘�(�m�lF�GT2;.��5W��_�n��f��-G�V������C9\���z&u>�,m%gg3�E9��#ƯV�hB������ؚ@v��g+��eE:�e���re��:IǾY�CK[�i�?�.;��"�ѿN}��1aM&��P����ƚI�}RY��ա{^�o6��|��0T��Q�a Hk
*�u��д��ap��$>*�6��e�(�J�����RW��P���Ђ���ptB�R{�,#�ִ��Tժا��FM��q柂S�	eֈګl �S� 3Ꟗ����M,�|�%p��c^/�vg<��k �������K��{�?�K�A���"�r���]`*z� B���a���/���i)����'�h�]�O�N�So��e@���Ű2�]���8�<=կ/���mN�u�̇���P�6�e��x����׹������I��[�q�[�:v
Қ�	��,8�r��$#�������x�1�
��P�MwW�G��U�5I����``��8��"��A�� �>>�s����J���L��eL,ۗ1�[�
W6�S�����0"�x΋.H$U��?�:*�I-��Q���ܵ+�DÆH�T7�Ս	\�Krٽ��.��u��x��$���ޏ6�B�7���s�Α�R��(l�7�F�U2�o�Eȹ�ON��C*�e^�`;;PN���6̃��FK+b����,ll��;�fo�Ӣ:F݂�h�5��K�~�����.���GD�vY�t��U	xJ��!l��z�6E��dqpR�w��:xT��ߞX����xǜ
0.ު�A����]����:�������8]/l�a4�G�Ȓ~K}]tw,a�$a��+c�=�ʮ��rGQ��L�=�o7�zq'8SS��N�|7qT�D2|pa�p%���/�X���Ē��<�Le��������(/��0X=�E@d:V��3���q�e����p�!���H�xc5·�D���˅viXx��4SkrDa4�	�̂}��܏�`�<�
[ͪʀ�����$L+A{����)>��5e�x�"�c�Gۛy*���CT�F}>��Z����s��Y;�n�Rm�,'�_��`'kmf/;Ų4�O�@���6����(]?�?f+"�HW�f�t-�%�$�pC�X�e��	2����w9�zvC@���:߂5`K��������Z�J�����vن��#^�\�> ��r�|��~F9�Rr��O�����H

��=Y�
�u�nJe�9�r�KK� ����(3����oV0��t����JB0-�"0@�6�C��-8��!e�	�k��m3���1xF?�t�5]���N��ؚ.��1n�o��e�!<��������mi^�����j&�*���:KB��rO#�)�������0g�@�5����-J�Ų.��G
�P�)�����a<o.��E���Ggs5�%��Vם" 8�j�W�qay�@	������8����A�m�w(='p܄}E2D�_w:�*��4I!�;aw#�d'7�v���T.��z+<�DLO���C�Ң���zgL�m��2�5rL��E����ۂ�7c�t9v?�2 	��1��	�k�[�vZj`F]���c��@�>W�*����g���:���	�!��{�=�҈�i}��d|�M�D��$^!�+��aqC07ϥ��[��@퀸I��k�5Mm$���k�el�7$ޅ�Ǽ�#��Ͻ�Q��2=����K�5�K�r:���r�)��c��͓y���.F���n�����B>�1�����+�C�f̶������.����o�U�O��F"y�*]%����� �"�t��$� ҀW�Y�_t����N$�k���x%p����*\��e��$�����J��Zo���Z�z5��f��~���b��*��wf�&`r>�X�@$��_nh*�Qa_Z����m ����� ��S���gh�3�$��m�>�?F3�����өҜ|��{������������ E-�ԧx���p0�j��$�*&c��=�NgAe��F�?��FzL�b�e_�VJҟ�8���k���=,�����,k�Gy�IWV�{���R���,:�@�[��la�-"�X�f645\<���^d�{;�觡T�; ��-8 �{��U�+˵��{\3R�K*��Q�r���;Bd�{�[,�����$�ߜ���Ԩ��!9	�9?(J�o}.�s�Yf'(&��4��7/X�3���Zx&T\�I�w��c&_����"��1����@!��EE�G��<��)�$�������?!�Mv�^��ּ� �-Jr�����u��G<��m���r�1�WY�5D�#�/c�53c�-�b�R��x��![��73�8���܎�3�fS)SP�э}����~�iܙQ���:Z�i����&�]/J?ؐC�g.Z���~Q�G�C�o-q�����R�5շ�Z����xecA���_���*�Q�_�n��@� �ك��[�7��z1R��CKe���Bc����մ߸�FE� �.T_o��T�QR������֙t�Ģ�1K��䶂��_ۯ�̽S^P�~>��%����{0wV�/V �gZi����g�cdjl���`���\М}��6V�1Ln�r�x�pˌ�6qqQ6"!�ެ5��6N0T�ͨ�+�>��b7��n� ����g�ͯv��p��-V��I�5̌_�>�$�f���/�1�9��#κ;]IW�߶�vVW��Lʓ��Ơ2�T��/p$�\�q�	h����*�s�`��?%�7w
��饦�Q����,f.���Zb��vo�4�M2Q&�A���P��e�߯N �(�@��a-���O7�\^H��tyq��.A~.u�����0n6�₁�S=e�7��w%�|�����=~+N��F�^�����-'VJ�p��M�-sr��')L"o�a���(���f^�.r�*��.�;�}�^K�A�AYhơL'7��6f+�5m��4��������#�O��4Ӫ�� ޸����B��[H:��f��3�e=݅������2do����~�>���8X6��9�u���+	��_7H�0]�絷�S�Y����특��I�]bZ�=�����q�j�#�Hz�h�35�M��_�FE�M���2~i�4_����ܭ�7�TW H�j�QO��w��|6y�C���U��o��֔�.�E���j�13�aV����WY�~�~��g֩�a�����(�b}M=E-)��F}��G��Ak��IÎQ�C��Y�~IL��3(��wM$����9e�{ٙ��X��>��+qk�V��7��~��5q�f	�r��$b����������Ҷ�7R�ZZ/���|J$Kl6בDU�:��lUA�Ж!�FS2ip�@)[��RmsT�u:��Ќ���3�sAxq!��4�XY� m�m{�۠F�îi�wڅN��XG�r`�G^hk}��?�~4�
OV�X��>v8u��ָ3��mpD�w��zq�Rjt�E-�xy�{�������n��`���������<�;��� &��� ӝ�iM�%º���T�)��HAos�Ł�h�"��5QI����O��`��VSh+�oR����0�kՃ��u#�vַ�p�Pr�q0���T�z�@�$��)��1+ɢ'm��|�c�hП�]�s�*,��zr1�N0����Z^d��^q�ϥ����8ިw���'���)�%�wpt7�?H���da}hc����{�09+�,4������=�*�U�}!'z~_��\ٙ+��x�����\�5���(����Bl��p���b�gF���M�g��-�)&iL{r3-��y�7n(�[@#�A�_^Ӎ���WZֆ`J���hƩpV.����/7d���k��*�9l 6P�p�m�J�8�"�b ��EUH��7 �r���$�R���ݕg><d�d��:�P��A:�ڵrH/��j/�	Vg�a5����7�fKr+x�E�%��C�2HVIJ1b?24�(^�+N��πwe�L�ol^:u{$O/�Vozmޙg��=�����B@�t��[e7[Kzb�d��r�>|�3d�_6o�Jm��ٟ7�T���D�Wf�z��W#~�C/mW�gH> �Oy��8�St��q;���u���A�2��lRw�;^����d�0��ˢ@����>Խ=�*��s3�g�Z�"�W��&�<�p��.�;z�@=@�5�g�+��2T���Ǵ�3���=@�,9MV.�D��?�R�žM��75Xt�i㑁z���D(��˖"!�_�M��9����O ֚Ǉ�7i5[s���M�*LA���̞�/'
o�u<� 1c,e���:��~tJX/k[��!�#�}EĨW����ΘKr�=2Q\�$��/�?�
R�N��D-���/W�_��E��&h�Y-�j�&9��J��сm�'�v �(1%�17:Oz�sc��PX�s�K��l��*(T�An�_Aih7;�눷��`�D�edDa�ZH�3i�y* �e!�=��gQ�����S�Hݧb(�Jl��P����D ����d���#7k�6�	�������'ȰO�=icPr*֌��1�ަ�x4P�GbϹW}
Bdt��<��#��
�O��r]6���P�����d%hR���]z��&_@�H���#MX�̈4����;&.0�A�z�9`�����$���Wr��O��p��Im�%xVz��lz��m�mNTEEI
�����Z&�L .Y��PV�S<�vxbyu�94�S�0���<���|!P>��� <����s�T�[��~�a0R7`��P�80���R��D�"4�% j/����hD��?<�9�*�d��F�- ��V���t�,�Z�v���_�9q6�z�In��n�/iA�k�T�QT��;��)���y�2^20I�R(�)T�i��L'ڝ1���%a��Ig6���qj\oK���T}E<"������Lr�Nh��$v�9�ޝ�á �j���i;��6u5��	��V*��J51��}�vvƿA�ה�}m�ֱ�-�"xT�;{����V���]�)���C[q>�������8��M�=��W���gH��-J�������I����:x���
dx��~.��mr�E�������#v�ǰS���A�F�r�O�Íۤf�N\����j�a�Ԏ3�"��H\G�gU#��6uQ�>���7�����V�.��@���`��n!a[��)�Ry�{�]�8;1�4(B| t�������p�zrU#}��R�6VĐ�P%F�`�IGO�61%^���� S5�U�e���(���1��`�^aΪ渴o!}�@^[��&A$��k�$|�#t�/�3z�� �"�<D�
���������?�;y��3����Ǆ^4c���k�B�L�+"'^�%ؒG����{���\d� cQ�3����͞r�y}; �=]�SR�W��M������W��/�)޻���~S`h��I�^����I^ZE����#SC�:&RP�{�:��- �:A���i��>N��I+v��pѽJ3*����B�ު�$\�=���8�xo�$NҢ�S�<sE��M_�u��U"��&L�sl��@'x&ΆI��CvDRً�T�h{8�d�c��ik�L��|'0#�6�s`�&����7�?2��_�P�-2N ASX�{����_ʹ��n������4�bq�fs/;�8M�R�-j4�z�mpp�V�Z�A
��ʤ/�һc���J4V˃�b�v��,: ��Bu(ը��C���^@[�bk�#\��U��h�=mc�á���IC
Q���zAy�����_|�/�U�pa_J�U������V6��ว��&��	�t�$iS�������Y�++%��J����uҫ����0�<�X�衣5�!1m|���xya�v)������ً�\"�g�x��a3`	�>lwM��fk�.�T0O$̜��u$�~��2&�s��2���p��
��/5%:�H��r�By��1���K@�?�&ֲ��d ��S¸:��1y��� ��U�][0�t|Y�ot[U����}����4Kq���Y0�#sK[LN�'�r�P�*�Q�r��jl�*j�>�1�,��v��L�u+�+�4��;�纤��_`�q!h�F�
pYG�j����p�rP:&���}	�L�V��IW���I��fL { `��
κ h�����d}%��������т�`��<|F�ρ9����"�~����x�/07�&Lg6��������y|�Պa1a�ԒZ��8���_��ǿdf�=����=z��+1+ft,? �Pl���Q��4�l �b���BʌtrHa]+����Ƃ���u��@�����|6�����99�I4°�u}����tg��Qz��&I.<n�h�`��g�j׵q������t����d�0l.Ji�{�+q�Z���������-�����/bIv��I`=���˜/%C���ǲ,��!�u�~C���ӱ�'ȫ���1X�Sʦ[�ǒ8�9��֤FO�.|���,S��I�ڇA��9���sZO�wU)����"x�Ay�nw�wf��
�%��P��9�wu�j�R����շ#����b�T��#���[l*�i5qO�����e���nw�Mو�U� ~�@�50k[����T@�p�q���py��P7�S(��\]�gwt�~��!\z2���=�O+:����=���vǋ�@LH��"ڨF������-'�Ow���<8!���ߔ�6��{�|���I�:ϫ,�`6�-j�E�&'��v�+�+d�ukη�^����]P�������>��F̤�����`$�⻎[�T�  �xOY�,Q}$��3C���ću �J�Jp�w_�s��%쿱.��}?�0�f���^�C+o����]�2��>os��B�t������!�iԟ���n�YT0uN� !�޴��F������5(�bd� �Jt�ߩ�eR"�i�
�x��?NӒg5��-.FД$D����� *����̺��x �s�Hf,��c�|�� ]�}q���;�y��r��p�7�G�ŻE���Zv�3���7�;������0$�������)��?� +�"�3�͔ i��g���y�gb�2�3�j���l�fT�=��8qm3����`�����oP.3VB�n��Y�cI]�J��A�@rv� HS���$&7�Nn
�R����7�p���$U����?:�+��GV��?$�Ԡ�/p}���S�ȸ'2r�&��ڰ�ۋÓet��LR�eԁ�5O�Hid@}�|i�3��뗶_j��훓pКz�\oc���.��m�3���f�	~��m���;k�Z�-�*�z�r���� ŷq���z��N}g��*���rV��ψ`�X�7��x@��8%�'5#`�bq�d�O]j$
xb3q��AD�lJʢ�x�@T^|7��K��Hy�=c:�jk�D��ɼ\9�޴q�z���Nќ��Įږ�2�!$���1S�\Y�Ե��oc4�Ɉ�i�o��A��>���X/���B�!}p��H��v��k,4�:�y��W�ԇM��j�^�7��o� C��(�'�o9�!��!����g��f8��ܥ�fVg�AmΉ�V�R@p���w��
�Ö�$��9�!�� g���~	�a����I>��~�L�^c�1��)��(��N�#��>gr7���	�\��ӓ���A�@�J4:��<��P��z7�1�r >'��Vj�8�jJR��!K�H��T]��S�D_�>\,�H���t@�O4��C��E�-�CV� U=�S,��g�>�I�n_I�w3DTEoJ����W~ ˉ���{�3�l�r��v��%Ȧ"2*��t�g�k`�q��8����Z�)}Z8�)Gm�ざj�l�Z77BnJ�7��㦱j?��5~I�wa@���%�bۂ�9���&v�� �um���?���hc��*UT��({��R�,������aI:��Pm�Ï+�k2�G���a��\�;�՝��#L�.~�4~��ϝ����YÍ����ߊ��G�	��HC� W.|�P���}� 9$WܝѪ�9�>�D���H�!��Z_pQ�DWEo�Uy$=)840����vb{��5>��n���*�3�P�dk��OY�(X#����H[z%������J�Y��Ђ���ր�U1#�u%.(�T�7�Ɣ4(-u�M��,��������}0�rm�m96���|9�Z+�~�"�ݵ!X1פY���B�t�Lbl���|�D�@���"6~W�B��3���_`o���(��>�ʞ�$���,�a-C�����G���
���ރLSD��WI���I��1�e��k��o��$|,z�p����� t����z�n<��i �r����w��2f�TfU���=x��x8ҁh�e��Q9ZE�x ��؁�_Mt.��Y7��q�:�r��O�#��&o�v|��Gu,WVG��$ ��u0��J�@2`����=/�[X��Q���b�'q�3���f���:����i^��؀4���*���&Z����"4����69όqZ,�%G��)ד_-���+:P!o2�P�������uk���F��|�pp��VL�~- �a��!�?f_K`ؾU,�g����=/�a;�V�OR�E�hG��G��`�~��9��3~�X��Ҹ��6;�iV,�x�_G	�����>���N��	�$���W�m�6�����֕� �m�����D�'xޗ�-�E��.�u��I?�](x]���έ�&PӍ��}J�=\/�3���ex'�LI-�A�'�&z�s�ɛ����C��|]oڏ]��}iK�
@ӻ،�8���m�ʪĦ]+2��a�w�7a�0����℞�{ͬ3u��3؆1G_N��R"�������Z��h��Ǽ^eG�G8�l>L��&�ל-�q�%=iR\�'�[�k�O:�G�pk���$�qS�+��^�Q�c��Hn*�['�^���I��m���},r�*1�-�%~D8V!Lo@��^ֈ]�ǻ�0�ى��SSr�u��G�晰p"7/f6�������d�=���8��+( �^"� ƭ���}i�"g�PԿ�%��-ೢ��� 3�"�`v�T�*��8�s��Vٯ@�mq��������d_���\eKRQ��$��!s$'�o@�"h�IF�lY���W�XNޔ�c�<��.��qU�p1���g�4т�}��� �"n�=�ЫN�{���{�T�P��ToM$+����&�Ŧ��2{�ᖰ=Å�~ ��(;�gd�²�@�YϚXZWmZZ"X�e�C�,4��e�_�C����5�{	��R��	������ǥ(��J����(����49�(;pA�w�����B�wU5H�u�[�
ytV����_�̶s X��
R���ݨ���&qz��6kEeFz�"���D&
Uag�^����t
,�۠cQ|�뀨��EL��W�[���fl�<�
s�B^��J)Ȗ���ʋ�V�Mvy���T�f��gT�i���/8yǇ����I����ᷢ�'�v�
��pb��,/.1�~�l�D�Lh����C��V���*��[8��72�e@�}���&x��bٞ)�}'��3Fչ��B(�!i�un-:|���w���W��1Ƈ\��h��0��Cg��ur�[D�t3�,�Z3��ҹ:����Ӱ�����q|� �W��b�v�Z��^�Ћy���)�XO`)L?���!����i�Q��N�G9Fa�i�GW�G;u��ɂ��~��r����q�/v�d
���z�}��h4[�t �fB�T�x�5�h�q�o�7�suQ��d1���yl^P����x���	Q�x��{6���P�Z�;�L����s��R��-�5�|@�B[w��oN���EiL?,�h�B\��m?�KA��Z߬k3"��D�������o����vn�����ۘ:tI+�Xz:Q��Ύ;FPy��1��<�IhA���i������险\>�y�Tp"��	(� v��DJ�J���@��R�'����Vl�;��u��3���	��CX�څ��\���/��p{Wq�El��rn����bGCM�=7D�M����|>����Z�$�Y0�kp�v��-�Y���ԚQK���2���2U-�F�nL��8�pw�^^��3	�I�Ӧ�:��r� m����C"��r�J7��.>i$@�3����n�,T
��7`;�ƃB\�����/���g���R�`T:�]����@72�$�"_|�wdm��'{z��Fm������
��)�y �0ƹ�Zy��r=�V��#������2��Ӗ&���꿦M��W�%�Yk���2�jK��*W�'xV�M������*��{�B�2�W���v_��4ls]�	T����U2�x�xI����`�_QH�\ys��ב�F~�/;�&�w����X�d�`�mxR�h��gR,�]e� ����d��]"[�	a�������0�yȞ��q�&��(L�g6���j����]����r��˙�?
����l�?���o��,r�j����7���a=Q��� �~�5�r8���Y�T{���;��bd)�q~�4�����Ŭ��طwv�]x���6V�]_|��֖U���cZ�{�j����9r�K=`�N���������-d���Gu������4���v���;<���Y � ���6ؤ��S
b �������<��V�#ټ]&�ӏ��kϚ�9t�wv|��_�*�L��S<�B7x'-����0��/����O�N ͅ� ͖��V�N��!�4�q+���?t��˵s�1\�@��������7�IzF���(z���ZwQ�e��<�y�hf�L1��Y�p�𽬴3���Μ`k:�a�M��fw{Ӕ\���xf+֛�e��8u�1�ѬxS��_N�x-� �odZ#nbk�3ӫ�x��aJf3h�����gerq8�6���2=���1�j��	��7D�q.h�g"q�Ԕ��嬯b��2�i᥼�g�و}��D$Q��k3���W�/�#2|��}��;� �r7�b]��\���"���%G�@���M��x�������t�I8�C�d��!�E~���̡\EE��#"=�1��1;WD�[�:�����C	>Q�>�s��v���A?ndhӽ����F"�`,�BIhFfH��OoA6�.ھ���񞏛L�I�3X�"S>�����z9�ǨHj�d�2�4A{���������3x�pu^���A��s����U,绖Oǚ�!�N���*�Z���r���N�<B���:�xJ�(��:��PB9y�0�xF()�%�#�%�CX?qh.���h��E yy �9�$1]�}]��#_tq�wlk������}�a�܆��_��3]2nLh�4�� �u��֤u����z�/��	݄��lpa%���mќ�_V{�qo�}�٥Ȁ��z�?{�o����(�=|5����i�BG���͢I�	�O}йAB�5}ĥ���(r4R��S;��]a��t�h����tGߝ�--��|��A�F�VR���)���%h�vh\?+��.� ������z��?���V0��!kʏ�զV*&
xX�
�Mf_��I7�s6�9H��j�d�����24:�gzZ�|��a���sg���ʌ�S��7��� ���������`�\ ���W2H$f��2�웓��ӗ+��rOZ껮q#���Ja����3���[�p��^:���S&3g�`t.3��Y�4O����X�W�:B�dEP?V�Iށ�i?1�=t*���<�ؗ?���~�r��;s�߁Z���
WrވtLw���:�:�_�~���Tv~;��+����ڶeS����rݮ�W B/��i8�߀)SY���z�Cd����9�w(6B��X!�w�Yj&v��,���="�q�p��͜��Y�:�#š�kUM��.��[gv8�����2��(��o���Y�:��@�����E^G�����fj����A�Ը���g�)���Ww[H�ʇ��, t�L�W�ܴzM�lL��l>�Ub��V��m�aJ��-%	CT7����P�5�W�q6:�)C�H��3A�`����c���l�3g��k���Ф~(���9�|�B����pP"8�J��`�i�_�!^�,�j�s���$�c7
�J�t�,��icPUZ5��/�9u_rl��<J�ٻj Ph��n�7�#�B%�>�,M�<���Z �b�P.�a��=�Ya�V�x���1a6�o����~�#�CS�B��\Z�m���մZ���@�l,k	�w�S7ܗ#\<��j;�S<	g9U�yzZ�1}���"q�sF^_���ua�Y��M�]�?^ɾ�<�:"���@x�GT��BKk}�5b44���N�GK{3��
���>�6��_*ҟ�?�L�8��5/��Ý��j�1:���7V�瞔�|yi�U�KŎ����"�*��:ޫ�h<Ϭ:6�hC�B#N�I�HPɧ0��N"�v��Q�״?��*U̚`��̀�tYU����P"V ����h@���~eJu���(?s}�$�x�Om����(��}�֞?����&&��"+=�"iHf��/���ft���t����נ��Ri����a����~Wc"۾�#p�4���r5�S.��_�F��$̦�{�]��s���R�M圿W�gމ�e��;=��_�hk�SO�ڈR�p�[����G�Cܡ��j�f5��l�k��6�z��	v�2�V671��'ĊQ�Y�;��L)��y�yHh�u{�T�nڄHCC�}��o-���@{O��+Y1y�&���zpMq&����P��e_l�8��-�8�ĵ�ݬi��"}B�<%�'��C��N3�C�^��X=Ooِ9�[SG�K�4��� �}�=V#Sl�%b������3^��C�C8�*�2����3�R��Q��\邃��W��	�a��LI���g��'��s/M�d��X���.���#r�{k�����Z�b팏��d����\��޸��d6�������;=��φ�<�MXq26�c�W�.����[�qL.1a�w�d�B��?����+�H'a�ę� (tǆ�nU�V�<=���6��ĭȡ�>Z�Mۻf��{0MJUj�=��+��������B**�����E�I]׷���:��>��
.���$����U�)��s�`�?M)(<�ū��,��	p_�`OJ�[��
L��/��K�E7����ט�)���j~�7���f�a�?�{2XܔL�S�{�	�hK5�{�WW�.�V���{�YL#���o��� �%�ѳrݯ2�@x��Vҫ���q���{�;�<�ȡҹekD���M
�ݠ�Ӓ4�a�����T�qX���5m���pqD-�M�Ϛ��lf��D���ƀ��E_,7ݛ�a��G��j�$��ۤݔ�p�N�{��� >��2��"���gœ���P�x��9ޢ�hw	+!�Xܯ���$wLs$B�ZA�*�B��{<�Ko#&b���
��J��|��^W:d{��<o�.�v�#��AHKR��B���p?��3�|с؝1��i0�b{��V/2���dU�mZ.;VO�T����܅/2��~s\\z~��Bu�.��-'�<~��f;��S(��I��4���tP����Ə��[ϻ��s*�;d1 ���,y�z�?N��%%��{�8�.�4Q2\���~�ȹ�������TE�YяE��*�.u]̈́[�?o���ϛ.�G�s���L�N}B��8�7���$:I����$x��a��m�9��ee�k|@����w@�7Jd�X�S�),�9:�����O�z���"����ʲ�m��-�nt<K��CdW2J��X:�~�O��P�����G�ǖ�y|���P�� lGꐧj95@;��hwry'c��^�,Q^�"7h^�3�z��f�����kx#�J0�!t��&�t;��	􏿷��衝�N`��0����i{3fahD���i*�2-�t1�h���J�����A�-�%Ap��7H� ]QL���gG������_oQA��.H�p��Fm��I%TZ�s&B����y1����W�ao%��9-V]~�i ��0#&��f!gZ{�,����,������axG��D�OӦleQ�"�/뎪�@d1��"|�r�6�P� ��k��5�J�͜(F��FI�QBD�2��7-���'��N��a8��Im�~>0�R,��(G,²?�*�\Q��;��h���Is�jm�/7���/�ؕ��wb`Հ���� <%�() �?<�!DΦ�8��\�6M��mT�c�d��;�T�q֠z,]�|s�- �����i�q��v�-��kc��Vo�]H�Dk���j)̒�^����n⥾����\��I������Z�hƢ�-*Uwl����Gå�.��sL��/{n/Y��bh�����ҿbJ���w}���i��MyY6$� ��hRbx��� ~Ç	c�=SS3�Ӳ�.�BSE���:���̬�z�U�O
0[َk
>�at���4��dl�BU~Rl�W��	��S�.������U�.!��c7�s�'�>$�LS���~y��kU����w�j�<����ۘ���doz��à�� ,9|O��L?1��|���u�Ӓ�ǽ�5!�եwr��tUmV�8�29Pp+iyl~D?��"��bg'�ՅV�?�־���2��(�ގ9�$-�Bs��k\)]t�)�sL�	FX'4@r�/2��� t]6v�1���!�"KI��D�	�N���
��P���,�`f	^,���HZ��]�Aшa�-VU��3�b�[�(k�
�bA���nް�[�A������Q��c}ey��
���+"N{ڦTW;I� �;>�8����א&ō]Ք�z�qӤEo�.�⽓Š��f�����}x1�g���.q��\��֣3��t�=�l�^�g�t�h��|�H[�\�c�25�Α����T��T\���������?� 1�@K��ڒ-�`���59kQ���c.4�Iuw�i�\ȭ�Җݥ��ٺ#�(k�bL���r6�ٓ���hX�#�JZ�Y�l5�ᣫ�̌1��.- ���-dR�0ͨ�ؒ==-��nyR�������w�F�^|�e�u;����]JDzn�$k �6��1��hQݻ������@h�|�����h��6MZ^����|7����
�--Mũ�6u}u�-W��1�+{�*��<h�]�8j;_�n2��4��f���U0�/J�.(al�h:�
йq�K�҇�s���]�z[Z�_�4���o���� 2�#M���=wR%<4z�]�g̱�؝�q�J;�/��"�G�X8���]��a^��(�B��u�`�%1�'�.�+�a�M��%�+�j�����sԫ܎NN�ʃ�e�B
ť��L|ǹ��5n�^�"H�����%�lA�$y��ǍTc���8Y��M<'-$�.�?�2�{�3#%s`-�7h&a�Z�[Μ�p�g�`$�>7���� �����V[�%m4~�n��hvM�Qg��݁�Ɏ�/�.5�T@ Hp�������*�vgh��i�wˠ�ޣ�Qa�O�#,I�z��c����f�XgG� �,�v�g/;^�^��y�>6,��ݹ6��/<���%��|�x h���	Wg��0(����ȳ
���=�W�ScM�m�i��#�]sa3JL��&��3�p}��Y�7�}N$3>���	��L ��Jg9�\H���tҒ����Sn7�ʦ�9;"2B*\���[�/�D��������a�LvV���T�Kt��Y�2c_�
\��d(�`�d�l0��yqh�DBmJO @_���q�A;P��<���L^��6�ZIym��M�.#�sK8AD��JU]P���Կ����9��Bz��V�GXƫ�	����#�@ >�c=��r���`�*{#iLG(>a1�����6��{�&�_I�ř5�\�:/�������LJt�u�\�an�7��Q!~
�;7�F���\�Q�]��=�8'�0�J5�սA�ψ�^��(/�P�}Z�g��OTp�+u����L���o�5o	Ju�qZ�έ�׶�0���(D�E})�#��s�o^6�x�>���B#qQ!�ҭ���V��!��q.LcI�=�mKB�t��&*���q� ]����Q�`n�9)��R[�~.d���e�K�~ �S˵���݆p;��TDps�SDI�\|ݢ�O�[�}g�Y���M'�&���rt��j�������5@�Zx���7g]�N:H��E�i���Aœ��\�@�Lb�O+1ϒ��hʳԜ�߸l�u�b���?��w�Չ�o:7(���i��Y
�<���;�TǕ����Cl�;�C���c}W?�~5�7��yf�N��1��/��&�g�ˌ�L�-��7�H�#�n*�X��MI�V֍�o#�H����K�Fݹ��¡4�8*�T0Ű�w����t�,K(+�a�'G��E�ō<�I4 �K=�H�= �������Fȋ�6�I��(�I;Ejk�#��"��,
���[��E�1Z)��@�p�Ԓ�������CI�o�Xl�rq�2�l�2-{W���n�:�&h����� ܱ��4 1���C��s�"���iKߧ_94�W����-�mK����W"9fE�g[
���F�^-�THLt�F����#�E,�M��n��wKɲs�r����n"�f�����fm��lz>�Op��4(c�������j��@|jݔ� W� ��NXdyW���kc����2��Vd����O������+ 7��_D�]�a�uOJ( ;0�a�հ��K#�q�v�{�K�;��!\�=mS��8�MN��%-�^]�ʂ�Åi��i(�(sk����9��1Z֫�y5��H]K�rK��0Es���qq�w?��c	mY���F3ǹ��z��^t��u[�|~��¡�6�����;�e������)E��x�A�%���s�=��IƟ<ab�cN8 {�V��j>a�5Z䁠�3%�zK��;�hPt��UQ_0�PH���#]	|R�dc���M�KB!��5�e�bt�
�@���~���G�� yGw:֘�/�9 r�Q/Uj{�P��Lн�[�����b9aT@څ�,cy�:]z\q�^ځLp�N(��Q!C`��H�*p�m�h����t�Ӽ�2Ł�
p���%�g�!S䬲�'����bx�Bʠ����|K*����ڄʑ�J�r���d��_ݥl
�[��|�i��o����1Jz���.�����8��ؤ��p�Ԉ��m�(T�!E�d�0����pv<�~��@J���V:�<�hD&��9ݾ�j��0e����vN��vg�=�z	#I{�qV�����6��P��N`�����2R�9ږ�hF#uӐ����U5`�M��q�tX,�eĳ��e��]�Å]w�d�����~dU��Mz �������S�'$����|A&�꺁\�;8�'�R�<e$���*��s`��%�®�酟�m4��/(	?�t0=��3C@	���TR��!�[���u�t\|)�g��a����I�#������~XM�6#���Se��R�?�^���A��k�*�/-h΀���$(�0%�z*�Sy����2�Zz�Z�IVIN�X�v�'y��&�##�(OS�4���aw�s��Ce_���x��9M�߸��w��>��]�ټ��9��]��3C*�'F!=�]���>���Z~R+i��~����X,B/���d��v�4��V�uR��o�0jkp⁤�P��m�&;�X��C���Yk�
����R!��S�^�DS8���r*���~���J�$UI:|~o�&|��|�H�6=*���C-�"ʄm�y�oP���[^�1`t������K�E�@|��g����ΆX�!dz<~�\�brN(���s>p����ٖiε%�������3ܯ;���
QEU�H������uZW֧��W��!}@4x���8�
��52v�����	�A�}���DP��7c�xC��In)atڒ�)OM}/�^�n2�g�нe��;M�����>t_0���lj�[W��{Z0�`��ڙ3���E ��I")jR�6蝤��G�Zb��U��6t���]�h���|��)�NLR�n�>�q ?�n�?��I����zIa��>����s[�.��KZ��O}�Cx����B�q�[�����E_"�_[q�fe;��F�x�˹c�e��=�i�@h��=$=6+��ٝ���������E+���J��?�]�o��pj'+����G�O_s�5S�����t���E���4�_q��oT�P���;[?��;��1Z]�5|F���d������� )�n�]�F��������p��o;epf��_<|����6A��Je��b6l�o}�:j�c�D�M����2UN��]���|����1�)��mf�*�\t�V%�n�;Y��;ɚ+rWv=��g:ؗ���1.O����xs��D�=���G��Ί�0X�x���F^Xu.u:�yt(}���9g���V����Ȉa�\�"��I�����Nթ�u/���Jm(�R;��^i�s,n�+X�K�,��!��2or����IT_�����Jg�i�Q��a�'�]�[�<�3�vdG�U��G8�)A35���J����\������t�zE]�idBm,�fk΂�t�b����-	�4U$�E�xg)SG��+qg[�a92�R���?�f�?b�R���s���X͘�Py9�R<?��"�j��R�&�Yw�̫t��6ó�Ձ�t�4�[܌�$*�Vqۓ"6�J�1�ޮ2f��a�ٯ��r�څ�{i �c��á8���nLPH�@"I7�$H#^�kUd<W~(H*���p�7�n�}�� �W�ی�ݽo�to�������5�߿��_�R��j},��A<�7��{��V�%Q)&q5/�5��K�URR���G����]��;��T͋B�'ݕ�t�XOh����31��<�;�X�g`�h���Y��o�TKMF���ǘ����@�V&��a�e:����i(E0 �m8�f�.8���i�7o�BX��X�_�I<SZ։�^��������c`H?���v
��A,w��װ��^j;�3�D[�;J'�҉��D-(�ɩ�R�m}{V;�꓋2��?P�|����o��5�ޛ|���7\gyV�G��u}��dt/�I~7��~mE��'�,���T�ɶ*#���6t���Q����@T_bnD�:���,�-�!���6b��?��z��~��@at�zP��F*�׳����Ȉ�ٰ\,��V��a��A l���<WH:���H�>>�ھ���;�B���r�n�x�{�����+��(L�K^4�$�� $a1ٕ��}3�;�l�m��Q�
_��cD\�sDן�#�(L�j:�Ǵ�?�9��F�}�wJ��l���]��w�s
>;וU��ױ�j��NĜ�BB�ԙʏ\����f���|�%M�Q�3Wݱ͉�Hw�3�q �ޏf�MQ�.k5�7�~RV=�ƪ�c�c�>f���t^�:�+�+ø�ql�~~�����l��q7MO����~{�]Q�����3O%�m@�o�6���+y�_��ɎO��2���9�o���"9�kS�(���B����a��
q�j!]�-8�O�)N�����ʆ/8"��Gu�~�,�
�aG~kL%g�OT��Z/����[�X^y�"��]�e,q���2U�/E�7i/�E���s�1� �l`�� K��#0dl��Q�w�x�ҥ�C��*:Th�B&v��؜Eή���{-����1�FNu�A�{YR�`�%�NV������z��h�==�E�ds��Z��"l֖�^�ŌS��O �hU7�dh��Q�\�*mjg�/�7�z��AU������/��ˆ����,՟VMhI*V�S�7Lpk��k(V��%mdg<���A&�!,Gɾ����7wW�r�\#7ȄM��U�Q���2�K��D�_�4��E���L��w*?���P�`�E�A�)���ߧ�a[i9B��;g_L�uE���|�A�$�ir͊5���N�>���E��\_7ؚղ�>�tO@Ю��,�������y8-i�Z���ټ��pZ ��ŌT*Z%��G�*:@�!b�����A>B�Gz��A&	ճG�*v�2<$~	'~�K����({K�g{z����P�K��^� �n2�|J�h�5񙲋���L�,����c�[��'(K�j�~�4�҈A�r/�IR�E��h�8����V
���`�4kza�[��d;	�*��0k]�w���΀�4\R�dx�=M�ǐ͇�A��@W�}̗���
��S,P��ך��1y�������y!�*�2��q�\6/c{�v�﫤��x٥5;�gH�s0!� ߪR�V��n:�]@�ۋ��	�[p������#\����5B^$��3�B=)�l��D}��k��m}�5��e��Z�gH����b�T/����ڍ���� r�F\�B�L�h���0g7)�,�c���>{t���eB���˿}|�����A\8L�P�ѿo�vA�$�2��Ԃ��.,����P+�R5Tr�󾳛��~��E�Ic���1�R�.��8Ш���C�7�ɬ"$���_�7S�X��ߑ���(��E�{��W�)y�p�g�S��p�5|QA�W�(����%x�.��u�s� _l����(4�=}���;�B+z65]�伮Vg�F���Z��Qy��i���W+���HN��KMz6n){�5�Ysu����:Љq��M��<�pX��h�������Ft�U�7��x���M֍�=2��펨y,��C<os҈�׫����]��'�<Aʾ�q"������Ez��9�It��ZO�Di���Փ׹���Z�@�v~je��K�C��5(5;�ѓ֕�:�7�������2�G�C�L4T������I�!c�!Oշ���|*.����P�N�W��_��TU##mT�������)�ey����"�5�ZD�6����O���a�
J�;���`?��G�5�}��?	�\]&M@�߉�����pT�����
t���kY�O?ڿd1�*�z�h� t�2��8Iu2��^^�k�b����>u=Q�)���YIW�)|�%MO�&�L��C��*\�k�Wb0��ѳaU�~�Xzʆ�������<�@�[�����/�o�I2���e7�uǘˎ`��srœ*1ۊ��Uc)o#�~c1hf�nf��G�����)�[
K�����!�b���޳���vߥ��&�?o[%IЗS"$�<kpl�8�.aTMg��Bߖ��d�������b|�|���-	�I�Nj?ѧ'��
���g�,w�F���PmC�N^"�L�	s�^t���o�#�����Q�C}��;&O`��`���p3��}��a���k_���(j�V��U"s.��H�a-z[���axξ��t5�C�3Ք�z�}�a����S�39;���0v�[B��=�.~��.)w���2�u����L2]�V�_rH# �UA��7BsUZ��g��C�I���������2��i�4)H'�[��7�1�2��֐E�$h9����G����	d/�!�N�lc$f��f�=BY�2����U�,���3F���w@Xhr�h��|SX��x㶞�D�����>Oǎ�B���0稲������jnل2r]ϙ��
Vɲx][��8g��6��s�Z��'���ٽBL��t[Or�%���������b�95nl:�_��i�	*G{�Lȓ�Byf����:��R��c�0X���e����������nlZe�Ѐ�����=Of�������_��
��Hu�Qta���Ƅ4�gs���x��&9�&zQ��(��d�F.��Kv����M��F?å�=�
*F�G�!�u����u��R2��v����w��J���Z�<I����9aa �D����uo���ĘKF�����߷��q��''�_�8��{u���8'���!��1�cm-�l^2{l�.��9
�{�Y�{�@�h"��aIL����+آvX���.��"Ȁ�j��{&T�@��~�]�r�u��BΩ2SvZp��"��8o�����~�
ҝ�6
�K-P�)~D����z�pKQ�z��"Qw	��U[Q��<��΄*=��Lr�ḑ{F:Yq����d<Q ��\����,����9�.h����$E�j���*��:�9�1H\?&�:�.{tar$'5���9�t��@�*c�ٮߘ�eDP������ �2�<���E�
+KZC1��	 �:�.��u�M%�hmmk݊�\˄��	���I�=/���κĢ$�#!�#���(���~�~��5�<z⽻��p���{�^N=���߽���t�����$h�b�'�v U.�~:G&��|���Pc���l-�۴ُ3=DZ�ČƠ(+��y^��T7�l��`���l�dv/y�Z���WhB��A���/�?������^y4� ��4TҾ�c������|K\jY{��������E��4�~`��K��~M*�F���>��\Sܕ�u�3*����j�RW�։��e��ʖ����(�9�O�G�1Ť{�Û|�������.�Bj��Sd�zjխ��R��9�!.��y~�B�~Է�\�O��c�ne��UeQ�0��83i�Pt�.l5�E�����~�vyM�NT���9J�Zw�X��ߴ=��2^�3	���?�H�P�K�?t�ǂ�$�gm
�*Zvn��Ѝ=��<�}��&��?����mJ�va���k]� Wy^�b���+y��$YJD	�uIĻ�������u�%@}<��Z0E^>7�̗�g��1@(c-N�o\�mv R��ұ��0�2vY��M�?�b4����{�S!����=t����1`H(b�B���/%�� {#�󤍊V0HJ��5� � k���Y��^Z"�½h]��푪����ٚ�Y������	��������S�N�$g7�䇨��v��)��|�1+���0�b}��G�>�v#1��ƭX�u��9�L�I8��!���,ys���%�4�\6���h��:3[�_e�N���!_�v���sv%�����z4��$Dx^�}�u��_�}���|(�S����a��O��z !�I�Y=F�ǇL�:�P�	��Q��uauIh����d��u �Е7�����D�f�:��4���u6K�CK$Gr��7��x'��͖Gk����cd�ȣ�S�0��Ac��,�����e�.f�D�ˢ%���xM�U'k���p�R��6R�K*֏����B�>�BBn�+]�Ѭ���<2��&P(,=h�ҫ�lo��	��3��:��Ξ"y���붻�����~��ST�J��Pf{�/��$�`b:�6aj7r�H������~��@e�{��J��iD�t��vĞ#��Cr>��90��o��a�\���И���i�1���[j얽!�]ΐ+�26P��i�m��E�T�u��2�}��w��"�5 ���:���[ލ�7j���:ӑ,�յ�	�Lp��w(���#��	E�z����ʉ"miY���-�+$�����o¶܊����(��:.�q�kRJ`�O���� �/!ю�,�kW6#\-�e�e�
հ�} c�qS3���#Y4(>}S5��ae���C)���<0\i���O� ��	�A�*���ſ��U��n�̦��K��e4f-Ǭ�iPnO�֡�е��2���D{r$�n^�/:������cUBx����<Q�Ĺ�qA�7v�N)5}�qE0��h���'`
Rͺ3U�����q������g��렻�[1�M������'��H�uʩ^a�%c�V7�B�_P >��w
@!S�٩�a���LO�6%tC[eCeG��o��^��JS�	�[溽R�4�[U'�;���Z�T*D:�w�2�(�7�q2�5����p�4��~�\i���x+�I&���Ç2E�ƌ�s��?Y���J7&"Nb�k��m��+G��DkkIk +�޾x����.Q�a�bx��,(��l��OE�������Q�:��8�T��q���xli��k���bK�6!�nP��Zl8U�wh�p��+�䘸��G�Y�O�c�\<]�IF���\���f��]tD8���)��:h��̖�sʊ*yq> ��%yS	QT%�A@o׳�,/���Z��qgȓ��n7<�*[r������l#�S'E^l=!��.��y�e3�%ª+/TղS:-�mw��6��>8,�>~�Gh�6T�2
�"p��x9H~�����8��GwOW�7Xɢ^�JO<cu2����ݍ3��fgb�Ԅ�l���9p
�:��+.s��֗�ڧ�v�4�XS�H�1oBAa�w������ H�9��7��kR�^k���f�S��z�=\v{x��8C���Eٖ�����o�m�>G��a��Wu�Q�˄����Z��Z����H*S1�$���>�0��0E�7�"�%7�U��Y���h��_��|�6�8 �C�5��j<My����~�ND�6�~X�߹�^�;��1�ɑ�&��Aٝ�R����b��-�H��"k�d�/co|�v�I��f`O�##j�����^�!R,�jU�!�����g���؜��qS�����Jy'�5�]�K[�E&�gE��A�T�JXH;��]�k�� ��fD�J����gt�>���ӔG#?& '�t<
_�(|=�M���&7���T;Qrz: �
��f��L���S�ec6���K���j�i*���I��Tc�E�E|���^.����T�z�s�u��� �4����!�lH�*�~��q�P]a����i
�cCv7�#;D��)���6�<p��G�S7S��TF��ISbI���#��m؎���c��j��_QZ��ؾ(���?4<lI��HR�d֞C��-NS<�Nnݍ�ax��NG'����r��D~n(l�M�:��+]�<t�� Ɣ����;g;j�EETi�	�B�4uS%�W���(,TY��Ka�/u>$V�������b��7BQF����K��ox�`+n���A�IF@,��k5��E��c��ֈ��CN��V�R7�����!}�(�3�DT+�EA��g�]2y ���:rH�����|�y��Օ�?��]����b$l�2&1�ᎀ!&U`	���q�%IO���s�a�T��V�u���x��eJ��-�3�i�u�R� ��iA~ûȪa?�{7�B�o����b�qK-����Na���Nb�=�nym���U��(�]��'àwi��Q�J�>HS�v)��>Q�����O	(bPX�H�S�l1G�0i߸&sp}�lf��S��}��}nT�k�Y&�fa�����_*ÙR,\~:2R��{X�sŧ��Y�f��z�i]0Z4���$π�w��O�(�B�-j={cη�ݵ�G<<,e�S�0��9)��b���Ob��>�bE&�@+��f]�.��>w{M���D3�cM�\t׳��KJ|I�"Afp�����2 1��i�7�s��2Ҥx<8X ��擸�3&(�yӃ��c������3�|� Y���\Թb���RjOo�l�� ��O�=�105����3�/+QW7���-���S3�S�� .6�A����}�%��U�8%("�~�/���3�Y��쟟z��)���@=J�1hdo����xw2�S\\���D?P��h��U��c��٥�[�����d*��ulP�����
�ĊG"��t�l��K�^�~@g��eѺ��E���6��8>��p����$W!F�ɰ}�9�M����{�=��ɝP���W1�T�_6䶎H�<�ѥ[e �_'��@ФP�zڮD\�����]�^��,4�2�HW�����?�S�){Y���o��&qetR�=��8X��6��DjNp�Bh�y�� ��6Z&�[�[�����J�.7cl÷G۟H30>.�,����ψkG�#�s������9	}W��zV67��{Q���x�|E�u.��"�?Sh�x�>O���\Q��r4�*ڜ?���7}%�;,�kv�|O�ៀ�t�n�Ӛ4��2��p�X�a"�[������A_�'~�O�8��`8{ؘLt%�[�A����DXi�L���M6�X�5�� (�chq>�&G��{�	�/�:F�V�qŞ�߭h�w?h���D wo���i����LU�.>���M)O]U��21��W#b���!�Z&�$Ji	i���@Da~�D_s�Y��E�/�K%�	�Z/�HaJb��,4\O�X>)+�U�������!.�� �h$ fZ�5�
��u�4���]�A��2��@�2��	�C���� \U�0|�u/�T�ռ�K�6˕�R�t� p����͜%R]Z���XOM|���N�#�b�<i:vx=�x���3��9&jv�0�N�BF;u����g��:o�1��%�"�ȫ��������dp<��Au�|/pȺ�����M��y+W��Pz��:�C�etR��XC�
����)�X�^U�ƺ8V�Ct���)@�
����^�Mﴹ��Q�x����*&��!b��U1W�=�ʳ�Z�h�ޅ��������s�ϲ�Q9�Zv���tZ��#0	PQ��]�QyPC(;�]��<�PU?��8Ɉ��IU�h�M��&�B.�Xcz8���,�9��1��u���2����qGĚ��ʎ�D��U�V;�����~���Y����Pk���2߮#lS�J�\�0�������ִ��ya� O��:�����]K��՗p�^�k��I��X�L�'�}n"n�A�X��2��b�Ġ��� ��!a�e��x�Hd����}�,�����'*��t��V8V�s��c5��F|�T���s���I35ۢPנ��>����t�1&�t��꒢3�ؾj��������]�z:�Q��X��$�q����Ψ1WUf�F=�Q����CAR��Z��27_Ѐ�}zt���l���>A�W��2^*-��8ȩ�d�*�<8�]�H���3)�2U�$�4K�z �u8E
4F�I`�>9m�A<<V���Est�R;�]�;3���݊gm9�b�%�̙]*�o��v�ﴤ~���a&H���<͜v΄����H�����Ol8�uQ����2�!����̱�d�����y��g��Z W�D�;5������Y�B���[�@x<���uC���B��%O�n��֐��P�e}�0F�D߽��J�ܰ[����
��tx�����윕�g�Ej8Sl?��%�
\��x<�r�o��߲�I�o�zT�
�bNC���f'�Nx�gDH��-�q�$�������khy>���dR��5��Ҝy}XC6���r�i961�?�Q���bǤ�U��/[�w���q�*&��=�[xB��խړb�t@"
귋T� ��9h�S�PS�G�zN�5�u��vH׵A)w�SS�W��ܺ��3�~��#���!��&i' ��b�:oR�����v].���D�n���i�P�����Z۠b���d ��s������rL*.֘"O;Z�5��FS��>iB�3��bUg���"��ʵ�3���M��k����^{X�P��U��Y��~kWMCn�t6�"J/�5��6�F�D(}0�0$D3$Z�.�_D<IZr�K�������Fk� �!�B	��J�T����[A�A���<����Ҽ�IuTj�u!�F���M����/G���p�ȪSh�:��/x|����(�1o6X��������{�T�W�`o���a�>Gk"�9)���rm��`1^-����bԘ��qV��?�����9�����0'�[Q�v��\nV��ɥE��B=�f���|�̓��:��M����nP�� ��Ƃ�U�������@�lH��3�����I���+��$��������fej���l9 �����܋ᛒ��3����ޜI��oMG��0��ȱek�V ���� 0�M��t�zP����8�Eq;�m��gv�5�y��-U,�OUw�6k��[d�M�d�Z��:������Q����=Me�?G]P-�������w�#m.a.^�c)AX�G�8�y���Xd3r9u�ȝ~ :�ս��3�������Ò�ns@�b�0e�|��V�a?G����1ˤtC�K �ܵ|�~"o^ I�*�l~hI=ʼ�Z��e#u��b�g�!�)A�׾��s����iz���
k�ukn����y�)���IAr~��=J�V���P����R:������7�0ze���~.qf3�#_�وd�����c��ء&�V�GL��xAƄx�wp��D�>r|٠ @S�P��F�1��?�VqP����k�$�}���M]E��D��W|^c�Y��ל#Q��d�a��s�[�����*�\y6��b��K3����M	w�tu�Z��i�3 KdCMѬ���l�}�уE��5A��l0v�3�:��ZA�W��E�r��.�x>lDv����I��@�E��L�_ G�c�72ǳ�@�o� ���3`7�ͩ���5��:�|��9(Vo�q����4�f�#��ύo]X�so��z])�LC
��*r+d�q��L&��@���اO�CmK<l�^�cg/�JK�II0����Y&j�yjq��9��}#��d�V(��ڪ�{�����"$��h��0?7��N��S�%���5�.*��ui��L��� �"1�T��I2g8��� 5pH
����Rr����*N�{a��T���z�V
`w��p���Ţ�D!�c+�5DV�P<�6-,�% ҽ̸к���ұ���|9����fz)@��][�b�ɞ�]P�H� �l�&0N���µ�{�-S؜/�s����ۻ���K�M�o�u�pP�W'�X���(S����i]:^+�ŕszO��#u����k�+�%�,0w:�5^�>�ڇ�!��9�¡��KCD�j��+
W�G
y.�#<�%�8�RA�X\e._�&�+ E&ڲ�8�����vu�#������۶IX�x|{����O�!�ɇZ9L?��B ���$e�bjC-ѓ�6�S�[y�i�ei�讍)�����p[�k�e�6�H�ǚdR��mT�����b!��arum�eS�֩l��.6tʲ�}>�ڼ�(�^�,ޡw?��Md16Ek栯�"�U�+x����p�{_sY!UY!)�¹��Al[�f�,S��3Ju��a$WP/�pb�#�Y*�PkV:��僘ְ0�<E:i�E����z9Q�#����"�;�y !���HɊa�EmY��u]���Ȱ^�q���d�W'�,y�����k��_s�U1Mn��7&�w�iF���DC��o��Yк�GUb��?����u̗�����cF?��Z�,�E�Qj\��g۪�1@�k��߻`@�>*6N�������b���P��}�xG����G��d��T�G�Ƣj��NXSw ����;����������#�}R�ys}��l7���6@�I���I�@̳fsn�$+�͇}��+V��*����5G}�\$�ӱm����޸V�7� >$$�"�9�I�Ԍ�� O�qe�?��ǘ#{D�H}4�����q�ls08E-��Y��;~��2s��W	�~�9TV2W���h@7��	^�?KK�GƘN�!sv�g�8��2�Qp�$�N#��DUW �E�|�[�{Ӛ�b���9��ט=,���$N�st=D��-Ł|5p���颐3ޛh�Wsb��jդ܃�Q�$\Ӽ��ћ6��`�������L����Kx��Dm�u�:+j.�~�2�_u�>R��@�W� _* �×�O��[�,�)*�9�`��hMp�v��D�9�h�����F����;j̣.�#���V�f;@W���T���B7�i��.)�t 8ݱ�cNg����Y1�`.�(6${dO �{�{���H��`�@b�0���X���I�{��u��Qhۼ�G)@t�b#�f��|�d�{AT���(i
�?�ֶ�\�wE9)���s,mk��!|��3/�6�dCۍ�­����v�
p*�>T-Ǖ<��PU��W��4��L��*G�v��n`�x�b�v��_b6f| qyb7������I�VC|���,��F�B8���B��<b��8�SUv�QFDsxv)�AYS_���T�ʒEݢ��ΠG�ۓF@�#�m�j(��l��E�'�`��N�g3���Fr����t!��5����-y�>�|\ ֙T݁p��>�tq����c)π8YrR��� S�?�w�u��l&U�K�A׬C�۵�1�����h��z�u՜��4�
ƀVc$�����R�r(~G�/��NW~w�q�����-�/8(뉫k��N����F	«��W����ݲ��	��������BZ�Ȼ�~�xX}�l�do���>�!��S{�n���KK�4c�
�S�T$�Y�����G�1M����n����9lM�0ߜ��IBϯ�����QT��^����a�8���~|�'ћ���a�.��5�/�N�����i�)]���_�)�
 ?������e��0�����q��+vDUu�g�m�3[��X#�P/�K��3{N�x�7(@R��A���
��"���kJψo��D|�"anv~t���Lj~��j�h}���N��<��}���<�|+�ï��}��_�-+KD0�ɬ,"`3�e�T�hi�!S�K��6�Y�! �]UwiA���	t��d�7���^�a��$#ca�U�Q�o�Z���:�8��Y8#�&_}��Ӄ������=wR&�
���h.N_2���Z�B��CO�0Ĺ�FwM�6q�@��F�3��Ի�����-��~m����M���[B���T��u������E�g�z���X{+;�m<a�v�f����X� �d�CI��*����m4�$���g�7'^X(����k4��iL���9䠳(n���8{٧����ّO���z۔�S~��*�����@�0��� ���l�PN�@���{Qs���^v����*Yd���5.�e�ʉ�H1�N�_Q�^2]��[���U��ed>�_�Cp�ri���a\]Ƶ�H�LoVQ1>�|��\����?|���j%�E���-.LRE7�GMG��8���'�3�Z�]��+9R-�m���L���&<�S2��@4���p5 ��y�+flŖN���~�É3�����q�D�
���K�˾A�g�����\f�$</:�ݦ�N��K���?��]�G����;+!�!���(��v�)`�<�����K�\��p�m���������U�e2���Fxcy���.
1U@�P�)�<��6BT1"GlP�`�q`�W�����2���GS.O�V�~�8�t|D��(K�\�A��:߿�ɦ1�ʹ��hK\�pX�5"�.C"�i*�ʁ�mU?7�	;�|�F8����Y*�k��C�)��W9c���d�r��4JPz�L��4
U���LzU�L�ĭc���e�f�Z���t�����e��N�n����K�}@��f(���Z�aK�׷]�o��
خJ{�j��I_7	���Ǎ,�{�O2�2�B�'����� ��f��R��/�6���|%�if���6XFn�:|W�.��&J����C���'+���NsĎ����2
�dA��ԇ0K�Mf��%���O )�����b9Df���gTȏ�h����~�+~Z:�E����S�5/�He:4b&S�4�,5.���ڠ)>O�Bٍ�)�0^�Y*d����F�Eͻ��|M�-�\��`����n��;c��[���^��U�7߲�<Z o]���aN�0��*<ɂ��4�O=`�U81�y��DE��=~�^��,6YfG�5���U/z�OUҩ��
-��ax< x����XS��2o&�]�r	�jI"��j�Ƨ�_�������~q�+����o�`��,�� <���<�Dkǭ�M�� ����w��,~!a7��� �1%��똑0bN�����'���D�R���������~�x��j�7Xw�SL�u�<���"���)ӿn�))������`M��IN��o�a�%GH3OL��>��S�����;Iow�$(�Ջ�ͼ�bUp+���^�� $�����:q�CE�9!�����r!H�Q�jֹ�C���¹I~���V��lh���*�צd%�N����W\����O'�:�DEO]M�#gv8r�r��_�${���fw���^v�\����'Y2��VG�7.�Y�����X�K���_���rhŽ;�ZK�چ�tbS��)!��_b�@!n�� 
�N�� ���b�[a���"]�:�>�c��.���	R�E��'G(�v)���P�D��>X8�ZϭYḛ�[�J��k�
2o���K��vܕpW2�l��l�|I����Nb�@�X����������nj+�.�}3j:"p�z�=-^�c1���.�оE��фM��]'�x`k<.��k:�xgh�#|�����6�bO7����_�u7a�����	�BC�s�ڪ��!�����|Z7ݮ��p7�9|H�#���*���Ճ��X�g�^��e0a\P��m�ϑ�ɞ:��Q�� �2O6'a��j�G�9�@��˾r���f.8],�7��a��I�H_�zY>1��c^Y����,x]���3��C�z�	��vi'(hѯ�6H?I �>��7��LW��Q�}Q����
�aۥ|�88[�F�U��Qe41��To*f��4oI9H��f9R����>�N|Iͥ��ػ�>b��B�
�o�CƉ�9)f�,B�h����6ecd�2����
�͐+"��VaT�h�����˯��|]���`U���*��x3iڦ��P9���>�L�z�;_8�N�\�<+>5������=�{M,�	+p�D��<�"�D�2��,WL)���{�}�~��.h�B��:���k�(ѐpɐ��f��/>!_&�T:"|�^�@{\$d�ﺱX�y|��6!�!�Ѿ%���q[�B�|J�� ��}ޭGF����]�@�
�kn�ATy�ۚۂ��c�:3f���.X̖b��p����SP���B�\���y�j�ji�sT��3���[�'-b���( u����}>X��/�R��?�u������\�p���i�8���@Y�lyJM�q��H,N%o���*��r��up�w7�̱$��sĳO�KJg �Y���d�ƫ��ٲ���(n�x�]���f)��>���8�P<���<���;�^���͊�"�{��x������q}@A)t�?B5�����bȐ2��&�	
����~��pb�AB��e�n���v����QC���=�FB���M�4xP��M��7T-~
���
ꙁ�<g�^��V��޸]�b%�6�?�=�D���겉M�n,{�RF��v�Y�������%}�Q&��V�5"ϟ�p
� �cAf��>���V�۩ʸ��`S�e*�*{3���jU���O�g�mT��!���H�f��+��I��.�W�3C���fD�*^L8�S���S����"�϶�;LoN0>�;[o��BLf[�x��6����ر?)*���bc��,xC��A�{3���
;wӒANt��X�z4|#�n����w}i��kV'Pm���ܰ�u�Hc��͇]�Ů* ��S��Hr�m6�\%\�]���׎����G�R�oh:��}ڔ�ۣ(Pc+�V�'��7����u�`���C�3���S�M�����V	��h���ϷCX��\l�,�	L��[�������$��UV���Xh-��ڃ�78�Ђ\�������ψ	v�eb/�C^	�ΥWy�	�C#�A|x-65��O,�I��ї䡦�Z�J-�d���glz��{e�,����[�Q��wϐ��^�K�)����&��@4�d����W�H)'���0���m�|�ܖ�IN���%T��R:`HRi^ ���-V)�-�,���ҥx�k�J׼e�bHM5�mο�)x?9�����h��jŵ��JV����p�ʪ��HI�谔���spzT.<8�����o��f��r�,���\����)Z�E�ֳ�zA���}��x���5[˓�>�e/n��"����U�����[}Ɋ��%�֯w1${�j�zC_X�=��z,���1?E������AZ��$��R�tm�~}m�>��S���+5)���$�����DӬϟ+�����]͠�aۜ1K�H�����ZpӉe��Ɲ�������^�Բ�E��ZU��~��ek�VMP�j� �8�b>�7̌�"������~��R���t��Ӡj�?.>L��џ�cް63�=pLg�m���r�{��6�=�4/reT헡�ٗ4�T+�5p{ہ��b�u��dϸ���f~���B��N/gI�8k-\���i�~�͔/4ϓuU�rV7_m��t+r9��^��sE{Mz��KR��b���8�-,�`���#��3f���
P�/M�pw�8�O;��r>I2�M۩�}1C�n\
fgxs_mH
��@b�4<'�^�A`�"��f�LۥydtJ0�[|AH��F[�T[�z�G���X�jq/�PD^ki�;/�����m8�>`���V�����eK�SI�,_y��ˑY�Qt-Ԩ�WJ�ٯP�F��=z��RA��PE��h���W�;`��^+�>�gS�*�ȣͅ�_=��ߩ/ߺ�~�п�����G>W��-��jS��������7���Lؿ8�	�P�:����k�M,$���������g�{��L�[�I�gků���Ǿ�.�]��9Ñ��4]�����-��W��ÈQ��e�!��,
�{�i t����;�I�1zD�ߪ11��j3I!��5-nҊ�-�n)���k�,��c��h�[^Q�51�N�J�࿜ʁ��A�Ш�Y�Ft�m�g����;��ѧ-r՞/R㢤+���M��)��o�%řt�ɊH,
�7T����|�%.���ʱ8<L���WY�	�
֢[��Sx������d��z3YI�c����>��߳�~.d���K.UE���0���K�V1 ��~K�bx��|?(�35�	�Y�ė]�FqFi`��.�P�������ګ����к���?e��9����Y!,��CG�0�`�JdΛ�i�����=��pA�e~�y1�f�l�0���f.~c�nK���cL 4E��Nzn���\�es/huj]����M+7��� ��o�Ňx˳]��|U|(�Cu��{�E��@|F�CI���D%�176�,���a�3��h�����d�U���L�#��f �"*�HfoKޔ"���Nӵ���-V`� ̸ө~	k��uމ�{5�bx�3�B3!��o�ߔ�nXRc2��s>}���']��>��{�*�<e��g[�)�Ih�vkqLY�����-t��)��Й�k�lb�PN�W�au�_�&����)�h��pW�ԡ��a�����w��']9�eX������@�n�fE�u�S��`La�^Z��/��^ַ�E�mU �~װ����}�[�[ԁڻ�]�і��\��SM���e`���_wf�
j2)����A���8�;7���+�,f�ٯ�s
��X���u['�5%����%R!��H��K����@�����l��"$�k�hK�����4 �9Tc?xg�X�1�xiJ�-�Z��t����3 ��\! ���md��������w���E^*�OFDEZZN��4��F{��g�XGH��(e����%gÔ}#���Zg>ga��&/���s�)[� �v��'�(�?w�4ާ�D'��v[`CP9lq��l��D�pW��y�}�x���-[̆����x�ಎS�m,�?P��N�3A�RS\M_����6����,� �M@Xã�?q��S?ab�����G�k�Bi��:��p���B(
#��0D@�]�q�8nם�1�ͅfp�;�g�W_<�x����� ��E"����5d\m�M�2EN�/���%�t)#
|4kuŎt�."�������e��M�/
^�U��X�LoUT�T�K+9Χą,����s5�+��d�Q��`[e����8�*m���	��B|ߊO5�*�?���Zm,�n��_�	X.���X��So ]/5�2Ⱦ�sK;!aq*xJN�c�9��{b%���1�-t�CÀ�h��5��p�Z�֭����vwN=��~��ڐ�Ԧ�,V��פ�g2�=|�uX���py:�5crH&�3�,3���^�ѴdX� oT�Y����yF�6H�2,>���^+��	Q�QyWm-81��h�N�E]��k�h�[�߶c������HR"RA)C3�t���F�V�IO��9o�
IN��;��/֙$ߟQ���v�����hm绑7����̋K䘇����ފBE�[�5�Y�����lۣ�é
8�?Qު�c��5���ķ%�)o�id2�;2�<i��nH�'@�ͨ �F�ˀ��,ゑ�c�$x�KU]1���F.��3��-��r&
����왟�]��s�J���4c��-m�g��E._��`w9�V���9ӁC9c (�y�t���Mb��q���Y���#D�v}�&��a�k_c#�a�񼓑^��9�mEm}\�,���/
`�ޖ�cg0xjgA�+f�*�b���f�R�W���Z���-	+��:��A���k�sd��NF��A��L<8%9���1��p�fT��_}&���������I��c\�W�������
���}Dޮ�?b�ª���v�/�4��e�5��gX	u ���Q٤(��q���7_é�x$��N�khxZ�%���t�cw�H�s/ǜ�KS�t�6J.��<�uS��#�n�P������S8t����]���A��	��N��	�`Ƚ3��VB�㎳�O0�v�M%̳��O�/�-��{ͪ͒�zE$�LG>�����9�Ǹ�V��g�N�K���D��¢�RlL��ឳ� �ʈ?�/�i���3 ʋ@�  ���m[l;���]K4�%�߭[}��"�4"�hl�I`of=ʧ1�d�"�][�|;WsX����?�{$�C9I�7�e�n���Ɍ�;rR�@k]!�)�q�8D�b�{$�wA�6�9���#� �������}(J��2�C�`��Od������� �����8LȘ��b��W������?Gi5M]��`?��in�6-��}DP�h|l�\�7F�k�)�U%��U��B<������2�'�;�-��)�5�悚�:���	7s�N�ז"B���̦6M��ݭ�\�^��|��:�B��m���SHI+g����olI�tE7!nX�:��/Ŭ��Vm�	�4R��uB����,}J�X�}�p%�X��M,�͘��$|�����4���C�VpI��>4��bR3a���?�[���@�Q2�;ІE{W8BǠmo^%J9��7mY��Ez�Aig�kTd�q��v�Һx�������{��ȶ��R~n>"Df$���.G����]�T�,�XR1�ÅA�=fLR��'��(vڑ0;��0C7Eѭ�ؙ�p�Ԗ����Z�Q�(���BZ�[�Cj�ZKr>��E����