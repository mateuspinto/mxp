`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13808)
`protect data_block
0USWSUGxovGsyBJteYpEoXRof0O89hb9chjBMJR9k5HCwy6Ehu4IeOug4tncZUaIFr8VS4igThpb
A4mS9H3jZ65cnLkCQaLpVEHhoFZD+VdJ/UWZ0RtEx6QbT+lIwP8/iXjbXFqWT1Pf4NCLUaYJjJyc
V5scHG3vjurQ/J+s9Xa7bzFzpQRxoS8c/nhJXlvHDaTAz0tZkknToBVSt1qKby2jMw1zo3FVa6w4
ddYDKNXVQ9O1msmUlvN7vjbIY9/AvuWtR9fubWnTEmIM48nlW9WX2oTru+HnaVdC72v3hU+qRJHR
rcqy8syrbH42JhRti3eTl9jjxUuU9igAhkmbpP6oRJ/RDNttDpoP9k0K152Gbm5NN0m3qQ/C6Ho6
i2ckx5NCFEbWXCemV2DXZ8Ccf4I7bNA+tROanlRiUYeJDY9FyC0Pxg1AROfX+BvO9glNfbfRnMoH
g/GHplvYgNbMbjNZH0psURCzEbK68ud1kVWI3NB9hU04pwz+okr0aFxbzfpX5c5j4Q3YiBobtPBu
XoP+UT7vJ3GaWxCUDVG7inBr2XZpBiwA/OO2fBPiyFscrdlZn1B1ur36Es2iISv4JRowfiR6w9oo
ePgKK8oiSUfXOEF+WX9V9SeZtC2sZoHxMoDcw7ZK+GY8RrOC6j+VIbsGWbffS+mEcMLSzyIjfoN2
cIeF4V76i15l/L1iFm9D3ZXUNXeoJu9lviyba0f4WyFWu9tWWteJ0+f1eoMO9D9ixmQCLuQf/ssF
a/W5ntutMogZExhrfSPq4XXOEC5Cq0vk/F2fjgb658kzTFcXI0uSWi2vEkr/WzZQlYFdN/Sww96+
dgpNnUr7tXeHUu4QTRHEXiQ/TOY14ZEsX1HJE0p6HT8fp3flZ7QKVX8ddv/7mJxsvSzgeMdFFBP3
UFOl9BdpvLFjDKgnwoPgyXDR7Li6UaHMelSwaS4tOZtc14c0UOR7V7pi2lM5bszR8Bv4ITmkR0A7
9uMNNtfwZjhXn3bnkDWREMLVxwAHkdyUm12H7tla7xh0Fa8IXQEmlJPzUu3HhCxzuSxLf8XZTwPG
2SAniXyTCQMq4XdTrRMuz5sDvX8X5ohcb1kjTrDfB9nv2l8gA0+KUSRyR7d1gK42Lrhq205/LQU4
O6k4FE+S04MduysvoZZWuLhrt4MwOt3mJEZdwWldRLpwX9N1estJJ4hkRgOtNuAIFpGPH0Mnlf5v
5ph7ilDDsdM231CbYFOt+Oq0oWuuDWEPhoG/WyznH0zA7HDQoxPmiH1NwwEVt+Njac+xqEldc2Gn
AzsGxy+6ZSi7uovA7CxjXS73iaeVprUk7MGDDsqFb4fLzuXNWI5EHMC/f8IM1gHWbUJM4vERMWAg
YM8cNv2m7UkPPJp6wxigvPpU7Y5tAMdoFpy9/geDKhD3SGdMdEDJrytot7zKTzb7dFbOBRqsMHKy
e1/INau+5jnn082WkeS0mLy/he8lBvGb8aJ6R4deWdPNWcP4v3P/ZbpaE1tVBOk4Nhwjc43yzYxY
Y9OHXR0Xrq0CxPHEHiBqHCjXhDpxVyBcfv0IESsVphJ7LzZfWVARuIROlO+3b0huEWM0jGH95LrU
e09l/7/cW+dysNoi43+R+we72urCDnsSu42/KhVPjUWj1kMqZiygOvzDb1QWk0JL3GiaA+Tfj0yh
G5kOGY/ZliEXAWnFhCBoc59xi6Ap+JrtkeZFhiVDgN3hTVnvdfzPJbuNoTnHa+qDdfN7d+0el73n
DGoH3PtcRBa15aBPi0PnkJ0r0nXbDY2oRvV+POX0DsvMNfRdwhT087U723C8fIaVW0NB/wODIjsU
T5oVB4i4bXszRqWDYoyKvCpyGzGwWpkKR7CI52W6KKxBntyUlK7ZCFzaPfvkcXaJCSJkx03iioc6
C7zALsUw6TyWpHQSIGzXvo//Jpq1rqln4oaWAuKbrhaPtqru5fFV4GBHrK/UkEiivl34E4UWUffF
Cm4F+8hbAEIeuZ/Z/+1hibaSG54cc8oF2MYRD/kSGOObIz6ZQKQ5B9C/COtGGnp+43ZSt0Sb2KEg
0Bmy8HUB5Mw6rhtTLubXBgVBJaFDe1vH16i4vFZnQ3Yqkc3NY5wEmXKdrCBItOJFzX2ioBtpAEAQ
mCWFxSCcGxbCh3uQjibHiWipmzxflRhvtxQQ981jXgvy4b4qMT6xJq13CcOtGqUcuO0FnCsSofHH
922hVHTMQqQzqimcD4WrUYA294gr8Bmy2QNBR2ge1TZ1MZhX1AmxVFrqayP6uvdjSCaL5fnLbgRA
1DErFv1+N7hMaN+8APfYyoEAuXLRUFATdqqv10qfzc0CcglwYETcaaE0Xyq2L+QEhyPLsh449ySc
OMT93tNSk1Zn9ZXFwDO4f1XSAvDVaqajbuEsTZCYOiKwhEZyjyM8YdIrMW5xTHiUO77TyT5qWNRn
m9Fz7HZIrmKPZ+mc0rNl7KLw4NxakYBsVVJQ+AzLfq47sm8v+OWjjTZs4ha6xjRqDhKBLQwmkTNI
wsyue7d2uPqM4WfGkH9avB7IblKcbgeFwkpvtMGizTX8JXohAW2sIwTrr+ifHOEe5SHSGMRvMrd4
0Vfar7dmFSDtoFetlUN/A4v1Agh/ic+8U9eAIcGR13zdR46ZwLVDc1kBI5M49yC1444T0oSplRy3
co+62HUISUiax3RUcVo1bRXxtUH+vHW7BLxWqSy3hGEry/qgTCUvslyJhEpWWfdmD2ZhrJNxHfTD
ZrnZwL+D6sVHpJuYVup9vm0DRF61L5hYVDIWQQnoN/amrPvJV3q4JpErSw7CW6L3i9D88mGvsLl1
uICzq4DA1qP2xv6BlNQnwIRJPOSwu1y4vpK+4JF4R6d9VBWUxM45bilw91s9NqlClAdea+YTTqTr
wZiQcYNrjtpPKYct9PxnnTzTVrPEZj9XCFIbnug3VcfHlZpMf1En06jI7MZ9xWtK33uiZ6FysOMf
e+Rdme28P7icpLi4juQO/uO+pqxw8jpFxxvEZcldfxc9iubiQ7maeN/PgMb+mAlawO2a4nMQVnV2
giJnhyCxVCYe+1MMwwIQ5aXN5bVJCqQaMOc7C4RvNOFuSUg2qGc3mPn2DOBfdHITyzDwv9m7wPCo
KeK/bx9kxsqvIPJPtIS+T7tRjsrrUJyQ4bJGN8K2HfEqyP6zb/JAOdiwZwUk8nsdRrvGnKgW3aVY
PKnliskY0E5onp1ZuL0mfdtjOP6zHm+f5aHYQgJ3ZAn7qsM1g8G2KtJRpEcaBauWAyAsCoMtooGv
cu5ZswRjgI8GMC5kH/Mxx+rMi8nvliX4PsYaxjDhtKcXsX5Iks7MsSlc/WtHKkjcsJ5tVnOK0CBp
y8fB/ZgX9Yzl6yFy6O+/jCIdgofrskp4d4c/9kN+o9iWv6KAqh7/LPu2t3p59uzE8bpddnCWVKM6
jm4fwTw3Euv2uRocnbW9sz0Lm/E/8HNv7OJxF0q9H9aPM4MsBqr8b+SyJ24f8xfE7UFhRUDxbdkE
DVS3YMiPqJE4CLF+PfXfmBJZ/QYGQ0NX9E6GCYioymx9DHiYXXZGk7AMp8bzRjeHVWuAZTIjnD+u
IYkGO0x9PUx/Ga7Grz7pB7g1Wejpigw5nDBEh3UJJp7dZTNCUYQVSwSc/iialfzop9wKDqv7Lax7
UNOY7Cr/LFWWgC/XpYqU6/LkWslHju9K8d0QVvExMgYDu+hTWhF9g9l5HcYzEPVwYAadkIKfLXDh
u1mpuSq57uj55LAEbJN9pmC39UFmqtlAV498vHzCTtGpoX27Jkc4zZcToUD9INMCe2VHpL+bJ0gY
0V5SQhcxRWlzTNyKvL6TMpzIRXM9xxKL6yYYXdY9CqzhsI4kEYj6rby+HH4AmUL/pOJ5iZ+Blpqm
rcPYI6xgQRI78u25QKXnjHSFnhpJn5WD4fAFtOqem0DPfDCG064hMiw1eT+SvwENTEdIKrl8SB8N
UHaZH+a6YBSk8PYlzfwwNhnxSfkDjKjIqoGKsKHXLrt8PFFdZL3fh/jlI68BRpAAlw9D0IrjlY1F
g+diDLDTp0R7ghQ9l4g3s7EQo9Am04mJumLkOLNyTotL/QaxFpJocfrrYNcDEODaeP1j4OnZ0Zbc
qMa0HGrziMF39uTOqY3jt1J2fpgNp3XUl5uXf5d+zhhkqEai/pjxKmMWXL+4OmyX3hd7W/JaO3zy
Yh29EXs9zShrkM1rR+EKrkS/NcHddeFM3RpzfCD1guNAi/zQc7Rb8B2jXsLXaL8yBlRgwWr8TTnt
6ilMnLbADHiOoMmB7V/o1prW+oHw4aHfcrvRFAlB4EC1Eak4X6Ayz40mB3wc3mSJSdT41WPXTsXG
j2kSeXObsFpDuMUyFpYN9aTpuUWs91Bd74Ntym79RgNLOFzIWRFY2qdSGHZMn7ce9YWsrmtHsarP
zfE5yGQSXZsBM799a+/JsfipiZT9sazHqgfLbgYshmCNc6tFoLfWM+QMbTj4HE2IaTNNzYQ6FwO6
jEwXX0XXPdkrX/dgsGNUNnyT03QrVyioW5spB12tpNJT1f0hOwFRKH3X+dRZHh3dGH1pw/ocoRJQ
q8HFA1X3F1EAMRYYn2BHOxNpyKtwZ6vHt+q1qlSnvEJGHjvN+e6Uu8SoViG9sZ0qU8+2RQ0gcjRU
Ki7VLQme+Zx35d15bMDdD5/9+wDPsBfg6i7oq0Mj3QPwe9jS29HZ+YXzB6Y3ze/96JqUuTQErL1C
V5myWLOlTU0jdCF0LL+G5UTX9yml18Gj/aLIzLEJa1g600hhGDj8srXz791qAXJE81ift4GIsZH8
AO4u5dcT7GlihQBizG7vmdbFLAzKRGh7oR4p4x6Hlhx1XWu0AfY1huKTIjWBxWJJG044KJgKm9oh
yl57uH77b4xKuTIt+9av7T/FdIC/BFoh18W7j+oYaSjuwmvV+I48WFtah4sK3x5VMYF9UT+DXJc0
MH5Bt5vMIBr+JK+oHdCSMo4FQjiFRQSgI4cYIF+jvO1eIVJVIWR3LFvxJ2ff59ArV+Yjfm8kDlPo
nkYxL97eH86eLiWo7q/NJe2HLw2nwRlJZs5RjPFhjSbq5b9SrevuGPcHD2wzITkEU9inX6y4e1tf
9jzcp7ZVs9AShBiHuI/7eID6SM/4HZUC+79DWPRTnbR6A6BO4zv/gludz46k3EVzBBvgYOMGVs+H
55yHRr9AhRlq5e9DQSZSSNbj2wJmSi8Ni+JGO0700P9XluNuzjxA5a0S2Lc67vqPYsezOp5G1QPy
kF/UHRFYqpYVRZYYiyGlwQeTGcEY2lNnaNvcCkrdm33Pw5yj5zXPBHiu9v1Gh/6kARa5iBi6+w6/
h36+UXawSU34kTnbfyFJQS2ApeNkfYz6te6QhDc/E6hRsE3Vjf1Pq5IK7P2df4qIYhcE0AAeOtV/
ldNa6lYFGm+2NzzxZjP/VpO9SMJ2fVRVlXWoO3R/A9i1TXo/B0ZF9aNi7LZo3KLQsRv0mXelo1tQ
JmZxawd1Z3NWIgLV7qrc3Sw8ZZ8MGZnQ49/ucCDpEWeY8xf9Oju8XRxvR5GxzKoV/HlZANiIOIsg
EEQ2vVYZv4lWChRvO8geA8hT9wMMVpFli9mK1kf2eESv/B9Ok6M5AQcEH8ELqy67ykCVV4E4w8C6
Gy8K4YBb9S6j/gxOOHlmxnrEJhDIOKspgAecAslptj0HPf+fJwHpjITTcr49QT6IcrRVw5cpFz4f
Z6VozG7pRFPwZa6vcoZS0Eo7bQoppfB8XHWGy8sdM1A4Ci+hLEhtYXzYhF8fPzFQc3PzjZEE0Whc
h6Hr/U/X4PYMU5cSrZXj4v8wSsa19qHhNPWZ5KOoYfTPNyLSc8BhSGrGjxSK0BWW8ITyrKbuFbdh
75wGJrojWealluEyp+bQ5m6WkBBmkY+lOvM/3QKmgYJVdCxHM851Rx/8d2aCybAJpQ3c3+Sdi4Wi
QKrN6uR9qTMuyikxnN+/mkj6r11MZtVPD9WTaNrXdAhlNtMp+uQEPIFfVNEAjgzYtrLYyevcJAmR
b77le4UUpT6JtBmjZdyMPn3O2KmNGfEPLWIpqxShwp4aZ2SCXckoRu3K8HPK93yoUIfviTRuCRXw
RUXexVJrhK0tWdpZxvqogVhR51o8RJfmB3MVod33Fe3ZvtOrl9GZpXF6bAZPhBIqmy6GbafyPwmc
eo/E9JbvQ5uicvUNs6zt7Z0QE6D9IyhFNAf8Uv47DVoPzwxXMmdR+yQArQuf0MzSgMgNX6zDIxdB
UfMnaW87UoTe9kx1yY7BleOQ57dgav7iQ6MaixtMboZRg3ZqnQbtuEkskT7Q+hWgjTEKMghTvQO5
dTfbLQwst13TZ0m+4BaxVQlLuBDVi+1uaEeUuaxShkfHyiEsH9o77/kp645sUMmIwRQML++RXqXK
skXvY+raqUOFC64hf7OamDCNiV3CKjxkczYxwWRYHJCVk3qzleNC1tRc0m+YDVSTSnTujDPXoWjt
8z7U7PPl8ZAngF2l6KGk2y2/iSWpI+IMwv0yfB6ElYdXNfIOHHg7l/wAgyr4jiNCNbN93MV0WxP0
jkQDLpFKPwY5Q65CMIuVsMHuEMGzSK7W+9O22+sqD+9nVtiiR/LTMyP07y/8RUIJgnxcUcWXVo63
mCwEJLfT/hEuoI5i6d6X1SZIXT7C4JAC3XGzrx9aVwXs3NooJsbqnY7BsOG8j3rU8iLLNhU2UmcT
5+IHIJpnSXZ/NzToyDV/SvTyuDK8hJwqpcgRpUj2fZ+fiW0aUX1xDGIAxjW9JA/uQitRegWRHgnV
G7Xuy2z/YyoLk1XeGlYeSTlJrRgEg02rSmJGkmWjRCzQQdj7E/GIn+yjbkg+uNEketk2qUDJYKyf
z8m8FZiE0kUxTAwTBqcBoVs4YkTQMYnA6dS99gP732Vl9mp+wqhGREZb6VkOuoe68fB+O6v6ACAY
f+4WvxnzSHa5UDWjF210nd3KEOBrE1mJE2P7/vXNTBn3kkmLAMiT+jqxASDv0aCBXxYP8a89erF2
ro0hQcAstYEDoFItpqxBsoo7bBe9obT8ooOkezvadvuTATGYeJROqpEO6sX4Ekr1v7qwfW3tsHbo
AY5dHLdDIoPKkInRKPC3fNyUetoSXWltGG3P3S9FVgRFbAbL/3jtAAxaBIjIa8OEFKHCIbkR7H8j
ta3M117Th3lHuNBubYLd9Bc6cFU7qVdJb9CuBAW8XEADUdCaKXVO8n+v0QBLuBJuViMMHW+r1QcL
/v8vKorF3kVy2PbCvpoVypr+Lxh9TlCe40S9/QGk4DhwR9lipDl4LVyvdInwl+evUEOx6pVtDV+L
umSCnn82vysj58rw9rhtiK6Bkzzm/MyD6z47LRonxMYa4I+wyc7OsYz2TdxC63MfGaEwVFm9w1NB
h0aqXpD2CgFILxdWgL8sI1E1GlYIex18r7YQZVMJV0s1dzdTX8W/EW6P6w+MgWjvD5jjW0FnPa9r
5BT7a33crfl2QGcFraEK9d6ecn9AQ78DdnVFTyG4kqgkFhFpSaNPLypolZ4gL6dL+WYE4QmIz4yB
+YO6lkH1WGvcaK1evuWcSlUjx1ddp3yaCz0e1rOQezumpjkhhIVFCW710hnOBUgjk3wr/EuYs0bL
jDTn1HY9ZAH7bkFiZ9/AGHV+eJxHq6JMPDQP3FRLaRWLBKdAyIGF/P9Ic9NNVZtb9e4nQBZIL2Qj
3FPiZXIbhNJ57H564BtSKBoj15wsXCzjtKuFKMVi/2pr5SN4icDU22QooDrZjxDziSqG1qHRD0DE
EBKfMXt9Jo3vPZ1yX3WQSsZ3tXgREUw4zvA6osM38OiEBmUVipohvlQSEij1SVeYUx2/uJ4y8qZV
5Tuv3LGr1le7XTeGqyHUh8E5o40MwR+gkRoBrZhbrZmmZW+7JfvuZ7Y6Bge1a6kLvTP8o7yM7c5T
AEE/i7Fc6IWUJHftUNadyDJPxplH0y4S0CWdiStgtF4w58Xi97Kydo4EsdoyfE2oxE7YBCnqYc8f
MkZYY9vpENw2138D9XvcyiIyT5yTZpZnprOIKK9rNmRkaFSqdf1p2VhRGygWo8fqrQxInRSh7Z7y
v8tdv3AN2qmmh6IOks96ydOnu/979rOu337TH8S+Y2U2cehwT5f1sEEU8J4U6k2T1xE3cjT3ZQss
nGwG9nu1IoO66j6qWb5jZ0JlbOIxtsGtuzBjprf7dEuyxFdVJAYQnvr2lkKJHPKCVNeCYw/r5mQX
QUju7ZC0XsTYfTtAlLvnpK00b8gaoi12geo3Lma5U8PbIB30tmA8NvniWcufc+D4YC0AtupCh4dM
Hixb5na1j6hnx8ai0escB0DELrXr7VdEjSeRbv5D9YhI1lLHo2AaoK4Hn6B/U+bEhQqhyh/8VQZj
YWN/iKRJmXKdGlzFimUl2GgA8aokwk4WZDI9uvxf7zzZ04CI34QEWbidEBv9CS6Ub50glBYEjGmN
i8/ldk+2n51dwQPcCTY3SN2H4JLk2PFumbe+CAzYH9+cPFmNPA+uqvO7P5BB3nzRhHBk1hYQKRlG
1VIrhxKR9YayJHgS06gF/thpfJEDnjzYWlEmBscfjEpDp97yppezcbPSa86Nvtgi2nco+AQmfDCg
p99a65ja8VsCi7wvOxqmH2prq6RYeqcv1irB847Efny187k1skSnsEyZyTDRhjTt6Hqj7116T5cy
gw86pCXTfwwOrgW7o04rB3N7986yh2kZdPPkDbDzX/VtTjpz0/TLjsOZuKSTJWVe4AJWR21Q25P9
TO6gj/jOyDtYAuEjAWxr4dZNFK6icKNIIqc9Lrqk9gth1sSQQVQ66CgCsJvHoBpoOGafyZ/32bgX
n/ktD7GOezVWr6EbWxFvX2cYI5zmqG0l9Lu/GK2ytD0se3N7Ifjz/7QFme5mxVhoYfKf54jNE0hy
9dyy7MInh8UOE17/JCU4RJNp4DIq8UnKejgouEnayTzUWBqj8UtLNG/x/RGpv8pjFYf5vpgXK7MA
9JCxY8FRcbmADAW/dLmCjZwrKLCWzKIW6nJiImuN8VPsTau5fsGOzZmK2vZG4/GcRKgjdco26any
SgzQcfACEwUZgWgZ/6S9tb4teVDUAWkw/XHLaC7XSs7IUKkxh4MZPqI27mQQfngYxYKPqqPN/7zV
SbcKryPe7JLWRXlu2R1xFpoeNS1bmGAbyk6QC/+pRfrSU+a5TrOg/dyjarRwLeTqC2voS5zyFrIR
+s6aPFAoNSuIXev6j+oiUUXvUSQYEV6fRyWoa5fPnMuNojUjWOWS6rAIFE9tQAJWSz1WELx/Caa/
C9RMMjaWaNdVNnDTlvRwxNEtvXdO0423YVsoEd+DvFjYPthjU1QY4hpDFcSW1iqROhgI+KmZ4r17
MQ2tewUUIi9jCfY/PbNAnqNtSEj8Z0mfYjzTzSWrx/2ZSVezkPywjl84LH754WD0VoJiZhqfvgxh
IqAmBt4G2VUCQFgauUMJtrqMepKUq++yGssSSuyrkKnX8808x7RlD74cy3YExvI3ZCxzEa0Hhl+R
9l0rtwzHjMt3eM7HI5D0mJj1W/0JbADuQmnDsWAZoovBPd/i15QwUVpRWhb6Evvvx1sjvUYBeAZp
+aUoQk4+lfsPw0AQzLGBVkTQScgprIetTWwV+r3Aywj1hgfNRXB9EiWcrwJMAOt5Nbqsv6BGIxuU
m3iQNW9MBy6ZelwsPWlEYabalxyaLKN3+cBkHG9+4qwuHZAGph9eZHRN/6DO/cjbRRHMW8l90ni+
Iqd5YZ0bE1wHz/GX/vtiXTbzD679vZar+61jOCTBliDWsW98+wC2vWRue/IMdSpp8pB1hBIDIWoC
W00OtY+Cu27g2EQmev1ztfSE/U/TyM7njPfWgsjcQmtUI2Ubd7TJGXNU+gdoz2DrjYlXbNdXSVoS
PlsbVT1gG3mgtN9eR/DD5ZkOtl9YzWZnhn8yEvB0tf1J/Iy5ViHoYQyQRn3zhGIaCGpMK1EKe0Do
9LpMDcTiEunMEVqhNtxGxVb03/GtAlocNPCgQ/z/DkZ17SoPF1JGWbCMLsReMSC6veQlzgPH+MSU
e2+gY3jAW96M5jZdj3ckHE9v6WWaim2iEDFXX03WWL6YNrgMTBMmKz28THzlVwVaMQRmY3DpvRio
vDmH9zXQGmR7/knkqyU90KNxt3WMDTAkEN3THXZX76MpMOElzLBmBM7TirQrhgC+GbWoTDzyD81b
CpW07R2KH7V3yRjegn5v6hNqqi5IEp6+X16Zly37G97Lr7VkAH+8JiJBhxZx7wNORWDmhMBdIqRH
Ghwaw7zcRFSM1cQxeu05rhM3/Dwi2XtjZJiRLPe+e23OGPq/T126Cax6HdvYwYG5bwRWy5iZwFaK
GTAuZWAO0Y635lSMofkygAI3BFsgWxcyqQuE72AiDufWDHGMwa4O4N3ucEasa6CSkkGUk9fpZDSv
bT5styBoXF9Th0Ghf2Z9dttruqyzZ0wutmeBqBpz0WHacVpPDP0uprPQDwzkKBqdlRUk6NUYQuW0
RXqcFFUTE15WRwc0u7VMXiz6QHXo5roGbhGsCk1gXtKmzU4rKs1/HUolTaNMA72w0Qjr77TKDxBs
SBX6jcNs1oblBEzQDkVlMWyZULbz67lUSIgeSdXpSxG8PqukzfskjuxolH7uUUljivg3gnsnH2xd
+a20D8w5vdNEfDkkSwNy3dp3st8HVruiUw6Gb1ALNWW2nvYk0FCZwh9pSe2QOcUrhpsvGU/IwuB0
OZbWH8RBto2ABs84Va+1jVP5sW4bPzhav8iXMC0Bk1ofr1OD7TMo3DWxnfuFULH0cXeMhwSOy9kC
W7iwCx+VXfZQ1UHOlpVjO3RJmdjQmeS29Yx/dOcyD1PlmJCqn+1OpJ6nZnHBGuLNOZWu4mogzJri
wZF6FIBWfxNXJb5TGIwNHMoeNg9UU8Ijmi/BD2w3TH4rFD0eUkMXGxlNTW5mrT55f4ZnQq/gqf6Y
hwtdJKMCD4dTmhbeqsNs2gRo3E1lcplRb42S7CIVZpSrBZlZhhaIlDiNGW0+Xa9028F9pLFrBOI8
O1oOFo5simVcUhcK+uKyziyDnR3Cwf3pUXv5PCKYYCicav5Rdc1nc+QrWvMDJHRKqjnrDugZnE72
gSDsqc1OAg7eiFy50ZkBH1wO693wG9teTlUeWxxSbEiIzY1g48ijfyJgFjYjvwsDiKuMwLp7qbWn
8tOA8/ubsdrRJfD5SExXnEjIkMiZp7ZVS4T6JaTSKf+W4UE4Ulh87Evi2/t8unP7kbN1IYTWUdAB
W/kUmbDtol82GkQ303OSf5SsXUcr6XS2UuiuX4MFPyd4HOvqaBPC+rajC708eXw4XJuFkTdIxzrT
IY2G/2mokTfBbstw6uIncRuypV7jAmp5YUz2EZoXHY29jpLEyKd+OTpr+iTTUax5vRCiZScTszw2
5U6jCIL4amECunxWu7th71/7iOWEz4WJM5mQ+S1xCdue4rLho1tK6lGxFBuv/tt4osnvYRmGXegy
KYEeUJ07v7jAGwPAPt94utJkB5J3hxnPkkJbitT4lijS+u6K/DEu91HOGqnABPE05mkbeP1pcSUE
gPXMQ5w+i4W3PHkwan8IPu2hQ4qSHZtD/7/V+v/l9KelO1azQOybmL08AA92vtZxYmuHhHKjyFeC
/orDzkfPNa41ySZGpPxHtoiVn0KsEwAa8Dmhy6myB5V51hRr5lQfU78bdFMTxkstU/8R1i7cGiF1
Hf5rActcP2kaTaouOIskKSBIC/Jv/lj1YJZyI+VxVfkCByeGf+CC3a7nnxuz0CN3lZi5nDMaxtJB
bl8gFNlx9BOExNB7otHC0DWWohHoASWgejS0kRmw5E7/q2gVR4usKUFFq2YjDtv3hpVRqupqpMuJ
msbLO//SazqLM06+Sr2cZvoev79DeDRaqOLoTAYK0kmB+zZiOBCjIBqxaT0AJ+m8v+VZntLeVCIx
725GeQC+EfA9e640Pxpw/WgedE2byGgqU4wTmGxHSksogoGFmpgX9At+EKKL9l35E0kHhOlHLalx
Afj3gFeUBJf3ZqIGJU6b+SD/Nilbt/jxnQyqxmaAgGf/RVhSoTKDanGBNnmlQbNnUNYBO9336g7n
kj2qgpJG+z0scnD7qQKvBAjKYu9vqV4U1Lyzqmx7PR3qOPAnoiEspXXpRhHoJLslhoIDYjtXUruv
gGWfDIemfWhXNJdsTD5zlhBE/cGJ0hr0k0B31zp+3CiR6EzcG+MC5spuIvNohyJAt0AOAq0TyKZ0
MznSSwoZG5u4AhqbDI1lrtOj7bTKh9ftL0Otv8PlyHcpFrzKXzk1v2LxLeLA+NaMyV4+IFKU0sm0
NP1xzZ/u7Um3tni1OT2kRU6bQrPmnqIjbz2u6oU5mvm02rvUJP7jS7JiCxqG+0j12qk94WNq+qT5
96lgGEiFrV33xicT4tCKXskb+A4G19B4sR0UixGkRfjkixQS9AAnzaoD0Kb0fAj1m+wQ6FsSQYvv
Iusqhgd4QxTaJUXUE4AaJYv4wTdbnF7dvSoZxMsqha48ZZ5bTvNe/15f/tsapUVYrSsb3wGBtc2c
M7rB9X3k12aaZ1cxAhRahyZxAuyzf8YSyiJ2f1rxqN1El6Q4UIqBzvAFgm4aI327H0mAhoO6vGSF
D3ZWxNiaQAe+VXcAM4OO+eN4eLjc3/fv4Fzpd+Sj4I3KbqWuM3Js3N+xM3yx4K/p/jx6bLjYIz+w
2fAZ6uGTwrUzktIaOluMQoxcV1APi0XIhIDeGtD4mA90+4HLK0/Y34gdBIjrEo/W61GQXNPDeZWb
n+gJmI0lFpkkNZkW4ZLJa4eN7oYT5DL1D3rbzyhU0SNOZiusyHAmywnks0w8kIZMDvfIFZU0Y3TK
fxARefSDaMPfcBqNBkLehu0+j8L66D9SjkyjwnKrsFrsxJOb633mVxfY9j+AQz4FLxsv0wmpUCSU
TCjmKl/fxEW9UOm/le6lK3fI/lJXCUxOquNvnwjbQLBA51iVDRCRELXROstKSh59xi15Zy2oYq4b
6PSYPh4yZ33TpqSTvhKUePuGyN+bf3jiQBjZCt88S4MyWs7bnefV0jnPl+UZ9MqruQxbR1gjE3i2
htI7z24Ro6kI2W8QxtCllXbkrXm1pu8CzI21TK93M/3v60iQOeuwwbGLLASyxAcAKrEKE5igylkr
q2PTTFrD0ob9cKhAEL27W6SXhwdpqg3hx05Ea4bpmtPg6NWwkz+roXMn4S+qGwxoicTD7DBrfTzD
Yp/Dq9N6MkbamxvwnnLKtJtW3zdeBtuXqxUJQn9Sul7EegCnyEfnOYoufTSH2Dhte1+glDry79sK
Jt+pqpda6e4eDWwlSsfz8s4c0/kZO0fZS1/1C+pbt/H9q0B80rusxEMMi6NfsTgIugzBIiYJmGU+
dx/9M+5I1nCGrobvPtXfZOFHRLBd+wc2jeZN7faWJGO7glKcVaKkpLDsufuJhnc88RSlDny7suPq
UFtcuQojUcqSPSnaNVoaUoZCZhGhhxCEmvHwg+nhZpQgqZ1IXS6Ey4/+JgVHqce/pxTMc/r59rju
onsa1OsBfKPQUYj4HXvtIUmOdFhbZKtPNxOQgg39+35S4Ffpdns1myhlKI8kC7DOZraawcC0B4+x
A5+IwyXXDIDMvDDT1qpERg6X55l0CZvO1MEOUIgmJuopnjPjuLSPWTZuW4xyVQAci+vaipup33Tf
QgQxKeZlUmHl0wheRtnYtePEOjewWXsDq0JmbvQ8Hte/1bdfKfFIsDVcQ0DEE0uuFG0glPwPYqjk
6cMWg+1lADIlbd8XdFhQ1joL15WaPKFjE0HjeMeg1jGAMkTvx4Jszl9Fl1PEDi3VDDUWIj17zn54
Byr3EfrgvTAQmqrn5QDLp6pkEc4+GvkiDnOnB1epcCJa1Jm0z6LtOJyXEI0CAOKicM+ZPH9krxT7
Ss3BX05Pxrvd3KpuxCnLJAxPV/AgfSbM1rb8h6zJD/1jLlVrTjO85Fr8ArMtGvMRQK5oG/nwbOho
qLf9N7DgdZwlQ5LriDXG05GKptGR651DfxD+thdybEurxF3+BbbA9jLIqgkckpV3NCmTG1a4+SsZ
/KEs+kWw8WjX1KZoG32s3PZ7SjHKStX5VzeytCIUR70ChhFhmOxvJi2kjB9fRdZOGimCBwp/eKOF
ZYgLOuwpN6CpwQ3f4WWTy8sdwR+1Yr7P2DOTMJU5Y7PkXE+AKiktkrR6Fl/Fr22zqDtTZi3CXpVw
VMYvOAfOfB59OV5cCo4Y3uz3ItXeBDZvl3IShKo7kRTwkvqhyJ/SSrNeiq+uxw/YniHlZngg1tiK
s5V6SWEJmarY9QayrCVEFxdpSF0tUJ9YhQHPOy6VT4ua9Odp2B9L1UPZR5Sd7Xlc+VonZiTvT6y2
S3iwB24WWnYOShw7FlF6Y8dnbUfVCzv+Qr6EgFYVYjMmveJO/wMR1ScM0Kqsa/Sy5l1B7bga0EgN
zN7sPOD8bmhPtkCSKy87qMvEbA/XJ31QECBbnzXfKe02E3kDJMQErAgzoiV1NVum8XH3ICSEVdEm
bmdBFfd0iLZygoAs1a6oKS8mu37ET+273cZmzD/MdSzw7Se0iHHZNvJj1UfRMbx10379dNUi8PCO
rhUZk8XiAQLl99ehqGdKAlj0xCaIjgPVlIjhjsyPuN9Qyu0D94XLOnklcQkwBIGwU4LwyD7EGK0r
P1L0PcTJaXkMa21s88a4GlmdkQTMfKNwBtnaC3aZtRgL/f7k48S1RxL74P9kjQSkZf9I9+s8VaXJ
oIX3WhWJ1bb3fbxE+qCR5qAgbnhT99x5/8IpQwVJdo9sS63fKj8NkWjNxpy0mcWCcan1FfV3uEim
NvRFRalUYtiudCYbRXLctKS/EY+XrdlWlXx80YT8iZRCynZwgRJgXHI3IXNb7xUqrqigk1p24x+N
9YcsYmtUDV+5QTFsngKA4JQts/RWGWGOwJxgkHhzCWQh8O8rr9OLrF0SxHpfqNsmggAuAcUiIA4v
VpP3SnwwT8FlsnVw0KGEjhVaCxAcBLAGMiBTrnEtbROmp7y687MQ0aIqnP/PJR6BoCiMy6sSiuuY
xhbga7/CwUJUxy6UNtusicqJ1xALF9S0Zdc/kVzX5dz6pK7panIbs4N4+kk50WIsQLqAi4PwbfLx
rJxGJXEFP6ey8cjbqoD9Tf6D/zGd3TkPB1NOMHm1W+iWE7el599h9I6Ec1r0AJF5DPnr8ZxkzyKf
3uwkJ1YMd/byy6g/k8xV1kpDA0fD5QTEpagBSmymEcNUKBdMIFRTVk+OxjOQO1wO57z55eFqrsWe
0VpzGwP/djk28yaShznfk3AyRhyIxHwUDMPtxp82uR8NeLQW10Dm4XuxKFncCYhtSbtJYocVCHue
3MXExpnQiQNg4AYn/vRHoULtGsRX5psT0D9wyFF3XfyQlK8ZBCtqRMdNVkkPScxqhSvTl6K6rMf8
j0ieh/af1kNz491p0As7BclA/TnACI3knCH1xfwnv75CFguwEnSMQ3tEV8nrNrUAV42fRHY+ql8z
kjmAdx6VdMctmZwuIpLCK2k7qNNsndOnT4A5yzbRfZSU9022ImTPix4Dk5+ZY0HJEf2IENamcqs2
4fsCSG7uB9ZWJ6zBJWg4WhX5U6DBnu50oQkbrwdFRJelH0NUVccos9vCHpJGfhwWMZ4emrohFE8b
RLCjI3OljTXZdRARCdp5Y7Bx4nTCqyga0qbkvHwFVTuahVmuKP/rxALBroGQhbkrW1I1zJn09mFA
MwwRyQD/43LuTRV2Bx5sDiKa3DGFQJrXT2D56+HVApdIuRaSR+/PObk0S62hu3Sb+iO1YfA+vsJZ
+cKW5BMFnu/M4rKudgFXWycQlU1ybr7UUmkNb5+2+jj4llWcEFtU7VGOAscE+RgBA9HnKbXVZHTs
1N5QCfoephu1gZhrTBxH0X3oSPyl8Flj4DOxf8LNYyy4e+EN4n64ZzAAmOJMyisrIG3tZnK+j9fp
u/seJfJqgHO1PxqZSvc3xpxMACFE0uNqZjlD+ubmZ0JzevEDgGYcJBzt1mplMHZHqGpDr2MYvdPd
7wT+BBPfNdPG6U4i8WAP7k7994RfiFERjO8cX8EPcbVD/lAHICoMrHtyL6H+vglsIGdClStyC0QH
oYzhGN2WGkrAL4alMopmQ9U8atl58fOK59+e1qU/edZbY6UinhHUKKQID2D1rckDRK1M9kamYxcz
UaPA+mYK8uPu9by2vzWsVDPgkkkN2JeHW/fMA2aoE3Khu6vHyUji54HM5ujei2QY34WCJ4m16+mD
PtuviGXJ0JUK3FbURISbFj/YZl2mBT56Yc1UxEEj3RNJpnJwKSx1fGWlRX5M2iyz6Pqt32Ei607P
Wz6PLe+ltOhFDCi6hLos3CF6aeDnFJP7moDlfFAKZUENllLe076GioyHRkuKU3KMiwZ9CLzNd+jz
ipweMAEb6OoKVGRjJqUjD0asFDZ19bgpN8rK3WekLzxF7L/X6ujUN7jZJsamJGevvlQbt48AfcFy
qvYD7m83yVSKfvsEglcj4DpWr/TT/LkqBP0fQ6NtXTKvzuC/mY0hUegvkct5vXlg48aaML3sEBpz
dkpNL91hBS+sxvA/Wbg1jqXD45NpoWJumrRsEnqWmPZ691Y2Pfts6DbhCj5iI9/RrZLU+bRFU3XH
DVH2m8YTHXd0G4Vz1WylZ3V+7fI08Aa5o0qPeXYnRC9+DVCjIqy00FiFJo4LeSyVJhpKl7vEW9w2
V/eB+axKY2I/WfH20UoUNsU2LTG4TPSuQdzney1A/qt5JrvAX+pUH1lP+z++vePvL6Uo2HWrtNaM
Vw88N1YRRQk4kXvpnv40CXYIFUJCcVEesMBtiKn3sEJHxhICyf1Ldzh1DDzMeuvlYLX7dmHP4WYY
fX/ltmYEvW5C3Y22FkkAGM5UxV4GSqItnA6yLzLJmRVo6JjxSbmQHuYs+OybUSRJyKBo4ySl9n2Y
pWUFpKYdsH21yEsviFxp6eQ5Hqsh3RqbKxt6DA8TXWQYPmZKFWt98GMKwJ+Ru3BodtV+APcQ1rDI
LhgeMR3R9EveojYtWqV4QlWLYpGuudBYYm8LBWBS7XwabUVJgnDyK9z5+HoyD9pWGPVL3Vg92WSe
bNrTdcuzOO9upgoMHpSqRUz3KXzm2Y2QaeFoMnip8fsg7lCEd1ZdHQ0MjDRIUzA9rcwCki9tW4WN
QcNV1KMojrbHkEnbg3SP50cxrsortENh2mAwUi9F5z0rEfIfmoHq/bLcn6a4a/nrjZmwo2OOdwvM
0rT4GKbfILLUuV72WVr+h8sHOsPQtXIBwHCQzmG+5BXXw2SrcSzDHmcoV8blE+etk7B/yyd+EtoY
9i3O1RGBUHEWHvn33Oc5ElgSq2fkKa2wHYBAgVjlnDdxlEV6nxJhw7xSDnhRiGYXwNAfB42bJMc/
tih9MpAzrA4rNoYhLqW39mKI9vQZRUCkT8OzjDl3+vIQd00BBVK6choYeFfwBI5OEc01YAL4fAbL
q1unbR52BUzitg1qTsLmk8vs37EMJw9lben+wCINQlltNmVc5cWQDIFT0yd0jmj7aH4leuZb8ee5
qhlP2OuITie5V7mPOf+x4DzoWZ/hsK5pvIX035CMDlF9lBmL9u+U94NQROAoJoKbjook5Z5aZ1Ub
gbtzWAXQ3fEpXXKuiTRQvGBOmaiu6BkC7rv3H/WRl84aVFoMJJpIKJUR8qyjEvTVc9kB7uIquA7q
09XsTVYcftCpZMBwF9M3HM9YugH5s2lgZouQJDPgymLRLJcexR1qhoX5EcvFpZaiQqRISC4NPfYj
AVDf6ybKLDfYOzZ1zFrhqKHwPAqhFd3KWUyFtJM8mn9iOSA5SqLJG29dsBDMtX5wfIMhGFcms6x0
FvH8lqAQPGRDHrndiuHo7Kqi0ZNdAViTjfsNeEnhNzGjJAFyj16nILWUAuAVpbMvwEomjdE75nBy
CrZTF6uwRI6fDUYhs2SrVbakRhVJjK7M0nfOLpRXHTLVM0oM9wPHPQ447Jjrcr4vHIOSOoVC2aVB
zAhWVgP///YyrvXsHSworb/+pM7z2mCR1W0JwuAcXvJdOZlQMNs5U0MQmRnGzd3k7jqCL+mRQA3j
TNbN3W0t1JFABbz+gHGn/matagPXWM6PVWVOx7OUxWikxRRtsk29+APgvzJ4XMfjD4VYlLnyq12K
9BVIDZYHoTH8VP4xK8aAtyBHt8VAUdeX9KZ7H+XGxpT3H2oqqShLdYMc2VUNz4ta+NgIM+ajePbn
a7J7lDwhoVPiilvGpwmyEEidYs68PcJtQEi2kljruTReAXTdLikq8NMy1u6xgL6zsQTN5e51hxDf
45TyvoUd7RlFu1N0l/kmDEp3x0aKPg5rq58fjHkHyJEY5acegcaHFQdlFFVcOY9lSXm0j+XXbi0v
kfqkAcXIoZxVp6j1JYU=
`protect end_protected
