XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��>r���ู�~E�U3H��,���S����:�cBg?Wċ�V���Jح1�ߜ{��@D5﵆��N=I������%��U��K:� ���i,����Q��HJ�Ck����xdh�_/i���*�М���6�������i�;����5�E�A��Ұ���w�l�T�V�!�A�i���1Gcv"
�&��Ar}z�=��9h�4�Fk�T����k&�7��a~ɾ	�����)��	{]��l���ќ�L�M�V�u�](�9Z2�^�A;��T���[C�e��j�� �L+�]�-睅��%��vK��l(^��0kx*�g�8"���N� zW��ڂ����fTQ-�a�r��^���?���_n�����CL,/
��(�q��5A�#��@��["�$��
^�(U�ݳ@���pT$�����r0{N)ʕ�:Lm�˧[�P�Z:�f"�/�.����+屎�-�*�lCm+��M�Mr*�,PR��R?��_��gk�r����'CG�C����
�N�����Ēލlm�$G&rb"������k�D��)�Cٲp��խ��f�Ʌ[A�� ��Hߨ�A5�М�8)����"zI�w�R2��G�{�6�	"�����%��;��k�#[C������̢���8}$0b���9"<`�v�8@��~�M�pߢ��ѺXQ}�hj��׎�`�^�b�sk�t�e�[�g��^T��g|�Β3��F@�XlxVHYEB     400     1b0�����3,�'��'b_=j
ED���UK'�p���F���\i�u���6�\P&󱜒�!�k��w]�����������>I�1��|#�v5���)�B�½�C9��s�F�/�8C��������+��<�%f�@�iW�4!��INsr���N~�U3��Kaie�^�9wȽ�W���Me�T�xM[� ��᢯O�ݑ���u��C[J����x��.�K�	��G�����!z"Q��O�O�3�n˺�9t���*�B�)%�,�q���Y@#ͱ;�B�?�)�g��+�ag�kX֝�u�u��ą� Y��OG�p(������_=��7@���QA^
���jDX��.���R�CKp���t��Cr7��sJj��e��ux��l�%�/l|��z�.>l{8�k��;��8�L��
��B	?��	XlxVHYEB     400     1b0�K���q��G��.�N"'�ҽ��1t=�Y$�~��:���Au����CS�G����y�&�n_����0d_D�UlX��4��K�1JFNXD�����l�g_E�[��?�@/ؑ^�Ǘ� �� ��8I(\���_�^�����/b�{�E74���Df�d��S�KtDbqɮM���Xֿ�Aݝ�f��d�����q��ͯ �6��I�=�_P�~���5׏�ɹ�!��t�W��)ɢB�ۮ��}�8[��Nh7�U�۶�|��Y�=��שa�\4?s�5L����XH��3�{)"�h��t{=�{�P�J��"�5{��QH�CJ�~�Z�^l˃��Z����%L����wAJ��x~Z���dȉ���<�>|��[��bP��g}�v�vP�J[E</T�v(+l���F��A�|�+�XlxVHYEB     400     130�`l-Ɯn�KEu�-%����(Ӥl�hA��Ƌ�䀼��K���@�n1N+�Kyd�f��
d�E��>��pk�˧��Dx���,�/Gi~@ �������d!��6Ӑ�ҽq*!#[xQ0Ԥ����ܭTo��	 Nz1=�l���\�'�����/��v���\'-�
���Y`c��r����ÞP����&0d�Н�zP-�0��u��9�wÊ����(:4Aؓ����w�_g��mn�k���,��꣨�yA�:A5�f���[�*\*�b0'��m�'��d!�4XlxVHYEB     400     190z��&/�q[��Mu�\�sVp�u�Mu�U������YO2�_㋍���RF /�L�������F�#"��""<e����'�,���I��"N1<���	��FD	1���g���`Ƀ�b5��<����� gE�㜾��Tq�O��dЪ^Q��	8m��� xx"j.�-R�u��x�ru��[��cTMU�b� ���-��/18ŧ�_͏���4��ͣ១Ev_�H�ߥRp�cQ�j��ֻ����q�'�9��$��*9���h��-*R�TTF7���W@�GND���%H�n��h�Jd��&��J~YÒ*>�&+�#sRNL��w�o�~A��WT"�m�Oo�]f�,x�2��Y���^U��>Bs�]M�����g-$�[�$�n�g5A�o���lXlxVHYEB     400     160/�_��A�T�]����C�F��)|���k�=�F�XnFf���"�`� ����P�8_W�:gI?2�g��0�&!��hP�|���Q�o5=j��\�{�O+�O�.��"�54Z��}��X�3S��ȩe��:����XW5�]����F��k��s�N�f��<W�v�����$u�N�|��H8�+�z���B�d��3��g���<$�/c�h��+6з�#^|^�ݢ�l8nN��JD$2��~���ְn���W��g-VTE@�{�,>&��5҂\Ò��}�&���Dv	y�)9���(0��~~ѯ$�F��
�	�K
ؙ d��Ă��U�?X��+�ܚ�|��`XlxVHYEB     400     1b01�!�O�K��&1��Gkٵo4UG_Ğu�4�D�V��Zd���o���M�C�Ut�L-��p�%~�4njt�)�y�Ɠ��/=H���=>w����~���̷��{�Y=��u}Ez*B�ӡ�Z4�-˸�.3�H��E88��4=#+ �M��Fd��u>�z":� ٣YkqSC����r�+@�Q��z(_R��>@0��q��<B8���޺S��M��CT<M���0PgX�	tC���Yp�?�#�V5�tc���o���L� ���\ �@��e]��/[�; ⾘3��)����
�"b��6�����K�0<d,��u7<�͒�?�#�~W�P:}��?���L�N^ѓ�W���6�x�55��1=�Jd9qm�h4�I�>];}Umz�hb�.ϯ�������iO�^D��T/p@XlxVHYEB     400     160}��Z@�n;���gޖ�80�� :5�a�OgCj�f�e��z�#����O�`�a���L����OWf_�7�Qvm7x66g�jw^�m��[%fuz2�G��M��-����W6ES.*B(�A��s���k� |S�'6Xy�K�$��J�ڐ�;���ܸ4yloO�����ZB��1��E�xt�M�E�fN�>��N5����r^΅T�1r�Q5kO��d=T���5o`s��	GX�I�w�&P7��-Ra�3�Sg�o٣�{�^Իm5e'(C�AC`x֚��жcfW��?��҃`5�E$Tu�\]�y9^�J�����t����V/�ġݠ�ߋf���ȾXlxVHYEB     400     120:Lཇ�(��U�j��8ǔ}.n;c��6J|�?�X����u�"{ !,�ġ����y?�l1��i�:��p�����aWCOA��\"�[M��{�	Q��B��8�먽6���+�d�z�&0Yi�Ӹ�&)�nF�e�����Nx�x쬍ɊH�d&��,��]��I���?&/[%UX�'ᗑ��1ڟ����	!g�\TZ��)���a��%A6����ZI�Ӻqk�2<Ÿ�4��½���9c���L7*�Od?�55�~D�1�n����N%��|XlxVHYEB     400     190"�<�Z��M��ww�B�;gL_�0J%���4�u��.`������S�c�p����6A}��	�%��JA-6K�p��� ᫇Q�52������`S�K������S�r͙T�*:.Dv=��Ά���%1<���ꗃ0���ӊ`�4Vh]9����+L�V��\��N��ͣ��H����pZ���K�o8HZ�-�f������V��w-�"��4�ĝ�S��P�޸Z���b��7R�&	��[�۾CBoa�K�T.�\��8"!�^�[z�/;6�]�u�,�_	��ຨ)+!��_h�c��^�8��	��F��n)a�	��?�s�N!n��XDHA4�I`��4B�2��nCP��d�C]������׉ߚ��,G@ul�ơ?�g�m�d��XlxVHYEB     400     140�L�(Nw��ɧi*���20eu��#'�������`�&Dk�d�"�8:? NS�{�
�s��P���a(@�\	�H�co�խ�t��~�-D��8]���Y��	P�3�&E��.�逨¤��L�>�����B=�ܟ�B7	�=6�Ұ<O�����(���M�_�L��R���1$wkT�R�?v�OV&bK`��қ�G�k/���N��G[Y� E_��U<��vgU���~�#^�M����O�g�����u�]������o~���`�BB��z駏=��&�̢R��+Wm�f��`DcP'4 �U�8+-[���XlxVHYEB     400     160���jס+$	�u�e�B�A�1��Ƹ�����v���Y�?o.0F)Q��;��G��X7�A֖@��!qu�]͜�ZϚu�3���	$$㐮` uI�mc{���F�)��b�^��ҿ6�x?Vm��D[SH� v�ζ�N�E�J�c�R����Q���qzY�W��3��J�n��>������˃:Ȉ���W�}�A�(!��gr��[?��e��R������Sge�b�w�)��-{M�0��O�خ9棿���Q(�!�dΔԍ��'��!U<;�;��J�I�aXf<��Yc�2w�ˠKk>��r5�t[�{%�ۑ����K=��{�^XlxVHYEB     21a     100�a��n�B���yR)��� I�8\Vg���0�A���-&cYZ�4E.W�C�b�9l�ٺZ��t����&s�34�Z�l$$�g��V�ҚW����Q���3���o��=Nb����z��������M7'���Z,$��
��@$y�t�i��W(^:��_u�v&��sO���cyv�6�C��d0��2T X����E\(�&oF��h������A���Os́7�\��o�r���;n��تÔe��?��m������