`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3168)
`protect data_block
WN93ustRabOsu4ajm/QGHr8/un2TolQkvjoh2y/yAB0xwsirjCbdKhnRC6tmrgo36vTBXoRR4S3R
CG6xIpza1vv/oZS/MIAEFhAqGBvc5x3aTK6XCi4ggQjN1rqIsjROuqDZsQkrRnySXa44Ij0dt2lD
0Xov+kmsWDTtF6m0sxfEfWiucZecqeM08ipIAGanTxjakD0ZFy0ybJzWrptl+wI7XOo1BSqV+n7x
ffA2nAVV2NsjodcAWzFpjAZ0vhwAn4Mr9M1MvlmxTRczhZOfSFSZ/w343r3rAYf4vDbB5Q9a7E6b
hAczYhmUB31ttKjcG22TJRFBtf3IzD1pIXLEYUI4M/k4RYkAxXfqMH4MEySZ0lUYF+zES9jJYiu/
kVTcRtdTbsiQDGLOq+fL0pAvCj2bA3L2jPVuTcR9AquKDkva4m+uIc54R2OtYYlMVommCTbm/1b2
RJMmk8XofxRkZlot274SnHIV+Fe4yYuRzD9DvTJQgpyi9qIyWWQXAGRAedLoN99iS34cfaeORFCD
iWZPV5DvdIsUR/6lg1STdutX8adxtx9EHf/wZNjZWR+SFsXe55uy54twIXXi5PuwTC8Eb2dPsdWs
AYVOjAPJGsiAWt2FrWIBLNQXJUtIhFYZOdso7shBQ3vW9CdRES2mknT0HxbKjUM6yokb6XrLJWaV
P4LvmgG4PBwJ4sn6SJ29juxOSxq3a0neIWx6EUFdGZrUhZ2r+PuOsUKYsvPztYTxWHwfiUfs1num
LbVSyd3zFnoQJqxgMbmKi/w6Z45LldZieNOuPI2fa8PL9VbztTN3x3fuGzkAfC/4tM3Rs2JKlIog
x66MZrR7c3DyGwNy9v7Tnuqg0eyXteiT8dMsEplPaeKy/1f3vWpRBwq1ifbezGP0o/7PVKWZaiWk
8pnQvvIQPmXvUbDSGaW0Tw8EFbLcGiWtYsZt+IQnXQ1eaUsQ5yekUpBPli5HGPtsjgDmQXTDn+Xp
F7EquDaneu8EGoA/OqXw1pFygedoe36jWDOA00y/kKw6jEK0QqilHHFUcPEp8yE9xGP5rLdBVS+h
b2FBDddoCvlP6x5GliGegFOr/PtHlo+tzWkzmFG2RTkfHNQpYs+JkbBBnnrHGpck/P4SvtB7XETt
Qi8LTgzm5KO7TJUAmYSJX8Gyhx5YM0F3A99frK0/bGybeXCQcUi0hWyP5bngt6gXymB6x53rczuo
eTMzTwFu9V9A471asKyXKwdPvH8ffjr8UjK9boulK7gZLViAR/oUnUWO1+f393g3jHOlWXMG0For
FRQG3Ls41r2nGgLNQ7ZO8B1O0s0NFDzcJQXNWCHRVcYwUDv0hsM3OMrKCF39A946xl0lZkI5NLql
peL0jW3WAJB63eZWeeIxclHz/7Y+4/wc6WN2+cgIz3tLvUT+YoJhvtg6ZtHXd5n179+jEOXqoA1/
vJTPfXmuOFWHUr2DGLC6W1VFeoPqSEGwVQNJ75RwQFrnw2hHBsup7aZcDvnncQzC/wKf2LYBaYFg
q0Xv7E/dlg2h4GpqqE+/5xbdzAuWVjB1kUPNHL2vGqnnsFtAViVeFYyJ8jr+TM4FvUVQyMKA2tIL
7PRlNcLGHBmQ6OOSvuFXejbL24/BKxloY/+Zw2Z1gO5GiJYboRWb9DksKi8009a9fJp25rGqyAmu
07pUXj5ynrxnxBzTiiHMWXE93MMDaq9yq99txr6k+nJ05kwCSxyisnDR4Po+CNOzcmUTrCZrEbdB
NrXsEBQkKl+/J815qpjEMolVxF4gTlXKrknfwb2eXib2258wvjcinCxWZWigcLKZJ9KFKULYQmEa
HWJVNIgHAK/8H7auLH1YLdpW0iHlvzKgkzUM4yLTd/YsQA4/oh/rA9I6aJIAhntOh/aYkS0OJNwP
8Hk6f/RTgqDq9tGfHO5OmShk1cVk/LNJinFpHHaZbmioQrQ92X7na/m1ANsNdVltBU/a4Q4XJBpx
H5df6Q1hnbqcbSxNoZLNf4J96SWuTYrhYNmXleIJ1gKGKYxO6PdH/pXgiDpkfFC26tsGbRc+OnEF
QNCI9JyQvdfS4c762lNsvQsYpsnrw4s457nA4YgxXH+6APLBTWOg0Pni8GIjKzC2YOirn6HFqxuT
YaD69UdfY7k+J1GkVZVCimWR+vgErjPMMu5lc3pplelYoyvRzFKe0T8eZUyRw3g+/QfaOXKJAQwp
1mAxWPzwTJpi5z8SyC102hTh+PV4YhpSCGAvZF9AG5BlZkGa6C56uDTTGNi7X9JVmRAcGkmWKtS4
AGdj7sUIhLQ8EbaVZcmdnh11ZojKa6CIcGVnxUAgHAOv9lAJ6IFmr6agS2l6csabxjjNP4haCBY0
RFAcU8akG7fawyb6iqfa5CGQfBRBBJPpCVvKwr7UO1uum+UnEII/Blh3/zeKz0GJwsT+Mvf7y8HX
IqyQdrVTE6WvRT/qX5/qznwdIyfGT1Je1I+gcyYiAmimAvfmzNqNamLZmnY1yBS7/0wdLwQoGUrU
Vz9FZjELle1ird33C2HGA0qdXsUnNTSUMnrpjRQ4bbtHAL8aA+5PcfvKxNXhLSc0HeA1DCPBgbBH
jtFAtMQTj0ejjzyNLWc2N1aImqPDnyM4gD99oTyK4T96SnhEmefJUcCaeiusgTWENO1J3dCpIsDJ
wBFqiqeiVX170QfBI8UmBY2+Ez5sRGnBn2h3itquj5AjsI1dTaWxVdGRODmV5/V+58SZiBSBJ+xi
jsSeGKa9XdDY2qVA6PpnW2UrpyoQQJm7XEs4ElT13ECdwdo9WdvS+ZXlyJmqVG4vCx2v3LKd4sXh
CKt4edmlu+jSNEDWUrPIWVQlwqVGEBkNOroxO2K+vw9sA93bBXGaO4YxIUx374JVj8Ztt3dHWW4J
PHUo4uXdymFN6dDkrXH22vMpiGm4G5hFuQ3GV6s8zgGVrYeRwGT8CsSihD0yzV2X8BW8twI1WYRy
FdoWu+sCDyiYxLdYTg7FwEHjwB0cdopwTT33HUNP25ACqW2R0aVX4LDUcmP295HaYJSKOhT+KTkf
kPQ+hYwKAeUPkwSCaMKTfhPG0htUtNB5AhfR+StvraNJLyuXdts2W7+NnG1VYRNICGWCZeNIlz1B
hClC/Of0DFvgKaqGrvvjRYDdD2deeDUbMZojoeWK9uSCVjWeZamu1SzlZdEBqqCGn0phmHYwiW95
Tz9XTPx54P+0igpUILAsT4JUQzWqpcFXKZB27LGlRVN5VsJe8griMMk1buio42v2dhR6xW4m4lQC
2WCQbCnuBoQkUgnLLX8Tu8UpOheoXtQfivaBfG+f1V1NJqSq4AWXNfcSnfgdg7GGpBzLQt4lDl0J
vhOhcmOr5aaO7LVsmjG+kPjHecEVIXRH4TpAbnpO6LTgQ6uV7B2EK7rGhB6tG3BYTVKwC5YtvUjf
GMiN6v/8PGjwrs/KMQ7O4Ui2BhWVgcJx5d6+HxBt53DXgxQz4DgxGf4ZJaxREPorm8yzU/W7slT+
57ZsCIPUN682FEGGD1ddwaFsq/uquPStsM/crtMEgQhD1/II1+OFEG0J7xdvlNO5Ypjps2nQUNgk
p1k8oLTOA1Ty5ZtKR3re3F/q8r3cmFLXFgDhyxr6bbtyCQAz8Iq35XMLu8dS6QyMPuPg7UiHrr4u
KEHqHbw+tJAz3D/CxYyAW7gILBCARiMPOYWj2HovMZcIGJ5oGclGjRUgR6VX0gIpDEbx253h3RIx
Ou5QJisUXCzbwHnnDYZUWEravwZGtkrtALe4+Frsz8xv2P4gI0sbYa7ZkgFiHYrySoilwhOHWwY1
RdF+zJkN9Ds43Kske6/94z0toC+U4x3/KA423o22oF+VXuS2FTBIjuBrpp14D5Y4zO7P+jfvnTMx
npwP2QUXjO+d/FUdKVhKERrbTRKOaK9HcytKmlxw3n0CgRoNhRsqND+ArBaRCq34wfNoYQZ0P2DR
+WmGhreeXqdh9EfuUUW+1cJO4sk4Bjj6345lB+YUOu0LI3mTss/GU7ajMGIurxIvLg6WNMw5XD6t
2SDMr+aBxYYF80zwftIZJKkpQNrbRyy7Ed9KrYOsRh54e7kSHJliHf0AeLxEygXXs7kHaCyXJHaN
lpiud279N1JH9zA8Tr2hne1LN+fqDYOQUPgX0pCVNMNIrZHAE9P+aHO7Gp7fw8gumr/wvwbaC8TR
SIbghK4WnZjBBpOUcR9iAs0Eygm5VF0pjxJ17FY6c6JK
`protect end_protected
