`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
m0o/a4mz9YNH/WRiKFnXnbS5LxDC+FXjpIznp6EsACcOjV4mEM6iUvZndrH9AipL6DDCXDDoQCZI
8Vlhuh7xjrVZGyKet8BxeBP4rbtgS+h3luG9BNs7WPxSCmNHEZRPFAkEuyKz7tr+Qhh0H7l2JmW5
mDMnRD+7JVZP535Ga0DE/78a3qEHyyvHDoNZHGvPl5JyyzZucpxRkcaYwfbOyFTBDUIxebnURgVA
ywU/zG3xPQJ41EYCHOkVZyba3KzI+dueTDqcvKHBWHdi5b5pkQCgThgVdg2sJvDwEUYmpy3zryh+
Qu7peKZ3qle/xittxhEHbfUwp/4iOYt4XkgUBw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="gNRsaamW10nxgnbPELbkhyV05DmW/cruYEfSd81gn10="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3520)
`protect data_block
JdEHZEx1W977umWH7OsTH7npHyIvoQhjWuWP+xXcntBkBbAAcMGnuS+5zrvcrZIuOiaFAYBSDnlf
6tR2owF46MubOrcESPvs4uiAGqzROanJUQ/mp7hnP7oytm3Tunw5iT7JYjEv+i6KeLodRV8MJWZJ
0sQVCwRnrjMX26QIab7Jo079qAwFfoE077McWWBFf5fXZeFPtdF8qxj5q0IDRXjKYMNZ/vVgGsZk
BmhfPtKNiuA5R+SphWZAmGP3pEBeITrOxH4AU+2sNnHnrqJm85g3HN/qfOl4ZeEmdL+mb90kVyg9
AWaG0Lm2kCEleTV7E8BHAOIpeYDJAMunrlCEdZ5SN79jTQsQXjro+/2Hi117NgKe6FBVlA+sjYtg
rd45VMEKbeF7NP2KAdXZwvgOrepHHMv6K2EZEudWHaa7d3sdtMYFvadJbU845kt5FUS9aECxCoNY
Hlgq6GWZsgBThHXrKoT5U7lEcn/PkxdGZVE3RB+dt/p5T7INOB/CEiWvnAIcX/3iGKTIdbzOASKf
XWjlmVv8NTRJoFPTu9bNzDGe9f9b/0yAcxZgrW+UvnANtakeMrufDpN9EAYKUTWdk/YgfhDO0s51
Tf3g4iEGUmN8p4MwONHq38CVBbEU86jjxWDW1d5ixW8t2VUUq4er2AdCvwqoYD6LPU4WWHF7kIkn
ROC/YfF4Pl8F9dGI7QfHZagljZhdxFWR8O9YbcwwBF0VRJM5i6ZOIpvGCymK65VTW/Kwkqza2pLo
isl+4Z80xVHDOUGJgl2q57oxTBLZaFRwzJDCUi7qYF4ckzXGncKQbAwagN0IGyHVwfza6oKvn2LZ
2gEz4jXGyuYWX6nJK+nSP41QS2p8O83QPRPvjGyfhI0EQCCyPuB31/Un+xVlx5SRKfsoj4/LChP6
fqMu2kpvbcFRO8KdFC3koIaqqvBJwDzwr+/R6ChH2iJR/OH06B7CcBQFMD7E6gSOrmGuRiFQNrWD
wo65AFQthpf+3sJiP6MDDjKxH0+nkhrcN8LCKDeAIQlsOIeQqoiYmN8POek8LlPThqeSS0u3yzos
hRtKI9v6Nx5FiiSSmgl2L/twnLTiuP+6+SdX/RBkXDkhVkCEFCdd12JS3hq+2xyPzIJCp/QpL1st
EyWASN+qL+G0LohVpKcQM14DeqIHfXnxQj1exPx86tonS/i5gI8OMAsL4qaIjWoVWjfiLHQV0nqH
GYx1UDNcFSmJtKnXjLezmXV8fdzGz6SYyCHOeQ+VXYiZ+fY0llP5vGq46EjSl9qhxXR1FIxhl8tg
hyYSgj7sMYv3lO4yPXqyT05EsEGr6NOIRKdkWYflAeAIMDpUOAft3WqE0mkeWSC9+QDzgYCPAIs6
ETScnIdC+zcehR3jO0QR76hkA4S18NeADn37o30BjXMLBD/EucWioDUBTCf4Ja31hTR2wd7mxgIE
xjZQgissu+xPf+nQhacy+7qpy0mvV9yMpzr1xIMn+iRKzi5kyWx6F6aDB9S1HIaNAx4FcwGCzZL0
Db1oU93TsmTLPvNf6JkmlqxKH/VuBTsYsc1bi9n/+7H7sUoi/WrzoFNtT0eZidLX/DB0Ck7JcxcC
piGrgpHQteBqqO1njXImM3bBWc9wmMbwtsCaMBS7bgstzmBWRfbtsIMMgAz1U/W8wpBnprR4RwPR
xdMboTVZhABjjuMple5nC48Rt/72jHG8YHdgdHIqa/FSJ78UJQSlISMcN/Vk31twoism7fQKylBv
5MiLB51dGI+mwgClwz6vrlIk+otF4knHaoOG0fcQVDy/r5CmUmujSn/yrQcisXRRemWWJ7UF+jzn
4N877Vw7PXiaPSE8OdN8jYLYi+Amq7GZrdJZw87we/g88a2fmcyiHdUlsrHiNRkqCR1i6BMDVE+t
o5GECJ/Se8dOqgynTlBtdt4AStgxzSKfGltwYxQgEaHjnmlipNyJtaRNEhBhlL7xQC9oz38N/Qlu
5YWFxUKaS2EZ9fMBp82nmV2fCKFMHSBpTAe+JjC1yhlBMWzwAeWVhESrTAIa6Uk3M01wC68FR8rj
eXbyMWMMZMNkti5i2HUOOxUEbbZcIb8IiLSegh7Su/JETmen+TIlf8iGC/2t75PEe4ulJ1/RMZSz
Px7RAEW9vpxvx6Aa1B3uj1MNdA4GrHv5Xnk8cEgRtZVqJH8sAJK8qZWGmlEMtZcl4LJLVaRDMNro
RV2qWmNNdTuHcz8n03zWvm5tyWPgNL+k71l7givcG5Ob7IzP8Dm5jNTi7YqdeaAEn7z9ECvJBok8
YRGkATD/Muxb2Q2CTLGz6rd0XVETVblLPavBW2AN3UNy/mt/3lNFJn/RmbN7dC7zUNqRGkC25wo+
ai7L1ijKFhZFuN4htPsRW+z38OvDJDOVcjZEZX3MiDHez05lG+Z+B+ZpmHLyVY/QHZfxVaOkNb+4
xynl9k12OBrHqzAqO4dpBhUI5/FooxdcnmsxTZuZRVdsEhehmidjxFFjAKDCmlDL5CORhEjGY68P
X4q7fUaVsmqYL+nryp95oxIqonLXCrfqHnKvcC8afjy0h23Znotx7qjAMDkRCE2Et85Dh9Mgr5lB
vuVw/WlMIS4ebvvC0UlkC2Qc3do6sLxx7DZVJGsXD9JpR0nASmpeZcspY0RWiLXackT0xBmK6ZpE
P2bsoLPMGNprxWvYhK6S7Dbm2lDnWrCtgwGrqsp99flCB+0sTIOmRCR6upaHagiIU+tV0zaNbQtN
8+SAv4T0bcJ19AQLonZqewfVfKuGkDhH2Q1rCFpmMXuKm7XepNbJD+4WxCOyE9vdBEt2OpyEQdDC
fU7EDqiJ4cpAq8R1RberPOG5OIRTZ2mapDTIUzI7tjX9dkTOmQSRv9tYggk7E3dpOC0/B/amJfo1
pOd39gFu8dxAoN/1wF6pIRJF6ygz4grTkDR7zMGQsCthHPPveCVrOGFI5mSS2wlar7+IhtD89QaY
w7FBRAQnsNeWquI5utXNMjK+5z3CYJycTEsNuejsDR/U8y27kiPbkjFrlwSZkjVrEnjIlp3wvUTz
MVXTw67SAp3vp2jVa9PAqh/9YDn5oaVlvGA7FJjb3yFmV9UyTT9zEmbvRPQaBVEe2cAHFkDD9Ikd
YPwg839Glg/aHb4txoiHaXH+WUXdeCmvHBG4VoVKO78F05T/ELISCjHIldy78e1ch97/DVfO+ZUP
gu/zWhZYfwtyuGOomUnI6bPz6uFJTkfHfLrk+FueWJQe++twtiMqOh97HoEHCTWgx9iW7lI2nk+W
Bs5wMoADmQ5XcUfWtoiQ1IhrWdtIwwWdYy2SsBrX127YXfG/yBEU4Vsq8UTmq9GrbLLmPLKNdWMs
NOoRe2iAggE0cRLVI6NII7C8Cs/k29HoXCZJfhVXMq3PB8GfFIRP6rwbCJqRSsk2QFspE8XdJ6S9
TQx85W5IE73uWvazkIEwMFoadD1+7e1mrF2+CovGEEvM4kpgTxKSfkF9FTjH1wR9iYqDLWfaUoPS
7WUBvfX3aupdrk9am56DewcaNYzrjUIo8Rxu1jX/+UCN2IJU+eO0jJt253I6qJIQ6j9mdYftiCJu
oV6tmnyDniaJfJZge1smPjyio6590x5vK143FnL2Alsu07Nr4xIeBrD41XXAnG//GxhrFexan3BM
MuNt4U8pzepQfm3/mLar+iSHPkP0/ffLKiffjHmt6WDbx8mkcfgAhVzebPgL3EbtXuxoZ06cCa7w
JQctpZTyuH0rG+IUbBpYM4JidAnx/v/XA4KpZu1+jV51dY24TyRby3t/lxCuFpNeeyCt7S8acs+b
lbE/Q1GWLkO7YbzgtzqPzqUyKi0eaH5xSYOoZiD/Bxwvb/n3gy1mTRY+a2zRvP5vxFDvRAX5UAAx
6L2vQLAIfWmVHsT+UK6qhN7xaYp90t2r7wQLXaceLr9NUdUH/iVYlicALY0ldtAlVuFlkSqo4Z8/
L+YgxbL++pVMBlKCWsfnYsrE0LBp0dhs635agJXjhFHpER/rpI4kFR7iMqfrK1XiS6rUiatPkq91
DID2AeiCPYvAaz6KPXH05Ml7u8vEgSHT2btWx5TMge1C5W6vOME3dcOAbMEDU+60FRVfend5011G
kyYH9rCNuFPRK/1Tuc4cFyO/T9LKHDli2L7UCMs+aGsbk4Nk6hbTdRqVXh/v871/F+13CPkxlRKF
EMLmAENDt4QpI89SOhY1/tQBm1OwkHmjKBfCXkqxCiEqh3yeqZ4YczmhMi9/Y7yxaJhmt+Qn1yDN
sDZnnfaQvwmwnniceZVPKuJAcHr5hGUT5TXF43PIOehPuuIoUWccqnghKT1PBR3SKEi/prhQdBtM
c/HmhUJK7UejvQpk4Tw5XdveB1YiW9gFXGiZN2ajLJz9SSY6oFWiy1m96v6a8qD3h+frKxfQEHD6
R/S4icVoGd9EzRap+cpyuxdbhBS4S+U0OPJd4vgaxkfgYLmRYgm/qz+sb3X8k++1F9O7xHHamxjO
qESzCTLTVklxJZhgp3oWPIdpG9jDo0zT6s7aPgQOTaH6uqLdD/JF2XoGz/LXxOcUD9ynL7DnN0gU
E83UK6tkUDUErb5xmhMp14dYKpFDJTC7KZTQ6rySf3Td2EGUs3jwrWH7gyiDq6DiNiXvCva3UFel
TIQJKfOcQPTp9j0m4GkQZW4IauQE+rzDzsHZple9Hpq0sl4gFeAP9it36g==
`protect end_protected
