`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
AAEKD5WNVcIRHRmfBF1Wt2X0aPEgP4Jr1WI6r9mEmcfW04AbokqnEB5ciHyFNH4+Xxv01TuMUfEo
c/Y8I/ONPsG8ilAYPEHqxXRurJMqxM40MSkJuLIvc6p5UfhbcT1X1D/5W4Li22QLnpSllGrsx857
9bXWQp+GNGOti0ioTnZqJfrLKelqgGT8TxcANg4gdFYjTGFHToey3TbC0V4N1Cvr2hlS2zjCaI8E
Vf2izsuSI6B949OnPF1zbFJooQx96JCFAu3qfaFmuXX/xckOdAoMPkAGspkEfgk3zfwks1k2t8xx
cwfvO3R646XGc+sRLPlgRlrQDBK12DYmVP6gJw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="N6dPAVnVD0GbjD3Izto9iJx/eROaUhA0M0mtMZaXxdc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8992)
`protect data_block
7Vz7FItV0+aAgN5/qRUqCu/Fx5mqliDZJ/cUQCOtzG3Yp9Q6c+8yryfgOWtd50i3FYVY/ZjP6LaS
+HohrCu1LSGmMgA2rsDHAi+k3mDGX89cNAqbHpsh7bXm0dmEhX0D8LN1+w1+Ex9BugPl7VkOOJ/O
E/UIzMmbuXXUtI4jQpRrR+1IP8Hul1o+4zkpy7yja+e832YyS1MwiExkIwDv6Ye1ZJ9p9kmwSaRD
NqEOcYeQN3ISNFqHmekJwHTTISHFdrOggf6XAVCxeIiiJm70S+/pphddtt6LWL55eoWT3TouAOkL
WaCJKFzyWL9PQ2tSBOjFAcsehHkl3bk0xZpScu+eBIr67MJpICDBsQnFNZjGfqU6DwAV5qN2yxkT
RxopRFdV3SjoGLOn/Y1nHYSlo95iCvrutHZZz5snNdlrRGLk9ZNgkphTIiFiHNhSVEFyiFIM6Y+s
YJnEYw7wkD3+W5jMk7CX79kz7lE0ReVKWB868dq2yu4SLulQfiK0pSTNspuRffTY1hb4gnein99F
kJGb/9B37j3iSGmd72TIVKDaWscrGFJZY84PixVJNNiXyvPcJemffMef0bNKo9y+haZPUAKRc4zI
8OknmHD7mwfFnexOeGfBTr4IrzGf8T24B0wA7Q+z8Ps9mluSMSfyxwO4TkP+NmRtzI+Tx//uKcFM
bPWvH1bauOuP+McWQffgbR8ORrlholODqdw1mIOtUDqOUuIA0x+sZsAoPTIA/xqPJ9GMvV/LgQJK
1pYQtUzJ6u3ATJ7gIYEa3Ga6/Fr7sAJ40xl+WP83Qu1Q1IEx50epSZFAyFkEIUKFOWrY87NWt2t7
NYv+hP80/dK7lPxwUPyjnfeWAplayCWuewhuORrdIgDZ40hcTfXR2/GRU+7+OasiUcNIbqsAw4bd
81YPtzD7KTvbf1Iv+6KqwBiKI4uyVbRevTnQMlw44j6c7JOmYbR4WM2BQK9yxb9zfLuf+B5o0pDS
92gK9wXsBu+momRYMUO6kXVDyhAHIaQN78k9Y1thAElEoDNSj3RlY58E2crMTr1UkhHJhi9tmfNZ
NJasxlQ7TsHrappFcAjr7U0L2Pj+sP/E+Oaj7QQlutUO0EHGB9G7hRfIKC8ujEuLgg2t5m5Yepto
FFKgG1Oy3d3tBC8hWdaWviYQHlaVyVoJIpdWBnXiTpDp1Hd6NSYAi3ySFVEkrjPVwqKVxB60t8x5
2VaM2Vp11SNd3zxRMFCkq/TKNDC4lnWy5/J2jlMqWKQIpBrBDOwIyOJHlLCzyz26TylrGjie6+OY
gxC0kw/wrXyU+telaq9grvZMrsXopPR0BaiBX3Lp66EOd7CwBbNs2PCTDtz7jJNWEkgYim150wf4
pewrmvXpXlgGc/o4VXEciyPq5pGjWt978dKxM627aV9debA+e5n63Ya7B+PXi69gDdvnSFQ9a6nz
iMowFRSms4FSURyH6eqTLvvTv0d7160/vxXrh938CyPDP8gLAGAaieZiccLbDdlF7zf7dt+TLsLy
hnySiOFETqh5x41wYTPHIFFItAWCoLB1LictxXtr/O99sKCeIk6JkyIw5v4b5SZVgI08flsjlVrQ
/JpX9sP+/fuChh+X/UwfvV+W04sAZEhwp2nDVOEFitWAUKZW4klYXs8TAQtuZLTGw1SMaIK8TlWD
R73WGNJ25Jp3uepZ4rtMvua7nmXu3TFgy1JQRzsjjjPOdCFC7mrpvDHqdtjySrRImyVkrSraXpYw
Ij4O92B30a/JjhRnRe5lNv1x5vd+LPPQ4Dcmh8fCvhdQfyXxoWiqTw/vzi1NQqsiXUiAnjLa+Z3o
mWSNUOui6jopzRn74rjWmTEWbNXeIrAQy7//XfAp8CyjNVNMJBHVbfCpLVbWLw65Uo/8SqHt8oQ/
ugPnaZqNyC07iELMjuot4ifnWOtXCeacd82NfrtHpjNXAK77FOfRYB/SnAYFPe44EsYU15u3QyLH
5yH/jwjrA02YruKEP77qwMcja3CCQYwheO551v0l/go5y98rrRjt8einUbVhhRdBT2/CA3I2tw90
zlihswTDPIHboRJs9blIeITEoNVIYMeegdD25Q6KUgJtVu66d4lt1+L9ubS+cnlHcdBFPvQSHlFN
cFzroNKp0oo71UyuIbexe0G3Alqw8XEC7L6c+ER3SRnNG1MsLohF3C2s/81okJggLzoBfhWaaDQK
GMZTqTtKGzN3SBP5veJJvwzvkRAE3QcU5/XjFck/fJzipb6huyVa8c6Lg7nSmmeuChyzA1OLwbCK
hpv3fd9vJ+bjTFAU74KLEI4iONVLsF4JCR/MIhLd2CCqSGmc8FnOpnVE4M6mYp59vsXHTcRntpcZ
+ZQpr64uWy/rDZa+8IuAbgV8MlS97u6Cx+cegQWeDHlkZpV2LSfTJPGqPUhe4HxJA6U0xahkrAQo
uQwc3uvjiL6sxwXxhgAsa1w8KvjbwgtC4x6N0YuhzhASrNVnnFXHyoBjqoRNfQ/N9bV48F/3LEdp
7yPMmtV1/DsLs/ppWTVNQNOfZ0TfoJjPaNAjg14NGERtF4WFSzOY8Cea8l2ryXc3UJCMWB9RZNc/
c1hBVmz3TKjRmc+7YE6gxN08q5KentnhF9x7mXiQ+oVm4ec0CDZ7n+5xuL62cRF/QrCbMFB77qe0
qJHQp/1cYGyy2FdyyZybf+iDS3POD7QyzjKERNo19hXD3F7fbutQ5fo/AYdA6LxAXubfRmKP66si
YksC15Z0nHWGRJP79asaVUc3ySvsVkKFDV16Gq46lRp1YagJEzIz6OpJlQXvrBOvLz1eEG1lsRQk
kj4wZFWiVZ0pmR+0huNOkvtLUO+ze4hpaloaskBP3DBr0HvUQGHEO6QRmzb6Wxf/kTx8+JraIk5o
h5Tpg338aNQjYmDlL8XbBuCzOYFZVo1hRBco5lB3VJM2+rPebvY/5d5EA1l+vAK7UtBf90enRfES
65FqwVtBgcwZ5TH1B5WP9CvQhjmKaPdfDIl4tCFhkjtPkBhzrB83m+xk4o5JJmlWxJNO1XYBpCX6
/PcfgoaxDBwten3BP65dN4fVvFMH1h8UI2es7gR1TerZlVvxMh/nTHzqKoSF3AgUGotmDTOBZ4+e
Y854vTrDS/QBZuRTKyTUzH85HT21YK1mgRs+vuFx3s/ezx55AsjWVNzVOITLcipAzgMnqmOGbaE5
FFCPIKbSAwAxGYMbXx7HE0QgrwUdOvYjE5b5T3XdHFjJB3MjPgr8RzaZVnC3bQySirxHMHOm79q3
9bp4+1nEdzyq+ucFRfERoqUx2nSfDepoC3OlqDyvICuNP6AOBJYWQ3klX1VCw2oIqs86uQizJW56
gOIR8LIjBfHq0IGV9w3dvyImN4n2/6RNeAGZVuYT+y7wdfyfVGRkl1Lph4xzFyeji1v6eCOlo8s/
QsqkJ+IfzyyzEuzTxQequBN4F2L845HYGBJZuu/lUbUlOHIUrnui/czjpfyxakq5oaWy3ey/MV7r
nnmxlcctWRtYI2pA7qG2NTQgjvpabZGVGyntGsaMGIiUMpC5O1wTs3nvKPGAckVuHTAvAIx6Jc4y
a4XtBh5k5V0G95tp6ZIY/5XBpoF9f56iS2MVmWlEXZsgZ2OTsAYq/UyPwMeYN1OVEZ/MTz97GPs9
ov1NXiZ6ozyfuH9Ze1lW4x+unyRQbw6lphmIB+tIrmXwKMNQ4SoKKO25DQLXNkKeVRrx93iq/QZ6
Od8zoHWXMfCsjw5AQx0LBnA6LtcZNgCWHnw/z1heHZr2C+NudGr5B+RcB8qtjKDiHxlwilMj4ztN
bflELJTq104ENlLryURnFCjrq9aQpTq3L23YdYn/Mu1qLi5J8ffggEv06BWkFZ3QyGwHorhD9oL5
T3kpQ6cXvyfZf3fDbtvdVyAJanV1yIrZi/JW7Bmn8n/x0izTEUctboW3p9fRbkfH2XNUgfr2P2zk
GwNX2kvhqUjBiQNJxAfdHBiA3c09ekvQUq8i5M/amHojXU0Er1Wnsh8YEiaslplpllN8XvYUYxUQ
MI5ucskc81jjGQIPceKFkWjdUi3HrR92a97vD/lo/2fqn6T2cX+4ATpDOd+fchJ8heJtQ1RofK+B
8KqKIb8tTafOAybsWVR31DpeParZjS9NnmmZk2DmjL8MIehbIq7A7N3azI/3wq/eAQhYe2MFF66H
TpqGMVX0Xf0zSP062rvV+zDW7FFIfhEwLPhY+FCMVbydwFzb9ODLVi+pTi/z+syeOnpD+hYrhCvw
D/yRb78T6vu82eQcEHMPiq4F3vfOBR+7XAIxn/pKEXTlOZwriVXjbNnyCw2CCJqYCgnfl3z8EbtO
ywBkncg73hveKq8s9LYR9cbqtl8eMbE3BitJ4eK5LQhlxQcwl7QUw4hD5lRr1nh+dBcsw8cWUIxG
e+6uc21C6UaDhGoF0dfZDWfGJWcXSgSfYKQcuDX86yJMsR81yujoKRnNGzOtk9WzUxKiBNTOfGX3
zm9c+VjPDsr184u27wXHNDpSwg7jZ+WcwX/hxFfFYtj+xYtViPoJLEqfTYuLc0grR3/E4ZTfcMOu
/RISHvLXl6fimj7kwGfwRB/ZWNjbKbZ/N9EKVv4sn53P3oD0UmmlCibaXdzMtzKgusc1kNmF6Cm8
IEp5I+YOHk73HyxQb60HjExBLZrneuBt6hEAlle63AJSDdYdd+ObJOCNj5VK9PV+6M2E8Dk/H10U
B06YHrAtn9t8QZ5Dg6GGDUetq7UxK2O4+eYsrNZqsXPyhBgO0Wz48k6L+3HLuUzRRz/g6s5eaplR
f+p75lBOd0+AfxI4U12nDZZikrtrahHn1UWyDOaCQ2h7sE8ekpQa1JDadJp9gw/jlAYuU7nxOQHn
5BSHa3EWeDAL1aQ5lBn/foS5V1BfvYzmcG/nRhh2QFofn4jaTN9IVjenKjR2OIYR9ZC3x19obotZ
fnftRG91B/g/Jwo6RCpczK3oiCK1+UqfRpbRGBVCjJqccq5L/fySMfEujlG4f0QF6HFqwuYRUIpp
QnCd755QX+wgUtgjhWoQu98pduF88pQLG/QHIT4JJvTlb9wpsR8/ApwNjGbgaRK4XGJ6BuDAzsfC
X0UbSrdd2TLuCzzA+jgoxCyzY7XPddn+7aNoLI6gYZEUhRgs3NdFJjjGKKUV8pMhm8QDSr2K/Z48
gunQ3bftNXR7rtmDJ/1upmeCWx/P6+Z6g3XZwX1itc+Jr6xUQA10n9ITSB2zFVyY8yDeWHD97UyD
7QHT28nEyk+9UGQhTzYonFqyEZoNNbAo9cr8Edi/AzoB6Np85y2sgm+K9Qkx3iumDS4kQsLUwW/R
Z4wn8D51wOz3RyvmDIpkqa+s/PR2u0e/faHeOAQ6z6qLyTDGP1YTrp77XcmCOchn9ZeZrqtAuDRo
+x7rdDJ8eTiZ6nWPN+gDFWiS1jE1MoKAsVx405yb9uB4Tp1eVcfk1mXf5u528o1H7+lMw74PH7Bt
ZPJkLsRctZBORdyDzYjUxJAsCGAmAG+bNQjvffXsdP39/mn5+k3Ype1CO6mDlSU105DPEM1FqkAv
QVv7P17teYuSH9HndJLOfjjHCZEiVkOiKiY5DEP3j2jdBKWm5tATfL9xdlq4YU+qsMiq4oJmOKbt
oc/JhOeWwC+rRUDq4+rlWd2ZZVJc70vkHPXtjo2FthA+bdbAUVXYoMykKbCsEc2aMzW08TWFGKCD
s3gGT8G5bFUeG/OCezhQ3AJSgj3LWEYmjPlGGw26pO2ZzUfRgVyPyC4NBES6rnd541mcjSH0ihQz
xWZsmqKaXdA3f7im/iEXDt4ufaEtS+zfVURKEoP6DJQaGqxpADRV2e4v2EKSa+MZDUEe9OdqOuOM
Fz6HMBLMkdNtMQXhCw+ehOXbrCM9RmxJgwiIA3NtckMDCgsi/yhIy+cRG3026F8y+rQxgKg47DlE
ya15HfMZ2Dc1amp60nhVaZdd7evQ/G62zIRJt57D5qDJpdRTUcfIDREm9APqtsnMcXG0TbC6ZjOF
u7FW0Lk0Vwlvz77+6QUPwuOWCHZjV/szi5x0a2Hq9bdHKWhjzNm0WyyPG8eYVll8mqt/S8PNB3ss
8ntA07lGDYOKu6fQ9a3LMd8DXiM3n8T2hvdT/ldHao32qhz1Ns2X3v/TbmXBl7uDzC86XEiAnVlu
pwD/N1TqwJOQ8ArirkDacuoCphcQoTQABGWlCLmhbhiOzm6nwu3q99VKdUvzK8DP3nV6FOIrrOic
m+2FEHqBhyyRZkutfCGvA2tn1W4xeP/Jk7xqkDc/Nw7ZHCsqeAHWENjTz1F6CpXGtfH2Y6X6SXLf
fNK2PNfkoD/2jN/b2WHrWg+re6nyrl2/qcFq8a6YmJm4fyliRWxSiB83HtXqsm9HiAlSseENtEdS
ZeM8V77g4xQtfVrKVTx+syfuLYp+3lQKS0+vGjV2dBzoFgjtKvaQpX+8wDlNMaWdre3eudHi2uJq
grIha8IOSu6/mekhWL+CuNREQiAEUKjBQOhWcms3DP1UaDgDK3LPw35lXjGz9P/vPMFzpNrrSj1R
41qelI/+Fj/RP23CRmqAStT81Ol5Pxj/tAE9wBtPvZzfKLzPawzMhgZQUv87HOlJGL13cAMUzUKV
shA29esQdUqxoXE7HWSh4CMYHlLbvXLiVhjbfrTYPd344q63K+SUZQVN6G7q0YYHc+pvQaAw+/PZ
DJjk/h28ZVv0dozDvBkSMsbKK8oegzxVlV2ADwYxmN/z6BHWwC5HDjyXNLrPgjGK0US8arFBBfJC
J66O4L73ipkS75quMO9jy3E+mXiB2nYbpD+qLSwRYGAO5Ea+3SZSHlK4LCGwiy5k6JerMWwq0MtK
1D4cshDL4D/U2q6oT7OTeJJcCnWHFmjUxruwZUxfzetsUtN2iro2B5IZLDXXA1KhQzTbIglb5SiD
wfCkQW2JcCkCX8FhVWzC3tSQJF11VcxN/Fowc9A3Wm81SNba+vNrJ7J6r1lqlyhkfNirkAyQIQlT
hpp/OBu1CmvvsWGja4Ry7uW5cqp4RN//Hd965Edsc48QqbGQkS+JtboeQX1qZ3AA1DpIDAMVYZtt
Q+dTiXo4AHWPoGsUJzWaKuE5EdlrKPrqD8w3ClFovpWkO+UAoFhN2J+RNL0mQYjfp/v8T99H5cJ4
ySl1qmnFTHjennesolxL84vIhrdZh2YozDtgt4pir+82NokagUMEnk4qYDgR/yxPhiP7tC6yL0f5
1w96Z5Ruk/1NA6IZ+Iz0lNyTGvahDvn0Iepgkg94w8H/OcZbxq+py8EzvkpxuK+4LvVSX6QGwZMK
WLlt2FdsjRCP+VYQKstMI+rOOAp2khc6HH3T6eDosnzYnGC4tikGQb+Tq8MfKyg++OsAiNE+ualB
3NIcxQoXQgEZ1vcca5h0hac4I5X+9UgRNGDC0SYx/oK9sxoAN8L4+HsYRcJWd+VzAKjpq5/pGbwy
p+RHq0GJtKu+zOwqcjQjXp/x//jfi1Kubu9RjMKtzBpYjzwlSEczJ24CTgf2l6H2CfUoEhP5Z/SL
clnVseZCE6Cqb2lNVPWU2bKdX3zkcUO1oCHYxFBszne1oCeRqwCKhDnuhHQF96JyWV3FPhu159jd
cc4slQUyO223e4nDgO5Y4/UYgZXRzaOP/Mgev6mPZJZ1tmd8Or5sZw36ShnagGC1KPVX0QqJfRue
SQcxlcKy7aJZ5NE06RFz0gW62ZeZ6CA+tKFtGxTa3Saj6FG26wR5+/zjqWdFRtTFNZaztkhtDCqq
Kchn6FEF8c5PDnKGGzcnmR99xNbQtS/dGH17EfZeiI6cA5nedht33+bSJ1TLvvAaF4G2veAbo1dW
1jgE+Av3dD3g7qlkaQZm4TWHj1jjUJZ5z17JEehxqj+esZ63QH8gbckddcY35c/ZEDtLRQPL9Cn7
gzkVgH9e/Ohv919gzSL6NAn1d6z4yyQ4kWpi5qO6aE7xQTOWJtJAprTAlsHaDAlU25lW/00WbpEw
fLWss+l/vRiYikz3ECr3nFEFldHhnZthHjWk7i0MpTZetzW40xjG+Gct947+GNrksPB3I6G1fZP3
bXx61eZd3U9kiRFAdIIpVZdmLA+YN4GPjX2rMl+DZDUBFHFLa/KQ7mGVxCodO8SAc8p/BNK4+a+i
2O164bgAKycAkV26SBExZEshM0ZKSPyHO1tRJsudn0LKy7ekQpCWfufKbHbLC+5HUPP+FfG6aJoY
MnDxiL6s6NdJOGdq+b7u9Inq7n4Yiujz+GfgmbsEmqihs069PTasxl7BU1wH9L+e7Yy+AVHW5kTG
KjQoMyzhiD2FUhslIdlQYz50RkbFwE+z14qriAYBHkA727M8hIkZNYcLlXYgXfKD5nk1uMqTvGj5
R2UNtGpdw5VGbS3peRi0TKzT7H/PeB+w4EhK5qfa9qBaKZflQXldLlIWNLD56/Nm+SOHK6MSDsHw
hynPBBP3qA5Y3BCd5XPkZNdv1u9C20+IDrCXSGCxuTkc0/1B8W6EQyWFje5wKrMXqiAj6H13hV8Q
CvzqR3yT6f5hjpv2yatxvNZDCbSVqs0DSkOgY+BlM8NDsyqszYZYRi53LbcE7g4ZncVGO2geHEOn
i0z8ejsgaIHLgTuTVqddUnCjU0YErE9GX6JrLC24oEx+oKX08Gt0DyHHH8JgwmjNzQ8xImqWaXBf
AYPGQUzAX6zSTtCbyjX4nxoTZzHe2aC2jvOxmcfEG8FdfBg9pRiqU9ckWk41EZEjkUR/IRcBSHuc
OhdHtZjq8mgd/wKwrYR4H4kqUH2f5TR4XDw0tGtdkzdXiWUdN8PEjpJR3lpA7K8zM1nX/wWLXo96
aRDbT2+RPz7oLxVWmqNeeCRV0oKjNuI3ZJiBugroQxKQFk14kNKPNBnBViFqby8PGE4J3BJLBGtE
nL4FgrFk2ro9tilHLTvKDnT2yPfj73P6l5RLfa2uCsB3tI04/TqYRMrB6MOLKKeXs6/pCESv4tNI
/h0ksPtE2dzfZGX/0DWfMKI+8lvu6fpFy7KdheEWenX5Qa4AoXFC3XMN2ylBGuwW0dJ06PWm9q6a
vtOuCS5725/n4Qm33dG+V6hgMfiHnTDHC26AvFOS1wQDRGeuubTQnWZFGMZCDDUOFlwz+1zPy7wn
Yhf2dKRHCBc0Aoeql32ytpwt9PlUdZ0oYH8ReEZBjF/VlPRvpyRd9QRS6gJLSBE2a/50xzH79Krn
vIh5WQP/21CjmYplNeKcctE0+2re0olneFtTyAnMhixHYXyECh4jpgI+GCtbebPxwWFX9ut4lUvR
WMcAY86gBb8gH1ZLhfBgeWaUUVhCMUZxRQ5UjeXwqsf2SbtIqiHSTIA2PgzUzGnlYcI9npPuIGA8
V94bLlwHeAa4vItrcKehks1WO/W2nk+ALZk1gtxS62KkR5ApFH/nc1v/FzNtum0lLOCrozhDjOIq
N6sU8P/A1PNjAyNTXZQYN//B5g1qbxDJ1wKUqHEKrb5y1R+A+nfhxIRStSX0mJUy5DbcmLRwdB28
EO0zwlTwTnim0feurr4SFHwL3qsiUipvuydY6OickSk+CqB1sdvyeaTxZrOxI+2mR9BeAAscSy5a
EZL79tbh/mJHdpBUz2oqAI6UYgpPJlmqVCEw+ijwk8U5QrqmtK1GPuJzq8qx+nyBx4L8TVROd5ay
sqA+hDYWIARCm4l1mH97/K3i5XKpLmLZbQQdEtwHxEDsl+JJtDEKUgBP4HRkMjLh0PWkMOt3emdx
Tu8UgD3mWZC9blGTjinNxcvQSSlEMILmy3b2EOGFw0etstS0eHJsGLE8TbxJam7SGsFBB2D1keGt
pNBsRadzBudO11OQ9qLTbm5dFlA+HNkXUWEYZbVmZiAjEJkbOWQ6bxCmxRlCpoujlOlRNxHg/BUD
6kHo9wLcos7ecHsEwFult7PcJGvQpt06gQvQH33oJTR2A+2eATYXFRU+fygCnKe73xBBccjwCwB9
FPKKazkgx2ya+ImEtSzcPGJFoXVe+++2VCg4tzsDC+Lp2smXL1uvqfgk+b/auV9vH8VjhSDFcknJ
JEsoWZHSY6OLjcbpihprEJQQaomu9YFj4/Bc+MZwZixc/secGww5AkmjrSnnOD/dez3QkA7+Fa8V
HNtkVBfMyShunkOUlGMDt96fuhrdedNw2EDiZy6g00AiIrEkGekXeKDNTyu9GMMHSAll6PbbtWJX
Vn3rGmu+3x3zWcT0BkTZQ48bRaMnK+bZGQd6s9hBR8XxE7OvuDeHmN0IG8qm+0Ld30IFc/PJplSM
uPeFAZZH8Xu2+hBMFOnyIAE3dVzQ+bEhh/MXc3jvJ4ACekdc4RLDaAbC287I6get4fOIBRUuqkuq
oOIEWrOgOV7HGrYUnPLBBnguGhZxou4r30GNAjNjIJik6cWY5o7ML5wtst/VUdELfDMd+fMeF7bP
ePmqCH5BN4Cwf9h0cGfblkPLart4dcDgEcCsa6oL9PAj/Bl2h8if31JZTCssy8zFfOa1KkEXzhRO
HEVJopCmk/OQPYNY83ct7beGWdE8T1z+Tjy/wayy9zlge68O0ugtvYGICzY9ulUeyv5POzPBy4DF
xemiMoiBVuyAbEt815gvb0sY7cpd//v+3XrqWoH1K5muj9PGNkuJqrdgVcR3Fbq6s+aqgxt3e1UF
yee12kTkjEpA2vN5ZAM6SaCFOvK9UAAc1GQh8vf5jcNDUlbf///YYJXsCAhVRBDV2F+OPD/vdcvg
L9dxUWU6j015dVxz1k8tMgJWGRtdYnY/KC9nu++JRW3ETc6Ytk77fPj/W+AojHagMuQy2ERfZqXq
bg6J0R4V0SvoA7JoMdd7YvGU68fxCpZO8gJsU4DDGnmgimEA02umlG60DQ4uXDY/+GHg/sSd8Gnx
+dJ/ONsTBk7V6FvP2bH+k5QnP16W8m+2bighhPtinm3mIIm3SQoQsNNl9oIzU/B7YsabTREJrNN4
9ROc5U7L3h+k64WLox/ebY+y7Wu/1HE8yKqOw6kp7MC8rG3KO5AJcvXelC3pbd+Ece1mvzWFLhr3
5EY12Ko3xsBkvOQ/Yda93Ji17iEWO9hdNo+mEdqT/OFAgTsCgR/i3Zzwab46eu4unfIVPDhAx97g
B0X1pY3k8Ddg/mGl2evpUnD0013HWxl07q8u4PcDAoXZQkt62CSxsLtGWS2pdQXbKK3l4Dn0DOYE
FAuzhgSYs2ai+7J2Kudt6YUaf+9DZV9PQmD6eRszkWDj1FtGJL7Ko1Kz50/yCY/PRyZRQA24BtC2
o7gKqbyDRUC6a+nUftgP+KN6BtuhfjDRXga91Vmu7jtNYBxtjGAx4D5XSB8AXl5JmyTVbFV+EqmN
4AvcmHjKky4edeOjzScOg5wavmdESaJC+gEw1sPlrbPpb6MwGQyGfBzAqdjfjLXZScDHSLk+SElj
avSiAhjUncXgBGEOF3KYb/qV5GdeSVBh19bynL2L5lKoJHvj3IYXsPv69XC1Hq1P6xlcnNYhbiY2
waxWu+FziAVACDUWv2E48N5uHCtqz9ebIi1Vudu5GXb55QBwU48vHA+zXk2KFRDokk58molzaZ6b
ZlG+4hV1/lh7CymNiAgtw5cfdILmA5GdwntLhL3C3xzfgDzoCoNGxrLXop9shU2VGLJBUbbN1tcz
qxzrkA/OWb/qeQaLgiSQ/JNZkxQ9hHk+DOsu4QOyNKB2yFZWMUOmcKFrarat0BjxCZfwiPJk6s5v
/FxBsj1FG92ksO4/Bg7LdVcF1XLpw3hdVKE6ASyN7ghh+eh/KXF+VhBP9HYfPgriNSfyB/NYQHc6
jfkai/0ey7RrjkIY4LnNSCf/NYxdi9rRkfzmSOSS/HFBYzdyKESyTFgZL4lLoTtSqmZZaqimzf7X
HCXJKdDlaRFqD5oDPJA5UzXEehFjuLVwNnPU363ZYJD36l7VOLHDez7VJ6CVQRhsMtzY2PeXBT4u
ot8OKet0fpmhcNVyAwnIr3Jgynw/7Ba/CpImlFX7pyFZuGb9dpIJOz35mA==
`protect end_protected
