XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��?yi�O�IK��'l��Y;�E_>���S�Yߴ�*r.0�$R�x���T�s��mDp�;5�[�</V�y"�Ă�`�yS �5�@}���7��O���V5x~����(ΐ(,��e�����X~��˦є�̰�QX��������B瀞2 [)�D�!c�r���}a� \�1	��$�w��n&���;풻������$�����Ϋ��A�\�mbME��E��k��$aPE
f���c���}����43t�t� C�T,m�A�)Εh��9�Y)e�jy!yk�JdN*u�'�I�D�=U�P�j�EN�8�@\���3z��S�o!D����'�)Y��_0|�������3�����!b���Lh(�~�MƂՀ�Dwҝ r��{7t�u�F���/�:��M��'AN�H�.S�������]ZE�A�!���|e��a5�i�=	k�I�
�,��>5�)�5p��RXB��b�\�=�ښ�șV��=��[ƱD<H��|�J�!3�*�:��E�p,c��*�R?r�)KIň�Òʈ�U���I<Cm4����Yx셡.}U�\6p_��h���@�WךX&����Y��D�����qg�a��[� @|�\@�m�X-�pA��ͻ�Y깇X;����{�����Ѫ_�"{�P�6,����}�n h�V�����LQ+����&+�vk-=!?1f��0~d$9q��j%ȿ8��W���!�������	{��a�#�z�3,����[�z;5XlxVHYEB     400     1d0�{h3�!�'tf��}�$���^������8��i�K���� ��рס�W:�1��̿�榔Y��f�_k�N���$�Qq����rm��9�&�JPv�K6e�U@��&�m��N�XZ���#��p�s�o޴�Q2� �x�*ןEz�%�OYc�cJ����Rz��*s�I�U�'ˈr8F>]{3*����<-���ݤB��48ԍHp35Q�AAT�~j�l��6�a���u��T�I�3�ď���X>�tt⁔�F8Z*95���+��W�c�N&�|�oЬf���; 繇	�����\w:30�g�<n��g�HT��:{�q����*����]<{n�X�A�3P�m�T��n>�;:)�%O���{-'������'dJ�˚؃�h�A$�eCa����ć֗\������UԄzg3������3�������gWQ�u$�mbn�m��a�XlxVHYEB     400     130<Em��l�c# ����i���X�ȝs��R�x���:ѾT#�^��݄��y���K���6?;��R�/9H�T�*2�"��h��>�+���	߻�j�ѐ(ׅp_�A1�N3�k�D�F9�n-׶����B�3@wXn�DU��ҥًÃY�&b�۫=����จv�EדN���e�KPP���0�ɘm��6�Q�c�N|Ѓ���Pݜ���f��*��Ё&!���@U=��l]�iT>��8O���L���_#�۟�����~bi�G�&�Dj`��KﹶUf�U����]UXlxVHYEB     121      90�W���־�Z�����W @�Qّ�C�!H`�b �|���`�ɇ��T�ĸ�?y�����?��dI�pD��l^��8�8�g�G���x����Ĝ���E�n��p�~�݋�c����	�
_�w�DZ�p���o�u�OB���