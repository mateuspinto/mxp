`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17056)
`protect data_block
0kk+a2nFZQkkBhPl39GppquPD8SpLCD6xSJTkOCVGX4AhiWlFpO9lShMcEsFh3q0J3kpTiQbSbgS
8x+bUP8d7m619wUL6mMgfpnG6HO7kkEfhFQk25xtroxt8HOASJ3LwSYuSEg5TioSFjPrpfliYRGa
niyU7pHUm+2TUVQW6o23ae0gxiK14Nfd4GohnxtedCf82DjgmKSJYcGQDEnJfGTbJd9Zyv6m9zrR
oj7zQNjQCHbTSPIn4TuobqGplCCHqBUtYmiN+Sm8c5A9ILTGd6MIu0ArS2VbjSZ3PuFLdJnV5P4K
i/jYfzGnt3JCN1yzVbRBIQWD5TYgCcIccKMRvmh6x7oZgittns4bB4nAhsAICvez24DBgrirZLkA
MwQXdbW/+sKfLmTD65QJWHPGjX5dCag1oyDNLOwl6YQmeIWFOU2i8NGjKcprz+TolyxymHO/M5tg
ZCT+4URmnpY3skrkk9r0y6aA9DwW/MlRAZ5aB5Sr8SddCljjQn/yQzjRkNcLvj65O8r2kbmGTnHZ
IUlZJmfCaV2+MS5SmqUWbHyKxSnCG1W+ZxWOX0+nURShmhKQF/bEn31HQFyPCTZ0NsY5b7Tf6ZFt
2dk/dsa32E2p0FvVvEifaS+qcAUOAiBmAjdDMNFctqLcVjNEt8STRxCZnGSAPAB5oN1i3z4YTbMs
crd5NLeEOSyqAKbmPplgNlcomEAGlAcB9Z9ofFTLfwKgwl438FCMx6zFLRRC2nPEZ1Nr4wLKvCFd
jaMwaZRe8kqPCyVLb0RSsqZvvrRT10VBA2i3Pk/fwP2RVmhBsk07GAj1ccp8/kZcmIZcuGQEY/ic
tBgbyS4qz/Yi68Qw5yD6vg9ngfUSD9C7HFZG86A/1FPqmvYTESHMfSVf/5hQhZlXHqfS2ZipL51C
KD6ir61GymlP4GDznrNkwiwglDtDGjxOAo1gI+uAdz42WVJVO2fGDEswKnk0nT0WH5ldr/gKzx3G
qFmkZQw1+2UiTgbUGir2cJzWwaFK9YKCbseUhQG8tdKzuDY3cSbmfeHIigbWbYDC6thp/Ozqa/AW
Kjk9UESOG1egbypTPLTBstbFPZ5QRyIglsaFIQtjnoWW2HDD0iqqwbAKk4NKET2aMPjf0Eq0RXxB
YpfZvZQwdxWfLiU/MPyMCLRhdw8jiQI3ZZoaefrV8UpVNncCRb98yql/yXVtoIlHydpnuEkD4eRf
/2qZzNZvaqcOMAILsIflYLb1nlYkG39oqJ+UEaTitt4d3wZmMbZZEr8pP8Stjvby6JuGqNE5yveB
igsRIKA2dLRP78W1Ni3KKbIROh9v4oOPH3aBIRjz2MSQwxvDdWDh9HET+QXSqshQdRlUUr0WqeJj
1RMBlY8QPlm3bnzLFoNv4GpvjQT1Wss0YElwSsoxuoUikWRBpAZVHy+O/EuxZHwPPFk2sBhE/PUQ
9Ptw5wuNPF+/+iSpwEf4jPzHvPJUw6FnHoJ+0dq51K1f5/9w4Cy+s51u8OEk+vw48lFZExWaIlqD
ZsONZ3HARmScqslcef3jVx1Lb0TwOYtLFjiT+QaORRPilsVNflzI/xS7gPzv12Y7JlBqxDnsG8ec
i29hLEzfxJt0LgJzaK9IbSwU9drNeE9nDLrBt4CtIILc7J+YIAXkfnZYauXz56Wj6iE33kg3UnYd
L+fR9JOtDbECCvREOcP4hiMt8/OYQDvoI3LWPYpAwB+onS1oWehZvDqqHHQuC88FguoNukAcl+/g
WQYgSTD/WcAxJ0DPQlTGA0uxx4eJWUgjgEzqXB2HMwIOMGkzNWSJCCT7GxA5UYGvi4yIfvzEquMP
mc0LMtsI2f6rSKpeCQFY5D6pHMJCp4xAy91ymWIX/0EcP/nPfRQjvvYLUAk+N57wC1Y/Qw1K0E2C
Vv28RlJvdFSWCCNhRMTsPmQl8SEGWBSEFQQ7DpoIt151mGyrYTdRe0dhpDGA2ibeZAYz35esl/OJ
2cTwYXfJPM+27P76Z1+H/fK3lG6sVcfqdfTHbabC9C7mf3IA/UzzihxDfLaRzC65HZ+wYssSv3xP
35ju9NtkXNoy269WqbGyCUYXyAdwyQcCegsW6OAjnv3PKWznCIRvIhIJWMLYUgrwslZc6B4+pU5u
uierKFW0nd8K8IW4U29YClTt8SA09Bs8J4LJsEtFJhCemtzTqwnYV45xxCWznYmnyAoQgKj9TwvZ
q9fefC3wOLFVM/kqSlNV7AEXvyqySHbgfcENCIbXTo3wNztcl1EWb4ycAlGnES0cXjwTD0juG0Hz
FELT5Y1jHR7ibloHZv7xBHn1z0TDJM/TjUswlvmjrDKw3wY5AslWJp5aQLAZMq/VByZHvTRWVBtt
2AROIuVa+mhqKREWcMRhYstq1V5cSEEgrjnycJH9pY4eA/Ttj/IyHgg3TbhCS3c1YEe8m+WzPrVA
fTCySYvEoUJt/jhbhxByq4tQmE83ApnlILym523f5hbDde1plamzSK20vS6arb0F1RmX4TJmevQZ
+Glkyf4hMxEK3NQBtqWwWnFV4rXYYsVjfkz5/LewO1z81lyaaBeDh5fHt8ckJo5OsZnM91BG5ErD
krX/pQ3FVcVboP27GVZa3LB40g/ZXyxD1lQiXHSbQvdeFEdJ+MYtpaBEdb2Oed3JjqkbIMRa1lGi
PCsDn4BSfXryH7ttTEJazXTYxOHOcAIOq3uf5jkaVglz41QPqJ11+obZ6UlM17zk8y72E/bn+Uaj
fx42Opiwv+6UM9sXV2g6JNSggfl03D1pGIGGEvIUdHeD0xsEiBJW+UOIJ08JeLFFf2qyzkVcYM04
cqpIuaCpz/ksTPkYbe+wCeIWMS12I69eNQt3ydFqxrdH5Ed9tVD1NsgriIb+4f560eU7uBpfM1yN
SfC7MIRqDuWL4l6MczMvMxrOOo529aI9JztPD4UrM9t3T+GYUiz2S1vlH9ajVRFYrvLJjEyS6oI2
ilge2d80lVZVHGt3RGf2JatrfuKrrK8vPm1Ju78d6+/397b/jFPsMiln4kaHVgX+Z+dd8fsHOJ7E
GmKbqRPebXXA27PWkQEvNoWD45Z3ckcTIvNORKq803/8hQgOmSJqncW0YS+VV7IYTs7S9dotm4/K
KUTqMdV+7jq2Mmi5BoAd9gWb5eBTdpjO1Coo6LqvxfzxB4wBM5zsDi7+NRI25+Ht7ditsNGTRjuW
0ktzUqOVSH8FXcEGnaravIa+B+k+b95aSK7xBXic9eliBwyas7a3H5T8JDG6GHnX6NniBASjTTmm
secofoAbar4C5KeM5QSIxMqb2rVArnyya2t/+0QzboE0gGgrE2iZTS6uc21DgGKo9aKmsrnSOo1i
hPzmN4pQq+FL+w/Fi2+0uEpOONHgddGTb5Xu3RlftxywztdnUFlE7HcdaJfbS+YbqECQEx+wZeCe
w+zzr6IP6fM9j56+HevyNyA4R4mjoabtA3s+WtOFFJ2bGKmqe9VJUs6AB3WcgV4UnlzVxXWi3+U3
ZMZsQnrU3PKbmMeDJ+gpHABfCK3l93RBbBfzezr5uJNBxwDdNEa68pXXXCTKgOsnwz3Azq53Odps
8lzFT4AMgcWpNHW/R9Q2bqPZKqjd/EhiWcpzeVnWIHhsGJBezDba04wJml1s2ZUmkDVx3jnGCmCa
YnvgLoB/PBRl0SBMpGNIu/8tbRaQjrVaerlEAcGEd5KAwdtcnoPK2TFekSBu/BX9fv8O24pocUpV
1z2WAN7RhRAboAjLkDbxCvVVqRNK95lHfchvtfDU1U5i3dxcuvKsug3puRh6IZqvyQb387DWRORM
SHMSKWYg4JV9yA1oBow7Iv4junVylQfoy45TQBr6ScT4nYGPFNoOi97Zm8usXIcrRTH6X0tAdA5B
uH5gLxbLdMoXpbafpQoAQ1CebsO2t5pzXRJiTR9iPI6GKe2yBJ8vsukTPXKYCWLSUm6A3k+JwAel
bnQ8LhYQVJPB3IaaZ7Z6gzrUs6pj7Q9N9Gf1x40zjd08YOaIaoQioM4SK3DYhKx5BY+8vD1HA7+o
bQIkztRUYl78c+itCAjYLNetvDumUpacUCRpa0RFW1Qep95j4k0+OTLl1nL7QNT+C979VNkXvoHA
hfSmbMM9ogkapRvco4QBfndab9RCgI8RLHoRTwz34LITq+QhqvDK2f3XABrtJAFxt76Jbqjtlsxo
9NoMAaAsVqzIzXd1+SNhUTpStjt1FyAywrASJV0nFafFgeAUgaH8c9yPz2wkGZExnEOlSExY+tL9
TbFBvWGDvkBazRUcgXIDhtgbOI8xoOdxC2MkziFIDLQNTgggOfTO+weAmij25wN7z6SsRRwO5HRj
1Q4Ba3zPzXzQPFNVqEKEmbRNniykNYnezo2V+vb3Wae+rg1L1djYljkuComR7ALLOjzjuIhBm1QP
sfCNKxS+rt0emN+gOA4POon7gJWkQB759L0Hs81QTf9pJHtfrRxCwstrldcljY2f+q7DjeLAm7sB
YDAa1ELVp5ouZQSVWYlii4M+hLJRdrQUcSHiT2/IoN84JllWIdjaC7560YwA1RIqx+eUE+t+bEZY
nEzFupuVzfPavwJi6EWB0kntaQOFS3N0hA84Z2P7luRXb4IafNyn+WJC2TF5Hkugs4pq21Xvc6Fx
Ywk+nZRw3pj+SjhFahwCZAvDaIdSXT9Frye+2UquQ6iGPC6nahG+VqWNLknH/z/Ba6JTyPKnCjbP
0NaKQ04ya3YwJVrDwgLxfpZj2sL1S+kX10HUPvaDQqPp8t3SPhRjLhwzxzaEUNMRYS2UKrcQKSPQ
OE7/4vaUaGe/YI1f6RZDsm0JygBFMAKS97WBmB+UiWvnNy1qV54EajN6GTkdY0AjQi5tj8NMdfWT
jppT/gpH/uD1q63jm2R/97H8Hul3GmOAsGj6P+Pdzw64TTtRUB5gPmM3Xp7bBBczkRl3qz8Cau6m
cI4iDf/Uv/6xvqDe5ZiytiZ3FrRCyWH1I6HQtow+p27ohFF62EOfXOViBvSng02VM8lb4qlmIQh4
sUXRquB1OepTDryzDBfSvIK3KtNOkgynmHCOMZo6hJRY8vx1KhZJGUPhBZCoJacg56dPolYcjPeI
oemCQrmhRAeZfd/1NPctrj8GALl2TrCPsGG4Fa5ExNTZI0BIjCyXuuCF3A+hbH+a7PcCNSq0Xfuw
cCUjKqnxtHFVISsYRXv7SVuaLJGYh5Xz0NUiOmmC1g5Yslnh1vEJjyj4vxvfq3jr1FhQxRnJ2LFD
KJXJ6nUG3uvxgKlOolGfXPW6wVg2VKOa0rCaQxRXoMxIPzeCBRqO0PkBzEEzHtvpYEqhRDXYDJdp
Kz99Lc4183BY5A/fKyPmd3P4fHAaz7AcwhO/2jxH5B/v6f7Sgj6POiWVvcZSverIhGhiEVwpxxCl
Sq00+mTsmI0BVZL0uo0p9QZ+jcjAZ6XNAkco5MuX8mTF6lRU8alBDN7oUqAtPTcuCab2TrBz9zZ4
IBBWnnyaUiB5NdG1a6m0omzhcritrUByqjFPznCOcQtVTwpi6sQ9IuH3EUKq/3nbdtZvmxV7aRZs
2WFvf0TZegpi+AtLGfHFPqvp37SpkB5Oxm2vNC0lOAzHyxKycf8fdPw3Onaz8ZqKutwDkvQkh5Ua
DqhHqb+528oE+Zel9pWzmgkcuGSNWpjTSlLvktpCuwe9qowqIWvRp96iNPq8dmqL9L4br52vYHqV
pDprTSYqn4Izb5uxSdDjroac7ShsVFL+9n4/gcZLKeMtFw1lW++VNDm8PKEcL9OzyexiBYVPNNyF
VUTWQP+/pynfKSWclXwPZuD8ycV823vIP2KbR7+RV1dA0O0fOrLNsg6ROnIdOstTTzOfDzbXGlI9
5BTogujHCn/aEgT4IVyXCR0nFYu6FspNujwl4S3rEsWv643U5ocEI0Dev0+469uGdT2a49PzmjMd
afZluh+F9NskZltZUtBuA+jcewLzc+qY/3+QYooUbZGWksbeOkqJmnfP8p4mLqnaRA3Ti0tsXK2l
8lzQfeifY8CEPDhGbevUak1M3GcXkYZs/JC+esjmZ0hGE9Ru8WIB38y95pDDXpjrf41HN61bfrrD
qEpfpsxlZCLkTrgzpVctOEuOWsHpGD1yDOZH8vzYuKPGx/eZgNXLEZ3D5JTTcalh4exzBNYicpEs
0DYY/idOpDcY5VnKw5XFOcmdnGX6PHokCR9uD94/ok2QzCty5UBHen/JTNlvwABj/vWXy7pr8lcJ
I6z46GDtgHijceJZUMazjIBy8KOhMdPztLdunqopu0bh2rH4ip/1SXTkASdl/aUo01Z8c6/y00lf
WoT9dJi0+rbIt5RqtCuKOJusj7AQUkh8MYOIAlZRNN0wuO9T22+WEIRsvpVK3QscvRQVJBM/mN8N
anVI5C8vpsZDE1tsXMkDNsC0/Sm6vl5S3BfkznEpoBVY0YWwHyyb4XvK6AigKYzOOdYT2vHkVgrU
oYIDNNidDY4GYffcKJKy3rlr0kpBpkowggNzEgthCkVDQBrXJrTcEeUctQR8m6opDV/4kAtc2esI
qxgKPQHA+VVI7xIsPBTCQwAtZxYjnWnXvNi5sGnNE3SbTui5/cMghIg/Jng0UDDxLOrKcuUA/vqY
BuDaZKxtk2yocqHFSqVmMGnzK9M0TRqKW5gkII2rpq++vlbEGl47lpJCSnhRT+vL/ledwVmVOrJL
TFccgseEz4f6B1sJv1BF7/n+2htvEVZ9ZhHPmuTwpNi0Cvugj33K/W0bao0L/vgZzoCV3xjmvLk3
qKMEFqiStf/mUwrp0ydSe3XX+IcFJK+kdmAspZi2SuFm+qqId3nR7o1LPCsPkkUvVXsm0lzz2Rcz
SrevFlgpPvi4U/979vMiNXDDZnGRg8qXDoNtLTF3G4pWyBKDQ3TIiIGYtpKSZCvlqgUr0fSJ85bh
e5xLT2ekyFMppENHly8EyMFcHRD3vaSbeY+cRNsnsNeSlzsi01xbuHZlbUgjkJkLpddpzJW2rVxo
MfbvEld4G+BnERw9Z2JUAFA0Ka13CFlGLZA6tq85QJhnQKchAu0T6cieu0u43IhF1q+EhHb7w1Ac
2pmHqqiiGTviLmpiOekK3VHYQRu1mnwzMX7Alr0qOAvioqJu0a8uHuP33/xAJEXNbI0Vq+GgNOg5
nnlOxeKkntB6lymzpu275IBN6t0koyWbExo4uGBjMXWg4f8xilcCOn/B/CjHmmi2AUDoIkIz7zlf
TjS1aVNAmFjFe8guA8TWnWk0Bp2zEKgu0F4VidlnVDP19VTmJv8Z+1pWVXxu77U0udpr3zLzBgPF
LQm2dRLvs/mT+1P0wVH6AO0oPkD888xf6RDIuAjiRe0jcG1csOIKnAVUFv6ZPZE1iE9u7ov9WLz1
WLc++Cll+4kOAqrdXvEHUInrWLgzobzfdcgtRc+jonYu+6pAyKJgbDBSYC5Q6ZKt8KA3tsBbESx3
c5/3Udpu4JgMuTSWr6pmtqk1ch2hMOYYnqt695G5FySUe75b8V3iicX83H1YJoEJ4nCyQ0+HzwHp
yi1ZDGIzzy3oqwofp5bkg1kG6r6YsD9VNXcPdyoleR/YISJ7UwHxBmXDbphjK33JE9pKKlvZAcaK
kZM7WWNUmSzafXD2JYGU9OW+kpIE4qFqOexRMRTQQ7G2LsvgYu8/WKpTRU7XGqX//T4Aac60B4Jz
xGgc9ChYVoICPZ/eCnXq8MYHmO7DOw0j8Dt90hWTMCpTyBvPCFtCz8DRla0RGEfgpS5TEk8udQxm
fMdifeiSxmVid4DG/sj7gbAsjrTDPea59VUvXMAF434Tczj+uHRbmz5Re7/p/NAAPwdp7FQ1+vaA
ngOzApSlDtVl9lW8YUEuFkt0BEv5s+uDo9pgLsJosaJ/I9zYl1YsSRTY19MeOHgNQ24wEFFiME0x
isuxZYm7Fzi4X1l6FmnaLL9/DZndfXKjY8OxaKOzM+BxcXEnDuECB2jgBKeiPp0q789S0g2pJubD
gM18WKHVgDxOLNztfa4PGVwcDPtNTvbyiYZGyf6V5o9SpT1bGZXdMbDfvxsqMeKjZy7Kt5n+6UPC
jBsQrDNENuWkNKIh/wAiZ6aSpDPnIcSdx4M9DpTKiX/LAciw4d5xUnBZsH8xjgYtG9JjQD8TgAdB
q11lsjVSoFSY73llorarOR7qdH16DfqwdsjkqSjHSszvaQVbud97y+KjBZOtIVCoKXCEGdbFzRrK
qVYPfi4NvOLKBtjtKx4fhU6o57AetFPizDI0HWmOO3+efM8zIBSgxyYbxAcu38UmJA01qKLkbQPE
s0XZhWJWSJbBz3XOZj0J4kLk+UnpqPDLvfWr+XjTwlnD6VwjtCPX35MY4UzZMS/bt7qWNmuJw/ZD
dePIO94X0+TBeT4kLFce8Y9zySkN2qkH81gn7AH8c4EeB6T6SdHHKDH64kVI0h2LdYOoOSTDGW63
sEwE6cjP+Dhm48PLDDHDAyOEXBckSGMjy70SsCzo1GKwb7Ah8ehaeNjw5+6zTl6jXejvIeNgtLe3
abSxcPHHmnV8wwGqLr1GLjNTm9OuhkXgRTo5wwXwEHrxgPXHnfXQmvlxi7uPpUd+JrvBO5ACcbL2
efMP1OqmTDGsYZS70667OGmnaPoSRKrFFDiJfl/nhQO1B6wAe/rcv0WgsazSvQVXWuC3ICfC173e
rOGpH1Y/32DXet4HSXbIsqawHh3nyVCc7Gm89ojCcQuVPbndG4LZTvAQcH3UGKZyVOXX3tNzKj6W
+DoVGV3tMVcOycpn/tF1TS3FWwOlQiH+qNZz7TDEinz0oXuFH9k6aSx9DFFeh5s0xMDKl/tCylbg
xUTORtKJTDxyvHhgEGZu0KWNdmIWDaVtk3fNEiZwo2wxHiHxE6UGusPzbHchWMinthzqJh/9dDUC
pPPG79JRbgHfZGtIzeBcOqqH9nVyLMcG9wBI7GKReGBW1pyH8xKealT3L1Oq+L/OY1vCv/G6kLm1
uM1c4fwWIxxyxYM4AZ6ctZ8IPmKQck5MeNgHlMPL2eSOZNeOvkTMrrWOR4FFFdN3BekOyvPDhTH/
Le8bAOGRdAjJFS0MZ1/3i35xdThqwVV3ERldIXUR/pr5bX19b9KqxtP/5RJIFNb2g9gFOfHih/nM
sF/ZkDnsY/lsPgvf2eRyP+3/N9p/oeuNLLLqGWL9oosWg44wEj9Jv1dIiL2OVTAjeC7uw7ARKnsw
hdrZgQdpFr8MKEUCZjNfAEufknC9LBfjrXMASnY5kUgoN0rrGT30XzoanN1SFub30AP3kpjiRJT5
dGYGPlYOJZ/YifXJ2uV7avM4KBfs9evPNoA0EMtVmu4upl2LKBFIi+yNUHH26Y+nv2TB1NDAtrIl
q4nzHHuzVBMA6wm3IhzgAG2v6OBkweBSISWr6bLhCWqQc/LTBLEw8dr1FlfJbVQLwQUz2w+YB8xk
WFstsJk0/TUCvv0h1ZN9d9Ex5RJhe/RpoWcQTmphx2D7wltJKRWvv/oL+neL2KEp6xeFbgJXhGlI
jXz4eqWS1AyIOjebMEw8k/H8AW4B90ofQx2u/SJRZwH1Ub9MFmnk673NTtLD9t1LTowN6syy0VsT
KYNpvOepscf/Nna6Bk7oOt9koFyREkGijYBHuuYFDy5GBOYzVsJ3F1lppwjzynUpjRXcOALwuaRR
9Aod9W6QB6wIoa6+MVTqBWSMyWoyEtrBBNTV/lGf8PEtnEKY45aiX95NCCTeTW4fKzxwyNnXj5W2
U6M1+uz7OEtSGsqSw0KVS2uRBcLzVGKGxuAmKnQeFf6d6yOAeZ8idI7iqGAO2QddOoq+Al1H0olf
iL3IiEwj2gl71PjAOV09P++goT984woNdIe2XN2KyvjZN7ZgAtF7zD0lgiJhhTXorN7wmh5LToP+
uhSdxDCrRtv8ggLak/3PPdaAJ64pP5+/xVdRcJYMrXKEHeU4Hlt7vfWZoOACpKnUuaw50iwcqZ+l
qHsUAtXIBgmS2OMA/taL3U47/cj0fMsqwwUJEmVy5+YYkjcFAL1fb4Tw7SxPUFuPy3yqrbO5ECXh
lcdR7jGyyrhQ75hQsD4c2+jAqCfl0O3hY2HdWGo0ljVImzXsG+Z+EkcIidzmYyxiI17TCY1y3iVY
y5QtskRE18hRo6mwugRrbNtkjhnBSn3rfOQKzYWx9ggeFj7NILnqwkmiIsEdtMqtU++kwlQaEoin
9wpDpUdy/svK8da8QP7XdaobCe/j5p22ALGYT+xeNWtXuBR3rGX7V4pgS+sq5NTFwtDfPP20JCwe
0HJqTgWu6EXbajBNtC8zwKqbK3PsAM2bUZVxMdY8h9rkTOsWVZgK16yQVuEiCYlzlvc+c1woD+dl
0G7R1C5Hvex3RVh31ySiotxJ1JHhTTYxDV1ut3+2H/25x6XKZgFVSalZHVFvaf9pUqIrP36OH4Mn
wyFxkH98a23HCtyygKtRjFg7YfRqubL7lkIAgdODGlF4uiqqHDmCyKBQ80TTyV5XQZ3YQPXZE2eW
Hz9BucnmcyER3Vx+RowXpimdI/xHnFwzR/GG66HNP1UUQ80SXVGJv4YdZO1Iyxp5tb6eup9q/cQy
xAr8z/yF6KaFeXdpkPlX/ql7RsnfWmb26I1YKQXCI/58fRXbfcR6Lmz2iSnSu5Bzo1EJZBOLssoE
F0ozEiZZDO3bnTeY6g9s7cbPVj5SsiKRAiYN7dirrYsVvCyKf5F7SnGdFs0Pmw1cw3Odg8qjW0ax
+MRmFpxx2vYH9w+aTrUiPQ+uFIBpwQRVvEOX0z+TOl1rbymnRdV8cfQVhCKmCcv0srXiTgIxzai/
DqLdtkyJ5I9M8q1pXOqNV5PGaeIj49ySTQCbb9mHgu7fVrL5Qa0FosKqJ7cogQAF9ykToJtyxvLQ
sUtvu5TLipvBfUDmWIRanjH/9hIvjpyqxUIYJFJM8qwb+DXBTmMBG0Arjb/ulFOocgTsKTxMeP8n
1rVchjPgwxQtGzhrjuZtr/kUclNrxPTuvDakWi8rAnzCpuUy8NkJuah7TTrmpfIaFQHhsqruOKKn
3ifXEMyFqj8OqMH909ErOQWZVR8X9ZxcwXeMhrw+6Zh1k7PSJlH49wR27mpWBQ4n/bO1O7nWiatE
vExODnIQlJK6YP0inG0t7lzHemzIDb/P9ZUJy5aNqfFhTIZcPASbnt0q/op3cPMfXWpiiAdANuRk
jpWc9e2dupNkhyxdGA4Gq3/+/rXGi5buW/QXU2INkn/jVPue4V3pDv2rqPJjN1niiFR0d94ftPje
NvE5Gp7SwbNcYAqhfZQ0LKzVrWIbmCcWlhqZpwP+DaNwdMZoqNJwn3IO0uvGiZPwy7kXWUhvjmlH
cBr/yT3p6nuaCGgTEg/9BCVpyLHOgJuR5z8ZEOfV+5RvcweIj+OHNBkH901A9hFCPyAv+rF8j/Tw
9wFvtrl1cm5ydCSmbwCfe1mYeX5sctVzrFq4eAhCFQIhJjqP8a2aqlMTgz2eFCtRHcPu6GBzl9bZ
m3qSnnCQxOqQ7t5PWRnqytnyF5WI8bKGlPPF+KnRAe605EzpV3kdJnUnhU3m+BCOnuuyrJ2Y/kIb
AMaB+pyYbBpw4u3lD15+6tXEtq5IRJrqog5i8sPzRvXE1zI+wF6VJ7ZmSHrjw6C+Eo9NGvfcoFXA
eqceGLZGrfeuUy/liynzL+HxPPy3GttbxkzXKYD43XAze4DEbQBfxrDUE4+zhFWl9OeCzeVGO24Y
IMaktw/hWT+neiyTJfHSo5E4wAl8hN0pctiZzUHMGxz5OThgombWlTqzWfMkZ4Lh6+1M4IZw/DNL
5rbPP8hguocB14Z/Nygl3p0qqswwHqdMRGBrIfrPYiKWMUOdS2UeKZLrHcgEzy9LQgRvcwrGU0Lo
3uaY6nnejFetEtLQMnvAowLTonqRTPkLZH4i090uKVg+VFT8eUVPkrVptM266G1bqaOQdEVT0Lo4
U46TaEAASoAu/LHae2YmaYUl5HkQE7aa0TJTRup21SblaV/prACQX5+L+52cuGSvqzZ9UkiLb8zX
Bab7jrcF26JXEzLdyzDwGErp+ZYBB7y6bWS8AHcJuzBx4WX3fe0hrvbrY7DKrArNV+N3rmS+22oB
IOQYSJB4GaHKZB8XA8PMvt0xDbR/bzorsxpqTf0IJe4NoGZ5Y3g/K/uWg3lPVnthjPE4p2c3N52A
zcmQwLfKfTHa5hIpgahf0rA9QW53KVFBolcBSek7Dv5zRZBZYxo16bmLhFoBTmZiuEHheAOdcurT
BI6Wk7L42uN//t6CcsskGEFQOP9LTwLSI06hIH/k0OvWQy4Luigz1F7ledGt+znuuJX527R3HQpa
s1uN/Glx71US/MjQbor/wqa7r49hUeuZRLIepzQK5VuvxSJJjXVY/B7WnNOU4GlhpGpPH7WcJ75v
UHlgG9+Sik0PFXkQyUSUu+IanLWHOgk8zAcBeIiha/DqEc4OoGPIhIezFWTsgiXKvc+tOrVeXmc4
1ElbiBdxqdutOX0nFEWmQVX8fhBWXDwKTqStbof4j3GZX94/HMzJuWirYqgeeMyjpDSaU0xDAxHy
H7jDRoHzPz80l8aojNJZUJJTTJZwC4jTvruyPTIW2LLV+qjzooC6SmzpqGasqxc7SL6ppK1bHuWn
PDkmVG8J4pvBfoCSh9xF3Yw08w34PonNbGBBkDTyQgBIjWfnIm1AkjHLXGI8YUaVvSWjorat8jIg
IUgpbaOgzO5nFJPY4ETaeDZTVYrSBUW48mNjpzcbJ5fzC09/ZhcPeGtvElELT7I7vcfsiFxdL+O6
R/LytTQDEhovbyzd/e6sg7i3r8QoLiQc5HRXcQBoU6DyO2TBpz4diC9BueFRojExNUtdKwnHz+RW
SWgjZAwY36YUYn3sCUMO5427aqdS7mhp0cbZ4C4Vh0QSBBbpSpZwmDnNyhLTDawPOl2JUciozOYd
hQhbR+rw3VXhT+dd4uQxc1MnaZSYe0tmQW8t5BL7mG7KofpkEBNAp6VX/UBACtyPRhVe7Xt+PpM3
lvQ3Hq60oCS80wxOzmQYRrhwGbn4B4w/Jk+JF/BWkbFqpKv2dMUfxuZ1kvvPCiF1TgjLcTYOR3Cd
Ng1kHsnn/b1u43yDwHzphpkVsl2JCwYsOHFK9npU0oVlSio+5I/rxaw6dYVVg43qAMC+YhoKpXq6
Xh7On+ZdEMq4IpP6iDLlbxaxwPge1LWVWGOZUvetkDmqZNGDEVk81qDHW9WzgNCohKJp6x4DJRur
JW9Nf0X26iOMVhLK5i+AyGZpJqpMvUTcKfCszncPMlav/p8wXnqS47EROBLkqP3e0OtdXqzcUUsf
QsqvY3RzJQYWkJkrJDjYyd8Qb85kQxpOfTp+SGpmeCCYAagwDivdwZty6D7dvA558ttJqZTgS5g4
zsChuz6nFSEnBQ/GJ19/H/TRmF5R0cmymdBK50/zqJL2c7Ew62GUtEH0mP0Jvf9drIFd9Btb4VOE
c/Q9OqVEkTkYrQvdxOliQqZh/jFMhclKDJLwzy1vZNreQTd/6m8lwaSfTJJj5SSWn/wqVpCy34+H
V8yZ419V0IEnb5FJymMrGnvYn7JjmdrnOeOXNau9636yYPCtqSkZzGmLnQU+piaaavpUU+c1Is76
ZQc4enlBLy6eIukrchoxLYvNyNI0wUzcqRQaeVYBG/+28S4+B8C/m5k5wlbhLzvXdPp9bQ5NhP+I
RUi+XS10vKLBk9s9ants/25e0nHRof6iALwctqGi6jTCHayVNzvDUbbx6OUc4M7W5yJg58rdvNWZ
G0aiOuwUQyVnpxR0UIx0GBVtVSDBMGviNtx2ydIUEu1Jl6QPHUy7RIDauSD7LXfPiiP5Ds4AarN7
VxxwTgFFIC/NRtr2DnKlbUxtAGeawvaEhg2OsOM4xOYXNnHbmpThEvu7pzJUsMHa9fvV64yY23jt
BU4sWhd2v6RgUAsjgoqfUMrS+Ieszm3MXmtFPw0jxlWw3ijvLQSEAgiEmrQdb6JXbNP5Qx9AmoO9
ag31k6fliRyQuo87B6QvtOSYC2zjS8dYy0VqGcDNBldBcx0Hxk9d73xTGQ5uijqGLG+jTPvMx1UV
0pnoYPsNuzW94WQ++Jn4fczT+q9L8SrRmyBVC1woZE9/pVGc25ZuJpoKeTLV/oI/ZQ38zfGMpO+1
crElgbzUgScZYmspPqvB78BbZYAgxSEYTJyrte/VpoViadSYmJ+0+7EIg9sx5JKRjWiz7tC62gRD
+hUpzUGjBp6CqTdSm9QxgSvJBeMrYugOPToP9/06jOWRKRqjlhwRFnIOYtoDyD/QdWlEHBeQbCft
5TOFFDp44FeP8CebenYCASKoFhebgPWvmbPmFyzIt6fT5YiH8FNBzWapnChxOEkGXESjc4k3FQsK
wi4RINKjW1q+qu455uiViz/SAOsx7Z7/HCztZCPcEftAHur9LX7wi//HaR+dS1VTl4NypB0ZUYXZ
vj2eiMohsx9h2IBcBOUhzRYDJONdGuImwEGaEf/7pf2LoOLQyBXTEY3G9nqvEam0StW7RNIMmry8
G+W9RhDjmPafrqbKTgq6Nf4oIKGRrJUwW0GpfKytpmDc037PTQWqW7CQ8nrgrzMhZF5caVlKpFVg
WUYW7XKhHcmKcgc/5am95MVyz2curS2Hbmatbg48UFYiPZSGG/Jl4Pm2Ct15JOx6AIWFwxmi5PpS
SW+WgwYhHzXzr/BSYuHhBgWWkbtCuL45w2IU1/i2vLepUa8egJsspC2qK8aR6dTzH7vTyRDqqehV
BlICPTHfX2OvO+75kFCebSMs6/eiPv9AqSYgvBBcuW1wDNL5B/iwtV5iJn5AEQo1HO+PUEEbACw9
HvQBV2BPc6T4PooY3iQ3HO2ZNvDMZ5MKyUKB7n78s0nomUcg0eip/PakYNoNijwmlAwk006OxoRg
geDV9Ryn9aYY428vCZyIBhBH3Momn/gPRiCGU/d1QW7Nm7A0+KDj6K+hBbGgWnm0DNBKwrzjLq4b
t9YyC77VtfMNEPjoIluMiVOY/P/v9OnVyfTMk/kHYbdxI+D2UBlbVrs3yh4RI33rmIcqLveu7DMb
TkdnBNCP+ZKxoAYP7wBibD/06Xh5v/Xs0Yrbs9CPqUHDbIZIRRqdBYxsDXFBWAhPdsnZ5O8eLPFJ
pQAvUYWW7rzbJVi4GOgiDGk1hIi328DjObvOqmTEwp5K++zt+Ctvx3oXuE31vIZBtMkBI4WFwmmF
Jsi9dnOmkWdCeYPrQvXyFInH5UgtvKOvhokYTTHpW6XPNm4HOapm1HpKV8NNBobUzXwiPe9Th4D0
jwX0BK3AtK/zhURdb/hBLorWadx7YRo+zXbP7Vrz4FyrfcvwQQO/bNMQBhMSSOk+3ezFctxF4qmc
Y02I9YsVdkqmG7/8P9bH3cRx97xs5PWUV0S9YwepZ+JQ28AgyT+pREWqBXCn9gYcdc2dJ4+NERnS
ZreuOaSo8Q6WqUfxC5pXf1JBY5Q2HHbvTGOvI5bNvH0cvfJZRcbr0bcLc3j8c3gB0kVRrGjG0Q+p
jg/WIpA4Xz2D5jJ7GWyfx9WX4nC7yDGBpk+aTkFd74eqOomzzQaSPTP2C5wrlKBJ+xBKDPiXxaHw
RfKsOSUxT/ScfHdk1EYnhaKNPYTE8BRgTlkGm4eF19ZY1S6i8lbvr+dn2D2IiopoEMQ7jlSkyaje
aLwC6/chq7j1UXs9SoFJO6yJ+8qSMVN0fdFm6AV0qFZmWnZBd6G/RpNDU7Q5gthUhd1qhy+VGMXq
fJfd/jhRFB9b9uvISgP5k/jeaXPWkFFVtEQxZZ+yUW31oAWc7z9nn9Tgs2X2SC3vgdYNG+7QIlWz
YZCIFxrMl8fsFzpYOQdKBKHY1CgXZ760NGeKI1eHXKbVLwgwkI2PKU9amKDMyNnZS8f0UmXYxBeW
lb++HUp07Vp8LinzzYG5J00BfJVZKEJ5sliw76RMStj1j95W4OHKHghn7dZqbFmWXKPe6B7wV2ff
gRpa+cp3Yi/g682cgTXLfcAOa0FD1Y/jMZQzOCP3w/dEVjsPaqgcIsCAq35AyZKbkntXsizwKcVH
t2pOogqNUECCwJr9xVrDCqwh7svhk+ezhzwGaBWGB2D6FJwEprh1ati3M24ErQF2cwU8y3bTeAoM
7J96jvBg9uUm5Y22fuzs2Lu7R9Qw031b+lsTZ+29t+IhvovuuQAQT41HhsDKf06TnIKyXkzi3mud
j2qi1OtsXs+HID5JGe7bJQ1P+erlaof/6LltecVqHLcmaTa5Q3pHrWPMV4PizgNFRFxCz/bY1BUm
evD5fZ91zFXZd51C4cy+f7nowUcYUAW13VC4qenNfSBSjnCgY7KKh7GuWkfBEiF4+wj980AMlKQ+
D9xqR0FQqMiKMC/BEFXAxzk+rlHlQm5bCyEGtixaddp/wXyso0ZldXoqQzlARmELJx6uygBJKU6p
PqvNUrjqq4PFwLuvexUhYjH2YpBKsuwiLMSfguPonirh4QAGXVqpBifkCtdmhANYLMDzhscvcSSM
X04roCvRekv0BFq77hudDOJqm5ZZNz5MLh0FyrNX38Z7HqP1RAP+4pymmFWLSSOHeU7nJ7dZV+JT
grWI9lbAJ7IXvf2ZJwHhHhYNd4MOVrOf+uMe8p1YotrImqzxTY0jarnei7UWB3+cjzC4OrVaoMbN
hAulMOSmcP42Zu/XalWASxhbcSPU4yWznI8ZLA0pbhH8T4UHnsCEUQdnwLZkgl5l15X+CJhk/8V9
/5alqU+Xnr0lI7jVo09yZsWUtZaLi0Z5/pQUCGJ41p5X/rQhVr3qAAtCox9TNq3tRikqTHHT7aK5
h2UhYSPKDgMY4ZIyCzcfv8r89b/SFw/034uwiyHn7T7XiFZ+6rx6rnIKyDLZ4f6tFhmePf2537Uo
VhYtSkFX+l8qXLERiKGCvPEa7Tgmhn4OkffNQVZXrCcUMVkQ2+jojA4DldV7wMXiWk/dVyY51Hcr
34eTRsiq+eub4O8FnaUF1vuyaGZPhaLk9KY0RxdcjlA/k+ly4gOfVSIjusN7YRJED3qnlhnOQGwp
emSThmPuQvB2ritb78TrPmbEpQMbx0ZvMees1wYDqhNKAB2PjTyJJ+Pvnaj8rpzDhI+CR9fSZQXS
RKri2j5AF0jtKcVBlfAYU9SZOIPy9Y55KRIPS+wkbbhN7I/jTqD/7KKRbKBhYT4DhxJUAq5qPGuC
8xOQTVbWh1YVn5TgkgRABGQBoJ67NrnzNcRuGpwP6Z8vEs439jR5ppt75IrKLVLpH4bI6yCYFENH
eAoog3FcMYiaFn2xiSpV04+jc+Sa9+xjFkKlMtQCC7Yl1UV5Gw551DEKMCJRU1KDw4MytSs8J0au
ECm0lbIqk3+ERzXIEEaI4Fhq5lA2lr5MrX4yqcALHzGoVLXX1ReZQVOQHKLr17Qpw6jauc5FgEK2
ZbggQJRy2ZIqWxGJE5eq3eSXjsED/lGubxnQJdQipxCg9hh7jnXjwEmMGW+WrNB8MVwuOrRmd+Z+
WtPI3xYdjP1wmDJBnBvbtvOzY/TO2aBP4uSGUYGX0Jo117Da0mc6UxxAi2zu6Bh9n73u6iXWkQks
OBOnbTAhnqZrVZKJnYGy7FjRw1Lc7PgmHzNK3xNIqXqbD1z8LyIeOLkuRH/aUdIFWmnUgUc1gT/v
xsUo2Zp0eusEh3QvIEg+x9OBZwJYfNIVs6NQ1Ht2Db0tuWr3bjZRcO2TheYKc1xxVJe6hKT2Gt/M
8+b9aA7z2vZSURZ56JdjxZEHF2Q3+boSVAoz2A9GY3j+MSnFuqnxrmjkWMiqtqXjvm5hB1ZlEJMZ
3raFuOt6qr/72jLfLtadHyXIqYIcwUKjPy+A6gzPLSVGqZqKi/+cafgsgmDFdFzoYi4OVoz7WbgW
vooe47NnwTY53HETmdF0UBPfGzKhH4+WKstFkQ+YjgWURX4Y+AcWmUm8gs4s2k9R4ebLu8ChQhZZ
/TE8SnDF3/BSiK7YYmwvlHygPfRKvkER9VMwREmXOMhHaszzuhWUn0LoBW+DH9AUi2drfoo+t6n+
N71cyjDJlefYPf+wRodO25c7LSR4bg4tPb/UfFdvoPxOBIcuOHXZhB67d6C4ws7j2w5H0a+1uNSy
G7I41inMbNyEPSa7UUsEwygJgqcZXETQlOCwxa66DfK9kIhCXAK7ZVsPmb6yiV8bz/PjfVlbo29h
z48xgxHQfyr2QNftCCAv8MxTscCuOhonteUDna2r8e8eIQdT9kEL1uMXacytFgXftHTzR6lgBUZP
eLPaGHhyljnWY9i2lcB8BeKk9UbgPdUJRsctny+gnb/vqQZboT4THZ5P4o04vTjJNWmxDHMCAJrw
PpP0GtgNrMrGbViegiPGtihLfbVRnPUZg8CiDX6s+eED+5MPON0gwvQoRDY3/cxWgavLrE5epLQZ
kr0ZswD5XtnPsp4T3gCmAcp/HG3kHBkjh+WJqaiBuoXWBw8RIRyIGc4AdUiF4Q6T7XImFJHXuK2N
WonBLZrKDoOFqJ2K+tg2XYbFyLDXBFq11v//ttb22UqXa0RVe5xu5l9V3ta6BWki1mXwupiIAmWH
OjHE54GtINCBRo+OAhozZdJLOGRTr4Hwp06t8JSewvb+8e1NLPF+5K7WMWlRS0s2k3xaaOGwETH0
f/TMfI77iNfxr+40BKvYr8BrOJkdp5rUEir+eo/cSi0oLV/YgDSjUFaKVVkLG+UelcVHq+FSyl54
9HPxsYLz9JPDN7U2uzdSbdKRiSpJNZ8t2ARuao9XLIm65KWIuvly6s5bGoE8IbQRGYBxtc4Saf+o
Y0+OjsCNl4e776Y5baY853UUdA3zNh9UnLvmzokdavehE7dmFzZHmfqbcvk/DftUCKaeWr/LrH14
oZEuAn9MxTCEKhoobJeK1Wyw8yWY9f3Tbkmt6fYH9glS7zVcd0Z8RI736YQZa9ei7EBw8uS5hiWg
FuZdbYDVap/z5RBylKDtr7XCZpLHlKBTUzFsL+fzceMilMkYOYg7DNH6Mau/uX0Oqv1pgcQ1MDz5
84N9qgeMFfQgLeoQHenYiIJx8e5l8Lp7ENHjk/t0cYmeRn5KIBiVtbvFz8TfgP//vuYNx4a65M5z
pRVK9ob1qzDPhAlerY2mbTTNsdXcVJsABjSbnZ3NB5LM5lzufXnFFLYy/MtrnEri1vgGkKBGr5wI
mbEHZE9geD6GrZJJhq8nmrAKvqiPv/ZnaAXlxVQ9xPWycLuGrzZjOI74ctRDlBi7SArRDn/YARyF
RhoQoxzqG4GCCqciTPZoUHdkjum+n7oxLnZNcRrl+LpFG9Ge2peSL92BMFtzF33mXdxk6Yg9cZIq
37PXx+DzwVnDWXS06ork22aHPUOaORu7XgE2rkHEiP0SjKG8k6nZeXitkvsSAVQvzoZ5mgIK4XNa
2yqRB+r1uZ3QVQYrYQlJ0yYzenI5O48NxelfQlxHh/ysoF7JcOEit+hdE+VcO9JDfy/+3qq4nVy0
j7zwrUg0bON2LUDMliKkOSt+joJW8RUMJnITVf/cU+ZWnGks3o6AAt2SZgndduqf2nE24F/Ydeja
iIHHrSlH2LsRVkZB3fKZNeuTssdSWPAhzaovfN7xCeyVlcx4CLhCSUYdgsX5wQ5cP0ThWU1S+Ca9
/jM+0+nfX0tQyIOp4qSeSsuQ3/ei+c6UBE7WvwlzohnY7unflf4iYFPBK/8cZx1Fynkm5L1AWwrm
zSGAT+6cDejZuJq/Xje5D8oeLZ4jy/b9SvR5jx8zvI752l2apDmZLSLCKbqmV1D/Fvf4ufyLku48
d6k/KuoUpgAlSWxegBSMsiCs5pm64GP8oPCZ74tkY0o9t8dCR0MA0pXONJHeDsDV9haUbEe+HFYU
45TLNTOuofqFFlR5k3vO4a0Pyl0WYxloFTPjM4ZzUJwOI+Uuse4SZP9J7yZrcpaLii5MTm5JHlRu
gGGpAPhnVuJWOD3NENZLSTqZdrZtjTxhUlRmJGYHCVArO0EutY816luCB0Ge6Q8/LxPht8d/89cM
7/ZMBeTBi4UI6Ch30GCgtrroAnutELLNM6affZMzxfJnfG2lKTJB5aiIJq/H435H86UqNEU/Oo/G
VkwGE0DL4WYsiDvlRgIkYNMUZQC06jgUuWarQ/U3eYTT7ja/XSOVSgBXS5ZV3NeQ1YlqnpGe8JOI
DzojqOrj63bzJI2YRWLJzR6nIx7f58+0aDJsop6Ti8sdM2oWk7DbIYf46Z1r47dSDa32lqe2bf99
n8Sn7sOpfZZ7qaEwR7f0s8EHqJ1CITeqOuBPX0Rjx7rpHpk6x6r3LT+ZOCEhbdBR687laySXDB1W
fIfGhUKD4h5GJHddNJfS6zOsObte5Z/5ugFj2znzw47IKoJlmb+BcVDBj6TF4+ppKaPacOtvUziM
Pr4KqYn0apMZagKFeWtmvjwiyeDI+Q4HZhMZAAtIzmAJ7AU4/oyuYFHQw6D2qB9nw1dYaMFUSM7C
yHHwgamsy9+Fnuc6yPjZ6nJ2exnEDzDprrrh/dlbJqb+Y5va6bPNlMsjoysvTPk3vV5lDDeXsL2K
lwxvzDpmG9ITYc9EhkL6kosY6SOxEghoWpVDe4qv97Ci//NAkn0UCACe+b6dUvNBXkM1RlMO0rwg
CEkTtJBOM3rEvMm2eplyHKblGgqGl8OEzbGa/OK+1xjuC+1eeRISkL7E4GAvQIVyvJU+XkY2r4xq
/lTPBpn7RpdKJHqbFtxEceMngx1jWY4jnbPD4YLaDz7DSARcb8CwkgTmaNFfwykq379XFg421ujp
GViDiRjJJPGG3M8tBM+z6ewDoA0GcryzQk/XEO0GaPSgIfq/wpbSEMj3aqZ4U1sM6APhHNDknmPf
LEplUXM3UWxyNAwo8XP9Ytto3KqAxUGiTFjxxz8p81udnb/ezamDtK0+3flJTiDMNwr4ZDA0SSdC
Pemqkfh4JCZEzI2bdfv9v0H+9OtqQ1u0XBNiy1JxEZ6zodtpt/PJv/cEucQbtchr4q0qFGfKlHXi
ohmHEIZ+PlYyHC85Phn0d46pTSYh7pEV+ZwVc32DUub+FWm8eQU3TtGiGM+mPtiNOrZxMT76DGlX
NN4FKHXVewq6oJZCw2UGFOAzov0gEyDCA64yDcmSaSGLtS/XPqhbVx6h+zYBNBKhy0W9nub0p2dW
GzmjZ0mm42TgNsDoUMkc2y7BpVjdwNTl3NOU7TVIHB+cUXkpEUGm1WT8zcvUIZvpeBqnz7G7HeLu
NFDK0l7SgO6AwhQu099pc4x/2P38VE+lWJOuIhrSb8LLbp4aM8aKYLhs5Gn+iQNbBEr5ptw8GfmX
oi8GxVkng1OWrMwGYMLaiu2ATSsqrDo16glkkIAeDTt6A66+YB4ByEIw+G5CjGFMgUTZHTryQ3qo
S8f6Xk7jctIJYDdCHb8WxX0ir2Lyf55GLl3xIIWn6hXvABMOAlD9GG/HVLnK7GNVI0sCQyMt0QTG
hATlWJ4hHtw1l2sMM+oLhOzMKBCorOxtt6XHUoTQDKYV7hkJZA0jOsILv1LGGcNUnXEkLDPfNN9p
cPDW5mJX2uvoXTOsj5U1UUBn29xM5KbR9XJcAqvJUpOwH4XQnTrh7cQrtHmi/37vxkEcdqdC7j/A
IwhocacozpjWTn6RSPWyiO+Qf+rwIJWZ2srN78NoZcTqy56inR0Lk/kHyjRutOpEYpzAahgPft6A
nrQT3hp15YCl3yNW9lHmeB19T1C34O48O8IMJRp4ETOZwtsb5Li6UrZZtXuTm/G+F/JibIva4GW2
66wcO5QOQNhlw+t8H4CqW25KKu5ll2bAPreM4itBYcufWUSqWhXDh8pDef+NxyM9tVLVa7NRDtcM
LQCIjFH031KLXu3va50+VpmpiJC/BDHeVWcExcGoIDbZLspezsZAshYYIYCWCV1doyP19M1s8UjY
8axYpIJjf6uN37Ych9u+Ab84YlnOA9ICLtq3P+xI2PUa4PxRS3o1/AdlFS29fAETzuQCKKsJwCVL
dXzL2pQEtihzX949gq933Gql98+zlx3qbkks92zwqmYeOdb5sGevaBt04CLVPF5s/72AlzVKOIAx
LmayjqP/aMin2R9M/KnfFXyXVMzlhVhwZa9e2Hvb4ANt1f+QY0p3Qj+SxwkeB0xskQL8Yl/2ae5t
cbHWy5GeomTQov7LQwH7j4soYZnwaC42Xp9kEByZ4cXf4vWIFpDB21ZCC+af4HpxiQu+0DX8Orb7
CnNCMmn0WstTzM+Yzyzynj5LPQA8RENwe3HlRcIwdlS3DTgkql2bKoGJdyJ0OYlGureLVwaQYRgz
6u2tNe69+isE7KR9QQ4fQKz0f6naN5s4ZLwgmJZtzd8eiuHqGHovRtatWvrKMsLDAKh6CfUKdwrA
xtYp4rAl35VrplFSpo62m92EJMr8Ol0exysYRNKffnjeoHTck8BTkKmWyGH0fBLWeroOhf/3EwwU
f2wh84ox1oyOTFsr9kj3yiMfwucmoMgxuYA+7wWejIOyESENn04kx6GEJ69IMIIk6dfCXsOi9BhX
z2M7RI54gZ4hIrVsLJaBWp/wUcy5dX5zDHDSabF/VeB2kOB+ReJfEKJCz0I/ox2kjJc5iO5WCmWD
E9kTf6ab1lFYgxKgEUJZ4Xxn9GEUMTvYFpIdYax/QjWvWy+SgGiGYeTkQ4JkVra95EkXkK1AuVdT
u5oF3Da3dbNz91l13FgxV1D3IRQqVN52YTlXoimgto4FCR6PuLVz0uwbJn2aIR4R+QCBAEp6BKkF
OyA5AY+lvBFvdf3T8w==
`protect end_protected
