��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l����Ol��v^w ���Ʃ֔;i)0��D��J�{���.�v_	k��tZON�����B+�lSAv�HWS��"��6h
r���}؁q��%&���#Z<$4�baL
��zn�e���8)�_,�!\�3��r�&�nָ-t�1��d�/�������!���Rcu�u��z	R��>���\���ƌm]��L�׎m/�C��L��*�#*���Q�)\yq݋t�y��"�ݗx�PV[����6�F��ESߡR�	J���c1�H���M"�f�xB��S,�q�� "����ORN�C!�¥��x�Iao���h��hiAՉ0��lV� ��5PŒ�l���.����((�6���<F� ���?~����^�CNi�\�h�O��ANy[�i�,vO�[E�XbS���<s7�&�ْ*�.��jFc�쩈�I�-$�l�_w��M7��sNT@�_���Ŕ���N=>7�t!�g���4��"n�%^Ը�ɧ�2����2���$6�4@��gؔ�4 �Wx:��(�L���}7��-�� �~FX��{5E8��g��A��ј݁ڒ��b�f��%�;���,���JM�{�\�* s,ŬG�8����o��|�@�_��a9aæ��dyKi���`a��HwG���H&F9j;�H��^~%⛅(sDHz,=�Xe�B���>V�s߁�a����>;�@ަ���@�,��V*��7�7S�}ܓ�K�LY��m���}�����E�z%*�`��Z3gl���rgҖ�� �Le������K��,���P��4m�ކ/Q���"��5-/Ҝ�\�d��,�yp���־���������Q�n���'q��:����~���_Lњ";��sc#(O/�~6�F�����D$P��SL��c�F7��w���٬]�B@�(��/�!_X���_Ͳ]�%�42"��S�6��C !�����,WW�G��xl�G�L�����Yb�|aHi7 |��0Gh������#mG��.�#s�}�R��3F\6y+�P:����Џ1�J,�ބT4{�ր��Q���p�+��Sx�e��Cv��N�$t�����N��3�� .��9hnFс,b���-o3�!O��~����e5�9o�
W�����S� v�[�s�]QqS�GZ�46��S���<
`��T����&���<;P�`�����HhD'ā������{�}��Ι2Q��"��q��ty륩8�����\��v��zpL�ڀ�A���u��h#f��`.�-�Z�L�Wڨ�,$��10��<��tGxm$�rOK��-�t�b�HV,�D���N�������0����$�tE�b
����j4S�I*خ%�i�
i}>�-��O��C�5@���<t�BF�w&m���i�~��5��w@J �T�CM�������F�K�v�*h��:%$v�E	b����}�g�P��a�A�bҭA��v�`� ec��Fq�4ɐ�����?��BzDa�G;Nf�Qw���� PH��/{��2�@���,P6Ӿ�:�d\��aK��o�@���R������#��5��_�c�R<�d�����I�h��
��;�M��ٓ����p�׬Ր�0�����7�%֘( Y�&S/,sz[�l9�U�G��w�)���(g~ͦ&)P`ٿR���!̶��9G��`��V҉#���
�+%�fN��1�A4枩�eN>#��F �*E��G2����N?$�*��G�0��ƨYv h6�T�ہ�8�&gƀ�8�9d��f|�>^������U�R�R���wT��{����!<Bi/�B5iՙ5�2a���ʒ�}L�þ��ܗ%��qߩT�ݽ	!+K�LŻ�\kg�$�3
��""�Y�~����
(
S����&������l��L����	tt)fa�p��/|k8��PA��'���TM�;r�ƾ�?��������������4��Y�A�N0�(�����*e�F�+��{��P�h?��+ۭ�5o7��d
ؽq`A�����[���b}��:��H0&/n�/��� �ZJTS�i`ē+,,��i���[����]�L�Y�ս2a�N��s(_�S�oc���U9U��P�#P&��X�^�FZ�����&�|w� H@�[os�dӓ%c��=ύB���2L�Q�I�q@�}L�ڙąX�+*H�:��Ѭ_(�BP/i<X�p�U<�9e�P]������QJ�5}ҏ���%`|A�m��my[���?n1iG:.�0_DÁ�͞��N�]�txO=ExcH���RA��^�:_f�4�nf/
(3-��m�޺��ؖi���A�r����
J��I]���T�~�+��Q%Ť�3��������5�x[� \�Q0Eދ�FbA�&�<���p���Ñ�����vWDm�5�ѐ	z�k�|�7���c@�,I���.�b�YiZkfZK�$�7M�C�j�������{��/gb"O��N�oOi�B�PB+�#�D���qVP;H��?�a��P';���\~Blۊ?
�?����S���dV��']>]d�JV���C���hф�<wg��V�A�'Q���݁�LkXUI[��o?�=�(�64)��vYꨌX�����o�%13 ��_���)��^q���\��y>QZ�F9�/o��Td3X8�
��������%L�<s��n#0���ֶ1�2�î��)�[Ia*$c�J.ӟXX�)�Fn<�|z��5��kU���;��l��P��F�T���b�?i�dp̝34���R�����\�{z�F�X�<(������&K
��s�C��K`���Q�{&��v��O���������PNoگ#̌��5Ş��K��7���Z�����T�U����аs�#�1Cz�O�A%�U�7�D��ǄTm΍�?&2�mT�3��4�G=z��!_#u�9���ȌH�7\������ů��40��l�?�G+�T��R@�2�%a��A(H�RL���\
-�@g����#T`�N��^\Z�]l\�7��h�C�N}�&ԦL�97�����H�>���[�M�_V�@��3���ڱ�J��������2�����n�`@��c�lnی�t!����;�dci�&M�A��0�s�R�	z~9X爷˾�v꤃k��T�>�� �R��~V�s:|ӫf�Ko5(���#�e0�jh^��i���V�����ˊs��3��r?�� ��| hD[�2T>�Ql��S�����H��=[�2e9��1Iϖg����_���2s2L�)/>��'������ka�\�
5�Blc&�0՗�V��I�8%Ջ1���hG_�}k4��M�K6� �0������5�8e�C���CI�^��
��nׁ w���ߏ�0�h�7�P���2��8t��U����D:dǙ yà�M���@�N�Gb8�����4'�TL��`eQ��Sba������OͿ���2.^MS����0��$xT��ؚ��]'���Y}hRׅ1p�'U�w��-�}�bhCD�VD�ЈJ�Ȑ�j"��2����F��~*JQ�j;Eos�����C���Īo���Jv��\0r�f����n�o��8}�;���[ߊi?8h��K�qu3����x��[�{��n����B��KtNc�m�+JV�CK<����I{�5XSH���QB����@C���8���M��M��@�1sTb��ź3���Ha�)\]z��O�ƫT��u�Ӏ��J�"՟BP���#��R��Q٩5� ���Z����ޘQ���Dwc�v`���HN֪=2����oK���(��a�k#�\�B�.�� ���0 Ϣ�[�`�`<[w�&m�#;d��l!S\��������aq�(���7It�sF����$x^k8�Ц{�X~�8֋Mܐ4d�'7���Ewv����&尵��p«�(�uE�ѦtA+e�9ĘNؼ���K�Cz�Bme�6րzb~/q�?���d��	�P��>}�OS���-������.-O�y�!�p�O�]���#�3���2x*���{C���--J���Q������3���%�߉F�����zF}b�����������٧W��G��͐{��8��^	��BK�j�G���~v��2t��y��ee�'z����&_ A=J��o�_i6�t��a�LU��J}��WQ�)����ȰVg�\T����I�6��3 ���!��E����N=�n��)[c=�&���Ȃ�H;��(׀�*{>BIW��*�[�s���In{=dߙ�':�v5�m�Q��~�MM�q���5�j���j�͌�փ���v�l,^�%d��Z�;5��0�N�U����{D�Q�s�tI�q9ˠ�U�㭴:�n�]@l��Jy����O���V�P����آ���VT�?�bW2xnq
�����М�ӁBoB��N^Z��9yKr8V���q�c��?�0:<���+V�[���ֹ8O����]k��CS��{�鯕U.���)�捉u)Q������m䈿D�O��B���Z�|S��D~!8&~��:�����Y����o`QΈX�HƜ��?;3�D�^���U��(5iCD`ѝ�i.��3d���4/n5��p�j"@�L
�&T�ŏR7w�Ƿ�\�����;��5��`Y���@����~,�^�-��q$��{�}\T�R�/e�Q���Qn��M
��$<���̸���Ί��W��w�S����D6��:����t�o޳@���!)�i��h�W~�۵Ka��9u�Z3�\b8�%e'����@�X�����*_��5SQ��
PX�/*+t���?�n����6V�)p&��]�L�9S�NT��:��D�ގ���H����Z����,;ե�j�V-{o��Mf ͙rG��|�[`i9F?Ѧ�|鉵&a[f�0ƍ�����'�yi&vn�P:��������y���}"/��e���_�j�/yZ�9A�@�zd1b���x;u�h�Ƥ دb�&�}�&���W����l�x�ͷ2*�4���6>ރ�t[p��_	��q����ݿ^��v�j�d��N~��4:��3��2��Mx�ݜb.�����M_Xg_���2_��M��t�B�Sh;�7�p���pDܔ��0Ҫ��^�}�쳴�;�a��%�̡�N��nx�lcw.������`f��c��M��h+VϿ�����~,�&)d���2 ��9r[�W�H��Í:�v���Y �HnE�7�#���&�J�����9�o�yN4_.�x�"�#��7N��L� ��`��gU��_�k1��`�����o�=��	儭P8TC��2�t��V aY�����%���#��8E{�����`��5�<�Rɷ��2�Gc�T.��ϭ@���eB�JI��5�?UF�L����V����#ٽ6�:R_������*+Hz該�gԍ~���4���,��IJh�0rU/���y�^�8Z�qmЈk��10K�S>�GU�I�����:�$)��2Ԏ�z��h oV�kJ|�"!:�u�?�����_�hS�a�U��)����iG�[�I=���Șva�'g�f��^&�3�n@K`�L�Y�C��qJ�4�WFР�-��4�e�m+�@y��`�9}�pBN��E�F��I����[&x2�q�ɹ�����SBw:�$:@2Щ�`�������4͋�h*�2�ؑ|8`A�x��ն~eEn���:$qr�&>�i.��@v<����L�ݗ��wr�'�S�+9b�f�v�� �>Q4w�z>�k��1��l���w(n���J�����=�tJ)��k�{�т����S��`�I�f�fQ����x�5g�^�&����`��'����5<�����D����ȯ���|H�1��V.>]�Gw b!f�#
��L˲�4�L6���:7������%8�����S3��4��2��/P]���<nB��iP"�Bh����m��ǮW��:
�D������"e��� Գ��z�T���
���FW#���0"Mp�HA�	����J��qc�!3@�ft��O�!�Ł�F�8kL��i�m��xH�F5�IHcǕ�x��nl B�!��{f,Dpc��x*"X�}��NI� �&��B��7S��^.I��bRX��K��/(��͏A�̲�����Hނ��Iu����I����9'����v�B���u��/Ѹ�k�:h������\Il
��� ���m���\�SJ_�3�|�r�)	g]:ŗ�����pY��(�4���̟��v�D�:L3��ą6��$�A���i�kz^(̵�ZM��KM�~���ZT��g�8&sHdu��E@g:;痫C�