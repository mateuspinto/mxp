`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
xdSb2iMjgZOVM91/YfMGxd7pxFdSV1OFf6ONi2Nrg5SjTC+9wuwe6Q50jOuUPLrllu+MbgfjC7Qt
MUkJTNkZ3qXl2XYWImjAYZZspoCPpkp5XHnqOWfcO0sbpNKeNMb6bTilHlFuoJ3AFX/JUPsjRQdo
lOVtnKGxa7TfAtBq3XRYfwWxM+yv/42Ok2obS8qTJSvpHlauMCP5l6c7U0/jNmIBDr9pVwAlA8vP
gAbr7Ueap39febomL8nCwqVuviFDQ24IwRdsps9xlZGpl6vJkoE7E6n6Zsxk/USqa2J1qoWi3WWp
bcTla+2yMhstCU3ea27rt+o6r2xhXEcGyyJd6w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="EbnxkuISmHD22yA7uecAqbGJh1j6uGyHibmbwuEkVUM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9152)
`protect data_block
EbSlmEDoYxmBgqwXRxMjF/W0DFNLgiPbSDawwATE+EniWOaX5Ug6mkskyR+3Vf9TvTUvFh9V4h/l
2EV3QXVG3A1t50wpvrBQfBI7G9HGOZ/8rgFOdzwaxzb2qDKx7hQ6BhzC3UZihTDnXItYDvSF01b+
elxmL3y1sQPxBBAeUx4N6u5Tnhr8Cn5ezA0AZoTqaHvHBa9Fmvk38100p7kPR0pmn0aQW2BRYMpk
Cxll+hJ8kcP49qcuyKP7Thz0idLCoQXef9iNhKYCMpiHmAlTVD9mkAr8YpnrpC6gxL5nPqj8eZ6W
TXWMaK8uaZ0Y+w7jDBdrpA7R2U3h0js5WAJ4WrPeR7KRwMRczgOWhtaDAFudeSZ+hTZrmnTrqXck
zm19cVAV6LeSGcInH0h11sDLi1yRa3luSlhHLyuhm6RxUqifKagu9V98iyxpYgDfvbXEhSSUDaRK
pvp6CkljlCjZe3oh1pxCUglWPeXYZ2xf7An0lPTFr36dRldVcASmjiUbs6R+9UwGgBLM8J7U8h+1
EbLhJQLJ1Xy5S/g+0V9ujHOc4+GnHVlWOe90cOt825lECUOEVhEbhjKUolXLj8fUn1vi9exiaCvB
VA4GEkVrpTvsHUfaWBydVKpmi27kriJfJnjTIrL7PyP+qli8ngUiPReMJBimOEbJGKsL6SLYVftc
wEXl6/Tac0l9bpdgngQUueOsK2zafMngihg8AwknWlUZpejnGh0Z5ZDQ0hLO8/3N30YBQbKWFtY2
GaZwIWtX1Y1ZjYfvWlaD1i9eJyfKdN7b2SXkWDclTVym5Jzk8D4wgtMbvrHEVYcRM4nyz/MNOt4y
ITOwMOINWXn/FOXlegQhEjGGXNmakdq3315gWkxDfwoqIAe6V/a/HuOgM0PGVl7mz4hBeUbTkdl6
T6+NZFxk8vt4UZT093YjOeBPLD2aCk/v5ADoHpw1r2UbWVgLwBWTzrtke+G/PKh54W4LG8EnxqEi
Oj2qnSgFaqnfmtP7zPCLp5ZhWFg7PxpNw9PcfkdjaFGJ7ahf8c9QVLfsNu6klXEMHH0e1qQRfuYA
NdcJ42hEfNb8PLw/wNZ9i7QaojFnF4bJicPMoF/ibYoEwnCM0cbfZGCE4hJSFuErb0KjBl8w1PiJ
PxOmdZsUyksk7a5jSPAb229QdZMnWpR0Rb7eaEJX4tVx6T4pAv3eJUaeB3MxY35VQkH5giYXNyY0
bNszgDKNwCuEvgbgVY6KsoeOxr7JSrmTdSmyj1LSqElFIwpnspLRiZ5itDwsJLUJf9WJasBXM2KV
BNBuOuBRplDGY4fH1E8yhWv8kRHyG8/vHGOr8SDoNURqODGVqLveVZIyDxu3gOk3Bvey83ENxVzj
Z2NwXLqmIlHXD9JnNJILtZZ7oYcCy90VCORRU9UeeZp8tfs9z5KjXo72BM7+tMwQb+DrUZeI+YTP
3kbhThWPcAVuqP4KR7xcj8WOF0EdQFg9rdDawesebjWCwKsmsR1o/Ww3q8rM4JUdekFdv3FERJNK
w0lWFHPcpUtSMW/LAJ2KAqDndoNBCRk+xvAtuYWLwDCcIKSdjO0zWHZUIr7+jF1e583RGk8lrlJ+
Ed0iFgm8N+G9QU2XfxpPsujm5AoG2TV6gJlBm6FGlx1Zl8ioZ5Y9dYtxBglfUcCu0NJqdOyatnUk
pHQ9oCfKG/jJnbs7PqoqEpg9kgvVVLUStpHThgGGxjT6OtBZst33v9Lj7bC6G1MuJUSdoKzKw0PH
gmNO6nb4ItbEkr26/J5cCWdN2+ZdDrR2xdFsRbFkuiVi/YeCRnr6lud9iFO8DNUfcucU3miLI0YG
PlR1di6alBr2x+QLmabGym5fJ782u10dIdFEAzm4nXAoe4kK1bGAyTznPqMHp81iu2J0SlOFQZy7
3a/6U3jptTMlmkpWFZ64TcAAba6sJkdiU9T6PQC46x2MgnIVwHDwI/wDKfC/d7BfwYKK2Z+suQj1
qdGryG2QJ6frakZ+vWdpnwZ0ydndk0SouVApPUoyUqmF0Y8pCYKJrgz21qx20sdmaHUYtZGhgxKH
S+8QoLRvChJfGoVKsHcZiDJ15/C4wbNKV/dq0tODZ/P7notBXjTuNsUtQn6rueNYx5m3VmFi1fW5
JwObNJVvmgSZdNsGsSXxSYgdpkVNlp4FhLKxj+7BBXIk3xZmJb7jaBO8wsSGVg/4/ZIv5HLeymYE
zJu0PNsf89WqX/3Jci0+XzG7vI2rkblDM71hvar0ax3x8Zo9Nm9mlfZD/5QSw1oX39b6wzcPeqFk
uhwSZFO1vSUcH08CA0H9cn2Ztd7u9Gfwa4huzkAM9CHaQrXBPxhm/l54KEQ8kHbpkHu4f41gGh0a
Ltaf7WchZzoURkx9o8L7Iv7grJaooWaJhoTGHRsBIcOb/utyM8wYvdlYfWKj6+a8LAJFTtf1w+WT
xF4Ojr3pSWRIGIkBmVRYHTfeBwkZYDRH/bgc4HL89NzEgvlOTz1yAyy27hly1e3BqW+lhZa8q7AI
r1SfL+gsnNOREYVeb0puGxnpUbId1wO1WUBeOxIottUjb+8cFk343WJ0X7Ln+wv0x1kYpm1+W72z
lrx5c5SyXM23ejMEgbCl/5MYbW2FXv7Rxfvx4VaxxCDObsFK8mHFKlrj+bjqGQ2t32DritZVdaMr
RiwHrOIHT2tHwwLlWUCT2pBeAOj+3MkEt+spsXZdlKW3w791E+BnYNL/cGp7WfOvbU7YkWYtbSmO
N4PZDO2w0YZCZn/Qvw51E7DCq/VT8UpCUwPjwjMp4/atbfzAUaUxlFEByHMTB/2ZtwZNbPX4ZMaN
PrbTBDwRF3ua0ms4QyPUuOXxsQ1KdYlurOXVIhFoNXH9COwUZTgRtp+SQ4SLW7h3b5xs+6RtCymZ
kK46waDw7nVsc5ppVGCodnjj42eclqsQoIR2HWNOfZUuTj1VTB0nswhhf9gCGmIk46kXrk/s019M
1H1fTXz46L83hww7LuX0K/AVfQ+JC/K0Qcs/rK0M1LsTWe8Dx7oM1LM0nQZsKjIF7AE7jf0jFuzp
hLPa2kTEr6r6R5iMTUhJvZRB9HCJrCfT5X1/Q8oeUyma/yUfrYUezZ0RROoLZxcYI1mWtGeTQoNR
BGeaeYkf/DQ8/nlA+Uiyzl1Vz8dU2Fa+KrMxnPIAiSfMheRqCv8NJ7sp+wK33fkahVSXmZcQZHVE
BjPHMYovxRJJqt+wE4wuZk6751guGEZWrt5287iuq7v8g/iubwLpKj0xnr5Gr3w/B0ysiOBT8Y9+
OcH2oFgh7JVHrkdglC4su6Xe+2S9r1WJRlLXIsEcsgFowBPHaimhBCQ1ZlujrWTO4Z072i718CSH
WdytKSAuAWigzyNrwPmskvameLEieSCslEKtgqHbMs5WbFPIK2Z1i+0JVnVArw/g/Vz+d16KNOOB
nHSFFEkSejPblig2qgon6kgyt/gD70n+w/rg5sa3OXi0j5gCYbqP+H6bkjgUwEBMfEGYuZmIFC/I
JcY1jvCf3GR4Ic6Rr48xunirlrTdzZm2oyB8wpHO3iwcmgGv5ibvxLgGNs/sNOyxjG6uFLQnf5bO
Ti6lXHJW/BriqSUzqIdrMLzuLWlZP8RPAK34KCvMyxKV8yizJNf3s1J8O/Y3u6Ku7F65BZ69Je9k
lnPG1+/7Ia2qnC5YMiIPVRIP/aqCCZMBwhi407V/D+uB1+f85I5jF0i1nL+atoehcUTThhQxwMPS
MtgbJF0oeBBbbhm4Te63CYyFSw0zF0AwjdfshtpmqGTQEjmB378O5G1GHSJ6WkVwq9dI2AJl5E0l
eROSMNWNXVEfW2uFhbQn9xABHjFVQQulVjW+MlRN7hSp1JniywVKS+TSBjMkQCFGBp9GUMGsAjOh
A/729nKvfFbLVZ0iXnaXZ6jPA4AIC2Xfvmz0Z2q8TiRXwRI9RNnj3rSN3srsaQ8khL+NA2C6SV87
J8L0x5xQCyBOi4AkhxjXuTGon/WMeX9nYFoOZ/kZYfKPg43U66Yezmp1avNDld4HDDxUSf+qAJrn
0nAP5OnfDO7lAHXGqLN+7mizwR30/w84+HCFGatXzicVhAY+wBVE+Bj4wvUMOrE0im02/oDlwfUS
3vA6oO8fCjBzHvw4DZXXICif44N7w1XlTlWV6rN7/6oc3xYB8rEzilytxgN1F1DI56SqiBxz/kbr
W+MmGIqFtR2hV60PIeg8rBWMKNjoVBnImyS7EZY+IA7yGaQ9eqJhcPKp6bKTP/2m6d1k3a8Z+hPJ
gVuNjTGWn05PlY1b/vAtdE9k1Pq0veQCx4hqnIZUxbfI1Bf+5bx0Qv0jgfIdAwI0tg4AUsFfN2uL
HhqacDv0Hl6LLziLY1i/2t+gVS1+G+yZZG+hTfTwWgTJqPewNFzSRXCsjgG+mr4cFY3qG1OW2bJp
s5ktaaz0n4J/ypyq6+LOtlHCFbLjyEvhSQUO84wDXw5zGDLKbcZNIoxbLPibiwbNRQ6QVT+r4eQ7
F5itC2X3hploBthmOa2WHj8xXXA/x5O8ysWx4Mq8CMx82c7AIp2U+ZpWWOn/wZnztsPp6X6fMlNH
Zqq1eizVtzoj3b5oyccZzhnn0RGO7QtIP6wMcUCNH0Q8VY58CpPqHYBSEPzipmeyQm9ImN0ETRF7
twvYZIqKLu3BDgsWFntPdZeKGKu5u4sg8XQXBK9re2tYnxuAhO2CmG5Bm3iRmGmZuGTPhVGraKjQ
Os1bw3B6tbAM+yjQdNHhoF7FeGd27gUXF0vl0KJeJ6Iz5xJjrDBqqLywwrr4hyGFs+vf3mWndUjt
ErW5SiYzyZAhPiKDULasZnW4ryCYHKLaxlmKtgj6qx1jEEsiC/KcyrU0COvzJDwKYQisxR9g3AX8
S8izAX0KFyYFKMBKdiP3vBTz4eTzp8bM1L1oXHvIQlHvomxg6KT4f+UIpDuU00DYAcYapsg5CWAf
wb+bsrTOuP+dqiWRmvYAJ36znV7gM6SD/nxgQRM73AIi5qJ9qqOI++v2Lbgd7hvLKmZ5samPqK3L
DqJZLX5Yw8pnUD1Fau9G66ylL999N0Hmks1EW/9HRt/u6rOyBJwpW0GpyO1kYjMkwl7KQmlX8qXL
qIlr+/CGXK47D7y66NWr28RvCEgeOo37cm1cXjnx7bpMKfZFImb50JF51+bufCrEMxXiU9mrpmIH
QhURAXkt+EL3+cVl8gCnRw3BicAIwuzjEKro9E5MbMEYTobN66Ja5QnnYDK0I2P12/4MQi5dKDWI
BTHa5vjJtctU8m1iYynhscd9uLoZo+BB+lkbMBe53bckogmFsDrkxAfXBlzsAyc98fxqSE7Bzf+1
xM4hpAGtOQlfERJBixctMXWFTXCzOKzsyX0yEul8xPwbdqfdTaggCGZau5a/0jbCLewD3EqjTpCo
I4l73FAWiO7p8rffyP8T/ckj0EqWU9gaqnCvXIAF6tDer8Kr4VRwTHSiVznWp54471Y9/iDDDLvk
P0sZuWf7PxTQs66/0HGcXCoUwshQ3x3TujvMPTQEJ3oC9y4RCBntvbJDXkJNSAWkU+uhiZcZHZ70
Zt4gUU9g5d+V9y/PsyIqPSOk2qd+uEKNxliu5xkeWxA6Zxof968HMNGOJI7U1NZXo8UewMVff4EG
/TRK1UTv10fK/be8sLW+hNiuQyZJlRZ0mNwZxwWtvhwozjfdHnMGWyTwkrRpezraNpJ42+GYUaWA
wVV2S80HZA+K9Dfj0X1NO1kGLncvqFpE+rspHEQipdg3diOAoPKFU3/m/3SaYz0A5ppvOm322iZk
Igf7B93E4Xs4Npkffq/+OsC3HERZoR7kRd4ukJsQyKgvdx2SOQr4mpF5mR4teqmA9xH7EY7yjuuc
1wY43i2iCEMK7gxeB4gLVrZ8TiF7Wtsxo5+jraNIHGbe/izbu7tE4uDeBZdvxlOF3mmbEWUI+QRY
UcB1stLx0/SQ8HFhrSaIGVzovmGM5hSuGNmaQBuj7xkMqae+IkprpbCuNPqPkRZKT40fU2wV6KL3
sTaM8KAkbqobZfS0y+NcqdhI2ZEOwhQz9SPPp5yESDZKZA5k9XMjuP86ciO5Pcmn7xAknNHiTaEj
GqNsnfctZkE1ujels4bLlYfldUT9mTEtTqCgdjoOZUgTXvpzbZfoa308MkrQHbxagmJI23gtH0JM
1CPCxa+kPgARblmrap9urAZnHR4blmQYLFdRPd9nDkG7Ony+zDBxoAGbpmVmG5erV9C8wn2wfR3p
GQ4Il4t2mNDmp4lqFGkMUfSs26NFP6azm7U1QjQSaC+bYFzj64oJrGEgJrPhjKwvxPixEvBsrM1B
rJWz1qf7yEjdgEehBA6j0qO6+M3ff9m2X22Bs+7zqwPyJqNn3LlVz1qtauTfhCMUS2P7HTq/JbsQ
88wVMgLghxcYCNed8+tuWZNDo3yRAymHJJQu+/I3D2GCD8LWYHLwlIEzQGGmkZLo42RJQONOl+k0
EGubVXnKBbvlfSXlFxRdED4auwd7X94OocuN+nTSjEzFNknk5KdesL47/c8zw6TE1KOcFBo4/sxP
toZobr2tLJCeSu9ghVUEshBFocI4waDl3RGHVvu5JxrlIlN1x7IW+9mBGm2G/HwO4vUCAxFKfaJa
z+ISZE7+IfBiFTLadmb8Xe8egfPm0FQd1Nm0e+dX2n/fzWWFhlpieKqLZLF7Hys69ojXZPi5qJX/
8npZprgfj5LyhJbMuMP8DjuTXDU7+a5o50JMEfdUgfYArLIc6cxs/M00ilsPNZKSJ7mGaQ9R5jjH
Q2nGwWUjYyWq0q7D0/ZpTCMNPRNRWHrLSVFxG3pgJpkcxfjSY0hHneCiDEIJjxbbtu57pTbdWLMu
mIx/JlP/+OpH79P2NNI5mONGc9BY/K+3uSrcI61kAbJE2e3JMw1WWXMl2yDsXG72j3AZpAwEzoAv
VPTjdV7brd940tb3dPvSIh9C75cYixL+VPhgPwCA8m/rbyzRBug4NqftY+Lzq1lzzSN5kFKQrik0
pcQ+PaRe7W5j/tPS5AZ+4zi2fabtTINwREyKjPRMEiEQyKJq9OfkX/9lRnhE1MJDLmfR8HxqbJGF
w5Jy1gWv8gYJxxZn+OpaLn2rACwq0+9gT1EipzdAT0b0yFGbP44SmYH5s1lw1ahpVevSQFeKCo2A
3t+kvyx2N8mDLdxH1KhZrQFYqUDidD9ZYHla9tnzfEQQGl8FC9f2WlhCHn0RmN43KdJR+uWDRwl7
OtoZHh1JUGC+mS+UF7BxkVNX2peDVr1LWYV2QqbsvVoOQCmXQsAxRrf6LXk3sJo97Zk8zq00NeKT
4ZQAtM4WB+25uIg+eYDnveO06VvGoQPldXd+QUNmIxPe7+BVpIr36nOEe7on0+txCi4ssoO2VVf8
1FRtWEQFeYgAbQqQ3E9QIKLKn5GivwVNaP3S+AuE4+AQIVblryzSAxoaJiA4mw5JKVMbD82Z5hhG
csziMcpllxqff8y4hYB6I+WeYNxxvLzR/V8KxxwskFMNbkS0EMDl5fdAP9BVUtJSVps+wxPnYjAm
QZDJhyySySl4Y+feFcEYXap9FfQo5pthrP6A0BTKeeKWspl2a5zLov6HP5/iwePZ3Wu4Fr69JOWz
NZYV2tAD5Yn5YJN4KzH0yUiYBOImU6aGv9hZPPy2KrTNnKmCTOsQ8ZEp8otESli7RYdwBm3+OlxJ
MceK3BD50jvRCGrzX8tAjvh58EdVNUCooKbstMefaS2IcZYVGUSzRbJFlP4yVs+7F0iudA7WHD0P
G/oUImm12lz4Ag8TOqgT/hyxdrcOEqdvH5Vv5j2pNrr86K5lwXRIbeuA1DTHP82H9OLo8PJ9EW3G
d5tVbeDUCUlPDLPZoaUIuepzE9BbgXYx9DAcHCQ6Zbxk8MAHUPn9SVbfIqK7oxfVksLxjSbNkmj+
ix5Ekj9fYl9norONvie01MXzf+nCfF6NWs+/WGO3EnFynCLQHCY/b/oomR6NKbGe4qs7mFPj4gN9
sZgvRjowhxPupRKr2SFpRk2x2yT67hSUDUHDPVlWFfwgGBafRqzCED/mAsxq9izCRd2SRB4dCz/U
Zm07fNu9i+C79hl4gy2plKy9dU4zqEjiwEV7slo61KkasNDC9exb6745j8ZMTDKoKoRVZCE+bBqp
MnSL9JsRZzZzRkJUSPumyTfFFWP9E/MW09RRF+fyrZjUlQGzygUztiHFlc00cKQ5dzGGPX19fnW8
IuGz1AdORSLczr2Yu2JX+uJbK8DiD9OA98nEy2GXDCvrnf1c0KiegNVeS0Q0NYesbGJwIyAPbqzu
7DA2P6HPWAyLGUz2gcULcRDNSLaqT8EIABf0fR8LuqaZG7r7/BYOiyyo+/StAq/KWNVHq0Xu4hYh
NTKvj9RyCbbHixsIN1+jV7dEQAlblzQrerYmE3XiY+Ezxah463n1DbCHAcjYqvi9ZR9bPqT8Ybip
/rVSwu0ttWc4gpw60P7oAI0zosdetmGS6Xvn5vB7V6h2eth3/7mk/B86YLwVbQF4vzGk2F6ypyvi
8PHTILDanGVwuiv6lhz9dwgoZW1L1V3Q5ZjvgtDdVikolImF1BpN7GQB1C0a++1vrgPMHDxdJfyZ
Gj5IDXRiriEUaro3zANTcOaSWBMKaYjNZnpAfTGYdhVFx0l7C9ZFlpIqg93rlCMo6jyrCPsIfTAh
W27xWzfB8L1ajHxp04pWm09QzMr86dxaKzBLgxqb+Kl++p+Ei4mBT9wh3A+3yvIMx/Sb1LO6E1Ot
KRxnxoyFD5y60XwjE4Qjnm4k3Dn59T3q2SCWXJvVHpjRaZ9q9VrnIS8GZfpXlS/5W9aXM8smqGdS
EnyumBuB70zLYepUdMdD8PDVigK9+/jGWLRsLPXgXuXZNM2kLqH1jQmOKeiVW2lznglraVvqMdTd
M+wuMOEswO6eB4gQhMh0BXjXPVuFxOp5Q3KcZfg8Ijijkh1m6I2iIuMVV2YNu9ZS8+77uEzeint+
BlFUF4IDNxlTkycRTuoDco8PIf8CKTmvNO9pS23H6uS9z/kc1wlCJvQ9Y5yXWDboJHJ0n1DtJSqq
heGPybKAm8/zDGN+/iUxCLc5XMGUwfKeHqgyEsV3a9vJ/DN37RYMn9J9INYzv+rnl9jFAXjKNaaf
J9GdPlQB3iDEEIfDoMhKmDBih068QeaTkdZ2EyIUIFG9cCCyn1+uWGR49gzCT5gpOCs+iXIHwMc0
RYRoX+ibIu+2fbTjjQpNl8WjLXA8+M47sMleU0uU0Pfxt0bmJKmAxrMStZaKspzmewOhpZrJzTuq
pD8wzgWOFajoVxorLcDiQpsA/bOBMM1rLpyLMquLR4mUPmJDOc7tnZuRwgyU7qte3jKS0vapVkLs
SchD2d+qua4/bpyE3oEyfjpoHQFN2OVpXVAPIpkjNcIwUoR03Jud447cB5uwlfvXSd9XRMiJjN5A
CQnXLf94Qz1TUsP7TcBZuXn8CuHkvpEBFbMdhAMpIvL0HGRuxule1Ce2YEzREKUi6ILfOL6LgyDC
Kat0YtX2OVnC2jx/ZMSooxzJ7SWLqRS6UGaqi2/sgWDxy7HiyGtVwboxKtGNcKuNomWxX1Dle0WN
jmghcGyMaTdrFZRXkQbamMkpu4YrHgib6318AWF7BgMuSUxeuSJ2id14b8AOXxytaOxm1R4PdFiA
ZhOdEGSMOR7wplcLp9HQwa9i/rMUnK5xhFbVD6YnSFFvDU+Su0aRTY+kBm5A9E/ZcLT60idQL21O
APPG+bPRljjq7jE2e0uG3t0c7iKTFAFdLlLc1ErikdWue8SJA+qwG5FodURv0D//6NVs+PcReLLy
c75hGrJVI4rAy40YvaVoW+xzNpWsmNef/jNCarU6cZnd2GRuoGnXmANfLlbdI4leldw/Y4T5FIGE
qR4jKCyxMo92khXeDG9vgPAiox8hgeMp4D8XtM3hblk6R83G2Fm9P9NJxFE+iW2rhbf3DyaGv3AM
L1QCaorRYfYSpUaI21hFWhw3wMaZzOvXDni9NRhEk1VJQJi7C4PHE0nBIrYDc731A9mz6PwpktKw
5XMBP4xeaeazF18pt5MPQbDJtBfpsUT34QDQknXTuOz3OJbxfX7jXdDbpN41DZ8VL32JqpAZbfql
7NgfCYnzlg7li0T7lmjZBqu4uoFnZFCdYumpP6dUG8KnNfq50gRrWyfUaF1Srp/MBODgyr6Si6zv
sV0kyAzaziZyBTvMixP/kfcQzLkf9PdhsktgJE82/jxODK0qfZRp0qFP5i0pabCmhg9oRu9U+EJS
1Ilw5XSNCpAwRrLJK8dSHaBFU9ICFhhDJN1x1YxfOoJw4AeZovvwlzPVCEoqk4f4LUGRI6pruUBF
duPFa3xdmCIhyGf/UBRx7XsNxBZQjqBq9Xd+C0xh98kHQqiATL2JCze4qgxZl9KhScZbYhPhrLd+
wPkqtaZp32CvNTFUlQYqnxHwPYRGtjwoqwV6mKL1PccDVfWX0gSiL27INkU1IkKo2aFtUlHW/Dy0
JkHxLjHi7gQuKHfleqyQ2iNFtAOCcBKOKHFoN7Ql1xKi9NQRJvTylDpXTob+6uIaaqR0V6lwYgAN
XjkVQuPlBK+gQz/UbzWumg/W74cek3ml3MKEUnvKIysJmfusxe9N533QsvODQX0/xAhTztlp2cJQ
tIkKW7vscPhSFztfhkNbDQexoUERol377tH3q/xJJN7GkesLOQZgIVQrvr/yUncNVIZvQ2x1nRMR
lIQiPteZh5dSIfN9jsGbZP577Nley6MhNIWnvo8ARkNj0W108spwlBZXBbhqaGvdaRtd/f4EPuHV
YQjy1WwGXqk8v0h+8woAWjmgpHJMJOXQ/yGZlUvuj4CesXtjcqKWuV6IcJpetr4YkSXEFkCENiTn
O8FvgXy5HDf4jF+M9+CU0oB4Al0di+az+WVmqbWQXGE/ejHSJV6/2Jxy31PdPEJ2iptvr2ob3esm
KEOf8tEc8DZ7eGuB3qo/kVAWwotc3nBvxazeEC6xmmTvXIV7vmUxOrFmEQ5dmtQm9WQUBFtDYooD
Tf6bfF6sYnOqE4OQQK1yk77DIMRoL/kE9IzdzOHRC69Z62E3ti5X8nAKFff72Lr73qioesaRLDby
000fQil6AsWeJBZi6kK0Po7tJO/KbgMsd3yXddMYhanWIg/Eg5pzCGAKMMN1B433szD+szJVPGqa
LrjSpmNs7EGD9maUlU9Y5t38ehdP1TOG84b5sK8d1f4xlLp4SA1JbGdm34Yl8ibf7MBYTG4t73Vw
NG0N6GvI8/CCqBwrcJ+or17TKQYAsSJZmaV0nJDXFcwv1V6k5OGpCHH2jcTlmGVXgGcGpYoWPlan
EfBGv2pZqunWt58uGiM2ZH1T1eaCHQvBk8EDA8VhrnGngCexT7TQI8/x0EHYIUuTrWe586OB5fag
noB3KmABbhl3jgaUYGuodxeNzVfzuehHYpOoSAx5NUomH77vJUtpUKMKhwucbg68naPJqa4VsIVR
O48UL9R4Ej7sZ0txPqYbm9s70XwLN91kZppd9OOGOHZZin590HTFi+l9KaGssC1oX87+/U+yuVRo
+3eUSAFIR87oDKDuzVjDfPOl6WLcza7bduTS1S+2+dgPfQm6cvEYEEMyUG9lkQIAYQWryHPDTDl0
vQTmDrwawpNu0CHNcS4eoLjFMBNKveaeqEdsa7sYBMBczPiA4pU2SpCTFicTMPE5KM2Hd/dP9HDs
XWhyn5tmZIo/xYBD4YtZi/jnfN3Ldxb9YEIF0qHq+SqqndX09/5NGmEkBbbRl4+ASTVsyyJL9KCf
xi3MjC6OHTJ8BNQt/ISQyKTsS2NK3fGa9P+WU8Ob5r+fICpswIb66nqtRTuNnDSOD16+9urJUmYZ
ihp1A0R233hZVPAg7SpRgJrr50lg3Tva1CytC48vFQtAt+jcTqr/L0vW9XvPSjeRd5nTpM2qjVDS
TXrZimlAjsaL8JjvDT+oiA/S27Jk0dkbY5JpDDiLU2npobERYAJnJrBM5Nkul7ubelungfsMD9K5
j6VFKQtq4nntlE1N+azwj2ESb1/Gn9uMQMyZVKSWc2S0OcOZ3vvGkcOnIb3Cgh36kGNk/S+L/KAb
rp4i7r5SqwuySG2Wr261Un5KDqqGeZ/oPc/c4poWEZxh1lKyENpriCHDnMp9upIGeubZWYQz33uy
x+JSWCJD6cU1QsT6QtRdWjhWzgs0hakmg6KY+CJggIg=
`protect end_protected
