`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
Lf+T8jydgI6xLSeTe2I399+YtaICoQAOhr6TEonAPHdQhLbse+DsIQz9+5FiAxPFrx4ejRE7J8T/
FTtfDOTGI8x5aJAxMNnyXKBLWc0XWJ3x6mgzpgUfNEH+XxF/Z5W2USVGmxgSQgIeMq8k8KBAb6Le
nwmFNM3p0R8QqvS62Sp7gv5fDrzuZhC72ZbHoMayL5FowWDtIsWTij6qwLz2lE17oOyejdrxjese
tYCWmXLZS8LFO2fLt1i3V1QCe7oZM3iAmLfcJUWfW4BfJewHp7r7FY+S2JDPu8l8FUj4nUXf3hdS
aah83+Or8aFNneBVo8EiN52SzXSvDo4SYf8oFg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="sn4oF8A/bxlB4FJLcwtM9W2CwhudbfCHi1c9TbU7W7c="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12560)
`protect data_block
HPTslVVlkMldWsrm0mJm3vagJz3m9e1oi0BDecjh9o3FNGXldbdtPNC8KQwZkHme3p1zYZ1SrB5B
Mu1HAW7n6qNPfGsvKvOaInxCm0NNtlco74C8TFTQg8NhbDedpY4441p4tw2kwh/VtW3kwaQFotjL
IxNmx1QpmiBj/QqMXmViMAgSeJFKdrAecWYZoHZQ3WbsfVwjETpKCbgt3UoVQz4RtR/9Eq6HCUYP
piQFBQyj4Uw6K1CL4kxwX7atd9IFOvlegXpV2cpMw7yp55gKtOOgcbQYehTBfQL+Lss78hwm8URF
cXImGJMBHlYpjQt+axsMNXbGfqegpmVg6/367xu+VtVDOXhJHagMydd/HB+3UuuQR99Qa5erSNBO
WFWKxEkQaZ+XUCFi0Mb6gt9oYc/3PjlhqDJCExE4rMxSnRaqihwoAfMpFhMUt/IPrpc4thnsE9tY
UVCsAMDD+rWzpEZq0OmFEnifQs1FdPPrT7Am1CJacD8eYGJpgNQIfh5co1Jvvz+s1Xox0YmF9a1d
53RYgnCxGv3PV4WoIJq7EiGkSC05pT6Hl7fhjwuiEwyVidw/UMWHAo5Z0BHyvEijKOvGC8SyR+o1
DQNCTNP1IrdVbj+Z/dFTBmDVPY2B5/uTNzzkMQD3BlASuCN/ZI4p98f1MTds57CwkaLyHZkkQtzn
3sbk1fDFJViQSY4PkPTpJVG4Qlc9k6GlOknYF8yKF5RcLHAW9v3L4Hv7MbOMjsbsh+NP2WpfMByF
/l+Gp6C7nol25/n6mX2Y6p0wQ7vU3F9qZbhM/8VqqdW2dE+sFoElXeSm09grnZdnZPem6ATaahph
rOs6/1yMeqtV5qY5E4UDaeWGAiO0X8idtS2LairphvaEP9+pCRPlBZaeI2iNmxK/WuVab3Z3rdKE
16OjOUa65d71eQuVqnAaqpggLAPWPJ7fIXsFE7w3ueM1iiWIIFtk3etTVBJWAqYeFIv7kR81spvw
0lRRiUJUgEWqSawhpLhiaPfe0B/Bui+R9MwyURZg/DP4/6IMCGnFFkY0VuCrEqs4rcxFIoUqhnRq
YjjRQkxZeEE/G0GMNxg10bZ9AJqYLAsBuaQJIjOL7+KmdhvhAX6hmVjIcyAudYMR3cMRcntrn8xs
DrGZIxnoC5CAd/4BWHfEsDia2KM921iwptKbBPnm6UqeaM9IbBpWyMvAzFfqVHrAXY72mGV+AOtO
miozOdnFYoSqI1b7JtzQgMpu7hw1ARVBOmNOcsef1CCy9LtYIW3L4acbfX00nOffHtGKqwaDLFjj
2w0Fub++OXiyDrCfNE99511jlH38s9xaiH/9zgsrX6H1v47oGTn4Yr3XXe6QvxCIkH5e+t0BXwSi
rJZYekRYREYOl+D2d3B6NgByMVbatIjXN5TQbtXARaDUqYgomPPizdX2f/E8mnUDG0eDySUXRsQe
qUPULdwy8yAqzyf8E12VV4htIlXhbp8EJGbCib1GzZq1J8V0SpHv2wquabA2sEaQzJgxYaVpCV4q
Bcm+WZN9szPAns8KRT8a3CYZmzEIJbikT5Z0Q3gqFplpecid/xA2EgRZ7wCSFKZ2I826X31gJOge
PM6Yrmw2uuE1sH1Y3dkh3W2j7DgvpSxLsQOoEqLwJ1XjJGr9PyVJW+K69PLqg537icoLQgQBe7MC
ehwHUozTRtvLyp0yr9QNbSA3aL90kRWdQ3bqWaP3FC83KfWny5XT+gAVpRsnhrIi4BH7ZhoHsx0Z
2l1LihHveMNSlY6zyB32rcDDEu+wtc5d9OXRuqQ7zN+we0ypNyCejkmJeiW9LWO59nGvLz3tQYHZ
kKDVLlA/A/qEMIvv7uMV8zeFmxMmp8egdf+yUrtF4T8feH/un2iCVHpfMtnGSb1XxLW1LLDJ5Qx+
I/GaECOdf7KCMoEeGrQdV/k6jg4E4SloDg+O/fhOq/x43r8tkL+hM445nnQifoDZZUz2g8JzZ2Dj
ahtL5eXetHOyByRHLxAFwk3v0XjcKnb6QNVcMvPEF8/U6ksbRF4/UBy+19pD+IfsJ4NzsuQ2kSiD
70U5QURPQcxCfiFPp60W0C8r2kBJlr+zraiWt939CCC/e5XNJ7s52cBcdTd/1Ye2RP/xoXFS4ZXN
Rt+FTdgksvhCiCjKqxwC4ZsQYO/AhcbL4d55mtRweQsHAATVt9vUPEMtRFnReQBrmpOT7ePSRVhU
Jf71/0Axd2397Evb2CZWOjJoKbtMisdhh2lyMMnjCdpIwdIbcGAORH3ewxUCL+sK/g/bybypchko
at1i9/fqdy+fdF5cuYXbyfEwtMOyRPMhpuRE/Gik12IGDcoN5COx4iUbC4KoJcqJZyhnquO5h5uX
AYXgg/i5Ei9BM7Cpnkgr+eH3V0D00tdqCr6ZedKy+J0VfVquMVlWYf9L+TuYBmYNDFmihtRd0qIO
MieCHmOk/i02njJI3jnrEuMzLPnv/cQOQRP5t+v9uW49FPDdXVA/q4mqOAT8h0HUMV1tvCRIPXqV
Q+4X2uQmWSJn5qOOKP2CdWSPt9Pdxq5cbatF2kaBptTUYY326HPkLaAPTiHBMYbyTMs+t7snMltD
TOJChsYY9woxus8YgT/el6fWxoBlf9uHdF9Foao9USg3sht/nPaBa8ij9dWkwQVcwrGv+400qdv1
N5eExkTBioNy3NGW5mTyPZuQWxAM0Yj4jJB8nINSCezmhOUDaQEuDAhWDcgVruG15S4uJqt3u0Mo
9sQr77DcJmx3a4XBL+QF7RlagOWBxk/YbVJU6U0/SBt/QUqQKy73MGnrep7w7q5eAqJpNyFejzyY
fX0QWGUwJ6zhzG6/4zB0nRAfCvVQsLibYtw1I3p5GKFfr/X69fmP3XTh78nIt3cPZ/6vCJXfV8wA
G6PiciphCylVnouZg4oqOFjXQH2Ycuyt4hzabOzU3PXAQUUQ2HM9xtASGTM/HmX77I8P+QOEv5dg
E0PNlKq+Z4ShRwPw++13mEWfkKRF4apwMN1eDA9NF265zdBcnBGnaB+kNceyR5kf/UoYGrEBxKoN
lsB9vWjKmSdqoXPaw4XievGRw764o2blAQFwkhuEhjBavDqyHgigArlkAjDk2Y+RcmtnEcDaLMzN
PQvrIhBKr2eQkg6b03rSSJOGOvagV9x9LJuzBYbnROKYvbpgVzS86v5zAZVYPYCl4fTZMWflAZ0C
hwLMG9e6uPTo/RntDzj/QWMKEaGCKxgLlxRhd5Im6OnWU9Sc5nshjU6jFvzOQo+cZc1vJZaT7GMm
e9EwGtcghBEFmtDeDHWENKfV4exmhnOl6dCHaW/zcp3oVFR/M4bKVYfjdo1Y/YB8HWfsmbOW39Yg
NPMdrG72odUuN0OuH68or7HX7FMsIBr6aBGIW0WKJPCyE4vBTWyXKHxA101bfhoASzx8FeFsnol/
lgLJzx3gdZAN158hyrFwA91B8MYbYhHo2VQSJU81Z1EyUovsGyD53a37w6bQ1Lt+NgG4XE8B3nEo
HB9/eEZ5Anfl/n2lNreeA3fzeYnPQjLaQ5X7OoNTAKAGdWENEA6KwaJjaSRBzPt7f23MyiNnHkuR
sS0ZqzRolsDMcbi8V7MnSRJgrJgOnhsAPEfgUHjvmZDAD6YGWeuYB0ICilpuWt2Jf9wWAInAoLZc
MWMSDpUXhmwzMlLEHCSpsbslT243Ad5qsKNrKqxLC5V0rPeIy7St0ioGOf820ydlN8mSsElmOFo8
W7bAghzJwrYaDRWxcJb+DsUggJ0rjbsgWb0N/MabIm1JVWHmQU/2wjbI9AqLqV/mHHXF0PjtkokK
7ierE2Yqm2y+ivEqP8aDO6yifigaTvRDKODzeNuIpyFYg6spRoSTd8IxYK0QSeCdxo5MR/aopD5+
QTTIfxcv/6N1DF+qyC5a6SJK3rJXxKUhm1Ehh72QzzAKbiGDyL5dhVbaSjFSnQ7f7K+iLNGWSnTt
qLBRn0wjGnbAGu5tJXPCfH213yR4Vt6CFWfaYLK8Mu1pn/uN1wLZx1zHN8IvHlvdguK5B619ZwRS
VCyrFjq1TTadsKVjWrxSGPfULvFYlmQLDLwwk3d64r+qj26gETH9XDmwGXbbwnYSplHt4F2yEGor
k99T2CmZaT8m0I47cEmSsog0dL7PJqauB3g7lG0JTWRCH35VQKQbSpAApnVKw3PqrjbD6vfBbNs8
v1UWNXoVSRRT6yHtPi7FX+H6y8CHQJxGb66IlTRcA4laMKa3qK4AA0myxHWNJs0+8KS2J0e+s9g7
35QqCPytwAC1R0YqChu/laRj7WX2Qwerr3DlmcrQLWgA3IZGnjXdmgrKZkSyTSC4mhA8omYMym6F
MVZjc7Tx6w7p09pJr6RM7F5oNNzekW0wEooetxOVoWDzD7/8qXUmJEWFi1sI92o6QQXVoHV5oqtx
EuYRD+CpMUVdcyyVJZ40so7k/5ikX5d8aRn/MYZdAoBFCUdmnU5u7whgJw9x3QxfKAb3Q+tW+XSX
tGIMV74DSrvdZzjpHyVipc6BrPe43rCkfWEUwvN7abFp7bfRDh5/scAOoRejLJRaqGl6xojwLNms
mBI5UmqrIorGa3pbzjszQ4VzR2vFTYp/A2NEStOwCahExzKtsSxk+jlzPEIIa/s4zmZeuc6sEziv
WV0nI1Xe9jJPlA/axkKb/Towg7jqOGMxyoIV3Kb2mfYalKtMdyIrzHok77KGYv8LOSmIhLGcvUHY
/sg3pKhSrY6F2jCp06KzNWrxqQxe3ZRKizRBk5AyDruEP81wq1nXQAlplPeq959JvIeFCaFaYVuM
ilFshKupKHKpvV974MjqUyVrFwtZ66C43HjZ9K9NOtCOIcCIlkKSmnDovdnbvpxteMaHDwPwM0eO
ac4vVUYsgFMfWloEK1xd8CtCraexh5xS/JI808Am0InbPJjxXOyyc8DHKD6W51CpydrPRa6iiDzr
PPlTS9ugoUwkgQRknST6813am1fNEz7jjblmn2zdjVLN8D5qK609Hx/Gokf27HLrobP0d68Fbm9I
q9dAoyLNaqXt/ydKyiK7jvFoA45Xai25uVErhh/mCAjQTH9+hicENHikeYniR7oM8bOgIOoTePQe
0AGp8VccZM30azUwRV0Llu6PD9ohomrygj39WMWtQygNzLKtXiK4eSKclZo2hqjIzztc2E7sPbGC
mRcT7loovtnchPZZVjqISStCIeA9A+cGLNIFr+Xosdrh+0BJW/2uAYdZGRMTWplgIA7TXrwkEnsw
fpmD46gX62SEc6HcqwxVTFuu0DtDZ9Hjz3hAIJBPZaYWdGMiGN36bkiRUKnTMUcOYhFJmXbOLype
cTANaAYNya2LOW9xnxbH3k9M557k14YtSqk9GC6v/EHHus938fUt75rDnbTUkLVOSJtnhfkWCbQS
Lstw1qVfnVkM8XS1AK8Zrzi/Ysa+BcSTrBCLbNv99S3u1MwPkp6uRUjTg3dzeLcTZEPFGrGHZt2v
2ZPjU3Q1NCJcYLP0GklKm9S9He+sa70yjKoIzovCGu6Uy/ml/UwuupI1N0jkgFRYsP00GTmE2AZO
IgXxuIljdh/gbLkNvLm9vfn0jN5JB1B7w2iLic7CKRUDl7lShWux9eqZsnmvok0y+kfa6SEwAwJc
awwtC3U94vdvoXDBnU9YZ5eCdRWni8Hlhc74snTHyEOaXuj5oRZufnwf/1zrcVsUhLfT+8EpBk94
N4Yqhf4gtTwTTt1IF1vrhLBurpB94noQdsZm+gK8TT3o7uierOhBuSeN5aOoZP+srwSpbg1sse0z
4FsmcGG9XRxyeQSKfPn1kqhwQTNnTLQOXq0v+BT+K5AGVTzJfXetH7Uq9eUaJfxQMUDkNL48wfe+
wChTCStJcP4IwmYzIO9ccyORc5CGYWz7XdQF/xptDKILJYNwKyGZ6KjyfTZMc4GkJgEhDlmUm1bl
5DshYSDCJjPsyWsCAjSq6rsg8In2IlrQFO6gH3yPkeqXRbeO6bnf1ExobdaYp3rlxsOicYNSLilb
b8m3ExCmmPnTu5b45ZYBxQ2sX4rSpg71zqEG3YFFyC+L+gdabA3JaHtgIJ6swg4Lky6+IolgQAXO
7J2bUq7XKKEb+bn0OE38tQdAdhxzldRwq3UunSEHuE4vVFaUNbNKp2nNIDRFjigcMgz5Xgj2E5Uk
oBSAvDB1mgKZlL+SnGuA1IR+mK+oMTifQb+zM5KrcYnwMNsi3I+/2GNUJrgdLm5rESisHH4EuVCU
Q071Db1FAOKFPcgs+tmuGjfmDBT6uJ3IvRB/qa0Ml9DOsDndGexVp+ta34ED78Oo9dENiiypcey4
8qgHB7x2sU4l++P5FEjhGA0DyUbs3jhhNHTVk4ECuXuCdJkVZWLQRlW/mZOrVQtdQ2Oh0gnOGkhh
yTQuhB8TCn1zeO6jV1uRb0NrIIcJEusjNR8Tehqte3ho0P534bTmX5nHXPcMHzf3j8zH+6mAPmxh
8bxiZCxbjY8gR32EfTjhtDwY0ny6theowARYpZJ4CLJd3UhIYCADSktElnzO1m5xc7fdmN6vePtV
0cH3zuqi/VnnMAxpMAsiUYn7RWtYuqgBxx9w06ymv0F0DTSlWtemyaqPRGrzo7TpCRWzMirs4KIW
e47VpVzswIG6Mv1IuAPHfWHyoZWjI87+Kz4RYT7VozL00cgdojd1lg48L6ldtHeyIP9Mpz0UoNbh
Gm4G1Xb/Xv0BwMf8bSuXsdzqCP+EqPpzXK+2kFqsb0n+r7OSnuwRxz3d9mYKJzZoWUw+J5DF2/XA
DyEN00DCsTHKt322UV8aC7OtdAeAeVttHGhPuIfRL3DEUiOd0p3QJYzrqly7NqYqnWf4jRmAYYCl
tuwXcU2NK1ZQLjcdC8pU+/93n1Sh5w3dyaDdBWvNWHliLaQ1V7mEFCoAe8HhkADHXcq8UiZSOSJb
Slr0DY2ATOW/5Ly7WC124rwsodKNKpQH5nTutLWEcTy9voVyNSfVdXpVCRJyxCcxHu4zrAmdEWKI
GOAHoNwfeDz9r82x20MzWoF3UcEvwX9psv7ppYxk4yIiAnNJgEWQxFLSsChSu0aBT+atSxWGg5nI
uVzK1aWJ5OW7vENhwy1I3Xx4rgYeLR6GG3pBiqLOcl6gTi5ObpG0m/UeMqzg880RROCLVnbR9xuM
JctMVDizL7zCcWcDcwGx4QNNX6amVN4bs9aIAtsAiY5iwvKVNlj4kgGLgUvUvCeAzEu/SIfr3KWS
bM322j4QwUhf5/zMhMCLd9l5TEPcLsJtMj4DVreOGny7xHkJ+C4HFrKWXzPbgAN/mqckH4T/p1MH
yt2TAz1SZ51q34CLI28z9JNZX4416p0ZQLu+ZUMZAcA1At1E595BgtvYHuTj8F4+9jQ09JZrnjvs
QDKS0zAuc7dxYr8fYK/YszRxplncqwxk+ToyuXZaoIWNZ8pSCIXDNjthWYvqNB4bMNc/DE19YMHH
hToEZL3JHzeFT7G6sT260HUUX34e9NethBYifkrP8pOqgoJPiqdxPTUhD9TtgvHm0nvFtNeydX6x
0E3gOrH0bfsnqCMxwkO26YOmcmy+GYcetTJvrc5MizQx6A9iguobrIkbCu4MrxconadxYAeIeU7U
7TfwG2Q4RUX3hkxOLyob6VXKeRml8usyyrDPpoTk/eZsW8vjLJ2h1t+7A/+PXUwpWP5lMHkeFFU3
LDxWMObziT9SPEd//nrDLEVGYnLAueCiryS9z16reJWcuQap7dzcY7etyji4vZpyj57y8271iqba
FdmpVBtdvL5H8d9rQq6an6YpKGP7THZhyf5mueZCSDGJiA6mL1qpg1yeMdAClBu/CT1+rrFBFINg
iwapzsuKRbo+nuUvJVZ51X8f5VSeybX2ObcXrkULOb2fqFsx6OZq2DRZphPNJ7Bst5JaMCtDKRdJ
kvOU8hXsxD/EooKaRjEYruDiObWZIIsH1IdGplAjpSe6jAtHJx16716ssxMXXY20/Suj3DsmJEQo
uWUqUqXk9kMnRvoz4PD8nFXoaCFy3/tfcgQ1DsAKCk9C6wL3nXplKrv8fybtLzjcGDt1gUxpIQW1
64pofdvo1cLmLAqvyGh4OEAx+4Y/PdUmZyVso6qkwvJlMDvBO+7lb5HMX3tqYejR6t2uDdCifP90
YzIxzswl8ORBrP2WJcpHsf6XGTQnIzUYTIs8mPS76W/gQa/hDsWAIPZMklyYOuXSksbdxLHu+cFe
lYoHwVEF3Z0P/QejIm/3nDUiZaSZi/R0Oriz4Izp0RZEPaqtVgBjGDtS1IqQO+CeetA0jxpH9DP4
SxD2JM6PJNAGhXpItbRbDQdgnLZ65VCGJonVYGil0HGKorufh2KTmtJyvwTjy0cgy5BfaGJenDDr
siEnDJrff/jhE453EJpJPppJEOj2/crG2blu049KdyzmLxonZWJu5WayAKwy1VW0FzArEZA0JPlQ
rTGAdame4UDjLZmGUs0WiIEkZRwVcYPwjE2AJfjmcKjX2mnHFzffgMsUdsyoIRhiOqkUnXAazekV
0Zy5IhSNo4GvUQWRv16SmVRhIP2XwY0I19SOTicKvoPiWVQL9udHSZJpDMu/8AkWlMa8vxyiU4g5
OOkSCmJiXCe8JFIuJDVJhYggAJKQcmoAjtDUF95RvihazBXhDfTVQp0wIY7lhNKzNpmA8lH8YL32
6DeDKgEuPiLYg/s3h62f0LY/JpDKp380vDJHSmCBMGvBpiS2Zu/k2c9TetAvKvzcM7pyXJawvJoN
n5p84exKzZy47C8teX5j7ijA36E9LU4kjg7KJDwLOQBXz0aEAKJiQ9BnHg1SXeN05ZrZyPRToPY2
4zhBQiZwC8EG1kwwz0LYcNnwxiSQ6NqAdfrXAbSKHTJWkdzdJw22LAbGEFWZKMYfuJP8OZHxzG7t
AEiLdjFvYvflnIODrvKU0HlsChm5T9X9SKYaFVSPFW33juyoHFLEjejuEas4Fd1dLMsO7zk/86rB
0xu/qdw30TrzuRDG0vgNI6BsSIoV3Vnbgt8O/SzYlTCo7Tk7DVBcidtp2hjlCYJ+dYNWxpsH2CTF
EQZow+y7jGPG+xbheVbQBdaK5kmNP9cJPCudprUq9DQ0S6K2kvZrGQThjLAUuFuF70uEAfvdTph3
Hh8jByEgcLE573TUG5xyIXLgJV361D/iSAiinmXvT/JyW4fYP4vWXsG8ilef87gK3IGcEpXLfD0N
xcjfJw1+XVZdIQWBWHz4s+awr/DJigycnmaqLDXGKUrwHML626poH1eNVD3JgMfe1XMqrpfV1D2Q
ZRYhoSPjISk83x8EkMJvj8MaFQMIxKtxnKyxV+FwXndTTdk7Q859wDNhV4lPSZ0iq8RN98SQmmvJ
G7cUoLP13N4zs1lgPhtwYKZD5xTt4Dbg5HiNXk9GGId4nwQT7Mx68KjetS0zh1MOPIlpfLutyf+I
yQcaWl56oaKQ25xdqhVF/6wZC8iFSrLWJ5+Bwai2xB0jzcRSKUt9nr36jh7mLuQET0fIShV7M+AF
JgMoOXpPYtc2dkB0XNVxUE1FAvGpDIJwBqtjoaj9IHTP1m9CR3agexXqyjQA9yf+qmFsMiwrO9wp
J7H/oyYnBTpeooLZBevEOau6TTVdhWnMFHuvsiGQ9V5jWdTT8vJnHt59zKl9upMVucGB884596A/
dz6ZgprpfimPmuLZUeThFf5qybCvvcDo3TTDVZGjbsbX2N8MERnz5jbalXZwpja9AdUjby5tXSw0
LK4T5c/ZfXLbkF+WPUydHqDh4p6BMlIa0pX2i8WxGJbVfUiVcueib7ps7MuO+KXVnKPBypaO0Qlw
AnqieaEijJHl4QXj+QaDf4YrvN9xddoqBeplD3x84PU9Be8E4scJngPszYQ+0t4ztkkxEY90OY7T
gbcnBspr4WwCPuTimxj4+3WqspqvicWlbl5g2z+WN50R7qhNe5DPp4uMKOPc7fMicxGlk05r04oI
5woopqg39ZCs1O0Jah3UZr9FG9pPaIIh0lHn0IYyWEKCt0Q3nsa5+O4X2PqM9DAl+Z5Kaay/t2CB
z1f/T3QC8RbT5gF1AO2zVVrACXmOxkY+Pk6LJhVggqu2CBVKofQW0Frp9Rv4w54kooNEhHcu2vgP
ZAco17ACoTnAcqWbioFDFgc5r9l8mcEUKLgCR9zMLV3kpiC/ZGVJP5xjQsTL1fny17VqV/eo36iD
+2ZcwliGJAFTkLWyOBtaUcfgOMCLJ0NANZ7Ub/FdV/iHq2yaCTZltjk5Z+cspNPhvW6Xy+V81ZMt
1vx9ljllnzOKwR1YC7yKhfwhdxnAIL/74Eu5h/a41fmli7QZg5ehh2YAfHD5KTJQLz7Cw9w9qihq
6nfy8JzbWxjOy69FOgECW2jn4jjhNec6y52XPG22wi4VpRUfZVpUiO1UFLdyRuGwap/u3gJUK7MF
DFO+IAsEpsFPeMD0/NkPXIUmY5Jys1HtkZ/XOzLFWazpJ27aLhUwxuRKL1qw0br+AnLAV50k9JI1
Afp/75plUKx1uufOsky/vHP1aRnUlHQBUTQo4ja85WNdeZXgZiLe57PcfbBPtnGfomhgqSGCNhZy
dbNZaE0C758OORXvDHuBYPL23FW6OChbj+hFMsIslEP06I8wmwfUEvJjmKGGBTmFgdSSV0HLb0pO
YUaxKA/gD/xvJYJ+jvE7X6wENtjrcC2bNDJlqv7YuR14Cz6/ZJFWaTDCRvZJe/py4XgyumM0bhCS
oY+JGdc2Rk7hM9RPS4HjyYSqv69s1bmeFSqhlZdgXQuiB8Hq+DD/kuIOBIR9qYsGwzZSXndsJsGY
LARIlFJIWddJwGaowzbj78yMJcWsuFLFPD7LwG1hmye1nXsgHcaVxwck9U+fE8iPf1Agl+XOfb8w
BFLtmQF8E4aKeS4vv8hg8aP2bYqSru63tctShhgcGqzWNhlDeW6dUOzuWiJ7RYVhtf6tZ8atHCkZ
t3Ve1telZBS7muO+0QhvVNitsdFJrN6mkMpOWwRi3V5ik3TmTj8IL7ZHd9NZ2T2/FSoNwfw7U5pT
Qv6IJQR1t0a4/d/2ckdvygZpFTgiaGIuw0q/Es++9FPzceKRZWp//r5gjIe02fTZwmns9MObBvjy
DhD2nbloMF+wv2mJRyUWgvlqUW9HM7wX2Z7YFUK7vjhbBGOsNsA6YqOygHb5hsS/eJq0+YfF5wCa
BOQ+lHDZe1zIMxVdr90lOZqdlMfITQs8s46alaGQAUKgapvJi+TgJN0GIbsOErpKdZehkNHU+Nqa
9+Z+64YslwQtV4k4SH9WvYfBD/R3EjILDWaP10elxi8UfoNaTovNbB+Wkpc2iLTQOWTXxI2KeaHR
WwcqQqmTDDL/V34d9ujq4wzhYLQ+eShJnC7x2TBgwb/E9Yy+NuWoQM7PzQI95t4nY5P7qTX/a3G/
RfxRNfapkzjIXHiZPcHsoXCedhyZ5yZ3JmILuh8e6wH5KeSSe//pCZlGQSilZOyz5Dfg5FSSLg7w
BonpzQdG85UyIObrB/bCyprdMQFR8Ug4nYyifQZPNVUpy8TCSxp84rSe4/rPhZbg6KW3cT2bGRkS
izFQcEZHLSzfBeSIppqT5ZfCIb5hB9YL/TMoK+lkR/9aOToaBimCol+tlBRjIq/sZde7n6nV3iEg
prmLQfW8zACT17BClz0hS/3nq3lxtRcZK+xO121xaT2YMoKINlN0l0bNHV8CJaYseCAcGmB7Oj5v
Bu68Tj1ZgjOS642Y+AFF6zvqkLC24M6lfo2YQokqFNtbhQWwOyIde8jgcXrPauu4ywjH8cripfgB
uhV03k0dExWpj828wwmPbWgN5COmdtE5tW+2gkwTLilJ9+twFaV0fKHff5KwYJSPMpdRst13pgAp
G0nicUe6Ssd2NJoRuA3wObZHAfQug2DtvZ7MuGHFcmom5ivvaIH8HBTQ3MckMBoal+Pa6TvoLO2C
e5Vs3WPiC6i1VgBASGt+Z+Zl0cVFxNAcBdUjlAp5GexBVtLRBkVYDNsRVKHAKyziXI84tRikzbRe
wdfw3hzb/XgQoFVOYGRnINgqILWReTWEKM2aKi/L7ogyapdVvp8e0F97dHotzMvKIySKEcJGWU+z
DBJ6Eytxk7f6Hb5Z1paTAbXNxuQPk2OdQ6hid2pGtjaC3zDoAe1qXM7glVThfO0DQeMmme0Fnbk8
yZF49/Irbmb5bvUKG7uza94Y6KA3/ytkTt8ON6tLH1dX2WT1V/VHQHPL/Mpc9GqaqHwKzh3wcnUn
dq3m3/oKfeMSyPDCYEn9PCVCl22V/hUH10Gu3yk0wgEkUuVFEO+/7dBs8t6i5kQS0/Pdhic4xAn1
IJKtg/4Ii+OQhRyrO6Vb/5//Xe2Al2CkUmdAanIODIADzu7sxw70r5jvbu6z6A0gu5KyyPUGxIq3
7mL9RI+hYJBqMqaa+085IYavwaQ95BRvSyUqtdjoEZCPnZBI0INHvI/FO8m99oefufaRm6cI29ST
HlTg4n1X0+a+h7NWwjYr1NYHV1RAGyt2R+zRx9pabP2qvNWsB8nDcb99vX4fY4OxQEHMfkbcc0Vb
1vl3W8hv5Jqvjs3UV/k10dkLgvVshMdo+cFxu73WcAs/EHA9b1NZ1/TGB5xL393dhAt/ZTMpVWca
SzEr2OE9nZHx8tl4wtFmtxQ4q8ajou+3EzsaJvJi3J2lcGFxljftL1/drUnELDDgCkS6A5H/ivrY
QPWqe29VKqC9SAabJ+1T1NIlgf9IYJ5ZCU1BUueLPbh6XplFNGnvy52t7VNVm1CqUOddsGbL+OtR
NGSd3+bGn6jwR6t1dyQrIrm2Bn/NpldyNr3SUHvDu81qtKneb8qJPw1ARxLaCxlD89uvU0yIVypQ
/COJCeDeyhVdOI1M2hA4ahFPh7B/L4F1sMx52uzTI70nnxZtTN/l2AXy1C41otRw/Ys8/7/McM5r
4UR6V6F92HjAbfaPAXWQf0bnkfqFPktVjKiTBpD9sR1fc1B6B3Jz3N3JHuID2wwRH9rqJWqFK9xd
LHQFGevkH+UfeVAACrww760scrXWXozaOiBZ0108mMw5R9biyJJquW/ShwDibdkAhIZYhIimUfbg
2ofLFqrXixJTH44Zj9ZElFfp8EBLK6OXGlEBdL9VCCzphLJ8WYwCF7Ew7V2tTCpaPgDvpNrXLJZK
CeS0LLffEHPyWZoUQhZpOoazW4T7hEKGxq1+eS4K3xcszdNtirveKPn8PTruaANyMbDaIW2kTG+2
Q++vjyd6oPN7Hk9c+3ULya++kwQt5ewTYl5GLe36ZLmQAREEMCH4q1hKjzyk8KhYZJu598ghfTdC
Pja9BbD+VaEaF/uxRFwedmS+yz81SxI95xhZ2wcJOBy5YOuPKoivnWJ3yk1HpvlYzHl8HYoZ47pI
/aYO+diNIIp7pq/9KKg9eij3KYs4hyoQxF2CT1sy+1bSCRaxug7is7GxYg5N2h9LiRWkku9IFM6b
z/yTzfJVaJohCVrgoeQ29Ejc8pdgk5eVKRwFR9O/INZYrR0ukuVgYddumWNVE1zawT8I2GRDnAX1
JBvYDYDeaO9RedTduEmxfT+PLfnko7VTgAOkcoKmHf9k1kv7J0sCWa2RSktDfAAzrit24e9S6B4P
sefcXw8zPvArmgjYuC6YAvmt7sAubfKEzId9jXlke7mZSKZ3G4bdlTwrj87nRNlMzRK29r40jXWh
nmrt034tWGlHf3yar/FEj9mR2Pa31hYdAFkMrRW2flw5B98W4OW4PmfUzlqLCJqpm0vMoF64cGxS
X4BXEQxNEjbNExgyQ3Nexv6ky6NRqIIlfdKtMDWv6STqQKoMe+tvBqklkcVGE2L+QnDsMsrG2vgb
Hz4JKjMkt8HL/FZKwqt4ELJXb+apo/8bWaqgeI9FYbczBF4rLeQpzUcysNAmKMHJl0gJN13G8AK9
W3dML/F5GXdGh1MnlViTh44pMWK0gZc+mFYgXfV2cqz10XcRgUgUI2RQjrSuBdLcd10t0lfLJ+hn
F/Yf9CrxvbB688r1ZLpQbMydbmklll9xTA2gcG25OiF2N6wIptAJ0Lqfkj0zjzMxvkRXmOuR0HVA
eR/Pq/6X9v+pQt8xLQfK3l2sZJpMEJwmlTimFupbZD6/SQxxyJyWrD1tF+ZRjQe+5x48EvIescsd
aGkVJErIDnvWAZyD+J6QFT62lGr6Ily5ZKBp05/FLXz+7VFwen/0ABohWhbONDyhJkU/GeUADDtP
eBTMZBjQmFYETNp/EbfgZxdJfmVSK/sfmNQc/9wcHK3QfdbT0iMr49/jTXnqw0vlXoWHFwcl/T0N
8n2vAieJysJAyS3JlhKUn9Kjm4MqDH0xpoJHbUv9jGLD9FNM9z3hPzoRGsSesN1LYGLeDY1ezS65
YRfgLYH5Ogok98VX7HWgVqGbhR4gsPSIlHMgQ5gBYjoenk0eYlf4iyw+TVhLyByv5yNac+iMQj6q
LCUCKM5WPo7oK4IXZegqgLYjjmsjWdQRZSu4EMsxIcngWSFNIOBfx4pR06niWxT5mGDTHJZbKgyk
qB46cW56htMWPbLE0eLsck4KXg233kIkX043hhUqHBCbR0S2D0HdhCLRbGmY/jTQv5J/XrsgNak3
cYXoCfiJFRTkgoLwIarQAfe3LLFxqUDqQvWadwXpNCemUs7IBJN8iFaak4D1GEpFbLh9LKUALfKc
XunJIdJNtSVj9A1b5xaBZDcvUzeoNvPx6gYIFUaFxaaLww+nfY/dStOwNv3LC0pivE4KS43cr8tk
FGtTN5K7vCdf55hXU2ZJNJQoGoCUB0x1sgFhosIDvyOKjjZYP1cvAiAmwvwjxENQOFoyhmpqUvQT
+KIn86bNzGxypjpCvO+fG/7K/w3eUQYPVFr85VG6sWe4MilNHJNtXPSwtjI8KpjsRZxrg1mcBu50
wWbINmPtjIXpZZftirbK7o5w5JsUvFOZzASD4FJ3A4YORs058nXkGQe8Jlh3ukfzBP4VnKPtzqCR
/ULeYwmt/5bNvuB/6hLlCl6k0ZhlXH8m5BiQOODPFd618iN6gjgZmvAd3uwiW/kQjD8fDzcT3x2x
Do+xiE233H5KXL8ua+JXKWlBf7ow+ZAYXd6V5KEtSVgTN/lbfge2FCk+hVh+MfX/ag7lyMPhGs02
N+WGPnITGU3krqedeMnheoTH+0T1+f55Wdh9Iq4Hruwt0B3NQjyLROnrQKNARLsmF1GtQ6Kb8j0s
XMGLHjuX+vb/Wr2yFQnknBFgG1lUgmfA547gJeZmFjJS4ukBqN23a3otbYNN4AZ3Dbib+9fIoSFI
OdBlgc1LiecoVk18vybirkEVAa2So+TtNbHOF4z0rxUGmuHFZ+GOXLqh/HMtBVdmLLedC48mfPku
aU4/rJH5s7VjEueTxjuBbnyNldoskl18lrerXgLk3rGzvWFUY1E1mGygWOrtfoOEP63QiFXvFiFa
BtG27kDgE6LQ4H8xCEtU3gsM709/jHjqI/9Sm69vEl09IvHJPZAOQ0njYXvQwJawQOlqj8Bn7XjF
WrAC/F7ZcQ2LWR+0SHcIaZvaOVTU2jFstW8DwoVtew63ZX8H/t5xaJk6tQzdNS8EwWc3TkSC+//J
XzrzcbL/yonYigNdGGhbC3oYQCRsoD2Vx0lb3WHz91Y6/z2WGmRuEDhTID7n2Uz0inlAA1dVkkYF
pGp9GW4xCddbCZlmohtxf10kh/wfdR5/Kiii5LwBu0zbG7Q6eeAjrA64h4URVaDgua7gbXE9Hljr
dtEXPrsidAnBgvk58J9lX/TkAHi0l0kNAgKmTpqBFUbI+q39TCeh1ELl/IFJeHLvlmR/umvIH8Ht
yUpa51gETbeJmAsFhJZyF+Nx2m15r6SU6Erz28BsEKD59zYXy5a5KtSEQqEJMhlnXB4bUoG5CRQO
dDesCV946emWnoafMTB6frwl9FoaL0O1x7WCypYgPmF1VKaO6ewgQ73b3CbTVQcgqiy0M/35wAOj
i8JTuKaqrhgRJNo2jurTDgOJeILlMdPnrSdyQUEPpPCR6TYEhOIb1cgR1C+/CdS88c+I5BgQNC7/
5h2bL3OqN8NoQg6cUYlAF20yXnBjUodZ9X312nyGAUuWwL9b7cwxDChfATG1B1ndgNy3sBdRW5wo
o9e+one5kHbCMF8rJBtTu8DglX2aChYUMkBm37rwk1ysFwUmQDx5yaBlPci6vEryt7OPDhz1KtbC
UN+ZbIiZKyFRt2UUz+dXxwRJCAqbOQvA8idnlzH5CCIbHFj0sEz6JR06o2zM9Jzi8rCLOkCPSurU
qTrPpsFFrsRCW7LmEpbLFH3rNAx6/RvmWG5qzmSDR7I0sOlZZcnwT0emI4deoLbWIFbRrWnAmoZ/
z3c8kU296umjnlH2WmkcbmB9Tgrem3Pq0nfQeDpsn9boioJ+FYgqJJdNoYuHmH1uegAlSeBczgPh
V/qcoqRDZW2WTVH+IcAB6FgMkAEErXi7foxbZJdAIC4ILqt4KBNyJxSHx6UXywIdhqq1QfvdD6zx
oyb/Ye4sQlw/aWwVxkZF7TdDDsXi+4Dia54G0E4zLo5DJIVwsOqp0drwTGOhO55zPb013dSPNdwr
vSCXPVUD8HrJed7dQOhrp3u7suMkHz4WQVBIGz5LJ1efn0yMtPzyM9nGimRV0uv3LHsSn9FmuCjL
r79w7pRN2QczvkGIo8FLd2xwoMFzYhUzq/11+nIB5746s/Da2Tjan5TH78eX7CxtphlUkm89wVMT
UR6CopPngDN8fhi0pzAGwFtpK7k=
`protect end_protected
