`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25184)
`protect data_block
pQRHoUWIxqKuR7Oc/9BpPYMgkwlKpDqVYX/5vP/PjHS33L1i5DVavrPooU2u8fIfbIcM8+amzSaP
BuzoTlFi4t1BLOgklc6jwvdcD3prApGU11ag2mAfv4YTAvoUfMvT6WtDkHYXtsmRuhwi8Ht6cvsM
BAql1IpShaZJangaKuq9K78Z6tRhd+2tnTrqXIXaIWngPPkWs9y83saUvumoMgYFVA4sDfVNFdE8
dY1ZUs0vDkD/7DhIRA+xMqMFLZInDrIr6qDPy5b99x1q0qlHkuoPpPuDeXbKfewRhW05Xujq/0Ce
J9MoEUEh3UOpjFkkoLbDAkDyEf8x3QzNtD8ZpVD5Rn5SRwywpErMD6MU6tWinUx2V19k6WFBHz03
iMKVqzTeIhtcTlDJUuYwmzORfcmqCfh2g14E6CUO4BgMnU5FXp4O570sS7uJyUga2kOYUqBUOs1F
0XRrxaEstyOi53wQVd4+6W7BL9wCgwlpat+wVd1FIliY/AwyLCXj5jnBRSf/Yo/uFbql6IYwcsWw
fYVuHr+R6J/MQvXWMpT5TY78N2WpfPaG6dmEaDft93Lgy/pMEZ+TWYaXSIubtnpQK1fqqEKWQrrM
h+RNb7DCQy6gMD4ZQyfPJAnJjFdbVGyRf7qNf+E6ddVdXZlLGlkCcZs7un0C/2RVVg05dPMXsnrR
12Zs1psWWjA3jz0RILPR1jdkA9Gv9GLXd8ycN/3st8TjZNUFaCm7UaAT7H/yyx8k+/t3cfxHm02o
TlRQBK9Oq7sSv48pEUWjaX4jt8g/0PoiIBPE8tQKv+RpZVXwSUnHlTqj8AivhnxrRCOdlwPlNeAp
6AFKrzShQ4BlG/3Cnl4EnJYqz1PoRlAjgs3DZ9m0OGd9q/OT44CvvtNv+v2H4YBwVZslj+5KK1b7
BwJXhzJxgTHVV4ZIw1Qyktp1FnK5Mjaucl9X7U5ZTRYJkBNjSd20tVUp5R8cjZB7pvpdtQlgF9FI
SyE6/i2ROKknAl/gkxQv/TlPSD7z+vYpvynlOLDEGxYXyyD5JLVSdl+DHTjhDv3ETKCZfD+Zcyp9
0AcRC+w3xalp8t+WBJW7vn+2iZRSjs0wVy9pHAotyO8M+Hz8QFFj1iczzsvPaOzD0DTWh38CW90b
se2RJ2W1w240e86XSy8ft5OufXWvidN6XdLN/J/guSM9OjvTzYqkaEj5rJJq+r8zBSvxWyg8b2In
Sr0Dh2mTHVI8q5rGA+opKk1qq/bDpwTO2Itsyu0/55Hi36Su/Rcv0l+XIn8u0+d/xNNqoUNDC9Mb
WIi7+dRu9PUaRTsnPK03Y+vhKMgW9bwuB2sB0Y1BN/Od6SNbyBAcmtkGixmPfWn/U8iZp8gx/10K
P1cA6hPHP0W5ofMIKGXdL2Zoagh/hzNA4zm6o3AuSYPFR0DbqWjb4mnn91oiryL9vr6vs/WvbNQX
+jUVljQeT5t17a2f83/n/kwrbNackMO/CTJlP7cvlzA1+W4sLfdAOTBlNDFTDTSRYnunuDQxDOQ7
9OYUshP0Cv4EGUqAGdzMRgb5K9M6GUU5BQbNrVQNJF8MAJHc1Ka3ByzD4DC/j2TQpqOAq8wZMzvP
fMVLhuuETkmg+4p4FA8XIkenTPtp0XhdKisGA0kwz+IqhXE9+iepllDRSUGK56QJ7ssmelOca1wS
mpzcX6AItmokIQhIlN0Es/Do8SMZZJxw2RobNiy8x9k0CuFNxsXvANNe+LsQo8d8IIU0AFZ35jRv
ORrj0Wi+7nqSloAf4XdVSUAYvEi6q53juIHRIwjSaExD5ACWwjVQeIJqZiDp0XX7js6eXy9lV9bI
Hi4exFBdw09KRNbjLZxFzh0ztF7ZgdKFp5k96yOwqYtTJvsLeQHaDDBm615yXVgNI7GQkYlSlvdv
+whRyHqVmvcdS1Iz+tdOSCMw3MTJ7+IhDfK2qEoqsL19gfmHch+uBP1+PLAuEcx+a6/GN2q7bGip
MwCJBgM68/TGbfW8YbKVioQDzkElOTCrDHt/wNGAW4ioTJ5S4e6wFWwvM8HzUPq2bzGNSHxOXJC+
+72Zoth7BHurBNfYsm/ZMYct6P8Rum+g/BHdwER0Ywu39qTPc72KNOd0vQ4DUEROioyWSdKoJLeH
fB6JpX7L2CovVMAW4LW+EtBLyRutEl6j++rtPEh7HRHjULTMI8m19fbZ8Gu/sctV8mPe+hkNDt8g
iWREOnThobQJBCwgULvmOHYRDAtXsVPef/91q9IxRZpkDz5wmok8TKNsWBy5s5YQZfFq8+Iei4C7
RKrla3FwdxYVs2CF5/oYViF6se3WY8nEhKn8pqyk/67aE4xJ79W+O17cXDqGhOnfWz8CaGMfFqeT
hJ3C1QjDrJ9zwpohIUTb9JMpsn/VayxInYcVG+pKwGs85UpPCjAqN/qDxj43qrhYUjR3KoBRznjM
OFWxUHBAmwtnO3bNLAICceEIZ19CZanngZb0ziJK4e7SkC1ekX5tYAgk4yEkH5z8E+EOrr9uycho
k6DaRldqhPrPZw01Rqe7CLV7IV8E4OGFW0nXAx8Zg71LymkHd0tqkOHiZY9VEROeXk/s7EJTdj7Q
CuRfbPRqCGDZPRKp1mnC5cGxuEaj9bFiluCTVGDjvS1NvlCQy0Q6eH6UmKhGRkQLBvii9zgoPrTM
DjsR3Rk5SveD5zh/yDqhdOpRex+cil7xGnssTISGG+sTfxF0PXsiXeHax01stEmoP0OBNGP08Z+2
EUc78lyFeoic1YYLdWvO0uMy6KGq18wu7BJJ3WvB3XBPEE2aaSe3OvY5j5mIouxGdIN1nJavBv3Q
sBWT7GCoTRgZjZ8Dd+BsQC94R844YR49S2ORzLHXgQ21NV7FDRpcPFyBP2/3aZYxmnHNNwA6SlLq
iZV0Qj6vVasHKnNkZdi1Q/SXJb/xzB7Ak8XV+d9Jd6qN+x1vwKO3Vc0Y5TZiP+Cb2+fi5I6AuymT
xgeRaiV8uAMcKSoV0v2mfwE+jTLJ2mJqolA7o74txh8BYU8VbeTdgtQR1zU769a6/IO8uYurVkme
1sSUFx7wFUaixBXxwairJNRnpWgETPn9UpUTsUw8o97z/SN9YNJ2eozGEE+R97lFwsnXwUKsne7X
RtBNivdjrWkMATjteUQWrgaHy/C5iZnn+zSkz2F8BbTW6bedLYV1RDdzq4lKoDPQJ/EAP9s5M7Qo
A2RNoYCVlOlL9v6qvoClqQCNr6jfrk/LN8SBMUBl5/a0bzTSAXw0HjqqodXwcbRyfOAGtixCvFvl
TMxYSchohMnAiYdrqlWm4mhuJdKUTxJxrKoUza0sij5osROA137nOTHHn6PT1Ck1HcONMhhTD2Fw
mEQcl6Mt7ZhTG9Jt/HseN3C2hdwGQTWSz3RECDW3g6hpb50W4m1rm5ETpMpIS0N/wAcOWuV6j1zx
ckgBR1QiDSqPZulDwmoS18408JqBuGExXGbA6DDD5GBLUITihVbVsm/ZeQXMwDNTVcF5bYSVmDSN
GaiCWxlrcoZ1tCNPv22b3mkZOYGEtz6oNPJizFx0rdShqP5jkg8UhQI6pomBYapyFWIqvUmhh4Mf
Ws8xt/rslx8PHGUUJjjLgaEctlYGWF6vBDBhNCjEjFVpfvXO7K1fWA8AzMrNHNaxEbHDnk+aSaDe
98fHd2paJ2ZbXuzxPJjttIN54rbmdgxZ7OI6vU37PT0vbROHbR/c8xAaFTnFhmuL4f6lW73X6Mje
Ds03sCyTyV2JTgXtjUXOopIi8fsN228+RAW3s8B7yhVDu2hrumIOJWLqRjQV7JhiAcCAwymZl4bd
mcjWLCWbapm3K0sgOlWt6MKgSm45Ga7hJ0cjXeA1p5NejFHyiir2yBczDXPWSQp2ObS1qi81fhUw
e/P0AvJHpTqLHJB/F4BM3zM7yNxX9SG8iR0331JAvFD+Zk+Mq3Mg/xus1NYr3sxj17Pd/vdgq+f6
yL7Y8SIgrUopvVMpa5VAZn7WIvZAl/w8jWkYKiSDtuKtINV91AHb4m1SHf6nKIMlRpBBYjsR6L0D
EA0+M68snEtXXBsO2MULLA5Lm58Ene8IGQg5WQgEKICT1ukS1miJEbWjl/oHWZzTnuk1SPdzzwsn
XdlDUN9r/xpF6ZdQ7LHZLB/YMlEHcr+e6xOSnlgqDnv7BhSjy5+/Y5ZSkODjhZzTUzBKRf627mLc
lZFzskLRwfkHoEhkpuxyKf2PJWAD7qV7QUeWWMmXd/DbBrQax0R/1jeW6fBUSckNf1wPdh3bNO9F
Bto7TDnp3C63u42crL1CILYT4kt9dJMFGpBs9mzCnd44KeyfxHtO8jE4wXUkC18s+5lOXGOLSg7Z
6pck/9ZuTGJkjqwLLLx3KymMLPFgKN2N2LJLCusglqJqGAUOuJstZGhNow3jBUq6RbchE0h49aU9
FEYCpVqPiiEO227zN32mpw1TcQ7fSz+kdz+RAUJgmwRR+0tuooiWKhZt3V2vKd0Q+CshPJanuhUa
Ibw7supSB0CHLx4u5gCeHrFuXIf+deJcEc60oX3EEHVqF1hPVcTaar0G6x3VA9mLH1VsM60cG4fv
2iouJ7akW4ME8hg5OAwLChZfBVCU3p6BhXVcIBe0BBNsCcpw1+5H0Gv3r79GqSkrTntwhu68Q+ll
ZoSrctBryT+uiEDFhJ49HsEf+r24StIpU3WZHn+9VhLB7hnEh7LNbcfKfcTnoxzC+wHgvWIahJlK
6HuhEKXv2aE4wU5tZZOHyvWK87Tiwkx61cg56ixhAg2BwTlgAGCsOW2MQ2u6/1FcwwIVTkYn2wsG
1LxjK0uS1OGcaZaeiZjtuCElyYDPEZvhZXA/MqOrMmHa7SmI0SRzk7P+RPdG/9nMUGq4Ps/U3hYu
8ANl2bmUJiuaNh4XwVC+I+pTLd22FrWKMpOV3+OkfLk4twwVh6cUWSGwWy7M6XffiCgnw1cjl1RA
5izTeAQ2XEp6B1sR0FOx+yG/8lXzoBLJpt1T3XNc3MkkqNwk/TYeXFkRTO05MW0ySOLLVe/S4pHg
Hz4EWWpoAQ/K2ZSI6F7zoolwr+v9CIJ8fJtUjO4bPVFIepusYRLMDHNtiPhQ9mSfL+XOZKNN7JI4
dp+j4ehqUt84FO9GSOyX3sFTfuABYxHt1p3ytH12l92j+8L8wxsbeozw6mNo8SAFgbGDqfB1G9zD
qk4hzWgDAFtXmoGBLsAcmVu8tLKx7enmjH9wDZ+/0jR+pLoGyuxVKu5XtmX8U7o4HK9IKy9Jhxeh
Xwp/EipD9IzQkp77mTMRGNQHjoebz1t50XwhQEOLjL8ZnPC/NdWrrKkZyce4oqiLE7r1AltsD3/9
M8KebqU3WUARACzqo2/iLfAozWuJPdTtDMw/18DqsbAa8xfTP2F60ilGgYvDzDxmrS4M2ETOQuth
33MBI/LQSZGtiV7EtnAkUf/nso5+d6NXdDyLKBzFNtASgdG6/a3F/vT2tgfkNhjuuKNbdmDs/QVc
3fwPFDnKn3w7Jcc3FblmkOZHKTnoRkHQlQ/CBT+vNeeL46b1Y+Fae2XfJMLCtwXRJbOhy+Z/tU40
QuruVMdbSQlr/B5lPcBot2EH6z9cEWxrY11Vb27XSu6WGUot4HY5Jo0OGbxvrwGKtuct6ERhFGy7
xEkIp5+kI/eZ/jCDkifIt9pLXP1mSY7KHF1fKnGMtOxGTD063hMje4QTWu4NuA6FHPD3E/ubhxqq
IYxPb3s5uh0s+c/R4s++SZ7drw+uuz4n6fl6z5jplTkKiVhjVkQNCH84Yt2McziLfCpjclktt/M0
/z8rzzJ+8/XX6POXWmCvbQWnoyqNuCadg8f4bqKuAdE7W/seG25E/M4+aULDEVmxo2pQJC2Wm+qm
/qOKPzBmkJMWKnPf7sD93y2qmguy8mpV0oxOPP2UnZEOmXqpC4A9LUOJ9PwpufRK9kfjO0vZZ6ym
rmdBkASVEjQ8c9fjNtLgY3uwToz9FCsUHCBh/Tp82iU4onb9d/b1fs7BRVAICsKYwdYDZxDTC3N0
lC/d//Qc4rBbQH9oySsYopsJfxorE9AQqVS+lmM/hFa9GkBFB/4Q9UaWnYOddoVwX91BKrK+aQHG
WTIc7KTWjhCVO9c1zx4nzlHzhTOm3gf6CpNOmTGQY4TQcWC7qo3sv496vskKbzWBoNmdLlwQmNRt
6cBLCuvPGpES9YP8NfZVY77AT9VPpBqMMG0H8Dnrsf1nuVQxcOnvthsuVIjAac/q30j6SMDinsMr
36dXY5mL4pvBwaIQBk6Ydlu00ofrn69AykX7RsOzglESeLJVzMzWL4pdQLeZt7yAnoe88OIEhGQf
fiCmkX1LL3JNYuMSbMPempoeJ0rL4BvIJuACDEKtJ0PgUYuPbS/iYsjD6eFc5qGbuERFYauY7/zB
mbijXPBmY1LU9EyiOltFFIbTcz7gCT4wPAYdWIDztnZZl50Ogpk8xHmzEv7Dk1eXSzCmkURQtlhy
Mu4ajq5lPpb8MKRcaXbxu5NDpJ6Uf43QL11KczvZBb9FfE8iFDVkogxud/0Dfz9Bz+Yyclw4fKXc
2h1IHJp2BfDoKS8+DdgADlaAtKaUBYbCtUczShfNtrQWEM+dtVncub1VOm5GMFeQVrpBkO2xzEYu
bSNfAoc3FDiVr2/ZM4wqx1HgcRKq51U7UL2zlf/LWBsSooYXLLF+szsud6aabuNtrO662WOcYMgA
3cbPMW04BI2Is3MijAdmPgq7WxVP8XcLFJYiK1pSW+yisUg1zfB0U8r5Yr16DCZ0YPWEGXMMu7wd
LZWBZ8MQLRGu6bf1H4Rl8RHxM4TJ4BD31b0ImsKRuqnsFJBiBBqHjMX2bDsOCXWxc5XEmP9vSzno
wPgRWXR5tQ5+Ov6EVLj5wy0qmQdUSDmiPM6XpNHTy5diTQZrbZJ63yyjZek5+hn5kG5R0vF3i7Ke
Y/czSAtoaUvrzz5C7CAinTakF14NAEuLmKw3qaL0Xisdq2uzX6iCpGmCiERyzopGPVhqdJ0iholn
JBVmXFSzleKqf8OKOy9uZuTH9GOuxMvWlTyOTzPJPPUzOafWSAZXDvowMsXtCUokOLVvEERRUBLI
+YwhH9UmKFiv01D7de/3+Z2McQ3MXLeNaG8SRDybtsEEQB96N5mYkjyLbKLcoChsDjeE3P76ip1j
SjX6KfX9pGBqWs252V2OJAfNXsvmCsn1tu3d2Rgh0oL9/fLhRyv6DMlQLL/dvvVGxKrqXtssdG/Q
kbiKEQDXZ6/Nk3piBrofE8WedrHWxjOCVDfeoKc3uscNUVHP2w+7/RiO3Wjl3rN2eBRHWsseRZlO
y9P1F2wCe3acfegmzYzBTG5/ju8DVfEK5OwdtD9+zvnab/unHJSUCrISgCSx8BKTbkdXatqHs/2V
lhkrNPumW07RoI/u6LPOJK06nZHI4ZHY6ZCn8hlwxcH0GTbuO1FqSPYSClM203flbTLnqmioQXQR
SyUdbBkAcMbHcKj5//9jtCdf2cxMpTKelArY8Qx16WqFRJD5fYIj5I0aKzzxavx7em/bMh8q+nXf
GtwvBx8Ti5BMzwKKxNRWM4OjvEjgzDIvXSFUAGzuFYaBt66K86FYBfg+d6b2DC+vaP5VDMQbLKa1
uKAbbwpceNGiQPqivPdsinkanm1BtWbAXcgsQ9aenFdHeIxPc2d727F6qbhMYRRsxDvxI8n2cLwH
8zUGDjtwtXGtbpVE/PWq0hkUbFsW3wjuPmRddpArnvqVsz9e85vARf5F768ly2BSfKrKudvSVSv6
gEXdCthbx1Qvy+B4gnmC1pwzMArz63T2jWHJleQ5N91N08PU8z2/J7knPsxnI7+iJEoIBVSbUlLX
UYAXhQYxW1tUPBvHawHhtmsfd6BAyfarPuISYzy+AktT5rF6yhvJpX34fjW574AI3XLQSe0g8GsR
VXic9xadAkrTk1QEGqoJNbweDF3XBAAebkShPhQB2d/SoY9S4b6cFWOfpz9FYXT3dAq3ZWwbwAkZ
TFQ6OimqjwhsHP7+9C81CAxPytFEsqd+YHJdAdIy8IKNK6+UzSUkVhgvAfKFZFjOE0VQmwcnRewM
/RVNJhYXxEwTBN2NUPxCd17IEVyaGreix9AIMT8RfP5nyBeQ5ukCIV1D7nA3AXTuujbB6CqHTaGN
G4mP6NpK4KRFbnrfV7PdBGWQPvwHGVxORbZFywbxfSMKAhGKhjENH3MZUhuH1evaumH0yLXU0WwZ
VBOMo5MFbJsrWeGLE+TKZV7++DDFsmmAXf04NvNXGX4+V9rqbtz96+KksSbhYCztgoxBKLbdjLuR
e18P60tVdXzd5LyiY/1VQSVFbbn2tSVOZBTaHenyVCKTf/015Wy9zKTWCz5wdWk3kTJcQXmiKWgw
nAbpPYgiKCVRSH++yfe7FQ/sODA9hU+mTaud/Q1iSchqxfstBQWC7fOCfZl/zdvaB4zpFXgCXm/2
qznnYYAlhrnvXHoWiv9ODaDkAA9EmVthTNUzZq6SctfLyYbxHCgobz2YQbN3uM66Db7Bz4lJcfla
1rsYDoKIYPf7rkEMPFGIaMMOnUjEOcaQFN6dpfOPaiWSAPaw5XlvTmyhOd+LqnqDcailqJxQzo/m
RjpnR6+UmewcuY6GKkBCJaP9E4krmledDMapWxPUzvR3iqBKSnnVBstyz5uuCaSMRTKr8FYKSsZ5
pnrgAeBwkBSnAGHIjzI38koQ03Xuix1FkT8HWGi0TFzYfEpvHQAk8j0MzqXs4p3ButHb5PGeF1TZ
JPEjjd3aA404/WlsCzS7TB8Z6mwLRvlqQJa6cL1xGnbzsLWxxpBx+funydNmtKrh9KQXilVfgreB
c4ddjXHkynDWag57dM3LQUJS8y4pm2dBTBXQLESntb/4vZ6nsXnDwpUN8j5gKyKr334szIRvMT+T
R6K+9pzp+mL/nUlBtVRuB5BLJID0MFoTRkhY05CQsurhajHJhKUVZAoMcoQOhHgQ8wAB0xjTsaRK
cXIYt3ZTnxPTe6TZpFt6xsvBH1L4xACUlN8VAOpQY7rdJtXXrSTxR6m7LdrV+szR7DuNtO6jlr3N
wLlefdns37RbPtB8IRsnpXtSnnSvbQPzjeLhfVYitNgMorWq58OMmizf58qzf1Uy5bYsI+mSrBrb
nHoT6bPy7jKFU1+3qD/jp9oF+vyPCOR4pPLIFw2OOfX2OuM9nk/fyyGBVgvEGDNrV7zQmQlGTAqg
8iAn7QxabCEJuZQtJMLZjP9uv1wGEWuN5k4daYiqYv6KVkRf0H5iopN8RDTOL8gmlSyHQZTAzGfg
DJLNCxu2/NLdEub/CuNYH5P+E7a+jmoul4ucnH2nE896VU+kQaW/MlEpK3lhnWlQOZQ3I9D9fCbY
eEKl3yAF/BmgRL6t/hAlSsUk7ze2sM8YVM8fRUL8QzfFNJudLdqAd/I7+CBKOIkiQONl3xExrtDP
hN5NY35fWoIX7PqBb41tgsi2pQiDF9Qw7QjCD1d5vsinzCwWo6eA76rKlMC0tEcPbwbknylZZ6Ts
aDqpcHSSbwfHvwGEtlLkmyxFqauiJEyGk+1aADuuSjoJC5jRYE1BjpZMJ2XqDLB38M2hTbKmgTI3
W+CXuGqK5pFKzGa3x6Op66m4P4ivCuv8XmfiuVM0baCFWUxAjC2c1ArIycZkRl2LhBNX2/yAsRCU
LwJFXA9ogmuYS1eq/Y59VwPBDM+XENqC87JhoVMr4i9Ma3yoYlZxiz7XYB0/lmz4TTzNQRyTUZso
pT+qp4fSDLNBkgbYLsiyN3/q2R97ubJJ/ELrc4EHrgZBwdolesB3kAKuwjAXOsEvByhU6EqE48Sa
Oz9nGh7heKBAcj/+ALLjcehtMOLNPfCNAF1GSl9I7kzCg8281p0tMP0l17DaPdNM3qJJx/qmruYK
RePBfB3Vf0W4ZjaphJP6OKytBhfqFGsgwkaSeoMgB0PoHtYXallU7IKFKhSZ2w7L4DuOVvZmT79U
7Oa/zi+LcjxlhGsSYywQS09c+5A3oGYeVti8EN2K4hNhzOlGhMpU7CeTqCU7y5odRuNyrwiq8/RJ
nBkV7Ae75Gg/EPtclRpd2Ny16f/B7ZWa4XGlWw+4p+/giU05ArNyMGcD2goXS/vPMzu+jyP5vNtD
1Is0em5Ii9Fo2rMmTxUlZ+0nhD2oz3fIRw5uh+xFxhk0s9Xdz63mKUjVToUjP3wZC5FqE4Qcle/A
fh3WTdzIH0RyMgqjI+GWWd4WtHTZB7YFahBbVHYIuukTfwUOiSHherx9Z69Pg5VqldqtecHZdwrr
qszZEM1I6sAAbHyeZzBnsQCsVHJVInQ9Aph2Jo8CpZjxvWwC3YyKT4PWDH2Gq3GTBwdrF6JHBvOP
PW7XRcv5ixwQli9hsY5G6GJxrte1lzGtITQwrVKLbcr7/JixH1yxXShiSMU6QsPlT/EFS8ahox2K
zSd9+Sz2Z8RLdcCUD7juiB2huWakV8IoFKYS8wtfttPZ7WAFf7Fq/paOW6NEq5u7s0xzp/h9lBJM
fxNkU0yyI6386Opg5ML1nIZV8eU0I1SGplDeoS/z9upw0z4lnZcoP7mjQgaHv72fEY+BYYPqrG/C
euw2oLfWHNIJqPCr8Qx9MxCGO+NHGLJGu557hdG3+0pkcxLFTvLFYQGV9mMUt0i+2f9QGKa1yyrb
COjxax0ixm1zfDXndnDtKrnqqiX2GDeuRRrkaVL+2mS1QURwHy+exngx8E2F7/FIScjlSs8K3E2z
+eYGo2kzgsCHG/5PSgMG1itvqJku6nxmgSmxPHhSTBR8QB8Zl3UcQwNgV3J2rForkq/1A7g4r+c9
etcRMNCagxCG6DNuRdHFXfyzLRFyJSG3h98N+kBwPXEFwsmyFpwhcbbdAAOdWsOjA8zgjk+ikewp
ksXrM+P+pZYwQ2pMOSb3OQM4bIZr1cUQfDkdNyx12PbOSbuqmOxGwgKps6YP/Q5NBCcFb0RvIzSw
MTn60YBY4HvFHHuxUTltxJNaKFEyign6Qi+0MdhykgxkvKG7hnjcjJPJxe5n4M+QKKHuWF58d3rF
PbuL15bRFgnf26vNJD3aL5JvoKK7XowbIrmra47rOFIEECMXUaeujvx2Bo+H26Q68Sd3NQ1X5NQh
TbMRcCh6tzA8J+fNu99S08XluJMdFUZo0j7G7AON82Wz34HOLM9E9at2s1AKusH5FSJVGMQCLGTt
iEzNm6zORlQWQY+wF/Wy6V0NmVk1DlC1J2NGUazxSu5Hi/39cvWf/8KOzDKa+IE4h7VGhU7IGElT
6l0AIufQTR6dGu+TWyt5WJO0VAgT0J/GmHsXblH9gtrNyDeedOJpXR7aO2HnZgnipt0VNiObpyub
hXHU35RDZW7rmAyb3K10hW7Jwur4mbmZupz6MBQjgFYoOUyym41Z36v/gnLBdXQqWemGkXQN4Exi
hf9gU+W2z71MdFCsSoGQxTIZBrLmz+4nbb8sKYp8gBegM6gf95m/iHoDvKhTX4snwl98i7rjRJeD
/401jgoj+Cwg8x+fvnRVCMA3qGBpTlse6JhzuIiqGFe5Gf2mCjOh9S9hSzVgg/8Ej3HPdA+S+qMV
25I5pgM4qTp9CuU0/QZuKxHw0DSi/+BmYXlEwGxrpqZVaBUxpRTew/GuYDEyZCj4tsGl7iuSR3XU
5Ct8o03lfLhssj9LBqErqW5PEzscF8pKqyl1RzgDGBjul9kq19oLr2Vnm8opnZpsZSaEaTQs4o8C
cxkYQFWahDq7kuGjl/5RUpPRdFUwF7wEnhKsITpjn857HFxZSYUNxPO6kXF0AghQPoClfcJVawaa
sl+eEZuuoutbX6PYEvapT78vgqHdBx+pIs+gCFV/sg97RmWX3/02yTKlzm+k3GYJ9kfvvSYNz53f
/fGO3bUjoQ+3L92tA9AZw5xU5gGxtZDyOH6yV2yUmPKF2uvFUV8/hLOHTXXuuS2/Jhl6egCMCOsD
L6tioHIITshStIC+eNl0PLEhqsDR2IOdeh0JviflMLRVeNpLp3s7M61xw3m8vob7VpsJw0hP3MV1
GZgj0z0tjxqRYW/b5891Fpj2peBe3bnOgUYMB8Zx8pBlftQf3vuzW3bON+DH83qxdRyCY+Mge76K
wFHDnv0SIzIfX9jKd9g1ftpdwjcnC5C6mY+r6NG98AP5INB+mk4exgy1ruMj2QbzVPUAOF0a5Pas
9HJQ8jN/QEViKPAsxrIkz8pDpciP9y3xr7EiNviZ6LDK1CNAwqfAaSlZBJZbYZmWZYfVKOH5FuUf
vFk9qYTEX8LZX0qwg5Cv7s6WPWpjkdu5N1cLs2APoiVtu952mQFnmN+j9R+abk0sOpJiXHE9/doB
WyTDd8VBLePLz1Enl0hAQr9nPW0yHEWQTR1u1yQ6YfecbOSkymh38T33LWtDt9asklXMbVFxosUq
X817T9f7DS4xXI7vulsmT3Zkzt7K6rBpdYN0TwOxOmstAcOe/SxQOJBjEYQhIoqmnPNEujfWTNb1
kSGPAGeFYsrAqWreD1z/HlQT78p3kPZe9jy4usKFPKZ9892t7p9c+KvgDDe2O5/Xqt8EgC4h87Pv
7Bha/z4o2E73ABmlIQCkPDsWp4QGHepDKmDeDpSMMjLsiFwrwV7ZwREAgkH0YHsQ/FELz9DtNucX
0VrOb/bm5C79imr44v4ZgT6tYmRSQ6iFAat//6NZ3OGQP7sXkkVXtPHOu1fPOQd2qX3Y69WLssfD
VKYJ2Vhf4w4uam/02gmbDyOlC0Lm6xUI48ukYTW3Na6+Yhr+aNMfkeRZEhDuIZEzKvkb5ySd1FMx
azmo7M/B5mJniNtheTplr4z2qo0CWMc4mZ4M/FL8Mb0pY7a/M+HSRhYu2VIB1Nn0yPajFxn1FziX
FuXcEUhrprqbf3V3hco08WghxGkeFGua+y8XZL4rUWCtZUV4FuKiMdwKxgQQNjoZSwhDbf/B2sLb
UYE92MHhwjuoGP/D/8nT5XVff/NQwNab15IK3y6lRrmD9h0Gnj23geE1N0cH7ciKBQbwxn/KxGjl
Eze6RYZZINvrIvtqvlUl3y3EIS4viIxWkYHYUwgsAVDYnQRfP1Q8lIfo9e+lnAslorS8mpBpphd0
lhXWbprRyFi4bzbZPvF6DZsitgll3gRbRF9MLdVBej6Q3pe+TC6TrSn9qWQxgP0kySayQqsGj5Ri
/PgzVoZndcIphcfTW3z1W+x+OXpeaoKQu5y0ulSSa2BJmjtbrNFZwaU2tdz4t34JlPZEVHi8eCS2
QTQQQN5Jf7xteqMbec2Rvdn53DvrS2crMiBG00ttie3ph97rW974T0tipn7gyE8jb6yB0jjRa304
TywS3yd4wLmZcDXpqDQtzaY3bdUXUcZke6lVyH9yEB7+QDAAb9c7x0Fhi8lBgpdAAvE6AHXJWxSt
jIb+WGxV42YOHwwoHaMb9XRouqwV9ScGHMJ5BWh/m4L3gpm8PVIRf+DyrrJS5GKqcxW973n3Rg2t
G/IUsz/zOZB6CjIuZgipBmUTsk4OipvxhTOFP+8WxaEIkDcc+JkIGB1LG0vbsFQpfaBcoV//3yXz
LZ9DlTRypKQrvT73VPRxahCaihv9xiHf0S67rP+WqOSMkdwIIcov2z6qZjX65KVjgUHNfa9WtyjM
b+50D4HJRfYdI1KmBqu1RrlwFHemFNopjxn9U8VJ3Hykj9LMwjyFpPFfUuunZik+b/mWtaJe5sXF
PI5m1QcPfTxgsp8iDRRaHzv1BjRqPB0m7gvHaCBU6wAiKkEw+QTe3K+4iTETbOKQYfymWtCNd8Bv
32w9bPKYCkN/d/eXmHtEFrkVDDFESYIpZprKqgWI611MoFG4dDZzMD82ni2VLMMvsu5udIOlUgHT
eg9VQh9S0v+5x3tFB39lpk+XH4JOzZk4sVfX7//fXMRut6+UIzT3fmmyVyL17dY1ewLaqdCg2UGO
Rzv66D5lZCQ+hXtvMKBm+5OagPALHuoTaT3Xdh55o+pYg9nHIbnEj90IcWsTLTcmWZNE1oveGemZ
s5Rbz7yztE4HQfwThCioo2cLCOUJkTk/1AXpb+Q418yQNRSLlGOAqiks7fpXNZQaJ5kO3xoKk/4p
mDqquxdRJLSoRUjD6c/E/hAChJfshcx7BfADPM8y+D0L3yl16Qh7saLuR1eyNTBkDUPIsVnnyMFR
poi6ikAW/zNi322u4G+BiEOBxMyzyVYJhffmRs3Xf/2AMqRIpS9enc4wkPjqhCbhOLUNKCeP+xCF
1OhKxvwlMiQ5znju5Oiza77UuY26TIo46P+f1VZ69ENUbPwozeaRM5S8fiaIAXuMxLqXXcG2BtVM
l1OD4K5+60D+O/TX/0wykrw10VWdIFrBs/EmtNcs2GzmsWpCUlw89fMCZYSdnWcWKPTNeIsTOIYU
0EPYTBinvhLidAcCohNrZVvJQo+T3Wl1HvwLslsYnMvTUOlU652upRcLR0LE0PWBdI3hJJVAwyHD
6zZODfhGfvH1pjyRJ/7vcsulB47KtvqyqFWiy94XNk8hsS2I1hLeOcf9ZIqFni6EF34BC65Y7jtY
4SAQUZWTDfMLRp7IzAZEGCYH7wEuYu0CdKdkgR12oFpBhR01Ha3OJ1ngbxKaTlnrW1YGqi36iqsD
IXJ5td8am4e2TdJLHElGsD3gjvVshXks95qAjT0fIeeSPjN6UgZXK1z6RHnBmfMVdVptarD77rhq
sjWPV7CFzYAXXRQoTw/wr7mlGiiwTHHMmoUzml8FGVzxOX9PFPvggBOZlO/sKacqVhFPI7RfNTyf
hLwBXEGm/Td6OOX0JCo4kW04WyICw/frCXq/zHG/0HZlNdHos9jK9n8yeoMFBGcJAbm0vJwaPT6t
lq4ZlVQT1ne1ioX1ATqU4VEF2R86UvzJ/bwxsc4iSaJL7lzKzlTRfMr6nBxCd1F5NJ2vw7gt1WGa
knjQ5PQ2Rua4X+Z6RheMM0jS1BBH6VI39bkv5vf79yE/rfkiHEpCl8z04sDylzvsuGXpCwuSlFn6
cPhmQPYVhKH7U+LklUOELXKVVAbKweafub6uZe/fLZxNfId5JSXY4eIjOADCp/p4UkP0EodkgFf7
hqXSXN2SEwYVSaVru8t+CuIrhcqK1tet4s4eVW3fWjG1SGgU+jCYtWCylZkVq3Uw8Gv5LFY47/Lh
hKopFA0oIH3HDmqDC/Sh02pmKVENJmXMIGv2oxXd2q+yacKfRB9qZVEytU5X+G9oioq5OKUwB0Wt
LKaJv2heNLi+2lVWhxKzErnGk8oWHqvK6LPpxoKOWVPzBdPwW1w4hWCAcfBltPcG6yBTOzCedk/L
aSEP4+uh8APNGYNvKpFJEjVflsNtrDKsHrXd0twWkYfdL4ur7zxgaROI1Ngz4CEUWrngzfKwh/KL
Tns4s6EJ5gxH2gi7r1lSvAt6WpJHNToJPSnN2w0n8zFhIufW4P09xyRm78k7JlKiZw7/W4UpLRAf
KDpfCZNhwKQAebuyiz4aoj/88/3h/MhICCWHw6CvpbsCb4ml+27ObjWUKlUC5mHEOqBj2lS92ty7
p5gEaouuMg3Z2dr4EvajK4G2OTABgH3bb2v5Q5UTlrK2ca0/yg96GdlrIpOVwMc9Rk9nlhgle9TX
KKA38eCqQgk57BHL9bGFHNd4OpIaPBTYAw199ito7YP/50SWD/eMpEqjK8/OfBWqVoGKRDJ6Nyx8
bFTUSsfanKcS57QBAh0T2whI1xWxxFmoIfWq12fhclP2iwaF7Cu8dQFO+NSMo8DaF9XgohQ++ZBI
Uev8qZIKGnYSgBg7BfK/sNLXhB8eyOdBOrNfGfWeko+fUGaUnvcyQoaqBLl4Qrnl/5XjLyXrBbPW
NgdVLG8Gv5F6X+nEQ5dwSDtBEgYlpH5/A9JRPpmMRU9TL1bZhc8rYl+suap7qcED5EpbeH9hlVAj
6PrMzjbaREX8z3NykHYDsURm/yT54L0bm1BxSQCCdmwOljeXr1SZ32SA9QDpe/IbRkGYs0Srwsri
vnld+vwzqa4vyJJmKjCgvQjNvvclM3P05m7OQOM8k8LRnrGsJGT4kJnsal7E58i1DxGRcnAdNBEk
U3vyPpBPIQJUKtjfoR2ZcistonXkq3V475qY+SznQIk8w8Vx28rS/Z6kCjG+HFH3mXP18uak6ckW
+gkW7tLM+Jvfma9NY/44JFILdVSa0K+OthnuVXHEpRbmgTLMSwczG+jKdzVsBWZ/fD27mrlGrpiz
o4PV2cq5JN75Cp7tUCXGnbbHZJJPWl7l31f6A6DKpOXOw5RSZR+60MtcXTI0EKwA1O6dmarte+7L
CGH3C8PZoKyI++3GQMSSnrDwv6KcEYoxt/ieej4VzSuCKE5ITYILkxxexhoXeEXOdyrxh3OnK+pm
tbXKExnvh+IlFuVnpnU1057ZkSAxhL5Qp4jblRZUbh6zkhC91IKHpvPiPmL+7gn4ox0b0JWfoKae
5rUsHVANqSmLX+7wiMadc6pp7BdyHM3qA1UNYSe8goQpW9yjocG4Asiji8K0BgQ3na77bB/0kYHm
39D0MmekzakusKFcVlkZ9ldDD/S/4jwzNOCViAbOPOHnDtM6R9O+3S8uab/uSqTy0wbJbeOVMtVX
MKSddiGayS++NU7epkepSltYq8NMOkvYaaW+PjRzQvfYmTqcNJRcbcfxVXFmTHK1Q4iwuJ1iuNTL
sDjY3h5w0GOKtmFE9kuAxyDQ1FJkF9BKT+FFHmR8FRmAk/ggTp8W3Bj/m37Y5EF5LOHJF9w9idMB
yXLU6la93rjaiCJMxSkqCiKJS7kmMoPU7f4+yL2dSJww00jJClF2vX4D7yhLzijtODrk05ykrejt
lZFVaEgdqoZWSOIY5yhO9qrHlhny5juXYU8fiPC/AJZN7vyX+wfvDVp6snTjDq8GDLs3OBU9VUW3
W9J0vSoyK0g9VAdcfB5wZHAXPmyrA4FHEfzQK3cuky49vl+SmDq12HyKlfng3Qqlqgg2RYFj57gm
fgWgE/I2PTV6qr57ViRh8vp211HhpS7TakSSAAmSubkgBhE8za47J7Y3UiDlJlbh+v+Xlfouc3PH
4q3gLuwTm8h+FzDrW3cSxUj4E0Y51McN9fZdDbroXvygPgVGAvXx8m72wFjLW0zyLusN5ycae7Ad
z56W5IfaYh9YGAsNd4lrzQxBUpd2f71zP9x+nyRdNDJNAeTmEK34Iu2MuHH5b4uRLXtCTxPt5T6n
94a1pMu9kAzl/v981OcPKf7DINrWng0aGQrNkJqZVYmecR5SeZReEAKqO65oxSsMZke6bEVnRu/t
nsB8jIRWrtBOXKFRm8WUHD2l73R3jwx6Ux6pCICAxpfPPJt5Sz70MfuGVRL4qXl5TWGo25rRkUxm
wsm5Oe5GbwO75FT4l/PXctMTARzMec3tuc91gjqRh/2uBMUkGQLt9KdJqnFQNvCIMdsyzNZkL06L
gRG/iN9+15NfhvOcR/X7QKQLG3g7sACVu4prNiHAk4k6PT431/6X9i6FF6wsSPlg3njveVIrEIRX
367mTYJbkEWcx7rlbflzUa1Ia2mn0PCOAqJSoQDSuXRufxrZSZB0J3BaKTxBL0MZo5qzTYIhB1/B
los84Xth86V3keQb+aclwVjiGVfukfX7PBtQWPAuNxgL569cvidVOOl5HbndImtXH1xDNxYqWKVf
Ta9EAdaJ+FfkqLepALpKc8kSQTZMcZfTfYiyiKxW2FXMr2en/+puylIuoyx8qh65Uhh5m1XtodNI
v8CCUdQuKCmw5kLt4Ta7mr86lm842/mdbELRgmIUWlY+dPQPadnY2ilJwTWChkBKN7kEz4nXTy0T
TOXgwUCqvvRjavCTtkqxDPiG/5PpTat6po+64OQrGlRbm923hY3/F8NY47FkivZf2yLAwh+8kcg0
s8pt+HkaseFNuoR9L8Z1fgjb+JqHbiAFNUGE2MruUx2ETuE0afltp8I+JxTfXrywoBMKEl4yQ5f9
1BVa99AcKwY+LqUPHQWg67vJZkvntdAj0V0UZjS5542ON1DE7yhh1zKR9LWel7ubOUAFw3WLWbFc
G+BgkwjEHfglONh36Ou92Zx/3ZkxVIPPvgzlWMkmmGniCvADPduScVmfzDJG0/9VLNDxfR2u6GH/
c46w7fHhC/BtM0pmVpm8CAzvehjS7XBF5dqWocOMQbQdtIPmDtBW3WxboX65/NVgdzEnbpOaJ+9J
EwM67N9VY/cMKRalaJY8xR5iKkUm89FJpMsPhjPTK65dw+ijjZE6l5V3QgylN6HlPc9360kBNpC7
IyKvTUblrqZmqXMlqG2B+/Jt4HsH0mmvgQM6xT33X0QlyAkW67psG45KEGB1UqWjuO2sj/6Sbv0o
iqCKFz/YeGhqBCZXraoESrtm1oL2PedPMzFcehJMgskJ8JxzsF9F8/Mwi/idGuIhHE7vTnuR5f7F
jKDYJzQzFy/oL0p9BDSupMo1zd+Bt3f4t1MvvohUmx1Up4yhdIYoXA1cQKlViMbXmXShK2X/LXve
lD7trTtURqqS59aCCVPs0aPqM3pgwh4BZ2bvgFLypN20WEIcqtOdsSm7SNilD4Q0xLcRWeAw7rSe
yxHuQYVysExNjSTtmcAQgJqhKrfjMYYKh/eeiMwkzwJKvlOIVcZlEXJJ6LXP5a0aoGK7QBx6iQ/o
vVYd2081CTZJ9r7RMnULVOc9qeoNLmpkPfGlymvNC+TUIGmJoRvgCUGEc2AVRyDbtpObbBz4/DQn
fBr49SoFLn2rjQ9C9H4faMfPiaGSsWCEB5pvv+vGJ0Jp4MuMuqYIS4yBWqqxVTX0/njzHyZD0eP+
I+WFd1tlgk/s6k64dcGg+JHHv8PakXG+makqTyg+r+ns6bip/Y2vRlaYcFN7NzTT39e7JAKNqnrS
k3W/VL+a0qTLXf+buSCMcWgcj0TJFKLJWTNYc+aJuBPWbb0NTfX4hICsrfpEY1Fa60d0Ov92GFR6
T7sCLAk7e8on+RhusgWnCqMAwaBg9jOfkVS4O9Lv9IpL9agAr58rbAxImj7KltY7W5IRDbhvDBpu
Eqt/SN83t3464PS+hWwMt8HkvekEbnA8UccKZp2ltUMCrRjy/cSHf3L58gHDQQCs5LdTx7wWgpQz
I9yoN0nM3mRN6Wb6maUDAHpB64h0grFjv7thbFDFWwNNzm40O2xYWZh5xdLCgMhtxN78QuFUbg9w
UEaYle3TMaIHZCprIOQXwhEc3cUkM4gaXD6yAD1V96FhfF5cYP/JcPZazpZx+TBg31/AbIdvXp4K
KTqhgHbDtyj2Sk5rPeM3NBYhnAOQIzlufPxW3n4Sn64DE3qmYRx33JFK0v8AMdoKFacvpxCWnxFV
Wsa2lhRxsRTXB8tcscZ/6+K89lLmTIJflCmdgW2s85M5uEIyeXWUyljdPK6safLmmRBCDvV4M1do
74fJSaU4aTHfc/Q0eFHgcuzDoRNeaFPmPnYSPpMvizNXNqveOIsHGJVzT1KYTIuAzdJZV8Gxfsgb
txPBoM2oyToqTFioWz9ylMQyyHYV+a4N56ocvjHDmviUxVTLNpmwgYhf82T5DQaTnEtzg9zt335M
fFXngpMG0kmmX3BjM32SZHQExRoDVUrZXfGzgi4XSRXhtHQkJ5lWkD1dKEYEnLlcwpD5UsnqTUSQ
QtprsYUVnssRfG0T0cXuCZh5Lin91+V3f8QeQeN3DMrYwCaCJgGGPCPSU5Z8+jdFmD8B6lH0N4Ac
pva5Jt9INZVAwJCTIKaCorkbeEIep+uV5T49uUvt989r5d5bUmrsxCShZYOzL3M1x1T98XWRkOSq
x4ulV8YFOAMwcXk2ICcvvWo+oetyEKo+CnWfVnZU5z4PA9UUqEHxiCjv431poh5znSP2tJLttgCC
PC5wtXHtT1YNXHxHhQYRaP9XQlVAaT+iJvh1f/pZlJWh7TVGZ9dzGsH+nE4zyM7L5J5W0kboJ+p8
LWbxLvC9sd4Bs5yHVC0GbSwuh3/Fq8Ykdo/T//hUotv3hAXIm6+f/aohHGI8pkSxpPRvCSU4cyjv
sMMOBbNzEfoJysPrZLdq50//MygRJ2CGAzC1EcPHnak+V5C9ifXjdGqdWEO6oCAw6B4T8exV/7vD
XOUBozGpQIXN5hgHjW0GmROkY+9BtAnFCZL4sS/3KEvyGf7ZjX/Lqd7Ls06ySi8c5qbfgUNnithi
HTKIFwA7mdMoiFW08iumNqufd5pYkOWcOhLiAT+4PKQkUD2rXnt3h+xbxkMIbPk3O1sxIYZBjdos
xSUVBLNMfelOsou+UiW4kZTVnsi12EaY/KGtKHbXmS3rBbyDWjmapt8+qMCpkmSiW8ubyz/j5i3M
rXlTbKsNDHdr5TyEXIaC0OrgALBygHDnY3MKkINpl/6FsK62hEbCBN32LU/lyL3rRjeI5IwlAnSW
e5de2dEB7KczPDUoGHgXcMjELQESB/TMVc6wa99rHZyI+AU0YIGW99R7DI8+Tl23Aw/Sudc7ARYZ
yDuhrmaT/VT/k+OOsTj1t6/DOlzrhJzYsHUDACtHqNSn/jX4pZkVk2W6oo8hTNZF1ei+G55KkSsd
R8KvITjnYPNzBQMX8t4i2gww78+l7uns4202pQJcHVFblj6qIaqpuQ/66GP7klFa1b7DPihDwNvC
VPE8cQ8SwTtqEUDNoSJGDA1RMxIVuH5lLhfpNHCI/ngFwmJd/UyrQb9MqjWgtRE/K1EJO94dVntS
p0raDZqyQwdJqoAHWfUY+8F3lIX1S9RuE0UcbUJ41VQ6N9VtW2nlwciKD3b/cUPJz/YPAtWHKVpM
4jSgmpZp5tfAmXr3yg4KuI/aB7QT6rRg4hmJY4WFkAYn3CYg4HD3+mYKNuUu23jK+6jPQHOqaMKs
NXVq+nQmOMVbn231mg6rmvNhh49Ag+8WXi0sR+cI0m+YfSbCPo2IVqzmlRQN+dyyC9gU0p4Wjkjz
0Mx+t88rsROyJDPIc5ZR0kE89GPZNlSaHICFI2EUfbRwhsw+Ff0u1Ect1TigqYJeXtXaZdWe6B4t
s1G2FVsRyFoEncCmfvHfWeFGy1FnUk35RIkAXpkdb8kWJJfwaMM9sb3KnBkR1oa0qjde+QN+fQ7/
21UEebOcn41O/7FsC4kR74OsJ6oH9VWqE07+dIgAFQ3WzH4RB6vL7aKfbcrlUJjb4hDHl2FI9U/j
1Rk1usj5cTPo0CTsviOnp8irjQQtrqb20Ijg+lmebdYNR7mnHYjr1yAtaZ2gzX67zSPyLwCOUl2Z
974ywHKsC7le/cl2IpFKJx0tLch4KYWSPvHgAtpNaoC1Dpt7TA5pmlQSg/tspuXTiHWqUFGQGdxF
PIya6j7qcp1QNJKLiw6SpjPq7VfHFz9boVq2jOtAkS+fX6nd94/1hnfGyxqSOn/54h6kI1GlV1ga
v54wVu+JQKg3Vf4ljDaABBEDLRXDFkZSGHzItqIzAfUUjfz3PVV17o3HfCYAd03F+4+Oj+9wzJkf
adPO775t9hvChrxZHcIbiraOZg+FUoBbhEqjECJ19/aeBjklwUyrNXrcLUoWbTMMqKWA7KckBn1j
0MVttW7Dzw+NPbKXi/U74R87u+9pdxe3Dkstkh19tMb7frNSeKh1OeFiDXAyZFz5PsyUDrgKQRhQ
+IqD4fhtwEsQO2E/Uf212MYwDFCwFL+3qzTwyuRXjq44AzqXx+YAD2HiJkmGwh+aP68b/HR6CaDh
bs6KrxDvqamOwDOlKCUlRnRRpqfSwWGwVKxqMttVtunRlnjXxijVAjfKkHHcxTFf8D1/pendP4VI
k9eeh8V7/cgHkcYhdHtypBXHlA6G6AZS6+gJ8AkPeh0WSaV9GMhfOhod3m7yvs+lMzH7lqOqD4n8
5umGTu0P/oUpKNb+9sPhmRq2t2hkpFrQmKenlg4CwGimEepqG965bVVThTlVr/dwOjo9vsytWis0
e4O81ucXPpUX41ptI4NIdai/9WfdI8M0Bb1h2Y3lLEhSKZg7g8KnrYLQ1OPiAIjTS3Gkbqb3BQ9J
/bsKiT225a3n+bEOVdeXWjMhayb8pEigI7kjpKX5ryvmLPQAHq6+StCzYmPLk4l8ZJet9dmH+y9h
ex/kYEWpAr10iLGgupYNqo1VHIJF730kbBnOtBKdNq1bsBU4Y5N8iBM5CzGXAP6F7sSYW+oTIEoJ
L8N4ml5CroaOXS+D0kVrWY6NHwwkG4ZObSkib03tneEVeIogd9Nrhxj6S+m51zEOnZAxWhhS49iD
4TH8KZvMko4N175f1Tt5qznG06YVQMYQhyNnU2LPfIOTXueM8rGi6EBw84S99twtfc60QnPOBBue
FTsejtFky8lSh8gLK7Ig1Pa3DvdvVdSrG7a9xzNt4xyraWgSvv7TZgJb5L0CASD3rmELobduq90w
LXr7EorVzvNSSrt+2/rMujLCx4wuk0s0Oaqbky3oNWC6Hk9KTOE0JFkfH6tOVG2nAT6uaYxEi8Rg
BG/s1jSeEAMHYGv+7CH9haTLl9ZKhyCgWvhK1ys7fVXRJdKEdn6ZhYhsO0//Ot/gJKLHBb4+z0MU
eHHQnPAKE7EXNLXXi8jIWuxXWV2wyE/XODXAstvXeTwstQV2g8Xw2DPvCJxf/SB+GrhEoxhLXWbV
W2vWjSftGcohjYzLP1Ha5O0hwA6G4fX+XPMt5CQG1OoVokg1R+3WvswHKqDAaPlPb5g9HL2J/JE3
4RNGUpJIzj36AbQZ9O+w5EwtY6Cv8Qb0vnHVhwQmKrvGWbw6iNCQsPSm79e8KuePnwSTPezgQ1OF
wBnxP+ABRAUnZCv3IcrjzCKIA/Iv1D70jHlzzkaZkozgAmHlra6CiLbrSVX9VTVPn7bj7tQBBdtd
oE19OgoKQzMxNI5WOk/mEho9YcabqRx3jRZBI7zvqj1K6wYWm2UE9BJwJBRP2fpKnoWAseGjfYW+
iNHimodeiHA7LfZo94nISwBX3x24CW0hF0U4Dh/YKZI3xyLb4QJtb6Zz42Wpi8xj4EchfPyA639M
qDmMtfLe9JOZEHcKVrgP0PPPXzmpdbRozuIo8HttDj+ve+pgvbklmkwgT8wkRjXAzErg3zAnvDDl
Hmn94hJHvXErN1u8Ijxwa0CpiP1KRF9XF1EAjSYYWc0tWJRMcBrF7EpNnvz9QnFEuBwBQqpeLVc6
/8EwyJNDK5wQDuaP398tMKg3G/bJEBas8j3MerGevN/EZwPJAQvqslRXpPsd9ebok6D1N2zwe2JB
lRThcWiMBADuUBWRN4GclAcGUZvRcmYHw8hUeIB8hZHhABho6WSak05wHmvSg45fTY6x9zzv7JuM
7l6iICPf+JyirRflK8Y9Qb9xVnvcp4HDGNa+Gm/2lSaFcNfpyYkFAbuvAuNPa7ZOBhTXkGfC6QH4
b1dQgx1div6xCDc2GYJnjURAo2P9Rt661DGD+Vdtwo0s9kgFfzJPxRrAxeP6uNFmjF+9HSpOD+U7
GFb+CX9MwtOh0bZy9jkDptwELaD5oRwL39yXnZndXhgfeQdIU2V4iwvJUKVS/kr9TwQuT2Pb1VEe
vpVyWjYGJ+ja5TtJ+ouoHKoi7wBI8SU5iAvNTn4O4hEy5Q/CmBzV5x/lpCUY0Xldo13HOYmyPd5g
w1ArtmD/wjQUrgHmRxLk4MMx6hdLzBRCV0Dg1arhYM/8g7jwfzG8juAbZJSSjcy6cd6BEGhFy5D2
Xxp4ROWIpwmrzv/6Fm9q142AuryxIZHPyTahZa7IQQv9JYegUvAnfJXZI/tUfhj7mPogpMWNhD9O
nUIs4Rz7SSBXBMp8gdJU0Q444taHBLv5UNAbJQuOZxIjWFyRUGobmaUZ2/RHdmPA3TSPjWLVWpc1
zJV7KZPQVaz7ztCmy6eMBS1MpwZb3BUj3ZIRYhxQ4rh7hU8rhR51RXNUjmRBTp8ox1bSqZe5P2vL
/Mf6tyQbB35PtMRNAJBpoD7x/RKF2yIyqxfyQ/umcs7dul/lcHNXa9tg3pdskfbxFaNflV0EIL4U
/zjX44BiTbvOEyu4U+mMMpQCAP0PKGahaLxNzhnhQS5V2h4QJ+9e60vLM1ks2lBBpBbt2D2DUWaj
aGEgkqK6IGCDgNC7HF5/Npqpw+3GtEIjnVWM+bs8SbCsPN0dOmXL6ysXcovXTHpCye9i+7O6LKQC
Bhcw4HbM7REN6OpvRAbHOPENcii5Rs6cDEfo62qL+Ue441EtNgTcN4BoVK0mclRMKAmBfNsSTV5h
L0U/RogIEpsob5tD/55QotwM/6Z1BahG+fxlf30OgEgil2YRBccjbEUunsgD2Vn6pcNfHBvazjYb
4+yjHkDwRKb+zhY1YvqckprYb1ZCXqNV6/ih6q0VX61Dt/9Y6Q7SMVaZXu0scdsqL3Q9G9KmnxGs
okGdX9HSYTBZbIZYJN2zF0i69CiYXHQyiRuRRI/4+m3TUppibvhmzOytEoeYbKsbZk0e8HJw8FtZ
sWqPseOiOoG8TWCwsv/eAlE/k/6cfC4cyHL+uLlLkyL2e9iXf1L1F6qkCwcIwqW55lZDZzpY+6V/
jCWfJ5kinWlWX/hJLD66h4RZ208vWxH8aCRHf9NkayVKpZJ4coMD0Rx0FUfZnVyYxAmuRQVVz5lP
mHP9VmZUzZYg8I58wzNJ65Pk0hlifeMRewdbpodF34Qtkw/s3Rge4Q9Gzb588TkDlJPZXCWP1QAX
wk+y8rR1N32YGGNshwXKDB/gCp8d0dkHFW/7fIlOmBVyvXkBinOderz5Q1rcm9YkgY4RL20DOlUi
q4WHCkZLRpAu3oijo+9CBVQMhdpvveKin9SjWmgiLkJp7/LOWA4JuYrL3gMtNgBTLpBsy8j/uTlG
gsoclJoKOuFtzXCieAXRmlDB3HdvnOFC760NQtjIXTvobgeau69B9/sq6r5nKmJlqe9URxaMHWnf
foXfs9xMe5GhNYf638xe+G2MLK/e9n44lzNCO7wm8OYxEbHvvWTVeNfuBZB5oLcJGzeGEG1zcwIo
YFxhOiFABuoPuXmqQWMdp1gHsSAt2EkoT/t1iwWS5mK6eIDwuTE02a8Q+oSo4vtw19cNn7umA3OJ
aJq9Xp5vCD2q6XpwgvE1tAnMAVzbSTHJH+MfxR2mZGArvJX42ZOoWT/wYaIPJJ7lQnb9YuEa58eS
V3ZlupvkS7wY+cUwot3251A+6jdIYGBMTF34Dhxs787yRY+cozmmS2ETd3FUWKFhTJDPspZUgGvG
66V8Qmfu+M9rs0aUJ/kGTIFnm+C+HhIvNTj0QnE51LpKzke0ufPFWpbW+nAI0Vshtphb+5/K4Im6
0LjJHF3F7d37mjh22rv0dRbpzTRMjA0UM2TSZV3w0qQh+yVEFmp0AVZM+reYlHdeA9zQ/r+4zM2T
s+noDT59gqMPGIfDcarVvegjmwporOAYzxhATUEYFCMJ0NlV0RCrCaSJaro+VJghMrt4DOUfl2jd
6JP7IPjj9ERDvIU5P5VowMpNNvyoNAfQmla5Q7flm5gbq6tXTUwUeTQSZqcF/3FHaSeCZS70d0J4
UIlPG1WVvVONMROoGdGqlpF+HsVMfAgG96TtHOS1tzhceaiivMCxCbRk8vpvgp6XK/FMgTBMxL1t
CiNEQL1hhyyyI0yYchGfdqp+er7CbiHaBA6sDk7mP5RCyELFko3Hegog1krU0IMFiCVzUni0zpct
wFb24n3MBY7hnyrrdgSqhStj+ULjtlhGBS6ZA9TOVZ5zvRtwkvdNEeCiMYznMHK6dI+FJsnujWPF
/84Emv4aI/GV7bsROumrictQAe/2DQcbgDm/xQ/EmVuvfzyy5CfC8BnYQc3pzRH4f/oOSxLsbuDs
yi6nXAGZ1txkDXT6wBxKljGjBQ6EZBHzGjjVw02Gnp2NxxKVC5KlOEZwaiilCrMO/MCCtGbtBIfw
Z7IOUh4FD/NToBUPGbQ0kIkUrmcDQ4koS49bi/oCOMFSoxOZStK+MZjiI0hopCu+cm3GaNCr/Mmf
N/0zFQxKC6ZEFCoHM3HKRD05OFjgqH0FIIWd3QQLTVClGe/UdQYtLuoOB+7DIKrmGptcq9mNm0bB
/r9XnFA95eQKNQuSIF9b1Ou8nHAjRDE3pT20yFEQK+Woo/P+gDMvDheiLavfZLU+ZFaeX3Csgbr7
DbHSHKhtXZxY7sHmMrgtlHVGXnVL+/VJPAaJJD1gReRFX3uun9ABaQ7/BN1X3hBm21t7vnhn3wL6
Nr+DH+XQGc2r2mm6ltzeqBLqd/LxwidPs3tGzMXtyEN5/vtmTj+IMawzdt58JjuQALn8hzpRRWaJ
MiqhrREtyhx+/ZEXSLMeL+OS6nw4lV59Nd9ASVRI0pegIejQdSNxQBZavfxNe/qg3o3EAFXrWsSw
d6nOK0Rbn2uLQavuS+StUhIezl0PXb0kdqYJTj4kskIpnwJJkqOnD92QFV+OdZzy1NTKNnbyqac/
YoOyHQY/z8vByPzvIlgpa/p+mGGdFUMwoWFyluMQTO4zVd3Xl5LNNDFb2fU+v+AKdnxUQKUgApfa
62fOYvpwDTBaWtc99QwXBx3cx7eNDoXvtVdkYrHyN43/3VX/8S4+lxqqA4MWeLVnKHLLOdKHmrnJ
WhIxbODaQLPjx9dBlR9XrNATQBUxTLnQPlUR790w5JcKtlKTLQ1vtSoG1655MKN/42EMwp6WPUnj
yt3QhtRvKBtgkPWhbTLlbKs5pKg5vTzsQ0i8/WGOqFVfIXcqcEgYyJWbbyj9CyUq8B3tLUQf8jzC
ZLmMbWb8PIMB3b4DtjXgCA9azMpTD8C3ewnjFgx4X7K1LEhljKfM90tCP4YBWWuNq3D39TxOILDk
Ey6J8/1lbX12LEo2QF3XK2RBwg3vMwo92fOletAdCMsiqFxD5wCgjFHavJM9xqC5nxVppXl7RRdt
+p/KTPSSHhjezsIHmjzxDLMnFulozace1CB9Zk26T1ymdlzL2AI/oKSZDVJy6Kmi3iV7jtHz5Q/R
o8ptHvz05hHhoqfA2AD1TNkH1Tm893JYvv41HJDXHfQ9c5O09s6ephMruMfvcIattyedu6SBIyPP
BR1sdX01knxZamZdsFFygtog0LanpZ/7N7Teq7Dmqav3d/iNG8zRO8RCSeYdPYk98ZjhAnuFwVu1
A9/0u749D6M20aJPz6gy34ARqMU1VmNWv0u/1rwcQijQsWZQFyUmMH+32Dfb7jH5Jf5NAvWcHXuq
SCU3C2TgJUg0FdHEMVkUfdDTkC7ewZyMY6omPkXJ6kzB1G5lMu6eKtM2TSYtoM7tKUB6/F7H53Zg
xzKkVyjyVFeJyzZOlaf+9/8RDpC5b0N5W2nUaoJf9fM99WO51JJ7W0e3QfY7BUre95LMMCbB1ZI9
L3bDHns1BL25k2CpYG7ccjV/puAWR603PddZ7X7S/5laV2A2O8NUq/18e6Qk6c0lcomAmIbhwJCa
lPNoPd+KU/ZWAWN8woENJexSvXVuAsYJNMqMS2m2W2C8VBnUQDiVGPMMcERz7Bpjr2M4xxxzJDFB
PMp2UlnkzPzPWGGO9bRPQz2ng9K2gyOlWiKWiuql5LeXWHUwcs0iGPYUvnvrmjdgRh9tYglS7gUG
ZweQ9Yi9cZZiMNAsXybvRD6+2+XIQYX923EyfAVU9MXFvXyNn8wVu3rmZlLSsC4Kco5BpH67cPOr
E2VEzzfzsAiXQ5JDJF7+6ONVKgSGK9vZAJRaYPhig5csZbqtSd901Imploj0l9XCOsA7UCNK4ZVB
eHLAcr8N8jpftyGf9eL+izpS1LtObS2D506R17fWr15+PdEJ7w864YBUH/ExY4cRvnAfg+XmS9PR
Z3PIDF8nKak0y9scZGgMdhces2RWJk1fLDFtHUix+ngDpEz6m7kiIzp0wVNHueg32JpYNM72RPHW
BHs7pU7hCsN55xuw5R7xUue3tG0qha4POLYrrnOhGEDX1Sd+klGxys8rmbXlOJhhz11vDe2hq6RA
lnmCa0lq5FJl4wlQOZOvHA3xDlI4jPnd1P7pul9QlGz6lTxohBOYUNnoijLdFIkZFv7TVgDXxnhu
Rp+xaxSbU7WHUNFujaZ3U1VspJuTmJ/X392vVdcsr58f0VdGxuykRjlMwNCxryX7MqolaTeY+juV
ngN4sn73ADyNVmVQoOsoKAySYoePy6+uA46L4OXiRQPP2caVNfoBrpoh1cq01ybrLSITPqH5eS0r
FyAucAdGBBfxWnBjfpJULunAyF6hDBBYeJNRhQUQFgrrKUDNbJt45phUpcN1n9RRMycaHpLwZ2Mc
fualqYI/rYvhivMCbObsNncGAzy6OQTFM7dvLgOjCQjSwfgDwGsQPRJ6Hz+DxoI+5GoiPoWgyeZd
npN87DT9RZy9SIZraUG0OWL3OHdZnuoSb0dIXdOVHhvtsvXl5kWt3+L3pdNkMRFj8d4P/pijVbhg
EpXbhI/Jbj3IwwDGf8VOx28YMWOYHmkOKcUYL+DezFgXLZCvh3x/ICoMtjy8hrioYcT+gegrpFV0
mC4P0jSOO8FnZiGLKSasiwM5z78QOnJgI9VIKzlm7O++j4YYskIlaQU8/mygRMj/oRp1K9baW/uQ
9yYZtSodHCBtEhJheuxV+46fsx/5ZeJ4FF7Vs7FdZTo8CYi1tv5qZHpkLeUPPFQhNmrEU4KudYYn
MFRkAjLu62Hb0F4X32+/a+ym0K4DQupQ679R12jDkcwnymXHa7BIbbLCpYrmTb4ZB8BYdVwS4QaP
861WwJyQK2W7q4UyTY5PZfFGwJuSR85qnfAugVQcqr+c3YGPfJbbE6cPm6gs3HMLAkP5NtNf3Bp9
AeUJL2bfHsnD4nKn3Nkf87Y97DWnrtlgoJYpU+NjT2ctUDM8bYAW1myBnzebW60cqhaV+DismEwL
1T4tfLDpqEsFqx/gNGiKPSqHz3SZ5bOHPNLACX8ZydMFcWf3OQiNNjQyt7WDD/K7uWFZW15+OaaN
yFRYqKtYUCIjx/6yt9xFyt8Bwqkpk51GIq5Wh92TqSIvy3szg5Nb9+cwfVqM0VhLeKPgOgmnSBl0
sRdBm/58wIwK+uVw+2/dbgs1vKtvPJPuw9w56q7QYktVzDp6sDL9fe4k1+f6c2bHGSCSb7Y+ZtuO
n6lri0QL7RO1RDvB+xTpcqXyw09HzTROAiAN51XhvN3a0m36XiwXOegRDaGcyPsizURWesrI8yfe
mMniMvR6aDK2feyMzhI2pNTZUMXYmEk6ZVCyK+uE4dBi20US+WFCoAZgAFgN2EMLV/sVW+UOhtbM
MRFlI1Se+3Fd2YJHuIcQO+aG8jO+AvCwSkHoD1j2GlOpvnEAvY+5e3tqgVJBCuks6mhT9GVdyPJn
JATM+xNjilAmEJPxvsypH56MuG+NGXBs/aTfc2+H7dqPG3CnP8kxc0bmzBCjvBLFTSA5lYArkJNk
/5gigWe6xuvGfZvNUJlSehAnNftry9CZ1Qd+hcLgWJQfU88LLw5Px5QSIBNoTOE1wC4+7+3YMfF+
feEDNAIVmcYuEuCxtLNS9wOhbPe1A5CIT9ooPMYGAuP3pYyFwgHQS+sdlFyEsdE9+GNcpWs5LsHx
3L8fEdOuOTKsa+9lfc5E96gW9LW98Xxdyd3KlFxzqQL8XkT4Lcz6l61nlOlvXLYJkY2nCtZsFO6/
QNBOnP4F1V+hRU7C7sf+UA6yQDqgFohOWFiwEYwPD1cUr86XvofUGb74wEN61HYsuYjdTk5sl5/3
TCU7D2hMrSIwWFFHa2dKWWB4+UnLZFHmag8ZLSkkDw0F6iNEFjw11AtsvFqFU1h0laTBwlJ4sP7Y
OcikDPAtIvMnqgAkE98dp9ulyTqt5pogQt2JrdNm0/mnVUmowKQibz2HxNlX5m5geW0ej24AsDi7
rCKokMi9hNk4CFrBHoAlm5bw+/gfm5k/BDg0rlR09TfDESE6M9GncRAcvi1PuJeUjAH7iNZoehJF
c7NRFkHioblvaOdHN0Q7LrOjjYcIw8/9bKtwvJ888ArxQlOj/Vvv1/Pn+NPiGAYWgruz5FZy43Bg
V/gT6Y1osKMmAVeZLYXBP4CadLh0gVJzHaOpfdOQb/m8JcM72kzuKm8qy+dzS90pJRZSEPVizbia
BG20if/1Fe39GQRWaq4v/ckgpBKks2p3PuiKB3ytYIktwF5MapJduiSkMEaQT45g+SVISE7XHCbJ
0aOCaP38980ZNafCG9yEbtDqA3b6OOYlKiYn00XmhAjuBP1QanKqBbAygGSqcC0TD2H2tQcvb7k4
HOG3tFbzDsqC0yGhuJZFtIYBvJ1iCtKMA8qo8espGXrB6Hlj6NWTG0q+0Z4Fnyp75SN1zh0zU5cw
S9ix6S9dfqNWT/H8qmjNHmtUPUXgH6+aH/qNZZgRp198kMMqJvhOdrvyWWuFvKDkvz5o5pLvBcG+
Y62LdX/rJrXJOwq9IvNN9RsiYM7+maeF97PPHnuSJ9LFnW+HDEC+rNC/miY2rSsgMvVrAorOXgZ6
hAd/1pzYqWwg33JD4MJI7x+37xpsnDh3h6fkGJUSRyPj+lHEu/823xUjwoGigJqcMPhPphArq2u/
kfQL+ybjX1xC/bWFfgxfmb6VBAgTvlLNXGWiAANcZ5yqzFjHhkWYZNThHYBsSsNVc4FL12G4ZMsz
0oXtIVQ0BKrVaKi/Ib+zZ11YDUKY3F96Nhe7uPhrWZLbTSPOroAbiGzdaDraRMraq9njr75o4QqC
j2XGeanhaMNxbJhDLlXJfd/vifvHz3K1AwUiWX7ELqYpIj1GS40iemETJr+S8gqc0dBEyhg+16nk
GlUWVct+jtprcUZuI8T4TiMikY3ZRX6oh5xrumPn99VfWzpFpMXmn0pWoHH+A//y5BgExaLry6ik
aGkjxYtUw6NMHz3ZgVDmOgkXGTlzEkop7RuZsX1l0XrQS6u2Qfx5kECWDD3pc6q0jZAfcMRCU8WV
uTxJMGnVSudWAsw3M2S1Q7gxNxQzE4hQ1fdo3SqI+R6Mxm3D8Zxycz9sP5C9D73uGlJ7odEMHR8x
lSbK0Vd/oQlcCD1rGImYDvd+uFzjwJ8hp2cPFEUKywwldF+18cApf0a3P0tXEUmtzPgrForjQ+b0
Gq3nUB4g0QvyozMHknHfccIcbzVxGRg60lprYF4tkV0Yln+jqPtZWRCFkX6477OcJyPwGclU8ieL
2IgS0m4F4gKwzMsGuzW01oE/v6qmeFgoJGW1H+MY4KpKBM7ubYSLxPeTxWRY01hYhHP4QU98mUss
Tf/mNgiCCn4w3ZPBa6vPJwDcsTaN1jaOwmOTxuRxa1QefZRarL/ra1LQZBpDKzRb4wKpZO8H3gb3
NPvKlIwzleDZSI9YaXjSWKUuFHMQZza9xDmme1DybjFOUioMELEHzZCfnv6lkDvxHE0Uhe9u9HYp
6rY7upj/vUpmmd1txBi3gX38IKHGRzt5hHn/qz+/3O2753l+djO+XbG/2G64oiE+PeQAf69BCpas
o4AEQZZwzM5KnJzCygg9LyvrrShL+U/S2OLYBeKF1Nj0X1EMjQhIweMTlRd4RnKFJmSdAniMt1jL
/h8NTFW/b1Hj6s9JJda+e1YGCbY+YCQlbC5xumiKmrR3RBlkm+owztkaocPCUp0xvzsJZ3Yq1UNu
u+hrBF/d/5236sb7myI1bTA0veVOmByx2OECPF80iu6m3xpHemBXZRLNijRRFRidrE/+s6o9Uxvs
UdEWUKSbssX9ZqTmE2Zsjm3jTA8GKgC5pp7+JvMtUXT3zXe4+KtB4+oO+5yZSwfJTj1ubNIHdh5X
xNMh+5grMAxBPdoINb5c1k5rkN4Sous7CITg3j3lDKLoOI1cmxsn0Bq1fdCfRckl0lV/ueFdN0mb
CqYIAzEcnEmIhhmAFG/JLPmMCEQIWQ2itXScj7SdCSqKxeDrPB4ZDbF9tmqTNEXChfvetk+BvZq3
9cLV7rpdsvnC073x+assDc2XrLUPLAq8JVxIDQjPUczQeWAEV2uV41Zp8vT1xyzk7yVXBFv/3Ui8
itQeJTAesGtnzztNx0sOR//gAhxeQmrNonGAzqd6hlXm3ADurtrEc4TFfl7+f6b+u8jShUYhGXUa
fv3OtLFu+kkC600y3n+1nEGgqPji8A82b4QbPLNuaV4G/sZwx3vpCZrojFsUNme+AHT1DiAps1pi
sTBtP8P/r+iyu1Ta/ZIURChWPz82TVbjhJ4JqmF50W61C+VFoiu5HiyWT8iXYXSycJ++hbkhfvha
OEsXSnysx2eveb72rFVpuE0NgX8eHRmObAJW+Xc7bGwMyZUKHpUVM5hDI8rg0QcyGXy8MJxP5UlY
Yb4LY7K5UjXHsF7f2SBOn/JTVhgdStJVZVRlblwK4UChO73U7inH6/8liT1+pCZrnaJgrLu/sPJ0
OAGO/PDBLuiylX3weqq0TpQsnMAdf2zap+WkEoNlH7xDelqS2e94PP/dQ9XIw75xvkLzxNSnBRfj
V3o3pZrl6ikYcCquyF+1yzR4gZZriK1FDd52UYgoSE/VvDrUnaesYqZrIMoiXCowRLh6SDtQITtw
WhbPzmqOOq4Pmy4CiYujvmJ+oNSZibYLXVewMTCbL7BSxiN+WORItucXl/zqqm4mMoahoX+90jv8
kdi2gPRIxscAKpgFcLcb3RzAJVM/N5h6VQFUSTnlwFtPMHADdlwUCg7pXS2x9mpJrlgZPhQIUlN9
rogrIaJSyph6plMDDHLAgjxkkTHI5eQBf52xhtW+35z9eUQRmEp2W1GkrHeIQPSzpymdkoyjP1QP
+9tmN+xBQJI/tUyDCuIa8ucVhET8JcsOp+RUt8wz61J7i27xW29SRttXNAheFOCG3vWFqWwxmxdL
P2aStSU8e+QUKKTlZDwwn+8bgUK39H62MLbFCWLid991orR3TxdcUG9ajDDE9MbBVXIOIrynqgc5
RT9CCvkyhfSMS8z9nmhtejcCk2rh3yXjMxr270nju70rnajtwCYzu8Ci0tSCWWofmcxXpq920oWC
6EYDhsoLINC/u7cBeDy+YxuX6Hdf8TuP18vVZksC2s7xSrzFKw2EHVa5j3MXu8k2AFCD4SuOU+is
1aySZO1yhyXX+OWVqk5pSVi/yJMGK94MQwNECOMbJxeLIIMtqBNeZvOz/ENodDWyEElfDf+UyZYu
PB0EJAT8l+Ngs8/vC0zwQxwlYMSBKwWzB5Z+hNMVlBfWtdT2b0OF9nyDvipe5KS+IUZ5POrSgabk
U0hn7DzsiXGeXHb0V42iIG/1A10RwsZRt7HAVIVT52I8yX+Qo1oWE+G+QHizxdmX/XwVyAaVEzkr
GsfMyilZ312LuWJvDjAD39mSDGQ5jHHdWMUzefGIDXtlvZPyGMt5ct9iYlGqG6o3Fu2Wr76IHuw0
vRKIhferEWNwn5LkBGLxPZILf6yaJnSN0JyVyuvM+/rT7cCYkEhGuifh8G/1IsH1M/bxpLJP5kGx
l0IcX6h6iA1b1GuhYLsARBjOF1YxaFxUQK/i/fStp3l5IFzUnMCMFMjezTY5hY7f1R6r/FNbUEux
hE2eENjWJlMkhHO+fhm3/IwIRXIw8hv0/K49HU9Wqg6KWy4M+Zty9jzp0t0WTM5bk+RguN1H03Pu
emOdeoc+vQI9m5WyCyTCVpYqAv7EKffNykBYJwYWlEeR00ix8PJOJmep5sbbauc=
`protect end_protected
