`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2160)
`protect data_block
gb0sU694jcjA0laK1vfw6ujKBJ86cKNfsMiRjggol5H6Qw5dkkM972wbiDMh8fMEQGfWr1wrPC0h
v8dzmUA6uSCg15GsYgC+z3vyp0tlcWsFYOj5mwsK49lX5y3FinME86TozjnbMZnVRsxLJAi+mPHa
BWNRQXnY/uLPICvVZKlZ+HXlEq/t64xL1bdKTZ2HPe5ZWLuqQ9VTvFE4fRge5+DWykZ4RbK87TrH
bn6otSFsbtj65eM3r16qxFUSC1m7CkLbo5YcYNdAm1W1sAwm6/oTzlx+WCeUkZ0sPrrjCzCgSwwf
y+1Xxk6TCygh7gX+ByhpbJQt4A/yRrh6VouhHLPVSm+R87OTD+XNBDS3KWaERkF3/9t2c9qsEK3k
FTsjHdExl0txQjKDGXzscOhK2OVSbKtGAuW3wwm1BrJYJpaXFO6gmsV0Og63LPXn+jxTPaPERn3P
YA3b0k3xnkA+/WsAhcLMIswZhdbd74C8ArwtbPUJNqI6rVpBtreSeKqNYZcR9SH+X7YfC0snw2AP
ewO2bHTGKFBVWOLe3C2VfsTvuBwqcJNk/f4Z0DXTRa+tlZqMBV020WCpdF0JgeHF9TPM0IopFeZn
2QAczDoPChc7r4Cb6YlnpKsVoywFibxvtZkQBkyJ6GbAniQoP55FetmNSHRXVGKFlyQd1n1pErEs
clhCuri48KFu9hh449WKw3dPI7Tda+LSE/HKktjnYjvuVo4h/3KbFpr67VIp7FtDxtGaf7G72iM4
JaACT4BGf29XH4dhSEu0LRoJyHkajC7BSht4CGvoJIFV//YHHtrtfuohlpoPrxrwjHDu6igBBACH
gbzxrfLGPrSn/UulQZhQemdK8YSKPIKm3W4KibobDI77XIyQr4mfuxNEQ1QVKzyUVhJWfuXYKoRU
bkO6OMRjcZ+zMuJbWnNlhlPJ1iwjQVH1ByoDNeGf07fMD2nCU1JnBc07GzcP8Vmpcpcu9xL19Q33
ahi0cYgMyBskbCmmRkTaVakb+JvquocpzKyLsMYHwKElLOtC6vNusVo1niRd3u1VZika3iqd/f0L
aNIrtQbhcLByI+HDY/AX9xkuhf0VbLecCH5fEb9WgVZHY2z2fm3ndJQIw5YMMUQLlKYTTXb1nEeO
2iRGdsmBYshUww8u5jhCH2fDam1tZFE7JRlYosCEtpTut+xQO5RlS4ZdLmiTrbSM02tSICIWV4Ig
3gStzTGlysCNSGSqhGTTZCVx1S0Xxu67GP1AAXuLYJxTEdZlh/UivCYv8qpiFFEAVd+vZuRVKvHf
ikoGT8EZnVpOTo32GrmLh0egamJEWEa3CfC21Gzh0hlduuIEO1eiivUjtYM90ki4ELwFzaYSO6pe
+mZQwhgwhYYS2w0RY6hZa2sraDz266CnrxpXG2DqW9icAofH1FUvnOUUe8O/iGdnnyuiSzXBAsn/
GRcGE5jqhC5CBckr0YXvobAI03AvmmWdvY8tERfl/NW+SFLcPxTKo2xn2bmYGGigHkM4SHpExIK4
YQmZi/1ov3weBKgaezUXtiS7+vbmSf7KdVdzBgyVDi45uqyclW8+f6PAW7U7uhp3CfM1d1NDo2Vg
zRNb+XJ6VBSk1s3wX3alngM728qfzfrTQSuIajKffzuns5DNtpx8+lfjFl9gEiZTLd4F56FWmONY
4Yf4+jZX/l7upr88jR8XheXhDDXudN0EVZwDi5XM9Qao1ywxA8dDo0V1EiHeQ/2x2L7eRFAekpBM
Nq9M7bUvTxvDw+Lg01hJWVZmVktXBXnFpWdIoc2RMFRzGJbXYWXZR4GEj1zKrVG9DAAMW0DaLgvM
2GPFdNM35WggjtQUk6UzJ3ISoNu4tdpKjKUcfJJwQt3+8zfJ0kij4T+2Dek+iZaEfObxm+k13Vzv
yqxHyRBJ/N/DB4kVPVaXxA4JOqtHoz5hV6RNVTCtAFICvKTRaaXYnTHvzAzlptG0oBd6pn/S1HNL
0EzaQNj3KcqFrT5OAVmi/A7AlC1S+5WOzD8uotO7S6KvBMw+/LLRLczY/HLREIzIK+E2cVZrUQfD
BbTHwcxRbD6EQ0G0jindklQ+Y/rKIObXPQB5wYQ+nSQfCwbIDhuHcvO3AwScC8BJmrV8u3yexbTF
AM2x4tdnqdL3LC0L/8a/WSVCzTkVGnN8+NpdE98Xn2NfHeM0zmK7eI0SJKBFVsRzBEdwXphGGsb3
O2jEMmvndxYw65J2karrItpn+cwOQxnFuK+knqUzEwUm3RVHyOXMOQQRKYxRqaOfe2QMTWl6xL6I
5S3Kkeqf0LqTswTdvhc7WQ0+BK8JeyUH9WHizxQfini7FzxkYwrCnVa6Ot3R9Tqyy0wXQsab/dPJ
qyYGV6GdlZKz8e1pl8fMJEGT0LaT67LxCX2qmqwEikRMpVQTg9mwKLPFmeyQ0YlTZLkuPSq2pxTD
jpgQfyVqicj6vx9ZRYfd64gcjLqMeWlY96NGu7VF61/Bb2q4P6uk7/t6vg0NFkNQqpDYuy95qk+3
7kEOi7+MW5ZGSFO7HGvrJA1EuPlwzYQJ1AYCKNH5I0zJnEzAM67JOdax1Go5fZeItmlPoXD/okUn
f8CY7eATu4lxLc26+Rc5wqvHOT53/QXcgY3TYnYdNxVkgu0B2ezb0E+ZzA2v+StvU8Pi1WVquDHI
MdQqVOHCOW+ouqY4Zi7QqNRUTrCDQEaLcz7VtbHZbnNvyM8f+qUH46zdsDY6CR/+r+xFv1q5YsAp
uuPEhifnk7EsWK19Iu8qYJn74qHruUyAlce5sQGJOLOy/CD3kX8otqprFyfvMCvjjCnkpPsCmE+A
TLKciIpChDcPJCN2vFo/xatOahl7JJ84I3TBwJnluC28RzNGO41hu/hpCqLAr5FBDoX/
`protect end_protected
