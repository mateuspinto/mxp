`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
vQacocEPGjyKImnnBzSOicBNr4LryveHGCa1mlpHfNwbexpLAuRfel/8WY0iwNJHByL7+8bqjRna
igI1W/+iQDQa2Qvy+6gXbjofEVKq2IAFHg7jny4q9LTd6U0scsHV1hP9XDOcWbrCbojqKd9pKxgi
rnlCd8Jqpp7klTp6h6/YLxn6UvT5pHXfJ458PhmuMfvUd0wcbPJTcmaNVAQbd3YarB6yiS9xVzGw
LYjMblDZaP/1SSYE+d7VFgWRFlEDrsVl2POYOA47syFNM0p9jrjTZ6PD0K7dIWF2LUwTkeJ1TDqL
xaA3M9qJvjrpbRkb8AO4unmCS3SRTdxd+jK4iQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="O1e4J5v/PWGkRih5xHV8B+pNexZYS3G/COJ1QxgxVGo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3520)
`protect data_block
6RwzyUJ40lngvj4Qtp58xgGiGwW8aCmDhd/xg3fbv7AZBYElYcRJhbn2I6wTtfYTl24wXfb1z21A
c3Ld7x71BRzwRHjdBFMLlBk80/tp0PPehpo2hnz/hpiSTUN+7DteSvit6PWi4Fh4+94vAKlirHuL
7J4ln+c1EPpb41g6xLJZDL2btXmGJRohosmi9oFIzqtpmQFCe1ZkiAsLDiC8Vo4Y+emAGenAV2Ty
S5mtlnMK7odqhslQYpRPykela590TUyeHnJRBx6PdTLugXhSeJIKVNkuYPAidlCfQAiEWnjpplb1
VMmHFqCfWj6E5tc+WFQzU/EotOwQ1vAn9xlF4EbHRrWNZeOHq9gmU8sDPWfHfmprXTfsHHI2uUsR
U57LFJMQwnz7I2NQfHvfw3aQfAhn05T7hThPevydecWB5QSiKFzgD812L/H+lHwulffdP4dLdJ+1
th3M5N/mE/FzBC/c674IaY0XBnyB885jWkeElpMF+az/84y2bnW2VmlP3Xr4+mqZVKTEhtXfP8Ed
EgagC2uTMVu4jD1vG8cOPGli9b9VpZ0jCimYHbez0lBiOtpLE5M7UzJyyULGaBWfBsAluE7Jhvlm
URzsEqhm5uoqs/Vjf6pi0tNcPxl617r5LrE6uE9WBlAH1KZr0uJRsoXuq8SKANkBczm1WoYkDcrq
Y0fQaoF7gfzk504dsb0XD+pzT5MLvu+nCYZ/9+CHXtuV2yw7Io/PR/ofF44hCB5okSr3b8jx7zAJ
927wy1Aj+JIeb6YljnXYDJ5FEGZNmEXJhhK+wWVyEIUAXwtvdQCXwKk+u3a+sZ/y1QJWc+k3Jxke
LqPreY7qZ/noWuI9hm/u+ovohjx8Ta/VD1Wf6SoQw+jDf8VQXhD8aUGrppMO3/0ashdyzruC5C3c
R4xjCRkl1pVP6Qm4n25LGeHibYSoz2vj0YLK8J8Iqg2e+YjNFT5v4UNMUhuJuBkW73ed0mTIlZRj
FmsevLw0kCLZCep1nYc2Zomz5HTGHoHq8fuX7993Du7eL8mfWL0kPwFOv80N6G8dduSXDVGpZlJH
uHTjLQQ1/UAB0S5VpgAnBRsO8Lq49G69y2K/uQQaLKhedde90TohGIDVXgYu8yjLZYOw67BIMLMF
m9bMRwgI/+fgs5rN7LYrGcD5zNy0nijxKMeyBuyhHWTAOvmkWRwdaWsWr6yZCN/iVmaKbqSaafqy
HcR0sZGRYiL7smMgx76J6asdrwwhaOth4hqqkpwoLZrngyJUawc43ypTCbyM1nPIsDqg95mykXOH
u5136fPSHqSTJj8kJzwoZ947zAIIY5WdOiRr0UhPFGlscS26y8e28X40DCCc76WheQfqZqrU16X+
/jStHo/gNLcvahLPphiU7UWNQDg6Hi/jfY4fziSSpLy/63GtGdQNioXuKMSIjuCJSe6oEAAWD/gu
gH9HgwuVbqTe6+HeP/fH/Ftx0Dqccv8NsotYO5rm/CVkOckatQf06ykFfB6bWWR37O7+fJpOGbph
jX0mC0oE+H54jxpiKNnAgD1faBXrvMYfY6wbK7w6nHmumZ4dMMU04J6cHpMi1LHiN49ct8mg2JNa
iStNd5ZbULBSvXtgRB7bGZCg4yRnXunzshblo74fO91Pm3h80Xl282SY0vGEg8hVH44mw/kCd8h0
3Gua8T3C9wZTTHCAlBk4xfxHiVBHANtA/7+omBDxIg1kHkFbTNVsdxWWbcNoFMgyAGKNtmwB2RZa
1zEWuIsn9LZMoJ3zm2g2xkeX64++zxxQadqJaLccwvrBV8hkiOwiEAYMM2QFsIUEafwDYLHmqZqe
YxwvREwUJpjJ15J48EXCgsCN6NxFPOjHOtoxLB+av4H3Q1p9qbf0Sfs877bvFfFqAWQfyl/0bgLZ
gWYECMI8xwdQp0omgzcM0nqUW/8O01EXdoKMnO9merktcNATIbu1XG28fuESgnluZXMMVsBpX+vN
ahDM6p64OT9/J4cM8zML/qswJ3472VlCwQR9Nb5tAnFFc36+tVB6x5hjg3X5g/I7xCNPOlx+Ag3a
N4ScDyO3pfMsQZmWSESSRFEiqbJDPHUbVVeih9f+esxD6kFpgZ5J0ka70a2uy6hJ6GQcrVlcuMxQ
5Ap1/WEuIIwLX/zL388Py8lfBQDaN03+A0tXs+e49uUNXM0kpPn/ioHwOw/fnSGUqDEdmbretkmN
0deMNyrXsF3jMenaUhUcbnq2Sf3YeW0Z/hZgSp5TKS2uNTAP/L9QWOsud4g64j0BbJaRpOC4qQk1
CKXAQrMshHr5NMsitkC3/Q65CRCEEmyDbxqbqsSA1HVfcT08sdgrYEjL2Q6cD0HipRoC/NbQcUzf
4do9ysCvsdDdpMg7MVIfwGVnLYe58V7qvOC+/EOi3dJIkpflDrTmhPUHwclx+3x4o3kfsybLzeMS
MbiZjVoQRBWjIE/RwCRVf608R3oYpPGt+VvDbPsm0Jo0QrOFanWggFBFnHNT6bHIikq25NrgtLM5
Q3poHDoO0i5pmMiZIdl9iLE/h+o/7BC7TuuUEhzR17glwzELbDy2AxljH2qeavab2miJu8RNRBgc
SfgLgZqu8OVSGCQGCFv1CcqgS5v7Dx1Zi2+xbAfuhVMeWbaWQN8yu/sm1c6ODoOJcMluHmqpv3ai
YBZoDZ5R6PuAI29NcRM3xvtNnuTG/IszTMNpGZoV/md7WLhqKbyhqDmt4d9/5BhsVHZKImZFcpja
1AlDr0UZZ26APgA9vpsGBqgcnEgAes+FKMvkwOVgwH/b8WjBAbBwR2Bvq9STVlesOI5riSufCd1b
ed2IZkyQmXd2RNjMYzJyfWrV2zztCo9PV6LqIjoHESzuUfozP/zVpmdtfHoZJ8HjU1+NaFhTqu57
H80G8nJekbyHj2U8TIgakRZ9xqYimJPFv+aTwxs+PMAitgSjq1Z+ZgrJSXmfnXYpoqp8a9zwaK0j
DhEmc0S7ALi9Cd2NgSpJO9EyJ+wunE7wIagS22RsVhJpzWzFW94CSYb+u4bUeuSpf5zy8Mh3MV3X
DakW9DHumEHqKhf/VscwBXfWOBSkhjhX5FbKgaWpqBSH2HVtAScEbhYGeeYUEklVQCEO4KezHrFN
ZnN9h2QjXN+TjUZ+/bVgS+RQxBtgegK1gdMi97qlQ/YYQe/hKVCDGfsyGaIwsS2WJ2Wut19XnFYn
GVXyIHYecPqiXhtpkaQeolCWjTuLerocIu7TmtApQ3GiAnqType0TGJvi61sp0aktjzyJVmzrUu1
4ywD5mY9yR2DOltS4XDTSQB4Y05z9oNAA2lnXmOuthK6+Dmr3NwupEWcHn3ZQX9YfaX+8+QbMMdu
8Tz1hHz7C9xXDgV484wxRPiRPq5xvaJAgeEFq5/Od6u93mT14I9eNA1spxlcy39AnHZ79gxvYuWo
MSCMYlyqDMGCp1NB5YdQRqyRIPvapjk3CQPcWIygz260o1vFlQ9VQPYZdkRV0lwXZV/XqSzhPXCY
NbD0kttNNfL9s+Wqqal21emxx5qr2XZnxBMNBEu5LYg7VQuCUHP7Qt0v7Lg2uQ546Bv7Mm2t+wS5
kKxS3mD3DPT1FRvLFlCzdoFWemC56njHTtiB8C9Ej2XspegFN1IZLXZn+7DtKKxRYwJHAD9dUgix
3ttO32cPUmKJJXthu9wznX0E5YBC6J3CGpEAv3BENcxYgKtcuHlgpHPZFOAdHQIxwnUWwFHefb8E
1MRiZ3D/OEMWwQ4Sl6wDWxc6ucODx9bnJSI84HNZNqktEVzkBDh6ZR7QImCr1OHm7QO9Un3Y7FNT
UlRhqqG+mxIBLocAmhqCg+/mREsbGxOEbawiUPM2KUZl9p+zRoLLnLHQtH81gm91ja3gAaGTcQVB
7lRNkGmu4+/iTRLcf/42AFLrbIm7apB5om6A7luLgTQon+btqBNslUouag61WIUSi5UFE6KDuNT4
dfQq7nkkvcUgU/TFGPhhybdwSldIfJWWAJJ5L+cvRqWeR39BmP8dLONpi51rrjfJi+HTRUZevOOE
v+ojOfHTFwe1QBwifut+Rxt0uUzRSalcE+AMRIwDp42aM8srs/gqwIQmgOqpkq1zDQUo1sb/GVl1
M+6hPOb3cxDSa8ofqo/Ic3MgIS0K+N1wzP88AxUD3sCdxyWL5pUi1c0QLfBNxxqcKSRcNMbjCz9x
aOVvr5ljLs6hyshisrTT+IkmDM3DhV4SZ6R5TOTFTzG8MjJLWo4gZ8yzxJ1xP8uTLZkIxjansU18
1Xf/dzpzi6KdJFmU7GDCacu3LIUWYoN5WMHf7XnTh9vk66dkcCAxjpnYFcBfmS37TzHAqFoL5ySp
JBrsVcfCzSI+NoBg6+Y8le6Qra2yYYes7fC3hGaQ85fV1tVulMDRh5haOTzhXX1hpXttLSW/Ua9V
G5ij3yXEOnPXRipEg19hAI/OdQ8ZjFtumdb1TU5VWSb7Z8lP9k0gW0iIQe0rwddQWyImoYO7iBAb
gA7SgZbVP1msA6fwhVH71GSb3W/jkjiLg/8PRi6RchbK5VYc9DtQGT0vkqmYU0sS23nQWxYmzISz
5dBzBhz0G/TCR7a83CP7nfbeNceGxt/8W2dpmR383IBpIgiWrSPqRcOl4mNzvSuCgtGWqr6fz/r/
nhHOR55M6kgPLpnp3XO1lQKw9tYELAgJ0aolw9COj7m4uqhDXdS+2aHEAw==
`protect end_protected
