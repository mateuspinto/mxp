XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���=
>9s3��-&0��٠� �L>x?8��|o�����<����P����Vn��g�k���٨S��c,����VB��K{o���\�.��a���� W�cD�䘑J���3}�6ơꬻ~G+�8���y_��*��_�NS����E��l�E��v�`�ڮ�p��%��JW�B�2�[�0ߴ��)�<���83+=��X/��2A�O"1�1�;�|$�RbEТpWS���hɘ�M�L���)��I���z��h5t�T2���(��V8���k"r����b�Q�K���n�ҍգ󜛿'𵗳�j�:��j�I�M���,��c26r$��U�xV�֥�DkN��=y���ߊ�4Q-���{Y�E%�����{��H����(E!IU
?�v��M#��Y���R]�/Q<��� `{�MX:o����FX��zPp��H�֯F�<���P<3m��
��9���`O�3�Z�������|jZ�����_}W�PO�Yb!Ңd��D��-1Lfxu2/g�y#�����	���0_����8*��	Y&�A�.�b��Qu�X9/,Η��x��/QNM����+���$�'+��o��2�`p��;����YK{�>�icn<�/�w��X�*R��%����t�Ap��Ag��FQ8wX�ƚkSnzY�N�&���rk�i-����4�~~������h���[T�*q�gK�Ok)iy3�x��)�j�����n�<Tg�T�<#���7Գo�+XlxVHYEB     400     180�a��vL4N8�cA�nM�$݋S-� ��K=PM{��k@}�Đw��m�i�(沈	B�{�#��)������:{ @��:���H����u�d��blW�0	=����U��ަ�<2�昪OcA�S}��tp��ꁵ�-$Pt_̂������;�	������ NL��:h�=!$2��g3J
��À�W�ܓ��Z�~�5��Ѭ}x�QC-�r�&U	XJ?��vpvޙ��M�8��;�}���>D�7tخ32FsN	:8�>;$d��VUN0�9�w���v�'�պ��_ض������#��9\<��.�WM�`������2����Z9�b�%�Tv���LLӚY�Y�e�9w��&J*u�XlxVHYEB     400     180���-1�9��2��>!ٮ�@�E	Si9*��(MZ�OX������,�;��X�==��Ǭc�
`M��C����wv�G���<4U���`�"��l0���F0��0���q���Ux/�B���|pG�M���jhN��6ϻ�L�a��q�H!��$4{C�
щ0�-D/��a�$:�f>�9����|�4O��O��x��������>6������ʥOl@���9�ܥSaw^c��N�ܩ�K�s�"�H��Cf	�����K3)ﱾ|��HJ��9�X��������̿Y>��~�0�̀^m����dJd��G{����˕)��;�a�k*_XO���a��j�����ї��q�v�B��aِ�DwC|pXlxVHYEB     400     170���"^�S/g�)#�jyT64
�*�;��Eփ��Mp1��`����|���O�� .��p	f)��Rvմg�E�<�_hB������;2���=�t�5*	��h�
� ��쎘f� Uc8:u�7�x���+��^�S�_�����^>gGy��v��:�8��������U��c�M�h�VW��V�}�ퟻ��F�"� ����;��ҝ�ɓᰳ�ie¼J�}�>q���!����#I1h�I�10W�� �X�P���0���ֺTE�L��C�\3s�
D~��Apw��{{au�����$O�)yB㓚��M�-��4��x�%�H�T�s�QSkQ���X����F������XlxVHYEB     2e8     120N���uκxЦ�����Ww����Wdw� 吙�|vg��ש����_1�e!;�&C*@8,�BIn����AJ(L�s�n@���arB�d��t��y���&��E1,}أ�T,��bdو��`ڞ���c����)>5q����Ao�Y�4|��a��5*�[��qxƎ��c�h�C;�՜s�n�4T��XQҎ�� �6�d�ht��� ҵ����`�RS��۩�սi��M�Y����.��ِ06 ��q���� �P-���:*fHB� cm�=��