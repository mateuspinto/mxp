XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����h5�\p�C*.px�9�&��p���#���%��T�8�����ӜR'PF˴W����ݠ���uO�D���r�eQ�{h�M��-�Y�$���m�-�3y
���KT�N
Mk���!�ڝ��金�%�NYa&_H�����"_
E�	Ⱥ"�ԴΣ�G��#4�f摯hxJo�z�c�l�l4�%�Q��}���� k���Q+tq����<337|OU,zP�u�Pg������-ts;�?3��[\82�)��AY_ݩ$�+S��@hLF��0Ww�[����m�W<����W+�i	9fpJ�l������;CvyϤ�^"��m3��K\��t��`]<b-��*�G�M\G��B�hBm(K�����h�s��(����C�u۳�g�t����m��#���0��Q�T�
�n�����_`� �\D]�ky�C߸ s;�'�WX�sY�!�/�O�~]�2�x��eu��|S��˺8���g��}ip��rd�C	��=p��
H���z! ݔ��9.������Z�;glnߘ
N_Pj���Qm��"$��v4��5���c��?JS�G�?�A.�Y
�8���Z��k��=���&X�7��r����G%:��m�b �,p�V�j��U�qe2\D%���Bu�Pc*-~E]Ġ�k͈Nd)j��rgh���}yC�lY1�Q�?3�^�Xlrm'h�!�oJ����Z�B��sP�������u���ލ�"/���y���_v	f΀i���3�vXlxVHYEB     400     1d0��n?�/�=i��5�·��a!���l�ul��3�f c�t��S��,��·g�2�e���>�7V�|žP=�i�}��Dj��^�g��A������E���Kv� ��J��6ӕs[�h��99�
��HDй����3<h�V����e�x�����3:BM��s��fFa,��c�l�S��!�����x��'��&
� �	� �A����!���ee̬<+��ST�G&�Q�+_�;.��cΨ'N顔���T�����[�F��`��o4L�_� ��ZɅ��N��]o��8����%�)�R��ʚ��c~ɓ�mx�,γĬe܇���FQ��?�'c�$�ujD����j61$��Ci�H�#��Q��wi� vl� ^5��G<w`���]� �B=@�J/Y=�j��o5N�������0��14�ᏠB���d��D^�;k�^4�XlxVHYEB     400     110�Y��5P�.�A�r?�S
dG�2��&��,�n��C-��J]�/��]�Un��-~�>ﭩ�X')y�5�h1VpʺVz2��71�#a��p�2��R�w��������#U�MsV���^]�?�S\F7D����N������n���-�]
�]��j_C\����rG�]�)e6 2M�$��P����_���Ϋ�Ap����/��k���w������}� +��H:������M@f]*�����a?�����x�ŰRde|Z��h�E�XlxVHYEB     400      f0 >{�G�aٜ'8Ld����T�������W�^�Nw���_��63x+D*�$��dVV��&�D��F�NK�'�>�YFE��Wj��;��q`��ɶ���a���<"���=�Kߤ�"��%Z�$�Β@�m2Z��<J�P�[���m��tsby��ݺ�'�����#���;�ϓ�F>��)s���b�9��4�4���t0~\��;��sY�6����v��)�T�~��XlxVHYEB     400      b0N�;ױ�خ���V�x�����,h�1z�̣� t��*�0�Yč�#N� x�U��r�����RQ�	8�|��oshy��4Jq'=�٦�G���no�G��M��aȭ�~�!�#��҂6x(��̘�y��m���D�����\�_hl��Bc��u����B{zuZsD=�X�[XlxVHYEB     400      d0]�,����hM�4������'���}�x��O/����Ež����&���UkE�:���(�ȑ�I$D���)����"��2qR�&��A��+Ò���ʵ����R$��8f{���u��0h�7�2��m�	��tRԡHޝ��ґ��=��LZ8X��si�4�):�ˋ�2��`JW�G�r��������N���E����(^��`��JXlxVHYEB     400      d0�;�aD#'��Kڊ��fE�s'��y�H�n��y��^7j�B��m$P���oi!��4�l�N%���J8D,���5�ڱd�J�S��x}���#���|`�p#�`x�����H2��:�Hk����mQ�"���=uy ��K����T=��9%l��,��:�)�r�����.b.�HXz�_�Ԏ���'��F��{��.��O�z�XlxVHYEB     400     120��}��P���]�?`���ֻe�X]�N\<�q��Rw8'u�C��;%� �E�&{��n�6m��\}�N���*�T8�Xaa�W�۫�����C�AB�yc�V�֓�@/|�:����J�Y1�ڡ�MdK�����aoH�L53�v����N?�����eDȍ,-h�P�/8�Ĝ���Գ����P!F�	Í��{x�~����#ԣD"���r!$
���1���b�}��ۏ�������?���^�@s����-fh
-�VO��\�S.�9=^�v�ؚ�p�XlxVHYEB     400      b0��Ѡ+�k=�ʌ!�h�Q�W��}\�)M��x ��Rm��Nqqt[�D�����w��Q��gh?[�"���n͛������:�߲���}�y�bO{>˼�0k�L�&���z�ezI�>�?r�����v���p�G��/V��)vv�c*Ԗ��6m�>	C�_�V�(�1���8Ș(��=��XlxVHYEB     400      a0��h�p/��!��n4.#�r$�pq��T����M�U�t��;�z@��m�Mڼ��UK�\�t�z�Q�F�su[�Z����AW�CTZ�!���t�`���(s����2�S/��_�6�����d�f���
��ҧ����!Q����|9�Ve\~-XlxVHYEB     400      d0	�S$�g���~b峩̢0v�o
K"1M�꾏ڡÇ_��=�R�k�F�r5rLF��i��V�-��&��{���$6��
'�.긭3�i�Ndt��j�7�Ѫ�yĤ%~�H��ǚa ���"�J���a�#Z+t�����'nr�o4R=�&�i隯�	պ�U���ah�<�$�X�8B� ͏/��ZK *�� �M�v�XlxVHYEB     400     180\-���B����AP���S�DΕN�w,j׏�%��j��}�Gu<��N��cD�"��؋#��!~W�П,�N�hp��Sɰ��11�&u��!�X�����J����&0��hȩiظ��~.7�X�̾Q�_t�u�X`9#��������m��	�D���Ѯ�j�1ڈ���?Zp`j����ӯ�X�x`�i�1���MD��)��W Э�]{����m~��{ȦG@���B��*������ �MFY)d���Fx@� �O?�׋�Z���Ȏ��1��le.�@c��R�'��MX����}p�ߺ硪��g�O�^=�*�jAc�ߌ������ܳ���ͮ��!-}-�U<4d��I92/	��kU(�*�����y����-aXlxVHYEB     400     130/�Y,������L�F=+J�M�I�UlP�(��i̕�2��V��'��e�;*=�<�۾"ѫ��}!�
�Ӥ���h�I-J�j)C5z2�&�њ@�H�Ulr�g���{z$��1n�@.���~��V�r����e�E�Od�wƇ��<n�L���&ecxK�H�d�.鸎oS�{��>N�	��`ۨ[6^D73@̎W�tF���r:W�U���( �1�S�\��X�{x�V��П�),�]�<ﶃg�@��_�T;tҳ�"(6����8ꑠ#�sŞ{�BJNv�h�	|XlxVHYEB     400     110��FN*~U�	��b��r'�r��2��Aڔ` ��<�i}"�I%}`>��o7�壑HnrE��o��j��@�Gw�l6�k�����d�L̇��ԉFe5� P��|+��I}f[��z��銊�sR��׼�k'%.�@�-�ّjCh���r��;"2��~_����JB���w����T�è�*�^��$4a�]^�*��9ߒ��=���G)#��V��	�0��E��'�$�h�kG��J��E50\������46Q3ޚeYv-XlxVHYEB     400     190�%^��	��������'�y�^��k:�_�yޥ�[{�y��M�a��Z�/�=�/$� ��v�Nz<aw:nƫ�0P��k�|F{E�N���27��u:��^ɿ-�_n/T"��	ΒF�e��"�l��f9UF��F;��_Q�s%l��p��3�(�#�1ø`���$a;fH �����QN���g|�ٝ��9f�l���}�
����g3ݽ�V����4��'��B���Ԯ��`JJ���ዸc�l���Vnk�i�.�<��v�����/OR̩Xesq�c;�{��G�+�������Qy���3l[���1=!~��3�ul��b5�/�Z������ؼP�����?�_�n��2Q�Q�|�i=�51�7��Xm�@�`�˝�XlxVHYEB     400     110���-�:سYi��Y�A�م�����}���i��D���%_cެ���b�p׵�W��EaĦ���s�w�s�<y�gc���ye��y�m���!����⑑#���le�!��)χ){��EU�l|��:f`w�^d9KX,8�]���ў�N�������=�3t���o ���
������/�����-2���z�d!s��:�z�ܪ��*_��-J9I�la�cA��V����l�PӐ��ׅo�t�TA)������ܗ{�|�XlxVHYEB     400     110�kk0�E�d�J�6�U���PbHߩc�*~`�ζi��a܇�P#k�����Ѽ�Z�G�`g�`�X�%�X�М�}/�Y
�0��D��s��r�:�QJ����T_L�Uj����$B���-E��n�Wh����x���d��=/,�m��rۋL6�)���&�}�|��Y�ݼ�>�ͧ����b������{�Ǘ��*@N����Ej� P�]�6��-Wт���&���MZH}���Dw�6�È75"�/&�f�~"�j��_LG1؍XlxVHYEB     400     110��D�!>�Y��ٝ��$n?���'"���ŵB�L�k��s�3G��� ��2,�Sݕ�렩'��-�''��7P��>�=C�6�P�d�=Cl�&����'�'��*0���}�s	 )��
�$(	��ϣ-f�%���=0^	"R�D_9G�nN���H�����ȹ��C'��YӚ��v�ů�+�� -�* b�HY�D���.
�r	Ҟ�5�،�]�P��y�Z��.�P��_�i��uI:�g�d�H��9Y�G\������Z��8d�8��XlxVHYEB     400     100�����
�aV9`�OD�E��Փ�@/��>b�Y�
]�5���)�������������D����v4{=H��.���\��q�NC[[����S�2�?y_l:��@�-�l㣙Q�pV��q�;�g�}ԗ��u��kk�N)VQ��G�E�{�3~P߮<�e!�uN�=Ҋ��s�6�[��8�B�L>�Nx}q��#~]���C0ـ(Q1�^�t���g�������!a]_���vf9�gl��L_E�XlxVHYEB     400      d0�W\� 5�q(պ��4B���d��RLu�<?��%t��%��!�\a&�Iь�����r��>�"0*L����n�V�GH#����$�+˯З:!$�幤#�<y?�zɚ�v�݂k[T�x�Vj�zsi�_壊0��	��ӟy�R�_k�A��<%�+W�J���za�*C�t�*��$���ֺ��
|KWX��gtW���NXlxVHYEB     400      d0�
��)��kL$��W����:�sU�+�n_~m��֚������%0��|�֖��1���9fET� �8�l��>����iCa�߶���q��q>�W�q���@����	t��cI���*�=\|j�WDO���"=W"9����J.�����3��Ʒ:u%��¢���<b�e��;� 6�{U�W��;�Ÿ����LN�����>�{ɬJG2,NXlxVHYEB     400      f05Q�>�YY�71�7ȸ�t|/�T�ε�h�Φ���Ϯ>;�"�co���K�Dp�`peROv��c�����_�&��zO�:st�OVd��9Q�ᰨ���Ϸ��;���ef�]bx��Rm� ��m\�y{ĉ�[�Y���lk/���o��<��=PxP,�^\+�?�i�ڢ�ݡCn%����ߙ�K��:�	�UU
W�\��0�g����74��T��j���S̔�d
��p�O���*�XlxVHYEB     400     160��iؗ������<W�i�o���W��(
�Ҡ��b�-��*�k�	&�p�J��H��p.-��X�c���-X������>Ĩ��L�Ax�@�xۻkm��i,�.�#As+�%B]�i�Ѱĝ��g9�컾��������M��$~����K��QH�C%0R�y1�#��;��$_p�1EՖm)�t�t���$����<��pE>�/�:�����-=皫я�5�89��#�:��+�[!7@��C'j<0�t��v�-v+b��k��K�=g���m�>�2����Y�x��O%���XeB�Y�� b��b�\�)O�~ ���ݖ*Y��5Ô��RR����8XlxVHYEB     400     150�"�ٿ��ݽJ�n����}�z,D�W`�R�����F��7j�Gy�{O����S������Kج�E��h���D�x|�R�+2U�}�Q4H9u�XB�sc��|T?8_��������g���6?ޘr�\��^�⥦4/�q~�5��PN�*g�~[�c�BGt��z�Nz~���ϸ�2�IP.��D(�gTC�T.']���t�Y7�fމ�?�1$A�q��	�pUJ�$ܒ%�q���v7~\��cj`�s�p��PЁm��z��zb��H�4��[Z��TktڃIU]��u���>�sk&r��}�"�[��̫�ȏ�A�����b���P�z��XlxVHYEB     400     100�����g�P����6�촰>{�qD��t���)�i��D�Tp�QL��s3���S�����מ
�c;1��6��OuNRֺ��1ĊmFr"w�T4���c�s�wD�B ��/e�� ��;�u����L�5w�k-Zu������S��/���f��zժqa���C0��P&9>>���*� _�C�5�-a���s�#B�N���{S?���V&�flt��>�$�؊d.�ᵑ@WB�ن�0����D�b~�XlxVHYEB     400     140��BS<�c�M%T�t�ޛ�܊ş�/ǒ�&�j��n-��a����Áo4רT��I�md��ɜY>�S�
� �+�W��'��ݖ��U2�cZ�Ln7g�M�A&���B]�5�,Q�@�~��}�Mw.P�5`&:�j�T�c�I�޸��:е�n�$ƀ���}�lN�����&�p�#o@�q-��Ph�ÖɄ
݈rT_^�,�N�ɯ���%�u�%n��f���|�Q쳠��_BY�r���{ӕ햃_<)p�h�m>�O��>�]�@��
��}p�HZ�5��n����
7G-��#���XlxVHYEB     400     140�?ߜ�&x����(��cB���zN~0}·�jo��Y$k60n��+:�3^��>���F���b����Y���JK�`"폭�yP��C|�b2 ���<��|x	\.;��(;�s
a�3v%	lM���_%@3�'|?x����3T�o�����_��"�����$ślf6уFv���J��iU���-�{��	�gjJ_#L7�n��Ϩ����0e�2�:�qv^�!�yP�rGG�ʎ�Lb�~�MJ�믌��]��#c1`����d�z`l�@�py�˰�Y�\|o�RHv�幦,8�M�}Ujm�ǚ'��
�#<��XlxVHYEB     400     130J{��}�.����㨏��A'jB��w��;ю+��s�{_�CCqU���d
�.UG\�\v�޲����Ӈ�aO|����+��p����DL�Α���7u�L�>���YvL�V2���O�:����ņ�Ҹ��.e镅������=p�_r�NW[��=��M�R=��gwX&a*q�=gE�o���li����b5v��S?�Ӯ�p/{��\0���82���Ys���~���
z�����$��aO]z�)B�%�r4�䍻�Gf��~�/dk)�bO���P��H����4~A��wXlxVHYEB     400     120�$�i�.�,�nR_U�'�_.}J����#Se�,Q�­q��hW��`/�]�p9�
Z���h�������S�h�+�R��˹yG��S��f�a�ޞ�"�O��m��X(E7"�1��$��m(*�J��=�����@*�'��.���a����KF5)L��dz(^�|$j��%O9�KP�(�a
��ֺ��NT�"`_��Ry�E�]2��|�\2���C��u	��ս�E�l���S�3����M��(K�o���?��dd�����؉�|>%��c�R9�.XlxVHYEB     400      c0�bH�ɭ�"
p%{��oV���5C�'o^de�K�\kv�fnK4d�Ћ��w4^z0�W��)���+�iŘ��Qe�a`�lu��P�Щnx��� ��Q7���A���m����w�{ʉ��[���=G�n�*Y�����T;�:��{�b����xL (�Is�ˀg�e��a'�s��j`�K�ɸ}}�O�q���XlxVHYEB     400     120R�3dޗP|�Ay)�A%�o���h�;�r�!��dn��98ιm�vH���ǖ��՚�� ۹̼3J6���2m�LJ���� j�kŝ�YoϮ�l���e���8�/�1q�Q��$�."��	�RW�QB�{=p3��1�
�6�A)��hEx�[$^��|��m���,D��y3y(�W`�Dn;��^���ē� 8,����PJ��q����S��ϲ�dj���~4��o�Y^~��*n��g՞��"ZL͗�p�
���Y�yZ=��]�vx��4��[Xy/�p9XlxVHYEB     400     120 ʩ��1��녏^C~���9P3����+��K�;�P��gJN d��ό�!�
׭�!�(���x�-"W�V����x�5��Q��o��:rQ&�E���yH�~�וu=*W��'���uk[�<�ۚ�Y#�v��U���W.�͛�:i�x�8*�z8w��{�n���*��Y�oMS�]���eL@������Csчv�����$�︿�O�R�	�A���b��^$h%ֽ�(um��/��qX�t�<Z�,x|��s��6�~����V1"*��0�靕�XlxVHYEB     400      c0L��m���v����%����,��;'I����i 0���R�}n�$�[UZ)�0��eEXH���%�u�,F�|���Yi͉x�|�ǆ;xm��hE��^�;�����ݐ�N��LI�On�Q���2\|�A�-�h.��[��g�wSߪ]��������&�p{��X����������XlxVHYEB     400     120w�o2,��gr�Z��ck�����Q('i��O���$�uǂ�CO,�ϳ�.��1İ>b���II�o�V�L����ou���h&�˼������f��P��\3}1T�w6�Ek�H}�.H���nfC��t����c�#^KyA��s�ntW��Ld���yG	���nC��ݫ[k����؛	��f���Jp����ܾ1j[jw̞�S82�AO��p���$�??Ĕ�0��2RhW�����s����LqieV��Ɓ��л!�}��+� :H�tR��-�tL�`�v���JXlxVHYEB     400      f0���0���P���%�A�=���ܗ�9�a���R荍���s�̻K�l�� W>X�"��Vr����?���΍����w�I�y�O���~�%���L�ۙ�s-]��?�~�g���*�d�e���q'w���T�9�{l�e �Z}�K.1�����9F�Os�ث��})Q��:W������u"����M��?�6k,�n�?�#itg��}+@ku�4�n 8�4˲")[�XlxVHYEB     400     1107U5�(��)�;�R!>�C��pt�.���V(���y�7�>22l�S�Ox�Mֿ^�h���Q��{Ŏ�����P��?�%�*���aZT̏\��
�q�m&�a-�u[YR�q���3�FYx
�^w{�d�|h��hx��Au��v�`C�s��i&U�;=�T^��2��������c���s�L�%�A	CqY�$xyf��cD
=$���z����	�*M��>5���8�Y{�+zT�#��G��5�@
��#q$xCh�mb��o�#�|XlxVHYEB     400     1207Y�زy!��}�Q��LG9�J�䔫��)|�6h "ä�����WO������JH%[0]r������o����]bܵ�mAD�`������e��E�=�dz�b}EM�8XM�,��x>+�2�j]�ϴk������&|��d�ͣ��)/�R]'g$�b-��T �y�>�=�@�n�;�B�K���� �/p�v}�#-e\+�Q���N��W&�J�S�eS3��H���w�|���&~?��4a@��D���=_ݱ��T�e�=9En��nt�n���C�XlxVHYEB     400     120QGh@<��u��s��BV'Ǻ��:2�=}q��SxP�+����;�]ٹ6>ֱU��к��xO�=��}���*{�M��?$���'���ye�&�FY:/�Bȯ�W�7[X^�v!r)��2%�f�v�q����$��0^�!�
gD�&��^|�(d3��_-�
%���82.�_(K:\\��I��XI)�k(�{�I	�Z�[m�&�p��/��~tw�xGj.6���`�^\�J���"���-�ا�e)� ��E���\P86�?e7�t���1�B��XlxVHYEB     400      f0')ʹ˝����ĭo}$��`GP�83Њ	��u5�IXhks���ҽ
���&��HG��|��Sr[O�Yt����	�6YBB7���-Q���-�b�LÁO��[P`���0����8`� �8slQZ���O�V(o�C�d�� �q������мq����8I*Z��K���̪ې�a�L1f
k �%�б`��-��U�'3bA���@b��l�N��Ƚ�W��9���_XlxVHYEB     400     130����`,'f�OR�9\X��2͚TC� �{�������=��˱�V�ɧLHd��vz܍�T�ֳ���bk�0�i�
t�6�j����TNO,v�܁���^�����*�+dڥB��:�E�F���}�o=��T���J�'���PXɀ��pV0�0�L5��n ��L3*_Y����f�T�A�DSX���:���0~ы��peP�<b5���۴��:��Z�; \J]j'Qk���uX&b/�[d4\�<MD�#f���p`~��<�����v8#	.�+".S��=8�U�;�ƙ����,�T4H$�~�Fٴ�ך�XlxVHYEB     400      f0�tX�z<g�Gk�>U����h�hg gd�ظ�FX�.�Sh�Л�.E��|ua�����D�eA���������~�K��q|����zQ(y��cO�T��A=���2G렧x����вмD���)T�f����p���?pH��z�l�W��J��nY����;`��ڀ+�h��t��[ښZ�i�~�wk<��O��2Ϥ}�b���	�}���u���r�bI�]��XlxVHYEB     400     150M��1���I�3�����1<TZ���PQM^)�4}Lh��Gv�J��W��l55�5�FdF���BvI�NE'ɸ��y���u����4�y�hqh:|����;ώ��:�4L>_�m^� x�)k��:���2��vČkZ����;���GY<��ϗX���MZ順�$��qZ'Rڽ�!L�Am�Ah�h���8�+G��l`3���c�<"�jVB�*y�KWV<S��۩ޡ��uf�"��-6�i+�٦�������4�nͩ���s������7��i����_��qF6R u��`�C ?���.���J�G��ό�׋����:��$��XlxVHYEB     400      c0B܌o0_�o}h�se�rq�4:i4%��HH���6l�L�j����i��yN�ꋠSu8�����wn����kt��1��=����~����p]�|׻nے`uy��Fy�����le@<Gr*��z�;�<���1�)!L>(srr��ڠ�d��%bյ�u�f�tdO�g.)?os�"�u�S�˸fRq.�XlxVHYEB     400     150e���;�Z`ܹ�!��1�>ൃNZ�&Q��es��+8��L_n��&�L�o�`VI�_��)��6v��c���-����$���v5���G�6����fk�81�2z��L��ܻ��B�N¦���|��[X�bj�U��Ձ����8�2�>qcG�+���Q0��w�)�˧�ר7`)�P�`�P��U+�5�g�F]�s1���@$.%�%Q�{� i���"D�΋���"���>@A��l�Ml¼��S,�)S�H�x�ږ�Q����ܵ�\�¡�B3��j�}������έ]�?Qz)2@!������so�B��lٳ�3\!x��XlxVHYEB     400     140�j�-�T7���V�(g�Mnz%�����U��q������L�+N9���G�{֜�d����� ����W���8�0��׶^(�Ң(>4��Q�2�ŕ��E�5���1)��)Y���]]?�m�,�rO��K��t�1�§���
Z����M�͒7?�_H/���Y������hq����*�R�ɂE> !�'�Dʺ%��/�r>��l�uw�&Քf:�&@N���|6���_�ޥ��A{�ȳ������KX1�W�ԙ���H�	i����JI���F
�H,�i(�����G��
���Ė�]Ǣ�f�Y�6�'��1�XlxVHYEB     400     100)W���n�;A{�a��.ǖ�U�Cz��S`=�}G�n�����D�SY@Gq�k�Xא,N-1Sq�QJ�ѱ�O��H�D�->���*�3���<��5��,/�����5ڇI���/RS&��TC�o&b:K�e#���=�*���pF���u��&��;܌j0���"5P�c��.�.$?��2�"��G��S�����o�@���jw����6�I����.���P�Fv��ō_Y���i��)�l�²ru[�XlxVHYEB     400      c0�bnqO��C�Qk9�7o&�}굯�?�>'�����n���g�����j����1���!�oiZ�xT�42ϟ�F���y��\�Si�`7�I���x}O������Z��y]B J뎱�����Bm9�,�bZ�9���^'�y�H�,�^�k�(�x��9d������N�V�LW%���`XlxVHYEB     400     1002���M?���@�����2�4O7�]ȴݲ�^�?�0-S����\=n�#K,p��_d��QG�8������>�6;o�kp�3�M��۪Y8��\�`�� #�u\[?�ݑCn��G��fg�K�?�Q�Q+��ok��������	�	:�W�"a����q�DTm��v���*Fd���Z�e0K��u�!`~�<[�^Z���q�<:5�5D��UwO�@���f�=�/�:�&M�Jt�J3JD���6Ќ�
PXlxVHYEB     400     110d�[t��͆CU��G��̍���C���=7�^���P�Á2�㺻!˅1�T�E��&�Â�LT��ߎ>�wQ��=iN;���Y�A(P[
_	��x�'x����j�pL��¹ǖ �#����X��.C�U~K`kC��C�}�r�?qi�?��8Yvq�=�Ͽ!X�a��.�u��Y��v�}ԃ#�W'"��Z�]�g���;3�g�׽.e���/������È�L��[����8�����f�#���sp>�ίm�5�LM�<�XlxVHYEB     400      a0����Y�GC �ݚv�ed�b���HY�#g�D�;{�Q}>� �VDcJ}Ė�K�ɾ�x��c�˨�U���,���|���#
}��n�>+;�L��MR>ВE��4����<�`\n�u��&:q�s z�B	�
ۃ��b�[�00�Z�B�
�l�0�C�	r�XlxVHYEB     400      e0}����ͧ �y���ì� N��~�A/E6B�at5��qq�0�Km��`g����f�<� Ĺ,A�~{)-i�r�	������D��T��=��M��-O&��A���qj�o�d�ˀ���HuSXf���;�|�xh����'~h�7ЉJ%�\+��fY���!�H�E��j�x7չhY��:�i�M���k�����3ZE#��!})?���u$4���-�XlxVHYEB     400     1a0�e�%��7�� �[1��~�n_/o��~�0w��J��������[m�?u��YS�\z^ecߣ�u�����+�@ԸWL�� �R�b5�Sv6�"�h���1*�B����#�Z t;�Z���[Y�G��L��X5�7+�f请m�Ԓ*G��n�{V��g��o\�����0`�i
G��Xc�X_cZ�鷶�e=��]6�m[��p����0��W~�i2����Pje�T`E�QQ��	0���!k*MO f�Q��Z�%�H�Ҡg�l�r-xz�?fT'��Ј��L��|XK�h|��Y�P���ۣr������6����O���v�r��8�Y`�rR(�/l�a��"��wŽ�>�d2�]=F�8W�.�W׭f'�EX̡�[D����sjѽ�B�z�`�(t�ɢ�Bj攚pY�PXlxVHYEB     400     150����b���r�&��1�87�G׽O�ZS21��wC|�LZ삇��|�g����yt��QV��aQ
n��'�w�Q�v�����.�I�[�j/w���W!E�j����� ��z!�t=PFlQ��B��-���[�Y-N�h�?��ŕ��\�dט�q�%L��� ��_�D�}�]QUGA�GD�0E�1����!h����i3>ɸ�&w/�~�ny�����l�H��M(svL����{v�;�8����s7�X�mS(��Q���6`�v�<UJNC�f*�����a�#҈��P�M)�jg)$�be�`t���\�e��Ҥ���B��XlxVHYEB     400     120�E��F��b��*�H|,- ��-��ô%Œ)��WG�;"�z�M���@=��_�z�-���e�^��2�2��l�"�)�"��F�.�0����bPo�Xa֧
f�<����ֻ�\r�ʡ1u�0�p����Ƌ��k-�+�9��d���(:��(��`���H�2C��@��F�A�&`���O}�E���K���ǩ���gS��9Bу�iy[P�����ޠ�Qa{��Ր�j<%�ËJ+��YH,f��X��ID&�L�lȊ���l���i-G��!Q�rI���XlxVHYEB     400     1d0M���lB�w���~���/�����L�N�`��>z$�QX�W�G`̖��VLe˕���if
㾹[��A�9��;2�'UV#�����.E��a՛`ج�h�\]��C�"�A��գ��NK1�3�D������ �@o����_�[���e>�\�����s��J��V0aZ�����>��j@IS����A
�g����+b��<�;)3lE//m�J-A.�b�I8H.=(������7�����V|a��y��JhtyE�Z7����w�<���{�u�h���q�B؂}�M�����8b�~�O|n@�#XU��:�^i�)�	�pJ�%�᪦`��[ݢ�O�M��:`��:��.�g#|}� ���ͺ�t9e�PE��BT��`T�g@��4%�r ����G˽����D��1�u���L���x���j�Lz����\��+XlxVHYEB     400     120�M��,&�zR� r�I2fS�������K����Ox�������!�H-�~.�` /�Y��T�;銿��(��P���h�Oz��	��+l��/��<�yX ��Iuԑy
¬��v^���v�r�L����:VP���̊%'vO,����lQ��w���
�k��Ĩp���	(HAS��4A�ů�_>�X��d�I�M9z��e�L��q �{��_j����{�s*qi͠�ڭ�%y���д��TX��\KM��I����hR���p�e5�#tf�3c<�"�i(�XlxVHYEB     400     100R����G|����m��t������01D��{9e��gUzv�׌�f%���y�c#�e;>{sr0���34,6>l�6����������`Cp���'�dy�.e���R.�d��&lF���^��(}�`c��FM�CiF��^Ga�V�܌g�a���c)���0�J���@/�,-�1�V���?af���K�܊��('���<�1�c�%f��]θc��K��$UyuO�m�.�ӡtQ�y�R9?���Y�XlxVHYEB     400     110��J�Y#7K1�z�c�_�����طYv�7>Ga}A��p�TW�:#=?\)�=��$M@nԦl�>�����/!6D���B���:]���4���ej��d;�:c0��T��vq�6�pw��u�p�|nb���iN�4k�m37���"'�If	�'Z� ]��_�S��l�'�c�N���j)ū˓��4�^ MU���և	o�<�r�ȓ-�%h�����e��T��G�aPM	�@eW�x%�Y�80�}G8�5S_�Wj��u�����r[w��?Z�#XlxVHYEB     400      d0q���.Y���'��^����:O������T�.�f|��	��[�3~A=Dr���ʜ['F�DS�"��k�����{�:�����5an���#|82{���/��n���U{��s����j�s���7�f��A�C��EK���ë#e�ⲻ��j��e�؊���97��F��
�Y�W�@���u�=�Z�O�b�֥dY /�XlxVHYEB     400     100 +��it��]@
$���v�\�J^}���.�KI`���=4�D�8����s=Tt�-1��TS����Y��ԂƬhq�Tu��<�^	�
����A�
)�h�Xi��ҵ�}$�D�Tw�0�ۻ1���q��@�s�i���&����{tX�*_�"B���5ʃ�Ĳ(�T�� � �7��ґa�ѡ��RWC�V��V"�ڳhn�PN0����ĺ�3��E���uD^�iפo] �r?Z�U�.a9XlxVHYEB     400     130�e�ֱ��16��M;��-�j�]*@s�am�DA3���%cV.�x���|P�gl���h��̈́4Ԭ�M.�ܬ���;� �8�#3)�פּ[����e�^�{�~����^#(��hF������Ì� �`�8�V{��@�
����ܽo؋����2oJ,)ԛ�t�R�I���2�.�JO���D���OQ)&�b�C�A��|���Pi��-�� ������5���J���ΈK��C������M5�ev���w�[,U��+v�Z�r	_"5.ޒ��I:�yO��x�QJi���XlxVHYEB     400     120�H�� �hH�����t|�Z��~�=����y�����662�����H��XfS"�<�ൿf��ᅥD�8#����~��ƪ�6��B5���tuC'���"qid�%d��_�C��I^��Yϖ�l�W�*b��g�>��zi�L_	�ҧ�:�t���p!5A=��_*��F���mt��zh�(9������S���V��R�w�בEuj���X'q���_c�&��s��P����-�i��t�3o������qq5�dkS�I!>{X[��i̝����9���XlxVHYEB     400     150����(�U�[���tL���V��=�ݵ�l6fϔn�eŧ��]�=kf��ɶ,D�	0,�E�$��H<�{7��0ۯFlM�-�:l_H��������:-�f�#􁐹k "&~�@����oFD�8�>]wH��OԽ�;;�v�g�95ws�xܓ��d~'4�lj�R��9c���qh�>!Tr��`�;���a�ן����5�;Ҹ
hc���+m}�O(Ȅf_7ʰ I�YsU�ӤF���*�g�R�m[ߠ�UhX���)����=���nņ5o$�ֱ�<�?ױ_��4�K�o�t�X��� �Zl�㮞?�~Z&���XlxVHYEB     400     110�bS����t�s�L��$%k�8h�Oj>[j֪�> ȯ���N��oѡ���������6_[��'��'���7F;00��X���!�CB�8O=t�-Q����X6z�"�J�'*��,��O��$Ix\%��������'oZ
�L�a��¦�����mR�8��=����ެCUǪ�L����?�e"Ɇ�)�F*4�:��G�uw���åf�r�g��Hcb@��Z��2��~ _-pތp�n�pۤ.#�5������Cq�}7XlxVHYEB     400     110���RR6^45�!	�2�B� �8-�:V^*��ֈOX�4���6�{P�z���֙�_OS�D]�4��.m�WBK{2�\�ɤ�;���2s�9MB��?������*�����@���⠙\tD��T���g�����2�L�\�5u}p�DA��B+���X�(��=2|����w��;M(�]ԩ�
�g�ZI������zЇ)��0��]T�g��D�����K5O�t'��<�D?ב�!Rs%�s\�z��������Z��*aXlxVHYEB     400     120���=��`:���E�m|qoZ���\�5ß�h�	��8�(�*��k�\��8s�6ը�Kg���j��LI���R�J��G�#�y��7�(Gu�E44�C1��\�!%����Wn�0w�Rq�x8T���5x4f�h Huk]1�u�i��2�p>���d�涼��t��{,l�UxY���7�D��LI`5x��b 	*�W�?��N��Xd}/��o5�z����G�c
���Q��v�̞p�u"�M
U�ּ����t�Q2Ƈ������<!�]$��	�bnpXlxVHYEB     400     100-� u�z2�	�kp=��7
�&�4k���
�K\�%r��*�HZv�A�ݤ%�;yHxF���΢H-��o!Pt��������i׷�e����W��h僺��X�sw�����q���{���Y� �Έ6��1�[5��-�[s>#A���[����6U��N&Kh�����P��V/���yj,]��3�s;��U9A$��F���SZY �����i8��׾F�2��:u׸RU��|A�Ƕ�O=�8ф��XlxVHYEB     400      f0Z��5͚��;��Y�=e%����1����[I�=�6���P�8��y�"��2��+u��AI��Nhf3����誮����|�q�0Ͷ���!zH5��v�")N���&.n��� }+�h�ˉ���ճ�B���4����s�jp%2坪�)a$�ը�lGQ�͇������|�B=?5����.'��_�+,c�^Btb��0<�Yy1>G�\��@�v�G��=��l6̅E�b�XlxVHYEB     400     120�|S�ue���Y���/Q���ٮ(�Y�
p���"x?Ұ����j��ˆ�N����kq�i��7��һ"<�©V�Q�v�E�L�~S�Ֆ�	�FkMbz|��QL�0��v���ӫ|6���Eg��hZ�0=����U�C�l�O�Փ)ֺ��eZ7 ��\��N��X'bD&�T��_�M#�^Do�Y�s��;x.lRX��T�'q������g|<KA$�W�)R��N:�9��=�*�φxi���=��c7���Չ7Zm*��+�I��P
!�0|p� ^�^j3�qXlxVHYEB     400     110�y�qC��
>g����Y�uzʌ�h��{�;�x��`f�S��ۍl��d��(o:�n'Y���ի6��f���\'�R�i��疩&j�~}�ڒ���p�>�4��/'��5��8�B�O�P��I����L���!�}��Z�<C���Z�=�L��@+4��\�1�����ԫ�q�rn�)�t�2��o�}5��g�+doA[B?�[r���K �Lο�(��$I����s�+�b�-"�s����/�<\��%}7&��i�5]���a�YߡXlxVHYEB     400     120$:G5�#%|���0�s51@	������3�B���������s&hE�?�_<�� 6�ۺ��s4���9����L�Ǫ�Þ;qc�V ��ab��*�X�^���in�j���R`V��O#�ń�n���{��p&F9&��QQ��M �&RN��H�7�����IWD��Qq����������4�1�&,�ɒ`�Sl�y���%P��Ԡta�r;�P��3�P�i�W���,��O�i��ϳoW�RT2	4�D��l��k+��I��i��ms��a��#�LXlxVHYEB     400     140����.JL��/�n#&}M���
P��k�h� iZmK���{ږSZ&�6d�=.0�GvF��_�	�۱��d7l�k���˕�%=9����d� /wT�$j�^vO�t|����(񓀿�pN�ۚ˿{�$���	�n�k �?3�@I��nRHf��.�J�즈
9�����|.qH�Q.�v����3O��G��*�L���p�8��o��܌��<wPlW��)|5gaUG��'S;K 1��|�=��vt��ެ�(˼BW_�X��g3�37���3�1��ޫ\���&��p�Q�g���%&dDM��V����/XlxVHYEB     400     140��U��N�����S�L�aQ���Z]��i,���	"�Yq����
]>T/�*2+���F$M��2@�ag���FV�����R|�*�AR� ��+sLgTYDhӜPr~%|�/�M���m �cub�����G�Oj	l�����M�gF\�꺗GX�'	K�ъ׫/+����t�۞D5��鯿eHC=�Ug��j�5�U<*��������D3iT�i�d��k��>P��(dd�}��/E����~;B��e��ۿ��E%�,q�����e����>�m���{zXJ���fWͳn��fy�pM#cozm���XlxVHYEB     400      e0ޤ$�&���0�����鼓Onj�x8�1ybmx�J9�J_݄���I�۹����W^ A�d� 0���6)����{ި�j8e+
�N��������j�V�CF|u���u��۬烨�֭{˺C�svY�Is���j��TD�H��k2ƒ]��V�2&`�St��|'��i�~�Mc��/s���n�v��L�&]"<��_<y�U$�'}KE��XlxVHYEB     400     140	����\����(����� ��P5�!*{U�V��j��������[4_��W��g��Li	Ohb\�2�i[��?�.p��\�~fN��ڬ\o[+6�1�B�dy�q%���6ް,NWC��l�8j�&�U���~A,��x>\�|�$7��s�JVy�>�t��j|I"���$�f��x��Z����4���VI�Ѷ�6�#�PG�O&2��*��HD�42�ҳ"����h*x~��24xӝ�f��XA����a����A�3Kϴt�Z�'�������w�Zwc ��ӎ-�5��n��vV�$�Ü�N��XlxVHYEB     400      e0:m���}�rRm/� ��#��)���n�lb��z���p|�å�ݚG��~&�o[MV]˃%�-�F��΀�Q2�Pa��K��N>�ѧ�'���Q�����ȍ�qwN��헮���½D�3�w�d�lC��� 2���:�(pgzv�4rtz(s�d��� n(�e:Ӛ6�oA�Z����)�"i��b�#T^^&?R6���b�$�Tk��`��6_�N�XlxVHYEB     400     190�o\�Ѵ��-W�V�v4o'�[o��"{���O���@���ǣ������;ݤ��o��ζ) �
�"U^������1N��/�]��-�Ua�;�b<D��=��5��2���j���r�}�<�8d������8��{2S��A���{ܤ8����_/���G�BU
�x]�S��������� 3��%ߝ~e!{��-�yr����V 2����cv^��U2a���vN���ԙW>�3lm�7$��b��BI!��$(@�A�sAtp�<Ku��s���c���IO�`�1�|�E(��1rO��I�J��R��%�2��Qs��x��N-϶���lۓŜ�40�mFMi3V�{d� �s�',�k@�z�K�����/"�92�0�XlxVHYEB     400      f0���t��Y}��oEni�B����
,ș(V�n��w���>� u������Y���Ů�����AP1��W�X�Jص���U�$�N�����(v��C� �V1�t�@ޟ@�u�ޙC��B��T(�58�<Z.�E����
���z���#����.��щm�)�N<�_����n)�2~�U��.�_�x@m�M��k�S�.#��1�.��uʍ:�=��I�2�J��Tf�lD���Ei�����XlxVHYEB     400     120�-��U�ڶN:+#%�����\��ė����lp���t[��'?��:6دx�)�;���'Ne��%�SI�3C5.��8�Å����N�t�����W�Sw�Ckʼ��e��*ُM�;���c�'�H�h-7�&��R
�XV=� ��Z:@�������i+#m��UT��!N`��������
������]�o��S�KI�'��nq�P8���C��sj��t����D�m�ZZ�#�� ���sB�睴E���ξ�d�U�׍V^H�cj�k*���h��T�sXlxVHYEB     400      d04~ݨ�i��,&�mp�7l��j����R`��b�z"yŶah8>��@'2;���(�4uPo��2�>��p>W(o�֨��IX�Pz��1�ku�bɓ�藱|���廿�r���'P{!7�ܘ��m��.Q�� ��p�)nq������A�~���]Xש�p�@�E�#�U�	��B1C�)�@�	1_��0�,��Rl��ӘC)�b)��r�XlxVHYEB     400     150���}�*
Q�q���8@���4Uk���_Η堎���?�� T��]�7?K8|w�]�'lD��C��DԥcKt���E�}&�� �Zt|:��R���)�S;�ڪ�Nf�_��1�~�W�-��(u��afJ罙���mҘH�;��<�Jp��Q��O-�pP��X*�5Yc�|MVs�s_^��&��@M����j��$mn֡	/Z������I��B6s��r�9�פ���W�Q�9/�&z�%���T`���$�f�nF=Ojpʰk��C4�6ۈ0���*i�}�N�I���c�e�FѺ�@�W"�v�[IlО�-TZ�XlxVHYEB     400     180Z�_�]��ו�繯+�a5	2Q\p9̇j� �� L]g��A���|�6!g��8�I�f�k.����F��7"|��(P�.v�v/�*(�a^w�y�_�_^��)�JW�}w���p酵	�9[ɝZ��9��#���>��S(р�1�Z}��Bՙ����OJ\�v��q�/6�B@s���*�#�`�����#oM����d#V�r��a����/#�1�]B��R-����p�װ�'ʶ�e
�6��h��\>,�� ֛�.�/*��ĵ��/z��\k��2�=ͣ3�i���rxD=q�� ,%%���z ��9�а�(�q�X<k ��bb
��H��o���ڵ���MR.�N��ĳϞwy���:��rb̻o�XlxVHYEB     400     120_�K��?U1�E��&
��B+oo����!@)m�n��~���]��t����uIj��·Z�&�8b�H�o�W�E���	iؠ	���GM�k�26��a��RN6��X%fg�$ƨ�g<�����x�1n�-"� y�J"��S�z�c�m-.#��^J:���μ�R�7rE�M���я 3�n�^j��k��7�^Y�
�ه�֝S��B�3�`�U]�^"c��\��.�mr�:�ն��߼�>93+����s�윸�%Z���νx�m˷�%_� �6ŸXlxVHYEB     400     180��a�f��K@�[��~�yݐ��=!�@ �ձ�g�J���@-��K�[J�c�z�N i���t3�yޢ^N�Kf ��X�*n��5������oރGO�b����q��;�p'�~)'w�CqB�k#4Ӽ�kTŇ����6^<;c
����{kL�j�zq3Z�)�Z�%����B\}$pJ��cgM�[4�Vֹd��?���?32�u)��^�P,�,�BJH�q�2f���ԛo���Kݣ�{8�������~���{�|_�@F /P���O"��z�g4�3�:�
}iz�3���>�{�-��ʆ�P�~����g������I�mL
�����;�M���J&��ؕ��X1��6dO8�`��ل{����F^Lw��XlxVHYEB     400     120p�z~$8+�s:����n#y_8PU`gߢ�@�Gv:��:B���$A���5�2��73!uY-���" �-	�Fz�Q�š�95܆hsX�j"�}�l�ى7�5�AS�޼L��ö��t��dז��%*�vs�4�K`ɔ�t�:/�ǜPR�u�y��?��^J��͛&�0"�Q4B����q�ƃ�}�Q���>�{������;M��s)����O�Oȕ"�H'���U���)*R6L��������1�P(}�x&�H�1>v�Z���#(�{�A�r��z8��/�XlxVHYEB     400      f0Ͳ���H���ueGNPl�v8���{�W$���B�vj��	e�?��?�_$�	H��
���&Ds�����N]��&s�R����K�4&!D#�<���}fD�;��(�n �]"���=��
m)�@Lě��A%��{6�Q�/W�}�\��70}�`CaZ����5�XVB3y��*ݛ�.����\[��t��&��\��g�E���8�0q�ؤA��ۓ�n�활i̕�2_XlxVHYEB     400     130	��_ưDK�(�Z�RBM��-jN�/ˌY��)�
R[���m����%�h����Ҵ0|J��'�Pzq�.>;����G[(!�Mi>˺(TG�v�u���o�Q_uxL����k�h(�ŷ��>����16�t���@�G�1�D�� �B������@S#1d�1�<9͜:��~�ݶeY�����K�"8��ɿ�è���s�I�,Py8�'��hh�w$��a��}P��*m������j]����l{:�oAV�S.��� A��::3$�[�p��N���A���XlxVHYEB     400     140��k��B�7��ɕК+����h�`��^F��!�x�r3�V,�S�rI�`F@	�p{���g�~͢M�1�bMB+T�	���*\u;��z�6yl���罭�ﬆ�1�b�ѥ���`m�@���5?��S�b������}r|s{Hɐ4�aZ݁[�v^~&��_ˀ�%�h{n.}��OП�g��ge�4��9Q�R��V}A`�ef��$K��8�ߦ<@+�W���y��D��fg�=���]#k�rm.s�es��.;��=�+���+Z8]l�?��Q�^X�G��}�wlR����5~��MA:��.�r�c��4�`E���یRtz_���R��<�=XlxVHYEB     400     1401�!���r�}_jy=�qd���u��SCO˱Z�[-��v�A��{PmРP�PY5���hW�ROU3���F_��rw�et}�Q0�R!÷�h�}���Б
�!ftW~��#���y-���7ctpY֛?e�|��I�Eg�W&�q"��h�٢����ET��0?g~M�M;h"�aIoxO�4<�hq��������|_�]"��j ۼ*���=����WϬ @�B���#���4�MGxo�u�aYԺ�������.{�&-����4Їw3��{���4$�q��|���ao�&�k��l&��I�j�	�ź��
XlxVHYEB     400      f0Y�¯rÃ���YP���mq����:׶�q��q^^3w{5���[hT[��@�Dg9y��?`�B�=���|�����6�S��.vv�'+���cw̜ZA� V���x��ϯkh{v�R��
T�Z8#u�L����#�)�b�������?�=�F�1��wZݭ�.���H�V��-�ͺjd���UX�Z��(e�NϨ�����i Qq��]n,=�(�B��n~J C�k �`�攐��c���XlxVHYEB     400     140D��rgF�b=��/����5:��({���{���|f��#ao8c	����F?�2 և��v��_&�+���U��6�&��I����KJ�;'�G�#�p��{�%���^c�VT���� ��x�2���êJ��$�<	�X`���'-�f���w{o��UsV����8J
 �<�����g�cF����g� 8퀠�Ȼ?�X�����y�i2���4�T��3�41	،!p~�֕>ɦɝ�k�{����`ozҫ��6@���ԭ�g<�]��Îݺ�BIEz��l�d��$	{i�Ф���z�j�Zjem4,9^�@XlxVHYEB     400     120dBQ�U�(�n;�҇��ţ������aud)#$I�M�`���x�M���z����dE}Y�z�V:G�b^d�4��Ք)"�����2���z�����������u ��<��7)�������
@7�5���B������Ea:��@�?՜ߐ�ey�d�� 5�qWm��w�h��<y.���^/\27�t���jo8�A59�g�X]׾t�M6"�@���*�Z���������xX���+?�#�Or��c-��f<��:d�#�T�!zn����XlxVHYEB     400     120A*�#{?֥�Ջ���������?K�:"�����W�Vr8X2^�w�/6�˰��[����o��D���S8����C�Τj6M\�H݌�8(Q���t��s�L�-�z�#4*�mm�5u~d�ݼa���7�kJ��o'F}!Y�ѩG
gƖ�r�]+�M�gw�n	��Z��>S\(����%L^�Є�)u{�g�氒�����.U�&û
1�/Ac�;5��N�($<��3�N*	�O�w9	k!��u@�o� ���{��#Ϡ�[�o菕�(��XlxVHYEB     400     110��U��N�x�"����-y���Rh�� ��c6-�����`�ţ�S�i����Y�`�6�8�.u
����Vh|��T�5����Xk�g�N�1�-��A\
��7��H�Ps�����6Xu%k	�8��XU�7�����ǲ����6�j�#�Dܲ�;��KȻ�z��yvn��w�k
�^z�lh��"XH�V���[f�s?���[��U�����5��
s��^�UH~�1�����ì�ɞ9�N��䔶�'���?2���XlxVHYEB     400     1600ϛ�MN�H� Gg� ��d��u�Ls�����w�|6�R0���$ٷ�Պ��m�#����[m�}�vb
�翲�&C��g�^��x7D�N�8����o��=�T� ]���#��}l��ܦ^-�L<�2���gRw���Ŧ��&��F�ެ)�Z��-b�N��r������c{��7@���O�3f�N��;�@��m�pJ�	*�W���
2�7v�DX���� D ����� 7�&5eu�-[Ǧ������|Q�rR�Ņ�3�0Nu���������kuX�C&ۿ������uk�Ϗ��o�[�!z��v;�+D/TXF���XlxVHYEB     400     130�"�>��W��X�ο��<F��fU���M�ܺ��td%�J�}����Z�Z�;𱋕���\����lLXM��ӿ��E���D=��vؒ�{���Q�2��kD�,v�TE�&-T"�74��Sͻ�R@zG�'~ �����b�Qp+�T��q�jњq�Ng%�za�\4y{��l���H�������)~��$��f����χ�c���=b$�$����W<����^�F�aN����pK�L��Α��精s���M�ʱ1����_4}���v�3+t��g����XlxVHYEB     400      c0=�2y쫴�u�?&�=߬e�E�b�M��&��-rk��دX�"��M{�P(�I*w�hJ� �kwʝkU���㥖A Y�k���|0�tU�D,O�����q(Ն>��Ɓ��V�=�j���x���4)���6z��N�S��C�}�Z�T�A�m����*�UyYC��Bv3�X;�^x7�XlxVHYEB     400     140���O�7bI9Uq�C�2ԍ�Or �x�������Qm������,$^�o�H��_Qs(��ȡ�-���?� ۍHۥPeo��>��lD�
�= jl����/e��V��7���K��UG��焍��i~t��R�{�8��o�o�]�=�Ϗ(%Q����#Έ��4N�0[�8��ƨ|�v=Q��qd�f�ި��NF���c�ǫ._+hs�H]E��Y~�L-K�5j��F|Q?�Px��}n�w7|�l��c1A��:�Δ6By��z�;��`��K�ȗb�&�Yrx��?�לI.���XlxVHYEB     338     100s�9Τ���̮�]k��f���K�����fJ,�s+JYY�:Bʇ�ڇ+}�<'�# i��Vaç�6��.�i`�����x3R���#��9�o�����
o޹�
B}�j��RλN�K��7N����(i$��ĉ�X%8����uqa����SmU[��)̸�i�b�����0�ߔإye��=/�[�zyH��������s����TLo_MU�=��{�'{�բ��F�F�&'-V����U��X-