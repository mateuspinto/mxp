`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
AMPLj3Pq9ubfuir3ejXADUs8xnt63ynbIrmvs28aHM/DbYo3D37krYsWhwODnuoVb7DyxWRL6OV2
xxbCLxdzdtBb0LZ9mxPMfsZ3qt+Iktv8i6F+VHUC+fSyKTyKvVoa7pNlDEvraJwRtu5rM5GkJ8s1
m4k/b0vE0ifOtOqxCRiJa+SQfPvoN2UGK5cQxDozRw/iOnqzjME0lXqGT4NevhcE6PXeNHfYPzaI
c9mWNwjsiIxT8oKmEUSnRyl//Dzhg+F5LBS+F1HIKYaG23OUs6EqVUg29AL5XSIALGOlf3WxS17E
22rwrFMEQ5ivBgoxqi8aStwCIK7fOHUVDW3exA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="k8kdmIFRUDlgraqF7Sm204pC5WuSt6xWBaUySwrTGAc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6528)
`protect data_block
Ztcrm2tPFqsvHrvQGwqnhikofCuLLfXRJHMP40La+eBh0Eps1K2V7AySXxm8QKNXypN73G3WDaZH
5U8FAAEfZXKooIB11260cgBSe0CuM9p/09rS8m4vpKVz4dC++pyrToFwpWtViR76Dg17mGbiJbLq
cy7JKu4pCVxsS9wXwd7Xbgj4w0HF4mDYztcbPotw1JDjjbjoLmQCWrrDOC44OKKts0ObGnGKs2y1
wDSrhkBSknM1wx3ZhYD+pwm0RvlGv4YBjiriaUzSoSK3zFto53pPEXzdRRC0N2FAW0plzRqIEsYx
jENpLdw/zIdt+2v+DDDz0HlBSBlj8fnHz5ZcDcK/K5dUBebUUF6mUgUjSx+7n7itvgJ3pbqriL1U
AeHVc119ykgDtV3w7ASKckNHkuitTSRlypKS64xAqRl/1NrhdHO50DnfrUMxbTNqPMpJl5tS9rcM
BTQW4PeQAz3rO/dlwyfd/dG7C4dLw+Y+EVbcvlt5z7D57Le1/we1VpRNvufnzdhXS0Is3P+Irdmv
0Wnxj30I0pqPPUKHLkf28kHgZ6crb6h+ov/vsyys5c6BJxbpov4Fhh3CLzUh9UlyZK6R1zX44v5Q
+yvPTWEVXad9GQYYBs40JDHAXbxJsI+5nskngeDqDFeHERFywm/VoX1ACaJa/bQGyX6+hHso28Fk
T6RbfMEJkmSy7bJjD04vHJuZPB1PcWayOrG/kMnDObcGHlU1WGnKKSuIEZa5crPl+cM65zuyUF9H
cNFBE8NZZ1/dIFg9D7IaCy5GT/VVlEjrepm4KoRr57APiBVmGLWJGPtyBLemzXyUVSDs6gpb9W1b
QNOvUX5YEMeoigd8HpJbuzlAAzz/TAsffG5P49VMZVsJIyedbJIZ9uA395hHzs2lXdpTE+8pLIlE
fumnXRikzEit23npASlM/6EE9OuyTw/IFSQpDtfImKExTohtjZJ4crrgCWibUSUyksCo7TVQRSyc
8Qz+36XmfkBU5DFGR3lSw6QM4tTpu937+Mcj7z4FPAOoI7C6ftxL6Bjo2vvLL9NzVAyPo+puRDNC
kjC3Mba5/ESbCHq2d7pdDoQV6F21YKeTCPJT+inagGLltWeVo9h0niHWTJQfEzZtaNgOTp1S7W3U
kOuYyqBrrF6ghLSM0QtR2tAOZV4S88f7Tc3oQhNczdO+Ko4vSwh5RBrnWID4iJRRZPds86t91OW+
8PWx5Ek6/9rdUKjkfv7fL4yutRFv6/yH+zHUlSzdFOq/MCLCyipLMkpBHjk9PqL/8PTagZGHq/8y
dtQiMPoE9845tGvPG7V2iw4igLvizhe2+XVSA+YgeSAl5EfgbSJey5QeLQYlS3Zy0j3bW+QShk6C
fDH1GNu+jiV7Jbm5ZOkEVkpzJDq+f/zv7I4gujXSfA8OKXwbrnh6ZV2dQL0kQ/4VqPelfLGI8OpP
baUydlVwhVTymHJ1UETlf0PzTFLQInLfEWEuGjm/s8+P2wPVPLp9lo1pT8IVFI59kZFZ4BGyRTiO
PH5cp9KtZu/JyoSSMkknhp5BErc98mV9hd7v2LSI9QtB2Q7dn/0A4DCSCDMwgkDna4eWehNQrI5A
Kqvc9okA/u9HIJbxsDeCoBL6iInT1JXljbkrWnjt7PEtxpiMiLM0c1PI2yvm1+Q1fid0TdYMOL4v
r4DnqsnWSAP4Iq7TeUKwwLLBA3DNjutR0YXPwSQtBUSBMduR9Rfi46MmtDHkptPI1LWdzPyrltnH
Z5ucEkZtwqlqNWjaC/PqYEl0Fw3PMLV8JzQevCxknbB7T2v3ZcclmzkUTx8zH3TuXhXKLV7UJqaq
oyaGbyKAFh6Oe1UcF4BTX8WUZ1RSDrUl/FIKkDLvEJjTp9JkBJfgZa2nkizArJXhya4ogwFqVt5C
wYcCfWiB2Bfb+MAzXzxAKX5NfaezNy4Cj0OrYtEv7EwgDlMNcsakzn5p319eUIE7bg1cvllW3beN
kaZXQI5DUJMdg6IepkvuhRDAPWrZIR2Gey58pxkh1VJl0GpIM68uZngKMs+nUBX+PLXl4Objo1qM
hARvu4K+HEf9pZKg3JDbf3VigIb3TrvqyO6tl9YbA1lBCRjNeLJPog5zU3BLzjZNAg2/Vwsus3gl
WHkbeJkjL1pp97T4gbcFcbYwVBqFoR3cNQk64d/J3J8xipUiFO2YUrkCAhyMfMnTt+AjXFT7JLpG
Fsj9Yzyn5nqpB0GU4R2zy6GJwebZO1uhf9M/xoEu2iISqaUZkyCoaQoJD8FBn1aaPBwohVCGGUqe
3wV26/AvmN9c+a2P4HfvD3EqMcOqNWoO10Azg6xQpYoMA8e6oSpkm8poP5QPalusvOii558xQPkP
sFtwsjsEYBQHDiZJFcJXuw5b1a5zK7DRDwQ2RD/bPgk7mN9XVoqn1wqXRg8MtCbO0uor2Nx0Oroc
BA/AHTXhGIdTaxbZ+Rh3Xpp7Rx6SzT3s92HpJFzp2nZnUw38n+nNdMrnyMU4g0Lyx6bogMp0vGDa
zMDspNygTstNAwzWqd8geGMazGH1Og1t6VrCYppNirir0yJI4Xo1NgtyXcY8H5kd5Z7sID00ogvI
C+BVJzQsFDKMl0ZwtVUhFwW3DWHhZ4quJjd4arXStU0VjA+C7mWUze69ShOiVadhHis5o8wf/AmE
DW40C6wJLzcED0ww5ncoLAjQHkHF0/mc8CYKelQtjnfv6rvDsVXkCJ4wvlgWohkjbhg9hQxZxiql
RG+x6Z17iJ/sjl2NPrTn48mM9lZdpGlzbShouKcFhcw4EwJGowXrnbEQBJHo1TWZzqnLe8pHT1O9
aY+txUjIlYcV+VW3rG+MjPxoMM4aiP7EYIf6kEbvyqIDdT88nrccuNrP1YEhsWmfk1WT5jJujp7z
a5aWujxmA8pnIREx0VrfkJ7bb2WG1HRIDWaWGWTgVWdvadNGruMkurdACvsBzHSsuUaf+AhXDVz4
U2AYbnlHuMKV5xqCNQEZAymNk/VUKw+PF02sDwbAQH/eB0MB4eIgu/Rq1TMcaU6IPVaXCy5XRBVt
JEX3VhIzgbCnTFGOD29D+mL6ywsDDlq5OyhBhiPS2gZ99gekZC490K5DpB4Qn9Eiju/P2vNHoblB
TQGt8vRSaWQDHeWUnH+n/t+7VZjwsY70I/H9mcuurDYeCLN3X3Lc9dOiIOr2faqAqRPTDtvZMuuF
ghPo/wqXVuxt+DHYEJiveEE8P3LPLCgn53acaO9DGw32VS+VZli6QsF2DUcl3dU1mEhoLhDSwIEK
2AM+MLJl7Ly8wP+o6NbLP3nle+kGjiwXsbjQmjwhld4HeblYbrbkvN4pnRvNsneB4eqXrwfKVkmI
t7dNLh3jxxDbr2mHHN5Smg3l+Kc+ubnxNCak/GoQSBe96yvm3ztG6CzzqHqTza14EZtE098DEWa5
IdbIeZcZssRZTiAasoxVf2PnoKbqWJoWdHU3Trbvs6OmsxWQbTBwtG4ZoM/LctaBuhh3yqpt6pHV
j4MCYa5bVy3NJuKSMmefw6KcZw99zQPxhUqCG/eg+W/gmy9aEiB37mYidkH1fg6IE5b/XRnOudQD
9OwSgqjyJ/AgSEI/thbirpSj4Sy46Q2mRIjLqD9wWk23IcRLHsWVZ17gNRVNsPV2e4vU5X9yIAEj
uJ/eiU2fCHT8jyh4UwnXJsd4sVhYmTQJL3drSZ+yXpXHnxuzNSX3XDBq2xpXJXNjoFzT0lBEYDR8
4bUHt4G2QEjQP+ZFflX5IJFqodtVhUfNYrBQeMGiB58LvfAxLuuN9pLYNAqttigBqmNg1NQVvVP4
oYnBtCiKHQIWH3VKKRdk4MDobJ3mdCS20hc9dMYGswzUB/DQYk3eX0xZc12lTrGmpi+V8JGZxk84
q/h+PtNve/Gl8IJFp/3EZ+seaGhMvySo8A4ICiRYgJi1lA55htUrZ8t+7cvU+QfDOHOPGbBZJ2QJ
oP15y7jLV/MUzUGGQeY7v0YUGAYUOti7W0E7rZl6QT1fWEe58cv8+tYoIqJmByD1JNHxqm/WzoVI
t0jucHXQuPdfnFXA7jSY+zuPBCKWUl+SHN8818twWIywGeNURhQWEd94wA2VVfBGg9st7Z7KQzr2
FnnKIChd5cEcvfxVkOwmc5GTNRf9fppe9/4zBfwBFcNOc+x8om0UHE+XpqFLXRG/BxMbHROa8Kow
U7yZe18sUixXPfxfUtNvypWR+6hi5o0vlQWoi4+XZsuvUSWakq+HtwqxCDG9P3tT2f5bkxlMGPF7
Lqd+PI3AO1tZW4CqI47+8YAWhlZ5BbdNIqijmXelhvWZ/gxNA7/Z5RdfRUzFKeONb9LgIgjzqnEC
5VezO4h/9jjiUl9Aj4Z5dvuslepDfrW1WIGdNe56j6v/gflXCaKBvUHhDXU0fOta4w1NXRRXJj7V
LxXdswWJAVPz5TFFef49S6198z8+Riu8GmsOeixO0QiXr4rRViGnw1qcVfj0LxN9PSgyDRp8X34p
dctjeGjhFXk9csRlpb4b4PfVMfGIowZiFSFYS/59RUiBS9yNQFpzCpqvifvyf6c6EgZ9E8Zdu1XB
iqj+ECXDB5Gbuo0AAqlWAJwJy60CDWvP7Q1WrcFKUYBRFQdrr3g1+JO0O25NYagme1kHJys3iCSG
8KoLF23LpGqr7W+Cs6z25X5g3ZLWHKFnvlKcpaCFMXshNlGiDrb4fezPwCf9yurMVe6JfdXgj/X5
TwZzJJsrmwe3boeAsOMXU1kos13E0LbvnepE9tHnl6Dot/YmlHKPkreb7kVzcZbFWem82Ub2USQa
dxGT7o70Q0mOrhL3BQjnzX2jbUbfEV+EFfrOFgBkLpEdhwfuM/DaYmlwGW1MdMgrrPDwey+a2TD6
rHJqnwnvmepNqVr1xFo+IVjXeCxoR1sF3ua0x6PV4tUzuYFiAmh6F9HQZQ4yUCwWekCdAB6fZDVc
Ao7GvluP2icaYNAXevY5yski65mESZ664j+zIvJ78AAxxpPNe1Zl2m1uPUPY0ZQgl6PJLxwu1nNA
AWu9jXpP6CFJFoWuDOsejteoihQa+mCyMhBpW1ZGh1YyAjhogfn5SRcefQnIvqlm7c4ZsSr+kZjw
dmtmk59gMLOyHoGMgPRl4WRz6X2gNaTSRVGAtFefBQoNYlXgYeFZ2QLeWTTfSqhzuWmqBd84Efjo
z7Xr7TJ3RMycEFXIE0G4e12aphz1RSfkrvmxQNYDeo4HVCnyeyxVv7mfWw6s60ECpPBFCYg8OtmQ
JsFs7Ki3gT5VN9ul0q8yEtD51CkBIVG8qr0u7x/T05xUsWP6l3MzU3Znca6dTvPHVMd+q2fiTl1+
X6R6z4w0H9tUrhff7m5uVvKhLDcfhyW0YoJ5ZUqMLbJ8oZlqPg+TVmK4xOi2lk+9xzvNVS5gbDAf
B50oZkwDo/NdjgYjREKTACSmt7QNQ9mouNToWgMh0plbZJNCmXAsRHm+kNhPaoAK1oxS47sBbz0X
dImjEHpi+J43Gj9rm7Tbf2+WnsCPCBkHvsZ7rWteEUhqJVchohVW0h4fTFy2hLQMeI45casnaTVR
+iTnSGEeNDD5+igHEFh+2qGn+IBP/dBjOgBwdw0TyOXFWgHKLmFRPFbA7p1zpVS3X9mJ1WbnHCXb
gJWLePgYGAJtCAPGvqvhB1PEYqitSyBqnzLY0nwTIsuS2x0X3QAYl4DnQplz/K5HlRzyEEmLWO54
zKrW2WWJ4PKYXk0BVVk3dHUJ1c79XpgzSUD69F3SPrt5KxH0oGd/Boghc0lN796coYU5qCuSOq6x
NFMf9/WYWu6ttALRlWDKIrW3bCXJqt9wKxn5v65hBvqdA6vW9G1N0itnWN0Xx9prj378iJluXKxt
poGeQlEntgBn52Sx8EKZQrLvvpeE5lKhKQTlvK5CR0TLI7by+ioXCRSzqdTbaisVtFhfWUslEyvl
N1cFu5El4Ot9d3+y4ARHRHF26Weo4VMv87ww88JplaCJbvBSbuu67PEJV3xf8SUgyNZ4BzrJ3RIj
Jiz5SXNMKU8Ebto1AuqjqU1W99dVFZEMWxC1l34BIjHISRXokacs4Gi48Owjsx3g4MJ458m4KzSb
J3ZnZDexTbpbUL+eyViWYQJmTyQvCiAUdgQF2MpUJOFWhtfVL67KdDlzvAph3Mywbqjm+6rNXSKZ
yKe3elFQapeMebTfqcFkRvOHDm22CHCSn63moc+a+ar6LEEPWAjyTve4OISV0pKT5T2PogN0xO/U
YtEdngd/9x6iM73KUlDQuHl6eJWQbgHq8IwqSEyzFcpbEh1M4Kra0x3izgFOXu66GB/E/YSNHzn9
dF6zMh1tG37ZgkWKninzLn+0HBRpIPfDTrbiyt4vsPSORyr7EdYSI/aWp5bDGV6RtukL0SjGpvti
W7+My4NGnHboMiCMUxQV56W7gzACtI5CxQCgFu7Bo97sGMWQ/VMPdHQUUAaPZca4d8JCB/nh5TAY
I4KlAOihwBY9jl9hVJ9cmumeScdsXYK9YTm53OA4vho7qCfH5PLM9VSKJ4kI55ACUF5IVPeCWzFx
Q6ZpgcjsO8q2RkjW6yD6OpReMFfrwLHF7PHO1FPIm8e1UZDvJWXKdd65zWV6t9Ko2SVGmoHXPpzw
tdRL6y4C1HFuhcnDpDHPhxI0ds2A+FvqIj5qm9fvQ7pkaPoayLxI+ShPi7pc0M/d9Av0004KJRs4
BFi9qzGu5FcfO8lH9XNA86t7BFTkk7Rryzq71IFbVCWY66b6OL9hjQ9XhEVPViec1HBBvUSfAbY3
CwDHajH6ISkVvRoOsWOm9GmvRnZCXKCiX+qxpQ5l44/M3X7CFmKb8djfZtjUd9xNevPSWDf/zoOc
ka90hwEWRVse2eltQM0GxJVvEbv94xEB3Ud42Wm/6K9EkADOg2nIT8gWUHR60qP852Czol4MEwa/
5/FkOKQ+1AOby3p3ScJyIgjSFa7kTw9cnX4DjoCWsAdElmQHjeGE1huvU2qtkF8K2h582IKkHIBL
cs18VmN3kFXz/BTPoRnSFknh58du1OOJxWmOZ9fIoFjqkLTl3T8F5B56HZ/Q8zfc2KGqrFl1/UFD
FJxDMVzMMSIU+CpALAMeFXzayjXJ1vhdvJtVB5bYC4NWm+z0QdpisYJxJ1Uo1eU0DpjrvPuCiW05
BmsGWN2zPeYhGAUJSo5hZemNqObiQEnjN/sBv2LbWztn1GkmgDUs489c/8Ce5SGfva5RIP/008tC
RsvXUMEr+b5oSNK7LR53tD1kjYlgXoIIc+bGlPbFSzV+1AHksVQ1L64yrOU5dkkLc02RnvLgn8bZ
rCQ20FYhid+IRYhTMq0giD4MlsRtavD0hnjXVObcyv8hlP5qClnvDAuLmGJwOB8/McDzq9ffGwlI
I1agzhb6p5qcwUg/3DeTEuIWaxGYcoj/B2SFYQoT+A5FZIn/jEfaiAB9YkWXizCnJ7ENsDo4eTBl
GJD/cNytpoATl/dlx2Jc8U3NS7uZWliQDIyCRtM+P1AZIOCY1kj9GI0ew+nZ5xQ8mooOZDGZYItl
ZDGGxUzUt6PdpBEtc/aPGataQajpc4MoQaa/tdFvbxB9DP/crNWxjbWadpZj0gQR4pitgtbvPLYh
0jg0u4UgLRFydCKxzoKNQn2EAgZMwJpT00CSZF18RAWdVSBlBl/gSpprzfZnsFytmDpAZV6DSPCo
IGxReHzB15VFa5cN8ugY+5RpOJ+eXEtg0u682+O+MHrBXJC0eTTLStyeHj9/q2b82h6ODFGdx8+f
mMdl5wcQrQHdt6rZ8CUWCmE3Xkj+F+muht9ALCLkS57s3NPCLTpnMNFd9v5VfC7hXvOBmpGfm1+F
UHT/wUxTDkgy3fN3ABfzY+qbOZbXIyLWn1oNZh/jrObEnRTlohKQVCS3bNPfyTGC/JrO1//kU247
dWQ8Vk8Mb3kfmP9Z+idmUbc21FFRuMX2vZvsP6NvCWlK/1EYX0o9SfyuFFWnfa4AVrtvrplo4VQt
F5PaOkmjc0y+7Y7oupjsT1sy7uyhiBpqVRFQfeXcRNN5w/6ZWdDm6abUbCEmtQjY59GD+J5oORmd
9g6PQ/lhZ3F4dy8Y6ssyOiD87P4VUZE6vW9iAHrqM00E5Voi34+eN9zRYklAUZGpPimWhlitWVYx
HEKNVGZ7dqLTj+uKsaNJAGFfBZB6A4/brvRgYVej8o+pOdIWGSgfIdfTVZ/h0sYaDf6h//QMivjY
dsnGdWa2GIntrxY7wcGOUHPlyKB6/Rm/EhjPEsK+mLQKhOhdpfBF3B8AJ2y7Jt5q3trXW/seYJZI
zdQ+qwnli4b5BvKczCy3Rnj5JwQTqNGSX3L17NP17d9pI2/VO/Bd/hnBwzaDF0nm/cJ35uvuGZBT
Gj5OkDoERbCdpT3IcQP7JUPoBtewGhGWv0ONKJN/DGRIpgerp2u5d/2JK85x/ixgVN9oI7X2dH71
/7OoclcSpojSoU09U5vsvF7wRchZUJrRbYt8VtSTGVk5xQNfRmG9hwSwITdejpL2hBrKwpCi0aAu
cRLPX3eftbAkN8KtZmURbwUQDnvfLhjSLh1AIusSyx3cBLKU9jsdwlfOdEwQ8xUt9gahmJX3LAgH
+VSvSwyM+Yj3phl9WnanN6iyEtE/ed5OlbdGag/Kg+bj2jnC3Wd9/Ws9Y+26cUU5r+h6iPNs6ZPz
aPqJr/yNGaFWRyfXFYPpsYRE9s8yutPG2U4eTCQP
`protect end_protected
