XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��2W�A�(�F�����*�R�Z�F��qx\� �em��'���E�=�'C$o������p���D���,4��;C1U�-�<,�Ɉz�!-����>-���M�.�Jtd��e�I.�7N��IMR��2[C���-]������J�,fTc'|�����c8��]	T�+��*�M6Ui���G,.�k�kFX
$2@�^��1� ��Q��Z��O;�o���>_I���WL�K K�bj2�)>vT�h1��6|w����,�7M�Q`�uV{�%�c�����U��Hu��'��星������ہ0<�P��'r��J�	nX?9`SB���0-�ô�Ca��Х?�Ƙ�ғ��om����۵�St�U3P�WK�9�|�����CV���=�bqjb�`�����nQ5�tnl$�ښ�\l`�2>b><b��}�y����,�~�Y�~F>���j�RZ��NY�* ᨳ���y��  �_��6�?_�Q�v�~�\<{G8�3�W�q���Y���i==��۶�ÍV����}n�������YC���VL����^��OQǄ&��,�8 q}�φ���>���Y��`wG��i��^v�El&xbS���h�XG>x��Pw���F����*���o���u%F���u)���g�}O�~h�j�eyu��5�u�cUP�"hM��&�P�̝���.��g�:�؍~z��Y�G �Wyv�
Zq:�ߴ�XlxVHYEB     400     1e0ֈz!
�y���mtv����޽���\�hf����6�T4��in�������xo87���#�F;��.u�1����m-)b����4��v�V6Y�N�P��:�&ߐ�':{�hbApfqv.H���P 2_Jhl���[�.$���OeSP`V&w�"�������t�F�!C[f�=��J�Gey�%��f:�h�6��:fM
�X��d.5��fը�PFwA�I_|6;D*
ԏ�*Y�i�9@O�c�aU-�F��z�_�r�J�̠��r�ia��k�yAJ���Pp����kk�`�J&%��L+��'�ԸO?2	��P�Nd���\`[_]�)]��;���
��k@�ر
Z�'2~s��>i�&���;n�t�9X�Vr��ۥ�:i�d,���[�Q��pl)�`,����3 �9�K�ކks��z1b\�L���'�8�@�Ӛ�����H8����!�.�y�Dt{nz�XlxVHYEB     400     1f0�J�]��<�d�CR�9p�s?3�$�|��67����y��@���-nY���Wa��"����ޭ���l���a��)~�w7�w��^?�n<��|J��~FjY���T��q�z��O���ɮF�@(.�|�[Bӷ(��6�c(��/�DF�n�����,aD��6!ӜIT�Ԅg��?`ʤކ�$`������h�6���x�������:�7mz��e�lſx��ȓ^�%]�)�^;��PI����3u�N��[ǐ�z���eH������W�Q&���������h���K��pퟋ�Ԡe�%F�I!~�9F�1��~⋹���b�#w3�H]���9���7s5��,+Մ-�ƢӠ��P�ɺ;��[`��e�"uQ������ ��ٯ��(?�-zc���K}*u�x�s�zH|�	��Ŝ��o�10�����8.�����iRsD���j>23:��82�����ŕ|*��RXXlxVHYEB     400     1c0u��}��U<�^���K;7p��>���G�1O�|��gf�4ہ#Ou�QwwLs9q#�1�E<,x��BUp�	��qa�֤S�<՘�W�A
~�Z��X��(J54�	�H��s�^ �:IM���:K��ǫ�w����V^�3���m��� ���7�H�XH@҆Y�Յl�j��m.X�Z�6	��3'�����K�yE������Ŗ�S����]��)^���8��kӔ�����W?���9~��������S��T��Ms*:�.M+��u^i~�Ī��h6�g^D0	
�}iCd�����.��JaP���-�ۑ���\آܓ�J�[� �ufSb�e%����l�V%�Ȝhr��`��,�C�#�wMO�k_�.&|]��{0�A�Q`r�Lh�6������.Y��)+'�sN�a�68��f��!�zb�XlxVHYEB     400     1d0�_"Gc�FG!�9�'B�WR�*��_�����4�SȋP��&�+�9$�}�#z��'�%�ߗ���h!�R�+�
�8�{��#hNie �x4f�А�[:�#�{S[S����b$���<y��aDŕ���������dqS�|��~?hq7o�R�t��pmd�ob:r=H���E��E�G���$�d�~�?b�ޮ`K���%1P��μe-Bm	�2��ة�.B�G^A���d�B��؏[I�͙Έ'9���u=���"�+dE:�b>���=��oV��"�غ�������ى+����BX���n�Or�?���w�yR�$��%k(��.Y��*eI�]B8둨���~��t��y�J`�
q��Ts���t�z���0���D�����Mh�+�d��u�]8�)ӓ(Bn�-�h\s �S'X�Z���8d7�
}�������@��l ;h�+�XlxVHYEB     400     200g;�yGj��{�(0W�5{���r�s�am�b��L<��d�v��u��/~���]���i7�J�� /{%�e��/۝���?�}_] ��S�֟T�E��w�Ў�e�o��\��%
���hB��k�TR��C�d��7[�؟���8x6E���d0X�Ҩ�!mT���,�H�뎢�/�7Fvdd�t����w����˶Z�`�<ޠX1jf�����~��7=�k@[Ũ�X-�A�2��;�Nj����C�s��'�/���p\ku_���B��Y�������=��:�d�NPC��#�#�=.�9�u�֎8*�th�$b/�/�8<P3�Y��0$�^jGlo�%�����qR˃M��(�O#Y$���%�E$ox�7X$іޘX-Z��e�pKx!��HT��ciaI8�F���x���/qX!�B�-BR����*�nϱ#��߄*�%������dX�q�_<Y�8�`�<-�^�д�g��XlxVHYEB     400     150�.�gy4����-����ӄ��p<3!�{`Q/�N��:��j��B�Y��ϐy�.G�=5�;e������ �����zF�آJ�O+F��- �n\5_��JfLs�i��t߲�:�]�������[]�ֈ��=O�J�>A�V�H9��HF22�d�zd�.YR�4�Z���(�� L5'`?
;BBD.h��O?,~�%����}Y�L�K_윎�}|9���gf~��yIRƛ��?+�C���ٹ@��&���LW�^�NRQts&�U�݈�YK���$�r�&���b⑨}L?��}����ڇM&����E`N��Ҟ+�l�ă�L�XlxVHYEB     400     170����Ӎ./X��b]�{�O��@gM��瑰%��T�R���jo���;bJ]��Ϳ�X����W=����o�2X��?�XlcP@��p�Z6�����h+��U�Y�@�`��K8�M	�n�}��sW�MQ�O��E�M/%|�6�ؔ� ��j��a�6-v�)�N��M&������c�A�|=�ǈh��T��-rFzx�Tj��
�k;��Q��#�ʉ��A)�1��t���  M��o~��V2�o-�����&��aZ����Bl����L4��H��L�����b�� �� ���d�rоA�6'<�������Q."��{�ⶆ��d~�e�-w��Qᇱ^l?W���Yv^ XlxVHYEB     400     1d0��w�z.��Pl[Gڪw�p����?Z?cY*h-��-.��:�#d�SV�i�9X3��(Qz�N7���r��H���V��^`��S��U���(C�D%�o�����C�-U�z6@�C��I�.�2�s��.�2h�X���11��p5?�=��2��"E��fN�o
����1Ӌ���w�O�H����F�m�о�1���G��=�u��2�[��i���*d,��>g���"72Y��a���15PZ�M���=MD���=/m��IB�~d�5�Ղ���Y��)(�s���J:=����QA^�f��0e׶ �b�P�	�{����qM�׊Y�׹���/��>x�o ��KJ�a9�Akf����@���B0Lu�3��G��`�R�lV$��P�j��招ꝸR�E_,Q�ch�T��QRç�i1�]#�W�mf�(�v��F-3�{CONcpe��nh�XlxVHYEB     400     190�B���}:v�C����)��f�Z�q@KZ^�^�K�i+E��>r�=̛th���Y�^%~�G��OzN���*jQ��z݇�K�դX�,�&p������<ݭB��a�G�1�"���>w։!������Ʋbh�p5T�������s��������
��:�2y�sA����EZ��@�n�=�K�VLR?S�2ʃ��)����6�S��8��Ħ�Z�x�L�i��q��{v/M^\2M|�epo �����1I`L0�X/͗pG�0�宍�=W� �fȁ_��
t�P{�� 2�aLC3[�A�=$�a�h�η��������e��Tiw[����>��|��Gb����g����s��Os�؂�4��.Ct'߽�x��P�o���rZ�XlxVHYEB     400     190�lb\�O �^�r�L�W!+ !��Y5��5�4���̀�\]��aC�c��u�#�J�j
AV��=F������&���T��V7}՘�/�A�R�JTĽ��2���f�^=���=	�{M�1���䴠�
��qC\07nH8Gvrڠ� M�A
u��m�9�?fůΓ����xߐoq���ɰ��ۦ�8���P֠'�����=S="��%��Q�4�TR�a0b�^�Y	��m������
���B���29�e�9k��BJ�'E����2�p�Ohb8������)}���A�ﲃ	T���K�-&I,��axE��s�L��޼ur{(�a�j�}��.[�@�&������FW�t���]f��{2ڴ�qm,a䍢����S�5&�72S��QXlxVHYEB     400     150��᝗�鮛 ��
�3��$p��r�oN7��Uf���F$`d{f�b�;���N�p��R�=�k-���-2(�7��Eё�"��G�7@VLj��[��<Q��9I��)i0�@�͗;3���$j+Vr c�x��Ϟ8w+���D�t�]�����VɅ	��q�A�0#U�g�*!:w������
������H�|}��(��3mJOk#>����мR�7�=�+�Y���q�D@BP�U�q�-O�#G���ȡ�+�@�I|}�%0�ɉ��:/��H�@O�l|��3W���*`ex}טb���A�6{������Exxu3>�,Ib�5�ar�Jz'��XlxVHYEB     400     150���h�����l�0�F���n�t���[�$x��ٛ����՛տ/�r�Ob�^�e��@c�������D��Io0�in$;�0�e�:F�F�p��� ���$`\y�eA��t��!�Z*��fʳ�ۊ��{*P��������>`]�~{�m������x;���C^V��>У�\����L��`d����oj��/5�҄�7��	'@)����mg�6�������������Z҈�|���p�M 4�|�g��;�<k&ejoD��_�u�xY���i���0�5}p�`kHAk�-�!��j�Ka0pW�|Ր���m��k ���Ͳ3�nXlxVHYEB     400     1c0	�c.�v	����=�nz��/r@znI~"�XZl�zb����QI7O��,�AJJ8��dr]	����a���`:f����P/����x�E��˦�W����}ټ�M[۩}�L���{���o爄[�[�Ʊ �z"��|��ӎ�kx� ��|��u�	���B�P
��X����&{a�FakGx+�x��	H�*��-��C�c����ZN|
ha^ZD'������l#���U$�q�U�oG'��1�|����P�m sf!-��T���.7?��Ԫvz�0�ދQ�]˟D������-Q��?�@f��Xhh���#B45�'1W|��&���2��!A{������+�
"��T���ӵ�̹Lա<����9HzG��[.�Io�}�uƟ�t�k��('0s�?��Qs��|;i��/XlxVHYEB     400     1c0W\��Dl�3��_�i��a���S\������Q�jy�/�a�+eh_6�֯�=n��4~[}П�<�d�ù��T��P�?�?
JD�ex*��±ԅf����"J���ڪcw+ �¿+�4��`n���G�w&�>.�m �\U��1����
B��W=�-Bw��J�hjg}���"}�IM�2C��:SE�{n��:�`�X6���Gq�E#> �9�ߺ�f�c��T~���>����>�D�'������UJ�Q�Z��ߑ�6�)�x�x�#�M�Pp���'���a����� ҵ$l�n��X���5٦�ؤ:�Z���$ +9����v^�"�w���NG<�
SX9���.T�/fcs<y�5vؐS�u'ԴZb;�w�ᡪ�z�e�#K���[�R��&�|X(�j;YO,2;��r�`�ɩ��w�[	���k=�n��D1XlxVHYEB     400     170C�����2�@�	�'�Y�l=L��2�m�!\��#7���'��2���d�UH�A�$�C����|�ƛfI��7��20#�d�����3��C+�l'�a��Wbϕ��[f�9��òv�&]<VS����m.���1�o�v����k��H�j�ޗl��� �>��-voS��-f(���K �A��?���%�ɖ������/�`<Hʶ�����1���vOW~s�ٿ��ώ�ͺ��	�s������g6�,3�P���}��JSк����(��v%nv�o���N��TK��]*Hc.lhW��|LG���a����j�
6�?ߎ����C���P�C"T�T��c���Fe����XlxVHYEB     400     200���(
��yr*)wzGC`o#w����R!�	c�F�i,��X��l1���;�`:���ۂ�dD\�T�:���]�q�g=-�xV�
����禰1)�)-����g�5k�9w�n��^�z��)���	�H8˂θhu���b��;��Ζ´�/��|c�e��4����/�.7?��QZ���A�*���1�k8�"�F��J�8��{/%��r���5 @���	G�.j�_�0&ۖ�/��{v�8�Un/~���t�ϙ	��4"��d"����/^�Tyq���ܞ��#D���:Jo��L)[EĈ퉍6;xӢ��h������_�|�7QTFa�=Ȁ�cx��wb��U��f%�6�z�Šه@"DG�sH.S�x1̓�����:�����W�7Q�����XT��������g��CIZ�oܽ��WX+�?񥍻�ip�eI��uwD"�.?�>v����@�ThP��qf��,�61S�΢XlxVHYEB     400     210�o�Y�!���4LEP��RW)�����>ؕ��YƄS.���5����d7~V�����3��o,Ѱ\�DUr�Z�1 �b�K�c>�n�K!Vǒ��[��ya\�?^��	����'��&���r7��?�B�]4N>5��ab'��X�`d2Q�
)2˓�5�S=T���2_%�5��)6��j.c��v�'Ry�k�)
�M�(XB������&���m}�Í
�{���Ȓ����D���P��yk�ݙn������ڂL��Yϒ*I�g*�$�A�t��Dj�"���A�)�}�7|���oP�/hu��#����`��� c,�N��i�؁��4R�{���*�a�eQٜhp��7��m�w��i���X��P�ڔ����G�{�N)��"�}��٣{,Fd��V3�cڃtqCh�	�8���\a
�j�s�)�ē�Ã!xk�0��e�h�幍5���N��|PR$z�I$y���W9�ͧ^heΦ�;������5�*u��XlxVHYEB     400     1c0^<��l���m����@��p,F�32��o���we���cˍ���N�ŭwmC���u%ӧ�ݮ��V"Lg�~
��Wt�QyB0M��*'��B��쑒uiN������D2��ȏ7ZJwʝ/�C���3",b�~J�7��s6�3��4�0���g�{���"ۑn�r�_m ν��LCw�>P��:�8��QX��#�n���y=�j
y�r��/��2�P<�&m��*'ZXx��4��$ƻ̬��#��d�;x�Ó�<em�f@���@���5��
�t�M/��[���yݑJ��'x$��Ua���u�\"�Jι�� o9/Di�zA��D⡤�NH&��,3#�8f��c�r�OK[�b�M�.O�뷎��tI�t�g�IZ͹	y���Ti�ًq ��~N�R��}��X�3� k`�G]��@7��E9�L%���E�����XlxVHYEB     400     160�~���!�=F�G[�h��ƥ�AB�3.d�?�X5ύ�.�{iE��^y��F�
Y�)��6�xZ���$�tO�ُ/fU�J7B�e�O���.@�F*>��w�*�rB�F��6\��,˺H�ބ.Is�x�e���A��:�?l������0�VY�������ݤ���f҄�>�83�#��q9rM<xԈ�ñ�m�x	�aMgaFK��UaBD�_��\�]-�K��?6y�[�\���N�ui9@ 9�Gi�Wc���4���k�� ��N5*"����&�zX���!^�a(�%F?m���{g���6;nTVe1����0��"h�]�W��k�9g&�XlxVHYEB     400     120�%�
�����������4�w/�y�����'PmFT~)q ޲t�km�{=�t���b9Ȇ�3"B�C5n��u��t�T�Ƣ�s���Ŀ_�T�O�g�,��_�c Q� 8��vD}����m7�".?x��.!Ou6�+_������x���6MDh�����e'奧|����)��P�G��>�4~�h/%�(?%h/w�t�fD9��"=Vc2�F�_����y���NRa�uR.�C�}�E��j���p훨㟁)�AE�s��{q}"�+��Ǥ͵��XlxVHYEB     400     160+w��^:k�
����;#��k��[�?���|�>�	ӠM=Q1�.���v�����$ռ@[1n���Q종����7h/�ƒ��C�ч%�/�Ƭ �������f�����Ъ�`D8����T������4_��Qu��e a��]h>nlٖ��|+l���B�v`㲟�O+P�-h�7�,�r���,��S�ǌ��r�׀�7����Q"�(3b;Φ��J����X�F|oݟ��V�C��6v��XC��L~�)��J-;�@�}��y0��'I�jnD���{����!r�&/��..�Tz��Cr����AQ~�5����㐨��flwQcx�XlxVHYEB     400     160Dq7�Hխ�l
������ �S��M��6VӞEsxX.��Q����&Z
F���P�b�GG�!��U_Qe`w?h)������4��31`��d�
�gm�|�80Cc)GI3/Zfl�#M�Fa���aW��6 9K�~3a������|J&���"
/�7�2�ױڱ��dM��j	��?��Y{� 22���B=J��a��|�w�L!x�@����b� V�Ѭ���JN��]rh�-����y���cG����M��˿������w��5��k�2��Q'9�1��/w��,
���orq~��FY1*�q^�pND�"������	T�m�]6tf#c�U��XlxVHYEB     400     200�7J��hU��^�� \��E��K2>j��ž�ow���~_F�*����u��i��Ei��lu�yH�8��#Q�6�dC|��rߦp�8��	CE��'("�I��;�q|�������h?#X��'fx������F�m�����5Ш�kl�~)�^�푉$$��_�io�4�ns�m�hP�m�E"�7�)� ��hd/W��O$بM�W�� 솜��P�T��'���;PA�!�!!�J�I�b��˴�"Y_�m��k��7���(��h���U�/Z�s��>xPm��
�l��X�o|���:�y鱥5�ghk8<)�'>�*�
*�y�M�'&���
S]�O�_2ᩪ15d�2���N�ij���.W۾��`��B�w�D���oB)]��M����^
�{�VV�]���p.�k�Z�%��uPƅF�5Ks�ԁ��ד�땛���^z62V��t�����[q�ۧ{hđ�W�� ��`�����JqXlxVHYEB     400     1d0��fc!�P=C�kMɱrΧ�"�_m�����/"xok*�l�x������D��IxpwR��aV���#ӿ(��ˊ3��������Ż��q��Ɋ* ]�M5������e�Ì����ۗ	��S��2RT��Ήw�A�|�ś�b�J�GT��+vp��UBĢuRA�BE��j�4�$"��(���j0�R8��FB�-����.�d�J�m���z��e�!�Up�H�� ��,��/Sħ�Vd4�`|M�<�xFM�:��1O7��^�1��e�]�H����źG��My�ލG��"b6{����ѳ{��G�L��tB������lQ��7�O���MQ\�Uu"�&�z}�u�h׬�W����\�TPD��!!�h#�5M˰/�U���7,�33�]���qG��C2�p#�Eގ�T~HN�8�~��*�l1����������[^HE�!Ct��XlxVHYEB     400     1c0���M�m��f��7^�5.M�5����
��6�/ɵX�eC��\�G0�)�@�R������I8{Fl|�	D?c�Z���Cp��Nͯ���_皣^$1��<G�KGj%jR�&��p�tܖ~�$��!��u
r��C5�%���TB5��C�T1�&��Ί�F%)�2-� m���ۣE��m��C�H�~Hu��`�ͱ�;t)"խ(ol�ZZ�UnW�R���w�-�.�|u��
˙A��?�H���Dv���>M�zP`��_JQd��(S	�!U;�}z�w��o%?��i�W����V��b*W�f� ��a�1����`�0�e�T�ֲ?d���,�>��L����(0�B�u�'��喩Amc�f�ZY%�n���jJ�4����\3 �+a�qȽ?�D�X"���-n �ij{���9�.H[����8ł0{XlxVHYEB      42      50�x���Z���Xs�d�5� C�|F��5N��b4��V8g��x�K�P��0���CĎ�����G����@5�-�a