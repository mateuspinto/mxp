`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
XnzUbaTY3qJGmYtdNFpFVbKX9VNVz7Gda7Nr8A9UzF2lYVTBEQfmVPY7wuJPOGgkq5ZctL1nH/Eo
v6DTa35DG9AI89XfI24ImgYj5mbqlXajBL6iUubWBbKUN7wyee5u/TAx60B9TnSpvXA8yyga+fb+
YSnQFbcYm7iTezISgldLoTducLHit38WsHwlTHFTJI9Sc0mJXKxzMHwJ/7uWOMgrsDcXgl5x81bN
ituwAeGWIO+cKAPcIpC+K2xjR39nPQ/zWMQ+964jBQa6uAvuQeQ0XnKpAr2dmMgxc5dU+L/rjYlN
PI8TFu2ATEs8ridvIqN5eBaYrqg52balHN4rgg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="MUPifCUK8PCHJTCTLOH+AA2//Cy9kQ4f6hKiges2WMU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9328)
`protect data_block
NpZAcxH+chTyPXNYRhwm/IqHFVpazQSJ33djelYR7m+LNl8cKo3Ypr7ZtONc2eGYvmfck8852mKp
dPI6q9jM19+QbnWgQScc7rjV3R24nDIQ5XJTCdZh4y51RC+wig1M5zF0nVVPGBl+twugfeKnUqgo
fCNRx6nts77ajkwk59X8lYPV9qIUEirzScBLSAwRkTSsX6QHFgpCpD2TZtPUQnblsNvTzxThfbui
EtTJVeIAqQqVtCZWzbq8NzogbV0WeYt+Ws7Drjc+xf7RtyYea1e0JJhWNmZqELlY16BDAef87z3V
fHcSITzC+d0Xm3swLKFcZQiBcVu0n79Tt2y38H+hIlmfR8NK4HpEp7Zbq+LqHe11nBTcgd9EOB+I
a9U01L1+3WnnjtHglh58hHawRY6dOTV+p4odf212F7/J6lRHZ3naylA/yZTfZQj7aH7pwXH1ywEr
BVmr2gNs8oywHWCgwbk3//JPz/wFbpfWyexjuI66BCASItX+eHipeVOWXA+JsheQ15hq2OJ5sx+D
PH3d2KQWJyCbvzc487USJsWqF34JqQ7egIfQGyTxOHTwaJUlpIqJcAZQgJwmMaAkukOG3BD0z/4l
pA3ISKQU4Jc8f7NIfFMDy0OFrEWIl34Xsza6V4pImJdCQN09RntsWLsOA2q8JwUwZKyWO63L/ZN4
ey52xdKEn2aQm8b2nvvJUOvmo/g48KSOjrOOYd5SsL4afzRzBEhqvjmkKo4ODKOlhyvtbVIkdTBU
iDTinTRQ+dGRnEuazeoUgVkkKu8Z8rhOVg4RV1v+RLdexPr0Url3BEh+Tv21lEYciZQlWpJFO5i0
LIBRLgQgI3eur2b/5M2f0WUoYhf22f/CkOanKUmgq3ohuWhyKF+fsEUHLx1YXMj3OvwZ3ATAmu78
Kwm3s1aFgSOXMe9Iqfx5wOEiHVrJwjQZfeskRe6e9J+BKvuVVvzDBR5//7aoGekvVoBObmFM5C12
7KtgYtShMyjnEwGQSXwZxShvX700IWlrgwXg4UU193rJAmFv4HzKy1X6CCtaBraRNTz5LT2BMmtY
zYOFiTGFw9UZ2JbRTaTMHy4LVUcvYiL7VhmSYcQvng44hhgzq8IX5ycCKit9VENwfeEMkkJoVdfR
XR7PIkweKciO7Lg90ZGJYInj6KV545TbDVFdBeE5VsYHKQ0Klg9A+Fz6FkEXNlYFPmXdKuqrRYak
drHM1VvOoLW9AamyB1O+OTrxmy7Toku2khbYNtn2Z2XpogMo6bDg/nnCr6EUSRPVvxJ9HhTp1Ond
MLy36bNcH6AHHNp6MB7QB9HeKSznCVnSo+I0fPGUp9a2MX9OjhxpLYDuMGV8tXKeVY/IxXImALyx
8mkXRTVOUyNRjew7vvwuB+Y+qOF6rg0T4JWu0x4M3n5BtAEgO43EitE+AWxUfWBOp7L4V7h9ooy8
g0D/mLP+Yrueoljwt0Pv1AFLZgo4oN0YJTwYNlMank5Pj+Q7WNzmbhHvjaS6FhpsnYz6GMepJ+2k
cI/RWnuKnszBTReQXdqDRgdcY15b+7wQ8O6KKtiBdIaZarsw/YLOo+DBn8+yCMCFsvg2zVYTzQ9m
CI/oCZF5mur5/VRcGJM8GYZQArxHgEr3L2MJiUWcz5J3fyZEOD508gexr3uvdryV6J974S96/EeW
g63C4KlnjVPRolQq3X+nhE7AAWrmlxQbALR30ed/fr8rw8NXqmh11ADEkmkem4s85yg/zpvIstXV
EUwKZzWBiBVWpc0OExa7BBE1qx0h5JRdX8Fo8bavMjrfj3h6TI66aRIzwqi/sREMX8jqQWQ+1L39
bLMwcQ6WDEBJOrbpz8qV6Iwan/lBr2CF8FVPCB60EZg8w40KHQ+9b24gPOHAzG0RLLpwvO2IFP8o
BvGSX0DDPhkMpoxl5sEhtec9ed8g5YMV6NsTx3F7J0t6rEfAU6YParpY1MqctHMbRookWW4TMeQc
pGFMjefKLOqThL4WZ4VgwB0EW+0nHBLG8JZBTEDFbZRo6vSjpgDIWYyxlK1SFHTYnSk2lVAyvnLh
Fyt7h3ZjWOWNJ54vV5r1LHRLELSMCce3G53nJfsrC4NrtUa1tbTCzzNNo5brAFjz/am0JkHXgcUC
dxG/oFfgpgwc7coC2jjcVi6XyHh+1xWz+IfYP2kWA1Gj87yYy8t2gqwSpnjHoNPap6kQ93pjxQh8
dWORVSbHOESJ3EHnZw7nOlwlIHNRa6dXKYqtuuOmGpXy/HdCA8CuDWFtvkqJEmHIHpeSZX9tz2QM
EzQpT/HKRowABnuqCkdLo5NakIJWXUfAsknEtg0omwj00hA80J3CE1pfNuhFxGwVFC75y/GNe9wT
SPdcU6Xx1bxFOx8I0KvMtqRcqXCNsZvG453E5tntta9P8nvTyIqwU+zxh3cq+v/zf4xfMGsxbYTU
A9Wy6c2IJlTkFHGc5hlnWr5IcYnVbEvXjsRGwWLrRIbbiT4TRv8hIF2FRCL7jCkWYPDvR4tK8q4m
shrDhURhxMoeAGfs+eMeRCTs+6jALJ+stXrxpYnDkbf2YapMrdcZM9630vy0UkmyG0zW1dKHczyK
QUoDqtvabiMriR6AVNRHcdH41WAJVwkb49wtVis1eUsr0Td0OIec2ZVxcdrXuafoTY0BPBfojsmv
f+tSzpBuX1Dw55pvuDTpyk0r1080ZRLlXwDScsk8giiPtAE8aV+g6+RoEf6e/Wkz2t42HCo7vnYt
WPBAPYj48HfLBZ9jyv0gwHPLCkWjaZD4YL5NCv/SRiq4p4wxZoHVIn1t2dHm5hLwmgE8HzozRpxq
ThVjLsiaae5tMbdqpDtXHWHu5kEn7wHHlRO2VJO5srk6r/XtEVz5RKHTTa+VZZUmKHGcgc3MCoTK
uIUt972IGJsvWzs1w0FuIf5+pB2x7gOa7woWgW4kBTdDueIWQs979qNpCw6TTQUxhOQf8zqUZqEI
yY0STyZrvnTjsodnyx7/Wi/fp6h6mk+UXg4ZiGmTRPmq3ZnQrXMLFzsyYSsPS2o2Yp2oULV13y0z
IOKQeTlTmwKPiiTuuxLjPG5MFpdZuXmJwAwA6UWQ0+lfGwcScdfT0xET2uAr8sb6zkJiV5yvbr//
O7wmhomWclFyRnBPJ8ReYGPO9kazBOfFW0Yk13GGGlYxnFVm9HWNOL/oaWQ903Ix1CiV5rSOMH7q
D7EWsdAWDhYcbBVq0C4jPrAGXee0YORqZrmkd2uwAGTmu8DDHHWG5qSHtU2jHN4IKXtiDRLb+M9O
gQr9JbOU4wijXGa1/gKWMEIJdKzg4R9/dYUP7VHHouIxYN+M+POen9CVMyne70t8BIDct9sscLcg
Da/PLGh0nNroz/3rFfw1Ct9sL5wgsI756rBFNdiAZXlLdrnS6MZmR6Kb/LBaLWHUok/dKV2EDX4R
41Rgh77RbfpZ95gB9zz4ZUd9aL8DuZNAlVWzzah8SPhs7+TDlbaUMfiokELRQRB14t+3Q2Q/NjCW
4xHJve2i3PW5Z6OJtJFCMgDGp3JL3loJba8YuQVY+JEDW4szdSp1gpPCuQCTaZQUrM/P5cJBIe6y
GFloZwamMEzZFdCYZapEJ8o0AH+h5OyWfxcQEP7uwC62+NENqgcX2na9UmfrA+oCG14PcFbOQJh4
yKp/I1T+QddN22WWnLkBeaeplyz+wX24ImFWFchIqrSOCb0LnZrvhwD5aOLW+pnVLsqiFPaIgc+4
1dwWDrhAACUxM5s2CoQU8+Eq5G9Kx3jr7x62fYe7bGSBIhiUcI9T6525fu0lqie2m7c+wdUsj1NI
rm1aVkGlcqFM3XBWqh+2bFeeavcw5y9OfGlZTZcuZAjdn8bQpJv8Z4WrU87aAWxqSi3vc3Cs/wdg
8+8p6UkoDOsWTyGZGa1mxrpHqVOM5dQWRXSI8rFDwJtwKcB6x69+f4jmgHO3lwUzc2Wq65OOFJ3l
9Ua1rUKhIyLvsX/rRtBHiAsxeKBNrbIJJQskkKcF0bmQ1tVjAvEph9CadARYtK5icAUpadWWCdN1
FvHKhRFi0JtHeHQm4xKl3SvhTEtGxd4qddn62i/dCLXRNvSILTM0n4KLAF/zxAKji+BAHQRYxwdA
evxTHLFQ98k0iSCK/bVcVuOwRSh/XTFT1LXfJLCN1c78DWF9eVNjfjkVn7Ehu08dlxvsoIOHYrNR
sJSyouIH30ySRd0qa7uA22DUBIaABZy4fSZkpUjmh9LSbr3pEJV9rgomQTaoYe+jdEIUkmAuemtA
go5f4/6DHFTE9CENQVvWY3htix+CUd3iagYvwGxOnqCedwmma4rTDHXnUV3igFOekHN05j5S4fpj
QQP05rt1B335aHAol5BYFJ4j5DKR/dBl2J8S8gJ/KWNNmweyda7P8Jn6p5UhmmloorKF5z/uqB0i
1qcmsN4BiIao6ueD2AjPN6M6lDxiHFmXxgaitonYntXCJQRH/o75yMcH+k6TJjEdiMiDB3TDjO/+
acpCtGZLCM6f3uNxCApkbx2CRN7sfO4SR+GQp8uQ1VOjZ4GvWDxX1/YvH3OnYWdPUp0RrankqOad
4epgGFyc91OlRcjb+OBfGpj/DqsBa8QczVcocF14F2PUNADxg+Bu8h1LRjeoWj0RmQnAz7HjRU3s
9madeMbQ7lVHdJ+VX5atvKLWI01n/yTm6afACaYO3seGzaKiqftAiOeTyRNsR+I5Dz+APETx8qda
RTj4I4468vm/gMxiDhNLF58WzJRQHqkK3FHy1e5Elb4iTJ0kjriKYv1Him8qhfn/5j8QwwxNC9E5
ZBn4Qe32b+wdNA15F4ts8m8YsaLoX3BUULJ/m5G6O7KbnuANakKPgAYwQ8WZV3BCPlDImByCS9ty
fcTaV/f1sqX/esL+WOcI89Fl1bHFjBryL+Rg/SNjZIIt95x0Cf3B+SCzJj2e/wpNO2f4ArzoEHSn
5EIma2Ex+dQAzzj6kPgxORqMCDc0byeK66mRENJubPOJPW65jVbpw+o+JJTxEhGqLooVhuJ0j5+Y
5a5dxqFFB2dL2fAAd3VF3xepxrXvOpM9by6N7mvjZahW1DSpoYPY87/8qmYCMDniNe1+Wxm52+qm
nuilZxu08E6R0WAkTaCBUeJXXhLrQZpAzm8sZpNT933RBLbSUQUb+W3Q6Rqlba5sIxh4H0Hz+UKZ
Zwx7xBJJ/rZMA/p5VEn6MmF2feTIjBrCx1xXHoXNHj10BVhId8IhlI+W8ukAYKlLVdtt5Co+aK/i
/Zkr1w02b3WB791LU80J+xH8VqEPyMM0I1pHjKm25ZngHnMAbzCGkJ/1862FEwA2my75j6X5OTPz
aY0WY0nmRAgn8WTkKoiCqtSRDw1aDWkpd89LvS6OJzwYS9MNTZVpWlsptKJwW6iEbEVW6M6DXnrj
c2ttl6veZMHnGjjtpFAn92gKlsbrgs5Vi/vtZ3dJvxmxM8JYt96GYIGEIOjf5x0vSrxEIqvFvgcj
eNz5YrcOjbM9lUyWCg3pxD/dxOp5S9dQSgXgUdpIUWxsGCHDtRg6EKeTL6VswmHfZggEv9ONyiLD
lNAaOJuyFoJvUz1Fb/nf2Mq2SoD/M/eP5AbwhFyIMEliXWU6A9maEz8EBRcCvvuz6vqa58bq+cmS
mPTyPhYq+bdZzm5L+Ud6/2heRkfEzU9zcYlBz1stIVE5mD6b9J2wovF79RtvPonbYhEVt+HEFowa
hysXZti/vKpGDckX9ifYbMqsym1HCMDQvnSvwQhkQsoBY6SeiR2bHWFrCBYC2oJDDw98ZR15nBuu
5/BTX/qu3Bq7aFcnpa1ewa4r7K+/xg6ud/FJlPTxDTy01IjufEVGih3TlsOd1S5DrOJC4H5Vlwj1
+yMSguREJnCqLFKBJkBxwng5Q/1KG5TnnHV8J6Vk1Lhg85FTR1SlapVvxGHeeUNsX72RjduYkm/w
LuYYmBkuBRZJLzVvyPLsKPLo4ljEqCz6YweXVQ+e93WQZjVhk2ryO92WUq/Ql9XMRWm1OA+30/DI
xLY0wYqLyq1iaCwQx+kiY4ab8pzJPkFlupBCpwmrsVGeNlp3aoRgCenDGwxpkbVe9JSl79OoPtCB
W0T25F+bwnsJXhigH3aq+Tmc/Y00NrOBfH5rm5HOxushexjMRAQrE1Mf5S4Z9VeHGKMliXpkI5ez
uLrFw1JQNa9Nj0kdxet34Z6DHbQOUBvhSZY0kmGDsXvjs+SPesU0NNhT1dVPSmGQIaJW3eXYRx7k
KcFKwImEqN1oSk59CnzRFt+Ej3uXpoG4Jj/Xh6egM/B0q+TtCoQO/shc1fPPEPFruDO/0yj38bqx
VWh8o1Ut2Op2vhJPhPPFPVmqa2wah9zvheTiCn6ndTtKhXktHeEe23pe0NjF6oon+0Bu8xN6Kiq7
KuXsHNmato2IOD4OIb5wN1PdZ29iZT4d3cfBnRUq6HN9sGl4vrPcid00/sxNfLPDAfhG31tEv2Xx
liHC9ukpcIyxMJG/PQGF1qmlE0beVN+rTsni1K0OqZra68zI5QC/Bh0ACRWrsybi0z/b4T/Ao6Eq
pbp/Hy2GHBEIaHvFIEdpN8iCgQBRlPPxlq1l/htHAhy5+4QNKdx42mfv+OtE0MFdMjhyRSD/QLkA
VBzUv1Gtil+HMzIWNXQLNTny6bwkFblsHmrHpkcFl/wuLCanySdrDwzRohR5dtbkLGxPxfTXYvoh
tXNxOmsJi48a+ih7txjcWsBJut36XykdwHFVdPGfBRTpdURxrFPJPliM6Wzk01MmtaLPPd4ba1sC
RnvaUdSJODggnrwBjG9VDM4uT5ylzRDh3hahn8B2ByUrgzw2x6s3wwCRtjCRmhHDqFJBMumS7oTD
uT7sOVwwhhX/pLFn7tkyYpAJtgQ9BMf0AmwJRKt1YnTmGxbsTXpA2YPSTvYHPhOUhx/NJtcda2Zn
L3Y4HB1z0YkBsW6SNsGX4UYH9sY5bDlmrlEIWMM2MzLh2uO3VlHq7RTxzWzTOZvR+Lqr03IURSdH
cPyts4FdCLvg/nmY0kRoyVOFTMR4DtDTZDZWWAvi40hEk76QKzEpRuGRa24dR4Prr9B12Kze5nYX
y2xhZBlljXw6ZUikkAV/gVHGo8oJb8u8VdrBxAyDYB1BR0Zs3+1hsMWrYqQQZx0nCp556H6fmO00
t5/G9X+H4LFCr9xlR0STUB0vTmNoIHGvyvyOgQbFtHLDsxkAPyRld0S1CvpNttWD9MQf7GU6/2SQ
IvYZoq2LUzjS3dbm5BnrB1WCKpmhuipwN7A/BCiFmKYA1bSuX8+oS9kCKxt4JgJwhmXFzCPumVmW
uo1ZH7FbJVJZ007do4SwKKR1GquOHsv4bH9Tv/5rAWZFA+rAWJDfDsmndSv4BQ4VQoLwIYHcWTrB
yLUN723pqfOjP4GdxdbSdwpq13Sf8wAOcfiENo9FgRnqsrcX37OyumzU2mQZsaBPtBkh4h0f1UuK
PQdRyBlPbv6/Kh7vfWlCLGzKl+doaAi45j5JGJAtExSDDgtqgq4XnTfVMH6cXxWIsTpl+JQkv8NJ
HenNf2SJMD0iwiJ9n1FqoRhWk+ZnyplJCPXxSuyMEIG6rMjp5Ti+7mffsg/Q5yo4dKIRNW1VJrV+
b9t4k1QAGKbY/EXEOUV8VdK0joBmYTVPLO+6cV6JW/EK7aG65QviqXuxWRZ/fZKIpnhpWDWHbQEa
fMkPiUN11NCn93QXSNR+/FBpRqUKzm4risQWMnrZjvXMR6TD/FzBa8I8Uqas4eEsTISzvZxuPNXO
M8kn7YinMUKXhLrUpIkKcUFfgWYDHtxatiT3baw1/iRCn3OpsxMpt5aglAb27vwnKj6lJn18jy52
d0kpdOWHBJc93K/A5OcMEaYH7MiGQPTqFxLUTcD3eBop0kn2MEzK2S8deLsVccBKjJjvOzjLkeu+
U1r+wGb0G2MyeOuojy93hDQ8uxH01w2GauW6jqnHzy4p0ARo0jnMbt//hqh8pO6DvwFI5ncRnw5q
MmvMp1qL7bhxV16eANrcsdKvPNp7k2iEG9Eo8i1u/GqLIbCc7E3UIpzraXuUD/vqDdRSKqNs2fNF
4WXL9dWifEaFSUbZ/NQx5i3KXGXn8Vbu5VjL/mXow1KM8VBBLLurVx2eSDZ0Fjy7byI7n6ZC6BbI
icp3R2e9UhRc0PXeq3ymUMMiirfK4LHR5DzEB9umtaNcw4fsNICVrUf02JqC1YpUnXdpdioZO4cS
qfydaXghQXoO9xoc1/Tr0SoHMBsTtcrH3E8dala1x8AhCMYH+bL86GspGgJuhkf767KsCuP9BPBf
JfcQ1QSHt3gHbS/nRVelXPKwMe6ba/3+db1fV9odv3+FjPUe3ZvPm+IdGnJPDnlWemHEOHj/zQe/
4xNtxnMfAvilJBeJ27dkeuzWih5930oNQkHWhXA+4Wu5Cdtd+n1Rg7HkAlm8xmN3zTpAk9TqqD2z
vOuuFH/2Dl1gxJaQiZZBNm+WOewMye2cIDDOX9qwdD0QbVfj3fOuwN6nHt9S5DH75xUTF/Nl9DHc
+I3qo4J63+dEql3ZWx3j4YAulBWMYWl/rAJWXhszTOiTQQC93xTWIg+rg3xYTIjeuKYIZ42n1KkR
Bt869C2UeNH0s36F3/J5dXu4I+D2ScAp79M8OJAlbL8qrKtfA6YIiD61sTAnFmgta4je0vkdMp/1
EEgVYWEArbELrqTHmFIznFktm4oHiACRVWYEQyX31vfd5zi9XdWk5qnDRD/shI1uqFcFQhQLn+rH
Zf/ji6is/CgPoYcCdi/Q9sJyD3b2QD3ycH6MYO6EX4zVnL+zEpO82hEPrRW0UMafCjakgI7Ljppt
p+TEnSpOdGkNHA0HSWX71pGSmfl0VGTdVuG18HTc/V8JQ6cXlphsLt26vGuFSkN+anMpkhhYy9LF
PbyXGMvKpOXov3jR8cvYqi4mmRMuaz3pmzJSncdjnbHUsIIWCzNBSRRhtPrZAX/kJ7/YggE5ceyH
qYZUrA7FfsbKzSk8Wo/+l38IX9CIGUNzbLcyGVlYjDYL0ewhQEI9sJafy+Y2TdQhnVPgjM104GAo
Uh7LFi+gzqMilEIbKiqwCBMBPDOElUS3R6eYKzcXJ41guK2LN61CPgjwOv9q5q8D3JyGzvlJA6OU
fo0UjWZ4XlP9jAbzV4OcQY/YeHTKJDwIPIt2q1q8Gh+mr06lfpyguqd85Iop3N4rQALWMX2F1+JW
WJlmHHIERVTYE8Nj2HAw4C0icILigICZt73D2hS+EI8ftQdixOTECX22Qy5ZkJ/LC0GawKkNRUhr
PvuSH3NM3iPTwy2JWQ0nIpIsv8bfuGjixAadCZCOWduh5A67bXCtGALtY+LW+fFSazbX0n0P4t0i
qQu7Zo0mpm6iHCY1g040TxN50EPBdooae7yOnhJe4GFvPeag0NfGzn+Q1ujNgMXFHBrw8xgqfRfu
H20HnHtE+M3vbWe/O/eEOUSjHeBApuWTl158HaI8Wd2mdf+1ddMlP1TurSR06rvkS6cm26Z/KIhr
rLKc/q7kqd1ZpvWCdfvsU2pTfNsPDVdxQ84gzbwRm2YnDhYxoPWP6Mcpz4e2Wtid6mEdpeOzh+cg
EPsa2Fwn+cC9qhOT5Q6JQekbIxqTc/kAnyIRmHKjseA9yJqbuj2mwFwZ8uyc7Dll/Gsqz2UWWutr
OEXTcBOT46KBdu70cfKRaE98+n+TUEygD+aMB8zm4cqOtRWz14p5ta8NQe/YBRm+NFmprXL5Qe9z
hV8cJpJ/xUCyOaccuoOJTmW+pp2Gpv+evnvR6vC8rvdInX96XYu+EeDI+UYVCwll4/n9r945e9z6
cBqHFJEQBKA9s/+DbPyWgNrd9T9wyVWjJgZnn5m4d3tzi0ODuc6JUyaamXNdJP1eIeyQ5amLZ+vE
h7LzSiprYnUGCPHiAostsoldfiRu9PM5ej1MMqlO/Ivf7gBrM9d1cjGbd8hYYWm2yAlHjkCoUVIL
yG0fFqHqMUyrZDcZi/QhaXrqkOvGiJOTeus+0Xh46je4+x1dfMdIVzXyZakwUou3jLg0u7yTuQVL
ec9PxPV2xT7p/GqL3wOKeanJ8ZKOPafPYK6ekLRI1n9cR4rUEI1s5ouHxiOggR00NpRiM/+euy4c
mVtnNb0T7P4oPrlqrTJBuG+kjspCrqMBHnfryyRwTse21IJjda0t+8wgrr7btzLESAd+YrmrMsdA
RuxCINdFzWPQyjWk1oVomkaWs27/RFJlB8ce+BcyKbxhNFSC2UyElU+D70yGL3lxJKfsjxneC006
RpkauzSPA0dVyE12RVeBEuL80kS/Iw23F5uE84DAxEnlGP2tvnGFfJLfOB+hsGDtG1PF/k3+T8km
wFY/sMvUBK/CHEYsVXogl+eHYYm/YyHBOV+4t3VV3ak1RB4BqHrCgwS8+RkGRBS6JIHVD5M0dLDe
wDA7DL6V/QkbsHr2/qLoUcOS4XNtbP429o0FtqBq+rmqigD/DYBlPPTS7aKIod2sYDvOY3U6m0vU
ANd89PigW+JOLVLE125HclYZpMs6knlllPJBVgT55eeVaDfmb2X/Z3qLLFVZoH2sPWd7XvZIHp3l
DAv4sXNn5j1gF5x2XzfK+vfv8J8jFH4E5m7nEMwmxgmgrOX7ghLwVBzWJ1ugZix0hl+bhpMP3vlF
n3yea1mpkgOgdMBbmGhhw+Md43OkmrLR8qbUzP8suGQA+zRoCVzT6FHNW4ziXmFJEgjfZyko65Va
ILgX2EllE5xJ3z5W+umZa+Hct9FktdPLGHCpQGMfZeuW+NCTGQokBmvzWJhFfkGtDFDymPAz8M9X
Bokig4whXkBAyltgfGLFauE17K4QfK+Xjh8Qp5lG37gsxlXuX5decBHruYB6btu2K8FrvOT0urcq
0GRNakMjumXjX5RKawQO8+EMlSkbULL7OuH5qOjzaVlCsQlie67CbxGZgoXlU1K+WrJQo78H4sEt
iUQk5QBDgXje90cv+KOkneOt2tao+wvep+/y5kLAxu3x5jD0pbmjHr93NPvTNscyOWoj77tOaeR+
rF/hzrk2yhBuNz650HixJJD/kUMJU+TV9UhoIxMcuLYix7grynwzI83E11YCFTrncll7YJHKRg4W
FfjEt/SN3rFXhiUctQGBLaw23A0PI6kNd719veGYA3Q341mZWvZlxzC8iOIcOQ4YQ53+gYyjnQq9
N4WPg7akO30GXbRqTcYOzSHqWE64gIj1v8rl1pHbMBq8FqIvOAQd1jKDZm8egXLpJzFLV1qR7ys9
GDM3y6c7YDtMV4iGDsVZd8YmLo1FFS+T5QQwBiU6RygDrQ0iZj3ORFqrsZsBLoIGkqsnTjP0aOYb
Ea3LocCx1E6gMRazwY47ubvpqk4Iyoe1bqK66+Y+kg9A17sq9W/u7ISx/kNvXm5vBpb8DSIzNS/4
ouby/2p2xM4VUqfB8g1DoWSfAYwOJ+rdOkFdU6oyO78q6uI4pGbwNB07HV5cJA8xpeTnJxLjt8dD
ERiI3aqbo3hfHsGiBXshVMlarYWjcMlfU2KMKucUFiFRnu0DmSL1TEIWRap64tQ67ITWlBm99RQi
eDWVSfpVmui6xWmVDXWi7q9q/XHlN+gn/JNUfU+aVvPIesFimY4nwfLVC1BhZUn1tCtUUW22YzvU
3QMt6pE05qDPxnLOf/YZcdOWKKMHSS0bZJ7GSVRaIG1/FpVaAZSZ/+A4cybWSI/4q/WQSk5eoybL
+0Ybdd7U9D3tFuCgTqV8On/hTNdkIAYP1n4kcvT0xV2IDzcuVEfR7hBy3AfHZlnE3XwUFElijvx5
m8/OIwxyR5/fFGYCMk6vaUAeQ2QOg2ZMix5cAiCPe5BZiPyaBdtTVTDD5TCUTJHKW4nR8anAnHZP
4bwGsywT4oIlZh+XnUFI2YcaJo4ZAN+caItY5pUDIxbxPLvOWt7zZRj7iTVLonYGQnHTbmD0SXTr
huQCioWHFuGok7u1Hl+dZWDm2eI8aKJArCkWD49nKHZRNJ27OeicFyNQSsOU+aTgRwkDL74OaBoz
+KPapivSv9ZtKG9ot58apLZMgIVhfH7MFppR1DTAdVSjL0QaNrm28k6tbRVHFCoyVAr9OeG1QSFU
FM2T+1Y/abB8xE4Biy7bu7Rzil5hir77e9noN3XuEAUnHl9zG0gfbvKehjxoDQOZXfYOAvJV1Dwg
wau4iNZhiYD3H2o6QXAFOMNFVMlHaE7dL8iQ1JhQGRVsV0ktyjHf1++Wz/sBksh1YzLIXtLazH+H
vTnGm6jpjFsUXDlQwhFBlb03rZlRydornLUzPDHF6rVPQVI/vVE5KkTllhwgRnp5hWmvZdDPxQBF
yYyHlolS/c4LfXMf1J4v5CO9b1Op64P60byZx+GZ8/JM2/6l6LeU06AaFnXr+SCeXv+Pi85JceCd
I6iSbvAA1dpgt3FoA6IzjGnWB+l8V7zyIvsSqwhpF2Xr48W3Pw==
`protect end_protected
