`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
nKpv/THrXH7govhJxOrX2y5LEDj+utqvFuZiUV/UqdIUWitQeSEkiJO1JX/BQeOhyQRO9FuVW9lM
b6kDnmslp53mY76tc2VfbsEhgYEB2f/mANGPyEA2F9EKLdSykd/O8W/amCKr9YY2UG2oopOtnv5n
D9XEjY+d133kE59CeO71MdLDkyrvZB8jpk3jffSuB+A/kD/2cqS7qIjJuVK3xsFQ6vSqzaL0XitM
JHBnwq9GlslWY+J9I0CP5Xmn1ck5Ty4CFYOrIp7p+sWPGVHgeRQejrMgKVX8GvbirX4rLpV0l5Wz
EQ/y/eqsfOb+n9B06NGP2Cx7H31ucrxJqElrdw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="31xZ4OSvMorFVswtwdAlX7mwcLHIl3MgV34/htK4Uq0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12544)
`protect data_block
cjHqMRYhb91/HB27tV5I1qlhwSbKmq6upzau1PYnNZAopDnSpma/D9eksRN6u00M7Xs3ak169Iop
phoxZ7HKFEhRFc2wkcLvCMIwPfo92DJAk+Tk4l/CsHadygpao6O6eU8qt1Di46tRYU3y1Ld/CxdF
ajh8gu/AJ99gdvErwoOH3xCNgiRJKU1esF7WUzDljeL7+WExtL1o9iHQDFF/5EnAdommiI9Ct1wC
3jOq2VBev+dT8t65aaSTGDHeq5IM0Lkj1u2ZG7D5Amu6ixfVFFOkKn6HfaXiEHtVV2VZPETv3ckl
/5csTjPlcXM4bzOlI8+HeWb6OK7ii8ZiuJVKtkujCjYR6D1IJXvbMi1Q45GMpqtSdPTA7YGu1Yy8
tcYw/O29//0EBlscorxoa9gaYkXrHz1GCegKtsA1FgD12wU5wEIgxSpqZA54ZSFmvhE24e6qx+yK
WdOxxB6Mh9NJ8O2c2V8PdpUk0xlgBneNUAYwBIprhy+rit6iq1DXTYH8NDo/NZXp/k9B8gMTr5yD
bQoOaw3ItOF9eI+mh7Znr0hw4aiGVPvSHm7WTYUKMmaIKKSjAaAu6IGJHBGA9/njRfO8RivOf0Yd
aDsrq9k3fV/f8DLvBbJOI9Bvne6KHacaLWPUV4m9WzIhuaADltLtRPXt50urd+i0R3ZwGsF7BRv/
VDQoB+aAotRIJgNAwa7I6nAU0hV5kkTcgCE0C15kbKYoOBITATIPsz9XRbmV2gDgIO6pnAktdhS8
D4jPFDMfjZBOvuZOGNtw5GR4+kvea4IUUGrnVSZky9FwltUoiVZNY+tqOD3URdnBrtlJHQ+fB4li
JS0gdrehMNmvmhxlIfKUk3DQGEIGnWfajfWQrD1zOse4nx2nhiXD0a0D4bKKnvCI4w84JlMVwqFh
A1GMZixZETuzNKPGu8RfkcjuOyX2UXE9qP84bVqexZj5kwtyZ9/LrXiJcHq2oLDLsokCBTcW7b48
yfn3P9H8jI7f9V6HNgK5l7YEMIyl0eOQTbJRIk3o5mtcrrUi7uXSyhuH9LAPkjACqqa3MKbEDRyP
R0VLoLNXf5qRZZuK7rEgpa2URmll1iAmVwaMJTf84VD69oM5mciwqc6kE+eYlPyBdvDHx+1zDj/P
O07mcC+M/NY0AIvbGW9TwHBrzdio02pDcbAFz2/Fq/Ew5r8qAs0ByQnK2XlRQZRIxvkoWF67tG0S
rSAyXJLacoLw7zLribXTi/7uJeNG4Rxw9U5j/9+88YZGjCkA7he2UVrlDYjhaac6uE08q//ggEwE
f5c2hnAf8b6J7wTO9sj2mHJmWtcvOj3UUDfzwCkafv99t4I//l8azFdsBim06gWxl5BUAB4urpcb
3pVm96egkO10PN0WX4kSONDD/JYD3sl+onizWBH8xIng4SUf7nfuo9M/4qAuRDD/YMIgpDxTW/4o
f9HrQR430uRR7a3abk6Bopt1vplntEbbf/bVS/q1KVF+SW0l0Vm1bhVQrfX3RMpdJFL8NtrHKdJ9
+5rCx9al22JPLORZDMtil3wOYDxbROAhvqy5dYwzOeVr6MFn39KZoaLJylSXwpxJsFp2Z3xGVGBq
Qa2iNyU8djEx0cWJJm6xmm1It7HBm16asH1RbIFpM2jVhDWwOQ8n+UT9RtgLX3h3YqRnOvLoeQky
8HIh92lXi6qrS2vaWj9O8TNMwI7ZIw+AkiXooST2Hpo53lXFj7d0e4Ew0+EYzrdDZ4pNTdOV0tpg
j037VAGJvv6e13CizXFzvqNodh3RQU5j+SFZDTw8CMum/ezfIsVuVjZFv812S/BOEOGoI/dFA+pl
gdoiWevsqG1HKq6BNgN7v6lBDMKz5lrgAMEvb1r58Ck7rg6Go51Z9+iSisJUXS8y/LhPnWj3MI/k
CohstYEErYcafzgLMUe5KMPbu85juoOwKnLSLHGSUT1hqyJbDkecccJDAqUD0Uh9Di1I8APN0xUH
/STtPovaROMDdXI+X2XsWbSPI8SDRabTqXfcO5Ec92Vv109zypn7Nxfk/q/PBpXyTW+n31U6A9R6
vyR8GvTGSdhhmRQXMjliRxa/bXYtj3TWxki45Z4fWo1s+VVCcTylxLlmhsIKjvM2WN0s8h82crXy
pMcmXzqCrg5YBYjc+BCFg1QQDVWTSKFlzq1fuNiIenK/FT+ta4F2InpgM5fmFS7ocG/klmcVE8E9
VdmHx2wG3w88EuJMi1LDQ+ba4cwIhAn2kYdIXj+9ej6ym7M4RpkVfAm0nse9+nGY9PN8ytifL09J
j+1vcS2dsLfVGApxIjnpHxE92zMA3nPnckX9zddhxdJcQU7QrcOx1JRDGsmfXbQSkIqZqYDs+yk2
DH81/9KudQGmde+xSLXFz7QnKdZsDJTP3zQywLaqFH57OB8vvhZzvEw2WFG2PmxBkd2xJAFK42es
G0FQiO2SDc241ypdSCeNjSPNZZsxraWwEf5yJrZxpSboux/gaFQz3u+ekvmE8Tvggj6GgVMvcYML
azskIUSXGOZfGej9HKhQGWURoPBUllik4EvKPWkvV6nRitNuqYbMNJU3GMVLximkX6ZHMIlU4Jq1
h3OHkLiXDp7DnIsw282pdvDtxn3FX1v55uE3NU3F9qfBSbAcSlaMu9neJc2dvQzB1FKIrmjpMuHW
9x/GJZkER76oBtSvMHPgGIK1GHnErMMCK5FZ8IPt/VnEfKJz/MLHhNNAejpV/g/HI/wX+EZbF8dX
vY7rKtyNVa5WHIabGTZSSEMDEpQwxCNkPaSBOmFukJ0b9c5Q+ELAjJI1VsVyF9p9hVWy+UN/Lexn
+VxobX9a+a1J401dByt8h1XQSeC3ueEMyXvzbSTYQODiTJcDAl3v/+ZpwrGm5KhUt1Fak+KKDAuH
B+ScrQkDUDe4rg1KmVYnBQ/lRrEHu3hXovu0nizH9K7TYml1yzIp3v8cpspUqc1SBhR7SQS2QdSh
xo1ljpL/fdEwYYtGE2oY8bFGEQIP4Xdntg8bO6DI63zWpDAflN4LfvtYqLxNSKdNDAkBJu5q5S4E
+kjmbNie6jjqByzp951GaImUXu9xVUzhMbon5eIOdOw0K70KS25/u6LDVm7S4yEy33prvzZPKMcc
86Hd0rbzmKlguGa/imu0Jr1swZ5xhr8dC7WSlOe7rLvv4Z5jkh9tewKLMbIgVwprkAajBmdROjZm
2465DhmZddNMkPNEjOEqOjOQ/2JqZcJfV4J+jSq5md7/GGHZzZgd8ILjiVy2ScofJIZDNY71IbRJ
QmSZyfXuwe7sVP6ZVGZpjdI/Ehn4N7guYWNeqtDfknc56I7N3RbhGGXbvv03MTHCrkbCVbgoQ1sX
d7JxcFCawU7G4VrANRBpGn4KuNRjMBEplRZewUzEvJiN5zwhlliQqy9ihsHpcQ1o2o28inIFJGvl
wGcHLgM0QP2JPi2ydh9uVQ+XoS/QpY6eay8WhwMKJYu4NXYTwzAWKJn+Rp0dXJEEuGnVErm4VERa
hTQBVTk1r/Co2Pz4UxxkpQDXTrBCxUrQcvR6A8tmMdKhytkwcT9HOGWEbIyY92UTrJ+PA6Wn4UkX
xDxu/TOQfYXTPhuj6LwuZaEmQlJAjWz4Bu8dPxh+cJOaZfoTWZ+/DdLJkoLJECPCOhaJtWKXPsqH
H6Sf08hTgtuSPPw0hPwcY+NAe70R4mEYJuwFJP/zuV6eiYGcQ2At/FVL2eqrX85X9u7fn3JiksJa
c3BJDRp8iGxv3YEUoh0bhQ6KkKV+PQLGWSgX7SebNROSMGBPsBKXOeNczgPMeeZ2edCf531gV/zR
wf1AJz44LBNaaDMZ7mP+mo5IhE/N51ujggv71hj7nq7NB8vOXRtXGozcCmpZvVqpdAEZYQlhCVyS
aePLhcsiii0Fs50HJSMQ4Y3Z4l/aZFbHAT6JfnojkrXcu+yyYJqKDyXq2Zv5m6IUBKCaxmRtqSC7
WekGnGEBRNP6pTXmbw7isaiwHagPppEVyVix1CCsDDa8A8EU5BhSVr0K4S2KIGG5E6uBzn1fUHXj
LXNq9PViu+rc/XDAw85osik4liF0W1tke+eI/HvcFiVdvC6w0bbAdc5UUnR16d+ab+A7/2+xhMyi
j3Ozp5iyGsfAJtBBDBk/cOsAP04iNNN7zqlqJFn1mWfp3bXgRIIMBYGq4dotGONtoN2WYlP3HTu6
VNSC5H1PUYXM6xmCtwRVBfUCDg/DT9isW/ymBnI8oubtm8vvlVEkfPFbwbc6gYR1qmMM6s0eVXB8
v3zaFIdrKIeWbGd8bqtXSOxOwLfZJZvVlPzfiQ6f7x5dIeJuuds2zGAxYux+qO0JfAyzGFA/FMa8
WnO+abUnTY3Pg+65XzKBOw8njb0I5ujX3Mlay5qOGeNnVKMlXEI9UpQvZCCElvxlROkfh6Fmfc74
qeIlIxJKf8J39q5A1Tlq5JOBUYefwCkuFzPESJP5Vn5qUgrHzMtQYbeqzyvlFeg75cqQnPMESNp4
RYDPoeAG0vHcvrggrqFE9udCaPV2cJJAJ29dI3Zd2a5K3nQb6wH/err3W1f4HY3Gjl56WoDPVFtl
zTjXnHAu1wRzTOutKvR/JjuIbN33HFBkBgX89h7ATk8YqMdTr0dCO55WmK1zXUneS6b5qg45j2yT
gLr/FzfKDu0dxU+kwXv47IM0TVrFn+MvAmjPMkXIMn5fJeqbN/rMdQTP43uUMdv9BUsDzMcmsht8
l0y8MW+7PO+o5IGRXbwtZGuFrnByj2GKBSRxMwFORUFOhP96S4YDmFSSBpgAuOuVqGwf3XKyiCJ5
I319TUvebnvPh4uh61XwwGhTOlx0iyhlwe18EhtwKdYYkageU5wXfQDHC7lrhGAH31iYRRe2bXdi
zf4r+A9dA9rnLN/lixxGwxjVwPVD/KupHTu6PxSmqUr6XfaFTCsh2cKrYC5mGXpjTnek6yDXZvoi
/62attZC9LG+SE7ahhjqtrNYe0rj7MHYkymKJ5cgeysxn934UqcPIlbgzVPjB4B9qtNun8pjos34
VV5vPwUCSqo0N979HujjL3LfvtN1rRjzd1ibMLh0BFt2tn5tZU/ICMEXDazfI57t7BMhvOmwEkFb
Qc0xOXDFJeWGbZOB3GbGg4O13jRq42HuEu+CA6YXNUFgsaREmIo1SaE0TZ/3TXdvzienLjzrzKNd
8rfPVdOuoboDrwoUSfCvb27D/UbfNUNfdSctiRRCOv0aXzeIKmJcx1MXMCtHbWdHsv6Dbg+G/91Q
rdHMhT813qS+zRLUUIE0Lkfly4kzp3BlLjaUF3QFG6DCMG8q95WuAtW91BDYA4AWOaU8w92Gfmwv
9VT/CPbH8FFV/FqNVGZfaGFcco8sPDRAhmY9HuBjS7Yt5s0imKKW9GWAuaHFAcqVpusfs0Ihj/Bh
ofqD8gpuLmShlIe0FtcwcHYRPc8NiokJ7LvQrDQLB27c27ntO7iMCnxML1PFcD1sNLFOHx/LuQf/
WC+qoofERh7nCiS7989jNTS++pvPQ80WagtWeDEv1vDhV40c9U8jjacyxWJQ5b3aI/G33jBvWtm5
WsGuzIRz3zeehc2HzknzgPoV2tN634SXfUaN/h2/8Cm96gg/RIMfLenZexz6+oHB5pX7A7yqe3Fl
tGiYEYQMZYxl0/W6Saj5PJzfvzeVAg9ShMAKDMCTF0rlUkAo1zjbo6f/NbKr5zEA+ac49cyrENOy
aonfLeye/Qp0Eo8RNH0wMm1cAahdgBLmlpb3a5v0JtNvR9dU4Fgtqb8BZQGdcAjNJoVE6H1ZzLmE
yzKesUOUUWRXx5LEV8fOKvPgBSEeYzX+7UrTuMSVAwhzF+aRRPzqNOHEAxdWa3NR7ve7QhOziD7S
MN17qOkLHBnUXBUHbo6hLGDWE2twXKVPXQLlt6+wcEK6AlAE9poniVUxeIWeNaBBtWy17rN0ZL1x
i3RVA04c7vw5EA1S1Ch6j/XiuNYa2bRMA/GBhzeZvf+eZvJCxpHTmk+gF+sa2LcLBASktmSHwqL/
ElK4pq7TxY7aLJF6rv3YUsGOCr7gLfprIwoyeZDPPJdZ3i1mBeRcdqv+/OpFuHN4hFuhzJwmAIre
42E27VGipLq6ke17oSb4gsNgpsl2cD45DEmyoJrRZpUYO9KzIyLPHtwWIacAIszNvNXSmD8CcQk8
QSGFW9b5jRr70AegdaI4D5+CLKxmznv0Mo7Wdy7pVv+KJ7tZNe9VW7vKY7evrjBIVDI4CeDmpPqL
joVaxhRRwY34FYqrZVm1K4t3EgQk9cXgO2A+VLPw7QEfbKKCOuFfokxhfpTwWtq9qn+NwgJAL8cn
byAdWjOgkrlPCS+Z1NWRVGzkK6BiMvuc+7j5355ZbaVG213qVBFraL2LjuGvak683dUFFBAsWkT/
z7buWhdOXPDOBbBakWxT2V21T6WsBL+D0H1vxv9kGcPWvpNgTgYAvOROwhQB+obzi/585tHwcB5L
S492Es6lj9cN5es9sKBXL45uVHXngKm4buos9j68IK/c93bwuS7w2gDG0HqjlJiSgPikYJRdC53i
VWDris9KGNKUT2WWw4CC3mvdMT8Lnm6PLTPvUxJV5QEUWF1NRFFoz2r4B1A5Tp/fP2xnLjiwfBey
WbqfhIq0e/+7iQ+dSeBrAV+z/2iuBVUYpCFdhbxBD86LV0mtjlHur+OWo1F6KEGpoEf7Pt1nFK1g
3RxoOtkmq4qR5q0hLTymz9IKnk/OwpJurFAvU1LHDE3uJFqtHA5oX4gzn5O2M1X8Z0IkglVtB9b2
F7zI9z8rQqO0K+TpRuhS9ujVi6rPJmDH88D1MyFIb3cViZbYY3D5rg+UfSWAkurAk2U2yKwUDNDo
MwuQWoLLnTL7ZJ1bZ5vV3YE3XpErPKoR+OkQA/0wuOC7rxrgUA7IYW6A2Z45JltI0dVyEPIZ8Uga
O9Nsc8Sr9xSwJ/vTe9yF87OhLrzQjPpmuzv7nHR3ZbXfJFl2RJG5TbzsWdgNr4a0eroXlczZxHWJ
rR0jNC/O+gJ6z57iCoCXX7GKazwBTxOLniZ/smjmzlZX45q5Iwr6a2VGSG/W9Jyuw9s/8o48HAoe
tXAnsurY6FAY5Sjy2yuodZXXkP1kVP4AS0MCIDxKTMGH8/NOH4QesREfJJ4a2lo+at34WjzF+K2Y
EFlzvtD0FpKX6v2ZrjJ4cyHRz12BWFsROuzuBPa7N2EaUXh1XJnkH3XTA8gTYwtYdsnm8ZXf7FOy
vhocOSMS0TVl5DAV+0uM0V7v5wXDHhqrnX8cg1Ocbr8qRNJNplQwRW7aoPjdr0izzJo6aLWUNWUl
j8dwCQoW2DbJA7597rMSMQhoxHpVN5eIJypIMpYK9WHos3f6ZyEmKfV8qiHQGLqacTkpH/uxIsIv
tfzenLzpLO2bdkANTn3T4l9HwJYwlcDZjUrNTJTCVWAD+eBQ4r5J0VbKRCcRZJeu/Pwjg6UmHKTb
3ah6DofBFg+GHS6BcE8hkq0JslBST6Jcgv4+mKsSQvL/HO6ZlCg/Qj1G5ga9o/jhnRiv5uNuT0XT
z2epLL7Ux1lI1c8t7aIVfthPIDRRcuM45zsnfQvIcJpfkfSU9yVAnV2E5DXhlmJBN1NOPnIr2mUV
u8cYHT+AY32P4GIaaLHh/M6oWphgtKlfH4L0mVmLgjS+DNwJcSXwqd8ginRYW3wnUIU176CZzQGo
u4vadxBwIEhaUCxLc4Y/U3a53tK/hi4WG1yvwL6SAJb2mIs7YhYohRVmb6nW+7BrVls71EivxR5y
wv5d4ag2pK51uwxp3tEVDx6HfUP/LAyXYpMSD/SJC3pYMVjJqxwqNBsKT9g3I1bdaxp8IXYvj7M/
10KX/2zT87yM0SkfQbVo8cf9yLSQO2x0TEiADiTwagpWj/WNDK4s6HgcoWCmKvnGS/nZvVf5QS05
56MjdPdRG/YmADbGCCH44T5iQs+6yTATnZuCn2wKtoRLWvYTC8nNEgDuZakHyhFT7qGBxlvlRHoW
9SCEwd3c1utE6JKzpqbXvg5kxKFE8OVXW+Gtctz2tekgbOuESMTyhPQM1Bu+bYWZm+3eZLONg7Ti
dsrHOGEVkjy/6eoYGKt2cNs/5C4eWp5ARs6y492bO5CqSHwUxSN2V4Ik2neIuf1Wt9B8v0ReKU8M
beKa1NaDY6pODMXPqhQZNFBHGZMa5VOdzzsOk8UjB0Vtirb5gquwjuvLzg9QgjCzlSf8uUCs2C/l
JoT67ytEil1gznQokD7KcZPdpXw+0v4EW/gAwYQj/JFOWPxkF/Mk9zqtSGj8pR3CYQg4QBuGwtSO
snoWwwf55ps5Ryx+M9qcFvl+lWiBjtoVpSIs8tPCTtYozHUMlIRDXRNkh1bxc1eG6B6upk5Xw3JX
CENwIl7xyCTgCp4wjJ4EW4eUDAB/JFV7Bcpp7ei1E5FNxQwc6kHV56xgJiMAale2SCM5tAKGfAO6
xdmP3HEEUhqOFnfzLlw4dl8aiR62kN3cx9/O+AvAjPIq8xD9a0f0WApZC3YIujcdoL4T5gWOH4Cz
DXTGO72IFywgapaHvSU6FW7rOd6+BikyRNa099jVOPyCxme4PPWbAHNvUfZGxhHP2FgQ0KfKrfQd
tPz9M8HfDFP8d8s+L1qezQhDX51/iw/TVRLXCxqEz2ZDvOi/EBZWMI27wSe/eJDno0mLRZvAlgeH
7VpPyl/yko8d1jv95d6NMCJd0EWK+/7Ye5JTF6yx3sX7KvSHX6kpdwP8Owb5hFBI1Z2FeClafsyE
cwH5/SpyVTWLgX7IZEggLqio/Cz8p4GA3fFOa0LFgLVhHLVlGoDNKD4SVBTTRjUY9KiHXrqWbsQl
/7Ejdr+RPe9ycHTWuS12fCb6A1wnFxDZyU5d0BQlD3xYwAceRQ5gQwUd+ObQluI1M5msDEsS0mGg
WvETFJuglwoGITNc0ELzcKJLAY7kJvNy2YIlH6aIvZPYKu8KAStP5ULs5Fp7bGeXDJKTAFecQgeX
M4YxOorlApgqGHfaSxtDGc5/UsRuv4JvM5tk5flPYK0lVqStLi6359ZVvxuuDKbIG58WvlofdX2V
+ZMqMTBD6VD5u6cA7yYAKuntkGdXVGbDTfx4b6/C2hsj/pUYzqgCptVOqdGhHqClHTRJKUNd4Q4s
1HLVIoWw2c/tr9C+JrWmRlMiV3GrIPA4VgYDUL86LkDDkqffmPtet2jdDw2p9AftpP7PYrOT9PgI
1/UPGLoor9grhL8q7YyW3o9PwtOED4YicbGSTqgj1hC5TPQsKAGdqu+5ziN5/KD7zo/PcJk2pk9C
TC1Uc7mOZSMGDyLaTv4jZJRJ214v3ZWMb1/Jt75pEcIKF1pBXNN9FWyY1IyeS+x/qUofrIZGnfEJ
h02NoxqExfeRqXg0kejZpMZrb4XKfNNtGEIPgL2356beZV96fZOg8VlkMn0EfUrCFe9ObxDMPHmo
iTXF7TP0JqOMPhSfrQrEHnC5YE2Ty/0+ebgRJDAZLnsPO/o4xDBH8INcz9eNEcfdPGbtTgLgjsRY
gkdzS48GOAPjX+LLLL9UeWURt05M03edFcjCvsl7NmrRKBYqMMsFIjFhx592QgtzMYad/pzw71ks
6rjVob9skiSbec/udBuNXtWT6iExhx63nq1ackpL/MTNbMObbtaOMnoZOhaftrytOaB+N+IbLgdO
pZR4/XBkyyCxlNMXZQ9KFNUk4/OId9g108yjqAMGOSeAIFUhMXYHO1zpuHPNknlhRBm/b44sV89B
KuKII7m4EJKJAiKuX370nkFReQKMoiqC6SPHTopjMy5xulY08NNqRQa/IQAa9Iy9JF73iRU1AlvA
fZxftO47CdOSqwYAcHufhQpo+5g9R7ooOZca2sLhkQN6pgx4PW0FLRYT7bbVigEcTVbEnRSpSEaH
tMLJLjB8adwdA+hfHYlPtIfTcb9XDpZZB/rWcgePxEXKLXPt3JdgTemb43DcKQt7tf9Di0AfJpJN
MUOaHo3BCX6rgwUFC0f6zMd/qUzN1C8P1FPkxPKlXUaxOzdzxZaxbb9AbHjqzZdt2kAX0sGumcgM
OYD3p9mYrIBAeoae4FW15jv3QIiDPlPMEvWTj9NlPavl48X8X0SCuAtCLVw7G9QpUYoafTfySDhM
/pTzCTaonIou300YAn2nQgtXoqWmWgsH09ZJ3d7xCQkyfsTghAvKQQLgkjEt1dUKT3uiIX67CF9m
ceyxrCoUPnSTc5UXb3rpqby0tpHxioXte5Y4PMw1puIMjBIjLG2toBC2WRQ/iJg9HSfhwEFXistg
jLOSytvBBUKTVMUjORuJ1RWAp0F1gD08UL3KUcbDfs2othuhuzYjQNU1jGEAN0ck3L31Ms2FKpo1
tJIw9pUwxPniP+uUZTwZi7nKZDo6b/byVCaqGo96s05a3vHw/V+Tt/wLvxo0oCKKshZlla5rywXM
2fOrafrqZ2pQa/lpRnCjBQqpbQbTyStd5som1ROcRRh7rq9yZg9kgOFj4x2xILIxwHSE3j5KhkP+
aaCFt8C3t4O1GTQZONw5TBTAfFrjX7RkOIlba0VuoeRIXTdUAfaSr3WGWbQ59OGvKaH6cGH+GdFC
iO0YAmHynMIz03xlDKybgtFVquPq50pBnTpl5kpKZDCYXbpQKxiSCannzsSnJrL444bhEnLNxzbB
IBDZS6hTFuUJ0U2XuPEGV10TxUhN63O5zStqvixjJEqirC4FaSpqJyvaZz6ZYj+DL6RNTUMCBA4I
ZPRHuWrxy0SPBBQyPatGBcSpO+xwLI7v7XYFachpP10FXBZG6jQnRYG3R0iozBfCCsptdOOIpYDK
qzZhnVBRsAxCAISZf5qQgfGNGEiVo41ZWBVq92vcOpiOwihz02MzEQUhmsLHXqa0GU/OWG62XB+7
zmPDvSJGbesv+lhQU9QMdsa5iYEltNWVamDDtROA6PDG+LJ9x8lBO/PWWPKELztldMmrZC/tCRQ+
Hb6yL3fvj824tlRggm0QK0lm+Qwtc1Xi22ZCJxpQXFi3kdlYFPT9gbjFBGZnh1Dg5uha1VtSbb+p
qL49JdXY5lYvITzTCpBSuCbUF5U+rd2VIX5Q01A2hxfKGYo6VK1EP5o+C8++xeKwtFAGZK5fhmJs
MXcqLr6vpXez2mt/fp50apyrGsK32fYMboYhRqCRIA/z7n+/2+ougACJot1EYKjxJo/h03uCUpZ1
8vrW19/Ws8qSUP77qTHTwvyJGZ+D5qhzHL3QRwYI7/eqtq/tzxj8xmzs1ZEHp8AFCsiSjI1Imjis
pjOBpNHtZ4tyhrAX1+DZjq7hy814Y+udo+Za+gf3VKfLRpqFWUa/WPGGzz/GhmlHQr80DpZUkJgB
6wZSUbtgghxAKscivSnco7clDanQ6rKHCjUJ58aZbsMeEr5XbKy+GA6VvH9X45NfTukNcvma8T7t
brxcq467WEU2SNTt+oWKV1neuxPq6bku9amjfERvkff8/iz8GH3Ixl6gRA1OWgHVmTdnmZ7oCPMl
+ean+xxqyxwIo8X2XwmKFZJHuTe0dC2su6v4KWw3ua+QEid/3GyL6b9WEMj7fx0tZQfjRcX2vkyd
dMuW0Y59BAuly19bu2IR8UKVDls2wyXLXFV9YRLXL/5Nd+0exVFZRq52hxpcEMxnvK1BNBUo9NaI
Vvy5/wEN0AGmMHhIg2lyGwKJ/hP6vaq9zGfjIoNYPKr7LoDzDTzsbAAKFkWBeqAKGLeucVaxlUHF
f6M+b9p3Ix0RlBWgz9bsOFuN+2krg3skHPZIkh68AgHeM2DK7MyFPgyQq0+1fTiHvkdgJbLUl1UR
Qf29JfIwN3qPRBJsZsGno2rd7np21ZfDKfAjrqwZkyOp3Uz2IUVCWKNE9GXPYk9U+V9V2laPKTdv
xGWOTPxc92zoYiF6k5eb/wozP95sJ2G/n0sClXtmMXJSRhvR+BFIJ0zqyiZGe9BPbOesRslZeVsb
Z8tLII16dYaDiJZas6JVMb+sp2l8Elu1ye8x5Yf/Z85Hlp5yzSQaAex5QD4vnflo4d7ydiLkyWun
w7JQuiI+5l034sObTExJmQ8ZQ3BeKVMQitMLiHfg93IOab7y9eI1M33kaHTbRo0cGgGkR/2TOWSC
snc6bpFSPFDzAW+3aqjWBcv7lcxjLXPQgqRPF3cmVrrJg12nEAPzcjoUeGzE9BigNwfavyKe7HME
vSV1Wb26+X0phmzK4RfamPUXTTH6pktFzWJ8wPRMU9KkceEyw96s9fsJ1L84N7wew/SHZC//r36v
+hMPmp8GEY+v39aD0gF6h2ypYBsd3LpXzqg8iW/WrT5TFPS94UvFN9V20RR7Lif57Yu+nPH5BxZA
SFdRRF3ToKGk7aOeZJSuZ+y68JSI3XJNaLS+lxwzENLawsMsx03xXS9SF8z1+p5TmaFvWj4qixCA
S8RXPhopO4aM/NZq6G4H1EBKYzABl/I81wzn/pxB4bw4Pq3tSWmrSuQO9PX9/qoY/gQD6Jgb+P3Q
h4oMw3KEUGWIV8tGxA+sLZJn4sbIDdNBZA/RihqgUV1+ZN4v6AtXNSR/MERZ3JNAeFjOPhWsKpDn
9PXO932k70j9baqeQxYT5gY5AvIJtEtkpqgnQmJ4QUgL63CFUiHvvqMq+cXLpLaRRHiowCiOvHyg
deA3Y8I2FRde7fbbw3t/YpL4bp/kJj6bR2g20n5qaSPvSMnQYN87bCCmSO8XvmkOwmZAQNB7NsDT
uOzchM4b96cGr1oiQO6T6MdhpuV8MYhW5sjivYA7Yx7Nx2yhWdPhsMh3mp/F/81NKt3GTy3wWPjZ
xTyhuNghp2n+yQmoyDiAnu6R9TwM0ng5sxnwAOj2p4GdadZ6Se2egzd+Ffqy75eSj5r/LETsBAq7
dJZRr39oT09xoG2jblGznr5lcT4jJeI/4vJE05iEDWRg/mwYyZXG6taI0+VjHrTce/3lkoesoQ2+
suh0IPhERBP4L/tVJ7vNXrrsktdkDIxSPxtHrDE/m4hiwt9V/hnMoPIXTtFVRCOmjVnyuiKBOeIT
Bdnlo78EbW82SGmUdCeSseGvbm8g7fPH6k2IRHjYFAIFiXCFS+KlefX9gv+w5+7ekb6209ulgc0h
hvROo5G5qg//kEfk/nH63ST9vAsMrnhMuis9adnS03z7fRWNJLFjDXwZgSmtl4JleZH47Vxh+GGM
lTtZoVVMq7mUmcewBzaeW54yj/h9njs/RZq7dTVRmguvP+b0Ni/42JiuYJpaOya0m+wsDJeNG9UG
V4i7azlJHREIFfLO2zfgSzxNSj9yw3WewqmVIJlWYzRisE4tl8DrN55GujVMKS/zvRIv5y29HBf2
vFMK4LbQlqPGkOGoUtHVe3OtFUxa4XM0ReJ0EbKppqICOEK70lDaD2cSnhRk+jY8iS2SkDjh4Wbk
/UDdd36gUKgRdbYS8mtidfgIl1eKErh1jTRImGwvS2j5uH18LvdcVmWgJArukMi4fqxiDifREPnG
Dd5MHIZHkiZoP6tyUxTHj+dDf0khQ2LLBP6QBcDdTcFvz8mcSFcBsGagInMuu2SDB6sQsu9ml8HL
dnLIOWn4HUFIe5n0Dw1g9IqFx+OV9zcLp0kFjROhc+iEMrefLiuGsEz5O/l5guuD4HTHu5FWvd5p
FDYcCcuETEPMD0T8EL9p9rnj4mFTns+DXZmE4JtGyqLaq6iSmShPXEWj9KEfycOKz4eckNBFrTF4
zQmL8FIkTqu/wSTFYgcU3SooTUhIt40JbFQ9JyM0scAck28R+aTwo7qO4kBf0h27ZL4MdHC503h1
ae6BebfFD/N6UtQMDStHhXJeXyJ9ackao0T9lTJOqevXxsBqQXoVmZPDyLis50w/tUYxvwou9Cz+
+/XzsUWvnsvLkPwUEdCfebIpB+c7jpWLDOG8RCfMq5ECtVrQrVfIWBDkfsOiR+EHZwFu6N3Uh7Fx
NUzYIz2k76bRQ/Gqmuv7Fkjy5YQAgNZyAZRi+kOMm1tXuzC1nSnWcvURblRoScTZ5qyWxq4UlS5N
5lwJjnqOEntGoUtuMS0HrTxjFUNxD6+FsCQ6hzpQRqH3zIAT5eCbgyQHAM681v9etkUfoQ+LSZwq
U4kdTEqmDCh32wmL0DzxYYfhYIIkj0hjkoOMjnpiQtJ0zPVvnJ8NE6QBV3Lq50dyjIiQF3KJIPQz
B2+jfvEGLWK9c3FpMh25q+jR2P6CoXeNJrhAabKUQEW2XHk30xe9dYw6LNgTUva0Y9Gi+odzcPtO
o3Y7oi3QexKV+nv1ppf8bLMtB68d2KTj28De2l/gA8Zxf5sRuidYz7+A6zUTIiVP12wTCSi6jX4O
pchm5XKrH/IYNjMiBWDT7hkNVcX1da5Ebu1DoaQb5cIV+tyCy2aUu+g5Qe5TJepA3jIHZo64sI8w
j2pPZQk+nj2bTP5WggY7q7lZAti1li5Gyrk4A/cTVbO3YxErY9dQpFFjUD9NQVmaOzo89yelLvdq
TsVMd8WGG3DHO2zn21J5s8fDeGZsOJumBDyesAoA0Viqf0lgHoQgzjcsE2ihQaCO+c/ZwCRDD8Qg
be2Av69Ug0D4zf6tw4MFwAAWjUS2EOUl/Ui+DMEMU39qWpRxfp3hpQ6PM7hChUgVGyBim7u8m5gY
B7OXnHO3W1HkqJTrfLiq23GZNSnQoEoCXQk92f+ntvgElolD8/P/pfv95yzccyLJ4xL2TicWvFDv
Nk6exchwh3rh30T3txFeXUeRpjATzojuqizbjWF4Ye+n8Pyz4EGhZ13diAwzv58su58CuHaR/2+8
zeo/6dpIeSW5X5oCC0rTT+/r8Ylu1yRtFcxmgJNwqTsnaDsEH/T1HxDpDDpZzLGt/03CC0dY95rH
VtKhR725enWRSK9kO7SdMyaZZXT78eJ0nfHhvBAjBSmoaw+eeqMEjVGI6EEaH1++uSifArUxnS/e
JiRQFbChuqbLbWq1cGRupPY5St9JuOqKRN/+va0Kwj1hrVGdPXhpSQnZvly1uAbHChcphZsGCb4V
FNGYzELLSMBdgg8LyhJkJvzXQ2KFbytb/NJMtdNYQCSOiSt/bxNts9Zcq27EgiIgjxEQUZzLnf0D
ssG+3PggRx02KpMpaqaN7sY84F67K6fwOb8GFD+C7hoc/IPmd/wUVoEzz0trprNUQmpO5jH/tk0Y
8DsqbIcPoKdsftPHqV/DWFRRuL3RiMxM6xCRXtlI48PF8AV1JUdjNVTfGN00X+MIs+Z0rT+MPFxg
KW0KbLiLggJr4ru76Fs2cbvNfEh89vVdxqJQ5xpLvRGr1dg4mgZv8nE2Ka7EREG+KOfNKyGNHg4p
RHWuPYMdS8JakY0kl2GRHdBchwkQEhNFXGGLGbQbN5i0ZRq/GezC3mDeWH4BdMhTeDQNq0X47oMB
aTXTZPtLPJ0YZFDyy2BHw7qrBDG0ELCi2KybrqO8oNBFuAVC/Mvjd7Cf3lURlH9/TVySANDjZIe5
6IhZ4/hxTqgyeuysP8YKKQHHudDR8oNWuIsIuL6/Ii4VJ/HKe9YL8gCyUpKBed9iBcBdUwTY9lTR
JVJ5Q10h3EXMAJp8i5I2/1RoiXEARMzVDAJ2jaHPsqqn7LICYiI5bBhBe37e8xEJ4Ef9UbuWtemL
DH9oEUp/VKJ2BP0E8B4q2ukjmIHf6zh5O/GhNx+DlfmMyZm8SssFNk99ZR1gLMDaTxYNqxt4susv
hAF/6zdeT9tBpDc912/3KvxH2lLgVdctdMkA5uXGAUJirFl2xPKqnoVmxVclIdtI4h1BOfEMaxt7
Nid+jIUU9yfY5iH27GEjc+TGMnDs3Fwf1krKKMTSN0I0b4SYXMeMZeR7RDG+xwgDmYDuRO3Ar5bx
XuYnHklf5xNnATXBbtBcFur486h6qJTZZRK+7OUfDyib0lwECHnpuxPKCH0qjs4vF4FTxbqjGCQZ
rH7RP5SiHN/P/hbebjqI8NZfhn0FlKUOxQnZc4o2IBjKfYd1ziR0QU7zCn4tTraU4eL0mvAYYkag
pRZH2QPoxajiizjfgkIvfUNi3Ji+G+dMoTT6JEyzOFoX4SurPBHIkCSkR5P2pzNwWpmcqvt3Uvrk
w9PBfxwVKmgHZG6E5nljm1IEti+nidSTfM5ziNgFsXHJN8wvbiQl/tejdWkpKwUvgijuumnwgMHO
Ig9aN1C5O5yJpam/Y6uX/gnwirYLHk9/KkAsCphYNArZi2aIQFBoZVVFTzCQT2P/CwvV+mCBsrfs
BkwNcEXsVpSnNWN7XHKrTkokVx9wXfb/5AtU8qZYw3zWzHeJ8MyWKcfTCvDWyPfsToHnpCEEjjUi
xdHUHTWuXDzDRH//v6tULPbwh1ttZnTOA2ZVQG8iGPu1j8/UV1+xFkbmiZ/5tStl9InsLNymjAve
w234uyDvLqisGyV/L8FsRDU5/9YeqLIaiZGyvERTsf21rK4lfry8eC9bNsO7hGNCVXFUxDJx/UL4
r5sGWCK+4klBwNaLse4nIhJneKHKh1lKS4yBkGwZJqUGQ0eQnaJkulN8GRXzH2seIULE6lXJN5oN
ml7d28iIpS6l8UTH2GvZuMp23WkRFabjSopkAl9sp8Mlc7kOyN3QRJkuPIeoJ48Gsh8BOqniN+uD
d/yiPaijcMwNrzUu6/JLWWDg019WWNsM80SJhFR5vqe1arm3Bzcc/w6UT8U3ohQiuaIYt3I2dnOT
wXrK9Z80URPnk89cWoHrWr0txwCdBsTlaWmUIVOz+xHMQF7+PqEEIEl5r+NkkXNHrwsDpTDibe2r
K6Noaw==
`protect end_protected
