XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��P&��}�l�I�o�_�d�]~ER�hC��b�a z䧒1;���O���kVK�T]�Wk���>ߖi�KRE��A�#/IlA�.	PV*��h���H� �#q��*��s/X�Ф/�2�iI��/��b2ۢ�FϹLe�1�L�`��~ByS	��i���>|�z|�=�m7�G�x��h"<� �R5�o�V�{r�H�ex)˨u�:��o$.X�/]�����v���k��9�����V�]Qr�z�~c�v�,,1�hx.�Ɨ�=vRUW3�s�I��y�m�`�L���#W���".��#��}���S�Ps��M�1co��U$�L�8�I�b:p�,9������ 9��=�Je��Sk��N� ���.ʀ}ڠ0�Ǿڕ��؂i�?��:��4O�[�b�L�:֚�����1��_�d���Qp�x�ٹ��Sysn���յ0���K������NVl�1�=c^�e�֯iehH��t&_]�p�՛Zq��y��\U�zZZ�ne}�8FoO�tF?lj�c��x@��e�����!��"�~ [�ƛ�y�����I�p��Q,Xy����fw4��q$��	ld�N���&a��IA���L����ڝ��1�^���xoz̋�3|�do�q�EԵW���ߍ�mc�E�c�F�b
��GO���=���D1�d]wYV�[E\��P�^��h��"-;Rb�% Jh3�oͬ�IU:�pn��-P�r���N6��ǹ��}�XlxVHYEB     400     190��8��6H�(و��ct��ܺ��I�&�3Yq���ӌ,Hm��|Z�#w���iy��(��{�
Ք۞\�v�Nn1v
�l�-�����QCq��[�H�|pd`�v��zګd�p;���g�`���e���{�C4�`�/�q�i�K)j{*Aq]�5��r�S�*i�H�^i�3�w������2^[������_6��v�+�Y�q_T�<�r�S�p�CF��4+�ZCp|!s���Y����P(�RlV�O�TE�vԙ+ॼ�U��Ă�Y�
�E�
�%�F��jN��I�C�0zE%Q��}]�N]�*�r�۲G}	dygGC�y5FN �D�Lsڗ2t'~�<�{��x�>Ԯ����lwg������l��Y���5��zj��ow�qXlxVHYEB     400     140fZ}��:�΀_%}�1�	�N�	)���������L���,����DY�X�;*\h�Լ�%ެ�?�p
gT����*灕�����2��ќ�5ݟ�?���`��;���w؜� ���:Q�Q,[�]hy��!��w���K2�.�-��VL���E$Io��U��J��I��߀)�˒ЂѰ~ޭ�W��f�y/�H$yB%�x�:q��5���y}���s&^�)��$ ��8/�kz�[��)ڰ��׿�os�T;|2�e�*�@�J��
��%��6"z6I����1�P8.+��U�&�������]Y�5W�f���XlxVHYEB     400     170�E"$�"���O�:	�{A�J�;�/����:a->�vP�-�)�M����k���x�_�f�ha�Rr'��s�"أ_�F�џ��}�O���w�O'��M�lT�Lp/أ�O�c�r>��x�}��;��:)ʷj�V���JhD瞣<�1T�g=gN ���? hսJ͞N/;�04?�;ǐ�tO��"�Ve�-�ʩ���]hq����L�F(���C�N?])�5�8����o�O#�h�b`c#=V�o�^�����)�([g�c�[L�/,qI�ɘ���xw�<�,��k�hE�޷�{]�5�"_Y}f��m�0=qc���	y89/�m���lbH���uyC��J�g�XlxVHYEB     400     130:���?��Y7�aRn~*�դm���F}�A�E��g��l����G6��ę�	��q�j�?��71g��/kٮ�����S�t{p�����@��Í�E�����ɜ;��]�2��s~������ѡL �l�58H%P�%��\�W#S 1\r% t��!A=��T�׶���x�5�&��|Z�"���p�]�4�fh:��.D�x���j�N��b��#�nhna� �=�1�cFH����n|�*H�%0b|��o������l�r�}��b��'�Uc\zh��Q�P[��2vXlxVHYEB     400      d0� ��)�X6��j*!n��r�/�U�d/����5��9�ﶻ�U�d�k��r��=p�*{�#�.]I4O<M���=Wlo,��Ne\�3}�q��X� s9��xT�JW[XЗ�S�y�5{O��d!ac�@��9����6�?�T���>ߢ�.����:�${ϵ:��A6���Ԣ��"8���t
h%��Q>Y/��_?�m�XlxVHYEB     400     130�� R|y����ܵ�5�V�Z!#�%,/uۦx*t��po��d��/e��{�����B�:*M�I�8Ь�u)��g|�QsjF��u���5�es�o2�F�C�+�킁NW�]��|O�_/�lD����:�L:�)q
�+�Z��NB}�"�q�#
(_*$Fg�/x��o�z�F��TMϦ��������'�5�a1w��tLL՜ߺ2���*룺�T0>\%����0�Ҥ�Lc�2�߁Hd���� �I:ȼr�U1�뿱)���K�pbZ�>E{���oF.GkH<-
��XlxVHYEB     400      e0;{Y�RݛY�Ec~���H*�K.`N-/n��3O�����"�y?v���$�.���Q��oJ����2د ��f�9���-����va���7���(��YF�E˯�*'�X�Y\���c`o��|�>�~�=�A5�(�g�Ŝ�:�n�nT EE�z��-�mV|ҝN]m�K���p=����)��QZ���n�R8���$I�55�$�-��XlxVHYEB     400     140�*���>BMՍ�|��S�+.JA��35���h$2��EW�	A��I,~�y��z��(��ֺ�+d���Zr0lw<8#�n	����Y\��wE�x:9��̋C�Թ�>~E�.��;D".��{����\Z:/�E	R|L��8��}rw��<�(/҈���B�����#�F�����f�A��Q��l?.X�A>���{:�<n���V���n+�?d�Ҡ��'�{E(7�e�k7�S>���~&���?K�O��!{Q� �i�`�ԮT�u=͘2�&��?t�6�N�88���i'�O`�Tu�UxX��Ta�XlxVHYEB     400     180��;}:��о�~�
���)�!����+^]L]���q�����Z{��T=�g��S����R���ljZ��c<n}HneJ֗��u䇔�'����]ԝV9���`aM��hI�7���"+.1�V�����EH���F�1�X��V����U��<g��䫇��iﭑ��1�;�zx5iu:M0��5��sL�p��-쵊�}�=!Ц?��I��r}�U���!#��A�'goXJ��(��zy�>�H��YRO��Z��t Pn��{ID6��&�C�Ψ#��9�6S�ȋ��w�.��mԒƪV�H���Q�Z%b&�
�\�{8�)fײ@@�HLg���u��6���g��N�O�Ƭ�k���U�
$�-&�[�}XlxVHYEB     400     150�6b֝O��"�d����[�b�҅d���+`�Ɵ�ˆ�W���̰{@�C�{�*���!��l�bځ��R1����/�/�弒6��E��/�{.��e��@h(�2E�O�3�#!Sa�Q"��	'������e�6��nm��"IK��@K`��B#7�Ő���n��|&R�c�G����"=��ЕN�F}p-�W]�^��L ��a='$���;�����)���e�'�1��f(�+�ל��Y�����|Nx5PD&B|�� 6u]E�ND?�v����S�9t7Jn�����~. ����˸j��}yӢ�?�âߝy������P$�XlxVHYEB     400     160.��=U�Ռr��{�[�����Ba[�s��'��"D�V�Ρ��I��O�G+��W��n7X��{�[��_W�$��`S:����}K�Q�*��Y`:}~�U�Z<|�XB=2W�|f��Q���x]"�d�㐽��0��|�{i�X[��͜0ۉ�K<�$��H`�N�n%0#���F �#�t�uj[swo����ue&�0xl����U)�f�S�V{����
F�1~�D+�ښ��*�v���h�G����0I���g4����0>��
��L�7����' �L��.�DF6PS@�D //�]�� >ۆ�~I��s��u*?��\e���*���q�8�]��0���DaXlxVHYEB     400     130�.��;�@n�m��N'JF��������� }l�
t����o�<����sU�)-��#vr��ڣ��Vg�ą����"%BQz�R���z�m�vWȷ����سa)�;������ Ph$q���p:�5�1H�Ѩ0�@-��l�߱ԭu����UΟ�+��T�,Re 22
�X)�[5��X�n�8
\�!�W71co $��^���鱃@T��LE�B�f[�mH�Fж�1>�bog�(YfoZ��(�-�M2������9F	���C��A룰�����_��n�XlxVHYEB     400     140s���ZQ�_�T'��{ӡ��ꓜ>=5���-�4k�8��Y���\��7��"�	�ƙÕ_i��dK� &_طd�lF�{G�K��	���K�q��M��8.��D��|����^���2�f��L�);��P��>��<ل/�F�W�������k �'q.rC ��_c��[;:mُmX�I>�p S,Xw�0�ZD�K���d �/��?���_?��XԾ๘;�x����]�
�s*;c��w:���066+��KN)4� ��Qp�M�#�Vzq�9���L�'���ո��)A�R�/����h�Rk8WE�v�XlxVHYEB     400     1a0B2����>�ǣw�J���a��I2��B��դ��P>ǈw�\��sN���:|v{��D�����|և�z}����Lf9��o�\�<S+b^�Uz�c)���Fm]�by�Ѣ�e��jD-��j�M��Hڊ:|Ҭ�ۗq�����~=�8W�W�㭷x�z�B,���2z�_z�5��7��<����;����>�3x��Y8�ƞ���ml�>�}]�#������+�ٲ����*�S0���}��ך6P�,8��"�=+���)��j)�i$�����C{�m~�k���b ����.��<���&�e�,:	�q����>�.�;��o��$���;�n�s��L�����76���-���1��$�޼�����s����`1���t�?��������XlxVHYEB     400     120 �nAU#k5	�F�;�Gx��n|��f�{��nߘ:*�"�9x���d4��~m�\�8Ѣ���m�h@�)f�$�	����>�v�s�Y>����%:x�*�4��:��4aS�b[qVo��(ې�(6�<��XG��wti�M��'F����i�֑���@n2�6	U>���P4��?)��[R;w�0�[�¿�i�AݨO|�E|5'^�F{Ux���>�0�>�n�9�A�00�.�e'�b�J��Q�moq?�n�:�C�܀,R�6�b����&d �XlxVHYEB     400     180�c�6�ϻ/D;Y��9̲Y
9I�r!������l�ݨ�s����gf9�����ip]�I�f���*���8�3�Rc7/=�я
���-%lH�v���
��OR�7���5����S��:[ÙӤ���aMf��fc54� ���wb����\2�17�%��	��H�gC,39�}��|��-�q^B�x�^�#ϼ�,3����Xvߙ*|9#0ŏ�J7P�QFy����eC�����n?��r~2A����{ٹ(�К����o3��Q+^@|�R i�e`�����g�$����ct$6JL��dt�C0��!_�0aL�7m�k�53G�
ӓ�w���X.f�������S���eiF�|3������>�XlxVHYEB     400     160+��ʚMO4�{R&6Ka����d�Jh�Q��P�vR�e�K�F��V�gN lݫN!���޾W͐;�����4�'��Jq&Ƀ�Ӓ����� !_{����yI���[��s��@�Y�ö�?S�K���z�w�:LDǠ,d��I��_�v�s��_m��Z�qԞ�sG>R���� 么�aަ�^l��Xʔz "�(RK��f��C/�۾Zb�q��he�V��5'�L�t��v4������e8�5��a����M9ca,sW�ڝH��-*�E�Qˍ����Q7�%���]ںK������K�����ق8���0��P�t��;�s}�7�}�1XlxVHYEB     400     1b0��(-7$�8X���0����T�0�1-��׹A� {�f4le��s�f�a�����گS���p�!�xP��2�s�%?u#�	���cv���d�8���_fԄT��	�ʩ�hr6'�"o�v�C����C�3���$�'��%r7��(�Y詓�B�Ac�'�o�BOC��$�c�Yh��s�g���u�A�h\V�W���e�j7���G�Z<�k]=˧��\ m�.eȠLR�Ŗ2�!���\�n��*����^U��:�/�A�n����Q���)��m�i� g����ǝ��b�Sa��f�#k�e�T;�R��gJ'Z�)bh��	�M����"p��k[��[	�Zcm����)�j+J�q����Ձ�I�,)��zdMD�e���'J�-�D���H}U��T^+�BgU_��)�I2n��b�XlxVHYEB     400     160KMlJ`�A9���>r��x�� =�����[�%c��>mjg�-�D�������q)����R���o���62xҧ2��;���A.yȼ�������n��\~��J{��Oi�7��?�Ro�ov�g�����HF�����������,�`��G�ftb��'c�DS=qc M�9B��H�5�U���te�.�6j�?ךm����a\�<�>���ݘ=��$�񵹊g�3`E���ER��,��|�Y�׋*f4@�ԁ�_I��x{�~#�-��\ Eη�����a�U���PTm.�yҲ�o�g6�y�{�-�nټ�����4"�7@P�@���:/<��Om�2��XlxVHYEB     400     130�6�V�m�R��?���ݚ�92���E��ok����8a-�On0��.�1Ԧ�{��F.�I�-#65c�+�s}�f�Ғ_��zm��Ϳ|��ٕ�7[۱p�l^b�pM�'�j�㽡PTPc���.��ɝ���ԓ�Ʀ8��/�3���-��[�y��`�+��e���L�	G7��L�h� 
_�4��#���U�#OBE�1�U]�wv��B�_�w2;GEɃ��+�.Rq�����gԻpf
;�'f�uQY����Z!
<�;��V�e\Y�ďN��\U�xynH��U�ˢ��i��xP{��XlxVHYEB     400     140�
�y&C�D�p`���Ϟ���;Y^�呌�/ �7�C3t�������h�K�2�~�����o�oL:#
$���Л���|�o���X94T��xi˾	#�{�H8�d�FGI�W�ͨU�򋫂߸ͮ2IjbRmҙ�c$+_�:yс |���	��U�a���y��Z�c�;D�\yo�ؤt�s���M�q�xU���&;��1`y�G�`�ũ�2�UNa�_ˌ�?xo	���9rY��u#jq3���.�"\�tw�,�9���N�R/���SԔ��X��%�?�V�lmm�c7p���Ṛq�Cԓ4	��XlxVHYEB     400     130i*N�'qء���x�7Zx�om0<W.�5�3Px�� �i�`��U{tT�дZ��gA��i��r���VO�(֗�@���X��h�v#�k�|��sT�!��z��s�q�>��ƻ�櫑/aCE��ja���HB��d����WlDYp�yX2/�2�x
K��q~
a��/�,��*m酬In���Ɨ���؃e��ڂS�7�(��/�I�|I��f�S��Ls�AY5��\��0.cѤӁ��ㆼDA�X�n�d,%*8�����ǒ~ omܙZE��?XA� !��hT��?�XlxVHYEB     400     140�i
�Y�!��S��w�� ��[W9�P���YqH�d����W\��*�+����LWb|��d�ܮ29���n�/�����i��,���^D1]����A��P���&GSIÆ���9b���lt�g���s���ș��o��I\�{����#j�$�k .�_͂'&��a,�&M�_Q�Wr���2�+�g�>V��mMgֆ�,Ճ�G�G��6!v�}�����q� �w�F�y0�
���co�3"F���������=�7f��ln9s�z��eؔ>FT=)����ׅ������c�2_�����
���q��}a
����nGXlxVHYEB     400      d0�I�i��F�Է�Z��J���m�2�}�d]v�!@�0��$)�q�:�洲4F��Va�]�!G���Z�"�m��W�.�j?�Q@^"B$��d�S�1�3<f���(�S�;�l �N�c��+�C���x�䴗�L̐䏦���4	�m�e��4n<��C��QAYS-�����M˥vJ����'��K֓�џ�W�իۯXlxVHYEB     247      b0Q�>������  =�(:�t��f�\%��5B/R�*��m��1�jKs��>�\�Ɛ�m N$�����}��&���w¥��u�<XC��>��@�Iܬ>�z6�q	���a���#�H¸1]�Ώ�i38¾.y��煮w�����ۡ\طK'�b&!��'�E�Dǆ