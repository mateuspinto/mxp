XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��;Ȋc��P�dEM�ȭ�{�>�a���'�gQ�j�tM��NM��Jr��t&?9*����b�D��N�i��瀴�3)����`��"������n�U�W$����;�^h�&~�L2b�w�	��c���y	�r~�$-'"Ct/nH4�KK�`n��K���.�]ڡ�\X��Ï�'Z�-�]���^X3Q�����hd'��G/Լï�Xɲ�5^	�Z��q��� z�q�<[/��}Ju J)O!w9~
��E�5��8��v_ZM�;�nla�n�
q��Ay�;�W*�g��*
��DݛGҢ����<x�
?���<)~�6*���`���r�}^U̱�P[��68;]ߌ��Y�R�$뵉���N�ub�9���TZ���-�G�3
$��,�h+����Z�a�U,6x�o�M��s?椥G���Z��W��nFҏ2�I	j��^*F����i��{�2M-L_�������bl��f�.��U��I��S�,��tݭ4�hư�+�N������x���]$�Uɡӣ�Qfks�1���Xq�i����� �>J ��E��l�2C1�&���Q�e����My��Ql����1�oc�Sug���ܾu~�Hͦcڕǃw|lf �������nıH�H���q-�.Ƥ5~�==Ǩ��L���	x.��x�P���a����B%�`F��0Ne�0���pm``� ��PEk����_�#)K� �T��DZ��"��XlxVHYEB     400     190e(��4�@����`Z�U(��b�I���N,�K�wv�����)}m�u(�_�"��K��2.k�
��E�1p">�)9�����FSO��Y�q��ꝗ'R{�J;8UA����Əzf'>_r����4��7�: ���%�5f���g����m��2��uY�����������n�#����Ub	;��,CFU��^V�"q�*i�9C�/_Ih�v�Qʯ�T��yT�u�ͫ�d��Z�)D��l~�����X}������k��2.xO�4��R�?�tY ����a�5�Y4�uQt�u�.{4A�o9@��Q��-ߖ^>]Q8��:�x}��>��m�'Z%��b� ª� b��)-��aH"���JP2ؐY�I�y/�<ɨ2<�1 �XlxVHYEB     400     1f0�+����!3HáF���6�������m�1��7�(i�mR�u,[GO�w�˰�{�p�����8�P��7�(�>�*��!�Ԡu�ӄ-��o���)P(��sD�Q϶16!u���'����Uz *lU������c!��\� �X����̠�)D��w��dX�9t�	����7y~RWusEL���y�y�E�66�t�����^���1\4��w�<40Y#���j�'W6�*�F��)qa3òٕ��\uƂ^4c~��rԞ�i`EQ�S����Ĵ0Y�xe�U�a0�dS�X�;�Z/	�EM"���!`,���(�*��@�O���<g
'�ءT�'�f�@ؠe���?�g
%t���gP;$X�{*l���/
�~&���
҈ ���of�=��y)&P^Cv�+8`����ȿr!za��9q~W
�-��+�L]R3�B�'�ǽ��<����?��ِ'�ٷ5M���̢d�"��g�XlxVHYEB     400     200���p'8�i}�5�m�.�S�e!�����T�%g�:)l)���6+�_l�ߋx�ܞk��"�§_���`��mP�����1��7bJN��;Ps���K�F��r�}W��)���q�q'���oQv����Gb�󄑬�c�ɖ�̡�"�`�-�	yd�,�w��pp�����CK^�"�$'�������I�+Ӏ~��瀇� �c!���8�����'1��cS-`�Ea�^��n�J�j:x@.�e�-���] ��t����\!/�fmX��H��c��s����4�	N	�[=n&����"������s�X��oo�h��3h��LXɵ�v����f�C��Ȉf��|�%����� q��/<Y-Κ��KgҪ�tG�+!L�"^��w4�gY�
��=���x�R��;�U`�7�Hh���4�}��v��3I��lʱ{�=�$&H�ƭ{��8�q��bM�!��;l�^�t���!":�6���L\P���׳XlxVHYEB     197      f0O���E�f�ЍՀ�,��`h�V�mg�v�/�������?S����[�Np�2g��(н 7�q31��I,��:��� �k�����Li�0�hi�W!���cp ��D�l�	�fgg���&��Nl����X������
N�vU�)C��U?��}���W��]&��syh��RQ�|x�����/^A�4��U���ޅ䔂t�Q03r+�

[A�~����pL�qv��zڭ�׫�F��pVL�