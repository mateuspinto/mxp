��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���mQ� ^$�k��Z�.d�/�1�<�3h)�W3
�v��Or�U�Q��u��A�z"|l�,�T[��i���������<�{˄�	}��TL ����퍢�� vk���f�,20g�|>S2�rR�\��Df
�F�{�4;$(�����΢����^����s�-�eA�ƺ��	���QܙIogV�����aFy�-ʐ�o�;z��@�C0e��k ���w5�3�Q�l E}/FO�n�$��di����@�^W�(��+�[�Yѹf@��a@�>W�o�	J��$U��� 7�!���:���j1���Br�7���#\IICB�D'���x�ޯ~
��ƽ��0�ϋ%u��C�����$����%A�LW���}�
�U��Ԭ��0���˕�v!9�v*9��\&%�eC&/��2>��<.���Pw��Z4[o��D��}�N�U/./1|&Wb b{�v�����H�p���h�(�M� ��QV���?�����mǹ��N���Wy�Y3��I�@B�D���b�W3% Ī����!�L��J�<�In����;�i���b� �`gk���;�3�J�9��bzo��JK�4�o=8� �T,=�-�:�Oh�7Q��/�T��ܕ�f�l!J�N���M��LJ��O��2%��C��-����4-����12�'�����u��.�8����]���=��w�XZ:�(����p�\I�"�>�Z5�'��2����!�h�D�m�AZs�iu��k�pҥL�%��pA��l�x�s���.RO`Em��9e~��,)1kt�'�` <�&�[�=᳚��c�{�!�+ji�Әi�K6�Dϓ*�ݜ�F���4�e�=��C$�/�����f6G>���4�zrQ�����,��c4I�uC�MA��>u�h
�JX�S�v��}�EOw>�@J��%��ONؔ�յ7�L�t������~�'�[��<���p�_��b�
�n ��c�A�_ B�j��:���G���yq?tE]��ou\7�t��#b�(�m ͕.`�wAk��Xe��Zc4�n9.d��������Κ����L�����zR0X�
��/'���ǳ?��ߨ���fhӯ.X�c��A�R�Y��Hw�Z�Y����|���y����o�	�lƧG���c�;��i+�@��+�f�����!D�/x���g1���(�����M��z(�mb�u��=t#a�
4"uZ�ug�`
!Za�����8�Ӡ�7N&{.8�t�;t���ޙ����)��>Wu����j;Q��,�k���|T;W9M���^��X��/U���P��h#�0�C��Na��y��~��@�E�b�md}��	�>%D���I_T�|Vt|�[g.%w/t��F��i�κ֡�����͋/4�%�&��H���a������p/#b�;�̂V�϶���tC�"��o��Tҝ�/�ԅ�v� ^������NgJ4�ZaO!^�:���2��Mj���Wϼ7=s ��"ڞ^��t�kL�b:Uz#�N���J0��ݔ>�\��2��1�^K��K��,J�fV����g g(Ӧ
F��X��)�����ƩT���T"9��t�$i�y.ÿ}5!c��I<e�|�[���[��j+�5H߂s�3��j�پ\C�[3,͵�sJ���y�}4�΍9w�O�юazΆ[;mY�Y���k�� ��EY�8��K{�D� 0�<h���r[1�!e�V+e��B����x��usgc�'����7�J��+���z�;Vv�K`�z���떑��
�G�?�������7��<@IO�;$rG��|��+y��I�)k�����pt`*BS������_�hV�_����Ӏg��Är|t�d`����p|yPdi٘Ķ=��֛[�2 k�ܗ�����&�,�4"���.��n��i�