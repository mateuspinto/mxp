`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3168)
`protect data_block
ELYIPNkxxYlmBG8acOJvlfwSZIwRo6qB+41yEzMgZo6UTqhI3apAdWVYuM1tEVKWKoYOoHWMKVYz
e9SKUB3l8w6OWcelwDZPjMmXYb1SOnl8P+K12MIycXaLLhMDsq9whIotDePHwJcg1X5KtX5j2tvP
+kvc84LsdY3QphFdw9ldhzHMrtj5xY7cPrsQnfigSBwhOr8/gnlt623yPQqTa62W7qgAvgI80rhE
veALlJNlVo5B9ZymtEXdcij8VIXSKKToZgKSWWkJXdr+pzUwxjgPbYj9GBBfpE1tWypA8wvv34yP
B3eT+u5ANAxbs4YMdwvZG8ezK20dXQuNsGm4Opur26YGa+yo8ru5MQURTeoN/QIpxQfDgEqmFTQS
vTR8yhMOxzkfgjBKz//AuWgR7jeHNVzf8kbdQZZbMBBLrn24MaVRvub0bJmgvCREhXsA8n11PlxE
6cmW+dVWuHKAaqcqNngwWf8JGimSOSQop8hACI38kJta9hPIZZM9YgMmbt+fwmgymnLpZeVP9MbV
8fqXZzbtkvgwMQLXLammVUohNEtI1jPBz6c9CESn0Zvu7DY4b3DZAfdBbG1G7laWQU57fN9SGMGe
nZ+BB9g2lbycsEryZaWzZfgAWNNDA5rQlY36/YU+r3tlw2ksc8cYbUZap3JOCKQuMGbyYemQ0k0s
C1gooK0Xxzuc5egnUcm4yQO8QveBppZu9u9mp4CaCoMrOn6jqIgg5G5RPKXIdf2cwhRtBdH/fHh4
EKfRlrmdIHT+95gpsQ5yZ+JAua7PIfotgTWWsur52LqIzZAm32TV6nAZp5xHX7QCNYtEc0zUbjYD
GO/PLL32GTO39fTahXxpD4RsoPr4OyXdWmSC1VQLTIL5FGp2wwSVGSJUQHiHAJDZBJk2jrusXGmf
QsCb2FABkHtf9dbck9FiQDNauk5JfkkPXV/Vnuftr4oPE8qmXAIgU0/lp2yYShJtBonr/HH/v7Hj
+JUbUC7KkGfuEP+pe0zXIneN9vaO3bqEG/pf5hLffeAXGMt824//nUN1TqWchGGp97NURMfpdlVH
HdF2i0HYi7oeuDy9yhbhYYTvgoNWtywHF15TMDp1mPaMlWwRJuUYRBVGSg5iKWU/qWe4BByQ7Zov
crC+JKjf3cuovnkypOANgB7jO78aQYIDyhCUKu/r5ZT7FSC1EobsNdtuInqVGkr3b1u0XcnAFUw3
GkdoR8MqXvpl1qojYexlKe2ky72gGckCeq5+9zwubO6Er7avsrOL7W5cDGTPcCCn+JMBDwGAY7lF
GJ+/KbWEGnkSMFevjrpe1te13OqcMCm/DIvBhT6sp1e5LDJIULAEOmRfceRe7TwjIka7J7xtmajl
mCsiErIT+/OefnjycJ2c0yIVTKMxA6fP7Gonqy7livSw6HO8q2Sdm6LNc1bd/lvuxYbgMzWaqNx/
M7a7PBmr/+d8UZefUP7lIM6uNVaIY0ziDzRqq23NVLY4WQ2xUVFTpSeer3UotlYcXZrE45msSN1E
C/boBAujVfbdmNEK7NtXVfsUjdCBz2LmhwuSC0TROCMm0QP683KSWhZgQ7cLEnV20PljfaVvoy+D
TIcTrCbA/T933q82fyCP/4bpjzga5og0eSvenQzZ+bi2lE48F644USdTlCQCb/dIC0F14oM9YoTP
kMbHtvrcXDWUTX3be53rceQoMXrZqW7CPoYOLQ4T3ZUjhyar7Rgd/R4GBb2EA+MZDBDKZwdaB30G
VHzwjVKonbpbTiGq9ui7QJt2FW394oLFpvenFeRh6mwZriTX985mGXOVYSEQH2nzjYxR2r4FJ0pb
JVT2DcDCfbxW3r4uPFF5HBXF+j98t+YU9i2GTd87ogmcBdD2ziRDGI7O7Vi73wQjRSgl3OFFB9Ku
KZkfgt43p0GJu6rk6hrXZYDSGABOXPf1+7Q0tBF0YaEVogRPH0dHZFyQ+hZfGvGiQLepfgcgNfjY
1/Mrm1H+FgCQDp8IViIdPwkgL1HZooy44hPWyIcC24ZyZ8dtLXQpsZHaKMhCNfshsbsIUxpP0I9c
7rPK9oB7pMEyDkA8UAy4vxkUMo3m/TQmJFe5piKaH1ncIAZbgj5ukhsypOKLbA1Iy80Fplnnzg5I
wfcInqebXJuioCpncgq/S30i8mVET9UM+GkZjGix7BCKAO1Sj4KPhVlrhzflzGb1Vet0DBAJiWZj
ZMaPWmV9bkw0shMwd/yUPecew8OSKZ+1IBrWMFmqvjtSjIF22mQfHgOI2SgvOXIsiIakqn/olmPT
Khsu97MAesiSJh4BtoSgxzEvnlsjER2wrSYQiVkC6wHRrAD4EpoKO46iGvd+FwkRWZbEVX1yN7aC
IZApCwDUhqKTELSk53GyDD8qDiyRAwCyHL5+Y8Zi2Hx1TLavfk5E/4f9jP4yjpeqBBvleNY/JsY3
t8mk6/YBzZ54s/khjWZgaQuazWaQqVdfQ+EbNvGEaWqaBfMUWBrIJHWwrE7QjyTREQDnNI6Z6y1K
twtLcljcEfJYX00WhQKEEXgRrxaZe6dNFvb3wUeCnVlEchmZdsadCN7xvVGBPzBtDWZyp/jbJBZ6
1u2l7MDPtuPorVCRLghtntp+ARu2dRW0u3V5+2KCj4FaIzH7lLJo6iDVUGHCxn2mdkaGCSP2XRlD
wgDLznQ/KZFcE43FS/025IvhAq+OnSFpvTrfChshEZXkLApgbUcwQXMUNNANs/7RSFrmg32HUkzx
VHK+qwubba1ofdJFdRrUcKgZgJxVSPWAgAmyelQRjv7HlEb7vDy06vKEcM22AXHVLSqr+ivOju95
yihf6Y2Mbac1dJeMVDjQTglc/uE/2NFiCzemsSYcG0x0xfvIfa81GvY/+TjGLzWvlIFuTrsm3QzT
HFzM/C+gl2E/R60ZG5CU3wE3eRlXTK5TyXik1+nkpmSrOKoenQ9cXKyaosiDVAYh2XYCMqYq0qbr
R8LjwXq14mEazXAEXoBVxRdnD0+xZGZApKYRUv7UhwXrrQ31X0Zm3uy1Tx5wYgagAkzE9Fk1jwlK
KKtVSqstIfhzlep7SkgjouDooAQtJBlK7JwYAd1/1vzB6guBtYjgxdIpRDnl/ZL1O0jqeiqUkPy2
uB7kiWiUAFdFGKJKKfcc8c0KUPoZsQZWDfcOuFeIzgqrG5wm5BAvWxaPHNBwWOP+mI1JTZ/6/Tzd
bSFeYTu2IVLi+tugnkFw74EYQGXhE6QLIktYHXetRm/6K/yRHMiOWS6MU8GBhDbIBar+UdGCrUhF
j8lszOOjauO/rFo5kVcybZHrCP7IFVhzPboHd3gs7NGWBGJtF6MBZyfN8rxqTAJB1K6E2wCXA7Yy
GtI7jfRgT0fd6yznLXL9dWaX5+VhfxoSz+dzrp4P2pVCsCCFoEKH2HHRe1yrAB/nqmZe5MV2JIxt
5aU8160fIHFy84zIgSQoS17y+Z9Cv8kxu31IKFowWXleeYGIXbCQ+eomCjELCqjPYdnBql8PISUv
ipiHSovuBecNwtea/OMQ9Q3Dg0JLvjC7c2YelQZugG9BMCQ6kbxuW1YLBnhbzok7IqhxxWH5k6Dk
0nA6Tw9vWAbhVN5iDqsj2Xk7aUyqycBfYN9PdBNwtBVsh0/9kaj57FX3nKeZ1GHa8d4UOC9qFDI/
kdfmdImMCN76zA8JX91p0hSe77T3ZgnEx5S4tXDRmwUxZuFeMpWmga2IAKC0kRcY+jv5UJ4NyG4z
2WxfONsc9EkV1UXy6s6TQJJmtax/h0056lpEg03fJS7GTodUAysWY9Bebo4fuJgAja3bW4B0zEim
R1MJ3f4b0M0TZ0q2MMbiC0jai64tWsZ5JqkbJsrzwYPuz5QsC4yagpjgdhzJWhBT2Gqp4CI2IFYw
OlWwFE8JzJnCZS9cvQqiBjE5L08Gpf15o3op/odTwyRYvfUoJ1ZhJkf47q1iDsTyfbeMBCsKudcu
3oy2/gCDc5e8/clNEo9s63Ilkwiaugf8MPsvvsWn/xArk8i5J6h3459C3GMILLZ5nrCLwGOSHn1C
BBNvjmMOdv8qxCjaSZbw7fzHd/CZ1Nu+TagEEC/+Mi3m3lHzgiY37FuTtUzaIUWdGyZrO0N2oDRv
T49AZ8cQTwMe8GI2Z/wKfrOq1bdKDe9e3YIlZRI6WLRSUX/F4gskOKLWSG3W4LxnpwSq5pazL5qp
UfC/X/Bk4uDmHthJZsesDQKyG65/xGvODNa3tHghhzo9
`protect end_protected
