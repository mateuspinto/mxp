XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��{C��M�~��	�'n��z��c�]�7fԑK�}j'���vu�����v]0 �>��p���$W��LN�(�_�D��∁�N.��@o��'��S��bu��^1��X�$���0�
�8QXzA��A�׾�9�c\0a�.2�V0���c���������;,��г�|�hzI�EuwZ�oH��l��`���QQ��mg�{�K���N�1vބ׃9Tд3�Ql0�pd�ï#��*���'܀ur3hi���'qM.�4
2���_bA�VC�/݁�p��	�8�\�g�#"�ރ'���1mg�\��E$\w��xƈM׭.mJ�-��;��3ܵ�Ȥ]|Z@���QНHH,�^���^�kO�-��#�Y�u
���A=�^{��xt�?Lj�G�)��m��,�����)����
	�wG�A��2Qp6�)RF��ӷ�9NS.OKN��P=��[y���.�KOQz-PJﻨ��*��LN���J�[�R0�jb�-��E�I-��{!��,���l���bn/�p{�t�г�dكk�[$�L��"�)=Z����
3Ā!8x�m�l�o�K�VY����)�c�� ߏ�;����Z/P�Q,igʟe��I�u[�Ő"�mˢ�\�����.�Q�P鶵��k�-��<x�tB��w�$�r�ϛ<HN��xu9��[o�D9��^�TQVvy�����)K>mOp�[��ȃ�|1�{K���D�Z%k�2��Bo;�
D?z�qYѬ�B��.,���	XlxVHYEB     400     1e0�'��78{���\�T��@���	�d�乕�˦�e���u��4��)s��haȓ!�ֳ��洟!�&J��R�8d�\�O�?�B6fs�M�W�z�����&<5� /+��=%1P@ܰP��5��@C<���~��m]�jw�����]nڰ3�����Y������HYmn�Zn=�eO;��2���J:d��!fffO�0�}}IAiζ=��k�*�����j?x!7Vg�ī1H���	SB5�<.�3C sn�Km����Vg�pyॄ�s'E��{�#��Wa����$�~
b�c���v�]3#h�' R�����X�S�������͡n��*^��p�z�����P���)�r�(�t�#��?�>+�v.� z��̓��M\Kʮj�b�R��!XI<WqI�{�����-S{��cA��G�[���٥��0��rܰ��`��'XH4!_���q�����}Z펯XlxVHYEB     400     1a0~�<�
p�9*d*�'������ku9�ÒlL���HB�?H��e�?��e��L� ���R��ؕp���#�*��$�~~8�o`RBx�.�m�d������_L�Xq�o9×cQY��3�{�x8�x9�"s,�cxdl�[�R�u�z����;������`Ѭ	9��+7����M�̦f�0ɂ��*�ϫ�EZ~�4E[M/^����A@6�{R���ĳ� �ד��0V:��4��[N_Z�)��!v �!&F!���c�cn������������~5��JZ�� ���j}�/��Iű��佝��s2�S��#X�>�jp��s�d��ׯ1�H߁�	��H�<�h�C:�����%n� ��Y��&I�r���8B�:س��v�Ii�l0���m~[�	c�t-�KXlxVHYEB     400     130!�1��k��ˑ�Q�$��2�H��^���1���a���X"��\G�D%�<��)Hjwy��L����6��2�=5���g榽+�����	��G�ђ�`���W�!j����1=�`�S,�KW9�7L��tR(��ֽ��_�A���=�-�Gg��6�e��^�A���%�`l4�33���Jb,�L�=ݻ��yJ����>�>�\Feս�����w�]~فA�.1������ZZB�x�_B9_����d �2 X����'(4�*�e��OlA��+C4o�NU�7UXlxVHYEB     400     150�6I�뤛zJeQ��3��x�g�&��/���B�1\ rT{���H$P�z"aWq��*VMiIא>�6��Vڳ�����B�������ѱ�ڊ%�7Nz2�k[!�//��*�&�C�G��8z���Q�9�Z!���L"�Bκ�����$qT���s�q�o�������럴������/ �vީ{d��\�o��;��k���ǼL>�\CM2%��8�C]�Qr�}r9�5�g8g$�"c����>�$���ر�^KB52��܎I�����^���������+b�!\=�~l�*&���|ux3���S�p�f�U�`���n�X���&z�+&xQ)!XlxVHYEB     400     1a0G�=�)i��⤑�OӐ��rβ�������;�3��kse!�\���w�'L_��3%�w[1*<���X�x`�ܻw��u�6���#+�X�c�ޢa:Ȑ:���<\��s��Ǝ=��q���pCy�jG;$G���g��V*z![Ͷ�e���-��S�dn���&Wu�K(/��K�g0�\��S.���v�}��5�q�ћ�st��i�@�||���z(ʦ��q���4սn��!Q�Z��ȁw�p
Љ5�0L6qƀ"�3�Ϻy�!!�B#����#I�� W%��dZj��C)A&�ͳP\� ur�LJJt�����92B��Rd�h�ʪ�~`9�6:=0���`v&�����i��}\�6S� ��(
kqC�}�Nߝ���怖�U��؜ ���8N�tL��T��AXlxVHYEB     400     180F_w�(�N_�N����n}iI�{.�%1A�����/�������
��c��ܧ	g��'����(����Mڣ�]�L�g<*��uf��.��lR  q���8��9Md>�;�2Y#��uڴʒ�ϰ��6�Y�����	x���p����c2�8[�p��6�C��R����m#>���dy�`С��Q��G�p�ef��+��'��[~�c,�[VWw]���=]̼z��2�8X�c&w��"�CL�Ԟ��[�(f�s�-RƝ��\o�R��u�)��f�ڧ=�~�~K�J]}���qO���I���X������d9�&"��Yza����s�=��c1&�s���s�xY�+I8+���,n�16���8�z >XlxVHYEB     3a0     170��R 9�}������We��Z� �$��w9�쏖��\�A�*�;�%҄���H
��-���)Ҋ'�E��l*A�K%����n���$tAƿ�V����	G= ����眹]�K5*w<tSB/I����5.K�D��a�=��aH�R���{��I�'���:AԬ����C5�%��Tn��n�-S���4�HL�?���i�v�U"+�_[g���R���̅1)!��`��@ �3��u����PDǪl_��:;�V�90����#�ӿx<~��/avdi]��R�d�u��?�H��N�h����`.:�e�~�7�ȣ���5'����V'��v��D�Q7L�����$AL8�j�>���M��