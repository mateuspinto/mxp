XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���	�ֿ��c��U��bx�L}V����f�hϤ[�T��${rS\ ���u�Ibi@;@����H�kU��-���`KayG4	<p�DJeWa�]>"_V���H[��s�7o5�57u57b%�
���C1���g3ًq�>�awy��qf>�{+2�D�wW�Y�z<�~Ks�!��T_���+�e�5�	�0�fA���1�SWg;�5�_�O�r�ؼ�H5�ؕ���2p�?:E娫5=_^T��=ɔ��@ �e�$W�g#f�u�J֝g��$�R�ۤopY^���4��X����F��ı��-�@6�{�{����3c$��Tu�I~���T���u4���/o���!��!��=<ɿ�݈�
�/�H��s������e�����G�<���nW;ȋs�{O%��ٽ��z�'��|�B��7�>��{�(�*aw��~��ڡ?ڵ�;fH;K7�t�u�0��=ߊf���Ŭ�G��Sk�lu7�L�|}sk��Z��\',��~�pl0)�
:;F$�+!6q`���κ*vkL��Ic'�t���_{������KV�ĭ�E���Y/}�a9Rat�o�ي��"�U�~���V~�E~�J�޼x7JH��1�ʌwda��u�q�=�[KEz����R*P��jlKs�H]2����/���?Ms�$>��2���0�����_ww	����%���5,���q������iI������~f�`���p�O�x1�����ʋfdl�k���XlxVHYEB     400     220M��CI���e�T����u��'�N���*���ԕS��Z5�����R�F�������DZ���m
;(�ϜN^F=Aп	��	�l^�۸>�=&�Z����@vX���D�p� [���*{1?$��T ⇵�ΨG
~�A�����W�45��.Ĭ[��gg%*ji��q\;i��Q��v?vwhi�N�����h�\�����u�A5�d��MN��̂���{*��wl��6�k��,���{\�鞞��<��5W�0��gg@*��T�����KE��YW�]���j
�|����T���;�K�xRt���}�0"��cnq�����ڟQM�d�Y�mv���W�I�9����KM�Z�����Ҫ_�MAq�-m�Q�AmR�[!�B�[���H"6woZ�6�=�)5$��l)���U�
�2d�_�$n�����z�!�=�I�5�lX�3��r�PJ���{Yt<j�Ɂ��N�I+��s���rM3�������>e��5�Q7b�%Q*��?$u�A)(&�C��3R������;1�s�}=�:]!XlxVHYEB     400     220$� ��_�T�w{PPs�{xdD�b�{��ħ�F�����{9x���~��~�0NZ��jД:�#��H����}����K��J��n�"���A4�K�3������v���c8Mސ��A�}'soa)��X}>,���qzx ��V����I���AZ@�G-�	�6)Aء�ˋ��ݽ*�Ћ�z�Tk^�5�3�|1��+Q��(\��YZ^��Rb���m�a�Y�
:���*ҹ����"�}�a5�pP�V��#�
U"��:ԭ'��FtA��ݹ�c��J,��]�Q
�[�cAk������ �9�	�fG�nlɒWY�MG����BB�C���6��h���>�?��%��{��������e��$�M�9(�v8����}E�~�&��0O���(	� ���0|�"-J��I ���J���c��ևn�bL�ŌXY�5�i�O��)�%:E}���vm��YS�� �M#�����὇5�k��Wr��<(��T����Ə�
z��Q��t��� �{x)�R_� i��HX�4>��XlxVHYEB     400     1a0�A�W���l#�<�f�EW����z�L9z����W$�;�`Rڣ�a���y�]/g�J����u2D<����.�3��è�њ��I����=
v�]�"���e~�T?�y���71̜Js{������4/���E����sN���')4�%��);_H�F��Ts#�g��\�Q��yD� �< 1���F��� �Уqe͝e>!��3�n�B7z͋N)�c$O��G�Q���A�%w�:����}fu�Ub:+%���#~Ƽ&췷t<�L#����<?�a�UJ#- ��A��vs.�։�c�+���;�yN�׻�W�<��3N�e�	Όfޜ�H"����/%�������6��rM�a���өS��k��n����JT�h-��KCȫlT�79pA��[�?��zXlxVHYEB     400     130���3|�%!�	��!��Amq|�������3.=#O�3-�9dڿO��	*��8x��*��������$]$��LE�D��U�.׵J�S�SQ�;��!zc��'C�Vb���y^Z�����c_n��h��;l
{t�t����JY>+�~�]�JF�'�Ŵ��۩v��`���\�!������ۧ�:��M,z�APY��@�N�����;������Q�lC��?� �uOҿ��+}Z��^��qI�*�� ���۱��bA���H��w����$pLZIb�A��I��;���dg�/@��R#�XlxVHYEB     400     140Ћ�B�W�T��Z����ۦ�9(^��D�fq��zr�[ڿm@^�R�:�����<K���:Z]��yT����G���Mx �:&�Q'��3����F��.FMj�̥9�c8(4(���g�RU��	�	�7C����婽��C�48�R�|�S�::%n�5I����r,�v?���}龏�\,�� ]Qi����y!t�Dś�e����I�!����Yܭ�KtU�m��,w�ҋ���8}/N%p��J)�����&��T��Ig�':��i������E`��@!�bq��{�?kqXlxVHYEB     400     1c0lM��w��㿔_�t�R�hѤW��?��m�0��CQ��l��q�"��$]�&�(�ǔs���;��w'�d9߰�5FA�g��E�+p?�SO��>lRa,�]Uu����g��C� ɧ�Rc-G7���9)�����H�o%A��Q <��t���6p(�{�����`�G2^���d�����b�� P�7��@1��◙�uiС�9Q��\��@,������Pʹ�wB_H���K�S�ٱ����5i��&�茭��|����d@(��K�T���H�bT�Ґӻ �>�*������sdH���tc��杧 N���.�Z!&S�U��w �����R��bU�}�ɖ�&VNg�3;����j�L����{�Y���/u�>���� ���S�'&�ȯ.&,�+*�2�h���.m��;���G�9�-c���G�B��D+&�2g��1��Y���(�ޝ�qXlxVHYEB     400     200�f>�����������@��=�~��&/T��L��M�,5n���&�#z�L{~�{��P�"q�"�Ū�w��(x�'F>v�����bx�2�Z�,l��җ����<^A:�t�5�H@����Q��x�|���K�	LT��Wa*lUsP:{�nWlc(���:�����3�%l� �r�ػ�u}iQ�/y-���X��r�����d�X��#\���D��^L�	F1�+묑�w^�����w&9�Q�xK��P�9E��vG򓋍Ă΃���L��j��D'c�X}W��?8���a��A��!��w�|}q���
�Z������.�����/�HvG���g�"��-�c9N�rً\M��>��,>���槜�	?+�B�q��*�4C<�9�� �zXe9�����P�^�98@f��j�F�碻�F��]���h9(�0�O���G��x��!3An��ʼ�|���3*^�H���q�.�W�OF�钃��XlxVHYEB     400     1f0bt�-�R�!w½ɨ�Z�G~^׻��N���E����z��7.G~w��oӓ�y:�� ͕-�Ӹ�b�?�Ni��1PRY���%�����a���d��������J�M�2�!�ڡ�:�Y|�6�g��T}�%!���UgS{}�A��j?ɽ���S�N�z���2�άw#�V�@�.�`huU'�pt<Q�Q>@�T�Ơ<�چ"���0O�^�L��5uWQ�ۡU1�Q��*R�OWfG�1��{+圞�8E>u:��m���#�M0D0ȥk�en�����\�Ү8N�
7ˏ���J��N���L���C+��l�;�����C�||�L��ώ�%ՃT��Pl��m�Q�I>�@W(K�G�L�4خ��+�Ľ9ۍ�Ɩ���E5Y�]��OK
M�+��Hb'KV��k(%��-�
-�ק�*�������	?&�n���wq]l��SǕh���)�qԣ�'�UD�sL3�,���7n�y��gXlxVHYEB     400     1e0�Ӝ!���>���q/��ǧ0�eC�6_��S�C�ZPv��#�C\��.t]�y<�Ni9[\l�[�K=>���B��7x� �PĽ'�G��+���� ��������/�:��>�>���M?t[�z+�)�S	�r��}�P��� �.���ld�ʹ�4�:��'7]"�k�O�����KMW�/���;��4�<g)V�<£�3��q#@'*s�='���fsvr;)䤢#>�u\��
 ��	Ia��dPU�R��L7��
�;+9��%@�`[�:�0݂�N�r�@���"�ы��d���Ź� ӎ^�S�Z��.O��AI�"��{������Y�F;�bZ�r�����:l�.��yĲ�W�Z<��� �:�$**�r���M io����]/�"�v��۔��@`H�r�0>�G��]?Mf�E�o~(�c���;��7 ��zZD�����NK�"��,��XlxVHYEB     400     1c0���)0�q�L��uU#De9yDxX(�����?�G��^;�N�D����/��o�P�ȥ}__g���5�/:q���M�z�̢c8@j��=�[�p}po�A{� �p]��w)�SFKj�"�Ҫ����Iv<��y/I���g�'+$��k��M��/�2Ъ�ʄ1̽j��{�ogDY��\�I����zš���ـ�<d}�j�Ņ���gS��\���}� �-��ؠ��t��Xٰ{V����Jd%��d�¹�/�	� iO��gh��|�Z�lj)��ܙ[��Ѧ�O���{�Ǿ[ά�E.)��u�QTTT� &�k�<��j����|�R
f0��+�9�ங\�suX(�8$&��]�=X��^`6�kH}.*F��vܟǱr)OY�N��R2l�!<gFv�YIġ�\H:Q>��.�L�.X���w�^� XlxVHYEB     400     130 I����x;���X����;/��b��F���N ���\VQQq;�L�ML�k���=�P8.���=Z�풻�J)��9�����;�����lܐ�Gg�[�_~h�g�&u��/~�MvI�M`��d #�W��|
�9'�����?����cr�6���p���٣C����lp#+��n���'�.�f㋕1�kQc�e^�򟵳��h�;���I5e���u!��� �.M�.N��1�$�h���_�L����J��.�""ݵ�v���+5����aFm�����zF쐅XlxVHYEB     400     170�l�0�\�l���X����q�+��{�%i�H3�S�ʥ;�䔭D��m+-�*)SN�ϱ�W���)S+�9e����U�?�Ѡ�����0j}�ݣV���3�}��*Hs���\����u��.��yi?H�]��x1��6Q�7����S\���-;3Wm�})��:����F������ +v�pz.C�N
��1i�&ۛ�=dX�Q�M��H ��>�l	��iI�Hf��6s�2Tcv��l<θ�V��2������U �b�MA���!Ķ9����������� �d�>��W"�Eb��?{�[��.�4KO�Ha)�P���K��d��~*͊99��Cp_W��_�h���Ϯ�`XlxVHYEB     400     110�����}�T��#�֭Nd�;�ݰJb~Y��z��w�
���jjȑd�K�Sy�M�@� �>��߷I�r�oS#���L������-��W TN�?�>}D�kť�'OU�N�v]L%��O����WQ��b�8V�.�_ Y$	G�J���g��F�w[/V/���2t��z\�UEl�H�C��1(���{�E��+��#�������=��߭�	���4	#R\���o�T9�6xn�=��J.\��GOθa��XlxVHYEB     400     140�S�Y����s)�΃���ގ��tN܆��ǐ��2�s�� 7�K�	��.S-�r��u���@x�`ZL΁�]�X�:�o"��K���bI+������QI�=��y0~���,�A��IDl�
<NE�>�X\�W�i�a�1&3��4���N�q�ϓ��� '��M�����#n9��C�q4~��\�j h�r2�>u��z\���N|���}�$��u��YF1cK}n�Y���	��{u�����ʄ����V�V$�ҟ�@���ZC���c�U�P���V�'�� ?��1�X�5��ɚ�������$׳~�XlxVHYEB     400     130�_�}g�K�T��M�u��=ٱXŖk
��r�GR�?���{�:�~A�_��	!9�����F��(v��N7���͡���ǯb1�P��u��B�P	o?����o�+�0\��v� <2�2��N2k�
�m�J��:m��p�	m̸�t��Dvc�ܜ/2my��,4f:����I�K�l��l��Sqt����1�z���>��aW�l�֗9Ԁ=�\�E ���u,Y}��t�X�deՃ	�Q3��� ��!#��<����$��?C�cR��=G@KN���â/2D�*���U�����&|�>XlxVHYEB     400     130&	T�v���p�.VE�ԭ���*�y�33���"ٯ#����^o�ю�N���H�ӝcu���S��f�N�"ș<A�A)��yd�Cs�R9�*zF�#v�?��Md�|�������K��1�I��2���o*�P���*�L����U�#�+��Ux��//JS�1�7�V��z��n��Ec����W�tI׫�#O�c�0��;&�q�0A�;�/���>'�{�� .ׂ�C�{ݪ�tX�d�Q��[%.z��q�5̸����1sqt������:j،x��I�5��)����8�{XlxVHYEB     400     150D^OmI���CizTh��1�4����Ht~J��h�b��pu��/�Rա�R��$$��*�By���Z'�&���ј�\*B�@F���D��Mk��6��jdi0��-�':��@T�����W�˨.z�U��Ս���Qz���aY��I��g�l�2v�M�|�cr�9߇��dȋ�XFBi��o%�2¾y/�RT;.k���Fq-1ℛ���
�����
'-h�UBS=帬qZ�j��6��.�k��E�`;���.��**_qj��!a�t�|���I�4yӬd�,_q��{�����p�3z��v�&�TG��)s2�imiV|��u���XlxVHYEB     400     180�0*/��fup�����~(��PQ�	ր����i���4��U�/�*؟ܐԓ�g΃��qv�#>X���mF���#B�L2s��;iʡр~Y Y%����@�d.�9��;�4��$�����������C�f�c�	@5�;�פ���_��D彥���^�NP� ~}���� �����
P�˔3�2�@_�<�@��'�T���A�$�U��Lf�D���#w�Q[���{��R��O��=<�M�5]Z��޷��-�Q�*���`��aӡ�c���2��!-^��)[�uO�Sġ�v�`�nS���]��b���Tv��z��ɇ�|̭Է}��:9���@�TA<�Xf,6�<3JA����~��XlxVHYEB     400     1d0��3e�� w:`�)��X�y�D���4}=�U1�o����(8�Ts(�)�fQ�~H�6�;���·"�$��hz���gMX4V'(l=bNυ�Pɷ{RtXhj��W�T�^.�5P�}�E�`1�� ��1���*�%{F/��Rc&��}�����񁏘�P�:^��%c��T�*����I��쇋�
v�mY�}�#3���H�Rp[�Hg��	X��l\�f�<���tJӻA#��z�S�B#\~�����&�\¢�y��Ah�	�{������b	]�#���*�wG/����	Kjzׄ�&8|A�<�I�1���B^*έ<�4�l\/����d$���)��b�yN���ᥟYΉAF���2�t:�YOY��GMI����֟���A��kza���3�7�R@ⱢH�k��4���qaU�e�VA&���zA�@����G2��M#���T;���l�XlxVHYEB     400     180T��5M�n�,�{qɭ���P�,���t2��p��u����c7��r����f#�$��ʢw�X�ͣ�e���=4 T��3���}"+G�%P1}�y��LA&��I'� �M*h��3��D�_�w�8���7`Wt�0q11J�@_0��#�%0��������>ަ6͛.��(��� ���\��_�,����OB��j��g60lC�6���l���uM���>0d6e���ܓ�[��b1��"m��	.s4{	5�
�O}�X�V`�AN��6
�jC�3�.H�$�1~��?05I�B?�V,˯ؘ�f�>3Ao�F ��Z�OSP��bt����0�]�:��C�� �*3 m]���s����B?��i�5�XlxVHYEB     400     150���w}+q�5t��Qk��2�Pu��k���.��0L�7�4�����2-K�L�<�F\)�zӟBcflv�W��V�E�O�1�ZH��'�e�� ıvGy��>�3Q����|�H�V���L��4I$nm��R��0�������r�C�/�S ��y��>d^���4������3����Q	;�o��b�ϊj�#�6����v�'wx0]����o�Ϟ2��������Y��7�0Dgq`�f�h�
_�zd�4�9��_�O��΄�I�����h|�U�� ��Ds�V���Hf.h�j@2�at�s��\�����o�L&:XlxVHYEB     400     1f0Z��,U�R�`ɿ!w
5%�n�W��j�Q|@q!�����Y
������\:��\M/��/��O�c�y%��\�+-m�v�r� (�[U��xB�4�VxƿA��QG�Vzz�3��KT(�$w"K?2�	w� *�zl��[igsC�H��Y7CÍF�߈����`,jX���j�n��:�H�!4�9��%,����)EBd7F��!��fB�ï�q���X�d�ؿ�.��>���w��#k����k�-����?.�a���͞���hh��xPh����_
%��Y�u;�*P.�͊��bw}5��M�)>��ͼ�
u������܃�Ųq���C���g���,�2NSR�B��������S��qD�t *���z�P�͚"�d-!���}:˭�,�a�z���TCR���y�?k�.�+4M�G ��?v~����佖�:Շv�pw)�.䅼@`�yҺ~�N�'T�-���>BXlxVHYEB     400     190�T������W�G�GW\�Z�C��k_c�W�!^N��揢��[z�?�G�X�iV���C+�D�kK�bp���?"�0%�l�J�Zm>#�ʮzq�P���6�'�ԓpE����SxK9$60{l�l���m�޵���'�(�f�CO�)hܷ+gR�%;{��Ӳ��`X�$����aP��*w�ҰL������� �M2��m�b�"�o��6���+M4a$�5>�>_�kV���BehD ;c�cm�>��M��w��������Gt���$�w*�hv���h9MZ��M&^@2����T,��_��r��&,��пq�~B�;�%F�/��)�5���Xر08go-����!�-�0Ɣ#,�)^����0)	V�F�7�9׮�Z"XlxVHYEB     400     170J8ј���G�nHa��NK���d����r��h^�+Ӭ9��2��Z��L6Î�4��~�n�۲JWLN��Q�v�rB���(w�&�bHb�1#̔k���F&w�o
��K,�q!�E��-1,.ģN ȅaYˇ��N�݁��j��
V"���OIdP�yV�@�fQ趻Dʱ�C�lN���		���?��09���|M��w,��J�e���@�z�j��n�!G)� k5�/�T��Ѧ��]��c���{Yeݔ}�f�O?=�;�G�8�k�+dF̿�C�͈�!T��D�8�{f�WI����C#Wnέ-�ֺ�yᦹsb#Ș�(���ש��%D��}�>/3�ݐ���H�я��d}~�u�XlxVHYEB     400     170���M~:(��tt9�����c�Te(�� ���]�,h2����y^]$ -��Đk(�+�}U12�@|��ĳ<���͓�2�څ�P���y�_�o��ڰ�H�h�{ep`<`��>���6N&�p��t��WCEO�L��T������םB�V�%�}���|}�P!��yR��X��e�$�->c/�HZ�% ���|k����e�@�7�~��S�_�Nh�f<jBL�-�D�%2�Yg�?K����	�uA^@z!r����J��5B�2g�+u�~�r^REUI; �
��lf���?Ŀ�+��L��ʓ�2����}��KY�	F�D_�@��ja�ڰE@� �~�$��!4k����~s�l"�o!�t�XlxVHYEB     400     110�!��m#�b�z��eV��֋GNH�A���M� P �!z �l���T�_#}ݟ�����#B`�.�Ő��;;7p6KXQl�ܮm����w��|�O0Jo"�4b�X-����t�J)ޏUO�Q�z�z�%�^
���Q6�o�-���)1�'�{��4VP����S�3d}W��6CtSN��#���r1�f�. ��:���Fj@`�{�!�ϒ�᰽�17��QKUitEK^e�+<w��l�V�Zr�$G�2XlxVHYEB     400     120����?�ph��w�����o���|��������P�o�VY0�$�J�JWpWuGHW)�P(��%1l����!��;�-|7����������JO6�D {�Sb95��'����U4�� b/S��.���j��:���ot$r[8�H�0%>�P[���g�s�Ӡk�'?�JwP��$�J�j��2�����������LI���v�b*-�?�NAI�5/��9�+k��T{���6f�KxRb�y	�+�(��
��~9ya�X���E�c��R7���� ��4�9XlxVHYEB     400      d0����-���d�]K��� �^)[a���%���n�D���&9c�
T��@$�P�~z܎�uL��]�)J#H��SUt-8ϛ�l�pn�接�X��%
+-��j���P�K��f�����'G�`9�A�b{���x����8r����F���B)���{'�"DU�u�ѵR���ۤ��i�6����?n��,6��=0Mn���ԥ�5���XlxVHYEB     400     140t�v��\����ϳl�(�Ğ8zJ���]{l<Ȣ栴����f���h�����z?%�Okq*�ARS�`">Ǆ��L|�e϶�H!�������'�H8�)��(u	J��q�s�?4x��equ&�%��%�F\��;p�q5�0��V��ޑz���C�E�J�((�v��Sx�:�M�=Όٵ��7#m�Į�i���W�Y��9R�o�}��.R�P�"���\@���R}�1�Ȼ���l@&�UiAWp�"�F���?չ߱������;�yz.��c�j.mn41�a�'?�%�����m.R��힕Jdx�?��ȓ=���XlxVHYEB     400     140�Xs�k�朋��=m����v�ꤎ�]bQ�@H?����2b��!
�m5��{z)��>B�2n���u����v<=���4�SW:���"�0f�F����<}�s�DﶨΒ��O�L��{�
�D�E��nڿ��I<zM�(�=� Ck��x��;&�~%o�7��pL �K���m�ky��F��x�E���Q��̞������W��r��ָ���{!k�$L'��۷e�N}]��~0��}���Ж�.��W��B����/�Sx��|!��h�|�i��V��Cb� �g��[1��S��:���0��ڇ.a1���XlxVHYEB     400     120=�kO���~%�+�*8x6�C�n�;f5�┶�\mo"�I��C���ڴ��������GZ��>��W/������c�&}�N��N��y�h0�$=�0�\N<'�C��X�8a��B���3� �/xZJʘ�;��5��+iE�QCR`�^�^m�!�5�T�*��4�>�O�)����9����+�Fe���C�G���1ܔ�m2"����t|��a���-S�$(�q�]$jϺ�Sߕ��/?�BƦ�_/��z`:�!\�O�h�<��HضRa,�X ��pM�XlxVHYEB     400     1a0����Ҝ�)�H�G2�ml�rpL�n�Nc#�A}V�o-��+��+�g�D�+|Bǜ��>� P)�nJS2�`���ȇ�]�!'3U��H�����dG��͑���JY�*�'����[��D�n�U˴S��L�{ �օ�:����S�2ˏ6��/��	���ox-�_���BX���[y
�>�c�^J1�	(��\aL�>�aL��@�ja�`1<xK#�ʹ������i��2ZE�c�2
��K��K������k�uk�@�X8���L��KQ�F��a������C�j��9�z��)W����i�(!�{�:��Q�@�L�ݘL�1��̿q@E����y޸m=�g����7ۏ�D��k>S��<?�>jU�k�l.�D�R�k*;�,���wx��Nq6��6� �ƴhXlxVHYEB     400     120��ߚ��P/��~���^���,�s���8#_�m���SIb�2n6��1�18�<����u������(D��]
�h��s!-�=���Wk�b�'��$�W���J�p"^m`?s�ص([&V+�!(
M����X��:�hbޖ�9�gqo���Ᏺ����\O������6Rea3 H�f��K?c>t����&6��z��0<|�� 뫫S�1�B���Z���9س�4N�Q�ꋭ�	�X���m�֔&�7�	
�!ڳX~7 U�pO�������2ϧ��HXlxVHYEB     400     180�u��0��rK}��T���C�������R�WT|}\E�Q�9�/�f�آ����ȄA˿=/*�6R�>��q �b���S�舥X��8�iRy7N����;)� �\��e�,D��N3��X��hwoks'�b��n�$��D�絰�j���]N��l�J_)j�o���	�ɪ[�wj�y��ʣT` ޣ���o:<�5o���TP�7Hw����
R).F�pʎ�,sC�j8߮|I�	��ْd�{�.���;�9���k�7ϩ�F�2@^�0�*c�ȵL(ņ�����$?�+�̐�<4�6�Dh*$O�-��[�(j>��p�+`��Tۦb�D���l���^m�e!���v�UC8H�q�D (�K��j��|��L��${J�H��iXlxVHYEB     400     170ۖ���M:���^	�ѕ��k�6���M��u�v�xJ���gDe�%Rգs
F"�<��~s���}�k��.~j~Z';�Ѡ���qLd���T�����=X+ 
��e�Q��q9,�L4^%�_֪UN[:plQC����d��m����c��y�-��:��n�W�J� ��yK����g���K�VCg�[�A1���]�:.��p�~F~ ʷ�6GE�p���$�����(Z����} �A�@XM���U�	��M�r�㒾;/�s�[5��r_��/�~���C9�M���AW��n����uƷy����CNbk���:1֞Яt���Y$s���>��Y�� ۯ��$#����7�f������XlxVHYEB     400     1c0�b��{�U��Ǒ�SG�n�Z�f���k��j*��E(���qk�����('[����<�m5<�0c4Ae��[آ �������@��gh]P�r�6�L� Z �ӥ�lHi�&�+�4�2�d2��
��1�c����v$[\Q�`*�ͷ;�.~s"_Sn�c��z�.���?3�cD�f�g{E+�rs�s����J��n�he����p�\���wMh�Y)	�'�vc�B@e�$��o]��+� p���[�XZY��>l��/ף�Z�qC.�/��]2��<����b���6��x,�_k�zYd��0+�5*��6��zhb���=���Y��S�xH/�D�3���X��L;\�'HL�I��|Pe���u�o#N����_��m��'l��׽Fc;$~�X3U�iv�.2��v�0JK�)~.;���p$'l���6?��OyL�8��D�A҉�XlxVHYEB     400     110�%x�#Q�E:WC���p,���C��m�B��9݄�K)��J����%L��7l��<������$�_O�7}�1ְ�|z�ٗ�S�?��-��&���|�~89�j�F��+K�_���*��YI+d������?��!6$��쵊08���4�f��W
G���e|�$y��s�`��	����>���gj[k8S�o)��4V����<�Ѱ�ƴ��<��� �y�9��������vѯ�1g�1B��c����$^��XlxVHYEB     400     170��Л�a`>62�BE8s��hᠳ+y�:�G�L$�z����,�,r)�*��_��o�&pK�1��@7����#��RsU5�+�
���a>�7r� ���A�n0/�{���Q���6��$�Kn����!X�#A#.�V�~�����)�$�����`�|�����A`�QT��'$��]e�k9퇈�TwMq���YB�=��y��aޫ�A��6��1=(��>�6��$�9J��@�-˔a&�2��C��ۏ}4�'®�o��x Ө9)�zTkT��9D+�H��R<|MV���	�9b�h��N�]}��h�E+gh�/fga)�Vd)��Q��Q{1^L;b �%���g< (�j�XlxVHYEB     400     170���j�& �9�Cgy^�����ͥ�)xB�B �z����J�E�hat���ļA�O�Q3n�wR�d#_�+����×%����(Bl|���9y�Qv�7A��e��lF���>���I��Xo���8np޻��@V�	��H��qa@�=<�|"�:\VA �����=N:A_7<W�!����a-V'5&O_4����5�����!�����17�-  �܃��lr�;p8�ͧ�������&]��A� h�G�)�Ƶuq��D�w��h�ȬO�G�=�懲{N��X/���T#��X�������[���I/j��P�P���!#q�0�Y�|��P�i��e�p���}XlxVHYEB     400     190�wL7yS��N����b�[ﶩ�*�[���}3U�{�Si�� ����sU�̍���$�gn��F���08zHb���>mYBli�V]v��=~�����|�rֶ�B�A�2%?�]�����n�|WmNg��+�-���s��@���`�4��P���^��$P;B��>��j�����kw����'
W���<�x��d��V'X�cg�:_㱩ƪǂj�NƁ�5R��;�M�}�Ҙ����]�֬��^���~X)"9��>�ʪd?�Jŉ�DW�����9�{��V�F'۶B@��`�Ih���y��8�����f@�� �bKZ����?[Q@i�nл#��}ɏ@�|Z5���bb����1,�Oڸ���C��N�UVL1%5���) W��q�!:XlxVHYEB     400     1b0yӵy�����>J��	�y�(§w�3����A=}N� +��Y{?7�b���6C��=� �n@�	�@#��&�����$�lD���p*|���k�qu%�݃�[��V#vf�����[cs�	�����R������a�H~�q�s���<�����K�*�'�ӭQ�	(|.8�xCw��в2_��<�d�؜Ae��r!��w��q��O�i��F�a��S��y�'ٮhb����D��퇶��:���f>|��4j�P�,x�:i��l(�Wh�_>Y���p��u�ZX��@⟣��\V�w[|�Q&
� ��U~;�tgUz���e�����D�
�|#s�Y��I_H��_��~3A鷤�w{g�=z�����k��6�"�&�$�W�kW��彠������4�V����-7�O�XlxVHYEB     400     1b0NY�m�}�t���`o�h�5&0W�9±�)2/�9��kGAc?D��\����lF99Sl ���V�4kA� 8Jx¨?�;pB	_u�9l<����Β���R�Pw���'O��'���-J�(���Q��n�������hJ���BY����e�����R�����z�6L�@��C(Oaٺ���>P���J'wޓ��S�iC��33��?��|i�x�5��^�沗����t�:n1����"��'3r
�h�I׼cp���p��`r�l1��Y�C���~
4n�H;������UԸ��*yA��_��i���o/�dȣ�k($���%z^����+�%V�#�{e�Fh���R���Q6;[z�B�����r#�S��R|FKk��"�U��r���7��z�S�9�<$g::���WW��7XlxVHYEB     400     1c0��CޱV�r�iی�w��`��P�{gX�Fs���s��Wax�Lt��0Kݧ	�D�Y%�B`7ue����7:0�������[��&�RnS�"8�z�_�dP�bST|��IC�"-��'�M���8���
(1��Bn�r���������h��l���c�'�Чg��^T5�8����nP�ߤ�`'�+��f����M�"oy\�B!sI "'�fǘ��z(��j�y�h!@
�J�U9�h�O[��JE2-9cy�SN`S_a�h� !t��tmU���R�	�:=Q��1j5 z�u�$��������L�^��<��b������Q�v�HjDڍ��ˍ�'ka��.��ʘ��ĔaP�J��D��A�:� L��p�X(��m�BA$0��i�9s�_�)F�걕�l�'aU�z,���p��Ӭ�,�6R��crXlxVHYEB     400     1406��^;��I�d��n!4]�w�2�՚eo)4��q�Й�f,ܝV�n)�����%�ד]���,;���>��J����K{
|s�&�́u��Bi��Z��ҝ$m 1\M��C���Ⱦ��Vp'�������hZ�%58�ج �VxV1#���k�2ꨈ�;c�Ĥ�O׾�ګ؊�/f�֧ւ����U�4�����r�M�*'҈O��.Ǽ	�g�D���=���žEފ2���bN)������[���ˇ��a9�����ta M��j�޶�f:�Y��!����xf��c���ݨq�&XlxVHYEB     400     190��u�p�:���>��J��f�mu�D�Ç�hI!͞ptW�Ŧ
+�&dEG�����BJ��+
{;O������1��~My����a9kU�do��B)1�F
���<�N:�����qeŷ�,_��v�m�r3(�|�s�:�t��.��#���_f1�+��p�ъet��0ZQ��O��	�vޙ:�^�૬{i�1?{�K��O%����Mc��q�K�&�vn�]Nw���"��TO���M:�pl�NSG�bI(���>K.���d=CĔ�Y�J�J'��߭�/����Q;(�}�c�I�R!�ce�\�w"��W&=�K��^Ap��� ��45��0T�hB�{Ć,��T�1��4bV˓��ՙ|�$��/�q��-̔�L�XlxVHYEB     400     130�f�E��J6��`�J����<,!tn���$��w�F�2""L9�%E(Bmܘ��խ��ߜ��S"*�/�p�X�IG�
�n2��2 +z�K@6l��ڱ������V.70=ʄ�~�(ټ���ﱂ&���C[��Y͜��6�A��9�U��Jc�·`IT�bA�@*.Ͱ �H�4	:��G�|��M�ZŒ�`[v�.�דnʙ��W�r1~����j�7>U�N�	{��|'���Ff�P5��I��!D��J�Sv}:$���/I�_XB���e��3n����-�[�"��t����XlxVHYEB     400     150vD���"�[lNċ�9��J\��?��XQP�h	D��bB���E��z�Ѭ�BZ�*��j�`�k����!e=TNY�/�K�7����f��b=��r�nkW��~!��D�;���tv�A�j�/HC��8�Ǵ����[�S'[;��b�&>7��X���>W��������7��d����k�h�n� ��P���>}�U̽w�K�T4���[Q�;,Q��:����w�f�л����Kq�CY��m���ct2��1]��ܾ F��Iv.�.�v���y��{E��>����.D�%�p�%�Y�Hɓ3́������UXlxVHYEB     400     190_��of7�.��<������Լh4 u���Z�l2� }ۊ��!+Eb��ߗ��2��[�=5a�KT�}��U�J񖪏���P��7�
T�0`�r :�)u�J��F۴�I���@Hk�fㇷe�T�KM�{��[3��`�gN��)���{/�,��G��ӌe@���rRC>9w1���7'�Vv�}z�����.Y��()o��[�������ۙH�sKi>���v_��
B\�hl����}^2cC�Ix�T�����O��y�]���W����Z�l��b�*$c�Q�����gJaUW*%���I�Ȓa�X�3��l4͛�������ac�b�U�2��"���� �m�i\��9,U����G]�A��������XlxVHYEB     400     130X�ڤ\�繇M܈FR�(��v�T�h��lH'�o�S{����
�H�S�#���o�`����`�S;[X���Qc�� /��6az�nZ��I%�8�enC�#�P�k�����` �ea�@�[oُ��(ג t�&u��ɣ^-ǝ���=�D�(�6c����&�eCP"�ۢ �H:
�u���o\�`||;��N �.�t��=Ί7�f�F�BkZ@�h'[���66a���ڙ�O"tSػB7l�G�A�(��0���k�}�F����gT���T�ʘ{�H/6`�eId�����ÌY����XlxVHYEB     400     150e��%�!����ݧn~�~��a�*�r/�hKj���i_m��F,���\~,k"������>���6���؊�]��:�5���{�TC F=���8i#���������]A��J�l
�K����K{cO%�a]%��OH�H�]���hq��1��&Z�i���T������R��Ћ?;MD�RrEe�[�@����N��"��4�'.�|Ûo9�7h,�Om�O�a��~St)(N��" |��]?\}$�k�*�2R�%�8*�$��n�u@�5��"[J����j��ҸC*-r�����V�	-��$n]
��Y1��}�.�a[�-���4�~XlxVHYEB     400     1b0a���#��O1DB;:������z,��AL�i��$�@1s0$��6?�]p#�k�!V%��I$w��f�&|�k%���7�uG�0�z�5�K <�~�g�u�K�<4��&E~+$n�BC��)A�h�T���*��͜����0�H�'�x'��vm�҃��:�%�*�@ʫ�F����I�
�>�4�U��i"v�O��2�=�".B�!! �V:�v��ܸ*IG��l�����S���)N�4f�{1�P��3S��Z���a,z��aLI7\���ou.;�1b�sR���Sb-jj-	[����?e$��Å�U����-�z~�e�lm�"���d��*���^����܈����/�-��de��v!V? ώ�<r��A�U�*[�2q�|�����4[]D�$�a2vG�����q�sXlxVHYEB     400     1b0=l�I۸V�v�5�BS��J��f�(�T��p_i�8�/lu�A�� ~)]�l��	�B "��8���Bc�����L�I/��J�t��)�6��P�+�Z�BP2�!$��F�<5���ۻ�Kp�+ I�{���:u�g�W�����;��C�er4 Pz�n����_8����fJ�3�ZR��� ة��6��+b �_�m]�}��*�uןPh.�p���q���8�2��cz�fr�f��^��(P��V���	��rN/X���h�#<)UR�@��1�����O���8ך�6��&/�~�����8���>��<]���su�S&�����+ ��c�M](ɺ� 	�u�5��HD�:��>�U�!�2@��p��d.X49|)��c)|Q6s�>��"��Ԛ�qϝXlxVHYEB     400     170���}[0$]Wj��E	&��"\ǔNP+Q5����m쿦���=-��;�N
�7���	r�8�]N�Nfe�!��2�ӄ���^|�\�f�m"�{�:�u�1C�_�!J
R�f�[�ڋ6���M�f�KC ����رcHP!��ƭ�B.�W6���t���C��BIG��=.��� �l�����`��D1��G����h��Lr÷�S�"8�y���P�9�V��ˎ��A�xvi�ۄ�N�c!m�-�k�C�ُ�?��#��޺{�nҊ�`�xA!��v���(�5nT0�O'��P���ovȮ�!J���^MۚVn���̦tHUcD��b�r��� �U�?3�Y�@�PlXlxVHYEB     400     1f0�b����3�|8$in�^�*�SCھ4L�./�� �3��E",h#�0I�öps��풿@/JE��\�����O�� �	_���W�O�#�棴�G�c�7��
��#P�߭�[=������w': .C� g����fn{��@�S^��~�\Ҙ]5����c�OV��A!^
�H��g}��p$�� ���<y+��6�~����x�	��������'K�4JrM�������P�ʼ��ɭ0�Қ�wW�N(w���� u��QkB!�|Z�Xu��+���r��0P �}r�
AZk?����س���
BMc:�7��)��
�Q�w�D�!�I�\�쀴@5���Y��g�c�EcX�����7�%����E�&"^�D�G���73��V��#G�wz�]�WmJG��s�_�o5���7�O/7��g�r=�v���[�@��%LX��2A*��|�5�8՞������������XlxVHYEB     400     130/���rgT�n�I�1z�	�ȷ��8�`�֖/�a߸ݸ;}�=`7����5��z��C�Z$u���(,9[Ke���KO)8����V�0z\βqg�\�r�;̌�)}�
�kd�"��L,��W<*r$�*g�ʱ��%3A�3f^�=�����k��;�R���kh3�h(G���٥��ٟF���:V��ž#i=�1���!+={E���^�?K�&G�	��#;�̫��7�,��`P�5�H5�Ӈk�?�^F��i�-�hW���^~pD[3�(O�~�w�`+���RzXlxVHYEB     400     190��ԛ�1Q�y�c�0���a+�hD��G��V�ְ�����j�T�@��m�Z/�x�cy�\Z����H���d��i[�mE��,~��,r8���_�ԭײ����ZXW�ACvgo|�"	�Y��!̒�� �������K�����U�N�&.�␂�Z�!v��Џl�%��nc�V�]Q,ځ��kS 4d)�����a��J3�#�r~���׆�ko>ͯ�HD���
~ˉ�[�jć5pkX��/p�xA,i-�I�����S��y����a�vPښ8Fc�ɻ��H�9���0��w��ԴY(��w��R��ݩ�M��^�G��Ao��`Q�" �e����nJa^>tm�O�j7u��*��és/�m}-E�ֈ my_7C���8b9� ��>	��Pw�0��XlxVHYEB     400     190j�� ��zi7=kŢ�9c�`=��-nF��O��ڄ{s�e��W��I�!��U�u�l�S*^�;�lQ��!�+}b˴WH$1;�a���G�95�gQbo��Ҷ��0�x������N�4����|,��iGG��;dV�NT�w�-�� V��ߨ���KL����p�DW3{ �9����&@�$�&�z�q�n���u�
�,e��S�͸%$���mr{��q���Ӥ'f�����	�1붶6��	: ��vC�N�;O��:1��_��=A�R��R��ڑ��(�dM��??� ��9�
i0��$X���G Mv��(��
	*����u�&�^��e�f+����f�zc�6��?�K��}K໴\1e��'kz�Wt%K@XlxVHYEB     400     120p����Fv���j1�'���A�|
��[-����x����qR��pV5��!���o��w�-���R����щ9<ח�S��j��ɉ^�2Hs�����/��� Y���jSY[F)G�̈́98�〛d�f%��X����r�!�)�^EΛ�[1�?�Ho%��3VQ����Bh�c�낇H;�d��K�VWI֨��昬%��x�v#��"L�p�g�f  � �A�A�/�Q�{3�Yhmj+�����H�!�v�"���`݁|��7������]��О|E���XlxVHYEB     400     170��1Aj:�s8P�{˅l�n�*���J�J`0:!�+�i��-��Ɩr��t'F@�T�uw�l�:��#��N&�7Z��1��$_��5�� {i�%�\���pf�m��jx���BӠv~��%:]�ٿvU���N�̥�i��!C�����ġ99$9(Ϟ�m������ą��X!��а��s����%�s�6�~�L�=z���ΌGF�#̺"��ޓ��o㌢	��ڰ��A�0hv��T!�p�*��BsྖuW��U�I�mD ���@WB��0���p�H7/������H�FH�R~$���#P~#�~�a���;K�29���8�gG|�8��4o��KO�y��w@`�8+���XlxVHYEB     400     170u�7)��7�c��om�� ����j+�����	Tmv���Y.�!iap�yn �k��
���x3Y��4����^����$ǵ�`��vm�B����[%��`���E)?�d�)���|oN1�����?u�^S j}l���3Ȏ"Yg��q��F�9I�7����7��tפd�ό@��b����M�=)4&."�����x5��rFݥ��w�s,���o�8��uY#�,���t��ѽ:NYT�q��B��C�k���+Nu��� ug��i�8e���7�;�O��;*����d޲�׷�;Ͻ����+[��ϟ��NU�ݾ�O�NZ�KP�g�S���b~�zڧY���B��sQ�D�0�XlxVHYEB     400     1805j�spq%޺�Z	����%e/�bC�I���Жc�����*��%9��_Q�x��b���)[ې~,i^�R;}c�#�<S�_-N6�j�ɿ���9!���z:���_ǁ��{���;Ϣ��J}q�:��3	Ym�u��R����_��K��&��+?�}��&\��5��m�#�4hoжyѬ�$��"=�i\�6Y9���ƾ޶$�	�c�[ V��X�N � &e��$�h��s@Q}EvI6�g��M����1��t�%I��W��)n�-�֝sI?"2�uq�'����f�T���`�x�U���Qg��]i��o��'�J�=��'0\nJw��һ�QD}��b8ڱ��b�臹�dMQ�l��%@�ľ�m8�Sy�Lڭ����[�oXlxVHYEB     400     100��s��鴣��2�gT%����ڗ�:d�Q�޿�`�ڬ�@9�O2�^�Ǚ2a�����d��)�Cr��k�w�O��VH���t����ӫ�j��f�#�*����*����Ց��qU���c�C���>����K*˹�X��Я���Va��3�Ah����f��3��+�stI7���^��t،y�P&�Ĺ!'��aFt�]�(���*b�v&������Ǐ��'���J?���ĕ�%�+� ۬��3�XlxVHYEB     400     150y;a�+T�Y����2J�E���gw�Zc�T%��y/�v��a��ި�S �"���0�4r�-�%t8ܖ��	{(zyq4e����?3L^5���)Ș�z7<h��W���?��	��HN���_b�;r â��$!�Gr�i�V������ ��*��x2��7߯�i	�I�-��/�� ���m�R��B�#��\�ƶs�h�>n	X��!��mޭC�d�V5���=Ժr�pFL�I����oNE�I&�@���X�8ɴ�6�\8R�������VI��لV��5�m�Ek"[oH>4Y��AHk�>��c�ՠ4�ճ�(��"[L�XlxVHYEB     400     150H�ר�T�������[��R�ۥBɅAn�\.S�C���m��g�Q]h���${�iYnD" ��iG��.�iI�Z�S$�tk�md�!�AA�_�S���ui�vt��e��"��dl+���p'm��x��l������v�ܷ��<���M���ߕ�j/�˘���:Y��R�}%�s�<5��H�a�R.����6�}0$e[F�P�%����Sr`?�e`�U�>fzF�+�~�M��#�١����/��*���ޒf=���ݴ��@�1 i��v�'OAP��4�Ib��`���%	��rF¾X�-歀f�� �	�|onX]&D{�XlxVHYEB     400     150�-.y��%*��]��S��c��-�_J�� ��F�WZKg�-l�����x���F�K��F���y�W����q>�Pk�W���0����(�5 j��Z_�8�)E[Y�� �8�o�y"�K_�\���F�m��ЪBU�ud��	V�}OI,Q!�9�
d,�|�k[�	�m�þ��sa�RՄG����^�*sJl��W����b�sy!�R>���`cn0D��Y�)�k���
��Nk�Z�/C�j�u�LG`-{�O�e���G3H���Q7ɡ���c�sE���L_H����9��0���B���ٕ.��� 蔸�Tf�hXlxVHYEB     400     180C�*�,S@��z0�S�'	�D�#*נદ�h�_pU�\�qE��Y�S���ׄbٯ�)�n,rq[�{1�S����v��U�4�߱J�CL�]q��#����/�&g��m��񏯏x.����c��մ&�s����,�ys��,�.`�1)�ן͍O�<^[��A��	�M����<C�U��R*���G����a�&k�E'�!�����'`Jd��"�siҨ��]�@�9�|�,�Mp���e����B��[zԵ�ln	 �����S[�)��
�#��Ю�>��'��v�B��m8w��%*
efQ�N�nLۣ���)f�zw��jc�a�A�1V�H\3���-�w:|�d���9!L	r�����eXlxVHYEB     400     160�21�n"��+ے�)y���T���$+:@<aX!��U
��nKT5ݠ�Uo�+H�[V�0Mo���fL�F��/�`W��csG��|+�;�$7�>��_
d<Ip��t�sR�AfQ K<YT^iD�* '���]�`����>�	
9�l!�h�5OC9��ʸ�L<��o���׵���]׳P����c� a5�h�wh��Pߊ7�Aw��7}F(��2��mP���ͫ���8�"єư�,~v 8�L�_M�K�-M��8���z���f� �&ò��J�,���
"�33A<=��`�2;��:���$����h D��i��2"�aD�XlxVHYEB     400     1a0�?8�1|��@��m�Z#�X�$�4����ws���,��G���χJ*(0� LbÃ2c�Qw���y�ڣ��s����X�d��&@{�r�t-5��җ�bNb�=��v+>wC�Fre�?�^F�Qg�b\��X_B�2c�CҴ48k4m��S����bQ�)A�Ԕ�LT[���RA1�+�U Z�ܾ�$\�ҒsoB��
Вo-rsź�#J�:��ʻ�˙���Wфn���(B���Q86��h�l�b�9�gJ�磆~i�˖M>ߪ�<�y��6)�[}"q�I'ky�N|ʰ2�g�Û���W�[$FZVT�a>>HT
�un,�����F��x����8���X�];6:P�zj.�z�L ����;tR �7{��k�:��(z���<	��`^��}Ss}<�wր���`J�XlxVHYEB     400     1f0ߍ������:�J�*-;��kQ^WAڶp��f�KFK�@aB�a�����J4i�ܺ~��;���m�yȵ��rZ���[1�Y]�X졵Ȏ5�:�/�8Ԟ����c��פ�2]:�+��4*�W��I�}�����OB
5u�gN�+��Ed�HyC��-��^����I�'A�p��SN�U���p��K
��V6%/ ��O�bvRݼ���z�V���F�6n ��x���ќ�w9V�X��~�_K����YC��-�7*�^Kڠ"9h�9[�4S!���h�: ��=��nv��^���v@��F}��� ��%HcR1�>�4�[X�z�5�	���b�_�.���#�c��6l�|�>�#�X���LH��]#t�(6���66�T~����#n挪�����$��6I%�R��?�:�A1�9�>W4YE����]2�V
�#��X<�w��w��਒�d9�	�u�~���i=z� �9MXlxVHYEB     400     140{�m �g;'?u��׈\�����B��g�*U~�s��iB:3�	X|�X�k8���	��	��!�b�M��u���S:��-i��$����*O"9��-�ǽذ�m�~6�"ׁ��臩�����f~�[�|~�(QHz�S�������o��Q�q��d��DX�^jS��Pakӻ�@	r�m��J�Ċ�����W瓡�'_�n�ҙ���][�f����7�&���CTv���cփ�����*�$�?�'�l��)��&�aKWs�k��� 9��M��Umg<�����3�^���y�\*���;��XlxVHYEB     400     140n.:�4|x>M��Ó)]<!�G�\d���r޷w�-Q�L����5�)�:�@4
�$V���Tt+WW}�N�evtne*��m��`�Y~"2�k��e���eV�_��dNk�Fp��A֘�4�k�0�ߥ�#^Gvj��(�4L,��#9���Z������xc�=+�A�t���K��TɈꁴ����7���~/ גY�味d)8TD��{�������3/�����Bi��ѩf�Y�@��lU\<������]�:��o�6�B@�03_ �x"5�� KW��VK6n$��n[j~�It0�XlxVHYEB     400     1e0����"�)�X�W̐nGw�w-Ɣ��l�:b�n+��-#�I:��^@Qu�8B��A�dJ���䧱�G�K���5�B�mY+���*�kA|�N���V��t���y�Ϸ�]��ŕ�Ĕ�y��h�� |._���"�I��=��T6�'M��zϫG��U�=��Ǻ���1[ #��5!� H���|��(��u�Z��k��)P���;g���\-�<ƨ
r��j� ��{6zƀ���By�l;^�f� �U1��Bk�4T8�	��+��������e�E�����J����	��'�z��)�g���<Ek�m�5 ���]�"#tG�.N���Ҍ����P���g��U��=-���gY;�>��g>
�E�fˎ����k8)��5�Σʖ[_�F'��U�����i'�L��S�[� ���У��/�*[,�L$Z������xd^������-rКx�>��{�\�gT��:a�XlxVHYEB      90      90�D�&���b:+��`fVo!�cl�3�XwRį��J��p�o�ǵ��)��������I�"1H��8��r�|.T�=v{�Y"s���c?�	���#�%7�I,�,KXm��V�c�����Br�|pi�b�a��%`ef�Y]�5