`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74304)
`protect data_block
4iC/2PKTKvNPOrwG58AG/DlwwHG9gKwQ4P6GAkluyo0z7FXOeuqrwvBMQyzy46NPQzqiSahCZRDg
RKStPLv8ex6uEckKX6MLr2xkZ37XKhh+C4iCH/8KS1ybGzndgJrh6kYu0xZHMRBLr51TMIAbNB9K
AfaYcyHLetPiSB2qGcjUaTVC3eIRG8GaFx5OEDrvjkGjwd1q9Qw5+/Kl75MYX4E/oagTqD0ayrH4
dju8qnwANM6h+keQV0sh7LzTABfyorHh24fiWaAkrqoVWoEWTNGqYNLF3kMo3JoBCDk6CCHFnywW
axDfV2XO/EKi830TX/g6S7G6DYUVG1cdloGgcMq/QkOPT8yrRt7zxFwB+cfdHgxRP0FzD78NbPNe
RJYSQlcDsqWSg6sFQ9K9a7FkS4uhMccXTVDYOwAR6Qs4thcGYkeEiuLROY37cnJnrX4Pln1OGY4F
9+5M2XGbvfLPUbbhoykR0TvRPaxz73knFIKEKd+OymgQKGUtEiMt8zfopdqUUwqRe1awWayoYgxc
3knVVttCZfyPqyGNPP42Gntj7Rvpl/AYzJEL8jcPlbAIcv5vzIQbcbgyQShnsoj60mgCQqQsxGIG
3nVXNHheEZQzv2JdWC2Ygv6YFPZ3CulFZ/AFPqpQVxtNFk+JwQO1AXFHKAXYHxd51JdvV/Qe6DDk
7ZVwT+JmHfku942Lhs64DFWWzBydP271jU9d8ZxsELuV1lYk2bwAuspBrvK2J2UnDcXFVDm4qG6W
GywTZ70mvey3nVvPgrOk8Ylt9gt0aqyX8DNDI0Hj4RkN/BkCi4ej9AxNglYofyg23OyJaLrDWmdQ
X3TLf2WPSPw79h18CQJnxx3a4TW6Z+PYmCMQldmqqYasr4DQFdqSK4KDGEsS8/uuSbWwNAcuXcqu
KQuNhqCZaONghJevF5VdTeUvxhfzXF81+mpwSE6otCh//Z/w0TVO9u80kaDhP36He3nrOuPRu07E
BH+YzeYeTMZDfuDFOj+xBX6dWiYxIPR1SBoqJNw8sXfEQ97X3NEv8PWXUAcREv+oXj2wk7w+O/1g
0Qk0AEXlm0G4LmsWEO9oKUEFPfiLFIvJGvldanst9jI6lHRFfXjsyNYTTr4+B6Pye1SSv7uAfifc
Y5W4d77+w1FO/qfvvnBYFGcGaYGahGqYHD/aVWNGQRkuR8JFvsex7uc8BGR4bMIc6zCLEqrk1fWb
hlBl5Di9JTw8bdgmtk8PLmpJGScS5tctdsZEKyqrskwcibcTQUDxjfUhWPE+ZZTtkUbzYMyQqLjl
C7B1rcY0TceGGBFwMPKtbSA9u4iIaNpYD/wSTo0wIQhkB1/cJFjlWnTRXRdnOVAmKyqSNO6Tbv/l
aCUv9AtdVwAyBRgWkaVQ31au8bdHrwPegcHf6U0I6UK+2cWVtCuOU5QvSbFxV32kXWzrNmPYUb/q
yqYBhy3iexuDoug2D/X/h6KNPMqZqGs6CzFq//Q+PFkVgAAuWa4rXgIXyl5g7iv4GDIrIbh543Wh
GeFktxU/ujyaGfRi2TOpdESGBz4KETUhENl2d2FIiUDTOJfJq8lb5g0oWEINO14AsBh8cIAWmRwP
HpkmGHahL75dY++lewsLPKTb8yb9n7dBvU3ndYxXnB86bH5Tq+nnT1W8K2iG/BWgipTVuP/EK3KK
vCFYH7qhAyBFqLaEkm7IYfBDZTs70DzkstbreX7uIccV8wo5digvTPKZVfLDcXDGcRLddKTM/7Wu
NNEUENw8fFD13p6eiXbQhVVhzhu32DHtDBGfT5OvUEO+s7MunuYUZTdzfyTddOslFKQKtBgk6ImK
ulPLHIBbT6iOP9Fxrk0JmC952irz7PVLgcyY2KA4zYixuLBVatfonT3Gl8G54c7Y57UKRGXlYWUD
Juu/Y2CUu6Gd4/MaVhnxgXzsqD1MHzk8Y8iMB3pYqq9Hkl4mY1iQvOCQx41wI2JydzOcOkkP6CmE
7WKNohw8l7zBxbIkS2sX3H+ZPWnFZ7I4r4++sEBNBihBxsRSQcrWM+lUwl3syLsAwfJls3px6wsb
OeN1Tiom4S/SHmnQeV/F6Ix7zu7kSBpNFIHU9OkUWZwk+p0SIVkgvty97YK8PZhKZnodJ3Urr7y4
9+oZQXjfxSNTmM5b4aaK3nx4TTS23H/QP93jWXzwyJ4ycYoxJWUi/UMkDr6CE73YOWR+yyG2fx5S
sSSlIAzvEwVzfU4jddaaCoRYemtSYJbqSpY0GsenvWJqMqrU+buqexD2yan126IbWly0uVmAYsmJ
9c6M3jOgqC7oZSzh2lxjlOK0SR9szuSm0HjBe4nkwj55vgJFxlD/Gj91E7yXaOS3VTMotuaCuvbC
hCEq0aQ8vNuKjDsVbo1eEzmZyDW1Wdg6BlnvLlR+/I++EK8lQCodfzS42xBD0ChPb+teRrr8O3+S
7L0jmduAQZbR/7WURUnIDQMjHK1RNsASnVHKaCJ4k2tLTA0VLXXiyTEfHxCAESR5NXOGiUIhtvDy
xPYMTX3GlAHfAdmjhDXnmsckjc1TmAlE67Nd29CvMU/7+WSbhxgUOl220a9nm+g6RffPANzjtIqB
SgT+E3lguoTok5HTgTZa17ulvyP4s2usYclPXamlouJ1a86ccn/x2jkMaXPqPV9DZ0GLZKgog/eK
MxD4JbIR7NV3+jeA/aFaZTyaFzsfo23Hkn7gmb2v37oMBc9dWtsHQl4TAGGT50LL318JnP5UU+u7
0/dw/IXpHihSp4SqyjHaAOGqlU7HDtybZFSC6Ur/qjEyXuPBvzBo72rhmJOC2/UOz4A6D2AGq12B
Sf5nBRODd4PM4H6ooF6yJy/owSrM+/Mvo/SFrKFSxJxSSInCyDcnXVjbGQU3c3yHEQeMYZFkP+5/
I1hqTzTh+Yk0oYkSUtVc9DpBLg8bjMfP3hKbecOq7UZ3pP8j9Qz2/ovbTTCchLcWMBGA7ll626IX
zkYJP/J39NxQJh+ovK8Lqcb9wXQqiGhwjgLmZcsnro90SxinKLjOZKV3EpltJlMXFFf9Yx6TrDSn
8NQltpltxY4HvZQ7vlkg1Zy3x6Xmw6IfQ6UB/yrrV6ZE6KMEmKRaUfzIsMqVxL0In3UFkarAa0X4
0wxox6Tb5LrzvWRyX08VqK+LYkdXTSldpQ2mEu5iQWCRmi64gpBChsxAcyGXQ77MysxKk5/ut6Iz
xeBy72DbQ5Tlce6v2tcLflhbAOBkx78Ln0X8Pi9s+1r6ui3nsQdYQcif11YsowGbytYG5pWWlSnF
rJ21wtA1CUYj8ZpJuokEoChwVnOdRHBajtjGrxEL4ytGy1FvR709uURUojqJafktfYSWNwQbMZut
9v4i2Np4WMNRqpCD00NiJAzmNw1LfeUcIILyOcpDbmrhgdrPtC5+fuDzeS/UC81DqdTu3/mdkKSt
UixmbEnmdMrR/6DKgv8av0WF3tMx9VE+R7isaP93q6YoaYJseNjh9o9bXzspK9OWrL+5zp4alXBX
VLfsX+oAevUjEV1YPzXgv3bE1yXhxJ3Z58hXMmYYhGY5xHFlFhJAWF4QFXCLm75gLImDMc+dPuwW
3TfIrGD0qq+T7ZZRmAL9aVyqWf47ddwaC05PnoTxOZhQiOufv9vsPFw/ZBbHJx5R79LnJZydCGuO
7ryvSnzlHHZTNOYiVWKVanUvNPzXrfX8MHRZ0sVFYMugncYYSzHO3S9rKUsbNPGC1wQfwlyMT67r
4Klb8ZzVb66z2/G8M+HLQ1c0R9Sn51h0YTjJjtbGd29VPJBYJRxzFmEFmGTrSNQ4pM462lL2s1um
vBfdNsLuSBpaY5eO33Xz2Syfu/py3F5iNzpWX9s6dDL7a9SSKkfJ+WwQopVTrREFyC4wjK/X250W
ug+HKoz5LUZEtq7nldVq6kjMdfPcqGqCmsM0OOpBfLsxg7r3LR3HCv//RdH840uXgZQGU+8SWbIU
6ZI2gUzcVC9uQPoYanI1Z6W4jBBRIhNP6Mu7RtiCOUjxSMtON47lN2raWf53CNGuDiVp8uYqWdzh
Elnwh20+zW5Q/KsUfygNXvejw9O2wDmmlyv5hhkUUqHmrcGqpKAjbp+lV1F1O1zTuxgFkyKwStP1
KEG6hv2YDw07+v4nLIvHpyM8VeiyPfr/5iP19wXZXhEmnJfS4qLEJ0jpcrbj2QIY8gIOCz1Rmwoz
x37sBDwNLa3tdg8q81M9pXI9NASXx8BC3aVr3HL50kK3NhIoh1kNsKJr79VZ9hlfw8KIep5rsfhl
xu+D2Xgvccc9mhNbDB/omCAqwRRpTenos5qC+D4n9lyOnexW4SrMLmeOyJTdK8NRG0wNjIPddZtT
FjMZ4/60OtWjt6MpgdYg++TtJBbFKgurPdUIcFQPUBpzl1GmCLzzlifwwe4wuRuxvUyPZMI+NO3q
Aa6NKNI5AvMV611fKTa0gEzPUVQMlOXLbSfPLReQ8WinhhIpXojzAbf0ED6rBfDAV9s8tR+JeWit
4rN+20sG9NEOBnEBv9Mh7TLSfNFC15ShT/V9EySScFh0NeKjJ4e4rWuefaN9ERDc+il4TV5RAalB
DmAc3kOB1Q1yjxFi/9/DE7A1ThMrpTpfiuVCJbT1bs3/fixSeKK+j9q4OR8qtmldRP+5pUg5g8vZ
D7NMsV0ta48xfK6j4DV3hEyvltKlRZX7RCFB/U+p2QBWxJtIgQ+mOqYkLnUyvWMdsQzGdr+Op0ov
LSG81dwFMzeOY6qpedOkjahOics0whti1ls1Ww5a3eDFxn+7NclluC3PzMD6m1Tie/ghR+NDhr80
XctvaVj+YejbXYlyK1VCObwlPVZ8c3qsk083YlKkQ3FghVxdcM4TH1sr4ST0l5Qh4DiUSPZdkYtz
XCorkxPjEwMQf7VnJV+FCH3ZaAZXfI/NjI26CdC8w/JNTMarJ3h0DMZcOy/SmbnB4AH2SGJb90V7
hgeZNaAvQZNgsbvRQ+zZrVlLrSLs8TmJo6O1Z0cxw9vvwPYkjEo51NmsrKXoPz4oNzUGPKDqqZJ1
uMwkeSqYEZhJq0qGHp5gNXc0Ci77WtxE518m3NhJ+ZM4xE80+WhijcB0d1qKl0JtdjySNFmMuYCt
kFnWROYk6Jry9upfgg0Jq7C4A8q5P/Q/cdz/F0F3QVRWY5k9jBMmguogpwjyGmZhiqPBB2wCJoQR
qqu5H6K2UwxfBFn47Ckyu1bBt3yJE5LO1EpSaA/ruGaiCiRfhIP5Yjb5QpcuBRhskr4HKRu6XJoT
3bIVtjQmBpE8xUP5jyVKt2kk7nhsTLEi5Es7JAQ6Go/g5Cs3v2ZNt9yCA8i4EoZHAIq3UXFzwS+8
75skN5UAj0REvhklBxfM8khw6TJbYoJEW7FlqZxXpL52t3t+jNp0LIk8PSBwd0syb7at+5+jTNL0
MQCLgxUlUraiVr7OH4mw1HgsU9m9t/N0X9Oq3t8q0qTLrqkBQguvTaJcFIKVYFDcYRDu+n4S2P8M
GAjXpLXftJeeuQ3Pxsk8cMI+snutkynowFDPPb3DExjZCroIiyDLzTcqZsF6fBPETraOt9G11lZv
SSpfsqZ3IxDaP4ujUCh0h/qB5GTk86e/lbGOEEGeoKJrxBue7hhQ/N2wfaRWAYNHe7b6VjZZmPtu
FFgApXHtZf5gut45IK/ITp6SNAWO0AyCb5YOavvmOnlwh4leFaoTeCFLvaRJYQgW6GdoibKca72a
JxsSv0u/zCYgljnhsDEd+yZ7vs/g4m62NWt01CIubnUd1C9FsJzjyvNFURAJUnHiGBgDBd3sj2NN
QrxevKV4eHJl/+IxWQacWEXIe/zUuxglGfQesuxZVO1zLInjl5CbO8KlWa1eIllLR6qE5ig06t+P
y9m4Py7Io58CYQW67OZke7TaI7tzTP3r465v+0bDicKPS0JURnDd3J0+Dc0Lcdl4ceiGHXlYnGJ1
D1QL9c/DdOffyW2qTWN5hci8XxEtANmTDp3nFKYeHoIpwLVBQHdi9iubfjqjpKQlNmjShboSPSlO
KM0Fibr0M0u+/u4TOdyioSlZlj5WRR28erKj6u72wFuS3EGFcspxG84hsEcwBVq7WexDSilDt5CA
7EtlNTHkTMW9FKnDErrH1xeTlDV40gor4fiDiadL9cvi2GvsOHSLPSEVUSBTB1Clf8ep6DRuwQzi
bStEIvghvlzeNhX2hEEmymSkYejVur9QgiXBFWy+U/myj9HbYON87wAfbJXqzRq1l+g0G+N2TS07
877zO3dc5oyOolunZbj+sH7mb0u208RamjtoyBFcsc284WbO62mComu/GFqdc1Kwi4rWWrjmpHLb
gLaEnBQSAx198gKjxl9Vqb7Sv1HWF5JvuXlRO5SFQ5LRFJAPMuWJKNU27x+oM8UVch/jTHPQR/mw
trVn1lGepOFNjkZIo2WZu8I0XthwWpI+j7iPVfGlF+qUtVrCUEu92swjmoaN0GZG428dLUUo4kM9
SnCHgjuPr8cAl9cqMfz7RRkLjW5ODIcR56LL9kstoV6oYECTbMFsi6iR9EGFsjoFnO3pcjH+kx+x
8gth+ZxzNNguSVtsd1eyk6t8xPHdA7MThCeD3ljmNRBZ3gzSD7/1WeZr4cXWOeEhjNLQcpIBycnT
u/OS5lbFL47P8heGfqQ6aODvTtWlhM6IZCJx6vG1vOfMj0ejydR53Uqu8SHttkXmybyeP+m3PyHf
dYivyMnG18VcQXci/zejNzLijM8u61nLsTzQ0E+5Wd+UjX5HT66z2CLNVuFQTEO6GugQPjvVg4A7
HxdfLczmCl+dG+APKJU5wBaU0tAY532IYeS7+b0xdKm5cwvC7r6O+f3esDzpoZOu7E/LHRlRfK9g
tSXnFpg1I4w1y4RGHMEOqK01xDfEhnslvtmmW8tMVOjFQqp9RqCSaRbtKVZ8U/yNk3PFCr1UCvbu
oIyjIGHocWEtTg2SrGFcn4utR8vFocpO87V+cON1iLKWKNJ7eGcL73ls0/pwXU6Lz8pbgMeqaecw
JEVdDarPCMSyTfo8dUHvypzOyY1/+Z/DxDtl5x+mgye46CWEHDletFo81TFitpatwT+S/hFpdUBJ
l3fMO8Gcsrz66I7FfQmIvBf/mBJk6x0bFCecL66h88iGH9vol+cLORx5oIkYY7mes4SV+In7EDC5
jC1+BjDZcHkpx+jmc3VMt9gJsGbY6ZzdYaIs/KB9Rfa2vlkZfEcn07QElLhcSIAVkR+WKBXEv4Y8
mw2HXvf61ws0GESbJN1vLhm63gy0zWMTLNYpISpYEjtSqTjXL1bohh9uDXYxft5Iq3Rq3mPglARH
qQUXmBs49Vc+6ByUa7N6jfYr2uCH/7UySbnB/JvI7LMMvTlImPlgkDi0u5kpPRTt3ACqMuS6wgF8
BP4EpIceTeqHEvqEHqgeMdAM0VVFR9flWCVv3bITPIA709MJATZsLqjelcEnvduky/CvXi80fgvy
/wan4e1d5QA/GLNrNouirIeUObLDDHv8QTNIc1gtqa0qzsCvHPn9BqqK/TO9fu064q33Epk7UcS9
CtqV/ujxT3TMe797xMWkem50wnEQezZDspi9Gc78pteqsyjY8KbTaWniJYZc2iFUZOfZkqGf4vwv
V3Hl8pARPZCVN+URcH0DrOh838lV+VLMRNYhB2t1jK2xgRPA8Lyh8l7xocsQZd5A+25vxjzZXDR5
kAFsxPNQAkIaGd0xINQS3WQ4jPu8iAckbZJADKrIeOJjlqjjxZbXN+GbsAsaDgTsmEVAHnRsypcC
lISbCBG0/yNmfWEAZ4fbOHL97FJYhWfBnrkVVXml2+8yiE0rMdJ8ohtdrZldRGsme38MipP6ZLD+
lzWBnPo5Uu+WLMq8Qp7+BMFwmk9jw76qWTIUi9uoYyRadm0ZHldLLUVqsnEHX6OgylbVJXMefCb7
KdULlADx44HdFn9W0aytPfjHJJ3uoy0KNFR8co+NLTFbor7SREUP1Wlz4s0jrArDkDbhCuo379PP
J8GTXDgm9eufkP2Qk314OFHgYdac/yfjGq6nzewmC+LYTZfEKKbjyoNuWzw6bdEpIkdgLF7Rhvaa
m17brhiE16kYLRRyVQfQJ7XKM5jg10v77YJB0NY6dMwks5Dh5AwrgIl3EJ7iuxuEG6zdBXi4XjoD
EAfrtVTrX8QHcryKZachS0FsImZJhJsGwYVj35u49Rji9kXMzH3fh98zAtVbCFBGlyNmr4qemrqm
u4KNrfH0LT4DLYXDFWEhbZxB5YugDxnaYRDcxdufQ7+wnuMhZAIBvLHuam0DAy+St0U6Bwi3dM1d
MQgY/5f1noM5dNCNMq8wg5aiq5vnPjteHig2vTMnLhCjiRpvfeWQfxz+TVitZGlRl2bLzpOFKIdu
TPJNJZtfYHAT86BaDFlXUwdI3p4aPPb0B0Hfn+DNXwVtvCLcXlxO5RnAT/8BYxRxEZ9GQhpMlhvl
IVmyf4p8CFEMy1VfJkXNB9ioDKp5ef8kjKNL7lLKQLRehDeXx8Zo5mIFLTjGhgnsyM5K3YacPXWf
3lwDzGMB5gA81gjMXCsDV/LWZ17jTc2xYz/HdtqV/TLig0FplMZoePZE3+aZ1ebSUgeEbGe+NmaD
b70tjQ2sxhGg9DFmV+QzqtRHYuVU4ihTWEoJQFB0tm7cNipn8DNpC9EWB7Q5IYhA8kEMABJNvcsV
LVBuqL4An+bMzu2crm90w1cnn3qkgbqMNBrbQ9khVVzcJEz2EpD6tmqnEsrmkvbioXJMEA0Ag0YO
mEO+nLfAhvOIAD1c/A2N0kIjM0gBfqbaNostiCXtaucp5uBkOvDwO/gskFotA8L6+KWCxGH0GJTH
7xp/7LToecxrLZSSsrLjxG6ZFA9/MsMZN0sOcM08yZx24PfE0c2DbmcRrDEE/xzSr2NPda5SDvaM
qp+IhoNpjRfGOxYlF6jV8DC2ntlrCl2kezYc0UvlgJ0lT1+oTbQfBSMNp9Jzt827wgQwd+gf5uI6
K2URsl6/TgnmbR2RjjV5aJkBwI3QQuXyiODYksDSOBff/Qu969Xkac3oB25jXAsgQBlOm17nGDwX
3RGTFoLB2jLkJulqnXCyt36vdqf4uGn7fYaSpZO1OB5I9IZ8jk+3Dvfcjqcb092osukrIcEcl7xj
3oblm5PWZEBnR2fb2CIBZxoTFlmCvuIshuEFqup1RjDAy8T0SSW+ycweaZLd55A10LMkDtcid/Hv
COZO+iry21Fww1ImFtW0kycSLVqKqiJB8UAdDFTLIgB6celtWiLxaZGdE+UntsTBKJqL+xnRBNJ+
Kn9MFqYj4lZ7JLciej+xUZUTPXdUMLPZFklJSPNFCB17yJw0eRAIL5OBvHYsh+EWjY0tIf6ivATi
4eobzOL0mj6krvXOJWGwNKRvcHYINYYS/xunDK/3oJIia4yDu6JeYP2P/Db8cGBWSl73TpiGFRrl
tGGIo6SLsYa50ERYGkt0JxNJgwOcs7NAfm0SzcGb9bb3hYKDefKx+59urhTAVmPryGFPehqgO40A
Y9Yc85q5N5QEf+bspbzOng/PPN+1KpnVhLg/Wc1/iS7H5p/X33usPR/OEn4X8KTOKx2fPjRzGTZu
EvWryDjcKnVDuEv7WsGB/GZOAINSydAvHw4ARjRZU3Db023F5NmR5EEVcnys2193X6nec2UCSPrX
3XJ2q5QbAdsm82nctNawTPRSoCfGuxZzzjMmfPOAXZrpZIq2FtU2rDR4YezzfZL3s3HOZEZWzFhZ
wlQ9161g3gHMJIjW48mybHO+4Fj8lAZIAvjB05cemSR5ENwd0Hi3H6OTDuuI9/o1CL4fwlu5TLe2
3ziTKC/NwSb8AihwASXEtObDlWed7G24Z+tslD0rvEPjGs/add0R6AV8fWne+/y+gwwUzcwdNaai
IsiDcvLqalTyoe4TUKT+aTCOfB6uQ7kRAtzrRUkbvizEbY1Rlm/RdpEq6Z0XwwbHy5BNT4KlYsjb
SETnE9BY2DqIeJ8sZkX/Y4CFWhKirQ8fEE5YbkYEkEH6So6sHK8WEYcfdvrNwTwjiEd8LciFxjMO
6Pol2jqPDy0fAL+A9CDW4WxqvCjazbDFJRkpF2Ce3yxgJapEIxLSxUbBmbjBB5TmkB9NXapojB5i
E1+g2ZGGjsRRhlqIPMjH0dk1KsU2E95MvXhu+hQVdnulLRC+L7AnSF1ResfnI4cHchK1AE/moKnU
DFks85pyj6bRDWXH4Ev2vIOwmCyMabU/fAukxn0POSsHYW6IXLW27hj+sUF7zy1DObt63ztOW30B
yqM8ADl6ot2irSL7zbXbCb37ueaEH+avIyADRs0MOgNy+QaQX3dmsXqB81ERsYgFv5bFZn4V7xpa
sMsN3rIH12uAoC5prZS5gK3VHcPNqfI/nvtXVrPvBsO5qSOpaV1sMmXhmM374KLw+mdMtlheS5pT
IFPXJN78I44N0QdqG1CYjPsb7GV6smUF5L5SnQF+gPmFWMSQBw0V2kE/ZZmzvUZhIu00+0QpA1fa
N/sgArxFvHXluTFTXryDJWQjCAA8wj1Nbw5h03ySYXAm/+0YVBDT2gaQlH8QhPZOPBAy/wkZrOfT
FczsgzbyPoFsK6MuI7qSJ50G06c+bVUGEJxy8UaLdUFBM/2T7JjuorQne5fBNPIWRVsx8gj8UeAW
G0Srz7TTDkpCVC8UH3+mPBg4yxj7uA3HlLDltAwDyCu1E60jHAadiwixGY7XDP7q7XuaHeziDaem
/g5L1BJeK5u3USR13WWjAnKBurRPCZcf+8Ze9PZCpynMrtjiQ5R+OKiyg/5gMXpe4oCid5nSu1f2
oQGlG6PuocxrDF40Uym3JNC537s2JurZke84PVWkGmoFd8pdlyvricFztbKbdI4S1lXt6CEidPUN
j+yYhjhlaVMuNhqxMPhCEU0QMrh7Dik7tO+3aJiJR5CC8qkcWkA33Z/vgOdwoFEsUBpFFgGc6HhN
1vgOWKp5V1DqP+jTWOH6xAbhkpBKvRxTsOhi6XAtU6wBJiBcdkDtMz9sgBywj/DWOi8GB8rmfg2q
xE0XB5SnJLq/+v/nffZ3zTfC3WoHr2s4Jek3QG4X6VFaxAHpRbfGFHvrWBvShi4Uf6cSuoQcOm1w
/cSZUUfEk8HIvhZ/YSwJMwwVjmNm277WnEckrKHcS/9QULrsDCcblqGMpJpijzEQrri3LCzgUmV7
D1NYpozqOVkWBhUdlbVVYOgtxo0ldPYeOwq81VKhkWhWJIwzgGM6eo42pRDuRREJWE2pwudcFFrp
fWSY7JkSvx3z+z7tgBQNzU1qWo5oPVvjJpf2Dy4uuzcLb1iE/FFkLNZEbpCQm/FPozFgKrU8NbRD
Q2dNwXCa1qVZJ5zH+qWi1Hnr5IeVKdGWifRZ1xS0tMlV13xFiNl5LFHX9KuomQpt72eYTnscSPT6
nyRBwWU9bDI6dTbvC4BhrTBK167oYQzbCUjK2qNDlW5SQwEqdp9UuzV/4TzzPCGB5Koiuh41VKMw
XbUfkNXg33K24mX5i+S5IgKv7rc0kL4J/0YxKy5weHNhbaxHQyPZfbYulmOAZxojYTbYGDXFUzkF
SdxRgtw5MGr3/tY2auZFdycDfT4FaO68mTTZQ6OSEtEJ/CuwGmIn909oQksf3daQbS9NP5pxIC+2
LLUS0csy5LR5PTmWnqrxkOCvTbGxm2D1aYrHOF/uzDKaRNT8RV01f+zc9CAolONaPBa2Wjcy2MMI
sgfA4VDAdpUD6ACTH4leN3KRdHqwxwdRpQltmSDkiArL0ku7ReqItGxp3OMGqN1ADw36gtBtBfH7
NJdodhKvbSW4jrFCfSOv3B69lES0OTtzJWmZ+nppq8Ano4DXxS2ms6pblW1LUX4XrZVJ0IVt82jO
O3evKfA1oZzU/gYRk7mAfBjgzNnm6WNtx1eBYY5aqnN8RcmaQIFrMtH7b6GXngECVsSetsqS6t+R
6JDHFfA8B6LDP0YylPPQNguwmv8x00jgsT3HavKQl2XY54EuHLI2iP0FCS8K1JMkiSHUXaMEBEo5
sf9QqZ69M1ccMBKdKwcn2J8gUYxiLGrAfva0jmoIvpcTXiqGveOo6ajaUPcSAri1IvbfiWy06/r7
Kl7b6LOy2Xqp/Nq4JG4KT8gtRGG7iZ4B8wl7ubKzC8N3LCcbs/AhLMv+kBlXT+AZPdhSG55Bl5J0
lFfghylWYu5EGzdqb28N8EAqCxD7ws4XL07ZyRtCASwO7rtOmcz0e9O16tuDuM4GUcmOvQdJtN+A
mIlh15F3Ym3AH+346TbMIU377J0C1npuuEj814PjokI6Vd9AxzMfWKlWym81HRRCc5VdtydKKCri
pMBlKciDUYDy3CdbzSSkfiktFKJMmjKStofKWE/sI74jfE5GOtKGnM3IWzM0u8ZyJ2eR/J7uf9Fu
AKDuUH8sby22V6kZFJumin2Q1mLFaOM7VOfLSO3ZMdVJGUbM8k/bTM3l1F9Y4pKmebW+VT4IqDZw
3jrRF8mTtT/4VooIeqoBdBWUegzX+oy4Ur8sGnObKgEH6/DiHTvOnkCH1uQxSP9DW8xHlMnKzYhU
Ogl91dvJA7E+UnLPT7rj1ZJ5v7NznYkIrVNseYmKGXGOi/rzjpTO2aU5vcUlgaOszjGYK5whPThU
d29UWU19Ia89twOJMNFr1+ItFdwag+Nog7I2mmvHqRtunDam/wYNUGF/FbFgfl4GaOTbXmzSsoXs
UXLb9k0E8a6P3ktrzuOmke1yovXhoYBXYUovsYkL/PLJaF9AqrvEWSQMmOqrstDtqsE/ISzynfkF
FrZrvrsRmZ2TDgvKjZF72dSF0AiVkh08JwAZQJl6/uMmbAOqOMV2qvyBaRQMFWlzZIC4MnA6qo4z
hPTJe9/wpEf5NkIaDBdymMQwd4osWfznAEU/Bt9TrSiqBDzgU2PcrYHkFiSBO54t81sbH1XTfVDq
KSbpMwiJ+arODHUpPcOy8daY3wJtt7kMGaCGUQSZ38iAszbETXCcuNtRAGqYg5DQTwfjPt2ZfrYf
ZaLW4KXLL0QffZkZCRuu6HASgaoy1lLDm44y5BZNDhaEuF28gOeaSPkbYm96D94Dnp0bYSwSJg2p
WcHkBFJ2tsJh2PS/Ew4zDOtRwmZlUYjuV4Wsn2rASRTnjqXPR4OFtG3QdUPsdmuuOUvy2aBKit70
YmmWAwYsSNz+YbhSNhi0p3s5Fxm5mlhZG+emTwdxbO7wZDeqOStalHqZsW30di0J6KHmAlmXq7Ad
WP4fQhwHZVekbDk6/1tvyXfhjxditNcgVIjTrtFdSC89KDgXiY2C3gBFV2wopI3UNSOEYIbzAudH
GP/lC+zBpeavqAdstRya8mdTZ5iF1+fJRS/uS+sQ7nq/1QIUn5BEia+8csGXxf0alyv4jO9VFBu1
EAHukFccQWDsltewqUt3vuxG/4q2PWAKvfrUHq8c0oYP0kcfY/3UO3tWW0kS8BDM0k48xuF0yFlh
HIAWDkGjp/asTemUDnCY19F/nPw17mFkdjsVw7+gWHXnCs3IpPBnFQABxAR/kmHXzrr9W/P9SELR
5laT03E6pGwXgkowGIqExKED5PAEHGG1GcKESyBn7VXfFBX2nWqRUQc4rClgZpy4OxGpp6CcfZIZ
brgHAiDCU1b/prC+lK0ia0pp5SYQqLisdW4kSFqFfOtAJdLaltJBclZFDz0H/d5DpHkVxO2dqKcr
efi3dlPBYebldYaFATLWuJcqnLEhch9ieCeNLrev/txb8yjYwORcKnCmT7Szj5IaPiO4pup/6PwQ
Vk5VWXZueU2Ycj26dxOJSGuXCcwoe5wRjFDBPmjcQCimCrNGPnoK/wpB+tp7uS8u7Yw3SQZ+aPaE
4LQdtNbtS9PClyGtcarqFNJK+adPzdCZ+GWn3d/WsZGLI1XPdQO0iaQVREHFa6CFEMMhdpYtkkoC
ZTJ34W6dL/NDmWf65B53DI3/SBWpzyMRrXHhBjVLZv7WdvfKYbmfj6bGlGpvlKfesmJ3fx33IeM0
zHc49NHMXlXCNzMP090bY9bDw+w5sgz4KRqcKQao+iUMa+dx6rZEUzy+mSCzMJ8XiWfcsIaLIZof
R8CeZ05/uV5KM3yWJ6vmgNDOxGvCXXPzcpu9ys2tBeXVYYhuxpSYRHxzW3GwAPEUwSyVU7tG85JO
Ei+oDt+CO8EZiNM0PD5Sf/taw7Si3j/GKkgZVC69dSOiZd9NCXcghOw8BRYxvkPoNdEPVWS15jgi
l57UNirF/VGntsNOGmvHXM/jKr899MpSd3cH1He2yHEjD0ZcPr+iPCd5VkuKFlKgVlyccWqIXJmb
QXfMG7JtQLkgy/UbWtrSFpuctB2A78JR1rsTVG9GRrQGcB4djTNnQz02AphqlzdS/8Q7k+1CR9BY
cpu7rSX0FYySlWGkxfe3OZE2pyJ/p6cc1TDKsisxLypo1tiZmyTX/h7ReTuzwRNaULlTE4qlFMAn
nbNHW5LuOTnpgvXF8Xx0D4EX456U5mLCqPTogHNkv4+O0j+KY2O3dPS2O/xPPjNyQUtpscDobM+f
0dvENQe5bvaIQmUYQDgE7R8qjV3S+qTTvihULBzpd+T8EZ4/JbOs13ZFA5zh1NOc1Te1b3v4TBeb
FhUy4Jad3i7a19JwROFlQgzazllZbrdar1Q1UerO7HObFmEGSzPnb8Ak4RtYHFsn420V6ZAr94PD
TV0GvNt3/H9CPoAfkz88GbeyohhGGv2OKfZF237IYMVyp84W6P+aUYQHlr0CBqLdyIs5FmJy+QUN
qGC2XywkAlQal6R/9Ugf1ing3+4kor19JEABXgF7YL+Y2LeJKEjWOcTGNvocAWNoA2rX3jQaIgSH
mOmMiQWNWEUmv2hT14tDeqvfu87cdAA1WHBtOfvc8cH8HLRlVnBicwFAnrZc0w3Y1HALKARQ8Ezl
y6I2KUpmkXXx28ZEh+OtUfERdp2evX/7x+6erZ4vuMa7VX/hB/NmiVx6/k2ZjT4ngJ6uBwQJU+GM
Q2J25R5ezO8f7iOJs2ll942YUC7xeV+Nw6Q+O7CbnsVs18+ssuYkrv924KBRMgr4lA1HDU7c7cQ7
pk02Oy/MoFiPhZDdJLONRE9YaRtugXCes+dtoKSpjDPzCe0aT/TKX3p+3q9isysLqsfzN+y4Zv8s
zRirqQGb9KeEwe5y5IPd8bUWlkeOO82e04neSt4xBL0Vs3IvnSLYMJbJPtKEu0peEiYg51iWyDcv
VCZRmfoUHSNb/7501vS7yUw82s3MmyyNnaCeEgbKGUHpplJg9+138BAM3vH9uc67kiOl0o3WdTs7
8dpsoM0by6XvZw5MSrq3Q4lSng6lt76mNa2bzQQlkeolwX7Ac/fZaQbaYVjknQM4luTfFe/yxRfK
zy5s5cQ3WKwLz9nq61NT7fRyaEHW42Cm4je+b4MvBeGgfK6hgzuHQWzB6+EGccp4gvP0h+dbqBvi
samqRHGHog4Ntwogm/MDPYoIajsuKMGP7p9LnbdQxAuz09f7TTjbqj3EXWHll3clVWEhGm4qKCCT
2SdIgCe1p60xCywi7frLQsLNDgdAZ9SqcsFe6Ndh01Fo4F48XIGHdr1dgT4cXQYxhRr4IMa+B2vI
b6jEMUR4TQ867giBaA7ucF/Texu5C0YPE2AC0hg2+rslUcq+IZw9rmSJnRyhf3eGoMIwLVxZF4+H
m8x9fNGzNVKyFDBC12C+pA8MBqJmNn5LvjFeCBuHgM+7D2A1axkKzAJg5Ahj8FPZg7jxSj6OXioA
2FkN21+lHHvwYIPQbHzAlgYuWYvJ12wJDpexqV+8jvgs135j0WYIRJVXbIB3rRegw8GvE+7Ty9ah
vR0YlqptPclg7zR8yKI2Xu9SoPZgb71/aD/Dv5NJPj2j904iGgQko1KHTIKB/JBM10+3dDyuErX7
ms5+ecpygSTxELl7IcCRoPn+vWl5P5m+ydEeuDPJDAtpj4b2ifPwKwgbcmQ+v+wlUruSo0GdLsj3
zTx40XMgLFvorsQep/07PJFQypzN9OQ0u+MgBwDJkBkwA2XpHdQrOXwSpwvwWduw5eG5PKEYyKq9
4HGysA0D75pSTQcZZYDhb3RJnfCtnzYVoi+zu6kTjkHwHyXgBrbUduYqpk4ZTN/jOBrZXPW1/0dk
gj7tiMb2yB9B0x7agYpRObZhMhhPFUjQ6dG9kcVPrBfsTunQeGv8HDohPMtSkEZrLMPQd5k4Vifo
TZxVIaNXPVhPxhUsQvJc6qMJ11bZsHgCp5NN+xn3wyY/m+tm3LThvbMtuSr22Rr6RpGlk80QwDg4
0+lHu3EFxfbq1aqEdq7ehWu/KK2EQ6lUu2WJHc4ufJWr76M2Z0beRqexBx4JkHCVCEAWMDGb32ge
mJEQdJGICZxPoSwOpZn2Nop0YL1fbneCPe1e/I9leWo0mnaeYDEJ42D+eEV0lsulHIGxMeaT+P3k
jUUIYDNSQPsps9yGUA75QLzLTLwssQZWbyrcp64HU//recilq5KSsMAuYes+EdfyunBlPiLSNqln
PWuWUI3z4Z5p0eXewJvL8FpFNi6ALHS3qt/yLWijhrR29L8hWVe7q/bMthfTWz9+5JnGal96eWGE
bjyAd5JwfXU7QxcvP7gEz5JamBLDygX2AW+Ba3MzN5x27TyGRwJFiwDMoAgv6DbnB+3w3cR9n/5/
ruwcW0eqgfIdGQWnzVdqw+/CQENEJfAhtApG7HeepX+xlvvizdSsOm3LYY11yuniI4bIZLJVUbBY
Y7Bx3U+z0jTSErRoed+dLFgn86YHqxHCYXedWZ6b1tdFOqDrKI5vutZtUwGxZ1NqRxUjvsFSmf6v
7dINBNSWP4cjbaSooj8QTF6TibtIX7KAf32UrtKQ/ELASsW5bdKTHA0NHyZV9FVe7Gom+J1dnfLX
8EiZner7W7sCdOwfXLxIyUSabYsAH8JLZvEGUklYe3Z4gsgoR4PfBf18avkogcXQfoEHFTkFmvNa
xgwkMeW9l1VRzilLPDeKmMwZft8LlF7+xDOnwmVaRPFR9SNH2Sy/q/yTcFwRY7MtDHpu/4rVDvyg
1f+wV5XFDSZ5jTRT0OWuzMtYBnC25MAgRtBgklYL88E64YUmsFL3LXowE4mrdcsFdv32Z/3+5ZAq
F0X+4hSB04KKInBJlPh4nnIAVC7009ffxBj3UF+Jm2dtXDb1YsOa1MuXyZUpDRvDtiAd+/XJoxl9
jsEm0mxSDBN4OzADSR13n4xFWckEVE0AAuBfPEMujbCsbp/pNj93FNo6ggboa9uz+1dgv8f40lZc
hRrOkaf9p0RhMSJeFR8EdVsQwaqkbkNn52vzoAs7xXtN4GIfXzbvAPrPjzhfMC3xeAichJT/nXSK
rfMM+NoWuF4CycTwkZT+VrhFX89jQXWKccbdnxnOdUJelRBdkY+DqkvqYXIyo/oc5W15R7msz4XV
391NETKzetsLrmQhWm4XYr1fKBSSpKhFnhYnURp0ESxWmIUIN1rkhs+1roStqgS2FxYDCaZarYjl
BA7xM8QZxo8M8KkRjm3slBG7A/1Hqp+EMaWHaebY+7bF5fOShSZfLfQw67hViooweREcFheWi/tO
XwZE3Xns4Mo6ZQbZ0dbmhE5+oMIwkADxGKJuxY4g7iZ9/RjSSpeEtn8qwMJGyTbxqKiIJBBjpLfl
DToTOFKjKXeafRUtwEvhwRUrzRyN26C7p/1P871OTibu1D7CPjaylwJ0Yy9d3dBTgUY/gVJfGpg+
XFhEnD/j/dwAXBIy08vIEyIsOUSTyAjA8+Z6wk3amHC+CnEnIR97aYnimmyRoYaU36DFWolXTSz0
m80INn7b8LPQFYvOWg3o97/ap1Uv+Tfyk/+jE1FDqzLhZsNMedBBg7BvhUyVNS8v1Wg9xGfMpWNI
Ix+7skkKfHGXppvJc3qcXu3XwFPhGb2rmpb0r4wrXlO9I2PCmk8XbwqduCCT8Pwtji0Vtju+GAXp
3CBFBKwrmZhghdV4Ult0GNw65mxD7rhjbliZ3OvOGobwi4PVHoJdC9/kcWW3i8D8mJApM2E4gh15
Pl7tIug9oBzLuk9J50B0ABhGT0CAkWNhUEEugTvAAfmFqnBfaoteLK7gLKhPDaXy7xG/gE65t1Gu
ACKkBF9CqzO9c3V6ZpQOWJE7crpPZ4aPiG2SiuVLAf/HYLSfjZ1OqlJ9HmEOSj7RqfkxSX7Uw6Sn
5qIJljtzLaCvw1UYS10NddR0rSgwxyI045YuaTZhuTws/9ubaz6dWKCRptM8lwqSFxlKM1YX9aeh
EJYf45D2jkf2BO/8Jqe2BNBs54Ske88qith5M4NSnq1zLg9C4sY9g6hPMN2G5RnG2AzmaK4P4g3+
U5pkGpsv3meKKR9fu88fxRR5EGImG7gfJ87Sr/9k7lCeqAP/9DXr3p5JXVA/NWtY8e6hApa0Y6Tt
SY+cNBGlSpfuYtzI6Uf93zdiUoNG49NCIyE182JsaaVG4WlQokmiHI+cW2lXeto3cvtPsVmBZKQB
K0xArgitvQj/ea3jcqdz36grpMpU/REdY/Yxj8ivzU80e04FS0MR6SFlTUCieitmaf/Czvg1r4Ui
I2LboejMVXt9SE1nwAdS2wkTGqZX4d5/H3V331+R/YTA2k3zIiLhnx931w6a6X49XwFI7CB3EGp4
8JdMDPVWDS9xoaj4nVZGKVc74n8DMQcuigdI1MnYfzGnLw6WlmvW+wnkXBLpf/RyGtYAiLbuvMY2
jM9WEiZGrjE6yJsNB/vdSUSNTUuMCppiQqw/qtD2iOjkZXTgPd1hoYFNspFp/fF1yZgb3jV5LO0o
TCHpSGWNr2pT1PQs6D1Yy8PimYVwqNwpzA9u4hpCl7BKDxK3KCLDcx20lArMCDTy8vaznvzsZY/8
bKSTrnByARjmIOQMLAm784LUc8cubgV0DARhsiCJ72QMNDbdXDgM7NeObvCU1sO7uoGmQ1T49hTh
cQTBYK2HopBHICu928yXYLlMk0NOsndKjB1CgFMzSK6UtPRBartvGdN24HJPkVicCqlyZft0TbXu
KLErccm8vHZ49dt2RK42ABN40Ty3qmgOssUoI5u0xaPMq3ErqyRBUWZWnQ5RnemypQTgG6y69zSp
ec0AqB4HICnFXUvSNwmUxQiCzxi8HCQUTgw9DEHJJ8nogsLaHciM5Jc7++NR/Xx94RKy++xW8rLF
mpeY4dMkasoBJ6rb1wsyO/+E3L/P16Veg5N4RbpR8XyjK2iU9I+Nv780t3CBMekm17P7Yq8Cm1dF
usHtK68hHiSXZcg2TtFajVJBCJLX10c9OYjNPCaP8brsfP4KK4RnT8KUWa72KRrV07vzM9hezUyU
jn3Xd/rp7pLpIOK30bCpxA4i0xSAwb8y7MiIy/IctNf0wdF0stOOBf6QrB+p9rAKh63AFUkMcnxW
GPZsOIVBdD9PnaKGw5P+wY8bVrKohjqHzaG9Y20A0OXpGSqu4ZGBtorlFJBSrKhnvP7nxVpRSxJQ
s52ROICxdFYdMfbffedVVedDlE0wRHoG4qbQ7r2yKUFxFJLnOcMkT6i8EBvM+EmaMHKOStzPJyiC
apHGOyvvy9Xtl9fxsHizhjI/K+s+eoleNUuP7wLbeYqOLxxNhPeylzDGXGIo5Jx7SK+WNwkGwaxg
h6QuTOxdQ3TlCuKvMmfdgIFF/uFVrDJExcJ8DcneAF0Mr6I5Y2ZdUFhh2rKL7UaZ/cD+4BIQrEfT
pfwSNPoFQVe3w2gBl8EBm13XZWx2SaL8W5YLGr3iur83bLJODUfPenGVlZX9mttusJQR5bqqQIXC
6OcWBqibWOlg1eMXieOMfU1Dsjru1LH0p0XC+klJueKcXH1Q6FkwrWz6xCRitG5eU1Rj0Z9djXNe
JpfcxKVUeEkfBRrsvcSHV2kDjObGq9KvXR2Z4SIhAa48kp4hRijkXx7Ol/a6JU7M3GjHFuptF272
8DIsL5HNw3rs6QcKrZzNA/TStdWjOspVpeyBnBUYoB4+CCQnfsIW3uDKrIaw2uljPg5bCmDso3xI
0cvmHUp7xWeNcWes7uhcTCLt0+c71+SvgCf5rnsrj7ijHW1ky/b0qtYIeCyUpR5QmSH6W8yScW8C
UY7qm6SZfUpbk61mvS3wsKXQQvY49A4BABFeSQt2sKnG/9zcECWTOEk0SpLKU0tM6VJgZCo3s77p
4ciT4GkH4Uyz24H4CSkj2UZKCQ5jf8lR02oB5fjz100qDadjSUZbfqxtg8qHL7yZppHCiqz124ZT
pSV6yPW0yEYx8qRJpkQZ3ei5mgsf9HIuMX4EceHKW5pvtRomRcwf2aIcfldpxm/SATf1g0U+OMgQ
KXnJtOKeUUcMNJvrise51YQP2zL8hDQQh/1pSo1r34z10LAcMMmTHnWtLS38grtMtRMll/aliMoM
RCBNQK6xXQJqleQOINNZPc26X+hcR+33tk814iyoY4cMO3C2RG9k7Xweib/6WoGag8SvaueX0QMP
GDbmpKNTSxoADl2Fnzy7EX9z4aE+jwodr4Vve4cA/ibIqIfKBrVjkmGZ0C4Zz3se2aU4Zzh2QKMA
nRNT6BE33YkRCnpTNR9aIgemv6q0ZVaGABXlBdq54gMm+jDKrYnUbbMhCVyAauJQe9+jOiLFbntt
dfmkWZ2aw9BDchOWjwILc84KW6f2lqB43li9AAd/HsTEcoRk9m7FKio+P8IaiB56ZuGt9BbHfBkD
UmqJWamRH9oixoqlUWbdy43dYSz6TkXwvV6OHbnqLmqp2FMJOO17QxogqSUUROIViw1as4n1erju
aG51o6NhkF4hWpDDAYtCH/L2SxmsOR2i//TBeyEFfdyi4TtV2jnht33cqjAGkEF/s4dVeRBlE1fk
UXEKkD2Dm70jdxIPaUlZvCNB4BokBvrPDQv8C6Tn6bwiDo+ZLmVEOeUYxBY97qTxkErWcgfzeXji
P9QjmqLEVgVZI/XwstkkWSi2x2mbTY+SlQmJ1IINMNT0iuU08Udm7Sv3VYMeecfDkX+ovvssXnmJ
l7Sn16mXswoNez0NKKGfF+5/T2e4omC+05w35rIQdl+qUPi3I/58y6yu+Gf2uGMomf+VEW4gCJ0Y
zSaTChKWPtJX7j77FRAcpFLLYEj70r62HHg8t8nnrY48sAftYB6WtqhotOEBcrK5k3r064waBv8o
Tl62dlvAYl+ouYk+A91aD77Xrkx7nvPgF1kBeGIrbpM6lYw1dxhpJm0fb4tPJq9qBVbybVnW0BQ/
WFpXkyvLG5YsMN08T6RXUgA+22VvtrZZEQjvT4DYv5+2VZLuDme64eIQdcbT3XZU58AX/xEj0uXn
LrOtKWiyX+KD+ccg+vJpuUzuMmzFXhhNa+ATJ37rMFSHc0jtMViSKiPgTi0LSq1VCXP2/za1iFXq
45SU5R/dZzDjejRDCMJNkhlqZGge1JK6/cXTzBSoQq9K0YVC0OolQffEui5ozhoE6a6nxHOKkujg
md+qWzRImtm4lNLT5xffbT3JpZnwkwaDnjwE1/3p2kOoi7IpJ3prlaYk0byUh9B5jbHclC3cHUuQ
6JEglu4TTyePRLCquQ5KkoSskD23/M9PJrqqUoUpMHmjI3fAFSgK38+OXAM7JpAyGkC5S2Y8KLTi
4J6YQMcX+OoPBXubzwFv0iWjmec/CMh9HSEIkWWe1MKhmw3qhXHcKAaWUPB8sNr+yFVnPAe4+u/H
Wvpbj+Xb+xFaAJxqAYNPerq8p3lkXKTffbUGDHIBmCnRnCIyc0VhF3VSE+pZEQSTtnFryTaWiPnQ
ypIPJBN8gmDEoOAZ7DF+6Cf/3NA+sBT40wqoZwI/IJFAcYgFMifVokA8zBuB3AyWIu5QWJ/Hx880
SfGDzIhpA728/WGW/Mp3pfSHth3X40dAgTrtBdxDzH+213kI5iVSQTDI50kEZU/jFjfduLYPG9Vy
WJN03xAZs+rJyvhNsKK1+VIiAO40Nb5IuD+cM9UYW+Pzqg8zoaC1DlKz8Vt/Xsf7V/ze/Z9x0HUt
tFeZH0WMKWF355TXvIo3l/2M+v2nFwPouAcMnOLUGOBnVZsZKLIksfyLknu5gGUNlHRcvV+Ue+lp
tsQ31DhPTzb4ACmteayginxYEJ1mo644jl44h0kYSh+mia6XGkskwCqUAeBbDrYMi/0W3hbu3YMo
3jVFFywQxtfHoyPJqQtiSBWRSp+sCdPCIsU9S4lbV6zk50P3GaZUr1McnRdxBwnOYPzBQ1Ceb8ZM
lo70utEQ3NpQWxrsZJaAKDjfpTmJ5CV5kt9xEcCNnHvriheMpMbY8d77vAYbR8BpTUe4kJO2FAJ+
d77OEro878LMFfL71yHnVtjc+n3+KA+rJhFOAydS9ZDsyYf3hg12XTXYmYPWDQsiz9L3+56qT+qa
pKsO8016O2lK9TlTQ+jPmQz51xv40Xb0PAnxvdDCZz2SiEnpBTCQVb1JBpH5QnMomHtwg1tfVQkP
xzLxlEbmwlcCN/CVrNMiyX/yiJ+Yx0SrbfFLJMsJrLaM4OGvXY5Yo3k55Qu5Zynhcgx01DE8dNtd
5u/kdZuxUIdiNGDcEPUait5CKUW02lYUSgy9RLXGzj9rbKvnfSFF1ftq7HVL8JNiliTPvmcZXXCE
lejyi0N1wH3JfDeLrFTYPIDrR3zVM+qMTCZ6Snd0LL455x+B8tQ84tGju6s9nNJkMoR6WEoRCCfe
z4t6Qnd33K3klIoNvx9uhW2v0KKLLDy7K3y3+s5ija0I84iDxoxs2CqchGeDq6r2QTemWGXvvlNk
Scon1YQo9mO1/FJA/A2sjRfn5O6n0TxDKV3Qw0FyqtAxtbx7VtyWNjsQMoGsrxDL0l2qhSeWgVDM
uFrTVN3fqPPH5YGETZ6jiP2oZOq/gfH2Ns7FhxSv7bodmC4ETIiL7JscJDeNPhgsI0blafGRd8pv
dEVZVJr/sn8pDZgIS9MesiDzkpK9BvAOoinD09rUSk8bUH5dFXentIr6o/qKC9owUyfYfyJYEy5X
i9mSUOC31iCXdlxANy4eNg70qpFn+eVtKiJdvbiK2NblHuk1V2l8j0jec8sx51AGIARAOjgrWil7
v4KaPHm7Z4RDvx4sHeBet+HMzqhaIQrUiMPY1+tPvWD8+ikuHrJ8u0jficblmj0g/yaM7eKbfezG
mAfXSgSOM1r1FLx2qEZEK7fv+hEagVxGtk0yokgrZ+xokvWi8LowuUiryd6hBKsRvT7JkGAGb1pq
SQ1RWBETsxu8n8LzMhF8TEtm0asqMUzAAWf2o5ks60zF6WajxMHrD62Xu5I3cv1OVb6YMRNWoiXP
V2sgZZLARUN+kDt10VOrZ+WqNXtGvRyjSpzG0ZJcZj0MxxocLTTmsalvOAFK5JnPI7PGQIGzpUWK
z6gk+jGDQdAL7nFARlQ4Na+A/7vJJJ7/sY6k1c7vgRfRG2Gnf6mQiRFlLKdNwRmY8Z1hfkgYtVBK
niHD6bSgnb0QMHmkKC+0Q5jInZG6c7BXpv/FVhEU8c/atdgHPIrOumodMN8lXRjZ4jz4OPZRIQfV
4JkDHVEzSofmtdgLO7gyJD/wLQwgNr4t+SLzgLp4dHZy2DhkPY+pHV0plIyqGXLti5am/8OG1xsO
K3JKebMreN5gY59trgMORlZV88RdL8zsmGcgEDeFWdEzDxqnQVLJ5FBZ+9mJbf4M5guJ9i4bkIj7
gJ4lvNSDDoE+hcrz07bgtuFyo8y40HXxlVBZv5pzV9JMijpMD31WJTXe3YwzQp+i+6o2Mpfi1xkS
uvyC/LUdT8i0nBUJJCtrmNBnDtHpP5PBCu/c7BSpMcKS+Z/mFMo5lyqtU+cnbDrb13fC/iuNe2iq
YJjhF4lcjO0OttPjH/3/NGUUyMKiw6OqBcxgcGBRFsi/XaZp0TC6xLtmP2KB0RjDYWk2odFk7188
GhrurROiZ5UasqSbqd3LfITdYstXq8hmdBneMjksLjXqvOmS0Qqf+hM/tce/alAIyBRq9mKe4K41
kz02/OPvdm+SMeWTY3MKEUv+7lYpVhzbDcGOjC50Ovq11Z4TyYaf3eHvDXye288eeFUk6dDqafQk
qqUvJ2n/S56nSWMoVPrpxtILeVxw/pdSc01fYCULrD44jpGRMz6OjV+nytQ+7Uc5BRrImPf4jqjr
/oWPleb2QZT7UhkzvNttOUW3kbaM1/aXpqvNXv8mrUDpj/e1YvNT76lUgs+zHVjgZ5NuLX0adqQI
Yka6vO4H1qduaDUStcaPGbROrjx198UMIo/WnUcTq7O8A9d6RaCRoA9gRyy5JeawiIiQk/F7v9sC
qpeo/OB7ULwOjsuk/nyWOQeGwguAgbWvSyrU2nnwYy1AOLaMMr8zHXx1qfqeZ3Fwi0QPasCDAHN2
tsU1+b2kERD6c5zU+FAsvW4ODXSX/xNZ2ndL1KcjYIAOcd7geHGg4/Ty2pkbKA6VBAJSnGI/96q+
pMlJLdH1dZuZHPu+bz8EuckctfdF1HxY1thOQZUnmGIrIRhM0tb75OUmNHK38XwBB9hhJPZx+vCs
44IiektNuWFFPpHbqbQx/6PgnrSKDmjk8Xz/Zm8w32WZmD91kNyldSiFSfhmfzYXsePIZR4xNFPJ
z5C3hur5Mia3xUuSrhxcXyKi3X6wWilEDqXgOyYs/5r76OxnkU4RUw/un40+IUrs8nbtT6kg6gKS
CmldIb2VwgqISOx+9OmIAaOEIW7NEuboB40fq5gvxgSOeJPQigTz2QJvq1UsLi68yUYVCK302huL
77ZyyoYE7QZeCrO7Uz56LcVxdFfGQnw9t+aacBovXli5p28oAFoWu2UrIJqhzAwAc2cuO5VwbCm4
OOBZnzERWJR9fu6XOIyYaZUM6MCRiesiu4uKz8tg8Up5KmABjefJEv5nuBU/6KNCbx7exR98+0fT
we2MPfiR5tAaziaY0ImtX8Jq1txscLByx7iVKCCI+nW6aUKFJ11N5/Jz22OQhRHRNcdmfnlOhUgL
+0e/rd2vPoyvydIPTxEUy4/e2DUluTV6Zo/o8XgBrhhxB5B+vh4h44v2uyL5RSBFy4ACm8Dv5q20
OfQFOjjnkddRCLO10i6vfOseZa0JHynQE2Mu4ZoT9GPRlDNM5CQcC3fmrrfDUCMzWRasmrFqxJE7
5RkbJKDCzCfrzznTQekbBRkNGAUOBwZMgruD7PTKmM8kGoTAVZv+X7zwAkD+Eh0+uAGfX0j78hS6
46gskldx3H7ccFJGWb/pkl6Dd6jKeRTlSZ600XwpZ9FLT7zJ3xnrEq1MKARp6VosPy7ScgnE59Wl
1UY6FrhbMQxFi2mPcsYRKhfqkkY/NZlvTdEGNMrjUQkkoWduzRpZera9KU0E0fDdhYwwmTwOjyrJ
Dscnve/FHUssLRQUA030s3eVg+OGUtDKVnBp5b7koT2qi3PPhmKIsrJhPQiGpNE3aEqtEy9Zacsm
3OhQjCAUJJpnHOaPZEi44gTzR+7gN5R2/RZWtMjU95XBLBJug2ChN8/RG9pACOx8TSGIU7SQeMO5
X/EosjL6b/6qkKWf6tESN15rMsmY7/He55sbr/9z+Gcbl+zL3NXywrctNK+TnsUxfBlMAA+D0bS4
8rnjQzQPv7RU7KnMqnz8sTLefUk4etd503cX4ahO8JSy4sMq7GNik/je9CLNWm6u7K3fAdNwWKMz
ew92W8jDfGML4qOnSACPMfOno4WyuQ1ei1dQq8oVIewAtB5wy117MdZiTrbpA3zMsrQ/k9eHK+yA
dax/09DSUtKANz7+iwu47ZT2XK+Cq6WVHv8bHBlm+YaWIFNZtQQsy+QFQguteXT0YJl1OwBKLcH0
oTqwfSdzNODRYIsEi0Z9xBk0l2uDVMJvSn/Z2fFPPIoN42nwjpEnb8C030h1xTCruUTw99/D+oaf
1nHinfzkEm82IeAjNsFjwmjHzu8/wjZSAJeNq3y8k0XFoTz/JKwF10Q330M7iGJkGTtPwkWxMp7+
Bpr+HQCVCxo1muW+6Lj7u1oJuyUShH/iBdd4/uJwKQ8qDhwZOKtCWY2BBj1ErjZeWKgJ7qUDi5Qk
zYbOIy6Bc0h04ACcsV1MUqULcVdSHpOkMl8pYiZujXMX2DmAH4y8XhfZg5RcJvhItD4ueWSP9aES
eSuOh+dtBLeHL7mVXJ4xPex1vd1mRM/LK6UjTwIGLTlxJ1++WcW9FQZz55xlqsQcarvqwYSyBror
HX5oUPfHJNXTNF2w3GXQsbwtWdoCMCXbAZJsXvNAC/ifh07ZpaAi0+9vRdMKIxP2W6JUV2cIr3hQ
OQXYwaZlUgmaYX9/uFTSCM+TseiQfYnr2daHwIJL+I3+5v0Yp4bT0SbJWEl2agwShNSXD4WTZCe+
TIlwY4he0l/5Q8Zr2MWQaeFv/OVfc7VqwzieLuBx0mOOFK+UWILeqBep0VyBXVrh9mVmMa5aI84H
Va4gwAfvDJkLWdk62Cs0JtlO9Ywvkcqr1Zdly+b07YaBBJr8Wez3lu7mdSdjudXYsqIExgjdGnVs
Nr0HqELRpXIdvy/uMixEEK3f0Iq1zlJfNtD5CwaFj0eeTmKYGCA+W3QHMzIMNIh48iKASSZ/LInr
8Vg7QS4NAC+3YsXNG8htUFeOvzxZlR3jNBpd73On6ZT4EsefznJ+q9YEkx2Vf9ed3V4Bbuj39TOP
htXbV/qCz0O4Rko/DyQKGCWEGAP8ru/91djbQkZy0sVKGN/yUZsta/eBVN/kISRalgbTK0T0y4JR
zhx3gnw8qLNJoSuKQrEiBbLhUdeO9cDo0skDEz8CPxWffRF0YPooWTri+07qUZBQOh7GBbf+dYtL
iKSrujCzILtrZPCOuHOvqGYlIazoEphAiSeBOEw7tBZ5xuyB9ZSi13jGneUO+ImqmNgMiaLtkKMc
83D5bVE80qXyTSbDXDN/10LyOcRdUNJOsuNOLp69EMjfqfNi1LFVWOSPRJT+4KPviLjBdkbgEZOd
ylHo9Dw+O36Xxmw5d5fPIrhxDqtaYGt6aWZ6UX0cB/+GdQOyOSUtqXqe9hmt24ygeYgFTOYmf/yO
JY3Ibz2d39TWbUP2gq5V7c07Dsf2+NNs4+tbCYRrbjDjWVXgRuYAOyhBDs2r4H35CtOHsI0NQuE4
+2LfF7N5cI3zczy4ZDAJJbUKuBzFKsRy5KZNchW+sK+611oiszC1I37ayuj/6Zt7AZWMTHEXb43a
vSffeXSHYVlQGL6QU0FYcGxXfacV3sXYIp555vx0ocEg++sIdKP62eeC5GacoTDFiktj4J75Q4uA
ytR8/RT+sNFgW3wbu2fXfq3F8djBVVayk2Mj3OBHkCFMyLmhbDFkwa1QQWlB+vE5kt8xFlsx5eSV
Cgtq1N9Mw/DkEV6DS6V8mQun57Lbxc7pvy3/I8o9XGajXCHaqpXEtEVTrupYzkpU9mlMtA5lipp6
HRmBWBa8wqNYpkKbEIc2gh9eg5a/1PCM77BHsXIHg9q5CQviYL3DCbJoaUHNLnMhAeWK3wQbXt8I
kuz0fqcHTo4sqSG4w3SyVn1QoSkazbSMQQSTfDK/PrA8SqdXUNdo1Vivj9A7EbY9C6xWhf/U9B5V
GVATuSxlIaG582UMYmvhy5OPXGr7z6VsZvrt5N322KAC3t69wamoq755e6Eh7aN+PnwBZUDg0m+X
Acb2VygyuZQvrKEQbM0VWOEftaQSxYAr/LCIVhcsQoFkRHvwjQNnAsFF1FuGeZ4c7jUJi7cg/V4t
HvnlfcLGOWrFYQc33ayTkI4vpHwF3L6J62zNiZzpx/69/BMkgYjYvPnlZYT6pCXOnNcrYCu8gb0W
AuEavwLdc4zx0WwTVLjxvpc56Fi79FjsqCIrL3Ovf7d4HHZQXRmtF5JtePfgGHuoFIRopS2tSMQG
k3JaZM6sW4Y+HfQrsyv6+UmXyKwRqw9Gaw9BiXDKSpC2UrAS/bCM0F3qVY96eouM0IYAAlA4dwbC
f9a4MICpBduNVmv447Cb55mrtUm2c+6+P8iJVci4AcN8C8wiSTDMfkUcpqKsx+3NRUJsS4EGokuS
V6KRndsgsYjCoxqU9cnYDFTj/mgf3nNOjON00m4uOlF2hTrW6Ctdsp1Ak/4NVdOqmwlSHccbwTNW
wzBQk2Jiv+IxqNFETaGTSe3ON1SFZrpGAUqeI7U5LqM3ugYjqY/38DP0kJ05+Ww6Way3T4ziAtS1
SUxkMpUBpGzFpSZ7ceP6s5RSeBlUnxGo2ki93U0Re4v/PewS47AsZiryrk6bQ5QFxydOOXv73YCm
WMnoa62dpemZhrD5rtoYgpWZjlmg7QnORl1jXUfDf1iNIvXL4HRBTOSLMj9ZAVPNeRcAUtAl9cDK
zPyIRdGkQWYF4I53/Lyt8DskkKBR/xQLixUbKr1W5IDTur4xef0gH9mafd4GF2sg0QAa2k03JHo+
bv4M8800RY0HQLVzwiTNynPWzjSrBG8w2iEZ8VSsUZBTt76HIRMqP5ltUzjGvj9O/eM8wSnTOhKY
z2zGzPY/+4orS+PKebfwaN+xgT6+8SfML+4ng/dfo4EIHj3x2OE/2ajFeaLbA4SyUMzjI0IcuNqf
2sOBtskF0jI/4jp5FeblNF5Nnjnc64JVvlU8kRAdzWl+VUSLzismYDwH+RaJ5fUO2YS4eaBXC+I8
mWr2BVQpCIjfXxBFDQ+3dSbOriyaSjk5DnAZHIU0hAgHMVMHQXW63fPDm5zCww2AEGbw3W6RCCW9
SJzaOkJKtwZ8ARTT1rOHpJM00Ft8AlddEu3d/Ss6ZhIsBGogb/3fpHg6YGLigZpeWI6eqL+yjHr9
vfct0LsaIAzqWpjWPMIqwObP0z5BJp8eGAZlzUhAotBFtrcqttZfWKncNQKvG4rjpsGeC8l0bY45
HmnaxytZI1wuyNz6mOyt8TvbHyUvA9lxA3HZSTFYJ85wdMwAyQAV7d7d0Wxb6Vf1bCKxAzVxK+Hw
nKtNBxgn2HOPiE14CqcuSTuleDe9zFWnzu1Np9s+oVn1vuuyCuKTbbJJOhpBo5ZEyME9IZuB6Ef2
D0YZJyz/0bph8Wv1jFISNKD0RIunAJxMULSzR5JLo+SSJnRdkSZ/cNqT7QYvY1ufr7YyJsf1mGRG
6m051l+JO3KkzqEerE9ZmMMmXGoM4vXOHh4HSl3mEVUzA6nKqVWP+OpVXK5zGodEVn5MocTTU0cE
Dc1b4zJ2E56oW/yuwpshnRHQHRoeHLGg0KsgizJuoDutJvZJRMHOgz07zDrxDucyoQ0aeLe84Wpc
RelK1E/UkciwDGcw6qL+/hK3Wr3I7lGxy+ZILoSLEVE6Sj8cC1P0XKujysLZfJJiPpDv6ESq1DjJ
Bymrh9z1cinyIu6biWy3k8RnN1Sx7ZMlgaDqVRyikcE1lvYclgfAb0ruVmZuvc4opSYWdLCmAWMF
Ytc1iIRT3Q7SK/5CggdjO/0hFG3VVHnBC9P0/aBJv3Mvxtp8QADMHdtQjypsgyrdHz7964/oFnNk
rK9ky0c5ltkGo7EF4lCj/xg3pKxzfpNd48/1H41Bke7xmEgLezYP/mHnn6iiiRn4ZutZp98WdKuv
1PHUbITOjMTiLci6Ey3IIkaub/osA2OmkkcX3XNwpKo+fAzaPcDn6iKefXSrQMgJxhxO0PwuWnYp
kkzXePirpiMOrCHnlEt2aOZ9xWQfjAqsSiXXkAnG0jqgKbVKEPhDTdG28JFGUPpHmY5SzlH5YYVi
0X5Db6vwrNaTYY1PGK39kd5tixn5f5t6nJwdUOPBMewohlThPGWFaLfeo6OCRlmGFujBIA9mT4cH
MzmwxfJqTcqtyqW4zr5QFsdAcg/D0oTqRdl5lYr2+n+vs4ohlpzVq1XfeGNOPmzeJN5kfO+ytrfw
SgBiVoN8bu+ZC2IY0jLOmMTD3/XBWJwBN4A/U75ukEW6G96obVDX3YTmtQQZsC1haUNYEtz5tuCr
EbktRWasYCarQtIngKJvsvQaZFQl7+/icNM073G63OFURlD2id9Y0ly/BYmQmxfWuzHq3+HY7Jzi
jM94lxYQPlb8xDX6xYN8QObOj86IXySKBULoQtVFxgVH22aZnxj8CR5Z7m08Tlsjc9y/tvDDEwep
pBTzUZSG6gGaZNsXYoqjVlAb4q7y5m9vTEslj+0prGr/aVBUv1RCej7FKk5WZfdsHRkp/JhdenOU
ZGoanRQBOLj76fxdzyI1PcYPgHvCZ4iDoi0WcPFDPN5mvPzMhwIj4ZljEAwLpwvcuEL2dgDZaT7s
OsLLfI6nNGn+U5G4gE3zWI8hIHmTUTrxJEVwhOv7T8PVQ+ZslAfJvo8Qoar/Wy6SC4WpKsvtw0HS
XpN1kkgOLbPGnaBfiQbh3oPOZOKyAo064LptsgqJ5Cwk5j2WhQGueNMviKvwV8ZgWyYpYjoQ7L9s
pkoLUL2efqikQfTwhmqykSAK1qy3KRtWI2rjioFj6eedQooAgF0c1eajL3HgimBmZKIFRfcEi0Wr
CE1xp22pChTT1oYPIuWQnjS3V+p4kpTpeVJf/2edphH8vqY2Z/uSbp2fxC0l+qwIQBCVV0DEYTza
MBGHMrstW1kegeMnSl/vPIYpgR0becsU0ekvlA4DMC+kjxlbFYt5bHFa3AlVbM6W/AqkotdTmVQj
JXsVh8t8GgmTpVlASy0FTOuYgJtv8FDtzzCbHH3SsvJlkPp+STpDZUKZ8ea7X6yn+9+nCtGsQSkE
b4+Kl2hwoCB2fDTfZfS+bQ6eEL5qgi70VU3GDXhhCe7X2XHO0IIuXTfSDkqekXM2uGWinc65U77O
+gxuDgTFoaYIVhvbHNTNqBG88byVj88Kjeox2Lv3FzjPgu8hLDgbFmEyrYwjUzxbMQPgXHGA0B3t
5DImmSFPH9A0tOuwY1FUhaRKSuW844TXnWwTADphd9nAd8LhlmCdzGXgWJzpUYXaOWlRTf0NwujJ
UrmKpIxf5IgSp9ttouv6GQkTpMc/sZUG0B4bB/nZXToLfw+0zIgUlAdoyPx0IMoYAMbfq+UY1bU/
zCzncx+n5NipLNUsZr8gfqc+4KpOmOLg7QQ271JaqNE1nmqQrdCZkFOqTUd/w+Fq1e4hmiMoxz/P
LS4JfpjP/PsO74Yxm/NYsMppjPiVjxaCRH76/RJQaZ/aY66wnFlFJ37dDxK/mc9tAxxMMeZUUhco
5lxOux/aXqzmrX1wzBHkKJP/cBAE7F9yUn8xrfaQJsc+Inm0yNzoQo4WEDlxkJiWOOyV7BjHuWzx
VYZGg0YAqjaPfESq35ETJ+zOYIkyhVi5SK3OKU6RdA4k5PThkb27CETy5RVtfRSIq/GCA86OAXf+
3flBNK+ZKBHSSDNPN4zg23C9k+qgDqIhRWUeHu+ziJodGge/RsP1IkqLt6WM3xnt3KTf/hM6uEZ6
RIMy/SuPPhg1gpvFT33bjrJa0oVZBwI7ZiVUkbMSMnm+inXtLr/aoyuHvNL30lmd6/caaQelEleM
ZBvX8fiisOunTz3zjYpGXYOWslZfTqYxgj7esGBQ16p7su/u+nwkLHotsrUET9DXz91NjTdKfDQF
/L91Q/qwB6CdR1orOQmex/LiVBN7dr8Hkl1776S8XjUW7wCoAkz0HX91AK2MhJUXYQC+EV7Gq1g/
WaWLtxa2Glrzs/ZqWtt2pdurcjS0jTg1aaZzq4GdEp3Dq6mCOTNyr+usN1/AJ4+XXtSrHCSh5pQd
WGrpCdyZEnyRXifEwn/HkWwjsiKWnmCU+X1Ns70HtbrwA9RRy1vZiD8MOWPje26N2O0k7Jn2o4cT
6DoX7SU1V8b/CbQm/8NZ7Xf9qF+9w371X9CJ1M3PgojBPD4pyBqY3Qjy+sMYZneH71blCoORpLuz
b6pq4NpeEoIwIkovgk0mWkpsTZXyHKFFvSpikzVtwg9d9MueRv9l6aHabG2xmhJuROMdqKIK7sY2
O2NkjAsGI66w2tjiaHWlE3Rm/RQw68kg6j9sARamcnQG3pm0Nm6QfIh+rdxBp35akXp54nkGq8/S
ULCQDn8oaazx35+ksMARI2zSPn+F/d6Ta2bdHkFKPB1BKbrdJ/LaZhRwMZCDq/X8IxPh8gizZV92
//Q4k1OpVvIVkAVroOTbFyqEWg0PCqxvcvemQASucCv3/3XWMTw57bCRG1I5nNwOogAlQurk06X+
VRbfCsAPh8lj53U45TeXVuVCDyx+vfhPveSRu9du2yzNkhgfsDjuc0J3iQhzgpoAP0Ylxvg4BRqp
ADlHR2tLUDrzCEmZbQY6a16TQtMkgKIn+hiby04QqOamM91SNL7GQVe4SD0q3zV3hFpyuU/8sENi
OcEk/OoSegVSzUxb0jdt8uO9812sooqtUNuN8+3Jj1lKCi2xtjteT78WTXsGQQ5T4qGmzk2IAqkn
U//dV6iEvwFIIoyfclNdrNOtlzN7TBFWrW12yBdu/KCk04DfsyujUmHgyhe1daX1DtDoTRWXTnQQ
YzivD8ubE/Nb2GsaTuAqOwmA94KCarjeJWymbmhjPgryjbCLCCPmnwnW9jiC0CZHjCEnrWvFSkm8
iIu6FDJ/vHTCSZSdNT7fnEapxB16OYOP4qayrkKzgEIfcwMHu4coGMClmDO7IJMzEYjTKczNgXyo
ptXfOr+VfYSwDj5S3NfVVw50m1MwUujU0DSLr5deRdxn27SCGvRorlnddLss4UuNZvcRZ8iWIn3N
aahA2nu71KgqDEWayLSfZfWkQbEjGLHDPlYb5Xb/mctTNftvcJeOD0Aesj03IT0No3LOqsISQewD
IuE5Fvt7eIR0XCrt1rPIAXHM3wQMLVGAcPk51ZIduLc9wgpNNmH3/+F6V1jnJcgFk31jCiDGW29Q
j476+00W2V9kbtWEWum5ge0qPP1am8wmKom9P7u9QjYWGu02sJ0PtzEa83/E8i4fEzBPT7aWM8ib
3CeR9ewKv1vuzW+kzUJNxV+8fQCH7ukWZ+qZ4gWCINlKUe8DkveAz+2kOhH9wqpA2T9/R4X9ouCg
TkYwOxmxp3TGROq9aGIg6uTDkp12Yeog3zw8x9Uu6PH0tpBQ+HZ/H0yQgZ3Hs8clWg1q5feX9k4H
gCVOVj+TwXKqUSLffH3e07SVZ5VFPelRWHIk4DxycaRHjPkwl2Bfl/lGZ2HoMzILEBSSMsJ5OUmd
yTnWNcgMnxlDjfcWUfH62mrMaC2GJ/3Gxq3TQP1mhvn5E2xiNeC5gi7UuixFw1qp+IYs4v6nEhrn
DArLiSiMUoyg8F0l83GqpHaVb6JaJ1JflUPZ1mmXe8fPesoKJcTBiSiYyIAYeeET6+VVjeBNeNZj
RxnsKKHpOmMNBph91UhgtTvv2Ga4TDH3fg/nfdfSSntN0TYiWa/PoNE1Q+ZrHul5CN29GzI9wrSC
LiC6LGGFrIxqjaFTTl4onBHrnse3O/AfLwabFWQpDOZnMRX/nIiy71RD8BfUOXdku5Y6w2OCwy4F
SMBV3fr5RswwBvML4a1bupkmEltFME2rJvfgx8u8BBcxdIJn67XPvoIXt3V8mudhIQO0s2eQWpiv
T98QWdzW/BNsmu8huKKCFGS7k3U0WbS/c2E+nKdeD+AQeQ/7MNlkosDeJFNPQEZFxP7XM+n3o/39
mOgXLmZISkFS88iA35eqenYmHVVPl2bXxjDU/pSt/3TfD2lGeBlsdmww2rNSVwWEaeyfXQggnCHw
2Dp7QuhCXY+Tw2HJuNmhNf5q3hzyzIMXDtWn/i7/8xUoVG9bYP1xI5g/pRDJaRmuP/7CF/5hXtrT
lE5KuLUN/V+h/hlYD18yMndG/lq+37TcW7nGYYVsIQHN25LITHnUObaFVXZUietVOTepj1Qt1iKo
YKmVKAkD0SmwNjIcyedYmBwgVsGGJqv52NIVeV5EpmQXIz7vGWSkSLoP+SfmHrJ67epX4y66pkfE
R7DVFL9NERkMOqp8BehYAFa9bCa8QVPDSGBGaJy/Dv+PCB8w4YMoliZIXWMddjsgGWc6iy2yfJot
exiiXzjBO/76xTNN1Pjx5Qk/7bT9F5OnCCi8t0khFzQm5RDVl9ZjcH6c5X48g8NELXFzbTRfgQMb
k0am5AKRvlm+eHRNV4y8vLIDcLT6+2C27c/hjiuKYcdL2bVG04kF+kerh2xzIWpFDd4PpTLKNo0w
a6AGFERE9MR3zXHFDT0X9b08wtYB0hWyl+ACKeG/dGsthfseewCvuga7FtY1ck6bwQjpGFB1chyX
7E3y3+RbF+YU0UJpQ3fS9Esx8lomX7BQ/YVPm9yhQAuvQ6RZjgTrEfLh3kxObUufKUNIKfVijyUY
Bu0khygJpmVXjofZALhWbEMP3kRmIYZpfoGWe1DTifQrOdUxhrmsXdJU3p6OkpT5RuE0x8fIIFiC
B7T8N4GwOZMxuGiuQ05L2U15g0segZdleEnlrlqH8H4WB8tY/3iaSsImDximo6RPxqnvr0928Aeh
AF7gZfhOW++O6eeZW+KNvnQV/xn/1af3Gd1H+xf2OSmNVA/PpTgP2oADp00o2R6iiVE0ZOy19rTC
8n2xe7CRFv/w/U1yuZRDADfbmJ5uHtDNBJ8ZuXf/4uUxsUCj4umCqcuZ4iPiKg43ZVh4GhltK1ew
nB4CyPwUobYpLcfACglOplxyUQ5UvzQVLOjLn0dud2V36QRnF0QVzazxHQ1EIqv+a7U+8v4Ejo5i
bApS0AqM6FUnv0luZhDInykETFMxPLeqyh0h0ugdbzjwSb80DdtfrpPeYSY25W6ZNCTFppfKA6tO
flVnIPQhjx2UZC67B1rVDP8KYBbrLMl3DZO9HrfUrchm+P9TWQdQEvvTUzrIRwLf97Wcvocn5nzB
d3ogdXfSizVkRQ7DbcZbRBNpxF5BAEImIb4is9bZMoel7Ts7FeyEtqYIFOllry8XF2UIgNBmrdxy
Fa2bfL4cLxMVudAbt2+s0ujai+1qC9outDHeZTlNHUlmuCvqiRxpxJbjEGAyLkNaAdtQClaCJeEO
dhqmcdGfCGNa5sTW1C4jqO8fGXMvs+iO6hRKyt+BdPzWamwtAJyt4xrvoYZjJN4AS6Z+JnJShRA5
DPCMsEuJEWCqV6QSSr/vLKB0cRjwOGUcAZ4Cmzh+0T3dH84ETQVhQ3Ssy9LS/xPdaQbtpLoJJkAI
7bVTycCVZFG01Pdhi54FxI8TAVOSUFZrEbEmqEOt+DJ0KEGpIht8+YmzSb/N2ucKAHGWtTvlBUKG
xrnriFeUGFfJYNJcNdQHtbNIL6x1W9RfsrtjHKeim9cw25M8p/47nLgwdJ4b4GAWbE2XpXy1ISqn
ckXNFK911JpzDSrHt/iIKtAqlZxMrMuARBzppi7s9RMxlMbBTpE05weHBwLraai91IAJrGkA8fOT
mCO50+PYX1cy0vpWB4rqspwkMWgSyTyrzqMcGwTX2AAm7p47J/GCHOI8Mauo1wZA/iuF2fnaHpkU
hXFf5cWfJ0grD7mRnnqo2/ataNo1oLxbKS4F4w1fhQ1aCGJxJaCF5rph+WaTGPQ/BT0omirfodFH
G51Va8yfp8vx+Um4EqhXOXaUeRjfIg0HAyE47fm60/MiPbmmXoByvBKcE0co73dYpkWFBQcrJcv8
a1NoTQwB2JHQt6WmqdEh4S+vdnWfsE5tWZetQmBIROBe4M88m1e1prZihhEUSWCrfHZsDWoWA3K4
yJFjuOAxhdiGchh3nNotrz9mDMbXj+rIa/niWsaO3KBo7lGe7tee0TRJE/SRL50UAsd/U+hapcPI
ansgWF4p8XD4ckqNvo0cVPlKrxg0Tca0oQu+FvbvMW8MbwmUh6wBSnr4OEe33DQsFo2M8tSWbzfU
90u4HfLTA0KVsBFr8spsANYA3laEhSEb9rgWyChp2BwwNseflTEHhhTEOrg2Jb7ZSUAq1c7wk6EI
wq/nqZwl5GSFm3lxd8CMBAdNlKj/ds+RVDI/ZeRI81XkqpISy4ypnzQfIp19Y83Y47vM1Ge2SDhY
+mcx4gZdfHl0yZIMvW6aNBpSwkIX5Bs8aMeIjLg6LiKbqS/ObgCxZlcAPoueWHYnfFUVZLRrxtNv
hDSastY7uYxUyQPxcgEI9f47e23MQge7Cz/Q31BKBGxSAaI5U0lUKQMb0nMKh0+TtlO6In1O1Bvq
hnf4SyWzDHA/Mw6Jf47veuMrQshxRcpKIwTXw2+a040CSQN6kl9CO9Yq92vW9wm9IhLndXtk3ece
SEO/rmNU3jxypC9PXgFO+cC019vub/dD8gxh0SGCzNrTQrlO+O7qGSDjE9ZaSY5JzMX4gd5yWCOB
yRGUIaD6NnkQdF1BOep1ZNlLgK1jVzxwBrmDc9y0+LELbCyjHPd9gjiqMQ1c77Dh/BXSqUCJ1U3Y
V6pmGkfJTB2wOIv3gG45AsAdm7ElHKoeQkSUX9W8gITyZkja6TcegdyxLR37rfjU7XyWBb0MkRLZ
MN0n/++2UuEOf+FwSgEb3Txrh5otEEnNsWsownAEEVNOAeRaQa21JPmPPvnTmVi6eO17+aMJEMEX
vvIX+3Sl0OMb9cPVsi8Xp/7YSbSzto2iDTF3s3YFKvOi1ENR3LAtBdWR0H59T5B38fEoK85TGyda
t+T+8a88FecHLhhWEmx1+Pi04o+OmmBe93qEYg0yOLEcLOSpcr0+LYI75HNUc384StgQKMri7kIs
BwOhIVlpb+6j/vBwLjdF8CzRH0mteImS2nHzdvNlqBwUhNlVyyqJLh9BiRXsH0xWZ2+dakICQuKl
D15XMDdRmFzb5ZWGWpKb5LKw4eSIPq/up3qN9ePw+oMkrFx3oP18nKj/Abl9yXTDvfjrPxwfffy1
hBlDcQfK2PlhB4BbIEDR8VuC/us9/vlSTeCL2yQKcQhYHxdzZda2cD8DcsTBMRk7a7NW/iMMdFEv
0ciWStQt1h0oHv6ekJ2wJncZ9N36qMthe/k+OyoSH92eQDeZ50NmXZi0EkNKek2NdBxWIGkC+j3b
mWXRbgurjhW9dYtrWMeeRI5OBcYeYWuD+xQGKeasYTj61+lcT2JAsQeyva7K8peRTCYFYrq6aA5v
/F32X1/wHryY5bYBPwabElywoNnA80eJK3Aje7kPQaBmMLLL7xsxFmXoeSYPJos61mneMTx+Io9l
LpAbzU4y4P7AF7Ktimi1FMJCvg5E7884c+KLzka7lNap4vLCXpQF4kg3Cu/20lwNf9y4lkvt8xuf
V1kdpOyEmpJRTDjxWPwmxX+kUcdJMGnM6KA4+E7/NLMphLdichX8YAo1XjB8e1Zuzy7x31s3VWaj
FSyrhPvbMrb1cRvydAvO0lg4UfSTqLR1n8G5EJpTvwGwq9MZqR+2yeldF8OTBZ3awRaPQI+IIwvM
d0+UTPQGrpqwA01LUwfACH6Tmn0u3mprH6QziXSIbBYp7zxws+GVf+zHfZKSoDHurWDnkw4INE1s
ZGRjC9gRaWK22io97ETlUisvdfDUx9YY34dBVa7PMOw9+LDbbaOj239ROR557ikKf+oi5NiZRZXg
O8SIvYebQCrJT+1HBboBA8IWR5WR5YG+BpAFhqEQeVrxzQfpI3OHa2f7fSmlhzbl/221rfA9eIEI
Cb8JhjtDCWaWAE5LtblLu08x2zvbgZwtNHfdURA8vEJMzCvph+BrAaEv54ANwDpsrkjb588qOKcl
T+yL4a8Bxa/8mI1C0jzE9taZqVRA2wsnra4D9RAZt7Jmk1pQpXEyxj++IQfKf/Qr0zGcrjc+hhnl
i2NJD6myULEncLFTPhi/v1FgGejqVEFt1yn55ogwLYdfIic9nqiUvrPBfQq4SqO1/MPaW+R/AvYl
5qJHH1ZYj2ByWsju6xSoQeZLYDFYwJMLDiIGaFcZN1F9s/i1z+6OomdI5P/2yxQvGiPnS+iMlL67
45rbiUnsgURN5Nd5sPGvmC3j18CCcQ63teBXFSErzAh9j7Vdk6VMwtZCapCRoGbITBP/16TwY80i
dYXbqepx++4RUbY8sl+Ofqt9C8wjs3H4toFdfwoq/UkUn0tvpEqpXa00FBdi7bYdbN45fd8Dh5k9
4XGW+66XuB4ZmsGqq3r4mwocMDqqYGDS5uC2YLxk8dkBgAF/RVME2lThshCklJ4aGCEKW76KwONd
GftVpDp7gywhbqT71Ns+sb6hQH3Ds23WbiT+EF+h9S7zXSw/nDwDQpXo2ekh7UWudujZXbXviFBR
6WvVkkjP+QzG89aqDPc4lXg5ItqHh2OEaEg9kGfvyKFtzB6gL3dbnGSeQxpEQK2rQ/iNCGxJOIwB
zVA/oMKzGsPVH7vrDhX57lspbjUWJL24cnks9MU6P/gs3Ixc0J+hCV2/IS2urBiVRwgmTCdqnlhm
x1ebiiqt+E27wfEfH/5GAKXxssnGzuhAVaZXepbd4RmBVruiZMQmfSlBWiJmAJjwYhTlXqETTn+M
1bbTqWVStMGZ1FLqMv9+zhrCQWtspr4GFH0Se+kBMDISGfWoxeRiF736ZdlnaUvtaS6rTT1edb2f
DDVJJGbUJ0yknmF2+K5J4UC3atE50n2CanG8nInzC7Dy6CLy6g/qEIdceX4P6f2b3h8LZdiNphCm
h6M4NZPz+zNpUAx9sFIZr/oCsIb8XxUDyq3qntdoXW88YdK7pwiYmKhREJxQG3LIie1j6AVMW7lY
wr8BH2H2YJxjYyJjIkL48sBlpcBCTEl/T1eRM5OKsBncuBgiQL6GIwwGelEwmbhRKWNV1SKg1pQW
GXe2NAtPeiEJ6TEhX8hMblLyGnghE63iTou9os9xB96sf2Ledjdr9MR9h8048GijD1lJIeFrLnB4
FpBEm58xkjiOayr3SCPyJzqnpRHEpqKch5JXLEP0MbECUu4sDINR5SSCoqFBmS9RazMRJN87c+DD
E0j9lBOWsb5dni/5QsXuUvbWX0B9JumWGJMIRj8Lt/uHHdwG43WI2czI8sbFjqkENm+kiiH/XzjW
AqHjOOO5Ym4jo+Iv+QA1CR8EvMRealRSAbnyiKPSHKSAQxcENJsBsFBykCtC4evDP/kIZ66zuXzL
ddNdZ6pZdHUJmo9aa0i5XSjTVF0KWNZXEz/FT+FweAloAZfJKH9O4XECJSNscPbtWqElg/Hc3nmI
qIPK7RGd2OCK+W/VdZtg1ynyN2Sgu1umI5Vw7std8gGBt0TGbFL4tt6326GJf0oCeyPHh8Dtz/9K
fqC6Sw3dBFwtUlIcfp8Agwy7+LS8jFyrWypLKg0CMF/7CLv3+yorVu9Rrrlzw8MPC5kGXs4DtWgk
LZGM3ZtPihkCX6HxKnMaYFLUCXyWKDr9OiORnMPYyGrBDHtgCgwIxX7pxqyhZHDKzKuibB80gn6+
9wE6KqFks2HF+bkv9xMGNVa2ptUgvL65zOrKCzR4MK4IWxY0hr0f1j1u/IeynWYYuhFNMFZOjnTO
WZRNs2U0Xy6ld6/WQxn0+XTFzF/4Ki4PTMDrj5X6zPKVZ+m+j+97vRCiB4dltwVwPZgP1W1VDTQ+
Ok0NtoAxbeVP9vY5qxIRF2lCnyQEDdtPTtKjpgVgkMUHYWfeEHBh9gHGhXhNZ7fhbJ5i7hsdgZv2
qejVhVmiVEqtoaejcvndON0hKVH6AqVjUYsaLnw6ypWMIfnHFeAv2x/Q42K/IpZM7QpZUFxF9wOc
wrHYsUsR2cam6u2q6SdnQnA5Ln18KWW+8tJ/5YtBEH2o/9umRHytW/zf5aZkXCZVyTdk06z2Hbfu
v0cBkGmsmBjCUPzlX/CTLdZ1YpqZgv1/1s12gEOyYfRf/chzPPBZuwwuuIJbgdRAATQ/5lLEq8wf
0kDO/jDJDlljNibg9LuYpFUbzGvCh2IIGsCAaac8REHtzNRo5HAiA+LhLRLjoMYWzKOlCKrgQwJU
+06RLBJYCSfQ+40k4Q0cH1xLKeh18E/xZvI5xRkr5ncIDA1np204k+2P6Ru9DkSQPVbvXdXXTll9
Y5eriRT0e+TmiUX9xNbQwqBNQRLfYgUWD5ecdByil7Z77qqenJ7oxzp3wOtcCMcN6Bl4/TsuHqLj
INkrTOPkm/jdkZjvzvUlzM6TnN8Ze5HeDsAlOedI4/YgTMKMQAtDxkMiN1kiUyoUfH1+Z5vDx3vg
/RxYCQYZFMYJK+PBDmewIf7KE9ftULXp5Y4XABBP+pSW7fE8D5qp2Z5QrAWCDYpgl1IeRp19YSs4
Kh9yobj2XCgWr7+Mt3uqVZgS66aLrGUy9t3aJ/drkKSIPOMlUbunGqcRCypRW5VPsPjHvshvG9wI
6CBz9KlbQ0cOjOaJr/Pd0HLykqSjgA6waHXlFx7FL8qJcTkTgX8xfhfWh0C7FWqdK4mBrgS4nobR
c8nuvdsDWJ3Qov1Xu2N/K55VDwaEvEOzVdenEHhUM3OhULz7iz6MhupQpApB9hBCQlbVFlzYGmIM
C4/7K+0SUqJY2tNTl3SP+bdX++rIVe6X7Fl2j0ZnKicF0Nh6oltTR6v/aWrseRn6gRWPStjDZc/D
wnN0LxyTU5tnVWt4sDE+mky4DYPb+5N2+tkhzIqh4UqyTvlI8eNV6F8y8GCKAoYGG5jT2Av/7sQ4
gAXc/J2Axf9I6qLOBVliSZU6zwI51OHFjZrSP0K8FcGWGygqrv7PwCb65Fbc2AWUyNoYkIuUOx8D
SMolzPkEaLJMdUExfDD2+ttVPvgpKl8zl8+LhSX1SQaboEQj5/s/+fKPgq6G/8wjbbKioLRnOw7B
oud1m9rFMhAzINOEq3yFp5NHQhFSAQ+MovDL2fuu/4x1is9OT+mJrpBwsmehFYTaNNciU19evK1W
k30I30UdZVemMaukJjs1xNeINURgu/JkrIhO8N8Pc1Z+VZ+cLRRmYIw3Fs2BbccrMLYG0ko+EKty
A4o+Aw8rP91D20EIfGrhhk/LjSqHP/QaV+40p5dB+cd9m9nzI4O9lhdbwh1UVCNfyvqoqcl5YhTw
0a/tKRadu5cbklmTkZlLropTLHRTsjQjrTLHzGBJfcWE95txmuUw/bDc5xz2nIQ5WzNIuXXQHH10
KklSTmlYMkUnCMNcM/EJd0CwU+kWtzODkVO9ksQ/v/El+bf1xE8nEVuIhDyuq+cpd+u0ztNSGwTP
smu0ddsE4kPRuv/tghCe8dvfhluFJoI+L7Sdk+I1Ah3N2j+iHCmADzzTHXeX9sjwtL2uy4Hp/vDp
hYfbtLgysv20IBUBIqR8v/TXeM59ZqDqhhD2m3twSfweTmt824xouLpMaZO3jWpEUrQ0TCRHW3UD
ZrZvjTP/bEXji2fcV6bhZd0pdkEBzF0ELMTqv49KQvzLzEQ6I0cjAdEXTg4uiPWRbSshjrPDEwyU
MaYvt/QAOPZZjQFlUEpcfqvDzDilXHtSl0jSTgVkxHIupywBX0LPpxtchR867iJ/huUvaoZ0pM29
IjIdy1iwSWaEtRkkdJEs+Ns0n0pIrUk74RT5KI/KSadB//FSnUA14fELfLORdUizPscOcEHItcp4
GUYRH1fK/24yqIcfTbvCHUDwMJV/rF3hgfcQFxYTOg/btVl9OXzdaz5W7+v79Xz9TkpfvWTHNFNp
u4FPVCRnyL6hxnQf56BUsGWAwfhS4daeE5N1j60tECSNGweSG0VnWUhEU+YnZVzcplf4uETw0Q6/
7xKyDPkdx9m0S7omuynFyi1ipY0fLImyd5YIhzNezCRRywJFp/2Vfu/GEkJ7RSZrXAXvQlBeZXqg
6ZPgAmIOgn+p6LdOZz7lES6eF8KiGXz469Q3XJaBlS+CzoQCQk5vPaFS5FOcqpZ3iKIHCzi/A2to
2TW5B82pM5sOxewzUl4Q6PKIQDvLF3u5gpS7Dx2hyI3JvBLdAp6TR4vE8txL5tn9pzu+sWqXOGmY
VLD+cKHSgFt9UuG267D+UEEWul+7Smjf6BOPwp3YCNEt7UmM9xUYNX/RKcppPyi1KgRI+IYgRuKi
6PnJWG8+5GV36PxNDdgDismiScaPC7jNQkiiiPEW57AmZgV6fP3EVGmUJasVaRQma10rvYn59yPB
UwoCWQnXEZEqQ1QPgk0yXKzm4qswloMV4KEOavC5g+jIis0UVnIA8R0NpzQ+QKfV8Tx0RUDUGPu5
3hO0xWnfevmfIY++gH+S+mxoQFUWaKY5DDsv8YuvJxfKHRN4WZ0KgNSErjFDQPVjYqe0OVSonNPq
L4mRXT8VATvocXSazjaw62W2Yc7zcCry5tFiFsNyjnPl4z/DkhULAHcqT5cwI9rmRCJM9gcXiYX1
57mkDp2rwTBqNnB5MGnza7eYwkOJaQqmY1jRJEAaI8fUYzC20Qw6kllngHkgMsXeFSuEVFQzAPeV
3GnXGIElVQ0EE9AkR0Y8yHo2nxu0Do5UlzMdxNipPw72h4Cc3V324VFlDbDKcGk92FWIlezq6bYL
1lsJHROBJT06zxpJ4CMUysc7RIDhCR2ofiwkgf9o7W1jL2E9PTdoCh04wrT2NRMnUMtnmssGsAHu
/0FC78evp44CiAGTZo3AVwHGOBIsjOT9z2W4dDip0Vu+/ZdhcuPNDVkHS+7XO1d4OTAbB8CnHAC6
5MKLsdpDWHBRni+BV1r+i/y3cTrZbN/xBZQ1fi9Vn7wZbSVWarSzBXzmSlVlTp7Dln98ZtCNFwPO
cjAiFLm1YKunXuWszJHkeaujJbV4lLIuKWS8IMcm4UB9X9GAcmb2jMKXYYyALim2duhYOQd1gZr0
PzwiID8EGwqGwW0zjxXoPoAXJ45B9EKi2MF7lTgRA2kh6tL8IBjYMN7wt3FxPsAQd3yVgurLvN/Q
5XF8KeM9UxkgqPbmCecGzgl4F8/J1cJ+1YyRiToeQYio4NZxCq3tYBqjsxyXDO1PbXDPFLiZ7PQq
dt1MxF2OoW4AGqsNo/uHfpNslX0bXM7RNg2DnG9B+Y14VMwgy40Aw3doRmdKah4DLMu03aRv8v9Y
U/qk7zZxaHghlLjtUKHZZ9hbYxrlSN4A/1XnoyGyujo5arM99f+V7QGRTW8fR0fJt0fapw/4jPw7
0EMvZhaq9ynvTzfWXdsu5of7bxBY4UkIvv8lDtfzi5ZlNgaZPLZ0t612xVqMD9TH7dPGqKxZkZRV
OFsXSFnN3p8ejsQJBpj6ZnNxomuOHqlFnuOkbd2j+yDGGzrkazH6NMl8eZXkZM0s4kI93ek/C99S
X1Q+zKAqgwIDjLdtRzjhF1kxhclPpQlT9ZlqJduQpVkL6kqGZM5iNd1bVGdNnjGcAR5LY/BLzHcs
B3xd3+ldIx2k75H/AFC5Rw25+igYgCftrtd930/iw0UKsnYBXjck9UcGLklMTuqw4sMOT5R36o1V
C9A6W4ya+PuOTzhfWAlw30sQI0vfZEB2nQYA5L4UcgGZL3ATBju2PCYEC/8mVySZc1o/DRjT46Pr
3ONn7gbxwZbsJAMfhlImpe4kLNo+qtbleLGuN+VtiMwjHed8dJaC+ph1wA1xHDPRv0kE3EA5SV7m
mTOXxgLrBwsycLArD9OASE8CbrhFOtDzlOGZqhXijo7jIH0v0q0oRWL6GtrNCv4U7k53k/dp/CnO
mcCVLZIJgBDpZM18eIN2PEy+u1UMQlCmGz2kSv9+CPgbDmW7YHBe0mgggvs/bDgVMQ9Yua/3FGct
WHo6P270fyKnKmtlNcBAuqoJ47uikYoLliTMSDWOBYB3Z+edzNLlAwul6iH8gBksWUah+9bJ0eHp
Fd2OwiXVaA+fCz2mYEgvbI6AQl9yay7hZJ4bQjADJ3OZXBdq51cKOQz/cs5ZpqmsDneKUzatcDvi
F47+qfruEFluHhqzhDjdR71EqGNCDHv1+0N3gIRKlFlfsEdKFKf+6WTmnaTj2TAKtNI1R8qh3WS7
YCifng1PYHHOCKklsSGWHc35585xMXP0nzCW46+bCGuDxECke2EezSnsQR4FwPNkG6lJo0IStnFb
KBVsknuoSNozP0wyZE0UvtZwLeduHI+aoSsGIOwRNEdCVzCFFO+dxB9l705QftBK6OsuCVSgwvz0
qnaIrOObpRw6A2W3/eRVwD3jzoXW8cclDtT3OTnwdtpYaqMGBOW3JCLcb7c+cYJJdnuB3NyQ5oRK
ZzM4mESL7PRH6egnznijK/qsMV9AsSCteHqZnxWSvzu0GJdmeHyq7yQeL17u85fsyi4/hXeUqBqL
+mw4eBjhVAvAFjWY9HRIObjgoX8LaTO1bIpfOecFYh255CQ5PCPLz91I6lbo1g8wCVBrXSUev/6Z
6V1eAw1pQbrA+WPZPc5dpwFOPM+bOPUrBKh68X2zDDJI5GAFkHw9qFIC0LVF/cawAgazyqhX7X7u
UStiKPwf3BxDWfeSRg7Chgc8ajTMQVBrSGdWjZzELpFGcajqbMCyyjZgbko7w5iGB0kwAmFkW9VP
6zHdwu5s3EghmSFpV3wezIHTjeIkBuDznDoyE3LaqCPspcK1c65AHJpJu9KAsSkBJZHn0Cwtlmq8
0evi6mBfc6z2fTO14DRysp4ZG5SOW2Y0prr/XQAPI13Z51klJ6AmZ3b4yjYBMQ10GgpR0Mh69qkj
FAHRAnfEctO7b4Lah+SwDxf+WanUeDiEItzVorrk5X/rWt/P11IrbfZkwtVaFyyI7GOVnletqnuS
ANmwySt/FLQbNnPSE0U+1CXvZD/Cd7ryj0m2y9D31pBj47DB9h0PdAKwcr53xv975eUoNr0PSfPX
GmqTI9Tc3LA+93Y0R5y8Hst5NrumYvtHXAe/LIjVXCQZKpKiDY155X1VmEorN6I3SRmtlMrmThJX
6/xVqJaJ/EAdgtdVMEzg9m0c5G88B1+4j0yGmEu0g0H7dz+69+vbaLnrr4RZT+lsnDTYQAogsQ5l
4UUkpM8Zton2kuc5X26G6EqWr637/WM/ggqnF0lFiLFSaDNeFiYHLRDdnnUasOp3fwYPURYsxM+J
1OPdBjLEdmXIgbvCGqNPFsX3BL5FFBiBI86PXe490ZfSqYlhS6rKXA+KE8hQTv920XADszTEeRWD
Kw7lFouBA5goSVffz3H2ODICPWToY8vmLHgbakvMe+TRdPzTKNUwsgP0j82miBMZRxQecnjHTWYn
/XMnU7kT9+SI0rv32Z8DjcsAhirc6URU7y7LyxIj1JZK7vc25DNwY2M/G95q2BGqHtPpneLdzsZh
rGAeAAnL9nZ2EOmEAuRs4gTLTtBGsd2v7dQ8XkXwDzvg58mq4M1q9FEfk4SGcDujhfzMB4ovJCEJ
xSyarWHf6DwHKrOydJdYQzTy1nKJ3mRtf4/XkAI4kMxfLXtsyZYdtr71TgdaNt/9jeiLQOBpnlmp
yDbuIOpgeTd0cj7pUeBFJDHy+ZqnIFaiOzHRg6cUKyhuHXBLlIscikM1WmFYoGnJoPmLgbjuPHNK
3hve+ctjrWazvdnnEdAhjTy1hWQvn2bV4b+eWGhuWPu9me5j7/bLlOPe847lY/zSyabuLjVo6of2
5gJfbk9L8R2pa/3GB12NzOV7bXrYMU84OtvMjjQ44IDTMzS3J3xNxfYc56P0jAJCu4PWwSwEToP5
y4LV68GiKZmkCZdGVtWJ6D8qQ2BXFwpY2KmBBXPCDIdnxMD/oJpKtALF8HG8GiQakGuub0Shyw99
lEzpEyE/5JbHocW9g8V2EnInP+kGPM0Ny/elJ7fKzEgfHlsXvBI/V0ghQMG7pVEqVeQ60pX9R1/7
L3uzA3fsRMjw/18+sI9FtktI8000W4FZ1HVUZjZvcXsNk6B1ePxCavlx9otvW+GnwzCPRqqrL/WH
k7Ozme2AtW+Z7CUnpZXugRZUkGvzIZ2EFNcaLod+UThKrin0bW5UsrzU4WLT94p7ePhBBStsmfU5
epAfpzFUOu29xApMG9F2IBdstlPsbUvOyKiqMbrc9EwndM/9SiYRpmPz6IESk40MS/v0FoR4VkT0
JusdXVugj/xakmYeke7LvZELICQPPVmLf9S4XMCRGxx4avdkUCDvnK5xy8xcerDanl6bhswVtehN
eL2tZCOw9zJ1dezofulIs1KcssH3xu2utuwr5OicF10wheKY5ac/wUqteWkZVTg+NDBHukRYza9J
dLSMfzzC0p0vlvBnFzlzKtnpopeKwaTPxEZFBJfIqBF9h33ayOPm60kncXX9p3H+8aHeaZd04IWq
PpBulYrv2ozG8ZtNKQgrP8tuFxjn+8iTA97FKmgE8eCmIbF9bQVB7sN02ok/+JFGJ2wa3tMmDggN
QyGsexk3c5oQE+i2C9wjIf/8ZYHxm1W5xqyCnx1Evv5XnBcet0c3f4w+eqGnoBh2an+Ocw5r7/SV
EiAWQtE7KC+A9DaHMUgccr93xsJ8yWFgmD+XR6IzgDAuMje6IJJXWzn15d11FfgDkpGt8ZxRyfID
rB95ulBTin+glbVU6EHLuDXMbmS5A55JCxJ38DmEv2RF6NpR+PeHB1a4IYjtngSw2uAXonzvjkMU
fNDNP44WfijhchQZG42v0Ez7flAncw4qa8gyw7Wl1JJFq9/j8i5PBApjh2+f3XP+vqQCOLbLaItu
dp56A+zXJq3xzNmIXECeOEujRZT0XWbJMThi4d7fRRPcpVY4oIViqMZJ527ms01qMKwi8uFyYwsO
jbLwmwFnUEnGlevvlpWR+SuTCkHexD6ASw1MFHjIVCoy/A3i3QA4jzKiDf4tgn4jaFjv5jAV9AyC
4JR05hi13jE5vD6aGK+ZIkSb/1u8Yni8zzQFEWb1lOfYW+M5KoNe/mRQ4sgBQuyrYlOOdzBdfPvh
7NQDiKbrDQuI7bM4ENmg/+UI3COyTTclSUv44EKdRpF6HreyjFqzaGwpAc823hqAqHFTCj5AEQOa
jBtzwlaAr28T3c8d58YNdxWCsgLUWbWORXeDIHtt8CVb27zjDHxkcci9ZSRtkUMfU3dyqK3VwXmm
8mz56o5MSzmptBG8tXRfPgc6oTWQOS0rIt4VJwvN9dvs+NNgfmdW+1OneWdoqZ/yChkJRqLzLRfQ
8sUfoxlloScvzAglccwR0Qxa1fSnnzDvdQtInor/E3z1p+0X0D/lt+ecWzepgz57L0OFDmsX171s
y+CN7uxYkm0vg+794Z7x+Sk85HJD26wPq6UEk6CBiM5X4VbXi6WXgqj0y6I+5QATH+NLpjym1Wgj
GpQBc/gtPzxcheObKTY42VQy3Qn+Cqnm+Vol8FC5aRjLniO+Sg21qOUHsenIexpZEO9d+bGqk/7q
bEzmpSXtdiEL4c5CNKeQJuira1z85EdW9jCpDBJXrA4UGvDpVsKcAsfm+wBVG/d+e/tP8RBv32RC
82EPVrHigqkilkIj1klASujv9dSCNDWVZzWVCIFo0Xo/4zabdGTzY6OLNw8JFrVFFMJ71d0z39kA
RqNqSmXl9Jt0Uaaiu8A2ii4d0W3s++9GG0V/6kM+rLsjiou/SvEF0rYDc0PvvzqK2HqRHcJzoj4s
84Icvrtq86jf5xF1d6c/0oZBLjD0ihgxp1v3DsfzIZTFciJb+M75BSJo27IjdPe4ZiU6zs6Fokz1
iqMhnG4Kv37xoNEwiqPiz9WRdM4zgs3Cf6sMTuiD+QxsNn7QBvuQhHjkALmt0zTTHAbhX0HO0SIC
Q8XZ4rv9wqONj0CnzQwNh/jFcuyoTzAYEpbPP8h33pOfxmaIwIYtgAQfN429SJGoj04j9Y0cv9q7
24uLUj2u0FGkWM/3s0QjbSrOhDsLxWGSGVCaOAaPK1AcBdAKf8DczSNmnOCJgT7Y7deQZqlwOGPM
yUUeH/k2H/zTfu0ZG1pscxE0RYmQn877NfP1FYU9xdOMOz5czY/7ToN8+O6aU+VndvhISLfETfuR
Nuite18m+8E5m6sJiCO55gvzS9ZZCXESyjvmAhppUoAQElarDo/pLEa46mS2zM2CjjH5fD0q9BrT
dYdyZjOorPzBme2AvbwjZFYa8gj55NcArw/0qC4ktetpNTtWj2Er5u0nY82p4bwlNSX/HOERn4or
/OrwH+qiZbCIHKyPBgT6qMjujN5fRXQ5d783Ty+miQZAxdSrryXgLn6wOX3Vr57i8yqv+FdCyr+7
ua/GbMes5uVrA4FCT7AuQLpZPRlKT6ioY47boVL+mhKRZhR62sOnYc6Bkrh9K/iODxzt4qAQMBmK
Rproynk4XsM+44B4oRUSSX3bQO67fDzBE+pUQdKcdVOa+PqTA5OWwGz8FxhBoOpi9aFZhRgTHBaD
RDFFDffIOkpE7y8xdvZ04bo05Wmk0KwMB96ZBzZHuknhDoqwTjV1UK+vVrIBLUOuKFNuP0zND8ph
vhPv06NJptf0Nw2etcrUviLMc+8hSEFcJwMWl9oMROBpJKfsaFkaa5iTaW5YgdK5eUgqeCULRrkA
DwnvSRhMiWFbkfdM6ffEna6IOV0DDVwMC56y//nwGqDfvU7aVZ4/1TL2qkqjpYEvFvyORK+DlNpl
5cZ2lanlYIQGwG/DhqF5iniPHnlgy2j+MLYr3Ky5cwDb4AntaqtfrIPxMe9PRXeaHq6VA8fhNA85
eNN/aXwEliuSpYQMLIpekh+mJ8QBCujYmzS7Q+oz/A6Pvk4/NEWd6ei4StwrfJCS5kASErijzphN
B4jzgzMM2pENykWw+1CXj4P0dELbM1FE4FLe8XD8bgV5ZZSuM2xaie2OvzaALpeirw+d5blUtCe8
riz46Cu7hqawiBCz2WyMv4JbEmcVfcAQlEXsCPlyek3zvxWdkMl0cz68S9ieC2CypN0Znq8i3GPa
B4p/GHSxMzIRSpbWWLkdqRUYRZ6sYXqpTY+XlkjOhpDTi0vKZUZ8FyGRQcOsSXccqjrTgO4SHTSN
5VVnZPl7bMfSjjnNGwEuCgCAnUKlwAhkAaQWBipJ7YSzraWjbAMH4GJSuSiLMuNznnOoSZ/xOlJx
lHunnE6Cv3IYJjZD4FwNxRAn4O2074weSjK9FQX4B49V7dLR+OypVIzRKfLJUmLJEEQzk/AttbbK
1Wl2g5UzekoP7sZGZm69yPfgi0mmn2pgJDjWx3s+tbx5ABhv0iiM8hAsKULtDpkUaA0y0NVguSUo
2L7Ysr1jDociZMzdNqZzbMeWaCANDpYy3oVZ5X17HvENzMhY35Vekou/rowlAypcFg4hiH+/pH5l
Y8a+/i5jwDHmgUGZVqJ38C1HfH5RSpu6mcfuJUmFV7vOLPP8oHeY72iIV5/IGY7zCntXKExzthzF
aJxf2YHNF3si27+QD7gqWjMMMAG1UtwA7jri5AKhXxIyHoLi/kFJo+/d1iL5n5n6Oz6Zobp6pDL0
sVEf4o6C9HFW8yYx68IPxds6O7q8qdu/vRQUWcEuYs70OEEk7krgckdqLA5PAqmzTlLArCVsUtAg
Q2j08lXapZOJWPkJ304CtAlHSNJwg/ti4YMvJHBern7cDI5QT3XkCwIvBGCOaqXBjB/9QPtFLz7d
5ZC/GKVMe1vp4u8W6uzKbklLYDgpS7UpLCnPlzqQp1gVG43qBD3Ksa7xCIHTECM3yEur9bWGDDnN
Y/KRss3csuDH6ldpNalNF1UuyeOvvwW0kugIiTT+5RncpPPP2UKMWyK5F/aQTwRV2I42TNPn0hlQ
1WPqFavd87fWHu7L/naT11f9JaGmvPSoaGRAVsQx4PdZuBqceqsGNM1c/tHFtr48v8YvU+17Ab9k
XnVIFGqwm8QlmS0g8jqnkrkOtI43EI+01rb3RjUYBG3JmI4l8vD2tOOfqXAdtiEqH+bdEbklYpDi
8ZVLp6toApMRy4D1oVpH6GbgACeVP7cyzs/83pjVs03Z3546NjAeygCe/r6ljKZnL5Y8CKYkfjFl
cWbAl/7eJ0FjRFzCYUZDccEBskcnTdVOm2MrhElsIu4/6vxqFw3Vjt/Kn0vFPGwhjdEYCaopZ1/+
bMp8DWZDLCsasE6d9T/JHZdbprPG7gDcmhzfXqgwjNyLx0apwwPaBh9tyFp0/hOoTgEbhHvXu3ht
GeaWySpBnG3NZuURcA6nVfyC8EVF+Y/byLpV6IzfCjKzeGgRL07v0ZkXAPBZIjr/S0Ea605k/jJa
ct9++3aVe4gJkz1dU5BMTr7kH9tJ5VOlnzR0Tfty3ON9n5/nvk26mqg1AEwrg6W7do7vHseBA4PS
O+e5QZtPPXGVUb5lyBQ+nOx1QyWryvgcT8VbB9HcVrLxGI9EpXnb66u136IPceSHbZBZyfvPPkIk
LZzHMHnNlR85xLLRI9Op68E9TWcThjrinr2nqF3JQ7DFsnXtw4OjObY5NS5B+CAcaI35EUCMZT2L
xn+TNtCI6qCpHLblD9msS9s7hr5FTAm83+oRudqi0shUjGmqsOLg/96SvGDE0nEsZprHo5LmD8W2
TwwOfDqKMlLWG4DKx7sOZDhpXlCIqyyKuL2n4R26O2HLma7WXv9DVpfb2ZcGS0is68WqvDohWu2V
9g0l/5FYSrEaBNwOjbuXn/QVjdjn5kqs1yclLWZdpIYMJOoP7BKLVTyzQtvKHjYxjbKupiPlGzUC
1Gy8UT1Bva3xNkCNxFPanCmWZVV0L/xnVtYLX5My/Ly2KJJjTTc8ZBVLBcheL2Z+soS40C2FK97z
Rt9/zEp072y6ZNJddVM3goHzdmzYX9mJh/xidaYKKyrDDJDeC+TWcs5/eggJmR623+PZBt3dPx8g
Pf20qmkf6acY64dwgVwzjwl/zK+LfZZ4EhOJMTVbTVz8H959ouJD1JoHpkO2fnB8YDGqaolmCyLO
HN2HGaAIrEcB4z2Lf2YqrjxTiVjMWwhvd6igc4x8QHOuJlJst8tSy13eVZSeV7FK2xnVPQtnZh2K
TTJ3BrGlaBkQZ5XsrwB+JwwS6+ymEgliH8/ZWM3foauR8zR5Iq/AwUtIX7JqLHLANMB0IhRP56fk
+bagzcUiphdlAgALm3fd0b642cen29waG4v3hAoaM8MxcZQPVp+YeXMbyr5d06MbSfmPCmTpEnFU
KlPny+uMlcQ7HQ8x9kZlrYdzHtg5Ery5cjfB4pinVRHSUCPcxkSaZ0e64HPKUuvzeBEsFVNSDR92
jIUtEyzmsZVX1HqQ/X3t+iwq4IGsfXNSI8gvs04xIS+L9xeCORN89e6xYZG8wmVdO4ph9y0yBTdH
a5Q8x/Z4Wf0BgOTuACCYP8uxKgFIcGqX6fWYFQeNR/x1O5nJskJeKPB72+j9XNVPG3Ll/ZoHMmj6
v3th9HFGvUUJykp+mBg5e2eBOC0+Oh7U+megrqSuHK7DcJYjWqW1Fzqpb5f41nyUJhimVVKCewTC
pqDZ648ZUlpDx9D2MTOPqxoFeuALQjdgVKWx4ilMGq4EFAUJLX2Nw7eoHZe0QKjwNEkERMi6RXq8
omBbdWpru3UmbIfALZ9RYQPwDzcyjQbpwd5jm6vZNck0uk2cE6egCK615AQK8qzuVbXiGfZ577sg
IkjYYW5KMB5oJLq4mK8HdbyNOjS8q+bXn+nELr49s5wG+1fY+u0/ceHKiNoOSfmnvS4PWLk8PVlG
ghitdQsvvxuORCjBC1+wK5x9xlORKiUJPdIfgllDBFCSOghrqr1A4neaFwUrxiXfPV7nIGUfZuzo
D/hED3e71xS0/sKvlzMXd7s0tZg5dT6r81CxM0xfq+rT9OuOdi63sS0bgP++QVpqDAXo2MygCPnO
UxPbMSH22pNV8nCJp6uiHkZR8OKneKqPipQLpQ3OChrxm+70ruvtukB7SqoOlcwEMYrBNXf7EQ64
yhHLxTG+P6D8XSrABqCh6OetAgL2OvLxH31FLMk6x4e9+2vW6UNLb4SuuZywqhOe76lGicf99Qmz
6vKWKHWZtR83XxVnZW28zmFHgdAF5SHUaL61Rp5j75TcNb85BQZUDLz+a+FrOGpgvoy2IYc2pTnE
gGX1HbnRv8x+J7UD2UV8AmLLAMuHoXpNN7AAH5XCHBIFDMXwL7zTdBronCkQ9ZXOZ3zhsUfJEDgQ
xrBRZzoOkcvXzjTJuJgJd5N/960WvvUAMrNfVs8s87zXjvZwc4h2jeBkfW0yj6ly2xjd54kyXtmf
DKu3faZqO4pLuFIyjo7rhaPMW4mvaaXXfIQtq7vP8aNe+AlizJzRYzBf8ZzyajHrwFZw+iE5FIQx
IXDYAh1gTa0zG2Gg2Nj/fXIeGH/JND+32bVfKgqa8NxVX+Q6IlIjRdqKjOBOVN3LIBCgOmCCJu1u
kurbu/eV6j+qNLRMmpzLlvVWmbIVT/wBOwyQzgpyBwnlsJyPXMNWDlSNTh8nsmKHLs0RsFsrwP12
MZjokaqftrKvnTRB2mWfLKPBkM5tNVMPWsP2k8Jow6ZdXfkbiZyRfyFoJ/QbVALjgm+LhUBqB3iw
RMKcJrgOZiAeaMyCKoUkshmABnI48g7aHxSzQZion4AVq6DTZKWc/dP3wApqD+fD0WungDMWaO8x
vrSCPZtxIS+GZUEvhaLWe1761/s/XG3uvIorqZKa/hGoqhbS1BARkHoRlYwgPO7xDPXwAKApZcIM
tPR3VtKr/7nYCF+mauc74GS67Bv7LF4TF/7q6stdMiOv74xM9/0rSoes1jBT+dTOCe/sSwp/qIXH
w+bvwSFdRwLyiOlbRrfDiVkMFf/arLmepqs83sGjDYxrrDiTfn4vwi1YJ30xhFWUnuzvX8pIYL5W
984DP/qBASIJLqtgHo32Q9grNsls0WY4zbRmPMBAz0lrQHW5It2kSWgoS8vNN7fskPTH08YS3XSK
4ZRBSeqpmDvjD/nBfbNnTj0JZOtTNSb1CQlzqO0UHiGa+UTdzaw0GDt46wleLx6XQPI88X6ljiPA
ky3qnIWElfRa6owDYKUES5DpQSjjxGxhkurXY2PmhwbjDg6fDKSoNXOqdSHQu1MXGbNQ0lP/f0cY
VT0zDbBVqTCLA/miJwBwvmim9NFINobB7mB9uwGY8WzuL312R5Mu7tctFlOI8MJI+jSivLs8eD2Q
/ywBte84yBxyrN4exn6dh/HXUbXHopqgbTO+HczbbhgQCkUrG4/SOn8USb5SUCkZbkWDldeWIz5z
EB6HQFTUkOAGSwtnXDxIrGyAXKvEABIxJSDMrYEIzzSjNjg1Mli75fpsygjwaEz3+o0oJKGrXXZM
36fcdk/OOsLHUuM9fPtn5UVabrKyb5LiJpT8nNXRqQuJUiTp22GddTS76XAHuyGcrlAssJnn8YfY
nDE9asO1wFbJhn3Gg0EAhds8wKJ4iL1zEO5aaitZXUJkwZHm77tA2aZqxOvhTsmM8S+CnKKjixJU
eurx23yvL3vaHvwhX3m/y7DdjNatFU46lgskxIlyHWeBLbD062qxsyf8hvJMtNiGYS7idK7bEobw
Mbrc7BHPXMymrI3SY3pk6RzO4g5FsHhtOudQcE+ekD0qNHQ4hFsIheV7uAZu/V7u5YvCZIADYVwA
fEAKfjZzULjp5UpKriAXc2O1Yjob2iAlyfArFSOfBZ+LAVW5IRCxOtHYC2z4awCU0GHiA1/1tOyn
9VqDHH/nbRHckqtlDVUvcEwFq5sGzJ8jLcIBROmsnk0H8Gu3mgcLNeAm7ZwDXlYZEZpdC0rTUEOZ
fzibYHR/8SwbR8WlvylBfiiK0pOXO2/Nea/4LK2Rwnbidvzhuo0Z1vIt7pyH3+qZ5fhx/OkxaZcI
phjh1WIB3QegPJ7km492UKAcTzWxNYDEcZj7uQkvETWCiIe0oTRp4CO7eNd3Wy4+Efdr7rVGHmxB
RFcvhceAUsKuKiN7hWcTw+XCsyrb9tPQ2qObxf8NF31v39DR0AFud+F2+J6Z2caBZOzWNYUZvflm
eTRAZabFs2Dnfd0XVwHRrgIjdqNoW0ISpJ6gHE29vX1SCYx37vDq/Bg/vTcOSH5y2iYOdPIuq0vC
/cSiVLgrr5YaXBrBTSbfrM9iwCKAO9DmNyq25o0khlPIXxTddf5CSHik/HzdRKn0ZLK9kj8UHqej
8hqQNxBPE7woJHUUulm02fEw64zsuW0kpzjptYd7+RUULb3rjp6Mc5ZihRcftxAUkUePB1MN0dFG
2J7Ns86ByGn7JX24i1eUK1h//PLBNGLoeDwLidPmDc73F3hyQsYmSzt0s1GeXbETQ2qJuKoZoW1o
ubKdZlau2HA4JZ8SH+/sndWNgX1Rpcwq9Q4V4e8lTpJAg1tz/Cz15sWr866xrUhYk8GQKwPH5LKp
Z0DFHPnMUgLp2YGHFXv6Bx+lZxqAqeRed+cGWqjux0P2SWlmtO3PrBQaleVkS4zvKIEblprwBznK
LxP3z2tA+KjDGVENWxd2XlvU2P7hhfbfatF1VKCFQ3hP2VKiUCsc9Rho6/vEe2deHTw9B8iaxmg3
HpiS+Ze4MHOpnzUTWRYQtF/wDr4IrB/WP1w7zLN2SARWB/Pv+WwCjrhZsQNJSs1rkZVf2U48rCyx
11MqA/UXAmoPRDseqVlwbUVtD9NCj9+j01WOVk87yYZdbZEIOhY5aMzRU7hU0OhFTKTFVjhmDjLL
dtl7U8slQ4T9B8Ks2E8MxeMJKriCGwKuBIk0XRiO+DpxkplSTax7QGvDiZoVzgCSbLl3EYD8VF1G
fNOkhHNdMlzBI22il7vzxkNvYRDxZsGoBp4NBuZaGVlVburkhxfz3LGydJV/ho8pBi3DpSSzr2QY
rYBGzQ/VixYP+13rGV7XTPb0wqg+EdwFCuevTTDESnFxYfKIj3DH55k3TUxEvcYDD2VVY8L+t0gg
4dFOjP1gAj0/w5wjfUDfqpuotUAtsEKw0gbxSxH46x6FlhhURu6O6ZWIuCYKwS+MwhHlWwX2OjE3
WfK2426SGNUlX9UCEFj56QifDQYUJ4irESePTospUL08R3DvlQMHLcbam1dqR1ocjTHBj1SwiqoC
Kh5EDTB3olXI+jtahiH+ljqgWS7ZgJMEfRQr6MAm7bR4Cu6sr9GQ/9CwMOGNy6YgpX94puCm5S1p
hjzdGvEP1WPVcQ6zSnxrahfnsMHOPf+XUctIoPgWKjkm1PeInxC3AIFhgBDdplPkj5odCUcqPC2p
Zznfv8/6HSVudQ+iuJzOLZra/rO3lHhEDM5y8csiDYwHK+129MngN7QFSY56Qhrsj+SuIqz7pZ0B
WuaetilCA5GWAGlp/50myQh9U3aXOkhvU3pOzBr30OFCaAfFm+MevZW12YP0XM000jSDclzO+Db4
W2NweHEMKoJKo4vp90E9XxwnzT9FL+48TuASfW/YFeoJeDWleickAuBM5uynAg7GMmdAsEuOa4wU
wjHPH+f9qJ0smzNOsmVQxhz7quOCjPLvfnPOmzUFx8Pfwv4FkWydePlf3PskuUu+cHvxxmgUnGIT
nZKzg1ewAkMDmoC3hIxoaHZc6fL1K/Ty+mpceOwq2GR+angunPgwt8QdUBovzJutr5rxcmd2vPIc
mXUR/sDV80RWUA93PODO/tN9LpZoyULcN6JuR/r3HrFqe9B8V6gt0romiXEsru0z/AFzlsBm8TqR
YIDAqEn+onI49z2tw+8aRKS2k/W7RS5jvtKtniANXRxvRbGGqX+/dp7dcufBanWDfww9YbtdTCKs
1vwy28OG9JzAT2Lpm9MysJwBV8H2WbaZR4D4eygT84AWrE1MgxQUhKalTy7FjK5xltN68Uxc7AEC
GH3Hc1d8coHXv5LRvw+MUyTrDgEsgP7o4FBQ48+sVl3fjrt4VitI2G2qSUSM7b1rqZDznyMKnmu0
JwxiTcTKVUcSzkQfDqCuxn3m0eSQmXLnb/G/HUQp8s4F36S7KE3CQ7qiCkcRHE/cHZIJM35Tv92I
7/983+xHqVKEpeS0Vg2pbLbhrbByElIHoIV+PljtbclegxA8kOqj5G2PPNpn+Law1noWl5T5PuwQ
90XXoPUlNuIBVDbs5+0ExFIo0+40OOZxIs4fJAH1ViD5lhW8lQNsGtF3DqdD3SVj5+RyytFPQ69z
ON8TmywR84gOpHASulr10X3oANsznplETR34TrVcralehdcP09pzx5npbGwRWhX4DBautLgFVxrB
9ciSaWRs64T4QqHXTTL9/O+v/07Pg+WXt+rHaNfcTmeyMSBeTi/q9ifezxpL3tWqunwJM3hzptJu
3PoiG6dObBTNO9JnSE6VwnQ0+bF1s/xeq3cWHB8NFYhL9euQDqcdVfMq7PM7zf7bDw+MohjYQ2TK
bczzM9yPXxZvWKUpZUBOATe1k5SoWy35BL4uMM7RH5KKhrUpItau4W77ix86Eu3tCy9dcqkeFt2k
cVSWsHpKviGvPeVl/g6l5n40D9cD7H98FHouGry7Cz/Yw00NNPfSDhzPqt/ZY0/1/MQxMoCB8zF3
2oyQD1Skj4JvIcjw9fOiLP3fkm4VB7TA13MMJRmqGTXPl2uKCEORbNwlEFIVh1HLXDznD1P6RKYI
P+UKtz+WbElj16gUoD82LHROv3rpRCBOXyla9Urv3hq/Ln9LzvNCPPJS7rjs7PF9hVzoq0/ScIbF
jQcKXhokbtBztMdSqF3ypamR6wgL9sDmauMgqLKfKkRt+MA7xu1+DCvawe/gbxzQ9WWy5zLUwQzi
DWrjGYwToOUfqWNVWmD4R4Unibs3MmAG6kPom1YAENq+0J4YYWsPobeooOPd3vstNSyR7YQIliMj
cskyJIji/x1BQrgn7zXgIym7sVRZ+6qyj8Xcqrh0IoFYkp1k1abiseVWBedxqVNy2DabcdMqPGbr
Jt5vItb/2tS4rHnqOSFTDl+9x96ekOG3qEwIgniiyWEMw/FA3MCoP3UrcRMZgknyYt+RXa63BpjJ
gyy5IrHra6LSYTOlDwKZ9ykvxYzntpGHTpOLFk0NNZI119lfnUYMCemW8Zenz3dT0Ur01GRNjVbT
GuGmpTQ3QpIELbVlY5UVeIAkzfixCkmAkVfx7q6gOOLvLzTg8QEdahaJdM+8YgZAr6Lb5Gx3Y+yT
OH8AFhcSv8kOtpy3taaFDtjkOWVR1JiVqxRg/kS8hMp7cLCVln+P/KuECcJEA8aF3OIR77fI97jO
CoWpxYpZcPcISGia6bEFTGXWQyc16VHNfVzbXw7jgB/FLEMFui9qcbGJkseXsWu85fyyTdfoAGcM
oXzYkCZhfc7ryp/NGJrIa8nzOI6S3s1jQQvbpAun8QSaba36mqpj/zFJUy096BVslPr5KwmRi1kp
T5Q2u3isDQ3L/53esKJPKeKTkzbqGsu31DwMUcNirXfl32vvI50GKpk0izNpbtXgYKLrSL4WVS20
0iMs1w4nJ6MhIQGqnFJuyUgdFH45S1sBEZSv7LC0mpnVXbrrKqE0UtoI0x+1xk7smhydquhQDtb2
wc/wqz3UKPKbxztkqRlILYpe+Cush7xxVFywmSaVXCTMFCJlcGJZ+czEks7qMNFdgQaqMDoVHcs8
m7SkqPnZInJgNe8cZDospyYD8ZAfZRbAwhmJrPBZ04z16QWw0go9fdDQfer9QOkLgjJ5gMtENrw4
0pQcx2UbjhWfcZ2FBzKkv60z205Xc4IAR8EnJ4bH0eAPgis9lLSKsxY3VJkWcUy0f0NT7xxbazT1
+8Z8Kb8WiluYe3WxXc/JeebVMRCk01jfpu8cLA4TqR/HtfzfVp9nDWHnh+4yY3S1fAhPdevAQ2EG
pEahA9Inrx4pExljnx/0pBrYxK44Xh510jrW1eLJe74HhjR5d+WOq6Qijds5joYy1sbNrVFp9ND4
ZNRenehn+zlYreM5bwI20H7MBZLLdU6WUKsaLfJt1Gy9eAHR6+TLVOY8dh09fIsn/2BT6KUAf/Pi
3lenAJ3aMz70kpMHkbwZYffsjM8A6JZtJ1fw1qnJVA9dBY3BhFs+Om1MU1nVm/2EahGadL3PqNCM
2TBS7zNCOQEeZXMTeo82frXAoxuH0XzlEzZiln9sYm3PUiobwRWiRlvH6EWMg9etn0vaWdEfRx8i
gnVrzdBSfFfkFDqDB31pQyggw+SuyOyBtnkKD9tI1qICaX87mMJmShgCyjk/ACKOMxXhQ15o2dPc
TnvGoOXCv7zGEx33Rm48sTzUI549wSPC58bjb2HLqaESlUxnAOqKLlZxP1GaIti0fERjiqAaok0i
bLHn9aQhpenUUk9wvLm4wWkaklMlKlE4/EcyAFUu24HNwQkQEKboeX+vNZ5xmKZnNEF32/fQV8nW
+PorfkuWMke2oNurvUthupGEQNXrOl76iZyyjCjCb/NOw7URbuHra07GZMx/AC2mcr8RRkBUAKt7
9rJs0Ukw6k9lnAVPNtrRoEgRam3JAMs8Ri7df0qzLjl98BOjTrkfrTiH9VeUHoRI0Mkifw0E+z6q
8LMGrjEagrACazza+5l7eJ1YhodwLz8znPlQUaI2gJNYyNq5u826GLSbnemRrzzUegv+N/BkJYHQ
E44shiefEmWJ9JqTLwkEIf/ddbjsy9mkPyo+ut491th1xeTxix8cBQxY4gwqGCzaMxwwi5HFdFPv
DxYUODYZYi+OCmkuqQWLVZlNwFQJ+1oWLyPZCGX7HaK7EA8hIE39ctZQojcyCrPWm4xNfiPO3tJp
ZMCZL50vNdeTjJeQFVCy7WxrjeuyL2B6NRLe1znIIYeGEUvWs0PJ+9B/C6RIr+08Tnh0ndoaOveI
mcKkTi1cgU692BSrLK5A1n3gpCZo5G3YPLBbtHySm3/PqgDPTPfUlxM+5XaNuj/0vhXtnDJDiT5E
jOhLfjUkMQpwTuvcgP69FukMDFhJcfLPuVUKyk+mIRQmAmh5iufou2+HgUSMZNMboeMWagGb1gAv
/W2LXVX4Er3Z6F1x0xTB8P53aEME2cFhpdeVhts3eg+VveeQNc59dYxgJ0fH0IQj86MPRstAoEe5
JpedjfSBi346zk60x+MGTr4DTLeu5r/rQreW/Rnzc6FnoXI4edFZ3ZbGhKSeuDphFSbz0Bev7OLO
wS8SghIHGtjKUbu/ZLvLRNNwVrfBrabCpE9ngOmioezsFu7JHiHQQdLQcuI/YKDqnl7tL2aEOSob
thZijim8XXWxifAxGOf18pNWs1zRStr+w9UzzzNEsTaHrXb2eNgpyRBM3pZZz4tE0ypbMMx5wZcj
GLABXNtCoA/Z+dqhZNPtXq88/rupJJMFMbhVF1f9gOH56FzZOAB3ZKRQo6XbekcruKlH1bFCVEpb
IPkBWL/zopvCj4q9LROQyDMN6Pzzzkt4Tz+L7DmU0ds2XwmZVqHmelfF4qYHxQLtY6z2nTVzXN5G
Ct5EF74Xv/Rn7unRwa2463LaCzaTCIsquJINbcL1T8mC5bPvKa8+VPteYh5mTAuD7EB+T5wMFt+r
PqSJ7zB5DQaYJmLSX8VCX5fQmOykpXhdmrqK8ZXgqk68CGNj76VfPtYEApCLOj/+oNwmu+7SqvHm
Mev6/mzsz/yuClNlKwHWkDz5uIxJ1Xw5WdUJ+ajVMrbsd9ROLZ4iuAoH5o1g+Z84eZxj0NVfdVQk
+xfvqDa8o4sCzr0UfvasNp1pVwU6/cV0Hs9d66uBud0uoFixg2CpzsJoKbKkD3BR0MhLGDraMnkA
kgETeGbmEmxS0sn///G+s5CSzC05hIta/WmFbbFxsQgksrrg3b4dtFWeLfv2WUQH8pgYhI/CUt9L
UYsy9wudvkvM6wlRE0yR/wfUZfh65qMhVdz2yzWnHLA6jK8UsQXM0HIpRheCggDSLzCZVhwtk+vu
i783SbOfjqfSVWGbH+6xYU4VeutYx/8x2jy+sWSYXxjigLQrsnGfZ+GwGZWrwm1Pu93LjJu93pYA
CW9jTlxtu4QNmzDtjKZKOI7A4iKuHnyaBgpc8aY2tMOFEhkuTXk0hA61O2WxKlXuCdaYI3Esa7/0
AI1enE4flJWtiqthIPG5nj1szVYUcRG0GI+LWVW8yf5ndtBAlCQyDEhw3idbxQ7lpaixe+GXuZND
3vMgMfIJjrI2g4SiAow2t+6fb6ulFgHPhLt+qvm801RvfWmhjUg83iHnwpSuRwupr5nL7M0dGKBI
Fvz1Y7AwjXrDW6N5sPoKM7oi53oeS84BwhI6pxaqy5QjHQnr039v8x6HC09IwUMZvNKteZaAtOEF
dPsPWQY7bD7hBiVJb1vzBc5y1j6PE33NSq7iEkfISqH/vHr0RE+z47F3yfQdVMztH5+cJMiemIXC
msTFfVA19y7T3nNr5cZzHesQkuP+oXqOME4GOhKUyOAWNHvFsjSWQm/9metn9jpU+aBuBRfakHGR
Ei9MSjeA5R59mbom7A/cOnNd8Kh7wDkxr/eT2neQZ4By0dcYK6VVjfGNVihPkfh09qpWeO5Kqkbm
a0f444gMkm/ua4neuU/iJgcUXDuiT4E1ha2dLw/CfGKQYQnu15PZ9C0nOXi7rTK8vlrv61MfQCyR
7I8SzvNE+UM1OsRG5ESDxnIPcYJnUiHo/y8LAPHNHoA27rD1EwDKenG20yKJMTCEEZQD9cEygi/w
wC2HY4grFMrUqPRf7bua7f2tZUh7oGUwh8vUnmNwM7NRF87T3FyvlWo+KZQdvUrAZfwgCOH+6lqc
D2cBAocG1ys2Fb/TGAey7aOzRQsX69gcpTQ7Eegq/5vy3ugnLFH8UBIxlIaHmwUjTVfVSYBe6dh9
+U3ZYbx9APBt+MoecR1ZD5SrVdbAHGmA27f0eBtooTtWKYezgx7cYP+5T7+UyMs3PXAQhuGIR/U1
2Pu6dBUNOF773kn7kI3+pnfdtpCpVuEfLcfMXevC3PBmt6aEHEjxzXjiExJFSaE7COd/LJSiNMef
+OlZMNsvRBGjsutmc1r/MiET+uLmxUvUFr3IZlemjWd1KxrkIrOiXSU8yEacStn0oFMkoq33NUGt
Cmx5mgHZMm9Jki7j9C4MWHSEXBSlpgPGBz43PxiWK9UjypYvFmtb0xhzPSOuwy2PrMZQENn/hBAP
M0RRquikBRFx8z++lF5GQfJYRnbyTNqQ/S9Ryx1NSisyFXrRrQSbUTVSk14M2OlZGnKPmwppfG3b
WCfDGJu7nBOnxweeS4m8vOmwRiwWVRqxUB263i2u04ZKisTH9vQGtxHsnls7uIYKqpc6+3tCBvC3
z2zXe/60dd3ncUs/EIqHye5PEOxQXkqX+nVg+Z85ExqyScaLbWAkbd+z/Wi76+xjjBns+IFe8X9S
SpRNS2dFWMG8o+EesyovavjUvfp0HsIxjuqQGE25yOMzDBzPfCH4tNwg84Jy3VnY1vSnDaCjObFz
lXcK6YazX+eUGfgjWhc9WxME9+bc2g+tJxT8ccVXan6Gh35cTsQVzW9QxDY8T5GKjZl6jbqFygog
lEB4cOKvWWX139OO65ZSs2EaKVdmh/mSL6jhRW1NGJMSimqYErwbcKXrd/SKy/DJuwhLWDpehhCT
fNS0oF1RE31YHFmBPPt+uelNAZ9hEqFyesCdxLby/1oIlPzqEiYeJWDuUZ8wrbWQ35g0VtYMngnG
2Fk8v3qsJzBadwU9rHwdqTZ687KTpp390olSEgDlMAvYlDszz3hIje3SuOmyEGBrYD3MQoZ5ScyD
xDGCr2RFRhVt10NC3rWdu/60x2LI2Fr3zmyzcBCahl/57t/tO2Kc4JZESHLb7pzZXYo3i3pEicZA
1UR5zsAZ1S5Gwzv5ERoQhyik5lrZ95njzwVG3R5fw4NvmUp6uTF7ZyuglDlEMWkiZUtouNy8yQeH
Kq1P5Oklb1r8DSrY6nEEeZ+JYuhHqIh8i6RK0SGJ2e7KSU1SyH55Z30sIMJy8dc7Vlxe1KTuaw1E
7Iqllbu4QfiHLPiFF3mwPzn4Mzy7QfM5X9XKoVD4rB/KHqSJqo+d7SwRy/LmXqFWFs5UrCJ4qZau
pB/5h2j977mTrP23ewa+SNb3e6GTLvRE5fMHV8r7UBdTM+oFxVCr4DrhnoQkfv/MCZ3oeRWFs+Je
ukCxmG/MXikBSQDk6jXX4RR+i1Te8G0pqeAwT7OZNgeBHxyxMCieYurybI5us3ob8LyZNLMUwhT+
bAkPp7+vmbuGnKSgssjEtWXVApf++Z0uxHNA00O5IA3nOrNxB/UxKt+i45FcTY97zoWZwXBUbIcZ
biEP/oSV0Swex3ToV4d3sYyqNvpisBkGFeBWgcbQJtZ8sP55uEt8Cnd/Lc7LnHr3VFsRj0uhmeaG
HYIpxqQgTEr964pd5jg9RvQA+kHzrU3UAkfslLu7lZ50OM8IuXomj154aMhRf93eGeO1NA848hYe
nzUVVgTB22DYJouB6AhKy6stz/2W0xqSQ/63N6nCY+MJv9fuuU8AkOX/YdvcjnVn5IcT+sfaevJZ
ktkD2xfvsxHGi1/7pnRI21iBCm7lvHhpI8Exzr5xavsq85MvsyCcfjAhxioO5aHiR1Xarsa1U0Jk
tv0h8K8eXdFO37ar6ub4kbyzS598Ne0gMkCe4wa9orqKhF1gNjzNOehFsiyXrNP0vhASDOsvsz3Z
i5G43SsXflPFCRuB7kZvJBfNBxvaVajW63ZqPhRQ0Gy5lVQowJguSDJuifyPhUBUEhHAzJpqpP07
L/aS01CI+U8ngu0iWm4ChP5aVheO39oKTiNOjM6noeP//UrPLJz+8L/DBhTApsdnOaUd9OfYjtIz
WNacd+ZJbvOIobSCwJuY0qiDtKuJaChPF5DHNOzw2uAGOmQWmdDzA7rDWYFWzlkqKlQMkHqmKPIG
VEdV4DWdFMCEw0voEw0kH+i3XPD+ufl8IdfcURlPJo5oHgpuzYSdxKooerzI54gXvozm2tVfQUEe
VK+HSBuXGrrgc50q3EmjNk/UCYDq1Cy709VGa30msuhP0YvhKHphqfQEgsiQZEZL/ToMOLiQ5q8R
wDXVVrlPwzfOJIj4DshMVI/qR+XOpc5Mxh+STOPHgJjEG92SIULpfcomlRFjfwqLq7vGfJ7ACJ9V
sei2IoeHK0Ag6R3g4fHkjs63s1GPqkKXJuKA7mo6udRtIEyTDY5Gq55O27GEpKrVsN1GpkgyG61r
35bxhRfTvUclBBh7LUsQtolVtf6dsNCy3JvcQeu2/uHXHuD4ucMCX/4JGHjgsD48o4y0qagVw8dV
59p8y7NBY6OwOQdQRscl4a06jBbR5VSgCrCDHbsWtn5/W0UpxnOg0MGc+/pEJM//dPI6mTnIJAAa
ex3Xl4Yc2SkH+dUB0QRnktTfnW1h13DVes2ybnRojfMImPf4thV1J5rC5l8F2MiFEjCVx/hdGlyV
FXqQXG8J/Sb1EsdqsBWvygc/YzROfP9HJKVv8QvMDSsIR8yqakr9RIKtveFYVGmVNFPkURGEv3Mb
kLQTqSeHY9j0bLDtSsXLvzRkgodriZXsii+3yOAz2vJm6ZLPdhXAl2wF+keEP0Tdg8j/CnHKuw7U
s3AnYiNgFw83OoBAXK5UN4i3lRY2iZVlh8cfuZksKsxJDJf9LKkWQzVv6rcdq4YsPxMFtMSIMXa2
3Uhw2ILFSfkKIQe6t/RqmcsAL8Ll9i3+Mns1W/6G+6KX5qYZZFhECTU7GPfGreAyA9OxTQ26Njiu
6tpq6AYLwMdHLMphr9OPaDNfwMTG/EcurkLXyaNsF2iYHO9OMquw3gCj8B4iidX9OIKm9TWVGJQZ
RgVzzvib4WtWkdEcnGncSFQmDJYareejwBJx7NMwKpdDT+U+2gQ23DgroER2HV6JorZMa0bHJkjJ
uMTojbqSuubC2UgIUyJXYFwikW33u19ar3rru6ctizyZfodrS5lGnL0VkOPJ0ebrtyxZDPI7h9UF
3EA1p3JaKU4aeTwsZeOoGx2zpxWgEhhFg92uNuhpFtpNjI0vRMxSNyd/+mSiS9JrGOy78rsYpHxH
jSiyT/FlfAPjnRGGszxvvut2MjSwPlHeAcSGidxR8fVjF43tyBqhYWCjCl9hwUJuXBAIJLEYRVca
BGaZmZq4iqolX4y2bptdOT2KEcniQwzUaUURM9hHDaxB32XSH72zAxHhYHgTpDi26wPSzZflLNVP
BEBONu7jXyYsvFHjH5/TH9v7JCm/bN37/E9i7udtNnOxjg/ZuHv8tQMz1LtBr7Np4H2ER9WteJd5
Vg9iX6xIsnc1HGYyoWv5Y3538RjP2n33crRX84B6I1UMC0iTxdcKUnLxMNUPHi7If7InqRNra4az
HTxX05fRc2ZQMuja/YIAgK17DPxXKtPl2Ff9Mk0o2mQCBioYTS+l35OJuQ/oTXgk2i2meivSn2cC
jPrjKvHzuixnJcOuz+YVTVTFLhCbs+TBJHAJcQaee2YvxgTqcFULRSLb+jEc1HvyQvsaDieDEqqK
6V9LVK7HJpYbQX8JdTzC5kHZRUZiv7Wl8zWhf7DAR+vyko2R/fTxm33qkxCamC5a0hYcRW+OD/t9
QUpZ7NYYvna+7HpDMv7kzR7nJspkEoVCdrpTTMmm5Bzev+mMSCbUdRXP1aXvMzjJXPik8Z6AqFGI
RYA1jgghtoiRdTxlQLUO1z5xXhoWJnkO8/T9Iw8GuhTwjFtLqoD+ZmAG15RHP1cPlgFF9/XymlEL
mT+nlYnjY/rajOQndXhMbYCIB9BUBHLub7ijy1Ec3D8yGEfcmsQacClRaHfpTGlskqL1OQkX6K0e
BMHx9Ykmq9af7vDPcblcDEepQMeTOLcc4ABzXCBHP6RTKHkjq9RnPHxpwLddRApE1dpvDzdWrApg
0pejx9iHvzJdrUCdYdUi0tvaPEretnC+C4JFctQr4K7Wy9KVykpafIXLqt+JD1wucY6/B/mshdTz
CydaTtX2f+JE76AQbOMwOlAcvs3TNn2SI3J9prU3fBd6I9xFlNkCvScG6umk5DYBJGGYlPbZKoN8
JsCr4XuGVF8EZxKR3ZzKOM8gtoh4MXo9++2gYhrnPBoI27LUA3a/RHC9soYgER69qobnDLQmnGzz
7J6Sd+dlFfvaSNZXf1qyRnVq8jk/Xct5i819HDmhV2FqJVkydvd0f11VkFkf5Ix7wdjniwoSBYXK
APgMxXAXCxx7t0o1iem4e2wH9AZtHyRwfstoq+QmP/xxUyu103y2CA1nBZ7Hu2BXdb2lw4xWp+bq
GBB7Qjs365lQFZ8GE+xrYfkzZWFF4WU3H4EgDrUXTZdIvSE5Qg0v06m/mZHknsG7bwYmJ1gnaWdh
vnhD61XPn1+2d/1Jras3CfI5Ie5Jy6I9qXfceN0TYOs7MNDDDUqXNOIOsyBntUPs89MtKdFlwGDH
R+szliQVwJ0K2HjpcpQu7z5/wFSJRQXVgUe7AG1geya8NQQ+XGnepwsmKUPmnXpbyNKHNeY+RAt5
EJjzHYLhvW4MEutr20W4NKyXl0xi0/fzMTEGp8R5Bo0xwEJpaR0rcv6bOmU18uVJWkpYDLppKRlH
fywhWN1hhSBMsWFsmmn0r2jR1eNRBm8RqEbd4ZaODsUhjINXlMv+PBaljkJX08cyqihlgu8r2dIL
Rum2/XYHVaz4VX63wz2+3Dmt9YPZNfRb7lQo3nD24GFUjqvkYwxj8jvEbNAPVmK92Nae/CwdhgYm
uY+kQUFm86dk/rWfHUuJKbB5JcmKcyVTj3l2wqx/GeKSKDkms5CL+K1dux4HoM9hIJ94nUNkzKHR
zkjarZo4VzXY23u9YSlOxNYeHtemuBJ8g8lysrgYwFqXYIV55kd4wlT3X3+vhZa5k3mzlLIAw/T4
eyhTPnZhy7Ii5VhhrUNBuEhHGsnybLzDbkzOYBr2vhSpn1TINOfXJfW0uu0DmrDgzMidfuqFllxN
mFv8DIwt43ly1CfsPtabuKiJMCY58AYBbYot4j2ozUEu7uE4eBUYkN+pcj6bv+900UaGX/q0UhX2
bhhHmgeAKfkqx6hBkcGeKYI7DFENtAkesoiAAyFO3l7aOy6VZ4rs34nIBWtIQ6O2IXDZRJ7gANmd
aB++vVUetj+mY/7CRswM+9d93qU+vGLdKdHXUoqNtvXuqfksIVVi5a3bwNlHbHylHISj/AIPq4cn
a73QVfjykHBlZ0hGQaFc3ARJiAUdtH1+Id378rUBkslXbGYGPbGH4tvl7Me9aEzjmvLv75eEfQgw
mGujORndxLXzPHFHrI7qTQRYdZo54GDDd/0q/9BMubTXjZbbFxU7WR8utJQFEYVCPrZSzJfzLCo2
blDZ0fE737VCAfQmRVI1HdAZUuA9uoB5AgO8QSiz9sjAwzeOPREJZI5L4z/OflffmOOqNwOOqpeX
XqPBcIWsehAXEFeqlIOpoR3FIHjmo7WIvaBHQU7SjwO/JBfLyacImCq4CMwqkZMT/YxgA/4DiMtf
/4rUni61fTxBGH6rF+lOgHZzQBcHKxicB6UmsYjYAfKnMRnjR3a3wovwX/kwJucaK+Rrr2d9k3yE
JQg+68d/XV3p7yvTeb2hRG+/6rzK6B4sKyko7fCs+s7ZDda5x/fes0oPdtTebpjOezhU7GTSAXNf
ZflWQCPy6TikRLOixrJrrIQZFnYHPYWPZF4i4T/O5VMvyso4rLx0Alosi5M/NDG3Yp2ugA4kf/0o
gI+kGy041Uzo8phxGCyceOnLzWhlcQqA3+vggV4B7nVvLMF0vVPVwaeqtxG521zcv1ZAGy4csBPP
OijtjJvBUJA6tTuLLmWGF6d2P11MhewWOTEHK5DobjkGwU2DCOj8XO4/DX+VpQhaRH/JYFkfwhWr
hmGm3Le1mcFcj5ZYkOrh32jZ5w9cejaGAGfhX+5a6RP9sXwFnVFrH/+daNZlKhXFO6iYAwN5R7Sh
+iYTTF/c8JVPHczixvq7qkHUj4yvKzU1rSXxyWM3CXZKM2ZdZdsSJ6WLKsL/hPsN5q0K7JMWO+31
KHp/1zUN7V6iO2R3a1rcm96lFMRBt5DXKwpNql25YqSvJNuygNPus/Yb3uyaivhY17Hm438XH3n5
FODY/F+FeiagbwAfJ8/Xkt0PynRUOsNgNGbBP4LcAO9Hoh7JYGNJFSiP9s/Z4xGUp8uPxQcMhgK/
D77mjukpHNZ3VgamVMMEraIyivwvr6160E/+VT7+/sFOYSL3YQCBfa2GHxPLdMjaYnslRwOzLJOD
oSjen2V12RHDh/prpVLPesJxMX14iMghcLzXMvjVU+y8uE6Q4ibuQ8m9yXUoTK8FXFt4PJNrJvOD
m3gMBlgYir5PBJCLIXNXtjdS9r9gPMkmVJXUwzHPIZniXttBgHo4PDv9ZroYWsoOlsgLXIDg+2CG
lWsIo+u/BzVJ5H6ps43SdF7UxKWfe04GIDDgXLQLcQV9inLOOBdhUy7dynhEXpVctnhy+iDVt2m/
6vdaTHPFLoD47wuW9esH2shvq3J/3an/+WbriQ0mXo01vE514LX37NcATnNkrA3AD8YUfv6UsAqt
zxGM7oFz845x7CLHd/Qdmw0ONl6sLO5b2snWqoIBWhDFZS0ok8eNQvrN7PGvw0cuNA0Z46mnLmQF
lT9gacGbXfGIEbs19/L//hMwQJGH8+lUJORO323X8NTRQhPVe82vbhwLGdptDhRMKPSYAHM1XvK4
rg5mPctT8fl8kq49wH+nc4IbyYs8PUpYC2ySwMvGkTjYIJdJcNnPcTTjzvUOzZNFwPNlOyKXDs2t
NVnvnurCF52ct0CKhRE9T348BZAp+wKzPrqHni+snS+2RHs6Gq6VqfrRTqJXkL0Y+ZfLhwdpegnc
TgmQTuo9yyM1D3FO6kQX3y6mJlaf1+4a5MqrtlESnCOwUtovRHa/tJAOKpNr4U4+S3CSUEdUz1iD
/NHtvN/7qXaeZ9lnKa8O7MeKy/cq2/ixbmInQ90Akn/V/LplNG+hBTYoXi/T1imr+6kEkVlI68M+
Cixr89+GDeqAJmwfDLm0UHRD73XOIvY2L9VOX1pmdwHJq5Nj6uIu6xdj47Us3rAFgc+miZ1NTPIw
V5kFHoon4Ajxm1emJgmcUOIkRi5exhYaSwdnz2YcR9FwpDxsDUFxkQZUhSvQ09qE2S8XB8d8Wfp/
yuGQpAIpzXuqBJ5c3N4/LPskzEy1H88rZmH3/JqBvB4UyWfcSbu2/IDPmPckkpza7Nk/qODb6S0P
E2+xK29JFzV/5YluIoz9/9PorunRfclY/u3QggLfyFI6vEqp5fYL70wSw5+saxfILuhmT+Ab7Wv+
2QD/amOmFO6DVbRq+B3y412MtCP5YUqEtS5J0xonnuTBU2SuwkJPDwNUYzTcA9JiBhCRDOSRedS2
M0GEuka0HGMv67UVHGxG0dXJMwzqFeg1HxXyLKNFtW7duUIoUKYgXUON5GT7KXYEmispfzvGd//0
w/jGBF+yS2XypcMqXx9Hd0HKeUMPE7Cia7LIv7dcE/ASVNm1eSCFq4mMzuEoqJvHouZbPYOP9okM
OhLgTnnceldntkLzkWi7SJ3YuNcAbHZnn98/HTHDN+JtuNhald+TkOyCYSDuZsUB+dL1CkPwl/PP
6JBYWtSR83mOMfgcDLl+y4/pYehth25FunFLILY3y/xlc47ZqYcZACJmAvGVoGXpsj20yHmVN3Ce
tszbBF4JhII/DcRAd5Z9ZIeE5wSL7xXngppmBA+YOReO7/dZ+hPrh+sD2CEmKP9fEX7AzH6AMys1
bR3R4ZKjGLmyxWIND7E9StokTkZMQ6Z7QbQXzF5SPrr8p2bRFpD/JBxbSCS/QM4Ias1X2pdI4oxI
T6cJyPS7s9XPih1DEQ3tlAE5IQXpkZMsAHaKUO4b21GS5Dh+k/F9CpXnQ5Kjl+612o2scT9fdadc
64m7YuQ9WjoZw8svt70X3GX/0dqL111ou7nAHYinP1mViiRTdiDAF9g3IXivNmt3LN7L3aHZbE8I
9JQXnBKK2MiSeWc4lC0FPUR5OIM70DaUoXBtZhOVk0P8ike+Z3OJpxIJ8uee6vvEHq+fvS/zqKLs
KI4d2l9rRqm1dDyPk5hJ6hJ5D9xWU15jTu7ippv7XvSL1g1ppSEUcjCC8LrhhXGgPt2vntwrPqxT
4anlByFLv1vO6EVuump4B9wabVmzdu1B4oWIMmUk1bsGaKBUGt4co2oU4cj2ReCmcLC+gmwmq8PB
i8T/m+dT2FqG18tliiHqBL11Ei1lh9Z5F06J3YhvICHainWR7+/XtR5DnFeAtuTFuZWwIImldnxA
F/S9vK0a8S5Kc6s9hc52AXE4CoB22EPAiR1+3S6aSkacRMl/6crOxgWINO2KDt+/r2s4L5liPeud
SjJquBoJUnDpYe9mCpJxsj8qqFVQS5SFH0JkunF1XXhIivfyADY0kDPeTn/4Aqmwj96zJiWFDVNC
bq/5aAYRW9klLL8vGI/RlHTOg4fox93G2aDNRoHOks4sphcYPV6BO4RJMsBmKsXxD/AUDqWA5YXA
TbIlxP0NjLB/ynPpwqu5ixukeiubqApjhyTULW9J7Qwu75IBArKRjHi2UvnzEhPrWJxLDOQb4a4q
6pSc3GIYWHjxClbcWNSknA2ei8ZAfjK3L7HoZ4DWrtM/X2sEq6ooaLJqn6Tt8mCn4RTKKABg38aU
pvkcDz5Ei232jHkyEQj277cIUWH0bvfP1h0CJBZlC1O0vMpnBeBszQd4RrkwcLHOzJ3u0Jd7YGwi
1qs9Zb9x/dzI1WUSoN+ik+3QWaTqo9HFZsq1sZGd2JoVdVR8mYVRf3uTYIBsV1lCh7ngfbLPgYty
CYf3cgYC+XiS4TFcnAqDBwzrfidxBfWmk24eLzmHFLFhc4CB/+rLD9q+3FVjrkdmj7QfhazT0eCC
poQcxStdBD54qgqgEtbD4qKYyw2Jc8PD7L90RP2uuRtNhlPMbmH+XdkYrMZY0Kkh7sJr7ZpGXfz+
X74tgttuubzbBlZUJu1DjXgszbBFlWtRJtmP6BjqRt25l+6hBrOfzCoHMMp6nUP6Fh2K4nA2ikzC
Xf+/YkFofb2tptTj4bzuUnDCn+TW86slrAjDyvl4GabbP94BrBrejZeejIlBbWGOGA2VQhMV56ng
DGAFZEjZdX7v+RRhfwKCmr+r6q2NVBm9WJOsH+1DyRWDFeiC8tZs2MdzbQvvAsUfZIc+P++ez931
L2A9c7yzfTUwB9Et8QdiuO97FggwZYc1fTYu9BCBBzjebGDmWqurzCtL27ffO+OyRK0eIKc0M+IO
EspQUTwuYQ7ccjs2wbZO0nMQlNBOBeqPCl86sPNbjYmGlEV6FD12yuQDlHtaW7EhcW9NwgBS5Amf
p1BKHqkjSMll6f9bCFGE0U6sG9MJW+sJXaypwB6igGzOU4GGVWVjKjW7FVNofdYutFfEUo9BREq7
2zdsFcgaKBHkAyXqscGikUrA9ow/ZZ83BPMjc92dtY9WnmWH5ZwJvOR4yz6KfFyv5wvdLtV/K8/+
3gUmb4bn95hKU/45SPr6wV8Zn/iTAoxVYgFWCEm8HGC4gRe2PUES0R9aoAud67gI81HBUt5iF5hS
fPgD3Zaq2I3MN6or8ZEIlIv09CqjKCHmZWysyessUbG7ZcnFkV8Pixsb6Tq9VdB9bkvvK2a5gClP
ysxa8HPeCIgi8koI4onnu7bJEgLZN4xoyaEd2epNf0KJNI7DidXE07FbK/ZW/bmpSUqvarOKFBzj
Fom04KbZv9bgTYGNIKe+xaw9b6d4fUz5D84xGwXKKf8aGk9m4SjCKXSSKCnh3P091VlmjcwvDsVD
L5ULnuW300RgdZq+FXmyJxwB3KGwUKkmtS3F/78UjuNLMotFo+8ps3xI9/bbX5BeHXQb4rFkz7Bj
rg9xtM1t0Gd8TktKR/RRexaRCaivGnF0YA23hHU7XZyZe++swUVO8Dilld03Awdr4AAwqypanrK1
95g3lQwUASASOyTqU7WqUrj3QYSPDTHZvnr9xCLkWXIGrfTfvWTeyuWCmDFLxeK/sJP2I52a5boH
EKso2JHGkDWgKxhXnxp70FtPu337yQcIZgvPIblz6McVj31HsWyL8A2/BfHdTmAQ1VWr/vjYe3g/
hoE5FpRJVrgbMgfQ49VDWiZEIucaZSnMDoHWXPSn3FWrD36jw+H2xw6lypQ/ygXnP+kXZ/AZngXB
DRp3uqSNhMY4I504TG6MzHEu46JPvrLp7cC2RUAlAocYn+iKeI9xZTzyRg9LIPlRNQp1wJeCyQo+
GLDceqFgnvt8Kr4MnVOQ/yh4uqM97bkxIWXuPSVsvvM+G8slXPO9Au2dIpIjH7JzBsBIqIyIZwpO
K7XUQdCCZ0tk/tMJQ8LSjKpPZJ9aneGraWjpshDJBIE3V93AB3viNdelwJ2pjBfXZccNf+rVSiAq
JSb2kh5dk3edZlTIfgoRCy5iy23joCuf91tKYe2S9StUNjjbmkB/AC5JJ6gk9tQdEZw15/owyGIU
QSo2jBUuBdcuuvC7gnr9Mvt+a9J06W3RUaf0380hbceiIgBc40ScXcwSMApXEXLqGoBA3C2xbUk2
DVsPw+nY+6Zzm7ZoCtsc7LQJmlBzel/sBt4gaxvToRCkkmyKwmkAWYoflLCDvTWasMd8U5YuGflc
n27jX0PjscrJy6wtQHyUwcqhOq2mFmwfkYXiy6gLMCLPqYkMrsdfAwPXpAQ/6ok7EZOD0URLJn2f
lnclmt5tChEgvmZ+3z4h19WIv+IgoK/0yp//mjzUKE08QoGxDmDOoeNtT6bIr6VrGw1GpJiQWLA/
UMfc5iAz8grDoKBSBQwqxAqhFF+d6vJfCdVEf81TYRcJ8BpYGl5/mUUnGdf4cjDjf+4vIz0EponO
ZSHPkhNQAe2y6tc+zqtThxRw9H0Ghcn0bWZp4wERzEMacdTmyd5NxAy+Avjs9YMfyCLbbuvh0jKU
xvlNdGuDL3k7Q6f8Z0AVLYicFTlwMu6CEgHD3Tl16WFrgSS+nE9B3fWrpuxCbN7zecFPoVkS113G
cavcqIY/RIrm9Ed7DS6jW6UCcYBJ4FjdWSOaeBhCDW9g31hL1JS9jT1/vCjlmZQm7OmRdZwlGNFw
DfwOcot3NXIq+OAKFcLulwqU3G3vq2eMSX5IMPkl3w++TUVjlN/hTSncC8XL0JgE8pgCp9DwQYyU
Z3OLnO0ypeMwQpXck4NYzms62dSF/69GN8cM0z+COT8aHKou51AolM8d0yI+4iK9YDWHjB1T7W0z
EIhF8Ojbr3cG96A3UQjvM+hbOv1V3ovc/WMVJFoLTk13qfFZAPV1Qb6ZSZZKx03/kylwitj80PJJ
hpn92ZJpSU2KlCV1voShZVgcUzPbeOXHqXB6M15hCIhHXG4hVCg8bxgEpFePA32PFhFgstYnQbqw
EMtnUtYF5mXmePTeUmUPn4XA8DM7IE9SSDWgiXKOzyoCL0bkh225/wNKs4nTKYg5uBP7938OgwHM
yyWYShU91YR/CokWUeJ+Pq8asFecxg+uzpoOuQ1pHq7pIWTLaVoLH7JucnqqB9XDDkyvugna0gF4
vURO4FYU1Y6Gq+2fyGuc9MyPLPvyeNKo1A/bLUS3ORH1M3XgBcxM+SJapkAqw0Zerm084zKLLQdK
fph5sC6LA1lrM5XMzAZwsDwvIizbIJcqREvL/RP7celtCVeAWk2W9d1N+iCowbRB4de+V/I45s2a
Gua+NRRDX29YzONL8o+MrJ6gafFqfkrJq017wfCF9MqEBfsDdsDcOSbAAs3z9/MjjTUAmyLURDal
SV5THyB0MqmBibn3b6yNPc+MAL8RtbogvBajSv+iGwywhQeS1OA938St6S0jJ3UnoshnFV17qesU
AmD1J6djnLMuMQNVuA9HRlMnNIGmHK0PUs5+dTSLkcuhXNIPGD/iiJxy/iTAKOwIVPQSuPOE264I
vWUaWbEW652wORYS9IvMR9VAJy9Xu5lk6UjQSU7LtT7pVoHcvlWoh9tp+J7rMBHX8HWizu2vYSyN
2QMzt7J+J7Fv+hQzIdzTGs75LsqIi742h4W1DYBfZbQrc34b+aVjT+ysL4OMNhDt7BQbQN57kg1Q
kWBFsGvaK7dWihOY5VbgHZJV2j1iS9bc9wh+NJsmW5jUPybHRC0rqSMDm/23C6OzkITXvH7BjbBd
pb4ULmyFIgDoAR0M6pZA5zTXtt1cn7DSb6+oKPBC5BD5FuMcELDjYD57Oq0bwgSKLSAj8GSl/4wL
0d7q7rBpIy3kSXva01jXof6+x2SeKtGPt6ZzJfLRIjSt5+s1D4vYym5Ujk2wx65uRy8otVEwdAb2
ZeMdHjplwkB/QztpIidecSRYzx9l1GKmP96BkJlzvBz6OAZatQmcYA2xN+HHw/zN2eZjqfybzpHi
IiAVySowe0Ge3tVLOPNWJPerDqXb8HifsxIZhkgsIlaZTqeX9qEvlgeD+XHRpHOTB0qxendTKRZJ
41x1IdFy8NjBUcmtC8D+UDfMLwq4qbJYFGVt5Puox63udmP+kposjZIKp+AawRvmsOK2krsBv9So
vHHQZhUy4GX4pV+JhzZ7VObFCE7ctUIlRKwaNtwkeUgylnUAlDXMsxQracVfxLZ8xm/owTYtsvc3
eMjrug8OJGFB2MqC/bVgQrH/w9FKZpa7GXtFsSRw6K3ByH8uHLASfzuvJExkOc4+WSHEYyICfZaE
WICkkONNPNJtbGaCpOmiGSkdtPohDtmffffo52nim+J6a6yhbJMOneRNNf4JIOTxZoltwunUk86Y
fOiZ9La60pdCLO5w8Qyx0eGp8hzH8xmh/ruyWC+XB94MhheoT4Updox1udzl6AiIcqlGrisctuI6
iAm4S141pagWxxycJ27cwBzjbvJFPl0fMb8VNUGChEn4rQG5B79JZvkqwsEc8hDzffS6Wc7pmFyp
HbhJwa6a/+ALSnQNECjJ51/TwCGhuCmZ1+v+pjUEoB1ONva2NzFwvpd/MqrgrLV1ztDOsRyULnh5
n2N/Wax8rkaqn0oTX4ghVkVvL/XHCbJqzeAEovGefM59hADoryU+mXTWFyTQOQhevv1Mwa1ZNXxX
ZBngsj7GAftj+kkKxmZ2usthpWUG2kJ5VpALv1BCBvS5uETbzTFZq0eGpoPPn3MRwplvsEFre08z
hGXh3Go3vuer768eQN9vOzh2rKEbVwphTH8EYp6P5IZTHeY3Q5pxk6ZspETgLbpPAf0XA3x4IYOS
wmk8An/z5oMfXTf5AFcAujwSu2ia+P/L7TYRhRD8igwgKqT7lgM4s91Iea5JqVT1jCQcavrepMjZ
emMxnOgRZr5Whv3BWYrP3APH4N6qUyUPPbLnmlRIpnFSIbn6y/UaAvqeu20idiX34HFQcYecGBNo
XIgFfN7TYQlLa2rOqBMCkruwudOe01U5xxQGw/MAGfPZXe9/aakApPLwwCkTSna+i+mG/qCH8TwD
oAwrbFTGK3RG+KsXwF52Sddrbwl+a1kfWw7Nt+k/GS0hwKYa/uC2H4kJFw8dXIwOJrmUv/uyDFyL
bGefT426dVVoYs5KApWd0Ogf17ZnAQ62MKq6gDDZ5dY/H+qHIM6fqD87lpPNkuRThP78nd2NB/6X
6zIFIemvuykaUkw/uAKr2i6NsUTiepSsTOD26kiQroWkgu+IJb4ZvFBydIXFq6jG4FZwiwXtBrD3
NI4n9xAJlE731ZougVoW5uaHnn3mCJRUhuNjeZjQpyDAjwIWaAg7jCM4rUM+qH2WyZ46zWy0NMyD
1wp8N/SWvaFPe2rwDJnSYBcSO7GGI3kNYfPytEf/3Bx2xHYE05Fpzvi2tnAVyvg00010nf5Co3Ul
LQKULllTlhBpucER3Qtj3M0KxSiKnH5KIB4TDuY6n/Mz+YOmHVWF9k0Orve7nAX5s/pG2Vp7S0sx
e92maaur8OnSl2oBvAJG/sPWZzVQVOqceQ3d7XsT7WwhYPJhUVVCqItGRgrmWitTenkEjIqDoEAh
sbdu3ZSpRNFzbFoxloEKkR09UrrGJHWDy8PE8HDZG7OC+eMJBNqbveERopf/3FYmc5tFdbjmcvL4
fU/3ys6pFOY0OET4TVcpewaiFf4xlCgE8HqZhrxeSl9lOQ9tjpx0yHKCU08QTFwZEREwabPUtnGD
GA4RWfhN8gUgyBkHyRwRRVVvUaBYTj8tZYmp4Sb50cVmbJRsULE/NeTkPZD5okPN8Ec3UKRxstbT
EI/AR+pmdYkJyKj3nbvVIqXzqdCwyLhqfFhiBnxt3KU2OY5SUosFYYIEQIBMxDMtdxSLiPyPg+WT
81QIii8+IPBbKrDqa3sUOcM8mGvrAfOh/m9kBrEizZLN9DzbT4liCDHiW38+TF+KqKhv2Bkr9Odd
AKNRkjHhs6amuXZ1JTcARAaDo0R/SeuiJK72da2+waxn5gc/JIrIsfQ1AQ34giBZGWZ7xExq10to
aRKgDz+sja4t098CAcApMvVDRWTuimn02hkn8/Uw60C7vksb+dVt43LtaDhuq3bhgLa5stOlaR30
l7zJodE9RQJuWAeKUhAHv+Xq3A9ATcxhg6inCgwa2HAfplFvLEzCQAI0t3Lekz7gblrOTxCj+Q7H
7aRBzWJecEzhx8zIZxxffoMn5Ifk92iiTrx7E8rDL5sj4uFIrYu0YOYeHcJ47DWf5bATWR0zD86m
amMcDwIOOziSr3vrq7G+sIAQvGDGOCANW2IML7jp+X2TUNIqBvGwO1wyu63nvtyG45qOKtvcSBtZ
DnJCoZVtlcYnWYfwJFx2aX8pdptx2V/od37pPO7IBZGO3aeqs5kjrxRBRzF4Z+9avTCIFAYfi8hV
ktIIL5WpbovhV9alPZCr0WYcr0l6dyP8wgw1oq1cTKB2F14RSJkBQT0V+HVFBJ17X5MJ1dX6meOO
J2JtP2a1Rp17gfWlgXKfYdZquhpUHCJkdcimIwVL6f7VuNySvsW0oSE6MOv7Sa4urhnMZRPUC9aD
9o2ZKTqIgiKxEuqlxMLr4nrqgM8MP6Y6U+B/8ayNw0nhSCqheqZU71wkbrPr+WiKp4wK5x6VhfH/
j/FLWfN4XelutntxaOfd1W9Jfpf47vrqYEgk8du7WrkDjUCdiQirlvBLKuzQG6+747LlsyKMvPK4
23sfluNlHFKS0L3HdDIg6RSn2ywgXVFjW7ayhbg/F0Gr8g7HarmPTo4xXo9HIvoYWoVcAPYz9mL9
lX5hzS8WMiHdv/nISM+xAqEsRFie7tX7/H0PkZomSTglMYmEHuGyvoYGuRMfrZgCkQsRwhtZYeJZ
+QMmTmmyWNjRH8uaWMWJJRmj+mmvC5/NozAWuS5TUecGcnvNGbug4nqYgDwK7O3tCIt7Va8Bs97K
2YnJUPyhSln4KXOtYi8dC1/963qBHxA31KoIV7iJzq8eqtVTJiJGNnQ4dj/dkFravqV4sACvJVg6
VPnAafYQ/wXCEI/FZn5NBzi95jmX9eLu03x8vG0KpESnTlmqK0EwZaRxRYaGsij+BBVspAWdb8RP
JsviG7ZNHme/OVHGdtuObEbEqoydLIucwSzOmGtBRJqdaez09kI6fq5VW7/FV5XBiFQKkvcFoLuP
/dPLHLC6J79D5LLgOHNqSDH6mCYYkm4AuaSMvqAQs1dmjddIFeS8Oi/MS1ZcTPMFHGjlneBl/2bv
dp28ZspUlPto/ZZlo+GkURlzOdrD8B5wkQgxG2PR/o0r4jNzxIhB50HV88hOlEPNetFXHsIR+5oH
i+KQX0+iPIhy6ZNQsBSH0ajt9RJB8XIz0kauXSP4YGVHZMmEZmzmA13luJOHUyq+plWu2BRZL+iQ
7maBBEC4+5xPznjD1GFFxRml/tqkmcZ4EeMNzdfGy0smk9VHtKkIttJ6oTlB08tO8n5hqNaxUXNM
mmhw83bxqCfxPrZiAg3F74QOruZyk8SWH6Yqz0c5S0vxYkMRdsfnawhrvyi731ZKq3voYGNTPGr8
IXlyCeeh41X2+u7EBrmCOt3BC17j9SQ2hJmyRxDnO4revArkB2ZExvIHmPq7+M84YAvWLcEACDVQ
B4bMKST2WwAutpanKpbggPf7EVcq8GHttNRu0SLhbggkLlb0sQ7yD6zGUQHtYI+oHTnUL7vzH/j2
fbhtrETetfmDuSzUiTAzbtYfA8vCRHXJnQ+aBv/pvId7BsZtM9WP3q00rP6p9kKwDfjd5b++nV1u
XEmVGtDuwaKujuKSC8IGLWxAPZjj7SFAtbBtelJRUXZjskCG0Yu35ODro5pOS7yyiYNUtXHG8oZw
u7K5OAoHf4ZBuciUZN1sWPOO4WvWwknb+T9EMT3PE6v0BKzHTvCXp90eAZyJvCg0SXdgAOOaHNWh
b52QKfjwNwebsb80EkjSKGjmAZd7vH4QjGwFj7GnMq/WKeNwNaYNZ8YZnjhi9X58t/Ys0dDkzDPO
ZF7kf632k0raoUsGBlQ/eTkAGeR2n8OB2dJJVnzPdGsGr5HrN4cBiuGzqHZEcb5nvKzuZtCZqkRm
L5JAKbz2qkCUZViQueEmVNDKpHGHnHfJFhry/9vLNInF9sBR8blf0ODXQKT32p/XfZ0VsYzBr/l1
fARWylE/85eHBM8bPejiCdeCsA29QMSdgcFgT7kb3BXZILx3e6bZz8LbUbprJOs8XjrJxvyU3yMV
yI5oY1BIOAJYZmJtlVVrdj6lBu5Zfu4qdmfJJDk+mhLz4LyiCSjF0w2rHfRT/a9/PB/QoMnsD547
CRndDwccO3J74NSL4WawonV3Bv0GksSVQdutKUlLRiX/SW18GLa9KYajZhjLrBGsDOObu5m22GMp
hBQ+0h/aNtwi+xeAieGCRWLKTButRK5Z5cVUlNyt856XWtQ7vcFONMo/QkL49cu1d74ad7k0oj16
e/e8ugjOH2EQZowZyeyS5I9AXTJXK0Hslnjz9QlTWVlrXidPEyM6TY+MF4RM6OgwDzA0Mjy5S3E+
RFn6zLuj7Gl2UMTxNxAB1BrmedajPTIsV1/0ANjevz6e7YttEciE5lFkO7H+nbEnI6SyTVBCJRV3
8RwYKCJNXmpvNcHakbmGL1Wk2SBY/3ygWAh+2ACQF2rcgAJ084BIdelRX233n4UV+vz1gPChtfAd
yrfUWGcfT/SU9roU6Iew7zzuRSgE7u7C+G0J0TqdS69p9ZTlIYF7BRJ1xjC3InLzcvJpHg6LZf3c
g41iTK6Sm18Hi36WinyASmTO0EDTd4ITFlB64KhU0IyJ+qyP7rI0wAG8+mlBLG0BODJ0gSugW6kQ
tABL4tgchlQGgBJjhsuL+0MW540nn51x8YvdbE6yrNSLTo3B5juQAEB7NWu4uflGZ1NTtFbVZ6SB
DAMpUkVkGxsMq2JBqEibwvZe480/0djSpwAL/QWa9clA+Dsr0PgMJGb6lnMd3MUZ5WDFw04HlGGP
cwSH3kT+J0hP6M/cEhJeK5FHIySj0opX0ewvFohO11lqTXwnSWY0G+O6V70htstcZwv9ahlj9EMl
kTZ+8vfj68iTXMFFUmp3iVX69x94R0ZYTBfq3mIVCxkqnek8Nm7U0zDzppqwiENT1kQNM6zAE+8q
hkwAwXlFcKfhkXMb1auajbm8Rvq4f7GIta2U3xB2FU8FmUmvAwPTgnM7yX8Yfos76L5iWOI7z4nN
7czSnYtdlz5t9oRY1V6PAkUG/KmfMlzpL5VQ4VveCBE9U1p1s1GA9eXx4xWEJOcX24MR8TeaeLVz
laGukiW4r9PwXLE1IGW/9fuzapheiAbaLUW6SGKpHiCYm6wcyns78+/6ehPuTNekFxRLB/ZPuMNF
lRINV5BVmFUZc7lPIQZHupZXW9GIFwnAYcwx5E9vMEEAAgiC4+4KyM7yI15y2eOD3HAaQo4Nc5ou
YY7nuaWhTVx3L/39BFrNQ2LdWVCdlOTBfr1fQrjDvk0Gj+9tjBCdCYgU3Y9g0xEwPIVqxzg9kPjd
rOqGbXR7Qv+h+P51o38OkG6HTtPwesxutmEx6B6UcA8L7yW+CZ1i7q0eF9ZQIHsgLGGczF974Zux
WeWbLoYxa17bg9l7UBvZqtVQApPfcS1G34f713bzKu8OLjQfQnSEOQu7C/97fymtLQnm1wMmPL9P
bVZqwAAmEwozr+oafi3swK6mNpM5gn/PWxDpwKHxDw3U583gdj/roXX9SBWVSQMozEAKVdBN+ILk
KaONPbKuZJa98eYSM+eTz/STDTcnpppP4s4Eg/ZPed2KVDlYOV0KviwQdauplsQG7vKKjltonT/C
A40VXVT6Kh5FtobIzyrWhu3wqqOybDXlD4XxpPzaF0Vnt9s+SMJJaRax1feiE4VhfBZCQRtq6Pe1
Kkp1ea0vzJ5b8WtN7CfivsBbhHL5ZgQyGUX0X3FiEOt/jOLjAtpS+Z6Do5mHe9OvjaKDUix9iNCo
2GFVgPo9EbgqsCos3xOyskuSPXCY/7wCxMnf1iEkZ/w6DPhzTg80EDIQIMzbmOFBl0uSJOMEX93j
GTzWzewfVXE19M82NML4+vITSqllKnjs7bj3OIHmvPdxuZj2ruFkOmzd9ORjlEGn1x3MLWNyy0M5
A1v6VS1WkJiyNSnNcnO2dKN/md1WwDMZerraIJKGnNDwiMW2zGSOHNIhO2L/2tZuz4EegcAI11tp
5nWPXodAEL+tcDtrACk/TbmYc85GoPpiJIwFWwxyvO/kXoA65JbWMhyj/R6CjGuBehaQXtHV4Ltc
ZgLfXsKeWpDKMvpbDuIquV074/PdydEuY9cllmpvqRUNA0IZ1bu8zUMY4TULQhkSV0EmNPBgPAj+
rcesDtYxbi58JPkVrmT5Wb7ewpGcAygP3Wjvr7a6BfkliuRT9x4LSndilQHFMBqWwG2HohUYack8
OiWLrqEA7ptKGYFLoJwYJcO4wfmnt6DPVI6U98QXitLL58fJaSpb+uo3CYz6NUta2AAoBoD1aNO+
PglU4rYGxizeMoi5BTXLUgN55g6Qp3BeyGYmS/Nr/Pjle1PaJEnW8McYZ2Dg3oHr4s6c73pnkHvO
I3i4M3+dSsPQLHtzp2jMqsp2DSyhzzjv2ov57SsgyAa/rgeIzP1EqIw3QsVfyPFD6fWZjqIvXflu
cIjUOBXPx+2QydGEpoyMRwC9N9H6uY2/1hPCPb0nSbVuItOvdUaal8rANcXCRKgJotE5zDNSz1OO
AL5Omn9hhYMWsQtkOjyaUd293CnTeGa4GAPCfws1qlzwhnlEL5H8jObR8JiAECwxYLeFcq4w7OhX
sXg30fEgpLGSEbSImoyY9Aiy77TkQtgkLjbWSRtbaz6nVN1VCZKaQ22vmSKmqoh+onEXMk/x/AVK
zOQBnai1a7qvpw8riuUmgpLaRxkFE2OgPj7aetxLaiOnzvHcj0FoFQNKdXnBYVEhWK3KLITz0c6P
OZRjbdmIxem/Ts2XbkPH650czlcIhDzk/Vxh7XXgIHfPbjNte7V535OxC3UjyiDiJD3sxQ4A+TAl
HLkY+U98gwR+isK8hAgv5sUuTGonrqz8+3AmTxFir9mBycDpoLVWOAthOAischF3untcve9LS0Pa
4ufkGdMk5YdEv0wVRyYQF1wCB54GlLn/OzwVHYCFqjPkn49iRrBzc3BI3sOAZddnedx2r42ltAtH
WW9EtfLgUfSWMn+Nc2G4WEa2LCqfSKLluU4N4IWQ2oKtrii+iOVslvXRQLl56z6C8NbBHIC6yMPu
gr24hfIrnmynU7H4VSRMHMARzX8gjNgs+pTh+vxUWXUbNZ41VttNdLmAUrwGnU5KpHxESRU64J+3
SH/zrPGinV7eCclOxe4xPP4rYy6tVCntIZlxHt5Y61W9vIQwfFnsHRGGNIllXB7SYkr58zj8G554
do0/4slAQBr0I1+8lIc4S74o97m+TkTAejiztrgIthFH6Brke9Z/yFT/tFec5/N/qtYqtCE/c2/I
WW4pTkSo63qqx34vPL9h6bAxKlU00yABmlxKgvrPZL2bfAqoUbYI3bSJv8PzjKyyQGAQN3+7xf1/
FO+kEnKk7b3g9CTy0KI7v4IwpomEroaCZXcRHZpCk+iYsX3VfDLBbRtAE/g94fSbjIZm1Qxjru2O
/UINJvUc5MMfZnOFWoIyQWnM+t2485F3MMB4a2gqCxlxQ3cFmvStZNIT6A+J1578tC0Up1OsZafo
UHaFh8pb2+xfhZHUDr0IlP4lWuZwbVvylbmd89lh7yVMsgZxsEAtkflxh2yrYS0knTgA3xNNHXCZ
XgbLNOKr0H5WHSvpFeI4UNFmhpkePeU5Dp8h0wl4BqwQ0mKBzx7bPLnqPQ5UHp5EXXteAvCB+wIa
rRldCpEl4nsfSowXhfeIt1BkHz769sDGLoD0Zcmf8GkNQ9kUD6bNshzl0omVYLn3kuGdvMg7w22x
21313HDpRiL4IpsbCq9P5T68wWHDh8Bv/vT92hBwhRn1h28Uu6l58zBv3x+NJUX1JbCVwyMAz0Bs
ZlQHaPGWdrL/Q6he44nMXRkBa20nelqMZ6BkmBoYIzGmWKCH9UdoecNDYbIcK42d+gyIDNDw4Q9i
3o6++B6iS5KtVpX66pX6qrQegRMTefKotHUXhWMej8QL5RD0PZdNGJz66mwnYAosA7UZlNcaxkwW
qrATWjHHxvmGLYEudw+aHwNK43seDlyYIle1W05vF6FRs2xShcz8ltXEzgJqA3SJnVhO8r5xs9cl
j5YmW0AN35bscUYlsNp6qd2YNA0lh6q9Uvhr8CGx5g+xtiDbOxVjz2RoLz0IaJJxWp7dGOU1faJU
ZV4pABmENRRr10OsWHKVNAtzlsCnoxdL5eGwzqryXwLMenwy+HOe3bSEQ1dw/RioLcMMt28z+Xc/
PG8HBazQQu8JTFCMhRFk9aKWdeGdlJAhgkB1E6nXS1jXCtbORducTfNXrGyNk0IHgWGjq6mzSQ+M
hFvgTgcch4SW7Oc3BsxhMDKiN9SXO+Zj/udUPGE1kqmRIV/VYM1HF8jFIEgiPAVEJddVVd1XsRaP
OPFfNlRe5MV/MaLAU6MWOqQsP0rWaMGd0AFU0hTvcsTVlI7i9udmOxIKXtcY9GqDcByqWIYUi/Ee
SqXDN5PHhQOlrxN6pGCVgvlSA+acpsk7ABAGkQkEW6Ln/lXbCmGzkUm8OUhr2yvD+1IdIuJ9PE64
nllRbX6wkufS0bLRqmSFEcVwusZb0bwgpgspjXmsMmnXIbnBDiqRFyQajjuO6f5jzyjCpb97dJtj
wb8moUiZ30M9x9LLEzSBf++Mw+6UG7fpiDSH3LJ699x5KZ1B9B0PXcLcEGp9k+fd1PGkxkMQPSAC
mtMJD11Q7LV6kOJTp5DiWUg7waur+58eNE514djFhL+LnsIxG/73IG5DiDlwKfKhGd2NDORiKW7A
GjZ6bdX4Jtdi8oUKO9Dmu+CW0MEl7/fUfpqOl8R7JXOHUtl5zxwRml9Tooan12DNGHK9q8AOfyx1
Zr+Xcn/7Re1wlFIftvcuUcVR/gU8PRJnEt3qrCC5EQgLn51LpIR0INj7OG14jLzcGknvqbQl10op
/XOJco9smjl3jyM+TOlfoXYTyPLyQ91RxcXtj8v/mmzS22ndWKwxUthGE/5m5SIDYgarGooXsXCX
TwYVvM7M71ydR8DxseCqsmpx43zn4ah66WBibjVcHalCY9SLPtm91RrMgMtEsL+MPPdhMT/C6PE7
WBZ/OnIRhDzBzb7JUAsW4sd6Slk7+3egzUZsjCadDkUYDNf4NvI/i8B23r13O419iPYzqTgG9skH
+H/ha8W7vqBTMAbTbgO8/MZIAsXNSWi21BpTmX2R42bP/fN3U7COtCTdmp2sL2R6Eun1N8tO/lJF
pYpPRV+BiKtJis0pdW6iqFcY8FyxkDHOJCo6kD89dbTDTe/PugSyR/5JxNHRbsCuSigSYssTo7lx
q8DsznV62cboQl5OgKi1vV227Zg6+yJr9Ug8HxHBeuiPk8V3vPmmjFSK8HNn+RFIsXdm6gw0+AQr
QPTaK4+f7oc1J1sAD2VLNcMs9QLt1eM5mqqjdtFaXrtvrmju1lVcNz4UyDVLlGwp1g9xhRrgvdzU
AHhXK18k9PI8KwMazHTcqAnvyz+NPD+JgetgSe0iSAaxJVBTIZv739vgtxSBvX9AHy6fK+BQ9aPX
HGJ0VFQjdYmJesMIw9YqaHYr+13enVAXKsGhxRBPzvKMzNrP2IoMCo1NRw878fmJkRt4xbG3PDnm
iK4LCJbvY7CKUsmd/DSsVuLCx24sTGh0Pi/8Q8/YAyM/zrzazEXqlGN/cAZssnDz+iJu5j6c8CGx
IX9VEAqAIUPwfghz9/K5jpnX+p9jHigZ+DmueHeIHwiUz5bOyPYrWRtANah5Gqh29FvIm1BekVtk
Z5mhqaC1R2fX3SDE8t6ZChzsb23zvoo3syG/lV5Dm8pE4gIwY0ftFvFNKMMZLq0elcMlgCCIMvjD
s2e3rMzGfidIMU1EJ7/ejHt65Tpfzzgkgbu+iPAj3Hh7n4NgUvLuhXhyRvY0WIvn6yaOmIeCHorQ
AyzbEAZbihTuj52Zp71Jit7yx6ZoGj8le0mby2kLnx9UFGDrp2pR6gqjybavljuqNXGmG1Bcmf6z
4Ak1nUfOxgA6kgr8kKWelONo2lQ9V1imB1ErAqHsjBRPVPJWJXG1OZmE8avWQxG6PsN3cOyJ2mDb
ZbhYrbEib2X2doca52gA3NRvPOPrkpXZ13Ud1IRUr4fx0yt3hluEl/nh2sXcQzaJBxBVnIarI+8W
bRYjCWBWJcxTRLDHmvlGmP838I+Q7I/Lnz/4J8tCW2MbAaRCwkwR5/YMcoG7EuMdn7VqKr0HnyFL
e2WRG1h0DDSBXCx0yOL4F3PuVixV+ZMlWGmZNxGnMfnslNGtyX2oTHQh+9J3gx6I7hbaKZNeWYEe
yRzxCU96eM8V6HzNhAUygFnhU76CmgaJyieKGjg/WvEmdxxqXBbYxi+GLMz+/OSyIphAQ5rwsDsk
QWewfqAUwjQBKP2UhX3mM5QjnzFMvz1s6xvHySC1ezYzdyEtHWjIkRo1KGw9XDyB3HzOOEJ+aKOf
wrRfHoJXfWQN7Ra1RGMqm7TrNxaVNkOrEGpsIhVmEyY0+pYIOyMwlmK0ej8xW0issboFMdzmfIwF
EMFlJFz013o4vB1GUVFgkoagKUwQ2a8AgaXQhBoSIWMABKMYqoYC48XUkVVGlmpqjSZu2/aWDZjg
nrMGgp+bHHA05DYqtBnAfct6WdQfccO6Pmc5a8A1VkAFM5dW54Xsp23177aY6pW/4RaoB27hPtEo
uuVEaaZsQzkKp3smSlr2wZpvFXihgIN6B9sUoU7Q5dN8n0TlPi0/YtTUGQJORNfKfvl2sPHWyU3E
feujucIqBxpfn009OQGXX2w7OcF/FoqF0Ky7d/b1SU2wAr1nnCys2AlLHzvZ1WGl1zl6hkLts/Wy
um0EmMuIbp2+gPJS3K8nvVyQ2+iQ2Oky8BUetutJkkwhQQ+ei4/T4m0RolIavZk12dBq/v94rFbq
oa8O+8Hf7TehWn09Pw9C8itExUrxv5Q97fPE9y1QzpoVpSVyfiCwtllUmWX4oTbOZ6KDcV1t0g2f
OQTsOqAuWnWkE0Sqdm3Y3E4yHxcm4Esx5zkeUymEOyB9PeS5ezsjs4gkyZJMBAwHSTOZAnRq5BOK
rH29nNcaomv0o5l2YS9qy46CbOeVNQKOtDyrrwKm3vvxGC30ExsML/jlZOyV1yKB2Q1nJpvFE8Yn
+vob/hn7K2yl5Djra9Yxa1alU68G8lZJyiBeZdEIJmC00x9Tmj3w0Fq11WIWJ6FH7j4hBjo4Ptx4
MjiRbVyUKb7xJdbQMnO07jZMqIj4WufSqFYuLvBNSArdBxFn9YNmpX9jKfZDxeyRXEYqt4Y/MZKC
MbucwQGyDzN5Kw6fjLQvRvUpuBn/7y3U1mtoK1yAeHlMS1nTkOCI3FBg6KDx9wJP9rELF8kJFNof
uRP8R6PRQWdWV9dmiUN97/cp8zYtdkSsLgWkIytUYPPf8ppJbaZZszx6ejx+7p6hN20AHtmACj+k
qZJ3AmpZJiDAv4hY9gbkKNiSKoumCicCVvdw7bRVfm3DueL3VAt/H3JiZhIFubmzOzM9IUPUqg05
ZzPMlQIZ/QYn0WCZ5BAr9kggrSFOe69ADmK5amKg8DCO43QRX9fHWKQmt583r6ekiE098LeZOuWB
jaIRxornPkcy9dQzU43653QvnkwAmk3rwACx2LKWW5Gh4uHjbS2t+ZEmuyoUqr7OlWodTXmTPfyY
taVqNW7O8PhUfHnzGH3KwBEu8dlsGh2Omu1LFTy0AFcjg56hvcgGMoglrHZTrOmkcgymJME7DqrZ
ScRlNjxGTQRhf5FSKWMfFgKd8CpOXfu3KlaCb3oCgbnK0ieKa7mMPr8I4I0Wbi15YQMeZF1NFrQM
w3BSsT/FMDOmH+HpsxRL78A70JW5n6i3PyuC3Ju77Uy5M3pHytwL6N7nEUSfiJsKOtpOjYaww1lw
AGGTpYnkD9+5TvGDMWg7lBe5gBu7ivMLmjWr2qpEeeynwATjbfZN8v3IQ6ECR0UHsP2zgXbnSV2V
SQF61T8XLq96TfaoiNBBbxzQu/RzV6+MnUaH9lJjfkGyeT8ICm1xrbQzhkDiJSYktxLBDW1vSfBw
30Z/nJaBYmTYX3Dt7ZGY11vtZX/YMe1Zxm2Ln8k//HFfbGn1HJWK5caje0ULG4KS8Q8w9xZECP61
WVkEn0x42laJXzJvmPZ1F4IHTdT+J+RyxolXMB4UkcZi/lgQRZncRc7TYZEUKnpazvN7ZolY6Iak
mKyD8Daw5MDaZje/WP+nK4gIGSTsZ7PSxjY5qq2gD0vP7DJckArWSVyoGrCe2w74iwGutzoefyX4
ktvSPdHgjceDlJXXkdkSUkDZ9NbwuDUPBRjUG9skVO3cJL8EmUmhElYF9X4G/2Xq68z2PdD3klNi
wOo2cWqPyw08ziZn4sda4MByzprzb/qPKc8aeKrazVoR8fueuxX4NN11PKIZPZDn+QjHi4th0ENN
K/nx2cg0zfWF0sSFm3r6obacG0DQesNmOjp7lb+UVY/tzO18SFznoRsnrFclwUMwaWaLmyWR421g
rWvMG5JM4iybVLnJzm8shurpGD19hfFhUXRNT0y/59jRrWhodFm8dbBSFOsc3a3B/dW8lUhYvc9w
/fEN+J7bA1N/NI12mubzx3QSEL/11GG7v84ZJMWEJbYkTdquhFgQrurGTara/AMVBDZesv0GL9nB
MV+ac6mq2oTLl1DuuYp9PLi8Am4jZIsqHZxqL1juR3M8A/L+ivsyUyDd+XwLgTmo7o56jalJksEr
wvUZmk+E3ou0CLzddtVKUWLJ1mxYxUvn1wbkTwGJ4vFdDCXpxxxMJDj1Hfvho0TAOJby04vePxMd
AOSlPjuQ+CBzwOTPHTeZ6VpkOtp6spOrkePeI+KIVNCvSxOEUZBPquXpuT8bYrWwn31ABtCOgCvu
pjyy18S+PXRFnacyq158+Wc2DsA4e86XeweegoaqDMdo57psdI8k1sVR5U4NOMMoeWsnim0lFR6m
+PILeL/RqZyfQnDhKEBTRCd76oW2IQ1+3gXaioDKTjlYUXJICyXP+tk8FEPmjP02ACZ6nM/mfqJM
X8FH693MK23H+Z8/2BPNYxKLX1OL3nMrbNhGYO9ltN70rMJ3MkvCO2uzCj24IllMrSIeSqE4bih8
651cb3yhdUZ1KjLMj87t0GiVjkwLMszB1J+xmk6wqNMRSN07oALyAsVqVUEyaCgI0/tiil7fTo+z
e0g63tFymS9jjYyR/B10mRT/ywdchk3Se/1RFAKskMzOg887AICtAsGnqJ0a/Smpa4EuSF6IB4Cf
To2OUmABURCpMc0h3aUNcwRlwwRztjZdQuW3cruxHL3zIms/Z8xBXYGXH8qMKNNhunCInXklF/Ia
rPeUAQEyYTpFoZOWzC9vZLIMNBr5s18COx+3hPASFZwAhl9i1HMT07xVpgyEqZ4Exzk+Hpa616dE
2MubYAYt8XQg1jqWOSgYbLpHo8B1K9qGP/ETuPJXr3qAhZndyOSB79a5ku7zN+2GD/SwkdCpafyb
h23p0t0fsSRnl1joes82TkDeZWHTSYSYHjXqV8JVjkWmtOWOvm2ex0p/gfd2weh45YhrpSaregGJ
3zwspsywOKFHMwDX+m1SH7leIjZxQ4DrbuGrrdC1pQENoRFQkH/6+SrvKSkDr/YreCUBq6v1Jic4
Kksm4J6VHjRrdKbS3ELYuoHrImOvGqXaTjuviSp0ncSsSVEZVFBHifm3rX9OPpXXQNPvPd+ufdc2
ISjv5atTeijmUawJmKtYobr+OYMIbVdVtoA86ALObUF2+Wq2MTlglGmLNjQGN+zGDsXQp4tO01PZ
99AvZY3+L9zj0FAP8zDIcUEwONh9bJynb6BePpXThXkfhPbcmHVdSchXuiJ9P2aB6RhVLq0evsoK
Ak3GmYWo2STLyHZbsxvnKQ6hwdzGAe2+UsbuWKKs4cnmRkxJp73vPbbJXGMwkbTOwbxjNIpbPXv1
FK5P1ErhbiHHUJMo2WSI3jy7YkShuJ0/uaBwSezg97s+dWoiJIpT+8zc04ckonpkdgQZKBRDPy4+
x7Xbz0HLjukcDDk6FRN6rE0slINa2/tKPCGPsxYSUmGG2yptHwsv74z5yQhx3oIcQwOeYvVEXtmt
P6vTBIrsX8+euOFcc4D836KX/Aw8+5oP73wqlN7UpL4Fq/W3nPjrLTWIfhrVNAvmHix43dPgoWkh
BzaJ3p/xEvhN8IOr51ETxs3LFHBDZOJq8T4YYS9RUb1GUQEzBAWgK7KXTYIn+VhJZ47P+EW67IVO
hD5MWkueD6HdsN29OyFLs4FgkzBoepH746nIn8K2iJHYVr+xpvwFa+e+Zxx0ZpMkWdAG4SjJbRVb
sGMNpyehweTceo5ch2/eQtdFTth+flRWweN5po6eI6fvIfA2CT5Jr5q5A2blJjq/UL8l+y0Fk9Yf
v2UQ9DlMCUKtesyc2j0q3iR//4RGcxt0sYHuCtdfNVdYBvu7RE34mQnI1rNQW7ZvxK5XivXhWumB
1+UJ8L534hzr5HdLJgOZo0oGy8YLYSrUu1xpCKFnV6zf9JEB0/a/CXJSuOeyFHFEeuayofWm1Qwj
N7qVyWpL9k7lqVt5eSr/osP8W+VAvFLXU1cF3pZoy5rrDJU3u8aKbSgeAy6FSZLWtGBD1lR3W7pC
3L7eU97SWbrdUPRGxgatLZzC6J4dwhG/JpmdbrUTbprGYW4yLqziTILSNwtpFOfFzGBiUGUrDCP9
BKv6r/h+6v8wtf84t+bJERstempn5hxLpQT+47yPOSYt4JCC9JB1o6Ufw9+YuD4zdTVUYUOjBlqW
8W61B+fop50O+adxeK7DpIYfvcmvhFGMRo0/p+rUsUD3RQv+QojFLYSQfLDUHaGZVp2CnBTT3a+Q
7ESFJRr7MDTU1Y62mCHuaJwqGjTtIxbYWazam6yW2XUwSdESWtncyx8ceeR6I9ZhlRibgBp8M0yk
bHZxnMqy8mRj04lsGmqPDYpi3BQEOkherioQkApHnBTvrg8W4dhhuI9pOwUF1Fk/NPK+IQqkVhnk
/ooZU5Cc6X8kXaWVl1qT9PGJMdm8mHhGbuNJgdX2GzSwTMK7ikh5pRemhJjlXXglSRIlGD3ztCnh
UKIiX6z5aOZBqimTxqlaLvE5bOVaOrS5BS2Ytn5Pa/ohB8taq0Cpa90P2aj0iFD5Vx1gfZxUz0lG
LQhdaNG3qJukfwgeKesmGH6Ua2QtKN0eMs/ymLTmJUOnC+dghyd/pzAm7AP1Cvjf38jM+3E1LZwl
jwUXkdRxxm0Uhvp5DQZHo3IT87BC3jUlKfaBiM4J63puy/sReEdttbzHztw+BB7XxaLqkSCLnhez
M9YnIsaLmtTA5PO9txptnxQaWQjO+a36oYNlTOrc3aC58+cK5jorMhe/6jrOqcDTtkTJ6DTweeHB
1zYgnizQ0v3bd5dQT5FqZm4rIaiHyZttMlYVAuAcH0/xg+wjGc6cAMzyEnXY708T6Jc6ShhpZCz5
l/E+AgwisTdlZ1wuOAzGDinl9Smmf/SJuYa8SQIbGCT8SZE7VukyZzs32YzPzplGit4nvDDMDJfl
fUjEdxwkdSSvcQ9Se15nxjV6ZeF7V1WzIKl8x0hUTkK58JDtSKBgY4SoKj4kEflVEvdPCng79b0Q
QmwJHczPDgUzXHqnTQrlBLb3I5xyZQQjppsp+eQ/QolxYY2/WP7/pWHcVNPXp2beloTB9qM72Jh5
GRqEJxr2BCbTaW5zveR1rCEDm5PX4vpm4LcA6QYK+ePYEHAeh6Xztl5jiTQO+ip+x90s9/IqyjYP
hiYIlSoKsQ7duN/8aWbUyf8KVXRaRRWSIqbIDBeuds6suMiEqIMDGf+L35xwExQS8vpNcd3USUX4
eDkns0HYpC9ZSwQAJm3PLiYvr3Uuuj0fhyIxcnTEqAVxEZ4KiIL7FIdHF5LrDnDoMhm6KiSfVuF4
SoozWhVmP4O8P0vZ/kWP24E7wtC7ls5Z6HXJ5OqakpD/dGBcIUt/wjPAP50BoTE4kjdeb6VGsTsD
KAmQGOysUHnFlDD4Kk2p4ZtziOZSihEX5GrHUaAuzzwGaO5mJ5+irJx1639RIUTtKz1V4B6ggIv2
zm0PYrFvibkAXQuLScvHjltR4QHuzFCqY4oSoBZEmNDNnlGkjKieEukPyEy0l0JV8cfzhRdJCAFg
N4IOOjmlI6wmSvbQ6Covffa1ASUJLpUk8cTRR4XBj3P8qb39LJ+vhhbUREJTTcleWQCx17yQmdQE
JsHFA3xgRJfbdAw6zfTbrJUUxPzRGZHY2OS7lG70M9pUexWhXjRwXO30iOR6g81vQiQ7n7Y9luiP
QADdgTqiF86WZH8FFT54cZUi4SHCfhMNj71Rnp7nstFqH88h0yQryDe8XSeZ1/eG51j/78rBDmNQ
vFr81CAFy4K0VJnyQvuhdE3GAE4iA4Gg/o6Ff87WWFhWDBk8Udy0YQekKh8LgCSFYXyoekbCrcMI
CAWpo3e5UIqs61s+P7nFxUPekov4fVZC4ypiFstck7pMH1xAmd4Eqe7gcYywaOM2ZOod28hgAhni
dYOyAJzc+YuRnztkFhgKNOGOc1Gd6fq2qeLo3GDRjsln60A/3vHxqhNxR2swWE3kKHpIDUUCBdBA
td/t5t94kiiJGy8+eiiBDCGEUr4NjPRq24nox452+3uyHxDY2bUZR/YWhectn+ycJULPMmpPtyaW
szjYWR5JItrQFefKlHhUOnGkmtaFH8+HMGQLbbwh3ImlVOQ281747iScgK6Eq6vzDIjMNeT6AaGY
JnSNOFK1tj6gbELSAg9zzn/H87RmJ5sZFL5AhrUQJ12kKqKBOoMuLChO3VzUTb2ZQGpQ9CtB2FWL
zsYNHJ13QoM3mKS4vsI4lO93DJIe3rZ7rnHT9Hv5P5B2OifnK6ySDGrhfNi2MdV1f84t6b0RiB0V
vxdyhXjio7KIdArOT5dUoUS7bG0crYSL4NxN8Tvl7yz1bWivZKeDGIV6OPlsDuaYxOxJQXhd+kq0
gmiiLhT77stmG3bhe0jwF8w+TsFeJp/uUvYqAtRNl87K1UCnt5qbrpkmehGbdqJgwjZ7+ewva2Nw
WK0anUITqT2DDMcHJ2/jvcfKGs3BDbAANrrVg8DaBaLm9UcExCbVqyDUnXFuz/QqyYakPsgmB3X4
0lDrwXfOHImNQTledTMh5rA54rnmQ7IgedhnaRLaNzB4aKd1J/lrqhnQbNFbd00crx82qgB4swdR
fd/eYltmsjo4TSAIiCqXu1zEqyLhF/XD1MW01Y79VjiGPUcml1qAQuS8v6KH7LgqqehiXNY/bMat
OPFGBCcSjpp+lndZ6siSao433guDxYI+V0QrUXovaWwRG0LLJqxmZ1yKl3E2tJMJN/LDulrFhevC
v8hVpvQjalKTFoCOREPOxvmBdecVO3FroZLijA3+nv2tG4uQKEgvjmRmgcrFKGgGdYaJ/0XPiYI8
ku+3NdZ4HU7MgraNuShgN0vqk4NK19PsfZbN1neh53e85pTFMfIG8cJfy3fcTvdq+yxipsEHKXe1
J2wtcs7SyCC3fPEgxc0qUmCWVCiVQzY81C0iLgGX1/da/X1fYwnXv8WAnziO0Ee3GDeaHI0wRvAe
RJA5v0ETgZPBjq2ZzTj/uOQxo2zeqGGbb2B6FDa4l5KJjKeiUYuGFoHLriNbSw1DLCCQDa4biJBi
AkmpnmvyktFGmrRJ60B3yaG1TLXIdae1gNqNCdlORS9w2YXS+6hFaRiAF1OgmfgwVI3XVQuauWc9
2pqA3hEcDFqwHciJbRAsqqZCAiyxvuGCORaxYYnorLq1emRSVQd6en3yzlm8fOhten1QWNwoof+/
Iw6JN49C4sqgYlMjpQey2QGXu9LZPp0VwsYyr16pl4TKRiiqqKjwSI6SnNfksggooVBObah+WVOj
P0vHCvaWKiTy57cGHNbBEFG0/ayLUKvuJ9wGQNP0AY9OisBESKhg3o+OWn5/hWgP/DuCCf3MUnK5
2CD/mJI7TIVfwFF8ur8pQ/8SCX/Mv8dTpWUaFt+LCzzvt+0XUbvl3wezpcyfZKe2DNeaGTOCE2P1
AcwYpbttD8B9kplgFnc1JSr+W0NjWh8e40MX/Oi/fIkiegY0qox7Slj6MU4/F1UPBjovpnoWr5TB
eJ37eukp/g61UQ1v2FSUP+OjO10pxpK7nuD5p6QfnlJu8tY+cx2aNNUcQunQJahekg22I7e39MuN
pFS+/pJBqn5Q0pcKaTFbnfT6j85F0m+iwxZ6iuuj3AYBBNyF/iNT8Y3OkR/CdKCLHuv5VbRHEZT/
FglwcCYiVpcHLyFVO+toadoQ6h53yxWfJqG1cbaXHlCVc7Ih4oLKVQPd0QNakNk0TjCML6UiDtu4
KyCQ67rKlcjWPui9Ud3dkySWn8m5YSvnLoZGpMIy7BKoOSOAUsiLvwtsvb3mktMuFLTHy61TI11+
oPQgwjYP7l6bOlcosduZsC1rYZ47+8Q4t50ej+xwZsDsK+EXadfxERyv7dCFGeawDf+LAj1FEINb
Iw/Jv6/DPEC/HcxMvi239Xi2hvplTqNb/+n1Hwx3qwZ1XTxpmyjYga/1KRURT6IxVfZNDyW1sXte
mEJskGicfRCIx2VAtQvoHsu1DBCBSZw2BIp2xyjpM9T8csb7zZoBfAf0AAGJc7MaALadTzyXNJo5
on/fqzCQjoiODFCUx/ETtv9bJJpcSykD2cX2nIA+yBlflccOfzHTp0Y6WpIm5NKILQSsk18MRkLs
DSokLTpxM9I69ZzvZpmtgxYgSduiwmo7IWc+WwCb212DMVZ4d6rMlXR3IS2FuDMdZvT328k3OStm
besmB86503jda3nK2IMfdZm7S2joWkhPCHbZDXDkJSKLwo5nB1VT6prVQ7jN8IwMy7hwxG0Gj4Lp
btSh5NM5o5iDXFjLhqWuTJmt3ch3SpqqiwKAqldvrPk6+iC4a1aDsOGIBVFB7jr1epaztMLHQCeO
1d5JmJs+Ye+NA7FIFA5sT9LTjmdeyjY1vOMILrhreLp4rE0DH/zSF0wxixq+fVGBn03Ndkp8J1Vu
K/PIrMY3LcZ9fUkBjdVS7ZiLAzTjh8bOhAO8dbvgOT7YLBMWSAeQmqtln1YqR39SKvzz0tKrFa9X
9+8s7s6Fenx338ovgJggAXWqboCbcjpg4LaIw/FPcPLzFr8iF8RaplttiopH2f+84sb+uPZzVLaj
8w/o3cfYnkwyyRw5cV6j7tTENcvR70HGVqH3NVXHrqCwZ1OrHs+R26Rmbj8z+pOLSN4gQ8zpZcRK
CEHr7zeIYUYnjbo1qYvlBPmzZE49cSimOW/EMWeeM4Yoe9wzheTM8fvt6uAsKlj82tWoFmeoZE4L
04mYZE2SYgzts/7ITS2QVrjXAkCqRyiE8XBVlRF4su7+jVBGSbfTEAitu5Pqc11ex7fgxF0oK0k8
eiau7hhGTRRK8YERIsqVZNJMCtPr+FrfOhZw9L7R8wG7mN93pGKO++s2mPRyI53XsEcQXNsJjdj2
YzGZGCgkhxYCmtcSvNi2gDv0NZuLtfkNPK9nBeu761wWZqnfJI6kZWCBdSNSPJR3FMXWh3KBamr+
pIhFZr/gJVr9PrgYlxn1M56YDeeo8rNCxuDSsQGBVqY4tmNXPuTCje06cHMTBEyVs7FFUE/qbI5M
t58efjfWWm2Bs9Pa64y9XjjY+aiPs05crtDhhAOu8glRoWrySP7wXPooHEkzRHPBoQcILe9cjjFi
QapR3ECQZUSfjzDDJ59P4gd/eZcFY2LYkgIdMJwZf9+p+6yOJLCkWykpc0ArNtKweNsKXkFQ3RdU
pn6jtf8AoqDP5WyjKM0bN3E651nDsnHz2FQP4BKAvLfpb1EeltYcygfaXO7jBkJJ2tLIWxhWcQKH
PdlnWrwtVCjJn0rqGDI4QgcmECFx0rGsM5vSxfc/Gvqe3bpp7pSonJFCzfGxvhu3scPI6yTn6P5Z
1iVaK35uxumqC3Szru3nxJ7O4H2y3fKzd1ol8fgTjy1zGj4afBQqAAVnOc0b4QV/sg2GUQcPF780
dyrXhMjd9yV35LR/sUzUo7RcdZEBwDU9t0ysQOV/nx1rpCEABqyPdqDSRNREpAuYpx0967qiqsV6
J9TIqalG01U/wRiunOYvmkd27BhAM3s8mCdC4bODTfXpkwCpy0Tr9ccIp6bXz1on501x01Le4uZ6
bLgCBu91BgXT0T1jpJUgwKZZcYj7J92oZTBP/JDSErTubxdqzY9UIS4eepNYW9W2IBw7Oh0CV2iD
eel3vKIrgdFHRLdv5Ya1iqKcrib1ks6TciGmmCOpP3MccytgXH0JWVJPOQ9wP7VO/rl05OmnJgXz
zEUkkx/47z3AJ5iGpM/kp9MDvOCQUUsLn1n+BEfB17xuP/YEjwOEksWjP3TeCuiXMbX5uxcu9JpB
6gzsJ/WtKONCcWj/+2EoCvMnOBPOe8Sa8g7CH9w5h6GToLDfUVl2XxUJRF0UmzJ8MDcpuLt6et/O
uAWpOkbd3Ts8wHm/Bp+XWnzFQRBzwzeF10GGQgghuGAxvJwUNlkvLs6zxt9mczQWHEUY8B+9ApNN
f3tcV83mNn5wolACA2o69sreKrho+QnKBvA86i3yKpkr1MuXLdnO+kgJBUb1HVUjr+P59AGNLSBv
mdf9WQWIAQZo39QY+zf2eoT9Vg98AqssWawk48M3FtvXOE/KTV2S9FaMPrgfOsMHGzkl79KEyOv5
6dIW5MDGEKM/J5CWHQ6xS1+/WXv7fMGfmUNgmhXO+HpeZETAvJrGBnF4R7S6Bjl3WzdTEzs+M9pX
LEGP2tvX6gY4Iei3XmGOh4eEdiDUBdgVuM1SLPcd6YbHxQMDXMS+fYTjn9N0c03e2UA1IpiYl3QE
eqKNQhFd/gd/qmPzeDobZDHgc6x2SJYPwDBGG8Na5ZdcI3cr/QCkMyhOsuej6iHvegn+/V56MFNY
aF0JdoLF2/NtL0UL4LFvOq/zR+f1khRYsm7yBC0GaiBRfP5JUtmxbVZIBtHyyPcUY18BImqfJeP9
8Z10yUlldwjLSeTVukkDpyk4KL2kZTUR1Bs2AF+D2FJorfsSTI0xMU4hxveFPdLI+4wQ2y0Vk6HK
hDrMEK2TmHOxcvI8CMqTWl1WYIF2J/9eFo0xjZ6Q1Yd25BQ9bTJOhIE9M1h+6nTXQwECgSbiR59s
sUu0tJiu0cW/WoN3QzoQzT4eRaKwu2ufqZc7obyaAi5zvRRpr6AjFpdvUTwo3njS+8+2aMgfIzL6
tZfQYJrk04LxyGnHTu+4XDEiRzuLW5vsGvkOesLrT0RZ3RpJF3inOWsJZIjHMX7mYlHlXvEkzAyh
XkitFBY7+Ol9XR4nO5VDU/vigwbW5Krs0OxIdnqtwE/ERBpK2Hl7ehBiyig4uDR6RaB1e2eNITZ4
wGoxli56Pgy+39tySeDG08wo73RKkef7uT0kxQYlE07vEbHJDMzvQTC1lXbxUOZNqUd+18qZjivK
hT/ecPe+Z1W1FAPzTwqCfGziEdCpIE3AZFuibtQJ8yeHRgfnNassRQqYO4IC6jexUPecrHXmwo67
/3XaIWtSeE4D5gu0TYvm0gl0teHT4HlEg8042jm5dlnrvOroKWyVRTewuY0srqQH75XZbfIeTB0V
5lr6a/v+DwVUU0h197yFdVJ3bIZNctJz7IB8cJUT07ZxxPcIr9cLP1cEErvCCgaD4TmOo5AMIqyF
JCUDWIqqNFXV2od0/6dRkVd6h1Z725eDR8qTkIDlVVsJ5RkKanmaj4HlXrPeEvbbBRZpL3k7ax41
QTzcVGK6D6z1xqomjUjQeQjZhMVQA3m2/YIRw0gbVu3FAZWDFucqPRsc0jNTpSRUd+MrxQYE1tVE
/7GY/clcXyt6cuM3Pe18FmdriA+tl9uu19W1MUwZ3Fgvo5jmTqIeVZ18Bvk01dOff7dfj2tdjRrh
Mw8lMpUwmIB14ddxeEVrWoBBNY0Du6rvcbR0ckUxpsXDswhKR6knyBCiRqkAvE9HfDUqk96iESdr
/nBnDl/Xsp8DMg4ohwpaXMYr98vU4s7KUeOLLhJpgGmKe4ja4TitFfZjZ6WJZ2D5yZOTm+r4yICQ
aomxn9WAR4f42bCXPMJZj3fbIF4GNSLM5Kvm+LOZf2z9spIjjZh2+RPi4ixb3ekA4UmLVaivFN6s
you0sNsmgWwM7WS5yNemhMHJKP/gFhKHqFIJG70KgOOnUem2DZWwxf1ks+jRlcYR6GrN3iObKtei
pJ64YglL2RRH6/WkynBmZTaaLzQPUIozxMgVRQivdibSKECW03d8PKbdO8V1jYgScB4HzSCgUmuq
IwC9vXFh4qdRv072lgAtu21ruSHZudysxVX/yoI30zSXQdodPq8WX6wdyBqKdcyEm1yM3MK2tGoh
EoZf5/0KKN9Z20kUpqN5/xQ3tnsgLwl5qqqUJeP6YZRAW7J69GVNA/9OXDZDUFdJ9OAdGgk10V9G
kSutfnuL7CdmorKM2vgXPMS4C7Iln4yVQm7Ni39FkN6PUgHlqR5+9oG7wBzssrir/gdQ7KxGtT/g
MrEMWR7Xr6stPC+UneR2bGk2oUvCBQMQMLwFB3gUo9zLcrDiY6AaOrMNJ8HUFn15e6U+eCqT7Hu9
l0jEbQ0w66JX7HCWQLVmLr6Qk1uVAMNBpzJrnIjVIScrLwKHTi46Gt2ZqLACL1x4q4vGd9ExuFkG
jOJYQRp3YdB8IY7KT0ZPdtam7JeyQKYnyubmD918sCr1qZ6K/yV3nCxiS5GNPKAR2lC4m7sfbgVO
Eymb8TFnHC4rB/g1ANDY3zOzWCPJ8C+QMYuAaDBBaxpQl3+K9xFxcPeT2E0UQxjjtMYjQsVzRNU8
uTXrxD5rUxOpNjGZEyH5XvhlDpYBKobEFU/V3bX67HzvuKOjaRnHIrMruyC1O59x/gaFjwOzLYok
khjk/wji/2KYC9AE/fufrwt9Q1Li33X/czIk8oRx+5IGK87XALMJXXUlxgwxEjsDgfguksTs41mP
RkOOBwWCzAqh+eWOmpzBgnYQCUf2DSwb3IAxw2HLSQnwsdH+iYthfe0UBL8NZLprDcl/T3OwnRmT
6xWGSpU6COUZH3pR3AX6etNpzJtjOLsay68gjUkAlWsk6cDcP9IwIKnffuCWeyl/c9uGO496iQAF
PJNMzuQyG9T6xlxkJsfdO5BH45N99iwAexQ3ti7fMt2Q8W9HA2F5ODxsrcAKctn92JJIc9KuwlPY
hzrZecq0kEAkYq4rZoyiUxf3IG52owuE+Zvh+LZbTCKOGcMTKa15pkSbtP+bAASCvTy6Y6c36AMk
P6upMPTqG2h3RByu1vClahEb6xHXlINHrGByzNicyb9ueqS1DIvjny+XKq4400HIF7cxjep+rlCE
icM0QGM3xCfGu73FQPVn64gFqM66MCRAu/0sFgrYqPL6XZZeyXxGUatUVwMY+pscl6nmAwseu6Rf
gW5/7LnLXrKhjo5NWDk6FbxzBK4tzbPKc7ysNE/wWySlL2CTgAt9Gopg+om/0omvYq18bghi1qMb
2HY0+KbxArvxx6aVc1LfRizvhqUlsnmx61jTgJNJuprBxfuo07XeLFZGWopPhxK439GlOWQxfP8S
av6BAp0GuiheDahZYwH2WlV7Z35Re/iiIXGkPmnp9AV4Q6lKK3oEHIGm13YagHg7R8rYQzwoKKxb
4ry4/p6ehYrZZW5ugeFk91nxc0mHsopxGyCn/cuyEDEIBDbYDqecnMrF45F4KMO5VW41iK9OqQIM
ei5HBVQ5s1EL7HmJN+TDZRobm6t4FM8MbxpdyOKPfM+W/F/9Il9N2vM+y2GobYeQx64dZELjWWjH
Y7V3i9pSgMS5TqdcNm3TGAYYzvzisOgpDGYD1GWu20c9dL1NdtMsvk4hC3ACvr/+yCT1biy8NSep
o1WxoSvAFfXXxx7UUQVIPpW+2y1Oam+eDXAiQ6uYtUUpe/AHIXO0j/2/W1kyGD/lTHD4yyD2bf+c
qHa5bR6zxBV6wCjQbdjcGxmCZnIZHndRuiE3N12byKehaDQx5tloZw82XatRM5pIQNvTd60At+pT
0hdJXafoRLeeMWiFXjuDmKRggomC9MMs5p52tNBE++Vv7GkeefEMildNPNMmn5HUWsH0uT4RUl8b
ICSliiy3310W2mLIQEiQdwUxu3K3vKnmYcvwpNQnuXvwGZfXAZxLB2lLQdgoqXb9jTbXxw0QJ75J
3Ur/D/hUOKOM8s/WtwPdlk45LdzJiY04LxvqZ1P8zZr4tBxe7EJrUQsdDg9wjrx+Y/ci1r4ys6U3
YbyuwTSnLkfy7naxqUVlcogV8ho2YydpOGvatlRaujIosXQ0g31Vm6CAF/OODjgqkStO254jKh+l
eyG0E0J7NH5M0Kgg/kmLm7BwNGvCNdr10XpnJ+sCX744nwBuZM+JiAYp+x6Kr2tOxeF35JDtjTBT
3zWbWvZDQ5yVWn9v4rgYs+6ZpKnVov7VVR2cvKwjMsPVmSIp7tkfPm3yDxDxxI4JOCWniZPMbtMr
8d2KB9yU9TXPnVZtEG0uh5HbP8n1yiQE7xUclDcD4mXrZwnvDAtMIfWww2EDMMhd+47YFXHrqpjg
ahcCHE4vt4umsyWsrhG+MVnDT0JfpPcMoWrFB2eodvrMnHm2oG5DyWgUrHjfCE2YLZqJZX94arAM
e0UWb0rRJhqhaoi+XssEOiV3aBzewNz2QXAPYLWD89OKtGib5PBcDowa9llch4XlcJT7O9uRkK2k
JhbYslzvw1efTS99XbO8qXRKRQuZEcC2Pedb7yUEo/P53OTu0sgpfmf0uNb+bR5cirQ5HY5WO4NN
a0Uhln6dPx/LzeBHFEaM3MOzTzmgfwNaYloR9cFAwGIi74g/xvEW529lc2cIxEEWsXSZiDMByGa6
SiMAx45YjdhegeiYwOQfamzffZIpgAfEtWbIvlPMxooLjPvkapVL7CZ15nk8clUSoBXPbGsBCV0y
FuAcs0M9KEH32uNNprsyLVo1X0Lx+jDa4XJgf/w2NUqPwovMTQs4xGJLs10Ckkx5BLSFrxxTBmz/
WGReen8HfghXTXFrWpqhM1DUR45U6x/jGZcTYi4oi2zzxrzGsrk1RSWCcLqOkFJaLOUx7XpXJUZ/
vIcEsLHIKgxvkVJEMHd15GrmvH9h3Gqyz0D0dXjqcuBRf4+AbXvA9sy6KZTw+ib0P4K+Jgq6c0VK
vf2Ig/S04SgYKhNTGMSJKad5S3fgVT0SZeCVqRaI6fcwf4ZD/GuwbV9I5wMyyrHFxVUB1YYracSr
XON9FzZ5KF7gAtgOLyXhtsR8woZoM6iRTsg/OTaa+Hr3d3FVbDdf+KCOSWgJD9C0LWKT+kgeTfpJ
fQ4xVWnS0KRi+LMhK4iqViPx/1eyJ1VneJn9Bh9pQwJ2BoU9m8MwzPjdUK3tm2veh5xTUM8ZSC1t
rvCwANXfyHc6BUMre+eiUF14RwkBhnLPMZOBsKotE8wISpyioI5u4McIKqugiZUx6y1xsHzgrh3T
0mS3+B8R+AtyQirUl/TwTMx4U7Lb+qJKQ7eiCdK02weRs/OOULDQcy4Wj6HOVSVgXKHOKfBu6aSg
RjViOwncWI0JIQo1b+PMAbFWt0J/CL2jWWTvrjhZlJDoTTcWK/s9FtGD9h2uJHUU+UiMzBvQQwvb
z2DFt7tEb4MJZ/zAn0lFEeeYij/jIZ1xz0xYVWAFCP2sFAZWwEVjqtV/0949NJNY48CX/O8Fdgri
wq2AMX/3CBAuErrzlathymytG65B23ZEKK8YtPz8vRzFj3DsAtsZj4mJ1XUpPxHgZhaVRaEPUxlE
+4IBZTkwGO6Y2azE3wh0we89ru96c4+Rnoye7tPKlG0uui8Q9A3DC6sBJftWah7dH4eMuzpD7nva
ba9LRdRbmaj4fuAmRkIU4CG1XTbNQsTP2bLL8HFrsDdTRGlKz3DwPp1pTvCf5uaESTWr5eNYq+Jk
f7RtS/t1jeGB+2iIRkpMnjH1I6sngI7z9X4JTRVV+NbZ
`protect end_protected
