XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���P�$2��S9�+/uӕɼA�8�R���
p����f�+�<�ء��z�k��	�M�����B]q�"eG����\�BB�]a�e��Ƌ�+<8�P��]���]���Q�*�$@�~����W s7WB"~$�p� �|�c�� ��B7Ln�(<�pV�Q�'���x�������2#���N�k�FO��֡�����y�'MyE�K�T��V�����fw�9���h�:�n?6��[)T���|�dj�2��Ͻ��j�FH��)����D
����Ud|b��lw����4ª����m�
��ZIk��F0�g��7�7w�`�n���},_�������N+�l��)�-}���-Z��ɋMTK=�HE��Mf�Ej#5]d�3?hC�1�0�6&�#�H�91�X�[r�"C>�ͤM'Y�����l�?��2�����):����Ϭg�7�wY����z1E3g�H�	C|���@�N������[Y0�I���b������1�lt�Q�q�G�_�8�S&6�,�^�9��Mv%_�x�29*�bΨ0x��W{i.����@��:`=�����c�����D�R:������Zω�}�'bl�q�2��5!zq��sݩ��4-7�	��Gr��Ri�&RZ=#? �
p�Ѳ�-E����pQ�X��GsG̀�%D�h��#h�w���;��%r�I۩ڣ�s�e��J8�_W$����Ҁ�v��%��S,4��ٽ�I/��.�M6s�`���[�XlxVHYEB     400     210Sc#��{�a`�ЋIi�ͮ����c�y�&a	�>&h��z!<A֜���f+ʹ��' >	�V�Cu�����ٟ�*�Y4^�n��"�Ҡ�,.��{JY=�����/[T�Џ�`!X$ﺜT����k:�$G�
�m�"���A�s7�q���*#�2h���'ݢ�1<#��z��V%r{w��9�kwO��gW������QĢkTBB/�����������ͩR����TMl�%�Ӓg��U.��6x�d����7 �BE��)��ݨ<���s�Ӱ���:��2}o�g��W�".O\�H�qƯ�'��4�B"�M�z�Jj�iT��XC��;�t�p)�A����}�8.H�0����Ĵ�e�~���~���*c��@8ː�@�I�6OG�0(�Q�DT������v�Q ��:V8�r����(6��x8�ns�T��|���U ϳ��$��!� ��D�����?^��;d�{���;�� �[���x�I)t%ַ�k��(]����������XlxVHYEB     400     100�-������+���@�f)9�D�1,@�j���CF��ٔ��?�h�ʰ/Bc���{�q����?�r���{���������m-�?�0�`�|��S��֣B�)�X��מR|����j�9�T��X?��_.}��U���i;�C�]t7���bO����K����w�	8�/$�6$�I�~8.Z��||KN�uA3��H�-��ߍ�oS�
t�㜌�����g՝+��a�η�����i�f��-@d�yqXlxVHYEB     400     1f0^v�k�{�j�b)�+�L��,P�8E��18��+�9찾�w����\�%� ^g)6?�a%��C�B�u�Zl֕w�m95h��o��P�mG��H&���hYR��ۀs'�E������Nv^.�7%��C�g\����U0�̪ڳOr��t��G㒙}B�b���,ѫQ��!���+��A�w�}����w�K��Ҹ���T�&��펳��Q��0%������a%d�y)�q��\�9>�$_'2��vC)�� �D=�ѿ?�%��#��<ڜs�K�b0���.��A��s2�xVǛ���Y��G����8W��n$lî;�㏍훪N~�	�l��ۮ�'��K�Ա�x��� �� 3n�]�zgD��Az~E�Bn��5�����8󱁓F�L���!�)N��8K��1��y��W�H
�Ի6L3"�&E!L����:�,=�y
����\�ØSP�Ǿ�ځ7�A��;��nȘ���jMXlxVHYEB     400     230D�T���y��#0t��
����{��vƟH3�_3$���������2�����8 *����i����'�h����/�P��wc�즣��h����V�d�:
A<*����Ǒ}������`F=>�2
R���x��OIO�s'��b�Z#;�n �20)9��G
�����nro����*��\ڀr���l�^$G�0Z��:WD����{sXil�U�o�G�������$�£u��i����V�����~����Dy�K�bї��$.�S�?��f�^�b��#��k4g�^|S�[�O	y�j&u�q�����h��J��K5RM�\Lp��G����ѹ�xI�	u��jdl �p�LOp��E$X�-ʼ�u�K�V��5<ֿ���<7���%��h@ Pl��~��]�#z�"���� Tj�W^VPQL���M	�xk�x���`��[�^@�[�O��+i#ْU2TO#E�j.1��ꢞ��O��`� �,<�)��G������ĉ��������}3U��1�&�]XlxVHYEB     400     1a05_ج��Z��a�F�B��->����}hCЗn�p�8� .u.	%\�'Ys�bRye�'m�I9�'�L��)�{�h��FHB�R
@�q�\R�x��4�>2zh_@&CS�A+�A�@
7������ɥ�[G�ƫ�%�7n�p�c�lR�e6�;}��d��R}v�����/kN��1�)B�u:0?�N��x�q�)&=��o`�cҋ��p�[�9����'.j��	��G��lY1��tR�cl��ϢYq#
	XEY�p��a��S�?���s���_�`�-?)��s�@�_+`�dbI�Re
���j�]w�N����_n�(#�@�/�ț��mى�[b^�H�����m.z���\���` y�;���%�+>/G�Ԝ���a���i�%�B�_VXlxVHYEB     400     1a07�����
���N<T�!6mղ<\�e���wDJ����S��
#׈��n�����Q�%��j�H�Eh��{�f�z	�	������֨�p�y\���6hJ�����R'`.Z�Jh��Kq�-I��Dh$��_�����<���Lc�~fw��C!��/Zc;�F�h=%���7��'��Z��G�#U�+i�yw@/���(ByC`~jȐ���hf�[�=�VN�Z�k'�)N�Y���E'��M��X���90~�"N �����C���^�~�o���d/�NN.9�E��͎u�Vv�����W��V��ps�����NՎ�������~�`�>V���`�?L�n~̋�6g�#���5$1ـ�>D�y�8�� V�;�CAUΘ���=i�y�I�:�lg�
\���[��RM�(KȌ�XlxVHYEB     400     1d0#7��Qp�ʁ$����2��%.@��]���.B�V%n�z/��[��\J� ��]�<u��_�	o���Y;�� ��L�!��2L�6Y�
P�j��9�^gN��J����h�y�&�<�}B'�u�;B 0�YYN���ɍ�7�-�g@�;�
[|���j��Y��uzr�I���Q���۸ �v��{��S��=QH� !�AI�X�҆��-6�
_�`�"h�A�kD��1���c�(x��0U!��2�{�B��0P]F�v2�Ĳ4�����p�d�+deZ4�i�)������{վiݦ�2�RYy���b�L�eR�\M$�]����;�^R�˷q��Eݒ�f%����u[�cf!�l�S�c?Q?�E����PI_n��������J�1F�Y"���*���Տ��	��3e&�m������} �8�%���%��Q˦��XlxVHYEB     400     170z),�+�A�����������1t�"�{ox�²�U&�7[��&/�.I޾A>ݐ9Rv7#��̖�-gH�S)9�s��������.I��j��s�<��a8x����J�E��XX�܃�p�1E�8�O�fu��_>ku�8_w//��e��n�`��Gl����2�t�%��or�������ǁ�n��ܧ�����V���U"�Fp����,�^w.8�X�,�X�L\��8
�����ʄ�U��Z���K$1������� �U��3���2@���c9<i
��8�95% Xڡ���G��j��ߪ=r纉���&���X(�'���j���<[и�Ԁ{�*�����,l/B��XlxVHYEB     400     1c0�p�n&f~E�e�#�EF�xW<��%鏖7�9S��7x2Ǯ�>Ɗo�3�v��>��k����� [��7�2��˾���?�'5�t�21��"��
��ܾ�k��֠���ӹS(�)H`��3v��ܓ�d�N���<����OKh�a9�y�8���y��9z�5�70��Z??}��x�?NxKt�o������#�F��N��|-�����c��'b��8}���J����s�A^ &�]��K�ѡ�R�e7>ј �j���j���C��������I�-���4���eq�r�2�ب*��ȫ�|����ke��/�M��F>�$�,�&�����>a*0(B�1ř|�����+u&����H0��,�n`�T�8����UD+�]'��&����p�T��'i	�Q~\H�U���{x�����Ÿ-A�,y��XlxVHYEB     400     1a0�䵉\U{�L�^;	T��+y�S��D��P>�8�BA��R��W�B�e����a�$��:�
�|EQ�8p]܎f�:k�����/W�t�!:��.jZ6^���}�>�#�x��Ok�������K%��z4�Z	���J�������c�T����"/��ٮ�0�l��y$nx��()$
��Cs�3���d�U|���1UN��i�g��I����s1P�G��%��9�G��l����Mu@Y��"9<L�����=v?�<�müu|�v�]�����r\��K�q�����G��=[q�.h�����wެ(\F͋rs�j���ո��T��*���QZຬG�*�ٚ� ��8^�ު!I,1�t&`�F��qC@�#��ts��z�ɟ%��ӎ31xԷ`�1W�EXlxVHYEB     400     140��x��#�7��-gy��1�띠��WdH���ٺy��WY^�;R�a�ANѬhWڗ�i`�%�d�+�&��.�����?6�����BG	��A*tjR�P|�e���A���$�F�w�4TPWG�ʘ���cg�HDq���^e�u�'���D"0e����q�C���i��	8�����^
j��+���l�H�J��F�\��	��y�]~��s�2��`���q�:�|��RQ�=�<p��H��+��s�Q4�����<�>�]1J��`Ck�2X�[� 9�Bli/�`p� ���2�Gh�BC��^��n�Ƈ��j��XlxVHYEB     38a     180���̫��RG/X�t5��sb���@�QB"�.%M�L@6�ю�5��=?z�H�7�}�ڔ��Y0�Q7!�3�~�(,�Y]�2Q���ifY�v��JK/wl[/���*�S����,s
{7���'�K���˸"���+S�lZ�P3������t	}q}m^�C���%A���V@��5��x���G^�DLy.R �)p
ߘ�%�����hփ�1&��%�6�t�'��gv�_�$0`M�)�Au�ct$k�'n7q��P�!�0H��!3C�Z�q���C"�%<_���z<&�-Y�\si�qz���	���HC���6�D�M�Q�,3��P�Պ�R~A�%�JHb������:_���"ݦC�h��7�*$������