XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��.f86�����* �b&|ޜ<N|�'T�@��8W|<�f��*�Ʃ����oi������qҏGb��$�UQk�i;��xMB��>MUn��)f�B;'������z���j��F;�XJ�p�-&{���#F1��ёz�\�zc?=���+�?si-�-a�}^�2�d	i
 j��as���R}鉒�2ML�4�D��{:l�� !$�%��,_��Lz��u�Z�ď�V?c����d�� ��)^�[#���>��*I�h8KN�f��������7�Ɇ@y��;2Z���I�`���M݅��a� ��E�rT᷻%�K����b��K�5�6���8�aP�Z�f�P�ӵ�Y�ի��|QR�ߞU�g�5ċ��F�+,���$�;��ӖY�C1�s�\����R=-!9fo���Z#�(�&����+9�ߡa,|p���+=)z$t�U�j���7Bs�����x��������Z���qI�sz�h�Xeo��O�8Y�-���*Kwt�����!6�lz�q��E��9[uu
V	��e�s龫�x_Q���e�ihy�W�hp����:���L�Tݸ���\T�z���w���#'ξ$��77�� �����v�?��p(�-�բq4��"a$����-��@\��m�D�F#��k�qj�����|���8�}d!�G{S9����*	;Q�d���4�z����u-����Vz�M���J~���g�*�A�#<�1%���s�J6���CkD�UK��XlxVHYEB     400     1b0�{��5�B]��VD�2֚��ɿ©�Rǈ�S4����{8������x6E���io��|fC�)IH���;d�	�.�sZg|����=ܮ�H�n*Vֶ���&01yQ?�D�0��W0�}3�����*�ȫ��B? ��;��������q��ۧK�K�V;йz;������%d#v��r^\5�=������^ 9$�� �q�3�$x!�?�E���os�o�t��e��ަ�+��,¦-ղI�^/ �[R}�)$�祪uXG�D_��&�xo87�G�r�ӫjcT�Y���0�4�a��Tp�i���&&n3������� z=u�"v����t���K{nY'�B��}Y^��}�t;��c����^��=+���9Q
7�͸;T�e_��0m��Q���p�������񡥞"�[�7��w�킢e�XlxVHYEB     400     130M"���/_]��i��*�T�P/��^)�l�d?raKf�J�k �g��M��}�,t.�H��M��a#1�� �ӊCip�WT���aq�И
4$ZL=�v��8�ĭ����#ۛה�y�C��, h7�f8"��V�F��r�ڒ\/p�4%���P�w�%����'���(HǑ�O�04�J�!�?>9:�uԧ��F�0���Ic�Fc1xk���_7��%�O2�f��r1,�j�@(��_d_'�D�L�3T��}� �T��o��t/O��-��HWe)J�A�]��J�{"�ϙoQ�XlxVHYEB     400     120�U��yC;T�)C+������ק�Q��=J�-�ڶ���\	!�D�RR�e��"fi�,�M�[Ě��rܠ�6�ľ&C�J*�Ʋ�g��^}h+0��x}�R4���/���Qd���в��PB~ł/��/�mʋ�S�ɷ��q�σ�4๝
-��m�"�:���
��l^~�ntJn�q��ϳ"I�������7"3���L��(�E�s��)Pߔ`L �2y4Rі�WZf/�'����oQ��=�J�|������f7�`�J� Gki*���~�C�P�XlxVHYEB     400     170E��E�P0� �1�/��s�z�j���&�X'���#]�Y�G�Ƨsh8:��m�m�!�ɯ����!!���CsĮ�#�Y����A�W��am|�e��� d�ii1!l��8U�Oy+�LG�[|��+t`QBAd����F�_��,����e��;P���L���� ��t:�7��_k���w�K���rD�����h�E�h�H]�?44����U@���ŗqKl"q��O�any�b=��W�����@�y%��}6�j>mAʧ��(&�]��턢�Gs�Pb�tQgGm����%�]�O��ϒ?s5�ZMM5�缥��6#�~,�k�`Z9�\��:�}��m6�DH�T��"����R�XlxVHYEB     400     1c0�iszqR`>���6�>��yTv���V}��D����,�#V���W��i0E'�ɿ�>݋�#����G������U��ږ��9�~-��{j���'m�+���߮1D�|I��y���qҏ�I��������iw��X����8aD�V��C�o�q����\	6+R��X����( 	��{�U�
��������`�ml�ls��\���ܬ3i&ŏ砝����=2����, ��z�]����.5�a�Q�%�M:'�@B��R��i�)v�aRp�쎒.�*��c�GdI͓̽v�=wt$u��Lg�y����mЕ�xَ��Ru��IM,+>_d����d����T0�7�b���4���є*0炇���C �Ȉ�f�3�x��̎��G���U�K�zi�?o��>��ߨ:V���ڇ,+���8h�|^غXlxVHYEB     400     170R/��cm暣�%���)�	�*�ּ�l�Xl���ǅ��S9��GN>�!�����R�H��se2[zypX��a�Ϝ�2 �Y����e|Y钺v�n�	j�^]w�H���{�H0����\ȃY�r�^��1��?��H
��$K�x����g�B��I�������]�\�R��9`���|E�������As�V�l��*:��	]��f�a-˞�
��"pa{�x�A���'>ڳ�~�����,�hOk؟�����NO�5�D����;lM�@��H�YE�yb+�C�����?�#�T4�iK����=�˘��_��0K�eQsX	�qw���բӱ�!��+�Ie=$<�3|�	�±׀'��} XlxVHYEB      5a      50R��.<O?Q-��u$ !�>�(&
�EZ�,�JE���K6�1�n�oفD�o�P)v;��R��B��]��������m�X