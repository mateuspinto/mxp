`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14864)
`protect data_block
9t3xACmYOlT8qwqqymHK+AmCovZjvoeVJ/LjPcGP+I564Q3tTKvr2rEADH4qLIRW9m+BhV15Dglc
sISYUb68e0QKKKVPsilwu9VP6L5/nHlqW4vsioseRpCv7N+zc6afNmAccoG7422C6Fnxo5tMLhaq
L1MYL1G+iWEy7mVpAeosHrn3Uz6TMS//ayHfBABWycIqyAHytcsaH1CBNWes6bwIYKCfOwz5Pcqy
0RsWWmUOzGdCdscvjbBagsrErDP3lKhH0UsTMLC/5/ZBdIfeMgfuui4GrJeGp56e6/H/ykneOYQF
dI1bRdsvIS3MLhIX2Y6HKbFPZa+EvYqQg4XGA9D9Wv66wZtbPU75lZnr4wuLtlrmhANAiLHQDV5v
HJ+q1sbyRCjZd1w2CA/Y4OX6jTf454HUJ7CwtjmWbw0LS3LqqTF1r69bZ6O3bfT95bFor/WLSQoj
kOhhqHK4khriSfoRE4f3EPS8Z/Ai4dh16KWK63Fz8IA3y3KvKSWL6TR7rjI10OZ8bJm57VG1f/28
WNB2OBPA2/xVJQOLNLEghNSqRvIp6jGgTXkZ2WJYAHuoEJKHwWG1GHoVYcRpseU0oV2NK2CXOxFx
8GntDFB36vA/ewr+sdq4ZN6KuQ4bbVmNskyWR6leOBs2Z6A8ucOD9L+5SgOcLFrcp38jkgHCIonS
9Ol8evLUfD3ldEdr4ZI6N+PCkjQi152DzRNTUj4E1RkMQKSbcxOQ+iXdWQGllPgdAt3r+rk0ZdIG
LD54ytx0vJsm+6C+NI3nBnnKJEmtJZWeUhJWv8Df/aq0Y9l7dheWXyJW9RUuSNd9/jkJoqBOYdq6
YyLWMOeIjIY/bEsww86nbyqDVBN3x0vGlZeKYfwwQf5KegsCM3UKslNapL+GClvbRIgcGj48WoXa
jNvC4nR3gre4SrOTlJwmEyE6pI/4S9704UdruZFVLd+SquGmpcQX03kvDsqNa+knb6UNttGlLtZB
wjhjNLtELxGg8GxdNYGwASpDaJuO/IOssS+Sr2cgm/Hho2FA1xPJdSrvJpXvDdXxJyCGJUp4fB4Q
wTlGaV8X6YihDrO1A+acPsDsY2K/lkgu0GP1X7Vwlc8gNo6hSRJfIySbdXqHPL5DwrzGAhwMrmG6
2p3Ph4eh7pgiZAkLRZ7G8TkXw4pMmd8y5leplDeIwV6j92S4iA8PyNwIAvokL2h8uq/HI0koNW2u
oPgNLTwNZuD8tT/LwemYjAyKIMFunTDN9P620fYoFvm8gkAcLCh8EH59GsGcIoaxSP0pVEPioOtX
FJpwBzgJ2CbvLXpyAXatFH6CAN25ZomEXCwbQWC29h1BSrRDgN83fjUcWbVKz8gvEAVbBVagVvlR
gTj1ilNx8WZGCJcKI5nKlgjgCGyFYANapUsWrQQ0+60LN3KEtCFvAI0BR6E1+jSxEZSkA1cw9qId
F8ws7EJSXfd5QTKqB2HCmymatVi8KqGS+EJt9CzocrkJ1Hum/LC4sDWbZK6+B4i+hfggV6VbV86a
Gv692g/D6NN2Fo3lSvgc240OJPpfs1/N9hWEaOT4pV+mFKv4G3YMVEEgVSWyBi1yo1ptsJPOpDOd
I99yICDT99IL2gjG01lonPpfK4gAd12ZJvkkO8YiKdXhyWZnnKJuL9lN+xcwGHqIc1BmD4tfc1wc
Ymf2+cCO8UQgDZvvg9h/V3tzQsWAwPCp4+7FhbDzbn6wwt7ej4CPu4RyoSLHKR2BPh3yrc02lmAs
G+mmUymyvj1UNpaycIdeVKqS8UIQqO6AVRcyumQiq67uTahBK9qaqp5C8EoKqbd/1yI87dPz3Txm
DXkXgT2XI31JX7uV6DpOdSLYvXha0qGT907WPmSvkZu2ctwZ5ugJGUKuZT7Ar8BlIwJ4iQLGmuDg
IZaHs7zZVpWyo8W34VZmRs14OeP4gJW7GL1tpHGK/kb9leNWHyfFFtuToY/dM+E1zZNgYJNLBhwh
+6rQi+EE3RCQPogjEbcJwoHEAxv9smLSsjmZcWy6COiC5tP7dFeR25S8P34O11YAoRjylkjkGKfR
mLmu66PPZ0SiAFno0dpBsh/u1ZxTTzgA6ClUhT1uC26PSTTwdr2ke5/kiEjaLT6VMuDqTMRePs1x
gDd9v4gg/YaP/ysE02JaLyhxTI1PtsUFBxCdu2QK8xQc38Ellv4l8dIiKfqsJtKWesE8t8Zki69r
gmdaFfnnF9sXu8WV6B1ibiXUziiE8Q+sI50vPsuenTF+X9owBCF5x/Zqgdp62Una4d75M72/ZtDS
ddxoeDI2TZu37DNDb/nSFRd8MI+Tc1zKAFLbmIUxr2hXk7vNOyR47Y3jyzXy8VK9dNJuqzlqO/SW
SSN3sd0YV8WI7ccqgT+vrk8yeka84C4rmXMnjv9UPRqUVtr8yDrn6HucWz545oVG2pk6pS3wjxvv
brhlnVy7vD4FOtGj29bdghwVHmDT7VU/o2m9+QtA6Yx+/ea9u1iwDO6GanZyrtXiCt0C+IK+c8DC
YFVH/BLJ3ercjkcfDFy1hupdmjg0UK9C+bUm8X7l6frt3jc009H3n9E/gb71lGOJk/17QqfRkAVC
dgACwe11jZ2evR7pP5bCth8qc16OYddC4176/aikG0sQDZjw7FJanfcy2IjzTFaVZvZZevDYglc/
Dz5WPLFHWkxqs6c5BLsobQau56FT4ui6tpKFigT796yfKItjjvOTtvJVS+awhld/KANXhdFCNvnD
Xp9H3bwrSuyPEGfCMxftBJoDBzsM5I9fL8zmyNTBU0gEEtot14BuzmzkgzYDzyz/pW8DMarzfrVK
5ptMxfw5Fpj6RRuP0EdzexXTXhedLYXfp/9BhGNEOiy4z8/NJqiav/BTxpxFjzFUlOhNkfyCh+M4
2FrCgF2bWUVhBc8VkxskDqTBfvDj5ktKWb9WH7MPtiPUzIje+4XFeUe4QPCGcaq9Ym0gSKna7btO
o9TDzKav88LqpVczUMFMQmjSRXB0jkSHF5JXqcRwLMPltowCOvED+6WJGYct62RFVbrXlbQa6Lt7
/qf5Re4DLHQcKSW69oemngw3CHYEwhySWvDMWQK2I3Xlo95jM/w9YCzLhwIIv9U3aq0PmqUynhJ4
wnzH4NWknI0mnr0+bqw0uM+RuM53krN6tGXDb/wgrExoyavapyVc3csDpnzRFxdcvi2+L/Uwa9K8
/wIqqMn0kCAxV6pLEzjamdllbo6dUwNIUtP6bxM6/1z+Lg426BdJp6OF3EIHTpuZKLDMKoc+MTxE
GKVqA9f4eUUl3Y+Mw1Kvi3TovEef6E0rm9h9uqMfrWWiTja4BCrhUbRZIslqXGvrpbVKntc9hH7c
BcveSuXLMOeqiPDPCyjPurD9+at4Ux20gWxaRGcH29KPchYpJdJ6wRKmyMm2k9fafMz1WOoJaJki
dTDjLpjHskAPViV8TH9ZCtdjg9VPq14Wy8tKBU0mdv1GVAW+2uIFj1LPsFSm3owOEg68zQp9xjrI
L6qIZP1KfvIYbVxKUgrNe8CasCBZjKj8ix09vwrngnxogi6FM1p9Vd7ZnSypDj61rkHcLFt3gqpW
zra4LLiFvaHWDfQtxNXPm/ZDN+fOu1DwWNCvbL1GAUQ1VZvu89YfenVSzQvUu4wPXtpicnsi1LtZ
z6VzWqmm5L4NwtCYvfd7DAE9f3+KGssWM4Yn9YZ04kZkYIXoS1JXJJBw2sle3mXmhTRMCN4njc7i
KUS+O/TJAlUiSD+uprEhDyCCiQXzf61sEf7ApMXJW2YfniwnxUuV+DewvAlJmmXXHkdc7K8tWflp
oOL+fcamzlJb448s91qgqt9gX+BNu2hRcdR8aAITCV4zWMD82aBXsg/yqG5Lr1CrRHKOJmRXG9CM
QQ6gahDholOyLHWxmu8kGiPedJ/BD6D7r/L551qWdG95yqPAk37nbDCQCmL2Wqw2xuxl78mQv9J2
TFI/MLRM3AXrda2zAJtpCkUwiwuzfKrnsafCO5H24SqLuwms598MxxDmjRkrYYOchbu18+Z4uMuW
utRxeJyewHFcgITnnxZYbMSGiJw0hnDPZQTj9ttRufZIhY1oXYKL0uGo8W/s2WTzaXyDBruFI7TS
NnN+Dp4c2jpXON39JhQS9kO4J38P1SVKCnDX44Orgsib6KIzdMkgT6aGh+GP3fiwUzgtzlWKBLwz
C/VMYudc3EOzcQj3EY4CUQjViROkyVB8wV9iWgOsApI0BzPangGPGDOIRcRN6nA3Qe5KbFGsV8Gf
2fVSdEr9uo9HrNpKoXssjDMeu/msDQpvqKTcpggQQKozVIY/IsUxAGFoXOMc3IhmDu2hJTM1+UrZ
cNsLlYMtMj2UGNhnPplfGTP6vpWNgbn0JxWByOi2TbbpkiULj9S+EAV8SNICndjvLzcPZaCEfqTR
/UGqLcLIjr3ULZX0xVxHoyGeyYIui6KTgeNqNx+IsIvokALwec20nKxulMNVtkp9O+NKGj2FCmFY
3v7qbVmdpRmleiohQrdM12F0GV97Rz04TJXcalRW/AGHwG5jw4npNt8iOHZ+BdsaudNLcXsuKzLH
7r+5FUHrNaSNwttHocLS0BJkFF//4TnK1w/nugCwW/+W+xAt6hRCs433kmkPGoIjUTV85cePkFYU
uOK0XqvNEJD3Om+ZH95pN5X9xAUk6BeWzKFvTp0dlHPFlbrs12yRX8oXRAgL0ekvMwJW1l8VZzIq
P0KhIIsKTH+dFEIncinkKUncz3Nu8hq506yThkDkWjvP8OxYfxLXCwy9G0DskuiyPzY5hkJ9qzEQ
rr01le95pwNW7+cC3oiUfVTaF8HJBVhOICTFJ6U25pX+j6YIsiDvs437JjgTDBGUYF797CzUAdvr
nEjMVpWlNL8VKZRxb2Fshzm2bn2rAHR40Xqg6tRsMA+DR9Bpma3Wnha+cUn9LUdWc5WbzI1u/aqV
i40DAfHqnJKzSnGE4oiZWa+ffk8bBYXJS85QcsfWvV6vxd6/n6kqa01pQSLy5bnz967dnoenq6oi
/th9ilKB6PyBgr7l/bxqusOB2Xb4ZB4DoVAdetoaVhtlkJzUGQo0afjJpDt66TQ+OtNxpvq3+ViV
9sLOJ3ryVHAqiqVYWJ5S6Yo86w48tGIlx0dTS1x9J02PUp71bOaBCYi69nzJ00TN5e7CGVrB8VZO
xAJQmqv2CODKl33z4/rb9sdhok5OSEBk+CEouhdh1FK0wzOjJAItYhoo8Gbr9wxiVkuPPLn29DWS
xGV5HqrCKDDU5cKv5YG2mh+idewlHKITR3RYefoFOnI5qw7zwYs67V/yDXP+tKhqW5PHuIK3IIJJ
MKUCvF0Md3gS4ZhKJlwch8eLX1xwgsR/lBgTLgEceQJNu7q84Asp1PDlAKMQNydLL4bGv8tsNGmb
xpauuFh9ZkOOoiS2lUyjdy6zhlhdKPvoldrYVmkAxkA1BhmTdRPrvFHlRbGDqVWcZfKnLkfae08E
13dGb86ANXnGJgh3/P9ySA3/X10p7hNZQc7NC+h4HqzAzjSf/YeByeLVHkvvHxIcKX+MVv8rwg31
xNoTYnH9Ryxscl6v+n9m66gFyOInoXKLyW8MkuoyVBdaa/AL7jcipoJk6DiW8gHabKynYcqUBbAW
04mlFqXuAs8s5Qk9l3oGwYieD7FRMZKdZSvY8YsgX6bkIf+gIQnocpDscPJYXQ4t3NymrrPfJgKp
xGzdUljzIB9ORgGs66mrUtAbg8dKul/0Q5mQDOWe/LMJ/oT+gpZJKyH/B3D6gF6nOFS5tuc+NbEP
zMS+95757dYYoHidj0IhvNP7J9yEI4LWCBpE9+4manZaCxZQ+ety5zbHuNx+VOfpMr7wD4tQaD59
91T1VQ9Ma2a9VYBIPRG2xRJUF15PRNvW23f/t/kEtR0Ly9M0U3hvzMOblasuYLQnsFsGMwt21VGl
+NnB/mKQifgLOH4Yh8sGmMyY42dHUkxKohC5nTheXQMvkGzMIW4yNu3dUlWsNZvP8HixNSTWAhsa
gRELP42swujrrgHOhZOiEVtrZZm6T+zWKKyv2R+OK2v0jiRgcZl4wpFHsty24YptmUDWK2lhhwyp
d22W3J3cqtYRIilgUKhjWHfhuB85mfGYguzcA2qxdsbNwCMeaOjPAsx+20jiI4JFZvPOCKgsmkZF
pvEVk6k6Jusm1DmDepDlD0XP1s+dTi4j/wIKf9MNwkt7HBxfEEmUJ64+cTQzOG9KI7Z/TaZbPpWC
/so1kD+t7dGnEaWiFykmP041Kspn4BZsW6S3iaSBGUjv7e9dMOuaiujVVjcCZHZWdBDj5f2joo4d
kpvIUEHN2s3bEf0Sn3GVgRtI3+jbzILWIWNK7Hkr8IaXSWkFYW2in8xdDd+ZNRXhf4oSQuxzDwdn
CpLtkKjnUGU5Z3E8F0EdDFsZbD9zLldTp20jdVtfCcN/qzDuJXXuIRlRvwdDo2qWPVFistws6cqN
bGiakFyCKvZzmsZYoth+sy1x2BOH4JBibYp6QqrUlBVLfe1SV7DoMvGkm6m07s3sgjClSQx9nUpp
ek32XbQtYOw8FG64zPyHOoLuBjgxe+7TfCW8K6odUiRuzXybTJ1xKJH7LicJFwRbwSgysUKb8bFA
2GRTcN4CqgY6zAsUk6Dq0c5zwwERNNsEf9lxBpqZSfng2JnQsU5vCoaLVXN6vlVUGwrWutufA3rO
oQiCWyhL4Ayz0HUE+ZnL0ImXZEhHmFQ60Xk492CLC+yygjbJO6ft29dtRVwB2E5S2wiseUGlfwz4
Tq2t3dqdD6JZuYrUCh3wg50z+33yfIv1r/+a/qT6RbvWOIFhzaTPGD4mMVFLLMCkIuhs5qx2Lfhe
gRlhIWcw5oOmw2GHnlQcGh80pvzd3uLbPPcLlHL+P1WIRjsDhGGaxCmRxmmupfRUazT41GPYsY5D
4Ay80Ohnghy+2HXWsyndtiiyXU0tIWsLVj9zHTKZVak0RhxmnGuWcPImAotVtf04+6EojvNbYYc8
BpFB6nDaZEDN3AIfQKZL94aqAMUFMKItLeZp6NXGIzSYHgcVTlc3LMDY/lK5rcRvmBt87PJV0FcI
X4My23VdS//ImWCLKcAWD7Rq4MjEXfAht71SlUZUBnhgVUz/GNushBPdC60SQ0OMkXjzdiJ82A9r
ElmDll2bANFHdRHhZjsfoyjXZvufXSWGotmtjfQYZIHmiAD9fAeX/os2OHLTqGxjNATRykr95g2l
jk6LB3VnvneTkmIobJ03dChjB4tmI8QvgF1QLL+fA4+hD8a7AidFfs1U0oC92t9iow3MLaNps3Ar
neaNBw6ZDz3mSGAzgJ2Rr/NRRvkB1qUpc1GCzr6MF9xw98Y+bmhf1Ns/iQq2nvalBuO52z82r4Yw
1XSrW9AmqK4LbIBXboQBG8ekHhGBmE5VfGQXFbn83mbTISE4MCr9ioXiC5oHKiW0ww45GZ3a7PCM
uHw6ic/A4336eheJzZCEJSL5q4CYIDaoW4L/mGkEBHoS93NKEkLqpkcHvLzxReoTPSdYWZcLqcLb
I55O6NM/bP9EG7oqAhyZD2l/Ud1u42zuPA5m1SkEqM9kakQD3CSPoSjXnHC48EFxe8B6vG8n7q3p
k99G3PRuLFrPBr43W18wy1uwYmrwMCQzlLDYTbJXKoboVA8gCo62okupwyBSBoc1P5stVSjdEgft
OXWMVxEy4CzbjW5IP4+jFLzHnIBXE9pczq1K7xhhcqt4W76NZtmbdxk4s6cU/x/JMmEqmJkRuJy/
88bA+v+rM+MyKXd8d107XFFTPrkHSw6vAgBi0SSMzHKd4eA+tOYM7Q4gCYXuz6D+/6aa2dzvuBub
ygZ07OKPts+Vq9dPXDzsb1heOdJFHHqGj2TPq8Z1e3x+/5d9f9EKDFhdr7qdzxt5hE9xGw05PhQx
qTmAf3kDa4OTIX98e+9DSV1x+I/1Rq8+0fWFI42TIffLEGC6hPAJqMIGggBatDzikUgBl+SFncx0
gN7cWvjD1+aicYEDK5BMfEd7UFzf8g9SbGMIVAMNJOWdPbWQohMXWozrRuVHAYQndLbGNn6Wh4bF
GbwnWknb+0Lp37BUiKcw2oBTMhJ6mRJaHy9tBxDrlhwiErzfiTc8JlOnJ7gVxFa06PibwEZZ9lQ1
/xhqG1BZnjc2ztnq0PNNAG4nKHtlZ36bIIbRtHc4EBxs1j2K4ofVtkIfoi+YbrFzY9CVINpeiRr3
tt3QOdrI7ZrUrJhQ2p8Pbrb/K01j6k3lojCTJ8IZ3n0SsIsOiFmMslCU4dn+wH/iWgR3Skj5d3FO
TSVOKsUMBvUIabUakAzWjVIb2A97w2zC3kYaOXqrJa9rHpGyf9T2J1F2nlbnzYz6WwursNlmKnJ8
rDFEXVLzgb0Tzp8sa6bcdFpA/orre67WqS6D/nnWJIr2pCt79vd/bbln/TdYgY1EnVLUhzMGuKWQ
jzPR1rzzFmryCJuJjTnSE07sUVlRsugxIy+Lvjza4ga6ao8tEyNKkoxC1+1UVv/FF5aLsPH2SSMH
x9ipeQu7PwdFFGc+xcLoWbJ8Yzap7m7ZoFF/X+RRIN4kLdsuLVo8j7v/7j+iLN0xS8m+fZJ+n8rP
tSwddNiHtqkzvD8WLWeGFWiwvZ2rioUxUAPbNMi4LR6xZSwBE+cYseQpjzQVni2uW2nODWCHbs1q
p+Nc4zXBPSJFVpAJ6mD05f9IrvvAcdxrSDv+xN/2vKNLFEE9Zalqtp4+G8CarDLnMviyBGqmwrjp
HaYzXECKgEkz0AVSewR9Mfdyxr8pzSln2WKakvldR8a+65TIbAcQorSzXLf6oM0Mac6VW4574RHm
SQhbHUfYLf28VTbXVFFDAY6ApWW9mzeI0j2yv/1j8pWUp4E2th7xVwURjToElBy7R5/EYNuXqnOz
mMQnbRJio8FrWT0pe+SFuG+DS4pUae5TXeRKCpUvoUSHpa5zm9uPqkccsIrqiV1XZYsTiyAMNfbs
neJplBoUQ3yfYMMbzD/VN+7uFm11GHXuIlxgtlKsJpw+KZ2t7HIG8xInWDrlshGVbFu1nhu4ycNA
yUXHknNwXuGzpZTtOyi3T6WOp8NzOugMoFpShOkw9ckK9YVl2lCpS5IcAvHdLgJoptr7x4Ict5+Q
HK56sSi1ji2FDoB++MB1fwdRtyq6sHQpEhU0QWaPYymwnZ/PBnY5pH74IelAFfnWPphgOS2mwv93
i62rClsphqGV9QSTLzglsR94wJbwVNct68F1lcKtDRJde6DXTuNIVRT383bfWY1RraA00PyW6km7
2KdCNCJM52WMCVjlPZQq5V6IBQ+8joyngXJb1cmvGDj7I5QrOOKv6rRupP7ujY0FjCoZ4oZ+rJ6G
IlljB+hv3ELjG8CqvnioUhCZB/stndbLg5y8GobsYVC46YOCiiJqZUWkc97cMj6DScSvGP4xEtDZ
B63h+pfpC76VW7uezbMNXhOq6wHYLPZ8XHO3BzyHn7ZCUkc3DVUF9RinUiQvRH2xukSt/pjrGEUo
OmX7/OpwMTV0bY+hvlbL5l8Mnp4GnlXFaV15P+YDOhDWllRjR7xQmpXk/tLGuz8tnLcasEhTxx1J
BLr+stsFadDp6xmIc70km4I2QshqZoWnXC5ei3j0/G2UwDcpNyjaPpSQEFcgjjxJNigH7ioaAXOr
UqwP+3SMN8tcDdR7DnTPlh0wt86iHPWoBhuBvOc7f0bPCdmPW6AKgustDLog54NZX4ZeBKMeHUXj
GIZBLV2ikDDe2yU6uPeyfDIzfQiLzfnKOS5TTJQw0C7tZzGPXsmE+fdqFNwbm+UkmZ2jk8qcNB9W
vkRthiA8qvShJEg4wij7GDHY5N7Wljlprz77MW6NDki0o+E8bhJrsJ1wPiVkwkp8wPCL+aEjBaAc
xECBfCaEYY0KylOaw8f+j6LTD8kh4afafHPm2rxnjioIAzpIsy3r/+vFBFsLwLP4yyJz9HQqyMI/
ZT4RHp5dNm878l3t9T8MHOt9+NY4JJwSH7D/AgbeN4MqIk1QFHDIPshFvfzBGFrOQqNVN1doI4nv
JGxEMZBgtkfOKUMfP5QrFRpogmx9VxUiVU2zPfl+6OJTG+la9NXiXGbPxH5l6/+OMfDZgqf3jjb9
QqKbcDxdNp4xjR7k5IOMs759qQ8394IakT25lyOuxY7m9MTESTXkHMVSSZx1z0AaAluCYCdOaKdW
cAWOIXnNHHNFKeyeek3MBLDLAi9Odz3CRV5JUgdi9ND8+ddaju7HCVijid0YqMKlP80I6B7FY/aT
coOVMXoDKr8zLUS0RjUFRLT30BnjwBHTa6a/tbrjwRvuyJzT/YoRY6rVszAFi4nZ8mO6YLoqDlg7
fJBrPKxfy/AdIyTYS5JqLp1bsrXpeB1PxXeF8tgugE2XmCDzznrFqU8K8iuTI/gBwAsJ4awiq1wB
J0z7GheR1x/AcaUBmm0Gzu2DNKbDDW9LMFcxjzpuUwvaiC7MnJt16bcbiEQ5KaGXiPpdR0IfyvMp
oy7VYZ/Z+qfYp00Nhb32MTZ7anNZ0XvNrkUFoNNp/BuggrnXZui4i0tWJKl6ZXrncIZw+2Bd6KVT
3ZoVdOjlREiT/kUTPKiMAmd+TNc2VntnxTAd64D4xeww+sdVhpghUrCzaYYdLBFnp+NIOYMKYoSa
FwuTiqE8aDwK4cxpgDGxHcTei0SnHItnm8GyebQ6NfVK2co7oQsD2s2dhl2fhAMvMe9xJBZpk63m
n+buSaEI53bFidhkCgwXN6S6MAuOXWwYgMkCzEaKmOsMXnGNe66IsZTZQj84IJpfe422vofG6I+H
uUK+UirtfvZUFbkc97n6WtQeF5EcqSzQqClQOhJAeREfjFkLp5Z0MhcVMq6ROI+FHw9YwkKZ4aCP
TS9XTsNnchoPrxywKarl+QfHOdpDxUXS2Kk3QIy2r8AGWfGNfj894BWSNgSg6vyidyn+zqa+sqN3
BEYea0W2YMet1HZ7Gdf8C7xeyXtq3lFV5DEzCdXbHjNnvV6CKveh1HLOkMq5cr++sKpwP/QxZiKA
eE37Kf2i6z3xuggKnREprJU9Ge/lwWTt5tWcJKS+TwUyDCxxD31la7dMiTgXJBJHJGkUiKMvlODY
XUxXdSHwqaWfLdJawVw49fzIAZKdXMrvChI0FFcYQ4BjPO0b0Xzkdb9hpR6GOTO7QFf34TmhmLDK
5GyRGWa87Lv+qCEuIojkaoXyS4ZuW9LVl/48+wIjYrEjUl5fRw+kqbTGWKXME1Tz3hjJxgTbNcSd
1P3WzrHgCaWDW2e95sahzz3GVx6T7I85tFditL6RpoeG9fAVgkTuPWx3hzhnEhza5VZnBQK4QT4V
8qFeF4LF8n31srvz/uSF8T6DZYYYPYwHE5DcXalqFwnq4n0z7HWhJwmEDPIq/tYhi+CDEhUItBz+
bE007dqGEB52BCA0jNx7+YGQdYkVMzsNGdS3oJzsKgSh7zvTtflohrCBWZwlDvmv/4Ig/D8BK90y
GiDcicX7Aa52KaK0vzFfSnAHfqbBaQFNGUH4GVqAIBAVDnhgHI+GIUflgfooGq/liVWRY38XSb8Y
eKpuXqBLPmhpXQ3OO0J0DTuvPlJeXX1x/SkTOHxWjVlsFNPN9JGInKuUUFaOylJpB6xIhqMtdRAf
uLF/YgEjsrLvnseJiXApog91Q3vU+tyws6YYLMAR51XjcH02vhY/zbTxVWrk8QAw1AKHnhh+sDz+
WxQqAIHO6J5aCN4ygow9l+l98JESjBX+afD8NRevc84drZZ4jCtGK10F6DLGL0xZUmF0wWb1J+aW
sHTmOof39+05/6F4y3zLj2xvHE3ThtzWSGrmzTJPQ8CrKGLfcjhEY2+DKCqs8j5MOlhqzI70u7hA
UVMFBBuZ59RvDoHyjR7eEO1u5qvgCcnO6FGhMbzLSazWBh6LK6ZLx7cRlEVER77o3zoI+QCEdlN2
MGIBGpAXv8Ojhj0izz9m5Vo5oQBj75K9PIOjwsG/z1c7SYL1bqBaAs/UwNX7e7g5EDnOq16Haxkw
X8lo5D2RY7CuUvhEuZIy9oleEk2+nu6zWptv09Hy1NXlCZGXR7CQhlzXb7yJEZclA/CqbF1fhtbG
mf7GaOib4Xss2oOUt//ux8GrJx92dEN3SQyXfzRkww5XIWHktuIRC3XmUIMz9gqwacy9baDfCV2q
jzDI6yGf44gNXJNNJ/i10FAFamq3ROpmwhs3rwjobm5tomhAP6WP9nGP2x9od6sLFp40seCSQPu3
8iqWYkW5c2aY9xmHiVt0uCPhcI115Esr9fNyuiiU/X9bEX3IbEqOGU60/gi/3ThKSn59DRsIfwIT
uQifzyK1HySRnFriFR7dF1hjxXoC4cNUHbYeUoQJ5NUmrhcDoPJfrJFftDYosdhvq74PFU5NjTph
vmpgtUAvkfyBXwuq4WRet3QEoGfaBJfOhHyoHww/sj30kgKL1mefYhVhE50e1K73k/1Wx8bG+Anc
g7CbcAWgFBoZj1y7nhql4GTac5SX/bUmlN2JosRtxDTAzM2JdRh4e9FIoP1WAGJmIZJh9zuuYoI9
3eAtm/UrXEhjHPXh0T4YaYT7/6HUsL+1rR3Xxyhp9FS0ddhgufyLjfNeI8tm12GHFIGQaMFaU9g1
dAo85rtog2sAAPhe54f+2eqStR0OykbluLo1LMcf3tTbeHVNtFla46pquTkvd54GczIkt9GTG5gH
jUpvhYOZKA1gQZ+hyawcWvm9qUNiDKNZ5rxyQhaB/aSO4rRCU+GsN9O5RLjCNyHoFrRR2BH/17rn
KWYNHyXarrNHTtI8K0p9R7pAwyw+zN5I7fhFgiIqhRCG1jl2ig6wvg7YWxTmusVKNAhkF6HkloQN
c74aKD8shRnjnPQzMh6OZpx1P8SWHxqADoeK/GijHcUlsSWUJEF58rIFH7k8gGy5LvUzdArGH9cI
UfVlxsjNbhx2tZUL4usku2awnNqv7mbLIklM9baTHZa/k1kL8PBB6ePOYhRFj/LnvyE0wKj1N0AX
tOCTwn4GSY0p2bl0D1Jn31YKRnXSGL2O8GKTP8psXtulTNCMqrIQId14mKSc54fYn/qulHlBezKD
ivQwQcltQfVP/KTjFK9dgvMeHF6+IsmQK2JXtsFBFqzVj/hOoXW1wGUDm1SkoIxmOmkppKo6L0us
Nb2PQwdju3thtdQSsCtai/d9pDi44/1qHXG/jApHSpRBmX9ey26wqNMUMB8WbvVbli5opRkpaXXW
kIlDY4uA8I1HU0YXutT9UEcFVEJwYSeEvuqy1dEeaQzY22UTWgIEEymTl2a+SexQr+pFN5VMopit
muMHRZCbCdt3/4qGbRPRt2EsNEAIJb/HsyDeWcwIdQ/QAHAO6g4SxUvC3ptZx1LdgN3nGFY+465m
6UzHYFBPtrcjTTJ4w66qHNmjm6BkwjYPLKI+5OhpNBNyPlIcLvXDfOygHULtKCigaacQXl5juK5G
Mqu513LVo9FRj6507CpITjTVIncgFpmS9Ys6QviBB2UiERzpirMA4aLZjS+fPG9fr2lymCT341Uo
Nt+5ofiQ+PGmX3I80N8C6y27aWayV7aZ4n4hM+lhpmfA2BCEo3Z98E0mmphSCehuNXePxSZhSETL
7YT+5RcZDyLp5sCfNHc/vckgICnyU9icKbbQp2t6fSfiIaRaeLo3MkQjDPpHvhI/UkeUJsXaiQGV
hqmRMg3GVUpdaG9jvdoyY/RA5MJTT0TIiWQB1xGrVwSEO+0mukNd0v+lDv1RuQ9fDL4v+3sfzD1V
w/jMQah53fGwnvVPDj3JIP3Vwok7rR3FdNw5Nw/N5gjrU46jY35dFiw/EQc+KjaLp9LxZXeEtLqA
b3Vws34+eYEZOYo2oT2xbRoOF+f0MSZeupeDuLpmHz9Ln0xf9+pY0vpHG7AYQbOhLqqRyk9HPI3v
1eTXbJT9cJV0U3SsC8GSigX9RXbodbYFYJOqUHHmkK+FKPPDjsDbDhKNFrb3aF1A5+WbmJp+GXKY
RDyGaUYeMsejki7BUV3EOkWV0IAhol45VJ/yiH0xjD8SHd2/7MFhZwZ7+kNurUq7ST8Ukgj3PA3Q
IxPrsaxROpJl9oajiqkd1JLEHmjVFVVkZT7DFL1KbLHiMvuvqRtpFFuYvUHle1ziKoeazLvaXqYq
AfHllza/hchxEg9TqaC7Es1vv7qwIpmfefX+XlNoRB/fllp8zMdW/mybZkYJrKzLQQ+6xWumadZc
7nK+KcrxjR2tb7vQ6LX3gM/5wsrUm/ua7w/d94gr74yg6kIJbJT+1UFOvCKIxVdBYkS5thQFh5QO
N7Uu1qW1X+djMLNk8ZZAcHVwm78vJdAKRyQ4rp74dithF2VcM9Luab5eEPZmVy7B48r+XOs5Lhsi
mOLRWtfyofif+BbgBRIw6GMr1NdwNoM9Nc5G7nvtHFccGXfI3xvbugPxB6zKATFxC1zKD9i8RNs0
XEHEUUAQYuRgAZCn7jvgV0fu5Sk7LtVTdWSl7z05XbjndbL61ahXljeCjTl3WPFLoJQ+u/Xnd0z/
ASqnHw1DKhEXh6N4WcKM+wrsMn4aHQHH04nLkXNj4txAhVsbRfAFZyeevFHARKD8sgJdiGCk2zWp
lHvCDb4XOELkmZ8DCYFcy1OPYp3vT0vQKqpGvMUF6eDBHnL3oL1lAmXb8MnqK/BVuS5kwEygTqh0
mMbgSWX2j+46s9xXKNn4qCFqOmoMznwzzZkEQBf4NkuEbephTJXOQKNqeYmdo4jKKqWxb+ZHY1DZ
gJvQl8yCmvOq+dZHz0G8kVlEAQOlMI6GtkU2mWwoBwy0R3yw7B4X0SwZJy1e9q7Z+tSJ6IdnmMgE
+hA5Dbte77qIxD9oPupAAfrvK7DkKHGx3AA2SMs3CmLSR/OEMiV3tEecnUmVSWCxs1GYyNH2J0Dj
wrhCseMvLSE8IxPlxck6XyZLYjapeTsvpMlXeJmiu8ZcuHyOwosrvfNwPDFHv8KMUknSinSd046h
9nUPUz5rGkP9FudMfTa0ABvP5lRXeKITOzc+EZ1vpqz1WoVadR936N0JjTub+3weW26wKrWr8uAU
VsfSKUtIMLy2Fu6RbRrTG4dBERB55oD6TUToFrofPLy5gQo7KQdm9wUs0Di/jqeVWVSKYqcsirlZ
v+BtqX5c4riRuMxO4BcDRKyxkX2y/EXYRTA1GFWEQAo7WJwzhnpWj7YrdhuEONRdl4mb9BkP9pu5
ieAQitwfSSV85Vqw5ruPgdsQyh2Kp4RAZqrjDO3pVZQqZU9WtgQF77Zcx5FzLwcop4xxD/4w0s2O
q7mbMrF6xtme54dufDqsZkBSxTDieisSl73mHN9Q8iD7Vm+Q6H3qyXftkBQ56ZbOIPcSI2gjrbHH
Ifol1w5ZEAE9iGl6VVJPp9tnZZGfG6jJbZ1TvzzB0GMpxlPfHMPv3XOVLhWv2a+EduhYzMxk5BsT
H8/lyc1f/9+lNJEnF/NEpF6Z6fkjxNj9bHy21aC9i6zrLwoBpKlDOULcqMYU27wLtypvDzIUMlX4
OHLPlcNaTNjnCvoaFO4CESAOOnEBpf8NlJjTIlBptZ1U0dHuUWlwAqmkFNGTeu0Y4QnqEEpt2Ofz
FlDuPz+CrzM3/GP57Krfnc5jHSpYi8NUlVMXojUHzwWGfN9hSRH9EfeDThLg9Mk98gUrp6zejaKw
p7SDMSrW2w3Qwk7Jel5rhR2kh/GVtr/zGeCtANhF09r1pUOcQLUfym/SWdKHJmcjDwUkx0QQ0wqs
9/3mHptxVCK8dbMcBQkryw6m+iGcFG92fVL01gdh7qHq0VRQceSg3AJUx7VucycaxS1drswdO36O
TFAzf408jPfLR6yL0fhLn2ckBUJBeQpDG4bzONxD2ZSfJmeKbgaDpXktLubZG457Y+3IzyKUR+rz
gDwPyMEbajxyU0yzwCbUyWXbCdVxUldbwyXw/peweRmKB23acD3YlJMcMtXSzvAbFrsrPXvNyEWy
CnQh7zqWefMwrm3nHlUvVvZPmYlwt+ntVCdei1YGbcnwlBBVtRL4U9QSXkh6XnphUTLNcYYPAEY3
9m/u+goWhB7KT6NLxWtJp8/eQi3vK4x+KDZuXqLeafiV+zYcrmYJ1dUST5Zh4Snc032YVGcfsWVw
BzRzzthmSVJhHFeXU0Yq0XsXLM3Z1mlN0+qfSUkfOjtgypcWSY/9oE2th5X9eu+DS357O7j0VVyh
uM+Db0eIO9Z1o6YSHRLXUQHLmmnJMbde4n1FCjPXLXFVFPPG8H/F9Ib3s3HpZGiGLDYcSTgEPyZI
WBNcQKcIgx1jLtJRyhR7eKyUK5U5yDPEPaOt7bCjsbUU9mJFZN0IEJ4pkDLg8v0cJ3WYhstAQfYA
rXQPAmSF0YFPv+cVBbEjpBXEpbzniHbg94cVHasoQjsd0c5855sUrkgOkg54Oa59qWpsObDndDLy
fyFPsfYw1EiS3NpY9GpcsDi4y/v9rh8WyO2ToxQCsRaqmWU7gSKglQrs48HJzekCQGcO9Xt/grQe
3t1IqtsN+d8qgKTKF1xxXRrgdQt5uwjc4roqB1WVbby+QhANN7CQt5ag8n4BT+zMp+zk98JlZBw9
2FNZ6BgF/hH54bc7vWxLdT2gGuOrqipq/33zODw2zGELPZLL56VRf79Q+GMKQ8pMMDQgA7mznkoi
VZyb9cu6XZXTaP4LwkYgR/eKk/oROUqbA92SEJD3b9f0xUOgNkolu90jnWvnFWDM7QIzjr6z6qji
FbkaWrz/XZlhx+DkRGFvxQlT8IZl1W81cQXyTUb+nmvoRlRG++1E0//u6peGF8OeGX8nx4+66iO5
c5R1R6Znc8Egm/oen4+MI+v9Ae4Oswzo6NwTWGm1smR0ZxA6GvM0tEqGX8DJzrPYK3EpgbfgPTAQ
MO8NkGgrNGZmgO5OOYRMKesqP/f+o67A7tN/Qy3ksNY5gfoTu+habT1Y13QTvCkoOFwXh9zykSHg
QlL62sq2grsSzJ5SPJh9B6QmdigqRCNwz3aZQ64/LmEJFu7WFUCfrjNiiHDJS9hKftESplpWKwz+
Iebo+Zndw9UnzvDMVSJ8z+sBupLYt9IzuUcgNbwrNPs7e8C16ZkUzkBo83xaVvi65DD/afN+d5LL
rNeMJwrd+ZoQoL+37rwqWYcir3ewdGggrEQGH3trvBvrLZIIuWkVWS9xiEwxgIGmu4XiKNqlEDH9
dzMtVjDt1KEGuenaPlvksUc1Jphg4dBDlRiaR2Oe6XTELX4aJzzFGfU1TvbH3hhivH2/ZrBnFU66
JIIGoQQT0QEyANK9Ooci7iyFQvh3VP0S5e4LsaKlbiCpo+9PSWS7SGQN2SJf6PuIAo5MKRAUGWkx
V6Om1eVkcvbzdlv6CFX3CrCBWCm/MloJkiZX+yn2+o6ZQBbksmil6prdi42HPB2CVB9HtDWex+Gj
uw4qL2kNnAPUnistJk+euLtJrVy0gAY5jiI/zlrHqyuAOtyFRVT445Y5wKuThiXuT3j8Nz74PfNC
aGtFFKlvXyrY2NZ1oFPRhhW2Sr2GZuNiWCT+9N6wTBC+LPH0datIL4FvlemihReTC+KdDdqz3L+a
tVHCmf2d0mwvAgNmxjnLUwYMaFwUqIrun84n3Mccy2wKbIgxJ9BPxzn3LU9Zfc01n98/LCkRbSnP
eAK/spPxQhtKIz8dopRS6aT5+TZbAY4xcJAyHUZDaN+TO4S+oIJmglwOcJUIoE/e6T+3zd1rBFRM
ONyTYD+RH/9mYfPxFVMKUR71DYviGX5WJ0PTMhQyeJuQ+Rq0+FHsMIcB2OoKShfA6ykKNyKGXZ3f
/wwVj+LHa8jmf4M8QzUkFFAjl1kBM46UbGW35S47Yf5ds5TsdpkuwVnBk209hyVn99+T4Z9m+WQU
K3rm31Xsi4D+UMWfPa6on/+Nn8I8eTz78HvlyY2FaZsHkqPFtkDlkbAI/GYZGQAOa6zBSfB+TB4G
VGGEr3hTg/6wyhxeckPsj20nsHhdFG8iPATIkO3XKpjL8GGGyruzwW+BBrStFVeSKztZED3lA6OC
NS28KkKBx9bZ8kzurNzTdI6s/+GeveBfLrcvvcZWg09IItcvTed82V/g3uC2MHp74A7TdSNo20c9
LQ1bLiK37u/5MhUmlL191JfaEwGpaixiGG8UGKuDibAmXw9vqs74e5KtiReNQ4nxo1JeTRRDN3Qs
DM13V3K2XQjsZVOU5E0mdHSNtfSYiSbi9zmIdOS7BiH1klVJ6tXSWwGb7sGROIeXxcgTfvrQdVRY
9oDfOTcVRhcKnx+txannZpiqg9NRstaPEQ4rikbU4Fep6O+DCDdhV5L3LpmD6aFeEBVH1nJEmiW9
iC3zdiilcuUveYPbbMB57001Eft/JB/peTS1yRaOubFKoSCVCMzLvXkHhotVt/MmUrmFBIQemN+P
roxJxBrpP1p6thjV6nx/EyzJVzwcHPUiezIM123+80IbPRPVdU/kea0xy8MoP6mlE5qoNB2RKquU
oNR+xeBZZ66SNZZ1VIx54F9z5orvdNg0ff25TwNLf5bk0Zo6oujqe/0w+k8N8kChNd+dq04lbqtk
+BUZoOmm4vMQ1FcoqisnFeJOANIjZD1BfCbWGxjx9eTnclo2iK/hMX6A5kGLaQUB+AnNqVW27tUr
rQXu+032WTajGhbrtIAcNPKpAC6frqwB+eS6MfsitR/0BbgQtV7CEorKCqZAnT2ZT/iPOOggDH9t
R4Tx4CJikOyNINgH7J992+7tpESQPRlIZxc/GQC/j54GHggXiMTenfmWuQVAfjDQOMV1el2T90jj
ChdBbnZ3UC2q+7tHrRyOfr+J8cQdiNrZnWB5qufdxNaoq3xVjcd2bwlgK891DDmbVi0e4yxTPRwA
LGSdKWIRm9cR2+UwbSxfcraqaSnJh7NyJLIfvZW3ZiZ4wAbrKHYj19lNkA2plLvSB/I/8MK+SDxa
BLuxsud7k4kLC1zAl//cONLxcv39eR4EGqjmDCyO+WVKSV907paNMMbzuhSQQV0Te8nObrd2kYl9
HHSgfuS095CdLFtsFvBpMKwi5PgkGwM4+HP+m78Gq16yC/TKf8R4HcmRITkG0d0TDg5mgGKWt9GF
BMATXQY5Y32i+qxiQ3ErpePsYIQ8TTXy5ubfpm1xS2Yp88wr1NVbSQyRLEGnSfBqjCg1rT0ujsGu
CF6fmqYymN0TtlN1HzrslZQUlX1lkYm8zUgFSLqVjz6cEXfScsRsDVVIO2D5u8wXorh/Q7nJl61Q
NhAnVJa9v9oSyPhN4U5VzT8pS0OZKZsd80asZ2cajHJT5rX/11XxzmQqZYy/jz2kXS3EgpgZUFuG
Mme7eY+NO2jn1Wo3Fg7u2Ovfoi+2IAhiMiTmWEB4NJTJVJ1pkE1AJ9K8H+pEWmKQX9StUZKO6r5G
ZKOTNR18Q3D/9Z0xEWtf96UJy101UtK/4LBZPhQwOA158RWcM6PfVOSQRk3oPlUeR5KPNSdVUP4I
4bp7PWk8KLxFW/2as31KL7X5Lbhk2aEFLmhzniwUd8SZgr2PCNkkUKHzmFH/RVu0Jed/X+WaiBDf
d9pzH6jYZbNTRqoZQehHqf2yNKSFfra0ZP4ae//DP0ypF391Rwqx0WKoVwRhnDYGuyiN/XbhbbYG
HhRs9mxBK2D7d692V/1NNAU2XKeKiMe7/msSNTgAOfMJoNN/MkKr6MyP/YZl7qST41JhS/8FVc4D
np5yMZ3CMupduGU8F6KYrzO8iPoh97fBL7OuhHUhBG/Ata7szjzESq4oA7x6Htcp57s8+9gcNYD2
9i97t8FB/iNkX9oEPchpqy3iA2MHruqkkgh9R0n6yTZtFTq10Tbdp0Y5ZT4=
`protect end_protected
