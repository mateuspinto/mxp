`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6256)
`protect data_block
FqH6wYbyZjhSzkXn6QoQO3RnKZ6+saA74Rs70naXT4IbnbSsY88MXgl/Ty5Ko3CyFpch35bvOcHw
lKpAebngHKv71QDjsG3zOxEVxacnr+fs1MOhDWud44uZnBFsWpJez7647fRrvVSZLpyfSquNQWsd
ZxrRt2sfU522v8+7SbA8dDIy3EMEQwOtDKQDVJdbYUfi3warBzuEOpz6H6cHOf6FP0fl0ofbD5ls
BbZWW050HR3lQFDYCc2BCOsmKB9pDoCmLfD/wzWNl675PoGeuumEqoQvV5lj6v/OYCIsGUyLJ4IW
ZaQUbX9mkoO5fXMCmkB9UAMvhjfF6SrHENFQr95Be7pwJ1C6yDpLzBKaSh9d6NqKcE5WXY2hh66J
EhDcHi6Q3ZmY1Y2EAiQ8yeSbGKaAc93MC+OPMdWmKY5s1x7v7J2Zqi7nV+qcuI3n8oDmIkEFp9pA
xRggu+glNjjWohjgmDk/rwyZaHC/Cvu5Eb2+BPXo+PhP3CjhoVG0f9s0FhgCLHiodbTXHEzo6a7x
1cWtI+pTMyEPEn/U+mTQmU28BsNlXZivRHnZEeRl30YMuRB0njvTypXZdXDao1GKCQvj8SL1c7Se
M/we+t0XFyF1lUkZlpoKI0OoUTx4kp/qxEzHzifbCHfJDTBR+wE71DPJNl5kkD6KohMeLz1ffOEE
cN6aSAVUAlU/N7tJQkO+BBZ4zydzT1nQC+Pdon2zTcfegGoOeJatLO2Hz2wtgHuUSYuD7wIC2fn3
t+ZxY3eP8sJ/d4UrLcvbA328vYZznl+pnKA2/kSFXadvcv+kLQRhDiF3BHp2r7F30OG5goP/DG9E
SQsmR8UlH1qwYmKt6toK3A0o4gjsPtQ/akVfl8PYPG1IaQb47491Y5eiuJmBERF96QokxdOLIPFF
0UvpvB7lbQbKZmcnlJ2tAUklGM7EKREczXLNsrtvdGHwEMcW2e+7vM8bPT9ejM0s7DIGkR7lhUqU
pzDfmmQh9bxkYo1ijbV7eFHmPptXtL+2VXL34gIXCqaYtD17cykYHM2CqiUfwiFlXfVekh3fhYmp
wGhWVpVEuKHvp7qSoRAa1HaQFPL7wqrnbnfT+KMhzA5UF3tCY5EruTpEKBX0my9x4TRYOoNkfkPL
9G454AfHx0xEhsUVy43Sgn7BBgg3581kLQs8tq5AOUG3ZumtlsIwthlGNZ1yIZTM84mHOz1ILkRe
0Zm7OKiP3S16fwoi9h6MKpbB5oocSg+EHx97njCQIU/X+7Obzk7KQIeDA+rtvhSwsRdXUmoLxunS
E6rgzLt53s2IY6koVbTCtLsvmhJ8s5hHqBmiJvZAbl5fyNRnqeAhrCLP6E8R/y3JQlLOZEZel6l0
4bOm6IzB6tu9xgfMuHfOzAC/0mEoMCROE50hieJB2RqKjihtirB2P0/hY33wIqVptjGiaslEtBcK
2EGQ3fYVmZOwWa04354VT3BngwsokjXfjTwGXtjnIs4NYYJTT67u8IukMtxQz26JHMaNvbyJlKlR
TUU1O1shS2aBwEjOrP8PNMeShT8hYlEJOdBrl4CL5SQ+4A5g06Sv3E2XbBdNtq1CMvTRnHmsECZc
Xr9wgZWZHfosM+9MJIYre/+LunA8/CiUAfR7ilDV4SjAIaqS0enlw4UoaRNtlmU+0bzHEpU7n3v4
6rfWGC89Py9a12hguCbKJ6G2Wtr3ZA1rMHPt/izqqWBmoPTCm7g0pkuSoY8/lBz4comgRNZAvOe7
gyyMBWHsIkA7vR8foSWle3ZUFY2cQJ2cMfKDHheq+rtIQRmVYH0em+Hk5DSiNuId3bZyFEBfREkq
Xam/NOcr3hvj4FNtZ92fF54QSBuL+2vK8bkUA3VamLvGi29IDt4h8/5m3yIKBuetOxAHsEJA5sl5
zMFcA0rGkuual0O94HL7Gtsvr6Un/hLs6EbXBF+P3yndG+OMQbRT/NMOqfg9TaBHKoDS8eJmgPoN
v9478vy5uPD8kSyaaWeBovApI3TybGeVdvRhqvMZ1j1uCzoAB9JeavC1PLwTVB3JFDHDTC1tghQV
MOFSosPBAwhncRRg379TcibmIBcQDoetWa6VRhX9yHBB4p/lFJ/4JESQMMEB5SnntGnWslOBN2hS
TYkbVObDcUgqU1T3sC3fGjTaYcUMzIGHG31nwJMEUwL0AXmDjEiZKRYpNT077g2Mrdprt85R5HYT
YXiOl0h3RV5rT+Yx0AblyJMrhAEShjaUWe88UWT3ITO3pAi69Bk/SzySPcfvcliV1FdBA5Lpn8G0
MpJU284vBFML/cQJKXNv3qtGnp3grlkXBlXJO2FzOZp1vER2AB51JKSKUknknMeTXwOBnrqnlJBx
uAYBPOUCKnmKDqVTNp8BtNw6ybgoa+ZMg3GxC3Z60I/zfob10Mob1ZOLwav1mbPgqClTvd3J0GiH
nr6SN92j2TT8CiLuvLSVn2SEpcCStAK9PheF13KoPLRfJ0+hQRKx9rHfcU0Rt3VYPTWR6HvwQ0YX
939bMbILjyjGkZEUinOcidIqeD5VoZN2dApWHCEk3/zjRPfQ8hLcFXkunHZMUcPTwvHjWSQrVNeX
AvqnVVZD5KtajYnsIfOxmTxC/CnC+A87/nUKKd5nD+PF29XvjBAvvwpSqiTbR4OMLiWbhUKvfh5s
QLDd7E1bkxsN6HAp/867I7uwCXKFVqYZysReN5Ho+t+tLaD0/x0ndl6dVEYZ/w/MPKFLRwi2Lpvo
jDbEcO2wO37AbUgYMcoxUX4JZNjnnEuo2x/GZUSLbIck1IgvMOPs1ZiWaKXrckmn7OJvqsG4s6T+
c8uvtXQN+HjFE8MXgHqzW+yON3DzRoEqHjGaZdiyM8SXguKO87oiUSdeaupWl2ubvWb4MN3TLygS
gFxh7Sk/nOrjS7V54MraWBjn9qwC9Yb9FlEjirEUO/I2ADxiru+ww43B4dCltUtIj2qUHNSUnupK
wRlXya576/RjlVoj8insCPd3CZEHmXASX8zXFli9s9Qw2LdHspif6DFPp2b5oMttPxgyVIAyfEIM
GIU20Idnv3qwV4OgiE/uvNJAP1dvMTvi8sUHkB0UsXNJsRMmbEyE3Hjy2yFeFy0MhI2H6WVLPSrJ
obRDjlHl+JCPZRYhW6+T+MUKXkQ/oCRCV49t7QnrPmuQ20YkJMZlxaqRj+RL32y0ZH4H2UW3gVVC
EJ85VDuKmgry4VFLly4sE6Qr9W2jg+j0muhOcAenB90cffTkaZuZGHSAt8kCbKBXPzTzq1soZY+7
tI9VUth3HVxriiqajabTrGGFTCC9vGnyxiv2/mzjEtutpzRHP0nAsJ4XRrUhfoKNryxYy1nOpsWR
wn0sjvehJ022kt+qw6y5tVzofaBsu5nc29DawEwy9jdv5qXUlGDLJLebr42LvXR9AAdSWPbd5RVj
OJ+sHfBP/oHDRNUaWM199Kwd0h8aNOIYyMdrySDFMzonly8yCKeSb+y2gdKv9vqXfvC+dm2Uxj5q
zELq/HioqzgKeJxIo0ijlq8WvXuapMUPvnvGfOj956VjekTa7eXJCK+GfvhQXgvixxH5djk1eS/A
C7NnKfmgi+x6YTS1sbCQL8NrN8AISgThvXKfFvy962oAoGqcGfHiug+Q+38Aq46TmX2arsPh2gVq
B/47t5nqQPeLgBtR+pfllJw2/yfPr2JAsaqD2lGrZ2BXRqZph1K0T2J85gGsJ0uMQmR/jdRVSSMj
DyO/h2B++CXlwp+Vl+BwfDRs3/v7SBuOe/upEy+84g1aYZjzSIuEMcJVFmlV67jz15eh+meV9PXf
SfT2UQ9QXlacSGcU30qBlOp30BL9xWDglsDtMKSGnRIt5g8GOjF5rG9FAmRThYoJiQkUy+C8Bj4M
HRBoNUzejX97Fmky2zATvTI8X2Cx25bgmYUzI88p9cYolrCPP330WN98HtYWLpIZb55fX4GAbVBG
3dWZsuY/aTSCDrcnrSAeiPW6J7TnW8FtOMcZa3XPGLH4lrdfkDWpq+qPPfMBwGCcseD9Z3pt9/iP
GOKFWApWTVS5O3H41wOS3z+E2h8wIn90evKam2wTOCW2RwgmwT5eLd8jhv7yktSDUkemqMAVWiAO
Gpd2ugvVHsoB2fbDJmmBjH3XlGBk6bnOPz0CAfIOHRK591C/eqNpz9olvFwd02IWt8056Ju0k7Ba
HMwWWxacZ1cMcsF7SIrUWdvIV79wTzsZ47axcYk9Tzr3SeZNdfo/fo5hL6+QR+6s7/vB+yeQSOWN
Vi9FSGaGxQ8BEOAkm5ywMuWMv1OOtA7uYIKi+o2SbbySNyHYWkhR6T8lntu5SwvT54NuGuCreSsj
RsKvN4nGt5BbxWEpKL8IaJKcGoo60JLBWU0gbk/7eoadxZC0ifLyRv306/LGDC/VbKxZP0W+JiKx
ACwth4+8+X1dpQP5BZLJflnIU2tnM1wKbOnS8EIuj4OmILY590xYdVC7TqLffPfWYdeOngSbNpi4
1/WH8lBLs1564HNoe7MpjkHKj46QdqAKAzJvDfsmzljAmGZRwINsEBCoSYJQyFM2CTqTHm5q6Feg
4XN1+EUgI4jPapJFW3Im71LGYxkWDRAmnPRVcZXL3A8wBVqlOu6j+llYmWtuXp0AF3oPAMinEEPB
Pd/JvJBgIrI/itvqWfJ1116UZb+lZIpSQexRL8a8rlCrDmb9jRXzh4njr8IQvPvGnb4EZ2LlwTJ6
K1oknuj3kBi7e1t8NeDMGbzhPisfphYnWWGJ4Hax2EUN0YFSOxQJp1g3hiXiHHgscF3Wtzaen0kN
yI6db8EdW+a7eoCemhtwF222PJ2dW31hzrZKuNgxT7T5zLTf0JOoeXnQVDp02O4NOP1DKoQeheFi
d0uZ17l4KLdfxcNDdcOTnaLs8H2SnwljNlo0vtdcfReBHuUG65rUu3ZkB3R5luqde3Wk6q4dgD3r
wchnIMVz4202AgI98/MvXBlPnirAVIKHXgOyabFcr+7al3XYpE018Z/J4IEtkKid368PBZSkpHT0
IvC1i6JfP4aVRdD5OMSfJGM+jQtt5weHsCrmNEbO2DSy9gUMykc5OntQk9CWYgVrVRStVtrxwyCb
9ztzN/6qdAjUarfsbG0dkTbZo/dE4K3c8WzHNP2GFJyVpwxmLImJCaTHkS9DekzgjRPeFJS6ptLI
eKOscKwGCmWKHjiSKMaeu+jdpx562sPD/niiAgwmV0nFlFc5Yi4zGf3zhtsUGq9WHMuQryzIJcq6
nSm6EFcQH84Y3eo+SK7V+aMxagVimm1nkEjxql9Bijk3rtCdv1rF0gAnrmUl6/oyJCEe6FE7+27e
4JpRMFmLKRrtFSE3kLNgbbt1LEHG3B3FYaDmYC/o50iiX0LqjZL83VP+jqzKL3mov97PMb60DuR8
1wxAvsjweof5ZJH3wU2MrslGR+HxtZNdjvE3h0pgqsZWgB7daWgfvp756aJkMTdwULWSyt2hceqQ
QRqe04PV5YSb2NiKh+aKGWPo1nDO9OB4qt9XuGOJz6xKTAvc4w1ZtQ5nvIiN0cKcL6OrN9CG3SZi
9M4P61Hrk2ALgcbTEY59xm+K0BV6afmPN3LeqmkwcWcfDqE9EbohilcRPeCF9qGH1b+gWr/b1S5t
DNNTyWrkovnfp3HiRJJbuVAW+FEXfvRPme8JXvdpNNbOb25o50me6ZTIvngkJjIk3FHYD8B7WN4Y
sFtQ464sufoV/GVGzjpbpw8JjLo/q+mBDMnfT5bcSAyrP0GyCF4eCyCABfuuHbSFNKb5ZEt3+fiX
brDnYGxvASJQn7NmGXazL5MBbED6Keqb6kBGMqHhTYDsXBIbo97my7xzzv8aacPiMPv5JqycYsUM
bxiHszFxadIOfQ8yx93C1pbR7d8/IhqGUabSLMN5Ruol1EeyNEUdUmgfQtxuPIxKHxmxXGTPRmk6
TfXcBQBENd+LPV6z71tABCVpeXKGBvPBs8YjGKKL8ddo9tNN260HADnsd5DRdb09VTSiOd9RGc4z
65nyR+E9BaIfEYEU8qZFuU1aRJfJmmd1IeIYlHzFPlC7ZemH5SaHGRcvJZ3fNA4ysIvnlKaRwb+m
ewoCLf5b/RHE3kXUvMbOoewrCQsXPLylAjKyjiPOywYW8xN5RqcpekpGdkMvgc57Sm/TwPMa1GcB
029W+e5j846nXExXKCVJNxS19RnhLGaRPrXayE/VwHxGnnOAbcxcEOubtmaJcqf3vGjVMrB33WO+
z+/7b+AsrbvqEqLCBQUihr8G3iaxb3izcL3i2aIiCgKjl3V5HBMCZVN636Xy6qbrcFlM+63EQaAy
mlLMCS+A/3HYRc4tPqgGFJ/pl8VMoP2NJaHKMynZhu3XnwtbIHUZkH4O+9L8PXhhvIFXiXKGrkeD
VhMIhv4O/+ReOgjFzNF9TQfPtLAZHIb0y4sm1pJPCX4oVVeUTaYi8OaPVSnJqEAp9di6TC9yPFYt
BCdnJ7nf0rAP3+14jQCvJXlNPPoqLRiU/nXvJk1zMixBGKRUR9WAFFhIjZejelQttBRzACNv1BEQ
97ynb2V71e6+b8zpZLJNNk1UrK1ivHFuhw9ejJMBXOeManOVkHpWNxesgoTUOgq/lnAP+uTLA0IV
oKXKtJ60OWXrYpUYnos3Gx0L/qqrFkFJLlkVreMeUCFVqjS6hyLGUyrRpb6W/rIp3RruxYdGFIxE
F0QHcO/6MdTOgUVyS6/IC/86bQ7ohECou5YCl/B8XqEcCPKjGPqllCMDu42afPjXuwUBn/am+jOf
V6k9k5UFkbTn06Fvps714dEDs3PhCsDcNHnb/t6xLApR9EcB8L25uJ6M+gL/I7a3unn42cM9r9Tv
X7mOoeVbsoLztWmZ7CXpxH7DdMfhX7v+0edDSsBXdK6hNgWZFZjB+NP21p+Rg+MEOPJNssbuq0Df
VoYFh1myGsy3ExFqyRsX1i23zJ5LGUg2y+iIp2qh4YfhBYby05qo2H1W5u/nPt25+EDSp41hzoGY
NNuPlHjhZjpZIHbJzYgOPh2UFpwDgUPMZDWI+RuGA1HUqScnb5Lpv6Qoo9Q+8TqmwTJhGvqxMH+c
oqIPrzpL4H1WTiNH1y/iBR3hfpqiUIH08o4EKuTj8txN27EdQovPstifHyW7QhCHmBBQhXauHywz
lM7zozqRYSnIRcS5owLAIjWP76vgVJ6C+gctx8zO+QYPgYDi/fk6tu1RcDqkPFdNy0Qr3BZB09WU
U4GQlc8yHgucuGaRsXaPrkAadPnJNBUfrDvkY1044ufnsP3hKTyZ4AcJ2hUAI29zN0iT/eFBq36G
jwfaDiLVpoFC5OJuN90Xm4mWRKz35+OwhyFLjqF/eIW1loEsjrYLK0vQ1aX8f+jQWGrm4bJiRngc
7QiGwvW6lxcNgSll+yx03FMp6aaXBqLd26IATxzh2E0H+2JtymZJFZD6YNNlc0xnV3MTWyjjqzfx
FV7BRCTWaIcgCtIKcJd+V/9MoMKmnoIZFx5oJv73PKt3fwIFIglNxghePkpeGWc51DsQVmCfEyFR
JyALWBD/vOT5fHJ+ewPqZ83HDT4XUD5+4UopdL0viDChG0q5bpIQRg6SRdQFC2rz3YvToH84n3n7
J7S5u9+BFXfJUJKfkeTMc0rWBcrjuym4oqlPuDUaWQhgTdZf7QVo1RfO6ndXafT52q8NT5GzklvM
zsWNFLCt+6dTDmipsqpiu+3lUVF9W0ZzY7AAIpwOzl2SYiOODCOSbY5oGmww6IXKijrQrX1thU5J
7fsVNjCL1IOoAmzkquqS26RSdqyN2ulqtb0+XjD4G6SuSiCVm7jUxxyjuNr/2GGqqHyOIcKYlzC0
+0baTF4x+4n3Ors8rVk7t0Z+DkVHDsioHlPwgcGln9syYbRlX2BNLCic3OMve08+MjtVdYe8TpiL
HYzqKiEeocZ7MUtH0gHzMGj9jCa9pgqnOdd5penKu1cQKJwZY4pyMlzkXs6RfmsVHEdq6ophy2Oh
9rwXS8edlXhcI4NIniwxR+h8Jy/LCRQS5qFazfCG/IMAJ6ZqOgfp9NKpyeshwwL8X2ZGjoO3yxQ/
t3/4esoXxCiu7h8P6dkQAUNxRPSnjiOrNc227JycNXhRkCXv/s1av2vy0SdrBatq5L1NTU8SJcyC
5xz8P9VzEIOpWJb2Be0NGpV1+GONAty0Kw6UIQqk+CJKDa5vekBKmejUiYzkVoZ6CDT6Uf/FeASV
z3rxoQ2oWK8pu+47RWgt0DwVcLGQ5zKNFQQbqisAAsWZmAZmndWYK2FPfzQsc73z8SP4svetmwvy
/TZd//pr6vUDzT27degRmNptCeZY1/L7oCUEf/RlKhz1dytvu4rKsCVbwA==
`protect end_protected
