`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
s+nIOjJ+84fT6nRW7Zx+GNnrlQI9pt4McN/4jWFN8XhRnDPggOC0VNUnofh+NGvCBFGRfiRvM84k
yjnM/IkwAxi7Iw/9gujLfn64Q140JCZFojGiwT3tcD8RszBqoo3W1k53zq6fGkWEAyPWcG8OiQ5L
2j69ua8wp9ecEhcYJ3i3lt8SsLMyjvZBWiXdrtRkkuKaFxATdcHKbQWFXSQHJd4CgFluaELAN5Fv
888+kpxvAlKHua1zNW8kztX9eyQS6RYqg+ECKaAdxGheZCXQ/wLpROdWGgWnZrqLFtP8c0TW7+Hv
LJ432nGucjFrxN0B+N7mfykEy9QripuiL/Kh2eO2MA6/s3aSvSFDZvCx1RTtNJA6vRpJ1zRClwzP
FC/xANMKBEBfJBC10/z37/72ZuQccQbVakTkFT76ew+JNdGqFST+Zw7DHVnhDPlQzmtCpy/+wct6
IT88SR+8CDKQDfbKsnB7KoCRkFjGhnxH5ffXdhazdlF8bLb4UeCmqyFO++wofiYZLR2ZWU6QcN1p
KMP1Zvd2VcQKY+bCq+n4gowOQaOMGKi6s9VvZ1BLEW/cCLvc+Nm5XUh6jBlwx9MvVcFgKlTE+p/0
hzWwoMm5xlF4Ak6PihdU5dMJg7erv7I1OpKqWbCHZxmb4yb3kJ5NAwzNUFCEHH8/VIJBTS1SpeLd
W9dSApvEmPcdCO1TY9jxZn/A8HjaRi6AurNlTh/ApV9CPqwTgt9sqg9POAm6NQfI6RFMEo7kMAwg
jdaDzhk8ljKF9obHeEtG/v7VFTDl0bRFs9quTBZWpfIpJYjftKuK6ap0/dP+Er0fv2zvhT9u6X2K
OBQaNDPCLx5YZIiC1LbSd9y1EefRz4VCdB7xJPYro9cDGUGfmMEw/1HSDh3DfLNzU/uQgz7yU0pa
YYJ+h90ZXQoDOpuvvH6Cc4cokM8o9ByIYFHRI4JMUeg470iTlmgHV1yq4HIXyseFbpNzqzcy1lU5
y9RQ5RKSJfYyIOk2x647a0O/KDPz7iz19YGGZcb/13E9xsRwqOGsmKp9c7gpIO+GqdOUqOqLpxCo
QWGbuwo9VKenQeKvxOWL/yCnrJWCquDuNkyyZeJ5IK6hYsZo1b7nD8j6REz1pj8oxcrLWWXh/CgP
2iVeoz6OvHtz2pfnbcJQodlSsMMEFylYJMr5FNidLRq1crlbme8AZ2fZDKP195j9OGZIEMIXflZe
I4v8OacViqjEUSuxbFB/Im0GPp73w/GBMLO/6HH9usovD+K8q0QsyYk2+/FvptPKaPHnVD67WlTB
Dy6vAMc9+3l2ciBA6qlosN9RMsfL+u6KyUaNeJwaoGPQAGMFFjst1Bo0BVvuSNhHDZEfLXrg1MwQ
teSRLy0rTamcIoMIAu4r7aanx9gsaMF/6rcbFBVAcnb3dqQP7pWdl+s00MKqhB8uSQeelz5c0lDc
hu0Txp9LD2kUs3knFV9i1+0Hj6thk7VQgoDeI4YiOmvcNWYKc1TTir8vWUM6+sSGKPhUq2+KTZwk
K/MxQwzoYGW8tDKwOcOzBVB/kRS1tang40IbNJuXYOiWVKmduWDIQeNKAF94ReyOcZobk9ncy6qS
hsLJZc4Fa7jPoFrs0tZwz+jI0YZmBkSNYF9um8YZIvhZHe7rcL5eYOQJAj29M3zpk6gxHu/A+XHW
1YgdCzwH45cYrg82PbU6y15nU2I4pSwdUFakfF/Nn84D+S5hZQhInD0ujb0JEJFVmwElJgSU1wW4
0bF+lhjIbpdjY0r3Snz9cw20JUmZMEcV8/FdQFVHzxGWWcjtJHfEI4QQ7sy8AYoIeN0QFDvwQk+1
XdgPHi8o/ndNVSCE1obwwUOtrKzcSKgE3y5bwkUS5QupyO7MOjz/PZ6k/Uis8rfHRsWlUSu0rCJ3
EqQTV83uK43W+TJgrMDa2Np6MVs7cZZzQKA9/Dn2FMcMdTYTk/9tcTm3T1C4Ffc9GCFwLbf8aK2o
UyEYj9BEtVaJu+d96umxaE5rVwQsq20QyS1oDezoZpzUAN/Q1vNzrNkKsE3oEq3L5GuR7f5Us/RG
9MjUt2R4taD8E2juio1CAJfmNpaJ2ODi6uAcsTpP3jRgTzWABaRv/nWpc1XU
`protect end_protected
