`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11632)
`protect data_block
0USWSUGxovGsyBJteYpEocafzmpvNR76SJm85fQVrcQTsbSXB95tgSzgSfH7MsHcZUa8dENO2tKf
X7gIWY0ZRil5kc7f/IhTf+020a6HnbHE2xoalEg7dgTlLQb1Q6h3LtN7Ewiok3YBDeoAys9/wkVn
MK8/uX1GnqBUwFWTl7RopcDBL6BxCYjRSj3EWstPeOBTp4CoOltOa437oJUQIdr/h9ltjUtm0a+Y
nkfabWs1DNt3LNbnPzBjf0xmhY1QMFuXItkchiUcyQf6ZFB9lmSGQW9L1gair24aPiPwus4DllxU
5MPeVozZpZfYqUsojuvqJ5BSiKmpkBmT3YvvSJncnwA/6/lGi1sflLx6lqM+vT6AgJtOXJMRR89p
t4ik30ycNZOcAzIFN2BAOYKLMxuXszZgQwI7NTcr1Bs/kNmXW9XjRuAAw31SgcEyMgsWROW7CxsF
pNIHbDbDlXwKLxN33LUt+pYM6GuXHIGitZ+meGZ2bvzkI1YE7TzKeNTitcbd/USJWpzsWcx/zdWf
cvcERrp6mP0mexSjDexqEUGwgZDYYylxoyaZFezpUS7iIMoH6D0dM8SYIY7HYg6hcs4bf8IxlJne
jFsCkc97G7+Wy8tI8D/xYlQbxSf/6DrQOdpA7UdeJhUyEF2GQLM3AzA10e3w9NRlx9DvG7HOT3O+
kmbpk761EIzZS9ERItSIFZOKZTAQvmd8SQkqMzBxKu3xsRLmKp+I+wb25hrrkDfxhK6/1dKXsUiD
du5cIAryOE7b3sB1artGuVxTyjV/M9lwynUuvKHEfbSxR4/naD3Km18Xs3JE1yb4nxTNyJnX0yMK
1MF04NK50BLukyi/15mFRnjN8RQcUvkZyPxPtHHr0ooX62CQo/PeXRyBQAP7JyeY+UlX9/ATxXay
F3QoHcYJVun3YURXsRyWvego6bJOyCpPmOHfINyu/ymkxQWsl4oAlFiYiGT9Pr3GPdB9rrzlhpOh
w9TQ9WjcZV2eZoNnyzUC4g9IGQB0z9GuZM/+Dq1TOphPgJdNMhxxdfhh+mmppSutlz1xSih0ZFEj
BS3/siClZ8b5I+S8alPOpxkk0wdXI/Twmu7YgUUvWj1hEWFmDPwE30MHis8+KeuV1zwtMZpky4JT
SP4qcbFn1WAQB7Xoz8/vPBQia5O+KFVKMW60WtZKbWdwVfQKghBWp1DmSV+h8POy79vD+1oFRzjU
vMHjLMPBBvDRxHvq0qp8jgFLdErnzPqlnl/QJVlXcVLl0TQ6k94xvVcCwwqGjo6RUXCbCCZYzGlv
mYYVtbQDYQ10TGaHyaOJmRzit6aNTXAlbl+sOi+Vy5+z632vKvwIxdPdfJDl561Q70Sq9hOPy9/I
ILEnVf1R+A5swfeiwAyrhrC4DTNVzufHXSDJ05DpJ6GUeoVeBAC3hC3F83Td4ycsjMhkP3t7aAcq
fXem2RjlCNEjXBzPMqRGQyaANX+4MGx7jpFJT0ZZycRLhyIoUy1Yg+PWmhoAspo5pRZJeky8sELr
Ju1+S3WLpi/lD8Hq4Lhyrl1QsXxL9vPatgpiOMeaA7lhxHyDvSQtpfH+IYYQnelwdBojusbjd8kM
8AWgQk00To+vBHRqWQDbLxfOgBI34K9sVEzI3ONsRwRai15RmLQgrtX5NNmU/Ccv4eMqfIgmD0EA
7GEKOJyXyp3QA1zk5YIeMorntTqBzZzWvsss+Cfh5Dea3Wq8l2Jlgebc8XLb4mQzfO0YZXNUoXfY
JMs4Yhwib4bBFB0uxulS4AleeE/QeRp1bh+4GKF8A3qBeMiHpsH7LYVyWzVkYo999TFGLcnFKftq
qu+pHUws09wU3AH6zwfHaL+YcCqVK+qDu9DdN/ExVes9IbgjcA92WYeg3rXy23W2SzgG/FxENlhU
68YPgjLu3J16LE/EVAZJzQdha32R72PagIr081Km7W/67bifulJr1k6jUcsDJejOAzN09IXky2BM
GFahgNPycbJHlMxwmHRvqmuRnezoYHH7ZGGyAGGk2H/KsmHdf2ddlnOY0vkrB0SoPW7rZj1TBums
9b5BVTT8fgsm6dZQev+k1boaXmXtIhLdYoRwiPC8tFZfmoWcrIuY3wxjWqfgqjGmtKJ/7a/ZAsdI
tTS0BRCZ6PcN3Gl71eQS132GnGzPmLs4I8E+GrMiBrakgZ5HpPv1P69Pubs+cc4UeNDwNHk8IQaU
632uv9hjR537qjSjD6DarOnM3HkUK8K5JEvVLD61kn5KwLqw6TAERpY+SZfOZ0wmPy34RIP0uJ3Q
nbgyDND6GW1rgNF4MjpkCORwrRRS/Lykt5E0OiPEPwBqMDNc8NBuIG3/Xbu9UUd3Slv1EjOOJWAu
W/dXsJwEHNRhIPtPcKs4rZSoTpwkn3ue938GBE2Aya7prIJPuo1O2JUPuAcJz2x10IHI61cuI7qG
vIbmyzDDS08R9MJVHKyJsTG8WRlzmD1lWQSzLoujRO5/Dcmgtl8JDmCth3GeUolWDxlTBLLQm6MN
NTT5SfFIRHnOtccnUTf34KHCPgcj1WKfALR99x4jPs9yme3hFrWlZTkrR6l0QytcbI34pD9wMc8h
RSIpSh9/ejjLyNW6MqHa0fI6Ep0xFb5DJxZmBbG+ZTclq9cgd2VbuTFch4wOTcUMLFasHwUV9NTf
BQgFkf0Vbp5z5sn777UQelRUUeA+dV6ncyKIIa0jobA5dnPKw2a7EN5jO07Sbkyo8p5srasOf6QO
n08fkF9SRemXfuF/yuQAWEJNwUUduon1Umw7h26uW2KC6XsLrPNsFO9jVzJYRFUXUngkjYgLXzx/
ArrvIKntBUJfLsICwH4n71ZgIx6YtIpItQ7wDQ+EC/zSOpMr3ofM2irtdOPoo83AleUyyGYhuE3F
MjHEudJrF6PvkNFHd5Ihkq2QG/AMaFWC8ws83wkv9+ZWZ/PSHHSHHpQjkzdpz/9iI34piWccxs88
0AlBUTboYa1Gi07vr9Tl6UN9rxzygYMHpMsk0i/+0ByJDENWgn3rN+LEGt7+JmZ0oJq9R7mJUIEo
52NU7J8fVsnZ5ybV+P59P0mTjt5Z8zMFa8QHMBsCdSo0DzF5KMoH+qbi01A+2lDeNQRoZlLX3lKa
RMTD8UEigB8jgIOAplZ/Gwgg10ThD4amXf2PSRVdkhPOHZKZKultNAEbHsW8YgpCnx1vteoNbUPm
nafi1mzDixQBsvTYbGwEorVCTJNAPeSyg0nsab6rmtV64/MJ3PavCrBrNkDeA7o38SiTCQ6hY9cq
ZtdYy+UJ5MRFfqmrV5y5oqKi4meQbnQEhsfXcnVwmGVKgGR2VfDrHnowKZOWGwESmPS7XhNfDOs9
lh4mBLsaXOAJNn0UqxtYcLoG09iE11wjqCOVvwDl5mDPVXoGAX1DqmmKNb2eVtRLA2YiU0PdFfxo
9SDh0EH/Zk7DVptEBrvEPl0OqiZE+N9oQXkOIlVGEeZ2Orm5BYHmLC8xwkD+Mw83dVhWaB056TjZ
5ljbussxyJ7S7ny6xpbh0MjE9Mpo6mrcA+1bz8bpOwYDO1AchJeXC2x51Ao1vNigC5y5VqsCF7u4
bEWh+9ZENnXi9/e5nP8oCWGAw1fPl9dalAY+DjAQKqF6FFrKX1go65WT/uQOxFh2/co/9QW/4OYi
2Q9/JLxwIRR1hJgTNONZbd6vYh+uDvpFLVi9QmLX+BdODr3wAxLavT9IEWRKjfxr9B2r5kHBmicP
Na5V8Vf7rYcc+dZKj6c5UvmkQp/5OP69+K5VIGcPoMaNoc87layi91trFc/Y98MphfzLtUqpzrmK
un/HbzTsBumzfORGy3qkyhokjkpiOUQj7MqOeuS4mkU+vg8OhAZCYrDTvgATOxOTSQA15aHLprgQ
tuoGG+8JK1Ku9DJtTIlSVdJPPzISUjrNhtVByV0aDziN4V0Y4TfVFqXFt9gYu/nhpzGgs/ejzg/e
zQwYfj/ul9hqgsIREJ9Lde7irrWoYfbugZjj94iG5fIDf4vDsJt4/8nJVb+xgFCFQoIhXKFjtoes
GiAsOBbqQR1ApymdqCAHPqLBe+fyMEyDmhZGVcSyumv6rxv/oNVSs4/usqlq9aN8Zw9Hdxuj/OCm
MjxXdmthkExac3LCCA1JYjH1s+wOZ12kXoULtVYvx4N65kXtaYLoxzW7tuyWZqOUuUAl+RCht/J5
pu0QQrZnfng5Gfofp2NZSsbRe027ASxVysaqpkT37iXiqsbpFuUySpGrcDL6dxeZeSBVP4A7jNbc
mhKdfdHb/rvNacc/SHPmhZAA3A0fdpR219aN2NV+vuNCfKlmMQ0s2u8CGpW5oUGiD0IAIDU16Ixs
y7e96IsmcsZBwm31kAorIwC0hd4vSRmdr2LC3BvupP1RhUy77e+k4CU12cr8wJKrIgnS62v2gleE
HRyKAIGLuZsi08/lV3/qzojsdKSO6TI1dY0C+4A27CqV2DEZadscTkG88yG2HrXbimldHMBAiPWU
MFJBm4fkTLkCmVi036Ub3IbDaCzEVrUzZrW87Z7XrOYPpopF6ERMbXVw9RLnJBFDlUZP40Nb4cVx
LHIf20dGequfvc8+Hylo3Ze2/p43EGn+A1ZaxsjB10qbqFnvLh2Qz195jnBzdwt6Li2uZKyAL4jr
kV75zJry4DBEzrId+LZprzytZYSntKUMs5YixP0s/Oi8gUjbQoYI1qeD97jkJbtoiTv/N+hvJtE6
3E06Q4XU0maFK3Z4zDXiFrYPdhdK+0mVk6lnTV7e6hpjUyjA8I6uNlmH7clY5NZadiRet8tmoLmb
rc0AYjGk9OU8SqQVSZLtsn4aEESm7xF3WHdH8Eknc+NWIq10mcaY+BFwNfNBNpoX8ZT/7TSg7esD
IOIcmIy7GRtR7Y6wTBeGBJ6MbaplkRFO4NvaA7k9+wfYPj6rnaQLRHuPG6sdmRl2WnGzYQDtG4QQ
gxabA7ZSuKCt/QSslfMK1YRQor/dTrhDhJq2uO9+ZGLHR8YKtseunZaZ3S7N0q50hHxSn0kT64QG
VY/PC3ZQAeaduzTTsho3qF7Z8HwKmb6SX3xv0YqInJaxqG242oU0H6GOI+AXyz6ItvWLCmUQVRCS
2plkgTCHGyXYNOxgG2T/LbpINNWyBc8I2aCRG5Zxmb8lCzsNonNDHw7PByZGHI6+ycJBshBnJwjF
xkuTa67L1eKXGJKkZnqMTL24phrZaDDz/aXs7TL5soNlyk/DHkK2l7avc++ZAUBNRor60souSTjE
bI+c7umYqi6dB+w0po0NImyYSmbTZgGsmW0Fo2go4GMzUjp4C4yMKiIspg2HFixG1DyvzfW68fYS
6ILHj262eCK1Gqb0j5H2A5jxrhuTfwORBIZqJ7lzyrE6h9bHIG0udh7tS8pbEbOHoEkYNfjmNuil
ctgioR0/XI+bR3HXUUSD8Gf6PAekrsOnbonWnMT1cCP0fpfbKLPtKYeg2bIRrBO13S4mxm8qeM9Y
e8VawKaNUaeQy89x1b9xDlImP1ynvwvFpHfyqQ09q89HifA0U+/NfFf1PQt/8Z+IvpilirjjAO+N
g/KADep9zs5/Fw5AmlUEvQ+z4OA3zi3vwk/Vx7i4jO7sppt1v2aijPY/b+epoU/9S70AZyHMmqlr
6JXa6z/8lc1sr4NaEE2d1mkiG/VZLBSSG8POjgaOnbXWhNGUahtrBAbD6A41e64jOGOGDx2Y6N37
hz0NbAV3Wqm8lzncvfn3N8RElD9GyEBBHF4ChWi5tBIkspGnRCYjsWllkBQzcxpyyPFA3U7jI9Zh
r9rA8VKSuXCgG5Ov+6Vot8KcISjWWVYLyCH9LcQ/mQUCQiLwvSDnBdnlZiIAT1DM0g4jIR4GscBK
N+LcDBJafMl1IH8ee54ydxoiyprjD+a/pfMpIaT+h+i3LzxJjJczlJIf+msJ1SHDbsu4rM3qILeW
gCXlcGZjTe+NfmfG8E0d7UagkiggwyiZQPCPHlju/chjpt3FaL55CpAQVPzQgkccJTQS49JyKnFp
NAPmFhIEC0IKi/vUDuyI8nnkB2pwrKqnr5KdlGQOs5tHvBquEy2csGSDtZJxF16QCgCAN0c5Iq8l
KhjFdz1o752/v+pfm8PkCpBWQfMAv966yRcjFgiVbx9jlpT4fFoVpTeI/rEeTbV7ZxNQdd/8ijJB
wyOausxT0jmUkZkIJrOXkyLPh/Xwai9KdB779ET+HT+CcqzG4+Fkl/oJ3tzCUDTjun0iaYBC+mF8
F1BAnl8axRVt9uRSk0PCAGCCo01huiOIUjd/t3F00pM2afndvJuwN9sm4Lu+AWRzqmFL4AmdfgTJ
tCq66/0c4ELJAA5vvHdr45wdZAahs+Yb3l3MqAvstxpoc/VCwuz4O3l9ABHqyXkZMcNRoCdM7OmY
AFA1a4f4f2yIxRO5Hu4oAlwaKKC1xCoxoXRwOLb4cEGw5w3rFWZiBANBRNjQg/ReRz8oFoEVpfbK
Hig3ixScDpi+JjxdKXQqWlJ5iN5+/psqe8CUL+Z7Goo8lrCXAG3TQxOstHFVSkocb7r7+CyVDFJ7
p1DHcK82XE3UvTltJ27zFZu6b6lgeyoj61eKnNkplGO089DTD+4peQOLcTbXiGVQ6pJe0Nn9MsiR
NYnT5KfyGK0nl8aIuK+9sMzHQXWnmseuIwfm0MFOGktLBbqvOeaD1GwW39bZe7fJMYOHkC6iVLEE
reZp9pRGm+S1KUEv2+4J7h6+E/zMtB4UJh3bq/C6/WPZc5zV6AyCxf99iG1oq+vvljtwqWF+mCgs
p4/pLfppcbF7eXBsSI2znue9V5AVUF6PJzaC4BtD7FkNtDILmtSweqMOpL6v+cSmPDWL9kbSZ85b
AWkx4lQIt5r5ZRAL3lnUCKZ3OqSzlqsRuZ+Bepr/JllFqSVJM8aET93LVX/omwSO9dYGWRADQp2V
G/FEz9H2XWBj1BES6ZJJ4ALjJGRVt0InvSpWMslTPN1Hc+JhQcyuYxhRHrSOUKzwaXsRbvqPGLgK
mBdB6xn9BMkelwfLi5XN7PgM7e67iBL2LpvUlPtTAFrf4jffMDo1dQUICqa1stZOXH0KgiIGh6WU
uzi0XRUFE5m6nFC4L8ua7EG+ytSky6lRkk7w4Yds5AHdU3ghd2/j/cfcuUIEKCpi5CmmxxisIy7h
sIgazI84d4RcXDtDtvbuqFgAIdzwQK28CfjNThuogfat6CW/q8gbI6afhjjAgLfnb/i3MjKbE+oI
JrWIaSp90MuyW8lJIQsSn5VWr54tNV3lg5tBE+tnDdTQWk9DMSUboOMwnawn6Q6DLzkKEVFsHbJD
GUI7Cg3QaQdlnf91ngwd4aH+y4vGk7ehX4MNR/EI4JkIi9Hie/JVIVtZFxIaGZeD7x4rFALIaFhX
T/IU5/W4y7N/xg0svRnG5lFlzDAWT+FP2paJ7yp9Q8XTDA6iMcYu2i+vlX5Z6KX9YT6PMErLB7GY
88zpWjzh/kktTvte6GDZm3+iAqwHJB8NGDovGpvge4NsYajTi1EJQ4/2b37v5SSzalekQfEr6a30
viNUiVW+bPvA5RrhSRTZFoSKFENFNjv32Cc2+RT9UsN2G4jVUmwhUw5lOBZ5bWeX0I6iOcnRrr32
fMuG3Xft+ZNMlbGhcW6xG59I/GElFJOvyBFPH3xdEqMZ56C65OmIRcjVVpek5AYG/Ih5A3qxsPuy
GX5u+3jD43sM5RApekWDKfhlcGKPyyKr9uAr5Ta37pTH80vGfJTJkdcZmcFmTruvCPCN9GXcyJoE
w+63ZBZYlFgLYuNhPrH0QUZ/iiWFVrxxmfDFY7cyDJ/bxiJNOalo+DjLWxZ0srePOy4g2oUC8zq5
JKQp+fSVuT605iBjuGivJbJ5ZbnJWyT35eOiFkvOoiorZ8v74D/ytqe6L6IOQo1sB8/6GmhvNo6q
Lg6yqyF3JhqIRFhJw+wSllnh5NUPBhdCVMVbYkYLU2a3jqslGmQBsegcDYDIe8M+BfPxPIau7pOB
2ZUACCdkyhm3kDn/asJjANFtOGggwejB7LB6tasI2bt4Cb4LA0ITt4YH9hI89kOg2S0vsOP7T8fJ
cHc3j87zxmBcUGhe6OCyLM77OT7TBWjdyOOkZ0kXJ0NrR1o12tiGq49XYA/5giOIh9Hpww8O55HT
yg9MIl9MxoGkq8TbRCwsZN8vwyoLN86Dw3BNwEGEnibJqqZpp/NepybR1qmyWHgOksLSHsCAg6Uj
36di00ETKZYOMO79a/u/il8+9PRMt8+Y+EeFyVjCFeIWUFCLT0Sbho5TdgU1pZImMbmTdPGEwlHV
B0230+DpmV1mI9A5pMtyx4D6YFg9l+shq++iLyv+HALjLaSU8X6L93VpILULeW/TmDA3KUiGf/iC
3Z0ERVe4MwHu+UPeoNHHYvJnf1c8i8x1n2Ab8uAHiR+9slFTbDVzY6kcOL3ULrb8YihKiuSuMvQC
A22i3q/S3kKMyyjFFU9RuRjedmXi/TFayNtDYQ+64fAXDUHiwrpXXe0LpuJXTCAZ1q7E+rT1digy
oVjcAHT6CfiHZ4ykOsw2PLguis7JHiO5BD8wURUc+3293103k9/PzuBrJfUfgDHDHHnSy7jT+r6p
C0mNTE36EBGIQWLcnHbgC+tmJGG6T1UYWveQrY0PDS0vvzD6WuI9zSAGF02cQ2vU4leiLa1ysNur
Hx/ItVnTPgPBRR46r0kgVjxPOluJp9psIwuO0cZ2/kK0fJm4+54+A3HKf7SwdFE4UoWMBkW7o+PV
Qo3bmaUwDMtT3cWdd6B+QCgE4kY2oWLGAiLxFmxRjTkIynbr4MuyQKEXtWjBWEb0xrgrkC/Vntzn
uhCVNea7Gi+7BswNT0J2N8B7x4J8W6LTs9m4z/yg1RzMPZb5Drxauc0T9Ene13QWvWSQsx9KSdFc
5ew1HGoHV3uHE8TsxGssqYwOvx61E3OAx4Ky7/wXAHpmHwzri+3C2XwN7volmug/Gf3hjFNCMWE9
L05QBtm+ryrlnqPBKWH36kvjG0GhL/EQNTpoRuRjuH7Yvw4plOyAFhxNeH7GtOyoqJBikTYoNNYZ
zXLWLFcgojU2HMuZLBtriz5pj8YE/nku0r+kxRzcMVeVC4W3jpTzg4rCKq96GKgkcuJx7WGsIiKK
Occ0nQjOKQ2pJAlBUsYqEBUaU1slE2TOfXMPFWaK5A0L+THSINTqK2tkl9UzbtpC5p1gTk74vraH
8nf2ma0KCm+dAP415Mxub6pbZI4KbsN8HrzHpVo5m2jz3qaZNCRlzCyEuTrLLJuoEzMKrXdpfdVO
rISaM+w12xwlGB43N9wDMi/MElCiU+EERKuIQ8aNyeluTgz+qBODHGYn5N0x3V/jiHiR+k0fRCGF
zdV+k7UWcF2hYMeGW57ojsLJaEiCMKOc02YtbjUFF4PW/5cVWHEvSCPg/yRZU1Wn6s/z6yZhi6/N
klcsm7Uqc8sh3awQrYjocSQ17rz5XmoUVKr5JQQytN2qFje/VZG9H5MhlelSbWohOAIQgFBEfRbK
ZzBXqB+yqA4p1UEtm5UjFyK9l5ErgBFTGkhLJACqw3xC/WE8fR2y2nfv9EKAhxMhylf+sSh3Y4C5
2btNKuFqmNUabeLx81LbU3hN0FSnncrIzCN3dBPgZTWIThvy7VML9N6z2Ou0JDPdvDDCz/GGHV6E
K0FXDbKsryMVILgCX0oFUPQSm48QhltqGa4ySRiuNUy9NIPFQHhr1Ez0JxghZoC561vlOO+O6pRD
U0iSI6kQf+8C4dtCkFseZY5ml7tIG7rTh5DqL8ZuQQscezxY2Y1r99Lv0edS17Ho9lh465vl2TLk
1pExnJjLjqgfsFpFI3LDY7WQrjMWRMG6y0tMzMHlaUIpHeI0HTWx6i1aGipIrUSSRklFYpfLwmVZ
Vf4lJIQqZcoLzczoFut474jWYF+larRVdOfEXZ5ya2wMuuuieov1etnVN33lxdAX1ic5lAIL3b8E
EPm7uGs/KZ1wUn9IfUSBRZjJc1y9e78+DSbsAO1v7P0aLzVMSJ+87134GdR9uAA5Q3wkpxzinZog
lOvsOGfqKm/xEHm0j4yY8+NzQKx34Mcg7EaEiyudwdCeup9VqITSLdk4M4ADvGr4ExuCrQCNFt1G
HvVA2XLcOKpKjT7rztU/XZCpin740lobCaHl7FhsvGcfsSRn8W7j6C+xfzgRiqqH8zsBIN0QhWYW
BvltfeMNKrZ2kagxQ1Afp3GI6eIcsCCYV8WEVGiSwAICR8/mP2murvjKbfuuXiF56J1MH1TTjMQk
Qwr0dw5ABIXmAdfRKc0Bpm8fBjMVNLfO80hlZ/5sbSLx7SBZIBODtpJw97Wv0jSGx28QBfXLIb5O
t1ly9KrwV40g+LdmK1teMoT/bldcPoVW2wJYEge47hJO7xCpCV4lgzRleRDR6b/a/Vcz8KrfiD7B
jfznfiaA8t+479735B6sYyzEk6CBLYEYR544DcyCkFcgOMu2G4KoCvmT1fdObQgUG3mIOpAQM1HY
x5vWowCGbqlAMmRU/Ql+ghw71aaM0E4WiO9MfEQ5REEe7LJ/aprb9cQFrvQqWkBGQpEY9j0i/59Q
3IL0y+PdBKG/5c8bneN5po8GbXWPME81ISnWL71rNRb4oxAk8SrlNdBxB4WMbErizpTHEmvIlzWq
guwBrAUa+LcRgMi+OCbZXtBHXa+vvQsqFxto8phi55TEq8U0FIns6t7HowwpUppCSP2+i7dlPGyp
CHAFlafFOacCzUDzUQJos1BmrR2RJ739mWHWP7vq6pR5FFWWxy1mQyW0YXwnk8IbYI3vMf3Gd+0w
EWYSC+lrGcBeR6oU21Ee8Z7vNt5aiIauEavAB8TU4tbaE0+hZdsgSeJtBvzYED8xEaSy3Kb5btBC
jbl5uRUwvsH01X6WuqT50eYhO3jQKHoG/6fB6pRB4t2tyCdHUiTIjkWwiJ8LAtn3ypgar1qrrTmK
BRr9n1TO/HwPEwQDLL4/Pw6QyPV7W0RqlzNKX1F2CH55AjXUbBPt0VwZH5Y7W4fDUxhYjJDeS+13
6PIl47JtNGleu8Mbcs+lU25CJZBZ/w6BnTqdqD+CxV1L7U+VlWlHHfMG8pPyTilKH56PktHpzNlg
qf6Zaxo7MKxixYfe0s/i69rFcT3e3iLZ3B6xTa/VIaqo1ceVlSq/NxaULemIn0A4rxvV1lh9HIDF
cKqm5ZeLcYBx3nD4AMq0ImVGJ1jGBi15o29xClMhfJM+KJmyND2A54Hd37g6JAjMi/cmYoZFusro
JFfUOylfJcUHp2oayO8rQe3Rn8qJDUz4QIXdLe3Qp8jWDEv0DPkZuC05MCce3t8XwMK7TIdmS2+v
ozDXyGh3Ib3G1CxNPsfQlg4LHXRD42a8qrH72f7BU2dAAJ7ptMXnC2rewb7DZjzKUCTB0Y4KrN7w
YDg/uJY7oZk5t4tA3vDVf+SC06AgUmAPllnl4X4aWsNztekAL6QvmMt/aXJPHC+iAcmbdTaMP6zt
po2PHVDylcNfCFe+YAe0OA3oO4+PXH/nsqwB/D06d6veYPtmFDbq8I6NQsDzlD3lOG0s2q0tF32N
b6lZBoJcWB0J16RIq54wgnd/l0gOXxRebwl3doB7Bo/Iyglk9mk6auuS6pf+Qb3J4PecekRxPAjk
qLKv5c+dp4E+ON1+6ldE6peutdZr2FV6mTL1k58uuyiMerp16+55EYWB9MUHxsvLVsAVKGCFEqBy
s/m6bdfaVBwz+um4+tMRsha4RXF8by7W9vuuHZ3AQ2wjjrAOJ+m9TcYJQWsN5nj66nfofaWR6j6Z
HNOuDtk2nIDhveIBnpHFgqJRdj3y+4uJlDtO/6Rz+QtQTUDC+DZtFwpM48kKRx+J2ni0FWROWdO+
fqrbpzRYdCvD5Ty+0cXXh1r5T0rc7au4b3gZ29lJ5IkjwrA3QIv/zCu06Obui+LzXmPQQcB89pku
aXM+lhbKDeSiqKAw0MuPO1udIvbYrGbC5c1H1ksCnZsUp6RFPvS14psNjs6wSilUTfdS4lVIdVcC
7G7FEOOLb+uKl6jBI7Bp8AnMI8YxpJoGPOQf4r2D/3TRn1q8ES8pSvigSXMRmPb2Xge46UOu6+gT
Ql02H1tWk0Vc6nw6XtzA/M9MW5YBHDx91fwSMlMdEz46dDKef5d4Cq+rUkVXYjF9KtMbnreqbJQb
nIgv0hnzyD/FZIqG0voIsKOMHWq0h8H8rxy40hht2SQaK5ouBPmesMl7Zk1Dm4b/w7TK8cT8uykT
JOyYygN/SkvgTH45krecEyte1IFdYqb9nh5dEbJx1zYM8pYczPAw69N739pbbg2rf53bBHOZXs+v
eNdgGRIde8dSPOsbAJouiYBsVOUEdmDQJZjVYXasUyQx1/dA4Yv3tEQwveRdkG2fVu+jeoEx0a7E
Z0A5i0Fgur1mx9nPUXTqsy5W5QCN0pC4QN6lHa6H5WWivR/vNe3ZSpkNwyrOXizyG6En2LYGeemz
wLpsuXXN3Zg6XFZXDlvckSAoAr+3ZBIgDiB1RZb0PvD7Vtp4jCl/Jv0yq0Q98djOUflcYoShD1ty
cZVkKRJFWqKzT216/H5+jyB2v70UiYsrw+/9zPkAyCTxj9GY16GJb0Ac+nGPckBv4/pPDTYysK2s
yQw2suJ1X/ogmFSVhN2iwDt4gGEnfTOnNU1hbPAO3Z98xPm5rluce9iF4cgzQrBS4U42O42E6ipy
fQ9Rj5mUgcnOoeDyGH+CRoG8fdUOC9D6Qwc/6NwVEx0ISwsZfjofg/dgrlg7RCEoOUdrWANCfZF7
ad4+fRQ4HpUnUErDoTPQDyCa1SxQU9JxwHrVvBOooU1FoAkgg/9dACS/3QCEo07EafTleJ/e0JL9
wQ/7nyuYNFTbJtel4gcKlKhE3iuie5ocfrSGUXiOcmiQ0Pt+etgJQ8/3P9yswIPLGmd4HWHFElkb
n/lqEeS0ra9j7gv8DnwzEzDqspKxm1+CarGLaFWwjdBRXWEQjo+z5U0BJu/9MjvBGYGBDB8vl7GI
axUUXNnOhS476FVelLpwQ0EvSHDzZNBfHZAoLPpJ75ht/mYGkAGkQLGQ4tk2kNE0bKBhHuSFCwuH
4ittov30fyHe18lIPDtmr/AzUo3GIjr0OiuFRf+l8dUpRCcC0jyg9xCiUzeJLCzVYpyOyuq3R0OS
T4GA7uIt+QsOeVFweMHVNfAgcC3/ugA1AkbLN43At3dPOl9FL/xHMGtKwfzrfpyLKFkw+lMGYj1m
1Xor5/7JrJRULocXcoY5FZuyj5SfN8E4+6w0SKpNTpeJ6766TraZXsGLfC8jSxBXnT+bg5R3f4M3
7hvDkTL63Jz32T0Rr6l50yTxqAHM19hYrU8RPpAeJNp1rlJomPf+UaxRHsvkG9vQXuHwCDsDHMZW
k8xo3p1XA3D6mjlLF/MS0G/rS+5PvgzzbXp0Pbkm6qlN/zqx5Q2n3cptE5aWL8HnTaTMXnwn9Cgo
b51T9vfos3X7KLH1Bojjd/SNt48l1bhDCCyObENHx12mKRsWqZWib3LEYPBD8f1ZV/yfJSfJlGOZ
5Ely3cgG8KeEzk3hUjVZ4534sbxtD+0OKJXUwr1wA3MtnUL1GOovVIXX/2Wy91ftcyO9hGzTDxV3
L+0pedjSUBvzS2whH+wJFDAmDYe8Hkhelf0dNqIBQiMBitf1EZoXebqO3dqQpakfrTC+Mi2U26FF
imIWdWSZ4GuaHfZZnBm58Gn85S+8oq/P/p3cOrVEOn5lvFtXhjtpSv7uMwmNA7jsVTJ3o9UfV88m
C5bsnV3kwRfPq0/TcqnO/gofqg4ZAtwXXpQzuaWphwqc3KmlErVyKqL9FcXIsRnZxhpI6DxKNSq1
RU7P7XZ1kLIVBIzy+4uiDb5pFTuV9FbFO8dfzlFKtqFFbrDjdfaofT1jBktbcJAC6GB6TkBRcPak
IDSyFNQvj7uSC/MLi8WW2XvX0qrVd9P9r7UCNLLRr7Ib6NGTNRMOj3YVsmj3b4S0JqxpKTkS52N8
psEX3WuV2HTkzZXmVOHZX8aUME49Yv1I4vpyfCWdJOQqRK/PFczxmBzXXSHJ6tpGbc4vqLjC4LJQ
kVTKXLWJr2biboLUteTmBktVQiCH+mi5SZ+aO8lWhwO3M9ZHiBYQaBOCegT6ukEYmjhbj4KC4LMJ
J3IwWT40tl/QoR0VjASJDVwtmO9un5N1KBCciK8BtYL6B/LoNeaQnKLRvLzEPnrqd9nJoxFlU07Y
ayBKDYOvwUsYB4v/A9hZWha6JgwE+dhDzaSJ9hoehewBHDaFoXkmcKCmUtLA86wrJ9lvNcGZn/Uw
49yXuuUX+yBmj0IyfBl8xftg6p+8Xp6yYsq3q9PoW/jTbTCCSPly20ydpDYBC4Z/UPex5zqVK+4G
kW3sQshxtF3ZJ6r3QTYZAqgdrSghhJSTqhmuIbVeKE0zLEH76jPkWK1RyVhZhRwtPMEUb6qjrKUV
oSM028pwGZq+TOnJo35aDQMkxqeOO8fUIGu8X3Q+Sz+Gp8CxEFq+sLT7roT5a8tf0LhYhLwKQzfq
6Jvn32/Ir++p4Cfw1270hPklGx2hbBZq6+5TsAnblWPxfD+farPJb1TT5Xt7FswdnnZAsu4VEjQ3
QEDPm7C9SyId5fNaC4QUQ3TBpnfvIJdKyHoEE2D81p6qYIWb/XPH6eLJSco6oStMRJ2jkVovZpkg
57oD9mBOZ/m58U2bGaKr4Fk/LpkF6ugQzMPJBgFuKZV9QKkLzGax83x0fS6vTH+QVMX259c1HqyW
Ro3TBKFN7eqeOJBnFTXjzE1xlB4ph9hn2DClzJmTXLuCYidDAuUBd0kstsLv7r6JQ4BQsh3UIvob
z/OFyIPuAZyZN6hKcNTra1WSBpjhJqb44snC8J80c6Iy7v6Yk7zkZPd1zFJk0WU89B+APvxKEcI/
MGJzWVLaY6PYk3ZvFedr40Ds4FSmkjWzVwNEXmBfhI+CTl+Ptr7+L1l3fQE69fBA86tHkY9E/BOl
LMv6GMYruXJpPh+weNdLtyWY/sBpAAae1uld8rYwRn3nt7CtFBjUT2IFPXzfsD27zy8+yYYpKGfK
3++SLLSOK3Gk04ZntL0vgFJ9I/70Y8/A9XHpiNv8rgYOtPrmz8kAFR/eqKauft5CIkWixsX53HOH
RCb25p9qNu0WQsZ5jZliHdnoj3XPkYvGx+1J2zsAqjodqRXWBIh6bRIUwQTT6XVth0Q6S/ZGiPbi
nnqsiy3ierhC9ndFZebQJt48imYICggu4PzWuTSfL913uAYapt1smq0UOAq5HWF145H6Z9nXiYfV
9tzgzprK/G050miwLO1+fBblI28nuq3lJtORXKG9OC2m2CzDN6HS6tImQTgpmE9D4H8NHt85SJ1o
DZFcMzcJ/fqbVWDoGNuBkZHiKbavJV0TjOeASqsF/pbcn7AKa6+bL8ScGZkwKmc4n7gk9pROr1my
K7o7CvUzSIpoDo+mI8X4bNFm2730C/T7rwYTOcoaFYaUr9fIz9hsxkgmVcOq92TLFaqf5D0m+W2F
hoSHIA==
`protect end_protected
