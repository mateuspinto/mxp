`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2448)
`protect data_block
FZ7VtM446FKLOLxSj6+L08ZmFgDCW/9GLgQ9zjJ27N2Gc67HIve1PICk+37n9qsbTL+egSqzy8HL
930is+f5uId3d27H0TsPmnx4VN1qZReVqd/IoE5q4a2sK0LikgH1iXxb8PGaFEYDpe5CYonBDXh6
sCoMNKsvuBSwWh0QXQrt15OUR9po9LC6fKrPLQAmyyPP33f2/Jp0aAaHu7CYM7SX+xXMYQ45Swqu
N4GV8Y50czzNrgdANi68G3sWQ4ciMfik7NP7eNkwn0Q9NzLZQmwc3NGImHt0j0uD3zITP3INgrVl
0Roh/G2iM1KWdtEKMmmaW/7kvJZ6CjGLFy/f6vjxZIbt6Lb/01yBORlHMgCA+Acb4gMGgNyhz6P9
DAnTRkFOpX4cCeae6+gAAXxzm0OIxNZyWciKcsQj6OfxfayDYflSytrqN5ll2HPSmIBQwjqACknD
YDnJnMZ5XODvP9rD4WhIvmbcmeM6Iy5Ee21lwOhzK8+mq7nuEZOYqa0SiLE6oEsfnRDEljHFwNLX
gbmE5H4e0cZ8y0aOjAPPe+QvK67uBXL+KbavQkLWr0Y2aIW4SR58VbSoJOlSgzMbP8hr0xeIiDop
OBvqC9VvhHMOe+3YOVrr9Ipn9wOQZBSLE6VVEY8kaw4sHV2UG/WcgDgw9xQjsNCDkG7AONik6ZJs
3XS/2MYYuEzWUtePdEorPx2eG+LEShTBXDX83H60rbtuLbFbeLl2dBEih4+t9pYIxygNKngkEnUE
G8sSHQWb9dYQePaUtjsAjil1ZBw7ElBJfu6t/a2sFhaAyG3TPJmT4TQuyUfDgwc1bByt0X21odaE
NNirSaKm5/hxgfZfXtLjbVQsAOropNVNPVLWaUNqlWlNPTPe5GPjQem0ig63W/OKvM/OgG1ocxBP
N4Ito/ivY8PJT3yy7d4trga3isYErn+nb8EYRDtFSu9akNCb1bRUjl5q+j+mol6Jq3gpsxD+1qkR
IO4rwUGmYlkRP27yyCd0MtTEWkYsKgf5B7sXNVrxWVsXZLdqjA32I7If+RTEj3xhax3LYymW+js3
6hsUGHm7II4nN8DQTpX1soTKT7Q/NEeWkJ0r41aCxfQ2V7n1k6HK/WVZ0F3fDwPd1bA4EsISOFLn
cCUcF9b18rVQBApxJwAOM1x7h1AHJcvineIFDRwU2FrPTF6sNiDE9L2eKJKGzrIusIkT1c+Cm9El
3RrqDrgJPkU3WaeGAxIlF+CKEQtnUpu3YKep28Fhrizl2eVi0Ck+bp4k0MTxur7MXcyffL4MX4fh
2Q6kFWjEVxG8WSz04rB/u4N+eWoR0pjxsXX1vDA/pbf2pUcdt12DcBE+cd2/ES5euXXDTAq7/E3P
gpd4ikV25dLAxV5/osmFVI4MsjIb7ZX0buG2rD7ySiAfplGwO2D1GMtVwR3cMabZ5L1T1oU0CZoi
hwLHgJvBTZbfob46SjBOuWHy/TB1zhhpU8L6r5sT/Fce12FHUAuFQuEKHI3l99/iqStMpvR5bJrS
2oD+wA1rKjXFWhZF/6ZyvykBHqi4cvQSHrRdoh2W/IdYRCv6vnoR56aIHYircJHkZ7Cv5HtyqBZT
+uZp7s3iYQJLfR6CA6PxfN9aJvbK3+N4Py2Ky/fuvpw+DujLWORkbQnQ5fCToz5syjb+RTZE/1ni
YWK9cPmtynxiioZ2ipdOAJrvDLiQu+DMGcxLAdlHFZvo1n8hW60luESt7i0PNfq1fSnll8v/4zBg
ZBPmaNjWttcEiSaNexN0NqM8DvTD2KrabhoG4hnsalG+5RsDjZhTTJi0Src3s6UwY4gw3agZ26TH
j9YNJEg9BvJIc2105ofRQfm6pLMK+ZRrRjdzxg9GsBwiBrYovw4Nd1wgIBhJQKJ5sFmMjMNnu7Zy
79+OvdFDFAZTr4l9vQfRecnUqrIg+SHWkzvWil+p2eVJ4oKwoG7wPESeXUdJfHLA2nBfRmGjadTh
oU8cqnvDTCj69s+5J47p3swOS8WibV3VziaY3b0v+nJqKPHgGvDHab3nz7+AFrAquWvpbTVXZZ9q
lQRGz1bg7Ek/Izc6haiU+4HDJOIWrOYEtd1636/zaEIwai+rgJ4mRCdWLyaH2lKAQKDiQIFHSB5h
Mfef8HCSehkh1xIZPKOMjyyt2AjC9q4Wf9ajcPm1zGov+qYsAn/i64YIP74kdmlxUcXqfaIQysx4
6GClBjGLNe6DyaSwKsBikEr4WKzXvDrsFrhj2jEUh+TClwd8vVFQ+pWgxk6I5LJgJkWpFHWdbf93
WNpOPAWIxKf5ewUgjSzWAmuxX+iAIO5vOcet95+bmJyOtI0bdqaMG/TzT74JoSG9jwikYQB1wWGz
NyIeSciJu8sHhAS6v2ow4LLNYXgkg+R/S8qfWhgms2DnWbamtcz1r07Wy8wOALWhQd6pD4MiyLgJ
F396v8ktpl/4RQwsTFfoI+1xSPTySOy+keovhEazxBgfBpgkxGAaenibJNyuJKVybKfY1J1MQHGY
xFF1AistvwUJ3kYNDRFwDc2DZmX6UhWlml1S2v/9hEv/0UV+iHe1OGDLvtZWOvE9JXFsG9b5tNpD
Zf7e1q9WTf+niJKyug/MZ5eVp3SQDyuRVqaPh780BCyFabuL5mg19fCMylpievAvA4vwuP9sCF9D
iBTdKWmHFXokTyyjbMSjyHpyTqfVuqxu7ta+y8zb7jY0vRRRMGeHfzRrh3Wklr9g61YQSUZ1BWfS
2VGK6roURcGlK76QQZuHsKJ/D34IVSYbRutEbzZpkLEhndyRYQ3SbdRtFU8Kf88AVOkpnkOZkftp
CZaVmwxwtFFGhWKeqLW+tamGYSrfVOYKRP+4nNcFZL9saIa3Si5bNdBE69OGGCsa2KwsjVvtSNsp
CoFeuuJ08ICGR9CO48a+KJDzLPkD+5DxiGekS3ix5OO0Fg0AmhOIruuAxxUGK8GrENmTYnT7Mvsc
V6AbPyoOmmi9V8ShQE8nNF8uG0thxbZou/MqX8sYrCIkxh3Nqwvwqoklw9smxUxO2rB6ohNal8Bb
PsDhCVC8N1hs6qzj64n8KqVOEppkpg4qC9jtcdTlaVoWEA3OAdqhtmx0BbcXOXG7d1YO8KDV0DSi
/HZbyiwh4udUGSdLVdUaA58p170D/KJM7wwnRC7ge0F2/Ry+SSaXBMDelLhViySRZk0R/8bbpbWM
MDL1L5EeKW8yhf5hx70xweCu5NBUn5oqAUy9lEx09TW15I53GmVDxrK4WyNok0zJW4q2xtCc
`protect end_protected
