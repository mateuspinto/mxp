`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3488)
`protect data_block
ROBN1lHUIdXw/Gh/2O/McZH3t6vAbw/ftEQvqMWjhDVfWPRflHw3fr9CJhYk6vqv5CMWESnbpPsN
cfWaGeHmP/GYkU32rN65BlNTsXwIadWTXKAHKMPUoGKB/cKbIl3bs7VFWNLRNTrnR32jP1qDl5+v
kRBZsSHlDtQTx7/kFeyVJOEieVihRbimG6Cev9zgV1fvvLeAV3OwuNYYR/PvINfrUXIXkHJ9Rf2i
5R3A53nIxivdfRSh9JIjjCLSWiXy+LVNM8L3yqC3LQwk9eHJ92wENidiw9nAYqS5As7onSvVJx/G
EoMN+uDfVKVYzmJDcZtjHZ3HNGvwID6ZcqJNhOKu1BkOSLPkJpsmZfKlw3jjYb5jXRODkvuQOxCH
g+/nzcGwytxH3ggloUjR5kaCkKmR5QyUccGSN2GIKqGw/D88j1I0PooIj1So6dV0UYHXHydukNkW
7Q6ymR+g/up2pnhz0HkZKdjqEXYeW8Q/WwStXebA5Elq/axIZ7k4DEoEaoQiBsLjlMRbEJuluv3a
/eNPD6r44xypxrlR10fhVSPCbR9n76Kgq9wUlfB07tLVSFHiWZkWl0Cnm1Z92XJxtvRTxa7/D9JS
Xm8sp8GycL/tEOWIDMn+qHqfqd7pUyXc63FPomAoPtkuteQ+YQmuEBeMYz+UJXh8XzeQg/tGPd1K
QAO167qQRJR6QKiNxOtfPYI6AIlk0N86ZXKqnQHZ3it698R/YAt7PKamwWeeZUdB6SzFnZ82TJfZ
KOePZhJdeCigyP00WoT+viOyERODHNvP2lX9ZoJMplKY576OA2Kyl5GuFpdP5c+KXTOU8KhfgVq2
b5Y46ArkoDoJfKtbU0+Xujd64TkoPAI8nfhDVNre250cpMy1/5iUkhGnagTZKtum7CgVFBovLbDy
OfOUyiwzlUKonFJxeoHeU7Gt4BOEAsD99NPXNCv1fVHFLktwWa3oJhyv3PJQzA5/guBt8vfAe6FY
eFEbu0n/4vEQ/I1X9bLL0ROs9s+TVcpSz4K0Dr8xIxCLhwWtQXXoJmhWTnjkxMxgE57Un9rVAQ92
MbpsWt9jQcCRRbeV0wuN4RKRywajccyUmCXhHWdNN4Lct5OYu25wl/aKVln+fC+ZhVWCO+vU06Ca
gh7TUXKgerkMY0bcs2yypRAiOy0OzHF2qEKzmajuHpzrkbQslJOgMG1ALEvOWfUsPLrhDDhZ87So
hMQsk7+0CSh/pL/Tnc/U+AP2mxYPnGpDEXl1+RyKOygrPjXJz7piOk85mZl7ErZ2yKIVsmlMTNNR
OXal8ly6cvynRCuf+KtLG+sUP9LmTWgHA68LwKpXQU0vQ9ixd1GBEXsGrUXarkgMWFhbj+TUui7H
2pleiYuNVP3ah3tI87hJ5CnVzUv2NNJLv3giMjk7UvcNEnIjzFX/BXldAOsbAHR1O+fO3qa6lxZm
NCWo1oVPRaSCqJvGo4R7XK11bjD1xwHWuSlntEGdamL6FvzNJlYa7buco3EeWpoQ2yE7tr9x+4JM
33+D3grs0KuIw361nAjDDQqk6UecEM1HKX9DKvK+Bw8hj0PX+svDOu+G1jVf8tA1aU30kcqKoX1D
YYrmBcis1N1ZSb6SpoXiYQk2I2JApUe+d2R20Zc7PSABC6dWThvTIfI7Lu8X4fNG59qVzqQ+hLjh
J/6Cltp1nQzKtaAaDPOytTGcI3dDN3ebsXizqNXIdBCDAdDaGrT5OvwGBiy91wyD0HPjubl5IkJV
wHhFYD0KrbRW3XiCvJwJkY3NYBCVcPlohhepehLoJ/5/tvbRah9yWKt6ZP+qcfwclzqBUdI4BatF
yNHOXwqxdcphxl2XbVfANQTdc2T1diyiY+JpCLLpmeb6se/izBFbHqGYOoI6JyAwFw7NLfvS/U68
hND3nxTBXX0P97pwTQkqV9amOdYgeyUjlx0gSiGwdceCY8z/109NQnB5K3u99HyzntWrK5IzBCtu
nVZC8tlD/kd6pWAWd1EAw8Wi3QOwkx9WNVqw+NjePk5o/vWlpFqbU93W7hzMkTCYPMk1PdqbtcXD
Zpx2i01m4uR2S/bHMrxgdsHyFHKgwwKSODefodCoGmBDTgwVx78U+kltzTaWVZ9d94+CcqpzawBj
/BtP9imXM6Hbgim9a7BFiKSpQcGtghFiAMOprBP6lh3zWZqzSWIQC1oPDAIH1FvHHr54BwRY1amG
Qm3cQcyEPvOQHMaSwDgsB+VxAU4auYqEiHgL+qDbiafGKEGlQGa+TNr3+FXF1nLVCGr0qSGutd+/
gFNj2IANpwDcGFq1NAvsrPAAItBJMFh+iZJ7sCbZ+jwiaShYiItQ7MR3ApXa9i0/YFAwaecUzTNe
CYZDdBv0VLYJruSg6q4ovv7GGUiRBncQWQ7b3Vw0dgE8os/m8tVTLgRSXktxT9QleazO7v+JfR7V
/BqQvRa6K5v+iqa8aWdt99HBc4yWlKEnPdxnWrTQB6YLBZWRYEAXmIDx5mtjIRy+ifCPG8XRCOj5
7UoZ5IkLdC8GRMWl9Ul6wp50OCD1JZotf7CHO75+CUmPB4NQKeUL5RPemP6kyfIhTbwQP2LkKXpD
GUhTcLCeYGRl3hLmm3DTOAnpRxtbGb7y4Z7lzhF5ZZ2FdJw9uZR17lYLTWZ694jyYtLkiFsAf6Mc
V6TvCXID9VjGhf1uCaYMG+PoW2sht/uZQFXGYpKi6nbd5kt/TqYvs35QH34QsumqAKyF1YMiYwpQ
/RgadQzIWiSM8rJauVO9tvl5t/Ro0IdAbIMXHUpJpvCMEyOUVjfvmMdQ6Y/1GNWPBApUHsVzsvuW
Y/452WnxyLr7IDnEDQZ5sdL1bBn3fBlRPZVB9zkHmw+A95hV1F08bMuTyuXwa/76ZAeFJsNvYJem
IhWQyvs+gKL9qnOf39rVcBVWWN9sR76xIh6kMMgYKN8q6mZTQC1E1VIp14qEkUBSBFmQTF6fB4AX
ID7s5jRyh6UFH0BWLKyunJxfg6kFqUilxU7VXTf6PWAqxtAQ1nqoFvFuc5QmIAHfzIvYO0d0ganL
vN+oXWWwOchhVMnBCLHd8yyhGFlhf1RXO55yZXg+B4SOspQHOt8/Eod+Lv5kixOTBBgqX8IuCrxg
b+5dp7prbHRQSj6XmZ4CsurjRglC1PnkQplLHtNKM8yanVXyGfG5EIMKzPV6sNn5KREmqtb5geui
1MX1iDy/ZzbAtP8jiO270NqyWSe9ctsMNG/iXbvPCVg20x4zz3LyDfNAdRP3VUMZrfyBkhq1UO7u
tEJmRmogFhzretQk0cWsp456rZETFjU5nZ9Spm9oLtCr0S6z5D5jUylgzuheM1RQgDK9DqAnCdFr
DHUDOG4aIVanVAiEfVtxOG4dALSXagc2muhzmD1O0ySAo0YVuTljj0eoHezBiaDr9BC2p8sXpY6q
opdAvijBhWBpIsyz+DxFKgnbFiIDwSlheJuOHgyEr0ew5El4wVf3Nfn3hdszzLT51rVIym99elUX
5kMGqW61J52xClyL39gAWhM9VagbhrKpXb73jVx7eFYmU647zdRUIJqRNW0U540q5Zmj8eMxEqV9
669SKv1mremx/uOagWwSZt4vAZda62P1kF81vdzxfwQiQQaQtScFEDOE3n+X/gbWlVPUdhFrxe5+
9H7M45wHopqmsWpjjGqLPQOPo0lIBhDUntGzVQAM4cNBR3MpHKd2z8R02I3MLDih2sZ2/Zlg9J+X
eJtomGvWkDcPIr+m4hc2XI27mK9VJrQ1mdrKEVIH+Z1SINp3Z4XVUcMyTI2p+V1niZjhYcEVvIzo
mkp1rIMF7IKzENVUdug109gAk2GHpQ2ItmAFEYS7EtCkxxc40iMkatFGvpv4GdWhD/HGzeTv99AJ
0H3wECjXZjrExFvbNs8bzw9MmgN7bwmPfvHiOzfi6ZFuCAD6ZOwjo52zexULnb72I/1Dr93TA4dZ
OmOmQ7X2g14B/jPca53mtHNHuW+/j5n2F4Rh07CIW5YTexfitIriCIEmjwa3CqHlj1s1iL9G1sKM
0sqh6O5IALzSXf+wHMAxQMZ1S1IP5CHmhnIO4A7r/2Q4+QVDCIo+8G7bz1nuBu+vu/qpw66eMlpf
p3QU0zggWT6Q4plOlLKjYa6dsYYUb/UX1FArr5vcwrXV71XgUHvybdWto95Pc0C02HLM6RDuJWDU
+/WLZM6nw2zJazTHpHgi0KjK8Zv6DDSwNt1uYaiDk1BY0qhbt95TwR6iDg2Vw3MGJWv2llkYlrDk
98kSSlPrhcmaIh5+Q8DMJfRfoHwRA3wpZ3F+XKiu5o+ixSd8ZpaJAhVNEtTmKiqyyArk44FDfB7a
/xuy5lRDX/1rWWDaZDNPR/g/x/m4xWCy01YQn3U4JKfz2Fz9eIHsxqttrXidjzFE5xiHRQvm3BE6
3j479cFDp8YOELzgqVMuM2BygP1qY/apMPNhvscGI4+I965iH/F4J2E4+QpEl4qrnawwHpCaMB4x
RK7Qw9CMbNaSukpRWpwn5a9MnA9oW7BnLMXMsyvfL1SrQcsnczRKWlfN4Aj9Yv+T/8eo0b0NKXPY
tUtau+NUXrxpmVHeJb1UMRg4NyGtHs2RQjNGClta0w63xREvr56D+XZx8MohOZnJxThMWJVgC8fv
qeG/Vbr1C0rLoUY=
`protect end_protected
