��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���8�'+ M�ҙjb3P�Ҍ<���Y�a�~O��2��Fԗm�!s�E�81��IO�s�y�Mfoo*k?#i�I��6����[�bq.ڳl�n]�$�����k�'z�ydL�-0A��4���S�0�S9�� ��K�É�p$W1-��|�/%��P$j��1��-��P9�Z�]�C?�R�ч����������a �%� �Ԇ�{oBB�L�/�b��Դ���/��;��^��[�k�w'm%p�u�q�R���@a�8����3�q��,?'xY�00i!P��1]�?�v���$^ש�A���l��a�;ɔ��5O=��A\
f�"�&��~<�-�I�a�Uw�&^ӻp�9���ܑ����\}&��,٣�v��h���v+�F�7f�����7��I:.���g]���a�54�甴Z %m�� DR�sP��^�{a��<��H	*6��tB�
��yHG%�6�/�ib��ۢ�a��^�*tgh
ߧ{�����f���yBo�FZ���m��h$"�;4�H@����_L `����~�����W�o/'G�n�<Ż-� ��K�):�����ea�߹�[�(��ԏ�厼��|�o�O���e'��x���f�?9 ̬U�a�|��3�x�~Zʾ
ƌ�<X@E�����w?�V�X`V��yez����s9�&�ն���Ȏ�빺�F���(Z�²<�rd��MKj7�NG�,��d��80T�i��1�n�t�Y#+�Պ����~��gUP|^�2�tZ�_h)'�� �t�t\�A}결���{CEv3��gX\8:|�Jҥ��M���+ �@�k>���\��G������7�/�Y,��H�7��ߍIB��.�p�H�*��F�w,D�B/�9Z��誧����OJ9$��w��A&�w(��O�1�~Ymخ���akAg=��p���X�Ԇ)G�n��?(��+@�q��_w��GQv}^�{��HCH��r5�.���DX]gX�l/u��5�(B)�ԋ\
Ć3ؙ���$zH��n;)�_�q>5����!C=�h�A�۠�ck[���l�Y��.Je~��I�5��s	��y	GcJ3?��5:Is�����Ǧ$�����\�Y�BO�+?���-���M�51f@ �/^�������'�h���}�t�Pr/��ңy��ϞwT����=��C�8o�i&�)�8	+dQBM4P!f>��Z]��S���%��.����΢?(�pCm8L�0��{�`��7l�q��ީi�P��|'A��*fH�㵵
D�%�n��uf��|��g��a�;`R�؅�^f�@�&]HBki���7��
ҷ���>��V	ԓ%9|�P|��4a2�L��gE�8<��\ڿ��ྚ��J�A���L^yF�.�)�ݮ[�%.�}�(ꍚ���gm.�A.l)�`���z<N�Q��3�V��nQ�x��p���I~��嶢�NΨ�/�Rb�p�8QfQl�	޷&`	b��?�X����Z�e��j�Hhj.�T{V�����)t<�HPO�A*̎�oS�Ţ�y#�P�1�|-8xT���;bM�q+b�4������"�Ry�+.�����O$�yp;3�;�B�����0���
������Gvz�,Y಺�"��"���3sOĈ�-���w�Y�(��w�|"�w�1�r��V��.E'�c	��I$��3?u��z��w�AS8�*��,�05���ı�x�T���S��##�G��K~��NJ��/��&���U�͖��VJh�$�Na�5%�����M؜�$��!<<���5��&���ȕB�<����i�Q2� 	���+`�(���/}��~3N�uR��>v=o�0�	�4wW��7kZ�Uut%�v�A �����6�O+����uޗLzX|�)�E��.7�mO�S���Y(VV����wr�a�zNE�Z�X(>���b2�G�0/��[̖�-p���ߩm�Y�z��5��*ť��|wD�U�� ��	
ē;p6\����2��ѓ�̋��e*%��з�xWaH�u��~��}�o_���w����"�2H� @�[#+�9���*�5ѩ���x��=����qp��h8뽰J��l��(���g4"�"__����E�y$.��~�7�/��k���W�4A���`��xJ���:��RR��P��ǈ��=�\uZ:5l�+��c�q��,�f���ۣ��=1�DJ��Y�R4W-k4e�0�5E2\�q�-_�y**cA�.�8��qQ�͇n����m�@�D|�|��x�������*e�0��-�:���fL0��1Ʊ_��m�"T-X�Sp~kp�)K�p=?O���1�@�}Ll�R�SR�?��]��r��H߃���r��\(Q�����d�R�t�i���8���TU�'"�궜H��I
�����f1]C������GD"r�O��S���䇽8�Z���:���D8�`q N��v{G���;n�r�憎$TĀ�Y=���=Hs�����fO~��?d�SS��Ȃ=ף��7B9�e�nI������M���X���@:���o���x�E��	*I�u��(��>uR��g�ʗ�ĵ[�.v)*����$�%9�$����IǴ)V��¼��z��x��$u�1'm���������%kPz����c D�T^��>6NU7���ԡJ�}jg���$���/�J���_j�_�y3�Lok7W)��g��C���j�D]H���vf�s!��4f���grJG<m������! 5�K���J��F��u��3����XTx{�qA���g�^� su}��k��5��CS��;7��.5�5~F�Q���h�HD]� ��J�H�"�Kپ��4!�k�.�e�?G���Z7}�Q�c��f7@ۍ��vIqa��0�7זb��#1Z���/b �d`m��6H?���5?�$�3+�^�j��P��Ц��^��9ʗ��g-`���s#����Mp$M��۸�?��97���ƹ>�{t��F�ƾ�~=Q���d������s"��#W!�ۣP�֝�<��֫W� ~�f��gn�������S%OP 3LW�DP^ ��;��j5�S�n6��S��:��&���.�t��?ܷH�������6�h���'���T<�`�Mg��,��q�I�'��l�������)Fߺ�]Lo�B��j�RQ��˲z��=Ed���yg�n�����)c�8�t��	_���;%oׂ������9}s��^��D�X"��Y
��XQ��˶��S�
�{@�Ģ^��B���u��a	��@
�]+���9X�<�A���^	�m�t��T�<�9�O��:������u��'���O�~ŕ��)�����kHWh�&�g�0!�cF4�I?�Qg�v5+X���Lf�<ͽH����g�����o�u�#�}���v)䌑��_S���$fe/���b�윪����/����}��y?��G�+��
�tE21����8;?u} 껎(��_�>����#��Waf��/�L�/aP�)o�Җ�Bq��c6�dM��3��#o���O�Q��U�������)����b�?��>���йwx�ܪP~�A�W���E!��n����b_�eOzҺ����g{���c��x8���P��Qt�s��a�,֘Ç��`�(�{�mr_���y/���?YX2je��{ȍE+��Hz�fZ�X��g���o��.��}K#Kr���d�P<Nf����=֜�'���,{*]�1?�uO�{{ڗq�|���~C���g�h�5���ҤG<���sŹ2Of��7�ą~��E�>?��5q&��Vⓝ�8.l�K���Z��(!(Y�o�{Sb�����
���uJI$%�܎2�u�w������W�9��@�2�Ҽ�2��n?�� йdE{X�O#C�p�ZÀ��{N�-�����V�����w�%��5n3���7���
��w�����T WFE(~��%�UL��E}]�#tnԲh�-������]����j�_m5M�`�g��q�Ue��nBm����}p8�Gܓ�8��' a�5b�cU�fBL���z������≇�ԇ܍��2g|��ʆ�Ў f�J7��p��p����)M1���vs �����䷂|2�� K�vO�DSS�o�?V~bZ�_�A�@���۪N��ˊ��T\�f!\�&���@s'�6D�����CV���M"�X��&[ 0�6��=ɿ�G�Y\��j&�։j	��<
�j�f_A #����CwO�V7'�5�=(��I����T�����G�.՗N@����_��z:�� c{�j˒0���Vƿ+�H��%��]`�!u^�g�>���`�n�9`_�ai�hn��?
r��&��V�����=�����2������8�,Q�3��W���@���'��	m�~gT��H�P�
���X��C.��N"$i�v�6���^3�0���:�pk�gx��(�
�3v1w�¬]f8f�F�fF�b
�s���fB�ͻ��qtSO������� ׿"-�oFõ)ǭK?�^?{)�� �08,󟫈s�7��9���l.�ȨO��Hf�uv�4ǁ�~[���ǃ���c�%#.��I'ߴph���6��c}�
ß���r*����h����L�Ϭ��ɻ�J>84�ӄ]�́�)���U�=��/A����̰T�(�c�=�a6�l�A�#���Q�r�kd��qH�bU�s�Z��ɣg�[	���i@J8Ua*.
D/5r]��;+F�D�w�4 u����~CK,B��xTV�R���:�݈��).Z����JB�{	WJAA�A��-��Ha�m����!�^^��r�z�{ ��j4u�O`6��ޅ�J�Q8Í1��k��I��]��= 3c�HDET�o���5c��z�ZZ� .�_d)�ʽxu����;d?HJ,��Ӗ2l��W�ai  �0BjiX	��~�-�!�Xh��5��0�!��}���l *tYK�ֺq�ʪ`JZ^Z��.����e��ߎ�k}JӨu�>�>m2@Fi>��꣬�r��ͼ��C�%�L6�7�rdB0
��֕}4_v�Qԝ.�X<`� 
7>V��͈��ϴ�"f�6���ܭ�_͵Y%ዮ����kؿg\�,�}�����c�D�/g��A����i-+vS��3����n;,��6�58%��9��!l�7�ꐻ���Qq緵 ���\K:Ii�C��s_.N�sp���'M_�S����y;�d��<��%Ҿņ�e����<<	B��N�&��HxT�?Ze��0G�;��6:6��#����*U6��������F
.�n����#j'�\�){ɏXmsF¤i��](M���N(S�k��Pa��2_�س�;�ﷀ=X�&	t�R�8d$W~L�&'�I� �E>��M�4�د��Ͻ�T�K��0[�jф���?a��u8X�8�ݗ����˫��^�BF���E���e�9��iP���)ow��^v$�D%��$�'�z��,~���oC�a���x�j�a��H(��r���h�L�|���Rp^��O�@5�5/�$�'�W�V;��M�̙����n�����+z߿_	�L������wM��V{���5��s[i�z/����R��S�o�~��ڥ�.��"���,�%�ův�u�l|��-@.�ΰ�!bw���p�_竬�ő�%,l���?U�	�s���#�pJ�A��	�F�=�r<Gs��CM�C�2?��&��ճzR�'���iÇ�8L�a��+��bqe�`#�**T��J�C%��x�� �����|~��rv�T������Gt�p�_�v_���cO"�ߵ��9�AL��4�Z[/)�����+�;���9��QӚ���)� ��.�J�Z)U�O8�O�^�g�.�b�v����'�^/3IR%3ҷA]�wf�d;y)eX�ѹq�ۿ������9�ra �]�6��m��;oc��Z̠'�����~��[��)�ԉ��+&Nw��u���L��6��Sܨ�S��h�--�A�|��=B�z�o�)2w�~�Pt�?��,&'	�������,7Dͭ��]���<����T�?oVnP���vĦɰKB���]�r����l�8[}��P�&�f�h�_'F.�NT��yS@F�_�	������/�%�
�KǗ�g|n��I�Ghv�#D!�:lC�(0��@ _=�@R1��Zʎ�t�W)��1y�'o� ����߮f_��<KE�3�%@�d;0�6unP]^
�m��cx7��A�
�]H(�T���c~��|��h.ş!:�Yb�ڛ w�gi�u��s�x�;S�R٭�Ɇ�P�E̦�E�ӿ���4��D����p6+��j�rt�4kܡ��2\��E1�L&�+D�L��'�.��   )r��"dϾ��^�%���\Ǘ_hEWb�=�Cf
����G�[�m~�X���{M;�F����g�z,�`����* {�9ܪ�-���T��b46�c�]&kZǉV�2
Ԏ�xaI
l��X/D��ʉ���u�VM#-M`T�p��|1�7��/��2�{���]4ɗVt)drY�I_��Bp�j0��E6.�ƫ��j��z:.�o��)���KYp�w��Y����ZdXH��a�Kj���"V�B�gN{��R'�����_e.󮻏 ��F{me�
��@��]r�<���	@l����ѽ%K3T��1��.�Ⱥ�p�r�#X�p�X�פ	�hqz��Y�c���1��?��Q���V�?��E��� �ع����f���MT��!0��!Ry�k���3(^��Dއ�c�)�ٳ�f8L$1k�]�GZ�L�m�����YHW)�m^��4��;���1�������I[����1W�V�<Å��aF�ڌ��k�a�2w6
$�^�6��^�e��(��Il���"��q*c�/��8d��G��`m:]������e�+P��_xh��M���hW��st�tH�­k�S���bWpt�bl�9�
���c+Ş���%w`�wI��X��Pb��Ri������q�";�w��OO�i4Z�P���/�P9z?��/2x�v5���ǘ
���o�e� 3�*oP�?8��B@���}����5��B�y��՝�4M�dڥǒ�'�a�#Mv���TT������e���-G�JV�X�w�"n��{�Z?A$��,��M�(!�
�e��#���-.qr�=���Rrf&��{��ˈ+��o� f2�s���E!ߍ��ى1�D�zYHA>yb�uD����]�1U4~���5"xp��$����Ə��6�4�;�k^Xn�����3��}���,V�/ab4���7�M�����K�^�`��k�=� ��S}r��[o�6�T\��s*�ˣ���[��.��YΫ��K
�5��6�6e"VXBU��l�LEztV��B
��.V%�i�`�z�Rt�c���� ��� �g4c��٥';�D���P��Frjt-��Ma�a�Ư�0T��@V^��#L�Iܭ�0�ε������[����"�?H#l}�ӣA6�E���*���>���_��箰�d>�&���g�8����n&���GA��Z��Kd<2u[�:�t�	��!�'S�UÍ>{r�]�����Qm�z�*�S�/�ᛴC��CC�k��
��N�7}��ޒ��,H�hN �C�/Z�66�KT<��3�����U�R�B�4�E_����o!����8IȊ�.��FMx��b����ry��@�.l��;��WE���)߱�ju������ԗ���[�0A�j�`�ⶳ9j��L����<=wV
��B<9�-ns����!݋������w�eue�M����^.�okt�J6�sĔ��EK�h=��L�$� r�����_Ӽ��4��2A�,������F�J��K80�>����#$������B8녁�u��4I'Ȭ��Ϗꪈ�X$s�͝#o�a�Do?#�	F���V^�lI����z~�vp�z�[s�J��")�5��.6���?����9,��/R�V>(�RC�gܻ�t��z3s2V��O
�
�W���T�u��L#Z�j!y~�6�ŗ'~�Uw4��l��n;UX���������B�+E�9��>�1���o�HkK�@Ex�1eɰ\R@�Q�k��f.B�Il�b�4OP�y��I~/~����f)n�
�&�������m3/��H�<Ykz��㞠����^�l���G��b9Ṗ^V�}�a�TnR9�в�a�w+Ro��)ĮF��H�m�2=晸*�!���cإ�_,4�jX!�o�<ɺ��)�e6���� �r�*��.*�)��3h�J.��Ud�k��噷�cU#���<ˣũo����[�S>=9h�' �2�EMq��ux��P�u?)*O���w"��C��!�Q����&N^�UYf�C�$3'�/8�9�$�n�<�'�����Zؐ��1�L�����������Mŉ�%�]�H�
�^%����7d��hy�E�7�٨���b}.bź��l�w���Ґ��߀�����"�+ݓMJ�9�����	�]5���_��Q�?�>2�L��y�ză���ob�}ib~��Z����iq}�#��!S4Qb�8y9�|E@Cځ��{G#����Ɓa
,X3����9K������d� UKxJ^?l�'j0s��1��-�,)j�KDN�����r.�F��d(�\$�n��	F�F���ׄY�ߍY�� �w=��E9�t�!�=̄�!�>T]��3��4=��'v*r�g�ϖGGQf֚�4�7PO9���a~�ຬ{Hts�QAC{����(׶i�e&�x�6��!���q�Y� �K�6�7[��%vyZ\&!�W����|>�k�:��ΰfp���F�	�;`��)r}��46i��"(��.�Z4Ν���������|� ����a�g��5A�S�C�p���s=$�X1K�[n���D!�茬�D�Rл��E�^����DnmZ~(xp�Jj�C�/᷹Y����=+G�Qínഒ�]��s�/Y_�^��c�B�;�d��:�+����~�P��/K�:��ct�z�5�Q��T���h��E�r��vP�v$o%~��ې\��[�W�zfdY�E锕��x�����b��P(Ky~{I8۩""�p�Z���B���������|�G��Y�@[�!N�LDL���m�4�&|%KѲ+B�$��|b�\u�^tT���[�aه��!�ez�XD��
۽S�I�Α��,�V��-K�]���!���Gi��}<��CH$��<�}�9�mC�b����vg(8�y��-���/|�\�+z�OIL��?��e[���U#�E�d��kX�ގz�t���{�SK����?"v����]��\�e'´�o4_!-�l�B���u���f��~
�W����'%�*�R[&�Z������ф��ؑ��Dq%�?�f����L�o��?�b�$�]̄G�7���/["=�_P���n�k��œH�
�z���h���۴�+�Kp��)h��I���A}^�2+��F�ҟq��J�Z �S޸#����bw�H�L�2K[�S��'�4lg/�{=J>�O��x����`��o��m ��-ȦLK���5����Q)������%�=�4������� ͞��4��6�9b:|�k#5bIJ �t~�)%�#鬈V�e��$�xiW�[�&G��/l}�v�[�����)���{��v��:���H��Q9YBx[�Z3*�\p	���N�o��������?��?��V�m����"�E�fU=�f)Z��@��0��o6�~��0p��t�{���xA�	��esȳǞ�=l��4��wxM}����
�^�慇`)��"x��g�ʢ�h�YH�}%�SF�$�V��ꌿF��U�E栥�K�1�����r=z��	1~Rւ��kNt��X?�Zq��f��g#`�*
������r�c����Z�͢���ځ.h �e<��'��%���b�������˝Nk���.�ԛ�TL���3�Cz3��f�����lO�4Yg2�<A[Sw{Y]��U ǣ�����g�GEv�
0�1��ߵc]ɔ�33�7.=��8����`�t�ȬF/�8qk�7�/z��dVaj ;'|D��ز�p	v��A�*�Qf��{�����äך\�\0��^Kz4<�UxY�e�����LF����/���Z��ܑ���*1�0D�}-?����C�z�z���S��a���C���7aXޓ�%iN�·�oj_Md`Ry�Ys(7��i�?�Yq��!����n�h�^1��S{L��a�p����(�
�����W�d��H�@d������)M.8������-"�e�?�q��u�����'X&m�9�����2U���%GE��/M겵���ƏT]�ki��_ֺ��� dX��꜌��T��6���f����c�'����2��6?�H��y�~��)�&�Na��A��v�6lfV���ZC�Jg�����\(��3n����T��;�{���_�&6"r�G���h$r�)��.D�������(����X���Lը�2&m�#�t�(^�|�C�����;MNG'xT�$ �a�1�v�X5>�$V	M-w'��Ur��s8E�S)-G�["
�N7��rl$n�1I0����uVm��7�}�d��7jQc���1A/Dd����p>qT3�^��O��<�
��"����V������|j�_�&�^:�H�KDp"uN%&��U�7gk���' s�g�YG��u��nm[d�@-C�~���7�*ӹ��₲ĺ��p�wL-�?����ԕ���4���/L�?ڮJ]�)O�!x���o6�V5K���*M�miN�m�=Y�I�q'�n�T�'��0��,%tM�T�����-��}���x�eP4֧�
���1I�Ձ�&��SP:�3�䠔k$I���h#XةrK+��i*q��y@#���I��Qs&^���!�n,�����^Q\����\7�l�6�9� ����L%����9#q�r����v��'wH�d��rBJ�O;�༘�M(�X��s�\4�*����&wa�-F��>b��v�����q�5y�2�J
����������ۍA��Voix!���~
�ԃ�bw����p=Q���mY���𚻮�����gb�i[�O��<%=�`ɨR�|�>v�)ª���Lf\ǃl��.�JE%�ݯ��>@��c�E���T�|h�96ic,,X�k�ں�j�w�bλ��LY:�/IY�zhub��\��J-Q��ո������!y�6I+��o�v:��֚�YO��w|7�*\��	ʓ�QU= A����Tks�SNVDT��6Q���!�$Y$����p������u�,~m���M%��X����.�G��T��2e?�/�ᣑ�A�9��Ũ���z��'�/փ���"���́�
X����{(-�8�e/uN����%U��'��~P*_���A�<�k�6��v�x�[g@���rEZ�{ ��x�����s���l#0�h&��𚵽�r�5��+VKϘ�v�7���t�FW�|���E�����5qa�V3�傅z�L���p�yA��1�lh>z�m�c�Vŭ��˩�gy�e����Su��	q��]�	�#��mG���|�ܔRʢ���Ԧ��zS��g�PX��Y��bىc�E��{����q���Z]����B;$!�}Sn��Ã��u��Z��;��=F�N�G�	=|��?t���>h%�/$�穲b�H�!��&����&�Y��{��*
E0G���A�d�����${�C��� �VM�NjGsQ[�Ԧn���*c.�X�����/�����=w�tv\ y�w�\k��G��"1H\1���Q<"�f�XJ٪2�32��j��B�y��a�#Aaf���k ��/H*��d-oK����O��A�9����^9E��?��aq��!H+�\j��Y��>U%?>�	�*e�{`E7�L�{�EU[�@�U=�?�����h�OczD���CR�.a>�ć����Ġ��5���ƕZ�|�+����X�e��s)�͗�%�	kg������mG�*���Z;H�|/�d��aє�$�K�(	s
�.y30^ˏ&)�@Գ1�� ��;r�4]JA l��nw2�8��"\~�k7�b1A�Zb�������&�������~�kr�|g�3Jۑ�R�U-e�Cǧʩ*LU�ӥ ���%�k��&/)IR�����{}�|�\�~!��{0��.�"��/I��K`Kh�\��%f(��'Eh���l���Ę�%ޓu: ̽v��o��V2AA@����Jx���1��V��,dl�Bf��>o��S�<�N����WǮ����ʲ᎒7!cT|dWS� Ž4��ذ����hm�OM�/����`��b?��>+�_�J�G�F�8 uu��������cH/]!�o�uM��J+e�
ya-�j|�:��͕b��X;�쬌}Mc"+����D�CȈ�߶���3���`ȏ�U>�������������+�����͸!؋�.�[�-T�f���%�l&�31=9����NeAd��3�!K���\{g_���N�s�f�݈���z:����M�X�z�ga8|rTIJ|@��J�t+��`!���a��l��ϱm"FP���臸���y�9LYZ�d��mg�Cyi�t\�ɫ���Z�MAz��V�H��m��?U���ȹFF��TթU�#\5�cŔB�ބ1��0ԟ�cj�ar��4Ô�j%�a���2ʴ`��p�
�j�Kr���k����\�|�v��sjX6��
z���6���g>F�,M��f���#ڝ��!��S����`�I�{
�~�7��k�9�Uj�\R��	Dk�Kv��ݹ{�o��yy�A*j���joa��@���M��R�*����'����ŋ@�O�e�W"�FH�mxn�b#�q��s��6�|@D6�"�RQ��&B��Cɞj�	gEUVSӿ���ʏ�f:��2�B�/��#a��l�i��o ��M,z�;a}Fk:޳���f�G�����c���Q��u�"#�S@�G���'�E��]:��Lr���a�=�w�/!��z����5;64�1lH� >Uܼ�$�����"c����j��7uE���,�(����o��
�w���I ��ky�����8�^kI?�lջ6H� h��c�e�zw�QLaD)��M�_o���=��k����Kz9��:S�֩0��,�jf�Y-c�\7���bG#�KnE��c�)pȠ��3��5�XG������o5�"I��~�CG1e������@�1G��3yiu�t��]����)3Gڪ����+�����\紁����:�bX�5�-�IWݭhk�RN*�����@�r���Σ��v�ӯ-��+o�7d<���Y�d צ�x� ?�?�5 !�%��-N4������5�d�(m�a��I���ҹ�?\�����י�G�t�7��g�m	<��!�	�L�����a�䡧O����&:B���&t�ׯ��V�B��D*)�e��>` �e��n�7Qk�	�� "YD�m	��;�/ft��9_���]/\��,vmi>��9�"at)���`O.؍�?GK D���8����#��{��'a�1�#�&a&�z~^�#a���8�&�'8����6&σ�l��ޙ���g���[���z���1k+fl��:��;ښ�YH-�ц3;aN�J�ӯ$X�y-�m-��xe�{���� 뽐���KF꼑���1̵�͸����oO���WN��S�
��rƕ��\~��-faF.r��.<AR^U��_f]ģ��?ĥM	o2�s�\v"n�N��P��O�H/�1���a��[�
[VL���.�%��+wC��:�N����XU�ћhڨ[K�0V<�֝w5�������D�Thj����`G���(�E"d"�ɦ���,����?���-s�]T`45i�U����}Y�bV�Qe���":�Z���	�K�Z�[af
��D��������fd�!��R7L��L ��������0/��dC����<ГN�ca����La�>˫�ǟ�b���Fr	>�o�s��G"�.�&-L=�3d������$�z����ʹ57-(e��}i���K؋���ə���<h������Ü-B�7뽲��r.z���|�["F�����9�h�7���A��P�M�웈_:rx�<�g�����A[ȡ�j��_]�k�R}���La��;�3����ƨj�̞#fv:���s��'d��Ǡknz6+|w����N#�ӊ�5���G��gYQ8�|z���RR�R��I��[vL��A���Ce +t��eͤ*���n*B~���q0>R�N؅��զ���x�F�S,��f�:�� _��Џd��rj٪$�iσ*���W�㖞�P�=��|�M�f�$�:zH��zWXN���3�ձn������n��MN���p�R��8���H\Isx����۹E����ۖF�W�����ء�����B�"����nTxa<�� ����f���	sŝ4tF���}ΰ>�t�OD_�H��d�H,�����w��X��%J�$:4!vA
E :�O��I�E`3�&W� J&��\WX#�9���/�|��C�Ưd,���n��2�w nx�9��d+Mm-,�B���᱉��BT�+�(��<i�8�9Q����(Q������#�`����O���$+fy��J���p���!���$?��)��a'G��7��^��z�	�{ ӡ�{T��l����S�t	��V�j��R7;c������g�s7P��ߪ(���6(�M_?!��~든�Hl�u����`���a]l��� ��y��3&�p�\aR�S/Ѯ_J=�*��\ՖtB�@E(�}.#}$>�ڟg��,����Eth�S�G�Y`����/�y_�w��7��@���m���V�\
��g�`����瘤��~�-Y�w��<��e���f@;gr ���*\�{��-V��3� �+�p۞��!�)b~/|� ϶]�����2���BT��ol�Pg�4F|N��_���*�E�x#�&\#%�?��3+x������_����<����_�`)L.��nݔrK=�
�0��!~��U���-؅��ORj!Քg�"��*��NO��/q"3>���U�ۼ�5�S,㛍F&��8n��"�n�gd ?��K��>�E��s{)� �;�^��G�+�O�v��.6��]+�+��ǃZRְs���i7NC%�o$���u��z�;+W�<O	6��|8�ҢWBp����xW�eG�I�d�Kׇ�A������bEף�pp\�F�k�]����*�G�K�j�� �.ٵg�V�q^)��D�"�x��w)���!�	�n��zoi�T�-bU*�s'F�����VgqH	kf>�р�
o};�#��"�,.�\Cº�����Y-rQ,3���i���]����N��0�?� �7����S٠����Sv`�'�O���uF��\�hќ��/3U �2��q�ke<��䎯}h������5��!za�WbRj�Б�-;;
QCK��������M�-`�۽���瘒��R|S3,y�k,���v�����x&k�����#D��I�S~'c�̫�}
���X?��M?%��@
�T�1P��~��Q9���-�$x١�1�g%�s�~�@�|Iz��)A�y�x�B�p`C����I!p�=��d��>Y�尯�KW5�syϡ�Y/+Of��Z��u�~+�&<�w�M
�#Ew��͓I�����d�g�!|��@�JYՔ��j��#tû0�Ϳ?qӾN+�H�
;�K�-K�HA�4������&��;P��x�� -��;9y6�^e�)�sfiq#�����G���13<�#6x*s����� �ӗ.�1T������_\']Y���\˱8�%I$�����t�oFŗ���"w���S�	t�����*��@>[����-���`(��3��<�@w��'-z��I��O�����p�����n�p(L�5cҸ����2[!R^���5��F3�5�]�N��B\`�H�"����dqU'���7���M%@A�a�14�J�ݞ]X�^�>U\��������9�'|�Sַ6�/���l	pc�Q�;*XQD�N�F�&�G���������Q<a�Q�W�������ldi��)��y$=S��C@�	*r��(~��/nxB��*�nn��(g���/~|��+g�!����&Va'����(ޭ�� �ܵ�o�*�R;H4,(�M]s0;�\��6��y>��A �(X����p����4f���P]qA 5��%Ϊ����kEH�B��~2�ch���G�X}����4>����"�5Q)?n�8�p���T���8��
,ġ*��q�m�1��ڒK!:��	{�����J���Z`��ź�\�+v�k�]�����ݎ��1m�?<���2�����o��a8m���h&;�+0�iE,�"[/鶲踼	#���e�@h�㕇�`$�۳�3��S.��'��&A�� #�u�t=U�#Le�#�u�Ӓ�z�u��Ŋ�K����-П�_h�0�wW���3N�ݗ-����|7�̰�/��g�g���̡Ȅ�O�G�6Z�
Z���~���Z��<a�X>�fj���QqR[R���f�9W�N=�&�lTo�h�i"�
��REAQ;�e�h�Kfh�0.�z�=��5g8�H94��߁��wdFs|Hzz({�Q��ik$���4��8��0 =�N�zD����*��QU�x�h�ܿ��p�~K���I�Ƞ�eo�-FظJ¸t#4&dO]�㗚�A/�B�S���-eWߦC����k���[��SG[x����Ep]qE��ǶS�\���,�1ӝh[u�N�akg�Z�X�*J�R�3-K�w���f���c[��)
�&��ϲ�"n/����/߃,��*'�-s���lZ-���VF�L:�-�+��-���  M��9��m^��·?גu����=����)䶀ڈ,q���߳O�ϧG�R���3kX���(�#�Ti�Ws�w�_�O��lW��w��[�:����	*�p�j%����\��4�dlx�=��-_r>-p��3��ur�t����Ψ\��;�7'&�k���9�t>6�OvTX��V��~&ñ�5Y��Ѯ��G�H�ZL�>.��	�}|����������?����A}�Q�#�k*�7:��g����J؜:$�=��I%r�2q�i�H��Q�(��G�l2��u�w��Zv4o�V�i�V^��.�����ZB��s� �2H5b+�̓zfY�~�{��������W꧿x�;�2|��8��*� ��1 .�./�x.�H���v܃�(6R��J�}��fGi���"g�����`g��^`�Oe�؇����u44�:���<�d�?����?�w,�ңm�5+�l����U���y8^c��4 G�_}$��srEr��j�i���x��}$�w��v)ߝ斵��m�O����Dlo���d8W��@�G-�s�T���#�[��e8A��1�;�B��z�1FR���/���zr�^�����HFmdeQQI�|�������l�p����Nc�+�,���7��b����Z>�=Eg��e��i��N1��H����&}��;m��bd�n��}M�SM��f.֘t�OL�o�J�-0�do�۲�L�%��֢�2����r��,+&7:L�RVT>����B��CR�%cѲ��x�@o��-�q��)��Z;�?X�FyN�, !�ŗ=fZ^>���L�6��ص�~����W��Ng?`�5Os0��S3��ъ�9�E��g�#���KP����i��w^�G��;�o�0��ЕԶD�V�	"Îfo��s�%���#�w�pm���|�\�ն�x���E9�p����i2q.� /��������k|����u�N�)¸��a�j�>r~`��x,^����G�w�YN6�0����\ڃ�����k��{ �Wtg����
�*��7"�|qHt�B��5Q۳�f3���?_�HO6f�7 -��`v�#W�I�W�6T��7zH�#���E~IV�GZ��䛈����ߤ?�<Ƿ~t�K�	����)�N�HI�Z��\-A_6���p�߇�� #�/y?���o��%qJv�l��ppD;<�3�����C� �!��<��;I�!B��r.�@~�:����Mhu���'�(����9����ZL���[ɏW���Ǜ
ضt��KY�t�'��a���¦	��k$Bp�'�φʘ+0��g�ɓ���.��MA��O�4�T�t���5���B�[�!-�ʇ�,K�U�?A�w����w��h���!w&�����9l"�%P�#����"O���"����}�?<畍�.��	T���� >:�Ėyz�S�#��.((M��=Q����pS�t�����%�l����2V���G@MΠ͠\Eg���epF`�:\��6��w�1Ϫ���w�x4.Su`�qf�;`"d�B+�z卛&��ZX�K�-���w�5qg����pՎ��!��1<]#��'yw��nMK_+F�x`���E�\���?�-�Z��c`7��y/tM�����Y�]��.*�4�"PXy��R?�V96�n��J��7��K=�]\:ΐǩ�1Y_���m��>�iK�ϩ���fhœ�G�� I��t<��ywk@nȱ���V�]c�b-㒥��N����x9@��A����u ̿�3E�<]13BrC�A�!A<I��s�%��@��Oﵟ�n��g��~N�PG��s��oOv�_=ܯ����T����_���iɑY�ǀ�t�~�����4{���6y���O6���O���8���z1T��L/�Wf����xE
��obl^���� nd|�K1C�}��U��C�$32`̇ܤKa�x�I���,aN�{�j��U2sc�����`)��9`�đ�v�@��e�y,m���?/�d#��}F>���GT��Uۜ�@ F��k��}�����h^>J��rr?�D��V�:�� �@,h�گD?B�УQR*ü��Is��P�Un#Ϛg!��|`�/���`{�(�Z�[1a�7f�FP(L��$�e�9+8��5���sux�����S�P�R��pv�
��r�4_[�%��u�~N�$�_iT��x��XAx��`�T�ccvW�v�/)"�!�v��x���<�[�0!��Ǿ5�uM��L=b{X¢�S2�Bd��c�C�Jd�/�GZ�^!�L]�9Q]������_�Q����R��\/�y}M��y�,Q<A"`A���\�H��6��
{�4�212��_��~���/M'e2&��i�e&5�w�NXmV1���Დ�R�]DV��ML�%��nYê�� ė��4:ʍa�� ̊}���T���k4�&s����
��
�O3;��AN#��PRK�@�nF�B���@՚ܳ�`�<u>�k����c9Xnc�tD@t�T�`H��MEk����$V��R����u�~��i�J�!9�����A�X^��q�n~�ZZ��"�L��ģ�RFy�\�	̼� ����`}�ܺ�\k�g0����t��=�1N"xy�+	�O9��\���,|m�5�ai�X�he1� �ƚ$/t���n�T�y����N��YV,���'ǡ� AlD�/�ϼ�p�^��iP�7���O����f/S�ؠ�~7D�D���.A��}�^[��ظP�l;�ْ����KaۀZBS@��˖�8/W�HAC�w����~Ꮷ����2�����y�H��[������#b�a[�D�w�7I��%�ő�W-u�d?eL>@N�+<�&����\�+��fK��$%Eۇ`���N��F����3��d�eWwo��Ԛ�e׸��Ŧ |2�r �8�ƧCb��1�� B��0�����h�(7q/�}j�.E� g����M�%�"�^�7��<�D:PWI7�1�>���+�ꯅ��^▜z����!f��s�\VHn[0��P����2���rX,ʾ���r���,hHjC�X6�b�[��N2�)�qQ����7/��qq<��Scމ���b����R2�<PVq>	F�$���g�@����!�^ĸہ��F(�v�4Cy�,�ʰ�\K��YH���<=�����df /H\vgV�ħ�/_=f3��AI�ܳ-��o8C��a�=��j��B
��G�s`��!���z�W��s���/vV>�`Y@O6��[@�w@R�,,��	�J��xkY���G���p��к�o�3��m��ӛ��ǟ��͇��1�A��G�A�l7���e�V�h�)�5�&��l3�hdǭ�Bg�|4PA����c��/K���^�gX5��;l� mt�D��k���sZ��8��bo/첵�e~��j����0-%������fl�X~X�G!�Q�A�@ڽ�J��2~C��ai�J~��u#Z��>���Ţ���C�v@�A5�	
�8�?Ft���j�zJ�^��_�ޝ:�NA� �N�ef���|�,�Ο����g���L�Ծfb&J�y(�F�i7[b;�)O����*�V<��=��6V9l��i���J���A����~��w�H�U~ѹ
IQ_UF�XY��Y���� ��[�U�V^@k�F���b3ӓ��[��2!�Dױ�5�1�
u���0 ��C�p�pU6�y�Qƛ���%�J�F�?����~{
�+����x4�J��h�>\d
Δt=�[�b���/ұŇ�����]��:m�q09��l/��@r�.J�|������q�{�����|a'���B���E���< �qw�o7�����"3��	S�6���^-D�ճ�(WV7��T|�!T����W� ��i�:�rZ�=��}{���XUGߣT�q��֢i�x�!�ܸS&��KF�c!�S����S2��M��a��> �VFC�抃Qw�NeU� 5Ћڊ�rAnc�D
4�jt�P�'�P��esx��<��BJد���FNX�qjPD;!�j�9�:�X�/[�9�U�3&�lC`�/�H5�+r�&Հ�oM�N��u�
�.vU]͎�~4c F�}��8����<ٲ3��p�01�	R�վ����'�Jɳ�F���o���S�!
7��
��}hN�ŏ��S�W�\��fX(��J��M~��]Y5"��B+�������Z?%�4�����e7��?�^�V�|�Yt�/�	������1y2b$�7hH]w=o�thZ��5�:�*ǔ��������/FZf1)�ؼ�U�O��)���I��p#|-ז����d�<�c}�����3�)�E�u�b��|%u�7/�R��}Ȗ(�MU�;�����~��M����m"���?��j]�S>�R22��K���+�X�ä�_��R\Jc��w�=%��Yp�[�$=���Ȳ>�Zu�S�#9�{��(�1r�0z����涱�*c�F�e���щqF/	쫉m̫(c��!xԥ�kf��6�r����8�Ʃ[w���T&m����y�"u��0y�*㾗xl�ܝ�FH~����6��%eQ�F����AL�[-��g�*,�S���"O[HXBW0�"���x:�)�֯��͕��EL�q��[���U�W1��gqzv�$���lf.�y�ߑp�����NpS�4�h� ?6=���{<��>l�w�0��F2#�4�&���,�^�7g���>b� �v��S��M���|%Î�NW'}�d��-0H�����X�� l���i����/���MJ��ŘDuY��b�܊�O��C�xl۹Ɲ��1#ʹ���FH�����'��r}�΋�_�Rѧ��C�: 
�jU���	Z�"��c���^��K����T7�f�4�}�ˎ��HsӁ)4�7���&���6�A�+y��{B~H4��_i~���XŪ�D��B}>LP�<t}��<h�OE�N��*��2�H�B�B�g"n:�^P%�J�*e^9�S?J�} ����ޡ`��E��@��t6�RKy]^E���,�q��	E��(�"������c���F�t�(���v�B���QY6�����]���d����������0p@��%��ס�[�� /��r�1�����@����ڭOC�@^^(E����̨�Ib&EG�ݟ�cQ��K��4i[8b-�ϼ�M���^�p˥�dB|��4�e�Y<�/ހ�����4�M�)�$
��)9@��4*��CeE�ƾL%m"ը%}lHx���$-���F��%��B�8��|%ߺ0Q��
~���1�'�E�Y�\p�mΟ����ߔ���`��7ʴ�B�:P��fCc��Y�J��p����G��;��J�0F��в�+(�z5�آ6����Nr�����Y��{N�E��ө� )�4�6�bmp�ͪls^��)"�V��ю��jZbH��
_Oc:$��$�����c��/��\���D��jx�BZ��I?��eU��M����cARt�����A��}��A7��� lOA��q��:��ã�2.��Ӳ!O�:��i�Ş�����D<��8�f����I�{�QR��Ӣ��/��Y�L׆m��#YE���"B���U�H���+�h耂s>�@�IL�$y��@`��������Z�������;�_����!�e�
���W�J��1E��J�HZ��h���>.��}ź|E��92���w:���Nw�x����\���i2�7Em�ï�X��J����v�I��Ȥ���$T<�M*S>�}�SSiy9�L��>�]WHjQL�l�J_WxkI<f_�%���}HZ�Y�٥Y+����'�ʠ��z�7��C�}g�n�94�U w��셥igs��:.�2�k*s������P�b �&���47w��A:Tԇ��䛻r
�8a�o*o�:~��B#��<�1���}��b�U�@E	S�+�@�O��3�.�d����#^�H%��ni��0#E��	V�R��}[�wF��"�ib�wV��_=\^�w^X�>�?u^@A$d���##�=�-JȎ�k�e��p�bo�MH,����%�	����ɲ��L������;�.��D�J���]��t� 6P(k�P��Ơr�hS�%K�����s�?�"��.�_�X�c�Rac͝8� W)����(��l���(�%fދG,ֹY_nodLuDf�Yw��E��[v���R�9Kw�ڻ�#r�f�� ގe���"w�fm���HY�!�z��܎Z��Cc��
��K�\@K�|�O)�w%;�@�̒�z+W�TN*]�E�/���O��t��a�H�k{����������K#�t�d�`�q�p6�1ٙ��.Ea�VX�d�lh�8$|�|L�_v�iBÝ�6�����\m� b�G��&w�)_���(B<a�ͭ�3'~��[��G�G��D���8g-�,/]�^B��X�~�v�x����(�e�Kx_�Ȏy6,5*�:���!���s?}=c��1�YY�U=�+�vVn>u2�K�l�L�h�}l0R��y?��՟rA.��TU�s5
g���lrz�H�Œdx��"��ȧ��ɓ[�:c=s�Zb�ډBp�sQ!�S⿃ �1���*��9j���#Om�`-�������@]�^"f�'��,�w�ph��ܝӯJ:	��~1�5x���`%HD�?c�������f+X~G�_�^��aib:�B�$��q2\�S��u�C����}�q���%�a���u(R�r�¼T����9�X�W���1��ܐꓱ􋴼;J�$��ю/z������ۑ�Q�4��޷�8ŉ�*��T�v��8Xv=IS�I�G["�����2I|Q�T�`��D*hg�u9�+98Dd� �s���S��`�eK��o�(��q0�q%����\��e梛�&��:č��WE>���v�09��:Fڻ4diÖ�q*	�/��?����\܇�<v�vR�#&���1f��*��b64ZG/9Jv�o��]cE�Z�AJ��k�P�Vߺ������W�@ycI9��H��Ǔ���V`$2՜
�*j��a���	�&��f�vu��Nt�J���m�"�6���H+}�r��Q�{��>2�@m���U/�8w�:� �5��	�^�[�22��\����^৅|LDΆ	k���;Q����\&�����Ԋ�&�}Y���f�z.�x�ix󱨂,2�A�SC�8YD�/�t����K��e(�ؾƁZ��_(>���˨cp�U�?"�!����>! �M2����MH)Hm�����;o7H�&��_�Ɣ��d�\�/�����sw��_��S?&W�0���rXC��Cv��q	4�Q��]<��iR��vm~��|v�X�!�@C_D6I����`���"i����vR"L�B�}��v��kP�fDgga���nϏA�VȟT���Xn����a�����[�R	%��T��M�#@b:3څ�(ۭsW�1���'�mc�;��]��������h ��:������:�+����~V�i�v&E�@�`e��^&r	4Sp�ɵ����qR���,��~]��P�c�[�Ŝb��~��(?n�ד�0�I��4�� �ܗB�P.Z9j�mmG���|�������5g��l@��:}0>��y\�y�vs�E K�x.6p��w3m1N#�����!#.]c�D����g~�4�Dٓ=ȡ��9:���l��]��qQ���bQ�"+��)!WܱiWG����Ŋ�0������_�'&��L�H~r���6X���}YM�Dvq���r��tN�OB�YIL���f�������m8;G�N��B���)�je\!*�9���璘���H��"������ϱ �՘WD)/XO���i�_e1�3 �W�ʃ_,9*㒲�k�l��F�>O+�N0Bz����G��ߪ�4x�(x���
��i�Z��|H�*�[�iM6>S����S�s��*N��C��x�Ή����&�<!J�O~�u�'.jg9�4w�-�vRZ����)��,��c20�t����k����ꗷt�)���3�Nd���'+��~Vx�M{,VN��Ȧ���9r_)4zd�$z�Д���JP���H3'ds�mςr�����s��Y3�邫&�3x�!��&'3ȝ@͵��5R�G�g4��Ya����y��������}8ywypk*�(��G�&�L�Og�'T��v�W��%|��q^WEϟ���뤉9 ��~�����|��g��6q
��<�.�4���a�Tzp��Vt��z'uɴ�ֲ����d5�d1���&����2)����v���p���A�o��_?bՠS�h�\xhb!x%n��Ku�4B��8�H^�z��-�j5�dgmdαO�־Q���Хuz�웺
J�zn��_UX���*����� ,O}b�lu�_�5��E�hO���zED\����Vl�5==�0r�Kݵ ���e�fVP#���0�Nԃ6M���]�K��B����p�Ԃ	h�-���՗���4e���"K@ak�B�xgR�&�w�+�N<�P��J�	��:[�?t��ύl���P!�h��''(6�F����� ���E>M6^�.,J)v��G Y��J��ñ/.ry�R��1
���Ev�#��'�'�)2�gj:A2O�|.�z�C�W6ن��D�U^���Ϻ���.�Z+_�Қ�H[�"8|49YB6Y���*�xaE�����6���Ba���ۯ9-+��F���3���r/��G)�{W�u'Ə�������U�RlO��������Ŕ�-�����΀f8x�dh7k�|�����PBS�����_��2S�-��9��?MW�	�I{�$���
x"|$��Vø��	F�`��M��q�:�|<9gz�64?B;Y�L�@�bx;�I)��97����ϙ4.	�DX%4�#��l}
�r����~��(no��(��ínS���G��X�}�t�l��^��: ~�:9���!�8�D�D�����@�0f�,o�(���>P��~��\�Z{YJ��?�1E�b�^��~�ߦ�����e�y����L��E|p&�}�.]���LʲYv�ic�����%���(A��FW�2��',_� 1�7_�_د��j[���� ^D��|��� 7�������+PK�s�u�z	��\�^�� ���.��9�1d�}N�e�ǯ�@�=�::I&�Ų��.��}������F՘a�o55mr�暯a^y��BVC|dOb��Y��`V3���2ԨMZ�!���l�3�_P��Y!��>]�ױ��:dMǵ.E��E*>@Z�*��_���/���6"�\�a��wN�n|��ҷ��X-���'�$�vD�T�aM5O�4a���l�yiT����"��o���}brip��Oxk��Ѫ�$و����"KG�ƙz�y��@�Bz��.�.�R\��7s�(UڭfJ����K�Hv(�5�A:V��"��Z}�_i���)n���������Ëv*r���*b&순'�pc�ɸ��e�<���t���|�uv��Ĕṩ¾�[?e�k�߃;�b�W�����K���1�%�}�a��-8����&��/jhK0+ӍNo�P��+\Z-Q�|t;?N1q7�rfй����hE����ƛG)�露�iX��D����O"�<��l��S�泓�n�	��/b9t;2i0��(f��U��RY��D���7&�$��$�(������pZF̒f�6,���X�n�;U�(��ڂyX�Q���C����^��v����o9��Cſ߭���$�x`�����l5�x-Q����WM?K��m#�u��L~^�sդ^Mw8���|����l��:I�,��Ѧos?E�՞Y^�2\�E��{u�����HX���ߘ���SbSIJ⒦i����uu.��]0뒭Xѯ�h\Z/:t�J�D��*o��eP���{�AJWߒCY�Tw����5�{������+�6c��7�ĸjR�g�����A�������k�އZU�uP��pB�����Ǚ�6X^lͩ=���@;��d�N7_��W}���G�Y�m������D8?MDT{�-Aoc��<�R�����M-�Fv�%)$w8�"v l�8b����:�>;p��6�E�a)�=u�I�6��B� !"M�;`�^��V.=�PC�R�<6*�B�� ~��@MP����d?��U�X	H�t��l~Ў׿`��?�p��J���ʌ�+wG������i�(&�t�j�T���i���!?&ZsXu�ms� 16�=���vPw��}���Y(���k5?/�E)��@К$��=M�$�:�Z��ۺ���l�X��C�@re%�8d���w'#7���K�J�4E�"�M7��Ɲ*����w~�wT;�|g`�S�Aɶhv$4��v��R��,��#�ϑ��B9~@������t�}��V��K|?O��_���l�R��g�%ԴJ�v-��B &T�V��!��^���T�����fWmJ@������:���n��Uz�
t�[�).e�����(��&L�<�8���s漢#����H��e,7��)E7z��t��{
e���n5�1oSa��Oҵn%J���]Q�E��',�[�vG1�Rn�B�0��? ?m�<`T'/��ѹ�����Q/�G	?�rg����~;m�bd�d"��,aQ�>�َx�6t�`��l�	�$��TƇ�خ�2^a�N�
#�%�l��*��q�P��yPN�@�!`^ת�6���C}h��-��fΥ&bO�Mq$g�cNIq -_�oV��'�Cǝ��	��^��!\���7l"�k�sgpZ����{��a�����x1Յ�ҋ��x��r+?�p2��R�,g�g_k��҅LX����k���ou��ҟ����PGn�ަ.�#�c}Öb�+X�;�Zmyh���T"C��Sw��BE�{���;-�r�n���QI�Fv�-V�7 ��s�MC�s���y�l���e��'h��1���|#��am,��f/>���ܸZ�R���ȁ��藍��l� �����=q��@���P�z��Bp�i�:�E���f�#a'Mb�]�v��sU:mVb�A���
:ޫ�݁�u�`����A\��i�3VL���B�sg�'�"�8�W
2���m����닗��e������B}3J�w�n!��	�=T�/�DY��{�ʷD4N�j$`X����gۄO	�����.X����~�#�^� Tt������#��]�shS���x�_L:R��wzk_�	�m�Bp�bx��������yG�4�g�;":!�������vT%LF�L;r�5_yAt��\aqz�a?����_Vsy����$ch���d(�h��@��n��u�)��[DDZv��Zpٻ��4��E���2�.��X=���mg袰F�G.<x�	��U[w}q8T����K!C,7�3�]������eO�}�l�w�"�ih�$���� 4��	�6@��2�� ��<��h]Q����5W���06J-�$�U��z.,���4<v����IL5 >��ʳ�R�R8��ѳV���O�VxB?��꼔Omz�Bj�,Sߌj���)[az1�X��{��L{���Tr�G�ԪI���u�3��չ�͇9o95�9N�Q����t���4�X���ΉGy�W~h�!B�g����ޜo*l��r�䁂�3�A�`�B*�1��ź�C�!m�?��1>,nW���0F� ��fsy����A~�Cd+�p��D�S������[ɥV�M��w*< �7;�M��1�O�X ^�������a:�X�}�xP� �ojfv���l�iRƿ��?��D�+U��7�衹C�e&ʝ��a5hq�WX��x���.��C���7�B�Yu?��� ����i������;�YP����A���t�� ����D"�W�ą����P��t�?�E�Bl��OP����?�%��x#�TY�%"S��b?�(� �X��,�L�^�^$,�
`��(�z�v&���/&�U��u��e`t#�A<g܅I���1	߿]n�95�����������JbQ�˅Cv?ۺ���ԏ������Z��Y4Ĩ�#
�o����n��c&���� �9GGT���C+�`mVB�Mu�v�9E�y��;�
��4�����-)���H��r���W�,-�ԩ:F�[�l��� QZ%E���Wz�E,XV��m�A���/4�b�a0�?�"�C:�U� Anԥ��aU-��GW�+1�7ی��T����7a�.��enIw�b��͹�*�_��q�F1���h�ɢ/,_�|��(	K6ȭ'��@�?$�=Y��4P�wf��D\��4���d!��pu��~�K\�^�/$�+X����fq�ɨ5�u?�d���6�2n�:���3���+�MA �4~ѩu���*5P��rP�L��y��Sy��g��{i��fb�����zB��U��f�M���$�9}x�j�ZM�Ŏ�,ux��#|��R�!IUs����bB�{4���[����ou�Gy��ƌ����;�5C��c{��|���ծ�<���QS���
i"��Ĩ�^w��WV�\\s\� Wa�^�l'I���u�j<վs(Li�
ݜ�o��J>vYP��|ݧ��n3I9w[j��5C��:Rj�[�xk��t�[�c�V���4{:�������a�W��Tp5� ������G�0qt�^��n�&����$_Ъ8FԹT/(�9��^�A(����d���M�ԢZ�A��}�y���ێU������v�����tt?��<9�k8�(�������qcEM����M����lwW��@!<���+{��yˋ�]Lx*��N�L�q�ʉ��D)�v���D��#��=7�}�wx@�ASu���/�� �e���F�&�z�S�"л+�>����O���o�01 g��O�_�6��������r��Qx��å�6fZu���D0����d�-����FhIhl{�h2���`�;)r��ߣ�a�a^�`���K[�����oqw���n���|B��ތ���ɢyZ���
�W"�\_����M(0�{Y��~��:v���z��R��|Ԉ�Sg�=Ջ���:M�"KMO�v�~�@���UF�.��djD�>��#Z�g�l	xr�j�^������<�b���jY0_&��$�{8�i������S��2��L�j���'G�5�!P����%@M~Ɠ~���o�$�F�s%p9j/Ģ.�0"�Bad/F�Kk���(^�C����m���E�#o|2i%�OT�P3#��"U!����݋M(�1�"B�k	��mo����FV"�j�[s@��?gp��J���
 j°F/G�drA�l�(%Rwt�K��dy�m��{f^������tHD�
.�&���`���H-�Ϸ�A;�gY6[#ܖ���1�h��k��5�܈�"��:�����{M_��:�?уZhs��S\��6�7� �ö��P���-���@֘��w2g�J2����Y�n���Y�jw*@@�����@�A�X<��)w����`���g>����Qڡb������9�(�t��2sJ�H���#t�}T蚛��[I/�(�9SL���J_��S
�&�W�i(��tZ"�����	{�k�'��U��LH��ۍl�J�9�p�I��o�N[��p�B��F�w�!	�q��AŅ0���C�*��Y���A�jmE���3���k��O�  �pHWޣ�M�S�F�Y��R̉,���'�2|Z! \oM� a�W�~�O
pqf�F��A� ��!��6SW��s�+-�FƊf�$�����ijwro��Zx�w ��S��W����?�P�~�3tLr�Q䯨�i�t�蚑�$�sPBpK�M3�H��"+�q58��>��M"b�_��Ʃ��d*���;�IJ���֌,�~?*�_¹��.�&��NDи�f�+��<�Z��������R�M������Ƽۃ! ��(5�$<�Db� ����D�B���ED�7�!�m��U۰��kwv�BF�����o8k�-dS8.�8��=8E��YfW$H|>���Wa����¯�N�r4t�O���Α��	�^P�cm��1*���*�,�u^=�������-�'Y�fR���\!�`ɲ�+�)�_2�d�.$@pBL��p�)���T�O1��`�49��<#D��)!��V�)�ԅ�ӈm��W{ܓ��W̴�/���T㒿�c��~u�DVx� =�y�ܯ��J��k�3˗�Y����P`��2���V�Ǡ>@-�Ƌ��	�^��3޵�.=��w��}�K��­udS��DDm�Nz�}g�1f~�����.}8�X�-����U���6C���FJSg?�����1�z͏�+��R�����y{/��d�|�P���_^\? *�륞��DE�#C;�Y��
�	(xp4K���IBA���%����G@G�'�֘�C�2���Ҧ��o2��HARG�����_�˦�7�A;�ӌ��R�v�q@�'_�%� ��G��Z�n�
�����>pSԘWp���G⤾J�C��f/�T;�o@�&E-�b͔O�d�����||*����W�q�H��0��ªGv���_I�����W�0���
UE>Y~P���Wɺ��2��l��=N+�a�#epI?��O),&�G��L��`a��Ln�Α}	;�$ő<H�Ɍ����E �ZwC�ts�r��gG�ni�����P>���.߃��L�AD�s�o9c
B��t�����G�;K���l�����x�H�Tu��KZ�h&%A�f�k9U-�T����+��q��Z ���j(�i������a�������ו�[���}<�qɗ�<�YG�pE��~�Q����w�U��\�X>Z�j����Z�yɏ��1W�D�6�c�]mx�@����"r ��������E}��u�`�1���ǁ��&�,���Fs;)��C4�$��LF��z>2���]aF�l��%��Rո���K�:��5�*֜���C~ey����B�͊9�Ik��P�1��_���T�&�uယ�=D]W�-$��1��%|�����lq�h!C�!���#��꡸<ّB�?��ߢ(WahN�נK�7�K�"X��E0�#Ph�f'u!��Y��T4Tt��ܬ�&�B�J�$r���X�B���KC���+��\[����"H�5b��vv�jV �$��vc��s�2���
`�d���8p
�I�1�<�֔9���v}P�w1˦���ej'��"�rv1��'#�Z�9��dمn	�Wvr��ПtK��uӯ�0�8�u��J�l�Nh�b�{��A�B|�^�ɤ��ؙ)vk4*lZ}/P[;�BCo7��WB�ٝ�=��}�ֹhU�Q��4͡	�p:�G�)F��~��ۇp�5����X�%'ߧ��O��cgG�0vV��[��x��=�o7`�Vd
*Vּ�t�N�e#Ѓ��ګ|F�Z[�??)���T�W�
��\��>���^W��M[7E8�ж��'JE�����vr��`iL�m�[��h����*e
��0v�@�H�2�M�G�0e�8+��yĳ8պ'�v@ؗ�ZX��Z�`�2�9�k���nr��;�0�'m�睑����4��#r0�c'�g��<0��pS-r��m
�(�Ke	�9H�6E�&ͳ �Y���f��2v&@��}��u�"�>��n�n���3��jo֎���~-z�@��ڠxXY�̋��3���*�;H����J*��ݫ{��ɥ&��2^9;�plb֧*���� �j�Fx8�/���Tu"��Q�dt�SK��ק�Ik���y�� ��$�HBv�I�p5G=�LG��JKU��=�/C���5��`�ap��`��aV���D�s	&7��`�WbF�Y���H0̉	�;�G��J,��^�M��sCb�@�[昼n5��^��s<iKa��S(�'A5��` c�{�Z�g��kH����`��?G���'F�HM6�����wY�U|�NC�D�z�8u�yAI"��
�5�T9.����p�]T�j��ɽ��pJK��4�r�rV�@&�0�;�<�`��a"�|����`?�)�E��FTaQK�܅9�_(J�Wq�H�ٚ-��aV�*.������������j"1BL�ϟJG������6�r�]�`���� U�oѸR�p u�����D��%1���)�p��Pv�^��4��C���4}�x:�&U5PB1!��R#9Y����nQĚ��9f���X�A�1r�U��dZ��(�&�8�0���c���n����G=��i4���OU��:E#*F3��6s� o�8��>v����x��y$�L/re0҆�ע���t:�9�w�}�ݍ"����_��io�X���Z��~$�Y��O�Y����3�;��I�2�c9��v'�vv�0��!���r�A���/S~���:�؟ڛ���V��a�
�(z�v���x�4���l)�S��gA�Ώ7�jւ1yR��P��{�`}eB�ʉv�qK���Hl�z;p]�>[�z8]�������,j�/�K��}�����Kb3��
����a�W6�|�螂�H�W�E�d�R��>ː��w�д"��%E[��R\B�n���g�R���Zg����j(浝�lF��)�����Y@���ǂ��5@�b����W ��"h�m���('6��E)T�t���%iK��w'㬣��Jj)ߓ�W�>n9P��r~���rl��]�2�r*��Cɻ�G��-8Y]qմ�-]����� xN ၺ4�o��s�{���3�ĕ��#����̍����$V0�"%�L�X�|M�/�4Uv�d2�do����U3C��A�.F"�@���eO}�.(JV���4j4d��f0ǆ���e�N`�>��H�lFġomly�H×u���r��K%�uf��f�����{3gB�8�r�N9����xzI]�V�NC��w�V��g��_$��;���9�g���A+k���\{�D*<��oU�W�Ó4i��8�nB�V�W��Ƀ?��Z�2���@���Q .�����ɩxc F��j=0�+h2:���;5��L-D��w���r�c��~�;�ਞ��ЎO]���B�̓�Ekx:0�z�'._ Q! ��Rٳ[.و�T�T��=�d���������\���P��bT5�i�To�����X����q��E�:&�\<���-�}"��@o�h�
���EWZ˰�Dt����-R�3���	�+kA���ٸ2t��7/Ԑ��9�/�ӎ��Pdde0,62{� ���d�n7~K���oi��C���φn�k����QRƬfC
�n�`
�A�l�Qs|d�b�;�B^��؀��1'�w�3�oI�")6yJe7۴;x��9�5<; K��?8�:��p�oK�[
���ɮb8U	ܺ����$�%�d�3����yq���A�TZ�$�<�M�?���r�E��A���SZ.�De�.���[��%�O��jk��T��u\ek����bf�����s���#Pp��oLԕ��|"��"|�Y��L�Z��|��jG�'4�Yq�6
(�<�)&*s�~dL@�4I�+DD<s�7�^f��Ji���U ��j����+��.���K3~�_��~X��qLĭ�/�IԦ����{<�d�����f~)���Pcz��"%��_�C��z�5���:�a
)��W�D��F��PB�Ѥ�.p�
t�ck�� Ϸ��j�e�Wf�>�0a��Ӧ3�.�"/��w>��r�Z["�����eyȻ�a��
<����bs	�C��牼�J�	x�16��/������!�==
����v�8�9V�A���L��5��ρ�O ������QD�����x�v	��݋���}��d��uTh¯�I��Fz�z�0 �!�`�C�!y<-��l&�V"0������������%cn�.Gn�:�^�����a]��
@�JK�!z}�a�S^=�W���ں�����:�4v���+J��+蘉p!c�����59�����FS�Կ�9��r���F��g:���/�|ؠ}��-�W�Pm�v���e�A�f엉:(]�Pd��C&��cztv=�"�V�Q2�x���?�7\��R;�~��w�lPQ���Zn�֛��!�D�#!rn`2�U��,�ܳ��O�tY��&�9~7Y���z�\+�\�Y,XDqb����˫T�t=��P�(O��
n��w�&�$���A	]߫�O�\��:�c����YX���'�����,~RQ��Q�`2N��7�x����bC���\������Bӎ��*K�T��I�K;;���|�� �$A����z���^y���b)��	�#B��o��YtDz F��J��K���: &[x^�� �/��S9C	UD��M07�*iY������;y9$e�'I?!�C�.\��ӥP�f���a>R�̡�/�"n �{S�V��^x��YB�'����	A�J���b�m��`�Q��8�!-�yF��I{�5����&b��<������-�@������(b�h,B� n�2T��Sz�>�N����*�`��f ���f�+j���nģ��llLto_�O���S�n��n�����B{�3�b��/UBJ�5�k1��&��	���3X��=��j]�)�J��
�rh)f�<+��0���7��`����$vw�����=%���.��|!pGŝRӓ�"�ڹ��t)v��y���Zܚ�0 z�9�#��1�Q=�H�uE��F)OV�\�ӷ[nM����6����Ö��G"�	� ��B�&
�T6������A�@�+�����6 ���+�y�O��L�8@��M�`?�i�i��~5<@E��{|]W���u��|H�l֣蕈��M��P�i�$j�G�W$b��g����p�����!�����1 �e,իT!%��6��)	�ֻ|+����tA|���Qq������R.
�L�$Q���S�fo8H
G��8"(;��b���@ޱR���*��CNH2=�	�cc`Vn��N@�>��+h3 ?�'E���b����5�a�	4�9q\���{DO�VӘ���	����s�3z�Q�Z�F�B���S����{
d���R�^��eS��a��
/��P	��KI�ܥ�V�61
���Iɟs�gЯ�SQK��#tr͉�Q�-,��4��w�O�=�Ͻ��Ԁwu��燊�Ԏ���$�gjYkZ���A���)w�Y�H�u��:�(����(Ι����6F;KT���#Veo�,(d��G&YPï����:5�E�m�KT�7���~��xb�`Mߏ6�vt�tibE��OC�ڬ�JսQ���u�"cf�=�K1�B�%h�m]�Oksƥq�t~Q��ւ�9aU�[ډ�#��`����#��ش��;��Cv���RC=�6e��1�d  �f`� �
��ҍ�������%�r�����5p�#7$��p��*�~�ϑ#|��K2&Lj/(F�^����9�jĽ�Z�
�Im����;��%;��P%^N����z
�K�]kg���n��q*�He~L�'nU�����7�o�1
���)L���H��$�e�ܣ �:����J���m����/��]:=�qU���G��C��	s<Y��f�zi�%G�v:ڒ����X����M4����(���ֿⲾ�Xi%�ݼ�b�p35�^�[Ӏm�ٿ^7u>�S~�H��s���)�I]�o&�$�)��c��%�.���G�2���F������P�!�bq�#R!5�:��!n�Գ��׻�,�r� �t��X�z������{L������îO(��r-�/��ܞ���%��b���p��
�w{\��jx�R�srM�&�ǉ�� �a:�����$I�b3���I���8{�Q�1���eq7?���C��������Z�D[L�����U�V��Տ��9	�]��p-�ϕ](�(�F=�GZB�GY)zFZ/]�K�B���z;�;���ȡ~���2_e��{����>Ez��+�Y���X�S��i� ����.�� 6n�{�I�����@G�]���0t�U2�Mz!�s����,���7�R�pl~�ā�!�����0�
�0퇞���4�A�������-�ݵ�$F ��+�)1�%�2̞l�)$i����ď��lP�pÿ�t		l?�c��{�`�-VI�4���%OP��3jю��v{�0L�������?d��P�\����;O,1F�>����z�����Q���W$�J�����n�>���^f�ޘ�S�����FDQ��˂���|ݕ��;8��#��)�t�
uQf�l��<a�t�7�n��\�B��Qň7�^OsqF�6H�@l �bS�)gK-���c�u~?=]��U�ā7�THK^�E��!�A�XA�* %w�x���ؚ'�?Ī%3k��k��m� �D��鸳���KJ��7h��i%��I���]+��4��I˻]�N{&Z�a�2�xH��Á��9�[�Xk���u�ph|����0�Ĕ��/s0��_�(R�TLe��G�"qy����z/�7���y>��:'ܯ/�	�a�Eһ�~�����߂m9��ج�����i����?����t��<���Gm&ظ\GlL[Op��~	_��� ���pv��t�-��dɘ'9,�jt٣4n�+7�����e�T�`��Y��ǻZ�|���b^��a��{�u�{-�;U�A�&�+l��t"_υr�V�-!�	�Z�8/���Xł֞�>c������c�8?0*�ƫ���&������Q�]�g<B0��j�����{〪����ۚr��U����U��w����m.���9�^U���+�P^���������IU��3G6�D�`��$�3�T��v�C����}!e�Ƽ貄��M��"V!������;b���2L��b˯����Q�b�T��u�*l�rS�r�՚��+�����bW��9�s:p��K��fQ�C�Mg�����A� �
�
g����J:��r�DFҰN��Q2�iݍq�L���ؐo�]�PU�qKĔj���NS����.����Ԓ6�޴�n��W�^�Pm��l�����4�J�\���s��9����3�p��TvS���.@*����pb���Hp�綶�U��B��%�E��w⊨��y��_`@�0c�����C���8�ܽ�F�i��;��P����
��{��֪�֨�Cx9)  �}��p��T	�Mv�wr��=���{^�biU�S��&ZtH��Ot�v\х� ]���]�pX5�� �����0n ��s�M��-ƕ[�XVl��Ԣ�0��r�-�Ef����k�+�.��bm2��7��O��,���ot�_̜%:d�l3(� D�SyP�u����s�{0��� %B�Sa��Wrj�5�du�x���y a!�^����`;Ov���;����F�:�O���]�;�D5��}������G�T!ϼ��y�q�;����G�j�#��E������ΥKH��͑D��4�z�*�#VY�L��L�3h���jW^|c$`��X���a��y��:�2Z�����~)�1��"-�����G2�,�㾞2h��X}I�i�>Ay�gJ�>�)9�m!i�پ�hʌ2l��[5	�O�$E:�!��6����+.պ�R��>;����C˝���ލ�|�K�Ms��!_#'ߒ���ß�M�ۢ�M��ԗ/z�o~B�
����L&�?��w�)/�.^`<E�Oo��Wi�E?��i����-,.3Slt���v�	�փx8#�H��>p�Y���~�?'���5�:��B�[�tX%רW|�	L���ދ���������iYM�KJ��W�]��0[`F���3��K��*�|cϮ�~��f�J���^]�w����5�{3G�:s7f��ˡ�QɃ���Qϰ1��2^�*�칙i`��������A	4ǣ��"~iRй�^��+as���T�}=+4����	�h�9 sO�eolr�0���-�(e�9!%�e�O���D~����%P��#�S�o�c�H���R���Mxk���d��L����@�=,�q�m ������Z���|�3��cpćԬ��s��}I��h��Tꂭ6�<�i���t(�PBKT1#[=� f~�K�ar�`�c��7��$]a��� �����5̀��	:]٢�)	�p��-z8'��z���l~�s�N�I/��r�0O���Ҋ<���a�9���%Z�l��m��q���VEH�����s�hKdG:�!wt�!Q��x|0�_A�w:��`���:*�� ���E�V���6d��8��Ͱ�1�L��{.�C����=�c >��������r�q���g�]9X� A8�ݪh#�U�}�5�ʤ���8:�)�5&k݇@>+����8��#3�O�W�3�rEvss0�7ل�`b� �X�p˱�0�z� ]���쓖$���(s?�f�j c XlCRW��C���;�R�B��G�R]��5
���?{{��:�E`�z��t�%��&�FB�~�a��ԃ�k�<�ƭ�~i�/8�U����1�����R�=��;���pE��?z�@�����|1r�n]K?�@6��=����\dǎ/7Ũc x���]R�R�[ܧ�z5C��ʲ���b�"��Se+}C�����َIG��n��5^�܆❑z�>� �[�y�f	�b����n������P�rK������O�L��� ��;Q�C��N9F�Xi��$��L�G�sŅ�U�� �r'Ɛ3�F��i�W�ئ3���X�k
n���o�����2���>b���)/qw:��<�#�\�m��`A�]3��K.o#��x\�-t&:���+C���tO|�,Q����KE�1�^8����Z>]ӝ����` ���A~���9��W>0���ø�սa�N/�&���õ��_�
1���-M/��~�s�(3s�aV��R��A��9rD�Mo���7�3J覮�6� z�w�+�������<zR�Byܑ����5�T���}-�&��(]��{V}�8��G�Z���c���L��Y�(\��V����뜫f�H�*�u�#" ���G�f��+��u�}����^�����$��5^�R�i#$��x 3��
6[��Oe������@���!&�]����Ra�;�J����76�6W"ҍ���X��}�E�\s�'vd<g��@0���}}�r{L"2z6&�i;�
�$G'�R��l� 6i�N�CV�����;�!
-�_��v4ȴ�E����U�Q�a��Jhg� ��QF��F=ۃ��=ܑ��J���V�*�K�!ͽfr��� 2���� �!Ǿ�H:2]D���n���l��%L�c�\�@Q��<�H�'�A�ơH7��&�)Q'�`�g]3i��vn���5��Xyھn
��h�g�K�ׯ�B <�e~����ġ�!����/�I�#���ëX����>�ޒ
��M��5-�C����i��u�H�� {p�kX儉&�|��P�
�(K��Ub_z�5ԚDoK�����LH�a1%Բj�w�C6�������S�����i��{�:s�Gj"9��/�rY��[L�E���<ҢY�#@:�+��N��F�Z�nO�\�VL���¡7�tw��Pc�s.ǐ9�N�|I�욺�E-��֛�}�?�YBIY>�/̟���W5��Ñ�Y�t��&o(
��"I�hR&�Qv,.��`�U�� �Cc�ֶk��*Ba�*�$��o��3�j�)�~�|�O�vX�aξ�!rYbj�]2n�y���G-���훨�.�g-�ɮ���|I�*Ve��>�9���ɬK���c��p�ĺ���k�j]����&*G���6�R�x��[�a�E�w��Ö��7���?J��i���ݡr��UE�K>#勨���QTz��Bi��K\3{T�i0oAb�8�^�Xt�,��ޙ��[m��21���Y���$�oJO-X�	*fǘ���>�=����\��V�kK��i��[��\i�t��!�	���`E1� w*-�	�Z���1�\�Rp�#\DQ}W��%���(��ƒ���ު��kx�����,{� k�Q���lJ�#q?JK�G��?6'�[~������MA�R}�� lW}ǝ������<���5Ϟ6.��	H1�%0Ȱ�Q^�D��#F��F�����"�q�~�|�R�D:�/~n���(��s�-�c��Ί�h}�+Xh{·ҵDU��G���~(����m���m��A���܊^W'�����\,�%F�x^;���,�5	��+H��!����a˺���k�eR�п�EGC�cA�/�ZV��HW�u��l+k����zjg�M��Aq��G�E�c��f�@U����d\��}�������y|�Lb�
dy�P��s�^����P������$㶼C�y�+��!�r�_�N5��(�"91f56.6���t�f��N�܃��ŭ{f���قC�����)J FTe%P�^4�ȻVƩqGN����s�����A]	�o,s
�B����MW�.*�f�@8}�lvS,�$��&;^p��q�� �t�o,��:���p����z��}]�D:�g�ʢT%�M=;5��v\����+kM���{�?������R����ݙv Pw���p>��w$5f�g���5|��]�0�u8&:v9o9���_ !�݃��R<q�eFEp����Ui��W%:�<��4u�*O1[Fo�)9_��l=1g�[��+��<�t)��I׭"�����q�{A�M}��B]��ᵉ��������X�2Γ���VȾ��r�W�8T����Jԧ҃v�����z���~n��3�2cz ���<��=�:�I�YW/z���W���I��D72������n`q&�<��P��5Q�6�)����z�lh2��>�v���om�a�d���d�4}���	S�.3ߩe]]~��R z	roZW��E���5���0/m�%L!�=����y}Xi�ga��ΒѢg]�q��җ�/'9)+Q�P]%���!�S�U��L��\(\͎�v�4?̄�.��:�ؐ�xɎV82��8Fp���2?�Jf�C۹YB#��.o]��*8f.v+��pYI�w��T>~�U�rZ[�{�,pxy-$��3F��>c;�o��_�-A�zKu����I�]��Cn��/&j�"�}�uKy#��_��.d��u����4���(ˉ+���\��S_V�>g�V���P`b5Y��W甩{�ܴR?2n��b"�A~K�:]X��p�r��8qY����8����K��.�.I^mV/X<�5�C�a�9Ր�L��J��S
[�´O�F_���\ʚ]�z���Q$���(�Q��Gf�h��RZ�q�w�-@�l����T��n�dp�d��r�ERԳ��{�S�L*,f"�R� �0y+��T/�)�6�=~�k'}���Rp��P��<��j�V�J�_�V@�|i���L�y�ؔ��(	[k�����z���8���[��I�A��I� ���"+�O�z23uf����e�	BB�����I6-�eo^idv����c�Y��e�	R����p6��6�Ɛ24�S�,"*4���*0'.�6�������5#W�F���+V"rT<��
�S `���{�_%9�_k����ݚ��P=�%z�JK��aI�6��u���Ё��t������(3�.��,:	F�N������<ˑ��b�O���UjV��Ctf�e'T9��4� H���տJ�e^�L8�7&��>�*��%%��sC7�
������yB������������"�O���GN_��Èy8R$�~ȃy��Z���N'|yY�v�,�ӈv{���+Xl����q��Tz�7�;E1ǫ?I�A��F/��mn�+o���'S��g�둅��w�_�-@|��T�cH� ������cɔ�����t���sӨ|��w�h$ ������`�d�S��~�\�E���pb�U��#lK���	�g	�t�0�E`�i��+���|�"������,��$+��z��$}&��%%ղ��?,��蕍��~A��pu�y��ڟ�q���'�9����5������a�!B���oz.��Ԉ�ə��%��J�8���4��b�#����J�.��(�x�[d����^\�I��#{S�ZI�ǙG-/�i��OkdNe��:xIl�*�3���y?\�K/+�/���u!5�\g���v���c�"sQ����Ym��3_��zu����g�����R������,�x5�1��6���o�Q��� _xI�@;�������	,j&Qqf����0^=
y�sőh�b��-�����q��S"}����{������G�q�So��)�k̶���+�L!q��[��Z��N�m��KER(E�;Į ���� �'��ONVe��	 ڿ��t��Q��L��ظ������|����$�A�l���ɻU{�4g8F�9ͅ��/	Ɠ@ ����ƸT�� .�A�vfL�E�X���W~|I���l�Hb���Omk{���'�:<��vL<�䐻�����A��}k�r�q��]�XI�{˾�G����|43��uK��w;%�����=�Ȼ�a��@F���<Q)Pd
z�5��kT52�N"�|L�������ù�{�����(�['�����X
��Xf[������$��Y�m��p��,�#�eU��Q��*�;!�����לH҅��nѐ�uK���ˑ�P�x����ݑ&o��-���5�i]��
3�'���WB.���Jo6qv�5י�J����W6��2��{����Nǣc�+|w ��/e�/�]�d����RV���z<�E�a�͒��I�aʹ��Ƴ�t-63�
�>!wq�	�� �ì���|��V�L_b}�	���,���̠��lJ�ؽ[������;u+J�}�5%D�N刨�<{4p䢐���o�&���亏��鲦�W��G��>U<t�I�ȴ���"m	c_c�<�1)�����B��Bk)^�fK�4�㛏�lf�S��J6���UV: rh��qe]���`8]���\��<���yb� D���ť�="�ʰ�Z�:l-��R�;׬���)�,��E�3����@� �hҭb`��6�տ��Ę�۷����ޮ�P���2N�SCH�jJ���P�b����L�����<Q[j �P�nĳN�n���l4\-��u�#<��� ÿ�[ֻ��U��.�}5V�t�An�>� ���s�IE�KQ�C7�$E�*T���os�T��6fØ��7]m�o��|4N�[u	v �ݩ@�/l�;qgs�m�.�=[7)B��n�猊ib5$[7N�����>�F��p#7�c%3Ҫ^�1��ʔ����x�N 	+0t�-9m��94�|��=�+z�H�:�ˀ5R�R�P-xp&��N��i���m�j�?�"���+��~�������R*�8����Ȃ#C�A=>k/&���f^���8�1�B����e��Ef�h?�Gj�� ;n���w�E��&(�:o��^�#Y�,�yA���<�dv��j'~�-�B�`^��r���g�d��	����ڎ�G�a'>���i�.C����2����Ԥ���c)H�,�g�ه5S���X�ޓٻu�Np��c�! �t���藓�|Ba�(@:]�zX�V�G_�:_����}�RPm����5p*"ބᇬ��%�ފV�(j�����2d��D�]������1DJcJ��Q�d)��1P�����1k�(���V�W��@�5�Y�N��P}��#e�ˇ�� %]��ʒV����$����`Q�GK�n d��^�j}��Pg`ă��ʈh6G'�?c��岽'���y�7��i��e�Oh.��׊^D6�5զ%�Y�'2� �~��8g�,��U���{E�>�f�^�m0d���=%⯯�_�t�/e�E/��?ԓ�22���_$����c����)��i��X�66�vp�G���e?�)c��}-�e�<�fױKa�����-�R����6��ˬ��"B�}e�_�H�BмH���}5��ll<8��b3�ߺ\�3���%��nu�!�	��ѻ��[\b���e��!	ѧS��?q0���[��?T��Y�'������@�O4����-�n�z醖.����&�?��B9ך���5�� ꃩ��T|`�B����q3{�唧;�����0B2.U��A�L��V�|5Bx��K#^h�^�[=]��vQ{��.Ѱ$�$�^"�Q�M�S����oΈ��:ʙ�!�jme�5��		��<

�p�z����!��i�=�B���w��.jv�ŗ'��C��I+/lD��,��9��
��60�6L������O�?%�7"�ٓ>2u3�Rϼ�r�1\a�")�P&��ۆ�Z��2]�����9^��
��9/ng�'�)@C���|�t�j��fb�@V�8t@ K�%0�Nr��2Y,r@�	�k�B
˔U���l�@�L��������tra*%fh��A�����c���NV������7j�O�p9�t���?���ZO4aa?D{WŃF��|�������!�'<ĕp]��_���/j;��˳FQ�W�����K�3*��e'+����A�H����- qo�0|j���廄 �6����sF2����OϦ��B.���2�ߺM��0�7�����-[��:�f�.P�d�J|Í��`�.!6�qt{��Y/�o_�ѣ �_�x̉�đ�D��� �2(��y�g�m�+Gx�WS;�͐�Y�u�22aO_��w�!��ڵ��냐�U��,���7
{��rZt�&�f��p_�yD���Ib��mo�	B�����W�q�c>�VZ��A2\��%8��l�,�N��Iۺu���<�,=/c���x;y7�V�[���(�4a}�b=Oj���V�5��b��%	�#������18�*NR��@��{u�}C����6��"<����_�L^��Uh�T��d��y��::��Ӌ�����k�!~�i���^���	��`l�l��#�@�m��1��J05�i��U���Y�ЖK�/��a ���'��<�����ֿ~�JP���"AQ���Ϳ�C�8�V�+��s/=/����/�](.f�nwi����)�ȅ�ڈT�J悡&O��{�q�l� ��/D���!�v�L�:e[�o���v+q���n��%v�r�C%;ℵ��O�ߓ��
b����I����j�09�_7��<�����I�Æ|ڰ��S�Ct+��SKv����|�؋�5=[_�R?,�pô6��ޫ�R��g�0��ϲ��l�!Eϥ�u�9}�����W_#ւ���>�2��BŬ/��΁td
�k �w�tn��lê�+����^5
����L� g��� l(_��X�������-�ʛ��y�>�Mv$�˫{�vap��1~Њ���QL��8i|��|��Je$�����D��o���w���w�=��l�1o�Ώ@P�v6���#W��le:jfB���~��\�!�m��!��Z&�J���������/71�j�K6,9��~�"`G]�X&�� 3f�R�F���o;Ou�|Of~5��\���*D��̀�I�� �A�J@�>M���3��{���*ߵ�^�y�c�c̙0��g*��7;?X��0�!��`�_�x�e�����u(7�i)j�Wec�e�����8�����IG��rV���EN��#�@Y6y�Y�9W �u���j.`m�=Yw�~���n���W/3)��i���WɃC���#���S�z=c?7�"o�v�������t���NNK��۹A��ް(����;y��ܣ�mǜ�ͺR�KT�=����f��~
��r����-�pD��vw+Q{���O������c.�I�B���e����׺Q�5t�}�� /�:����m���i��ۡ��n���Ŀ���Su��	���$�1�a��Þ��ۊ��X��M�c�:�ݘ�M(�{�W����0S	R7�/w%eL�Y��YcvL����:��XE ��Y��N��+G�ҵ���k�k87�T	�[���U�HK��k.�C�9�(����"�����vQ�V��|��?�x���Jʛ�D���1��y]�wx��@,؇���غn�+���4o�-�J�hs�3�e���q�}���Ӭ����,އƚ�{Ȉ�!? �{b��1�l�NOY��}��t���5�~�E�n}��EϬ}ǝ�?'E����Ҹt��_���
���z�#ϒ�3���֔�b��wRP��0�ػdA�Wn��[�A�O�����V{�?e`t�C���"���;4Փ�����C!�;f�2�7��&�d�}�q���K�1�����j���sh��*-�8����p�Ol'	��e�E[��3�T/Z;�PD��#Q1���u�z��F)�Q;X4�auf[��B�J��^���AMyĽ��N#�T���!�1��������h��V���vP����X.mQ�b|a:sD
�����8�zꅕPW����T�L:��%���3��E��y�&?������t>{��eA6C/��������+x"Q�?|D����DPF3��S�p�2��8h�t�y�3��ܸ�mD������ ��NϠ�X���'�h��F^ۘUs�J6�x$��L�$�YZ�l4cm-�ѝi���p��jjq��#�1c�N����d���&���Z��t|��a���߰�)"��rH���)@�����B����*�G��l�_�-1:�� `M��N�5Q��8�&3/n@�S�0�		���tfB���o� �4-�AQ�(c�k��?��������T-4ɕ��RB�ӗl��W;����j�Ғ����u�� A�~v�<`�0)�R�>��!fk�ˡ˘��f,��z�l�UB�,�y9P���w~�I�cv\v��9@Y�����Bh�B.�Z���!��D��9~}����.�s�^��C<R����jH��5���R	n��g�y����T��� �W��ꐉ{�έ9�K�Ю	>�N�,�c2g]}�	����㓳��3�2�g�X�!縩t��ƄPc��K�7ؾ�#�9Lz��ޮ,�f�l���wOY��X?d�H���DF�"�����d�j�}4�i����w?vS�p�rJZ�����b� �(���NθPn�yw#Dt�a��8$_�Nwn9x
X�9Q0Y���/��DSU\�פp5gn�z�ZPN䧅<
���A��(��M&״. m���+M9O�VU��)y�݌�Π:B�P@��=q�D� ���h��I����{b�?MY���̣Jc|f="j��Z`�%�^o X�X����tG��a�zR���*����d�i\%��j��
؜L"���m�[�3�4
���=�e^n4���5���3�d��������\��  �N!�X�SK����-�D����\}2�OCl{Rx{�sx\3g]�ݺ����X���c��P��r�v����Ah/HN2�U��{x��?�;BF Y�����pz��<Z�x�Sy+ə��VO%���/cw�T�#�_4o ����=R&B�dª� m�Hq��}��Ο�sK�,���2S�{�^��h<�]�pk�Í}� �^��,��8iD�6t1W r�O\����(.�͎��v�S��ʳp�X�9�䱆Vہ~�A\�zXo�WD/����&���!���T9��U�
��G&��BVh�)���c͂�v*\����6��r�"�W����d���0�F�ooe�r��f�Yz�C�ɵR3��E����DB@��RK�m0y���G�b�/X^}H�-�{4C�]���t_��Y��5v�۞�I��5�̈́ �R���k3,W&��d���Ҡ���sJ�Hx��|W�/A#���¡-G�
UVʌ������a�.gf_{{GH���7zXÅ�u$�C�N�R÷P�f�Yi��x�Z\���0��[��2R����]8�z�и��%É �k��"��EU�� 7k�� 38bZɹ�\a��������AcJ�[�n�S&���e��F�H���%��A�Hވ<��oF�� �#�3�$nW_)�	3j��w���{9wL�p�<�,]����o1�Nf��u�Ł�����C�._�v�sY����7�I=۳z�{!�j�81��<( o'�3/w���:�$��u�
�z�����cV�,`�:��7e��R�Ǭg9(j���
s?p���Ip�ˤ#�Y_���=���o�D�cϚ���o��^��f�d�/2>hi�p#�@��l������.��>�Ű�(QP?��B�>�c��C?kdy�c.��X�os��zF(��9,3Df����S{ ����t���I/#u�(\fG��L�W��+)N"7y)&��A�h_���<yʑLU'7%E>m�䥭R�)�&_���i��5�q�bLhW]���dϵg��_	�_Xi�{�W.�&��a������c��~iJY>2�����P�_o�7�Z�l#e�O)�9�s�����Dv��l
��`���/�t7(Mþ���~�o
.;$08�Am�@���h�p:���	Q����I��ϓIh�Æ��.�� �k<��ܔ%�:mRDp��9�_[��֦�J��bRES�i�W�L�O>���^�jLT׉�3�t>n'�7-�a�LN�b��7��![I�x�k^8��*��:��4��!��&ּ\-��Z��j�y�%>�ԣ�:��ro�G0X������Sr�r��fHSAjCK��(Z�7�擥ݴw3���rHqD�r���p�=y�z}��q�宷�z�T�6^"w���4�f��?��j.���뮎�Jې���F����ib~\'�}�y0u9%ȩ�b��'+�/j�"z�.�-�U	��>h��Ҙ��(Շ�6tG��&���_y��u����Q]����0����d�U��ۯ����(���"�={K8�y�S�>���!d��B��)}���+#y�������mT�G4��~.�ԏt+<!3�܆�ŞH	��V�C��V�E�e`�}5��k�9r?,�/|� wr9I��B	5�=���:KA�K?o�=�DAZB/m�w�jT{�����?u�if�#��qկZi�j��ғR���`�,>�_'p�����W-��2u̿���� �1�>&7{�=�n����X,�Si�����%����r����6��Ye��.����^��S�A޾������T
�0�y^��һ��L�/������5�N҉��bP �,��e'��~��f�ߢxF�^�&i�H pɢ��ա��aP��p�f����Q�K�ǩ	W��s<\V�w�����^Ņ��b{�����S��q�4���_sҰ�$F/�J��p��E��hQ^Y�.���M-U���s�Yf�|�ޢ�dIQVD���;�2(�EwRU�Z�x�R)��M����p,�>NiF0Y�ި�V��(n�����ʈ���<し8Y6�H�A���`0�j)w�������bm.���!o��W3�j?,�e�!�v��v���߿��vp���O�xH2B#����r&��E�Dީl�{Xh��M4�M7�ٰ�,ˡs�l|M&��z�Neu�%=�dkF|��^�*{T9wL(:�v��i@���v�hYi��$x������-�l�a�p$0�vi����\���,7�!��4 ŀ�Jo`(�o����[�
H\<Hu�E>��r�*U�ZgZ%y���>��|Q)S$崓͏;S�c�����a�93{�%�����[nӛ��8f0I��|��b+/,�^�K0�XG򻠴t����5}�\o�7#�Δ��s��)Q���$;�ZE9��pB*���[���D����J䒦��I ��ر�\պ���wR�����}����>=9b��s��?n����^�c_��Ŝ�ͦ��WwAub�
��h ���^@д��#�ŎF�Z���f�J&�ml������RӃ04��<i�G�\��T9a�%v�Xi(Z�m[��^c�sN�j�+Q��J%�6hH�z�? ��Dy� ����Ǉ�qq���i8����6̆�G3�[���h�Q[H�����j�@�؆�bw���P�N��A�����z#p������p�ρ��\�]�^yM���@�+��1ۑ��B��|����	�>:8� �7���NÃüx�KY�8�202@ C��$�&�s�}�x��9�%@������I��p	_w��I����ل��x�T��� @;9`�>������WDX3d�4��k0�y��/Y��0�!�I��*�A�]��w?\��Vņ�+�gg߇�0>&rh٦{4�!Æ�N8}���KV&�:nzz�W�!��|�ʧ��%/:j�?	Bm�Me�`�O`��7>�����Y�	���1����M�����Ö;w�����Ԧ �
�@;1�_�y_Al����I���n&�{U�z�!�D���ŋh1�>���~�I�'���W����sY�ep1��U�����#""�2CL���塕���]����Ac}���|ȱN&��rkxݎ�}?2�T�:+�����dt:�O�|e�z��&J#��+��&�R�mF�'������8ぜ�ؠ��Ғ�&?7�(��ջF�q>��W�W��7v��$�Uu��Yw4�S�˙�e��f��ZgV��95j'���󱛃A)ԩ���H�U�B�*�ٕ�z�ARz+�+�m��1��srWߚ��@	�}%�"8ZR��@Ym&�����V- ��	Uys$�����õH���W���Nʭ��E�ƻ�4��ؾ�}���rU~w��f߄w�l�hFa��~�g3{;�ԁ��r���߯�B���-aV���Y;�6J��t�C��X��B��-�Ӗq=��|�eY��Q���TL�"�d/�m�l�Gt���(��	���t�����}/�4M��3��M{�*ngϺ��������0(���$Ѽ	�|*�;S��F�覉o΍2͡a��S��J]�>���uQQ9[�G�Q�w��b�<hR�X�c��0�����Uo���lMa���:�bX��jz�/af������2��j��m�ii=�J�SÑƽ�C&E������]��
Tq���v�&%n���o�VDw|�� ���xAt$Hb�!�_?�q�{rU�;>B�C��g�`�b��4�RT��\~?�3~�Qd�	�.�w�q����]�v�NO;�5�>��*��ו��	Q�����ʛn��8�ӕe�W7F)�sZ�vFZ>�d�v0ҳuҮ���W4���a]u����g� Zo�{�M�'��u����X?����^)��3AQ�"�,��R޴��	�A���_��N�7��6ٜ/�-����7���7d�X^�>�
�'��\��`�i:]:i|�\��x�������$�������wނ� 8	Cr��8R�t y����F^k��v�gZ��6U������8ҧ�
洤�v���i ���"�XG�
Ց����/K$zEܿי+�^aȿ�(m`lbh�Z������(��C&��g��Z����?�$!�?��,5i�HF�r|�B|�x>�2�'�:��2Q>�}L�����F�?�g	��X^�����	X�.+��$��ڠ���e���1��]���n�"�L�d�4|��8,-�\4�W��Yv'����@c�4`s����3u+I�S�L8�o%�]��li���1�l��e����*O,m�;�+�]�n�����
��j|�`�e��W�qIY_#K��:\�l��gUf�`��S�&gI��`7���=���Yd�+�npf�@ĕW p���M�乱.�[�b��Hx��B���V�yK���֧-�b;S�'2�p�U�<�`+��<�[�3&��&�( -����'ÄmY3�F'���P*�|�v �4u���T��=T�2`���E_�R���*��3�wwjQ��s�-���вLO-�1Y&��5��Dx�0�Q�:O3��*�"���ڌk+F��[ekb����r�r��u� Ŕ�t���S,��
�^����.'�"\,��ڌ�u�����K��H����RqaP@;��z^��uI�s(�_�B;����_�"h����9�>��cD��,&��JM�\����S�6$Na4��N|P�pg��*��fb�B�=�l�pX7�sW8�7[k>��Te�v��B��Ӧ��ԃi�?}$��B/�$G�>����BCK.?��G�N�7�H�����/s��m�@��(4���0GkF���'�w=5�:��&������D�ard�����b�=��D鏫��?M?�V⺜�q%2��-N5ċF
2"����DZ<<+�}_o�}�>���P��0T�"�<Ԍ6��FÄΚ{ôMeƄ�7e:����x0 ^h���@��m��	x�ǂ#�. ��y9�<m
�ԙ1*�*i�=������9p͟I���Ѹ���l�o��&PfE|Y�)�	Q�τ�$�� �*�fz���;�^�q�(n�����?����W"���NJ������e,�Ƨ��2t!�=뉄�9z�ҍ�?Wc;�	��U�#lPI}�J�yV����^�@9��@��N�����u����CJC��Zf�V��������[��ڳ#hMH��H�Q�;����D�市:��Y��$6$|�Q�㰈�/"��l�UE�������ٶ�`[�����C��������H`���+�p�Fް�/�q�Δ��w4�ep&��x~�j����hu�q�X
��1�����*a:��N�����D���=J�w��c�*�#��v��f<���o���5�P9��.�U����QM �jg�>M�,�����=/�*�o��û�`ܐ�A��ZC�@��8�Š+@�`��c���� ޾\����!��]�/]�o6�CR��m a`��PlTxALsN#�=<�1���� #�}�N�����sk�p|P�J�vm����=�!L��vvy��EՂ��pԱ�V~�@8A�;|3Q��*e�3���qTt����5�H-�oӊ�%\��~(�%q�QAڶ�S�2>��o�����a��8�IM�C8m��J`�=k? ������%�GS��}�l��f���%�.8n|�_��y},$x�jC�� �Atx��Zժ�z�0X8��I�?¤Ji��u�"�t�r� AZ��h^�f��fϢ?�d[��^E����%���%��3�a9o� ^&�~:�2�:-8R�Jt��y�b|��}[�N����"WE�R��T�g)}�uݲa��"�*�CS�����P�>!���ǉ�+�<���	p�!�/u��������H��	�����A6K�~h"�0K���J�l7* 	~�1�i���F��s�Zai���N���ҋa��;��4�p�i�ٝ��Ur,���Q����l��Z��Uu��1��X��Z7>6��7�$��s��n��͉Xį�@���;�XfM �P(E�ܣ�O8�n ���X��S�w�_�۰y�r42 ��v<.K�pHr�efF��tY�pr<��(|
�7;�k6�������h�v��8��d����2`X���9l���u
��a阿�
��X�:��)�.���lT�͐�7�gSg��������F�J�I�.!T�P��S^p�z����')��y��V�� F����^����������~;a���IYkG�H��&=�G��K�l�O���'Z�$m7�ch�4�kw4v�1�˪)�4C]�q��M!�Phx��
��K����]��?�6Y�P�r,�c�F��q�����B�KBoH(�v�\a�D�ѱ��D���Y鏈@���C���2͵�A��U���aϩDqb�%X�?�CK|�/ѝ(#�m�<+	���}.t��WB~��,�����g4��+,
09�W|I��a#i�'X+�{.[�<{Ⱥ%#}�={�q�:W�����AU8�*Z@9��-[]A�?uj�w�g�����t;H)�)�_���G������pg��}�OL��Q�c����ǡzO[��?G;l0��)Q���F+�t ��^6��o�H3�k$�r6���!�¶��$�Y�I�Ј
A�ԙ70t�~�����S�R�S�"��ΈL]뢍7Y���t�H����L�ҿN���տoo1ޕ��� %�y�
G�˺���{zO�4Ưz0o�E8A�-��ޮ޺J��_AIe>��f�^_Mޕ
V3�Q�~�ވ�sލ=�_�VAu=��"j0�f��c��|�D��\ţØڱ�ɔ�VzJ��,�W<�H(s��[O}����7�����d��Q�#�o��5E����~0R����k?���-�2�HU)� S+C}D�J��Lޜ�u佉X�)��%��m�PD��h�V��Zu;�tA(��6b��N�va�d9�����`��^	����AKO� �L��-'/3<�2oA\����K ��w�p��8ѣ�={c!�Gv ����e�ջ�۶?�P�aWr�0���wQ����6��&N�hx*`��%��d$��^��7��,��fv~�-�G������C�a��
��>�@�9�t_��љ�l>a#��������0a�H���:���J���C�Լ\�
�S��6V�K�oo�Ԫ&�V��qd�F�P��7�z�#C����w�4?50���P�s6�I^.zm��)B�ʔEv	�O������h�N�hT<H��e�a��I���r��Pѩm�!P��o"g��;gl ��6d���(%�aQs�8.T)���/�<�����o�с�ah���J�P�aנ���kkK%��z|�dvsf���'P-!�,�@�˿�\���G��*4�����]���	a�յp��U"Z�
����3P^���KA�kBZ����������o��t�7����rq�̆��?2{"�<bpU|��=��DV�sd�~B�a|����^H��Y��Fd��e�N�?+1��u�	A:�c�Jv�� (y�-��-z�^�$ZA=Q$�6h0����Z�8�����;!��*�<]
B(WOE�\rB��x�@b7&������8��?:2�%ڈ~�/2�����8������7���̈�<�O� 诰��Q��x��׊;X]L���^�W�ݝ�#j%�Q�����c��I�����`|�0Cˈ(*�i�14�?�t�
�8�x��<�/��'2FxlF��	Ĵ�ұ�mR���"�����9FBflk-F� ����O3[���/_{X[�`�(��i��w�>j�3i9��@�����d�f�����NC��+cv��b���hj>z��3y7{`{��*�L�RYJt=�4$���bf9\s�\ݙ�>���Ϥ"��vS�89.��<���r0�k�:kI����?N��l	����C� ��6�Mq��+�2(�6F^Hi�yOVLi���=,|��l�	��&|�3�0��޿i@��J*��
���ȠU��S*��R�p�!eS��e�~��-	Փ�=��a����MO�����@jĳ���+�.�p��,%���G��њM�8��'03�<F�Ka>���j#Â���d�Rݒ�(�q�v+��zz�����t�w;Dw
�&��C�FV�lĥtjC8I�檉��7V���y��Hd�3D���e�*��=P��c�q�W���,�I�(��$�Ko"�������O�)%���J����Z�G'�ۅ���.ov�PY
��KC�9l��)�aEYZ}r|$�͙��=��!A�8ї�{�:w{�I4.�~������{W�=r �ڷ\\OM��X��~�����Ɠ�`B�_�k�'�L�i�,A�����TśE��zƃ0)�� ����_���o#Uv�Ĕ�b��a���<�t���p{�6��l�oc���n�׊�� �a�� ŭ2�!�8�d���
�2�lgz$�TeG,�vw��٭���٠�*������Hz/52�������������i��׃˺�#4��꓍�����3�q8���kN�$�{A�h��-ŋd+���^>�0�e�
�[�TW���EN�RR$�Q�ve�ܣ��٭�v�l�U�ƢgԘ��/�4^q��@����ʦ���f6�	r���&ڪk�K����_?c�G�4��'GI*L���Ⱥ�>���s��8������&o�L���ܲ���q���{����0�i����i�@�>�.LbZ�`a︮�p�0\:�z�Jyi�����+�0�1��4�d�n>�㯎
6�L����K^,S�|k�#���л�E
]���)��R�q'���H�]�� K�6m�ã��	7���#��T�ߏ˄?1��'IKw�þ�[��\�S���'eq񋁬jq���Va8���h���#�R�ih�G��gZdP&�����-܅�~��$mG��N����`Qsh���hs��H�ئ��:hs���?ebd7}0����ZtU�A��C1!��d����7�E͓$����?�� ��V�ki����|L�:0�OQ&�W���&��S$*��RY��62�f[�q�^��)N�Wg9�#*�̳��TnX��5���/��>�p̘�f�\����b�MN$��kF�T\A{ɘ�4w(_�eִ��4'+[h.Q�s���9�WЭo����d�j󵝋����V��\�Iƨ�5 p���~^��I$W�����r���w]�ǉ�?�YJ�kt.��r��ϲ�m`δˬ��@����N�X�)�Q������$֮�=�K�خCa�����AQ�ך�`�u��x��_ۋ�h]�H~� 5�W���~���vh�p�
��%�S�E5řs��m�];u��pM�a��!�� y�%�,+-n�E��\I��� ��2�7 �?,A~a��wU���d-[�D�&Dsq��*Ӛ�_�_/��}��s�d;*>`N�rrƳ��,�Jf9a��90/gy����C^$Y�i��p-؎��K?�Ơ��Q�*96ˁ�� #]^�J9\u��� ����N������1(���B�i�#��p/ji�܄��?X�-ߥa.�J��_��[�lo�S�U�t[VW���>T��A?��g9���������1q�&��0B�wt�0V�·���1�O� �w���+���*�nP� >/���ro��� `݀��JP��47�.o:k_���dݿ4 {�E_j�����b퉥��k��I�^{�@��=�3����#��/�4O����`q�g-�sΟ���&�01�k�b��h��,ᝦٜ7�ey�)o^�8���cNׇ�s���Y�5�Ǟ��N\e#kb���; q9�@ �8�lLa]�G���o���@��M�X��}�^�kc��Vz�RY���O8��;i#e�$�����j;^{B). �Q�k���"������Ƭ%�
�)�U��[��������/�oɸ��F���8��\bWG7�ư�7k"���oR�Ŗ(D�4v/�������wP�:������[�ڈ��:l�Kg&���Y��vj?������FynKtw�Tnje�3��(;�͌x�d�ry��Yy3fz�@),#.�l�q��`�K�{��|�X�����2��T��ff�W��M�B�i!���6�ϴv�	��/=�t���a�Tx\�.T�Ή��kb?� ��u�3��ql+c"�P�u���f+l�}m���l�yME?Z�"6�&α)i`Y2s9�(�K.pz�[A܍S,TQ�F��7M.���`�����<V��s��7��ѡ��$�R&�ݗi�z�y �r�`��%@ɾ�����R�d�Z�Z����{Rs�Ͳ�@a��U��~?su1W�(����1���LP������)1�#r��S�im5��������Z
,

��������ur΅�^�]�s�qG�>P�vySӹ�e���w;�ϓj��j�64K����qzH$)�ZDs:�{��R��'8iA �`B�����D��F�L�%��8�
��9�!��/��Ґ��U���9p���O�?p�m�f�S�oՔ�ٟ'!J5�n�S3��==�C��u�ZGQѪ�w�ձ6���:g7��h �V=aY^��b;�� @e������ �ūJ���:մ�ӭ���("fX�VuS"ǚ�$��o;���h3k�	ءa3]h�}w|�ǜ�V�.[\�S��~No�=�S5�My=�7�������:>S���b�3y�s��������tp�&��d��|'|ڔ��_9M�P<�b����]�����7�B�%Y���
U_�ج���4"M�'����Rj� �������Y\��O<�Z��(��/& ��k:�ɇ���)s�;p5fS6����:�ԬQ3E~'w
j��
�P�<���I�+�s��o�.��-B*�\3&
�i�PU�MAK|�:n�#]��I#O��7���q`A*g�S0�U���q�z�Ǧ�@t�N2������d���S*�0]���� ��M�u��kFZe�7�%��'�B��%)��T�+2�|H��V9r��,1���;P��q����P��͛���&�L��,R�߽n$:���Eq-[�*,.�1��|3��%`����udp95 ��p��p'M�7�l_p�n�}cx]�e>�N��F�oYq`�N������Ҋ��m7����:�rƒ�o ��ᭋ �}v]SA'�[\'��?C����B-3FC!�Z~��$��Tg�> �E>�eKF�]��+���s���9ͯ �w���E���H8�����Yk��@,�׼iQ2?g�8?J�zEj�0��p�9{l��#m��:d�YōQ5%��J*4�!a���t�hD�k8�>����6%�����)���^]ӡB`Hu[Jd� }|}���9q��x�zC���J}��n!���RY�=��Y���d�!w�I!*�R��k�",�x�j��;��uF���Y0�2��3f8x���GR�=re��d�RH��x�
׶�n�����E�q��֒��ŒW�~]�>#�J��pp�D5�W��i���������=?��۽[6�Pehy�
�o�iI�"��`b%e��.����b5�Y�R[NH�S�"�-�̦gW�aHo��D��+{�d� xw��|��U�c�o�|S'�>cLB!���#�v�[��@�# �����<)GJ��|���S;j_~�4��BQ�_7��0v=��ҳ���C+$]g�����ɞ��ޜ�������941�3�A��k<;i����
�T�;��y) 2�^UD�e���
��>��|i)T��e�]�(�n�*tK>	k�=�iq��zE�3��M������O?��@ �S��	�E�\���I���������r�
��C�E7��9�g�����"�,3q���,Eջ!)={�+����d3��{��C����ZN�6��?x��^�>��4�\lc2x�>.+� =��'`[<�������ۻ��G���	��������A��dy�eP��/�������s���
6�^���N�jd"��$��H_�%�_
_�s9��F}���)�p��^�
F���c5��"'�������4���������s��_���0�����d�p�:��hj5���һ�&��Xv�F���10g ����OUl�{�-o��_����.��8>���&$ޭ�ŉ�=��6>����S3>c[�B�����8��:�F���B�v��ʔ���Y�7���3l"����۴����Xg:�ʵ{[���'�;��thzi?t�![��,�W�c�Tg7�t��"�^#�&T]�,�}�fkgU��[�Q7Y3Z�H�1�:E�]��|P��d�f�̖���yU\N�[N���ŀC�D�,��YU��0�I��:���?�� O��ڠ��S��yhe^?V�w����wJW@�J�!�Uq�M����+���)C�톅�M��\�ʶ�u}�E�	��}�{���,Q]9���k.!�ʹM2G{�4{6���2�2�IM={'�N��b��C�U:���$�4���@�<��ws����t��>�߯�x�}��,!���#.���*�'��W�
�K���л�(�hi�<c�hL�ԙ�!i��a�-�3[3��;�pmX���D��$���*�m�C��[넔����|��O����'�����t@�����+�-+�k�Fu�P��7��/�&��0%���*_���83w'Gr�VE5b>̙|X*���5��(�"tfG����������T�<��;�eV��Hj�"ki��") y.Lv8�Y�m}��0��l��.îo�4��NR�ivs��	������'+��m_c�;k~O��p�߹�?��U������Q#�W���R���X�j��;'h퀩�k�}�Wޕ�ް��GZ��9�E<��o7���_�m��ḱW�[��0e��F��¼�J�}7K�|�ʒ��'�B�&(r��q������ck
�4Rf?l���* 3�ɟū:��ZK.�m>I_�Mn�O�)L=��s�Tj"�:Dg���5�����@]X�f�ݎ��;�-ˢg&�%j��dU�ƅ�H�X:l�g�8���sf|�E�Sv��ga�F/��f�0��C�t��)W�����a�n`{���D��)CU�����To����s�pUx��-Q@QJ{���ם7^)t@�+�A��v���y��K��w�nt��?G9��v����g|��^���RS��\�/7'Ѹ��g�b�&`�����	f##>��V��K��Rc]�^g����LT�ȞK�oA�%x@!��ɐl��(�# .�.z4����x�\7��fC��O����������/Qy[�3������0#�8n�TE�\~G���(��F+h ���^�$�6z� ��?`���1ũWK�!^ny�x,�
���>G<�LT�����j�_G�R�M�ǻ�Q�B��#83���Ӊ[����%�4J��O�+ȟ�l>e����K�#��:1ܽ�㢛i]��(GQ1��w�~\"�t�A��&+���Op��\J��{�ҫ���D���Ձ.�;���q�,��Cǁض�@��F��I :fmS�L�#�O�c��N*�?,�	X��5Ψ���P-�d	�qQ�1S2�DT��0�����k+�sd���ʶ�v�����q�+�"�x����'��k�%C ڣO�J9���E3F\�m�bj�M$3K����^@ztr��tW�c����x�ͬY��+D��c�������dH�~��EP2�N�3����X���KYm۬��В�};Z0BCr^Ok	�'�aW;�"Z2������=)p&�hfM�2K��@�֫m�ZP5��o��p�����2��Y�\�q+��ς�Ŭ�e��K2��h/��u3��`��:�b�v9�1�䋐"T�N����k�s��&}��"�x�;���P�`D�<��!)��?}�|Nwa!Y�c�������61\��x9a���9��X��&���Q,�M�z�+���Ew8^�80"o4�5�|faѬʰ� &sO���6Y�T����$��3��)����ËńKE�@ܓn83}�,�lE���eB�X�P���YC����Uz~}&��4uf�"D�\�htMK��@3@�]M�z��	�Icq<>S�'a|�_ρ��.�+zA �~4�z˽VWh�*D�#�� �a�@�����P}��f�淙I,�H����o�8�e�w=��c�~�ėxmIc�q,� �ҟXY�,�)�(t�xN�>����p����1�w�Ĺ�O��m�C{ҝ�+�p%����n�h��nI���5+O�c�/�YB�k�b߭<���K�Y�b�c�jrLz������k��z����&þ�.�����om�h��m5�\��#�CM��K��"4�n����@�g<�ޠ-b��3~�~���Z�E޸S)��r��K��2���J>���&dK��T�wv��Z��ǆ�|S�K���<K��;O��y�?e�� �}��`���c�M��v�P~k%�n3
�c�6��ۛ�l[�pw���o����x�ކ��O;to�H�%�%ͻ�chsƖ�c�	�}�����@{������G��N-y�6��0�"Bˮ���`��ǅ��`c#C$�r��zX!"���|����J�q�}!c�N�i$�=�@7~U����a~�z�{�ǈ�K��F�U4a鵴Q�a����\g����G����Z� �O@9ɴ��<z �Qr>�[��ѫd�"��4���O]-�!��a8����j��e`�|��
�)�{�2��^��ہ�7<$��"3�Qh[�>Q��_H����JZT:Z���Q�� '��ܾ[2�6�|e]a�UrДL�*�������MRm�,�Dy�II�6Y�h� |D���m�t�b�ͧ"o�r��p�~M�eKw����8��52q&�)�:�i����a��q�:�,� �+�u�U�>���N��7D[0�a�!�u���)��OL!���jH�3�+���S���֑{������"��X�0����shf�\��{��^�-�'k9a��L�C=T��������p�]}�,Dx��$24|p�/S=[��"�����2Y���Υ��m��,��d0�\�d�K;�`���=2�S�$�dQ|��e-qJ]�V����)�][?��z��5�-W�K�0:䓡ʑc7g��XF]͒�߮��������J�2աP_��ii�6�@-�0��<e@B�Io��Ui�x�|V�iz�U�x8�o�R�O�0<�M�z�2F���m�V��Y�����qy]�m�xb�wl#"�wM�j�|���1}ǫ�.*��ʧF�X@Ѥ��PW�K��.�N���@s���ǅF�{�=o���q�pT��]>Z}(�y�'���&!�g}b�G7d�l�1(6n�S�͙�#����b�:*>�e�剫�़��}�@!8O&jE�#{/p�
��-H~e�J�x+�`�Qv�ØH�X���X^��c�9�,�W��iE����k=��{�g���е�q��s$=���>5�Y�>hT��u�3����ʉ���"�Tq��k5�L�j�䳦�7�]��D�|���^��ﾷ7�R�W�2�MY:�2Q����Cv���Uf^-�E5�@��d�G�s�.S��ibe^��C��e%���x|�+i�&i��
�wS������P�2Wx��==/2�	{��օ�a.�ʝ�s���n�A�:%���W�Χ���A �O�Cd���\�siL��}���O�MU��I;�J���^����$��i9O4��g�ŵ��J�,�^s��s�8�U��D�Ǡ���G��3�wx
\|�J4�-U�H,���ǵJ�#�A�>\��#.z00�C��A2/���(W��Mxr@)amM�(q=�e�ܱ]T�HD|��D��b�Q�Ѷ�n��q�p�pB~��V8��B�*�5_�g���P'�/M�ບʖ����D�f�ck\ �6�X��#wDZ;��B��q�"u�r�@ �-|��FL�-�R�Pp�ȆX�w)�ٵ��!_7�t(g�;7J�,�zO���ً�/��!��D��3ӆ9PA�]h�k����̤^�s����i�NG֢��#"�F����aBԸ������M��p��|�$�.�2���+��y�Oi�Js8�E�;�e���w���l�L_���i"��>�,���N�Z��B[�j(��LC���eJ-�Z	�f��m`o�}!����p;.��P!��w
<�n�ܑ�qK�DW�_O�#�w�)��O/�'o��c�Z힝02{`��K��8��m�z6InFˇ�I���>z�A�
���BA\�ylh�[�s<�8V,Y]-pƄ>��rO8.�B�ȕy �,�j����=̇BirT�)�P&�+�u�"���d݂��x(9��T�5
\���za�ȝ��s{0�3i�s�	\Bgf8nb��F��!5Ѵݔ�v���L��K�Ǣ����oF!Q�? ����=��\��Y@�%���vu�E,���yt	�>�p�W��[���A��ƨ�7�^A��S����ȕŖ����7DJ��B�L��?�W���c�[�bP��@��A�OL ��E����V .S5)xd�������<@(=М�!Mlt�M�!���sR��NO?�.�XYtM����@|jJ5f���N�����_���0��d���������+��Q�^�n;0���m	یk	@��$D�hdW��n���%mQ�6V^�&H�M\X�E�ɬ��tvv1���۱�I�;Wwn��gS��Tk"��V�5�Ei�
KA\]��M�@�P�@�.��i:�}?cT�j��gTƋ��J��6��`Y��R"�mG.�?��ڬ�Q��������T�m�ɘ�����)��>軪bG�NٖU���j�l��Ϗ˙ �#�Ł���f�$��:��fsJ�Ԡ˺�K昖/ �h@1�s��9,c���#��j5�Pǿ�d�v�WN�\7 Nv�RϻC&��J+Lke�}�.��3�h��]��ߋ���́ɞP:p�AX)����T��+%6ᖟSޤ�]�B) `6�(Z����|�=���x���ل�,�SJ�wk�B�lW7Q�#�v�Єmz3�4Lj2Փ���$̃{�Y�"\T5*���#��iN�샜�����d��P�ꭰH��� %B x��bg����Q�_9��
�������V��+�6��e\�m�"��Ub9Կ%����[�d��)L�yfke��5�`Ͷ�����1HXR�Ǡ�6.�p�J�-8���Ҏ��^gg.��+�z8գ�:W�;�Gr6�x��hU
����AM=c�W�I����O ��d�P^;1�N\����6��r�X X�ŧʞ/�Wv�ֳ̛3��F.�54J�����P$]�9�7J�t����ԋ�G�6O �I�ė1�"	6���u�JqMڙ�<,?_0���xв����S�9�R��4�k��!YYj��>|YX��/�����ة#x�D���b'
�$��� O�v�Y�_$�g�H�]���S+�!c�I�L�G������NsS;	ǚH�L+���6`������Z�ɣ�0��,���*��H*���1�$���d�)��v<���RG�:��^S*f�oJ��Y;��m���)�� �%|1ԋ�i��j?حؾ_3��'B!D�.�w���f����V��e��s� �.�u�v�O�@7I���A��ߤ/S�?Jx���z��^����u� �lK�n�0�zښNfT�{��K�`8������y9ow�;X�g#�ْ٥���@v��B�����47F
N��J��b_C� �m����,r�HMm���]��5�Mm���f��11ж*����*F)�$eo�a&ѭ�QEu�r��)x[P�#�2�ˆ�-z��=�)yfFE0M� *d�T/�݂N�Z"`.�(�$�aN�10(T� �2��#l��o���֎�l4P=<�7�T}�!���M���`I�~�4��xp��Ʊ�`ua�ocɯ���n�,'[�{��[�5��*���۸P����5	�d��01S+�}�v�/�����+����'��K�Y�N|Tu�h��V������G&5u��m[�i��\,���#;7�	��Z>�^��%�p̵ 5����T�.����#��7��l,�Mi(]��U*�x���]X��ܕ�
�7����~$����Au$>����>�ر��-��qX�%�s��3�.|/\�l��9eR7F���䦦�E�a�r�7�|��v�ַ���\�r�����b�Tb�� �%J��C��e�~��ozO�J�b��[���gr�xjMm>��o�m<�j��鄍+�p�X�)���E����qYD��U4 �f���"m�`�V�}�P�$a�����Wq>�ݭsn�N�*j�.\��(��m��?B�>�7�8�Sw�%���)��{8MYj*��y��r�Os:!b &Q���L�]�E'��Cd�,
�xם&�O��2Usxя'���5u�ޕsl�l�y�Gc֖�܊=p)�T��w�Tnv�Г�^W����E8�]�	���].�[�g�AW�zb}�1���ݢw���_�p�5�C�C�%�f��jn8S�N�j�t	Wf��逦���M��G�)�D�T2��\`vf�� �jO����n1�awx�M�1�~��X/e�,,�x��F����٣�?�N)?L�c��k��!���S�N颻�������rk$Jm�ԏ����>,<.�*~y�v����9�����t潣�'1c�*=ڢ�T<Ÿ����3���U�	�L�����U`6�L��⫖�K��n ���鐴��B�y����qEFh�rƨd��S4�m�S?	��� ��բ{Q�R�[\�Uf����*��@�!6���������c�����g��+��B,��i0V+��!�	����w�![+�&P��mQ�w�r������4rx�k�7�Rjc�$�v�4aӹ<�Ho�_��[Nk�w�@�%��1T�A�׾����"���j\�b;� /)<;����6l��֠����2��bX1��"uZ�}+g�7��tax�����������O��^˵�2�Mh�&��Iv�1�(�9���*���f�{�l�O"엪m��ǵ��?)��%�f��<�RxC�Y��)��r<��n@�g";��lll)���ŕ��+6�Ԕ������L b�2������h��՝5n�#�F�+��/�N��,��$�wy&�N���y�����.OXB���P� �#:.���*�k�f6�YoQ(����_E9�XL���F���4R���:��&a��������XQ纎!=k�=�6�T��b��F cp�GJL��� �T�����
x����Lw��*���xye��Oř4[p��k�/ܦ��kا[���w ��W|��]�ֻ��(%[�ߺ���y�Hdy�Ch����#8��{��u�8�|�����+N��+�r`���H}qyp�+���rq��j��M�:�Z�$�5�$�E}n��D'��|Ԩ��bAr�d���7AJ�*ץ�U��A��=\�* ��V�vh�� �6o{�9󸛝|)�Т��_�66RiQ7�T���q��c-|�.DwxG�M��hP�%��S/�]W����ܣ*eaUR@�Z�"�[2{ZmLCp`�Zs�R���)�#���@,�>j�%%�.��8bm��^�`&F��Uo�|(�Ĭ
��������n�[s�j�<Z���
�C��
9�YEiǎ0��a� xk�}���A1.�NFe��f�%#�C� �d
���K�`���.2���m}����{��q�s�{1�G���^-����"��o�f�{��`���[xjD�.ӽ���=�=��-�nA�:.D
י��vn7�c��>%��I����#5��e�T��n��U@���/���;�A�}bf��z�Ngl��;�M?�/R�!��޸8x��M�AVN ��b�E�~��y��[��YD�/�K%]�Tzř�4�H����H%՘��^D-��(aU�j�w)�:�+Be���uX���;��\��*��64칐�m��L���*�Zy~�c]n�
NB�������6wZ���ۼ��Q>ƈ�;%8o�Q�d�UX�U�
�`0�wVM�,�����L�Ii�
C�W�=��"eX5=�(P�b@��������L�����	v��T�K���{�����cE�H6j-Ud�F`Ie���}GNL��gb]�>��0�u�xO3�G���G�hY�6ћ�zx�ܛ6�z�i�(<����Ƞԣ���\��c����x�hDI32F gR=##��r�Y�  ���7�Kۣ�X�[f �n�Չ�:U]�5�\ȰV�%x[�(����mYŔ���R�4<c�[uCV�+6Qrjd��4��?,�F,[���V};?TPp;۶v`Xe�a9�����%DkG�C&��l�P35��~|����p�3�}�T�$e���y�d��)�D��|Y,Uq�#��<�J004����0��U�*�ߔ�e^��t�W]��_	���2����8�_l�ˑ^���nOԾ͐��R����/��������kc�����K\p�,�1��_Sfz�	��ܦ�����f� �)F{"f
u���%��q��qM��a�0M��Hcx׈������pH�gt�k�gLo��6�S��Y �-3
Y�6��mG�s�˟��VR�\b�W�WY6i7�E�����R�������K��q�f�f���f^�aS���7��Ģ�D��l)wO��5�t2١�E��t-b��Q\�үe�?gmZ���iYUW,����1�z�>�o�Ԏ`�\��j�`�(�g��6z�R�}r���+��t��j�ˣL2-��d��T
�+��c��Ѫ$1��C�k+�ͽ�T-��Q%�,i�`!��f�#J��È)zڜ����c��:���dx�zߌ�g�ws��܃���`�fY��*!��95a�5��+:ߕf�;ڵ}F}h���x̯־�Oǋ�0\�`���nvb;P�U_�@�Fz9��Ψߌ$���>��Ǆ�&@�s����.{��J�1��蛬��������b�&�nD9ʲH��.�-�a�+NS]�`� ���}ڇ�jg��z>��B'_%;���$�<̕	�q�E�R�����D<��`�V!Jjh��&3� �׆|o;ʨ�*SX��=��F��+rկ�`FS%<B����{|��^&a����,�0%���W���W�N�d@@=�)��Nr{���G'L'�d�EW ����Ib@/��p�S9��0�|k�lwn#H����ٶ��%��eIv	�wǳ2Ac�I��{E��	��_������I������E�(p�G�;R��i�A.�A~��܁qXϜ���e��s!N��<���u�m�kt�Q=�k�!��H�<�"P��8K�uN�Q}�{'k�����`wcNƸUW�t�����>��ҢL�a�+8eN��ԭj��8�z�����S�Oj��r9u��{@aY m����(��2?8�5��a�ۿB��Ė�)e�����P#+�-*���<�<�� ��S��S.���Dm�� ��>Y�kǖj-?�3�xwT�ϳ����M�_ �o+'.j���;�f#wQa�'��0k9TM��Á��ӿ�l�+Ω��[�P-lD.h�`��"����.�9��y�ߥ(�A����8�%%4"SmM�r����SQ�W�yK�e
G.M!֩L���IZ�6�,��j���7w�8߲���/�Db,�����C�Q��ٸy��l"�l= ������^��}l�� G��PA�����p��$���`-��I����Z!��V�q�1��g�U>f����R@�J�)��FJ��g�"���/"E�ҲK�2�X�|�2u��Dd�����sДu4�9^�d8��=�|�~^���U^�f��#�g�����w�Ǐ3wzQ��[��ə�c���V�Ư CX|�BS$J�vI \rH��f	ZTCi*�^�I���HCM���
���:��]�Mo�eZ2}�A1ga�H�.���-�h�6���q������^Z����a�����b�y�7�����'��p��W�ڥ��sohiWS)��]��m`�P%Iѧ�'��-�2s�2|o�^�����DS�jA|�W&L��hqUbu`���^~�u�z�����j9��H!�(���q�%�ַ�3�'^J�`�}�c�V�O�|�P�h{0��+���f��
E,9y
UЀv7�F-��6��׾[��Ay��Tع$��Mؾ��2�tQ�&Ye�/��~�G�H�Ic�a���iڧb�m�H�;m�yl�u$�g/d��"3M�E�-�F6�8��vN|܍·rl�/�ρ]d�����AX�`�CeL�Ŕ0)��d�2��><�Y�!���E�J�k2��ڇ!ϫ6���K�y�\�xt_��x�^=p��R��J���5��=F�~$NFY�Jv��#����H���C�0��	2Khڏl0Tv�a���h������C ���SA�e�C}���T/ۙ|6�L�6�����9aK�z)i���Q镕c��F��Vg��kH�fO�Xc�Vf���&�hաz	��$�.�:\JW�f�������������@E��s�|�d)�/oC��.e,�/
�{;^4>���X���xdɃR�q���+9`�}t�=����iP��v��D�*�}�I��B
	qͬo<'��ѲQ�$q���j|�[�����љ)eGԈZ�8Ym�m����3�[��CK�h�=������Ԑ�Q�AL9��Iٽ�R�� $sC�!G�;���23��!�]$rχ��ԟo逛D.�,υ.����\�]�1^cq��FN��:(i�2���?+6٫�27/o�C��n��o1%86	�4��h����7wX�t�H*�I틎� b9�W�}/Fަ�}E��f�F��脬��e8f��������m�rH u��ɡ��{��+��/�"͍>�]��	�[���_꾏~�f�����l6�Y-�QB��h|#Đ��=��L�it�T�ޠ/�[
�t-x�iD�9��2�Ђ�@��Aؓw��6�\� ��B=�K:T!��sm�Cgk"O�v��O�g�ZV>�,Â=��Q�Q���G۟�d޾'a7��Ԅ�6c��)fRѣ����,,Xw�GC����7!��u�k���9>�>Oh�?��]��d+Kt��,�s?v�3�]�tT��e��;�����%j~V	��.DG ��o�%����m�uV?{z�����a|=+p��V�M�e��{1���kz<�n�Ш~�wn�YV��O���(0��6"Q�ts�G�
GM�>��V"��"v���z6�Z��4}٭W56p}-�28l��o뿽�9� �)���+;ng�n�#�yd=���6-��]T��_ķ6#k����%�^�$d�>�9�WF~@1����K����fB�X�]S��iI
�K�DYjAd��n6B�e��0��fS|Gl�3�<�������E{aR�ߣE����>�S��l6r���j,tyPȟ����Uv�<� �h�!U��'��S9]zm
H�oR�?�\�w+��18=-�>���0��5�9�b���L��R�X=n���B�e�,)����XCF&lσ�g�ܸ�F���k�N?�
�0M���U��B�X~b)�jcȿ���Dʘ�a�G��N��l�頵׮���"�)��Ͼ�@.��H�x�����I��?�y�QLB��y_Q(�3s��f��s'���?+JG#}���C��˭����1-��{��o���UI|w�,G���U��~=���؃�x� {w�Eo��0U���,5����Y�t2*�XML�p��%�ٵ�����'w!�?>�]����m1���6�VD�v4�:�����*���L�?��2.́�ʇ(L�d�c���	z~^��H8!�5߅���}�0����E��0�=����V���"���v�wT���G�QJ�����g-K+?fK��P��g�8�E���~I`օh$��9S��@��Z�j���xՠ��ҏ�1�=��	�Uw%÷
��֯��s��	]�!�uP<櫑��U��W�Hw��C�V�q�HBʍ>�b>�%��%��+J<��w:(H���]�??W��e.�
�Ԑ��z��dr���Ѣ|ػ����hht�ay1������VOb��P�| @D����f��G�M.�U�WZ�'<YB{(ޥ�r$�@�ȭ�݃�Vw0��[����=���5_v	ѡ����D��/���TY��!�$�:A��t���ؔ�\��;�YA�_���� �{�5)���󎦦�^�$J#��UT�d�����~܆w0D�YғP��0/��>X��0I
R��64)-Ur�=qlC)�.���)�6��,��T�Г{��sk���~�����0 V'@�9h�[���TR�l�{��["�nO��Lu:wd&�֘
I���Ŧ*�K��`�R7Hq��̜����u=����e	�x�& B���@	��Ï�jP�X`>��ިN��u|H����P�3G�Ɣ��Fnj	���+��+A�D墨��r�疫�;��I{Ci
�E��;�T)�,5;�C"Oڥ�}%��jgIf.���.����+9��>e,�*�7c1��TJ�kmVL���4;RXB6�p���n�Z��܅F< ��E(ݝ�F��6퇥�χ�y�RI�=N.�7@������$$Yb!���5S�Z"��9n��z�"I�!�����i�ix#I���G��Cx���&(w�=��?�x����1�Ϋ�d��	 a���Nˉd���A#���{��aW8ŜՉ����ȪLe��C��RȺ�8�M?B��θ=�1@�ʥ���#�
X'�O�͐�
�Cf�ë��4��޴�:�C�`�	h��< zT!���>-�'�/E%�9��"6� us3f���ήB��k"�]�qa��d�Jl� ��}��}v��U�S}4��� ���!K��8��>Q�jt9P��{�����U���q�%R��*$�1<����zT�C?�i�ؓ��ڻ�iD�g�L�̍�[,z�ܧ>�f��������2���{��c+�>�]"����i�DW�l/�	O]��&��cs5z�:5�T�5yⲐb��܅ze!���I�$�cdqԱ�H�ּ5t9$�@�<t�7̘#�%Y��G���t������~���#e��K>�<�� �$���2�f\��5�HtV��i�u��5���TԴX�ªSH'&&gw���щv� 9&���7��T؋��P�ę2��F�7ҕ���T��)D�	`d)�I;�$->'�7��Z[�qI;\m��ը���`"�P�&P"�.��H��Op���}�Pj����W4׊`W([q���3�r����5�C|����f�� �*�>�,�LqX˗�S�� �S����r�MB����ً������#Z�`ۺy�8J�1~a6��	���IX�B��}� ;qW �J�0\ �l���N�y���F���U%{�2�-SԖ�
�X�������U��#
�M#Kq��A�z����טɝܸ� ���Mvc=&�U����0�ْ��JX㸳^�eR�O���R�,(��	|����@�[�.|?��G(я2(R��h*8- ��i�?�e;��׀	�;����s�.�a���m$V�L�������������M���q���N-��bQp��VI`ܑ�1X�+�{ei�&�Ѫ<
�u��#����太��+"��k��&�iS'�i�m����y8H��饼��1\��JKM��QȀ�����[�4�����hNr����j2��U�E҇�/��W��9fg�5~"�q�y��a`X�B��ݰ�}.�-m���b�}|��:����[s5s�ɠ�֞:d"?u�ה=O��ƈ�*�
�V��nA�N��&�mj:��<��>��YJp5fg\�������Z��!֤�N��0j;�A�s.����̠�ʎtM`r/
�J(�L0����[^!ܙv�����F	��c�G�@z��+���q���a]2���R��G���k�����M龼ª�+'���'�E�JoV�v��u:�`���޻�u{^!nɯ�!��\�y�����n�v�E\�����8Nv
E���e+�Dv@(;�^C'&{\ЭI�,[�2=�B��$X1�!K��}G/5�̀$&�.����L����EЎ�����_�(;;$^[�����.�Sz0�>)pa�5��l�U���Qݼ��$�e�b)��.t��K�aω�WIʠ�$��Kw�X<�W�EY,�뷃ھ�M�C�ѿ�`b����!%����˟�m�I�/�B���j��F^��C��K��m7Pw�`�M��R��[@}m�kI��[;�,���_����q\�c0t�0�k�A'�`;K���4d+Jf8e-r(n��m_<u~:u)F침������إB�@^�<WK�'��7'E��t�3�p���<-���|��������$lDض0��a�[�o��N�y�IH�U��ac�DͅH@ĭ�����0ae���z��rpX��A������
�I���>SSs��8)Z��RzQ�m~�@�d2D�K#v8,:��ܡF� �혴��o�G$N�14Z�ޅ�K�8�H��le�}ך�Lwc9�V¤V��N�UgW,���@�Q3���nj/<%��\��El�Pw��7VƋ�ҵq���BY�A|��*b�T������~���que�L���UU=z��~�6�)��0�U�.���U�+��R�����J��1k(���W��<"�yc�UNPҍ�1��.�\B�Z������4X�(&�T`(ӜD� ��'_� � �WAh�4ܩ�AG~�:�#�|����J�ݻ(*ixU�Q�����'�So������`-!�m���cK�>��^OO��{�H�G�iN6$����O�rő׭߂�q�6��M#��{�7}� GEK������A߃8��~��`!��ZE]� <�_ғ�o[a'K:�������/�^�Q�(Ëo#�z]>_�Te��J���c$8]oDN��R�ǋ�bo#�mA��a��#��ωp�+4�$����͏|�[mG�n�thI��%n�ne�$:���x  =zzQ��D�Ow9�T��3 ����u��q�Y�	;���^�ps�&���xg�^{X���S
o�]au%�`_J��f]�=�[m�Ċ�3b��,`�۟���w/�ԋ	��I�{���Q��a W�N|�B4��l�,����u��[*�W�U�>NS��pdD�}H���i�uLo�أ[d�m�Eq1����ڌ1K|��䈌e��x��Y�����?\7gz�B���Ÿ� 5+��<DT��?0�܁F*�͠} �~l�c�)J_3�e��%j�V�)%��2(~иث��+X ����X;�5;Q��y9���EIF`3������P	��M��-�H�J��P��H|{-s�#������ˤx�������[t��ۍx&�oF�t-	Ȧ�Dz��[#���A^]ą�ة�^u���>���:�D�lg��9�������{@]��}wB������K�P�3�7����A��f���ߜ��#)�t��2��*�)�p�v����J��R�����s�@^�r��1YI!�7K��RN^�;�.B�k/�'@�X%����-���F �����}�k6��c�)���'.X�0m�}��+���B�UvIٌ�b�+��L���j�悌����e
ҿ'�-`��h56�T�(�� >P�W;,A���w�]��Xi䓓Q��>�F�@WR6�7���Ǣ���m#�N����C��K��*�DsF��	EPG�ؒju�`��8��lIN�LH��B/_ǚTb�4�[�#���\��w��	[�=V��vӭ&���3������?ݲ������Τ�9�GE6�O��� ��H��3��/��e�X#i* �,6���Ԛ�k���^@B�?yV.�;�	���,(�/$Z�`j�F'�C��x�ɕ-�o��s�l^Y�Sl[5B���ʬ/��Z�l�Q�
h���G�.H�������KJ&z�8N�!������HF��_/�QnT�;��^%;�?�G�sd�gHB�!^�}ޛ���o �M�:n@$lᖛ���*�3���t�ѵk���(b��I�p�����і�`E�2=U���b����cם$�ZK��P�xW M���U�h���g�oj5���A�8���V���Q햓�8�gP.���Izs�9��įLƝ���K����}�/�6Y����ɾ���Ҭy�SS�c_c�"��z�_�,�8�=�>�m&�`��-��,�v���P7��7	US/�Ga���*�l�3i��V&�1��>�{�h-,��s�h��!�I��D�Au=�GLnX�@}�\-�#*����WR����P�q\���(ƍ�5�O��Ư��մ�5��� ��.+I��7��4�m��b����Zsx�j���l�IZ'��<x8o<{�I�M7�@�b��X�������<Azk^�\ ���y�P\�YOA?�v�lU[]<?��i.OKK1���Ѷ@	F�@�ҡ�w­>!
6H)HQ�`���bC@[�Ts]r�Hfò��K��"�n�6����z
$K;_�b�5��k�ySɢ�X�7#HG=ʦ��ɠ�F�� \�ح�2��������ۀGx�@��1�j�mU�#!��?(Ҷ�z�F-n�����|ގ�f\z�i2���T0�3��ʪo�A1�.�5��7�����D��݁_hDQP�Y���NiH��w�)���4�o��L�Ӕ�0���Ri 1�O�BɌ��>M�O�8q�>I�d��qY��6�j�_�B��L��u
ĕ�H�����U���QN�����MŶ��F>ɀ���K��O�*y�sZ�`���FE�T���(:~`�S�M�U��̈=�G.u�M���1��C�|�0�'&we&�%G�2��B�c΋XG@��b4��2L�*0��.$�	o`\a;�Gr������%��\�!;~�5s�r>�m�V�Cٵ��8=r�k�).�6�q��#͖��~GԢ��G�L�H�u���(�J1r�U2�+#�����mѨ�Ke&"�R櫭�aBvs���\h�3K�LٶsC,t�qQ���q�[���[ǒ��}�6��bm?�
��Nx�VCE��d\�����Um���ES�6�W�o_vB����i�"+��e
)�坱��J9�sD,CLN�7��q�|;��{
=b�����X<E;kC�'��T����H
�Ղ��[�Yn���w <v����W��* (�����Z���q���yYK^�'Ǩ�i�d j��Mt˽�7�h#g7�B������E2����*|�����B�xBI��mb[�i&/�]�
�,6�)@In&�ɼ�4"���1~�|±�O��9i8�q�W�)���QE^!�¾�3�[��w�6߿�L1���/�a)	h\�v��@���V��A�2i��޴�)~�����͑E]@��G���qX��t�.c�T��1�p���fԑ�1�E#���W͞j����bb���M~�m93��>H��pO���J�̀}��~���MSN� :M�A5�ni��Ür�Q$��Bxw���𭐄�>���;V}�M
��pY���3�(HU�{��S%6֌B�q��gY�ؘ�ϕ��b4�\��8>G*fym���	Q~T�,�!M�{M�ʷ�ɽ��1B���x7��H=�_��8���f�i�I���$�wSu��rQG`v`�-��f�p�g^�߳$51�xa�v[&R'�膐$��ʃ8��c�k�HK:��%A���w
�¢7��Ǯ%��+]/���|lD�Ro�Kz����!���4���()�YO�mD���,#�K��mg\�� :����B�I���;X���[�b7��?Ś�Ө��F� �"Z64R����I���>P�����zj^�T.��k��SbH�ׁV�$�Q#y�DhWF+�;䐑�Q`�H�f�Yd���b�z����������~��-������kW}�� ���o�cMP&���� �T�c�i_d����+�kL�ρ���3X��*���>땪�	�{�5��ZMMf��;�<N��gDk1��
P⢬��}���7!;I{_����y�ĢIv <Z-�T��^���j��H�����r볚�{8v[b�J'}�&Q���5����Z<����9 ݯ ~��A�, �]��؇�Ģa*m�E��TB��;��|���C��9�{ܬw&��T�?�"���%���,�[K�E�@�9�a�O�?�s@$v�q0�#�A�`	zw�L[��U��?������֊i/Qg�0��ϛ4�Ȉ2�bږR��R'J[��!59�7� � Z�%.񔆼75��FU�H�cޘ�[ݘ��_�Ω��z�������΋�b?�r�h�1P��P���:�r�{�#�-\���_� �mYĥ�s�3�c��ҿ�Ц僖�F٨��j'���,�������Ƃy��X��Iw�j97�������W�^��I�R��)2L�4Z�s�D��_���Vx��u�ќn�������"�oIq!����3�D˶]<\mn����F�]H/��Y�֥DP�c\���3�y��i�Z�,l�̢Ei���"��	��z�-����rl��p� �@`���w�i���OJ�h�'U�Io�,��J�1��e,�4�t>��> ��6�R�q�[M;�
�6�.�a��;o���I>�{]Զ�cyEO���n��K�TJ�9�����*��:�r�B�^=9���aF���y��Z��Lz��1�&�[��%�0�� �%��HSPK�]�����B�N���Vm%�t4tD�[P��iZ�d 
�}�S��C�)E6��h��ˊ�WLU�7`��
l���F�?��%I�6͚Ob��*F=���5�Z~)��X4%1u�+8�6�6;**����[֟�N���8gZ�W��8�m�>�|N7��� ч
)�L�$I`��{`��N"/�2Ȏ�m�E8�3�:��bx}�sq��#�l�p�l��%I���SQ�j�Xr&����s��`����cA��Ï2bj��LJ����Qֳ,��I������hm���-�.e����%�1D�m`Y��H��w��2�S��Ȓt�����@�a-�8()�Pab��
��ɨ/�b�7pk+��� ����-&t"u����f��㺄Ф�vn��7r��+K���Z|�4̦{J�6�@L�����rT=�����2b-@:?�,'��l�O�v:��N�"���I:�����\3U4��J�*g�B�j�nL��Ttꄟ�\	�t��^�/�}s���	/��<�4L� �!(4���-,u�~�4p�����(��������1��_��x�1�#1y���eDD��[��!�!��}�t?	燊��srU�|���K�N8G#�)	�y���[Hۚ%�Y�&�M��m���k
s1��W�Yr�����(\ �y����Q}�ab���A���n�{����F����?�?Li�HhZPc�aP'��Ї  謸�m�}�j�b2Lɇt;͵������Bdg�:�q/@��m��w����
wZc3*v�9%Q-碋~���`�J��Z�;ד>Y���}��D� �������w���DT�	�+�o���FQ�:�'!9 �k���g�� bC[�	D�����k|�M�
���֖�I��ї�$���W���*m�zT�H3]����O���}p3�+����a�a4ߐ���#â��z!�ILM�` �4uW�F�h���4!$	�AD3b/�1��1H?���OýN�`��Y�� J���۬���"Wz<������|��Zf�vRw��M��5�����*H-곹����:�T����t_��q/g_m��u=��rP�7��ۏ�B-\�m~�n�
Ȣhj{~0���
/��W�Ҩ�Y�XJ�����}��3ک�'t�޸.��[��"D��̻���M[��^��(����T3w��ٻ��}-��`c�CD2ՆDv7;$����̏���=n#���2�L�^�ɔ@!�(*�cg=u��Õ%���B�ݭ�����զ6�̼t���Ar}$�{	�i�{2X�bR����7ab�%V0�U'�-��gV���_�'$c3ڷA����MW&;����+T�����Y��aS���Є��%Gaߐ����1��q��gYt|���4�^v#�A fz��NPL��e(g�k��ڳ�gp�<�(�S��8�FzMe�,���ń���8Rd��H�����sO*�v����\�X~S�Nz�GK�$B��a�����ŋO�U�&B*w�+f�dƉ)����wB��Uw�yMQ�W�} �Y���}�n��h���]��@�H(Vd��������[������`|gѢT�<%��.��ډ�+�=�ρX�DI���Q`�Pdi���.�S��dx9�����(c��"���zB��v���D�.�I��{��O���C���|h7��=�N�YH>l/�����귵k^G.�
$�ڿIpjaD&�ԁjqZ�Ѯr��۾�rB1�}�|&q�J9�a�b��i�h��Ć�*�R~���z��,��D���Q�_\/�d����y��x�>FH-ks��5Fia`7	���	M�h��1Bp�zw�����ըɨ?��4¼ V\�~/�D n-��k�̇����,�K�"�-�ޚK1a00���Lb����.�lˉ����"b�&'7?�f3��8�Y�4�\�b�_~~%�$s2p�R����ȷ��*h^�o�"W��LWՂK�Q��MԋF�P��`m�S��U��}x�eƬ�ϩ@���L��xυ�E�X�x�t�S��M�y�[�G��_��Ę퀅�_�˲��_�����Sd0'%��v��#�E�XI�����F¶�]��#4�@�9�09niy4�d�������7Dϱ|��I��!�mU^�kl��$���j^�A6���r:P�;�H0U���0Ol�ۜK}J��}ڀ�'$x���@e�RqPݰ3I�(�	���uwpS@1h����:�d�U�K;i����������\_�+��٫��N�m�n��'U�!�ū'z�7�"�x� �%���"!gjO*��
���ӕ-�������ܑ�Q��Oɾm�R���� մ1�� ⓳w!�Z�N_���A�6d�����56-<�ןj~��o~*T!�9;�O��gX���������<�RA��S��0�mO�X�Po)"�����K
��n\��P��E���>;��%���.�m��Q���q��,3zӡE�/ʷ4�	�gS3zF'�5e�>2��`1��眢:G��n������QL'�:e���%(@�$��J��lE�ħ���[)D�2��-�rP��&:UM	_��o��΀�E1����������#*3�x�2��9����"�*�@DӾ��ls����dq�5�qG��/9��v?^��~��o#���M��
k�飠�e*���þ;
��&U)���%��"!Z��:�	��z񴯒�)��w'H�g2�u$�-u����12X�BVŽ�� �<��,�wm)ODt����x����G�o[Keқ?�v>`']"�5��n�k5�Hl`�ӆ\mV8N9�����Vh�\+�g{O}����C}a�.�����z.e��ṕ�)p?'��+6�S��}]�Gy��$Ub�����"��e�v���� � VR���)��n�ƈ���u�2��'�9a�Ꙓ�j>�(@��T��V
EXp O�	Nۘ��*Y^���A�a�"��*��sJ�]Ыa������}�u8��,A�������B�?���I�L�>����M���`ظ��i�4(O���DSF�(s�邮��j~���Ä/���ܙ+���$�#��se��2`��a�t�>(H3<2�ޅEJ����{�������~�����~7wg^�gu;0�HPzQf_5� �����3��S��h�g��x@��xxj�	��;-���y���r{K �N<����E���Glw�-#cj��rr ���Hs� =��\M8�nN�x�C�$76 �\[% DO�\e�;q���(� 雈��j��5XNyLK��U������تG0Nd�c��\��B&��Ǯ���j��z1a��䉨��L�)�������1c1���̔����BC�K�6kf��!B�Uq/�>,,(����O���Z���\�'�_�9=<�ۜi8�Hsf`wB�`�F�ȗ�β1˟E�S�u��sI��?�+@4H�����A��3ƙ$�0$�*���Or�g�0�uh�ڄO��@��El0��`��S��g�tPO%��[��!�����%�*HG7���ʞ�mN!���o�#H�7�%c����6�cwʲ�4v��kY�n5����V�#��d��x<�����LjB7���X�7��z���Kz�]ele��Ǣtj-���5�=p�]��O���j1�iu��F*ᤅ�#�	�i.�Z���XהbC�:�RK/Z��c�f������d��E�ѓ]xT��c�=~<�,�?l�G��k�W�7sS���ȧrY��8�J6k؉�u~kq�p�]Y��^��gnbw���D��Oh�\����(�5�PMy;P���ZG}��X�#���q,�?؆ω�����/S�)U�H���L�\5�C�gP*/��	��}1�y�a�����3#%��!���t�N5hs\�������0 Bd��#�!=����:'��z$��
	Kw�}���+�I0N��6�ʣ�8"����
��f��뵔�94T�=F��հ7&�}�K�q�h��F��2��Ji�����E�U~T|�k34�T9�*aG[�&�����e�՜�ےx8یݬ/!��Wى�G�vO�w�\&Ͱs��pva5aд`�b@m�-[0K$��� ]=1ެQ�1�5���$�"���S�VS��פ�)��H�S����(@Gm��'j��.���W_��#���1P�f�E�4�pFܕ"s���˝Փ�38�K�%�n��-%H��x�"�P}���m��D�L��|>���6����{�]������a!�H~S�博W�bĳ�L{� �����yD�"���ô�a�Q/��0]^�V��9@�Vl ��>��y�FR�I-甛k�����K<�����/��a���Rb`vm	v�]h�e�
9y�|i��6E�@� ؛�����v2Σȯ7����d�L�����*���0�����k6�S�BNr�%|_@RP��~��ט�̿��4d�5ϐ���KȢѶٜ� ���Ӕ�({��/.�"�l#9�M_^yI��q��{�q	yl�
\S�?��Ͱ>�k&�Gw�~�8T������q{�De;G~d�"y*- �TSW��Bc~�F���juPQl%_~1ɛ���@߲r����@���:'�r��o��Yh07�!�Q�����v	�	G�u�=�m��G�G36�]
<�7�p��0�U�p?;�\0Ld�5r��X(x����[��mTC�C��HCk��1?Pm�.���r�"�����$����n�c,�.����
�O$�]J�͕.E�L�ER{������ѦL3JA����I�kM�ME���@刐�_��h3n�����j �#��qr/bĊ���:)3�%K�m�iB�$Yv_�­���4�g�$��|U�cp ��7Θu*?Ȓ�*�]?*e���c`U�/:13Ea��*ENV ����
���j�P;�V]�-�I�6^$4M����T~,gdS&���Il��T��ɢ6L��۸��ߗ�I��
�J�2�̕a��U����_Ǯ��Wէ3�\�Pܝ�V
��ERȷ�a��8�ZQ�]���;L�H�_����aZ:�sX�.k�I�NF?�w��=h���W�wV9G!����@!*���S(5����ɿL���j#��'������+]"���G�C�b��ԪD-��@v-�v�V[��(F�e�,N ��OF���������S�p��.}�M���������A��o�T�X���_�"���C�<q�j�vf j�TM�sn����R���i��s�d��򤮸�v�KX�8��!�J�g�t��:���W��D�=�Ԁ�XbhA�T�p��q�Ѷ���{!t+�e�FI���GT������e�5OC�q&$}�N'� Cw��S��:h�����e��v�ƽ�ڳ������G�����s�h"k|���*��+����M���[;w'e�<J�؝�M�0$K��4��M	DU�,�&�5�4�B�łj�Ǻ��[��s��C^UaC�����ŇA�v�0t}�~���s�C��=>"�,J���~�Ei�ã���,z�0 ��η=�Y28�m3��4���S/NQHd�p!����a��UlXI���efa��r�ћ���u@�hol�Y���E���)���A��D- cDZjY��w���jS�H�Es)��A��1z�(�ɓݝG������'���U �dg5��9�%C�-�G
}�c$\+��r�z�䜖��|�M�&�Ak�ԐNeiёM�����{'Q?,5��h��ÍVfnm�\`�"b/����P��P�i�����D��p$f�)�v�h�W�%mQ�9r�첌cy-�ʳhQQoK5�Z��!��[���l�w�	�gl��+�ٓ~��?�	���S��a�XggtJ�<к!���q�=k�V���l᣹�����.�P;5�a�(�L[��s������'�7~Ik�������W�ξ����d�j��-��bp cw$Y�վ��c=p�Eq��\�0R�^�`�(ٞ�"�M�yI�����b)�kjL x}_/����~ͱ����������:��4� f
oH�{T���LSTO�R,��g��^uP�T������{�^/V�����i�2��K�g���A�ߣ�o�@�G8G�ǂCɥ�^�����dv�+4�(�K�O�sq�< (�}�1$���VB��e&�*�xA���K����^�1�P�v���s�el�^��r!�Ax��~�p�Mрn.F!�^�������-n�^���k������i�����_��x�eQD�F�:�5nf:�t6�ʫeRo�J#!�eC�y:�@��a���|.���0�ހ��F�v�I��*L�Xl:����uކԃC��;��IRد��.��斋�⬊s�u���]�'���9�:�­�t�舂�jx�R��+|�ب�r)��,��F��W	g��u*�H�Yͨ%�� p�C`B�e�o=AH���
�#(�������T�S�u����`;6�ܻv��� �^~�,��׮��������V۪L �W��I���Mˌ+���i�]�դ�yZ�NaO���h+J��a*�l�4��89}�k��&�gu2z �-�'�%#$��٥E�8%W�_�q��Jz���n�h-X5V�|c��6��|9���fS< G�B�0�Z[����5�R̮[>��;wY�S7��*X�b�����8�o�����SΎ�!�>�����cR2z�D���BN)���������+/��%��:�iB�r`�h
ze *.�@[�
��e���4F��pr~��D��꨹m�Q;���P�5J@V�Ȧ�d�����f�V֒��������y�ۢ��«��ɜ�)L�,`0�(�^�쒿{�w������_?B��뿤�6)51���MS���E�!��L)N����O_����*+f3�"3�a����Y.��G_l�1WAn� ��o��P4H�w�}�v�Po�����Gsʢ[�|��R�vo�K`j��[`}�Է%H9�w���=�
/�ݾ;���L}ל�ɸy���0ap��p����Z��V8�.1��8�Sq��mw�U;��7��{�r��f��4���C߄���gL>�4?S,U,4����r�v��IS���2��.�q3�����Ԇ�ɻ�6��p|Ut���CA�DC7����)��f2����2�*$���N��Gh��e�ס#4�ge�0�#|����,�(�4+�Y�F�Ԭڀ��S�;�ٱ�A�oG�T�����W�o{F�R)x{K��*[��Z��3�ju��{w*���a������򝐈���g'['�\�����Xz���CP���x���!-Z1�)!�����ۏ��CSr�FE�p��:��-oO�G�l�q�߉Lwt\O~]�l�CZ`(�����7<R?�}��29{؆K�4$Y���Q+x]Q���6q�,n�LkԲ�#���B��g��(�9�R~�hdq���@�� ���u{�{cq*F��W�o�K��w��O.��z���J�]6X�	ߏ��
�:d��� z��uc�rā���I�׹G�8|��#&L_Ġ��v��X�!jA\��9����v����$��xK)<`��N��s��&��z�^���o�B�{5x0Dl�����ewW�i��@!���饬X���x���(3r���XO7�_6:�j\U���[+1�+�t��G2��E���	c/��؟��^��'uV���gX�ޞ_f���,�Ǣ(�M�k�7���~�2��JF!#W���Ց.�rn�>�`�n�,���
���dq��PpS�t�}�s�8��Z�?�#bo��t�d�r���q���Xr=sI��ZiQof��^�rP8�&�fho��./#������H���IL$2�}�1l��iC���{����̋)���\���O<�!���9H,*�h�MA>��	����9du<��y�t���]U�KD3 VC��:�W�
���T��r;a�es��bY�k��K��^�T{�v&�a�����=8Tf������F*g���1�o8_E��nkh.���ǉ��e���i�@٠���`i<���~��=���c��G�d��U���S��M̕�5v�g�.��[,�J�V����v|Ȋ+���J1�^
|�D���Nө�ъ�+C9^�b�sV ���YM}��@��f"RVji�e���kf'DP�d�w�q�=����U`@��L��b�G����o���I��ID�^�^f�h·ئ�kx��;�)3����l\D�;�^�N&���N��x+7�B&��+���JE��U��Ԛ��S��oMj/hl�eGv��+�H������1>��2��ciy�{����u��)�`��	&��T-��]ڸ���ѡ&����
�1��U�8��RYt�(��`Cn��A���e����B�t©�qyx��j����F���uz�ܓ�Az(�R��z%#���p�K�^�H�EjAٽ�8wy�������<��/������恻��7�7h����-��V�|i�k:�����!��y���S�o~5h��`# _m�6رbƎ�{W�"�5�m��i��?B�0�H%�p}�.i�(�ؤ��C��v�P��]z�.��oy]��~=w�y���>4���� X�u:��k��<�p���j�F�N>��������oM�����S+��A@4h���;આ����dT�*bO�v	vٮ=�W�Td���ㅶ1����Z&W�|��lEMs��n�d����au4�R.���>u7G����9-�N�ph��5�8���[���5�1��ʙ�a�)v�<��U�L,����@:Q#�{.BH����χ��I���}gE6��8oh���y����%��d1B����;�
*�tĻk�Ěu�ed�To��my��Y3���Am%�[:����C�n������.��<7��b����-���N6�V ����8�4�w߮nA!�~�ή#뫳�U�u_Y����r�
����1lc��Kèj' ��5�2��OTMs��p��\�?ꏤ`
�2O_�l��4B�F�7��
��YyC����+������OsR�^ώhlq�`���*~���~�Q�ì���B� �O$7��7Z8_����'C�~�\�}R�xC{�@e��z�mt���3�������bu�6EO}��i�d�7X*�������j?�U������kt��P��ء#C�\Kg)���dSF��&^��^}�~��]y$�g�P��R�b����I����\�<�f�}k-ܿ`�Ϩ���F��m<��C\u��?Y�1�� �g������	���w����=�)��&������6kL�jX8��FN�)Xk�-W@/���PV�A�|�]h��u���ƌ$ $�JG���)�_�����ƴh~��r���O��%�J��Ys1���Z����� A���O������Ŵ��z�����u�18��D�l�"��!�"^��� �s�x*^�idC����,՝8Ř,*5ŏja�����;,kٓ2����y+�����{9�� NN���_}��Y��x,�@���E`���r��3�x�zBq3k��
_��� e"�Ź/:��M=!�*�C[�J�">g���.�M�z@�pw݈l�n@T0���k�%�a^@M��(���Dv��^E��E�ۚu��oO�a�C7O�OL�K�]��܈���}�������F]�=�<�����hp}� A4��j�I� ��P�R���涢���q���)�x��˳�$6����G�kG�%�4�� �)�fp �]�+��W�� K���A�iT����{���u�V�[�F:�h�x�K�Zm�_��m� �/T�e�+m��X%���Yx���=L��{L��Ln�����7�<�o��hC!�\oy��~E.7ȆB��{/;(??L���(���C����97��)�޽ʋ��fTq�����$�R�s��\�� O�57ec�����z�n8�����.�N��^m(�>�x�([���W�LH�o��]*�MW�r��?������'q�1�a��K��n�/Z!b[���5�q3���&���u�NZrm�<V��y�!�3
ZN�� ��h�[�G �߻n_�y.�&����E�?�k���C�2.j���2���#w):��_�9=��B�O�Hu��Ղ%A )�����pKN.9��]��Y?:��A��6sɊ��4���ăH���T�2x��D�^�B�s;� ���S/PփNb%1�g�ϴ������7{4��/�}��:�
D���0�+6��g���(��8B���=VǂS�`�'�2�̫.��@S�����N�u#��ӷ�*��*����6�a��Μ�a"YC��ּ\����ϼ�T�.)�O��m�v�Tl��ZU��!Ol��I�����T0?��:�EZ��Wm�ӯ��Bh��Y�*�Yx��2�l\K�Q@�Ct�[�C�_����;�e��"p��0@Z��7�/�k���S_��>J3G�˰�n1�h1(�d��$N����*^������n؇Y�k��h�(Y0"�����_. ~���j3�Ge[qc���
��\Mq���)W�/�6�m[�*%/�!���#�eN+.\jD�b�k�9ָ�7k*ou-��V2{8�
�$��Qp��1��i-�bO��g��Ur��dU�T%� V���##.�Z��`��YRuހM�Nf�xچs�`�P��]P��Ay�[#j˗�5�-�n���:���������*x��	nN���M(=]�q{[�Y�a����"���UVF�]���]�����C22k�)�`�����݁N:�u�� qο����@DYϥT�?"��Ȓ�d1�k��8��ਔ}�1��L��V�S8�"��1���%:����l�<3�&P��vr��3iU_��9�<��3�a$T�*��D~��՞V\��)�ޮr�#�]؞�����q�]�,���]Sڙ���̈8������aA[*ПG�"��0��>�E�U#�U��o�Y�zu����E�1��z�T���x���h����R��ixC��
��O�V�\,���������: ƅik݉��H����	���s��6�E�xڮ|� qrŵ�af�.�=�u{f�#G��P��^�^��$3��1��-��d��6�@-ѹ��8�X��Z��#�� X>|(m�m%I��i���?��{zk��H��P�IPޕ��M"���eϧƏ�3�Y���Si�8Ϡ�a���9K���ge1n��<�l�o(��DQ /5��#�6 TR�c��&���LKʑa������g��P�-C.څR�4��4�_���'j��׳���b��y�ʷ²���`c��k_�7}��l��¡M"��?4����R�<O/!�Zl��YC��"�~}�*nMW�u����'�|K/�D�]����h�w���/�!�df�����.M���_�WM�Ȧn��\+O��@��u%q��+]����r�a[Dup�le��-�n��@���GeM��e�y�0���