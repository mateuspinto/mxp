`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12192)
`protect data_block
0H/MXe6IVr16+b3n4HufYH4A9BjdBzreLpZPoKtQBfEmcOVyQRjqJzfL2us0d/9QPBT0HifD3nxI
IadB6ycOoIveLkCRe7hV8OKHUU2KMQgdKd59/tZf1v8zzJSLekhD9p47BXM7ZpQ4ZKRVRWcjXfG0
TmfXfngQ8EjmuSzcfRWr0NYSNCwnnGSkBY5zhjuwJeMRft+gs456fhwsRXz1DY+b9v71zsEZzXLD
k85fCOugA+LRLI1QJ//Z3wK0uHKu0vWV17pBreKlrKMgw55G9l6uPu2FiklMmx/k084O2UyDi1XQ
heVkw6gPNcwVZtFP2TBm2ScENR19c7du/lg/c4lHpYB5Mp2K8mR5EgF4tsoaV8Ou+r0INiG45iHu
XbgCoobJH7hrZ3xGcK4RPkP8CaJbcwu1u/DOabvJ92qDjyl1qi1Wa1hISIPuvwMDqgxNTcxDFeHS
4WSxDGbTuQtTNYbUiAcqMhEdXGXvtMYzXJuSCl6bxMzFmc4vuSCpcIG94quJUt8LCR5opSuJQGPV
67IMIvi2REXUsS1I20JJro0013Sr6DaP3H2ULitaqM5TLcTB2dojhdbUUMcky9pypKyepqhiglD+
vw4dqsv3nphoOAakoT2mun3vneLTQDcaqRi0TQK9cL7gTUhBeV313O8+0+2ned6WpexzglNuyDw2
w0pQRu3Z/J3UbSZb8c88ZkYQdkd9u17Sah7NY4/tf4goXp8IufeInzIaNU9X5hbAq5+HS8soXKfu
CwHL8ujViiLzFIAWDaCy16DGVGjAnJ2H3R7NcEUZtm4VOf6sonky62ch6AXQmy1RmfhTv5LLT/V0
+myKAKADv7+GV5LQp4MYjs+SC567husRbTHQ9VGQNvRcVY3jXmyHWFdfhJamm/DoS+Wb/UsV3EKU
bJATsAAZ+w/meFOYH6idBsICglyqjfZYUcfK64QB1k79NdAdgMF4t8FRS91cJ4PkFZxmSaDPGYVB
MzKEcM08JvZd2VyCjSFLU3WFeSHPI0gd35U/xEfElpEou7gUmqp+rxTcpK3sIAi0BNkJwSqHEjjJ
IAhMlJcPJvVOM1bG+fKuHGtjp9+rbhAp/T4YR9WtjBXrbQVjhnOCODTFuYfuebm+nqkS4eOTIA/8
29O0h//jfnRCMvj6uCDCSpzjB2r27i5950G+BKGvDL5JR5MXEtUeHxQhtThGmEfxlCqG5QCusMTW
anDw0Pt49bU+ACrRQmYGoGZRCbPQdL82IevccsfE7kkfqHxZiy8dEsMayxt7/n73tc2iqjTpuGCT
FpAdR7r4L8J0TnObSsE5Z0hxrBryGgZNJshgKaF07dMfnTygD4GqWqQJ6eog/fR1Dv+iFu5jujZF
IYITrp/oqbb3uuDl8xxGWa7VNPveyxHbYiHkn2XUZPoEaC3JJcbhIlc47Czkp42NmQm0cp782C6U
HI3XTCdvn2l1zEyxvD+M16eQGeEcvcYACvUGcxJbiaJ/kJ4iYDhNvWVo6G6Xi/qnALvEB5v9bblP
5eZwTKdljGdCI7cjwxAyXVM3QsKItYjHrpocrC6bS2ogrdFVAl420lYZXrnvjP2LQxUO2RA6fl3v
nZcAorNQIhNaPzA4E/P5GEUDqzw88ZPIajh5afzP7LIHHXaVrUdihPBGxsXXE40LcfHyJI9Pe43r
WL+ZJhlqP/5IOpACWuXHLHm2HcRxv8ACQKT546nyMGVtoVPJePXt5vXu10B/+axBSUkxyobhBowt
+ROC74le3nKTzbVpuQuPGRq/3BGE5oyva2MGBvloV6WDTdGQfNl48m8Fm5zseaaAvqd3S1QSvQdg
ECyiElo0heLttIH39NSzVfbUc/Ym8ariouKRm5d1sNEl0GRdJJfpTV+J5VeOMg0R0CXG2yjHv4E1
mbicSWhKy3DUjA0PDvN3cye7J4ujUt3B6pO5KkPeZFRJFnWvWzhPziWcFZVeY3wKUvJdQ6uwb5o6
nFIDm9mE1yK8xNYiPk4jTROmAdl2mlvJFdqC57TLZWYReIiQIrQLRDnUdjBuSUuZRPkZ8fi7lBKE
hN7r7BPJHTbCfetyV0RB1XgkmXspacBX99yAJ4QQ0CL5DMW0tAygw4p/edln1Wd7hkKxa53albLD
k/PTD8j6BbTCLI7lB+VA9oyrLVMwDACJGP1o9vsbFe6sGdI+wmO0KIEKlU6gdNSqoGc/uDyjt4ZI
shqv9zgIa3xI0N2kvGijtnr8jZpf5a3t13z6YT606r9X8kvAuMDygS8m8rh6qVKEaavSNAo4MP9A
oTGTutZjFmKJbsWdnONAoFMFAMKKBYmoUx/jRdX1eIEEPIbdy8SwcQd7z7xeJvOMqWvlatGVmUIa
2VvcTfcZc6u4MEtG6iI8mo+iHsppGJ1I5HRrdJ240UL1ZlRzkEbEFebWkoffINtFZpogJHukaOam
u/iR8oRdBDHpCZhQOG6hbJZfvIeUuZjNctg3AsxCClGFSsaOgAeNMCxxYPfSmzEv87aVjCZjV8k6
KrMkMlAk6rsMCDmCXQjAsd0A3OGDLRVQ9yhAwV0QikkZjw9aO5kutFZ8Af3tTpN0iRL/gZqJTaEF
E+FXHqFjR3NIIqVefaMmtJXmGIUWWDyplFu9i2s1VshPD3vA774D8d2+qiZBwIVEgtWVfnsWRXJo
Lf+KIAL+eYvAB8XUnBZfLCCeO4azioHYywZhHoKA7f0h7qU9Jjhtvpi77kLHhACjgol1/t+GpaeY
7p2XwVPjjlPw22dIOwALysA4XM1uFyFn5M+A9orrCaw7cHbXgPksCPurBzgRXdTehIeVjR+K1wNc
U6TSvwuMj6n7Lw7sWbB8CKwwPYqceh73QgRqDI/7OeFKGnAza6NY2K5LG+jta/rXp2mh5kZFWAWj
IAa6d67agdU0Kv9jS1GJBmGGK0XEPTG+eu5z+2aOWxQPqK9A7GbYCv468W4Ni+qBm/owYGoU2dmY
xyGOBQ8DtaJj/3Lni8/wjUCDQ9jcNcdM0truuXv/rcrq379f45NVyvirAPEXpXRXoAodYH18SObA
qkrnByoDFmbBeUdLLKD4T8Kajrb8GBbEE8ryDCxRnPeF6ewHXjCrLChkyAFXAlFUGs46LIm5BQgG
x/4CgWwSWJtf98Vnz8sT1GE5HCh3oTTlq9CVoJeg9IZtidWX2I/uDsUDZW3sAXxAjZCm3oF3XAnJ
aUoUV/IOVKOgtR5+JUJ+HeUrbKv3gmjG80s63urx8Od7sYqqONZtd1d10f4ei9/b0Tn3Gqoih0kM
flVD2OsYSulsMiziDRlkgIdUqXO7xDwlMtHA79xlqzgFhVD9NXTgfx0jHPPfu8Hmhr+tV6gdrNEx
corvJ9t5Qu697x2IIiJ03h+bhY5Xf9PKQrv6DD1A5bT/5wTWuZl9FhaxjvUzTG1Eru1kosrf39WT
otzCF67k2i/LrnTT5lb5lIkys8UjHimSNTw/CT4MOmxSZL58UUSTftdhHTP3IdZNu5QE5F11cbp8
Brb+unjgl9qDxtth4rdsz5Lrv99lRAn96lw7mIQ1zxWV40RUpDvM1A0gHw0hYbCMUNEraIbGvzbC
Hct4qO3BUOm7vHJ4jjmuRcfAeX6XSJGbwthSPwXIVIIOGAGIrP/BzfR3H6xpoUvX+u1mCWf1Nl8u
jjH2cXePMUsUEJFhx2bmhqiKX3/ug+NBD99jCzhZltYlwgvlFvUexA3NdMidwEm0n4RpWi90vJz7
vQnAEDBrUwhA0vvp4UiIj0swGr7N4oN5hzpX+hUuM8lySEZ4duejlq2e02HScLBloiqtYNUVAwrg
DGEF4Q4Dsk7dTHm2HPAzFyRDBAZdPLTng4Fg7zlza/agAOa0b/SgDm0WrSY9T0JoLPHojDQNw2ZG
5Q6JLKW8DZuSYj1f3HXb4zCEVABDPHNuz7+PhWv4bkxSi3V68RyBKq4RqQ2fL0ROHDIQX6k4rQde
kMoVwTlv/j61UywzBKA581OTsnpxiwjd+6HmTHh4B5432LKdvFXaskyYMytNcQiM3fZpJ+Qv4pU+
qaiWiKOj9/o4C34gPWXDXw0/4NsFO9WmElvU0DuA79PZOJZ5JAEgLxVUp9RFBQeICbY7Nx35kxVc
s+RrLceCHQTLVYsAYyIqHrpLsQk4wpwmlx+i6C3GsYBFvbEEuuzb1DWj3bNsbT/QPAXhKMiJ29F+
R3G5IqwnPaH5Xo+g6PHUAnYGjCWEMjSKS0BI6SVp1Dzo7M2e7ojNS0TZ78GFjhqjLpd5yUqsnEOc
UzNE4eeS9/CC9bxb0REzcVdBBalCf1j4bJtIEStk4LvZkTdDZzWJQwEAf6PAFnPbnk2jNOrVlTtR
wpiHXaQ/jjn8Ulo5fi5fTTBsgC2NdGgCaFcA6kXZ6Ln+FEbG+nvko7TMn7f/GzQT+dGsaG5wAcx/
1swKKyVw3RTrXLVihfsWOlJVwXpJEE4URxybuGDm7ajw4RMtbxYMmvdPffppKcLvfcZXdOCFeC0I
SuCzqRPZU35u0LXg/AlmFmrNEd1x8WKWN+a66kmzQ2yH5YCSwf5L1nMhINX2r25tQA9/zmNstmL1
pMJiC08TY1HhJxu81NuyJAX7AYhfLFWgBF0A0y3n/JtU6vZ1tyKvvOvYa7HCeNoDerhtvEgmA7Tn
k6Q7zf5/KidWSS14nmpEx0LjFlZKCCosknojZSHjSMQ0kmDCkcG44lEkudEWFw5r3b3aJ0vJY5uC
1yq3hMn8cWUOiDCfKSR+zItCqSkHzqNkL6bD2jWqLPk68qB+Wh9BcamyWrSe/jFp6tgoEV4/dsoL
yY1afJZWW2f11ynaIyV757b9tWZEyN2yW8XckWI21JZDZ8u8KjKvO2LUsUw9raXSp6eZ5pFbW82D
k0K8pDdjYT5104XHTix6739+GwfGs5hXF1K5HUz5s6+6MNoGxiNk/RKYyMwgSL5069C1QG0uLQSQ
UXTi1TJQTTwHAEaiVajmNC2pQ5+a5obvVGBepPJQAEpyyJLFgZWOa1IHo842lfd5GPsprv/fX1X5
2A4OjrBeJogc2MoHg/iYR5vwcFCtYfxsA7OXqYXGCVIn0I5sDnGTB8p29J83JKQSQrT36FVRlNzh
m5B0Sq6KIHW7eMCMXdbJAgbBoFVBMYhK/WEwINJOfxnkh+QnX58kOpL83uMP2B6xWl7ZmwDM8WmL
v6864HXrteCM/ojDzM9NA1pJF48YgV8FFC8IVHW8O1CVwXWRLshHJaF60aL0QUEOFugfiS5U1jWQ
esmdIpoe4XrDqOXSfv+zLJ0zOsg+TtZ7+QuZgAiX28khpR4kShztB4Pc+S3lbkBTzV3xX6cPlU+h
LO1ppuoa5TkOPop2SAbS0PXuK1y68SNbEZz48Qyl7gHB+O5hKxlG/IrIgQRQBHpNV4hHtXovf62C
xuTOsIfq1/xk/BW5xKryvhJVKh4OXeEDPKF0ZJEJpjfXLmOX3RyWYTekAcgqZ73UoqnLllAHlIbt
qHrpxBFdy72Ke0qRNNBIysn9hOZsbA9AStF5VxpvJYBVywK3RVk4Aqv9WP0yNx0AAWkImZvuPkWl
bxYVfUIuZi4T/WmqYx1/0bfgWZkBwBAjfnoZwCM2L0Z/HHzktjqF/IffkELNNOD/doryxCxVuBh/
AKTucC9/TmYSTkQSaNCapWUkBPGM3ZPmQob5CK5nzpYWfPWF9Mwowphi5HrjA/pOzDhmnufVoeOQ
JmQsy3SRm+HLpzJEzTiQ0jwQDknmQq9BdvMGGvNLBph8SZOdrPwFkWVgdk4z5oJLJggTFyOTspvf
ylyBF0/ggvXRDOMDBu95e+FPrZXkN0URHpeLbbCHoIWbQt/m6no6Uclgnm6ARZLniX32VqXs3i8p
fxE28F7O46Ni7WKwFwGgfx6ASNY2AihrZG1RlcL23CLUByHVoFLDPvFcGukJigCP90Rnb+lNEwGK
JUPADfZiWGGEf3cWFcaFBPRYj+tH36CmyCbFOtaq3aF9hSrPX6OZ17AH6DfbrLVp8e/SAVAUZqa+
nxf+4u/+a5EYqDe/cy1vukItGJ36kRvLrcTLZEnpKcpFmG+pzdP3WBfr6ORXndSJ6p2uDRlgltYG
D87dDB6sj8l6W/keULZbecPmMvpXxzObxAEXPAPK4dQx66Ev5xdgGZtPvBoUf9ZZ2MrkopNKCNd7
Fzl2xDzL50BmQtpZUu/zjsRiKgEK1j6VgqrMfns35ysf5NVBD5SIWIFkNoElaO7ak5SG2M5RobfC
4pm/cHJiRU7r8D19M/KcRACdE+B3I1k4t5IlX5rkVSNRQm85TMp6rv3Xr7VmLmEgurinWZeOk5Lw
mWnzMieFLUt/SOKETNRKq6rNrDpPkNSrSvnxL5t5z0O40UBCJ0za2P+F4R0VUd+5WG8FWZvOE/pQ
JG8Qjx5y3kC5b3eIGqCCkyon7LcSVzHMM6UTB+pj7+p7vaTi6cBPgJTopLhX5rllJP/hMOg5r0qZ
NlMLnlLMh1VukUkanjdreZNWrn3bIjXXARCU7f+MV25+wKlWto999Of4goUC+7RJnf+2dSYXRiUK
GXActG4EBeCSUmQA+fmamrTNKWVblTazueQjprHspD5YtCdlwykztmSX24ZK4Vtq40pBetwl5Xl2
sJ8iI4fTj3f7I328EqL9j+YyDCmfSV0RrEZJuXYN2hQFzoUIQRCPTgIghef+ehLWOrimYjNd9icX
YLCXD5Z+f7K4qcxGbt+wk15jxnp4+Ks6Lir7h4lRUaEhGm7xxpXvS7IRVO+ZnldnQ2B7RBcyykPF
gOP7TKOGCqloND3CoKDWmyqbRKW2lPG6vyCMUa1px2PV+i+nAHFgb0ca7C2WlapmVMViyRWIS4rl
CwPf/90+jnzJa9yCwnA98o9aQ9UGytA/6WB/uL4KFR0Fq9vF/PAzuy+CoemO+RKiU+sS1u5HxIDN
pwt9YEyLaOsOAgQyESZ7p6Qyc55Bp6uXzMt+jlqKagDVWKoF/2gE8bvpH3X6QYys/8SLLuGEG20L
vYTXknSHB97DBKX1DqfdYC2Jwvugaps0echuXR/UsBzHnDkIPvseXN8ww5OFkZexn1trSTKvUGFX
pZ3CzVsddEFrCcjdxV9QOeZpc6qxY+xxqTdv3G8BfCpmyIKNTUanzyTtvf6/3JtzL+PAWOBhIShf
ZwRBIlYmz5kqXB+7hqd+egEUvM8fS3Lb6J0JaJ95Zw9qNWUqyDuSHGCGj0DsNGWFsMyyqkWIrVun
w8/id98GFcQ5MELPJAkm2uobcWV0hB+tZUG965ZhPH12KMfQBmm8AB5EcE12RkT7f8/GSjfCtYRx
wN/Hfx0XcIXtZrjjSb8t1ezc2KZfvJ8zUWy7fokAIljn8MSj9KAAoXXVua//G+if5DIQt7s3Cqur
fHGlDFLLLKqyMY5wH5PcTiWHWRHiFvkHnxs13BVHhNsgYlRkbEkY9+cnUkV4UYyIxlZ9xqrgx5vZ
9ldSjzbVbPY2iR98h+YhSfx7zLA+RIymxU/gO/3Q1147BhQPbF5e5ys6z+OqvOG4J3wnDACC4UXF
D+xvlbCj6sbptUpRnC2c1Fz1ehIrQim9D5e53/0Tugw48lLlGe6YqyJ5NOf4NntsD+dNLOZrDSRe
fl3FO6CVFeB5/p2WhZFxDHtdimNInkFQgiG5cWRvmkBOsUGMYVw0G/zGQtbIEY9dsAlvDrW4ssJK
0al+oRw5TgeJ6L/jHTObivsbRyqNvil9Snwbo4pDMG6m79C6aG67rA3l/Vi+bJ0MW7RsFORVOMvg
s8lkNpTYxf1L220o6MePSzjCVTnMRgOVOsD3lsad8POThHAUyvTgnM0ugEaicvbBIxikSBULYtWD
tD8o6rhRlRkiow4V9Hx0T0qJfDFnWnUimCmTgH8acNDEDenrHXPpQn6BaT7jIM4DuwoQog3wH1oT
4KYKUuYfm/wHrU3GzbHYM6TIg/P/Ba3nrh9O8IY7GTY/q+BxjZaReTun+VWY1xJyZnWL3rs7NgXd
Bw0YIWa7n50Eg8rttGxK/wHMFfYLlNqedYmCMscjUx3RvnPjDgxJ+oPr97WGq3XuSTManEzmUZB0
1IUefKIGjKQcBtZ/9lDdFdRNU7/tM5UJC03PwSPrATCZo1FBbvrxhm6HNGoo8x2zDGRV3ZONuAAj
EeQhMqSD1ZzELACIym4/aYOlCn0ocQPdCAENx1Xn2gGb2vWFMbTbZxfnRtKWXbiumqf5dwRpnAJV
enBbJWMSk3a50yLXj52a6T6Su+f4pyJGKhrsy+QYfTQuxnXRptI7E0blPSewuMIdNNmkBqISQLGM
BHwRqd6QuIf6oSv6AMjZQu8y2xhJLw0E8Mbpx13Hh3FnGeDZ2J071XZ1ew06+e2rOH0wXeCAwEJ3
WzttL15Z4j5ddCNrtans4U7kryXFUtbzK+iQnohmasAvWUk/U9u/LtGJOjzL985ftJWhj94uwLge
wW72apuXDKXqZN26PD+1bWyA0gC32oZDW6xve4zQGJxEHNvkIU9UHFYrmlwui0XPkuj+tEdzpWoc
47YZLqo5XSjYSTCB07x8+2qhTXEDUgQBbzHhxAn/f6i4YUYyM/JYNOOSXKtx5F/+Y3+vRjLZ5kIe
hqBlD4QHAlhWliSDclutezcXNI0eX9OwljS7QrgSAeh9QqGqIsZy+oQpQLsAMh/Qqh2xJpIeiIze
wvqavWyvDgN0F37DBvYkwLgYU1XRQGM6xqaVk5hcMk2Cl894tXzLOPUddLhYsR3vWCD5SCs3Bzo9
h8fD30/92uJ6cZYplNC4Ng6KJjliYMQ/O9AcHB8HlyBaQZgj7ky3E54XiM6Vz6J7ERa/hd/6P5hp
wr/27awHr830Gc3aEK1AP5FEQYMZ0HWyM5zHUnW2p4wuhHY6M+xbaBP++zeiyaEpT7kR32tG22oD
salogziY5bScN0HoiKnC9fFtZSJBLvo5aXY2QWFoI21xadNVN9+K93MiURofstfmLoO4g3tDEehk
D+fnDhlGIU/46BQeQx2vbGXrIfB9Ec+VsFsfbjgjCYqnRYqHGQzF69a3tP3ivfcnJCwPuSd/QDS8
S/16wQv67XDfFgIQK1Jr+LUAjPXtTZk1V8Md9C5UBFItf8rmVtcA49YPClJKbn0VVMuUMuwnI4vl
UqX5JalNS+38owXRrHlloCJETpKgvPad1UHtfCSmybT43P4wUtEANMRJTXkH4khGSsr4fAPMSMpX
pG7efGOlAAir3Oodgu4D8kutayIBHPzWuj8W4GOBmRcsvG79Gm2BrWFpECy0nqDomasTtI0K4rYK
kL/44QEYzsVTzZDp2MYcoAA1euxdA1uNamdbhcxCcX8hUipsqETw8DqNIw6muVtup+kQEASH77UG
Q4CuQ4DFG9MwR18viE19Dg0ZRwSVMC5vRKBo2MrXOFUUM+Q1AAA09an0ZrivKPMLgmQ9FmhatT1s
EZeOxnRPq5x62CtgLYdf1+U99SrpJ8J3ptSsLhfkRSW8o+OIns75JHBPJKXFEzPf8+uIZZVOAK+Y
p503euqDxIo4g1fgeEmjc6oJh7PrcAxYmN3ILDj3TgiaE4DYxxsjRlWXlH7sWZqXlCnDlFa2lhwn
v8Rxg8WvnZZl+y+pwj/iI6/I44/LmOf+a9YrHMyYkcYz+CiJ7SfvBNGpdkud3j50XbkGKSsvXqwq
I9qVt6GALuTnlCw0AR4XjsDiezfQSdWKMJ6dBjaQnCbNIGBsBYGUEhz46oM0ptKv6wC1dpWTrO8l
XMohWZVpeSsq5ITBxfIeY0IMXxD6G6+UJ6+P8j4inW8bYhO6aRWbyN10daL/WrYy27MVyNHknxB9
HWKvEnMTeft+3+wPLXQUWmLvnRebbDqjnQczqTqn7ezjPOY0aUal2IpqHGIipqRWYYvxf7TOvsS2
+qUUSu9Rq8hqEfkGdXsAfDc3saNFSiG2PGZ5I+LbrBRdyDs67r1+LcfDr9v0zd0SsBSQs2OVbnLc
VfG4djv4fyjDrPGArSSlkOcs2+vrLeNE7nX6+hmidMxCmltvYXffzo/7vci4iSioRlG7xAzPfULQ
chwBgSHzEc0yv4RaREu+6sp5t1S9x8C4pl9vqaw/1rkUusqvLPdFIFn1Vr/fJO+5S6j9P+ln24NE
629jzqyVIue8ct+6ZPZTqtileYBB8EDQ7hCYBCN02FUsmjjucFv2She7HHru+DVKXKxYKvh/TzZZ
vshTl4vtxSZLrI3b3TpnZgLM4Cdha3b+U0kPowSNyHWT2VzSBgXsfNb4E6uVl6ENBVF/0PqvWexG
i+fp1+h3FohbMa8ZQ5shiE6OCJy1pEKuI7ykQ0Y4kTRQor+p2tNSdw71vmslzfdYO7EGiEz+tuth
hjPeKiYYFGyJoTd7e0YCO6xJfl3y4DHDz/XSdzrmJYAMvtGB2V95XbGij4cDLcyjW7ksL4f8eh94
zbuoACQBchnx3qye07pnv8yl4naJdbqqQXUf51INVY2Z1AyZJbj+ag3e+h0tIuXkmuK1QidkQYYV
o0kZlENIOyzjB9KcUq1jFwKCntl1h7PjTGYjhErTamEfB1L5MgKFz3q7/LuGvRcJvZUpcHoDnK6h
qAPKd+sQ7uXzoIllj7KjSniYGo8s1VzzpFo+y3KDCcYpJeJSp3HlvJqsE9CDFj7EYrrtlajA0Ogx
BwKKo1Wfq3Xy6GmYfMA7JQq74n4N/sjwnLYGissW+0A5sXN1W1p/wzXfP1+a8mClhIoxbj/kgMtU
kF7XDeZ5hrZyiJmuLENjk737M2OLNVsx1cAv8kzGsN4mPlyJYjcMJJiUQrfjw6OLY/hIFLMKVQQG
+q+4YEKKi84639lZQ2hOyTIr8BmylYBtkSctlkSZvTnTe6KxxRBbFmXljpIl3+idPd2yPtihjGFx
5sQXHroYL73uBebxGEmNEaevY6HpXVoMPiI59r3/ZgVpV1a1N92DcQsV2YnvAhKn6fLbZW9nAu3h
Kon797vc41QITBVE3lHKYeNLVBozVmsY4SWXrNtzUllPQCLmo0QvriQc1RkGItEbnOY9W8dj3ByE
BrWvQ6g+qER67Jb2HkEFH9qgN3vsltvoF69Fk1H1Z3WrdqH57twW4YezDSJeKJiF0xSwWba3ayvi
u+f8AU1/ncSCAm57zuxiGpZ9DqmqkBQqAMDqUZ7xNY2S/YYphVgpKtIE3I8iK90BFtiN/ZJTWZYl
fZK28h/DFJExF9sn4TkBl/MkpVkztCwQyGFJjW/QSUvY5Bi1zSjpi2wVL+NUW+d6MsnpJ1/S/IJp
tGGjiGHv4hKPnq2F8lQm8UDtGsZIyhXe6SDkFwYItYM5a0RnQBQXcP8juwG9O0k6ABfdhB6JalZh
AIriOmphTSOgshrCDxqy3NU2mG3Es7zSYaHze3AUW2oViqDdNP2l8VeZHiTJxL9SnAdFZP4YmEAJ
2FaLOqrrKV535bX3j5hFvEuCSiPyuvGLFrYjiJgJUNm8CkbOdXnUDzHjft3Aq6Ks04bnzZtXvIro
OdIPSCCXW3/a3fZK2t5qCAnSRbqX5HQYklJyuMcIkzr9655IMu+u4xKL2H298aQdmHSw2pL/f9xE
3uGZD6IKB5hLIOjZY7sx9kXj0Cbf9So1vJm9hpXzVeBZWmnAh/NC3zYg/wFX3WjW9gCUYY3ixcP8
3ISczIt0n5Ik0xdAeyB0Adwi/GpGtAGnJpcJJy/Ojr32LxOe98qeJOCjMVy3jHwwEMTxJU4di0wp
aVJLNRBzxDWzlXvsRgQn0ZZ5AT0ZzBH0IZhs0st0FhLK80xY2/6lixEROOefgixETR2jFB6k2gbW
BtNUjrz6OSvYKM+aWKpjmZCfLBtkO1jpOYcRNppkKnQogdStyT4DrJ0j/0nfYOMAdziwkzK5cVq+
Mhtr0BNjjrr3Y3mFxEXmmTkP5EPaMmwpcqwxqeiV2gaV6govnHhnUqDcW45ub+ch4re2FdMqZpT8
vHx2uybZHNNcsOPjxZdBA8laYHi8j1eoKizx8tDyRRoRyO6UhJuiZRIXKvnTZLpH5Wf2VmRaaYt+
6f7hm/pCK1aMnVfcp2+DkVoOmtCwA1dZiEmRF3lrUHAAY3dTDcZRgk0X7NQSwfvNgsydtFz582ku
gjFYRuwhySVQ7CBLjqGRvuwWRwmbuHiU/0cWtIYCGKy/Hpk/R1uAPwCZDK1+2ng72jkhYnN5gDWD
JeALqma6I2B0V6MtuYIYaI5Pea809ROCRpw2Y0YoCIMzP+BZehlao/gBear6D0P+6AfXOcjdIXlm
3QpqYDN6MB7fqf7XG/ZwV1gXO4iDR0mR0/G3AgKbySYsar2UesqubCGViU6HXOp2QI9lA26iQ+en
STq7T/Gm1HIv8phYbaMqETbmX7daDYb5pzpnDqmZ3coDwfsMy6Vs1B3vXVH2NE1A2JZw8RWCqNZq
yFah14tWeUlpt0g8d6nsNmwl2kerFo9muFAQmeqkhVrqIGfplgTmuso/30nfrleJ7Hi8zUypqycK
15gfBHVI+iwerlZMXt3E4RzdpS9nYCbhLheV8YYkuEp8P7+xRjRvab/RPlZ0rr330+f/47pYbC16
666f3wLQplNBO8G5P8VJYnDFg9CrF8lf6vHE1DCauUw5qUakyiPPqGX5d+GLuKvZhZu+j9QyAxQY
iNcHkaD7NXqUzLLsT6IkcKIEiB70RA1SMfgqVkU+AoZ06WuJq6Wf+cdVZlFZY4+ZUFvFqWFEPW4c
CjGj4ps86SjvCrnro0t1jIuBv654x116c2t/llFa4zvHITMy9WMga4Dr7fCUAd01xszkk4SrsNnV
RpxzgFKorW9gcvYfx4x3CsrF47T3vD8jOkOpWF+lT60f3HAT5V7BeXRl9CTIZe3Pj6/WHlCIvurX
iiDUB1mWemTdq5YVQsleHFnWhbdPlCkOSEIEeh3n/3PT5m9IgrmMVW8nc4b/oa5Cq8fcAQ8ATX6J
YGLnD0k1yQqjWGqSX90UHa0zgQWspfIXBYIg4siQEC3p/0dIW0TPt15xxPxrfnDVBEnHYp4NFqJX
UKtD6O8ig1bEgSQzEfOiwFxSHAoNgnSVXkAv/3wi9RM3WrVeu+9MpqEgoFZD6f2YMZ71RJdW4Jok
rWfu2DAeruFkiH6Q2pyNwGJGYEk4EGDQYlUP0umnmBS+zWu2Q9yc1BpyWooWBqkOmqu4XgdUkSas
8NBILgub1rAxisP4tq8CkUgnSoTOeJdm1YSeqwnZd0DEplfy6Mo6nOkL0ccr8txWOhIpW/xvukBy
eZrWEGNmGs8YJrO4ZBwfFSg0vAdlezZZqHgk5i6uzc7tf80LHkJf5XWz22aKnfdmo88ehC3exumw
wrr7pJNfpipN8F/n5rD3lzQumsMgUuayV2x6YRXRfijARmPiD6cO052fhxZlRATycZ31eVtLPOfA
DYTCgSHNOP3DYRQ/yg+EB1aqrsJbfRZ9I5C5DxzAsqW2Ec47DKfASpbTkhzIvEeZ3ux8qE0yoWKm
w7ppS6MjMoGWXdhCOX74Bz0hOLWOPIz4YXLDQ5siAHG+5qqwwFo0xykMFaYLtZcsTP86baIgSjyU
BXzE1tyBZpU8YeGuX0ZN8QRvwMdEWVwdFlY/vlkWm1oaTneQgkKhU0dip8NahMXL4Ik/CqBFhjLR
/lcizQsZHL+cl1nl72LWPgs0QMEdj8DfUUB7Z9y4kpTiyvw4qavvoZp6UUsi5YdPJqu8hXD98kmV
YixzJzIsxCBRCkDOjXoQ90FQ/Z9H+jtqtT02XtoBdO6gd28vVTDkse3wcHU8g8HsFsEfJ6hb1gYo
ebyW9cyrKId6wjbrVPu6B6CWNPTZc45eB1v22yBTbGV7YowvvBiv6FC3ctGIoP27Awm7umbTjdvE
L3d1hfB6oqHDKxyJc2D+334CWHIeDnfa/bK+NkmrsIHXAgHYTQpFIblacZxtG4ru/e8iXz8sywm1
IpwRQsUQCXOZAGFPR15PpPgcGTC2uD1htk+Znoc4aapcekXsLGy+ZgLPft/6lOFPjgu8bofblD4C
6aKHovmNhjtdGr9w1z6xt1w9ho86ApaWJgAkWdxBJaRcYq4AnCKv+Wu6r455mz4lF74gMRZ1ZBvw
Eq8YsTX9a0ellNg3eTne/xh+5q6jP4UJAjH+fmXqWJb9hefliiOcaU6yO5DvzmT9JTxZQRMFkYCD
5mY/OjFgLayFxDJVrh5a6fKPRw73ANrlTV6l0n/DAJwenZ6lHNYCIe0Vlfp+SfROwcCzbIj41Ufp
kgSGURq+xXR50eFqkweszTlWxX7RCWogcg7pIau1+bzUlEIuUxLDqm3ZuJmuc7JCf+Tp/ZQG1oF/
b3QOrcbUjB+YA7O5hTtnVleae22q4Natz6CsuB3GpawzDa7jOk6EQWIW0SejYii64e7NcKgv4ppO
sO8g3AKjG6xMq2O/inY5ZRCqUi334vH21hqJjVVxb9XqgOi6jiGNstpNtd3ICqiS2yw+biPI7BSQ
HBZTtnXNrkmKNaDBzIeKXecTYTbpBBw2ZzvF430u4+r3BT2Y11gbCPd6o1ec4e0+r5dbToNSR1CC
O/gnwN5JX3GXzGeVJw0EHkPnKKyaC2Ra0VB1RR0cxAsBYj0lsECnAYYHEFpQF3vVvjMNgY8T4Bg2
rLg/Br8pVqEbLD8nMQVy/h6YnQ1p1Mo3z92kNjch8VBuuXIY/684ynPhX2bVflEX9MGGM+EjliKu
Do4TIWcVLFsDMjJPjSXWjPhi8vBfChRa+oD+uIv6D1LAc+DwwScdfyUIVBKswanKRvjgalghIUjy
yPZ8/yzsATxNZC8DzILpGRZ5yTm6bmy9ZxRXjH3+ntd3K592RtP8pjxCVRvh5ZmcRyPpK/TPcq+u
K4QT5ajQECnGr87jbU789fZR8Gktw/KenXLq4m4MRebaPQI9GrNx54RDbSnZVsxbzik9zia9+yxn
LDsBwC7GdtcXB2+LemJMyMr7SnqifL6KKlvvUBlcxUANaVCnfRMCVn76Jfz9OFWa1gSPa690jxDl
RTlroZR4UZzaO/D4TOFXht+MOMYqPPeuqVIb/IqHBcrPzb/Ym+nhpmWQWci78eTsyA+0Y/U/XDo4
RQryANhSyQaa4rd4nDFXPRhje/ws/vPycnVxTPWURnHB92JRTTJlhrsIPgSb59MyMrcovVAfixYs
1qu1vKGcopEyjoZHL8mkETORekUGIrYAD8UYrzSi5WGRcut9i4dmjkb5jBVmZUN6+vrGcQSI8swt
/TzZREclAtrcqwXLFN8qCaXFBeLWui73nKUJUhKa8JzCUdzeNgrKGueI6yvM5+ZIR+kIDb5wNueL
FlZoF2lksAGVkE7wIws3ZsGSb5gzJ2DpX9IXo+ooTqrDcf6SS60sMqKy2nshTpCi6dpWejiCkjt4
07Kw/vbTt1aoz3m7b2QWJVq+bTG/+hqHRliHdQ3eBELA9QaZu+Zr7jeyirdw5jTVE441clA2RaZ+
gLVHQ+wj4CeRlWdrTcsT0Pa1JSuMnf7hAa3KgseDiNChaeRD4JUSb09ge7S8kWvbKvacc6J1kFw0
uFu/z8jd/r8BoDYefeBNskIpLu9baQDVlFsZ0ogBH/Fm27mB3O8cJSXi654wdX0F5wIwE/4Yed1P
yCTjfOK6fVbdFV24QLxyHiV8P1MsPrQPwas/iBHOkZabfOGTyigKxmqcRuG47FHfsc1TIrU7r8f1
L12ySM6y6A99i6vmWkYK0es3aUEulwDnNGuxj+PIl69GYpHuAC7Fbn8MVAscXQGEExQK0iQwT/WF
8S1MxJ66S/xHSPk+7iWOBxPBKirMRExYQebssQOrtSeWgWuMaIIfF7Tl8Ew2kk44vLzehCi4rJGu
ETs3oJ21vsp9I8iPy2YJII0SRkvhH/wyNlJyEU49/SREUpGTNxnP+OmJRGdBHiIPiKsZmRd0/rrO
fx0wzvWHcNGe4ebGVZaEdBASe0wRO4kmQf1CIoHBli9bQT71b0aZV83luKyZHdd2G6hGYLfuX1GX
4TMzizWEIup8axxQBh9W6IvSXxc2dqsqJ5ghODNFiZ4XdIZIYDDF2QAWOkCn8pXCC48vmS2jaFxM
NuE+tTBMXdr+xOkPVi/yNucyFm2HPEo7c3m1W6a7YXgaxMWFs8WT+gF788DHMTLy3c9UrJqUDpH8
T7j0sCsRK39aAvnGgQ5nJsn7m3KlGTYelIRzxWRm69uA2VqAahpCJ5JnbtXnSTSKKI4HrFM2zGUY
nqgd/k6WN4J7JimPx8uTodGf+/RV/laeKToDKiJ8kUmYA6b6Yntx5XBzofhbkRZE1NwP
`protect end_protected
