`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`protect data_block
0USWSUGxovGsyBJteYpEoTgLPudcQL7WKkpu//hi6TrqA7+52dzwSByTrmJFv8vLmeuvBugWsQg4
Ybq0ajV8lw90tdj3OQPCNVE6wZs2H/Aaan56x9YmuuIWKiBFARmspxGWj6AGyQ2jA3D9nwxCHDg3
KzVLdVX4e2vJf3o9CPQpJ+DsbAZCPSbo5brDaR0PUd16a4ReTh2u4ZqF4v2RJPBDCWyU8eMqpcea
BDY6BvxqYutQhi/+5kfZUtSf+vJr9m6pC7Scyr1U9GctvFRREaQ5SAhqFLx/J91XmJVLkHbKgio5
dMHHqm36zDq4HMuedLJTyLArxnV+HVEHYig6SylR1JNWcdpcthHlC8fV6N1dcXSXk00ya0cjPnDF
lrab+tsTUBG3yYun3sEWLUZY8bq05Dp3Enabl1GPs9NABgnaZBAHAtA9j4pkYX6juAWZnORKvLpK
2eyC5YuqiPKmcuK5rFFTZlMUwQuCVryDyzQyNT/3mPYllC//RbsXEB5QgwJnq5TJOv+r8WKlRfSe
Hiam6QhQptC7VuzUv1SJOq3HvhjkToQWf6Jf8VeTOsrrqdzmzKpi+P4e1hp8s9boNCN3hhkh5qpV
iKIV8UWSdMjVJi3XHRQGWSRaSqPDoR+dRdliR5zjivVnHEz3UeXCZj1OaJyllYHKObTczITxbjXh
lOjGx44h6YuHkdWeCCoz+pi4cZ7wRIx0X+iJivYxm0nxxDPztFoAqwb1VOtA/QB1sRMBL1O96fM2
Xz7fjY3GUZQvVtflWh4yPyJ+KIsl5a9Gwu8ybcNJnAJY+u4kfh0eFF4jxL7yoROFYiWCIYntMLUb
MiJBeLuPvPaFbxGCvXKyXKDQxoBJC2w4wEsQDcu6FeFVhXkLaApKYoH0GmehAlQhZ1YyEK7tugPM
MPY45HJyZ1Sl/K+WfLnD85A0u4mqEqfTJ0D+s+avO5SNgM3Llctqpc2xPFZgX/0ILNdq/a9f4A12
EkwPF4/AMiVvIqZBhWOS3kk/hbCIKmt67xusa/N8BbIFoP8UYS9ebpZR9EPuV+cDckQPkaCsoy/L
/unf/0Ptq0WKNDm8C+FgP6+DEZCrW/H8h9c8HwNYQaTOivPtEx5hAkGyxeOa++JREsMN5YI5haxr
JFml3GB2B6EgL+JS/sxEJhVs85O3ECDkZqCcSwliZd5H5bNLqpfxsjrEzFCwuhx2T8fLKcYbnx4w
5qK2qI4M2SmirbHdCm078kFJe3oaXpXQixCVSUSFMXaC8FXWjoJrAgJtAdoQe1VQPJCguACoW/iD
+JbuVBqm4e/3084ZURSJBkUutDsWaod624DKoyWupYdzlTcMrehucPspeYp9zLUihvKsLiPuLHr3
IU9h6gloLyMng6XHQxB78y5KRF1V+dk3PA004fEzYdPpETpjKepSyCZsXTWv4ocgiZ7+HyeQbGo7
DOGWIoUh3ppnutx4DGyulefcwabrr8ZII+QOFabO5i1T08ABafW+dVZaZidIMTv5yhU9em62LUfD
sk0J3YHKw0xIMWZJXGqaCY6A2fxHXYlx7AMthyOVaulguaovoCpEEC7CEi+2Hv4Hfm0jrZJ+GQiN
oRkFKw+pYqs6AjOGdHbGIurBhztqVKrbSaZR2XMEWFNnlDpxkBH+sbTj2rFfgoRpjA5dtsUMWpBf
uvJ2ta1XlP6sad7BQd/LCyAUxKN1j2/qMq3nI6prDs8T94rp7uzYDO/DAzGrl6b2mgrtmOQWFeR8
qjPgB6pebuRZSFObZ4VYI3LZDWOFzBYf9JG5hHayOMy3SSJJMv0UXpsj7bGfbCBpa201drM2iIhV
MDIMCPEvaHFmqLicku6aGLD5Glrv19H+pdcYbd9/uUdXIqJ6hAJoY2wWQ1R9Wk8cmqTH4ASfXjpp
9HclzClPnR69Sc9Qnhx4iRZgI0Ij64a7Qh9AfzdA7lsiORGwWi2d7RNxQYQwoTVTohNu5sU47Sre
/JdQ+wrsDFoBuagFHdUgRKp1chkPZRNrxy4//guYzAl6QbyPSYnvUQQu0qNwOjj/KIu3dilcUaA2
M6rQMkzxwRnbwnjm9rBU60y/SV1mkH8y4niZ9dI+IYVy5ndMeM3va4R1Pse4JmopLF8ecwfpfFor
QKfMEhux61h9b+ApOMBcx8BNWFNglBaZ5T/MQao6UYYDuxOEeAWceU9zEFCkJsQzLZ7+Z9R3vo/h
R3eMpIxIreCGt7t7G70JpXVushhMZcBuWzfWK2/fGk65DO/CzzV576ZkVfWqPOPmwBn0lXfpq6Dr
XTXFdsVTVBy6NexqlQ6DCcGX3jjwmUyF8ZcxnyxBcxg2XTm5syx9V9/MNakf2s3tjk9/9M542dCw
Tm2P+emSD8tbOXlyR0P1dZAJ2NCS+bnY7eVc+zGNVkVRjVn9XglKJvm0J9djJO0XP9bp9eB7Ljsn
glm9Tnf2xD3fdHLNKi/fNsREoYglYIkDhc4OLLlAMvPrkAK8kNDL5jU7sI1nMNEiqELV4Bvuj0e3
ZKtyMzaWHbO7lrdQRvPDVj9cBa8GD/Cp5B4+fOWyLY/1CYKsBs+jt57aCANGLfA64lutMDs0uDDS
BN925GMdknNLqcO3WneHg7Idc3DrRiTfTFpZqUWZanI46wRemOWG8MUBFpL03K/GA+naawqIeHfG
qbxYroEP4Z1YZEkkp5kRMaT+uAkgy6ejsXMEnM28eInAkLFehYHzsOc+XLGqc2dngfgCf89hfh9D
emwcapCHIegeD6WvZd4En0FaJJwW3KGss4ZoZFCyFEnE4ynK0evMy6NqM2JGAEp306RXiTZ6hejW
sVfdaQGwi7Uf26pNisj0cLYmiS8lWtzMeZAUVKL/HcxmnUKGf8360InGSLsuzfRvondOmXlzvViP
Wrb3kPYRr/M8vnwlY72swe/clUEq739zdeRaKx6KI5VQbSUbKHXRDypwoVIVzg5edJ4sutICBH9S
c+65ymQKUsQlQUBbUuAsvDgkEjjZNI1IphXKBuQFgOVT5Ihm+O6iB4zDUhhVrG4oQErCboH/iw/k
PN9NTS44wFVYdzmOoBr+YNBKc+L3GtFwQ4InyM1lbh1JWf5YrHGQQpse/LQhlUOoLzR+QCp1nGO6
4/VvvqnNfbeifjp+wTOCFXN6Mj0aQwalUhGI1fdoIYWDFbNizOoOPVk7sAKEJzwVRkDGZLkkqlDm
Ld8SZo/SQ51wmddrxDp/TmwdWm5S8VerQ+SU5p7jUD2OWqOxd/FyK967/U8/6MfqpvASsNGDGmNt
gzSo6SNdrFwkDP1ABSLwcrsZj3SVuqwMYEYNfD1xmM+rjBAiNWX2vMZDeFWhavNYfXZ9uoQHcw4V
UkN5QEHUS7gRGpkxCi41P3DGbINnpz+AY2r6bd1usoWf4mqkHUoIKJDw7jtAmqGQRmMQLahLRbzJ
oO0TQhTG2V3bDm7RhWKlG2Hhj95RIBbiZ/gtxq5/YxhfE5jSrSSIYtKRMOetE4pISk5AvdgPtiQ1
UDSlnKhPI0H/m+YijawcbSJP5Aaj9eBcGc+ATJ3YUJYNTA6aZ6DivpJxGAVtf7gvqDeuAK9qAVZ1
KZ7Txmgx12U9N7NtfgLveaXkxtyflfUUDgMTj7uWt6gywOLbLS6IF+6/CHvgthLSbBmx49S79Guv
FQXtd7sbHE3A1A5oFxllgV794pRwMZXgXHypfu/0+bmqWMxgvacI+IISjXvT1wNXhLIBaam6t9NP
pJmmta6OhtvhAMOpXbM1QVvOLVbrpHneu6dLZpyCfKlMrM10gqN3VTqCQlRcTMSoTg3ckhC5Oc7P
Qx+b2Mm5DTqGO6zX7DazprD1GiIGHL0b4iTa3tmlnTq714E2Yqs5Q2zpwSMnT3I8cq58hrsCCeLL
DjsMCKeeULPomhzvoUlokP2J7ieEvlLQ1mUGHlqLLjh53P/O5wDqehfN2uOuUMAaTfwQvxipYnpt
3ry1u3R6+NkK67W32Qz1qgRHEOoiDys5Ln/wStjRh9MrFQd3zIr9PIDTFngJ25j1n6pAV6lVj+3z
amepQ8BWj6VwLLvtgLr+gRpbhI46WBlPY94VxSr1pKeGRbAinbX/ipQem68g4EWQQBW3Ae6JiFsj
WfM6+Rh9gFNR1CnXrK+gnW9HytIipFJtOLHvCjUV6rqX7ftr0+mY36FOEz5aZG0H5wGTmilvfDPr
MGU0kl1GhN/h2sPPBwkV4aPZ3HTOL5k8wkmZi0rHhZNEhyBrx5AgOvxxyznoAIe+YMkYt9tEamdl
nGrqiakvIwsuIpgFRAeefPetJmld8ZmQOMqcZQd8Ag/DDkOij3NNu+jajAcizUxmJY7SuS2JFjsx
lWcMpwsLFA0r2J9/JciFOfCITgqXw22V7b+DNBKlvzgfe2xvFTs38wiPtEsnp/P9XPdepLotHX+W
g81HTfFqRj2mNguqpnCDD5ET/4waXioWoQNiBpm/pVkBW7MP/EBC2ORMqkRWGyN8xfv9UXoY6wix
6lXVEeDT+mXdajRgsj+0vJZWR6hlvvzg2jGSnbrsV3sPZ534iwWRvSH4KlOY95qd41VwG158551G
Xdn5VJRvKOKqu105ZLFqChWrBH2S51ABTY/Njuksnir91nrz2ETlXzPBl317UVQ6aq4nJQNC2Flw
RdLr1+H+lWA9eeprchI4loJb8hLIIqzv0yVr
`protect end_protected
