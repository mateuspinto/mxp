XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��.>��P�W����&��p�d|�lL�#0�{���G�"tuZN�Iq_t'h���uo�(����Z��[8�
��їAY{�&w�H�k ��Y��4]��w�q�WZ�7�36�5�

>�	^��>������&����9(��z�	���Xao���(�OD:�Ɂ�����JRHq�'�Va"��x����0C��P��V���J������:4�ѵ��h��b�@e1�f텚�-���uLhwQ�������6���.��JS�9^s�cK���=j�W�_��D�|���9��9�EH���ð\յ��nb��,F�N�}_ J�^�p����6FWQ^#n��q��k|�;6�V�:�4��O�\�р�_�1��P�ri��ގ��3�����ݔ��tG�˲'���v��7��߰�����@1�x|�`�����]�TĪ����^��j� `�,����
Ep�-Hr�t���S�Yǿ
6�ktSA��M��m�l�(e�
�����6�)�@�w�JiD��Z֌ �1W��g���32Ɋk*�i���w��+QT�'cX�re�y��F�S8���ͯ����4���.ϧ��,vc��Ê���8ݏB8��U6'0�����Җ;�~���>�­�X����8e�|�-J�"����Ҕ�[:=�� ���xY���#�K�}�n�^�z�%�x�|򐍰�O��J�%1�'�#�c1��LԚ�=�f�;'��u�+@5������}�j��{�XlxVHYEB     400     1c0V�]@We�E�%M�S�\��X�K�F�y?q�/}X�uK:�ȑ�׺�TP���HV�8nuM	�\:5��,����_�&�����]�KC�4EI7�s�H0Ș�"��Fo(r3�9��X?����>Q���G'ӔW)�3?.�\��&j�#���FeDh��%/q�h]�S�a�yY��Z���8ùb��&��W�`���LpA��X���B��^���� +�$uIСP4��Q���ԣ�F��YR>�/�)� �T�I3����
�\�l;k����evI�1��m�v�- �3�RsV�d�4!�/]��G|�޴��3Gڋ�!�	Ӏ�����8p.r��sV��"̳O'$ǣ���ލ Q�n]�����Yt�~�Tv	��te~ZWNvK��̝	C�h���<*�m�s��G�&�3@¬��q;��XlxVHYEB     400     180O�5��uLK��L����F�Zò���<C	�ɅK�����x�[�:�^�Y��D��Mt�8C�_�K4�7&m�D���7U+r̆�߄'?�qf&Ey�M4���� ��(Q����C��/�g�@>A��w|}t�o����7&B:��N�������k�cM������F�F�`ݭ.muP�'��81� �!�����yP&�8�N�_Ss	��Qqű��YK��G�_�L[.���b�@>��}��|V�KG�=Q��N2�^��_F+�����������t�dQS�VZ�	����e�Ω�<i���]�̮dM��.D�R������u^-���Ƅ�=�{}t��R"t]�/�r�u�I�f�n�[�XlxVHYEB     400     150'_g|�!�Fi�ڛL�7B�y���m�.��C�j�3�h�!����"r�>�&����f��/@>_G�6�^��i��/Ƒ����]�EZ��p��c��;%)�i�i0Y��M\U�/Eݏ#,��,ˊ��d�Z(ËOO�0�	�?,t��@V�U"w��+ϱkC3�������(ږ�7��L�#������s�LaY��`����'��4X+1��r��`�B��	).�z�QW���o @��P���V��)ޑz܄�"��.Ǥ}ե�ę�����֗��imR��/��wˌ�G�k���ĞCW�L>���9���a������C�p�Uqh��~�x��XlxVHYEB     400     1b0ecT�&��b�E��,H.\qP��q��[���	Ef'|싓*�DL��D!@Z�Wi��]����۠P�A�`�"���D����Q����}���p6��Py�p~�q%�T,L^qf}��p� 0�x��H�^ s�4ȁ�����K�.��ia��E'$���"�s,{^�ע�2rlY�����/�bm^��r	T�����2�@��!f�z�I�z��ҟ��t�����D�J*C=�2<�������u>�O�9�����n�/*7�{�N]�R��>��5#��j		���|>�L�#��2b|v½,*e�e�Dz���}�Ni�%��߁�;����=��ρ�H����
�Q%�q������rP5jj��U�#�Մ�#w\e��%��?L�3�x�U�}u���`'��A��/w?�[�4g:�4�����_?�, ޺�wXlxVHYEB     400     100�O�oŒ���<�(�I����T��W��A[K�e2/��l���)�bF�P������g�ߔ�c ͦ�&����������A�qx�Vij��ZPvFX�+�B��h��tVgg7��}_&y��:84�|<}�=�۷XrN � �J�c<��Z���.��gP���C�������'�:����=,X�X�o⻈��9CtK���n�@>e��䘯넵4Rcp9⥚�O੄�찚��̻�$t�XlxVHYEB     400     120B	f�90H	�~�\�L�#�C��c3�7���E��rd:A���n �$�A;V��-��	��-���9�$Hη��a�j�a4����w6��5[�:�W.M����:�;�\�T������W�C )��#��Ɋ}��v�5��t� /��󣴟?�|�*�����`�F�⓼��8�����(`�<?A�t���q��0�m�M4��_O�� ь�@��6{��	��cT�`f�q#PI	��Y,T8��B����q�2%wB	-��x���`�fu��:mD������XlxVHYEB     400     160���y�z�E�N����g�7�8uˢ�kOe\���5J�z[;`��$V-�sN���]��$�Z�����yB[�'������0b��Oi ��
K�8(=����rUHM\�ⓥn�f���)i���8`��\a0o7B�L��f�O���a~h`� �b9ŜU�C�!���F<�H�?e�e##�j���Յ�-?������M[P��� �mfHS�c�e�W7��o2V�4�tA�FVA���Q��m�NN���\�î.wH�����T4���
�}�GE}���g���P����3 �GR�?���: -4��Sr�R�����;�On�q3*�sC����;@~#����o]~F�XlxVHYEB     400     110ф
�-���W��Y�o�^��e�0ʒ�b)�HY�x�[٤�\p�ˬ�2�7z�BU���Gm��q(���M�'i�E�[�޲�R0�e(VO"8�'���O ���	؟9iI����;�T�і>+~���p�X�{=��+M�O��bE�Oؘ�)��c;qB�$4p��2���90�c�.c՞~Q����Z�3տU�w�F���^���J�	6�gs�ӓ/�ȅ9!Sڬ}}���96�5\>��޾~�������X띴Mf����b�#]XlxVHYEB     400     100d��z��zq��O�~�^����!ĕ���(��_ۄ�`�ǠK���r:�iMR;g��A'�&�</��d_�wX�O�n��^��y�Lt��`\���Y�6���
H�E[�i;�x�Xd�R�`��i-Z=��J�؈�݌��Og+�͗n	)��^�6�1J�yZZNj�f[��"$��t5�>d�%>Yd1�ŝ�2p�1(&�r�W�mK�E�L��<٪���Q� &K���('&-�7O����BCO�XlxVHYEB     400      d0���0�K�kh����,�ӧyZ��<�:o��B���~�;T����
LnH�j4#��Dw�ݎ2R_P��K��� �����IiCț5Z���|TBJ��L���@�L��s׫\E�_���1~�ꡨ$����ֶ���T	ѷ>���?_�S��m��2cQV�XƐG�*��J����d����Y�wՌ�È=.����i{XlxVHYEB     400      d0�u@�H�E�Ү����������G{�K��(j��B�O$����2��4l�rp�\�⋿�����g�S�G���d�*25V��l�(9$7-Q�⒃&DȦS	GC�s!��q���fxႦ"x�s��O��G͙8��AJ�֮�2��`��J�Q��"Œ�
�;�2bj�������9Z���Dl�۸u��}�Ls�� ���f��XlxVHYEB     400     130��,W��$�eF��_��!Zg���/lԘ�4�ƹl�{J����o��>C^zξ�l~J7����U�y�e��v)E"��~���DJ��������?�9�5���1����c�>c��p���Wc�3o_e�$���pD{��5��� �t)����s���S�B�7�m �򔨸��mE���Da�����sb�;�I��g㳯����[�κ@�.{c���@����k��y1p��w]_ʦ�o%"�-AV�ȳ�'�CI2V��	���P(��G܆���祿mh�2�KW�m����XlxVHYEB     400     150���)���(O���'.�D��0aoȅ��(�$��"0n�]%�(�Ѐ�D���"��/��Cel��+��A^ƅǆ�DO�w�|o�S#��ٟ�t��8���$�;���8��HJ���c�ܬ�9)V�w:��s�J~�1�f��y<x�vַW�q>�(�7���k	Z+��H��H��sZ����y+:��2�"Z7vR���e{���nT�(a�wDΤ����c�{�4dJ�n�Ű.���5�b_B�"8����*T+"}���X0��e�N��͢�~K��m�lF�����_���Izu����}��Y�Dۿt���i�����<%�XlxVHYEB     400     170ߒi@~��KV'�Q/p�� N�ρܔ���������8� �7� \��~M�d��I���K(�Lb��_�Pd���8/�o��5ߋ����|ԙ���B��:
���jrexN�5Cmvb��n�N�RQ
j`�-I~�t��>�ʔ�}�s��e��x5_Ǜ�S�$S�������MWc@*G���M`�������J]\�?NH�Ԛ��tb[�$D���v".~ur�����*�1ywj��5���K��P�|tɇVg�Q@� ��ԝh>%�-��nTR�D8XWn@�|��T��1�n�n�k���?�ٰ�lJ����'�T�%��a)�RHه��\�
-FJE��B��N��n��XlxVHYEB     400     1902J����4hЗN�Ʉ+�/�,^�M���5�?<�1��Ӹm&�_�Z�^%�,}��(q�����i�,<�4W�J���:��&��Y��:68��3.Q��eـ^�;��@;؝칟x��yХ5�����3j]���l�Q���Ϣx�NE"�ȬY�I�n��X D��M�s8�/3��,�=�jo�)��n[Ĵ}����Y7�����_f��c!�M�`��ج�m&���2�X< �L�(������r��zmg8�����T���\��YUSϡ�$K��a�a��17O����� b.�Jr�]�gJ��B٩�`�s")4l��Q�WGH��8&�Nq*&��|`�{�.\���hkѴ��	�ۇ�P��lO0<��u!'�w�ԌZ�ru/n�XlxVHYEB     400     180 D�d���RJe��� �#�Fi�pM�>�}���!�3r�	q���u0�#���/+�g��jp)���[��X��7���S�6��
SOg�@/�<կ^?��x�1��'�� ���<�4�����r����y�j�PP��t���3rU��������s���ĿH}4&�6�<Q�%��,s�7��@��U�6S쒹,�;:��$��sb�G�@(4.�u$#QI~B=�Ge���D�'a�A	�X�/�jh���K4~��e���lDɿ9�]����'��"A�H�B��{<�R�p�H�dT�h1�g��F �� wC-L����rR�&�(��b��A�L"�}�3m�7Ο�w�l�wX��e��}PX�	�ӂf�N�u�z�XlxVHYEB     400     140�o��L�[�	]̫�����Sx�'l4zO�vP��DJՎ�o9j��x�ޚ���
c;h�k	Vbo��^�P9d�I����b|6?L���޺h�D�<��6�M_��\͝�<.��,�#3?*���	���E�:���SS������暅����G�� u��6\q�:K�3e��A�ie�2B�vA&��%��A��*]�i�zzG����S�v��&��lA4�W8ԏ�_=RC4j�Ƨ8?G��F;������0��x����� ]��n�U_�����mc��ie���7�cm�Y��.XlxVHYEB     400     130���`6�{���t�Fy&X�k�����4���ݘE���y�!��/)�A��T����-H)�l������p!L�i�[�QfN��iK�Cf�>�)�Dq��x05Cc+�c��hl��bFWDai�G^X-�B1ٖck��Z>�[�{�cQ��/<��`�����+a;GB�{�ug}��U1^ӽ�cj{��.ma�J��O�T��pz��5 %��#
��n�>^�O��>4���2ք .d|w��I; ���\�oIn�N�I0�r����tF�)��Ŋ΀q�����f>�R�XlxVHYEB     400     1703��x[�\d�.��nE o�|�wD���u�������J�7
��T۹��6)����Iý�k��&o��F4�nU��CIsC��h)�Ֆ����P����8��8�tE�ݭ
�`�M�R;���jW@#�A��@����~�#�oV�QHkI,�z@Y�=a�l>O��D�&]b���)��14��J�>��JF�������>r����9�����07�����k{�������0gacG'%��`��)����N��\��Q����%��tNg[��fk�0��;d֥Ia.~�X!+���LC�u�#gWj��2$��H���fV���dթ�)��j��)����1\��x������h����6-��kTXlxVHYEB     400     120��|�!�m�ސE͵�%���w��.�=����a���o�Y��.m��f�	�cbɕ3/���V%�����
8�����r6�|chdw"��r ni��h^C�1�Վ���(���;�s����)�xǡW�:��	��]�0������}ٷ�p�_�b�I"��b��Z'QCY��*�Ѭ1q���������ҝ2�-.[�k�v�� �,*A�@͘Qt&l�-}(��=�`D�+K��C�^��c�;hp{8��qY����� !LT�+ N�0��G�XlxVHYEB     400     130��ַ{����Hp��{b�Z/us���d����Z�+D����+�IB�ڀT05�o��Z@����!�sK��.��a��SK~ߕ���j��xD-Zwx?�j?f�,�m:/�@�����!9���G#a�#3.�/%��W��TRqw"�M`-&��^�PJ|�n��*��6\>�UM�c"{X��-$ ?E�v�G�[E�ٯ>�������;��\s�!UP�Q�*���6�M�r��䴘ݸ�b};���h��ah@(�ÉZ�UL��iZi�LðZ�ߥd�����L���Q����>XlxVHYEB     400     140q\�_zk����ګŰQ��ґ<
�H!W�bg���XU�?R�m�=u5�4һ�q�����{�&�T�Sm����4�1[��+��� �h֣I�pÿ�I� �DD3�	�ф=����(w��+�����4{��-��w�a��7�a���s��O�E��Z�#N7@9��$�c�����@H��:��F|O��%gwP���E*wgM��u���b��ʂ��M��d�a��>��Ճ)��o����R<t��8n-y(��!��+�'i�����r��(����@YHP��f'��j�5̦iRɛ�7���C� 9��
^ҡ�9� 8XlxVHYEB     400     1a0��Q笾	�l��n@��_b��Z���e盧޺*Wi̷��[�N|�Yj��It��"|m
��;�U��<�#W{�i�X�o��,�9tnveC��^�aE��Q��A]��8��_V��� ~��\Κ�!8�B�����N�0�j�Nԡg�9L�6��-�����b�A�t�U�.Nzy�R��I)c��g+;�߀T�[1a��@^4�O5��Q�M��O�:�o�b]�@H\�%Z�YMP��n� ��yݡ��1Gpcg�iQ����r!�ꊔ)z����b1L-����~
���b`� ��k/,c:�Oa�MW� �zƣ.�I��w���F�'L*�_
cBkR]||�C�z���сw�x��oI�z܉)����8N�q&O����&�@�*|�ʌ�c��G�Z9����E�*G�XlxVHYEB     400     180�0�Zn�"��� '���*4�~�/����'6�����Ӧ�������s�X-��ʐ�]�����ʧ�$��1��WY��sw.���<�}p��廬�X��͙���rXa\҇:�c��`LJS+m>�:t�d[�7Z���KJ�Z]����k)tپ���q���5�@s��RMGl�1	���@D"#9��sl<���|�W�Y� L�D;�=��b�����W�Bj�`=`:��|Q6�1W�K�q�~g_鄫���~�q>ǉў�(��9�9,z�U���To��(I���Fh֍�� �M�����T��s{؄�!޻4��>��U=;��;�cп�gu��	f3Ő��˵��JL�����q�ѲiZ:XlxVHYEB     400     170�"s��$�X��aoL�s��JڅҺ`�9J�����󞞵M�$����ހ Ά�SƔ�zv{V���_a�������ޛ��6��r�mq��*���>�d1��>���xe2+fL�
�"�pt�y�]n��dS���/5>^^��ˇn=t�F��ۈ��KsF2��*���!%���F\�/�H�B߫^�@��f�d���\�"�T#|>(��v�Ks�?�,/;�������^��{ǟ�4yz}�(G��-m��i�)��[DU?�u3�(��]|�t�@�ٔx/jxh�r��1{C�Y,���n���QU�Ūy��z�-��QԊ<���7S��I2�g~�nZ�1��s�q�z�XlxVHYEB     400     1e0��e �u�]S� ��
<���8���y���g�~�`D&�þ<�7}d?�	3��#_O'cTIB�V��<�ϛ��P������c��4��"B��o&�'���ǧ���Qm���	j~+j���p��%�/'r��el�{`�+xu��R���.�>Tχh���v���&^)Q�f|�N���4TVoPh��B7��}��,�p�ASҪ�_�N�n[�)jJY����"̱�h��F)���Q���l�4�A��6h'Z�d�y��ʑ��/�ڰ���á�:�dX�)�����2����ʣK �D�G�_PW�B�c3q_�l'[�@�\�=`���W�Q	O����������3%�d�%i+��C�wo8~����f��,T�Nɭ&0O�CL��C���Y����П�izΪS{�]��)oD�<�����:��K4V�g^B�V�FK-�����S	I"	&v�
��;���bTXlxVHYEB     400     1b0�����γ��Ê��kf~�'&�e�i�e�x/�Vmd�jGO�b��ZH��I�N[��i��/�:cHñ�ku��(p&1'�7����&�蛊0E��rNH��	�g�:�K�{��1�WK�ul�)�c'�vS�;��Q'��tK�m�O$�&�N)ٹ&�%�Q���-�YhI���B�	+$R����B��s�;�!A�]=�V�(0c�Oe�����t��$�VW��"8��m�@�R#Bnwr�<��CĪ�����g�;��N����,R��:F"O���� ҁ�����f%�f�Lm?�z���.x��q�G#�Ӝ�v�ZS�n��[3YYhV�X����D[a0M�Y�8�IqtV�6O����R��F���vd����"����tN��`����5�y+���t:�w����Ҿm٬���XlxVHYEB     400     160x.�&O����Nh��e=o߮ QFV�2�4]{X���6�s�ן�b:��f����%�3�ÕDJ�=�;|�&� o0�X�+�_����E���P˓���Bt��0���!��Q�G��U�+F�q�~k�d�wo�I�%���@�8Zp�9���I�cmh�
�����/�>�#�����qԶI�Xۑ_��M`�9�4�2y|@	�ؑ�-��T7%Eg�^��������s{*����W��P�EA��V��������	h�e���["�X8�,Y��������`kr�6�@ql����0=FWz�k�`dU��1\��Pu�@�y�goEM<B�A�K�=�QXlxVHYEB     400     150�Єd��]��x��@���Nּ��
�N,���r �H����3��fYtp1`��$�z�M���@��),�2#�sH&G����[��ÜW��R����������w�{к����qB�q�B![�H1��ߐ���%b)|P���\����K�No�m�WŦ���%�<W�Q0C�� ��%{C�9�(���M��L��
�{5ɠt%=Uj�c��B5�u�@D��x�R2agG�s؈w�+]�a�7#9����Q�����t�tinl�O;�O����ܣ���5�e�M�m�G[s��So)�˛Xj��:O�] -Y$)��XlxVHYEB     400     1a0��_�E��Z��1Zo�����=+P̦��ێhD��UOڬ�ɳ'GvW�Uk�2���� &�At�"K�(��~�+�dq����^�	(��:���uX��eq2�1c���d����z�����*�f}�K/��ph<��Z�����y�ő�`��F`~�B^y�5���Tb�\Ձ��bأ;�r�R
4��ݝ�w3[����猢@Ͽ���XF(�r�}�_��hg�����P�i�0�U��@6��0�'��I���>cm/�?%�x��A����L�R��#:��;u����]`5����C�E�}9���!Vz�=P�}t^9�ǉ@�"ۉU|��ݿ8ȅS���v�G��dܨ�NI�)�$��vR�P<��(/X�M�v|��OM����N�j4<li�LW���Q&�牪)��v�,��XlxVHYEB     400     150��
�hH�5Y˹I�q���x$b\li�!J�a�! �0,���-v�.�;���˔�#|����T��0�r�5��d*if�1��mʖ����s��57��Q���tP�|�*���<��&��)�ߗ�F�������a��ؽ��c��-�kMo�K$%�y'j��׵��%\����mǨ�v��7DA��FGL�o�j~�l�ŎR�ǅ&�1������ۉP}&����a�e���q�ꍟ�eٶ}��:ؽz�Yd��o��N�W�SL��؞ƶ��MwX5P�5���Κq����+���f9���E��#2���x2���9v_?֏.Z7`XlxVHYEB     400      e0����W9��ܻ�,BQ��Գ�6�`:�۲T�S�^ټ�����)��YFW�	Y���YK,�g�n:+�$U~�98�k4���:��ه�~pb}Y��z"D�|����ֿ��b�%����]$23b/j�����;� ���Hca���X
�Su>GBj(������o>U�;چ�!�S�X�n���$I%�SZ���;ᬃׄ�1$R�
ILd2iXlxVHYEB     400      e0����f!B f&sr3��a�T�~
{n���R:��{�D+�M����kԐt����EߘLC#�Kj�?-�>#5�Mé0�|�j�j6� ��C�k?/*���'#�B�<U�t��AMQ��M��-�̲k��Q���5nyL�9��M��(���H�] )��M8f�,���^f�f���0G��S1� 1ԋ��ƣ@�
t0�H��)߻Pw�  ,��4OD�w%����XlxVHYEB     400      f0�h�-�R�2Mma[?�$b`��%k��QQ(I@����/7?��b��u���Z���6�z5YqB;�q'އ��ٟMп���;��N�~;��$O�>����$��TB�U�4=�g�G�7d?:)р\P���!�RW��vjCt��̐*�74AЁ��˙9W�1�h}�޲Ej���=pK1 ������(�̵P<�\6,�-�˪�b�0jKKʟ�dj3�s�����XlxVHYEB     400      f0��N�C}�a���|�	?�@Ć�v�C����ߦQWM�G!�"���s�_�mU˷��/U����ǿQT�bgd�OC�߂'����(m{ �4�Oi�0�U_\�SM�
��}�����ݾ�(N�C7�:^F�}u۴ҁF�7+�9���d꼐j�<Y����q����=ui�ys(B����,����x��R�U�cH�ƗL�Z�u� kA$�FJ�����~/B���'�N�XlxVHYEB     400     110T1�F��M)٠GA(@�����<�?GQ"Ls$��-�^*��+���K�����g��Dn���o4��e��M���)��o�,��Sna���������TF��o��]y��TǮp�Z���\
C"���	��4j�|?\«��7�X�O��T�d�i��>�Q�X������AOd�r>�x���
�v������R�~��%����B�~3�]��O�9G#ӫkk� �0*[��UM��z�0g7oo��|O�>��H'z�Թ��]ȆXlxVHYEB     400     1b0����/�?=�E��D�
�Lx6���|Dl�n�n6��?F�9��e�0.�uk!c���o��o;p�0����C�JN�y2b�VƐ��{ۉ_/ %nM7�p~��)��`�x��X�Yq��YmI��z%�H��9T��ѐ8�EZr�S}�F���k$�a#����S�]-���V�	+��ԱP��Ǝ:6���"��{��fJ�]�ػ��ֺ���?b�q� ��N����!��2�����V�u.~�
`X~Y�
���Z�f/
��	r�7�&V8!�Q�<�'��X׽.�'7^Z�Ǩ���И�An�/PY�@�����A�5s��#Zt� �����{�
�<2%Ǵ����u���b6/{_����j���A�o�7�P��(VGƇ�;H�s]2�2�DZ�`xU�S��S-yXlxVHYEB     400     140#��X�B�GQ��Q��E�e�Տ�;�\
o�S��	����V�,��%�\BQ��qL,�xA�f�:7�8\"Ҧ��V�6�ۡہj�|ǡKn��7.����ޫu�\+<@�=7I^�����Q���#3�e�ϲ0����pM� �r������H��X�n:��M���H�ᮩ�԰�yh���w�
-c�'�b	NM^��Ȱ��V��^��a��)��?x;�>+�w�re�X�X�)��RV0�����n3~��+=���xd��J��=�3��Rc�0꾞����κB�d�1Z �I��pB��D�XlxVHYEB     400     160��
J�,��-���49 ��s��|��,_����&����q~�=�0A'��hŜqϏ����m�@E�6X�}�������h��g�E���4r��YHѤ�R�}�]�Pϫ����݋v���1�\���9x߫�]�d���(�ű��ޥ#�C,�n5@-�L�s�^��K�\�y��	ID�
X�J95N,����4���:�Y�?���zƌ�0W���U^������PB���%�mV�e������S���rAg�͙�)+�4|F���YT��4�p��ME��7J�~6��R�C�[�_5	�I�cͤQ��e�&����+�j�L1��� �轋 q��v?g���XlxVHYEB     400     140 �O����wo���w�Ĥ�q#�׉5H"4��]�j��/ɟ��G�7�<�KF*����	����9#�H�d�2�	�`��~)gQއ�#� X��	[�%��ӧ�7���dB�ÐM�>��o��i6��\��U�Ξ/��ZB8a Ġ�d(g\��,Q�2f�E��~QRw`����W�+lU�*M~����4��صS����m�/W>�Ҝ��	 `��ĕ0���y@���X@F*��!5��k�s���7�n�s=� ��3%g���Nk���N&g��K�t�����Ku췬:`����]��E���Y�]���nx˹`��XlxVHYEB     400     180�a֓��s����;���(\ ����=utl�ҕP�Н �� %��q�t�p��1���k5�Ɂs���K$��ŇFZ?)n�y��C,��U�:)t{���K���&X�V��З�c��)��ϲ�P���ͻX;oi�5�7�Q�K
0�g���[y��rY��d;��O`&6�_0�f\���0��)�\��������ɛE&Q��S��äk cw-\'�/�r���t������נh4k ����O{�;~ʷ��O�lk[勫�}�TZA�yQ�̔��_Xa
���'�4���Q�Ҭu7�%ģ�̝*�!�e������x��aHŽ��k���9$�T�sXD���!����U>P}�A0ܮ�3i��:XlxVHYEB     400     190���mH2�ܵp����j}�?����h�J ���L����B�]�Dk2�f"g�����SO�[#�7q��
H���`<��y�MA���t]S0��^�K𭘕�v�z�9l��Q��;h,�����4����*z�zf�=� ��K�z5��2�W���v��e:N�iz�o�^�Ġ����Oa�V�#�>HK�V�#��E�n}l�߿��VI�+B�5�(㱊�����ܡJq�	��Mw�Ny��_���lE�WV�^�����U��6 ,y�^fIH�v��"W�5��+�0L������t������_�26�``�pi�F��;葰}�I�Go��%�N�����ý;8QVDf���5[�Ⱥz����m����/,V���% �C��EK��$+��VXlxVHYEB     400     150|!.R=����8����\L���=(�f�������C��(e� 8p�T���2c����e�r�he�j��ئо�r<)��[Ry�vI�mk�rc'F�?�_~��ŧ�;�s�d�ȷ������92�P���:�pxgU)z�|�$��v���cqs4�2/P��<9��+�"z��{`n�]1�9�U�f��Jo�D?�k��|ߞ�b� ��J�cb�i�(�.'H��-þUs;�M�n�G��<n�Z*�?(�C��S�S�������/Wu֥T%BD0"«�x���i
�/�
��Tz�5���H=�4�F�_���	rm�����%��N�QLXlxVHYEB     400     1a0 �oS�����y-ϋ>�' ~" �*۩���
D��}GV������άi��;|�b��ض�Hup����(-؝R�~������2s�n������Η�o�L� �6�?���^������3

����䇖Q��dۄl *=#�#(s��w=1��m�pq�:=c�DN��x6>��������:?����%��-z9x�՗<[Rg�0����a�-0���/.>���1�Z��HU�v��X; ��n���@�S�:oUث���9i����=���l$�[�h����/���$����6�1�Huy�? �1	[skܨ�'�JOp�u�U]{�־.��f�3�O;Ra��w��X��5U��s(�����0  �N0�����|�<ʌM�U��ӆ�XlxVHYEB     400      f0��,��,T�]�ԚL΅��.��VJ�0���V��5���ƫ��6�ۆ��\ u#]u�2������Y��0~�f�����������<�R�Uf�Pq�1�ch91`�}T?<�7���M�}w?���Hz�DkDV��o^�Φo�"'e�g3^gG��a�c:7���Ū��<�L���"U�˭x�+]Wk~��-�o��<�G��լ2_q5!d��[�n2� �t�%�U��XlxVHYEB     400     100��P�_Wg�\�&�� ��FǺ�\TX������>�m^�m}2õ��&�lu�~�,>�}���:T,�j���Y�yp�r̳^b�� �pW;*����3��|�GwcA��p0���: �q7�k��!ȭ��j�a� ��ڦVQ���=���p�Z����CԔo�$%�C�D}9�x���Hl�Ћ���1�@,�.ٰ`O���'�}�y���?�pl�/g,�@�7,�T�3�\E���·��w�$� ��O�!/_[XlxVHYEB     400      f0�ڤ�΢��k�y�JZ`T��:T��F�t������=P����v
����J�]le9�ѻ�!��%t&�J(�ݿ� .M������#��?kWJ��d-z��jK�KJi��橣`�$�p��r�S�p�p(�c���@��}f��1�@�-Q�<�����|%@0�5�H�huG`�e<X�,%���y7�/�Ҥ=0���]'�C('F�1�E�ȟtm�GS�&On�XlxVHYEB     400     120 }֗�o��>��/$��w�]��0]����Hs�*��b���s�
]'Mq���|�H����W�x;�-j��S*u%��X+Vdy�(g�*�$���ɳ�7u2&TO=��!�/�P����+������j%��Ԅ@�}�>7��%ئ<�TԀ{!�x���L�*!�*T���=C�����w���:�,��X�ѧ,y4X�#�UFD�£���IQ�l��1�!B����?�'�4B�,�^�{頦03�{�ۖ�xqZħ)�@�/�[�{��d�/�@6���XlxVHYEB     400      c0٦��|��v]��5�k�j���7�H!	C�Yy��s��J�b$S�S�Tk?�kk(b	>O�4����P�ď%-l��f��ǌ���m�����aO��v��q3��i�R9ڕ֣O"��Л|����l\|y�,�=٦<|<�� �|��,�a^��݊\�Zt���r�W8Z{�(^*Ȱ���_`��PXlxVHYEB     400     150@��J$yʩ���]�̂Cv�pe�Uɖ(ݕM��p�}��ʘ��}\Ȱy4���U�R����`%�Gy�o��}�<jĜ��ͯK�@�|�p0P��/y�$W̧�&�	g
�*�Q6NK�m�8p�zEX�@�D�����Jf�ҹ��YNb����԰=��'X���
���Y�Y���L�DQ2�i��bt$�� ��֣ڿ�q��`ʹ6m93X���������n{tR������毯#9�����O���7�&�w�o���T��6�t���}R� ��H3~�Mkc�Ԧ6�U8���_�+�T������Q�d��0ũ�A��5Ar�XlxVHYEB     400     130�7 F�pH{����ʊӎ�1���"��ɼ`���#�L�C4����;aS������l��b�!�vqr�������o!I3�c�����1A��d�X�ބܶa�>�b�űB���k���᲎� (�8k=������M����������m �G�PqF��-�ߜ=�.�щ�pJ����(>঑҅C��?��y���	\����A/ϟbA�ي�A`r���=A�<�K1�=���r�K(+�I�]z�����������"S��l�:�l���/�q捋i9~͘b��o*=`ŀ_E�OW�O�}L~O�QXlxVHYEB     353     160+��k�)Jb�V�F0�*��tH�q���)�sW"� �=p���x��X�B1��'*j��Hp݊ �[��ă�U���@13����R.�|ؠ<�t���G����ǈ��Qƈ��|��pN�WR����wHpIr��\��1c��.�9�.c��aOzz����v��c�V-���=?�pR�3��#/�ב�#f������>��N3��2dr������zҖ��yx�F�4���*SZ�Ǒl�{�>�5��_},o�A�7?�wh�F��뭣X�S��l�V��=�F�Y���2	���/����Z�T��'��wU0�j>�wg�
��Զ-��[�KEU<�