XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���=���=�9Df��TW�b��HU��`���#D�j���M42�d����j&�X��x�A:�j��1����1��>�B܁@{cFH�B�K�∎�<��AT�����H�|DRfdJ���4�&��-�g��z���gט��o�F���S"��@��5:�F���鉋
��q���ʤ�U��\3�+���X���m�^���F��5�z�"�)ўs����ƟK����L|"���ad:z��93�{�t5@9y?���WbD�E�m]�qK	r�� �~��?R��f�����B�q�M���oaL."qQ���d����:�oES-�0��-�1:Mg�ƒ�k9_�\�VяsXJ�B+H�Ҙ̀V��m��e���_�����7`���]>C+>Gλ�8������4&yV1�;m|�Ֆg��0e���ָ;%?3�m$�	𸬡8���Rq���j��75���J8:�l��t�l����<A��&��<`�imG�ja��x�+Z�9��i��7f���u�[[�<	��L��~��3X��쐭�v4k���Y}}(�����_�%����)ԭ}�P����_0�f~I�6E���>;�o��=�^92O��=N��r�����Fi/����3��[�"ˡ4�Ҷ
��8�
2� �ٗ�u����
�a�����ֿ��dK&��!ӹ��1�S�W,�k%�\B��x���ǣ�ŀ\��mk9��>�FgʒO\��Q�;S�\����K��,���i�lI����XlxVHYEB     400     1d0��z�6_QT��U�$��*-���G�;�Z@A ���˾H��W�%�~�V��W��A�o2�'���i:���T����­�+����$W�z��+��Ku�[s�C9��*��!1�S5���#Y�ϻ=5^
k��W�4�a`�XJ(����� Q�?&k���l��(��Ў_��ZRI�EՎ�hm7�Q��kjb�p�d1��ݺ�b�m*
�c��u�˪���LlA.�Ng7e;���u�1Oc�>0��8Y!V+v%�����8.�sF�`Aa�RIw��q�e[%*W�n&E/��4�3�$�=tD)�Ku��/N�<L��G���O&���
��
h��ur����i�8��<���P�ub\k[���=�UNu�.w�9 �|^�9H�H�*��9a0�XDyr困�5�e��/���[������b�����k�t����<S[�TOv��XlxVHYEB     400     180C��(�"�24��]!���)��q�
�hn�8"1��4-�v	�S����>e�D�tHE/^����X����!C�5���r�QIq>cl���Gww�~bE��3|Pw ��b���F���~̈_4ݢ��8a?%�XE��%4H�Uif����Ąh��f����2|׎��Y��q?�MM�i��BXV3(K�!=%���m>�:Q;g�=N�\�+cȞ�4^��\{��/�y�̾��@�DGw�Djʘ=�U <�'NG4���f�9���vg����w�q��g[E��vBL�q��Y����M�tW5l����]ǟu��K��F�ԭ�/Gc|���|�S~xB"F>��7��KSg�􀤡ˇ�8�|h�I��[9XlxVHYEB     400     140/����Zfq��cg��t�.n)q6@�[�"�F����������3kx�Q��Ӗ����f:8ghp>��%�������y��ۜ��$��ԨMʕL��i�:��m�^(E�~疡9��ٱD`�>x:k���D6��<�p~�l{�(�	��o.��ϸ3~�	r�g�1��S���*��sp���� ����'�,2��s���op�~�r�	��IC��@Z`DQ���՜j?��� 져/���1�?�S���n0�e2&_`l���_�``�<q!�5�ޘN&h]���JU�D�`�k��]���*���ȥ!?��c��XlxVHYEB     400     110dF�U��Tdy9�Ћ�@�����A7���X)����*";o?��������d^d�,���Y[�؅�>�"O�d��t�3������}�Z�F҅jǻ��kȕ}=��T�<�@3�(%��r�����֙�gR�v���{�!M��7����m�v��u�T���R�CC>����pY �� ՛f�JկH���g�y��C]�Ek_��%qE%l��1n%���C&Fp�>l��"Drk�u��S�=H��� ��!<&��rdXlxVHYEB     400     130E�G���{��'�*(*�'�'5���--W�524�<Al�@��p����ɬwwD�����}�J�Z�� �9����
�޵ۑn�a붺�l,�g�}O���BDR�*ɖq�49��\�"2,��Y~�O�H
@�v�z^��׋c5�,@�� ?�1_�2w����H-��o�7{w�ԇ��̍ϼ#M�l�G��훰u�;��q?�����9��*p�N��(Kx�{�?N8]�	���T	u�Ӆ81�IEʅ�O���Ι�B7'��+MpQ��cP@K�W(�K�f=��q/@XXlxVHYEB     400     150�V�`1M�<n���Ÿv�+$���X�?Y��Q�F��s�=�֋�X�!ۂi_R�Q�bt�!����
��J�i��EĀ�����.N3���\�G�����ܶ�.����E�L4�m2���rv�<��!t����(�Q�np���b1�rB����"��my��
+%��PƆ�����\=���E�!��\?н#*�b��ג	�M(r�(R����J^lI( JBabb�V���때f:��Mb*?
!/�EPj"�J������%�1���'�Cb;Taz�����W �L��xq�K���׎W��'�����|�_���p(t�jg7�ǒXlxVHYEB     400     100<a���$���n{P�R%ȈN��c��X,H�U���f�3�W� 26���'�*�\i�?��Œ[F�c�Wp%������[\`7r� �ٿ�)�(_�y���m�ݚ�{ƭ$K$�۔�܇m�6����9�yā�Z��[���k����N
)�e�~{��:�m�h���Y4k�+v�2���`��̰�h��?eL2���8nT�2�Յ=�g�eI=p�fҩ5���.`����;ɓ=��H���9��MXlxVHYEB     400     1c0���V��������FW�j-�����+hcޤ��$���2#糪�1�ݷ ��$��*s)�������ÌO������Fth��F(i�Ie���s��)�>K�ܺ|df�tى%u3h����r`o9VӠ�C���6_���V]�i�)�=�ǭS�Ѡ��6�����̛VD�����P��jD�Sf�u1��T41X�}5�h��*��J���fi|�IfADӖ��?���	��������n&�cuz���bdk�4A����ۙI�����haj���`��9lbII$`X�-,$�ݶܲ�sxZ��Y K�,8�cXG�û-!#�CK�wg��x}��q�Tl����� ���k8C�k_�N�i����$)��"*����X˼�=P�X�V�=�����`��C�� 7NypA>��H{\gϴ���	GqwC���QQ%�XlxVHYEB     400     140�#g��#�>*ڕi����~�"��T�dh��7kßZ&"��4MH���'
�7���_��: �gp��b���?9���F�yݲ�:T��L];:��a]�J�詸���f�e��$�l��ã�$�&w	������k��>��ul��j�=@L�@h�� �qO.Oi�l�Ζ.EH�ڵ���m�ی�(i�Y��\�fZ�U�R3�{����j���p\�wGgd�{e�q��t�E�Bō.�!�4λ����7�c���lyH����/�@��x/~ס<�9C�I�l19;��M~���!��d�](���,�XlxVHYEB     400     1a0n�V�F�	�kJｪ�Α&�kHZl��[���̏&���S�Ŋg��G��*/6��i��R�������������������;�t�J{���l�0'�D�Us���O������'��6�N���oF�Ac��d���I��(����M�\T��)�D��uP<�p7�e.�����"�pIX�����>���M�!N[�Z�6�b4#��meïV�Uv��r��ߘ��#�o��bKk�ڏ~
i,n x�ܭ�f��C�Cby
4?j�2�0.�����ͅ�b��D���7�M(~�M�6�C�O���48E�����2MUv�ّ��*f�ș�?�
p�lXF��8i�Έ=ߵ�Cbˈ�i9C�	L�!����,U1|�����X*�n�Tg�/џ��|�=N�D%'XlxVHYEB     400     190{����n��j�[:�K�<j覟P�郮l����Ɛ��.���Ֆ��|_�='��Ǌ	"�[Z|�)l��?Q�����f�2� �U	\�U������}1_5((5��H�'yQ�OC�"�5�
	��:��Ot��?�6����4(>!���D-^� �)����*�_��͚��h����Y�Wk�Â��TU<�N��S����r���6&7��������|�a;i\����ň,Yk�;Uu)j��g��%��~8s����k�:r�.n�:�XXu�+%������m�1���'U��,����n���_̙H�jz�.����(�����mJN�lk����Z�]n͌�g� �n<�j�*��{��d3�����F���.�:�Q�\�9�鰯�XlxVHYEB     400     1f0�x���D�6X|و`��I�ߎ�l���kO�?��4�7?�ӄ�v�<�����N�����\
\�[�-��M*P���:\L(��.�P�l4��p4�� ��K��l8�l�<g�!�<�<��I`�8��0x���4�oGέ6���ٓ�c.�����,����q��O@Z2O� ����<*��U���f%���w���컷Ɇ��QK�� 8?��	��_�����]���Ө>��4�XS�\�&��/vO�+Vj8^)�@0Z�^�)f0u&W��]���r��wDj}T/k��%�9���3�.)��4�S��͏��g��T�����X'�M=p��m�!�`�u���@�:�*�gu�(u·_Z;l��\��m��^�i�-){a�*uE�����}���ڰ�N楙����(dЩ
�f��/�lc���Jl�N�ә�6����;�bcg�����<�#��K6��;�8��[XlxVHYEB     400     170���T��Ě�ie*�é���P9 \b���A�+��|�q˟`-p����5�D��F�R):�_�?[�!^X%{n|;��,��@A���g�(�x���4��˅#)�Q�դX��:��~�Dg�.s\�Dc�Đ SO�\|�@��<��g9��$��}�1
�8}!�Wǡ`��ztb��ۖF.E��^C�h�r&��<�K�in�\�$Ү�Z�i��!A�R��_� }'ħd��g�A&8���B����g	�Jc�~�����Z�2��[���w9H�X�x'u}�+���Y[c'�=u�,��Zk�Q��3&D0����4&�L=��h��L����T_��Msw�Z�R�Ao��XlxVHYEB     400     190�.���k���ۨ*w��Rr�+���*�3D:1Ug�c0U�2'��+�$���h��8���I}�;�;���e`<g>[z�D��3��Ё�bDp���E���O�|f���L ���X��;ԗǠ�	�ξZ����F�=�Į2�c,�����f��@b�`�"���{D/�b� �9!bQ$����~O$RD���0��:���5��2����x��}k���j�9��l ���w۩{k�]UD������75 U�zZ�e�M0�_k�4��K5T�F�΁k]���?*��1%�H:������5<�ڀ��6���kî��� �q��q����k$a��Z�Y�+5�bw.!�X0�4��O��5��Z��i�I\�l�,�>�(��E>�C��-Е1XlxVHYEB     1fc      d0�H���o<t�+�|}�Z�}�6{��nP�����-# �aOO��x|W�rS��D�%䶶�3/��y���Z��� �������y��s����`�7����+
�Y	TZd¯`n��L�PO��F�&�Ȃ������|��Rү�*���L�/���y���/=m��`C[I���$��������^��X8�f�s