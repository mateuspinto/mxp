XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��u7A�7�ה��˺*]��ޗ�N�G�2�7_�p�fZ:`���lP�;�ҥ�0�ၱ��D�$�4�z�d�ؕ�3G#�A�
2+ �*M}кi��?�*<4��O�Tb7o�wD=��Z<v֙B��M�ʈK�v�pa�>C��3f�򆯉����J���=����pY�UE�&_%���n#��N��G瘐P��k����ځ�G�4�����c)��:
�C���3J���d��2*��ι�`腼��q��">���w��2)�c���nƔA^�e`��j�0�/3/�p	8b?��*Rb����c�mXk2��h�`�7_�RL@�����yE����}]%�Op�U�G�Z i�>Ǥ1�K$�E>��K�<Һ�
��s��E�%�AՀ��ǳD�K�;QOK_��[z���ՙ[ �T�kD9=�D�m���Z�J���<:���k���������ө��,?���g�S�:rp�{"c�N��М���
yr� Bz'��*���	�\�N���0 ÕCc��K+���O�i��	RDL ��ҏ�#k�L��}��S�zӷx���p�z(H4Q��[�Z\$Wrd�)�Z��=�I,�#��M�.��"�r� .C�W�%uG2S�n�]u��� ��u��@(5-Ql�34ע��@��5�/���_cN����� �y+�oJH� �L�����|�{}>E��!h�y����4<ܳ=yO�����߻{�0ݍ�1�Q�����m>��tg��I�����wx�����镥��)��ڲ\XlxVHYEB     400     1f0��[w}ͧT�����O>[v�w=���9mO����+�����b�G�����=~���D��X�� Y�'�+���>�:Č�T�U����m"F;)Ф��Gx�6�X����w�PЋ����������=��"�1
�"��% "U�����ZB^�j��~��V��oAK���:EdK�n����F>��>{��/�Dd�%n1A��x���X;�g��,!YygIf�K����c�����qL/cd�j'�Z^�E�9�j^��*�co�F �s��I��o�J�|l���� �&���E<��6�Y�0Ӹ8�g^>㓶W�k���K	�v��k6�ϩM	z��0j��Aw��X�$Ø�| Ρ����fC�(C��cXL�	����?���?�l���I@f���45�$�K^��&�t ��"puPѷ�w#���eo�ќ����� ��_��ɔFL�p_V�	x��59!�0XlxVHYEB     400     130L"�Ի����8��G��&�/A�
P��q����
g{4ey7d(`���PpH��ȗ�< �ͨg�S�`�&lW�CF�$/}�G���:� C��h�a4W���כ�ff(�K��,хl%"�(����߹d%��ɉ9Qv!�S�!b�SԉfiNB�C-!1\�(|CQI@�k��L���>�w���ͽ��@���I����{j%*���CQ����4��ס�W�(j���V��F&��U���W��ĢD���3��Z[�nf~�. U1�\�f�x	h�C�X�2A�m1u�'��E�mYǹ��JXlxVHYEB     400     120~[�{�剬%�rj�z��87�퇌>U����.fGF�}���_�AfO�pj\Ţ(�{�VMENL�J9�;�$ό�)�"��Do�� R�N� Dl��� u�3��-G�v��mGӠر���9Y��s���%%mwT���Q�����#vۥ �s�ZR2�]�رX�֨��y1�V�8�w�H��y5��hhV�8F���4h�]�?�ļ䀺��{�"F��J���M�rm�q�����ZM������v���Q*Q��cJe"�a��F(T���b���}Y_�>xH"g��XlxVHYEB     400     1304�2�YjV��'����X�nXX:��u��O���"�3�b��f8���lj2'T	"	Y��Y�R �	�٪⏡U�_8q���e�6<�\��J�A�aa&ڵNIax�DB��M[���IZqh�{%#���Bel�@S���}�����u�x���eR� m�((=&��$4 ��*�h
���7@x���(~BS�)d��,� ��7y��ׅ�����\
j*T<)tԜXX���
���g����93��r�]�XS\"o �#�Xi��|{J�:���K�s�84�L��x��wr�F�aX�eXlxVHYEB     400     140��o�L̬���/:),[z�&*�x�AD'.����Hԏ�%_��{�'2zH�|�z0�jI��"�2�Š��4�f(|�����L�	O##��D���U�E�\3�D~�n��M3��ܣ���s��^���vʃTN�~�����B6�4T˥�b�m��f�����$ݢ� ��Y=��rWFmK%��zS�:�
n����Q(�1]f��� �d��	�_�j�C�R9��TLw JS��*���ݭ���ewCډ��
���➶�Ŷ}�_s6$��pZf����Q��[��/QK��
(�}�<�.��#(�2���g�^�� �XlxVHYEB     400     180��K�j'0v�`Y�0H��k�`Pl\X(���ʬ�����B�&p���秱xq��S>��P��Ղ"�)$u;�a|���ix�K�6�~��_9`�̷��?�;��e���50����b�+�M��x��@��M)7�w���@џ�mæ7��H��3Ψ9�^�"_�=�>�.� l���P�!��L�$�?s�ͭ�T�QL�-�HOu_"�`<��\: ?�;�c��փ�-d�>�z�58|EG�+ʢ�p��9������!��!\��qV���S���\�Z�Y]���p_}�`t�N�I&��r9�e�c�,L���:�&R%�/0�#��!��h�b�wbV>6`��EK Ea�����5��`H�EVY&:1XlxVHYEB     400      f0n��~s���8���1־��0�j�ۇ37^�^;�����?���1z���B>Q �Ͱϸ����f�nƶ�O=�M������qW�L��@$JzTVp�D�n���A�Cj=�Sv�<�H.�-:#��؍�4�=����;Z&�n�Ʃ���>r��dǒ����`��Κ�X����?�a���/Kl����aL���G�ܯp��Ya��������8čet�P��^�H�,��5L��CXlxVHYEB     400     150q��u<(!g�t_$_{-ɪv�����CY.HSג壆�O�dVd]��tHz�	��o~��S1z�E��/��%�k��V�:Xg�g��y�z���2�(A��� ǚ՗R������\��%ܟ(�\.���N�#ޠJK=B��0��E)��c�*��t�J�>���E*��u�L�&�ݸZ�	����7T놏_�m	�r	�c;-�sL�Qy�
x�@z��m�����zu�f�㞔��ԛӛ�t���,��:�a%UnёH�h�	�{�鋴��s�V�))S�Ep��.,Pp�$���|R㞽X�5t�-a���� T%XlxVHYEB      b5      70'!�����Ջ���λ�v���G�|v�A�j7ˎ��U�w~�S���/K�ɣ�g���3R�l�%�o�N����	�Ҙ�I�]�S��'�Ro��QqJ�G�b��6�=��2��$#