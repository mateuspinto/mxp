`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
IeKsF4B1WxwZlSYR/P6oaJdFSQoNihrnnI4R0o9Pl42IEcgjOOEP24CwsZr8UzJbtiNue2YRjQw1
sLoxp3O4N8vpxTVNeGkhBdLW6yhi2C/A+sFunyRtFTgS9LBpD55MINIXFbARvBJS6xoS+gDoxbKt
mWcxlQHjJMpg5eEozEirRufRQQep2HEh6EqOvITdTCucD9EpERG5CUG4zOiyk5QisP8rdeOtRArE
/YAEwYOmqYuLkyvCXmoagYejfzh+tmYXcaB9eZkTltICqveHET1GyLyikPP/gm54nixOQZoLRym5
QW8SqXEyQzrrut6qYq5Hfr/m5agQyO5UIPL+SQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="oGHAcwPPvNmcIabONr/eEJemzCAEvwte1K7egdUOyVc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
NTDaaA2fxk0HqG18DJRiEPl7sN04KcH+R/XcaGtPHPvcwzuHGbOJX82MC742BXa5Shey707VBYfD
7sqOHTuBS4APMa8o/34nCW+KzZcXvPDEw2e/bhEC6mnxL22V3v8mTZBzcAt+t1X9esTlqNgz4eZL
936yh10zekmdgIOfZNACN2E3D6PASwohPqd+3g7beahAUpsF1d27n6g7zKvxV8HG/cHWghcxcHVc
sDT5fr7xN3gUGyzRziilsz2qo9uYRLWmF4t5QRoFqDhWrX8GKx0nUvZEtxXPw1g8WRPt2uo+bWpY
d6o4IYlRQ21HBQY4o1NyETzT/iISHcPpCNopON4HF0A9UKvtKXFsbxef3TqeaURbf88dNUdEjkJ+
YquJtLjxkpszh8Dfx4ZG0Uvg8Bu/HP5htVRLZasdfX7Q8ZH5SNdVJS19Z2DPaquJhHHC635dsl06
OLv/H0BoHPWZgZpzTI2E2l0rjOE4ePasWoQNS9wWW4ecM62gEOsLtxhqsOpMOF0F09EdssRQnROK
yXOkO/9mA4BF4STPSOBPLKIH53i0osICHcWQi45UfQ3Ge14H6cTygHGAlBe81kWTybsjdZcY2emT
2hPmCn0co/QObozTTNBCJI80N7e12bVcJXiJcKLa9f45tgVzpJM78pV6zlCRaK9a5OU6sjm8OLVv
NF2nRKNSqiV1NaQImPrdK43ezPz0f0SXex4f5e+wpzErmTz4d3Cn+e73C4dSHPxsfsSoc6YkBFx7
+8nNBMHt7NCeTDiOxbtUBmr0N3QrNrVHr+LOyW1B518JFHNeiQew0HncqpFW171OwEVChVXhAmVQ
8AST/3uJSHRTPVkNiwm8uUIi+s7ONWH4q5k7nnnFtuQjmwdqMFfjropDzyN8AVLqtviLZu37Hm7+
TKajT7Tu47OmkWrMyxlsGIRIsOomVeaA5uBoSvwuagq/OvmhTHZIncwceJf0jHCVlEDSIIWFDEbd
3xrVzG4VW4O9dZpcJEqgaF5l3Gl9RkrkKfH2ybk4jYWW2R6keT3Ex8H3iw2ZxjFCBSfOdi1/HMHs
+sFIZk9ETfzmpwnmfCZjL1vIovkxDFOESivZzQ93ajYvVHjo9Ld7WaLb6fXJKX2Ps8YIgkzs/eH+
gaWT38+qtCS5BHFPqw5vr+re9jD66SNufJvvFqDGSbsqP9NW/I6ja3mKHRJLNFkigF595P9BNle4
/BcigChuuq3stwgxuw+hOzFk5f86nOy7K92xsoxoNH0N4YARSXggkVuOI7rGRwaMKbp2z6DjMB1W
s+S/SprtYFvwOKagI8ZlbHlo1e5jmMjL6N04TXZ0p9qSBz4ZYnQF7XNGF9h1b5FHMwvdsC7byasS
boCV848LncTqX3tJfGkYiO8kRjZLE31bFROkkzGlCp1JS6wW2iSe9YXpemLwaICYe2TcWc6Jiqq3
CkqTrvIx22OBREBA0W3ZJ/AXIkkrJmOnK3JhyVdjDJBPQvngG1ZguYgWeDwSucje7XlkweDKF/2b
myfO+mU1mSC3OYx9KLMnHxgh/ppVNNKum/mg+cUs9pw5OsYTCsmgxOakUOlwhVDYcQWqAyaRxbtS
0mM5um1Hx6dY2rVxE09uvksd9WICmJibhKXB5Sc/Yc0Of7PA96CfwTEUTGbx/JL8irhmGAsUga3w
dmeFOA3cgZ2IGhbeVJiAqd6EnK0KxCWGfDu6wQaod5V8r7wAOdE5iJdXBh2WqXaP4jcde+h9WUlE
OCjoWsfxtzHGwJtkgG6uAID2kf1ubvZaCjcejWpmU2gubFR8Cj1kCY4bQNCT5kBHcuPy1RNijE5m
nNCWKsMdxsypg8scuIEuPOcN4u2OfoRlprlKbbvIlKBoQou34mWsVe2RBLbBvLL7y8yRJHFq1yWA
J2qMp3q+aLfDUHhT6zHbAOMxjsI4yI0si/kJz2lRokTmoETEY01A7whu5PKbudI1feN5F7SHqej1
ji/z16aph8MaoUVm750vtUxlp/GA+6SX8v5uHB7qRN5VImmL3UFRDE81eRN8xd/jvk1EsUS3Otiv
xfcHU4Off3xU8xVIqwdLlTBKADZD1uKHQJrSkGlFkgcCD9Nm+s+O294T0qncS6D+tRyb6nUqU7Zu
ojGOKo9+t0a2q2QFHFIrlJT8iZI5AxR/H3QyFkXgjF6EwD0XcJ9A7PXcKKs1GKJYJJBqFUzpr8a1
gU5xdjlpsMwNPi0M8WhGzXHLG4bEVqsbvp06ht3wrznSBSnI5C0BseC55TwmMpJPhsbCvR7tb7n/
T7gk48fU8A4G1UlWEIuiiB3GHZb3jVNpq1p9sOJ2vGt3FLMfV00t9RhQs95D5vxnAnlluKtUHzf0
QkMLpX98EGM8xDTtF/Mll63mx09z2Pv5fg8d7DVL+bTK4yhZR2c3QrvqhMsur15dKWQqiTGWR8Bn
KWfyA/kkbvcl12Z8SYdwyQIK++LLNan8RKK5fzUftav/YNLiaInbQ2t/WfLT8ao07gE5d6n5ewvP
VUUx8lSdgOC3/5dCxnTmRELwQieLyWVJOm7zHp9pzhA/+g24zf2mwNvtEB56E/nuxaNmX4lH9YPD
SsTsYGKcZPWB3B4hP6QTBDXiYrV+lJT12aA4R80y6ID1laq2xVzUAqqElaQdRGoTAROg9b4ebrDM
ac2NDhN40fG4fBzh8ozkT343K49KznxMv38TM7OPv84COueXNpaQurYKaNJXEoWrX2uK56s237Bx
nq4u7nrAcPgudFp1cjkY98xmSuFT9KEYEw2S1Qh0bcrugTWUiUeQzChuxW5i77ku03D4rju4G8Eg
oi/OkBndHQMoKYtCOVsWO1PVz87njn+rCBmzgBfBTdXbaf7GIFZn6XmT+zfFzY1PKbNFdWsMo9N+
o00zLi93a1uu0mY/eKraHwxtkOD9y1x80BaaboD0WQ6ctbfeOwp/7JjKQ9dt01ZyxkQAREaz8PhD
pGWgFdPK8oA3VjjCQMVgWGpzl9vMPhnc0ElGBNF/+KkDidTB4wqKjY+6t+Kc1HGdur08LS1gBveb
ViVBGjapNo7Z5eEjux5eQGjN77UeT9LKB//2034XE8KGqNUCmLBKYTlJjymsGbmmq+q8grpy5GJf
5a7OQYiL7WkLqh+j1hD2ylyfesaNRcplfPrZI11Ulcghls4wUTnKWNtHGTPNtNIsw4sPv8qFy6WO
Fk9nkK0FdkmuU+gkWjljSfEP52Ck2JO31N1M2BksRCzfjqV/DJR3YU/bDAI35eA1WCfpzG+ZvoQ1
SNEA4/Zq78DH3C4TlLJpYaJfCxA9ADL2dH1eD4TR8cgHZllA40NeF/FAME7kbXQWC17Oe1PNfiX3
V8wMxB5DTzjB3Os490q+DJ0WVInWWEQc2DRxsTkma3LDiiPkn7I3NDJGKndUiTVSP35hAFSF5eJ8
bMbXEIbf4/QZumrR6hblXuc9iYCkg+glK9ZfyNUvFzlxJ34EBHmw/gidSJi7miOrvMkEKv6u0PY8
mkh8Hxo7Qghmv/Rtnd/2PKFVFm1Te2xxoJFBwgnTrdi1vRKmnhECO4jIVsYEliJiK98lq+rALQxq
qeORKF8zVSsNv4X1QaausnmR14LIYz+ffFazB7mr3JGKMHl1s7MkVRHvZm+1ZK9YoK9TirCBjuWi
vvdDvjyg2L2BDa+cSsGWXV5p8qe1geEMAC4ReduYLL/lRmjWJ8hOzYyRnyItMofT7Qkx+fD7qGZv
uE4UvFO+QzR3g9c+k174sVWALwHbfRAxPKQDnPd4txMCwM7JKxzCDzOQ16pfxudwMKfQfAXppZtY
U5kAtOFGKMywkRn4VMP0fcZ5PPPFKLzcScnI+kix7inpuHUC2z4f0++/VplkasQeIDdcFAeZ7TFT
m7icdNpSymgd/k4fL/rgqRfgvQr/5ZKfe7LUzkl21v/qy6n1X8SH6Tn8bW/Hk+K9gh+Inerep6ky
o9dAdCr2UkCMc+hGF44uehW1E2MYK83g+vYR40zNd2CuBODB0u3wlao3l2v6hp0HmuOCP+yU7gSi
DnIKknJTZv+VdnsG2EHB181ONW04Q8RrsPFB+UCasT+3in1MHhVlt1UKwzb8D3NzOyZnLpeWgqEU
VNAgrlMQsJGeB5UYV3gM7fs/R0DgnGAceZECuflXWw9wIU+sKulrytrLfAEFp2nwUXZBCytOTkl+
B9l74THzhrAbMSmNYQkq71QezSgihYUrYImDOPE41gyyOypw6t8y1gs5YFgmaI4w2OwmTp15Nmlj
zj95wjnBEKJ1wdzJkgz7v4fj4yTjlWZQDRuzCncQCBmNVAtOR5lfcCYYLdOvSlpjprZmvgJ/QNak
g4lZqVqQ/fGvLXk/RhlZByR5CT/7hhH3cS7T26Pmb5f6DgHRwXJpI9TvRAo3gFVRNPoadUwVal7t
adeOoTL1YZf1V4WsCmL2Tb5fJvHVMJbsHbah6mXOC4KFNvyv619e+tzRkMcqI0CMft5fTFEEHvBq
A9eSL7U3MsthG0aaHMFSujoxPO0o8LNnlR0tETjfx5yFe+icA040nQUV8zES/x302T6TE6HI8pJE
UvVvtvVhSU5bO2mN8WIw/whE85sPQDTMdoZLfZ1EZsNDFWAWlC+tnVGEGcxTuuyh0SS5wUPR6fSu
VQOIFi7MXBZwMi5XOFPtcvXRylgUtmvYopyIHwu1JTLukvUFNHiCT2oDlET5+X58nwKNxsHm3EAj
cfsCb4jFH2Jqm3JdAyNKqG/Hf+T/VLGfL1dkjkelztA5rOgJuu7hwGNKZNCRdmNmDhRlbfn3Viwg
5MlPfkau58+af+50+hy7Ld1SM4tO398rMtC+YzQU70mXINMvGQo5u00Fsl5B0prx48CjGnlTQS5S
sI1hP/eWvTBTnealgCyeTEaCq2aihKey12x08TradMX8uf56O/YI/wRYrFLg9CHHealF7Umk/uCV
9aomUDSDm0Qwmv31LX7ngEsDV/5UHUCAG9jWOfuxLOjq8rP6CbfrSWQW79cbbI37qk2lLCiTvwgR
6y4SJifR06MrMkkN96+s7WZa6S1k9gFuoqnf80jB05CDNg4ZcfC6PCeQ4rezb/KQc4KA6oRGqAQo
oY7gATEjEe149JIQ0VAXMdtgV5uHA7Zzlg+TR3lKdCL1FZx/H0gTcDHQnyVDyvSel3/eKBCKAv0o
YZ9B8v7Om2MWVKucmYcbjl4qt/QbAgkYVP3DDg4KLNzdRw2azAYkFmwS/0LT6yxzflu5XyZ8aXEX
UPJcqqMQN9KGEeeCxnN7CaxNk9LZiBr33h4F2diDfPBdZixuLNjzBivE5RuseKr7F254TDruNaOj
T93D2F+YtCgYSS0iJvGH3yjaIyUwSzuoeVN3zzjB2ew8g3CcSZSR0oPJ9cFdYIfZcXPOclvBl0Ve
PM06ILYK0WhROk106BvzCqRFNasCzz1H2JZPKFKigjHqxRTnRygKvJG4B+rBf5S/HYtuH5oJzmPI
BYlKk6SoPdzWxS7Yiw0vx/pnbby2yq6SH5jGszjHkx7AtJBfcoE8MRGtYN6nbcAQC/96GRVNbaZq
4Qq3ilcRSfLrpNhUFdb9BP/Tmht+Uh4GS8n8Qj9OO+vo924QhBM7/gezj4OCHMG7p3ErcBnTjabw
6Ublnaa6OFxcj/07tVFuMgyFqTz1cbXp6BpiuQ2Z1Nh7AY9hbFlRlwQ3RFLaJiV3ah+ACwp9TZtH
Kyl2L02MpXSv86KhVUA1w3wBXIFY+1Hw+K36PKDlkl4DrzCRvB2FP3ge+D7nrae5JpU+M40wdaFT
KWpjdFbMBeN7bOxWhLxAH9+gCYuoPzbw66e5XuL61RGaw0CVZ3pKVO+XL1mo9+ik8ZtVoOubZIHk
rkPnQpobza1elkYeyreZKWnj2MxLOXEWUuLKetlfgMjTKS3XVCbPgytahbkO+DfwMRrzAWdE9G7Y
YmqCyYo52d/cAltD/5kGSkMVlXGgAjNLMG60qe7Hc4EElHzd3feleypCUDosPoR6Z2OxEVjCb+bd
N0PYqbw0jXpMF5Va/BuBGNPl+lecYHy74Va2DXXMyedP6ifcUnFolcYBRgGcbnbuLrp3bKMdX5aT
LKAIGprJ+7KEUURjDPF0Q4r49g1KvOS+qphHylbiHveOT6OAll34o9p3DOH5jTz+c2ylPm4YKZI8
qwRiA8Ssd0ELeMz3NbntCEeeSGW7tNxaB+Ud7qEpIu0V148rjZPKgPLJU5MuoBOyx/wZG3G8NKH1
73MpiGQXJHqvvLuLePuiFOGYZ9kQTHJjvdaqh837jZNOYqdB9Hl8FVIiv7oS0BSjHnfLOdsuwKZk
O+vWUFrrtdB+kgfv1i4yDV7JgFQ6g37CvdbKxjginZxPRxWsxSRUF8mcImWuHIN3Vb07XBubAo1x
4tH+00j6AWj5re9o8snCmqDzRFXtugPKBX4q3e+5xVAXJCAQ4eOoiD6B6MWyIw4GbybO/dzvLRHY
sTG+i0t+seWPRt0xclPb9JiQaCPcPmhd/NjOl1GCCRdnsx5vMwuOiOiATDMSa+xgg8YFUcP3LC1p
avKWHLRJBOLmzUAEuthuE4U6e1E/9QpaZA9OlL2/hEzC3xptPUSdCh8hacNnMPIoTUZA7iKECB8R
wYvYK/Q/4KZ0vgOhKWTxQN+SJhlbAZ6R871BgsYY0VzJbqSoBiXIXE1QkieH5aXT+2iqQ4ATYewZ
bgaVgNeyQQ9WDNuUmRJzy+uIM+lqaw+XeJnOmfG+DtPoHWYMZSy1qrewTmXpaU8rw97zth/aNIgc
W+uwJ3JjAPU9a28k1jRVWjidwrQFhSvdE1QgeztLosBlytWAG/8N8nw7IV0DSPSK+PtgVJeyBxE6
UgAltOsTZJEczeTSDlxejxTQzM1vJgXZoDOzFU1ivcKVEI/8O68pGOdOfFkZDA5BE/q7ItmMxCao
9sAOz9NsvFgiREpqMZu/7CEz1qhZ9KzCSTGA/w/5Vr9S7V85cTGIxEgm+lfEOGQ8CUoBu8I9k7yB
PsBRmqeeRphtEDKZ9kckX1Qu4ofnBCBk+K2ozt2h9Xe8O8ThXWP6D2ow2LM0U4jPTgZVnmOB8QI6
p+RxwH7KqBlLGW5wPgljlE9PvDgmiv3rIHC8BGF0WAMcjNeSDLX8KFPztkuqYXpOQU70EGyKvJK7
FJf3mNCbndHaYQiln/dIEXWars9w5ZNVrY8wvR2wT3p8HU6+gEaR7SH9Eserax9KgtxhS5JTTkzq
kSxPluz6ceKAtCVH4ClUAudyJFCpp8GN5GDm9xvs+0Mc8djCKbNHkHRUoIpMlviurElLxiwOBH8t
6s5ob0qNq91xud/K0HTzrJrZ4H40nMofKgmb03TgLac4j96gvjqBKRXAoE2ZA54nP1bfPklzJogn
7H/H89a3b8m8lqSn6BPfNUWQZtSJE5y8nbjBp+wmxvITDW2oIYlA3zhBkFMaxax1c2Srwbjwe4Sj
0BlmoeD31J/4Fx3IT7SuRO0BLaXDEPLZJJl+z5MCIJA8G316Zu4u4i65ScBh+sya0z0AO6uUW/Xk
1QTulqQIQfDBXZzkUppCcJYE8RHEtzXxF3IMnNNCEUtwLPPK2WVpH3qvEUSsrrrokMc9m3V2kIOE
fInPJM38nJhaoMW2lHnwonJB+q4X7ACwb+lf7V1NirPwgxaDjEyBWl0K46zMFTtpeVQSMbXSno7a
XOdmwnB0JqmssDnxI/E/O6arBZ+rB5JVIY4XIjp4Keic01YFTNgPiTF0fqQVf8MyLbfESkYyOg5W
8A2aonEx8ZMPFJl9T+Zfropt9lWkHpK4BS71nTXIOgvYR3nOA3PexEc4ZGH+opeBcJbO2UNmEipE
vkw5ks2YMmRc4+lq4/VfQALoZ5XjIbz+TC4IOkVWfSRx2k1mrLMfmOhst50bqbAtmkdctaCYZWKv
RJycQ/M99FiDRaBtzkvcctdDb/JjJk46jTyQJV8p/Jp8yS8ORPk8gOWO6hnPSKOmdyvKWKrbD+QN
Lb+/160oFjNg95qUHJJUH3A+KxxCAV4H6b87sCpTE+wsQfFtYSkQjqk4RGnRhshRyR2IVjcqPe9v
/nBY269Mwx4/H5XE8UglshFZjAsyrxU65IrJT62gUkyyUYGNiQt6UQc3x5erCxRCgruTPttAb7Yu
f5Dl7Z9+JBxaHxriZPmBJ0eTkz8cCQaYJfsIiymbuPTY3JDF3bRWEZq1Btv8rrgfQhrqrC5eR4rA
b/gnKSgV50AHAsDOdIK+piZXDkL5jVTMO1VZS+beVQ9Ia4uq8ku6Idg/Y9k+2K3Qb9vuW7+qvtVG
mAVOEu5QFSaXv0RewGdAQxBtdhgGrTU43mDg9gvO7B4uVN91LmgCNCEnWaSR3R4wFD8isP2Qungg
SC/uEsYRMCJbLliabbzM6MGZzwAVwPB6S6VoH5W4FmT0NRvKMiobPXyQcLInFw+gXZzj8QOXiNgi
Ji9GJnWMW4NHbTYj2BjDFEdCZbJnftz9PJnw1CQkE0mSvP8HtLOSa5R11Y0a63WlEDXnyF80E29g
Soazi4kUyMmhfv3RHukcqw==
`protect end_protected
