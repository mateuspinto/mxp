`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6256)
`protect data_block
zCtMM5MVlY89o1+WJaQBqonMfawtbttIDXUY2TVNwTiOiWHTyhGT3fQ3bmr/SKXY4rcEKTR9R+Lm
rvZb5YvkDqiYLMhi+sgyUR+K7ozGHCIa0T7brjCv25EtVAGZpDIvkNlWj2+FULJzYKOSWVYg7Ia+
yE+zxpfhkNY2gSlYGcOQOcmk0hSzEncv8XubTirR+MiD0XxtCJ1GkMnMD3YUvbQc7QY76N27BUaR
Mvh1t7jRQT/LVf+cAAbthgfayYt0Sy3I21a4a904ozsHCNWHO0Vd7Jy//JUExC1huT4hAxo2u3+S
bI7Fo7DIu8MH7iMNMBscLUntdxDqLcInH8Hs0B0JED5dh77deKjMdSClhlIAJGXKEDHMIZV76Jwo
j4YvaTBlqhT61/RICS9ymls4adFHRtPGF1RAeLep3hFwGxpO3aQxq/YKK95TqFiVYiO+kBPXrq6E
jJLjXUtxBN4SaV8nwOhFGWe8y1xorclSWvQlzVl8NfGo4ax4a6Z8NJEqlPRUJ6R8DLKVz9KKPqcY
A56OAGXm6BfSHBILOPTRRMRQxiQUZ9ALrk6xxttNGtywsYM4j6taYfwKA3wR70YfcxGJJ2/4/QLc
f7gyUPT0pwNaghUO+ZzVy5eontRuY+dfggjO0qRe4TZioB+9I0r+dsTY5GzdFlus5faNfLJRgDvF
ILf0bknLlwfyYLQPm3imENc9Hk1OCsNDAtiFpDmah12gLyFnzsgyMgOpasE/gkqTNq2+aZqVJL7W
Ims+kbm20cy7Z1QzcyKqDUpqCfQVIZkNb7ucD1yqc3TFn4t3nH90wXwM1bBPn8ucGp9hf0CLri/w
/dIdlNLWfOfybPWP5qp2sCAsS0Bj2dLZwx6S+cvOt5nbaGZP7Ym6/g1Y0J6hNR1Fvknszcs9F9Ng
ELPm7ZSK577OyAhUONLQeuaeJkeErpBvg4vbxAQQC4lyg5Uab2iJiyBvWxwWBnaDI4Tg1TcbmNfJ
J3rP2cI+OZMyURZZSeXGgW5EVE+bni7QvFdumXFne4n5HJrnx9QXSFtYRmG44uAI5ku1gZhh3yHo
QxHg2JaMrUlcR+8oq/wYhbsKq4YwAweyaz+7L0MR08oMBvoHe85WTsLDnOfR6+FsklxDuI8KGFbC
bLcfBI4OedEMVoXyIOIO/+lTMiGAWluLdnb/yf3vy8gEC7/CJl2XUpWZMfzR/XHQO1HIGaUI8rJG
WR/M6DEchflTTrFqL2JmmpsZ5DGrnUe29sd55bW1r3hQi1jp01kPtdPH/WfS+rBWOc+KXRo+lFNa
6XcKpIeyYQ3ju2OQHUv3l2EwVL6T3mR3WnlCINRO46SuJrikgiIUNVuY45XC4yFUNkG0W0j4VCCF
wOUcX0fMVeh8bw1vhy2RDzQAfT8veB25F9nrvlpRauqUO5vXyIzrITJE2bWQQAawGKJdugRh/9Sz
aQfs3rwD8Hg1x0b242ImcLCI09MmfCNxdYKHtE9t+HZJgiD5gC502wDdgKHfat6EWozLUSaWVcjz
KSYVBi3qZXoXtB0/K4V3fp7jnCnC4XWLbqRh18H6fEuH8j4whQcoy3ubmCwMdhwlUluBiyIwhZgZ
kc7/I/TtIKUOG6kpgP31AmgnsTqBOU2l+zh3N4POI0LTz5WY2NsE6oKMb6NHnbhl7x5vFFnwXwtH
kfanpMACJ9WSErQGqY1K0j/YTG6bKyAvvR3RtcMPeFk4s0pdkiWCZmpJuggxIB3PdJKn/IuLxgG4
1OG+/LTbPBiKjHnxs5jgXjbXmN//XDUromRtikcqkr4WXkhACt+4+KYmAXDwaecSmSlvVRbHbS3m
MEabZyJHS2M4x4BIDLtoIAno0/bvwSlGsYpSZX8rtM4qY0E9cP4ZLmObIk90LCJqQB/2lb4IrRHY
jMOwiRfZBXNzqvFJ8PjWiLC7ADNkBw0n20bFRE2ayDgzQeHOZczcW/quCCtceDtw6TLExp84Fn4E
YdF5FAJuYY92yNnFwe5gnG+xL269cuxUvFNS7b19oG9u2GlguJ29sN/WRGGe/bzfalL36tymrnE0
nR0hY/0Y9GDpVb6FsXEiY/EKegGJaZ/x14/Tpqbg9FzifuvFR79sL39vZQ7LUt1MmFjaXntoBaVf
QDG05pWaTKKYxbnxaiiwm+JsQbpv/Nx9ct2wWgWgeccUVFtcPzX6PgTVJ7Q/5t3EAHuqWoY7gcuJ
rgAe2KYMhNEVMJ63mVdH2wgDupIoB18766ZyOkI2eQ7SwoxDSBzYZn23VmNzim7HQC4GEYLOfNL4
sB9oIf1ml1FyMPJaWqcSI+mer0LqgNUFWQu6dwO8qtn2ZEHN4NPYDpVNSOtEDggwGpWTRwqUl6Ud
EbIELyuQd2Z4pm7Ga6UqgVVzREKHo/DXvU620iHmjjswjyD4TnQnf1ENj+PqHAmScawbGhiondR4
Bv9shasuHkLPhOAWLuNqmhM0e5fHS9if9MnX/OG93az1zS5iFT01htpsXCpXO61jSdzLkxsw8jBc
V/kyo76uiepKiMngUoFdKdK61K09m63TJos0x0pijbzCtUgNDSne85+MWD/I9r7j12vMMx+dxF1z
j6jdp9Oae2LhQCgq83/tPrA2E9OGZsXMVf++WnGVpcCmxn8XRy5n9btIrt2+cWkxNoprILGKJYi6
YeiAisQNUb9eUTKU2wPkH5Kp3+8vUgK1YfV8Zk+c879kvmBin2opN6LzMvJ0DYccVafjxx4MHe64
iQ92w5kBdj+vv9fXcXaAqqAde2l0vi2hpGABXIUUjfqOxrOO/pqecTfZx/wzkrG+/7pOfNWB9Abr
aWb+UuIOVu8fhOKdfco4G+jlXhay4HXSkygKUs66EiPSLDRaOdiye/NpPnuker0O0ukDmNuGSemK
I9t1moYWMZv/mgng3kNlvt/UUtqZF3yiLPePoDb3UhrnBR7T0gXbt74wAzg+SOV8vBKxPKS9swJC
2KT+v853uNKcB1VGToNAWvCcbKubjw92e2rMkZHTy8spSS0wEd9RyQHPApPBWz+wHjv1QNOmcH1p
Iaohw2wfZw5+TnxzhnRGZm3Oo9u8jXTbI8iVKSe1Eey9LWCj0BJlt9iciTywLujc+MvzlsIH1Dgy
KgHiFH+1UouknX3gSr63VZj8i2gVgj+B5KJLiPApRFOW+ditCpBV3QFdBWD4bGhuRpNXbsm+FtCM
HKN0I2yrTlEVDYBO/eWJh7k1buxk4j55hgONeERz6juKNMQ6uWY3Oa7ko97fQEfbrNXZ+h9BY4Oi
yVW4CMVzhXTkWpPlhd1WwtN03gJkoOilWvATB//7DSycMUo34Op/UhTZnJvfyGCcEr7xVO9Z/OLg
JjCL+H70iGa7/LTD3PvKDAMWH65piE4HcAVmnNviTB9Fb9CPGejzLKc+dhh9CaZMNtI8oINCsSO7
DFAUSEez5vB8pV/C92eX2C68pfd7yAs/q0r+a8rVtWcLiLS4cdTC5lZwaHWIPXXBVmbFFj4lYf1g
A0mvPPQMlJSZ7VxcphHODZbNo9W4A+73ePgzVQ/7Guqb4JiDMcN0OOJJbjEXPQvC3ZnspoIrhhsu
gExPuiujKQyzWeHY+9WEyn9BsMdWimoIS3i+pH04t5wohXJYpWyA9BQwLdJJzO3IMxMp6PwG72zh
F5Y00Vys68KI2kFpkeWaU5GON/15/Nalx2UtiuXz8SGYm4bSU5/Qnl3yFPtuzMMD9new3jif6WeS
3dapF31AypZCpnVynxtzTaPehE0uod4dlzobGpZyTC0mwwuPuiCFik16h3P7hvVru5QPEkoNwJ34
F4+HlW78cufFG3IeUcg5e8Zazh6as4AsNh2qWoYzzzjb/IS6aLiBhO6tR7kjiUj0kiFYme6o0miq
oh1EDA6tdBCHZX09CAvQhVleyOdwG/fdKCcpVxGB3UGGLnqrxtwBjzi20iOKQDOS+2W7auP+1hZp
xl4PkrwVYGRfrs7rbCZB+gE4Tn0bEgj6qY7/68tfR5A+QyVjsqc+SYZ/a8UKeNbi7eLTsgAngg0d
i1cY9HDRX4ngqO2UphuaI8gNudwvdADIpx6vYFmb8XyukOhCil377TP1f2QJMjFjbqZyBepg1sph
L+TlFCdGoweO+iOaQ1/AeoJ9Uzl9cBea/0499/5K6wRN7JGHmMWuV9xzLZVVUlfDskX9ZK7HHb0l
JwwwAynchiBJ4Pj4EBx/xbEf0JCJSrddl/0baETPrCgrAbVsKksdFtOnVOrI6GxZWkYYjUKMLbFT
B1gEKcJKLBGjZ6YlaNCENgKk0RByzojePbtUZjEGu1h5yNV/jfQ7Rpvtas36sc95OIbJZota8gn6
MGBwmvISbz7/rPwWO2egiaUt5+rFK1uRMbJUbBuCzEAjyWcBsBWARox1dXGB5eGixu/uwr7zLrSh
0ki0IF4FHGNReaKx2zlWwhVkUqN6xXe+Wka5RpkWxUCLNxCFXJ01NgUvNKR+tqPicGloBnwOGgHk
1AZYlr+euBmsyXVYKa6n4J7HN+su+GqbHywIR43F8amqGfmjCrPJIte+rqvC1ZPIdkDD47ua7Dsf
LZJo0Y0TmGqpj+NbYDqI3pDe33ypPtwUmphYYohg7+TLjnb0DH56aQzAtaH86V0rCSox2X7ot0Ss
J5GyQi77Hto8DYk9zPexqzZJNLNofN6Q41yPEapeZrJ/t9evoNKt+8dxi+5FPlYSdYyG8wWC/C4V
+ek2HWgDtXLwJA69K5dnyLSTr4P+GGWEMFX2Myxk205/VOjN5YuDqgrkbdBT+KNO6mhDTT9IhBZw
apFShTHPkfaUcFavQAYVjbsVGbhxQWFzrMgo37RuYNr9/Wg0EW8sXbtadSfAYueUiH3vdWhiiXOD
tyUVIzuBKokrkcM89SODqr5iopuYbQU5aLihQGmiWHZGOKdM3wfV8rkRxiJ54bDCCRZ9lb98BjDP
CpFRR7CpEUoHLMo967QglMTpsI7rVc7Ixs33NjUfFkrFnbJT2c6kWkpm1VwY3scKBGkWKvHqshHP
BMdgKP+SC+lnzzGrC8UKQ7YSFkDIOypnqbLicb8XiHBs6mBFjiif9Aop6immqnRxVCW8hHGl+RWY
HSVHxicJm3xAF8a2yDeXD9g3tSwV3raRgyOo9IsHPN9nsxZrZD1Txf5P4XO2vaJw6L47eZ3v/wvg
9bWKH3wcoTop+Pvr2LvdAJy4nQNZ3UlDCDGJdviqUKVj3+VywE4LPkV91LvBsOAeLfMs2wbMRZ/q
0Dm+iWzuHkseVYZCgQfa//K7tLv4XmEIF3K3i4lUnOGR/BWrKBMFacpNfYLSyv4+glmxkbfXvJxS
t/FmU7l6KNTH/EU+Mok8xWMHJLnkN3GCQ042Xt44aRC8sXtE9Md+8nHyYh6xjtXRv/pIf2CO4+OV
prMwuYnH2IN00rTpD4JfbZhH/YgovHnCeYsbxqfg5xEQzD2f7aRJf5/PnTBBTvTYupLf2MYxiuyN
hles8+k6Eq5MJD7DqJsdbfXxCPfRgE4CBQGJdPSbS+HjmzwoFagL6QbQ0WTCCVa5eSsNbWqvqvKK
WUFMQTsDpnRrwUcsopjxAVdnFgQKaxdGF54bXTzaAPLN1FJxCPeTDQtdulDNiCTurH4QGZkxPxWF
4bsfgN7XV3Jc9gdI7KAAAqtWzYBe+dVdib0jfP2Ho0nyXcboQm+I1o3bm1zNJjmf80pOAaIWgjN6
nDRILC2+o7raHwm2U1+3r4RYSkZ1GbR7+Hyh5xx2ymYtAf4TfRyAI50X5EjO9pkwCTJwdbTFg6Zu
0XuiG+mQNZQdsHj22I+4LoCU+/ZSLWkiayBFLzeQo9x/mFhIyLVY5PE7Uq86Xk0dlcMZEGqaif3g
1cdwwAg4VCLdo3fxdQZlxuIRe9q/acF0/WHM8QtHBV6Fr3kq9B3rl5dPCat+Fg71Y9sqRDJxnrOU
RBIZso9zhFn1VZcLmO1NeA758b06aqq6nE8yxCkUxrnfp3pYpe84lZW75ilVw4eNFgzz4Zi3MvGH
ZH/cdvarvZODBggFxvPhOAJ7FW0eEMv6L/UMXOyMQMP7EyH+AheAeGGolYSjdtVkr4CNME5g8r/N
bYNyVAqZYF9Iaav5eDNQFKOepZ5OnLUPCJjNajaVHTQnmWDsXlyOH0RZf59xb7f4JCJqDH8Fr8qw
iYdsOOfpgwjL30CAbqU3NyZfGofoURsSmqXu4pdwGZqsBgUcy3tkkluLQvoH+uvBqPEtx6/nzaKR
jxmCevVD2fNijyl8sYhO22sykPLRBsNezf7+1KzzghxkDT/KozeUD2lqRjOANy2JDwNzBtdXdBXn
VQ1tYlIzseAZS4kPhg50vynvdnB+fil5c1/r4yaW12rHrPuL/BpHJsai+kG7aBFU6G+LJSV3JCY9
JRRqY/185KFpGhDBFNrBWzKmJKjcbjyrERK/o1SNLYQ7nUrJL7tjC6xL0EVT1Z16JhvUHd1AlH6N
wX0py/h8usnWHwO+MeE9ywTIBYE9PWFuAuO7zstNeRLqeUIT+xTsq9poGlk7l1bCXD97tl2I1VB5
a9xoEIJpL7UEiw6qyMdX1oRnGBSeVpqqhje3MGI3rN1W8KBOk5GnAwSu1sEsW8AdEIopk82UtD1y
sYLOl5v5rzumr6AElZXTB+lSxFHyBXl0rAvh2rBSkC+uzNWqKUjynt3zFYEaepSY+FW7Ge0WSd9H
uSLHCxljsP+BkQKKyfBsZnW0qnGZa56ppq6sGnYjLsALZ2GvocPz6Tjp0dnxb+xxez5SG3Ocbg5Q
iyUxOMXdwQwho6+K+6oUtICpn1KZyLTHbQjun042zyDQUwRaQgk5uoJhTD5YsL3i7iVd9zob5NKz
jTYsE9bjiwYBp1GOrSIdKmNNwTNpDFWcUILvcxp9yo2gZFZTYALvEBjF5ARtPf7UipnB3RBhKITe
mu9cXxaG3jVbrDkj6weY+4AUsss/XHbQ/DsahEUDojiB/JQfQudk5ndh7RkrmoiGtoiV7UKaj6vk
fb1tZizhvUqQ3t2dKfezOE7jTEFODuzRLUJrLu46Gwhqrk5Ng6rf5lAslxvYApk+RdHv8PCBzfIX
4xSDJHHtWqyjK9TPdlF9jMtjhO5GSlGumHshAHxUITtaGJ5kFJsdU6qeiy86GPHI19GdvpDGKBGb
QP9qCURxC1kJGLB2eg8qFEMZEZ04IBxh5SHoRmykqsVQ8KaLm+wa8t6E20C0XLuOQvm2jzBdMwVV
ghV7nnwnzsm3UxDKHVViBANJAZ06sq1+aOY7o7huUL7MxKdOH1n8V4VRvlLCOOcSB8PpvdgbNprX
4SdgR7TDnoxkLbprdMz7uhFR4CcKv5quAihbAqg+UF3gum+dO82vySDLZs2RVaPcK+3j1Vpcn9cr
8JskXZZXDs57oGRPtfTmtckRO6egWkG0ge8DCrxtmT4YzM2EzRYLzRClz7SKSuL3baudO91Cl80c
gKMEQe6cb3V91e7hoQjQHpeGoYopanUUzFm5yKLWkXVAyLy6hlLbFRcXJVjUGKhr+49nKEo+RMjb
W76kwPpOTS0ME3tqznqn8xbVhtENmB5WZxjmn5vMsF6T1YkG+PewafBmMwHQTPnn2VLX8POrSfKT
i9cfwpqbjgvqlQ27tYtUlZNyTrWv/c+ZNlff7PVjH+btvhRS127GT2Zj5XSA1FMFVMJZcWADCgED
S7S4g73Vj71ufb3enD3+8Xo9W1xIkb9es1La1hGEW6W8jvXBnO6KYqV3xjx5WtRYfW4BZvaLIMxN
kZbO9s+2HEnzp6ClLC9eJ+P5p+4Ue/IYVvAGbkwZ3D+8euL++SfbcJJxrrgHXKxa+d8WqUrseOAQ
4Uj3WgKwdVku5NwKoLhtBuzFFpvLfz7/5L6z63T62FiCt73ewDCYXnmOHa1CXYaKLnCnTUKiho9+
jyzKA5+716xS7yqsjbd9cL015D0zBTcjxtW/M2semyGyeXbVXL104X240vXKWbobHHCOJgL6KIir
j/RWaGc3IwNTyhqHmuVwTZyNdzhIzykmvigAmgJDejecAOPXZJdlVfWxP3rajo7AUj+3zK/ksd18
uYeXQ9mEDU9to1S1YrHcH599MRtm5R8n8ZHw2fsCgB7TsZ+pT8cJ4aefmWdkk35mOei9OueK+gnk
ddAHrzR6mqgoG0oxGiHksl2E1gRHYkkbGonfHgqUodwdunCr1EHIPEDNS55q2Lhk3JJOBn3s6SsY
Z4vkwLmWk4kGOTTs7CZ80eYB7ImKtgFIng30u02WgiBeM0h9mFZluLFVNLRHYjAkktYGzp2ZXhRQ
Xr6nFCnSXyhEa/M+In4skVd2zZHzsuMao1lj0NuakBMNm49HozJLzExaXA==
`protect end_protected
