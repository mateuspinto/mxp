��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���L�n�����68ۇ�fa�F. }?DЄ��ٜ{��Hz�(�-�Z��k=��n��R�5���K�:��.	���S�Y(>x�?��6�e�Q>�����ӛ�;�;�3�iE�mDS��wbp&$��wMθG�Qb�
�[8�y;E��B�sr���K��Ċ��st��5��΢uR��4�|���x�.G�F^��y��w�o�f�l�dp�3��@;I�^)Pj]^L��|c�#Gt"|Ж�?���3J�'��c9�����&\� �]=4'����(o�C�Աr런�UfYh�@��3M��
k�e��:|3�אn�	�����s�1B�I�g�p�ÿM ���V���!O���<w���?Н�U���=c����֟փ��3b�_�������1�۟*�{�0_Л�+=R7m��g�Ӱ��|��yL�to���@wh7�u}�A������"x�ʵT)F�I��,�6Go�mWؕT��62������&n9<��xoI�tneF>Wb3��Zf�*I�����=���_��.��QmY�<�!�g�x7ΰ��º.)7�/�.��-�i�������j�2S~��R3w��S〣���<�Č5�ޞ$thK�ΰ�{fC�_�N��&���:���� i��x@�J�=]�E�T�'�Z��4�w�a��q�SA3��y�������Ӫ]mO�^�h�8H�}��;щ��� �m˶�q0(�?1����]K0
p��7�b��j�	?G2x�ڇ��u���u�*��4Ӯ������~d��h��V�s��v��ٔ����|M����R���k�n����u'�g9���}�ĀS��.�by�ہZa)��X��/#��Y��R���kv���|&�}�����Bř��.
�v�8wS��_I�,�0z����*����=��e�M���wT���c�܄('�馬'q�8r42��OZ33!�ԃ벼Q�#;,#?��~٘��6�Ÿ�<9۳g�YK���M��lK��ʙ���V�ՠ �y���;jƤ��e�M~���/��j˼>��ߎ�����s�ª1J����˒g	�5m��BRr�!��~�Չ�z���� )�"&eko�	MS�x�j� �0�����~�U�zɻ���*ϡ���z����;�fR=���,!-�F����'�z�Q˙�޼�=�u�an��m�|,b�����bS�24���[�E8��k\����5�%f��}"xM'��@��]�k�g���ws o��*Dp.)����j��4x��+Kv����;����%8�Gg4Qd���\����J>�,ވ���V�!��W���Ji�P�����W��Ʒ�`�oB`��jO���2������wt�������M���c8���x|EL��wۋ/�~Q톲�1p<���Ǆy�5L~��@8T%�F1��!	�)�H5/\�"`�O=�ԊH����r�>�݃�8_����f]� ��j/�!u��̔�T�{ �f�^�We�@=�1�[(,�@d2�T��n�����H��T��]�v��%����+@§�R
���Z=�	�h�����£�
h�sQ,�<f�>����k�Ƒ�tp����	�a?R��(1��P��&�H�K�����Ŵ�q�@4�	��{�G���|�HC��m��}��v�C8���O��Eu�k�Vy"�*�ׁ�5���"����@�1� �� m*H�6����?z�%�[{pl'��;[i����X��0ѤjQn$vZ��*;ƕ�
�X�_t(�B��7�M�����k�����(l��u������ÿ�x%��{�'N�ʎQ�/2l-���%$6�Ä�:}�)]�O�g�{���V��ʸ�͌��)}̰k��+>�懍� �	�)�=L�����m���_�q��D�+���̅�*�����5Y���w��6��`��YR5?&�&o�8�P����*V���sƖ�F�d��Y�]%!r���~Z��>�0B"�u���M[��.m�H"w�T�a�e0�(���|rn�ߓ�׸k�A9���Z�f�� u��iS��������CJh�:�;O�/�)�.D99��q�+Eϳ�
����K|g���}��E���R��jK>�V=�7l��`���Pt��`Th��ovK��3���$�aJ?�y�hAbr���sXޚ�f�E��b�r^�}s�.�r��Zx���65w�csfj������.�z��q
t�q�D�d'%�Rv�p\�~T��)>���w��;q�\�2��.�um�_<o1��g0�Լ}�$ȶ5�1v�n�݋k����7�fJ��w��k�w�)�q�+4��9��)aְ��EN�����WP��\"6��jtڭ��\>����RO�D3B[|<p-�{^B3�d��:�k�a�?hj�S|=|�y�Gq��]ȇw�4s���:N���u�T`�e�4Y� ����%q!W������n���E�ۍ�˻�w.���_�TX����|{釪k_^��}����������_.�����^�D��U|1�H(n΅�<d��%�3	4'��J��C�ʖ.����PX]#.�L\X%�4{S6�:�+��ei=���D���f���͋Z'��sO��Bno�p*�2�X�䗣����s�6��d���5�"�BԈd����$Ð�v�R�d�+uL"�3ZU�,�2�?�Z$���W-p�V>�j�PV���v��U�PۑEWM�"#rS��?^cO��C|��@���2��';�9�s6pv\z�L���^���	�M'��X���Sǯ��$�ΨlGw�մ���p���+���c��q}-x9��g�1=�|�І���L��E�
V�Ś�������$P�'�x�4~Gɡ�O��W�"#��!P}�@�7y�D����+l̿�9ǝ�Gg�tA�(r�}�Ү9��b��@��z:;Y�����H����H5�	�A�ڢ�%�)��c	�OI51P��GC-�Bȕ�(d9�)m䐺�3Lr�HmvflY�U�I��m�T��%S�>[�/��A�z��"�ܸ�i,G���n�*��+�ц��rc��é�e �ըPl�K@O����ZT�4]ܵT(m�z܏���hy�1�1�WD�7���	�n�g>��P�X���$'��aw�9�4Ƨ�D��E;
�dC8��+G�֒xy��)ٽ� zL��Hn��[�8.Ũm���`<���I�t�ST[|F�qj�����y5~ꔔ~��?@���� g��h�Or�v�׈�L~cuG���5ˁ�����A0Z�;���i��D�A��^�7�Oo�V<��)~�@%ᘏ���:x�o �ڼG%�vjt�����b�{^{���0��]�_�:����\H�gL�(g4$〰��" ��~z��Pj_a'�׹��Kc����f2tyxv;d� �\���9�"�~��LJw�(��G�H?��ҺG��W}ey��Y���(�
Լ�Ԁ�Dףn���jDN:����9���!�To�n�{�Ҩ<b���E;X9�a;��1RT�e�{kJ$�p�i�gY��Ze3V���E�����bA ����������6�'	��3�}~�qX+�C���7�'@ɣd�\Q�|����J����6'/���W Ne�Yۃ�y`��}�M;Y����ۀs7�+̪�l�֯�<>�\s�$F�I��Ѭ�:Q���?��f�/�r_�;N2rw��&�S8?��R�t���خʍ�Y�dU�<׏�e~�h)���]{� t�_�� z��s�)��]�!a`��X0]Gʼa��$�<��i:���~��v�՘fC��eA�rˋ�d	S?>-���0��R��2 f?�����	-�.�e�q�$C�:��@
�yU��ȹ(�b�e���<�(\ĜPi��x���3B�䪺�ʟ��{;0� ���
gU��q�?�9�s �� �ܶW��0�(r8M`���������ax�x��cW���&��H��ս&�V3n� 2�)����F��P�NP��-�F�2���d�:7+����o�Ssf�/��*:��(| �3B!ۊN}Ƨ1d���H{@b��mXbӅ��܋pW���Ķ�D��Q��xa��Ar�Ï9�=��c����7�B��W3�kjݮ�����P,P�V�ҝ8+�꒤�I�x�E���-��C���	��8�L�M�ݞ�7�7_O'�������z��d�M#0�vҰ��*}�)������+Lj�i�Y��1}Y�5���˂�����M�.��[q)DB:����#����c*��A�-Z$�5.�zA�t���E�̥��N�u���Fsh�So,{�H0mM�c#l���I�W!�<��o��ree�M;��Y��_Q}�3S�3�"�$]Y����Zg���#U�T����d�Mu��fS� ��#������r�~��@>��Ez���_��i��9WG�6}a�=J^5�Ly�5E�h�v�<߾V00��a�=�Ւ������/4� l!(:�c#�q;��HߋUB�毥f+
�$���F��?�8���p���' �;�Ϝ���)�HKݸ�,�isN�=�'��I��a~1z�}]��x�֤�&Dqʖ|BS��Z���(��y��*���[�@��f��tf�P�-��I!R�*s��������"���)���q����<���(�����< ���	Qk%���K���7���J�v��o�Xh��`�i)�?���I��j�
CW)~~��1�,M�覺F[�+1l({�>�z���������}����uz߈�.H���]c[?Ix* �U�I�0E��^�p���c,[��M/�^��_eN���j#uK�F��f���G
Gۑ��'3'x�������,�N���Pz!`��~]���^�ܥ�i;�t�5b��H�e� :�e�mҭ����[��&��E��!����h鱽I�Yj���r�����Ϳ�U1���@� �c��FiO	N�[�S����:�x��;�z̍��1��>�ѳt �RX2���C��p
MDq���$)S0��.|Z(0ǆs�u���K8��K����������%��E�?��d�xMdd\��ʼ�6	��Z��"�(�9J`:��Ư嚎�=2<Ff^k��m�?�A�6�w]�1�������b}��}���헯);�)~���Ŋ�5�I���5�i�PU�|�Ws;�����<�g�:ݳ�&�޾
��\�D%�3�@��U���:��h�H��a[9�r���\,��>��pE�O�_�a]  ��uU�8�Pe�>��H���)/�Xd�Q�8��A���俥�w���S�m�������3� ���Z�}�������,��Zi��ն��ˮ�3�[�X����n^ �y�D��qgt��rU��e���WMԴQy��oF�;����@'_;U�^�d~�\X�=���B�g���ђ���xè������| y������,�����&몠���Չf����r�A��+69Eu����2*㼝c�>��;<\���\�� ����2oJ�2fﳸA�1B�W5�99���~��;����k�h�Ē�³�}l���G^��z�B+Y����?�=��"A$������Mj�Y7��'��>>�ٿ,��Ek��V�@u]���.{�	,���2�Ty'ܰ���ЭءCp�9 �0�� >=d��K��S��ޫ��!�����}����z圼I�ZDQkQ�'2�tI"%��i��p�j�8�L66�\r����ۥ�މt܏F]J%b��KS��_��oD>��h)lwZk~2�ȃ�>�;����%Ѝ�����J����z{V{$�Ak!:�O&sNQ������$���Xl/���ـ_����bi;��7�r�a�� �{�$�$���,�����K����D�3��rk�Xd�z��Sd��#�W�n{IV�&mfO��h A�}�&&���{�і�B���t���+7����-�`���|���q��<FO�wݛl73��M-�*_a:	��B�1q�!�`�����l���He���q���&��p��	�;�j���Lp�w�"iV��Q�6�"^�AC7dv;A&=ar�M��t�p��7�}b����rA�����5���5l5���H���PlD3��Z,ۿE`.�Fp��U3/$⟍�X ���Į��i(hڣ��L��A�T#:4fb��N�:2i =����j������@�(�G�+�@Bl�LpJE+���;��1�I�[�t���qчFyr�
�|��*�X�Ѹ�f���x�{(2},2���p�f�/�d5͓��z� �;�ow�C����4�tsc�+���_uZ���9�km�]�/��ߋ�փH���xv� �������.A�����jcޘuG��8��%��(_�<F�{۬[�{%�iJC[��l���5=Y��@ak݄Nd#`�Pn�A0�����8���ms#���D�sfh_97�]B�NH�Я���001>D��8��?+���O�Ú�k"��$^�G��s��q�|��g�����qR���7�X ��������m��|�A	�WJ(����+H��m��J����r�W ���ӑ��t`P���%泪rK|����	&;���y݄J���
%��50ctކ��"ڞhF�>f[Q���b�2��K� ��
�#Tj�8���f����ڮ�!����W���`���^1�G%���������H�f�"��� �*.	��$�,k�ˆmV]w���0��0ίӀl�J�H\&�q�n�^�]G�>�tQ�fh��c��|�]l��#��r<���m�WO���n�#8RW�
��//�a��B�m>�w�5��S���x
�")乴���-����MeU�"���E��΀c����1�2�i�k+����8U��L����<��*���Y�������F����0C8��y���fXuP��~��}��Z:L���;�ʡ�n>�a]z�1�vH`�����A���&)�D+"?��<>�B�po!�q��03��8����`�f0O��cN�����&�b�f1�t���v7U�M&,�H�F@ҼW���Z�a�8D���sҮ>s����f���9�;����p��e*z�n�3.ά'����Ѱ�Yd�T��\�-�"�I&��z�qcƲ��[ʵf8l�H.A�I��՘S����K0�؞̘O��l���Sx+����һ��������X� 	�2�I��mH���K������fqY"�ם��A��d}o��H�\������,�E4����x���?yM��6L�'p�"�9��D'���	��Е�c��u��{�ń��_�`G ����c<SC2���p����	����4���.�/��Pp9�0�V����ʺ��q1��6�f�C��0��9�>�	����dMMalm�	kA�+BW���E$�������x6Z�o����:O��c4��N�F6z��WEH�Q��x()�n�c'㊆����O��3��+C���EDP*�1xi��D���ԁ	1�&����L�k���CT��J���2!��
z+ �ϲ2͢$T2�nU(*�A�W�Vf�w��ڙ�֓�S7�-ȑ�5Y`3���8X�bxWۯ1�2<y�"���ً�2�/�x��M�6�f���#g~�ݸo���e*��C��8�3C����`��!~�$B�Ojo��B���7:�[��S|�v(�o�ŗ�&b��|�ڭ7=�(����9��ɽ�\����!W�׋˩Oà�&Ԅ��`F	2��둘��f�KO�\�BqkF�ڀ��?{�
���@Uj�[�!��S��'��'.�y|Ż�r̞�����Zu%�^}�d�/bkI\�7h.[�z*�.%�	.Vµ���~ �P��1�%�!�Lc��`C9��Q���Ȯ8��|
&�=�p#�1��t! �	�4�g�H��I+R�9tx�F��׫�ٽ�Q�*�.51�J�N�lOzd�K@;���V�� ���I��w�ܛ�Ҁ-X:	3�����K������b�n4�����&6�?{���&���!{>��]��Tԡ���U�/l"�Yi�,<y���T!V/B��''�����L�j�+�Tx�R�k�5��1�����n��+�t�Gb�P�k���о]��C��X\�k���2aG�XG@��J�g�q,��4��
r=K=(D���t�F|J���4(��A��gG�d3MO��c�+�y��ii���&3�݊4���D��j���i�X��<��8��ȃqؼX)�� 5)Y��T�2�� {��,Sɸ{H�oS��[�2�H�#��&��I~h�����|�ӊ.ϣ��bc.y�˂^���$��ޔ�YT����ħ�d�H%���0��<��ӱ&��m .�$=��1��Q��
u�÷��X�N�{���T�x-��2ē�ms\�d{��e��V������"�\5��]<7�oL ���-�����D9S�dȃ�I<H�Y��ǈ_�yTi�5X�r7@կ����� -�b��M|V��){���"�?��w�l�����M�ܫ��_�w؂�R����]��C�cj�������d�����dT���,��n��M�O=�}*�I�Ћ�˃I#E�����A��9���e�g��4�i�s�ͨ�n��/l2G��C����t�j��ZcHӵ���}H�X釭ӟ֮�����X�8v=�Z�m}[�s���˒%�f��\�-B��{��ɇ�{����ǒz���ү���-�"�8�F��W�:ˑ~�7��7�Z��!��(�˽Ei� l:{���.E���Q� �!�@��B�IH�#��)�����N�a�U�uo�H}���L�.�9�f=���-�y�^��ˏKH����sYZ,�)O� ����3��-�a��͔E�������ϴ�41�Tlj��'�$���po}5f�O��e�T�I6��'��-�M<�o����05�i�;3��ւڕ��"�Oaw��څ��Mi�;�L�V��뙉s��0�^$��_h`M������?̇F�#Sģ���* �Y��p��O�OUU�Ux>@��De}3�=�ũ`��d���)깆�0�l��<����rz϶�c��v@�ejƿ�i�,g%��*8�L��Ɲ�!`E�Gyf��{Ln��":�����D-��3y|��e��.u�5�r�u��~�	�d^%��6!��	��6��W���G��G�U��-I�3�{x�5��U��j�!	. ����nn��=����
?���N�6�C���>���{/��¥�)��
���#�ަ�So��Q��$��t��Uvc����=���iv򞯹Z&���� LA �����$T�1�����*w �+-'�)��mL$,9��zaXE��1?�bf�����!��GΩnofo��i� f��CA�mW�����M��!�	����t� ^�7肌HI��nrO?�p�S�8.�k�@���o-�-�:`�_��)�-q�szG� ��)���z��XA�t��m�*���E�ii8�ev���n�no��?1�a#�=��ϥ�wZ��_���9��9��H5kw=�R��m�*�y%��䈝���_����9�N���S�H�X��XZ�&M%w��\���.a�V+@
�� ��?Ȁ�N����`nn�����[�r�4�������z�be�j��Rl=�Ͷ^�~�fAh�함�2I ���4�e�]uШ�]���Zen���)�{����O1X4b�n(hn�^u�Po1��X��B��O��Ԉ�G���q�`�qw�F�8�7��a�t��l�����:�k�%]����Kc���X����p7��a��y�ଡ଼{S+ 2���c-T�`s?��ty�rG��'���w�[>T4Dn�϶I��8��9��4.��H���Q���``Klgv��A흧��:Z�Ц��Y֠p,q�!�ߢb5���"���C%>V���]���򸅦1���	��Y������,�J���Dȇ�[���P��#����f������*��Dl��[���K��ߓ�%p��z(��Z3����^�m��D��/�>b_�&T�=l�	��3���V�N3J�[��ދ���<.���((1��*nu����Ï�^�#��E�1��3�e��{}/<�s��hE�J������n�o�a�T�ط�+ ��rr��:wI7�DY��)�@x��8����<q��o�0��Xq�'g��	�fe�̦S�����Ġ;S$7G'w"ʱ����;�>Ifv��cl��O�z��4��G�H�֘���`!�6�@� �h�*�^�Dܔ��x�ڦ��W�I�s���M�8(�|�(�9�`?��PK��p#���J�qޖ����Nk�};lF�u�Cb�-�N\�R8N]q�/B	o��3A�)0���Q?�F�\Z��/2�?���E :d�� ����̘e�蟗p^�ȱ/+)P��8j�#���n�#��XYr�N�п�L����x�&�aޔ��? jP�f4p;ߴ�鲚1'� )f$O�Nal��
�g2�Fh���i�j�����]�qtZ`)�,O:3O��*��&!�"�v��7ʤ�iVA��d�����[��@�-w,; ���Ӛ,�M�&��t��K��,�)#�w���yX�ڦz?�;[H�����bN$�heV��� ���Y�Δ�v�S(�g2@���&�Cp�����;���Q�Y~�����x)x�QE�*ڠ�}t�H���k��',�	���KSap��������n��c=�e��,�:h��� ���u��ľ����7�T2��T3'Mon=�HlR �y"kS�ؼU�����˞}
��~{=yő�5�]v��-�M�(���8�m�'5gmUFow ��G���>��lX�ދ2Xuq� h��I$�G��c�hkE!
� 7V����<���6b3�r0�Q�KFp�>��P�!���<�N8�?�ߍ���z�y�3���'�C����-�^�}hGg3~k�ۯgJ�eD+<e�>�kȜ����!� �V0�qb'6�g���^	�O����k��y�2\�A���꺻W#uE��Q~����KqIXJ�Q۾�D5":itZIv��b$�k��+p�r�� b>�v�k�T�k�� ~p�)[��f���c�ϙ1ӧn&��Sa�5�i4;�tßǴI"� �-{��zd`~�l���?:��+a譜�:�|��n�.��}����Uɫo'e �<@���{�!��C�.O��,3`�B�<�l���6���b�|�n��#�މ�]��&s���/iZ��lQ�i�&���V�v���"!�Wg�Z����E�o��"�����g�8Ym�M����
"�[4�`���N0�;[ԇ�3y���/K<V��M8���a@�+���<ሰ��Rt�Rp=����CK��.�Dw�QÉ�m��×rF�6na*S����Z�^�1ɩ3jY�iH��7_���ak�~�_���G���uY�H	}D%<�?��/�c���l<�����[-��_�b�'�@^j��2��Py"�*H��:�a$��X�0�c�-������y2���R�"��x	�A�^�8���*K�)�j�/���-s@{@>kyG+��ޗ2s�w��G`5<4�����6<�}�Ů��������P{�J�|,_�Uec�G_����`.zM�l ��o��|1�ɸ�L!?RFT�w�\=T�*9x�!`���}���3�D�,�Z����0�:\�*yo��� {!��w�\@�n�+�CùXR""ح�31kT���ϥ�A٣ е�;/!&g��"��O�%�s�t���0� {F�}输��r�,�a�_lD�9�$	s>�d�9,Rer�U!�Uw�; �pm�����O�T��ғk��'U�c;hT�+�;4�mV�m�� ��p��r�!r�/���,��'�(U�-4��p��ym =��:��)��>DRjލ���E��״���� O�"n���O�SR���Z4D]dV�Bu�B�o�%�O��-��`�Y�/�ՠV�l�����^!7Q֧���ڠ�1�֚s����&wj�D`�.{X/��WȻ�a�ɎB����%���zq�'�<lMs���]&��y��Q��(4�11%|�8� ���ü��rM,G)�%S����A���.�r�>+G���0�r��ߑ������[���q�B1+E�qW��<X5�7l���L���$���	�p݁��ܤ#4)(R� {#p���[хO9�>�3����P9���y���a��Я�A�,V�]y�י�c�>�M�B�	�I�R\�Y���"�|T6�o!��:k_��$�m��`�Jw\o}u�%�S����<�ّ�wQs%c��(��1	��eؒ�T�����߅5���3�+
-83a�����(]!qЁ|���V��~��O��6�T�FzxKj���|���f>s�4��W�`"����=��j��
��Rle��~ 6�+K\:�?��s�/ жPSf�tۭ&��-"�[�M���{�H���b�j�Ұ�g/.V@-���{5qQ\�OdIp#8g%uL�ػ�����n[%�Àr�LT7�-��+�3�ϲ A��� ���_I5�^2~�����~0�:���d��N`��a���R�$l��BM��t^�}�F��	��t��逑=�!��ϬZs�fyh���SO%BM�'���:��3��������ł:~w �����so��dk�ӑe���"�4l��B-�ug��ե�|�H��¬D�﫣"���^�>�VQ`�	�`�M����kX\챹Ӳ�/�de� ����50��B���_���<c1���HԄm��(wO���������Z���C�bA������q��$ْо�r?�,N9$���(�H�`_�����ԅ���ղ�7��-�ku�X�h_��v�8�z��9$bDt}8�$�Ə��{�۶q��w;I�nb0�X��J���
��jU���e�����l
���/�*ṵhE��T_/OO���A��!��>S�*w)T�v:�>ǡ���膖�4�`�� �1:�4혻��vZ���f);0���'n����4n!�\��I�e��N�ӷ�I�9����8�A��5��h��i\s�М5n�HH���=���3��i�q����5hn訩##������ti*@��ϵUÁ���M	���^3`�Vt����l��a�et�~cE�ɣ���Ѩ��8�m��_n�!�f�����66���B�e0��򍚚�>z���+�&�	㐷_���J�3��۝S��F����m���o3F/�y��v$��?n9��
teC�T� TϻA`K�Mo��'f����q�(����g��'�eע�'����nQ}�&NY�LT��K^P�/*ŏ�X��xr��|5h!䡛)�祈6��`�R��Z5p�2�O�ƞ��}���pH����E�	�kS���y�����3��8I��W��,٩��Q��$_�$a�?6�@*;��q����p�뤍3�7�i;��ʈC�G��q+q|�D-���r���g�:	��ɳsdd~{T�;�=E���xC�u���J����xJ��%M���8��mt����2�0�#g9/q��O�TgiRf\��+I{X���Oл�W��)�W��EZ��/"V���C�?�e
�ST��[aN�@����+;d�*?��!Gz���N&"*�����
�fL����G�T��9��h�0��0E|�����g�&�b1'N?�5����<wA#��\�؏f���	|�z~���֢t
�'xSP�����	�@(�{zn�#L>�s�����Au�%V���Z�Xi�_�6�tX��a�{3�W�k��#&{=8?�q�z>�(�Se�a�,���pO�겙�����)��|��$�mhh��L���o���K�I`p�~=��.���r5dQ�����e�������V���^��0��e�ٳI���msdIx~
[ڣ��elf��2����J�C��W]����.�B�ĉ|���b� �Kw,�"/��GjY�u�@!���]A5e(z�����h�y�[H⒒A�$��n?�=
x�T�P���z\'5L��w�d��q�ɵ��F���Q��#���5�A^���a�omV�b����י��|�%Lx*�8���ZyS2�׃��Sll��""Y�dB�XLe��N�w8Y��e��Jz�;K��J�)O�]�1�fp5�~,���<��t�w5>�%�:)
Sp�'c��4r��b};偓���ՕiN�s���n^�G��`��C�i��frvO�u_�
��k�ߧC����_8�7���f|9	�1�X�`Wg+�h�oY��5ܗ-@;6����r��17�d#N��K��M�n���%uI��&iCҩ��M3]\�<_j/+��!I�*�1~�&h�lJg�=,��}�o����y��6"q>p�lY�=�>}!�d��K<���KYX�}���,Q�?Рă���3�T�!��n���p�~4�뼨��mm�5T/Dq2�(
gl���>,���:O�������~=ra{h caw�@�wp���-��P`��G��jp�}���U&��F��ɫA�T���m� ��U��eD&��Yc��zY�la	���o���F�	���a�@
.�B|J̶Ꮀb�6+�\��Je��s��H �{v�b�$�;wA�d8�3���;o��H��
�h�>F`k-5�lBi���\ͮy���h�e�G�%h�����sz{�W�����uE�=�����X\ iv��t+o�t^�k���XF��P9���*%�f ��]Bb)��x��R� ���Qu"��G� ��9�떖��_��%1����|W��V��='�s���D��"	��V����U}����*J8�����"�����52:G� �V��ǻ���-{)�N|���Uv�nM�tk���>��,�M;��������h�r�}p�+n�h����.݀��
;k�� ��Y}����x7Q�C����*g��>Oõ�Ժ(}~�}7L���Yj-��w� ���+�K��ҭ�-��7�֤�M߲�2
�a�5�^]�p#M�>�A@��)�/�ߋ�YJ�=i��h� u0�i'1�Y^ڗB'����`����!}#ZTzO�&B6A�<?���;��m�q����%0��s��ixۘ2�)<�_ER�GtY�.���9n2� ��}GM��M��AtU�ј����E*��I_$n*h��J�&���Ć�8
���ک���3#��8�:��X�=*{��}� A���+��^Ŝ�0�,��5���B3��C$�z�|��+��Qs�)��65�Bü�	yVC��U��fd��4��i(��B�덓+��0�����-<�p����$w$�v�a���$un�R�Og�u)�@����wq���wݡt �>>LS��8���
�DK��C��fq���j.��'d������VB�E���'�����\
hy���ҁ�阑v�"sQ�lL��%aA}�Ń�n�oP��l`����Y:��� �3��52���+��?�ź3ú
$��4�8���*ճᚓ��e��o�h���h!z�"�pD]�����(�֮AV�î��X����:h���܃�U.?(vm4��N���jϨ���Z�,uc�T܍¥�/�Bq����x����
�6Ot�p���Ѣ$SGJ�8�~e�&7���A��.i�T����ئ��rK��F��jK�&��B��<��u����$� ���#�\R8(M�����zv [�G��T_J�g���us���~c
���iuuy{�ͷ�~�c˱���Ĺ�ۀQ����"u�&z��*���l=�ٛ��� �lE��:J��҉=����Q��v�<,oF�D����L��� ��QB�x[�%��$�3�Gm�����d�O�]X�]X��$_ziRN�s�P!Á9�g#�
��m��oBhW;��(G5���y����D7���ٱ���WY���)���NcF- �br�d33}��9�c���+0O'�@����L�f=��A/���mw���ӑ�/ڠ�X}�7c�K%��Y���;B3��I�d��>�	��M���+=���썐��P(�����$9�b�U)vj�:(�kk >Ro�˝x[ęS۸)Ю�9����9M�4A�vL7��@�~!���%;�DHr�"H�r�œW�����$��L)k��.��Z�/����;h���i��殓��Y_��pZ!��kL�:�UR��BF���,Fr�-'{����C�A�ez�$S����<�豦����YS���Յ�=o��8?�)���^0&�����Y���������@�����έX�uU��#���v�#�!7+�}��Ө��j[�Q����>#�_Ϊ�����W*��+�0JDGʣ����WR� X��PD�L4�qdˈ��뾔�Dn1�-�m���~::�l�ȡ0:j:j�:f����پzn��jY�H=�.-"��MM7�@���+��̧s_2�h5U�f��W8�\1����;íEX;��:�~���������{4,��}�$���%�lP3��gf\{t��Ma��2Ԏuqj���l����58L����^Vt���u�
j���նRk"3��Oܢfq����]IL������t�﩮��u��
fxW���jK�u��}����r�a�w��X��ߏA_�i$�Av��Kxc/YK��M� ��%r�z��Ê�,�8���Qs�� ߟ�]"���;8�r�������N8ʐ��[�U��(�ة1�Oa����2g:�% �.\-�p�=�ږ� ,kV��X)Y������m����T�n#�����4�t��Z%TCO��-}7�X�+�j�ΰd� %�7�@�t�X�`V�To�;U�YN�v[�j;@g��n���&�$qk%S�1+5j��!R�2�_Y�tZ�=Lݷ��𚽪��!f��J,�o��xb���s���yU��w�şV���%dU�m��O�]���m��^�is�R�mB �����Sbe"�9�˱��F�.S������m�C3X��LT���٤�EN�k�^�p�JĂ���	D�1�A��9f�T)Y>}B�LT@��9��T@P���߅������+S:T�'���o��