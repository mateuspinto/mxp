XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��\�@���)+��M�vkd$�g["H����Y$��҄�Ј�3�p�p�n6ko��we��АJ�D���.,�Q�ˡ�����Fφ���7�n�;�xå�F�2�=�Z�oo%�C�����T�$��0�PE����A�*���
���܏�l�ٔ�ϸ����BNo=��� �C�}Bc��Ck��a˓{N4dk�A���-��#zcâ'��XQΤ�.�N�gp�:c�JI<�p�?��T�g�s�W��
�4�4��D����ơ��;*M�v���"�	�.�C �oc)'��ḀC?d�P ��1����3/DA[��9of��M��bY2|*$�!�d��t�O����Kw�~\\��,���ݮ�_,��+ 9�ݾG��t�Ձ��0���vՐn3���sΟfJwJ�M�L��i����[���(�xr�XDAN���W�R��3����/��bi�������T6���'E}G$�P?P�%�- mj5�F��қ�G����?�161�
���@�?���/,ʝ{$]h���] �̧�N!0���;u$奾�_E��[���P��{��M]X�l������YF��{��~ȶ��I1w�~A�j5��4hT�s�Ј�C�|���l�x�� �3GGf��u��-2���Xj�]�(Eha�r�-P�A�c$�_���r���%�)��Yd�8�{'m��K�T2�v��! ��5�~Y[K�	:���R*��&�OӟY7�JB�+`��I�q��1���9*�_�r
<XlxVHYEB     400     1d0�^�pQ�kP�\w�8d؈쯪��v�P��:��S ��*O<"�h|��SQ7y�G����:!��������%��B���'�<��1�ֈ��h���:�X'������M�FsA裡8?�C ͣ�Sԓ4_�2�H�-�y�N�BQ�?�E8��1�1 ���7���ƶ��#����/�(}4"!�m��I�P����"�����}����&��Ln�`�������F��i$P��?&+����U_C�z�
p`l�u��5�����/`�UEI��?O(-6�L��qT�~:j�w4��X9������0����V�#(I�q&��t@x#��G��5>�Vcvٓk;=L�/ʪ8��>��i�v�GC��bI��  ��k��TXTcW^}u�H�=i�/Q���= ��1���T���S�
^#� �K���GX]��l��ZG�6s� �/%���*/K+?(
7<XlxVHYEB     400     140��Ls��X&Ϗ��fκ����S�r�XkX�g�o}����0�,�S1�d�̫�`!�s�<��-���e@�x�)z�E���oF�("P���-��C��Y ��/R��1 �'��\P��C� n���p�����B�>��%>d_Ǜ����kx�!��l �`��"~�*�
x3
��� ���m��/�=�%~������LU��i�*S뼀�����rGݑ�m̿VH��>C0|鹐M����)� ?T�{�4�Lb܂0�2��}'����a�5���W膲����C73�����'���DĊ�?7��XlxVHYEB     400     170�@"��E��1��<�\������"T9�#8c�Ҏ.�5���uv���{�GM�{����<��Mu͊$�E�6��su2��XK��~�Po�3�1��a��P5AT��ǽ�"K>E(��8��i�(%<=]�*-���i� ��`���-�D�AX�``������?Z���	�.��}�ңQ)�����/�b�����
��v����E��NuV~�|�~q�;��GZ�����XHAiO�v`��Gh��{&���څ���r�3J�DS�f��d�B��M1�@и>i.]A(谦g���xR#�	���_�^>����h�>��ʖ���u�J��JQzF-�no�"R5E�]m�3��Z�&���S7I!uuXlxVHYEB     400     140:R����vs����#��c�o�m6�l��_��X�p@�"��pэ*���:0AUP�_���*0�!�I���/��~���}HYe/3�R�Hk!;�v��M8�[z3��@��~���C���#��V�F~�/[k��W�t�Zk�� XH
��v���hV)�%5P�H|
�¶'�k�l���5�{��t>c���vz�0�z��-�H{3���DA��I)�{�7{�l��B_F��֒GKZ0?<r}�}%Ur��jh��u~"A��f�ۯgxvcA?uO�m|�����ҫk��/d�颌�b�*I��	� 2����\�C��4�XlxVHYEB     400     110���[�١��\��n��.*c-❧gvX�U�)���.����=�S�˻�`���kQ@[���~$�}�և"?�p�6	��2M4=C
��-�Nd��$>H����Q��{�I���\H\!�H�;0a�Nmo���'=N{]��D��{9�zor�1��u�SB̰`��d]]���;�0�'��m�d�����"��N��P5J\��lShF��o̤k���������E1��0��1���W�"�sb��E�{�h��	�陀�|�M���,�oA�XlxVHYEB     400     120B��}��'����~������xJ����HQ#+���\a�`�Q������[�D��U�IE��a}Yy^�?:}/9�~US��,���^ 
��s��q>K:�����t@���lp����[�7n
e�9h�0�!H�J�/�W+
1;e�XL���J�)�Ii�Jמ�D��,&E1.�e� /��{���:o��'�����/롐�x��f�<�.R׆HN�<.�8hn?]?v��~=E-n:��_�LI,B�lb�ק\y�a�u�_B�3�	�\�H�x��UX�XlxVHYEB     400     140�2
Z���.gҗ���(��Gn�>S+���g$���Ȃ�^i���=H��C,�-[��J�� G��dR�?F���X$�8�SX�VaO�?�I-��L%n��SP��'^9�����m�m&z��M!����$��#:jS۳Qh����QJ<�@�jQ}��� ?	�	$ק��^FD�D�v7PW��m6PE���ܒK���Ô��ŘG����l#�/�9��>k5ph�7�y]�Nyp��[FDO<җXEƴ��CP6����;N�͓A[��j ��\ ӌ/vQmE�����]�,z
Zt���w��PA��ϦYiXlxVHYEB     400     150�~[���Q�R���������������Lί�R�gk�4��
�h��nȹ�j���D!��DԚ3ƭ��x�IKJ>�W�E��?�3�ş��2㗁���;�.[��
Y�l|���4rQ�b�
`L+e��G*�ߗ{�d�梁��������Ls��G5w��c����31��{1��Ed2a�u|�!k֘��h�Jk�Wޠ�3���G�ү�C8U�ElF��~��d5����$�P"R�}i���eѸU�E���Z�P��8b0�F&pRA�>,X[㷦(��%.w���ҽ��M�>�/xK*es5�-o&/�gߨ�����X�XlxVHYEB     400     140͑�]Z�u��I� 
W�h�A݁ώ��ri�H=��{x??d߻>�q���W�,;�{�"N������h�4R�%�X�`�i\�Y�*^� ���c`B�=�|�3u  s߇��b	��~`9����ݸp�P{~�lk�P^��>n��+D܆��1>(P�kw�Q� ���4�-5���O���#���Q�β+'ι�*ς����h��\s�4wzz�N�� ��,C����fMO9�]����'-��E�����ۅh��,"����1�:P`jր�X��L��2v�^�k�|ȕ�X�*�J��K�vxu��d<�V�XlxVHYEB     400     100R�OX(�~ե�aRuNRE�|,U�A��XE��9f�&�U����&�6�	��&Kg�+^��dM6?�S�[��j�b}AFe��N#.|�5>�6�8mH�S`��%�)��4�h�AK҉����#��A�[�{�K$����~.Dbr�P蚖��	��MG��d&���)^u؜o�l�/6�u��G�b��HK'z��.~m����>m
W� fi M�`�hڕ�p[�y��Bx8�	�w�%"�U�>�x'�XlxVHYEB     400      e0��c��^���`����2�N����'I��	*N�����l�s��¼�$��D�8b@��a�e���}�D��y(͘��a ��A��5��)�B��e��#5�P�,�S�7�4w�~����KDB�{�q��9g�џ��A����O v���y"��C{�qj�St�5p����TB��(�c�"T��=�220�]�Be)��_��ሰ��^���1�XlxVHYEB     400      e0*���E�IY�](����uX�b�{B �
�ໃ����{�\�[��%�~^�paƘ���4skN� 9=guwo�a]�fl��N�:�T՘NX���HE߿6����4Ji,�t�ƥA�*H��Z��>_�ت&IՐѺ:綞�N�[n�v�Nǚ���kmjz�v��y@2�<)���ٚ�-�.��N0ݬ������7�>�OΎ�!��Ҍ���F>��8�
�:�Q҆�XlxVHYEB     400      e0��E^�5�"�9�Ӑ�L�����1��Mp��������#� �̺��	�k��G;�g�%�FU=�mpĔʙ� [$��b���<1FSqӝ�3zU��U����Θw�(�A(7H����}9���:��g[�$Y6N1��*k����Úтs���C*�| ZMB���w�#��,�H���q"?c�3x����$bM��b�Y]]��g��Hi�}CXlxVHYEB     400      e0"���is��*=����s�ج��#�Ph�l�Qn'TŠ��-�~�����t�oIp)�8l.T^��f�?�Ʃ��͛�4Y��z��� ���߿6��7<������D�c�o��V͆EA�,���%p��h#�O�4l�cX�8J�^���P������C�HE�]�a������Jd�$�%��A��֮:�wUj��$퐋)m�B�v�թ;�XlxVHYEB     400      e0�X�3�y�#k��契����pA<p���-�i<X�\�:������?W���W�
��d��G->XS0lm@�:�E�dM�Xo��;w'���{��Lx�`1���y�>'gʻ��g)yuA��?&�k��:bW�~?o���
�j�=�?��+�(�w�9�ˡn/�v���Rw"m��H����̒��ܶ��UZMw޼���~�O*\S^��u�F���O	\�KXlxVHYEB     400      e0ν�B��8m��@9�V��ktv�ޫ���D��+��м;�g�A�r��T�K��
Y��$i����ȟ�T�9���w5(�ߨ7B�Y��/���a5�P;fh�ak��n,V!؈+�7�i�<2�Jh��1]]D�-#]���/�˲c��k��i�Z�� I.~2�/@�E�����ے�Rt�9rP���"_��f;3�ߥ���٬����R�c��@�XlxVHYEB     400     1c0:�G�����&��C���Qp{~W"ۗ���_:;S��}fK-/%�o^5�S��;(������io��߰���UB�HCЭ�"��%Ej~:�
̚IAR�XY}�h7/��y)z(Q�1Lqh='��m�[}pܠ�)-��~bN�e"�aZۜ�d����)��_(s�Q׈e���5�N�<�V6���t�ʍ�g�8��rr��d�1T���At�3�P�_3�dV�?���~k%�U\�r�QF��V%^b�v�Tzcb�o=�G�j�Ƽ�%o`0��G�e�~=���é�<.	:[m'�A]�^��p�.�(��q��� �Afi�T�GƦ�NdH�D�k�tp�r�޻q��:͜�I��o�pzsZ:K��;Ȥ����#���ad�є���L�	��0�|N]����W-δ�FR3"]M�Ay�n@$��}[l�T&Wm�Y%|+AXlxVHYEB     400     130�l��r<��t�I��B./V
Ǘ���L�8���� ��&�^b��5eW���J�ډx�Ჽ�nJ�,�&��Y ����y7��dL7��!�z���Gd��.��ݥu m���(���!�
��������C3hz���./a�{��x��B��/+]��E��@Wee��4t�ȁ8e�mjh�l��2��zSؐ1X%�emS�6�����(��r���X�x'"�5m�d`�� v�5�5�Y��F!�v�Tm$9� L4.ɠ�&��(X�SC��{:l��t�; ��NM���F~AҒ!jXlxVHYEB     400     100x=�B���h/IF6[MAU�9���%X,�b�yi�,�y�m�d��o"j����]�3Ą�S�I{��-�8av_��Rxt�x�؁�|��b�Y��<���1}ɕ��V5�|\����R��Vu2+�b�ɚc��1��5Y��#��s5�����O�J�nb��]z��;���n�A���=]�c���0p����L!;4Ԛ`>-���a�4�^��q�?����q)s��$�1�|	�;�R�d�b-�XlxVHYEB     400      f0��@�MfWf
t�7�8%��b�u_ɵ{7���&�I�<d(@���, �v&=��|�ղ 7�����*�G�D�J��TX�$!{�Q ܩ�أ��\g����&d��b��N�cc�v��%�ZB�JX����RŃ`����o����1��͖�G���w"3J���+�Y��mS�G�K=���� ��U�[z����jTڦx��P��G�o��M���ӐR�A�;���gXlxVHYEB     400     140�_|�����P6���UR�g�������LT�-���k���z��^�v}&�԰'d�A�}v�l�nT�/Me�eb�p�P��5X��1*�F	�P���FM��T�O�(;�%�ZhĢ�����k��DX#��o��	������X)�Ҵq�xm���D7�����j��)���n�-�3�H~��y�aj�r��w?w�Z*N~Vd0�ݑ�c�@[LHp������ ��?c��h����� v�K��qEq���(Y��o�g	��(�.�_�����N���BXt �l
Uo$촱L��wq�ܤFaacj��/�#��Bx�4r�XlxVHYEB     400     150��{e�6��ǌ�����ԤeP�;���5$j~;p0}���٭(����M���Qq�j��fc3�\����s
[A���0X9���M�{VMa�@o��@XU��MQ�A�]|��dQ�	v7,xT�ن�����$h���{��ry�C��A\^a�/��!ϙ]��蹒�MЪ�U��R�	�g�F��������L���!�_�vg��~��'�b���/K��Y���_��G��v0�Ȕ�Rd�ՓĬaљ.�y�(H&J�U��!�*���бn8�&��o���2Y�[1+,q��97��j
�TA�/H+_Ӣ�1�~.�+�ɐ��i
؄�XlxVHYEB     400     170��N�y����tJY��b���{C�?������}c|����n'�{��L܄N��R����jCju�	j�M"`�gQf��<��Ձk�<���lTF����]�٫Mc9�!U*�0)��"z�S�3��H�q��@�+����?�'����%"��EG*>J��oF��'y{>6�[��bG[s�	D,ײ.�"?=�Sh 5-_���AT�G��'z�Q_��~i��~��-�z�l�z�� O_��1��"��I�5;��NT�!wj�sYv�=�a�͟�19K����D��0�3�23�D�Q��Jx}mZ�V���URq��:g9�7"e��H�-W̫bA
 %�au$"�6S+����2����XlxVHYEB     400     160��ɛ��c=TM�7���w��g���urS�S{��o��M~j�
?u-��0;3^�� %��1�RLE�[�bÄ�%�հv6.�e���Ω�|�S0��oǖ�=Ro!�Z�������V��ɚ�8 ���Z[Ė��I��
SrN@(]G��W[)v]'���4!_d�\��qHz�6,��F��G��E��E�Mb܄��a8�q6�"`��5M|Z�����q�Y�f�Jk��[E�8�O�ӏ�U�٫G�=!�%����ۈ��*���h]	`�
��'�9�����9WO(w����
��)��` n�պT�@�Z�~��%�XlxVHYEB     400     180�{� ~�MH)�,��ܟ05{"����@Un�茙��e��\9�2u�0���,mh$<�����L @�j|<��t�$[��μ?3�p8�^N\�:��Bz�kb��a�#>ί0����4��Y���埣�"M�92�����V/uVL|H(G�=�F���J��J�4�e�o'�~C�!�1쬅
�ɷgo���5]�v"�W������"f0�:[��.�,�4�6>��S��5���>>�&�!K��-�P� ���_�����ZE1�sJ]�W��4����n5�$K��ÉÐ�y�yjmj�s��U{>���,�(�J�Ec�j�X)��kC4x�vj��7Ç�M�m�U������Bl0��cG��cN�k?�إv��_[�|�XlxVHYEB     400     100�u���~b��`�#(݀c<�U�ڔ����,U�z�,4�XB�C��pRi���M6��Zﲲ
�0�[,B���i>�!O�jzs�vjW-����/"^�l��EE�-��R�"z����_�\[�&�7;�u��yj��'@����X�/Թ�s�8����Ea���r?�*�k����E"�t=�%޵�x�[Oy�_ǱB��E�Td��}5����� i� �H�5�����a�=���x��1pER�Y7KHXlxVHYEB     400     160y�ۮ��ܡ�"<>n�13�2c�:���g$�AۜX��\�:!=M�WӼr�8��|���"ݪ��	�)����c��\|�z�&Â�E>t�]�T �Rg�)F>����Z�$ד2�|lx���_���@�*����S^DVҮ?����$�sR�*s;�?����HKP,ĕN�j5Yߑ*��ƴ��?�3Ķb4�}�Q�����tG�b=>��l��.�QJ��7�����{���j0�J�~���x�b�w�\�ԙD����܌����8V 5�e�r���J�@豸�T��W���@�%U��Q]���&x5��֏��!��7޿;6]����;X!���_/�G��@XlxVHYEB     400     160����>�OyE� y3b�ݍ/��͜ezM�\�n�E��ֈ� �S88�9��!�+W�'R$�AY�.���N3�jv���iX�$�`-����GqZ����y
�mRt�F>�J�-��s��\�Б�=������^;-�I�%Wz�Nq\Ywu�GL��~;��W�������&�.6����s�c2W�$�U��,('H:X��7�{���-_�PBe^����G
�xĽ�]n��%��|����1�w��|tT/R��؂ya*I1���6�nXf2���)Pj���b�b��w���w�/=/$��lE��.��q�_���,tO�Z���b��8�>&�u��C͙�&n��zGXlxVHYEB     400     140ֆ懴�э}t�?J%���6��0��m�-�Ju�Yoc�0��f]����V���5Ԯ�x�A�g���^e������:�f4�Ѓ^�Č*~���g���]5��4�Ř���lbZP6�O5�0"��>�~u>F#�ć���v�CK[�v��I�=~��/�������^>e�7:�ea~к��o���ʖϪ���S�aQ��V��+'�jtӉ��ݜAb�I{y�̣��i��Fl��3�^�����u��I��{w�1V`�}ǔw������g�GזS�[��F�O�/���"�f�K���!ׄ=3�yaC��j�M'�PXlxVHYEB     400     180>���
�9�Lpv�V�s�v�>�@)�m�n�9P^/]�2�3���v��N��%�)�L�{�#����q��(.���Z�%��h��Ɍ�8��N��!�������Q�&gr��PBp�y�<E�I2�a���,�jع��p�U���uR��,�E�i7���_���.e2p���|=�}�S�/-�^�I3�����%%�u8���e�&�iڊ��@��ާ�q��+:�q��ROt�����9�1�ټ��T)Q 	:� ��W�ݸ�l�N�wp)6�7�PԵ�6�� 9�C�%$~b]�9��0�`lv�=��[���(T$^^f�����,�c�L��͹��A(���O�H���;���������y�'�XlxVHYEB     400     140H>^茥�� W[��+/{��@���'UÚHe��{��l��>c�S����^ͧ*��6;��S�.�"L�;�Ku8���9�(������>���zE��܅���2AnY��iw�����n���P�]K�[�h�"�ڱ.�"�sM��!m�<�+����~��e���:�R���j)�%�t���Tq��Hf���=�F����'߲��������唜�]sdȷ��~֢����st.���5P#v3�o���S�~!�am5�X��$�X�s��id/���
ZƧ��+���EÌ�n��4$��qp�ſh;�6XlxVHYEB     400     140_�8�ڻX?�!��M|�3�j�oy��x%�rpK�e+y%%�^��b�	�e^~�$����N����AE�p��1YL����g��g���� �B��ʍ�?�/Ex�+�0'(�ׇ�܌z㢼6X����s�<�N��Sk�}G��Ez�s�1	��[��q���nᯅ�̵A�E��m>)F(O5�$i�s�MS�P�E3����B�u�pQ���Y�x13�W�Mt�k *���8��1Ҫ����/�W�^.�kȁ҆o�9QY��uӕ��Ͳ�,���렟ܫ�rh�8�>v�B����o̿�	�GE#.�6���+v
��^�OTXlxVHYEB     400     1305��Ю�t?L����:}W��>����fG'@�1%����\��Q]5Wt�G���\�+cy�p�lj�Ɗ��I�]��#�H��5Xk�9���PC���ߌ'��4�_<��7I�5����&\W*nE�,�Ʒ:]~�q���2�%�{h��s*��\l:շƭp����>H2�~���}�dF�.�S.�g���I�a�]{4N�6��w������ڃ�G}���6y��e:��{�&蠚��5k[bb$�k/�W��b4��&I\�`�; �Wt�,�M����=w��)y^N�XlxVHYEB     400     170��ٙ ̯u�+�%UD	��8��K�Tw`M�t}��O��#�b9|�6�'}�ȳ��U�5(�����z8,;b�'�R���җ�HO� ��ݜw�$ů��\�fI^���_\S����V�#����~Ǆ��Uw=j���ɪ�
���wv^�sT��OC��d)^b�I�C�k=2�&��*va>DUw��j��?�1rt:.p(�3��$�3p��:{�7b�v����H�
��o��6���a�����F�t~��^3[���J�^c�B��X�_�ꗑ�@�길�#|uf��.)|�C�� �Bֺ��:k+�ф�}B_����3�;q���K��l(�L���@�FmW�7m�XlxVHYEB     400     170uO?��n������r��`8�-��׳���i:��'F@Va�{���2ƒ�����~����j�+�Y�	$l!Kl>���N���ݢ����Q�b7!l�&���>FI��
���^�id�%�ǔst��?xO�<ğ��22���Z4�4�J2U�8?_������!�4\(c�B�CR�\B�u�b�Z �����J4��i,P��,����YY�M��t���Ys<��g��`itfS��v���Y'[�m���O�FG��gY^.����������^��c`r����/b+��Ћj�6���8ӊShI�	��z���T�Y�l��b�H�˒���1i�r��B1�o�+f!���^���&/e��)����XlxVHYEB     400     190�-Oz9�@n��M����ǛA`'�>C�(���d<�@/K�q�7=K�����x�`�gI��V�3��Ei���kc}g� /���� �`?	QO]A�;�Z��Vfo�_��@���X߅<Mnqu��5K��������+�d�)�<�����y>g��N����l�����Χ���G����GB�8�����S�b2���\�x�����_Vj��GLם�@G�`F����[�ׅv^�,��X��Bm�7�=�;D1��T�����y;���x _;k�O�p酕����߂�M��g������D ��Й	��VWy�2:l�mʓ�a������ �}|�J�!fyFv�wMw>'N�q�Z	��iЙ�����>=���c1��=���44$���*�-��XlxVHYEB     400     150� Z Ź�j�cS�o�I�O\#>M�ϐ�&�j��&���ڣ^|��=p��j�����P#��iI�U;�X���?�iw�g��?l�_FT�r+U����Ot/��&�}rѣ�FQ�uk]I�m�*��|h�q���
�g�j���w3Ҵ	�*�-��&+�CY{A6,�g(�y[�~٠�)�T#�/ ���r@�7��/D���0sf�g��u���83����[K+��p ~�0�!R���X�����8���647�_����}�r=4�=-�8&mr2�"JftXS�pPA��v|k���)C�����{��L�#!ݟfN��4�8s>XlxVHYEB     400     150DQflr��������X*��A ͅ��LOC%�3eg��y)sA�	�+��Z��+d�8��/&\��OI^�\�q�Gg��ϼ�<<��h��!��Zk�R�|�i�`]̜.�iV��~{_�ք	��ð,-���L��ͩ[\3�����~/IZ3;PH�c���Ӻ���%�0�/�଑wV�b�4�����V�z	�O6�H>g�H�Pr/���,A�cO%�LU42��v��0Ÿ���e�ke�)��P�zg�1}駞�-%�ʓ�T5K���_�w�ch@'^�D�S��)������Z'�V|
�s��>�L�X:H�t>XlxVHYEB     400     160;Z�5��BA#4JP��훬��Q��	�@�v�t��"E��	�T�6ӹ3;M<s�c�9
+[+�I�-L�c��^b�2�g�'�k_j��S�
я=PM�RW,�U��1�PV�B�BXW�<��h?v�9O�?����*i(Z�2�<K�'M��KS��R�w�c4���� ��ug٦�,�g��7M}�C7���Y#�'�[2�\k��u@O����ej������%����1GF�>��|��E��U�Bz͉�,3_<����������~�0z=�+W9=Bρ����=��:���K8o�Ԗ.�XbL�zڧ����
�e��n�;����Ng��|4۟C����XlxVHYEB     400     140��|0�U�~���;:/��Eq$�����Ã�i�a���<��(Z��P�n3�� �4�E7ًis��������;��7��t]_A�V�o����T���	�{��V�"5^\b���Gi�UP/��&���>����������7;x�C�|���OJS[������F�tZ�_`t%C�c(��7B6�.W'2A�5wz༒�37��M�=�A4z}@�[9�MA*C�yI���i�~���\���lN�W��~����R�sQ��H	 =,2'8N;����`^G5�@��n$�'�.�Brá�U��T���.:�XlxVHYEB     400     170�I��iT�G�/����8�j��@�^�dyv0��I��3�o�kתt9vr�o��J�|�m����צ�gC�Μ�g#�D��]R 
i��I��&�J#�iI25_TcE�X����:.69��٥t:�k��7+8v��"�/�>���:��)?Gĕ�������h�+?J��K*��V��-ԢǠ�8�oj70yz��*��zE�r��WCm��)6��2�ig̇H��BK��8��
�\�I1|�u��,�Z�ގ��_�I�Z�	-���W'L�0���{��j�Q�Y�����`�ְ�_D��k�O��#���ee{�
�5j�%z���I֔e	t�������˄/��p ~0�+OXlxVHYEB     400     150#�-�&��~9�z?���Vc��Y ��.�-t9(�(���i�a�aX�햳)i��<����˶����/�:�F���Y�h@;&]𵼦�������ه�h��>k�;��v�܎;'�jX���؍'�P/L�_*�ZXH�:�=~c�J�#,��D�'� �������O�����_\pim�þ\�N��b���|�����K*A��5�J{��Y��6�����1b2��u�7c����+~1+LL?r������>��a���O��h(O�������_jgqX���5Q/ e�4Xٖh���U��_�AЏo���e�~���P�Ć ��XlxVHYEB     400     110F�\5M*��'�������EoQt 	w��ږ�e���Õ���wpv
%��xH��=x��� 2�e�ٓe���5jXL/�N�Q�SL�1ͽT�S5��}H$�F�g}�r�74�B�b��<����r i��O��t�K#u����\h�U����r�^E�oF��C��Ƕ��pIÐNS�J��K	��u�uh;����܅cYJVV��E�� 	��6|>�cZ*�ʍ�Ks|)� ֲ+�� �M蔆K�����aj*h�c�֕�<XlxVHYEB     400     150&'���I̜K���N%e����c2 T 
�|���R��A���^O�y̎oһ�݈�͊�`H�2羧�i���LדQ��[�H�4|�%#1��WI�n�,Y��y��2���9?�� �����G�]��u��ڦ����D��<�+���s�/����|���<�4��M��Z�l0TY�l��.���Y����Ln�'�3| L��iwS<�
_%o���ӨԣQ��]�5y �[�mHSNC�5��^q{�Pbu��8���nTH�Clf�Ѣ��.��/K1�.�+����~X,��M��s����1�>SG;�bg؋�Ȩ����.�\m�XlxVHYEB     400     1a0�)wd��80�JB9�Q�]��w'��*�;Χg�aR���u8
҉f�	�_5���h�{��dzX����~ľQ���5�W��x��d2�}�↻Zc#IbpX�ż��O����*�m6p֠�=�2&3���}�|DCOqc���6�2�����g��炏K��ͦMaT�,C��r~�eVn��p�0���{�����a�_������q�36�z��S�H�DK�$�z@�v���5V�HTO-�d�y����f��O�p5�F�j&���i����5X��h�@�mpF��_�|@eM;ܔ��|@/Nx	���k�P�`�b�R���]�(��Ԟ4q@f߰�<j�:�Ġ�Sj����������������J{F����ٹ��hZ7K((%P�{f�"JXlxVHYEB     400     130dr�OZ<jY���z�K��;Rף�z��$���(����������S)��~T�6�#_�GQ��1�Px�x��13�����]?�8+ a`�v��[�k���؂g�A�\q�rN�ݚV1�Qs�$���X؈{��S��o����<B����2�xV�^�F���p;uW�:Ye9�=��#j���S���W}�* @�Y���*/��$�%ɳMO�< ��HߍeDt��$9?H\���	�h�õ�7���R��dC�(��XP�t*�DO4#���y����@�a�A��:����$?=.�գ�������XlxVHYEB     400     120�,��#?7��5��~�u���ń�G��2�VsR&s2�
�MɧY6�p�V� x
���制���_9+�/c�2�>9�a�홻#/ȱ��I�'8��ZpoD��0�v�̋�?Jwg0*l+>l�
�.(0*V�x`�5K�Ѷ�W8�	|8�ɏT��-M�ϣR�u�N��3�{���fη�U�V�\�L��u^��
�I�qa=n��
���*��p-��m%r�R]��1\�AbHϼ�B�j�<ƈ���Ou�0~�<�m���W��������<[}S���=Zm�<t�C�XlxVHYEB     400     170�c�R�\�vK^��������E1����57aķ>^-<�h��S>�C�RR��,�wI?E��]���`�+����T-��$�oO�1�Y6�^�nf�6��6 �"�>DBS>�C�l�x��,n?᷉a��(��@��Fbn_s�i���YO��&o�P;/Ƙ�C �jd��|}�H�j�~k��^��Q��p?UPJ�B��DĹ�{~���G���Mk��2'��[�m�w����B�u��;�����Z���zw�l��C���z0�ф�܍����e��9���SiR}j�$l����+_M,��sc���7DBAY`p4�w*R�[�rH��q�s>��,i��'!��kDִ��̤����w
�w�XlxVHYEB     400     160��r�3��h,5@a
�e <�$.��->Q�&2P)ϊb��%�~�3\�$�D��3����z���z��sd�2�65b�׫ ���;�QR?�1�B�Ѝ�����,j�"N�C��{������6�R)��J����&z�nC���";S0�<h��^�/ ȂA����Qy�|1J�z#��A��.|3���k cD�oH��̪�ӭ�iO�A�JNu�B62�BjkySw7GP@�{^�^P���["a��&�Ht�F�;�.�g�ܘv?k��*t���^��_l�+�m������,�k��_�Q+*6��Ӕ��lH��q��l-!�%��b��T=�U9P�EXlxVHYEB     206      e0����'����A����5��\f��(�kY<^����i�e�q��It�GR��v���2iA+s�_�t�ᯠ0	�4���d�#��J^Ў2//ׂ��� �	5`����[��X2��4��^v.��S���?��][�.��=��$��ӹ��k
-��R����U��E���:��O>Ft��3k�x+x����X����r��=�����(�>�~!�U