`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3088)
`protect data_block
iyygw1agjObBXyU4WW+5qJk8x+3kHe+pqHt0TR+ljZVelL3V3P3nI28lRpXJ3nGzI7nNTFmVHUbF
hx3Ll1WtFUnTNF4Il3FFf6d3d1mU6BRKXIbpH2HYShHo/dcoGLnNaNUWQJXywZ6zxS3DsxADlhH5
r6yGvl73S4USdDDoaTKy9Q/vl1BFrFw0MiWptaO4dxeGGFmzHr29wk0xjCBhntDgx3AV8YpklQ+H
fGyIK74qwpFdHPVMBgrgjiVZjCS0xcmABWJQR6zRKRHAJy3+6XARkY5T9G6uY/rmB6gNDplmg8dx
rqHFoWfJZBdxNrgRQ0GN+OPCvIw18jVO2b+u0Rl8c9hm3xOwevqXsJL90wNwW5b2OS87KhJEl9k6
M2/CZgX0UPKlEMa/OSERUL0mfFEkH/oe2rxEXC1+PjpubbS6CWuh21/AXjA/XHynhGnw70q8qfKL
4b7WxI2flpkFMQAI/hR6Ecd5rQD8wPEM0Pd3MLxEsKFBT1zkiRzH5HaEXNitywvYX0VZa/gao/cQ
8lG12J9sJvdyuHUVFZW9+afUfGuGjagbvvSDyCtefBtwj4+LU0XfAiSLYxM1cKzmg7r1E097L+cc
j7IUQs/Ow2GorLh9DNBjUTKwj7yixdVyqm8KID6jSh9IQ8Iqc+1klhJXFdQMdUUdqCONJFpH+QMA
FBJzrS6xuie4dY29B6F1lCUwT2wPDFiDffdeC73TNQtiMyUUyAnTmuvCF1YWACV6xJ4YeBGcjOTb
yFoVNCaZOa8r3yGkYlATcT12XNK6kqPKXG5AmQsdSH3dwbj+FqD3hucU/R4gUMxAL7yelPggVEvc
lTQRwMs3J28pP7s+jaCVY8pX/ZTXd3KnYkZIEgzbWXjANG2Vs4Ymga4kWcSYim2zFvXsQQQQC8yK
3YGu94X3oJwh3z/IWgb7jtx4wEHOGwRXYLxxwO+gVJn5L9f/YmUrhKWZhciIisi5jAYHyJGJwSgB
sfhWuS6UJrYtvhhJ4XTFPAFFnuqyI85vVWO3cwdq2xbk2GhftYjUUliVzX4u/eMWeqdBujA4YPAL
VrPXtCS7Pxvrogt/ncG0DB1KPTspjitedRwSVuCOyQhOtip3PGFuk/DnkRx6PhqfP92ZJTybkRl6
0xIzt+nzAqj1aML+1rfSfs4zH4kO/MMBJkHs6zxKvEfOoKRvPxegkPADG2/GZME4yx8AsryoGG4R
Pfz/B6VTN1rNy6XbCBgXXU7jyyWg/qrk9dlyd93KoZjIvDcdFcg5/oEQaKYl43kJM4Mq6j1npMwj
kVsqVLxwgjR6uS42oVCfBEu+oa/ewsK6dVLTnbpu3CT9UeBjRHoc0H8AB9tfUKr9bDlbrAiU4DMt
wowxa4ZzKnW4zjq1K6tCSWDTPGYSRvwYippBEdsMdjb6BZ8Od64TDIf89MnZ43okLM0k1bQPZbVV
ri8DIpCRI+b+kcTk5h41fZDLaH/CMfVpKQbL4PpY0mB1Yk9XEtgOnerfen3HmVZ/e7xaCvzWSv4Z
uZ3ePxjIj8Wraka6yozMr3kgrVC/jMzGeAgMR7VaJz2GF4UZQqbbNVFEd7f4gn2MhKNGh9y5EvE9
Lb9ntVBsjhWy371FD9IGjEHwoy2mxehvLFhb+IcdXabB7QYSXS3Tfp2n9wjeIxEXGhfYJf4ZAqP4
/tVKixBMbjx9Dqr54szED5KWx0ZuTVwmv1r3ZUHo3ZLtEyVUc/2SugHMvK8UavyJyaT/Yld9CLzB
nGNAMovaH/Ix/B+4dqOTyN3fb8Btbjw/XiGyAGjYoPEmpGy3qz4DNjWuBdlD5NLedoRHS7SU8D1f
DazDW5oOyvnQFIj9lbKyC5Wm8ZJHQJ67ATJ+8ldmR8yKrlOph3wC/is9PJojkPXVdYqFIJ92pVue
vfcvdCl6wacH8XUymo75ixWUACVulYfM4gyW/Gzpaxxki4wmFzM3YB2wNAhd/wtzDPkrYKT51UbI
oKtTgrKFxKAD7abVOSj9bmBsVIQNZIU3PhVbbPBBTROguZVv213GvQNrPIzhRB+z0MyFgZYjJwWC
jbsam7uuhZJ8DBNqxeHsgKzHMucMHSYXlpAS7n5jVEmGV1WYW9r0xQpHNh+mHXVfTNneGPuHMWS7
3i/xZnshddkpRMdlbUMdNNJQJ61sP4WIFD6z7ol0CmsNRke0n4qEpuyPY5JvgSFpcX3QnG04Xe2n
yZ5Qp7hbZLZsFyPTxDvE+jPQR+m5uEdVU9MbKrxYh03Vv4bktoz+PL3gyjifNnWdd6Jmyyoq9wpp
ugvjJ0kZ8TGJqDk++KDzB7jwTLMiX1KhJxCm2FM4B424vGXbkOsPKxIj0Ptl/Ck4WC3DRAJQJZBc
/gRmsnjjolpHdqynS20PCeBfu9uln5pK1z9VL3GFGZ8LYwN6C8369SjkAYtJRqdaeQHkMkgVXvdt
e/A5CgHCA4cdxdX11Kg8at9CQkoKLizLiQ5dqocH62WrRYdVPLK2sNe0VhGR231QcYmF1TLrmMdr
qD3G++5P2iTOuE80X42CajWdLZIFFcZT5on5hqTa0BmLuzRHjLoW/3g02Cl25Vt19xvSI9AYTnNP
dhzEqTuS68ZKOhKIdumFY1FGG4SRDhvrpIsfOmlCYPJIQUyZJrfiimJpScDxyAlR3UQisCMbzN+0
0jIKcJE6Dw80BaVVtANu+z4QglVx8ch8Mf9CtyG02UhUGA5DEbz1YbzeLadjYg0cl/mQGq5u6Qbs
WQ5YjshfIRT1mGdq7zq43YqbWqMZxkQMICyAIjvcjUMD9pf0SM1RwSJYOBJbBNW1BsWX17IcRuav
GzeR32j44IfXWTX3ipil2dwBRVx+O/CWoS0RD+vgwWJBsFU6D+ZExXQDnykE9+PEIW4Yk5C+pAL8
VDaUnqJ4Fu5+Vph7ERN8c5+N91zsc3l+L/krOQrh6XG8ouGMKdQMPHksrEvDYZyMvn0OTsQ4Pjq5
ufYa+ntyEvg49YeDt7bYz1poMSHc81f4t4uUiDRxRCfp4xQuwcihgnCJshQnZ0dA8zUIyxyecFng
VjUyw5NBmJZc91pInSW8Gn/h9vwk3WVl4pK9MBQ3Q0CKTmq2lH8sSLQzHSsv5aFcVE4Xapmnp7Wd
EKc1N8rVvZFO/yEafCU3uy3bc2Y+T8sFRzsdPGtjVO5dhfMnt6zybYz9l2GH7n8+EGtKo9D7ca/j
+P3FsIiXAUMBjS7BY/03cm9FB4mpovvJX6KFIJHA3xk0R8oBCZBADof1ADfsoZWa0PNqJnr1MXz9
kGO5uuz95zbP1CeseZMDDcdI1hizZE6jjpEODqkuI9kUmSX6UQo5k/9XLWaAWeVOUx2w0ezPg8dY
NHX0zRhm3vNXn2E307TqLTDpvMpVw4bDfcnjijK1EO7N6QKOzaqZbNsW1zY7fRDWs7qKdY5wXL74
6o+Td9uU7tf7Nb7h/X+MrZ6z8jnvsbpBJGii55rUlhxPT0Ea0wESEUlAlHNytUi4MpyMx3B/nmNy
XoNQAdCl4VKfdlaWeg27qSMY9e7vKJjVW9exrG0oWAYb8hsItZlMJFULFGOaJ484SX+X5Xb2q54J
/HM+UQhHX6ALuwILgh0o8hGInB6I0Xq5ucDdXy16PM+Y0yUNozmQr7PDi8w8FyMNvNMMtTtgTjeD
4XqPG+o48egD05zHPMOnLzeXV8jjKIcfIwyRy/OQc9NXWo5gb9MLtMZlCxgX/UvDPvs40GSNLq6E
CpF8dzqvjq43gLZCvxyMhdE1t9jqxWRQA9ilf2xyxyFOzSlrMfzBXBhtvSG3Pe4ApTF+ppdOmzIC
PzyZ+7GT0sbv4jSS9WSSEG7tY51NpHh2RadDluRKq1I8rePa+jh4PkwHLhErZhUYanTC+51nHgUU
Dv428L6C71EvqbgJx9yxtyaIXzAMa/wZZsE4sOROZRXx/A6u2Z+zBsxu6a5wmwrP66eCmCs4HbK5
jZ99DtMYnIFjBXjxwkYlxoYGLh0LkGOZZvltaTL/IQaIHZTiJ1GCkjRc3iu2lcY9IDBGwW9a++RK
1dAsNhTXlSij0KR8rTcw+Thez6WfFPjzVFyO6DeKmzJh1OMYM4UV7awBwAEhCzq1xBNxwzsb9GPX
Y/VmW2gULjm57g==
`protect end_protected
