��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���8�'+ M�ҙjb3P�Ҍ<���Y�a�~O��!6�:��P�W�����N"\����`��l/:w�V�?�$ΜA����Ad��ٕ�.d΂:ͻ��3A'ݳy����&�������b�}u�}�5�G^>p,�t꺖[�������"�x���k�����eԢ���{�,���|�'�N�UvG����g�F�sJ�k��"���3� K��޸��Y#`��L�p���s��+j�(�uN�0f"�������������V�dV7Q_EC%�c#���($����0�o�k�+�����C|�8M)����K�8%�7�8)}>�A?*�@���>K���︋dx����!��x�|I�ηZx���	B8oV�c9Vs��z��u<g���+��Mn�W*�S��J��f����f��L=Q�� a���6N�ms�춀@	Рչ:>4x����*ҫ��ЎT�dCW�"��(�7��Hl~���u�Z�LOc��n��L<�?�,��ϋ���[)wji�r�UG���L/���j�wKk�3œ�ҌW�I~�h﫾;u�.7�w���j�I�&a�6)ǥᴸ��]K�&�{�@<Ob@WÉ�9�Ϻ�*f��F3�@������ʺ�Qpǟ�3]gR�>���"3W�i�R�"`y�=�������7NeA���L�r�� O��L�[)���]ԋ�7l���]��L�;yH��d�ٞ���A���V��������Y��]v�/iN�I<d�b+��4kk��5�ߑ��=f��9m"dL�r�!��̧�m8��aS0�m�X�(qҀ�������\f�o�{9���s?���gR�vIh�[�������n  p ��2��ޝB$�4: "�h�G-eϷ*�6fc������{MqU����5�r�00\fxnh��b��̳���}i���;ӟ�������I]]6�b�$1��
��!��X��Ϙ��ٟ��x��Z�X��I�p�j��G�V�]wxŝ_:����#ܪ��1yM��2�t���6[�@�`�aQ$���r����!^��G�C]�z�@�����U�0�`�
ǰ���&������>�٤���]�&4&}uu˔�e����~���������81�&>���k
����zJ��>`�n� }T�gm(n<��Їr~��&�ρ�`�𺆙�����2���F�ԃ� ':B��W����ONz7��yK]����c�U�JR�CB���+k"cJ�:���X"�.%g n-F}��A!��Z�WK�#v��#[�Y���G�P}�/�"�r KA5ςcw��Z�#TY$���,�_9x�!r��΍��hј�K�*��zC��ۼ����)q�5�*ףG6�kc�q�#��z��(IC��v���+9
�6~v��
J5@4��*�t%��x4��Z�K��f�:(�
c����a��-���1�_bZsx?Q]Hg�~k-gMC��,|�ʹ|]��ٸ����%r�Hu>��;[�%����H�Hy�"h5+�5��r�_f��W�M��Z2c����,	2IO�Re�'.��VS���u�����\h0s��s�]	���ҺV~� Q��y�:���powTZ�)hfS<B��k��������[`����¼&�%�Jڤn���ؼ��84�&���I�.E�b��Wn�8J7���fd?���5��~��)�j���у":��&~�*��CO�7�u�G�m�1I�~�)k#9ecu*�&�3�'���z�\�CYJ��A�6Z3��m�.���'sy�t�Ž�xCX-��j7����l��E������gH`X�P^K����dt$��3����b �)P*{���Xa��@gv������S�X�#�Ĉ�#�?��:e3�%�?9�]����7lKs�U=D�y��H]p��K����=J��~��Y����8b����UHL��R�7�R��hy�S���i���Ø��3����<1���{z׉V��Υ� G@��L� �g�fB/~H�[��a)�+M���$��T�[Q.W��ǔa:%t�}��kέBU�B�yǼw����	v�xU�cՔ��X����!J�l�������~U�h/��`�}-(R� �E��~q�F<���0��?(��Iϗc(�����<�=��ߌ��,)�E,�YC�8S��>�*�Ԋ������H�>��ۋP��8�${:��7Y�Q�6�����mΛ=�C�p��eo(LxR"z+�u�8�����GɝO�	�Y�?��AMJ�[�8���C�}ɵ�\�'��񰚯��)�"� 7+���2np�̟�1�ARj���<jK��zU���6��g�ƨ�b5!/��.�M��<&C�g�R��u9'w����[B�;'��b��2T�GWh�΁xV|��M�Q�A݉�纡14c��'���B�j|#��#�(4+ ��w�r�hD��c���y�t�a�����o���P��)q���Q�'�[5Ɍ顚FF��?m�~K�.T�3�D/���wQ������g��6	*Mqi00G�D��oLm��Y����s9�a�&�%�-䥞CrJY����V^B6��n��c�ͫ.�0����$3O�'�9ZV�h�K�$�T#�iXXސ��j��B�>�	ə;��>s�I��$�3�������U����!ĄsǢ� NYTn��Q���R�/�u����3BqZv�C]���1���TL�Hά�r1���@���c���9?xQ`���2�[\�{DDZ��F6�X� ���]��~Y�U'*���(J�o#�.$�z3ŭ��f�ݡ�;׬�B:!U��>�N�$�D�Q~�))kկ[PZ��%�\�8^r�'G��*
�����;(�v�|�^m���k���v�Ft���4�:�m�w\�,�i��'c=3a��$�R���,�D��m�$#Y���.'"��[]h~�wT���nA���'@����娣?�^��GƸ'kÈ1FvA#Tgd9f� ��V�x6�������L�ۇCOx3$O���?����op�������"���'�2F�)55���4'�P�e��TT*v�W��:6$EMi�A)I��s���x߫�҃Pʚ�w��L��t��Z���/�s�QYQHG��4f�<���x���Z�o�[��.�`4\�m����y���Qͽ������x���+�+�Y=�	ҭ~x���'F�#{p���1x�>�!A*��H2j�� HԛܓDf��%���v���U꽵�ON���(!���M8Hg�.:�[c"�N�S�@����M��q֎��[��V���e��_6Q@	]D�eyӕ6�JA�2�7�hd5������t8o*!���&�0�XIH�7�%oj{�D�d,����>�H�s���A~��T��6y��G�"&]�� �u��m� juj��D)TK	���,<�� �@����,M��*�ϐ.0�%#&���o;3�:��q`��,����<� �[骖X�p��7�g�kU�R�׼S��;C�������u�ؑW�X�2v8�����݉
��8�sṠ��Q��������Fl�����GP )]cV��B����sk �KU�(�$$�u0���R�����vm�����n(���^z�C��L@V��о_�4�P����V'^k�|ib���ɣ����T8���%����R�%�TΪ����4�C�r�6𗈏���z��^�c���~����X]�,ob��-���du�R��\_�J�6�:d)�Jv	E#���O�*=�2���ǵs�2av�2� ��C�DN�ҝЩU��Ø"�k�d�la����(��	x���&Ø(dq���7�̢�wO P%�\�Ծ�)�":E� Xrhk]�f����Ǻ���[�xQh��ݖtP�7PK�.�i�V�M��I�R/�'�[�%����T��$�<<0á�=�p�'��) ��G���t;JI�p @`��d���|���C��.�$'�*#�G��[�yD���_��w0���b�^qz���̽c�Y��N��Wq�#l�!1_�<�O�w��{lK0�Gvax<8%.3�[?qZ
��*�1r�0��K���(��N�6��!�����1�ҝ���.�l����a�����7������;1����2��c�]�aI���W[Y��J=VU�Q��@��?�g��P�Z���	�v�VU�|R^�l������BNg"m�:X�HP(����
#Ϳ!��(���Oϵˊ����V�T � �l"������uWz4L��5��$��0�h� ;f�?rA�ن��Yh�,���5f��}���1|�C���l~�~�,�L��G,W԰u����>���{�#M����?0�%�$D7�NG�:�ઓ�Up���V�%Nq��F.
�u�(��M���fb���E��)	�����p�[�k�S]t:%r��2M�j���/4�����b��,������C�%�A��Y���`&8Cn�#�F3�C�x�")=�$��~B2VC��(�h8�8�v�t%|-�o�bL��׃�JDU�0�S*P����+��qh��ړ�"��Z�}{� _�
_6Z��k�P��X@X
���`P���E���+�o�3m/�N�P�j�W!�R�@�`n7��)8�;-�v��ig�9x����Ց��r�6; U{T���F-m5�(,����t������H�(�f(IH������9�}_�YN2zt����6k�.�m>���CYfl0&�#5?�E�UmC�x�V('�{�V�e��[5��_��T�U�u�yC�L�{p��8��*�u��N58|�	)�9�C!i�@��b��7�����o2�H�RL��$m�N��3����4�݆	e.�-b7>�3���d)f�|S���Y	���Q=�Q7}� A�(��a#tM�5!��У���Xk�H7*w�w,џ�b}�Nt)�x�?Q�! �Tq��>%�����3�� %��MR��ō�e�MvƢ�嵐�Smٸ��2=E�d��f�Q��9��B�ORQ������9)�Y�u��ѷ�V)�/zpcyn}�B��Za&"�$*%��f�7p�����{���N��Y� d�-��j����ƒ|�MF�\�t��=�_�Q�����PYf�u���*G��)�f�J�l	��֍���zXR��F��4p����6a�+G.)2�}j�ʧ���V
n� �\W�5@�8k��mV���Q�}�l�[r}�O��'�\R��/D5"�{���Ν��),�V���Q��!�����C]=¡�8D&�Ā�r�}}!ۿP�_��(��:9�t2.��?������=�>�a��w��2��������䥑�ݱ;E���OgA���ݖvc��e�O?�5���,�
tTɸ���.���_��P�z�����X���d��W����������]�*���~�sZ�r3�hc��a��8��36+�qj}k/-͒^�r��P��lˆ��\V�F;!���;�����~%�y)K3�I����`��KA
:�����WH+Kֲ���ּh ���D�=�SD�R�X�g��5b��(�߽�SK�;IcִI���$)@6��)]'|W���L�fȧ��f8�t�y�o����Vz��څb���b�r9�0~���߃�ģ6މ=�}w���%�w�M����pQ�����L�q+��G�} s����x�l��� \W��U
yW鹺�A�B@7; ��!�g�X���m�L��&��*�Xt��X�FQjt]U�K
���9�@m{�ւ��E��<��v����Q�Gq�'5$U� �3�x ־�8�82 ����7��S2��E�3Y%|�5l���V�����<��u: :;��<=�����QG���t�
�����b�A$�0���&�������=}i-�ց���ݧ_��?����EK�(`=�CR�G~ƹ6HI��:�o`4�f.Ji��(�0�qvh�']Щ#�+�ƭ�	Z���:̄���J&PYp�IZ�)"{u2P�$�;#�����?�U�3&��э�\c�`�Y�G7q��<h��8朜e"z9/���a���õL�o����2!�m ���⹂�qZqv;���A�tiCW��~{E_/|w{���X#�'>���U*�"�ނ�YJ0[g&���+��>ĻK��+�yG�{�x���Pf���h�S���|�kcy}� @�ɭ������frݝ�qoA[g���	Y�W}=&�)͞��XK�2���W�bX�x�Z|�N[��*�G�>���k�E���vIkq�_Z��,7�0n�h�WU��,Cu�����Wƺm��fZL]%�eW��t� |���^rL�ݦ��ڳ���\���/�h�}�(b�������[���s�(ތ�.��C;)�J�<j�X�����/�ȴY�XI�Wf 7���X��s�[�t&X5&q�.E��"ot��~��+I�B9�fbR�I&yK�փ�����(���W��\e��2�����=6+g��� �_������^�$c�LG����k8&ͨ"���Z[�Ļ:Ԣ�Z�N�=��L�Oڅ"XU�����IB0��S6CX;��~�	��	����jnkN\�G8)&�A;l�}/Ph��ߧE��긨���������^����C���ڕ��tc-Nњ�. ��wdZ�9����k?<YJ�I�C�5ݓ�^�=���ʞ���+�\1�q\Gs8�*�_�%dO�D��>-��S`z�i1�©�3��`��ݤ�$�H=k�'J�ɋi���P�J�x��6�En/�p˩7� �6M���F��a�Qs>��t�--��$jɿT"�1�l�[͸�:J+)V���������(=�{!H��O���h��OQ���l�7�2��w��I��8R��=�<�[����c�޽�����K��2K�rbv0CX~&�����E�=DT�/Z��1�n���8Sx>�a�>�.���G���1>�tM'HJ��:�E���6���V���4��q���C��D_�^�9�x/mF�U�x+6M�Z;^��.��0�	������Zn.0�+��Q��{c���KγR-�a�X���>��E!a�[��$l3S�k����F>��R����-9*�܄�s��������T���f�"�8?�S2���'��F�-}4��9B/����נl�B��b�|`8�f�Ǒ&�.�>�B�K�_�m5Q��T�:D6��=qS\�o�Mر.ø��R#�ڧ�{ʬۗ�"�i�3�V91���r��9�H��e��a�����T/q��>_D��=��C,F��K�Lkپ���:�������,G	�L���h݃��wVL��C�QZȏ>��{��˸�R	s�:܌6�++��EJ���b:�FNU3�����V:�Kj�zc W��!,c
@v��q��.4ˡ�e���t��vq9]zH�Ir7U>cԱb%1����$ ����U]�����y�,��J�*��QF4�h�y�/&����Ȥ���u��~��a�C�}�=��}��{l��E�G�'X[M�q^*/�z>X�(�8�ShBGES	α���o�Y�*n������y����vڥ� <�n +�h~�e��6��%R_k �G��|n?Z�#L�5�V~�G�Y]G���S���J��jF��f�:�ŭ���}q��`��_��<i��%]qs/2�jx�i����<U���B�t�E²іTخ��GI� yJ�J��1Ĝ�"Z��������U�Cʘ�ڠ����Q9�DoU���{O��F�J͹�����@�o��v횞����qc�N����އ�%fk�'�^�*h�S,�ד�;&���綬h�)2�9�QO��B�7�'ƞr���	)��7H)����%�P�:'0M�����b'�!f�zh��[�Z/�ז</���rE�>C�U� ��Q.��+����!,3�Rƒ�f�C^e���;[	鎡�iIH�g���ޫ��`�~Cc��:�����C�am���+:��o�Y5����f�?���
���	��!-��BS�l��C���T����WOH�7��]9E�,�o=A?}i�g�[���h86�5N|��Gқ���~��]߿�B��nN�.��nL`2=`�zv�m� ��(���yl���}�����O�U#��Aƺ�����7���N��a�����v�����
��ɞlk�g�y����;����"��cb3�
V���IÍ�z�7`���7e���1=YT
3�p���q���Ƹ|��sq�SJ��+:��u�!W������	6q
0��
,X	bt_Fμ��wκ��(�hs�f�g>�ҳGg�	�O�o�Y[�B�,�Dr�;��b�}Wΰ�J-��`B<�_���gȭrA7�u����r�H{E"�5���:��*�$�|b��B��f%�Ե�0���Cx��v@��gC��hX(�*�Z% ����B��p��`[Z�b��W�Z���2�DTEGw��G��yM���X�� �R���KJ����ּ6���'�78���̳0��
i�df(�4�������%��x��g�dM�b���3$�n�K�y:��'~b�~P�	 �s
�`�i�0$@�n&�����R��t�ږW���p76��66������Z�k�9^�$we�ҧy6M��ܼ�B�Ȏzq�갢�7���+d��Z�"A������w�9��td`H��-�Ni�����,�i�MeC�{$iO$��\
��/����}��]���L��
C\L��I��i�n&�k��u+� Kg��Q��(@����xt�(Bg��i�9ym~ɮ��*�[:��t�3g�ZGK H�,ޣ0����j�����#����)��1㟴���z�N��{I��ȉ���Ć,�y͆�����`�i�˾Ɩ��i~�T=�}�x�q'w=%m����Q���A���4�����������N8
���>��CF���b�|�Q`_�C�^CLZ`N%@YO�0z6��\�8ǐ/;6�1:�'��{�N��g

�M��7P�d�������vFK�s����}C������+��}�q�SO�O��'\A�c�+���b>V���͠uq�i�&���s�k�����ާ��Xf��3����C[C\���x��֞��p=�	u�8�xV�-��A6f�y��C�Xw��ͭ¯����O2mI&0k灊ћ�Kw�R?/vK=�\V�aZ�>AX��]j�$A"���{_y�Ѳ���I�s��=�p�j6b�o�����ݴ��f��.�ߩ���$�vz �Uټ
�p$�(�~'/r��T�J��Ň�zeҫ�,�������m�C��+Y�ֈ+�S��n$Wɔ�On6=]F���kj�-wS�������|.,���5��j�
��c�4,囖Γ���c?��}<!���$�8��5�ttf��_�R*���/JVݓ �j���O/Tp�YQ�D�����M����v�
��'���Vd�1���:��GSA^EK���}�楔�Y�;��[��qbt���fT�i�����j����%=ڛ����#�X�3'6��:	��Dh��"O�S>bSh���1m�%x�V��@��E�q��'%��y�A��	���ˬ�M��g�o�y���~��ۅ� 4�����V`xD2bP�|Q?D�1�u�o���m!�����ʐ��*�T8n�-Ǆ!q����n�2��Dk��ހ76w����?�`b�J�s�W��@�<Ӫ�h���.�(n���V��k��.vJwl����q�r���3���)�$�J��:�=34X��C�q.E+�h���3z?.{�s�E�H�&��n퓗���d� �8M{���1������ض�^1$�/�d�ʡ��� 
E�e�~����t��%��>n[���7�<��8��'��e+k������O𘣎�uIp�[?"t� �Y_�_�����EW�ɳ��Ǟ��4H���i�B��Y��Q�j''�.i��q�� ���� �>,�"�Kfy��� ������Aߌ�jT-�S���!����$���
8T�!�jѢ�Io��S�A��_n��l�z���Ҋ�F�F.�n���0߸{�q�ʙ=5����D+
������&��TgX�����_p��"N�x��G���%Lbq��%��H)����;���n���v[5GOp]"l�W܅�yDJU�:K&�\"uclg��"�cXk�J��0 z�uJq%m���>���+JU���B2��!�s�^��US��-��h�,H*Y[H��զ��
�q���<Gd'y�G9�u��]ހ�Z��$��
�%7�1޸���A�G��l����[
^�����ܶN[֪��Tp�$��N[��O�s�a+v"��8����4�D����&ҡ�C~6r<)�f}�[߀Æ@���G鈱&�`��91�*W����w�Cy� ���h�p� ����4,zO{)�Ǉ�Ӂ~.�[([� ��(���4ajsC\R���BP*�hVE�n��;Ow����K��+w��v��.���N��hN� !7���������oe �v����!tA�SźdNu�Ͽ��|Zw̾���l~O��Rl�-.�P�)���
��@	�}��G�]��o��8�6��t���AM�y��fC�%��2LN��1\A���]>v2��o��3wɞ����9,�V�"���p�%��)𺙩�c�����J�d�%���W�/+Gy�>jAFo�Û)������Vq�*5����gX�E�0ԯ��$��g�vm�[����J,�V�s�������kW?��Q�ʕ(P(�=�6�^.�+�����"y��~��CԔ�푺���#���IQN�׆��Nnx��+iɹ����*d;�����6rC��NO��BN�����?��Ly<��ܘ��L�c�	���s���3/��e��m6� vi�����aA\���ti�)ĸT��7���{�P����@g��}�ٜ!�w]����Vl�F�]�};�d��Y��z$Q��/^�W J& �q�s�	��f8B#/R�t�5�F3R�b�AHpJ��P@�G3n>��l���rL"��vMR,��`j'�]{:��up�/��S�\Kϣa�U'Sm����N�Uɛ8,:��lR+��S�T��X
�q����3�>L7igp+�6�q����z�P���`��G��Ӂ=�8�MQz��,�`�u��Y����]:_Z�}�bΐ�m�<�i=�|�=���/������ ��Da���:梸
�CiX��e��r"d3kD����x�ߖ�������^5XĶu0 \��{9&�;2.S����.�&!|��j��P���8	A
�q� ����M��V��8a��nz�
��»%qWc�Tש��]o�u�%/�F�η�d����6��+��eΠ�+���L��z�}"�ީ�{܀͜��Aɕ���K���O��1]��O.󚑭ZB����V�<���6��'�X��::���b&>��B'�(ުw�_�⽀3���Rn�Qr�u����{Pc�]��0e����/�F��Y���X��4�Vf�~��j���Ή� ��%�Ar�}��Y.�����+�#�C�c�L�����m���W�Q0�î�яv��V������9�ma�A�HDuu�����=��$���o����e�x�m���w/��D�9d�H�[j!�����l�,|aAc_�OQ��H�e��å��qDG�i �nV�D��ؠ��&h�#�qӮ�!���J�'H
P���<����Lo��:�-k���xT)i˜�q����V��T�vR�V��ˇ,oIY5�I^g�6�������W9ҍD�Iي�:�M9�<��őG��X9f,.�J���t�1-7�����q����JB�3̶I^:���ä�K�:�L��9�����S���`�`�a&�8�����'��t�`���I|(�;㿆!Wia$#�hw@�m3u��js�����%���ysc�y��B�j�8ݙ{�'������X�I0qXE�zV��ߑ9��_����͛_��"��$���Y`×��4��r�����x�sK�^��)��~P��A<��9�^�]F�Ǧ��> �����/6]�B��+��E�m��dG��Z�R��6����}ӽl�Vֱ\&����j���-�H����}"�ӄ����AĠ7z�P|��{��ݐP���P�M\��㊨��_d� )_��ɢ̍ip˕�+�̞��;ɕ`A���?�F-*�?z����O@2�5�Q�~�&h��.y��G��倦'�v+��E=YB�+;ѷ�/�΂)�B禶��؁`�7�����Q6'�ܺ�3Vi����`p����N�^rL�l�f;��+Vؾ?��f��ˑ׽���LU��2�%���5�P�yh��'�J�����|{���aB{J�������0\�Uc���&3ZI"����b6ʄ\�.�^L!Y@����J��L�)G��'y�oT��*ˌ�,�HW�������"�� >�q_1�=�lU���	Ӕ�f�B���d�j��l�H�a��
w��GDW���ZT�����T)��#p�)�|p�O޴���k�A$����ss=�W)?��L����֮�}Q%�u	t��W�Z���[��ͱ�ɞ'8ϼ p������؅a�%���W�=H�o�׼�p��i�W�p ���6)�G#�,���[���<�����YhBh�G�:���v�h������y߶&�	���a�\�"���fC�}h�UR�(;w�R[�ɠ���>��vd,0.1ܭ?W�i�����	�?�G�'���ZE�m���������˔G�0���Dߤ��P��
�,�~~5㇁�5����ꥻkxW�F���I�'5��R�CNa��c�$^��9�/��3ICqc)X�+�k�%kcZrL<uǅ2R�h��{���f�v~�(u6I ��(�w�T�Δ��R�O��qyO�?\m'��/��H$�ֈ��KV"(�AE]~�[_l)����彨H�GjҊ���JJ�>�آv����;\?w%��n�y��<�7�;	 I���l"J�*�KŠD���Dh}��}R��)ӵ{h/i}�F��z�����TcN�D5.�+^S��VI�뙐~���[��Z'9�W/(�$�l�':���E�)��(FN������s���u� �n!,�txN_
�nY
g����{���$>/����l�zP	R��Е`��Ѐ��'#�}6�I�Of��@ah%�~;���$m�c��&l�^ilb���ù&ܨ��ֺ�+e�(ծi�P}�YwB���q��4 ��^�=c|�O�bj@V��������C�ް��r��a K��>A��ɳQ�y��	w'�v<��t�v#���Y���.ͦ	*-3��
��2�?)V&��!���37�֌�4���]`,Fr�*At,����J
�����-֔w��8�_䛘�Q��Z}�) ���:�&�U��{�Z��u^���8�6B���V�Z��I�!=�9�<9��"۲mb1�$�Ӆ���q/ײ�i��д��4{�qٯ�qT��E~���i��>w�m���mgcs
��V[8�>}c<^4�v�bo���v��m(��a�ܽ]�t�xvq�������G2tU��j���̊������|���4f���p�m���~ė]�I+��߯l��,֚ŦS
��kLI�]Y�sLKf�Ƙ%�y�Q̅j��BI�� �F6�}l(Q�FD��u_�c|��o����k<��#�EsѾ��Xl�+�j����ɼ���mdopfw5��F��<*~�^$�a���0@?ᓁ���ut��$q��]� $�m*�9D���R�܊�om�R�� ��&�����e��o�
N��7�Ni�z�@��sjiN�Ol��E,Ёh��a�Ә��W�z���PɌ�E�wQ�7'{B6�2b��m~�#e�;��9�`��%��v�YGW+�+E<��V�?9��
�N�G��@*S���T��3'(
]�]����#��������na2E��)������$WR9\M$聼z9���RɃH�x���.�䇲(�V�]��+t���<7����/HZ�i�a�qz�Zui���ai�a�Hס���}�P&�5gѝ�fyܒ7ڢT,3�v��P,7���2��mc�l�)Z�{�o#KlŜ�5.kts#GGɻO{�!
~���3j��(|X4�x��2,驂r��C�5�ȊjUj����1�3�f/4�Κ�c�p�!��m�����,&{�?�˟.�%�5�ke�5��_H�S���u��`M@8�ֲ�\>룜�O�^w�T�%l�ʺ&�9,�$�S�T; �2?䋻����7���rS��j�kN?�h�
��L�C2u���hJC��S��_�%�m���*�h,�s��%��b�{PH�Y	1\��J��D�t�#
�Bs�/��D̢6L��ҸA��W�j��ӿ4����r�Z�r�X8ko�x��,װ��3��-�̭����p��֯{$>�p�6�[71��Nߨ�2v��7~0�ѱ��4 ��?��@]f@�Mgw<�Px�R�>RQ�B���4;�!�O�*�-b�M���ʇ��8�6�$�8����0����߄��|�l��Іz����LW=o*gy<2�W��^U��n�!�T�w� B�能���qGn�\<�J��h]���Q"��)��� 3b���Mq�Ek�y�Թ1!�i�2f���j��w�e���j<c����7�/h�d.��A=�l��H������f�����`� �i���y��r���P�@�O'
9������D�3P�z];�l#? ��G,EUG_n��C���nh#_x?d-�A>��ԅ��^��
�h�	 W�z�N�����]�-�YD��I�Eb�`�N�ؙ繷kA�3��~ju}|B�×H>�����W�p7��J�Uk�{I"��?�{�f��n@F�/d:(�/s�N��(	!�m��aQ;��~4�����������Q��sQ�l�;@�U�MxL[��8p�ȪК�$Nr�
c������7���h(���V�r������4}Y�Wr���r�>��Mut��I�G��&A��	$�R�	���1��$����.��B���I�����Ҋ�HS��.����a�Y�v�ʈ��(���x��������>�&e�6nJ�t�����b��D q��,fܝ��
�#Ls��)���6�v�h�`�<��ػ��ptǺkJ?���<W�w!�:�4$��F�a�#�,�y(f�O|0t`��MsL�=�[kŮ�bc��%t��r���D��?�@�����B� �@��l݉~�Q.�|0V;��;LLa�.�&i���\]��B|MK2�4�D�Tl�52N���`����w���̱V�$��}��T���S+D-�6S��$ǿ����J��U��f����d���u+�d~��A͐����$�֜2�{���:�T~�NMW�>��قE{�̗�p��#��?���7�O��F�:�.F�A�R..��T�$$��m�l"��m�O9G4>ܣ�/o;��T�s��B+���'A���؄�<&>�tg7k%!0���O�9_��i!y���'l�F����'��7l��� N�^T|�X�@">"�����d�Ʌ˯4E"����)򝁼�-d�g$��iN�����
Jg`��,��yF��Pe��'p�P��Y�hA^]5Ďe�d��[�k���ɍ6��v,pl�&��֡p��vY��9�A��ý��ĥ�X�'�㯁uE���5^�USP\al�&ɟ,e��أ�I�,��a8)/{
L�G�/�\��֭���cP�
�rrj�(;}��.���rz��d�G�~���D�.)�x11�6Sj�]�����I��8��Xu�l�y�R[k�ѷ���6:{8pT��	�/�(��ٝ���&�5Y�G�Q�3��yX,���k�=����9}!�/� �F� U�ޗ�M�i_hȊ=U�ֻ%τQ���^�����N'�Ǿ�Q���*��e��ؒ|���d��t	^Z��8ae��U���D܋�_����Ѵ�'��l7��ފ�S��x3?��'�}�V�,lIo��If~hY��U�8���
ò��>��2ޗ. ��g�|�`v�a1Ҹ�9�_�h���#��2�l�
��G;�:�`c!p��ж���%�e ]�!�6L�3���B1G��VnJu[@ �
�����[ĸ���Q��-s[�~�t�Qe򎈒z'*�� .AO�,R?A���u� �1c��N��tWcF�"\�J�i>`G�f�p!�lxC���b��4���k
H��P�j��i�[�a���\u���D��L��l��S���4�D/֠仠 f0d=Ś�t�w���WΧ$j�����\�j ������g1��� ����]�<Q�tP�(�-��a�v;� ��U�ǻ$�W�FEd�
ad�$���_zL��$F%��;�Q�+K5��4;g܃bJ��L�3����dY������us�tT��)�C�\�1¯�%�݂v��g��3��>���\#�n�6�a'�W�e�7��K�ڈ%��:�|_G��b�Gf��:�\��X�i��aɱ;7�fy2G�� ^9�Kj:B�)%G�&k�N�zc��R�Ab��h
�:;hM����4��8�?v�xC�ԽD���\&1���/Q���>E��vWRKtɋ���q�KqY�� �T10kd�˵c��'\j�;[�1)��"W(�|�j���0zHMTu-�!��b��w ��ll��E���p��x��Loz׌s�����vƷhT�����?�N�?�!�o�w�,���)3�7�U\��^�dX�Ci	橈�l���
8�$cN��`>V� �i9� �
����c&��?e�T��O�L�]�����s��,ik6K~i�>�J�H.4�Ǘ�Hϣ4��?��PVR�A@�f���:Hn*-��	[/�Om�����')2�4ch�?��AmkpNښ�bo���|��B80Q�3�i�˔��V�4'��s�3�����S3��S����/�����s��2���o���N�
��Jm~Z�]m�	�9�x7̏K�*���P�J��XTMt�r�g��~��k�����u��L�6����-K�H�M�r
���) [�.J��//L鳗��ŨtY�ө\�<�dr���Zv���9[�`Q��4Q��Cmo���l�f�.>K����w�N�к(�R�R��6�KH������tN����dY�+�#�G<�g^�;�,Qs��y��<�N�C"��`��f���R�ʽ(5��dgB�O�8E�uArZ_`�F4%ne�sp���_L����L��'K�u�������xU�A~"���E6�Da��]D(bˢ8X��N��b��e`�c��2Z����Ԥ!�#�=(t�?L0�ǞZ�I�.f��p�թ�ܻ�w�`������_̷�$s�ڵ:O
�ki��	(�kM�Y�m5-e�����jž�����sn�+��Jϛ_��u�p�W����ץ���㺸�ǒT_��P��8-�_�ʔd���ξ���n�o6�Eo�]@؋��;Yx������Әf_s��Nvi�x�{2���\Dn�P��*������H��)��0�������G�YT�!�h.�/���<J�K��
�j�A�w�A�PU6#y;d0�r�Mn�u� i.���+�Ϝ�%���?ED*v|�S2���\ۣ��c��h{)�=�C�<_�M��0��GJW�s.�4VB�88����ퟋ5��틨]��{?�f����iK�S�N�9N|��	^\UߙF[W�B+�bLU�W���Or��h��į~M�W"����+��Ӝڡ�qFIe�^�G�l���q���']��D����k�ϗ(�w'02�\?a�̹O�a�xEؓ���A�ޱ�f�l��&�48�8`,R�Gq�껮2zn�y�ޒKU-<]9��dV巎	>��*g\�����h�;����]A�I8&~�H�ڪ�ֿz�?�X�#�b�E��F7O�r�@��se�Vdq�Z����n�{;KF��N3y	N��������ۗ]E.6��i���d��0��8m�і�@m�Fxxf�@
j�L��tk���<P+6�-��}������'pR�5���8���	<L��O7'	is�qS����?f~˯�I�ltp'�.��N3��aD��+�9�E�A�BB	�x�����V��F���f�,�-댲ކseBߡ���ݑ��c��p��=Q�6��x�6#lg	��zԻ�gθ��_���!ŪLڤ�1l����gZ��*��,(ļ�$_��[�Ɵ�~�c���9�tb��*�_�ͫ��H&)�0�DC������4==`��"�.6�|���q��2�a(�3}�۝R��M'*���������U�rA���SK�5�>�\�m,g�d���s�Q�0@��ɍt���{�S��B��G*6ص�9�9��S[�Əgt�RGB.\�ߴ�/ҙO��߃�M���	i\��g���9�s�t�p���L�5�����8H�gH!�!�r��t��ٲ� wSz�P����4��b~0�m��8�:�S*���š�<�!��YPl#���I�lq�h��̼�:k���xjf�����V�� �э��F�
�pc`�ߚ�HM3jF{��ե�+�._����e2���4�'q�,t����s���MNF�[ƻ�B��q�(�1���>�P+��k�&�-�����)7d��̩��Ӈ&�\�-��<���B�)/���zm����c2nA�,%�����T�=(zFT�P-Ks��Õ7"X�	@���9CvJ��
�M�,{�l*	�k��K�,���I mMP���}W�f�!�J�lW����V`z������h"n�O�	A���^��#�;&-=]��S>����z��J�oo��ư�l{Pvv�����)�xBVw2���`�̔9�Mk:�?|��l/��W���$a��$\&�j���i�ǒ���N=��&�q/V�5�VXEW��Ԯ��`�l��D�����/!h��{�"�U̦���a=�J�J-�����ޫ4�{�r���l�Vx�{*�����Wa�0��V�����;������v,�k�ٝlm+���\mf�������e��"V�ҡd�6��A6�*�'�\�B5��)ӧx����J6FR���8L8%j�[F&3��2#k�S0bS��Vp(	��S#=�)$�e~Q�G$���Q^f��c���'��{	R�����ϥ��h��i\���T^��p)x#�Fc߄ �r���^`��l4��1���2$A�ڽZ7�8b^e;���R7eT�Sh��Ab���))��?$����:�G������<��l�R~�J�G�&�VatE��R~��U�BYΠr�6�	�do�F���j�ϔ�FdT�5;@7��![0i���g���>eP�pTd�5x1�&���$*�u���x���	��\�@���|X_[�f�������q����&����j�E�21f�	V�[$�ߟ�;����m�*�bǜ����}p���'�5�Xu?X;'�ozo���@Z�4(�\�{�n�nAנZϔhz�܋a5!�U
ҥ2��Cb(?w��g3��e=�]0�][�Q1 �����m�?U���˳ަZ��yJO����`2�M����)��X�� ^���8 ��Bh�2�ʿ���2l�3Q��ٛ��u�������8Ƅ� ��e"���h�c�XK��ɭ���(80b�����N�\n�Nϝ_�w�}��3��4�_$�.�L�!�"�M���D�����{q,fj��WK<T���hX����"`^	2�����*N�Q!� 3+��l��]�"�|�E����落�e�G�m�5q��U��%�c�-A�>Ǽ�� �x���8�&�|�,�
U/�k�|����)%/d���J�ZojM�ߨ6�*,zsYH��Y¨�h&�A9��?S�U�32ڧ�)����8)H�����r��S�t���d0>�@���,�,1峦��(6�|�W�tM���᭮lq��k���c��|�����a���aʽ�k)P�J�G��~x���5�����G�#7����' 	�� "}�KZi��_�rLl9$����_�9`ܫ<�@�\]l��B�|~!�0禇��"��o���@��|�Nop�#�{���1��%��E-���(��2��c�Iԁ�$~��f���HO]���N�� ӗ��7�2���٠�ɀh�;��O��1S���~z�΅ě��|d���t�`L�� ��:��VBXwJUi�)�~Z�!>�����a����i�G?����	ի<�'�,�rh6i�,"�`�tO>�KRg�y�K7��,J�^��p KP�v�ȼ�B�/��^�!��p>��Ї��G��SmH3�(?�[R�!��f&�2k��J*D�;��Cu3����)əʺ�N�y�q�}�8��(�RӒ�AǊ�ô6�I��������2ô�Z]��|V�4۹�W9�t�D�k�Ʀ�E����\U.�a	r�5r}8�yo&\Y;�y��/�J��ë�?���(�![��*�n��2���V8D�8q�"��DT�ܖ-$���𖖧e�ؓ��1���=���_�G�dĥ�R��H;Dl���j(
ɏZ@��8��͑�!�f��4�-�t4�w$^�C�~��PiQAhE~�f� ���HL��L{V�;68�&���C����G]���u���:�ee�U�pG�jK��^�S7N	�>����ƌ��9&���6}��ǡ^���r��V�=��&��	�42	��"W���b���&c�*��$h^ J����V�6�omޘ�Eˍ���j�1b��M��hb�p�f����������;���R�y\�> ڪm�Tcm�o�I�9	����x��u�d��&�6ʧ�&%�hIlx;�V�CP�_��h�N��4�	���/��׎��Q��&���8�P��1+n.0%!���R$���u�5��㝁�"�'p���j�p��q�|.C`$�� ����6B���%R`3
�A��'|˗6���A�����Wv*���oB:�����k�]&���B�*��|��N���	r\Hy~lM6	�΃\�b�3G�+��4_~��F�З�%��|-��b������XE��0�z�V۰#����s%�i�f�P+*s"�T%� ��#fNF.Nu��?�Z"]!5��[{G^�����\��H�˥��=������\CIA�r,Xl�гW'����w�!)Fw�$���	ur`��u��h	��h��R*ٲ��s[���P�E�3�\�|�&���J�yp���]*p'�h p�2�=�-���*Ɣc���3��<4���%{|�N�n��ޖUf͐<�"Bd�z�M$��	�qh�@~��jW ������렡�ʼ��w^�.}���W����ؿ��H��/�R����Pq�:�n�O�������&���+����p�k�Ƽj+����,��h� ���ԙ^�}{= �hV���̞��N{t�N�`r���c9ɪ��'����m�#P����>�zn&� ���^���)� m�x+�vd���)ۻ;�8H�WVZB��ᅾ9fb��%r�Iob��
�����Ţ��t0���MF��o��J?_ݦL9�94�xv��^t �c��w!��2�ʌ����a�8(���a��~$Hb�5�������1�W�Sh"��Bo�~B��Q���� G�dJ2va��+6�\I�#�/<Mg���4�7�����L�Q�J�xL���7��&�lr�Gj;�6-T�}!�/s���!5yp����`wo�_��k�]��B�[x����I���D��y�Am���y� �C�mky��Ѓ�_W{#�g ��-+TS|�:��7�WV-Yo�*��3��W��'� !���C~���P�遪)��	�m�m칉���мC�����J�O�Y�f����H��P.d!f?��%�en1���hI��9��
�K������1��m���(��89���>�N�	�WT�F�_�b�`���N�UdH�4�:���>�Ć[�:���F�5�(��I���Ԥ�J�N��Q{x�l-���K@��� �\��O�3�M�^�шv������xסì� ��@7�q��i���^%Op�+&0Kg���½��x��bڵ��/ۭ9���xK/����V�����R�Z��ӻLΆ���FS�������(�[z�WKV��׽SG=���J�5L�~���Z��,}�2Ҫ귩��El �g�S ��T���"R��d�vʣ0�Y�Ϲ<+�ừt_M���Yo&����8�^�m���LȺ4�J�h2�׫a	�p�ٯ,As�-{|M�\��QRL
)h��K'"�%��s�!�L���f�'p��WÊ��+G>�x��~:�+�w����[���n>��\�2+�����0�o����y_-y����}uVE, S'��`�,����ȣ���:�Pʪ��Doц�X�k�Eh��H0h��>;#f�E[�:�\�S*Cr���\��K�^M�5�����9p���#�V\(����k�]o¾Q�	��I�R��:���!ތ��M�da�8e�:h����rw
�k��xhv�ϓu*0�w&�Ӥp�O,��,>ÿ0B�Y�;��z���^��`X����X[��SK�"�i Ļ�b���H�5E��Ҽ���w�S����]�w/ݜ����j�H	@�	 �C�����Z"[��ؙ�W��$d�$G>�2��J��`)��ǂ5;I�0((>��
:�(�L�k�Zp��:ɔ����GPf��/���79�Ot_|��N���7�i�.���.�?��ާ�i�g[g�ȅc��!H�K�o'�͡lӬ�y���µ�zPN,m��^&��<��2H�j>���N�/!}�P2�y{��rN���M�7Ԝ�n#6�5T�����Í_?C��Ӎrkc�d����S�,kX�oo._��=ވ$m�a⌮mC"sӹ���U�^	Xdt#r=E�q�$t�8���Ԣ��M�2�\�ムE��	f���%���6DV�aSA��h�Ę�o��U/������y-~_�����1��k�2Ш	5��	?y'��u��8�c�
��͵���1lr�"�[��"����=�7dl�|������	�U��'���m"�_�����2E�*&���{�iK�SA���G�(Y�y�s�(ӗ��w�o�D�!<x�ts����}��8���%�JUt#+��U��&��2(�����i����~@�����4��?�A�;
��L�6�ݯ0=c��S@�?�Q��xxNN<,��\5䑔���hz�]'��J;���k!�.��X	��ɣ���9-�1�
�&���1�+�[n�3�ߥ�D�Z��n��_��̆���L>3����KG%�
Ѽ��?��ִ�UI�5!��a�����i�/7�}H���l/J?d�cLJzǬ�_1:��vEeP��M�MY���䋿��UB�`�2�v5X��HQ%O���.f�,SQ�����z�'?��w��
�)p���V�/����Q}I-�5V6=���0�#��!�\y �uoQ.�Q���V^���x��BhY�g�ޮ�]��q�KVd.����ݲd��0�� E	|!�}:�j�k=�\q���L��v*�2��h��8����Ӹ�nfo��W�7Ϟ�p��A#���D� 8���9O������d9ap�5d:�)`Lf��c�G���*S;�		{�?aZ�ᾎ����"P6<?�S�	5)���0>�7��ܚg���VM�tP~����FT_	����eoV]��i���g�G6�`��t���4&�{��o�@Z?]�U��r�l�Sx�4�39�E��ꢑ��K5*����13�m��E��
��y�B@����y�nJ���&\�+1�n��&�>e�%�[�����u�)��T�����4�n��Ԑ^�i�����!
�l�r+�g�|Z
���!�FW��7A�JM\(��א[N�+�~Ȍ����[HCg�؁��U��V{s���Ω�]�k�t�}�c�~+�t�[��'�Iv�Z L_(�I$���:Ő��v>���8�}��_S�Xr�8J��1�KU3J\!�W� /���Ed���܆H;[R�懁���J���'�+[��,˃i�ŐH�͸�G�0-���i�AoR�j��g�5bH!�$�ю����-F,\ҭ(đY1�f�[sQ�VP�RQ��hT!���ѩ���,3<�~St"P��¶hȝ�����n�\����mO,GrS�p9D��7Q��2�ay x��3>ЯB����ꔂ��ֻ�$ċ���y�"��� ��B|�<Mi)ފ�.C�����YN����'\��		H��a������ȱmD��G���1�M��Y�}�)���}U�� G�$p�H:$��%�A딍M���×�(��`J���Ye]M~@��6c�з�X�Q-��Դy�Չ!q䇳��x��7:�y�"+O�d�Z�G�H���;���q�6I���Lm&"�_[�v3�n�~�4���ziW�@�Q�ц4�8�'��N����m^�6D7�G[��v����#�z0BR�>�4����3v
d�5~�Ht�0��Y�SQ�T@����V�H]�7*Q)xA�oP�w��37?��R9��3Z򭙭�E)Y�6�O��G�?�?�Uv�Ѥ9�x��jg4�1#̜��� �S�j���>,��S?'�,Д\����]��<�=ǅ��!B<ѶӺ P���>�ǈS.E�+:�0鍄�.��e��).�a�Gl[���Ϋ *��G�驾������&���٭�u���Aϸׄ;$�Ϛ�"���q/Tf�_�4�(��j��'z����-�U7]v�W�d�����[�G�-��7t}a���o63n�"��j��#������F�ڭ�T�O���Ӗ����L��ȹ��zۈ�s'`=9,(���hv�l�!��sTt����o�R�,��*Cl�����(�cg���&�yT���a�q��e�]�E��3��95��Q��ߕw'�A�#�*�p	}��Jn>�6��l(�b�j��֏��5�4��v���<��XD�>526�>�-�R�$��#°b��Bd����"D$V�|Thn���3M$Ui)b"�b�%���^P��*��~��M����%���(�A�ϟt"=��M��}j�Dڤ<��y
�Kƶ��̊�}���h��S�����A���'�ƃ�H�r��뭣�P#�Ϩ��bN�<��"�ҹ�~����r�d%0w�X���r���}�R�b�F3�+��1\��<����R����O�ϥ���Vԗ"ә	��g��V>:-�'�S�zhy�Z��Vp��76fC���'��2.g�1:�Jw!L(M�?��@�ڃt:҉w���W�	�D�D?L;7C��2�_����s1s��];���Y2�����i;h�9j�A/H�b;[��%jj-L�^$�Gp�i�5Ȼ�x�����b#���;��;����4��@Y�%��0JP���K���[�O���ھH�,��b�?��+�$�R%�=�� �"<�B�iZ����US& ��΢ovJ�h�urKAb��~����e&��0T�Eň������*d�d�Ȅ�*�&�]{��l���7��Ð7�|wm��`�e�7%h��&��l����8>&�XS[�j~�t��_r�0T��[ЫR~�{��*�򓡏`݆xBz������܀�\�"JH�[h�ݱ]�Y�_H��bbVH��!�����S�(ӛ^R<��ˠͰ�n�B�x��i.��@��4��\���]�:�����َ�X�:�}�G�A
3����h����r���=-(F)E�(^$ef��Do��C�/�yo��eְ����-c�H��F���$��J ž\��Ĉʺw(����y���#�G��4X+��Oo*i�!,���1�7��?�\O�����D���h-��hנ�J�x�f)��Hq{o	/�lj�r����Ĭ����Qy�9��3;��D��	������c�)ϱ�ɮ%��Y�>���mùX$$�٢1���@�����p�j���M(16�P�}���� �cxѷln��q�d=jR�/�鈾��I��CĶ�m��S${p�#c�:����;��O���H8�޴��GG���n�(>r���'�(���(����R53F!�S�	j<J	�}�&[5g����Q�V ��y������ _���5W�D���_fD���@�2�"��e���@G������&P�Ú��"��䙵`߂��P�Y�wy$��{�?vJ�\	xk��ŵ�J{f��S��Sk�o/�U��e��.��򔎎m�A��{�,ݳIR4
b�)]�ٳJ�^O�ɮKg�˯��#��縙	�z����X#H����UE�;�0$�"��`eY����E��u�Q:�VZ�8"���c8y�]s�'�;vih!�Q��Nd�%%�E��j-҇�H,n+u���G���u�X�41z�;L_�Х�{��oA���k:�Z#o�k�bV��gV���o��(ȷ���ar:`L�m�qqet�o��or��F�����$��k�JV��&���j�!DC(�Q3�sb������ �?��n�5��=!}�����p�4�ʺRU<�F�}��9����U��w��:	�������S���zŖn�kkC�DT�E
�.u��
b,.Q��@�Y&{�ʹ����ȁ�'��L��"�&o�ދ[%ߣ(2X�"�d6:4,()==������:��������2Z�ɠ�\�v8ܽ�d�썇aO��eX��5��r�2�f�(�H%�~L-<�7]�I�f�����c��F���Om�V�F��&a�JQ����<7�GZ7���U��}��`�Ђ��
t��\���Z��	|~:!��Dx����ڏ�
̼�1�G���v	f	�]șrJ�E-��v2�6��m�I������l��RԼ)?Y��K�h�	���$���G��k�����e�4w��`�bH�QVR+ʆ�s�+��	5���u���?*�i@}��-h���e�w/q�Xf�]݃C���%S���������j ;�ߣߺ��oBz4n��JAmѹ���+D�<��>��->�������B�s	�yg�S�[7w��Nu�R�P>��홖>7"n tǵ�Ǩ��������9X^l��I9k�UQ��;ء-ލ���?�t}���7�Z[�7%�R�x:�T�?���;�F{�,F� ���{[f1K�?�x��J�
�o��e�!N�;�ܤ����j\�݉��K�V׷/���������Tj)��^��`�Є��ٳ�g,|,.1��b�-�[��/������`a��3#��`u�쁂gbF��N��cn��Tf6��E�O.��zm�"���<�@|�`S��\�2�'�t�,��0�c����0ue�͝L.2�ʶ��7c#��p�����]
�N�.�!i�n.eДc��{�a��#-�!�	����T����<�m]_���8�h���J��8�|0�8�t��*4�������zyr�2�юe�|���<uF��<�V枴�Y�DV��R�M�37+>�$F�(N1�Wf=��H7 ���~�&�;�r��"M6��nwa;�0˹�UA��;'�(��U�K�h�!*�\���n%;s�A��:4N#/&�ݵU-������=�Б7A�H_G���/3�Nڎn&Z��~M�.loN"؄4��n��yFT�]`�XwA��%��>�Y� �{E�8�;�G+�u�V��x!+e��#�maե!�b�X�Y�iP�ɱ���O7r���;,� g��g� ��Ta8\X�_mA��[w�����;��.�l���ʺ�#���},���Gg�d�j����ve^��{�N�KI����N�BD7���%W�ΊQ�HO�b:�J3}�qIէ�y��.�T�~��A�v\G$�d�����K59o�	>��������'�@;x�p����<q��
L�b���� T��(�� ВAmcr9���^;�?�H�Fy.��Ҙf�ݳACdva��ar��+�T�i���jJR,�L���7��;�3_q�@ϯz�������s����~@/�k\�ق�_&­��+՞C�J�p�?/�	�NI|�%Xd1�#B�l_��}�l
5�P��.=��4��q�i+�4x(T����9:��]
]����m�X�f�(�Q*��ZhQ���4���3"��պ2�w���L��Dm��?��8
"�c���C�-i��K�'����f{�M�Hf;D�{([lt�߬Ա���s�
�ZY�/]H� ���ߎ�P|���<�2PW�����ˤ�'��	B�|�� �E���~��&�ho�7��o��H���f�+3x�RB��*E/d��["����. �Ri��mv{��1���_j��M3~r9����<X�����w�'������	��͑�:�]�àsҬ�+r	?�9�@�7��(��S�03Y{#���{�pd��/��D>�ŷX�[.���};?!���	�@/.��	˘���v]��|j�tY*�Kw��t�+8L�|��:�F��ݞ�����0��jcV2��Zb��<�����#���W�4�Z�S�mn5���V&��#<Հŗ'Z�����3K�.1J�B��̝��<Q��8���b�!~��g.�Ww,��[HCnpl\.N�]@T�r܉6��ؾy��I3��M$��fש&ȆV�[9t�w�����c�Ro=� �(ɶO.lQ�� �Jy���X�Q�v��H^�|ݯ����rs����^��A���c�2v3�Ĵ�#�k�L����aK�Q���:h��j��d!:0�c��"�k�q���:e߻��N
��J�� ���+W�a�F�����ޏ�;��VAٌFW]�Y$LOY�f��{qy\�kȅS���D�qbXkd�]�f�����^������jm�x�*$��ɋ%�A���S\ǹ5FZ�Cbr*���U�f�v/���$UV�H:#A=����y��}0�R�U��0�����}$�*��8T�  �78�}�m���ޅ�'�3�RdU����=�����k	2h��|�bg�Cq
�f�"k��U���}�9��v��:X[��s����\�N��d�H��od]�˟�yMo���>��d/�%f�������+K�s1���I�YF��@����M�!���XH]���+)������G���Ћf8��fĤ�{�x��Ĭ�����)�?5&�� �z�����w%6�Z����	���2��NP<���a]���X�J���v@��-�9�e��sC
��!�9��y�7�Pz�e)��Π�� w��K����*}\:>z�}qP:����H�@�w(��$�>��VJ��1�
f�MyҘÂ�@�|:IT�kA$���ǚ�po�O�����O�����mx%�B~� D}G(���m4Śv�c�OZ�v�&�2�Y�DOe�Ά�|1��e�|4%(�l'ä�k�
�ʀ�!��?����y�A�|N��|9-=�|`^h��Zi/f#� �
� �a�F�;r%b5`�(����Y�Y����{:�:zgv��E��{�o�4�)��q�>���F���
B�&X@(&�Ģ���I�=�:���\���/���e;5��_&����(�����l���#'�er��IW�j;�!�Խ�w�X�S4yH��|�%�F���΅��9zF��W�N�Ƈ�p&���I,o����y��s3I�Q��R�̘'��z��pY�\'u�0M����<��Kj�枱�kא7g�r�����-��+�Rk�G�/�)��R�5���?I^�Ԃ^�C�{1 K�ݜ�"�#ɨ�3�y�P4�c���T.�xB(��K;�τ7�k�z:�5�n��l,�5�
v�P~�Ӆ�(�,0�����ޟE5� �7�ʪ��RT�-�9t_�/�!��h	 �c���9
��~k붏�D�$�ӵo�p=0�Ք1[TW�An��I2P�d�!ZɈ>�F$���dC_E{��-����'��o��$��}kQsZ��t�y^�,5>?�U#�QJ��eK; D��[�J�����#щ	�&��3���{�ў�LD�m�a��Z����IT��L��ϖ,OZ�|����T�DT��p�L��[mA�5�x'�隆e́�{���g�k�#	�5�%��ğ1��ߓ)^1 �]����4����W�A�������O>����K���m"�pBʬ�>�8�`���@uY��/��E���j(������
q_�E����@�U6���|\�_?wd�����U<O�^�7�8�(��6H��Y�N7'���<�R�gBLUxb�1g4�Ďm��H�H�W+T�"�x���zR����a_z8N�gNʏ�2+�ɛ��+bex����K����ލ�q4l�}ϑ5���>v��p��U��j�#<P��n�f���L��?S���{�f��B1�.t\�q1x4���ٻ���q�E�M��76jf��_::��1�-SI��f~cJx�+�(��.���' ���bl��fkz
�i��5��yM�I}d6y�L����Fħș{�O8��[��߰Pp|y�vu���˭#8,I_�w��P�_�r��Paʳ%��j��@yݹ��2���w�8���Ұm��K�u�])��j��<ƒB�k¤O�õ���(P�+�[f��(3�]v���kF
sW�8#�y4l�{�X(���@4��W���1:�w�A��
<컄��w��D��g�E�	D� ���Yk�(PQ�V��od�?0  =��{X�����ղ��*g��>9�Z��Z��ѻp�-�12�\޴�K�['�@�5�ٽ�+ȵ�Y��T�f<s[U�(�j��Q}>)a�z ��%w�R��a	o����������d�g�l�G��VQȂ�@�=oꋢwVH�O�k���Ӽ�c_�`B�{�r���=�[X�A�8�V�(���)&�_���ّ��CE�<rm��
;d"c��
7l�1����6k��D�q��E�u�� ޽�J����	݅��@iMyv�[g��`4���������.���q-��gI�����`<[ڊ^S	��G���;���{ػU�"&SQ��0������P�g"�Dr�紳��bd&�1�u-dmftz� Py�o'�Zoy)�FZ	|�y�}�~4��R!	`���>���#@�+9Y� ���E�׫�6`F�!�H$�%��Kc�'�j/&�����������:Ge��"���QOJ�v_7�o�I��9�O$f9J5��C�l[-�q%���D +m��.'T��:�셚u�i�n�b2JE���qt�=����2���#I�l뚮�¢qpƙ%��L#��}�
,�C��z�O�/���7��k�%�Q�N�
�F]�{�38�[��c_�ƻ&��$$ K[��z����oH�]��������z�؞h�`�>�w�Y�e<�az�|�j�Ǥ�$E�K����Zo�L	m5M�\�����]�][p�< ��6��v�-��4��%��QLS;�F>ͱy*����Q��A������(p�B=����W��M��o�J�"�_oݶ�(˾�Z�����l�ߠEw^��۾u�%O�=�M_��Vb�$E91���G�/d�^R̶��O�a ��P���=��A)�<��T_��I�ֈ� ˌs�w����cj)�����ă�[����I;���er����q��'F���Mnn��I���*8�T���L��#ޯH�F��D��EC��7�F�@[�ƅ��Y��M'��zO͂�ޔ#I�)߭{��3BB�'�x�u��a 5|��0Aƪ��)�X'�9��S'�Erv;���,4������s��z�n���	#�3a����E�q�۰�4�o�
�׶U�i��T��H?�>t�k�+�(�%�:�$5�y�667��ٽ_(l���z��Bx��h�n9Yj7� ���q��	A|�t��d)J�=�C��t4!'�[������{���������ɖSqb��6-���(���X>��q���.8�	�>��F�r����xq��8�맢ž
�lOo��z�����̛8w(�񈈰p\���>	���֧^sd�����CP1�	?���me;+m����~uOѨD�zt���VX-P��(5��&�{�(��{�%n����z�Ay�&�C$O���]n5�lgt� !�y�c��9����Ġ5 �
�����$�G�a��-�էF?���3Q�i�� %U�������W.�j��#r��)1�\c=6�/uX`0�_�#F)V���t��ƅ)�({��ٴR�f���Xe����er�MΣ���^pquٶ�'o%��c1��ŧ5^��~��o���l����ԚJ��>�����1�5�����}�o���r�7��S?��m�ܧ&��c]0 ��x r"�����
ד� ��A& `m��a,n��Ry�Z83t�:s��F�|�>lt����!_��lȒ< 5�;�tK��@�#��?�R�+}P�X��:�Fyq�/�Q�*��_v08���WUW�\q�{bX��u.]�����M���U����ՙ��ZP��dRB���1" Ζ�Q�?�s	�����f������{��7��/W�H()GH"�:�7�4�9z����_nL�i�cv���q�:�1�"6TS���fAX�zv�BT��o����B�
cr�=���j���Ĵ5	����G���|�!�S":���}�Vr��KԆ5@8����\�����Ɇ��p'Y�Cݨ����X���>�MP�=�F�����]s��F>;�zAh*��L�z�H���I`�Ǖ����t+AB�7	���� ���D�1}��$M����gG�'À�L�.��mw+��1A�izm���iI�����Zu3���q�L_�uNQz�?�˂p!����[~��Gt�k��)]1��6���G�|HU��uc�S>��2���<� �"�G|ܬ>�� ��IW�m���.s���G�4�=����ds���n��A�������0R�n���6���E�F7��N{�r��"5��yە�f�a���0\+�a�1E���p3�^:�Bi�JC�g[��+�hl����;�GMƟ{(��u���qu�*��� i� g�T��u3{�����dLާ���c4�H�kkOv�#�vڃƬ�Ęb��7&������7K���0�(��B�h��yד�b�6��}CG��䧈�/8����\@Q64$�Ax;a�c�x24|��ŉ���$K��Z�io�W<��k;5����N�K �{Xz���:&������æ�FŦ?7�����U�ځ �}���#й>��2\ɢB���q(�U�w���PbD��[��:(�j���m��_Հ��ݤz�����DiB�q�7��c�ܶ_��Q��o�I#��~/3A皖!��.+-]�Z�vV5+mKHl@�d�D�����>�f';�k�ݮ"N$���F|�V��jY�$�J�����5 *�����T�m�!V��)1^x&���qȰQ�=H�b���Z	�Ev`x�hc@�|��v��m��4Zn����-R�䇕'��K�W%5�/G�KM��OI(��ն��{oD���C�������9�K����;1lj��s�n�9�l�����5}��
�7��!V���x����Q��rr���]�Ǩ��N��>����$b�hw֪g���%7�L*�pN\ċK)��㯌/Х)4��������gZ�/�JP���]=@c_��0�� �������
�#�o�<h���O��`= �y#�8Jxȫ�}(BL�Yދ��X��(�٭7K�pxuV,���)�Pz"uv����Hw����z*M��T�{2g���o�""��������'S@����(6���l-��q��iY�W�+���
�:����2p��J):��\���kD���/\���EO����g��i</�q��.��Z��mͰbk��-�ǭ�G5�����(��h��(.bxߴ�cyNX�]��m���աwqr̛L�� ��ݶo�i�#<B-H�]is30s��,��r�R��/��س�$�.��_%*����k�S&�JW���)�ʂx�ts2�i�`��*�?e����Z�,2S��]��K�t�΢$�K��DI۪�T"Pv�\�����%�|�z!���V�����Ja7S9��P�P���1@d���X��9�[qSu-~�����1�����O
f=9&�~�λ�ǅ�*ջ���5��o�=p��������s;��*�F�w`�t���P�[���2�M��MC��PE�b��DC�X��ˆ�;o]�
����#S�B\��6_;�=�
c��$Íڼa>(,c9�{Y�Rm.sd<0�������!���ܘ���.v�<���F�,vV0��顧�!�mi�InPZ#�6�j�Sb��:(�U����7�h\���Pػ�G�"�BW;'�LJ�\��YJ��w��<ٻ��e�J���O����� k`�i�t�b]��S����{\���z��?,����8�!��$Cr��F��pO���ET��a�U�JSqQ��s�u�x��R\e�$u5�mDFUM�a6ؠ y߁Y�rKP��'�	�O]4�W��/��F�<:C'�<㡟WV��8�S�Dp[69��ÿ�NR��m�$�����$���#�}.B(��>���:hw},�b<��e�)!���'")����i\g����@�Z��A�ݽ��;��.A��.�;�ܽ�56s���D{=����q��%�!F̥�?�c)X*�:�t��`�Q"�ӽ���ސ}-��ƚ�bp�3t5S�̣e�S���<�jR�;^��(��w&\��3��j��[��6��kV��m��1�TЬ7�����Fd��G6}�S�T��qg Ώ��@`��\�_hy�(��z	�Z�>"F�Wb?*؉������`�'���R�αG�8��.�����L�Ѩip�$�@��84�yC��;G��Hhx�;�*s�X���f^��ŗlH|.��5�`O�(��*��-��t��R�4�s��O`)i�3�<,b�LƸ�x���'	�P��/FOߐ<&+I��<`�q����5X�_,2
fܪ-o�	"�sê/%�=ƠLV`�1ݸ�.d�Ժ��H˴�tI̧��9�󩶭L���A�z��<�"��g�w��y��W� ~bǌ�&�r�Z>
;܈��0��+��O^%U4��Y��뺂��a��U	�!|��-���ߝ�\y->x.�CCH�����>MX�܆�"�H���p��[��'�ܓ7.�lGy�p�<��:m_��-%�p��M�j9��}�^����u��ޛI����F���0G��K��g�bhi��U�@��i�3TjP��J왷�q<ה��>N����5Uˇ�[� �h?}TB�A�U�X�o��rU�E@��l��sM��[eP�0S��dqG�Z��=���ق�ӣ-/�ޤi�B[&�I�T"/~�����<}�W �U"G���[%)2�.���W	��\�A`��Ɛ�R�T������kqGB��nT�(��j�)[��ϔ�"*�cw���g*�Eb<1oʂ�̗�٪.BE���G%,Z�T3M���*��
���֦�CN��DT0��ʅ����?�}�=!�N��5���~�S�`]��h�=�{1��4�����;w�f֌����5���K�ɘ�,���7��E>x�j�ESq9�o�+̑��7j�_��S��L/[y׸�>	�u���*]S�{��xN��sC��8J;@d�6Q��6j�d�%<	�h�4	GqX�|��t \�J�fE����f��0'��3#T͌1�����hI·0�p��$C������iޠ%$2��`��'FS�t�mI�#��Λ�!��:���ӞQ;��x͋�#��YgW�fb�.)�f�}8�/�XGs�6����q��J������l�)[p�:�
���r���Y����>����8 �/_��]"���v�va%<�ǜ 6��<s`�	����Ҏ�V�����
���e���<�<��xs�%B#WA¯;0o����JB+�ʭ� X�������C|T'�ve�21���9�*ck����":=R*
��X�I���bz0��ʚ�n��9�7&U$��X��؊���M�*\��~��Γ)c�l�xR�g��$����;���P�*z�h6���~�zRî��H}���ՙsy4�|O��O�&��� �Zi\N�w���Vq��#q� z�,0\���ĝ�_��d{�[���sN�[Cv��o5��-�C��oS��r�=��ۇӾ�����K,-1��w}_��+����(ӫ>G\o�{������_�������мi��H;�-����N��i����P��J��%�3��_ܥ���7���`��#
�%^{�y�"B6��`�y�fa:h�0`魮���t˱����]I�?a�
��͌�����.�<<��괔fP�υ��]��r�QY��3�4�!!M�`�:��/K�y?p[9�p�ݠ?�rE��qp�(.\���D~!��4x���-/��T�Ѩc�w�$��SӉ��A	��^R�MWa�*�[��M�6�-�>��VϹ���w�F�A�qo�^���f�`B;[���S��u�V��aw��3��e��Ш���y<���< ��sa�Ã��`!�����=�с~�nE����'�͸:�[xrzU�ː$ ���,��p�aA"ݭ�.X��.;�Q� ������\ȝ�heٿ���?`;
IV6�D=i^W��2LD8�6IbU'���9OR�N(�yx���΂e=L��en��ˢ�\�<Z��N�s\g����k�kLc�4l$-k��uDg�Ĕ��i��}���UJ��6��*�����������⺅}-�<��vc,}���U�͖�*KM���3-q�it�Pa��j�\�� 	-Itǈg�C�ڰ���P�E��~ts�i	��G�#]4��3�PR�0V�O�V�H-oZw�jdWn@�\�]P����",b�h�u�������/V�ʵ�{⫅+�l����U�G����`�)CO	�;;mHv�v-���[�!��	�ؿ��;�S?4LI���.�X�Z�f�MS+�x���V�𼐖�_A�H��T-vv�]3y�J�H�יu��]2y�ȟ s
ج������nr�6>ʭV\濉,3Ug���d7��#RȨ�,
���69�eJ�]˂&[���T�NC�K�[�;u�K�x6�8r�*��P�'�+�^ǋ�LT��h�Y���ݵ�͊�N�3�ɣ�^(J��[��7@K��6�pyc�*�ϻmh渟�L��Ƶ�=>�K�G߉_� �؛��]�V6�����x��},(C!he��tbt4w���F~�x�&�7�F�ʩ�n��W��#�²W�L�n����&1�(?���]e@7?�7��Bl�{5���jg׷����E`���I��.�bv7(�L���f��QL�hv;�F�^%`cu�.I\՛ڔG���A9�x}����?������:�i���N�����J�I݇�n<�ě<F�-L�_䊭<�
��.�D����<8q귦�3��r*̡(�>�؆6�I($�D�x�]*p$�?^&:�����4UQd�9�Oԅ���-C8�h�7r�	��g�`�(�����nP9�&2�1nh��{B�낽o�^�v�ʵsO��H"j��h��ˌ���3ü%&�	��l<��[��P�ݗ]��V��ǉ���=%���HT5�R Q�ő�!�f߻pi
���Ƴ%�/@jB����E�� 4���\@����,|�Z������K_�f��+zK'v[&oU	eM�8fy�
�kyphg��u��/����4wH�9�t�{F(�w���,nO��:�]՝�3�v����,}����M^�x?��*_5fI%/8}�b���h*���!0)�x�-����ո�iT݁2�+���0N�*���y�z�>|5�0.�B�e;�j��ÿ����ځ\�Kʥ��W0,��k\8=(?����~��U�,��ar��Q���j����bf,_�c^;�Mš+���E�1��)�>q��E�� e��6�C�W�T�j�9���K����s�!.���Qh w���u@VNZڼ��7CҜ�8`eL6�D��e��ټ���RN�fV9��j��Hy�b:q���Q_OP�0Gc���&�1��Wb�@ԋ�$�~#,���ں�����UD`���+���M@ew��Br�o�x��@��=�J�+�)�K��1K���m�q��kY�/��|{�?�>q	t�3E����EK��<`��+���V�i9�kB}�A
�?Hj-��l�6�e�Њ���r�W�8�sn�T��� |..�{[�ݜ�SSa�y���鲢>4��^�B���Ib���w�{%�^�P�DN�;ƟeE���;&��kfFѰ�$9�&�T���4��d�t�(Wms�y|�U�Q��b�-�I�}�Mq/<BNq�&�*{�a���ǜ I+iAO
��ta����J��"Ｌg�H��[�pr��X=���c�\)�gx��R�}ԓ��O݄EpS@�#?tcj��Ӑ���̮��.5��)����5@
e����9��˺0����Xk0=u{
^����wco�(ee��u�V8ͫ��� ��'�"�(J:���|� ޵¡,Gh8��Eqɾ���7*����>z\��a�w�z�śv��(5iV-]��ŠȢ7U�強FL|�ˎk��,�^�kt
KpUb3<8d{���tD�xP$�~��$0���"�����ES���^0�C0I�f丧��NI"�I ?��8�JQ{5�:������vq{[�7��X�`��0��4O�~��Ae��k�N�6���yekԱ�O��vܵ��+��m���Eȓ��n��#����s�l ��H��<�zʔR���[� ��H�t�8�#-+�Rl}h0C@�q3��t���ڠƱlU];Y��'������i8'�aa�הn}V@���ܶ)��l�4���K�&��Rpk�9{���L�������cL���e}���5��J�y+oX��]�Hsa7�>��$-���F��emW7	k-a��yk���U
�/��������	�sF�U]�x��z��\�\`k�U��p;�ݥbz���;1M!@�g��3���,���h�	A���ژnN�Q��8����ߔ~�}��|��p����0Z�
�n���	I0�KM/�j��I�����0G4�^�������~����-��s�-J�F+�̀��K�����j
�T��x_�O�>}��q�`a]Q|xz3en[�������q�Q��l:2����:�~/��M: ��"��/2����y�	̹���[�&:�n��1re�>�h���LbY����������6m��C�4Mٵ"g�v��O+@d�<�m5=�̓;&t��ڙ��I����`���퀷m�Bro���A�Z�2�͔ǭ�Z��>��\���Gne�B�'�S����@'����k	R�I3���(��1�����j4�I_~q�Æa����2.Z���0����G�S�݀�]��Ո�Q�ҕ��~FB��C܎��G�ݓ�����[��^�	��R��RS|��N��Y~!.�p����MkF����[��V�R��������]"�دV����R8{r9���\�Ї7%�,�����}(��o��P���S1L�tS4S��S^��qZ�t?d�$��RO,�u��|�y�n01���tZ)_�DټF���d��:��,�׫���@��8���g�.���
B2���֡L9%�����`L�q�{L��T2��l�"�
S4R�qd��~2f�e�~w�`a�T^��v�p�&û+�58."O@۲�RX	ϖ
�N{���"QN����K�MA�^2p��D��  cUF���Z}�B_�st-���]���Gg��˸��!np����N�y�w���L�3�ZO�Y���Q�Ŗ�§�I�Srk���*�K�)[�K�0��w,Ѽ@��bY�<����l!B�@@�F|�~Z�)OP���~�6��pu�aR�I����I{�fkX������g���G3��O�XlO�pM���?&� ���{�U�#�3Z!&���O��{���в����k� �Gb�k._�;`pm��V�cv�F���rRx Ո�j�|>�����ŅF@*!HC��&�x���86?y_�����o(�W.ۍ��'D��V�Er3�v�Qc*::$Of�#��*e�v% tЬ�W �,�xY!�	IK����VN�I9����0G ~�aE��<�t/��s#��S(���^����e�.�S��O-G*�%�������#����u�m�-b=J��Aޅ���l�r�M�U�P�'�.7~�#B���3R����FO��v-n��Y�6핃�@���Q�&W��b3hEa�u��0D��� �Pʪ1�d���+�<o��3�]�����������<�#��*L�p�OG�"D���Q��I����
, a6Q��Q1#>U���_�oO�;q9+Eھ�a�|g~�l-��҅p{����ܙ��z�P�K�vc�)�nE'�������&-|
�Cڡ.$����=P�G#���W�
'=��>8��훜�sn�R��7(hh�^W���d��ĳu�d�	P��p�ޤa�gR�d���Qɋ�C*�4���ZdL�1������ْٔO�^~;a�3	}1�{��]O��������x�����t�+�!q���h/ ]epC�}g�$x3̏ˠir�T�j=p�6���M�RV,��C�3pD��A"�9Ԙ����H���I���U�"�Vj�_���Cv��EB�3��K���<nG��qCnh���'�B���1��_�2�(1���������;�`mTs�� s�r$��Vt|�=X�h3g�9O��*~�䷎0މ5t&f9���6h*lڀ�
i�o%Ⱦ��$ll���O	Q��z�&�����$(���Ȍw�~�1A���B4��?#x�-�F��%95T"Ӣ%�&�t�`�%��ˢAD@�W��~���;n:JE=���H���-����f���l�3�����B�B��|��Z
����( �v�(e)R�z�l`[8�$�F�i�[��w$��}.Hw���i�K�=��Oy�i�7(0����f^��NbE��^R K��Ȱs���"� �R~�btfw{��M��h��뢆 �G����,rn�p������������k���C��	�(�of�\@���G�06�ܙ=��N��r�d���f�����M�����#���Y�=��=~��DN�̳��L$���=����P�N�X9¥�� |��d`����%\����D���p�)iVK�����A�B�.J=q���_�:d�C/�A�Paa��:���W/��Q����fգ,m�\��a�_i���q���ܹZh�*N;wo��C�f�aEtR��9�<?)���<����!f���ݘܭȎR����<v�a�7��wۊ�>�,�w��<�7�M�O��6�!��"d�a,�7T�)����3n���a�^�ؒ���bH�6�U�I�K���8����������{�k�)����0�F�]��u���0,�"C�V�K'[����A�"�X� X�+k�B�ќ��bL�� �j�<�DR}Y<����>1?��?������b:�8�KMǰȧ�-�"i�i�M�nߛ������L�Uy�'�� �����!���sL~�J�/���*4c��3S���jXH�֠��T��X'�G'*��g� �=?����c�[A�O�aE8�YxOh��h�ߓ�I�G����k1�4��vO]��J�8�g�T������q����� ��%�c5=O�	�-�8$��h�T�S�S��0J�r��iVחC��T�:'����NG�]|9V�E�J��<ֵ�M�:�p�:���1 ��P4��L���ˎ��}S����ҙ�y�8��I��8��P��w�z�5�ئ�θ�J%��1�K��f.7�4�F�չ_hk7���~K���T���/�yQI�4+m��m#K�Z,��%(� �n�S�X��
��w����py�
�]����&�j+40�4aq�fe^�eM�Z��W�J��}�A�@X��$�^��Z�A�޼�ȍ���L��!͛e@= `���ԯM��Q]���d�I�4�7���Ͱ���I����ߖ�bd;gҫ�x�_�f2mJzA ��Ac��G����cs��(_��Nd%���LC�����	�qAB@��ŏ�h�:����D��Y�?ϕ޿�w ̒|�&?�El�n�m�<������~�1sEY�?��o)�f����tl`���Pyd�J[�N#75���;ڒ��Z ���5D�߸��3x��сt�3�eXh^�iM�����@y�-��g�	hi�/�A(���s Dz��wɮ�c�`l�����]?�?{*���Wn1(�ѕh����d}P�.��-5Bо�+WsՔ r����ʻ����4�k�y�|�L!��A.�}��[q�9Ԍ�k�+mO%!�	Ò<l}t9�Ds>��/�2��H����j{���r�� �\i=�i�F�x���8o�*1sǅ��>)�*�֝ĢCS? ���Z��!9x�}��� ���9Oc��T����������x����XUV.5����/D��̂�5r{�I�P+����3皛Sle[��#v�G��K��k�i���jB�$@���' �x~��+^F�,K^�$뤥π��\Cŵ��>x5T�/��ro*���֎�����aF�(+<�۷gj�Ȥ���e�{\�S����TH�o(�:(��,�#N��Ǩ	֓K,�O�c[�ߞ+*�%�6�ܲZؔ��
�U.a�\��s��8�D��_�_r|E�^0�MC:� ����{$7�t}J���*�#�M����׳M�U�N��s�R#��H����z@]��d^	��0�e`h�{�C}פrRP5�2����X2���}^���tw�{dIҌ�n!�_Z!�eň`gq�Ǉ|����9�������r5|�E< �����}R��	�'�!����cd]8����b�/�2ʜ�G�h'�ͧ���rG�����!�QO�݀�.��� hYRK��51N��~	�ǖg{��AҕV~sK����e���*^�8!� wY3oGxe[�,��n��@���¾����\5�fe%���u�\�7���x��uʹ�܊���	��c�D���Y��jP3��'�Z(g��Z[�ka�b�:�^�c��
?)Fx�����'GO�MM3�$"����n/O��
��{��5s�9"�nSz����8d�&�0��9�W���͑q�c�"���F]
8|�m�˯�nqF֣c>i��FXiQ_ё�c%��^�KӁ�^'���O[�˞>r�5�Z�=>���F�m�j�^�sP���ѐp��ü���<:A�{��4u7�{�� �"�K��4�F�����D���-v��G5.������h�;Џ�!F�p��.rC�U0��]���d{��!����k�ud__3�2ت`
_�����U�k$iA�#N���q�Xz�8<b�m"or�N���^w<���GX����e,:v��:c,�
�P|�c�(-�lC���V��s��%���caXj���R��r?$a?"RJ2Q�zJw��� ��~����Z7/x��$�Y~
�Tq���;7��l�5dMyc��+"�v�뚙�*�L��'���ĵi]�x�)kVSZ����1Q��6�o�4���zl>L��8�Pi5�����(��o6��.����T��,)��������.�#W��vA����LnJ�D~�vڧ�C�ȧi깢�3���2k�*�i:ta��}�Wh�3cӽ/�k�x�IS(_�0CL��# �ۘw��}=/�����"��ǚ� ��ݍ�HR�,13/�����q�l���0,��:�Ah��
�m������
���Ԣ�.:|z`fv^��"BA��h��DP��}|����@�2�����0+#
RU��Z�8[Z����k͡]���+���WCbZ8tb��&�;sB׎�}�
��#D��H���׺OѮ�H��ƶ�&���������*8��� ���+Q��fO�;W�}T�px�:d]�@B�{Ä��PE�@��V>ta�K@�k��D���q��t����;S1Ų.u,	���i���DgO�(M��LsR�j�h*x2�}5t���K��x@yn̹�\0dߚ'���oQ�ͅ�CϪ�|P��X�`A�1u�xȎ����k�A%��]�Xڑ#�|�;y���mq&u,6$�����L���qL@��XŜe�W�r�+�Ʃ����oIwt}���J<e�c��4e�ڿ���aRBuCv�^/��;�8G�rnq�$�	g��w|�e�̷��#��E��X�Mc$�>V;~h�&�%i7��z�2�v�Rn�9����㒞�q."�"�Z�uT��OUn���J����`�:#|=\]	![�&�Wvki�~�	�rF�z�>�>�= N�`ϳ�n:�����]7�!��d�Me��{A���9�]N�h5��Qt��o����%�<f���`�7S���j+�c��X�J�	��Qս72�}���g��z����-�0����`�8Տ���`�Q�1�l�����w�?tƄ��H-Y%I&͉J��C�p:s�J!W8�T�EQjG�:�7b��\4���bF\޽��6{>��%v`a��7��q��i�)ɣ7B��G��>R�P��<x��xBa��nsSy^ڣ5�G��r�`F:�ѝ�Qi�o�+W�ȗd��<�<�{P�M�� u�{���"�2=��ǭg@F�pK;����X*(eK����ؖ>~f�=~r5�+z�f{O�dN��F��H�mO�"(�_���	�P%�Z9x����*b�����GF�9�#���
cX��
���(.M�b�m]'��&���װ��6n󡇩��ML:bJ��Fr�͏�hPP���b�T�����no�f�����Ϩ��a[�g�)�#J��A�3��HU^`�q�=t4���a��ߊ ��k��N�����%��/ �6������Nݝ�*�nj&s�P6Z���WC�4��F�E8���ګK�u���~R/�
j��,1Y�!^��:�\e���η_���?�g�@?6IBS��[6YY��E$�z�Mc�t�����⹦�Y<���+��`��Q���j�m�9	[	���]���E �~-�w�u5���#۩�77_g;�_�����\!JB5y�k�(:���@J'Шf�|J�qxU���cY��q�p52��SGi#[�K7t�k�I�aU�t	|{	|��/_�G�������X�^Ӄ�B�d�LJ������j��j�nqj�á̋��)��Tr�7f��楂�#��ayFF ���[�-0C�Z�qB�6J�Woָ
��bv+y�rb�M�g�2 2cf<�N7�e�$�s�U��q�vE44e)�}��,����9:Q(>�*��^\�g "^b^xe�♱#����35X��<���[�6�1�d��k�����6��R_߉�x�~0��G�mQ����e�����a�����,;�=NOG48�??~>�Sd���xmlT>�����;�� X�g=CC��Q	s6�U��[��҇�6t�/~������~��+�����qRF�:h����[n���-;MI[�6�FG�	�'��l�,%�U떭�k75<�a����D^�+�s��3��D���H	;��:ٚc����
��b��\C$����V�jӯ����\ViP�,F��H���6v�����p�(���|?v6�-�,X4=��%���r�v���#C6O����}��E��I�?9�eq���k����%���ݿ��E��xhaĴ� ��	*��J"�#�,�1��l�/���B��4\�p�0�W=е\Ƹݸ�O��F�\^Ң��1.1����4,a������/�Ѹ�=�f�i �ʨ��'e�������-���ask��B��
~e��EB?��\2�MR\C�RS�UV�\[�u�U���篞Nx�#���J�TG�""Xh��o.��ᝳ��biH�U�� �ןxm�se��������j����7�+}Iv�|���W�o�ߔ�U$O�A~l�����]Cm�*�����^%�hc�<����j���M�~q����#��9�;�v���]�����NQ!�{��C5���ܜz�l��s��&�������(Vl��gC�>�Z��<�<���QM�VGJ%��IR �����,$��h�F���ɢ��u�J��Z{��/o,�v����~�ޕ����Ac�^V�#?�� ���*���)~�"s���ovfl���
��	 ��/�HKVQ,UX\f�ɏ��b!�9�Hk��W*b�`��T>(�'�S�`o�3P��Amk�V�&��J10v��vˣ8��>��I�L��msPŒ2�䉚��/�$���Y �H#L%�Z�����K��f�6�� Y��M}Ş�^zԸ����2lfc��"F����;t��E��Q���bF/�֠�7+�Q(��B�+A��k-]��N<��� �TH�?Z���=���� D�T�=.d1���vD�7��#F�$����C�c_J������nx��ʟe �i��y����c���p�Q�@�d�{c�����C'�4�C6�U��.r�m���asg`������Y���4s���pә=ѓ����wX�I��5�|��-�-7� 4�q����蘌�8����>��j�$ �-0��ϓ���H�M���b���=4'�P��z��vɺ:���Et������r���̣�qt�
+���M��ǚaN�!�	��kHNҸ������5����oS+�,|�TZ�k�zC��h"�nb��Y��Ď�+0�z�V�X�
������ܤ�]���
�E��6�>��b����c��*QH�2�g�ŚD�<+�]� 
hѿ�Ҟ�uB][m��ɬ�ډ5_����l�O��2�$��(h|Il��CNqO�W�&ڿ��΁������y�Ь��:�l(�v�f�`�-��%PR�r�b�����M��/6B���2.NH��1��d�~���l���:(�"`�װ�f���Ja���V�F2���;|kb�o�\�C��9��F(ׂ�c�A�,�d�S0���H�58�-M)F�"MV�c�G�[���������8����P�Q9�H¾�K�2l{+�Ya�U�u���¤�U�Y��w��T_�X?gGiY���[�aJҟ^7:l��Z�ɍ_���$/��N�<-�u���(M�T�~��,�ٽ�t6Z l��W���L�iE��Q���w�m��K0��:� ��i�w'ᘿ�eMR����k�88
%��$�EN����N �U��wCz55dBz8!�r�IS�u:�g�F�A��O�e��m��Ni����§n��6�IrfaD^��;6+����� �s�?��S������١��)d�¸����[��+L��4 2��FTH�Z��C��x� ��MlR�,���4;�.Jd<�D��43����t��L)0't2��_4.�
�lwq���d�&P��ce�7Q�	6�kI�h�G��hZ�Y'�1rl��y�l|�O�#�j_R�#�K��_��daq���t��J�Q[��{+���I̛��O�2��AU�R)~�`�����ُzq�*"%?���@�`�dqa��A�. xS߽��Ɗ0�v$J��1�K��;��?n�'������`�l��A ��#Ʋ���!��4�}I�%V�J!>uô�Y���1wS�li7�b!�s_w��B-58�H̀�C�[H���EI�����z�;dI
x1�YT3֪�'V�(�pN�.�w�WI7�e��KP�n����4���G�;IH��3n�Z�}` �c�
��e���ہ��If���	�Y����F�X/b�mjv.|U�|8?���2��%K�r0��Ճ���o�H����Ν�GX$�7�2��a�q ����!6r{��#��0{U�!V��{mT�p��^Sg5jz^��{L�8d���	$��8��'qby�Е�x��+����q�+��Z�X\�,-Uji��E3(%{�\,?21���a��.@'_�~�%���j�}���!ᵲ,�S���k�O����ɔ�٪��*�B�G�n^@2g��vX��$�xE:�}�D
>&��u}w�Uyr\��a��h&ڠ�#2]}����"�:���,W� %�}.1hY��� QB��N,��`�Ȍ)�{�����鯬���͍�1�����+�ڮ�k���N[�K.�;�Ԝ���^���ɬ�|d��pg���-_�^�J��B[_�L�63��E��?��;ʏ?G��؞; `
LC����I�3x٥-ʈ��b������ԅ�'=f�ۋ��,��_��?�H��`�Խ���j靋�d��5I��OO�Wϻ�z}��xNG�կL����H:m�*i���9
��Ob��˗bT�uz���L
�`�rʊv!#H�+�i�P�4�@
�n'�.M��t���xG��0� �����X���""{_$ۖ8Hı�
���o�<=��p,��ٔ�������9��S���ch�R��ܜ���<��C�|
�MW��ZP���ҕ���1�ɦ8�}�}�#�z�M��JuQ~R;!�th�a�U������G��J}$��u�;޾8�50E��i���F:�y����K��cP�醼_�6	���ҴjFA�d$~���C8=$�)ȒƢ Ձ W���4%Z�]X6�t֬p;���c��:�:�b.̝#�҆���=��VP�-������M+�V�"ˈ���l���JE3�չ��3���a5��B������!Y�4\5M�MK� U�7�SZ�AJ�i�D��	�|²��6rA��X�h@Fy �vA���}"b�'4�Nۦ[�4�����.&����E��}.��ryLZ�eh#7h���g�Ӊ(=�Eg�n��2=��s5O���]��H"ոlʣ'r_��Qy[h��*�c�����q#KR|ʂ�}��/��&�@͞zѯN�i\.���5�"���N���I�P�%����E�fBRf{��||���i@����<T�b�{�U�O�d̮{BW�T����w����$!#ЈhJk��i}y48�b�7i����=�գ��p�B9��Y�|�C���z��Xz���9���u#�ΜL�w3taI����4$��R�6lU+�#���g��Zڗ��S�@� <�x�f���N�bmo! ��pI_f��)e�Aډ���<\��!���n���d� �*C�d�t�B�ӆz�ۙu*bE>�άaG�IX_Gd�w�����b�Q'�ly2)�`O&������0���㍎�{������K��+��[�qS�d���$�~���L����Eb�PmY�wW��ύ��Od�.����B4G��lʌ1z��` LDGR}���K���՝3���ʅ%
z�n�/#�Ѹ��~U{��G�@Ҁ�^l-#�zm}5zA&s�Ϊ�>@J��E�L����+���=:M���\P���G�	�dW9F��1x�T�g����}�ט=EV�V6oݼ`���Z�{��ˏl�̃v�7�b��w�/�����Y@,M\bT���C��r?7���_z�͌��V3{����&r��ys��C�����US���	��_�W�4
1Z��]��1����̻>�`]�N�FI������I2��j�y&�lY�'�� �TQ^��<�B�T�u̲yx6�^&z�VI1�C5O/p�n۲�B����r	)��~�ZQy ��r�D'�6X?��1�v �^�	���DŽ���j��
!�4��Sɒ���)A3�a~��I��!u�弢ƒ�"r6���"ILa�� <�&��P)��/���:Ħ"!�bg)��pjo�3����AQs�rǄW�VG�k���Rs��ʰ��Ӟ��O�\CCӾ@������~5�RՀڊ\����h2|wfH*T�G���B�/�*�L��&��خM|/�ʡ�S���kG�8���lՖO�1<��͎�`o�X��2{&|ڤ�D���0��k�:��FÕ��z���vC�ܙ�z�+P������I��+H�P��8��`=W�G*�J>��/������_��e�5_$u9�;Vh�T�LDK4���}te��S]Q�RxdZ���B���y/3�&��4&h���vH}�u@ &a�vyULtl�@D`���� �#]��"_����k��gsΑ��`ٸ����XD�`�M E���iÊ̹�s�tt,�����F�܉�ݘ���S�Z���GW@�t�??d?\]ia+\�*A���E&S�6Րȕ^��9��TiK�RAW,�T�g�����m�.b�z祖��Ȉ���jV�����CSK$�F�%��o�w�i;�hqv�5я���b5`6,�(�\�� jCj�:�a�S����5;���qi�6	�p{�kj�٠j�]@�9e�]�P�MB��Pk���z��X��KE	�D#M���K�`��t�_��1�%ú��T�բN�Bog������Q�|`�W�"
�k7y�P1+�
Pӊ�9!*X�:��N�Y��<~u�&���,�J�m�kD�U~�i��W����t�T�J�s����Uˑ�����yOMZߓ�IꁥL���$�/V��T�%�ꀍ)���q��,���`m���	x��"�HvQk�>t�$���� O�r�E�jj�fz��S�J��ᙠ�'2��]�=�p9�j^���m7�fEw����P�a�Bya! N��q}�nzw�9�&e	`-��hgѓ����)k�a�l:=6_F��ޭV E�z��������:S�TؓiH�IC�ȗ��s��S���KB�$xI%����UD�p���?mt�J[����%i�q#�":mq�����r��Z�Hbmt3�+(v����Dw�(?�J����\�@n(��!}B �B��eG�Tv�+Qy$���v���[e����Ҡ�mI����p.���x; N����D���w�֞�) ���5����r��VU"�m� �!�1ڦ�3ZRxѓ�B�`�����=�¹}���������,�:�jizG����P�ίՕ�6�):Bޞ�Y�n��5�d:��b6�q���>j�/oZy[G�c�f�����n�B�V��V����я9�_o4��R��k�h�5�Ob�L�t��'�����~�*�� Vb�Z�I�UC�L�\(�Z��{�5�KV�[gR��%Kl��.�N�y����#H���N�s��&����9쮌�����¹P3��Zvˋ�d{4c�)��A�c����+n�s�+]f>�)�j(�A�8RC��4���;�Q��j�^�1�s��-���֙ǐ(��܈��y̓��D~�i��i�����0B�O�邨o�e�CC;��'�O��Kv-��9G7D`���d'�9�$&�Y��.K��0�o���m����B�I�a
$�D�`-s�̻rN�S���fN��T��!=c�dadٮ9	\�E����P%�C�N�Y��a��l�����.iZ@.�����r �f��*�A�7#����n$<0�O���Т�(����K��D�z8!��7�Y� =��<� Q���
�G���,dVGB�r�����Uo���_O�o�j6�ƝJ������d���yZc��n�����uG�8+�5��� )�ƃQ�9�!�t�!��
<��wb����nn=JCHX��u�c���9�#����8�U�9��\�EH��j��G>��C�#ؗR��=�`3�����.f����J����"����~&�W:\^f�@����k�Cr��WŔ��z��H���:�w%b�Ю9��_ӋkBO�T�ٟu�\ T����LjcG��t�R�4���j{v�G��J���N�1�%���r�oF�U@����`5j&G�\�bº^���eyW�w��V��R�bf�X"3xQ���._B(�u�Ծ����6���Bޕ���g�$���C���&97=X~���h<���5lb5E��.ʑqf��L0l@$" vv!�8s�|D���n�c2;|"�S�z��/�e8|�%�Ig����diA�ێ*@����Y+�[́9���
'ϩ{�_7ٮ+��	gj:��
�8P�0���mT:a������	o�8P<f�Cb=�b�f��t�
n���[=(�t�G��G�g�4<t��za�ɤ�bQ
o�n��(fP8�7I��@b:!��="��64&�p�t�H�2~��4C�� #b ���Oa��k�	��he6�	E7B2��5�,���!8�0 �����ɘk0��Ԧ�Z����,ւ���+���@���$�)� Cy�QȨp��̿5D��YH6RQ]���j�F2��t�1�Z�4,DY����T���tˏ�Y+���s����)�
�=�!oc`	f��w�;�_�ZeZ��oIߏ���ʖ��G�B�yl��#�\I �{�Dͅ�q2y&�����Z�C=B~hr�b��|�u�m5;�H,
���'�2,QA�%#ã�rM�`����W6z}CT9��c�-�,�:,����9|�q��k��a�Nsq����i'�H�Y�V=�����p6T���!�֫F>�>�K����Ki=F��U�c��
5�{F̒�l��+z�V�A�A�T ��7��2�$�7� ��R|�C��,L�g�̀���k�ő��9��Ġ$)�������*�˝v�~�P|L��!��}O���4��;_F~�$x��EU��+j�^�����,�g[���Om�k} "YD���\D�C�ܐ��.J�R��n�8����]2��g'/���a�I�8�p�;�VJ�&���$����W��X�<���'�k�t7��(�,VB��?9� ����5�߱7�s������tm*KU�ǾEY0~�%AЅ.SGbW�Q�� ҙ����]�m��nQ�c��v����j�f��>�������{���ֳap���x��,{#����<�r%�%�2Ԋ�_!�8�T��y*E!���,����z�ʧ�6H��k^?��E��0`8��Gܟ�)\�C$�Z����c�d(��a�ՃLg��i��4�W47��$,����E}��L���!������ΰG���hf�V:�+=�W�3F���h�:Zl)�mG�K�8�=56B� ɨ��Tv��<c1}�~����S>���B_\"����J��"h?BC�	~���|e��Դ��}�h�ɩO���X��KA�G!V�v���<��0�/�tO0<k�MJ���k���i{1���V�KU�#�6�J$/�kA��&�����*χ|��?b�Τ>�󰞜t�2ϡ$�n�S�#�{+h@.�!�E9�?G�!M�OY�|�H����	�~F�۠�ڂ��!�z�=��%E��̳���8�&_�������e�ȲBM,��O�v�'�rP���"8R.�[e3��us�Y�����z��^Vn�q}�}�4h�W23޵�����������b��χ�<0s�BFk�m���������~}ᄫszІ@�Ѯ�=[o�����8���M9t��1��ҷ�.'B�}�p�;t,�RU�F<{�xr��O�%.��o�O,�)"����ۙuB�Z��X^r0x�`5J���~[�/��J�	���H,U�X�;ai��) ���Xi�^Y�#�?`p�*����J�t��Z�E\����C��¢	�+��)�@��x�������]����Ï���4͛��tU�yj�{O3�n}�֯-N	��U:�ڛym���I�~)w<S���퐥"����-4�no�;ghd��3`ɽV%Qi(�W��0�ug�+mOJ7a��{�ӥdoC#������r���Z$9�
�����	 ����CsӛL�NoP}(���W��KU��f
	��),���p��/{�m����-C�}�%
�\��	�?������� .�VTnQ_|�Y�Q�7������yWbt�{�vv���s���������g+��Ij[���G�i�d����gTI�{�2�a��'�]�=��f�����H����n��V=���d�P��O�]�1�S�l:�dy�H��_�-V�ٷ�m��&��9�zp���Y:��E4t��	�O_<D~:.#�n5U�Fk�;
�r���"T��x�y3��8E������9�}���Mi�c�����V�'�����{=��B��#q2ir���g%��8��p�]#�t
�|��Sf�t�u�������2=�����>���JD!�Us
�!xG���pD�/.!��m�����8eS���F�#y�Jjf7�tL���`!��: ��EA��A������B����f�m=et? �B#p���omr�Kxu�����_S���X���W��\���6^�g��>�	5�i��K<��i�ȧ�DT��b6�<�5�åy��p9�2:lT�����s6}�W.��!� D�h`��WSg�{��ؐר�k�����d[J�ZnR�&Wb��e>h��/�i��G�xM'x �y����8��{$ڽ�H_��H���ݘz�>7��?�J��*	�\���Q�#�k��Y���Z=Z������ �u6�}�XgE=b[��Br�c�ި(�X��C��|�(���H�_��� ��T��\;Sx	_�A�+6?ޱj@�0�᪤6lǘ���w���[\{ʺ��Qg� ����3�δ �ԿB���[�S�i����/M�o("LE���4L�D����Xv� �Zk�ֱ�/�gg�d��_{㖡+o������zNi��o ;kˑ�L��KC	�9R�����]�E���)��먘��(Z�#�Oc��o�y�f�F�s+�xG��u��֊3�{_�"N�dkK9>^1Kbr�F�EY��t�����m��#������/? `���m�^�>B?L�����z��(��ܔ�bC�u���}����v|h��Rì����a�)���q7	��"}��� �,F녵�SB=�fR��/\eМ a��aK-�3LC�4�"�M2�96:	�2]��|pC�R�煣=\��}_4�Q�nCui��wP���2јFJ)a<DLJ_�p��
�x�-�'�P�MKM�BQ�ۤ�-��`�	��&�k�,�pD�����/�ן�A�B
�I���E�[z~!��Q ꎿ:~N$�B��y��r�i�2�;k��Jg��pc0�8c܀�\�-�b;�F��L�F/ׯB�($��V?���N�W@,��R����+��~��R��ج&���L�s����2*�5sK��ٙ�a���4Wݴ��T�����I�Ș㛢y�A��6�]�i_8��p���QK׷?B F��&jϚ�&B��#Y�We�6_�@�-�Z����k����j�ǫ �KI=�\���'���2�_����i7���D� ����Zq��n�
S3�g��X�O���u_�#���H�72����E���^@@k���n��%�l��J��cMl"5���W�0�0B�%�Y� �e.�dK.�u��<��E���y.�)h��Y�>@��Ő�xĈs`J�o���M�w�aRx�NoZ�ߊ(Aȝ(v��sz��s��ya�1h���(�%1��g�����,�aG�Dk4�?��(P�#��`�|�\�A}��0�jp�?���dL�������)��=��b�rݜ�q����n���YT�yi��JLt�q�0�&cR.|�i��D�p�{�ɉxHo��3@Z'�#Io8l������ �X�7m�8��J���;�Kُu?�b@����A��$Z8���¢ ?�l$$�7���=j��1�73���Tg2�bt^���π06 0�(X?)J� 4*ୠ86j�Ȯ2Bd������M�+į�;tTcS�f�ǖ�#"!����d\�w�,��p[�}�����A��R���s	�i��0�ݨΉ�g��~K�?3�v����Ƕ�ܟ�k�4[i1�P���2h��@m��z�� �e�G�Wg$�y
�.��^�l<l���f�9� fT(��Z^��N&�8L�L�t\�d+3�\s�T�^���WMgM<U|����U/������|!c�*�s�Y�o���l���Y�V��9n��uH2S��0�#i��mK��������:�����DT��kÁ�^��J0Ԇ�]d'E��<�4p��ET��p��O��!w:U5FZ�<
�$�ȓ4�D�>���:�*���x۱�y�j�:��ÈWՇ&M����/�V�ơ�`N㑒��`o���!������4�x���:�`���t}l��cD��\'@��j�u���S�����3��M�g�7�8B�;T����vd�Y���+�ݬ2�
��P{\O���6������A��n�;>�+�KqT�M�����6�~�����&'�9�ruv؈��z�!��r��.To���Tx���,	t��d�	��dc`�P|3��e�9c��]�x���e�X���N����$�u���_[x�|�ŖX�/�16�ٹrmύ�1h����;>s����k�]f����W�,>y��b�Ԕ��2��)��j�t�o�$ȏ����>s�1�IL�a��W���K�4�}(�2�T��q��ǝ��zwT3�ϴ�$� ە��OYR� �� x!s�:�-�ɘ.ۚ%0f�1�n��@�0��?�̨$�_�'��[wE��\������"���vs"�:۸��` ^i�Ź[�A�v��$�	��.Qa��LjK���L#���KZy��Pɯn�*�A�!=eB=�9o�	�%���.G�Wl�w�X[�J��g���5�s�������W�DN�����\���M��#�=|YXҦ�D_��)�|&�v<E�i�]�@����LI��	oq�H.A?�{OC�j���b=w��2^+���a����@�?�~Y��$��ųի���Z	0-��p��8�r�{��u���jf%l(��)q	�/�y�Yɯ��BZ.v�M:/�ia���!�Awo��v?�d�O�Ǌؖ�6�T�0�R�	��j+w=\�P6��5�E�������]�[j�*1�j´��9%�k�ll���1ə�!'��d?6>�&M=0@J�#ssuz|�
�O�P�R�P�B��Yix��8��@GLz�����ϱ��,�-��;L�u>x��U{(DU�÷���>�&��K�
�L�ĺ��Z.
ޢ�B���������k�0R+*����I��d����N�o�_]�J�!C
��!������ �*z�'G?|>~��Rpc-	�n���3�V�2m��Y��X)e.�Hk	5>���٫a
��'�y^����{tlX�l�͊��D�Nڥ��s�{y��������s�u:�o_)o�k�5�ES�)Zi��d.���P�؊ߑv�T���AT樊���B=a-��C��ZbQ��&��4�l�C-m�g=���w��LI.k�B���8��)W	K7N��6�&K�Vl�<��M�]!������"�e�^�I�=T�`)��`���=ƿp�u�:޵��(���M<�+i&c��N��j�eh=9W��N��my�C��:�8����'�������8~����������0�o��J������nq���+��s����D�ҫ ���E�W�uK���c���[&\a�[HK	�EW����R������~����<�����]o/`3�O�0����V��r�>��ۧ_̣�׃��Hk>�I�TB�֐)d��͟±��|V��%	A����5+$�Y/q�GZ�Wk�)>Î��`�i!�+4����,Ó�yD0����k��r�h�c6L4�����hY��9��LM�D��Ũ(udg�}�FK9a��2&߃Ƀ�3V����^�i��L�}6;\�čY�f^]��	�y��Ψ�u�)G���V�c�Hv_��SO Z���M���@�B�j��!v\���MHk������&a�T��"��1��E���Iȡ���1G�YaQ9rq"��P�U~rY�oG��[׉�б_�Ut���'��yRL�҇�ld'���1�6@(�
A�a!韍}�k�F���<P�(�zS�pX%QV��O��`�!���%�T�Q|��m��R,v�J�C@�x/$Tu�̠���z���@��p $�&KB���c�\$le�<����s$F�,�U�.(�*U���呬��8JZi�T>~AHL�ʚ�D�G&mj���������.���c�#jJ����[
�q�S��ݍ�ȳg۲쉘���Q'~O���j�|�G瑯8']|T^�*�ή
r-�
'��Cx�9l� |�;pS��^����@�����{��s*C�/�Fy��3����9�[����#g��8)9n���w�_�K�kxY�Dr�*W#T����*V8I%����ة]�������r�����?_ w㞠~��P���A���UZ:���
�ez(N�9<E���tn�XE����}�M��xWV���rB�O�r�A���.dW���Qx�����!�}�!�Mm�-��I�u��:�� ���Ud%3�#���*�u��MBS�.@���@1�է<��Iw&=�˙u@��ޗ�\�'"[�o��M�T��'Yv�j��<ݎgx]+��i�?��������5K�O�F^ȏ���~�ڀyD:��(�rc�]$�:��y)h���'���e���C�c�'l�x�dL�%	����]"���	@r�Z-�����:UW�U�n�w�u���u���{J���Y}�"��=C7���*�w�nM��q\�s�~�+�i.#	X����mX�j$���	�����/p�=$�"�=L	���1�:e�G�K|R�nD<��{�|�E�����@H�����3�hV�KF����+WjP�rNtd�U������[VB	��;(I]nۅ3�SJ��}[M�Y8��6z�d�J鱗�q4�/���3�E�� ��##�v3n�5+z�pc�2��K�e��R6)�9�BfZ.�GU.\�	��T8�hs�F�4�u�Vh��ߨfO픟ۯAGX���v�m�3i���|���Am�8��Z����`&C��It��x���0`G�)�\d:y�Wߊ��I�t_��"�Д��,�����#�
������H 'xᎡ��ྣ'���r�e�����5�,�Ւ�씀���H�CK��`���%d�w�ҍ&C�����Y���k����3T"s��w��N����+�wt|�2���H{��Lvz���\�L��M�K���L_��<U���ܯ�JmQ�H���l��l�>�\����t���!����&��9� �E�}������9/"���
TG����o5_�$��̯]���9~�&4���P	_j�s��+Z��������\���p���N'0��k�����ELS�z�U��r��D�TK�2�!_
�㚊��⁀砑%��c�� >��̭v�T�l)s�`�8�?���h<`�N��+��-�8:���~O� _���'�Qz�Y|�z#��jF��v*�ڠ�U�&����pƮ�K�~��}R�(X����5`��o���``UW�-�w޸^p�,^�$��&P"�Y���}�v��VjJ���u��	:����Z.?g�W���A�=���97�����Ӻ��L������#vS/�*ȅ�ȇ�t��e�~v���]9:P"#��:�J�+��[/ҭƝ��F��!n��rX��$��a�jj�K����T��@�p[���2ށ,E/��ꬡ��]���1��l�լ� �O�Z��{A�-b�Q�)�����|�?�l�ͩc��7���ag���|���s7�Zy*��/�������8`�>�!��"_�T��������u�ˆE۠�064�&���s*h����Z�}ft�Oڕܬ�5���mmR�s��K�܋&$%�ގ��{����L4)�矶Aw��F̑v�����E�%~�%�F���d�m�����X���D<����&o':� �[3�����?J�T
�����6��A��)�nm�a������ϧ���{\�n$��>军S�$��z��?]�$��j.�8?%��]�N�����\iaE�vDw���e�Y<V1-�>�NxV�.�������A�+��٥���� ����D%�Aqv���fƌ�"E�ɿg���f5�ݢ����J#x�\K���h�/x�y4&�
����,�s��ƙ��5)Gq�\�P�橨3߽T����ռcB��4�)D��m#\4��R��]��ʾ�%��Y\��~)i8�4G�Cc�S
%B��	$�"�s��u���ԗ�>eD=�o���NM���2^G {z]�[*���>�<*���D��~��M�}�K�R�z��RW�����f���^�;���Բ?q*�g����&Ř��<R@��ⲻθ�/�R��աfc���b?ڙ۷�8���M1��Y�4�J���c'�{�3��d�c��������o;�F����v�T��?�B��\�z��s��M��`�5��L:^���!.����C�W��*���\KH<�0�����D�z�����P\�!y0�flW���8;S�F�^tI��2��G�͸�!zw>1'n��Z�yRْ�:B3����c(��5��ң�+m3�M�����{�MB]/L�@e�ɉ�_�c�͹�sԞ�/`�DG�)�Ξ:�L����-����7{X!A+�j��|lu�5��G��\ N��E(���7�Ca�^��`XWJ��M���r:��q���x��Z�F b-6	f�p5�D4\��8�Drӟ���86o�ء��6�n��S?���@m;��K�#h���}cZ�w<|�j*ː,ga�R�\�ͫ4�T�@5#�s	;�$�>��:R9o��7��m��Eq�8j�<�P�+Uh�`�7�y���h���52���B ��������n=�#��QoŎ�X�W6cU0��<�1��ُ'y���w	�~��>�$+IJ
�쏳�ڕ��.�褿��P��8}�l�n'��@1����e���F����UE�k6�E�s;�,R�vy�D۝��ф��7f��\+�]�+;3�yu��?S�+CE�M�OՐ,�<�t
���Qa��Ӧ��N٠t�J�|�P�]���T2%W&���杌i�,����W$�&��]����!xz�ni���x	
�z�,]EQ�;��	�'�AG�Ed;�:��@�_�_���gi(�$0�����D��hƼ�$�l3k#.�4i�q���S����n9f٦؎�����ŷ�w��Ds�P� [��3&?P�cD
úI%�� �%<��33,�a�6�&A~�9:�)��a|�Q�m��M�$<KK򐮗�����u���B�S�\[79��ĳ� �	�!0�Q�`+�jm7�\����a?�`� (\-�6y=��*I�؎���r|�%�BNi��7J���}b�=��d��=Zy2��\�4m��3W�1\��_l��MOC
k(�#�ۘ�S�UY�0?U�GH,jY����!�|���+��c9AUQ���#;KV�I�KSW�<D���J�y���pi�BMtQ2 /�����a�)�H֚ғ�F꽆�k0�:����JT�����-6��ɎDk����a@_�^�'�{Ν�XǷ�|>�񻟠N���l����sg�J|E��S���ekUx#��8q�������tdJ�|S�F_���>��pĀ��P�p�'厏t+A}-!`ݣE��pr�~��1�cug4!d�j��	�p��e�Y����H�j�i/W�v�t�����0�����Q ��(��3�5 ���Q�t�5��Ǐ 6�L/-YƷ� S��j&��뱪&>���r����@=�1����3�B:��d~w�Ͷ#��y��q&҂&q�7o(k][�����%P�ۂrثG��)�)��V�M�:!#�{|��:�Rn��6�`���z1����X���GDGF܀<ٷY��n��	�DN���;=��u���+��)��,�0�ka���H!T�S�g2�Q�C�F0\U�� &yu;�P&>l@d)}Ͱ%�S{9g� M������������<�WqE��Z�9>4k����;h��'���6^��89�r���Q?yM�j�S]��Gſ�F
�q,�mY���`�8�H^���}��t��<��T�p�"G�4�e��#1ݹ��b�HF0�4���-J��|ȅ����k;G���:_����⇻�⤶8��ԡ��؃r�(i�Ey���A�l=�9��P��V���k�����5D���Wq�1��N��/T*fܻ�;!T@4(z��r�g+|c�-ٳ�`<fR<Ҁ��d�B>T���p�c�����&����*v���ҾsD�}�F�^bc�����-�K�V�H��jT}L�� \�}@�i�1�=1(H�)G8�v�y`|@�.Pq^����ՠ{>�~#���2K�w��'op;��
C'Զ�U׀�P��2++�K�J�lZz+)���+^���3��۱£�p�����]q�����[��eI�y9��1y�Eg��([h=��=QM���=���� ��i��?��(�z(��n{"�����?�(� �������������s�4��띨�0qT!VY�IꁲL��b��#R��R\�fƙ� ����E���"�N&��";��/����=�^xP|W��U�B5�g���S"υq��u^�Տ%���������	����u�ưL��[��ʐ�C�� UF��E$�RdNO�W�(w��
�(�\�oK_���bƋ�\ uP ;_�G�2���Fv��y����Ѣ�p���w�:	�e���V��Η5P��~Wd ��RXBpqp�R��nP�c\�0 g_�I�M1�Jyd�"T���.1�O��{�?>L^d��y���m�wHw��),y���ޢ"2��R�@+0/ÿ[�/W�.�̀����wuJM���{o��[�/Kj	���|������@PA#��q́�il�Ҝ<&�'1�����A��gռ�t��+'89H{+s���`j�JA!/U��0(ut9e4P��3���i,�j�_�́4�`���[����m�5�X����"���v���T��Ņ�� ""'��f��;@��OR���
����+U?��0�Mzb�_P��.�,� �Ǩ�J�88�sJO����G)�^F�J8l�|�>̳�����*%2��?�.�|!���|ȶ��͌��;�"_r 7�DV	� �>�D��������rx��	}LdZ m4�%eW�������D>j���1YGnN�t�hp�o�2�� ��K-�o�N�J������X�m!ꐙ���F���"���FO��9�{� i��gM��� �8���,�L޲�rFҌ�����V������>[�$l^;g�#���߈Qu{�
A�*tr�p�$��[���t�XZ�/2+��O}H�v2�j+����@�p����xh^3��˴�n�c�Vu����j���\ñ�jH #ð�SL;��� �u�ӏ侂u���'�w��p���������fhJs9K ��̧ͤМˡ�.���C:+=�����C�������fL�����W�ߵ��A�Dw��{������7=To= �Jh/A����I�n3�%�2 ��J i�,�<Ø���7��V��8p�鶁c���z#!m���B��ՒP�c;�Ͽ���:)�蝙����f3O׍��S�ũ�������[hOe�<�v��_Z��3
�%��l���;gl����aǼ��a��f��#)�2k,����_��鬙�]�w�B���>����?�K�3���V��O H�qB�;�qL"Xrx\��pN�]�b�����E5�撦�B^�'Q���r�hB�����<	���{\<.�'�VJq~�<�����Q"�G'|<{�s���Tӡ����f�Bܤ䃪Es������)B!�~���ƚ���T&�P�xl����4B)ڿ�lf��(y4��Bi����+���J���y�X� ���E�v��k�ݗO�*x�f'�c?�6��rP"x����K*��9�0om&\�3\X��Ɯ%�� \��f���9]�������b��۸d�C��}nY�4�8蘨L���_�J��%�SZ���J=�*~�/�J�֜_x��!5O:��Y_t�_ ��f��A��@C�տ����-�}�_��7Y3p�D8q�7��-R��_U�~���R�L�`]�2����O�~3���8hkvE";���!���vg��r�^K�����R����ϬHM�I�ꪇgk]D�l��MA4Z��ᙒ���u�eB�+��7F	���g
Z+���J�E@u00u���ͼ������!��l� �����e���ӥ2���CU]zx�|B��@�_A�n>��QQ�]n�:��������՘)��6`�Dy��^p_� �NQ��b���?�A�8=T��\�#:�C�K$�8���>OY���w��.�j"T��+������y�یc`��
��T����H?09��~-
;�O"n�[�Su�z�Ym��9��ŮI�o�q����B�[j�J.�����B����l�Jk�?�$�_�K��<r
�Ծn'f��Q��ە���%<Y�K2jP+JCol�#�
��]���V��[(3KT:���ex���������I����ea�>���9��0����^ChZ���<�1H2"x������*
ڦ%��N�zR�p`���_�%���@���˔�7��!>��i���S��Z�m����
xsEGD��I��J�Q��|M�/��`�Y�%�{k�/+��"��	p#>����B���ē�������fb����>,��VyA�J���gպ��֚٬P}�7j�]�6� �԰��D��M�[/�����١AM� Ct3� ���o��V,\u��g@׼Qc�ݺ���Q袘��ߕ3y�	>���｝��ȝZ�X�:f�]v[!�J�5�쫦����R<6����)��｣t�+����V��%���l�zs�=��	�s��x��qR�!i�V��[�d�$�����]-��N��zG���2��J��C.V��I~E(�d�T�h�ɿ���%��"��V� QWDv�Jj��0��Lx���ԡ3���ߌ�<9�F`���'߀[{k�!/@�$?��s���b?�'���>	�7���&����*�,*���dC���N�QOj�~kW��L��?r����ðp���?�p���b3lR#�Ʈf](�#˫�����Nܭ-J;���=������$0I��|y�ޓ�J0RK����~�9�*�*�KqCI�Q7y����|��]bϰ/�T�n����Ѷ�]�6��0�XG%f��S��)X�ax�E.^;���tC��d� ���HF-�4H"j_qڙs{2��`��c�4�ESG��Vܰ�45�����@�$���	����vf�2���d̆�?#�	`�J�<�jI����k�j=�oa��4E<+ſ�d����F@R|���ܱ�S�>�܉>!m����ʩv?➳d˥�[��>�z��1�ڣ�ѯ�QЄ$��8k��?@��-��s�Ĵl7l��΃��0.��΍��՜�� ��nc�`�p��զ�]��������={�<ܞ�>\,�y�奴���,�z�qq�\��օuŘ|�JL˼g�������̨���7#��&�)�A%ؔ��,�.T�!#��"H�o�g����[��^�IU�����ҭE���E�[&�߆�"#�%+���Mz��⢄wg���`懝�-_!<�s�]7�r
_%n`p]6h����H��3f��␧e+��V����/1��vZ&˂����v�.�α�r���;s��������Ŀ�����tX#�|�II}6�K�Z'� ��o����BfX!wƅ�'�ج�P�%�b�N�ՇD�i�d����q&6�p�Zڱ�ɤ�K�R3U���@B��-�V�G���>�Hfg��t5�&sMr�cjҊ
��to��G�jw��Rg�9o�+�6���	$Ia��ɽ�R���7��1��j�<�ۚ��ԀZX�$gj'��*���
�U��)j�[�N8ެ7eYPa��Fݔ���*�:��l�Q�Ιm����WDeTe2�R�>58�Gŷ
9��.JQEI�aI��
�E��b%ƶQ����~�}��{�Ҹj�}DbJ���T�;�^����_�Ir(}��k����k&�O)%�xD�MG�j���e��C���t���S�/</���2���m���Gt��]���4-�	� "��s����C�i�z�>�f�=�U��>ĴS�ٮ��/~�@�FAWQ��OX���bߚ>�`4��z����!���	"9:�7d���1f��lI&A����N�/�Փ���2��hH9P!�&�Ý�������vOv�KEta\@����^�-,�1.�ې���x-��5����K��������Ґ���=ԍ����.��l��jQ�h	���*YĨ�4��D��pK���e;��.0Z@�p���] 0�uݼ�V�2g40�U���Å��s�L*�AB8"�5a�v0#���g8@�UY���A�a(��M���2�٪w��<0�2�`�*����0��<P��6��`�	��0����d4�t���#�◒�����+�G�d�*� �8M�H���ٙ�jMz �mB��L������y��KA�òD�^���(�Z"�����A�Cd9������Ik,�wuC1�K�f��Q�-G�T�]]���&���aH���?���K'�en�ۯ�I����9�Y��<-Uԟ"��2��rc��hpL�p./�~��)���}�
�E�y}ۢ������q��$���Q*w�%��������c^�l��dU@�q|C�󜿧���7�칮��.��Ҏh�VVI�A��i"�;��4�t�+��	qU�z:�Y�ycG���F?I�i~4c�;ޭ�[FĆ�K��׳�@���A �w#�OpA�⢁�۠����s!����-�(�@oOǻ@gp|���sʛ]��3C:-h��z�0����d� L��ydQ� T��u(�������Z2EN
�G���ca9��W��]��vS�N�JKO"5�������k��Pe�.]���M��#+���eU��	X�K�.�L�X<:}
�`kܑ4�\�m�9ңrYir�]"��r��Ԙ<:����}�]>���
�9ƖRB�8%��"L��b.���Ă���՜�wXU�o[�df���wG%�Tx�yK�9�'B��Ɲao�Qz%m�r��\HRP�G�zt�ɵ�����8 �k�rٗ�����Ga�2s��b�4L=i��3w�S�m��W���F,:Bc�93Qt����i�nW�&'}��e��6�l6��
�ć�>��r��Z��
�������>��g�,;ϣs|�6���ֈr��8X��Q�9�|���+j6��Q��hpܭ+H*�я��˘e���C���3v�qw*=3�]g�Y2�8��7��gEam�ǥ�L�1 c��N6R���A�	���3lL�)�[Y��u���W�K��=eB$[�86*�
ت32�2*�n	-	���p�Xs֤�t�ܷg�ٖH��c�@&k����I%�����{�uʹ�cŒ0	
AyH@f�몿�l
̋����p����cq#]�a>�)__$*ћ�Tu�P4������A�4S�2�(� ��*=��r+Bg��,�W��	q^Ѝ�}�s	5�ظ����O�)#N]B���Ee��0�ʥ*%��A͟���K,�`�Q_�3#�x�qTILe'��H��FM?��8LG	��O�1؅^s]��tR~R��|Y���ƶ��H�5'�MY����7�"���;Z� e%��Zt�8�r�׋�E֯�O�l�Q��T��t�:d���3��f�^���?�J^z^��E���f��TX�<��@B�b��:�O֑��\2�<o��z���4�X2$-���Qy$)�T߄I^0��|��|���m_q^�7k�N�Ұ�KK�O.�n����9�xK��˦���]�Ǎ�Њ6=<�}\� �X��ĺ'�B��*1Pf�5?$�����w�ס��*a�c�6fOAGX������	��m����[��F�ε9
����qm/f�N�m]����5�Tx1p�m?�C�PVD��o�+0�(S,|���S��>�$D;.T�:��x
EDD�{�g��s�w'n1@Ԑ���8e.�|vQ�����e�����/�Z�n����3��槚�XQ�M���]<�U�P�������!Э�s�a(��1h���a�Vebk*P�b_ 4�jbm�`�Ū�n�A�c�0"sT�~��(�vQ���j� ������@ =~j�0:`��!���j��{R��.��(�b����~O8���;�Ԭ]�D�sFdUj}_`��&ml�0�c��$�@��
J�Ɏ�pH�Ϻ���� ��6����b�UEE�8�$�T��mz�9�Dnv���^:����A��k��w�ֿ�s(#4�)x!��X���m �m�v867���8Ե3�,�d���*2q��N�`�;El�IX�Mv����E�=OC��kp�0���
.� �=��gstV#,�g?����.��KՈ+�M��s$�4F��S��]�>��)Ti�A�ڪ��Cb�>���`�}��f�7�[�O��u?y����G�٫c�[1UH&-g�%C�����6�6W�'T�u ���̮]'H���:�
��Nu�m[��}(<�a��76M5�\L2��s�)ˡ|n[K���'��b��(vѠ����&X`�;����O�(EWQO�Kpe�s�|,�/3�X�	\���=iU�5y���&Nϸ��s���7��D������{�F�Ĭ��׫� $.�l@�F�	
^�U|K"�j��;�V6K�M��P�Mj���>X���DU�R��~iC=ژ�&hNXaX)A���&0����AJus��ҔQ�1���|/d��n�r�W\��
u�5[�l%0�Ж���f�{�z~�v3�C>;E�:ҫlD�C;jOQ�߈ �L߹��X��	�T� �{�\N@u:�?�����(_m8�B���$��Ĺ�����x�`y2~�)l�(��@�w�`�6�5����c�6CVX�bO�%V8fT���N�>���Rb��N�ci�)F;��Ј���A� �����ġ#��9�����}�4P%�x6a�WQK�~�q���:՞�L��x?/S�|���2��|5a����Ȫ0����0�o � ��邘��]H;�s
�����b�&n���s?��ں��Ck�7YկD@ΖdY�8S�<��g������5�_������K�)�ЂX-d�!�Xb�2r�6S�p�k_�idP�y��.�h3Xui�7�t�T(Kq�6��0���F@��'����41����R�@��Q�{d��!����=�1Θ����		���v�k��vh��`?��6e����y9x���3��n1c��T&�zMb��������%x���6e�s���?�;��K�1>����� u��9��B,Y �hJ������(q&Nt۰��Y� A��r�g88�VuC*���xd7���@vP+�� -�~<���Z&�Ѝ�'���q�� ����P��]n�ڟ��Ӥ*�cN��MHM�澆���r�o*�/�
�ä	���!�,���Y���4���ǳ�ӋV�2�s�u�r�rs�s�p_������(��;�߸=�?�f�?�Dc���J�@43cX#���-�g�ϼ�����Y�Q��4������x�	�;w
 ���z3t�f�B�s��ٚ�����@@��e2�R5J��Y�����	u�� w������8�0�/'*����f��'L�&H:x6��̝[�1F��X�g=/f\��
w��N��*Ⱥ>� �(ZբT��S<a?��"�;?����1��ȁ��nVM'��X?������ފш�W9�*�T;�i�]�Q�0�̺\�Q��ik�,�`~(�Cv�{�Cqe��'v>'��KΣԼ|�(��J�[>r�	p
���x�c��՞FUU��g�m����G����y�L�ξ����}�� &�M�#����L�v�y<�nF5L�߾� �b���?�L�S�fK�ʳ*�g��`ͳ�{�ç����|ӝ�D3�rR�X�rlopMPn��w6s��s���@�:4����4��x����n�~�l���X����#�ђ��ZGMس=��Z�Ӑ�N{���n�gסJI0e��{62�=��d�Xڇ��l-3fV��5%g�1�T=�x:�cR:g�)�����v�7����F���7e������+��{����y[,��
�K_�.����T�)�~�>i�k���Ē����o��(��'��M�3�|�[Qp#.��#�|ZP\�Q/dԥ�S4�E����
<�b
8�Æ�4z�8q����<FcmD��qo�9��$طS�ɻ�9� �Y�H	�l�L�|0˨�T:�ߘ�Nӯ�_&�`sMɇqs}1b(��W��I>&�Y�~}{S��}�@TϟuL�S�d���i�#�.�����l�Ҧ����{2/,4B��h��_�\��^��ֳ�Ø��̹Y�Z^�C+"�b��ۯ��^	�Ľ5�7�p|q�ؐF"�C~�%�b�u�(%=��#���Ü��jЀ*a7���l��H-��p����Fࡷ8���u������2ׄ,����w���\��ނ�]���'7a��Z`�qg�v:3��O�ro��Xk��s=��@����
Mi���Q�r�K�Q���n#~�Ǝ�9��e6}��E����<D�YF.O�;@�GIX���09�`�߽�Qä��L�o��t�v�v�:ρ�"!� �u���qe7�:�Dj�jDt����i���1��۷t�h"�m/W�ndt�B��~��b۽����~�1Tj�H��mU��p8�,�0}V��'���?��ʗ�]��wT��_�ɻ��M^3 �}��u���ft��&�p\���Ыq�.��U#z��2�.��A)c�}^�����5#c�r�$�#�[��� �/�������	6ty��T��6�����9��.�����뿸	6m�P���tI��_h)��>��IA�|�#�X�\:S�����g�9�C��-���)���O8���9W�3	��z����zb�S��<0oU�1'
���q  r������H{{�ޯaS�I=
��(����[�~1=�����e�Xc���.	��M�`��d����K\�Bc�8qng>�z�*"n�}���m�y�t����O~���D����}f{W "���*<����
5����a(�ZX�W�=ry�< �饻���fp�:Y�w���݄���\�+	�q���1��-t�?lu~ �Dƭ���s.A�1
ߞ ��Fy��D���C�4'����M%�7|�*����,�`��[�݄�6C�X=���Lm�ʐ2;�!�tf�sb��8�m���r�v�Ia��r>Ķ0�~�8tL
�3�/���z�sQ�ئc�D/�!��ٚ3ө�,*��y��^G
�.��?6�"� 3��AP*���]������"Rn��,���t	ě�-e���eA?@��l"�9П4��R�m��i��������%N(��))*�2e�m�S1;��ɽ��z,����
�տ0�
�K��i�j($v������*�~+2�Y�]2֖{�\�^+ba��gwV~I*�P`��϶@a��\�qB��R�e�� W�T@���WF���_i���g�N��T� ���.HW�]zQ�#8x�A���{+�P�����|>�7�`D| �Ҽ��L��λ�]	��j�J*��,�Ra�ɺ�(�.�S[�y(ط���!!���,��Q�������n�������:h�P���E��2��d݅!���k,�����5��<6�a>�=��1Y?C��c��,���lw���|B�l�ȆW��!C�n�
v=߭hi�/��[��k��`9A� X7�I#�Y@���{� 6A����y�>;y�k�.<�E�X�`���5 V�
��G
��]�+����۵���T㊛�p�/�C���C��T8���	A��nm�@r��u�8�N�x�E�b�.\��G�?%j(|I�މS�k�����-�\C�N�����$C���Z�cd,;�m�(pƥ�\���E��u_3���AιEx��s�(F$�[�԰�l��݌�5��0wV��_A��q	R�ѧa=!��)�T�3.���'{9lJs��C�v�d�^!ˌEaaE��it���r��Ϙ�\Ya�w����S3��"CjP�jX������D���ոKΟ���K�lu f�.��ʅ�/����ũ�^/>/I�@�J�V��J]��	���5�t��}��;����r�7�����C�	�M��zٺ	�nW(]�+�(7�j!���h�D9�"����;�J��rp�3�[
�WL	�2�E/֡#[E�����$=vH��=���
c��C�^���&�
�|��K|���7/�6�s�:u=cf�'�nɝxi��!r�&Rx
��'*Q3�����n�S�@��Q�H��i�Q	}=�7ZS6���f7p����PN����kQ�̰���c��ZH�)a���� �6qȿ�;*%1�~?b'{p
�=C&lF���q�-��ƨ�c˹cqJt�}_2�(�O�Z�}�!�!��R����Y��6����_�=�x �3ƫ�w;]�W�W�dr�D�-ܮ���~}��	��x`�c,�zc�D�6�Q���z]4�eh8�����90��Y�h�����]�Y���
�!,Ϩ����_�(���X�K0×Rx��L���k����`��}�2������u��Oѥh�C� ֦+�J�l��C���ͽ���.�1ǋ�|j�)��ue}pP�G.���
����Px�Ri��M@�I�3Ey���P��%J81��_�P�����+'���I�g��$ _H�k�|���t�8��v��Ӽk,Ӟ�e�C������}���(��*�e��SŤ��XɝL��]����!���v �<BbE���DTDh�뾽o!�jvQ���J��k�B���`�"s/T���襙�Hk�k�(y\�������j/?�nG�y�?*5��Q��vk�����Ֆ��s3��ԋh�y���QƾM���m}$�e�K6�	\�w+��)S$�	"^FBע�$ɏ,d~�m�b�q�Ai�0�L�C�z8�ِ�ʟ$ ��֩��>��LY�߁�����g������'7�7�Ҷ�����(�"�����	���[�m�}��p��N��M��`n4� /	��A��+ܣ�~�2��q@Γ�D���}&�H꿭	���:T{��:��q+J���-IK{(�@�]�!N�@z�]�6���Y�m�

ft�n�r�";+������B�=|n|/��/�s~P��]����i����^�a�y��x�ODj���D.y���i��Sܻ�7&��=�Ea��&�ЖR��؟��j�*�]�^�;ĻC�L��a8>3�O�m�k?+>�eKe�	J�|c����[\ZG��#���,��J��G��0�֮�Q���ԉ帅^N"#�]͗�����Z���1���ږ�OM��i@�|��R�ֹƫ�Ki�H�)�3�翔��)>9�WC��K"؆�CR��\Vn��N��H�F���eM�/�c��ۮ�z]V���xO-�`k8����2������ռ���]H���Ċ4�?��Qщ�RI$���G�� �<V�c�)]'�(_"���M��=Fy��P��io��T��\�>�t����{�;�?M̨����@]����B�����p��lT�pZ��w�/G�)�g%��N����d��e�W~�m�I�	�p�)o���}���Q8��r��U;\ӇqӦN=�N��<臄��d��=���_���cj��$��ԿcQ��?:.�N��ċ��<�)��Ə��j_������o"B�s��F�#�;�Sݪ�6?�Q�D�/oX*wt����V����� f��ϳ���-=�jRk��ؼ�n�����?m�U(7��߬�6Bl}��{Y|�tf鲂΋� O�;������!�0��1St������"�1������I9�vESk��ecezR`��){��Ed�����W4�^(�W�%�W.�}_��a`��9�t���m�����D�qm�XC��8u�p��Ua�
0-�U�kb�N��s�O� H�+=�����7zD)������]$��|����b3x�14{Ms��r-�ZZݢ)j�y�r��6p�x+g�bL�G�c(S�n�i�X�o4i̠�p�� ��AA�S��9���]�t�a$������a��_Y CVnK$��v�Z������{��)ͯ�B{��A�dr;��u ���
!nn��S^�K���]�n�"��T ʦ[��>�,�3�Fzm?Ⱥ�s�Pbt�v ��Ȥ���+��Z>>�GQ�;����k3�I�҃}��-'�����%�����X��t��Zď����E����x»�ok��@q����NV���a/�~�m>��Q�B?Sׅ䔹����ב��2q8YΝ�s9�l]���w�ܤ�n)׹t=t�.�n�!�rb���J*e͛�ML���H�$ez�i��-�Us�.��vȄ]0�v�pp�H����M�>� ~�%�;�Xk���Cf4+�4�}��t��KmI% �c�h�S�GH�uRn��	TW���_������r�e"��e���ae�����޴.*�5�6�1d�ސ��O�q]�#�*�S`.������K��4��@d�Ȯ3Zb[�� ?������i�͒�������9`�*�#����҂}ŶfI���l�?⒙7�])׉$U�Ix����$�X2�3����v������sn�n��ؤ`z�g;��d���maG��ךh@ņ[E3�{eg�29��jK{�HĴ����	��i-g2����ң�E��oFR���NP�S�R�5�9�:Vm\��"�O%	#�����Z3xA������K���"{�F���5�o_#�8eKW���� ��T"��ܑ��F�I��b��9�Sm3'��0�����/��A���˯^���5d�
Ҷ$��#<�Z�����S:�'���"��朩�5��&;5����@0�܄;f0/p��Ӗ>�Z1ft+�8ڣ��ya�R6T��u���	�ȯ���R�43Qd����&_�g�س�&���>�lJu&���H|�P.��+$f�����F6MB���� YZ��ս{ڭq������8B-[��yF������Χ��� :��rk^�L$��5�%r�1�8������gxI͒��ʚp��(`yӫ��$����$�V!f�
t�=�l[�+Y/��
�����7 �����P�X�JR�v��ۊ\T�?�Pť,_}����a�O��,�b�֔�Qz����D�O08���Q*��j|A�v�������i�ȿ������$�G�d|�Q��zTp"ؔ[�ȻO\�?&�ѐ`�E�TV���.�[ڸ��	m�̮�
�����0Jɪd�ߠ�p'sq��elў"Ym��P��":e���R}�mʊ��a�q}Ȼw�Snn������Y恅~�a�]�}c�g;D���}��r�X�m�7)IY�e�/?D�<���+:�-�`�������ʅ� ������AS+���/O��
�H72�0I�nǪY;�k�u{���o�cN��olnVQ(W'Y�
V<�lYR �.%��qpl��zA���ȁ�`�0��b@�(��Yh�<�PBl'	�%��s�q�͊B���
5���M�[\����0eT�\�e�v��iA9l98��#j7c��,!�^�����j$�Ă?_,�R� C#{3���/sG D�h�D�Fk���O��cP�/�ls�oث�ZL&<̜�#
M�T��nֲ�
�zTԙ �'œ�?,�����q�j�8M�����3q�7DMv��&��-�x�@��jҩ��9�$*�Wfn�%
Qg,Fӵǐ�r�J�nTΟ;���3��ꔋ��G~ʗ� ��A�5��!��}�>#˸|�^Ĥ���sY�J��b�+(�F��Kd�R�S����b~�F��ة��몤2��[&Fu=� ��h��DB`Tp���O�#��y�(�;�L���_����h�n�kG��Lr��+4������v�m0�����N��}s��c�S	�{0b�l�$��=�u;�wb|���x�3���V�KM#z��J%%���Z�Aj!���ܦ<��K�-a�>� c���( l41~.]�L-[|��t/I����R"4Ri=-®�vs�sötύ����$��)=�ڹ���=ʎB�P^[��0V4��KL/�������Ӗ���ø,o)uw�
���.�͕�%�GƲ�}�lW:���ۆ�'��ǭ�l����A� ����A�8*�{��l�O�_����2%�dָѢ�K]�B���\�����f�L �kv
�Gj�m�`��NǸ����i����&�:i	�[)��� �qG��C�	a���ޓvx�8\��(�1��I��[@��Xؽ�z�g�=B2��w�9��,�z��Z�8]G%��J�E��W�o�1@*�����՗�9�ɫ0���`�@��x�^�O\��Ƕ�:�!��Ժ\⃫ܛ M��d�ϲ��ٻ�n䮗0R�T�DXM���X�D��Ǽw�D�*g� ?pL�02�9�!%���rk�ICu�)�C����[�2�UGcjBֶ�<K6i��#X���֕�>���4��ϸs���D��x����?����0d�!yy/ #�}�"Y�$"�j:s�t\Z�����M�0��G�$�/�������ٮ����$�L����`� �2�]j�*�קx?���a�/�,�Ƽ�������D�kWo"�+���c���Y���+��z�>�l�p��Ԣc��|n��m0�;>e���.��-�R@�_K�5]���]/^eu�ӓ�j�}�z#����T�ϸ�9������j�j�v.�	]\�^��H0� >j lGy��oo�L��`��7ϫ����/N��l�r~��X
=��BΌ�
wM!�:�ٱ|P٤.��@'��������w��#1Q��A��~�n6Tm1�d�5�.����ŢѪ�d�B{��ظ#p��ύ��5�	O���N����w|��gسDX�R�u��t��#�d>��W�2���z��jD���f#g�C��L��m�O�1#C*�~ۯ�0X�[T+[�:��gb��-z"`�]�p{���=���=A�י���B��"��"�mj��j���] ZP�嬊s�8����ő��38Yn��HvAU���M�L��\=`\�|�����2�ǿҋ��tF󯆴Y�I{Tt<�z��<��%\�{i�WJW�<��i�_�F���
�?�<�`{C�,?T�E�h��<�r�l�dMC��,%�]X���K���t��O�ːĩ��ǲ$d;����3��+O<��|݄GCS7�!zd�s=9�'@������hs�d䦝K=͠)=�6�2�FzC�����x\��$k����p4�r��g���_�K��H
������~)D��F�{+�V�\�HH��(����%�����Q~C��a�m��V�0����^��6
.,v��D��k�*�j�@�uN0��9fg�J.�r�&%��} �]��~r��e�ȅc�~�hߟ�X��LLA<RR'~�Ɵ i>��H� ������^=�0�?Zh�L��)���Ӡg�������J��^��1�Z�ں�
W�7D����7ZIՄ`.85'EW�"���N'���p��.;��LYF��SC=�����s9�r༞H(캮����4_�	X��}$��U�jPGe���*��/��N3���UҖ�n�gQ�&��)C�d���¼����k�	A;�W�x�.�=��X���U
���n���7�?��j!�$���)_^���M-����1�M�q`O�	�K�{yn�����W��o��t{�`��X�m��Ȃ͈a��Ms����9_�J��������Ïo��㉪�����mV.���ׇ��,�Y�7�J���AkU(��+R�&��<��?p�5���C�k��.3$Ή��o��W�iK��z�cX`����.��ŬW��b���W�,�w�zq#���7�ڑ��,]G����@�QX`l��-�/���υ�hj��;�.n���@K>�?O������4�U�xZ��t:�`����i���P���-S���HF�DaX	+1W�r`�O��`8����g�����q��Cv��ON �-s	:����Wm���j�ȵ�,qo����N���0�'�X>[g�۝E���5z�`�h��%(T�������ˍѷ�Uz�'�.ޡf~�a��^�t��-���C'&F^��`+�?����J/�~	��1���Λa�6��e"Ҍ���9�0NE�F��~���3�%��EF�mӇ��;Ǉ��$}PVh]��ŵ��i8��g�W5��n�1�v�A�j|sJ�;��I
����5�s�b`jv�^7�"#�=c��,1�J�j�T(x�i=w-�'ׅ��Z�����J��@tVu����I��9!>%o�av���<������ �[ �_A�������D�B(��B�,M����P��k�R�k��<�ܤe��P<	�K� � I[]H��J��P�ѥ́~n`�f��i�L�t~5�"MU����ry���O8F%��� �Z* �J
�/�y�,sZ�����5B�W��T���;F"��Ƀ�B���������A���x,�%1e-�Y�,Ei0)�o�3E���Y���-�mj|fE�ʂHD�D f]?m�ʲw�6?\�w�=⶯�+@JyQ�B�)�bnM�o�(�X��%��8�Q<��?@���~�0���<��;�iO�Ix.`Ɗ#o�Ӣ��dv��<y���+0�|�ʅ���h@vê����-6�q�B�
���X���#6ä���u��Ȫ%N��8Amb�ru+��T����U=�%���W�Q'����q;%� ��m�ڍ9����%��Nh��vF��H�#�"ˤ:/�gQv_W�HE��߬kE�+x�G��Y\�/��Vq�9�y2Yx�����Qݞǅ2�}ƃC�X�����9)���۵!4��KpᆡriV�v�SH���o	3�������n'鏘s��Cq�2�\7��ȋD}�����&U]7��1�-�,��A�(4��`	N{���3ȗ�̩� ��Qcb���˚���;M�?����}/*���GflҪ�=�ٜ&H�\���5�ٖu��`��e�:-�AQa��t\/�*���H=�-�j)��םZCB��/O��6-���֍q��ә��:M����3�����n�����7��M��Qu!ڌ�C^LPZ�#?Z��������/�(5�1~��,�-n7Z��i�s���*�����p���gH,�}~�HAd������L�F�T������"�l/�;jӿa�Z��^�y��.�`F!TkN��hs�RƼ��w��eT�r6�R=��Ej��v�M�цg),�E�����b���T���B���ɋz���,=GQ��?#�uy��P��oq���`TD�W^�%$]��V������]�D/i3I��о�OƦ'[�f�F���M7�L(=qt$�e�.��O�AQE���HB�~������A�@�;�,h.b�>ML���ڪ��2ay��%剪0-�����B�ژ�*��1�����0%��V�qtt�����
d���0��FzY��n�Ӛ�^�k�V8��}��J9���m�l����ĜB|<�Lht`�����|��ȼ����b���t"%�%n�����b
�$�"@*�ӻ�����aI[�R�t���L���g5�`x��"B�n�E0B��'�-s�mX����Y�9��80�I��_��&"�gV�9�)�Q����檼�&����KU��J$���V������-/�"T�s�V\S��΍��ei&��`W^�K| ��d� ��-m�Ea�(��_t΢��X� �
23�<�g�*SҰg/Zv	���1M�i�d���e}�
�u7I�ys��:j��/���y�R�(�wO�gn�F����VS��i�*Ѳ�ݖ*6Ӫh�������eVl��]9c/K��M�vK�L�����
�_�g�{�U���""��3��+��V���	�VK1b~$�~����N�[J��,��"�[�;���B�_��b}Bw�mCm"~�*�i�wG>��m{ln��WD�E�����{l�&��<D�7���,t�Iӕ�Q�)�}[�$����?�_�޿�k��{����E��a�V0hU^?GHv4o��F�J��*�����N�C���e)q5�ن��S���&d粴O�� �WeX���(o(a�s�Ѩn�a	����ghy�o�!v���Rfn1vz1���^+"M���m`�C'��j�0˶Q\�5����<t�`.�;s�Ͻ>�J���SNX�H�8��c������0`��������|�3�R��|2H���k8�U��^��p���� v����3��?
���%�*�$��--$j8�鏐��فQܰ$4?%����,�h1`��"��g�mɸ�i ����$����������o$Z��yИy`�38��HB�� ���c��N\�D���2M�՜���Ye�5�S�ZPp�B���u+�ԍ����4V,��$p=#M�/�%ujz��jr�����*���
-�$�^����S9�d�Q�~�� ��e���2t�=E�	��W�C�Ҧt����������~�?��P��O!���c{�U1�J�rQ�ݝ����&��I��4G�*�.a�u���ӚC���]{�M����q��,<�����t��b�wu����m>��c���AG�/?�C���gC�����笇��@���G4rS%�j�q������~	���t����-�<{m(���Ji^�����H�Jv�����Sޖ�>��E&��U$��na\��2[�j��� Y�5VߑY)@��.^A��z�/Χ��4�R��w��y"D��I��Zo��yܷD���kȭ�MNx��V�0M��q{Hh���?]�E�K��:s��!^�r~�XeK�dB<N
[���-C1��m���ӎy������������NB����BsmO��Us��\B/�n1%d����t�m��|H��æ�������` [�ф��Hrm�hN-ā(�Q�{��ZkW0��|1����Md����'|߃�d5���~0�a�͔�W�)r�ߜ�<+nm�+�#�"���ӣ�ON����hW$+��_�����b3���}� ld�>�� X�,��IU����GX��{ɺ �/P���_X�Y!�p
��"�5sg�LP}yd��W��:�[��	��>�<��Ao��n�'l�5K�C��<b.N��"�[�U�e�x+���0�㚉�ͻ����@����]�&��;��^��ms8��s!�|)[y�����5G1yW�4�4Q�`���64:���`�&�,�p�m�����u�t>�g���	�#n4��$�W}$n�Q�ezr�x}e�����;��XИ�}�z�7����%l���4/�:���� �C<_|N��1�M��b/���;�wp!�I��t�deoSѝh �e�tm-��4Z�a�1�6�t��>������r\AÞ�:�Ab�`@�)W��0:.C?�E�H|1�����ߗ�q��U���u������9�v
s�Aм�?z>j�B�s �6M��V��8d���V��k���T]8��ׁ#YEN�)k�ő4q�X�(O�!+����zq����F]��𺷮��Q��xi��3����lا;����n��!x��8���Ph$"�C��R1�׵ 1#H�l��3�+9����m�w\}��Y̶:�����*��]ToF��u���O�� �X� $���ƀ&-�@Rf��9y��G.�L���Ki�bUQb���׃����IT#��O��T�Ri�@��<�|����7d�٘����]¬���Q�h�
-�1
��'M �������p�R剦<<�Em�M��G��]��
/���YXV��9���-�Ҽ{袌��j��(W��-&j���BO�b���n�C��YH���C��֠��3n�12�W�P����z�>�7�K^�"���W��G\��$�"�h��f����?@��R-]�T ����
"뗈ъі52��gT�'���r�K�#m5�3�G�U5�Tx�_�';��B'����$0�̄��:dj���o��%�	��2���t�K�P�!0'	2i�s�Gfό�~��uṋ������ Ӌ1�<��QR*��[�x�l�d��"�p�IdV]���'k�.�����a�d����;����(h�KoC`w�7�]�\����/g�Y�)P	KJ��e��*��nBiN�~L�h9��f.�B�z�� P���P����U/@���eb��&����Llr�Vm�P�"m����6�hz�f�]�Y����W�QK��P�Jt�w]��4��P�v^VtY�aȔ��N&�� ��mJU�Cz�KWYj����H��Z+��I
	�L��r������j���_ η�w�������w55�"$:ac�Ɇ8��Ʃ2�gys����st~�*D`3�{	T����n�_�f���8�yR�O��`Z���҈)w'��AI)S�����n�7}�M���c𤭹��嵔��c�7F�=v 'c��ŻfFf���[�`=�Zm/7ň簯e�w��d�H|���y��ɴ�4�$ȉRb���B��c:T�g�'����Ao��ǢjY���{������~I^'������t|tT�Dne����qkضd\�IB�	V򢲴d�#p�/6���v=F^9���$-�����x���Xݱ�5+&�;��m]�-���ՓG'7�m
	��Qq�dƤ�_8/M�N�<7��ꐎ#�73!�v�%Т�B��B�Vb�;��bh�$ �xCw����� 6�A��v�ΙY�EWzu�q1͇���@Y���Ѯ�&A����l���а��q����V�*ouB%H����gNպޓx�dԸz�Ո�2�Н%�bA4��b���Ri)q�񊓪�����K_�8�j�߽!���֒�'�~����������F"�̿�L^�"���{�� |��k�^�:q:)u���K(C!j�Fr��tWa*��o�E��D#��������`�MI�B>f�x�F���b�R�Y̔��������.G԰I/�*�RH�}�����'����1�;�G?ֹ'o�����E>`�*��5i	=���/�����^�@@���"T9�F�K>u��dߋ��>�B$�#��2�<1��rf��Lv�1�IZ0I����y�TĴ�{50wc��Gr��
Z�;�I�&�`��t���W�Le
��U�~ !Xܜ�`�_L7�<Eq;2���b~,wKB��j5��7�m��9��\BPpX͞<�g�z�L��������N����Q.:6���P�,��}k��)�,V#Z�Q�BnYB��'�\ ��w;f|��'���$��Z�춠����.�DI`~x.L-V	r͓l�Ҏ��ʍ������,wJ�X�Yd>�)N��9NK�7��g�?����_]�8/ړG�.S��1(, 09����R�0��b�4�5�N$Kc]�Hz�Cqnȶ��qJH�즮`��DE:�_�S>�}p�T .����*�)3F=򟴱�z#�9�8��M>��C��򁱃��0Q{��	�����EO�[7����5���Ub���RSŶc�bJ�1hb�HV����l��V)�y<�Z�`��t�16${1������ͦn[�po탳��z��97dh������ِʘ��s%��q���]�\<}��Z">���~e�*��)�%���6U�OM�d����"�D�v����@3%,)�7'��b�݆�F��,�]Of��LzB���d%�-�����fD�.i�����@��Y.D$�n�,rD4-�_�������!.�J���z�4�#S�?�C� ���B�j����?��i07<���`= �gt���{ѵo��l�Bz����6��l�p��U�m�]e�kt�ig� �beq�&�))����=��\5���⬜��z,bXb�M�),xb~=�0tm_"}@z?�;�.��9��z '��r۠j�"�gQ6�ԛ!$����I"M��G��=
�U?pX���"�)�K  ��|t9�����̛a��q��^7�)�h���0���;�Oз�/N�Ĉ�����D�k��C��^�H�M��5t�8�T�F&��� �*d��0���8�X���dFUGT�n�TM����g���^`���νXC�8ہ ��l���ֻ\|Y��S��5" sI���`ml��+��ߊ*ѰU��q���&�ǵ�S*�o��'	�A������~\}�4��&T��F��OcBV}�֏���M*%P�\r�P�@��K}��oS�|�������z�ƥ�;U�_Gs>?��@��+zmP�p�N����h/�!G�b���K���r���?7=X��f痧Q�Z�&�/o�y�雬ՅC��liJG2�t��j�?LUC� #�W�v�5eur��vWie\چh6>n��hnI>��h��oʍvEC%g����|�/3c�D��bJ�%�#�MJ+��htNLb�6���F���t�JA��(�����oC�)Z��z2s�����K��=$(a�?R`���l�[�&󯎃x{��j2���.�c36�_���?v_y���[Q�fAט��4����F����<*�W�#���ޝ=�l��M�p�7xv�	I�U��$��#YY#C�����nK�T�;��E3��9zy'?ʗ6�OUU��p�v����Q��ys�,��*�,޲����Ȉ��Qx�e�-���_<�]n�%>u�ŭ��	�#�(E��}q9�Ҍfߏ��_��?�_�C�C�W�^j�94A>)�������O�8��� �|�A,|3?"	ӌw��,S��C�@~��u�dt%8�ˌ�q�Y�1ٰ��p���{����k.;0��c��OtW���w�J��s`Bb��hH�}��
Fy| �R>���K�`�28�\�~�M��N9���	;z'��¨y`XbE�⾡�b6��v��vA�rZx�/�B0���Y�&��=�N,�p�{f�6Ėޑ$}���2���3�l7�ɝ �O3F��N7w�R�r/&o�,�$���@���0�%�fD��$�Y�?R��	��}�Ύ�[�a[?�X���9�@`X�g`��g����C�<%)Ձ�k��E�1��j�� Bp��W��L��r<���T@YS�>&�a+6h���Z˄�{q�\�ݜ�����MFo�Y���֬�]��-�G��PV������ots�x�aޞ�X����f��V�X���� �DY��r�M��x��F�T=U�tٕhY�zș�4Bb,PSMDa�#:Jj���@��mR���CQK���T�҅�*��(]�)-~���s�w�j9�x�޷(��&e�"�q�M�@�|�%�L(��M��Q�3=�O��ߛ3��^�7��<���T�h
�RuXlc�9\n����OX�ޥ*z�`/ZU���ҡ5(o�o6�� �KL���<�;b����k���k��"K�K���o�'����YFC�����8Ħ��p�����1pf��u��
b�N
z��	���-������l������0`oL5�tI��(�����O�ӔP���])���e��ʁ���4[�W݄����<?���E��@&���`^U�佋�<"�ZN��C�h.)���E����[t�bف��`M�N?��SM*�Jp�j��&w@燊�e�r�_���M6�Ͷ^�� �iz�H���a:P;Z1�e]�s�����v[m/*x[<�{�#
Vz	l���3"�X�vI�����o���<A#��}����-��
�yE!+/��3��^k5��y��t%��p��#���4+�<�FiH����
\�8[݃��T~�jf!�˹e�y�/tЍ���+���e���搬U�R �K�����s��8,p4�α�s�p*�$D*���l��@<5��w�7󘀯GH?Ѐ�l�J2IqNH��!L��S��3s�[��wK�/�/�2'과��?R���{��DB���N㥎�Lޅ�<c�y�r�E�]�>��I.~wJ�囆O�����jY��L�����d��2�n���ʕ6߃.��� �Ȁ������V�Z?�"$x)#�9�C(X=\�7ƣ�o!���w��������b���`��ml��2�9�8ͶFY.I��vn�y��b̴�\��(��N?���I�b��b��,�c�9�ޒP�G�f�Ƙ������c�Y{m�+�^��xχ� ��$�ބ�/ځ_se��J����3�E�<�}�R�t2˿L���
1�A8�Ґ��nW���JR�")��v8����B:�.n��C	���U�ܮp\�'��$fk8��?�2�P��NA>��"��Ǥ��D�Pp�����&�ֿT7�������(s���	��( lZ��T�]Cz�w�o���E9�Ã��W
Օn�1����DBC��}�u�`~{�qV�L�9�Φ���wp/��Z�1A�h�DU����9�6�@��!SpB/Ǘd?�r�,&OqS驙JK��>]l� \�y�i�3�g��"~:76ki��=1�?,�*�s+��T^��d�����g�:n�w��Z(�J��'q��XV��Q��YN�K��`�A�?\+�n������G��WaP����S���k���F.P�.0��z�`u��[��b�R,􁴖,b4�\���B1�SNGA�m�~J�E�4Y�����Q�y	�%�VnԂ�u�6���v��o�T��U�;�5��<W8
2�W=�2�lw<��z���{I��\��0�Vu���PlB�9�� e0H#>�� lqS��|��e>�N�w��v����{Lp������t� ���l��y&����/mm�o�F�P� ������ɝ���"�_^H��oT��|�c!��ܣ��i�U]
����kK�V��(�}��W�Ѓ/?�����c���WJY�RE��t3#��.��g��r<���.4��L<	�aΩDEp ~�;��-�����w{x�Xod�f��W����^V�?5(�x�����/�l�����/�]Će���O-����"=\��p�Q�|}���wS�iIi(v �5<<\��;+�s�_����@Z���H]��g�O�a4"%?@�����H���߹
-~����r�	����B�A��k���0l�yi���g�ҟ!9b���e���q�$��b��$9q@��D��RM6g�L��:����4�Z�7
��c��D)Jɳx`D�H�t�A8&�UF�ߚcw�	�T\h�;�!sV_����e0����a�ޱ�Z�	����YXG����Y.�ds!�gG�[D��+�Xf��9w�u������?:[��<�ˀ��鲉0{H������ȑ��w����)��!cFQ������X�G��⫥�y����A"z*}ڼ�b�Yrw��>	�h0��܃U+2@21&ڛ�΃��%()��v�&��n^C-m�j���P�6Gc�I Gb�l-iG�нIS�.-멻�sD����ً1oW<��Fs�_��u
��v'��J����ܞ� ��j�{����Z����W�pr��4>e:h��2�k͏=2��a� ���7lW�=�=X���k�FP�� ��g���!Xg�|��ʪ'̔(bO4�|�U[���gFE���T,�Oa�j���f�-�(�\Yr��0KX�Y �)��k��<�MWMӝ}�+�9ԡ���z6f��=���E&L�R��{i�Lv*�~�)����� ��B<�����yV���s�0�~�:|�\�`�T�HL�>��b�]�uؑl�K�nt;��u���j?�����G�8c]����wP����wj6f��ȶ��E+t��o�lIe�8�k��H>t���n7��<�+*�Ss�[<����WH_�M�`-$��j�)�*l�d*~���M1��@B;����M
��y8~��/�\���㝯]�J�-����z����I�}�h�
��3]��R3A���7)+�祝���M���]�޺�4�.�Ղ�-R�x�z҈|垡�>�I�ܻ)JS�����y����(���E|�$/ۏ������B��iDxQ_��p!o<fg�*��h��{��a_OS}���%���E9��	B��\J� �3����̘�
A�{��Y�V8u+|sNGW8�G���~8db����������N�� ��j��dx�Q�·��À��mA��s:��9}���~G���q��&|��X�R�Bz�2:��9@��E���V�y֯9�_�-�S��TIX������,zIB�-p�~��A��ó�2Q�������;�U�L��V~w��t�dI�#+�ib�C@����m��9UՑ	�DwZ���`Сf���d\��0��Jy�@�͂��-�^x����r�#n�?�'�k�M���Lܦ�e��豺�&9;7@�<8����Q��OaΦ����>�2$3����-�2�L�5�$ ���O��!�¼S�{A��\޷ş���[7� oG-�TO�c�fg�b�{���أ��fxF2/�U�d��.8\s%͜��hD�O������_�ܕ�U(C.X���M&*4	�0����C�9 ���1-i�4�\��+)ݕ)T��N�o�"+z�wSL�>\����xȃ����S��*��N� y#���b�rx7�<ejU p��	U�
�E.��m�:�GA��;q��yDb��Z�:�!s�'�x�E�X�	�ݽtlX=vW[��d|�'I�����A�N�<ǒ��R�Ъ��)��K.�\��lB��
o'��	�B�s��j3G. >�i;nc*�lFך�[TR�IN��ܛb�r-�����%���R~���`����x��y�A�d�[��7K�w˱Oq�Z	�;ʤͪ��jo�2�Vxl0��>S>�}iv����;n
��^���j2�4B�].�gۛ	�q	���R��3%�H`\D'�n�f��q:�������O����0�)s�0�L��sJ5����~�?W�>�N��ي�o�\JḴ /d~gP']c�R�h(�� ��W!��f+��<H�2����V�0�
� h��`g	q)���#Dl�7��.N��q��X�p0��q�Ƙ#G�C��BF�P�z5��K�f��t^]�ww��A��0��cCc7���~M
�`��	S�2�S��
D�D��7�6?�B������J���C�O˶`,�Y�h�+��#q�ĊaDYy%�h	�1P��Z�=���p�WT�������\s|�$����)���|d..������7�+'�����|�SP��6����}[���h�bW�IW����}r���D�+K�IN���ZV���U�/狞(@�>��~R�w��qBo[|{#����%����_���X�	"�|\K0!úH�*�,��E�$��65�/rWk������4OY1�ME��^�'�
�5mB�)��<ͪm�f������=���c��I`�i-�T啕�����c�(�[����� ��B�f�����;�D�('�IvA]�0+)2B^����ӫ�B���Cc3��r�#5ga�f�������-��X#�����s*��ϝo�0�p~0����P."dE�1\�ćZ��Y�����-�/�5<�avu�� K�-"���ʨ�-�
��]Hs����vD+�De#�$���1g����l&m��I#
�iM��� ~���'3�x���>I�t�M�B i���ß¦�b�o5�r{<1'X<��4Eq�+:vVu�m�>�D�q�,;g�!}�.ݾD�X����j$6��Q����MaR�Y:��(��F}�<������ ��1�(\��y��`+�z��]��]�R&�g����%���K�˪`�$�_PTe�>D��̠)��X�5Κ�����_��?�Ҁ����̯A�����).|R<�;IuT7���-N)�k�A>��Y�S��Z��2��X5�~�!���>������X��!�d�>vnS@��#�?���ޱ����G��/J�t�
qF#�m>5��y|"s]�o�����Y���?�-�p��̛e��,��R��fp�#ŶP�'�#�J�ٿ����DHC�Pw��e���u�(EM�b���ƣ6N� t29��A�`��w"��(�t_�"0��$,��K��2P���ve^@ ��Է����v�� V�o�%�ɫ��y�+*�� �>�ުW�����6[L�����w*��SQZE�m4�p��Ft�@!B�p�g�ȱ$�^�ȫ�}�,T,��P��P�Y�~ݹ+��t~��"12nAJ��lq�A�j7Y��wNN[x���3\o!�r;u��:c�R\�:��Iol����ɀ�:��)ܖ����%�����Na�9��_坚���(�����}鰚����W�t.@�����Q��
�n���!�J��2�z9(_ʓw�H榋�>�&�3��h̤��^��'�dN�IU���elc�v����� ��(�.�}�ZE��scy���6�c��&q����;8<V$(^Z"&�P�J(:��{Ч<k]�G� _�����H�A��V�uW��X適f���4���T�e�-��9#�t:RF�VTҔ��lh�BJ���Qop��Jb�-/��T�>��^Px��t�+�G.���yl ���آ����U�>0އ��C�k3�$X��%�2�m�B~UH��']8Ԗ���b���-lNo���N��T-�o��k).h�Wߛ�9�h5����'��o=k��d�]��� Aڌ#��܌~�Rn���L��t�OʃZtm�=tGU$8��+GQ�� ��y���`,_7i�l�6���c-nz�[:L��n)���E\d�ϱ���(&���Z��l�&3l�ٛ����rQ�JӺZ+�=�{@����T��d5Z[��w���tx��옳����*�?{�+ʜ���v�;ʼ���<&�� R�ߙL,e�BBFP]���^��@�C�{�@�MQ;��u��Ep>QduR�A�=|��Y��W��>M�'-9;��P�mN�g�Z(�����}#��|��m�l Hw�>�픋o4��G|]8��|��]f��~b��6d4��d��P�<<0G��i�ǘ+X���|y�SU%��N��g%��,���}1q��3А�R��i��1w��I�y�6�t���!u6��L��ʵa,�pJær������.��g'sC�?���ic��P G}{��n�Oe�oz��~��J��`<.0n�ę��!	��^��b�(�bh���z�9!�jJ����uq�F:g#\�-�#�d�Q�h�?��,UV�Чy\��u*�DP��7a�5$d�E�B� �9�V�}��m�-e�1cEf��JC�0��/ |�Z�ܯU?pcŧ����<�gy4=9#
��ߟmWk~j�^��'(b`p�,](Md�ؿ�2q��?(vD�y��h ���J���Y!n��
�O#^�o�!Z?paIK��h*���TW�ފ4�_ ��=x�ĝ�٠HHn�㣳��Epl����h��R�qt������B��j�dE+�d!{�Hژ��7?���aM
�#��P��.1?J�T��BRp7��o�k"�a�ڡ|G�#`?4(?}�M�9W��QZ���ڲR��L��\:(����j��١-CA��
|L��#�Eg��$ ���)����_��\/2����M@� �1w���
�T9���=�=ǣ�F���O���