XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����鴎�5�ENX�m<QZC�y̽��Wo_s�AO�H24Nf�6y�cX��g5BN���C�~u":>�2�Fζܿ�sͽ��@��kꕟ��>h�ƾ¯= �$�����Ė��O�G�Ս �ģ�U�\�YD:`�5��͊o��6	�\�O�Spe����ؕP�pE����n���Q,�?�~���7u�E���5�'��P?ˤ�`�^T#�S�#G%�n�RR��]�������O�:ڞy �P����ph	�fJ���xF#I<�תtm���9x��w�y��D��<T����;�TA:�࿉����5=�<��X:V4���j:����u��`��c�޽�5ܩj��L=ܶ���Zj��.t������j,:��p��~�
��b8����?a
a���7����q��Oc�B/��z�5>��E͎I���1��ʹ�;sB�Tÿ��W���r=�HV�Hr��U9^�|�V�a�M΍�T�\�,G��Ż5��(F��w4	=0�G	���A��W���<�'�mmA��yj��ُ=O�cC����^RWC�$k7�ts:���Ds1�����W� X���V,���3S�#���,_��Z���.�uL���0�i�`��?��]�Uq?���k�y#��#d��o.h�ӣ�;�&>%-�"��']#V��{)9ߛ�r{<��Z�)�ћyV��ˌ��5��ؽ���Y_�B��/b�^�'G��^e"Z;A���x��� <82�XlxVHYEB     400     210��x��6=-�Hկ-����i�Ab뺝�l�,�۠V��v�辷���ע��^�$PG���v���Lx,���9������77Mtȓ���s|T���X|bjJ�C�02f�W��
�YD���k����v��$ ��s�.�-�Z�8fa��ko�ЫC��^c����R ��ƌ�A\8FމL��ӡ���z�(��7�T���%���E�B�׍}�U=�||B7����gl�*�޿YrG#d5��K�K#�Vה�9*��=��B����[M��U�X���Kߏy��"����1=�QO�5�s�8n,��َ!h'�ڏ�����YM�3��_�vf�9�>&�����#}���u�	�WKǂ 8�"�
�����
 ]�`��$qG�G�Z�`�p32�� �*uct���!Դ2�_vRp�?��.���s���Xq��< Ww�x"gOw��I�0�;̱��2!Ĝ�t R�=��K\��(H�ŋ8ݶ
�}Rh8T�,{/m��Gj�FuXlxVHYEB     400     100tY^++�h'.�MQ��̚F�a]0�
ظ�>�n^�剩ҷ�BD��E��&��5Z��dD��À���kP�@`���wj��}��Ֆ 5� �.�B!�)�c8��@�Tǝ���~_�L�.�@u�(+E�a�F��P?_����Z�Yr .�l���^f�֫{�����aNlԬB=�G��jl�Qy2�`����9�ds}�S��^���s(V��
5��&�1��m��xlB,f�.�����o����,{��-�XlxVHYEB     400     1f0�%DrK�� �S�!���5Yt�?%@�z�h��S�߯ 3K�3v��O�b%0YAڴgi�����ΕY����U�uԙ7�e�K/3�B���m�Oփ9`�Ȁ���&��e	�*�����-�A�hB���4��g��Y8.�����h]���Ƥ�E�fD
��/V���z�#�i�=f ڇw��f/����&m�T4iz��H��`��5�c���l"`�?���p,��~�e����w5�9��a�����ǊW��V�4�g#th7�M�C��Yuu~:zܗ���d�Ã̙c?Z��l�Mi�S������C �U��o\�LkD�a�/�Y��X�4ؘ�w��w���0���m7n��U�j#��eo�6��Z6�~�.�Y2���vs���{Lĺ\'c�Y��q��G�x��ӒXU9���J�[�+e���WA���N7+���/�w��!�ट	8��Y-ۿ�@��˜9�(�ܱ��U.K�Tv���b�f,�I.p�ʮ�Cԏ���XlxVHYEB     400     230�㟐ipe��n�����!�F�����e��1/I�@����ˇTOl��#󃂅��#>crn�%y�&������p+W�u=@bi��HЧa�x��Enh'E�K�G.<ْD����1V����_Q�㴨u�[5z�L$JM���='�S���7!'�bB2{�\�xO$͇-q\� �"�ţ��a4��IV�Pӝ���3^�]��R�nf;1N����F��Bg�Id��v�E�05�	[��ð��(�Y�Xي��kR!�ӵx2��|�(*�����'�����
f4Bm45�hU\�ިZ�S�wA��J�
Ӆ�j�������N�h�⡖O������B�����y���b�h���(=�v)�$����N\Y��5���VȮ����7Cl�Z�È��"Ɍ�5n��Hj� �*�������&1�!V}Y����R�lsi�U��&^e5����O|/X�ǾG����3i��Gf�B�'f�M��z�'��~���?1av�%�]���bxM�pUn�L�(D�cFy#��\ʂB�A�{�"0��9��7 &F�XlxVHYEB     400     1a0�1�qv�������-��u"�/�'G�q�Q���).���Zc��yO����=L!:	G���d$4E/(_C^�I;�wٻ;��CL�˜9t����t)�6S�$,Ն±��q��A�v+�bԅ�W7Z=o�D0|7�ɵ�&Ǎ����[����j�k_4�?0���ч<7�����[����2�����S��{���:�&kg��R�~�|���#K�L�:�!2�:�@JFsy���F
ߎ���z�R�Qm��� ���1��X�s>t�z��ú�jXs%��q=⠛9����t�#��OR�s]H\-�~L��<j�wk�!��N�i��>�{��0]����L=�=���������s�D�K	4��t��W��C�˘h���=h������t�XlxVHYEB     400     1a0е撫���K�.��@�z�]0�v��*ʸ�}-g1:o(֔�T��U�4/͋FR�aT�}�ڂ��c��X��b�����[�J�.�X�*��A������%�����M�ȸq��ʁ@F��0V3!
���u�[�3�}Ӻ��y^����{�����F�mj�^2��Lo8J�qNC׳���G���i��2_e.x���x���g��.p}���Z��՘Z�"J�k�_��^n�r8��_%��6-����,X'@ud����K�ɷ[�����Q�X�����Fs��	��ВU��Y�$v�S��e��4��:�����.��l���TA���ug��fZ����̉yyo�S�E+�k�L�hY,��i?��	]�J_����!��E.)q\<5�hbe3�%XlxVHYEB     400     1d0��4�f�ZI���D����]X�z�F�T��K!x$ ��4�Eu�G��-)z�8����l �w;	���lz4��|���OB�ռ����#��<�_Wz7�\2j����%86����&���q�S9*h���l^��]�_L�/@L
��z��y4�9Z8I��(��7�M�5$�r�r���Bޛ���P.*V��1�=\�i�ڳ(qt��t"��ܛ�+{h�٣)�s��1�99������X��p�@g�U��*�3yժ��	����):�f�K쾳f:ydDM��>J�$ԥ��h��O�$��0��o�afiۅ�g������6�@�J'���z��T;�K�H�e���W���K�_��j�2Y-K=��p�ύ����M_L��~�oG�t�{�� �κu����q� s�oX��OKZn+�g�֦a��6i
m<-�(���!��!��;E���� [n�N�qXlxVHYEB     400     170�<+p��= ��ς�=�kw�c���������ׇl�-��so㣔k3�51����=j<.P������i�!�s ���ɭ��'�j��:c�S'��Ƕi�t�M�c��{#�8dX\~X����XkB�2b��}���
�>I�;�l'leG���F[R��z�d�'.�n��p���-I���d�#%�����釱���G�g���(�?�r>����!�[�1t+�;:�ɘj|b�.@��0�^(�7�/�	bڨ�Y�,���o��OYO�E2�E����s��]Bh|$�HK���NA�����.�Z_k�#j�g���<6<��*Y�_�_?O&�1g���P��s�~R�m@X CЎ0�����p���cD��XlxVHYEB     400     1c0�3A��BZ�lB��z�=;�̯���b����e�hљn\G>��|o�"�v��ɜ���[O"��:���+CAqR��a��3�ĕ<,�G=�G+A���)L��)��>�˰GRi�����ŹTW�2�m~`.�P���~�Zj�1]�{e=;+�0���<��!r�D��=f^�$~H�pI㟽������Sn�������|�9������/��Qߎ�`���j�r���ک��W�;#�wg�ܚ+UCת���c*�ulb�>g��Er-���{1~��?ʗG�����n��C/��R��QƏ�4#iK?z��̎�W ����B�\�&���@�L����lZ>Wf5�~I�~v���b4���	�e�d{7���!J�O�T\W=��A ��խ ��exX�����đ�y�8�m[x?'����z2<Æ	�jXlxVHYEB     400     1a0�:�`�ɕ��%������t��B�F-"�S��u����v[���'I� ����m�=Ϻ?�	�[��2��}�9���Dc�ζ'fq �����>�6)��	m7M���p&}Y8�$%ݻ]zNC��˅?w���~G�� C3!�AƼ��z:��Q�!��$���]@3�D�B"1kp�;j�m��},��4h�ye��e�N��hN �Y8�ZR|�����"S�Z�ء�w���N�!$�j�C��ko3�~ē)�Y�5 "\�"���S%�]��K��3����cm!�R�Y��t��dK��P����I�S���K~�B�e��v�Ky_�j�W)1�7��.J�?�|H,Tq����tS	�.H��d)�S��)s��_^U� ��gm�]�/
���*B7�XlxVHYEB     400     140����29�l�͒��%�ݍ�s��IE s=5���Qd��@�2+B��_E$hu D��${l�H҄�c�s�� p����ʝ�֢���X*�9���;R:eS���f~���/�(�3�o���j$�TlĐ�����C��\ȓ��ML4��F�h�9[Z�:#����R���u?�K)�jGa����.L���c��5c�����<�e�DG���G�VzN��H�[�t����c0X��i�k������]��Z{փ�9��}S4ǫ�B/�8?'J׹uQ|I��:�j�YŃ�h3��Z��ڴ��9zXlxVHYEB     38a     180�2�G�(��~5r�6$����Mŏ��=�� � ld�$�iݢ*�!�r)�D�/�
��W����@ٝso�gZ�
0���tf�J�xd��B�}X �k�x�܅ˋZr_Ofk+J�s�FX��)�;">����_N0�ۓ�&a���<��@�K����ܧ�ܶ��~L��5|S ��X���>��L�qf@Dc�XT���@��D$S4�O'N�j:��w��X��csQ@[K.53}��c��C�3��\3����t)�מo��9^�P���� ,F���+>sY�*�Ű��>�Q&�BR���≌������ݐ1Q���H����D��Ga���>C���C�����4A(�xv�Y�g}w��[Дz?�>�uHKS%P