`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
XCcNdJlvr28nqpHqYxsYe3YcwsBAZxbASOyIRKv2GlBMkRthESaOkoDjGBLyLsMTegDyWkFYX3Er
Y85h/ZNyHIl6j9Axy2eNLAySXiPZtu9Y2JJKjQCTgGClaY+CdaboG2R1nFKzysmRUz9sPx0R0cvq
7cdqTvnYWCWrrqd3DWIgEz3ypbWwUjb9798+ybXSymVVTGmH0qu+1VWlP77pzwMtV4EFE0Va/Go0
J5zXU25fsEliHpkz1DqsVsQsqznlWjz+KtqbVUtRlsCpe0Q7rSrO2PBvLdx7I9R6TIUeMAeuE8vl
09ZnQOMpoTfA9P5AXVZB2Lf/iWsNsV8HCvSqEw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="aUuxJWVvqwwQG6pXQINVFEi7Rn78JFA9Y/2o1SW668I="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12208)
`protect data_block
HMBCVi9mGE+/AVcFmcWbVenWXRQMm94dxz51OF0Lrz7bNKYXD4I+K6PfCyo3+7zyHgazYTHh5dOZ
aRxDajpbUs/qmM3w7fZz37JUwkvnPCBdS/2lBZpaCYHh2LzpT+HFpeEgPyxs37raT5xE3Fe+IjQE
UAVc8baBJEfPYalaKSKgXW2dyjYAIncmH/Hqug2rNFBR6p8+7mruj7ySvQ0YRkyzLuDw0yBIXFbn
KZopy+0juZeQ+grh38Y/MZhZ2Y6SJKsnxW1AACiZbDHavcunBbifG6Sw6goVkAHQO8v1WEDE9mc9
wSH7E1/0MnbmT3fUl8/Ck6rOCvGU6RW6f/1eJGd5UvhCoMvyT7iFzNKRCzd26TnilLdbZLLaCf/f
U6ZcN4wnGmQluK0zHohazTviCtfArCpEszojKDLHvanVHa4lJ5erYpdF6OfSvxKiwYaQif2TvW/g
I+0MTecOx/V2Fg1vCalRxyhFb/seGqSq1HG/QqQC0ahkqrHlmD+5KywCDwtTQCngraiu95QHBMIg
aGpreTXoqnKKJch2VBTE9akzIqGOByWcOYBKJc8By5Lrq0zfELIdw+8AvYgoYdInDlq/VmS+IgGM
CDn7V/KQ5U1zhGbewXOABRDYPh/qnatMpq7BMiu7BUj1805zYsPdxWajkMmWb9ov6MN2x+FqyjnU
s+yyJQWOEmu44JfNjQYNPuLpBTkaee+a7bEL+omPZ22STA523f32HLXSHjNCf6v0HRTc1wsiI2RM
3N+0XaCdeL5DXvLqzpSVTzSi8m6SBVPOgjftw+vDkTKp9+G12AZyGdwTeJ+am/r4WMuTZnHaB9HS
u2ahgoWzuj8CizAM5K8Ipa9yE+daDmkDpAcgCE+4gSZGVGMlbWQ9l23t5IMceKTj/7aAc9PAyPTI
aaO58tpKpzkM5y6qN5hVXHxkvz7n9UaYPiYgX+YKk0qpCpGQU0BZDmBoYKoy10QetMlXcAgWhE+q
zLXdcVMWx0/gKlADpOs3R1k3viItQqVW2P5P4Fw+SQOUa+XWSE6Ti2jVCofo4putC2XzLI7HcA3P
UOd+M9mfm6as3CI38664IeoQjlOi/2VxDpfcY08KE41BDmgtPt1CsbnF0zNFE9OgaWztmSykkJct
yluQ7TG16WqCgjfgOFSnJmvDJLeC0uaySS4sn4GiwycVoY6XyikDq0EZaMbkn1cOiIcua2w81oG0
gADnhRTHdpzOuTr43wKFDUsBSrW98Hl89sfN9wzwVCGZwCsa5BqaASRr6K8s71rc019QSZ3gPy6i
3pzE9BAvTxPpnD4yJu/86wIvq1iHoxesCiTmFnE1eru2juD8lniE3D96ZzE3H8C7VMlE+SbGw2Jx
icRPLWdI0oKePwL6YlIHC994lBEPlrfseWi3pA4MA9MSR5dXeMYad54RBbVi71HCihoAL3NitjB6
OwJr9K8dd+xg3dNkKsyouMxEsmhoYLBmiatMp1YVth6N3a2P/jd5NLXobSbnnaiTDqQCp1SR8+XC
Btqbp9+T8eV3e2xFmJo7dPokXvavQOfl3I09SRivCdmFd+CkfMz2f5YsyiaJQXXNDl8h88IiBu2E
SD2FenvVgAp+b77OafIHn3YFAtL8177sEo5P/q7qTglm2d4ewdRcnt6dpgEr4TLYNw7tey/6YFab
JECVjQZxy14ynFsqDcxyKxerHh2nu4hxTQ29ea7tkl5WzzIXve3JYPabmVUyfTUGfPgEeBjNlVPg
5Tih1vI8ZSzr1pyC5nQKjW/YwIyWzGkt5QvpoRhPMc964DKIm0JYJk0erAB5zByUFutaWa/lrcbD
6P6Fm2AGlSaRzUqTBT6ZssTcKEuxrDMK1kTzgjVYkY1AgaIXkMSmi8yb/s9+J6fZwc4RyL5iSTQ+
0u+VDdU3QlR8AelCGGZNgvyDyzI58umNYWzOpsIKfphGw+l6xJUFVDVS0CIGjntexBehIQufjuNt
hNhGSYfUQk30qLUoxxttsMeFyoMgI88ItabuWInUH7qnttsgXq+XPMaCnyG9B0UH6si0oiF3YbWt
KefMqs7tXHWrw76ysFByOBKHrt1WuMJsqP0LppPayDW9ckSkK+KCUPEwJCB1ZrzEHoYMrGEfUnmo
/2BPA0DJjBvVauSXh49Br+jvnaXHwEkb6dhdqsEYOogaoCXGA/72XiSgH6gzyVmX3XGalTrIpLNJ
MoUdingORBsCGusfwNW6Yx8zgEIyba8AmDfVDDqkanaqbZYSysxlGprklAEwr7qpRFpB16I46OTs
KP3os1HHvhUD20zxBxGa1MTFKIn4YXpHitnG52Dx6QeKDAW50GTOPfloxT+4vJ6QzhWrSMLX7Zu6
tULrbOetCC606MomPL7ASckNX520Vdle4f7Q7ULmGduyZ1SpUUb/GU1o2juHsyll3Mgkv1ApKDbu
QqY08qOl4dsPAvK3HsyeVT6K5EydBbFrzvAUNzI9OgrXq9gfQ3Qi4AnlMqw5dfnapBEJSHhZC3P3
Q9coRz58bQ2+x+obsE6H0LI7mYx5G3OzFA2R6oxyU4B28UfocAoczfPqh8NLTSWx9bnwgi6lovcm
DxdSB6k/02dioaFcsYDo2Co/Ip25L9IGse/2aV4EtwoZ71Zk9DqUUkaagoLH6YIbMOHUSHPaJwGb
OcoFcCIfCKiUrZOAtCZH3cMiQzR5H430+fKXTeLJULHaLfkq01pjXlSdp71q1TONO7VQ6MYuT0yZ
iQhNhUT9dcReNocHuB32SWbKiSseigLp3enThbQC6HHN5/XgLAJ+7ERcvbPuPVZhKg7hOFuMroWV
EFO+bc7JMkjWYhchO+mR8v+xnt6FtC2nTkKBsBfoFq+BCjdocimDpIQJqdcifKwKRoMg6DinwYs5
63udU3cuYZWoZrI3APrfHH5rbDkp+AzIXaNII+Vgn7TZj69YqYcmplB9ICwm6lUxVAEvC+ZHJ8tW
0u+Ejo9XLwH7CcK8xY1BtVJY+5UOySsvkKa9pL6uBn3dQ3LlSeATvehr63sHs94gKFVRblAWNbCM
6yhFfpeDmXEw0bNWAkISVyBY7+CPjf2jEh3oUd6mPg5hYoS+i2F1EJSloPluV1+E5H4SVkxyIwBH
VauUtWniZI5EwOU8fPca1gjKbxdcskE9338IoU+T5w54szM5Eqeiidro/BOmX92jwMlAk9wL/tBW
6UCpkmjXwaYXqJNhCjKQzC38bMemhVctQfZMJBs8g+h7htNKExJ8RWGls8VlOwhRgD5Jb6VmxvTH
lxKU1pHE6QAJcocAebfWKaiYyCXb7hxiby6EUAG1kFKpz/XHirKuv+Fu6ELdQT/5xbiybv8SKJBn
GJf9w7v8Mub+X0VIk2BW8wc4nJUGzOH3iFmiw+0+gX9mbAKojgJZiB6Z3dyhwWC+NyQd8elYiAYw
UNQQMtz/SEB3WI/nZ1BavclWYbBS4x0hibfBk8VXb/7I5JQ6GXHnyamqldaeeQ+wggBCS0TvRjOq
XwOPdi8+mFRdRzZxYAFJFRKynnjMxI586iGLqAnNeu271aICVuxoUL3t9JNeOfv5LdCw+yuhJX84
iw8/Gbiocij7CFhZaV7Gdyw37xaLwk8pRVhj2wII1C7Oa870hVJiQ8aLKjy69WUTYBc+Hqt1+sKS
NOjq99Y++jJHqU/6f90p/HhMfK0kimsGIU4qKK08yK66P/ywwrOds4BPEn7I/c1vQalfxrsx/CDY
Oin8rn7Sne2az/waw0ymZ48oYn9jhhd5sEbi2xQWlkieoNWy6GYUc5w6j/MhZU6uX+11ZbIzGBp2
XguG2PZkTeeE0xvCdADb7nj+NcQtKnL4mhHihuSnr0bpW40cMUOf0yPbLCtZSHDsAyVWKUQ8Leo5
8ODYlNuipHuA5cY8kN04dXNOu7ABko3TioelqZDdhJrAlLLi60ZSJ7tG1B7WZ9q/E/KCwu36CQB7
xikcA3okuwXDa/fWnhzj4qGH1OjiIrreCOwbu4iWBAy700PPiOiaeFRTqKhbjOa/vlhhJtNWXtu9
42xi9B3YKRhEFKlQp36itUrMyHcO64slqJ/1uXwU+NGaNSJgtevTApC71rgHc71Q2pGgacJUg6mF
5lwsjpGHW7KYn6ei2KS8uNkdRuZvYmZUL2s6fiWqZj6VdTao1OzUUPbZBbT+Ez2JH+c3L22HHepE
Y6GEtVUz9l2MzP5TqeetuCQMFLXC4h/Y4U7CC/usADSHaitiOIR5r8PAxR5wdRFRxjL1hvpdC8JE
7W1QiUWU/La1XZfIebSCyDLmSUeZLouYwXeYQOuOj9H2AFajle0zEjHahRZsNYoAZ/luf6z+Ze7h
EyiMFZO6Xs2D1b6mGan5cc1jnmoOVWyrhFtVvkHCzFN58zu2sUfuNev9yDlaL8bTY+KCWnXYImBz
wCHmaUEnPrbhQFp8ArBUPKrtTT0PFPs2df1SinYfNWKwGlif23MBf8iH5CQwnqSYdMbBHkoaBAim
Dc8PjWFM0flozMIVQ/WFeV1nGyRYRGI0iACdLaPe3d3d2owXsJnoplmbOLQlQqQDxmKm5afGUk2s
FCYg3q70vnunWZN+RNfmYeL6ZQeKngNBc01sxMDaBWosvSj3lD1Sg6BxaxctSXGFv6WLe6n60m9c
xpsisuJwCSs5neZGVhE5Sj5LMLzBG39Hwaoc3PBO5WUY3Vie8a8V6FH+1wvOWuidxbyeaz5nGqQF
6ehEeZbTDFJyhV2igU6zHn8cWWtkmLRrvOv6g0B9Eah/nKac4409xfWh3HpEAcyK6uqbB8Kdf7Jc
OoUp0T+cxxom4kvpsXuX2Mn4QlQmG2+Yt+wQjeiLfWL0Qr3GbN0tGCwoAScw80WN48ShWupGWPmA
KA1TQ2Gc6Gry2jfk5d0/FidsU6kqjJsSVO8GUgGGvcmAmsoek6DbZjSqFudiWCb6CxMTRdHlOPqi
5l6446n/LyljfrlhR0HmM3UKSZqfKQoFz+IHTj2pDtcmOPJa05/WqKUvsVBMjZJWbA8qC7bZTeQ6
JFkDASH/ZYZOpsPEjTowFPM1ZSAuGzAHIwjmAS8RQeJYL7vBMqfLdeurz6FQ0S0RwFZj76NLNcQb
gmiC4kGBMvnTQ/nREVfBlp5Nlu6W34GO++WGxfZRsjZcfQDN+OF3/uusRAPBnhpWueNIKKrfbfxa
0qnPoou5G6uEVSg7U63fELW1rAVF258J2QUbOGd5kpkWFHaBZ3J6eGHPG+AWnNh6EjAANYAiVX1b
LUVOwnh4Gxgcl35RkmS6PgxMwj7R/o7pkHX4Nc0RxRDrWzRo2AxiKQvzVDT6mVQ+dUNaEGVRg8hP
YN88+Zvj1+fz9rGsxGwuof62xfJjy6bSWM+/8cjGR1CHPgrgMNLFI+6rjeqWlMwBh78yzLcSMQJ7
CV9b17EHkbpj52ztybHNqcKUpa0drD9aceAawdUt7oxmJNxABKtR1HwiNJyTE8ubw82rAxkMkhAo
JHBmEzFMhV3SDZc+FuwsGKrLAuI/9Jm8CSnUJk+g4+HHl9BbuQeI25ZaXi7eCgBjwpVI9UB2B7dL
nyAu4udjb55UB+6OoIR1EMhvhRZQLIZLhvxDRP7T8CnbGe7U+Z2/L8mT4YLJoJJkhyTohpwWwKRH
8iXxVwZjciHpMXXKwJARtFzWLRqG/kclVrZAOHnreoYYJcoqwrgoHaGKuWof5WPmJId2a4SJFoqm
u/owXLFnkTYaNrrGUe0sBQ39ETdL5T9xA+3/7G7jKURt5vnwJ+8CxbbyWIf3w1QlMoLAKEfEZn7g
Z6m2uOV6V1Ftx9bzk2VHi+AW8c3gkMbRmY7zf0aY13ZI8vRlOiWttXMQb3W1YKbS2jxhqV/s2/K9
pwW0EqvA144AOS8+CET/+wvjQ2+mU5ibIChXQ2vRhgxNjp47wNmLA0A6f4ldtaw5FZrJhEdIYgCn
fv1KRyCildvbbsCdyTvsiMpTGzRdqhXvs+5BbNg+b+weV6xjGYJSJP3kvch4v0cxu7SptswQC+7M
oSWk0gmZg+pdczN5Ipu6hzcF1shN/J3Z7bZ9JOfXXakuhegeMxbFfGsbDpteOICxOuNtY5FVEdBT
BUBI22D+Recmk6M9qbs9IOfsHFiAi6WkOLxPdQctZvkzRxKHvfbHimvZqDiLqpO2bOxunDQkPUB8
XOmIezHG4VUSivDK7Pb0eQF0aRH7K9hBt2UiLMejJhYU2CHIDaNKPJpQ/OG7oZkhWkaRTVG9Fzhf
H3VhCzYIKcB2helpVWme0b4GRV6xb4h7sKzdP+qXuurDiQa/4egZWCkoMDri+rAdOJFg22xS7dc7
pLGVk41Q8QIWSH8UkYa1Hk6qszyrkUbExdGjzB+0Kt1q0DxfpZScL9+PgWvj0btUv4M/1G421sN6
xVSCcV3JG/sZQLdJSQggJItCOvYEXWBpQ62So0a1w8TJ8vQFGDNMO/b5M9SzyHU/niN6vCv0wc3z
M+r2ZKeV1uUYLly/uVmIHQ7ebo3zMXAB1tm6+R/HRoHO+t2zzwsRIegK6qbwaZ1HI77t9SI5zUeC
Ce8VoEW6akctXGEI1z+n03l33emSa106OUdn8NS7LN3Mjl1bOq0bCtAfu6BG3XqkdJvMKxrb33zA
QOCJ/lHuW/ZPAvHobxfmhjGLOqP5JHyglDf/Fmd/2dVfA3n5LMCACbYLJ5nbQBjppizvSqK4EpZF
CtqCqRCSb0TYEHmtjn5zNCQWN6xJzsF+imKgsyyDcnp+B/d3kPmQW/FO2X67J4+a/Vs4CPEljKqJ
Wztz7/rc5fM20oV7/Z6k5JfGmmRFEH5WwSbOxiahrD1n3s/6bzoopPNLALCCJpuPGU/TUkPPp6uT
PcOh7hV09qM6zvwn/eezzI1XgUW7qfad28853BxMHjWVbLXpPuafTrrt2Kb4WGJNPn69TaTue5i0
Y2FvVyBthE9kLPOXCP8dvVavUSOHONnaWqoyYEAMdx0AxwUsMm45hEOhQEUKDsCLudbt0xgEhehQ
m/msNqkIOTxgIxhv/YxptWptymiUnIdyHGcBrUZBfnszNFvs/sZt7gQfu/NGCtQc3Dg+8ENj2itg
hUp4uy0a+23G4PZghp9DSVDE6kUIWutSJuNSXnzpbgYKSNQbf+FOSHAKBgAyhwy9Bs7OISbB3chD
OmNYKk7XUj52CIaAg6tXF2M3aWW7uyizdD2GheZsWZomzz7ebwcSwqfRJbIpCztRPfGhV4n/swHR
i5eVp27t/01MabwtVr/wKfv4fAenMzL8KTwvLVCXEsDpR8JQ7jLZRUiTRT/363M5JfQHEzgNtkE2
+cSwSOthTrjVm0xUioJ5KXhWaTc3/yBDkTKXf2c8PdUF51J/nwELdSy1TJE81T+QLWdhXxCsCTAv
V55bGtvpE+xDvNC4gQZ6D08fCfQNBG9+3IkLXv2MXSH1FfwFqNfaEMp4r0h5ir9xffITXiEllosl
zDY+CnGlI5CLXBKDl7NszFQyXBSPCqP9u1LmfyXeN1dQJk7uLuGwQVR7lw/+3jv53i9sQZKrdF2B
hx4Xg5jd081n2B4Me52+CEAVXg+pa3yuB0B42yZT/zMcp7Hlbp8lOSPHNLgvOVNlXYRciT1dBkXz
SNDOQ6kiNFTFwArsJID8Py2hEJKaMuz9ltE57FN0tTWeh1sexbsUQGGKGMnYKip3yIefJbSYRAty
GkEaXTWCo7v/5mr6NtrkG1n2lEfAxK6NeyLPe0FjJinlt0uACfd8DtjOHM9A5TDIQvLo3H4SD6WA
nDu1ZKqx7yyPXgl3j1TzxPS3yks+7y+k5xms2TyYswflPRs9p0NKQ2S/s57kqbicmPKV/gS7zthG
hXDfJIxb+hsOC4ZxJ++3YoCztKGyyuQ7PNk7/XuGTOWIfPV2a7TEIaF3FdK/qybXlm6960ni7kJ0
/DuVRmZSkYOKWKDg4S1uccqCgjyHLR9riNK5uv9IdoLSbgh64GrE7bVfs7gsJd3vPja2dLxg2tSZ
NQa/I6gr2IwdVJHCf05/PGAN+lK8FqJrDKkOGccge1pS8ojluaXk7TWgLheuAQ2N5wcWPXZzBlp/
bWhxQnK7XucQmNyOm+y5isa0MwrqfnpEFozh7aaC29/SyK1b+pfe6Ss3/RjEPBragL5MeG647PuO
gS9M9Ji/dsXkMANP2UXwuMIdSUy5npG2L9d1PaOUUwKPMoHYz5VNMWq2sXX9BLwRQckB8ONnXNjG
8RJJOof6O1eT6CaMHQapzA92s6O1vA5VOLuEAWnaepNJS7INeJSV5O62S4eq7DGyx+P/ujB+u0Uf
HFGcJycDYrMZ3IpSdiW/ACf68nG0/qb3r38kwgZFpdjxIJgmOJzpTU1QHmFPJrQaCRBnOMSx879S
+gZHEJoKrQZPeeT+C+a2L/y/AzuroXP+aDWvEfdSJkADTiDybzQYfyqrFrmyWEOTLEZvYb3TXQ/d
PS0pepHYuTGhRdsWDqEHCzIRfzEAIlBJBu2UKhE8PmPmHZNrtMatJm3rpjhX3TqjgO5jVVJs92Q3
ZrfSR2WRGQMgmd+zCXfXGeNm6E5ArXFSHrCz0x20NJcPBJGvGSKF26/gvDqqz0nKP87T84ZxRFrs
Nqi3pJa/0XgvEBEjXFC6OKANLt71NvuRXupAmGfWYgwQbt08he9sGn3ewyWzhTGA7WWl2IP8MzxP
hncghKF0500DOmUzQZLCR//xQGmVwaGg0yybRTGkfZzu6pGPMf2db/jMxJ7luYdoDCDSMqCVziKx
46i0FqX3VciztKHAlNImoa3lXMnnhk8vs1bdhC5GQQN8XIMjrscaItsRmAOCsqSD3FiNQIBE9CSR
GKRnFoC797dpCzhT9jrNnJC8zSKKPWqBy6eEfmTzxpPiQgXrLoN6hL7EYO9XZMwuZQfg+EpHGQ3i
X1KO+9iOMzhjI/YmDYX7yoNLnL4fdxyXuZLxeZtxyhq1rY3gn6CbdRUXUseTN0hAC9ZGcrH7FEy2
896aPlgQxO4FvMs6odzK1D10D42Hzg657Ex13NwKW2g2U5oJSIP8PiwX+kDB+4FW+y3KOphDN35J
NwolrUXISwR8FpKPbiXrs49KubQZCHeaxXmj3TV/yNNivmYbq/8/Kt/qLPlflzsxPHIpYJT6taNT
UPtLktSHTxERqdvbc68nPGJhbWy0P3/9PoJCRJ2NOfZmLbTz8TKeJqhQ1uCH4EjeSrgsshGqAcib
PvQyd+IBrydf79Yy2yoiBGXDnQeWFUodu44NXDsBwq+CJ8sLOuSj1qrwfRkG+h9SYQT6W4nA9KGi
oUgKs5vGF23EtE6v9jbJ+SoBpdHZhQl2CnunMQBJY14RsEPgy8fEjWVQBOlYabCreRniYhuB1hjI
UTGhuma77PJCgkaEHFyIaNootA7CFYQCw1Ut+2KOot0R3PA5vxLrnU+qCHgj83s04j20vJ46mafI
mSVBtY5zfJ0Boq3dQGsB2/G3rFC+ngLfGX9q22RIEdwhu+WTVsravhlvpZnCGjK9xhIYBisFJ4yP
XtQDEo0FL6gF56FFKySJ/DFCTFEU7Jez2xBa7n/dK1WKymNtSzRx5QzuVVnCopIUJHjvR42X6MZn
+9ZaUYS21m1OSAlfvIKxJCzEQC3VJHqvWf17p41nqQZwnTQ778p5/bOCxmN53aJHNqjXE3mpOsra
aK4QTXHbXzy3yHC+WL6QBQPsXq4og8IuEJMIbZZyLLRpcbktaoY9GCv8IW1xQoUcnSCdOJzrWAyt
roao/gvxeb55tGr1SGRV9vUpJQXjr0ARz5P3TzkBRQ0He72jiCpwekSEguMhXRy4QYV/7FHC8oO7
kox9f7MDDfKb0cDCWisq1ogWtAluq+7dNl35/YTpBZ7b8V2eSTZT0wBlcwbXama5Hq/J2jFJLMJc
hriQEVFZiN6XomlmaSqbNeTzkfakor98GUCQBNAka6cnYmLW5vXgF3Xa1HpfatB+o6ZJi3Ve49a2
HUrUf9mux1Rb0/0rvsms2dEFQdOnTuDjZZrINsSAR6RDjL3JfWVbGrIRe4O/BDu2QjgmDa0vCccZ
msNgKWfclTMzO614zUrazJfr3UkrNgjxCEa9DqswXhXJGyb7PrUdMizzmNSX4KIVaFqm/82SI7/c
w+T8HLObfHA1QU/Jxfk/lGIDwwkNuJ1Kio+/l1oRa0qC/wXtCyiKKccoDlJlpSSXCoerqQtQmw2D
ze32Q0B8+88ipLTikyL2HKnsOARU7E1HEUEUlTVAd+tofOQHJpV/Ia9g2gA7YaPo9gnhAn8THcwJ
MKet6lXZbEHe+R7OBQ6q94AJL78hPMFsY1bl1L8pA8GvlqahIWzEtbqkFYzjOhN1OPSl7NUC+lTi
aX0acyAOJ2iC3JLNWqUhbwNueHsi33gG0+dq2j06JsLkv8Gpjv9NAvkoShspddYGnYfPMLBNvYps
hmJwgN12SacN4lEYVDlebkbmM5ZI57n2bkrWT8/ES0nX1e6txrDOaryl/l28UIQ+lZNoaAwThIId
kN89IF0frwX8e0l11oaXqz7Y7M4wwkjjfWbZrHMqaMELJ1Kmv67CmFZ3K9z42w31q1uOPddz7kN0
wZhSZtLEWtJQarhjUDYz7NT8d62LzmNd6967DiRiqvVai/xwj84tDd6wnaBQZHU8nksqdKoFcCR2
hOPtOzAFB+C5TX9NsTFWwvpo1VaI38j5BADZLxcUpuCZxRcWJGbMJ1kAO00ZPNcEr15U2n+/HEk5
5jIjL0FKpItR/uhnUVvNk2LjAFcaEifJQ7OHzaGz+51mnm2YXZlb64rElRQKKD1RwDxOG02uQyQZ
ZB4lPbKvRQ3nYK5WEXCj71L/7Ff4eQGbWHgnJCdLIvLLF5yESXY0BJuNQgGt3yJX0+2wVDn7nD1f
I7bd+mYasCzGgKJvyuErVuXHlIgWxs+cBpSAm4E0eOU61amYAPuWFw2HvH1ePyxN8czsb6lVeCKc
j1Nv8Ub4Yyj4Azqnid6cgd8JUCacRayUuzdEvzV6d4UHSMiFOBPjS1I6PTXR10dX14P0uyQr7/Ym
A0Nfb9p33HodygoWTZx8OVW8HG6gNB4reTl+gkZL+Eu6kbsVs7Y/p49TAdlE7tisxVSDhaEMhCa6
f9GoZGAsIMHeiAza48S3qPYXqkiBAIK4oxl2nmNftYlhDx/GMRM/xKQKrsXT1fwmVTyYempPH8NQ
nziZZVJEmz67oCpw2Gf2+aT6hUh85/Re2bKg3j/9rWu53b4vHjifvh8zy/UQxGIjKB2AEjgXUnoe
cr05LQCsK7RQwFwCb5eNz3Jgjy6xTgr5+PIUechBxNe5MhkHHwiIOGCN4nV5LVvN7CyzGowEXy3a
x1rnrZIncOKFoa8wpzpPnxZ/19jHgp4Xm/Ig2knAHWp5sPmdZuU2H0Yiy+RffavKw0BMtTa6S8Wd
AnEW9BvEEhACXiU3FiMwJN9aX2GiqSmBGm2FgRDVHUOyTZrWBes7uGmgGL8QMj5p8XH8bBi8NPMa
gdcOqo5OvHE+dk+buMG6h7O7wgMCUcqVIVZvzKCdI1sws1R13u5Vw660nyA0jJMUrVQFBhAtb30i
feJRdBTLyeIKGSft9YdjArdtt3IGHfk+Gt5OyF/TWYhNqfzI/0PAVUf6aMLcTD/E7BAMgBJiJcKR
yVPFhNoywH1o1mS5f4rVKy9RbkoiBT4FXGoQmU9u0QeRsmV78BDC4OE+k+/rFC9/WCV0Qg7AW/l9
pn3InIfkZfpGFnM+Fs/d3e50AfJxS/bZ0izGWIjoyJw1L+0/zB3S9kRcBeF51ngMxhFJ9nQZHSDL
TO8fU1uWrwqoZNAHgpDD8Px7Dj8yA7wbkRghuV+JLmBuD9MkJ/NBxW5c++GBm0Zim0YnL+eAAMlQ
s3RPxpndKj7zYKrfALj+LE6Dzw7yenwjzJOi/pqXXocpCpxKfN8phPyAwAC22Fmx4ppCohm8hWee
8zNd33wNkG+DrVWhzWdy4YENRXP6UBmagWTYyTOF0sDAfneBtIgF77XBTIJ0IkNmU+EPAoLDDSPL
g1wwmp8f1Wxyg/IKuaLQLIJhEJUDJfRFjvP/sQNi27go9nKIoGbQLe45QxCvl+5bR/cpJxEOicQJ
6udRxOrJTcRdLQiWWF+6WaFnnIKedrAYG1Lk0NE/dw9pFMI5DiXbrlUuY4qxfIiM0vouu6tEQSKN
vCLo7bSpgtwXJH1oIv8BMxmDe8FoHkVa/AHncF9fTVfy8KMBBhWU99R3kVswrbQP/uEuEazwArc1
kJW0q7CtJWSt192BvBOdWHHD+UgltTrxB36BDLFmKDTwcVJ+zKbBm4d0PFdKq1YZAkD5AnS1nljH
jYkvEhtcFfeYLxJFma93544omg4DhCZGvtf+LAt8DaLTlwBidZ8IlcgyJ+YB+702CSbEEROlXo9q
aUwPJm0Hv2FMB12B3ZlrS4OQLrKlWlssmOOY+mzMMLCdsTcXxVfj7p/+CZAxK+dZll8umAgDOqXY
qG9dfKbuuNsYnnyn/QwsLUsCSTTxwcC8ny9RMOaekOQK4yhSH0In78ta4Sa0hAabPoJXewJzbmBb
KRbBgvD8RpldQOtmxzuTpc/0+Myph0BXR/QIEwm5fYJ/BnG7EgX/Lh9901UhBStW48XDwKvtJKWc
vxLZPKy4Xh4ysy1cnZ+Z+mtJcD/VWkvSt0+QvDoest5zgLMf7qUolaG3c+0AWi5Hv5DQGNuifjP4
DcskrWfyPB1/ekWVd8p2mAJ+VsA+wl22t0nOXc8zLrvZ/3cuK28OMa2n2HtfpwgOcN7rMh/KC5JB
vlk7mAqWGPkk4Uqtr8zIWVU/JcSeCkiY7xHyitdQ/S/u+XbPEV4+6UJaI8vK8WeXZ7okkNTxWou0
xYauQ0mzBS32bOOKHBajlXZUaO44SnhDqp/OLIQ/Y/S+dCx7uwVX/l9f+X975rpLfznsqHpzxUJI
H098/LvJXmcEink4/TXUxObEY0hP9NqnfeTGwDzXhyGIy+OEdnL2/C45yLwszYGlrVxqcrTXyFLZ
9X13sDoMaK7CGTVdARuRF8P0rjYAoxLrrX9wZpzyYOEIXFw2p3rwu9dS26nOGWiJpq2K+EFWuyep
NCJMu5duol+JfDOWT4c2M+D3Qnl+29X86Sna628/Z63jd4RSXnlraynHVVCVBML4avgUxqvek0ww
mc8UllmzgJxht0zHkpZLMQw5wkJdIq6fotz0oClEwdIiXGczCY/wR8Uqma09gTOmJup6wGdcQV72
L7bMAilZzDJjaTosy5GnAJCS3dx/E/v2ivOwxYAkhoFlf/3RVISWNkxFnnIn4xNdpWHyFrTAlCdQ
sTH0CPtCiwfS0EFZPdix8LoM8JkkbLid9WOUPoP3Jm8ZdT08sBwUL0VPKNrqTAJQN+mt5gIFX86M
lvHllP5OM0jVEeSR9tVz43ZBxR0OEqQMTYEXTpPw5tAiozkwD2jJ+OCR0bWviC+QdacQFhrKkgsC
XWlgtSRF8y3Izjr2jrRtifYRn4E4kf1VM2v/L58E+4MfZyG7pB7aUSwa/oFYi3hyYFDTqws7J7qr
+0Jcr1PF4GcYW8CPSIO7eZneu7VwMDPvbWyMHg7IUe3otLQqj5oOJ0J2fuVMpL5WDqk0HPr4iX5q
rLBFIzWz2vT9eB1vAH2exInzJARlJERMJ5SRs6uspEfpfdnLt4jMjnBk8fyEI48wioYHv0E/ozpK
bdmixHw53TxeOTFE9e4dk9n3HbRay9dWn1Dm8wvEaTQDinObGj8GYnU4YdMf2VITr5U5n4wdjOx2
B1724v/zj2OQU0s/lfZuVKsvFAtQdzHmS4maubAqnsyWV7adZtHC+zYjgcMFrIIA7GtEksx/iSyY
mp6S1vW4+1CA3suiFoMTpGGPOJaOUAdGxM/8p33ISK98/DrV46fEZwIvixJtoUiVeuwWmUMHgQyA
7vwpQ/hjlSj70riaSC4CJA1VQ+iNlT3SSjnzZZobjt0fAlmWAo1UEl5qlYayLuaczzMEWH5I+Toj
T8YY9frsVrwSIiYoq1W6j0hLCxzdXArtCDBvaoGp/DQSL3qdoFEiGw0SbZB5N6fmQTVlZzckUXSe
yKPbIU89Br+W0S2EjxPxb07q3i5qx16S65XOcFe1cKskdiPCKzODDXjFm+by/bZod+Lvg4abKuhs
VHq6Usbm8RiNcYD1/1a7tad5bWGQveWBBtbNAOQQGs7RbBE76QYAasIIE5P7A6jtLlyxk4ddatMG
YQ3Jo0Fjf4WwlShxa1sEVmsCGdMpBPvMJ1cW8Xn3NeRW3lj/yiSnE+xK1lT7QNb/4DNcmKZwQMOh
xjjr5Ccr+RdHX0UkbsfrOYgs8AhdO5mnKdWU3IIJOXpCZjXbVdI28hUCBdTWgt2emORWXhLYdmVc
XL1JQ86LyrNI/UzQfml9Qsy1NhYutwY6UVxrm7xm/x9zg9vtx2kjPtEJZWngh2Fmwn4HA2pVMj3d
UeWhbwrPJTiomSsyaEYVrXYEmWf6Ahi6uAT+5qRAcGlKrJ8BEoESczCwoe9UcubL9UMIIPkeGxys
zGjdTFnLXid5kpemFhbMzZ9Qk+pI1ZCf9wExZ/L2hNQa5R+rBdyV4awJd5PE9xZACWGrHZneN98s
kwl5oHsaaVYUGj0PxTYnf7JH0Ih/5t0iih7b9ksY3LGrKlAYud0ykYVT2bIcQEBw3LhPNhC7ewCa
INBuTxDNftnZMsQDAixEhl/rjsnGeS1WMlWL5KISHbId92lMoXWt2FafoxT4knFgiOBsMnBN4k11
TAxWei3rjCAgJjypb6Igmiwm5UAVk5hmZ7saB2M8R3g8ais1o2ELrUPTXegDC5M6fg4iUwz3AJCq
LL/UUAe5HzGh1u2+sy4GfxK7vJD6jfk2hONAOpRVJ6ZKpZQQqRLE/A+CHyfrX4mY3I4j6VMFea9v
spwEcUW5hO4UgoezZQKiUal+rVxvDRLflg3rEJ8tWBoD5lRtjT2y+U5HlOSf1KMB6X+3JeCQ4aD9
lPLznvjnw0xUY9qu20IkXBV2jFS+ZI/r8C4b6/vm4Yi5AO91S0Bomyi8UrhNWqxn31pb3rwh+r2O
Jq6Mec/1t7JuYrm4GPq5si5JpCzlJa1Avo9RhvkdgJG5ogx4LiVcilVsvMj+vrZycwIBAWh1v+8F
eMJl/mUrCboNMiT+d/Kf6k6bsLmk+L7ObOeAYbhrBHe2U1JUf8KRRq07eR8/uWwYblfhXdvNyMUT
Chjhi8D6iHVnjgkPENT5I+1zYbj0/vKwnO3bhaZCk4oJtHfUVp208tQ95pMa7COVWne7h6xJkfzV
EWQQvnz+Q4g68PZfhAgV5Ic6sTz549baB9zgHmN2qnNMAzWXxZfOmGLo9tAPGlW7EF0+jn4ZBEWA
S6Yvck7KRW4YWUf5aU6NFGbSzUvHciA8luxFgVt5FACPpMDp9VR7CYPb+aPfzm/Kkec9x6th3ANw
byP6b6ZQwLuHvnaTE06cQz6qenJPpiSyCEQPFTvzb6hSiIYYC71bIzPw0vMDyIn8khEycICsx+BV
Wjtzx4/Gy4M0PEXtsar/sF2UlHEi4znX0IDcISpNaSqm18ljipy+9HBF5dClfxhv3EY3vJLIRn4h
zEEylZzgCPlQH8u361t/lU0Ng1lBwHPFwsf56WSGaRtpkBnoGRJNBw30K3u0df3ICgDx2+j34oI/
VJ6CFm2VQl0NY/9WUd2CXFnidXJX3Rof9jdIr2NtyisPVID+2/BEbgtrZYljcOHaqQks2UabHbJx
8tSSNvqvWqG9MZ1MTB+9fo8/7BwHhC8VHpNmVYEV9zXWV27gZVaTARNQdEOdX4tj8fjtSmdllM25
gWXq7SSbJT8LFPFZA26/7lz61+TwJH6khZ6TLGqAmZpEODQVvVlk/Gnh1ZLRATppbsC4Ew8CEhKO
X4rxMIAcUwqPh35ruFSsANhktmqhr6x/0tYeUDOdSui5PSj90Onjx27QtsiH3Bymq4KeTVozyuM4
2yBLyu9TPvS4oIo2hrnsP89KXoFxe+UTUOsuMR1xh+ATgqTObDI3SNSvBR6jV8x71O2KdWdWi7QT
NzXZd9BqDtd1NX/2jnLKkay6T8SJhwGgk7dzAN5ddLJYv6YUz1t6MPqg+2xEeki69hYeiGUSDWzM
Q+r6CUr+xa5d/WInP2wxowpOHQEkTaGAciT7mEquGW3o5ANioQtRBswzymQIZ4iANC+ON4JSe0Ah
/2qpn7hMyyPeDsX+LpwCI3LwwC68caE999z8uIl6iX1AhAUBwFp1b3pioNmXVy0i3mvnDib9yb4a
P6/kcu3/qiaVFw==
`protect end_protected
