��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��л"��D���ȗ�{.�.�[�L"�I]j/G�1=��	�2`����!1�D�hB�Sǯy=0����o�B�_�!�F)�$���{b�����y�!.�+�2&�(�F�{��&��Z�AC��9�:lr�l��u>�/��[�z0T��E+��ΐ_����({�*�ؓTՎe&���������+Vj�����ζ�o&ߚ�(~�	,��zH�u�UiK�!��`]��e>ޤ�%�K�\1�{�<5�I摛���W��<���_�H��e��r�<��6y+�e�ٵ����ͨ�7�Y�r�v��ה�Y��Wd��ӡ��,��C����g�ċF�F���[,��~������|b��� ��P��H,���v.���J��%v�Ǚ�i�1Z���ժ�g~K�+���p b�*�l�`��.͟��%�?�9)r%`G�A��B���e1DG���#d����O�p�s�Q/�R��-扦K���Vg����7�w]Ҫ���3k�M󅀵����EF� �Q*Ǐ�@���+����/Iָ�- �r����1~l�,���i�	q/�=[Q�>��P�2�����3�фh{7�N���+�v�,����g\�RC�J##{��o�Oţ�V�ٝ!�8V>'#�վ�Vԧ�}�����Ͷ��Mm��s$y@M�[w���Bk�j�b�������S�*H��]nOuE�B#X`BS9O�f�?CYBr��A�-A�F�Bɘ��y�[�*����1�vhm�9�<;����2�hz��������?�>�5 _<i�fpF/���ʼXB�F���x`��9�"|��	��n@(` 	����,�zb����j�����O�R����A��vLB�4�� 0{Ն���nu������P�x�6Z�wT�7�������C�eQ�^�"���~[ZvjVdj52�gC�����#�I��C�h����\�R	F��&��z%SϦ�����:!�U9�_��t;sp�Rk��(�Q+�ԋ.˺��m�#��Z��$��>��>��ͬao�S��z�;��������d��5�޾��e���}9黖�[�x�>榳��C��k��Gtp��h��_���N�?�pA���u庵�ȔaK *ix"5Bi��2���A�ir�ht@+�js�����ȡ;��ݡ..��QJ-��8����ȒǞ�X"���GQ)>�(���Z8�٣�^n�jE*o��{k�U)�G��ܖ��A_� � X�J��G/��f\tG��[���K)���U�V����Å0/���E�(�t����$/�^EUgn�y������(�U��$�a��������<"����2t%I��Yzۍ�adtؕp��F��`�	x\c"���#ĸ��2�n�����,���ť�&`?1^B��r�%5���x@����7��( y��\�����D$�W�j�i%_���x��y0���yytˆ��|I�9k�U*XX�P��R���8���6�r�`DU+��o-�Hc��\�p��=��X�84������8��z�b����OY�{"
�"��*����Q6��S�z��F���$�6��d���� ��}���qSAcݢͳ�<�4��s��x�o��A�<��F�W��'���P�R�k��Ä!a�O��������+���[v�<q:���u�����c�� ��%V�o��!θܡ�;f��иt��׫�.��g�=�3py_ذ�L����3]���`:�i`�M� ���h��2�Mr��ږZ��KܭG�
��)�x ��,eMK��y�K_�e��gq1���b�,�rB�ݛɐ�ﻏ�iz�s�F�
kfRA�P������~�`t��yO��.*ea3-0םc�����i?"�4�s\��'�}��}���<f�H.k�&œ���K"�V_����c�����׳�%��Ȝ�y�����c��*,�r�L] v=REJ����t�R'k��hv�&ެ�א�/�ݮ��=��c�'���
�4��p�Ud�������z{ ��Ŏ(U�9�L��gς1�k$"�nb7��9Ҡ���m���S�-