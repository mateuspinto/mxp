`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
dJuHBZgGGvExrGHyqxUwqx3X61EOOyYQcfx9Bq2q15c4xYei/yN45y6YpCpbIQIN7IDQTD48sTz6
WvooSAt9RgpDyMU0Djc3ztkCTLrZoHHzfhdY9xm4gnQVWU7XuvP+tgJpune6GCsHS5NHA95rcZFQ
vP7tp3ENGFbIue24+1NxbkD+6YysM+kU67s78doqb59BRASBK7b0o69jiOHmR7XLupLDFt+tEtB1
SKHAnpd+sUlzmbGKRO/7PANBlO6HZHSGJLoMn7Z3BtHYAnb6/p0nFAm79ZF51Q/whAc7Mu1csYi/
ozdvLGc5LNzKUgMf+eQ/ekTGYG6Ea/zIn1akTw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="PiMsLZLwx4/XWaxbyeARhGTaSPVEvXzrZbHiv48GTVo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2160)
`protect data_block
WUvOCcdPwIQ4QBPbFAsGZsX7pjaQYxDdvuMnOWO5ZyvFPjQDslFShfuPEERnwR1EmNXsgJw06oss
utWzBslj3Vctyh2fteW/kO6bJRjXM7IYcQ8Y+YOk7v6fRzDv60p9RhjWqr1V3iZANsDQwkP+7BvO
07kiiLMHWVUjOp4FVqe3v5PcBrUcjipiJaK0tkdQftO5wPT3tyVgKnLROWgk0Mtnqy175pCbUYoF
I1xx5ZLMwMzsfvtx7W5vV8gGfooIN81Xy//B9PCwM/hrN2GX3HMslJC6uRTd/Qs1jA+ypuGOxJqJ
5bYxWefGoqA025DdTw61DnWZ+ztRyl6fAGh6Q4yoxFq+8K4Q/Yy+ObBd9Waodm50vc8DUCy6SeWX
OIRPWLNVujdT0mwfg9b4na66ghZviEh6BYBwxCzTQIol4A7KGkHSA0rdUxo2YSlHkX+yLnvFjNHx
f9Svntp3BLClxLlsHPeTBa37qnnKTzxHW44iBmechJH5HnRtrfoihxz7lsVohBDj7B1I0RXvELtJ
YfsQ7Wv/uYfsm7EDoQLO/Lupu0WKHOnjylXPIYjUQMcW/wEuRi7rewVzpUR7wweEC+g5bwzdZKn3
2698BIgPJ9+JdXm65Jjo3ZfGc7K2ET6OhpEAQOSnWnq85375qHxtk2/T9J7nBgkbumesYSs/O/FQ
CgzpyhpGs05n9psV8yLQiXTFoZtPcbVQZUhg+LN75pJiWhDvxebnY5J2z/GkYtV4ykrdx+SauO3l
mhjKXj0Wb9hyCjjlHF8Eq5nUw15gSLNWEF5lAocv2S1BLGKi5131jxt4WxeTtaJPORi853/6Cr8y
pipdSwXbAFO952Od2sBX4MgEIBjmyQ6UjPjp9bfE1X7dESvmJrmfvr7m7YFMLPbx5wZVl/jRkzMj
kOlZKWSrPiqZ371TdF1ZLAIpFUOj9dXdTpvYTasPV5T7480luNEZoqc9CQnuRUUj5Z5CcEr7ZUbP
ELATqxVTnxapPvplZCnNDC83IOblRGx5TmPrkvJSq2Jd3J5b8cyjxxjFtoBDUUzsrDc3kZ66Jrhf
3IemrzRYyp+u1EIAr5Ri79tBhrktuCZtGP4ZB0ZSwCMZrC2ymrFGbR4EPhSW8eSci30+bPb1rnck
2FS8PdDXsyYgey2dr1DCIwYFIDznYU/HXx5ekJwtpItF/K95iDWeu3TkSnjTjQHonwxc35PdRKl2
8hG4qk2NG99OxKAeNsJYd0mn9JNzyjDb0/UtVB/hu8lQedIRwHbXEurdCoXhxr8HUOFQRhwd3bJf
GYL42f4L4PEVzpJMQL3hXMTn/ZyfI3XGsM+W7aQvW4llTmfOBkTG2Rsr6z53Tdj56DizIiSy5NRG
7xrBazG/A4GfMcrJ57inUjkI/mgoz8nQHOi+i1BqbuNH4pej5/5jzBLuOW6yG1P3bo+4zNrij6aM
TshaiWouNTLZr+SRsVqkKLo+5/DQbfKbFVwkMYlkFh90DVx/NbjeZ5ShAdS+erWS8saGGLjfBsAl
UJhKnpAo5H7BmzAinx9pYASnFiZMKmm8PQYrVOIoweLl+eWLaYBtNgFkESM2efVWAYsusqu5UjE4
TpD+FkgRtehmPIu8a0uuSRE6h2muRJhCUpWfdyCzCwPyrRQPt9TlepoV8F4ny/Fya1hkH6Hd/f3V
Eb7vODtOwEhUgvdaONLa5elVCTTaJXeTVW2uI5O0lBYowum5b/X6v0clL4429SyXjv+f4wAEOCiM
PmBoAEZ+SzZFFPJyAS34OHK3eK48c1Ot/ReCFT0xIBmuRGOZakiuGvviLoGp/2tOmNpuGapwVf/X
2KVBM96ATt8Pm1UROHGzVAaAQHKW1LHpwAWFBKIYbLxxYKJf3JReE+xifNsFRw31kixieadlnC/k
PAfGswxei+57ZrcnEoPauGnj2E2PwsCWPvlxu/4Va/lJHFGe93c5/qqKurla1YVd52yczVaGNgjq
sHpOfXjgGT9zY4o4liGK7qaAO3u5rvFQdPo7SPh14ToVDVnJab2Ui8Ogo0lz454pQmJle7/PVq6n
T0D+eyFeVD/kmgXCzXI/A6yt9RQkUdWYgBgy1FkyURHOiR5oi3lZ189p5rpj41es2pJE7CzDZtQU
coyKATa4iaFIElxAaaYT/0XcTgDouGjoDfwjpPQWO0cXKZIPKdDag0Ly/UrUO4e8O8/Rm06nwIsW
/DEPk6we6ICW1dLHS5AFj5Sq7JfOPDk5xR8q7wXHtZLdqd5RxvVRTv3kXAnEhZfdBWuvtJ6SG2rU
i9mogUR6DV698nwpLndCw3zdJGjxIZoFS6CwdKFbQZgrLBTKiSnl5tuzgSCKxjsoeaGOKiSuf68v
vq5bmLLUyRrItP/Lvbvpi6k53YO4RYi9MAGAM788G71Fij/1UvTa+ACMhX49GXk3WNuI54bWPRrI
76kfiiIYtz6YttgUsHceEFUoLvoqc/m1CU0UvMF2DR5Z240wAeZ9IQlxsMCZWqJ/Bm3OmOiAX/4U
N4FEkXBBo8CQWaGqGOQB4kJhB7699l4H9DBbt5+DyD/h1elvhyESRC9PQ0O5zmN8DfzEnmFc4E0y
o7b5PzsQcXo0oXHz6VGaE6Yn5BD6pxCB7303ZJ5aBgCmdHXemeMEzW0RE9Ct+7vnYevELY/6A58e
Fj5BVZCDDnxQDXcHeHP0qR0qUP17efN2f4nFcxP7tbuZU2/Fdc4YPdGqFjITDNmgHbGq7HR60Yr1
6e5EgHNkAHLZiDr5cs6JxPUIFdu825LVxehW0mgr6EIPgWgVNgnIgUWnmPmWvdvE2Ta16Ad1ZRRk
ju+s+eYuiMXu/g0hMDXRvBki/PglnHvDp4BQwcsd6iN/bQJrBJCUP8c0QeE/x1vZm3jE
`protect end_protected
