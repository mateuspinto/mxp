`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10640)
`protect data_block
+B209a/ANTO5nVEye4bSopE2xpvLvIjbp2DDbJx0gVAUPT7w/fbAHcESH3buWL8PJdcWvIA1TBUW
NR1GrcC5AuLBLPbyBZP0hjZ46vCRLe6c4GlMkxijxc2unT3pE7FBjdsNGi3GPcJDPbbKgj+ImBil
1T18sYvVmXXJnPZtTS6edax8FGWJIPAwAs/QHe7P1CqXKm1u594XqhRZ2ZQxVNDIXdS9eiVz6SBd
98h4ak//0gl4YuYGkw/Z4Rd6bzlPcFZRpBgtz7Wh0yK0bIi7c9WwHY1yj+rmkPtTy8QDqFWuD5S8
2nZA2dR9rkzAjb+PRXjwPh9V2Fk0AI7XKTe24t0xXI9LgiLJnkntGw3YwXyixo27+25SB3QvdVke
bjq1vZJ4Sjkz1ua+3SqxlvEsTR4HdA1bJ0T5ZTvC0a22vB+3Wkt+VdPnd8WALBRZ1PYBrCN3pIrb
MyQF96ptS1Tqxm8xiwBZzMAC3sWWs4vYDwWMuLppc2LQfuopPPGvsVjA0dx+B0VWD1mj/SIYQomI
YkYw3SQc+MYJbnWNnQZHbey4h7Td5Bo44jgTdasz0Wz8yIgxioRr+g3Lj++xQiHt0iz9EG+nYS2h
dsB/cmDh0tM/5FlRMr2Fi8XGAhw9EOqYGt2jlenu1HPp455dvPYDmVX5QJbkhU9ISASitL9ZuQsq
6XVjs7lapq8KwaAJOtRN+ONNjZsGFgddSX2dLvgjorVR1rq3i9u5d93K27uY1VXs4vnYjo/BenlW
x7MJZDJ9QukEcE7eIv8Qk7LSoyls7cOwrZS04CHrysD1AD3QFZgonW90wSNEoMDHvb/g1PiteqdG
KBmAvrCj/H/1CDTM93rbD5jvGHQNoCbXhSRHbkkAkBW2H93bvRKEwXQCdg8yN99bwY0NW9EeFRQX
nO+CFW14skwhbmBDb/p/twqoNt/waC+CFlbI3aFeFxPILDmyRG/mdv0/mBWZXjmBxRFAqfbY9oWz
OGxlpGu1/eJKcsMQPkTApVGM0TC+cLcj99RGsyhtyn2jdOWsHnfmlxTokDqnU4DDbFHxBaaexgw4
tNbUF8rMU2seLhbgKDfj1dBqh3aFI8g8xvQEmjjCmuyIbHrnb0sJ/g4/04U8CeHUPo7sZnBWHGPB
U1aWwvnW1fecpsXUQRmy0uLicCTMOnzPV6LgNxuTnFn0BChFszgF+AFdqV6pJQuxWZqrXPmsVuk8
TR3V7uj/dmGKaDBUtiiC6FxWMGvKMJhYlQ3M90WlEKmjvgrGd/ouDNCVWZBs05BjhhATkiiT2sN+
FODcv+xx+P0TgaM6MPkhBv53yibpUg7i+Edp6df1dyS491h+wljhcduFE1IbIkvA3YImzDif9tG6
0gJi82FSWbqigzV6olQCW1NcpP0kx5kQv1uTnomU+K/gUJVXPrAYAZBheu04JapgZZORBMR2NDeS
A76Aafkr4hfAWokWJCMxFvDCnLal0Q6Qo2jzONN6F7tCgbeKcNY9P/ltmveWmUrSoQfPGiYVAuS7
WxkZkjglgCjzCWTmhuQSXPofH0aMIVu6MDfNauqFK7gIQuVyNL39JPbXv0sw9cOMsXcJPzl118EB
3v2bOe27CHDltO+LnpIpQs+kSOpl7HusWmoJhSIWpc1TkebtE7qFImdHMaZaJtuDII4+8P+DwhGF
8CmSBrhkwvVAxuIzSeWbac4ZIOL99QV0Yk7/013Vim+LtU4AqOWmcq/MGgwdC4SyrQch23haWtu5
DxTIC5N8P4e7BWkjOqnc/XB91hDmgt1yQQVpDOi/9JlMzYNqm2MFBRx2Y2K9AaIXJia9SXpjUabE
PetTVS2Lv79Ov242Tvlvua1D5QNSPIcBCb7n/SB0ruvaBNEhMR3LavNh1M+sfW0Gv6Iy8KhPdPZG
3RORBCPTa5n2nWwQLedXH4feF1XAjQOa+an1xjkImF/FKtUsB7MkDKoH14EsuzfTUX2GHqfjGfwn
sdXD1sAaCvdLfXkgd0BKHc8zWXJyzu1x5DbmZLiKwaZLZ61YIuyvRelL1USJieXnFqhlCwdiihYJ
03TcU0FZbeSDq/MR8cYvL6+l8Jwmhu5Z5US66inN6u7OmI+Qo6zV4xv+YMwL/Iy+d2CCL6K/cLJF
NfS5WHBr4KOUx73vHL2RiyRhNfjyrGSNoaVukOBl2fmBucYlNbQwB322mqSQUeFbVUlzBjMgm7pq
vzc8Vj6JthhNdgy0GQ3eO/thLXTb+0hsF7LRvP6fDN+GcLdTDU54PceFK53J840KKbQGpNpsScWc
KOfq4sESygSQbTJmC1uTf+MH4znHtwkxZzy9gR9Wlcc9nF+SA7V4cKfqeHrvGVoQAv5Q2QAdbNXd
qTLtiMoqsB7NMSY5Q90AWmvzeuqdmwgPz9dMZNkzf3Ynxw1U5i3nxJ+pkXtUK+c1igNDAAzNkAe7
Y6ITysEbm3rnpFUEteITDkv6+dsBjZK5uNkUZogQQJ2SuxgwPyCCoceUObShX9OTf542HMidSMOq
85qO/0c+sRnH0bQak8m3rZS/E2XMlgyL+xL4vjRRNQICc89K8LpRBxe4n/8SjMBRMFnkpgdUWk7q
KcSC6BqqrRWMIUdhRIymj8/LSBCCmwDqP6Ym52j8QOlTtTUKSxV0u/+mdTYazUj1gIqWr9On4vRL
NIgIJp2QjukVyb2d5CdCRAM6hebg6dcyX/ZB17mz7IWgphfyRv+NkRI+jM6MLAmAH0VQftk3QJwv
NwRDEqb9Ci9dUNIncA16Hj0gqffv+17kWohpiAegqe4AKdZStC6cJPstZQPGKYIRsS95+BK/HgIj
jpf/jfXwN7+aN2I/4Yf/Mf2k30zJFsWFB4xdqt1+0iZ8XB2cRf9Crgen4H6K8n9qsCVe3lRAXVsh
QoxbnWPsT3H3Z1OXLKxdFyH3f6FkhBcJvWwINVVsHv369bE1Dn4tAvkiKG/3BvXCSOLEAE9J+FnW
E0z7fB/rcMiYsPOcHC5qXehqcVfjIriTGP3XA36VwDvdPQvMlyaNMYJVBGWVSbpv7gaJ0/gKG4ND
I089bSqO4YmexkSGS8yE09kb2osMN6nqSL5Yh7ZQENplrcYuT6HxuMke4SkERZ/cxho4kPXqPdmy
gAd5vt4ZJr9SQFWdrV1PtZD+E+02Zo4ito7uVix2vF3Vdw4RwRH5xxENMMfjI4T4GI75V/9P2yyL
YOCCu0OJffD6NILRLtwreMP1SqRt/UDOqGdMS90ocuauP0LOa5buMgMtjQzv+VRYv2aUxVgK1mmY
hNnhZZmIPWJ/7jEyxH4CU2qQmyyvY4/CknCA+IDkFB+HiZPf+rVR66VHEUuYZMra0uH6FDmk9h4y
Mx75E60pe0InZIosV+cxpB21667xvtkb2kyvs7cdPonFZVu1aV1KQJxHgZit5/jOiIiuq6wE0De4
RplpUoovd+vqQP/49bNCiu3sHQsVz1VWHMRlSMF+RuBNE8siawMgNsfgkAPnFQ8CyuSUQCcHnBda
lIceYwWscO4GzeEhG7e3GAWOQ5AE4dls4XgaS+kNSKpJCXRTjDGkSDsjD66sdd9Z7fqM0USu/cjA
Kv2WcsZSGunWSMMdJPuqI0IzYpc/FbdZ9Hyim0jB3FPq/WJWingwB5kJxq0DuKSbViToHB58unNH
DCSm5zzZrROe2XdpBZn6KdDLmpyuR2ocTzHhRoMklrC/XEgLi5FY4vQOubUVGjK5JbHVRRJzmSOn
jmMJLh6jMLwSLNb9H2ictHzilOVNY9Oi7XvdUym9PUe57C9HMnV3FxJOWjfAYXwZ5EluMAHP2/8A
qpJL6xH6dCx9dNsyVGE+KoBg+RS+cL34ccYlyOPW8MTO7kViY3iiUgAcQ/3WeDohEul8BkNpaSNF
xYiyf+fv6UCDVFh+0/4x9iH+ejknE08RcKnv/aTAg9RGzXetLJRTK8woaJ3OXOpLAdmfwVzplfmL
8hMOa2HNNv9yRsFDwXOhbH7Hv/XDmIwPgSD8StwQldGzINpLj9lS6oOjPYFhOoOyFvRlv8sRSyL0
SA7jlj4YYDUVxPhP0UG9M6jufjncAho9JR8z0B/OlL/o58tgQLWZZ72rJ3PKRwPB1tK90H9G3GDo
76RFw8uuGaN8U5i5YnDeeVDU3cF5tck1GL7sPT2ODOMUceSFfgUZ0GsGHy5JEJuDHnZhCm/pDhCX
nynsgWjwlyV66QVKXTiQDGrUKpSxSpIfDyVlbcUDOtE0vmdSTDzi8ancfb2i8Y5nymSueMayj2Yp
lwLYoMezK/ksOHCttZ2rdsv3ax//MbWd58YLm398VPTGZKARjAOBEfas0PopKimOgpPLSGDATRYK
O7JTTlaTQsuIJCEp2qhpFcJWrNFDKRN8C3mZELRgF9hIxCye/YOgDqzawHnVe9o1KYJgqU+uo6YO
H9ZrX5eOE8WOubqSQugBoO6YsRKoAYXTO+ABDoO3OGyazoovhY94Y0MCK6tUTjo2wOvkVj3Be9zo
8oHiSUQn65u2TMxCZIf6zjZdX0lmDEGra7PqqycVE08KtxpTxIUgv0zDs4F4VBlGu4lTLsnUlITG
/37cISnnJgcG/w/HE7HNUI0WPQsNC7VBSBRer7+BFMnY4jNOPdsx+ngHd1D3I+Cgvf9ozu8Wh7C5
rvz+HjI/oV9RKa61vAtN3O80eXSYWF7M7NLqcErAdbvDISpd042K5J4DgzO8j6+EPAJPQzjWRfrz
S9nQ6IX2PwB5v8MYt09Outjh1FkzrKBPS8BVJI6Tywfeu9pS+Lgyflzdcm6/NlYvkRO8DupDPQRz
+l1lYUQySLIA9XUpxFQfq7j1gSC/dB96YhAOsVIrY2q2OBML0id0afYVNYPez5BO9BznqPjh7rRo
vlE0urS6ysicQFepeRM7NQ1e8oAAJZxzh71R3gMof/Q84GmmMt8+YAc7bAQUbxi1fVs7A3WHDfc9
ud80OuqnSbwrjWrYqSe5QlTfg+qyG2ENfADL4sgZYJj08wYureuakK3jq3yEpl0PQHPfFNZAKd2V
vHqiBO2RFHZMYv83k5bjixx4sa7mSi3bH/0EL32VBk+MvmKb5NWBSCO392etOZ9El0Y1jXjjdhWO
8qTTqO5sAM/yJQhJz8dJQYI82bA0ge+D5G1IxSDOX5xZfriZRUp4qrOp/hz8w6xXheaFtrdKEJsJ
c5LVATgapP3t5Ovn+nODKnNijbO3egSAi7moB1BVXd+9eVpXJlKJuXuMLuakputl/zvyRZkxuvB1
A9QQ0iGr0dO5efTrFn8WDWQpo29PZA7m/xAwJuUBIapRDgwqXr+2+/YCJv+znmaA2F9/fD/I21nL
X0Fi2Lfec00ByyNVPWJhoZxbHvybrvbw1+Q20qaiTa3YR+KThdHymMHpGAItXQrfR510CS1/vRes
LoXMwjHY4JCqSmkSG+WPadC94BNBOhPGlXrM6/8oJE56bpUBeyD6Q/Oov+ozmfLepQkXeRX1E0iH
527ROQjYhST0zsqxQ9PLCX1w8/eynWLvcg/PEMD44f/IE/y5/W7zDLcT/p4oq4Q0TFRr2HR7oJlC
PF7S+G2fnaEBYHbpLjsONnixDDqcIrlL4LLIbGb8aXoMPy0KMKfdRjMYoWyz7mn0n6JV0PJgrbFR
koIBLjA5o/Q0/qzpe92D5m0YY6DVCudER8z0zYCu7Fj7Pi36PUKDI5vINIrh0GFjfuOaA9ELUINH
knc08acU2Ta4SSq2Ud+NBc9bm7Rr2gtgQzRxnzVLOU4OnwJ0eB7cSXntkM6EhnrFcqEcs97L8mFc
ch89qzQF1VQvLb8pIYnsRKu22kIDwiuo9lLy7NSGi5LFhl4n8SZIBId07rFizwHqPjhdZL05HVsQ
xpd1uE0qct72kOUyOJweIITnGf3ZLnmxKR1eTl8PSVCVol+56YPB1Q5nhb6ov5jI2lne5vyeTkQL
Bi9tGfEDnquyJL4lmQQqOP2XpYzJltx2bUjTYTiYUtQWsYXDeXJkggaxgiVXVKwobJTvQxIhllzj
qG87aTfRzXEhM6ihvJ0fbJgi0zXfWxheIc7Hos4RcT+8hEsH2a0SVIv/JhZ+dLC5vqHsu0fAuNMR
VoMEg4pmMk1VYYZk7lfyID8sKxvvr3YmlTkaqQlpRwun07hWK99JmFTEGY3ReQgLrbD37W1BIyM8
teY+n2cKe83Cc8qEhBosuMdIagXPghfg2rB3zBRBFkxRP4lhYPh+YQNQEZEhztV8w5AtBUF9NpUK
QCZKG4NwXMk8i+3BXnaP464D1axErnbQTu8vXRr6+ensnkBDfylrta8knHtSVVB087Ohhl9+MPgK
m6cfDRRCQoAVxqwMSW6gWL+vtrJQJ4Q41qmNXqJbDMqClfLTGATsQge0SauyhuixvY5C1PNU73uE
7cFYDYb5f70HheOdOMVHgqQBSLkEw02ZCGphdAMw0fBbDi9H3U6H/XCFI2rzPIw0snp82cLMCGZu
D7k6yImSSL8dIboQ5T14r1lzzlXmeiP4lPsxnf1TUUo3tvNnOGBCOWgayki1EvWDp1ZKNxajQOhJ
o4QeO6UckIjCwPP8WAMpo+w/ygh/P2VqwgKU6I26P5NqQkF5NJI92zIipNYqPTnfwegdTgLCzaaX
vOp70o+40B3FaTGshfGyE7M145G1/XodzsIG+8EnxVtG4Lh+iRJqQvahEF6DttKZRzfHBtUiY4sA
LEMu4bc/HZ+lPEATTGdogkD4ng7whMlJFnubN0zikg9pFmzTBgB4wlun4Mgqwd4372adE/8r1ldi
H2F1+4iYOvjcqKic3gLdjY6cv3dOGHWYX/3cfzE1O+og+ccCO7IX8jLk2H8+qHIPZZISY9MXUZw6
5qQH+ieS+4mqop/wNnvyLKaUM91YvBYMIz4r6I2qc/2/Ztx5mjKlm8+XOHy0bCvqWvb9JAM5J1Ul
dKwAzYLw/kv3gVX9mTzKJCi3w+Sxy1nuxBL/VaHU40xv8eRvHtXKIZX6rADwxbmA9Ig+LmMS4uyi
GPGrvxrFIaCFaeP74SyKCNqjIRTjNyCpkJ2/9aJRFTBGhSVuluuyt9B8c3CNKZxZ+u7TgzFhgcZB
M3IsyDJ64S/dVKsJBkhU7f1HdhtSTzWzYKYuaHk+qGlKCffgccMYgAl6hH6Fq8aR9MbzofnY3/FW
xWCp/6TeLS3wjsm11ZEOpEmVD2Ub5q9gTjUrT5kEF7ob/kWNFFZ3uhDvqCZrvPXBNxWrgn3ykXP5
rnLChuhSXSl9gApyxnEey8d+XjTp58IXdmpLDZ9eW3pkAQiNza2PvJ6YJa3kx45UfDojOA1ypyoc
9i0Ynu0/4pB51q2g4JiUeHJvHfM3jdiug1gaHnWfFlbfxDjxhMmBf110Z+uYuyZOpgbZzZ7aZGT+
UcVbzvjn+zLLFTq/BchAgUTVSM0rA+HKAAGMOJYHQ/5xJGSLlElM8zkuMoBYvsctEGqQunXegwpB
brvEvk+3o3JuaaQz+sH464Xe+rp+vjQCv8dzBEkJxMpHXkS4M51qnuBd2LDlwj1ntwwprkkOoXrI
b8FdVzYzXGp3GQunHRjO7zrE6wTPaLqfqmVSFrd0uyCqrLMkSdlWkD9ytowPTjWEo9GCMuZ69cHt
rxJKBEt0Dl7g1IPFSrvmZMi9ZGWRXeVIxSHOVkxFxXn++/qErWaO66IMvxXFoxKgvIPOOV6S0n4R
kyQwZG0pWPsoQdwfxHessPdEFNcOg18JF2h7frU8lIkejqmLMBtk2C5Q3rjfANk8YG5foI/ulBT4
yQWjEbeJxuOBQx52WBZp7Aey2D9xbNwjxhnognjeb//a9CGYOAJre6uNoKyF9AIzFd6rekD30WQN
MTKZaHxeUxHLpulAE5P0zdsyht8PoI7RrPzL9vunTcNMDAAQlD37cNanaYJRObJCLd8A6a28GN8d
Dpr5UXUVyw+y6sH0Oqv8r3DGzrlxkWoXvI/8I2i4iqpKpdoOD6JxvA3xs5wFShtc3NDoYgRgIslN
3n3Vg2BEXnB5HRqkbuxvAPztI/DnIIiioBmnad/SSM5IifNTcDz3djaEQlMNGUE3GeVyU6ggLyDd
yDMRgs0GZOFzIEAzsM6eSnJhDnSNWdoWW7e1R6xHlHRED0p/1+ThG/+lGNm+zt1r9ZNQCzVEn0GZ
e/Wu4BLCMuZqcFkSSxxdp9Sn4UngUhlsC5dd1/AQeN/DLUBVhVKY9rpsEWi1y8BFSsRhnT6yZk1Q
qeSAF23I3pA+rCR7CkKf/0FmvaYfy4SUOdR2if376+cKpU6Obcw0/VDSeBsb42vgF34a0zSU8cAt
l818zeaZ420dthM8ZyVkLjIJIhLE1Grfb1ttjxm4npW1jgnhay75TukQRGlJQJ50mvQd6ub1W+G7
4YcGxwtHtz7bH7ebCy9FyHY7eLHGx+MUqg0n1Lf3oe5vEfYzvIB4QajH9eQsESv71jlvM+4A/Pyz
5Ej/v4W6zdUEl1qaHysVyCakC8Wp0Y1Ot4hXfWCCpAtdgNLTD4hGxX2ZYHrh6OzLHSg+nilzMm6E
DgRVq+5PbU6EqywGxIH1Wm/jfCM6CtAoTzi9rjiMq3t5YZfvMc5RPk3EU5x90XxOSqchg8UOdzCA
OUF1e1CGaMs5kwEsKWmW1O3uVmgGNnkAL2EEAkhUU8XuCS9ozUGKl+kZq8m0G0mVXW1xKJ4ZHDIN
kQVluE1lOEsjgaZDi+8aajPM7eCYuYizcL0FGkQWcVdepG7unwtGij3RWZszITk/R2bwxymcF6ja
YuwB6zp0BRBGLAezqAJmNaGlgAMQVcXxLQ8RV/wegxu9kxPj3yUxyiHRJQrkUEs+zRPTl0GI88Nj
V2ErfH80itfSfe6iANNNWt5Oqxhoa836wy2OfQfJQVNB4K8WArTrn5UlQ8L0nOuUaG5UeIJUPBhF
koxIfG8NtXg9epsaicKAFStyRkeIANsgptuuOw/XaHmTEiE2h0kfbTuWCUF/HcGLIllSmbZ6JfEn
XPq3ZXyVvEdUaSawefgxGnKJ74Ep2m+iCtlJ9nlptm6RNYHLcWihxO46MSRnhsPGLbYZIVsIuYMm
spwNKr5WXZBkNFI+K5y1Cb8P1WDd9dDtplmZ7nhCmJiEXVz+jDmD5NXZKuLQFzxG6YChhWWIBaQg
PJ617lFgxfYYJ9rDGQ5j4DZ7RU/U/Rr5Sq/78/utbHqNVY6+dj7q5MhksVB3c7NQeEIJMqiMZKDD
lb3qRaymF3M9xBGdBmOryp0mGOkxdXN4TLc0lp/EwYaOMiETouwBUnn5NjoOsaR82gb9Wq9N6nWN
PoMy+C5mObmnDfTIwhIyAd9EzLrTJEk1v+Z+3KIQfXjWCtcNKMbes4P1bHJbzv/yFfgt4TVBXqmU
kuizHS0Rn/GBec2u+I69UHsfdnaS+4ce1/ke0Zln4Nb6SoGfAb9VlZUNcoEF9RVSvhQSXVS7NyaE
rLR1oR8HCkD1ShpVE4WbJwW+qbr4InSiTg+CamecHdYpr2N5CslHdz5D/JlqH9z8zh/0BTkhfWS5
PsPiO0BbWy6dHEc5EXZnkycZdvjLSB79MAdLxuKxIEXwQevrC27EsuHtSSIEa3vmwW+09z2lwJ5h
YnSlP9EApBSeneP6gHAoUJaz/nk0m8NYwM+P/6HhE5Le3Ar8lpkjOQ9OD15cy8YBih3UNcnu/L9F
viCKSfAF6XieXJYnN3XMbYXGFxVIfOaJK71e/HUfhn4Uz+BKorKc/M/sRh+JfAyX7nGtrPiuf4wV
m4knvLEBY8xBgN7IDKVYbEzv5LYNcQCaGuQgh5yecoDFMKnLZ9by21g855hNSrjjtDfvkTItSpZu
2NiIzXF9LVX35fVDDeN4xg4MriwYOr2S5Z/EnCuxdRFAYYwSRZlO18+OesWAv3iAaqxSP2yfskfp
mp0O0Kv4J7/uyzbQjJtm40zl7dX6eHscbgjN7tCd7RN8mYBYxRzt4App5NCfdR75McAGKtyg4cza
tD+5CF/GH2VUcNd46nx2U05g7IAH6ZeSMWExB6a0r7DDV5535bUsKZoHf8olMkCs54UUygITxt6O
sz1XJKLk9VHf4Uke0ThD4r2uRNQvetLoTGeOXhswE8TKZExDy9UbeI9qf9QaAtjMxwek0Ae9EYc0
eEP+CWrz1hnWJ/FhoAf6d3k1BOeteR84z/HMmo5H0z8ZCvz/EN+QVOk9u43DCzJoW+rjQz3hPcG5
QpbVCmj5wbz/nx216jbQYX4nwozycqpg/GXktoNu5fNvZuv1OkBBiMzOBDGgejrO8q1+3y9iD+N4
n69qmTFHhqm1QX7Ay+ZIZD0Idvz1LMEdyNygliCQa7mAcSYu13lLkv9WrtqJMaNQ2UHOR/Da665O
BGRJSR4IXgGXlLSL8h1HDhg74jK4u2dwZz0endm748YhdTw/CxDPNCQbiiDgnR2tLpplbjbrZcwW
tOzBqMgDwmvZV+GSA+Zsu4Y+ESw8Bz2DTq+GFC06DnVKQNut/JfDRor2wzF61QgagSRO2vNYoM1q
zN6TMd1RvifpGcGjSYHNA0PoVZi2MQClcVFniHJrn523FQ2wpG2ksLHp6/RGgGhy0hUdm9y+Lh7Q
YrX2zmAkgBKnL+s3M/Cmq2JDyOGgGz65VkDp6AqBW7Epj1IPDqBPK9qbzs/cycfvjhPMEiEOGdro
jBz/TXj+I22jvA32XU44rfoiDeA0Hg5oc6Cbu4EXN4YfAn9dYalURMbF8FgSO4W7sKgmPh9Yo5ML
H68ublxOHwFZbvaGx8YsC4JLjeEIZx2lb3uG3j7wxsWqcHivY0maBHQeulGDZ3ccVsTNldXfjKaa
vFqXnyowABGj9wfui3ifErLz9gvk9CsRCrZ+3H9TXAHWJGyowbsQSc6GKw4XSvdAWjIXpSeXSkbR
3dwTCTUoki3XayaReLAgPRSzIKkY82T5Kv0FGooMxafq58hmhBgZ9dt1eJr8t7HRxrRymxRW22K9
MraTu8JjoMYK9RxCJox7hKDgPX127EW4q5XniKNQx3KX8WTK8m5ztGNvEx8LupU7y7b81wq+lG/D
p2LouFkfBRsEFzYw9nrJUuJWOmAcZyhQ0WRgqhA946HNGTmIZg4pg9KcBQOKqpFQD4Mzxa3G4CLh
/I0LJG2DUiC8hvCJsRfegsfKD+A1TkrZuRVmZezosIj5AVZApSe7lwpH06MhADng1ulGeSS6E1GL
DpMY19NdFLcFAp/KEUPsMOwe2zynxl6fI6Hw/cHuJiqVD3oIR6GvZ9z3i8nhb6QOEQgHiLVwj5Wm
khV19DoWtW6CXEAemQeZfAkre8T/+4V2WYcusVYDUEQOva1Tj6zf0VzsqnEk93veeB/wrEX6cL3J
tss0PMvndf+SA4aO18xa6TeEEtpPA7QgyktbDS5DqAafIq7RISvSFEbplVhS4nUCYC/FIKNw1iGC
LWp/usNZJTL1IktlDH6+608uJRLqtZv7I2nmMwpaQCKV5/VDOxpqplxbRDp8e/+pVHe3euRHTn3p
XEwrfDlmBiMx52zFo0RCOqgk/DKdZZp0Dn1f6yGGTXxGp0hPmwNWfejjnvTwHviECYR3x75YBnDl
77fUpTuvOB6ugCcx9VHSuHtYKCo2Uaf/QsMx5U5+j3/eOQJY6EJEPKwgY3TdcgHYOufaDYWXkAnA
kotDUN/4DmO4Wru+JVURv1w+/V1fVAqUM20hSOBq1dmZXHW8+H8X3mdl1fCeIFPY6ChMhqq/Pm2J
21ACoRcb8fvpXT8FTg9Zh47xZiBAADUhAJ3AOE6YkOgGgYfPil1suUPNthCxRWC7u4TsClpaAeVT
LFGxWl1hIH1hCD2xzKNBgXJ0dwNDW0Gq08U2iPsLrw7UGXBSTJwh/9w6FWQpcbJkPa9G9nx/f2Zb
ZrkIPOt5izFtnyu96Wk+DxvfhkUaMZyLWHyjM3bv7PesDf3D51GgRwGMWt4UGF0BPht5uuf/WkMA
1El7zt0BJWiLZqflUx3mCIMXB0zue0Lt0XwLGPEJeQcrNMdUojUXuS6OPKLTp2dhdKjlwIqdmg4t
S1D2Fqylgjv2Fn1UcaoYyyNnxt3VA3DJfPfzHylC1TwTq3VzotWonIdlqVSumiFEz6nMoM83H/q8
D45uWG62YqiF/acvsU7q4suZdvKVCTAHvl9n+ArnZjBayb+cXxQg1mI0R+QRXywrQ8fPKUCqypxZ
7OMutGgha1GrV33yuDO4kVOSFZqVTnpzMiYk3xAJIzbibgvM9TZHhsBYPNKZMxhmsrH/ncrILn3E
jMV5BRUUJ42IhJ33DwaY3+MqJoSetA9xOzSyKL6Ob1SRjr3u2kNOLbTjKr61IFj2r37s1mZPiOeg
JP1U8bwm7WOCbaRnwMY6pPkh5oPrNTn1UoJOLA0eqy55mYoTjek28afamL9Izw1lNyXaDiJ3sgY2
SPkPs7TAA0YFVN4sx9iE81+zw0Lli6xbsaJpj+7AilVD/yd388jwoFlvpPY95bxNwPPb8mz2nwJ6
5lWcvpuDD5/nBWu36sbkVNl5yj46Bh30f8QWwniv5rjqsSvTWpv4IboiUn68rAc+x5wQ8IMymF1z
GBDm/4iMqmhYK9xtUcYgC/341AgylDykEQuTSlKKcC9Fb+YG6TrEsj6A2kQrJiR4aiWaQVnLl+W6
FIpeuAOTqHVrXgWYzzuxQQf5KK0CRfsUH52ViP1WpG/FmOPzI2E7XX2gHvLtQ7gBiA8S4fjI/HSm
r4fWCTdmxfKx4zr4IucvojfSwFZ2M6GGkrJrlHa2jw4oHKYc8a6bMI5A+i1w1ZoL9CPp0JaAIrWI
CcUB5lJdu1QI7NamZtqXaQnBKX4ziL7xHkcyFO04qqeDfvjKWVNdmrwk9oZdkjjZkBk2OD9ansqH
SO28n8Vzo0O/9eAacuCVv/Se2XavABFr4MOwRJBW/d5ZVwseaSfNuJpQuQ2ud9BcI9NmuEv/GRsh
yahNB2U1odm5tEXORQR3AAMGRQcV2OTgNlfjnmgxLY1dkNY/WDKC5NsvCFeNQ+5llHZ+omNu8q32
+PIYLPDwTc1BlymiGob7HChc2umUFOtNLHNf5gcL8V+/QLJ777oGUT/mUu8UMfV2kgsH1t2ufuTK
gUGot3445K7z6Uk54qosy7SZMaW+DxGsHLXtj0737Fdb+X2tuM3R0uSoPEKpZveIjlfzFAGRbHpg
f895a/FVCN40yTD33ZlIWh5QEnhYAHRc2iJyWeFo3eLQnAb1ZH/nfV6LQ2ggkvu6g1ARo9c5onbs
va0dtETEHx2cmB82l+kHyQL+aqC4gsPBjYtESCa9She7htxww5OZtslV/mcqBsVhr+VUJPnD/PVb
qo4z4D8k6LB1UWcwrpW9y8WV4siWT3AxuOG3oL/ETlYcT3jY0cQveoy/WTjhPIgIzJPmGGCv5P7g
7ihT50PMfNMSH7ktI6Hk5cz85RoYYF2qXs0bzXW1oBDi7vj/WIXAblOj8o7sTM39hu3+jIQInKlQ
dWKJFoiqrnIDq2RVyzbA/FYIvH12mNwleyWdnCH9n+K0q0NadUbj4CfvT2IWI9yFwLv/eIouod3X
QLZAL3sRA2Agwuwn45rDAq1vmBYthXXUDdf1kLOyZSJZ8myNhOuaqON4YwDE00nmJp+l/razuN7K
thzrOphbEDKbWFCUQp+gdZsbcz/wbeyMkL29Ax/NW/KdYBOkJMBoqC2L5THFCl/ICIa8wigK4G7J
K95i+bpTdPR7r0Rs9u32I1/UwH1eQXmXnhM0fqpKb632ZL9TR2mi0sClDF2cNN2NPI0Hnu6kvZ5G
uZ9Kd5npYsCud8YQ/nHBPmdlpGOYpmemf/b3SlqoW+i1Vg6JDmjoLK8hI5te/whK1uSNChv6uYmX
eQ28L8hBiTz5fNc0l5Eqi6KrC2CdX556cc3G2UBD84oEXiqEOmaXhK1+sP/Nf5R0B2jslddk9+uf
we8Yme51jtT90gGDV+RMn5Rr9l/iMshhStqXJ9tCgtqUWonDyxG/53mSIal1jyrk3kFY3MjFmU83
GX6C/lkwkF0Fydu1r+fPx0merUZLQ0xqmVIU+G0IJqDsQG8Y/u2nNaqy5+vwRGINFCKJcU5Ez48C
A7nrF/iaUmiao+RUJXqAylbwuO5Rlcs/Ihh0FinPwTTCEqPG2U7JbQz28OKRZP6J9iGC0gFbtgIs
ecTDe5bu4DlKt1gaH0BnlUKt+Ne3Y6uZi/mBShQXjEsqNMx7Wss=
`protect end_protected
