`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11136)
`protect data_block
ENeK3HpQg1FhPE8ioqyGP78H+XuS7d9d/OOyKqEEWQebFdVZdWbJnDm94BDDADlInGY+48O+OMSy
8huXzoaKqEAE8N4AOKol08fObpRQQofXRICYiErUPS7ln9bgprhnCjV2/NT2cX661ykxeuXItFL0
yc3iwKNKw4U8wnQHqUCWzFwMqaRQYlLamYXCQqm3AdCIdm/xW3EQUHXWUtR5SSyKK8G7pcqCixbQ
pfgXTpucdt1owQv8br2eX4xfcuv2pblJesq6BanAuMimEqoa0WagZGonjdxvKvxdcLIQuBmIOwN3
2SsMo9v45FW1N8A7LAMGfmZTPPGVBY4x9sMGmdQTPt5smjm8W5W63CatltxeuXTTLNQwA2d+djii
yIAMRVX15cMgjK3ttrCJv0SJ36m+1p69no+1HafFqv0W5vz6vmmUAsAlmR3Gn4aeQjeT+PWVDcAU
g4E1Q1JSO6GpiRyLkHCZtT85JGB+xHjykN+HvzPyu9eScxD6q2GQ8FIwE/qcc3cloZK+i9pJmNsa
uOJcOl8dVP53X2DR+4htNcRy2kvBNu7kJwMOqrmIV8Z+79mXrfxmYmPaVO8l4eBJ6XP+8UuOkqw2
C+UWo0Yun5wCuLeeSO8to3EOWWPTGeQXnnjqweGSyo3a9S4mPT267860Uq6lSQTuSuWKnJCxF7GG
mE93ZA/6dEQWDj0kD9Cpi6oM7eAbx8NPu85330lJq/qj85RMcipMvrqjNlgBe43Pbj0garXb1PHs
dAyOlnq9ZtQmiScvuXYsuMgkn/Gb8vyUu+EeIWcA7KiDMPkoJa+CG/ezLc+S4wl09BRN9I5siwlW
bEsftr/tuo32PcMk7RdSpajYhAaiOJkSQxh/CD+sp1DXMHZM3HsVpGAelKxaDErvRssf9dUFvHjZ
p0IH918+A35beLBveaA/KL8dyMiHUx5kbRdpQ8jtR2aYG4AOtAtnsgqp5icYgpqK0IPzyPRKKaYo
8WclHs4B/sQAvxlo0r1i9uJNOhtnyKkxF+uhYS6tN/HqFJ2wQv58IWC6l1+DnUrHED1BXiS3qeVC
TAXmFbeCa2ps0zuYt6vK6n78KEpv/ROCTccoS5fSESwO/zI/12NQmcXVyKG1O/HFjt6TncpSwNXR
BNnTfUNKdE4swyEyGhTQ+Mh5h+saS3Ng+yBAg6/l3nshGkgDG7DRhR1zaFFb841T9V5pmRJGCyTe
Xuncd6nYjvTxqOdYaCYQaBGWzvxQrFMU8qHq+rc4/Ox0P4W//r6B8rE2EBSdFaLj25+RTb7Co1lV
xHri6pLGMQhx9mTG4qVTmXy/ZPvyjsIrJ/q+KN2cpoaHr5dtn0VhH5vAPtbkw6TrXtkifuauH3EH
aDLk/eqtlF1EqyMuO1HzojXHGWxkqgQo5jPRFmRTS2gOiVmKRETArgg5lscEHQeWhD+ZsXY4MoVw
dW10iNNuGm95QpnwYqCDv8rDrYK5AqdNw2PzEgtFFc8KqYOj1o6RyA2XRZp2xlLghlIZde5QIkUG
i43lJzwRJ6AZOqydtQ64gAtDl5u/XFMiscN0fRSYFyLqq49VX80F6Y8F/JXNBJYLvCHHA1An19MT
Jh6V1lEUqyUQH1pt+KTGALhMgPPHltvESAE8zJw4QiUY/i4DV9egqemrJ+KQCGAO1uVJUgh4KkCf
GY7OSO+QRlo2MMPeT2Skup182b5iSn55uGScdpfdBnOrvCdv19ej7PssoLgVugDB4KLZn1lYapIa
iGh8qo9/ZMdK3R+56ysvMCQL3+kqKu+2Dl6es3AO0pL7YaxjRcjybR95p2hvL4UbkBWhuKrExxwX
eVBSpBvS776PUg6zG8BvTrKEhvyKsqOmBcv+FmqPdHxNVCQmdRhPwxyKY6E3quyb1cNnkbf0K3Hi
aVSdEiB6bEk3Bf63Ih0jinnOb1Z9S2P9bnd55f1lrasuvGePQtasyDcXoinSRi7IyhTROiw4KDH2
GxNIVa9kDHNn1F6PwhN0ggmRVL1VMYwYaCmQG0qAmZ6yXFEq7zFd7bFqHA/LJr6WB7YvjTLoCcc7
JbKnuyWmchXY0W/m9l5PHret7zCcbhNHEt4ZZlP3cSqX/A5NyrySygPtJ6PWqHJIX2EuYk3Xu2Sc
NMXjAYRspt0KfmC2v7iYLtQWgwNiZNED2Nb96cmsZJK8vLOqU7axtFA7Z/LtE3vdOryCMBV3QDOi
XQSD0oqfync5uVgKsgZXWV5NUAJlRjDgoHX/skw70WhjosKzGbE5QOX4T1ExaptbXnVCywlcV6+4
WcAFspZEiskOveJ9ruAH2p9Xfml1btJIpogCvtOalPaezFrGOF8TqwWPtih6qccIRVMSRAWpA7s8
dpcLIXQRo25JTl7qJ4rsqJ1zhqWRzK2s7fGi4TC5K9AuLbb/5X4iECA2cPGEgcCfoO8A5xa/aB3n
EbHVCp4OmLWr3n0cDMgtlAJsZs0mBos3AtrcJyK7GAdhxJmqLLsVwnw4tdRwt6k6trNfWbuNCXS+
zSYhK565b0vtjDIJbGrRGjhNy6Jcg8SzZy8tuGQNt5dY/wDtiWQEu3wes98/c0ve69TQJSrrHVdX
yrRuwIcY3K4FjJ94v3SztrF0T8+fRTb2XnaXTL/E8bpJFxuzNc/KFI1BFuhI4VosDG9XQL2lITS7
tWhH3X39KIsR/a6x6yVBtFKqRS2nxLHXF8UDzXuJPLbh1g+pcaiS4ADX4HEJKY6H8/eelIYck7V1
xB64O7nWZj3SdHln5tMJ68ydjimHYck7VlXT2XjP/IsIHNSdTRPCs+9Wlk7Li4cJS35aRTClIoKW
mdrN9E0KIYwgSKIwL6rBddrPZyZz6Q9SG5q351219Gekt0Bi1W7npWad56L2t47rOBNosHad9HeG
X3D6CHpKkK+U+78PXsekDvCAd3nd1Ks8PRy2Cg8mceFv4sThHdZMzZr1Dq6qCUsivOMzeshnHfEI
4nXMHTHN1+nh2tHw4KdvKw5aU69GV9n9dUBz9KNky0LqC09YTS04YBzL8RymRisS7xISNsyXLX3Q
KAKzePWOZutvXFEhHGhou/5tJVISkxoattU6ZPRHrF6PkehSQoSK8zcbzcotn8n9EUUQ+qz0Y4Vw
xSbos4qpS8+T1m/Loxu4c/wlig7q+2KRKieOigMY1nCFopdEJqwyTM21A4cQtS4MaCLZTY9cnu2q
dQZInsyBoy6A0bH/VRcpKkwN7JxCLOVp2bwo3P+k8bZ23FrONIknK+Z/WcCWiW7XRJ7MTvvBkgpb
Ln/6YdBeCAR7OqwAzp82zLA4wQTeNa62QgwcsuyhMiho+EDoxmi1LqhRGnTrnvTktUubkp3BGJxb
Vja4gQ7TXkLbKx3BhbocEemr/pOcDV9kqUNJOEOynmIUezarIuKbrIbS6TTkLU/wfZLodScujjYJ
8QUYaf+7sbVqkFBBqcbcm9mu8QatapCaOYfDt9kkh57DaFFVGdDTAPJO6V1OTRxi3EyT6iSyu0dd
iterjAM+2ioUDCYnRcfq5/7/ZVgV9Vfy/7cr6UM4bPiztxaWqc+8GAuW990BZLsBL6rxwCfRIy+g
M7fnnvWqiy1tvkUM94oL4U9M6SRAtJsvguzVqDTWDtSRX8/QetTpTvMwrsW9LLZ1wkugMbLUwaSc
m9oFeR74+w9JLqSWGnVbWgfOUb2z7NdsUTN3V/yApE+JEyfcp+zpinxLhSPdCcQPaSF7lCijk7ut
QRAJwsmkObZ64HeHqDPapyL5gsKz61GRzbJ0+sy14Y900tuDsPJJByW7zvSva5Nl7nM0F/JSJWpq
Lxg3EyCHrhadVc89xG6tEqhmWi+G30E+IxFESO6t45d+P/kXZ4TKUhNKRXnzWtUT7UD7C53V4TF7
OykYkuKAs3xfHBm7+MQ+np3mnsh588rbVLenzOrLtwY+hpYiX4LsoV4pgn27WvpIT66ejU0Hcz8s
2jygnfT7xc5gd83+saDv1V2/etzzmDIEjJzFZhLAAO+cGRwYP91fpZxErQf6mc3Z57hv4X1vv35I
0GnhmIfIYTx9bMZrfmpBK4ek/ko3r8AuvkvBffWJy/0uDsx37L7fHQEzLBVztTxmN/pLXckWf97m
ew8VTnWfbt0P4Oy0xURj0ATnlalyxY1iEB5XrQRyS2o2EmRovrHgLDXp+G+7QzLz2xd+97juGmsq
Pxre6B/IWTD7X9z3nI942czHIvmXRmG2CGtFb4ZN9eOKuu4gO1Q/EfNm8TAGH+HKxeplLKbQS4kQ
G541hwUhrN0sZ2a3UAVSEzgR6ddylt+G7y06/QGCi3ndeDrxgmgROIpPq1kEG2cu7/s+jTY4Vb0p
ZxNiY1p1a3Ryg8uwMoQ6q0g/65ovCkStuXHWzDNPqywp2YwensCLImKb/IYNhGpr7y47ecQjFdsF
2MBLd4H3poxNXITNKGFysoYoiT3bCcsbnBJSABmKfUUGRQw3OpA/jYnyk+xfGRAX0K9n0LJKNFGb
SO4m3FJGFpZBabjqXts/g3QeuBKy8w+NbEvAuiVaSJJ4LT1lg0yUSEYz/Ac5/ezUAUL7DYfcEfB8
vYotiIDcLr2IFHYfAqcrHboPv2ySmMuFxAHWYQ1oL/jhPi0VA4rVJ2eDfHWJlMloDFgeVqizXS0l
sbYXIwZQ0fXQpQ++xAVHHjpBCuWIVCp/9KAKR6K4avakK7xZp6AmRYg3MOgnZdx9zCKZb3Qjrudz
QniS4fbiqDVrak3nZAJBWJGWfdyG5vkht0yyFTeNsTAD+S8oz7aeJbKpJ0jEwWjhRHAUkX1GhxTS
QJoRxNzmlmD3zgi9b4DHIURQbD/xjURfzY5Fg3M/fG5xi91LgkFqwMVMXXMXW4V7H3p1X0OBHs6X
nW+2cBq1wyZgY8MGU4bG4AmaUFRMcLb/e8HSkrspfTUFB7cS2/AaYHqC/1nercQz3iu61L6JZFGK
isFVmQqWh7R8MDWmFCrsl8AkrxalpLO75Nk+I6fKw/oDzp50Yla286XpKTixTBDbBdpE4S+LSoUj
gZrLsOrfFAG1YklmucLXyHqoys67MISlUt4YYhfSd9ZQhxhpydlbIq8XOHrXoiH6wb7hoP73+ccl
ED/gYo/Awo1WoEiCJrqoen7yP+ZX717t6Ac/x6EeCT9D0/LQKNF9NlHDAwqtHTdv/Q9t8Nj0Q0X0
BrQbp03wh7ONvl6cVsnSTprvrCPUHU7krtRoMcyZKIEkULGjuwRlGPxlVbtmJmM3z7fCMIwDLQK/
QYtxByeAUUJGtLqY8tuLwKBGmNxYSEKkr+TpPqICmB28s0eJkcu6OTVgxS8XAPSe8C6ePa6i3tN3
ZkMbsiCfo+TLLuTQuRWpvYWIjD5mTw1GdxKPtVBcDVxbEDobziD7iSUD7pi5x2+9/AYLumhZW5ww
uQ+hY+FFU/O98UO+ekAJ3t12hTR1F2+ZsmTU+yTvwV0XLIMcig7d6h5pkmv7UGS0xvjRO3M1EDZr
8079U4yU9eEYyEMlLPeeb06xP2mwXNY76pi59YUnRNbQpTO2CjBDxA5XIcD6aAWsf70Zi9Uzi1E0
h0DjRwv3NNd6LpeLupdVcR9HRsCP2yRhqT/VKlaQYi2MUs4WiJffGUsQZxonoKISo8rXzpkCLt/o
JuPyaSRN1lHgypqExpcWhB2Femexp7kJEqL7OU1dc0R3Vhsi3ewjd9cFDeDs8oD7SrHgD8ooc1Ee
lHU3odVSJBqtVMqflT7CGVuLSF4wEzcdtTg2V5jBTcxHumPPRTpQxt6WZ61VDe9xRwJcAjW9+nrR
BjIfWHVIr6Q9PEmOvXCMkIefiy9IJkb79FNowBOiDBWe6lj2m/paOgwZiGFHFIzMWOPRtVcIwYGP
IP6oKF2W19tutGA36s1SRIfRhlw1l/zfJpnZY7hQupXQAlMEGxTWbVY3T/NMvLAfDK7uOf/nnTho
Hg308DBuQ8cw9cfkOxoDh8qv61gdHSy9pDDRdig6ZaCn3ZfVpqTBQOCvztjCWhd9sVzwqQVh2n+G
Pfa3d//EYt9Q0J32A9ZbOewixOp78blk52eolx+wnhkSdslIDQTYfdHUCfQPrYy9nc3g1y+wx7Oy
SAOK8IKaWiPgWi32TnrlxBiX/TGuivzt0emJyQgYRz4QTM22nUhZl0W94ZpJyovDwidNZAUsdofq
j3n16YFI1Bfw/7NNd2kv8Lb9bOqT4cVLXlLPmhkRt8fr0qiECOlGm7UQe/T+NG0MgMrTbzPXk+1O
oZyz5wkLIK5ZFVEBlIidUJMVOVh0ekAmyoQwY5ABM5Y84mQbtv6Zzoc6auFDQ5CBpITW1RvuiTm7
s70j90jokTNrIAajOnEq9zo6gVFEAOC9D+N7/cTRliTLWVGUJXg9hOHad9YxBdibg58RKvRP+OEZ
cFMJBgKPxLOsdYK1dFUz680R+vOwc+NLWrz5RK/BChdpH9+p3ewnqoiXL8aC/hIcEhFjwPkP/ygR
cJkDtOe+hVzd3a/ehna2aSB5UUNXur0Xv8Z7aoeQ0bM0ZtO80WVtLc2FP89TgAxXbGonomqGixj1
GPiSwpSUcIA9z3yweKywIcq/etY2toUfY5kcXfI5fTNwkvE0kS7X4lxAQMO8DN4yAgQTc2Y5UTeb
5qxR0nWymka1wYIiPN/siqr+nXm5lGBUQ88iyj74FKIlJOntSlHKyc4MOXE+mYYxlhl08011c8EK
1P0bxgHdpybDn6xl6s9eKfdAF5im1I1M1KWNTME397+OrqXCDro6tjgEf5jHUQ3fGohq9M+Y5MGQ
sHRJJgGFpOOFzWKfpCbJ+vKN05dcRdUeLRzYzU/qI/tVcd7ZrC+vd4oGlVYueBxmCivT5Qvkfh/4
T5yV+cqQYeZmGQwz9MdEo1bGmgpzBTL5EKBrUB1RZmntKfYPShpUZezmGMlq0rdsMhy3DF2h+9/g
BE+FXm5bsMmQBGPyKLp8RKdjX+j5rlMCiC5czqLqIm1pKv6KITdsmrh8zoKPGM4pYkjEJkfu/hxu
U38C6VJNDwzZNXAcvFJY11CknOjm/aXxXd8ACfTBA5Jvp7eZIT3cRwzT64JP+j//ZsrXI21t9PKc
pJlk+WKxj5DGbNGByNXuAPY9vEhMKNLJMhkuBlWhEqIjXQirLcWk7O7+RWgP49RFWQ3yonKxEUDg
Z2rR35HGjovs3AIsoTX/+uNSD1iYidsVwRol9eEfbozkxPItJFq2Vupd214n3ExWmoT0PKv2QkLG
tew7BO5up/ecQADH+nuo8Ryc9fWEvgxXK2tsAhKWC8elSzX0D3q+dGC3cv6x5aSnjJX25KPTnCQF
dy9vI79y2UjYjX6fl3vlhl3wjZgl7umWgbmYyxjGYTzhRf3l1HqdUmBmLlhnnkDIzvC1TFVrb8II
7fzGTj7ZYhcFOquLjTWd556sXPKA3lm5I/kxKejph2toTjEDi887BfX5vhGR2GaTaGFe6U/55yxw
6w529S6Rl6Um+2rz8+Ymc/hDxqy4MPS9SCGTyeIUxnBSi3R+gEQmnnBgZTSCoZBqPJ0nf4SVQ6Q7
CjQEc2pKReY9dCD6j1vGd/mLthSyR9YKC5mWEvsLcOsU5ktepAAZYLVGif+YYIof/d/JVKCBFX+D
Chyvvr7Mo6HoYbxlhN5hzI62+uPUyXYZJSpMzcUPEXBBWC3j+OKC6ABd3Kd9FhynMeWT81Zyl4/K
8NSTYUluGdZMEjC4MQPun7x5kX0NSJ27ghoYcDdslNKViWsGrYzdTT43jYKqETZMkpSAKyAx+e9K
c9qAV4S2m62DDfwJc3TLaiJmetklRwZKt6Hq5KkYfbGSX7G7xmbiurmWray7IIAeh40pCW9Pt7EM
ZQH0y1qwqz1J7VxV/qtN9S/z68uUDCDM3iHjyI+guPxf5m06alGY1dy5JuhR3Xby24im+ZQ8XQ0s
cjgjWXnVgcmKeTOZem+RDABXm4T7+d2OS+0p/jb5sKY3HhjMSUCgskz5ubjCsmfdxFHCzouKWutc
YnrVtSi9JnCufwJ8sZYFx3wCEPOaVmgcLlgWB4diNgVU0CQPFetkz5dfHLbylxgb4bNs6s0Kemmq
Q0vakHKYc+D2N/iQe+CFwwQk7xMRPyHWHxPzmKUeJIW428zJShTIkiNpd7m2ci3SUZuUsPMTZD3e
Y6nGuQi8obRdWL0jrSCmDBPbkvJyK20q8rQvLyPMg42gESyVL35VbvRysfgGDTZwknoce4mjqGqo
8Ul9vTrWBRt2e8NLFEUfewEuCQjkctRuzMAP6MluoYjinvD5MG81ww+bzqTkgBgg/gvJaTa+H9jG
7MmNr0tmJPfZkO9h2hS/8vqFUo/EIxxba+Um3i/OMn9Auumw3KyY8YXmcyl6Dugo2ZNebRuLcJtk
1sl/yFIjRJ3ZVXt7ueTiQ7HjnDj1G6TCoCFQzyA2DuD2x2Cp1rY+VpcsxbqhMThMPeQKq7jlAncx
kvROdcZzNQGwKNMGi6BfQAr8f8PnH/PVQ3xbFr51XJ+gv/1U9eFB81LNKfnqoHejLvVLgQjqmpp2
M6CLqGW6nOHfu0POnY997iFbe+SsNNI4jSqtHjJvNyFh5sCQ9hOUApZmAvUQfiag4H4cTSzNSOtW
uRmg+ivTfzz3Y6AS5PdfKtbGdem8iklZi3LH3vasyTinL48KqphLQqoGCwM6w+Hr+W9Yu3jhpSH3
2l38JuAwvNTxfXbF99anYGz/s2IcDyAcDXgl5QSnuo7Fnaz1KPXGXnAPN1NMdflPEYnHYPGSu33B
OeBvlc0QHW/1uA88I0fKX5g/5bwPCCsh6CwRNHNJCpfKVkQMkbuPE11HzyiOze2MwDbyfyGCnSjH
VC9Pw8TaDRyQchUtP4iucXAI4okXXSismVpa13AycptpzGfb+23WXlEiLS26BObbK61Dn6mEAwdB
uM8euWENYSrp4hEotjfwat4wK9/pyf8X9f4YIWk5fwonVKxJyjnd8dmG8ZgHjunwywaaPDtFui9P
FE5HkEwBoI5qfylqs08Rh6JDqNVpEAB4P96UPHpeHM92YOg44YXGuAJ+IHQHCWUTgp+CJq+hj0eI
Jv5Hf6Xwo4OOrxZCTdHK+s5TJE5wp0mvmcPkX4idNfcEmTwhDorOH14M4/RLLbob0XPV547qERyk
H7SBLPEf0Mqzs32EpgJL6XRtHgZtwPCvqO8cyglQi2e3NWgq3BWwDEU9stDmUfLlPCylvUnuS0kg
CYQdii2hHNQpiT7vKhBw/oFu+jTOTgWUU/bVZNY+fMVqdxo5LuWEI2WDKVldzTTOao7nXFeVNwXU
HqJV8f1BfnBe57N7m/n95BXC1rvt1lCtG1zbWb/fxtrJdDrhl19zWLy8q12riJ3/qxy44Hmy8E06
EuRnZG/Nu3vDSNASXQYVf1o2FQzA5yJojM6b1VpHJARpmCg1UEkrOp1IQcVltAQSu5hvuH0pB8n+
cpLLB+3H4w9Qs9YLU3wnTlVBf2J6fdTtxe+8uJlCLxldabcEE3gUor6S4lX/ySM5EILfW8ivTron
f8AvqCFEjYDz/MsiZTPARyvizFl0BHImvlJjTx4VU+2K4ugt4KoUPnGWcFx9MMxsT77qRTlDxZ2W
Jh5ze7IMdDRvglneo0RELztIuiLqm5RSj99unjS7o74r2bXsn+SeKn8KKIzvJvRiKRZSRqjGjKpi
HqogmfZXjtTWm8DWu16ITlHzSXWfujLASCeTjxJyqw7Rcm27gitU/tOAslPK0cQpXr3W4q71XJf/
FXrdYF/FCJTjfh3BCHkM7uNLorRff1g0x0GPtB5fYb3EjIkjVCtiBENBEQo0mZjLjLfxfToXuFaq
9BFHsDkkAvQu+ubfs96eey4ZYR9WqLWbI2hM7wwd7m+si6v2R8zaU7vpnxfU2OrlQaLqf732ZLia
PCxAdWdmTDMMp0yto3ohYg4400FlrKL/tbPaCCrpDvOP2yDLEJBuWLLEljvyMMZ0y3ybKNnJRrZG
Bpb1vEgs7HzV1Ab7U8iHSD9GromiKmBrErs8I91m8658w7lmykKjPVC/0u9n5x4pVtRRfzYMG6N4
yFIWQvmvXpXWZAob3MsfHq6yuWL8apkbbOma4kD29mB2NvKRmN6fWD9Pc3nfuELsKv8CUg5rLV/r
f7/SKTILMT6H93MNByYZ2wida9KULr1D42HsFp4rLXnJHkT32DH9XD3MhNfwLWLVVFFXd8Bqr7LU
BJCgdhDgL3rAZ7oXS/SEwCrvyce5wy8XL1Me/m46jHfs39lSlq3826BsDwCZgscu87k2PDW4EPNo
AZUdQBJ3aeTMBKvxOqC2gp1Y3JKQzvzXLr3tR8vhgLccV4OOUCZ9fqQLExZmc1GdrWJ0OqUiHw9p
QoEzmrNDP5DXo288o/ylT1BvrntuHc7Kg8+aqj9MLYDdetXAxkJ7dnv16snLcyj03jVxcqy+Xisj
hRdwhxygkgxKPtgW74zi/vKIzBTmw+EQgk2Y1PT2hlSB+XaxKiQfn8hu6IHtyMY4z2458NkVFutt
FTgfyIzUMlew6PlHBzPXQA6MIujJzZFTqUjGHib8JJSjzNzj7rJpH/sgK3Z7ErAtNfJiTrV5BvKi
/XDW8sYqc0XfdyjSVkX/1bTaSty+AIVtbcnbjeKLCwBKQzHcFSaU2sZJJh59uojjIugeopthot7p
0XmhWxDGJrzFMwhWcFkSiIgkG3oYKIFplKGKqgrhnSHodnKYrdKxxMrjFjl4JrCEaT/Uly9g8qpl
mvkMm9Lpsp2ZJY0novyTOM8FecRSLEMkJAV0kQRzZQH2kYC8M8xd4SWaJWe19rUz0AYx2LiSTSQw
lvPOXRbn+E7nkLYnjx3pwahy0UCpUtdLdD6nWee0wQQLAq47N626usGE7Y30sD6Hdyso6/QBuCI7
6/usY5rtCOLvMFuH/oI8Sf/PaxeGbz4dbtKqqMlvUkENZv2qhbC5Q9Y9H6hA/ZK/v3h//iQj+FTq
f+cuwBs5AS7SLTmujlsxAumrcJBdUAlGm8ALdIp0FU02rj+6ltDe50ga01L9Mcs6Q9vifM2bRpQ+
qPtf6VwfITUIUJUvyB8H+oicLGNMGuYXffClW4w2j3C26hxBKri1L+hxB0Vi6ibck3qKisFC6jOh
tpeg3McyHVW26T4xNuowcXAn4P+tcYcz3SOrLnqboKDIvly2S9OromyCPPiZJfnca9Kj1olGIL+y
V4Wcz9Ae1l2wBodNLEW8NsC0tIjVQEJJ9O7wnbBVY3aYVZ7B5F2PHPs3M06P4bKtOW41d2LvHOm9
uw1xojm/6XFNfxVKPklvNw7H2Sw8PT+0ipJA3JqZvIU1z/34kE4O5HrEsQ8RfeFQ5ucQLGkmxmN1
KILt04+pEScD6wRUOWPY9c98Eu1tk/2Y03BwuC2F732IkSgC4nSy56fXDQ6q4amzb6zGD74URcxu
Kuqu8LHhx1pulMZcy+hiYUDfiLskR/G8DDrNHjLZOUDsPFpHqkaNA9ytY/UnUttXj9TNOENJlUTp
yb2xw9EgGFOO3CVvRsS5cvYTcYYvuk9d/fDynDMYBMznbectq5S7pd+cDU/SZ1mIN7mA574VheK3
wXUdYsgnC0WHreG7KlruSisy+15mvTYM0B96O3Ae9Hwa0uFeSSrmmv8PQ9dfZEWf9k+oUeatqK2l
eNw8eId5H64lOf5RynLO0HNwoaiilryOhMR63capHq1kepYdzjr9B1cQ7iZ/Pg1qYeBB0c/Dnwcc
PzZsuenUwPPid3nXrJytDgCVqyCAWI3iUChVBkjDB+HYM4Gyjt6M6926F4WybRfLFHg3FWmgoA+Y
AljkmbdCyov898d3tQ6eRJT5AXhLQnrF5s7BkYiH5PmIGFltvl+9DDdkl5pOU/RcS7RllkOKpw1k
O5k5lxwxdzji4wDgfh1BNYT2vhWby9pkLoJ60D2cBFnwjOO71iXZVkNRyEU4NGulNWAocEhnaw9/
TqgqKtn/YMh0f6K1fdDEWPxNsOSzXRICzUmRWskHupxYddqFz+2ok9CFzru/foVzsyq9uEEoWgwX
ZW5C4je4cCQwba25Vzb7LZZNb5fPppXjWMQ67FAFWY5ppoJXh5fg20HznO2JA1zrrAogRmF9jaU6
+xQbyQb+pTKIoCDzAqWKHsJyd+aeB/2gevTvdqYSmWAXMWiKdod1I9dP5h86xgk7EwGBU59RxtBw
dxaPRuC2VREeCFrL6RxQ5pgit1b/THny0qtPwzDhIJkpN2bdlcVQT51Fmyg5gnclClx2rIs+Ww2f
0begSh1A6Qk92kKRloe/7/k9Utut0FNRR16zoY0naN+7Nwpw9hS/jgFSt4pu1l80leccD+6jXzCy
f1Y+kEU9gXCqpYLK79d0XRy3Yu21HIGKswpACt/qeL7GIcTBDmIA368wRlBRzEwgb4fhTREkp26d
mdoxITW6Y8dQkdGn8/ELeylDk3Y/euujb/zmia+4zZAyeLOQAmWIPfgIY+nfvrtb6H9t3n83juXG
Bs/LhmkrC9JPaROQcTsVYuP2/YwM6nARYA34IsURkYQNsjcyD8LM7FSLnvx/z1abuvxYD6X4l4tQ
3Ou/wQS9o/x2EXDqyM/5vv4i95WD0CIXXBIFGiA687b8MhwTNtDPXYCnkL2XAEQ+fy1ErFVO+ERL
pKC1D/ybPeHuChIOl8L6L486f089FH5u4za4vh3ctrg7WylvfZHzIiGBHNgiScLBTeupl5vN4mm0
jL9BXDoNcSwOoFmsCL37NMzXz/Nfu3fg0uCEJ5/Et+kYM8VRNwh3PI60YUjcLI4e9Feuj321aTiG
oPCm3OZhy1SXFeaK1DaFXWncrry86KoV6QFH1nZOaDoTpmQuFrI2OVeSRIgeZ7FQKGY7qDsIdB3v
yGIlaxFeGJO2jy1bs3/8dPnoQ384iIQCMNPqERYh99WtSd2j/DIw9HLdOb1C1csw4M5ecTL/scMz
R53maO79FZNTG2hvUPLGrxUGuz6Ok77EYLr8+y+jfzrDwNFARVdyvdpg7p49J96yI7yIfJK8QNHQ
zVfcAFUGI3haOj3JMb6BoEVeoiHqqXvuOizrhnqbkxrPkYu88xSk+hfcIsjM3A01o7N7LLHGOevQ
IX84Vm9nsdyAN9J+oy3Y76GttTGXGJlUrOu4WgB0/csZlWJjY8SLV8HNc/DgdVzIgt/wnu14qqp3
zCOx69hSxnZSZJhT1KOzJE7ux8iZ6izG7tPwM0GDgmQY25tctT7M0K7vez2mYcxabWbs9foOFQON
7pffzOovf367i+KFWgFk2vc935Imrx+4asPwP3WHBN6vWBbekCMlusIanwQ71q1HGejcvYTSOfT+
JsNWHxpqTk3H8WxUD78j2t7cO9GMlFhPjzqQIlWtTVesz92eK8nyzPW2GqjlT9t3jcIlePGVTI6Z
FKDAU9O93BavkGu8ZY9ifl/zgHgjvdBV70Cq7T4HSTydyRHYKI5epsEu8gffvhLdJ7GvA5YY0Myx
q7kogkKp7mdbgKIOv+3iOO0M1nbyyiUz/SHjrSQBhlxY1mY3f6/tX7uDyngJ+RP8c+mksTPClWN+
jYsOes8KKIUghFZvMdwPTE1ej2woepmejpApqDZ8zIXr7RyaGl1uSgV0xQqnIm5u3c08LeBl4mta
+izI5IXo37i7r0ObpScO52syObW85PrOXbmRwLzmROSx15/NS8kHaXqV0Ku9oGyCFaQQdGvX+c+p
EumNUBCmhC1FnmKO8YWdisH7xNaZZ3O2UcqCj13w4dZMhrQyGjP7xefj7cQzYyiUZCzB1O4Z4bxz
Mtmwxaj4PsRLniEBZhyqLUp0awetFl4212e6pukyuKqvMRSC9yWQzznckPBrteDjcQYDwMiPzC/H
bB9EZbvU2V1PH+dG+JkQgOfLpvE17NNOmR9NbwqSzqmj5zk5c2XXEX3yNwEAL3OKtEyyWwKUUpMm
DSfAO0Kb7AZ/Eqrl26N34shR03rfKzxQ9K2CKyo89Sul6jUW0K+fKGsUJtRxPgiJGKQi500ra0PC
N51aG66r8Iah43+8CtEl//9439+Ou7IC7U8iHd9EhZJviKNbOyXxSl9VAPl2FSUOZ/E16c1wKPBQ
YTwcuJ4BfR6Umtrp3JmHYOi8tEDKK3JoQb/LKjizwFJg4wHh2sUbvFzSz7DS4y7NWGk0WE4E3vSZ
tEv+2Ho+os1pEU1M1Dr9RkSj+U5awHwrA0USbQRGZbWzeJG2q3CS6XF99hSaHPy+H8/fLK9+7hhJ
cds2VQDltzCoUCOZ/08Vi5vN1ELo5U2yGWuobC4H4e/UuOdA1b4+wFuxwi4oeQgJ5jwHUumtla9w
ZQLUAzXeIYUjYh6QXUJbrMvtW/ycYM1yxUtt+PoiFTMUl8MBmGQqQjWphXuI+5BLCAzvLE0AlZm6
6zU9C8bZe3lrHBoffi/sooiqdTnQyMsxf44TS5adbg8nXjXCScj6J6YO6kGekV/MYW6X/vLleAof
nKJXjYdiN8hJfVUkoGqvqbh17bG7cLrvbr63SwTis7llGkPHZGQ/30jL9TSvy2MWMdKdrXwI2WTC
+tVYGt8xq4KrLUiZV9zGoVPB80AF9c2+xc1nheBbw2D5TNuEazi1vKvYfAX9M5MRPot3FSYlKyPY
AcQfwEJici/ARaqdy3dbrnLxfjCzoDgEZzlOcw9PbFmPCAZQZbJ1vX0I9P4A8vLB1/13goILk8cj
Qu4atxg76iMFy23lbjhApFEboXMqKOOD0hej47ETUwT1jnLyxC9idiCu7TyJK77Q1PU5cR1aLZ1O
XRYkpcrYr/zeIN0yxIV8sQUNkBMba8eDV6CfjSFgb+UvpgJ1vo8GTz0GU7lNZ90sL83dQIbarM2s
fWheeCQY4WEoMp33E3C7+qMlVLfW
`protect end_protected
