XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��g?�؁O5k8*L�|��F�ت:yo(}q�t��F��d�8p�B��κ~������ϛ'�����xO����Ģ۸����;j�����E�FS�+��,�0�H`��>#E^��[���$Md~!��k��Q[X�0�lқAH��"��f�g�oS4�h�f�,6�ȳ�7��1�`
��L�"l]ph����PpFإ��[C5?
�m�pS��3xPjn�}�>ej*�8�H-�Tֲ�4���F\s@1r�X=.m���K�O�I3�B�����@p@�V|�rx�8x�]9��9�t��,:�ćF��zY�s�S�XB�xcC�ϖ�t����2���r�-S�J��(+���8�"czq<�y���/h/-�>.ZX�.��3G�5Qf��Vl�?H\z^�K�>�8xk�"B�Yڗ�F�c���S
� D�I����^��Wr�=/�	+:��̣�T�H�R�NqmQ�4q�c���+)@p΍3��^N�(X�q��\��f�ղOa�j@@~�O�k~���y�,�� Uy�mU"�O���Uk�VY��.��]eD�˒TQ_ɹ�5"_�`u��^iB��xt'�F&�T�F��h�&=�hHRm��kζb�{����OXmj������lK��JE�qط���4�At�jEBփ���K-׳��#���˾2!��TWB�����_�Q4D�~}�h�<R� �Xߎ���өٚ�]H+�"�\?�<���r˗��)�r�XlxVHYEB     400     150��9��RK,?rҊPF�6r)���ޓ����e��a�>�8L1�vM�b��h��}{I��n���ȣY��Q)NO��	c�+��{fV
}����k{�go��!G}��EY���R���_��DW�u�I3��ԍ`@���ci������[��(��L(�e:�f��³,��Y2R�k!4E�M$j�61ņ�T�\3j��[W[���9�8�,� � WvY����/i�wo7C�~Q��|����<�7r$`:��p�Ԑ��Ⱥ�.rD1�	����B�mK�fb�Bm�?��1-*��G��6�FJ=�
�i=\B��(N���p�j%J#o�3m��װ��XlxVHYEB     400     170��=�,`7N���T�q�0���1�b=rY�2,f�;������)����vN�;��7�Ecd�'*@O���������u7�����^sP��ӥ�����lWg��d]��9:]�����4t^&��o��?�z�,���nÄ�=�� �d&��7�
)ZL:��@4���%i�w�t��O�$�����g�a	�=���#X�X�(��z����'���W�oo��Y�������g�m��/��c�tM-���>dI�)�5�r��X;M�UF�r��JW�{6�,�/�\1K�����j�L������%1~����p��s|�=d(i@�O� ��i콆�ѥTy1:�&:��Pf[{�^XlxVHYEB     400     130a:\̿$va(;x���� ]�lԙ�����W�o\�8%{���pӷ'��[�9im� k���"\l�;U�����_�p�S�᷽=��;dʩ
��dՒP4	�
�$'3�ς>��ߖ���q~����`h$X�u'Mz�t5D  �����RH4�Yf$^��iW/��PYQ�W��Zx?:Rh�)7���L�C�u$�v�H~���˻)��)��w�>	�7��}� ��y��U�������kw��S])dӎSa_+񞇐f�94��b��-�4m,�������+Ld�yϵx��K�j�XlxVHYEB     400     100S��*��A7o!�VQ�,K���.4EU�T�j�o��MP��9ƶ-��ʹ9�P�&���z��x�I�N?CcZ��d�nNC~.��lkZCGL�q�]y?����	���Q	A�̖C���:�mKh�&f��A�ou���A/[
��[�s�����g�D� :_=���3���qA���g'/, ��jnj���{.������'�l��% �ݲ�)�x)���w[������j��4�G�D+i�.r�C,XlxVHYEB     400      e0d;<ۀ��/9T'��<*�"�DƟK�^�9��^`�)�Ë�q�ֳ�U�TE�2^�~���;�6�}X. W�'U��@
1W4Ap�d�0v����s�5��U�����&j3�ʄGp�O��Iz1�^ɿ����? LM����A�V9N����R�:�������-�`�e�;ΞX)p�j]�N�$av}qx���I�lN��Oa����T��[m>l�v��>��XlxVHYEB     400      d0}��[Pv����2sOP^*�[�<�F ��̌q���3��ŗ_�㋶�n���X����صA�j�,`4P��i�#�<D�[E���H	%��d���ǰW&�n�1!pL즫Iܷ�[}�H��2Y'�{Y}��ȏ���ǿ�TC�A�T�:�^"Z������C�c/;y`wH�h�H��~��HJ�F�$�tWpRs�@0�:p~9XlxVHYEB     400     120|�������6e�NN<�!�D�
ڵ��q����*��z�.�`��C�-c�� 	�p�B�B���~Hl	�=�LV�"-��8���
a�kF�э}GbN8�zk��ġθ�Ah�ٸ��I
.����7�ӄ�qq�	=��,J���A#ؑ8��7Ky5��!Q�!��F��|Y��`�-�Q-�ϻ�W��>�ÒY;��W���'��@2ǻ�@P��_<�Ҏ��1�c�V1��;�t��G�e�Ű��>�v�b�w��7 >�*86�A<�{A�o2�	XlxVHYEB     400     180��y�`���'�0�ǯy�9#��B
S�&��/H }�M�v�l��w#��l�<�������v/�)���v��y)�Q��jޕ�s����Xwc'��e�Z_��#�S��O��:e��2����u�e�uS��S�ٕ�ݍ�_��9�� �o3��0v�#������y:���D���f��aG�&gd��B�u���$&����Jeg�`fw�WK=�b��HT,���j�K�|��E�U��;J�v�zG!}���DklmAY��f�X�H�gZ��n���w�V��+���K'oY�3�o��3���*�INl'�f��\e,qTȥ3��/�G���d�p��F Q(�j�I�U����f���5ST�&�ìqU��1�B�XlxVHYEB     400     140�@G?0��u�l�It<�8�0�yqͶ��̳�̔*�5E�D���&ȇ?�p�4�U�ܨ��U�=�I�v�0}��V�w h��E�f�vk�q����%	0�
~qy�^?5�;"@�X�cW�6�2��G����F��ڇ������&E�u�pG���Q#<O9S2�o{v�hҡ�,���w������{�DTKsiaZ�tjcO\Ze�7�a�H�����f1�9Na(CkK���Xʔg���;B��Jr�jF���2j˼�W�	���[���G�����{��T������jr�����XlxVHYEB     400     170�	�Y`R��r��{_��Vb�71x�+CIY��dJR��R����c��G��o%�"��h�k��)�|���^_�x�A& �L���@�A��C�����u��ř�� ���\R�[e�@�o��TѨ�vJ�Z�|�H�����Ӭ�����6��(��D��T�}��&��TQ���������;�b����N�n�ćwz#vLY|LD0�q́7Đ�:���O\����$EHe0�;}�=f!n/_��V�ao�Z榕v��$3�[��Ms��25AS;��_�w���	c#��Aȹ�%<R�"Wr0~*�� �x�Ό0xA%�F�)�hgތ
�[��0��{��B	�g� j9�XlxVHYEB     170      d06h|ےIZ1N�.�W�`˰�?��?��K$Q˟�V�Ţ&��u��|� �&�Ơ.��=J� ¨Y�� �G\2gW�_��IYUb8D#0H��8������qs����w1������&��ByA<���w�~k��%��Q�לʔM��!�,�?\[���p���]gb�]�j��С���N��a?��-/��@WL F�f�W� 