`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
GwkQ4iYCzbNcd76q3dBNkM2SRaPLt8meyJ693bsGNhEPMfFkFt0i3SwUSuSVhe4Z6wcLTsy+FaH1
mjzvzO5GQV8yYCA/Ers84fe+3b2fJgk/ob6QyQ5z2LZKSjxB5/xKzFBxf1S0m5Peqv6w7yA9dnE2
WXCIox+MNdtuHv7cPKLzwF1vEoy/pRZSbxg9K7NayyRx5Q6oKpIW5r341KTkseT5P/mZQV1B7nBn
z6A7bTYVzuy5UJWC3PBwvEmzmxaFzD4+ONS69I5SWbAwH8N5IWcjEi2kKE0p4ZbgminhD2ZyzPKE
Ci+va6fe+x0j4we1FOjTx1fTOSU7YY9WEEDdQ90Z3DwdUT/rhJ97dKK8jFuoXKrhos6EqeGi6lbD
dJZICas6H2hdmTQaFIeolu0HAJ1pPsQ/g5FETtVWpHUeyXZRVY61xDEOqwe2LOnNtUP2AX5GvcdG
idd/uRG50Bih0cs90GBLyoW7VnauH4UVzjgkiOrfHp+GCrJccNTaMokFZ1Bdq2wXYVsPah1o2cSs
JdDPnLzJVqpL4Bson32teMKBGu0KH3a51vxNU5xOc8FKTJBH+WTe+RbpTZTX2qqkPg2Ub8C4wQEO
ccnPUxh3bzyUZaF9yse61ttjAEVa4DNQJXi8bv4c0kR2uwCFesmWzZX/GQYZXfABtDpHjSV0S5PE
OgYhIcnyRVhOR5TWlgdoMZ+o4SnWbybzXlJh1MoKplo8N790sLKzxvKFHogtG7LGzKbS7wga8D2s
kMUNrfy2altJ4hXEuGO+jSE96aIDazLD4UsgVZYER/TmLkNR6EW2XB5cWGyV6jR2D5b0ioZogfj0
U2kYFeGInVC17EBS2xaUPdUredCpCoiFGep9FEBaPBFMIEiQZMaqaxQ6BpJgWq43vF1KfjrCafp7
1eitoQD1OO17Ioo3ryY8ZtRyJbtEmf4fBdUdEU1q3TDNEfIfs2WAxxwCEiMz+4KcxtE841QHIveA
VZoIW678FAU5zQonThSYaeNr2Kyfy3weVCC3peVYlyZnsq8JdBBC8HH0kS4l96Cdt8Lk8q+QAQHo
9BOvljBjNRdsz2L/Kc7xvExtYkaWKSNx7xT//LHQgd681smBRg/p87JFVoBPvWgMvH0+xtiKw5oM
+dvpWLYHEp6SqE0Y32KdJD3XWsYpJeDACpcLszJSjiszNVZLDa+ndv2eoCYPCZ/Q0+3H6c6tcT8c
WkuA05yLwVJV611VzcKiO0NmdYqlWMfl0dm+fQcYAmm3YX2cNytBlV65e8UINF53vNudGXqS/L/Q
1IF99b3C+3sCrtcR4uJ6UZspeSlZxlPQzvnWqhBLJTsKc9ijJaDuP9xnCENw8b08LXQN7fuMjg/P
wABw5yCxVo/igZSYVqJqxW9MIeCFtB1fBjmROjltqGIT4UBg4GGmAUc8t7bYVWSyze/ZnqP7Yv5C
h64Q7b2B+5Hwc2FCYb1ASDVAqc18rjRG6Q97OQocv8aQpyMZKt8iVDLg+ssZhrmyQAlO1xH6D8bA
Az4d0V3jHB+WTm7XJUg+X9UIGnYyCwj1b7pPmwvmWw+8XIJvple4HRKTPZBUrKPadHa7yYrIx6Bg
6+bjvF5yOaELiG72TH0w4LO8jlWCSlHvPfNhx1vRSr/eigS06X33sj5MTOdtUA5nLKZhBvCOQdKV
dGOH6PfWoC1VUkeSzfm4G3XfLeQwpK1NDMAWUYCBylHtfeaO5jMD+1fuFMT+jJzTAUTOIH1PvlMx
4S59hmSNo5dkZtMgg9mEZGB+PLoxWXnUqFFgKPIxvQTwRfV6wD3IWCxjcmB20FHYq/Jb2VVO0h1M
TCjWR8VB4cCZwZ43SsCvpvH8+00Q7xmwfOwfQL9R8+7flh2cnpUL9TgkNwa4bluiBfF2nV54sNDF
nwztrgVnAlFo9Cepx8yyxxqleOR5vj8aBVOpXHr6OHUN89HFNn9+dbKVC83besYTkCnLLBo77hMr
jA0PQYz6+wLRJxzyHK0RyFdMVPeF0FAE9grLMosRVAfvAv+PStlTBJZKOMSVwPwoiwoaxXz/dwfk
2lNtVBx2HSloWT54qMd6WGJdqatEuDDLWFU8kV+bgKQFeUaUFJ2vfJvVI/NI0K0cAGnRGpCcHIhD
FOJxX5vosUK6yVjlbVZV3c6Dzy8tSO/LERQnnjEwylv2pQY88Y7FLS1+nB8/n0xK6WltyFAt3Hbm
C8dEGpERbNvTMfhXVO8wGTtnsztf9G/6OsAHhttxID7mEOyLrdAJojy4wJmL5w9aVsTkdLF7y0J3
1I1Drrom3CnOlgl3oawTo7I5XeBV3eJR3xx5txsIuwcl7scGER8I/BLPzt3vfXYsKz+vhozF4KCg
nO0gCkkVJsfpydyxPEW1D26pyrmahR/zUQCwitgRzuFCujeVM9OADmC0ZQbbVQaJLNpF6tjoguCQ
cFHGFHJszAUe1AQANM7KApkoITLHtCpM0xbz/ywPHqNah4Nzn471Bzi9s5zku6I5z0L1ZWxN0enc
Q642WP3he7dU4Ie3xdrsc35OIIGr9loY2s9vzPrn9OWvWooErivC8VM8Z1+WN4mh0+CKdNKzzgf0
b/sRllGyE6Vb+SNeNaqlIkIvwbMKMoou8K2Fnq2y99S82KG8B395egt1IPwQErJDXu1qL2QatwAb
J05FP5eQmwdtVtG9wBN+hYZnHkl6JA6YYDopmW5VxSjadBNOzllSZg72Wc7DvDpQtwB2aDCQPScu
v3vQUKOfIGUcEAvENzL1+MJA43a+CXb2ofNN+SAlHIlmrG1EXxpPaondpOPthdlHYUTZzgzgJ+gP
vP09IyXcdbZ2dpWv+v4fAhSoPc4CkmqZ8zdCw8iZorN4mpfdRkcodytkmy82dqKtalDoCnq6CJ2R
oIrNv1+GH3uehn0L5f/ogpYsyrXExNBLmECM4onW5vzJMVPIoqBhWQV/tkC9TTkkD0V5GscplZG2
VTyQ3L3O4GwyXHmcEssqo0YFrSd9ChP3+Av3r3WXtPh599ymljHjAaEr3CaQrE2vU1PVipLbU5KM
dtSGU0ROCt0pgtn7NkD3SayPnh+Ky5GyMbQIeJ1eeqtY7uzj3Cw5wr9l9u8Yk/rdVRYSDc7z5shL
fmwewh/5mkpsO5HI2qqZblyabmLd7Jf4G4xDIk6JWpqNw850zHPB2le4s1KDk/L0ur8yTyka20+n
UnT5/q2iwWFtQPsFJY2eidtXKjL4/x06+mvOkcQRom1hc8/v7X5+hF6rciojknqs2YawkjThGNMs
oIgcHFAyhB4Y0RJquHSVUXty7CTl1Ki4i/vl9j3cIxC0nGx+ARdBPjsiPYSu+peWCRdHYxw/ypd1
oyVgGM2IA7hl2jq5D7IYyECgMBhvpxhXcNgFDme5GjhhXs2jIkwwIiqPLfNp+F2EsJ0VKQhCHFD5
Y5HaJWV12Xja3bRA2R6o11XXm6SB1IH42YPHVEPFgsEvxdxkg+S7Fm4B4BodPZRxDDtSx3UaEKQe
Vm0jJx+5myjMlKF1t0al+tkjObDs+E0c0JnMkNAhQ124qZEtyIZTOVGVbJDDqnlOn7eivhirrvvG
32veT2PjgsxEYfxaxl6DyTsdrqIj3cySDbgTl/0G6HpPt1FthsqyW790JGn6NpEff9ucG9iN96yU
B4CsRdZp5tCKZxuqcpyc6dU5Gf9rmEIi98+DyYPaXaYqnukV/yaLTpRgSILuHdJHSXbpy2ycCdXp
d6kQyOAelVorc090qJb7vcp8Pcm/IicXwgVCgfJEO8HV2a0Kim7wvZlwPInoMOiD95whmhub4Y9V
tvLJhYrBBC/+c4Xd+esdI0zepFhLILJML7DSSY7YOC/AfeB/GblBuci3dldS19f4maTPP/u3piS+
8iIcjPXYQcJeT2sI4hMsIZVSFOfbdAWBzOO66R2Junrh0kHKOuJX0YYNnxclIc4RbpQKBa/SP9U7
vHTfo45893lF+8SEHkgfXSHQVRbTVY8WC0nLY+1ANzN2V7bvzmXR0cesPauyH34Ohafzz6Gea58M
BlxuHGvCcGjBtjnWbaqnTtBd/Wev5a3X/zkXhuTs4KjdEtfE3uKCi2zfxwKGVBIROSjHkuaQR2ls
XOD0k7g00FeeJ4b0F3r7HfaeTUbllZwzJj9UxnoKL1DzCaORNzAdDC25Gh71sEgGFx86+3xltVwf
80kTAJbUDZ21OQi2qVGQzkRsVWQAQAOK72XZynUNobXRlV/UjWhH1n+ZAHCs9WQOdCQQvxG4FVfT
K2q5uU+uFB0F46D+NB6QvnNfFJ03t+3nURtSkY28+7pt9gXERecYEfh5FzLHUmWSqDbRcnh7NwoT
AQyhoRgFqOCkM0bJlY1n10bdLHMMse/r8XAEUms5qPwfFk1n0rtxU4u96V7W3zIkKXNsDWYeg6sR
s3aT5z95ostpQN+MEhVxKuhI2BJUoWn8dJJZVzIN46jMbOyQBa5MC9VIJdsaATBi00UBcW5FVE3i
FNYSgjQ5ELWNPEAZp12K54GkBcI1Axi9yb8UTwwD0+/BcejYfsd2taGIZJOv8KsEGkHHtUhHH0zS
bFLXakTUFvT50x0bEd0dIO5DGg5xvGZLm2x1kP5x2TSCVNzaVGrGjcwZkTN3JElU2TNr9pvffHOt
6bWSnYlrvsMIAuYEzLCH+cLFnjmTVAjyrqD9ulCqcs4wD1VpIlaYX0esx4QjsakdbQGupmOlnMCO
SWqZItElFBBnB9tAAyAvn4G07rZT96/nFRzalD9PfI7gN2Mvc8oxhSkFc9IyA5U3i7HHMVH3Rdwf
33UJfXYvGEG06LBQxo4t4iDLHgZsotRW6yuOv6I86aJGFpL5iPv4DuFUzmbQVTE88IPq33JQYgND
3HOnCrWo8cHot1rKenNmyewZRYXeEk0kMBSFRn1Hr4H5X4AYTb7qszA2JMwDWaj3wVjxSwuxrumE
alfZj3BNgkDTvrqKG/86MSEsRI8SU6EWWMAkVXd2tH51XGhPMxh11eLxwSLH7d42LAYEQukYwtZf
t60SqOz1S5HqxsEOD0c2b7iAY1QvqyLXRLIs5M0wPcsuU0JthpduibFogMiXn+NuOVH3nNPW/7fR
zd7xkonTcO4vxWJlcjTB9uxvADmxYi08krvQf7YTvbR12iIZQm2Z/MrhyVbmhpMOu7qlxl6DxbPL
uENYdEhA+lrq+Ixrr3ZCUUBdNWsmVOOHr7yMSzAuVa1f1ncKnMfxmwya/DBZq33OIRyXPll/ro4i
TsGTLNMBaKCcOySZaf4oBpUCD+k99RtS/nQDh2xDcNNaG/Qsu6aKntuQpkIC8OYVGk0lARdxM3na
bwmszNr/ytl9OIaCZPM9ev1mCYD4IvG1b5groMvxzxKg7S8JYIOVThKH1Jg13W1AnDbxpA9InWBS
0yxti2vTpqkhn3jwKMcWF3cQ69E5nyPDj7okRHNWTT925QbsStI/TWe5FvUjnT/tlibUu7T0ad7t
rsebz0yxZqS458LCdPgbwhL4O4TIidekmEwgUkZtF11A1V/JBDST5tPHEBblUiSHcsLWZw0pAGZr
kMx0FfnPK1KNT5cLO7Ui9bacbiNzl5SFJYaXdyjH/ao/KiUsQXUN0zuPKIvWLrLT/CvUzipXHXl5
k/ZuyVUny8wmbt8mLsLkpSxmiVeO91NUhVJLDRfFxPAchjEGndCYFb5idvn5NMjmx2n/murAYQ96
N3hM9K1lchtC3of6VYmB4Kz0dwGLZA13XqrA3TxlbyvkBiydw6Vv0PxIWuV59MnO5HYR5OpkMs2u
1rKPT+qWh2eKKWnabAOdIclpMK0P2TvQ23z7y7MXMweKoIzPxr04RjPf7LUTk0g2K3NKfcuyGkYZ
t5WoW15tqeXbO0BKkd3V6COPk7BYiIZQu6hUraCcQ8a6ToBDPv3sk9Z5NRgoZHhNcYB1G/eQQquy
kNSTrKwz3Rdk9djGHca12nNlWmGrfGQoO8iqbrLCgh9OgdDCEA7ebeZNDp5mFjK26JdzEL+Z3BDB
E7hbTjNuGdbTHY16U2uMZdU8G1eiWkqYymFhQo421+YI0fm9rw47iRGK9ER1aHodJ17SQI8wIiUX
eJHUoKp0ZMgQeQz5/ZMCmqfQ1fBBK8IVbpMdIa27i+s9j0SUdcwXBc8m4Xg12AKmtLh/B4m48/cf
WTQMaoBuwl7niNUFspcM5CwnSnCMoa1Tv4UVUMNGfWh9QaQa9fEpoodgXGrFqdGqIpCh8nmuU56L
pOz/W0jdUeYMv1iU6F9EVGqe8zMxfTV0v65ovuT30meorPI8aVpMF9l4Tapa79oIvGheLSPvBiiV
BHH83jwmDbwAyRZrwsftxE6ZKOurZQsgRQEpLX/FMT3p0DFQetS934aYognPlEd+N1T0hXZ+tFuA
IkSOi63n/DwOCnmMxFv17pViZZWsCpxuzJAns+cm9ui6yGEbVhMX97K/a+hJIAjIE7ZUcgpuAKZn
EjyY996mhxeQmMLizm/9EVSau+pU0KE0mEhlp8qyhlYoanM1fKg+XEnFcoHmtFZVVcSvSUn9XLfz
/PNJPcwWbyd8E3X3uo3mrYRfcxwAQDtHypZf7M5xevoa0LrmxHFcLHa4PFZSeOiPS4OKTc4YkR97
RgdPAFMFUIl2TpSy8GU2eEQPsWn7PyamRqeuNhwt/p2LB7t/+ihSq5CUlt+S0oJRzRx7041wK1LE
1q+ZxGnebCv5uLc5VcHPMD59egarxdVDwsdzo86cJINKLk/gfbii4RA5d5we54HW8WScuGkSVzTX
SAzbTA49gAzPFxJQNWPmTRWuIAKoDYuDjnS8aeBUHtGo2kAQGyOvXIwlkqnWVyTYcLE3Z8ubSH6n
Uru6psuyer12gJTOkysNAJ+ocRbT1w4B21qJkujKjMu8EJhZ8Alpgnem7Pr8E+jI/ewCNO8vPGNv
2s+4uQiI/6RqrlOp3t4C8gK4qRGpRN14OxoefMut4C5ifHqpBzcgjeHbEyB+IxtwOmQTMLc3jgJO
fZhBWe2Fg4EatlYQGmrS5LdjyOJRNKiSasar+Qmb4UtI3tco74BtOJTgC3OFii/X0rBTWeDKcSyN
dBo7JUWWU+DuNB8T3AvWg7iL5homx7GySKYzqhwfxjqtcBTepSv+nwUUmxlo5tomSqsDlk1USDJ1
qHlVckvLFxqIUWrJ5TpcFAigV4Cq4tWBUGWSNMq+UaCg9+gP1d7Ak/MQq1TJJcumJVUTLKtWDm/X
dEzZoxbcdG/NxwKk5A5MUtkSHp6W4VrNzOTroJxAL4RokZJyQ7SFQWTM826p7D/5Mk977zvUKyOZ
rtzVtjTau/dmLNAIZYijOBGQsF9xH5myPngGcwbnxH42wd2fGMZhHGsWgWgZLQF6IsxJSgGHqOX0
dGslfLK0lMhdc818H5UjV8F7RL090+JOSk8AqUdXNmLBax0jK4/z1VNgbksCSgkyzUMDkALi3Q+U
/amVTiuMH09/EP9KPmQpgZ1GZvUaz63QUz0czOgHNNeR7+BLbz9AorpilRvNC+RrCIWVskI32Lq+
vdmO3ztCHtJwbmk8JaknYyTiKyY+QVq3y1fKoCpDCxFlTLRswJqYaLTfm46+6j1Q5KNGVNWTWB4s
qrm8Q07CMMTKUB5GJIyn+HJS2OS5mhbA3vV6IYLEFVcfF6GUoOkK3Rt8mgc5fFC1fzTkaFEY5eAi
Xia9lARZUnrgQLd0PcaOrSPz0OHesatzBq7dKA67KpLHjf+f22JXl6XuhRqH2oBN1daxeCCrlPSC
x+QHGXDJQO5suOJ4NVfIHKR63o2531tk/DUeJ5yEmg5be95xTbZNHTtFf7VjMqFoTL2mZseySdzL
Wxlio9RUb2NC22W8gRj/MRyQpj3y6ylavy+y/8c/Yd8jFpSyfQuOCMryKbKJ01LeYOTcImkkxQUf
Y7I6b7T8OWQGwIH6aHcPZcLbtDHf/1w48kzOFc/S/++NxS5lreb9ec9h8cj5Qa6W6x+qoFPn63EO
Juw+9gPFOowQ5HZnVCZPskOLZeaw5++9fuoH2eQEKPztb+HSh08rrxIk74o3w/wzCwtu0a8/C65K
A5nJgHkn9Ns5SjgQBrUGtcYkgjwerdUH6yNcduwqdYzTm+m7oa0M/Z5O6nL/wQEgCMUSuwDbG7ZP
xcPwxkib2HrIISntispS05EK6q9nmK54kyt/uJwCcH0kgR5CLO/ncksmxXgxsDVi9gfOOLzQhEno
JEhUdIYnSSMB+qzY+nHUEKKGLvLEY+oIB+ij8lx+QnHnmS6DD5s1vYNjCrQjT3DWSnkPFpKDC5el
uJbXT/OlpZMsFj8JegMYDI7BfWm9WQDKKm2N7M3v7IY+hxCQNBvWAT3NF8t2Sqkdqp1E0KredbLi
an9+0eFhzlKxiB8crm0J8ICOtc63FB1Mx3U46ThIalVvOAmPHoKsGsQZqEWl54H1/zTXzLVEy8lo
91QRigFRtpGlipjCpXfQQEulry0lgJDGMzJoLJUUzSg3club4kqS/ei0Y/UB0+uw1w3uPerz4DWF
26ZhXqbNIffvLwAwol5hEA==
`protect end_protected
