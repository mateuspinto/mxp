`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3088)
`protect data_block
0USWSUGxovGsyBJteYpEoXjW4Bbzd/GZ+16uHdoRQNgJwIQ3HywEcNH8JgLlUunxVcpU/vEgcZ5G
F8yJs2/fjnQ5cu8n8IlpXKCEmrYGcpL4u71759qKRm3YPpJjDeJ1xTd27HWLCQb0Apt9vtB5elkT
s+tu8WHFrFCSxNJ6eYx+whttPO6QUAMW6sW3KQyaSJpb+tkgwtr2vs7Hr3nAqnTwJx9FCSeGt8KO
uNr1pcFB3L76XmZ/zRqR2rZP7j1Mr3vXadGnRbkdjfApZWVslgEgGGlCdcwOSTBezJ4VOpRXDk19
Wi7u4qckDKglnTysv0vKC9kKRr2RyYmr5JoPx4+dWqi4Jt9q0ocus7ar3QS1ZYP4uyVaQ7hfCIc3
UlUR+ViKsAFDiGpBcrGrwS2Dykd/KPtSifGUQD5SSrSp8LuGlcO6Z3JT9K2w7nYcta+1F81gnRMZ
cDEnttJ2ovZWIOQZCIdAMAQWYejEQY0ixC6xzpVPaxv3Ym3lnKMffzcB59Lr+tZ5K7dlpYzsropa
bC6H5R6VNo3ZZc1Rkxh6VTl13Qq6VRK8FY2JgL6f09X7LSuPjrVlia9sU1FGLZhZwE3rFM741Dhr
oZyq2OZxg/FujbrDorr9S7tkTfQLy8cafeNNsywWFXjHW25zfg0axbBLaFek88RRn0dq+6cj0MGG
wS6qSQ9BZCh7HPNLRb9GSd4O/yECinngibErivnVj2Ei5XTrPbdkOD4tBYXwBUgXVRg9sYFRQpTJ
+LTpacGiBFwOd60g69XN9fiFJ6u3tcsW9dUTaVG3lJ69c0+f1Ykhy4dm7vrdnrxauKSrfOSY8QmQ
KULS6T0v8LIUBLGcGhiXnPfuUnb2/5MNZvOcIrBTUKodpLn3333t37SpkMr14onYH9TWdJexvSwn
ngdA3TDXbEjJ+4CpMJMmEHFwRLUQKA/FRFKy+eKGgixX0Ua8cPTb1DWDJKlv/sNHyLhaNYWZnBLG
HtB3l3YbfjJK8efi3BPPqm0B2BH+x/zyFBG1ODfJfXBjwso0P76hvQM6gRdJ/2UuWC/XzRjR4Ncw
fd8sYH3diSpH6hFnBekvpKUBz21FDismSjEJq433+6J6wZQiX05w9Q9Lx2Ba8A8Xcfyvzrpk+Gql
+JyNccymDl6dSUWTEWBu6726s/2DJgwCYwGsfcecENVSfsqF2n45kBjx2tODmiXQqB6OIjL6rLp0
2xwwCFF8yxsg76qMhRikBjQsBfGwNkgONlWVWEdWOuBCXSp3j+Ap7SsyuHbEegWKDzrFtQoEEx9x
MA2fQOVJlpAYKGjAQ+ciRi3FRR6PZesKOxqBU6IHW3qj/ncjtOiuG4REiQqwWJRJ0A2w/Su8Prq8
SbaBbfTjaF5wcuSJZyuWMrzJrqro18cdoYxU6lGGinHoNUsO4EFI6DYYnrWcSYBTTp5D9EuWQ3Ji
QBe2EXYQwBvIS5QY1rA55pjesjts2IGPeLrSc34KUc82X70eFI9LZkIbxNcnw3X5kvmETmwyTMya
tX9vcMuiRkgraS+IcxVBMu0gEQ47RifUrUYd+l6M0XYXYcg2LB0UE4gzDeqH1kJoffBcCyLKzMIV
7FnWuWgmYIW0JV54x9TP3Ojg2/2j09sKd+35VoY2Va6i6dsBAEtYOp6pPUhlCiYsBIL19VnMrk+Z
xB/YCMUS7EH/+fZThFYTg7Aqf5crRjwtR69jtRlysDmztfCzNgAcFk/cW2xU+H1kHxuTz0CpnZ9n
zxYNFSeJkiTTACqz9Zf5KPcZzGTZPWxK3hPlETYmwnHqri+WUPerzMwNMMuO4Ttyxe85cAzg4lWu
y/apYvhWch9G5zrxxfank4nRDibjZ4QMccG6zf+vRlCTSzEmXL92AM4ctNDNKJKDsELi/3zt7Jgo
egkPKR/xUDU0TM7OWgapA4ztVHNf3Oueje3yXei+u9Lkc4f0LkPK1w8nDImSjw0B0gCQS0/tSSJR
g0oSohgghZhs3zY2pO1U0wFMeUNHlUF1l4EgFwUboQhiONzUY5yNPA/HpkVzuddKMOtjYsuqpcrT
s1oOcbfzTyIrGJJCztboqKUbuvJX/9+9dV7SSZt0i5J9GgwuiVlVsXsRKHWNWMAxFXU+BGrvLyJj
NDMf1hnE1zSTwmGXrwMT0ebSYskRtn+x9P661BOtEHeiyz/IJVT96Nne6DBfM6+YjKgb3qs2JZfe
vIlh/FqJAqmglsvhxGBPSZU57h82rEjDrWfEw8kYn2gFd2WoNaZnOt+x4DCDsu6XHGKB9uO24x5d
s9MqDAo/78kT4KwcVvoQ26iCdAwtq5zOmmc3u2RuxzyBEUozRFh2w0BafFkt6p9q91ZrADn0xnqd
YID5NSf38oDOSocCMNZ8b/cIaRzGGCLBHP1leYi6LRk1Y8SDLtsgPxt7TbW/9LQRAXrcMgy9SBAe
HqfWMf1SKKHVpAP9TYC1ImI82eQF8nno6c9yVfxyld3re7ofXYwIEPE/mo/vMCucCmub7xJJfXkY
Yistq8nw+1pubW+4/tCWhLZPg1p2sDThgPZz/dyEqUBn1O+ypITSz42obMOlqL5slH/Bco/c5akR
PdGbReU/4zWIkZcU5mSyLbFNJ8Hg1TD1+F+Hks2xQnCmMIUJTPBMlPrUfjtK1RrZ7mL73krFkdvp
KHzRijcfbXgdTX90FpO9YoEg5FH7l8TmTl3I5otqqGdVY3HH5Ua2J3KomSIVWviDrIXqURkggDoR
IxAsXMPeMwJdSDE20pQX8tTTiiZa0a4QZ5Pz2WKP7c6FZIQnHn/tTjdZiaoMB754XXsdQGXP3ntK
kV47jvIoiwJuDkuj6gcGTiQbibxUVS35RfZovmFBFY8MQtF2GzEf/ZKsrqpyIPyNsLvOsvp48UvO
mlh9J+dCNYM3hWWVcOJ84GfSf+iONXGUaNkHiyE54wXnCd7qwopnEGYnl/uh756vr76JDGNgSW6x
1UOoeGmEaCxeCJ8CMoTuP3/sZRYhsAYNknaljYyCE7h7oe5uNHZPceqpgQYoD7HXNQiqy8t5borD
02U/nvW6Tw8Esou9dfZx5jcF8oGEc/tKfyY/mf5H3QiK6Plw2ah/VU04LUAlVTdf7DdvG0bxpkvY
qi6KEWxfoqgVI703qlsROkNNyxxqRixtfbyOKDw/62oveK9ne7fyVUnnVXCgS7dJtxHjTdRaiXaf
FOpzijCWV7TTDsvRCt87fvfEAcuW5fsYCtE7o0PJBFfqQSwyoRWzwsLbVCnwJixexaLH8+XuXT14
wpnKu1QMRQH6tVSTAGt231eIpfGB9mDgYzMOYZfYr1Vt6r6chOh47PsRzAw8tn+DDUtGMTZIIvms
njmRhtgg/L5fFP4nrliamRvwrp4JK/iSNz+FXQEr895CN+zc1zDWHsOtOdlqHAYww57V5h+9E9fB
2MGw+2YnNf0r1WiRs0Iz8jQR8XXejY+9/j7mOfrO4KWw3y9QXMZsJLMV4CmvSm4KRAoDGT+Z2OkI
cE3o2HCa7TgGgl+CYWg4j+BwaD14JAb5aXCvBSAAuStpDljjHIP6+xXJl4ctK0wOIOeHWfVgjxmY
3EPp+Mb1P6DvJL0W2YvMHoaYEkB0nUWR6hERNmCL2XNBUc6yvlSsbQmEA+W5HwodtSsF7jMub4ab
LnVZe01gQ4UO73IMwGL8kgxkW5mZr8n7w585FRcPRP04ysoa0PP7+YO9tN8y2AxN1pHNITzevLNp
950Lj81tE0uMPfqVe3HHxswXpQM/xqZ2085Ie8a+aCvqqLSp9ln3rqp9Ii9VXT+r2udnvBRYNC9u
BZn6jMDtLwoHNValXCXlGHsThyK+PztRbqf96TvWZuFWamNw/QURrlJQTCzRuR6Nh3sHGWN/9JTl
9BjVcm69IofWjy+DcJVuck4bTJlKfXP3gWdJg5PBuK/WRoSSY0ZqPelxdcS5PlTrm3bmLRRoaXgk
++vFI+GTvuSoEfyZ3PfmMXtTg4B4mDdWD9/wGIqv2bC4/7DeefNw8f9hz3B0xJ0AKLQC83jCT3Vj
nmjLASeie1FiQShJciXBIerU+gS3AiF+4yrirW+N3cTnxVdAUU/BWGKFngF/lFGi9sUOVJlSJoY1
kLPg6dac3vx71Q==
`protect end_protected
