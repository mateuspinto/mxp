XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��2aL8��\�(u� Hȍ���:\R���P��u:Rhz8�sĆ�U�jM!ٜ�26��5k������H���#��5켲c��xu�ފ~�|>7�0p�aVe�~A�ϣDA.��c��k��Ot���	�[/�O�&�KD=3��Z�Bm��a
��H�ԂL��ۈVf�)u�l�Qg[ù�4�h�\K�vc��k��*f�v�F�4i	�H��Vp���5���������F`�y�>X�B�0�+�\rP�t�)!X�����^�[����`�s�}W|��omMK�w�E.�m�m
��P���%IP^۫`"|��5Y#�`!�b-̚�	8�P�uZQ�:�^��6�ցe����0o�9V�?��_Y�����S�o_&�yT۠�Ʃ1��+_��@���pV�%�:nzYE��	�+g��	6{&��lK���4Uun��r���d����5���?�����F�Z5��� ���j�
R�"��J��$p��	�\y�'��pq�(�J�-`�G��8"�L�f��ܪ~)��R������|���vX����H�Kᇚ��B �l	`ܤ6**�)�p#�	/<�&��ԆG��l�1�NEw�L�;��dM��d��?�� u�����!��~��7S .�*'�ɏO����F;��e
Br�����Cfх���*7h(�1����F�'�(%�[v�k�v�4�j�H5~CQ�>Q���t���XlxVHYEB     400     180��5z�� �q0�Ūoc_��ѯ/%�S��,4�5~�sɃ:�޹Ⴟo�%%K�	hY��O.�xZIc@p�d�\թ����a�v�����FH����m��,�W����;�P����BA�PMyb��+&�Gz���o�g�Xͺ�~Y���]�.�K��3����]�8.��˳� ÿm𠜃��n~S�5��R��So����ch>�'N�lI��?.=b!$D�w�ʷ�f3�|���� 3��,
�2Q^�|%8!@F
��-��F>k�7'�s�c�Z�Ǒz��"��ж�^c�tH/�X(�pOY2'��!Fv����j�M�%x���7�/���Ϧ���8籲�;�2�`�"�ʥ����ÍböXlxVHYEB     400     160/
f����/�T�c�rzX����3�����
3��W4r��P�.L����m%�^�2�ō)Uk(�������:�kյ�5��j�l�+�����欇�ZY���� ��Pb.�қ(�T:�U5�翻��M�ea�Q��$E���)7zz� �Z�Ur�B����MT��S-��X���	���3�e� ������6��K�&y�3!���W�H�kz�3C�')��$4Li=��c�H�/L��-�9�?꟥����`�ᄔ��.?>.t���9$g{�1A��)���M%*�_��6���4Е; o�����;s��W�n�m����nc9tq���>nh���%XlxVHYEB     400      a0%.�ƣ������=��d�:�9؉�V"�B�����/Az�<�T�,���fN�Im<q�kk�Wø�	_�Mp��&X>/��Gw$.�Jۑ�>)=�ѐet���3�#s����J��NUٝOZ->}M�������7%�]+ͩr�����3���ϔ��XlxVHYEB     400     120p? l9��X3�G�J[[݄�Ӽ��<�c�T4���6{�(�H�48f�T%�f��ϙ����n#<BMmO��~����4b^jD�M�j��#� ��Q`����$�,G�1Y!D�Q#v^mP�پ�_c�`�qW_L\�:���D�#�Y/�l@t=M�%��VQ��J[]���8#(6Ѓ��$�V2v�
����^z��m�|{˲l�w�2)�+J4yQ$�r+{
CM����!�#�����ؓaǚ}@舴\ ��ސ.�H�09��{�FB�6qJ�������޿��XlxVHYEB     400     110��[joߪ�~m������ʞ���g�Qα��E�Ɩ/�,d�C�.��wǜd�)B?RH���P�]�"=2�}@�Ԕ��)4	Ȓ��ƌ��٫Ë'��X�/��l��|���AvZ����#Z��^�n�qW�P*�{��Df�ͺ���(2�a�"Z�p���7� N�XR"�`B!?��.�����.$���gT:�"Uj���1n�F��Y`I](�`])CG9{�����q�%��3N:�8�Ho5�Z���[jK<��OJgXlxVHYEB     400     130�-P=Nǲ�Aw���2{�>#sh+ �]HT��Q ��~ZQի�!;����j)�����
�u� �¨9� Vm`�WJ���Y{�M7pW.�ſ#b�8a��>mf�A��������)�+mgީ�0�^�� �����ܝ����X�v��<���Xgق	q<�zz_u�gzeu��5�W�k��E9f�'	'g'
O���d���8�����*���mrPښi�$E�<,���fN<,7Q;Q7%A�.oa�TVv��v�?D���z�X�E^n�_r+�NPm��}�-�����L�e|XlxVHYEB     400     130>˻L�ߞع�L���߳��M>`|]8��>�����m���=	B�Ɔj�������h\��<�u���-���d�(��@�t�K?�r_a;k�����q�F��Ï~a��F��fjlF�.e�e�����)�X�Mم���:<���M��w�����ͨ(r8��6Vg�u2�|���4�so�xڒl�����o�`Q@�Z0���^ �`Tl�^y�p�_�B�B��Ew�N�5b�C`�Z>�0,˯�8o���7���``vD*eo4���
X����ʣs����1��N� XlxVHYEB     400     120�|�b��M��š�4���Z(���X;X�=��!w���{9���a�Y���i ����p�#z��o�*���:T+�\y��i�2E,���}��(7S�����KUm�B���ឣ��uG+��+��\��#.�!ysB^w�;y����Θ*�F#���w�#TQW(�`l6�j D�����B-O���j.R����n��}�JN���T�Wa:��qPm򲍂9J�Vsi����'O�q؋�Lv,i�x�H+����x#|@�V,�p�@�#����B9��XlxVHYEB     3a6     180H��!'��z� -�Q��F2q[�)e�0�)0���6)/���j��)�.�k��7�O�t��ܠA�y��22eUd��gDb��Rk��8,�������j��H_<��~�I^z��|�z��j������l�v�*���S�����GR�LHt],�������S�x�E��Wc���qUyujv�4�|àާ�&�� @-Nr:n]WcW�)��&�^�#R�?�y�u��<
B(��3�p�Y؞N���tms+(\L��&cF����p����("0k��i%��O=Rj��
`�7��`��������&Խ��b�KN��(�Y�g��y�o�����L�l�2
�ԩB&Ob�2@��8����x����2ꕇ`��;�Bn|�Q=