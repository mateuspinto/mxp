`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
gSNcb+B6t7GN7GuV8VFQz+lvxYR9aDzRHTtJmnzYcJOiq164tH+/FKaYLafRnuMlo6c7VbswuHyv
7r6cQnYW1isnhmm0NRV7uuMIy4UkugP3RiD5EYsUMTyo2MFrPjI0+NCx4Fr9axnwhipB+yNixTN2
TF50qwXCmDtfeKIn0S54HRYZR/Fwwv4ceWIqNjE4JMkMYykbswo845/UKL39g5+afr+VDH6X9RVo
8tX3nNnL1Q9CnlD285wv26exNNvi9pf5xZHyzDMjUYg8I5XLa6petg7dnWj5BHz/yxzd9Xlq3q7L
rqk7QsnzMXqQATUKCR8W0OzU8WqJZK9msFMlQA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="k7nEJs2uOqvR9E70Gmc799QDm5489mwfI0usGgDHaVQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14880)
`protect data_block
93ysQJqMcYmoMcLj+ZS7s197JggpnVjM0oCJb1OLO7y4dveNKfc4U3GQa3Mqebm9/W4WQJckgmmW
EGnxAcV64p/oW0PUVLb7y3o7n4w99HgwZ4upbpzWftC00036SQCIlYzLEhClnUClYIrPHPzzRo1J
YxwXw0yBw/4kJvSZy3mBoF/Z8q3SxnhzYaEfa2DPbgvjrK0qjWk30AwjLu4lZA+gg93JcM18k4f0
L0ybc4cKeBEZ00Qfd/eqfRNsJXuK5b9OGTMOfi6InP31FzD1C1a8PONvTIaJmfCRuYhNflmTBtQF
ggEq57llWRcRssegDcqpDpIyE/iR9pykBDlhqoq+ewJ7arDfXPza9S0ilP6muLNwrHgaOGwtBq/q
m35gtA/I7D+85+pAGCHsBG+x0CciCL6CP2/Z1M0jLb9rd8VQRMd79sEvhtTY7t2bi9VG0iqEkrE4
33WISyYhylbeixfhVNLsSa6jYOw76HqoFZmGYTEoMpjnM2wW7C1xcuRXuG1BwbUfycCdV7m253Kq
6xrZv9xZ0XsjSAQSaeCV0hfUX/TLeC4Ohm0eCUZaQUp+SAqhGPD42ZMcgy42VbSgiWwy5WHNCi3J
9lmg/EdErttFKUNuyWeLBXPk38S7Gs1h424a7WzxCQRbpDH79EriyUqWAj76leF9PEKXO6iIsoNo
HmYBjDL+sZ0xUsqO/eMxNfVT0JxdXM4W3x/L6nm/rpaSOiDFafbkDaepD9usZox7w/9Kd/jNOYd/
FFf+xt82JhI/sq9W0XYupvLij0eH3LD7/q2xM9PC74S7Y5xS/EAt0WXA5UidtN41TUdG79DSPf8L
4GAFvc1JcBI246gFblaFauT8uxFg7GDPA/1LUidJveho5TXyOzKhZHktyeTp0BLoLoXFbSiER6i9
AjvA/LGBZhGJ/vWH9IVKK0Pc+FjJNxgoQ6ObZ/UuBYKUtB+6t57HOoOIzWDYdxgEilWvZSfA6W2P
+JjesG4vnB5fosZqryskgjNwo1N9himS5hcukfPCF9vTg5uRWo5LsnCe3m6vXKLyyF/Ev5xhRf+o
Zr/ElfpZoBy/u6rUmT+Ca5q+iOKv7eKc9RBd0nSMZQ9x/nIfei4zQRQkYzZ8sFxPPZOyDj/73kVF
q74sYkzHhU+UO3ekbfsaa+dFovBEPyQ6eSOH2Lww/bSoNPlk9hcaSdCsS3PaO3eHONbQR7Ukozeu
66WuULSYmNuOB4f9SAgKRQ7ybhCrJI+JxEDeeDuWBEheeiO4YkcRldTHKn8cM3YaBXsEdv64a0/i
3V/9x64GGo283jjWFJ+QHPFgPitFI9WxZOaYnbqXew/yNGXNXphvWb96+FtABm3GXY68HqcH0Zkl
4yqyi8a8TrvQZZ1A8KtPP3WZrTBPc++4LWTnZyW1ciTVPMSD4846HzloMWShlQMUxc2Nxlnc57fj
kCSTKTh/Q2zuYOR5xcx8yMMYt2a+0ZyBv/633w9PfJCbGBgY20qPY0Z6mg1MzL0OA6ibMGpZ0HNX
hIoZHqCaOIp5Mse0UEq+8Nb3CufymQL9v/XoMuYAslXIPMu8EwyV/fNq022flw+/VUb945hb6N+/
1lCEw8epgrYeEgegauKcjvYMWP02hMObiKGNb/MKi0yKoQxScB0NpYdMWpaucx7aTKv80mwFhs4+
XnTJRK2fJmzJznBsEH8uFnDzM5rqThbtKOe5zZPbHoZFyohs/DXHYpODEwAXB9tJAx8qTK784XzJ
HGLt8qQTTrPbOm1UAs+AmdiaedUOW+PGu/jMx2yuKM8/A9r+/bOP0g9Nbu5WEvov2LWoY4Imk/Hy
Kc7ko8JuRRL+IQd+coSzWMkgZh12OQahvP3hYdDRXy6arUoKNgO5tksWtuC0WLqhRO1Fmwtkruxo
9+Sa6zGWo10sfDHHCre7etvT7KsJFPxTfrpJLzj9jLMi1tZ/KY8vmqNYuzcziVq7xjIW+LR/tZyR
IBVWZdHqOKWac3I5zT6evm9hrU73hPpRYgowctAo4c3GHnKvgy4LMjtlbi1addYJ0KUsV9iEmUTH
dXRa+kVy7aKDGoARQRjBM/OJaZn+lWCzTlO36IHZWzmhJzguIgaflzLgHnvgOJSWUh04JRf1FFRO
xm/zJwk8DG9q6db6GlsSQhFa3BZjTRwrBeei4LRuBalIRF/nSyf8ldZVLZ+UhDccuEjAQA3QIgJe
uqxQgjoNyGutbHxq2QDVXhsxEucbAwaaga8Q0G8FEDn5QqimGP9Kk/XnFRiVUyNXjygwjbuK/E2z
oVCVfq2rt29B82GtTWXE3jXsQCf4OL6QkZPZ8UYSOqV/XERvhxxuzFLP86luDzLON8D7G2CQWaiM
JIrZ23lWgwpsm2I8qd7uPTrENp0IA3gQfbPw3JEn/MhRTMf90FxzB7ry9RWwj5roBE6F2dTamp24
ZbdE17VcTn1UhUfdCeSuI77OXvknyQdXkNsPiKLImaW1LB9BsBgEC4vIgikSE5s4HlkSoIeT1lI+
shO93r0QbH9zRGt00R8nY19NT//CnCF6pXLeF79cUwrQfLVlj05/dzjv4rSzPyFoKtTL51x8JAwe
Dd+s6EuVzJRe4pIDTwMsaRGipO41xBFCnjIgsFn7OZisE8G79oKSJ8YSLjErXXyACmeXG7qIqXhV
TQXg6m5fExVexIP+6gtYXXsiOGv0eBlr+730hL9OAxgBlJCRSmwpY4aJ0XWwTqzpbNsSqzsy3ciT
lUmwGL29UQxx89jkjaXHJMyIa0F9hotQM71RCa07Lm8la7gW20XOOSgR5QmWoABZktBDZge+t+Vu
eYI7D6pFUyX4vPyyLCrNZkdsnlxxbBEu1ZA6BDnst/zrB4Gu9um3nMMBc64GrP0UHCKqszJJRBhn
qyoOyY/FvzRMehBM6HwgZqUsm9xg7zPHmTnSMmLKof1DeVcuYFapPNK8oZpGSf6qRwEHY+d9/I5C
HCQsCa+dDgVUNPN8zxVn5loUfshvSfFIUk6pZhweN8Zel2Vt+BAOU/iTFUMt/spko92CbRKTbyUk
GA8lJFe+N4Lf5gv8aOr6+A9OHDHaCIgBK4GKuwEOlGCJy22wQViWCr3gsel/m/q1DAmGCnZEeEBi
gdE/g0qXg6PSsIv0tlXBfD1PSUf1xPMpycwH6YFy7P7xUKaVTtMlr53k8YMBVM8h7gVSckYGl38H
gGLsB/OgxEVSh6bRMu3AZYtYUwj+EqnFb/g7w7mfjpIM2aJCU4E9z0tklkQmW3x3Zm4Wfrxo2jfT
OBQCLGu+HxAC8IWpwzURYU5FwLZ2Fy9jBdQaiT5l+lIy6givFahWm48vMRtkT7pdwdS5L76LkNlT
V33rO6VGHSAZ1kQ2FHmPzAKJobnDkHLFKZFuBpwkUnPPymhcuNKEt0tFQClNZ8rYubvIq+5OrdHi
Url/kqP9pfxnVg5RD/s9GVGvD/IaVngMyr42kVSaQDn06WQyoUNO5qctmkNMhspLWSsfFCQgO2vZ
NkDN+RA47P2laFJ1Oz+RKkSh4lN+lRTNNqqwwdafwWa07FsSfMmG0S1PL2hBr25kdHx5hs2ttr1/
OQY2dQV3/Qwz3xNi9QJLSF8Fgd0aJkTGynOKOGAQlUsvqxC6y+gC+xiWceXd2qAs2ndPsVb9F/8+
p0MKCIt1AA1fOL+FhBc5BtMeyTReUp6GYZoP3rLFjwPiJBdY+a5+nNjVr+BaPWoGCyKEqG5ojva8
Nn2N4RuZoS3QAwOp2esKXMayCXfNwc9wQQF15nv3bGkzDQI/MsH9BMQWugRw8Gvnrwf1BKybm8ZQ
aBn8OX/4BfkBwDbtgEdz120kF5UuOgPYuRQxhQ6G9tBFcdHnNzEYYVdhHRe+v09qmC5ZykaRRdgc
jZZ+Cwpvwx7aUNcrxVi4tOWM5p778I2KIXsk7ayE89M529pkGLnVCE+EQXn3NHtxzKGXkL2BD3UX
Icf4Z2/0dg6kPAuPhr1Fcu8lEhADmm9VFN7G8pX+NTxYrAtQyZAUsqT3SsReenlaQnsJwKv1UALD
5BHVkTD0u5C/8rDnDhPJueVGu7DhlbrXOXVWaJ67i/5cPy7kkSFyLuiKMgsgjNEFLFLC4bPM/kBW
w2pv5fOfyOomacaDXb5tCeasLl0plov7OjdN6Ss658UwZY4dBoBwviHOwxU2ZXc5tgoty3sq6UDK
6HI+pY656GaNnY0BmLCkgEFJDGhLhVMPeRjb+8FNTogmdPuWrv1m4pm4X0H22s57H/BJoTvF2LAM
11kLoD7tlidk+iHC64Nxtmj3W9kWPBpE/2/ctBos7e5THa/NBdNVi6VGSuYD+HSVFM6LXXgXV7Ys
NTuGVTGpjyiVcINkANMxgRxW0Jv0au5ZKUg7hn+H8pS+Drwidki+FXRdUcwJ+AWKNlwd1vYI3YgB
tWC2iIX7LD6xO4XvjduVd41PsYv3d+1JIwySg4DVhbe7Xm09HLiIBj9f2t6qzCpzSctLqKZK3Gef
llnexBDWLk+V1S8GPLSMi08dvjq+r00EhNTzSjM3Jw4gNS7/cbkc9xB1Lp+FFcjrgu+ZHqlUlRPS
OxW01XphMZyn836xTPE5DhtoIlAf4vhAbhmSiCpReMbFjhSouJSBr5zcg7G4ahcWLcZg+sopwenS
y90eYG4uWlTetv2/T2VbM3tcYOqLup1MYw04kqFy/sWZCnajmBPoK++t0j2qsspzGnry5rWteJzE
5UnglegxWcSNaKFv2O+CwkzSy1Oft77gmsPKdt2eO1SM+58PAirpgr67RjD8GB7P3R3yes0QDV4y
a7gs8VooRVJ0uKTaP8+lsezRBclmRYxH2O5T5fRDDfHjcTO2IeHFt+XTgBVDV5EsYif6LhknMG4v
ytez4yibA+qhBhorbhCzLAZBEsHFsIAQHIHEwCL8rL+jsS7Opl1sTNKg1iCU+oHTJGM6oV9bHlkY
h36ix2L7NGKRZxDNUyWc95SIl1U56oQM2bOvEdMESWaUpJTrBbrac7Q2CMX+RIsURDo2ZPaIbNGd
WlG2dCwqkWmruv8qQ5d0JWBSOpDqGSRIOhh+NT4/MNXOgEnAlGWkuERZYr0m/FT9n3F4ZYENOKG2
3WDsWT4R1I1B/4Rg3mRC1Bearzh6nzCmhVB8aclkknQtwnrlvrBMzpfusW2jNfycqjcJBQwars1T
OKgxU3cNjKE7STUlsopm/6eIrv9AY+VpZd2yTgVVvnVi8OBC3hpuETI7AZN2dKKIRFAuaCyrobW0
5FJHDqztGI63myJiEnIejoA981FoRtXy+hP+MONquLi9mPOimfeo5lCNSRWIGwYnbYxpwsOsEtFE
fZV4uYWCOhmd3aZLHGUZMgkyLP7SCNzIm7Ib9MQ146FZ19RmYgu3Xn2H3yIBmGqYfXNJexChxRuV
GgwXbVEW47yvSDFIjwb1Jje5oAwbapbIaKHlhj3YHezrI0XpQy3QwwDiKxLElKefo6G6INRKSX4M
1b/1zaE63W3heCGpsWZeIDgjoqhTW4/Wi8sVHZGoqpNXaAT3y6Hh886Ok4pijDpu4hiva1ZGwsvs
cOXFhqvmF0U+egDcWGkziz70fTd5+QOGwWs65MLISi8mZoGX6v0JipKgbR4O5qIbAyji+dpdJQd1
RzLvRUyE/jLVhn/V4bdvdNfPbz73gxig7nHr5sSv7vPkwiHD49yCzilpiXjRTUgbduASnE97GQKf
um8ewU8mwqGfRh5c+wT+y6T0hY4LlmM4nWe5pVUHrt89ydechUf8T0gz9kTed7foba71af0szPL/
uXbon4SDqS1feKy1+3Xwsr+qGcaoZY/c+LNuYbbOqjVNH3MCsjqe5gaMbPx1Ya6nDNkWZaK3XqZ3
vAUZl8PGHa30ES08ch4nmJNZKzGQ0imC3FdhYir15BWQDzCoTt+1FZN69I4iOpB8CivP2O++9Mrj
O5PHyKVPrSt4DqhC7MsNr/9EuVDoJXzZDbvuTiDVDcb001fpdYOjT+C6P3P5pqNX/KXl1QvTWTV1
xnmTvSIExEH9FC9jNgolcEXA01ft99SQ1y2PDf4SkZgT2mAZeqzlIxNkfkZP5xeGWDUNlWL1hDf+
MKvHMycuUxRrqQBEBKm2178YuyZ03AoAZ8jQQp9F24uRBdj3v0vwUhm7BPk5cptWbWclSRjfphFl
gpdSH3eL6UbN0q9ufzv4mL+cKz/gYDCW5MYL2Tr9H3p52cQ+Oex1ImpWHkEBsd8N6jGcoyrJSZNO
HO0d1AmKII82A/1jCx0e/WA9bo1bw0QuHpz0AnkX6kEYqiscvnETxu6nEa6xhjS605cyyWsdUP1T
MBVkr5+iwPN7RdeLPgeHyxENmryWWyDvyThzrNLF6X8vAlzViZ3f5pBJT8B+ks33/OxlU+3s6zdm
Mfg6Mu+6gkxXiUBAKKHZatxrO7xogLMlZkgjKrdPoJ3OVvJNxrjDBPzej+KClSK14mr/rBe6zzxc
DbSmHdn27xRkAXcRD+dXUmJTfHcHoXAbgSeXE2acpO3+RsajC9lwNKfXZ+z3W+Bq1h+qqVkajXyH
RARafmMNpyOHIPW5klnsKzRkwClA1MzJb/eWgnzHmdTX5Gwdlumdi2pPF6IBU7gc2kc3wv0FIBWb
BOtbTyVVyReqcjvapGtsIu7FQdiQQkVZcIHD2TNTuwvwgggSrHOg8ZmP9iGAY1Unj3nNLpXD6Olg
A8VriLGxeim7ZToEyugym4AEIlMCYdexBwSloM28tsaC6UqUSCcuWo21VTPwznQkCbs9NK7Awe9l
7Haj0WpbHJw7uLJzBcMVJPDEfk/y6/Zq7Q2p/XcbtOeR+SmiS71PFi+zMuJMSIHxtNdl43i8lrLY
xgA90jqRlZVNC1+vrhZXxyQ8ikz5p3eC3Uxs4IZAOetFmluv+UscJWc1nxFwU2j/i1L743zI6CfZ
YNA7ZYwEgXpyvlqpplZhTKYDWegorzDp1Q92BRrt77zkSwDOLu/BcWzcbuJIoiX9j2q6P6gPv9lq
OeNyIp+pZiOjnl2fcMI/Rf193TA5ov0plXhQdCV7XEMyW5NRcjZ/Adem46GWLmm6h95kzleI+nGq
bPfx7uGu297GJT0Uz2MjLhIZ6Yfq6JL5Dfw+u36ts6uAFf0wz+c6yEgBpq8y2B9FjGnkFOpiGqX4
0yRULObIj2+VfPR2myR2wPdBciOHDD0yb2xWXTRey+pXy6DiCCzgQkAuSGoZ7eE8Wjfn4yMRMWsN
0mG67XR5Tvu9ctNaJAPCUvd0NnpKMjDO0BYo5oDnA8SiBt57CaCiAXTOJMdIYof8pwg2tzkfDjnu
Osu261NvDFH3TUhtL+o1tpxofkjitB5Ovk3TBtNv2hzUpIe+YhRv3eraKp7W8WwdTnk7odVa6RCI
fQYUXl5pi7ln71WLfyKT4M1j6JKawJynVXP+JVvTOq2MucZDwf3n3F3Qf74gh8mdPgXU5eJa7aPU
2jVzLB96xqMiFCcypo+5/zciiOkeHexItAbKVaLxYmcxd//bpr2rymGtDNp+E5G13N3lepkLTx5Q
jNWJ6T90jjGHxb56ySRA2teJ32RhQo+nuH8NOkW2lCO1e0/htV/XeglMxw58Sd5swHtemSTtHBB2
iMhKVOlWd/98i8wuR9UXlFvYpLoiVoMcOz3PkMIYfhgLZg8ixFtYNKg+HoUSkmZ+veZx1IjjgIzo
4oKetrUsRfv0bVIMr6+GwHpIP6EEtHH95ZQWgWWZajLN0lzFVbq+J6ueuwhb6q1wHyPIrrrSwZ50
QRdRzkoZKfQTUJDkRuWiKt+06XEik6zpYoyPn/UesnbjdoK/4DbIsgy+6grYvOPwmgfLhCr6yoWg
QPnx/QOlMI4bv3hUj/1yUdph8YA+qCAv9pzbXnDE5iQpzGL9ktS2nRwGkTmsF7aLl8g7h2MynvLP
I9tkf0bvx+lkjXReZvka1+H/ryjm+xrNzlUa4gzyHcgetTRf6j00apHJa6YI5Jq7Rjw3Xls6gqYC
N/Vdy61UVyU8CdxL2F1kmfGIAdcrKw5pDazgWiZxhFg3iyTHf0L4Lw+pr++NY9lCPNKhu399beHN
K+pi9JRG1nvRHlYgahqxibxkv3zqWdmYtAktlku38BLwaGTPcPuN1cxJgajfnv2aG5UtYtrWRPz8
dng/pQ5Mz1uMmAizjq3bt5D0FTHdE+nS96TxyXG2+tyAtLvW0Xhfvisct049dP439D/ZhT0YFjaf
HAscbsSeMfR41XF+rHXUTcrGvZ0mc4/6GELsLDiddfTHBLjWTvb+vQpO3vITSatbpf2UbudPDFf4
6SRsXs73M2JpuLOmwCW45s73DwHnv9DdCGj4gyHDhSLiOCS0K5/49/N+2AuviMyIlLipbhviulLL
S7Ot51Y13aRIiFn37IutBcBCqTJ1DvXAT1GsOnOFj6KbSj/9P6FPmWxgIsTQjTBOkwjeoLZ3LL9S
w+WnnOGwDhbKd6Gwpw9BeGf3lxMdTq30tLxGpNLfd1SE3VPbqEuz6EfVhBGflHlZnDGfysGzs5p4
Cvi7QIhWli+tfFxk2RBaa6EYK9qpssdy0YMR4ky4XmmGeQZKTLO9TzeacXkNCL/F7SqPhwlTzWYd
mL9Saac39qbwEkTlumHCz0PuQA5X1ySSgq0/2UzYb08AJs4tpS85XLHJOCdiflyQ8FfudzkEgxdw
cwfUiKtDN5YWy+z7K2nWYLbvSq8Tv/Wb/iaPq6UIVGLuouPl0fOKiuPHfA24XykogJVibgCtqPp8
0BfTnl1W/QrqAyA9wAZJWTmhToT97bbqjeUBKGO3dZ2lX9a5916jkG1zHo4ltoqL7Zbt3U7cnbNk
0joDjap+IGzayCB62TeuniG+HjIWaXYDi/Krt8yqMkdcbaaAQpXARvcWagSZKZj9aDvo+XGbKyAs
D8nhSeGk5eRhTCJxexvQdsKxWYxpIgxZJyWjs5ZxfwusuS4PYhA/b60wH8KaMKT2FcUKXd7p2VxA
m8T2BjWBljPB0uexoz89GxC/txI2EIMCi1H1ZvUKaZca/573L4q6vQEOWNiTEwRq+JA+2YjA4krs
ZbPDUU1Ok3URlUJEUkdRBXz/8fyiTTO3sp16GrIn4+uDZ00AsunFvt3pTRmezdcPc6Jq+vjUkWnT
TZMtrmEkgS4GdmV+/3puZMS7Q7kLOgzunya96sgyCO8CCVvYF83hE564bKVKGxFkSSO2N2n4qzKt
eq0HgbeqS91D7NcPKM/gldKJFj/WyIMpyxafQWV7VHo7JbHLX8H1A70T4i8DRoCIjuTZBMybmc8j
csIsPGVzojlWNhn/HMYRFi0nPDn1qlaLmHdKHDC16EUqT+T1G8ORhFsR/IRGQJfW12ny79jszI+m
DcV2j2DOeN5kuPBiENOXqOA7orU33YFQ1tUoH5t9VSPh4RwZ695ucy41pHIvlPUc70EF1pf3D+Pu
fEDJGOcWqOf+doZrChtGHhsJDEfN6lWyDS0vVapG0kpADBvUCJ8byjjApf0iUbybdZvqV/JlO5lp
bUBE+4/eogS0XpVkrQuW9YgwsbuauVua7nydWkAhkVZ6XDlP/UDFbwYdvneqSJrAHITY+GnWPETv
TUTjbwnC++Vw9jiESAfubx5iSf7w+pJn3l8bXwFdMW4IsvlINqweRX3AEG1UkD15XUNYLmQEafd0
kDZ7mMo5whEYbbZdrgZVdr3EdPn/SYXKzJVyaP/KpGC7qr2GeZX29rv7nzhDGbEhuMUE8fdw0K9B
9ADxGJvy7BowncG7Mw/y9kn7Zn6IQq0/HiaE0XcOTTo7XY5PYU9agm9kxsMVMZbvRUimP8CvKWOZ
gSlSCOYkt9rWDEnMRRO4Z4SD0aKPEFTtCaPW2463p7lHBzfoxtH/Oce93ybe7qufNpuTddar9mwT
CmpjwMMSHSIf6RuCvqofGrHUdzbp4aZKxKvhSgT6PcEFVnix1TKLm67YOeM6mTaWIputYRE28hkE
GoLtiw6IWiShYpO+akSV17xw0CHStGviKnpkf8Xd7nN2bAZBLOQ37vWT/UFb3Dz27Bq7/4NJg9uM
keD4wFWibp9MU3NdWtr7RrSNL7SzVVT/RsVUQgNecL1sd04NfSqJGx3ycHM2DVpOCmMSHzo1rFOV
OESuyJ0ud4Ox3qeofs7muZ+nji/oh77WO5zRcYxnMgQnGPOAOgIWCTM0HjXNDGPwFtU53BZtNwFE
CABtYttZj64W2zSVXUyWuh/WWUhh6GWWVM1rncu1ajT/2O/jac63U9yT0dVVGKB3RtYrJPyxq4DP
EMwwTmyTLwMh2R55U8V0v0eX/p1zOZ79q8J4nQfdFIMvoUqXBWaDYi3RcCpcWc4uqv9Nb3hHZ/Pg
0eZSfjWgfo0OZrSVVIpqbW3lRqGwc+PLBvJcENvgoxEq4dZDGnvSOScY/Dhbm3R21I/7lqb67I+7
6AK8OQXkGSgP+oWAvRWqJEHPsJcMNyNtHiyMIimAAHPYZR6mrCT8Qeg+W2p+dTy1y/6oYilR0gMv
+fgePcUzkBP4J0i1xs7tDgYdahcdcgcIlKxVAX/crohPKGgcfe1j2wWIIZ15xzvw2v+NT4nxhdl4
PlzPCAyf/v+cyQvG1NJUzvGRnHjKPma4Lk72kl0LALJ2yJN2enyE4V+mV+NIp3VzymWPNGfY+Hi0
zdYLPaCH75JCjLmqLww53cN2RmVCrr6yLylFrbx9HFRC/LlWjFpu4E0e13fmpyO28k1KZ6sVQJqE
N6KuLnPG6/3Ba3eN8KykdXNA/SzZtwX8RXecgDW0x1T+0eRe6eTPrKlXbxlLiVV4a8o+d9L+58nX
6n3O4zTux4Op1iykNf0mbFBljQCD0QKPDPyn12pTMjLgTb7lv9NsZc4oCBjDhOxWl0ZKw+AqXGt8
XhjajQrpuLAVIP9FD4rxMkmULVdO35ktPciKHa/VGRiIIMYcKwBTnT0DU2Yt7HGm9d+CmP2QEqsL
eqrAPMEqQn2G/hvoagPbI+DAaZBc9sQB7J69hvOm/4gFJh12QzmpEWcSRKLB/HjzUfkScfgzz5Ue
mgyzczQD02bZtobbpVeBYiefaDJToaJn6ehWPNTGEgCzIKQxpBFVUe1AuBybYfK8AWf9fTKxMQs+
vrRIuUy1s6UWqxnQhjr8oNvIbGlVqjnCovGcKWZOBFYcgZnvSmgrL4Q9uie6J6IOH9w37MaqdQF2
fuWC80orDcSNQFnVZ0YR0dWextwqqpVjsP9pu1U7w5tHcruJwLU9Wb4pINmpdhSHwtVld3kzJ7YK
UY/z49lnvnHHRc9tndIbSD+dU8bRvFsbWf0pHeyBtO4SHWi1dIDnzdNFANMscSi/DVCS/psCdyIs
utBDnJpA8/W2o67oYXOODgfI0pnkv71neLLUYMZST2/qa5jLinLahbRaKBjNmnobK+NP60WyK9XO
DnLaYBsGajd/NVyjWGOUOS9CAbi2Fzk5ew4v+H5rkbzgcMiXCReYFCrYWykRvAUtzE/Eb/gQkBxG
aodMACRdrjT2ntHhKJIMDG/J7oNyF3o/K/DzWgylwi4/wHkHUgPYrvOFL0ON9vF0TIcjqWxQDVoL
GzroxPgIjbtk4oJBS9kqvJ7YatLcNhs1UeynmN+WIOTOt67/3AYdxbsj56NnjHu7BdAk97I0Suib
Krpq8WtiWoa2rSE5QKOosZWFuQxwHwaTq5zRLJDJViDF+uADV+jwBTEuUPBkTGuuf+4NRqbbscV9
jOvvLvidYUa/1oppr18MLmfzGU8uRAIE9oU+QgQurzw+MY1KLF0xRSWf+Eb8YTXPZeLpLB34ddzI
TzqL9PJdwGdiY1s0I9/Idgk/ydSBbwrzCgIoasKtL9xgbvM/G2FWG64VvXMjG3xQdj4Dncd8A1xG
gFvPOseMmtEJWJ4lVG7B3c265+/lN5fB2NbC4FJqzyc8+/i7pFo4pBXpEZbH6o5NOSOBjMB9/qzk
7Zpe/AqC8OmzHeruz2fBRIRvDhOsRhUSWz2jY7f/lxI/IAmFRhEbly+6bLhHbI4+arYtYybrwuYl
34OMRxpZsfu4u/9uutuR5owFFZDAbcE6YC7pHaQ/w65BVV8aQoUkz1uFciQXTkHxonpP//m+bBRG
cmHbJ/mxefoa2QfKcrhl6TOhIH+PT8y11/I2/cTnh0goypxIO74JhoxG9rnNFq2FG9Un+ygi18gP
2giAnps3t3NXV2UGSE4xk3iyCbA+eQexV6lHSEtQ3l9aHn12lb96g7mJ8woRf2hFF9qB6MZXRI7W
jcX4cokz3JcJJNHK4G2qPz8qHneV63dSPuyK75oPd2fufa1L6LzDno7Y3zjOJYrSluA87nLgH8Rv
LasCzSh1QW1EJXidTGN90laNeM1mX0FDZeCtiEHRZ8mlUh43Sg7vO6iX0t0GhCKJABXojbu60Xmk
dDZDKtUnDiiSM1+9QGjutgNCRN2yKtfHwA8u7EDmkZQXQZQ7E6iZjAuCjE+jSNavkoV9JggPwQIC
d0BAkmO0Q02GX1HsnvL6+Z+TU8m3CrgnGt3lPpvWr+k7u+lN7BJLyy+8bzkk1lblnQGrnToVM8Gg
98/X9iDFuOiXk/f+LHfxt5hR/tEDpOWC9pzkfkyYNSt6DJ0d0bP6lb2ZkV+Mhkhrv9OOd/WVImZG
mUgId6WpU8e9w4lXJvyOVGbN2q694jfhjvvTausWPszt9zu4jcp9KTRFYbu19u4SKbf0fPQZedII
0tfku3RsklVCly5XAboSClfTrjnT/v/Qn7sUPFgkfZq7f2AXdc5UJ1WJEe30lHon4VQT0Yo++U2z
1dqxteHKUJN9YRAT32kykiCMzoay92c+rpkb6pu8EvjQwwGufLWuAbZ03FYzYfcHqWYobg9BzxDy
COzmxflJvDXpqS/570tSaL/zP0GzbtlRKTqLUgfQcEWKGVThCrC9fREXZPJYpAFLLr2aUywpKMHL
zbwAg8TbXiXgkMCFNU2z0C6J/r1DKixcEOvEIbcwnyno/5OyBpD8RCuE6ms8aLjo2nZG3BIM/pFn
ZfIeb6fd79K7+u3OvD4LU0HzZGDDVCQn23qp+XZKkINzZex2pRcSZuiPvbY062nJPqQOjE9Gs8dz
GHJsNodyjqhy/rBNltpBio8yMyrSWgx+ZuvCFmlFZ9aCVJT3i8TXPPq5QKpk2fAVPjjnyeCIfMcZ
F523CwmeN1Rq1c7cCGnMtE6eAKVuoPNrEpQ+cG2DpxO8TNiCZmjxr8DR97y9Y768SL3pZymd2cDh
uee4mVorjjOtyYWZAeNxrLKSTOdHnX3oj9UnOObwfw5WULww+C0lve6i7XZoY2H34LTAIEXjFC4l
pUo2GwghaB4qCzsWjnVO/ai3yKPfhEgs+7wgQ0MRVrIon2wtrbMBRnriVnFOjhbmNH43kz9GxLFQ
o1Zz2q34hFAPMzrP0nhPoKdPGLH0rx4AP96mz91gpS32UER8QQb5aAk+HnqfeU938wDZeRuJt1LM
XgvwQ3YyZZEInbG2FE6GbMEKXmNw9iXEu/3+UadtT61roVZg2IW2OkRgqq1dstPHjHbHMeFNcUbd
q5NRBOtV9GtfucJc13WzG1MHnaDCxWTeljoB/ZgJMTIaaT0zeEvr0wDyXbHaIXx1GG0MBRCRvEYO
ym74Rg2geN0BF9h8QqhIpJa3eJkyQXxDUriR6HoT1deS5Q9v/ohPXbB1qFCg9YZ5tqM4qBx5jZIe
dWilEaLbSYntuKD+UZgD9+EqD4I4+IBH4a9BNdnTnWgZUhqQGX1BYEQN9RmpG8CAVzhAHXYJnYrA
0vlh1nlDzbcF59trxY4xiVQp+w6ACq6T8KFwnIc4rsIfjbj9fsWr0nPVcgtBqvuoHZDsqh6WrQVf
+tMP8fhwYAj9DjWGyGnUl503Y0qFuAAyg5rKPYNSd9a1pZt5zp/rKvLhhKu3JBn3TYpZtdP8PG99
6GefQPfiK1s35QI+BFZ7o2AXynEZuDuf/BWBCJXZ9J8nPKKD1ECGq/UTBatf7gAIrlazwbjv/qtI
hT0LHjRDKX26W3Hl0ODoBGEG7OR+8NwD6qEFS+X2zTVirdxyf9VmN+pBY+vCxkZdalFCtyAShzQS
7PsdAkHjNNJ53AYOK+b1kIYtu9ZsgFlS9GQVm/WfTF0xaAtazlmkJRZTXqwo6cXcoF3HJkza2420
A8bYdb1K8aIdEhETUEOjzncHcFcLI8qd8JLk+I/KXnSYJcPdSPLRbguv+AC92+yHHk5Ql+j73A5A
/+C1oVBDa5gYCw0B0tVx/qHT9LxFfYsuRB4VPOqMAYSjB0TN17jmyd5LeglX3L8YVq+QhkRVEZTN
ZAkWkFii6260Qw8MHDgbO24B6CInwFb2+yDJx3dM34fQsKJiQajT5OjIEGwdwzpqcWphcSZizyTM
hyVsMwCyeuo1ztcMlbBM9xsbl6X5o8X++RKIEYSUPRYQFaeJ+fHpTTBIoNWRriPdpfet0hLcZYDq
8n70349P08skPbS139L1toNBWcMZJ0VNV9hQ4BbAwwqa0CkFT1y/1DELzhJTGmtA0Ga0g7w3YmYo
s2xd8SSWGdtr4Npxjkj35aFxPWishDHxQS5BXd9FWM61324vcqIW2SLPpFtUutxQJk+e04eDWMOb
Ho/pDk0G67eWanZpDQswPnOF39Z7P0C9mmk9lw5w9ZOMMIz85oL9uwO6AkblFKHohZOg+6fudSsI
UAucG6JQ5FeEy9PpzQ8kKamhtTXxQb8O1TqPtHS49+mjL71kPdvtTKdYvUGTIZwHlFGAFAjuASjj
nKqUQqSjqvHbcs/rYPpL9UJQIbzoBThZLrZBsYawCUejdOnvjSXYxKOttNBuDbjWPbtvunyrVzNc
6LtiT8BSiaFLNL7PWWd3RTsZEA5/eFMHCbMsYZdl2VS09Rb3YWhzf+KtoCmJOHIYviEeWw0hzVRb
Xufx+ehDMAIfjBee2+q0UUKMre91QcWRTE63Lq4iqnoBJfIoyCbZYfPm5zaCRXhf+NSKzzYAbObu
/0pikuRQZmkG7d5BVh/ByTVPLRqDii7YQ+d1MhpROQWHKG2a0B2lG5BWD0KfGpd4fN1iC030opHF
rJdVv6oiVqJbwiG40Uu1gQQKDr5bguqWLF8DP9jmyuRjTuJ9P/pdxUjiPq3bKJGrKwPiJO3GviRn
aO9qAjJO3RFaDqT2/nN6vUU5eNNWovU6CU+OL7e8GMdbTBB7Ama+g3klNqNUAy3bbdQC9f30eX/m
T6iLsWYZX3J5ZK/m+2ESOAIkR5agMKQXoLt4GT0u0maxxnf36IDmdMD7xWMpPcrk9qnJSRcDrYKy
mBQ+XembJngG4SPSk02NiDjF0RY1UB2Jk0fv6G7o7BVeSEVUAUTvy+rNnoA9Raq7ZQPhjPTYzoPf
a/ENkfdiCM3aI6orQ2GGflnXxcA/S2UMsClDJbcpq7h3uA89XHSdIQchBzhkJbZZeMroV4mKEaAT
ppN/hhXtSM8u2q25lGk5oednvkfOC2zHnROANcjaOnw1aRrg6uZ20Eg+f4+ndO4imiIs2p8Hp2nc
K/U/4OZWt4BKKVQXn1dPi8wbLTCxVkRwNYL9Qv7idDa6NILInS2uuDDOr9MBC+zgJ7yLlWLIQ2CE
OTrARDFH9DQnwp24j7vzGbyKRcO5Zk+YQcmV7gfKQsda4d7fjZBUA8zIliE/xoZ79dT35BllUs5c
Q9fhJ522QRSpnrDvZXFDfQtm5W4HOFbhPUIMFz7iLxa96CNv455UVYr0pQbOcrruYtmGVeRnp9/z
PXF1l6WBIWRHdZniq1nnNpjzFGjmkDxsnEV/J8spulQzGBcpxg4H+v2QoA25FwTN9k5jcKiccgmg
1Qcw94vDVJisLs/s4ZktZgLb2yZIkYuAhPGqAl4cKvfpN4kqb3aXaQ6QMGGkd+rOoi0npbXc/Z3Y
ExOI5S/OGIXwP+eY/QuDvDS0pHwswRxoIyQ9sAOdQU8L0VsFjrpPBV3WXiyPZkSc8y0pGcugNmOW
D/RdlEINaRdYtRrC/0CZleViyeSodxaOp6iXXpCwKG4YmerdGLs1yLlWRrJ7IfeoVR5AmUzJ1BKN
NTXfvAT0/jT5JFAguOEwCy5Q4qMAr0zYYcYmUa2BH/4w7bj5eOuRuKdjUno0A60G0qvezcLXiPd8
1w1b5fTHt1dB2rb2NvYECh2J2bVvCZ615RQPMDKKL6TZPjKjRvdqZcY2wbzZMv796iMvTdOKX9MU
SGMDBelyg29u/QOBZc71zqylU8LfXHKt96AMXBJRSco/NR3EHoSZyMRY7ahKPdx8VUgLprktn8BF
Wt5k5h4TozTmoGRP8Xi2Cz9dZISwZcBZH7UL46XQClSuWXP1OdH/KoVVQMS1hI0zm2D6P1Fa7t+8
M5/GKx2HRdWKr/xUlIFsFWfN/Tp2HHfgq8BMRmb6KvF0x2dPpSNHGU7MNBUo7Dex6kfwmUvzQuQ5
c2PBrXcXfoU8tPGUzVW4lZaJtbrOdnRPGf0X3kwXxC5tvLLsg7TE6rRlusc4m7alLLYBFi+5YBVz
eRbITT3zG3EmZqdrC6jXZFaj3lC4Tl3tshxi+jbQwZqQdXSYjBRDRgayXqR3vm+ERXZRI4m1K8K3
ACJIKYQlVxrDKukPnN45MRP9/TBW9bzQXXuFLNiqR4+L27hGmwUbdDAKRXZt+ZnKlhJ0iMi9C2O8
wXyPye0Qa7A+EaGwkD3H75CxHKQjR4lC1a+B/ry4Tf3rQda0WwuJMLPdT1bjb2iPmW2VBVpHACDc
pmQhjocDIBdZV/rzLogXbS2FZiZafl79HSJEME3ZeS8O1EGqluk+KU5Sd/CLbqygoOAonkRtKYuI
R9AmhDWpoU+DZcJnhCLOmfNKtY3dVgFV/yjbWKce+eCX6G99Rnx1cK9VpKv5YqF9bIlFCWEd3jp8
4EV1T8ykrO0FC/DF7Jh0cjPoqQ/wF71hka4Eel0duHqW6hDHMbSjI5caIA/CyA3fzBkNLVmu7de0
t0G6kmMWH0TSmVSJW+MyAm8QnDP+C/qqhfUmzFvhpF2SjzFAK40cXgYDqqehgvrNq5bboqcyis7Z
LqEnjlnNUSjFJX/UEp3zfMCdmgVxU01bQGKB8pB7ZgUQMXO62TDObxx3AYwKX4YsVxSHuH041vjg
VCsg4hkJxOAUdTYUr06ZEq2bwJbCIqeL7W0MotuYpC3UcbYV27WzroowivAZmvkNAMDUOFL+s2r/
3GhbIP+gkhvkiqXx8CA4bb4f8ySbicYIK8F6XPWOvBla00jDdB7F0Bq2xH9TaRF0V+PgA2XTy1FJ
mSJkP+OpPLUjGDqgs34aPHsW2NarQR8VoJtaIm7k9k9Iv5sQWsqW5pupH9CAKMuURv6gPvGAFF1P
Hk6V+6+v8pYC2buc8xw3ZcWKFWpCKCQg6dhsKdU8jnXgJurMUNlxxwBPRXj6Isgs1kWplwsiecar
bI6F7oD27JvVzXEphzqHd5edpaoLsfx7Q5agWVY1YFzV4Skg8a28ScLLDGs2RyXW4UWwARepKp8q
2GieyEVrNeSPRLY22lvJVH4OOrxY2J0x73m4hYf+O4M21bAw9p7baPfet+gD/bJqbcHLTiEXt3EB
2qcSumDJO4qVgQRW6X9HcQ5wvI8AwX+BjuPtaIgw8QPsemx+SKH5RyziFBFJ5573iNcdRqHOr8WU
6nx+HMNPyJ2jUc1+7WTVrEbgpJP0Q49YXlNzkQTTLrodnmpNulv1kIFCFBG3aCXPQGYY1v9hv+ce
kvV/erCZ6BHMtpUvH0gqb/hzz3MCWJ6LLe9DhOa81+HSdjKuo2NQrelCEI7gwC1NvfezfbAT5qIv
u7UfJspFDl3g6ZMFeozbwal2Zkf9I4HEhxQbf3WVAWHGtPB4NiOxv+aR/FQ4vNT0N9JA56UU/Sx3
z0Pn+E9qN+OxtZlcYDjepZqRK7B8X11dDjoRDsjyEGruPESVyNeeVjbof3CUflZyjj53sjZqZbFp
fWducQEUvuqIdusoI9SvzmxKK2bTCjfpcGTpZd0ndYa6axxax6mq5+uuJS/OqD3nn4/C2GuL21Cj
xBPFWdo2qOrg5NhT4R+AFu8LNSP8+Cy3scCyKp/eOSJu7HITvLVSfqrZ8kDbuXCUk62qlI3X3x8H
IfCuVtgbDGeATmcTBc3dNxZuWFrY1AmXoHOjEVr4DJW1ZqWK+V9ufuftBKHuIu7TDyb+hLnvRls0
+yaxMlmcAnmrTBqr7l5bDgfcut4WEOMCpkNGq7Bk5ON5QjrR36VcCfLp+eJkOIOxsJ9bobbsVo+Z
pWI5aG6INbjFOQPvM5aWQqczbGMcKhAA7bVkxloEOvS3sT0AuxKif9jmdVlMYCfP0Cv/OxXxE632
XLgkMl8oGfBnBFFo7Ej8Tq04vAciAvVz78YOKwpj4SbrH6pIAJYJtIzhYgGKPWXUNfVRztHmKOmB
FWNTxBy+4s1LwWJ7lfpKqxQoMkSrA2BupYRK3Y7fzK8J+FLLh7iHh4yqATOvtJN2wWGiI7RXVxlS
kLQmRk2/J5KLpmOK+a9OmthB0Z5++UwSSFmyZiLE3nAnmVliXIJaPqeu9HRdYaEJw+r0i/SILWV7
PV8/ScKuVmxHVOYiSw4/g1IodL1RQvd5Ixl+0ZqMu2qRu1+wNdb4aMl6QkStmJYPPKF3Sqt78cNv
pyEpX97NCVRO8HFQ30evedUrZoV9xI0cxE5YcSiiXLm7/vloMq6/AX0FBYI6dXNL2KJraTUNGYtm
Pat1jZfMRPy4Dj9WwE8rCGd04DhxDGMLg9eSIsC/pbD9BsaoMBXjRi8nO2/gTlG8d6cWvljyTEcO
VcF+JveePFhS7dGps0IbWl/ozf+536IYToefjxlWqwaU6L1QM5GTJLEVpaIDBSkaagyJGiRI7uw+
RJaYBPBWmPdhlQwKVgDaWUJbwrsQsviGnb6H8uuVqjziw59xgYhHOCP/EhLyh8WfuKzQhf6Paar5
dIPerOVB1t4vcvyBjtS09nCUES5nQTdnDHb3uxU1YaJZMF1qRJjzTWos9lTBiF/SCPuNMx9/GP33
g7jzWrv7dRhGchmVKxWdKZCFT8ij6kLPsLvR/kYWaYlPpSWeGxzlT8SGPiMK6wp0mYBn2j2XwhNw
Nb/t6L61yvfOSVT5DLLb3GzJplHFXVkmLCZRA4xYKdOF7/ZKpbQbER2cyCF12wf1DGdnjI2QeHAv
Ko+GWdnbCOUkbbKX8ovbeJm4RA82sEcQy/b5VwI4tP3VFOKOQ8nhY6y01RJ7U7LhulJQpjH23h1L
KlHLjrKKDW/pNuL98a9WNCdsCRzdbuOwZvXPYedLhpBnG5qSVVpp+8C6BVZBAfl+/3wDpw3I1aky
VrhbdeO31ClxdNg5Si4yy6fuUbvGE0s8DJJHghxSbpLw4iFIBPpNHEQZltXE1Rd8p/7UyTdTNzd1
OQUxp2LnXDOwSEryS4BWWpBsRMbku6OOoahUxhFrtf+zor5obbRn2NhgPm24TAxC5YyuNVIA9LMt
1MHiU1WgfJPS9jwtfq2WGdoLwvaLK83mENZlS8swWPmH1uNB7ofskZusIbKSf0DVgB3bW0Yx81wa
lJteyNmHod0Xb4Q8+J8Pd5eAyVu0H9FOdgGGHLdK+8k4GpP6Wt2d+kCrxcTPNhHmBrWl0wo5iqlO
/p1poE1CuZOSXsFUoUqjP/CImq/RWgS2qTadLzjRd6YfM3+NZwd1RVG7sr/BKNm4uamJbSG0CVi4
F5LL3+fp+78KHOpuGHITX2D7aNHGM4dAwWbwfacyyPEIzBYbTcI1l7OjQtO0s3P0lTeoUq4AwpXF
K3wnXrPxGtPTrmWI3XqOKX9EEk9D0TvwT5GKnWW85UaCAIiRBcdJitYxmprpQzIXx4hD03pGMvIy
pCb/
`protect end_protected
