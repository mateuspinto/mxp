XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ˇ'��څ�!�=&��	� � �K�<^��g�v��d�����񡖰�#TKw�!L�%[�H��Q5��ZO�������ׂ�B^:�|ˮ�%��5���X�k�-��z��D�@;��2U�5Ek"�^͐�5�!��7R��ܜ�G�����_Dꞕ6�I�*tΥεWZ��"J���w�K���oJ�������iS�!�Z��^T�`���∌�4Ϋ�q���eO\F�5!۰�B@� Dki+��R,��v�.����Р�P2V��A���To�Z	�	�P�g�D�����"�IS�C��e�6�*Ɋ&����b�����-"Gv�"I��M>?wZD?��	_�S��m�Jϲ��,@��G����7L�ş��U��	����"m���9�;Tk��X6���&:|�����xp<��O܏t�#y�+9s"��<�z�^(b���&�dyyz�DOn>r��iƶ�������[2���J��u������_����H7�M��g޷�����H�m2jD�ڍ�.j�< ��^�ұ�l�h�([$)�P��3kY:��+���[�N�
f�+�AA����㫙	�<V¿�55?��!�����a"��֭Hfme��^�Y���m��nC�)�� 3GM�l~.�.m�(kz/R\0�WS�:l��y5k�=dP.�`�����̎�L؋mi�}���p��G����[�ޏO����N�9�4*uv(ӟ%�%�s_I��
��H��0���c�~,��c�n�;[�-�xXlxVHYEB     400     150S�Z
��q�WPB���
S�<�0��/�y/�M4�R	0i���BT��QP��W:Q��Am���
���d𰥝�-���A��zM��1Q��=3�(���j	�˺"������3��A*^��sL�>�8�c3e���{Fd�!��*��E�	���!��������[�\�����J�U�0��ߛBe���a�M��
&�5ǹ�7v�4�R��O!��LOgY�
�e�uP�wi���(z�Ƙ�D[��z���O����3P�Q�l���J3��r�W;}kZ�yy�q`���rf>���l�/B�����$��D۲u:��b��^Z(ݣ��XXlxVHYEB     400     170�'�������'�#T��Lk�������B�5b�~�J��{'��ϖ��Z@��T���2OG�t< hHG�Gg�W�g�Zk��W�T���,��ғ)���l=x����]V��P��#�Wd�>p���-�$�;H���.�"�yN}F<� ��S�4]J�.�^��݉�Gy�g��u��k�]�6�0D�g뗺�E�Y�Ш5Yڗ�tlf{����5�a�rrJ�%�f��(�4�������'̿8
WX'Ha�t;Z1� á��L��@�{E��	�t�ȏ�h�)����I�ʹ#�R|��uba-�E���܀d�z����6̧�[��*yO���0��J��]��B�v�
��*���XlxVHYEB     400     130cs)�00��w�H���[����ݒց���+Kq/ő�n$�U'�랩�:�����	Ǝ�Y�Qs~7w�2Eo�L /�e\d���e�w[�7�S#��W:ǉԅ�9���L���W?��]��W�W����ϫ�PoZ6�t�F�n���� �M�����&��q~�T�����\�0):+� �n&���u�W[}h��mi	�T@���y�HB��,���I'G&)�Sj�p@�bvb>�C`诐��-��Crd���B�v_h9��/��tI#C��F��P2�m=��|��;���XlxVHYEB     400     100d"M�>�"cS�M��1CC�"~;>��$\y��w0kZ�(���W�2��?(��fsI������a��;R�Q�E�r�k�?�����6�j2�M%\\��YZ�SVr��@���57�����@[%z����� F�F��[�o�����:�Y8Q���$�[ъ�(��Z���o��)":T� ��Tؒ�`f��%D�G�C����^t+��.�)�6��@������8i��כy\j�[$tw������ܖ5XlxVHYEB     400      e0��8���0��wN]A;"���b�I�#�Yʚ����3)i���fv*w @�"��Ym����H�4����r���È6>��vt�p��Ƶ�	qꨲ��Î�~B~O$�'U0���J��k�۟��B�y�Ko҅��
LB�#�����;���p0��I}��&K�_���AA��YE����B��R�E�G��p5�3��O��-�Ea�Ը���e�;(�O~��y �XlxVHYEB     400      d0������
�R�%jA�{<p�=��Qz�4rQ��9`eқ/����c���Y<g.>
R�SCGN*2����5jL(Pf�c�,��w`�='FY>P�y}qdY�z��ޓ(~�%�c2^�8A`u�G`��|L
�	��ȵG�[���K�$�:��S���Q�U�����T¢��](���e�!�F��s��!#�i{]�W>�]烛��#/�?.���Ý�XlxVHYEB     400     120��S(��piL�������&V",�(�g8h��%*Ɔ:@u'	�GI׌ML���2�m�'d������~�+w5��e�V�&��]Cr�r����ɞ�ޜ��+r��C��:�_$�m�'nS Oy��vQ�c��������:���#v��o����31D�6/����KPٞ��&Nv����5��X����� ��lKz��WtY������m�)��a�y[A�����č-�����$���B�t�[��Tw|\:L�f��h|퓗����Fu�XlxVHYEB     400     180�T+�9_�F	4��tnVE&,�d]�O�d�(�"Ȝ�!�܎�(2Bu�Y���m��)H	L�BV���b�igJΫY;Ҁ��,	����g
~���N�+5t�4��k����Q���ͭ�Z����8����GR�u�i9�._�>�̶���3�I+c#�v�n�����8Ӿ/��}��M�[�r8i��D�Z�ͥ��Us4ZS�)�:74�C&�)����[f#�f��c���]h���4v��i�T��jD���{+��SS�/�:�X3��q4�c���Q��O3��*���ށ0�5k���j3��׃��hRōq�4���~�Y�y�0��H�=���ǩ]Y���A��7�� �tպ؝��w��6�KXlxVHYEB     400     140�ۥ0��bH
Wc;g(���f���-R{�npu69L�TH���
��%��G?�!,��yzՇw<ik�P��/d����^7h�j�,��������;3۞���9>R
?������~���T��9�60����j-�N��>R�_�G�F�n��Odn����a6�T�H,��xK2���R4�<�N��Ď��)��j��:��u�D��-ܔ�!*o����B~T�>IW%K�LO��N�O�~d���>�"�cg�,/���8��	����?��x�kF9,�_����?�8�����i.��MV2Kc!A�UX��r�aV؛XlxVHYEB     400     170׮n�M9�It�{m�,�}0x���/Ц9��pQkJü|R �vx�+�D�����!��"s#��5����#�ب����0�$����ϩ�_i.�Z��D����Q��%},#1�;Vi�F�Xe,,9G���r2k��N�� ����5Â�Hx�duj>o��W���[�y �?��լv�d[�'�_Z�q��/<,LW�
�����Z�  ����n����.��×/o����iu�L��K
"��x0��T��6��>]*�����`-���@�P�}?5̾>��wR�\t|�4"zHQ�)�ef�w������}+�j���&3nⴊ�V�4Gk#��(��� AF >�?ꂍ
GXlxVHYEB     170      d0�}QS���I��h�(� O�p3f/]Վ��)����D�p��%�[���SԄѭ6�?9=�l�z��sb���y�a�0�1�8
07v�m��i���C�s	Vr��i�k`� �ǹx��9�fvR�g\8�g�0���1�嶕H0@�,��הf�����5l��k��f���x`kJ��S�8�L�����ki�h�dz�`s+Bw| ��{