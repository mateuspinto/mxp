`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3168)
`protect data_block
9vd2JCBZW1Z1akD9Z1BQZDGdoVV+odk0cQe3RJQ4Pl8EXHSrJsLm7j0eRyuKbRo/zpht1Y1Ksk1M
VgPu+c9T3hWmoL0tuvEBrtyIzVdeYkkjP1ApTldSnxctfBqtf6OBePquqqVeUyEANA8yv4V7gLeC
fxklGxJgbUcfpsye3XmS5ux8t+agkGJDgbE+U0Mu9g49zoK/QWh/xz372l3pmHJTO3MvfAciW/CS
JHJg5xV/G0SKAnPTPzI9Je4eSEX2e2+dZMNL4g0WQvAKpgop1KBoKWn2vozWrPfGbvcmDBKjzLTK
jXD44qImg4gzt2mu5/LQpXTnalxGj9WYvGKtuTdb2w/BMX0/Nj6sI4bjltCmD2mqCkPitI5B+STk
OD2fH71rrubYOlPv77F3eoixz6ncFVknJ9RnFElRxO84wvTDtF3PUr+/xw3i4tdlGmQcwWJitskG
twbyiRml+vxYwMkrRmTbSO5tJYTWCg2qTJa4y/FPKQZeSeZ+noLOGFn+8mpw/0IJT9/2Anl7d906
AIvin6wD3mzGM8PPMGHvkCV6Fvc3b7BkVIeUT2gWuCMAANr12AnuScuvyQy4U3d3p9RhbhUnbMS/
TFbYzGQDWxX//ybZl+Rkq/7cWy1PaUxqzcEOreLqcB9txDer/+zK78SAI9PFj8OeIatr29skCpSk
E08VAeF+EpUDr3zk8wAGdjYHbv/TfB0nlBqZQLagP6PDYsl1sFL0xEQgm+ZytvxfY8qsvPjpcaMJ
OB3oG4bn1l4Nd6Wk1/N6zLgxs6EqOiOO8P7IFH3obk/HxNUXLWXNCKdMqguyXI2dbxJvgxsTByMe
GzvVPAbyPprTNWMieBbgD1OQMj0KXGkECx5jhoDP/h4JZ5scmbIysQjfkvPWtrK0nTw9KiqprHUF
m2wodM7VDLafVZbudsnuHk0Vj6K6+Oly3DyY/rrdMIz6TUxN0h5yXBGnjDcrGT+k/CBAIup2Oe8b
38f1zlfK0U0PQMZkdVZF4AgqvZg3sxFUkAD63xm+tpfp9c5yxsPxQMGdxw0wcIv0Lu097d+bMYGN
b3NzZe/RYOTx9SFC+Q4EyZnGRxk4/1qXIxR6tz1KCvvUnBnN0KUpho6TKGZeerajIOqT+5WQrjvp
5Ca//od40cjJ0KrriAvuLS7KMbnkCN7fJrfvTOoOr5lZizyyzDj+MgmnUCgjOakjJ8jOA4UwMDJB
K2akdb5ybHYsUZv2rRM1Y3/QsfZNza27/GsolrmYNEj0M7qsA6ziOtWT/TuazMa0gALsqLDUkAXn
hq8vrK2xJIo8/OPT3li9sFmCukvQTSd/wsh8vL3Sd3zhn8QHCkGXKdjuhdvRqO8L8YyWqve6xjgg
lvVa8YsKUfkTRONi1Z1TGwa9Gn//csrZSEKIs8sm9lq/q8z9+svRQNLZmwlsrtsMBw+wpblZoGEC
G+jLSlzmhwDg6zVH9zvb1HAHiTvJeqyUXhWhxcjt/W/6HBtonm0bfnjhkOqlJQaEVrMfm/4jA0Hi
vBJhFz6Ytfzg7PIH65kfh6KKPVR6h3cwQhAD/b22rS/CNT7JK/swUfG9MZW/tdo+a8DZKnALwG1g
Q5vCNjQB/w3rDh33cU4xcD8bEPE5tSNHCz5AMr6Q5OeFEBvEZrOzpmjHAEShp+mWe7CJ8Hxm0bvH
VVQpcQGO/QJGoHymRe+ZqnqGfAiTKauwOpmxVr+yaB0fQaaeK6J9PqAC+849E+UsWlLLm1TKW0Xm
2INXERySpDfy1dQDOATS3Y5mJ8VlGB5NrCUKCdjyOy3uCVpk7lpp62c22cMLhaN/cEmvKyj1t75i
dSmvPz++PRmiNdEfWFuokEC8R0mj0iyAtB0TJi2pH+0pRbPehq8j8gDeHlC7XRjgtqmnwt127uny
sl1b+P3WFOV/xfrY25H8UwMAvzzkxBL/1YLOhI+gFpmIHZ7l2jZG603E4njxo4/w29TEwXj2SbzZ
R3XeWzVkP41SunHcbAjFxNz9S4HV+UtT+897UUhiu6oxTIuyHGlaoXakGSEFpXoc7q6poD1Picn4
NdUDG/P9ziq6SaKsmRz5MvzyiiMgKncCqqY6dpoD93LpgK5jx3UCaOGU3qzvpFxZJqT4RPER2Uwi
bUpz/zQAwivTb+V3I3qQWX5BGtqiSIpPySznjxuxGch47dgyHtdixNNMe7ivoe1GV5oPo9ACdIoh
mruf4qrgU2zN/97lRm2QJSzltMrIFz8mPb1u2hxBgiBma7J1VSa2HUTtn2OYhWClMBPILZLpRNEE
ct7/CUlvKC9R8tEIzv49EVD9O8I0rEVeWYaw950/07TUNXvmuYmweOHIfU77SxKhkhD6kB7elXzu
YdX4CtGJ3/KK0U95DD4/9wQc5rW73kd2hYHGXtyBLUFczakO4qzVA29QUaqodZwpi/L2OrzZqdCI
ofO62YPWtvXyVBe4kMOGGzuBfwyWVlSaPzm49LgrXWOozD+QIsSPf+WkXBaf1P5yEfvHA180+NHI
0HRNJW4g95gPeDeV27zUWhj3oP1sSxwoOqe2yp1XWCqOENXgzpPWP4/tYc0j6hW9zZ1nmT1U6oFQ
s/TKcECD7v70mMEMJ5ujbzzxd0wbjTnBZmYYilpQmUFkXi03+jI5VmNN46gnk0MQTEQ9tRvZ41/7
qxznXRd9XmBqtj4vJlZBHzk2QI9ZvoGR8z4mO+wBWOgpgQQ+pdrGnC57kXqBSKWyeEKO6TCY57eg
xQQOdUWmKT4X2QZDEWrmmS9Ht2pD0odDWJMzFgU1IVsDWYn8VFcrd6Ypc8owG/Iu3wSGn+ZKFyi4
LYu+hY8uI5Xv9eQeUnXdXPnvAbsg4i6jPw555oHEZ1+w+MBlFAJc5Ae+Gdd0D3ajDmjxkxp6fHPd
eLhFYbS8I9/JF3PDIg17cDVIchuDJhU59OUDvLVaaOBlPfd3lnRNMTceTX0HH+oApOwJyj31fKzH
DY9DntWiPMgPLpi7CzZJhRByTqx2VDGeAfYQo8ILs+DHzmg5/L5DIyUHmiyPCJ6BM4r3ZSsZpDYI
Llzv/tkUlQ0FGcX2DFF0Q9WlVtJdbArrHn8+2mJ/dwySPd2vrR6ngsu1G7MF/ZL4IOQlIfHv6gDM
gMUU93gH0GS0rXvykuaIummEFDp2/DMjS0BgKZYgxf/35ylulKFoEf21nmpwWZlf/9tz5KnbtYbo
kkqQMLQDIxljGz9kko1d4ux9k/fGaFx33PwPOxKzzQbK5eovNAJK088bIjWhNum3cL8v2Ksyr8l7
PXCMdLA78+RAm+/xRtCMjfNpdgChc0n+aLSGNr1NNKSBwOyiMW1GLXvPo/3CwpHZei/Cn/igLLxZ
8Ys7munEtRMOJJOMWuydvfu9HIH16a028ChsLPRKw7CCGbXDxJcqc36gjgV2g4NnmeWUDN+8hI32
q4V7K0aKXe5A/AlHvUwnOrtEA1TXTknYdIdIcmzvo7QGtE2CbyBF6kQJCY9BE4BTaQRRg1owqElR
Xqb4I7bvuLG4Mlc4YpPPnMRPqR6X/yxoLVlmBbKOzziwHhWALj4Pu/Iheo/r6AXCU4MC9Qu2j4TB
8XKsy++WajbLYPHozW83pvdK9n40zYyTDFhunAEdFQcBN307fC6wohCDCfIyaSvNH1eFypNU9Xvm
FT+uA+SDhTuuwxdUkBs+rxqmXnbZUm6zR9woVVeEa92kNcolhOZSny9xRroCouZWKMU4WvfDvoj+
qRLUgyUvicker7wVPMPitkb6jZEkLMBzZPUxS9okQi+be61C+PU+pb47DzGKmjUZEuF8ml58aLZJ
9T5w8yjxxXhDcGYqCmsXHuR1QYbJXmzD8LOBQE57W6Q9AotqdgsqXw6HDgOg4JX4daPtVGi3a83l
udhm3kQ0K/OyPQb2DW+3U6NMjxR6GIHkUxoEn+fotnzk3CItA2TuDFHqjqXO7ym+Tw6nu1GaaekH
S+m/NFCYu0MLtKiuEUB5tJbgdxKOdd4GfogyaY1Qbbudl2y6dKpHxfSLdb5qSG9tEIYT7G4+QCDH
YITcJ95XzASH4FMRC92gc+mZ4mfA37P/MOhjqam+2h4KQL65NHR791i/fIGJdSUB5zO0tSaovMIW
ud2iD2SV1E6PZDzk77GnhHbjcPBwBB3myIW2Ro+fkoGYwDy3sObNfLXClYHqxamf+LmcwlAZaQnE
0M+agm8FN31kmibMtHFTFQgeOT251qltDTqfUsSANwMj
`protect end_protected
