`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14864)
`protect data_block
BecqBaKAEEbggU/iuxdwPQ0a9lCXH04zodob+1VIyJ2cR1JqEbeQsHn3pDVfOaOhB/OOXzKyMNUd
PyE47onI1Q7KvJdIZ+K9NmyKLu+2cTcNTA+5pahnQWFjwGKk2ocA39Q7+96TOZxQQIpZPplbjMw4
A76U9/1248dlT5ytSqVM11fCuizeKyIkuV7AqY18UwMrzzb136aGFMqZC/s7QKPJ6xeKmHUnTuwD
6fyqgyubXgton3I4hAfw9a4mIi96tD/na7ZqUIIe15OZNdcRBkiWdXOVanYdfZHMaq6RRr4QZ+qM
rzu7dsx9Yd/bqcpFV9yRDZXvRs92GPNxvXA6w0wSGHiLWWBPrivE68p8BQCS7Ae2EZUlg5iOk856
jBkx6ngYbhO5rdBIMAFP5eBLS9DWCada8+99tn8dgkNOS9U95ttJqRmPUq456qDLuUmKmCoqoH/v
yTj129zMictT26JDxvwLBgHfGb+7kLVDdj6HIsQFihM7lNwxy5C7r+HgZ3ZhoH1PeUe7OlrOGCWi
tE0i8EVf5CehLTPE7cvaPDdJ2rX7YWGydnybYK2HNuCX5GZwz0dB5+j9TviEWRVROHZX9Wif3aEE
mKf6ftj5Q80iiWtPp32CRO8w7w54BQ+ZI4UU38RSDSBLph4iQw4QDgQ9MDz5RgKzRkjJnt35UP+U
AWHYuncXOA22s8YPsKm7Gxjv7KEhz/l9mMLbhZj07u+NfbG9vJIbJqf9bbA9bMSiht//E6Spz97F
jpyTEf4zhu0XXWML/KcaqRndvh8Ajwr55ScVizTMb1Hu3BrYmH/hrvCsr8RMVo+7SU2OgTdxiUv/
oZus0QTxsyyeLWxtsOVNtmEuqvdZbePZpK4Hcw4aVgV0teXl+OallryLc/eVV40i//pdAkX/7K8Y
y/+Al79pOTF+pnMRKIIHD0PEovpczaPqWbPl4Cj65Eg3tiaZ3xZeppwD4IIEVkYldRO5IFmFA5DV
gze/9L3sRF6YFjhoPXOhyI5fhelQToG5qV9ac1vEoVz4s5F0RcdCIlIE44HywSfOwLaTIAOLzSRC
YookUCfhecntDsoSV7qYFQ7Jj7XWvw4T+Te4n1VLICGj0hLLKO3ECDU6DdIhRuuqzbM3QmAMbRif
1qT3NC4+2sZj/sGrYcc0PgL9xRNv6qpz6CbbvcRBE0ggQJDw3GeWF/Hp1uVtbawYoTbcJ1wI8JSV
lWsKzeqdyM++J8yDqZhqL1/HsS80s/6Qn67ErGVZQ2wYBUBN14LVwZc8f5th1jBQmTLBIULYMV1b
dS5MuqYynzjD2uiC6F3/18x118lFG1+7xVdry9X2EhRLniPwpE5BaluxRt6HAvpays+W7CVKK2bP
SnckQvXlF1Uip/qJv5mVtE4mWx2Bnjv7wfoewh0sJs9GMBTQgioxKmYMSORAXZpXpEQMPYK/fo6V
1bdNK0ExEGftqvF5+fc9yvkxqyNzOPXD3uSEiK+c9pcrIoGoFIpJgv96D0ynOifSu+3ubdKsp1FN
VycKUxCFlvcbxvMICKtdOfDOaL5p219CjmsYmubrR1jcAwtLIIfA5j2NVUWUZ7JoMII6E09C2zC0
Ewziv+nFVRfn3ZouaIkiCnmXTbWLHfXy8QojWmKohJzDSf01hG+oK6TuORqccuO3avm7v3vJcQ5w
M8T2CXMM8zGKhZbdyLybpC70h380p/BlCnODXGeCnjwqsJrVeBbbRa8SX7s7CIQTDC9WWY311NMW
QvLNovZuKVZJdHoHACVKs9EVPXomTzphf2XXrG7giqOmh0B4CHSaTxmJa226FTFqAlWop9zgJUI1
aG2V0fqDB1PTjCjKcqL8OB/laKdBdcqLVXaLxQ6Wtzrz0mAiOL+znBK49ZqiwLJc9Iat8cUHdNte
5RuzPISH8F/v7MAGc8YPe1j8uRe884OXX+rGdYFKSCet8zvNyux2pHpAdl5rLrYtC+mA0uZtdXVE
xwBRcQ1PGvv/MhZols6Nt0sUP8a9tSLlnADjJBzhGPkfc4awx8seRYie4jDB2WHms4jd43tCw14W
KJqVkoRsKfWamrECuHWiI2xwx+KjoTj5oRaZcAIzp1b0eiyHhvdoQl6NY0tCImAmcVkY8LAPMRQn
/9Jk656lzktN8v5YXl70I+fhV3NrjXBnwG7fF7ZSxUdF4FO0PfHSy56rPKSGWh9BNW0UXmk4nZGL
lfgswB6myUPLHSP7k2PRMkk7piFBfTUWfNjPExZUkEF8bs9YwcMOzQCF6lgo0pQGzbwI+RRUR4Ee
Mb8RmQmiRVa6umgywmn38h4TJNfgvm7Whw4H6gnQtOLpMG7d4z24p7eiCVJ6j0Im7NbJb/QzufAL
7Ezi0+9PoDTn+tFJLVTrgOW29vMwjgctRal9tHFdVs20QGaXzo4OJ+4F6Xr7oeIo11IGcC4ITGiT
VPw3vEnsVP/JkY0KYuigxjH1dt504tJzs3w2J4Cr37Y/GUzdNcFpTG47jB1unXXZJH/Jyd2Usraa
+5aG0Yyn8zK6ve275Z92YdXIR8Xasju1WW1eV0H4uvKQ+uAIWkcNUUc3ec5x38br2/O/spP0n9hh
CERgWCTS+SbauryRd8dBkmJap7ZnFA5m/0uFbU2JPMpcsuT7GhGJ7iY+laC9h3sxkoiCk5uaxKQB
TQ2VbApu+1yntmNtLne0KGFSAYM1nIGHgaUnOAVGBop7e3oolM4A1+s1bvS7NJPlWQ7IOtc1MRDN
QN1yJdGdeZ36gDZBPNbcONj7JCpReOX6p/QldkNPd3uHZZs2eyGw3XMnE5u/ECv6/d4t9+0Yulio
po/Yhhw4mr5QsRSy//RAHzH8mqTkjaNWcj4oDcoDBZYXALpsr4pXDxe0gVm+C6pYLVesNUUzutSs
O42kgPRoicXu4HaLUnJ2sIBb9Ui3eJEmkG0Zjs2AHJwipFiRrDwt/75LJPtOObBnzgQLz7GVdi89
MI52JGcTr0bFMR4uil5ty0juJLk9ybrIHZcb3wLWnt1/gATaroEWaFMNHbe+sQcqoUTQlDXa7sMM
/NZ610F25eR+klZDGBKziH1hWgvmnaEZ6LFEn1KX7MwiobyUS9kLp8MRVeOILQIcdXBGpqzMq3x0
LlwBt8zZ9Ilz3AXvdtXzJ4L+sxXYlk9nPoXYfNyvAwiw9e/mu/tr4QI744IN0djJ/bar1h8PRf/N
rFjBhT8bCZI3BY+bqUs+EyRU2v0zpkO6z+j02xcZp1GSUU47qEgyW/Piyp3GuRHI5MXiN8whaGyZ
llfcAj4G7ofALKbI5V1sj8ZOGmROSDkoUcg5jEP1A6kn3V8gL98JvvLa46OlMiZSa0KjbZUITyrj
OUT7s37nBqbS9Nf5LkX9Tx5DTsyl4nvSV9Qt3zQwy3SzTUoDBihwRWslI08VVanowJxsgjVRLA3t
DNji2hW4vV92TMuFKyi4GegIJ4uqAEi4C6MUkv68HH5d23GT2Er19T2VfdtuxJTEIlMMHdpGg6hI
u0LIc5l4EDRI1UoRhvyX4D9nZm8F+wpxF+5TGcN3XR60+hSXt7RWcxX8FVAFcerDsPnbW5GKBi0L
kf/IURh2rzycb/bFpVE3byLM6QyU5brJm2LUmjodjtuhi0zlFMvuor7Bv4lYfJRR4qzts/sgevY8
4dXTRMlgaGVwsWxt6YEOFPOGlCNm7dm4QWntOOjWOalV7ev53rXwJ4AFuKkk8Ua2fgOjG3gfrRKp
YeHjm3GGhyfWkTbpPfYgHOnbmQ5apg7mUnXecNyY9yCptlhj8tciO608V4Mwy2rmWWi1UfYqRVjv
ZVhm728RiTn81bNJyl74Gk9cClvC8JADv2uOms6Sd/rsbDh6qCJZ6RIkaO9Wk9W3dcVtPDY3IBwJ
BoPQSHTn9XdulTXK0dHlMrNxpNX9la7zQJ0YQF2auFhTQL7/u26+1cn8nJraIAbvwkkyhWq6sy4b
jjBL8GapRavtPm3Vlf9Li5Jrabw/axkIGWGNlSERd4l7B9YA+SCa/cmfXz66cZd5JJw4M4l5ModA
ttAcbd6hG/46d+OYyMoV8KHe3BSxtXxU5Hc76l7dH5sruOfKDm9F4i0+APEBAzLsWKkSPGxR6ZEU
4ThJyqRD/wSlgqMfOC733mntIiFrgMRXc3KlDHoS6nrEVOmQYZhD7bK4VNZFJSYSdD27jwkYMe/9
KTCRhUvbOsGWZ9oCZL/M/EJkvl1T5767xirGrd36aFgKQWhIkV7sWulLiDnx4cl0cpTjzixJYyB+
YMJFUDAj47YdVwpOq1iHD12x8+yPNKmmNu5eWk7CZPcd2Q/dUWnN/pyAhuCZD46S44A8djncQMXA
dlheUVWVKeolGsHODXS9Wd68LjDwKU4Ua3Nem94L7Vc0JEMU4TL/qUQLKW1VAUN3dtXE8wPDuA4J
+ITvtQiHjZfBrR04S8j51bOX20qt6NSVTsX8oU+vQZe3bNAkSYFrIgzCkMRDHQFub+klWL98NYSr
gG1TLEkNh02tzakrDTPdA3t/Dlr1A5gudID0WQlHfbuuAAP3WGuuQynj6zeYuQREAk1fXujrn89f
rWzdr9DQhLbSAMUxwiHA0A1voAqLbpA8pV8fSVINbNw40gaMwgkSsBtfDgX2JXfH42bpO25PTmcp
ALc7X8bL0BYmIgUGK/EjnBg6O/GDV2uPOG+h4LtXGPTdHWoihLjZeur/NlUqwowSwwvPKWUh8ZZb
ceQw1bTph5W2gAtrc6hnU3PYQNejYoyX/kzLE0f/KwqRmFzm4WFezaLBEgjMfsDiDFKtIYLULSg9
klSBEjnYduqLBZbtcQvobu9wWri8QEykeYDv8hC8q0lpLPjKBsMG563B8Pv5Nb/segMA9jRE32us
QDc4ib2Gb1peVzoQ7B3L7i8bTXED1pgosj9b4joB8Ykk4/Ktk3lCxReC43vDfzHk42XnT5PD/BnQ
sAbyvGgiUTBO0fVAsr6SHChNtCQePqyeDuyKTdJ0n+0hK+Hqb4hKkS7LBvIffA+HD4yx8vgt+kUc
+hVxZhUxA40LNQLoctzmgVSikh7clgN0TPPFfXtEyN7vieFzhZm5rbSJtukWbbGn/U9UynmbkyBl
rJh+SaeXbkRY4iL3caL1grzBBchPmWK0/YH9rKV/yUE2+hX3DpDGp1PjbqN4cfmwPEd8d5etPZ2B
/XwiuWlLrjHO/216fv56T2I0ZPnoa5r9Kkj3oxzno4pZjf37RgK0BSzqwoPEgJ7G5x2LOJz+engS
upo0nGX5UlB2pUJXI2vqm4qFuF0tAX/nJZxoroe8VabMYWovVCAztlRhjTqV+ql/ySOGKTdOVzNA
AXjVssmjD2t/6mO28dtxYdFXEktmD/Y0sCTQ2DFJNnSH6P0P9jEBW+6WvLk0D9yvlYiIXgnHkebG
YjSZoIoTUQRpblsB/WnCz2UNPmMIaWiM9pDwHeHmHZZacwf7e77wJ+J5NlFHxA55jA2gif7vdb+L
1169xQ5+mRPhxrEuyBYfrNlqxC+9bw3HnvMdCL/HDiUZAg85WmIqXbxNVuu9zsDx2PB3cqR9uNkc
cxkxzMhShSar1RRtsoqFKeLgHt+PPe/h8NbLjrPU/kvdKLKfnSF2nHusiRwbTH5UlsSX4i3kJwSI
YsjCljiu0PogUGORJiXGwi+3oac3Q84y3EzhOYFNuv7F7QTIh/hIHy9ONOI/O4yNlDGF4CBog7t6
eFdjKMLZ3YWAN+iQ14V+R52EUvfdW9/nHmeBXM0Zo8sUmVb3j+GdVrcQyPh/qIsx6SgK9HA836kr
k1Fnd8eZvf6q+aaKsr4TClU+TZgrHqbgGQ21QSq4Wyi0ZM9jGL0AaybDictlxvOnI+P7td7Igz20
WhQrWBDBVKyZklW9xZRenaB41eGl/SOTLKMXbw+pLwY+G6mbgFE/Hs8cCp3GgAgul7C8ZFCgTSG8
avGULc+WvMK4/prwDZNBMS+WEIIir19loiI4us3wiHPKaDdAJtHn1AkioLozcU87M3N8GKXHs8Yb
0jvPnPFR2QugezYnRn/I5Q38IIhi/PBR/MJhLV7LHEgKbx3iBHCCF0WXlqVlMJmBD4QaNXEY9KOc
r3GyVTUIG9aPLWNzREFy0HBifSA8ZGL5nbKsY5MTFLezxkHF7Hswzp6OsGNcVUNerY5nfIoTao3v
E6C1Q/AXyGaYkIZqKFVyag8UBLV0ibTtcdfJAJCPYVMQyND2f2selcwAoM8qt/anT1lEkPhyHlcA
b3E/yW1eiOG7JiyL1JmvMmYTlYzhbOa9KdKPC/d0IKkMeo94m+vdq9guCK5J5wb4PdIxCABjXHB4
gI9sSxqle7HmYJAG8wH1351Oxd3s5tR75PE3+AeFbRx4XiZH7+oWkji+/DxrCZClO7P4TR3vjMTK
k/H1irhU51yyT+HQTCxAM/BQQCDuMEzFGTTdrG/2+/ChbZXot7A4DpGhPCymub+azWyvHDkS8qSN
t96PvsuDUq2drPJN7T/aaX+XQ8eZOTnF6FaWzkctXHo6yQuPjAA1TM59o65c/n/zZUEJk994cpo2
GrBNOjdhvuvmsvmszG9j9QbxpepYj57SNfwnkeQ5ZubkeM5jY7ceHK0YC7lIw6BXONS3+l6/Z6kg
YrrqrR4SbcstaqQX/aFUPxYURFaGOg0+oj/Elq6IylzMCf7kahF1AjXLfWFQaGSfa8d9+UY6QysK
KpVxHsJCtToXw8FOA7buUguFUb4dbQeAvWmHISDy5pCWdbocRQXsYXk6TXIqtWNlcr/aExxPVqZd
IzNbT4o3mAAIxGYK1to8Ud4T4Oh5WpWkFg6N7Iedt/jMTOCc1EC1iK0IfWrqGmM2S0Ss5y1FmnxH
FhyxQDbqTborJVJYss79j2l/bDq5+9flJm1jz/LX6fVrxsD46/16+4dzJ/R21MIqzMYOXwPccsqm
bZ2KvEX03DQ7PIpJrTYizryQCAJ4/7+6bCIQ4YBGFpCQM35tNH9D7vRVzm3F6JmYi9RiCvv3zzoP
o7BF9ZlNX1qFRrfTzTTqm1mZnPozdsw32kayJBRpp01DKwC2aZmXMYiFLi/nEh2nvSWIcoodKCWL
kBWRlEzxPRLrZ25TscgiBcTvEBDI14L4oQndHUD9ZTOl+wKyLL4T3lfKs74UMD891+z98XoG11tn
jisdShvxRXk+k3FWKwQlrFp652+4IfAWdg8cdrU3jiZqS53PI0RBhiEG2ApzOjNp/+gq6DO3Q3le
uuZBTFtOh5gyVnQkAUGL3djdEyWrOvj72Zj4ZfPA78OucgYtGQKLP0Jq5tU++e7aVYc5iXrsbXj7
iYu5gQpuLUdNtbf0wycOFnk4mDC2QQo/8YW+p8uK41L8sdf4qe+P7QRwavB2cuIuBxREa7yLDwG5
eEyhc1Y+V3LgOIJnywTJPE/JEN1CEK8KtLLtefJKJEHiH/eNHQ6AJGHCeSBUTgVOf29fXe9k8ZV7
wXs3VPmbIk/n7bQLkz5XN8ZEvr41GG4E00eHP2SocUrP+NDr93/waQvweSFDmfacUGHb3Objx4gB
qB928sCYoLWyWsHuH39FoD+ZNse9iLYpTETJKRR1+kkahIIL/6sES168nDLZbfuxINONOpDzuT97
O2nScd2Xwdwrp4X2/7X2sE6kmxaJHTxZxIMoRUC7ckWyeI2s4cNyCv7RVABQxXrKxvaQBCqdM0cE
fKlqyaIR5WkJ+H3nU57uSS+PLejQhDLg/S+Y2ziE8aJWetkvtVEBZdJzfNF0n8nx/UPVtobMcMpo
p42cfAnWJX5rTdEjosS5a4+CiaADd5JUI3OKpYQbLW674SwDpSeUgwmBpxvY7NOk1cUiNzAFF3A+
NPS8zbKFQzM29KqTl/iGBwdjD5T+ZWigLgW8jnhTXa3BAVmDndvL31BKq6DKNlfLIlgXJisfwk7D
Hw6e2FT2gnzEzmGKjOhEYcqUruT3fpKgKpKKcz5M2dY7i3zbslmSXyO2I+65kY8ThR0o2n59l4T5
MEVudWXfbq0YFPW8NpIbCWNRo0jKFxtymVZf+JknOS6r3S571sKH5wHEZ75F9+GWgz/xLKaqZBkI
b68RrhTXBkDt6PYI6XCSZfIY5Fj3iv4Y+E9XVvDOcHeUt7yD9CjUSG9XFZeFt7Ix5ArvcGPmF09W
T8f8K82JfR3fGM+CkZG0CFA/hWokEaVKaFO/YTZpz2FyNewBWefYnopSeBK9MniP/rFqiPUlNcmY
ux/z+NAgJWW4b10rIbp9iiiR4hv2U8NmB4L+Uo5aTkHxcRveer3Tw/S+Fk9Mu6h6FwvFS0nNbXoO
6QtSeJ30PbpwdKMDdWtOXKO3hwJbK+wAcZdDje607joRuBPY7GrVpVcWmMsM5RNN9wnMosLtpt0c
9KMzHqowFrLgqHE8qf8lP78HS32yddyhYMrYtwHsnXwmjHGDKk5KeKq+05cAXKrTkg4h5lIgEaWS
isO54ElGVtPY1EH96/KHsXXaX6feG97O9CjhBQAuFEmGDe+QFp4xRs6Nq25TPRRZzfBaMH2Mw7KP
MZdL3KHB4HnLCO7TpoPq0ooNfAVSt7cxYXwJs9O3jmdU2MMNfj35YwlSTkjaJOUawGbpa0wUJdDu
Abe2OTAzEWhpRhwA6/tUxZ9hHcPfHX4vSOkkeF+nV3ad1YcOhSlNP1GnVsLoqkTx5shh24YV8QEv
O1kB7HGmc2GNKNRybgZL9LMShD/rWGkW0LKEml3xkTLYr/wRwD0acswlK6YOIqKSn+9vNfu5WY78
H/9mVkOXGTgXq3p6vZl9lpe3IkDhpw4TlDCYaF64NWjCmVzpNDtg9LiNf09lCfNttD9WfBwCdchl
skEkRrpWLipRAY0QQGi7bVwcUX84Dtq3lSMyhOzkjHM1KQCIpGNfUJR8jwE77bOB1OnzwliQwxZ4
RQDHlMvg/ZR1NRPoEC7rjtI/U3JIFsx1yQz+YW75hB8P3DKhShY66mUDuujBHK/hiMGOFw5CEZLt
bvGVBi/B/AoLbSIcGAfepUe3bj81ZLhA8+ap2lPg3n3qKYt/z/5pZ9iiVgo6fQuNhfsFBzenb5rG
BZXqmZaDDmTR1H1hxhSQnFl2HHvDkG0BWlCOHin4zMNXbq4jKL/eXz2AfmwI9e8dn0WP8EDYwfri
MwukuvxWmjJRt4wSgsV4hqic0N872PPvZ98QjM0g7VGs/2/9fPjmP+irlB/8qB+QC0wZWW2HvJL4
VygWGxu1zhgCB4+ZvVF/Dt0rTtg9k+B3MGTtl9bG0AGj3TyvoHdFhRlSvDITrLDvho1l3qfBVXtK
iBXcOKL2ecHNH7uNxfKJGCM1FeNJnD5ZuDWaPFk3D80iQiclDrvbRnian73Fyfa1Y9BQ0CWGACeZ
GLk+qzxixL3uhYaszTPwQRaBk8f+UKkRWRh9mg6UZ/PpMuerbWCzi12k+i9Dq/HyaORPFWvEvSYS
QctkI6IiPK/wlUpmIBZMEQVNxX1jd6iz/dcjsw8V/PlakZ38eoCKcBabZnYMU/FsRm/Bw4NLRMfr
T/8zKiOngRrK0cTxH8oW1zD+FVJJg54ZnwB9D81YlVvyykmmaGofruCRAefqlM65D21hF33lPuS7
PtB60wgZHIm2QQt+9hzU9RauqfNmSwlgGS2OMF72Cs7WHSqi0k+VRWZRJTUPPZnJ3kVn9nx2WmnF
D6Zu/NzDVa+x1fUNy3jm2m03uc5r+G+0Og47lUbs9ebkRscfsjzyGN0/8WhmZiOv3kwUCSZ/mvgj
3GWNhUohEOX2LN+rvylUEfavhkn5l27nhm+LzQzegTa5xWV3eZjc20DOASdDEWhTCybAXBxXg7cU
wcQGwN5sYaRljuEhkSVNnwRO/uXRWDZrnsLoTDD9Z9aFbh+xVB3HYzoIOSPIdFou8mNjqQB9ZwjG
7UvyXLunHRAuE8RKktdzsrK0/bPUKsUXkiq+/e6AGmzPr+cxF+L7tvpptCVbhXH3qqLs15B/Tzz8
fL3jMi1bCMVMlO72Y/Yw6uzp8jpt14S07whSFFmTrdvkwuJZpxtlReKvJ8u3VkWQDD4R0Z6sSB2V
NJy4Zf4KjT1w8sOpm13OZZA3u7gsd0zqUPJeTV35QfHVXmb1gLxTd6An809NQ4SroZc5RvjiITjj
sMcaJfvJmr6XbdSPPeUwPUP3dDKXOtvSdT5RXbdEq0YDwdgUGt/0H15cFpK5SgAMWWSgglY35JKC
1I6ZdqPeRZyFu2k4wRBAXrCEFQjU0ziXn2yivjcHBYHLDXdH4Fyiutd+7CLjQ3CIB48R04RU5kVt
6ugI0roPEA/bVuun42FZuzvxvt18Wlv4rxM4jwbmB85fw2wGnf4C6QeJM1PEsqeC4OhHDzkkxLjB
r5ti0k5MEsMzlahPYdOzI0wHt8lt044eIRWYn9Mo3LwedDfAqKGHiGfy3snYcR1CLgU8K/7C+s6o
HKtB67P80byzYgLp+sVoy5yoKRql3B067k1tz5fwdM2IhCnlV03FGjrfV3jdvYqE5FVdhW2zQ0ZR
UQUUJW663pbciQ/vCedkB/sF9Ia/78w5Iux27djGNuJN2HaItc5WtKkcJKKSsZGJfAoAuPIJrmbf
mgbeh4zWUroyoxwxFKD5Ijl/7zwpEWgaC8jP+DoqvBjuLk76u8WWnLGuXqRphtflu7+0idtsRqtp
zSz+OKAVnR5uAfbccKN6p790w8Z1FSBVStbgUNdB+3o5qj6wDohjWvDBGwdEOp2XKgeg1MM1znqy
4hBOw+3OyMEw6hO008PPJhob9sr10x3d5NPRyVge9g4qa5TeehDEYuHw9i1Se2JW6LGn9Yy1Rmp8
u9S6D9eV1ZQhfBq5q1Df9H1Kzdsoya+1745PpaMLF71T01nU6I/mpWiH73Nu1tJc4B/Ca7ZIDYay
Z6/ksC1NYTWbTg53airfe93AEwSfW3o1rCD2bdok7KfHMRC0vS2/2TSV5KQlvBSdM3psHHOcC53j
QHSYkskmwoY2n1SCL9bgS2R1o6V6C/+i5qdU0pQgyUztq57U7TbF4zsXdWrXy0r7GADruC/sU6SS
nMpmcLC0bP3qHFtrszS+kUDPGlcSdZXezTSYp6ryNbye2zMA0RBUZ/TJk5DiZ1JzaRjRayXfwSku
h5Amsrz9jqtf7hbfE3Nq/WTqwc09VrXMyejw2ZEGDPNVGrXNgnsQGZw9WlFPqTYtIlsQmMn5zCcd
HtS5FdEXrpcDT7uywEtRiJgMs/ro/Vxkh2fNkL7PpCfXsSYy6csZ3rSTKMXBZX14s5betxsPdfVo
qkmKYsEaGfJmRf0cu4x18IekyK4GbBEw7i0+2eY9bJ3GO9gdfusmyQ3dO6YiWxGQY+4P/Sowqg41
8V5WACcrZGewrd/uDRDYTQuduI2FcwGll3Req9g0GBETLFSG0WNtb8/7HEhPXn8VaF4DKvKYfcoB
8V3FW00wS7L4ecupNGv51lNdXJRa/DO1kX5LRK+8CGAup8A9ZY5gGAazHzvgQRMXGssmEZtQ9mXa
Dq61EgFJ0DNLVyglLUA8m5vgak2VZJckOyC3RgUZvWIsi3TF88u+y+frCNx5hW6J5sQPvGqB5SpJ
b0fRo1CoZvnYkJn4f8Vj1BJRwDRKlYZmVvtMrM9p74ZRhzahe30xbnLpt5z/yzG1Wet5sfAbPSXf
rXJb/SwWm2PlMkUWZwl0h5u3YML6y6uK7r2ixMfw9xX4QTR6KTVmxK+yFz/QCC1bVdUvFMXkkkQm
7As2CmwzCrQJc4zxaSZ+vo8QTSzPRXNs24IQQAJu2tJJY1XytFK2QyUHee2IzS+qpzuNRKDtOUlz
G01r6jhwEz56v8E3z523CKJJVv8zuxuQ4K2eyvPYrDmxlIQIO1cNh1v1fJchXQnNTbfeYxBb2f3s
O5X9kNRCi8ZmA3+2OtUj82BK12VSkvMvpFtaH48m2HycM/v292yt4rUQ5X/8Fp0c8bkwcjS8fdPS
bMwUKvpxHFcz6KlJo4050QT0Lrf/q3/aYRcMZp8uWqeyjbzwrbtM9HFafGfSEQuocUMxYHv7nvWg
ltqFhBrj6Tt5lzcC/Dd4JfC2Wjx+hghE2VTC8TrJXxkgvcHgEa80MdF7b1cbmiAFc0fGCv/1yeg6
LT9lvlUQ33T5hAx+oRyrFIgNosIrbrgrzTJqW8RFRyESJw8n3STW6jtbhZIh3qzE2IMJAOmwB5rI
HE2HkppdvakWvf76WZFYLXclAH9XfC5b/KQI2DWjd6b5WdoX7E7LVfdXdHyGt1Z+T7e9264g0dPJ
HtxtSwesAxJyEVdW9Zh4/i4PS00ADuZuSWtWwx8PtlT+gSmJxAF7m2y3PK+YXCtSdR0/6KL1Y52G
MTmByM6816jSAvuOTpPrIeTpHHSm31A248DXOv9xXL05HFTpyze1qbygHsuy2hWxdqsrWsX/eV8M
/zYxblNAVu/by15a/WZG6gSpacvHdIHlMS2ap5vg/67SarLEbh3VrtnOsGvumYqNinKmD/Hsi9jF
TQmh19iH4AUcRt0rujMJRicR/dVHqBLLVRQLmlIrHxOQzsF+doKv84ZjqBvIwln4rFZbNAa67y4G
ncogHVVL07KwobaL2ZID4t2Njw068VsRBjmxNqJv5UlQZi3UwsjjbtFMkxBRfTDmKB/2CPBWR2pm
Y/ERmJm7vKJ2riMwyPAS2G0tVFQW6nsrc2i/FJcjjHW8qL4MRdb4mBLFJtqNzpUo/NGpcKEgUNSK
jmdl+m8Xx+A2oCqmAGZS2VXxF+4U9V3HPLf6ljSK4cZA/VzUj96TX1I4h/t9ztizfeweFp2xDh9U
74nlkn0WZa6yxQphBzaI8yUTq2gvXJ2hj68ww7UgZqpuzICEdvZySwo+iCmpVegaiH4cbND6R+GA
7/BOnSkve5TAAgK3c6oZW9ro59w+wmemeQjSfMj7nfoaqSZRW5KO1SOUkXlC61f6qoiDaNnMCX1E
j3RzPf4NoLsPwCtFdkNAXgAnuD98wDg+l4zbxTCkbvX1gKcfroVu6KWYnrIIiz2w3F0jVhMZWI3v
axsthjDUsWgSmIpuawPf4TGrKZ+BDFX9vpGzK8XpKsbziq4Vcbw3dw3DRwsd4W4gXGiMgO2n38Hh
ElyZSDoeqVefgPSWclM3AGQBEDzO6orecHfKxa5+JRsoVX7pGFfldIkmw1mZHji68a/dnIjs3C+F
OE/v74jM7TkCGOfgd9Eqf05NTDEjS5xiXMs/bhq9QF/kA/vow931C92Rp+c6itvmYPBTOddwMR/G
bh5KriGhpWxq5SMq4RFD+dpMFrZKJzvzv5n3Nw8C2fuwFcG4066W0Hq8CUNIfGDZrfex4GmtEjKL
DB6krQMyXG1Qqbv3oBDtoZD1+j1DtQl7g9yg2VqFwrwWghMPBj203E+eHuAlJR0nvCXC4wMd/XgL
D1uvj+u5ojzP/wuYv3IN1M2N9IaRRNw0Ai68zRujEgABiBTFh3NITWYqydhqMdVbym0F+h+90Od/
j6rsVWrRC04aM11m2ZOvbEUQ0QltKPlLNF8dDb+xAGSLgzfbeEM4gXkIarE4boc5BMsp/LgqH2oe
MqMyx3yMR28gJ35kVnJT9IolJAMPYAkusNWtzQRkzyPjrLO4aeGCoAftWQLq0hnEJeXq7o+r+T7Q
UmHvGPkgooi7Tv5mVfS26DkFajkZI+0eNwAwZIZwskfwSPFTE5PeqYhyXp4UAEgNlQ1bQT8O1DMq
UD9edfjNSUVerGdJ0cXelQWgmomhhdvtE0KTrSBVzsFS7N4maLOiD8QrSbC4HDHTcG107JG0+n1s
4p7xeo+GVGqTU8lK48b1GLNTxNO6NfL7I9M8P7kDw1pF5gJ2XLAm1+9+uc9hqPf5Kt5rpaz8nsQ4
BV20LOrzlkT315ZGP2DM+Cnqe28w0ZojHikoEcugG/MeGH7PAi34DHv00ZtE05HzMgfs0Ves/1zS
HDw6EFEUeUnemSTFBv6WW9INKAM2gR763I2btUW7imfuRDP0DVJ395jPSx3jtHn1AvATk5FDMUxJ
yu4S+Bt+PBs6Y7iThMc4kzj2cm/51AlgA2PZKd6ujPXSu7ryneI1PJKZjENzRAf0Du1w33tQWd5w
dhofZV0CpGQHrKvTv5/hHCCNQMAbaH3zaAfQm9SQtYAhlZD20KDh8Dr29tygJbMGOFtbdVM+QVHi
huEMS4imeq10o5wyMBffhTMtU0N4dFCiQ/qKJv0LxxQksyLBliJLDCukaQW9q7J1pbOHFUVWLTQr
MQCmu0FvvnOzrocloApcVJR0+APDsHO3eIvI8IW8jU+w3ecG/YdyHaz6f7R5xLfEn8YQGnmf3xXv
b3o7Y3yA2h6f4H0GkbNLHpsLdQqmvatrc5t8R9+CdT8gUvJghLFlHzldO+EwVluBb2PD6Zk0w6no
660XQOheeitc5oCGcI4FydyNlbpbeJhyr6LDt9iYuRV8XI+Bj0ssJUcxO9IvNtGSZ/7qtVR5OtLk
qCfUKKpyTcFT/kw/pwg7RZzhxfERnnNeC5bvwXdZIUWKpRP0HXhUxFp92ZmXNz0ydtE/c6eaNlPv
azPxQtxnTkxur2pl9n1cMaVQ/tw/jUCK6Jk+kL6zmzBgfG2Qz/Ej8cmWDQGeiO5bmC6FUp4FiwAm
dCAKhnfrryt69HusyKbEevqy60m0Nsba2ehxxFG7AHOcTL8JkqHl7BU+e2upPukcGzc9jXTEby+a
BcdPGc+PIPxg3tD+tfTcLhJV1j0WfCLPB3R+7UBPv1gGsPDUfm7WeHxT3ARDclKO2/FwMmKkCnfF
uhZv4+jjp1asijKdpkgot+7UVtawMpeSwPjbnzHDtTbTAW2CDRo0S+9LPF9uAnmn9jIozVtwbE0n
l5pF1SAAlRgvRI0BSLNBzZBPuJbkmP/LnJbU3NFJL+tMqND8DKqixocy7pOQ5swrOlysRBb5Y4o/
sgqIlgObPhcqP9FkVvuJF/3yPn99O4lInZSHQ1dfF0jqb82NZ3hWN/2Xm0hyybVxZs7CvQa9entQ
+cFUTygFAW6UbjTQkoxBk5epU0cNZIsCmh5MAUiKLi2nhGHWszqBF1fTjkwfdYF/+GqdJAPBKIb+
vKEl8RSX8MvMxJ2tlC128g2flSpjLNT0B0pZryX7dqaq1+sShv8x6kfv+xNNqygNH9JNCyiu1Pu0
tcfo1lZC6Gj64ryLb14uUgpSFMa1L+2dKYP2+9biXpKylOXWJUN19dgN+FxrSF49Zn6rUnzQEHbP
IABdPLbmimvUSN3SrjPfgYy/yjlXTK/i2RdzWg0py6HkcWNIsM5wpayPQEdxlZ3yBQfhUrHpVeIW
oYKRxqKfcYpyDN+VyW6dRhrSp+Ay6MDCRDa6GDuWlSrqC20FZr9ix6MPpsWQPz55uc/0S1jm2stO
O81FVaNhxXQksz2jsUCafXpmcSJf7rTpRfzFE5nLcw8CmLbHq+ieFgz5A0aHsfo8KUOJ0c9IAfvt
E26QW0x0DBTzHFrvlPNbu5zFSqkJBO2KKrak+GPX4/9W06UD4m2/SA11RzBQb4tzV+R7nSHIR5Jx
QU1trwGj7OvSVfI0C3W7di/4XnlpQ4RQ6cYg6alL0Uqgjrqr9bBIXSRl/aDPqJ2lBr+dQdu84Tsh
l1bBSgYF4U7hmbKjBR9r23qTt5FrTPCbxtdPJ6dZrCdDUNydb6yFZ62Yz99b8F1LtV62x9G1MaWT
53HSB/kfgAekqvQajP0r4hM23ZF4bLCVsn0FhjeZhdmMBYX/myC43wlySmvTnyNE3c6geTHXwE9S
1DgFSvMfNEcNdyLnCTQ7zXEPq5eEjxRw5aGsnXMb2n+oaq2A5guHxEoKb/3J4yzyNgXm1vsxz6EC
axwshvv4jOW2A6JlIGQE7gj3+zCiXpL/3bEwDx7V2B0Js68xlFvOPhgam9AU2mzZlzYWoTX/6DlB
Mx9Q6KnhDTg2Lvfs7UBZS2Uul1JKzW0D7TFiVl1+LEVmzXlBcxr25xJeO8q6lZBD2JUKJdShVVKr
6tb/BjuHAQCRCcLUeHdFFEOHj8wPcT8pDr0pVkxwMTUrFGxzuge6lSVlb4j8tG7VwPn9Huc6Erhg
aAj+K1BcTfj/jDLktwc8qSB+rTz2oSWrwWAHytoxFLo4Y4EYbk9G0Hi7xs1SivBENHl1kmsL4kwH
GTDvzHqOsYWJ29DA/CvozTaC2R+GpHLjOwAi/8o/ug9ynbXV1HKHLLAHJpk7lkvXnrzaoOf7bQfW
qqjDNAAxzPsWaBwnlIK3WDYcLxhuVA59qfXcsJjPgkB/5lMLqacpTvu4+WN8vaX6kA8yZbTWQeBu
wsDNiG4RhesHgsM+fZihvG7F4ZEyQZZvYVG+yFsR12xSy/Uqryl5qKRaTAnfKYRkdM1Exu9We7al
04NP7QW8fKZqdPhUVLuZRP3TPpLTT3mXHFBGSQaccIfRewfVUYQ1MZ72NitN99gNb6rZ6lQWxIQp
s3tqYg+hfHV6L6xIys9ly8uBlyTUdDdNIaV8+sGgNJ+p2DCyoFpdyAOK+oqPmpcM8SHY4NlRzr4k
Cf+JAbX3982U5NXG6gE4UupnfcNpcIi8y5j6Wj/4IjuPozV0wM+7wqC0jMYdTQiGf2Q/qjGQDzZl
VLRe7E74TdvztieDvxSCi0jT8aj/uqHioYC9vDcvDbNRcVTmOr8sV7lyw2Y9rHVz2pyvZe0gnGVo
vnI76xcNw6vUDBh50UBNxrrFWr2agG7R24dgAmcuCZvvmyzeDYdvTl5a3AWgFSTnM2yijkKSFPMJ
iGnMGTZAhPEQxgsgRkAUXg/FXhIG0NNDgEVOmzlw4Vtk3CZypAblSEjwQPc+4DHleYFg4vvzk5EX
34H4rlW0kD3F42Ml0UxREd3kSYLR9KfdlCJUUj5HUN7jHiODOM4rLOjagT6Iro6GECNKILZRg9sB
OnM3bBq033aMD9x0hGpS8OmgPajmEzp/AdrkWBUSYaXzVZ5K64/p0sI/1CDLACQXas3DXGrJO7OM
2k1GRHx6Z8IzQyyRyMLtJQramB+hVGai/nbGirZtUz6sz3YvTMfK616w+wSXVVVtEgSjCEr4scuk
VbEtLEnAkS45bi2W6mq/KNw1qfxavW69WTJhEeDYx8UDSRYykC9wtOtY2XUtQWE24E1q04UVby00
GWKaiPMjvn68sjQToCsfyFXJ1feq6o0orjMTVCtHt3l5h9ZlZYUer15UIlXTnHNvF/5CkRENaI+S
0jNoesLC5lEV9YjWkJ+PCbbFlQU0GpbJlVUDbdtupYcVSFbah/cYwYgSaQ5hy7wZr1AiKnP8FjSn
pPre88Q6+5Nw39MITYf6PlLQp2i4aEpURwFi6GcVqQajJ1WEzPfjOjtSTBy3qm+UwpYWVWFT4Xcg
D2wo3BIMLlsZ7P+Mx1BSs7cAIUSbqJ+kUj/rn4L1qoQZcT6Hj/fB5y4Bd7+WSZdj0++J9YGbhRXj
frDvlAaYhblP4+q11Q6vCW3pRA/he3KGSLnEPL2K3Jt7lBJ7Fe5qWhiZAbAzpuq0eig9TJxRlXvJ
LuMaJlf2eBOgYVqNLBnImTFh76nVfYljftWmIj381Kz4/AcooAl6tUq3buAk4CmkTyovAmdEjE80
0dV6BTKRIv0FCvol++z2cPp3O9rZsjsNZgaRxGEMDrDAaURCQKtYr3cKdxrTLwMEgXA1HLb27OZk
55E+oNQgMhdA3PDumHhYfvUzn8ns2GLlRR2y9gono6NX+auvNdzg9ILMf3T+mquh+nYKslZku5yR
bpVQx1+q79zUkQA4NXaEsQEMKGgd6a1Zu5J1uDpyyLBb4yUc+tzYVxw4qGWuzfHRjTVLZFhh8vwE
NVdIoEClzRax3hHdozpNZOAd1wSh0J3MdhdFaoD+9LsPVKLOkXwLK4qrQWyCDvtT9oN6JNc18sPl
a60fccKnEeSmt/rfgXw/eHP0OvHsVs6XNwQg0iwnvzumamVyOSk63majqpiCWrAFEpkj55/1J4nL
J09tagVZE8d/KTIpqzAfXuC7SpkfWl7bBRAPQPeDlXoXbOgrGxm0/fm6SEY/9e5D5LGI7vl1bwv7
vVDo59Ap9QjDniJkF/2nZMRhykDOzmwaK8fD0RWLYntUdFtLnjkIZSG5P+2WCN8SgqZplyaDMjdX
SO6leDboKNbo3smr2FAkNWUDjVXRZfyPNFf3YscyinfxOQ9gF/nsCO4r3JIqNMJXcK1G4/6hcAiK
6Jbr8ZEqeXS0lBI/0d+QMsCeKzWxW1qTFRn+FMR9rmSWN11PS+QEVAGMYb52JlvLJJRmdR3eb/8e
9pX9kCMtaM+ue4v9FYb1rpfZZlPBeS1bwfGEPVREK1H8VCJWWywckz6yH/HI86IJkXn6IaOcbVA3
sEAB++5dYYQD9GrAXx9mi6ye6rW4vOyfhHtBlOlCi1CXvCzZPxoAhxUZ7bFMbvkKH36oiawgjnVq
dARRW9Ybri2FDbwWuxwtRbAx971wf6bp3ZPlRboFOtck/RlhTxJFO6wWcgUYd4KauC8ioLTpHYbR
cQheOoKXLgcZ9aF/9UUnZ8/SYGGEMknQYW9NQdLw3Mi9nfFgC7DUrfhunjClW2StHJApg46pVGYy
VQ4S56sdFh2zJe0wDqThBrnF/w5Q1ELh+M9cM8reJtsb6ti53uwO45k82zGhs5a8woJxlWazzcpO
ly4zBd/MmI1c/5nnvnBByEID3DTg10UYHmTq/yOpYjto3w0DfbncXK1xIL2dBoJ4JJnZUJhfCKSn
uRLXnjrDcpB+DitigPFy/x97L9L3B7PqoAV29XXj059olq0fO9QidqhkvcHK5c1xITKzwxzLIMEf
y7ROx1Y3FTOSJJt14iTbEDDZaYejfNM2Nk4//7NEJVZGsjNfl4D8lZ9vq+vVJg2xG02PpwgSeLgu
48T9hXx6+IOOA2c0TqDCx50AZX/hN26Huqjqq8hvbnza+tXz4o9Uy7rpA1/HOxBgIC4mfoTqevKW
/rITUHKoLa/c/Ae02mD9wiQqURUFkgzaxsyEGx1Nb5OIv3/wQC3jUwT1JROSNW8QkeZRJavn+1zK
MoHj02eWRZep69vry8Hho2qzdWdwFotMQT5dQf7hOXGDp2DLCuTF0JMHkFN4C6/3nfVDV4z2zuOA
v2o0P4NI3+eXkxSMh0nlI3soOfhWXAqU01pK0zeKz1k3XEUvGO6vZvn2bENa4RjUwCoLeEkIaMO1
0tAILyYfGZwhT9a3Phnv+xnoTyOwg3GbtrNJ+cLUNPqhc05Clp+Ug5K4xeCZBHwXzt1lboRgQUy2
BO0Rr1PzUuOFoOXGaPb0gwqhb66LUa3MjDCBrq8Y25I1VXIYbDmkkwVM7pnXIR+BUj3YmgeWrN0G
lYa+3HCrBoAhArW9Os+cutKkqSE7dlU+HXiyLH5AEzev8ea7qg0U0Kr6fRPlB6wUcya0Ed29MoD0
4Ie6sGVAKxmicclWoTv0t3Dd8/Fz+srufqZD+SIygbW44j0RBaYQ55+rY6ZqpyUi4OhQllts424y
u3lXnVh5KGaGCOjaGXwVQVlxb5/KxrgyxkvWc/PPkD5ohdiDeL5x6AbSvysk2ukw5Mx+0QEp12je
NaBgHilaU7ET3yIuUA0vLritmf4cogBKUEGTZ5ef+8LWOtaKqXOZU1J3qWUDfAVyZndHTaq/FFxt
2M4o0hnsL1hebvhy29OLXHsuo/5tN07KGEWtQKfYI/lgpF2rXaF4Q+1GtIra2lSuFB75mbfONJyJ
pEfVr6TuFRPjsrEbHuXHfqY6PgccIMDyljhESy8Ob8qPdCV5I51dMw2w3YoTf8Xu8V8qZBfkL3U6
vWLWnEQcGjUEgYxg0gE6RdaD3qGBHPBcUcXRnU/AgLzNqrddOTON/t6uj6E=
`protect end_protected
