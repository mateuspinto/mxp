XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���2�M�6£ZfǪ��D��	�S���Y����=Wc:������1�gT�Y��f�Cx`:go>��~$|��*���>.*�ݿ�;�[�R^�`ܙ�s`�@��to�b;V�'�֋�,����]dD3�4EF2�t)l�
�9,��>�._��̢����\����f��*�_��a�Ef�Er��6o��I��k޹���
�&6�����d_�'+��~�
o5�̖��)���Oh��6��-=LkI��Ly1�R�?3�B �:w(�v����͹���g�vJ;����~��E�0�ĩƃ{�<d�J_�;�\w�=�}�s��cϦ��4��ǎ\��������;Sd{݂��П%Y0����^iw�\YM���R�3.�Su���@�V�A�5+bjy���n��v�Ւ�lB{�
��p�<$�U
��\Tv.�
�vƵ�35�T)��f�<^S�F�ea�⻙r^���ߴ32���E�oa,S���.�p����2����GV'�p P�F!(����Sy���|�y�e?;�e^X��kf�D5�w�T��"�m� h{��3S4j§)�I����a�;O�tĀ�]k�YR?��_1j�' �Cᾭ^���$F�G$+����x�fC�q�d.Ah�_^u�ӯ#G��`O�����GcX� ���]Ѭ}��O��Ȭ���tÊ,��J<����Z?��)��v�3U����5��`��2Q$qn���=��� [�@��ʶ>�R�mT�s�YC�:�1ܗh�8XlxVHYEB     400     1e0�̓	=�I�4N:R?D[��؀1�|(+`<����v��v�Y�q�j1�Å�4
��2�@8���G��3�":��_5��@,��}@/�$.ĩI���b���ӽ�w��o��'0�E+Z���,B&u!v^�=YA��珒j��	�P83��Z��l�6SVy�W|��]�æf�?5%=�x[�{I�z�èY�A.�R����u�`O�@�ѻX4o=� ��3X$���7a��R����3w6���"0Nˮ���U���-��X*P;}*ά��hh2::D3Mܙ�v@�|�@v�C��z9�QA\��=����g�F<�I�vԬ�ө��ɍ�@=Pߢ�q�si�E>�eߜ;e�8u�?�{\4�~���)[Iu��Ŭn�x~��B�4'�s�ۺ�9��AZ�=�A�6���>T?�ŕ�[,ĭ�9��~�5��b���mԀ�dmґ���쮨���*^4ܟ��B�R�XlxVHYEB     400     140��Ɍ�M��3�@<����w����Ts���51�9���>�G����o�e�~:�_���U&fT�r
�x{��RAoQ��4��N��/	�Hy� �Q4�ְ�A#T?�P�zXm3Y
�uy	��V���-�]!Rn����d�E���/��7$�;j�%E���Ys��e�KkG=4�Fu�G������;l����p��B����1��%S��nQ��b��W
���qY���
S%&�����-Ow��A`��ϙ<�'x6s���^�}`?(���@Q#���������k966�F��.|��gk8�	H.5O�z�XlxVHYEB     400     140O��x+�:l�,;���L�RYC�aJ��rt?X#� mJȬ�����#N�	�R�/�	)���K�G�O�R\P�Me��z�1��e;�(Xv���g?�}���U�X͙�?�
��%}ZS�P�_�!�Cr;6��̲�����R5��g.s:y֗���:�*��E>T]�>ϱv�7���Z�W�^���s��ۮU�w�U�eN��}��!qA}��D����Ҹ��\L�,�xl0 �V��P�Pf|��J�+'�d��H�ȧCXZ���Wv(�X%%Ga�ON�L1ɶ����-��(#��QbZ����BgGXlxVHYEB     400     1a0�YL�����ٌO���
�TCQ,D�8,.��[0v������_����`��Z�ޖ�S�e�2�;�\7hc49��>nw��'����;�俳o,�G��������b�!��� �����$r��{a��q%K�`�����y�Y�0]7v���h�w�+�PN� ����e�e$��`�I��_��V�m8��ʕpjT���X#���.=3��{�I�t�@����x (�я�y
�O[�v�a'�Og?Y0X��S�i����xHᴪmcإ/�>8�<*x��'#��0�f�f7�R���22��r�J�m '�,��Y��g���j�^7L"���G��Bu�b�I�\9q�@GH|��b��gk#�I��A��A{�W6{�A��)���0���7XlxVHYEB     400     130Ǫs~/7qcq�~�.K�vph��9R�z�N��`����M�i�bj��F��R:F ��^��d�ٿM�G�g��1�G�w����6�;�/t�Ak��ф$>5�D=2Ԣȳ1�b���un���� �;3otC�gU�������)�A]�'��.$�x�Q��lL�~s�'��I��h���W�q���O�z ��Q���]���2G ��E�v�v��y�oW�W��)~~sǝ��w�V t�T�ӉMQ�y�o�S�o��Iz�s���إ!ë�ݒ��)�T�3
��3!��X��b<�:XlxVHYEB     400     190��a��yE�+��]'��rBpx�$�a(p��<�韃��fPl-ׅ�\qF��M�Ok���`��
9ج ���L��n�����8b!m���d*�����C�MU�<�C���q��2�3F�����S�7
�ቜ)��H�<.Ln ��ֳ�L�+�$>��C�DL�lf�G��a{n��0^B4+�Z��{�g�C�7� �6��w���D0�VDO8�b�A�u���W��Gⱃ�晞BBVY2E~m:�����ʇ�=�k�Xֲ��Њ�馝C�]Lsϫ�}c���`�]�H�G��܀ĝ�ƿ�Y�=/~ �w�w��O��~J*�l�����4z���$Axl���%��l���>k�_I|tH��̬SL�rڳ� 3�O�fr<H�������j��XlxVHYEB     400     160�7�n��Ɲ˵��5�g���X�uM�SV"�0�(=�[�5���B>��t�X� ��P�5e��|N���oK��|ɒp�+���	�9*�/X"+��=}7�o����ԝ���8�l�J�/��>B��G&�F���eN���FiӜ��;�4��m#_l0���L�s�<%����c<�7�I���V��}ݽ���O �vf�>��BW�+�1b����W|���d���9 ����چ�>���u6s��YT��j�y�=��� b���2��-fYY�}�v5w��ٺ�3
��"
!�vJ�7|����銽2O���f��Җ�3:�<f������
�����?�XlxVHYEB     400     150��-/f�\ͳb2��I�6�w��a˧S������$_��P� H�WI��NH�W�P���O�.�@s����$���̓���D1R�ļ������ӕ�������e�)DM�v������
!V|��ҋ0�w)�o=�<Y�	)J͜�i���z'܏��l	y���%�bX�ؗ����(�$��<EK�9�I�!�<�~wM�;��	�gl�%��!s�[�a?���:��{bss��-������¤�G�]Mc!e$3�#��q�ECt?(H$2��SԢ�GtI�4�F�4�3.#��s��=��ct���Ώv)�{�t�9G|���y�9XlxVHYEB     400     1b0�&te�Ѡ�Fܲ �l���s���6hʸ�ϑۆ�p����2wZ(B�uƎaI��� ���2q�o.x��� �0���Q���*��P�mn��g�IٕT�So��ɟG~OOB�N�.ȟ-N�/��k8���_��+�j�"��;v�ހJ��=���CCO�\V
�F8IC���Όm6�:D�"�ʚ�8 ����z^E��(��iAȵ�'��5"Q.���pM��i]�/)-�k��1��E{�dn���e�q(������U������n��ͦ�.�����������A|�OЙ��]�i��fH ͮ�������ј��;��g��ӗd4�y�|`�[��~� �������$Ij��>B�BDP����Nd���;zz�>^eR]�G`���if�Լx���@�Iӽz��10/�6	��E�eXlxVHYEB     400     1d0QS�3�d�g��25.V_+*���2���l�(`�\qf�@�S
�3�������ЯpUl�\������Y�@5.�朝��~�0	<������*�fОy�����_�i�:,����9�w���n"4*����mA�e�6�$9!T�!�}��yS[�'`X�D��� �@�5��D$~N$L�mY>z:z�r�e6�V�h�eW������h��b�F��1�E�=U��0��r\Bs���77p'�΃��T
fv_��>�?i�M'߬8�i-Y�m ��r�.�����r�fH�Җ��o�s���II�(�!���j���>�)���_7U�c�,�3u���YY^#��N��$/�,�"5���c�Ksgt�&or���F�S����إ}�b�/#�_N���4!�^:Z��b��vy���W����F��F����zٟ�gO��~��d1�@�XlxVHYEB     400     160�[5��3T��4���A�T�6q�`b�[Kv�_�>m��0G���|�����Q�p��O�j���A߰.�l�P�@K�=����#v�!u�r��l4����>��ԝm*1��ɼ��pv���*b�������S��UR
��,�4z���ԡl��[�5��� R-h��#2�/4;���5Ydw(}L�������4w�)W�I4�-�*Tn�1�ƀ�W��-��w¦��^QrC4�� �������!�;���kذ��LиD�܆bYo���f��O�����% �;Hpv��W�xTZ�y�S�V�u�F�vQB�Υ?��X��!��L]-�9�$k�XlxVHYEB     400     130n�׈��w�၄?| ��ۖ򭌁p��p&�(��~��ǈa3M!0`b�q��E��M��x����:ݬ�*���'���xC�I�W���-zM�E֝���aT
8P����[&������6#�r~�K�)���A��<i��>:�-{�{��M�害)~+$���aM቞"�Q�ov܆��� %��:�j`n)�i�CJ��p��e(���{27�z)��|�)��]����*�8��U�އ����KX�r8�L�ψu��t�26��nY��������f�sr�Ɇ>�^��s#9 *XlxVHYEB     400     180�j� �(Sj�M��e����)t��@�!I�W���	y��j�v�h�ߐ�2�{vh���ͧ�ɦ�P�$�3�.S�q��~^��&�|b��-�uτG��M���Ȳ�R�o�Ԇ�$qM����<�Y*I+�T�f��C�o�ףdaLɩU������lu�K�2�H�����"�}$�t�pg��/y��li�g��o~m�<��Vj.�~������T)���ri��+{x�_މt?�P3#��6ߔO�~`f��-�l�a��` �}����.)��������!�"���� ��PB0=6�d�DQ.c����@�E	���ߨI����ʓ�t��ޭ>]v��0sd�Rd���iS�)X� ��XlxVHYEB     400     150k�2��|��CbXL���P.����/0����11���B����u����\$|�Uû4�rx;Hr���zpG�k#�˫^pi>coHoA�x�ɂp���A�f�#)��J�)m���$�U��w�&�rjf�	.�>��t�����CWT+�����2��jq�w�.�w�J+J�'\��~�f��uE��2���x(���s�7��]���|�n��]��b�@���SJ����`�J��I;.�Y]��G�V�Anr(����-n�{��#D�!X�{�I��	+^�s����,�}����K���1E�&w7��֢�E�_Ф��-������XlxVHYEB     400     120���!�jgUNP�P���}��Q��͐+�C��n�9N�ʓ�ب m�K��M�Az���n���N*,����Kwx��*���>66�tHRP)&�*��׋���.¦=�O[�!	�Z�ZN:)\!����c:%�V�TN`<KU�j�3. �Z<�\}8�\�+�_��l�X�I��E��tY�?�풥:��hׇ�zF� s9���+�1h�c�~0��C�L �\e��#���"ܹ��O�@4>����W�Ii�,#"���7�	�0s�:�}�&o�os�qL2+�XlxVHYEB     400     1000~a�D����>a3w&������cT\@�E�����#���C`5�O��o�����2�6$J����U*���IYӜc_eJ��0i! �ˌ�vop�ʤ��$�gLG�j9���3�.�H!"w�k�xF��%��12����`��6ڌBG�s[V��R޼��&DN��^8��)B,C}W'��IF��d�	V)2$/Um�
�ǞU��46|0K�HEw����T3�Q,|�Vޜ��jx�+���� ���x��h�u�XlxVHYEB     400     1a0O�=��	�X�2��n¡�CZjS�����Y��j���X7tQ��Nz�_tX��(��1)�g�X5/:%�-��L$<��~^V���VfxL��Ͼf����5�Xa�c�b}�.��fgF�c���e�E��L�j�E��E�\�\𙸤up緰��T�+�Os۪+	S����/��a�֛q�Y��F��X�H��M,=�Z?ڎd��nL��f�7�]���l���(GЛ�u��v]���qz��x��B)�p�-�D�.���D��:Pq�E�HU�-)�%:��t/x������#Bn�o!i��b��,ї�~���ݪ��W`���4k(��PḣTbp�#ąV����%m�^�@����sډ��e���u�,�ByeH!�Z]q������V�U)�u�!T��5��׈XlxVHYEB      27      301��q��Gm)��k��u3��؁���F<���9a���y����8b'�2