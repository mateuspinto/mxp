`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
ltMulJUzPQcK4xsz7mxZjNW/8Zxxt7ZYm2oWBw0vBPmgjfB4xEzL7OZFrJeoZ+fJtJRlDr2SbSmJ
iNyYQkOQCpG7tecLRF47WyHog1luickFvmPoeGDdH4FrEluZLdBibxVZRBUjq4gQe3Yof1Kt30ph
MPli12HHO5aTJ5YKdw/qm+bBQwwb/2IuK3iKUspfVTSuMT2wPGfnwVkZk2YYE2TbWCE/6NxGx/KX
2mjXJ4ld7Vg/sqEdE05Ir/q1CGSeVzUPkJLPycnsckdmegHx4+/7sS5Dm6a/LBo1+viHQ/R8dqFA
s6GFbgGv9Ba1IIpgwTgDWSQfaqivT5ka5uxcog==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="GuEDz80mMMAYwTbuxD4wT2KjYKR0Ww76mro0cqGSm28="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18000)
`protect data_block
+Sm6U51yC9h1wUujKIPQMlB5hg2pZyVV19ItoRu/hJ/zVdgMtclzuJKzsaxa3rv0YUtS8xXo0Nwm
GZH+XeX/J86fXa/CuL2+sVUCH9KvpuKM33ESmWOJYL1R0LQmiYm2Um/p3GOOtk0XkwqlxxM1g1Gj
sHsBkO0CynYxv076svcXaDRhXGJp8Wpvs/B3mPtLI2ZgUCecUfAqbJrQOKq3d89Uio8UrTADp7Y3
PJcv9KJcZ9g9Y+bSFTQPup7vAXX+Qm6UeQOxwJQkQ1lsjwZx4TNEiUJioAb8zxjgUkM3JYoRh8NX
2/AKBFrEN3H/QbJ2LvpbPlpe/J6bqeNgRdsBNOQKRW/uhMJNSL4auB0a4dP/wTQostDRcIoXqpOE
1KblGp4tvji3vg6GhNqRjg03cZVm1Sdosrxlpx+Xsny8GCLVWXZZhvYOI+C65VrSynJfM7mVmlXY
i43w6Dw/V2WWJaK4w+I3EChB4f50VCzDtMGHABJJ6dcYZTgNRA1tWn7uldQ+St1o+8wXOMsOJaOd
AT5VgUqMHiqoRKnrU3ubz0SkoWi+avuD5ZfkeJg2uun0dv2iFsCKoVtqBnrRx+ThU/j5JhA+GWg5
z8p6iFw0t5TMwzKY9gObYg6zLh5qS3Ltqpr4USGMxcAYu18npmnSjWdcrBl6WSZV8sFHtPa6w56u
XrZVIfPrNB5xnfFBgmqmtrYu7vqinTbuiZyHuK7VTbrtzhjZZ2l3pz30G80cxz4vY0TwAs3X4MJW
0yM4O9kbxALKfaU9HTrOwPMFktL/85EUgwSPbbRg2UZBrhUsJmWLt7DB4C977K7zzzhFz4AYzKsd
sIbG41jkZK+HBJ/pIbokuTVrEjK0B7ism7WP0J3+vI61gDhV53mjrjtmwLh93I96DAYKC3XEnp4Z
K4VjwQZbgE436nNbSp6JIe+9gXGOkxKPcXq5/3IJzGy0TrDDsav2k5aBb6HJiJaHuH2XgWsOwIq7
tXrrCXQ64cIGRzOARWsa+9HWruvnrfA36DFf+Oktt1NQoDUfCiajFjk3LFdCtArnoBWKrRctyRtQ
zZhVrRw7eTU2MfczQdSzZfqVEZHg02vlm7P48nwPFguEixq1lgRmKtk+rDGFvTrDhMaulfKzLBVa
/mStu1ky65Kvv/bZ7fG7zsegFga2tUYk7zxfs6H7Vv473CX+ZfN74NrVtdHAGu9g1Pb5mgtNvIBm
ALHJf51dT+YsdpVfK1etQvaaf9O4l6jqlsw/tXTF+w5ufRUJyrcckgJIr8VzDPgI5wDRKvrfHpTC
BV8o9kQv377fIPbOdv4vJCOvEM7ef9BI9EybXmbexDo7eCMWyqodf5Zsn5xIHK14SjFtQaDs7uYw
ttXepBc70KEF30TacBjsYVear6mLGetWUfMcMNtBY8+lOhh40VzALJepp0YvuKDJh7RY99+oqZV0
8yNYdVdgUlmGlaLicsEG5SyY9y9AxhUwepH7/yrildKsyU5wijR64P4Y6zKMgsPAh0JEccjstA6H
qFd3m+kU+pjNmDTvR34OhVvDyQv0OTZi976BWj8WeKrcjQqWV9ph5ZWX684HuJmjf5nQxHj+Cbql
SpMVqxxODF8QKZhi/qkYqyBNoTpHPctNFqnCM3+LXPLmUFxO/CqIGrUrSXGX43sWvzT7SInVRDby
MtPvYF6EAardssIH1u6X9mvOGVZqns9NZu9C8I4wml8yHAppeLlGJkg+laZ+51OCEI3JKhs4qsaI
KYdC59O3/12/PQL+DikpxmGQRESC63oeW3X/iZj5YnphmhbuY89o0OtdxRIQS0viZGzv/cXX0ZF6
XwOLf8H1bK3WSE8C9ViVOAjwyGwE7VubBy0jI6kkwSqgL8UGLByb8Q2KHDkTpcPunNYz6dbW99ev
Ddwtmfza7oOJ69v8r78zdS9Yw2FVI1e+O9MryYPKZHy7y6xh0ZgB3XO+eLdsJYNoCS2lom+nifHr
G9bkZhaplk85DzWmfaexj6FEyVkytIttC4MBn9k7jHWxV4dji4Pml9LZSv2FIlZFKmlsHt+XnLrN
hWAr9rg5TueC8RxLJVHjLlTqERq0CLgVLqDtDJOKgCBqwS+ZMQMXGDDKaMiP46yNvMCwiN1Bn0Sr
aNETFmTo8xYSwv6fGhwgjH8IUVhJSNBdOPVVnL+PTq9wWh9nXUeHGiZcbnm22vcIPvNSpR2CqlvU
OeU8ByR+atK/zJ5k7zp/Hs7m4/m0BYfv7amxZd9x5ibiymxYmrymG/WofANOixSO1CaAJAvCUt/0
iBdylOh4SO+pLbR2iqVbQJbLczp25XmW51VcWKwjIR9OKYNeEkzt88sCmxZzUA34P98pdnrDcpCP
8cv8Gp7Biq+Ftf4wOQDN9vojO8ca10qijkG32p8ZBgqxAf8SVLlJ2BII71nid6B05HGiD1UpAVWr
dRZQHAJnatZvBxGfGT3lwTxQW4xgMjhYlnAMjVEFxoHH6HtdGiDHJbd/l8ks+QKwgREUPWU7bqnD
sA530WlYrh6ZmUDxIXbI7An36FGGvtA5T/7pStDaESltcuW/PyaYZClmxju7TOu164GPZHxh8Coa
JJcQEC4N7WqM/TcJ0i7NmrJcqHtaqTVKiCjp2BScq7HkRtNc88jB+tOjEx0rbJND0wXwmUka6eBI
nwdLoNICLiph+E2ecBrWBvXT4Sk5+2CsYbei9qFVP4uIKSZXB9pL8WJlEVNQbb+4v/xFQK86espE
qnRnUMvxGqBB5YlYXgQGAprTHIZAju01BqkORbSlMVhWL6y7czwaHyMcijfJmrDLnDiEeXcBpkaE
vwJ4QNBBmYrWfypaBGHrhPmBtFjZUDz7A+lfcnzwn2xxm+Jf6REJOgaIFVZr550BplcKbpbCRBV/
wlfc1UGEO2DF4qjvMW7PTNomTgRvXZNIn7PtwWVbgDPW8vJI2pn5uOmpeTR7WxV/4APGQl2JaLTa
6Utg3+bOvm0EascZg6Mx4C2S5j9+XXTDAo0mEcSQTwo5qgmqN0QgvdaKNtLJ+fMyltXw1OLm2v3G
pFlMH56oZEhkrvbknfbiv50zndWrZbLmlj81yYqr5vJzgMWNWS1Qg10gWPIRnoKQphnEevHdlTTV
a1x4ztvz9lnk0vTWyQKzv9YJwWfQGkwRRX3otcQ0MqSq/OiuD3PnXGC2FRaouUURfmaDP0FLhwAB
gN+08Md/2cjzCZT7RnY/6Nu2t6XLs6WLo97Uf2L2ti51UG23ehOmOSVAVsbed2cvKLkXaF+Y+eby
MXLd9qepTus4oHvxkwMNjq7Ot8OpasWc7U/fT/1zTddJzfy6uqd6AZPaYXzBaPwBSm0lMv5hp8V5
7IVxd5ce6zgEEvRc/NvegOia2HNHLE3OCoMseo4PuRSQggdU6dGMCv15JYR1DmqniPR0/EcNUUBi
hKuYCcr/SkHlQcebL0/vu7N9NBZjm/xaAmHAG2YW1ZW4cV+KpSTIZWmR5INChyLAgEF+hGq6olIR
Znub2Y19JFIaYPda7me3uhK+DEmJgOOpbHD6LCu6v04NH9ZTYEwuKzw8jHwbl8aV4Z/ubWVCtbH6
BNZb3BKCIwTnWobtvzjT581BKCvAGdm8kAeO7rkRyBjnX4EGh++O7ESRY6kGJ3AFsq7tZmvaq7u0
uzXTUJShoMG2qNjnJ9F/IdgViEnbA6d9M35mdFnW2eVyQpILOpdPbcjAhzcUlvu7TZdq+1fh2BK2
7wQVAF2dOeM8NdP4M45ygDW849jTQ1X6+UCZ1npAgxHpzT7Tg3oQnfndi2p/8ek9kYxvrVoJL3oz
PoxkDTi1JdjESTylHNmoP0XZHZk/OofPIWFGly/RsAd5xShn+aOqLBQ+MnPTzFx1MiYbPF5bb/WZ
+/u25503II7E/+FkvoFNQPsOleWzlMlUnyQ5x6IkUegH+OcRoXFznPe5PqpbgF9SecHWWN8JHHpF
pIhSi4lZ+65/pmrALUsvus29B+F9FwaVrWx8/8yLJBM0dQUGBoIYlsug5dxdxyNpTkDBJV6/lhmF
SvJXgVOzOLRqYUEM/rbdMBfr7be81wVBEP0ngrRgIZ+2o+CYHrZNLvwE8UIfTVaNZvl75Ccu1Gfh
GnUEISLjRHJFCSGDwxWv1f2MMvKn26tkDqp5NRGpeJncUgX/xlJzszVyhE1AAxiI3jJ1LZrQdnfd
m172Ka9CjH5NNvMlK1TmAYUlC4ktmjS+0Js18DgZ4YKi2wdq6C8n5puuT76sD8cIAuDj8O5ZpbwT
6B+Sz4NNviJu4zGi5yoXTQTJzBGIAM2bJ/4eeUUQHCdJX3FTYWbWnPhSOM7DCj5uZW0Fz2gkEeXX
93r8FvZX4EApeicI45Ue8jzm/+rtpQlcpnGv1PQ9X5Eu9KGpUCvFdGA1NewbSp+wHXuoqwgswef7
lxlzs2DjmkRlOsv5fvMxKVMM/R7h7dXRIqw/Xk1efb6bnNtsLs1I7RraejsyHDmoOs0goVHoNFkP
k6AogPbU9Er1koU0QgRgtUb0L2FL2k3pTdy1c420fx3dA0JlaVkcBfP9PX4Tybdt7fSLSDScqu+D
6b+DFU3THt9O7HdfbbdXGB9cvF6wgW6Bmqa8c/QvwCaWFixFgqMMJn/d1PNaf2uizC2vyu2zbtlG
G0RxG+/cmFQvlAW8waUvg6IgwpdaTJtJFGCfT9+Cdwkmu5vXC4mNjZaaPVpTlvuCUP4uimAlDvk9
2ilDNJ146ajLNbWoFS+7JDqiCKjSXnbfzIfq099wSzcxePxlwTG2Y15RI5ZR4aUfHkRVIavsm8cd
CUq5/Qzc0DeogPTbxXMVQj5Lwn0Q4I+nChdjki2a4k+htvvX8IlOS2all7Ls4JVcJJUMzvAX1z10
rT8lnoylb/MnpQHe3FREaN/PIJYD+bmg7Oxr2Y0av41fdY1SKeU3AemB92rcNrBoNadVJbteKrKo
krVK0k14DgWWLmTVLe+ZIHyj8rwXGXRpw4+X6Dejx1JP1kTdkymPVOABjEMsEhPKhmRtiCaOhkFF
Yec9mvpkpNk/8b2FAdEfybzqzxLidL+Q1spFGpt9PC2RZCyD9ovYAJ+2GQ3oPuH14kDGiaBMbMIt
/NpdZnFw4Fav9czZ9k4/m90MIuiPfh38dZgRIT3/YtrGRRUIj/KYsuaCdYJQOQDJgDesfubmyDsk
pm13Ubb7BbtFUdLWEUq30N86U7sR1l7b9S6m6v9LrMYdjFKDB0yCd79zH5EsG89ulw7t/Xo0tPWz
FZVM6bJ34T0zDYvaUjwvGaCUCVT1dsGgmZvf6n3AZoIXoMa9MwcTGo371eKZMRhXHP9IoWkFNVYc
P7j7MlAPau5oJPItBvHqVXN/wrL0NBRTRtyHhBQbMIl5W6rjbr9P8KW0mGjR+XPRHDmuhzrljbif
IZoqu2LPj7GXRz7VxOtQpu7kEIgAJgvn83tFGqy4gK9XWQyMOi4r+t2+kR0sgwwm9pcskLVj7XjM
gDxbIjvRFcoDlIubb9Usrs1LwEvchhqLP7yAin0mlcxF9fW3ZQaSEvoHkfsPbhEO0jH8feIoIkN7
HogTgx7ky4K9HuJ0zUgmve1JGfziO/qWVp0hsdbZvjIlZPJDcdSTYH0UhLMePGH6+7vDXbK/bSFK
QNG+HNRhw4uYULNQXS0+NA42RU5dP25AAvfiymm+ON1amwDOBH4tnVOyssA2Zmsuaj7kqtCE7Ogn
DsDSR36U0nfBLY2dbBO4JUQH/7b0BcSw46IEm3EvVQT/r0HgVJlH9GdP1laYP4JwPNagwqkkNIBU
OAYuEuA7uX3AtC14su+Io2BBRdMeUnXe3SFK4sPV/ZfBxGinKxDJztM6rSnmeSgK85NvRDkD196w
IrLAQ+b4Mt5aFLn5Hs1gsicvHg8MlcfomZR3+R4p6muz3I64SV2GOOa6vcirW4B3beueg61j36U6
DsE2vkZnvtbH9aKk1x5Iq6OdmXlEIkBsZu8zHLaDrmbJGRg/vgyVITksyMRhwvhiiTBF7ExDZEu5
PZrTeSfHLuST719DvL65NUhu6w92XoSwYeVHX74VDnNK5MH3y7UkA9hZiv3g2tKkrIgccDsp9ozA
DFdyBUWIpLxQ5FMAO3CNukEd+BSSW/FJEcnkTfDsC0ks0zFwi9+Z4dNnASpxCSWFFv8iXUT1JmWO
I1afAOLxqpkWY60OSgSVAJu0zlAxEZxxPxZjt/BRtJ0ceMBi1Hn0QzrrVu8Mf6bJuT0xhe99uy2E
Jo5f4fSULcMGRg+5A0ScVbyK9/mgjsIjnJaeXMcG8YtdpCtGYDHJ77MjBa0wh59gOPwTgNgg6Iqb
z8kCJaHFwKBJoAxzcf1GTuAzY76B/gfxx3y/i78fwlE6k6zjxeyT0hGXqdUEH3RWiAQE1+WMwQ6g
tOG66puUjf4I1YmM5MbXavNgYlq7lij0uHBMICeF4h6ykcqfPuj2wUeVTDlS/KhIVl2N3zHDNSI1
Z04OS4o1NTlCBikJKGD+WyT15sh7Q8vMK8OkilKjGfXy3XlxsenMhZ4E7TT9cPIPK26a0A7/I1+W
guJjqvZludO5zhfxb4rmhipFBgETeYDO/9cPDrpSnNdnZcRZUTR0Q1eoIRDoKqclGG0daggrO/kX
b0c9bMjrMoP2EvwFpfIiTSrOjwaqo/47hsBiIKKohuwgkqjjX2yN2Us/24osy7SrsKenDSPUnLpX
JKzKWvYQNZ2sluoM7rDIISCEqvf5+fOV2uxLnMhXx+J5XWLWhIbEQD64DHDY4aiKX3gjnKL0Vc4P
eAjqDUDDctk24iEY6/rKz1oBcW5TpIcXxjicdfxOboiaYumc2ZEbxCGC9fLbxun63sygS2ezbeWx
mkziaWjTSCCWBLk7TW+4C+zBYtAvxyVCcbxxXLZAmCZpxm6Lr3BddGfmSOWRciRKDM87EVKQTXeH
KtBrzh6KFJcwxcvBDpm0wUHxkEOvZHDX0y5ZIcHdAlC/moZ3uqDMpRG/dgzoBiqlVReXbisW/3/X
q9aM8VsI6cXHxH9OQyOh2iUYLUBx6DaM5beGMsLyqFzXLOXsX1txkCGa2cagOoCV7RE7hP6SJO9+
jKwA+X1ygNQgw1YHxmoTx1mgKK7J5f02J7n7dvP56DKd+B/vGNbT9mp7McivIozxGOEHzhh/FjFe
vcpZUH0ixSgDutAC+PY5zHe9Q0Nwdav9AG5eoaTLgeGRKe99BAo+BXqyH3H7/nq9cPVx5ZQesGX7
k4FhHgujVdQLZ/f0SIM6koUhm2rhkRui88R6EzCFI45OVQkUH6AhDo6tbDeC7sIxMrO2JzhWf21r
Isqt3exv9p6DGEUnAYcLHZzRMNNomR6Yi+PVirBv3GwPQT71Rf3ZMGMVht+abGqkJf4adZwKnJJa
IlxQQnLI5IQuqF85pc6WoA409O/GY1kca7bxKg5e6BJOs2f45g36HEirToP404SquOVJe6y2xOYv
VuRddBkq6v72HG/W0+V1q1pAlVF2pilwb2/HQFFoK6BXZKweDRkPyb9hnyybsU92yKyTElGKYWvi
9BM8tRolJ+0tMo8v87MQTOPGFMk1Cu2+GtyEhs0gNxrPNdCZ657N7kljUbDbnj7hBGf3js+tCIL1
E1Zy0eUVexW6V9NpwmczIeBUJnGL9TlBPNj1gKS4E8pUDoJbIa4Z4hIL1y24bT7I8doco9P6LR0h
9vMPIFhw4hsbk3/j4KcKz8/oFn0FP5FuNKD2R8rjf0ukG2XqfooNbgcZ2jtjKCbihD+H/hiwGl1k
eHhKvHQrhDtbTX9r1gCj8Hvp5PznGlxSE2JVIzMNIjaUMD3sRVp20bKtpCQB8ArZdivmcoH2+Ve0
0kcqJi9dRJ6FSB2hb9cL76hM3V8DhPgzEhuhubdMPbgfVC1GzvbshaOu25g+i8BfMDTdS66Yvmbq
lfaoJTWIvTTP3YHwMbL36ro33O9tRm7F9Kv/nOtVfSD1NaAYT2XNj4GVijrHmIwFjBmX2b8QqWb+
ycxREHScPYLCqHOAJbhZrIOU255n/uZ4B6wkiG4A3+lt4rivJ2IHWGOv9CLR7dAHNq5yYm0IRXbX
F08BA+6LASuEuvHs2TQxbuWPeT8zc+s3IpZPWZV1DPBXcQL4Ke/kLgKyHCzT/rCXFTJ3eTzEc4si
LpHXyVHekOkfc3m9sdzqC1VqIQcXniDnvpgCpMHLZYlBKf41PY8fKJHvh7MXtgpFIyrYw0OFjORa
pVJebBffwXK+LKH2aE7uYd+30AfZIKKO+97morESBw4x22DQx3bMKTWAWT5j0zwumeN/Bn8GR2B1
HjNtXq/faUdyMi1hG/lyFs8TiEQGzKmLA9zV1Lokbwzm+QqR9d/dav6n4CYHQdOQi4Gt9Yr8igxf
JmM/d6dJcDqBI/gjthabsAvbOxosrhi4ugmFAM+N+7JwTshHjnZDIuzcEsE6ZMOAi2r26YKW+Gfj
0rhLX+LZuw6O+NUQ215ZhK2cObplrtQ604yXml4jsLNhI4ZXSoblmQLjNHtD1z8EnWAseqxYi4qV
RwIr60dx3jMsFjqrkA4MR+yT8KRsQQi359RmL4l2SuY6iqgO+1ScT5YdVQVWselMUgIdugXu6N2J
sjvl6pu80SWEEJSK3rb+ukz2jGj+V1nnYVrCquQe8G5TWAZEAZYxt3SPv2Aon4h6dFAaaKCWQw6Q
mMbNjuBQoYkAXZosrwQrhdQRcaEKBb+R7I8SNmBHb+BoxcL30pUTHeesoBFXKr1msUMkfKDR9239
HNP5ju2ASLOpMx2oLtEPjWeJZ3sBSSvw3mYqtxwWvzHxJ0KAOP8J34j+XrRGMIHNCOkdcAo+8sOD
mbct7U97nlTxiXga5wiBCTGdSbczkSpPA8JTp7P+VH5lKaAtf6HAAws5XzeRnBG7PJpi1m1fgy4V
jLLaCjse5uksiDDJUG8wYGEav3KitAG4s0yMQtZ/sn2zg0dGYnf8Z4DQGuWI6H4ZXBD6EL7rC5f1
ZagjOG9uQmdaxTvQYJBB7GBwYzDifLsb0bgdT7vGNUnlrcxqJajlIrnB8Nu1xfc5RJRA1jaXyJ9f
4MXlGsKqYShf54AC0xdRifeJrJd1F9BJBX5aylsXrq4BhMmL5tjH7UWA66o4HWkc0uG8KXu6fpvq
doWYYYn6LZU9MOQan/jGArwOAA8gVgSEYF8qqDGCJQTT26kKkkUYhyEuN5kNhXfMh4SA18GphIm6
oSyv/F32R7P/yZKgEBjHnNYm+/IGCYLYT2sGnDav/HilljKlRH7Di7H5JOc8u/lOfcY1+UKMFNHD
ssoUUPh0KxuCvpO5zkiFby66I98LKa0pZtd/j36G3Ym0FeKcGoSragl8jqCeNa2est8HScNaGbgQ
jxhIDCdqplgM0sYt0V96IsDyXKJjICXlOiwm2Lha5nVZfKlLWI5es/vCj7Jk25mb8lqIgiWDmXc8
7tSW55bMTEqZ6inKb7JJ3MsAa84l6mYV2C9vDJ1LpBtHZmjfABPagmvoY4hqf5x5biuw2Zz+Lprq
IHCN+4cmjYpz6Nrgtfj8YiVXRARBFq1Hp/VZTLVghu0hfrgYjYPj/on8CqkDNgkpiAcG5q65t7r4
+7sfbCWwFMuPKoD/10RTPSa+ZrxhLE+MQTdb0z1GZuCWmFc4ZZxNsFru/u+y5a/GLHTnNr1+o0Yb
vMHX7wcPtD0Bh7j64HbttFF9jmShF3wPyJwnfarYfK/yBW/tINqlVZke41AS6TOGpv8AaXd+WRaX
yjmVbNHfRp/6J2bP4jcxSSw38ABBcmyDCxk3/WDufS/zOCJP1mQLYs6j1ss/QJDw7sIDWgyO8oVE
0WNV36ljREZcsMx6yC9LU8eARfsNNh6rpqR5PRWcp3CCCCoP0wBbyga0k1F1Bs8EF0n3YyKZ1ha6
P+U7eJqIJi9/eJ4mNH4N1iwMAkH5WN60mT0NVm2L2sGzrh2VuqinqlrxKg/xfTwQpmBwtvHQ9kXD
/P1AI+/qOqv2tOOiv/8+YVhEzykPnuhNAd8Lu7zk9G5tk38ied1QnVv/ekHY0RmxKFnF9zLSvQln
+EnIQn+VzwGuqzNpq8kAor4N2+sW+x/a6j/CAC8zKBDefXRSXHMlZ86IQK4eDMs9W1lGJpNCQ5Eh
aKMFma8YybZN4XeI6lLvfEi3HWNiCDTAMWkhVGNFSi/nFwVBmYHTUNRLQL1KQCiPyaTD15KSHCdm
e4jyTq/eI97VGUfZ4pV8IUisKGYD/pQfm7fjPN35O0X4dRrShpLdOiLYCPe8rqHgRt+m0jY6IpJa
+Db8bSmuMt+923O6b9MNZXQEzmUZj/wkgTnjeC284clcBCZEWpMDTFPcHX7Sxw+DeeZh5WOx71Cx
uioVYi/nwJKMhPEicVhd5/FSjOpZWMwXHR2uIR8vOvQ5nCqfmCGe+QxEOwydy8CPV9DiDG4B62i/
2hVv0iuy8oQkb+2LZvF6hTDKr6Ccnhk5KOJQGDud/lmCNd2z3BGwNF3CA3NEOMQg3hKx7UlCs5vx
oqz8wTtmEMScgTQNhGh86Yka+8+Bdnmmd3ZlgKQOsHkY8pIxziEZQASasQ2CKpJ1lB5o1ZWIJd6g
PnFwiblCYG1po7t9k/odfqZlq5l9mRLDowihQP1wBINsEh3n8rXsHcijOBF3jFVOvFRALRYmMrBv
Yqufh0zwHjKJiiu4ECY4GjAmgznCpHWLQ2DEcBSYA2/9NY5rZPteY+2/92Ak5QZ5Q38PfySex5st
EQCzNjBjDgpbASgcBy9GGYzMJZqjuyWLozCco5hvTo2WBXCYxeQc6Mxynnr8Zt9NAVJZbNL+PJuo
e36fOZQXuwVkmEogHN6ScsoncADrvZkR73kA2zspIJTieChYmgPR4IRqGnw1+ON1kupa3rHWN8Kz
vs08AQs7XnhHQGZpRjom4Be1TP/NXSvyYV79971BkMI/bHOPrhII29Lb86tP7EqsnrfmHkYTkB4+
cd8a9BENzjjmtvri1F+1y0qdsPt67IC/n6xAkNSVSzzNwhHzJVoxdVNw6rYO1q+1B2rW5Svjwl/I
A4fZjZHfekNiyS+EDJnUdC58ND8vsfG4YE4n8tfcUla+s6WkTaRCBltQdTBDmNUCeo1V/Jc1mhmE
OAVGAGpgimPi/+D75NOsIjK2cU19m/g1jFwuxFXitjE9LPogNjdt1l/vlNLh79URqUOwqIIFG0+1
1UR1xJg6AoLyI45ZQLfkQzgM3mZyiTAZf1Pi7RTiSuYDZdGqHibsjNWf6GxJB8B8KNd/4g10z6SS
pSWDaElXQO/YqM/fqAX4D93edN1qb9XAEbkmhSbfk0FDQbmjzz14hIyJKasO06cNOQD5SOlRZGAh
Vc1sUgutfcNUAGLqyGnV8XiepPkjD7egfr1nqRffazgyJTnuw/k5qz7gNKDYQD8YMT7ph+Xh7j0N
uFSms5FmfklqRxJsJW7CCSIZGT6lPHf7TS5AUvAr8T55yK6Ix6u31vptg68RSNFOp6fEDur1QtzM
kAH069wGEUgsx5cAjuak7RDQAJhNhWprZf5YnpdXpT3fdy9AApeX/IbbMGiu8BzxoVX495YMfQJJ
+QoyRFYYtEs/LT0FFSh3nQ5dCqwQ7IyUzP+01EOZnnCZ+1qmAVp7ysc1n412WRc3fT2b5PwdhQ7P
AJBci96HoVPZ7zUW1Kx0I+ejfc0WA0sJdOWQIreeL8RgyDRVYIwVOBd8StvjvExOF1ecLmqv7Q7x
PnYDGI9Tl+ZJxVxte886NEe1LRyHOPou33LmAtQyhDErh0m7ym0za0lR7JeDvPtkzMbJzD4CjqlD
Bbmdu6gEyKDFA9+M7fXhs8gsCuP44cBYRACvUT5eKXCQBt6xCgdWXWj6OPMlMoh0yMOICgJi8SX2
KjSHTju4a1gUtj+tXLSl1vnU5dayDo7/jEm0yEWF5MKrZaoifpv0/jponj7GC1JZK7yXjKhipdwQ
Ij3u6rZrapK/bpZ0vyfJfzbBy3IbFnTTnMj3KxLug7alp9fumM7MCSD3SlRCoYJ7+Vnsd4WRIWLK
Ya7/qoIhbapSMGcylJbJBIFz28kBkgV1r5LaHDkgRcPWY1qM/owKvRLiYcdDa92nuMVAFsGFrHuF
euf2rVzrNuw9uKbRjqMk9xiP1qsFx+zLX1q9xYpYPDFUdyW4aO86+/Fdvo4K5vTqAQXiIBb4zaXl
SdRZeD6OtbvIvAFC4H8I1+sa5jER/1X8SyczYSQPlSKjkseeQ9xWtrohsp+5amOmA21IjxrscgPe
+WU6mkdgPFVBvBHjbYDc2KPyfNTGcvpEStyV110N428iCYs20sdfgVplJhvB/xaJrHrGBHSBNdEr
7a1AeNWU6l+g5uOOL3vvD0tG5LUM/0AJjoxomx6G8SRCMvQQk7XfckYrQuxCbeSR54DQ3XUdFHVb
WtpMUwZDYalx5kxAObIrnopAR4ZIwdOXuo2m3u5Z4nPZjvHAjXhE3jQJJyWsr5LJ78TXreMb4KHd
2BYcu/Z0m5Cbqv4Sx7kFL/wOWeSq3+EozCIAUMae8sspEbB6A56/cE+ZKjbRrO9F3axW/Q8Ps8J+
+9cf1CPnoLCroIznVMR6QlFSQLN/ScqawLtSeZBzNdH7MoRG80jsNRSPM13KvO3vikCq00jIiorY
VW7q+bRoO9z99ds2wi4MiR3lSPh2x0Lkih9l1hxBd4AsnOQkNBzz0R+Nh8OzEcqPXXL5e1Y8KnuG
BMkkKdAbmcANDxPzfjEN503PJPAebbF28JXpv96xlEjb2QEdq0k7pzlTIxQw6HoZLYyTrsx+gSe1
CDZqXMf4kp9LdqdwNJe/UGPuW4H+6qMgmJZpQxlG1ZSnwp3ai32cchuS8AcLXqrXc5QilNlF5SQj
NWuHT6onUyYLgr8arZaIaZTb0tANtPIRqNes5TwHWSmkf8+Ij+jUGN/ni2B4rOmXD7u76MZ22ppf
uez5ExOQm4zMh7CJoRBHOTuHbO3r1yQm1piS95pPPiJmhvI7T0JvqRjohIV/BhYqLM2j0yq7oYlh
9FWXiIowg97I1IxQK0vqULRR8D2izmFrmUr1IprscVXQ/Ru8W2BWr0U5PlNQBtd7Cg0j/5KN1wRG
rraiDd3TEBFJHeGC+8x4bYKRPYM8MLQfUtc6+zLamPpXwvkRuRhVJVrCzhPfoDNg3g6q3NLtKTZv
BVw4ZO9WPnj0bJpgHjB7HuYFR2gMVpWRiMQocMLyMdKTjT4HCiYzdnWRbeZhFWInmGmHjXq5rpfZ
Uc3EbWcX4icuT37Armtf3sOqErxzd2sxV/KEjj19LPy2SALBn3mtmoglOgmLpFGbmF4xBHMuvwQW
+IU1SdFQJs2Y6tIk1oxd3I7eO7lBZEWtCp/A2HURT5RJT8FrWseq7E6/xNzhZxEV1G8klHH7M2gP
8omG0b4PJhkqdrl4dPiHm/2bQq4ry6Ntls2InmLB8vkITVvzYgfayALYjctp9hgzxvg40+QwvswZ
8lP01XSsY/mfdMvfHpGRWQxG2uufGotrBduo892gXTrnRLHORyndYRiKy1jjBGO3VRApskJSuefw
tepiOiydzdEYlR7kDZ0xLExldnDWiVpftdraFQpTnzwOjJhSytJavnmrEOu52gOTfn35RBPXW4PT
RTMLRdV4b/8uxCsAScDnpKyv2msI6gbNUakG4Q+KGVHUaObUK9Ozdd5u4cbD5vTP+r4WHQ0A+ZAM
7tI5X/2nmU4QGeksKYTgBKrQJ/jURvzzD+HG+ufMruqeeDRjFSXojRLuFUQOhcrkY/0eklqvgLSN
Vkfvad2q3fKhWUKNpgzQjx0Rb/seONkFGvjiIU3Gw0pC1y0MzGLQz/NXp35f+sSmr0VI7/0szeyQ
Vjdij9jIy7UfcvV+nR3UHYRI4pTGwphfKwUNRIA4ErFHfvoJQaAj+hK4QJA20RKWRcBxYj0Blq7s
+bCRh1y2EVGz2ldjdndb9V2oBf+GjX5l0LGsH8xElaGrGOUvC7kN4MzjfalcgL/J3E048631Lhp9
JIihkcbao7rd6PHZ8oSHBpo77zD+onIcRzwJxXUtOgnM3R6K74MNu6h6YjEw1I3A5s3/2rGFTsov
K70mdNMGgHOYbtgnDNmlL0t7/UVrKVUn9r46RNGeWwC9rWWCEDKy7/ONNc6rD3y8eAKlgqRPRpZ/
oC7VvTPTYC+a1OcFyAAbo9W3GlSjeN93AOfQOdNM4lOB4C3T7Fw6u0Wn41uV9lv35M7NQbEFa9cp
YAdrtnPppaWrdE+FT0+P2TtZICxa8dClYFQdAv5efiRFf5+Aouxv9ak2hmcaZ7NTHMO7sBZnDl0F
bV/UfNBvsuPj50S7/UyMvWakUhgImHtmhvhJ7stBIr7V3jICjj4cYz3VXm2SIJWMAmZA6EecfJ2s
dG9qzI5h6Q/z85r81azEyAPDtKwby7L+eK9kIdWCJ8lErYoXMGLM3tROMFnD9EPSNACN2nBU/f2t
pzMroD2gh5pO5MS+6ltVMGXNrO2ZsOb4FjxxNdYqpzhzf1aaSuf5gG/WnsgysmP7MIZvDUKu/IXL
CN96GH1t1rieAc3Fuvo36RIUkAc9wkMMYPpDwdIGWRUT6aaKQG6iHLvxwIz8rIhmb328zn6dAtzC
kRChrEeMrVb+p9YgqdO1mzqjaoojr/2l0vUZ19szuUiSzfoespB1fGQYu2OPsoeefJED2aEPz83z
wO4WbWQCeX7WPk5t3GjOpKepKsHI4d4+yPkf+8sCgY2yCzc0GEI2vjCFfekUmXBN4XOg1P19jbV8
LhW/1NbVdz61tXGglEMWwzL3TxxKbJt515kTajKZFu73n9E942/Uv/ExWRMI7ToavyWbQHPG0iwT
nhiuIM7P70+aI2/S0vXw5qzwFGsMNiabOUbh2hqVRBSniidSsIsC43DWFTWLe6XxOQJOm7zK+bwb
TUqp52X6wLHqJAUb3Ce5kv2LN+hqZlT5uEcJDApdY909NQnlFix3D4jEKcOZhca2FC07fil8yREa
O3DbL9vDRC5E3EisBpLLfQfOWWqUCc1dl+S1sDIkpGeW4s7Dwp5cECW6LNzBqdmCIbfvibG3UT3X
daVHER/qulMOhWaxvdCB6NqgrZa2YN8ctxqRSyU3YhwLx7W79mibwxliM9NvXpJHYPmUqZmZ2Pho
v/YKZeptkuz+nzgxGXjiPLWgy50hWeOS0TcvOOomxa2ZuYXckTlOg75/MUxKcaQhJa96PFnFtKJl
nUZu5jQexRqXMxKzMhPe/VXX+c44aiGCDGwZDwV9CCKlJNyhFdGiRv0u3KzownGXOz8JQpNWIXKn
25ID9MDxYzEzbbKN/nCbqd/WX5pZGocVV3lS5AB4iJnACMSui1wdIJTLk1eBpW5OAA4rX+OLz9KZ
Aes1gxCrRp36MIpTPLMo02iGjKhbq5g4Lc+yXe6pFyiCC/dx799Lspb9nr4lsRmvm41ud9hoYebF
FCkys7O0bjFEl0N3ebeFQdVSn/dKxfC2pruEkz/pvPmLN5B0Qvawk2d5i9ulypOfRNEuE5AogFOC
KbaligZvwD/rk6QXKYMRQm/9fhSmyy/QnN8ZRkX/JXXJjPPm88T4g5ZlKiD5LwIQGbcLwOBkNt3S
OFV28rjxI8gQOopVSiMzzWoD9Um9o4hfllE2i/NUl/mhoeadBvBT95+ctkgSKH9DomCGJyn6FfN8
n38utfO/7+h/VglDUsWINOPIWD8OByZ6SJAowgVoOgaOQI0uSAsk8cDwlZKaSzS4cuP8Cjx2YI06
FLaCEJrjoblfC5QE2W978D+O2Ztt9ZHJUOiHXbuMhIwsUM9HyqUkWEejyVJQn+9RvGwkhiXlLGOO
QKZuZezCwb8TdBT/BJR+tdImq3tzVgHTfAbWmzIMRVWulXTAvb10r2N/PUsDD2dr3knSX3V2K+0J
jRIvAL4FDpJzx0z3nWE6/e4QRaiBFwyw0Fy1tgyVl2yEkblSrlHlAVTjHW6zSMWqJTcdXFlTl8Wz
qpyOTmw1T4jf+bC5vRVAXbXJc10zrpEETxLeL33ECDadyhJ2PqZGTbHjoYCFCZJHHiNy+mbZaVKZ
gVxktDqJvm4WgyWr/nxRKmjHBTpl6g6NHC4341DhJQdG9Tok+ORSlIgUx5LtbdcFrwSdCNEaN+yG
rY855lmpHSF8UbBqz0kCeO+1f9laxvEa4V08m/boGZKdzDek1F4hk05e2KeUAFqr/Muxc8VvJv+t
dQrh3poXEhAedzHLz96lhyuITWCupIi4ZktCxHKrK7CAIf5TDzRBwc19+VwEBh9NEthMkSwDdwkh
seCcDfQ+kv7JNkBXVfWeoiLV6+BE4DWCsas2UfAqra3ItRMMCH95SvvflQWM5Vi04N+Ya6mGSrtA
/POfLf7FURgpaDrIFlhfYC9+kYIJG7qCh1EWeqZb+4kVoxA675v1EK9yt0s431j6tmcr3BmFLHRG
rLYqnJ1GZNSDAjWXj3OSNDhpD6XFgZ3MpOM40uyEQjDFo7+0e7o8UoJvGOwx4B4c9/L2OzF7DNQ1
fCY7pEggS/Gw8PF68UN5n0T3fZPSyVhnAyIAYKG8kaZSJLTca5o3GNBZgr020Iddno6uURHfg5/Y
2o+1ryYTsz46f5LX1Fedo0J+JtuGpg4+u3UCeO3xbm5Z0qVK7xCQnROUe94EWYJs0E7y8fdc5ZNU
Afhn3lWFUMSwDKIKpoiRieFbeJAaO7BWfcAB2NngIRzqHAn8M5c03iZUr4ym+xRvWPjYfBsEAwSM
UByN7d6HwLqDCGicyMjT6EySjGXv8BSmLXaOGOmRrURMEHGLCXzVe2kV1EQVyafy3lmxVE1dZ5/r
1mGE6Q/glAR52k5M/G9q2KeAoUKk8xC393HSIL+gjEIVLyo4Wfv8zjiS2zoI5Y7dnnWzqPjgKY/c
ZOMaeljHsIhjRTY8CkUXrXNIEVXNgJdx2ONr8dhNCBpsrnRFeBh+SfW6Hysr+4nuqXWB63Ryo1+O
Of94d4BrlbyI4e2lvLQF2rILxmqbo+VMPcNprHVZOnkVXhZlEm5kUwRx7HAtCMelsaSb/I2f3JJW
4heBQSqAMt+iRTu5djN7sijztx4mzj8P6KBZiLOBZo25FjTgi//VVMWtgFd98jt1KzBXRfCcG439
/llWXAzWkJxr/BGYYxIXs1WbVCtPopFv669635/VyJ8nTqT4odkdlJOFIBvNz+4CTeHdmm8QIKM8
CLvftsL+H5KXh72WBDEE8MEkhbPzsGQ6JpSt1cbnvw5FGwV93ztfKgpVIW9G3YCQLdsyLhoV9D0K
qTH5Oy8he4UTZqf8EhlEYfQipmWTsNNQszFdk/Z7HDqDbHVgmjmjChY+0aMsLP8flcQ+o3G6/2Xv
MYBNdaGiDar2RHesPXdxFDF3mnb5RXpcx58k2YiUy2n7K2FNSLAznCO27+hUVeNx88pVLcKeditH
nqRO9AiIhsDHCL9hZW+Gsm985I6fQl5xoBcYQUDR+HlsATqcaZazMs5EJiwGZGnWYIhLnDdq+vCx
NTWcpumNIBLzIoRDYYmiV887IJSiQI8VwenbOI1cfCFc3jmeFNXncQvtdiEyDv9eFyNedC6hdP2n
aMDlrkJnQG/K6XbDhpIfwEbiWGjXLWUXfyVwkU+tQgEbIJ8u9VHkmGojPt1JUTadSoDFXup08PEr
0/a5sSZrfrv6G4yMsL70kyISjYfak4Wsaz6IjcFypC4AdyiHisTjndzGsJz29CvXts5+BoiJLBQf
X5L0h7pbxHvoPl6w81hXPYGRA/7ogyDTdw3WfwNqdJtdgQVtYFhZG0LBNlfe1K30wrrq4mQgWFzn
MCdxHp1AGNpkgIVuOo68do28417nOBDLgFKpK5sSWwIW7ifTT0lE5nrLkMQDaNZ01+bbNb67JGSv
po+IZvsq443blRLzczh8kEjBTOp/h9IQhQg8gNAO+6GxGc14BjuS+1mUinflSAXLur5fF23jpAa7
2WZBz59qki6aZhU5zyIRjo5CKHFbssA/yooJdKoo8XNg9TuQNZExZHuGsBzMVauN6L/bW294THsR
q/0Gr9BLJT04nM0uRNLdGwTtimV0AqNIvxh1U6TO/6GxXLU27+1P30i84mOHBOVoJYoBS2wT37Nt
TPm39lIujwp665/bVhyilfwG8YIREdbG3s5J2Kfo4jnCaBzGp8TWXn7+FgzwZsc03ksS33XvkhKn
S+216r0cWXVnXiwPmnjVQ5Fi57ObX0BdySKVo0SUeEKw9o+61xMi3JHnJ9zaIkpXTMG+kYnJNe2B
pYR5+6Ml0Ar8zoGwtS3tl6EiC5eG435I9ux7nRDmzaYwlN/jTZN2MtJsQFDUNu6AdhKmUYUcCzs0
+a5YrSNiXTdjXorfhKIjOxzJ15OPa2pNIZP40cFKDHhgeSONDGXsVgeuBJHyIroj1dVfVl41eUmO
2DRzfdsgD0jpvaBlII2Wq3bck7nNbd6amrM6LJoIfdL+wEg/tUmJkVEJqt8uPOALxo+eZE/jIBFl
uYT2SbYDhvBVIAnIVDNP4VjI5TK8Iayn6YxkJIUbVefJvZULw96b97xlH3MvmRVXD2jAZkkIBun5
HCPfRgcH40Nhcox/oszeCov1WcdWFBwWenl3+V7suEJbc4BGOVjxpWPeDGFLYgxd0RCjk9+r4+rf
UqqxxTFsM6O/tZbpUkNYk0czc+Y3MNdxliXSQFBzRtxwazvuab8clqK1Yil+vcDVGZylIn+DBeih
6ivKCz005f7FyJW5aZ8XddsK2kzgXWncSi9sFe1AyH0XMqQWkcQqYAvhh+Ij0n69BMBVf9uVbKmD
nuFRF/7C8FGdPTt42QrOpOYzhk1RPyk369RsDiaxrSj/qMTkCDnq2yYjWsCznb8ZDlAnzJvgYGgt
C4r6i9d6i2miuFxjwW+1UBsnZUx3Zg7P7pIo/54Y2nM+qy4RXLLC09JlVLedReJFLbRYYEgVJ38K
E3PCX9NJQMIzIde5uZYTze5MOBWkG8VwZUh5SNaZEceeszOnKGUiMD5An3fFz28J4WnXspbhVuAg
uJFlFjdg+oj6rz9j5sa0zi3rtbuO82/kHBGT2aghEpZTBIiiIq6h138bbiIcycvQw4B4bxnKWCmg
rctj7Y8Q0BQWbtY4vfBAZD3a/nv8lj5XE0V/p7sIOLGrw/Pj0vhLEGlZ4OQy6fmYuCvzjIew5hDP
K8qDFSnuSPK1+3jZ2p1EVV6edNFVeLTUivS/j+q43vTJ4JlbKcsr+DXujZzOpT43D697rXSjI9OK
HCaQeOLYzE4esombVBfKd7u6bgw3160rm4/y8YFQ/0DVxQD/hok/bhCIxVvnlPN3gCmcdciDvSnM
922/7hspK3VW0MNazXhFvordXz36HD4/KH4ZhIsROEq96kg23t8IyqlnFmhCc8hcsbFEqUMbNryG
SN+Ta6NahqEXNP7rzGA5A3wtaXyJx9/domajvpdJXLQT7I+ZtoBiVB3HixvW0eE4z8YaAXoWf0ah
1+nuMqF5g/yjvneyR1M2sOJzagYuKFu+lwnxuUx8gjYUhaOtbSF8JuSOQ/Hj/OHUpkDP25YZ5kuZ
fnM/G41JEvLw7DzeT/+VYbvLeCvvWnh3daFrlstSY5GpJ9O/a8m96FQ2gJqpj+E5moEBR9J9brkD
1ILbep49BtYnfRLbRyxEEclsph9RLEu49ogUTghqkSAROWAxWssnaFyNZk5f3/3cbSvs8o2NnzLU
OBApw42E2ry/dqibd062tR/f+3A7lNP7t4Non6sH64OEu7UTNiPaSXldOZnJmgegNfTtoXYUxM4r
0W6+BcmRyKeGO490XxLaiHbIzyl4r9pPUs3sY2L3tmWe1S73+0t/NNzzYSz+sNatKofwIjl52Ean
F1wj1VUQf7kGIDYuAYYFr49oV55iQjeHRIen0G81eMUl7UWumhFT40Lx4O9WZl/9H1/D4AZ6gfr0
BhfQlU/xnn+V6m0UTwPxW7n4IuGVw/dLLIO+H5pX7/p4YyV8wDFAAgil0pfwxI43Obw6pDIkT31/
W1VXaHwNln/j+6j1R0O+tZg7x6c59aK1DVDtyzsNh0bn4ca5OhxHI4PLHkOZ0Ox6jqNAMzkYlffW
JGpATk+eM2JEOEbeXpp2DZ3yU2b7dAencrtekdrSPjHgbZcx40rEmpbW3Y+1LFDlUBpSGJfTjCN+
kWV5Zv9WjOsrZnWWG+QjkNPJuy7u1iVW2tiFDVHUcHoG+P/kCwcjaBLszkfrGonF21TCcpdRUfTs
btM89c+CNNKui7qQNv3rfUPb71yG9YrU0z0NLpCCgzKopI8EDqis/eTAbJp+EqW/SGjbWzAx5lE8
gAOPZEtOrOiD3/ks7TwiBeFe6536Y7uf7VDx7m23eC+vcY5aZc0AI7WQoY8wknvLZLBahc23tJXS
fCs3xgJvcSmogJs4xwUWykIZwB4BOVyYyXFVaaUiEyaGaFfXG2rrSmksw0K0drVpCpXnM1iMAFJ5
dWHw5Fe5K5H2II5HxRct8XRveMRDiNHuhqL2siashthmxwv96Fv90tFpfn45+D1UaAOnTuKxpu/4
xsdStDvjL5AZVgMZ+VNJpkVrOBzW45ZgYt9QU7LFEIg5iYXCvry583GlXVCoUFULae1/hPqFkAht
SMJpDpgxPIlwoGHue6eo8h9IsRQ4A+t5WmO31Du9DlREqc5zABjQqAdgdmQTY54Mmux3xic6oLSK
hKiTS9VIp9CO4HkH311wu4Yzc9D6/UqEqScFhMxYZo4SMReTRSvg9St6Ui55xNcoK/6L6uvq0cyz
Vb4LBrIdGFztjWqOzs2WM6vHZAnl0lZdLxnb6UrEFIXf5K9bE6W404quLIxaLq9dqgSX4H6uORiy
EZJ+mUmdfJqyRFIJ8RAF1mpaMMXot94spOXAGd20lIIAvMAgKkfPZ4oDb2A7oFzz0yotWpiZOwom
Uwge2PXMXyjkrHROD9AMGFm29GaeqjzvLR6d1Uqs8q+4njUpNq5g0KsZ5FCLx+34vb6QFbyFjJff
nUmkJv6d8KTN1ud0/wIqS2mO+q/o4GdmRR4nzcUwg9G+gzR5O/tZ4UHfl0BUMY5LYdErD1ETXOA/
iOqzrPBsv//h8tjeWSqZ8vhg/0W28cALwU2LGoZ80uNn5PPZMGCaAI3SMR6yG9vY5Y/dxfBjuLFz
43mjlX91JJ7gfMEF7Dm1OvWhmKAjCJKvjKLirg8gc6wWeOJUqGWNZqk/Wb6XF5sx7wdwYHDiJlRK
l4EjYpDBvvJ3qr701kvOb1/pKXIBWxhWx4T3K8PdMNBhTlCqnltH1/wyaJWacTOtZA+bdGYPaEul
kH2gXzr0HFNzHCLRw64nqy6ToJRB+T58eYhDZxOF0u1C3oarbOe/dV+nShvkgCxhBHrHh/Uza3Yu
gFDGFw1ReryMlkW2CN+Np3qO4jfUeNnSrebrKOZ/vc6Y0LJYuojuAiy//B1Zm2rv60KbYFzYJDrp
yiGMrWvD4PzQ3SX6mDcfvX/GVWyYBbnyJyrB4xuXHr1Ye1f//ZxNSyxLSKKYUFjzlTSMBnoy+uR0
cDIVu9hKKYF/R01cKqj5xx0GtwYfrrIjWM/FJ082giHaIzmWAevexnXp1HU57TuNUglXzF5CGNzP
ItGjZ8AW3faRPNYKWPBnMOPbo8dMX9mkefhB86qvB5iVECFBg7R0AUbrlsW5elYoTxZn+4CK9pCZ
a6Yu0hBjtbwaxwOd0pTqh9eeb9kbBhQnLc14uSEmlU9vL4xy3kSEzGa7e8iAWKRsEmFgT3tXHeii
apmcdmCOd+ELZZx5M3KEllP+lh+Z91somaLFp5T9j8y4WXhSSQe/twnAAV/q7a72A80vOFEp6AjO
wVo+DsCB83dFlKhi4taIECjmoEKr0MWkT7gbyJ0uIhEw5Qtamgh5HzQhEmSImNJqKNL7Q5vkFYFv
KBeOCWczKHju/NtmiSOI8ZHUQSYwEIxU0vqsg8fs6p7gwH9u9lYdyBEJbFaTJoVCy6XS01te9CUu
Fm6bu1OFbBDLozBUshbMRcnSh52K7nYzV1kzQj+29nC4Ky+G7Nmb8JAz5mDK+k61IeFUY45kVnSZ
VwDN1zS/Lqu6JtSFBvwurUTUcuvTEU+wPs+lH46M+ix7TGV31eFO4R9WFp+EwqRe60bXx0jZeiQi
6hNRssCH79UPZXc99aoxqeaD6vZBYWiWb3xMLdbiMkGVE9dUeAzxw5mRDu1vtZ6F0cVV5de9gKln
h3jgRx0aOArK6rrxXTB84dOkqwbYoXVlRGQb8Itv9ijT+KaPPF/gptuzSPgafMzcMNMvdZZquXDG
pcVApfcL01CPUxonRqRyxE1KvRobcAzLj2GhxeSD8/A2IxIgDNWGUOxzmzRbTfIr+nBbDuw7iDJp
sqa1GtZ0ebWy1T1FyYEgrRzw4iYXMNX46VpRWQ3GRM6ozC2RO/YWkzmI+uHZOdA7EM8D8nUu1Lh2
Kuh8wfaBfpakoasZu4FY0CKNuBt70PcLhNHxGiVoqrtNR7ljzdPC841oQroeUPN2A2cEuGM7qZqQ
1yvFmFcthSZzxEL02E6ynwePnC5aTc+qwNDYI337rwZC2tDY/cRZRgiZSSZrRwCTGsgOKXefe8lQ
888LgQWe++CP63trmL/Rn+1XerwuneM1juv/v2pT6cppm+OC4WN53iSzHl4x/Zxw79eoFc3v17O/
w8hSYGVzR62QPnNev+/b61Ot2bvQrRnT+OsTIT9y4QGbemevmnPW85FFfby1NFffo8f3/PsEuGQd
NNvX0kCNhJQHexXOvV0EIhLHrKPruseD28vUB3tXo1Jbg7a7RTyNGROBQss/UOku4VU2oMRK7Urf
I3EOriq+yrdRY0XZtu2WU5iSrKxeAmjI/UUp7q+Br3XGbSlh89CPYsxudlwIV7j80h1b2Bm/BLEf
H8zdDUhxGnO54OxbLy5LbxFkpitjzknnkv/JuvG9tAUOy1ZHxhVIXJyB0RWuE8mTrplnAsV0u5vT
FHhuQhvxiGMdpwQN7DQV6r7PF95GXa82kpAJo0SxjkEP0qJNhKZ7AlB3P3Krk+6t2d3CAd9r3zZM
YHfB3d7WG3Jgk1eYCnX+lTfvH8YPlidiVLxT6FhxkUmH3EqiDuhvwgOcyvNJtcM8yPFNvYpYbw1M
Ywz+1ROXuBuRMG9IhoFH7UATA5i66QGl3esnw2HcNYZU1JxxtrHY+M9Rfs6ZGIgdmssqo44qRd53
6rnntps2uOyKEjLHGysA5fhnWz3vMV1TXfXUjPP9GG7Wx5aKzGv1UJxLm+tUnqRr0rlRaCo7MWx8
QA+QyeDzXd7aPSfLrlqovZV4LcFGjuul3DTx4XByDJmsDteKfxXEFZ7Jak+R10wCzzTYHlFSIVPS
dbEnifDB7Z1m7m985g89IWdNepAhoCvYfbzbp/O2LSkXyE2d7za7lopxstEMLdISd4mMFe5wlNsh
X7156TT/UJfaHSzUtFfCSLf+PNVW/GNkL69kdaeEZVNYaU6bg8kFl1o7TwBbQ2ZA5Rpv/v23mz5V
HpiXx4kp5dctD4Y/0TwMmYlO6AL8Ua6bWjTYRTOY6IzwqhwC82CLG9QgHzEBtoLWC19S/ro/7Ik3
lNHMZOxUIPV+TIV50ovBMtZwrwbkPzGWi4hMZF7zoEOkEhuOMfajB4mUQ9+fLBo7/qaCJN4DIQrH
cspYDGM49r3Y/vSvxU0/L8siA6hl3H1/Tc7fvwYH7oWG8KiKOInDmyvsLTGWYW9wKJXsCdKe7GOJ
CKaBtGvCDkZ/vfmYeXkM4BHuWqGCxUYpvNvg+hHhKADsCSAbDZKDveiP1B/YTbTQegYSnzmawEam
9nlYGKT6lmCMSb8AMBMP64q03sHlvJD0iMEAcK/32lMKNCcCSqtbiKX33RzMkOKj+VvaydVT2yG+
6g6Z/Pw0aSWn6WIlK5g9/8OYY53lbjaN5N3+hO3lT7K7EW5Wg+DMeAvwfMOgFQma8n1cGWlxJMqJ
q1to/h8C6Xzf2o6Vcak7bHycG9RdIHd+/2MWZT9t16sDqMDXwTcKUYOLv2aC
`protect end_protected
