`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7104)
`protect data_block
OJaFm+21xZnAlSDea5llZz9S4LaWvCI0zU4Y6+EnqqGCsLVYk4WMBLgWn2fpqlljHyPEZbTIgB7+
FxFvlE2KulF4cgUjRJ9EpDPQmw9Xa9wS0DQWjyPO2IDDHBSyjvvag3libi5tgfTb204egMAWI7mv
kIWuyONLn4uykaZvIg+XSJREQbCCARb2yCfHobFkR1SyDtzkQTiaDKH5deqJSpogNQYkpQJ+uOeB
75Xo8zgpY7IEjcXbOlLPK/wz0Ii+V5+aZWCM01pzMMlG8tjA7FW9TrS/8WU+7qEv8eDLjRF9Wh3T
b6rWSwrsThyLdVIo+IPtrCqPxMvahy/F/xqXIvi2SIFNc9IpebR6s4+4MfmWBisi3pT0iGzWFbr6
y0TKqwXmOkjyATRLSe0cb/dzkSIbV8SvZImSgOXi71LysdpCSkIJMZIMd0E4/bYPk4VzTQSnlZUD
Nv21kMrFNXDihByVAM8leMjOvifAlCID0leKe7RaCFROp3Em0Hc/DZXiLeH4Xmls87z/7CMfflQi
NyGSqsp6bSMZqYRRAsn9TT6USYl69j3zikskwENx79FYjCW4aXjFtDCottnBp0KvYM6dz8i3ww/b
2L937Nx71FXKgXRbdfTpahcmEBc2a3nDXaK98qhxqLIcaJUJz7jFKLWDD9RBuUfNYACZQyX1mV9q
GqFlH6bwmM/9ZTBr8zPIDhqiLw/YjPDM3FNxsIMWE4WJ8UmpIbjFRx4rWv+uN2hclS0WpSrjW/1/
6QcnzMnymC4YNzwqjG6vN5GSRw0YGWO9ncbQrM5gwJ/zgfVHvyzsN1W634DiyW9LbDU/+zO3pTmE
KSQvXsiBEYbBsExzN82paimVP00ee81FmY9HCLbndN0resuzdXv0/SLuuFo5B4Libhs7r36nauz9
ouTOJGfJ88AO4a5x7VVsYUhrEFDGYpS+tjGo72ca2o8W0hnwEqg8Tsr/vqOz1TgSHwDavjgbjaNK
MNNKGLn23DMeqC2cErOXItcWuf31jckPY3JBEaYzs23niK2hjX8MiUkzzgDOFgMj1cBnOrAKg8Ch
1xRIxmduiaRCkF1rId+6poLKlnO9sWoTqAvYrUo5rTf/WMiSXCzl8xj5VkPXvG6/8cY53ANUqlcJ
cKjvEPs1QtYbEUMNwD4UJqsp+qa+RHn6s6jfvwBmglyeH1LqspZZaVJbfVQUUIStdTcKrdwiLOeu
vqp81sXcMbFSz1wLryKxWdzjLGb5xy0LjVrItnKEtFjZj44TM+0wYMExYs6Bgi+rxo05aIvG26qY
YWslz22ZLORg4jT6pvZMYb7qQ4C3MqUxIGILwj8WteK9cHFpU4ahtjVR1RwJIXZW/pnk9fosgUdr
EOPgiuw7iw/YglYlHas/tUlbiYyDT2U92Dd4SwzUc+sbwBdM4OGWjmq4YaClkUaWRHu2d3kW4NMc
Tjj2pyaLs/30j+87/DLuL/FVr9iOS+IoQvGpsS4kLv8PpeYppZeAQtoqlewPescuyCsGBxhhBisV
Wpiaj1Y/uyvUKO4JiqEPcKSufZVrtkvRbWjiXLQMHbgTNSPfG6Lo+uh3Azsuel3bn513Uv5oAgT9
0HjGd6UMO1VopaPvNHhIRgEAq983e3X4meTLIz0iXjQWoF437ubxdXOuPV8uR37HnnVpWA88kebf
RLywz49iIagVUrejMZQk/b0vme2HHuPmgDGxsVH5pecHK8kThuoCiNAwUmzbZvsDYFTXkfHQXimH
HvsV5Otl31VjquO8vaSZMN1we4co+P7WzCN1x5csK4HNqBnaEfb+0PrHNsNyZSHBy5zZgY+yFkSw
YI71jbO6M19TxzMOsnsXxZzWmzSXHCKWtkCpVAIJchUCRC8DcnsPrJS+Sar/C47XMLHzZAN8hSUP
MDIpdH/nmqjpYVO2AwdSPLszSRks4dlqnHcYLeuIN2/s/TrKfCBAvcue3hAaXD2WcAKocvinoFEu
3zgyCFwpqOM7H3WokupACWCx+mmhc9Hu/LZ/5WmHT9ZRNMp1/0f3lVeQxp1/JmK8WLeVQQoilFkt
K4wbnd/0iGZ6f0cn/AVt4lmsWIiqMa2GY+hvOdS/5uF+3Mrz7iKvd046jcIcZoemDhXzbeCtc2Fa
43F2UbnjQVESUuuVYYeSZRHZg9Z+mGluo/6v6mN5VFfjHpAtSc6w1w504DrqZ0Ab27MMX1ttyHHy
4XPbqjeqsxt3mh/IRHhj7gn1qIwIAMai8nri3I09cJZ7wijy5nuGWZipMz+sHez7/hlaM+c8Ph3u
TjGyhKxYWBOIU9sUlY7OBns3Am5wJb2x1HsrcnsP52zhzhuIn5adapItC8u7J3E69+LdhgTaHiTP
UW9NKt8N68MyPnRBfwlfMVGmReXvZV2BHtgyL0Syp4w1ss6+24wNiN6BMyavIVNw4XN/O9lJSq+S
7O8EoWuqyGBlzJWYOpzLV7c6RCnp+N/Vr1CaXHqnOU2S20Z2JhmKnkS3qP+uKzYqbowCbY4N6Uec
4uJng06xEDjGc/UKkgmvhwwUNYT8AyvQPgwo4/TQTtnl9jfEgbOn2dpyCMoNp1Ndr1EHg3NbV747
+gMWO7KvBEC2SaKW0FlyDorqAilpZJjF2smUk65qCdhJzyutMnkfahI0mBK/mg+jadQgkwSsqHtW
A7Y0TLoYEkDQkTi4bhK1XLWKXINP+IPU1oWHCfgpr1ys8qVskpZDlchBGpCnX6hrxCGCSXR/HHYq
E74B1G5645P/hMMjHXSNObImqvDWaVlfAHiYypqU0bwWGhokzXhBMamXIJgklQb+g/SfA9Otg5KM
x15UZcFqb9mDrMveb6zso1xbHeZjUJnq85Ma5SznVE1ViYvNPHQNn/qHYn8+kmFRra0TomZ3N9pi
gKZhbowQR0R7Y4swMLXT6hPsHcGA+0k+QJ9tUrulLbKL0TA59hYNooszxun80+rmqgu5Xz9Vd6Dp
Wn9neVntXQr6eNseQMZAk2d0Xd2Mmd5NUryNEINbGBTs0czKVUdnCoogQG5FKNN4kF5wR94sMtwP
PnE/EKE4iahpoLY6SfvfJZFBTzbTlVrp1acEaQL2fOrCAx3GqrByubisY2/B2bNK9hP9WjSXWlcc
tfn/bixJLiBmUfrS5Na8UEJSr5oucCbt3/d4ht+GB/OTe408FOU/ByWOmxCwdAfJS/I7fcvnG7U2
1Ox/cRwM+xNVLy+pGK0U5UY6eO3+t6TQgWBruanv2tk+mVj5wo9fmsGV1AsQ7Sf8TMBonrxPaV+W
sLkySid/Sy8QhLH7Nw172t16eMkpoiPhoxhixsVbbc0RDbo82tcduzwSws//4CacL6H5HyXjvLJD
OwbeOjMbiY49eb6AalqxX+aFUW5e8SVOw5/CHJktnHJKqyf02VZscBOyRKoo7FSf1Hz1Kki2y1MC
5WQSWj3u1ll1MBdMfsBuaFHj7cJL2APiWfesrr8TsOtrTwIste6pFxFgV2eePS2jhyQMYEkRsGpj
HL9F8bXvV2Iq2aJgBwUkSXmwIaLxLQBZJNZs/4Iuf9w/4/QhWZvL1TVNR9inIGWWtEmoyD1aujd4
PP2Ou5Q0dQRCHH0ihtw623ALu8rY/liK+MV04RxIxasb3KbByAFNoa2HSR3Uz8dqVb6gjb3+L58J
RvmurkdnWXqdOA4Um0FYrX1WppeOsZ7iA06Rfq6URrc/AwX4zuZ3+NIGc6lsngN0qesgDs+a3551
dB5B+nS/LW6u18Qg6Lf+oGdZptm52U2nKzcXseyDkfijzFCylwIRzsjuDxfMvxwTCmBk5adMPInd
+9k3Q0R2zyJm3GrwC2vgubpDehFMK/trSNt+Rhx/5J5YY7MZ3mzYXUL6sPG6uPnhGCs4zdlqgC1h
56GpdBnzT/nN6IkHr73T3Y+qy7Hdjr3eVNHsAz+jtS8qTyalu/UeHELlYi9RK5if0TdupviJ0lzH
o1Aac4XJFi3QiqiHAfA5ek3OtLCbQ4qIrvCWF49/BuTFTSsaJz2qc1HhXbd2tRgguhHkADqP430A
WP2nEpg7bvEXqMM0J/KPNDTTZil7Kj+HErUKpmwKmEiSCY8LP8Vp5bO/EcJS8zihZ5mRlATzfqwT
5qQJYOHW+oHErC4Hl/MZDvGXGvs+2N7ZqAOFntFma88E6mBF4dt6ego/yjWQxeaAHblfn3X6ObkA
/CSnDmnARU8RhBm0FOW5A1ii41j1wojA1PYq+pdCZqxa0tUoFm9QdDVssYx2sfKfWInMxsb04Bex
P4s9L7xWUZPKo8ROdQ3HAwLYSqSW/OiK1WTXMemwRXXfllewozTp6plRnVjW383GkI7RclFLmEuP
Xh/7NPveYd1blqVzISdvMAbSV6vlxCDOr4nM2eeW1tVllO08ijlfObIy/u+P+CnNkJfQPSfJuPHl
bo4mjuNoTg3WF2sro1l97A14eDAFQNsu43kQatXT7c/7DbLRP3YtSBVpoW+BUmhrj6rjLxiw0M2/
uHWW8xzLMOHW4u7F71x8oWoenXixuBj8Ybb1OluNgQr2lbvQtt9KSNfbF7+WTF14sXuXbKpwhWF7
vhYrAWtZ80gCFhblcVm63kKAk9NFl5lqFfdEWA7Zo32Qqf8RqHtZCjZtxkqt9SG+5V4OP2O6ulPw
IJIojuIy+Q7NTsMlhFA6ZxbcxnqRoYwhV41MKy8QQbPCA39qPb3ayTbvFwhS7zKAYEpKalrEF3m9
wVHQ8ZsTqkI1BTziA2xh5GD5YTaRfhBnIxkBbYp9ivEoyAswdtPayYcDBGkfJXfbRjn7o2UuWAzu
VPD3xUa9iOdytbO4xlJZxAN2Mm+2mgKmCAa7Ikc/fI4naQj9VyhMVAFBkPRYOshKWMiUxYMNz2lx
uNe6Aw61NeSiU7aG49uy52u2VHmOVlPqSkzbU+Gr2efbMm2z6o9ZPQ9rnEjyBvJsdH4+22lzopBF
VkCS/FfaqFWT2tpSoxfaZF+7nPEOZA4FnGWjF/eUzLyvVS7d6h0oMWZV3Wbk/YyUroQAr0kP2XdX
Mc2tDwB3e/35zAHxhL9KOUkhDlqfS8Cna896NsDXTVAHGIjy+Klz/jsI0IgUrGwTaUa7qIymDwMw
i5yKynlj5WgNIufTmpULw8+gNmWTB1tRsCygucZVOY2ugRUqmjEhj3qv0cLP97Ww9+VQR6mEPydN
MnMzrqiBERZWHFsJzPMeUa9RB1UGI5PwQc2np0UnqS3l45nWOwiNM0+1MwoKGSbcPTObtYrF8PhU
35Pv75bjmW9YUng+pI9YJUhJFT810Eh9Dsd/s08OCQznzvsP7qk5oAmNKKVCOnFIWb/kxvmwhiBw
slHrP+gmStnpRUaRHWdinL+xrvRHJfNwawjeClsZVpjMMWz6GcNTaZRpC0i88aQ6u6R8loHfZmeB
Tew6PTACpzzPD0hmNT0LxT5/+62ayJAr9pT39n8wJlctuPVztGe5qG8100XxDoumxjZ7iMq15Bkr
rtyJOoqxLPCmINZBrWzDDJfUuN0J9FdN/CwMd4O2u1GksqFb8tMIcmLQvmLjip23RKeG70xQhuKp
IBxiFKoGH9lY0baDttoRcSWDROwaUKm48adhNNHV8Wxo0NjzgeicoCjtqIWxhxLw4B2x6cDl2JuK
48xOdz6nxTTwIsm6M/dAoS/3oTX3zmciC1WO2jgIoplef3xkyLE6qlitOqgzFowWOdcQmK+dVEap
HW2iqKoaRJkDRIqFZn78IKd2qRcOBfgp/HX172jEPLYuBd3m/f2GldXeuYs0SAqjlhZvtAQdFA+i
U9uxxxPc9lzTL+O3F2LG8dfXm3r0E3MUZW74yK4SWghr8q/byfAMqvVjc/zHq4a3Lgwv7mFkZfBO
1fyEB+F543T1409tDSsKxuJRT1J/EUg8C/NSYPqBHHWq9Mb+qhCHhsrgSgIisoPofVAWcmu/NB7S
8Kn6AdhX1PDG7FGWmti+06kuqRBy9t0EDBdKDxuKqyusIdWbU2lmC6rDhn8/oKrmddE6Hck9M8gq
36B9iHUlbDlaPczqLn1MCbWsBM8cgL58HeHjRXufVgvxA9ZGQS2hhc7Cxxqdniga6U6D6T+a+g7w
lJF5JRrTuYZQwFGp8YAlAXHh/DtHMuhd0jnyEkHtjG+sHbZzTOTBf+mskiOR7EIGNsLLo4aYwshA
C3qkTcyod7vurTwU+EYYXZ3BUXsE4K6SBwaB9lvAE/2YjS2JuytFKEYrq9piF8BdwI6YUOV4rg5g
cjnRU5878DbJ1EYRhuuGtwPJmI6LPGk/oAJ2u0aahreC5rmGwOkZ+C1+1u7l8rSV4sSeNmqVdH3W
smO9ZVqylSPYX24xuShrdZGkCmxo+3N6mJY8WUvT33p6kWCNo7N8L3uzHkuA0nripr3EFSMLqON2
VVhGMHdneLCnD4NjsATXBPYfu3X1ba/gfwFuwXkeAXiSoT85iMIwih7eEejv4WiVv4rpA8CJdQ2g
W5v708GCPKspbMekW8Z9xy+dJjiyuNfLX+vdBkiXPg4H3dnQAskTDt2utFQwRawWrJTWRGs1S9BX
NjC0yHxb9sKbx5v2vXwxlv5QcJQbnk6nS6OlRsLusWlLJB2ACmKhjfrMKWxv7Fz5Z83Xmb+bSZ9U
T2leeVL+RC7vTywCQDEM8kipXCJ7ag0eCFefeCp1x7aRIhiFi5oOTdUGcHojHC+5KPt4eyXLZcr4
Pu77aQ2V236ny3XyPvtLG+sMTScSwglXe3lSsnm0VuwfIsVKDaVM09fgrIXewFxIsIRFuDmtZZIw
8h0s1HZyEppm7nAshL6/5vNVFTufMSZ3y8gjMWQeLsW7FQqdDDGYU28oMGeZomnYc88PhdhLcsaW
+NAJ166JIQo/s6rcfN0Ei+Lg6Xp+e6LjqngNJywJQnD8w5WRdDcQGeRcB71hf+ZSKDdJD4gm1dtt
w95zsc8b2wb4Jq8sd3lx1lBPZCKSC/Z+44gz17H/fZ+QP7q1rThiudUTkciVacMXGcsn48NkodCv
t1xpiO/vEHP0HIOwTz5bNZfkdB0RBfT2FovvwEbIBh704Au0AhN1PE272ambtakPXnUtM9woKnt6
Wr4T1lVpukkm/QEBORWU5H6H94LZCSF+QJ8rc9sPu4qT5Ns944HhWoI99tOrFvrmwlg8IB2xP4gI
gK1+oUSxObBbW1CLdz+5j/gUaRey0KIUyf0tSFYrGQGvjiwY8CPro2rQ3YUBSCyUmZHL1UQwqEa+
aaaBVHrOsNsOlobinZ9GH9quWfyToy0T94+LZpKtgsEohSH+7txENBzVxK0kkz4IE2MYExT40LcA
7EutHgaiA/zs+ifflGmgOXWyW95KchQnlodfsCDc4k7ZWiugtcAiCo6yGhJYm8kXY+aI5/Mtn1q3
bWNvDvpMQb2qdLh7ZruZbPK4UfhrBMqf+AZ1+kybG9oxq+Mw72eQ782XX+z+o9HjYE2MLLMpunkE
aWCy11QdfNg00hRdREVhX00B5goDxxaRfPmhDRkYY35emPZ0LfID2HXBG2+Uc2tDfh/dRDhP+94n
NeqhY0ED/92gcmBWDmrNRl06A63yyCmm8pF5d4GyyYmLcQYqMaJq2RyriaQycokDywUGkddKttXA
4Sdh00S/AZFT/Y1O1BsqOxyd2ZM1QQFxLkRII7xRJ8ezj4MfMgWzEr8prBBJewypF5QA/GY6bdTC
cvcpBpTUm0+syB+0lH/EZQ4Fhk5iqZOw7En5C2Y2QzjgnfkM7qbgYDhBhFgBnPhUtnnZT/W6yFb+
YJCmzv2TaOaNd928XvQxrU8WlSPKYljvfoogEkcSFnM5hOiUM+Ov3/eK4wjlBz8Tw4PVtIOlc/Hc
Fr9HpBt2rnFM1dwfePjXtr9fzfF1VfVGPbxESXTNmBfKG9cnSg8fOkScBqf094SYFheKIXUuGHy8
eKxN6jWlTlL6KiQFbNDe8Q6nlKTo/wH7sbvU9Uz7VbT1KekFW5z06ffhjap4L9nl8posFYH6EBhF
1P/uMWvJ/VxgAYFu+XOM8JyPe9Y3zcAryMJgYrBc+WB4rHvwSAyKvZMR3iDkz1z+T8rPVkCL3FBB
rSvFadhlcCZrgj6zS1ClKmbGSFFC7d9iRRucOcNVixPGJDwMIafzJafD1J/NO2hvPCcXU7mtD1bO
m/3QnbHWE9lBkVNkPHNwt3wEZXmTyKJhZUbUx72DaUMwKpOufDy0c/y5RP40/n3kFaTUL+b6epKp
Eu+s7ieugwr2idTSTfJ8QWk9h9iHt1/EQTgzOiBVQx7YxFa5B9VKij0vGwmvpSiemNlEAaxYV1g+
Cjo0XXg5S8A1RAxZbeO8Yf9ClmTTY+7cGOgaQKdjRotWR9tdIlRtA+09guWf66zkYT1cMn8BOzmZ
P1NooLy0sfQPBZ0kaLrqANTSb0sp6cJcI8D+LQWHoOSV30/qNItITRe5SZRH/CKBPVxuo17Iymyn
miq1YOCI6TVATFFTqTHMfI1X3wQ+Kl+SEQieygQvxyW1zHK3nhjjFPUeNTgwat/YamR04fVNLgRr
H67IHNx6EQfS9p/zqgfrPNUtGlJVIKAqjdw7dxkYOdKbsq0TrjnP8eYlKyeZNz36aM/GYdpMAq98
XGepQbBJESrjOn+OpQFK0YQTAV9x7+Ax8WUvLfDu9h+T+fkejLhHPaQT8xViy9xpqBaYzg7yByRy
YA90X0AURbxKGivf7w+/993ohjM59UCmDXcTV/8w+/8x/8KogrrKUlB0XfmOe/qHMQRPHWENaJeu
9ETIC1sg+L2+BoboHDEz1M9yXeDmxQd7m/64e9ewD22l+3fJeCEXE+1LqyIfZ4ojRH/lFXrdwEGl
iyppbGxmc2LuEoywuOfQ6t63akkXsW3mza4AjJhQ2K4IT7IAfulvzG6A+SM8hVslSiMa/IBaRWe+
mumNJQqkV1zsBVJso7KV39zwJb1cfmHOKafNt8xUxGcHsIyfoUBL2t6mQa7cdjxZQU2oPiJ7NbFL
lkeJ+EBdO9AyHI7lXnU4qtLOR/+Y/QUO7P51pcIWJAerJmT/vniS4DxGke8v0j5x/I6JUl/YKSA3
385erHskY6v+BnVmyoUP61/b2C/WeEH9zOOYKakuth17uy82HTM21V09BoRznu7sAsiuy51cgchG
z+62BPSI32U2WZrqsBaXdL99WEgnQ95ZN8FAPZuErU6GxztPDHIVSqYUoHyQq15eKe8JCHzwUQX+
QQlcwj1UxTrUnM2+36voPSCflXvvNdUqGdEdFWUuK+j8+lE2P2EvXnrDxOVle3cRtiRWRwG5QoF/
mtBlohlDuTBSqMjQpmLfNllVfo8D2eWXEnLSIZpabyFpQ/TqumL6VvAP+RGE/LuMNSiym4sHB4kB
XGLI34h4W+KuOmbMXz6XYI8j7PsLLrg9irOZ63N807BmA286LD5OBvZVcJd6lFGqk9JwasG3twn8
38o3UmqchUzzfW1AwGT/lBNLBG9TXi0D2cTTaJ8JRwEjh61z
`protect end_protected
