��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l�����¦`���B�B��l�v��o|O�6nXWM4u�.ƶU<x�D1B�B�Ȝ���80�[a�T�����#���I��n�˘��/-��zۈ�<������R��`�?aG����D�\�h�G>�`5:��A�����ݷl`�ڕ���d�s_#�/:lTo��E�J�]]��7�v��a��_��ghq?�Dh�ɖz�6�厲�YG�|�?�F��<��Y�vP5q���(������w�I�U�Z�i�n��K��_2ڔ}�9=Iݚ��!��o�im��%���u%ٓl,�$�jQ���tPJ?�p������	�q+�i��f��������W��B*zE.ՏՁ�O"�:�3�50�C��T��N�x!^�9i�x��?��$bv�b�෧�AY�@tV������!���J�h��4F��ja�@�Jb���y�eM�h�}1�W8V��&��
(�h�U��F8>����`&�`�$�͞�0�<��l�aF)㑀i��sOT�is&>��:؈{�"f<G�i�渾'��Y>$�K�Ow�����ɂ�$Դ�m�����F#l�C��,=tx�l��J;��o��I���۶���)q[�!R��qǰ[6�&�y������
�5��Q������1�9]�T>����O1�k��弓Kt��r\�o �*��T�5�� l��c+y���f��Fw`ǭ4���Y�!w�jU�����c	
2��*`�@ޡ�L&�a���Q�L��A����E��gӈ�P�I��, E��A0V����2��\�Q�s$S���M�����vxaj�W���#٣%%���M׽i�PN�ⴡ�#�t���m�4љ��-��SW|�?�ʔ5�yc��*8!�h^�U
Y�bQ�r� 6��p��Xa!�҅��⼉ڮ=m�h`�S�;9:�X����wr$�DE�����
pP?߃}l�#n{,���j3ӫ����x�&�m���g��+� ��D�i!�&+�Jy��rE�'�c���̹~�v�\���S$c�(U���2$'��3��=�}����k��� �U��=2���&��)
?��&�/�5�x�|�~`������ �cO=e^�hd�]Ch��#
��?����Dt`���}� �{��OEZ����Օ��뺙��K[�������q����$�}~b+�g���.����Lk.���@ +G�����`"�]7=		ȗ7{�ॱ%n��X4��gٔQ���r=1��#w�:���>5iY+?md���EN���|��}�ƶ/���.�,�Y����Neҡ��!_��N��z��Q]��� b�<6����%�+�����1��wS�!���r3
���Y���f�zv���yVuO�Uo�V<�R�s�@��?���3��9�A��l�fm�0?rkI ��؏Q*,�����r=c�7� 6	ժR�i������`��\�C�[|Y����>�x�+,ӿ�G+�/猪,����Z�9V�U7m9U��q)QFN��Y��LzZ�W���S�W����IKcY3)�A�a��!k�ĉEu=D�-�N���^�����62Oizؒ�My���Xm!�lX��X9X�(dE���v���31X�p��PV�r�	��WM?�֖߉���ȗ�}_oby!�P!��F�&|� 0�N`p�F���7�o��I�!�̡䵆i�ޘ(�I6��S�&����k���ĭ5��r
,��e����[/���U�����	���" �ݷ�N��<w��eE��ܱ=�T�dю�V��*��q�?�< R͂���T#
�#J1Ѕ�B��6#�?[|����.��v��t�(�2�N��T�!�P�p������V�z� ܼ�h�����}�|RK�aTMn���P= liRR��d�s�n�y�y<�z؈�^	�1���ɾ�|�<?p�1f�(��y@L4h7a�xKK�1�]�~11�i�l���z�ȵ2_��l����lm�r��K�%�z�S�%�i� ��M��x����0U��\��ȣ�|)/�;��4!]�F����W�A�������c��$[�R������`$1"S����ub��#�e�w��b-n���h�Wؕ0�O���}d�^X^��6�'2f}J)����!ޢ�BUL�D�QJ�O�ⲏ�R��5rB��mG�����`K�"� /sYF�"����6�q�����L�MS)6R��p�$nO�{�����4DLY��XLkv��0��*:�{ �+���	,�Ġ�v�:������u�����u��CnR<����=b����t��ꥴY�=�uk�g��-)���f���*q�N�-8STE���o��F��V�C�+40MM�th�s��$�p��y�]i�L�7�`=��\������ؚ ���X]�04���t`�%P�TP�JBβJFB���m�O�]��oo�e

����Lr���+�jb�W.�<}㙁?�}")�쥢�1y��Hn(SU���H�'�����b���� ��A�ć�5RG@1[Јϼ���qV!�}Mg(��\��_	~ª��W�H��i� �
�z�z��e�����?�BIؤ>�*9)�Y'κ�"��^�b�i@��*ŷS\�����f�K�(N���_���H�5��P���Y��<�7������t�֯Vĥ/��ݤ�W�`�0���G�f���Z�Q�Y趱�<*�w���K7V�}f�Ϻ�H"��b
g!ui��wX�ZNZ$W�VE	Yy���h�˝8	�t*��!���U��ƺg���6բ��V��[
A)��,�a4�Y�!��w|� `y�k��FTrw5�4��S)-T�.��jC�������YAZCt�Y:��62,VV<P���� K,��F*hN����*v	�J��a�1���E�|'��6�V���������E�0M�\�R�����Nc`�;�CC����ͯ��?�A�y��_p2<�� ���F���.t���4���qv�O >��K�h�H+��͛����v�C� sn4RC�r��U�T�vF9$RY8jү����b�)0?R?'����n����%أ�ܘ7c�c)���F�ﴯ�����@s��<%𛎇��Eqt�А�!Q�X�G[�jk��(�Xe��J�x�Q������LeB��Zpk�Z�3�)\?�[{jc�NHg���u��1���<WkcF�3p�mb�O@���3�j��-7��I�0j��2�-�5�,���'��U�j�d�(9)��y������}EQ��5hY����,�1ٻ:����!x�_��U��ÜI��u[X�l.���{�$,H]�n"����2�|5z�MÒ��ƻػ5�)٣Y���W�R��Yi�Ϳ}���a�oZWq�J���F������OR Q�|�)ұ?�.��)��lNbX���)'@?@n1�|i
�<C6�0���\�5�S�.��C��������i��l���HoL��'a�~Y��D����Hb���U.a����[X��XĿz1���P��@B	�}Q�
!�ͽ�����]T���ͦ���ۀ����c�/b��(q�)������9�z�#�Ymi��D�Jj�յ�"BM�������[iʐ����(���Jz���y$�S�0X&�sL������,���J#4�;�m���Ǵ(��a%�����:"03����@dIN㜁����f�@pwep�ᨎ��#�F���~���c+[/I���8}%A۽\�v2�'�Oم�LT?�1�Ns)RC���iLmr`A%�PH��N�")!� ���\�[�-"Y��U|�T��{&ԭ��J.�I�X�?X�+��V7_�:�j+��T�V(�E�(��6w���/3zkp��.%'R둍�bJ��4/���8��z_q����qB������q ��[��$����	Շ.3\e��a���Ł�;�P6qbԩ�tt�]��^��kB[PY��g{�p�n�I�l�a��t&<�:#�X��v(�
�?<hJNC�O#!���ǡھė4�5����͔D��S��'S߻��u��)�,f�u�6�3�N�vo�e[&#�����o^ޣ;EӾ��Mi���c�ۤ��d�p�7ރ*�h`��>��MrZ�>��X�;�C&A�e�f�I�� �3/�	Y���_o��+�=��u������ݚ��{{,i����[�\�HuY!D� �|+rL���+Ա̶B��s�i����o��d�Rj�n8����8���[]��ㅘkya*\�Ϳ�+T+�ְ:x���!���)'S?LI���z"Δ���p*����cݥ%80��e`H���M����N`L��劼���z�k�xe���V�_�n�"��t�w<X>����ֺkx��ɴ�r'��2�R3@69��|ѳ��p���8�&��V��V��!��x�SF^�r"�Y� ,��ᵤJc��9�_�{��T*�d���)I�# ��Iȇy���0Q�������,c� �i��{�L)��0���sv*:�a �`����5�'n�	?�fa2�r��hQ�ji��+�*�Q��]%����+�.����a�߄��a~��O�?�ӵ�&8�۠�ʑXv,0&�.�����r�t��n���[�b6��}���b���m.¢��	߬�i�O�Q�����m7n�;���*'�	�2�m<�=c�!�i8�hv��?�<w�G ��A���B,������E"2�#jI�	�>9���༭��B~}G,�����7�p�,�9{EIa��;�͖'��v>N���0��?�1	(:"Q�uA��Q�̦�,=�a��W���޺�o+B>�sQ��'D����0ls��D��E�Ȧ�	�D��?�-��A\��Uojg~=����}߻��Aq3��8Z�.�E�$qOl�������T<f��eu�m��H�h޵4�$����<�en�D$5ų@3���7�ݚ7��Ċ��e!E��� ��Ox�[�bQ��0��~q���c.��(��ic�i:�Lc��"���o
����
�"���G�.N>�w5�����@a��C�'�h�).4���Cq�%ŵ�0�b�.��'J��Ӝ��|Cg��V������f-J��@�x2Q��M�m��dLg�[7|tw��m�XU/~�R�P�QH]����by��&���Z������b:|�i���d�bփ'���8E����;��7�_�����6��V�L(L�o��d�5����1jo��;?R{,8�)�%�)T=.{̈�l)FTR[���\s���H��6!�	�\nO��^5D�0\��f�?�7+�aa�P�ec�d8��6��E�ң��KҘ]��'+cK�@
@[sk}f"����W�74�8P�8�Y��^NF'�	�j7�j��T�HSy����|H̬�ap�-���]��� L�D%�/(�|�Oȟ����|�>�my��)����mE�jȤ�vy�ր�z�/'�f�6O���R͍���M�ϝ��$�C�&�3b٥��:W ��H��9��!�p�_�$}���4)A�0��\%Y����]�qa�0 �VQ���|�F�֫ծcp��,
���̇��&T���IYQ�W:d�4�Y�7��~9ɠY��HMua���M��#r$[q'�Q+Yi��!�#�@��-i��i�#��ѵ1���{ꕸ��d�H=�m�17#?	����x��m�x0!�eJ��S@�KJ��͏D�0�M�r*W�D��F�E8�۳�D���bRJ���+�0���Hwa��5�޴r���7l�G�]"�qUR([x� v��y��$a�� ��k
y�&O"����\PO�Q�]�U�<
�JN�R������k�e����L�>_[$B��=�8��0֘��8��ac���}��|�}/��z����|8V���:�X����ܝ���x3m�B~�l��s�I�G	��0��)4{- �2b)��LyZ_Rb�d�>�������=v�^�޻2>=��B:Zz�# �.xl<aq�w���:�m�q#�������d-v�</ʹ�),]����#tT�D��}�sY��{�ᆘ{ϯ�>S�4ק3h>�5���S��8�a/J��2S�����n���c�=	tJ�����f袔���8���A��_�Z	�6�����f	�l�AP".I��x�B��.��9�YD<ݫq+�4)�p�Na"�+t��?�6���c�O��Kr���h�Ġ�1���,3���K��Z�r��z����R��_��9-&�/mZ�γI�����*]�k��K����NJ�2�]��c���r�¥�et<��=�b�"��C�\u-�ڍ#��XJ��Q�v��f�R�L�8�'�N\j��^^��q��V��S)�_DlJQ# ń��-�IЦ�U���>'�,:�:�$�rZy�֎�u������}�9����k��xd;&���<������۾T�dY�S��5"r ��/l�Ѯ"�It0�s)0�a���|�<�
 ӳ�]�$) �����/���#�Ņ�Ś���:3��ˇ�+��ELT?�O� ��d,��k�5�<{�6ja&;>���
7z�\4|ߑ����s�q�*d�,����ʭ6��r����v�I��'z%P����z�H��!�ą��J�"�f�Lï'�tp�v�n��}�e���jw�=ӻ�{�|.{i�N%�Gd ��V=8�#�R��)���'�E[_)N�]��Qk����NMf�M�?B�&Bc��sO
$$r<���̀���z>� I�0��{�]%�ӈ��L>t��~ ��8��Ym������N�%��ŋh�~x�6D:��8���7���@��LD�J�X�ߡk�Z�)�%蠳w��UF��ΰPWB.V��^��I���9fg��j��E��|yU�u{��Q���K3,���6t]ׯ���w0d�	��-u�B���?s8za\�*q婮Qg��5�6@���(9��5Ɩ!�I7����ݷ�H��O�E��]e�@��<o��
��iU����*�# ���f�������=xu���Ÿ����VƄ'&$�T��\��	p_��_��p]�N,�w��3O�O?Oc����y� �ac{����V4W�%�۹�n�Ն�·'I<�!���.�D9$��W'��|.�*������(}u0�C��2o�ʃ�I������˫����"m?�q���I2 ϛY���l��1�:�!�i��j[kV���0G�ӐEϾ�z�n=��S}M�;����{�d�nWpI�m���)���i�� ���7�\h���=ШQ:b�8ش�B�d���K�Ma͂�	Ī��Jg�"?7�("@������!8��5(��˾�]��w�K�~q���f�2�$����+5��k�2���HN��xda4l%�����̭<������UΖX���b�f�����Q����]���`#5*���r��u�A�!��Οe�,x�tj]l�}�Eh"��{�Y�e�����,M^2�[�#bX3:|��GFh��FF�t$�~�r�c"�U�<2u])��X�� g�`z��J �x!�����L EǥaD'x��g���T�F�&!��LV<L���
�:����$�sE!}�fJ��/{��tʈW�oX�60a�����W���t�v�ƫ{#k�G9�$��Ώ�l
pO3Nј��Q��L��o�R�'f�9 M��|n�����y�V憁u��K�L�=+����9<�>���Yj-��A#,��n��F���[!Ӈ��L&}�H#]AW�A�>�d������8,� �yX�@���]l�jGH6�?r%�rA�^iX�]Š����˖��Kc����mD���0Og�`���_��D�]�H��"K}������|��o@�q=�d�!#8��f�"*x_L��ZLG�_8iE�5ۆ�U��h�+���e���{>��MD���%�T�0'��H:��"��+���w�[=���	T;�k0�o�����"*�U���X[���n5��k��	���8��L���5��2�4��%p`��d'v@�5��-A_m1#�,+1� 
��D�h����.�ϳu�j���a�ʎܬV�W��/��a�6O����@°'^���T�����U>��o'�DF�gЙC��U�����/ ��W���}{�N%�iU=�`����&�9�],���~޸*�f�WE�1������9��I�����t\b:�W=ä�X������!3�#߫Nly������e��I�B�KG��pE������zB�C����>?�=��k	ӆ	��4�V���-��47p���/�M@�PSjy��o�syOv�b���� |��8���67��,�~�lKQ�����\��7�7rh�i/��
t����g��b�Ѕ��R��씁�y��E��ǔ��Qה)��!iϲ�=�>�aͫ1w̳�Q��2�wy1B|4)�Ê-keƥ����aLEǑ�u-���TvQ��/�F/T�,,��կl��p]�	*�K�	�&*���'��d��:����IKE��@�6/��4�˻�w9H��+�O�sH�9�\�]�G��o��tf�x2��jH��N���o��I[�:G,���^pj�`��u�ԫ$��еY8Ĉ�?��h���pؒ`cGԱ������t��'�C	!ǰ�`Q��'u�S�B}_��Wzh� rd,#g��zY�.��M�Gć^��?!���(<��נ��
U�$	���|�x�<p�~�*�9��N�����D�$��?��8�oQy�U�aMz���Q��,B�Q%��+��!�E� �,�j�kD*O�1��-��r�9@É�q���l�b�t	�\��S�`���]���Cn�'�,��$�L�e�g�S�3zX������Y]�{ ��J�=f���{�/�����Ns��۳z��_'>pެl�JP�iƞ�z��z���S�&s������8m���n&)�|y[-�O~��熤�����<�P�/�*?�)}��� А`~S�I�]�z�Մ�x!�3�E�FY+�Xd���R �~�&脙�)�fF�w�'���3w�K�Ye4ʠԏ�Ң�cs�����d{R�#Ey��������V"x{J�w�P)�����2K�;|U�[��ñ�YQV����a�V�پ+Pu%F�Ͱ�,�<�D0k�+!Gx����s�j�s���s[h[��F� ��V�ؚo�v���׋���fGz��Ry4��3�en��\��X�ES=�^E���^T��� o��ǯ�� �ǆX�2�ǒੑ_G�֧x{�z�����?D~uc;�6@��P�[��3K� Ρ4�I�H(�\��OD.O,doU�Q'.���ڒ۲�Ȑ"ޯ�ΜnJL�L�.N��:'��a����c�����Pw�d'&� ���˺� �b��u>:fT�k�-�E��L�B��<-ʞ�b,Y��Ӻ�en-Q�������#h_U/�*ՔǇJE��gs<p�²�3y3�tx����<�2�������3�(S�(�A!�`�L���c�g�%��`~�<�����Jaۊ}{���� )�Sg��r�)	��.hӏu�\��6a�-��/��k�vZ�XK:������ ?�_��ˢzM,Qq��L#�WF(b�K�� �7]���&$������CK���9E���ct*QO�T�����z�|��Ũ��
��Ȍ��v�����Eq(�Qڵp��AHP�ӎ�>�?n�û珋��W'Cr�J�ʽ*�秭�t�,��8FZZ�>Zn-[Va?���8��c�V�6%�|�o��Я4"�k��s���/�ղ����.a��g��G��0w�!/���5�ëO�Ƣ��yBl ��p��Ud�-�5���r4vl��������V��䩂�}���f�j���+��̸y�Y�{�0{=���L��`�4¥���̀���xcP�C���9��r"\���H�5��6V��h ��*�[��;s�5��˰B;� u���o&�&I	�p0e��1E�1��Eʗ�<�ǐ65�4�ѕ�¼'��_��8.DUׅ^�`^��P��&K>�xa;��^5t�e�`�V�=�eP�z���2od���.K9 �F��W�sE���v�Rg����mGˤ-�A/Tf�J�GP�D�y٬�t��9F�u�tec' LD����!���RB���%���c�4���s��נд��`>W�N����Ӗ�o����mMtx�@�V\=3.�|�aU   J?wDE��?qE���=�����pՔ��"`)xm�`�&�NGs��/y��M��1�����&E�àL,y��^ɮ�1�'�l����,/��d! ['�@�k�928���DFl��E=?�Q�T;8���L.�iЭ!�,\�.����%�����c�C��x_���<5��|\�"�1�2&4{Ѿ^�5�CP��}�}����؃�����剚Y5�t�9��O��G�Ҿ��8�~����(��:([�l�z�������_�  EQ$a�!N�R��8hx�Ҩ�?n��t�ɠDmFHsf������M�L�a1IB�4��L�[�\���#��[�e��c��ܕ�m������!�"�h�G��r�%�$TL��:鱡�d�9�S�n\Qg�+��OGv">��ף��h: �Fm{�����'Pʮ ��7q��- �$~��B��#���9ߪ���%=�l�{X7���3ԮI��j�&P��g��}o�C�9+!S�^q���-�`�&ad{�_ʦMϦ�k	p�����
�����\
Ǚ������e��-,�>bm�d���P)÷�QX��]J �<���ȱ�F�7a����>��$|�b+N?��� B�`���8ۀ-�/ڙ��0(c��ڼ��5�R\��';|6u�l�}}�9N%��*�����
.X�q�K��XZ$�A^)J
-�=��.��u�uc���:%��6�ј.\(��ֻJ2%F�0� ����q�@�qv�l��~x��-��dqى1&���bG�v ��a�2(m��r�/aVԹ�醌bc����{O�p�
��i��*v�RVn�d���2˻1�Q2��� j�at��T7���,f��*ݾ(a��U�3S`�����(;�����X���K9����x�#�^�2�sB�~�DV�� E�)Ҵ>������$'Dw�����x}w����Ez}��bG[T��+�M�>: ��	���.AQ�,����ձ܀�?�t��c�a���GyĦ'c��߁Y�O�Q�(����є��8sc���_U����g����yM��R�� ���jS1���A�@������A?s�ؚW�^ז�|�Uq�G��Xl��x���ތ4!�h=�k}>�O��&d)����F�,�[RU��&z�����:�U�d��Û�H����\��$�9��Xt0=� ���t��mM.T2󮇚�U̐�����K��*:Pj��r^�B<�?�T.����:�xl�-�p�Di ��f��c��e�1"	i����p���j�7x�Z ��c)!Njr��ţ��\���E�+(�IKG>��y�d����@vп3I����#~+��Mn�v��b[��x�Ҹ��w����U������@➝�Bq�6WM���7iIC<���D��(k���m����?V6J'T�诜���N{��e���c*�t�;V*���E�FC����.��U�X�ﰚV՗�7��z����J� �J>�����,���'S+QV��{���l*���׳pU��2��"�������E�@j���������K�acļ�Ji>i���E����E�������
�(\bn[��yX<�0�gI���O�L�{����^��r�lɋ��#�'���q�f^�U�M'*7t������"�)��4A���̌��ٻH
�d0�{��ݗ�_��~މ��f�3����j��W��~9�<'�?tPɖ�}�gKg�a��D%I�;K��Q<���p��
�h��(�X���:��S�f\�.�C�c?g��>�J�Y0�f�<�;�,Q��-��P�n���Z��	���l� 	�Ę[J��i܈��~�y��?�a^F[5�y ���8�ry�������kM؆�	�8�(�pHAWTx�qM��l'�a Q�}+>|^�K?�*����E��m�9Ԑ�<��S��сUR+u�j�6��v��r}�����l�q��"ߥ�����g^���w�*��ŬHZ�JQH�D�1֯ �'���Aq�N������h��y���"��&MH�n���.�.�^$Y/���>��c���b1?IÿCT�q���[��GRٟi�T�'�����d]#��ȴf�I�R�'�v�#�c�V��,��3�7#%��eK�
���"�_�f�����q<8����Z�N�g�C��vZ#&���5a�Р'H���4,���{�Bg������L�`�O�E���5&c�k���� ����,+o�v���T�'�˥u��F�b��I�;�h�a�%�"���r�\za>CG������*�
�z�݃3e?����	N��G��ʱ��jpj���e��j�:�V_�e�����G�.��T��͉�e_=��`�]$
6{�~�̪�� P�"b')�`����ɩ�f"�T��k��&��������=Lt9g2��E:e�q]ZL��36�{��O�Go�b	j61C�p4U'3$%�Z��Zp����`0�s�S�B5����rYR�֜o���J:���_#T�Wg�c��X��%D�lZ�"�� �*��G�������%�"�y9-���վg�~���|W1E�w,��c9Ϻ��H�j:��퐁���i���]xR '�s�:��Ƒ�"��ѥ?�|�\>���w󾻼�d4U$�4��b����i����Z�K��q��s3�3u�Dˉ�ލ(��FE�g:�6B$rc�2bMB=�iE���]��m~M#G��F ��R2�ÜV1��h�5u[�Qd<��cf'&</j.�@���wQ=��^*�r��S6��f=(���HD�u!a�%@��Q�2��Ak������7:۱�N�q��p$$j�`k-��b�����ԍɬ���`�k��Z�.���2����_>PC�3�xr���j�y�ǚ�x-3�иf��k�?��Y��5��sg��T��6��l����X�}�ٲ���-���?���������&k���˞��l�t���1�Yn�5;s�Ɣr>���j{�ᵞ��)ȉo�[�7AW����0:yr :�=�ٖ��No�~�I��u�p7Zq�5܉�6�Ծ|���0�1�����D�����bY�:10F��@�l��3ݷr_jx���G����d�z橘�H ��#���%Kɱ#�"���[�}3��|Tc�����΀3���m<^m���ز­�G�=#������k�!�m9�z_����>�22	;���ð��6Dr4����j��I��9T�N���P����z���rm�(�Y�z�f��I�'VY�ڢ\aB�H�H9���n�;K��	gS#mPx� �WXϰq����O���[�m�'�=�0�# l��ٌ挬�vR3�
C����oh�Xi�������N�Fo�g�|0�7s�� &T�8��q}�,��}��;W"���lQ�john�#�Dm��\�[hF�i��VV�|�D?��xݚV5�~��\� � &�՝�"��Wj .�"P�9��e^~dJz��\������P�a��,��F��I�U�Aa�<�o�on�F-@���钝����*`]�"��kD	l���`N����[��OcG�{�M.R�~MI4I�#x�qz�f������k��l F8�8��KgC�f.wn�oc6x�:\��QA��SK�Z���L����|]Q2�)b���϶�&`�3�ʬ�t/# �,��v�G?)�y[�q{�F�l�l����b�P�Cvj��P�R2��t�����lQ{���T39.��Nl�%�A4�WQ�ݰ��gY�m��%���~j+:}����m��F����u�������+gY1�̣8��V��98b@�1(���	�^}�9��-BPዄ��P��Z:������6'^Nq�F"��4�;Ś�ڼ���ߋD8���������C�^�ł���ܨ��y��� �TtO�4 S���Y��О����0�l�l�[�n-�H�Z�D	
�̨����4�