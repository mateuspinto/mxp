XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����$�1�����:��z��ثM���)��v͉����	�.�wH��i5���ם���	�Õ�d����-X/�����H�̠��@��m9���w���CZ�nKl��|r�u�����=V1�K�P���ހTi]<�����&{ه��yJ��A	_����z���@���3h�����ne�:��հ+�+��� p	��(+~�n/x�6o��e�҉�y }D�'�#�<-�����ރ.֎���@�p��e�-<�<9$Ytt����`�v򡗈��K�����~z�WO>q-!6���ٮ��f`�����e�8���X�?R��Kofs��@�mY��m�Ӹ�O�K����|�%��1��WI�7J��.��r׌�&�'[���Ҁ��gb�u���,�j�"�Od�+��*���#���}K�7<]F�����efr��O�)��\6y"�\������T��>�T�b��ᚧ���owQ̶>x����?��n�7�B�u��P�P�}=�o�R�$Ch�,K.* f0�j���a��>�_�u+Ǡ��r��Yˋ-�9�$P��@\�V|B�b��C�v�nc������ă�^+P�GI�3�?JNwr��4�cA��z3��'��Q�2�o�7���5�"J�`DG�����o�2�M^J�^�rˠ�e{����jx�k�!`�u� ����kU���<m�b]��\�I��3D�I�����&c�V�������AuMYE+���XlxVHYEB     400     1906�]9Mw*����A��,&{�"L���8x�Dzb��z�I �H6��^�!��<G� ;�����?ڷں���&����Z�S~p�r���� �Ǒz'+�-�ć� ��Q�!_ֆ��`D��(�Z�"�8�pwX��}�b����$�q������"��N�^IW`s�|M�zdF]j�6�=Ի�hf8߬������b��-+ �ᄯ���Z�T��ojw��e�P���"=��ޯ��_�}��.HZ�(�cʉ���n�C<t��[�ٽX��B4���7�Z����Vd������d�rb�6|'~���)�t��~��ѫ�}�P�6��d� ᴣ��fE����WXYIL�9u+o`�}�� 4I��j̚� 3'���� ېXlxVHYEB     400      b0�s�O�n������g28��m��F���C�� ���u�_Ű�R��KJ�����������������U�ʰ����7�so��h��M��A5d}���/�^��<y7�0�f�N�pr-&2g�Բh|%..����x>���ޫ�`�#�u8q�,M7���O=XlxVHYEB     400      f0�K�t51՗u�.0����P�����3�S$���w{�{⢤��}�Wsj��-]�%�a^{�6]	{�e��58ݭ��x�=�M5h��_�9���`��mu�{�99�XI���F)N4�Xu�n��3 ،5x*��3��<+��(.F��jK~����./a��͵�:nJ�6���ܾR�����w�_�/6a�鍩N�ְ2���>��1���;z�����o +��� �j�U\N)�Z��XlxVHYEB     400     150l�#-�r�׎�v�
� ���3�vl��umwJp��)��Ά!I�&� �V�]V9꟩8��X�P�D���o]2�)fK��71���-��crd���|�8��^��4a��L�D�XV��X�����EK\�ٱxj:W� �u����Ldh� �ν��ꦅ�
fYi�7:�2-���}yi�\��=���ƻyS�e%�	][�0�m������w*8q�;�wF�6%��)nu|g�ib�+6��A�-��̪~�P<�UZW��ܢQ��@��<��X�V�]�T���@4xn=�>J�}�`�-5��s��i�G̒���O6�(�aY��Ϲ�XlxVHYEB     400     160�Z�">r}�����B伈T��?��,��2%�Ā��c�c�0p���o1as���`�
M남R3����߂�8�=�N��I�I��#YUl'~L.��� ~��#|]�o��p��&>wz<}߂z�ʞ�x*,�7�֔�l����ߘ�,ƌc�����f:�&�|i��s��Ta����6�wT��yL�UKȰB�)��ok��@g$]˦C��T�S#�����i(O`f����l|����kԆ?<f���O)TsI;����ʩ�#=��)6E��H�t�P�`��
�36�NX 4/��:ٜ��8�w��R�+A�� �����R���ѡ�$m1�%����]��j4�XlxVHYEB     400     120�$y,o�0�(�uV{дBAd���!��߁CV�e����/��F�q�,���'߽�F
{[�c��n���-U!�G�1b#ߨ��ch�.z�V��X�.��*f�9��RТ3���/=B�����y�?��6��F�fi����~�RΊ?����>��;WH��Wa[L��̓06�9�Q/�OC�<gR��;��p2T��`�hv��gf
f:�D �w�/pO�����	*���5k�H�G>�6��ة<���$��6�Ɨr����v4,R!V��$am�.^��خ�oXlxVHYEB     400     110W��<�~]m�f�l�[�ٞQ���M��l��4�L�`�rz���R��\��!%U(]BiˉuBhΏ��(yj_�>@	KF]°�WqÜ��Ã�h:iG3�N�;8q�oх���?@t�W����%�{��/|n>��Ջ1wYԇg>���C�5��F��_��(����ڒ�#�������|04�"=���.kϣ^�j9�	䦁ʤ3��nVq�$!.ǰ9Hǣ�3���"^�������}��ǲ��,�	�u�̄mA��)�`�lU�XlxVHYEB     400     110w�C�/�H���\����M3� �S= r1��@�>��;��̙��Qu�Jtͷ'8��f�[Lu޸�x�����o��e��TC9Ŵ�eG�P��s�w+X&�jF,�����'���k��
�c�Х쐊Z���0i1�t�Q��x��óP�$N���px<&l��#�=j�t����۸\9md�pM��ot�9~�5�u�yS�a)Q�c㙚�f	���K5��]d*M�V��g|�~���F����3�I+��:��*�XlxVHYEB     400     130�.�笵8��J2Y8�9�E�on�$�w�l]1�{<��i�`��O}a���z]��s�-;/ �g.�������2lcJį`���{R'g��_"�o/��y���x�P�EF�ұ<�69��]|(�i��Zr����2($��ߓ�^m���:�Rj9�ԤQx�ng��?-�yQ����V&���`�>��\av���Bu���`�#�&��&T��h?c�Q2M���%�	��[�L͵R|K\y�m����R@b��C�&�����]�J2e�6
H_���4���8	vb���&�Q���XlxVHYEB     400     140����%�mPf��@bI{�3EPY�Nݹ\�[?�����S�ļ�m�s����Z����<ظ~���� �V(��<юh��-}�4���ۨ�H�����B-ضd*���a�	P��p6$���*p�����uwvF샜��@��w���������Ώ*�ÝW����_(-ɭ�k�F8�T(`9�̖�I�ʑ�D�����5��/lJ�@������g?��l8Bn�H6��T�����%�VK���zH�����#�T^J5���fT� C5y?:z�'�$?4Fߝ���{�a0Ҷg�[�T�diܪ�KH�c�=ēXlxVHYEB     400     100Qf��tN�a��z��؁�u 'az?��*����B\>Ts�?1Q�K
�U/� ^x��ɰY�R�7��%X:�z��?:R�:k�9��'�w%�����Bb�GO�DN�n�L��]Ag�(8�TaTz�&�nZ|�("|���`_����o�HsZ!�6��B����h$�P��!mY�ۻ��a�1ܫ�^�g�o����e%?X�qw�x)�L�K�H2�~\��b��x�i.
�V��$��0�jtl=�̉/vb��X&�XlxVHYEB     37b     140�H�>z����S�/����rd�KI��m\e�y紇�hB6!i�;k8��\�$�������G���� E^yC>�g�a9�[����݅q��Z��W�RӉ�%�;�z��W�#�Yh�J��>$hL��P�'R|T�M;i��gE���!�[F����x����_�5O*��K� ���8��C�]�/�^l��ʖ,<&�V������.����1-z$D�:^�sý� yF�ت 3�V�r�m���T���v��ZT���s({���fY� ޲�Y$�"���y�d1�@�n��q~��K�5O;7ޱ��@��*��q�