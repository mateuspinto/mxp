XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��^��;d��ô��l�� ��\#NAn��3�n2��`#�kz�J5�a���v\fѧ^'��"2��OVL�B��6����c�]=C���&"��.6���K�~�!Um���sv�����P�<x�)�GUR���d�L����M>9ѐ[͋�dH,�;>Y�!ҳ�)#�_�YW��5u��3�i��SC��m��u���ɔO3H�Δ�3pA
2� �^u[f۶�we��H�$U�OLp� ��;���q5��Ł��� �i9�K�Iyt5��5�5
T4Dw%���/����u��6����7-B��̈����l� N��DO�-#��,����~�$�|�[�ξ��ٻ�EM���jAv�R�XX\�Ǘ�;?z�6K3'��n�U���3�O_��ӂ�1�R%�Ʈ1��i����>
j;���2����V���ha}�����vِuw�"QmV��L��0�K�)� ��dW�Na˸u�}-�;�b!�u��� ?��ieڠl�7�uS��)sQ��B�+eڻ0�x�6�W���>D�Pċ{��yrKq!��.z��Ư���Tu3]���!�E����-�����[�$/;L��<V�	vR��6%�t�O0�9eM�t��h��\)��z�Ֆ��eu�pv08��Fl,r�'$ԓ��5F�>�*�s26�И{�̐z�:��MC��0Ct��H�y��(2W���5��`H��j�:M*B �g�z��E�9��I��O���RN�SHNi$栞e#���XlxVHYEB     400     1c0P)��sy�$��,W�Mތ�)�Z�=L�2����<U����k�aD�wd�ص�i��i�݄	��>jg79h�� ��\��T-��QCǲՕ�t��'�a�םfD�'�'F�+�%ZLκ�;!�l�ΧO�����쑊Lp}B�w� �f O���t�T��1'���EX���3�N�������]Q���ל�&/�����wd���֑��;����笒��n<�?b�#�5�C,|�?D�*����ED	���o���+�R;pl=�㦌�uGWKЇC�Τ�:O+���:8��LLhb��C�Ԇ�Y쪩����u��PN\��Ӄ��7�d��Q��ܰ��͹t��!��a��[a]���XH�6d�8����K�����pǤ����H��M���n41r��XQo���HW���?U���P��;iZ��T�5��#YXlxVHYEB     400     160��a��w٦���0����yCM	=�)&@��V�Ќ��YPߤ���V��iw�h2G�؞�mȋ:���(�SP�gj� #����������5��"9!�ؕB���������7��w�ӹ����ͷ�fyCr16��3Q�	vuޯ�#`Xə�70��Z6�eRB�n3�e�w��)�s�Z�
��XMJɹ�,�O���+��3��$O�[�\��cn�_�cs4��l�.�,G�jO% vhu%Ai�H�fHQ�b�M_�
��Qo����:M�L�v��Ɏ���	�l�y��l�fԇi`fbg�X����z�D�3�<����Ɵ��i����ڙ�
3b��2XlxVHYEB     400     160y]�e)LN;�W2?G!9�$�+��6꽷�������R��YЖpdmZ����'�(ݹq9��G�?��7�W�#�C��9��,L��M{ԁ(C5��.'�q��Zu彜]�X����{�^S�X7S߷iY\�o2��O�Q �+
E�� �����ՠTu'�.���Khx�v혴u��mt;Z"EǓ1̨g�lN����&/��R��	����2��)����3�R�tmƁj��K��lu ˑ
���������n��VD��hM�����To��0���slT��"�c�V����R�$x"C�8!;,�&?2�^�XY��GnHl� ��"���W�|X.�[XlxVHYEB     400     100G"��Ǖ����Z���[�R=oɬ�z��4��_WFQ%�;��'��|o#X��N�4�Z-���X����0䓐,7�������C�F8�64,���js.��q�Q#�]�����������{��1�}AH��-��Nߑ�kY>��G,X�9����b��u�)A����Q����t��S��OOS��*� =��X����CQ!�������l)&}@>IT p̵���U�����eF������~�&�P��XlxVHYEB     400     1a0g�]B-�/�J4=����/�y�&�9C.����wѽ�{��7�.Co� ���S�!6�����Щ$�Z�uwV��hf!�(�l��	 �� G��F�/�	<��"?o���.ĺR�DبDe-�@#�c*��U��� ˟����U�T+�����>�|�e�7n�E�~�K�r|2���(�����?�t	�y⣾��p�z������QL~b)H�B�T�VE�1�}l>m�_�q״�6�s��*�ia���8��
�P$�>�šRD-�*fyě��NRN�d�Q��ɠ��C��3�a�T�t��dV��˻wl6
�d�F=�k�=Hr�q�v�"Ąw� e)
�G��ɖ}�]�:8!�?XusD�d�����.�O��~�V�Y�I �H���W
�b^�2`XlxVHYEB     400     140��Y���~�9[#g�5���ʎ�`tWKB6[�@q�Y�s��Y��"�aݬ�
	!�	V�*��E�"
=�ẠU�_K��-�0�2,|�'�@���}�������.��W�/+:���M$�ݓ�L�({�$+�T��[i;e*��F�6\�.ߍ����Y�<~�E���T;����.����/ئȇ!�pdI�qI�m�%�e�a��2����><��Sڵ_ �ZIPv��>��z�5�\�����0�;�C�`i�N�� �c��h��
�z����",�	� )�����V�݋G��ͻNO��V��]$�4h���P�M�]XlxVHYEB     400     120��R}���9���=�C�ׯ��r��q�LC��e:��y~:�����>���MJ�\�[�bU���@Z��v*��v2T�Z����ꐴU$�(���U�W�'ƅr�x��
3#C��pڛ��{e#�f�Ƅ���|E��"x��#F��.@�/>'�����n|3��G��T<�h���՟@V�$reX�6e}��'��N�M@MIoU�������{$��������N����`�߅4+p�<Ma����·{8J���+	a��34�ae孄{���XlxVHYEB     400     130�F�'.ל�Ġp�>WU���Cfߎ::��]��`�6����1��1�@}40D��<z�6������a�/@��?e�6�5?�8%E�޾��8�q��G��G럖����§���/���*��r�`P���/?���\�w�=�taENi�����!��*�����W:�'���+yK�a�����)���lơ_��[���{`�{}�Z����U�:HB2���S���2*\��A� � 
�p�#�;ȩ�IWkl�v.�b�2%�yҫ�Ҕ��+ ��#��As/��:?�Ǉ�
D�ϜCAH�XԔXlxVHYEB     400     1c0Y(gW���2Q�J����싲Q,l2�d0�m�N}��Ef�A�ļ�n��w�p.n`i�1���ֿ���#V�X���0�����<U�=%���j�
�����?W����4~���ԧ=(�j㟚ϣh.,#�F�I��#�#����[��-�?��H��[���t3t+���;�����C#�o�o@�ꝟ�f���X���31(�F�P�?�&c��$�H�L���v�Я���'�--�Y����?�]9�.J��wDz9L4Kw���F���|�K�;s�;��&#���|	��ħg,0k�v���>۵���:���oi��L�v+�Od!\Y����iU��j�N�'�s/HqO�wjw�T�"�ݧ�&���Hy1:�2n�
��R�x9q�ad-�!W�7@��mҚ�L�&����E+�s��g�.��I�gY
�>��WzķXlxVHYEB     400     1a0׫��w�~lm��t_�������o#��MœR�<�N��|�	F8G�G2V�@t�Id�.q�����4�>M����}E�~��.MO��������2{4�f��	R���x�"�(u��"��'@)�/RF�
'	\ZF=$E�:r�D�=4�Ķ���n+hN��������:��+C����?���b(2�?�c�a��i2���]�q�l̞�^h����|���\~�֭���jL�vAv5��!n�}�X��z��ɲPչ����L�8]�;�r���3��E{Ub��]��ϛ��@�et׺<��(ɼ=zb"d�Z���G �9ȞWK�C ����W������`'h��Ȫ�q(���o�� u�Q�����IP �/�:!Z��G�1�}��_%3s��ՠ��Δ$	�k)sY�XlxVHYEB     400     1a0Y"�Y�ކֹ��ס��k���D�S/&���}�P���é�Q_jH0Y���Qv�*�����q�ӯHkm6���4iVOW��O�/$u���ӡ� �:i�^ݬ|#S�&��R~Z�T�]���P���� \RH"��rH���C�q*16z��/c�CvTBܩs9(���/���<҆�@�T�n�" �T��q-z�$	޿��g}��݌���*�w�3ix�\�jiC��Tb�P� ؚ(%�����O�i{�"aa����ɦ &��.��XzNw%
��dnϭ�i�Y�_����)7���E-YF�jU$s�S�+�xg�&u���?�̟,[�*Zz�;���]� �H�Y>����8)O+ Y�܌���hAD��%��Mʕ\?�k䵦��;>��Vo�zb�EB����.vXlxVHYEB     2d9      e0��/�����oE�����C�Y�S[�E٣nz�3���@�-�����q7��6@��w��ƌ�b_巭��Eni���{`g�y�����p$g��S[U�B��ɏ�SEA��`�ڲG��~߃R�AD�O  Ү��G��p.�;��ƕb��5U���c٭�җ�Ǘ�wx��>۟�W��8�7��\^�P�mgec�K6c�T�.�ՋG�q���Yh���