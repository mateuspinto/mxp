XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��No/q�/}��]�ᕚdÜͬ�h��Ψ��q|��C~j�X�˯m9�� ���-����6��FPX����.��fb1dƘF��vөs�\j�)q�0�ȃD�W�`�&��p0X��K!.�H���^4k�>�ѻ�)�U.#A��0�h�&P�X|�q��x����Xd�Rd��م+Y�G䣀��8I��\�W��� t(XR�&ri�{�1@eyM��2�t���:�-aOb:�%v��_d�������R�f����Ѝ�$��Œ̿�c��B��%�=%�0,av1~,.���s���i/��{}um{�zˣ<�F��Q��2w��m���N*�u�Ш�z�!��ʃ�2�s����ޚ:ŮW3>%��:J��n��F�����"�7���<^=��(���x7��ox�LGԠK�*��Ĝ��ˢ8��h7������k%����y �\GLJ����a�_��]=��#(f��H�HW�q�ά�2�+��6�: t�3�����j0\-���Q�yG~9&J�0�6x��p�I��f�N�PAt�&B R�n��5���~#^h��Z#���wǤ���<v���{��CF�M��i�N_j��Be�Ei�Or`Ѣ��n�{N��<E�ッ}��aL��:�������W� �Q����5����R&�N�O��q3�Q��>��E�/�̡?j�"�Z�m�`ٟ,?\k���ZFM{9�41/`�'�T�G�[ڑ��6�"��`���f���թД���XlxVHYEB     400     1d0�ƪ�;9oC�6��٭�Q��Νr��k��s�E]�J;:�����	��g�w|�����u5N«�,nUkg;�Y'5�B�P��KX�$E��.x�z
��l}s�C6܃4�K��t*Z�	�k�����3�xs�����n�@�x��9����)ݘ�(�+������$���=_�F�E6%�98ЕjW���xa�t�F!pkIU�C�n� ���I�W���?���샆����#��3U�ak�g�ظ ?�-`=g��K��n�e��� \j$Q|A#�J����$����iy,��
�r�s`���6�� J�*��P*X�'M@ԎD���mhQ�����Vl\��,,x����	�?.-�o�=�IA� I���V��~v� �Yq�O�}�U�O5�M�(��y����!\,4C����W�A�nR8<*3M!�e!'�Y�ŗ��'�T�?��X˦XlxVHYEB     400     170v^��������5o�(/���XI@�_q�k �)>!܃T,��D�c�$s���^�(��&�;Ƕ��+r�$��8Xf5��y�:Ecj7A
��w`߷}�<�Ԯ5b��ٗ�X���y��^'�I�X��D��N��A��h�}%Rؑ%���ۧ�b���xk�/v'��H�hK�V�����N�!]�8�;+8�G��{x�6�T<��Cӱj��S�T�����Y�&��RbtP BZ��VZl3�����K;�ﾁi>=��p�8�4ri]b��uLyq-g�H�(RT؏3�5:��3Bb#�Bv's��oԩ���1�����]�|	R|x�TƬ��ſ�
_l�G����,��u���t�nuX�dXXlxVHYEB     400     120.�Me����|w�.q�4��,e�~S���*���"yV[�߇!i ��OE��gX՟�s��C8��/�b���_\
ϫ��30��%D�T���TA���4򑂤N�/�Y��,�� �*��zا���Ó%���/��S~�e���5p�=͒��o
:Dp�O�YYυ��
�8z//������ �����C����̕Zn�
�`��	4��k."3�?�!��˹a��P8��r���$M���h���#w��Gr�Bׅ����`b�OH�Ҵ��(W6�� ��W�XlxVHYEB     400     170%n���h\L�҃�UR+2m��D��4�TK[�,SUXwX�b����{�|[����  �O� �J��ГB�+���,5��b^�jNrVÅW�b�^�(�}��G_��ȻM�b�<�"����uNU*7E� C�K]6�˾���u�H
�f�_���+��lR�=�����4WW��V)r���s�<���l{$ƢƋכe�2���:�nM߂곋a��k�.o�������P,5���X>lЅ�C�IkɬFː��K*,SѸ&]�?W8H:^Ǿ�׃Gs���8�m93l��N�?J��
��CC��]�IQi�S�����n�Y՞ٟm<n�VƧk�h �����6�eXlxVHYEB     400     170�5��8� �k}�ȡ��g!bBR���QA�T$�v�q�k	���kz��r�h��'X���* ���f��BW뗴ab��TȀ����m[�U÷M<W�Ĺ`TҐhOk���̓�hcb�wNf�� xW/Y��aL6��.�VЕ�k�^,��AA 戬K�b�E=�[��Q�������)��+K��0D44�WIY�D{Ttw��P�~N(�Ű�������?�/��z%F6�y����I���=Xt�������F�o�a��Ͳ$������q8��G��gJ���<�����L�!Y=�Q�B� �.{����c�,�{2�,��{!��e���&����l4�O����J�d�
V!f���G��)hXlxVHYEB     400     140P�mL�Wۗ]�h3Q=C�k?.��H�l:�b�?E����.7�y����©����*5�I�b ]�ۛ	�"��S� RG&�
72EY}��+�S�-+�_�~^��lA����ȝj�Ns�F�
e]g�`�5�/�~�dg����7	��OA�"�M!ޑ`�dL�U\�x ����J��ȵ-��03h�H
<������8N���5���"���+C��bW;��0)�i9Gi�bb+�&@����H�@��ƴ�5���j��B�	����:j�����6uZ+�*rN����fg�����*@L�4G���XlxVHYEB     400     100Y<�CBv��/�w��J�_�ݑªз/���/X5���|�V�N�Լ��;�������t��+mn���rgBңV;�!E��	�0��x��GL�)�r�]���]��-���Q�i?e���a�Rl���Ǉ��8�h�/�$Z�����Pܭo��{�v'ϖ�f�~o:�d���ꍀ�Rki���7�d�9�	e���E�o�X����q����Bl��h@@�M�zV*�HT��?zq�8���b�XlxVHYEB     400     170e;{���������U��$ �X�.���f(�����w�Q�/-�8�����_�G�V ���?
�{u��3�g�]���ɶ\|�{9�+l�	[t�
ʋ<���UVy�ҝu		qW�o͝[���:�d�jЫ������5�n0����������
7�"�4F�27�������x�]4��E�BGl$e+)J�������s�c �Ʊ���Z_�$]��26��jK@���Q'N��k-��@�>����{���
cT$�'��΃*8��Ӳo>{Oe��f?���T-A���A��AB|wh08��~~۰�K��Sjܰ��;�<��i�&�5�2n��@����3y��xU�sY�xXlxVHYEB     400     1b0�'��C�ڹµ�ݠJ��?ڀ��W�f���O��O�pf�Y��<7���<�H���䐫���&p
�(�T�h��~�'z�
&�	���w�LL��
�ԄG��eJ�m䌒k�0~�c
��t��������\�r������G����(G��?��~������%7�huF��QQ���i"�u_&�W�t�MgJ�_W��<���"dſ(h&c:D �P�v�
�\�$0f�7h��,�8Xh��m���ԪHA+%o/u�
.�uʮX�%�]�	zR5.��-�'hE����~w����Թ�ۨ��N��-�)�aX2�3�cj4+U�������, `���zzE��\�<���I�W�@YI��yQH�Zr$Q��Pg�7~0F���C7�ٜc®���<�RJM�����?�j	9�sE��P!XlxVHYEB     400     160rw��,���(��o�Kt�M��jO�H�5���c_��|���}@���������t�r[0�<�����vK;?�u�X:Y���)���sGeo�O�MrDq:ɀ��T�zb��8^�X ��_�ز���1��J��]v2B�0���3I���D���J�͙<�/�꛸��� 4�&�1��d�=�@H+N���5����/�ꍦ��tR��R�QEZ�K�`��b@��̊�q�J)2�,����Ts3_U)��%��!L�x�M�>����+h׻	!�����n�};�[�~odK�׎�H�� ���¨Ĝ/�ऱ���ڴ���:l�&�j��XlxVHYEB     400     1d0�;���a�[�x5�X��w.���v�r�{����.��\f�E�w���h
r�jL��\�Kà���`r��jK�u�-0�$���o��'�+�<�V�T��P���|�X��>,�#cY��G��ê&�ݴE���JN�:v_�:��d�^��|ƀ1�2�ؐ�`{Cyj4�3V�3�u�aY.j 3�>�*�F��|Z������$-��-�}[%� s�p����1PiC�4w�lA�97�O������+x�C)��!�A��ǐ�E���}R�I���Fb��9O}%<Q�}#w^� Y��ؠn�yo/�����ͪ�WL	i7s�C���g_�.�ͅ-��ë47������a����a�&(���$42Fg���
s��V�uIل���h)u�Xo�/����5�|�D��x�"A!Kv1
��L��X*E��c G���-o��ξգ��XlxVHYEB     400     170\�ѷ�6	���9���/�t�^U�IEzI��L���$�`��q�G�}z<R;ʝD��+�����%]���}A(ϏB!u�fO-$��L���\�Q�|���4��B4��Y�U!�c8�E$h�qkE��י�8��,��$��Sp�WX#{������}IT/����Ǥ�
�9��*��*{�l<Ø?��+Y}		0Keɞ��FAo,;��f��������7��*y����L�qI�1u���ְP֨�Y��o�3y�N8H�=� ���k8/���9&��
�e�dn���w1ϕ���!��/.�xA�:D��m��<D����`���I�ê57]V"s�X�P����!�S7fY#P��XlxVHYEB     400     160����F�>\�y�l;�ϕ������M36|Ɍ����<¦�;d(� cpT�O�(SI���+q�.��:j��`��pGyǝc�$��R�o�\r|�r��ַ<�£�[L{�EĬ�\b, qV�Ķ��gT�|������-%M���)ЙVa�}nO��e����æ�=���FH���S*�Q���U�»�)��w��4Lu\�C_>��h��������GؓJ���W�2~E���3�R�z풳�쇰�Q��KG
7��2��	��8�j����t�*�����k��9����Mx/�)Q;����M�,�ȍ��1B�� %�v~!��x��q�D��q�C�XlxVHYEB     400     180������:$�(��)B"�@��q��6�9An����8��8ibƊEr���~;=�@�b|�1	�,�؍�QIa�o�02#�ҙ��砧��P@#ډ�dm�f]��N���/�;u�ŗ����|��:_�X��W#>��V�	��|h ��a<���I�����~�l�p�>p��"+)�-J+�=~~/���$���t�����h}��-�h�����c65���p�Xw����W�NKi�m��M�?=c�����[.�M�HzqA���pvh2d}m.��6�q��A�:�9�>Q��C�dC���N�?/��:�c~�����c�����@��K���EP��o	��%N墛���c�"ip">E�����XlxVHYEB     400     130�*��7�d]��Pܟ��(98/ ]���V�x8O�H�|n[��In��XLZ�
�š	���@����p*
7q��T�ۧ،!j
m5���A�z1���-)$��p�T�~�u�����Z�{v�
�>7(��|�C1%��G��0m��v�$[�r�m�-n��  ��p�m���<��"Il�e������s�.R�ЕS֥OӲ��^�Q&^���w/�ؕ��OJ��&̇%1��0�����0En7'�h���� J�94B�Mp �o8e�n�Y4��� P̥6b"�RRw`º|5
I�r����XlxVHYEB     400     160�>7p��|R��cʌ��"?��E�e�S��X# ��Vv��V5���[�&T���+�|T��I�b�%5���zt�y�m��e^�s�3J���FW�i�5͵����"��ɵ~b�̚a��S��@���������+��?�ټ<��x`���V��#����AW`�MI�?�3r��U�	��$��Й��7���p��/���|*�L�,M�U���Xb)v���;d��VxF���Sف�Q����mWD3��LY:$��\^�b����mt�"I���
�7ov���r
����p�Se�:S�W�����#�-R������.��Sg\H��Gc��Yz�f���XlxVHYEB     287     130�N�a�0�l&p���M�IQ���3JbȜ�8l�,�凯�.(>�pAs��0>��&Q�U�����a��Jk�	�{�^>ߓ4�!8֍R�D*�
P���=�BTlka����[�B����Q�������Q\��a0�u�C�� �o�5���>�o+�Чt?��YK�nM8�^�8߫@�<��iH���ϩ�H���1���!g��Y�TyGF��$E��#:�qױ�3�z�C�+�[��t�B /!�:��?d]�Z�w��&?, ��6����C�t=�6���_���(�Yq*��