`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12016)
`protect data_block
PurehZ63j7SWdg61YbW+tRhaNP8GcRJGoYfLpyvljAId9FDnO1tJjtfIdr+IdVHQEHzBGSgq6GpU
b4Qk217E8OPPRgg/wNoCNmAg7Nt5m/DktsMAKx+UzB4P12VsyJZGZHKGwthTyriG9T+j+4KqBWhK
9XgFaQYcfSGZ4YczyJSpixaoml54jDQtrNWeGfEUNEFPeKEx5rrKGqH2k32z72kNrB6msGfuZhw4
dUm3T4pvs0/e8nhG7Z9vjxhHQ8tQBwyvI7/dX8seVC+KbDK+b2wEvgrenzmhKDAGTvD3sLtMYmeP
wTU3F3Hiu8S1Vm2ch44bqomKkHWlcWPNJOkY223Qt5d3KRfjHNCgBcDSYvLrbLuLtrUvvR2TFN+5
oby+ymFnN5/y7kW1o/qxmVec/qYuJG0Tg0EtHgDgCbPmU1EPY3n6XmjlMI+QYxJYMzOrWljRHH9R
j/E/lfVRqDXPI1Ng7dS4ZbvR85DwsedhsI4MkJIw3dHlTD1eBrnprotRaT0VIDQC7WIrSVeoOVqs
YmAzsFBlaikHyjEnk8eKZ9o8SlgYniJve1Ifquj/spDLaxa6S4/9ctF15B8CZM1XGb5mrqAR76wH
4ztaB/kCcn9UZsD0GA9vwp3VlHMgMSA3og3GhoNXpo8yYzgY5mHPpAHBXN+OQMRcvlz0GV54b1p3
39DThxLOGxN4gqWbnMslQ+s2e+EP/XZW6+Q1Ss2HUwiI1SIBYse+e7FjZ72QMJnWWYzdaZZiWPIw
zuR60uK2hcjFqaU2M/SzdUxN1YTfXFVOSyyYpQEx7Gy1FxN+mhLDj0fLvAzBUhcfRB9np2pKSMw3
p49MZqsV0lMWs3XeUWCMM0G+zxTJgnE3J0wPv1GsG4SQrChhKu/KrY5WRO3VKfcnmWxO+X8IABs/
iTSdyrlVrcDU+1XRLTBYkgW+99mFWosj/Vb+ifs3OoLkZAytT5V8/0DKUI0go+nPqZs5Cic4ck3l
8zvd+waJmV74YSbkZ3omnnblE1ZfEE3gXKKYUv+DmHmKeH2NSymMc+Wzprytip5WPFginxf6r+ho
q6lYvN2v4F9K86pDnOntVfBjpPRhEWMky1zdaOZRUhSRmxPe9HctWaheWF3TWLrimvifrqlMNYhG
B2KZgsjhlJ5Br850SKea8vqXo9XoHYAHPbJqKLFfzh5upo2muwrw9vTFtr2ru1p2Qa3EHlG9QVMp
VnJprqSt5VqlM2J95Qgj0XUc7iVJyVkcegm8oCNIDDSv5yKhshEvolt/UadLqowoXEknlIZv4C+b
th7gxf4LEP9u0VRqY8GuQYB7DKd48o3zYVGBPsTisnptrVpKcPHLonN8RIewt3DfJkmpBVNaMHde
Btc5b+89QbQeiV1L/ObMYiYAwuCuLHZJXxb1734gN4jL3o4UmkuVV6EDw73SW1ok6GaLPqq6CaRg
ecU3sNJeSzQBjhYzYNwIfa0bXs3Karw+CQoPOtxDDtrhDyskr+xolyp42mgz1onu257iizIRU8wM
vRXVKZRXbpRl9zUfKRx3p4YheB3NqgIodlh7ZP/hQSCc4gF5U2X+FMhvQVc1Ep/l8Ih0Dgx92BUk
uT/WB0najfX8GhicwypPZTR+3CC+MTTEY/atzYrjLt7QRILuAuYvYzqJOG7jCJOahf9/Xtts028X
zQsX6D7lMM1w78yBydJJ7ju/213TWS5lV96C0mfpnRaKzIiXjmYlWwF6clsRNUD/8s1ARZ4swZC3
jD7xWJHt03WachZALv0xccyqpb5HXs5uM/eo5a3gGIeTlEOPBtJ9tgvOVLGJfqefgdCZDZH9JhDr
d+GtZiRZjC3pTJOYSlzEflENN1DMULywyYjiO27DOS0H2LhyqdgRnHLIcjdTJ9DSerC3RT17MqfX
G/rGisEqFJ+STMHbYSc5ziRowfp99F2njqmVwtx41Tj8qrB7WDQn2Fe/tVOainPXLs/pbnH1uoXZ
H/3iCFGfBbvZDf8NEdT8xMWe6rjWCMsbdlFEQn906EA++q+9J0wgJfO4wfZxHxTcU5NYFdsaL6Ck
YoehRUbHM5TSz0bDIy/sCjdgyV+VdzcObWT3MAnHXmej2Utb1q3O+eUIC8L5ABZCBf3knnsMr+Bz
LkcBAUzyC5vNtdOm56owEyQ1lsY4Nh+k/qTZMGjjgUS7V2HsSaq5zJ0H2IdpwHVRrTZHgOb1n317
TeYwxm5hPFEtb2XH0EVG+DO0kYjkp7u0FIAmjSHQzSTNuWcriAcPtgfbGMQmKaBd721SJ3/Ovmk7
Z/jf2zwg83FbhNdCKkiBGvkNq+MxKCZ5h8NxmBpNb7DTpy7lj5d7ue1fg3ycKxIlyIxlKbRgvTLd
6XTJ0tOGQFkQsxhirURIaY8h+BYDJZ7CL5+vCCl2xmyD0M+QatU8nnVw4vYe/0WWmQ71SmtXXNOj
sWrUkuT4H/ETPJT6j/lCX+6rFFqwX5f8MQ93EBcmy8CMjLgV4SLcKq0EkdtWvazrBoVVEMdAT5kz
kY4HD9iQf1zLkThQa1i1gQOhwp4QORhXJuCjBK/EiL/OCFeUE1AQHx59KSalp/CefgRT6Qn16wMh
UVVPI2qgeXmK9r/wKbU+kEr8OI7C6ag+RjGPLQEzq3PX3piALfPSCusHSZTn9FLFegma1BPEsZbu
yawa4UC4QW7Qva3+spWukAHPEc/1k3bsGtTK+iKhyMKXp2Cie1gOJY80+5iSKSsa55xsVUYTcR5i
cjtRPzST5+JyCTs0wkzrogAWT1bUWHDWDp7QsUGqtt9G3vxiiSjwRyEe00itVrN7t+iWKSctUhFP
AbDivlPaI5yyzhzrn9Fy4Ddr0UAEB2lBtfvBHSLAj/ldyIAdItwv9UZ7xZ7pXIBlVFkqjFz0cZqv
e9O+d6g1RP3WU6jQuNsmBtmtLV++mT50DbmzfVHRPtnyCSaL2AL9fMJJgr2KL7xTBMcXumpTFWQi
aU8B10829RO4ba27Uvdn1EBGbWOnpFTKuJ7JcK/Mi+I1fVzECiPIib666CZl0et6Nrf6swXxt5dY
XtKd62ffkqjbhmw98DAX0EZExyQtSPF0THB4WrbWbwHgwisZX1vnjrxP6XbrirENjh13o3j8xU6t
jxRJo51xsaGXAIygbjEwt4PiRDoM9eqrjyeDNWyANPSSDEwePB1Ha3RbUXDVq14akgMtizCiedDv
bh55R9FIJ0H3d3HfnwFqjR0XzbddsJ0AHrB2XKusCAcYQlbAroG3G20aC6NV0S/CaEaKvdRAsIsy
ZA6OBwIKW1aZJgEjKx/sECn8+YF2WxEDaunc2LzuZgfj1Wo5M9NWxNWV9bbXp6Mncxag4wimK24Z
gF2XChWmOlIl86sETKcDGixGDUZikuxkBsWfcxOHI+9ANQtZAgFJhwgq281pDyeKPEIQscs0HfLF
cMVDZisCJQF2kdg1q0ZbabAW/9B7BZintPRGEA1BUayEEmaWfHiKFRW2fC38lcOgHiK57rBaSLRO
CPhDnE0Ql3RIXdsBj5yZ4EtoF2z8MXR4Qx2aLOpDL4IgH07pni3AMYg+vCbM11GQx5FwWgQU0Iun
5a1666nF6yZHZVOozSN/p156hHCusn3eVCUluQkXygW38pZ797bxc/27uhYbvPFm5Cg24kys4j7U
/hsj4Q541b8yc6cj2LndLwxSb07w5ycypIsRqd0zpjFlau6hcA+rRlrkX1XMBIhfmqppUnPopKhW
SD+aPnH3C6Cn8DpjvodwYIsrN9N5Dl/2CrJHKWyLd90bBUFwXuIzuHwL1Aniz7LLY2N3rHS6wEaZ
JC+udYyQkp3l75VklEzho/i7RVrasfcBsvCL9mYpF4tQW3gWjv7EWiIygneWIkMDubgptIsYk+B/
k1taNKrpZ5iOP5sXrXJVwwyxQbBbPEeTA+LfJP8IUQrP3D/F3TK1AMQHboEplROV55ngaflDl59/
j5piBXtq31MjJiQH0GGxHdzvaBD6MftJXd+GUxJELJnm8IP9vSA7HJ1LbXtLwTEtbOAMTWiMbPgP
I4im8pmlro3QT5NMuU+KqhKfIZeTdFEay0uqAhi06dkpok6wvY/aIHRDU52G8ChVJw+5NeRDnhde
sqqPNFdlCGcZ7uR5J6hDkxGxA8tIaG8Kz+S0n7FpxgZwClXEWwA2fC5Vwqxo96ES/4jshq5Yyix3
RPMSiZqPDXaYq5AwjHs4xAazGW+Cf2e2rczS1fAC0BGiIv1mg/0M1Fe222lYlgFcBCzlJfnfTYxa
HGxRAVcklqWTViO9iU4NvdW1tkaGkKAl7x3LHx/3lKhVopDH6RKl5ICgAlzrB7GgvX1lPtXkQqaC
EjCr9026rvacShBUdpGb93ixYWYLoaYkW/1TTLfmVUL9MsR5UCm6CahbtQmC8TUIQ+K0EuoTTmyi
03P5w2OAUUcNtj+sI/dOon1YfL4nPQY2iON1zxdPLbTuQ5uskZtKlyCo6iWc7/T+AgtUHzDZea6E
nbm9AUxl0tgcqjULEbe49xv/Cfihls8MBdsaZXS0WKGQaOeMMjrnAajRlfDIBPpRT4PqG6x5YHwn
jlwZAfYUq2e6UwMAcHDRSmyx/WqwkUyhwAqvyofEskQSYPV1xlk2GjTrWp1h5ZYxMKgplX+3oSse
fQZsjoJsBIfBlVBnD09I0WJETC/nzTO3ZDFAwI461btV4fVHyNiBLYQi8mBYWbWEXgWq75VrW/M7
e+UWr0vNTvGuvfzPqIwpjXrodbg799lLZeSCvQFkI1CcmyPVpi9yI4YmlCV+dExz5SgZ3yah0aeU
mPnk8q7hIaOs7j5+T+xwL55AK/4FJkDTBIuhos0TbAA2BYkIC4ew+5gHDGnlsaYxry/SCK/70pXi
fBWAV6dyzeIZeU5wop1E/NOvgMQENaukOCW6a7RA+U/jhd7vOksT/NvvH/6Q4fXRrgf9sun/KEXL
cDwajw+/EaO7J4BBesJo5i7ghOHj1OapfQ0CxtFF+ufWmJYkm7II/Fh/QRnIkQ0FrW0kMDrDktXp
f/jDrA3Vho4E2PIKhrTyZE2CVZD9sd5t+IvZprij/Mx93wwxmRQrhOfMw3kqj/ldpAdTaCFdKDIr
/JXZ4fhw9K43klq2zg4QlWhCQhlk09Kpjea7TRO5HncuKwXoHvmNvddBiu/sOmg+OrD4ReWsjlYP
RnAmGFYxt6FNyMj5x3cK/CgEpWFlE5XgaayP2dsrfklhYP/i8s+yOiMEdNNx8SHt6ZDkCGVPLfg8
XVZiZ1EyEcHDIZjUbbHNLm7MlKFDzwJNKpjjDy/HbcyUFAmAFh/w1wZk8Ba/D/GyVvrqVAWjfTZH
2D0d7ee/Gaa/fN+d5tAzmJvaJsnqnOHr1/9l9CTB9qaHeSbbA79pUa/30TfJwrbNSnulMgACA36y
ry/C64VnWxBfiygjefvxTurSxEECHQv//fuoThgta+cstGhtjb7xX+YzXCNXgq9Lx5vDQ7aMDiGk
2ppN+B8hf4D14O5AhXbAH2DEj6UeuXADEGfziEWs+yH/l4CZ0k5XVZbZ0ZDWby6CKyoezzA/a3CI
JLPOXfoMC/N9KnsSpnK2cdQzBlt/UAnPwYI7a6iTRaGNw3kAJ1E7pN4zfw8LLqdmmWLu4SH4vx6t
XZPLUg/tunCYWgWuI6YHVs1wrJhxWMwa67ARBvuQsfdrw1j5qmbkKLflAOaPqw9YF7WXB87aAQC0
WKHcReZ7jMaQEXj86ndxXLjC0fWRuQy/UCVhrhctIBLURAalwfSvSYCQG7PoGoX50+CHUmK2DCVQ
cuijp6BCEfv3JvlPJPYnbh3HWJGovO4SSabj4BzplNM1NoXWoJyu5kG8XL9fTWd16160GIFXypJI
yGa9trX1PXmZuglq+WdsMfyLo/zY6Mq9egsofgJ5YFUmRkt/BpM4fIBnBWD66ZTk4U/OXp6VsME9
vx/45SLhyMPnV7mpEGcwW6w1rdTFgmAxVgsgzckC6nouvTn+wP6uGGBqEQwGKwJWrZpOxNG7gX3M
JIJ7hXr8QL6YaJZJoXbSIeE9jKK3pnhD4/JQyOXKoAeJiYak9vFPGgPGwQ993UM696WrRtX3gZyI
Ng2FJPXjh5HI6RtQxb5JwtcFRU4401DoSGu4OgYXq6WYKE/PFoP8B39BgtXliGwB+p1Z0YP+hJhZ
mms77SG13WC0xWyJFp4QU/XkVIxwPKOMvc1yJ8gyHxoRp/IfKAjbccm/U+C+Nt2Zs7GDWS1ltKNg
jRbP39xH7p1z3hAEehXA1FX/MehCxwAMI0RgeSISdZ0EuVN+JH9jnp9zmTQMEeqZqDSTRJWESLGl
v91gH2wRNgQvk9mkx12ITdlj4s0sGGVqw9POmXGArfGuBhYYwgkSjfiKFwNHi5ScCSi6SXbnAJJS
Ybunjs4isPeA1rLNKiw6uLCvN8jB7ANRPY3iaTV6v0Y28CVkzSmvFghyO4+jFuKAtHdAuuFjNV+1
fBjyyt/8BUAM+Z+jkZusGulxEpgkU0GUZKxkm2OchRKkDaIBBXkxFWqSfS02DCT5Ght9uiDBXEiT
nBj9XRWVMNGc1vrs7VAe3Lmcz0n42+ZKdjRO8j784hpE/JFnDGuDN5/IGnmRlnslcV3//hGy0lgp
Q9rGMyiC+sMBxhmSkd+MLC1X/xgmeiNUMD/3TYREj7MaUOMppNxXYEOqDO7GZHVmWugkuJz6caPJ
jl+gOStpZ9ONCWNX+l9Qrk+4ICTuAwNwSPisJEdRsB0Jk59tSQnto5dcOcG7QHahm8lJJ+tF4EgD
0XL1TwyQNDIfHH0b0dSvB+xeUjA0r1EzIK2Ja+NKBoKr39uXmjsW48OuqcqfvKjtusoKuAoFnpzr
JS8BKW3sAUgjnPlEVGFC5e4jaJxtbPbC3mfAQwDHiqIBkUY+J71oQBg0XA7Rb9NsHFKgXRorp4P3
NRxwv5+KhR43Xf94w3fxoZVomN78A4AptIAmOcUfkcc9WuuiZh94dwegUySIEzxTG79TW1S118do
HhB0riV7A6WjiZSdldNuCtLCU/foWHLcuO0ZVKQ5bVgEiWLKUgVxl2h/NojkLseeGJud6iHpPVkH
XDRX1f5XRwXClHBX3t6gnSd+jS7yAru3/hbmF+ZPvvpOElmsv7Cc8gvhSNK5mmQ2brYyQGGVLBNH
lGw2jB3elDIesacFPDSDXRgRXxi8MzqI+RwJZUTb0YBhv8BU/TUFH9K1AA+2+teN2XcS+MUxV4Wz
I2nLuYegxYc6QUPFXblCiNgBwacrC6wPP8RLPJ9GH1scubqipJ3YpoK0hmf2bQpXGxjHSf7MdgcD
P3IW0zGaho5D6DkKG55fCGNr6NO7fg6aniJktKXcPrZW50HNkvte+pD2V6zy36Gq4dIOXtfinzAX
d1ZHbhL6cNBXWy1qJ+82LSSPf3D0Es+4lIcn5KWWfs2qL4xN0u7kkwwCEHQjTGzp5g8HJWP+iu1g
W4idIH6pjTXhxKK5D649sIUr4SpEgnsQa8zH5V9CJVl5dYTT6H64iD6Ur0hAi1nml9ExC3I+vaTT
0sOU0dFEoLYxoMmbN9tLhIaIkKKB9p3E877egD+GYM8ahyJFquhCAWcwalGocRj/paEKRfQAxwnm
kRpPNDNnZhI555qom0fkbZAKEYhLgXtp0d3z3kRBM4xho3YEjSgwR0mkFZajKq2bOjnYRC/fPUlu
GuHuZrZBmSD/86IZdDBBMYHGtaOLHJORbUpc030FlIBiUluXyLjJkLEStVi68bGk1go5ixV3/scY
sY9y4dOpnXg0jOAgXBxlIHcOKJw4H32l190nhzi6gF1WM8rqaGP9ebudTnGXGwrjVW05Rwk3liB4
pIauvm+Mgiw6B1NwfWnOfb7n75BCWipYX9huCckROQ0xh+lY/rmbu9mcMNQoIs0cKUjYyRwe0ucr
mSMmbVY65XIo8B7BJWSUU5p8YyxVXCDlHGAOMUyiQa1RxVl5KhhUJ+phjWp2B2CSEkrufk7Qeg6x
aHZoUcWoKEWNruYAKm9kyd81FED6xDlicOJLbwVl93XCgPAFstSkZEQRwonFxxY+Mg2OkHFY/shp
4BMHYXoo26HWq5NDr5hl7TZeNMVGb9eu8SNjiXHl1bQQ8qQCdR6gTWzi+Ek/en1a7f5L/AeQU1gp
Pyp1K4BMrrzF2Qi8EQrCReNHR/+2m6OEDuRT+G3aWxrQV4VtMRZX749myRxSFSPXqtK2fE8lRD/x
rEMWkSxwrn0S8zYwYp6jdj5wcS3ay9QHv+YDk7AFMumQ6kuFrVaB7igEb+aPwPNICG9ZZ6Plzba7
376xFAGU5rZvX7hMCR6FuH0wcZWRnRSSA3VgaIyVXjgSMEV0wLFHSRYlc23Ac2HBegvz7AJjqOKr
T7zUpzcJDXUdF+yVIEW2l/2OWxfPLqYQbM+9UiCm5ArCQK0Y8E1uqLfYY1H9+wJAKnipkERwHlCy
jD1psKZRSXF8j0R7bSD8coIXvYb2LToOZesucHsR7FuYC5Iswc1MoE6rZlbdSBfe7LAnDzsbjpVk
BhSwypBar/Hr98P/yjgSku5amEFGaoAEwNgkXvn4lbfR/jkzkvtkRqz9Up3rYBo5Yh503Z9PRG4V
24DIU2i2A3d8St2PdxE7Hotu3rwaRC2Ht8AkObCLQvTGUyyrDmH0BhMgvusi6g+MOaA7rkhce4qC
o9ZQB0vADZYdOzIhgZdEFxCOUrrk1UxqaxzkCU+3KGGIhfNg7tDn/vRNh71RFxlXJTKLKjgj231B
znZKR1TQwdziR9DHfXH3cH6MYKxu0bxIfxzlzmFuSbAbd5RQyNYQ2UcDM1CStwhcYK+ck/zpi2Bd
wfdMENKP1ySnDy5IihpI5hn/dmjtMVPYvW6pqGMUJAZ5H3v4VpX7o9VMgDkLpgqv3GgygqdY/32C
lONhHvxoP075rCQYeFL0kq4Kz1YNQ9D/Hr5o933CPqqU2BCcPHUIR50YOmcYMYE3yfKFp8pqKMTQ
M8B5pD14X/T8oMD324WqLNmpILNSf63dWhJI5XzdttaKRm9gxXwDy/04tOiO9rguOLPg5vZTEdz6
3bHL/0QB8/Zp8GiwNn66QQLzVhvMRTAOGcaBTP+sysJ5v+It8EXU6BMHuQwZ+VXZVC+krsy6VM9g
6RRWOA8XnQxXuqF2pi2r7Kvu7CjhwcxVKK6aJMraJPOals02McH/JWlsahWzUcPBin4JbJpfQTpz
BhFSzswV67q1+fmlmSQpnc9FOUYBVDuLpzNXJXAOgcaHF94EjekHWFpFnRDtSi/U7VhhZJlMsURH
BMdFAWI9MWOwowB+EaJHS0eDnyZ185HwGNh1R2+styBUkCQEP9xbv6rvh7TtPgVaM1xblqnMa65H
GOeUR8SWlKkt/vHcuJ32USaIjwO6UumX7XQeI7zx6sQEnMCGoln6MGsJmXy3lqIIy8bq6GHKTM4G
nTumyZ1t6X/iRjK/calj+FbEClI9JZF2r5Dg7F2D0/iEa5mZvRoJUmqqnHTn0bPnmPosBTIpNqEl
PhVbsjLAZlAvmZR0C5t4ZPPIe1xjPDPYpBjCKoGeaa6wslX7NoGzeqiu5af30ejsDZy8YIy8b/7x
6o1RQ9bGYYEZmkUSGPVxL4A9Hw+aZR772D2TZmf0f5gLZIlcfv79n+HVvAOOYS0b2+C9fqUKbOIm
GHdkHt8Gf51DP6fBZfc3xlV3EUBnsanidMPCE8sRgpCp8xPtKQRi03nKpuXDjQWqlpQ/XxI5g0SJ
bJjKX8tC7DyoEPZL8VDW0iCz/fJzCzhYwfkth0D0T+Qek8iuj+ZjnYb0Cae6gXrzho+0nzOC4h7P
y88zI/eQZeQ68b3p6Uv9hWDoOJJwVvwo2Aaq81MUqA7MD1KGwRnu4Z96zKr+/DbpGXyHF+GkB/zl
/npY5Q4/FP+KgOPXrEiVxdLGCkTm3OnInms3/honE11GwI8xbGaH2yffjOyjExKoU5613Yw9Lprq
ccaifrnVGv9XGxPz71PF5as4A0mgORKLvUi0KE2ltlx/1EdnFRA7UTY1hdsHoxdJJE0pKoK8iSKd
pqTgPQn1/d3IKa/Lvk0F8t6lishjCIMPZ3URmK5xHks9U5j0E5fOOZfcgVpy1e8ndaSd4/GVPJPf
7NYvDQY7xPwn1Oxsa/jZj4xK5cadsBCx+1pgjc+qU9FNnlJvy/y6//YuC6vNI+DCsnzEBwfR8wxg
H4s9nK0nJRazQaCVGvKjI71cgiULal4Lck/gYrNTxE/3huj6GyiamTnyKgor5F56l8b3D4eKF6XC
qL58ueBRdRK+cq7m/HpWx8798yZ1Y5RYIBVMTm2KdKZzzSfiMZRTwA0c3T1fU+B/NBQZ33h9PwFx
SwH1xcDdbPMfAVGvoZo9o9zXjw+O0jwk45qeHx7/fcYjtCuCWQX7bDuYWcPtXYT2fz+kzyN81dBR
rUQDK7kPWDjWoqBtr0Qpsoz19Xcy0yEAVbloMSupA5emuwQsvCBCdLC4mjwmp3hqsPfxYTHGupcJ
UWoG3XjQPeWwuaSJZ9FoTs7WT5XPFOjlw/KAQ4ETHGE5GiCBjlpnLEOwKJz9G7RuTAdFC5eT9gCF
kcBXHIwPZSF20R8Pn8P97fcX0wPL+uUkmZbfIs7RUAsJAfmDw0q0mR1Se3KDCWRfUYxFaqaIHZXB
UA8JDqQ9Z+AW8k4CB7o6zJf3X7qWwtT4yYXxT9C30GRZ+ma7LugGPMloalNg6Tpx/9Sw4/71vB/7
b9OurWnA32AgmjvpJniwkteQpU/UgKitCdh7ajiCrv/OwCn+X7VGIE8imFZhefwSYh06saI9i/Vz
NfqZieygC8QKQUTv3RcWOa/et8Zk9Z33t+XP9Mi030MxFD/6dzawma5iKjlueeVSNTbcrgRfPwB8
yUlFq9BUlBQYlYXT+OPwheOCw/K1FG6QC19jAn2syoTDlpqpAwy4e6GRzd1x4oZxhhOKiFzkDQr0
huYYalzhVOiQUuiOTAmfpKfriIatAc7g40WeuYGPET+qwJe+ffn9LMdkuhZ/b43QOrldB6Gnfbg9
zzCpNqz4tYNd4+d/zvR6J14GCWU3aVdpCkcICA4ZkT/oYepFMRA3AQ/2w+a9onoxlkedcpBe6nYq
zBr4cvX1mcAprdEnGxeCpFMa6RC6+sQYOk8XWgHzTxhoZTnMSZa2Gt4zS6dy5p3pGcIapZcmnfFJ
iDp9aTawgAbqqs+POWnzI2gD0ggmIRkxZZWkIENe90gkov6j6bM5Iy3WnevHIuviFxtMPwXs3iKQ
plkfbXZ/rpfIaD2mNCB1lrNDQ5UC7rysIdiGvOL3mDIJKxrvb23HfICJ3Uujrsgp2cARDUiS8NdQ
OzPi++L5laf/b15r9C/caIJpcR5oeHepusVTgG9iujCmkq8ALW85u+KB95yPYOVha8W4PJbCJ0mE
abrmsfW77V/1oG2I15nTVPZy76gFJHR+8rCDzVn+J0VXiIJ3IH5T3ty3zX7y9kdc+Bz6jCEi9/L6
pWqb0SxpKdhFsK8NCS/3MUCx6PpVrug6xEuxyuqOTaaMCW5sS62kk+6r1qAaUR0I4iUYlMxU6453
wo9Q/hMte4FbshpdaUv1MEsQfUqN5I4lyuI00Dqhs95maF2Q8znrIAAx04L07sNwiisXTbxbgQZy
N9Vfi2OLWYEG/LnptPErC2jZxxQBqpCVpp6OBUc9v0m9OnAkDNU1twsEOdCGpQqbnncq1/oDJPzM
KuAkWcKiYK4vgskvcqfW3n7RwiY+hPCx1nKig87a8ZjminwiDMyst7uQuVMbRrCQfCf+YnpJirrx
2QBtRQ/GKUklMdb2WJAjaUEr2YIw4ogEnC/gW2KfyVs/jDLBOE4fSRNYowCScjiihn6Ky4T9R5a8
ub5zbN76It1DcTUQ2jFW4eAiGE4Cs7EUDwywX+MQsza9Jqfc0z6drIgcMYfUzDUOifRN3dAM0NFK
AXOGLJQjLcWfCReL+dLDTrl98VSBGA32IzKWgLJ3lDssxZnGh6cQRMoIOBX33ISZCFyA+PEM100c
2tUDsyfo6hEb5QubZJnewXc+z4oi+cdKkE2EB+dhn378mcsDJR00PlVxePkNN1CPgkFtwgNd1yPv
z9aS+BqfC1K/DNq5dgBCSRhd6+t9Yb2Js7SPonp6XMISUN9gXnS+16kTQL6DCtbT/+umXTJDoLtI
s2fpGONa3N0jVp/GKWMNus8S96ItV2UElcs4e0RIzdTroGiY2z0/n9XAqKNxhpZvmF5mDOoiwX65
Uz5l4t001o2JOmVao04i4P7MavGj0MCM7GBOtBkePyYi3Fp0MbpYFjHiXZlBuhlBOZyyoxH6zSqM
v8tDX8wB6ji2OP19rMbjwjBGR/V+Z7lyNdNereWprp0lktIaO/ZzX5Rm3JguMRGr+LQAQ2+GCGas
XQeBsEGr+31dd05cmWkGIkGptbQZ+QOeZeBpNQ+PPXa8Hb6/y8KJVQxTpa0A6wPFcIsk2PzQ7k6g
EGKvF2TQ0AYy01MmBUusPrdXvrVHecrd6hd+1DizryartQAJ0K6D2mM282fFCQdQywuOULayb+la
QFcAkZeVpYuxREbkKw1PIe2CliyiGAvX/yS1P/IuFupVntvxUO0ZXA1VvpUB6B7X2Je9s8q7AdNB
7Zb9D7IRUPbGzssrvJAH2pbBGbZ7me0vzQ3SQvYX8TdR6nlHJCS6ZNJpp6Np3sauUZSOxpbvJIIl
bvPN9TyPmdbGAUqthM8AdjLeSAS8HZbAV/BdN0e744aVN0nuqThyau6En7NsMVKdmHGFMJjwdoi1
Mwmu/1G07hJ2H/CUVwmXcVKg6tFG7lR+bGEgUCGsPCmW6VWlDukDY8IkuTSG/JLbWl/ACQfr+KRy
zac8o2XhuhBt9mIKFr4jgoAGh7kxZdpkOmfGr2M61Rm+NdZY12JnLyyYVumbitz9KU9YewiUeUcw
s56+WMplZpN8qsV6DcOcTg16Fi+FrRioKzivJQZM7fsWBZwF9ndW9DqwHfIIxkHAtsIpNmuM3ttD
A4qSuIngHTpKY1lzaquDgp3m73hkIQcZdWn0sGi3i2A3NODEZTytIkXWzFSAVRW2z/PMZnBBGLmm
HgPN5A3swLyUgdLXfzlcpb4STvUafBgKkrH62VbiNtGCRoIljo94X642L0h5ijQjkgQdqVxSAGCV
+/VOl9CgE4u5cPkOWpy6qgdMZHSqpDPgKJUBuxkyhpf59spXmI8JC6QOtV8wigLMpjz6rF8vihxb
DbmmOJf/Y2kG8eR7mDZ06g6xntRJYF7tCoVcqjKsrsEAEDjJT6nTGDnfHJWYF8yZ64TQ+uQLK49L
m7x1ZqP3tnjdCn7TGJ/ftl/RQxXr4Riv26ngIeqXh9bGZKvtOrehAzLCj8f9+7I5KNUf8Z0zqzXQ
F2VBoJ6V/ReedGdmU+MMGj6W0RlKdpKIhQOsJ3hWBqOBLrXrtC5/se/uPPbMAWUpYvJLD8VcOKa/
C6Jsa5vQJdK855vAjKFCCgX16rGeXUgrZ22FZ2ZgUkisqzwcqATSES9o3HIZAS5twYgtmHZ7tStd
w0fWeeO45XEdvq8H4ygETSTywZQYRTNL9GK9FGD1huBnwQ/bwO3IBowIxsH1XKXCTZkJ5bgayJv5
d97DOoAPH00r2qbHNHSIAhYLB6YlhX1szC8hKjpy2+jocR4jvQoSYo9DoRS5Sxgl1uS6WvIdCtxz
tS+etqE3R8ttrJnu26EQc6XGEkizt1L9/q+uCqgYepa0OMfDSoz8vkVu3aFc6SIA4V2EA6Bc4Ijc
LLwjU86guOjPY36FK6drQMiRy5lwMurhEXeurX5GSZSVNL3RUKQSu53XbMQQfQdw8EHFx1YTt7oR
8p4JhwZVWKpkn6tMOV6svPcxoCGrij3DA3T+YbiVrMJqj8Y9+IkAhef6D17DYJ7ZRzTEzdk7zKxh
PlqCu+WptHoYrgi2UK+2pir/JKIZZvpmLgurBHwyuvmaI0ZlmWGCa2xGkbf4Q28CUauzW9lnCqyU
Sxur2uYhno+T964rC47EZv7X+1gLWfz7sVmmYk/eQ3hvOJ4fXxz+lpWanwqy0BOjOwcOtVl7MW2S
vSrWKjTyxDX4z1S05ku59Z9v/xgVeMfuc5PNiju+4pzNk1R483iulLSs9GQhUo+McyJYsRSFF0Gn
8q19UoJuKrGDr5iLsVYDUh2sDgbuNE3e7yJziATt6v0clfN6+uUg7rxGjbrA4W8xVUohrEIX1Lhf
KhCPb317KuarwcpCl9p60AseEYN5ToxXYZMKKSXJ4+H2BcIenryX+5XN8dxLt/GeUm0bD0gm1F4g
/r64oZbDp5j4ADjW/L4raQJwDVheCHhKqtnJ0Iyr24OR1FLW35/2SNClrnRnGvtLWiCObKGYyvI0
eVGf2BCWI0eUoe6KtP/oBEV1yiQ9S5FBIwlj037CoH9C2PJZ6gGiJuqBD4z2caLjfMQzL1GpXHIz
2e78pZqJld26LZ+ziLSy1IQQ6SNyTcDBuGCTaxDepkIWxxNmT8H54tchKrixnDrbUAanqb/nBJfp
xVlZeJEwI6qeAvLqj33G64I4ezf4fRqDoBfX1uhWwaiRkfIanA9UBDiN8RDtnBaSd+VLd7lcvq3K
uBf2ztup8yut3Bx34XMT67SJZAkL1iZGDcteRvhiNIhWbte6+93jLY+Vm8IMYDFadkulq/NIGsun
sUsqOM2L5xXHnrUk2h5XHI+XqS0ZO/EUsHSAJHur1e/KzEGq2e+VvWNQecEQWmYLZn2jrw/ZmzA/
tp+klD4uzjlYaQbhf2BO2WV4tR+dzESIfdP/SiXj+thcwMTJ6eR1Z01VHGtWJJPitINkAaQhZjnA
vPYViMTeorqAf9yMBcvw+lSHZKqXRUdsLWV6cfhNeLH7aT8FcbrH7Q9WlivIoT3jqhDSqfsHVZvQ
KUZRviufg9UnyCXnMZKWQm4OCsOTCRo4r5JYZcOybrWy3KIsMBzcu0jrfLelBnBYBfbja4xiAodJ
xZCRiQDshnrZnXqm85th/ywU/UgVZZ326uECUQ1Q5oTGBxHKsH4PeSHJD4IhACaVgsiUsds5RUzi
J4CYYpga0/8JQTDbozOvVOjQlobmIdYGOYUKhmY7jlzr1u5dLVzOHPhp94+ISFtHDayuSDtTUBaz
1flPHeJEEAaOdsk1QMTgP0TZqeEkzP6o0HoqAGx47prmFP3CfBX0fpI9sdAOulXLQ4tUyU49mB8z
FRvP2/9kE1ttfv7aVN394siUUiN5rcxyFmRlA7l/wMEYm5NqIhXmyQ4YCkWmj0h4oPxY0PUor/4p
irH7qSj2kggpY/IJ4HvN5eSlahPvQGVfc9u/Jm+w7SZXA4wjUmoISonrTHIVF+cWAxWcRXbF49yr
EkoBeo78go3SGAlDmZb6T5zjl8+VHN587rIKvJxcgUuboTaaXCSexahMfIZiZpocvBl6io3Dsi17
kpcSoQylRJRLCUERxqltTpoTmwLEeyXrbK+UviwOo1AnCCTbM57a1d67dxGABleE8fZmXa1gRjr+
yI3bI/kY3R8u4ehoy7Jk0ToXkW+IQQsb6IumXkrAHBsKhMe1QhsJ0VQ+14igUSZ288zLOcxv0pry
t8H2oGF/oyhXlBpAkF7Me150hAYWYHeH2kyFnaguHKPqq5vrsYyBEUBaIhXiCHxgALLAI5jXR9ha
r1E82h9oXV3s7rEw1CzgPSU5S9YJZ0KOzD1FAmGzmP4pyP0tFpk07ihtzYJpYOk90noRAy/loqq8
ob7UxkEhC9+RmSgoRR+/V171rSTYzw7lWFeSJ/x45nRvjPGSzdes9iON9y2r1gMQvOvKFr+LZp1p
S4FJMGDECfo6m+4GwNpgaZJW4d+UxWha0VUtiaDKxk5OMw7E/u0eydmu08l9DM3Nogd0Qq6P+hsx
qFJPNVLZJ0B5XgC3173Sa+bA+lBAiz79MoIeDMpBbFRcQQeQ/oZezxRyQJQCWMKIr1qm+dVVmCQQ
TqNIc4KXOkVhnyRQk/TcXJDbilgDarXCal5ra1m8saqeNNfgBscJkLBbUSXRYQ==
`protect end_protected
