XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��D��#��^�_���Q�>0�Hzn '��1cC 	��:#M���NU��v�*���]��;_�O��O�=�[~E�i���j����Hx���D<������F���K��w�b��b���{���"�-"�	��-%ǟA�G�Ea>viΡ�`��L���3P�v��Р��k�.�k�y��!�#���ݢy
rCmY�a
�G�M�Ae
��$����U5|�hw\�+��l��3�ԡ݇x�a ^�i��'jz�q��ؘ���ug���(&
�%��Cp��ҙ:�i�&I�!�O⭪��D�Y{��9��e m�'�d�����k^�56�Z
�٘�v�媔U�on-�G}@oϖ�ƚW'^qcE7$�>�%^�h����U��܆<��*��(��>�q{A)�-��-�m���)�#���83M��:Ʊ>��j�r��Ah��b.�Kg	u��e�����9 �'9������I���fș��Iw^�G2h"li'2{��� E�=[��hGq�`�3,xֲL�i�N�KUI��c+]a�/��B���9k��m����Otb�z�i9��&7,#��Pk�'�JX��ߤ֭������h]Ts�X%Ҍw�tD!%�؉}!���|rVr=��{X��eZg��B��q�Ml�k�L1ڊS]��v ���2Rщ�.�[v�j���+|�B��/e�U������1!��E�<����՜�(�UAeŪ*�m�%eh�)ɓ�\�Zb�qc3\p�v�MXlxVHYEB     400     200iVp]�-7�=П��Z�FL5:Ѩ ��22���l�4�WX��r���j�o㘍:�6%Yp�-?e�͢)6�5I8�]��Q�/�c�T�=���3g�u��ˍ�&�0�}B���:V�i��	[򼸼�s}��fFhְ>I�� �C�юZt�(�@61��dS��.�'X��Z}�����Jˬ^�G�z��ן������B�h��j��h^#�fm���Ò�5kQ��Q�8�^]�%�ݺ=�{ْ:�!!>8<�N����B]c�΁�� ��Y8e�5:���	�F�-�E��匭l�d�z���k�:��2�.��Le�vX_=�4_48^d�M�0��[���ʄ��~�9�2�+!-�4�6�x���Q���1�8@��v�9�]��Y�۪Ɨ�
U��g��<�d��n�O@�~8�Vÿ�"C��\KA��&rM޵�'���/Rڜ�w�Ȁ(�SQ��m�'�Ȧ3�/j��R�����^��k�:�p��e zXlxVHYEB     400     130�?�;T.�f�F�Mc������@��-g����k�-�*�7�ʕ�zPā�2f⻔�	��~��\����Ak�����ƹ���-�o)ݷ�۵}�%��"��Uk8o��� N`�o�C�SG�|ıƕ*v>��QB �ivI��҇��v	���T[�e 0�}U��srJ�i��(���E��-Ap ��ݟ�U=-@3�[61`��c��D�Z�A�S�YC��Y�!O�	��(�'g�AU,�=m�jVH�LC)<�A�o�Sr�B}�o'{Q1��{�9>2�����r�k˄#}��G!�XlxVHYEB     400     120A�`��U슜�Hb�x؆��k'���s�6��"�G
ZJꈾ�Z��&���"{��W_���QM�r��_����25\�pn�R�a@%�XP�(
�9�Ͽ6�g���S�d��C�W�n���~�D_�-�e5_(&S�T�U�\R�ױ�J�1�ʌ�naEn%}I�FU5�#q^�Y��'YɪK���� f��L3�% ��~1��.���!�gg�{���#^����kD.5y�ʗ���<ao���! ˔�p���T�0b��=d�m83����E��[d�XlxVHYEB     400     1a0��@�6d>1��CHv���c�l\g�cZ}#9���i����T�X���/���!P��8{������j#zݙ�3m�fBW&4ɘ��;�O��k%��p2k��*���.+n��[��,d�΂��|���y�t��&C
I�G[�AMBe���)�0��Z BUxA{�o�A1���	�T�=�fTjD�(ւx��E�H�)C�vK����]� jpVg��j�Tt⭸�Xf��VM�Z"�b�D��
7�p�Dm���82&����>x�I�tN�Ƕ�+5R���C�3>m���\��lvII����������Q��ch:��Kr�����]��ܙ0����i�,�/O�F��|����q�����[Ɣ1���ۈK��1�%� o�e���T�J5l٭�}�^#���-�]���XlxVHYEB     400     140��4R
�0w0���.�
��x��u<UD�Z�L��:Ď�f���4�x�@4 ��I��Qd�kA�=��t%�a���۶��Q�a�oN~��*<�{���Z�@0�����X�� 7F�K�Ϭ��Uwۈ�>�����ǎ�E1m�Ё��Y]mIR�J�FuvY��0���;�#��ۈ!+b��?�bp�inRg�^g��۵�|�[�}R��P��3&*�h�u7)|lR�܃<_<��"���8�.e뉄�2ȑ��=��"������x�������]�!~��W�@� '�Lz��?��#���ߏ�%r��6��B�m�׺�ӿ7XlxVHYEB     400     190�`�0t��f�E�*;���p�	��k�x��X��/V�<�8���(�4�bf$�<0���+~����q����wLD��������Y
_k��u�q��N{<r� �r�ˑ�݃�<�T�4�G���Ð��l���`m��u�4=�/�KP�����_���7���,�Ϟ�<ؘH'��Y�_tcy���&.Ŷ�l1/ֆo樢Zy��M73��
��b���� >d!0��|����璃R�t����E��6畋�_\��;��m�M�u�Z�k!9:�c��е�%�"�o��Q�%�IJ��8�݋ה�=�h�rOQ��0FF�<KB�'o&���Wf��7��]Ng�b4��CX0�ɘ������I%�Ǌ�bH��[j�B�XlxVHYEB     400     170d9��I%����@��Cޣ9xJ�qn�G�g�Tk�Ӭ�� ��6�/���5�Q�����l��z3d�໥M�aT�g!����b��@��D@���N\�!��������G�0�oUq�K�����q(��´�0`�$~gA����[�ͧ�;���2�L}z������$/�x� ZEk+a���ܤ3���#ƭ�R���hM��y?�����P^˄�a��9'Ea׈�������8\�[d������������f��#N�٫�^r�O���" cX�:�����_ˢ���|9�3)*|������LFMH "����� ��/ge#����I��9��Ҷ��n��[x�1�b�k��;�XlxVHYEB     400     170{���ȹ�)	�4�~����\�'3bt4۾�iᗥ����ev��t�y�k�R2���O5;`�\rS�e�X�8� K���JC���^�Ơ��>3B��]7�Ǣ*c����ZX��m��6AO����ԛ TR@)��΍��K�9��~j���G�I4�ZQx���n ��ggT�1G`�%lD~�(߶�7�q�(LsP��u��>���m�C�h�/ƨ@�-!*<f����̤�,�_�|L����9��i�z�����3�w�)�_g�8�.��I�D����}��[8/7����{hU�d��1+dU��+�[s��e���4�������a]�������A.<�������?XlxVHYEB     400     1d0�j�u�uȫG&��B���#�`�<ɚF# Ra6h^Y�k(��Kj�m#�_X�=dߎg[|�(1��UI��k܋�TA�n�-�������e����B���,W�����R�<��J 2Ųm�Y��J�]���	5}M���%����-1���jq}�ե�F����֏	�4��ۉ�����.ɪ��[�J-���	rx�G��Z�9�؞�ک����*)WM\G���\��� ��A�H@X��P> ��m"��08�.�30Vxn4���i�,���P��O#|�s���U�X�q�ǕG��>��J�$��|�9�ᕹ-3�㓒���V~�V�������:
���/�;�.P�s|��>������`<���&6rtO+&E>[P�V�����OK�����n���'�y��vz��/ߒ�#�p��[*�	gd���97���`��~�խ�XlxVHYEB     400     1d0
�����UzҜN�^���
����*��3Lb٠s��y�f���T���9�R��h:SVw�[���\�i������hppR0���J9�6|�	�=.�ӊEu&��N�U���#�D�b�>��7y���V=P0^`m$v���&���`{q6�P�;�Q��.�,�m��IH�V�Y��F�b�~�^z�U�����bߓ��+�0'����f ����g����j�~�g,�0'-���i��K�Yc�99�~K��<�u����K�GT�Oy#��$�#V�2q��Z-�)zt2$}ĝ��x��t
�["Ԥ$���c �/�j��Ц�s���ה_�H���!S�`^;2��[�#��/�4����/qP
ۿj�������U��ʷؼ�FJ^wL���?Ж��(�d�R�h0a	��z��.��7O�)��]��x���������]:.�XlxVHYEB     400     130���CS6	�_[����n�/L��lR�l�N4h2�~'ma!
%w��ˇ.mv3xⒽ�5i)b�EW�j���'�g.XM�K'%^����0�����/����1�m.���g�v
p2��[o��P"dネ��%��*��$���9�4J�w�X$��5:t=�$մ���ܵ�K�����x<�����~g���)ŉ�3�+0��(�D��>�Ș�}+N�����$�A~?�ޖ�$U~�N��C��l��c,D��-��_M�@���Ǚ
�*|/����w�P��N�@?@O#K�J��:���[K�XlxVHYEB     400     150�N����ʢ��i59M���b����3�Q���0�8��@�p�V�<f��sQ����y1�Ő����y�5�"3%4��xPkՅ�GW�F�O/5�q��Z�+�"�J�>����&�G'�����5|���Ȗr[��+zO�b�ó��+�ӕ��C1DO��4f�I5��j��켒,^�E!ƿ�\�+��ź��4�S�߆���	�x�_��!��,����?�ڿiep]��me�T�˜C��7㷴ݴ�*�0ieI�~��X�>C�y�:�V'����fN-�F�h�;8�f�fTP����w�T�p�j��#әr.���02�* ^`ޣ�XlxVHYEB     400     150n��o�]q�h���$H�J/�u\W=��Px�Hf8�q�K7VIv��.i�({��
i��(H&��	�&F�_b4����P��p�9Y�S#K�y2~�_����چ�%�@fڎ�
���*��J�s�c�D�:1	U����Bf�T\�.	w2�k�ϕ�`�D�i���䜲R�Wj��e���0R4�B�{M ������G_��Dw8Mx�91�4�}�pXtmՁ�r����?��<�;_��0-͈���5K;	�a;n��Ց�լ����✝�k3g=�b�g'��� �����3�(�=�p��;g�g~��Ȍt;�E��n��XlxVHYEB     400     120MS�a��No�T#0z��M�%��ٖ� ǇQ|���3��6��I�`N�_f���&�y���qŘz�}����{���㟡�;�i��,ݼ8Ab�i���Vs��砠��ci=�t�m�T��h_ n/kZ�VԌ�]!1_?�Shoul�� ��e��ֈ� ��-�o�NI���e6|�]����L�B��tIM�e	HU�`��I
k��5C_�ԂQ�o�z�w<$J�o�>0b��V����eg,�R����!��g�xp�-U�������#h��h���w!RXlxVHYEB     400     190 �Ϙ���D�0�!�������֖�zlr�}��W۶�wk/�"��nG.'�a���%���� ���s�����~���&��^�dG
�Z��_��n�U�J*$�*�\��ߺ&�H���sJD2���G��F�W�O�D�
�M�"N����;Y^��3[ΙO�3��d�u˪����� 6zI��⮜N8���gYT:Q�~C�j�O?�\r�Ҩ=N(��H�'�d�����"Y`u��to��%�2��n��d�fJ�������}-^�f����v2C.�dw,}!E+���Cn�~^�4rD�d'�P&�g�;� E�<��%���j���Z=��P��ȲY1"�����((7&��U�9� 	R��e�6�;��*Ṃﳔ��y��X��%XlxVHYEB     400      e0�9�.�ve��Ь�i���*GX�8M���G-]CTE�SJ���C�a�����z%ͺ�:�'-�zME��&~��_���Z����- ��D�dO�ʶb��e��}�c"B��^oPE�|���0Jwj�3��+mT̡�oa�~K�!����Aͭ��f�˲=����O�!8{i��UX����D��'0��=h4D� �MIo�6� �f�����>�T����XlxVHYEB     400     190�.@�����Aٻ�t��杈T���5�D�0�+��՚=cZ�iZ�D�I��Mخ�el.(��g���	��z��ӗ���e�˶�����4�h��X��$+;���Y��B|�)�
=��8��M�FZĴ���X)q��+��U��Kyv�Ҍ����+����� jo����.�gǉ�Kk�?��ͮ��Y9�*2k������t�f_Z�0I���+p��m���8zm�,������S�E؁����Ch�Q����!0bb-��a�!Х̛�N#�%���?��I�m���F��a5��rCd���Z��-�?/U�<�lb�,[�����d�]~C�U���y��^�QANOZj�2�9j�0�Ȭ�-]����N�v�H�4XlxVHYEB      c6      90B���(IjzwZ�_�u�z~��0���5G;�����U'*�Y��3��/����t��%+e.��Y����d@�t-���(�rg_M�:\"Zy��;�Ӿ������6��D|c��1d���4�F̩~1�"P�S�%[