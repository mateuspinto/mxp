`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
xJhVfBWYX9WSkAtNPQq6tDFahbZBsh4ba/pt645cKtRObjzdiEJx75DSuRKU2MDgfdXQ0vj7mDyU
fs5wvbZGxqW1VZV2o+Psr3WZZOmgI/TY0FLO6H9xirL1DnJPSEsM30lCdtgcziL2s5pzlUel54n0
f+azu0hHvFydgJEdFFA+0kI6lWzNLKPc6vFIOX+aj1hZKZm62ogTk6+R3O21HnhA5xEyoIwh+qFR
NGbhzwPrpuhU7SJBaLm6OKNN/wmoA17u7Z7UyozKu8HjN+nHoKJynKRMA8qGom8YpJw9hXQr7/eV
165j+sMgjUXMy7z3nEGb13DOqOoP3S6YUpe9wEhnakYfHDQP5kMq4hPI6rTAgvu+P6LQo+NTF48h
wCmOthNoFngCegNxdOE8do9m6xp6Q9QPxEfeAYZGzW2RBesJiO3jJTUPphb8kaZWK5tcdRSIBKpw
wxAHsniatV0WWaQYXm2ekKJWGsDZhHQXD9RkxlvOgMlud9HPmADkGaj+3S6bBe0sxFXbJ6jgQRFN
SCweg//JPEo4WHE4EpwJ7aZHLUtgoTQasV1sl0EEiyqYFcGo/wGLTXWBtRPLUcSmYADulwvLN8Jf
5/x3xv0+VuggchU9Gsp8iH1yr0nJSEY5AE54dR4rWr6+yx2d1tcpTgaB9cuZN+sfuX8bbH/fhefq
PcRXjgDi8aI9pea9av0cRmi1MJ1hjGTqA4TlXyvjczD8+aJW9VoYzk3LN+X1F3rBMpLPuvq4UaRj
MQnYxazhrmozu3KkrmYPNuUMLPOp3s0hF2J46t7HzmvyUFORRJT7iyb8le0O1jd4FUNc8Y/76d6n
MCy/tH7ROEUHL0GYiGaA5By/JtgaCN1BdCKv8fx3QVVaTORAahN4L+xw7+E9QNU9TLVAe84iDjku
lSbzdzzK8zaqybKSFxnH8aw1GGEn+3TnyV6hXzDBmFRh/x5LNMR/rCJ+GtalVyD11AS81+91uLPw
eVqhdeOTO6IFDn756gEVx6nEXgVu+EEEEzAv3HaTQKftx4KnZgaAr259dVHOtdzK9hNqyyUIPBvX
FsNMYkfN+Y7CjiWcl66ILu87VFybYJZit2ph1PmsMQmrpdrHke/F86A+FDxjvhFufMx16VoVl1me
g9BRrQS+9ar8NvO8RQjVhOV1UbHBF1UTFr7R7oShfbgGGohg1oEWfnFCB+KvT4Jgklc2QC4FnyUD
Jf8NrPkRV7e358JcxoN05iF67ek/HgXH+bygf/T7RAvdbKkczph3CjbMHb22xvjGln9U4Ne4lG3k
/DQuHfnHGgITHTd6T5MIJZkr/v0qog3GppGL+94JdygUYeYa226VzbUT0MSzhKpHN3GntJKlDQP8
+1lm91TH8rzouZr6QCwItxOyL9XE/HoeSxOlZlyWj754vpuSK7rJzXLOBmXgn1GVeI/5Ifd59JV/
PZx1urwj8Bpwa5aaPXLVajEg6TItsVrjRly0RbAQ12f3MX9yrmZuVQ5bckP0sOeXHzpLZ8DuZBWm
fOWXh/ot7I/8CSjgoKAdh3Ue1oLQ9SSz41WmXGqVUimJCy/Q7fh+FULW9a6v/h+Foj01OUshB020
lun6cWsWTODkk1JsZf98EzuaROBkAZJ6iNKeUV7zer1/faYaWBbaOzRp5p5hfTTioHZr+kLIOwRX
uCjgGVDpRNgGQGFyLMXGxZeARyXaJzee2on0p2bran3z08tjTsE2z7cOzhf3G6B895bEUFrBf1gf
vG878Cs0QBtp+aMvskFTe/cvOjMXsTYpDKjqRtKr1FcmkR6gctyccnm8ylBON0R9bYMN9J3swJ7D
aWagAOzI1FriZ/A24Y4LapeVQINefLjGhQ03nmW2bMd3C2x8hp09J/VBx6K/UR62YsmgQ1QcPOP4
Q3J34ETMRnM+1b1dQhqHkWVOrd80HQq8cCUS/ZzG6MWrXarnAd4n6djVsCAVgTN+up8gYTjXs5s6
b76X96i2S1ipiWB+fzNX3M0nY08bjMCncUviV2bNiabzX91L5026vM+xHl2DeI33DS4CCI7On+lm
hhHusO57I0Yv0wb81LV01lYlvs94JeUyaHClqYi+ZxXnxyIG1fvWd/EOyh4/
`protect end_protected
