`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
UZLE4dl7cQKA99HKN+eydu+swJkxyuQHLYNZI0u3Sgfl6Kw+UTmGllEujvCgqzjsxxjOu7FZa7ym
KzQ6dhFFfyoLMewJEdXiambQ8q5DqjpBCuTWdlYTS5ZiLIKlHeR3odPwLeTubhPPp481DVUHp9fR
biPt2oeSoAVEtAhDtr9XzuxV2z4LR8eC8caynp6QD5nbdqcDScKifTwOBfNIrS9FclOt4Vz6JsUW
+jTR6ovFj+/qeBUs59mOV7Gklzqbh6fMTltU+2heF0H3AL5TWieGhdj9rC657T4WNVeVHDuYS/nA
rhL9hA1Plt1wtSkB/BOYimo7klI9n0OQZjBQSw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="WBairtn61ClibG9fgY6nJdc2+B+Ys8B3IPB44joPzOo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
uU0BMYPHAnKyrE5VcJb/0JLsbDs8q06ICsYmbmCMOfoE0P65JrXGgiEFQm0ZzrYnYalyQA2pAGvi
VY4tFk7tcTx7yjrXHi5JosZ3UguU+wzmMdEWgtpUOYrzh8syIrDz0Q+ayXrJo7UysuztMzmx83NA
DBinoPPX8dY+u1zLeROQriZuiXnvujaQMU0JYlvU9FDj3yK6yubj7dy3ctfv9ciYamoN0BECNItR
Zd/AwOMe1GZ52AX+t8dWdi6a+DOxu2Y5pZSIb8gn6xF/vOKqCcAE9sWE1LQQTKiQIYj6DKclnLoT
Nj9rd1QuNm60MRCaX3U2DXAjkY0CVqYwNbfcPkFVBuT++ml4Q+nk8x+DTADhoUjQJ6aYRi13dMEH
CRc2JKpKWVGXL9hvM1Wxv2AALXOvCkf33EpQnSCyyE3rSxmzRLAjyJxj+mDezenyizbk6nvWk9L6
+NurvMmB1+bJz8HYN1Ta0kMs1z4MpGkULCJYFv74SlkOQXjdbMVtsG/ggsVDWx7ZBHSXpc3LbSNa
OCDPnPDN9ccVqRFROwU2glnFzImsKMM2GtE3Z83hb7jyVivOOe3Fj1FM7lMlypQePmT3HRK5wnKS
BRJYeOSFw6IdL1z1o3KEAfgQFopnRWFZTOMZcqUzNdR8arHI5yN6V8tGTRGeLDTaAEBBGj9t7Oh4
sqrAC1hmDUaaDx9A7wqKuiocH1m+4DArEGtMtWGEt54JLSi3u0cmjQlymORtfGq1CaX9eh7WYO7W
A7CR2dmH7c3x1BTcSGjNNaPvPewq5YPS0fgnsS6KRyj/TSShS3GInd3a/RnJLnDco296robRXXvz
26uvxSJdmaZ9H3hB2yx1Pn806RTHbYhmwXX5wzlf6RkPV7Rv4qR3sDShoKf0jmsHUU8xkIzULVWe
geTx+jndlfdhrgSL6sGUDGAf2r8q1ELllbpIikaxSqQVDLDM0Xmfz9dzYuPVihe7N4NRk4KtRU2T
9E34rjhy5AprsIJ7D1mUiAjF6nNnrPLAnZgnTizHk1roj7rPYZQdo53M9MPtTrFBtfPCVRy8upR7
+CNWM2cKI9CKAl/OmYtmmaE7qvlx5V9ZWpMgGgYXpxcTP+6A/bsYjwQZ9iFNRTNEJrBEfuV+baEV
RGOX8cQ/Wv2ykAVAr9nN9Rr2jV04MiOnHNZFKpfeLjiQ1yHDwxfDDoChYriRQfk72dRRTQYaDVN3
ZrnDKa8CVQBRPD46ZwNfJUOnJxuphq42TdtecgiK+TzyLH+aonKl0yHgMLFAM2NXbJ9qxYjh6CMI
T/qrjeh1tiBO0vOOrc28yLMFyT/g++uGLKJOz62gjL6mqIBKxGnkUrxXO7TGV1iqbErdjZyUHtjL
aP7Pi9P+2zyfZvmy+FsBOFCMDD8CPlqvkFXMT6mVbDC/Dk394vc6cM3SpeQNLDOqOHuc5ibFrnR3
HMrcPekU5TRCfnEE+Alfqk7zSTIxMAbbL6kyXneNn3+vuMBmQ2/qsjL+JDr76KAQFKltQPm2kX7V
QmwL9+Fa+NMQ8d8r8ctz0KyKNt7+casIv/Eg2wskaLHAG3kfP9iNHzHasomTi5T7YC9Uh1FOzarF
3SAZ6dH3XHerFxqQDkWn/JX0/uMgSCPDCqvXhepcljnKHdPTlMx2YuM/lq+oimuiBdWbm4sK5qbx
zSRsBiJkw/6XoLYHRtJ4obwY7L7UpWY/Xq6c0EIJzzaxLu9hXird+acL+alvNLXqxSDiZJGtjpA6
j2udspSDguPM7c4BN5l31NaDmplrmtNTwn7kfhLQWeKmYIsM4KmpEbAGu13DXpgVWfrplTfEZtOo
XS2btXVqiLPRSGr4mzT0rvYVM0qs5kpWN/82HFBq7KQ0p/KNqbRK05WjAP3tjh9zdoTdC2IxoErZ
/ZjBWvJm22x0kfAVbWKdALtJlC9iagQxF4i5lRDQ3cLGgk3VgoCR03cYEQDclsnd27fWwgo9yawh
VFLcW6xTztlE0I5cRVGcECVYGA2algliuhwRz2+8sWkIcNCfIB46cCz/4nqP7vSRES2A5XcStPQO
/aF9e7beJYB+jAiAxmUwlJNHvqIk6BwYZv5GsxGruqwAyQHC+MRIU6azy4Qh
`protect end_protected
