XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����nn�#�>M� j��WB������Bjd����Q�
b�eJ���k�=�6(��%FA����)�"�v.Od�Q��r�G	0}߃\����ce S���/u>&ꁠޒro��P1ߺ���CA;_�X�JY�H���C0S��2��7���:8v E�]��]�^eW-�2�T�
�_^K	$�`��X���M��ٵ�k� �j�� �P�D�%���K���2�:<Y�:Ĺ��j�����=ozD9٘y.�!O4�g��?>��XtU�����44���?�;@��L�곦T��ԐK}I�Z��K6211ĵng�$Hʙ�M
P}�+|��a�iR��0M�,��a�4��e�}�W�y����v&7l�������J�sMl��ޭ�"��K��@p�� 3/-����F/X�.�b+Ipwʎ�>n0 H������p�Bހ0
쩷ݓh2l\����Ւ�©�	���Ħ�ҟ����Kh@�0R�7�h�n�&P���E+���Hȭ���
�S��lC\�K�,�+�V�4A> ��a��-4	]��m�V���s��$JN��hy��O&Ō@�ƿ�)�r��i�jTQº6D��n�i�[�6�
�u��P�V)v	5�o/fj#p��A�*����T���z-v�O'@{Qn�jo"	k�)Y侣~�7Z��������^��{Q���А��؊�����v�#\�	}��BŒ�&�?���"OI�t,.X��T�*{$x�j�OS�s�l�XlxVHYEB     400     2406�yvV���G�c��o��[�mk�O���7Mu����G�ҡN'��z8�!i�4�VU�vx�̳�a3� h��X�9t�d!SC�ObY������J�/�(C�/�����b/��"b�L�$$�諾g�Z���4g�~;J	�&[\��|���e!"E�U��?x��ˎ�p[�ܕ�F`��(��d��q<#�4�48����	��b��fac�m,/M�)iPK��
TC�=�ň�������X&ts�tZ���=��X����D5eU<}xF�Jb4M?(c	�������G/j�.y�Co��j�.�+�̓�ZL�
�<�j�����������T4������'�+Ik�ٔ��*.�K�S^֤h�����KK���`�������3���x����#Ao�%�@QsS,e����qs-�Ry�����U��-f U�p�3'���qs�A�/�jCb`4W�K�Euކ)ޜ}�A�F�����[F���ڕ�+�{�`��"\w��U�9������Tߥ�;ɿ8��82����x͍���"�Zi=���* �>0y �w����X������yxXlxVHYEB     400     210@�1���Gl��? ^8�t�Y��z5k�$�|�B�%JP���W� ��,!��+�&�|HB��>���g���/�x�-FdQ[�mi�\)D�x��v�[�i|��93���X��P~l2�&L��нA�i���G*��c{�‍�Cv7ɟ\��D~�)����:�K�*���QG�?�h B�𺦬fM-�ѿ��c0i|��s����mNsQ��!���9�u��Sh%��F�"x~��tVw��?�J��m�
i�)��"�]��<��r=�����K�����@����؛��ΔP����R$���� ��pܵ9�]A��� �7�g�'�P&�/�}d��G���]p߂��Ǵ��X�gQO�Y-� �H�\옞����|�\�)ߘ8�y�j�CȕS=�a�~HX�~�&:�"�Ğ��\ �W��9	�ςl�8�/:����X�.u0��j���}+�^�=�*!0��~�b�_q����|�T��횉\��Ar5��7d)�"��s���L2ASjG���øXlxVHYEB     400     1f0V*�� 	h)�+� OF�l�?8��Oj +�����v�[aGO�V(���8���glC:ru�s��Z�{�.�.>A�\��R���EF��Q�#�o��I�S���Λ@��"a�S�K�o�0�^�6��}�d��߉��m|�l��4�
O�pO�R1�����')�痩����&%�u��o�%���wFɐ���ts�	 ��v�!B�Z':�k%�N�l>䅻�s�(��<�]l�e��;\�7��V.%�%���]����P�Kp<ɢz�|��,=��'#���������B��}�R��@R�Z	r�9D��J!��q�Bv�7���k�EU�jd	�F4� ��_Uj�}�`�.q y�S	�⭷��eo΍�{����
U��(޽�V���^�G���#y9s0���
�l�F�1� �e��`�L�t�O��R���mQ��iaV��=  ����oI�*JF�Mȑ�i|ea�}�����]���@1�8XlxVHYEB     400     1c0t1�����,ވtU��b�Ƣl��2A�����B�+6f�C;^�>=�+]%�,������'d��j�<�@%e왘���"����E������[���z5�_�:�4���W���L�^x��DO��v߷s-��Z�O��9$r]'������lVN�,-wO��g���*�"s��s�擄D�G���<�4DmL<��0L��u��u4'�A��uI�G�e�%��i~ݶ�)�\�)p�m Y��zn�tS��:d� !���B�7�.�Dm\����@�d�+%�9�hV�P�i�{�*�9��$S���+� ����x߲��xk� �G�\�⽐�۪�����]�	_�����`ō�u���`:���������O�Z
��"N��T������?Q+��>~���g
�0�]>=Q�R�Z���+�I�׾�~i�IW�X�lUsjzXlxVHYEB     400     200M�*��"�R����Չ��}h %�i�T��6�'�u�e"o�{W^7(r4�Q�U��V&��%F���mU��f���@���v��*����jdy�E�}�:U�����A)�A�:t?E�����c\}���5�lg���1M�"*RMG雄������eB�k����Q+T�H�-�l��-��T]�>�������ik�W����ñ�f�V�;?�K:��Q#oS����D�
����zk��f�ү��qk��"$���ɱ�l� ��C���������4R3�A���x�s��X�����5�ѣ��  %fj=�˭�%>�ҕ��W�a<r����������EK��ڐ�˟<5��L���s�em9Q�)6�;e[zѝ#�������r�ST����¿�a.�/GoY����O�|�O�tk�zɢ���]e�[��(��p���8��Yl�$FV��(�o���h��F� ,�qɤc�|v{n�Fx�����r7���|XlxVHYEB     400     120�!R��2SL���HR�B�77��L��ӂ��A<�G�-��lT���53�Ā*k�<k����c�3�L\⼑Pd������$ܣ�`�����u�L�����k8�h���J���y�W6��+�`(�Pڄ��{�պ���
��J1���R�]z�Զ�Z(M+s���NX�������|
L�-��q'~�٥�?0uxN����d<>F&rvԱ�E�H�C`Z\2�ك�@z�G<�q�pXx���=�[�F	|�D,yb�Gmq�����V$^(��v7��&�wXlxVHYEB     400     1a0+�*�Ee��j�LX`��H��ϸ�a���ib�Wr�]MD��JV�d�a=�8���V���N�7�1�,.o�}%O�ŶJ����ֹ�L�����n+z�Y�p}e���֤
�m4q��Kle��?Y؋ݞ���4����N
�3M��_m�&�Ө{f�CY.�ڥ�k!�(�?Aꄻ��gV��sC=M���*y**��E�?�^����1/s���C����Y1��4��s��Y�� ]��96�/�f��X��q��T��q&��=B���5��})�aI5/Q^����KzC�<��i��P�َ��\���J�8?h��n�ŗG���i4�F��ڨPg�Ws����j��ղ)�4�O�3i��Q]�z�Ǚj�*j��["�7�4'L	"�XlxVHYEB     400     110�t-�4�����<�VW$Y�S6`�x$^%BI�eR]f�v�����[ͣ�O�)� �]���;e=��)s?r��ӽ�]�Ԓǧ�Xr�9PMӎ�֜�e��ť�[D����T�pWS������_�Nz	��Ym��oyY�Cq@K�B�RZ��FX���5�[�Ɇ���]�eJ�#���+��F׾5(?���UZ ��eC��b]���om��-!�h9�ʃT�46~�gg���묰 ϐ��z�������I}�5KXlxVHYEB     400      f0J�T<�8�ģ��M���ꤞ㦳&��jYd�eBY�3�/�=�6�YN���$q�[�l���>&׈j���ԥq��L���LQ����7lG4��g��R�ٳRkH�h\�WnBs�4����{�޺G�1n��4���6�XF~��2�����(��ck_e�$�j�7��k�	2s�B�8%�-j��-�Hl�-F�_�����n5��X�8� ��be!���a� 98�$:����<�&XlxVHYEB     400     130n���r�<�hھȆn�����k�zU,80���s��/�̔�YY
�6� |��4ҋЉ!��Я�y��Q�>i�7'~�']t�����Vf��1�O��n�W����j�h"���A�`	�mԑ�7�m��^�"�j^`��*�}QWr��T�P�<>.�
<�^�GLl�$_r��ktG�)o�f�Ŧq���e
!��VDD�(�z���7���\Q:vQp�@ML���;������T�-s>7Z2��8v�^c�I~|S�rM��Gq�qE��$b;�a^pEhΡ<�uG��eܳoz�WRH��q9XlxVHYEB     400     130c4��h��8	�fb��T����1 �\�ѐr�����P-Ӫ(��"�����e~���߱R��e��xjt�p4�!��"��i=����`�,	���JzQka�u�d������T��8�w{n}�;�}�)4>\�3Q��LaGe���a�#b�;>�E���~x���/x�i\�[�t�C�K)V �4�E������'���B"҈�e�Vs��a�8`!Yb�ө������\�����)m��*?����Xa;��K���R�6��*fi5nԛ���n��z+�H��g޸>�S � nXlxVHYEB     400     130����k����.�R:R�vb�:�4f��oG�}Z;�[ޙ�� ��:�O�H��6��萚�P=�ə ���5uD�>&���7�H�k!𨳑��������	�goh�m����bqi��E��^hR�-EqPn5Yo���d�p��챹��/7����PR�����6�<�T�|}z��[brM䏧��x*��]��5~Z�yΣo�0�ppQ��^]��{S��������{e�h�÷vG��\����W���L��}�Ru��}�p�Ŗs�:�&7?�C��$ƫ�l���|��2�HXlxVHYEB     400     190p�9��ہ���<G�޼���.B���W�l��ٱ6ѳ)^nw�غ�Zp��]dO� *Y�U*�/h�N錐\tٻ� ~+ZxB�Ԋ�'p���N��t�=r"�ll\à��SV\��͖V�V�Щ��&���X�G�t�,0-��n^Sl�6�uq�T]Vg�AD� 07.�چ� �ln��˽���(0�F�W%�:>܏p��d��}��K-Z��i�"��=8�s!j��dWqg&�'K�'zbQ��F��Ƅ����=�jFr]���f{,��&����؉�X�s;�cو��$--����M`k�p�]�����*'��L�]�KgFx�x�3��������<A\l3ZF�v�)�xxpy�	#F� ]ݛ��A�d�y6��=>��XlxVHYEB     400     110��Ǳ��ׄ[�q"�''���Є��X�M��yaQ��/n��:����,�݈�j��P�ӄ�ă����BO�[�h��}3E�6���:��%C��HJ��pol	�h�^�?L��$�gv2[X�Y���o��Z}��Q��oi��&�{m�e� �đN�IK!�ѧ��GP`�!���Q��H��*������OZ����\��h�0���Дp�2,m�N��	D�(�9�z$�����ɟH�п-q��O�111��W��p�A|@#����*��r���3�XlxVHYEB     400     1b0pW@)�5=&-��m<o�Z?�?�ë
��엒t��*�	.�S��6��5'��XK�|��۝��|��%�g#�.:�h#���l��g]n�?gd���<>(>����h>I���� �X�dL'{��>컛�/ć��)\&�������o�ݿc
�c��(�ii��O`�T�dy�O�T�J�~���S�E��s&`��3 	@2��+X��׉i�'����[��H�8I^��m��w^q�ƕ 0�-�C/��tt�BX�se�z�Un].E�L�����2H��=�~j�"����g�w����_�3\l�Q�J�( SЎ!k�2�i凡W�dS�̆����9�����2�}y�hĔ��� �L�r���$Wؗ��e!59`��IE����)K19Zf�G� �Aaa���@v=^Em$�"���	smEXlxVHYEB     400     190�pn��)w� ����s��{���U�p�L���ߝ���!Ʃ*��i��/l&�fv�|h1�� @ V�(���a�q���ʚ��~Uͪ���VH��x�L�f�n�ߠ�`�=`Ԛ_e���i�ld���~��[jX��
"������}g����=�A�۰Ībb}�ꑦz��%���Q��j����mLoMA�"�$#�%�o��참�����%�{���=�SW�~��VF���z?t�8�B��m����#V�e��!�Y��Njƨ�lA����|R�⌮[R?�3�����I�/���Qمn�]�d�,�I�p���3�\FU�r;+�c}�m�T��z#R�WsV��Iϥ]z�����ɳn��U����tǽe|���F�٬�XlxVHYEB     400     120%f�@�jZiP|m[aZ�=�F��y=�����B��z��u/t\0}�pAhs5�l�3���JV�h��Q����I=��\��/��dG37+��4��vn)f���f��^T�=K�4��T֫�n;���;u?:�-���&�	�9�ϋj-q/lٱ�;&�A	�������K#N�iqn��Zr����W���77�Z���{��󩩮�� �?az�6�H�HT���"��UQ#�pCa��=s����y�2�65G���f��b�F��x�"�;���A��V������j�]KXlxVHYEB     400     120�(��u��ĐN�,(�:nK'ba�Ŭ�!��r'�|��r�-n�8�iݻ<��:Ԁuc��5� ;�K�����eF%y��#�\"n&n������L6��,|���� @.�j�����p@��PE0�!x&�Դlz�Ϝ���F	���b��g��\�v�X��ʽB*���g,U��ˑ�j�v�i�z�ԇW�3A�6��G������2��:u�����}To���#�W�as�$�W`��'���B��'�������Ds}�M��K�Q��eD�W����eB3&U�XlxVHYEB     400     160�r�������&�n0tv�g�+���h����EJӉ���Tm��X:�ϝI��~L�r
��U��/���I�G��Nq��C����O��k{��֗����X��;�_H���*�z�,��n7a�7��;e;&625F��#��kv�%������H�S�+��)*�*�^���ٞ��������}��9�{�~k���3bZ�ม�w'�hE�n�uO^{�RxkSkS�u�㰋*+L���e�����I�����wa���cV �й�'�g?z�x� \�tU��ty�ALi�"�@��w}9�;����y(����p�/s�+������R� ~a�])0�XlxVHYEB     400     150�Gnvo"��~��j��W趱Bߎ�����}�.�SrTB��e��;� /�^��v�,��֋\��e��������KUy�0����h������f� �[�
�Yq���BЌ`�E��$�]e�3N`6���=�OX��Qvoj�W�yo���0B�<H1�z���%BC[9栿jW�1o���{n��E�Tb01��28UhSȌ9������6�"Ge��+JV!����;��~�E�ETl��?�d��ېN� l�T����TT��z�~Svt�I�#�j��R7tI�Z���ʦ4�w�O�X��%[�D{�2���ؑ�ӥ:�B��i�0yjw���*j֢XlxVHYEB     400      e0R	����>�1YtJe��~�S�8һ�p�	Y��6Y#
$�2U{��}y\^Ժ���p�����5��߮�.��$���?޻t�V%��u&��Ee'�����\�Xu���+�	���>T�����Xq]#�.�B����������`���yGQ�	{R|ɪ}������_'��,�g*t
У�-;��/�nH����^�ŉ��q#���� ��䙛�XlxVHYEB     400     130"q�M�ۉ�:'s*Wy�˪��h��\�B�ER�lU�ҴX��էe��F3��MqU`zL1Ƀ�ԝ�:���1D{�v�zC���7��%��[D}0D�P8��SYMv�Yet�����/}�EX�'%�<��"T{���@/��ZaA��B�c�+����;g'����k�z�M$x�T`l���Q�;�C?<=���H��R��h�k�&�I3)�i�W��|�4�@0=��h�A�$�p��U���h���Y?��(��-�=�e G�g u���>*7�bE���{kP�DK��XlxVHYEB     400     1403'&��r�i�l�|n�'�9~U.ڮ ��K�Hn|�����=S��s��;b�%d�}�>V	xKO�)(*�W�_'U����W�H��%�Vҳ��G���z�9d�ILP����C�i��hc���f��_�0W�lY�uy��k��� ��1�r���禈@����?
��z�X�$3$�/�ά�=$dP'�L\���UySn��O�f\�,���e6H��b?WO  ����5v��d����&�PJ�zȌM��n����^㪂��|���[?!��k	�g]À<���ji) �����]XlxVHYEB     400     150�*�!;`��zj)�Y<�v-x{��*�U���gߍ������c�����ֶ=D���Kh��<@ݖ����'?� �_���v{An�f�/C'ScS9;@���tc�a��cvT&�p[*]�&�Q*<�/#�SqG�f�-Š�<��G�P�����~���I+Sv���Q��;���_��!M"�m�"�h(�Y9�
2�Bu ){��80D��L%a�� ��g�d}+�L=3dX�����f��Z;�w�Y/�Ev��8���i���pˢi P���K�����N��s�x�kʨAm�>x��`��b�WU�����9��Y��Մ��XlxVHYEB     400     150���H�б|�c�ۇ�@�lvxy���,jnpꎞf�՘�Ѥ��i�ѧK�x��3����sS� �����#�����w'��V]�#�R�#6�?�_�-Ȣ�_Z�-1����ۮB��R~�Q2�̗��3�4X���D����%�*�c��� $Թ��mg/{�*w>�V|��P��Q�'$\�ܾ}��l46�jU9Rg�^�*Ǽ��']������%&����Fm�n�{���X�-��ju�`�RT*&)e����I�g�L�W�[(�#ik@D֙^ڌ{� 4�}^��-�j��8�ubve�C��T�Exb���^;Ӡ�	���#XlxVHYEB     400     120�֥H�2�q�5�z��<����+�Tny�y!���;�]���������t�}a?���B d#u;D'�p��s$%jQ2蠆";��x��Ej�;8SZh��-Ֆ3�2=Ӟ�`ݏ�k��L^�&�o�0�Z?���_ݙ��@-��Z�)d��u��2��:���?��!�EV�6.s�mI� W�-;Z�~94F̀EN*��sA�/�4�st����ٌ>3�����vd�D�,�%p��>G��� v`�^�
/;��0�N��itp�*f���+Ypn�L.v�3[��J3XlxVHYEB     400     130?�3�V"�5�0�"��EG��,���ߨ�~�Ғa�P�N7l�o��k����Lm�D�y�B2�����Ԗ�KOH��z}��6om�6\��*��[���)s��c�}K4�;�Ic[�j{TD��Ήh��b��< �؅l�y�L6�����`�f���@�LC Gh+��Ą4�=�:M��,
Jo��&d_'p�QZ����^�����8�SK�4�=�����޺��z=H��\��E�[:��b�M�9C�u��շo<Y�<u�ȥCu�}�ނ�<�?a��̸kXlxVHYEB     400     140G��->{ԮE3+����IS�mN��/�9�4Ҩ4
���\��|�-������a�6�gB�:N}�̆&����7-�nƀ�^q	���d5(tG�D���֊�ܞ�.�i�h?�Xb2�)��"G�w�ǿ=%���YRy�S����G��F�M:9/���ܥ!�9��#���g�V3a�v[fJx�=��5��o��:qm�����V|� ��57((�f���J�/��e@wł����Y�S�2�<��O�T���&K�R# 0KN�{U��5��Is�\�n����bl�����b�*Hb�i��,}� �]ϋ�#jXlxVHYEB     400     120�W��y3���Zl�ٶf�$5�����Y4��21p�'0l͟oА<.y����x��(��Հ2B���O��)�*�!!�fkB`wb R��e:I�{���`ϭ#�?$���T�J��1{�+�3)ټxX	]��^���zga�9X>�U1#�%=Q�I2h_��>�5.�!����$MĬ|ܑ4��wײ��Ӱ �P@���ɠ�Kxt�7�K-O?mv�it�c;\�|�+L�*�\+���D +�^$��T-/���mK�9wb���u7��@��!&�9�U"�XlxVHYEB     400     150�&Л?gq�P�f��o�j̓������ ����.�=V7�ç(i��]����O	����9�3�L|_�$�(�[cq��<�=AJ���N8����H���0:,[]�(�ڏʾXğ��(ۿ�Y�	(���'�5���_���:W���ƇQN�5|2�PNҫ��nv�R0K w�D�;׺�ڀ��8�����/�T��~��^ �����nrp ��ܳ(�Y5��a���E1j:�&��XW�s��6�s�jo�]c!�/�>����St�l�����/����m��N%��2�}��� ���z��;+��vߟti95�X8��S<B��O9BƥXlxVHYEB     400     150wq]�:�i)�gO�X���O>��G&�N����Z2M,[ ����p�:����7׮��+�J��n ������L��#��$���1>����f-��7�Ŝ#��X@�ő����@��5`����8篺f�]��bcF�P�d�x5�@��$3�hBͲOˎS���F�Vռn�wkē��ݒ
1�T����e����犔�̱�%�Iˆ1���i�=
����7dP���j����jȉ��}�ޜŊ�y�@�,�5���ڶ0�lH��� X��1Đ����H�d����`�SP.�,f�XT e�`��,;�ż<�
v���֚�n�����XlxVHYEB     400      c0Fq�% !A��b�"[�5]¬\�u]վ8�A��-7�u,r�܎{IVbs9.�-�q�^�9(��a�w˲%d0�l�D�7�+�ѣ�\{�U�w�7�Z���9���
��w2 �)T���m��ń-�@�G�#��MJ���Xf�T��;,���ڂ5��b��?D��%�!�[n�h_�;�Q%�s����ϖ,O'�XlxVHYEB     400      c0g�!g�e-|�ZR~`T��A/�j�`�7�l0��h�DDnSb�^���=���v�{�k��z�Xtי���N<���|@�m��9��6����*��H^}��V��YJ�� A]��z9#^[��]Iӕ�/�6<��sY6�wY�Jx��5�%`	 ��� �(�/u\��#K�_l�-+�&�p�&ʡ��6
��XlxVHYEB     400     130B4������ji2�C[���Ti^p�n��nM�nM���Z$��yTH����h�Υ%]0��?��ߟ��kO<M]�H��U3pU%�4ɟ���!B6��G��@��PKg��o�P�7	����5��/�(��;���C��0�[��b���5�!ҹ&a�"��cI��	'�4^���V�001Aw͡*�n&��?����MǺ]zZ�`�%����Ek)���4�3�1�� *�:�4J��k 3�&R^�qUL��=�ɽL
���y�C�p~��e���d��^݄��`��8VXlxVHYEB     400     120�$�mf��$��N^���ny�P��ܯe�������v�.Щ�� ��~~fosH勠�@� ���Eʃ/�PU�����Ƣ�B �Y�C� ��AA{K����dxQ�C���Qb+9�3�¹���ϲ,��`��X�x�D\�^Յ\��z�h�Y�!<��1��������I����R6R�=�j�Ir�D�X+� |�ߕ�����?4�?��Q��5?(y�����}� A<�NWO���|�	ԝ�̵�	�ؓ�I<.+1��l�k2ּ���������l�;Q>XlxVHYEB     400     100�;8���.(f���e3��o`~э�K�tJt����w�M@@�B�}�3�����h��z�p�J���˒�(��&A�R ��kjܫpؒ�eP� ��aJZ�0C�u�k0s�e*a��/�_�9��������x�GG�!EdN��1DU&�J������7�~�B��MthR�,�@����v��U	}wT�1[�U8�+tH(tp-�c���ЦkXe�p�$�ӵ<��xޛ�#�/B�L+�J����}��#UXlxVHYEB     400     160>��d��v.���(�����<4�guA*
3�v��aT��B�э��$8��&����ꖮ�/���?]K��}�K-����|AR�PerJ�ee�(R��ä� �/�b�WR���x
N�%f��1$qdz��5����?5=�jHJ��F�jf#��e^��娉X��
+T��蝎��+Qf8�y�t`;��4�3��WN|K����gW�k�ع�o]�|��SU"���,�����̧
Z�x�>Kq�_�Y��͵̮\F�(�{7�`�Z�qZY���_		Y���
�k�M�U8+������[�i<�� ����c��W�t7����($�s#lP�$<�n�{Ce^t����jZ�#XlxVHYEB     400     1c0������L1 �>��g��÷g`���.�N�G�b��&o�i&Y�p*O
�]`$Nir6���Ց��ZiTN�}X�8}iJ����O��V�x)B�k�}�C6ꓫm7�����R�3E��U��Hl%d݋b�m\����ܜJ2��S��s�
l!G��FS�l0���_$ϋ�0�&&���'.ux�}]4'��b���qI���& M�MT��TW��ó��q�t��o�b����nB���=}�6$C�a�7t��i��!�y�L������ԯ���Xǲ��j�A��]�)h
�:��Y���+U	踁ZA4*�<��HF(���w��0%b�z�<�B�� �{�^�a�b�<�t��˒K�-��أ�jo�}�������U��{�Sz�F�e��Y\��%��7`��p�~����V<�$^~�������񨞎ދ��2��LXlxVHYEB     400     1d0m�vv���Z:pD9V�&�!>.��T�i�����Ӏ�#�0���l��Ay�%��>'=0���|�.;C�+ �t!�XS��ט����zIP�ع��?6�VD�t fX �]���{��SFd̽��[�f�Â��B���+�y.��Iǚ�(�� ����ϰSfͽz� Yiߚ��W&l�ˣI�t�����:�g��B�0���	>�B�4|`U��s��2gl�l5gm#ůn��� �[D�	�<����%#x�5���_Ok7oۋA�..�W�ۈ�K$v��2�ǿC��7�F5�xq�dm@:j#��QAij�;d�2G�����V+��X}8hs��T��W�+aS�ا=o~��?[�x����qg=Sԑt:K�'��X:����BN�w��7e7�P�] 2%X�m�(t��%��e�'��Ys(��qK���~��H�,�� ���L5W3[�&���Ẫ�4��XlxVHYEB     400     1b0��������;�{9��$Fa S��"#�'�!��v�3��GI�~3�bA8pۉ^�)tr��e��Ԓ�~��eVt&!�d��q]�0�ʂFs]�oL];��˸ˏ�㽠��,���:�l�0s�_�g�s��#�8�{�����͔J��jh/�+�����S�	pK{v��,�%3�#�wj{3`_c-����W[n����=t�����D
��7f4��|���L�Q��!�H��>���V��I��+V��ǚ��u��!ZʤV�Ģ�B�y+�U��1�{j�j���Bi��b�3qde���C	�:�\�2�(������Kر�5� lNęI�y	�h�@*�(�i����JV�7*>���"^����������b���0��m�����8y̩rU*��ܚ.�n:*2i^���y�6XlxVHYEB     400     1a0;��"K����b�L<t���:v5���̎��4�HY9q4�+%#�1ПAx0r7���4���g&�(���,����1�gr���vn�(�"Bn�K�`:i���F�)+��ݫ�׉�����mp���l�)Ga^���L�T�^�u��e4�e,�zaC�/�@4ē�*�����9���Ž���/j�zR]+�^�U~��+�ayP�۫yGr]��|dJ���2)R�0��Ў�STM�_b����/���iOʤ`��$��ր�[���|-����?�n�%9k��B9�䴺?�CNΖ@������9Xm*�Js��ab9�$�T�m���}������+ωZU��Ζ5�⏆-z���q1�d�N1���l�M���"�i��}��l<z�Pl<���"���d��m=����n�XlxVHYEB     400     160�^Sİ�2��a��b�ؑU���pL�þ3T�p��AB��1������I%�!`Z#OX�_\���;\�>�$|��	��L��Kduz�_��8��*��/-G���]4�{���Aa��N����hk���d3QO�Z`Z�WVb�L	bUj����N9٭Q_�h���oᵴ�W]�k�Ԗ�ۍ
'�T���Q$���~��+���>9']�4�#�����KM"����9��`�_����{Lic�����:" ްb�f��ͅ�.V�{�_���>/�"�c/��h2���0*�e�$�h�J�_t�_����=�Yja<5�A�2׀���Y�(��������m����92XlxVHYEB     400     160P�s oS-�}Ec���6���x�u��v�]0�]�R���9K�o�U_ ^|7$H�R���1��dی���T��k��+���Sx$�/I�4����dL:��Nla!!De�E���I�GW??�vF�iW
�r�NJ��g�� rԚ�t��VD�S��'[7\��`A�x�	��\��+~��n����iS���ޑ��XP9�g��#�!��®-�Ε\2Ķ���v�iRFj�oDh�S4F���Ir�,4z��m=��f���<<��IB�chc 
W��9
gV5�YH��t#�J���A���M�R�0�l,t�A�	�M&n�\.���3&���Oaz8XlxVHYEB     400     180x�~k�[vX��]�L�CG@Z
�!u�*]��
nF��ͅ���w@t,D9od\F�N۲�CCܐ j�  ]��_b"�Dd�a�`4���5u�؍�/E����s�?yR��5���q��j�0�x�;~CY��ޛ���~��_��H�u����V�9�MZ�����r%&A�vH����<um�ls�n�2��W����������e�B�ۢ��/S�^�P.yY8̓���05U��T�u�l�0FTv|?*<Az����s����[���Sg-,Zf	F�J-;���o�L4k��\���}�FD<�ԁ%�����.�2*�Ҿ%̣�{[��U'G��5V�]��6���L ���AÅ���.�AL��tp���F[�!���1�XlxVHYEB     2ed     130�܎9~>IɗKfOĹ�Äh��v���5W��F���<�]F%��#�
Z_atů}~�Mթ�3b$�o�Ψ�`�T^�XU�k/���|y��+��l�{��a�7��-6��>~raA����Θ�kW?xN�?'r�p�M�Y��9�{��>箱�3Q,mw��&��wy#��x����Q��͍�:ħ_q�3{mtR"O��?b-(��Nܓg���	��i�'W��`c��w�+��]~|��I/+����
�W���W<2+y�⸣�%�G+J�>|�]�?%s Eޑ��36[f��ۧ=�u�>�@"�