`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17984)
`protect data_block
s1PSxzy+lgypEb8bR31/BwJeoEHGfHH/SPkO+OTO4OzfsjL7MqfAGbTamlhV30ohl9wr+A3wYn+2
lzZrdAOGxYO00/etZrTpWrJwiGPAGREnnxErPAVL0vGMFL+GFJQiAPadhEJkRMQKHzXzXtuRDZzp
4rpksXmcTqIKPTjS/eukfP70AxnzHwSN7sxzi25Bihf5LXIwX/F4oK+APVDfnWXoNcZSqUzz46Ke
de1MAWhx9Y49OOb63YvI7/PIfceKMMS/7bAEKiRS50ah32zy9lI2GM5zFSA+uqcV+pfymRNtd+G4
8OTClO4klKa1pcrX7YPfyCezphJ9cCKB5u2hcK2qGqS51EVGcfTJvSiCGHowcb80/a8EnTtYI+PD
MuupeqZj8Ueg6Qv5ioaqz08BrQTRKhuF1JN9fVFUz6v3W2/XZFWbLen8S8Z9KQC3WEFiPCPRP3MP
WytyLAWJ8VefVjkZDWZ3nt95qBiwjsgPTx45tgs3Ug5ZUoM2lUVlt26M/e9bj/7GsisVkzpogjrT
4n8/JMJmLfb8nroF8ntlFltLUWmWT82BkOGzzAXzzVPjWpPPGoWniyzJcxvnUFRU8M0w4Co4lw36
JQ+qxEOAZVQL7z+Q5b11T972HBC3tCB6Vwr7wL8QD1nfESPuxau43w5m+n/vFOjq5D596TNPGE8z
hmlSmRTFV5wz3GuagTUyZuQEVImW7qV/T0tR+GKyepjQuIn7Y46C3omN1WRwHwX/aiTQOvtS0Vvr
wIvd859LG4CD/QeS03VHM5xuurRZM2zz7eNV6FAus55SXKlyGaR9xTirDZj8RbD6UO8k15aSu2aQ
qen0C6blV5TqStWerUr7M29Z1NUf+VeLitTtuXdmG916M7pUvQlyY7nR6ZzkaWgc09CQpHqT+eWj
tcPYXHMcWTaNqoOlyRmyNjCs5JLVh+viZy8PPXaHQTORy4CavFwtdX6//grqCH3Y+/fahXQoVt9o
pcmq4+7iOuP3uei7O7rYQ4quBcXxGFwOmBAs6+igUoJJ5g/q9pDKICNYkGPRcleR1t8Ce5DNmMJr
GeEpN6dDIkZ+ZfzRkpQmwnpvLaFbIYl+O6qq+vwLlKfPwYsIh0tGzPqtJK7I6e/60kMuj92K4BXP
mHA2O9oapek4vge+xB2P2A0FcrjrQFLfU2YcdcAfIdv5u03qi4HN+XTrGFHSrAP8yONvIr2VrevH
sheuL0NffuBZ9FKZYKrCDx6vg+Wk7gK1I2mLzcHX56S8NM76sNs8kU8llodrEZUHFuVi2aQiGoM2
ltJ+Yf5Glk+9gaoMbtmvWoC4JbHJ9ymrdfBGPSitu++ncHo2zxisdiUS3FZBw14lsuKwIDEJS+A5
Yzuvr9YjiR90I51xC6UIztZNeL39iRY0iOvB0TFY2FMopsCq/3NpQHgbJCoaMnKBbo8j0cUPUBv1
9T9AsqPPOXF7DLMnb0hCGDYd0rH2xdUlOWag5FF3EZPMyNdzDDMoW7PxwGwOL93xZo3MwAoGBNDP
83y2G8KqqBbfDxzSl7i26A93eEds791GPIT6lewTLm7KG5U7BbEPHu89bpeadAjjfBUq+ADh+z4l
4yvd3j+5VuDU7tVpngudjaoLVnGWPF1cRYty2c1Q2P6pFCSDOgqREx78FRjz9uxJAlU5w33bUXNe
E0BnN+HaAeZOAWe1s3PZ3w33rInqoyq/gymih+UJ6GLerbz328LLagZywNIzFiivahNd09NAJTJY
vFqv2UsokpqGqwULSpCFjDszraCnUPqzkdTfQxj6xSc5ah4HahDdS+vXZ7xQ7ytWZJEIkKV6r391
w5Yd8E+bMhuoTbFWnQGfroeehu6rT8bX3Ct3VlBsnEd2GUYFtG7/Q2mzi2O99FcaC7cK0HAbvoAI
CLUygvd8HvIqJi+23M20STbVnegNnp8t8YkpPH6z2yzB9pV17VI6ImcIlp4b7UOsRzo827xT1y/Y
DzNdoXwtI5Y84l4R0xuu7Rj6e0by7ElqQBlla38RVEG/F/98xjJAForzI54G8iIVrC/2EdRuVFRY
la+LIbJM9UK5RjaiuaxX4IbuKtm9RjPGs/YCX2fVmX/6seLadM8Ohkj7LLtbFhPmVbYA4DqdqyHb
A17s8lYWL6oD+km1p7FajUbBwJmXSo/KRUoRaL2oNV1ECW9hJI82jikPLtSjiuy48uSICzGvtU4s
6Jsi77cmOER4Xau8dQnjx18o88Y/JHLohZ501jfRC0g0S0neX7H8rJcSKW9ZMJg2dMeTt2m3KlGU
ge5pVu/P41dXBNh3mbMIoeGopTXKPBXcgx76Dxx+hAxSGq5px3riGxwhbA/JIQK7PYq1kMNZeQF1
DDYplN4TK8At61nSdo6c8Y8aHIwg7O6GiurIZ7A92mB0OZf40/sxAiGywJX85ad0JCfAL81xSHBi
bVrbx3VmbHb8VoDPjYPM5dlb/aj31cC2Ehq6672ii1HPG0DZeG7OnMVgCYFM2guDvYXG64ocZXo7
WyGErOurov/vvHCw/XDoENGaxUYUdztHV3/F/nxgJgjYThyRS6++hvr8NswveZKdBOKLUvQzRpg2
ud4malIbsRub7NPIkbnfypQPpC1ljHLvcSX7SmIuYrQGnqatIXIOQfoGsxeaXSMwyNK9YIxF4ou/
co5WzU1lc2YYMflfNRxctsa+otvVKwV6zq3NkFYTDLzI1iMYpxeIGMZiETlbO2xN0ee671QpteWy
HCX48VgM0ZdKL4yXYzgrRFgvEGrIqAd1CMSAAHgyybnhw4dIoFgULNXZiIYWOutH5Z5649VmRxrw
VibwerG3F5ZFA9K1P6HN4p0137USF//sBZ9E1noMfN2r4hIvIxxCchWrRxm+oTqbLF+iCdbs0gXd
rq9xTVN+CXs9CzdRhTwfJiHs3yp9V49dMJ0CLziRdvrE887EIMDIs9o0h45KZj0RtHb6j6nrHZfq
x9XGm/fJ4rHAnvCt4N2pC8OdtkAlbvXYhnn47G+cftKl/Ed6swkXyNTEqq/umJytzEvHZnleGEzz
hpUgcMjKDUilSt72OcMhfAJoXY5YrjjrnKyY9rO8LK5FEaVg5CLDQGNxT3Zp0HSrdEu7Zt7qUMfm
bgB7zBEZBn5guJVKQqvkumPEoSOa5y80NTgwBNHdeNpm08oDmH7mULrhkAOc1U+80L3/R1AFoJZx
JSE9//LCDlVOOxX2RorLtybr9Bjf0IC07q20s1QI6swzY8QOsBOPtz/xavhxi1XvcBI6b8yZhyUA
oGtbL2+yH/1mqJxw8YQQK/v9X+8k4d67KCFerc/mbXxi/b+s5BxGT8QmQb2I+FgVAaouw0cJOlCd
Xmk9od6Wm9XEthRjQEZsYtUYDfwrfiV52inFbSwpNxFgSDMfQ4kZe/O7OBOMUAkUFpQ2bKzkp+kJ
toJ9yDbHtnMPnrUZ7ymKtLNTKl1omSnDr4zef/h/H52LKTJSWttrCBE3cGDICsbmVNTrYNVs+8P0
/6UEed8LSaMwWEPf/+IKYnEuWFCdgSD88XXyzejEUUTi65WR8WSFrFHSvzHf8o6I6EHKf4aY/u1G
6Qn4/gR3pUCUiJhgPKU644xeof6SoEjw7YoYuLh5hKufgqs4avM9f2ayAu3Of+iApd7T/OryJj6/
kMDeJB8RaqalZkJZqZhVj5amp4enzLc/vxqnZD4ow8S2MR8xR0zqyHJCOU1SFqnglX+/Av14IG7r
btfEyEpSGwMWnFqGrQ5eLppTfq69d1E8uEcj+/+ztXEtVYLsNB+iHXvNnmyT33cqgj52cRDdp/BO
5t2QJU3AjOSdS9vahaaHr5DvVFMpdP9xjkR1TNOjAuZuERYPm2wVGibnq5ebcU/avcgoeAkjsgdQ
SoPsML+6jzmOKNI5SO2C8wqlHHZazmLgIRWDb1R5uqc+WYiUGXi45q+2e3q3mTeHfPLsDS0zU8Au
jPCEaOIpvnVwM6oE1m/0FDmyZ/RWKi+7c1dkzW77/+FViVlO/flz1EApQG4WKuQrhUcnAvXP3tQZ
tgZns1lJzK8+UNRS5eVD9zXn3kjXVcbOQ6XCwWQDg9iHTDfNmgZ71s7+XVAW6E4bODyRwWa/ZSth
egDjmwqVWmJdqRDxA8vWGN6nMNq2TmGVmHG3S1GMpE5H52bwnFr0JpoAm5Ao8fXi/TCw6bj8YFAc
Vvu4mwYhJoxawxeZc4+N36dBmAAh16qZ+DIm7+soxh1Dd6nf2h3d39eaP6mY2NpSy3lCLrJgDEcT
3C7Qh02jvowqSAFsqZfXXYTbTvsk4MWSlqHNyy0tJwkRYa/f1XotljxQ79lD93epAGe9EuSd8LE4
81trPcTGGX8nzHnGptMdYCYVlCt3hMMHOshEWtpdlxaG2LJOWMx8WTtF9H5FyrRpMpJ8HAKFWFn+
3KxDZ3C3HiJxmICCmprRUA1VTyw12TUG/qLNQngrtw+HpsIvJaV58HThJeDSNBVBZzac/erCC515
7JkfJKMWCxwefdsPQmclP4jFgFX1G5dWvZQGYSvB5Jzj48I+6vt6wl7fe76kiuzR8FZCUeHLr9lj
EkD7BIi6gfYEikdId4W0u1RSjn7s38kDKI22GKhQSfmIao9JlgXAxfFOOOH0g37snIcapWUoZIEe
4KQSw64zBsv6XLhIzZmUko6YLcSmsxN15PHs0AnNoCr2V4SyIew810F/YGk0L0TM+TrQp+k9J/aB
epC2Y+GwChy3n/1gZQfQXT5WJ+oV/jLG4D2jh9equCLg5GaWzMUiy6lBU1Pc3kYWgio3UUYUf7Q/
FtxgfWCsv9YLLAZH1WGICR9ag0JG3DfGwK5pHLs1FHhQ6EV7al45mZS9WYhjcIQ5BzEBlXJqlZWL
LrVuYnKdTadzuXtDEs4X3EW1gLIGJl6NbyLpFZBG23uTE9sNk1QOA9QemllS097YZQItv9UqEFvf
roEQbk+egktrU51nuKPsq/lhGVvFdNOJBR12J3E34V9vd71kjmWAvP/15Dvi+hNhDsqSc5SY7ZjC
CzzoENavTCZzN921OracOplewfqQCsg2sMM5vzK6KIvXiQYMRpoThEZ7h5/553XAnilmhvWcjMHd
AL3BwUkWeaaJVR7dgL/x254POCNhsgcFGCIPpraK6KbBmnIVBNmabPHb+7K38wPXfVX9ggveLRca
fre/5HfpJ88MkDzJkGufXGi2Za8R0h/MI+GlFwI44dsJJRLP8z3fXf7v/42aAbO+hccEIkSLxvxA
VranfqWgvsaN7DrqDbcxgM1gJOHYMdsX5RpfKiFfxnKEx40WFgeHcR4tAciYjrNtMgslvelcCanx
Z72tLR4H96NP0r4v2OZr6kFbwNAMI3O2xhuDtS31wwfn8VzGXLTtfj3iZMkTpS7BusTGCPWKe+8R
nXKtpb1Z0jlTDG9GCkbV0akzkW/C2NFWIkASlRA0KVdfwCf587S2ociF7jzutFaF3GJty8IkxAfj
HMDqUVKLVU3K8aNAZpJZQ8+B4GU5ZSXL6EWXF/RyIFP6hcls8ori9KbcvvbhanV8K9LfqoXsPSty
dJWF26x4croiZ3J95Vo1e/dTfJ8ePlWDT0dW9crpxDqhdB8LVYctCBnPm7xOhT6Ezhs/rwwAk1GM
eDHxY6/RwZ+dOw6Ajw+hdwcwTrqvv5EORgczQrUhk9xjNH471BvY7SGcZaiGA0QIR56VmjjVG8Nq
S19/YlhtV718GFDOuX5k8Q6YoH++f4ckGMDNyKTbeOowEuzat5aMRzp6tytk5cRLJ6/OcknZ1xiv
HoSDZP3tGy+d67oNSB8lvGn/EAqAk1uuTMG3hcFNqqDn/HRraGOIlTl6Xcq6XM/L8j4B4GzmEbsc
Wc9oOF7fqrTWVAN6WDLGNrJe5E1Qd8kfDEv2zKDWelR7M0hldhCv6DOYHPdcVjjUJcCYptEO6kcq
/4wLmCgTSdoxCtO07I8rvhPkbX++O4ukIR0L6uITTCwIpMfFeTU7DS6gLGfRZXpCz3oyhmXcMA2U
IrRboOq9/yqFU4sKC/OspY/wv/kxP12wXU+CK5Vuf2AZkEDmkcxYZ0lebt88HGE5rVvTzoYB5Ud8
8lRwFx1TywX9LCXQpHXMCtDqO7iQUzXl6zwJdgt6+3gz0TiTpPxiuDQGm+OV1fwwkF1FbnsWDJ9b
9P+M24ocfJLT43MNE4LqflDAijS0arPLB0iWO9lkA1ewP9UEB8Df/xUPqoyBSD7p1PsAepnubRQK
Q3dzuBjkJc8mZVN03FGb3sAncxksp/e7WIIRYJBKgF8f8qkvkh9sRTueSTizZW+yrnmVm1kEwssr
0xpD+xnx1f4N3Hg+NjEMx6kOtNGZf0izyyzwCyh4znrX7vz78YkDSKLGcLnO+EabI+Rxkl5EapMD
Ie96Y5S9DInsRE5OYPLsqQ6Jq5LqV0KhyE9MUwYz7AA4mXWPg3QxgLkYYQ0+N/yLcRHs2y1i6Bwa
S06MRTQvKWpJ/mzsYCGDslSXBia6AVod+UeKwMiy0VfrVtSgL9RpRuVI6Q6/piPV5QS+3OboqK09
F+L6YDzzRsgNG6PUe3bNaC20+aBD6vC8Rei0D1xovkmVn3/eoPjGhQhwOIcG8wFHGuCm7E6nX9HY
iJiRRToAhk64KiKbypmeUysjO8WBq4KG/PvmtAeWHeWRf6T3t4Sw3IS3c/4n+8ezsvskBrWJgOKy
C/xX3Vr+jO8ygc4JP8uCui9ygvUgwmUHOadimqyWGlC3XPXJILBLN51nIk/XMn+dz0XKNqbArHgd
bVp8f0SEo0+3UAlERs28mlJAwClGJoZeKLMxFHs/6zwHGZclyZ4cTXVFMEZaZdvfp/4kST1VM7Sc
pPGcHdE588Wg1IvoiVP7mGaAGC4oScbj6SOfoGJRhGJFnIrmNGpkmXIbqW89EYWugus+6fi5WSFM
0llFpW19B4+DdnYfutYf9NlnmOgfWVWATHF+eiFroSTJcwSrdr+DanlU+BCretkt+0W44AncGkh/
Jn52j6t6IPVepKHRtHTotUCyAKVl820dqQLi61Kxx6WeXCy7M0zYWJJ+6hAzmQF5pRymijEvRzp2
1h68p2rPQR3EfE04n8i9p+Js7A7jUsgwK61xLnk7zkZ64fIovPk77OHL3ciVjw5XAO14i9fL9KeG
tCTWHgOl+MkZ1AHS+2BXsHIMaK+0MKvCVRuCyPTJyFyMKY5YotJmsST1+iHTI3YbIcumiYHYTOhG
s10E44Gzx3HsoC+S2eNA0ribVbPjULu8ngS1wBAspoXyVqLORppy6VAZnxc99QRJEl9yCKEB2GVX
/1bozfbW5eXkl8GUYjbVFc5jZKeJdOTuyFqXw1Tt4mSCBbhvpPiltlSUMRCWrBmpyjeLd80WMyWN
2E1Ff5LAALKKu+H+GrIUGZvumuTqwKiRwZtCt7azecCz0Vr0+ENNJR377VZhcdzlzuzd7fDeyiHN
MUc0NZXabW10M1ffdrpf5kwXMwKq1Or3oOgp9JeI2j92kXuGWDeJSYfEqExl4eOCPi3tIdLQQTBd
U4Ok4kfCpZP9vko6wH159NmpCowlE3YzTOESA1N7JlrBAV92ChEoVHJkeIwYCVE/jb34vxAtUntY
Bc4ReZlwBFIhO9e1xCzCvEBiteh+YOqHzHVgj/DmXZRluvTWCkVIcOeoQ60uaPDSoKtQ05hzQ5N7
aJt/pZGTSU9+8YufKg1Kp12NnOlhd7gFFD8GkCP8vypbsXHBFdiZpPY6SvEDSxcnEfyKOkcKTJ5p
d4WzXcM0aYOAU6/D9JeyfDzSYKBAEoQJApCMX3spVlZgntNKSlufpYP0PY4VE7auer/y3r/AbpWt
IrpLRDPSOS7WDsx2qpn0XW8Wolp8PXq4xZvyT/20a+m4p6adLmvp7DULSqA3g3AcZnEWwOHdHbpz
JkDCKX2U5wDvcv5XpI7Xdl02kQXVpJBE8c9gvB+xuHOLV7FZ34ccK45wrsgC8E8mvRRaGpo/26hq
ue3XquK5KBicguk2VY/iWDKg2BCd6+nXderGSITK7ThwmWIFnUjMdf2yIKkvbf4OSzHeX8oyZwVZ
zTS5q8qYLD6+YuFkN1j8Zwm1jEgAiiDSbiyJpWQpUzEVcASeUjIqalah4EZrg8VslfXYoAdUP2UG
21RNOxebhelPrWZgO6qOMSI5REk8uz/5EizYFIRGBrHZhULBkFmC2Bcf32UY76QHO24q0/gEkvFs
1LyyPGGf/t5WqVmBowi3onxJm/eJQlkDu32AGMxZ9aeW+LcBPG49rC/YntlaCUGie+a0oaY8FJ/C
zg9/rZv84SMkszbyHbLtDbFD5GhzTeazRI2puqTAg7Z0xk2L/adi5qvgSbLkMBzRxbjr9vF+VWXy
v0LS1pVNLCWK/t9J8gd/NIUtBTY17HYR8bHr8gSwpYJIhpcy66PX2m3qaZ3rLAhEcqNY2NgkyEw4
QpV+6D92bWCB21zR59Irzo5SCw2E9y1CUf3ucN4YasgGbH5rdtxRLTOCMibh2CfJDfLytLvdOwbB
mU2RjgDx/OhkJpkzb6BCgLS32oW4E843/0ddnxbDmy/DFcCckZuKtoGJdJZfoiydYvLp8UT9igKx
ScU2FXiIIJOWYftz0AFr6nnZhBhqSvLuKIgsJ/JAuhQA0ZTOy6jP1iXNodficvvtW43vYS33SX2p
1KGGgBqnDg3HTCZT8M5OgyTieiBCWRJK1052gkm6CUYY8gxNNDexUiVw31oRCEggu5H02IFEbP2s
cJ9EIVUM4kCoyeNGTqjBw/UtgNW3NfzA2BrQuXvhVLGwnM0o+Cj8UjxkAqfO9O6+l7sSKagVXEbC
93Vi8BULoPfF8/xGwUTe2YFLdkon3yGlECoao+3+Mtq9GIy6UCebXGWliWIhiLGOOvWElMvstHd7
nsxlbjmL2O/iyphCZYSGqxJIrhMRP4ZNe6I+4Js7zNRJDUNXurdBM3KDCqzMjSlhNuUx5VdXKIFX
h8veSKFeOqQ7yPF9rKgSmerbtU9IriHk9l2rQEYC+qIrp0IZBhwvFhCALsY6ZjggXYAHSeX0OHhW
Trt0tyY+pxr3vRTd6qnv1sKlnyZuae8sNWu+69HSAtOiSG/vGEx0IDOq05WeifCVHhl2z4467CI4
hnxihQtgdNAS/nZbNZIDORulk2xJqdWNtG+SbIeaNoBPEpl8vy/0GueFtkdYA/hajtuJ5QGfeOZk
M5tMk+b0MnAs8jyfkAlfZrSBofmKY65cRENxwiy8OFraDbb2i1N3/ZI90TbDkFZPazywfNJhpOR+
CrppH2XhpqWAT2uPRrRRr1Lb8sFyu2MEIBTowa//P85ArOPm35F8BT0QL6OSkn7EM153B/CCQis/
QEMA4fU/xkpEQ2tgNJYP4+rV1AuQvfiS4UvTebmoakzpQSU2Xf62rV83Z55g5d6KGUZ2075R5M+g
qUSxOe9kjWsRUTtPWscC1+d/sizYDWSrGWoYsd3jy7iMb85MPF9CC8xkTxL/ymk2qSfzA3ul32fK
B+yzZDjVm3Fr63WRQapJLNY/Y0pp53uc8/x7piPk93uxlBAnxVA1naO6/LNT0x17bDsBJEmWJyuS
9lGDIFxnFKaIMX5/zY6lgw+1GvVqJ+gtzv5WegLG34wEZJxMrU1nlvE2o5CJZHvpvXSGLOSuHkqg
KjXZlSLC8tWMpA0Harv0l9ik6H+VIwobb/Vra+RSfiF0Km6ST93/9FttLN2oxH7J9AmvVNZAfr1n
6E/zP/wQwlUbI6e6Fo3RK2tttXULEB2ST4lI57tMrW9iZPxZ7xTXDEYjJhIorMONW1WvHjLQOoaA
fGB/IlcwNqnJ6h/5vxY4i3WeAQMjpz/puptVY0HgNeFnu1SgZHYnesgbI7Q9Xt6ZpouxZXQZ2kB+
hLDj8I+fWjuwPwy8/LwUzVFLxkImy/sPDrAmU+hmKPLx5mMJBLWom1Bh7ZFKqnVWXtY3e2cbpI2y
mW4BGoHrk6/RABYROWU/39hwzLv7FiQ/dIkKw83gXNoox0VQ7MgxX1gmnHmuIraxiM0uTIfPB1Oz
nza0AVzl3PeTl6GosYnCP+4ta8y6inwW5YDZGwKTOn7XYyqLSLR7xNhxh5qLTr2Kpy/Eoy+gNfrx
0W5LpKjI0FjSuT70pYqlfZqm84aTtAZJYQFdknlak+Bhz60uHHYWiOvwr0R2aPy96jDlqITVBFCr
MSYk6BEDKf7QDgZb4nEpPj6iYtUDngxozlmWXt+Q9L08slCUFyZCDWIE+Tke7ouVtFRsn/BELLT3
cGb1SHj3KnLvlNJF4wZ84PcYidkRFosvyLMFI/agFAGuVoSwIj0mmqxTZVuz0EPsduQ0A83J4ATL
5CnMF+gsV1PjyR0HmBd36zYRRXuhWnZqjF0qWju5cQE/yrduEcyDRdPV3o51VMQeCoQMAR2mWLvF
Ei2d7PUW1hpZcTT05bIyZ5sjeJ+1+iCUj4ujstQoKpK5/9EZfNPztPiaB68ui2WYKHbzjss17as0
p+OKDoHHfmWiTy4PMeSNB+rElrOggR3ixD9nHd/lSpH7csexgIIWIX6YkotIOZT+GF6oTt0obDdN
3qhJh9l5tkDYv02u+8lqljspK7OW6FtOqukBh5NLb46cwCEJqk8plJP36WpfLn+X59V6Z3QNHTyb
lDIAxQ4hTOPqVVWG2WNZmmrESjpnWJkrrQYtdLLLq0FQmfd0MaZpshmbQzL9LStRf8/iRMWOB06M
CoGgsfcHpoU8RNPg9Im4nUz501rSmwXINmFiJieKvTqEwnVmg8JYjNn1fXBnnYfoLrEWZbs3rLNB
PMBQYf/BWXf1O8laqDMH2tCfSzhNizMOLZ1xVar4y1HJ+MrhIGur6XtoaUn6oMlv9b+E0bvSZsjN
cMBb3/pTlJITXn5KTOhFsgFrUFgmCNRnVyWIC+F8pQ5Ohez2d5Ns1LangBQjDBC1dLn7iczhrfVr
nb53WEz2ONeJjJMEIzTj+GV5G9e04jVS5DPElM2dDiofE6vHyaH0fC1d+tz1TuRK7VdNx8zjzxTU
37A6hI9T7E4fH0OYjCdsHM/VEJBpaaJox/zt6wdPwfG3jrZosUsszHTcUsSI7an0o//VYpa8ao8O
83Rva/Tb05EyQXy5CtJi6Kes0R741Mpf1risftU59mD1XlM7JWA/s38EP/MajhA5FbR2wbZqnJ8e
GO07raC1gABtE6SqUocaADZgwc8W3D+m+/Yvuo/VW69K4DsujtkWY7OBT2ReRNdNDnDBU2Drwest
LTX5qMTpTVHym9fi8Hrv7yQWiWmf28owpLZVLOLfYDtRPjT/k6I5IYut58chh/erdTH9SUQfDGQW
OFvShmir+Qto/0n25Y3Js+mQspDX8BOSd7vDEdB6h4UE9l8AHuB/qRfQGP5Ga+Hs5mEhNWGXatJF
VZbjwHYzIQHbT4uSU4VpW+JH92oiNtp4fkuwURRyjAJgErhMnoWGoa6Hhi7aYrAGCNMkSL3FtmPP
645EgiRAWsUkDkh9hW4rcvPMZHJa/+io5ABquKljUg0pTHd+ZjoDwGEskqzGOWfN4KU8C5tEW3MZ
yAE5f+UnNX4RZgIZi1zZdfd9vqCG6LCP9tmAxjR8yY7t6C/jFLsj3mdSJso6cfbjpdtPTwBrdeqe
nTRQ1tE/LE9ArzcL0KSMiZ+LiSqWxEQhAdh9B9yLrgU0uRtn8XAPBk1bZO18ZESKI6pmlS0WRqds
ZmeMpH2E0Fx6NyEYBO69DHp4E7e67Qs+sYg+AftkJFujSDH6aYVyLzsinXxJZ6DIOyp4adlXvDNS
zj8wg2QpU+pOmcGRe/m7MzXZp0gqVuwakkchCYxLxr7EXrOuNjYLIiM5LmOAHkuXofMtpuF9eA6Y
QnigC35dNqEfguXm9fmR3T57Iv5lRd+VWZ8PuTsPbpCrtWYDyw0Lkqqq3xfjTl4r5rO+OBVw6LPs
4PCCDztLmtvTUq9KGoUWESuZvM6HSg/Om51opm6ubvpLQq6JeYlqE10WEgP0e8E9YxJ92PUjo8Rc
FnD3UtG37F2ezkDwjHFDFHZL+aEuaGVvGr7JP5flfnJUmgQryZdHaH9GoAeGbthMOBwObSm9OhVN
Wr2ReAu/8bJbqxSfkHFFIVIpbwLdsT2awOILtGKM7oZngUzfGCydvshdf6Fifw1ZI79vgSyfMtgB
uACH0KzKxA4th8XEVepNSf47lquzTUIF5ca5hwHzQc2K8iRt2oBMw55igTLm+vMmez7u7WavtjUS
zGxAut+VZE2tQfyBI2zJCFdAfuqdKiqOTeG+805mtA774r48eaWWTlphkJElCW0oEBdgzyIB4ObF
D35TRk2rMHFU8f72LukkM8nLxm4eoTazgnsvhxDA/8ypqpi/wc8fZSM7++RSl+11+LZW6DexhNp2
dqnXW8F38HIdVici5xEkV4t8eE8mOpEz7Vkm9NcfR2t65OeO4eC2PtOc2e0aELxsaIYYGvqOQxYZ
dsqJEVxh7wAHI1DDmS2JuH8y104WcBNbf0xHUdcHKnQRls7lhuFsy6u/UHnR4705XfSHAD2k83iu
Ikups+FNMfiDgXZRdvXGkgrO7qia5tPXn2fXjqMLkLxgVXX3vlsS3OhGcnxiTIef7JqMVLqnbGHB
+iq11gLAM/Gh7Z9z9ysnq+Qkv5CQrVmtJNPqaaFEQAOpC5DkkRfKkBnOb7gzxSj9wJDMJdPX6q8/
meb8n6sBlG+Px1G9wRRCHXBair4z+czpCGvsWtufWAFDGopXfCwa/7EpsGtHIMoXmd5DLwvvD/13
2BUL1FSomeROF4cyac8F6Yei+jtpZqwyxJYoO5/LwEZbJR/b4J9gvvbdp/B9ib47vAiJNPB9eVEn
p5dpCkTac32Hv5QHa8EmLG1egYH4bPNq+oG2mITbHH47sAyQNqyUyp4EmLJWRUZaysFjNKXUZuMb
vjV2NEjsEEo7VXYthzxjucCtjJtiphjSgFGb4uBi9gI6KBd/2yC34/Nqpb0IhORmc+fld+EV4EXL
ZLx5YGGOh1nUUl+CRfr2lpqq5Qx6/WejmxgcpwN0nlsWO2SgwoUrpboBV0ASPr5CF9Lo8vRJQJyV
dqcT+Df//cRFzo3Ln2HZykGsEwDDTyK+tDzp9SRWTTW90J0f57+OazK7bea79g6NJ4Hcbm2HMH/N
2HZUlnEiLoARb71MrZVPqKoUfbCiyn5aocSqXYBt+PW5ee++0N/JWP+kD5j93xEl3J0qVyMHLwDx
Y8eUHBkPSbuECdaFKEB+BsSzYVH+h049M+yQwFekGQBcVFC1y0OTz3Ui7AhxEq9bOA6IsGJlqV8o
4NDqPANh10vqm8omtWsyvdRMSLl32zxl6pm2BXJ6Ja7LntR6jRYAL3l1b09xulETdN4M0LqkR8aN
jgi1IP2q85vmBGPicAwcXwcgySbBPMdDProtTHwSv9tn0Mdzr7lltkiuULt2QxBTnpZdq9JmbVcN
ymcb3CYJsNduOnUdQhpT+B3qFXowZxRb3GespR5oSpjofjSj2pwlzhEo8+l6W2DzMxTQi33eUaWm
JdrK1wCkP6KcZsN4homQ0X9wBG+tSMxCvYt8QSF1+RzkN/sFVv4ufRDJAJpu5hRVLH04IS34mQU/
O4zI5xCbA62+C1ML1JpqqxfwpPLk9qL3Owmvx4WmVtEN4qyHUfsbWCmaFOuYzzlZoS5Wq+jTLffD
4AStPM4EV0q7vmHFmKGb3TYhnzX4++BYqbI8kH/sYTvM2yUTDaksaW2+rI+KiHq6pTmHhWKgFwj6
rQRvCTe7t+bxLR2xgBpbpj6EUQql+TFwsGWAg69B+Zhfuw+/jziTe8wqGG4Gay0Ut2LyqaOpHi/5
f+3LUNrHWdKP8g2+Gchao6sA5vAtlj8AGz7tR+dba0ZH+aBsW6BaD4vd7/eyfPVVFr1CFILWWpUC
NORGhLj14kv3XUj12co2UcwArgeVDPHRq4DNaCZz9OOoXki4y9+W1shSF0I6qsY3nGHZxjz56C6/
/OpXGCckfFKaM1TDGvbuZI7hz5b8xWjseP/HFwRdq6yt5n2FJggnuwXaoKfEwqdVf738vvW2s62D
NSFr4cCLDFKFitP+FKmmsL/VKQR1T6hOB9QSi46o5Q0t3ereMH6JHplnCGc8JbXohupHA5D+yEo3
V5bhrHcHyJlGb5jG1yIyvuQFg9M7F1LhJTO6pnOHOQoaC1IdPN5OxxiWNBbV4/CIo56r+Qb69aE5
kPge7HP1MfAFo86+dnKlZtlOlN0Y4yKW+K2hOJSzw51KfgrWhVDcEjrb+LK0WI4wgjPVN0uuPqFT
IjfHWRvzHLdYh6DgdqLpm8h77d1jQ+faeXEojB9Z2rwcDiSiKlL1mnooT9TSStGVLEj4PZmUjA7w
s8NZwYwycun8WTppmipPIBsQOo8WyvsFBrybIA+x3IelHSOsWS+/YebpULP7iKtorcaCZ1C9H+Q8
DE7X1yeHNkkulp5viWng4RCABU93yz/fEteOI/DQ+IUnijcQOtDk7bECaLSVClAfbJxCoYQb5lJn
4LfXmI7H/2mZsE365ZlnI2ywD/MML+gpWPybmlU9vRSd3fNf27bz9OBV3KN5thjK+PR9CxGJ3G26
hhBy8tgZothE30wc/QvUCGi1ZibwPgTX1EblEInVyAX9KddI534yDiHK2RyYy8/czOaWjHNoq4cZ
viX/rtVw5j/U6ZQzVtSBv6peU3GV3Nfvj/ykrvQbqcUpcb28tWtW9v9+ih2jxoiAOgNSg3taQyoN
w3fgwsfIRRWIH/CYz4/XDJzaUzVAoRJxZ3FVvgvSHiaQ7PF1+s1UIi1RaPVDY6H5xkvBeIRlN+XK
7L4sDlif6mRd+yxvfgkxGTv6IAr437umLYFXuqD+D3WOiRwopvuJuG9xNBy8+AfaCXxUXKnv9LIN
gNR10TvcKVF15L9RfJzAzfAbs28O5ejToO1CvQegSbs1n4KKuT5TU2sK5z11NR7whXGW/2B9n562
lgxQP4g9LIpVEEt/+8EJf1HlO4FEPYbTwIksO71KkxUHuxE9Q4UCN0BCbnXYThAvRbW4sjuLv4VI
PjqD2OA0CrET2mmVUA4cVy5tEkp/ZQjkEAknKltRCpVHqT4so9mU/HZuVPjRrEsCxtNXvXeGFYA2
TFvliseYXy2XfqCgMPeKTE5FwObLDr7As4YfHn8naU6IltwpmKWL8AHStPxlw3uqItRa9xrMZq7j
vYBleyQXiYYoyEFuKTzxj2p+gMFlfTSoRxSw4RPUmsXO3091n813pG7y76nPR4wR1F7DyYZQ8mt8
VKT20SwD4CH6S0sRwF9ekTMi2RuG0RPffgQbO/GWavwVjY372IGWcrG6H9VyaOiFY+bZRMNQLhu/
EyoXaYmDlS6y7nH50QDs0lHpHz+PmXpPLYgL2ExBou2HHAaXTHvhbkf5oZ754K3BaXMLI5MtTzrs
J5JCdBt9oeaAmnX2mwpm4pW1b2loXwSLuXRZB13o2vuICAG7KdIzCDkYNwHuBDcrQm29vUtdP9kC
9lP914w3LjBZihEAFzyBJpq8NcwcYBUoDGAOe5mPLldGsJke0zdD7iVjcdUgF9U4+y3T0toPxjKU
FiQvd0tr/xgStKOcXpn2N6SKFVD/3L62Vf8/elpwP6qoCAWQvNZfZnNmMYDt5quDMUOufcqA3m2S
CZZ5uWq/Yny+Uv1RF/mWGuZOzORyIr7Tev1EX4uqdYdmka3NaTCcq3RwDpVxzJ1+0ZOejqhVwbB+
czRFCz+gEgG35R41JZBkgB/r80SUSPUH8gFbXV+oPwMXdDWLXc2g+XBw8rcKxLR9VnLwvo317GsF
IvDM6joq0NKEdDP1gODtpp3iaNH1qkGxXzeceWu2fLRNE+Datlwxixzt4X4C50KmXt8lmkZaUuSR
IcBNc9YSJHbe81aWzZrGbE0yM44dP6//FOH+Ae7+PBzmy+513p3MQ4a68jb+i1ZJ65uYvwSHlLMl
kwPw/GI8B60Ru5ITsMgUCViL32UPLM0jioAtWlXsXzAFS0Ozi43eWF6UIUvO/I0UTMVWHif64R5F
SOOXzkmQ8StKHx/FEisPxXu9Kjl2J7shglDs6iJP3gXBMb59oQxvIJPtizr87oqJXrpYzsNxIEP/
JJghW6km/yLi+i6FTemv9Da2726ztvD0dlnHd1jl+cNvxHrhv0xEkUh1ew877GD1tygSgDSKxWcr
iHIVZddDIBea5GAbDlZ/oEERRnavnqbaYfDrhhzKt15SqHUjNE+yQt0iDAj5doshMhcAl5mKFiZd
MF91/M80TSi58it2UpVxtnyldjKyFFJWDG9WNc9skLqeVcX4+g/+XKvwhXHWPsgThwbok5SYwBcA
risTDIb3azFgvWy61NnILPHam1tCpYFGxT50IBpraohRIBzUH04zPqbe8bW053nb378hBIrnHOTO
TB6sSk6+oZIdt7e2hwYvXmAlrMhD4Cfz103++IT1SOYBWADlrQlcBi9jlr+cVgBDDtaYIsfvLmqd
6wU8VkPDbH97+V0flJZyeEI9KfGqRK2v+JrMnBgclWNsG/mqW0wmC2BC0Finlma/GiEckRzoEmKe
qML8T02ICkn1nqvUDsMmESxoDBlT7U1olLhDw5qNNyLLc2jAWvV53880pwnB0js9CLhHBO5T0Wfw
5szOgXjJVoaXEu4lZ4wg2H4wY6uJn4tSdYRSQm7XRyWRyrFW74+iVCfbXYFbzcQsv5xCxOyS4+Jt
sgISmieHhh+gVfiXvFQOVQusUTc7/y3n8vLSTmjqYq/REzGmw2GZT7KFY4kA4ZtL7uUMwEZ9+U4F
DZSdHh1bM4BG+1D0kglNmvSDC2Q5j20NqMKtBmKpfNxy8gxrFUMHvTDf97Oo16isRloc25YEvN61
sbymgk8Y55TEvHFdckWCdJJbNqXDAuFCELlJEHjIdMstUQyq1oGbXr/gCb/ZGYtloe++JrNFuDeI
lguljvmcNYiC94tiyfnIo1xFjdT9+6NsH6dSqjN7vW3JF6fTfUrjOr+yablZGKMMhzMlX7VDtuUl
Sz4dEsv22y6KlGsbCwwvtghuUOS+R6kLkZhLiuLRHPFEPsjHl2JIUI/PFiay5AaFn0P08sINMmYb
Epxv71kxH9BWzu4FRI0MsfCK2muGcbV2sHQ6sg/K+8gOIMIY41+/RYuMjpa8gKonuiqvD6sfUjNo
DN8joy5Rk1OOrFQ8jEQWr0wc/kRXp1YQYaYzqQhV6aKFCSgq+Oat1WBbYwN3Od1hETHPvfC2j5HT
uk5yoYGmd1LjpLUggHDsMkvep+SjFnTG8XFDlb7B6d4eO7kHHyn8xRa5k7fZb6BbQQty+S8D+JuG
HguR8WsQuMmvtwhjzu7nEcZnQJqTLWIwcaZei3Fxvcov751jV4LxP9kY11/Rz+Yk04WKBwyVrDRr
a0A10bqTHvowooMWt/UVTmZQycZoMBYhEfA3ijsrNmsXx3AIkCwhf7BLb+nclkbJSKanzENVDgUc
sHTw92dkJhIWTiAG3WNhtgk1Upxm3eQMp8oo9EoGyf5+J2dOBoQQuWxyqoi9t7L1+QidweIHRLai
VbH35oWdmzHrAtSD2cKwZKz0tsn5iKy+ODw4rxgfztiXlmVqZaWl+e9K2DAczVE4GrWHWIp+6TkJ
3MsXsFejD45jEFCTZozlcaHLtACNL+tOYb9o/c+IwcHa/LoQfXrx63J2oamP9q8DaMN0f7yU6a7R
hZFwF+d48TdeWyUWDwYKEV2lMoLI2ED7bfdpSQDYKGDw2+4+rQ7yj36QLuA5mhiS4mzDk9KlPMB5
2HExfckidh3U5ClUcd4/r/OlYypbtbpBYuOlTEs9UJGMno0ZvKMq0fUJoI0Dt6nYJPnfXXUMLZxh
wFY8ZfCD81zu6BGzGPnQULgNDBhMlDlSYHrV77X9TwYCgtSfzfuvY7eWua2j1zpn9BxPEKR/kMPG
0P5iOP8z22vTKh6FLyBy0UDs0kEpOsiOfESRvT8zAgvfqyqoRHfDtvdtbr3RVgeJ7Tck3uJU9dqG
zmy9BUHzCr1cYUcYPX76pYHkX1onXFuF0INLcLJeanEY5DPSg3nmoWpiNILc0m4xuSIa1ApWN1Cg
elkCodkURLVtJp8eq/26dPwcRBoJU/fhvbcL/34Q8mi7yD4zh8HInCtPkXxHSfSVPaL+briSfemZ
z6pjk80YJ8epOQRtnMt0r7kqRCNUc7bMZy0Zv6qa8WUW0Pe/6fl4FoUr4AMtFucUwVcqisC/joeK
0wcwdOk1pQ6t6KlzE0eRVfn6bPKMMZs78IU4q7fjmVO9TwfunflgbJOZzP7Jdm6KuuhSi8ZJ4i1Q
vSfa/vgYYZEcAhr/tTqdCizGucxC1tQuTsIvUTLO4sFEzws9ND5rpvkDSNW5wfBjkIJrzH7c759v
1Itkz66X4Urr1JzBrfJqsVrqo8qMYxmAdcohfEPpDTn9IsQ3UhfbmRPptAuaQB4lPMpA881H+nhW
nLb2qCiDxudiukh0m2UccVGj54DNQzYQmsWbDWph7T9BWnrEgXm/ZsJUcr3i6a3hReirbx8p+4oF
Wo+bbqoLmEADb+PwAFlMaSVNFYwcVw35ojyrJNp90uBsL5hKVZmr7MGQXI9vU7gwakR9TfRzAjZZ
6da0Jgn8+P/y6SQB+Gy7cOjxvNvnRipWP3agsbDMr4MXb6tlQg5omIrVRsrmT4eaUcVZ29HrKHP5
PudZ0Rwp+bXYQVgOZ1dFRgdMiZs2DPmu4V8rcpwaaoicuBdo5cpxKLrSKZVPUI/5mkjNv576+1bX
nYn3n3qqdX+JTnm+pr3/epEkO9u9k2TaEMWcr6lcdV0NpGcwN5ejX2iw3laY4tB+aiEM7MZsA/V2
2fcezeoKWpG20AfyQQzxZNcva/Xm/cQpO0pcozZ686GmZPv3sM5kncBXSt2Pn8BHqCpUOSOE9kG7
uqwrS5myH3Iu4oQjDfuCD3cjel/tylontmbv1Sn8fiQNMB2lF6MPujK9esmwSYpd0Uazbxsshy4x
B0ZPoP4MrX8sgWkh9pe9s/TZ5deThYn3g/r6svn4chhfWizkt7FDK8DPsBSX+hmskKtApX+c/aye
GTh3m+m7FpFOjlAeopdvLzcq2ZW0E8HhW42bGvjuCUBOt9bHz0v8YfVtfXgLjkbaLM6Di1LZN2gB
wOmNTfFO9PM7LepVLzxrwHVs3B0kDbS17tBc3cGbY0g9kMvhXv0c7wGSToJEiP/aIsPxSgCTjKiS
tJYTu9n52RJ7y78qehBwoxWMusVRbp0qj4g3kRre6CRb3c6xAfiyYwAiC+wJKkb1nrjtXL0JAkZQ
zxdCOtk7fKjn3F8TM9lDMY+3C3EsXxcBockRMtL0Ni+XT5Nn/hJ3yTNmqn1MZEuGEM5YFCTYPybC
YBP7p/7NVI9SFfsj3uacUvTN2vMCvYL8SxDBuTiZ8ACD3huYu+US0jBEiPDmNEmr8T4Rb3aO4mac
Dv3kDpO5yp2pba96SggS04sliYFKQB1+b0pBPnDXVB3TiutJwzIP6KBa2MaWIS3obCI5oFcKWRKn
D7B28TlMH6B+ScgtKRNOmzdGb3Z4HC8hiD/G0j1FKjN9oii1HX54C7dX5hsZzk0ZgrR2uoCRG7Av
S9A3l3Jdur7t+JRPzxl8r+nDcjW9zpOYL3x49FMai6PFMAVz29cR6ceE59p90nOwSsR4fjArPC0Z
NjRU3IMinPa2no87IeBQWn7xCmJQ7EaHNWoBK3GDgHFAJjTRsxmBPHPcQaffeYL937wOvm5GX2Vt
I3cjTNHwIFHXC0LaFYHHODVPzJyJVMvJ5r4iYPF0By6R9WjUOpDick01c0vKJg9c2Ty02MYbUVhz
J4W7VsWyEVa+Xys2IEB4Peg0/2xdytUBLr+pNxZW5Ea57jnov/NQnMtLTPhUyTF1veoKRIaWkRGw
Il59K4YQQRe1jePl1x9g1UEqEHyr6shwTJgYmYWtIpm1t5s6fVXLSVdNKyiFK5xFEy8EvMNaBRcS
Z6/Hq5t+zyKZgTN/sKbt9gy6BceD+ez7wRzspol/4NzOwHqqJcqAsZYiOD3n1LcANWe0ZFXmHgmm
CfHGcdrupLKiPVqEpW6GGrEB6ZJn3H+N+QQLffEoldrd9nKH0rrglH9EGl12KLLZG4AAmX9v79H+
3D+m2m2khS2d6KHtt42cp2Dm6pKHadYmEaN3yZcgdou2LWtKkFJhYb13QrNpuOyqcPWx5EYv/SWZ
68AeQBVntEXx4BCLW42c06hmre730zZatXVFdKb/D3WnqqGQEqAkfVXTSTPFzE23cm8z8lQh42Y2
YFEbPl3EPoeIGDqELNGqSXZZkw/xnxeUk564herHjyhpMnrX5tci1BSi/NZyqq5YU5h/IxdRWtb4
Q7YMNx7yKlUkqdbkpvnNSPHYiBxmlmjkS5ptyiYCqt4DZbrrmDkLvPaWxg2LGgrJKBPPQGVmZoaX
32kVYftPxWCAYVw4gBMn+IxhmJ2nMW00Xs1JHeWHXW1XYG0pud255pnbuNXEUDtRtBD2FmQ5/wel
Sd6y/mBQzj6/NImo3zyEsMRk9uSgawZrASyWylusYEcN7esVmMMSlBW4fuAS+C+DsJbjgTrdI1D+
N+Dy/JTsz1wEec1DYv5J7hzlR81Tfc0/Ih2NPUnY8XQ4FNRYD/OqjUBmRb6FGiZv3GfujrkrS1pJ
cnHQA/asioOzoAGuhjYOlSlEGfjIoO8DRnzjxLRQWC5nhJ+ASv1ubZCU9KyJ3cSU8tlT6e5y4WOF
HRTeAR/gOYr+Jtvf3myYtklTLJI+WTeed7b150igWkYXRCY4wG5qP+B2mZ2H2fp2s1A4IPUSVxYa
EAmM4TXbzFGM3afZ5TRLmmJhgY+TW/NuJiszCdAf0WR0XfzRaIXr/L2wFR7mgvB2jo5T/bXEZhHs
13bTAvw+5dw8kgoT/12GT0qzn5ub7UtlkeVvWGSJ16TjE6AYJw7ZFV0BLBLKNxZMNkFXOpJHazx5
Od84S9B2Qw9IuUSuJGbJmwvq0b9y49X4cZRKi69w4dMQhzJ7DIeWIA3BwleaSO9Ge4lr1Fm+V9xN
5Yr0QjVpzZX8DzOXzNDBtcL95NW0eClk+3gg6OCpHWKCkb5EYATtHo+zyM0/8Hg7fDJkepAQ+K0o
wlnFVjqmxSDGRl+92nAlg3z89/+fBXxaH2fbYn/QGO1SYRXBiBsT+tgGeP9qsPGAWTythqvbj85S
2JeEX0ahLOilJQeHD3VvxafBTjDbyE5B5PC8uSl8yN34/+c7s5nuZaTWMMbKw/fcM5raL+A/yAle
n6fljbdo0sN7Yrse55Qfd6mfcfjZC6b/tL0wv/Kgs9czZm+w8dFqGxHZm7FOFiA8SsexYP7Lobt0
sY9MsYkieNBRjR+TMFIc5GmZ+21gp8Is5MSOiVo3qwLYrucppCIxqTb0trxYH+7UiW04ni/aBsqK
ch0co3fEl4u1qY05DBnouB41xLanxn+vJl0LMuFMeopYZc4SdjHcmmloGgKqC6M3AATVVoHlGfIR
lWnqaTcUQBaAyLj5rVJr39PFjLLc33D0uNdRiGT1pFA87ju0CR/axBApS8laIL1tGM7PVJjkW9g5
T13aVcFOsY//vph3b4j/SKsrbTL7u/4WIgCFCj0gQlqtCm5D7XuAPSkrsFIdGFTxtsuQPFV41CHq
sGACnV3M0IsNtfbeKwywBXQhunRBjd8THD/Zd4vfDUuD85wgu4pOToKq+kuwFtiuDZDHILtThd22
8Eq+MTdJqjb5gcS048TypTuAuJekU0AYupmz6Lou8PpgCeHOd/Y2cep3V+7Qv9hKN69Ib1KEqtkG
6AXrLyEUuhIq1+dS0yZyuNYRV7iPaW+jafAUCh0yHgSxV/UzXt2eccZeLRa1xLW6so34kicMnr+O
geQdtBbNir3YBwPZt2eGo8gGDeoD8jtuyDvkYgOJpiTM696qgMhxI8tNrvyqkdpwV09aU8cTaCrb
ltKz4iQAwTuNVKDpNjGExUuBgmERIPpjWjrNkHIFd6G5IHCMFH8eiuiu33Q68VOb4y49pt1XmBYj
Tn2zVDMj47P+udIeyHbXUAKFBPHO1GHuZypi2n3AbobLaQrWQpxbXfmFjeecU5WeHqjV0VtbO8rm
jEr9a3uIgWYe3A6bAD9M4TAYmZfvR13nMfec1ryR29yXFyB6KNgSTh+9SNg0Cf7MYFEPgjekHkEt
8VzNT1QUUBSJhvlWIlV2nl8TSVRKVdXGISWxRl8Wq2I4e+Pzv4/bfCnjs9hkH2WAT04zfGmrLWa9
u+07ak6CWz5BkFu5AWCI2cf65BENo+e9eVCuUm8ccr0ZkGK/vsaTSOmvPVj4ZRrn3Pej3pK0ZyWG
CsrcsxbVMBF3P8snLHmDLe3yONPJ8VIj7Bf6OlwefWGUyqpvuFfIiaov/DjyJqrDkTqSQzntwJj2
3yUmf21weHnLXD/jbyzQQo3E9dWnkObSXTVin8fvNVgwtO9MR3cTMwxasyRq+MMPASZXpBkUOzTg
OEPiFPNyegI/p9oV2TRaCB1rciL1o2IGVRxezylpK7o0/WOUSvY0pgZ2JRCIhKMj0cgcLmuJOZfI
VfAESxZVIV1tQqQi6+yIsuo34TzdAH9Q7V3E8VXRn2swAztoOU4jNlU6yUHAXFo+AOdeLRpk83y/
v+eURoiRTw0nW6N/YZQVPBt47SvagWAD1PIpZmqpsUWMm5ugLQ9kFvmuSE3hSfpS8gNK7ZFm6Tpd
w6bTJjn8gsH+srmzk/cV0XMVWHpxmcgH+row7/gY3mZ+KijKfPI9027z8aPasGynuXngWhO71zy3
BX1N/aj85qCugfQVLhHV8sCY6vnjWz35v3dojCpx3L4db/783+xRREPKLDP5Fn3ZJXFcp5rxEA6O
XBeXV0mhjERhtOF7vaEjWSe+SIXT4RDIVlR+tbpC9Kv7o7gyZX510KFn1qtJ1Qy3wOkgXp/gXy8N
pTtiXDebg7//ycqw0Gdb2bJDSBWIgOFA+1sKEU5pDaHaXWU2ycqcMn6hPBfhkJJs7lmIgZlfHUtk
FFKUgWJ4Z6qzl3a/LuBw5mqFIbZAmyvTuY5FcjWEJN0/UJLdlQHCs3U3z1G5MzgyG+FExvc2mZi4
e3j9ShAEtysBy0Z4vfoNkRWCZviWWm7iemr9rlY0kmk984L3O8Sou3B/IospDYN55r6kb+RbeLg+
74ZzYiemwa32Qny2j4dB5hWrdIg3CQauZ64f4VX8xCEstRMOlV3amaCXRfrylrDMaoowTaya4v8v
MjfJRtDaMQN+BZUnRGhozSj/Hj8E9aLMr+53cebekQh+ribAdlblv+Em5edAz08HYXTCt5HAdKBq
kvYo+TEbgxXCRtt5KAaMEkB2Wdu4ov9CTwC6Ag6iq98bSsZSPEF04TlDtiuBtIRBe6LBHJsasZlE
dj7A7UKn2h3ZY/hI0QRgUkEYKoUVln0JAG+/0TSjoKu0GmAZeVaXfqRCLIIIRk0ssb5pC9veQCg1
0JGO9tYLQDm5PAqVkbzv7uWmPJDlEdzcPSRC75eCGz0FxOj50stqRZ2veishsmMlTUQCvbxasDeQ
LqEfO3QQVyfPPk9TPAXV8Bb4C7XZJDFQJb8vXVmri4KJhCr73oUmhTQlQsITOB6Zs0e1h1fiiMvT
HHHmXq0Rq/Lj5dl+oWi4Q2YJpd0HkhzYTjFyHW9R+juYwUFvwP1fu5zYVJXv8i8TdWYw3Mjsqwfv
rwrEjBR492gafz489hqQ8NMmJDSg2j9jUdE2HiLzgWoh/CnVZDcIfAsL0m3vFyx2SQe5Pmy6Sbk9
vGKLaUup44B9/oInY9zdGK82Porl4H98m3YHoEiHSwxGQkfUrhmbCNh5JQ5zBgzbNKMniP3yBz0H
QLIFiYTwBLsKWtP42DreMFMh9rNlWqovFL3F2mvjDJahgVSSM4TvDZihqHrHZw++US9WAZ0gs6vQ
F700bgIvcGNpu8iiXBVD+QiKBdYFnW+wKPZuQCw=
`protect end_protected
