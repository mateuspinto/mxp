��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l����$B'���1�5�i������~�S�$�L%�<R��P�A%�.X" ��o���g�TR��F�X%��/�O5R�f�h�|{�9Z�y�G�L������i�3�m��b����ZM�:U���w!<Q�qs��؁����2�K:�(���_e�2�~�����7Vҟ��L�2�j{���N0��������l8�o��W�ښF��\}�`���տA��z3K���8�[�,�J��PJ!�s�!��i[���I3Js���e��
"vTOV�����=�(<��Iˍ�zCF}d:o�u�h2 |�Pϴxqz;9?�FhA�y��X)J�%`���Z�0ı_iƔ�vh�rA!qz���V�\������Z]��B؂,�.����k����\�}�ֺ0�*�x%�6���6s�`@�%��x���:a�+¹PQQA)8���(x덦�l��}í~�%g���y���vN؉�b�_�.�2'�h.��
S>��{RH������K�%�z�%�@ڕ�>:t��;�L�o�Ԓ&`K�τ�S�B�הiEa�D��:Y�?�����6���l2�'jʱ��:XoC�)��0���̶W��OM��D �e)\���2��\�H�v����w�M�F:�J�!�S��b��X���n��tȺa����։;@U��\��8��|G���O���*��d�/�ӌD���i4�n�ΟT�]�3��@�rD�� `޽욿3G�}��,Wi�Ҏ��ᗝfX���5u���8�pܡ�7t��t����KmN:.�>V��bG�*�1ԨɌ-�.���ʇ泅����Xd̤z��šb*�A
z�h��~Ү�e1  [;�&�O�?x�B0,>�y3{!���4s��h�r��kR����2	:Fb
�N�9���]~+��v66F���Д���C)�<�Z.W�ƞ%s�5߁���/2LӸ�9��~V"���q�eK*Z��~�m�9��4Y�U4_��-�uV��æ�P���Xt���$A�]֓���W6ş�u�j����up�:@2��F��](Ф�D�?2��eb��+˾�$.��\�_T�eK;�O�O��,�:V�5�n9���.�!� R9v]�4��J˂6�>j8Q�����a��Jl�8�C��YY�)6k=O�5e.'>h�#�O�
��zP2 �:�M���C!��%�ـ�c�u�nL+sw��϶�?)U��]��i�8��	�TK��W,#H���e�3sC8�7V�z���PL7b8�V��>�K������t���:5�o�Ri��Z̬=i<�M���7ӿ�T;��׃��v-��y���;Q�m>M�%Ƅi*�R�T��ǋrC	ƋM���IU{X|-	�=e���S(UW�
,�)���@��tl"5.��[�/��_E쪘�<�i�Mߖƾ>��q��u��� �B!����Vǡ��*-��/\7�t���U��#b�x���ҞhT[��B��+���b4@���Q�-��D�w��wZ��cV�-f�F��Ԕο�c��j4`��B�l��n&-�w��p�p��˷������X��'ن��駳,�s��O8l��H�f��F�'�IX,�!|�;���#�7.9�-����S}$�"���-�Uw[Q���K�ЌrV�T���8�C<���\Q(I��[?���]9��D�h�Іk���]�����`�-�ᢗ����(����O��|���}D1#�Xv5�O��F�կM��B�o�'Dx--��峔�*Qw�P���.�V;����>J���w��Y����f�v�52j�)3}�����T�Z}5�?�Y�"�;�T���@�X՝J��Z�	�7)��S��������P���Al���[�/��([#���~y	����ũ��ѩ�T-�2�¸CE�T���M��z���M[�_+X�d��&��obi���+��1PT�Ke^��G�0���X���\���8Ŋ��׋ޝ2�2�e,��u�\���-#�N�~�s�@�8���� 0�:�k�K��Դ�*N�Gy�3q��p�m��)T�B/2��~Iz�:��e��C���L��)� �My<�x`P��ъ�o+���^.��}�fz�p(��x�S��f�%���Mw� Q�&p4�a���[�ƻcD���}�!��\��+�$�M����M����c�Lt��U�aX~�^D�#)�X6L��!��Ka�[Q�!A$�g�G��='�X�Hȋ?<�'��j"\��4��q�=_��1���+)o�@��ւ�ܶ��mR�K�
]�����d�=$vI��֑��6d���K�5�W�XQ�n
�?{-��P!܌,��7h:������DxYmD��|Xn��I{u���&�b!{���K���b���n��'Y2$��di�h��{Y9)Cb����z<N/�����\�U	�^��haX����Ɖ�ބ���8d|��3F�"��G�<S�����
I�*��B��v��� ����\�b�����B�aT�?(uZX�i�f�x9��4���(+2�ϔ�9�kha��4�@�����Vۖ�.�R�q��5��qz�-`'����9_�NPI���bQ��'^����b��C�2�Z��&���Nn@�\J=4%�z�'�K��v���q �?�Y�R����Tぴ����j�j��gؚU��P��c�e�c�j"�U&�g�ߤ�����|;*�,W��iP����^A�>�_3�{Fp�R�9��Z|u%c��ve*���C)юvx��2�Vd!��V��4��2����P�p[p��Y�i��?��#=��_؞��ĖX��r���t�+T'Ԕ�=�f ��a��F�c �M�8t���и�iź\(0�^��V�������V֫��n1/>w(���砗f&��cx[YZ��#H����
�9���(4*�"1k���c\�̗ �F$q�Đy��\	�ဵ�¾6X�𹏇ۀ_��Z�і�:�q�7��n_4 �a����uBlPS��pE`9��i��w'���X[#!�_�'�V?]�P�1�N]�+0����W���9�F���x���V
/�W��9��θq�������}�x%gx��0,���L|����^���_HA���4�P�IH��o��E�L'u�F���ZVAH��˟3��؄��Y�x+1ػ�����YI=�,���4Rږ����0-��n=���,�����^�GF��/��d�6WR�.9�&������H��J��Jv��1�'�nL�E'N΃�W�.H�(�+������� 㪏��}1H	r��2�"��0�3X�YK�%�!B麺9�v�����P�_�W=�/j���RHaSb.��R-�t�����ҝeri�ґ�0�0x�2���r����g�z��u�I�h���/1N����2�}�I�8K�^�ԡ���ɨ�vW��=�ۘ~8Wkm_�?;G��%dr�O�`���0'l-uI���0���?�?�!�J�}]�F�c=3�c��7�o�\����1�|UO��g�