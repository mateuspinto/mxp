`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 50912)
`protect data_block
Clhazwkz4lgeC2yQFCTLEsWzuuhjSabWTcqzQOd3u8PHNqly4Xli/Uqjqf5XZjTGEF/Epwoa+WPB
y6EqC0DOj4luSipZYNhRWIyG16ggwnwZf6rYBOJG9emAllgXLFF/40ZVJBcRGWHPU8DXG3yn2CYF
obGcU2yK2oXyezGlgcR7tOoRRWVbYACS40F/68q2aG7hUA6EvReLvNafhVvMU9ceFSZ0flCuQ+Aj
O49AEnvqqBQiqMDuA74brtpnnIHDsm/mHn7IMO2iLlG+FMiIeBmBamBB8jzc2p+otGNLN/+YWMYO
9w9XDon8M9c2sFefRyOczQoZsIESB3DMmO/Da7oaqbf39XgDnC+oHvo5zc3P33uW5/OyC1+DF2j9
m3lSzLb64u0gX8kljXi6rO9+5ZfKHjU3XTG7PSvwOMPra5GexWGMcE9Mvs5hCP0Cl5Wq42CvYPRq
2mP9/tY91Hx3MGINM+OgWimXxVMiZ74Ur8VCUMZW7oRPbFuPVMnmHwQ960xGIeUXgyxq9R+sCnqQ
AfT1CcNpZ7MXLoiwyfs3yp0d/P10fMsaKZ4SgybLphAdquk2u1b15Al47tDQFAGu9kCpxz9/cPSU
Jho6xFIBdToAg482xwS+tzSCU0swSoIRVI4qyRj/E6Xp+eXNU1EpGRu/8RRdCMeQjTM33E+dSRYL
lLhTGzyhhmRRdtFa3hfZGMJiEovbp8uGU2tER5u3HgXPjeYXfDXe4YV1mcXcUpahRFOb5DwnaHlQ
IoCvy/rgYyKBpERkAaBAJwNKqpIdkmag/QbK+LkyjWpvGGuIbhP87vJ+w22EULEeKf/sX8Tcjt26
MEAppw5ps7WuR+dVsgbJWkLEWHnnYLbJImPQVHuKr2T7g6jTFm2zZzcQ61aRlLJBjJ5bQnIEu27q
22Dk+E1Pigm6qQ+o5ygQHBsrQBvrNXiO95/sEF4sn+qCU1IHzEOdSoTRSEXC1RNBnNYW8hS2klQS
9mXMWwzXKAC+5dso2nIi2Vk8EClUfaVC/IPRAh4yau22lKa+k6HDYCqUrLkVPsBgZSbjfucyLPrg
XfQksqmrpZSthz5yqppEElgq5M2QNlWXDKJC2/gX0SeE9dY0Z8uy3KPxinuX4V2eYUlcDJ2mFZJh
Rx+z2Bl//CFHwxEYFkaxVUSmTLMgeYtXGwVLixCcgfX1/rOFenDk1lrAYQF0vJFbkDlNME7Sh+Vk
a6Lax09HybR6DF9ypr8cBeyETtE2LWWuUxJ2f26y4ildOWH0hAw+6ChzfvlcBMgxWESDN6Zu7Qlk
CC80qlCh7V6ElCzDm/puJofYBYIXp44w6xcTxj3H/sCDHwfd7TEvfrbX3i+s5vg0Soa0rgeWAT/6
JVurg0y1+4NRrX8XNIll5gTOtxcpcwjLp/bz8OZHS/caCtNSuOcicTzMMFi6t/JKo416s7YekQb9
wmQv2/Oa+xdv0gd39S9iSARO2wJ3T4pCFllbclSuu845OwIYfSKoz6stXxf9o/0NLdoIvx4Mifsx
oiFPn2fIysnOZ2eKVfRmYfNuLHvyQ7/H4b4ARiMfWwlxfMajlr/Ji1onN2G5QDt6+k77sHLfU1pc
Gap0x11KpoE2oEMp/KZ4ZQublnaVRMyVWJjM09v0vvE0nqEx7GiODMa7KJcgvsi9S8ncmNpf7LJs
3qNCQSYeqDSeuSt6ECMoAXCHW/r2ASkxXqxDF3sKwvWtF8DD117IgrZTtbQpkRCGNZNJErCzfbO0
YjOURDjYpkaVmLbcV0K0huhmhnbePWXWUhe9JYr6Tev9JNYT6vQptv/5HHWVerBAG24fDgGuQUHF
5bEdex+egaFvLj/P6dTDUvDw0UBeVXdizW15zzxPngxAb+n6MI6ljV5UXNUZ2oLdtzZzDNJtsEqn
fXoEZs3IB19UiFfIOOmWU9yTSQaX7b6FQ5iBr+dfWi0A+VeBPP4ND8Au75k0KSUXnox/msBY1VPc
deh4BxyKf58B2PCPEn41UMXOSwJ8PvPAm9hFyo+0vcg5R6bGXNtJyx9wid94jgSlV8r0QbaBe0ku
YlCv9x6UJ7J1YIZGOiNhqayD87BIGc42JWAaWna2OrBlytZkgldNR7SUSZEjrcwHz9deOjss7ZOu
mvOAKyRjpb4c1G6LZMiMckYpQ5cT3gOZl4PmIB4RlFJFmh7JyRzJK5zDuA4uFOCh6REGUU3Ivmog
GWNuH/Xt48AbT/eLwPsHRREsetBZIjDoLOFUjsQAH0KDks2Qd6F8NLqCU65XSWrTcoc0FnjS4ENf
pNdM+XRd13eAOmqnkQoSrFLcBVOAF+ea1ayPeGDfimetE0GoyTvFDXrCU3VoPwIfVHn4eHMwMI+v
RLypfOo5IJ6V249F5Bfi91bHOmbpIY4cgc29zosODNXH1jpXBqoaKQipz9/t67kf211AA2lf9qoR
MumKNtglqGC0fFGls9crDcADM/dDiX4QgV7R50gz/J1e0z4XSYuntQwEsOGLzwKGgPQ7NMLJSqM0
sNzaMjYh9Lfjow6qAMDFHNoaemQi+pF1oFJpGdaJbwBg+0w49sAKq8hv18CpVQZxjM/SpMZfJuI4
Qm5FW6KRmlG2xrE1DMgGtjrT6MPdhRzl/+dW8lZHj8JVfgTdanOLJ0zEL2dtWOpqq6IUeJVg3ZYB
2nVCPB+VsLbdXZgOdwuKo8K5pwJFA/1hhYAEJrIvh8DUm7Sk4q5z9Agxh5hx/MYiq4Bmp25y+HE+
FUic+dw9HO+76N3Kp4JlHuF6LWLCAyxycyKHgnkGCfdfzMh73N1p4s9FE+Lt7Drz1Pu5SeG1yI9R
zhVgc+n4BfrExia3VfKq26TH3TxHsSG+93o4h5RObXLbJfVEIy4yrFxBF3SBrPjpwAgeSrnecp6y
3+LPQX/TlB36ymEWVc1u/SBlhNgNicvqTuFkj/pfKmEB3tyhtX9IjxEbCBOpTWg4h2t0Tp41c6lZ
ReTpBjFtsX8YwfWyMYuA4MAXx9csu31/9kSGe4qs0qq28Qe5PZRAKr5xRzg5PFrAni77KaFBVVPh
Val2jUQKsFiwlMCsbGfR6B3VzJzbcLf3G3FYzskL9W1AcackR+IiDP01g4XOTw8J8sXkUYAbBqck
vrtPz/UJLgZAV5SsSF6rSA6Oudo85ofDIHaNVcEZB06YWzqAB2Ykic/uCjI2a3vrsudAV5Q2DuQ/
IpoxMxvMQg0xjcTWUXyGCxQTx8OHojUkm3RqnBuYb6BUJGWNb3NLjo5ELDQO60azdqWlTL/+qhUU
WSAbG0X4O6bsSlroJgpNeGX3cCaLsjao7VM5XYe8B+Cl5utV4Ye52W2XDwy9VEBn1drYMImar4Od
WWC3WqMzFeNAMc2B8Ju70IYZMNr3BhuNWzntKW8GD5623YCWHhijf3NsMw7MEnW81gmHNnbEoksu
80MxPp3bE/Mw2j3bUMKMSG5aoitiU2ALx8SKvUq5K6nR8LLfwsh16Gu+WcyiLqDAWAaKSC3PFu9c
G9QIZDHTYd33SRLke6ukeV8JLUMCiEYeGkaeEdHI1lEblpdzY8+Sg0WGZGGiu/gduzqEFKFg47/m
KOTPMYi6b7C3ZL/99AaFGQctZO+uVpC4oF/ROyuN5oiFid2cQKfU4ODAZWDbz8zyEqRzwHTV9w/0
faI5LgAD0YhQpQM6p30RtBGBwzRKlPAAqdhb3QTWlwvO+6USlW+XkwuNmqekah/bFQPkGf1Ck3eT
MhnYeZ4ajPs9K1WiCSu1qpf6Q6gze7F2KkKho37XXbxXEvfZM4JMJeeQK5xHyfDR/Z3Q7FcgVYnw
6/m261jwuLyjHluyE3UUkM8GBhnoNOClA6qTGGtNrFBD9OA2gPBPFrJRP0UEcCLlBl7w02kdUeDT
q/f6f5wnFAsWwq/exunTrGYTn9/Syop3yNmfQTvJaUXBL3jtG+Zi8pwcQs5YN3BPTeQdu0bUXN1p
8br+bhuiscwOaWrmzTw/EJRl15IGkBtvWhqaBiDbxIn3QGhqkTn6M3B0206+GdMt5NPlmy0M4ZiQ
Mza8ps7Kdf2XQMcn/ShuydUbNc08lTBoPdbvG3LLD4nu8FgglOk14gQjd74lLpNloos5tPrZOONI
4AT0bxHRQdNM1JV0jc8s1H86knZr6jMy94wwzdEJI48fILsiObjf5CvJKZAbmHYDSAEvhiriEAJH
+dl83VpHdxVlIdQ9yi2r/Z/MfMs7n774so8PvLy8j6zI3tPXx4bbJ+Iwvw5+NCGuuoN25RKjmPVN
NFmZ3swvNTsI59tioGLg0n7DTZrGItpRYF4h7H4LXISsZko35/BvsHYMl8c/B89sfJvyZ+LlNEcj
M8/a1w3UPs0OnX7Z+zISKkALuKalLOCzXjQYnY2gmXumSKAVTZtMwFpApqBUj2fyk/xiTsQo4J8F
A0CdmUo2GvzsUt/WMv4eHmfSndhJwTeOL+fPPrZXQD+Wdm1Ie2ygb/sXqH55Dw8K/o2qxxOEyJIA
aHrs5UWja1IEPNE/JSv0LkDh8MLS123w5ZcWNoGnpM3WC1sJhKgAJit9EsPOVC9YtgWd7Hht1l9E
FudLnnIXC6CJzKmhLI35p/CLI61Pg3sBNDP4LrVfpbPo++gFRUiYIodPmFMH93fUwwZWscbiJKFr
FbMifw3nLxqC7ZGWMLsOr8MVmsNFkc3X3OX97tadhmlGKX4Al3a9aMYfPq4DWXQvTLmJkDPREIlr
sWySc08Z3EU57dMz8fZhmpQlSojWbBgv5QoAlHrebf0P+p+ZVExo6u3FgkSdZ/aQC9rSnu1aEAUx
YmOlQsOb8SNfL2YqxJ60hovqLjxhxoGttumaAk9zKQxuv2BYQBUaFG0Z7z5J3+vc4dcc9NI9YIEF
U4TUhN3/wEdrnBn+hWaILEs7hW0tCw0+perhr0J3gHJWXteDZBjhYqm2KvvLoEBw8fNdyQ8Ik3vg
6B2V+prK6Hg1INSWgx2v6pWorVmte8BX36COu9lt2ktRrpD6FLmm0Jk8t+OdfveyLo8mTPOUDxC5
kebtkwR4ZkU/tCpzNj6dpuI8NAZ6l7opQugRsJ5mVq4h1py7/n5JwPWZKBAOnMgrNh9SJS06yQxh
Sw1UhWE/r3/cNGC2TKv/qDlQW9UbkE7Rm1eY56Zx2wfOSVLJMlY6jQmSXgwJ3rjKa9jmh8BR2+HV
JvASOVXv6E3ualRM09IQDA8J+8/TUgnwJ7Gf9pHchd+8Hjyp7mbla0buUZ1oNLhk0COtKtEcxPJq
fYqREnYb/HfmPSq+HrQIg/3U0w5vuLw01WEBPWdPWoxBxtSyz7F5Oth250heNuxNv/j3GGZlpbVE
DAt4W/nGUEUuM9xKBYi5q/Pdq668aAkYSu6kTdc2qHlmMWbSW3FTl4GyOKKByNaEVYOKlmB7k18D
wiHVTewJUe07bdU5xLGXhAr/EBMap01H9QBBByU7GLStLvLdHTNkNwNeBKmEbT8P5NxfRku41W5f
VXW/BasRlUsHiM0t8ub1ajla97y9sJQeD1zFejmuX3dR65Xv1I4mz8bMG0HIxiD6xTZCaMKAtDEL
lGqQd+I6yo09r1HzdeOpWg5+PV9YIShIGA7gg1ikvUXZDtixE8zFuRbF7jz8S3hcPdqmHffqNwqC
HtuFX1tHF6e99SOAcARQLd+2NHV3Nfr123ZEF2cXfrsM03QPeLMdBHzTRMG73fyx0eLztDla0GNA
o9737hlVIBSvPOfkOlTREP+a9fMgRm4rovSOaZ9VqDTJfPLuuiFmp5U7DOKizVJ1jHDTUIOAGUqe
Od8hnk4x5v+W0f4kzcEU8cw0U5hWOF+GWfUud8RB/sjhUfVKlw2zBEVa0h8GV4raJpxGBvzjBW1j
BXY5QIIyYg3a8NHD1oX21GEINZHzYDb7wN99UjpmGdACs5NcgVcApnCfIZsKbMLdJewdmRnO8H91
i8A6u556ERTbhX644sB5ykMPsXrRV+LA544wif6wO20b+Vtn6yqpvtkEliu4o38iDDRnRKE8XrS4
Cg6YnOY2fpC7CYIem8Y/LC3uRjBgUAAp9yHfsB45PCzvKN9dOheL98qNY0zY3w4PB1g9km/7Ri5A
yX8dfDBDf3nFGYcIS4wRIwToRS/wu4L4NCGiLWe8yNapDSfwXjRvhBQ+ygfwjEXQ4kycmT3KvgCc
wttXJAy7/e8UTn0FfjNdG6VtTuzYPzeWxaJBuSEX4NhXbjNtH4lHnyo47V0FNU5/R/woLfRqiiAD
YMcF4InumOXMoEtweOi4A4NuJyM7OD91HA1jB2rmjKzGzt9BWgzEV4ypr/50AFheRM5x8+HtlTWp
SzK3VH6iUkJXPY4gJbk1cQ2CHMcf9D7tE1JtP5IyNYM4NWyT1nbGzspwkcZdmoHCWQm61tpQ0Eh+
yIs7SuSBlWBMS/tt/r/gKtI88XiZ4TFfNQlaXYKTrhdQ8kuFyabxb6CoES6v26W5CucrsKr2L/3a
cYQfS6k2p1GkFa5gBASOjdzeU/WWbOMGHSr2V9mpwJXVZJo4KkBrnumn9bFhYlBLdIvPg2NRhq0w
HcP7T9PLWEpXXxRJ0qin0S2EbgZ3XGZawUOAbsIPxL67IzHslI55aCK6vVYFyNLMC+qndx33yfoR
R4ZlWzyHdvT0On0I08ZGoatGeGbzR3bloGhwqYwQnDEyAfNoCeZQFEg0TxOrQ90VGgXp7YfVWrZn
7I0iK0wBMhHaaQlz7OkO+e0P8kWqARZCoZbSQ+9rPJHYnA0RzgSxDkz+IcgcMF56HO8Q/GPucw+Y
g8SM8QhqNKFe5loHOzacQL/1V8MLqGSIEnFhjXaArnM8nX5I684Dz7uxCu11TN30PVA4slPtGjE4
DWw8l81aeopp5wc60YXYoXr4qTkgZT0w+Ay+YXZcUgbfjeHLbsfkF2YCnpOxg5tG5AhI0zffYGIi
jn8uwWYNwNZE3ECoJWnAtBmoa64B01CnlGBVj81bOewa1GHeEt9KyyNxwuxaQIbk2NuiNuet9XL1
nimoHw5Qu3ZWblaqZKho3FRvEPKue6spdBhkl7FMtXdsmjQoqEavTv+RvdpRBSueA1nMrZa8Kfjd
bAa1hFsRqQk0pxTPExdAnrDxl1vjUk5/VfTKEb7O8TbDGEoILK4lA0syE1A+KuA5m2QcTFFSJmIV
Msu3bqG7LMudC2ZuGlIJZtWb6RuVJTUYmo+MgVAxkdt2KgGHvoYQMiIl125PesXv70GtfJ1qUxEu
g33B+Rt5wbQJ4cKjFekzjokQdmzez2Hkbe17xKNgRZ0CHdjEzvBYm7kx9hCl7Q76OcMrRjM88zYZ
jLJf4f1p3M4xv1JqE23RqqagJRBTmwpr0S9ZyRlC/Vd1T6Eie3htA1RAvXJ/Qx/kB0FR3kDuHtFO
k62/uT5lBzLLC2q5grSL170Wlx2f3J3mXIzZcobTCNQN4VNMcUXFoxlD/8uHCo/705SppKCTlqXQ
5XnlkrxzYPx0oPB6LphdDj4qyV9zSuqqPUbMIbO3nhn3YwmZaacFt61+iySp/D045k5XSjeKoH9V
kXK1yA37VcrF8hluSdsx9TOLum1vzdzjC/Q4zagZVVxyHBL2mplP+tjWMy/PczZKmTLIp6e7hr0G
A+vP0sSMvvNGhievPagJLwqHcq6ZD4qum/WCCv9GKI8jCVNBpfprt808wuNpgv1/QpBsUGUfNnZ3
AaIWg0qxSX1mwsduCmv3T4iNrJDutqPZN0a97l3GqsAOZDRHWwOfkH7XsGj5AqrFAtOsQ1C4CGlE
5wUFyb0wSewmWTi0tUTHlOlZSKptkQ13sNhloc4ojHbnGZk5d0YHgxwSAhooaPnL57uMzgKwCQiZ
7LEhTRxFX6P7WiqsJIquEA9WUySAhPA4Vh4XME0Io0qlA6Ag4hV6HhXRKLgB6nh0YcppL/+oORx/
r8bIXNnyMA1NZL/TG2gNkfxzWUbd42yiDhSggKccI+FjPUZKpwXMjgc64bQt7nagJA8AWV8yCrGn
4tcK0SQ5HDNe/K5zNhkyWYxAlYs4D4UoIRb6GPzvdkA7K352KiDSRygnCmv56Wkl6CUYEKE2P0iV
lmvjHQPx8FcDQj/5SKrktijUs2L0IpwPTTpZ/dPVxCgxayXTHunnpIZHfavT/tvU8GoLOIEtBu+r
7TC4Rym/BLzNpSE795Um4a7RX4vYRIjw9RE/RS8KcggEIKLthfoIZE4FalRcmA5i8r3mYjWdvjp1
uzKPoXwG8ahhTCnxVZxngFpiXx2ICHGpM3xJ00CB5pPS0rjyHfMBVY+RJ24CB5rvSP9LT2uLEEdj
6/RWKrLFhKvway4DnqvXaCHeeMkgvRYaWUx6eoMNX097ayIOgMynRMBAGA/pY31PN+nZduzSJ3SD
vXPuz9RMS+S9Fz+niU+/Jpyqmihy80Bx3tWt47uRMIU6n3ED6oIWeS5+qJyXGa0LZ3bKj9HD4xaX
ewSGtnKslAxHO89gL0ZAkTIwRoEvXL9FPLd4zGbzv0Aaj6ElxQst10iTyoMAqhTl4UvHBjkNGbhk
EtAK3l9UTVGaoipYzBC1TNrzzTE41T/BjQ/7psqz7+ic8H8l7SSjss6R+zs6aXcBROmhTOJIVfW3
tnnnJNXgnKu4Je9b+PQndnr9izm99wsNMc5teSpYYLvE22S4bLYXsMFF3BCigfYlba6kB8RHsJqt
zZXCpC7oAE1EjRqQrJowJJNvLz+ROxUqI4tZ47gohgJnSI4KERDTSjvUx9NFNMXhE10XmJqz6Rvn
ECde5wk25KjSPreMy0WTO4+z6neo1xl5rhDgUqA5tt8EaxupWeLerb3VmAbZEFqDqfXm1dtlBwku
P1dt6n6mNZYf4sicS/3rDolfz18+n6LWBbhca4TTYBpydJz7dTUhCKRDDA9D+tPspiysCXqqDmKY
wgXkCkhZDd4WFI6Q5iTGQQsom8DXZTPHx3+/Bn2CeEAJX9tI5VA+8zB+WIxakgyZ+ZHXXprnvwBd
lrprEnYw4kKZ1rht7J+4p6+u+WFg2lCHCEcMf+/BXKY/7xguarV6UyPjdiTBfZWVRFsESSvkGWI6
4FCL00Rnr16dLnOqbb6PHv/gBG/0e/ui9EoLKCZx3nCZ8PNWE2j4avTrPt4EdiVhk9eT+dxC9meQ
OLydPArBNaNcEuxNuj/3vsYK7qNFP2hGm9GvV48PRVF20MhFa8ftw6Uksg2gi4b07MpZCYBD4/tL
61sERec0hkJ/ZXDoUgl52NaqALsQBYui6GaI15scwW9wP1yeZjE5WNk0DbgxaVRF/0APE7Ja62Tp
1eYbIoo8XtcV4iaEvVwMyebynXGM9CiDGhp2Rzw+OS8SiPpYcjijQHUS9qkFSkELI1C//ueFbolK
K1lxsEuhdbjMjZ07KwpSYAm7Hod9QzcWjyRIRrdyPWpfiFZss9eeszlid78k+8Mf4bRx2bSoDY22
4pyFXDFfnH459wsRPwa6fZpZy1jgVQImE1mssq7j6jHtcnufiftnQKMAs8esruVfpcBWKocsCpfp
8/GRmtbZjtUF4BEj0Ys09fNbIAgObAbY/YsSFjKK2/aiGsP+5FMXPzKA0e5NJVxIYyeNWZ42oE3B
rCTGlA8ZWWaLB+Qt81m6xOmvJXYAg12BBFRcayNKzuhjWoMo6Wjk91MTqXj4/5irAdnKCPTN+KGZ
wLOrDY0dge18MAp9NeJ17zwFXiFQgGJZNHysVoRGBboNrz9bN2uQS0tFobdy1rxQfGAqUUvBxDbF
QaklgS01HOBVBnxtRFk5UnJOUk/ytqI4KwwZGOEYL8TE79o1B3f1nWFpOMl4X/Re8ejZ/opHXHCn
y3KHiLGICvyqOogYzmKLvimsfapHJeZ0bui9dSGJYaKd8b9AV1bYiIyWh5lG+eyZLZbBL0Ej8aCB
Nu2iAhyVyPWRaMRy1zc8Kxhwh4OKE61cSrSfDBctAb7SFMJw8QKcRHZs9vhXRFuq+MMJWJ1sH8An
gxln/wrUyJbb0mg9Uf/0GDfm+i2DAfF/x4mwIgDQVne44liaetKyZ2K7jCUS03rmMXR/4osZrwvY
In6UABMH7fUKHi5VO63W7moY7XTX3vhmJK0t/XggbLG1AuWUgqzoXxr3XoykOwSqXWtkPJvO/kRi
HDa1ZA5jxmzb146E1hTbJy5R5qbCjhWvUUlNnXAp9VVAODvGcZsi/gDsaO0QpmQRTtsFz7NS/ybD
KMTeCFM2R9yMccp3iB+s0QkO78CWt/SKT5jsMrhFGA+E8lrGrWAtgUGWIr25p6VmsvjIswOODW/I
bECMn39XaHrNb0ceE67fzISjA8Guxruizdj8E8ftmg4Sczxv7UggmiyK1zEi1Shpns+JB1iCj2uk
2YnzYhL0ALNU6cAIhgDUmrxrmkRuW/Nc0nRsz4nRtIFaDCjz3uKMgE0oS4bWav/DlYywxSHigK/o
ldC4MVdDZxgg8RowMB+VThc6NZiKHI7or9jLyPbDysdhbmzwyMT9bq8uyI8hl/PIMxeYsBha8jCs
A43zFrXwGuH/NMy+XrHSAVEqkc8Etp5j62wk+gAPjUszwHIB22DlLkueUGlmwWH8j8xaRKIS/UAY
U86s0XwQF6X2aYgKurWnHXcTLt7q/XhUD124y/XrO5qBD90d9cXq+eEDGCiz3l+ez9fUsE6WLmYz
5rvcfAGPKSepWvPNnU+F/YyHLXKaxTf19LLDuyOK0M6suwUsH0GpjBoJrBiM7c63wmmnIqJxoBCP
mDk+jl00W1qKCuK7ul3ue98vV6Mg38766OfGR3Sb1e6FLRCyc/oSljNBejew9H2F2QvRlPgGow67
/jrBR1KN3UZKuRY8jUWqYrF1iayn0DTZEViurZ2/Q2OqU6vKRCz34XqqtGUoG+5qaiLFldSF3BHe
eVlwoKcys9WX+Qt1rHpVSWxvR6oatm5HNv08mrn7/dMZXsXwBXymdmcSH3AVeic7psuZTrk/cmZr
KLc7V6TSOKUMynJ8mwz4CCtkVnoPaHpCQtbxRgKh0EXycZHWdU9uMkXNAEHE+8pBoRXoT6FzSMYR
gH0BT58U+kVGNCQIJpsynvoeP23KhtDrTcLa492PJ5qhP8+cUNOQ3AIWWJAqlkIlbWodvMNgLRGS
kEhgjNKGo+ZrWxt8Q/8w3wTvA42M/GXQZyC47u9qQMohJMKMrNxhQPIchtpLqJrqMurrWg1ZS3Gu
Y22x8F3gMAas0dIRKRxbm7I9PVLKxAHM507Ad2FXd6QHG+lV5SY8YHlqe516PMsjOd0XLZZIuhvA
IW8g/9XQfxPZdUmew8cslRFvTwpYC8s4/g7PbqZdBoNcLzXY6ce3Ahwfc/kIc9iXXjNULqu/ifL3
JY/N3ps3OAzlRT9jdogye4TKiMME2Hlh126iwKwfL8VuLPLa51ZFhVDFMkP/LWXhSMJeO6J2Py/K
4BeuLpEeuCk0ka0HifDzYuPI6/Bg7/tJ9AuZkXbcb/Edgvz1gcyuw1belDOaJvTfxj2hRjXVSVCm
Gg7sN3MnUG4vdAjQptKR/B+v2MnBrFihfxR5OmL+hy03lxX3MXLxW7tDPw10ovteX3HJgIaa6p9Y
/qR5F80sCLAjpcXSPOkabcGP7iVdmWSaiQJFrInu9XaRSHk1ww6YfPz6IpgNbvkaJLVqxFzczd5g
eKfVsVHEalaX2et+uBw/OBpUEbYkDnwmJgzYQnrfm/lvpzlhfA26Jd6t4DZNXMf2k0kr1RjcBIhk
tiLBg3hYX251samoFC+Cg3zq8Oe8Mqi3DXLpwb5VALnswmGt6yWToOfP7PDx7vZKfHx93vLEnt44
Uj9cUhs7liUinHmbv82dWuFwrybeo2DNiJVLQGxupJwT3dZW0BIv/H4OA4rEg8cd/oVsccPSqx5R
q8rqD0UjNNiZpqtN7/TxlM/cbsCoqQiUuLquAjH6Q77f13r0yOecJTcQts2R8Ke3oq0bvn5+6eK0
fG0DdzWeQcltKAhSYWeXWDciDwvqqfiI7uBxVXFPVBCGSTX1H3+P8vQKyd78MZ1ToH9S2vYXLqAy
fhA5ZPS3JLBIVIOLgk9mSU2I66iFnAg8+XVkxEADy+ypz3G1fSylqAWgZ91slP5/sVy80oFF8kbH
eSYEFBuXxt3cWuHu1MBEIzaDlrAbYg3NQk01ZZLfLDkbXbsQBkuSnBk7iCpjK5oDextW3piTj1Wa
3dF4zwn7qRhIWex4oY5LcDyjMIghF7dTnadC9kyd8KG6cH+mDuGZo1fwk69NmSRxvuP0laLMIEoc
tjKz7nq8Udaj2s7ShUL64quKG5ttMFBSQV45ThLjr1kZKiHo9OXXmjvVVuFI1Uw8T0wtF+jC42az
AAh483IA71JaQKL8wX26vWP4O9L1Tiu1bWLvXPYKYA40SzRxcpVr3El7Za2sUUlQ9n+lirsrrN+1
d//uJDkH1NQK2aGe5yWbkTy3y+dGewli1laBVNO76AYj5zmSufkO7/+Dkob45vGGd+eJAb0aQ32N
ebBKSgjBRFCFw+hGlKrl1yGGmRhhFYXACdTYtkcm7ipSO93LKfJzl+fUm3C9AoAviIbFOVYB1AFz
DYfYuFaYcMWebBMwATlTqe5tECftuVLCqC9NbENIM3MhiR7Z7s8M+pSPc2HdC+LiQpc03CZL8Mxn
j7g7Drh9DHZrpPpqHu84cUphpsp6i2bVVFC9FQjP7P8bzYsQUEAyB26J8rknv61xgmbrSGRzTPSR
GAez/CXOmvBvo1VQVmYssMGW3mpjdtKUk0RDMXf7JI22Qt0g/9PT4fvchI/W5gmGRQu6+cbaNVfK
KRutrBlU9AGv0nGrUz47rsIfXRaYN9ButyxAuQRxnUWUZiY0JfVUvcjVI5p5D3yXHWGQfbc9G+Wf
1ZHPUDSUf/jahf0g/tpSzkaDgNUzrThWqw4vgitJ+DZH28LDzsWOQ91S4ob2dWo5d/84qlxjoNEL
vRUzjDDFWbN1/+oIIrbdtG+AwM71AZ3C/0IKOCPctpR2E2ZAP8TDqw28xIod5gVNYZXOdhCDWSyA
qcPTZrVyvJZhsjSVQTFe8uKj29GL2IqnCEh+dE4ynAjOm94hmgDReItvyVHeFeJQuf/y5qhbZTze
agfYZ3woeeT+hoox7A4rJAGMUTENkH43gmyZNC45KUgPtDz/rmvI7XKdmb6vhJq2SZr6QljDhnnl
zbB5itOT8oh3qQqUoX4nCJc+xjBZKM2ko+wIOd9Hmfns9EoeN6CUif78CiCdmFU1akCeKcJHcobg
Qm3I2+D5hj9CEvAoQH1JfSYrTwzeAKPr+zwwVPxOshbxRgCAlKXQKFa21zUe+Ek3qCBfhFKdq39N
YisoaP1rKLI2Hm0iCh5u9oT0K2iVszrJp+FPCJeXn+x7XVo+bFqNQrBZzgoJep5xf9HBN6gYiqGc
ZtR4GPWmEAEXtSSHOatUbA7gdtAlhGtnXoGmlAPCmMo253mDAaCXCsfO5VV20EcfwUgSWuUR0B3v
YMkORGGxmmV5Bc0vNjs0lPxK8Dq81e85Tt4GZP15CyKo+NCgW3KsXb27BbYgofoJm8Fcc8bdHexU
CaVLmTMGpD0+FyYxCM7IdG1gRRJzpJ4QqDri6nfxueF0ekHiWM1T1CUbRQi1Kt8NDfdvTyXbWYsx
rsP/uyCVQQMQVuikyPIzsZPvSMcKK+LoohWUabnKkFfNvkEJBBSAmGHMkqbmx0W4OVpwHEAQMvFV
VvWbEJY8ZnEE+NMEKrE9IovbDoMPcEfeCFYX92HqBx4pknhcu1GE/eDr+F7sF7EjtbWFj3OnfUW4
EQN/Z84eH8+prUg5dJU/TMeTAaEXJf89/RVwlK1X6f+QfHA5isQ7tkizn7ZB+g2rCicorsag8jhU
kTvcFMTqMdL+5OpB1kMJZipW9MLlDY1wNGvPKQAbmFcfPOF27XIel67Uyv1NcyU7KmGsxzYVVYS1
NOq1t38dpd6w381sydurWrxHWFBuAXibz9rLOBObpME35NtrZ/2zodwQgz/SDFAWMUZ1nrwba5jL
BsRogW/Mab17aSmz2Y/wDC3hmvtTV5nK1Fim0M6/rAnoe/AiyfEuaQ4lSNLExZByFdzvlTM/jI+x
32PF7+n2XRC3vBxgT4vwugnE+uJ40/5UGOJgLTWMTWnqRz4hIZ2OvOoIfTTqBuY++e5QUGUUuGXy
4/80Lwfp3VOLnuYwrTSkNrTJuWgqMb8xdHNc7rCaWSbS2gcqZyqPWom2CCkgnpAy2/qM6K1ECklF
AfubanFfxssBp+8w+3xIQmzcNwLo7isuPexW04MMKAe/916bz6rd2nZy0hIUDRqF+tFLpu8uKxPG
QcEi5V3sXZ9wigq8AYjpNtMhiilS0saHQ4vFkbIJxTXsakCnjSw1CjMe6HTO3wM3WHO1pw6qxJ7z
mg9d45wqP3MVKj7fZp6S+y5k2oVY50Gp2AEbik4ceGl75jGd5ZO72zjVrw1f7pPh2Ht0U3Mcx3v1
uHAC9D6bnsfRT+M+9Z90k9kxY1Q/nBCbNyUs/pp+SiO11r0idu1efCnytl/nupduITctoue9M4EO
sTtkZQLc7+31R12byjV6veRBU8qlyvtx+Sqehrbe3E9r8aAcJ/d2dK5Ceb6KyEsJ/RYapfejIlHA
zs/paUkSqQIkGdH1UH8ZGYoCA0SXtIQcW4SXprxovLdUbIo53WJDvI+AMRwzzfBQIBmaKSiM0NNW
HBph0+hHr/vTF+q4YdHJqYLnuf3ysMlP9ZD+6cF31ja7E/tkDE1p/BuGaOiYyFU1feJxNKt2Fp+E
VprZmmujFcLjW7I32MNFjIg2tHz226tTDiacjXaf7eY2X8Wud8IJkMCKpoCNCGyrHkNlisMeXfi3
PMOSiIYo4JZu4vKv8ejatBNlqmmbE6fDbKw22OtuMXI+XvZSO7I8x9QLRTTRXqraKwdGd30s7hs2
5xnSPQSW7iPdOL7RbD7pbvL5++qkF8MEsVdawzva8Nh7B0UyFqONCrFsjfMDWfZDO9JpM6o7IHaY
grEjFA9/x6FZ4jzu1o4yqVCLAGWvnFVhZFHihesUADUokmU7dgW76A42LbwSP/33vvFVCvK4+DSb
HV053LfrerewgwiNPTo9CeB3xGIytlfqD+KOPllG2JimUCIJLm5xQd/YBAqLKVoSuhUDbTeEWF6E
dh6lsSGkeYnoPfFv1AJ50YkqFl9hBeGUEcTl8k6hvlB0KfC45JliATHbWn1BKf2V0pkDHSmmzv4o
2eIyF53Ixu71u+XlUv2DuH/mAien5ojwyhLGCVBUUd4JLxP3Wd8iSVWolIiwaQY+Z7sVbkYgT1oy
b9osLI5qqAivmW4RdUfjtM7dHwlYQwOAo0QpWVFf7myjYGLhvSbidUPbMYGQ1Ci+xGgSCTt1i9pc
tqLMvb+t9e7qJsMWnszgHOfVilMICsp86TePB9N8WrofswhM7Ypf+IGlY+DqZydWn1n3tPQGyet3
2XF95EoJqzwMqKtB2tg4hi7PBlCkJEgk9zUI9kIf0vmyNtIqobjVfYBJ4X6RwIrLgQkUoFo9hXZz
v7bKOMKfagpAyVGfzDUcP2h/nqiWt/xpx5mJAJm+64cfcKdVfpZa3+XMScckE/AR2vbypoNqLR9M
plRZ93RGLEetu/jIZZ1D2I4fleVVCgSGYOXPH/VjYsBbBtx7453goCMBwPHm1i0JUMI4B76zwlKH
p3abZUNin8kmzmwtM77BYKj2qE8E1vmRH8mVa2AnV/Saj0FZFjFZz736IyRpymm/VqmuLlaMGJz/
2Zsa0GaW0bd21ugkx1zPrp40XaMnWhf+a16gTgNImxhmhiledbXwGsDPjcY2HtkYA61JXtjqgUN9
bW1lnetCLznzi51SKmSFs7lQ5QO8ovo1D0DsxnA3qRbBnw3CFx4GO/Leav6sWfza8qDC8BlCk4+O
gCj6TJSVZzs780PDzBm14enEptEFeCLxrREi9q2LOHmq6MVV5U7rqEH/rNZgNyT4MBjNGze/TO4M
leb8js3eZYHcD+cUG7K+yuQAc+WPm8jU7HElYFrvtPU4moMnQhutcwEXJLxUBHe09QMXGrpWnYJf
yWTNUvc1zdcafA0bumnLv7XtbtTC4mlivnSQjgPkorOYWWiEWzoZAzJOaNAOyDxflGCVTzKW+l3x
OklnSb9c+puNgX/POtnwA3QrKmQpSopN3EmXILECybIUMfHRQ2Y1xa16w2yjXtM97bFHg+hDrjj+
8r27SvjQvJOa6EBxLKs+LyRNux6YPLepR3W+aUoW1uyeYZCy3rl9xtMHLZhgss1+MMQXL1obdR23
TDZRPV5Mp/jzoYyDHwHl/p7v2YABub3eMnXma7ljHCT76IL+YwjzPcsxJjdXZxoXCXkJHdFN5uWq
K6IFaJvEiwU+0fya9VxVqEQkmlllrk1k52djILP916QnYbYlq8kJmFky6eVwLmlx63M8IhBgBkek
/3TZrFBqfT7lvAH/xzV3zlYGAO+GEnfNV1ZbIBKA0OZEqVPJU9UOocemCjv9Pt23jQ7rq0P415db
qEu7WFwIVPs0Lfvf5aqHAkTAKf+6We0kQE65R+uJThR4ga4P8UxeBehUSYBNTIi11SF7o2ZxxPNp
dPjgnFa+kBhDPUgbbDrbGi4OfkTbek/QybMhJb+8abnMSWltKp3KTLPawEoNyan3NYH01UdVYZna
69biC3IpQOvSHVrq2a/9rWhleBYXueBbamBpHqqmY4GFppSJAyvDUPImx8oYLb6FwcL+zGHPn2/3
QDOkr7QPdFcma5Hwq4WBF34em0HySYE3nxHT5W+lYgl0HjVl1FmPgiCLyFQM3Po1eFR5oewuM/wS
qYlve0IFSEuQcs4HPEFQAUwU4K1ox/MdEgZhzialU5oHSr+KhuRqv0tWp1096zCdxR5aH1NBHLLQ
hZPabuVzZWxJjCMiHlkh87EOBiKc1MJh+J0tr09Zt+7UFUc2HQH6UNUWzp/GzoAZGGC+z/FMYTG1
48CWdRd5rPJKJm9aJNF5dSd4yZE5cxPqo/VeCLCR/zsW6COs1Js/0hmo4IptV7e7Nm0C6+6ZTeiW
BT+BaS7LcsEX6Gogjrld0928SKoowvJ2yGZuxnZzWAsKhkPlIfcT74npf9mdWimkXKxk2Y70VPrH
dHVvXAWRogiS7fbR2vJ+kWsuyOPsg83gK8fJiehp7NpV6i4Ptsg6gRrJQbMKxCXcjtquLsQpPDbI
305Yx33l4dSplXdQ1Unic233dtISiR6jNBdi9z5wLv3EuKUcNCdj6rrAFbac4WwvPsckSEfgLQRZ
aVMPMsGk0Xj0qkfdCCjUAzLzPiUhSLgWUvwiWGelnbmXQORPv2yX7gR+IVHejUSZQV1Qxo/VHSBK
DRigBSVwD4FSZc9Eh88JJrUFq9tHELwK9w34P+rlu0r/MYDdjdTL5qzAzqjBHptMRzj/AwJcJJPg
pVuXrfHfgdbamVJ2+n1ctjdAAXG7rkimhjOvmFc1Pq1hPz9zLTcb5D0oyCrwV0/qhGLAnIqYxfZY
4aQq0ayqKqYKgHKboHD+LAcp/j5IXYwK6YhLLbg1qaLcMHLC9CA+rveTxegScUCAEtvGktocvvlC
G698+WLaavdBk8OEM0/BnG74vhuh46B8s6WRT2iTzOXzJoTyT9pBT2cV49YY5Y7OJrVxdj/r2Az3
mTVQwpOLlCWzC7jOfsdokdQHyWujThRRuW3a+EscDvRAzmAOwQPy6VS9/bIVD2ATygQx0gAQ7rmL
gyV91h/we2K1xi7iEK+wJcy98Y8COYpZCFF1wLDrPEKY8jErjs7cQ8KYb13jk3nu3hc8Z4CyYIgm
BiFvd6pA3EpcO/tVirNRnUXY/izl2bNyRHQHttcxy0A/7ce3aUMEnjPlzv4CVATgfuouGfju5Ezb
uWSE7z1HCIWr0+In99lr1kO9VS2VzEtlVjj1+GkTJjzzGazWKb4srVft60HavIgbP16OeuT2xBAf
ubdYTPtt3fhygEIqz8YNkP+kjFMne4RyNqmN7J2XdK8yd3gbnz1L0C/+B/XHDISyiAwNyspSe4+P
3OM+JuwUb9dzx9IoFKyr9Re9yVMEnzclhANpL9f1GrS55Hh1YmXVIIcOZZ4gmgTz/fMaW8CoA/6l
99nW3Y88X5IC05E+Jv4sqLWgzt5j/EMIbm+WsEBA9cj1KwCzDs65JL47deehy+WGUCJI/180wsbo
dZZ1xPOSTcIgOIXQfTnWNH2XNMj/rwTXKxsus/7UTyl7bKjfhufBICb9OXlWeLWNNJo33e1JEcjL
mGROaM22wq4ndsB3UNkXVFw7oi009HJvWLM2rgvMrcFJ9fu8F/DDDnH2e4Z/BDLiPc3JZ2TBFUYE
Ll2K77PkgoQ/E2P82KibJI8lqjUqAf0YRVeqJrHG9SvrTR0ZmvwLTaw52r4KFeHKo5D8YcfK2JRn
+nxYaPgip/M0Qh/HHrAN1a6mE07G67Erj6KcrTQQTrr4G8ZThZ0JuswBXXU0hREfkKh+nHHUxfD4
TsqcqELrog5SvuwrSynSGEwX5HPd6hcqH3bn9kq2UqkLO948FK2YtZSvesLI3XV8V0ciDCFWUT4r
S2rX2Dn7y1gFBT5ipvgYaWv6GXXiHkRy4gDCSvGt8HazRCrsqD5hchj6uIi9FU1O6DMFF6ytL7LD
kHp+cTIN0h27+j/zwtsXfxULCbUkCPuf/LoE69bROp8YDGuYgmYPBTbWRzvA3lD1DtBYRQVHCFqM
zolvNlRV2ChRhd/jcBHm0OY9OvzQc/XL6dfuLVcSbLAqdyrFhA3aIheSLEn0idWOlWGDRunUadFN
ej+baNaox6GIVKM/AMZmJ1DGbObH8s0IKGqAnzABjDRIk/lLa4tZyvm7n3E9HwMVOtTSfrcs9jH9
y19DBrHHJuZTZxowng7jyV6JB/M7ByyAHNuFk9UfEDxq8z8VAcNbsIbAj1cbGMskOinFb1pa1hyK
3XH2eoI4/MxadCTRvdbKKh7ITSKz3m2iin8ZJHEraiiMleucJk+qLswHq22617Q+LDB03EY/0hYy
CE1IquNdCl9uC3bhgNqzwLEdPpquWDzXVUqauT1dJY8MhoKp2V3qIOp1zbTOWQU7VTnVh4Y4j6w5
jv9btdHaMAbdko92B3ud5+yI09p8qewBerUoKslCbp0InWvCxe4GwWqPmY7RiVwOpc9c67bzribY
uRRCjew3SuKmqiRJJBejR8e0yUBlsJSk0Y2nXBGCTy/CfNwofdh1gaRJC6nQgbNd53akU7/GhhjR
vfkLfHwuw67t5/V24T77+1kEZrqk3JJoNLJQKh4CsPomZXzxpsTkGPfcOUhn3fBcmWxCcwlFAmqq
W8cLd93kMzc39uDxgGYHwKQ8CPqjnyDyjESR7M5QxJTbSNEACzew3NnNuq2wt+FQq2PNVjzH7X0I
CnPYnUsndNi/bUHqBSHV0R+fZ2SJWQLSnr3oJsLjp2XWG3I4Cmb/DNnOG4esmatEqTriXcguNQT2
qA9yNZLTXt5Vpo1ACqXlFlbm8aaRTz/+isVMZvIbezD7PGL7h8Fljm674AciORt3+dNUALC+i7Ff
6fcNfKRB9jOEn/KgZemwBfeBGu/8yRMAazynRtu1fzOPn6bFFRKo/mMTSr+8poYPkk5y2hQcIf+r
96oX10ixOamo4/dt2eoDiqEewswHFVvyzUSJood9k+8lvjM+n7Q7cDXZReaIoGQsuuRg96XHT6AR
kRyfRoRlg3h0eMAuPE6c1imL0Df0PxPLmreFEo4PEXtpasLuK1TIZ914eiOiEFTfSZwJf1NTYP4K
eQ30B/EwFHSDAcXfm8FIQ0x6KfiRAkWpvlTpkHqcs5NLnOwBJpK7YNsF/LhNCwT+VfYxxbXf+EuA
iwEnM4FyxyBPJmAABvWnQqR6i1e0egZMF8QNbNfPJvHtZuxgBRJr36cqCoefIzK4pLNacUaHgUkb
+4jwRgfJaNZv8oZzdj9MDdNyv66HHpjW7DZR9FsOnSgs55rehr1O0zsS2UYgHdsEXhZ0sh87U+Mu
e+cO81fnWLIKbGBEsaQks5fWPrYPsNFs99FhTdSAZ9jnnRDsqNWkpMCOXnTH49Hv2WgsyuFn+kdc
p+j1CPmhvZ0onBvZ3VKBwLRHJNONBEfJG6/HfqlhjKwMWEHt0/vJiVh0VhKareqWj772QTlJw2TQ
BjTt71jZc8y9s7zqfGBhMb+f98WH9tWWsAKihFPCeVada2ncw0zJmaeRDhYBwT+z3oT0lFcdnCET
nJNPJPJHngTvMvXt/81x4YbufgbGe/p+smcbm2DWo2zE4BXs82L1/eEgP+THZvjk9C67ssHrLru8
1tNjf+q6YtXpPIGDu4o82KsGed825IYfTXRoLbGvEVl63Ol/86qYOOuHHLDhPN5pHdA8yEfJrGpW
yXvcSo9vvq35PiJCdD+D3hOjOd5TqTkcQpZCLhocu5yCA+lU4SfwdPDqpAZ2cSzmbJw2N0GDIa3g
ZPmwlz54wi0uRSD2kN9MehT98TMN4FPvnkywX9EEcZrWGD89V8mM5ff9OhoG2IY868+9E7EKt0gb
bcFeh07m0C+WY9x5th8VMaAh9Fg0NPEDg1M1jHdmRjIvFOctmWNZE+irmjT2sVOBW0LkQWxpBeiV
HM7WsLDBFZplb4ozaDarUVy6Tzind6rnM0148tjuTQQlNnNdh85T6scM1s8pSAJHpDe2QPFNn6KX
Z3oMvdibuFpd7V36hXfGI0jdh8UIj8bY87Ws3ubss1v9Q89MYcREVa0uuyZceHFx8pn3poXtIjym
5fFAqzHsqL/EPwrNB2sjnNwBv+fPsK/AVzdWZbkRimWfMSLCYvnwQUzxjIQBg1GDV+16iWmdbDvo
0kxidhr8VKLssiK17N1JT4YY+N6ioEPaRKbd4DZ4HvkxwhMDOBVF1B1kcDOJ2rrARNEsDgacLhCe
Cz+bjNpLpPFT9MlLJTXexnisI6Jl5lbc1tm+cfsxBOsFiMgN/5KqTVZUHzI+e/WntR9vIEMvHUXo
TFml4RyYTzQfPlFnluo9XFpojDK3FTqXuZuFwrNrxJWoFH7YyqaVCglDWmzeLf52CAuaQ9f65m7P
5lq8SI2Tc1hFexj6yS7JTJ4iMbdUKuzqS2CXDUuEc/FWXM5JZj7XR0TZe6m037To7QXkfRj2ak9z
kGfJVaTU5TtkpDwqE7AW2/zuL8lMnRgAkG/2Lx3KNnV35eJydDuTzdays3EtUlP5/zTJr7l3HJdP
kmp+sky6pk1lJyOA6p3NlK2W70faU3rOa04EH32M2YI/9mPw2UmGU2jfuXiUiWjXWyKqGIN5TAqQ
YPeOD4BSM5V4W1z7B5pYpyrq9iDJRNlh1XmVpRcSsFDr0LNpcO0MPctZuBccxIJBHpRY4JXRsjD/
SqTUPQdMRQNCU12SFlUmijFDkWoedCnMFL2Rk5WBcVQmcZG+Obg6WWWypE81gLPN0wiW2C4OertG
uhZylOPm1Vl+qu0a+mmc8nkeI5IvPHCWpSNbI8KGUg1B9z91RDNWkpk9eoRAwsSNXgBWb1Du3tH0
QHaCZaYldk0bUmElryniYVV5Cr10UyRRebgKD3tdag9uUyuVQkQBHnRT13rxg7SIqGkGyKTJ6tMT
8ciU6gnItFrnsw0bexw6Qf+t/HDKSDIXFZEvVDfgzhnatW6G2PYISz3hCQtqfWrjRdCRNgLQm95o
wPV0blEjY3tGdvEDebp9nEoSe4UockYS6wTi4U/0K0kO0w7dIZ2yBjHrPSGL1kblmhAUJnqUD/8f
g18sMweYzud7BFW/yckuK1/p+99nc/xX3+tBPy8IQzdt/28nCG+pkJqQixVz58aSNS6L73m9bLY+
9mOfuydrwsty9/admKzeV5jJUl7phGohDAx0sKyYGy8dws2fCdMRvmaUHj5YA3LwZud90julesYu
b8ecRqy8f32QEeaZ8YuejtHvUMSAFgrTB+2sW95UFz78T3K/Mtf0NBLj8aLG0HstndFoJJbXcMKq
o9B2aGwYyHLUYipFJhIIRGfH+3vHVcrstt6GZdz/xUvss6Sc0CcKodKy7dRv7wPzlaU4OiDDqT9d
9lvw0u3YVlO0+q/zKvOgZeGr6cQoot5GTtmS51c95gT2gbi1PjAHTeVwbvJvbHgGzeeWMpM0jlf9
jq6W7hdz1EpR65AcXtOiqFwVw2hBcXSib1CWvUcMxqRvKUrymRVHly3/KwXZonm/1EH1otN3Tvyf
FetNcqmxLM5LmXw+AzXxqxlVDjKSBJT37FVMVCPd4lYIbXHZGBCMey+miQ2UcKUcyXanzsaoqWuz
tSGA+dOepJpFeCnoIUCVR94W9RRpswiWAf9VYjsfE2JPLjxIsEW+Po2vmM1siwEce+xrWaza/5b2
eSSU3YGEYd/ihGLeftSAqxaG7O93+uGoocnvLwqxxZCbmCCasB/dM6fCmqOKtMSbWM1DuEjAU553
gwJS1iSgoPEKxtjA0RfWQ5LQ1ltBe6J8GS3nkiAKLelGrZFev+KARvvhPS805dGOc8nhk/Xta4ul
P3c6VF57VqJVmUJ1jKcecIgU7n9FOWlXyozAomb4jVAfzbgkwIUmoG/lFZwwWFHW8an8+DluQt/Q
vhCoc99nbHlWwmIl/WB2kj5PDuCnVHk8Iy9Sbjqo8jLboJ2kMN1p+uAQ1iLExmTvx0I/BTBkdxyl
DlYy+zi40CiPAXz7t7qJayQDcnIlguLaOhd2xB8iRpRZPCdax4R9VSNs2D4C45ezQU2B13dngAEU
r/vOuK6DaddTcBWBN/GTvVbzRjy5Z+/QMuMAh2udxqnPhIvy0W2PUc0KBbDuAAgybzlWnr07kqkQ
JzW7miELOwPrjskdluMdvpzoCpVXs5U7D4+W2YxQi3OL1U9XtDgKYTdUyi3rm5NG0yXS9HZyVAKW
dtCJL0nu0EcDTgMIQHBKTDZgyWKYdR4k9KSUd2xydhJlMkzopOazffG/KeqLIJF9iDTSSVt0feEg
RtX2VsIJ4huwu/D/Cg8XpNMenw0nBJhHqyASNHiVBixw2zT+Si8Z2elTr0HmUzFq9vLNtJ81vsQH
t/RpLc6dpU+S0D+1HcfZ9bbDkJY2iwdwxtoMqwFHT04DkH2KbKqmGFr3fBLJtC3MgQNktg+sWz51
0EEsfPr8cKiPKO4BP97uEE9LyRjGazZJuVFzfPOoXFThJQA5XYc/8GoxnEAJghv0tkl8WUX+w0Zx
d7+W0Fa7mTKOyl8rXaiybYzYtat6cDrS3Ffw22Rrb43KFh/Ix9w1uErciaNVfFCeNuoLDQRWXRLi
zsj9ATCLDkYT/8VSCqB5MSTz+SI/U8Jr+9/IW/TmK/v0/r/Ys8fqrX4I/UZcsdgm29o3TEJ52d0E
TIp19GawuCMJqHLUphvclWIEwT4kdqu+jESu9z56Jc+8bKpNS9kC/7wUBav0mP+a5jjNxkpmy90s
F9RDcmf67qlitOhVRcIbpjyECpiIwxNdL2OIoc1SP2DzwGwXilCp3nozTexYIMHhdSJbn5KKQy5a
7U8Tsv2CgggVNxzCsC1lP8CVYduAKxYZugy5D+g9u+uV2GIPpnDImnM4fe0A/TAigXnvISMkFKw8
tBNrwUQp8NjyGQ7+3ARVesClpr/xGgdPw9Hiy0zTQYp2ffS3rTaeDyd2UqaeSTWqrAUR9NA5muP9
psNnJz9c9XZXcJcobmrQkM5j5mvikrJqZLAYw1edIZ6qu0NJOkToRMRYRU7S9G3L7GjKdhkkKI3Z
9iWuLQqtraAXCm19R+G2uWeHApKNhPsO25bLptiihT/+eQwPmVujytWJuTElasBrXYPc1jVwHXzR
aPwt0NUGNodkN/J+ppP626fDu6Xud9xEZ520fC1fylzGwslVy1JFGiw0MACqJgBt6+qP92nx2NcM
62dIziBGOE2OTmsFbvMHone3kyIF5Ze+2iXIX+Ow08jWyumzCVIyzGE5GLpLN/GsiYvjtQRW5Tme
D+x6l9IYX5FVNo7mgRHHKCMw0EhKXYNhF3PshFhNQO4CNkNBeTLEw9DpVxwjRC+75fYcTcs7Kn+B
M9YnufwxB4PRgN3+JxXSbJ1oHt4gZYXb6vEQGCZsm1FfPhJrpDmbv8sA4FpD+vuYmezPG507icJ8
ixLh3Kz5HQUKCYWOLnIYP+9UnwKFbMTcWuaOWA4FihjAF+xA10wpSz4i8RPzT92ETTHDNsx36WHe
Agj9YjeYcYbU8Y1VheVnvqizTgg1NYzIc+X9vz/1DHvxmkCoWWY0IhyVIBHnIJmziLCPDS5ZBq8W
vwg3S5Ix12xO2pUw54G1eXXrdJIT9TR4rTlxeaW6rHeZErRTLjckbRbWvlO11bgMMwPvsAkxb8r3
CqJu8pGM+QdsxHY47NRoLL+ByPb1fsTclPOpBWIh2oF6Ukdf9+Xp0142IM0ytPW4c6AylINvzmWW
o/HHGbcdkEV4U4KZ/RpfxIrgdQBWdX4OVNE/X6vvxxElLu9Pdj5npkxR8MIne3toWS3Oe8lxqArW
o8vn/l0lzjBiOTgsNxP/qme1pUleIhnHeR4WUX6hxGgPeQTHb+LmkdOAfzbdcg2LSRzJ4oa2s440
kDWkp0pkDpfOF8nnQJcnYUT6XcgZJB3iGZ3ReX3Y17KXJCkh7uY+f+mhZI0acxZ4/1s1HTTrjfPn
mboffkLvl27kPYWiTPYbfTq6NbF87ZFVC40/b7FCCI5K5VBGbL9BxluTEWAh/D1qQ8yJMFE7CBno
QR3CJrsISruPMtggSRR2O8/a1UScmlY5nInIFJy1WvCQKIwwoqV2CaXB3Iljj0r8aa7otCTpVfGs
UVDv3kkPOEpK0X/AZHzoE3cYPEg7VQ9UU/Gt0X9yYLnEMeduTjFgClr2Ie2I/sXeDu5hmK1JnRIG
uYEUoFbaw6Wce1akh4Da8Ek3rf+seoWU23L3Vtme69wd0ugmnBKMbGHgVIBxraRmFX3L0YAXyG4k
ZBqMs1Wd67MoITd1StWKiUmDJbLthBCVFkGAHuS+eBCdzkCmP9x0pZlaDfjtXC0zBx8FHGv0axSs
arECLXufv0RZ4yAHnRv1M3bf6jOTUqMYHTdspQ/8SvDn5MD3UpHohEMhJElmpdLVwKf2bmzio0S6
DcAFxzwc0XlBFdmxKmi8dR0VmYbuiyDJD7SP1HKgkahRfFXuCjORDbM9qPkUAbVlc1K/8WTcvd/X
e5abp/G+WMieKZqHhxIMfw0ofULIJ559UWBDIY4wGnnbFz+rqFTF9EuJ/ZDciqHiKEe8+94nt5zf
2FxRINzbpRF+Arzj0wKZtgUCns2yFfCZbzfvLtpXY6rhIwhIRD0oMCICDo98GDqjrCSLhCWozQjG
xrDMCi/Pq8r4JFxBF4cZAq5CZNLmazLS73RHszHF01FaWpbjmQem7bPvvcb7T/R52+R6OjejdDch
YoqLvmqf38tVUKo+4ERy9dZORK+BhkNYxTF6tYKZJXRXQ8TtQKEQJEF7rtvT5ifpiirMpXlS8Vr/
XgcGAcw5U5Inox0QazLCFaz342Z7f33ZQDB81SOk/zmbvaW2WDEvRecMrY4UbSVqdiHQji/nksxA
lGIimuD9oyxr1rmzW5erhG4k34c/+DHq26X6yl+aTHPQJ5jmm2JctjhMLKb1jxVuGiVozBhPqXUQ
0aXUu1FYtYwZorQ4sok3HP+9bbh4RWo3rTiayyrBKbO9z42cdjQxCEK6hL2wImYfq3cVwbuEkHNp
vfRrOh/95CAnnyAzimflzjCt0FUZDTvVJ7s1gvRN4eKnWexvmP83bgEPGTDdOPghi+2CTpCwR8kV
d1H0LGQqIupagIO036dObIkfFAdAHc/lAk360FJ8RjkmAhLSYIMgmrI9LDCnDngN7/Bq6Vn+jL68
0CcEyUPs8tt9fzfP3D4l8kY5vPEWjooSCN8zcDaD3Nw2gxTwU9m2OaeJJMlIZL5eGVM/1GxSzpPS
1TH13zcTaNkZftrS+ohmDzsk1dmCtEoHEv8jFJNpZObdv8K3u3LRRx5244FpKDIikHwXI3JlP45z
bYeLGH7tkre0hHumoA/etKhSSA5R+cZUR8/sUnjjtKoklMXFqvBb+48rkWNARuJAE5HCw+4P+485
vWX3ZAwD5FKWE6l6YOW1zN0pVDsOtaxhuWfpQb9P4mMdoLKC5H5gyV3pDQDHWJkzJfxprrcsXVLp
IXGDXgx6xTtOHMPSy9WueophpKLU3PzxLsSnZ9cDByvo0pq4iJEYrE2sH/g9K6MjNsJSe+IlHQ3w
2VpdNUslaV7QLVCVfLeefJkaUkPHmt4YyuWpId+eqWPpmSJ05hftmRjWUz60raRjCq2ga1yoWcvR
IuzQppK1I2lLN5Zj7cv1wmV4eB7Iq6V8aV9WoSAs3FU51SYWM0r1dB1QfhzVvNrZEct0W2w6uekn
PxTCmE1U95/e4jpBLlOLb3/BlLxMjijjaXaslcJXHzO7dOCBGIxScY9pTXW9YsunCzX/vjEmfyiy
/le6ggogAzauaCI325Yw1Yn5wJsJfnuXA2iUx4b+Hi679j8fKSKeDNitBkerpYbiY2PWDzBkjz8l
FS17YcF6YNvUOdfimP+FLS4t8sY+mxldl5dm9R3L2E6lEGoZNE4g3JGeWTDMysUzJWXd/Z2DOcjG
3HEFUVS9+pI+mHM96rx37R4TRzTBR5AFMQrWyeeTXrEqyAawajD90/11VUF15KOQx4lkje7YFQi0
UjN/J+HzTRWl2SYK7HhGXa9oXSa4KBJ19+XqyryLAz1CVTY560tDVyA376LV2n27wsFX24jWK3kz
u3Be5FE5R4ypAXEB4RMSRvziBCX+SaAQ9WoETbhi9B+609g23IbURSJ2fSG6agjSKFdqmwJDGd2i
Ad/BfKlb7inzij8z1uuE9fsIk5KvVjGiFc7gXI2Q6fNNDkgVP20a0VH3Q57zAT4p6KTsIgy2N/LZ
kkxt/7VGbViDkQB+5Uvqrt0+Q1Qgq8EJAVBhLiHbHnbhSZQacPo2N5deZtf7xRIQCwVz3FDzM2N/
pz5cCUozFrdaOfKGvFeMEytR3fbQmCIOONfAlgDXDRyXW7pfB39FaDZg0f3GNDfsQBK0VvTHzr4+
s4rRBTYQU2Lip4ULmzvO4lF2j399qW5I2ydg8MXGT7CfutWuLqSyhwnpMhoYv2Ids9ndiz1/6F1m
oAXZvwCZNwPl6zdT7pNFfhzt3hMkUqdV/QoAaA1VM3Vo5fNWliYwr1gd/3FJ3yjRuPT+Fvge2hyt
NxQYarJpI9ye4mJaLpeneKik3krbDdFiD5NzMmynx1vrJmgdEYS3+Y7/0Xk55ThJbdGA9ma6P9hZ
stXJdbAVcbyPIwarQomfSE2mpno4TR45dVl+u7la6645HJyfIvAz1Hvzk4QBZ3C9OMPIxLgm5/go
o/3MmEURcYVF8B/KqpjB6tSZ9xBgYLzddou2Jec3CyZxVLstl/DsHn2RJmXtS4rftQRxqW00nB1m
RHhtn/7p33iCxWtC9IS00G9KTCksDIVR+VtYKssPl9bs4LM2JUGJDAYxvOzVxV8emEEm/8zl97z1
ff45bH4ZGzC11ZNbBBcSR/qYIbURF4eM8E3iIh/u1avII9gqjs2hbYEa15yWbd7p4TAILhY8cBBM
5jm+zW88ZAzPN2KpWgPYEXiEdQhgJVWwv02XLI1qPmngKqkqT9P9JFX0t7RANeULgENojvMVmhH2
XSK5bg6c5n76E8KNkBCdQB9bMWkLeqvOon+pIqyO31j5/ExsXqgd9AUDtOwKhAK0dSKTbrvH4tr3
Y8fAEXgzbQ1kQ3+e0M7XmPQ1y0HRAzdn1WmUGIhxdB+3Cky5cizJBZPV8CBc/6PT69J2KVmZpWMC
nd9thiyCmFV6t+bozsnkhPMBJ/Lwil6wCze2J9LHzEGY2crlHs1Kwytu00f0tHI1gYSpuvWlpm/7
nUk3VjcUlVJN4J/Gr2X9hdeRHPm3E/BHsnKl5NcLNHnpNhDsuQ8qEXP+CDM0O/hPZCeGOa9MgR5W
DPHdYMJ3xAfxMoynaM33dr9huqRbkgXq6zTAlZToyGE6Cu36WcdcCi5s/7Aqu3+/nuC+kYPCH9ZZ
goUoWxeueGPIWST1NwKHTZ3lH5mY87fYVvFVF30mEKfXZClQ3aMPGRbsgae+8S9UHXoGWQGqJ1Ti
tt8OMEygeyKUrF92U6bxHwxxjBvoMJMvMDhU+fmekQ1beFYcCACZTiugOi6P04okzcRx9GU2mV0X
xSRNkfv7ZCNYK6cPToL9UyLpRD5YLKJj9RvxNOQ5y8qkAnxTlvAAv9tfdU2MjbLk3TJYpOscdddb
RahU+zqPc/gaInnm+AniKUOnbDYIsLF7qUUppYldrhD0Y6SDpGA8ubbNZtKc8zyodfSBLBi2e4Mj
gAKVrMtMoYMUPZgd58QY0LlfXLRw0Ddeb7h7JVDocubMixR6KIRvXyhLQ2iXd5hHlI6XHPSdNEtV
t+9fvwAw8P582ZxgqiC+Tdfaj82wv44nIuKqBov6fPURpn9yfI2OlqXeSqL7uDDurOwhy8QfjJ+p
6HBhoD6oZUC+Tm8ljSmbnljjMTVASb5MbfaTKYyOHMWAUWzXfRLXiz44wo1bG9caGtHJbB1afNQp
ozi1s9lrtxs3A+Cq652aShlFK1yOFyne3RewNRwNkDw3ALLMFrbdr1vX/BoKHAFhSlgj3CUJNZyi
eBY6F+VrUWvnm5jSdx3uHpKvJo0xTwcKnIoHG6qaxkLtLYVCXuZTWxk0xJh3QpQIKP7J2lfNesDF
CscWyvKfIl6nMRH6vtNT5+nG70R2jx3PIOpnqH6pxRCa1M2twMri622Q3UC6Wz/02rb85xL3Bs83
qDOnJ71Vuv2pebr7KmuNvsLTQnz5q2kxb4mYE7c0h+FZkry8gvtSKmToHRMULuIn3Z6eK4MrODk2
yczCBBByliAsf+eQsYtjJ2JCP+qJSg6fWO0fRN6cX2Y2FClFpc9ac+TSTWBX9M49vuBJq2VYMa2Q
CjTMnlSNzTfHE8q0XwaGGp3KEIQ0F+gR96vlHWVGuhtYgXbYW6Z55wrEQu4hiztEGhRDW2uEJqG2
tWAmJnivhGOSz6ldhz7leBiRAbn3Vqm6U+lQPNow+Ci8ZScWhmdSBeM5OPh+NAyGqjre7+xOng9q
cfDy561dCnsCcHibObllLdSX5nh+ozndum4WKJZPZ95odKAI4BOlQURYkzFYECRMY0WOd7kOXvcN
po3IqSv/kUiACXrB2qVJ/9skikX8vlFqhk/P08SQGiLxf8KxgYuq3mmyftj27srlRQ4wDjMhaPF9
Al61u/eZdrXBFn9TPUTdyrS3ah3+0vsVWy5ptQeMXDbSgY5r4p/vz4CSdCtrFtkPt+A75bSoWJ71
TVJzhkzqH+8HuZG0d/X3DUOEoapzrcT3ICzYvtc9/k+ARNV6B6GZ4QGPP8CnKl75Nsu2w18wuq1Z
AXXAU3CIEfF3AeulZJo8VdwPyHTq+NYJdF1MlkdFo1kQ81u9ibjInjq7Wkabg9fvalDU3IqhCfIG
8YMA+VX65W8yREWprcHzv0ucJyYIpFuSjL6ENzOMNH1DkZHFXk7G99+jHgTx6T4DNui7YQrjxEWL
X9Dsv8j0DEeEsXKiszFAG6cZE2S9kwCwdFqZvY4duWoKxo+yoT9mChhI3BzN0gwyN87BNjt5ElJC
3AG7CmE7CZBzxRHKrknhOLeJECwO315Ye46uZNPk/J4L9xEa+KBAYaTasz/0VxzBp/06mWZ0xHUk
7WbMfqUsIzL5zo0+ZxXRE/Lnqed2MQMFvE1YuE8KCIEA3DyA2eLfklwnRoVH+ZsfhQpVp0w9zwEa
eLbyK0S4sLmtPOu3u/ayJJG2nDjewY5IPQUgFQF39KUJtD3OxgYqQ++pFHW7blXRoWBNxcwCSXk6
XuEz83LzaDb+5iEUymbUStAh7/vz+7oZY2mlATLA3eWht1txjSiRA4hKEPjcAVHchNh77G0EpvwN
Drskv7djIsRDXsxKEbK8DK33xCa4Bso647nFDB4WRK0qBPWAu8fGPiQ2LHfvHlQT8HF8W9+H78SS
8qZGj9Ssh+LfqrC0nj/8Zha/szu95O67bbs4jkCwMEbyhTgLxC2aFNMI/ccbQ4hGLwQORFPBn7bj
b6tY8HqSXgYp2WjhsndVkrCjEH2VcCQOjXX9Uh7SKo2aL5hLj/Lu7/sceguA8R+AZY101oBeTtip
yAoRVFGh1oKkaMB7QUpem2qCuxPIZiRbMN3mIiVK+YEd2us3abQAtEmkEvzUJLFjQMhEFxq2QQEl
RTdwny2mYxg0QfTOEZDbN+3Lr7FBpu6bk6FFxwjN7b5DVLoJWymZX3/8oRqgz/qeiDWmLPN+0Lhk
RX+SmV9Fb7ADtQXYcT2V5qcQMMY+XeZXgMDdy09p3F6bYYvYW5Ge8mKR2hoshL+LoFsOsEec37c0
HoIVxFdHzrP/DNOKlyluVO6H9DrMiRrAd6CHH5iV6JPVtqQf32hq0/91Wt5lVvhqC8iIEblSNy31
Tpy1BghuvhfGPKQbkcqb68QNF2Uw2MIu5aKqTnWbG6i3bK0gCOMicZz/QwM15PG7n9T9pVldhfcz
WrrQQ63XmDGDOlC9Xtere/KJjtrrxr7N0oLm7+/9/ECBEu6vYCbe3V5pY3+cXmzigsnDB63SybEJ
Z+P76a71z68CinXjjmsHSW0kLy2k5LslFF6lflfO1SpdCVPJqwi0FUE0CQukEEbowoyya9TCiQQK
iPM7HgaSzdzWiD8jsZLZUnkQ4ZdEZ6DWVuaTh05yZxLNgL5JliOGsKcwomUwhUzwiHeH9gsD3m+p
d67V6V+X/zEMbAJyD4UODt7fW3YFa2x+BGUVXNXZBTjWOPeJNhKg1C3s4fuAts4plNFMJSe7D8Zo
KzhaWHe2rGUfHiKxIsKaoLOdQrHo+pDUc9LxmTJFO7zFsf7csOIFNaxQ5tO6+d8u7gihiHJCojpM
q6vTFnkKUjRVt7jneBoH3Vnr2Xx/wmDk5OMa81LK8HU09gaZj/Pbl2BNDa8wWRpAr+jh2dVDXpc7
dq5JUaRSSPs5DM90lankkbHPqpI/JVfqzqYrAjz9HMaTwlquZKLxsW7xLWyrCJ2zN4DA2tnaOOiT
M0m6aIZJ1qETes0no/FnYYzPTaviM702SBrsB1/cGDg89gjqVA+kPmhZtPIy882Z+rXhoqfiO53P
Sb9yKK2nBUe81V0DYQ6bfL/lf2ergCS7k5THqFR/7nYXXxaBN9KrjIrq2BD9mNPpTjQfmEME5Q8M
RMq3WWyb+tD45dYo4D/+gvrP5IfJpkoo84PpW+X32rONCdoJf4SjY8MjN4v6u4Db5Yg+Q7AKjRSx
IoEW2oxVcoi0zD6dfGwoJKMIkHob07jz+/0fomqZXeeYYQ9D0TPqx2X1clwFcXU8i5dkq8Vj0WBg
E8Ha7SzI/AdiVuAzukRIFVil/mncluBt+VxX1U4U+KgwF9RdSrCodLTzKLXffIIxcCSIkbNfuj7u
ZnOO5K2Qj+wY3iYfY0nh48aem/WDYmg3Fw/eVksKes06HtySsVgCMoTJO69D4IYEInTtiLR34bpU
xfNhhq+kmtvhF3owqeUKAQwwa3XF2zpYcYsP5rH/ZLWaOA9t7Qr0S+ljQ5dnYdPtzTfBoF8mGi5N
i/tBqeDxed1uXs0XG5ehGPOv9Uf9mb8dluXinTXClhbj+BYg6P4mOKwuKJzpeurHaKTya0HrdyCs
Rc5CG/Un5XrN+4wuEMmrGaO2l8N05wAdwoY0WkYff21l3DXKzX8ZJVPP6Z7eWDKOTkwqXq3niBIx
h72RbKciRkOdbeX0wk0kBJjyPLeXJQo7lMlgl336mgCArzXbPL9O1gyImaZHrKnjKocXB3HxeTHD
eB4IhlNQ8LH9pF6nJl/fkIeELR5pU1P3Fp/xsCploNQGO9/Sd6DyqAG3lZMBbd+FeOrwrUygOFKs
vm1ts0kLP5b14LUreBG0JgNjHEB7HJsbPRbOSLBTtflUmyuyOyjul1Nai4SGiE7FGy/5Rx8VAtLf
XBsXRva3Q+Dt7bbeFvRYPqnkxj2SlzNAhcs924HSDQs3ddM+LDJcTvHCGZ9WKP9xgLizBJa5b97f
5DX3yLEFMFtjwlQ6gburFcLQS7cElEXE1r6u+yPXsOoNJxIdwUilzZuRCAJVlahJCAzQhlI5ZzNK
ot66lIwHjQUGIZONqNbHWsJNZFOQ6TiLWAAx8U6glHsDTKyDjCjXvHZhsCRqC6bUeDRoznc20pug
1qvyRqOBugKo9hVdZHFTJpd8nCtamMEPZOCueKwvQ4F4teQYxApNiAoWLORM1vqyOHlEb0C4EtZ2
OIVInNE3iVyE99/gswLim2g2rOzXod87v4xuUCN+jIaBGiNHk9AsvLXaWE1qBoUDBvBQ51zSY4Sy
fEfwNwL2LgCeama2ZFZA5LDT9eYPOu+wYQ1exKTMkPOf5oI8KH/28Zc58/9rggFMzwTKQX/FGmDa
DnrA6LekoW1T07AAk4xeDcgqUZEYJhYvLHJvCDgE6gIwpU/5GaRqUO97rswwVQIqDAlRYWGx2iHP
4hJOp+BjdEutpdx6pzEnWO5mnMEbTV9/T2Mq28494KjgtMBOd6weDPTHCV2HudicObtFxOImoh/c
ad0vVQPjYP45wNMUMFGhbMdrWlrAHb3sTSSRHgpD0yJ+d8Q5/np1jf4UJZVK1fZrfDy/NU9OrG4L
fbnNWaHaZIpBpWN+JR85dfg0m9FrImiQYxYlor+oBFaLw4MBM0T8esEpwoNHbVUmvSHqxCLpO33B
HdCInaMQOI0fri2G2es46oqL737aiZWO+9QavahxOjMwZVT/IFRrhCozDvdL9ZOiG2LmQF7DRMDH
exmiLDGMx/aCfO6KQIP/fzrO8r42SmfojaFbJ3mQLgbLeC0nwILk9pnpLAghUmxWQhxOMOtaqZZn
vy8MV9vP35loMfr56RcZZXdPnaPpN3oJ6blIQpxSdzuSvFiEic5LSXQndZYEHgWGAu5vzcVxVecX
XkGhvxJKl6p6To7qmJsZ5IPKyLix9phLVjcVeZ2mXJJEeYqY0zMkmDqVn96g/N+n2Fmysb6XLj/+
JBCet3/OZyAfddUMpEDDfdBwhbWh1j1hsMa0xqwdqzGh4a3rTc03rWDPAG2eZhibxfOH0Q470nPM
WbOgu5Ano2dkpSztNFd3qBKpJI7Hfsw8xBVh5MeU4iN0ggi5dR04ErTMFS+Km9k5M/RdyMzvjmpI
pQMe2hzn4Gg/w0yMrypdh+lUd7theAYSEQNi7LJvbqZfwTdRQiGWs/YS6X7DhYOyLOzvet9z2XCA
U75DkUP+WExa2Gic3PcXPGAYEt17G3D1hDyBQGVHW3qUuz3zyTwSXhi8TGRf1ri5ey3BJqNDODxv
j3Z1HLaNFoMz2zof0udCx3DLMkWVOG6l3YnCSZnOk6dSpFz7WG8wI2s011FpyNbPuF16SXCQo2+0
0q8A44ChZ6jndKVOFTNwJb7d1+uYAkCyfy3iZBz+N0yEBwG5mU7InYHh9YFfcOsSgbyxVkIgeanx
lsdQATjovImos0JAiCNmDbxolnR/4ihS7hhyyACqDF55ZRc9AUTCOGvK+q09SM7TTQo+GItpoi5g
o/GCZeACkGqyV+vzwsDXr1+JtWevhcNPXW9mtMRSNRUbgj3tTSPsajcGaGcLdcn+ttYPE7rr8vTz
mrKYRpjKr9M2wt1DBeDQpeTuS14CFlki+5iv5BuqK5OPeKC2yELSX0LbisVRSYKdxqkXTfEKJclu
rDo3UCzZ9e+9Z+s3mmzzifPXuOlNbvOAaJqaJrQHMiEXT0EdwchKi4ytW5uajn3368xWyaI+xvZ6
lAt/hV/52oz3Uyvr+8KHMWArulYx3C4boE3BWaFRX2BNbsxap9TOCRETMOGALXmbMiKMVqSYdAu9
avEgpapvfKc0aoURW1zrobFdX1eh+ZGGQh0+SNRJIKQ3lQczPOdx39B+4a7aTzwWZuY1sZs4xxiQ
IU88y4XZCK4epRRBOCrHGJdCUE079czePT+w8w484b5LxrREuewtjAHYDVXLLbcfkDozk8cIipck
WXthB8q9uMMTeQ9MnQv/fee95defJt1v8qwyGKKWtRiKXaU/AVAZTNZ6U6iJK4NodMqJ1huJrW8c
iPNyXDzX6+Pr9HN3rZZEmU0tuE8wtdI17INCVwnzkdN53Tybvk4fP1him5qpqNs2chUrcMKBR6Ys
pgkZZo5yZhtEeZM77vmx5Ha3YFeXp0G7lQyDG9bxAxw6tn5Z42oj0e0CEYWlyeIcTu9a5JfYctuJ
Vq+NAUQgv1bLmnSNw+dRfJDa4dmzus8mS2ENP4Cni34oWlrfjY7NlUgK8Yyy//Y16kqPb33xv5Ri
CRlG8XCXujogYkOn7VVhFymNEDrC8dUTocsmGNzJov7v6Jx93qyhTodl+zcth9mxohTf+0dr32e1
hzKW5sV1PyB6cq7p8USuNodEsIjMKcn1rW4vrw4d1JZl8ARzfIrgWLMjMvS6EeVfX2e+/TUxuNpE
Psift2hDhVE9Vkgx98hTIMcx4TjV4/freV0PGs9xgxPDoMrDm2kD8eabK6U5onH9QTYFuYZoeOEW
F69azhDgasUvR9kjc/YGnkjJm6jMShhrijkXKDGunEgebPfzGxQOCZBzVHX5+JpgpFetx/fX0It8
svbhDkF9oMFmPrTbeOlEnxOhY+pQCMPXtRzJldRRZi78NBcDDHySEZXbcoX8iJ/yDiv8+Z1xbQ0H
7vrGAY6ZMb48LZUgwOZDJoCVU1iDRtGgLbLJboHYAOLd2tKlNeB8lbO8C0oQlS2NRLvecEJ+BPji
G50cS2sD1ae31pw44uyWxs1unRHecL30B9oaQQtE/XopRn1uZnLs6Ut9b/eT5NG0bZPm1jPIYnTf
lb+3EzB85qGqwMjxfjy3UusICLX2qSmKsT+hbTqoGrRbFpQM7MT372g2WWb5A4u5+wDzZhdgJXX3
HVNflrl+grPzBuJcBpzcwXh8GBYNwce/8WGRNF+9qrub9cbE5tu0zSdTxQfQX4TBeIcUJpCMpKCD
eVgh0DzVy3eLMlUiCMtb+n4EyMQlb9rMiUoCGZgjpJZbkcfI0fDzqtcDIigkMQbKt3bZVCK7yw5o
jdC6scvS6oNDV3a1sbGf934dW91jhDKbWG6ucXshSwPTBbM/5B5l0IT0Om+EeFc/ygj6GOxDiYU7
7Nfy3ZF3n6CuZhZnwMRq8QNTbGKtxZAb0AMBN726V7lyJTJGLrZ1M3bSwgm6U+xcjjQ8DHChihpH
XXVJmuRnRF90kppBRD3wRQy46ZVo7bikeQgfMDiz7qnzurFzWztd9m7AXKU+yWRqr3p9Fy/X2F3t
SmyO4Kl8ScwkPWF05MbYCQPl9iqpbYfAVTotfI+lHCYl5iIdrzVITygNWX4VAxBLJL/swxZkrb8u
m/b8rS6EhJ14Y1qZj8/g5zf67PRsBbngGQ93PTfn3MYSRAOK8aFZWfTY9DWOpDwy132X7PCDbZgF
Mw/dcZTXoTZEMVqTLYvslkLSD8lk7O21J9hBOLpPY8ZWuix6/zq5kMIBLfjOSJKtGU6WupNg6LUw
LoncSGJPkpUm4iezAZnFdvquf4/X6/lfOXpK7fiL502WS1viCJz4AzrD6iTVnUFfcgEv9AG+ntH8
AD5zrOvT4rWwE+JbxWpY4rw/IIIBTj3Q2Pw5bccRgcJG30uQmx5k09RGM1vdk7HHfNKDvXOvDEps
3XXwe1uyizI7/cwrapY9Q5Dlt1iIAYCvQD/EwNvTU8hphKtPsI3uzHe3eCnCedWTaJdyDoJhOZak
ScTvwVvqbbl2pfj9MMP3hW1z2wiwOE7Vr3RrVgnh4ms0XaJ1tZs+/LXif5IECpt0VesFKw9RWTAQ
k3q5DfkW5uPlpkmTtyV5sjLYzUNb/kI9nJy+v93FoKvIXk/hv5q9sopIcFulTnzBRQvKN15eUSWr
fMY+SXNn7xjh9pL7scOxa3Gafc3weu0+f0clsRPzSRMvDeCgtAp+RsFfEcxbgxCk2CZKTdpNDI9f
nKoL8921dV/s6pzQcqzdD+9QuC5Qc0xSmInqRzqC0X/CGz7tANLZs3PXiEwNoQvlIKZxPMrzZhpk
ustgbfXuK/HGTtyq+zi3OV2XcvbI3LCsQ8n0iVO3i0aU3BnaoXgET7EVoOubYlfuFxT1WuCLUhFc
aTJZKJ40lq1Mr0iFDERKyXygoLPpKxLVIM5mMwLgF5GEcrLcLInVbY520Ox95VVi451IfqQ8yZFv
KtCIzftDTDwAAHyhDedWl+wugU1c6zp603jUZ+iWpwggHwjmjgixK5MXENpv5VNAu0UnonVmwA9j
I5xBk76N1z7h+zGaUB8MwIGw7eKUTScPE12xdlZusxqD2PS5i+QNuTeTTW7B+lQSVr1p/NF7Malc
jnWfaRpRG2iDUyfHRqLrkZTEU3TZgRD8NzG9hHJUpi8M/LcPP3VdzwF5zYtJbKP9BJzMMASoSjOi
dbZRfNpniUUsmKmn8QDHYYPKlwvJyb9zyEHpsrLpObZnQHdnJOWil1gGE8w8hEHBVrFfnkOw/L++
wgWg+GNk/ty1WNILyXnh29H/55jtyJN82ZuRdId+ZeOEtxMm6wIX32g7UpnUhWgnrgEQYbEPnUCT
bOgMRu69iMUnKB7uNIym6leZZ8y/mafqud4+7wZY4q2FQL9FeN0mmHD16nBnR2cpT2+DzlpCIfs7
5Qmbu5x1CuL8GVHx6Sm3T8ifRHUFxXoln3vKdEt3NGXSJeugW/RDPwmJmq1BpWu59EUGmV0TDH15
qyN6J1eVF954SthZQtryRAZehp8Pm5yTFJKVEgan+CSpmM3/teZxd+nve1JgDWZ9NcVgfHtshctP
8+svDizW9txAfe1YH6bjI95JEjyoekyzLW08QpzfaAg8YRAhOtPB6Vtr8jYhPVYj2hxbvA2iTkuO
XOFK/gCTEo+N3HXY5A40XwiPi3dk61ktNdVhXSvyY2wJTqTcEUS60JSZTnTq14lhv5UeCo7zo0b6
5MtxdhnxdFWbH7URca1AvHbvRsRwiisTYBbt6sWYM479JwEnNhfeROvUHbashzju2hrb0WRWMBTp
KBs5iweCvjdKjxaA+qYNAssJGns1ngjwTvnZRDx70D519pALtOoVJ/+UalGHe+Kkf1A7uARbwzcS
c4rufU3dP5f2lemxPLhH/5RV5t08MmoF5anms8fX3YoOZABjq+OZcVGExmC2oemXG7fSkOV/njyC
A82SgR1Dz4jZNerU79J6MgDGA6uPK0ShP/chrfb2aphURjavvCxdAAtAyAh7NbAFxwVAD3t76T7F
+dmBcHzXRfnD84D9zMinZjInMOzC/JnZKJtq/xtIex/LT11+Lf2fGuRQvoUIQuiWLWe4AefzmOZp
DHr8Lnpus+Fc+IMYjDB+rr5ubH71kw+DLZvYWe6AHPRPOe6yLfvsmIHswis9Ndlfpyv8aYVfXls/
XWkEgIwY+TfAeqvL0vET4/iQwroZ0B5IBiSo22rV9CIQqNgSy5IcC78H2St3+3qGvnk4OrN7IpAQ
u3ZrjSadWsW+fjw4qAe+HNlDHzl0z2QFkxCHEyPLQ9vVsTL4BdodftASyB7w3icas06pxct+nTaK
rSvcsPqSI4124kJfb2jHSQ4g5qcax3NXUuzZEDpr5lfAhBo3cvvRSzwiZiNzVwHx5BRPaoC09jFn
NrZLcPNK17vChocasEK9s3vWCOMNSQVncrlQni26G8BOdCoSNcq5zo2Ef8eLuU4oiIJif5/vjULC
ZHRxXg3tTZsz2KyKyNPLWf7TfYdQMz+9yopOPfSczRCn3+CEehUNlZTd0TawtXb5xURUxTDbSAnE
6FHjQYfYhzgPx44jimspaF4SbEPIqkg/932TwXZMD3LRU7vvZauytV7lUNL3Usw1r8GQPEef3q+M
vOPF10jWssQmZZUZf1NmSivKkZzmeJfpFT7Tx2LBi6weYwNkrSVo/CbbgGTIHwytGkyTP8IXgxSc
ib5vyVH6dyoFqIqLjP1DNa6/Rx8tpZcdZgx1QrqunlfEdVU59gsl+4imORmrr9SA9vUhWsf6iwoM
sG8Tq5IZrhUSosKzYsQKeijvqhBeZlUEEAlvpIJJ8vNSUk/69NaI2m0yLfJLNauS+LXYkygCS4+x
T10Ay+Jt4WAaeRYSVGVcDfOB7fJ8+u0AKsz1OdG5fBJem9hh1/l+9HAF4mLEqZ4DXvdVt67bKget
BDC5X2PMHosaW45rKMSzgjfAIBxXGtlyFDGeB4MXsRRCr8cvw3fk4n2VPLv6u2+UNHu1xWXSEd/K
dCp999B7AbxH9+G12n/lk98GwnAo9Qmf90iT0d5VU4m6GP/A2tCjmVuicsAsSVfGYKSqyVFWLNZq
76y9c9WwVIWnePHy9qNCnBo6yZ3fNdSwADBAUEZ0Gv/qyb1KRr08Ir+MmviVg6JD5tkok3vpQ5S1
GcuTm6B3IB+euYC9ToX9dOAbknhBCQPm79F7RV5UiCE+vRZaqiAqoKzmmQMstVamCJ74qoDc/n8e
7FtECnpRPORb87kqSR5RPhlhzxAbxBskKRZLX4yi/99UVRxqyUg/+1mFE1jsQU1fmzmXw+sM45Xe
+fqoWIEk62zVbFzM3Zqe22724jIQjt18IKRm6zIQGYhopeWY42inCBGtO6MsB4BsM7lEx3wGb26v
ykZvDmnfiQAL2CV/kqXljfPq7yuJvGuLopOpLyxgML2nPAQ9vpf4M+z0oH+7M0KEYm5WOrQoTfns
jEBIo5kVMLoI/tIoyTccXhwzOiS0AgtMOhZ/n/q+0Q+17tIdMc6qmTZvs7kxOASWtb3ORrCxml7h
ey6QijqE1fDtZbVD+w3PZ1nB7EHo7q/QtbwYGSVvpZ7tvhrj5O5Q293Kvl15yc7Hdy3GWK8cygN1
IbMF+HmvAdwMRWboXVcHaUkf+q3GJEnCCZdvu7D7flaSqEzGQgtVVVJwvPAgT3K89E1C86D0hmPB
ViWEc2h8qwciZh2lQNiBkRqnu4Z5rTGk6HILc2BPe405guWr8l6mWYlbuFif54Q+orR58qjirqZz
07r4TtcDmUXzZyjdcOYpQFD3p1zZAczVukn86QwSLEAD1VtSUX0aAaHu5snQ2ekOhO1FvYBGzbxG
FPqEJQqxJXNMoZ/alzXGNW+g5tcf9AY3kXQaCHeJx+ekOPQES3gwdIifl+yaD4O5ww0ybWuG65EG
ggt9uhuPk1Ilo7jocASIgwJM8rDdzLqd0y7eq3oNGAzWb88fxnwc/P7AgOJEIZ1iMQqXkrVir/HL
VfMAMRKoEKjhiNMhKcElEx9AUCora+tEYNdMQwAQchom6kD+32+975ICueyj1GEaEHqm77C5KQh9
DMljD6a9rQWnsQINvwp8kOI0a+qeAzp8CULYXg6+ddsypHQZbNupkBmuJsXs+El1NpRikrAV+wL1
V/d9XtbeunsaVAjSEyOONcg4dgrGzIFBxXiO7HGUsctjklDSuwm5szho9D0Jjr251R8/LyOUbEEr
3tPjDXFFZ6ES/KvDCudkhlsmUwL9RvTpLL7YlWO23nTFHT3WM3vyuQMCa4+dVAzbMRe1EnxLggQ7
iNieMIK9Ws2dC3oxA9CCR1XNRFRFs1mio6lEB4U3xNfC2XlY1QSe8RvZle4CxJp7OJbRKLQ+eu+1
d69HCsXA0PyEnezwCfXOvapsISsUX/8Qru98RAE7NqYQAQV0yFxbnQiE6IGNaDQoU0lwNWosijUa
8mGY5jscFSpYqXnh9c0gItyxsiDXanzBhnIbve3mkKbCb+Chb2XXu8/W69B144HGQFjnxbU/QKU1
0Hvg+lzwycHOYnnek9dVHnXIaiLNTqhHCtekGuBnkl1iohFjkW/sivmbUzbfJuHvCx6gKxwxfrBp
G6TvePfTsLpq4fxQzeUyYraHrclM/Kfh36AS0X+WGT3A+dpblXx9BCR6u8BxW6DK8ZC8q6ClpMNm
CaO9dMIeLpAiwTGIsbAhhewzEHWa+hR7fuqoFcBEITFjKjoYgcxa2w1sIplILpVgBzXfUN+E/Tas
SzbUm4h1Gn9oT8bUCgnTBQs9+3u0Feb3inrZmATcRKxLINJY47Rm6b04GGT2PF/7XmMoGvPKWJNV
31IjnNTReoTaAsTN+WfQzp0q3Adc5og2AoYWXKYdYZlKKuxD1ehvy/d9LXJ5YwdwUTAcA1zyVVog
nVa1rSd4bp8sjAdyVXrzw0YPZwVlQF5cZfd8AQCkkUqXz9Y+Z7QrOjKBu19i+4OSg/71LuXiwWgs
DeJ7x9mf/orPzzTshX6eHXg2VgjeK0BYfXPuwo3QtqYNvCdFSoDUZPdzuPjxvJ1Xt7kMntQ/d+nW
VPftE2ah6cjuCY9d65WwzPeGVtl3Es0GEpNRzwU61/nIabigArAxnblKdrErZzrZj+TDqpVBeEN6
J5oIi/RR0yH8b594GbkP3UT9Dd9rFk102Z+olgGHd5UrXTqvPWXhjwII9wSM18wkGFu064tRA7CH
cplfXtXAyil9kOxxmEYIrWVI5Wf9xFzUvqsNbcYm1Cfd8QpsTXeHgeXf4VrM9st5qlARuWoFZMLv
2puFFgN56ol3PlN3rOImfVlfyn+NKahjFCovwBsUnX4RxT8DOtyb25Cd11PMslMm5iOoppdwRJ6t
KXcYKKYD/Hp3s7oNcfsbe0AoXLx1LpEBgEaJzhjt0ixLpdm5x8wXKyGrdYcsLaXehs/lraPaZVfv
7xQDrg8YfOtvMG84mZcJYAG2cPDAhpkgk/zz4S/bc4xjmAKevBwxgQhMCPaupwRHDcF6B1twhzSE
nWRlmrKJgYxBcY3bxPUt2Bxv3jusggXm56fIJQ3Pj8m1pjRleVT0CTP7Z4x7hU0tJ3Wm9BsHHnfk
QYyHsYiUGtCSoouj0qGMnOLPXZc9q6QHUGaYfMVxuFeWir0+ldYvNqU6bunilH5TfhmimlMbcm5e
EJTJXLmpc562eYPMhAZnDMy4DnHOcmIj12ZNnpe0FowuJep956tq0h9X+zKOebvN9rllIwjRHusY
1UdHn10QT09aWEVRWenX+PCYRzZKMVxwSLngHQuKvn00xUNuaTIChx4B9rOWR1znRONXhNltcK2v
XTeQJpMsQWHkcKsMqhEZXcpIKlH8Mzxxca6aTflvfHNVug7+PDXE2sWPWhJZwVnJerkWHwYKgHYm
hhRWFbEKkwvWUIl1+0Cz9ZAz+cdYWJv5XtcBkCqUBi9C5LeV6HNQ3XrYxxtp9ZepX6Lu3wjUsqL1
RXAyNt+tIAF+NMSoxcB46P6KNRF0uIxsqfRmUTvRm5L4h3Ybu01KIVWIgWbOk/D1mrIuLEPAoACb
welVOWQwoJXcl8/W5r2DggB44+6em5ZIo1C6KrkDDpCT5h1HrQnhjQuCcSZmIXjIG6tGYN7FT9gW
E9nHIcreWKw1/39ANLdtSZ9XSOXUPE+VZqJ91pQME/mQHQ5yKO3hggtvc1jzpRt4YRV1oNTExyyt
G/HkiX/U6GdIST0peqA5ZX+dEgs2ZC6Yph4f68jB02+yajxviBJR0TzTc6xSDFnjj+ZBflRf5FVG
HmqCk4fzLdHhmeaVKCsJgGyHq+vn7qbgB4R5dtmC4BzWwzRvxrbfMK2jGXDHlOOYmt9yu3VN3Bvd
rJ7L1viDWS05lQa+8yptAAxi7ccxzj9LYdpTD/VS/vUmfzWiLtwf0wYX4m3oW3kDlkRSRYENKqwy
ScQpWSOPwSa+nmFJZmQMwFnFf89IZ9kRWIQmKf57gjNZ75H2CFDzNZ1XIM84TP4Kyk/vJ47XM8h7
/zEEDMtTouqxO0un4mM1bXdRdw/VUEHVbtIeUJwEO8MqUhFJtS3Yv7RTAY2HM5tCjm3UVGV8G7RP
CJHjUpZqG3GPOH6fodXOJcn2HmFr/oH2uqxCLqYyekGFPOvG1L1noEwLOW8nIVcYKjQHzuWOvaI8
Nt/4qzG0UYEmz9j8GjYFJajAP2xQy1xQPkr4LGFMowsU6MoM7Pq71avRmqBtUEz65i8rE+nxprTJ
d7QlZ9SwbgfY+gCzMHpLKPf7pQ9l3JRW4sfabnhokVF23EwsA+2dqd9aISH4rpCBWA03lr4jv+Ol
qqkKH5xK4F1e3n36tZ3xwkP/4lDwBpY5ajb7aWA354UTWioq9/U6CYRDac3RtIaxpdgu6WNqNfaU
1l8FUOMYt7oYea4ZY8GCkFu/ivfGzjOsR2GRvrYnTF3Pm7rgeY7zHTm2K4Opnz9JDtAQcLV4vSDp
kBVRAdXvLR767hONvzrXViJ+8psVTq8HkfnAnV+9sEzHOGk/ymBnRSsJCnv9Gvbn6F1zr7ZCn6s+
g3YuWPZSDpAs/+8+uDLFXaL/o+zH5uHi79B4Wze4uPmXCGsxThjDEJVWu1KfKfVu98Sz/DBoNoEM
u1Qu12M2+vy3fyc1wdzTXm8l3vLis1NFsflJfgrpczItBWlss1TGKnvFQRnAlLzc8cai6lRHLRWo
dzXh3abt/Yb7AzcIr/STdc9cr1H0J8HpdSXLQ2kc8PxLJHqtyJbLEESynI46t0dzAAu+NBS6QJn2
h7p2AB/8fhmKgntEtTIoYKyJTGMrxZEvaA/ruR1czeBETgnPlXayRGQ/bJT+IjpT6NgznIR1D7tE
6DfeUJXL4CTzDKuWsGvoKugQKdG33ieDzzN1mH9TJmSkxcPLMqvY7v/+t1UQERRo927X8IvjhXW6
3pK7JAvHHdzj083u7Jfq593yWvNdVilBCrFynb8spctlgnJHqrqRvJDm2sFTC378SCIviLNaXUdw
XvV46plpUgrjZaLbHLeAn4Gp886xMkftz09/i5OGKqSQYzhfR49oByBKibt2CdaBA0+ve9J2imO/
yK5s34P1b8LzChRQExdh3bxmQY2isZ5/ssFOKMbfEhxvIpR+43dqaha4pb3AmL6T01CdMxi55YEX
vPcv8wiiyvz0Vfp8ZlWETN5e8T8ebqA5HnIxNcuxtRbVvPgtvwUTclot3MqU5iXS3Oe/mWDerCzo
tJi0GqaQ2cXbD29ZjXuhW5U2iKI3rv20PsnAWsoXAGJ5Ww0sTR7xxKQoBAg2a8yGmTEOnTCxtfxe
PDEpB7xYoqXm+yAUq8/KF1iEdM9AEZH+7v+iclkdW4z/Tu5+sv57qRvBZfAnxD8s+dijh/s8gIy2
7ZsEh9U6g2MF3+EiiupfsZKuJv/g56OFXssjE9COIdcvsVFnSDDMqyV7/sdIXW2cXwLwJobSWfBR
HtKrUdVVnBx/r6UJc8ytInDLtBeGOg2eCzzpdLAMaKC+ptNZe7QSmmN4oxluohiVuB+M17szkXgE
2ta3gAGs9SujHkXObt9B0xuMn4vhN18oEmtotVPk+M6V5kuR0y6j+a2cH8m21uHSsIcdZE0gk3Uf
DOrDFGMA7b9pHPo2XylVWkiBUXCj5ZtFZl6JYAAxV0r+6O91B+mypVuPcg/+A4O9e9AeHjVzwphm
fv0F32DJYS2vdQcU29IQfNseH2WqKQNpsideUUQczLwHatsy3vlVVasiF/Zbt80sygbdDuJZK9Hd
9D0sgQjL/PA0K7FSP53f5XDeD18BklToDYws7lnWr6hrjNaddzx5oh5Ki/mnbUpfyGxGHv8ZXXZV
N7nSxa7NqOtrxkXDjk11aGyEOounzxjcTNibU70dG8jrjamdzhdoTOUAkBspAEpVuvlkqLlTAl4q
WzzIhmpY+mMv7/ESH6btxaThl8LYsy3sYHIZRAlPgXj3UQkc/dUSMEeAgxpEdmqAlEPKerWn0kgf
Cv3MRKM88dWkLxXybA3TtBeC/c21j5xMPnQkSt4GKWGmheR7fZDK2qpNA4D4Ew7RxE9xDhYMhe2V
c3/nhmCzeJ5sMCi4SX4rZMVVaJ8SGZkcjFWbveOfFmAV3ygXLV4U87ye/Q95Wk1I7GDvKliiOBtd
WPh1OtHcJrSwDypD3qa/8nS8fhlK7kvRjf5mb/QKX6D1QS7mdkwsmzGEuVxbFPQ6/66+tJLsumsx
pTYaJFZ0yB+1dIT7GjWmvtondtd8zC/UyaHcdf4UqWmVSNn+QICsLV5h9WaODFfKg5kQzDJP24S0
MmkspA90F1CPEcO9VGiIWnG+ImjIp3rhScGkc0eYUyBNH8mgpgHLWv9X67hFLRgfVKLIkyF3oxxo
S/Ey4Inm3Grf8kF/jdNwIKBxQf6ZdYDwXA+7TPuFM4SpNU5l2SlhLFD1snVZ+DqsNMtpUkRbfyGA
rjezhOCRMzdM78zEiHlRkXkaigtNCjV7EVvUBWVFaK0faqKJqKYN6sLVzFSHvmgKgKYE3fB3sx45
Z3Z2s9VvY5lkkEMm5Orj9WfajuFnygBjhL2iFGRfxXBpzbWMSFN7Q5Mx16U961Q3GQOUyI7gzfJ9
7O5CqdF+CMwKISqMKXNqQoTrb2e9zqqMc6DSddftsCxAxC8/JtZYUISlQTWmETcPdM8tdzD00KAj
WSTOA8kyeAhHMVSMVx1qg7XRfjVF53Fn6J9azfKguWrZG8HlfxN/RARf/NevEQMg2YCLdN3bIrvx
G9olxMg7JhhNu2QRl7EUE/U3jcNfCMY5C0heP4MaFuJlgJ5d9sttLHPxBMpNO2Pj5DNITshkuOoz
Y6JFIAx/Lga1V9lxc6YP3sH5IyzrprBHbY6Q9f8/druVg0RQFumzfoBhFpNnzz7rt1vbwf1u9tKL
7DC1kWe3JPOZGy7kUg1S1AzgrjP4C2ZpM0MfejpZq1X8sVMWVY2v7OnZw7r1fwOYTXS1ZHUW91+V
jTNwiPyPiL/EW5nFmNhYPONS/4fRzNDZjfmI06v1GGhdLkP7kCxlwTOwLt6c7rCmhLxGw6mCPrVZ
HjBKXCn2xbN/20ZpktbQd+k+kbCUKDjEB12cjb+oxssL8GRt+jI3hCUKN5GBBpBYFy/6e/GFHFq6
wqXopdSd1Z59Llix4UmVv4nNvfndpzFcvPIenN8RY3LPbDtJchLh5gGY2GFoN2z0h5Sez1QAnFXm
Hx8IIPiOxB2DpAtuvgtxCy1u72zWM2gPLul19eOoxZcRfXK0BTQkfPW6yRo+ocy6tL+w3gA7I+8T
7r4amEjN90wBkGbsb5pGK5wOrseZeK2aim3cps3KFOOX/030LrLdGgGRlGRhcB9+OO++Tu0c3F6j
GzO+99KLyfw0/IZAk9LczWdh3v7DNbX22+YxPrulFYT2cctFwbvSqiSS+T/D6D+Cf63ChbJhfzv1
1ePbyvnDc8GUkBLFgs4IIfPoCbVqwC+qpC8/7kA+PQLa1jA6ALX1NvLvqT+mJmxvoVJDgY0ijhLj
FKtPDBGyJc6ZBfdwhOtaueJcxDxMzSolACvoU1l3FC6GTxhao4spOFBhTOGpOBICO8yalheb1E2z
jhWcV8163IuMFIE0knsGV6h5A+CsMpx2z2h5wXOCjP8ZWLJM2sSExRY42I5R38bqTIIUqX9BHj4M
L4E0aX5HT6eG6Ob+V9XNzvBBpDl1oI3ic4s4vRcm0hTKI8gowfC3yxd+JtmsxDFd4s8MgTCrrvMn
kNxOzGXOT6io2VLJ8BSFUOqvolhJpaW5C1XxUx3rDr1Mx/w2OKvS+NKipVBnpWxsoAr6RhiQ9rD1
3o5Sb6+JH9XSAMXFacyk/mh/4WMVV2P16qs6EK46JP/qOP91BPfPOZCrodrGz4mXH6hVuEGILAPv
n/2PDgJM67kc13Kf3ZkXWYu6Fwe82FQmHT4nWFIB2We0XIMoU1eG31nBTj2M3nfTgXTAgtpUDB+J
5awG1Q0iB4128RrRmWPTsQoHoHfa6/pEJw1r2jgaRUzVskT8obUc3ED0QS1/cESwdv+w+6F+nGbz
IDY1q5unGg5tco3+Lr2cS+CqdQ1g0zEhjRrgpNL1blllLTVxrkxPK2+u0TXuSDXDtIwqERaAZHnB
5CCG/N8LfxXPL5mSCWty2DTMwHxcormdwo4mzHUhx6zr1g9hvxJirKLurrhR/2esYUxZUxcaSib7
cR5X89VWSvtSsZfiT8Dvj6MHqBu2g3kuu4omMMLxTD9tffL11zcrnF/00gkk8Iz5JGBFmK6hF14g
uX6QKvLn3gXnw9lHHdYDuAIhi5lX52a20r2Q0KI2DkxTuxQM/1cN/tbc6nhLVPV2hIzD8VRXTis9
dgPUI1s9g2qiTvSS7o91eKQM6r+D4MS/jRyZX4htvcPb/Nmd2GtKR906MDgQVE1DX2vtyaD5WyGU
uIpFPoWK7EcQtV1WW3UdSnushU9yVn/QnLfP6GTU9H2yT2Joqksw5jBBcPWWadtS0gofnBkiYe83
2MAn1du/XSu54IxRUbh5oXqhgCohh28I4w9UqyoAnLT7Mal/VaLQNVMVLbRSFiNUKQ19n8kD5SKr
NaO8qmWS2xlLwamwS7go021nriJ4k29nua+nNRRwjYxLe0ylIlA/EAS6ohg5lhVX4Z4wGww8kyBI
9b7SU2btNlogGDt9koHXzs2SFTcDv4a/d61lbCyItv93DFFKg8vWd0GWrTVkIASFO9f1zi0cdx5V
hsr8RhUeVbda3X4Md3WdncY3z3tDCRVN5zjnyrw/4XdpQKE6GAPNSNCoea2ItWxVxJwSyaLomVn1
lY7cvWVHKedYL4m7fpBZ+mgyrVbrcJVb0JRkSKTDmL62WKTPvIZtGqqC/t3yVI/sXmxAWvhmIHZZ
SFm8TiOG9jSOHSYGjiQ78mmodoGfoz0Ksxj38nuQAYN+0nAWer/VohJxQUGNBpgnsrmKbpg2aq1K
nHashnHi1msWwctsWixPr8UuNufgqS84LDsztWzX5ruiN7NYqA9M9EDi9+aHQyj1CGVFMUN3uedG
2xw1Ru87yB6CSrj0zhvZlq9MY+Dr10zrc4/8jYaiJjkNQxjE51RvA04QXlDIESOrgF8Bp6bmnquV
o/Ht9B0aa5hjBTg+08xISyYGMg1h2VT9qhFU1e4RtxdHf0yKIrT4lfkysnUHX6IfYlGWMrJmL6eH
oxlBeloskVhhz+//YZLZgP5xak7jXik1nkTkCK7j5Nyiyjc7nb3j2KnRj1j6xH8rwcFKbncr8K3X
6nH3rrYdFD/7ls7CISPdF8zgU9qFsH+DYO3SELVlsBbb2KgKqP2tvaP48iuqJ44CHCV58hze5RNW
XQX3/lr9wLSmqYHWP+CG7MFSGCPz9U7wBLWawo78xQJ3AaZMLGif/767ha/qZT+bsP/+UAn5dtQ1
lNc21r3Jwu6jXSPApq0DgcTgItiSghXRFMwXU4md85+OhpsH3kBpVfgpw9Y+foEBa/wjjt8W3O98
2wNOWdq4iTfO5BIbAe/AEJWlQXdXWqwnGhjS9fBgVPi08lZjHqdlxyoQ1fGtNFv8neydCeXjQYtr
a9ywyC51Ou8Q4jXBlSFO3gQ1OGdkPv3p8KJXEAjymEyLTy8ekcbWEaeGRQ6x2sFF3fmYFEKvWP0M
tg7Aq7UlNaYfE2EZPiFaPjer2VKYqX378j0mik7RfNIBo+dYzcy/PUq5ybB2q0vPYzKW8Kas1YOA
Z2iLNlrU7zcAxw3yTtQMrP0tSJr6mkw3tBSWZ9bArzwAaSrKrdF1fKjnIwFtdjcc3Khf+/9KxOWe
3F1W1pltDkKfcuWR+2APL1H6ql4YWM/HwtDPi61vDi9l1JD7bQglyU6Xp2hs4avjYRskfbkBRIp2
jvlv5M0MEgnAhuxvlfzbERz/lefdcJOamoRXgezMiKUh+FIF+Pyo7/0QlD+t1oOXoifDh3jEfytH
28Yv54MECVPQF8VGPs0OxnKwfuzTm+6ylLRIxV0QaSjPJkQdf153dr/s8XyRgXxA0E9AX0Il9kW3
iOdBFbe2/fpekYkRkNLN8ZL5NCJzja88DpYMDRs2u2QNexDsjPpoItbSJsdX0kkIz89W13JCtJt4
VZDGxMGROaBKeD5JIFdBmcfCA+1oYVtiwoCh7u+FgKlMHvwr1rV2U/BDuLgbMbmxQ2kO+KNrZJVC
a1M4URObDgAPZrraYCBaOxiv1VOUz5thfEs/XD+rmMURnhSv7NL8I5YT0WdqF7WS51ui21blAUY+
4qLbdr+KANk9EV6O1akxbBDQ78lYtM1Pg5gTFLCsbVvMkjBT127PJ0F7y2KPpdOoOQq4cOHIZmeV
mR2TmLpOBbfYmLgkJ8yeTMtAbDxpPB31j5lmVSlvO9jEBfI04YenrUJx8ZcDbqFXHUjusCbjbpyw
VMKZEb/tSd8f6tcWDqBJkOxWc49FQkCcdpbUeNGT49X2IVUxWwH+6xCMNXYQu7oaf1rdES8ECTpM
d6vq84R0z9OGHmuGBoavk2ogA7PZzkF5rIKh3eL48l4DtSMCxYch04FTpkz+jHN3YMOKMi7Js4+L
9hDR9CL2OUdD0QaCoyuJpsYxYfYIi3ld7gsT1qoiONGrXfM/cxf1ZMcAtT/RqmBVCnK5JOnXbKlW
mmqWpXnxUZSwFWbjILOIcJ0xCGh7hBjn5lPJ8MMgLQeT1ida00fGzG/Fo0VGxycBn9YW8ozmjmFc
b7ex/W3bI3VMar1S+54Wb6agVNABBxjeKamjxZ8eWxTIKOn0Pz/V5j8BQnycFKKBiGjJO0M7qriH
dq7pUwStQ2psp/fG2VV6XrI294zTMEJAHi+HBUFMBj35+/4LX3UJOFGVL2XdUG+VjEa6WJIZYJYh
p/5Y9qqzWw1D70T9dLUhAMviyosKo+v4rlDJbY4OJmkFzmtV8Ve2xq7gA0E5lAscfC6y6acf1Zue
oTBuDQqGyddln4DcfTDcfWyB2JLnmiGVM+ZT/5AquVej6dW1/xCE/oQI2ODQTO//YvsXIYdPTooM
c10KTZvcEU0BMc3Q/vvIvXWddW5JYRgpHKlIoS0ZsVvtW+KAjo2lz/vbl01mUjjW6cY6Ye6t20EQ
k2tOwEtIJNaRduzFrGr9L1GLExs3uwmF3KOjPXLVxc5MmkfJ7A2SaZN1Uz2psrHOQGUzkyMzs7uE
zm3Zjh4UOVIwFTaTf0ITa5lJYNk/zPZQBQjuSJQxJEs6UO600UGXDTNAz3wGciJc0afpA1wM2Vfb
x5zfJNoyxXJ18BeuxQK5lICd5nXS+vI9stHaN23lLJTn7TzA0GS+YbpPBZ1ggWdzRcdydOrpxK1P
AhV3ViwWt9ngqXITG32ex69h/IwH5K0GLMSMVY400S7cSaSL6J9byfGmEbY9nGzIMvkp36ecyRa1
HCmpG+NemD2llYCFo4yW6ouvE9nG4OyLcZ9caWKhQFBPGUMCEERIajOKz35z20FeAsw746ZvpeY6
misFCnXSHYSWf1/NTY8nwGssSqZCnYVKvykVTNEO1V29VZzeLdhGJhrt+FwrqKundniA7OVXmPov
VU7kpbwGzjOYjhMvp5zjWXZB2NhlQV4GrjlI7fOj3Y0vuVGlS5M+/e5ZfW298CDpegJY/xZG4F5W
+js+YdVi3YyeUWhzIb9vv8XZvvUT1MSodh7xDm61AGcWstMcY1urRsGBEWR+/2fkaAL4L2rvKE6K
kTglHGHGY8AivzqPywdj7DfOTqxL704pPsNC2n1kU5CxbdiGxuwTSNIdqAKlklFxfhUfnlZHUWYV
Z7mdKBLvEyHyZf0c/jlV0U5I9wvvgwkhdc13LcJaJMRnYy/6fmfpaLQW3LSZDC1PlO9aiu1+svOr
E0F5N5kGhE3Qm0cHOxT6wjIFAPVcKCGtroLq0tOzey4nYEpPhQQWyrYlQcc6v7vYhWJPbW04Kqg3
OzUxX9638kDXJrvMdy5Oja12S+dLm1kV1O7dYhaVfWvlXx12zCEW6r5L8m8QNyvRoSipXRxZqcvn
M3KsMPhD4rrxDgoyesDL6KFArA4rqt60hWpHwTQiKhn1wpEAHRxaTDJJkWukBCXqIyGCY35VfSq1
1S4KyCY+/5FeUTBu9qhYLfRV9yIYhmrk/UuugPS3aLaljSXw1uCLMvpT/0LQOWguOK84kbQrduMq
v83HAAFiIyDNQeZRI6IsnVD0iXOHzKww02+ktTUzSN6WvOMjAnyVPYwO3We7gzwJ67xcFv19d/Z8
jOGvK+nqyuWISN79lDSMO/Jq1nzf68O3lryJipMQmoj3kA40gvhWaexudruElFyj9SpGW3rSDmJc
eQiG82IOg51rIKce2izL8vrTz/ttiCvVBaeNnoZB8k6LSdzENUZNXqK5UWuCUOfnjOkriz9hPklN
pAkEyX7V4cFHjg/SP3w6p8P2pafY8sYU0JGAIpT1ahDVnrEO5eMK9XHiLV+nuuBVVdywX6j0ZkCs
Zu3NQhi1k3JbniVuUbCV7Oyt9Vq2Nk6qt+t0bfUmLvSmXRY8wteqXHTsn19JP7Akv070gi+FqGC3
jcrX0XIYc6DT+P8y/sASOcIUabbPBNwVxPGIIcUtBITySgRuw0L1g6l314LyrVnKSWXK9i4XlWAu
h1G/1/cfD0tIPWxzeLQTf35NxyzGI38GLlvtWp3FLGb6Cy3T7AgOA4Dj8wzYPpgOsggfS9pzDX7D
tLP6VpXD4kipNLO8A6dbQCRB7YOA8WQ0Zbb+P36CRMS8b4x8kxv9bBLDyU7uy4f5U7NI/a/sO4sI
0mjyhy9SEuLjvK6nOdbG5R0cab+3v7puEExYuCEgrHdQwVhTgIog/UYmXqwo2oNVGLI+dvNBRztX
ZGoqc/2dtcd6gpdBpXpZMPUy0lu8jdL/BI1oaodRmIQMfqjiqVGD71FYhiSkYxmrB1ntyIfroAsV
VaZ+QjqWgQHgvmxlgwjBDsNtYJC9Ogru1k3LeGhMkcAKeoPNiumJ48sHcKc4L3sUv7OLgnjGxbxr
AoBa6LUHr+twaJsk/cqHDaxwaiIn6e8kFcWekqAWVQqJjxMJrJxk6Qb8TthHeOYJV8zTmUeir3aD
jb2DnOw8TKtC5pM7jc3/dflmSn8U3Mr9vJ0/gj2iWrr/2W67XurM5+l2u1KxWiuqFsflwEKtRRm3
kVS75G7b3A9brfFsYw4LRlZWKuorR5Vr3w4GGRaI6zDWlAdPSu7xsdN6FatgY9LQvtCjuj9cxvpd
nNh/ShF1GPo6asgXu4yDGU2wrczU0zbSs+sDpNel3cxyfcChTu0ifQzu5sm9/i+8G+xb2H3jrR+c
VjcMIT1Orle9TOKgsp43RRBssAPGfKAD4eGJrmrEiP1Ws51imLn/UEDjidiC7EwqsHULEPF4WDGs
vrBBp1ew13D6MyBsAiE6YcqssO8hWgiXkq6zaN11v9mL7lOSgSPhyGEhrdOMfs/fq25AQ9H0u7Xq
JEQ4S5tdWhuz3bGD6ncawzacV/YVpde3MQVdGYjuVNvTUWzOop+SBZIhOUSwpVe06jiapwD7N+if
YvCkw9KqLEp58h5wupamNeqg+TskjsfRYkgcqfN3VDMg9s2Njelody+Ht+Tv0kjWmtlYswF1QVKE
CyDyXqlMstamh1WR4AEhL89FdKnRlCOyuYdyMcEvifLrYepaa8dscyrEhmyf69ttxniDxiHspE6d
6/SfyBpen6xssADvTZoXdZ+jKaQa2Q+066DtmSrayjJoYMmZImOI73KkEeO7HPWfIH+H7SlbS1mL
O5yB59oTbFx/cA0M4KWxk/y0bkZmx6Oaiy2qOi0xtFgsx9MbkJQUUUGwhcBjhaUs7Zws8MRMDvJf
CVo1FxyjHkNcoa+2Kc2h3eu9YJuHK9kvF3vx89/hqbGdMhBJSbQQmFcEoRQL9QxonHeTFcc8FC2w
PN3yPrUUcS/mzAU8nr/pWy6Mdm1cVNoxoklYruasE2liRh4bAgGHP8TL0cFdHsGU33EGkGp8tR0m
HSzmQBz3rb8DyViurENGY4HsKrUxqADvBa54JHmdnodL6hIFFP3ZnnLCph5FDsjC7eQw6dsyTYfj
PZdsc/tJv11oYpUvjF4VUs3jZqPEuCq6pJN9zKG1peAMsEEdQ8cr+wAFW5bP0QwQxUPUAVpM0iND
+RyMTmeKiMfa9wvoLpB2XbnPqsPdVi2VnkN8g/ifVATB7T7u5Q2cszCnFc4b82R+RgFwV++1NVYf
Dr85BJe0Xc0wQMkTVxmu1p9PA6ycVLCpcWY0/VUfqSyUw126gHW1uZQnDx8f3iIDsZZ+cw1KLeYe
jVETrxZ5v5wDMM1iFTJ+y0tRadTohV8l1qng5SB5J/jISSrdXB3VrBuapx+Z+x/l89SjrYifgO7C
ehgteRcF6HonzcDfb1GRoFrIGeYBBWuiysQiQw05qsWeqg4WbG/YOmwdsiVeCUflQX7tCg1NagEd
UCeH+UJdCcaxePC7w5JJ08+T5R58mEFtqte6JIIHJM+VKHIg0PDOB2Q0UrRf4SY5cVLBG84A3skG
KVNZtqjFxgEifhXfZO9W6UFIG4VEIcVvYl0Jhfktb6xiUgtvbzki1fiyLars9bFMaFLGCMY9V140
2XyBN/+XcRgsspfMrkn3SENZh1kflVh5ttG6x9s6UXxtqG79WqzLEAE4MNBb8hii99sR9a4RlCR7
YbuvjAprBfomHn2GwAVQh1aQG2xzumkGMXAcI9rEWCBvaiKPnt8YtFmQpBo0crp11hrxb40ww/Rv
XqfKC0aVGAO0mEJB+IpP9uz+RYa0VLKSEB+vqXWbxzYingQwIKyFsovBhsRZBvzVyyAb7aWyHhIT
f3MtDK9Ygx14d3lJB5o7EptxYG4TaVt41ICoFUXAaK58KDiV/UL/AXb6OlbxIzznzxEJs2nGkFn2
obwQHYYfbYADawJwD5k2umCBSSkeFWCuJfGhXixPx89EftvCnBufJ43Oigi09ntDQldm+dASz/Fj
efubGz/kHdLjLZWD5PAxWVyfxPQLq7AAa4jLeG9kP6uomfo51g9vJYDREfFJdTQ6mpiuB+B+bllV
hINOg4smigzlOGMhsKcI0epTNyi8WlVODq8/JKKtJldrr3g/BChx+l6gQVOb4z2c/DCpzaueJ975
3juw6/Ric5HpQlOgqzDBfRJdM2EeX/lvHyo7fDtHE0pWK3S5IXDaSbEWlhiJtFDQKn72HlDXIlwd
WwBoYTObBeL6AhRuOQtPmibNZvUIIFQhKtrpx9v3qs43CHAXr5ILgY2w9fKncTVNQ5px/rtQFHBf
2w4SybKAcMEp6vibXUvPvMZ7Ubzj6MchsmZamaFQdLm3LNsGw4izM9TosTsZ3i3rIs1F9vBY2b7I
Vz2K7JvIP14dDqYqEvExlSb7cd8PB6xQzs0oFkFcZZhPN4Fnf/TwoiqxG423WCZT8FbtJDfYYk25
PRDaaZaTmPl0aNeWCgXrkoYMqSamlbE5v1VrpK9VMGgkAK8uqwjHfJOcgAqcOET5aTis+SZo3535
cGrrBtwLZwa9eWnovnjQG5jADBGRqOI57al4gk2tHw0NamUzUGkNgOt9lvrqJ4jdcbTPLBAzFDbn
oA6HWNDnDK5VEfhusjypjLE5Yx1wRIVdMCpxwIEPqNhq/1Rds5gQqKhujOP46NVJP02PTpQT1LGJ
8d1e5ukbwEEPr1Xyo1oe0a9zUimikcZX6Km5BGM0rEU/sApNU03s+cQc6dumUUMpRfwatc7t6Ifs
Qkc2YwyXofb4QAXw2JfjPdb3WPjE1g9x6tpASyhTPvV8spKMI68y8HPay//4OLZx3txwrJe9bABG
b2myGClJrw2KKMAm7VS1nCBeCZYVktnEJVnByYyvVok+/TFqhb2famjihRG5sb9PLB3M66T1b10o
R5bKVYjUfS//KBgvp+ZX7WpbBThtOuDHEazkj7LEjsrAj50a7XNFzAUjIfg+vI/HCyfi5s3QdQZ+
A6dcVV2GZpza0xtIBx3JQnwQkUqBkaD/SNwzrdMds2z4b2+lZqfjbEta2yPQjIy8WpXGjDPpYzlA
BeZ6emntSPU0ZbLRYE31B4lzkqDjHwUtLX2AQB0zGVTQyfVGAKnZAt0rUoX4pCzk+WK2CEf/z7qz
fmlIqhBHfbUTenjodOopFw8IxO684CqZeNpoZ/CJgXS68twcwMv6tO6O6CirZHqQd82fAdbZdjfL
/sufeJbH4KRs0B+T5dWskxRQ3bywRRPNhpTj4deOIlW+dNTezxbG5m+L8a8iT1eUqwo42MTl7ged
mcwmexzBbEI6sfM2zxSH/jnaG7VSNZKFSYvj1J5R1phO7kGuawf7ze3J8Qp9L1FOKx32x21raK2G
7SFzAr837gHgLvvQLLDqjeU+BQq+l4rjulO5R64DG0Q7RkQwbbUE5wVwaNz5LuMoUMxeC5RKf5Aa
XbAdZwe4yQSmgIR346ehGktZwwASsfzk4JIincBkOR/xHnd2nQi0kKsZqzCFotTINKLH/LiwTG3X
IK+UME0WjZP07E6ubkv4mkDGn9QwtoOVAsxmlV1+oka3k4bz1Xhdi/QE3u0J9wGnBj0wpdRLIn96
rVtJrntpgYWg48gyQEt0tpHrqTJS5Yf8R0SCooHmbC9+MBPpLbCzctruI4o+N350w22SWZLO0M3H
HU5SDj7FdIr9IyotY4vhl5O5n0zBoZNNEUC3RgD+bm1O/eZr78Cs9JwrV5MJ8OPzRT3ToHO6b2Z4
n1H7mKKsIqcsqwH4NzRKv1LmiTRaxmknqEEA5cPDMNvUx2sKtUJ6aRbgW9AAG7G39AWwMyBsZtRd
WMf+iCGrQAC3T6suJPkV/V3nfuWqoV/krcZdDgrT9FtON6h6sU2F+OF8bTxZcEAdFxx6ZrOLx0JV
mM3VxW8QEe4VkB0GIurBfVrrHYUgRExGgDQmEg7rXFOuTydOkp4Ff2VeJTUQxc7lUF1rEKJw2w/6
NUVipUm/t9WZoXvkmeF2uE/cN0wWDm5ZWPU4AY1DFsaEtXtcxdZ+Vp4ERM2WzCGUEtB0qEiwGgf+
1RQBqw9hl4rm8aBwFYq7IQK78x6UgJ5N+fN80bizulKAWGIBKrCHbqNGAN5RYrqRD97sarJokKo1
Ekr5VZYOnI8W2cw7xg5z+oPDtm+ukR3PKEklSgmKPrK79sbr0EIgXwFSDp8frRiaQYz0obiVVT+2
p1Gx/hgzKQF2a6z/7EmLrFU8Fcnr8/epRp64sYl343AlR0sLUGgbBs5IOiJipQd03RJfPt7+vzXG
V/g0A85Ik6wDeGs95j+eisvrvFLPTRBw49gkzQBBuuuWnGbPRdMzKE7y6Q4qJ1o5ZCf6auv6eCe0
5CFJngOGhCb6CnznYlhqA56lh1bHFxWz0Xi6Ixi4zEBqjOKMnmco/G8mql2TnyJ3bR2F9afp9II/
Ql2qLFJ1ezRNag19ilS+KdiGuFKNJZr0hfzpNG6ZfXK/ITfiO7OECL8ZiWU7A0pZq+Wvakkkie/+
z1V+eCNwgVkHdLkOTCoR0HsgVfMlpU8z+wJXSjW8iyzmPTqwtgKd/fELCv0bJ5ylz0dVaifT71qU
ahqt6bZ0UEj/YWKQUeexS6/FAkg7Z0lkbuqK+Ent2KbhH0fF+GKuYH7rei7PU23yo97qasLG9LfT
6HHDuBoOHuhnoXxS40o48QcAVQJFLeG8DSJZr4c8+YrEjUBbr8t/j572QtCyS6d7CQ/iAZ2IjQl/
SmdELN2dOGS/dilSMxPkoMs8U1oioFusZ3KSqh5hvIlc62bSMwYR7DFiGaJE6CPrbZV25xvPgMM4
jA7jDCOCCjr37mw6EDsvZ4eob0E4wK6bMtChNeFA6gTRubR7sBLZbbkvj6i8uzMfxvKilWpTVm1U
PhIF897CQjOm1UY7R0ijjI+3Qwt0z5e4deos6FFwE3L+/EebD3uuxrj2QTEW1uPti5g7OgerpbUg
/r+Hzow2JcQ24Y3QK90YpKW6UTsjQ4ZYmm2/yk4h0lIDLKQnne3AQsOV8BtAYBI7avz66USF8nN3
fGMsukDt/wXt3xxIoeVkAPvxPBD2ENfHB0VLT8uzCqQV6YRvH0w8w3fOInDQoFqDaZGSCNabaiva
0LU2dmpMTZ5Rey7nfasMHFQMmidjDsRvtDzcAqs7TbqJKJP1bfQsMUVUGiC0esxP90sutRrKBxgH
KewZNcwaEZF0Bqu1jW0rXxm1Vhy1sAnXLpvetuqNi7QOU2lyl8gY+LnT0/jrGkgxyjVr2eF1cxuH
IvVXmqAzDghgVBwaHrMxM9/Hnm2iBUSAnJa6BtIiYWyQtgh+iAVm3tMRahBxV2k/VMRRT8MDLiny
JsT+QmjD0DXIbgXBDs5CcmqwNhNTIpLuN0cRflNd5KNc4q25NpgbYrXlkC3WjC08J047EsIhSobu
bBxrCVzNcYWsrZKaV8AqjB17Go73KC9gWvfDpScODrfrr467Or1JN37xM8am0IPrJGCKBRH1GSjQ
+RDa2PN+xOUmbklCfiyhhZKuggca0FR5XM1Fau+jNSf2f9VXunwN7QymV0V4WY7zzvmx2CWU1Q5c
10uVNlR//3URVJbypQawokUrNYROX00ImjZy4hrr45jw19fG/bHwOjXX1JLNFjOfQPyZ3KgZppIK
ZbPPjzA4MO/UbttELpAJ1AqBGSVjwRiUHwMKuL5H3zRAySImtgi6FZLeffqAMoaot8MFdYw6Xjsg
eLflgCpY7ECxWTrYjbA/UlyiYUn0/fIQSoBBBJUYh1cSy/RIxHp8JbpEFqpB4hSHDpcuPqbG44xJ
gM7phtg/gvrdFMlko8CtclhjjFxnRwV7u9oMcLns7apsjnl8Qkvus8puet6h3hUNI7+pztUKhuMj
eOEeqjuGGTOzbIFWWff6FXOldOuKHAPiCec4qjjYU1YSQUH/y0GDbTlffIa0tJ5GwpZ1fE8Hpl02
6kiExLQKOLcdMV02zSB+RO5vdZsf9a1Ls0rri1oVarKu7i+BDE+zfqs2VRdh2euXHTSO8L3JTqBb
ZBuKALZs5Oq8sbYImXmMSIghhU6tkLTxRO0H8GRkj8EtoRW4ZS2kCx4oEvJZx+B+SbHbMib6JGBM
43OzlChXSOo05JIa+5zMlJWa+jWzxSggNveW1/33rqlB1bDQpGMKKjO496dcbMG4RqUqheT4iehg
3ofhtUiYuiZGI9eNrxlVUKF50sYzhEBCMNdqumtOrdHgXf5d/PdF1co5fEFHLZADl+nADRaN3BqS
f8sbB2K4B8/IGWYUNQ3EmYuBzbB+7ltvr/pjV6qCocy7zoa9/ZS+eyRI8VyM3hnx1AVK+25remoX
18GL6Nq9DJnsijoOsJB+SYIOegh+9Ar0+BZyX+Mif31v5OJ4r2FpNqaZLQaZIYMsl4XFDTj/4tsz
wjCbujsrq9t26YFyAQKbSramZRIGngHUyHQRcjyWWhNtxyEn5NsojRGMEBfXIEHnWPV2sMsC1InY
JZqNkHDlwuOKH8Apg9HxymjeHOCwTI4+SJw/b3ens4j2hV7A6z2zJsgKxRDYsB3RHDelI+qJ3hGO
JxhDQ66vhUVaLae6DRUD3wtR/Fm6v/q4q1WdZyOJsAer3c7sB2GhMJaqZrbKxHhkDlHuYEmpUKFY
wqaqWRD08wWjZRo3+ZUX1fCcIcD+SE3IEUaJfBmPCq/6jKB1jIkEELinK2FQsvpQpyL1uOpaMvJI
ITBXLPskI/B6nSRB9UcmCzzjFYI+qTCZmbjL+7vmkm+drDFhP+MxoQQSH6azjC5qXEd2otcmkbcD
LeOlz+806NQfzpJug1II6ffQ8K+jpKIYcAqzbw6zLq91qzsNTiKgdWAHlIc9vr3pJgbCFvIKMBKc
Z1/12ZQ3DX+cpqpnAOh0TwIz3VuRA8JvV68JAoyEXbpNY2n1plLNoLPMlk/PvjKv5+noGB15/YIs
QLV+lLV85IAZsHO5St3px8UljftxMTbr+PhP0AYpueOzJHSvX4ZGlqhUAEctM3aO9xD0W/YIoKn3
Juhs+NBa+2jKZg5QHgT/VAXX4s1qj0GxuvEKmv5OJiOkb5WaBIBru1Y+xL5tYGHyu/nfC0T7oruD
gK/I2tvcgwfKTVfXJ6/0mU9CogC+FJsc1WZfLVP3HNcM55jg3V0Ye9Oh1Z2ivhJ5s/URFkg5lZ05
4D9+RTNOZaCPwWiARw2ix5UJC2ydnMC9usbqsf/L2PCPLaRO8zAEbOSfLTPcPdkgQUSYf8KT3Gj7
kQoeTdPqU6ch6J6F3xjR/BjCQNmD5fUZ85hFhC8F7nhjXO1C4MVWnLQc88j9kUhY5Xm4RdP+RHqe
Rlb7QmDsvE7izTupxgo3EHBu16HwP2ayEkkRXJHrMPgyIq+gRIjJJVIdxTwvnCVQqgoRt/kWPPV6
8AW14GGbKE3j53P0/TZhQKLr3dFn3z0WP+f47XgeyfO/IBZEQ7WxTLGyLI6+GMGNHgGDk8pCE1Bt
l1opinmY0lZmrBL8l6VifbZHYS1ia6Z6GjIcccvtwDsWu2+lZQbwx9C1BBQU+tO9cbMHuulKGWjw
72CceggWsO7wALOv4Aar46cxERC2H7LPdjfrHf8oIASl77tawbcLbOoCjAZOxkvES1ZXc2bSPeaE
1z/KrALjyDOkGfTSX1IAyiQq+SuzRrb2bdNGAygibJeyemdv23Tf4XOpW7IGmKz/hHIYIMtgSWsS
B65c/AM0FMSDX0h/uSGgVa3nZvX1GU6BaXerWJHInhRtoAqNcXI8aQqXsYEjMaFLMk02azN0lqE1
tHkynwGmMVQVBCVT0E7cbAdt+mSLI7ouKdENacF9qxdjkvNz0DK04RDqhGhTvQhw6kzdKM/Isbg2
XtxACDoryKtHfJC2RiPVi/DeUBQvUACPr4E2f1RhYmRosw6KW5UuHE1ZjiwFAZM9LS9SeGsDOvNT
LBXBkUr2FU0BdDu9jHwR5xTWdqEunhxFoaEFjkKbrI+aRQV0XC2ShKLUkT/zYiqBoaphxgWfc1p/
Nfq+N2mpyyIyB2Je5WKJTmdZ73HCBMeu8B5/TFQD/FEi9BsZnBUwyKSSZeZ6fexqzgb+LR8JUILN
PQSEewjKw0ku5D6bmWzSoAxm83saO2XitaQEg8woZdHTRvDElBslPLrIV9/TrTRhI2HPgz+CTP7J
4v/lupyWDrgt3pZl1MB86GrCXiXcgue4XgbfqIR45qrdo+QF0ZO3JhNRieB3Z0mUN1fqueKM4Y31
IRKun/wbT1sMAvT+oj9DPWZuiNeP4wcJvfOCv359H6UiuEqxqUdaeG/V7dG/RWvCRnelTLSPLYQD
UWiRpDOQDaCLkRW1+nM6JU1+EjXZ8krtKmwGyE6EZmy0t6tnaH5iNcLPIVfDZ6/hRPlAY28MUZk9
yjNGqK6A0Byn6wumKRG6uG5KW2vGVhXr06hu8tn6YndaQ7bQXLKPJwRALGE6Ml6bAdjyyv3Z0BEx
rR04MxP7EAg+cY/AZNUIhas+48zOyqFPqHAs03pP7nB6gjUt1HWBc39gvhe3fDCRHw4dREy6LkIV
03/VFWlBab1MVwd0RdSiN19hlSebS/tEsa8HPGhaMPpgArOzcVyjzaIuxjoV6PWpcnmSv9spV/V9
rZuhl5c7wlI1RERepBBh9GOplUbsGtIDZua9HUk2dWMgZu0svgWKSR84sb2GOLxZxwTvlZEm37Sg
CJ/5UkFV6IMrdbnKq7ZMYFjMNdx9an76/7pfhhg1//vWPxqJduO7kiLbgojgTFfsCs9vjRtT8Mxo
CzPMSr++a56vANRDKZd7OJ2NES5UaRTitq+OLXANOOi6ybFaV6vsvCAFs3A08BWXzckAeNtpqYsw
oGgzJ1t7vwMvh4LPmlGFLgNXTmsjXbpwmsUPz38n/qd2mA6yaplKeDVtC2qrW9cQnNGIRANPdqaR
YEoX/kgbjhHqMyXJCmrf/+CwOH65YJWYXw2e7W72KP/R38MGAXQzIhBsNJ3kIWk2iGdbWh/h9U1s
Uu2yCxXtgYsnwMJuWCk1DhQawuCYbrxf6M93sifkmIGy4BM3WWZyAuqF8ZG+AP30EdPWkV3K30p8
//zsdHOflhwV6WQanSeVk6a6cx8Fe9GtOk5Ke5JmupuyTVY0m0WOov8tR0f9cy43aRBL+AAi8GNb
hhAsYMBb4x2yV8UPnpKhlLMuIfmOnibvX6mcYQwwXzpmZkjvHrL2Y91VHEUl1QW0hzrNVUJynzWc
mqWDCnTnyDMFd3c+8gmSwUHwzGOtkHwpT20fNgZ5+AgIbVssE7byqgDAF/4wGv2hCgs/sCPzD5Mr
7xXSBt+AiZ8TlZsWxZUYlU+oD1goeKr31hvbdOlyFc4dYzrZ6hpWsdoPHGpxtm4Wp6PnVRoCxi1g
Sx+8ueb7lSr/Omjy2hkVmI7690Z3ZwDNEF7ZvIpIYR375p8x1SgenzWaFcnWMtM7gq5x4ZDZBLOS
xFOnMC2XeB6vYZBxFQcB03QsmlgcvCUzg1deuCU7ovDLEenvFhlYG7pM9qC9N3WENyrGISCt+vy+
3Otugtm/bbhM/xBHZaJkdLjs9k9lF7shCcMrPY7L34Y/poAOe63pPfsEnvGNQxuu2jXYwJQBy6wE
P2k7c22/8msVweKCyJdNQkYJaD1oNX3u9fgJ/sdfVZc1xZQXbnBfKlrgIoixf6Ws3RdQMdYyBNfY
Ku4P+UIgWug+yyrOhM/iUvUMeh2NqvnbPZ/fMeOGC1ZzM5hFcNlkUi5HCA/MLPqoH0h45OMUwhuN
17OtkqeECTG0HiqGlTowTzCgiwF9YBiV8qQMnMPuJPNm0BdyZmFzTqMf4wUHi3qVobkUUh+RQdOJ
gF5WL58A8RgIB3Sv3NRra6HaZ64nITHHeORYD6R1S5orAYNhqzQN9h5Wkot0VCd8g7ov+e6EoSUD
aFhcZVJ2+oswy6yKYTryD+AdP7J2N9LBnJKYfpp/aLDZwt3Ccs3UmP2E/R8/GxHRFag1l1/q9ECm
/UY8JUEy4OGLl7yfqY1LKZe0yzwhm0roDWLwSplrzpbXh/fVKtkTy/LwKfcgLzn2hsdgraqxNIxt
Yd98y2jeAmtsUsueFvEMdkQvlZ5+nEH0kcwAuBjVFyigT95lGAybaaACaEQtg9zhZ7BzczhmwXdd
5FVeruHu7Czq5t1MzdvO9KXIC8cwFWjkeFt20z+byntnJ609ZvWFsB0sN/ecubpPcWKXcSnfbqi3
sWgggqxgRUheEnZcW1mShrI1JhdqvXjO/f6ouW6h6cJCDEhYjT16tbdJfQpmcghlzO/nZkuxkVl+
95sDsDQClLqgUf6Q8MG/26BXFpSPtd++udI9qckGVij+y5pKVf4ou1Vilr4yjpId/uk7MkuH0jRe
Xwos/FBFkQfoLyDMfdMxCjdXJYQL0x+z8lYVULk9yQ4QXiUlpqJV5jYo7uHiaBoS3k9TrqJpNXYx
ncjC7mbF4xvt/rBb55osrhZjmliDxGH9aU4JNhK20948HQCb4HRp7TgDA7/wIMYK1wbW2use71YY
CfvPClRzpmfnS9B0XQX8jskQzGte+JX1lZmCAWxFr4T0nyGTjYdUIU47MpbXQW7xAwIvsdZ7E/8Q
OAZ9gZtN9Sejy3kS8ode2a0RCrSGWTS01A3yJ6ON0o38iEDHnrBhQe7GuZn0yeYWP56ZMFzEbzPg
smNgV3u/uQMmt0mP8kBL/ZDs64HrmIMIlVzOqmcpjjytX4xHVLf1taJ33OJZf1iODADwxeflvJdT
RKAX2fnXQFvhvHZ0xYnitgZXB0rSpNQa/2LTZLIdo75nS/fNd8m/eZetHzDq7JOYZQn/VMjXXpQB
88VYPB2iyV8TYzoYbyBbELC4SNEqQjnyRvECIZXjwTbxfDfEvD8NTRzEl8QCcfiiwdSdSePbG/iu
AQFEJ7Qv2zk6zRCWBSNTj8Zh30/W+dm1k5qt5XMInvjM2c7pa5WqnpvgsgQRu7ft4cycUCvRSfx3
q3m/a7tzsDuMlWC74J+eieS7EHAZX1S7Wskd4oXjMpU/+//e/CA4Wc3G9R8tgO3iSoADYrwAPqbn
gCbj7RSJajmqmKPgqXu0DnWpHFu3QGMUywFoSSwJ/D802O3xaZYpQhafAEeo+XWXJgIA6fMBQcwD
mKXVhMEVYWeQSSUoEdrcTsrsVP8gPUIi+bxYkyNAy0IFgSQ2ue7kv3xlGDSoUvIendPF3KM2V/E/
olU28WxXR/sEeTm+GZ1m3EA/CBMYeojOEqktyXtQTpfhxj4ZVNrcgIXQhaBADsPiLjDCi+mDr9dv
4D6IOzfrTlcKy7PUGCQbTHQ8m7QipYUQqM7iqqrD/P4jSXGtRHgRYblhiw8fAXEAmWQuxvcRgAYO
y+sUW0f0aOjolghCOVJlrJb05uJGvVuL+MChMmegWrDYyUOWddmqhTnTp9puZ1icp+3bcPzTmEgA
qaBhN6sxs+DD/VSR8y9FUQz9nCYZqnC+wg4GScEDtEuiNp3t7GFoxRZScSsmWcqkOCqjF9Q3W+3h
EOatFKco94LIgOdpo83QEVI8aFdKm17uvo5KdPfQI/B3i+F+00EdVQ6HqqoU58tXap1/eOmoxDKb
Q0DYYePnaALF5v/O1sOfMjQvbS7IRNa99Q0hFQe692Gk51vNIhVmNm0SWinkmNpzm9QCmlXNbZbc
pqdZNCnviX5kZOVG9pH3IMzFo8pWGJZXv6rOGfrf0Xu7bqfyvmOvQbyW26CGmhOhQZCuDTo3/TUa
l3EGNakCSPKhvRa63xBD49a3675c7QDi8wHGcfr3ZM4s2N3/VL7CRst3OA1M0KUNgR5IqvfhfOKp
b7oCglp6/x8Yw24emuJjpPdexQPRI94pf3aO7LlUjbFXqY/hJh8Dc3WL38vGr9HeTOQ6SPoq14Qw
Gr54WcLwnZuuBse3MrZfzTvkFw4o9hgRgXJ99oLQ2k6OyWS9lMKCVoxdVEJtSwSKM1rd5svTrloT
jSXF5sXFtkzAKc/HQhNLFIcrrcJo6O5k0uIYQeSNoyKtloS4iM4x3yDTwXHB9F2hepMkaTyTPC11
dbcp6nLea2p/vJrXhKb3vz/S5TY4RFmdmOpihZeRV8bsJvl1T8T9Xq4zM8RDDtZzAijD1ZcawY9p
ozMm1iUuhwPwzUuLnvfFn89KKdaOPNFafSnviDSNnsmAaYMTH1tTNLGi/HrGlovwe1HOtpxWzpas
e2/GUD/KRFlzSYWCgQRqVe9sIj903QHVHvjT0RPioZXhKDEpUKS1LcpMoKA4/uX2ViWkqWognl+I
GRvyTQI+8EqZMNUrTf0+s6ciwRy4D9VjdjT2A44cd4gprH6nYpzNX4I4fBjeHzmikGWjNC5SGdAo
xINFGnGielv13DdCsFKJZS6Lw6beIzWcP6hA2UK/LKvtBWBi3KFS/gGq0EhHnkqTHT1RZ4bqS5IG
niIkH2iH+R2gfB8Zy27utHF8ye/V1U7av+qrU7/DEH2qyjXHAWLlDSC7VFD/OOzH14P0jhjDYkDk
WiZ4bMOyvtD5AxFsZGitwQ0eEXIvAKmZD3LSf9AuhmlauOxVWCpo/ZDI1YQT9DvHb/W/kkgdcKkh
Bsrd1URKO/6FFMuC5V9foT77U5TLCu0c+UwBmBObY8FFLIZS8LrIqnU/eDeF6mKDTp3dagIQlpuf
CxSk5f63pqoj7QnriE3bl6qElDNxdEOQjBIrzdlswuHLsoV8mLJOuyK8+kggbtUB/HfzE+TjXJOZ
AITB5HpNrxiL0b8QzIqaW6HCZEgNlrkXpOLlorqQ3Nl7eMv1iFYxTSB4HY1n1RQK1mioIhmWuc5g
PnB2yM2jGRthylf1RPYfflpU9RBfkxZj5su6ZUpJJOBfMGQC0iE+2WMfGMZg8eI+SV2MB7z/PZIl
cGhg/iOXfa46A1rO7tfxv9wMMlHdu0BOk0aIP21iBQV+4TDYZhX54/6W0s6CasPoEkHF+Yth19WR
SjBpC89BiM0mUtEU7uZgNj8A+IRPuleSoflrguz2BL1Y0ipQJbH/T1lrUws+UNulq9SgncT/kobQ
0dKFpNDn06fOdxRiQQBftEBfv0dFfZLCh1IsbJgpctA8e7qI3Q4m0INFvDsiNHuS3CkiPxEqbPvw
42RovqOO6TWzJvz1PslxFiO2+TZSAMj6xxAE3Y+aWo66x54kn0ZhVI9aK8umzn7cor/S/RjznU3z
zr+2q6qkI5i6UJ+YzIXxcORBIEF6PI6cWvP2Ousof/LfihvZ6cDKjaJGQQi5MqLC6XWsoQG+Cv8V
wN3LS11VTiqrF4vlidWn4+oei2HEIXBLS8gK207PonUQEBSFATcwsQbhP8kYUrPx8k6ZUegZzmTQ
3zIt2MoI4NUobDVqxv4IdeT4HgBlfrGwbTKHTI6y3VLcpnWXlXlFLxeA+UnsFn1aAwFT5TTrQCgR
8+F8/QfuctxbK+tVNQu213kZzYH15tk5Axh+MEu3vN+1rFNbQU7+WWnRb1/YPE9jpspJF4JlAOJa
ajHsNUn9ByJL0eVXaFDoKc1RKspper9wOoJMX+ZnIjWHWLdO1QJ+kuN4/ZxStGtHJXup+Eu6CIZk
0vHpCu+X+KpGvsKrRpHeldCINlXkrozLgbz2x9+xmBTulalBSmnrRAcVNB0/7wDwersQ+yp5ELQi
oB2ezXXw41usNVY8LHFbvwzsV1Gz4YZN99aevLTpT8smktDOdjvMxdbLBkFgOTa5TpO2xpkh8npM
vakSAclGtiQx3AsayWgh/HdYqYfjk6+aN3HGihL3fbC07aDZcqmaE0RsPPjUmy5L77QDU9VY4AjB
cPjh1xU/jVos4oddNwPN5UAHID442i/P5yWW2d1kOmgTqyIhiILCkP3YDjmy9KtlbOsB95bTi+Rz
KW/QbS05JDAmRPQRUMSBeUS20314/ZtqjH0GISGwiy2efDZpnxI4XtzeLxP0NG6beNikhauBNkdx
D2gsv8sy21Y2ZkLsNJXyFeYLRrM+s9bu1kSrhVMjdmVSFMlUKkaePxphmqBNCzA5RmC/WRd4pjL1
ziqi1bTKafYe2/LipzACJxy3THQMOpwTSWGtnYoOD54ZGHHKqzGUtQUMkP0aGNP3OGXKgjLYzxsc
Gd65ghwy4FdE+uZDR37ILbnczvMhZPKcXQxlsEj498HMR4QPwfwVjyaeDT7KEzxuGgz1sipH+D0Y
1t4L1hG/BsrEy5+c0ZgvqWiyPmXtFgwrxOk7hQteAYT3PACPUWNJ7EmogpacLl8b2wuKzQtBOCou
qDq9FA7CIg/QcdrZiuF1FumkqvvmyYR3ogddMKLEIzQKI0Tv/fueGutJTCjhZUbI9lNo2W53IS3B
HhB8gmTqSOh6eupzwdRxH2ZH7foHNyI26uqDZmU/ig3uQSiqfpYa17StNC17Pf5cGN51XNngS1YF
6TsNMRiETPVHHZ3EbH3HZRU0/MleDZVy034ZxNVMZDT/MRn3yZ1SUgO3DgBkHYTuPBMFNx8vAA40
chJTwgbceu9gZlAAO4GV4tY5n9MHUcRnB1RbOk+Jc4NTr7QjOnYd8fcADXU5fP54rfAeDwTxOCdK
s7fPS0JYW8o0sehosipGrJZ9Ol4pCBSIZ/gu8xSNG1XyFjOZmwVJkEfht4J15x37HWdIxIvLNrOU
a2Ujx2al1YQmZLV+CgVGSjw+3Lh/r2GDYV4EzPMknP8Mq0S4kZied6ToD2YmIZs/D/JaMIiUEwGL
aW4EcXl+BdKNQhydjRVYU3z4pGS2rJAG6A6bmIZ9Ae+ipX1m6DmVPFhJg14AE2EFxPMWUr7sB7W4
2rOP2f6M5mNKswK/l8TmBnhZhmPUEAX7osYhiOMEcKoD62G1O6OYYSlz2JScViLTHo/odwlpbt+l
5e5KYIUdVrntgsJ0Z88CGxk0j084ToFziWYu57Kwm3VhNemdX9kl9SkHXl6lusJpwO9aUAVxKp/R
/VQ4XxAZu6C63DBtcehBq+gIc8Wt733uXfPC5Bo530UK1beaq2tNIi+ihiXzWU5zomHGu1GHsoxX
wthRMH3LrvNa8dlpNkguN+Zgfmm+l25UwJe6yIGeo+RrdnX5VdVbC+IMRc1Pld32QM1hkNgnlv8J
9r+l4WiZSBosvjeDTHFi4yZLcc14hjswSgOIwVv0jsmBbHFtZ6jLHdMZtm5czT+kUuxcUBxvCxLN
ll96Ln3NB/au+bFPG64Qluu2eAwSoLbLr/JKelmpoysNGFd+LLSyWPp6skjSIcBTmEJ8G2IsnVgA
tgh0XHXFR9xhR0ZMmP2a4Ov0cd6YBBv1Gzc6KgKRdm5ZKPYDWc81q5m01AT5dDOMkFXrLudw8Dr8
oVI3N4BZTVLAXS5apDlGMddIxC+1TxR5Rg/0S7+kAld4Lp8UYYvq5mlNIo0PyyWdQAlHAlX/WfjP
OgguhYGW0NhiDkYhK124+44iUQJU8GnKef7uUC9EN3kjouqW2K3IB7t51HulYRVY97mFi1xTN1NP
isxMfMYXTtIZCUkXeC+FAdYZWpTJ7Fof85cZ97/8B6obFB1U0A9gT6FZOMexB6LFEco/bOGGkcZb
JkdszxDToWl8KGQaRe0ZZffFNXCZjos/OwLV4Bq8/2Km320Bd4j1LzX/75pkd5ttOKs/jLGQZXgN
C728Aa7SCQQ97w6zEnqT618DQouOlH1iSC/qkLmvi1FVrF4xs6OwDb+I3mTWkIAt9JvhSBDv8UCs
mS8ZsMqvoLmF6U3dKl97M13MxrLuX8hfUbjHDaB4QorkCVQ1NFYh0SclcRJI9vmS8zPbcV4I6gWp
nMCT4SYTN9qYFHwu6mV5fxbIN/8gWO8tXVEa12CyeTew+s2M2JgYXX25490xxHUvBSDVZwnzvliq
1B95KlVxxQ9fstBAj6/gskABN0OZvKG5p9Rc79/U77AiR2MpNXhVf6b6XRxKvDvj8l/L1FZmDOdX
Z6pt/bg1vaoH1pbSUA0B92dDQ2B2m3TIJoGrhO0PQAsB544GU7kxm2oMXUfDlhaQKHiS9ZhMkk58
629A3+VS54dLn8b3NrnfyrfOs54ZajL1lc+JVq19FUw0Q2ogvr0N+6UgbKTnhcCVqWTOdjGFdEUu
a0opdeEw71EkOzmx+gQ9P56As0dUSihiKhcL8Oa1qP88InNUgnruTUvu3+4ZETMQkXUOhxYDgLkn
wxvMmQAJGwkdkdjbPAzo6Z1QRrTvhJ05gViR64tj8o/fZSXDKoVvPXaBxeU0cRffMjeIpznwlTid
/tL+LNMdxZMxRRiLZ7Xpz8sv7RTwt17HP+L7DyOWBwPO1nXXFidPMKuGSsTh2B81ptZMj3e8RvAE
OZs3nYCuVG4QdvRaRivOQ+A3lPHyOWxLxsx7vECd/QGlMiiN3bxDh+nB9wy4AbZ9XlT6k92iQV3i
DXtewVgKCGp1LMw6v1fiAcla0+mBZDvrwE8xVn266dv4v5X1GqMAxYl3xRaqMO+KOF++1qmRo1KE
+FCbiV2uXAl9sNBiidfnAYqHjTS+f6P+UbtNkgPE/ixVakc2YfDCFi9dZMMPzLG1VVA3anD2rmzm
gmjbf6J4dYf7HD0geQvEgqA7WPJ+V/8/6l2zyyOh2QGVzaYxqIS6FrdBsDqXU/XHCL9vJCT/fDfN
Q7G/QhgULfzGZLO7ChRa6Gagk/1chEwJrzDkTQk1DJ2GrK+IriOc+FyhIawFNs73v4Hrj20qZI7l
2CGdDBlDuw7sodLRVJ9QMixIu8OlctOKSuBVNsnA+iZe5OJYkjb1Wp4fQS0vvf3994S3LVSH3k7O
V30Nc9cd1Wjbm3doXapvLRYf+ql+2bgcqCqFXzzy2MmGtorTz+JEc88xzb83ouspLS0YlNBsuCAY
lMC/fVPc5zSHYH89AYg1j6HfWDTrl1XvhLkQLO+46IrMvMJcM0qnusTAG2JIkuUWmmJJDOT0tEFN
JfLK35G9BoC9dF3BG/x/Bi6g1Y1xEgzubNtUmf2ZUpfuiIfFWEemxIeE8Lfb7Y/vpqHR3x/Y4NIG
gcpHwqhD7WsVhG980SiKYmFpUbp5egNdXJSMhDqc1ULxwFAG14M1FOIxmLYhyN90+EtgLeE7HCVR
+6jVRC+WA2xi7ZZm1qzpVWcl6KBM/F0YKDbcR3deKYcqsEDbcU/DABWtWWTbpDrCu1XDiChcHAhg
xxDMvSqJWjIDZ9A=
`protect end_protected
