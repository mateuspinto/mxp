`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 98560)
`protect data_block
0USWSUGxovGsyBJteYpEocc2z7dSGq3StaT4cUrS5iZZeactdHia1f6kqYgTi5RtAokG7jbN+akH
Y7IxiSd3VNFI+Err07xg058PDbbP0mPJIRo1Z8zMin7Mdtr4RWrd1MU6N0afILC8H0hobfSFOU3x
FzxaEXHoPjAa0JGQfn6Ne5B9MNi5EQboRYqAnCMycE0qUKD53qlWpU3Ife+baKoMoV8sPw6oCgmv
3fa+6QIyeprWB8K6nL2KWu2TkMmjp19ImJKNpcGrtgncmAzLlGhA28rZUR0B/C3MPC+9rYKNu5WR
Qyhc4dELi8WgsIiCqYWJMfI+oYyUH6kt4K3eGIwhc9FAfThDMdIj1JpwoM3MkTqXGMZR5VJ+6dGg
X5FBJg8K9ihXyTga4mmqnFqA7BXQW7kI7nWfNQzryxHGZRdUGTvPd+xqIvZ5JzfmHmwpmM0TrO7f
nQW+d/nEHHYwHggXXk0E41jJnGttRtf3R+1NxCM+NfvuejtNo1n3zfoe3iBvYPxwc2mrD2ZH7lEQ
ESnY0SFXn+shquvtL35FR+kpkrHUp5pz2XRQI/SeGJx3tr5XHr5V4M7bhG5aqVUnHBUFqqsUIoc7
LXjVg+eboHC01f0wlUEEaEjGSFAt2TObXS6t2S9g4HQ5GloGUEqC4yEdHF6HYpO2yChqGJu6Y53q
EtGNThlzxtN5+7sSDx/ydNQoZp8NvopxBlmZDQQhraDJqZKdZQpP+pTNY84z+laNzVCBrv5epaN6
soT+/zu6WC/CEndVSq4qz6mvg65QhPLUHawA12Yca3klJPfALC402q/XmvcZL+QsUHq6A3OvRSu+
ABmcU6z8Aq7cHlJhVZyA7WsBI9TUx63v+zEw5URHEWp8aRrihI6kGClNANx+l316xDwdeOwOrfbW
I+QQEs0sZfKbdmdrERMvDGFvVAm2zBs1dkb5SsbEDgolLoAycUvDtpSpmx6aJJi7g2mtwESLv+GF
pmFYHPBaRKB4nfGL1+NgPghBCj3fJIUFTz35HHb8xZCPwMGQOS5/h0syA+Mx1TJVlFwGUHS3Xy6/
76EKcZlWJcZbmRla0SDyxTYb8HLk+rSIHO5M3/Zeu8p1RoqYh5GlLzf87EPAtsAknTbjvUWKtd5H
EsmWbCyI8UsajMGTXBVmseh2Iv+VcSXppAdIR+GclObwUlY9Buc26NVTQhbQZ4O+Udrp7XaEo8it
S98qymWON6j/t1mLW3GJWPIsUo5F1knjNp517q+8191VB75ZZR4NcuhkrpE85/Wq1IudFRbpQIvK
koYfENvVhMNj0zp+q17ywLr11GHOcoVsY8kP3A7Kr7RJT/nCQi7DTOtUW1T+68w/9HVkaLj4M0j6
F/NNiGCqGKy6n9kHsGiaEGOdc8B8cKpxwwuue26U1xZYpt4vRaqrjuUbQGagtkdce0LwT29ySvrj
8vquwb6Ahslshy/2DRDMvMACTG0aeoC2mgwUeWofCxfM9xi0WPhyfXoYukkqWM4lL5Qv5c9sNzKC
xJCIOFyJERSKKsUkHnCIHXIgUB11XWu+ExpkbdVJd6yyO/8U2wvvMaqHxDbTr0Q1YMoUGgvOE56e
Ujdg3uf178WLanKwN6C7wVVrB/m7SMaMgNHnjdM9EvLI5cCQoCQWsk0KPqY/THY1T1x6Lrq7tbOM
hnz9JeL14p1+XpyBjhz/2JO4EQufduuBPfguKNQAWX19e+yVLmkbKRK/zG6rprpdBxx9mX4ML6E7
cWXpaIMr/wUki1nurgg4G0OL7nezOYOsQc5gA88Z4bl4bWxqcDwL/Gx9lPUKnw33TAHk2rSEWxgx
mjXZdRHGsl+fGZUtIBOxq6RNxycMszFf8qui8i4JCY+Siq4ksm67hiCAg3DhnHQNlCD0jfL+8ekY
ligVJ6wSs/Kjk0n9/4O8tbkneyWUp7zK9MEY8Wge/igOd6A1h1faQj2IDaOGqWvqZzKcpXtXNY7Q
ktsCyxAdPdh8UjwXbhy7u2bQoHLnqLwZIjXVHnSzZnAl5WDHSF/f3VJnFNIEOSsW5p475pev/f+X
g/wEz4NueexNYTEaqG75L3A3iCHFWvlEOaRA0HBgMB5Z+AMomQeQm7nOj34erU2I46kYH2H6d3Fm
vQYSs8/32sFiV+9vne+31uhnejVfealOj9ef8rlpQaJ2z+IbqbzQkn9ehm/ulZaI1xn7AeiVlJ2J
War3CexEwJhLLJxBW9FhTfzf3zvcRab084Eaxe0AxsH0lj/XHmnc+EJsf8deQL1RFLB2z0U1JGCE
ihJZ7bOo9XcmRM6aau62YKY76fdxCGjCpjIzp7MqImMzaEUdzOpBeBfyF0oaoQHaW4rU5cvWHabf
zWYNIQ6HImJG9cvaPtgkubt4KJB6sp9VgOIRKgMKhVyIGR/mUywoPW8/KfwWIfGF99/4U4U70auc
hAkahhwNUl64TAuoO4yaiZsxdv3u4AG1LDX1+QFWDGWYp9aFrqeYBGgtGfZiI2WZmoQ5za+sh3BS
68EKHl5loTuM8phyUHpa9434Pa5BprmCI7/tpG5KOWBZ37A3yIUhXEGx+IvYAiP7M2jxiAP7p5Ck
BBVXKcmfyWroXJ62psjg6p3r0Cj+vTvhp0fLgEM9SiWTIJvUne4tOu2dJgs7T8emi6Z3buX5TJDB
uG662IZTXIjanCP7R2GycgMX7Rlt3vorbKElLCrOnb8YJM1OJ/JiOnCWq+ZuyRtAkINBa6XpwE3k
/hW79V822Q43Z3OlSUE4zPkoSGvrGcF86RZ2Xx8pkYglBWZL4sA/4EDEMtCZcO/cqMJjTO/MYy9g
zTJsTYIg5wPbF2551gn/HP98ABrHRN/Ty25zq2RkyiBuw7UVVjYKEcyg3C5EknLcF59VQEzlC2sK
jgiAwZQDWI5+aAuy0KP/6BOhJGuoMAk2e3ta7l87hk3LKHw+EvdB5Xae1i74agRaEjA3igv+YaAP
Pvw9SNaBGO0mE6l6nNSm7Spk92kR37D3FlGpqFlE6cAr2XvbKgpw+Ci4hIBnqUrKHZUICdPP2GqX
40vdRIqbLIOB6gR2QIxd0w4dNOb33fSt2/zDg1byg9eA+DDl4H2tU6QJRtoftzZ/t2ymiKvUHzKQ
mCNPjTOrOGXeagt1CbMCSkQy14hkl5ZlGLsltsazBxeBky2yKqv3glEPVeJaSsHFjGTed/oXnGpI
Q+79Cuy7/+wZX1HKorSof4LX7yHru9GZkW3i2UEN4rEp8NXYFbd334HUi9m7NVWGYMEZpIwkuyY1
O7knCNbWKwJCjb9cxLb19tHhWxrc9qaSNf6oTI7jy8ksXVyDj7lqolXxj0RlZi8aH2RCtqmiigEA
abl+4lTuUQs8xDmJGA5FwLN2VoM6oxVDDogB+buJ7xCtAiK+jKPOhB6K+psu5LQ1tjqdNfDZ9apl
a5QsnySdjwaMzxA5jOqQBustRnJSnk3i5FIZ0AR62A0qd69pVHntZpe+i8o4mo1ipZ7woAQNcnON
ovpXN7cvSiPf+Zw94Nq1ZXufgg8aofB8Kehor7p1DewchPPoI3BkaswxeX5A6DYbHRvSkFNwQRoT
lb0OQ6MkTykDEKg70ph0PBm4NPlCuA3G8pQlTBeO2j5C+zCneQ0RzpFqSAWBN4ww7/tRRuOciLmQ
gLJSfagOZFfcTYleZ6dVUcyt47svhz0Ie4OmsTRxeyt5D2I02Mut0nR6doAdtxnZbN7h5XRWeo6E
cse+Cyqu11UwFo2SLXtrZpgCY4KXEUm2fa9seaCFYnBe4260bjkM7oXDwbWzwEklY9gCrMinRzIK
NXd5tNDGfCZCU9fubnGvbbKC8uXTE++f+6Z/T7kiFErdEG/qBlIUSPEn5AMdRH19wrjXPOrJ1vd4
amUdoYh+zANt+mNGPuNdqCD0sdFpgI/jLbuU9+vaeHJ+1O5VepTdE/mLkVcjw4Vg5jtfzQbi1CPt
ccu3/hx3o7/zXUfXKOhssNL+9nr/e4wnVEyn10bXxTl43rMTLTuo+NqHQ2in3sqvKD7qpw2lwPsw
9SKpuIfaQafKNvWkv9uO0fopZVO5WlLP3Jp9wighdqBoiMsLDFn1MGHnS8D23zcT+Zyb+EY8tzqN
uJ66D5eZZ5ssDHCElDD6C6yeSuPVu3dKVhp/n7BpDLx1HstNvun/L46xeSVbgaVPr1OBlpvusr7g
q2EtUiAA4yruyrBMBX4D2GlA7HT2NHyONOWo/EIXoDfXm8FVKitD3jKySbUFaKyckqecRYtTRByP
7H04qomdzMLQQERsaALTuDaNh0tfiNVymHvZ4J1Mx5681PBCg1C8uqtYbsSuRw984dngbs8HAuvM
qacLuYyURYLBv0gNKummQstd1REhiv8D4OgFi67LoPXZMxVfHykHVqknFd6TQ9hNuGugabKNdkDJ
mAH32xnNNTqVii7DZkpdcXYiJ73gI64FE+KRaB+9dTGotz6vt2Ov5pTwpSm5Wg5InYGWjsp4OIj4
yQAw7CSazGMx25ziZAfeAULVyWgecUhU2nGDhN33tIDAkhML0x8CajHtizU+gjWmu/sLJpHDyahj
Ifb0v9yqEU6VHnlFtI+rKZ1IhoT/jV3ArvDU5wQxzOcnrCKWVE/7Lax/YDkV9fGkVz9QE52KI4Y4
Nuo1ET6atHemd1mEElFhH3gw0kg41o8HbNt5yb3kyR719aceGXX/mZGw0B2MVrVLBZ6SRXBNgsBK
xufHTpRsHLSr6qLrKjFdEZdx1GZ8jYL2j8hzmWZHBray7W5CIZ19SDCXPC1Din1pLiaxf3VHbFad
xTE4PQgz7DzbqsqOmqXhrIfNx7rGCnm9AsyYI1tqPSi5m/UjJqP7ZehiHLqZy7lzCif3cqh+0KNW
tHAN6RvpEBN1PmXJpYEkuEWKuDJmcumtULCQCbous3nedNZMCevnbNzmpvcQ662VxEWuGkpcdyj/
ORr42DW6y7XEwDk5h09vAYn+28p5ko5kWpJc4aPt59mJHUzae42tWBA5PkH9QeVmvFk6bZ+t107F
l/o1GO+GRYmtmpk+jHYKF3TOsY90sn/mIeWjYIKta7U3fXzGe6jc6/7ccDgTfcC6K1RXvGBtVoPJ
zzicqP/z28deYOWqILgMxlgj+3uLS5mcPrOx+hUZw/28wu4x5sID3wR6QrBo1BkEv7DvTlyFEHFL
DHYmmxdYE971PkWFsavOsSGoVDu/kpi5egZ1555B5SY2A7dCfOt/4xgrANyMkb42tr82p444Eari
czegtgcKD+0sYMy/Z5jssb85KqdaMXzbvGv+68Pq2qLSqw1qX3A9bUIY0yjkURzFIqmX7OE5iMdK
P+aZ/rZhBTaqZgeahtGbHkedEyj05zbqvjMoujfrl6tIkRI3R9UsxTcg2/sxTfCIVY3MXwE4Rpjg
hq78+uDzma2I0YO7QQ/YtYiv9Tkp5EnG6LSWb6xl/OtpJa0MFO+NYVHyXNczu9+u+LbiDcvmAb3N
gV2UMZMnTZYOoEDukPPmk78m60ZpC+FTIXFq2+6+cdKrFvHluE4cqMwKqORht0u6SnkMp3NkYy5p
1TfWCILdqQwis3wlBhDQA5J1Zq1rbzfGolgZcLAQRb8d4x45nPEuszvDk5wkAxGkbNT1qDGS5zqt
j8rOsKpGCMqa/gJgczF/RtIDosGTJuSClzjjQv92e8CVzLT09O0ujF6Fb9KzZ9jxiGGW2GCSTO5D
wdUqqdYAEeaGVGxiCUg7EtNsqQjVulAkFrytbIGd9wVzmRDtINkj9KtR5Ez/8eQN2MePcMY7n4YI
AyV1/ZN7lfDks0FWuZammNwmOfY2p0OP8FxWowSJDrNVmdbbfzaMuHnZSZSN4U+sbzRQGFS3Crod
cjaadxnvp34MyiqeVRHq+RxPsJ/XbQgEisj07uR4LYFyP0Pc8snVzkGStChkIRAA6Pru/wo1KRZG
cTDXRTpmwk6my1oIux6TD+tB9yEMC2NfJLJIPcj/nbfC+Qikhmgeu4Io0uxoG0J4wcc8DrDRKUAO
AaFYccQaeqgUEAKqz3KH2YaVnGqzUfFecGRul7NqcpZmgoajizpIgUrCGPqMl9+KfzBubtjsWdCH
/SNWg9xJzdu44FzOZ47iIqx47Uc32vWWi6udkFcZiHPMfr1sT3Ws8vY6yFvimbXqSf5pRWZAoZpj
YqMdxz/Yg3oNMtjj8kZ3nM6I3FxLu/OCrhID3AAXDSymj+IHPJnXeUQDUCA9fTLzJiBQnOa4j7Bo
l5DVI8WiiMO0eqlVfsAT0V7XiFOA92jC8wRnHBBS+/GcBmO9cQX1/Ifbc03iSDTYywcY5WtiZgUq
xRCEAkXpiwEil16QL3PdO0bLiGio5FepqBJCaIZCTXrRSK4BN0BuwFKljcXKjISsa5TOmiMRyu7U
D2x8Lt3z9Jn33OcXcf7ia7BkR1dCJUnco2Q70W2/XwNuwKbT7pqVWoEjVoviBFBMP0Eyj+4NpM6u
Fg6p/VRiV40X9tudvdt5mJ+4m7PfWkd91YEx7p67KwEc0iIBtWcdelBfJeTcAjH2bB7kKZOwRQ06
69e0D+xaDcD/35twUTtgagzrjUnhL5sMiWmgn7TvD07VjmKPw+jQQ8HUyXolzNbwAmlOu9dvnxBH
Gqj+a6GdvkGvkQ6Sa+8RyYpTGLI0dxvx4Uh/qi2ctejiewDqfA62PgH276TIFSZ9OTuHy/ONxX1s
la6UzHunTenBf9gWUq8DFIdW0424CsimxjXM5jtFj+KDgWYd8I7xrXra8kdsNkLR4+pq/Ppn4ysP
r6CTcSvMP8Cq1/rM8Tvr1PpBvlWw8NHGE+A5Ufrp6Bcr4mwEvPMFxbB8/zDUxY6iOSsAiCJFb9gS
hrFi9dHL9nST9RRHHSBlwPe03YhHTEMFpw/WGHpST4IUQKX+Im0BK8b3JhHcEE1j/RPal+PlK+8b
yDP12AvE9pFx8Gnh+GJWMlYREKvSjAb5kwHFQIBj/K62JvTduG7UvB5jjtx8fiLMpk6k0h4/GYoI
6vhc998mNEX6szlrMYeHNP4TTRnY9zZxk7hW81DGIT2PTEjl8OyuK0sYQAbHRtar5Z0IR+6qtGbe
pPb28WVx4zLLyVKQpnECCPaxlZxEqw8c4XOCnlSn97Z5+J/1v6lt/2yjMna0kxMeWOnx5j1Jy527
8qlUQPHQglxgDMFT6nMXHyUbGZudAaOiFIwiyKm6Ez/iVNVsw0Tlx9NLKfJR5AdHqMk/0Z9drWXK
jcuFviMxO2bZV2ioXWVT1hUkWsgvVbBMCVBRXU29AFwqjR3OkNrSbwMqF96Cq6dPncbnPjm+LaHx
FJQ9QNSPKOgtqG4lv7Ndxf3ueoQ7tph33lKLPXIJemqfmXuckk3zkZa+5JH3xZKj8TNA3XqklA1C
/Yk4SA3ROi1QvTu2E80utQMqxJq/wO52woBKaINGfTiUAotLb45gffPAXXijZZa70xuc47nLRCCI
UrRTHr6yjd5CyYUtL0EkxW6SX82MT1PA4S5CMAjSNwU9n1oHp2YbiG6qgVBh6p3CL55+iXI5ftjE
awBiu2d2R1LENRWSLgBDdbXNomIPCpq3p0UrGvuGQ9l/WE/vP6+PxTQTnkuXfgwcyUMCKVipEYbJ
vcCj5ndUuXXsJkkUMeCEs9D4JMffaOv4dd7o6IG7JlRZBnez8boP/lm9aGAcGcdEJ9WvEqvcOhO3
+oaPavXVH/qJ0Ibkwhh3CbqpDTrAAoR48ZEPYriR6rRNBTyjgiSDhbpV8aUSHdx+W/y1SbZT2TQP
VtUsqthZAJxH9WkmaAbRHuCeMk2EWnaWHeqIhzYQ6tHZ7tmnAwzHVU9dD0Cri9k28brpbnAUcJYb
K+N7m2ns/bY/pdIIlZis/h+/vACGMzh7x3WWWJRmqcTQgSxQbUZ7rsuhQkXRMgKvwr4W8+FKosm+
9cVI20Wwep8xwDYQb+AZx/icAt2KrwfbS33xIza/+/U5jADykbI96hajp2VRCx0rBfTO5X/GmZHd
MSOZSnsKQHVXPR5+yIgZQJFKFMvz7H28gCzpTVWu3DfmwCIJsB/O20nLK6+0KK1W2fnnSqmUB4T+
KyOJF6e0Yg3GPPsLg8U89pielBJ28XDhgvLRZqfgoy2jYVwEyWJn0mpfokDCROf/nuGeo8+qdX6A
slhi4BvIxcEubO9lp8vPjv0OBrSyo/H8p75OyRO26vGC/IU0TNzd/xwJ4mUYnS8wlRJMI+oYIlI9
jjbwNC1IkVXJqRBYwZwt5WZDFOyWgxedm5bzWbvMhJujj5zTRKEsbSmgBhOSMRqnf0USV4lc5Kpl
gWSgswVQbyj78/Wdu0q63leP2PfrVu0QrPUwRHD6hrXcwmQBIfTFmI+Z6jUtulID11b2TZyx6YZH
vRCXdGEz6em3FWO9PFOjov8Z3EMQ3bI8bsKdX4LTvu5R4N2cUxuHtezb6jBUxFM6TnX1n3uLITXg
369VdT3dDgXTpieIX4bJH97jTF8+tfYVYAPCtu02fZyXDm7et6T/7EcKmi5Sn+MugezHdPL3zhIF
hdnXwH3xqwbkwKlpQ10jLTxDMySw6ITfJY85br9oCMWiFgErucMZonJ5AmpnePui/wCXROCxEOjm
AlYD0UA5mlMWfSJWWN9QrMFx7apm1LNfMwmpf+ZflkVRWNKU1ib2w18qye8znRirK32TJJCN4zKO
oGNrJMtN4NrkVc3Ud3EXRJzt8tK5rCcyl2WzqIWSssfZ28oMLPZgwjvVbV/C/4IUlH3IDC9lu6Gn
7+Z3Lus7cT/fYTIaBHkoCV2Yb1m4XIFcl6VsFgnUnC3/enlld1xTs5Xz4kODouIU+fHxrtohq//Z
IhzulgiyBXBHj5JfgbvsOPgKlvjbm7D9RzqapWFaKi6njHWDLulH8frYyqbJHcPOlMJmz3nep4Az
iRsVVBF2uo+ineabyTQBM/JaR3qISBtfYk7//P/9HIdHdV2l3E8vgZzX0ZDSC/o4zyzc200aM6KD
KanCO/mWXEOIJdh16c9fYcR/hxKQ4Di9QgmrUac1NtcT9zV8Dwf1x6/Gmnp1oEeax87R9mJcuVmX
RVACLT6LJyuDMXwEaRlkhD9cyRWHZeWx1TFeKCeyc2GqRz+bt9TY2QFn/owktpm1xkFlTtaM/Mwy
U/AcCUdCEZtMWY3HF7qNNjuKnDZxmQ9wu9F8iDUvznztjMIH9RhbfP7eYb873Dt6G1mPiHyxdQ1E
wkvzKNR9BcWZnlW92vTMCCM1nIrmugvFX5ojp3Xnx1uiXIP5Mya92ds4z4UJ7xxKTWT1r3KcSPMh
BAOTZw0CPtb7ZjDZO1fY+k9h529qMmeFTidFRq1gVM3VLAFofj/mjDxE1mhhG2GcucBtf25vFhWK
QFgDxdeQNE+OAtkNk3jieGyN6xJF1Gh+qHDnxXsHmcCteDAVXH5qjPA3k1DUaeqf1sP0qbWZ2hYo
t+5zs/bQ6y8RBXk0RIZkaB8IHqGPxNzeF6VOyPxHGBSVD8Qxojzel0a3gGK+oPDEb122gheh81JH
k1Uc2XxWkBBJjD5H6lBryC0WfmOSSV/NXU1WyLB2O8Ooh1wTjYKEtJo9fUdyRmHbShk++lSYlcft
QzZFwuPgkOKUU5ONa80RYcDhY2MAd4F1gBm67KNg36QNkqHIbDy8B/Wdklh//rOb9LqI/PqAc+37
E/OCT918blVYbrHWXoD/AONSvVKWtQNsCRE25rO19FnBa/aVyFBFHN9PRvyQi1GUKg+ew/sgOXF8
7MQPjI+3kJQVooS2vW0pe1c5ddooucTfXURo6Q0N8RekxDThQF8BlWIixM5j6vMfj0scyhLXHxLy
qN8c7zqbz0xCqSASaqO3Y7EN8zUJOvPYZnDvdkOHbHEQ9ULHutvrIVwcl2VpVFDwuzERujZ3759F
qLNbbjA2rrQhfIO9J8Ylc2azVAYdmakS/CmP/ZXr1dboAB/Lqk7AWXo4O6SDp1HwD5oUt+O1pXGo
BI6WhyQ5qOA1k/7stQuitqAp5xjS91TvMLUn5NQNjDyiAyvCqL/Ro+0hasDI0Jp8TVGGdmNWC1cU
vvjkFF7YHAkylsvCUzIu8Wn/vdAaYV+E7sKH0+KTt3FTQVz2vinzbYD1wj+fvJb4beC2Cz6bGuj3
O8pYplABkbRrpyUmCkqcK7tIOz1v/RjnHQdIdsbrV/u3NWXNkeaRX0jO/4hucgFJDoK+ILGnwCxn
bA6/ZKts7ReT+YrMOeX/SVEa7BEL9Zmmq63MToUVtUBdtYw12g81iPy5vKnGNmuIk8Qz0bzmRIPJ
cBUWWNfIaDCYHrnbyXYluVodK0RmHSaregArQk0QAbngQg0KivgPwt/tnJGV1/qjqXLl0yS1HpIa
GvpG5UQy2gA2+r42INL10q1GtCHNCt+Q93f08XHvoy2Jtn5CrhEe+XMtAsnhTQUCq7sUiC65gglY
nxw4E5uueUWsO0hFYAmVpgdHQqOa0nTrAjSHVgCodnsc1kPHU0O4UUHP/9nlikbtrKIOLpbbQWof
vx8pzX2Oyt23hgooHeCrfIWMhL09H5XzS6jD+NN5MYyaBPwsZLtxBeG4P4KQLed5PtZ9u32tg8AS
dICamaGDKrg83eg/u3QLjpDq1xk7pQqa8fudf/Gy3P1ydp/ceXDCdhnnkF+Fl/V7Xpp059LpyIcS
eG0dDJJyPU7ABNOmXyMxkKOTyYH6klvxnUfbc0g0gAxvuPnoe88b1Y0tIKjgyDznwDoOFdp956I9
XbW43jhhWqNQAIj1GZjrt0vizuOTpdfrJDkBFDQHaMl0KKxCT4Tw0/eKYuyenvjaro4hIusUxX/o
O+PfHG4A/7O4JIkSRNDn7RVs/ldE55ESfb1NtAmdz0d1Ckq6HX82aTf0H/BTGSEaByXhyndysMlj
2sZ5IOB4VQamdsg4tueSuaDnFymCEcGy4CrRRqdcK7Zbu7sinmy3o7RQWE3f6ygwt1ddjfgPrUf3
0vqebBQiLhkDsmX/7O5JExrRaiRx7TUUjc7SMzqySABMoVdVXYxOdLznsIgO3/r/Y+YJ9KH0IxYb
d/P4iP8FgpBh/IHwlLrg/kFqrkP0QajmeXPdVbQyL7Zrj3PCFXuW7u0IdfdVxyAN6HvrYHjRnXdv
pIHrOHQ4ipdDZ+40BZzYQzjK5ur4+U2zvjpGGZLyElJW+0VDx8NjJiMK4aM6O9VkLIODCD6h/bxp
/Xk0f9lbfocv2cU8M53hHC5J3yvwO4i2xB1o4woP3ipsAU3Zxpcm7BmS5Bh6Al2YlqBGR5zt88Nq
DMSu2HLArcCXFBLhyjNB2MLq5pBMr0MHS/yYa8gSMp/3qTFP9V7p5Dtobbn3p940TdH0Ms3c+be3
LkyyzjFrbHqxEYBYXkbu+tshwoy4jlV5YP+c0dD5qZU/aFT+Q2RhtSL1s5gWVTp1DdZmQ8nQOXdc
R1Cld5jMdBx3Ql2xfoqrs3FDxka8r5ZYP1cOxpdgLrjIvQVv+CgntV9pn5KqIJdjFQ4+7kAbNTd0
sz6INFuIc/mt35EOY40nFk3aXZZwkWRSwXVWfPaw+vDK8KZ65iGpU3C7rGZ0M43GTiB/vailYYwm
/mjNkKRku99AmoTXsDD42LNZSu950gzRi5eTx9EHlLliZb/zMdwwIUwqWpwcwI0voLQar1FYSeSF
gdVIojvPDvc8mIEcnydWU57WG3glxq/lXs9UEv3Ox6iVwejz7Apu/Ta3kJcXFUK1QFWzj2lM9ZvQ
b7yBZ4sEk462iCWO1yb7wCRbIjbs9nmGLWI3N3VdfA8hn4PJGDlk8r2qLybbizrjBUZ6lvXgfkK4
/DI0W2ZR9fmGoPkCxlSpIDT228hyo2lMXEnZz8PcTLmzNtw+nz0g0xIm6vkwkssrETESn9bL3zeo
FxyWld77XI10fVDff1VoXUai+nZz9PokP7o+xeuR0IuQ7AihqeG9iwOS5iPodhxMZuikY+mk1b7n
7e4dmCQbz1TNbdpg/Y4YfphVQvfdkKdQpUAAb9mjZUaA+URyCnGv4od7Ko0cegC2i1G3tjW5/9lg
UU9p10WeEgG4j2kibmWapERM0RE+hi2QjRZOKoh5gLVC6/+n5hcWk2WvF3gR9LpDjQmyFo3QUAuC
Cc3zO4RvkhGrQCb73kZsnZZKVNHrdAK2eWQ5JHQRkEYdGxYHuaGg5F9DXv8qwtH24rBGfni51fdq
16BxdRi/d4Gyf9qiLaczQFCwtn/lJh0rxEhQhAKJb7CGliMPXgN4ZxmFs+hC/EQ8lzxVCXBkeL32
A4EImQptXsxWaPw3q7m3o3FFsdHx3gGTEMEFFl2ip0gTrV2Aem4xFC2EH6SF6PbtkWAMYaxZf6bH
g6qRbxmaUdcu4WTEflgxvkuU+zyAUWDjBRFs4bTHHsgCwoolNY/Y5RRZzcSfquLLCu04CAxCRbLD
AvrYH/vTtDSG+hZYhQUakkQFgSJC9U1dEyIeUndiX6TAj6uXm6jxZ0GdKaYkJwCaQeDEWmZmVXCu
ptbaf/jiKcH7PDLURab9ezhA1WodqTIqyWJTeIlEGXRP5UNPBUc/AQajQHW+UGnNJPi18cfwRFRW
0j3shp3JSr4uL+quTDVonbY/YaryG7gS/kEcBlcPf+XBOe7y2l4xTlOv7RmTGvkN8VabRvrXuqo9
oG7nOrWzUEfexrKlXTs97q4ghKlegM2b+rBblsXhdAW+uBQJsRVKXpUEsQTxrUlNodUYIwjFjlZk
zXzWxpWgQu3MN4K4e5ZNJhLBNsG9FsWnm3g7vL3GApiw5JGyWTdWC9x+eWqayAkD20rE9FkDQhFD
lY5w5hhU/3s8y05rdccPwd9OMJw+smaQMxo5Uj6sq7ZLofeimK3mmdL7KYsoMZb4PYLzqOegvVe3
jUkzAm/lmtl0zqR1PhP3AQtN/2w+XUsLAaT+4D6bJ2MGDkfXj1toFodB5HRqFUQmZQTOA49gScxT
cNxOmsujx8WgkmjUTWKFMUtqq4MROVgnKiVeYETe3JMi55vg+Ehm+wYTURBkfE762a6uE2JFKUgz
asURj+NnqoAJQZDRQjR+0z7aq2Byoh3NfBxNz6ywLeRJk3cJpqMTDQbjCSj2gXyJAEAMvjlnKTR+
ucgt8Le1KqqqQYiyFG/uRXp1fFkeyQKoGL2507WdN1aNKJnH3TqADmV0HtL9kDYjkM0kMKKI9KjX
n/J2maCQA7YwQ2bkfv0r5hNCzW0+Nnps81GNrE1CBlCJorFvRun/bFui9Om8OE+5q5AQxUlMNhN3
UXd8YpEGUiCOhIGbj9MVcMZ/NKYeVWv2ys8dfak2yLlBW+XTAZHCZTgFGd94c09EQFyFZOkh50Dl
hUC5sDd7/lx/fDtNqRKBTOE5w1swwMsO1rriZTCaTZf6NXlXzCRFTOK9h+CQdFAOEHkNEWQVQ+VY
eLvoivEl2Wo+MUulbCAT2wQvrJCsLqI2mgXAHe5Bckobztq7wYYacXsptCeftt5+LIAPjXeNOETg
S8QpxOwpVnSB6ZFoiXYsBAqxz4N/5QYHHGGyr7pJZ5uuxiVfYs2go7svEp0Y3h0LgabMWltE7ZQw
xUwOf7PExxazLOsio+SWEbNuw9FJd9uqucHW5iY5V8LCh4/0GAuwGSVQu9IhBy4q3Dq8IiwhOZIY
+Z7N7CWtbJM1mec0fj4sRYCpRMzFWf0G0AtHCRm4d0MEga66dLcIcbWMFDI/1mZG3B6a+5B4Th+t
NZo+NDlqXYoet55cDmyy1+9GRVFSd1b5kPmOoTo6nhGAJwbrK1LPYYhpAaZc4LSs47eeBHmuEJ+Q
jnQg7YEoXhHVz3vh9Cp9IKNCLFLl3/015c7XeEw4k2GJB+jqwULlJ5YXs2d/OwDYaDgjEqdRgsT+
Uir63tR5MZEE6ppJmSf3GpziYrC7tuJtnqm89ixQXQu0j8to95P0POGUWUGMUf5t382FNwxNAlIU
8L33dG6XRc36AkMMeDVio3yJRibm8vZ83K25bEK05zXD9KrGouHedKYw84JvVc6wFcxd/FkVviF/
2Hs8WjGaMuzjVSsOfgF6g3ISNiq3gVa8Fit9RhjwOObfpKwUtsk/w2w4YCeQn45G17xLsROVskfy
CxB79mzf43MPaaeskQDmBRWQkitxzKr+Dcizq7f3PJk3b+LbaKvc76Iy+Zy0zQNnTpb8X5QWwdgU
j5m8x7iW7eKNO2tbfhGBKYmxF71y08HVkynWhQuXZtEMuCT9BPXplbo0LyJNqpcLop+bGTDxWO4t
F7vwymzRwnLgYHez0KlMSooPTPG89QtjA2fDumJ6XdI/JGlo1/kEH8tt0MXwSBFkEIXRNAtt92eI
xpOXUcNwt5ygSUydSiE+RzhCN0eVERnZ8Nm4Kfw1mXr5B/+Ht0WX3gcWQvjqJJ7eL3UBGauXR907
fRkv1fQTqrtVIg8khud+jTpeLQHBUAEj+coObbO4IqgWd9ZglpoxlFjYjC7dfrPFxuoGHwm3rq3x
fnOVmcZYEfFiEw3XHp8vX095mJ0tJBDrMaS9VUCRodLLXVWV0lBD+VYYyOeFkvHk8b/yhLH+EASS
+9osb8TEaKTAZVLzIPGV1S+N1QiHJXa7Cv/Gtl3w5vH1Di0MFmeSSr9uu+woegopU8eRZ5AKvHvM
GbSkijZpwlcJ0i3zrJCBsgJZKuJT3ATVfig3VL7seC4wax9CNFI5tbu4e9U3xjD2TTZmgE9C4fDg
/qyGq5VG+X0z4wqChjGED/SRB0wLUBNdX/3fqWG2+Czez5b/sxAC1NJXVN7H/ByNPc4hmaDopyZm
qaA4tMKSdVrU8BX5LtcgtoMo/8MF2L8qd4k1ktEPvASUIy9gZTs6oNrYyTby1hMZnhzgSa4hWHNd
CzqlJXy2pneHzbLEIvqXxBcE18cBPG2yJoBVWpy/Z3LUBHm+i8nLFfmGbO/iVvbKvOoSEQfUR1t/
BedznnFEo4P3K+/aAIqRQLE05Rdds463QGd4Ow0JQV/cva+GPMGVzPfTvhCqDkCWd1BFo52UYCk1
qGVhluvsB3wY1g45mEaunO8EkJ8rVKAN9yDtApxeVi5cnd+YJP7r3b7H9fBDFQA4BosMpqrD2CY3
H12LMGIP+1jw6vjN8Pa1hUEUEOeCu4dkXWhm0moxQp5Gq3s8JaMDTAlwAIctvcyByZ1vDjszjVMy
OeWFWx5B4Tz7xG/jlG2O0mCM0wyyvKijV8vjX4MK8pWKZPrjwZxycrVGYKknvk6PP4VloNpOfmiN
g2lIXKNoW3CzynOiS5Ua/oteMO44iHeA1NH6jR4F4xKbmulUs/DJUEojwXXdREUiwnhwtkuta5Lt
rFCDQsmprfSy/tkLngkEmBfzm2MD0lMtbJcaDCI1ze0R0y+iBSiXTNHoXZTHzb91GW0L002ULAGa
MxKxb6Eb6U2yhQUbpDwh/v+DWhLzN3To8xLP443mnsFa3P77HHmVgH6rADLtJep92izgkJRde7ID
LvOggE3wvOVqLZa3iXh6eK96W8BsJ9W5dVQ1Xag/iV2lzm6djvCdwVRsZLjRyttYzHo5cyC6L30k
JbVqOZ3xMEzcaMy240IJsI7uAX6E/dEs2WJ1TSJWhezUnuNUpmaj/ntpzSZoI5fSi6g3uYgQB2lL
Zmt9kXv7WE3YhWzfMxHXunnhBxHja1MsXEwmWoktwXafw0Q0RNulYYgcRKUELW/4h79745pTvAZu
KvBRvkvEBdbH3AGIib08434RNFzhJ/Vksi6E5S84/OrtA/ZlN7QPgqR6yEpUKJMGb34CnQljWuck
7hvnuWsMOQ3Mr9ImvN445heZJzS1QM6uuweV70QQ44yALou+ca31BISxOVTCRv3u50X47+oNzjyh
/D9nwl7BfUPXXEYj+wSgUu9BSBLNmElXFiwNPehcEdhCRmrWdJnl09g9vTLSrRuWBa0rlJ4mVojn
fX+aU2f/qOW0pLYUU4SlZ5n62QFcG3SjTuUSRk0FloW+ZH5hLySFtEqhmYA+YEu4soiSBTG6CF4M
BgIOBNp3k1l1fVFUcxklBpNHHHKQXmISEGFAIszWeANUABp4fQPg2aqp9JJ6w4NJCgTmKm8LMOyL
3t3/WwKCD7CmbPlPmOj0JOOp8whHReLRcdd+E9WEDH8Th1G5YOnLeMWo+ktkN87qwPQ6d02joHDQ
B+6RtDS7kzUzAicBimOOXboqAfJjqljgEZ6GmjqS/RLBXPHW1JP/PCGSA/47XTpnuNZ4hRJzlFxd
2dzt6qoelC4DZFpn9W1jbF22vSpcgICW2Rep4aAQHV0DfaLzH5MZ6RWXzCyDQMGwmDjNtZokA+aL
f+GoolGTrW+6d9NbjVjw4/m2rarOZgwUc78kKsq5urtZBgZECwEzmnwE9r5o3eEvdaMWnmDH9b6x
bMa8Tr8WMw7iib+aZmfg49bOjxxHJRy/jwRl16+5M6Wqsq4iRfUUN8oLbAgwwhm2oBuh2GIDw8+q
rbNeFKZ/K/fD0rL7y9lsn1yOOYEjuH4jne79GUZMZZkP5FbcdRun7AENWYjuPnM4CAzZeA+xfQ7o
PLz9tZBB2iR5MAW+BE+JDbpgViQXxeCiN1mGSxiQzPOxC9SUOW5n1+GQ9e2JfUx3BZcUdD7NDKXa
lPB69g9GakGMrJG458rS8sJ3m8aFsvFHUbgxHW3jrfVa2SCJJrlEsd3P7yHKPP5Y4anuGfSMsXrh
jYm28wFl4gNnyIWrZmSJgp6wiY3fCHOs2yfbqsIz3FeHUyFCpYBWlwZOySe5CgYLz43uDdNBH3Rn
sByT6ZejRWuVZRRwx+9Ks+k+LgM0GzBIEpn9DHHI3jgrQ3GAKHQ6BKb356xZIgDSL/SdqRRDPZ+n
K4OfdShIpaISmiJH507lmR/QFVMojvSc6u5MrZ8JSzDo6pH3cGtNAxWr+JL4lVDgW359NFPto1LX
XkQsbs4Y74HhMrRYBYK9C+FLZ6Bd2Le8tfCYWR57mYpZ+k72MOEM59q5bmfhBdlUKVxKCMUJh63D
K9hwAQB+HejaD2A7HpCwhtGM5sMhNiBQTy3fQz568uBzisI6iexaAcxKkT6sYIcBKPKhsubVcqNo
gUW8hEuVJMfFeO7SvJy+ROJ00sin+Zr0bxoTicNNvXr/FSxaiTTsT8d8bp4EhzqyUJKosb32/SUr
2rneDe366u1R+0SRV/9XGvWeiSwwSZYt2RuQcGGVc6dtu5L1E37qAg6O4bFr/fKrLVpYXAiYSLPz
vVRcbk/4qo6ywg63JLUvpxRTlojcw9N71wEfqrsu7Gyuf+65YP4p5qAYWw7nKasBXrzx+4aQYv/X
eKQN8r1gy2+NcBmoJd+0FEknx9Z9jmYtTqNjfxFrRbTjDxBTxmIegltYFxv08lharwGr+gFhAMT2
JI/uUhaR3z1Gqo4X+LWQ+ZgbuPkRq9TBhN8kRuUiBGTNWOmfEqCFQVhVFVvT0+X/T3B61HN+/TuM
T+LBmtlBoIv0mXcXxPmhUWgf5qxITu8tb0lkjfqAk2aqHn51HaWVhh0J1GJldJlnRfjjz6ewVnkS
Nn76SUGTQWYkS9rX3RR13cWYq4K7bdsUss7g9D0BIsWJbHAbqNv54lhpzMmuiCblwDQax4hzxnTh
viDkRYTn2IT/37OtqY0SOECGILnGtwdVjLxgdS8LZAES8ndW/6Yh9y5jqLiqdDAP3gJJhz1An8IN
JUXuPfN42/r1xKz+jkzTJUg+1S3RX1Do82iOd9RQKREHEpJBK0fRa31lq/6PiBfJrG1Q3G2ZN2S2
9zaYwhMhHGNlfV6d9xyAQ3CWeitAzNlJ4rX32w+jfHPes464WiJVUbPc6M1YK7Cqn3uMLazYPlLI
YE4/32rhle7KMFYwX3BOP0/RrTzKFYL2wBao0oQpy9MZkcrmntpIVXS1YleMJjVbqfchztAhrGmM
YTlLHyBUaZdck+bQoMCKzGI8R+KDZOiyO9dgdvO6IoHMAgMM2Lx1Qc4qtVr2P5se9vy9NpRJZLAj
tOBlEP71i5q34cMpc54xqVEbGFsNzeCcjn4ZvBF6Tc/nNvdRs5kfK0ySbXteys55TQpHtypgZVAa
QHvn+0xKo5SopRFb9y42AEJK8S4a6xGifwX6MsjgpCGi5BzwCfSVpKhjYdR1WjQ/jB0nzxYk88OB
Sghk+raO7s2MBVC6r0lk99onk992akfE2YFdh1ycDaaMK6qbDWbAnKkfVMXDmIWoWJF8WjAgh7pQ
NhsRgqgSz20l6l6O45+tVIduvbko1CbCZMu14W+laCW+mog22RGWzgiPlaUtZ4onFtcOdAjcWt0X
OVu4BGYzd3yhBHmI3yd9PbM2iiwXKNmklGMLH+Akf4IxyhZaaDGqAEYRTnYx9lqnheS2UpR0kwe+
JepGrGAQ1oawfbe9aadwHKLHwnC7GKCC/hp7BGMKf5t0nOEssJFyCWkIP+6VgQgHEg76UxCCMhrp
V7l9/bOc2uthK7DxPESylu5p9ClmEvheU+c0f+Ess0xA45ijvJ8oPgwVk2DPI86FOxzq/xdRZgp2
QmNqE0HN/WKzh7pu2nbdEc0Hgq9Rhbk639WZMyLoRevjPxkh6bscy+SngAUZYNtXHEdJ02MNbSNv
1mqtfKsALnVJZJnm4/3n3bt24UeKCjqLmDWqnC3lcchhliWhWUjprHDC5FLbcpdlrqSmhescijjx
Y8dLPe2QBct5sUuzuqyO2v2IxpNe7L/LN4vZFsEoCyjM3aDgvxuecf9HCVQNsAul5TNZtGd6XsaL
5xic9VcjOeDTYDsRLBfsAvfdx+reqqtj1QPQCRwjIVN7vSGZbZOopk1sG4yFAsGzqMfeyzGq4He4
1H7tV9O47BIDvRDVGaEDi7xpAQLdmYqrZF6FP6ZZ5x0kCDBJbHt/iHe+mvS2Ea/lBl6c8W/jgfm8
ZxGaPzvLrAnr2MM2HD6hztdw0/2WxR7EnLcIk+H86NPc/gFNmUnfubhjWreXxo35tXu8AQ5Js4wY
1Eu7pIw928MN2h9HcIiJUf9U0tnLogPeWs6F9ldJ2QekhcG1a2+nuUVe5XiCgcVOEB+3ZV43erIz
qsiYmCZxlIQ9MJrE0zInU5p18ycBianM1/lz794sQXub0y2ZMeMUxanJQqrYJcgtP1YiL/ZB1z2/
to+PT5xM3rB3Z3wxM+UoEzY170Zm42ylJlVxsGkjWo1lbs0sHHk7xct71fvI59iRaEX0sL2N7mNN
1ONKHoFqh4bOVpy/nk8OgsQmXBT3npZk/Psn+DgvFK0cs6DTGpom1mQ7KXyJXzOb4kj8T44PC3Ug
CVcVUDlNuAxRXNntbA2QKxUJnF2i+vNcdxW6qRotk1yZ9VAGYQauS62luumCM0FausFqlUg+IHsF
+AMEaHQi98Chde26OPBw7rrcHSjtJFY4AtI6uGMQIVDre5jjUvwPd8It7jtRHrxBB+E+yqwUQAQD
dUaa6BBb4mcVxithR+wNa/tj+b7K+zJGvhNQcQtgLC5CLbO0ELqo1g9pUMmJu0UpUNkE3tz982rX
4mMO0aB7UBPfWtQJG9HVqRQiMqj28h64LPf0O1AwUIyVBnyYCpFke3kPV0X8R5ic6T5uSo0UT70T
1cctIsMQI8xQjKwirpMnDwSkGWOvTm206J/Dn82jbtZdZEnMKh2wz9LploBwEf4yrYULg5gqGS5a
+Smfx695msPJDTNJ7qMBXh85MnBrGYKqTPHczAdS4WuCEnLORBLFyfPzDD0NMciP7opzyE4OAopf
rGHA3kYcROiCsMbKtoatYdktGgUKpTYXErYmhYczP4KRPDv6gTptzPt8Jziqul1ZETNsxhO33XRd
LNoZJiWWIeCo1DYs1pqhZgfxx0Bvf3wXcdWE3Ol4Co6/5zhzDwIqjGNUKrtQ6xVkTM3CslWhJ+bW
vHCgS2hPoGwR/ZHTFz9AXCseRE4yY63wBdn+Zzshx+RI3m0ubZ6fDTM1Qd8oh7yeCHf3s+acWyZe
bhRt5KnqvQLOP0Bqb2lhJJV4/0j0E720HhPu9Lwj6+x1oLO0OtUJhs6CLSpnLVIU8TnIb923yDAq
vFi4TvLOHs2S+muhBKCcPKRFGYj76CPk7j2LO6fJroM4EXa7YnRO6shH+oSfpIwi/rq2z5DiQbsI
OfWjYcAWcq7RfREWrOcmJ1MBB+OqdxZNC74nbSH8GuL1JB6ViyGwGKvLWBxTA6yRZAAojW97K+X0
X8ILekmm7kDr3R+Sm9kJuFMY8P0nzz4IvElygRy34EPJtB1qbjAtvughGL+BGmk0/qkxf/hzr55K
FBljhDZkFAewMENzJAx8vvlPzdabVKV5lqv4boN6k8DkvrGohdDsIKVlimTGgc7Hw2vp74fGF2qh
z/x7HJnoJO04/GEhG6qacWIfs8LyenRRfzcIOZ5z0T+ngHj7tGCP9AMJNDDBtCkMXsB08IRljCcA
CjHEWfq95025B7dk0wQXlwDCJM89cQCprC5O6VY0JdtGzCi4JOwqN5FBjTDusxeL9qcK1shQ6ztN
AsbXW2pBVDW2A3NY5edoebEyWdxxEy0/J12SW62YxD4NLWN7GI7sSK2R/UkSjZ0Czq8gFKlTtf0t
Dh6XEPpKAx8z9EBKJ8kR7KmKUFvhR/2TtWE975a9ngy9OiCNmJWZXYg7crL+7Ucab/wRcKXa75YI
9pGTNmlnqoxES8XAjQ70qIFWrVETKdPjB9kexZSecZy2bPN060KiHSKzQbHOAJGKVDN/vyBcRu6l
riGhpdRD2ODqj5rfVXPDOTSoQZsAbmE+S8ghJ7cS2uTCMxb7tl/j0mFQvYT/4EkxLKN6/63+8WIA
hqP8MYaL/DFxR/CUIZWSe6+Rd44PIPtkhi9Q08dVVbfcFx0hT62Q14nZgFdnoNd0AZOVIL7WrZ+5
HELmDdW1VwMbt2441wX0xGBWILdMdkNy3w9S3mlhCFv5fo+ipYXGucMUoM2fDBDIPTqrjCnOslZW
ewiLKFTT/wtfurDOc8uDbhnVKtdfLDJZ82iYS9lcH2x0vY65wQOYk/229R+pyawoIZLB+R10tc+t
xiWZ14WnNW5YqHP/jellx1uQp0d4Exc74DzBir0QFihCOYo7f96UZl1P0xhw3xZNrvWoFXRlAYg4
G5TcQBNU0kyCrvtaoozDbPc+whZ5aFEsGaYQ6IvXtlvAwWdUFM8rM7n5M07qGOFfITDLDxncVu2j
fwIpkQjgVUl4aMcTClrcAyn0y5FmYT7i0Iz4KqWnQ8PVPxKiUPOESlqNDp04zZFH3Oo6fwBtmdDI
z075IsXMgyaZcjztCIww/nLpLTsYTlHUrTTdzUUC97eri0pgPo2KQPwyLeXgU35/XDhXOQzNSz2C
HjDczJ92MDJMDH7nMfntxi/tJh7+H5R7aNIJbJ0Aivn7goiw6mBlw0djuCut+T5xYZdfdio+cGAL
kDByp2Kbwz6uaNUN/+IRA5yGXK16u1WQaXAjsoOoWT7GTR7ONFyPw+SWsEhU//AxXkHokbm07V0u
o7VQbqDSqAhqZdbAePzlZa40HxpYCuPraW3JgInU3LYN/uwcCIriJ/0wLsKXU/ia0ec4ZvHoHMQW
Ntz+XFNUMUnsd4TbTL35Q+DYLfy15o4o+NDVCAy07qdxEczTWQTcJksvdZnvTUPTlOv77m3+6l3X
YElt4Fv0V0siBKvI7lyUM8uUdwKB7FjwBQ1gKZOydCPoW4ZQeoQVaFCFJVPUIfUNlJlPQeTDDg8V
kEKYb4xEYNUkHQji5XmBnYUYizwSFHcBdX3v29nYu3ZCoE7rfcbRrFeLfkLOODZb6DEXbUg/tg1v
doMyfQEzOGDjIutLm09cyDrZLPTEfDtJbt3AvJTPY8KsY2W/GE1TgoUEp/yelFjUE/JWsctAdrEU
UzXNgSwafnlDWZwqCATFTUoZ1FryFkqMDY8VOSGDxbnHjEVDRl2PO3RRaS+s744rGYnEuD5DIQJH
iz9KpMh+Fh+uHL8xXiC/QDdmNTZhvOdmK7f0gpV5NxsE87UHDi3k+oC/YL808rvq+zxKaw0SJ5v3
ZbZxDdhputZubiIKkoiBJ25U4+c40imbNa39TzzBw3R+tUP6ELBPIEWGmnABwC5Y7Ni6hLLTJ5Vy
jugmHR4UCJwcd8JDz4c7ZzoIl9fc+DxYWv/ISHzATogf511g6JzThImYSvXM8izK9ewMPs7LDeq+
uaVO21IRGatbTjqCODNFcCPFjY0ecf1hN0loQ4sQdYy58TvJ6QJhMsVmwDTFWNNxDWdYlT01qbZu
uFtpCQAftVhSsQhibYN7r4v2Qh7mW45eFkPj0vL0df+PEGUWD+DIYWD1n8rgdEAqaPrkXduTdrDH
gTGnCSwjK9IKV+bdolMAjJVcqN0UHrktdAMMOya/SS/CDh+mCeP1DBO/irsub7j481tV38TjUHBu
b6Ab+IUHToGv2xarLijEoxSjMqU77gqMLRCyuh8Awn8bpTHv4HWMI/oYrih8PGeX0sB87CB2ruQ7
dtEkF4pSsWfMcS8FjfeRhq0FDAn3F5ugGlvPTNlLWw6fQibekpKCEK3KMqJpFK6JAhYEY3SBCOd/
u1xBJtbulcCIWkrkle/Ui80kXCOAJ/OPbnYEieYYSVpBe5B1L0BWreOXpx71W1RqktEHy63Pszw/
AJmLRLyjyovwO2Ht3OJEbynAu7oisw9SLQ7/l8LDkszhMr2BWB75ZaGgud7yOqj4i9a9+ijwu/AL
O1ie4wll1tHnFcmPfSSJ1hO1pOzR0Ss0nBAVxQEDtdhpGnSnLuyiozSrxUErZQ5lBeRHWiKcNpvc
R+hRbUJz0yupsLHAzUWXGihX7afFWDoEBuMP8RuKUd85hOcVkmwhTl4MZh4k+beCmuwAZV4Y3Een
vcV1NJFxMPceK5tR5ryjqpaG5rrblMuiUhXPrculZOgxYxhSYu7uKcwXqr/EAjBDQJkd/y9LbRLY
8pPWD0LGIAPH7T8MbgmXUPPEtyvCMRZr3IR90V/j3dDZUvPP+CaNmuJOaZs/GwfDbYMmw9gAl2lS
C3Lwh9PW+wYuz6aSE32fJ4qGSlr85pABWuayVZjAZ8+h0CSDH8Wk7d89H8wVAgFQ1e41N5kmUZnU
H4NuzAznjOtYN9qmgt9ZeIMwCQIK2NS65DemKvUtJbscladCNg+nKpDF491SjsDww18uyNjVL2xt
eZh68e8Dv8+DQB+YTHSUk28Z281JMuI989YEHy5zL2fshUaFwQVWtp0fPoTGaV17WdRWwGUIFF89
aBlzbWhIMLtjXK4DKFu5e4ON2EmEUy93t4J0gnWwpSGdbJ4ycAabLyJBQMv9hVd1qGqAvSfUwO6b
g9uPzP0LovY3X0jTrzNc7futtMJlfke6lgAgL1ZpvgODkZZ+pN9ZYRdu95+QaX/n50W7MUdN93fk
QiTvY7HA7mjd5YBvdF3HELB4hXtikodjfzbQdT6o27xntZIzXicrh8uAtNa4fEPq5vryjRiMHXac
diEu7uQQjXOpuaboxwmm/ydECQNMMu8Dy6979tDyBTaImloLpcYJg85IwLF1tXYi66F2j/0b88Tr
octEmt2BA5EHwKUzIH+9oKC9QTHQXebqtYjJEyEQ5gyaQ0cp22TeTbMwBXsU9RKf9iHFBX1szHWZ
USqMUHpbBF15bdor6bA1Q2/LOoybyxFNSwlqDtrD6J08ZDpctSoiFZFNhCOVmtb9IIuFSKjobP7Z
NRy/Ro0r8qSsW5UcmClr9QVZtXBJz4VPDgDtyVy8xLwyZctS8NdWcyWlHQm/P0boPifAoQN7EU3D
0sbut6Cr8hU4yawPYOMEqBbJgynvaCp/qFoLjnWPfgLaYYXwkya4aJOB09hzfCDbvhieeP8qBwOK
Gw8WJtr1UKv2VRWPFDe0uumm+Nb5rmAwePgjjwWa/GOt201jUvO1IpYZ3onnIUTD//av4uaxPA1N
FCOyIOQhClsfShIIHDZtftbm+MRyAj1zv66ggftIrA5SXsgS39YXP07lCtjspIZ7G79HpHvTjM+D
z4IpQWrZT8DG9r4DfIoIdFIolWpHx9MT/D15tgYl86WhcBpay0jo4iVXSRzEScT67YvDo2Qv6/3k
XZCYKNipNN9Lvj5XhVWoC6WWqrx62i6G+FJtmwQOhPm2y08GGT73BOmnzDqvxmn286K6gkWHu4hB
arWQsi9JF44AHSQzAAy+4QvxD428scU6eUnNmKJ6UDEXZNHDUE7dwFGDHo6ooI/V1meItyKe1/Hm
IbfAJY4+kesAVfJBoAiqRGTvXR5PNqhxtiBLfY/HWHWBaca8RE2fRZ0Lk8v5I68EKWVqFnv9GnNl
v+2htl4XhVc1D/pp/8LrN9285KqybD9JzhAuPV40UV9hMF5asfJ2D9SOKqipPsctgAvBsbr7zXy5
dlbRCaPMGZfgzcqKId3eiQYlG8+3KPYYW5l2JtCSffnWDDdzbzZNzQC+DZpng5Z9mSEab0IPI73D
2kqTIcuLzK59bIV/Czzrqdry+yZGxrI6s+Gimq4VFds+37nCt9zPCrYGwOca51QI668cpBDLDioM
Wdc+zAET35qgyYPU3I1TAfcX+c4Iik633ZDiLGCCMUG5ICDL9QlVtv6t4+VdlwZzhu5G8dNP1Wng
eSVtlTUo8Nlp3VkyCtwdC86AehommqT+qx+api8TkrbOEBimy7ADU/RukQKqBVpDCB/tIHI54lXv
nEJXYqpbY6NdKDkd9CEOCFPyHyjnJIryQ+ZMPjxESHF8lWFKTEwdRGK02CC7CMuueiYxlQ9u810s
5CQ4R2uZCn9PMkh1Uszt7wqj+ypAVkfNeFc3EP4/rIWxq9JpmGUaHldTCupTxCeE1ubcVrJwQV/1
LUVrUS5gBkGXDjpMSfIhxvA+YVdBWdr7k0Ghmp0oSvIOpwGsIeW33FkCp8ziCKRey9CFRCkVmM77
jV62LwZ0QiVQd51wzY+omxuv0C7vnEJXIolZdyQ3bNqtmnz5zFRfWd3ZTXgREBIFsWQVDk1yXlOX
vI7n6JLYuasSE3+R4N3Ob2Wn2tSPva4koBsl2tTeY1eOU3dfLCPaBPwmwvdIeHa1izMq6B9g3m6A
14yfqYFjzJHWDhMcH8FjEYjiF7ytH6yqNWNZUFoUALlMLpCzlNw9jPVuVJpwpgGWDqwh5e9CGtwV
9ebQL55lpBzTRHJriXEIn6xdunWrUDaee602Darw6mxfZSy1T+6empjQM0KLnKvMwp8ZtC7Yh+pi
f0xolhC0izNW7U4KyP5dBUarLeodrWV4EeyG3VeaPCwqdqXOraokyUXxE230cnDaEkBVY/gsOxHG
2gJJHKEZbTQjnhHQuAAdjcaxWuzqR86Z9vA2WMr5pX/Q3G7IO1swNJfmZQx7GSrTucy/FQCIfuty
4DjTZWoQF5p9nA5Qf/evygFIpGl7CnskGfDZmlt52uul5gKNHE7H85lNGV3Nl2aHf2SGt4EaXPNg
hHJMNllwI4IKdXMOrbupQmh87DTwfJWGZpNRd7Wh9PKx7t3LP8xnQp6zt6H5l6LJeJjI2ajgzq+J
JmcDmetglvjsmebePwGldt9pIG7kKbjk95ycW2aITsOt5pYCu8W1vZjuaFSkF77grlsAykIzpWfk
lQ671tonTog3JvL/QUf+bFwAdbjBq+QyTOUJtU4TkL3TJWlniHfCMgxh1Tsde2Zp/zEkuJeqElWZ
Q0uwUQcR7yhaaoKFQXYR3r9MFAsM1eVgKyyIRxmDHzPxrLhDMbFmN0aqHnHDWHtn5bI+4Lmb+mqM
wofD/if44EM9oe8PqGt9Y6yKJNIG1X4au6AVtapQEVDY6WzPLu5QwGrELZ7q1f7fIrj4km4SOHse
8o/AOex2T5J1+cQbboOoE4yZeLZrKLNpEHiKXj/cA6fKsL9iO8PK2CghT/pif4O7vfhQHpM8KPVb
sy2aDtAnfZdjJwK164Je6h6+3XJ91dC9NWoS1oaH7OB8k+C9BD+J3KTYTaH3WTKUssDJ1cnXYFvm
AeKUDivD6mG/M9l/FvU8kuSp43K7UFMTAbZeLCSxTc9cwu4GocfHyunLOYmWeKOLXfNHnDWEP1Rd
L0ITRr5iqrye2xXaGckS7ah4cKPAZUlh8M1wzmS0ByxAd23FrLCJ6816WzrjMZ2OQNvNXJmHgRND
rK/D2GFfhSR8StbfLz3/ttY7arvmCdF4XZRPjiT9zp0ydoRfQ7Evg7QU1W0bjonMVJrSJKkqpQ9k
uooq0UXKG3B4D5+2cKI+RATvhYZmuviH6caLijo4SpoRz0e8GVXcHluSxPd/t9gSTpPmmtlHPSgY
beVW8+U83719P8anLBbIu9vyFDaWMxq0ZTkEap9Vmq+mzQBrsJ3EKcoaMk7PxUwyvoIxsQ66nXT2
q3DVT2Cv4xQXFMSOEmOc8RPwAnm08dzwsnAWV5vop76562i0XsVUS+xBxrURMASt6315QmWr+TzC
p6WoD3U7dpH/fDbxrfZaul5agiQ6+mjStGnyDlrMjW31yWA2zJPyYeWMRW3WeItdPCCrsEwISyOv
WGSlZv2ZnOLnBSNFbxMqpLr33NBK9xRS2pVdk4qEVv/L1iU/Iq8fI2u5RcFus45c6SsIi4EaTpJa
XwwtBXuNcCMmWQ2y6fDUHl+ye+K4smIs0KT/UVKGJwDaN08bGQqaXVP9ZoSv01mqUKEF3g9OQbLz
zM4M1W63qRJsnUOEDX0Erh/Kc9I3MAR7zh7wO5qC129tiEV2YKietfM9IDDkj6BESwFnY4YN0sfK
mqsYYbi7l9A1E64fYB+YcxSz/YXjKjG3VbmG+C/YrdhQNAvV52kZGQZJFMiY+UZL1CsEIAGFRRty
r1qw5Gv5b6m7Av9FhRqIeNe+63TBhk2GffVgE7TFFbFChY8KZ9Nfqbhx79GwEF/IhSS/VNH2+qsv
zMRXCZH2tKQM8z6ZwEYUSwHdn8jFG/S5OGZ1RSoEiOrrLIplE2+3EiW+viDPCjWZz5bPbkJkFNQb
QfXNikxVBeNNaHuq21Q9tdJAGMM0x07iBRHAI/nQRmS2BCyOsp9ozE4JT9/5kFTXwysHbV6f0NaM
B/ReQ7ZNHWKP1/MKTogzNCFXFqSbJTl+/KKwwBN1CX4gmTcgRNK+LkdAM/+H5PfnF3PwRE43IArg
tbKMsuLIfxA7NpFG+hLwwxgBMHQgFS4iOUwvZ8m/rOm/smACAAysVYtAHUFDvyAkr6hNOMcALvL9
09Yz/J9GWpEFwQO99OA5mCjPF2mSfuVwIZrAfN7B3Zk4qOHMnbZuPM6CnGEmT4GvTnljKIIaFxcK
qMqZF/xUHEc2yU1CZVnR3ghuAiwsQV45QDWm6Z72oUOu4bMGBC8Phmgh/kFNTG0FsdVABFC5xcLE
fX6oU3GK6qLGELqQ6xa0tQiPROpCTOCm6bBrvGztRPCslL5SOBLV1KGiCHqWEj3rHqYf8ScGfg1F
rWX80MHPPR9owuR2bLxHPPuOXi614CLD+OOXuutIhC4vXkYUvsI0n8t/kRHboFRUj1amsCNS6iIr
x/hWvTKqyjT+orYjZoGKG80mlGVq+v21M660lbBmHZGgPhpfVu7v2YUYiK27lZ/duD4E9tghfyaR
Fhu3/1isRGikLEEL6an2gIUCchN++AYfzmlSF2whbwAqLugLzCLDqH4zn3iUSalMnA+/lMbTZbAF
tIdJ/PUQra6kohWr0KHGUONEM4AQNXs+//yK7LGMIRQQiTqKJBBGEV6n1mQpmp1uDgOdQyH4cU8u
xgjHO4Jhxl1xJDkbHePcWG4ZwXxC8OhO4J6TUakEdtmad3EcASJRkv+C8sNCMYh8mplFiP4PTtM6
2HCaYm608rXVq5ujlu10YUGSSHz4k7OHCS+XuUAFRs2Uxc1r1FXDh8q7d7syWIHIlpsBRH0xVQc4
rBG7eHrXmlsZ+ZMPYptoRpIWeVuNNqlWHT/kFHUpqyY34kWOCcHBcB3zCwmnlbr55DuOwN4B5c/u
SW1l3Gohy7yDXSSgrdaIsRmWUM0nVJkEQH8guNS4nQMF5PR6eEXJGE5kUJH+RCWZV00nvb/B0PKZ
TPmaXxuwaYop/j9cUo7e+fEFrB8zFk7+FsUJF8ItNPHRwbRfUZXu5PyO1TimP0Vqc7Y+89JWylHE
hJzSMUGNfAL8lw2SDIQjYKCGEO6UuShFBxLU1Tf4mrmd5n526lkz6/eLp3ZDxELz+/xhdRfLDAah
ELkXnMKSBcPRVni+gsR4G8Kx9Wk/FtFM34ujeOFQckrCPGwTMfFSAj/ePqtSqR91BqGKPh+/NlZd
1ggRj+YTMVEjCdKN5vy89R8gvVQJ9k5kXPwuDZCkHZPjG8KoQBL1UgtbYqIJM6dmzTtWbpVrmCWK
c2beg3ksBpVCpa+WdDuWx+7WIObG64+Im5wi7f2F8NO5ITTAKmM47uPdGIGNGQm8eTh0+s8/3Ubl
lFMyRMzS2VTRuiiLyfBqkX8PTRA2YccFecFDgSFyMQz00gxSciV7Jt69B946zY/zUi7N++Wo5h/e
92ZyheHt86p1rzK07jbFCTi6W2UxhqJWMt4NvfyzFzmIIWXKRnvAHkwMPpZN9wihDuQjeR746wOH
v5VxF7ozv7mFgCp/XfkUDue+JAfRmT2bbF4cgQb9SFeDhAzsyhk6pcvXB4ntOYgh7BXDfDj5bnna
rlstvNGHUrvHTWZsmLj+rJ5jv0Y9lIDexQ/dExYg71OJ8ySUuYNZKnkJxh2toGhcnujpjFx5hsxm
qOWTtbhOQqdh+PUdvUe2oUJXXwjMhJIfEO6GjLYztOVk1lo7BfCZgcScb62vP+at8lQmV1io0Ly4
UQUFM7G85KStIJz8Fu8dtsHzwk7K5aqWmWknNYX/1vMd1uZxNtTJogLKFr9tpy/2EdZp40W4zZyw
19y8JMY3LC28rnH4i6AyNpQxm1G8HInufVZEw5zwWyAdpPLW+OEXnq0S6Su7xcRR2mNhh6W4CM1h
HZzp82RMO1yvn5exI3kPx8CeiSHok4DYx+e7OR4LePE3KrxJGUTNiwJUfntQUO53VMjWOUFKtb7O
SJXNLRftyu4XhhLApSgIeEyOXkVkuyFtKilxa+FAETKh63IH7enJJdsoxGsanIs3Hsm0UFJajv/h
3GTRS9K3hxFtcLv5wzWsECw4/NQGKiWVlXkdop/K+T+vCBxiGKfoE66a9mEfDwgrV+uER7QMzUBG
LSCyI1uGfVFGG+3mGv9/8gQEGx1q4RXSCLmmg6V3SL4KYEAn5dKun2yFQe4zyFP/l6S/xQ4HQ7Gv
aKvLmQ+TwfTE6IwHWYbifejRTxBOjm5YOdYAs1V1ajJW/0mYW11f6J7TaBnZG8Jn7m+s7yQqOFDq
oDHV/QU3ieO0SbxD42yaBAmvrF+nxtxavX7YU0ZaMtikTvwRBuM+2BCg/MG4STcCX+DbUnKcimb/
oCVVy7I+dy6VlMROkz7YtZTlGk4AISk4J9rDP3kpOyOsVTMnBq/kGogj7R4TRcLgyHgi/tCi0gwL
Zd0hqEKt8AuuNW8ORKpVeKUqYQZh+iDg6PKySmQlYXlm0z6d+7jY4PaG5fW2V5za+4Yt8b8uvIGq
BkSUZ40OtWLCVVWsVlnG7oxSAYdNusve8ZbJt/NQGni9movWXfMOvhz5ZTxrznz7UqRC1e+49UF1
jBbkeOy4Df26JtHWYXJct9naeed87a0VfUdA1mmmVhwGTodoSgjs4WJBtkzPu3JWavq0rpsDviWC
jK73OY1U06zdkzRKScJ7l9WMTrPHKr2UgfUSKq2odI4Gh7XqYN3lwpUQegb2vsZIjTS8evzVQmMM
DUBvJrjlxlQB/rwNxMbU7fRpgCOXDYDbVJ1z5OZhSapLHBUNX5eao4iiL4LuBUcCvpmgTgVhQj6C
DLtTUBdKkLXlkGbTgrrzopCpyPTFRdBdNMxcp72Ty9GRyBAvFCmLWjdGrcr/QeVGOYRxnwGY/ont
EmioC/qCO/7eChCqr86oGNCL6K/Ul2SYJZVDewLk1DUYHbcf+/qgyWUmGoeoDa5BkAz34PzDMBWO
MprAyUaodjUtfeTqVCVb5T/mFCJitV1zQ1Gpj1MeH7a7MFVNDmb/WHBtGkEq+KOxx320m7DUq3s3
Qtd3MrKRv84QPClke7QTrcw9bKbe0efthf+Nvm+ASJ4FrNQtwpbrWOQ8Y8aK+FQwdN7zYc/A9pyE
LBcXdP3dOX0AZkG7Hf4FpuykIY2G/Nn+/yfwcw0R15X5ZxuBtOxsSo9pRUm7XK0y3voAngdaHfu6
7ZQJHs3eiXVUW06RgUv+UDTyweWlJIBuwEOLSFNREg9tjT6hfyfGmL8HGOeCQZDll9Uhipcii0Q9
y7U60mgTnHkVhgvp1VjLhkesplaKBP543DmGZYOlsu6M0ervW3EFTG5Oa+3I5qZ8MYUnmLB8soTh
uwbyrlTrErqzjtu5vxMsElR4UXhWsmPtjgrtS6KbnRXvUghDpaThBNFSh2fzT9ym1yhOgpw7XTEW
17G+s8qBD1gKP/EN0FaVBIQMtIJNKpblpk+i91VklqVi5BD6EKzWj2zqpjkcV1yWLYOfl9aui9g2
HNbYVtBHEBUEfZq86/PL1yna2L0hMLfrz1a1K3BiMJSeT41IrIvZnRKvKW54BcxCSwClLKI/Zzdb
fz5Sk3MldJQ1Nk/Vg0tp82JT7JrYhEyBKEfqGvulljNQMF4pgc7KoXMMD+9LzoVP3CCqjZ3eMFGN
aLTwNtiBhtpa22mL1I7Ljcsjs/k/9D2tJXSlOH0n1gYQrD4YldrL+tjxAgGX8j/VHw2VhsYGuR01
wPKbxoN4CkLDXEX8dXUVjLyrfLE5YAS+iZmPYc8oonsbw3sS7LCjX1W84qzMQdCVJqyJqDyXV5rT
OcA8RV9nIMSlpccDhiMf95Qlq4ef2XcRHM/dT6w5qa6e3VSVt4H27IEXq5Lp4lNk9HbHaP/rhFJH
l8Hceogsg/iPWKnE8WePj2XwzoR2na4nkZdOiM4j5UdoZX8YTxxAhopJ1f+r5qaOF2rXXRJOFtjc
7WmMlXCPyVTZCEZDC1bFdi4H3Uwow7Kn1mZxs9e88SyV1B/CvJKlA41ZE9VJspTA9xvNEBHqeXrE
6OBAMS0IqX9UkhODwkd+U10MbHZjGvTcVF9sTZzGG2RdeC6gEjdn1o9A8fS+7CSfvs5fh5vaALq4
hv95yqY+qnhVbAA6ZeG3IKqBKnJRd5tqckz6pPImHnlzYrze+4oAHngQsm+1hsE74BpPRIYYSIyi
BApHOwRm42igxuU8XtfCcWYOZxHPCrTNNeIDRIwyq6OyqVEBBdwOdZyG08i7NLxk7/IcwmgNwi+Q
6kT2ZqYJ5dtz3ltlYwdGXLTO4KzGyYTHqtUy4YVgp262xVzvXRSvhDsNPxo2Q24UYcmPt4ssgmRp
YnmlOKXi/3dPcWFyiXOBnJvsRdMBFBW61EeM24k+vr6gcEEHKFcGjdG9Z1gzprbXalF+XuTZyS69
kXnvAWqgGv09aet9qg4U8xQWAh3IyzaKwPH9ZDzZQJwtL1mK6eXrvAy7A+oomSulnpYvLh0i0yf9
2pPH6rdmzSlL/LYl46c8qw+rrs2ZUG0qKUZw+TmpPhPoC7wnI1TAZACyqi8TpJ1qwY4z5t4dxVPm
b3u6fTjePMSGsFN3/auqrL0EpgfoCjtfKUzvg2frOfqRZZZF6b4bjfkQm01i3MRiktzJYx2OGYNU
25GqnJBaZ9vgX+i2zTxQ+woDb8lkZ1qyQJk+mv6AmKq0oNyoSchnlig+k3uDbJMLYKAfNlqEJd5n
dzDEwNQ8KAlRRm0ci6wOZ8J+PGf6nlRGji7A/sy0bg7UveozubYpyDD0I4+xDgHdKzGzHtsRYI9c
0h7jM0tkyaBHonWMBIgRPr/zI5nkADvignOoNW3gVN1249Lstt0tAY8CpeIhuQXqjXQK2IJ4c0Ve
d+gD242ymZTO8kMv9vokq1KGeq9wIlkMQbRZJBSoqNAKyZ8CQkfl9ibXeUZm73tBHY2U3iBb0nQx
jNjMT1WsXtE+oWfaGQUubh+zFao7jh/aeR8GfR+3G7tnC+oY9vsp/SU95ArLnDKdkohWRFmxF4co
KVz4Zau69EOJ3DLpvPVBjhaOhhWJC1q5GQ1elE8Srd0JTJKtRjPb4f5u/3xGuklyN5+q+fwrL2A5
bE7kb0zWD3Bsayb5wohc+i2xaZ5NoMH9Uwie5Q5s6Q8CQHSKhgdKx66728AEcpppuFAbF3hTI2Sf
wboEuh5UZIDugRHyn4ejlbnPheQKTKxlJVHJ+nSGHvGUB5kZwios+3ddPcSeACFR+ZiduUex8snh
OCvqkiaQSQvzogyA5vVjdTK5hxMZELeQn83AeMnaSo0O3VMBDY/vglTHLlOPiHtDUkLp3+3hj+jz
RlklROKAXflOlbM07k411Q2aQc7RG7OJ8zUvs6wCee+qiXOXJCE6K4QWOw35acxlDrQcNaFNk+ax
KrwXt9pMAdpTVgM4K6XB6s+Hr6J41Ocuwa/sj6nG/d/SfizZ9mY+i2CWtCPtCeEqZ2qpm0UYOXX/
HMeFEZI1/IjXGYqDVqA//fN1AP6fjzKz0j2UNpvsvgHamdzlDs3TsUvOe7aeVDeI29KTYt2bLeOa
VoQDO14y9QHbcdAWJjMXgMtfYLcFeEekPuTII2kzNXwWEWFJpyFVleUGwNNnA6W5Al26MHqOuBuc
n26M2HFje11dIa2gHsSTWTCazFxXSJ3XOy81B65stqVEw563/PyODajytFQUk+R9F8qwKrzatMih
XDK5N9qwXyPQ9cnZhvMkApDuA6if9/dFwTFCdcJgf3bHXZ+y3I9YV2fCxeUiRieibu0JfFA3nOh1
waMju5xyE71nivknBL5WR3wA+3Ag2t9TgBLygyecYtHECiSsecuAbtTxxs+kKRSEQPODvHOHvHCY
laD/AyMEutrKgAzWMchS2A9gJHKFxX8GD1r0OKGa+WsrZzTCMDt4Z9yl2eMEBJbUAsm7+yJE7YE9
QO3rflHA4Y1ONj7X4w79GkaOlpisuc+XsFZ8sl5x8BFoTUwC9aniXS8pAtWoha/FhG8AJlBW1LjB
PIFp0RfD3E5IGcyT+ybQ6Ght11iPskvWjH2vSpXaI8P18i/UKsPwHhDWPCzyz1O/lmgvjkzUDPWb
L8+rIWSaBNHRmZJgqLFJ0nuNgOwrhhYQAqW/VXNsEyIpaEa1OfDL2kkEsYPpYl8IB8hAm9LrlWJF
t5c/gihksTG/I1Vo4NaO2qjOf5fX6i5nFnp5RWlwDakY2BUmae+y7ClOk/IKplCYsrfqldsmIWqz
ajqbnv5WZkHqD9xO/1vGf9ft0t2v8Gxe8kDZvaeIaVDKp51PU6Hv7qR7+wLDv+g/nf8X+U2Oguwj
Rxhj3rHjR3JK8uoYIr7//98te/QITrqvUKAdE+f9yy3h+WoCFiw8jQ/iWU54dKaXbIusz4a6Zx5Q
2rAZ7+G4CqDniS18qAaD8rIRuugYbo3Sa6yGImrGctzBKjXRMcyBGBIv2q2rNmAw2P4DSW08vQgP
aQIAAZixvWAJ/DVhlHQB1l9qXJiJF2nT0HWFmRRcS0B4VuIgQbDxqLYPs7mzaeOAdVHKoiTIvR47
sX1/+gFA2xQ4WyfuNIfEdNYGU8PreKwmKlHitKwZXgUR5NQGz5orysxyXsZblClbJ4SJLsot2Tv5
AReTZga2c0X5TKRLYYlYnJOfzg3EF3xuXtIqYKzrF3zCvft1qry2DFedEdlNePiHlX7rJ6cqx2U4
ciFGA34JhEgyo4cOWh6tdyFIxI/9HkXVHjhLPEnvanU/FKFm4GRAhelJAMsA39iHlxdi3KEuzQAk
YdCLB3LgNKrG/GSvDFAh+ExJzg+jbsOxsHLwnQaHP+01NdPUHOSJ0hZ0r9xzf4tyccvpVOrE+6qb
aNggaJOGcEWdqu8jcFyeU2XzjuZKjg70Lu0DYnQX3O5fysVbOOehN0JDVO/4uxSVLsQky09FB/Xa
JjZ5I1JX/rO31axxJFGW+K+NIkM4sMlI3+EJfXrLB2XKoagkc8QoJbeBLNFoi2cZHzHgn9lmOMoX
kTlwofSX7Zp00nnslVmMO1Z4dnUWw8ZS/LcWLzF7QdNwHuKkqeMDYz9qGPxsPP/XASUnzwpZOtUZ
19PMMcIz/YPWvY8TRUymSeu9QxthMbKCCf9rp3DkNqm3xloPVFt7FD9V1Ywfd5YY/ziXlAz5K9C/
YffmoLiHQS3pumNUGZREFAZTYVJy2FR1gtye4b8Gs2/RuE8q/kuaJkjw0+SZsRt6E+pubdp2kbmT
6LNfajuaSAjUJSWGVAKNsqs/B+P1T5MqybJCM5LeqmC5pNvJ1fIWKYnLk+0nozJGm5Qt0aRo3ssx
auKV2irtx/vZkmyrXABa4Bzk5X50UYAKusq3vbmfxee86kPROvdzqcPkThdwWzs5d6DBgdlYf0Kp
/YMJBkscpt5jMxUf94ooUaSjx2Uk2iIWv9hulSjA9mv6KfUIv9FMhW3xueLP19KiPiLTU+Sr/eOV
d/o/WTQYXJNdFs2wi8A9SQ6t3GwqV4KS86Mqajz2gMhzPxG7p6p7YIufgIYXg0kEdcR9FjMgrr7u
OjWe0lS9mfchHMddPZDmwF06zcoLIdwvEyWl35lphLy6IfpitxHoCnCgDsdTVhmUgaQ9XF7M/Xbb
ClApghhg3hcJEc45eqz27T/QZpWohTUFRFoFBltooSrue7vfRzsF+GsVnelSibBd0vBZZjfKqo7t
nk366btr90VuN8WivUg556ymUuxc1AK9bwbkuJY6SE9oNInA3owUmiZbjVpD5Ty9IfA28mmr+YkE
URjDryJ1pS5VYBPgoysbbdqxA1NkR9wvgadEqAtNMYtzYsW3UW6YsovHjC8IDAIvQ4+0c23dDefD
R/cfDozu/3dUmFchN2MDI/NlkFYnUBRwjW/1pp7pDvJzqVmpETKMT1mdJygLrBocdWTUmGSkHel1
IU2qn/GLZ97fO9Lpt0i1/A6DRJt9B/oBlzn3BSGVzBHcl0Qc2NixQ7j6uKJBPdAweUVu6j/dX8Do
IkiF7hxdnS6fFWeKYkybbpJ4fkxDOHmJDADPExmvaxp/YqqUyubBD+r7G6HNwpRyiPulSMAPbvC2
eJspCfBLaWGYA8SuX2bRY/qx673FkTfQff3nSOvMw7wf8uH5xLo6nd0Pl1ilLoY1wZTrpNMKutF0
MhT2vPhiIGQDm/WCl3R8vygfSTD5SaII5fXfkK5bq+I5cLhuNV14WkoKCoSMVSvKB+zRA90FzvF1
no7k6xV1lLlg0+7qjflDGmOnTRXVzWaGsv8+Vy7HpKPXtUS2O4ZJTSyLDg4gPTFE5b0SlnVjFAxJ
VxCHp9hX2UOLtF5kbGtx8iFYSy84kFcJa9EetJ1KTTX73SChys7kpjYIdJeTGI8yoxpZbiu9lPDw
aIvfp+NTEliuJj92ostXoR9A2RfIp8M9nqw0QJXdfA1YkFsDkYZtxhKaddCthbuV82/SO8ttBNX9
X/i1NhbHqhQZznq5Tsba5q/tDpFWq6UHsAbJ7aLdzGn8yh+T0AcaJCg2TSOPTmvSdPN+5EPf9evr
BD4PJjMxApSlmmf169Ogdd/s5qdL3TgoSQup3N0syPhTK4Fm8TsuuQ9QdRU3RhpZKI4tr+yWGwJX
lPFzMYOYcbTzeT0ALSf+FjdYdPNsFvw6X/sPirRIydTNLdXQk0vbSRgVioRT7GsEmm4jGkFA1GbX
yAPgnIlXCHjKNmNYwvOse1HkI36q1B2qHdcjnomDw76uknD/P4vG2xljPF8COC7gZnekcka9kfIu
pGJTTsKX+x5IHt44uZAjyW2CQ+z9lGST8mrNwJMw7RxHhpU7pbV0x/yKld8qn/1dYerknc3FyKdI
eQd3q8Y825E1ihYLaZPrt8gsAccVgGALrwNXdPe/gmJ+qyJj8FjzlK5+kXgRzAl62Q3ZkglVvhF7
O2qrCoJCT+btZQfDG5rkVjTZI/Fi7bdQUWa8YNdY7sBFwg4EAxN43MSGrfj/rd3AvAEede/xYfXr
TgvtC3iWsPj1CQyqnatjHFtlC7c/d/fkcynt/XXxaLNMx4BrimpIFhXhlGKr5UpOZpjetw9UytE7
mQGuogaiNUE+50n1pA7uZZIVA2g30Q82jIzx8AJ8atHoHLszj7NJQ7teIC9YiObl72sgTyGr6DWw
zCCkM2+bigdtZIQiR/JhU4Gs6pQNhYWLKHXx57UWdo4oP3AOfp2L9aPAiKvfChsQs+qbIuXAXI+W
LMcpZhZY9KR2OrV192h+Nwc7QoDI+8VR/lKQzp8lUpw9g3zjvjIar9ZoNqdujTKMQuJDwXhQ2Lbc
C6CPw0fkh4j32c8XKxEBZffrTla0oJLi/z9N3/6/gBfLMkSeF1pymVWbMcx98d/VxynVIaMO5JUw
wJbI9qh/HJQQSrm1QVjEepNwdryDnMbQ7zQXj6R3378oO0RW8mbCopRQF5AV/H7p/zJBevm1VrKK
ch0vCh4x1ZbIPW+Rrnjn4n130SNCwAmUtskLkM8dLFLwc+dvHOmuTSzBYql03qdYClJUnTNzlHzm
mjNTmzXFX4c5n/YXHCMQ9jhSb5JGUwCQV8OGiOP3cpUOrS/oOMbB8Xvj6xvoHfsIaK3ZL4d2vjQD
Xm+FYL1f2VBpcMKS18EmLrtS6RCgwOp5lDbUvK/bOpLxUiObHjvNmL6GdeiwPLVPnI3JV3xiN6az
BrFKtWTb2wFWB6rK8wpysoh802Ogko+t0vEy2KcVhjJTkBsglNkjxaOa7STvFuemcjc4SuRF8oWK
C5BU+1XTWU1yEn6kDP1SrmEpFl2AW8yqlYVLbgbgixueh0ujUG7Ar/Vq4DBSe/MyD5dBPRoFVkee
DKMAG2RyUvU/Csfmwi768UIxeH4eTZz8ONck4bATLCQNRH4R1IX3PfYDztIjBVgDnluwkQqQINvV
H0Ok9i1ZOPN+A0GqhsZRA6oFHUAad9AERc5+aXRUEbiQzc2j9AUpGnh40W7pSVIG0uMZQSr8LgE8
dORqX+UaniBjLF0lTX3BmL2bpaEviSouC7ln9gPpzRgBZhgZwk311poNTQlpvdTZPh8oFex+AFhY
N4/sZFKEgqBBJC7C9C65uunncTxcmIWh+chnlSDqPnwuCZL9CT8ORp9Y2B//d/nIGiBB2Rt0D2Fx
zd4/jpd6Y/tY8CxnDYgRRLdVAFedjM/VsT8CqlpV1fGxdYOcYDyFdqtoYVdOKzKGkCem/7wk9U9J
cCTR2arsFtSLTfW0tBmWKhfwPiZO0jWr7yc9UkQnqet1sfC8HQ362Acl9eXBFnGFr2r1W7GjpHC/
hiGd7GkqLLwSg8pA1asqM7aqXoBRl/aWK3iMnu1qfk9D8/4SNHNsmRNuV/K+Dsz8mX72xygkhJrD
Jwza+sL0H6OdvryvcZTRcyClZgGAAvMxh3N8tAPkqMW2IpRtsREgm3mBPt7rf9NmQUGMSzN3PoNb
wsBfuKdlKfcMMiVR/W4fcwmTcF6/AXUpqFVkSi9AF85VVWjNg/8iKOZ9//r+k19Zkx5agX8fkb+w
VsfHBiq9VQOS7AMKk4MsLVduFx1LK2l23rjv7SR0kRUdJ93JtnfSrk74de/Kwm7BhLKM/U9D706s
kilO5oD9iq36HotG43HXNfr0edZQaxWPPWF2+oj97/RtpjofuI06g1dZ3DdqwwzoGS6l3JS6n7L5
rqYXv810KvXgvOcU+xTFmCcwD3xHKa/5r5OF3yu/arowWEo7s93NAVRxkmdX5gAR6U1mRWO0Qj7h
1Jw3T9wnpvLfFvxRlUC+T1oVr4YSQvyWDxMoA+HWpwZqNjw5fZ0KC9msCCzUUYmcgbfJKqGSxMIQ
PUM7l+Im1Jq5AfNLkyBDbsjf8bUk1LKu1HJTT80L32tknw/j9wuHUxelieEDQF39MPcR/Wb1WR9x
Gd3CovTyPDSHIT9bgNdQMgHjratjusaUCJthwyTXLGOanYejfAwghS4eRFQ4r/ASabQS+avicFd4
gO+ZY3EPgC7iJvvLn7yen5JfgNo7TD79GXS6s0Dh19QaEQkzRofGiFo/rgOByiIE0ZWQ9IlQRbrF
ZAFP9uEqSwK5auxVdcvaG7VfHb+Gn1WG1qLtxsuKNy9D1BJNdiyRBnyiLwPE03xVapFiBQ41ENpQ
OdIC+yEc5ei9Vk9tZaEPOl2WxDZsqhDINXcLm19MGOwHIgmh+kST5ps1h4kQCkty+GL4Op5915yW
6MhlZ10pjCcHSMz/L8dV4N4n7T+tY+0hEhyacRiQZmrYYw6mOV8zvfG4eP8N0/jhs312/qiM1sc8
uTnjCwThOMwx7qn3ZgXDSb/mimCXL6D8TCX4SwJWaqrWgFAdB5gpBg4/zk8eXOpEPSnRb/ORppf/
OCP1POMhzxmMgqBKxhCh8IhToawE8wAPMlDd114wWENQuY8wf+V+KfuJiBfZ4J+WL47JecthJdLK
S5v+RV/S282htBwtdFK8em0i7UZNfLE0TNgCbG2eYu3Sk+mt2ST8Lb94+6kaZxqwJZWLk7BQr1wj
Dwq6VvEiAst/Di6lF68IXYPQJj0WjbXE8CToGtXX+ICyQmBEnNpuiPxarU7gMEtV9NKXEiA975/y
eXpyupstvhbl+rr2eTfPwG/cPmxeJSTD9fT6J0Bsabq63zJJgf4pSF39eO3UxbUVFsT/CHkYLzV/
V7Oy3tYoLoYaZcQRPn/nxvfDHgGmTyzprwc4UqNiKAasa42ppiPpBrC5zVxlKf0m44Ra+mj3+V4/
xgcF2vzGek/7DEbgvfAf2rHBpfikyLYHdVNwk06YyQPnHiHUDlVw8rDnnYc/CKbi/R6SMa3Ciwfa
6iqF76C6i/gkoipZz1cCNl9HIOXCqcociZHQYUfZuAQw4wLYEtGAXwL/z7BbWV7bm4al0vPlQwWI
f/gg1WSQQUW5kgaJwVGLwKzJ+Pd/nOGWfcXeidx7jBTzIfz0APMylAbikmU+uDjnM+M9Q7Ut/58Z
X6klMC6kS7cWh+jfj+727lSjQuzH8Xxw282RXn7v5aD3at3LurmcoCSyYGp8ho1L4PcRE/X/TC1Y
LqR9fd0d9tpgTHawM9XusxocdxfA5FoqCyjK3WxH9y9tApEE0JDi3eclEqYGbs1qNvM/yDs0HJtc
PW2FuMb4xm3d7K3ryw6uwN9ympuk7oj9XsckpDHyqn2GNaTvHN4jU3Qjh4checp/c9AxSYXkNC3u
ykN75aHdiaIgFHMDIQxm4tEANSO8rS8regvm7b4MitvD/VkEU3PY/+XjKoRd+l29koZ369tRH4Qm
0X0SDS5WIUv8g6qvvQguzbLVW2cxjAqrTUteRIDJuMK9GW4wyBHHjaJaW2C8BKYcDk/zz9qCQ5t3
ScDYuoLzV/kgaUcLcROsCTn4cm9/OyaYL8aas3PUrOl6z6vckhhE60DevcIlaiNO3TGibmYyEjcn
RHQtROx/qh0yMVBVIScVobHtLzFFxI6iaTszl1DIuQLFBNAojDhe2TtsJH4RYl9rqm4P5ZVysX3V
4PiYuauVtf4Ilog3Smc9/48EwNRY0fNhxZ9Tl2rYexSLtam+Rk1fZG65hUczZuGcklpw3/P2XafR
hZhQcqFhGOq2komV1gRyf6hgfVa0iuWdV/hJi+dlxquL22d3oh+wTCl6SPS+SjPAVaPGx7t48xgO
3Vs2NyMSsEd5HdcVYVY4I5slSPV1JnaWiSxBbn0I1ErZqwmmiAZ0i4SQPxA/L/qX1r+buYpMq4AP
AyZQjmbrDh+sYpobRvQTJuNWv9E7FHqWrizyPA9Z/RPdWoMLESg5oaS29K7fjM/aU7od2eaufyFh
FWRkfrWOCEdgYYzXUqVBqS5Y80Udj5nTn3UuFKF5JHFn56bwpQPoL8tmgESyWHo5uXTA4dsTBj2U
JZUV9OMJzjZy1fEQ7+m2E9dNklhi1/l5OfX3/QGKwy/vMwStn/fiZ31ENuK6EKcWncd85io9xPYu
8ORntdPPMIKh/pKStUsO9W+IrVdtFdVd5alNY/z4xvyikALF/JFGHD10LZ+mjr6eOdExry+59T+p
F6ou2FezCvxDxWafGIe7P/AZ4bQUt1sbKovIye91U3Fi14UbnxnZ6AMrjXioUnNWHcbhxnWSpnIs
DgosRWVl5bRhapMycculpc1wVivyOIqT/wIIZDUukwYx57+iKID/MRaEJUFUGu4H0qItEVzhWCqq
iIeB48aV9TnEt4Jszq+TfcWqCKszr2eW2LEr6j1k8ScnI1l6XvbdEDezq7GCSb6BRaaSBIbIuYjG
ymTDy+N3RKm0apT/b+/RhP3gfTY8iLX2VQNRQZB1ZR4D7viN8iEc5FjkUOIZ4na/CyibC9LneZ3e
MYUZg7sREiP/MxBBQsuQlENmFyX9llsBR9euvKwoiZFyYbfheMAmqh5VciMHs0pnXZJwP5UVjh2y
lQUp56/1r/mBfMI/uiP0cnGrQ2JMXCbv0ECyyzo3vDGn7UcZSMo1grzCWC0WkCE0ckEKwBB4LwBo
0vwbDRwSTN5iBHFZwSEWHGI+ZM2K3amkS7DOX87EswTjOenbGNNFd3KnFcfdLHX7WBNRHM1ebK+Q
IvJDEMCt3bfH5ogsnrQmaXQwIjvltoLdztTM9dJ3Tks8aaszwpSJ/Pj2WLv1hOQc8TLSzaOVc03v
Pe1v1Q5Jo1PG0EdhPDkS7kVwZug/AvuZhFLJz90lWMElY3shBZN/TRXWYWLuR6HWcOKLmH+zj6Nn
qoPQD+aoUafIuiRKLC5WdiISv3vMevG+45e2NTnXVhUS9qauAcV0dyk8h7MPzYP9EfdQS7mOIyxD
zCavRL4B3fxO4NQd0xAld9apEaj9LI1IgqvfDGuhkxEg5we1Zuh8T7yNZ0S0UdWqvd/t9q3NUlvH
AOnbqHvd1BGpy51MCVvhXsjXPgUvjM/3y6eQ1+aauH5awHB4KzABEO1Hi8MTRIb/as1wZJbgZ/TS
SXclzH0NYeM+m/dYch6NhPgofUuAVprM6KRVJKp1R4sOKRr/uXP7vB/RCI51UY17TALFE2RGLwE0
z9xV6mAE1xCo4JHygp0fmtDEh/xr1hLOH72527bvGPp0lWNc51sf2GNaiB6AvxpGuG3/YJr0oO5q
ojteOO9YS8FJnStyRXe66ekkHcFSK/4Fj6q8CTWJ9UpK4alWvof7wBDyuvZ1LzXf3gB3+ve8njSe
GYtsvrGTZoJsLkZiBAwBmYzbWQFpXWaFFYG5Sin1ID6yQRRKB05CugykxvlI8j4IoMkhi9LlDqKH
2z8lomJav+gXaXEPVhyIA12wB5RZWYP82cD1co2EkIa3QXeE0dbPP2q1glQRMu/UafFWg+BuTKqR
k/P2VvwcBvzSLo2FDc8Rdot+NAbz7C78SwFixwpF0RMpyt5RzBYzxG8l1TDNlf9Vpd/eNi0+7nIa
J7jQjUhIPbSUwcA32hY2iHFcJL6NbAGIOo9OV6/R3NyYEUJG7Uaw1cPge6I8NBi3+9tkwvAyZwvO
/kZAGGZ+2Lm6Yvaq5M45WbWmwgsfBQQ6sctISNC4flf7n+57LYNs33KjPd/+kWoFhf6l+3qTCIHv
l7lnj1qSaoVUWk46M0meSLhOcybt17RQaQAe4wiMdlNck+sIKoZ4zZ+zsRErzp2JUU1IoiH/9qfG
H1rhX3hERgomrrguLiS9OQ5trk83TsQh/g1XLH2V7ZUEhazx6v/1RnboIdbahLNkaoeKEXm4bUnp
TwTneuFPg3aptDi02vU8+JnjwwIrmZXzx/gCheI9pP14inTyvHnudmA4i/kygWj/sMf7IcnjUHDd
QywxGg8rgQBhfbDApc/Z1ZSGgtlZikt6/uJwVK3fn/H/E/WgMs7TK0eCcu0adtO1EC/00vkAorRp
B7zExDQSo5AUAhpFXRW/Irge3rUhAD47iatmPZeDd2UaS7EmDX2H9UOYftYLK31u6zF3v9Ox1N0/
k+Hq5UjiPL9LWDRgGCn1CRMFrJ1YvZguyQ9NTKWQB+qRGS1+s/tdiBSw1QHk1sDvMC/NFiWtBNOH
bLCHUogiL64A0OkGQhTQO/43UHMZnPfPaZ3hPWXHs4FSmE9a6uYU5DT7pOXWJB3xt79BhCG3Q3Mx
lmDy7gSrXaG/cLpsGm9efUJFi3Kaleyb2Hk9ozWLPzTodgvVj7Vwb7LwmO6LZrDSpV8xAm5Cymfy
ZB2ElcgJ3llaPa3kS9n0o3rj+nVOmolU1qvEV8hC4epGNcQYTutPodbzg2rk2eyJNHHEKq3JjO0/
brrWkGJXId7UB4MwsiJvV5J07gY5c6E2faUm+AQLOtIWFMMdAF0QQQzZK/2l3ft6//ArdAYQ7+XY
LCUCpYnnwjaiStW931NT9e82ULryMLlwF6oF76clDYSy4bRivFTrjpxdQgE6dsRLyke/vy+qPEZU
MGKXP0uE43D2YSefK+uRAxaZEtdBWuQbw3RKOVvVVcFW7Ui9u+Xxw4xE8h/J0Bl8h7vTT/OunUbG
spwLae4rl/V017cc7Oj/MgxHeVIwmaHTUogxbxuiBgBPM/L3dn7pH8CmR/Dsg5JEg8vaATtooOF4
grAkwFX63sZ31PFnPj/qh2j/I/lcyJ41TX5BpwpCzASYe3INsWcYrjr/KOgHH23eHSbk65Z6b+8u
iUSCZaVfyhrkaPjpIDOqdsBy7rfNN297zeBKlYKmiM1/5b9C4jx2BDtxulggXXqefPwjT6tbbnZO
eqmb4DOt1zW0MerQcpoQj7lxFtdpcavErWLLtujHNjzZj2sx53gvvD5pJlJpGOF+6bmg+xHggKqv
N5IE58CIMHgFeJGvUyhkpY4oZIEBw7nNYMWRk+5H5rgGmGJ36ZRiT1GwTAeqadfr3Ly7HcG5CyUk
5bnPneW5rBuyEzHLT2IXcDxtYKJglbl1YpfyjgvzWQS+4mMYkL6Y/jeorAXvctEmTvk+BROucPL5
eO427uMytQ6WTBeejj7T25i4P455HOJogbPi9j6IBH3m/5SAJXuXy8xVdKHPadx1XwlMvymsxy0n
r1uCqnphNUJBJpSRozx+yMiirbz7TZDWPlNmRDq4C6FhTwViy0+PjPPr3wzET9czXsy51Af8SxWB
lELQMoWqrUhTIwKcP2SQo0Kav3Cldxt66uvV29bg+el02e5yS5ACQ5JoJ9VaWVqQmS+DcYPQHbd2
Ugi9QmEoj+cf3q+SuNBFPf9aBxL5UC28cwiIn8iIvn+agywNXD+oQ3SHmxymkFQR4L/2cIsWJrDX
3u9cUWgXnJoP+0WhZVW3GoD2OD8EoYdD8JGARC1oH1dMIZ3mbxaDhZmLJ2W7E/vPfe22nATFudVE
aJxWtintrVr3bAdxDHFew0F00rjKgp1jhStksVGOriw6ZlC61l/kq/r4P+AxTj9wVkqrMs70Hncw
ZAD6UPxwYiKziu8t8RM+YJNIAGDV1PDh7C+14KdRMSFsdSu/Oz0M5Xxt8KakmeucrriIfmZC/PcA
GV7YtF7OjpdaDHYwaadvDCVvXnprSMXVNCn2aOdueE6nMpFDHhUuJgBK9t4Lc84/Q9zirThpQexX
CsOYYhTYtO/jOvFyaTrUOMdNK24nQsWu7OkKI6rVMpdD7m8AFSVZGqbxx7MdC2btnojdFoQxC8+n
+PPmtWDm/+aFTXM42sZx1nzC/MWd2lPh1wvH0OWmP+qSVC6od4W07VOPsca66u8JWnt4bCM1Fd93
THzkMSsBR/I6lj4X009fCAKVYj76sQwpXql/FptgcgkZBMSBr6PVYp9YRT/Gk3ClndVseCsmbDQ3
AL22PfREO1/Sz2hWh7Zm9074Jla0pYGqd85pu48Rbb1ZQkp1OdJXpYLsHHmmXKsgTPNXQvULR1IQ
V9dMHZvBbAt8zHDc7yeEIDnc02p8WWOR4DaHuS79Bqsd1jTy6wfC3N0JjcZRUItYgnB8Af/p9t+N
yqzSmHhKML870+S7kxvq4azw3xln0qg8jlCZrsunDesDRd80W0xDdW4v1EZumQQgfHSgvkkDrgWI
FtWkB98rXnVTK/RGgSndXJ7SmVVMUQY2+dSsym/6PW0jtiXIrHfP9ganXOUYuEzawOdgCaleu4sm
baIserzg4FQMCYfPFTEIusxwTmr2gJ41wJEB42RY3V0Syxl+ezI4CaQzCxpUQSwNzhw81eJzd80w
B2XwP8OnetVQaj1DNrmI3XL9dog15bFq0i9FHKP6SicA8cM4IRStcZkZikP/nT4T0DQw6eJip/f4
mfs8ON9kDLCJq5EszoQYONVlzAFrUCxDfeYFGUOMuuEMCBgMAAKI3W/+GG9iNF7m5P1pXGAakxTt
o6KHe1SQbmD8DhShAxWFHNvL0+vK3LXavmdoRMHMbWpZkfITkW7Xx9xEffbbCU6BZ/9C85sIYbVd
NcXjuXlZNGjEvn72ZPkFO7zWl4wcD4giTXU/fh/wVn7WKcTkh5hJKKkHHsgZoRJK2Jb27TNKP5EH
iu1f8PtClbvNqOpO9Z8hfq0WxFS1rGHRdaK1nuKmIqHQofj5o1o83VGkybQtSmRmeDctud6J7JyG
Iu4pCXJA2rWgsN5rwyPsavPrN80XqLmMtZ2bxx00SEk8iaiSA2bEA4+7Ay5VM8fforjblS3LbZbY
5Pac+ER1i7v5L3SLEhLNco/2E9IUJ82lOmQ01o0i0jJQua+9lzZf/6qVrzf7ASRFM5j3NOgW4Iag
5CkC3PrvKM9+fy6mMhqZISgO4Ox30bLtYN3Km8aVNaPnCVmORaLJT4Bmy0wUvJZIu6xHLPcxCdC0
kByV0lrFwTY2q6jspNvPmwFGWnWie6H2zwWcKtmxLlDG4x2t89k7vyl9cyuGuN5TUJnFn9KS9Grs
KR8ld/3XxGjxRx2R3VGy05fNu9wvavumx2y28jVnewawj75hPg9dbctTep5SGmXUeEAApTo182w1
6FAb9kYaMj7UoxyAf8gau2o/wfnYhQFXHFcQFPnnXN5tuw8JHQCoq5yQ5isC4uPNlYDIzXw0+Fvs
PZllDHbEULVnYzZJzpaFvG5K9O+nrhuZlMxp6o4MwIllTumuUbaouy3w7XH5BhKwT4tvDoAT7xS1
RMuTgy5JvzevL6xUZkMM5btJRiSnrdfQXY/RfN2tdAfffA83zBOn2C0/Z0c96uXL2pQWkMCAs/RM
oojj0sDu0ERG7uxiLkoJfx5RZpgHjd0O6NHm95dfjvtSz8eePCLEEuOIG35I7C7J3lgxrOV1wlA8
EkZKvahHpM17eCcSgy84UzlPqIzAowyA//LvBr29xSUa4e0XApkXeG8NjyUlo8707NIy8cCXQh7y
ZwpA86fmX0UxdW6q4uKG58AiKjuj4ux6wMenwQ1vovsN4pjmJs1dAWG6sPDqWLqK4rgfCOwIbH0e
0R7+BuLqiXzypkRny0WUWTyscCfiyYSv7RJpON/xD9F7HtNczP85fL3TLlvGGczbC0M6m7U0DFyP
cVaNFndg59UmyLO4nu8+I9kjcP8fn3sKN0/Axu7UPvNUuD63hFAdH8cN8aIvedq9UXUzrphMoFRk
eH8MstTi38lfULcg8ppJjCbDWi8XYbpGbru42oUkB2WmgFpNos+w3Z2dvX+DWStLjr5i0spPZxpn
ljjIcZY1m6UN9+AdugwNh+uYswkh1qt4qT+7hQRIML2RB2AbgVpcLwAAeUnmKxKGpgFhZutRYVX4
0lNAXh/d0LARt6Q9VL8WC7ttndXVzVH+joUc0aBaLZCWoNP5qGzmQOx0v5opMbzoX0jMpLE1AckT
mPQD4FCN+Mw3egC6MIf1+ukGfi3XI4n5wC9cRrVl3nyKZkMnlShYSHg1BQTKx5EBx+3pPu60B4M6
wDiR6MEGnYUNiKX3MbQ0XEpNYyuoPPI8WjKcFfZDybmjFpv2pR+Ll0LVIVIvu9H16IidRJQaY+Fi
xnZzA5H4GN8m0sddksbtc82unXl+QbHm6D4iNzswvBbZO1mX7oqtDj70w6FlIOXofAXKJzdJ/v9I
AP95yPhA1TxgM3DqGss95KyZgQyMWYz9UmhV1JEUYB1RPxMFPM1mDZ/dquBRx+dZZwYuy911+lcC
iwbl0nUBCl+SbZCDAvFYQUeUhFM9YG1+fDqOLiBRcAqGxJGYbS2wEcvLdy7OZCV16mRnGuytzzW2
1qNZnF+39Hp90w8S5FHAap2YA0ip9E37Pl3JDU/gLOtnlSriNO1f1XNQOf+QHBjTl+YT2qmu/6OL
KWF7cj5onxJUeJigHqgRsWz712Borv4jpOt+FgRROaRgl5MnNGPkcebz1WflkbHGpje90i62K0VE
LLS8OawjlAAlfwQHRWmjm5nRVVUVdrv4kEiLJoIq5XM4BrAnp4YAQ2eRK9hsFvA1WbnH2jYKK5vf
0oFjoRNeYSoVr1XpGCtJbRl/Rbpge9fFyiF2L1PgeUlI+uAUXC3aENEUMp/PPBQc873LsPuSQQX6
BrmjSxfM1PyRSLt1N6odzEFJTmX37mHCDscBvEMpsVpMO5tczWfVn84hXNiOMW65IMnXTJ/JdOBt
kbCrs5BGfe8mLRya82QlOR3IULEjn5dLsxKCM95Nc5kM65yT11WWmjZ4xfalgZZKbSBLsWNM/kpL
Crwb4skEOEMHUhawWNCSYLutM9Hhge8rzUuJYn9MMWV37a4XVO9jsGtTvk4IMmqyp4oRGWQ2Qya/
2RqZ10zNlzui+dQiHimyspvfpeXUjMJe+pVdpDFV2QXBDRh4BTjMNf3sCJ8GzliCOr4LwPKzRbx6
E/fY+Z8OD+5fmSGBqkU094I7sdFcTaNP4N/wYHqjtJbAqVAJZi7S0uVAn2oy5V43+nP118lkd2lL
fWCYnkfY11DQTGWcHkOALI5uhOOCULkAau8SPGsFBS1ns09+NddnuOudF5n/zdrlXkn2eXTuduAa
CS3LwnfO3ZJ20K0oPl8SLU5fk48+J8wDMB0jup8nbW9/MGrRohwmUfn76DeEHqWsvVJra5twPhMu
an6DhrMm/rEAHQJRXwL0OHAzySMZghn/nIiBFFmUD5h/Lh33xNHORKyyjV/ktHQFwhaRKbRg40/s
wXKlSBoZqHmOf4kkIflFq5nw563oV+bqzXZg2ivh6/7t5UL6yv3fCfweX/QYbXdN/72ImbtEuxE5
QgbiMT5gHce8TNZBUFcb7VgRcbS47MEEoZmmPC8PXkBvhpbIYKh53ki1iH8uaCjZLQLi5KhtAovo
A/iQQdhk4MW7Bel4H4yJVkX8b5qIDwj4QOH/M64J2bwsdwNPszWRnWpEU/vaJP60imxyvNDKIf0E
Xoe2pa5UgGkrHoN/DbquYxEeyfcLZfEnTaJCXxHWB1bh/vVtbOO1E5QpWXUrp/CvEZVaDlrP8muP
Ro+PV/3bAr1cjPIyOFJz1O4/0gg+yWmPW7dLEaKMwLYsb3Vlbsx0s64z2U/rfXUCKdsZbPtT3HBO
Ur34yuMMQ/yVvuzt7ZOJIzekb7SKUKo1hkrNzLtUjcgW/rTQ99run42qCVn71dAJ6xTZwAQI+mqI
Ez86sgeYgGEithHctz7PvF5AbPFpacSDQTfm7y2XQSEELCC5I86xH1VSU+NIMdDQDLfnjQRK0Bax
3V4KIeFayo3nSRcEhjOOrro/RnhiGdgjDrJvVAOC+4Fzqelneg9/1ZmmDzNACqx3GK6uhK+mP/ce
j9oaGOWTHoXQlcUOSRhKRp4IxcIOif+KT589IfJLT5/TRC1xHv35hweYpp8bwG9VWhZ8f2saRWHY
zy2gFyY3/RSS0zCCB108ABFZnIlC7njJIu59+x79RG9xLkTOUdbM6TscQ79vMWpX1LRg8YXlfjAn
pu8gVUjq49eLGw9Pi0sSDHF7DjmivtNlaiM4Vktr8FGQRVdrkazlgaeR/fcN+jcpcl9Y3InzEe/Q
TxTtwm/v7pwaNEYIbnN8+u7uXr67NsrWkyahazMXe1iAG4s5ymbbbq5/eucmUpn/0x8o1HWpnOgb
mLnfYY13l2XctnYwPogJU5qhYEWB7AYotJ0+kE/yi74VFmVkCC/qJhlxNDUrjqYPY8kZEDk8rzjf
19l2/gXG4tYT3wLwzZs0f5xwluq2A/GUCixwGmA6sKsGYyqOGVjXwPsDnK8wzGdSH37U0pkYLnQz
wYnqYUoDiNAqkXLKD7K7Pm25hXyBrwPg6h8VVulDVFILphFEx/qIFBYBwl422fxHUifHgwfuz5wq
ZtNDzyjXh/zYZJa1l8u+SyiaKj28eJPDMFKBWBj30cx1yqf1JOwvKRyynR+iFJIn8n1qNMNHNu5J
3wHla1aXI5++j9fCuA5atgTpIrg8Qp3kL01ceKp/jBKMgCPdYZ3b5hSzbxahL1mwiMWM5jtUcIbn
UxmetDp3hH/2839ihj7clqv+c6i8HwZxYOD/O4sfInxTjYHMr8I81/29sLy4m01/WOAjqwEBft0g
Vwu69GwO78277uKWfksyB2ST9Zc9FqmQf89KmAr7O2grI7eMDmlqW/NJI5Pimd++oCVg7dDNq/4Z
thR8vYATYwrB8NULEt240mgo5Kvnz3zcCjPibQTp3B1TYnHmSdXWrJiy3tkvLkhTBJ2FHutpPIsG
3j8gBAoDtsJvamu7k95Tr8KDi7ybW1Ry+oDbjp39PTVicpw/L6fFleQvZSsrrGf+helx6NZB3wPC
NURGMs6dJTXvY0kOR6l/ErxGDFPQzcGLe+gTSmxcDz0RyNW+19A9m4v235E1C7kkLedxwqPQuobV
cwUtRXPyq/VhpFEhx3UEOKMgoNwZm72TPv/ILx7hB8EGjdQ5ozpmXT2DywUs09EOydedCGskLPeJ
ziK2rnrpv7Ceroe8in29XtWOdqaHb+SMev+tB+GFZcogrMHZ8LVgQXcchuKrKJXjjHfFE0sv26to
/+ehiT+JDCGSwMEJqfFKheMYkwMWpfTpGNQO0Ptmu2dOUZ51oHwd0IlzASToaCAT0/lv6OFfHo45
YgRS0bwTgSWAVvJWEnuiHnmQWX0dK2HxNiVOVIRAaw3yrejVTReAoGhEzI0A7X0DnpmShNhHjVzC
hKyn6NQQNZ8v75XQwKOwZFPHVgGLyaoHATrLjqreoZmEAVG9LvYsTEZP8S34qsoDJlWsjfHZaIUL
pO0ErZaSpBodHN3opGOUd1yP0+pnB2Rg9WULghTXhxKsQis2ny8ONXXOrGHhJf+uIzh/ymXT27MW
8Tp7hOVcZZk7Am9JNOIEnlrAzQhKc2HOo4i5MW/DyQxuKalkpS9lQwUzhURMTxjtiPMRArZAewsG
2XTq3T6U72eJM6kIEX5Rkg7vFd6J6VfpmH8NzeNHkjcjyJe5+6g0R5YRO3JJW3wI/ZFUfjHrNDBD
we0mV93oyN0Gv0yNtwZ5M4R4UjuEavoBK/U3UUfX5mI9k7Oc7op80WAYx5RQ6dAfiYB7QHtKtKdS
U0UjUhAAo6u+Rpfda7QWgRjEVy1DC/tdHFOIZXqWHvestCTAIALlSfTPSnW5rtYQg8DSkNqLzX4Q
lNJ5kf27bQx0s+WSMaCOrzCn9KQ4aIQUnXdeAhuwLNzhOA5TAuYl38vhA76I+QJWX5XjrEzKgiKY
wVJkenOucPhKmIGWbImbnDMFqfV3w0etm4w5j/po6GhSF6UxgnUQw5nulZr5hfVjRX9rhBfH+0/k
TvKIPPC/vGquvo0LlG9YQ7klSrMY8fwfcfzYqN57QbkMk1PKHTRE+BP5c6NjzuNlR3d1g3jStgNC
Ge9sNc5Z077GE33+phAUxqxqAmJJo5vqmLDVi+XNwe2NlZ6giKjCJLdjdz1R6y7isT3M9G0S5tBM
yEvWiatFYqcY/gOp88Gjam4kAJCC0iSRojveFHaC/WGTPNONdgyxS8XsE5WI9O22ysUvjYVAZhO2
x2JWpHzlSwRdcorsRm2U7tMz5YIPBNAjUV/iI4qyw3fn224TrTc6mylxmlYatmBo3Xzd/TekiNRT
zJ7xwmyioXRfAdMx96Znl1+QOXuqnu9Dc2RYY+F5GqvelJBzDZFx91UxjJ7Vj2rJsi5bvmnJYbxz
DV7umq4m5RMXpxclgIlrgO1nmjrr/JXmglLpUTl/i6t3Lds75oxsr37QMrKjyFlF2b1Q0ZHNYAIK
oihX3+KKJkz+L1YowYwTbSl11/idaHKvqrfSrWRV6QOaNH5+4ywtzzK4Zt4xA8TcdY8wt9LsmMuL
FUcSJOKev5ZGle2Yff2+FX+WaCstiGgUOFDPu1kKfmqlNQdLPsvh6HNs1mZkhahCGljGzFQxmjUx
tSoeuMD4hUZRPMvuR3U0rzsh2u3C6bBCuXAWFOu4gxo+11eqjwj8fGMU2YD5M/3fJCY2JDhJ4nfT
UbEPy954v5/FW6pz0m1dXyYu1asllEND+57vZWj1cYo/HMFnF+chv/5+LlaOkLEUdTGA1CMxT14s
e8zHgU3WaPR71tE/BKLQ8pLvQevH0WFcfIp3nBQTGN/5eUfW5moR7FFmVxkKmRwDvGQe856hLXAN
Xoj3eJqFvk2q15wwM/O8Pd8ZXsg9CPe2sypp3qDsBebehWpHYdpf2KD1iBamj85wpptQJkpei+lE
RzzI37kgv3uON5zFMej7WjyTdFAjmGgsWrvmfyrWlZ84OxbXBmWGvBpxmrIcT6yCoerHWjbReWlF
xACuXYvcgFDLQUjR9xDgH80Gg9FH1MCaBODsqoSuKhCY70lm7tk6ESqKKEk/n9knaGp8H6AdYqoh
p8Z6ZgkgYQIMCycyJ60qhCJ+CC4zTxQ6977is7V6JrbUfdm1wp9gQDC7L1PzieFZBACey1uL+2+V
nwkpHF5rgyXEl0YjddSXai4RiTw4n+64pA3RZYy3EoV/T3xYV6BlIud9ChbfTFwwQWhoulMbUma5
NDwkKlq+m+n7OCKpgPNzXhmsn8VgepDkP5BUKfm8VQUokiK8g3RU8RYDCgwzehjirsivCH9pp2gs
gEXfXqOnYsyCML+Pxd1KmiRGbkxXSnAlwkd1O3xpUyr6cYjcXb6surT2rl48QGr6S1jAJkWAzO/B
PCZ/vnFdInj1gPKm2FNqIp9uUP1OPW5gLWphYg6cPkLizVoWsSZKKVmuZBpV2OS2XFtgbrAQlvh6
TvkqwZMtL6DJTqJ6LBjne+sTJEvb6FzaaygoEMIKhlmn1lBgdzl+8iSu+EtTP8MIH3nRfvUsVKKC
FYhX8xHLliWMmgZIgWgvwGjtWPRfWwjZlXwHk9sa5WQVd33N95W20O7qzxJw10GYwlZsadjKxnLw
WcJ+UuuRgZDzd+T9cfAAE7eBp6Zp9Dj61mh8QMevRel0afrB83YLkK6PgE8O8EtFccKHKQcalRRm
eviVth+wGkhvQ33cZHlRc81DTOiLWYUYRlYXKgsBbZBBEZro9ZAL6rkOJcneuYqyuov7jUIeTG3+
GaDY9IhXvM6vNXak9JMPn3IGh+UwpS8Yxg5ij3yy8vwY6+FjgNf+TU+8oefFPzuCGpvVZcJAtIjO
B3tF1KxuiMIq+WqlF6AYsLMt8JrXCjJ9Y9wWWsqp+XXey+2OG/6R/A7rBMb2BG+kJl5Bzn+w0Emp
C0LHc0b5pdv+sBbREIszwldpAcdG62UwEUHWSBT2bwqRL/BLmxFmr0krqd1K5DZQbW0fw6UuBQpJ
p98mv7oGGD6I9M8pR2sEPnkQHwL2MU9Vrbo2th5tb8gxIph12k9fcpHS/Vd89dTDLD1uGTXm0gza
EiQZ1WEy6qqi6I6HSR/0ZgBCO7ft/kjywv4UcpHmURvNAu7FPSjJpltV0cSsVTdwrGu/i4yHw/Qb
VtKqqzx7kakPf2yeLhADWIRuzGFLYj0Mxt3oJi9fSHb7FksEFS4d+GiscqYk0BjPkuUmJCjvjdsL
wleF7n6UzRwbjmou991/jwBC3AiYJjHRbJ7+aGyP4CkmeUugb4Qod0IyDZ4jUZvYOA55bedtPI43
yWNHY+zRaSb1giuq0ALJfQkjyz8m2YhHNBRxjwIJIHOnqMpRpFamukGTJL5GpW6JAEn+h9Kj77YL
YMrtqY6g2/8moe1XPDaK284xV+bYHcIA4iZGsLLjmMAFjcwe5swXKtTaSMI2oOwCbKb8352rXUl/
8MSEflH79h7tUNR4dMblm7GvgfzYyn504fI8V7seaS0xH4YOyld1w5CgIXzBKcT3XW31odubOZj0
5rXxXT9TF8Yn3ZbnZJhbdNuQzalelwO+1Ijb90t2Q/i770cbB8BArtLAeqUK3bSH2Cvzmu7udxgA
UPQUpIjz+RWzanxI+38RSHOMw6Bpl7EycpCZmMJpdHTPmn6ppCYmnoECoBH0iEE3BEAdlfK8VFxh
rc24mUlxJqUHBNuJqhoUlfZ6q/VTGj8uM5COuI6G844Za3u4wf+yTDZYaVQ8hBWIb6ZCeSOnb+S3
eUxlu9OnlPHabBDCaq9BokeujQLOfIO/+cCwzJ+wu4/BFbrm0cXS4cvwGU4oui9TpKdrS2QisdF0
zl35jcKje+FZPuHQC0/UtOmmk0Zxu8gFO0Vzyc62AYkwNVaLL67OC8Dcr06ighCpPMyMIsbMc+TB
vbKs5F7UvomSG2mWISX1cEYxKCRxtZmougRq0/ZIcS6S4ZB39yjYpK5UGlCfw9xBqrXbg9IJCqpX
pd13Jgk+4W06sgBgqWziqwx2/ylIQeFSbnOVS1OJfvOYc4c7SZNP7xSfokHisDpeMZ0KYuhrkRVc
qEbcBtbmB0D2HL07nIWo5jh8h3PEFaVbOrsMPOr+yi+1AfYOMr7cYaxAM+sNYulccecxre4156M+
55l4kYvciMK9chqbL9DEKTZHgm4sGTmfSBPK7J/g58ToM5XNfvymFZkoSQu0GI1ro8dohHZmto7C
kIQVmsELk9n0uZGoDpL7TTvzAHsSNs4tZ9nBlA5Dm3gfS7NYdGa7clF7KcKkaQMmcnGa7p0sIFce
WfvdjkcHYn/dZIKgj136hI5wrhjVuKQ6HxYWSZA6GpTfVOTuyO6YJk4bLjam29V7uK4avfI6f/F9
X3jy67jQiCi4pSN7Gzco33k7WvsNHqLIDBcWDCUCSH3b7xacNL4H9DYLQih7KK8eAxte8O8YsFWd
OrWPNgwV7tnDEI8jYte+scPkFvtqmXPvOotAxTwNeg/r8bEW7sU1XSNC6Zv6Ip2RA9anYzykBzqa
x+M97Ex2fxqJIGVY4z0NQaeAkm2xvDaaBxN5QrjeMJAhwUHSbkTBwS+1qTp1QGVZYu0Cg0ECPj20
02TdIpYfBXg+MRMsk6ahE9lc7b2ow/6YT0SnPrXnzxl7zffv5FYKwMCTjtbeVQJ2CuCOipLCDaHP
AAENIKCAbbVIPDn3wQA+baRnZ9aAty/8z2A1PiWoSLle6YVg3tzARm6Ohbgef+6qYoHLsKagOe44
8w3w721OauhmCoSyWQs4XFpbh8udz8wUjPQ6mHt81r/SRiHFrRdxSikka14q1vIvnsOj0retx80Q
dD4sfN5kyeA8SzbG49C3mGvd3h+wYJVEpqjuyQJoDzdk3boHWdtPkBly6nFti71uiUclcpVSp6hb
KhF6eekA7+Z8Hpu0WL9O3+wZHuYeydJddblIXfFiSm9FB6K4sFQc5W6/xmRYj86ODn3X1pXFgSVN
jarFg3ZBFN1q+qu5OpbZ5LbyFm6iwLFBY7/Vi9YyD151G2b/VBJULKIvLYecshMdMbfwKiSYlqNR
T8c4XIyQsj+9y4kVB0Zllj+/9NakD/Wlls2fLrVfVbLlFsI7rUghzFoM8FRLz/9EtGJejUEAYLRq
JOYlDVwDPbIRjNotczV3UQBUZLaCFqgyaxGSSMMF+ZEZzqrE8ckWRLvP3+G4rJNd5PRJ1yqNicWp
YTCTN7vzQCPaVdsANUNuuqTuwpYdRR+NBeVjvGYfIsl0s75R+d/XZxWmGQxLvWUA3v0f/QTySa6Y
FK84ur1QDIQLslx/VknHn9Mi5DbOMcKZnU3GSuPnwdBB711ivpge/t90VAhwvPDIrP/HT0DzJTZK
1pwKuPaoHPApSRY7jtJnIFQq7A7+aZVqzTNR97IKPqxP1Ijt25duLuQxCj5fxSuX5tIWgwbhawBm
V3HzZMH71PmHi2xsfGODNn3L7ciBxthpxMrcUTu7Up98tOpAcg6jsJiHOSNwceR3H9DD67h/X/E0
9QUzFW9JNOm/OqdnX7+LsZYwDGGuPct6+ihUqN9rHBfHmtQJ44OcjEhe901UvERBRiEeRSGVomAG
zLXqsaN9zQ2GhZMP9ZcQyrGGZrErEIDvrGU2FUPfAumU+zsazExsJm7rylE8AyYRe3QKdeSnRa6+
sULpVoHGYfYhJvnlOlN7wI8eNVV9bjsxcCgwbhWQUtwKCp/AOv4ZIjaJuDwgyI1bSn9EBMM44+MV
fXdUuhJbRgSQ+kWvCdZJqbTU/ZN8brlcT1klGVOxxXOVr2RcvQS3s5mCwVUQz4kEvcSLTalDU71v
ikKBy0qM+a8gX1c1NVxSElg3HV7Z+MtlsZbld64U0w0qJ/z7pONj8RG2U6F87mk12k/jooWhZ2Rn
YKqJ+T4FlrR+QMmVBfXsF5+5Hw5gUZk2jmIInczjIYhk6JSmaQmQPofZnjPy6z2ynwXAhJTzzFS6
qahVhZ7AeQLntUm4rZBqOgecBldawJZ57ursx1E95VU29iPD8uHBbElozXf7L/EfjF9hHIiMXeAq
cZD0EcRFBFuDLPSYJYJ0qUi+6vPFF/D5AOyvZ+GDHOeKrMWqKpA0q5mpsoTYvZch6MU+jEn8yByB
cI7tcJLI5CGR+SXIMqoxFk0fa8+n9Gm4DM/WxPvhha00XG7xqZA5vOJGbiZFAoNhvQTvLwvISIT4
D5uUBWZIR/KJz/Cn3rKIFmqSLKty/WOoJh3ZVlFKEkjFqT20SZ0EOMj/a3Qy/B7ON+9PXZcfTlJd
W/uH2a95/a/wDCa58m1yA5E6uuwUzUa9T0w2pxdxIJuhjd5bkHg89yxaUriaxGHYEOLcstfZzg5p
taNpxDDV6kJ8vU2HrtL9UnZp3TsU8lY4i/+It0gYoUxXGeiz4PLCcqtFx2s+WMxaG7CeEFojfVdj
7fb1ughPR55Ha7uub72+JVma4FsTZ3JqBXqBGVSNPbHuAD2Xstmja3VZ3NEOFuviftIGpP+UYoNu
kyduV6tlfqoEYEFVVtfWbj0mblFyOBC604njYeFyNPSYvFXO76sD9mmxijpyVqKPFwDdkc1PNm3s
XJLpSlGXMasFTBJZHZEvmzrjd7LqhOuD2XGsjJzcuCmVbYsx6kidBSDrHxLm3/q/Iq95j0QeWZiZ
1Wr1Qjz/b7yAQwHh4pW7Q9tJ/2cd8GQ41d7f2+9llVOAWK0EYQXl4S9AnokLnRSP5/sxddkU85sK
bS6W5tQbI1srnxBgdv/9drStaGes3EgTJ3qdfI5HdBv+HWgAqBp1O4hWaRKKEzd3F5vtTyjkWXb6
F6t7MurVqkqJrhXXYerqUzDjLEUzbnc1abooV/HSHTzk2R4tz0YULbA6nRKbwPO/jNU43oaqKzWq
qxVffJKyqvVTAnhjjDn9yiPUE2Vks92uEz6CYYj3ytbT4YaTvMxbvyfScx6YguBaR/4fmTFB5va0
OeCfZ1tR3FgI2VpnF2R2KtgsH5APBtskAm9l0pKzm+tIMNzx8KSdYXXsDirH/P/dsTn0N3nGq7ma
EpiisgDvAKgd7+KMVMCu2ayLUKJ133UQtgZpAPRFtKOGpNwDH0bgNWlba9tF4seaQ0bINQ8JdWRp
0C7+3uid7S2rdW8ipvTIIzZ47nRxbiN7ukGZe5O08zKJp9Xz/YNtVf9y3WQUnBywFQetzscpckaH
qtuB8pFHua30fMiTCnAzZxfwU32SHciLC8aL4AYf+a/srQZ5Ubf0Lb4jyBJToPu69tWJPWf23kwt
OoATdvuUN6o1CGC+NrY33PwVbnvrI9Z4KH1BCVSn/nyJ7jNgjgjKLq4hNLr0demdHjtoKU1SuoVg
jBVN8q1LCGB/9dOejrdSe7/FjjgRQode6f8XH4u9e/V5LQFE0z+BLMQGZDO72/2Nx5b7KXugUe6a
S+cKH+0CwxuT3UboRSXesDqUVuXjj0qPA+HrO7yudxtNipxFgO9JuqxJyEV3bbl4JfDF0M2PJp1c
gyVqj5nucBTiuGg/0zoQMf82HBcDRDydmwYaCNYc7ACGTIGrrJidHnjvwmfYaGnTTELtSJ1/cRts
s3Qo6Uea4M3QAhxpamCHMcOTvLgFltZcXWbXBe9VJtrifbBL11v17+7AZTevQhwThZqOTdmuGVFy
ekhdTuy0g5146dGj94MVxsvFWb5TuCn9Dr/xWg+nTO/2vhFnOV+UyRyEr79BoVLqOnv7eR7xo2ua
yTKePBEYbmPAeEhxE+yoezxi8Lr+dOv6eNnQJ4t6SIV7pqVxcofvdtx39lWcYL4IPSlLPD7UJGy7
wPvs8hqqECRkBTIUOeG9+qi/j9Atn+u8udHmtdJBeGFi65seWNOFT6vXZLWReVxdlt8DZ+qH5n39
PiL69EpKVGvSvAn/zxwXdYSVrnJfHTGYB9myZw1+7ETgm+XjzyI0mOfyj5n7+InwkQ9rBuTvIiLP
cL42FQiGleemfxBFBn+Ht3pwof4HYfm2Ept9qsx83Qq2Fl96bgq64CsQPt595uNqKe+WK5ydSNWn
ZDfXXVdoH379avZA59TC+d64RhvLsyneXH+XiPH/uuxEu7b7S2XP1LsdFQO7RT2rVCue8XJEZDau
V7jXpLoS7K+yPo2Klz/f+fCnYV10KbOtm7sdEtRz8rEcl0PtXUrjW5WCKCR5OVD49ly7yXpxvkca
0nH+sOmvCfd5hvcYZ0HP6v2biEzHlsJuAQpUb0EF6zfTY0gziS44LG0RdaQqTJyb1k3aB01ANHWv
jeMkZA9qj3bKnSu3ihuNXER7OUCGZ+NG9JD5nPn8WL4xPoxZNyL5zsXBfshgOTp3b0O7b2xjrvER
daUT85aEUxrwVNlzlVFTSvmnel5ZdAInREQrjzMNuwuOzOdD7ie+wPOUKThtMmvR/C1uFor7G6Hw
EBIp1Hn5gzpPG/azxFCxr3aNTHBvJ2eMDE48AGFojRCSqlRfIY+prnahbYoHmIiD63gG1b3K8XNb
4K5sUaPBA+9dqf+Rr7fWyqvp2jTaCEevPHorgDvB8BNcllKIoPkc2roVYAEHZVGRokxgKdXegSkw
RqN4di5HqCL7NJcm3J728P4BSwnDwPFvJqmUYJVPKFazS5e+HXc3SLS+LEkpAOErCGMhM4hcOj9p
t67TcV4SqmEJ8tzajxQQA7fYDFkWK6Lx0dmyCboWjYK/2JggCWF/wEw0MbvXsEry3hVuVN8jbUDq
eBVoyNj+KOOmD9BRBzsPXZz1Yz7log+ScUmn3VDejykTjdesVlszxXh8rq3igz85gCUbjiz0Muv+
3k2maMNTRgQJfjrGUNmpH1OvDhLe+xyNs/c3AWwfayaXjKE54wQyqGY1LRgphPV7TFN5OexoLblH
09ij/ZvUIMrjeZnAOWBMrZm1GTnu5QCTpa1gTJ2M8g3TDnVnlXR5pXvz/43nOg8eyOvLeD7Nmutl
VxJlwjCXg0BBkYRYDZ/ybN5qviiZt7lALTuU+LCz08GL8aq28KjWMz2S+HdzojO1WCCciX2XfBlr
qBet2xKslF/mELs1SUjhiwS8T1Oo2VmodukSuBCBKnMHrCo451mo+k8+cKpkRJcqTe5m7kfUabRa
w1Xjtr9CdkIFvMdpeFcAFeDMt1ZiGojbga+m2WGvwfV1EhGTvKj0/+L4/NBWNrBRI7Sw3keQWCH8
1fPeaqkZB8nBOX2UweuqrIx13BRrcPhO9hCkZMoub039OJC1DkzySrrCUssp9+BrizZlkpDdG0OY
AOX+OHoIytJQhf50cdoMWkacfoGE6yYWDozFmqaoa5mc23qekLFpu3msl7x0CpMIuq/jbS3mEihK
YCH3B+1i6uT5Pww4usXi1Uij6yKiyS1N/Ul/PcmFwCt8wcksAPPZQ79tvBZE9QoR/G6dF9RreLvO
x5XiQXDZJf0YbnmKI4yj9aI5YIO63ha9zjnWuieZ2AlMdrSP0MelFNwqwi497YoiebqdjHghG9+j
rH5c2q3L+jQD55J9dxn5K3SzAOz4wKE+9qsd3nMt7S2Z3OolteLuBfvgKCrjwWcgdlsAcrdmHfH6
XVnRfGJ7u3HMX+Zz6sK95Y/gSvP1alRXh9Znh7bZjgBwr8TxJ1JZTiBlP0FpQ4RsAs7NuJeqZ17p
0QxK4Lwc3AwCJyH3nUMdm9ZOoL2Nu9ohkDoCrUB8KfAjZ8pUn6VIQju8p9fY6UzU0IWKUcvw79RJ
apLYk3ixiiLAhJjdjvz8q3W3P8nfTzaG1P8nL9DrAT4+W7bJngMFBJLudkC+Az2Uhv3fEGt7Nxdp
5fkMtHHVguim3ZGIHHd86SxIpJ7EpE45eBuIbA+MR9emMC7wbdwPJfnF4xNOuXEFvreXSYH460zH
nrclvfu4eozlT/DRCMxIBu6ECfrg1K0McaNad9j56DpZ+DhTFqbnOOjl5tdmWN8FNWO+pVEyNqqP
6akZN5WjaC7oexOyQaZN0QbXpQQ10WxTfDUTHPVGHgCCZuYRO+HetK0AJy3/+oSLN2uI4fpvsgpB
EIhhinZg7leqKPJ27mPeF4sYgT/jyRk85n4YCZWlMqLtS3GMciUsJrj4d/5ImaMKCWD8Thb5ZjEu
BfDBOzau5tcAP5b2tfaWJsVZn0U+ufNJsUDkHbWkVZJQxR5RkZhLuTMt470i572xa3O1G+gs5ev5
p9z7QS5ldzilAHiqgygZmTphzO6Fub0NE2Tpnb+I3PF6MRwuN/wc9PcBS+P40561olKz5cMDv3Z7
PNMRd85yHVNkAsxhx0OIF4s8Q9+CsRRXB0F3/cdJquJSc2qKStxGbwekkOEYbDRgSWBI5D6qG6Wj
8cOIH3oPSxyfQYPRztuzADMYZkoYEn5V3GOuphD3gsgXt0FzTMp1kc+IjlCqGWjBmruq/A6Ov4va
f2qpwPNyFw9sRL4ozTevcrFmCyMt1KU1LuUrF8W8+251XtWLq3JOJ3HKgmHwCQ2yYxiTxQlwCMaV
vuT/XrYo79x5ikAwFYAdAMMegDTvx/boFEM+l5EFUUoyp994CioKEqALdEmQiwBDi51UU2C1LmWx
GD4i1Vu9yFzo6REGHXW5W9LUKAntFJPKp0mpe4vpRtVAoXbGq5ii4YHh9M12y58GI9pKJckVm4gH
pXwbyQW2ouqyyd0CtpdoqjGgSexSXJoSCaWWRGubgftGbDraAvhaMUzT7TAAcV1qWDcznrjaj/pW
/oW8TwC6Pvn3eoFuFnuxjJa9EtRQHfGMrigOjaOTgdCvpkhI2LMNAYOBdJduuDU4Us5dpL/qk3AF
8wVg+Jh1HlYWMRob/IZyHpMpaJh+4r8BO/RamPRSTDnTQj7SIjOBnL+x13WzE5coqKvc677mFvf2
GgZr5AdJsStmcX0tr3oHa7S8hWxJ/CCSOILwxNPrtjPHZNn5T0Q61PtGjYJFiMOW2v/gAUTfbj68
qGfhlGYujNsp0maZ9m2kvuUo54ZBm7GdkgGvlYWCZzBbFNPbq4BXcJJFseuncLIx6iSnGD8/opT7
Bs7XWZkMtIjDJnN6C/dvpLN71nuzHrseBN2hcHG2Nohg/IeLiUK5P0JERE4RAMP4Brhq1fxhCtr4
wZC2Ocw0onOBpI2y7spLFhmRpTZPtzVJklrQ6Z59jyGqfdkKow/s2hRfNO5/16xl3ZmZDZNcNswd
RDC7pp9KtLPjmrPJ7u9Txf0v2W5CBWtC+i9BKLedsi1ANvYUeHFrCq+0pDZ4+1tW5ucmz0Wju6ra
SrbcpobjqoY9C5cGC17P0wLUiz9qt6dnJCdIDuVxDNdvcRrBHHQGvaP9npRbpn2G45qGItWLgfR8
EwK/kNeBYTHhEVXr7sDXk3l9SWFxUUxFjCjawdU30xcBsmNy3pe5BrWYR3/NMloESuQ6pD1A05AW
kex3bn2pGM2aVJF2aJ5Looq2OVLySeBX1+7KIj04ns29Kode3XwOfU3Cm4DAPwuYMvESCnK+Vav7
e7447Yrs6vbDazInPUKBZVwEavWHcuAZmMkvcMfgtM+jpUSRqdYEKugvOYr1ehBsdCtqV1YIy8Gu
iBXnnDjftiTTZpgU5Kjf9GVVASXTdQaGh80NNnE422C6Kp4FOTsv07bVn1yjSJt/8ihpcmNu2Gq6
5lY+EeTssTDVLoZJv/crh1k1FSoc0XhmTii4twXZcIHezIrIJ1rdVWQoK9cxc84JhsXot9x05CZD
ZoEAVSAEX4lmsUXKxIyiyYXRVsGEbyi+UQQHzDNMvX8wQf3430QnpYhOIGxzWEMaLxq/070AyDx6
VA/IvpXNVBt96Z5GvZmPe4264drtIMGfuIXVGHW2Ky+Yf0YoxfPtQNHdoF2T2dYPmWvAAhQWn+vu
SWU8WnI9rJn5zaZ983YEwbduZR5VO+ydAZuznUa+YFrmg6KUVtcY1DycJo/XSk+6QDer82iPLgxj
wyDUorunZR4d28hWJVIGdoVBEc7PMBYjEqx8QXmAzfTv4MPlzNFwuFCXsulgxbnvq16N7BDJFLA0
wDj1spR/FLKYFfc0pCy4PUBwq05Nbk54YxmD8Zik34LM0SHYlPHL+oiE3KdMg45dIx7RrjtfR1rd
Ob+YIwz3r4fiJW+TE8Md3neRpVgrJguLam/uQx/UhUj7xrnuoFwWQApPSYjHacexdcwbMdO/hZ0T
+A5QaqvTM+/R49dKw0fJQ8MAI/XOM/o+9iZGIVDHiIHavTGCF8br+4sPtX33aaw5MXNq3kNd8BXA
1Ut6QDsjnge3REFiPI8k9fDwBJq4Ro1Y7ANweBb0ugqvN+HuDO63LeKabO4n0edVq0LzSeKNua/6
VSeiZiG7KYhKyTR2CWf8Rd5fFMtQsuJCSnl9ht898KRlB1FUc8xaXuJSJZFCM71TkTSK60wyB1yG
z0tasKwbIhhseDuTzq77IGzBsx494j0NH0lDKoJjUdtXOPOp7dlVan1P+OTYVvFJAxcC/aQqCU24
dX3QRh9JH5Y1OnzDHFNch1W3wBQ2UmTAzPh+CADu/FFuz+agU+/TGEGax9CIFL7wC55Z1lk4kOVA
GOKzN5b0LVgz4CvUCMdoTXxIvpg8fs91LQvPkYTfOJcFIY7DMKUxGUwQKAaNY0ghUmXzv9qglPVg
yJEawlJ1kPq4kYe27tEHPqJNta9K68g+V3TMG5QaDAx3txNH26G63kIo4x4dat8WEjOmbBYpNY77
GTqBNE+C8ZYfsxvN56+f+8QjB6t2nKOmZrx/E7oqt/GDj9nED+XGzSIySn/UKCKZAcPO5Dh/w9IY
3rGRFJ3uKVVG6s/INCUvmr+X1iNFEVvERgvYG8hOPnaSYiTYwbfrliRQCIibdEtUIcUJoPtCjyTR
vOhuaPLcviYp/xRWLt3NINj2h6HRgWQJvdOK4Ry+MX+Zy3vB+BoflD9SZAfGDANipLaa6sTlPsqH
STHNysSgQztD2mAl2VlFeVYLRzUm+Q1a0pO2LgSTjcejSQ1sySUilytIlsvYxqeU2C9qwNWHc2Sa
jMZH8AFt4mEGtwMmVDYK30VS7nB9TqwyLvX+883ytocYNRE4WH7cso5W8+rRSNPkWbAzNs0dew3Y
ctN2PcFKIpWNC6pRxtLjnc/KFQ570ERg9q6H+Vqsb6rnKBnkIDz51bdf/KA6051Rol7l80JnWNo3
gEZ51zUqErxuyivsuez+vCiLhhnnNSRl5cdXL4Oke6DpJ86+nw7B3iKEieAS4TMvqv2Hw9iokM8N
0PXO+Py5MXHkAPPRzcEdlHvi4uNDNUk8NzuvFjPCAYknHbE3qy81e7hbxNCCXevdCrEUCBx7vc42
T8gCA7MNdjKw6wHeVMJV1PsRtXLeVKqtEC6FaAdSp7w1RjbfV/zTAwBl0wLLJVU963A1/tBpKfcN
8VItcESDItuPgDmlpRs/ZNq+VvGW5LKKp+N6UkQlZsakm589Z9BlTniA/2kl8W7KaDquk7h1LCPz
lSZlBZSnry84mWBe4RZmbCeXyJVYjSorLWnf+ncar8+grjySJev9UnmFQ7rsfXiuh6Di/528zvz+
2PjJp/eW+qoQi0WryW+Nin7ysUoPPgWFMyVb/AYBFRFQXZLtD5DUagxDIqvUOueCznelgkyt8qIM
PxgShplqtLqUnGnTybEAxrU6YOaw+4GPXvQZT5PcVCqXVIdsbKR/wf86Xfq8oqfzQr4n8sYrPsaC
m1JZsJqCGjdwwy8vrKhI0fP9CSbK51iFeYJgAm0VloepHBwHKDxEIJYiISPz43DztaxDdd0cOuhS
ZYwZ6m7E9gMxqr8VXaG8QzHLnWmMNkQJ8CzOAfRTviilvVUxCUjQ2hdS+1rXA4889r127hgGygIF
3pb8XnNU44gleW+rYCIYwCsXOZ9g3cqqPJjHHrov92BP9s+vLwG3pGoH0G0YYY/i/CKpofN+lluT
+2vbt0WeADMVxO3DdTWATClS9zTH5u3s8KQai8bJjARsWNEnRLrY4Ubkjx1S631gffYB1+K/YWIl
OYGJKBVN1O2MorKvxnTWT8icna7SVxjhVPwIaGqxY5x3nR8F2b+ISI9TIUmHOhw2SLkIu0/t+/OK
GF9+5mnr1F4yVIF6SsEIx/c5ofC0zztEX/RwPaOVlMJIMMTE85FYE0Zvs559O86LVpkbEhEEOYek
g8G5OWB3cYAoq30IyUpqZDATbAFc17M4ozDpHGP0hR5NuiRDGztQRMMp8A2FFQ9iyXqwak/AxdRq
vvQQ53eA3UKYHYiJ3yy5G1PZ4vbQES2T+4mmkoKRPRSz9dkcpPkUnlOaKAfjn2knxVpEHTaBr+lZ
oAv8wT3ODoxcv1AxhhhIzXi1ClmNaP28c5iFSsiO0WAbCY7kpj5QPHckqjtdmgUllN7x6D+qR68N
WwaJmgm3b94XRrUJybmWlft/29nN9mM9aHih5kCOFSHVSWQj/TClP3pPFvK1HkDge9EHFDNFrat4
k71FHNu5MzsWmC+oGnf0f62sGFT/ABklwlFTGdOyCvzla+QU2pEJxa6Yo9AWTXfevC8Pl0S9Durf
FLKNwlrv+IiAeLLecgz9yo5GS69WFwM7/oO7FE/7frP2GFNXfTqHIMq6xvnsomCxIDlB8BSPSt/Y
nj70UIQc85m4Mc2ViYGkSvu/jyll0bYVGi1AkmRIQZZyyLprzA3h1E5Rvsui5LGW+IblTm0hgFCd
Qqx1dXGCyTAuZetohnekoeJ77BXv596Exwb+KEoBFWuwVrdFsHwL1L91ppCZt2Scj6NzGpECcmKa
ieKXqr0xbyxMk6GPV6aOkY5fBrylC6Z6RToitsKHRUtCQrAKZV88k0mWrF0y9mq1wGoghSiEi7Uu
KmRBgAzUhUf6n+cJrWhahiI9vWvSrWgKhW60FUmUp+DqJIDt4nRta3qAFYrHk9GfaEiUK1dxmVch
hQ4SkMT6Q/zCjqcfMVP7A9aiYi0tYriLykIrOq4aXjw0DtSgokmP8wZSduc/DoftdguYZRAd9Jbg
p3sfbbPdDkQ0r97H/lrW85AEV/yAymtpd7Co/ZP17PNseOouoH2YpG5peZvn4sbFUvl7v32FhTyA
y0v7o4mWyWKv73cnofA72DE9+ktp4dgjAwk0dW7pCw51Cf/7z0DcN0MYjiZyD+n1SoziuTPcSbrA
CGYsnb8xE//jtTHNUQweh0kDwC0zDTrgzqYuHeTGbUIAaVIoEA006FLiRQNeaYuMi5usaGRZ1Fw6
6GmUF8NplO2AjJS8bxprN09qLCmnCxdkl0Zb7Rxqyptv1k3+bA4UUJx9lofyrgWQWr2SBgrVaWsr
OhW5ejdyYh2HW+zLyY3kYH3NT1Q01OZWBoRZbFgHpbKnk6wkeGHstXw05nHd4o52dlyGJY2EuI0L
/8OOf/j/C5YH2gDG2iG0ofR3pagYFLwLvRsjJ+j3TOLdnCPkKzEPx/Pr46guanhU/E/jnEkVpk4F
LpI6WhxwSU+Mi93scgfWoPa47X0CbHKDA/+Z2rKZcODZlbw7UH1sVi6hKODWf/rcyLkygnELAvCI
DqpDfzsz9c347nFaWAZjXvN92M7pltPssAGqipcy9B2Wp2UwbMaVJzfQgNaMgStvjjnCTo3LO1GY
qofby5xWzHolerVHdhVctonlYGibibgwL71KXOqWgMisFtPnPuNpV9rxVA4Ndw/ShkomwcHu/A3H
oVB0enRBa14vKA9QtJ+rEX4FdSjcEPYaw001M92tsxlBCE2EFbXacBazF89p52FDzKdWwT/rBa8H
VEP+eX1Y2HioSddEygQiBbA/ZnJ6YR2zwdKwuljlZ1B1KvCq44BEZEtjsi9byhEFZ3FWtFE87crD
JGTgrBOeXXn0wo4vxjRTsSzYEMNiyEM2HsGaa2/hPMI3Fy8pLFk/S0kZDZ5G7eBGlJiGlTghUG2B
O3+lQ06BRlsAYKhLBzTyjPO2a5gTPbFgVmuAsOIpmWIfJzMKTAyH9zOeS9AE7636Dgef5OFrB3U4
4RxxsEVhKhtDJfCYB1LbDJjGMOTzZUWgz6+SxGJyROi85YjGrxApNUtbnl/GjOE0PACOszh1kAY7
mEMBwRnb7zksZl2T9WUS8CxB8+DhsQgC5SmHfBiiOSiVV76zfp29nSCUdGE/B3LC9PpLw8FqYj9x
5uZlsUhDc8RFpzQ0w4jhaXvaP04KupcSUwWNInnEVexaLH5bb78yI0MuPz6sX0Jfh0nYjJ6fSBkD
gOnqFcMu531CViup/NOw2K2N3aOLHBj5abgQPD6hAj0r2PpiLbWZQ18P1LH7t5Vdj5hp4Q3OEG+G
OCHMyKR8WGJVndsdmoT0I1J59+EEmj9Ky++7h0Y9uqVx5MWQBrxmqDmZqymXUbqHGJpkwEdn5GPQ
NzRpoetr0wrKpsigMgXSn6LGhXJwX4x7FW6Do7Fm1aXnwbymbfMCitpcEcYLRmmikA7m8em21JYe
6evGucVgS2SWqUmbFUSfOpl5m33bq3OG2nWS1Ot/yYloPFpuLh/C+Ieek2mV7GwRT6syOt8snHBE
N+nNS1BnUgGEkAigQim47RSNm0j+1Amb+Jl4adQqqM1288HZ6RjF4P8FkK9LoOih4/RmPA5aYwcO
KIW0mSOl+sLa3+FOyHRQpVtNtromd2IOojQDCXSaa5n2BGdm13boNcAK4rNp4C9kIPTFGmxWBjKt
xSNLZ35fU4Xum2nm0DdBq9Xn10/wxe5nJDq6+TWlEYHAHwhX+5qCYFNqCn3GOKU+oEa4+uB0cV1O
Mtd+5l7huu9TUNKaiXz1GP8m/CjLAFjv3nfnOoLbNmeIxNqi87f+YZbMAec4Ka/nMjPUefm9Ij9O
XVQ8x5hpQ6BK3lbCFtrVrsXinm/cNR6/diVGSwEPp2KOr+xT1MFJ+1VbOTRxCvZtEDToHtm+DdQY
1KoopYwMZlrLD2kDiXYbDvUOvXJh4vBziQEs6Rp8gZ0XT7lEvhDVjR6k/yg9dmvVvGz0G+t3ZTZn
ewOPdcnkGEmbv6n1VB+KIDE00yYY9oTiqNKk8yIf01CsKLZ4QiOISZBbr/9kl8bmEWEoNAXBpakb
XtY61CLqQ0wdiyB4xp0RI9vOueIbUHIy6J5lhu50bZ2hr+tucQ3A0+4VYw/nhf6Ufp8Prfum4rvp
PdETVYS1EI8v8g89Z9hMVeNpRLO+yNBfHp6ENuDsl7pYn0XRA4YfJz35FnYqGxUqrjS0nDkdEqRf
8DMa6EZF7iK7uwRlfiYU0wx7sgEanLAYazMsOkrBNdrXC+MTwuSzdyZpDIk30nwJJhV5ETfK1E3a
4S2PPKHGHLS5RKkqhLLO83t0srq7UvVmje+A76Ov3oaQcBXF3N+M6frN9sG9c7veHlualzYwhLpJ
IthnJdXZmktjqynytaDBc1AyfKasBhmN2bbNRE8vASqFJjPlWaIeYDwMFOZHndkfEXCkJ7Y/WcrM
v8yUb0jARhvDoCds3emV/7DQ5y/Jf73c0Uy8EzZpHo6URURS/kJ3z5akQz54vgadNQTXB+ndAUp9
uJ6i/4h0lgTVDCl+qxXBeV/Mn8y4J7504Yv8DGzTCKsiNlE7UdSj/erjmjxRoBBiZUpUpqg3N9xu
CXYtX21AIbWEJOLJd5rt1h10oRiZcDvU5Bvp28PPQWCGvC9EBIQW5RwWrV8jmAojHZzdmSwwooWw
fRFeGlmjD8dtMV05Q3+NhHrNFW2oP2y8R9LqLTZJX/esAg+1xsF24L+qDU2QR2WlfL1ASHWLK14J
wweHG5K6L4znWXvOPsx+OJDA4MiSWc2f4O5KN5Z2cqwLwcw9DLd0zrmC7Ngu0Y4oaiGC+E3bbaIu
C9biLxbJ7iAWRSzkBdn5wbC3YZ8CR0E2keLkPQh+zjR8sJdbFXJ5zV5IbdchqX5sCTSAfJh5qx2z
0SkA/4c7+ZuW4gfpEYhJEIGW5WU9c1CG29VWpa6P5IvqutEHLgT76iDBW3OuKkISHJdJR2hHueXK
witzkrMpuE74tO6dNzB4qlUgk0N4TFG4w0Uidb1xwxc2nqqVBtg9FyHGlGTY1pHNz95q+7HoC2bL
Ij2ew2MGMRroWmsKMM4d9ULwmofKpeC/1OWwW9jmBoJKQgYR0E5BAZq9//kFRfcri13rhuVloOHe
JjNYmZPzuk+46kKwYWu4a5my7vnEZasSLqAD872/tn/WwuH7WchUb05RtCu9XS5EOg/fvGxR2j+9
FVkCKZiYEZjC6xMU6Lfkm9knxvAnNyXFGSp05A8WQggKQA7C+DX8kExqKLU05dkDrIRgA5E+XaWs
U8S3WFs8t974v+zfkkLuu+4mi6EOIc5mpedTF+k+HeBjVcAS+Yq9AFGbcQfguRvIa6WKwdTlmZAB
OV0R+TtDO0aicklS+2BDv76H/jhOUyJ8DEZ7wEfICqPs0jLf/VptXuTuddf3thv+FiN+zz010ZzW
1KwDB0G+tkboE0A76wN3dB4Nv3N8lweW8igntWRTxrtTN+3c5jEPHFO2afr1vTzYpJFH6B38mSA1
8DsTWmrfcTUhr5eS6q60nAEiSodrVKV97aHtukcmoeLBLEmJzqtKUZUPOnaRG41hiKb4kEu6Jh7L
uFlneaw3AHGfTFGwvx89DkVEkY/HXnNEpJo/jMTjk1iZSu5jaDIqDxQykpoXWRRyXPKtR9aQ1gKu
hoJCgxV1Pk252fmRIRxVceezTe22Cp6lHaJ1S0+3hCuA1O6XrOqDnJ1j87d6W1XKFGxe2pRxoq15
pt8BkxyszwjUrXftA0DKKe9jHdsZnx5HYwII3ddkwPbHfGy6GJ+6VPSoVvS8D7I/yN5UmhJy5S0I
MBhv9rf19hS8UN41aV7AfM7BSpVvhoHwlYccAHazxWoV3Zx6AqSWE0jcZQPkDsR2AWcoCgZptZeb
fW6/7rYbnxKDjiYctBXHqZZz8osuxuth7YlWhvMZSOBlvaBJfpSBJOUzStu6oeGOskxwUJZhlQTo
FNId9CxkYTZnXXCCwr7oC99CRvrcZNRrqnFUyJio6+Nga4CTuscbxycLfrA220CxQUCbUM911VIz
8/G1SAJVGNgYMtmYrEcRdsCTvcSgCCq3hTGdGgJu7KGbFtcKUijk2qCul18Jrumj3e4w6ujPH0EN
SqKjECT8zF9UTPpj4tNRCjJ9e4hMEnu3EIbQEB/R1Fpi6uigvxe6g0f603BExAAnJWFRPbBdkpsc
NCVI1JkVmx3fp8M89gUttqgHFIzLlFhZaoPVEa9VFX+gozB09zovxW/9dpWYb8uj5WRi+rfkNOrY
uOslYdd0iJUte3YujhSDcl5qD+b9mosHLDrCWQ8EvlZqd4PaqpObCv5P+/a6SYPHW0ezctA75V8l
GEOutu0srNDXul2M+MVQUfDg0TOZgzjBTcxjomXhUs27V16zDA+SUjsRX8bxVs5mkNxAXkBTshAR
YqWcABrXLENpj1V9U66xLZxqpEkcaICiWydAgZA+v2Z/7RAd03pj/yMkot5QFOQyOnALbWw+VP+Z
+JVhVzMSaTIuSEThlpy3zthsXyGm/5npjJ59si8qBAXZaTUR414lM4md5gtsBBZBY6EQRXaGqqhe
VgI10s9+s2g3ZJ3ZIL8PYeddA/RLwaebZmHJfKoe8OvyJI8j06DqDobddVi80cGr/w6zEi4buoJw
pRgemSt6FvPu+CWzMWiYfP1PEayBG4MdHojIzW8aGBQsawZVa/DP6/DtKO/vvcOI+hr9Z/bm4V37
bO1XVFj8ceVV+J1tkhjnYb3KX9k1/OClKBlYFb16alsBIweiGISZkVWx1OMolCX6bpusUlmx/KJF
vemhW0dsl31c1+vCGlBgLUO6jZwB6T8sfClUOKJDoUgyiRjTeyQAlILc5F7smU6WvUcFRXpYPc/O
qG9hbJtMD1bCnpvIKtFJMAzTbsIowvMsTvIuIhjxF+FRp2WWB1A3TofixWQ5/HkLQFFKaCbdlOXw
QyjbgesgdvEUjJweWHQxbKetllZmzyAo0IXZpiz68mr4fi0NetwRfqTlGJKztj45fVkbeutvd0+7
mls3jd8X4gu4UocAAALWyYgLRiHqTqr9M7SWrVBRxkff1ebiZpznXaQeMn72LpNzc3NjBjpd0Y+x
5MDEZCbe+OffzmzEUSW2NS+lPh+FrlF1kIdN7EjU/foQGQz1g3/Ge52pGWOytwmmJtEdVcg4Sdbf
ZxsfZaftU7Lz7qOofAKtcc8chn3yx/PTONMwj22Zsh1xi/XvFKWb/g7XHU3uMF/YT88RTtyjKdNj
sKWsXoJOdLwqs3Fxk+OW5yMyNVr9eVXbts+MZCdp+OztyM/i299IfLSl0b97NEBWkH9AJ5o9MmTw
49XipiGcXVCpX/mNX7yhu+zpk1ncx6DRqFdhLUeS1gMF0KDoBovKAkutn+goQwOmhEHCy7etZym7
gqDPYENMV1XQ7loozIP8+b5jEH65LLg02Sg8SQGL8ECW9jsG7PW1d+L7WKcQSPknbANKFENiCDSW
AVXBuClq1num7fbFb2HZzE0aYJado53OgSvxrSqOT64hMMZYmF21MVQ+qST6Yf52EWM+DakLP9eD
IKxIo2KCNb2PINTFtUoC6uGdNv7chXcjS3/Mj+NIBdlg76Lxn3/7uBrnBy9A1WZeofzetOvhIVdf
Fa8kdrnOM3xz9uTLkVVg1atcVYKKR7biLYsmXecXP4ZQArxIjjEG1C5z37Ap/X6YlO5SoAZ6FnIm
XTbCv+SrjK8uKIoC/6hsTl9deLbsgTLn3u5U82g3gk3hMW/MVi0MATEWcrhmgf6pQDLAP+6J7sc6
1uZHnXkdwKne7EkMgzJUfn7fgdOae6+TUM8ImvkruvXN/OO9KKaoJaSpg70sBnwp39XSUfVXpJAq
lypdTxulVlZGk2OtKNrTf1dRy4NhLydJFt+YcTd2yYMnSyBfsiuRPQQdTG6i+1AU8RcL6ViLFJPv
kfyC1qV/TpFvnl+rbvWiKiALY17Wn9Mb549TQmkRl1X9aQ7NtJyYIRZhrHsj/9cAMXSuAth/EoWR
+5eGS9hEaV6JZCJH6LCynSu315QBahPvLC6SZqlJuBODuq62+x47WoiYorOcHvvcXEqhPFdQimHK
tibR0KuQPYlaRYkGPY4qdF3atrMJdqN7TEO046iXmknrA4JynTqdUxTCOVaQt6irTR0HpNs7iaka
mOinlVJQvvqhl+wtrUjIPrGceZmlfAa0HznFTDfc9wY6AnHf7N1M6CuhY1WJK0v0CVQnwAF/anMd
Q/WaGGV48EuusQMVN9jUuuAC2Siz2xJMaQzjmCcJKJ/zk8zhRTOh2bruubmt352jvvEF1KYLwafL
pp5GcZLIrnXsqThTDxIkmFxUBXY/08RhXFMG4l67pB2GIXLoFm57ARGLbOiAcFunx5iotq6JG7PI
kf0OJI3uMzQHQiZ86FP/pvKLu/bUpXqwr6A7LQyroFtaXMi0xym/O+rZaNrH/gAwmZxDRjMkPzWM
Vbj/jJx+LkeaKEHjX0Wup4aYu1JIwes+75ljxJ7kkorC8hX3/J6ISM18HDA7xCIONjVZamxl4oJM
nJrvmd3fieGR1/n3wGQz3DWnKlSb99x8gCyoa8KcCpcoGWmLwUHV7Gdocsm34aI7PcX5/0nbFXAV
AK6qx2B5ZSzCW15Zy21aH6gBrLgmrAEkh4Woc5fRZ0M/aTFzr047ncc7GgydscxPgqyswT7V5oVx
6zJ0zvEf6/vmpHiKdrg89ofiirLcrCyj7VNaPvhgKMBEEVqKIPq6QOemcObeUwHGgRvigQQ3e4mr
n6SgW85izdLFIlkMkblwZPtiHNpAzL2M7scSE74IiwkLtRqnrQVgeJQHHxlNgXwsKjnc9xpJwbrX
/0mTZKbGQQx7jjhbmGFJ1KXs+DR9sySy5HnAt0nnoNfRjTI3JRhNCt7Mq9OIr59Nn0VErYhJ4ES3
nkFRab4eULMfZxMi9NFOG4oCi5lPKFd9uck1ybDKhiLhe38QKBy7RbKmSVX1G1mpCaLgkrdDBLBq
RwJQyO+S1T5DOjUf6arFOJfv62Xp8Yc/zz1tPEAmJxlEHQ2SeybDB7AOzv/61W5rcXNClDu+1DB4
hyXvobclUkDEgnWqMg1+ImSUuE9X2s7Ce2rcO6R3wTyRbldN9/JmjoyireS6T2YcypyxVvCj8s8h
HhcgNVssz6/2B6QPBa0rzbh3UeYosFehJMdrOQV4xwoi2H7j2Tw1++tpPi+lt6Uxgom41Tvs79iS
xKG2o/XrP2D3ZtUmcfFBbCugAsIQ0WrsCWKicyzlmY9AbkpKXB3SbcHevFtwPaElgojquKV596Hb
AAnMZnn3OEznl4M+P3PqSN6pqGoNeYDm2Go69mDLJu53pxyuSNoSW2Cc8G4/ymJecaRqbPirQsZ7
XdT1lAZVoLIArdTCvIzfDyIffHogRyhTKfh0+1Zf5SPfaCEye6/CrNCy1/WhKTx1JPo36150YqDY
YR0ovx1nIW9oul3u24wXIDCU90C9VQjX6E+tALIlpl8tHWMMFi33qvNWnkiZ7b/0/JLaTufrw8G/
PtnkadmYD/fcVym28t8ImV8m71WnHuCt0baLgkPswC3qosfkQZJ15pZg4bgD73gtViFaWvQ+aMbM
+t8xd8tu9VQH7QmF63obBNEkgEp0FBesG0qkeSd3fcDITLr1t53qY7qx4yDIE7pSRFVQ0C6XohVh
FoEvLJVcGEL0zrA9jO9ob7y3UhwxTUFV+lQRKC8QYlB+h8A5/S6WCkQXDxa7CkO0dFXAKsef8A4R
f28FmbvE1G+cSTrNOKyOvtLsD7u3HtifX5Z3Yemn0LqEYsVORNAJdEihRNb1MNFpgZF5BiujZor1
Bsksm5pWGds2G5TM32tEs+6PbWJYIV3OFfL4E/xD7DFDzgbkzlqGX3Pw2Tw4m3H7rY/xpqd2rRP8
nHHWFVdP/+3xyt88PWzywhuvcdRxH1vuG/2wfgc/4ghidbcCcuohQuFxVXSRq6V32WRZ5mFRV09A
Hb13L+O4ZcwZ4BGuzTjhZoGnjmnM+0KaJtW+9wxzp19pqb6HZSCb1WOZgQoyptUnlVn06oTt0497
fEZgK65Tgao/gccsO3mNIP58ELAriBgND2wiUIeaxJtlQ0vjjUINMyzP5723VjTuVas2fOBM8IJ/
Uk1Ekmu2NckNv/u9gWvWQWSySaaI6nL5y654MQdveLN+4n8znz32ldEH5DpyRYJxcXbb+bSAMTDm
wVtBiQiOmRnrVxFFpegwgh5xMqyjRwUfC1zPE17VwiYF1/KoiLNHTd67kMif6IVr5G2+sc0ZAD3K
SWX8oA7mY/fygg095lWRJ2I8e4b7qb0Ad4ywbpaPaEj+A6MuoTQbVftkPWyNxc146oC+OEC2cbQ3
92rLZEp9CT+VS5+6f1oEN6qwLVuwfq3low5p4YNQLaG02yW5aYTOAtiArvcUNn0PaXW4OoRRe52t
RqVV2HtpiWVPOjjW0QoJlhf2A+iEOgMHkkkzrtKbMiyzdvRE10d6vHXL4mEpFaoEFSjrqsrRVa1L
4Dz7RYadyjam5ng79DJfFq4HfUtCJMZ7gzj5skGnqSlF9eoGk1S3Vvl3vhp2XGkqgO2jtBiWnS9h
Ln6czfhmUCd7tXlhswDq3mwXd/gVMFMSjCWsTHxepq8HlgfP6xMRdlqjxEP8fIl/qmGCwQONWE3W
7v9zql2Q36yILAYzTTDdOZNPBE0w0NzGdXgT1OYdwgrJEA9lNBqTheh5F+/TP21KtYtU6qV4a/MN
2IEgHl0ijgnyUpbQoG/Ci4/UHdDeLEMwrPSBLn0tGW2JHIRkQBaIEf73GIoRYVOzZb7I7oP/+AFA
pxRLAYL+ZrSqVhGBw3kHXymwsOeZrYgwefcuGWr5Sog8g3uEkNd43sHboE8uwyo4Kj+wmCVpTd/t
BKvVz+EFaquKf+BA2MSSPvSGvxNiHNXW9zUpyU/alcS3alEiKc4v8bL62YuYD1Goo65aD3M8WqZb
fc6SkdESCDPavGZzPJeZnc90b+enCO83iAkRxtbTV8YscHe33mt4JaEGOVSgHRMcr4xYQn4Hh1rF
Hrq80dXs/mU7F49Y3wgVDaF4BDbXu042AmR3kSH7qOd3H+cg8Bl/KVy++5mQv5KPdPcacdLQscMj
KugEBbQvwA0H3mw/oY/cniinGe/v5MwEFmmopVdokSaNtq4ZS6yGz2LXNVNBjShiguHfR16uH0ei
6KmAV3kABxHu/TgZkaqTr9TGhcQmhMUOa9BkTv3iCOYJF7eabsUBOqqLfUo3z+huc5Sw9MXR9zJy
yZr3VgQFgR9so/EFu8HceaA53z3dmOV0W3bYh3CPUW65bz1TV7/0oHLYmkuqOk+fRnFbpnwEiGFR
aQ146Ya/Zw1kwR7xXGM3zF7DjNKG6VAenVoT8HN+RDb4bRIJPEWAyb9+gDi5qKFCLfJ3fcDqX5jk
le0NYnEeTByqG3m6+lzO9vbYuYTiZC9jlobJeeLZlb6z8b6nOPmkvDSGHg5oNfv+zv7fAZVBnKxA
N9rVTVuIrL2ZjrCvDrH4aRUAPQwtugkWKmvYcSIZixjryqG5riQp1FRVPGpzFfiT8Jxq8EeqwR3k
SIMfNj8/dsNuWdF8RWCsTXv9/Gv0dvMUARk8tq6K1UTZRp9B7mUWL9wkbCzDfDnWeONpS3LByCoC
MDTVrPV06fOdfr/cLVObSIDmaD/QujYdcQMzyPj35ij0BazBqfdX3TN3O5TIEnbrlUrk2stThWon
1RUZ71zIZqkptHPr+qA5hXQ1qx0ZqPvefe2VGFTbcWWkeIC8xMgl9uSMbfZF393xGWDjJwSEi2D1
SHPSvcawtw3WfY5fUyV5GYEkHwAVcgMvIrBRFiXj+D2PtX7YN0mBIu4w7htrICRznRwAQbplflNg
pzBMBTj7lm7I72/hPPKgsZLFKWvKCxU/5LXL5uGzB62P5+fCJ0NiRTO0ouZBfWHaoVeIIBf+4sBZ
woRxb/5HbWc7An458bHcziQ6ii8Vb8jc67VrBluIoWDXnahUp4jM06OqgOzYIQodb3IY8NlUXO3X
jxIxQqqaw0erx3T6UulW32ZnLrFDSdlOL8VC3wCEaaD8jr81yu2iQnRZC6jJz3N3cqEi8eR5cslD
YQuymIbuDwuKCr0MZrE7r5jGm8BazZiI4sVhTcTDIi6tj4MP2lpIskmUi8OupbqROU17fkE8aATm
aWJvxOqUu3qBvZ82yJQSzvp8Pxit4fPsCd2fjEw2OPCvpioyyBd8u2TMCIYQMIDiIhKjX7c4tiSl
znV5KHC+yim1Rz8G88Np1YgCFFTSVh41db5uQ34cWrrBDEjuuqxrvysef0zjEP1Un29UwgzmZd7+
gk/QeXQT8sYDdOXC5WT9iENrDfJwAu54pEaQ8kt9NH89s24/vCTlC50ttPZMb0/1NLPF+O8Ucomm
0R67kal41jCxhSwswg8oDWfWeQcYeWAfcekIHJKCCE3/W5wPpMnJqSv89lpnbX2BC75tyv5BERTM
5Y8KZEC8tFJAoXJ2nco2OpvtczM/+wWYE9cTpdH8NClBTWQyAy3SGQ59z1E+sgWzgDhmklA08oE2
3kfRO5USO8H9CHzmblfV36ro6kwaB+nQR37jDJvtTtw+T0iWQxCan5lirWQ3plXDRF7ZXiXyIIIE
ypvG+bOTsCRQYZKlmck5l4eCCKL31BcLGfiCdhFalBLuYibMqGf1qjs8n45z+ST4aPtpXCPPxwHL
hqnQMVU2MTybfNg0cp3Xq/tZa7xN44IIHxpk7+PF9TSS9ZrraOi+odCvmPGQ8eNRNNqo2AKvbNmT
F247cP30wKYYl2eLs1s7RGg0PerZI3mvvT03v2Qzatqlc0xPw4SD/6bC7hK64F9G7IEtp+7QfIdy
Rs85E5kEVqCw/IXJ+0VoTl48DW34X4TC2QaIPepQDafesVz8JRI3FN4oncKl1n1L32wPNkumIAi1
bG/Q+g4ePOiq78yXBBQW/mANoveuwSWcv7v78rKi4z5svKxMwwrRjv5Eg0EJL2qBfyWoJW58lzVi
7W65znvb2tjc9ZyiL44H5fhlniEK8Co+vITRqGThum1tMxAwaNNIVqxs8jOvVHp8Gts0zvv8CyA7
uAXbUhH2CEH9G82YqfVux7jMd7ByXCEB+hGnJh2pbg0VAJr90hp5uOBfMCLl8Ioh2UHck2ddpfde
O3L6lp5ILBYtTvDWRaNGS/s4s/3AzPteUK7aE+Q/SENRYdaE6A5oBguOSVwbuET0j5WzOIwLJD/m
4eGTNR0t2RGz3waGhauHd8xw1d2iRb++wObJ6sI0Y7/hhp+YqnPRswJ7STR/6GT6iTi57CxTpXAr
OzmFLPYLgtvSFG6AT3bAoScHNul+1LHyV0Ke6AVE5sufDqknAkKNo9+iGNaEhg06CwjNbvQXHTvh
f/Lk3Z7xdhuexQUgZBsfVl+7h1f1Xw/IdOrN2oMO+2IT4SA6yslxW3GZTjtNj8jPremIMjjvApPy
+U/CCpA1zBU/3IP1aOecB5RTge1BXKUseWTegblCl7TOJnv6zFccz1UiMKa7hFiW0j6MFZJvRrgW
W5oOc/0TZqKJErIoTYykuc3uIaGZfzS6IHff1SQMQeECeY67DC+xqbDbmAKcd66FGl7FCyNACNGD
tXiogYuJPsTUglJZ6Dm7uyOcuMLoI/oMf8Nr/UxxxOzzHWIOiBBOuMQwjgQ82z6X+74zHiV90R39
PJXpxKFcobLvOA1oBJvyNkspzhDwDxraFNyxy2qIHIySr+nneZwa9fjRQA88bvcbEo5auKKeq8q/
FkDXW4UW8Yun5V5pmZyLyDxLxvCI2qKpiDckRCxwIhLJG7eQAaZSnhq7ic1zrY+LGQK/zmerm954
ZoN0PcAN03Eodg3AKsZa6oSaN2UzkJex7+kuVnwrS/5Pa9OcNETMNrM7lrBTnfvQWKhUTYBVW03S
Soo5q9KrzNX5Fz/cRC1VuDWu4uBjYxIY9hg0oG/Csda+/WmRYZRNa47K84I+SY9eifBdivBVhCFb
i6t3FpLU6OsnkEEWItgyKOq5xo35LIpZKKyNpcJEs4bEmx+2b6+IMOr88Kwhy0WUZSxQy6Pip5Su
BJs44NmogrHtqhN6Gkk4/f0Hp6IR4ANbKCOmlNoiDOE4Lqi2eikR/MiOcqKI1vKYD0FnfGh1NJbc
EY6v4lXcMeMXoQdC7DkHImd8T2K/zYpGC7whhlIF3p//BD40LGra/FSppNwaEUaqk0vgAU9YSBuE
dWbm72c7TQ+0ruPuWU20VSHfchulwC2/4NnG5rVTfIQ0GuiNgwbrRrPrOj1llVQi8gyMEcMikwPL
/VhBGcYSpaXeIUFtmzldT6TI9Wkr7dyi6+NarkucIJmVyV1ZC4dEGxOmd/ANp0Cjc5zT+c8Bi85N
xHrG6fyePeLCK9FBen2B+2KyAn/e1OG2KL3zy5tbkwZSIO+qnKrHCmtXkkc+g+MKPnqcna/kBCvD
8zmk/c+I3cZKT1aMWi6UPU3awHEnweFC1g10YaUJTHlpcG7h/txKKbHzDj+1VP0aVBaph1uJTCDA
LpWYlx/wkbtsiQJjsmihR3t6rBWQ8TIfcfwGWjSqs9IeBYNaIceAFPieQLhuoY8WIo+TjjAHuO3T
1ShOYqy50bLSSrpSyinz7FKr4fxlTnWfVxJKavJwgePAFfUtS62wf19/hUFK2SNkcF+fa8RVSSql
iU1GXUQm2QknNFyjsz5EjjLwjgz8mBKme363wwmvicZyZubeMKjjhIzJ9WaqLbhtN6Q2ol98XDB3
i7nKHPqFwNIma0CUqhbMeSBQJX015V1L5R9qdxXtiWMpCYNVu52fzCwVrBImGJOLE3qU3QSk1wR3
uZPQf159NNqHUuoZf4+t+d1V9hTZySaRh2gUkOoc/tc7F/jjTl9tulYrMMYFbtQR4bYHaBYa/oWb
GBPuJKxixDyAhqC3ruqb5nXSU53b/NgUucR/CP2pS5zceP39/tgLmPU2jtnKcIdikWwMIVlaf/dm
kgkxB65Diw+k6kM1e7aktTQ7HfEB0jqVBdN6CAgis4gD/BgbrfRNgsZyp3RAWkzpJGVexUOKaB42
gdZeAlA7QyZNCVMQb4yIi35U/0dzh1WMPsHPB7iE1PYD+TizRkTHC1JeXTODOjfrernC8CEgQV7G
ndi9PHRPrTJDUKx3/Si4Y8ZLQjGpX0pnrNt7f7KfY317X3JZ05d2d3N4+Yc2wLYSzj/KoGd8yPM9
4NlIslb/jJua4Vc+PCDDEF6ExduexB2v3AY0su23E2GU9qesMq1aTi1T8MjZAzRWxF5dI6wmOy+c
Sex+3i7GIHOW4W+cHT4SY9uwJqECACuIWjxI4fOBs2vslQbRFmUMlLaQJ5mDKj9Q57t/+QXkdS7v
dPIPS31u/23k4+9B/s2EznQeLfOFi+W7b69BjD5g3cClhpsx2Dwk/8KZy1nRC0M/8q/PN2Tt952l
JZPOKpA+iENfswvR7yQMa6Tr2VOsZgq3GkgUj49lb3SK8g0EKMvqy0M1kyAkGonyQYPfxOuuGuTG
BsQ/clczu9XDii8hKk/AIlqO+EVIg/qWKlDWaCXsNYVJOUGkDuG2nx3Xt1hwlC8P36Rtfen+4zNh
qdVSEKzSh+uBYKQ35qdZMFs15CXvRS50+WcmMvBUg8ocW7tCdDi75WS2gErdORpcJu6gs9VqLPv1
LAuulIds+1TrkL4+UVKfQAY8sp6/OvqY3CwB9yCXH26jk4Yydxu9bCBJnbYh3slml7/PzWu9P20S
VuTZY0EMJdX7Sx4/njQfuGC6yXuWw7fcz91lA0uySiM+7swTX0G0ug7EuBY7kiqhhfBLh8758J4d
TvN9TI1pCU2OuYCtMJGTz6ZiTkCqtLrvdmjqB7gnIwq+VJtfM80TWCGvpW4tMeAo2POjgxYLe3BP
7548pHZEJCfOF2W0e+TK08zvDZ42sS1340bHJiGS62ydxBL+iTfWvx7MYSchDysY0pdVHdkHKXAJ
VMTuoWmyMCBij8+VJe/uRA/EoUkRcAuS1Xd5PS0MCnxYhSuFKACnmJ0Eo9k33cC5kx+r5cOzeHRb
0xWjTcgZOPzyDp6BaRsq0b4qfUKbSlO2iVC5S/wNaLtLY7ajxQB6cs25YHTriJnaqpus5NvPdc6b
s4jyTeibhymTsu+nI+u9ioZhj9qLJR0AaR3rGJkIa+S1MeOg2wKUiILBORA7ZdaDizriqcG4C+xo
S9XGPxJKxMUJYESxsQvlP8ObGhwsSLxllWDhck5R6TiPKbk4FUTYCWX9HmBm5Qz86mrvLzQipRQo
3JLLZ0e7NBk7geK3vBXWTVYbOU2BFb/IoayUpU8Mr3Yu1kYcssyYbS8zISarZHdLhZwgGtXK+6td
lDQl0g78SG6KntUMpYLwTPed6lcHeadTIals0SqeMMtlZZc0jKRTQnuDhG1x8qTVvsm+1O4fNr02
5rZ4/n1kXn2Wbkm0NGGS7Ym7N+lyGHIsrqC1koWvqlPKQXG1ji4EN8bX6siIvXn+ixWsrxPMq2QF
YUPsk9dyBV+5mRKT0fQ1SS4CA+vWNNBGwmt3UL9W7Jf4b4Q//QYBlj+ik37dFOLJz47s1qWc3LfW
0FKzLyMpJmbqIcDmuBbRPO7zEOeA9yYPvO2S9RJ47zQFvUS1gVNtaK88V3MThjOlGubKTDVhYMFO
7p/rkjCoxYBHQdWFmpmK3SnpGnVvf8eHwTlEhBiwdJAH51DtnEd69Tf2vD8hzxaLEp82AOAjYAjk
Us+UsTwL8CIv2lkROeITgCvyhESzJc6keZnIqoJzDw/lHR1kRzuCpy7wlhqk2L3mQ+35GWakbqTi
LVPgNn5ug8SzjOlPVEjssl+CpuI/J1Q3L6GWBrAL1iHP5xUiN0Hh6ITQ5x41g7Q3YhvKIwPH0s9/
8jJUEWpHjPK47D825vV/Pth9BdzMh480pjq0yUxxJpF5xUsTlnDOPlczwv1apH3+m882v6iDY2SF
8x2H4o3xBG0B0wsJqfT190XzDILbOWdeNCk16R1ENFEPqDk2niC/+clADp3/gYzGNKlUgRKsk0AD
HheXkQVOzqWGqPmxkBFTb0BHdncL4uEyxmhEdHQNxDDxQ8bdSbauXElsY11Ypb1TN2/fzhYNRvoR
ZaJ/5IIiMAxgTi+2/+NqbTJqtP8U3/nbGGtDyfZ5G4CfBEq4IJUnzuBv355h/Hq1/8zXtTMylRYe
3/8BjTnWXNAEyD+Sc0N1FIsfZ9W2Tj7xFNjiCxawYeHsA5oD/ZlM7f8DvymSzk+cT/6CVi2DYOjR
2ZfHvRW6grDiQxFotUdHpDodTYeonDOZxBCOlNNAi4EMSajGsyQqr4iDbIp6j5DpGRQhm9+knNaa
v+UMNN6F7UYVhIDiUDkQ7lmG1QyryowyjEGH7sagzQbzIT4eE0c5ufQNxsEjFS0+FkJq7cI6n0L2
RyMpM4HIwms3SB2EEHTDE+VfszLhCbYOswSu7w4r2GBoZmD6tXkDE3rC3Xwi6obWJnQk/p8CbvJI
0RIkTmUyAhwnEF4FQw4kF2u0QdVGdvbHjGt2SE24ZtiOhfdQRuBvP6mE06iaMJTMpbHIOpOZP+7b
EnqS/OgaEsRKlKU6ySkxMhscUtoIKy0HRCJJspwM/qdwZ9kM4ifbzl4IztKH1IDj4BTg5un/COsq
WrK9mIY83OBgDclrdjY2hpX8+jCqeo2ZqIGmZ2O5iMe0myiNb4RmJzfgyfrr6WGWucUYlo1c6Nqv
T9MMGDjppGm4BdD5IkE9jm9/Ud88mbz09bldBFklKmQBImDSp4AtuISSB+4eZEC2P4zyTSfM88sn
MBQmcmLDp0erScZnfEHAsLH5gTXdtxBwGRkCnkPIk9w5PqvuVS+y1CWGJdRJe5f9AAvTux6bgs5I
vXl83n9QKgJ2exPFnW7DcWJTT+f0rE8wuC4s+cVNJ1eU8oz2aLCeL+0jFXeaUSXUkbo0s98G6fmP
Ki4CUEdAgTJC3Q4uw8SJB8pRaKtyaLbzV1Jlu71XISJdtzcVNvqHVuw7tJM2cNwgTnHfoQkmkdLK
N1LkGn6UkooMhpnseBZdGvVCplAHaCsjBtla7m8B5+ZxfIeyc+N8Pp+cmQoG7HG8/JIXDbkGpLia
iabyAH3R17atCff47K7D3SVgZArogfW1rhhITx+g+WfWAr7tEFJTRY4CdqpimS3PoQEyOSlfJjgl
RiUf9/Aj0Mdyawex74YgdJDVLGOcybqo9LSAB9B9slQQF2xwhbiGH9vd6CpiIvuPp0wr3/VKYcFA
si0e7h4aJWdT3G3Y4051p5u1JcD8USfe8vshSH07oLvON3dEorLiKtYVCMKnCbeFr0tlWpEhzcA9
ADwRVCTjWH3Oj3DEq+m9ZP/ayhP4qWMN3eb5VLxMLmKWymPv2uPiSLMakHP65N0b2O02oWlwEPzA
HxKZkwP5VvLm75ipEhnMc2f72gH4V9RRNHMpGZJjQQaprwYWyZdJqtDpyAFPArf3v8VlNPE3+NNf
KQG1k++Az94gzrpwQA1L7po+fNwrtk71rEUhcDatO82obbAI/99gPA4gSX3XDQlsjytqBvETR+Bp
beRHxGgNpjAejMsDkwooRCKBPfC1c0sUY19xQw31A6UaGYj0EVbXSBlaLucDVYOMUXoPbvRnRcwY
dbX62J6wXNPUvzCpm+ZZXTAC8+89ByXD61ajD0OnGjQtBj5+3bJOMofB1ODM4gZHQMDlIR6fqP6K
6Lqi8kPJOFWru+Byh1eP0N75lzKN+u8scnajk2hJNTa56kGb+eck4b5Na57vQgd1YQEEzkHTNxFA
cuFVieZOUKLnN/AZMeBrCgQOaWyJCItHreEQKqiJIcEtPQfWterZ/ftE6LfEpM/l5tssNsN3qCv1
wzuXHGR/PVnQ6wMaoALNgDKXTo9orhhNXjYB/Yxhh/RBRKfmFis5/F95P0MnQVHiIuo5oQLGS8Gt
kScAfrsNW4fcKKA7wh8LwSiDeiwgcyB94iXU+VqgYADJL5a9Jnfjkx1nIniS/9GBMn+Mb+3POp9E
F3EHHT++GsekzJe7z9qfEpiF9/tfXzmCMjqsTHNO2qKhAEP9rY8MOMYY482k/Eyc0gHO4yS68YDx
mLvD7Fooiex0SgnwPiiu1byLCCEoLe/DlrsUeahfNviwKdz9ipUFM9fzM6MUQ/Hdi///umV8Ikin
91kQeLGNGC9ZF7iZX/QLLKY7OQmYLTRZ5c/A9GEjpRjCH2/VkdAJlxyPd2BzOhctrWue/JyYWvZY
yYcL9v0dCClt0efr1vMhwmovhAAFIN/HaIkGOnRt5YInW+O7o1LQ0lEasxdcA/vH0wjvo1DwG6u2
3IB22F4Dh+AE6qfd0HI9LUadhxhBFhosWkvt7vJS1iEjK1zKCtOyXSxQ/VgXhBMj1ndqIetroWWE
xSMWJ7sS6q+LSTyad0NkEe9xMmDLDELlTpuFWJDYrz2TORTR2xFdK9NIPbp4Ur8WJzgmv1+bcw4A
suAlLX7aYrJCedUL/HNSdl4uSwHrlwU5Otk2XZnFmkuvdXd4jQ2cy7mPeqMdwzFXuHIvDCc/xVwL
83zATARVe71eSkv+FFDccCPlbPj48TrATlpc/ZBKnzIHwKFLvvt0CxtylTj/4OdrhJoLBJPs06sI
/ijqTAjvFimsH1Ua9EN96bVCqGjY3SXfOmwiwmeR7SAt4tP+DgAu5moktSXuYk87aFh+655jw6xD
Ddv8sMmohbqeQoqDdYfT+hA2hewe4eegn1AgUJruAd/O/zBtGBZhYGM2/mxzhxXtsLlWBYNpZi85
Lq7Rc8lOtJ2YlPYn6L/vh2BF5pVsSLuJXN+L2TFeShSs9Jv99LLgeF6HLjNKvsJB1z36yIsZOuAi
tk/GBQWuFeUJSQtXyKnal2MgAG5ajJLHwrPDJivou29lE5vnUxb5M58fn2BwPUF68nq18SDFOWzk
sxizA9u2qlPBUTQU0lSWUUsIUCIkAS1Say0o3JKZ3tYUCf+B2XOxLASJbkJTCUPPkKB2gOSlxyTT
cgUsy09cA16MEftAN0cBHwBc+ggf1oQoquZ7QIzQ+GYE5fhoax43NF7EJ703MbZUWsOY090fhulQ
fVKOeE/fJa1ZoG3vHbt9KN4/vc6yqDomtoKwYIUCGSlmIn+PVFw0v0RXRKtNWM+ehlQlCRoj88P/
p3TAj0pKLIFqG4j5Bdo4BYRFSVPMRE5JTn0rM9prPgQIzAWUV/R8Zeqeq7KsiWnOs65yIxpADn4a
2XbSn653lg2OJl16MTMTCi6tOdx2vrttYCWzBduc+M+WMNpQAZU5oG7QpoJtnM33CsZY/bo0ZRYl
U+qV3zJBkw5031Tt+fo8GHDwPJD3xl+/lMic6CKrrv33n/4vG5kARItI4cOvdoUvr2ap65Uk6J0O
n3OOpzMJailVTCuEWW0jb4CT9XKbsgVom9IPsVQsDEiVNHZ1oNc6yyp/RMAzL5Qh1BhRhk3CxP8L
PDswYnvv7Svu62wqfU537v/Gqp6RLhP0Z2VH+f2UVzfiHms6pwP9DEU7ZPq0mpWyoGwS6oqqiGB1
CWg3731oGAYW5240tDkJuVcnr+UvQ1OdS413tXLnPpZKe6O6Y16HTZnXFGQG3aI8f6mvcxByU7Uy
l/ifDdcvSNvqpI8Sc47/L+nQdzYHUbHy5V89LhbpWGX4xi1tv9bHZ/+/ZSjoFvuLLq2o3TEV7K4d
NCG2pcb7N2aEjq43pWQW+XxassnsVNVBvnWEtocbZtl/9If+1jXX0GMVIeM4aD/e+O/fEbWzUOYJ
hBIShI5nXD+zW9vOo+afw7E5eFcOHlfkFLE6d2b8VH/qTqjEWbgO+/eQvTqeS/K7CHPUswOcsgP6
83MRX/d/9ql5BFyolzCrT121wdeshJOCc0E32we3lxG6M/J7bPf+6rWt+WHo/6T5SygMr/G1uAo7
i0IH19axeaNk4xdPMoNk0APVYskDgRrwYKd+yiD7fE/j3yec76jMAr1z3h0uxfzHjM4ae8XSdhcs
25CIfDeO55YMjreOfhSoW4FvFg8+xp3xnk2FBKMgN/jA44HP5NwX+ovt+6DlQRS1OB64XUPAUtAp
fvs/dPGFzQtvuNWbM32vnNTOzvA7dpZXck9udS/Lw81zAV23ytT/C/M7NCh54O5FX8kHqLkA6fsQ
zpy7TwKiR8XFyDwOHg1K1GKG3pvJmSEcol6DqLUX89yMBylqAXMSHAFab4P5fTFwfVPGNtZEvj6E
rsA5RQlP9VrYOC52Rm3relnpJXn8YTnZQ4NH1uFzf/X9A5FrJBcyffjVVqnuoDxYn3C/W3M9fpfQ
nd0cvCrHTCb5hQsHk0TQelffrrHzWAgt1HKXD7wXJY40Y8t1SGn69wN60THP9ZGY+FL6p9lH6gI8
N+lXC0Ao7Xmiw9w2w4STxAutZn6fQlntIT9n2KEK8h4lszYrmq2IxjKO2XCx8pX4gyqOpUHt5Nlg
0oOuuX4gg516lIK5H3qzpU+L5SV44c5iMuh3yClXnztaqIgm7Lps45FybusDucmcsPdxx3pZFgnZ
3PfNlCIDK0Q5VcrGJeGApC6+BPvgeNtB2xH/tCoz1pIeYBLf1ZzBaA9Lrz4wDErQjXYUtW3t4Ro2
HDnA9rW7deQfJVkW6zKKrBK8pq1SCgvjYzwuOFsp+KrqNG5g/sHnHEoUKHrrT5y5ufK9lENrhmPB
l2x5r/RZek36PT5pQMHr7sYiP20BPOBivy5FnL4o56+gQVJPv2D+QCjtoeHvR+vXFb+Ypmr0QUGA
rXlO5lfsjg5QVLvSL1jdA/4QvNp5zo6tQk2toDt/xM4ftolu8P4yUJ0vb5CVdg6aSI4G8eZbYj53
txoPSSzSiEkYWX/dqoJKOTKqVZgSYEgW010Vrcd7TAVx+kfAHszDzuW5c6+yEgNjKx60dPE6Yhfs
q6YcXgdVY0WaAQcUKvfNtWSJ5/j7mLlEtBMPZnVhCDw+/K24CEfOuNJ5taPp0g6k/4UB/4XGJYZW
CUSFYlAg95msV17frRF9bCXeeosxrSDoDzJ2quLCVGKAVGcHKP/bys1mwgl9aQBggVWwLohrJgqE
yUnADBw3R0GdzjxDLENnz5517OzqE8GRvvVH+lQOeP/aME32HcT6WC7rDILoYFYrD1nMkEzd3+TQ
twq/NXSwuuhTgcUlNrC7G4wC6s0HkPUe3PyxwGvQOqjKFNUIuJTr/a8IbjwHkIHpufh7/xvRPJ46
LnLGy2SVwSJn1ODVNudkC3s4pseyPGmTW2K/bpcmFWf+iP/SzPaF4MTAuWpw8Hlxi2nVTEsnD0/n
ZdVFBMnD0W4p8lrxENA4a1UznEyVE7JQvcMRQiui0W8HiO5UkQwyjNTId1OvRa99J4r0nErj+04r
EvnpcRAvqe1k5VGBhER9NbiriUAeMIHslLxlt7ggTAqctY3tIwfRIbVg9cr/CWyRDCSZKfH8svZi
2qsiniB+KIBU1GLVxlCkQF38puNLqnLVrOH57RUOEWMjA/tI45Ay0Rk5prebHHu6Eq8qPrqJ1aMg
rj1J79SEdxZvhFmkvVbdHeP2Pw/Zugh6bwQ+vUi+u/9b9tVi/2UXHo0+O672OvcGECLC15cOfcoy
N8EHyorZw1rwFttduUeC9oQ8mDy4gGdu24/iIzhPL+PcRERJ3ZTsa7dCj7ix0UjN8+GEWxI0ZwPE
VLSc+re2Lx2MxROwNBFsRl+LO9wojZTyae7cC30EOWqpihngyywxE3CjjDbRODLfs/tpMqksXiYc
DsFHuwQOjFABZX3LlidfdBLTbaQwTtaHXjygsxWAjex4G8Om/cCTX10UAQdYoIqP9/emZ4BPj8eS
9YBkiO3BovcS1vTul5npMs0sQu1wNJxKRP57Dxb8eADJPJldRuT/BLalifOvS3NUULF7ljt2TYvB
9YZUKbjaRiGktPfnJL3X+OAyYMSOQ/XdLPh5WbFgB396vFD12XTn3R6w2LvTrnQ5WJHOJli/DA5L
gVOVfnv4jWm8jmpNI6VJG5S58C8KJAz5QMWXMTV07/1T1zLyWiBi9zzWGki6XizCs/m4zFxhXuqF
mEEjXRil5592/Y9haip0fGiaJ2dBt8l4klgrnw0ArIY3KMo3nnwx1r/lTH+hgRo4teB2kSTpwBiy
sn0QVeYlwCLUNVWbudkTdTItghpyHRcDutmGZQGYoun2Nk6VTKb5A1Ks+1VT4d7O+3qu0tWpE62v
l1LIkp+pU0uakMs4E8ZVG7a5lxuYPtqhpRtw0QRShuTDUh9b8KLCNUGV/hd628foSZIXZ+/EVYz3
1Bit4wNkcyXRoOjAPl3lwAZc9rFg+zHOBZnn/TGSyC5JS4D/K0AXYnVBWyPDkmmVCjSnQfsAbkzp
2/ZbdVWuqOLn8iMbaDXZK5roc8KrK5XAeZoHgh6Jq9JSSysdHpNcQo0k6yMqPsrUmP0CddeGFD0z
VgtYwNaN+IuLgWZ0BLieG7sxih2kGTd7cfA4t2PabOoUMhAAedEvCBOMfYL95drgL0OS0uLH3y2R
ECKpVFymOz/aJ20gDuzaF4eA5kaqZ10OQ5O2928mkxLVPL5WfwHyEQ861HXYUm4157v9GW1PYJMO
7QdBBfie3yHW3WBXE3GQW/A1F8RaUCZ9OFnaDSaY3gzZNZkk7IjgcWAzVYZw50QN+/UlKYLfalac
dfOFNG6AFagtjNKQUSYHdXBOxvZ9jYB17+v1J+y3lDWHQQ2Rfh5/BYS7KFHampfe3mWyGD5zGISu
PXwxtwgAaUQeHk5UgEzyI/DFhBpzK0wBIN3yizUTEjuPqt038t+ulefweO/2TWteEPBR3YYM0rEm
x520l91hMJAlRIAnshNpu+YIP9+1PdsMkT3k+/cgW3n0HfMXLgXBT5JWWL9eygH5vbCIHjTybmz2
vbvexV3nkEaZf65iBbH/zgkkRzpWlN+5oXLgq2Y9SmCxgpCzMIoIv+oBA6ZKiHEQoVsiltTYlifd
RUqpjcTAOv8M8vUU1woHE7mkUASYdGJhgpmxqimrxQgaOEBdA7RCH58F9P7j5J5lcrypMNBTzWG2
vyULh95baCOunyY+rqWEZvf330DwHVKgAs+9GZsP92AO23tLuESg/Igl7E4Q1E2M/fkxAaw+AwxR
0tVdigO3UVAXxjBTZOZO3EW1dK9lllTZrrT1wTSTmy15eRwXTqP/omxJakm93oku+arXM01bbh1m
GKh50XPtOG4ZHsJcDUnRxjRvHmS/E4GGHdxReKDhCpZ8iIXamlpllcRywgsrbMDjyuR1rxmMWfGw
6avAXnTeFTH7v/hkQL5fl1j4jr2QEr93GkSKZC1RYL0QQafskxRc3aZhehBGUkNRmPCtcnLXNdBR
WybWZTRnwTLd0ChsFSlr8JtB/xl4bcF+OerpaKGp1R8VrvxI39abofFQv28lGs1LKLEm6LOLDqdt
KPc1nLXzUGTgxffsF64quQGog4vsE1zjEj38aQsbeH5KXZusrqnZptYgVrKnhAbTXCPCnOgHBZKI
/YH/dTPcIA6lhzBTtrIOQDeIgfr6uQswpGICYA+CZdfCZ1wbRtUWInVSGLDajLmhjg4zOnMfDwj4
KWsVphZFaecQ7hPeuvn9ZVeC6gRAn/IliztSvZRvDKMqMFFAjYSAn1CZqs7BJMl0I9xcEjD9N7af
i+gbNU6beMllVwlI36Q/SkhKhUEjJCh8gMLchkDFj2HyT+qfYUsnQTmz1BwTScQrLrhzmJi+pYXU
C5DGLbrW11N+bZDHNvNxec3Fm06d/8pUN+0W87NzwcUiW5+glhJlaTG9gHzUmSx/UKXWJxiSpbWz
Bpq6Cd+/ywengLenToT48kDyAOdL6zklyW54Xdt09qIxx7Vfu54YM6P8VoE+SrKT+M4kOREXr8Fi
nZxMW0/Akz9vzrX+KIkHEl6hgv8jAEveEKVWb6iYY9K7c5mlAPV6rpY+1xx6saHenvmf4gXuIhQR
uTV/iclkkxcQjHF3k21akk9rIP48nKtatGWyPFa4brGB/9txKIY3Z9vS8guhYbzC1JSOOBlfRvo2
nC8BWqcvi9fKxGajkBhNembUu5w9W7eCOqSPmvTpadmUWGhLPaGPmAVDSlO6KtTUNbK+hQDSrSiU
YfAIvtklMnlB3rRDujMtB+UIi+3qGA8tZ095vpg8+TCe1PVi2RPPIxz68rs31+7r2B2F+QLGM3EZ
rSFrFP8h/zhlhBe9xTok0BPdqa8L/gGihQEpQFKKk1lq7x/fP902a9KlrefV1qBaRGzRFygVorN2
mdAKE/1CIMks8u7AzROe+MWg1o3HLQqLNYpl5/TZGMkVr4TE8t9xoDyWP1uchjZ+sVE7c+wjGAig
ylCqUjx1SbKeYVGlsyvlRgM+hr+oaVS55Q/3U5yz7qR2kQzvTVhxhodFFHxAq7j0l2LM9b5KglQy
1kqzQu1o814SAaSRUXPrANSh+1XaW679EwzCL36aGIqM05px0xZP873EPXIXNBnk/dn3CQm5g2NZ
npm58pH9w9GDyiOBAFGv9Ry8FALV6EbKTSf+XVQItyygbZOG/e8pYhogsvH7nW36XFvLwwN1bMZN
xIeGfK4GVRr5CMH/cCRclpJpfddkhj9IA614G7skMTQw6otVCUf3FypAEaFblY+V5kR341em/XQV
ZUBsPhZ0f5DaCf6MrcPpHVoxljlqNCOIR82LRLmkDJYWz7dI7rC/4ETbrP0pOGlBHECG6CVE1Xiy
G+pUQfqcBBy80LJoIOguCAWh3ttCmUKBRHBGqehV1AmO89U089uzI0gQdwJF1gKLhI7KNDr8nS7j
syZVjWRKm463CnVoIZoN4i+MaO2+gvtE5fno2tMAYV20VYdX8qmt+vCcCYdWEoVpN2MQZWIn1Cmh
Bo7Cq1+kifWz/d2dp/viOm3/cLVVmNBi+Wj8Fc07BPWGnccojgqv6mbTnMSlQrvcm4/rqQrN6CRW
1Cr4ADQK5hUJ6yf1D8m9PgoFowNhHvauoA5RYR4Qv2dmtq04yUFj3K9ekz8NAY0X33J3rjAWGnxI
cxok7csoOQZ1jMslOU5Eq9JOXflql2eAkBVvless9Vj/rRiXVV7lw3+agGbIq0w3He4wmcFEG+Pt
hgnV7iXetDAvLgOS3pO8caJ14Dp/cdU2XC3uO/A9+frDSHWwbsXJQtC1voto7E341aGykvdnFTKJ
DoEe3XEfuBsY3XCeWeuc+HdIq6s0S14zL+/n5rDCSMCfrmCAPk/nj4KB6En48EVOXSaZGrJKvrWg
JexpPSvj5OkUbaAhXIn0ypYxGT+qTEXWGeArHMB/VqQY/ALSeX29YdJws3+4k1XM65iEMtpROBu1
1fwieYj3URWqBoiQRs8xAduhYCIuzr9PrCr+2T1KxR+2h3zOxL10kCAfU5JpSGyYDkf2Q0KcJgEh
LDlz2btfeYLQ+rurtJVIMe1x4cWGNwxhSGw9a2xwZXsYTtjbiv/Se65+BOSXbGHde3Q7gmaO4Vcy
pyUjM8+THAy9HvzrxV7OE422S+BjvNnaCE2KW4B9ATkOyFaYBGhqarHswly+XFEpYfV0ozwpm6o1
BfC5MsVDCOPATV5HxJNFR9T+65+6JxjesE9DtVRd24Q5DwmrkcADS03vMV4IFMhe3vUCF9EQXL/S
aoNzMpUd7H0BxlruZt/jSvaDakBIbdFrRmC3QBHQ9VurTB1D41c9Hce66M61N1H2qWzBfksoeISw
j+Lcsymro34pcysv33hZAA2vLotuhXsP84gVzD20HdykvWqapRS01bGt2iZpGBIo39OxQhfVqZfa
m5lESZvH7dygxepJshe66T9QgGDfElXpOCde/7v5WCkuew0jH+v7b6FqUH7FW0V2VZDQ8rX/4F6i
qF0VoP8W2ccM/YXw8wKgT2nTVMkTqze0zphWV5B52SH4uwvvLAQQ75Vbtz+oCFzQUxt/FGYatnRU
gCQMuRD+UJAksNbtac32AWYlCvXm8JAdfmRHLmu8/b4g/78L2EW4P1pbpizJzsvXNLz5cxmF/jd3
nLEqsIQPTef0utwkFCm3J3UCyoRkWNhKA5HND0YcCce2Kn9GI0KeQ/KnKg8SbBaI5/bdgzK/IF2K
lcfi9WrSIU6yrP7yfq1uLqa8hiUawdKo/6cVkmdyw5fFmX4ZE1Cq2Qdw0VMmKVudy5jy8NAU/FyK
q1oqUw3nupBQ6CoCWv1p81usuBLHsatIHJ2I6Y1TIMfTtEwhnnW9+wH7IizU3ON35JHECoKS0Ya/
gxMj73KaP3SNvBupYYXhHLQNmAOtUgqvFk5dRsD2FGjHv671mSdC3tJ0kMZ4Xh/w1NQ8EovpZVlx
EuFB1vZ3e42s+8Q9YeurUtxYBgSO2KwebL/YYMRnTwhpji8/xDumEWqSCvyyNJAm48/EmKDQjrPZ
PoFTnRolXS/9Qw9yFbej+4HWXCJTN+Fas1jzqmwO2RmvroZ/yYp59hCfRgv7IeeQDROrkqWaijat
VAcF0pSy6fWV9IkH8fmH1HbjLoaWB8kSaRzaPBhiJ5GRa3L20yFpS5bUn4nsvYpZ7MLsW1tpP+UJ
3ZtQRx30lK+OVG1DZC+Ji0iP+6YuHyj93A2HLkIAa0rE+te7KUCkFFgIVZcoZcl3j8CcWK2rJfnB
Ez8MJyu8mxmxiLRwBUGVAIxESP88T7IzeK0TjI8quCWzim0plpSN1qsHMzml3/5QBX0jiGvFPAWp
+ZUAv4s36+TTKD0/cfm0fw0mhUK0kBFDUd2VnZzyaUQrNDkimo/vKqJxnPoljQl8Lb/gc4ZGeI4d
PSmzK1NsC20o9V8WQ0yaEix34jE4//k1qlIXITdAPr1ayRaDxPAXuAcCXIR5OuHwDkxGcrpSO26t
ulokXrZVxlUVQPsEGndIDKnQRf7luYMiBFOxIZ2b/r7SduAU5IGthNnlikwTJY6/UIXMAxv59WeZ
x+pG2CmnLpqvtY+k5WJZs3hTVp1xpqYHsN5g1Qspmv3nt1TBwZkaxUBfteNZnJ7fSnDtrb00fBex
3H2BdYa4RqEOlecDTusuv8BGjb3bqi4iTO2vqVKLtKT661J3x4WQQXvtrUZY3tKGKelfudJSpHbq
2uYevqS6H9CNVNVZd4u1Oim9Uwb0+ttWe0SHv5t1zPN9M73F6IdD5MQfkzxKSQoe/3aHRM1TImnH
qExM5oPhYZizWnANYK/n32j6MHFJjKAu5WifREXFlTG7oM0bNWUdeUcMW8eOZVq4jc7XXUOTeyLj
Q+dYfN66DL6iFb9Dt2KIvXfeTZpUGOy6xkGO8ppXpFXUNsCK5V6ZwUWVqis0STDrOYF/n6F6CDR8
UUrlJmNZint+dy54BihS7b8imyZjzByGyx+cyfiyOeshxf8VrZTPZ6ajMqjUtaIWFvy79La2usAI
VqXlHfuC62gFhNDWOfMqZgLiambsa20V9aaNIvadIu0HfUilAwP0y+e6sWRW6l22fg0LKSINL7yq
KD/Rw4sXGI44nJxsf7Shq/v4Jfe0XZUK9EjCM8074pV5thZ3uEwHZtskHuBGlRdGMNhYkHh5naan
TTQDXTH/Ig78r7ieLOccQiYIp2tciA6WMZGfi6ij7aRWjfO+LlX0QzfyUuTK9Ode6cZipY7S1rvo
5w9LnIuouLo8aHu1WRkmYdfcjpGsuCZcnWTFvfb68+tMoNHOLo/qYOe3T1+KlimKbuoCKcuQyu0x
OW8cQ2gGbmP4JxBgmst63qv5+amA6UYe+O2dHFI5GLDVSC24rxYG0pq4OCb5g1qj5TjCCpsGVBog
MrKVxgtI0N7upaLDABS00KM8O+83tPy6Ve+i77w/qOaU7q0pcyC/s6uHJvBFdfP5t719CO3Wv8tO
3XCrSxV4VuyJaJbXAqP4OtCS5hNCzWzOY6yk8zsTpd42XXvR0DgxtEw6ePcGbtXmNWoI7B+cHggm
t7A8JE2nGKhrdJALtreWlg0EScEiHTK+L9HKrhqKviV1K9Zxjk83ikmQ2Bzc3kzJ9gNuQBGqWWCL
3UaFZcQgZAV/ExTjnycXOdBo+md6GvUkFdP5bmbCdpAyWI4yycvKDJMuI2i3VrUSfROUG2658P/6
+wNpyZF33KGg8ptL/p10PKdXwuW6JvX6kBdocoL8TVgnesj8CXwn+pZ/Ewf82qcsKtJLEvtd4l8P
RZICfcH4ce0py10X6PkCF8X/oZx+quT/1hIOx7cb7Yy9OqTdD6BYT92XiW3+x5H6B4DEL1GpmGPr
Nkaxxebh/tv9ht9sbGBd3nDQFtpH6m/cQ1l4Qpo+eRzJu9ttd7esgvESEy1lkhjCoSV0JYZn0nr4
Z9KXaYcKq4lK3GWEKCt/8G0HACqZjKg0qnFJ0gsi1O4d6OhKtUturbqQNgQW+xxhmcpG1dGAx+Y6
KtH7h0pkhREhJeHkf9eOLiXrP9KPqlYwJ7nAdybKVvoEfOclXG7Ow4cLYGs/gcrcwnimxiwnK9e+
GJfycWJQ0oWWk07SGVE4exY96zq2Ed/fyPX9ZrTfwmE9FIfQQh1WAtT+yN/9pSDK6cOAkycAck3t
SzT5e4IjMD/A1a5pQXM1Kk+b15WTmB+OdrFx0ft+W4K/VpPmimZfUSerVXlNnlNDDNuChUb2Nqli
7CoVRw/amkjPb/g4EojbZFDrrMh6LFp2L84jGZ9s3G/ZWTd024teP2TwQxo6JgvZY5AHSniu3mh5
QE1c/45rd/TFgXPvZpUcmcP3adcvgCimftnHS21FiG6CP8p40HGS7RB8qFJusRdPgwa0XvR/+CBG
f6CmjLMc4OcJF23ASwXKw3h8MqIsHiUytqFDj7L1AEbsS9/2PMlvKxEM6G+/7dg43zYOamDk9JEi
/s2lxFfPD9KrxtcyzErTudeMZ9jRvij0gAj+GWELLnxPsy776onxZQE+qUL/GHXapbSiG95CoGTR
dRKoMeslUVSGIMusoluhu/eZ161ulfX2z1NLNGYbpCVi5bL7pkAaApjwr5hQwZj3x58KAeVINhyd
tBzNapvrA1C5QmweGu7Lpkx6IZzGtGhGRJJFZb2g9Pbq2O9wPuIAKaYJM4syJNcNB+lF0ug8o5j+
vetmYnOgZ1A+fiuQbC6gIcuQao3jxPqDhmHqxrIO/PS8QLINKMabAnQNjLnx9xXCVldc2miorL5s
65dneHBZmRCDfq2zR++5cYqhXP0WLJXQ+/XiCJrpxUXBjvdMyaFeD2cJX2dW8Uf3ZToRR9nkMvh+
UKedAeyJmV2mpUetKnLmdrZ1w3Ma4LXjudVjbS/9BSpjaB7yV7EoNO+pZP9EABihC4FQU3Q5MtTI
7cNGUMvj+bRpRu9PcqnLx8W5b5QyLDTNjgfygjUMlANZ/a9quJ/To4UxKrxDTwYOFU/Rph1CfJSM
/PcUNntDat5eo2FjiJpvjWhOgDUfjsVs5FzZKvHrRy46K3N46u8frXTKo1er6cGqpx0Lgcqxj8QW
qYXkTvGqcgZjsAjqFQhpCVGSCuVOO5wN8LDDbSnvb+ZraWqrFytdvAK/q+jDUS/fv53ivZspv18o
qRRoZKb4JZGdKUWsGE8eNTjYtBuZQVx1Ip8UtgmftIz++EHgkbwb14YDzDclReBDSYi9aM3W50lm
TMrtY1yfg53WZdUCod2IS1fmZ0FyFtBBKzG6LGtdVOnw/HKBjr8DIE5trjEzkeP1MWYxmG7GAYXr
4AdGXwZLCYq7mpyQPEg38jt3t1c89bOmsbezIo4/8eTbJJRyGPpen04FkBVxSXqbcgFnWgxqdlnZ
T+xbvXauHlCDQ3EFIDn09g+0VqixieWcxiY6GzJ/w+5I2nu+o2FgE4X+f6AdcUnAvzbgAZ0WkKhg
D4TkN35gEqZZDVkSIqrfJkh71EM0KmJL3xzH2wP35kE0mQKEyR2b87ZtYoFQv02x3YmM87Nn04Ce
0pdKdmr73nDKeRi3QQKxeXqAeghdt9H8uZEg1z/KPbd5iKZIyvgZeq/ixEHEQ06SN74cerC/jdW9
2uS9eWsLUWrtwi54eGhLAUuDwyuApsboEw8QQkrO9XoQVJ5YpW1sotXqjpBABbzs1kupaxCs9YuS
HQ2JipxHdCxr6MDNvBFjtmpCKoO6p/5dc1nGAhcDCYfxoucm6/uOIfltvdehp3s+7QkZKe5c3FhS
QZLzxqIpg7ePpkRP4fg3Heivl1YDkI57TgWiL6NJDMThr2GeKNQCyK7g04UR9E6j8khBd6Qoe5Tz
MpwacpmimfAu4A558eml8k9Gwkk3dGvHHOqsSNY2c7me5fF28NDym2IjLdM59vU9T/wddiqNpGVe
oWQ0PbirF3sFi8qwRVl09tnpPrBiW7Kzc5rEsMdKQDBT0/aB2q1RgZ0jzSU1kbPopBSKtvibxrLn
irYLsK7cBm5RPUdSPG2tbn5TR70jZxbRfUZre3KXPR2dVyLYseE8/3h7ORD0SAFsycrWvHwHSlSu
sjclIsAaH/yeTi5mwm+KwsRNptvf9cupO+xy6x0B33MTBSVMcmiF6NwVUV8dXBV+a01AaGeF3Wz1
qmRXOjHMLWqItmvgc9KupOTAVvozRrOinS6p/fPw+3PbVduwh1eXbrloidzpjWwxU4z/gY0DLnCh
yGw7WT2r+ctnPBNGufNxbBUgTmHr2yBhfygBqofqDjmaklwwCj63zA29eS9oX2Xov+rtCcVrZjip
YjRkpVIDEwOPQt5DHEH6Xw9HklW6qCxUdHuWdNRNm0jHeDW1QKeg+P6k71WeEIfavzQpVKAMGzJ1
kaaCbn/ZBadtDT5q7qoCZBygPN00zsAF3RF/z15Ocis5lWv9v1bb/EUj7mwi2R8ofi3RVh5TWLmm
8psC8mDFdAG+HSRq/LrXsGXVLTZSfkraqEZJf6xuLTlfWSu/DWSaPiOPJqE0mxtpYEOj0EddWWPZ
umtGDbKziI1L1XEQpOUFRhfZgIs4rmOXgMDogQ4MBdKGJCRCUGfaFNaKgiU9hkA6xxIhAkgH0fPo
EyQBag4rYJgfPLBsXW8zmAmUhEeVvbH7lrlGUEADppm4Lev2ZZNrsHXjKtc+Gvw8HKfLwLy02yAg
fW/Ys12FeZD5Ei9OGkY075TdLnsyDOdtgbkdkZCqTgtT2KukXSlkRRkT80a4NgWgZgaJ+OD5Sb66
PvKLAdsQoPrqhGZBFnJJ+kGOxoj3F0qvANDfxPXx9oV8JdxgXbCNX8ubSdIGN1XTpSk8oD077IFk
HJJ5ScWKYIt5iKLY+lyvhjPIsjpRL9Zf5ZdoZayP6Aa7DINKidLM+3a3a08QF2I5PqAObUX4+JJO
YsTeKAvh5NZ3m5yy3ORprCaDgGvuOImEdFX169B2czh44chytbfh/VWP64V6E55JQLeku86qyVRR
i5rtb32G+ORktABoerz1SBkQkDQOmceyiJqh90F2vwNnfTy3iOm6Uwqn3Zz4VbgD7QEmK2L/tYRc
EgUcs365EKp9fnWsO2RrdalZpLiIL778XdOBaKO6yMmwLDPQCJRoBdQ3kZgxsDu9Z8vq3DUCzoVd
KIsaD6R7weo4QN6Z6qMvxXvDnxHcvjL5RJcYQzJwtcUoI3WuRjxAR7/3SOZUNQvTIkkwKoSA+MpI
SrhrP1eoyRiVMXmFJcSMh86CG1MYLSYiD7VfI4d5E+gpcLxh6M921A6n6GjVO2Hx+6giHgP7CNMS
cPwmmX2QHa7O6aLjuPqAS6o09RGxp7dEplie8OMDlnJ4ogYl0s+BD7B+WjoxoRuAAmV8ZcyuwwUS
SUyinBqWuuZFyrJ+SWXaks4b4H5AxeVs/pLH4N75eXRu7zBxrllsMBruzSNWFDqGThbmcRYGCWk6
Rjgjf5tiRF9CehfHpbpBHQlNLfclHBKSpFrTmEr9jdPdOTQGEUprrh9hmpA281G+zsvt2lh0j6g8
p0tL0PqR84X9BLqknYF16gZwpY7q70Hki+ZcIGik3i+2rBScqEWUgAAvW7WtrjymH2yDJTTxV5v3
BfPME4myA6K4o9TkB15OMKPJWM2ynsqxFRcglNu69FowB5X1vcvA/ymdgNeC1Z6icPg4ffQn1hWn
wM8a6wa6jEDLMCEw7c6B7w6XQE8VNmgvfHQhKLQd2Qjms01MLYTxqcpLNJW/PBBm20aBjWgh1/ah
5/46+Q2v6SznBa4whzYH52IYGFArGnd02fAlXNUk2Q+HOpLim37ZCo1eXvbCSruVbX12gvSCSs1T
0CUPmpm9NthGX3MOa617V85n1i8Evyaq9+w89hSB6m9MXx4jxWUmZKi8k1xdVa/5sbVFduDjdgTg
+bIs6hP9eIE5Hp/ynHMo18tYXgsQN+vWs0cZ0/sjk7Y5XUtHBwSCEI4I+lP//2oRE9ggsVGQ3e+J
prH4gkPLVvfWU3RUMXIKDcyMjcVA6Hs/Cb7A2VhQz1xHy3h1RWBeELhaRd8CRszwdYUXENRhnEFH
u7O+dNgDJL7DCWCKVA3m703Xqm97Skjb2dxeck7v9g2CUJYzH3Pk34EgdV3mecGFlBScnMyTSQAh
nt56VSvWoWg1xZFOpKmdejzCMnwJ1eeQYJb0bCOK6q43B9Bvv40xgZd0eshrZo4ehXF4WIKi2OBI
i4hnJa+PeuSNMpl71GgmwFjplG1mqW5ygLuxC6VkN420+VD8R0/zOf+q0x1rcjVqwvu9CfYnmwWj
ijvMpkRguYRfiVQPcrV0mldSKYrT8A+KraQ2B4eSjG1ksZnY3NzilrE1OysveoaQWyb6szCm4Q0x
g/064R+st5ydO7hVvc+yyOw+RH0yuvt49hehySgKPw2gKam8yv6AWvQGKFiTmzZILuTXm0WmreNm
JsZtiJHTJxb+dLbn3s7y21h44u2LDGls4sTm6tHL8thzxbikQzhWOCJQFxnuwFF+f2r0pF72g9EP
4UNGliVyUlbJ0URRVsDh+G0NQ1KEc4/jXppNSETfoArehfI5IhJqfc2DC1FtBH+MJ+dihlxOBshl
xdBYtuBroq7JfYLyCdWKi7we7aNTbvwooRFRtHeK8/YiVHO9vPl2Rc43wrOtBlqE+c29A/VHT9fu
q3QBHBRuvvJdrAlYjoP4ctI/769PmPtDOEJ+rTki2yj6IlsJ9qmM/Ok/bDkFmXRQUb/W64QEe8bX
TVmgFDSaWuJuzTBc/LcUJxj9WeUsJULT6rADbjVIU535hhMs73TdkHqZ9KYRMPE8xVLJ9n8vwPen
RyKft2ELe4SloAjZB11ozAk5k2buZvawoi1tKqEB6D71IfvbI1XCsqst5GAiR3UH8f8666jm8w41
z8KnUMHxwIzWVPE19c6OQ6b2/cvvK91/3h5YzUOB5yWoa7CK7VLz5IiIZcm1inYtgQBIio8f8C0Z
wJMtrvwG47pHbtff8lOApgv3A0fBFI+JIP/eIASW1jdZ0tRGtXktOCPudkH1elxhqPQA2V8icpTh
S5dcmNRFtM5PtLVP4rzZXszZs8yr77hA7ke7uKY58AenOAVGH23MQG66rdBJaPUPhnLOwsqXKyGl
xRoVb0aboVnEGnn9wnBDcYUttR++37PO8KwpD2hzg5aKhGS3cg6zJ04PDmEsFLMS3sXq6594edub
FUpym1iVPMl6B3AfA72kVb1GjdRfGsD0rsg7DYA0awGvT23QXgMw0bnMSP+bcHmFdIwdbai47MQr
D2i7BBDUMn3P+778WoZkGV2Ow0M4oBqDfCDY/nhan5jqD0cn5Bcf4v5cMBV2dbx23vgyeEdpRzd3
a+QwfnZ6HsnyPzqgtV44hWKdFFbONeJlJKPpdQdkVmtxzfVlI7yDzu2G3MAa7isFb1LH7FJAGDu0
GrkllXI6K1LZUnGWTyMiFKlbovljtJRV1Za692G+pZTF90w6GgBMA7lzyfR9eFIrY7pHp3PK8c0M
miOWEqKaItIlmZMhP2hXPTWacmMQ+Oxxsc3Q5SBE2o4MXEwmELIW1b5bSRezIpXN3Ox6Or7fm+Qq
nZetocqY0I2aHOMdOv9MAeZYtkFldtGa5/ZJ94zV+0lRD6m0dzCNuTVi+rNc08JdOwfbuodncWV0
+HJQ/6DCXQw3Yn7XL8lwN3AbVoXk/kjIo9y5d+mJEPPu02MhBiFitX3/SY7LaPnN8hxumvRI9DO2
DvWMkxlLZOhE2Rl970xW5uKD12iSJQtDB3QHZfQydTnsFCw1d6LjJ20jxzNmxvD3vDel0RSyHHge
6lG2iwDPODqV9uUNL/14UsGRIjBu9SRPrCfAnN9CzzYBvhQzgoD7SMvh8/rawE1HOBFYESzZ8zb9
BR9qsp9YkVu+qngZMU44qr2I0wWtlbwFLRILku8QX3qMOzXec457rCt9ScpFv51PX4GEmqH2TEbK
TlBjL+ENs8JBXkYRyk/QlNK0lse+uzYWXNSffGS/YeDWQqEonn1RvYSdKhGchHc8anHf6CkxSsl0
nw7121Kpzjo93yN3u5NFumSnzyXHM+Z7Zt7kJ9tZcHBB+hlj7CgaDU5M9Qs4+n+C4YE/8rY1PVhm
5KIl/k1Ych0l2sXjPDHFkAgyccxq5eCAmrI1mmmbk14A1I4Ph4lm7eWGADcalkkLqRak8vo1+HuK
umR1enBzgTuGr41dqtLDutQI33Vb0ubjcqUuEXm03CbzRrtu7BGybq5zzybebBk/G0rYA/jed9l4
eRD7ybT1ynE2vUzWZRLP631LXuouAj6bA9uDKS0CbInOyWccvCIg4Kjv4wIFUTd/ci25J8A60JJ9
qxtNRBnK23ZAIBpsyalzM/geavyBJF2ac9e/4OEwdt/xeWb8ganZxxoELxPSyU9ywkWbi6JGfXV1
vG9ELA1hBafXwa28L8J8lEim0taXQniTKNQHY+3+L2aFi+vp+uOUjmmdgKvu9qiTdV6DDMpMaAvx
bKhZtiHbEKJ5OC5GeaKzh1Pm7BrzCSXvwb9ZrmNGjEgU6l+1hV7pdtLM6C2r/tNVHE7NexhXbSb7
o+BWWr9gDxVhmLr+SmDDU+yfdJ8zDJliZVxRZt06sn+eFAZw69kXaNZ1dhWP2jSTdbQMqo/TXQz9
VmpRtx9vorwPrtElsT48OiEvosQSfPUZzZ5w0maSNrN/2ztRAGCL+qjNdIF7P0w01ZEGHLt+HBkr
dg9VaemO4cfhX0v1TgFvxfVan/9nZfUxsF6Ph2wuQUjss+e4E7y1miUQEXkN9/JUkXI2yftjZnD5
GNy0lw9NESnLsEH/P7b+K1O72+fJj7J2NSHfLVEmwIlvvQT6s5CXH2luGESs3lQF2ssB9s0vPlbE
1C5GgbF9mLEON1pZJUGb9YiHD7jZVP70alBzQwg29MvHwtpqv1LyZop9coY3W/+dYb7Bhzab5TOd
8VabhEgVWUXJCoPLgM/flgAfJJnmjoULULbVcxjvy41DkRHjgBF4+6jEWR/sZidJWlDoIRcmAkGR
9Q999qNChzdHXjoE39AmzU8cDfeWrgvahnGDEwy7UJPoEuE15G4Tjq/SyYrAcfbGOM0jZRBqKdon
z2HHeVDJodv7pYPhSvJW6Gq5EAsg6atHE/h2rDF2R2eBeYJm4QPNu6OojTvF3WMsXzCP3twDMIF7
8LM62uD5MEYACOuBXQf3VQaemvAhsXRGFLitJRK3y0VQ+FVZ+BAezROmEzxyzRDJDj3jllfTzvCg
JBl6DVSksYb6X9B4P2zuT8u+h4z3pyoc8ZuFWp634Pn9rfAngIl/LQ2P+4o41KaqwaJH37T9rMrj
8UzrZ7sMv9nO4P94kHY3IPbN0b9n3fydlyYlomAwaz3TJ5XWFcrAiXdCfW/BvU2CYJQC41sz8EGX
jmAyULibTwO67nCkihEqx2U5kE2R5EZghoaHJ+wTETtCC/ehCVmMnFI4Uqqp7QxOgZqblLQZiczj
+6uAsZkCMu1h55S3BQLjzAK/JnX38f3M75fR9KFe/Wd5q1/T5/UnrlhDzMWcsaniepbwWKtSCXc3
e7G95wiQr4GFtXB7Xke2FmHwLza0E68VqWTTD1i4zzYRsAdCTbDt6YQeS6pP9TkkKR91HFnroHkS
JS6n0fr4LJyCw0S68AyP2TVzVxT3aq95KtB1/bIcP5fGL2e8bQfJuSixj7FLUO6M7BoQL2o4I+Oc
xjwXBhWaU3uGO8XED3Fk0IIUIzu/qMJGJsg0+oG862yM3ZsWxvEv9xih9oPeDCeXzETq3wWw5U8I
eQlawFYs1cRtExjZLrXCNqGg2yglSHk+qfUsbpHxqWMC9VgyUhvDRjDq27mlxK8Io50Druia3S1Y
Lb9tMc97INZFSlcZkdYE49P3wUtdUNjOUAJlBLhnUbSJwBf7knYCKrDLnAozxIa6c/l4aGmHSV8t
m+W+dca7UiSfG1txt1OsBMxvUd/XZkqrSBt2gmIfCDq5bsnVmxyeoyMiY40aR7Mo5c+TtqJuzQzO
7TxMeSCJlgSJmnoDMU2u3L0bKeScBKE9x7CXPLeLypzEnMGFE0r9Gwt6dAo/NRcmuTbufx8jUO9S
ss0uvPY2ZdwcU1XZQ9kR0JZuyjudKHocBp7rTtOyn3JQA0C6a7vGioqQW62umIOcQNGRc6WbCYOE
dab6ZR+YZ+WINLJ+ZpczPFRXOrvrX3YwTRqOon84VgUEZ3TxyVt0xUsDlJO66mjv8t3N3jPo+59S
h2FktIWRjVBpeIqkTZQsSQU2EZ9MRGOvcS8rvPg5IuPhK6b5GHO+EZujI+wVnWmfVmNmgRwf9W2F
GU1QkawAgI2H0Cip7wzK7P5R5LwNKJ512JTYhaa6eX9PaPrdOqC6fbc5YCjlmoSznkR/AA0Y2fwD
wl1RWRysTWr10GYUWXS+nRK+qb7CnW7uY6l1HQpZq/yYhlC7g8PagpNlpUwe3lUTJgXr1CVYOYCO
o52oqaauZPiCIluUURGx4hpFZyzGLXA2TL29YkzwEb25h7u30jvHXOvZyVu9RKCRk+sQaSHmr1U0
Ahi6zduGhtF3bpFTag8jlwjTRrvWAiBAVRc/m5Q3S/D4kGfuzO4GsUCj9xjHuzmPgLow0duZ9Z0d
4O8mRHbspOh0dw4bcFTIT400cFiB1EBDanl8cEOkx3ZbtUNhZ2VFf7War3qKbtG1nKeBhJZtbY8U
Ri2qFfWr/rz7c6FdsDYExAPU/08VPnpo5ufvxMUOEehk90ZKke34JNgoipeL0K1weyDLX4SvrySd
/bFw59TpCbVq6D9ZQPnMcRyIuqJpASkroF9AN0iZ+9SQgLRKAntlNHf9VrLUQldZFqoJlXfc5dQ3
P76x/U8vrIROhbhfubj2ZYcAqvSBN+w4lbH2RykQtFOgCR7/t9I5r5Xmy2u4CB6kFlwBRZTnyP0/
uQ7Zz/MWGDsxlRyNDrIPVNomLpD9hvgXTuL6ZD31mv/qTQFMtbNSrsDFXu4O2GpNwC/HNtiHs+7c
qdbrgyO93Q21HaWIDCbqsEpURvroP8TlRn4gK2cF/BQzOkKV7fafGD+z3vL7W0dOqBgw9FPGabqb
6WQAEHWDOMXil4cJxgwdlKBCBqf+8m+jSX0dBYGw+0AGTKhbJGusfEBD/PDmvAqlDRjq1gcAInIh
fWhS9jN3ZAzrzI41qo+slI9mm1duiVkm04ePDmH51bM9MMmc+o3HzojfN7Lx4+M9GH77uaFpW1lO
7OOdwZR2gMLC0sD13fFTIlxh3cJRCPXPozAVeoWqad6hS/1GyGmktzNct9qGIhyanfVZiF2lQ3dy
aG9p87JdzxbizRzz78Kjx3sZSMWwpeTcZVUPQnunLBuEWCvXqPT/fDxeDA4n5EbTuRYGaCexKi9x
yQMmN80GozkNWoJwnfzARh/TdLg6uqwXIQi1J6RDAzRTA8/aJ14nvbcLMdE0JaEjRhwKOTzmEdqa
2j+OCXkkcwpoLltRmO02QmUYbc6oZ/EUA8girCqp4UUHQDHtg5hVOe+kWHNCh3L11dTTZh30GBy3
jn5IpF4jD82n9ZaFec7oHwzmCJ+d+uuMXSnKqxWCuLm9geRwGAyTaTt+zEZlXI7ks34ZK+HMcKD2
ODyNJhO1gERUoH9kF1m4gFbuqxyumdS1LtxFbbrfGVoHhtaelVLltfOqeBmBNUWg359QIjPse3Ds
W8TXXSJQMirqlxea2zQrqh9+fUkF8DJbmO/s5+S3RQYO4VRClVUlD3OdRrUmA0QJ7MAqf3NkkzYb
st3REZH89MNxiM2HzmWl3xdwFw0kfVTuYbaLkMtAE6pn9bYyThayBCVeoqkoUACDru0P9ceQv2sZ
D3pCw2RY1KgXkuyVqoKjpSAEiPhcAku2zUWlkiVdcmydNtFsMHBhQvmEA/MpVfhlWe7z//8DxH2j
PyZzj1wQ9fzeOT3PLQWJ5xmwghC26Q+yqmTKxZPxUw9eQk6DBmcfU+q1ZZc66T3HVpAcZI4sSrj0
AclLuLzk3ka2zK7nYjfC9e5ssOGUU3eoxp5E8V8nifPiJWReuY79wSKxlngGKjPq2m3KPkbDbB2j
pDPR5Jg4LfekjE93hGB56icVbfL0EDFTkcSLAxqSeVU3Z6UOw4hI6iesyWZ0n9+x9W3PMHUxUfaZ
5+LyZrzPQy8DGgdearFohQiHvZL+B1Ife6TTXSn+JO2gd7LA6nuP/koxFVNtbGB/QvGJJahryEzX
XP/hreeaz9fGmAtnviywuy1sOTAjed/4+tPoAdDt28H15VQmE5JcrIPw0L+ApiPcGwlohuqI36uy
e0AgnfkF5ZotqliHCho52DJIFIwfv410g3Np1s6zjrkuNHOsF/bMj7UwxUu8V7ZhcABWs2IXpl4J
xK0JZpRMFD7Tdo5FEmLw3+qiC4mN7ujVK94n6dfdaDr/KzVvccxY2A5cS9mskFELvmri/PdKhbtr
tNCGLa2pWZtNh2vRuz76cXBv58hrgkhbMf4jjvwLp2FJfnycsesBdk5Z09GHMpi98bQPqeSOwHSv
wSNOyNZ6mfbGmhcBvqEtX0csrfk+wb5wUyiLL7PKuR6j+lBYn2XV/uvx2jysjQpvUXlfl/p2GwER
3NCKpJwaybaaE70w9ExEj/+ov+zvQaHkCydNWbFSEioiEsl00wm4TXSZFzy4RPeadUNBTHVmQ+so
W8PTXToL3kafN1ylqaNikTzbI7eU//TKnxrdLZQJUz2BV2/ScB4537QSQ156GiH0OdE9WxG1KTld
xen3EJ2U7FCA6n7e0yWRPPzHvIbdx+0iDtA62MKqj/OjkrFkvTdmjWjWGKPCViI9I3GXRGjh46RU
ZVBNf96U8bost2EfkecAAEM8LrRlJ8AkZEF9bjcdBfgAULHIdl5QG7W3KdmErtr3iryBmw4bZIYP
3jLRqHOlP7hDhQ/emFzv/r8inauw3RrqtXi9uLSiepnHu96ZfP7wWpKpYCQml3GALHWZrlz4kBO/
znW/onIYixT3eNZTqJzcPCmDew13ZmlOo1rJsxQttddK7S6rlpAKAUWXLCGQj0EirwudAKG6G8io
o1c2x/73Aza/loqxMWL4BTn25UXMb2UAHlD1ATW96bBIeYrEGtijYZjwikXebd7JlHKlTfFLP15d
LRZjMc+44p5e5Nq4Jp1pZE/rd9qKGzjhXMwAdfGIINpirl0hkdbctTRnzJDqemH0KHULouuQKhbK
GPucfY7P2GKonp/Fr8YHm14g4laW+jS6HOe6SqtwWrcqJ0Wt53ZQ+JIfF2JMIfa4Fl8h/jZSXGbb
ePPz1TxCcOoM0rqkbIFE7n3Yi8MEeapLOJBwISedX6I2rMxS1K9u4zRuC4oMYfZkTjuvs7hscJUG
5mfest6rdcu17PR2PBh2IXhmkYujnmcWv89o0ftQlXICS0XhaZ4ZfA4ukYUe/Ejaof+8at01OTew
UKteN7GF+vcV3VH9AOqJmOF7UXDlDLTdwmOcEJR9NG54LGyrLC8AGEMfYmAUsPI8KZxZsUAEHEA5
8q6wKKGvLDtKIKF7q35TpDadyI9psNfzEBBE7wnUC5WboPN4cvLuWrYuEMkELqXC7wJ8Lm069050
SdDrmdKLWwL+QZmvoJuIlLL0vMqL+RqHOsT2MJ3L9cf2ZyCLGMZcfTsGR64anN+nMwZCYJsTgiam
kFQykWbOr4aTK6oxcfqur8m54gOBtv6tAiu7/EiIj6kFCpsCZafWzoIEnMqaEz/+corLor2tD+is
W4w2eIZTyNqavPLGQ67ANXuYTRqHzG0/53IGPLXG5wTnfJ+X0DGtClkSVjJOj/6ykFPP65tGbhIf
APT/SVQIEteULrf3QYyts8JBAwXbP/rcdM+Dzx3xpzL8Sa2o+xnTCkidRStepvPFbovb3YiX0X9n
KGC5YLSeBJzbOKtxZyzlktbntOjYC6USGMnFMeaZRJK5Wh+EhzC+rhuNADMcXUFNRLguwghU5m2Q
TtXyN0F7D/OuTKkDZhhJ3VZUaqHUYtaH3eV/g5JNHT4rXmxiPeCrd3A5qI/RhrQqtmNVtf00TDTv
b/TKMnV5M3bG/KfbglrybMjthsS00BU1URwkSBnBbIH6WmI+xIlLR8AcFxjBGzoQ8p+WX42Q2vtD
uknuftQTd/Ylw2tz/ZMcoukmAs8084btQFhLImE0F2+v1jvvLcIYrZBDSOg76xtr7yQd2SAF4mDw
tIYcpwoytRZEdDkMjkwkGV/spSfZcJ3x1XYLLu2zBWrdwNRUnJjZApW+9n2FZrsXq+P1br6YRmeF
YhhLxrf/CBKtrZyqNXdGgOsX5cxwqIvVoe+QycWu08jvq37PT27d8lMgO6apwg4plnSDZo3wG+aF
hmnOWOuAN+n+XlTVfM2KMVWWJJevSTSZnN794dGtjRlZr6s/IRyOjazVdwX/RaJZEZknKeQ63lnv
X26kwrbxHOqrLAUka7kZDpR9GYlLkSj0l8nnhaHQN8m7be6SpUQvv+zG/Kg8UsWAnhadiI9dAIhA
0AJhWd2upfE02zzCug4NYcgHMd/T0oGZnbwaCb6UdUgEsARJI91aNYEMhk0ftNyNmh5bj2klQ08O
vyGtOieJNG33eh2hB/P4E+7672CQV3UeNd2TwwWw6oeYgJSK9HlpBde3bscO1hWn8lusp4v+gIyr
+EGl2YnQbDJOt6UlnG1yG/Nj62pxGSIuQ96k/VygST6YI+pdKAaQq09iJmEkrbWJWuQHNmiThwpN
gwyvU5lfxEKYmpvsTV6xAmrjthVz1sqrNMCEi607gwFfWGfMtunR1RZiPBKabxGtSDVDhkEl4QJF
8uZwUfjoTS+KnuBkixbkMr6jzvfHDGiA/Yg/XL4Pj0aQbYGoaMTDMhlKv1nscqR7m7T9OIJj5Cku
fthxd+og8T5nb/T+3Uy/B/PfV7k/7/Gk5Av/6szK+O/AclYEkZ8CyXWvMd4a6KGg4r3DFDYI1UXb
5oGl8UhEPgQmtxBE8JgqTr3fJRrkr/+qr+NU74Tqc+z+wZKFB+rREvJIpK7ycWfyEDJr+IDbaLoq
XcqGOyzo3hVcGl8uNP28NgsKdSRiXB+nVaWCbc2DnBovhQrKQr7B+c9SKPPAtLiyzA2cCJ9jtv73
7O8Wql1fLUamBWUqGp+Z3nSE+6L7XBknxO43VDX4PvVifgnFMoTLvaeW+AxudmIL9ag2C9fMGRJ0
HHXMiMETjxISa2EzYfSR866kFJomkpvpEMRQZuI+gp+sxkNp7ICuCRFKn9kVVEFIv/m/7aJb3USk
OEkXDUeRX4rd6TmZHjq9An6A8oijPdPWiOj2Wfk6WRRVpMasobMlYR6XlI3whFZ5Rm7ilErsC9qK
pHynlv+b5FqgBobbZzHKSFNKQK6+rnrd275drzZkEC+et7Dj/k71IRRv77dWcq5FCK8o2F6RUwMA
ZKbbGvGgRlBuTdZrbd2u0oCR84dvoOIizXRwuL9K/fsU0myPsid88UGw+qsmVBN2QNo50cGLy23o
ZlrnbfhXAhsnbg/mz0c9rnxGd+/Gs03qfPKO9K7iTcbG2BGkOWYm9WnHrgK8+4cJI1X3lAG5BKqp
rpIMODnwEPf1MJcsn3yjFI0WOEajaxjYP+MkIS3Bl2fi3KQGOtP0V+tJD60AJl/EssVy/HpbRlYk
/+sZ4WUIxmIeTF6BBJl7jiTsAkICwIjIvGbNKDqGyr/2oSu2GvDFVO6l3VIwO0zoE5QtuMu9pWvJ
JSPGvnq8Eg4MHkPwmMOP5HUs5/RwozRMHFIGgatvEt4GhPigzASap0SxKucbAfOOe2ARVwaDESvv
Iv6VfbORMPeJT50hqyBOr40F35u6rhtp56UK2nnainMwk1qFLyfaw2hDLeFBqnGdi7HLWPfuJEAW
MoEbyIh0CbnnqI4LCVN+BT8MZKwF6R4uz6l3clODPT2T5jUtltRT/5sh77XHfsNkF1VqL4ahYRz8
LrzOqNPhEpehBkTAPSYkuZa1+8JvocrOlszesQTqKB5UZcrTbuN/vUui9XDTLbeWQU7JrhlH+Z/w
yBj08uFSTaZMOxzXCWPN+ZI6WsKMpGHCH2SAYsxp6tDrl81JLIxHHv2e3S8DdRnE75T8k8unxMHg
zg6hzEhtNpIs3qpblDP4NgogQIj2DHbmEufEDcmLOpzSb1GZM4ciUJmJlbC7M4m5GgvVwXnKFlp2
TRRXAuEvkTW9nc9MH1MdLPfr0rRjSRkTfXjRRypVSCbISw2jp/NauHLYVuxi+PISWwONgSNSYE1S
PycYYbAEJjjHVtBz3ODYXsK0nwCaPd/0PQnXHRHd4PS10whP9e1VXoFBZFqopoprx75B/vqelo0W
apxRvvB3TdCahvFPNr/iDDJItMii3h380X9zT7CJxhaLXYo+pSzTXXKvINcxHtloXYasBT+iQbup
iNRqDcu8uy18AKMCde1gRRuBmGOeyrLREm0OF8U1/90vljkne5kkNh/rrZENRWorbyjN++sUvgYI
7lQd2XTs1n0KIo57XImx6JVviPoLfDeJGD0YV0Kk61up8bnnd6hDpYMkXCSgLJZnzOXwl0y9RAd4
vb/QeH0F95WZWQj/dymRXah2dSjZT5QFD2E13gIemzrUb8fs8Dvvb84tHBYo/w9MmTdjf6cnfJI3
+l1IjCdMFE5vn2piIZK0q3b4AInX9Wrw2foyDwpiDKXW/5r2Xx47OYcOyvoEWbit/Xi5PTk0ERSQ
3B4QoaQvq5wbd8lGNhqKq5dzKrwWXo3qqQux4V/WKuNdxkYN52/iO7xC/0vYkaU31w+nR9FF8pQv
61VsMfeoAsz90tGGsWicao9oHYllsuLLxfAOk8GgS0sXRaABK82EMvOHFa6LPU1Z5ZgG4wZD/TNp
luiurrMcMfq3OT/gyYZD2NIxmiN28hl/D6+ch0t13aZ5Grsvfq8Q8YnCKzAFAhkYHiJKOff8zRGB
en1MuZ2V6bQLewP8zMqG371AoK5B8RBNtN6bMahiTeO7A6FAFbiktEmZKfN46S5/RCc2vE7cnwHC
Eqc49MrEsYAaFnvg5EtJnOtPe4pdn2JPz0DS3sLzW5Nw3N6koopWUeEY9P9IWdLOwV/DE7vKF2oB
ftOlreRtSe0N0ExHTGyfUzVus8CuLl0VkfAfUymk8jisMqGPq0Kn025Gxf+K4cq06egA7e7XImGR
FsD/pDMab8Zalh2XkCFmWuBHYvecsaBRaR3cumPVsIYEtfZAwMEYuPw8TibPSnsso8FLl9xuO6Us
SgwU2/lQmyDsFbLsfBZm4g4aaIUUVD/2amxwSJkxZrUL7+iQvETzmbZd66RuWd0Igh8/wTjfP+Gy
Qk6CYfZEziULXbtQtbDSFFl8hCW2r6MBOgKZjErWXeRcOtXzvJnkfVgauyiqUWtHebYbQ4I4klOR
Y85ChZJQ/ezpsheHd9+XIWoCWwGSsncRpAUH16tEI7cXLXiwl2fx2cClUH9YTdundIrSVUZPsUdM
M84BDzJyGO7Bid72cz1nCP5uy8kuoQoylycKiszdmzvf8iQRZcBC4HbEdrVMYww0dpaVabHgQI5D
GSklVS2RTbzlT6YWt91X8ZvtdEnwRgkXpS8YSAry00W/maWkPmWzJN0PA5MgnpfJYnzrb3eJQG4y
WC7PDOi29pM8a2Er3qZybwfO/l4ZXsp2brsBWZo5tFMzLB0lm9A7pYMrfQ5ynIK2CybVnW2oAz7B
4COpNMNhsEBgY7Yf9q6osxalkjZwzb5ZgM3XmkksL4Bjih2/Hx4dnYEoEELB8bmszZ9CnrTLHTlo
QiVJPxzeUuFS3L2ISNaSjX0+uUZdSVkQIHaKM98/4u4iZOubPGUqmXC0r1cZZE95ucYtANvpSPhi
eGEyAR+/xPvCgRiYA6RKvwtnROqevOSivcFwf37yBHr1hRxnesRfFlaP7S6cufxYwadXZJc7hPA+
kgjilUhb3J5YPHYk5C1lADyhyxIeCZcdX1zHfIZLBt3JP626l65Y1uReZl0zFqNSuU/3iGqME/Mm
UV7vZ1NRgDdiz8ZpZf6qXd3OXEra+CIVcEgtf0Ig7ohZ2vhUnUSvh+xF0C8h+wKa3eJgEh6QSde/
bIaK0dZXI152f91055PF/89Q1sluNdX+Ns+FR6JyA5tFkD06nYs/Oym1yEG1FAVjr/i99R796ZN/
mG7M7N23OSxLgUDbUmaAjgCrvv4HE0LkR3aFXRh3shWBb96RDmhMQy72pfbJ9MYoCKvyxg6izl+S
SjZMr2eId3afIbm1jy5OZ7hj7633u4Es/2BlGPpNO9auD0rd4bhuLXCbejtv5RS9neSQKx65UGgL
r7OFd6dzXF7J8+8rOVoLc608L1is0rDtpojmr6JwhDstn2MTDj2RFDuHbGqwp+Qr8UE/xW2SdeuK
wZ5NWiC2KHC0Pk6r/Sa3Pm2Px7UkQfX/oMXZR7XJRxjFlEld21Yuwi1w3lPp+IAVRZxDZWpEdrx1
gKzCBVs2b1qN2AGSd0oO1kAAmSGKIzqOFGZCY/EAv/vY00BHqVSyeJ7lOp+5T/XLmfI0/QPdRA9y
wVNv+ZHSGMRvR2x/QUzZb+9MVsdwj3WN94EVTiCFDzACxz0+kx4wkD34o/hAJPfBRVD+5JTjGPTZ
nWWLmkTSp+iLW3x9Bf9D0wJojvr0Hu1BwfmWt4BI9/WGHgq9QbEujJG1Yn8TbVFtU1NdDw/NL7P1
UB1o7QlBlXQ/QuQ/6UULss0+LzQMvJKVCe9S4ANW9rTy674JhUaka+reUi0mchuePNGuDFipfgNW
sUUdcgIcUhsymalmtBYYguol8+Dzcqn7CjsyI6hZBSN6hOu3k0Lh1ID0k8YJD9y4H4QCjQMOLJ2c
mbY5jKP50L1TICczmiFuaefcPe/fhNapeyvKOCc84RCgfzeA1LwNMg1ubadrekBMxgWLx+sgn+jQ
uv7093cZtlwsumZ0VG4OlwCBWZ27S2PgoWc4+BUkoZolO4UPhvLEMbI7ZOWNr//VM8MhqieCxf/S
b0WW+2c46aJPfeuZLxq7tdmJPmyAwun9TVqxIzAaE/PAhRaEaO+KuBk193Cp6S5ACS6FqkWMPbMc
bjyTiQO0SiALfQPTiQ4ZAAkvl0epYLghkV1Gv8Mfm16OeFgBSJwKy0zKkKoNseptEm5mxJ8yLtRl
oEJefatBSaCY9Nsyp8F6MCGX64NvRU7PHRcZX9nbd4bjXG0uACRY/qBBqTPg2N8EYqJKBAcgVclF
aFH8Kbu26b2N6obYLZrQFfrxvoGaxO7OAZSxv0BtSxnHpWG4QxsHK8CJaUVXpXhvyZkCIkPJy8Xe
jhM0hqRdNp1doORetKc7euEwf7e95oEPXyYcnWkfvc6b82dYdTfEPC9Qta2Q2Ct1IYpoSvcCSWlH
rOdGRkK4ZJhXBjuiYZC55RY/kySxPZUONIA0s1WyWy/8L6ox2TrfxumGmw+MVg/X8aGgz1P5Jrrz
8j1A/TdrmgcBDXd+STd1XPfm5gWabAQkyqcJbXf1vVzbwRimrcbn6XIt638zzgxAfEBKqWNfkpa3
NotlDtx+IWn5T3/UlorPgvBABOl21jaRI07q45lpUVvwjgby6CgwCqX1atdAbEbAtZyQ4wJBenye
ajWnKx40RFPPPULHNIXQawTxciJ6vf66v4Drhb7PgHNrsYw9f6R69kd8Lm/ouHF6fbfIgdGoM04o
lxvHU3ym+BMOl0PYLCM7TaZ7xu0BGN/3yZhne1/cgMfnlRfldOrvP03BOKMl2EGLZlFQ69Qt0n+i
SfAo8KC+hnIX6nrkyKIxp+RPiQC7Ofiu14nGlAvNCl7MKAWweI+irUsNnCptNeyUbRgwbTnokWow
HIQxS84oJdywnYS+asWppm2lY+CfsFtsAYJAmMBKf4Xi7OF6ckM3wgB4Mb/xRk78kCvZkm8ey2Rk
fMrSJc06LZvnIfb/7XeBJD4CAKVDtN1LHE5IRA4rgiuv9PL2Hiqxb8mBIIa5lpMZ1hlW9K/iXOhs
HuwfuMuAdrWk5KbFQSmFVxkhl7G1afaUefvX1kW+AWovlocS8MyqgiA91u07T2dV/Q7E0GSmOF7p
lNrV/IqKLzGtTp/73U7XdklnwQ9ZvvA40aRm9Vlj2JgCRpouzPgnu6H//Zb1UO3w2O6JtdcW+lLy
fHbiR88H1MM6RlcKxY/FiXo3hU+umvP1HIOGwiyNgHgTmRNeNv2TCiZ+23sOELwQrQRBvFwAGVVH
DOGcVRNL6mSGKxRADUZqOmysIrVwlkA1xbf6GO+hY1zu1/jcP2X5lDGLfYKgsZkze6xL3qqJHo8A
ogvufUqXoK+J+PIHRTuGdJVJMuCHIh+4febNtkmZ/DuYYZ/CGGDwdTrBqbhnrIExZolI+POTDWeu
LWYIvjqLUAm06dTnW1Z/b2oFfBlwUvBO61Cwsb9G+BdFuNQDGSVMqqcOa9/RbjkaqVgJhay4XDm4
7Wa5wZy8H8JWC91oCCyiZvVwEVOAWVPRvbcIEUG1UbGaNdDwRTTXPoH44VcrV9i20C/+ViBR0cgA
ZE0Sp2jGO4Y4nBes79GguI8WA2IIutu1jhRmu1qImGO7jBZYuSYA6rfXyfRe4yAH4s2o5r8i2+Nl
aoy7a8j8OfAuyl2YTTqo1VelweqAygGaQ4xJaEhLqtJoBaodZeY4xpAbPWlkhv+Cc41A+Yi4FdYI
xBMkAp4HvhXgOJiPEkoc1t/tpyi4eo6yvMiiCsTmeWotEbFdw9CNNrYzCBP54IVKLds13uI7jWMQ
6MphOnoxLjSWYQ9uavHWMU1mFMfVGXwUUPbwwZQhJ+R8W/JQ/K0MfSo9l/KyozbABhGaoYL4B4c0
hdt7ViqQX35emdsMUioOTTKa1dZE8Sepq1BtTfSocI7mBEtgNvYwG8ikvimTiyFAPGWl/H+ViYAz
d8fWf64FStzzS7KU1eysfbgRwQq9pYgCGNkCOkvKyHFIauRlIZEsmG1Cb0OcvatThxra3PzFRmKR
IYo6QzRnIQgPgGDHknhdbvTRHcZ3I4Bol68bjyApkPa9hWTaM28OKW/moQNhBAKKq4gEKd83fYNC
PN7Hdm92TBB0sPP5u7yzP69n6Wlk63a1hNH/ICoz46bHch9tXo3vnlZU6S2dqBQzsoQzGYAifkz1
Aq9OpgUVUjnEZ6l6hhLfNiN75VitKoicN10z3rFxbg07llwdi79Ps9+//undTv8X0IRPC1Pye1x2
e8Z39bv9p+RL39qJuiUnxeaYHjOgge9FVXm6FDksA7U2iIIH6POXKVX5tL1s74QdLVbpkbnFwQ8Z
JGu9SkNw3E9uvnqsj6/5bJt7FBMAM6HLYymK4zEjrjyxlqvHyclLvckUQajmLagwcU1xixDvn4HB
tExvz66NI+o5/Z1PnrXeb9NDGcEY5Sv4ozLBiaJJy2ilVCz9aReK/34mwTisEc1IPKoz+kkvPmOQ
qp/EzUofidc2OtPae3rypSBzuK8XC+VyqZWLhVmJfbbsDe0hWT2Dog2Gp+nyyaNwxzghefw201wV
kF3jmclEta8k3yIEhjfrFR3z8eep+KYgozWgeDjHaIVzSRWjn4pt58CxvoUFO/SpXbWu2KJYULTM
bI7NaZDId9NcSQiKd8LBt/9uRNbYft53sCLVY26Hn23QDFoxusXv1rnuuBU3BheA4uu3DQuQqz98
CH8FdChU0FRMT7vyo169oJnzNl18OTKLo2H3em8xJ5KbTR/GR/eB5gZY6+ViIgvtmo8ND7+tyshb
bdk6DO0AQ2DRUjKcRVXDCYEG8PXh2oJHNyMgSXq+MNc+MG95t2Ry8ddrWDhfNq2CPLHHj0HOK2IX
H+MCv0taJZNvlonNOlaQAFhpCst78sSLUpMyHuWJzqVUR0PWNSEvq2Pm2K6y/kWpqlfThL+KFq5v
ib4yBDUNdl34ipzSdO9qO3z6BZ6NwaLQjbssc2+M/4VwwddBOCvW1H7U7s9oZz9j51CNeEE16nvO
tE27Qo9ElDn32+a8qrrxMN8DtTdwWTG6rIP5zJpOJj4jhEsungihgZp8GxKh4FNWZcdI/isOr9ph
ra6glgUFrdfFAVtH6BslDhZaYWVZYgo9nkRSZb0k6s17skW5qQVaQ6KHlVZ9Vw0rBJoOqKHLP8+U
FVqWc89Wj4Pcd6JWJ7i7lDfV9P9O68gl38H7rN18wY9hSdHJVKej/B4pXDghppYprmcOBNFqI46U
xrHvwWU75avAEoTeMi8jBbpBfQL5VKSiL3bTlA+HwsEc1ogJ9ZeLO8xwzTDgXSmT+wIBG+dWRgnI
mUePGyyirTeWfCcm2994D58t2k7Sh26gFGt+54VT06fwQuvtDgvDip4lVTGekTu7Lo8bum9crB8M
rLwbGab3PcpbIOoVmWeeX7MvSo18gUZ1i2BLrdNkdrAaGc2ZXAXYsBO1e02rGegnKfZCF3ZxSs+D
wl24VpQXxUZRnNFFiTDKt8UdQ626n9rK11YGrLm6+vTmffWCWCLE1KbEs3L3YvJ3aGbJ+aKd3w4G
R2y26OGbr5suiCJt9fU24qByHnrIFYLjRtow59DfABPMV6D1OULfuJiyuH9reEWNJrJaPlr01WjX
0Nf2PwdToKeWVaJeOvFyC/4wR/E7aXhJS8pDSBAnJx0DK6ldPFFlyvu0OBtveWU5mdjTDlZkNfYV
DSMVMX3R93EQ5dnzFh23wtkuE89WurYDYyj+uAaOoYuAwFcMlvDUuzB/SjNYNkoRtdXiaSYGcyiL
C/ihPshaQZR/pdLkVn9IzRBIEzLWdbx8HqJgdhNzkAQXbjsVGviILmfTdcPXkJacLfxr+x8kWVO8
z8EsDqg11g0RgKD3bh71HlaBq3RBke0mBeuBX6CElWYNkVR56XkQgqFpM7idOPGCB8lfuu7RtUMk
sRdWNcGHxPH/9O5DL0WJppdSviTUXAyP9mA1ws1lgdT5sZhqznxF0K99FGfKquaU3GBk3E7iKBoV
FnxkfdEanFat40AmBE371+5Ugdt4ph643UTEg7xhgZdXedLwvlAxAv5/CxIyqaJ1IFsvDmLrW9Sy
Nu91ZZ0+2V171eb05l3e5kKdKSRXEqiDEoSZvHXHQ1tgP62CmlA08N7t7CMbdhSeIxe90QUSTlUF
D6Vanx5RaqwHsaWbH5KehF0DETZ0SNST5M/GJCaxc2mGoQeLKqJhP5NMvi+HoyATAXcF+3hOwQrv
9zvgb4UBFeKbRrWqPc1+QhGCbQXtlTtTIdzXpvT0gTPxIU8CeSEqrBxEakhhemd6vYcHjftozLXe
Yr5SjxKTs14cuLUli9EWzJATelu6y6faGIVAT8DRqvaeSoIBKdQZhUxItR3YNlnFJY08bzEWWx1C
3ASitAALfNi2pQZoMiEb4NN97VA52qfNnnRsXHd0+ai1j20iv4sqlvDF9+gskg7fH/Gs5fwEJX2U
WR6tzCbTnQFAk9HRyfmXM9Ul1cAjb1X4wQfmrq/latI8bsLI9veDWf8ui+2IknySfoP/lwCJZWnl
E58+k9qs5xdA4lvOXZq4y2jTO9llJAa+ighzyzzIt+IBuDtQuYqooAz/KtPpR0dKFIH6Mx17TguL
KeuuOJNjkIo/5KGG3/4albKIEAX+s6LtANgnvQc1oKPZVodjwHrFS88/uOS0yJhXR12zqx55hGix
oTN9nE1IAMnQkgShnhW5LUGQWE7S749jRraBdt/V3P3m2XfXsmK6gQtNSXTUk9ioVtTz/bk+Ya6s
EfrrOIP1bCoqJ9j7m29TyYJpr+HDP1SRXirg+c3ci20K3O9lsEXerbMC1oHUjWPhifwkqZ1tB8rM
nlmjSBiDpWC9YFLdsUd86XU4E93qPwE/ua6JVW+Za/kvMFA4DOX+yi08MWzHMDW4sHLxX90x4g27
kKJaY6s3yyy5G9LerOLlDLB4Onz23mNhL2apjSamU1FURK5FWtRTWc/LBWw9M4K+yIRtHfNIhiFR
LyWBjRpeO9cSXlT/rjCefAQD3i1qsNJmo+vAgBGOCqm1YhGI1glszKQOQU44lMPXsi9b0BH2Wztm
50Gsgsu8LLO2LWRwVZTEMqWmPdxYpK5UYZiWSOZQOfhmlm4XTM0nxttXH6MmzTSRaTsDSZCXg7A8
CwjcJ4pAKw8M2oLSxOH5KwsXEhAx+x5L+QU+7wjufXRXSeLsmHIx9HC9IPY1IjaQPJIs7pDE1zX3
5PU7QrUKsDtS294/8rpW77gmoAdlWvJpTWEY5gz45WCejN6sO6d1QQdGp57mO1kbpa7+7nz1aVkM
iAXUa5RI83WEUrykcITt0lnmkMR0wI3INidPcvh96g6qzZfXwIgZ7CR0QJJ5mbYgtLByXQ8Rhtzv
URp75kOT5bxNjruU++xxf23oD47VeRLcDTI1jV3K5UC9LUyEi101vvcutyL6DLTLf1cR9tBi29U1
Nitd/LxaKLCPbUWErPsOH/zAGcRJ5ucK0iFhwSiFlroqPFnkNaNLAH63wzceJn7QMEojC233NmSZ
wQV6hlKED55trCWw12YuV+QJTK9+imCVbZ+0NiZctEO/7usG34MKVHWn9hekfMwJCkbIroVGSUNs
OWEAz2nK4SYLEjTrQh48+UASguGOXxY+Wlv01xJQSEMmZK/lhsfF7EXieZ+pK+POyY5P2/03uYgk
83YO/rLl2MJUDL7WWMOkpitx3zQMT9WEaPYvamii4Xb0NMdDwmhA7lGXlNwMajO569UYM7ycfVa+
coTJvQFMrZBBZr4fKFTPDVqmuKK0j+y08gtViIzLCFxwxkh3BmbVSwNWD4RmaxiPebvE29efAiqq
U7h58xStokD/m2ChkRv+1HCz0bVE/gNrx09d2fsKCsrZc7Z183okdeRRxntHC2GlKPdX+kRD1+r7
yXoei7I9R7MgjSZpI7of7G08Rcc/9zSrviMrDfKC+6URY2MWe09ocG/oR2Oj+2AEwYyDcp5iMsyh
28OTeiuv13qLuBJHHS7lO9pS7a5JVPVPQ0I0UzZ6EiuI0kBZGvFbtLHZ4HuyJm57PasqQQDGcxDF
4sOxBHzFMYpoZSrV2+sHsnqwzua/g8m+R3UC21c3hPXN3U8iJZFWPdgUEq2rArV6es/bY7pwU84M
qW8R6P75z2nPON62j13JQ2H3kF5ouO+c55XUI3RNNLl7mUYo8NQpF0bdyfWst/fa9p4TX0y4gA+j
htPE4lGm/izR799770IX2yQ96uhESJg3pkB5xVvGsBdlOB1V/9x+2/CNlpscAuRhGEqIZRXhhHzy
43dj3P6hI81Wblbgl1+OrtXqAn82as9HzfJk2QOk8BRCYZxFMs5ASz5b4Zof7xKvN34xB5hbIw3R
oFCkZLJYmg2inJv5thEQBFGzF666fdNAMLwPz2V0Ec5VgB784Y2+lxsBBtRjuVJKm+uhv2xzeJA0
m0wLYHQwxMzUBGlgc8LnVWLeVa83s7Th4YJglPmtsaImzFm0wS9z2aqrRcdPoCjqSqsnuON0eXO6
l4NKCfqkTFhdMoyqG8rPF6x8catBpaaUK4JJIQDUpG6Iy0gBQ+PL7vng6Zlz7ZMsto1cFztMuJNz
1LQVHWbpAddv6S7tzWohYM9VwVM5yik270pU74GokrS78DrcqMzpXrdHLeIOiunB5EAzDhH8nYER
PILZyd8ieCYmybIuxdmunBzt4Vxf9OQyVtceo+yUWdGBqerq8N2M36zzXlX9V/cS15G0TmjoWHcW
2NMQ+DYTRh2sBGwMPIVVBoXhbJjUHp60HcVtXNlqMR0BxCgFu0JD8FmUh+54UYq4i/Kdaash3VaE
s7WdiyiKM63wo/Roj5mzzaIkHkP8P8/DgjzHYRV0Fvua1jV/n4Z98FuTSCodswQgTZEzAVzinccz
F3MNe2ejP/sp05Syka9ET7DtaqlVeeOIx+9aQYwmx3OmXlyRfdsjNclgwyHRWmUl+RwG8/EITq4A
bRkYg5MSsUj4JzAV8MFmB+yE4Ihpd48IjBb0Q2jqycN3VdJeTQeZw30f1/hiemE31D6A6Ws+k0RX
zfaz/y2dWyCz22bAimfRXWFvf9XGIJxdx9xXAHATwDMzn5SEZxDnYP//pRHi14xy5dFMOLyOntjp
LCWRRK9zfBmeRud9ultoZmXK44DL7nv5S/UheS9LVZsVnEoh/x2eTZGDQRY+GQOcN2AwY8LtSfxh
BmMfZOiD9KA/6RQuP3oclEDWDoZ5cAlGlP6pDCwpWiB5FOwNQFX0FZRuA6wocq5FXm1iEShjP1h0
U3Ob63klr4DCB0k4vZQ8+v65muS3gV2oK3GfCm9NgRqVar/NGgyzkKSFzFm+UevuVABw0bSSHaxR
B8EwOHckvzSApMtN7lcAQxgZd/7pflJ/ApaPi8PctxvT/2Kwe8ZCenXjMALZh3W+N3Ja/DgRPH2l
DUfDJCka8gdBrzVkIOiPIUtdAzdktqYansBZAH25cqqkv+Q3w2OIpywsNpdv+Kl8xafz9PGR5Es+
NdKDQAkST94/y3l56Xqnn/83Tze/jGkTQk2IupjRaJ2/kY1OhT1uXwF/ECg0ySrzCoEY9VuYLQ8G
gFP2/pfbOEX3rerQtV3M8+GKlZtINQgUTsQQ2yYj6Q4vPRyZFgXaaUXvDLpQTYBwgr08v1ZJztQo
TY8tFCir1qJGeMO2HnetLVF9Oaub5GXXnnkGlf8v6ssPtrBPLa0J8unE48rqWPtsQL2Ufmcq2Pkk
Wrh3XYiStKyeibCrLk5wuS3XMq281gx6GIaWxOIy55kU4ZYeCHcoeNHS2Hd2dFBCwFlsbigAvCab
H/9oBTwKWWjWEv6EGnhzfNoB+9dcKbQMHg0c+GKhpyAcNO+29ceGPdN/4ZR047jqeFOWMMEeTFM+
y/DstzPtVtpqXLcCeEJa2lchkkifDT2mV+OwdcRmtC+ylNl1cfYJx3tbUkLNH30/mCXNzmFQjo+P
2mu6NMSEk42W0ZYxk8bbYWy1y06wbazAOrHkeDxt+Wu4hfNdMlCzI/vUYWW20MQc3WM0nlGI7HXG
iMkdidRj6DdbrI84uwedmO4Zw4y4cA7TWzsTguGJxHX4KksUjS109OaCH2c1CfuxW1bGsP8o7v+J
XgTL8jQiwgskSyIMfutwqLn0vSR4y19I6hmBOp+W7KTl0kEGQD0OUlSNdUJELdbS2E37fqq8vJOW
1DTkpuhuJEZBL7Fx6TnWQnEHkSHfzU8RGD0wzI4ouDCKqP21wL7eZC5Ns6jkPEuHqowpCoDuWXfO
TTLTYSlG6aaYpVyQ5YPFpVW7jfv4C3CHZ78B04lDJ8mV9/onN3DQ0pJ4VLT4pQWoS7nJau8A4oCx
VxQhsEN8nZ0Z04V+olnr83y2yTCPqsE6qYtlTZV/ZoWhDufwF5Y60AxaXrHgStWVgecn6JRNwOy0
ye7jq9wLSe35oI8yX6qg+3X/TUQwLeaUsZqZIsbidszzCkWytHWs2k+Acpi+MC/tC/hzaTZEz3fy
Xu1AvUKspbhW16vEAM2zh/vSGOctOQRjSH3E98zfJC9YOAQA4oGfjHNAGP5clzyaLncXP1CHfILZ
9Pwvo/JB+uMmuFbr3fDXWwsL+brOr5KxvheDBAjqGVgaSbpkeDaxGXPbh8bDNAIFrmYd1DSUz+40
fn+f6jF76h2IX/nUqmn4nX4cRGYTw5ONumHxfh5tN9G/2ivqqh4PPboNUycN1i2TyDBomkWEhliV
7UZEnSifXWuPVSf/uIisXNeNrF7899nHxmRT9XIlp+6d9KAQKBfBkuW0BaPakuVd7nZpY/Ka0eih
mUrr7FzF3pfehd00fAeNeHY1rIfV8b5l81LWeUMvFBbzBTtpKArLwqaDZYSV1AdqtRwVC7Hd1qKK
T9lYRJILrnKhkVfwHQULzGSCbvRHxlXW8I6YVmpOqv0MlgY9L5JbSr/vKzW/xUvBamK77JXhaaj4
mR1yY65LT1wFdGixOkFy6Tf4vJf17vKJvz/nOuQvSI434vxtIp3nug4iurr5ETSHhuC0c4hr+kVS
lNL146PpfaWb3CctBq8bx+LptmExU3JNORnFPAqzelz1xzw33lFSik+oKuJSNMyIYCZbyewMq6RU
tE9Uog0qfrKCanR9PSSM5YAjpIfgLL3/5Cgrit/FqtdGBZFSVGFb9s9QpyudAksBw8a2CSv8oN5M
OPxDN3AgpsdZFkpQ/Z78Wr1tElDQbPk5elxmctpbKW5JWfxAZ7AwSKDbkC6eSUmvuRby+S15HhyB
nHiCffw1x68cIWOGTMvGcczYhMT8GU97os63Cu32RIByVJV5BSkkKtgSux/51q3fnY6P8DuWJCQK
Ne1ZqkPdJR+R3Es/v5V5RgvlDIDz444oDSVF51JBUxIj+SR5M1kfjC9MtUuQIslIiYZRmu58RNuT
iPoIzltNdF9MF6l3rz8x8dFslZOwsrxrInyP+1PkMllZGxfj63MpYZLtkdS/Ye57AJQ/9YrpBRnA
8GEAXesAqFoIVsSSIYQPZ6+X6R6U5BZvi8LFyZnn4Y3BlE+A0UNhMK7kjkMaDCGvH8okMPxGbZLl
OoMLNdhozlIgInAsJUKgHCVpauW+Kj/EelLccOAg1aUY6+Ly7Ol01EDNx552W+pETj6bo9wo2nvf
0SvmGbV2PiR4z9Q7+PO5Ep5ku6W6EqPdPuBvNq43Sk9af8cyCoCo1wKqGpYOY2umuR9SZ2Ig8kvj
R3Lq0f4+BGt3Uxkpec4OzOZENGvr/QriAnOzrlLLdk6Iy3QHwcHG4gsiCcDNnEOdDoe7i32LjtU2
beXO+SJz+Eh+Zcs0te6ZItWTBb5X4y1J9H7vnWGBpO2xtwbqa89BcQS/ImXUfdiSc9qZQQyl8TzM
nFj48d2zb2ffB6wtllYZVujvn3g6uvYI6I5vIO+pbzezZsZ4BcIW29sclea2s99bmC+s0CgEdHDR
ZZfg80Dhws6Aw4iX5x/vj/iJHiSo7DIJ80P+CZlmUx3wo2DG5yqBUI1dh9iwh6iRtk4Y37zr36Pz
/tfIEYVeB4KP9eMyvZgXSQCsy8u0p/lor/XRZnMVNRjcdZw/lK59BUXhUw1zR6E6JtsS8UH610W7
evaHClUE7uIRf8WqY9rUIDPs5auguicATteTvwE8GJGC4l38ku70fDtGYJBWEjM9A5NHFREsOSRW
s48FjRd7PguPCeAdLvSU0WOnMr44p61q5wp6J9hhhujPFhcet7pjfWzHKzE+49z/7cp5kxQnU5tB
wxweHNnESaoVzeBfKuTJ3Gk+jwVrtI9DPsdVv4+BuSHxWy6G3kw+2CU4OSiaghyx+ghtosUyIbfX
dPAgMSZZ6idmmr/mbOm+oWW0zKR1Orjxd4F7Bu/+DZtXJrsOW/RpkdDGkU/sWpsxDoWoH/qXow6r
z/he4v1ngaUHtUUx7odTnb8lCMX06a/9zCcEH29Y/t+i189hoVaZwDv4LozTVSV9H6ZTMDio+6xH
hzqk+K+qIavSdAKZwH92xaOZNyaLnjhVcksgjisJaGnNOdjaYvIZV64tchJtjsmweXVCdx/qnMMR
nKe2NfAL/4f4YQUA9vVDcc+kAj98Yz7K7UZu4Kf9j08ctTDKQ+4Qj2PQ/Zha226eY0IOTXfERmMJ
xur/AAV6P56hpIUVF4+vSCgneaQo4Eqi9cnw9GMl15ARazgBuOh9bVKETaa5jEeRSkgZB2GOqHZN
1NlEVV1DyQsXpgwa4OH32kJGfrT0PZwEVu3s3kc41H6ubIkUI/UH5UYRNS8qk1tj/u1w/QlWU1aE
oHr7Oub6WkqnGkGLpz8c7uJp4qgcKKynhB+fLp7uzKSB4X4yDD1KLfbmPDvKo8YEdY0qMRxso7EK
WZqFISe7GJGYoIuHNjRgQUxopuan66QD9yfndmqxD8ZevQJZRksNAKZkc2uoyjyX33bYaXEZkN1r
FoS2Wr4/utJN57NMx5VRrGh7lmVVYovp0fJCI914v1H8h6c6Bwpd1zADnqi14pSyN1DnVB/j6w8/
/Xg+iWvmepbrLI5cxSjjjqbf6NG/cN3GCTC5oEaZwZ1mG1EwokjsnYFdQpHtcEdWvcfipGEME22P
LIFyfLVLhKb+i7t2zovEaDoqXSSd8IPBZ7yYarJPTNYkFTfEyCZOdL2lIQSvcewVf/5oOxkjLGue
W/QDgvkzoRVVzUikxOfdqB+QMh7ClZR+9ueF/FWjQEJkyFj68/Qa/4H9lKlqhpKvSHVu0r3sgz4k
ehoVtfNgKVAbUswSosdc68KCuS/DYMFdWZJjUXPP5wWxCr4EXiS+6f31bUh+aa70cDa8t1KpJY13
ls8UeMaVm3PesKJQPsW7zJvCjJcwmsazAI2eObKy7m6qffBoC2S1m3avRd6BUSq6riibmRTG0dvW
7hk5CXoUnESfzu4iqp7cQOwgMu++ROBV1DC5VqhORoqg6byoX+FhQ4rTiMU757/Gw6rXFcm/TNWt
zzrcP/GYRTA2UnP+kSXJNW1ZCCOYzZdbtxiGMR3lJjnLMAziO/QMnlRSBVxD6VGoFycZXlqedTDO
dwcgeg+eQQhgANwISQAF+a8NLfH0zamrGGd5GFreIBM32NTW6tvzVpJPi9AsNGYpChc3PqKNOt9X
VPtZavr9ggp2BnJrVd1aiCNn+r9hU76N3xCmMpDg1/1zaEXVoEVZ6pVbpqClanat+D14SCzrOulS
1yz5irDtI+X1vvkpbiKUFya/oLzzYH8wy12HZV8P5eJXN5sLO3q9rrm0tc2k2kg0nvB91AvtNiEz
iIgsFgrG8ZdSmzkC/WdjvfGB7mrB3OJLnOOO2v8pelX1YeBWHgYFkSyu8LrQKlSfsBGIdHfDqJ+l
6WmtXNnS63ODqnxsQp1dzrNkHyzjiBN13gX5ZbzRFY8zdy1uYFLsAhq+p9xBDzZ4X4Fb/VDAee9v
VsQhvxXGZHT+MBzQT3SW3Y5PPBWTY7h/YP0dKnE45Cy7PECuIqQknJM3Srl2lJCruuMfM1vV8diT
QFk7gcuEZcFUUeVO9N6keZbztldKSdnAJJLAtrN05iLVuDHZz+JmWQIesMiV7FFUVX2R/DGCh/PF
mwmAGd9ekdFYv2gekeGstsTMwWef9hn4egNBwZjz3eUhiM1WVJ0uJ9m9s88boXSKhJiXVmQ0vcFP
imiyYQ+7tORc75W4LnmlK7JBmD6gmu95oKCD7DrXh80Cv7TfjJojGEiXL1pEOdDIzYxepVuobj7Z
1lGL/icIEd+5hoefZbY+W8NtT2sb2zjXfmWDzWDVPWUhspcdJgXdZ9tKvbgs0WcCbebpH7VORFa9
OFCZTkXx7BRINeKonBYJOjG8+XXDtAlsgm/KYmgwIjXm+FjmMZPQs3sgFhzCFHM2YHTHYza0Gr0j
+GSWCoeJYzToi7IU4cWRtNs4Iv/yZwY2p07nPpPSUxe7gZcvb7RVM25FjyqFYEFVifrDNPfIJZRz
D33irfDLTUk37LQkjJgFlGzXKVCGO6YPBqUw+herO6cTaKw9ZCeYnM3URW1NkkrHGo4q/UZIjjbw
zYMBasrzpEF+bcFLhkpIZhAFETNbggHsRzQhstKR5YOqh5heyfUiz0h+briSPL3xmyzpbaD+Bcgf
0h78+qt0HElqzweViwpy6i15hJpWWHt0myfHlLdBLijLY4iCFD+YrXNhhxo03QIM2VnBtwJEOKOZ
8wdqu9bczkIb0TX5ZpKq/l/DWwixBtdsFDC0CvO+gtJCVRXzXhIkSlaUYyMkUgUaaxkCZGzkb/63
TB4qF76csqwWlqQqzugddxWIAFICcz3JbBPt5PpV0A20B/P7MNgOsvyAjlvq92r+fWR746U6jCu3
aLEr7CFGoGezPiVsU2k1+Q6dRCXibFggtv19zzQAOXT66/T2uv3sfVZu80ry8zjbsmrvJGP5pfFQ
rZNB4Ntp22u+Tk/gyIzeuFiB/5lQGkHz5EpUf+Eh77AAT1fDsnE7UqV8706hbaHdqMWHG5TVcH0c
CijsqpGpVGZ1Xin20hV2Phxs7jR/NpJtEllvpkXwkDQ+IDmC/mdkPkjQFOcJyaJjfyn9TePBtkL3
WU4H9wQkK5LC40v/5Acu3ej2BVAXyScat6fMmOgcaHyIGnkN+/NcNxhzVxkyMyia97nh/MEj8DEQ
PpTbWxrdNuH/dP5lreCy2qDOiZKA51KYAR/i7tZtj8C4m0mXWaKjlufxgpNMevI5tBLs/ww9u9J1
VroPBmlr16vMREgAq8JLvFdx1ICPM2H6yxSrVnS5vEVBYfbY6SvCeThO9Ti5UDJJVueusMVRQrRT
ZcUjBnme5hI7Ep+5WWX7J0Gz0oKjZ46PuHQoANNjEQ5bktuUDB4NOPMloD5HYaubXMiDPGUecskF
aWNuRzx3FNcKRpjqznPYwBL4apBgu7nyvcAsMpbm1pWaa17egnFP3QCxvfUWnrhn80WJNsHVZN60
kOofFNl6uNrQtbNET6kLHBl4PzPEAyf1AGVGyXL1ZKVuMGiZc8R+00q9cIFx93ZQUUYVS8z8H0kL
LauhG7tWw/BuQCoINhoWybQEM9/BMaNihjdbs/P7cDs9J79bQTQggtHCJwKO8rlMmg40uR/l90DG
dRwBMeHzl7LZq9oC6lObkgpfoR1WAQOdnF09rNPcxcNH9yhfLmQlT0tKInZzI7EGQ8qBLIaB+33r
7zJk+wB3Z1XcqYBKuyMXl1DOTYzL0phYwfJdXfGgDE1EFHLM+Y7rsoGuw8+zsFH1RDof6LvkwWJp
pJTUqQXDjv/vjD3/159IM5hGbXh7QmC6ndgv9c6wWaefjnOwUoJlCszB/AFPNGGIf0zEA/wgkKz1
17Drp97BNJZHrqvTycvGlLoUL6oZwiQ1anhIuYmYZsgOBsKkPmD6J7N1iS8GufUSW7g/gKjO8yQV
DYY3smAQWeprmBF+doLaIqQHC8vdPdd0qIsX3lhQrvgeGn0RDrUIiVy/O810H4zj5LV7E9VIm5+n
u0bz/wm+4nqBXuSQmyXMSx0jsSCyfZTueHOh+28O4OKazR7oZaTxSa3letoRne2MXRtPwjFDSm+d
yYL54uYNG4txr/BfJj/xOE1rSGGyPTdrHHIZeoIByQ+J8yXK8t//ghajaIV7vM+KeH9LVDKXyWE0
DxXXsgBOkF96wJYS7tjO0GJoyP9scUE2z4CRn8R8sSdLFIwdzvql0H1NbMea0EG1B9OLcKEji/BK
lXhwiokuXmn12DxawMjFGnzpBqK27nZr7cGZuFv+bbPd9bR54Fhzc/aEQ77E0QCOAEkezA0/ie4d
J2EGtNNk6T4M0M7vQTz4D9SOnd+kJZTd433+RXrQIfi6RLHVy9furAoLK1ANoE/V+RCCLYRnm1+y
xFT9AAUP+9juZ3/1vWnpRj7dU4vRs8JrjIbfyUM4RDdQmx7+9sX+W8W6/kT/c3UFgCnZB2pv63pf
hcUdVxmRX3+ziDLnCeTRM5mYTNt9i1LDRakTpgxl7v3PTbNwWXON9gXC/ra30kKo7c+8yuLXHKzI
PUspqdvL0NEjDNV6dn/OSHT9EytNuKaz5qiaJ7ZKH39V6HNeqB/HCUh6DRprDe1i5+DyZKE0n/B7
k2WXoMLHnyshCuXURSK9qYsJEw+oDcmHGMPesLGPEPsvQPtXrQGMbyY3GhMTH6DY5WqRHqYElyp8
xlETrexGWU8UkyaXgdyKjRlRxUHsg+iN1CNR8DXWgvfmToJedcvFqaRU9JfSFMV66ykVqGnnor6Z
wrCF3Q+oz/zvSpTw/UJuUZiLvGjwh/CO296e3fApEYW68YAcj/8xgFPtKFKod0nmOYgwv/i9NP0F
aqC7TDLTOMk3IMLqpGYOvhTPP7of8z4w+jmaKVd0Au4nGn046IkPTEA22JNoLVrMrem9eb3fYr6G
NDsxfcqXO+injQzt//5SJwIUK9bfT6SDG0z0mz3T+i6qiJi1njUAAvTIosCfJJ+ABhJZhnJAnciC
wQFEycdDJ32qmSecMiZBtjcv9HGrrsz1+9YzDE/3mb1egP2GW8eYGdSsZH9uFIWLe0cJ61aYrMkr
W1YHGUui9FPvoiBYZ0be3vhIRvpNOQhkgkJ32fmDisVuD6siGoiu5w/2PowYc8AFmffLtJsi4sfH
tluFzxzpZUKho2xw0C1kY1tDtqYOYhJS4kcmhlxp5IWHWHrsXsIBszQcyiTKGwK9eMSPpbs76FJX
Z4UAJOlSwxj+/niuHzrBj/pey1jx685ggZew9k+Fy198EY97hGVoVTpnRpugU+392IND2KEwzlH+
uBNmdzDt87oXhJle7EMXFeJ9Zk/gQtZ4wBLBuVGZEmbmTccsn2Xdn6ytFHuMkldyzJP+YJJyTumA
hoyy9SRe2ImUvojXEySXLygR3Peo1+qhCPagwdFMO14oBj4K04MM+GTRbaYxz3bmlwoaJGHRz0kz
EnIh55T+ZjqjOO7eESx/V5M9jZQggK1PXJ32EBRh/uHlG0IcljtGS8OmaU/hbaeX8FKoelh9kJYs
VE6QwMNsFzr//iMr+eJWEcYtyActgLN+VEizBhl0R61QwgBgk34rhibWRD6xFBVWFo4di15hj3XK
UZ1T95Vjdq9HB97gql0OCYIEJ5klrho2w28e5W92xNbIP8DcpbrCJ6EjXXb5mFqRXx/+n/fGXhsW
s2BSwE6VHfOXeR0NuS/FCdI9K8ClMVfRwfU442aqfsnkdB0S/fJTKvoaEH/nBDH5eZTofmdSzMVh
44NvZNwdi4YEanov4rwTkb8KzZUcxyccKhhXcPQ7Aly8lbKjJAxLEZtH35TPfrBnLAMZvLQdh685
8EVjB0T+ucn999RnGx2tcXfDSxNFl5AwgKh5q2cvcBYuIOpIEhIptGvfZxbUtrybnHAfFYETeu7+
pjQ/50oxaX0hIoXkzIlX947zCE1gTwAYy1hUJsFgUPJR9maZ1aQrXZQPT5wZ/VcfWte2SOLgxi8z
GfIzoCSpAhGg1sn8612D+k7Qvv0L0fcrbUrCV1MtL1DHQFUAxmCb/0rYWZC/4n3Sb7i6y1ByYq6K
dCxZX68H+bgJ81SEPV1ULM8AnhFTsuto883lckxZaOawfBVlzKM4inguz1zfo2rNXeZOQ89SRzW6
MR1MuEBEHiqVwJb+gCVi/GexIW8csrSvOYAQOfiZB0wUAzgENYZPr2QOLA82GAppRwlVi2+R9+ct
SQCFR1Rjv1t9Odz9OD3vFLpztkEqQA3Ry/zrz9DPAV6xQtOeszcCGq9RUchCA2xAIDpitBdoIkaL
cNk4Qszjuy3Zmhys8zFExpNRVsOrYsSiHumsSNMo0NjXYBFsFDaKXrufElsMDW8HcJt51arnpUL9
N1L/grKGB5bt4l/gjK3MptfPu8VGmlKXPaJtC0s7JBHpoUrgXtlF2AhU/1nARhWB0zs7Oa4VNhdg
HSo4JB1YXahpiADPwYHQnyL5NkMsTMUux7Pm/4SKjoMnAgF+Cmpm1LOqPsWuL9RDiKAlQNXRn+BI
zzEqtsR45gBlAXttVYuJkbXIPG2iOW+5y6zZmY5QQ5Mz22KQV70wHTU0kE2HyiRVZ9qyAGC/ICBS
B6gRXQvLV2e+lZVtl8NI0dDFno0BL+VfNKwcDpDyjB9ua2jv6oUwncA/emXlpok3O0evDyAYee8/
uMOB25v36e1ybF6UyDi+8qmjDvii+7AKl2SA9JIoHeMUQrYMysZurMFhGGDglnsRYhWVCNzyZx6y
w33h415e52LcGdPGDz+uZN0j8JusKmSV8sTKnqKCN26WS9AmFy/s+BNTDFG0o2m/cSJZ5VSjSZFQ
yd97B7vb2aJZ0HSR+1/K6kaGVg4GQq7pWU5Cjflcvzx92q39Is3BWA3rZquqWyhLUFhczuvRAbE/
8v88yJwSYtcyre97IfO8vOtmsTlRBYrY2Tp4wxewPiLlFbT+TsTSsm7/2PdvRqsO4rUr7PaZN8o+
ww46/yQJ5CzINBUn2NkIwR8GtegJc5luBp5pCMCdYkaMWflydlyS7ujLlByKQuAVhpKsnAJjyYxC
gRj1gW89TTIpuXQsPPHYsuSxmSvsnvHj6itj6LSJ+nOhcfIqvFzn+39Vh4CUj0aOK4hFmK2548Lr
Hntz9h+pkCDNF7Ctic3J8gwdGc3mKABnzzW09t1wBn7EvClxuk7a+tpVGoeN6IYtKNnwIayZ3tmG
DwF9DPhSdLZtYNvHmjJ2Uq1h9V9lqLYV1bgYVu/ZymrHWxCGeKonEShtJJXt6ZUQ0xdLSQUIum5p
ICk1t4LgxHG1d3if5Hu1ncFFYjgJ5COwCq+0dHtfhXkArKxYFpOpFHKb84ynxmLun0md7zumZKZo
nCm2qhVWWf9x1GSTdjoNQ1TYg3nDvHJtkjOVV4uVkmIhmnomBoe3ruAxBlGkFrGmO+ebEaTfigZL
DB9sPe62X6ltpns0wDsJ8OMojn/001p75kZpGJRXpg6YQfvPJKOe0XIPMKEifymJ52PkTp10Pw1y
gvUx99QJhT19AP3nhx/+xZKy6U2bARIlMXPMIItfx+JnvDP0WS2gbjbpKWX0+wrTc4bV71cjDy1a
ifan6/OHE4YMm4WhtfYLZUtLDnkTjyokVsEBryUj402AII2macA27sgO2fkDhh+scn8pqfXwfQ+9
WJAOElPlQqd9BE/A7jeS+dw91gz8830BlirZIE2ybSm3FHhfgz6PwmNovywTYMAIlMv2w49PI7VH
0LP0R7qdV4orr3i6B6DjkpIfhcs5l+4EZyc3yc1dN/6gmtOlwBHKLWa04gF//deVadS9Mg3xTGe9
5vktpcXOaREv9Flw9EEmijzjFG1Sb40rdg0uq6Sb1vKETjZqDe3djToXFdfJt/clSrn8GFA5OSoz
qLsdwccgt31l4v9jX6x5OmeA2qy61bVId/tdOY3oazZB2f4P5hlEEwkBdNQM6KVTlv9CdoMwkJz+
K/+XocVTsc5AIut132PA855uuRQPbbaB9KC+UTHC6CKmy/6LXLCjmQrFHiWK5L0a+XzzjRg7PiWT
HRUJPuLuVOOVwjAYmUkAoUIyGUJfHipZAzGWg+iZqjHyjLcQ6V6FX9FEhotPhx7V7FjM1V4mps4Q
zWBSn/1FA8m4rleZYA0LVFeVHvUxrxshUdlDuHeB3NO35hjy4yPRA3+jmNnoT8tDupj2UTd9fQ8n
TsGADiz+EnmAV9a+JsG4Dyx8L9CWFxR71hsbFPcDEwAF3jA9R+SkugrvsVrLWYo6P/dsiKc+imcx
ZCNudxo6r3IedGLXrt08Y8pVRbJmsZwJGWH+iW+nCTqGAMy0GskZX7wjT8M4Bz5Uvpo3TRHzudfF
iQMEMYxv9uYCSsknH/J64ASGtKz0J/qmoxszIrIf7bWXFIWKKFHEgIIvNNoxWTevdcRKWDeeVVNt
j9YNJ6LYb+0Py+Gu/ZdjVP8jUxO7ffZDjTdU/3UMF5GHFPIBTRhCO1lR+nXDWiIj1gICp4MYCEPR
ISCQMn3qGhm3VELRWPtYpNOWoWw22OpvxvNIWtAHtkiTdyEzHzK3ByPKp2EIdYlGofahhz63EEix
JZkwRuJSeQzXgLALGBuOa78M9ySZBE1Bug4GbRCRumgaH3H12Jcvl7rECopOE/tW6ebH9V6i1DEI
ATrgFP+iuqQhiONlp8bDOuAp4+pouMw05XLFqYMkY/dyQX6MY2XsnS3pU9t/oN3k9oCasEvo1Bt1
6t5qJPrWyWEK7dpyXDdVeGEPSSE1ubiqFmYC4PpufBNdcTKVz6OR5+Pr7+XiVAQbo0beqXD+XK4E
UPMjjHO4NffGv9yoRATGHmiRHCZ3lfhhkulenCkp6XADl1Jdy3HVzaJZIsTYMSN267xR2SziPzy8
gNG3tHQeNTR9r9376GJ8YeO/MYaWkJidDGqza0ZKl9nk7zOs+JL2kfVTzdO+OX+8Nzx0yyIx3iEG
P3K15FqB+vjzY7oVhmxQeb1bNk0xKkyF50Lg8ids9tXk2jYTrd5Hfqbbzvm7FzhZrJdDs5j04g7K
krWfTL5XWU33NLZdf3wCPrIo8TPVT6f9OVVbq1LhNefm2aCk12/XDS8zWtR78DfMR1R66b0qW6or
OTKHf6/37yei+VJcMj1Eg/m753IGua8ynRWSjzAwXPeStfMzWZHTwpbfgrvrbUmuWPxnPYwU2n4b
Cz+7L0X17m1ihowPXysbb2xyZ1DMhU/tvLWS2Yj+O6z4TUvcWOBnfYql/GUGcCmMpQAUEZ3Y/PGl
U6hXYuu6HlX2O8yGvPkvZcxFYroTabYQZhlCBo1BvCeNQme+nmPt/WlNw/5zKLVNlqPU/RktBWke
ktRulKZkmsvtczWWr7IPzG08ayrhpfX4fxrDZFMr64ul5fNQa2XyaqTINDuLf9JMg9VZG0/jrgJD
tXg1/T8kqz1NYnuTPiH9d8lGbyydGkZidk60FNPOGF3aNKjLdECsvN05C4Eeuhm1F6QWGTzapM49
BX3k3eNjjVq6xlWsy4nqFPkZhDMIIGxnyvY+BEeXHpPrDVgVYwUnmjiS6dQSmiw05Lc/92WWa6za
0V4WT4twu88dfi/WB/100xbz2FViGcumyo7Jv2uDpJpGKMA/17MlLo18PyM5Xp0QlD3pHUR5JRx5
wvNHdy94Y/6HLx/SojKCzqJ7H7bGjF8r2Yz2UWmPLuX0VKGNMarvraOxfhzDdk+JJjhjl2TyW9d4
c9BEovRPLxBsGuKxe0wsUT27X7Xh83QoWXB5VJpVW2OSPZwGnz4JcDkcNfupTe9X5Vo/36++/Eq6
/L3a52IGxMiSyIadUjU6RMq+mghww6Ldd7m4broBHsnBEOgGg9E/aXzgK3SIIE9mwn39vSHXVRsE
Aa9ASiJC9NGSMvElgnicvSin2SVIxHfcdpfT0oeLZwxysx2PAmGRUQl+fQxTy2gx5jspl8p6rBWf
y80pKq2XhFD5SW92JkDcsAdOraas9zG02egN/2YxlmeodzmJsCnm4KKTe348ZVmlptmXZ+0QKuMS
7kPC+neoSR5FQrkWTELE/zdmcYRNCB8npd9407J+xJAHJZbvCVXFp04KRq46Ga5PNUrNxNTAHqmB
GFz3bSRGn2T6oWI/7rmp6siLQ5AecBJCVmASGv/7qQuB+xdfF84Uv0I/lpnHxy0rec5b0Je+MqZJ
yqBNMn4TUD8XbuJ+URTVtW+n5qkpp4j3Jfo1TFBpxiS6Y3LVDto5B2CEw45Xc7Yj61XGZVHAjhJc
jZTwCuDmrP3iUpZokSP1it4upSpKELavWQYCJxeDLjTeboeaOMWRHTJ/2EzCQtAP86l2C5BsrGh+
WfsGO69hIxnuweo6M0HzQJJpNzlp4BbSqBSkf5PcPEunLVzipi5HDffYVmu7R8Z+/qnqPeOoXNMp
7n4gwNmRPGGhZX+6Ef6NcXdPec9r2tm1f+P/jjQ1pnbF19bNkHI4OYi0jn28BDWYpn2T6eJ3MMLt
BQtg9zZ/6rSi5KRP0Bo2CT+WZ7l40kOXvh9p/kwmVEa77j+Acj1HTBP7ZwWmDYOUmbqWYkOPAqKj
nhiJ5cOAvVo6JUCQIE/+8U90wfIQGozBrFL1ivg4G1WnA2UifXOzndVJEppWoyLrFU2HBJlT1s+P
hjqmckQsiEACzW0PS+oHJlUauFSrbdJ8NiFxipgBdzCzoaATQ+2pKy1URqchPnrtJ9/H4CQqLwH8
Pu0qsKuX7p67Uzi59PsluKqsp0uBSPII7UvOYAqtZiRrzCkVA8Ot/ec5e3eZ0O5srVMmjYpGnHV6
6BMOGutLXTAY2dT2h3XzkUadlnIsrA/2UUdlRSfX7gUKLqDzU0IRZ1Feyb4eZSw/nT/R4AOitc3I
a5V7i9GIoT52PJTzPxJF7KLXAUGSn5zwlpRK8T14BC9bHFFWQXlc+9fD33vsUdkBdOdv1SL1APJk
YKVwi1q4CWO6/j6RtTss13F6Wcximd8mzzrWRRtjjl5zAeAr+PHC9yZLjNIi0Q+c02SjlZUXKcxN
rH3bUJaLOs+DNGw7HRXORsM4hUhirhdFMEsdotYlJzETAqAw5pCnVRpZJ9mkr5bVXrvy6TxFfYOo
EIz5/J03CpB074dpy1NsQH/NDeviZpOOrxx0SoYFujpBkF2RLhsCZuZyHUqEwQ+fKRt39Iixb+y7
+A6CLbLXrYqto3IrIhBcX3sQDOHkgW6SwRjt112LWPt5Un7j0ouQxhA7Nb/lYIwTK9MKAFncJ0nT
choCCZ2jk9BDLuAIHOgSQ3iNJTJQ8s6eO3XKGzgNgASCrJ1312WbiwSyT3tOh0PEH+3GkJU2+TCk
FxWvZULq+k4U/ajRLIR3pGWO0r8MxM1DK0pgJ95TSydMqsi42ZaepenfikczkIs30cm30m5mgrdP
AkRaqyafE4h5S3FcLbaidcl5630dbmWeQ5XwtRGHw6pQ1v3Y4rhhaYqoI7qz+S/irO4N6lPqkywz
NtIUBUZSyCkZmcEVkKb4XvBBELp1U4SfFCNQJUHu5naT6Hu90hqbPtkXxIgRXsypwWrogmgwjiE0
Iy7ayHv9nv/IOSkUbNUSHM6766bLabs+uJqYmwuQ4k6C2CvmXPw7i7CeDrhj8kdzbOX1mojyq3p0
a+E+b8MHAlh7l+OHkuJEB/hikiT33yt33OAx6LumLf9jmf4Tb6UNidVhB+1566H5PNTwCPXZD9M0
n7mGfsTorF0XHmVuIAr8lLaNmws5GijruYo6VocANNgitSe/9f6edPV+RanT5EYKkQmUI0iQCSn6
NCwX5i8Et/yAJJEMjdFhzYn6CCGnPUPTPjRk1g7hisjF5tn6qistUoPFb2mMOqIYdAmonr/m6NjA
DBw7SsbHhZTK+batWC14Wg7iila1XTo7Ie3Vl7a4t6/mMqfNTeRw9Y1unedcUlCU03BO1giG1aiK
rHsQnIcTNuuABS4ZXfuTaDrgBm9F/dewI6J7FSz1Iv/K48Wpuc6qMDUeduygiv2xdgcbhpgJAEn0
XXST35PBdxHOiYjuAk3Q65QowLjvofvx36gfJcXX5EZcWJgWeXEPAf9BzUhzFOMqS0BkosoWi3Nf
VGITmF2C/IWRTgq+UA6fpl+8DVgmJtQNeRN4qrFflbJT2yRG3CO0Im607WcCWpOnINircplwKcmO
2e/L5Y21nIdyEth7ysK60vlHPY8Ts8wn/D4oAImUhAeLdWL9cg8gZUhm+ndvy8Er8uHkPSU0k+5b
5iKDa+1sJLQPJN+/MY6pjNrJPfqfBIbUrw2RR7da4GBTfzqm4cLeOTZ8tqbjMnvZgUZ7LGvnsk01
wcE/IDAnSgYns+tV7HExpCr0jOehjGyM48anpFyeIVfKeB2+0Q2Ac31bTPNpF738STKypaRgC/4h
Oy+2gxIlxtbndG0vq2cbqCjzehsnNqyv38dT8kfC4rrWh+OTPL53MQRxqhX+JdcjgoHFEqsRInXI
eB0tFHj4+HcseVrP4YRWcj7bKaCDJ349cy3AO8ryg78JsMOgSkO8Lz7BgkCT3moyr5SAd4QxdfFq
X0+HZ0uvMGiRBIjSPecp7n69F+bUSx2DaULy4o6wwqyIThJj2pzreWshsyV1h36+2mL1PXnx65CB
OueX/KxJJz7x2zZhlIeek0lbRjtPNo1YUTAN+Ujul6DCjpAcnyBcac9kprhMpL9rV4tUviXbRAG5
kmUyLUrWy1yY0AN7d4myGjHQFKmX8E2jn4jXD7szFJ2BGc23fNPYVhbnsIrEVKtWGbzw/KVdyLvl
Iskkdl0UZQa1X2UseAjiKGlxDyF+l37y1SWheayd3/M9rSQW7Z/AAigxSBEOUsMBnW0AxI60hKMj
Xkzi17LGhcfVDbhC472/TCdL1hg2nmHPo9dYZGehIV7XwpJKgw/afwpFb6dz8Tq098eN0599BYwK
22Kp8tllgrU1Yyue8kwt1NJ/KGMUs/3E/Wl6pXOzzqY41trhWxf0o0XIcUFvV0YAw/NewsZU4xfb
gwhIYiXiWmfAg0KrAGEsme6V7GubvbgwCwGW9HsUKyefCMy0eEtcQ/FS24RhR1P7s/xK/oQB+6gr
hhW6tKljd2IOmMRFmrsrqhPk9/4ISkXQbR2poOU/gVzCKAQC4sKFzzVJ830j8A8eXcCfHx65JQ7E
e/vYAAdfiA3Cbv58GhR3v+QVvP40nrPfo5QoC5NmaThnX9/ISMkUueBhFbS5OwH0gasQUseH65/P
5cjQ8EmE2nMrZvw8MGHLpAY9G6z4gxgAJBa5iVF4bkYg3rgfENyscJGx7oM19YXfXCx+xK4ZtEqh
yq9jwpXkstgFUTAv10ircugB9rCqBiGRwAvp01oCDM/v0StSn5fxLGEuC5BHl9eM5b1QyWoIaq9G
fT2RZvI4D+H6qUsv5xN4ZmO/F27qlDQ8kolE3YZVJtITtBTFLixWfrkWYrnrihXrSvklvgzw4hDT
L36IGe8FMYh8czCO9XEI9Wu+zGxn/WkLzqOeajL8YJiA5Rp296WUg2hUu/0vrUrvYbWG5u2tN/T9
Dvyb0pMcYuV4ROKgYSSsKnIlgKFBzc+9wIIdPjRjjvO8Euw7B5/Qrp9CJ6SI8XpbPMjJWaMUL2EY
cg6K33RC88IefOcLaaHK6Xq9UkunK8EoijarHXuz/OeqK7Qeed3TRdojRpaq7OCH6VqRjnW4JoFR
m0eskxgcmOkM+tIOAsEDHhm4LDDEShC6ECqwX52KkbSBSyleYiCZq0K209xX10HX8ZFrVqFnnQ+R
UMrMUPnRkQ==
`protect end_protected
