`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14864)
`protect data_block
EYVKDOxjvblJY8/QBf44y3sHkbw3EsD7ii5ab6rUTCHKDXHNfq6PWogqaidiEk80cD9qDrP/uBZZ
2lerK57cVUKdfdThkoTy/N8r3AuVHOUyggk0a9WP5DxqLGW4k/VPr5Zp/jp4MQ6H6taAHv6xv90k
gyTSg85spYmwzyGBtMNpYA26mof6ki9jnxvzB4/dF1UL2oGP1gTS5HMGYhczfcXer6v3lpbxV6D/
xoo3/q1HQPKJMhXkb7lpbugl/M3OGiYiImjooVjTc0TflAmus6G+U8hUzdc5aak76hdym1N5/6Q+
ZnlVvizd7cLLlkr/33P2iNhGBDRwa5m2ZI5dHCFwRGEyZyiF5wtMO66f7Ll2foUk2zj2uTgSnuzd
XdtWsPGb2behzfoVNfnMAeY53+3kkOfhwBA08LghCjgtFpFrbTItoa/e5vJjPrfYEhSMwdrh1FeO
P385kz49vzIgl51nX6CDSkmG9a17YgGdhBLoa1lx8TCALvvo/PUCPYCrrdsYHGErpskVOBi58zwd
XveJqLlEv9Z2B0/k46cENtTz2+TC6bvm+ia0Nu2j9xa857tXdixINHfzzSI9prcO4iaBa2pqqi6P
sCwe13oZuKFboIECab/i35wGyB6dvjBpzY+Oi0oBShuhb+XbKhSStEHznOjM8mThwk+0YZKEFh4V
1I3FK8wRPfxnaEZwirBCS3V8zXJKH4j9lteZ2bSNmxhbO+Bn4TujTLpGLCYwBpku/ej9bxZmuKq+
fyOrFA08j4E6pHrYy2U3w+L4P0gg1j0IwjmSDWmxBS8FVBnzmoK4pwx9jpCcF6EvKG+N3O28cIPl
paEtj5WSGNXGib64jWHrY4Epvt9csaBXKkXUHyMvOrWK3ayt144IZcxqJ2qkRnaW1fl3KJlb4mQ5
PKLQcCUxJXZYmVfrbMLdrkboqF4NUIjQG8ICYLoWBFWbwgL04ESSm9lN8GMr5Qrz4n1+YrytTV83
IskD6aubZGsTJiMFUiNS+l3sO+yzNWaCiHG2TezDeOr8C81gOHGl4/j1JsoVT3IrE6PJ7oQ4eoQE
3XYQqCLzmtIEZmS6ceXDBf/j2u01LQLXjMlijjODKsMYGfly+tl4P0JhZ/6NnVuqnGHwTTnyvQDf
utfD2aYQcn42USiY/yaIo6A0cV8go60FPnhxk7OoGrpPT8gnQdxR68GdC6ZoYHxHkWQxzDmr/GBj
maz4HJz5BZoqS1yFKZKuqpCwzfjsyA0ejUWmWgwz1agaReqACbNVOo/NRTw5S2WV3dYbf2Gd3R2s
s6W5pnlaHIPOWKLoW7cJLPNQdHbjbhsfWtyXrhYCCONy9AOWr2yOcMebSrQiS440Fs5ilyVkL/m2
hbDS58lu0DeNJWt6CxQlJWXzWGOh/wmGNzS61BZsFTPpQQgJBd9CrLE4FrelaOuDpMxqyPpYdEah
Qs84hvZODX4ym085AFQ7dzWHo/AuIlmIA3iRGay37mdvTe58zGeD+lXgz4DsFh8i1lbmFjfTJuqE
f0bjoF3ZSrcrIu5swqJrZhXNtVt0LyYuaieUxzh0SFQxh7SfiQ8g+oD8MtEfTxZEExLwGgNupFsn
1KOk73Wcbb1xKvaektoFkNnt5gwO8ngdnMlB1BYSBAOqu0QQO7UNVRJitj4RVn3zobpK7W7ZVj2B
Plh/gXnRnuRTVBVN4SpTGzvB7hK7mE/39dK0+KDpcMGTYyd7BRBmYaMhuzFtA2L+RdKdI7+5b0ny
j5LgO+waQ/xx6x03272VeD3WxhwE1jC6oIOBDsqS2CsSRr7P1dYPbTbY/Lms3uogb5KXLWez9MwR
l/EovDMmMLIcK7Zels4IbSqhbIEJKM9aYyDCUOodIWkVIg0FWEfBlRTS6X7f769DFwbec0El3DM6
WycFrYZqQPIvDyvD+5nI8+lYk9/T1YlPh5Xfoyc6sL6uwnnwREYCbHigLdREabNn+FJAYoqD26dE
gS8jTdX/b/8vt4KDHCDNW6qyJ2AjKKmmMi9MLKynfGSdRHqF6RW119tf8hoejM/nNgNtcKE0vVgF
tCnSLrrFBmyNvXz9208ZSw/mrcvUQkhoyzXYDbdsSvqbo/3c7vbDxlKFJwc4zfSB0+X6KcwXw483
SvrPebT5ss3KZ+reCXmJX4auEa70W9lRa7INfXPb1RNtgv3y+REwK7Yv2xu8J+XNCHjFVCCV6wtX
cjBy9Cbp6E6EPKs+Distr7/B0pkbCU/s8MsKQoxHUQ0S1hIsj306DyrofPuKMrLfICj0oRzQFCJm
6UydHMoTng/ysokGMsGNCTFudT0JkZ/S32pB37rLrV8l1ivBZzCMqooET1SmjG26pYEQJjwTw+qe
BgT9ICHCxywJp/OmXNNe5TS3myZOHaH1skOXXIefCGxJs9El4zR7tDMYagQC0U17rGGJhSyBRh2n
D0Z/BqkcvaHhlcU21KU34K3wJyyomC6jGk48nwxZvIAMk7jxQesyYA5uDcGvLWMeVbN/kAHiIPZV
+osSFJrtgfwDQ9XZcnt+8i4bIlq+EV9LJ7XvgvmgHRtvoiTj7mb1eRe0jtNDH5IajTb7b5j5exbk
snB187iSsSYtYSXEgg9d7Ksoovaz2B4tX/+xnz9XiIwVdZ1NbHIlPG5xf1oadkv3bRzZv1bX3uPw
A9UslDNsRxYC4WxRlqTA3D16m/PbjiVVnhgE6XOVbxnqV5PmXEVWRBHOSM7gv4TdkYfeY92STyvf
KW2Tpu6e1AC/UALcO+vsKuVhA7ZJmRXYnMXewIFTJMb8hU2Ht0qrWo/bGetsmw6b697OI0NBWWWT
Cfc0uO/rplwOjKfHjLyk9ThTabWdwpA72RB4Md5MJNowFxmyMFtF/pFo+yQHwJPflKdTa7VfTb+y
GpLi241N6kCmYyvJH36U3Qom1HqKf37u5AstzM4yN0TyD8yh20J+5MXsAw3lMZsd5+FXHe5qONxE
oFZKz+HDp92wuhtcGyH3sSNC5nVPt2Qa+dn5Z0QKMcivcBgxD/xZcBCAnSHCii1Wei1UWSOhLKY6
YlZYQWVeNf24Wd5h5feEpMHhdABRbp6UsXLn2CemwOHnMX2WqNsmWHVsk/W3U8ok5nMgvLRexkq8
qVSaaUpVTsTI6XV9a45TRqsuncDRfwKlcV4R5o357dX/WHTuZgIBtUQ7ABIq3Hsn7lcvNrwlRDeu
ydaV2h63Qcn6I9xwHSPWsIpoA/WccTRO7RnfPdrXxCspeRyxF1gNAxoODjPK8j772RkTOU6vDLxI
vWZ/r9ZfCW0Rggb6QTlZhGqeBOLAf4+1cbVvd7gYSu6yCyQ59R8tG6SszUfiGl1ME00ICyIdK3Rg
RR171X+l2DFI4bpwl0zMhnCsfqOF2RycOk9M849kqnM6E/Wpa4APrSbTIwzpdZG6Nj4Dao+UehPJ
2NrGZEBUJDEUgcjGAfDNzLgPONGbCkqS7oMholBETtrKVtyUfoOvktLbsYcPxgpXeuUm74K271VT
S5Teba4OItHWUjQx71gb4BIlT+4TM73c6/q0M/uFfL84y1qoFiJvAY2F49Tk0PEYRc5W7Qum6zJ6
6mf+E/SPWd1023eSj2TO6YX0hDyqoS6z8NqMhFlMJecQLdhnfh/0bmvuu03oVUZ+MtcQtRfBuj6K
8QR6CQymDz2SHMwwEp/ulVrTrkc1hsaY3BaOaPrAfHeFfF1qh7+9lJVq6+4W4AYhMUGv1OHuaFkh
bRbCp875brtvdWIqWT1cGYQrrb5BeWdw+43slSTuUTwRIdNdMWwrl8dk6O5HKc6mYODn9TgxOyAy
1kNy9A7KMWdq2aI3bgZLINYVQ9TX13U0L/NzsJByzMqqceMEPgZGWbnf3sqPs/lsWoX+Q1/S1Snh
lAyHuxdPHLHZpfnZrjRP8dcZ5MkNTNfGBCXqlv6AAeIg0l9gwwdHoyvT2FhcWntrsU47+YrQLRwa
5QJi1xdUupXqw3jFZ7U+UGkYgdKxhrrewQhfVdMN9h5lnHuQWLq29SwuHJB1kHqejGUl8tdKYso1
vexkx5oZSQlruG3XiPyVg81uUft5jM48lDe9omnTSQyVocARbjqEC9vADZDfR98F94Bbd0Ynv46h
LAYK1Ss464ppS798Xl361kaj4vr+GxNm84gKig1fhKCMJcZrhtxdCWYISVP14evP18vcTYWEnhKF
qruD8E8rE3CRLCiZ9XWYweDaK9DF1tCv0Xank+4Z1SBhmLe5Ki9TJmp8wjJqzIsArv+E1wiepkm7
uZcdv+42YoMo6Nn/gAnVN4JBj74MAb78US+M7+nrwfPWgQ5uYPFGOeBiiChM+QHI5cpDoKWgW+CJ
Eoajk/SY1ugV1yBHtN/ev1D2ltJUZ50nWFpe9qR1JMAsZz5FQfTzo6N+EkYKKfU0uWV3zH+9qrW3
S4BV3rHUbmZKl0gdXBOLCF92rLC+HXNfMBQ8kYpYyG3JU8lqdNRXMrnUIGTu+UFhS0zyNtqzuPln
cvW5cdmpNpqi+Nt3u/PLuKte7XEzckk/JJXzhbdlb8ye9SwKd4TDbyLl+fvk0kKAzIhgB9qDYdS0
HthVm3uxw8FV2ZrngtdR86rfd/es4W4B4nasAtzeVoqnepqkXpWsprEFX5mVtlbI9znyFkalHX6C
OdZxfpExZd0yjWjiEeSUrX6Dw2ywLm3jFtaAIQhyCo28lirCircVuzCLL9HNWosnh3aFhiSr3ez5
IBSARfxaS4Cvkz6OzHXxlx7UtIojW5qtXjAJoQChUEulUlPeys6F5OcB0/K0UW+R0J5A/7T03DOk
yaO3iEhwK9egCsmfLIxJ4GiE/i+WvYry1QewxNdNES9pKNL15tDrmi+4Uh08sCWVfVeqBgm64yt+
mhH9IgBHIU2vZ2RxvPivIT0+OIeP5F1+1EdNwZxNx0jTmaRkqh9+HG1402dTLGB8zZzuBYZs+pU6
owTiX8xgYuJfspRg3Ar9DMX0pD3A1HZmmsIRvSODVnNiCABY1xqQzbRl/alJm5E0sZMb89ufatuU
aZBE1hiM9CEn2A403ChehknNnNC6/wXS2PBa1m7TQQKN/bXXIZqLEK/x85QMCWeihosEJZ1CAr3o
TvqzHzsmBV1WCL+G1S5JEZ4XwVV8I0+JVIHImmthwwl17gwQFK+rdG5W5J6QDbs/gecnte2NvXrC
x5H+o0oKdlbXZY9Aw29ZADmragy5s5bZybVaz/cRzZ5ra6huWZaTjHSwQ2NHST+sm864TFAKJK17
wTq/9qlfrXOf9PpRBVv2PVfpQStS0mgjVb2FnRMSIaEL7vCBJuBx6G4xEHbtE7d1Y0QB8/kE0YBw
fuyMONejtSPdbskt56zVyoNAOHqttsSuoQv65zD/16DAMBaehjQ5EzWrTM9q2yYK0v4663ch2gOt
HCOxAE69rIp2wycGB9oHXZCaBMrGvfcfMWavcmehf103aw4IjvGhDG2ubbf+aqFa1zIo/Lzna42B
VfdFnud7xPF50XdGc/7WVH+0cQ634R6x9bWKkyKtsDPu148F4/lZjVvekX/WHIqQl4rY3fAzybzc
l54wAtGnJBac+5bXw8LZoO5GTtvowsW3TGqKyfRcIE2M+Q5FUbm3DAgxXWoTZuyRWT4LzZkFuJhL
Ymd+PXcu+EoDn3t8EIJB4H3yGX9onzXrrnm9KTBEplTnFGcbxHycPinzzc+YLQvHMUy5tfSUJo/t
9yCWUA4qvvxnlipYJIBg2e7COLYLgOfbZnNfUg+9mkiEm+UfdXaXkaNk1HZTT1ShQl0BLZhCJHfk
QQtOR+Gypr3TkH9v/U3FRrV7nLZJnwZeYORnTvN9Y9TaaQMf6YGIgxldyF9S5kOsFApsSyqNoJN8
lb3pB8WieMnofzWyqAfTNBQdb6m7neNG/udjmLz8SnaFxDAoeNTEQNmXakTOyI5UD1ThFnEzBVUq
XXgLlUcEPFPywGDTsZCFO4ohJWBQRvxUVu9LsvX4Pa0db3ehWYoq9ulcqEP6QmPgEBkxnbGheL28
jYA+vKcMft2tGBXdN49Tk6X98PiFcsNWbJJxsdz9Itz46X4bvMM3518DcVnt12x82k4SC0LMDxLq
yCJb44rFq9abt85R3bZCjsGONttKUrX1J2Z11ROlpbu2zv4h360LsPsHNHMeg92pK1wTFlW/cHHl
BGs24uGv0Z7bLLfiafo2ilytczBNSTzD8wjr8snpqyPYnWTMKyrFafowkRAxutgyZ3XcJM+//7vo
k7rzO5/ADO8cSfJyC7p42gP0Ow4vrxoKzW8kmJvUbN1akjxKwI+AZQB9jPCSJsOU3SLICX2s4uaE
Y7BV+t5aVHEkbIzKyACBSxgGAq1f67rP/xd6sWGiOifa9Y9XXqueuTc5eak7iFKi/dqvFQLmilQ1
0lsVpLclwUQKBm1xExi1wzA8VQ4J9DEGk/UcjJvzkskUSVMCclAoqDB51tuhl+/QnzpXAV8qr1To
8rlSsh06AlWuX8qdmbsEWvXz3+H+7130ZV5YgTogp5zHtklCocaHh078RTFOu9/tWhZtlT7eNQfx
UaoNZLEyamCE1yp2fHNpuTSuAB+u8hUqw67RxvavNLIJ7IBgg3LX5xNgoLZViZljbMwyHThexD3F
yzpbYBekIt1DpyabxVie/lC6bj5hNgeWHCIJYuEYTUaKWoTBEZRLkD+zg+6Q0+87kzxTL6mOQuKn
MS6p1bRLjYWtTg4x0XL3sXBQz/5RBMnNVUq6IPiCvyE2/oxmon07gMN1hShM0+GXBykrodaAMWze
uJiH6cm3cxnT5P5EyoPb8fzTe8JY3BZS07UXWQSUijLKpCPpSuVNK+hHs1ALwlxeQcMzLYyG4SBL
xxFxKUYSffJXPHqcEkqYt0A8MdwLoE6gRmCIODHxP8Ouw1M0kKj/JQiv0vx0yZOzJQiyyT1LKKXI
kHQ9UbMvEDwZiyQbdXU0eEamSlOIOupnACPgY+E+KJ09cmcMe6Rh2L4f3zZKLpynxMIpNbHycaoa
WYu8HJNiGQpVBVS9af0IhLKrzNqRbAorgdb0orHuHNlE3dKXmhOaB4EyncPAIKzuFzWPeYEdx0K4
/SlhI892k1asqNDVd3y/5inDBrYnjSIevncCyyRMAQwDwgvtpcr1k3/owW786BmpLmtmaJ4yim/N
0aLcopgOz+Ajmj6dV8LcHnBemE/NBtXU8N0vxW99nsuaJbMN14WlQmY/yQVXhiyE6tmDeKVp/De2
R5eI86tjGFHayFMt1DR2HaR/1bP4Xf7g1Tyz2d1NKJDl63BE+j4FzFjbA/cA5GCqEPQUgCbHU5FJ
XoXJCuQYiBvU8kdVGMI2qoBJz89jpwnYavhNbxQbqsAvV3ZmVdYT+YWM1oqVjuAvdOlvdTxbZSPv
HKif60FViPuLDB04wusQA3wCU46I6G/de6tZJnJZCLmToOrByOlFEQYwW9+Xk1XNsdJ8h5iY1nvQ
eJaQpqqTNK1vKcuUxsByK5YluSGzcKy82rDx8iJpyAuMJIseE/qPp/EfY6n6s0eylvlw+cVrkv/i
yLzeOVl/mq50+Pkq3fRpvmqtX0CKbUWTelLo52pEZti5X/EKJC+jXtXhp/MpuZf/gs7QX764dYbe
4KrSq/4Nl+aBt7jiHzO+yDsIMvyTj/HaNoT5DrYWQ5PKoPST0XCDB1bfSN6nWcw8MOXQwFuYBaN1
gn6z0KdqbMGIKEJzZucCA7IiZtJHjF7cyiS4dmyDq5nFlHTC0+rrJ1ecrmC/c7B0+v3qnOcATSvm
GkpZXpb7sJFamS3WqGU11rpozbSxRjNRUEWoXkPUSWRn8GWlilEo5cfVaWhTHfShaZaeNhLZTloS
I9FL1DpxZGoc+ZKGXxYjt3IjiysraT9wjdW69wtW7SLLEx20Y5KgkMtin+1Le7qG/qhbEtdx0p5N
htOAhegywVSTJQ1t0i0MzleNrFFitX4GZp5K8VY3P3CnmOAt3I8s63NaElK3uB2gqvmDim/PZmSW
Nltr5hz6C0RWQMCkYkJjYbuqWGSiNzsB2Tybosb8LcZoVACAVQ8dJqHHvm1j1hn923+pl9VtetG6
QZ3Vq9EgXFGWDi99C2xwQav2ZrU1FhaqSElIrqoEVKdpYToa4w5i7k0hW+vwXIsvE+kF/0eF27fF
l+rqcF7h9+00nbfxeoU/2wPYiA0scN1stb8SHicT94vCt+j1D+HlQ9nGyz1tESpUCyedjbbkj+UV
zwKvbEbvEKaKTDRJVvSKzqU27QmGgKJe0whAl0najl3e1OnTLizz+hVyJ1kTRjiQUaGT5GkrmfWI
ZkeqNY1xENGPqPakBft5cQAHyZBOL/z/du5qcGCkqjYUv2uQgriRAMu4LR7+QoQv87RHjvgur91b
/4j6H9Q7Mrh9YxKo+hm9VxAeyJzGnwt2EYvtG/OwmWqefMzgzWCj5xD0wkd0WQ+si+hO/nu4VBwT
9fyglkP4ehRZC0LFhKjEx8mZobHa3nFpTIpf3KQEkZSSTZFcmP8A74uTRgbRlv477re4UaPxNyRQ
t9Udch4c1t0UgTWyG6NSYD07o34kFOhrIueTwCu5toU6FaRnFtAzAz6kzGB0JHGKHgR2C3qz5SXh
q4DH+yHcVJ+RbkHpdJqAKnyUXNdYtI7I0I7VW23MCIHH+Azn+fAl+EFjUzlZS0QZnLtwEaNXiGa6
MoDZPG4cR9j9G5nt5oAu/eXYebmzNfITypCKpL5y/wu2PPxC+QZ4K6UX0/e3fy/S9F7MhaqMVKKw
Rvqo3pvMSBrc/PDHszEahfEk08ouOtBufx8QzXkjam0N4epmuS5+hmsL0tzRKWrofE62LP1keDEF
3gbu+xokoVj6W7kPxM0K0GRkiPqSXaJU656k2g8TIlcWa/Rg5vSM/WN+dHuz/IRQHbaaaWKpszBh
pYPNWHp+LLj2lzOz6S/qdB9XEJR3HQk0hK6bAbv/2cwjNxA/6NrLL/fIkPPryNXw4TJQSmTDV2nc
FfkRWERXfFf23Hl3+9VIMho0voJxKAwvnfdkHjSzHj3nTT0+0avKtFCskZ4Oyo0ZspBXU8c28E3r
o82azF6iarYfXL1a65GXhRShEndI7aDQJZKbzuNmSXNRGJJDYvCorCtOzhTHF2P1IPP7amcqCpox
OvnPHLfldg3/0ZUhyinV1m4d+Xr66ivORfuvoS7mOBPf5JSoMUCRD6h2pMJtHl5zSPtctxmhHfVX
qr/d58svwQ41pJi/TurFgMTN0cCmFK4hj1PLdKJxw4ARhDZJ/Yz9+roCtJzUMOGBRPVFC+rBwj+f
Q13oM6BU0mEXruqTrNs9DJorx7Loislf45T6sTgHzVC/ym6x/nWlkoW8xnOC+F/SJ3oCef6WFyXZ
sn2uZrHu8j2/6PaDbcAVO/z7iFHYH7CHpkU+qxXJtLa81kgxxNVEejr3M41kbX5DxZUbKVy6Hd+b
L2hhvnLEbPRRH5VJZYETLAixYAIO3YoYaYEI7nZWMfJb3D36RSN8m9q3dvOfhrloemqD59sJGYDi
RkQoKG9I9p/V0OLNd3lg4NcNYt3nCaqEJ5awxjF1FDB7a5hTuzIwgoa/Bq7xFXHfrVzgLNYspUu3
mL+DHn0v9wMEH9KafWZHgMiR/5BI1lRfEpwjdLzEgw9Vjb5y94bjZ+2EiLIHbD8qtWTlA59ivjqm
xwlhVISeI56jAS10byPEY5+bvNqpEfbapV2oI5NTrimtrg6obj29CuSN9p3CD53Zmg6GZxA+8/ns
vyxYfP50swIZUkFwJQoDAUdzzLTUPNh4XQzRl3P0BPDV5Pz2nAHeOX1EchD7BFtT/IEvKhjsXtUj
8dOAo417LVeWCdQ2kprUPigmhqflL86LFCZa51S34Sqy7N2QpkQRy/BIo2IeJRM4Vc3QJwO5pSrA
Hse4DapKqs5YvQX6t1akgn7mgA9Q17I3Pxb7BcPZWMjCysrxWF+7LGuXpnpLNi1xJU9cu6jxrOte
iuQWcO3UXvY5A4KYusZPNz66Xqc289SfB526la+N0o86jgJDEUPWfKuas0PkdqEvWfdJsRUmFcGW
oD2G7QGp0bCae6x1kSoGALp4xRzNy9hp2FO9eGnQURCCrciEs/pgyePJHo9VihboX7MZj5Iymq3S
JmZ+sTWRTEOscv7WJQqDzhqylrKUUt6w0AwIW2tPQLsu2no+AH2wEvENbKqxrk7rXUWQM6U18yxM
owAZtvYRwFx19Gd8QZ+enstdbwTwNS2jExQeHtm06jNIFUtspPcTG6HUk207YrE7VUeoo4bAdIRi
r0sH1XaBqNHa/b+cNPMabGoc3qCXZ4g7zpjN6SPKZAgM8nUrUvopslWo3tUkduAJajYSGv9rdo5X
281fRRrTMsddqmeY66azLdeIItLu1z+Y4UCk16F0Ahs0YiCBgsLMy0E519UY5WodIP2ByNSyPwM8
NZlEZPUxvW56BnDQFxXvXN+YDMZ7KhJHUD4L5yeWOslFZfNkzIQVGTKoE/FbRisRsrynsL9c1hva
oguY5f8RGyWCOtPGIXDCMacDMr84YrZ0kLd+AKwllX153D/7RyJSyt1cyV3xsLyyWqkDfo3IL4fS
6atNT53sKB+Z1iQe2afmVEFu661J3DqCiC2a1UhZtzkCccA5FOlnx55zhapAMlqn6K9NUVvdBKyN
IzBdR/ETXbgEdIGnbRDivIFPmlmIVWHtJWYUpTd3tZvh+ln1HJmKFX4bgMK+GhpfdO0PaCde666B
j8c9SBdmaXkqswoN41twzqcn35Kld2y4CLyQr7CLuuTudOZ8gelojm/M6o9hNIczgQHUVh+YQlLZ
XycCRXygCpQa+qzErbpg/wqO8NDNR6A+WhEQYjgykvUxEWvZBiku3W18hFjZI55tMF1qJB/Zq4KY
knhuAUSdpfxg7A5bPxY1haw98Enruxe36+w//lox+lgvpP4lt0W/WfEZJWNEyirey4qe3KBrCeLE
+KTn40NFcPWi4Fav0wPiJcpeHa5o98CXnbqEYJmKTARqdbBXE/8mS1XELpJaIWB3QL24cFVEeE46
PRvOLb73Feres0PpgHzVPUBMEyAM2xhRWpz9KPG79/qEUxQg6Jyr4viW5rqLXslm3bCdq2cTFN0T
IPt7ADL7g5fM0jSovgjBurU8a2ZAu0KHjo46SwwbyVU43aW16+y+hGKQ38sT5T3sNEiZruQI3zdA
2VZc0B/cWUUgsbgw7UoSi0UVLnPvEBVIUkOpRsk9Gnnim08fiM4gN0jliBjeXxnvgVzVbvpXyUv/
UYTqfa6l+wOZksLE5q7Pyj6cKbreS873FadnKR9CRuuqJkNaP6LsbnLJROI/DZNoxQQJGr3srR4r
oeDyt9wQ74DIPkp7Md0fK6skP0fOJtTMhT/3YoSiQIfMeerUERV48PI7ETvK2yHm4or/xq9VDBmO
bAsDQITaGEYobNSAPB2+DhSznMdMa5NAtXxxmGzBTxuJZD4Xr818CkgPo3YigMo18jxF40XkXz74
5zo0av4WFhWslAHkVD3/324/37x/2yVKoYPnY1PsiADU50CZLzbhO4Jh3TAk2gNkuVTZvgvN92nJ
jV73kjb3pb7ccUbOwHBGf0f0WlGqgEnQD2t3qTH8lcEmsdwdWz9KHQCQsFXsU7r8iOVm/5hpPavx
fpaCAYXP3XXQkTILC53a/bSUqOVRqaItk8SN241XJEQLa7gKzcgFLD+lAqoPi9tK5NWImJsZnF+i
bos3QHUzjIGPTKeSqxQ7ih9KS1jDa+xKDAO2FknS3eXdOCZ4pbpiW2r3zGRhsF1ohLE8eAhnzd1J
KDSA0VaaDeWuACOA69BzJIPSqLkAbVPzJYQC9Nf8WJvq5pCPhb8NvfbXbbY6zPz9o70Wt8XsQyIo
/4OsQdBWv1eFjQwuUqA5A0zh09bpUgt22eT8AYJDFFrp/HfjUC5QeJ0k4+GhsaoQsE6dfRIXR373
C93m/cqOGMCKwqTeaRWBC8gTAHodJ5HA6bzQ4H8eWWx7IpzMMFlfHqyovi2S0AX6/dpC511rI9OY
Z/qyf3PGgFx74xqpqa0nUY2ZtaygH5WWx8MnXA8z9YE+q1Y8RQ6rwyxWXLtQZPwgPLKmfezVME3N
OhUVPrrMwfLn0++2rvvMv3rTOesPRziRG6l29jrF7deqsNfUfSSfi7yNTf4nlgIy64zrpERzSKaY
BLwMLGOoAN/j+j1f8ZuG/fIi6I+ExOqXVJgxDZOy1wJens3iZunhKXwXgMX/pb1Gdn2YpwHpd1Jn
/VBsKqEWJ7sCe78tX0pxD9+48DOHmz2fmdiDU0ADOnwqbO1dcV639fWYgPzkyyFb6LRu27vl3wkM
Hbh1u6AbwUFymERJwta6vFXr0o3BEB21ObmvK/P4k2vImNV80AmQv/x6qQRXhge5/4+7HmfMChIk
dngc8cl6iqTabI3YD8XzmR2UJYV31UTk4M2787x3dMNHgX4oX0rQJCf9H7ryDsD0ziTajWrVlWdG
e0es0Edg+IFAvfp/EKItEjIcnKnqTtOG8lCcM1axkuyqPXmMA43GgOFsBjS5oYkflo8JAkFrwRa3
V8LTW60Ta8erTp4i9jkvdsI3xcZryz6s2HOoITntBqT45Tv9gCzUJzX5gtdrTxyiakCnYaHavm5w
Rve8N+yJmin38wql34p2aRtZ9Xl93CI6C4//nqWCTVqu993UqQeOj6Kcgp+/Qw2iamdSiuLVMBME
GjCmjJL/UEOvUCHTnPo6qFHgqPH+klZN4SaPkr8dzqUasjQa03hHTOemvZwR7s2dYICRSWPbtNzg
Cd8Do7nJwzQ9TbGB2gdLtaPwIb08x5LkPhCrLX3Lfaw5LGQjX6cFiWIzQ04Q6C6FeG3bAVvfXAdA
/sY/c5+VK39pICF1LWoASQL3nPHFw8pcIlC0X3LwX904aECqlrD5Msl81a9iSDDuX39RDTHghggS
Enw9OCBNqdiiHLqcgfU4cxlaCOJQN9zMpDwF0MK/HyeA/6aTCakVMVJ6rbEIE5V03NFRE8YcshNX
MAfy7i14sMfnDxyz1MBm+0kPDW7Xag9djZsNNzE3FvoT1OtvVqQTchNhbvGWC3wwllwAf3f/tqqX
q3PKALYUi9ZTxFya3C/fgdFzEUUDXzHhVOm+CYmKLfc2G4Qg8ho0lDU52I+Lq3fYbc6PcIVX5mK7
DtKKomQg0j+sHtsZsbErL0KNGOpVULJl362yKGOW5aAOYjS3yaH6Sm4pK0/SaG2w8GYn23FiW96R
pJ2kcU2kY1t7Fh0LxASyye49evhvPTKO7X7eZEPqKxk5W94beEQoV63x9W8wOl5h/dExG9RmxHGY
dnwWsCcVnvEGM0Lz7Au/Vm+KTmsPLmzHcAOBbuuzlpbWwHeRSBuWqBs8WiW2rXQC3VFtaDe3+ZY6
QOO7LfMcKmn4gFzIiObXih+9Y611nyX8thPsZPYADCLElVEjPEacF1YnWBCRKytK4juhRX9kd2Oq
/04j1BX5OLGtQ+WjQ5fyeNWtKtHnZdOsC1qSy2UFRu2a6eArxTixtiadAg4nEMgk9WckOC5oBNrq
+ZFqRBIz/Z2EQgdo9P58JhrUHTf86l8EzczlFVZqCl1wJ8qLATTlbCYAAXTecGbFdwZ3Ty7aiD+4
QO06damwiGLaJOnWkTTuyGtYVIjUVvCkAoSOvS1h77/9uq71JcQ7W+5uq0Qek0ydgdwfopNe7VgM
58c13co0E69baLycPVW1QDAIMz5AawMfiCYwzn8xQQY/5UH9pdav8dR9KQmGaKwxCTX34j/gW2M9
s5hRgI2ag30Gc56uTmcmq3+/F3Vqrup7INYSDBXB9VotLqfcymdcAhCTM7dH4LR/FlhdPxAI5za5
sdWcfDM0tWk+7DLodlkKLmNZA8Ka4Z7ssaFtYNWpfCxJFaBbGdWn8y/MIrfP/SjfRMZQbdBVboez
WvTlhT8r4I5vDWGnM99tVoGy4Teg/fXnZ0q2RvNrNM7V5/bA+GOYhuL8//eJ/IRzO8IwGB1e8CY5
W0l8dFPzraxkJfDCs4TJfZHbKRAXV1d9LcvzjmiQwBGPwRZ18W/CoBSgpmk6cHCKGiJzCIZu9uAE
nHfTCT8vIhQyMeQEEWUHCNoAS65MQQCMXMsUFOtkYc69mOFIiAdZWXIrA9vr2HYnd3LXQpu4gU4H
YgAPB2xE+A0J4cy/G5OB2gH4CP/PtfdeS50s/yuCz8qqLr1HDnodkuPT1Z+ZF6EHdTg4MuvH3Agn
DYSkRdJVBi03qCz4PFPoA2yrg4Cf1mxEec6eSl2l2nHLFLK2CQ41i4K7O+1VprRdAh+pHKIMkgc0
2tTHwIH1YJTLCb+r+6g+rSn54U0UHqnicfuTH90I/y/L29J7OVQLN+BV2j9tZh/dRP+lcCxzUA5j
Hl1fowEPaWUiXsc9adEmfj8gQBP4F1kgcZozptqhJ4EWweSalKeYqN9sRIM5PgJ+fhI53inPryfA
stGUQ0PNyh2TPsNS/jor2yRJkd+JsJZlzsTIGfa/I25xXl/4MRjwWJ6f3wAjzFoQ3eBPbYBKn2DI
c29jh6jC7dVuejwWq8EdKUgz+DsQLWbHEDO3B9ERCUmCIy1/UZr3R+w1Dx5PsCZ6HkyWoPM95Bvt
xztmX8I2rCeyuWrhxhXHuGZGkvyGjP5E8FasBfJnl7rKwtHGon967KMcVJqoqObUNn0FXgo8wYdB
6gx6K90Syon9D65NKfzirA5UZim5VekMvz+lSKvfMeVeLY7OZ6vW+egsUxcJpBBlCyPdgcIp0PYP
rIuTOcVmmyqBj2wATZ4nZjc/5+pipKpSERfL+WxyPXVr2+3gGfb4ob4GcMy/mwECT9VF/H9gn7f5
fXS0hri9SijxXniTJYFKw+unWRb4rYzruNg5i5R00l094HNlYJHqgESZ+h5vFEOXxw3FhJIZ7MjX
yeySheAom8nD1MVAL5XaiRwTU8mQzVFWjOqF67c+0Ym/6VFy8FBAl9NC4YEsZ/3gC+9FqS9cDrv6
nrMbt8xtIOuUotd3z4wt2y8L75nskrVphoJ8Fq5w/nZWGbIB4xKA2Gk73RTDs7A9RREh3trRsJ82
gg4PMy+joP7ITzMVPlq5pzEd13IPhzyR1lt13UcVUt0qtumZzztiNPJ+baV/4b1tBPe/3kDho+/T
HM4s6n4NEPNP2QKWmVh3Eieys6Pj6gloKDffDg9exXnH+wRPTif3EUW1eEkM+fxCtnEY6cA+lPM/
Ig/aZ6VmkIoPGE4EzwgNqMcNd6I3hdABfU/RWDocq4v3eIZThaKvVOZFHJtCiVoka+VfAnfiZJCU
QNOLJuQRghvNGbFM4MiceWtGXi5v6dlzCPVSCuXD+gjH2pTVSdMTtwUYY1kSU7jpBtMoG+9dF3HK
vHYKBp3iGRl7GBBKHxAPWMnp7ihwmWFrwaBUJxewISxWxrgDOPfszIFsa48wEWTfH1OcI6Nqp7X+
sJa+07+oipvvZH6ZWtRf45+jfzWvIpPaPTD8cIlLaTWIxJN+0wYYhnpJ0kQRHwhYBksALTsRTWFJ
YWF1wNSJza++rXguUDJ6/L5cJly7w/PRcEEWfHvG+pMa2r+6884Fdtgt3XRVJmVPXv9dvVCAyCNS
eC3JWPbX9FaNU/9PGP7NiYSQcj6KhxuHukfEBuEZSWybDRjDubtD5yDHaW/4qCfyHSOdWKPDzspy
lDMqFItVeQuT+pt5ksr8dI6pUbfPSlA1V+IuUqC816KnHyn11S2mUzdSpx5jqTlihWQMm2VP6l1X
taJ50hv038N3xRkl1fq+ewM/zEKR1okwK+cvlKuZZJqh5PQ0QG+qR6UE21vm6kexozy3E9m2kLcJ
LJe4qMDhzsi1xck49ObYSOD3l3PPbMb8UiHnLBj+ZMTpM/yaNxif1fTI9oh7BknDkuhurR59eY3r
RM0Bt64YYT8IanOsQmyOnfD0c/qAtkhKYywgigbh3ONJ1NqR12tlNQ1LOArSOdS1dnYN8Wq6iVxo
zmsh+y8je10qqlmC2E+BfPLq90/Fkx06hENsIJq56PdSFU3vHRhjK22+RsQWHHjNlVt6wwkW+Rrj
Y2NT400CZnE8FCmDWEuA2Vm2OWV4AV1gvXMDv4mgfMMGCzGYCAz+vCSpkblUiTub/scyJlFqDL7b
vjHLyL0fC3oj6+aXc4mhFhnnOEV3mUsQZ/1rfxFOb3XL0azBYqDTn7u88SxbeNYb7e8KrmhI63Yo
55UMVfWJNVrAMO7ZOQDNyZ0T/gvNGU6Cj5nVONxrveAp0TFi6A6uhshReJ+ciuuVNaZG8XoILvLk
WHyAdCqYMvjOQM0ex5NMZUAKGwpzekvopYLlq4Gu4rBhMmPl+GCxFALJ3ZVfnl1MWNwpt0BOHMkY
ThzewP+YKl1FwbSrhd0WVpRI2mfPdVNZKvJb4n8kpC0pAQkHALBLvTXLoVmmxqVU4uaPNim5Lw62
Q2YQ/ng1c8B3q3NgR/ewVL0JmAbAgNHTd430pmTBIurz3tR1QXcj8xSrwLJeSR75Y9OX6sl1r7fh
pPhYA4r0lbKp+ys3DlpBSc+CMcW3lueM5xcchd/zF+SN7N9gBGEA3aHgnxMdfGb3enWZX9dGfrkd
HPxzuiaWwTQMIwxAfa5AfoXiw+A41ULLE3JXy8h8GQEoDZwlhK3N5Rrgtw5fR2mriN+3i/316Q+O
cZyEhAYT24Hc6MAPdR8Zrw5IRuJV4iGljbfq1FLLeds/eSCrU0oegQrYxgmX+UnjI2RbMrufEShp
QcmCnrhMENWyaxGF7wDQGOhw13Ug441l04DR4n2kJILxUW13LGQiG7B9o6lRRpJKzNyQR1/diRLJ
nxKz4zTj9ah2YlFgsj6tsd5Ky4PqsEIUJkg6X41KCkVkwDV2yrRaKxQFCbPgtiTNJN3mMtEOiAxd
WBmTPYOAhBkCuk784k1YG5L7SAEXbWcn1xrjjDhkITB4Gv+URJLN/+CpwAc0ZSjg7GbUbHXmZIqC
LSdo5mJqEVTBwdUQGcvKfJirNbDXUOKAj77ciAVC8YQxeeP9BwTNlCJW4sqESuiFHh3aYcTG9t2i
mzB4i0JXbJbYzlMHvF96VBE3WrjSI6o8+rcIKgLLF+Bg+DCXeZonytl9ur0nIGkxfyYdoaGq5YC9
++l3LBXtwa2WJKbYA4bB8pU4zZNioCPdEzu2fM/PZ3eYRlHWCjjUELP9/lq+HS7nYPqLa2oPn1M/
mZeXz896GfsZSRwvnspDg3JKL1w5/jN7lGR/dfWA67kZhnu+0MRonizXgUEcw7+/iDwztT/TJNgS
sOxnZHXYBmPzfBe0huTLSMPc2fW7F4Y01C7OP//uHWenk97uOuPFal4p1O9CVKnowraxxSZ1PVJE
Llq/WoOYGm/Egji24KzcCtmI4yZgbirt1H0KLlgnOPhRtXISPc9zlIR0B9eBctKxR0pXPIC/YPRs
rWycssURZZl7rB5yoS5TgNJABRYB9MeaLu1/OUxrMmh4pKxXIVUKEKtokla9jyFFAZlFvDnk4rKj
P+k6eSlZlsnUZ+XSUXU2hxyY4wyvgf5r5ROIS4m47JLMcJ+N0uMuKKxpLXv2zB13a5Ifsk++i06S
N4LWRj8lIfbmsBXQKDRKXbBma8W6de4jjl0dQNVe0rvvCbOOfUmHaqV8DeU0jZmKGnTBEyokQ1wy
tSkrsOp5csPv4bhUrEJApZ8i2eb8rQhKZ/mEYBB1xzt8zWFQ+PNzBVEGn9rudlik9ItwxQpuEcye
8u6Jk8QUstQY3RXCcT/vmzzhsbnCecMIVcTGtkyB/WSHNN4QLjHrCB7+WMMpLIye7pQKpO5xM1Hg
Vjl+hAqAs/ma3MshdsKW7sKMkdG6q3BkV/qjGJ+WqSi+asHn6hKukmIkkP3njDK0YErThuywUftd
TBxGLKcwnio+e7fpyymt7fzDYIMhGkMJozVzH67dhUHKrON1EwO/P3b9dqZgtOvTn78AW9qCzCkp
FIv5lYO19eKrM8Y05ojrXLJvS7bs3AD+ErSQEj2ImvHB2+GihesVxeUXm8jA/khcaeASIeF5fR4R
re7FQr2efXX6ya8y6exlMq5EQsouYSAknpXdcDwoMbIRY4P6pNNA3gNWLLS2m338MJA8S/YVG4wN
rANHJhzTLlkA6NAH2AMtu739HFZSMg97ARQVl/0e2ze6QgyhzlSpbPKyBebzAk+WUtAZ9IBMN2Eo
uEpuhV8zFYnw96wMbloUN2UX8JA2Ai47EGjlw9X5sT21FhUao6Ux+6OdJ/7+rT6dAZn957235k7P
f36xLHqmZ0FqLWW+F8bceaBc6Fkt4QUN3utfnWhU/+Yk60Xmg5iaacLtTHnVJyYWkl2pAnQby+hM
rab0X6klr8dIl3nMFWyppt0gRsqTXCB1+PEDlCaxRkAw6NiuL4JvBpFRfcqMh81CXpbFYg20s7Cu
ivtJAlRNr7HUzW7rPkBcWEVPCt7ugzwydkxnb76S+FTNrir5XGUkk6vuuKDDDShBvdskysRMOdmj
Vm753h08TgjfyC9t6ZY/XYgNWS6akD3n2ykexPBx6u5mo2fdM6B2jDrxljlAu9PEiey+5V5SkVMU
HUpqi2y+jmgueqmf7jWBTreSjaT2cFmxUINYD6NEupyl6tQi2ejjf7b6pcWrgcFLJLXqhP7prOBo
qhE9r4/JKV62PPvuCINr70X5EohsHk1Y7YHuZl+ndDT+zmxe/uKhFwwFmo8drSaQiIVgYykrcZBe
8PmNf/VngIbCo+/nww9C7ZQel8djlsUBsQLLM2DfZJLK0TS9sySr0Blq8a7kADy6ysvLhpMvgIZQ
lN38kc9JYbj72yTVKjKDEPbETPm89xtP5LVL9+aXhLC+g519W+4JuLlJd+l1vB/p3P4MQvJuNiEJ
vmhKJrHICb47SbBtoLseAsx8ooqLNshCnYGNjgsR7pTgINdslM1ouoopV/zhhw84PRhh+iTF6kRV
E4w1BuXS6o/o62E3s4ONI3jqeeD/IfiM/2KzlMtClaxvZGJQLdvjBcJ9UAPDxoAllVupB361mMcE
FZ//HA/ADdmyDWZJguQDZ4ooFqoMT3cfNDqwgWp8t/AggAwX6zWVTKHBAOwoAusX3jV+r67J/j+t
tjTMMTld+1veROcyYCiV9Wph1uceXNxq2ICey7oKUkBGrsB3IHT4UmB5YwwBnfVquzgzQs3CXtSm
6YpQx2WtdxLsNLVcn6xhUK3KdVH9wIhsXk+blOizQ8b9R5+DGSUxhGbT0yc/ch3Fu3c/gFp2IqYs
41Z+K7PJTDeOC2nXvh8iIc9o/emdr2Iq3rKslkJgveVmaUOkpiIQAw+aa291lfi/saZrQAbrm6Co
UjrExcVjqoTfzPcAlwchPcL0cydc1t2XV8kCaLUfCT96OQQE6TTz3LGEaHH8ytVp3hIyNMdGHZ17
kQfrgz13m6oV06vNY/nXNTwYWo2LtduyRiXsAAA6alCnShdnOUYnaLe8W9xeKy1BpwS4SykU5jcf
5TTMpIE3FYndyJtY9nCwiJqpgGFqyWsumN4RRgzMLs/1B9cf8C0IB9wYvBx53zyJbWkXGqWfNylR
uyOfj/rY32SIBAn4QBhb/0aqTZ2dt7N6o3Fu5gdE+X8p900sIyK9iWfcb2JMpYR5bUpmHwbvP7cR
osTu41BClcob84lY9G4+QfL8ibLpQMxcDODnMOASAD97J9PF322ijNxu5t74/o0zQvMaFHAjHZXX
XhNfZXyYIFljh54RL0hrzhIMLczQfIN3xSEvPDnytDDMFD+cUEJsMYw787ya31VdJYgqVFpap6aa
2u2rxeukaMkJtSuOSmTgomCUAqQtK1HAWQT/csJYd30+IaEwR2xvxr910Gg=
`protect end_protected
