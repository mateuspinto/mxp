`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11136)
`protect data_block
com6RlWXnZXrWKT48UfVs9sW7l138Em3VqPCd3QZ2N21qdPsmlOZzXfaJ0OSyCVDzJRLkwtiH4/9
vCbeQ9j1nc960jRav4KhLaMx6pR73ujGsT53oq86uFv5slorQSK1v5fPQS7XihtLLmtelO3/yygJ
xoDeC687bCkF5tnKpyhk37tP/Zy+8mgrmuDTVSucVn17j9NXn6oQC7NH/EdIO6fcAqb3WNkce1ch
fpj23nzFf9aPmgaiID9RDm2pLWNKm+d55587rrC3h4X/qoULW3p6LQd35rtzNOoeuymng0BuzusC
QKtfTTy7jfkdnGKfx6t0RXA5p+DXXd5i5QejiIwfyytcgK9DFHwCM6HrM/DyCfO8S6v+guYu1hl1
mEjkU8kNhKx8NGOcehLHC2B/KD5efymc1/6pXZoOYkdX30okTIgag5iAyAo984uBT6gf0W8PfFT1
s1yXAHoldXTRVKxSgKel+aa/A/1daQTxrea3saiTDMVohWNnBhsGdNjeI3CilNVlwZ5McmFIj5E9
at+2Q9gt6/kllXA0b2+IdKt7YiQkiZyFEnO+Aj1X//b3jwshrjXuVigDrEIarlEQxBRpOs1VpYPv
KzpGaYb6+uV6TAIL1IdLLd95wmILbxaV4qdbnB8375uhHprw+7OxfQRZkREiBLW9HLh+eZluF3mX
kT2D7rRpTUuxrnQUke8Gtyz/Z1HvaSm3LvwZ5pmBk7YbYNAx0ZmjtjMFIvP7GAOwHWL6LS5JJyjy
WWNkJX+jkWS462YX7u6Lnhp5jL+o/YPNMYRUP4v6i/UslbBju89GQrN3+/QiHg3qFKqWuF92PZlj
VDeD+eed5zL6y6BUjRxlilk+h5npyMBy+vl8VLbcDBGDdVokWCFSGWusFa2aUN2iXs7i61WqCwQw
A+FOkMVETEDxCidOD/WkFiLyUGgfjHwp0DIJDvD7R9IyJurghuoDTTy2GqwlunybjkBIuVHbdnrM
xQCcKSVs/xC5NVu+3w+Ar8BIvC6+5bpmkZNkMDhFQ/vP1nAu2VgVzQUviAveXqzcjFByoy1CrGsJ
XrN+3hZYNd4MF5ENFmlSfsUQJkV/kzZEyFzL8FtWBEn8bTPXGTSNpa6fJSfb7WEiE8CpLNuXBU3I
jKSbCFRNbQENWAAR1N/7lyAe870FD/rbvLEgR+axM7DwBdoDg5ZHxaKsGJbjRz9i56Ov/VImAPoZ
2JCSO3Oxirg+UQJjF1joPVXC3HTw6zy4PImmOEPAUn+u4qAPHv2nSGs0rQFroSW3V67acBqMgAwN
la87ILXcDAKhsvj+6+BnGlD0T3Q4ZMr0kEVEgAw6ogMVqjhA4PHTOTGfK6cWoEwK/3x9uqQejYbW
1QRDZe5wXwDVLBZRpjhXNdQjV3pwNoETmubsftnNB87dWevU5EgZcAOjxyKLd7rNAKMjAoz3Ca/6
yANZykglA6jWJmoqQSNsjWKlSkN8fKzIgMrMUVxzXX5/CZ0Y3/tNAsitxRCjmxampJsaviob+ii/
VyZyBIy2NoIwaX2ACjeVyhxTgZq/t99d1vw8YwVILwBlK57cDIE4ndpGT4DkvyqBYf+SJbLtuzA/
komKkrRNNp7BQexiTK5q3wqTbiaYS4xnSaDhfUOSWB5tyWUDWbx2l9ipQs+qIbuOxCtqtPO6/Io3
s51SXnHIPu+ysdb9oo2b+ZyLXDNMONPQwD1pNd0zOuaehrKPKPmUnvo54hxFdNuOryKjwVxPgs9n
dpo7BqOZOeGdjvqTzfMExXV4WUG04Bb6wHs0iOo4xyCkcseJ9QPv3SHBepMJ7p1yGlZOpawxVDYl
MhS7tjetjaRCUVww3ESDdrX5bTjm8RVCk0PJ9ZyDKSwwJyhgx3FcDlGXp8C0Bumc4mkYGmGFLnJC
bB239x6yWPlVBYKLXiZqyIU0CB5wFNoGOQJmc66+EP1tNQmkrUy0VLBtHFklgr2kh5F4Fb+c4uP9
nvbFTkPU0MM6tlMkHE068aYXX1BqRb1iwXndNwfj0icPCfnDH0fweMB4q5rvROfMrSrTKlwvTytM
mbpBEg2xKu7l6l70sk+A1MUTYKSTJVe0OLsJmJQhmU8LSYagmxxwJ5Oi1luwl81iu/od+eGXWJXO
Y1NvjGWJ9seSJMS0gT0Cy6OcGsG0rPvxuSfWCeNmEtZLfELL88GSymsjUiAM9N1uHNYowThoZKId
+4bPlyVFkYDQAS95t4HU9U65Bos78drKU6OZaxMOxKhDUPYElUJn9sI6e1aM8xSHzySe3HhoYePb
D/SKRjmMbH5G1P6cFDEQw40FKzIU5P0qi8UnEFu8d2PO3CmXKxH1N9R9QH+irmdvQDKhsZpCaeP5
AF9bc6/eIIHV+OYmOqtAnrou+8noO88fDkQm4hxI9V/vow6/jIau1CuTmk75XIXMiBswBBW+K8Rl
Hj7zC2wGwmvju+E6p8bYEBAfENN58lWDkUIF4gfpInID6sHhrlemeDjDEdWl/h+aNcuFl68jRc4X
fCw5dXXHVkYX76zDwu35aF5D53PUwBRuWeYnQS6xWSRj+RW4gInFvdiyRoOHyjH5NrQ9uvoDCu0M
yCUrOCzVkaikTffg6+7hAhCfc51i1AvfHaKltkdmJKHCds5IlffpzrkT2CupcBOYqiHhB3LpVcKN
5aze+KW4UhMXAiAO32lwLN/3/ySwxTLunia+yLvNVo8bcWMznFGmWCCZldRWDCzTzrM2TJRKmT+V
itGgFJmKIirfGMEsU5njmx1p8YenbbM51ciZmWGKwia8EpcFBayAPr1kEN6yjqvqDv4e+2b/q9Tk
o4WZeCxSCinJWuRE8ZtAduvNsOPhYP1qOzg2HYX8BiKEJyPjYQxBR2XWVU6BifXWy4Rw5og32wG5
SUDqFrg1WrCXcNYYoI58Ll5Kk2zILE+i27y9vAYieN1alu9s+0YzJ6G+w1/HITwHeYMoEG8TQLmm
kkrXE9MSR7Skw5+oDIopXZN40O7+2n42GWoOa+ZrS6jxshili4A0FeB/rDOCJLFyenxHvdYKarAr
QED4pkD46/oVO/mF/ggAYbFDP4yzEM+AYulU/33UTfkvhl8/aiiCYyr7Px7X+JtdVfZ4cQn+NRQQ
nx9vnxUmGSToTzol4U2yPHFs1Gzg9/0C8m2kul/bh3+caFdGJhWn7Nin1pNLKmlDKXCh7uhMvIC/
M88GVMHsZlumC2naLHJExylCOGVp6kkXAwG5U+n01RyPZZRzJ+gDlaASFHaaWoWWAIsfcqjTvEup
BR94wFS6hZ19fMW+dFKEtXy6VJXg6/9XNzfh2M2RACHbzbDlDSw3MN5y7n7ZGX1Is8wvC+y5QJpT
IWqXTyJXSzfH9pQwgz9Y7VcK+WCiHzWAm5bAnrzjdkiRIvhl3jfT2UG8ZY5RYL+J9raRkUd9/KlF
meahtW9G+vm89apnI/qgi+zMmBF8iiNNntRIVAvWPlD1yKtbJ0Zn51+JFLxR6tTt32sqi8qx3pY0
OpvGwoad+gOsyQQTFsvpvWj7M7G+IOowgvUQ/CJsqkmOG7qHcNJEb0wnQp3Pynb/ARTVVV1MYpww
d29NjNiqGGbqwXwJfP2c4rmZOj46JsvaOpARksYoC44vP1b7kyn4V6qDyQ8xvt08jFuOiIp5PPkq
u9/77fWwUltaMf2v+U3Wm23umVkEoHImfUFQQRZjsxu8ydy66dcig2UVc30iuD6k79B+bRSmmkU5
WPDPeksRSGeO+F6jNi30Qy4yYsGwH9q04LdtZH1eHiwPRFP5y4qYIfSiSYmnDjs5rsQp+9Xba6FP
fHeMBzT0qH97oo55+5NaILPWohje7aWBudRVwC0v/AQQ4SZF4RSLU5Sg0qFcOg64MgObOk4SmcPp
Zv/KtDJs7tb9/NWqxfuQlTRhoA2QD+RH+y0TIegv0SEc5HAlhxpV/ZMb/2+XNi7trwdJbUxewCW7
m7RjC5OAnJm3vAN6KQGPOwR/FnfJhtMoBleWw9fm4Uugz/Uvg2D3RveV39WcG8+omoELRSjqu9ah
eAf0JY/8q0RosyRS9NE/lT1zziG+uk1y+EdipHZflXHRZ+1pbHj2/6SBdQG7eu8Zpz3t9sbe/a6z
snJ/9Y1g9iZoYmbmRRPzjJ4JSdWPvJqDiTMDxYb4BPNKbkPx7Eo0DzgDpLR3VwUigXweWnqspkgJ
KEqFGAoheZyRFRdLXx0fc6/EvWKNnVxln19bhmWBifK2LFGIDBfZJNHE8HuOHlz4BmeTnKk2q5kl
ENJkaBP0Nb96Dpq53qmoWQGZhBoS5R8fe0UehbiLD4EjMTAzqLPQJZsFtc2GgHq7aPXa/pvYkAVV
7IjsYCirYoFw52+LTJEX5+owZgnd2YXtCz9+CpUgCFCUdaDKiBE1nZXJPHj0zpNKgqrFkYmwp+3p
dRifLKHbG40uLx0Yv/MMWOrjIJTMeYzcebkO3EbaSjbU50gyY2UzWMEUizWmoQnJF3xOku3BMN5B
2haupdj6+wTQaM37Q58pL6El01erdmYXfHrFhdfVmnTR1MTh4A+jbB/bRiucEizs9aqEfc3Mhq/N
uFAECV+x6Rj0SQS9pb8jxoJq33sV/m0DnRLfpaJSpohr/exSuCViAdiDvowJYeGYlzfQpDTfZqVL
YCU79Xfdru7psrp2yA2GmswaJPLYNazrvM9o44RObhoDmq5DE0Eiw9YXtxmwaLK/NccCO0kqs13u
6BOfODDZQuNDh5waf6bnNk1PrWUZCmpEL0WkN1Qi8h8Sw5RdUvnIJ2kC85+4ax0hKegvH40HTRYU
GuNFiW7o8ViuvKKXdM0C4MEgTAClz7xpfoZwiWb6NpPJ7RK6CJ6Wgjcf1qbOkkL4KobC3rU2kmy2
p/tmEbuQ++YI63WhHGsnQQWVBAQd1sM+v9RMS/AxdVfDouBXqG9tjqVTugqeMMychKXjkVmlnM/y
YbV3PWjbL5GCbO2ErT0ZyqQscRKil/KiZcqs6GfCHW1B0CyyafdBFtmgJpzcz6ZuqWDeA+guJr8N
zCyrGSCsVSPuxh7EkB3YCjej6twSPCowm/VzeKMimJNYJqAlmMsDannBVLPIj+OOvulqTRHL1Pfl
JgcAZy0ct/UgJvKHrBxggxaTXITOOrQ8lgCLlUWrs7LAAyXr0eAbOQujWch5eIUnJ7CNo25+pVVZ
dNF8kQCa+SpC4f8z2FV/Dc2K/pakBdHvgbclre94tI7HubbY7kpyUaHTEjdNpjuz0d8g06iVV5OR
gDexQ0brxJG1OGdvP3B0dhmTAe/2YEx2AED34fxzs8PbaQpHkoSVDZvydESLkXHXhnkE3UxXTV9/
slH1fgOakKJpSwLLTCtefHK7UnDiVH8D+ULcRuoyH/gFV4uAWqdbvDK6tZdWMw0nwapzU0Gfh4UE
0wQObBfFggLWiM6tl0ycNxV3UNxhIF0JPk2TQv9cPBjIAyjQhiNtWCOgC+GMI2uJPWlEmVgrVzBE
BXAWu5qHsbPgWlRNyLDnewE/4AFkm4yPvCRT4Oe6ABeglcb5fWNZbS59YU7XW0zY2EMWca7BZqNT
+iFWJ7GoVzbefuYT7gKUONZ5AYQFPH8YRo/EmKqRdHtZtOsrT944Y2q5FLfpv01zs2zE7jP55k2d
rf5wU5ZfW+oG/cBhFO1If8hcO+IgA0JQCctptW2l+QDpgXvbv70MuLTUzS87YTlk3Mfbk9AAGfdB
GZKvahN/+mFImUDjV0rXn4LoG0BtoHWErYQDVrNxPjOjqHJrEw7A/lLPBjMjPY+30/AuviMMSBF2
5lN/Z4H4faaEdrNyCLlaya4y0LlvZ9JRvMYioRYxR+/qzkCLAm7yQFgSema40Bld3/ZSHdU/DoQ5
iukKGfZo9uRUEpLM3hJRQnxW2kqCRbIesaWCaTPdjLMlX5rrmI7c8apwKttfrAq18piTxmDsQqgx
ItslDWPVvKMEAqL/gIHcF4IJhU6ZicDjnKt4+IXRooWRY62MxMz3Lrrp9kxrhXEsvN9VX8mDuGy5
ud/JBHNlO/BBXilnEwUZVp07FFTf2AkUjJv8uEr5ar3xV8MJVcYj2N43/Lv96r/Eu/5G2+sQvxHh
1W2H9wyvL23cv4W9orzmw6mlmnjHpvFy8FtZ13WTNlGTt4FdcfA2iw2DIN/gVlTRZgCIqo5z+b5v
am00+esn0C62LO0tRSiXsR5ieGBIFzEJMEo+Kmw4yGfTA/6/GiJ27RvXh/+DtUSV8ufLVlixf+fQ
CIOgxvDPZ+9DEwZvYy1uguwA/ip/BUAHjmMyXyuCdgCKFlajHVpNh9S6mkLEWk5f2aCwMLbkU10w
lwv+1a0tsiL09m3qZl2i2+o9sR35Fp3/LG8MjamsW9Dq3k/yzSkkwSLD78dtiDkIerF/NJDNwpQr
9GvW/7YUOKWoBGALx1tzPiYn9yOvGqHVVMms30+49571aO0aMl46J8ZIAvFAumnjtgr/xztrchYV
iWjmeT/tzH0HUaKpz+zUn+07PrWKKk133u/X6sx6k4rEIC+eaU3A5KMHg94I180CUDD7A6GJXgjM
XL8voejKMRoGGsoQzWzPtnevODUQvNIiQ/yzJxR9UMzt967w62N6BnvNtoENyOD9EoAe+h9J4LHV
Wo7IlbXNv3j5i0T+bhe/6XoyjFC+icIH/J2vDdrtqc0bl57yv9eM+UBFyegysbDRGRj7ih+tXBPp
utTR7kMOSZvSzdNK9moV8amtmkHgndS64yWAWFhuVg4oph8HORZE9OHTGPgZJfX5GEoTY8xD4asn
IeOkaEwpgyA6JMDvKxT1p7CqfeC3X1N+bmbT0k7JA6SktdmF7xotCl1P78X1U3BcXpThyaUvNCNd
ITty0VnFcpKXxj18avks5wx2h6zwALWEj2g7l8441bXyYhvzhpNvypZUOpn7F1VGpSkRzoR9hfWQ
Ti1mwUEPygBulGqKGx28+1YcqcMt9ail/DfkBYBddclXjLk7wZBb7GZVQ+7FAoC/jc8h+Yg/IvEc
EFrfa9JBq7AinnOaxzLZhlYDWSwaWGKTMRwj1IPixUxiGDcbDpXvL9pmQ/gB6pPCE3PcrsAVllgn
DzTfioT/GUJew4mlVgNmIayRLp8j1PPhFIlZxDBibz+ORtUcSoil4X0mAv8GbALxqsEldrUHkBDb
xkZxSRCCknWTa1cEGJIDiTb488NXEJBd7V7BOLAWmrJdcnZCej3vTF71T7UgJgO5kG8KJYlimWL7
UnV8+YN81gATtkCwqYZcSKDwcMS2YskjHP9uvpsPLMRiW+FK9tnUid2642/13/lRzSTr4Lxjghb0
9lSAEwMz15xC6n8Lyca8y1RDDtpFcxtdquNOBI/SOEXmEwf654u/BNj7ZPPaa9KBB5/FMqvpPCDy
gztGZtay3FBFvkorogtkP2EXCr3+UZUSbbgeYt/MtYehgB0U0TM2/uZekpKyBloWppZYrpJinKhg
p9IkL5xqjJ64tnMY8A9woRF31pFh2Vj2Xpf4FEHPCKga7pyZiYxdWkZ0HFeBd+nVGr/J3Pa5ADUx
zapWGLjDh64seEvcl2566ATXNvuTTLNOcAQxyew/84sNdwHSaMhr++GIap3tF9Z4Aq8nNJQqgQrX
aOYzCSpO7S4a+saiEs90zDp9sjzXu7u5Ghk6e+ILSTQYQ6726tUZ8jWRt5954gbtY8lCPq1OinzR
AZzHu9BFKsOx+oOWXRUl43XeqLKHxC7i8/XPmOEkJEPoBnOTBP+9muRojjfiX7L5bVMLVKYSxCEd
qPpvlkozhRkOx1r3tFRxclz8/BkqRgyUNCaLhyh+TOx8b5eeHEnq2PGBvTsJdS6sfSSjpwE5wR/1
eSuIlo1rvbNuzcwsIt2PDN9EzeEz29s5HWlaF0m1B9SGXMlM0ZSvSv1Th7haucxwg7vhGcyjQ/aQ
UIWBYdkwFlmBjG+rrJ3l+OHAxSDw2V6UKICi3ym67qmKpQRmZcFuesVsuwoOFvvtv+CjMQdSr5iR
GFmGHpp3Yvj+PiwcZDA2t/3Q+bmhY856eJ5NKb5e8isPqBlvMTCgoDXhqBIRDQ2z791P3yyG6uka
rx8GxsSmqcqQm5SehI0DK9OcTw8f8ACwtqZhumz62VCuW4fXKsSgO4CXoFG6JpxY8RVpSOe2mjcZ
HIa828TT8/0wNWHU5XPboG10wWhwkegRkQkgplTRFLM/VDvMx3k5UiBlAflsvloE5DgQ8ttbwdIH
NY2evAGBlxhHI2gsk7PRjexuz5nBGcZcp0k40CtveMoKAGuSZwLQTS/DVgP7NbyOr0ai1cFTXqHX
XwLWvCPoWg5lkPkBpRVNSUcsjtYng6deVBQauMpR9ms0k7rm4ToJa/rfCkUyfj7jTDOKJWLbVKgM
9f6slT6mY0Dds6ZTrFGMaATd6VR/hoHoQnAmbmTUA8Zbsn3FNiZd1gVmYzbV14Zls4v18OM1VOCd
vIhiTIGSChzVZiH/gAMsqLYAoVooU+vVxzX/ITTMxsvi+iR62xOu1ECnm9JWrmNADCRaSr5TS/xG
YnQzgAc98ok1xys+qpev4CPTkP6/OfBWGDYNKC6HzZ7A3rd3m8lU1M+Whhq40HpMc/VWrzIPYL9H
r73MWtwqbJOd/ANHO+Z+Bf3f2FDMnjaKUpJs5J3BoemVBxl07OZc2E5oPiJQdI9+HmdI/t96FazC
1abwsj8QqhPw4pFcVlG9OEn+aLXVGKajaduAwdFmP5H0XxDjFI+QVfRTAApurVdnzJ+Z0u5leYMX
FIxW02FIuPM950E1ZJmcWGnEUI1DT+MlIVAH2CIRTg3XG2P6iLQHAf/K9a/IpDVuGTT6/RpBOKWp
vq+HpxigKwTjl6qL/wJFNzxbw6VZGvEJJBbk9j8/syQAsFvG3hoFO2YXpnRDEFFNfz3YAe8clkMX
f8S6Dpao/qFpnETXNTPSMqExUVLqyQ1UCdKHKd7VVlg/epSvChqdOC8U0eM/O3tqA9gX5MaUWIkq
RJPJkaUgjr9EOncytbVK2HZeys+Ftnr75u+wIvjO9gmziOTjD72G6FoNCdiDJ0/KRC1l0xMo/Jfh
f+riud4MRpZPcU+NjvXaqTvPDbiSKFwjyJ7HbJ/GoKbcAz5Moae8fK7cEIafxwoKAu+rmi57eRcG
DelkgEtL63BClCesT3RfB4QLtsxeVoPccGDDy0bpOn1Go68+ZvJ3DARmDhmX6Hps+sE2mDw7RfeI
oz36ezqFu+EVP1br7ejCSvK4XUeS4Z6r1XAGMhqd9yZDHd4BNDbi51/urm+svFH4p4tPwhl+KfYD
Tx7uNjcSLjKLgkIC3ZU34RKjKpxycPwpn3Fxy2OfRmNhjmy2inWnfrCGPljtjqLOfPh1/8jG3WD7
C5EBDaomBt6UmIJv1vcCV/2V23ti+BqjvcjIYl2W2E0FqVU/xAVvou9HVJB64V/8L9twpRpG/P3x
eVWepxoNrXIk825UawioA5QUv1QyxM4xw8x2NPR1vXfltexFSeB5Zd5o+kmjPkoRU7o096vz6S+1
cprf7vojxzK7xVf40O0nknJG1511nFA/UOwWRhEbkr6LqbFJukI5NaxRlqBQr5ulYW9dccxmJisq
tpeIGvMUcc9cf8gf14E9FrdS86rjX0zSdfN7GSR7Y9fedXzlWUIwgTQhq1qtLmAdafjCvHDLfJM+
Nq5em6RXo0uRRQs/NkVLEY35rtE3EM2/G03EFIQxsl0jThbSpYs+JrbCn+jLKkfoILBasq1U15r5
eqLWtjSrtH7BeiNxz2ot6pGCqG2okUVR43VUVN7zkNUADixw91QtQQpvyWBKrGQazxeUrqBYOilh
rQGtfS8GfrMeNJIhTAF1SMc6z8NVa/vmH7HDEq0TDodQNerlw0JGMOHcRZaikXPYWtO6ApPM9pjD
daHs47YoybxxJeFSgxjQaCQls695UJhwmMpRscyO7lTmimST4kkviKMcS2LknPAGAnePRyTvlgAv
NH3iHCogA/jUE7JbupYR0jTpJzrwURAKcUTM1HDtADP83scRkiCBuShlB7g/AanlWxagpNTA/eYg
L93cKM/t8RjHFUjocBjPMVXa+hP6m64BAt/blH9vz6kA/3XEvnvAiy4a7F/skZ25DiXfMZGPdxV7
sScyEGA88q9ssfhe1MRDYCIDTwNwyYMVGc74Eb4ia9Dvua8HLZyGKXiLcqykfORxQPRZLhvgzBiS
OdpqtWu5Dq5FIWKFjg58pJoIcTRJx4CDGIbB/3acWDI94gepgA3baYJJjr1I8Yl+6IKdblCtxw9V
a6sCprGRftKkyvmQPe2MmO2+LZyrraTcfoCzykjo6f/Kn1TQWySPVjuhBHu2wDn++tG/PSFj3XET
pV0P+bezOV/3oEIILPcbSTDZcLQs8liGRpxaIkmCtF4Kpiic+W1OgyCNQFjkxi2/0CQPwUiKSDCx
Qgd8pYhiWRvpNysTCRmJECpyXn+W++vZql3x0id1dYc2HjAYjYGSHKIpsRBQjseoy5JCup864JFb
KgfTUV9MaWTnKh9cCBA3KV3QJ3KClX78e7NHMcqMFT9rYx+PQWY65WgqLQq4RlQV5z9u/wO3BNxo
7w+m/rrVA8n7GOg8yyMnmD5dscYr/kedu+av7Xx3seDc67b70LW1Rn62c7MS9vVH/IhIiGu9U2eo
HomrfNptIT8LJ8SSoER9O7KrEP9qZmnwamKKLfSVqylhdXPsxsVJm3pK4WmSqDC4iZID76P1zFnX
7K9nefKQqQNAN0W8l3vdN+ve7dUL7hestUjKaI6XYyMV1lYJJeG2leqxFJabg/kplGcN2iSvGeuT
k2UYxEW2G6eNVyoSD9WB1HaBseBS5UVg3ydI5f/ypOA5lGGMbV9txn+X9z1iurOYJYcJUlNHDU5K
7W42Zb5raZ4dAaQXr728zqyyRZ8tlWthiwyM4E7I7ZVSBCTEfsAy4DWspWj/YKC4PFWdxKbUCfGR
siPXuyxldoQDu+hS+5Wjdt7YFIf15oOluNSQVikVy2Zl1y34GYfq4cEZZvm5CJnJv0ZMCtKklOxF
qLmINVgx0ouhIBX6qQIA8nQs6PixiDetWTD+heJzAhvsKl7z45tLCT4KHxAwwED42T/ugToK3Awt
SFb0CCgCZ0tePhS9v0JXNPVO4zzLOyOOJ5fBknfFizTQfplnSlc8MVhxxoY7EHaygitipGNQpAhL
ziDS7XkqYTGLNnCsNXVHk6FMextbv4J9kjsUSXS9DL3nh/IJXmOjujIM9Xl2cbhShD3oiKrdiBrU
XZYEeCCtsjbbLjbsQHGzSYASL7xtNaXNKmVN+hHPl/YBf2TB29G6+eZHhbQ7rA5jQzSZlit6uzZb
qlS6k6ZWqyYtHlG3E04rFWiFXQf2WKStz2agak9wEW3uVC/B+50X4YfGpzQH/io1TkN1PAQARV8J
xV31O8E+tlyGbtfmxWKtaqc62rCZu3R+QPy7AXBtTadipoWSFwOX/erRoSR77dWoC3z2FPfwxzLm
fxvU4cfumaypBjl1LHmhj/zUnx92J0qp8GbIpk8jk3l1jXi1Gk/hgQoZ5ZCcXJpXcuvMmYcrQVAO
QaUMf8u5SvIC2V//+Wp0vZPsQqfSBUHNrb+tisyyMxlh6RlQXK9Cfjn4DkQbuqMRoqARWTPAlVe+
3alImayalhDDpkNZpAGm2Mgv7nVRrEjUFIzTurB/dLU7PPRerXTlUn/y5cuA+P9maKgmF0ozh6Af
xoPzm1s6PxUnl3jiCj4yf+Wc6mKOrcELyIgLwxoVUsvvLVzpqIckmFiQ5bFVUWPZlKAC8E5WqyIC
CND1WkQikfPTvgAP413wPkVgoSjreBYpaP3hXCK44oQXd9n30FYfQDqgDGVoFI4XWZy1wLhMK6Lk
nRGzPY/Hthr1guKB5AF15Gbilih/GLwDrt+bi7DwAp8J0cAbBc4USeAVsQRUFE5MJ807zwfB0PgX
Cdb3V/gxLCpwh3kJMpxRU3CoIurbNce6pOhu76fdfGt7HB3RkIkKvs7r5mHRjUUpPvpKnjfcKjku
NktEJubx9ukJhtTAPAWMb/PHUDP++MsFbuC9UeFE8ITjQiSWCq5P9h2axB/wlDgJFdZwcG4tyN3k
HYIeSXmBenXvnVK4gnOzVW3NyRKoHeuujbfFvVD8A+eZILMAR0kza8YJNrzflJ8NgWK54qPaGKNS
kR1xCLHAbOTp1gMr1S8y0eucg9eMScIYsUJxy88ml5yngVmdcUD96qkazNc1Gelx6fZF7PcgheZs
76UayxY9mXhKuk0buxWYohPmLuDpsRoXc/48FJq5G/EYxHgMHOMnPeVHEOu3Jysox3Drh2o2ismE
tVxpKV9hhPLluU7jUmrKynRcF33hQOxNppb68bnHyb83NSUPpsu+eIIqF+ZBIX9Evy/BqbVp3jEn
kN8/ZmmrGm1H2XTEoj4XMUvN+bk0+IOMSZizSW+39YV66pSr1otjY9Rsxhm7LpoKRPv4Td3QsNDG
OdW9MIsSA+4pWWkhj2QJyhZ70KbDnfzoKEB76KekM8CywZHxEvK7vZZNoUE9bKfzWqE9mdT3LDj5
1r21lU/KZojSzLbcmVwgWZKhpwTomC+fo9zdwy6wbh34sV0DmyH7v/l2oNOIIaVC89/LeRi7Lw5K
aak2KiAwhQEADdLU+d+J8sytPWUy3hszGEFr+/RI2sOtMPMjS/9iWzr8uNaknnhnmOnAfdJ3Bg+l
6PItR2lw3gjsX6B0/iM+NAwDe/9h1H+fjoLQonhGotc7nRvNrfIyINxUeqtr+VCIlBDFZlPP5+uG
T3Sdb8qJRD+olttmXHDzgBIxhgZqwHMdQRlFK2jpOBf16SgdcAExhWNBlCsNwlMfzx0m1EtWDldS
knbrPmPyI+YiIikpElJqV+KV1OJc9N3Mm/Kc5Qw3+768bCTjVUjhiMg67cVjtAQ1C/oZcGqg3xBA
Gqfv511iRwk+lpPiZw3osOxMCALXmZ2rraGl3V6sXOAjGcuwbBXyfAEPnWHxNuLt07SKR6Hf9o/h
7ZbAjJn26yE+b1Xdbg96ux/fmStFuftkrpKTQJxxG9X6yxctgm4KtUyvsAj8ssn3luFNuSIDEhfp
xXytUgNOcuY7CBrqhJNHKzBfLU4SMCFCstafzKbf9r60nn/0D56W3sgPNR/iUYH0CDAHIPzDdWhB
luunXKT5O+ZRidnJMzB/ZKPw33pxGxwunYNkvFEiibfDODlVEX4NsernK9MsU5wVOCtrPf+Ewjjn
H7diUoGoFhEN8bycmlYgB5xgIuiXukwqcPoOOisKH20NxdtvG9tdGshz6Dm4FAMow7gfGlrlnJTU
fGCeda3RovN5YEVTtXI+xwpNxsqlAUnUZUTVu19ddiOL/wYPWvKiRaRxZAKo+Bn0kLDzc1oBBqRX
fC9wI36WFkLnegMrFFhjgaTwDBs1V8SCv6T8NRxx75+DPn0QK7tavwFFvpMOxlju8RFN4+jtgNzP
HBniywO5ySVMMBku07gGIN2czfWjk3CL+YbXimnWu9rday7V4OiLdO/pUhiBmNvjAqVxGO/EPEsG
xDShorSUkRp1ifUheQ0ooBfAjXIxJ+pEX5xP3My6Hq2Nq1BoGVGiKMCm/eLIquiP2p7FK5xoZ/Pg
UgacmQZYffl+8yXWDezorERQj4ows5s1pFZibLiBDmbLllRFyv9sTNeZrPRXvIJ8ODruu5jNt+My
ezDmQe7HxehLKbtTzIkmRXUHGaCe2QLuHqt0kCClFn+cXxrxNpE+pBUWa0m/xo2R+Y1x5TpPzFT5
D+aKWJ66ZhXJStpxH4GRo4MKBn9CtlTE0WRh9NDVXggQgThVH3kI8MBvl9IlxAe7TpmH1yxSbwQC
2BGRs6aXQVPDBA1V3C3nOVmd2knDD4ceK74eu5Be+Qk1cZ/WKtj2nuJk+l7Q6/3QMKThU2wBBFeH
ZWYRIKLY0iVUQAy1pPxP18khOzZFKErzW8Hz1PyjFKBHxB1f6CZf4BiJIn2OwsWmtKzFhypk5NfK
TjQ4dFw2EVGe3nBTN1juuX6AUS7rxabzvM8ZF0juiSRLDlQzMNg0SlTkBS2WsaOPWH9+5iXJD7zc
6nL8eChZSwFJpETi2qXI5kApSs/4s09C2PTUQrfZdU6rQDY9XtdWqE+cDl8Z9XtkcZ7rR04HRAUJ
EBuDTIMD1h08s41vcPLfLyeOpLXl8KdeY7XfErLZQlGi3E4slkPPdSZHJPnS7p2oWXQd9bxCd2QS
+v4DB4wjGGP6GlxkrN+4K7+6ShSoAKg1HZyesune4yp0RdbtWx4Z6gJoFk3438YJUcpoJ7gIfk3N
blSzBqc+RL/LR0PQugH6gJQ8XJ5RlMk+R2Lug8QfIp78heVS3xAq3f8Rd4ZyJwCyEII1h9doWhSn
5o4m4LvfxMS+A51ClT/oxte6WU1AGiSlmJCwh63/KQMYHr4GtQmWN6IBE0pIv12P5cMzu8qq6xg7
h60fUfpJ8+haRcOthzgFOq9n+M4gLWWwp1b9adOZXvWqsHkienj9WRS0dhH27BbXQRsizAerYZ8/
+3zWeHOly4d7Mwji5NW/ozfdLLpFfddlIB8R8q8g+MmLLzBbA40kAUHqHovvb+ZNt8ksDEbRqnj3
pyI5omq+pHwUJ5c+sltEvf9igzASrJbb0FWLLtCf3od3J+nW1mtaxtf3rgr14ECg2wrxOA2ObYU4
R7twQ1VzlmmR21MHNHnBcggrIFFeXWo9Wqb4/g+SzguM6ulleKPSJuoENdSAsu3U5ZHTvzkcScTJ
R/9LgY0a2hy6rPpQIkAGwi8dTUA0WwQAxVT2/wpt1yukxw9TP+cRKWARBHfec5WGVNbPxJVwHLo1
cSs0YLgcxf0bF2jexIqOZJMK1Glz
`protect end_protected
