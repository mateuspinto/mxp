XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��:�.жX��i�	Of����ڮ�r�U�[Uw0�H�d�̱�J�?'���8�v�s4jɽLG�>f�͔���U�LI��ĄL�Y��-b1� 3��'F���!!�_�>>$I����J%W4�����G۸�=MIe�0���Jk��Pş�Fb�Q�g`6��5ǔ��Mo��6� ��3���SNt�jm�
�j���o��SIf͛;`�X�׼��1}z�N��[���I�v	g�ܟ�X��o�4<
��Ba�@	!No�$��:�s	���H�xb_[^peB��gd����x�3mM�$鋽�O��8��ʞL�?Πm~?4�U�t�>��%�u�.@L�m�Vb!�O�&Ռ�;�f#a2.n�����yoLS����({��;6�a_��;�����`�B�U2�ɻ~���k�NH*��<9�?z�|�˗�����,��gU����	)6&���[<�2��(��ā$-<^$=)$ѧkd��t��\݅��-�!,+��0�G�~��^������FE:��@)K�GF�惻E�"�cX�	$�Ů�T'���	Wuhn��<��T����.=���g��������)v�pG˹8;p���g/\����<;�����D�r���Y���Ϫ�������2K�saپ�����/�st	��h7Dg�3]S��@��^��t4��/
��4����	����
1�gÎd�c���`�0��F
���VV^���,�c���n�Akث��b�,XlxVHYEB     400     1e0!�R���e��$��������o�eC탺�NjM��'?�
�f<H�T�¼����^F��Y�!���,����`�8§�X3C�f5<M��7 8�rL�(�㮅4�_/Id�h="�B��GAN��y1��e���F�B�hŌ~���A΅�J0��%oľue�g�A7�#����Ox���u�� ��j�m{I�c�P�4k!�̘qDj��MC��ո�ǁ��?%m�6�0k��DH��_l+Aa8YY꼫%�EBJ"�dl����VH(8S���q>��95���U(9�W�pE�IVZj:��Dy���1x)��t���V��UYj��d��d:^��O��tP�,�P�C���Eo����[��\?��)��6�ϒo�G�m}�^[LIu�afS4e�)�I�b4
`����LAܣj>*� |`��s�Z�,�f�%�Q&Z�X�?�r�}�Ċ@/�.�vICXlxVHYEB     400     1f0f3a�@$�~�训p�MpH�1�����5�	���D���;]��H�N&J����W��)����2W}S�%��W�wX���5�"���m��� �4l���3�5�m[�ϐ� A��y�O5թx�q����晌�#����UZv\%�S��2&"]���x���F�q%����k	l�ֲf���W5���#x��s����
7����Jw���f�6/�a5*x�`p�o���&�}
�sn���!Ù�`��Ԩ��WoS��p����-VjB�i&ϱ��lE����7nsw�a����]����=p���Yr��[�yNn��}U�V�8KJ�h�i�ڕ�tj������p��#c���#�M�{_o�$T��' #k�����l�#�8EZ��"S�������y�8�ڮmi�_s����H�7K�l,��D�i�"�����sz5�F�B%�]��X�<�S
= b��R�����,�1�B�TKA�W���_ʍ�XlxVHYEB     400     1c0ϥ��`6jF�4.:����̄�龶~� ���mǘk��?I�y�]j�d�] aкec�dh0��`MA�^�5�O� �	mKg���R�))�g��7Fv|�?��Q��M+}ۇ���H!?������+�+�U��a� ʣ�\����@�|X%�p�C|1�����SLt��|��;[_�އ�7B���n��	ڎҲ��v�Ċ"����Z�:����>�����)e�2���c���nz2��}����u�oC��9���H%t}Л(k����(�{�IpQ��%�Sgz�3���s��2��#2xǢ�?3c�)����zN�0�1!�~Gn��F�>�������'˛���L]�\|o�39�� �������ɹ@���'*���׹D��!:�!K]�ЏY� K~��V�v͍#.C���<��gct�~Z��cLXlxVHYEB     400     1d0Sr����)L?�
�Ü��ߙ^5-@���w~�`���*~8����Ύ�"�=*����pS\u!���)R��CڑTі�w����U�htmAϠn�4C蛾����2A�y��^��9��L�`�Xm	��,�XvP�H�J+��I��s%�#�m�'��hVtq����LBJ�ը~f�DG�Q3���#w�AeW�\4�C�B���G�N�N`�V�P	�
!W_���EgaI�z��P]�B0UΫ�sg�9y�ZT}=#��v��O�7:��\�Z�{���ڰT�ٕ��S���f#j!
�2ʜm��Z��LM)�1?��TӠ�H�&x�To�l����O8u�-�x#:�"���޹��͎��/=*���L�-�^�VS��p0�Z��ǎW�-�A*z����M��(����%"4�휊�qtIh�qB�8Ԑ�g�N����ͪ��&|�XlxVHYEB     400     200�H�,����v���3�Z�G��@Ӵ��^�yP���f�Y�&s���/F��'۠����h��:?���J�\j�_$��H�k�%Ogݚ6,�D��U�S� q� �G��,�v�hn�K�/�3��A���I��X�Lm�.t��<�$�dUJ!��O#R��^IJ9n��R�f�9����:����H�v��*���Sۂ&*f\pY8��Y�A2�|������#�ȝ�W�_G����sPaQ`ý������,���l7Y[���4gw����2�5K���eR7�p��u����k�HR�{�k������J��<h�vT���r�Պ��6���C_C�#�{�s��Tօ���+}���[!sҀ�_��}����wm��G� �I^g
��bz�4�o��[z\�c�?���6R}�	��,��`���z���R�|��F�J@��w�xn�;{aɀ/�1!�Z��r�3 �|4�w��f�☨�C\�#;�ԫU�ʡ��#���ɭD�XlxVHYEB     400     150-r �ef�����I$��Wl�a0�X;c�����X�\�������=$c)��t	�ACy��?����m�	�����{6���N�����[w�q��Z#\���s��_�D�Yc��թ�y>���^mN7�z�* ��N�T��v^=��+}�k����~9k0��*�E�ώ�O���A�K/2=N��<��""	���2�P>_�=�0�%d�eI�ף�n.0�΍�37h����~�MB���o����%h�K�4+�E��v����S6��.R 9"$Q6����|y��@}qbA�4��b.��w��B�t���!����v����w/gY2d�\XlxVHYEB     400     170A�f<^ Mn�m|]R���}���>���$c@*�[��H1S�����U�?R�w���0��x�c�UrX;9��8ʗ��3tE%�����y-��T���^ �/
��#.ȅ�厗���
�ȑbQ�ނ�8^�'��XQ��F�~��8��j����Q'�BuI��66�];so����|�CR�g$U�pd��sw@>V����NTQ+���)�6�\�b��}��oU���"�ϓb�b�

q��q�l�2��Q�1L�r�_ t�"b�Kߝ��`�*p#�����7��; mH�����p�m �������V�:X��}9zM��D�3���Y}�e����JqT��#��O����Vu]XlxVHYEB     400     1d0���@��H��smN�B�EQ��麩��h>�N�iU~�/
ڈ�>`q�R!^h��ϊ�q��vM��{���f��r��tn�(���۪��<~Ul.bH�:����G4��(��p7��M�o�H36 0gbOW9�3�gA���א��oʂT�2���һ��	�y��*�q���0��������=�SJ2�sLp�?ؕ��@X��І�u�t����M�w7u�ʼX��Z�K�ó��X/�|�YҌJ�̰T��8�9�<�W���{jJ%�T�M��нG>�	����}�H�R���{	Y,�����B�-�p�EJ���%�:�ʡ9�0��(���#f���p�{�l wxH,��d�ۏw^PX�UN+{F�d
�7UX�wt�7n�u���@ԹF��~�n��맦`'@�`S�	o�H�#d~���gX3i{����g��� �]�"�檸mj;�G�!XlxVHYEB     400     190�Ko�Z:�!Ը ^��l�o2-q�j��h6��ו`�Q�N��0d�tc����-�Ki�2-��B.-:x��.R�2z��s��g�xI���m��m\]�=0~��*f�i���]�=�����H6گ�g����@S�0^dG�Р�����m�a&��|�)��������0uV�C�5n�S�L��l@�$l��7�sGa�"�W~�q��ϔ�'r���ԗ�8m��(\-���������8fLN �� M��VfP�%R���G�m��ȩ%:0�	e?����"�P�4�b������y-����W��lS$b��Aĕ�れ���㏮81;������*k��
PJ`O�+�v/P f�rO��m-[L�}���WM���,s�by.�mp��|XlxVHYEB     400     190�����3��\3�Y����#UFs�����=U��u�� n�;`�y�$w��A����fU���P���b��Nǭ���	�ؼA���/���Q��H�r%wKJ�=�����뢾�g8��`v@a�A��|���X|�0}����P��.q+0��C*U�`zuf
��{�$A�L�´�z u�����V��?b<B٦v�<�=��3��9ݩ2)�u���x%���U�0N��*��˶4��mEL�9=�6�i�����z8���?*�8�n��?��g[[2��T��r	%氣Wr�jS}��/Uq��#�mU�=lN%����l��1J�3����g�1�eƓ��:=@y`!<w�p��?�]�� �N�35�@�V��5��C���JI��h��XlxVHYEB     400     150#'��i���]A.�'�I���Go���\�5rdx+����f�������HF�`w(���/G�:��=�_tf�(�ک�C��������`�#�,�ꍣw5y��]��� �>� 1��1�[�q��8��3�ɵ	���>��.�V�����ļM��(a��O�i�p̍M�m�V���(Z�k1}���>�@��F2��\�Ʊ�#�}�J0������v��P~]P�+���T��-�A-���o�oUyl]ׄѳ�e�@�I����%�\a_�����헽���CFUD~y�
� ܳ�"��tt�،��g��y&}���G�������XlxVHYEB     400     150�^�U��[p��뮦UQ�Q�	m���Juf��@V�9�@]�x�ݱ�nhY�W�� �d|�2��$ת����|,8ดžA�^�?�e�p(�b{�x�\��]C��3�(ېy.q�_�OH�_t�ި���˂̯�6�kQ��C4��ț1��������X����������e�?Ao����JHwf�Нv�D4��;��exDx�0��De>Ӄ(,:���
�(&P5����.(��� ӈ�����l���m��,����p�Mӭ��lՔ�x�)kV�d�?9C�PX��
q~L^��BuU�B����^1W��XlxVHYEB     400     1c0<�*'q�:��.b��-!�S�xn���L�|�>)�EП�(׹3XUd��_MF��pt���e��)�l�J �f�����	� �2�_��*h��!�,J�Ȅ�疆r<1mc��0$�t=�Ҥ��&T���E�47
KF�H�bxJ	�?�6ZuvĚ�@Xh�w |5�WV2}!a
���A���u�4^����o�C`����81;�Y�!P��Es���r�_mavf��G�����_�\[@��]�֋BӖ�M_:hg�3�#dE��,�)���1~.��t�1@W#����<�%{G�% xf��wW���yCEƳjc��N5�[I����Y۴=/SA��,*����+���%��6�wz���_��-���lZ��SW��$4Z�j�酼���9WK{���e����PNХ�V-����t��-���[����79@��M#����U�A�,XlxVHYEB     400     1c0ԍ�W_gq�R�ᙊ~$��P�҄WE��[��3��X�fx�(�=]X]�d$*ĔY��f����,9�	=Z�b��Ő��&�y�4��p�����]��Y4x�
j}�a�<!�Z�$ray���w��p���9>��N~����\�H����Q�r(Z���� �ۤ:xGS[}�����)rk��:�J�6d������,��mӿ����3N����?�%0�Ng
��W叝EݽA;%;N�UՂ���o�ik�<Fx��}<�C��U�p��2@.�{�(a�/�}dI�vw3�Qt�&K��e��(TQ�d�_�ݍ�W�ʵ2���3�/�ۿ��z9%Ӻ$Gs���Z�-o*�ySp��Dl8�L9�f9E0�(���`P4����p�p���^H%!t�S��9� 
t��/���u�l� r���2 q�}V�s���@������XlxVHYEB     400     170t�'�*�΄',�s�I}�>�Z%7s?J��3��@�0J�Gj�l��)Q�>�J*�ɓ&��X�9���Cj��[6���l4�����Tn�D��Д��lT�2��QFb�=�"��'��P p\���7��8��%��)�<DZ�>\���,O�OP���F��b8��Y���H��v9&N+���xP�d~%z�h��v��Ok��~C^SP�\��5�TPoA�!/	+�4� ���5��gd�i�)�H�O8P�;3�٨�+x�S����D�
J�7�y#I�~�F��&8��s)h�������Ys#ŉ�so_`�C��@q
iǐ0��`�H�~���<^��bG����S2�v��q7�UXlxVHYEB     400     200�-%]����An��!d����D���=�'aŢn�$<\M-���%��.*�Y��V�˳�4Q,�{�/h��I@���֦�%�S��Җfa5e�+���FR��P'���]ߚW��,ON8硖��`Fk�>l�޹�e&���:O#dO��n<�`8D
S�j���Z�4!y��$A;�p�	��G~6o��_�HEDi�x�W�6���ۊ�ի.�w�r��|�+��f��t�Hn���|�� �x>Y#FE�_�q�}���e&#r�*溙�b���B�0)�a޺�*I���2��'�@���`����L�Tid0�d���*�sA�*�uռB�&(03����p{F�zZܤ+���v�,����cx�A]I`Eu����o���<0W\�u+� 檣n�/;ne?�u�~���.���T�CKq~��D�i��W/l������	qSU^��BI��z�2e��.�sZ�d���W��N���`�<ڔ����*"����XlxVHYEB     400     210|M_�,_�V5�c'�)��h@��s���{�ƽ3���&�7i��ʝt��=j�h�4�P�e��Ġ�s��$�!V{�P��G[���bC$3�O[�!�>�@Mz/J��B�Ki�ź8f�;y�^�5�����I�{���\W��,]�s��CO<�d��#7#�7�|Nk|�񉤪�t��0�el�x�:�QJ�Fy�ج|�K�O�[ĩn̻�b0¨$��L;l���"뚉�[3A������@��CFwe��к�ݤAڝF���2ϳ<�'`VZ�.����|*�[���BZ�NN��`�!�k��Q�T�ջ|�)� ��]�� ������+{
E�Q)1����Ƭ�����)d>l�	5�\W�w�~�a�h��.�`,�j��JZP2֦fܴi�-2����_~/4/8�9�@c�ձ7auD����Ui�IҚ��"�V�J2r�
�e����+��z�i001ea,��ě�;%I>����u�\%�+�qJ�R�p,+h� ����
���XlxVHYEB     400     1c0����L\��2&d���l7~F�&E�L�;�24j>t3�7U����՘*�~EM�
0"A :���j��'��O���%�n1:�Jܽd�$�t!|���d�¦k<�h��w�D�4u��u#X�s�W 26z]Ka3�9&��t��fz�҆�o�~���(T��Fz1=iuX�91	�D�Tn�����Y���[�_�7˶*�ozM����{{B�yr����rD���_g����KoT�j����ݯ],3v��/�t��;O���#\��w�����c��)n����;�-b��2W��)8KФ��x6�I�K6�r/!.�Y�wou��x_��Qc�s	�uWp���Z����pS>����-�A>�v��xږ�k��Y�{�GMԷ��	��\Lϻ�$�@4����_�G�^���]Mศ_aXlxVHYEB     400     160�X�͐f8����U���^�ǅr�K�`K/���-���;0K_)�����;�y>L�B����u��}*.���uf�p��$���Ω>ǿ1��Ez�%����f��ڬ������sҨ3d��{���ÈZ�d\]A�?f�z~L�
�EJ~S�J�����gl#��3�xVIb�*��Ӟ*ݑ�[)9cl����a0��X�U�c?_���j-U�fշo��#�b	�f�e���>c���Y�(%�,Z �]q�����M^�=p7p��2?ܓ->���r5\��5����`�ߞLz�Xi4)�$�/W��t`qq aep�E��%��E���K���Yn����t!]��)�+�XlxVHYEB     400     120�#:�`��	�Pl8[�+RcV9�4Ǥ�Z5�{q��S��Br��ڧ�Hx�Xo�d�F+{X�C�wa%�+�kҦ;��-_��VC�8�(;~BB^�`3Qk!���G��܂֭��%P��������(]��e����-�v�[���=�i}����J�5�7�^��bE��}�$�=J'W���u_ߢ.�^=�T俅��	�"W.0Z5�$z!X[��6�g�k��V/��&�z��"��-��a=����>�6��s
�I\R�������ϙ�.�Z�e��2l'���XlxVHYEB     400     160����>�Z{���OGh����Y9�;U	�;���G�0���3��A�P��̌�����á	�:v�-�i�r�͟�JMH}a�>Έ}���[��y����
BP#@@��u�ά!�C��8�C�f���lgl0����Ӎl�����p�Ȗ�D�Ȼg��W�Ύ/�� �� *��Zl��yD=�!�0ۂdCL�i@.n��q��	D#��]��e�}�ˠz4���U:�g���z�����{�Qx_��?��V|H����n4����M:��X��d'��/#�ѧ|��O��+����'��,3�P�OH�uT�];6�A�	Ȉ[i7����R�VY��&5�B�G�{��ةXlxVHYEB     400     160��5��&)��j��uC>�`�'�̇%�J"yWۿ��6���u'�G�&Ä�!��Wd�J�:C�Y&j�5 0��3x+�L�x���Y�'5k�`��vuG��#��q1��;���u����[X�"3�~ɧ��K�\�qrf0#�4�p�FH�N �P �Y�d+�)�4�@E���o�}��nij�V\���Ds���ϨQ��Mī�]������2�'�X|T���\�������K5�@�h�D��z�sI1�D�,/�H��d]��@�^B��>�W㎹�S,$�UA�>'@?1��B[Ũ8l�-(Q*�N��E���Oudb5�ig���{]Lc;Q1g��ݵ�XlxVHYEB     400     200�z���<ѦK5Pj�'�qqM�Mø?A�ػ����I�*��g'��p���>̂�&�\ PSq6wߝu���	i�ǳ�vk><��ggKC�R���/]���lC����-�ؠD���	�S"��Z�S�A*�v�/��T�.o�O;%����5j���$�����s�g�ŠB+^fG�g���C#���\�^�/G��p��̘�l��v#��ȍHp���½�-_wқ�ÿ�Y��y���)��Q�	���Q�s����o��V~[)��xV{�Iv$���B.Ly]�4�����f�͢�R�����̏W��y�Mf/����������qFV,�3f�����p�%�����=��ʹNi�H��g��o�W@@9T%?~�~��9�8;Cܷ\�
�J��{�4�E��5V��8�h��J@+�ʳ��ĸL�j�p�;�e�8����uqS[��:ޡi��9����9�ޖ���¾���q��;X�?�3XlxVHYEB     400     1d0RH��FK��O��k[��=0�C>/����	�4@����C�����BA������Pm���̖�݃L3i(y�聟n�:
�d@eV�R$��٘���_�؇�i�>B��\�"�R
���ӏ��A���"�:��ԓܯ �"���P�ܢQG�h����CX�u2�jǗG��7��fP �61a�~�LCz�!�vm��BNχ99�L`C�*���M��sS��*������W�nn0کxqQӦ��lp���̈tv$&5�w�� ��}�5�6ܞm�#^������b���d�3$ �e�"�2`_7�qȧ]�����B�y����H�l��$|QX8.��%����-�[u�X�M�
+�X^��kM�ჳTm��;8le�{cJ�
c�s�� P�YBB���T˅���h����	�����WA	��b78�����Y�BR�+�o~F�V[Q�pXlxVHYEB     400     1c0a��+O��%�) Q��=�$����Vr�1wA-����n
Vn�4����T ��&�~Um��x'��%ZL��:Q/É؝/D �3����,���_A�9f��H�W�����c(b��q�2e޴��\�9X5f����R҃ ��S��d'�O��1g�R���b���d �	�1wufD�
?&w���E֧=��
�V,��ɜٴ�Yi��K��� �uꊯ�OuA���+ #��x��WˤC��d�ң^8���M�l��OM�~Hs[Hv��Z9��r�\(�v�73�'6�6=g{�#i����q$���~�H��2zZCq�ej8]�"�m�xގވ}<�QH��c�KN�Zr�~_��?-���^��3�If��ө�C��\%u� ��F|f��Kf�'+�UU4(�Sg���� �ay8A˻�3�F��&��XlxVHYEB      42      50��?����+�W?3\:
��ӴڲX���5
l��S�u��K���޼{��%*#�N�R�������6�`ʰ���� ��}�>�