`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8400)
`protect data_block
vLMJd0T+YjvHUWx/FJZcBC51FA3zdb5QiElvZLIxUB5aoq1QGF6HMzT/SDyttn+yUeifcDUE/kFP
M9qM44YscpPria/4QBCx2Ijls2MTPjG/lkypKC0zu76d6oqq3y+ovSDTJxmuPregOx6UyvP3DqrU
pSVxZ/vy4SqLHbfCm0rZQZ28qjp2d8qiEIUmNY4RkNskvJNIuLO2kIdHJjwVwGaz06cgQszRvH0T
as1C095gxIXv7mWAZ7OQEcOLXy2B8OPiBIgw/Tzc59iYvzJep+u6pgWK4VJ4SPXrFaHorAkuIHIA
ZCu6QUD8EFgbPvTQ+Xqnf37rNfDix6lI8BzUX+/Qe8STJMAk9s4FItw7zy07m70cPrvUt8xtqugI
V/FnmbebO2zMfVBNeEufRa048n/yY1tysZHyroxRFW4dIgUZyCU8ppkJDELyMKS54VyFGXGZ0Ri0
Gp1cpdwukNnBqgC2vARlKXTQSUg9SErjqkPvTVkdifPtBfZMnMSbn4nZKxWFuytuT5xVyfiXhX8i
Z/0JhyFGcLdMMpy289d4LSBxzzQxoipRcm2ZSqyLoT0GKeTYZBrA+YXec4B3SVn9zPM4TO8V/90f
9DZqlFp7bT8wZUWRgMf10IEF71KCD4Cp4ZZAsp0/962t8er3XNXsM94J4JnS+4RzYUiH4WaoiJ9O
TkdDKpR80P9/BLe39PvxPbsNqkHtWerlCmavSZiLuysuurCVA1ND+yhJhZFdfmzI4Eqzpk1pQ3JX
ZtCdiElBc4kSZwDxpw4Up8gShep9H+w+bWJ0HEggihYs3v0+FTy25BkhM/kJ+30OfPXItrdTE2zw
JWbkEKNxUhm+4v0du9Z05v+rcyb8SxiFe9LpwpTCeu2AqrGjTGLrB9isI4LtLUoRa9x5ARdrI2T5
weya0pJ8wz/klrzaq/khHwN9/4gpfdwg+cEdvc2Zdkv2IszPAD71FUMzKZEbB4AH7TgnI0uDhGDL
XHk/z/r5BjpheK5GVG7lgxEtcmkU0Bth/dP6wzZ6qs5Z9p5cUOEDJxsgkA3vUVEOL43xvlhi2NjC
qUWe3ja0vEIvjEQI7PL1umadsX0urzvLtc04sN+XdRSpasWL5p9DeUpYRVbrvarnkeQx1ysjGkQJ
FmLQzVO+QYJFHV6OhpJCZNRcenjh6dv6KQ6MEA7azl25KFoBSt+EUC0OmRoZPIcKqD0M9/itTrrc
NELU/WXEWezEXuVFkdJIuygkATMFpqaf+C+TtQWiVD0h8kpyiLOinrxnB6zSf+uZIvyQrW1gWNf/
s4D+ly5Avnalv6z3kInMh4Y+t5M7DFV+MgW/fEO/TdEQkK1H7RnTeW3H6QNo4JkC2YZj4Fn5N3eu
WDVsfWDsbZIvwcHZuu7oP0reCEbQNxDhtXrjkAzohxPGH/aNaCvi+C/b2lELi7U2z429GYpnOfz8
xaadNsBMNHgUuql/fMh55rzWrlteJ9r6PSSL9znaDRZn11ON7WKEk9r9aH+deF7Ql6Wg/9jbsYax
0fLS1EMyp37bRgyP3imqHuLVwfV7amUBTglRvRQmM2XXd5OmY3Sdx6+f+6EceoPU75DW78tWfleG
I8CCsK08cYZ3mGkVj39YfFkKTn/MxiD3Z4dL4vziyx4Nmxf1eGggi3mie6Q3EAKy6IanSM6BJ3Q5
RcHwE2lWlYdQJASVUaSlckCEZ8H2Xdcgt3AMTLZejUXPhe9VGrsahbfxDHAPfkT6tRfeFHaVkY4j
ua1cyVJfeKeX7xC/dBLU8dNZOq+k0t09DQ2WAiIQ1kDQS9/50pCmgClqEK+Yljne49/hGcCffr1u
CEYNMOpX8dQhUdkV5UTVj+aP00+5lNCRjVySPv+WlFUC9F5fkwhdmwDsCEx2ZO1ZuMJEgwq6iVCD
O/L7qyFGWVeawlg9J7HZIKvZnj88Y3mCY79NjsBC7LkdOVC7QN44NezLww04pIrX/+QiWqtDaxcx
t9ibucjTijSksDAIHtSjHspf5ZJmtvK+lnzwkqwxqP1fzJylkJdIDrgxf+JSYp7bW0Y50KVW/7V1
Kr1uNW5hH3GpGTwAIKK2/64M2PZeT8OuYNf8+P5hhBgy8+F4nC8s7HUUkp88PZkgw96E1VVIK0OF
roB9vifCoeNzdxO73ijPqR45i5Gt6TZ26/ZcOfo7CnZN/D6oHSFZQ37XaJ6UYR4L9bavXpCG9pLb
ShhmRkofdIVtkEMHlWWAR/EKXZXyAZB2YVyBUWIosKcVVs+ti6NOwEcGVTFV2OF9WiMBy82UQXJ1
VGo70Pq5OUJIOo5sBFXd2FU3rCWl6drMvpTdUcF3r5NThIfsugoYvWgKShgee5WKTGGQcDLKyu5Y
pQXiq6SFgaPrg9h8KQe9TNTL+WBJD6w2kQ2ut32CgvdYpea5lu03V4Tg9KlVhOtux3Q8JkUbvVbz
qv+RsgLOTuqXHfDIDgiJodjVfUukUQSj62dEKyEB7W8NHcefY15ZBTy/O18Sex5iCUolMW8K50jP
+v7jT4jd4nSLLuioIZchf1hgzid4feykDnA6G0I7CShfejhQnX6EsyMXlkuMKRz10/2i41rZaY4N
BVEN1NuT2ytK279Vw64ned95JhGKdxjbLMZbYkXEyVIcwgpEjn0nRhZwNGzHvbsmFsS+Si8GS8FG
dwbRgmXtfNE8ybL7wl/LAcchLZfmw/Wd8NWsdXVPUptIrMylT7YCv56GEyKCckam0sOabwlqnnYO
AWbgBS0xGdV5zHqbw68bS9nct4FtSLs2zXfQ17IRMfUn2+3rzzOw7SJ6dJw1u0GnrZoUS7ZsKF7A
+cNQEmPFc7X2EStqby34sPItKomeSyjWtrKSZVE10VkokOcV7VNbz+YuQuGS1MmRtSAssvPsQbwc
lf1VeIu8aLYTf6bhMLWNs4RD7bLB6+dlj3luh1H9TcHoXVge55WP91Nt7lZHiniPK/BTZ/Nk5hoB
XZHbn8bfH+/Y1q3qZbkoJiGNjfqJFasAG/Q/slDgCPZi2i6HQA2ZmQSCjQYHMh9428GznJRtIQhQ
D8DTDucY7nMyYRanHxL8KjZDtncFmlghVPPEZ8wiAOo4jlGhcUU3m155Kx8ypgl+OWNyNdh1Va0/
7nDx+KXqlIicq/jiaxgDNWHzIP2hBloVsDvQtt4kOs8fiFu4tAsEB7zOvHtUq4pZroXc+NbsVFky
gPwkw4QlUvFUWmiJk0bdcZ6Expj3MkZg/sSMsMA8k5nd9NqBKxN3vZmLeO08p/yKHRbwKO9Slyei
uB2CFAqEvFmgKSiREC6VNwaZgRDuG9eunYMCUrVBZxKwcev1qgzU9QC51zRKgSxwwp8hqx08tzsw
P35mum4ra14hge0ZiYys19aAazhT6hyxHlPDdAa+Qg3S8gdMgUgjgZQR/Rt91J1uWHbDnpmZiROO
XPiQYXYfXXiEtksbWb65I0gS/7x5fjPJvM8Q9BxM+b1l+dwFrmU4cn+GON1NUgDxmjbwhil1vD/s
udYXx6dHowJjGyTrgah/72eAZdotPER5P7lzlDVjhH2tF6q2VsVxL2CdtzrTwQG2BRrU1Dp1hCEQ
rTcbUuoPFWSHpWSh1f3RqREg78GCSBeUWKYJyNij+G0Efm3lw15KmY+HdZZIRap93LjfdrvxGZJY
9R/Yzu8lVTS/ovmELEeqBfHxFmTs9xlaw0F77Ux2g+3XkpWTuFC7NbchFGe7KWIGBxJsHUuefs2O
0x93cAZD6tqOont6l2JEJaNERijSahLXa6orT31svRgBxKRnBMtHYhq6/ug//0sTBIqFivR2W0d2
RzLZB8m4kV/Y0X2H7w521BZAV99B0nCnrVqPLxnslTuvUt6gDya2ePvcBklho+QBfExnuM5FpmWx
MGnEkU9kiiOh441MQyT/a9zzrfd0yeiS2gPBPR+WTbYKxHsQy7y1ki1zzbns1NlMURN6qwcTHNs9
7g+VImsyBjJuaPWdap5Ykm3AUWHmrx9+y9E0HFgOIeVdJBQAd+k14FLTUjAftdreb/JmbuPsGcS7
KYhMS0iHkyQdYnXP55wEDYAKFg0hKyMcey3tWzrU6jKRhREpbAA6y1A5G5O13I6C58auaO9jsu++
gAULbPeLeTxQhbglClFiM4dpCCr+6R/3pSk8DCMP3PS2IbLbWTDIWruImPjmSWXKFs5qYrMWWn5P
izufjhLwHut1kUpw66F1prtaBXBvBWKgINLX/3pN6fCBOkRxBPIlJLYtKeU2sqoxaI6HZUjElAaB
zNeyfoqmkiL0o70RidpBokN98+CCsLcXva4yTX8oNxFzIZmjsin8uMdNrxqa/ZLRBYpnJR5Qeb1O
9/rofiMcwTyGV8xAIjpTorv4ZB0mhno/IIoFqHhChMg3teGYKSEBf+2XvSfnXXAvA5JrNNcrAawh
uWGWfIuWxG1dIiMQGW27EEfFhTTjQCFLL1zQ52TOie9EnrfcAf+GorKKsjqyD4ApIkfansjzvw9+
cPTdAAIDKJaGmfQrM9AIIbe6rS+DXzXC+PkbMclOrZovX/hl9qPz4od0LM4ETj9/VctF7/e3V7DY
C5j6lEw5dPTTIe7QWVpZ4AGY2Wj7Lfn7hFkDaNumydaXtAo7ed31rL1+7orhobFZh3gL7+rk96fO
VOoqCQsfpE9d4IDcibnUkN+Mp2J3GyIMmgh6LX6SSjiDnUVDEZmmZFxXbX5zGEczxkkGaDbznrJu
XMgE8qNm/BdJ9NCm3FDne0HOfcBxk+F20QbU5eBxyj7J+JSFbsF2G+woASISFMGmTL2MtcNIkQa3
So4VXMDmuMzHyXpH7Sxrxk7ch8Wd2lrH61FdUq+qUfAozmEKCC6XU5ZNLbiApugR8ejlDSVlbNjF
bKPA7UMblTYACcLmjTGRLvsrd2EC7llJbzp2HchY0Dz5pP6E7lJyHVraIt8s0+8tSGi93zNyVjC5
sBbsHu+coDsggRlF0k45ivwPoPGNBLspVVeyd6T1tPpn+PUBI+MdBQJaR6b79LnbeixqftUnquVR
Xc5tcazGHsIoHTzq6Znoei6WpHbYn8Wqb24L6C34p1Ag7fquMm3KlKtsA6AfP4BovtPBVBfSBdyK
cT4Yscdy9r8yn6G1G7oKlYz/60jwASNhHpWyutMAfTeRZUwwqeGgjHEzcwvbgHxcVdG65cY1FumP
H9EZ1zmGYHJ9jfBy2IOmUtbInMIg+ropybXHdVw3bEzSAIRVk8jyNLhELV4RRz22FnAmSL+Q20uX
OIe2E9b4ASR8R9NBQxqkprJtdMlolh10YYzpvSblWVTMaMQw96m5asjvjTfTSDELEHjNtRNYpRWs
Ri5y54tD/6LhqgncuOnELCPowBM5KTC8ylwQK9Eo6sAr4Pe0kp9ZutZazo7W8BlaQ1eLE1PwieMn
fRgdS11+HU4/vho8q9LpzuT7manv/XTBFTpCsMQWINmdP5oCr9ffgQqOZnHFdZmZcQE6Gm77E3ep
RUcn/Henfni4z2aD+15b4QPb9EvEmBVUkLvgv6kzj6KrLpZ/vuQjpPfmg/gZQtDK7rg2UZTb0lkv
QLeap4LqShWPQwGQT+0iCcSlRwN0gSr3bBK93cshZZiDp8G4sNG8xpMIm6CPDp2La07sjMZ9TCpF
Sr2TnQpSLtc9P5hDCumIalqKEC8VdCAcUzq4Nwsun60h88TFI5j8l9a7bLXGl99M4RVGVvNvqxxN
FDshWLiuNBtnvow7dGZEQy0220Wv/jA91EvCBZD6L5pfpgCt2tap7e03qsEqXYAylBD2Y4L0grDl
0b2Sgnj/jSwUE2HfR+g0RPD9/x7ySbZVltCHJLyo02t8Cp4D+ucm3bAWygjsBJQ0Kj05uTEc/aNO
5qP3oup/kGLldV5GC2LlKy4cK/Z4Nrq+gfVFjOl8YKoLPhYAF3MrRxDXmIu1HoShmB3azy73PtR7
Q1DoqrSav24DzS1HDwxpWxe0uDMyS0vSueLq0qwscFwAj6LfIcBkAhyTGIAX1C5qeNHQwRxVVPVA
VrvwRijHtlrD6gBcefQ+QeG7kuyIxrwoYHeseoU63DZ5WfH7CxBm6+UEcjmg1vjgWhi7cpTZKtsn
aBWcfI2L5gtUSG9gtpQVIZEsmoXfOSQlfJ2zrgvDGe7LyzXt9qJ/cM4XKUM6Zmvfri6CHdVEzwng
/ch69vCbPl5pXGnEeqXN2wAucEuEffsstrF2Uv7xHONvw54Ekt8SCmOPNNLgg8VJK5ziqxaAfOvx
x5BIXb73JK/8nk9PJPNzwD/TPBDlhYK4uyGlMFNcnyaQtFy3tl7uVcT17DtLoA5RLZbyKTSl8Big
NaYlwtFBXWrO2HYEzFgKX9UKW5A4J38m0pQDtK5yc6Us0Ze37pC0aClzTs0zMiDckFFx5fsmnIkV
c1GzhuN+n3GaATCkbMAtHLPdR7M/d5r3E8Cc+8J4YfDa1hxZ5ApVS9jUq5tJhx2i1bGQoUEFDYJd
f4er0Ly3I3OHrHx/bbLYI91KPppMejSqP+SBwrwWHRG6+XkUgFMrwrnD2TmZwo21YIQAQFJloRP0
ppcqqEyUUFkangGAFJasv5+mhxc+NFe3NMOcQx7rDhCxyj3L3ehhUOQZFc85J3UDmD3ZxpYsDLvQ
B9Wb05b+hw5gazGz8s43nrPufmmF6wgw3j/6Guje+bjIGqWac5ja0m0AFUO02hOsb7xv6MIEmjRu
2HVzdJRxua0enE3pek+1XLlSEg52/H7qpIlb2yq3FAz3KGN8ARi/hJAVM2iV9QWOf2WBf5XX49os
KP28VHvAKA2HNJ4B73sYnWu7Wc69L7DkFOh6h8ugY3vRH0awITfcnFCk7ERhMjBQJuQ6bjsTN/so
qJrR6byVdYZCjbB9PbZYRWsER2bAq/PN7Nuy8YLGzmg9qNBrapJXkvKhVm1NIQ8ajKeiqEIEAP0+
Y3W0kCXFbsJjCu+PUzaDcrjQphGP16pKcYW3i3mCZc1LbCQO8UsExnMqqqvD1+5q6QjeqdzI8FFb
sTXHZkwGoekJFoDXit2fvfJs8EzX/eYqbNgE/fu9JJD9o7DiS/LsnYvqn6UT0xzXttI/ktDQFY1p
GbkUl1U4AVoBRyzypMTugj3H+Ribzmpq10rQ1EYsoqkThzRWdv8RPz15vE9GjQHs81lyo/pgU0y5
6UZY0Wq7v0qCc/YPh/c3NMKrcPeNmnI3llJ+2uDQQuJ4OyksRLAQZF13xf13tJYCUKboJZgZVzBh
GR/uZx52idiO3AnSNiFzxD7I6askBTPcOGWffixEtc2ZckaaHcMnHe6ow1XKSuGKJRcgvOShNNys
EpYpCa+DkeFT+PzULFQt23lY0AhNBhlTUdnfPgT8qWtOtw70V/ymkZpJ2i41iu4dp6qfNbnx1N8P
elUyku1Oup/4B7mJIGZYWSNXa5eshMQkQTrwAuPrPN16dJlGAeN98wGUJHeVfwfUfwRxVVNzTkS1
NIWp80elOzjiwKfl2+0Z/X7cUzdCDyA1FMt5af7QJW5wRGFFlTt5f4cHjJS8J/YotiCwrcchHx6P
ujw/NhvdbaJyjk4trpFONrSJVqjVZjgxaH6g0H7QzzGg2hFXOfPWiwfXjXVaz0GwgEj5LvNqwwML
uKu+lPAGp+Qgqkz8GIFiAYKxPKoBE46JAzmXiapgZ3Hg0tfNty2VXD7LzgzNr/UnrseeYq1r3seH
MOOlKfZ6UNjpiCC0nLz+wTi8aXf04CRpubYmMV3ufoxmphxduBfwpugzBQSakTlERYtqLjupVFgZ
nrkln1Us++l1ZLchFaZ1+mFsiwa72217Z+1ELOdRrl9UBj73GAFLED672Kyabc7ALRmkZjItTMot
UaZbRwWZFYNyrTDrPx4OCrQ6/noPg09oFk5xnGbUP6VOGvQqVIYZCP2+NpGGezo9zmgwKjDsoxqO
2PP9RjobjKeYZ04GocCcxxncR9L/a277CVN0a7eMFR0gJJ8K32MJknha52TP28s40KgdKn37qkhr
BSGiJ13/YU5PanTvgPsxJrFT+3gK2VkgfDqx21LdCayQul+E3tM5T/x+Tk3KbyenDKf6g2hOmBy9
Q+/Zd5KDS+NZJhrZoGPIrvJbFVBn9zWmJK1YdM0gOaAszG5SevU7IW7ed9Mk/Pk3jO1sQlNY7dRJ
LkqEjk6WCyK6xhv1LyVcKV4RC20oIvSqabkcT1x/VhetUIwUQ5ZsVeHdtGcjENFJ5LpMICBusWl+
rrYyoA7S3L46mIEdthwVmus8aNb6E+8anZOtxcgEUrsNjrw7W4PrJa9al9FPwMb7ZLXI4/qaXah2
LaEcVfpuQbUEZzuq9TepGyXHglB4xfDGP/ykImL5Gu0zvwZwFKFl+UMrnawrPB/Gfwq3Iv+mWucU
ue+hRf0R4nkG6i6byAxwB3hQpQ+Ep33V9BW0yACr/mMi9s0zKsVubvOtp6w5J82MqDzZCgZnc32N
2PKnpy6HXEsuOGUD3YHHNxnoCasgxvFbJJzK3oVeNNDy2aZXwNXuQa2L55K39XCxCY3il24tZ2bp
4+5WYJAtgbTTFYNffnqLrF6ajFgR2Td6jIff06eIpWL0TnzlMFmuhFrM+yS02qC/5GQ4glReETjD
IfDk8eeJZ0fSIwo4ZDMR9cDXUia4P/hV9Vqc6lXZJphFqpW7CLaXQnK3vKHDF9HCztgAHZb7ODrq
wRSisF81ID5EKzNvGaHWbToJ0UibW6pf4R5jPD286ucBy8Y1GPFu/zVkLDaedMzM/t+5czAbm7K0
vUqsL6TS6iAsiVGQWQ/XIJVz2zwZAFfUyrXg6AIHupnADXXR6NBxDOJ+I2bmBMRgWM4xh3SZHGpe
2EOI9KiXyxVJyVeIlkHwNNo9j26A+P9dGxh2dwQq62oSPyQcL9aGpLgFWGxXiRz6rEEvJi4XBJKV
h8CIKx1Edwn0AZrg3fnv0BC+EIZulWFiZClfWMgcZBTtV83HUY3iLbiOLfpOUysgX5Gl1aODsG71
1YAxGQpYj0Dg/q7k++osUQuqZBt0IjM6awLMETKKdITJ90B2+JlWMZNdDB2gN5GqSQ+AaMVze7jB
0fgRyZLRq6rmcOKVT5ih2YTHkDqz8MnLQ6oxOLqPQFPQIl7nl2oF5LgE3IwutBHFJPR8Zql6UfsY
jQDShn0qXFVaLxEDc82ATvdrKVF35vDLmEN+YkVpxs1WNK60hSV1iKmjL/vmPztfacUND2GQbhzg
NOP70GS+kg010GUtXO8g10KIjOdcI5wMrmXt0vH3GNb9b44p1AeS0VrFJ5Bu+Pm0BOAt6sw8YDuP
Kdm+8Rqdgab6EfdDj3GDk5KaJyaoDZQG5MNXV5c39/5vNz520x9EYFQ/WlCVKn2IvlJkDrUdjoNW
Q8D6Hq3q0jAZdEjeE5aD97S4UcRocO3Ok4zFdvz672YlGAyO7NlH2GPX9vZ3HpH3dVHJdI93hdYy
0Y5CYDVQW3F3DNHVqUXjszZiJRlXOqhSdZPayHFDYgr1d4MZUB2MZUJ3xnjXixxuSc/0RnQ3MesZ
axHozKu/Ym5fI4+fHUj8tCa0TiOheat5bVazBNPUGaoCDJPigc/PgQA2KnVeGFg+S8u6cGSLIft2
F6PM4vHuw+rNhd8VvJsrByxD+th29+ql26lthArYJLQHVgMVxh0YhMwkCRJ6K3KvSciyVQWuiBsC
RX/gb+ICcaovMlOrZicxQGB0ombk+gXG7TkyBP2w8ggrWs5oOgqUFTSunxmtVhwnwMwTBNaWVo9X
OCmGxgW0wMFrPuFzm9wLiHXwacZYbU7UnxELez2PC/RAsx/u6HUCvwP8hgrnZaP9kcc0K+Pd+Dz0
jrf1zNS4aarzxtHqMURu83G1HYe+dEzrjBF2Dg7Y7gSzz0H12jb2seb1VLjlxn0fu4ZCD+0tGe1z
73rzglIHkoKrDn+EoFEDbITiQahTGWwT1RSrEHjGIWTpt8koRjQPqm8mgPykWxRfnZju0D8E2hu9
u609Iy3sW1lkYLzsQb3jHtBlWkKprMlwGwr/BHrQWGYt6+9Mc2EUAI5ya4idyaVQ1bJHuWoqvoVs
bLDP9BFqLaex024deIbIRltEW/o4jUSqauu9LzWgPUn5S212WGQfaMsBMeOwPAIii5uzRw/wGc6c
R68yywbu2U0BeJhsStpkhVXQxES4ikEe7MXHmTDXCM5T4LWsbFwji+9BhjYOBqNiOcTrBmaDbkD8
SaRlcsDf1oeN40EJfb+ooDNqKWD6rjc+K4fJ0OAyN4E5zx52eyaXHUdx1IE8hOuxSnMjv5PXM7CO
MWXjFmNXxTxEbDsYRQuKRrHOblvW/d8uJHn66iTHpIL/doZltOY1BIcW550CmN1CWqBsmDSXyUhq
CtZtwOsekLLKf872n/alPAywVk1aX/P1zZ7sxXFz0EdolY7SDx3OAk6Csz7K6aMjJRTTKkLDtVQC
Z0SHfZjf3/4JBwpnNy7Kye5g9R+RkR5IMo9WaaGlUIFrmdlk7iv3TjYSMSMlvJpr9CFyYE25GwJV
RJHtloGyVZQzm3UWGBI9kiaf4TnO2x6d96kwJ2Jb9QnzLeI9l0H+m9BjK22UinNIUoWm/DPgrd76
VufUj7cR4+H4ROuhVS5y3gyf5xB3kBMY6Mp+HTeN14C67OA1BftWU43fCFTWXW2u8FbM5PPy2BIj
9qBTgxcxjIXNcLhR3WVMc3JSEgTF+yg7ITZhFPlYHJZ2HrmMTP5go1dsQrQ2lA8QZfEZqSsjtaJ4
2KHOEEwh4+EhVZ6VvQAX7m6ytQOD0PfdNjWfnk442VZjMUBtDJHpZFygWy4queYKkZ6rmuyARa6j
uETs0gfba8klBwyBuSxEtZJgCYRvA/r42L4nssrOx1cv3a0kj3m79cvLN5eVBn1KUvn9Gj6pikk5
68IcdDqpYNt4kCzpMoCGLR+6FW+XQBq1hvsvcYQrDtgVJAUroUJRo9cZisCb8whvoQZJw02COH7l
MvyE7pNkrqGT2MjTK4H2458/u58HMPttrFFnDif49VoDnt86n9jpFsFZGwW3+aMmWCGg/bh5p9xp
TliLDyBZRI6PSe0pjD1IfJjZ8YXWpIrypxweZr5E07O0Jt8M+OnWbNBJLkuql542QfhWgxf0ncFt
svPDoP1p54tEa4xyhR6LTKeJNiu7cZkqLqymUwB09WPK6+n+bBJiMFxX7+yaHFdfiq5FA1cXrubh
LEiIpV7mQYRsEQVc4oNSwJx6Rrax
`protect end_protected
