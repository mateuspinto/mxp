`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11824)
`protect data_block
tDVqp9hhUZx52CzVq9IlJXUpSj045BAeFAzxXPGCpRU8MaYPwoiFKI6M3EaeHOHomXnZkbAAl1OQ
zD+tAaun1lK+N6Po89N0SuQs90vAYJt1vgaIOXc8YhtCsdPXNUO3/jqdRRKW/zquSgp40Fmi4UEW
h5q/yIZOD+oQW/AqXUa/T8d62McHcPLjBgiINL+zsnJ3bYBu2FwMUdiLmzlqnrHS01s8n5jK1Ys+
q/wq7Vg5NroostxLCLXG5gay+w6+VhNiUki1qAywl0wTga6e+7jOCoNCNuBuYpeWFsgPpk5kbu7n
NMB5eHQyFyupaBSIQaVjDqZMJhXUUsg+qtccequDmF7YXk8Lrg7BM5YYpidX8yse8G89eUlpDwhq
OOnDXALSkoay291SWp/3o78okVuLkaCKVRTE0Y7sUZdXM7kAXck0g6kakW73MVrwUHcFE1/bSskE
Ae7yeJ129vWHcP5tXT4mI5f/NtGKt8md4/fYjjRoqdsllgh7R2kjoJ8zKi+rjMy9cYgC5rm2YMaY
G3BO4Q/MKJZp4R7i+4dd3Lho9R9Oj78U3ZyTxwccIsBTHsI22Q6KbD1d62JFG+gIPpbMpGLXM5l6
DIFQBFgBIhJPOYhaf76vvpVEEmYF348Uy4FW/7r0E7XR3ELs+425p04D5a/Qty6a8UBIGUB00THL
SQwHGbdMX5KuswApTtaUX4Pm859w387eruxFwrFxKeiWgTbnLHEm3K6+EpFpHHbmKa3x1HhdbehN
h5CXBdGEDMbXwKZp6Pw9KmTmOckM8kMxPyj4E9QYh5cpHcOB4zUjgKGVBIMbQ86SxGuFSpDjZ3Sv
bHgxoEEXyx8clKXzUpHvqeS3Oy56JUSNz6eXGIcMVR+DmuFS4BmEfhCXoWNrdV3ws3s7rDgcLxHV
xIBFACvTz7XqKioeERcfnmY9uT9Wmv/jZIYEbs8Ai+Pj0K5Lzihje2/fccnTpDaTbBoJZqkrLaDp
rULicM3NB5PEqba4KWD1TdlNB1nbx+wG+H4afJp3X+uKtCelt8o61Nlf6Dvy1Zk1GTHQO8hr/cDW
tXzxupiCO3fYMXLJkE/PKLYwWHct52mqAaR/lWl8KEHVSVRgaza/YmOVHMT0UszarF97iyLwNQKl
IXjQpx1NXglNIVFfK3cfqrvdtdP6GL++Kn00Gac7uhsA9oehSZz34/MrRWkMo/Nb0c6OUcq+wHzq
2Mkro4UBow71/ksxBUwm4L0lFwyCJGcLc6quZbfZEBuJEJ90Ro2v+V3SrtwPEI959d6YrYWMw3Yc
jeCA1VFIZYYYlR3rp8U2lSN21B/T1Uq9N1hiR1ywyH7YXhjp5zpBdwbDUe/ZsazUBOBjSRIzoBbz
MdQLxH5w+UKHMsO4brDFGx2pBRjY3HL/l0xtts36udRwKS3P6y+66FsGlu5fzPnT2LDtiANlaiIh
JouCjAa2rcqmAshLiV4ewMykUXLp+C9x3AekxfXrYE/d+I4kdo8r0NB3Ri6xxd2/wgXgMBAJ9SCQ
tAG1WMtl2XzfOG4/Gifxs9lnaVSmsvrPpNvBTHpzoRt4a8XIBm35Ly4iQFV960s/BSXwEojwM8dd
mdSWLeqj5/0l2bxl5u5wqu2ryNiBZzm0cFOjLypXLmBiyw4xiMgduLFq0DwHpOpLdyslAn+Y/jPx
YAxK1c6XHVTx3lUlrZZgsYPvviVkQkVbt/22e9NBnd1GlODZF9Ea+MGGS0aC0wPHyA5srflLL7Lv
dTCvmBF7a7yP4TJMFgMEE5c7N0oX84F7xccDpXkKNP/YLBN2Z2yMpDP8sZF6uWVW+azOo04aoOxf
vhBt2ZduwkABH88q0go8kILWBzlKAjhdr5iFVv46ST/L72pv0Wz4pAiXqyQOAXnGfWUk1w2CkWZZ
HPl3uURBxDISz4GKRTnS80/aJhO6FUO0kokLZueA8hNSiFROfduLy5GPyKn+ao+1zIa1vLfY1mIi
Sv/7WqceSwnTFa7a9rG+KqyLIeS947JGmocqzhNb+Mwc2rApGcCM8fS8wEecYdTQx80lAseW6bQz
PFrvShe/MnOAyoW6ipcqZ3YK65unT69JKvWmHax/Ml036fcoajGlOwlYHDTWbNFR6UCH484c7mbJ
0wQWSoQqhJ+epYNOUrcyTaAKUM3Ut2CQOmsisTlhjfaQbTb+OvhGEBbpWr/+0m56cBWT18FJJHkq
eqe3vQm8Ig4DiKrqCPp9OE6aavA0wlUjS6ZrYwygzb/16ENEAJPJUdgsEr92MWvySKvI8y4DBNTO
0VzIE4SoLbdBPCpeAmLC5r3Ujgl2AXiV12OzoAUf/IJgJyeKKSq9lzcM/4pmH6AjKgxiys22m+v+
sCZKctrklBjZKxvd0Psbi8/thGtt3Dgvt4pZj+/OUl7ZwTuvbk+8ZHv9ms7qCUcSIKuhuHSCkSq6
K4NulcvyaSRIkj575pQclv9J0puItv7w0DFSN49zXacDbhScjy6dXBIDR4V7YPxekyjN8RQuvHxw
GK1t1FIMmLPDRXVNjj3IEeCfGfR0pvm3jpf2vHLVVOMiE528Wzx0ev0NN5dkcG7f/MusNs+9L86v
hf61nJcO6Y8tAUnNS/D741q4pYPL0phNVX+/ZG2SzLUw8wcAEiD6hBrDDQwl09netIza8ASJa1oE
NVa8v6U2K41eZi+XX+KhFf6i/8mrOA4Da+TGwjIVkhqRZaQ6mdi0+ZftGR2as+mDMelE2Eme3YBu
qKMNAcMmpTH8Gybvt73cFJCGY9ni2K7JGkd387jUfUykSjWDIe6JhY5mj4Nz6eiZet0ayO30phSJ
dsCav0pbbT+B1leZZPZHoOVr1qYBqT9iwjcrDuqUVM883pIYC3I7lXlk9JVHxQ6H9AjT3y7cgsxt
0Bzz1d87b1bDvBR3B+XQbluo+vvNgi6nhVx12dNE1+GXKaHUFAIQPIKLzS6/WBzAj/VctYwZ8cie
Kzebr+mZJE0c4uChMtiBOQsEo6N0QFynjXDuSOEA9k6kk+mzxZWYW2DGWGzqYAMFdrGXyqEFUv0v
tRQPDv+gLNI5ldwemUzecMmJAXdglxaNnZpoi/jiE26EH8K5zdVatskKaodzSFZBJ3FKP/ZM0xe5
9ZX+gIniid8klElrgTGjhrLa5hFp7X4nCF5gqyOVcXiod+bMWC5NQ9buVzPV33qrKs3/EXFt7c1Q
33kfj8JDJAjS2ftmvEH4Bw9weZLqqay/xGkb0D+7LIKN2M2Nqs1Zd3rnrgNeVaFC/JCu4HmXV4At
cIn043exN2Ziry4lYEZnB8ZIkdyMM99eDpxUyCSOOTBq0DmDXgbnNcVbii9RYnGhghGXp452jyEp
bAoaPb7bSpy+v1tw3yzTzKU5j7hau43ZhY6LNaHIDw0XlpLyyBDucJlnX3oUSAFEbgUWRzG+8Gfl
YtZ028aK525OCA+6a/lY8U+vMBVPZ/iPaCNL7V9rtSdSJMrFlBVx1/IONZHksOKTv1Y6A7FHcziG
hlTIrQ+PszSI174MuXWWd+XjQXtqBIYxxSS+s4xaf+z7AFKoeulIur4dNislguYrsTqm7Tm6GTOC
CwXeAnKJopMWaGPI+IrRL3jWHXIpQU+3M6uGiZD3nMSJXDe1ffbumkyDFwA5oMkkC22hnXvGes3Y
WL+3nhmLOMj399gyuUF+OLJxNl7LLgN3OYB7lMPj2HmMMh/BWFFnoZL8Qj4OCWy0ZNiw5ehtFYqK
bZpk+Kx+lVthwwomwhhtVuKRd504ClRYqVTmIP69Xo7TqHLqCaQakFJr48R+PVtHcEoZFsZkdgP9
xqUk7e9CaErnjxEY23Km6QOsF8mu9KUYFDaddF0k0UTqntqRam0LrqEkDGrpm79yQpQeW45N2RAh
2sbk8Q0no5A04Ea90KuRb66dzovXODooqGyRjvLMuCio/JVTBHsuSccrsZusuyXYjxALheg3UwEq
4qAUDfz6f/W8Iqdd9YasfS2Viu51MPpL4ioa2/Gd/wZ63HqMvEU5SC+K4sNcaSdpMdTt6oW8D5pY
2IWyqVsqImVeOt8IBJRlmb8HSfKzm5aMnPFUGNQVwNoaQo3w6JA6TI5DjXfqwbbGCGsGqvvEG/1e
CevWUyCBzNukm4Uii2i26iUL+19sMGHMjBUqda9YclcsjQxwTvdVuLzXBFQGvAzNPvaxFSRQoG0t
eluwkcPrD7uVnZmMA3xUwMU1wUdE8HS3z1k0DLY4TC1h+iJToCbmQyrIW0+MXE7GZrOBtVX1luBW
ggKc85ne0d8R3hUkzADPlE8LfXodMr735k1SujVGOvE8UQHG7dP5zp6NE0XjpwnTIhbbAl8y1zpv
3kZ/UNlQanox3uDfHdSS56dod9Ppc764z2G3fjNMJRLd1i4GlO1J13SUZwA7NO7DaxqSCCFtpQ+Z
dHcsBDH5RlRjvs6vNkBFtfc7MisMkYymHqKnfySxYBpCoh6bNUqSPBWDe2NVP95sY0+7YfvbrbMy
2eCX7pNEziV50ecJvt12rM4YBRDB5WN7012wB+qCkPIP25pF3tW7Tu9jiOqvreCDH0mCeJqavaVf
Nt1KVjAxcg+g+ATy15/j5uZ+NsWELMXgVUc++cQYMxeYR7kkshjeELNTBDCVLzClUoq2LojAWiKk
/kj4hnB4f+x5dVCkeBXRglbXBswTXwoG8/SCE93ZEMYRW5YZCyHcKlhm0Ul6pyMJrpc02tOGUNA8
GeJvD6zukp/YUY3DvEuu1mMa33hHqzklUx7puUqDTfiEQJ7qbJ50KJy/E/0F2K4LBawtupVskWJZ
wcQzSOuPimqpf7crdn8quFvPw/KrTGPwWUB2nDczwjHg7zYB7TPPyT4utSWr9SYlCTBz+EkAG1LU
/nqQBvimCV4L/I+luEgNmTzv0a9rf3QKJl/WEqGlSEb1CgyLtrgMraAxGibzsUJSoETRaUnz+J38
xJnFHSGE3kVwKZ2aFBCb9144pLCPTgDHTGuMPzGMlDg7DTrvGlPvnLb6SdcItI/ja109bZfez3S+
8qOSMIpsBJfbc0zyqimHhrNXkG0mB5GVPCo16ZezI0UTFcvgSKRmMyFwP3HEp26lT6a2H+o744HC
su0yvRCk541rKrnQ6oVzfghAK7yb8jyaSdCgoatmvUK59KiJZpyJndfB3u62AARolzYAWiQuGIAf
GBs5NVvJJ0H7bO0zgVg0CbMBmXSSvoob7Nv/aCTCPSMm2bjNOdu2peTe0fhL1jeYTctQVWRJ7PJ2
z8iMiX/L4fpPj0Hipw3d8MkX4NAwzrnSVUd1pwdC/zc9yZuPoWbtJrX+Heq24T93jO0ED229DgQV
cKWy+htMDF5D3/Sn35tNXG+wROq6RWcdRfaDJB1mBJpqotEEWhCvFZMkV0MHpI9G5StkIX5AVihS
L4s5DSr5n4l17BjoSeOKSW6K9sOz8ccAmbJRLCb5GDV0Js5L14Cwi4to5yVsBgBAAvgYN0mgM5yt
Bx1tMu4K8j2cJom0JvrRI5S4a3j4q6B7RXn16uu/z8ktnpOUZJ3yD4onfSxjDhx/BXxXOWWoAFyJ
nH0ZKVvv6bJtDiu3NXSpsucdDgMUUJVVbsmzHceOA9CLMc0V9kAmWsi3Cf6QNIYMJkLB7l+xCLOs
Cjnum3IrlBhsTwDVvLHpdi/dnGTDpZJEgsZGR0ZRxsD8c/Fb6u9yhyygqNXO4bxIWYYu8gEmmkfF
4n40I2ajOca4x7rMwWK8KwdV+JoYRA+uNB/lkodVYxxOriwsFPgoOqy+bkiMWG/eHbmLqZexpXU5
TJAX+wzToQHnpIySIKO1krpQ/71sCgrLB4J2FaFNpZy9RK6WfKVEzpX0aewRFpJ2iD9v20TWKa3v
40OefliV9PBHCQsHTiEYnBmIPLpmVooFZqLLem4R69vKbcqdtOECGP5fW9EYTywDI+wdzfZIaIhy
ilW9fPE7mNyU1ZwX9iJ5Qgp1KxP9Fw3J9d2qVhVyhGA+Ppwu1cOynxDTBa/j7icykHe4VJ4Jn3Qh
oz0wVnaHlHlIL5qpr17fjBMVveXgrPbzoQ6NNVM9x8FdzX9BkzNCVAt4NHQM1545zQhSrpkFUiTC
m5ZjhXX/tHDqnS8YxJRkvJrXGaKEdOGwsQwsy+P89liZMjwT1kXvUcHBRZZf70d/BVJpu5sx9X64
HaahuICBfCdd7xaXkk6WrAM5eoDlxKtchm35NTx1I3r2ZdOnwsr8sKpGip8CytScwBvrcyuKj1at
FSvTNpYe+O8qpV7302VXM1/qTksIGEdHKi1qq/qRxOU0WBQpDF2PlPmCc6HAZB8iZeid6B5QRhiB
nk8SK/jwJJ3vU7QSLwE3EYXFW7G1tmoMkya0PQCGgVimMvlDnphk5bAo1xmJHhY8GRnzBClrHFms
IPP+dCuBeEzmPWZc7z9f9ZSle/4s2vs51et0DgOxhZzsIexscCaeM2twvEtIl86WzzjCwvSXpE/2
/4h2z27ZKaZhrRFvfwfj1CKZNa1LH5WcuVg0/ivE6deIosyK5nPSmFvQqaHaSG0s7Lyaavohdk4z
qcpmi1Ouhm/dQGtQbzZ6VGro+IKjvaDdxTEB2GrWoGYmERJIQFb1zCb73J0m48klnPQ/80s3moKR
zjPduFfpYegZr42D606kiYiElkeGQW5ybuuEdXalvK45HBw5I1hLC6MrgcLGGGXokgoFNzgyjHeu
dAiMJNlnN9epWLY+srkydg5+tCEci24HaBrMfT01DScgmzyZEoQU4U/qO4Plt5oH8CNFVLuBBk3o
S/wYR6J75MdDrntzl1E4vs+asaGo3bo4c6OCLpoOnfh1EI8OtyCWyoVeIYqiTCjqV/zy+fNeWMS6
76WTlnOkhwTKre/oYwH+yEqjqszPgvhJMtdS4h6N1rgtezjcruix0gf/agntALwNpPNPg/OMpJtC
nu5sG64oCta50Fz9WcJt6CZOuz6xiJbGjNMaxNVvWwEwSaE/oDDbotDcovb5ulE+Y7bEU+kZ+HNZ
CayurnkMDGTRjIPC0kW6EbUKLHV6CyCzgk6PElvbfgf2UF+AgofWxCL+SM1SROxBu4dYMnycYTSb
pO4Rp9VUqQEITKY59B+ZABOv+EhES7lvVNeGumukKZnSDM6XLqySbGQ/0l//k1mJEiu2c4ppY14v
RVSK3EF0caCM6E5/1lit/rw29oaVmx1FQy3e3aZCRmf2H7ygreery1M7PP+lswvJ9F0/bHQmJBG2
tOSSby04J3TyZfSiiXe8bCB7JL22V5/fjQHtv55o+5SctbgRc5J7JvAm7H4G+tuna3JxNR4tWANL
1qdyYc4w+WrlJsD3m/6qONq7FzpGEY3JuvJCFnPZf/aWmpiky7p8GV4KsQPMafSUpfSPluz1PRhN
nKkxaEaOAhxark01uSmzqg+8S2MHgFlhOtdqT8ackjK7M/f+MD0t8D10496mLhFEzvq9IOPgKEoj
3Sv7wknZGFdKX32Q5Xki/qLLVv/ND1sBh1baCRPjARqd2sSoSP/uWvD0dP2dB6sSvUtB/obk3dKu
q/3YH3oZlxYv5fCR5EmjlBKbTyWC1YSQ+p0Vj3AaMRRkhHp03NwRV0QlM6T/J1Sn4nzfS669KCSJ
Fv52mn3j/cSDEixdc+WCE2fx3TOYF0oCvCDXeLGkpc/7Rv67Vs07HC/DDnj2wjRipWgwb+d7Ii5V
QnNxunL+TZFkqWGWa+d3IllFHYgZdgrf+fwssNY9jIMMeKsE4pu99amGpQ+0uIeWqVU3fyHGUQ1A
+5a6pmxekeg/PWcP7ZL8iRyvkX50PxLjYrS0vYObNniLH+K811EyEnucglgy4IdvAOdM4trCE76J
LooKvrReMI72RudNXI81II/8DH0AgoTlRgiz5KVl7uaPY3vTqtuV0ej8B9WfeXwQA/OnRdPV2VWo
mtpVD7yrlgC6naPasniEK9LKQ1mrKdczX6n2dvkLY1YwWfk4Qbp6F47DwP0MYlfT8QuT0+tVgGQ2
DIoaL8p8iwkJY1/SYNZz/uWiXLQllloMF5dyDKrysxZ+PUv6R2J1f9RwzmFp5raAvPFEM/znt+5d
isSC1x7JlnyO/ahwyY0vaegxHj8aU2NvwZBEFfQl7xfPiNc0XCya+2asHj+e6/Sn2i81uZq52oI+
krD/FNn/x6UNWdwxo9xjQRfu/pyTTwa0w5b4cVE6QbOYMdgI+9r8w7+a/GuSRQvkR2uarUWfMQDS
n3lR8mYCS66i573cptS4wnRAXFkHl6aMo5BuJaVY2fEzOduiEzOgpWvT9iJndrLKrp9fAxI3Izfo
v49bSAEvmLlnRuLRxDGZO3Py7ovRVL39pvrMbaTNquO9awblQ86uaMzoFyxf3CXBDgct9+YSIruE
BbtuaOKgLoS8rnMjsPatgoE9jonxe7awP6PNnFo5yvGVHggR9eDVZvKRyC4SET6a6NoNjWdOljB1
oK0fxt6ofrW0+U6ppZkuVttveo4RxMTnIEfIdaHGLh+znCvQEgmHhkQkrKFUHGHU5m0TS1FTZQSv
LAQRJoI0AECB21/w/4aWL1Q/mQ3UQS63dPFt/qj/s4m3+r9qLbgkGu+Csd1VyRcjgCuEC/SqbRbA
DCs6Bhv9YmqXgcuPtLWX4Oj/P9tXBuE1CxFG+S5hb2xoTgIe4wMV4CaUJtX+fBeIgwgxqQ1jYJm7
5vrfimyxMEg3PJ8XiloKPxacb6aMS00hJ6E9bvTnvHAG7mFUisLiedhJGoXpebRG50Zv9DV30Q1y
pAnm5N7KUSsWXfcVtFE8Wd0qL/tA/Fj40Q4rINjRkQgA54UX3RjfjxsVoFFRfQaAjGjgYX8Crx9N
lzxpamG5NiCotO1WzjR1q6v55HagyUn9IhhL8ZJYARel2kJoCixwq1gyt2qMoKw1tlw6s8pNVl6G
iQuInDNHWkJmfqqYlHRG01j0m+F2R/o7jnVhGVka3cbLzxiT1GUtSDi0HqIbvrrs8z9jNGamYasL
b7AYBAx1P1FES4eOY7AEPP2bE9Ym3MUij0uaTnwryo9F38zPhbThiBaxJ4NDiGVHWDzFEdNcBimC
75lNCFP3VRuN8LrTct3zQa4OFqlPrV6rmgAUGwwx5tAq6+vTwID6Uf/GC9Os2kYaGWk0un2mhSOj
m3Hd+fzJ9L3IaMrGcoMDMK6vqRfom4lkfOGaVf/HGI1zwquUA8LMi0jV18L9rKqsYPZJBW1bgQ7Z
HHzqAwEjrBKtP8qXMGxneFteXJl4WNFL2Hnvc6DtOxs6VzhAvajx8PDegljPUWzdQZO8z5sLuYVd
pLjXBzMCGP5yAJeu6UQZUIWWwGXHwZA2vD+OELM8t1TvLoFKSGHUj6zTV/3nf//2NEjWMo/2Trsw
Yy4UwNeybdKXpYIOPu/ktojVfp5HlkHDsK7BXpFDaQZ8U7GER1hImSyQvkSXF9gb707umaBSdFn+
IiM42qxwQodTOYfRhmInkp1y8FT65dG8hMatQcHXs9RyoYB90aqg25HP2kHSzbY5DQCZMlQcRAL4
fshXQ6RYdRm0dF5o4oitIQz2iRVusoXotkaSL/FtN41qyLEBlux9mvxlrqiZ/68PZMEusVmPazDe
rfIz8VaDcWpY41t00Qy8yEY15imazrIT4rcfxbyMkbF/34KT5pAoU1ZyK9zQ8GOd1U6dmrkfg9mG
JyYJi2RANxTCzP70471MF3R6dpr2bmMHe6YHoXyBDndKRU7ZMgW9Ff316GFNddPRWYsvAx2ynKBR
LOlZJgFdDk3ueagHgj/f/I6A4z9vLuCZ2b5f2ANcYbD3pFLp7HM6hHRTKxGlEz8bxfIfyY5RW87y
qZA+rKbCRTgNMVyXk4sbz7nKl42NBiYhZsQFkN1oPf+YuPOo5kf+tKMtr4gTAHYbzF1KlV9jxuO9
NVzPH9kpyfQ/bzuK/cR22BQFqqmHANdUQnu/fPDuP+tNdDv+GOBWvHGSwGCA41XkLM9djSXjO4iW
U3AJRmOBLVJWRrNJkr8JFpf5PZfFZuujAR2BbwlK9GBgiU4FNI9arAs6xaocWvNqjb9/blIu97uH
fU3BHUtyOuILC3Skbnflh73+H/gmww/GVvdULaTaWYxT5aZ0qCYx0kcfGPfzhnNBj7YDoJ00V/Za
BrLQVpLoVLCZTNOC1cdi1b2PMix7+NT0XmNkoSkFq5KBXVHq2TREkM+voCTUEYamYUAJdoPFMoQ6
6Qt1o0NT4Bw+W1YSQoo4BOQ3ejr7HOPMuUPUqdxcqvZzRs7fznQa61+g1wIaXckfGGbuQPK6C3ei
Y1JJVl3wgHEQD0koR7xABboi3MxtcvsQzw9DLNQ92x/t/6T3Iw3sl8jJispSNYT4Lh0V3QCS3pPv
5cfPkcNiEsK42zceyE/kaZWqwNG/vq0eP9pdtKbxR0fJrcbiC6MPKRbchp/0MoF3yvFMYf4BZ65b
tytw5aCE18t9lZmXHQcGBR5LnJCHljCFVuUDBQqxuEHAHzH+5Fd55aX+dNFfjbdCvJJtuZ8BpSlk
69aoNK7m1O02ZVuS86jSh8MKj+Y6JVTU7hWLVfVAfLBiZaIYbl+MrYQ/X5C4kaNekSM3nHa+UmIY
JeS4rrgXow5x7X9/UrQq/A/NZGfdMsgLyKCPa0PmkZJ57ETCYRuZkZfu0M0cw72QZ0spFgCZ3iF2
yDXKNg3bGfc7Sr7LzyLuGBH8z7npGdV63EqmdBqGr0q7bGPJyDjXnMb7uWBq7TR0iYzZfHcpNS6w
VZGGrLErf9xGbHb1oIfMHg72qzNMWLLdtzoeW4mq45v7DLjt239zk/U9jz6/O/973gb0EHAgD/C1
fMAqJc1vIsSbmOEIsddwRj9CvoNSkCAY75WcKI1r1/hco0IsLlw1pBeTfPFd6ibb+kozW6+IZ+Rv
INlJxAtWyQL2Ij0q91VaUceSSYi0Pot8GNwlJI0sBKz3lNUMr2b+IUo12jRwN0fa/Vzy8VTFeu5l
8kKxbgxgGNQ6iDjb/6vslMYSzePmGJDh9TZvNkWWtVkRM2HoCx57VjGEjFrItDrh6Z2CtIo5HgXI
Vw2zjyoSopk63y2KxBvqgKDhW7+gun8H5R38si/Yl36CAp6aqHUOrA+TNOC8irTG7EqyAPFy38PU
fqlnRTG9NHssAVGKTL1n+2BFSYJ7zahRuVZQswZZ0ZUfwl3YoHgXbrdlEBzJBZw1hIc9xF4+QUi3
AS+yeMT+Mru1CMDzAWl0MasLNet311AndFRgTEvtsCMeMwfPwUIuENd2LKBz1JqWxPM0Lcgcz0tI
clAAAt9pDoihphpKv2BOaTh8XbJh+gJdOm7GcsqOZXaeWMMbYpi0DVxFLb0gXXXHIkOQSYz+1D9a
POcQPqD+uZ03rfkVPf5ES3lkipwMyOGmmh3glmsgfy+ZFoCWW7r9KBuFVACkeYUqPrm4GwSC9Rpx
XKkbdAayAH3wgLXAzOyGKQygYEwqev6tIiMR0NExpl+Ype53bUWvzdvt6LpaJJlzR2Q1irfNynhZ
iC5oQwsxWUZYjzjJIASusVEXyx3eBvGcYsfe9x+vMGKGw613CrHJzj2Ev67s9DQSPsXKodTYE7b1
MyJfBzGL/Y+4Gh6d+7KLFTNnRK3uaPCSKYPajah0ANsjZs6LyaFf1PUPd1EVcCbcyoEP3JWq4AlC
/dLyP9/MDcmD9NMifpdWCaxPzqZ5BHWnFBXvc54VJ4oGUDVd023fHdVnQVnQzOtCwQjr3jVUuRXI
aNuu5P2jgI8Ck653CrAa0ErmfzGO3vcy/qeNKtOyLeomSJdL0Gg8l72Hth/EPEZbytt6Aq41knq8
09m6tL1U1e1xUta6X8RzHaBLjLIBfAQWMkkZmCCwVzS0yoyZ14JEZCe4euIs7xSCjRWzOnFaHA/k
q3Nfm1T9dHWChq3CBA+WvedYtbRfs6eIRkJxOQQSMwHrS/e2jzT37uuFCEdx3LeIxJ9MXbEvsWXr
KBHX6853KVBItvd3NtmlnMkOz9v0OMbe7fD4S3jl2ZCJJuquAKTdu4IqoG5zdx1HHIVkvU3RoZq/
BbvpFqCDDdjh+iA19WNcbDwNmcEvMK3F/pQCuv4w+aohk5u5tBFILtL8noVsT8dmzO/fryg42q/3
+ihTM9lEGGzCJgpkO7tC1LKxzTC/Hy4fJEoJ5l8z1I3UkOfLw8wyiYHBDSx4K9GvGr153n2c1O/u
YXRh+zXXCMo78yH7ZcwWrs1itGoFd6E+YcwCv5wa+YPWmByi0UJMiMO+VxFfcKXvkVz9/ZoDCqGr
FrffSERx8ZGZ6LiB/b4aEK408MhRWQMBO7j2yb5SGRzZNv91oXmsBg8HJ3rFPKdd1afKTFsDG3yT
K7LhLsh7IwUZ0hAw/O0C0Y8QdrDZTkLzkCzc2FY+lb6rrdm+w48/fsf5b0dM43plpqzxb+PFaphH
W47ijfOaJNo0tm/eXOODmKKqsoe+Aty6KkKPU89M8jbztT+Lx/B5gnRYG1dqxrbEX2j/zUnVCfYq
o3V7jXBU1S/JyczWsxDqoaTRPDEoItD7UORwjPRz8fqCwjCb969mbR5MHpiRpzkgAQT0VpJ3Rxmq
dhENWRJQFQ/gwaUWAeAaHYVirfMj87Ji0VA7ZCInxgmqTO58OWyrC7AAt4T9yEZrxjIlvvg06X+B
PwhwbRT59i7RXFwAv3HhHzASDXortD+Sf2fIvZfLcx61ZFv6V1qEJqG+dxxuDYSOgbdO3XFgwrbE
mMW8r4crfvH6U9eEhHhYZdA+9+pPMSppw6pDmQ0a5FUf6fPnGFLkXIEoTvRagP9/sMAJ8okb8gKT
NWBI82KgilNz8cEGpmCXbpQoUugS8JlxxYeCL9fIdW0qPJNDG6pJf0c4BlEbjLWw9CwOA8Zx+7WY
BythJfD5jzMxV3hMz6bfCoOzTvoKH7dcx1PWpKxbC3jsVDb7YpkSY9xgywqTvmLAAntZjc7ARI8w
Tq0eLae6NFfmm/eTi+JZJ6xOG9wfBnY8b28HZQwVUY6djEkJbCEKEgn6vm+t+rx1IOMnrE+Uin1L
HrKBctiLCZUQ1o4fwaWL8qLzicfdGy5jBk4xm+7fxSOfg4A1l+jCxmmAc48AN+dIPZFfhmTWAoI9
enuJ+mgWaouK5dhaRf6PEa2EF4piuqRXlD9nAXcpasi7CCcu5yXUuWhJgDOVnKbSyzqFjAyLZXCP
CvhpYovaCO+3U3AT8s9cxNt3PRsOkGICu3Y36f4bLnBostmkZHksUVWch/d5ydyX/g4PWxDpIpGo
jqSEhWAUbSdJV0zDxKxHsjnK6nO/iSEah4IQyg6vR518q5NLXK6ovOyHrfvAbDn18TSSvBaXa/1U
NlnXjsgcgVdtTaRI5ubIzPKhAZNNHzpPVBh3eIgvhfa+/KW7wOQgKBuhYSqGhVJp63lofDVlxTx5
iZWAucYI1uhu0cLoCD+o2MgdzE4SAHaEvmXyg03/ceDnfop7x3c79P2PL3wo2XZspVqH9mLKfwVA
ardc48zqj+buorFgbmetGfTj+0OVnwak2tNqMdsHaNOIFxe9b3F8wQ8SnAGi29RdJwZ6EEHwnY0d
us43U6aYbA+52ibvKGIaCYqyKd3S6jom5ho6Ly/e0sPHs8rIv9bluLZOQhWqo3uGg+x2zKI8f/Sk
iO9blV+MPVg1+k3dTZsGnDaSzMTaxoQG7OT6abIA7msTABPJWNax5vZ0FDgrNvd3GZanhxp4Omnp
IMmUrure3Un2RkuxFFrXyN4wmcnhZNea7n6G52HYKT5mR/14+4LtZpP06Bm4AY7z009ctTQ064NQ
7BITfNrALC8ARiBBdFAM/q7vrIoPmNsezQZQwhMylTRI1Mrj4/gI1uIcMypxzmxbvp2bgxZP7if5
tman0pHmIyy2fxgw3S6+NrAqvaEH+t6CWV+nfxtzgm1c5qemRZBybHG6pIRern73jTv2xgdXUwcq
DUVwyU0p1a9PkAk/I2GTE8KOijHYAFPlmKRxEj3uPcNRYxVIygFV76vrjIrH5ud5V6WSruUXgy1b
RPAGLD0KYJWg0Xic5By1YXfD5ABL5+Wp440rOY+3vLh3+Bl8bs09n23McbyCgL8Gvt7zmKZf9yXr
MqMEwijRD97dDqrJ6IH6sZl5fBK24CToBDZA6Ycv6HeAqKHbujyn0DdHMup4wkGpLq7/wkdQYuia
wT7Ei9Kf6bk0SIbpwMuR3QQa/qzwDhvmwNHPtKaC1n2eIi15tVaImmp+n/4C8qOM+fnNxefCebkI
n30oC301efvEktesCizLloFqJbJoSQrqofxf9zwPa8YDMI5gOk/DM1djcodPrU1Thy4UKGRBOYg7
tMbU5I7DkeauXATZ90twA6oyABx3KrvcOb+GV9P0+rIgKc/r+JD7T/5+uPmk45ITk0wMc5OQTqG1
35wf+3WSHtRHPKMDgFWdSt5ue0greXmcd2Wr4i4dnHzw1lmsoOx2MK6aFrZ0QHbfJCXIHrhNXwmN
7KZYrAN80Fu3U/C4eGs0Lx3zncn/JgLYPbY4XUfKUQEj0IL5fHIHquWSFtdpe/Y1Bk4RJwfm6cBx
4OvJg0N9eI8A5z1+dJiFu1I3kYNtzzhnnZzczvCBOobwYWJ+2Z607uymbmqDAevNWT95Cwy88h+8
uO1vK/lPrU9wKFV+ckU1WFiXDAPMnLrJ40NUHX4kZ8M6veQqbBwI0UzdynVIbynw3HCfUHfPvTit
Z5+/9hIusQ3AEjgdd8a4+w6bt/qCCoJdTKyJK8Q6yQ9pWXidoNYxqzMQ9t6D7DRij5Ti+6Hrv4Ne
GkQRjX2RFCsK8XTB5RI7xcoyP8umT53vUahLO5Gakdz5/jMh/dNHO2rG2i/8MU3G/CoHfUeuOz1s
7Kt7Ae/L8RkJYPTbi1/jFeqCq5KkuodxKTjrdeCIvmr2ulg0cRZk4u4Kkd/ETPHWosEWocxMhGRL
K0d5JOdak5VwaMZwGQ6jarMJT6+BC5G4CL0dTAX6aSrQQ4jMN/WrYPUBcuKmgc2zdONnGVXqHhMc
1OVqjXQ7/ec7w6YgS9eNfeCiJctpXwK0mrWRcDZUZictWkeq4jT5VLGE8N8aKa2qfHm60jBau1AC
bKid88vHYkCK1RIcnvc8tYHEKDHgfpWQpj+Pkbzs82qdYDF0kG5+yeFP0ONNFR92I2GvE3tPbXd9
E2FXsr3EfMoxWX4yTu4Lt0gHXHrqTOHNhgpoWBb+IXnuMvWyiLBGCtWQy5M9JmUoiW6juJmd8poc
Y6pr7fY5Buel6MUNyYWDirsdTnGiAfTfUCC3UBduVWTSe9cSDqXQF21mWuRWtwb1XGoq9otIxIFb
XIwOW6xQGN+ijgo2KIO7/NevKgwJYAxWeatQ+7JaGDRkwt/G5yc7zeDAw3+tYsDNTaejw9kyy9X7
EtDNg22VZfQ29hhEais5TnaSIxO6xkIYMdyPKbGYhAqC1jYSb3qKtv1aNVvOc/iERZ7jK/79ZTqy
BlEtmi9MDjVex9FEpdQPEw5O/VxtZ2XXaogEstL5ynuY3g8aLc4+QBlFi+cTDU8bv54Do2uQP52c
ZXGVslQv0xNMs+xGl6GelAJkCmbyr1NS2uUgoIvff1Mnoy1W+snQ7t2W6CVwJvPKhOEFp0TlFtwr
ufE2AvW+/YCMcaR6DKP13FpFtlqITFlokkyLft8jVhYIZkin50HYg0gBDMhWapNvydEPyVdi3E4j
cH+uGFleE0ahF2UN5OBFlmjS5seQU0sz0emMC1oe5n5vK3rDvpYDPdY7RXBdQG7Ss8tmoJ35gWQ1
GHXeitVuP12f6UkaphbBc/WhraZHl9mAlA==
`protect end_protected
