`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
fPgVN3gcwqWmADiO41P0g+Trmtbr2K4yERO9ZqcongU1ib+RTBv8xFDsK3ZjRk3zvwO3QcclDPvf
R86eFNguE8XAjVLmVW4f9TnCVCf3SNBKQ2GrwOytQMuc3kxnnI2qemMsHHywJTxmZVGqqmlcfqNH
lPsMlhWOeMoK45wLsBvQKuUn3Ho9EsRCqUKz1iENSHOmXoBukG5NEx3TG5lq0sao8JdyjIAb3loR
Jxr80M+ttlc0t8QmydJ+2ZwGdjDc0eTuGp6JpnN8ID/OhHOKI+AoQRKqk/mOBIbvKUCdaURvjOZr
/7T4lHY391/3PpFSj6jifem6hNd7a2j+9o3wJA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="5srwG1qf7UKlxAPQJxOyUw1xVrTRhWQ8XZNb84h7fMY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`protect data_block
TGolr1uCeN1KJhISmFhSczR77SfZE3RZxmKve4IDTBlPoLlanY+xXoe87CELc1O4TmSL8DpAM9dl
q6567wysz0SBHBcJWf8W6NBwkj3SmvRsSAsYccJftR0j5wmx6vInHrMYYuOgNGRuXFSg5XkgeiCn
PC4Iwgu6hfIULaI9qNJ+zWSq0slIFkqCo9459Ml5daDfRsXSD1K2jcKvHhy78sx7qyhnBOZUPtf5
cX+NbtC4BnR8ixd7MeKp/uj2F2xGSEHRwk9XyNfj0xZ0Pq70tdBUwyh8PEr5UZLlMTD9QONZFMCP
s/xlioE6hriQatOXcRTW9ikbnC5mlg5pKEGQeRBx3K3wEdkFu2zeccQvUcOnnbKR8VGKDtU17A6V
F7uF1XgTQiLgZWWfkrci9+iYWxVocmUTyTvWO4CIizt6I9C0rU5edO57HsFlWqv9y5jH99FQsxJk
d1BPHWhyEFzdbcXkMxLXoUEWUuXLM24MbTlKyAryv3+lntJ7Yvr7+LN+y+yNGIZjEg2Fn2qJ4QUd
zdC0JCmTI6fyRFHGgQ5bgUUhXapACg+ntJYQWDne2eG0iD7A4mW+4jAAMNx6ZP77XwmrYl/1r1VY
LhaTrOwlHDhllN0Y4fFpEnEKxIMFNtUNQCjYYO6n1jtUyAJFo4o4zHHdKtUGjhu5szIJ81JywjJy
9vSaO5AV25n4gUosSAbVNIMImo4FPXuo/It8L5EFa3EHTdsMQrFM7w8ANGxdLo4ahjeqO7V3QMsY
pYRF6ocM+Dp23Wii9OyjTtxIGQAK0UtKh2JrWKgspXI3HHav6M8RvKgMUozyiKDWFunVEyoWwGzu
uZsBU1/s3tgStwAf620OvkL6VsT9rvSJ2YZEIRPk7IbDtmH7lUVzOyALI+Hz37gt/odfo2rRQWZu
Y6oPeCYG1DS9Kc6OiGIo+UJfoeaujHPxfnH2OUklkodmQ3qvq7TeH2jwrH5A4JFPUfqHbSfDNzQl
ELt3wyzRzxCmk5iPg4JQZUi+0NusoSx6uEO/ThNy3GtwsmSCcIJVIXsM5ogefqFAwVcLxywF4zLp
5mU/AnaDUh3gzyJt8NQVZ4QujcYlAIgLY2/U114lys1vogAFrNnsIFGtPhdPUi3Lg8LoeW6PbFm9
c8ICb76brkqT1ky98Mf44+MJ1xcmT5x5cb6OceU2r3FNshINcouD7uDNzA4ZLxRgZ6OWve0cVTfa
kdKtsrGYbEJmgJsXqbVQQsWZf/oxQ9hfkvFS/2EewlulALlc+RxzLMUjJUxePAUpjj3bt2Y5CIMU
Yi982I2dJL0TW91bd7gA05IYx0gzfm1NYU5nRqMZaENH/2bL9KVa+eL+g0UoUUSyR0dAwMan0MQC
m7NwWzMa4FuT1mGdUYLIDD7JxHR4SiNXN6BJ/lyntKs2GpDtvEht5UMzRzw5YP0CW+mHJ8Bbl4os
f99O/8Py6TORLhWVapl/e0wECcU2/MwMOWXAXcjVSbHPnKlAyZmuFnt7WSzYFKqHF3cnOvrG1Zlh
Lg5V1RGbkoSD2jVgJ5awxqIdvM/Nh004L0EGc6Jb/bb++4lp6mzarUD2TqVCtAOludjLKSrxm2Rs
NXUcbI46b8jm+w3kTcVivukDOXNtV7LfIzAecpYg7DLM9I+B//1F/aEOexuBo8PlYDg/IY9MTSrj
prRrje/GJ9dqoZnUTpcAyEwEddT49PK4EZLIHaRfROWZijNRujl1fFGI9zK6qhHnaH+jflEnnfdh
KjMYG86eV/w5Y1T3DK2NYnLc3glXXw4YMusXb6F7199w5oMZCusTJSmgZDZ/12ge9tdRNnOM+gHf
nAzYLQCLwTjW4WXvnELFMPaK7PLP9nJxLbNApUP0VbDs+xuvA+9M3yXUR6FA50EacS6jDysvOCd9
j6nKwedp/oG3MyoTqWzG3Kljdw+3W6u2r/kMNm0EknrPAtpdC6QSnrX+2Q9Mt6GNIk2AuJQPfUeI
4/1DgoTugqBEsuSe1SZwm4+1BFgA9EqvARsp8kl9+q0cA/d1D4Ed9FsPTFuFopD+Md8LE3gc1AKM
mwzBmItVnzJi2zzVdI2v01SlkdTt0s/EKJiPifSEt5k422kRwrsAbZcKV0kUTGJ32mF8wfmMJOqu
YjdDS+1LwUb7+gSRXALVYj+JluTqNL44z8+Lze3x+aTmzPRqrK2kyuVj/+ggr34wFV4ap3RJzUH5
vYsRD2M+uulC6T2glMye0YgR1kfbANrNMHJXluyrJPXFA5EiQSkk6+HCIo3Ui0qJYNtWrmeMlRvR
JNQ9hDvy/58JZstj1LN6/bPR7XcysXJx4Hsy6VzNFmll5Bm3dtF9AWZZHV62VmeStjtr3LwZ/dlP
Jte6JmdojFYpraMqwWoMyBYUzeR1EcBhO87KyxEcFRuQ8S99F/c9ECUO8Ozlvf0wm0bdhB+9jfo6
CQrtuWs/u/G5f5qyru3tmSXxjSn44YMaMjWNx/DAv7uwGppdegkQxCF3Nt5I1kFZFVFX+is54vOV
XJojyHDPbAn3ppBahBVBmyp7apUJbw4Bx9cNghinevGDI025olGs5GRkkIWEuWfjjhTJWAO+zpbq
c+NDI0MhTOClMrXzcTQrjUpzCebOpQ3BuVTkGMywRdt9ayyrq2+yo8YHFfzDIprxLm2HfAurZV6v
dqtVAVpUKWXxRdE0PnmglrFrDzZ+M6HKNcgy6nH4Qhe2J1Zq7bOmj+DTfe2ym/PZnlZXY5BxMZvR
a1trX8zfjtrfPwAxedDzWcWtp/NKJGsAoZd9jl6I64nVvpLmC2ddc/ml1K3xuFd/jPWo4F5sBkBd
3KXjfRFL5lPyjaj5pqMogpyM3xdTIkCZLqviK1VAiBlHChnyeoG2Kwnmy6II54PINAVIq7nBiUBN
zLSei1i5uZX29QWQtfgIp0d1qe8mpBzChtW1S6ciyodstbOIJgT0hVux4zO17/63GqTe/oeumaL6
fLDgWZsZ36HmS6eP1ZCAkxBH+Tvimo/YmG6Z9GgU6k6J/+CkeUQ+bOQRpzSiy34NwScINhneEaxS
Y9S/pqT8o4BwxMS9iHcKe6eVW7PsPMyzuMSESWtGKo+GyJtavUOFfgfHjSdj7x99oweojCcyc0Y6
iRt5GWBpsYPhq5m9Wde26vi3DqPzPtuiiqBAKzHmD2LreDRkBHaNkyHZucDjXxO1w+UPXCbypgVP
Ia8ovZjPt9nsrl4SHYRlbAkT4zhC/UrhVInL/2ynu15/JCI3JfDM0aHpudYDpBpUEiNDWx7m8ChJ
OZBMDcisB14vpnH/zEufvS9vbPNdVuV8xO5jZ4mpXUOwz15tZry9Yfq0hWF6BOgIx1fTOyPPU6QV
cudrJEF5Xz6HHqOKel+TOYo1ICoPXpxa/mEtEps5zkfinkPhjGGo5WzTbHZnGNrHgqFksWp6h/mQ
QyuWvH8oDzxs5R6jhQLWQ361z9yLmfiRc8hDWn/L3hOlFB9yWzan0bz/007CVso+8svEmEWQqE6r
UIu0xdI+H4vpkF8QUBAmJn0n+5x5nE0b/9ZAy5XrfxkOddpIVur1uP5dmWVZ/YCXdudrI9Cj07U0
hqrG966T3twdgIc/CSqKBSKWg9lK44i7mbPCDIiVGQ0NFrdjeM5CeFA1obDvNNguLR8mtldCK0cc
f3lnPMF7NC0vIKdoHERW7QB/QWkmpV/Rzl4Y5rjwPTfGe0/KuK2Kg8rr+1TgKlyBusDEa/w4qfO0
nxofIxy2KJSheO3D9wC9NBLK0nUsMoalqpPVGAkI07Au59qAP50IzIGAvfRyA3uc5gJDDMJkwTec
HJQooP/O7Wpffqj1VK+3QYt0UJxLLv3Q7V6g3L23Wr/YIwbYJMarNL4xbbVoKgvcywQORJUEj7uf
g3okb4Go7gx8POUuOXzoZexxka2COq/56OFdjf1SLm6rWSm/WwqDGnnE8Rtmd76tHeWPsvWvzWEo
PqNsz/wnZ5Z7GMIzK3yJ9yYPmiTvMzJPJCQWkzRR8Biu6DWOE0n9DTMk2kuybcFTEGkOsSuKYSaO
csII0Z7wdl0QOA1MEvhpqh2y2+WgdsV84mefJbbnPct/XKPXw+WrFE2c1YOSK+VQGTuo9at4DX/O
aZSZ6+8FtkG2VovRovdO5288+abJFkbgUKG9IkjVO20eeWYl9hSjmX/2vRLOAptEm06eZf69tG/F
8zKitefy5vz+mWF6bV1NOvhhYgLKcgxo6vmlIbe/xvhHWknZgeSNbLOX4DPCRbGFoK5TMjQZVGNs
xpgdQQUlaGzx4ihGI6ZQyFHIQdq/ArBuir+yUzuX9MbGyIvOcC+r8PRNlr2iLxonhOTvRHYZeaY3
PVJq5oemOg7u+eTesAESkl3EJTcLqgiXY2gOzBpizjvbMEY6vgvKRSaJOL/dk8jwEZe9z8jrbCPf
6kxgZs+Az9tywdkFn3uXUW8/o/m9C8vt0HflmTMMwIoJqnoIcp2lrGZCiJNvDu4+Pilb889G/0Fk
2ii2Nx2k2I57fQllfRAK4lah6aeGalewZUlgbjv0MqZvERpWsw3E4wBFOSNNJHLJnNdBo5/nKRPC
woV+RdoRTt3A/Rvm6LS/YvRaP8OjTnM4LdCuAafHsulcJMdZ+7oycbK+csvNUiMjDfUIQ/WkOibh
R9vjsyU6XA2Xrdr0VO04t5YZh6r9eGNHEfoj
`protect end_protected
