`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45824)
`protect data_block
agpykLWEGc826hfOyA/U/HjF/q3R9vh0KniVzkanOJsS5QKiRxz5SLkFzZ3JuRE9SzuTjqqTihrt
a2/1fGtSfKShxsfiBf+tgCocR9gi4rMx7bjpk3bu33cByZVdiMkBKr2fS+ksa2xc3E6Kdw0OXPQd
cmFBMfX45jjm1lbG8upiMrfGMmRIWlVj30PomDxBlpWJFDBRw9rcjFdFBkSKqHGM13zp+kPRVw9c
+3XiJlVmb5qCB+pyfajyaMB5rvdEFl9FnmrxpgPjB0kfEMi1ITGzqZr2YKbf0SO7JmtR1y/jbLpa
M+uoOeBVOMYO6xx+DAQ24R/sgotcP30kZTkJYEkUKff1ltwSn/xtUomaWFSRJnTOFBfeH6n78n8w
JlIvrIEmO4BGSo6vzDElpy42JY+/GS8/dj8kVnhXPeJids6wKogxeT0UQNiBOJk2cFfR8ir1j9fz
cSj2gfEXKr+me3gIbbUVwq0s8eFoz+znQ8SHYfonSivk6Bg324Yc7DX1v0miELFkn9rrcyJomb4F
VkopoyPhiX4JU46TAYNfXRl5FskzvY0TFpSS5/EFWKy0GPg+zKgfQvwfBhcBCocnxbdUXFW3ev8o
jw1bE+CgYiP1whVs8jz+qeHCLzn9vM+cnQuR2C3C3VIBCNmaua2jO3ano4z8xZN8S1Pxqvvgt9CC
Pw7Em+sPDGGCzApzhaZfl2BSSmhpse3cq7sEutlSFCKdHdTNavc9w4jb7jF+dAFbUwVpNcULSeVV
vfb7HaervjtEDKA8EOnI1+2/0iK2iFm2dAgjhVFjGq1xoJhaUD3ytE1TTGsZzsUVFjQcjgLlTWTr
Y8sJXKqrVAFptXXsh/OwY7huTqtGoKCl3nT/43fHxAc/AORn4frW83RMNZH4LKNaWRyu6IRYaCFj
c13RB72zj5DCr1xfNIWWxrIVFcrn1uzl69Sw/MbK/KAARTS+Nksw+c52gYMuE8Gpjs4hke+vvuvc
x6JaXKRqXUa5kyUEbjE6219Y3GQcd0IDGS3gbBRhdeiT3xoLHM2nTT01mdRnI6rArY6a4kVvkr2w
Spc90l1i8AHEvhupDQE+cyibstqOaFmxOW2VE8r+7KNSikBUtk7ckglaY++5iPzCybB6W3Xw4fPc
OT3mjWClJ/fzmvC+Ga9EHsV/F6Zzk00+Ttaj1Iq27t1RiUokFt4n9B+eeMXlHu48gbK4vUJh01qm
sf9rNK8digpiAiQMfMbzZ0DKOS2jafl7qbErGigsUBdghSBU8n9sxZVRDzqveI6B3YYZ14BfOHHU
dLPE3su4mY0hNkYBJei5+zt2dFU4VeE7FtNqxvwjzm90yN+GYRQpx/9a8PEco/w80yylLy3p8hxN
mKMpGjIrRGM4QYrpr7NZlfwBVfiTu0CtRfRc0LEM4OiRv/8oaK/EB0hQeoaIv5ElmZTHcFkuwAu9
NC8+Goa5DiADRJFxQsNmLO7CVB7CiyxMYP6nLorIyHuR63q+gn1XCSF3lvPnM0MynWRmMIR6SCzh
q+xuLfxPOIxkfrer1H62RVBSg7JF2SknrgqNZ4wCCCrZwQnoolSZyjPJad2PFIbX4J9etkZHt9rH
VDz+abdG417QwbjErPToVBqpjqL6XwRVOiWxS9H5wqE6SqMDaXnRKM18oQw7QCE1aBwBp64mkYGL
gc2GLkIo2dXbYj8GvyWfuny8mWOJzyD8ZtOIJVf94OJA5EkBfrFWLUTB/f1kLbr9KzL/zlsV287/
k7yJVrxLIbGC9Z2Nu7RTYZzja5tKDC4J5A5u0Qn/hooVlUGHNzyWOzFHc4sj4m8O85k/hKHmYr9t
wJtwjgO3IONArAJ2Zju2vpIGoBfAqEwhzOtbe7/yDigP+Vn/J739s4iy5cHYYX30Ol0ZL/abmaGC
Z3Ph5X25IIjzybywB8TZGvRR/oCVUN0oXumcM1TvHQnQqAanvsxIV8wenKMUIVK3siIXihY73xSX
5sCH6jfddcAT9tnxExo63BvsG3anY8FmRHfNcGpF4R/TCn0M49cm+pUfR5tZ0frnG3o6JMsdM/47
SejD5R8XP4EX/Svy06zjnwc7MuEx2iQDlQlY5MBHHHgpADF/ab4akZANizRMwm6LQUxNYwv8V/wZ
LPnFuRNAuPioutZpfikENiErTwFZ3cow2zdCpb/Vtv0aNV4LnOOjfoWqVd/+Y59gcylD/mxI3n64
lRRDh4/abfbb33MPf4OnI3tuAoKZJ6JxQWeGV1/xDHXoHv0bsrsbXA46/sqgZi8sHmmBZSr2u7cO
T7ieG1LBlUyRS6t1xPnTcUmBPoZAuSGaIbU3sqVpp2cpIvOpc/cAJ/6yArT6fI5AavDHrRIz07SK
WLpER2Vn1L9TcfikPMX2z3UiGazFwy9ib+foB04sNBhUKav4Q8b2ZQtHMzFlvB9x9o88l8+anQU0
NN4KsvdoU41r8NXW6KpU7Ascjx34BQhxxUWomc6OzrSsv8aKs8y3aFjwtOcG6GuJKPYX/WNDWhGn
DFbwlejHTRiwuBwWyJ0r/wEUh+IYrbRMlsjlBUYCs/9U2/I7eWkKe7zNPLF2BmEt2NsICD0wjAY/
JjUzo66OqGtg7XmLRfTFtbX1drcn7dWBjJrk6jNGyr6XjeEaPNbMHR5t1ZTmAhf6iRBcpij/fhNs
NxeS1qfFqMnC8VOsxwSEuyL9jVWsM45uq+SBykAcxghFSEP6sgDBg1e76DKNVVvbseYD5reRNVnn
V0DOn/WH0CfJTZdBWKTSE4C9oKZjAMOwqLMPPI73Pc5Exp3bqtuxIzmR4trS5zD5tBLr9WQCRCI7
/QRm93CqHEaQWOILxGlUhTHEGPhTOfr5NvBwPjP3qYS7YUn3G9bEGBIBkYn1ngXymiJIfDhxJbm6
ewUINcaIPZcjzCc+WP37dHAIW39HoLdGDC8oySFx1JYGywmTu9b9Uc4M4KYKAqfDvEcBtmi1WbWa
ACoEob07iKdPUaDz51TU5pxHZk7QXwQOuLp7SECnGrkNkfTUTIZNjCEITY40KBt7pLHDQKTDch/L
KamNkrvVuqiLt8uFqm7KPLqLfLldTnr1j4ega6ctjSZs5lA5PDVFgtpFarOBzXlZ9b27bHNinrLG
2JqQ3FfmuGy/ytwYdW3EHblScdaqH6sIMWaPmRg8K/AL46CyHLkuf06g8OyuS5slK96fTxslG1wL
2hl7FnA+Bu/R/+tr4qsgo9Z3fE6yzMaVX7ipFtAUYGVVxjN53fhRPppXCo4SqciaUBvv00238t6R
okNZFsFtbDwtn9sgHMqQnoz3b8oT80sPLLQoMmXvw72pelN+/IuUenLrpZtvwEyAgVPPTqafNAdz
URm4CFcZ5nrF+WdwWcrBR6pkJz3n5x8G14EIcZ7INCjRCylmi2OL38EF7juZYukiMbW0p5nG1S53
88avjjG0zQo/LLWk8Eaq1kYhyz0+9hScR9+iWEx+s+sepHRw7hUWxHLJ1wQ4sNfzRjK5IjBQeWuY
eAhZdpOBGcuhSy/dF2iv7ad8VTLUaXmydNAAzw0EBM822ySiLKCu2HTJFGqVbsZUqDG5MofqtN6E
KChCcFGUXb8WXTyAzeEdfaaRptqkUxVQkOWT4GmIScNqtN3GzU+8HbPZKHHW+lVeljcuPscXjBlJ
rf/eoTSZ3YRD2TtdYInF9GLFm9cC6hzqwge2w+WS1QS7E4tzbTfZI9d/bYYmuqBn/kFFyGbdtK5I
YxlNCGvM7yuOJ7cXErDX5xGQrUSB/g5Tsjmxatmki0tQdWiyh2uyaoh3WfSQRk6t6eFka4ZeTk6P
iiq2Z2rqRx8GXK53/Y/6rPf6OYqgoGHv+cUiJBSlPhTr0B5XED7gEgBV3volVDTqihAPJdazb5TA
G2I4ac+OqMBptBlCkwzWbC4vfuMPFpNUq5TKBVWHBPT/weI/nXqItVzPTNiQA4fIfRjJpX5uJChH
dAjqANpVZaky4wtMo3xBA/n0wEeWoAyvbUBohRo3NUOcYjA20WNIXgqCDxHktondKT2hb85/xg0c
8J+s0nTXII7yG2usu3mMMkztSekDKuSC6q1MPXAkaDW3QtAl2CO73F8OGY6DEmJLg+jJInCdRo9B
i9zjt1p8c+dhQSQJiZz9gSg9xpbNd0QIuab6+ckmfKjZp4ryL7vX/NLy+TsulEh8hYEMwsGDi4ej
NZLGuH9OH6qXJo7WmCmT22dMQ0ndr1wVLYjl9yKukoaenAJ/T5eUrHt8Dc8pYDZ4qoWjdpyOcR3O
0+iaB60h5fxMt0JtzV97mTQrAesUZEpWqkGsASCBcBbLce7rCzv5WN8ZJpuL0SMcsNcmGAwdKHMf
IRdujYBYR7Mdmz9YySeSzTgPOFPQ6cK3CGS0v5cbJJd/MOme155D7xfniJpcMwiY2GW1FK+b9X1l
/p4u0Ke0smYqgfv70nK1VnYJAq0M3g7Q4Np1WhxjkcfUEcTA4SI+aGAC/j6/plcgccNGrM3RYCL1
neB8w14oHJlOYwDWIJqXfQIJ/Csk/RVQLoTPnejtcaXb+uiDs657zWTSaKWsfoA8TpD6Uv9/RXqt
LQUHGJ0JG2DSJvyA3I8PXpfrpNtaLpdkhIb/GEgk7P4OMWnt6yQsSq6xH9u034KNvlywNwB/R3h/
334C5VgwO0f5SRqiGVFPiKEy+h4HnCQ1IHATkB25LYEtGrCuYHrjHA+SeD51kcNA/C0ECJre/DCm
YxU0aURR7lkHkceoz+jUkpneYxqA7R3TM2Ippwx423XsRfjiQ2mvUB4INN7ZRLuOPk/D7+N/b/n8
iI+GvLQ5NovTkJP5P0pOFTEQ++52Ztg/fDpUxXNYtA+EIe28rc1FHinqfR21WRafH5wyWfEX0Vgb
ypW2HKjncu0xQ0fVULS5dBPBUqMweGv+i/A+VQvsOKZM6OspSHSp1GQdrlrQyprrhnKbPoxsrbe7
jGb0wtD1N15/eGG8olUsM9XSPYT+cJ9+S5TOGd5NqMvv2l/QkPx1mZ+Z3xOwFSpuql0sFWv6ePYC
jpEWa+2cDUUPcuFfxrJfSieKMkvLOCCL+oPsSLLHVm5KHEcYzsC5xDpPNpD4QvYBBwV+0KmVCfLe
ZXunJlt+rwuCekdsgRvpcjqLVGD173mA2/wMNoR+Fa+pBH69SXizF+Z4mZ/HhM4RXeNPfVqjDJxa
cp42jGkyM20KTS0Gw/j0RhJMAy6etIm4FSQldmMHsFMQsx6i7pKrDOZTBOytKwWy4mgZpz4ZUBjc
BpGp1NRQHZFv3hVICvM0tZw1hV0YgA9faiNwEzzPKDv3C+PkxawH7gT8tO9dfVH1aSIpuBWfWAHh
o+oiPFwSJdcdfOyIJ+U1B4bFRlug2pwHVxn7xFgx5XK5QVaiQnrXA0yvG72iwAuKAszDlkGRkkF5
/JJ98aXMDgMLhwff/SmDArARkLrQpssOOkJsvPyJBMmUkNP9dosQA7WcuTvIEtfORljgBpzU3Y4i
lzm4X87LXTT4U+lZIL5vFZTNkYqOVgu4pbuPxdwg6przcH5qR1qFzReutj7nrEjwR65UIRkB4OXV
1HRXWj7SMtnGZ2aMTIzOlHOzzuguC9KQolb4VktZhcYR1zYUx9DSaN/Gyr+We+miduchNmzyBckp
pAUerE319IlYNlHUgF/pUk46vfNbDY1CDYbOFLUggPp0ZBboG+X681LYvgCh/Tsnq8sSLAtjTJNl
rJEy+GKWozgeUDBrQTeZvCccG84r79N2BKlumVnuPBeXxakZoNVQ2co8DEqB5pxdVHUC2zba2xnP
ZsQJ6/s9i0iNsiuvC3mM5WxBn4eamo2y1yF8uuzba1ycx9xmS7e+WigHDBo+8PZzZuxCe6YQLWkU
Alny7Qzw79gNRSfp+o58McU5tZcFURRJtyBL18XJ9LNPHQgzyy/xTKHYa/v2TL/+SAtSHB3hecFz
A9J9jRrTuqCZt0+kyAzJy4tSZu/qe3G4yhtV9ZY3JQE+P5J0qhHjOVafUnQI+uV871cYWYFpumUW
2cuyupvHizISPMPz0DSYxxfqZqpZ5BTnnxEUhQNu8GfylEEsrHgoYMUWKylhI1ap1ra6Bp3ld2me
Xoc36VH4++7peOrz/gK1jcqEmZDe6AdG5truojp9gESo4DUvli3FbhsZ8gy6js2PyO43fMj4sSzG
2bVo6nfbZGuwmB291kM2oaPYm3jAK7eO5kEjwhtJsRUgQXnRNUTaavuqoKtA8UNN88H9tHbR9SbL
ZivzQTNlZX2dhJzX+c1H8FpRajSEYDzbs86nBtteAX8etdEHbutIFS1nO2aX3WOal25uqvxLzGDM
yOWDKOZKObkNud3Aldvt8H5IeKa+R3OWogXjXO985bg4TP3UUSlo0mf070l19KFBiGe1sTBr8Y9T
19CTZ62ao1ggg1YP22hetL/JFNSmtrvL/hrGjtn85lBUowUpejLVvf2Ini2L30Zg0RiYydVVjB7z
tmkZlvO6QCpnro9sb1HPmcsubaNrZ7nOcXsyujVRpeMIWYhbdCtxkNF4G949EodTBIpvIRQeWK9U
1i6YrxnYLJX/BNBuhJmwpfraQ5Cpn6imeDz8wYauvqfDahMr89hWb96qhZC6NbTecN9RlftQ1fTE
4i3m7oZcw1Er1KZb+hnaOLYuy4LOBDPo182VMXWKf6vmpMqXTn46t6Sk/Vjs9nSX25DI1+u+P6Gl
CWThLw8rW/uowLajqYwhdqvm1YyAhb8ZSpSa8UlkryW+eBI8VUb7R8nw7O1urNW2YDCr5Z8QYuzO
aJzLj7b3mnXAlkjv0wtbzCEenbqLKcvd9Z61DfBVQlmwbG06/zlZ+r/PY213p1j7RJqZCaRZ2RC+
o69BGrXMOB5wQ0savw7VjndW8jGis2tORyKBOTYB5ZRm9SIFqr7/kH6E8F2OF2EXwICDQlpzsJgA
l7wlNdlzNUOvad6MIpfYIEk28NK7NAyGaPuaqYxPZyc/LpN5dWFhJJzlE/f8l+3gRDF9WjyEKlhz
rgyRMjurVD4dwN/2QrSTgXa3PPgn822Ps7u2hM3qFMoc0aZBs35nQ6XYmhqRnFzkKOX5D81jLS8H
jUlsjlC5nq8rjmWK8apmzGBeRnTJoiLcJHLDH758woH4qOsDcyYGEd30SfqHLj4YGFO1qoudv3oj
h5vwHuh9htt6k/utVYJ091GhlxLbA2ijGvOVHnmubw+F2zYcWiMMHIxx0B/6YrbNUVTVq8Q3xH7v
dryxM7qDQkz9HN5PVLPaYPyoVsT63WA7a8FX4j5zqxDybcC47i9QZKEcVAS8Fcrt7CslEYqJFope
9zWzvjPibWhZE10XLwQ7nS+asCzAln3gqJ7vr8Y7maIN8pXGn+4uWul34qblqN26KT0zrvKQ3NHU
8ETRrBNkl7o/9UM4HMLx8ijZ/05PzuQw/EgnuWQE2dC+rDoQwW6Awu989v8H9+8VSx6ymcAWfg9e
hOCI10iAlm8RyUtM/M23dGDIobdtvaCopi1cIdBdQ2rICTXqcQ2x2Zt2NJNfdq/vwzBzz9NdMviH
VXEubG8WnEMVmoFKDFjJo+3enRubTqKevWvnZOiGX656Kq/1Thn22g+I7J5dYMXnqrGKHVUaeg7M
edBnxyrtUDlmCS/k49+S58OHc4nLnirqRmRE3ZXcZ9pnebGlNncF+YvfJeH2mvntba6zJyPaFZim
76Cp/131QaUB9lxjchS1Iu8fA5Q1Vevea7Sd1VzBr7WVmMijvXXYul+G0GeTqaucYgNHYal92NN8
7XFXDtQ6i98YiiQW8ZAMs/gBIP45fn+S10GIegZmX7xCp0QsomflxuHSYOsXJ/BYrFkakBSPmyTh
R1xVaihq+JOPTgCM/NFDXSZATM13FXdYjun7w03kQ7OZ5d9sdYuIAjlP3vj95HgW+WEEmatUxYU7
YsLg2Xs3Tk8f6N1wTEkVrzQhXtjdoEjbJM/Mazm6fBF/c5xIs1sw7MNM6mjLrZK+BM4teIgo1luZ
Q3BSVZNWjN6NbU3tRfxdUljzS6zWCEhl6DsolyafQI9xIM6etmHhKjfv6a41a/6zAOeCalVDy+GW
myi5NDi0n5ZurjhOx7VHi2DiTp2G5aLXOcJiCnll/ZVSu6MHyGuIHqM9sjKt9Jq7NupktGfy9xIB
sKKQAeiARvCpv2oncvEU0Qu9Om0CGyC1Eo1v1bD3IoVoCR3+967/XCk+6XLBqtApoZ7Tn7PzecCT
Oo5kH2EoesTit6ZG0ri5JDOIuR2mWxuS98vMVifdvBDjSNIBU2vdgm0i47ggxfrgHo9YCPK2TlOj
iCklT2iAU3qqN6+joGLT8g7zIFcJZxMjJwEgUjTD+xpkQNQBJRyGUNqYFw2wSW1ioJjlhfCQl0PV
toza1PQQc3XgF4tEsWDZJmOaTpMpy5mtBwCaOXftFbOHZnJXQOCcrYJMoZPTejwnMWtHB4LaJAHG
yWzT5fTl60/CBfpBKJVleIskVb6X7eo6PNu1RJyCI7/+6nA1sCXuGELqnFNp9L29iby/jreA0CKF
824CkImaHI+DmSyMegOZS/m+ujoK0qTs8vA/GMOyZihloWH8Lh8048fnAZna6Hg3eZcvRFMajmg0
rc0wLomtUBMtlGl3BCpYXI0/3fBN2aX9/ZwlgcVyetoCw9q3Yifs6fk4kJ14PVvsCVPmNSzq8Vfj
pCU8aWjb1aruoUj+3OZVkhZMSASJEu5X9eqO40UlNsbdhq6+mkg6evXWhWwn/G+XvDqXH7YKgLAs
OQSrB8j6KVvwv0R+oYQZO14HdC8pn7JJrxPjt8xW7NFG5nDw3nQfAzmEt3Vqv73x0Ko9+VpmGB02
7uir7hFBsOG3Vpw55jvApkMAEOZxdsCfPA50DnlmOTHLlXwZw3EY+tj1ipxjq/Et0/xx/+B6jK33
DdHzvjRNnnt1x2mLPME0ugm92x0bt/H8R3SJs22TwemyHM2fl/oTfMmNMwxVN7d64s5w27hPL3jD
NMAXXx5TvV/Ac8FYeoXqMTi4h+jZYYuLW4kOxkmdam73sgCf1M8FYYtVfob8tSxQ3nBtZmaf9Duj
qe+y/R9O+kJaEpoowEqruNCDka4Zmkxryzx4ja2lWIk0RuQO95sdmpDGL7Lwz8RmMvP1mabzDk2G
k4ygM3H6qlmDYjbL1jVIR8/zFD1YC6POL7+ixtTz/kEWOO1RQbNpn1r0P/bGwJc7OCIbEbMHe1oh
1m72rWAr8NfFHU6pdfRtxyMl0gYUp6Pv2Pt4s6eZFFA6h1zFFT/OzAH02OuUYAOiMeSdQCT/M2Jl
b5i8KPnEAhMP9mUQRrr/wQ9biYO37W36kAh+f6pqZ0cXjECkCw6M9J6w94CaeISMYwEoCwMHi8RJ
rCwf7sTm00+nhJjFH+fuoKayXBbwTDYhtBUdb/HozTjEOswCzr72SvRZLZ3UvcdfFgtsak3ophL4
HmAmbXzwh+9MYk2dtcgh0uwLTN3h1tBGSKriy4XSyrE4NWflVgPanQJlWndBD0VBjDuJvF1UjhSO
6t6jmmr3YVsSVs3dT7WyB3LTDVLzwsnSkyJu8vi4X9Hz/CJAbqgwM6uR1xQV/HBXaT7MzK2/e/aa
O2Yuk13bG2dYtJBcT5dIhqwuemb35l6QBDqrKiDnw84/E0dQ89UsaJ7mVBndKn1N2VY6VC69GUXu
3ZreuL5V09yzD0uLQIWpG40j06Yw9Z/RfBgBmBHP3+iBw/n9SURdqxb7ffS946hnaRHwlmhrQ482
OQgKDvwvR47WCUHJmthMMr0/SbZ5GICPRL9ijh1/Tup4b3YINollvS8HT0ABc+0eYG2Wdq4zMPCd
0LS7DBU6c5cT8nxiQpgg6cSBvcAvNXxzLiHrb1JB/Oo5KQVNYSvaXlV84brUF3JCKdAchpl2FI5B
4DLJGUOXex01+YgN32rZ6V/vubnxOXEAfshf70A+dvhh0J0feNG5xpEm4ryPZbwps9TOy1QxNSmQ
oFi7ES2f2taZ6+ZV+7KCSfMDFawsDwTrxa/jImTORjjto5xmFlzE5hSaehYlRmbpvp67x4TyrMHH
YDTy3T61aJlOotXoe+s6gy/qcwDNPApJxtRzxqSTw0B1s9kJlQuDIPyxxm2svZBCnesjQx77LGQO
/pN+iT2ASNPZ0PtXbI+8niQs/5YNjmxyEDzfwpIXmiLomrZTiz7gtQvjfFUOLYr7LlpHAcsNsmvK
YvPrGosGmx8RxzrgBF9ejmV0Vw/KRsYd052M48i37E71lSGlmnevEdrd50mtZf++xdb43Jgr6Z8d
SelrDk1ZonyU54wMRRGs+VHl0yATysPr1EMq2M13wbz7yDEKwe+Wqtv1NDgbZedSPNP8ZOC9Cuql
peVod6RTJM8rMJdUHq+77VnW6DrY328+xh60m+E13QfnsU9zAluJ2jN7MRWJs2MdglqqzMMLIRhl
dfhWtKZBumrSU1PhkybCy65XLHLPmuq0cEWB3LVOufBxj0CUJtLFIxZIzurVr7HTdtgkoqOrhWJv
qzOe9AGB6NdYuxnZemOu/6B0/Bczt+9qQUjknqqXb2cW2rwKXFGERF2MayqxG1W8JrdJiRJf0IO9
teRDnlT8TRP5Y8lHqS9mkSlrxcFjsfT8+iDwHTh4ZSoZiFQfyhoZGkEYZ36j5f1Geildk2rWoIy8
klDtmLLxqJzqAnex1C0PYSuscrH+sNE64ZT0jBN65CDiOmthTQIOAJSznzorGNatdIdjHruyJzOD
vidUXvSHHu0iDQWZuVPyRd3cL/HupufpivoSfT63ZRopfPH1qW5IqyYTMiB2Xd44TLuc6F6eUCvL
/VrIUdmBJF8jZ/+MnNVg46KW800X2VhdqJNJp3YkKcBVNJir3JKOlnDEJ0deHp0pbw8mjmtjPCm9
3di/yzsjj3/CAVBe0GxeBLPdMH0nWhRw/gBD3t1rofoZnvW6DqQGY2PdQ3T5qKg6o3cNR3IhFuWI
Q1N3jbDY5DdWkGX/0lW9jo9s4USoC2hRLZbP7ViIqhJUAt85VC29ctKKr77jJXOX+NlLW1rZ0OTm
NAl2UDjmAMFRbgLLNypRPc7KvJbm3GVXy1AwHPulmjuaaZ1x4RhVSJ8zUbD+BG491PqxS6cB2fZx
rI3WP8LXiKIpCqZ5ZxLJ2zEu1WC9htrxYs/ZwR8/E8zNag5nXNaqCiQRSUaB5l8opSyzyPTUTdtP
aJHdTQQLmORBMZl3BfW31E/SdpWRmICh8Zw45j6vbXT1CJJt7QnkOzPoisrpuvULNWGYD3o3PLnW
1txGgXPutnq/pHTwaZZ6YTE3TT0mdOshhQJKgxawuYZP4jkiMY2fRhKQo1ZBWWMC9AjdD3Yb+oOH
dBbUgHE3ekHLLRdBx3GUNfqAOmX9RuYFFOfU0KhdygRLnj6g/gIxqBTceIUiKLP2CxFQYfgDfy8p
iXaNc8fkQpWhUyd9DQll3TBOO7NWw8DTofLc6YxLl6ENQWs/mxG7907lT5tJdYe/K/WLPlQr/Ixg
23uyLp/j3gVy3F3A4oP5B1pKh3fatZ7cSYVTUy6NpOR53Pw60ztmaqCfxW032YxlFcro/Yuic6g7
XmWu1F5DgUbzCqWq3SwIOfrcAoJqcpRPUsVe9d5mqTLAcrSRDJwVB0ZkYsX/6U2IJ/6IW4FhanUB
EQaF4sTALTAw2vq0QjDIybimkKQeZ8SL/VaoPN+W1T2zTap4a/j65kePd0M9UdAy8LNo8pNLocz+
Ih3TeK8KnoXRVT9Sdq2W/Bfm3rENrzRMDNdqE53GWIqFpG5rXCPhujWLekbz84ABVIzVVbmxNoVd
6xiWvXrtTqPfWKDhr6bvrNMRY77giBHxW975kK8KfAwpZwgnmBiPy2K+zdw7SmuRVZVfTdKTK0OE
n+wbqjS/OwYUizRhKPRy4ofaX4weyjq+eOxViiH3nNGL86wmvjN8m+mr6fqL3AD5EHUZsQUMUJpx
34oYm1nec8lIaXDlrNU3fu1H20U4X6r+KBYLuvuHFDC6C1yPzJzaPubcaVfdXgveT7JPf/aZYnyQ
ZxwVEn6mDQw5j4bQCl3KJUD3skds8pRoKzGzMs8t2nYA7Z3IyF60kXNg6EWstdth/bFhDLoWJ7rA
oneh5b1lG7bCs2tedE73x6QzEUiBssEFUJpPEfba99ktp+EmwisJ5hDRFoVJ2k8PWq0DGM7P57jt
PoDT16KFZW7CVdOhoaeEaVY8lXIFm9pEMjMByifiaDy/H3I6DwjC3FOaspITYN2uDG7dN1eM9aZI
6GwxXvZhvHjG39lc4Lwo4411bnjrPvk2nKLoGX3cp1mQME2y+7L/FSehK6yk2/UdMe5EfRnyztUZ
HwtkdsbOCqt8LM5t/fGVdOS4zZDAPCem0cSIOMboQ3XOvjUD5g4m+ywL5uFgTOvIMFPrF8WSHewV
oRvSUCY1Rt43R439+vjGfWbWc7nAu1rwnPwiOyjAfmfU5e6zWotP71tdwSkejnrKyuFU86kdxqSr
g8IJFztWbc0YxjzZCAV9HH9lujFCt7oLQt3vXDgVTzaThRtJhBmbZL7vWr/kO8hQ3+RxnfMRQw3z
tEE9CysB1MkZVZBqM2A1WjUHiUXoyNuZ+7eb/G7acoVAOAEfbVqtpVE0OrBHqAVGNsGGha7s4LFJ
XzZHncr/oMk/7dHPj7hczU/QLNGmAHPNrFZJjH2sTpd9wQCoWRknGNFN4kZDLCEH+LXB+j4UiJuY
l3BDcNc29XSEDt44SXpfOR5DCHD17AREY/BMHhZkEjbPQu2QSN3U3y/r1j0g2lpsmnwwHhBz55RT
GrZfaSMiR2Ey/iqw1gut34TFh0d53KC8T05120EkfqzmyNIoc4WhlS7HyVVWUP64vaWcyRCeAa6u
rC+WldZQeiN0VxE1JRoUbB5VUWHelhJfYk7a2WmU/P4jNf10E9zt56P2U6ibEDrzTmtyfLDVWnqn
Yhz1S/CMkQEmCUaUwZ4VTLiBbCx43yiolzaCl971y6IXTXCya828wVOtI26n/EVqXaGkfUlqKGZw
/U2P/4Lk2eSlaQmpATzXPIgVgPs77jiDN7fpuUDGws9QSg1wP18orF7IOVMf1FcHFZfw40t829Wt
U7ryBEYyN4RX7RzMjG98fgMIuWFypLfEs6FQMTLjoF9pifZntTBTOgPzDEn7TbSYlW+T4wkIvwXo
OXGNru4QiAtNm3q1s9IkMilp3gQ+Lovp81Yk4y7GYcNZ0SsHlTIHyzZeIYT9o4a23Rl0IcjJVluq
Zu2qU6KBo3M5xQvuvLM+1ExqmSfIsgl6RKPp7LdHdZOrnrrUAiIvKOxpkWCeM9eYoouXj4uqVcPz
0pRZyqpPYiTbDpY6/3w2ngaUvGKExIDR+hYFTiIJ2qBqEfkVQuWM1UDCIw4MKDjYHMwZumROkbKL
VqYeHaeBCPTRdejjds972wzAyDSrrMkoZyUH252QBmjlCpP9VsQxXgPYeJJzFVPWxlSWoaEvKfuL
/sn6hHk94j/wZfdaKPasCue9UR8kG26SBmaQE0l/6MwU02YhsZDSGJnnjEHGVL1T7zJ0nC4xEWHe
2uTnUqlXC0Cio+YCGVeddKmrwum2OMAtjRR+3votC3wf4OGVGq6ENrU+lvTQclAENIFCfUg9pwaP
9GiLE2tNEBf6mdF133B0AWJ9qnFm3HyNef2ofx4t0Bn8/dFBrGWQfaaW3pEd4YcIH/Qsijjqt0xe
R1g5GTDBxLOJPJxP2rK74BmuAmKGYk4OiXn1V5fudeTvxdLxveVa/REUbZzqo3mjNU/fAiZ8B5CZ
BvEJuSVLKN5X7A3T03DssWpmjKlJvq46PyjAgXild85CL117ZWrQNBTajzxDL/9WAqFqhuSNysjT
lAs/YDdYbeZdPmjGn2edlbnA0IU7puI2y2qlSPgN9H6U9bhTPfKoIqzUK4KkymQuj6dD8o7gIUAI
MvP5gKkUKi86QLU8AtesrpGSNe6gcksTtA1hRxfvGH9sKuIAvOdY8mxbUkYfpia/vVPC+FaBrUzL
QpGr3/iEOagbxHQdRQDvql5LUgvi48dI4rotEzhkj2DJnr1y9vo2wrIwMnf93ZrYXmBNV/X7LpLJ
SwOOpilF3/u08J43oJc3CCy82R0fyjJdWDTbMIa8f/Dhygc+7PsK+TLEg3ODjZkW90UcDQVVlwuG
Q29oT8gcmQDipzWW4oZSpFxD1+2CAxyPUd9Tj4CTANKwr/KwUjYGs7RwuPz/xfPqaPNis0tUe7k1
+luPw99m+uwIUS48yjRPR0rN6yqit46RkXBOgcfJzmbZQ/M/Rs8VJzWvRuCR2mHs6nbNWie+5BkG
GCPivsUzEa5S0t8vY8U0UFwvDyl1hVWXwz4Pov9ow2TA1DdTdkvUsbu/+O4pUfxvLcjoIKx5E2Sb
9VgM9NI0Xr9RtQ/G+DIIHFkgW+HndWnvU1CbWVX601KyFd+LJ3VlMKJWOpdnr+yk3Dj4dYQN/hmS
WPAyqQzokh2Cv1c1wOLuOZpdF/tJi01hG70GqM36SaD8tRdF+SOCc4wS1DzdFXmB8eRmNXq4vYwG
mwQW3hr62IKP2jCnKiHs9WQ8+9a81w3jdWFv/leDb42rTGPXAJh5qgMDlSV74riLm23qBd3Z8fHB
Q3H6mfmrff9WCyW+6v1UBLmiE3ege/45HNgdc2dkP41HOfVn3MVEgQE2UDG0VpDiPwU2kIyMg2vh
2aIVP1SsCMjlJU7ouyek19YP/TmeM58yZY3ngpT86c+GA0+Q2NtgrwRydTMTvDkQL8XqZL4Do9Zn
uZTgl4ptYKjtPINnnWgFe3ja5LNRooVlxztfbvbm5mdEiV9iZBy/shHwJxKx5CFla6/VfLMtCLy8
5blNTGdbCwEWKN1WnIt5WY2ScarFFWcgZAnZ8ND4FaNiuMX2zW9U9gu+ZXjkfL8XwnIfq/4yTRYj
hII+dDRTdDt454BXqgdBBx350u0rcUHVt2aWoFjqmQEYGW5549krCWjfb4fctQdYblvyiZ6iuASt
ZBMehQaF4HntAHvZpJ04nGBOLfvOpquO2X64CS04cQbTp9Wbx8Sxafshzpea0kTTfdcn/KLwcHSE
mxvfgysP6AADFmx1bTFrq85lzJrVTo29Sla2Wwy6Z46ZYbzqGJoSY9qOoseeZbU8334H+5h0Zlh8
HL9/gM54bxPjO8ACNt6r1f6Bzu47pMbSWOmRI614hZGsz8ksgnadeOI9k2HOzdMdnBVrjZ+AXsNf
APg2TGm1v1q0plIJVW1NIqbjHBcRbFXgT6nyF0tJb2C9pY1LvCC957FtI+kruxhOOUNNroZ1KNap
9kYbzY+3GH7RZYJQpEwU8uREAuIR4m/45E54ICnDOsNsnDzBB4vyrJ6akVL28S0gjMD3C7w5XXwo
swrK+ifBhM7ahyY5eygJqm0psdHR4taQP3uP6ESk7oG6+T+fSe3IEDSoCE10CNC+cC63MNgrOshX
sX560rS9kWIpZwq0VRHSPkTyRZnNtYrzyOC4hrq4yHO8YvlhrUgh3eazL0b6/oaYmOCQ3yudH7+7
uD578gvTB3/gAik5Tn0Hz1sQWb2R4d1yGsordA8FBYaUnWo1ZUkwdkH6F6tN8h/wNP9URXhUoURY
Ci1nVEig4uCXwiQKL1cNx/OLD2DmJ8onAUiDRBgmi0O/EQLDvJGpAKEp0c2cnMD4v3uyL0O+LhfK
7VG2UZV+upKg8Wjb7b5qDHbGT5Z8PR7AtwAr3f7FP0waiAlHQCcL9xkFW8k9uKic4S7A1ig9le6L
32VJvxtE+L1R5bKkwym/XIBb57Ao46YgFtFPn+QqPeXVlNFlLWkT5SePijrcJhBHUNhY64YSsxKe
L6cDCDKxOdkcr7qOlr+jNhBz0z73fo4OmZYCcm3hqXNQtAIDChUGawAyuIQOm9UZst0XIclTbnZJ
KwbLOmBlsoGwhNLv06m/7GLzwrVRixrNGCkrJw80xqdAN9iRrzM6wpY/0GxcbHPN3p0WUbHtZ1/+
OrN5b3e+7Ms6i/7zJxdelZ+QrOeSjbKNH25orIwZKIfpHO/qWD1YXqLQ6wmoCdQjjS693NWpteTV
SSQbYopzvVxqSoTnjh+QD/sZVv13rSSCaNPvActWNwLO7Tg1YfAJN2GAwIBQN/SU4p5pZ1qQrSIK
8saIMm8hvg0jANPYrvHK7cWsIK09Ju6h47y/zvM0HwBO4O3t2KNJOL2vCF1q1nGi4xlAs0vyCA77
92rZSn1OpcU76Wa5g/0QLQYPC7j9XRSfdLnuAzo5KBk54OC7z/IYe04fiq3yPRA46M3vapsM/Khf
Kj8SuhC8JXx1eSwBxuFc9rjkYsU4251F6I3UD0aWeS8KemtoQMebifrhEGWFnZY6NPjQexZrEOm8
X1L3qgmdjFtZa1G/gfpD4B4mpJi95G7V7lKHJ9Sq7fVmvf2E7YOU6F0zmHXBACwcn1APOTol5Dno
E5lXNvxz1GPjOnvqXnIy7xZXKntg/goqJAXErHAF3BTREVxe7EwugIIWgco6JUc+Qe9oV26iTz+h
KqQ/PQbAh61Ii8YZDLG2J4nGGnXukDTzDgEUPxG0JAwy1yQL+Scpzoz/W4sp6tXik2v/DwpyabeF
VdPETFs84OggVGNfuNP+uxbTKCTfSrLfSJ0M71tqOvkbWgiElwLqTFO6IWWNLRFjTyiVdk1CwieG
CmXgi6RE+2nO5R+v9fk42aDeaL12c2DI+axuLtgJ2fe0ezta8D6tsPUomrA0NjeRMbihwCy3u7UY
SWhNYVDfWAnGnzY05zTBEOwZtD1/h/OPsXFj2ZNFhPDDaVxVaEsoeYTldGIfJRzNolNHkhABIOwe
Vq9wsauIsqev/fz6dUiGdaYVsErUayhbEGwwTTPm3peyZhKkaMLzoD6e3SduOzwBHXuim5izS6if
Ez556oyi8GmQmyA5CeeDWFtkbxRrtD+9RQtgM4ZH11335/S9Nb9ZuoyKkzvI4EFU4QnIpOlrIllB
C760JS7qV08TOOOxvWWJ59Z+F4DRKVYtnmU8HpdekUjiqeiQ9ELNTnjE9yCc/6a0q/jJYuz7USrP
m/Vb5SpDskdWwfulK/O6hIXqJg82CDS1vYh/4qErwyjQhM1V3ZFtMtSD9v6X8gL6WnDKnKztsanu
QtVBEnA1fd4XfVEqkHew79AvshtPJdeNTroI9ER+l4Yl1zXYCw6ONo1WJhS4wfY+NW26+683S/Q7
8dLtBHFtDJe3V9bxOTQ2uTrT25Q6HAfqIppSYAXg/2p+PyAbUKEpl1iWVBakbkHo9411BVvpHHb+
uccHxIRBhNJvaTkoukXWHI5vNFFuT/OZarJKn0C2H52MFk67eD0ZYU1UOPD2on3ji3FnEorDLBF0
K2YSERk0i6B1HR7NDMGUzXfJd6ebZNP147nlH1h3YOFWcnQuXKf7uu2B8O0wLkDPqvUPoV3+5fNo
6Yz1WESihsweLeIbhZ8WNgocLLQGjS+HsW941byVnrBE3E4+Jt6C2uimqgvJNgRXTJok87DCxuda
WusPMfnrcNwr82cr4JQ9SzjETpYDaiMyF1Kqcxp34yoDFLe11+/ZTAShGu3tcBTnBmP41ufS6A6A
9j7F93nVflPISciwn3ntfQtFHhOaTEeoXIMtxPEDlQslwFfk1knzERjY8vmPs8DGVPaLAvTAV9oO
nUCZidrFFtijugvYEUQFT9TgfvVefwTRSn4vapt1tURvWrMMb5R/1jVi/R6+l8NX7m8PfgnmTD+I
VUjql9X6zxVcJ7+JKD6LBTjEfP3BIw7Lp2NoATNTVVagTlXGzmsXjaqG3gLA7fWod43NdfJeKAaV
lGJ+u4R/SstJ11AhSQkG+FVfsHB8XetYpWvFoE7MEkxksO3tWcBvf3sXrojIOvcGP31uHN4gKeTE
eeim9gaUPrr36QnmaYPY5H9A4ar9zZyFDS0XLGh8F5qT7QRaAle8EdkTjv97sNvPyJPmMcVFh+XO
pCd1oc3M2EGfY82uFuThj8hnM5eyp9UYMba/xjiByz5QqCoXgQszps2zquTtFLlrSG9FHZcygiES
EJFNIeNy62khy4I0vQrQN9WVYMQXcCLAI+QVPJb1Eqx0CYdhK51K14L2niN73l5YkV+zWWMmDPKu
EmUBAv88VdfuChdA+5Tv6LpgtYCdg/U4YRvbcBNspB1JU6WHkWLzh4TNPHbNI4v3xG6a242Jh/8Z
wP9CcyjZG8n16e5Crp61CCjSH6ONZ3WV/WNPXM2z0zhWhdG/5+QrmL2DEBzWLtwSe78y/kEtW7pZ
cizrqkF1EoJERN235zyftM68uUDdgMhuP+Q7Y+6kBDWH6V8LjA1F+boXZRflvcaumEfmiayQN3sX
AaYbPmvyQ5vALGetqQhQDKRUqhfrVSx7fmNNbLzUuiu54eeFWJQ7sSZ3e+np4KMDjJg87NUl7DJc
/ytWYfzqi0iewp/D0L9UVa9KmXbm86oYbmQa0oPHEmk+Sc76J6oQrMXWPK/65kjllBaGUsYYUt3/
Hn+jN3vzu7d7A30kpr/hvcK1OvfgQN5j9bBr+mQtrbc5HNNwPoqjf3N+DIcbrRJK14syO6fdv0wp
iUgPkueArCtjneGZLTjlZ7NiAe9qiGBr09AGCLzoM9fNjZg/tP57B1MDOhTdWbcDGK6Guk0z85l6
fgzjt55CNaUBthlztASxSkpMzlCB/B6Bt7mEPiFRSNoxkXzWH2AofeF98c9MBkdG1ohRKDnKhTOn
Gsg/WlzdroufV4i2zL7M0K5/fUISNi09XvIi9oliin2+PxXHT3H6B/BGqRqC8kY3dcg5cOKRxcZu
tgYFTrZemqGfDYJb9rlY6tW9zrKt445cbzYvqysrIF0SdFHMKUKKJGT/WXauAVt2N9If44lPGdDA
mff4t7KVa+X6XDmhb7fAnLVQy+2kwpCoqKbN4Rl1y7Ke9EPJ95WkGq566I6BzsvpxYS5DSsUD26W
mEMwMM+jahiouNDTy9xY13T9XarqdaqOGbwHiUZfiHGXdsEImf1xrAGiR2CBzY7lVhDaMJ+/YG9d
jPKEkxZ96Bj2VyAdyuzlB3P0cdNeedpxtTKJVAId8LC2x1YGrxnTo3vpJjji6s/tzhj1LUrifmfc
oJT0eF6BHwMu2/Z7YyZ0ocTJPKzJu10yXQehocf4hO1gjnRa4XbM+vc17eZr4m2GDvo6HjIVrQHX
hNupfPCKrgj6qysAteg5wcCL2cjZl79nyUanYP+pVqOs/GVcJpUlqbE5rxIaArPMR9zjVBX3oTKk
O6ILooY3p5iEkCFpbliEcZVsYrA3mkfy5qRYLEKvYIBBh44BlLOYBSX4VhVBX74IW/Qx/mrnw+Ur
48LmjD5nsusHau3P+Fn1pGUo9qSq+aEljrfYoLrW6t1OG4l7Uz+J5l0y0irF1GsAJnnn7e/LrA0g
+9sjcM/dXvx3TygUms0j1AuF6lnT5DWoT3vnFIazYZRX2zLriG34YtJjkmIr/WwqGPe6C66u+W9/
MB7kFgU5rJYxEo1FLuWmEOP2rgJyqfpbi2EYrnSjRwfnrxINDNQJIDy3qCkw/gZRHal9uW055nX2
5qloQzGIILNbMCaZpdWTZktqor6vKKvPVNqKCvGDepyMJ84DwE2AmldujatC3RqpJmhTIqlwaSbc
+TEyYGjRaPzNR58S5ikLrsdqQwwsrr+djsV6mh3y9zezGYIRCmdS2NHokiKgrrw+j/MAa6p7B4FL
s11pQ20aL5L8VVagW4JFixELygrE376JV37xaxapbYPRzFCw99yKw7XQy3Xebm1UcA8q+ORoKQ+d
61iOmm+2rOOI1eCdxKbqRgUMN22EKk4hndFSearWgUaG/5avLzxa18CglWctg5DCpOSXH3QCjrXf
aYgF3MUy2x38D+lc0BgnpMh1pCikf7l/yZgAzcH+4rvIBkBneUm7LWIrDtRVIuawAt5bGC2/c2bm
DxvM0q770OCvCVUsS9fW3D2yygcVgebg82wQJZpVQiQ69IP2jEiQYioBfoUaCGpGsMLbjw4Zk6Xx
vKM6phdK3OIk5TPshuZ5HHv5LeNUYGesVUmfSaAep5AkNTYXHYSlhTwPpYAt96BUxYNAPQ/Jgqs3
WajBGuS9el9+8y7h+P07QT8/YvubCMrW++jqREh2x8S5671JEY27mAvtZTE6bF4kAD8rccY0AE4I
l6Uf6a7V7qa4Ac11hq24xXbpMM4vKC5tHst/rDu1wSD1mJVJw/VDcgzYl0Tn/kC5PoPxM5KeC/EU
W6rFnVpGtPU1Uw9yCe7ev0uNAUDkbVPInE84JPeWrx1q33PaWkStSqDxXzj93mPoWyIkeGOs4Bqa
L1pWxHWoycCk2LtrOBxnnHQx3sLDVchYdu5jCvuzFgP2t2uNlTTwOCKmBIU5vurvtXwkaHVb/Cbj
WMgR+GLAG+fESpv0zkf23PE5VtgjVOs2iFiqBb4tk1tSyJGC/wXuk5h5kdFQmZljHABURcQqmO0k
pqTcKE2QfB1pLvpLwQ3MvGUsbv7dZFBirZp6jWdRqFyNbEzMFsyfRGITBBBb1wGYLgRx+5nuWNmo
IFm0hCsbE/Hi4msa0jj6NcVcrtb1wSw4dCgk8cylTnH3pMuQTWxYCna+fx2cEhN1x8nSYeJSuZ0x
5UgfqT0DOhDbqnhmaJZ/8jX7x3z/mbqlsMs/B0YZfBtwNaYBrg0H9AITH8ViaCkWgxzLy9h6BFMn
STVznZEWIJAqcHZgdIgfRRLq4hWr0LNcJj0YdsT/BXZ9zBxS5bcT3BoZOEEXfrONQmYnRtNNvFJZ
OjLHFKkwK1a2UaNVjipYCmiMRz69bUEVnarEx8OtSRhZFeqc1+x8Dx1ssTVFfkocndn7PYnwkWNm
UcZp8EIb9K8Zc0xy+PzM06xLHnWkJ+8o5nY/VWOZAO0T2MYTsbT4CWr3ggNHpaU8mKSTRUl5667+
pHsDILr4Vus8/hTvy7av11YB7JW5GjstnyyF5z9/o1Uq99xBm9VIO4UZ2z6AZv44piF+ZiHYriaX
NbcMi0tonyMjeTqjKlDlu80I1Jp2wOl/O83xwy7Xq4kRhDuabmPVF/fhb9ZqLmOPE2PrKYWVUqWe
+hDZdz4/VIGPORKjEqzCUHuApOog7ofICK+x4c9Qgig4v5mkLMJTRt4flx30ULcGHHHY7VUML75D
TKd+/vIFC45l97RsdTAYzsGOvwLYYS4fTwV6KLb6bKSsFThM/3mf9FkR3VVSvyeuMpdAUbjEZ8UA
ILXemGanXVUrZhnNhjsdIkLRlebPS/MT7H8koq9nV3yOcK2He+8/WL43wlukE3BCPYng8CjlLPmr
w3wHukVbEAoPlWGNQurX5ojR/RhJtbWLlIeV2ed1no+L0ZsMXi0Yx9M3LBQV6SQ+FngopFW9LKTc
+u5Oicjtq3hErKrWINldx+0xGrgn0RWzIy6DXsi52lNRcfiNvHCPsu70LGYYr+W4VFk2N7vLyn/9
5qnGBX5g3k9YDn7l5hlUhwewP+uHOpv9yNsURbtLnRppHMxFjAxmrFnS1PDXYwbwhMqtb/sQNoUx
TPGTVar9/wtXBgRV5+CaGNZCqROJqxPYGC2iOL6GBJjCDpV7BKrZhUxGUUFLASPQWypyAGcIPZrk
7mQeqx5LwY4BJ1VhBl4M+CgkLVAnMyOGtUZZLueD7Xb00OPtyqANGZEdVp1MJT3C90W92h0Mcgp0
Qhw0yLdfNYTb/LitPscopHXHItTkSGKiRdlWqPnumETTJxruZdq1m1QEmKCxrXkIP1/s/D7LSAMH
oB9WdhV5a+dD9Xgsl/eAn5ty26z0HC5RLKPn+aXQ3EgfTwCcZx8zIM9GQ8vtoVk+1LUBNuVCNRxH
soF/xkIiFNxEB+TjLNOYwkQXv3MB66geuZh8Z/abSJ//HD9NKKrwYx+z1GMAIi+0smD7PMpHXAZz
09DzfP7qYYPIVFSrRj0FFe+GC5uqiNPmvIlj1uIJ87mzUhU/Og3v8sPEWCSTa0fAvVMU9vQzspvo
a8fo57faiZ77c+7SVgJDfiFfwtbK80IuFfTC8MUMbhn7phTRMaFINn21kDlHUjfwMvFtgfyON6qR
LVKMtqXztp3a4yGavCMMZJ9zd92qFquqVYKk6eSFfwmWA3p8VNVV2cFlCteCWpzQ8lNRRfXcC+JB
YuIp7rvk8sAd3xlUgeCaH4qNnb97HGYoqqynjFY1m3q6Im+jHO4MmozxvhwsCbGUHUFUgTQCZEVR
UsyAYjiMKkvzncT0BhvMzDI55VTzJi5QSpRcQWBckrYOHit4qF0czBVccTaq5HyMfrW5gtjtdPdg
rO7RHd055MTeiwGAvQ8iALhJZCrbTDbcMWEWBEtJRTvnUzXReDjfLf0bWDSvB5RnxUbrp3fit13D
5FOgOeAlkwLBIivS9/Vh1xlz/hGO1/J+JBmRCLKLOIjvA1wojHc+GTHpmuZBBxYSh8yLq3N2IXNo
YGgm0yuwlr/s/bTBy2Rv+h7m93DHWEcm4g1GOmdxqUEv4s5pPZ3rulCXEgniT22SOjEWIhQoks1d
/Vw8AIjwvNNGbCVg31SQZ2HIC5keoEdXK9bH7G7FefHkoAXflwLc5v0pONHwKKK3WvxhIZ+4AcHT
LopEa1eevOEsP7oRAzmP3434T/GJQJW3P20/x4GKeF0USroPi9/dukqUYjDUOGHxXy/7fb9wg4tJ
Ox0L5g85cbDx69EheiSRq1j1wPtTmcFj+QZaWTp1rhbLMDaAu9T0nBE4DBTtoO6JLDGdY78tkNp1
SML92dchW1+6IZ3dRJwt1jxm3CgHEl6NzMFfOdp1VZ+P6oYxvQCXeAkpmcO9JVo5BXEaPxPDPSAQ
ZUk1KqAkqNSSKy2XYZrT984zSZ984CZ8wmCM3hW64RN7EcPyEotAIwU5pclK3ZFc1DV35uClzr3y
ts2H4kcnQ4hVFXOkrzsHWBM8jZRgv4NsdD+WZxrOZnEnNfqzXiz2LtJazi5o4S+3KpVBXo7jxXWe
2NAiaQw4MFakK7yf0G3Z8lg5u/xt8Pwyv06mGF7AESSyk7B8w5lcunY6vBX9y1LOcAVpvBbff+sk
jhrCtq0wQ6r3A7fEZEcB//DGs5EuTXKiqpIKbBchZNUzR6guLhVfmhYNogVxoLXpmp415QC5FbL1
2rLDNuW8NARStYTyjvAWRQlE1rLXqXOpQ7JMT89Mo7mAhmAtWkey34obMlRiCEbAQvclSpawAygu
XjyubfCHj+bUK1hMHoTCUGSKsH9mfVSc2BQf7y61mDW0AkQbkSFOnrVFeWCPANp0C3TVcwwqfStF
v7c1X2BeyO8QK5+ueUABIhCxtP5k6h1OGKu/0xJPH5YyL1gGNzsJo7qxV4WL0POJSBULXMFeFNNr
pgEGj39wsUAV7InjIVprF1BCZwvMFVs92CvYuC+2j3AuohIXnjEV9z5XapJBciF2xkLAHDzAlU+N
UuTcajt1XiaSBCkR7kI/4k99p2lkCTYtSXgPX4Q2T+M8+oGwIkuReFPicW/q+yJfaDQK8l9KDksv
mo5SOjWIb7yV5BDvv75wl/kM0bHoWamI0ojOLZUhiJuAsxmgODhaKTeVPABV2M82sp/53oUKZOtX
G2sK6XJKOIh4mpTG1RidjX/3MTqJvD60KBX88kUlqj1fldEVBxLQuIzdJr8Fk/TYxy7FRjSl2JCX
f+hjPriAN6Jd6/5G4zBtHO04DNHRI51PNqmrg98Z4Yc2G7Qx8byiIbgRkneI1MpkNlcG1RnXuCjS
OIv7cSMrv8V1sHKfvnHycirP9jmw8tWqqfsWxN33HDMrGdKzT+bVtxKBltJolrYcyMrY+8RX8sFv
rswypgxy2DCncbC/AiryXtjohE4e0MaJ8GVPkQixVRVd7x4wsL6hFnkTF9rH4HQ8QLWwF1rcuOTm
8RqaBmmooy+bBs1ZyYWcSYPKGwWY41vkXvPjg/7LyBbsHg1QX/MwLp7+f5VDeUtdlRXEpOok7PiR
4wg1wjgATuEl6Le8f/uaT25T66YiYqrfwCrX1i934GhkMZybAIvjICjPoqjF7Vtpv/R49Ynv0+/B
b3Ilk7BrcvNRRV1rjaaIDUlRaT6pbC92AkrY1EFCJAosPsLYpSLgzXWcn/Kn72DRoyG1nNPXS7+d
kZ5y4D1S8lH1EUq6aE1+hboxCG0w0MFWr0LpbEI0E7CoZ91wApDuYMsNcgRvclDXx1PwJQF3nIOk
W2UtRhaCQetAXQxhKzoGMskejQwP9S+JXxlaSTV9EFQ2RM5oH9T6u7r6drrPch7Dhk9tdtPEjC53
xSPfx330kOicuyZ8SxcvQ8MVIWKXguExlH3fO1jc9ajeNaNlxZrENfg0xStOv9ijOwEWzRyG2r00
ynpLsKUf7/FC9Nv/S7LJI+E/UtLJwf+XDWig/PrmygJt0ohQHtQWmD5U0GqzdMemNvM0CVMkr38Q
SUXZMxy1Y3jzviWdJx1DLe1y4MsH966PQ1U065gN26vfliTyQXDbcMWut6LvcepEvmKCuLoFjhZj
qHtBxeH0rVe3lBZ2fNThoFwnITWAQ7nmOBEyxgKbbhlZ1XLtJ1r8gwOF1bEgzr8pSrA6bkk4Lq4u
oT81ccsJlq3jDrmFzG1rlLwnrNQqbgOamL5pu3dsY4nbFQnTbt4Nle/NBjH2zK1D0B5258qTgLsG
lgaHD3hvdZClVIV0p03zrBhtUWsykEso2DL/Y0IMzI6njIr180pHW3DjFd8lAEY4qx4nLs3CUtlH
qkao7EDQ9uD0PLiTokmZoheujKeDwbBwpOFbWPdyU9XnEZdzfc1usu0xmw8x5MWf/0y/uv/uMDH6
fDiHBIhlPT9Yu6o19IfPj+PgWWzI247S97w5IDaYdVGNKw5gEpp9eJVbi7MOBgH2wtY04vE7crjW
SlGgsibebVRN1lDzeWvX3iHW2Gvrxz6vhxnvd3QlzswOd8ECx38cuHyNU4CSvrzhOiBnoTLSH82i
x9F9FDArlLa7vhmjgMs4lnOk7wEw8ySVRmEcccPhWjrmhYUgYMQkee3IBzeK5/xlLvz2KidgIiZ9
k29myOIDrDFU+uwKaluTGYhuxay9EPmfI5Tt+EXzs+TjgoFWzEKvyAjEk4ckQhl5bkopL5WKLzaR
WOpu08J/UkmH97vObtGsqHOdbhvYIrTPBbEnDignJJZdlGr0yCu+W8K80/Bk2Z3lJc7P8kQya/gl
2JzeIoesRH8/3I6mwPATyXI8kKLq/xx/JXXMlFyi6cVIfovEvED2LofEtgaF9T789g0INta/OA8l
xgk4VSYNfux6Gwgytpk2E6J9XWs+D5AHexRMvUviYukjMEEV+JKEIWAFqDyufiSBt6tm1KZk6Zp0
E5QCDSnSTWxBWDlbNHIjnjpyVqLLLFSYmMV0JBvnlDvUbJ8BNGkts4Kt9PhHXr2jC2qt+ZNQt+Us
9Wvp9pd/whQkfjwFAqG0MF1yoFYCCX6hrdMC6B3M0c83n1gz6LjwOan5+XJVHngSggSb35Qv7+AV
523oKk/Rhy0nAE44bVWBq3aBi+/Kz7GGuRHKaxtPXsxcnwwkCmhUMK93nMh0dQRIozMyGF01mBZ9
b3OErSA+fNqQ4PuC0v8gcfoBiVBV9uP8vW0D4bkiBq+bXzzcF2xEQDsdZAg5zzRGqF8oBnbO9y0/
YHh8wU6M0aAb/dIgE+0+rpB1K3kAgIaASOkMMRAlcFM54kHzYln7r8ftwM/9NtpvzOx1mn/skEiG
lAasUItWut2o0qgMTYusw2rvB5ZaNUgGkZt/YPKFSW9srBstxfN/ie2WEJXADhgO7RuUyhpj+F81
gp2snCbiCjGVl4CJJiCWht5Wc5h5DOIS+hpYy5odv1oFfuRi+jzSWOP6DY9Nm6zbvSpNTQIQbvm/
RjoUp/XleCBKzHsU/hdTweSOJkZFQk2sN7mFadRanKL8bOT937D/wQktW+OSlbYy9XNgNK9/Z59W
AoFSukrCGSNy8lO/peoyvVKvyJb75ZxxIKMor3UODQxyeZmNikjnVZ530mU3LRdAm1KWnuosdrx5
XnUnQmo8gAnl0e5JiD5pT2Gm0BMUJ1sTGrBNOJkVrOMK/HhWNaUgf1D0cdaKmN94uBp0CzB+X6gD
wfFAYn94qVa8HBhERX7uLda8taQMECNuoPdd2F2NGx5m3yU02tGU3zHaNKH9yQC38C4rdOPSmDPu
17MANBFQwdbzSjgOzoARxpaxU0+vo7/uSN3vGmFHx50GTF+W5fW8BXhFJkG7Jro/vHH8oFnS3llp
U4vDjpq1/IxusJL30P9PDjSkYCOx1/oDPjOEtfIS5ycx/u8fWFlqA+LdCDy8xUneZm3I37nbMl4H
MHltwJQBaAWOFbtOiGD4cIAfmdbZ25t46tczSH8VJAwQeT62+ZsgG1pIN6XSlBtbN4AzIHlrg5yQ
HB2RgYRYm1oniGUw/z4mS+OGC1jhZ63r8g8LvkSwB0HDricnaNlLDpmXOiIDnSd00Vye9e4e+EH/
gJCMe/Mx7al/6WNSa/B8k44MbzmiJF30bCwRVl6doi4aDPS/Jsmm+lLbwqfV0hUcPxdoFHyDckxf
D6uLhto7UCDc0XGO40yW7Prk0A2y199Uz/E4GuSZowSaJHy1PXzvqvPDd/0iLqgw+Q230eCvk9PD
pre2DX0lVomY2iOENrAlbq5w4pipyaSbAWln9JDztbC3Rg54OuLm4GgTgmK+4nXbb5sKHvkWYexD
LkkqLm1GWad+5Oxg7egmA8xGg8YqGX7DTjbQdhDUqzZr1uVLReoI5Tex9RmFXEvsuFrkvidtOdb+
tLmL1vAtaCo2c3m4ZZGFJfTsaElPkmWHzlDEj+3MLWEuoDvU814Aa4tML1SAbpjhHftLadrkP0QF
Z7XV8EM3RKdhOo+zXONTXaPDSEKH3oFfn8nXewYl0JPajh56FgDbfxa8BVXaEhyWI5BMAfo9WNVl
PjwBMROAJ78G8XII++7Mz+l07RveC1GhzldDJRWtcHzw4goDYulmNYbKtZ63gurEhKeWrzXjeMYT
djCSP2QCBuI5/Rkc4MA/W8VlV+tT8e7jfnkwBE0D1cdBF1VP6wi57/a8NtBS+3bvHxycv38g2H3m
I3wN+v9u0uTzUNJsd+1ypB8QFbVv2TZ2/PUW5is+kOBSQ96dbp0QGrNTj9BLmM3xpTl2lQ1dsaGd
rzbqJKk+3mvTrHBUmcXIRW8zKsh0QXSEelPJjeJn8E2Yx/y53cDtlFvMbfaS7azs15Ix55Q5Cwec
PNoVQdRkNx45tC0Minujw1OA3BvBGKE5BvBhdRjHFUMfN9sMjARj5ZXHsTWjMxprwqj6dVYZmmk6
/1yekb8spGcroH2w3tR2AkyFGf/4UJoy3lUAo3HLBArOKg1zmlL02gVqsfKa3BZBXzTKAzmjHEP+
xruMIghtElrEG4302/AlqP+nxNx7WJvSaMsNTgfOnF/0yiQ0/J+rifelMSHcysMG4WurTZ2JpF1X
CFENF7495orBaCs2/yF4X0hAJKrdxucJsGTD1pVZi6OumLE4YTaUX8mAqcBI7DYSrEw9OvmQAATr
WH4/96kkCtXoMm1KPBsb9PudQNHihKT7DjiU6YbFBWUXriF+m0bQGISvQohJfTl6jJjARaM4sAJd
86ET+mg6ymIyj5OIcoKocsqgXfeQxiiTVqVPabuHp68K0Tuwhhah+D+wNSlO30Pkb+juHzIeKoj7
mb1wVHPc/fwP8gzjobU9v/Z2TLVkc5Dg0GOif3+8HH1PZRbyWAcItrXa79lUuJK28sGt3WBFUNkW
rwGXdpEp6qqZbvQn0AS+gyQyff7t3EAkHPWdggINWGzYo8SF375/LRGr3wSngIb0ldo+A4AqJL4G
C1WVps0TxDD7O9LDA5fjp9qct3flp2Drj3ACHAtzT9cA5jcnIoI0RsfEfi6eMBm6Kvh0qYGeMEix
FS3/pGoHhBvACk8kZXoaGVCRLUU6cIrsPljTlH9HL0UH6nh2EBaVNf8xqNufN6ODqARHUgx5nP+N
qH73C3cse+XciNAXPXPdt50OiXdPEIkw1wLoTMEkz+vuJLrqRzRcdixydCsav+iujPANEoIWla+M
pecuIxsjgubMrjiRwS3FXs2d6yFvZfMT6dyDwamPDEU97jeV4An8ET1NU5k3ytPwt0+6NwGxro5y
Dx6SpsWBuaAnjkwDhGpXkZS4vdh5Fc9U8OILT2JjHojHVpZt5ccUmQ+9bygQd+aoNEWou27cEMSw
0DIqiDQHN/izbvgckljhDrbu6p4iut2NXuPsAnTelBcRQw6oTqyaWWS/7RB0QhzEzXLHaXNve4zD
+rEVlfRiV7+Z0NO28NGvqTDFwAcayHkT+yZ3ACf5hIvKH9ZA4oqAUjZTC+qi2AblDY6Jc3TUfLi7
qb8+eaHb6EFUgkrrz1tPO9QAou3yYuG6zkP097YBIzA3QYSgJH7+FD4z1MAu0lfmq/mG2U2tIP5F
zIOFKpW/Ic+fnMAKBIWDpU8+cyvuvZBjkyxe02hGue86YW+3CPQhS9G5u59jPykdH0ZoVPNGdVfZ
0Y05cxFlquuDwupvMcTx3kdlvDK0h+mmuWu9MGMXwUQKuY3NnRSnKwsEEPzhmlhGF3nqF4ylW17Z
W3EBIYq6FCui3/RblSD3n1VlZMM8Uez8FfIv8SvX8zMCmg932vhm6IqtWpVv4ZUTRjneRVndSUi2
Ce0auk+L26eO8oRcxuGQPhZAyDEaSQ1aFQ4yxvmYPkoHAynbHh3EumKwqLHsfRYyUfOlxTbBm7aN
G9iKHK72HJgxMFCOfHlTEl6CcYCxy0hkDT02NQh67Y7PUXWGyqYxrvKIWQSVOBZ0lrN5IIInoLPL
tmIPxcwFfsVSD0pbI1BIGFvKbJ52XE9mM7VIqHlWfewFes2HbndiuGwi6rLDMS8l8zGRm04GzCfF
hDjZHX1N5jgEfkENywruzaJ5/mkTAslJN2Opx42jr6Ajkza2MWjSH04f7LM4F4fUHEkQ3eqOKiGE
zuPlz74IMR1823dDGotgAYF5R1uS0iXPXP8NUCOvd+LCq7wPZpknPeQH4mIHMEjaHfTB60zooSW9
2o3OwG2Lgwf4umHkzvpAvooQCtSDEJJFxsjsS/agxD3OcYXIAQi2sSFoeXHTUJm1r+fS6prqRZj7
r+W9whMk8YXn/qsAPKzCD4Q/9Og7iBXd0o2OZwF3gXzGOCDhgyHuLTSLiZ7V2l5LFfDy4rNgdv8P
dw1S/zUCmJhJ5t/N8UpycMegKQrhMHxIMMwZmDwNEO9fFEW3qMPbz6/tXQMIVxLbf9Pqmh8reD9a
ndr8Lu1DVvrfIw9MT5xp4D+pQZbBjy7MkMkRVHu3eJscOZRQ450k00uzKcHjKxRj8VjzLw52SooZ
VemDJ2FS5DZHHW1KpaJkjdGANXLEdx1Rnx+y33i8h446UVXTZGPHMnG0cysE6jS1nAFx/SEesPc9
+JVDTmTBKd1d/4L1OkyRHi9y0v013gbL7Ns58cw8Odf9u+Dik/U0WWCxp4eO1qQnQA0W5HcsFAtq
azDXdd67pxYWtzFlQe//yW7Mhw5IDGlv2ZBOUGfFAz+C62d/DHmDdWitSBXDfjzf+dSEDwGqYfu+
278ZEsq9YPiPPgJf+iMVi1zNZaeK6d/sZp4SO4++1RGAcqYbil2wsZW99fUByrh8QmgpcYWlMCta
vmPV+jko/F/Ovrtmik71CRyN1IemeoWpEZTpjm6viNcMW1hvtKygM4B9oDCAqMldnwJ7IzrdYkRo
9hhgIQCo7NwP4ERh6t1r58WdGCRkYM5UBiXOX2adAIr186eTiaFyaI7PgS9rd4ufQoQipRF+Y6fA
rpJNTr4Sttk9XzryNks6wyda8TcF/XY81OnJ3U7y8yhTgiUPai5AYT/K/hajfBJwJS6SKFLixSJH
W22FhKuPmwPAZdzQ3GdNMdgQeZ4HYnDO4VAPyMqtAK+mTVB1S6CC2VRuY82yTwu/pxN0iZqVsTkZ
bReh//BwPbVc+Xye3j5GQeChT0/J9UZluKfbrf7MnnilxtKCb7oQg9a9LqpkVy74ryD0pahbLF4I
vvCONCxjA9QVFsZ6R6MPi9gWOw8ZD9c9LAgw3R/1yMV/yDqcBJdMhew5AA/h2xLlLtrtMJ5OTpUD
9wUCnJR0eTPy4TKMFbk5JyXJ873GiUsmafQ5A5JvAcP0OQ+fyR78aRhnZm5xLDRXIqQFlV+Ng9EL
l+dyQW3w7S000dCU0PgmMH5tarNMxeDJOaftnAlRxxnMZsgd2hs6sunsFn3MJmT8pO2LUE78YMUB
+bqeYIFJlHBVarPbpzNtWWVq39l8+ZwTpD4JvJ/E+xPcHXWtHC+6+dubJfX7FM0mhl3RtymXg2cB
AYhWTlMNbvXKhUV3v4lwXxBVMsZsG2Vkh8jZH5oCacHT5iNxEMtEKIqN84LhgpVCxWY0F2QL2Nr/
wUIbxJoVo/4UBp+zau7qk7I9X/ch11dFPud/pyzB3N/rTuGIV3aoE55gzw4GCtxroYAUz9jUfNxV
TkFeUZ7sqoIirjkWdAUi6+vv0HYXInqru8Y/P4t65LVZ4Osr5LkmLVL0/nx6O6S25mHIb8njFWAV
SX0iOHwl6XPkUkHHc2eSkfDKLa/kfQoQ1X4coU+5A5nRC2J7Xb61wo4hbG5Bvk+YGOHKEcosgTVO
zGwjFGutiOwJ4z7fOsryXBf+PswcyxEYalhIx7Ea4vmENo53WDpmLNjA0JgodE7jnRRpK6QMYUW+
uYonB8D+XFYS6HgBudlTssJVq3F5NYub8S7dQD3KKsjsEFx8WbEaPkCrsVF3Uj6XBL+pOYEMXQYl
lPd0jU30O0vqXBOYrJ0ZHGA1qUy1asXJE6WQkEAUyQxBLDuorrRfXIU0oZtQS+cGzd4Dgc+2MXcC
KS4HcThCRm7uYX5fQf7iawDAiYu2ptX/PIw2S/88wwPbbRJLb1IGNrtAk9m5ubCBGB/obIr806sx
65QJFZSIw1bDeolCgueBSsnqasIMZZvFtguyS77MZAYv5JnOL6ohCTo40lV3e+qNtltCOWboVJGv
v+egic6BGU+j7Y676d74BBFCRzX8y9XpLu8OJnOGCAcRGye4VlR1D6n/JMTaT8BNhV2DglXsDh+Y
/P5v2oFQEv8QEOXNow03sGkUf9WHaxQTc6xe2t6ok8vpmed4A7sjQIdWIoAW/Lwg8rK2JhobIOyH
XocvEYLcpwLHwf2ItQ9T9qV/XsphlboeNmWhEyjYju03t1JzH9S1VDk8i2qtF0wam9KLBvA0Tfli
ygOifdNs3V2DmbYz0APbc3aN314/CbLF+FB5ickaptqGMJDq4MbP7ZQkB2et5icIhjWHE3hyPJr/
5ejhdL96SV2s9vHyIQf8kqMW5QY1cw/p2lnZrqgd9eBpi5HOzWcL+R3PnY/s7yP8gYsqxmZeo0Bx
HmDEjwYn8U5BytDlexyQNSphbNyjCuB+zhpFRJmn3/f+VALKqH4wzxYMEWAMc+o5K8DzhqIwXt5H
QKkh1dVqmSe7IBpc7emIrA1WVWmdG9sVcE847TCnCK7Dwj065ir0wxHjfmLOXad5mPHAyhor+XOO
POPh7A/pu4uaaTElTa6Tk8lLB8ZMKCD8xpiiHO7XJugW1cQzqtIEq2YoyIYYG7XVfVpNLaySF/tm
DmF3x68cYJzCR+3gs+8mV8je9/zojNXKq+Ne9Ut7EfDHyRZrWmc8AqDu5EqZfB33kOlfdWx56R5N
JP+VjGqlQ8VHD9jQf7BW1tFn4vPOV9/SUs+H6JSbhYcFAGjy0qQc0P2XKzWw90I2L8uq1nZVY7Cf
/xUg1a3J0k2oMwjCcw0wqySJrkFSwh6Gt3gxjSK+2K01dlhj1jgnblBn+wA6h+TqJfO6eU7IQdax
hGyvH6rcCxQnm+anaWFrA5+Nk6NLK0HqoE0d9Ol7BEauhi+w6vDhDBoroeruapO5jcD5tO0plfYk
veD1NJM/zJi/tgrHzvTy3+dYwvuQguUcPPYvMXgnnHB3zd32sTg+g8WD/jRjs9aXPTDYLhgFt1bN
gvBW4R7VTxwwuigq2bCkXY66mMmZjo4G1tblERJlvC8vXIrci2CwUmnU+rF0ohZrLHtB2BwHv210
G+yklsIPYq0CKQHByLFA+FTWdEIR6KEw+LvbykpbY/bizRvYF9cq1hcG+x2kbTrbcNsyRCM8WBAW
GxoZjCGd8A8S7327oNxiUPOcbdxRmUXrDJNt0btqFTXl95WglXSK+5pPDQg6pxznKDyd+by+Pta2
LBHQr5bLW03/htN54ZTJDBy2PkBNhz91+6bIATJWEHjfUS8PXFqLe0kMgX6moeC/vdYRssh+otGY
EadpfpIf/qvZC5osyo7i29AoEEAv/erNjdFfdSQ5wBMNETCsmaLofsiE/+U9xc1aQqcrfEnzqazK
CiCTskrBDIZn7M5ZcdIOG9Uifkkd9zhBOnL6HOc8BcKTcfLeXoNrC1SSBMG6VhuoH7O5BC6kMFQZ
JenXazO3CifoDib69yX913LvQ45ap6aHAkhp4uMIIm+VfdMDrLnqFqjdtkTlmdKjVjE8CCEn5ZyY
J6gDETzQTg7PJmRuBF9IRDdax1DdGgXvk+nFyPPayfhBHUBsMB0B9I7q0aPyQDhMjIF3p6Numnw/
o84GeHNqkutLo3MW9QMv+e/uY8KQOTn7JTFIYfcwenliO2bZUOAz/pw+y5NRLb2kDHQiD3J94VcC
bZdlh801DDysImCz9So1wEXXSRKxLY73NjXxfMtsPV4j4i0qSgJfK7MIrhVhN0uuCdMGg4j3V5Y2
/AzivOhmGMFwji+tfqGfqPi1eBvujLcbOUEJ6/yp/1E+SR5Qppv0Hu95l2r3Mscyt2KBOzhnhUgS
0lcKRWslg3caVTr3OjKnrCF3l1lsSa8nk1cHryn0JLbVfmvdAIQ7Bgulb/zTQB3RJT/pYavObMer
y50Nmy/XNZ2Jyjy2aTOqMyEntQTj74BRXQKxO2WTYSdj/WyTCPlR+2yMjAZxdfNCz5C6G9Klt2fW
prcCEbvjgiMWk8NTe+tBjg8YcETutrrPpTqNK+8hB5dD7uGJgXYPc+xg34czdKMNlPeVNM2vnd/5
L7RfuPHTn6loiof4QHDqJguBfAH9LX1dS6fzhjqOcc2pwk1yNdeXA0+P9x0v5jPckes3+pFGyz3v
qlCcflP7yyk8/QAs7rvBKe8RAP2g/JA5xAcJmJW6nkdbhwpf7QcDRjgdgCi+AsIWq77L50KTvi5E
etJbtFlrEfhbGige9O6Kzs16DOoktwjA8ym+kFxE5CkV4dCXUfbz1dnXXovINyVmx7KOL/cPrjPg
b617dk7SaSWh4Nr8mMVksLFABCiuG6cFPyoV3tYUG0+uum8seR0Vprgq637JaRMhirM4+oIL8JRn
0Di8Zh8eMXBeAiDllVreZs/g2BTkXzDfmh3lCGOyir46ZviDeZlbB7zzVYDkbPSRy0YFHio0CoV7
NjPJJXFpcA8NSDcRupwXioIS+Ufb0Sc76CE98F4PtlukXyv3z4HkpFwQYzK231NI8/s11iwla9ic
cyMlwUqhF6Fpe6goFYyHCl65bYh5CD3mOiahiFkprVM13yuukJl3cZKsvX0CLXkWcgHfkg+yLOSO
nWpK8K0qF8bgCoZI4h2irFSmkndoXcxFKKCNWbuhGnCRB4jItVQ14lweBEj1laevHNih6EVeLzz3
mwSowzDGhnq7AhCc9M41WxgE/9Cohyx2/eCWAzEbO/9Sl6v/zWQuJ/GQjzs6nDPnnxwGaQb4iC3C
kJVzYWTtljfo71GOv25siMNlAQtUng2MKIw7IEIaULRfkiBUnnFzcIm9x2smPJpw01ROC7hsfUrV
dLgCp0f+MpUTC84eR4egA107ksIVOzYVccT/rgleHVNN4TEOvwXhYMAyWYWBP8TJmVFcgUFWY/5n
hktzlC5kBNLPX7JqfMSF5YScZjKyP7KwBtK9bg5NjljGUIdkHQkehpgN9gmw0qNk8eyXUlxhND3k
AyRMhJ5/f7K5oDuXDGPxH21mOlYoNgIXyDxHWhYJnURSqa99nWQ2EqMY3uybmdPbLLAD7ozTFiaO
B+SQ84d+f8zO10XhJyLNmb1bEjy2H5G/1fqwvQGodmHe/Mu/m1GG8Q3Mg920Fn+oUz8IJiKP/H78
lmo35/ZX7yXEt0kkBxpQInvQWvE3mOjxoMGQwHRKvhPgfE6MS3erzFFSkgBSqi8mUMI4M0E/5GsU
amhM7D/BZViVOZCxSV7++Zl98tnRO6SbjoyIpwpCnvHAfRjZRWL9FVEKxGdSN9Cf0EmJJ9dgueqf
1J7IBLVhHfbhagv43zIP23LzmPyEUc1uGLPdZQ0b9b5GuulKPvcDkMSvZOmIR2hpmfXz62nD9YFP
Vtod26lLuNaOjUe8/O1IBTtflNjTW5HqW3gAlXZqeWus7ezu+sey3sGD9u0tPiWoHMDj9hHK5l1/
qTzZCLkqAO5m6N/ISPvjPpvkCqfkX2CLlAb++v3KWHghc86YjWaUSkAx69GdZI+PAfPqE/Yzjk/X
jUXzFiBzH9qzNc3w2l5gjABwvbvrAmPp11jtFIWZ1EXwTo1StRB0ORYq5lmDHZFs9n+y6G55/mv/
Aa3wHNRn+8aP9FdnSRe84KYolDZc43+DVPCUV+iNAWtVKJZS93LHgXEHtSLoJjNPJkrJ17B88+pX
7lZE7ecBqJErct9N+WgbBO/9f0QnHSDnl1HBPho8/i66OAgjwhFNWTHmcxW1iwR495bAY5e7YqK/
3FEbSg6f3o8pn7nW3nZxxn/7d0GMpCNbmDwIY6WlTDLiumhBf4mMGSYSqgRlrhRyPxoN7gxtnCTc
NXF8rN1WDeWc7B9fIrRAVQs0EUoh6SAFqU65fwyKJ3xxcVErtkOc3RvkjzQJkp1L1Y3AbHaJksYE
J7bhcHc6sYfxDOjFY/FdPraE+GXsJU4o2eG5hvHj3aXUCwTcVQtMeyODEE62mTGhCzv1eIrEIh+d
jz76ysBoK3pD4PxvQXoS4lXyQJyeznl+DWxkI8J64i+9pVUyDLksxtrEa3weEYC8DP68LGsDKf6J
CHUlf6JUkepU93eWGqmcTG1K/N1TdtlZRkCfuZZTIWKx5uzVnm6nHSREZCVwCgGIBWv6Bphev4W9
TZwObYhYdca2nFbn8YClauupNyDOE/pmrBY4G4zqOG8PLtydX9FlzF/u1iXd/z8CgIm9BXoTxzK3
zYqpAIoC5zJt9gKu6UBDC7MQnS6e0A4MHalHaOZDp5j43MeGAaPINtsxjXNK1RomkrUDD/NTMYxI
b2gxrgxCGwcYHWYOflUp86K8SCLLNj5qGJ1Qw+de1SGhDqUi9PHQ6EwJ+9XBZKkbz4+a5SKF4wk3
MM0ICuZZFXEEAHWWT/T9gwqEWFpp6ewbbxPC9Ii08H0vxaW0rHYRG/5Yq9FqM7WhtD53JhaarBnr
50vJypSCj2ou/B7B33jPvyE6gjZQxS1VYl18ciacPxpcDmZeBA4nWCF1/359JzajXZiPi1+TkLEB
FKHGfO/E6Ep6Z97xcNy8bZI4ioWfBNnTAKLNS6V14vC3YqTJmX4QK9lGzSkRbQcsPysovVJGtn4I
a1HPbrwHsTuYUT0uGFZUkf3bjrFckyXJfQrufQpLhdV3+PBsundvZ1BANcCE2V1KxKh5PSpQFCdC
roR9rnpS78nALwAzV5Yhqd4sdqoDIM+z5ERfzobx4dAYcBev0XVaC0j+hb8KcS9Iq0ptll8hOjKZ
6jSKVgL1ccF9zmQBNbtx9R65zFZkBRufTI9bDbEF/ETHn6+lJkoWHAtDw/p9SDoh9rSPJAR+aGRG
eVJZoniczOQVC/bPyqoPJDAh5B5lqXID16UA8c75Mzp7pkvL1WC2d+0SEnhqb19uq6vQeIcccG7A
G27jDjXwOgRL7WDjmNqxC2DlOkpu0DHx0aum1kp24ErU0yQcPOG1WONrEIJ4cdLhkb+u9WGT7hnw
0qx/Se9Z0j78ZmnKezgDO1yZLANEfLu4GhPExEKx6u6VyzoR5aUAJC+uPLYP2GJEAZDKSCj3XGmO
Ry3+bg7mgR+Hg2Ra4wRhVyZTweb/Q8Tw2UXVwDQrxzRHLgzw9k15WJrocHjyFOzBEBpkhEvRHmSo
LnmnAaxk6ogWiHMLvfiyWmTC9N9vMbIfVxfqpD2t9qw+Ehm5bVQaiEhc7IJHzAXqAwxSRdTa3HiI
g/hbkaWwY+fw3uAxbgfVa2vOMOfAYjV96m35a+I45Ieg3TJ73ZGOzS2/54NKdaPWwhftdMb7jzBk
RkLkLY37Cv4DwUDS8//nJu7B0e1KWp1Yvhvwn26DestvrnS9z8hEpVTaDUxrLJLRgbqemCAdqFIX
t6c4hIOWR7nnWg302g/MU6Nfl+7Fb4R1uZHcmKN2xYRCZ9K6J+erfB8yfW5zHWfHdft0YfF/ZciM
BbxKrlkCtnnqHOjgM8KyDOpxS0w+hgGcHW8SiLH2M7ot6Q+9lwcDyaVnMDJJQYQHbJhPJnpsNxSh
PrqcnRdetd4WIRX9+Tv1BQyBO63PdAWWJJuO2TdJQ2ZeKlz6SSCOsj9nNA/tJJC6V4xBzqjEPlOz
5cf3nepIKc9SAnqPOd8wGbImXQtarBHye5rOK+EnF0rXeqouErKMINQsvFa8mjXIgQd4AsNJW3Mt
JL/HDvGdt48HWwIgQSQwG/f9UYsBIWllieVYVbWUw4xnUKkT2V/1IIskVvcDIoYO7nNapjCnPCPG
o1Ggca1lPxqrYQU7XqskCSmFRPlhi1qbZvA+6fsnKH1NIAnxGkGbCPrEE+RiV9AKS29TzAdcDxF1
bpHOb9pSQYT7XxmFbZu5F6R81GdAT+FpPNXwODJlNtnPenkuqGRgmFGxmh+65X5kAvP5AR3MWxAo
CPbgILf4rSe6eH6REZjv1Rf3dfmBT2WAGMBxczmXlZvdZ++WFfiw9TSlvhlds136FQrARvSuR5bI
xhvTuagLx8BjszWasbigWNG38DoqwNcWZsLsOL0/3Y9wPzdYq0cOzS/Fr+rf8b5Isaj/SvfvoyAt
zT5X5kEcAOJpWYiDa2TAgOkLY3EhFkg0/mr+BQaUSCR1Ctgtv2Stav7biTPc5KQL8iamHJvODgA0
9D5u/7/nkq3JAeukTx1YLAYOkQG3/t/xfXNgNvLVhz4lqhhqp6kurlBdT7aFm6WRFynHipE/Dhfo
JSiNKyaGK0OtZIFcaYtTtXPiSD2agFH3qpgcG/es15fDZcUJ3As6T8FQnjNbDIFNU3od8rS8n7Oi
O7Uj/Oqhsqyt3CMCqYd3firX2JntksSGPje5lfpYhCU1aQyExo3Y6TbG55v4MMZ1hmqbWDsXawfk
9zIGKxAkK4kl1x75CxT1dqEctf5AzoxwkPN3QVua1FqEqQI5FykOP6jTvznegAR0p+R6Cdmn/mwC
qLGNS1HP7lTyX4ceBwrM0pEk5dFZefXXbJSB10FadkHMzcdUYduf0eWnKO4RlC18keZOjWX0GqFO
US6NbUEc9ImW1upojpXhK62HUm9Nnqh71jCGSAQHa7UxOLCCSxnZhsTQHp957/ELnGQOdK85n34N
AQU+E4CZFfwoh5aKpaWUFujqorsA1F4vZX5MiJ7L4suXMoSaMJcLnvRbIiT5qNz1BdoitWycgORM
DBh7E8kX+QSZWvq2gaUer7BgRqBVl11dxYdSm7+e6XH9HrwAvtiPbWtRLUWCbUPvrg12YIPaEv4O
SL++qLP1Xfg4UCniObVikBh4rgGgp+/owopAQCw4jR0wfJX+YyKlqWIa/5eDaUhXt7y6j3+0R+gw
1bMqFAw8K389dIBZ9hqPxsPIwT26lGkdsrkW02NK8eNwTYXARpsK39sYwgRwom7W4oI93GWPRyZA
x7tI56cTs6gS1+oZgqCwHhY3nTCw1YIQQirv+wscV2KIVA9XYfgQ6vHWNgcksJJ9AfZS6Oki4Ftg
dZNjh4PtOBGGHLqDqz+qlJo61ZZXx6w+Lfo73FZPILF8jEPhEDCMVPrwkWeTU3pAfP6Apy7oS8nQ
eNUr+xUZgrcVCItgXTHHbZJilm+Le9tMS+nuqRwnqnUzl2dxWB3a6ZViIgtTONNE14GV3pHWAo9w
2GrHrnGtf1+L5bQQQNzqyviYqfsrZAK5j4IAhgIJsily9Hav7bs9wlkEJ+Yg4qJkvW3JT2zOg/jn
+3C2ocOEBhs3TOzqvurhVlrCBPrzAcosK1kHcrPoOMGvw5AJesQFr10ZIm+NZGzkRtGPSRfbKc1S
Vs9/rlX13l6pP9KsxGaqPWNKWVH0mwLknWSqSO8RaZ0g/41Y/Quu69NBDAFb8fj2yz5xUOSsyDuD
EqPwW/2G8/njbCzzrBoRiYSPHo8V3hQaF0jZ8UePdt/K8jyvoM7cHy/ug0X5wahbwK7t4n7WOMYr
OgB1vQYc/qS6NugmCc9b2ono6u46r4CNhnnWNxx7TzhxHxGiM5pdEmr/2VZULd4VbQbC54Hbqe2r
NIhDEjZYFxCD+QBFxbvIB58huC7vTqUUq74A6qRk/44qhl022VbH1q+7jtjvtl9MtFd4/cUW6fMV
da/HuVZk9kpMK2kIZm8Yw4wifSX8pwF8JPmonY7W8OLhsqySViM2dgb6NLFNWr3WakHYen3LlxpJ
FGAh1esMDXlRrmgHm3AFchrliqvWo2APkCFWyjID20PsgrcXfEEj4FJray9anlp8OacLM2BDtg2n
066FPz8OfQnIRc9Rhz5cUfDRfYUCMTFTy/Kxq0mF3wxk4n8wYNdNO4fpobma+yBX7qjKr473c6s9
qmiHjpvHOUfiXb6pgo5ml41hAcK3O7fBUqvfRQG0/MY200L4T/lKpyPrXs7tg8obqR0G/qiV2MnA
ZLOajtayswuBd03YvQiZKQ3lcWs9r3Zr12VwSx5kfdn0TQw4umKjO1tErYDmK/T99MIOrAiBlKeS
JEm7zmvZlIOgZFKtx7J0p1HW1K31eMFh7ZemWWiioWbeUC+eoy1c0PPoWPoqGzqJHDWkWmUrp//8
MULoUvonVtbyJuigjX6O1+Xp4XE+oyg9LVDgd8+Y3axUz7yh93N/E5pGvxrC723DFIENmn9ueZKk
UAR4DSFvVwyWxA5zOG/MM9iKeRzDKpKO3qKuHLFTl9qjm8y/jH5eePsXQcct8AYrVnUL6uoBGRBg
xguSCllkfS6trnLp/V0ytkJBd46wOAIlB875nGLiJLVSwqvlZ1gLKH/bVfV1TcAQu+M1Nf+Hp0u/
NDhzf+Ln2TCMOH92Bjomsv2A4bXv7E/TnYCsRh39jaN/5RiVdXe4Yhy4Z58dBOV7F3BOiRHx5Ev5
6TItcTbFwPP7vFktnuUNHIQ/9fS3DXXcA4R1yswG2pHXRWN7EAQhoRNIhT40ml6JjxZqc7DXvugr
IEy855mSvxLgLWoO7bH7vOFiAbAPPutRO4qVQ2PkWknUCVwvWTVtpDLCOjFVe+tuYWoVVMvExMY9
GJXyP5a4e1JszHotAQ2IFZtAdby+vbY7HwH+ATSOUOe971GEcGWB0MmtHtvuh2pr5dzvfcqa0RHk
AjTLnB8JN1bWQbteC0MPwqCWH4nSadgDQuSECttKULhrhZAPjX4MCwfwQVi8cyjUfXfPb/MjU/5Y
5Mr6r42E7aLt83hwJ7yyWxCAXf/W86sdkHr55rK0RkPZ7WNWZ2M+gjAbB+8/rRrci7YnxgvQPRyL
ITJ6T7e5AJps3nLkPPGkq6zAB+H1Rmf1/ZUx/pYzB05R6Ydcm2IMibJ9qxhH0jCcMgn6GyY/dODx
favV56Q7ZwA5A/KsMwfmSBXCo4neQM1JTlZbExy3nJV6A+AiuYJr2SlgMB3p+FACDKhaHiGHaURS
bG4U8NPvJr4nhnq0Owe6jlpSqXAiwcj62pZ9mOYUeVBIgvmDSxCAlnnvkmQME5Ka3LIrl1IFSImp
VjpgPtswXx/nVbIab44dOZHKNeNHpp+iuwNMP+o+VmWIAi9LX0Nwg6szbXL/pwIPZquM96VCjVAr
1NKTNZzQeCmgDNj9e4sEgfHbZuQUA7UIFZdXAfIw0BRp2i/GKCR1Tee4+alz/arWhYMXtJQ7e/hR
m4o60VC8/Glq4BTHtPbkji0ffytXIPdptwFBSvxwPiA/hVyj6G0IUT4SZtdUfs/6V58YecetOngG
UjpNHGE5bPdA1XTyrjenxLAJtQe9Xrec7dlvv67UK/YgROqpDlXgZNSQvq82EkJIpgCwKBXPE42Y
aKKF+6wO7ONAk2LzF03SAvF/K3LJMndiC9u6Mlw/AzWlxgNT+66v3y5jWYuHYDPxhJXbVO7fpeCz
Op7R8BR7a/jOzEIFXf8FWA9NS7eKdisyq+4tFQr5gOJiDrLfjkQ3OHT7ckcLzQMb1/MxT4UrxJeW
BD97Yvjsq0R7HvhyzxkcLvJcZWhGOx+BkscCojKJCILP3x74ugVSsNVnaZ16DHLg0AczM2N/MaEt
PTRl2NxgSYwua5d3j/M0olHigUGHK7Wm3RxeBRoPDEjDtJqWJSs/UekGVdosCVGHPnDIPg8sc13v
1hXo8qOzrcQd/CmcyKtyPbwawqk9PBUmDsH2rhd5ttjW9dtqJgp1L9ylwH7Q+/M06ZjNm2oHqtIx
WYAbiXb6KUy+Np92vXJ3Ml37IGuO1weYnG9kGdXQXQHBcDbQcKtN9Lo6JAARWzvbFi31q0OBgeZf
qSjJ+l9p5KjIUOq7qK+k8mIDzJSO/2j+7p5MSJk/+R5WEsv+jyVoWn/+VQPRfjGou0OpXfrCfTf9
rH1qfNxxLXxg4mYQjgxoOFjITaMmcokqUd0R6/8DXueHJmrp/ViSnyInX+s713cOztJYc59Hljor
qitRVeRIwBgTmQkO7NCzMUOVXk9c+XSLJ1hNU3KuOmncYhSwLLx8DA50t/GGRRe1XsoMh4GjyNQ0
7Qq9ZydEjO3zX5vul2oGnO5wq9KgNj1ZDQlCSnUlJpIuPZuRAVHHgFCNBVluDHaQFM48Yte+AQhC
FOn6VLtreaDw/yL1/szaXgoloJ9e2+hskOVv1AaugD/xzSWE4u8os17/EZIai8dtKzQIXZFiOEMg
I7CiX5iJu2SjA5Ubo+xBlXjHEe2Bo3E1ox9jVq1xlhGu7FaalivBwrWvgQRlcVODexotbU6EP05z
Fvrw5bqXB97ZFrXh5QL52yJGItPr+6oXavkQjqQHCrxODok8PvRoTGgn5DDNzYGPl3H1R1VP+FNj
k8LcSym79pXkPwod7HJ0SOH3uWXWRow9a3XQgQKz8OH7qTasEuxVGqXl0/FD91movFo8fs+rs9A8
oLLUUwHlkyn8PUdtzOwWQNQfvxfrwAf7OzTk+40ekb6KY2j0vjb796fQJ1/PSsHd0Y9xJ2l0pgam
qyTx89SSUU18y32EWlPmQRBSZm7f5rzY9Ymq6NRSx0VddKg+3OokhvoK+QVKPKfabh03jwLdMDAM
rCDWjhiSSeGY0+H9dMRsxQe/l0bUgG4adJsfNSTHGQ0Gyk7KhHHxpBSBiLUIu8qIAw071wKYbDQL
KTcVNQewMILH+ukaoRAasuyY+GS39LQBe1rrpTzdVH3OmOoP2wjBXqAfe2bdONZypJRBtYxy0SIz
gC8lImg/BjrEKEna0kNmsjFtf8n/zB7ypNbk26ESNbwiRyx6eUTgXCyAY4iw6mIjNHx/8RPUWIjt
69IMpGTwdrMM/RJmfJ2GgNjLDUgl7gF99ZoFoT9yTm/nPGC+tS/VMfV725nOCcLJyeCNykZefwzt
bajaeVFtEElZkNqsax+IN7x8X1HFsK3ych4fpRDvTFUS9WsGgrE50SjCxQHR+6/VYCGx32H79D0T
tiuObGQ3/V4Xoif0vuRGMQW/tmlQMZPYKDqK3cYhHUIf/EI1lRbxRQ4lfFoOQQM14aYnmWOQ+NF0
Kup6FdeKzc/e4Pm/athYCwxtr+cBzI6jk4kj8SzqDzlex+S1Ym1E6AjFEE1diWlPxLT24DgwsA/I
fVayUxGeA1mY8Yo0BjEU/4p2vpQzITotcySoRxLlK5Z4msWdNreXs5MN+euSGIJ7q51l7fNKnP8Z
2FU9ehorPYS23NldF7YMtIC8JGcLFuml5M+yZm8DfFYzSfLJ9PB5M69XUFP384AViYD0FL2MFqEt
DjXwp27vPYXne2LBYeb3UrZac+xlIvAIK17D5xiORFr0xRMaR8h1ro5fyCpztDNJyOvndRJe6c+i
Lj86Mw3fJ4a2g9Wk9E43dYpD7PJwD+Lc80sDEltFGJC/IvxEJes4sGh6zRW+ivGAQV5uzcCtE2Fe
BCKfChrL1e3aTqQrbS5t2CVIZoymhVqq389FXScKDjpA1/l4ll/zGpfZeykP+L5WjO+EMXCOvMBV
LKIcgBejhisHhpTq3tmzeJBF1xHh7F65b9dyzA+70NA7EFAtOKEknY0dR3kcsFlGBnuwr/GpjKKv
BjFC/OGJN0Hp2XwoC+AjSGiEYZ5dPIuVv4P7tp2ytgRcd169CCc72l6068912wMIPsC3ZlZsJGGB
3rThTxHgLrhuu0YMNTGdhPHkVGOAQS8+qLKnlOhmt3v9NDH7UFwN8W0G/gOXMjLWu9VXvf5KSHN5
69i0GT01EjsOcHovtPS/WnyawZsI5ZPtM4m2eDfC4h5cjgOh6SdIbN3h+kTE3PncedslrWmL5lS8
GqTABnsynzRfeFu5xhUr+bqnRGI7ncJyDXjlGghcnWNoXEw4mIx0cTKCY3XlkDJkUnTUZTblxp4x
8viDP7nKe6HiRInPvPocFUAtKadocohCaZ4sT5fZCtewKGlnQs4gFciTNTByhjmpjZPCNH9xBvm4
9ivRxyX4ywhodYobYxsYhbZ0nmhwOjrPHzxPPNPhnjzI0WitCUhyzoXehazBjSbrgp7lmZzFy98J
uXj3tdBOZrwwXGtUGwj7wlAUmGy++NRlK122sT/tYnmm5K/zN0UXy2v1ZZdyb67H9z+C0qsAzHc1
59Y6ELu3lEhT8t8AocwrDkM1dgcVJGgV42UkAA+DHrlRYZf6IXBxY8a/z+pGzRKZUiKuIvANdoJo
8vL1YcmNae2x9AaeqrbLtNzN89NGi3rMircTo2+qeNVR0pMZBB46AMl7lFKiY8b1xU1zw+h/iZgp
FUECOHIfpNsDtdx6j6eVO+icW3gjlMgFRdR5ThB+S+MKQ4ESD6Gu2z0k376gK3NdPHTpLaBmDBp2
UOqdxgKNVo4oX2O8Pr73Du7++qDOC09fgxMTVvKbcDz85TcRaHP0Z+tAqj2UuYKHZLwWj0gIJjQU
eQeTy24f/Zdy6FbxOEQmZOMyImZgQU/XaOpqaCprS9+0vXR95gD8QxyHw064uEu2pVCfBWwjZUdq
n+cjggSpvP+Uxkjth6LkdHeYwHWkdOoHwc2VqQa0r/QbIO4po2POD7azDxQSqjrgCs1NuOS+VLTW
zg5j4GHgIwMG7fTZrRSHMerNqJKSki0RqKDwKKgNiHP3jQd3ofo/3Pj4Vt6R5FJz+kcqPRlWlH/K
jUUFnGf64s5Vs4y32j915hkJRv1Ceh4Ad06VPoiGFP8/nj1taYeF45d4z7ReU3xpNF6X+vqMG/mP
lon3Lv1zLetGXaVW+P/KF8dGq5TWJy1tNO15It0oAefMEoKYF0Xp3qcF+MrSXvEsaN6+f3ToFkaR
apeXpfa+1iBzaRPILE8ZpWf8S57ZujTSjNKS9A70BDfxff4umqSFF0pR1F1cWpavwv729249lUQW
89ayZSPm14J2KwU3TI8QYkBn7ETX3BXbCnLKIQ9uUPWC0CC2+o9q5hXtyO4LJK/HYF08f5nGIcjl
L3MTHuUA1hT0SVRP9oLl740lQDKkhX8DLC41J8Xrhmf06AQ6TWqwuAuOg+CD9pDTbCf4EOrdM0vk
T/qhN1nRi8tf0630q0iNgglKX64lUWFCygJx00Bn/y7xUmgZoOKho0gJCt6OSCDXLG8kPrJ8KFsL
znAd3C8tGdt+6plxCp2X/0eKsTZLJnfFCirzlAaLMCKtyVxtiwUt4MoI6FlNvUI02/L0jJBpfg7y
V8yGxqUzGbQ0gdpxJ34i5tu0M9Fiv6On6XZevw/42uul2xfC+/fYMA2aYMlin+zr69ge2ogdoadF
cbaxM2tabAZwWIkSsAvnWZpJRyWCCwXGuksdgCF5j3GbWiRoLvga3fJDdxD3NsSIoUeFblSm3E4f
kEKOjAT3aYrfvGO1OzhZAY1ZGIj9ZsJjCZlP/xEhhMrQn4h9hMxKP1rIqyQTJuCKigwhoFc43nou
t+Vs5/BoZOmfwVYYmqY1konojCK0mrarBYfd0JUL9ACibymk4+3RW/YLCk9fH1lsWJ2NYnZ0ezIl
igOvpcg4h5aMQhusQCRIM9fsoN7DJj0HKNKiLVkZD9Was0HezVQRjs7P4JU+tQchcGZEULrewCwg
k7MWZUg2afm8AJ/bEN3ohF49FxSa26M+hDO/aItdSga2UemKlmlZ9C54eY+9G5PXNGPwWq4gpKLe
2B/oTSr1FLV3yZz+Q4G4EBaIkLrtnx38FTWSS1rzHWAqV9gy2Smz9pct6MoO5r7NxKTjfQ4NmPxG
EEOS56ey5/6h2ophTwoZ035YfnNsINOfQaP3sueTz3BuXoYPTrOFfoc79gf8YGcAP+QBrX2rrj44
eKu3At1D4Fqaldf0/cbuzM1A14FfQjW9xggxyofueMs6eVdTc4w2+qV+Q6i9f1uF8YbGoVkeTN64
ievHiZVqI6KsUms+XlHwIFxtJDh98J6/RRlI55JKUfdbwC3uU6lVaLHijOHZTAj+oQSXoGdv4VVj
YG3hZHsbDZ439pkbx8x1yXoeyRWDP+/+FO0K4dWp/7d5PxrELwWKwsiiKUyK1FtxtIKXLYdv7Am+
sD1Klvf0hgDmAaPR0PKL4bPyO+FvNRW0JzBQ+JufQMbt1pEFnBCfeL1Ix0tFcwrcir/xABE4nQ0m
lXJCEaMp6bXbR1tuQC5XHaHc4f+4cy/HiYxbANmgu1A7aeOPrk67fsbeTWsSWEPMY7QUcBykTLpK
H8GF/m4Cba37WmKpxsF/PnoCupGhVYr5mI0QoWALah2cNirZG7bhD4q8RoPb4I0A6J1YQ8s7x3B8
9cwxpRstP94gfqveY1XDccVBIvHD7r5atpaX/mIH5X+Y3xl3b2BS1MvpnEWhOgRmv131Ym1L29wc
Fbf4dypbBx2JrCbi2HbkhDsBfikFR1xUKPKV2TfBfDNTlheEkc4D9A79/7mzZRraa48gm3V6I4XI
Xj8/WfdVJD5EX3rdXLl38DXKSkWKR89e4mpA7sZLXr/BhU33qAgqvgcoB/B0/h3HoneuLWyYSykx
9c6OACIyDJhdGTjFtSz2rZFyvWuQiPQu4Xiv8p9pSPlMdQ8LBBLUwe1RAsNM2FN9mzJNiKuPcnpO
HduLvuFb1x4ASgCdECX0jcVzL1k7+7EaiGROCWLaAFFSj5jd+vcagCVLa3wO/JymexlRKM50vc4w
6uHn6FHqY7uZ73qplW1VYxixMQiLYYC44v4gAF9Og7DGY548RmGOyP/kD/XdiNmvXplF1BVc3VSK
r13Ml4n1pMvZ1Sv/7JhZ/svRVOvheF9+DYNQzod1ZWGlQKSC1Gf9o0AOuK1QBSkH7tseiYg+1VGv
HBElyoLxL3cEtM+Gh4EqcturLXIDY0m5noGAtmPA1UQLX4JsEYvZa7Kgd4d0VXEEm2CCjGZiCMHc
nqLXhwphL7wQRjDd43doMCDbrBR2JkEznCdN4X4eRhZ2rAwAzO9DQYX0VnVd8fkKfysY+TMJWwqT
WJzURd2anr7Qog65xAsFEALtzBAswRuwbIRCtohiQYRZ++86ddYJs5CGMRYKACoTa2gDClr8joju
YLVM903czl5Q1R7671Y6rmgeo2HB4Oo+mO9xNEdfIcwE5zeJadNepplZtcBmPzGML+7vVVKrt+9g
i7CwGwkr1iptVBnHXch/XZoxEEdgTDy5PpQF18KYmip+vNN0XObi87WKVRjGsL8zt+t5taBJ8yI4
+/0U/V1Ex7/mBgiToXdkFqHKEv6HUKOQPTEFEeI5/qJg7vQwFEcLB3nIKMlSTe7MB7yi4yQKcdOB
q2tBmtwiR6n0k4JIQmDgbgg+dJn1ATlBcPwappkmllWPqSzy40BJOhzAzGDKmiue8iKpK3PcN24C
gGodPTQE4nevlUJym1y8AILaWi4cP6FP3rNum+65wOW9mLB7nno7UURGLhr2YUwt2xt6P3ztasdU
rG4v4rTMebyUm8eAEp39UiX1DEipM7vb0eE7xd/MqBY0ivjwVoZlSmNfkWmDTPq2LWHG6gCaxRuJ
y4xNwe1jfOtzMgSmttsZPBvzjaA2QayJOk2B16hYkgbBmS+4SbfRW2QkpCX5EE4JZug/5WW/EuzN
kLP8xjsyx0XAulC/tcL0wzk75c+iNwqeDUgCSUXR7BrkLoPSM30/jKLcG6royc2B7T2lL3bhOG51
1tAmovSOpq/iRERW/5RwAoEd5bnB1jKH7jYBS4FYrgkV9umdt+dYiyyKRLVO4AwRehcu1DL7Ru1o
RNSgH1iJKDWy/Dkp1cjBflT7xX4aWdXbGsSUGpSewAPpHyG/XQtyty2hm7DZ28oEAtm8F7gfx/eh
JLA9WDPRmU3ntann3KLwLkiYgzuNp46pOcJQX6388iPooAso/NWHqVdDc27qK5mY7NKWfeIZCkdx
tXRotXusxk8VJqXnppaPByMAwmb7aY8LdBaMuJGbhYDtSxAJzcELnEkUTyBPSJGIQeIvxbjNkaWi
ZD7/RR4FvtzXV11XQ9/Q+7nsd8sD1NeuQMYto5+kGidA1tfcPhi/kfz9Eu2D8ot7CjuZ3nSXcrq0
Wogz0Ik4qUDrvnFKfx2BKGaeZMvt2hyj7+RKDUvtsifa53xGLdE1mU6yplvavJ8lQi327f2s8GZr
WEnjUhN7kMDKcIvuvauAoJKHcVC6NRxumAdDzcPUJg+LJtEt8cXvQ/UNMeeY8IOZtBFhzHmQSioZ
/bpW9NAt6dqNxwcN6xMYraFcRia9nQOVytyUcheimql4dUnmbn74NswnUZd9xBkhigN9NjOGvoOy
AYpVF2p/DYKMdbMKE6aQXTJCJSoV8cdX6cI/H/ahos+OsG9l0tYERUVNTDX/VxILufYzX9gfQ0wY
i7xfBh6DCgsBl8mRRwTznqZ1vXH1YWK368uv4Yx8u4H+A/hzKTYjyj4V44Ni/6palG+pzKeyPutU
5zHHDk1xuy5sJ0EicUTFmJZ3XYfzCNd6HOlNF/CSq5IVVNqyNJZzwqQ6DE8kNZzSOWbP2dsUfD5V
WtJciu/qbOAkJKBo2EWeBTmAob/YFjDfWyuuoGDiyErn2N2tHAKShSvkBfhogU+tlJw2YGj1vmc9
3udM0pp0zYWVaM+PZd+U2+fUWycX3k0u1rfTnY0Rxb02XFfg29TTZWw18iVmcBP5OVyrtVDyjzv9
ajJZe0RD34iV/Rz9FmT6aUI0w9kqALS5lD/EXkV9Q+pR+yNv3CqfcmuhMmQsK6n/epOPOrs8xp3q
x0Sldj+AHJ4YIa39czq5MuZQGIhcwwG0u9jntLlfOlbfm/oBmfRog04KwCbRsrQVrIrEC3l3j0YV
fBUYPBfVp6vTWoFjuczLq1N7dNsVVtEFDkMGz5WcqqgzJE+8kZe5VvPwwQBq9KhbaCxVnXp6jKj8
AgHVSAKlKtgw2plxyzK75DwtSoqL8gLiERqFxthYz7chx8OjKYOOavhuz3LD+VrZ7tXV5rWA2YAl
1PYzDKVJbpfSLdfEL/ckcYIgGKky6YN/zTX5x5vSIeu3TYpbMjBFtxJAgtxttP+QPN5mmDHIG5NJ
RPEwlQe/Qp6Ux9NoI7rhmXysWi6nrJwftM/ZiZxEzNPj1MkuFbQ04DdmbgbBuX25Sb32tT4hqdy8
EB0OhLGIypVyttTKK972olGYCVE13h8ZLcr/B3SNFxAQB7nkr6CJ3x0Wxkf6MtJOiYTS/7Ee4jLj
L76CgIAZLZRtTBkUHSMc5T9hiqWhzHQCBzVnFyNYV68Ht4Hk+3Wdli+p9pvSrAN8t9U97tHICaU4
Y2u26q2hrzaAxZY0npTO/2vfJcSKuQQ6efC0shTF+2lLfBWPWTRtb2nWAEdHnPpPnzI8MsdqmzSw
EwxwbY9hcn3ZeRPXRWi52hWNgN9xSeqrmZiUjZv4JuHipiMgQXIQCNKdzQkxgccJFVUzT9njmlEf
ZEl6+FeDf4px514dGyUjSOFWR91V50ZSgttTU4CJX+9Ot+FkbIqYpPgRcqHadW0zA/Wach3yNZdf
9IKVLb23+OlhkksBw4yC9lv9QlLyyTQT5K/e4XAsR0h0t+xsB2ragxjf3YjIjLaigz217c0/k57R
l8DAfy+b14kinCO0akeTheeH9+Imez4ZWGCNoO+Nr5Gn3nFnFR89lTWCsjNvmh+cRrlYCcwTeIrC
0i075jj66OF168zBgcxqmFigcpi41y4t3yajMfVZLmO57wmfIy7EJ6qEihrhvl96SrzTwKFYcUe2
dsVpRwXya6SRu7Ys4iI6VDZ66uYCxjjZ/4QgB1sQmZ29gnkxebcmfZcmG9vZ1jYsoJ3qMVIr/RTN
FgUEVt4oAwNi4stc8dwNRVT+fl/VSkGWqSeMu7sS9WA/UZ7Oc8tjnjjrJgNzIEZqpNi4hQayDlBy
/hiGX847HB7XYlVr2N080q1b3uSZ9PNjuWNTvHa+kiTtdTjkNUzQElRnCoPbJ9M4F5JLRcR3IOsq
PBIFtjjc0FMWcznZp1qUkxf3/phWYq16dqY2WT0mOhXdiLn+6X4UBHz8l0vKxAu/gcqi0dud+5zX
8/1p8PPvw6vGDANQJMhkcoRV1Dl87RkR6+bKvnWf1QkLRsRMf6Aceiv7qmDXPaVzy4YgI6LVoGVH
ABdY3I3K3ZAGN3i9NXSwZHFBJPZ2P0ZmSjtj0dcAkOmRRwwpPuE07qZftJHj80BW0K3whQqNWMWV
A60oMbB2huF/lr7z8qLP9F3O8gXunBbrXsu9ISG1N/vyTwd+6kTtzWNJPU0rzSN7HS7q0CYlLLYr
PbmpCSLIGWiHhOXqPTJ+oYrPUhD/j1XHQ1unqedUY0Sbo6ZH7nBT9SYLh78xskx7twXklcIZd6SK
xltzCvjsYq7DCjROhwSQAqSQfzBSv0eoI9oST1hKXIXwcunhKvZwva/dD80gDYFj3QJkj617AM8A
8eigrcv1IWv6WK3ZR5l43kNJuhDBei9bF97iOpwGpRvs9/rzMepaaxOFIBSxDG1jgKgwe27p7BaV
k0/04aKiUAY7xbL0eLiPbo+8fSPQROaQJp05Dkf5MQxmO1a8X0/WweMe1nVWRK2lzFJdqUoJBtzj
M2j8z0Hd0Ze7YN0GSNY6aNDTia16YTZ2BpMYd3V0HPic1bqb7oCcpDlk1LhXCTLNDpOXaWCckIA1
nJusOlbjZ3vWzw7ex73GNHeBltmGmdNIzQvPlx8BWO1y2d2e2Nbfd4TUr3lfJphc8rv+vbj8yBvA
7gk+rtD5i07pQRVu84LbF4Gqw6P7sSH8Y4nlK+UtLBokcWhkwJ6+YziwXblW3WI2iVFE7T3qufeN
IIQ7oKDdH/+pjvOpzX/3G2sBBe2uOPuK/nefG3qNFioBUphhpL9atijNlWq72mbqZsNV0z4KrG2M
3nW5rSDZc/H82XiAbfMkw7Synm9b+XAZJTK5qHentQegYLjXgr3gs2g0ZGuTvnIFXM9T/fZpDZBu
3M2/gmf3sMszFIM02iejrBfcGug+xNIZBvhu4A3TfdeOl0Yb9tkNM8Vr6f3ciAReba4zbD0LZgg/
5LKJSW0pHsVYLsaixdEqFQ7gc5dHsVl8bFgXxNroYXI8qF5/p9bvQpfTyDCUW3Of3/Y5O9CdjRpp
kUVIa2yk7JPlf5ILyW5YlfOC43dMBK96D2eC6uCCAgr9Dphj6p6PQ4cu2EYYVpChzmXtPkhR29Fw
o/eFqI2zs0kNFeF6iVmuk6+e1yc61X0h8Q4r4LZu0g5Xd2o75peIecM5wYDs3szn0loKKtZTHlHK
tUT2xdn5iLvjhnQFd/siBt9WEYBqZMXcJl1xpT1AHcJZKOz7IkLHYSyzvJmzF+YZCCwMr3xvGmBS
l1CGe/4HzQZbNbLcy1sbZu+8h3fniqDc2I/4hAKmzdGtgx9zEC9vnBjveK4+hxDPTNaPHDmcS39h
zakCMdNV0ERcifp3GUMJDIIPdo8N3XUZeRIN0YW8Rz6uimZV8AmhkgxNajAFKrmAACKtOtbW6rNu
6KNmPCNbPtqJdqm0nj4TodlEK3kZRkH5hPIuOo98peyDEgON+yfKitzMYy7ptvoM8p4Rcw92rxgV
Y4N6Nr0RuUZQMnAr5ewE01RRh6PHcw5IsUdeqk3nfxqlG04ZNxiWgpELXDJxSCApd5TtHCWrSYDm
2Qr7M81ZwuhLlYdpA3ESQ+d7D8qL74HqvWvvnAZQqCI4m0t+7naUny93zA8LKRwIOXCqC8jsi9Pu
bqs65FqWG2Ab/W/scQWqXh2v69wGx75EOM2FxGULzpqZRAf6X4v4y1GsMhrdM1XCeDs6Hn3FGW0h
j247Si0G5QKm6eH9dygNEYiWp+nPCBsXQ1x2oBVWd823nzyYYEkApogQgM186pQvgneugHUFQmDV
vdNjCmtsdQQu8EhkSdRj0c0YEPaB2D9OXHFto5zvRbdeZxGlieTZabV3btspdLsiaLQHT/CNuKKA
uL6JMaz3MwQFcdllZvqsbqkCXyPLSSf8HaV3f96OZZQm4EnjwbwzY0phMD3qptlk1yaIWHS6TwIc
EUYlWhS3FB5kLXH5LocD2+bamdCiiVFB2cvc6HWZNOjvw4bbG2f4F1W0WZQpxIfRa2Y5CG8KeRtf
IGJXpmLF/21dtEBO90/BxVBdP5DzJYVDuhAC0F2UcqHqoJScDu4RhSBsD6ilDLOeJccqFW/USnxQ
vDHzZ8eI1ztXrygZdXntAXtnee6bfD6rwlmyzJKScn1DagHMZ3QBdAQWZ8NbmtmJ9uoSO+wEDNYE
BmNKS7+VWxLQOzCEuJJP9Gmsk9YdRy0NshMYdzpc9u8Cs85bY76RFxjyEW4e4txX+pDc6hnYHz9d
QNoUH6tBCFSpmCBtKY2Q9zKTpRdvrM/NcGULZ2oQqvqRzZ2SUZebpp4IkyVrNykp2C/pw81U6+WN
A7+gvKp3tcKsylZXwaTpZaPSFm7w7ze2GyzfZMj2WxhNssGxt5IYpuwMaFUi/OvH+wyPVQtg+8+p
MjGyjK/7wWxo46fUO9hOj1V031BVAEApSopSri01i/hlMqz31kY+Ghub2y6pftwD5/PjVHJCqq/e
nyIooqTHdeCUKy3WHTDTaR+3uNICyVMuuiLuKWPdzkxc16K1FXCXa4mtkPi+eQ6X4lVH+aIZ3/1U
BBPAzmQC/wmfENTG/To0uZhaZ1wOtE6+96MFwlFR/DjHG9UetBJRPjL1vS+JzVUcygErEUl/hqQ0
Ft++uM65HMreN2HY6KVPAzd0AfTiD4M6vu1o2gEbPTWnobnF9bAYa/m3v1Ykykoqk+eJ0QuIPA7z
soNZ5s9qFzR/ocxPUy0JsMdT29rpP4D8PhHx4EbsQOydcGsoEWQGafzOCKjEaWg3qIG2TWuaMgZI
59ufWutH5KxeODFUv+7cebCpi+tMtAfQ814N05Uczz6AamiGM8z5ni+I+SW7TD5QgFAV9k3Qbw2X
3N4fB4yINHVSEYdD+GtNjABqTJwpzQAh2W8XnCR8WoRHkZW3Yd9mQNfNiOEMrLjobYvisHVqV2Kf
BPVbFnx7TGVwwJocpI+Sf78LTGoqyb9ijWDqsn1Lkw6My6sr7E9lYrB77mVo1jBQlVqCqV8IN66f
E/MHoTLZFkSNZ+lHB3+F4gZEvlYDOzLX7OrN5hwapdJYiMSfIsjWdpci4EW9mUa4w2r8IILYvdtr
dEEEmFNiC6Gid+BXVwPC6cYYCwSBGVAX9DYhX2QGTE8FON5ueA7S3jQq5QF6yvDz9i5iRw1D92WM
rz91uXT3HnwxZSHpS3P17auzHw2pXdGTa4OPCzZ3Zzh6dXNwIjBrYl/i5Koav84p0DaXOjhSiktf
C/lHtAaS1muCiHtudfqZU6SXCMPDJreVzw+qt+8fEi9TOfElQT5KAPj3rDLIAIYmHTcMHaC878he
s31TVchw1PKG1OShO6L5/WxgmDTw7fupCfZadabfS5jcNMrolkUIcclQl6wc3zOjS8PaaV9bkdZ2
a8ZRloat5oIbAo/15HUCNIJZn2BWk8HTeunzgHByPAPd+9ZB1xzL+ROd1Li/W++DF2XGCXb0tT3P
1OBj3dKCqEWHVhhRP/a8xm9IQs/gMm83wfKVrIn/FnYgX/vLjyEKxrtFi4fU6MXhiKuaRIYfWMMR
isf9DnMs8c4o99IiDY3BCztKwUZ+lnWt9ejIy3QJIw1fxZ/MVZJccoS2cT5tKakbYnD+HxD7JM0C
9ypRDQHsOygijTWu7eYLX39v+bgl1rzgmYwG4LoAdgdh9nRgjFJyJp9PH3oSX2po3vzg1zFukbD8
LSLX5DJI2EAFFDvh84q2m8SuMvAsnjDGxXLShpqFLn8YKYALgYWPGkdLlTU3tc7X5+QuxO1y+TeO
+ktRwa3ZxT92tfaM1fq342hcDIYzHQfemx4Bj6Xsf1di2/74DVeHqOp3zEQPIb2CDG7J7QSKYt0c
sQ0pcEZASsQleDDL8qOra2fI93ojTAWGhs/U9hZurF6Y/3XdIeSJyPdzTfxgviybCLMtkzxyKRo6
R+IH4K4/qZMJCq8/TufiwQZg/Gbk26uN66yORxLMYzCLt3Nkw79c36DlBQQtFsu2RbpTzlUGgjrl
c4nCN1TYMb89QlVVdoHnwCB1HZqbbF7/s5JglftSf0TX2IKla7H5zJ63u1uVe7mPIFBwlUA2ACwk
EEA1uiJAndcC05pjvNWVZQw3qXHcpXcLF5QghFxtFbmJOD/7nokNqWSkyNtU+bq47g6o4evk5ct+
d4mEfqIFSvGWxDCa0f2+7R8Sgdfd9U6ZatdA34Mg6E1CKILdQbgbgcFmRUwbSO+6JLGs27o2CWnz
nxjBgkx9Ssa2nZA0y92lZsVN2l+tyCMBW0ruY+9Y07vjmeH5QWJQpVSOqodzElROfI4HTssh7AtP
kJYdAU3+5tMIKxMLInEDRkxjVRbzcfRp3QFAQGIdLon3HCwxwYCgTWWfVPpx4Tj4YEKhAIxh075a
ksrIP+7sFJjB/KTcPgbCH1S92CUE71XNKhgUAslE/Q2gaVrXtnwqdtr04YrQdj3JNZJre1PWLfVu
P/lg5ylL3SHDPh2/H0T+0DC5Rq0/9NucZcEDnbQRzvD+m+y8SN32ZZhOgGao2FgJAvMw+PDvoMuB
jYS+ISaDV+PtsrFx2jK1qFCjfFvCgs55J5URcMOykTBMiCJrnMUeWOvHAFwtW/GsyPXaEBtOcxXN
ExqScXIsWJMdcPYbTo80sQzQ0SHLa3Xon1qRjIMo5buCe1uAsNlMbjiwbSppD8iWzjzE8cu8AVnr
ihQQt/39wy1TYySsRg+h+VSvLw0VRcY52/ycAjalWIRLmyLIvcMu8GVl2pk8MneJbb666p4E+f7O
+lXd4eVD9xvpumBokG+hoxly7DLwGHbateWjWA9Tn7PJcRDaKoLJpVDhExJJA/6gNMe46s35+rl+
bzj1ApWGyn79f0mhPE7Sx8jtraNpHPLFzTD4cXZhxMEgPHxLOJrHpVGUZ2d5s4FI3FQRO0HBfF/7
09XTEQ+Vdmy67t1h58B+hOnpy1dy7GzZ/RRpumh3SgZ1pDbszWRhsclck+OpNSvyWNLNYZOBYAKo
X6N7/i3VT0DvyIhXhc9jnRzByT2u98+BjKuxBOPBMJLhtuse48GdRGmKloeMFxWMBW2wvVofTKMu
ClbQ33bNHggF0mmR6Jf2u2U2v7fSmMIYw2ItyZn/YBUvEevu1cfwjJgYQW+wBrb8gMspEl5E4rej
qGXIuuGG1SlF6TyOkGMOGfEP2NXslPz6Jfj85R2YelYS3vU6Cew+Is45CK8IrUrgseKqx7n1ozJk
Oj87ioW4+Fkoh0ty9GuT/xOs+QJ7BVXf2eN3BL8z7/2k8Kh8w4VyHiui6SvA0oHLoWMP5VqeCcBt
DZkFOMF6Gkp8uyGsc8yC5j9rcmx+gVq59C7qSYOJaJpnT8rzMRkwdmM7Lcw4RdTV7aSpcrMNqGyp
aF38f780bj98pTFWuSju4JGi/cEn9fA3H7R28kRmNW21KMai6Se7xXGSlwtSWEWrUHG0kmFE8IuV
bYFULEuM+v+0vDEUtp0MJqu6tfpDRSCjX+Rn2+3dxROwCHZOAUTh8ca9kcwbovdn1o2jEFTxlh12
WcervzzfdHuVDby4Uofz99wL+e02aUS0lN4aOIT+VoqqIlAStd8p0330VjyHVN6B7LxyM5Xcd8h5
umlVdP+Az+GTUDBEoBQDO+/CQk05G6q0MOCujShli3b2YGhWQTbGTAlVAdGgFCvXaHaG8oXJjrJq
nTp14bvXINY1rN5AcPmwuBCS7XowE4+X6MDYN7IGf4A1w02MskdSqykO9TuU148ZQrBn/6xccBwS
RInDB4/KL2l1P47lhVkSFMzY33/UoJWSnLiX+mySw0tSCL+1i34WnP0K15wwXeNSyQhQdNAVDsAg
AmZoHKOF+17GVilNO4a/rkxO9AYtMxYYpqRGIjbvjO9kBSiQL9KRp0pB+c4eATixbxBptGIDRT/2
9rEp960v67aCeuYRweLqtXAGVV9kCCQY9cgSFbc4EpvwBSRSZRSeH56BT53amOvsspDHnLzJ1LSZ
LRQ8x3wZdAhSxWcaZnYHe8pHRaP9B21/Z/f3HXXZmPE9oFtLUC+ZuiX3psj9HvfUTO07gYjcxQrF
AzftKMQkcAp9/3lO34EFhsvZvzS34odG0Ig2r9aVCeFqYDBqzLbZX7aOO0CUewgXT/pxS+SjQQpO
83AzzblWcqdM16e8hATdFp7E9TGTEHVQaw3T0c0dKDOOjI95kawXA3zQF5VZobsy8nvuemMvJPLU
tDqZPLak5eQL3xwogIrJJrnmS8Q/+KPljA9af/pi53JX/rAeTCXXuvfT61FpJQGwsFnTEJrZZdym
TbuxfywQsbB5/HB2/gD4Ic0H401cfRKpN9pSvBegBLX3KzjEYaiOgMmC3JNPj2f0Sc0Euc1AijJO
i55qwe4qXES2w05MlWlPRq+RH9Gbo3aOKgnX/qI+wfeFKcQwWTzcCm7yTw2QMjTIP6dHFhS9bUIG
OiVEQLbaV/eX3D33/oY8uhLknm4hdIeA9hBDeyyYo8QARYTwycVSvz6lTWkYDYlCuC8bxiOcA7B7
ylycRah58B8ZMm/tiLYDzS/qKre1kJa9i6u8wD9p680GOp3yAg/wDELmKqorIS5TrZ/XvR42Spgl
bmS1swbDOmPeDeiDOtNMRg9j25JDC3v6nzLQQmp6SuBVP/V5RXcTx0qlIJt2dcXku4LrzEbRzoQg
/q8WImViKOC7m24OqF1X3+mGfc/xWd5VBbcvVTQBf+nZbMKODcQDnhn5kqxEq5CQvXALfbXKYRKy
THH/8dgkqg2cQYEgHlkefX181a6j5exdaj8us06jRS6ayYnqVRGhECoVMaw4BH9ZB1QmTlSwTzzN
OzNf8gwzc0AjDx68gqgAm7+V31yh82c0jdvxaCpUkalgeT+gGOGBrYoRL2ex0ydAkAToshGx5p5n
Cx3MX5nqAFSQhKs5Yevc9tIDcYhEp83kf4GQvMXfi2n9oVzU6vRazLqmbeKpFNuNQQSaC0sq57Sh
Dlp7WoFvuZuwT1lAMxeNObNsELkjeRnTUZdtrEaH1pKlZFnKdvDlb0z8g+XYo7coGq5dSLG5OiYn
0RwSGQ9vpFlhthR5duI9FKdQmTZV8jB9zR7IjNv5Ol+XAauZHX62vZ+9FO7Mc98Jy0TtQ8rMCl07
ojSbVbWcbGuEU8iM5gj4iuNwmLdR2JlbwZz7h01EYdzwIA9tLK2zm6mUQwpM6E81I3w6vrW3eXIk
plwwNRUlGldtcknjbzqfNw0LAzWynTLfMLBDjbk33ZYnXNVVhVtBlRiU9PFrBRNHgdx7Ktb8m8pX
jKMNOCzc9UqDGx9DWhqCmlO9RGT3JBUFHOAmRJaLN3uJYKV30WOEQ5kdTJcNpkgaTbfpF1cQvsd7
zUNw5Ck/35SX9I9ZKI7NxwY63KVkumif/WhRcK8L4Q/QAMhdOgl3K7xSLdz0lDDDLteFb7Mn+Ylm
QFYOjxngDJXN7DxUVAAvqI4naOqHpTEv1QnN7dREgd/1wRTk4OqXBgRGCwlqTh4DEugZtxC1sE1h
MRa8hGxZMscDUQop4raehMu/FMkgYU4tVrNnD/IbNDn8mKlNmj5QsVLXhqsn2upJfKHvQXaYLFiX
aanaH9DpClT26nCaAZ6fypN5OVTpzYblNA1YvTZY65zidkajGvdtiPirUDHWacrl5EEUT5Vqqzdv
zZfylz3/yvR4VVffyWw/L5M1cNofIXjm4fSMtsnolWQs4QdyUUJa1/gIhpeRVwpjEWvTxaFA/jPn
88lJi30GK9JGWuUzMeu4BRXXlTJ6EngQR7+Qy/hebtvV1wNplRkLpPOcg/P8pyZOtDDIc3J2eH+u
a/PwUeXrzv33PgF87sJlaiQFTCe6wmg2QC3QUnXEq/UuMITfI/XDCGDkuG85Prk+J1fYCKgESzCJ
3Jam/sTzr41RBb7CXwBuCruQydzK3R9Q628Ks+DXJuI78OrFRW1lHa6ZrLDXNkUQbR6zH3ZKk1H/
0R2mJRRggf9XyRrBI3v79hMR/JcDmzbq7i7xfnw2E1nJCCMJN7sLRU6d3uMSvQ2s7KPNkLYaOb8D
a7sXlLdimNnOg4zXgV4g2OjdPv/zsB2kkH2cO9oYPE15M8t+lIOhgBVXpZHemaE6h4cpQXrKUpvb
V9wd/bHTddVkV6/sQoj8KyACAgiALaDlKJJ+ZL9JuDvY+F+F3PBUqoI65IOwM/oFIZ84nxkYFMUA
EsF0gHc/g0ohHn/zHPmFbHF8YeuCox4y22XlgZZuTRw2agpRxBQINjtV3CYqA14RMwo9ZAoBGyX5
F+khibLqJYEMnkftGAShBs9c/Hcy7E06i7/zl7C1Drh/iT31litOT8OWpQKYvD2yKXw6H4YpnkGm
yOwYhssk0nF+13C4BHYdlEXl0Jpt/5Eotcn4nRv6qsRcGXPXhwVuyRn4MnT/7reJ4IyLh7x+USB+
8l+B3Tu/rEBwQWXtJljmdXpNyGZYoyQeQqQiw2HbAet20V7tFNE9wC+F0UQJNDmVQtCZR1wnLuBq
5CrE+cd0QRjbVLwVj8C20tYcpnodU6oniD2g8PHN9bBt0WGcKkJ4h2rOSkdG9MgJgR01uuZ+aoDt
+K5c+wAIiHjdYQLSqIVpzZJDbaXl9P/qUSdCcVMG/fSfgqm7EDFYhS/jEJ3UMoi3d8EMco0Cw0bw
L9RXUrefCdHsiAqWA/6uNZKZF7xRy2mlGbtfI2cE2HCv8sjnLiWnWvW12MYsW7EfBDXR32hMTnvJ
byNI2muH5FRm3TzQWDtUKOw0BNZB7bbDGl+RyWzmjIQEWxrukwYwTXsWloSQh9+h1bu0ztgyi2Uu
cLDHNdL2jtffenxXIXGYip5MPWH0vuznLipklAyPejEho6iRTXj9kxD9UDrGHnLULwdqaG+dsGVP
RHED74d2QGQKjg59GeRBIyZ+gDbUN0YymDRoRfvdaFt7kk4xIRKOzB4VtXWXBkPbbtporF9NQ3nb
eRyjmOmcXdMf/QOyg54TDAZxvu0AHKTwZNCoy4SDaGCpRMkDo9phg4+EpEf5Uec+1M1BnVx0vnbA
sbGGCtr1Rtrhj+kNu3ssf7WkgA4N03IrGNXsWq59pYQKvKFuKzrvm6ktt1NdBDyOGvo51sHINygP
obCROEx+/HCQY1vNbWx0bkGOgmBvhpw9mmsmlCvoiBq4XrQJl73SIfZVWiyi682GScki7YltHbCP
mMW4KpiwJAiMI2L07XQRlB1GRCCrNdOhFxNHXiUIPmV4O5tLQwTLy4L59nfMXrAkJTEgrory2Q6I
UdzUhIQ/+jcGUFYuTcS7YFlwF4Q89B1t+draYt7TUcR585y8ktw49n0xP6+M1oJbEq/bfXumAUxz
4Pg1tU8P24QJOk9huE4VInu6qywOdQpEY1/SVsS/GS/kkqsXQ9nRFjQfKFSaJfVDmMOcJeIst0As
CSEQHjxKTuqRL5UPEIFyhFZubE98SN1+Vs0Lp7IgTKhCZSArhmwbCJP50zD3nlLFqH/NToleNlxg
dWfn9MYc0t2xLlazXOjKjMTiYD6+bhLeI+vL4ZDMAgAnq4hVWUR3wg5BHUXZi6QRPZwSlZV4yawf
RXehyOuDF40Mn7gVqU1z8J3wCakH9lgURJJv1Mtq/4v7BzjIytTEfXy9823iE6H7IOGDwxWRfduI
3C5AD6XqlXTBWQfDAA871+ybOlzAbAJVpKl1p0KXq0QHXoBUiMf0ck8qNuO8e2Fs+LIm+StqYHZP
jtZTS97fmARPt9wiJfhXAmmSNm7SjCMfXXaOd1dkIEz3v0S1jq8v7vt8IHKeRZt9jznBs2nzoy4C
Hog3qet6KHQIrDfbB+llT75R/6GEHFgUHn6JAqLIP9Jty4QEBudfj3n8HschQCG+Zlqy/N3YZ76u
ShsirxhFCwNZ/44EzgIotst1MvpcnprewPrAzu1atKq8J7f1n6Fubm9BGSzC741irMaOpcE+BWmY
eeAD5JalG2MZmA8KBEtF1uGRQRTjPcKhWhSFx5QU9WYrIs/YRGaCdPb1VoAGpHp9xsxjSSt/iTMF
nFDAX70Nu0327iKiZPCL9rh0gYbU9UhZ8mSCjEPP12K6r2DZg7Bywt8iQ9Ma79vIG0G4gKrkPS3S
P1btzNBShaTyAW4sOleFtqF/gNGssEf/DmyTD6KqHHy8TcF6zE7o3KWu8rXToaTy8+/gFxSqCso5
4rCP/KoIiloVVvyzOH9mm41s5yRRphic4+ZSJ4tJKZW407wLFS0a+JKYug/Zv20WQEET4FO3rE0R
QlGg7S4aDTWw2m7Pvqqb9v3mILdTAjgvs2t6pYldcqaTB1YE70a+dV3vYhsSqL1DTrMw4ny3Oz6k
GHHRuZ1zDd9tLeE6W6qS6pYyuv87UaSMbqh1H+aLSN54yJ4fED8waP9N60vj86PrlufMwvzt2sE7
T+EMXyr7YqqEFk8FL95qVic3l0Pnu4bWSAUdML1bbPAcC8a+7/jKUb8P7j4JkrjdjIE/LatkrdRt
Gaj/H2tZPhx1m88SfdnY9cb/EhCMxK2gbxkb5kd8tLl0PuXmjXD2iq+YXGjrSXp3ETb4DZv4svYB
Pv0YLiHmJ8u/fKkZX6iYc79uR3aDoiNwBdKJ8B/LBi83zs1tmu43+RFZLshr5sJ1E5Y4KgDVta3B
IgZ9M1CiS1vbb6v4XvtF5YgP7SkufYHrPVnKZyQwylLpCTZ3LFD1OwDXXBl9BmMZk2HouLhSp7F0
r4f+xA6aaLuyFI1+Y+dJOwb9YNvBn06gWk/8uTu55669dF/VlHyYPEFf8stQ77m5ElpChVNpRn3y
KlGl1/gT6+oPhKjpONFy34L+hLPcz2hmGC6mN8LZtSqDeo+c/VN0Ob+AfCAeOCWiFQgnW0aHd94c
AOzcphn19I45ncWxv3ExIZ5xDT/cUoLwFbxR2//yajY9esJJ7JikDq2N6u6aREj6eBGBSuDkkT0O
PhDTBJ7LuVRFZmzgY2rim6zcvLHDhxD0k+vF/lfZhp1YUKyqW8JcQAKXnKnODBQ7nPzoweFRkXL8
NdaKJ0GgKN3uX0PJz/4rCTRkju1tEd/bXVF2Ry8zfQtKX5zsDT6EmbUT2dM7OK6PVXGjr5YL5Lwl
9InzkDqvUAFLZNsYnTfexTOx7LkuYpoH9o+rZNCSJdRPOMFRM0U7ih6iBunmJdO8lFx1WJO+Iead
VZaGx29y6Dz4Uf66vovl/mUAdB9XyTM3e+/Sd4/6AwJ1LY606xRfWmfZujVy0nerRZuKNj0Hv1vk
ig8nm5C6yughRNyGhuI01dACfj3AC91kuF93S20HWST+htrrjuTgY5yHNjD3HpP8JOu3BnnpR83Q
NjqsHLm9cM6dfHQxR9tHJoLmGxg8ipzoNoc17juefyrVYmna45rtOjDYjFKAXYRvoKv+k4rx3nmW
g22JhM/db6ircE+XJlfVl/+O4iud1Sn/Vnv51V1uJOWNrZBDwYs+0ktnPYJYI2JEUgoHyyjCarxK
rSoALUnrfT3BUyotsVzBySAjhbjGvTyTpF1AZiX2K+u5YiKqhtkdONH0/JFIB2eoWZ7qXkdTRIDm
9z5SS2/cTmsu1DoiaIN8dhDD0J3QhgzzS9v5SYa3apqiGyZ2q6DjcyqCXTv3JJ60Z69rg7EAVOND
JO74M/7wC15OQnUWt23PZ42wbyfFy1iNy+JTTzTl84vBVSq1TvrTe/v53SbZbkOSUBDbhavIa5TO
TzXmpPAexBPqAp+09LvO2NooR7/pJSSJkNtBuygOv6yQrdoRnAyiQ709UPmznH+/dpxFtEGTDlOY
tAj9GBzx8IVFfkzXv7QYAy1rESvgj76U/g3GzX6bpIE0aBmqLleINeXzKX4lIKz+cxaBL8M3UHHy
CH1SPZkeC3TmTZKJvyLWDJY+mc5VZXlZ0HNWd8o4TIHI5E/EFQTfdI09Uz75OW8Eovi40x97zMDk
ol58/DNM515v6XffpT+/vJv8P4oASVW6zso2ogJXzL75W/Od0xzZLnaoDxw0nTfcNA+GOi8nkJrj
Lq05F6W+TjLcS7frjZMx2c0KhkYoXbJu3tVizX2MkFbZ+bIDyap2iSOMYeMww0/W9ncGB4v+JwJR
uqfPlHtg163wn6BOFe+zIMPt68bU6HRehKFWTcdFQeas9IsaAGz+0FePFub1ZSKLyrds8aF4xTZR
3e2lB/M5Oujr/rQrP73hx2YY10O/VOXSjGZa/z7Xa2wM+iKxFrYypG9/nY+064KcQhkKkArOX1WP
eUPABcS8OTG/ZoD281Dxb0sdDmXrKccIssa5h2D/TVJEskYYvQkZiGrJGGGbNvaudZk8F+E=
`protect end_protected
