`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6256)
`protect data_block
KqW9pfxrIDJpH0Oj71uQFWrisXRDIY7Y13o96we9//2H1cpYueRtk/std5JRUtEug6+TNBgWpAn6
mw6FVxIwYLWbhE05voxeM0A61Nuuf/CtlfP7eNlQHPFWUb04KUNW1a7B4xBqiBHah8BGzzjQVFlq
ImAJsJhc/TqKl0LIA9pgggozs6sKgc6jTcQN2Qc8xJbONLfoP0OKyi/jo3nUVB1AtZ4tdeTbetME
+F20/Hx1N793rtOhbx+/VWwXSOGZXRSvRnfDCXuNr034s2D8kye2T3UDsiIE4/aJGTgiDG7L/wWx
DB7NpkIFBnmgp8Rvp/XzcUMSIyGOJd48BYf4VfPoITud21/L7a6aGq+NR9jF2emHAZMqBS0QX9et
oknB+04SPiG5C3QUW+1SmrOf4oQx9yWsDOf3YLbxz3Mkj2kgfteSkSUuQ+Fo8k2Y6JmLGka6FaYu
+5mzOPcjb8+iMe2WNTEcxkaruJ3jo7yTk4mSVUOKL8fb5fKGGQsi9KEBvYoCH4oGwRIDkYyXgG/P
Sv47wIB+qsYgx1927IbrbTRsLFJI41taQMsjws3Ba3PAyBQUKWdrw3jJrwRlnZSnDURHAuVv9uKA
qhFtKqS9r7gT1+HyFE+TroO+PJstMAFKJf3/GlYkWj9CX7xwfK2RnTetRHQsgk+q/RkgZdtAhrpO
k+m5zxKAIcaWd0hB/QAt0yEUgn+CZbzq3t8WYkkpeAPvPuKSVhhk7/HVo42cjeEWq0J2g8kSNCNp
N1TCVwplJUjD84F0C1HuM+lA5vW6qorvX7LjBhbTwPWI4op/iEOkK2kSf3NJxi2vDAZ4YHdsNJvH
KO5HLqk0SBH8CZqVMGUfmqh6hmHbq7D0uq2Zag1dxZd5gshFJTYf36Oz/gShjb1nZ2G9lpJ+5fW5
MfySylmJQzpYM66VMx1rBvK8kH807n5XuTssojj+Lbo/g5/xtji7MIBgBOvmno4WLKDvlYdNGz+l
YMgvFpPZGtlcmugBdXZCI2P3MDb+z5W0aM2v7tkBBYuDDZ7p+aDqwbQ6gC/UQ1VPeXhC4n5VEjC4
Ozv6OZ5uk9rNvl7soiKyhH0DVXDE3NhATjqWIc1clOc8tKvYINPvWfeYHqIYMSGLmPJ5OY4d7fOO
E3R/c8xH/5b8FfS6sFSDs1A0OjkW2JUvntzTnRcX423eaFseAtXsmYk4tjVEX4LQBeyPLA1o9d+h
bGXb94dFBUqFbTQ6tAh0ZiBds/RU7/3yGbuuwcld32JhRPJC9SBvJ85SWpmxkFovn4p1DdekMhT2
Tihzyj/HhFErQAF++dXbo6AJlLvnQ0m6E84loEa0ZXiF1QEQfOJdW7YEV7eXqVR5mxnROnAoR5p8
ozu8Xhn11yc3p3dQw3NDc4Dg42oTQ/ClV/6cTulGp0VZq9BUVrNpRDg4/PouwrRnEfaRdqWzkqBl
3kDD+Jq3Lk9t6RjdXs5J0OSlgGG95bsQePXz5TDPx1HVOEjJKM7c4OWlXOeOal6p65X5LvlXABN/
ZsT7D9GiiH9TGorMB3bPuYenSRQR5y4RKwjUKDyCEuTWll0R45F/NsFKha6ssSDDJCQEz+Cqd45c
SqysAcloLG1sgJMHewNrKL5b2dj/iOIp3aKNVeKj2fXRqomvGCzr9iGMXgLRxR/+qj+JXn3cCkY9
Y2FOxzeuIVAOOwQNGiSy6VkZ+RGuklxmf6E61yBI1T//LdcvuHvJysICTQ7jKz5acQLELtRQisp8
f/JkOE0nzwdUO64MnZxWVD4AfcMn+rALoJ4+YPbexh8Wbt3MLxKDYheP+RcY3cVZtwy83jx5NQrD
OzxbEVm3i6TUzil/KjbE6P9kHSZJUbOZ2CY7QFYAmdMSIfzUA725pjnRLq7m11zoTfY/m3rQIaaX
NgxlUmOUEMNg5M5F66XQpHAi5dllubc+CCat73ZB+Qqqe0CbLOZtOo2rl/AfNcVymQWvOdj+XLAb
3r+7kDEJIiM/OcELU2hx6mLFv7vqjkWogSY0oryQ5oNDrTG7Vi+RKDBu2oiyEGv0YJCdNdzTGmk7
zXCDZC2oJQQf4iaFLpySTNlRuNb/2U7okDeiBWu1PGKogse0B3rJB6beCHUEOeUo2LBwQLB5hwOa
8R5tSVQl7tiFoh6ezncGReJUHTROumypEKuJMh6M0AfyGnNxIjUG+6n0Es51WGxKtBlEI0LhDi+G
4HVkvx3dhFAURStFF6w5ZDqU6ZlDVxo9D4xeWl04X378yQWMLkOpEmk6Iz2Bq6wlRi2kVSl1XnCL
o+WMhCdFhsBecciIp/vw+7uhVv3/HclxcQNofJgFsxSnp9mP4hFaFoKk79om7VO0eG7gifKheKU5
fYGayZsGOFjJYqAPuonEvZSRxQOYpSHlT7GmVC1mmnUB1/aZ2qkFc2nzwkSsE+LSEDyn9FNVZfsp
A1FN7v277k0GOTCjlS9vlbo509fHW68JdwGKLTsPZpCN9z4/xomHIzcCQ+5Su2XdjtAdIoq4ZYJ9
7U/nhXEu5YanXC9LydRwQjvi/sThcASGi2jQ1+90CXMaZTOxCeMuOWWreozYwTENdNzHSRv6bouD
tUdTI3SqeAFA66pjDGjXTiqheqqT/Y5G+tZTGIuvnVJsZ1hQH+pPaLGv7yJn4Fo+9vA/8XxI9OBK
RUvIlGpaKXO9AJdL5XXvvvKF8KvQYSG7rYsH1mn8gmRX9TOXsNXOpzPKNCJ5VmLEvOd9V9UX/X9c
zU4AOPLIZ6EL/4NBgQrg30AvCA7DevbXsQwxMFHZ6U4DprEWNzSwmBGbqWAgzW40pNT+cUKDkFOH
73jOIxy6M5cxLhT+1iCqeN/1Zo+VHv3uMgp2chEnkOijcuFk4SyG9QmWIszfI7y7Z62iO6Wv3cdA
kvU/VBpBjSufxm1z9YQZErGTz+DiiVETSFPZ0UFm9hc0s00MIEHmvrQ8kbyynDX/Vda/Ss8dpryC
BF/6/iJdT6cM+U5z4Rxy1cRrnS2WeKAoCvnBPdjSG2PW1wjOMwie6jVfrVNKLSXDAT/s2o9XNBOy
95vY/pS6YxX8beP3zHBB7LX06mVlBk8J8gsDcbteP7MAVWgaUguVc+BYzssgW2h69WYvhEsvA+cD
6ogEw7YH5iZRMHih29t3yvqiE4S032ftBxvfV/h0/u7MZ98Xefx4auuAugGVslIA3CY2jSLRKGK1
hbF3oJysLn0OHEfBU7fNghrKCQJF036usTvK8gGCSaIEhD9KVg5V9z6QI9jS+l2KN47eDRA8RR0m
Ty/gNBXvEEBfNgTmXbxsIYWKPq2ICUj0zKa8GNX7vwAYB8jGQxWQH3J/Lq3x4fjzFoHcPkKKou8J
CzWs7VbCqGLt6TMWZNjMF79FgRega8gUGhDszwAWjh8yWktDHfm+9zpdP3amsL6Vk636sXKVecEf
kXbJwX2QFdLwFk8OM2jG6WoOByqJdE/yGS/M0gvsD0YztV2PZbIp/E9x/PY3A2Jj+3EAUZdhyuIT
GH4F2EgZIYt8IoTGTLtHBRHb3iYVsbfPCvb9PguwRk+xKYWLET/1hdcL+hGu8aRLp4SAsK4BMidg
O/rzmutT4NC9b+cYSC6EJgEZ7hd2hL7qXMMn1ILPJ80nar3x9EawjAZ2MA4YGXll1MXBXr2NYFBD
JrWBogDIzYx2++O35b9T5i4vfV3mUmqK7C4BM32XPa+r+L9ZTH9izx0TzVDeDTUve95iqQNjY8tz
JEWnkPZnfXxPJv09FuQ3sE8Moa6FbgMMUGUFc6XotIlyH3PLpIrIpIVNHuGs0l9nVD0z9wKxAsOl
5031rY2W41Eb5V3NaQxlzVwF6J0ABfTWbf6DHugDcB/zpIy1yy2kZ4M+u6Ob8h01sd9s1CIvldyx
NwFYBBkrRaVfSOpSjPFB3kFTITynEMjIBvK6n5jUmKm4p0Ic+z03yCWVXGYcylO9nIqx6juwbE/j
ilTlN7hJ4WcYCz6OVJPD+sQPBiGo1FFqTBmi8jZ8BuFYgj/bH8f8G96pRrGeSqkGvNPSVzm/vkJ0
7EN5r4cBnteoIwSuso1i9MpvJUS70ty2hC8YSxVQVDK7BIG222R7EgR1hfn+ouX7cf5pEoGR6zdR
/S2HLKH45uCqakSXZXLfIbbSGDlTfa0aqUkd6dXQLCPRMwV6JFojHAaXgM1cVxNnZp6G94bXVR0G
5e/PmDNUWbqwH/2KSHwHGP0MuV5oj4unbIBgmVJJcX74dGfTRUmcHWOe85EkO6yLnq6rLcm5geCW
qYG2i81q7q2oY1pZ7S7qgUOOrqRrUYrhPcCYuxKh6kwjaJMqEbztOhSz8kkiYFqd/wfq3gzulws6
2MaNxr2Kky86sPbT06dOWrzW3WaCCgr/TuLzyZLTnGCerw1hhqOdTx67NhwnykA43JaP8aO1tU7+
fqC+SOOw8uUiE911+AljSHQZfglUCm/OM/LD01Negpwcomz4sbw+zuNJfvgciuDLB9AqmatEOHSG
rs/4m7EHqwODb32tLpc9g4cNOmqcIYAv3h7iSmYmjyl0W0JlEfOfyDIZvtvt+8SI6YVYF6eld3D0
w0zbCKZ9LNYrOWMKtz8h1VKRJwwuvkFyLNiO7lmHwy5C2Y28AoP4f6oMkHWze8ssHqKMgnG+G3sx
Xma5auDQEtqKbweJL6OD9xnUR4V9/PR04ld3QR6mUmHJjQbHcchkgwiP3tz8Iun5Ltqmq4m8r8Yi
yKFhWHles7Jq025FbLWIULCK0UZ2vHvUve9cqvCTiCFBNcy796+pNXHWVDPRoHYaug7+dsQH3Cn4
9Y3mOh+lUb8jARe8goIwDQSTJ/SSi8l8SiRXTrhCmn2elTk5CXaHv47Gt1A4wMVZBvxoYEf3tJhm
w7qtS1OwgeyqAEnROj39qiGQ0x1kAl4TN09Oeq02mCQbskMzpU/LYUPCVJ5Jp17Vmc09fAu3Lhtd
Miz/7it+qHhs8B0HH1IijVJR/cP9OTZkRms+ZklAuL9cFf2lJrE32yoZcT6VV79XU/VPsQNTpftv
J7wpOl/Jmed2ys2Qrxovyq6XqQhEs6vL7uGviUE6Ls4+3IRZa8eCV11anGPppU9tlxPGPH+zL+Kc
CpyfxYu2ThnUyzb1I5ViC/zECh1ZxcCQluZoHnvVCHiHnMb/uHtjiNk4aOsZR1mGlWGmjuFL/GZv
cUAY0aj6AQkvljWpP3kC+MPidcCZD83sfKQC25LzaMrxsatIfTH5oLOhPE77w1kqUWulx06Da5qu
4zOdx2+mgLibPHbTGdsb2zrCNKUrXo7jPkPsd0PGcefvVqARoHf8a81r3+sNi3lhVV1IF9xzFok2
7ECDTJFLO8xn5YZ8bcWvF6KpBt0U2l0o+6kUvDmpf0Qj2VhUBhFQL5gJIiwU5GYyRo+JW4V5Qyag
esnC++e/r0iZq8Bhy9p8viVA8sUvOzk4p5HXHoC4Sj2K8H+4l3lYuYDVZ/tjrGK6Pmpw9cRSBqnM
suZFCwN9uD3trahrMrPEhHcDmcEbdT8XVaFQtqIKhy61Ev/8flvmn81CJS2T51adwdtYPVDTmmCr
LXIQKFuX7DM+0+UtuZ+lNmG438RjTpQJGDtTbHcVVL1p2oMZ+ioxGg6QPuFkHRK7DeiJxUesofqL
Of8XNmi1jprXoE3XeEUvJq9+jbglacl4WOcll/eNxVADiWUbU913zldx4nHuhYDGAdGDUxJpFbji
DnzBGDCqQ/ZHV4M3WsMeiLWhP4kmZ9bNI1qH61yu/ZsrHb+nmtB1Hp2jTKp6E4kwoTzx6CTDl14F
3HOgfKlg6Vod5DClIVGqfOzPee5t7Mk50FkmlFlDPYYfCbGiEvttg48PGJKmvneQPzCp4zna296R
BFUKlAEHJ1LZjMx+MCx9aXOQJqvTHjdvE6QxrC2EfpMXVR8+zzk+l7WPpxFIfx0V5WAOCijfZU0m
fU6smWcg1Wvu1GDswm34ytKV4ciMxUawC8xWEKSgNyXcDDGF0y3qZrpzJe5fdz3CleHmkqzJGwhm
76r/QjoT9obnL0sseudUdS5B0LjBrjrlBmWYKXqjtABe3Rhg7McT8SOTYtEQnpG5n08MOrD1bhS7
Hk8WiYSr+r2lfy6j1OnxXzBSaj1+TNdZCimoaQil7AzGvH5nEh/b2cVJEK4QyyvcHrtlZ03ce2Fs
2flLcaz9P1B25LA8F64rVG7llSBh4XhTa35V1jEMP4Nhh/QKz5jey1dD1rU+mHJWQlksHQibtbxo
InLcPvcT6IuMbdYqMDsadVVM27YpfRq/C8abyE8AAzdm+J176tNDnGehK2r+mISzksRWqVswiHkq
WYzh5XFjto/Cq/VxEe1fnl9zEkpzXcBvxIGgt86Galx31c19WUqV7nFv8WsWasuI47gjwvO/KK0f
993aPfppQGYlp1ltbfgN6pRRjtOUkuSG/fGhYLhD89rl6UsQSPQJoojqT7fTsyZXy71zrDv+0feh
TJLtIcpqPIM6XUGJhqeiyhkUW084dwv2689QXJZwpZN5jlx4qSsCD9R8CfkPTB4tkvt2Cs2Rgtxw
uvUo5iA9Svpd/ykPtTZ2M51PTR/WU60to+r7LkWZ40K6YYH2SerMQwykGXRGeIKJbXRqD6tnt3JL
L/ijxFDppCkZRsubbxU23u+7/tWmu9OEBWRXxH0YIo0k7caL7819cH8IWgUIcv+kcqxduPEm2QMu
TzWK4QAhDHWSrP0q74lj9ek34a/evZdegDiQpboFM/PjbrpBTWmUFazarfxR3e/bbh1v1n/ICR8m
ooocFVJ8SxDnLoaMQNxnmmD7ctGdir7xxG/EY/MRHfdIEo0BIm16MMBl0zv/t8Qmd+Wkckm8vYIK
LzsQCMmtGUYlTnNRMZke14BLafOJjlueaNHspFcGpOcrHxBILZe9qEIVszBX96lRIK8vSNibFrx3
0f6MeMv8ngZZa4xIC2SKTbpWMf8yjm83W3IQuG3++O/xujadEzbWnsk50EpRGDZT7uFX2AOmPurW
qBfoNe8JxAa8Ow07152FdE774AOx24CvaHeg5Iy4MiUge8vDJYB/ayDQXFN/VnvCqyAA6+SohTni
vZknbmVROeOhlYJEhAp0rvntPhFvBvGTPASwcSz22OGdc6Kl8fG/XQZPUscvHUCFmx8nL6JWHUoH
SiKmIKlsRo3Y7B8YjXklL/t3BoK83FCESZl1I2LzK/ytoUpv+pqG3K6tF2tvDBVquXA02ScVCeLw
3QjPhI6PByuJm1I7vOJ30tu19DTPT+ckS5wUcPKzpMqmJX6E7rlasUjve3J2lU/glob56kT6JpS9
hObLR9NGTGl0/YE6fTcS6353v7P7Tt4CZ1Gsn9FVK1kZ3F5gp3aWTrk33gUrOrWhl+AJM9YVgcVf
RB7vrMh+QPxtEcasJc2bS6L2ml7D5ZDAEGlDyIjoK+guIsA/2fGPMjInYjxGDHvVjc7IYUHpe7Wd
TO3FUu2jc0HxaXq1M25KifCdNFJbgQ3XWvdbtsSZdMuYo7lPTlPJHSKShEREmjv6o/ARNwJ2LdgE
RjlVIJvJlm/9cvtrxG31gcTVwsH/4Oa7l/MbziWAcY36TmRd9vSHBhdy3O6zUs1f1QG7J5DGWIjl
iJS3ZvuyDTiFtlrNyxFkf7gvCCQELtuMSGbhKOo/Bu9F1B97hif9l5VLgYJobyJe5QhGS1kIkdr5
bnqPXZSaP2bHmvke2Jkyfy1IL9sCvJDjiFWzfiK9dpTvcO2FgVpDOL/Jmxv5fa723t6zlaXe7ydz
cQ4FUIyN7Lcfwtnjb147066eZK+34JSqIzxGIRXWoPnp7n6yrBBrJqTGaC8/JBAH87PEDCMTSMr8
BNJxiv6qq9iXAPzbubAOmNUq7c5RSk5vHEI09LiYNT9KtwwUGJZK7pE17pYOjlWtGde0FtjlzVDq
oHZEX/cbUwMxv+sAASCQGZfcA9UacVFWmDqHWZap5hFSt6x+vKFFaBvCCf6COp3JzK191nk0TvJi
ppBm9MjpR0RPqvL9Nvqpzzj5dWbHG7++lbs8MWFsKDrB4atz61TfTmzgtQ6vSp4YcpQkJY9fEELE
wcQfA+GYxn3uOF37dNBJY0nrwceWUaNae5QzQjTe5Ja6HcapRs38PleCcLv5OGFsk1+OLLKHaphM
Tv+XX6OhMrhX1BWVFfKldkFK28OgaYvKo/XxIkmQb0smyb8cPjgLQaXAeVP6EXNhtDKKoO8+H31x
EyiLrimNW3lRnDYFkUVznsQprA1TpUGgVChvYYDAum1MgbQ7INr2PfE2NK/4UPilCySdu8KLS+xr
N2X8KMGokyZvCSwxc3ET6mwvrPhc6dGjLi4UCmLcJGO2Bdr52eZHRQVaFQ==
`protect end_protected
