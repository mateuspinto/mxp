`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
XM9g1ps/vcHRKHBEgSlzf44aZmanTqzmwIdkiREfx0uyuEQC3bLgeH8V7lnLwQqg/81zsvi36fv3
k750ybWOWjXlr6G58qAe79DknJKiMrlICZvEawOPh734nkgP5eRaBR+B1eqCfyiou2pUhJfTqrDK
Bu2fSUP7jWw4MOoe28Qul0vfJwNghgfR08CZftlcaQXYjSR0TmI8yODsElIhIlVx9X30Qux3HdRs
WBYQxwIwsp4zB87fwgDJIpKYuqyYiKHjRQRb/5F/41p7ix/3vMpbierkEdx97j0J1WAY66EchmSE
M3vbUiVtp0QFabvzU4qE+kjlBrYmUGBxv/xaww==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="meZRCMEQk4eF/K9FEhXsPN0NpSZqqsTyVLquafuJN3o="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
Erq2mIWOXAonK4eMgFOYPxFtxiqzOweRIZzFwkUisD12v5ovU7mHnaqIpJiBbpzAXVtbDE3ROTvD
3dN0zwvZWhAiWeHF6Q9Io+rCPd17ZzbnH6++rpSlkFOvLDybXormVpk7OXX/aykv0b0O6GhT5DR8
fCoY0uHWi5TU60CnPNDkCAFvlQR721buwIL2TRlXwYuzIy6UGX6X0+MH4ahnsLMilmAU2rVlr7hF
XQQsnU7i4m5RsIFUwf3Lg0tRol0qO/iYY9CN3b4GItVwU9zjQrgNIuOUX8fW6N5XGG8bisWUj9rS
3/ZmyQEAW8WR9drxyStmu/JiYvWCAvUjtGV4MY10szdNdBfiQ2cq709AQATOoaJul+qGCWxZB9wG
wXd4z7CDTlciVnVFFzNuSMY+r2HGGGoGdSgWKg2D/NQJYiemSrl9mkhhVMxFqSWeQW8sFP4hasi3
SSKMeLNbuLjUokpF73IULYW9eMjul3bg2FerUrjysx62o/CaO9uYMYiRpYtEoksUcpCLkO8gGSUL
ReO4JVsYS/rge0+4ipke1dI/QzdyNG9YUOe4CSbHqo594z7lYo+Yf5keUiY8RqoPxpUxfA3aZcB+
7ZBXTJlmikdZqnBFYGB6bvME6a7Y+a1BEIfBnpb8jwYHL/3InY07m201u1GbShcU17TPQF1fAN4L
11VfL8RA72qG8yrYthzBl5GctGQASPzZXx45Q73Eg6FF04+jRtMGhFXgnL30CV/ouw/M8v2ome0T
g7kMwJgM7lyy43HA4lStaj0rSj39e86gCUX0lb/a4Du4BZbk26fiYqJnTdV6gddkoVsWU8SbUkEj
Hz7nAEcC652eXGxuPF7tNki5CSc7DG5MCOx1Sa3JuvYJTaKEAKwPo7V1py7BhcUFFXfyIM4gvbw/
XeMIDSKyZXcWZGqAxiNTSyBG4Rn70L9EW4XLyQlSO/qx3Xi37NzOOfKMC3yMcfFUME9ofem1TkVJ
gFyO0kjGd1VK0jNd2zlZrOObhfsI04hcRtB3DormvKCEEn2bQgwjMemgKHWgnkSL79FzGZ3jGoih
/CyDyLdadKGdU7x8Ok+T7y22XpjUsX+gT1POQyxVwxLCFgKVzKSTPSW1txUJgC0/xCrkZzGs2m+Q
QdhUNvUWbRAzI1bW/a0Wvs+kPV8lhRke5a6QgCcO1V8iRK72oT8l+hVR5DrRS1nDNEt0/H/EshLx
A1q4f5QuE6aFfDVZUcVrWjAAAXrIfTnSIwricIevzocWZXfyLFOkOIJgGRhydN8dvWeuExO6jXMS
RSsNO5KH9WucV+IkO1oPCe4hC0/5oCiWQfn5IW+JnCkHPE2IqU4zNPH2dd8EEdxdGd0Itb/1kBAa
BWsk1C+R+3wYM2UDSJa/37vGoB8TUh6sxtIZC5r+5Ui0aCs//khSUdT6xvCeeSfh16Tpi2S3c2mQ
JXS8NIK7elcsLP/AODH2L2eSlCIyfyj+BHUdodduGjALVWdgMnOIVMkYfSfMne2pI0FAz4DaP9JG
48JaoMNHwyXZ3iQEiBTWtTWbwmBn4kZ+tP8099xVhkssKKr/1Dp1Vw4DuojB2VhVB+/PnEGeGwG4
kIrTWXvPR2aDKy5B+RnlXWbT7MsaN0cINHSzFtt1vHm7dCjY8DPgQWzeLrLnKjIbDHotHSVyyhjK
bnN/2tMIH4U0YTIy2RrRefttXhOxoEOPb/gF9Y7TsPCFTd16kaL7ZFtybwzn6rVQpo1otL/EmeNV
5jcxVJsfkuEDeOyJKg5lQvrVUhkrWTM0QsykZW7eMbt1mnww0px7hhiblUILyOpA1i5u7gfJhSJY
IePs5uLcDYVS6+YrlMzTHB00mvCKlUaI0VjN5FhDYE8eRRghmGjrKFaqa+a1+FQJZ7rmbLzmmy5R
WTIaz96inVPGnSTw/4dVWE1ntpsvI6bnVu+xiXdJ+HrbVzpAi13TGm3ejePV83nJK0t8mDrz7c4N
lR2i59OWPEIDox5JP1422KLGM9CeXo74EPMPP4Y30locxArZGogcOnrxB/6Wiq5mjVbir5G0IWfZ
nKPJsH7L8+SM42eHTmzadS6OgxkHnnJezUv7Hkwh5EVUNAXd1/ut9gtABP3v
`protect end_protected
