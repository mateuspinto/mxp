XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��y�!H������F����ǆ�7�H���O; H��\j�ubsY���y.!M�H�$ݠO6��<�S�Ĉ/?�}��V�g_�| �#�J��X����1Xg���㗚��J	]��d�Vp�a�G#K�	~t0�_!V�~zf�g��1F��Y4'g��t�q�	�����+s�i9¯�A<��05��i3ȄT�8��b����W�/h"�c&~t�P��e����L�邹�y�x�c��~��	D�+'�ՠ�~��5pZ-�**�����p�8����pkE�����q&�@��Fan���[��+�.$��g���H�ɇdhk} S�#�Cg"��0,���@��|�k�>~R^�׼j��a�/~���t�j%�d�P�U��jL���v5 �W�G����:�V�Î|T�/���HDa|;`��;��c��d��ʣHm�%��Nt�Q���0|��j��;�
��O�`rO)QQyx��m����uё 8l�<�y�-�A#g��^�y�Y�釀m�7�"'�{��'�j�w>4*�q��z�tL���"�z��Evyj��kFa	��d˽��e�x���4N{[_�/Hђ�3s������kӗ4^pƞ@@�i��$��;����zbnQ|��{䥱�Ľ�Ih�������w�g��gco�ɄM�
z�4�^�蟁��ae�O��#fEV��J��[&�:C�1z�؂����ի�P,_Ș�^�ƣ�6��UHz�9@gkʖXlxVHYEB     400     180⍪|[6m]D�3���y���_��}dl,�³ߣ�\T�����_��J ��Z��^��{�wM�ң����+��9����	��h�󥂠H��p1d{�i�����ޔu��y�^K㭍�d�\�]�G��Ԃ�Z0��4�"T��9��B����%�T�!S(k��;��O�}oq�i�\���Pi�{��n��+PP���^#��@����?�Q�E).RX]��Ա�Z<�i4����*��3Q���s��~�>��{��ŧBU[���3Q/�gF���X9O�@7Iv�>}�`�jB'�x@<�iR^����QuuR��-⭓��j���iď:'��Й@�*i����X_v��{���_	�h����N�P�-+g�wXlxVHYEB     400     180��=���%-�W��1�kd��D4�h�?�\�֒���gY��r����~y��F|r��lh��d�%�o�4�^~�=�r���j�s'��R��ql�q�و�1�4��$�0�A�#r��t���jn�t��x�A��?M}"ry��]�E�;j�о¢�� �-�� S
e��)�Lœ�5g̓i!�%�OA�A��Q 
��b�����Y����oЖ��4��Dp�k������%���O��b(���{?��j݅��u��A�yoi�@�݂;�j$��O�)�Wڅ������ ,؆�`t����&IJ���ހ�[al��in���ٛ�|��;��|��u`~���[i�$��}�N�����r����u��^v�a�'� rfXlxVHYEB     400     170����E���8Ѿ����?/���
�W��~#�1�$������x��ʓ� @�M�N�k�����E(���x�䬙�:M�%=��ސ���WLݡH2���
����zí�I� >��x�j�tx0�kj�	h�`���X6e�\@��˵��s� ���/%���f�|����(.�0�Ι�����`L�R�b��S���	G�X��"@˯Pop=�(z�M�]԰�WجEP�i��"-*�����������z4�E��]�������#	i�g�	�!(������EbS��!�"��*�IFxL���C�-���9i��NL��G����V_�-b���?Q\reO* [�n�m�'~�XlxVHYEB     2e8     120��au�g3��\n�
럹?��)��ˉ���\"W}`��-z`��C��_:�Xۆ����Oy���mg�Zs燁E,˼�(>�U�iT�wb��K�rGY%��b,B�^��]���PNj#�.��\�V�ƺl���ס�@s�3�*�7�%�� 7�P�&B)���P�@��`�z>"Y��'�)R��geD�Ҫ7��eXknb��>��Ԛ�/mÈ�?Qȷ]'��c�P*��#�n�Fz�`M�e~D�4��f�:�H�Ϸ��1 V]�H��'j�W�U$���ʍ�'�u��