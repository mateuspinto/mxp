��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���>`��tvM21\3�f5���d��(���ו4�q8".��<�/	ĀL���ߧ�~6��i���OŤ<�>: ���l��(��n�9�P�٦�����7|�O�!'c7�9C��(��Ҋ�V\�A���Z�T[d�K��},���ݟ0%�f{s��!}Nm�1�fOeH���+L��'��ߊR��Ӑt2��K�a}"^$�d�@+�ˣ3\�g�?�RH�����Z�O����S�oW�{�"�����
��f�h�Z ���m��M^E�Z U�OjYB�5�!x2��2���.�^�!�.r醠�ff���j����A)�#4�+t�/7Y�aeH �Mg;LcK��c����eWaV�P������������� ��ɅIHA��2�Ϗ۫%9u�u�;������ئ�at����u��A���A�����Ƕ}�i�J�5(��㌩,&��z�f����X(e�k���~)_7;)K�(7�=��Ui�J{=��p�+�Z_0/�G,e)ȯ$��c�����{jB�á��C<��� ՝��O`�MȘ!)��SE|�3�n�{������;d����y�RPA�Q{������GO7��>��K�E���C<^�!6�A�g2��o{����lf�ه�^W��R��������[��`�@�0e�r3�G�h�;�܌6W��wh�M��p�z�PH���k��o��p�+!�/A��G�>���xe����D���W�G>N�e �@�<P����ݔ��΄{�q���߯�N�j��46|;{h�jG�)Ko��a��U���I��Z/�)I�+��V
�.�Cr�&aYa�hI��c0_����{�%aT��q�Y���g�V�T��M����Q�JI�d�`«r�?��l��T[uJ��>vC\��0+6P�C����(>��_���+dZ�u(�*�YϩN$��eZ�vńա��o7C���+����/��Y*���<�x�UF0ݪ�wۚh�e!�q?W�����&<�� �D{��e �#w��w�=n��]y��Cn��o��/l���+܄0Ļ�,h
]þ��@������#X���O���9큗�z��묩����*���h�����H_WQ��Q�V3�Qƪ�`b��Fx����P�l�;����wP������]"Rr
��%���G��I��^�����~�i��<��1-��@)T>�0S7oG���Z�����������$�\��jfX�
���q)�j`���i2��E����/������ksv�b�t����$�Q{����CB繎zH{���f���4�xI�slC!��'ͤj2��-b�-�����=��,��ÖJ��ot�ޛm���%8��y1O��.T6�^���w4��oE�]Y6��S