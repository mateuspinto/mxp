XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#�4 $9^G�<��D��y�"e%��GQ-;�Wʳ	��U.����]���� ����w4h>�Km���[���bk�@����F��wf"��.`?��k�4~M�>�A��b
��"N����ia�0_3	�Q�~���r�2xi8zV�|���j񨡃�D�c6�z��#�<{�X�V<r6�w���R7`e����&b}��$���(wޮ��Xo�bN*Nh�}w��	�x�nz��v�- ^"Q�#��x��P�9�v%��D�T����tP�� Zu�n��*��jI�s�u�g�OY	��mD�<�f�'�<��ß�>�Nih�s����{u&/3���Cqd��չ��+"�!wzP�go�X�ε3]3CP�#v�	ŦT�!�Υf6^�^`v�P��϶�S^gc|��V�.��Zfc&����OyA�6�.w,�}��R��L?���O(i�=τE�c/;�7w�D�$GM[Q3�ٖ�vT�!��^;��k���� RH�f��p~,vy�]��N�HZβ�[��d��d=��.��9 مc
��F�)/�߿h�Hۮ�T�H���B(����^ɚ&@�	�\����3�+��P�CB���Y�+�����e�`��5����A�����ͧ���IOP��>���g�n̊����<���-/�ڪ��/��D]G�U�*��o�03�=�-��:�h��l/;�;�,uQ���2Ȳ1�ݶz<(][�U�V��U�@�JS����5���Њ�urly��,��XlxVHYEB     400     220,��<�V����p\�>+�g�S�5�.0xC���`��=�~)������o)YҘ� �������5\g�6֌~j���dn!�s7dŪ�u_��2la��W��KY5t7\?�v,wj|���%�g�U�-yԮ��2�������	�t}�I :�=�%zUU�>�.6������t����#v�T�<����*�J/���"��[���K�����Z˲%��U��U3�@8�Oׇ!�Y����V?�A��.�D1�5�x�wMuP�I�^�c\ ���ը���ia��낷�� 4{�<R�B}QG�%�3�]kM4)���\���8&`e�#i �y�ׅd�v��Ԛ�,�G�i��x9<e�,�9¼?5r ����~m�rg���)�L��XS8���G}�1���J�;C�Pf$^�st�Q�o9IGH�����x��_6|))-�gJ��o�1�0@ iP��Ё��c?s����|�~�tkE�HN{���Η{���2
_$>��^�o;�R����H���Cj��}�z��&>ؐ�=̓XlxVHYEB     400     220o�i�%$`uF�����6��\!y���u�Lӆ���`$�P-W�u�Ř����zm���>�`~n8��/sE�N�h���W� ڐ��l�?��{�B�Qx��^�/]J�r ���kM?������sc-����|;u]���旾�[�GOtV�K9"i�ɍk��;����3�&3 ߽���.u��e�?�<�бo������5QB̴͚�� �>uFg˥ꨖs�p���:�j�!��\�*,_NPN��C0�~r>��H`��.�M�y~�GI{W��C� ���� ��tJ� ���)\���#?�)A����mʨ^��$�����шm��{4g���|�/�uM��j�*#7sԆ� �0�;A���~�q/3�;�[\F��3���������>=�Պ˚-���,�T��+h;�r�(N�ۡi	�d�X���ť믲�X�y���1��ټ�N�l�gu��}o��˫��|��h�=�5M)�F2K�BA �@���d�g�S�KZ�tF_[J22xAXlxVHYEB     400     1a0�DI��6�_uR �8�s��.D��A��<AX��c���i0W��Q�֕�;\�玘2j�m��̫��8P[/�u6hN)c�,����y�Eì6ɥOa��,�]o�7��T�.ZS���q6�Hui;����]�v'���|���X����'�]�qm��t�C�/�|3���"@FV�����Ǔ�\�W�ΦQ�t�N<[����1I�X}ɉs-�	F^����]؛���<�"�(�H0��e��|9y��X�?��7�ۘ�O��N% 	���+T�����Kxfw��Z-[�I�3��_��9�1�]˞w�N��Pc��1�,�n�����E=�ߺIh%�qA�$ Qڢ�z�\��杭�7�BA��1y��Z��ʋ�e�<����3��݊w�����)�XlxVHYEB     400     130b�%,��{�F�M%dS���[�|�M?ƹ�_�&�y��S�f����?�9��ȃ�=�oi�;���� �B>���_{0r�%Lg�6�[�۳�ʌ�()�p7�h���E��ķ%�m	�ctÆ8�ƚO�o� �(����kf���������%���흝Ze����g�&���_��)գ���ņr�+p<-"����WO���p�@�}&x�Sgm��L└�ǡ����,B_p�A?���Pr�+�j[���ۯkҥT�A��Xsf�"��k7���2��/�H��� ��gJ�y�j�cXlxVHYEB     400     140a���z\c�韋�o��8��2�ʏn����a�4��X�u�m���i�X��d�a 
�;���
�h�R��kLy7f
hzD�>l$�`�2 3�/q�꣈��kc؎��z���Cm�T>7��;J�����Y<��Qps�b�r� N{����PK' �,��Ya��oOu/M���.Ye
��_P��� .,�G��c~�w%j��v
�m�a�O8r���L�:�`�xRp��i�e�'�)�IL�����bz,Ka-U%�c�_Ƃ��b�H���=�<@�����zF,�F�� fQ�Y{g���'9&��XlxVHYEB     400     1c0�Z��?A�s�OR@mf��B��@xHijgf���-D�q�\��.��������a�~����\7˱2��(9K~��A�_�>O;�� '�%e�n�ɶ������Y~/�� ��

;�ښ/74�Y{�y.KR�͆���l}�ŗ) ���,5�(�n5��L��Φ	U��ڰ�_K{�[��Tf��އ���
OhDn�C�*<�F�l�ra(�.�t�i��E����U��
�@�",1��x���l<��)���^ ��(�D(��d��~����?0 �Ը���������K����k!�ɷv�v)�Ю�:�õ��홙;�U�����i��Sf���	\X�v6�r�I���5��^�3�W��#��r������]��1�$S0�����E�t���-����}R����3�����H��cM%��AXlxVHYEB     400     200L�Ӏ�'����y����)�Q�"i���v�6�:p�i9��N��F�-P�UOgeXYZ�Z[�Fyr����$��&��`YY�����}j��m�e���|�^���P�=�&*'B�����O�
��������)T�h���{��;���2уѼ�����1��G�K��#��~ɒ��~�p35� D��H85q:�񅄚�j�VIy����s�h�4��᩟nfA���7��0G6}��b*�R���֎��S��Ex�M5�r�)��?xqH7 &�hU	@`Ne�lGH�*��S�#s����o��̓��'�<>25��4}�ￋ^�OC�I���5�/��m�P_Ɠ��N<frp�K�LϾɔ�
�U�4,�ݔa=�ˌ�1����re�N١�����,����mu=��5笕K�jF��2����lA�F���3��Y���X�)	dv=��tY!W�X���@i����v0��㗼�)}ko��ix9~�-Ë��XlxVHYEB     400     1f0��	+vV������3����w�ʏʨ)�:���$�c��{�ཐ�H�M�0h0�_���4ӻ�HG��{O$|��XNfܗ��T����-���r�T-3b۳?�<&�����q�۔E�Z�{�Ҙ`�H���{S$Ӹ�c�*�ja�l0e�j�͕�����4�~�r,�閡�����5���sS*���`����W��_įL�!��r��D#%<��:Y���9�9m�D���#��ԟ���6�Vy���g�={s5�W�j��:"�^�u<ؠ$_�uz*�,s�xQÞ�kH؜���5 ��׫`�
-Q¤ݨ�8�G�bt�}{.d�EA���[o����IY��s�R��"�_4��XahE��e���oc� `�h�����ḱ�5%��m
��3��#��.S��qg�q��]m�d��qa�C-�6��N��YYXy��M��K�j����^��J�b��ڂ��W[�ɤ�@�o��o7�XlxVHYEB     400     1e0��M��B&��X�jhM�I�(R��t]]� ٿ@���������v3<w���܇���#�C��H�i0��݂�+���!w�0�y[}�9��SN	|f|�n+�7��[�-�P[$-�!��}{��ŎF�m����Y��DZL�?6�(�\�-�d(�w���=� M��I`Sd�ŋ������k:{w�<�v�RV��/�*��+�M�/��.� �%Mq�7^�b��,;����3UF>����ޭ�� Eo?d4�I��Y͛���
��Н�g+�y�/S�_�rFD[�$[�v�S@1.�����Q����9���kA��*���$��,,��O�4P���к��k�����:" ���=��`�x^j!k3�R���.�RB����g�ˎ�e���$Ůp�v���`�;� ��Jx|V���8@��s�%�w>yD%~�\[�|�\�D�( ���:7YG�m5�p�XlxVHYEB     400     1c0��>Ě�\j����n$�7�t�!t!�>J�aqr7�F����Yb4���GR�է0�Ff¥K�VE���+�7ٝf�p��⇫G�4�̒�x��%�-��Sڪ�3���]_g��b��i�]�%�7�[�%�&^��W���GKr84���ڿ�?C��*}�׫&k��N����*�w�v�7n��˭�T":�))�}���O���V
ꡕ�<��RY(u7��̯����6�U/���A��'m��}P'�;3�$��u�?�	�:f�Ւ�CN�w���u�CnQp����N�9=�j�$N6��fP X�<8��e������:P&��^	��k�9A��7��8���IԑS~�n7i���O��ꃔG�\��b@v��q�o�y\����< �'{i{C�	],�=afW��]x���dW���,R���-9�aN7�td�MnF�UXlxVHYEB     400     130B�:X�VBW�7�-�;����@^
-wZ��L�B�k��ʘ�2Gu��ⷪ ��,��,�bi��ρ���\�u���N�WH�l�$5)�Uz�ʜ�S�H�	(8]��yr�����B.¥EEV�%�H�9n�A��J0����~�5'�P'�� 8� 3�k]8�⎠Z���m�_v��Z"KIf�ȸ��3���V��z��b}�VTa��}���L�ם�� y~j�?%��?�-���g�v핤uƉ�� ��x%�Evs �m�h���Mu���~t�z��(����I��M��U6���z��d���<ɳXlxVHYEB     400     170s(�mv^��:8D6���tI4��l{7v����n���"�Y�)^V��i���(�xt���u Ï��~���z���"Ϡ<�.>�t�ť���3S��L����%�J�����`�Eud-�F��1�G*cH�ã�2���\e<�jts�N{'�`�Z>�͍����X�3�m0���:[�aQ�����f����g�=jC�y�ʂO(�Ө^�f����ez���:'ทqS�>fh<��4͈ؗ��3���.%i�d�_O&�䍬J����s@M]^'��/u��;P�Δ0$�B��ɏ�"�zw����х�� _����F��6�������u>Vq��³!���rs&�"-��$�XlxVHYEB     400     110c!�5�PѨd
�X��	���%ʟu�襇�w��Q{�=��N���|��N�y�Ώz4��q������S�J�8܌=\i.�D~��މ�{?\H��8���$6�M-LP�]8w�Vt��e�7R\�3:����\���Ǵ��F��%W��~j���B�82]X���Vؙ����iux��� �u���`��/�o��"{��7��yr�]�� q	�\~~A�in�&��T���� G��2Uc?��9�)��@����t4��O�?��XlxVHYEB     400     140`|T��?%���Q��z�n����&}���A%�ܖ��YEXA'&���nkHX�&��h̏�-���!�����c���5ݑ���f�V
�#�c��'ME�tX+��S�=�9�XV���9��v�����I�m�h+2��W���l׆/��uŮ���~M����"hsLM	�p������P�*t$�U)�X|��Q�S���An�\���Ї�Q����l���|��bi�۩w_R�Jv [Ȕ.9����S���X�ۈ����`�Q��ɞ�_māS���6�0$�����ɡ�����<��tV�ܿ�"=XlxVHYEB     400     130�^i� /��R%��8�wqʾ�*MŹm���7	���W�۱���C�B���p�b=��{.�MWA�*�7`z"v�Kӊ�&0L\�
{��D��2��\���|�I���>n(�!5�)L�¸ihf���.B�@!�3��zql�'lz9����
]{#��"h�+�jj������������'���5�+�7МI��F;�5�\�v2�����im����.���~\�95���t��}�\�(�nYu�3�s�������m�p�!$%ى�x~[N���T	�WY��K2�;$���)sR��P��XlxVHYEB     400     130�u���Q�����D]�)�p&3&l��mmLi̮��'3�!�73 �<�����?F�t�1-8)xE��q�Ⱥf���ڤU�~;����v���$ʦ�h>q+�t,ax��Ȧ<���voE{�YNJ�g��:���O��1���Pķ���`1��lv��,z�ͦ��HKH��2!�Y���ek����E^bsϱD��Yc o���jR����zM�J�4��I�]k���Ǥ��0�|}�����O�X	�N���VŢ'vu��vw���X�٘)8̹���y�=�+ c�XlxVHYEB     400     150�_UVH8��'�-1��� U
ҫ_�&��^��/)kuFW���� �X̵��s���A��0�����ac�X
�-!��}(aO�c|oi�Ä�A�iL����i>'�8�5I�	[CH8`�������ɣ�#�K�W7��0��BB�S�8^���ϖ<�6��,D�sOb���4^p�^f�����1
t�#Ow��؊:��l:��'=N?9E�n��٢e��dVy����y2���e��U#VL�:��
��Y�5]rL9Xz�BCt���GVy#X5ʋ��qO�R��L�Z)L� �Е�޷ZR���&�����'<Si0����XlxVHYEB     400     180�#/��:g~\���i���>c�}�W��j�׷�I��]�{#�y2�d��.��Ҳ��dDp�UISc��W��:f{�t(��i�Ϫ<tt�P����z�2ͨ�MvH��*o��w�>;i7�|u7���J����V"O 7�'�J�Y[��{��:���-�|܌μ�b�����oiP���5�_� �o�!R�Δ̥曳�%ޖ�`��~>�I
[[:�^�q�IԬ��j�� ���s"�^��E���3�I�w��"�֑�<�*�V��X�Ng�Cߗ����GW�	��(W���1���/�ؓ�7�;SӴ�[��\��U�ݘ���Qc؅c����Q�>8V]�g�m������}Y�m�؟�!��A )P�|��"�|х�XlxVHYEB     400     1d0WFl�\>T_<u����WT�5]�ol��G�_[�>�O}� �A�Y�77*	��f��0��ј���>�g�D�|��*�8���3}��ձ�.�ȣ]�	�������ޚ��ì�I�.�S�M&ʹ�z�9bc�J"~=��n;��Y�,Q�6�@f�C��Ud���P�����U:�t��ȍT�����㥜���!S��5�Vᷳ�1Fʂ�M����WqNY�(F�ZUA솲n�b���J]:�Q�Oz�?ݕ�I�}�r1��~%tMHr���{��6?l��[�pY�0��|¬,Y�iS����a �q4Ump[و�X[<Y~5X��ʲ�V����!]Aj�Ҧ*�9hQ�q[b�\O�I��'�
<iJlE��*�#bM�������^QΜ�3�l:|�t�����.�
#����i�8�T���x*���5�y��hؠҍ��v@XlxVHYEB     400     180��}��;UU5r�( TMR�U�L�I�"@��Cy�	����)|Q����!-tX>���!*M,�B�f���>����A�1)s��n�ֹc_��^��3f9�J���Q�Y��6�W]���F��k��(�D��IG���k;���W��:C+MAF2q$�3D��.X�*��U�Sm�u6q���յQ���9��ɼw�j%W����e�it""��A8�\��S��%s|ri���i	e !͈�f	qr�2�Ĉ���̐�S����2�m��o	q[l���&\Y����xZE���ԭ[ )4x���L*��SS����9#��n�O%�A1>⬝ᵄM�qb{�@@J�>��zo�Eb]��vGdGEr����XlxVHYEB     400     150ͤ���K.)�Z�b��;d"aW�&��+룚;��dܕ	�.� D�TQ���L^�ص�8;�r>%�	��it�C�]*�A�����R�u|kQ��5F�t�r���j�Ik�ϩҍ�P_�C?.���
&�W��KY��T1!�]��'4B�8���o��d� Ibr� �����
��
� w����k�mE�:�臭�ZDmma-N�	ɪm#G�/��4�^8;��6K1��{�ȋ1�����x}R�د}���G.�7	1e�H����=�_�� } v�����ʙވӮ&����>E�!��h!P��[}��=Ԫ��"��=M��^nXlxVHYEB     400     1f03x�~�TQY����X}g���$�h��m���a�\D��Z�^ջ^�|�ų��j�k*h�2���;F0k���P�̭��U���&�{Q���f�o9K�I]A�U����	sbMZ�#�A��z��c�����(�������A���?m����	�#݁�x�E��#��w?^�g�	�ITŋ�sԿ�Y��=p��>�m��b?������m�%Ѡ���5�.�*�i���+��w��G0�T�lv�N1V��� ��o)C�R�� �W�#+��Ɛ�m�&b`�"Y�Sq��~���	�8-�M��Ԁ}^(f�ĤQ����MFh�,aR��.r�c�Q���4�P�}��Zn[��E����T��N�Y�0�Z�?Ց�B�T�b-��\i����UŠ�h_��I�)	^�B/���f*k�O��L�:�w�y8��\��Q�ܰ"N{�������5k��^�g��ʘ�]�?xXE�Ĩ����XlxVHYEB     400     190��^˵���a�m �D���mx��9Ai>�Om��;4v��8�Xe%�z�Lb�ú`�
�&�cX$i��y��M��=����!����#$u�yry5�dP-(�#Z�­�%\��%��O��Z������L�I ��x3s�m�D�>v��	�5�c��n6s��׺����/P�az����u{��Z`;�v�X���2�+g���A���G3x�4s\��L���N�� ���u��ZEK����$8G�1��~R��~1WX��A�Z���X��SU��_�>��'d&�s���N+�!`�\����ۆ	>��-|qƴԌ��/����9�n����˔nF�C���@H�*�ʕ��[zw˔&�D����Da��:p�[1���.��F�iCXlxVHYEB     400     170��B��a�g�7P���~��*f�t��/��ڧ8�=�,��Z���y��-��b��iD�y�i�oLtBͶu1%�>�9�,d���@����xj��)@fy�����]�KG{h�g	�������õ�A�j���Q��%F��V���sj���$5�Ac�(.|��O�G�h��G��Z�zZz�>A��)��x	�Պ�Z�XD���s����lےJ0\�)�@`�~����!�(�M��O��R�ϫ�j@��S���b"YӋ�� �\��~a�H�X�$Ė4+�GcW!�V�f��RR��E̰s�$���޲��Cx���Upq{��CT�����b'��pB�$9P%*���qr�XlxVHYEB     400     17046
��Zqٍ ��	��_W��Ȃ0˱�`���`��5��EK���ʃ���Z�!�I�~׽y'���F��<��G^��е�~&F���[�.�J��6�CGi(�p�f��ح�Tx��-z�#x����"����r�@*���������t�BQ�����ϵ�wa��kc��6����pr~���'�Uz#Pc�CLM[7��F�'�`f��D�¶R�"���~��,��.�:0C(�m�֨�ja��P�5p%�V�P ����$� 7��#��H>����G�)�KA4#G�:�^Eˡ�)�V��It��q���� g�q��ύ�'�7N#n��˂�`AL�Sy��#����2����XlxVHYEB     400     110{J�ԡU���$�w���pX}���d�}K
jPn�42�l�f*���F�����,|�)�9��y,�x�����n�A���Dˇ�<"c���Y�r�t�����M���
�@��m�%$ՋN��.��z���I�d��K����pN�Bg���h�~���|%��[�>�隁�LI�N;�T�J4G����ţ�S��8"�E��dq)2�c,�w�0�})C�F���������H�0Fr'ڮ!�w�;���r�����
G����XlxVHYEB     400     120#ӈ�@ǆh��'�Z3�'	��m/��tf%�x��vJ�P$�l5-�_Ҽ�rZ�!���Ү�&<�R��i#��a",�Æ�L0a�͙�h�����-~O�$,Pd3�^u��JM�;O��N���>�t]�9ȉ��;`>$���5C�ϐq���ܕ�|v��"�1(
tp�0�Y��I��io茺A6�E9����A:'x��5v��\'��"�Qֽ�>S�]p���	���ݔ�Z�!?l�BQJ�p)]*v�*!�^��V_��(ˇ��(4iY���U���ђ!u�?�za��XlxVHYEB     400      d0j b���'�o�#I<��Y�Ejeդ��zX��g�~��?�v��ҥ����ٌ��Nw0#�9�������x]�J^�5��� �}����gQ}螌���i�BW�8/i��.���(��."�!"-����"�ڭ
��0�{�q9Sy	��^�.�}�l
���|�a���=SG�J�b�1(eL�P"5��`�$p���pO��9Z�C�zXlxVHYEB     400     140�!26e�ϙ��xa�|>��\����׬y}�*�\�tQT%Q�`ߊ����(��L!���s�oR�&�|�	=\8�?GEq����o��(��]�2TS�{�K�jM���9�I��C�%	��
V0WE�z��CF���؎W)+���r���Ѓ	r`/tb����z�C�dB�e��(�j��%&�� �� n:�~��=׮�O�G�RM����}�wꤊU ��h�2�@?�%�R� �� 504)�%�x,�EFz4����X�_��ub�_�Mi��ufi�nt�Qf*��,���Q�f����FTXlxVHYEB     400     140|c$P�IT+Ф��L��k�����Rg��ޒ���>�~H�E%�Rٶ����BFiQ%�;4�_�)N"�5{h�AQ{Bb�
� wU�+BI��mQ���@H31�7����\ �d��d>���UB2����Nr��.�K���aI+���
Ǵ��;v�þ�W�b����1���P���	��`Q��]x� D� �t��vSQ�?h���8�K9bgB�	Y���xف$�f;��mi�T��9]E�t��(\ K��5�g�s�R�k��8��
e��Ff�7�S�^ �)-n�Qq[�#���쨮�@�-XlxVHYEB     400     120�~�c3��ś����jM��v�|-eɖ���ND��VKΓ���Ű��g=ޕ�~�Tc{w�R6	/�,>RA���s��_��xU�VD�n���S��s&��%_ʶz�k��k�h�T�C���x�`�'A��?�2�vlW����m��ӆ�i^����z+��zb%=���H��P[t��2a4v����ӭ��p��,}p��AX�i�bPO��Dl��_~j|œl�2��v�Xd�P�����C�,��(��K!Z�3c=��Yku��<þ�zH*�
���XlxVHYEB     400     1a0_4W�x��h�&�?>�D�3c�3��w�?���fK���+/-	Әa�k�G1����»\�8�Ia��p(O��mmڠ�B59�6«dԸ�+�ּ�O�}O-�ʴq�_�ٓ�;j�	#jCtU��p���	�Hѷ��P@k�j���7AJe/(v�N�1�b�2�	�U��//7�5�i��84�Wɂ���ɇ����&�׌�JZ��u)+r�/7pd�B���J��?OgƧ=�׳�q���2U�t�a�p�.�p�&Y�a3�7~QTֱ?��6�iv?�Y�!��[<MI�W��Ӗ*�L��,8��̗�M��6ڐ+�{_w�e������%<ay��ǌ�O��V�����Z�{��j��lחo~�ڏ�!�Q�q֞�`���u�!)�����O:��%{���<�QpҰ�XlxVHYEB     400     120�^��u��RL���M�'��I�����HA������
�ۂ���~%V�&�8&��jҏ��>�����$*�I�8IL<��I, n�q"]r��7���#��X�@��Ǫ5�ڞ޿��`�� �Z���ѣ#Yq+�<Y������p�S[������զ}�t���6��o��"��x��%���D[������ך���(R��i��И��ȧF@����I��-+@2���R;����x:�a�L�QVi�s�b��B���n�Χ5ą�1l(��w�w�s�5�XlxVHYEB     400     180_�����N���1*�˥;1@{��B�T�l#f-��A���G����`���}%HoK|!��=;,��b_8�8�^��mw��@����L��S���UC�{�d	���k�=O��|! ��
�]s;����s�f����[ ���>���� k��B�����`S��1�t��.�GS�{=En�h�=�����(},�J�?i��Vz���d���,^�����w?
�<���u�2I��ec�PY��v|b�AӅ�AǢ���"L� |�7����|Ѵ8��������oZB5�ԝhG�j� ��- ����c�Pu蘣������-�wdc+�������Ż}�`�r������A�뫔&�y4B��x�9Z�h�$�Y"#XlxVHYEB     400     170��٤`WRYe#3��s�%-[�)���n�Ѹ���5́��u�������]#��g�@��9Ne��,�A�	Unr��c�����t�)i�~TZ"u~�G�	�&�m
ʘEj7�7n��i��G�e-�������3�*ީ��� �\��SK_�ێ�Y�Ջ�kW�2��f̙�p�j��|=�nnb�ݠ��r�"��5?wդ�@����)�8�N�5e��q� =q(Ӕ1VEN�`����,���m}�x��&I�Fe$����j�R�؛���l�uyz;:zw���s��m.S{^lW>�KsU(������@l�_X�M����`���6A�r������(n_�0Wd�R�Le��cqHW���
Rs���XlxVHYEB     400     1c03k�u�ֿN:��k��!Y��HcvRQ��j�z�e��iE��i�g:�l�Y�m~��{B�g�l�w:��C�
q�����^\�M�k�C��&6��n��d�1�	��R ��&~�����h�K�0��:8��-*��+�<�WT�9v�8�]�th��xht��`�$�m�H��&(��&K�����S�\0��{9lt<���r#&M�(�u/{�Y�(�Ue�v�(�O��%ZV��مz�8�R�R��7z�DW�n�=�1h"���b&KT�)����й�w4�{Z�>`>E��))���A��bVJ MD0?��V�s7��4�+��-dW�8����᳭�#�ߌΤ�b����CF���XHw��V�{%s,�P� �%���YL ��3(���0���NE�����J	�ׯ��^����Z��[XlxVHYEB     400     110�|`��x�J�[F�o���]����Y?���q�K����:�z�V�*@���� ܯC�F���?���TcI��T�M�鰀�4�i�`������;)T4�V�Ұ`�����)%g�������p���]jvo&����֚�Z%g���� 9x8� o�SHL�T���Tw{�D�v�.��æj(������d�51������+���+A��SӰ�ȅC|�.��
�̥i8Z���v�۲f	D��v�4}�����!��;�}`69��XlxVHYEB     400     170����;F�e���`;t��kXGx+���R.�8�'���s����.��#��da��'�E���;z�f� V�:ёK��@�|k�a��	�o��j�'[Hs��_�؁�a��}�k�ѧqޯ��.'��t͋3�;��I��N0p�[����RL���>���O&��ޢu�=9[M}�QE�=	�]��y��sc��j��+w}�v�q'V��^�h�2�����8���T�j���K�ƶ�K9VXS�޵.Ca`bc6J�|���� 8H����ng�X��YIٻK��NY���d��ND�s���=�c4S�c�Q�~��a.�eGO;j�%��I�*��<uy��.����(݀��͔��M�R����pbsXlxVHYEB     400     170:qtq��?�(��Br��/���FI����~�oJ�0��m�r��h-�Q�!I&�� ���6�=�9ǧ�\a���������!Ċ�7������H�<0cY�/#3Q~�%mߖ��&OM����dZ,��r��U�����Y�*�4!�E���`��b��yYGL�Z�Fl�����JW�إ��V�TH ��r�j�+Qs�i�æ�BWҴ��
{9��-Xvz]�l�7����<��ϫQ<�լ�c�0�7~�Kn���DD��m�o��=fdPb���)���%i�&ff1̗��T���2y�-{Ɏ2�a�j{��?��uK�*�rW;K��v\u��o�G4ԍנ�w�%XlxVHYEB     400     190-�r�ڥ$�1�mh ���Z%��_g���Zmh��><�#G��4�����-Xr|mSk!���b�v(��c�ǫ���1O!��荠���&�Z���eER;u��X�?l����?S�����調;�?-����x�$����څ��ft6��S[�{_ ���Do�a����;V��\�O��p�.�_��TIf�4��f�4-�*��@W�΍���s?"oi�t��/!9\��V�Gԋ��l��H]B���g��_���R����}ގ �,��~���x;XΐT����4~#	�o���p����Ik���h�H��� ��Kk+K`? �����xX��J/l�+Ѯ���>N�g���H���V��l|�c���e%7�
�K' �����ZXlxVHYEB     400     1b0X,[�����E`���5p��Ω�I���z׳����j�9��"S�����ٔO���k;��G�G��	��n,�?naH��1c[n�Ito]���J�o�kK�*u~�U��rN��b���\5�e+�-����J�T������l� w�)����\ޣ�#������R�Ox���V�-|��+u/'E���н�ݨ��� �&�]xdN���O���6�$WDQ�9��M2���i�\9�3�I�^���W��	��v�H�I��ԗt7(�X�e�Mtӛ�aq�5"e��gSÇJL����2�3��C �5]�{�ܙ����	��4\�Zr�o�Oy���>�k��{q�cU���_E�[U�$���g~gb�xpN��;B��m ?��RR�Q��U�.͈��h��|����d�V�ֶ�mʅ<�ɩ���G��XlxVHYEB     400     1b0ga'WB�l���_�BV��ɲz��p.�XZ���I�$Q]2~�g�b-�m��c�dL���^3mUw��/���C�x��MX�����NI��U�fk�o�
�t���r��(�د!�DLH��g.dҼ��Y͍��Ѕ!�h�R&6h�$���)��l�cՃt^�1&���tx�B���o`s���yR_����`�R�N>��|�j��A��7=��lM!��������G`�P�}E�p�@�r nY���%ȡ�z-@�\ߩk�Q ��ЛY�9��{e0U��2�h�$�P;:Q�����J�.�@�!L9u�����Iå������ܗA��Ry�Y]�wF�*��mHm��.9a��X�B�fM휰��^�wp���P��F|�5�at��	lZ?��
gNw� G��ė(��Ġ��S�5�C2�/�XlxVHYEB     400     1c0yp��j������@�r��?�Pm`��ڭ])�����0�
G|fD��ߓ�@{��k�r}2�|$�9\��K����­��y?:�d�{�l.x��e�����*��C�e_�(Y�t�����{4N�v��7�2HH��C��Le�����w�������C�� �"�׶��5��])�j�����%�th��R�fݐO#�>B�J꼤�&��q��(�J��HTs��X�Q��gXB�n�;�F����4�R�.8j���̯M�GQHجC!���+kJ��Yh�ڻ����J�C��J[�����;B���s�n
}�i��h��.�@G�gկ��90Z���.0��F��q��+��N�c���O6������x�e���-p^ڱy��@�޸��'��$k��5��5,�^th���-��(�5��ބm{�:7��"gױ����XlxVHYEB     400     140�d��i��j!�rxIU�Z4If:�+�*KdEГJ��wS�dq�M5�	e���)n͸f@S����ù�oMk��7�}r�!�Ô_��_Ǚ�F[��s�'�c9mh:�g��P̴���"�}猅Wv��~��(2w����X�BsD�Z6����5���&�|�#�tyϩ��L΢-���ˮvO��H� V4�\��s��*7O���'�$g�r��ʖ�N��{�� �t��T�f*��H�cTϟA�_W�H �
��>��E�"�N���Lb�'D�?�ʩ1Y&ɇ`aI7��֒���a�Z���|lpΝXlxVHYEB     400     190-���ە��*���z��
ύi��� jG��N�6weT
���$��|��Y�e�l��]!C]GI��������ܒ-�݃�i�BM�l�C�Ă�:���tQ'�8��[GVj�&�f�H��Z�9.�M�ъa�7��r���o8ņϦ+`#�Fg̻�/���.L_[F�Y��N�����|��:\8śn�O�L?��R��Y���j��l��>:r:]7�ؐ�k��Ή|T����%=J��Uw TB���O=L,�y�|4՘6���g0���:�=��U�tR���F�U��j7���$��hn��z���Ƕ\8��f�$>O���)@LR�c�����<z�pW��?�B�=������%�
�N�$�[�HR�2�k"	Q(@�r���q���oXlxVHYEB     400     130�n�yµ��Vhf�'Y��-�\���ԡ�NK���W.FuZL����Rkv�<M��ο�w�o�����Y��g0����t� oPϭ$����z���;��,:km� �݋l|c0$! 2s��F��t�cs]��n��G����▾9�~zp�)�~:�tP��n�u��h�	8:d�ҟ��eQk%D�淃�}�֥��$W}Ð�v��KI�3�3<����ňr:.���QN�I�X��3�������`�(趁-��s*����9gAK�{e���M�t^*A(�J5��^4XlxVHYEB     400     150��ID�كb�b��>XBq����kA��7b�tg{�5H�߃������'��Rd��;��kF��cA{�N
��wG��t&�h��$D���ݥ�c� ���:�+e��g�,�7�*�7A��٫��~�v��N���p~Q$�Rȹ��.�4<���O5	L^�#������-�[JZ��tK5�z\Gԏ�~-'��`�� 6�}�H1��yc��~�F�HXcʹ��k��TXW�����f�P�B]tF��Ē�4[�G��iF���8�/���1��Yr;cU�&4s�X�u-z Z�[�z��g��ྲ�!.��!+��_�J��գySXlxVHYEB     400     1904tN$Sw�R��|�c��j#�wdK�_���C��Y7^�շ��YV�TL��؇=gr��O���4�#Ww��7k~�,_�"�Y�w�Q���S�$�m�/��?���=��*5����@��/ZְH0�ǫ���i��7�+G�:�_{՟�E˱�ɇ>�銐��/M a���h�����8>
~� ԓz�-nU�ȯ[-&��� ��0��^��yTB���
��%�[�P�pX�%�p;��7���m�<G�7��Y������IZ���q�9^��DMĹC<����h��f'c>C��{�[(��o�=��7?�ϼL��p�=�J!8鼆�������;�zWP��h�r%#�m�ZIv�A�H<��cgI�f����U�7�M7"�奇S�kr�	��-}]�d� x9�XlxVHYEB     400     130��4e�#�'����2�I<�K��f����VO�}��?�)  ��|�·"�w�4�����	c�_�ؗ�`$hgd�z�h����>+Si�o���:��Y�V�&p5��d���a�l�*�rgC�`�u韪�EL$>���Y�.����������{0\F��	ۍ���]<�%T��1�]֞i�Ξj��"�]�=�'���fV���XX�p�h�pϘ�+��k�j��+��9���Zz�ͭ�yN�kp[Ev�:�`~N q�C���S�r56�KV��)c,�E6�e�|]XlxVHYEB     400     150���tڍ7@C�w��N��<��|Sƌ����O�(�R���������",C�/��{|��?�K�_"!���l����6����H�q�N�����I�P�զyۨT��´����ls�KI��/�ߴ#�ffx��[-2�g�,�Ң������ϝ�3u�ghSj!mI��;s�mJ8����瑽�U�)���hNT���J D^Ո~ӕ�eR��@ޒ5p�Ԟ�u6Y��8(���r��n��u/$��Z�Mi.M�h����la
r�J(�zSa^G0쓸:�j�p�nĆh���͕�Ǳ�t�,u�Jr�^�-R�XlxVHYEB     400     1b0��	J i�����GJ9G[j��u���y?�4ZT�	,&Ge�B�	@ø���(��V��L*�_��m�B�]��L�K�u
��I�Q�S�QR����/�a+�D۪��ԏ`/ w�j�_�πl�9o��=�8��6E-"�0�4ˢ~ �!�1Y'%,��%�K豣�2��Q+R���y\���ơ3�1ذE\��Qb~����+bM͓K�|APl�e_@k�8�D_�)�p2�޾�!8A-蕻���r��ҡƫ�-ݩnT
0s��3� �I`"U��}q�ԡ/ ;,��瑙y9���M!��6�/\�{5����۷�ܱ�\��_P���O�L�C��菉�b��xm3V6�{�:�|m�� gwcTk��4<��Y�s���S|�y�{��@PvZX�
0Ѝ��;��*s�>�T����XlxVHYEB     400     1b0׾��l
L]_8I��.�|�H�����8ֳYTe�\&M����p�C�ć��mZc���"�/ο� �M6���_+׮��"�mS$�3%IF��F����)��o�:znC�&p���~�Z�&h�W~���m����7�p�x����Ͱ�7��"��I�����w�.�� �~�9b7���2@Ny���� �Z˔/�p�&����;(/-9\OGUtk?a_-}4O2��+�a���򸪖��ܤj5<�6��,��AZI���$"o���y�p[A�o~c�TYlNj�U���G��qcF�Ė}��
%,�����&�J`T�੓zW����Iv3)�O��{�ܒG"�3�I~���d$n]Q���*�̕��^��l�t�;z��튝9���*E��&'�����������
�.4.�����f̭�����?XlxVHYEB     400     170U[Ւ�����>�{ u%g'oH�2��VD<�h�r@��l�^��|d
��0I���z
�`�1�lg�܋�77����f�V��Ε��γN�����
SR��
~�>�4����uy����M�o��N�qO-���|X~�{��U�/pz�b��YU5ѦUH�^���`�E���Z",~cʸΔ����U�o�px���\�|���Ԫ��%�g���7�P�1���mK��C�#��2u�_g"9"8m3��%��2QC��H����X�j���9�	�F祬�-�^����(���X�?7�7�wD=@�D����a�t�o��1F���F��$�O�B<��կ	������XlxVHYEB     400     1f0y,g��Y�o�ZO����:��i�O����K�:���.�Όf\1=ᇳ���W���v�v�:�c,��.28�^(c�ҺxP-���_)��A�'8m�r{��_	)�IX�����s#����iWeI��S�F���Fs��L�"�Z��>��8H��*Ri��?�^��͕qu����ݝ{̴\�:��ߤ����.\��P_�h<;C4r�lS
�:�D�FN7�o&g���Ҡ'�{z���&����mɤpR`&�x�<�����+��]i=m��E>�L!�,t����R��j���9���T�mÞRy���r�`���2���8�p��J^��pH��h�H����{�	]{�J��b�~�b�)̛�8�I�e���/^cϯ{6r�Ǟ}>�c��1�Z׀z`X귔�H��&���r&ZH�%2M׿I��G"�}�ˊ��z
)ι�8�(��,,{���\�℺�T��7�^>�3Q�Sd@aXlxVHYEB     400     130���Hd��#NM
��d�uqՄ��peŽ�Ry�� ��������R�Eti��G�Ё��vQ���գo����Y'�:����'3�����S8>�x�z��9�衈MKhÑv涚Z�up]�݌�U�}N��U��B7��Q3�!"=%*�H!B�fy`��Ǿ�d�g���ϲ�E�I=r���B��֯$�c�O��;��~�2M��F�8����1�6�QW�5�޾�	I�6�� ^X���U�nչωIN�@p��ۚ�*]=b�����I�@���k�ZڽM�ޱc�g��P7�XlxVHYEB     400     190%P5�X�.@5?���lN�5A�'��fKіg��Djװ����	J��=UJ����NWP�u�&���%�H��2�cW���x�@u���H|YT�ڦj%g��?
��'?�/<h�]��_L|���"y:�^!G
7����GJ|���;A�!G��>eF��<�B?�b�m0���`���`����Q�lY��#DD��Qso��\X霿������Uǿ�%����Q^M������l���}��t�9�-����qH�:X~s�V��V��b晃�������jn�&j|��y3����ї)ãɤ����C��~�/Ό�
���HK��$�}��hh$Ϋc��=�ŵUi[vf1�V�,�{.�����2�i�"?��u��0l� ��v~WE:XlxVHYEB     400     190D0���\�Y���ݴR".�yL���f�[�!~֪���@1�W�r�|����c'Z���9���A2=`9x�~܊	p��E"O߳�`����������ŝu��Lp���ӏ�K��d�
�iy�Bk=v��A��B]K���t2��s;i�A.�/�K�P� ���FD��6<�xoВ�*�F'��p!�Mu�������6%2�����tqfbK;oc7�������Na��7�����\ )�-1[�c(�mN�d�,(I�U~��D�ф�z�0Q
�x��6'O�_<�
���u"$�H�D'F��+����]��o:�oUT[��ډK����Z�G|\Jl������LW:9�u8+�������jS:{:����J}e�BvY���<��5gXlxVHYEB     400     120�O��'��㶵A��E��;Q�I�ZY@�ꒄX�ߟ�q������������"�t�r�%crB�3;'�jm� ,�0P���_q\EW�r� @�	���:.�t~�����*e�G;�+�cư�{8#W�|џR;����^�脂�)�����'�*���bm;C�l�8��$ʎJ��z��M�R�G\�Mkd�W�;�c-z����y��e�&]5����@����Q��c��zZ�b0���b�/�^��j1��9�q��gŭ�i���XW����L�k���M�5�XlxVHYEB     400     170vɇ��� �z�ԏ^�+�^�GV���k�g^�E��ɢ"����$r�,Ǳb��]o�vb���/JOIn��+LJ�YD�n�j~%���_¥��ȼ_�ۥ��s���)�4y���G��C��pJ	�?l �����A�g�ʔNA7��I5GJ�G��]��0-�}	W���?Ϲ�RO3�=y��ϑ�;C��*�&q�(�Kj,AbD	��tS��%#��,�ThB�7�|;�n��^�����3��>���U��׏�w��Yy.�Ӌ��d
�L�s�_��/t�Z��Y�-������gV|����^���Ƹ
��.�.�q{^��'��f����&Y��"=�9����XlxVHYEB     400     170�V �0�RN��4&a�)���(����B�80T�������x�eW;�-t3,�VuJ�H��H��ɩ�����Z�W�W�H��Q7^�{HAZBVÛ���*m�뇩߭���"A�k�z�[�������qt�8(�ᣘ�d�����#�t�|d__�TJ#�d�����jrRD!u����@!8�/�k\��8��rEs5��FMP��2��[�⁢��������6O!I��շD�� ;��߸{�0��K���"I!/����^���-t�[�g?ʩ9�?}���a﬙��V�4A�=Jp}��|��}�1:c�2�Y���zڲ?�('�1��A Xڥ!�g���������0� K�XlxVHYEB     400     180D��*;M�<�M/���q/�]��{�B�@}��F���vy���5�g�l`kvB�"i���~��XR�M��L�@�+�b-��D��)�T�o��Cn&�� ��ہ��U'���b��}!G5�ܞk�m2�X������J7C�G(�S�3{���k5�_�AE	m4��n!Y�I�~����)
����Z�]v�G��g��܈�%E�
f��m�2vFX�iQ �8?l�4s=)�9�آ� (���;�
�uJ�ޙ�F���~��g��t�([��9�?�8�~�S����C��FS��0ܸ_������\FJ̐�gw������:��o#�0CH�.Х " ��b�*/#�|�J_U;U%�zXlxVHYEB     400     100���T�^���Vj̆�8>�8��W�VLҚ�V��n}�#}�b��kԙ���_���(�D���c����t:4'�^���ky�����E�>�F�ݭ��@��ņ�.ʛ��9xA��ߖ^��U��˻���uOy��T��J�����Z.}ܗߖ�ЁMEg{ɖk-ַ�d$��P@�N+׊�l���<�ۄ5y����F��p^�huA~�2��b�r�N7���ft��#hJ�!����~��A��IV�>!XlxVHYEB     400     150(Z�q�����A�zՓ�0N��a���/��doU]/���q�������7`BY�K�D3�1�F@��<���>;�r�~�dȃ�U)�E}q�����v�;��9m$��.rw��1P��Z�����3��A�W��Z�����Q��8����=����m�_���,vv�c�ZMU ��i��#
�Io��+�����8��
,�����U`���a}����k�Km4��36* ��5��	B��9_M}�\��A�y`���s,Y��H���}f �����)|ɞz�o�Ӹp���b$F3���a��%�hM�����$x(XlxVHYEB     400     150`ͷ6�(�7��'B���Dv̰����И�K����M��-}N[�xSH�Lt�1I5�%��MR�6�����a ;��� �Y���3~��N!S�����PA��B�T�ﳴ%��C�x������Tb�b�r�d&s��`�ݞ�zw嚼e�c׵�.�RqT#�K��O��j0Fc���!��j��[����Lѻ��^L���R��5Υj���B�fx���@����;�N�����s�`hI#�cɨ�cc��3��x�)��t����6:�O��9]�\�[g�	��p�D$����02d�ҤN���Rja�-[�!-���s �Oߑ��XlxVHYEB     400     150�3����=�	�_u�Ĺ8B7_���R�����X>N#(;�hD9t��|iA�FL�8�@�x�'��Й���Vg�s>6WJu�61��S=N��ⱔ��;l�6��_��z�aK)����f"&Y�IeH�0%H������jH�mQ�ɲ������M����w���s[9}�^3�J!vy<��)Pc�H��_�
V������O9+?`./F��QB��ߛ���8j�e�)X`�I!�
�}INk��״0�A�Z�WrW����5�@�5"��c��"@��؛�74c����0�b@J��y�|d��;��#`����M���{5�|S��XlxVHYEB     400     180g���9Zj�3�?�#[V+Y�*���#����������Pi�h:,A��a~���/9����Ϟ�W��O��E���ж7���	�|��EJ2���c	<��&�':�T/3h�L#1(uYD�M�t���=�I���O��餦���Tл\/�y� ��R���8����28�з�F��
���A7v�p���ȷ\:�/�u�Nd�%!Q�TG8%��.N��0����YYr�M I�<<���Ɩ�Q�5�3��mU1�ַE�4�s���b�=S-�H==��՝S�9S�6U�����W&���B�HW$�}�ρ�)��E-��y��U�.����ɮg���(���xD���7=���h[!ΟJy���
��j*���
�
s�XlxVHYEB     400     160����Ƌ8]&��3��ϙ�uI�d{�o�3#��!�Y�`!п�6<ۼ
E��p`&�"<�Nm4X�"7��V_�iB�ߪ�}r�V�F��?Qyk�uJ��]��� /���̐[@D��ܫpS�Ux
I�!s�Ȟ�A���pɳ]ƺ7Yt�|_F9\RW��n�nF'q��fG�X���_�T`O{h���!!��� Ab8T�Q����5ߊ}vF�ꂫ�P"ݽ��`;qU(#�1���
UE'k"m���.�V������[���J, �h~k����?�\���wH���\;{��g�2��E�G�o�N�)yn{��M���g��.��XlxVHYEB     400     1a0-<�,(9�"�H�8�Q�.ȧ�Xp��2>�Ep���q/0y��3-�pk"�K֒�	6ʙ&��_���4{�fNRAd��dz�MN�rڈ�Ae7Vw�,���ॻ�"�����-��l�����D��z ��Z�8�|�d��H_���׭�R�CyQ�g���'GLD\8�/�Jd�+S���Qt?�m�r���M������R��*��я|�i��J�.����\��p@�H�����S�ʫI�j����p��gW���(��ƙ�ٓ�m��@�y�A	u�y.Ӯ|�A�"\��79����v�4j�P�g;��k"�Ak��t"�
q�$UCT;��|�l�\��x�6#q�~\!~�jRT݈�С:�*��-T��kp;��CB���'ʝ��g*�2�>�XlxVHYEB     400     1f0u��&�9��v�L�S�~�U����dcpߟr�Cd���
��Y:�k���c;�Cч8�m��YiZ�oc���z��Mʨn!Xns����p�K� -���E�`0�F�5Mq�/�)��e��Q_��H7l�ۈ���R����M8����:+�nu����7OnyO�k����r%�:�߰�c
 �=�.�����ӊ����͜|zb:>����=#�9*�-�Z��*9���-��N�J���0���/Ln�;���+4֤B>+��e&��gt�)��PSV�:��.��o�7��� _˵#�N��+9�{ �C�ekI��S����ǿǆ�,�+V�h�=\_�'yn#�q�6��mfq:Ѫ-@A�2���>�On�JoR�Btn���s��gS�2����w�ͣ88Bߥ�G�K$�����Eb��t����"�������}��%g�����	3R�L��I*��7O[#)�
NW���y �ɐ≠���?�XlxVHYEB     400     140��)���߁�:��'N��F��e�>O��4Z��=|�.{H��269X�\�7�f��3�������������C6JNT��´�i\뉠�Țb{��|_���ܯZ���wʱ=%R��O����wi�q�
��w1�� ����j����e��g���y�.�+��:���e��r$,J��*��s�K4y������!1�\]�������-��`Եw����)�<��@���1���Y���@ ^�/{���V�k���<>���.E@Z�`������G����q�v
�DK�t�K��.��RePtXlxVHYEB     400     140����rR��t?���hm{�ϫD/S�	���X��O��_3�fT��P���)��-p���N�::/n�O��4��L ���$��$| �q�̀`�$C���1�$�[��@>�cϣ�p��$R\ϱZWuU6�Iތ���v`o~�&n�f :�YL:f�3a�=ě�*כ���o�#:�>i���ǵ�i췺��ڏU�8�~`�*�T��Q������R�?�7�bE rˬ�N��ao���]ɢ���v��i� �3�V�Y�O9�� �E���?�!�����vʑe���L�Tn��t
�I�i�zV&�XlxVHYEB     400     1e0�BLN9���j���m����P	�Сc���s�9s'lwL�'9�(<Fm���z	<o�	��M�#m�� 5�Y?=7>~�(�*�i���W%-���)��:������(�NS�X�Ys�/�H��'�4�����-Wk�c���rH(>"fޔA����H8���"��#N��~#л
y(]�s{��?5��~�9TAf� ۻ��?�,eB�:О��I�Q��H]�.w^@�X�l124U�CU���Ć���Pz��Oy^դ"|^R��%e�s{��)�!sJ��щE�d��_������%m��m��1K� �������L�#�[�ܷ��XQ����,�H��gk�s&���i�w�ȫX�QL�w��.�1�Jb��cxkj��+ЀFz��5pۉ��bχy�Hb5@�W�^Yc.���ʴ��u�폒��K
�J�����_����-m����O?����0Lp�ڌ�v�'�I�XlxVHYEB      90      90B��Z=���.�����#R!UX<�ӓ�L�n�`���1�	E>�h����P�pl,�J�\\
A;�@e��/��p	}�bmQ`b6h�}'2��E �LĳC����y�칮�\Rd���z�'��+�Z|�=��~���G���