��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l�������레,��tevGH���P;W�!����������6��cʔ�6d�2*���8��*i$��S2o�U+�����]q�m>*��V�WV��=\��Ë��5��kP���T �i"O�����O	B�O��U��I�]y�Z�.���h'�W��B*�f��c+��fGA�>��rpÌf`(�c@��a$�,���͙p7B�"zx� ���vP��x&u�>���@lI�h��8�[���i�5S������̬��:�E�ҥ��1��o��J����7	�j��C�c�fHw�����k���peA_P�.Hc	����uS�pl�-Ԝ�U8����5'@��3۝C8+3�QW<d�g8�Y�D}Hm*��cw}���*<Ax�7��S��CC$�t�^��be���5�;W����W�x%�r��{�W���Զ�5=��|����� ����,C���Knm��mu7��P�;����@$�(bZK^"f�z�&�9aR�	�Z�[�<ֱ��_�1)����?�kx�� ��4U��>>�H���ly�e2��h�D���O'{�W`U�h�d�vi]n<oeC&��Ce�fE��+ۑi�b�j}�-x:oI�@sP�T���fr�0ѯ>ڄ��_@��{�F�V�8f#���u?a>���*���iA���P�Û�b���XsA3_fq/�zDد�-|��;;+L��`lm�O���_ ��{E��9�a0�2��$�����h ����s�n�7ߙ+>��<�-3�V����ږ؆w�[ /sQty��|=1��E����K��̪�&h������G�De�rċ�Tv�=k�)b��(�ȶ��x�h2�� n��q����p�
wq*S����VؽCQ�0p���U�*<(��
����)��@�phg����<4�b���.+��CT��� u�����A�S��4�)@����l�?�1MtY7_x�j��v�ƶ�$ΚGn�*��G!݉�x��>:Xy���X�Z��,��w4	�*)��X�fJ=�,�:`��r\mN���sa�h�F<*^�@W@�X�&��b;�oި��jC����~�+�t=r��n�ѕ|�/�j-������Txi�6�aW�,#�π��n�����>"H�8j|UN'oU�AD@��Ι��Q`a�Cλ�brH!!��K0y�\���/OG�v��o�vD�LVA���?����#��L#�T�Y M�VEguְzd�]/��3U �lT��%d]���987%e������Ьh�&l���s�N/>^�t����	�pa�t]pE�#F�s�ւ�%�NìTk��7�v�����o��9�~�GAf}�c�Rd���R�a˧��n�r�i�>e�?�k�To��4st�ut���O�g��,.��==���P*f˭ ���պPV�Z��!���=t�⇃ժ6��W��\����h,R�Ą�X]�����&1���\�W�F>�?G�6򁫈���#Z]��񚈻��Q>�<��;��cĠ�����ZQkY0��j(% �M��9�{>!l����̥�H���S�xMw.���%=�����%g�,l�ֆ��W|�Bh��Ȳ�ʥbQc�WoZ�$P��>�=��� ���%�%���{�W���1&��ɿ<��OU� ��+�'nst׼S<>Dm�������DØdg|����e-�@�ϭ=�	�A؂{���[T��/��?t�4��������gaƼ��X�1c���6�E	o��N��|~�Թ8�bH����w��h�}0A�~ܠ�#�9��{�'�%����W�p@�g�Nu�mZ� �.T�L����ݭ��CYٌi��,/Y�e�}!�λ�Z^��7�����K��C�r*��l�	�#��Z�Jۓ�V���-c��]���y���ey~�x��Y�xr=�6�O��y4�uZ���%װ��K~���z�{S���L�����_ꀂwjd#�s$	�H�CP>�S�"���y�Ē�4�n� lR)��VHQ�5�\�����$N�$wuU�/�!���B���<�o�t�8�E���G����U��<ΝN��$scY�Ԝ�rI����?���+O,��ga��2��ڟ^b�w���̰n�k�S��m��0��Q�f}�}��}po)�,��F�W�D{��)_#��s T�ҁ��6�����L�Ȏ��1L�¬�i_�T���1c��@�Y����~�����Z�ح}��מ�q�R�Oݪ-h�f�S��c�巳��*����)� ��'j��_�p�׋k���=Q.�����<��^0y��LPj+�A��^�;��i�3�Nh=j�l0��u�8��pw>xt���e��p��ϧO,��O�3�a�+}����R�j��b����es��K?Wy{�����l�R�V�m齰Gc�Ad烆����EQ=�rc83���BͰ&��$"����1:t���`�$&���}��H�P"�N��|O=<�~.��⺤~����o�ԈG*���i�t����e��$��7PC�1x|s�2w9���1�cT���MC���)i�r;�l�CM�M�����iA�ʴp���-�B'�T\� �vm;k3-|܋��3��_�)�pt�~�C4е����>L��c�8����~	��$��G
rN�_�<�j��q����_32J�a��ڛ8<� �	�ʎa����K�/r��)+��d�#	-���!�:��6tY��f!�Fz��.Hv�l����D�&q�Тw&s�/��v��/�>/!��\' B����s�R��i �0�&�|���^�~�T䚮x�JT�p��|�B8���r+���E�R�8�´z$R#`�g�e!����		��ܸ�:� }w�wQ!�J^F7�a)�\"["�Zm�b����՜ղԹ%�3��劗'G9GP\ ���p� ��/���Э��m������.��	�O�8s��땽�H�c�P2���a���X�t�<}������B�evO8-O�Xd�F��� ǧ�ҵ��X�Q���Zş�Қ�:�-�9�	�$b.�4�=�����<�~T(�Fͷ��.�5��ʗV�S���p�� �@.Wa�κ�'c�Q���p�r� �N@J��1�'f���Hݘ��[6�'9T:q���՚t�K�G�z�U&�;�tZj� ���5��n�N��q:C���5@�wT���O9�� tM�N|Q�T�қ��S�2KR��-��MٌS��S�@��ޏR���n�C�y8�ǖw������*s꜊JS^�����{�h��a`��3���䪬�v�&¼q���ݠ7B����ȭ;�n $�Յ�/��Cn���#u�u�p���\��q=cȯb� ��`�W�(/��Pz�С�4�	�����b?��6���TGuh��}��$Do���{�R���3Bf#�2�ؤ�G_�QR`=�.����L}KP.�5��xx"�=��ޣ��r'��8(��x�6`�=��G�{7|��̊/�j�E�#HZ�(�7�?~B�ңHc�m��:��b�v,����8�ܗ3Fu�X2B�cnW']
�7uH*פ�Ꮭ�o7�I+SOe���7�]G�t�/�w;��x�5ڊ�}?C�]�nN�30Na��|m-�Q|��~N�����yk�!!!�a�H@(F�:e�2�]�3����z�[U?fT�Ii�~&�N�!�:�4����D��씗"
F���� E�l$U��0�vW��|Q�x��-��;��������&6�Y~���2D9D��j����ծ�c��;��]�7ѯ�]\o�N+�eZ'Ԑ����������<�����R<�M���y�
G���R�?�
S����R�`��7sSNE�qD�z;H0uř"4�E��j���xٯ7D�Ꮤbq��M��}��?yUgJ9�,�] L�Q�����.��z�)�n=]X���B=Զkl��
��3:Ҥ\P�h��OB����1�aփU�}�~�)X��v������
�I���]�qnr���ܽ����f��A6@����U�{,����ݿ���6�*܈p5'��G���{-�Cc�vnF�i����~.J�������##�XA����m{c
��$�B�g��Y�P��iW<�!�:�������D(�".v۬���ޔ[=z��D��|\)�%��ڻ�}z���_�W��L�֬��C����,�O���.�,��ꥳn.zD#ڝ�Ts*�h�᦮ڛof���"+��to+�{2��3�,��h1OO$Y;��nƬk>���xl�9WJ��8T@�-!:N���p�Hky%���Ƞm���d�/c���[�i߅���E؃�A�śHua7F��1B2�9쿎���+Ca:��Jm��N��� �u�-jA4I5�R΀���@~h/�(Ɠ7u�YR]s(J?����W�󾄸0/���4	Ϯk܊MY��~��M(@�R�;��T�zG]����.x��,H��}Jm����=ֶ�`I$Ή���a���NG�K�F��B�0`vF(>�P�Rd,I^Y�@�'(0��w���X��C62�,v�B��=�=��6q �UǄ�Zt�#0��F�y���^"�u඲�4�-�	�6��1c�(�6�>/#��a'�7Wi���Y�
�2��DJE@:%�;<�b���מ`����o� ă�V�U���qڝZ#�ϫ��G�wP��W��6L�� ��j����o3~�M���V��5w�/��)�� `���R�J���W.AMd/JX�R1�[)>Qk<���� 9�Tf�Q\v`��E����Sf8�P~��+��4n�l��yI|�1��j�Ŕ�<x�S10�#��G���uӐ8GƐ�i�&�l��3��/g{w}^w[;Z����� ������(�)#qh��k���\��m���&4,%@����9)d�zBa1�N68�Xy���WK�5-�.��� ,߸Q�*.�� ώ�n#s��KL7s�)��$=@���_�:��,��(�r�y��ܓ�5�X��$O�d!�h?/�`�@�rO"�����z"#b�m9����?��ej]�tf�v[� hbG��	��3oz�p*1.o�[�B�W|�n���ik/�õ�۩�+���<������w���t���8EyD��.QEؓz�����;��������F@�i���{)2��UU\��{�\�Y�m���I��~.��/���Ť�rx�MM���[�t7�9��[J�]���?�����~�R�J1KZ
�'���2��%mqXզ�z\�*��k\2�!�Hh~�����\����)��ȅ���F创��ɍ#����k��ӷ���Xp���lg-{�L^�i�.���7��Z*ko1	A��l��S0*w=[t�g�pe(�=O���GJ0g�(�?�L�n@��=��Uh��u_}إ�%�Z��9���B�3��E"�1�YދF�����H�w8�p�G��m�;�����%�&�T����r]��&�I�~��=D���D�A����2��ºْ:A�펒M�ء��ּ���)-���o� b7��4��,_(>T��� Yq�w`]�*D������Έv"�bt�t0��U�2Au�|g�X c��/|d�d\4��N}�g4�[��҃K��j�����_�����w�*��g�̣t��@�TO{��u�'p�"+9��i��$���������T�%a!~�S��ђ�a�k`����S�zAr� ������l߰=rP/`��E]�誌/�<��q&���i~r�qn���\T�T�[>l� �X�Yw��AD� �P�.(�+�V�VkG7]�����d	��>i�����^�r�N��:6�؇S��	Ki��
�1~8<�zN�<�q�c����$;󹖇-\��ǸhUq��߆�^Z��!Jj����U&��0I̶�zF���oYmjכ��ʌ?˽W;�G�?ٝ/x?q7G��}�w���x��]��;����3bj�>�H�z���A��N
l��F���՘@��3��CvB{6������ٵ�}��FA^W��г"�Q���ϥ�j�9��4�l�T��X	��s�M��<�N��xV�w΋b"�8��f�Cv<��;�a�zC��|�9�O/Nx��H�a^�l��d]�<�%�q09�<�����<�A�쾱�P~t��$�\����)��]ԕ�Ѡ��`;},���w��ĥ� �.��ފ�_�D�)np���J:��n��=���F���a22\jA�b޺6r:2����_5�E(b�V��6�jJ:�oUҍ��x�o�'ߞb��{�ҙkk��ck�J�l?�����Z��(5�p�m�RF�g��x�#����p�@r���NSr���e��iȉ�0�˧��JE��Ӓ/l�8Jܱ��I���%���ƛ���JJ��Զs�Bl!��a�"�X��5�!��g	��#�i%�M�p�^�bcn
Qg0gB+1F����)�C�!"�:G�F2��i�[��:K����GԿ�Hl�}tgq�nT��ہ� ���8Q�߰����3}��� �]��.����BD�$Z']��U��E��j���uc�HS��	��p:��`-k�9V�JFJh��RSN*�����)����R�(��\R0����**����|��x(;�N�iv�sM��Z�X2x�+�lo�8� ,�	+:�
jNE�,���p���
�J���܃`�����OɔK�#�0�ϸĒM%��{���������D �A؃>�T�P��
t� ߻B5l߭��K��qetj�t*��C=̛�נ4�:9]�nP��)��75��3��J킰 �$�MY��Pi#/ ���0�i�}	\�^n��1X%�ikc��S8�����t�iD��VW�����J8��L�c0�,f�[a��妄	�'r#t�q�L��uB�M0tCo�V4䩹��w:6�:�^���?��C'�oɝ�W��+�b�u��R�w�Ӂ��%�U%w��R˝�r�)#/ᘬ�d�xT?�%'��Q�`UrXٛ�T�Hi['�ޱ}~������2�%�B���>NM��]`v(��ķiKn���_j:Q�I�<9�2;�K!��-�`o 3�irP�T;��|�J>c��f�����k����Y{%Ҽ�n;Y
$��+�NJCq8�6�+
�k�(��Iw�EJ��o����'�~����mN��T����^qmN����Al��:B��_�����
�ֿe@�,����Y�uP��R�X�� ��]�(�ks:,/t��*h���W��(��G���+XI_�q;�
���\���x��V�d���=������n'�EH�3�g�;3s��`[�w�V���vd�� �D�6$1��H�t����"D��"�|�;�W�xt3p=�L8>���3N �y�s��$Y�Fjl���([�+7�w�p�G���4�����a�r=ld�yr�����Nn��}L�^[��/:��[���A�rOi.[��m�<����<M���ED;��� >mʆ��W ���@�OM}[ڒ����D\��h�,�K�fU���HڳBu������F��;��E�(U�`?}ͩJ�$Xw�͡l4�i���ٙ�\N@#v�~Bbt�~�J�w����	��7��{-�^>���04�`�o��7��N7���Ј�U��5]�s�SO��d�s�F@A����v���ҮN:�5Q��� ؼ�|�~:�@����+07!���
�;�E���l^ZJ}QC���b�:�qm�p0��q��7-o;�)L�gR>	��TSc��KX�f#8��NbW@sF��JQ[Ja��q)(�$��
C	����`G�ɀ��e&~y�����G#��)ٰ	������4�%�n'���?+�B>x���\�͐�8�V=����S��ȫIHv�_&��r�"XaESޯ���!4itb*8��?!g�^?�`r9f�e[�(f֜qz������'m>�2">�SՃ��~'���T��-�P��cSv���A }��I�o/Ɂ�
��p�D���Q�'YG9��X��ǽjgn�!�/�7k���򆞅)�[�4���w<���E�{��>��1 �ut� �:��L2Y(	s��'��nh�ş|�b�B�m*�W�wϊO ���NJ���L��V���bȆD� [�8�Ȑ:)���)�j#��>��;�k��F�s`P[п�p0H$]Ny�~V��K��e�⪖�z�Z��k̬q�H^���K��Ը�L�xzw*@������I�UZP�:�q�!�h9a���XjclV��7��$Qrg$L��1h�.�;���ѝs�[] �k�S�����͓�8���P9�$
����u'��x<\��� +�&�%�6��r"��'�����c�ӃV%���Q�!qZj��soH��yN�\M!&2kkb�m��c�����(�@�{1�\�߀=����S��ڹi5v��o��D"�4C	j��_����5S����6kV3�	�RV��e�6��!�Ŕ�z��|�"IT�&��8S��^�l�W�hư��{0G� �!�b�v���0�K��&Xޝ��&s��A���#�p�P~�M�U���ϨA40l�~g�Q��}��,��3*�2��9����n׷�3Ѱ��%�*B5?"�`IJ�]��5��\�Zްv)�3K��0��gBn9&��һ{#�����T�������uܹ���� �-��v���W�ɝkO<=:��q�9G�Egh�V����� �a��B�x�����g"�<L!����PZ�yK{ۥZ���g�M,�X>vm�#���Dwv�|��a�4j�6��16�5�d��JW�0���&E��Ӧ|�r�O/P2n%3;_�X0-6�8q_)�M$۬�S�&�=�:�_�!0�$� �4W-�HaT�]�OS?{�Bi��n*~\K�*3f��Ɍ���~w$Q��K�,$���z���"{���lk6�ȇ	��Stg���a�D��f�z����A�f.��8iB�Td�W�u�M��Q�q�{X�(�e#�F��x� �Yo�G����pk
�o,�aʶ�v�����~���Bx���j(�m3�G{~���7�k��y����+z;3l��S�i��7��xH����'�������9v�,LQ��H��BrP��r��
x���<���^���.Є��fJ���!�q�;����M#��]�#���j��g*ċ��4C�P������4G��;��&�L��

��u�:��������0���2��f��k6i�1C
����혨kA2%Y�J�̉�e�9�B�ژ#��\cY�B�2SS�=����Z����������ss�pYT�6!2[�FV��rT�V:9�������9�ˬ��u��'�/F	�yK����SZ>�@�4�˿�X���Ż@����T������G&Ka}k!!$�-]�/��bh�6���N-n�)�\�M��l��6��%�h��+�٦�6��7��N*0{��Bc�i�L	}Ϭl~��n�9%zX4ia�`��0�Xg^[���^(7��-�љ8�u�ҡ�]~������p�*u#Z����*�����of�$���|4�����!+�s|�������:�F20�RC&��?]JGO�x���b n7�uZ������ޱ0�(j��xi�n�&E���r�f&�e�!�	5��{qo��Sa��<&���ֱO[LN��eQ
Sn�FĴ���Hs�a�d�6a�mp���(�݉$-i���Z������K��L���Z�P2>�du��F���2[~@�q�az�oT�ȻqJi������p���lo��6�LN��q;�ڃ�D���1�/����JtV�a�C/ �be�
is]h�}6'���/�!���ʴ�Sݬ��qpK�wݼ��"Q�f�	����x�T$g�������6Dߍ�������p�)H�?��1��,M29�x������t�ՄZ�s�C3W��vա�h�6�ԯą���'���)<ΧV�І3}�7d�f�N��#gb��D%=�J䗿$�@��m:����_��.A/��ۗ�$\=n��A�o(�y��Q��o�flXB��x�>.��[ZD cq@�j�$	��o�,/N�E+V��B�c�����ʼ�joe%ZrX=���3cq][J����B�@ܢЄe�$�:sż&�h��~�$P����H�)��QA{4���.@'��f|_.)�a���%�ZcpZ��lQ�6�	��M��D
�}!@(��o��R:g���} f��wL��"�g;G���H�D�T^`	���r�K��T�q�n�"���z~�Б	�XƔ��.4��N����7����2QT�6r���K�]W�2uZ`�LB4q̛����'�iD����c�C��C
8{tO���*B�����Y�'��k����4?�i��)ݙ�,:�N��Ұ&�{ec�@z+�p���'���p�����7s�0���g(]�v@�A����J�-?�#����`�y�Bw��x�	�8�|�;��a�Lb��͈��O��4�^����Qx�5&��<0�>wYͲ95Q�Y�F^�o&v	6�y���,nc�KAh{�Wp.��)�&����,y�i�7?��A-X��Z�yV�A@Lo��h��e0�t�y�ŭ��a.t�'��d_�&z6r���
TĪ��y�O��#�E;�J�bIĤi�f�T���