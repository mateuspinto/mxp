��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���?�;ENU��ڽ�/ı��Hb޼��~H��.�d�g��vo�D��/���d"�|it`�N]x
D]ܠٜ�:t62�<e��&�^y�P	D�~f|���}��B�����HAF[��t]-�6��p!��i��l��uSbAƕ}'�T&$[Q��u����C+#� jJ�P���k&2I�8��3h)���p���6ڞʞ���C�<H�`�`т6�.Xħ�����y�`zG��V�bÓ��]�Dt�W���0��=�����2b�m\7tI�v���=Z���G�zj��g�e�t
!P q�ޜ5;��r�S�O��"�d:�2��﫩
��(�8܉��Br�~
il�Ha��KB�m�ZW�s@�vX�z4*���<~��R }��ڪ�e}�ѐ��OU4��R����NJ2��Y�
d��Q�!�d����6���O��(Cy�c��ⰷ�_:և���t�u���V�/�Su�,p���.g�	`�?�� �1�Ĉ��l��5دQ�M�!Hq{�fBe����͖P!���aX���sD鯠�h*
��*:����a�MH����a$$����1�8&�!�=,���X��uE�}re�<�C���"��~�n�e���O�dq�\���0�8�y�����VC�l(oZ[|	�
k��s(�7���}sW-u����
QA%^u�wBK����l�� ��?P�r}�^Z[�u[���b���/Z�
��,��`h�-��
�m���_��
'�M�O�k׏+e�ӱ�t�l�%�y��9��sJ<�"�e�\!�O����o��?����9���
qT~_9�~.$�OƝ�`�7`�<����&tM��} -�x&T����t��)�[V��b2�ڔ�*F�����f(ƅ;(�ߎ���l�.t���:��	��N��i��K0�����H暍=���a��G�Qߒ�Q��J�2b%|m��@���"ܼ�Z�S�V�9��_�xr�|q�8���en@au� j�e%j��G������u;Zy礝n��7r/O)x�MJ	t��F�/�O���	*-r�X��kdX����:�������ƝI�_�r��)飳�7O���7{iJ�WJ7�L$��3,��sW�}�\Mkbk�@�4�FǂGA۽D�C"�I����� T	oe�����3X)����]fP��ʩ�\%����d�a|6�rEM��a��_���� ��K�y9�pT~���h�G��ۼ�$RH�)��$՟G�'fD/)_{�Q��G��a�ZuE$�CtNM>œ�cC($� ��M(��&��(^���sĺ�8���9փG�ɤU�QNrY޲?h!����n��?���
��4�� ,�#��xBKۯz[(��:�ŷ��
j�rUџ�'��F��ʮ㲥�p�3b� �	s��1�棉/��\2˰Lᠣ�T	�?��\�)���p |�%�6�%�a	ʚYm��#`�/!��jm�9�nM�u<~Ep�풱�\:I�[�w��l��Z;�3�L�f�oD�sm�R��'q}��RO�F�`�!+C��T���;Wlj<�w�Oia�~�S�����J��],�����!s(��|���J��e��P/g�^4��&P}��� _m�U����Ȥ�L� ���5��J�t��l.:�m���w��_�/��r@ȕE�ރ�����=ɵ� %�J�f�
�Ӣ����^gm~&W}��+�Į�\�1@���T�͌��2A\3G��"����d����̹fP�gS����3�:�W.@�v���d}��� _���JOg@<jY��{�N��_U�힕u���y1ΦH.X�d鳛Wi�A<)����?�R����TI�TZ�����	�%z�~�^y���=�cO֜��?���shgpj��*�k�\�a�{�D�;����%����x�1U�� `�^��\ ���2�+.�л��ꥒ�ׁՄBo�z9+�f�)s�/�1�Lg�GN����V'��l9�9� ���͊�8�j�E����!�y��Lغ}��cW�6w!+��5��s�
Z;��W��X������ƧٺP����D�6V�%�a��ls�Av.Vδ�n@���9l�d��<�k�s�Υڂ�,�3Y����n��"��?T��I�Ӛ���ģ_�'��]ƥ���⤄ ¿�q����N�?4xU�ͷA�r�p_mP' M���	��		�^4NN��ܡ&r43�W���۝�Gbx����a���:EZ�L���5E�0����4r�۰hR�7y�(���/Rt���0���F�
>Gy�n��Q�/��jT=Ж(�P148E����4	b��ͺ#�f6̸��^�XH