XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��o 4Z�*U�Q���#^� �Z��2��YB�NY�W0y��S�@*}f�C��#/?���y�i��"&�ݡ�#�q�.�b�NJ�}�V�1��d_�Fg�Y�ُ���ʁ}"^���.�dq7��&	{��~�I�Qj;A,������yi/��~��1�(}�T[�}����`1^OS �=	�m!��d�ᲡY��I+p�.�~lB��^ ��f�Y�C��`��ݢJ��f�Jv�7ٽy�%�g��ܹ|��d'�߭�����#��C|^���]��۽^V��>������]�
]��������n|�����ڳKOP^�_5<�`�%8$FQq��o��v��\�}�춍� �v�Bք�8|R��!����cG.��	�x�YZ�X��a�&����A�z�c�����V&A��̘:�U #xS�؝2VZ�c���K��}x&�B�uػx	��p4���o��EO������gߚ'�P/L�ko�ԃ	��:��Ac��W��{��uZ�*/�8�C,y�n��
�W��|���񷿂�(ƭm�ai�_��g����0)�ؐA'K{��i�ٲ17	�����%Ǣ`��ƭ*��#� �|�7���!/�1aY�[* �P����쩂�>d��at��4f�
����}FI�a�����=͎��o���ך4��jы�%%�@e~(�O�,'�8��D���F�_]�ßt
SE�p�lvf���)0�Q��M�l�i�7Z%WSe��`u��XlxVHYEB     400     1f0�"
j�m��96�d�e�n��4����N�A>����#�|�PidÁ.�9
?ىv�U�MOt���Zɏ+��b'�O�~I��|6��o{l�qG%P�'�+L����Cք/�36��_��t���1a9�z�X�L ��~��)��R�K��3Id��'���B����R<\/Z� ��'U6z���&��B@v� ��p��cl�,�}�U��.1�F)S[���%:��\��kח��O��b��Y�ƃ�#�5�Ѓ�F�"��P���^�>��2u�Gĸ~�:Y������i~�
���'�f�jBʝ 6qss��$�L���OZR��C�xf+��N�KL�~"qR]ާj���Z���k!9�ql,�:����=<Z�"N��2v�t���E�G��Hc5V]�l7��&jjsO#٦�T߂��qa[3X�eMf*�#|�&ӄ�g;�i��E�X;�O�~�Nz���P���
�_ߌXlxVHYEB     400     130�J��[�v�VBq^��{/�@�@������gdQ	�^+�����'Š�e'�Vq�!��ܧ��՗�y�;Rhl��)ޢ��h����&�ꁾl*�^�o	߮5��Zr�=9��$"�F�uT@�*E:�嶪��f
hq���;�\2�&�'�Z�Xg����TO�-F�Y3�/ui�X�������}oYv��I��>ؤǱ�~��/���y6c�������7�%���}��/x����W��?`x����*,P!��.7ߝ(P��a0���yгo����ʚ%y٬�`N��;��mXlxVHYEB     400     120+��>��ko��͉R��0�)�f����]�4a{gE�2u;��'��������v�Yn,����Ud�CR�eKdP��l>\3%��x"7sͮ���n��Y��`I��0����'��ȡ��W!eoȴ��\�=��C�Hr�,g�P������0Q������<&��>��-!�G?aT����8Wu
�ܯ<�;c������C1ř��O1S)��-���#���GG� ���S�"D+B%4AxB�����ƤL�s�H�����-)" %�	g��m�lK�:XlxVHYEB     400     130�t�Y�������kN���#��=K�l�6{��#��6c�O�	��f#:�d�J�d>O�v�s�B�(�Ԗ�W{�c�0��V�z���@^�� ��T�%�Ta� �n$�R'OR$��̍�1����h�M�=�q	t��>]c���a���|�z����HB���v6Zb+8P�*���Ќ�&ɰ-���3X�׹���v��t��qS����CJ�o�3\�s�:	��1moP7[~� �]W���=ٵ��)Y\�e�`����!��ծ'���Bs�\o�������s�XlxVHYEB     400     140s˲��sQ)m�/��)N��`jR��X,X4�$�J�o-`z��<I5��;S\��lJ�u ��s��Sr�5~G��{�}Ȏ���p'�xL`%j�.�O�Z�ޭ��~g��W�
��[	�{��]�g��D����7{.�D$6�:��6'nK`%>Fآ�.d_�F8ò������}B.��r7f����_[K0QE�n~b
�8��*jZ�X��h�2���O	^fJ����U���L"�]uY��\h��ɟ�jD�.����\�'��|�º���98<���zL۟��|b[5Х�tX9&�~l�t����ӗ�XlxVHYEB     400     180��tH����
$\SD	2�O,���O�WV��oD� �WA�Q��(�w�>��r�+Ҁ�&�,�j�`�F7�& �O݋B��� .I�� ����X��@B3o��?g�Y�#
�ϱ��0ěX�><��?od����H��:$s��P"�ń��eEI�j|��5T�ND�9����9ִ�V���}��-=<,�D3T��d�lG#:V� 2�e�$�Uֺ��;u��}��xѩ%���a�f��Egd���u�"X�,eP0����/7�I��{���WD���7�%�	sq����D�8ђn����4\=)x�+�6U13}�h���_V�]f��v�'��1�y�٩��-�V�2E ��Dn�S�(��x�L�����~%XlxVHYEB     400      f0��U����������qr���K3�[�Ȑ{i�BU(	I������]a	5�Ƞͨ����}����?�UJ�}��o�n3�A�EL�M���-;���Mk�	�d��(�Ӫ��]� �fR�)��G�,�qMS��� ^�Շp�P��`c��#Q�&AI'���:��K��.��H*�qZ��.
����۲+���Ak���~4�O%	�]4�z�	��[��_l>���3cXlxVHYEB     400     150�%��4B��~Mg��>'[A�a�Œ�L�&��Pu�)J�Kx�k���+�{P������X�˔ x���� ՟��P�~#�����4����[�U��7����p��+_Q���%u���q��i���O4��^2Cz��Cvq7��^!��d�
�p�x<Ŭ8�r�8h�ԅ-���pA	zl�����24��t��%bM��W����Ѝ���k����284��Iu9����X�ЇdwQ�u|�b$6"+�*{Pd� ��K?|i�J̝*L��Lk�/;���"^��f�|Nk"^�៟p��%ge�-�ɵt���)52j���Y��`nV���NXlxVHYEB      b5      70���Ⱥ�x��3���y9����b��2t���G��4�N)@oJ�žn�7��~`@����@�������K��?;ph;�n�+����Ŗ�է2Ї�<[��1���d#,�I