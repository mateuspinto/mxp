`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
SmbuuegPi8e+4xmohtUS8RiE/xH2lKPy76RR754MOUjezFXBZd6R08WLVwotjS1aL4ck7BdZaEUX
c/NZ1+2K3BF3gl99JRBPHAKIgl9sJwb6MDZchIF1zYAAhEQaXJ2UT8gqF4jZoIvEVkoCISaWbZGZ
nYn4Xn/pWYJAcLX0Rse6t7jRA7Dva2/X16QgLxDd6mRogknRoiLz0xdy0jCv3Nkrb2ZBelvGQHIm
yDmdilq2XXuoTmgOQi3WCxX9WjcqvDazI2GSYPAFMYjlkTHIrz9fQWmt8LloWdpU6t2xV9X0BWxy
ysdlwpVWCIyZpG/Ti/1yu0iMxo8c5OWevaiTiQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="UZAYjDr1/noODYE9hUZDyu/kSjapD2neXhmkbhv3+WU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 94592)
`protect data_block
4/Nu0h3WRJKZBN/V4c+ZxPJ3nVss/tks7f7Fi0k+t9TmIzT9Sl/MukK7Qb7CPAAMVan6WIDMLCol
D7BvXAvE1KM1NOpUDtkP8pdBImBpZy9EEammweo3NDMw9iX9EmocoQ0llB2Bdbe2mS9Hor3aePFw
VlRcB6t7RtImnqxp+mGbGjHHQSio6CslEmWEsRQAiq1ukzhrQXXoFASeGbGWNunlyWEM1cRLcqpI
t22+iIQ1f+EKFG0GHfRCKk3DOY2f+GxszGnJFwKwJmpOZ640x47B8Mu9F44W+MP2/nyFj0bpP9OE
Z6tEosYeuwC+VoHuWH/FTSVsQ5BKsJma+UbZ8ByIDNQpz4PCIuXv6xIoNuwGKFhe8W3xk38Te76z
DWxVx06FjakU/UlSHFo0k8BdTqx34kQnA0+9q72eZMg7pQlmui4Jd2GDU/za7TpNTOxP6CUJkqt9
LIXtLuBV1GcP8ytjIoBBGo5QYFbq0zk5gufzaFZmsP/kukTxzEz6aZKzCP1V9e6+dbEEGg0GLrVF
+ktCvJm1mY82v222b6rnhsCfGfmAer5Lvmhc8x+DBKQP4DSb2zSZgb80Yo6HfXWllc99uYE1NVw6
K4XKbsUicfj7ggizHhCUocI0S3ty44OWYjhfwByb7retf+DgkXtI8vWeeZ3BFYZf25fVpRdC/DoF
bBgP30fy70sMLqBTKT8fgmWIR+hN4uhhNvqf0+KInP7XiFfpvhB3l+p5kuoymyJijnongKlW7Adm
DJ5BWS+EbBDE/KbfaTMxMbLmkOGNp5puQ+LfDHdSXwj9O4oViw04V/3GEQGEOQIUx7hBVjGRY6jU
ra+pl6UYMC5L6BRfYqP9mFlxD6OwiNR3n7bDfA67pRY7OAqpp8eH0v7NYNw4ZlMk+qFHM7kG85Pk
JJ+j8XHIg0ncpMsJTf3lsJkzOALO2W/e0mywQHapZV7KIEJmkvfE+G5FyLqEelouvG85oK55X4Yy
4NZ6dV4w0G0ouPWG6lsNfs2yaREUb6gpmMYHHmbeS5NBSEw75qevJnQuwvzD1JAlS+lcbu2l+Oes
UdccAt8uMk2DadmUw0D5iDkzgRpRvdw6lZxPFGFi7ypc0NMyKnh9Fa8/Qu1LqHGyfnKH92zAO0kr
EeYeppjqUmuZhvsbD5irm3faLGgPigN2txz5CkeC+uZF50GYo3MD0KiiZJJEgqfgWLY4zQ+/PxGd
F2kR6cRx2egeXxE5WSzG6i1QvTc1swPDul+a4XlEbE8EK89X9yM8vu6HDZj0QH9e8P7d0nXDeUS4
QiwRiyZ3AJdqZ3IBoGNoxWWBxomd5rAZbNq9gg+sqYCIbWqHMEreMXwMZO5v9m1ilCpQqaWBSP4h
OHNgVL+w0lJFHMvHKJVBItJxk4RhvOdM+srEgT7t1c8EmqgacHNiR9D/8NhCYw40NYR8DW710Wbv
L4OUl0dJDIDekgTLrGxPpvpCtXqEhRcMhrxxDQlvyaTwevU2twseI7ZFIE5LbFAzCyGbto4oIiI3
jLAN57Op+A9hBxi9dwvpg5KmuCnYnjq3XJLFSFgZcxXX3/I04PUSacpncQptGOttkN1XR9jYaMLZ
du8mFuy3tXC4KBVt/GZHsDuhVpUK2yVW2/AvjN7Ec4+mhyHfqORj9Z2qNNeErnjQFcNLGparCITb
2lFM8VYpFak655/xJXNgY3SBA6UWvOlyzHkbpiwakozLn/9fmMF5qQwwqPoMQp8AGq+eqY/bgOjW
ZRhX2QDt+lDwrzxVm859KiDnPtFonMo/1uxsjUyztFgRF8bqTRB9HGT5CY29AbmSWsUJVUUWP2xE
KHERr7m/5E3gGJiNbbDVXQzKUdmQsSRsxypOySW4eDg3Q4YVYy8EIqOPvZ3srLDZlkDiYwzapbOr
wTh9L56tGB+XJ1ehQakal1+8uFMSQNkKBYiQXS/MPIiirZoDD3fPE9chhuR8/wK6SgNkND/G90C1
bZQbWX8YwXWmet7HCrhgVHyzIZt+7z8+UPRKYAi1JmzEj4Z7zjprdsLTa7onCH5z6oUM/vSfwy6j
/24Skwbwo+Yjrzthy+xlAWjLR5Uv2InHPf4Z2DVSEnIa8/Xo7rkhAFFJI4O85MNt5udXksmqy1bU
L4JgaDTzYfww6QVduq5SoS49Pjkz43PHSmax2dwApC9TkU8E97kOulqOGb+d7Zg1LGtIMN13ilKB
A/7Rt/sCPqXR35UIwmzopu3+9su6GgocV5fcnfb2Sc+U2jwvU7RJTmDZJRW6K9MTJR21nkTkP624
aFGvJEBruYq8WW8nLjvvE0XqwP/R7oKhPweqPMFVUyA5mzDnqt4kHNu1HWRULj3PjKVA5/LOtpcg
sFyTjHKLG/64G2EpqFTX7/mIClh2+abWprztydq//mTmU+8LgToD6VRqA8IQpx4YOqkr1dZO8mGh
SdD2LD6m0BBhGd0CNTqKERaTefJ6hsOiOtRCSeSJjKfSg0HEdQ3unlI0swDsHRMVlFwUs8zcIr9s
sSFDibuYPM+STiNPAsVc1IPQN4RFYHm698BUXu3mbqNZy2CKchjhBd657AsqSlRkrtICCbQbbEX7
cFCCg1WaPDzfSQrpgqX/ynGufQi94qjuFQvgFKRLvPMq0fg148gBcvaHbvvYty4QUiGZFfgOsWSq
JQTLfNnm4oUuQl2afKoo9AXQ/g7L1pQufhTmDqsG84EI8veY0Mt+fTX0Mpv/OHGaDfW52xdHmVXR
HWyPlkkWSWMfNrLpDCU1zF5I5/xmhZ/hy2kYRs4oz+OpYv56YwYQf+Y3XxDkR3RoXHJpefN/PMAe
HPwQ1ZdKWP/JQFW+VSHN2U3HrkRE3Wa7d6oC2d9loHKU45dtwFshEeuYVKk9nvcne85GCBlriwi7
7q+IpHtOV4AMe61miWBw6B81wNQ8ZMrhE0rcgOqR/n0TDGwl17ycLHAUaKqVpV6JSotCIrTwG9h4
r4J8BEXpcW0JCfDofOm+FfY2C4go93gUiwT9gsfTnUD7OWBTckgmS0X9RhdVmlYQUPy+FWMq0Fkf
Rzp4O0L82Y5GJwe1BoJM0O+RXX+BulgLf/rcfm7qKC6jp9yHjGHst3kExmjDQTHzBadXhiMGhdY4
Fiz1GT2SQQoOSMsYbEGLTqXgRq+LXqAdYR5q5ff7FNuQ6eGIUNk5+f95mw6RwfVFCthF5vdO2frK
Sl8bprH6JqFvvIdsfqcYUM6idWKWCN8OMggIi+sXYYS8h9puRPkuVM54A+4uMzuYLHT2Zk6CV3Wz
u+LuwT9ajxGkWZoTqrQq5fUaAhta4g08N3j0T0s5LqhPySOiUbOcxF8yC5c8uDgnyuFBbT4QVJQM
qOr2BpqReI4AEW7ihWnBUDAxw+i/b+XgwM3tO4nBUx+1Aaugj8mFGeKpuZrAfTjObj/3dAqCcaYv
G9+8g1QvsQ0dXAFHlhoDvPxEtoADnXGXU+gfLfs/KuCFHzYjhSzLodtiAQuHXNv920eVLFu9jf7p
UJJ1lfP9O2rTNVZY43PHKEJEjVCspe3Lhc5GYWUDPViHtvzPMrUysCdlWN8MUi3i5IzxX5674Aew
h7Kz/FO/DGLrATJ9nDseK5AF0QwVb+DPJ5EJPBiYpJPWexOHI47STL1J4l26zFqxlfA7JLajpgvW
mhCfygk6AqoZCyr6P64W6h5jHDdyP1Suh56MGgORygovVFZmZLunn1zGBokVVfL2eKEyE+oJT7Eh
KqxBf7owfZgbjCz95sbHaCRoQ29uTh7hUC0u10uym5Cy2UwdJjskBrX1vAdhTQ8XojWAL7Mu2FB8
Y/uij702YnZTuvWx/4AErA1aOXNJOBRwC3ksKwvOv85n5tGUlS6/PSgBR5uVNYR/YWVSE/YC53WA
TlvC/lUQLe+RlOdv2SJ6eAPfaAUX0nQY+Y98n6bKP17R4E+kWbwuqHloqXRIBrI/O/w8ZUe3R0LK
Xc67Ig2TSEaYCkhOzoS+BasY7xoGzaAHRXH5T8kyIC4DFBo1ZsXvCr5I7MAXL+wQkZ6WHM8arXan
hhOfjRs3twDtDd20nOLyUFzKm9mIJ/sVym6iDhoYMGonmr3DvGLWUAfEJ+gLtqixqb+U4RwFqdnL
O5uvVLhnfiTyA089/zQZsuH2ajuEeV++QPkbbmOo3gr1//smVsm7PnzC1BxU+WlBfGCYb/AJsy2C
VF6wAAyEQYIYKx9J7k5liSHMZwyrw3gUpiyaIc4lE3UivwMTvQekL2OtTTzcb/G4J0IPeJvp65Yx
l+xl4v7Wd+WhKwL4nQm8Wj991uIj8icrvp/oXxwN0NoEHi9PhxaGWZe79sxN6vAO+ELA2JWSl/jP
jCwT4VgnTUmdXp0RUvC6/qQxtjIgYq1CEa/qRWOhL8SUUODaG7oazuPd/7/GsYaBrWpBcfdC4gW/
H6MCcm8ZLpKFiHhHMYcthAYzKW2S0i1dRLECPOcMu5JU/iu0zGc6RWQ1x0WPdqaPAUpq2HATCoPj
coW4KrfdjOrxiVe5a3q8emmaUIZt3beE9RKVCJRXwN5+E/rFM315U5iXYNtcec1BWgGCKWswUcES
67kWVPRx2hNTj/QzLfNBFWdhEfaRo5vSwxrAQouXjga9rrqdh/A+7d+u5JhwO4QP9IsgIt/rlbBJ
XABKQzaVUSekfkp+O2BD8EU8UmZekpoEuk0cXkDJpYnsfF4MqgVB0my7D2NaB8mk1dorL1Y/IK32
Rl6UGQrGQ2UjOo1xsBEMDV9KFLLdhFAzgSUD8KbMtzk11MoKiORAhVpch5l95mtycjvK+racASwO
GAnQuO6BkC4HOsUpv8Ocnq4MaYcVYRD4Tkxmw4+/R72RteeDGHYY8Oe8PI4KJxL3bqa2t1x3iMWo
Elax0O5QQ7TnRt/h3D+t/JsfMTLzaiElnBa4ZUgWybp4MWJ0otV+NJllv97tNj2kkuFrOkd23NEL
846Dy75jRu4krVzEOS8MemLkZq/ELRGKVAzE+Z5UxBIwuHAjVeRUwzhSTltB/2vkJUfWIuAra2Di
+QKChioJnCc806il1AKO9b8Gt9TGAM4X22hZk6r6DFp+FhxJnAoN0e3z+/NqXb3tFua1cyjuCUPv
K0mS+kb/cpKNldJsIJD3N219DhcjZ9S4rgay2J4MybVy/Mj39bg+7gSsOyUjF7WFa2LJd2XlA6er
2b/RYd/7sbfPuS36b4Xena2H8m1CFXi81itJwMSV2UBtWcWlR0ZtfdHU2qfmWSzr0Z+RRLO4ClVS
uxhgoOzajtKxINfFPVP+QRl19W2cjKt9tQ2Cz1xzBphJ7aV295KUqVO8Hh8WNmOsvYSRhKQPlobc
HXjISZcsnYMCe4mb+yBVGz+IEHqxtngpjPu1CZNbspIGTI9AKaL6zR9HHEdBKJTWryfbCbNOaO//
5ks7aqZfx4zERqFX6vOBcKNWa+jVhn+w/gRuXf66/lPM1HdvKKr7pOt3NIz1e5MIxmzH/i+bvjTX
AXKS6dvvp8L/E9V5iXpHkQzIQ199OTfzKSLHRiB9j8tUMG4FzrmtivOzCrlrkK6f2uneL0DnPVvb
TbhYfIBGRtQnPGLhZmyk+M7GaBQqqB5vLXzBbDE/NNA0RKVeL/rbNL+Ibl01Srjg88SQr4uHJgwp
vKh7/hvbx+Wlp9XU+9GYHJmRrq/vo8RzY/vW//bCHiBMZuBASE57l90E0xa1hD/dqLmTQZrxkx5K
oge2dD3G6EINzWkle4k3QQX+LwArlawJiwlToXcEHRLLL6+iQ/JGmDxt8QxxHVLhFbHDwGfs5OU1
JBTcxexEMGTNLHewh4JOgGYfBee+drLjNUuLuguuzn7NbNPLkpwGt9L/naO0mPYGvMR9c8BPQqZj
OH8csXCCC4e5awu3L31cr3Sae1se+jjitWdq8SphVBCFGEp29wtJAsbHVe+Ku703SZpZu2wmQxv1
FJFoCNHeFNIl7tS3ozXiU6LEHx7YjBbhU6ZQlS7OqnSuPI806hCnmWaFhlz6SCgArmhB3OyoC9a4
7vOVWdUJ9cq5WJn7ZkHA9bVJnwf+G1ejUECVjo4MW871uSGWChQei9zKav6qajb6m2bQjDMbDIru
vja9XAhZL1m7gjKsPoNDD+9TzcS2g5sgs/frJFa3R5JxrWAEU7qCX1fzxREtdGFEqkdo5oLSsVNg
4aRRxsZUF4MM6iF/Y7pF49JKTlVUo9QnPlXLNxbXW2ODdv8vjduCo9yFmY39i7GpVea0Tnnqv5cn
vchPNNsugkRMvfx1H+5TFKj8z8uXpqlbXEPIhzW0HH1j8L1lyKX5lprPVLLrWfXucwqD+R2XuTCW
eHxYT3pktqSPEscRTglA330eq9QruDs6UouUhUJwewdHZbWuD9DzY1kx8iBkhxXvKmv0jt7Frdbc
dkFvbTyAj1b5OTT4DTDS6JUXLIinjdYiwS2bAc24GORXSGaCiRnNbPZgDD4CdNqPfCHDfDG/lQO5
CZv9/LyPWJUbMfehuf0dJ/YFCqtA4KobMSx9+0Yb+ZnDv4dZG4jRPlys95PRUcjoa27uTzd6nFD+
N4VCndkqj6r7d4WKhiRM5HvZvBzBSU26DWXL4NeUkysK54j0ZI81e+D6uJhe9HxPwcLdrFxJj+FL
RDwH/mkt/EIWvVssWNJpz3JOjKEM1n5xCE9+S0/pmqxfuG0T1JgqxXLJTcFo7sCtXM02m9Hz4JJs
G2HbDSYw5Zhg9wAosIczzlBvGKRkMA5TKrVw2bnLCMGqMOhBEWv0KwwI8Js+DLIBd1xPmMYdCpEe
7v4khOAWDHATOq3CVLGDHt8i3jnSkUw6KCfu7BBvYjCeO3EYxp2ZL7jai5+inA4kuKw8Ozxnqw67
pG4KcAUSCuUX1rkl0OlNmgoGFEr8lwi4CPLbKLUko4+0mHrtfc/pkFrYlyS7BX2fkyzAOPEO/Ohq
HoKfkhnw/uxC4u7CT+L7mQ9V/oCBIeALtKyw1zqRep1AsDORXBL2j16uH3vm9jecgZcKF+ILLs05
gVeMleTrfVijNLwzvM7iWgXiev+L7u+8damvNZ8/Clc9/qJ6ANC00nlyW5zvQA0IPxIz6n9C+SL3
HYVylsrvdTqGZyVm1jbi3cln4BQIJLyRwEGNy6j5NRND9/YoXlrM3jnR+5lA1Z53fh34WRUBmBvZ
PCRZvKSCK7Ulm0nTEzRZn5wT36E+ZmyD4jVzCrHRxjzC4riTfKDihT28bwidOZIok7wQE3MrnOhb
KaZnyIhmr4JkKO1did6ZDoQxwRqB6XVWHmy+nhet4Sm0NMyhSQAn4alg88mC3W5WsugBBW+xeSIs
L39So/iXpRfebgsZ6jxBJDmbosPVKcmjgaaGpmnQ0CboRZarADrFurWaRqdY8664ztcJATQSc6hn
aqSPu9TkTdsVEywH8PyKI/15wesVW1cF7kk29Hv3/5eXzycez+3GwGt7XJpRiM8aJDDMhEwoKPLS
y3k6RShdCnwd6PlUHyIUbKqV/pBlcFg/9zOh1AvaUR2G9QAbzuFEhIAWoPNElroxdofeCblyfwXG
OsHpI4An7NwAnUsAwdxt8MmGeESFFnfapVz7f89hSVkik2zrd/qEYll748uw9pkfI6rQzXy8SCgJ
8gjcZ85J5VxXv02jYu43UXkTgtZ2u8OIR5ewSSocAhqP/9b+6CmwSbUoF3hnzvii5NWf3BXoSzIR
1JSNGY/hm3W2zoc7NMWsYlwyuXtxMJhg22x36N1cQlchy+9AMpZiWjlW/gQgxBkjAFng2ydA3oHO
C0Upa7EiwX6DnzXlfgGlyjBVeqMnkvU8Ahv2Q+fFqGuu58OtlgLYN/7BLDw1JOXDVBSZAXFCW+A+
c+WHCg4s6TobqGYQyfmbT1+A3aW7EZ9N0Em05yqzXm1VFWmqyx/OnopezEbHizLS9yieaf30hPW9
AWGlwvEu3DV27eu9EGqn0chOujDoeKuly16ABUcOwRZGDQHSOqkHpnhgkJrSnxU09oOoS4MffruX
JfqZDfGdcl5UBoLIZqfOuVo0+LAGSQJH3QdtQZGcmvczg0q7KIDFPV3CgCjwkI/1Ja+cYEyIyL3B
PE/JT+dnwf5BBlKjB22HwHnn3+iia/A3DoiORiwR14wRj1gT6qzImGIYI7++/1IY8L/sI4Gd8zYP
ehdCULU3zXuL9Xu7+xo1Dl8Z1dSopld6tOCsN7s1FyIod6rT00sdsx6DGj1LLp89qZ1bB6t5YEq7
Z+ifOxKxavebRCHjxhMd/78hN94zsFj1RQ4pnvLBsV0QDYxMnGFpZ/ig12JSLKxtTDYpe89uul5w
oOi9MHNR/zm49cnctz20GN4gz9Eb2gFLrZpwdX/TkTu2MN3GsDIe/tucEjC2PWW0jy3IXu0v9yzg
IPuJgNHtmhZApiBHNon2atxPB4bvnc0VoBXBQUdOAFhnXeBfq7uBetGftvE/a23jlUJEOYhDi1RB
WfAut6xsNY3OsTKbW3mj60+BC+2oQzjBc4g4ktESlnA1dT2wwjZd0Hq+NX2GgpqJIsY5eHl0ZA/n
HX9d42AgvtgNdC2U6djfSUlRv6vbJnX443HHSVozaoZL3MciRtjkWaowLDGaVD/Ri7WsMO263bXg
zmoQJgy7pB5mIgo4KQenDmlFFHGZEme6Np7EFZtiLVv8cPzGd3/JD/8w0MMwlpDPH/qVoisqZqi4
qZ+4CB8ezacVG6QOI3b5M/15oUjro4ZMDioNMNnr1kGsIBp4ZPF583Ky7y3QbNrc/ne5P9ixyzlU
qbSgcLAtN1XPASzgLgEWCLE4kDUkMhofzeb5pAcxXSJiXV5SNcLEDJoy8Af+VbbmrRkZa41D52lF
+cX/c4tEQ+gOpP4LDSsc6OM8QnqAVUVB95kTAB3S0Hu7Mo+Lahy1bmGBxdmNnl3/vTskkZBapRbx
hoddcL8QmtYHvEvYWMEJPzb8rAIY+RQYxO4wUhckdYDjKQJr0+h5g+4RmFLadnlgOMMIyxyucu44
e9WcbeDRldPVNwpKbSySnS2I48a4uzGM6CcH4aU+xDTNOAt8QW6fUrMUQC1EjoSFZ4ocsGr/ddOs
V3K+c3k3Fv+8oLrm10OoHC6CSpHRnrQ0J/rZD9aNYTxMK1zAsCEchtxboGnOvXIqUhYOfvennjL6
Jnu/3I+a/GT/MkvEGrHgR/Qa5vMhubPWP4cLJuBCqC8pxTzLTWfOMitFARZI4lJ4X+11wVQIz5yt
6RMBhY+Af8QjOOnm/sZbsN0C/T4ug3Gy50A4lJiDj7tLTMJ3/PWceQU3DXHIQrKxZX4Oc22dMg05
9sVEynEukyipK219c/fBHg17P8wOvgRLOlr4pArEq1T/Rc3BVpFI6gCaMCLcAinAz3h/aLil5pM6
b4x9jFw+gembdDug/J4ulWthJhcgbo8+DyOaY0WELSsoP5N/Xnaig7u/NIaCq4EqPvkGkNp1Thgr
RtgnYwtfL53W3zFHqht95Drxmf3UG9Qo6ythJv3El6u84cfrLoApge2vtYT2m150YykGrIX3mFcG
245AOZ4uF7WHj/Q2cM/OyE+tBFCzcpbi2jeGGTQLy+Vo8LriAQjEKkt+bwMMaO3IsxPMovGNXz7A
Al66B8OcWEXlVaTZHrxzU41zYJrc3HGqV2TaDYz18MzsUEMHqPK0RQDof/c+tyt7x6iz7tVN5lEx
cgXqxHRPjZcWXnJAWtwvqhkyKDN2gWbblSgh+/0PnR2x4qcmSU8rE47Qk/ls1FDMwAvktILoio0j
p5ucw+1UNJ4UvKhiAEd6YTFauO/zf6iLBOUV1yxhgHJoPJ9/RKw1nQXcFQu2mCQhkBn7gd5qHVye
qCZt2rOhNnKCGsYlB7Uzjd7HFZy4UxMvPDp8qYgQtMHXEy1kYe0dK7u6Dt5+IHYvi6praABDXPUj
6sHeQLJ3t+dVOvsUoY8CAAU/ODIk25stKcv3ry7FIuudYMX0XEd+jT03J+wzmcPJCvg2a5bVkzzg
EOmixoJuuUGVEU1D7869yZ5DTa50xdolQj/BOyYKLVuAEVosBzcJBJj/2o61SysJamuVt6iDN19C
THrEAJEoRGriQMRFzT9g7ydgAfKnFKIStn8DMMxw9x4p4A7TpeQ2jffT73x/c/75ATZXIUXssSWw
im0TXvo3lM6PkO+9qvcBZUZ8L4EPyxHHlnhrT0U7D/y4Ok/BVXGRIzMOGx0vkFUGs2Du8n7eBqcX
uHte/1vVYON25Qpio4kEycE+CJLH8bTUwqnsHAhNVW+9DkyrbKOVrbFInoPg2VTirCeAu8uAijN/
OWQYGBR179O9gFAEj9ovfMbrJ031+Ps0cMBKtTL3T0dgT5K7Itj8+CuWM4jDSuypZuKJQnPH4oGa
f9ZZT9FfzRot1NvCo0By9FLLYfP2jcCjsxgkH40gDIRJhpq/hqCU8Meun+ICLlcmTO/Cku7DunBC
rtnpUg7qR0KeE2qj++cmcHRwBByycXvH+tf3toXfo34CUxF3FZpZm6QQC7JLp9b0JBRGRBOo7Gak
fxzMGVYjTumxP0toYIKTFz/goWIgNDnHeTC/xN74zcJ32CXbaFPBuNpw8BKkd+vIU6hYNDV6KpW5
MIbDRolRyxMkrDN0otddqJrOAOzoe9yn5e/1sMBBrjoeLTCXsTZAhAf1EiDaXNwwvoWXrC0dmncT
M946/UByP+P1Wec9S2S3EI1UVsRrSAup9PpSijpjoOM/9RuZOtcXnPq+zrL4ucgGk91XH85Jt9T0
TrOjnMs4DLtUEegs4NOWIK7swoKrThIPs0lDtzOnWg6nR8XKxWTwIGyszkxY++eFj/lrycXFyZ80
W0nNBG1x8Ap7Aq4L95xkSxkmDwzn0JW498bq4BoeUUTAjNvobJ0MwZlXcoZWDFLNp31yOLJUgevz
y54MEXwk/0d2G7qLXE0Ku/GPSoLJwCBc9CCFcqBk637eHRgBTF3E/wzocKjf/qXsxBG3Otq3Y2wV
fjhHhhEMGmkyCQAjDxdBawH9WuQUTw0aNH9L5N/jVbIe7hbIGhEORAIgkJxQ+jP4igS2n6veyrgA
WU0uyEKlPNC9ga0CtwdTdMmc08xiIWYwO/aQqzKFhgGMsNVkmWTQj26nKO4hAc0/+13UMZbT12FN
RwV8Toacwhmgu+mGT2zMlxKvFi15cle0CuxHBtghjIIOi02iH+lzi0wrIB3gPZ0CnWoBwln+EU3W
usPCe7MYWmr7Pc6NMK3naOwzBcQ6Lq5uKRsnsTphh9x0zl6PbhM57N5DvevOzQc7QNY0AOXGk6Ic
drLTTDXUrkTZog6KHH3Qu+1p1zekH8pAheDFymsaEzQB0k2j/XG5rH9KyIO/8ePk2JENztfN6YMM
nobd/6FPNo/VNOdKNFgNFCTn+0brYkTNX1+S8m5k1F1r6O2SqfJx1KzRUQCOn5ofgo+dbBkZffmg
EjbszhGNpg8UTZ81JOFwKP/3GjfMB6fiLrdbYCkEqM+uNOPEqf30sZj58C8QOx4KwR/2V6liWzsh
UYOWH/o51JxOZl+l1jqOTQxqTlDR7c0w3tp36pRzy4MvCtTi89tyL6Lrxwawuue1glPTbD+zSaVw
Q9RDLgbCbcurnITdhnUfRt3V4Ky+GsNk6CY2KvgVpEtBePibk90iP9J3RGb62grKHfV3Zs4cUgpl
pdp64xnP54rifWVlYJByFYEInGCH0Fj4g4mRbS92JrBYaqmEIvdFps6T8lZZP2O0rXgNCLxGroIC
6R07vi6CZummnldue37G3EeYp46bTNiY2JZdHazsR0Go3Ma6ohfqetPaRAKFJBmzRw2RmyhvJmbg
d8i0qHciAaQz9k+XzIxWZ/q/rLGHlYbv1OBIqE6YFmmj81035oFAcFaBI3FoC64oY6Eu9E4/GvY1
fwWKpJR1Z6WZLMSZTgl/aV2/NXSfuw3DXQFrBtdAIDDQZqf0xogGv5Mzzzvh6L5iLfsM4PB4065Y
6Mrid/Rinwrq0OIoUvxPYfPnK5mDo2Xr8bD5Gu/+WJg5U4+XWFNVLidjOrX4AzQ149QEt0ZUcgTP
GbQ/lPvf/LxrpEDKeR/y80l2kiFoDDM5+hV0jAWIYT9OC7JSNw+gNNcirSP6piuf1TNUQCaVn1qx
utlCWV13SND3nVFg5U29qjQRLG3ENxM8+WZmpPDrie5427U3V8hjxfnxZycuncgiF5y9QgPM3tkM
w8M5KBj5sDpNLXwiV+NM+QNZgjcrfECGC33anMhe0oHphr9r475DBiLbAUwMQoHD3co+9BRw0J/x
GAM0r5yV9PHlF4sFm9hcMp/zB927olqHF4ujVg1qO6FI0HnK3J2bXRvofNzTYOLRHg87wLpogvsf
ON+d8bviBZbSzpYhx05Q+GmzykdL1ljAToDak33Y3IoqoxnByIsX1zTGvuPplea4LqcpwQffj5rp
jpw4IcvB41PLBCkFONzRBqLEutXOAj7p09mijSOsfCWrXOgLgq/0PR6KjLaWmJlIZE3za5+zG93z
SPRbiQCD4iZAK9DWXGpUY2vONgyY2vUUC2DvU0KicCq2LGY7rsMs9qM4vTv8iGP8MVs4GDe2BA4w
EZDAJpR1H55EqBh6qPbEQcrLoD1CJ7YaSVYo9l2vckw9ztx+khUdPJilCuig3GNYxZadWom5VdY2
IaLicJuVXEARGrLzID0zyMcYraBJHmHYKXPXSLsFwJZ/nN5juP+onNBIodhnU17EExpHrdT3YUak
T60vSlErDUSZRs19VeO8M4UXA69efLB6Mz/VI+M/UCxTY7cx9376bNYAWHlcuXNqjBwmA9V1uNQ2
8q8QCVaNQ20bGHaFQ5b/DyYyAfGi/Ez76PVGtjjrCrl7HwYwk8Tc8a9S88Eq1TRQDFuAOcjCpJcy
rnyThqVD2B7BDZCYhGdwKsFbFatNPKpS/NBEJgtHz2+WtEenFCquui2ba/b4rbK84YRidwxxAKVb
/mfei0z5ipZhGS+P5lcBuq5MKflkcobd9oKCYNRmieQdQx0A1m3i5aF1spW8KyHvHv5AcYMmtu1R
MEgM//hqNxGxF+amHpQgfamobDQxkCYmyaceoWzYXi9K+xOHDKBKenzPWoNhnTdsoiOyzG1uX31y
+VoWPZZ/onVbjVsQ87hico5kB6tge9zRKWroG5VNdglGYVRZjxU3ypwG1G8Dm+3wHIddqYjjSJIC
Lm6eAikwhgdhfvmT5QqWAkoinC4J+i+tZRjaI7nw2zQ/vaOqj5tXrH4dIJVlNNB/04HhVOOtM/PV
AwPPhOP9uQR6w3ynmD1h+fYxx1zyf4hJyy1cZv+rtr5IX5M+20IbvcEpdgur6pMJgIWP/dC6+WJ0
o6IGFsI1YU02beT1MoRCvodFbKBDYrHBuW9G27b+xRyOxnZv1AiUN+DCcy0xVOM713jPaF4fpkKg
gNaimRgYDfl810ekqFgGUGERBCUiRx1U2UbLJG08GHQGUUi2xWk6ZwmIwyGmpxTl6P/e8FQuchjI
vgRC1L8ouwN/sFK96VWcwPlfSqnhKOsTl9Y7uaQ2l+7aqQITe17Mn3OmfOt9G8kv4vYi5KQJqYeV
n8BxpDrGq+6a9exTyw82BzaLsiwiuldSUg2X1aOViyDstaEcF2+/lHT54db9KFeTvjod5ZSXm1ts
yZtzP238VrwQiypeWM/NjGDjV1DbSzedx9DYkuBk19peyzuS4x9OXqdep8VmVCeGk1FA/HjKSKcK
OguKwzxtdV+GoOAWc0NdkmjOTwWbqlOZkplYvglSqram5x9yfzHf7cBKSql1ybxClr1sgRTbXKvp
K5TXz3Nsq1JUy1ruX4n1zHeChHWfY04elIwLkxXDpzeGHO3+0kQrzeqAxVsqbRAbkgG1eJb9sdNo
kI6UACxbAa7Vfo3J2i42dmMRhnWzcHL42J4+o7vjlVRPXSJ/MUUpaqwJMTQrqlzS34Z7FTWfWEkC
s0h52xO18Q58cZ8b0HfytTvG1gG1YYfmraHwc9X1yfMoZUlHE2fsHkFJkdVbWO9eoSBvY5c2iyba
k2kThVu9Ox5zFhnjYKn3EPNs4rttnbp2Sr/9KNhu3Z5msaHqWH79Xvd+5ISMFcWef9r6fDKiZRth
SAgKkzxK/x4SbgUM3CcTDxnxXC3ZUU/8rinI99D/6hqkJHAxO+m4/F7dYtmebFt2UolUqtlVqjdo
nuhGV8UlI/EsGkaKmHV4QAEFR8sFqfMkx8NzfKdE4NE5EoXonr92xueX3ohvn1n6ANmMqEd70v3b
05Xtnh3t4jxRLjPnnTc8Lr9XR3KTvgaawqSjmBbjUTn5KDNf7hkS+E3EocuIQiwcQz/ZqU6ey4T2
Vyhpv0fHMbFl2tT0n4KlJuqyL/ejajYbHSb6Jj78dqePAnBYo4z2h6IrSI7RxQwXZSVRSzVn6oSS
h4oCAe6dTAe97xOtD1SnjnWqNc0vsZhmPy6Ot0KNnw2y1042pfdsc4zzsRlkkVd6TOqUwBxMaOUe
MXM0UQC1xndVtReaTwX047ajBDYORm5ybi47Sey4uFM+Bq8WNQglsDK7KZ7KbE6J8rga0WmOBxIU
8wQ/O87RSj8ElONWHeIciHMsnfwljAX6NZpVwJDl2O33yfZECfViuTGX/QqccCxUHaoLRrUFsvf5
yTj0eldty7z915lphBxWK6IppUF4Q7hTOsPD0QtPQy8ah4hnKNfJye/OZtH3SG1aDtLXLfBiSTgk
erpzz8/K5WIMOfZUENSsbZaxqA5KWjJQScsCzAfYk7gS8CiB/93KisLAnXbvugsCgjsGr/7nrXpd
SEyNuywyMQrdmxcJJRqXX9UdONB0E4pi34xpGkSXb2/ufDJLKG3EkcIe0L4SJBqNIrk8Pk+f2poM
tmXRXsaUffIRB8NZffbJuqFY65oahdpc8+V10rp9vGd/B508ofjFZuncFPd+ekP9UM9srXG+eBL3
7VFHatqIgNyNeksLfXmAtXGM47DoT3QvoP+ems5c8QgQ4H2MTRirYKGWuUe4fhi6ekWSGqGU+QbE
PEtvAPCIrxGhAXbTAWf4kjGH4jZ/J9Zc2D9163kb55klyU7mUCdWg+Yi9V2Tt+Kdn38iylVRUgXg
UGDc7oo61vxkGjgv/cxSGdeRQLUUUjNnGRtUTPrC//b1namZgO+ZfYMKl1bPKS7azJL2uaCq64A8
OXZwnj49OMRioZTDuzT38q0UsIfVKlpA+KvbQusmAdRdz8JT0jRWOn5tLCMqLvm3skK7FDg98TFI
E8ac387gKXRyXC+3yJJ0TxRCHXS9iNqHblmqn1vPJY5zE7FbRMDC+jkzWwYoMsM96966tMyPeemW
Uct25ZbZtFNqh5mk57ggKYAw2dzqOR2xqaSGsK4NLUVuAjentbb7ZaxsUGZkCaS7cojKTdLnRoP1
loxsE+zAUHSAqc7ryYfPxjLKiGwQhnJvuGX+MCV0B2It5Gb5Qxzr0fAAo1Q9jWfNC1EHp0KE0mBz
XLGPAuoIoCgqXmQqwaHWTP/aG+SMNtdBTaDpOp/3R/qoj3IBKBuP8yWZAbuT3IflNDj+gVieuObE
eEfodf7pimw7HqTPiSgEWwTS/KINFZHX++e75U2ylnyXbqi8zWy/8Sw/mjbaErJ1u7ymQ81Ybsdy
UGvRDsm4Jjp6W1tIU1AeCS9zJfgAn2ROfaUI5H+xIJoqTgOu6Kjm4f35K3NG8RMh4YhL+C50mZvH
MvNP3VvFAbq0due38w1RPtUWEoCvyqDS+YKt1QBETRJtVbTa/5JdlEf5XdH5sgbmSfPpMp7NRu4A
JS3NQ5iqgzX+fr2QBdEStZywyYQxp9dJJWTZx2uL1gMfuafk6m+gO7gSdH7hmAM5oGoOvGaE8gIT
ruQOhrEl46s8m9GcUA4R+D5y6onoqVar3/TXxHv3E8ZZFAf0joToJajvaRBfKs1gPo5Cvv9rERwd
epAkEZ+SeWoQAfJCASjD/l9YRFm0Ak2dKFCEGuUL/nsgHrG5vc+0iyilU08g7eRZxAcxrka5AFJO
4yu/RuTo2se69jx/nC8+G1IqfOV//xX91S9qqvJuJhHvmf345ljh4yQ0Vl86JhnQaOHZDRSx0i8m
R3HoFU3vw5MPB6dGjQQL3I7p0MJKbdsupLVwhgshC0Aysal6a6zAInFvcJtbJNriSXKDGEG/dGRN
9C/ZR3RIN35/ut7coDw60XluVW38tu2D+ixb/tasdFgd+Bh47IT5i17PdPdLMkp/68BXbqqjrwJ7
HHt2oYAUWgviavl7iTV7B0s/gzQoW8L7FyN1Zmzq75ZcD6+dfp151bEnCTj3r1/ra0+4ujvnllri
bDARqI4RqlB/Xw12VMvbITCCVuyMSF/KdvdNxGhT9LaCm8BY+cW/jv6suUmsycGY3dEflP4ZIkAX
oNHQJXK+8vKHMCP3pH/8VKitUf3+cN5ql6R7PnmmU70/94BMEaDyjomjD3Q1aydjTq7ncpw8MWa+
QCw0zWcAau95tzBhJISKEy2EmgC+8iyECJKTeVWuI81GOSfC24SSWWB88qSxizCkdei7b4LjDkS5
nJW6VbGMhZJ3HsQCI92Iny+o02jPctX9TeCQYPhu10yE/XoGIqjK05VTj2vQQ62/Jxzd7D/HT/YC
ye2izRcg4R3uMbe064yAgPS8VTb74FeA2DN1RYJ5WSYt4Pq9fpXyy35mLCdTWEZMNoxipyFqhtr8
6L7Oek4O1PLHLut3iBFRulZ1LgLamuelkjeEbn7WORskklAxun8YjNdXzrbAFRKPBZo9bZcVC67N
lCqu9l8RXlIUfg/aAkBAr8/js6Y9jkLLha5YB5yvN6RJD58eaMhCOrj1N8HOewniXdR4jbDsbmXW
ITSd5muaXywUIgEZZcuvq7QxG6CyymLfPn/nbL4lmYT4U8g+L2O8NVktT635xTSIgvQ4mVu4ePn5
k6aV5KnqPadosq+f67ohNb5VW+DscjUC4rv8A4LjLw5/2J0bCGDFoAE1+LgWDAFtfpCQ7iUWWeQl
3ViayxyGaVWjI1qaPyOYlJAd0v+7darIQyR0skjpyFLbEbv6qE5zOt25QQyAgOi8CKi/4avHc0os
nkv+5imiV3yym1+pjkzxt6uzn4hoHjCes8H+hqqHvHnzy9zTFCtNeb0+D7d5rIDDVIGl/4GGOJFc
MXijcRw0hnxKVeC5WIaOHFlscgOzu6Hry7v4jzSGQ4/xamIMc77+utfK/K7jioe0aQsjoAMI3mK4
rlLPx/67nlTgO0futViHz+AvLzI/v2PU+tQOsf6JU4cx6zAAzmTm9SMjyssjVB8RC6f3cm2Gfx4V
UNQZ1PjG+Q4C8DRHrHmk/Ds4go3TiMpxqQPjsEX/fdrFFD7+WWkAjTGRztPbz/mDEmFjzXSXlkVV
5To3vXLuffQ9hYjTm/mVjsXRzirSlE437Vmhcm723gEHdn9+Vs/eoxBlH5cbVtShz02JrWPRSzkv
jyuQn8V6ynGmGiCxx7o1bP7Drc7/mH+CaoO2Rf6wFl8GxVpQHqYhgmTI9czVInVk8LfA6VvkUK9D
/Z4tLs4m/9SEx1nvz1d0CrpqX+Kp2f3rSf3JiJGZPUt4i6cpFrMtwMDt/zUkkhhSIAXFSks+jVu4
CwREGlRQbUHIlsI0a0xRTFU4gnpONLew5Z3Jm5eszEsxD3gF1V4+lz2IWv14oHiJYNhdGNhf0lLp
l0GYXCjMYT9T3D2rPHB4zIv/VmmeFHAL18kgME302rz3mwzf4G/DRyajlGajZKHel7ryWVYosEvs
fsU7qbsiHXZrY7MVlf7qQatPVdvbc2s4vlI9p4e7BjyB+cQrxvLqLDjbTjcK7PLKXptFL7HkAUWp
tBdhiqauNFd3BpFoBiDQyvSxX2HwtCZhku9axbwDn72/zDWVtiIGjIu8c3E7rD93aTGYI5N7N4XN
c/qQAyOd47Svhb97FJjdcShJTK6lLtbttcE6qaifVfbbD5MziIk3ZyttXhPaO7Ma1czvVdYlNy/S
QxNDo/CI2ocbcqFSntn5WLbz5ddXEwPPNv+avN8Kzram0CF9KDQUcqjR4arop7VT0fqDgjyCXlm/
ATfKujkvqvL6dGt0SNoHFVdFanWKEcCBDarwGHcBZL3qtDOb0b2YxqLV2dk9M9bzV/15MuFepM9a
nx20JKjZL5ICSQmAm+T1zi0j85sxkke3LAGdp+Z1CRnmClV/tMwMXAJVk05B1mXVca/dLP+Uo9z3
/Mt77yqKTF87+9dI8syFtAtP1wZk4yb1wJ3CoFvbkxVpAbC3YD/t2rK6lvRPetMMpLAXqXqzREkz
qIpx1xXDzD+t1HLJWD8tUzlSXi9gbWZyYU63sxstUnu1fvbrefNLRGT1kazUiCmZbtqHzux8pY35
Kx3VWxX+OemLm5pYUUh7e8KfMCM07+Qgvb+XU6F2a3uQ/0NREnnEdd90QCpxtxQLk81WRilSeiDW
aFSh0ifnUAlnKmIyuduLmlBZc6zMWoj2nsahwUbjAPgAL0bFL8zjNQuQmmVUFLNGdKWr3M5xhcHN
EC8EnxSAOFQTIsKckfmN6ke2qFI4f+CWoSD1RqfZ4D546jmidAp42vs6PPCFl2L2QIMUY7e8x7b0
3zKL3/TjTPc9V5kueNQejHfCLTLTvJjC1hGaPqyuCVZA3HgxsLPKYZzPMa7IIhC/0n8fOE9Nih6p
UL4PE16Gop4Z/V3pnGeZrkR90e1r8ScthF8l01cB5KSH7PBDmaTjivcY2OoJQxu4jmH6ugfjk1mH
VaDIPguWlf7qensCld+uZdZRaDT71XNpZ3FwTs9/cFr3VakVLnjqSnXDTkmYea60lVppitNJTuM3
hCGcqzjrzhA+vUIxrE3fEJ9ecATvSuZlU+UNSTaeoo4MAVzGxJtC0CzTUErfqKN7j0sdTXywHi2H
Trt/iBGjNHd5cIuPf0Vs/fRVV1VxV4g9ddVzBRf06NqHMXerdj8XMy31cRdGVB5KIjIxuFiI5yl8
j7K07n6+e13BBLWUXzhr16jmu6/5vu31fddMxoMr2MTpcte6fdZX60PjMCW/Ll5K04tGOVKkuCyg
V/tKUY+dIt2Kf/MyKGwGpAv9jFfjynVZDxj3Lmbs7XgFYtArX4MhgAB1t4TKIrr1jL9Y99Y6+6lh
7ey6fc9InJXBdtdeyu8eyXQzLcPMFXRNSBf2QGUJuK3HuEIZetK9NF5FCl+1N9cJ8TvsOHC8bmMa
t/+ST+OUuwmMcOecxcFdXOqdgEQIIZ5wO71UlK5Qz7aOsjbhZvzT7CV8CuIQDE3rLLk1zaP1Emyv
R+NQxYhf3f2jb9UxC4+1+3ULpj3alOZSDN0uGiQ5tD7mMY4myN8ix/HOJtkB0kuh3oFhJDnLGur+
tzw5duCUaF8SBxbjLhChYUyq1Igql7cozexcAh6WlsegRmX7iEpOMScGRXex6KcX3Tgs8tcpn2Q/
rylZ/55puJOClwcP24AYwUvu8S1Z3bWEzSy0OAPmBosxO0ormueYDiuTuhWmC/pQAM5G21aEjisI
TD83cyK0T+oVM6AeCCZFSrJG2CN1etI8jtTg2Y1w3+R55AkGeow+28FDmxIO2P544hPwNRzimuOC
CLCwwTkahroPKApdzMyOa+3AnPBpPW1rF+M7fera5E4tut3X2ererCigPn4tJNYe6rcM214Hi/KP
UDR8gfAW3FmvFHaD4wa6ej5iFfEf8lvdDtCZfRN+gN4tg97h7bAvK+j6XWY9auT/5aOivYWtjv8S
bv7F/w1lkQmSssMfaRbDudEitNYZhyCNecyfyw85D5cgOGFEc4Iu+9goEN1NJRQ6vN/q60KiWRc8
IEkolhZ8bSE5YbZY0fwa4m6ibveABv5G2OJxEZPYykiy4rBYWjmKTh+GQQfoWbewAffDmkhBWJTC
juYwIdCyTPmmJj2+wGS3pJmLhYbd26lULR8wlFlSsrgT4YU8hxkiE/g8PRGPwKE3U+Lay5TTxHDC
joGObXmmolphSlJ/ZRFf5z8SdLb0N4NXxzlO85RsG6uPDyI2GNKC7uoSNSdKM4JU1pL/ZExgb0og
FQ2KPWh9ZFYRjx8ZNp0c2VtbGwQsxhx1chnari5XvEeX6ZMNIj+bJ4Iyc0xotWoIS6ni/kFeLsV1
lD4/jYXyqOCtxgPN97HnqniFz0TUyDEvP0GSA1tPrGVVYIocFAJjlBRMb1lwX5KVT601di2xlyhA
RYInhWqGuSTvguG9vGQlO3h55WXjaflUhFEqzkR40p6A9dLL4Th+2cRZThkpjiJJAbKWX8T/8muO
Fn7L8IRnG1f4lqoXuZe2TskdUef8Qb0ujxY3gwkg2/HhucSrab90DBacfy5aXRDtPNn89rbwc8on
45hzzABP8VnnFDO5+PZNwslj7zd4f62PBj6bjkBxhJ0hWB3Xj9xOvuN3qWpmku+BHKk1kdH5ZXVS
o99I4e1DjkGpCjXIDbthoWe4ATaAz7ZIX3zngTKup3fJ+SaTq4PrmzfKsqBdhkyVLeJDNIWfcEZw
VcXap7JLf/vARAA3ePBxEgHiiyJQzpwxKw8UmhMtUtlaLLm9qfFW/Kg1KtHRqxq0vIY0F/OgIiI0
q0Q9yfvNKAitvTwPhsAP/CYGk5C6xdIwg550NEsQBR4ru/Appv3C/7ATuTUZ8Pj2qzU0caXmf5Xr
CfwLvkRFcMglEZBv8QcmI+Hys3UbkuY8esnFBtkM7ir9pQeAmvbb13wJx3dhoN56/l7m8Wo8xjK8
4gFcNV7GSW6CgcCng4h//xzcBFDxDJMJZ6fwIJKMQ/BN2wKmPLs9Vz93/JnWl2xscPgkf0JPbjks
aXAU/FZX/qksQOetn1kYjkXGJ3GSLU8cHRaQle6SoL4pbYxCNgsUwU7u+44aJIu17B67qN0QHruQ
iAS/D6SkXrAdMNBl4I5iOTZEl2AWE9ufkgcYa6d4MlfiAgUF8IvYFqFs5GfY/XhpWYURpdMMFiVk
2HgNMxGDk0xwSA2fgFO45vQitCpkuJC+TBH7GIMscc+cbMck+HmzP03OZUFJ2vHokbSuwvyduNpO
c7OR7htRrAv2nZ5tAfcll2HQCmCMgYR1OYteu9OEP9ytvF7JFIVr9uOlPU1WwcFlgt9ODySisHY4
MkFsjxcQ9BjGoqgRuR/DwmSNSm0liTj+Ccl8mLJbBS3niAAWcBcvVn7qIoZ9PXhzJ5CPLRh1dwlI
KMF174pIRael5mj4XiSMcGa7n8+tMU5arukEY4o/ZaqnoervYJAFQtR/+jwMB5v9BelIR10r7nwc
kCbg4fAZYeU9PtjcFcoD2l2TKw09fyBakqu8p6/U/Z3LMhisUn6WTKbfSToeYdRxeTm/v/tTiDpr
KrUlscL2FX8N7QKXlgbgwNf+kfo7w85jXD2kHz0GyC+NtjHnleoJLsc5kL3g+A5mSTmuBfM+Dcz6
c3dP+tUe9BH20IgxUdPKtvrBzk3XsIET41hTbwVc2xu0lKpPZ5cHPDCHr6eZ9u8OV9f0MBOSyFg2
NDNG4M3fnZ7cJYhxXbjsVliCq/UnTS0fBpP72c0nGkIDcWnC/JvyERU0zjePWrClaAqIJy2azX56
4jrM4Thjmr30kFK0Vd4DQQD1OUSUl4yknwrUfYSK6yPnoes0LcrK72Na9CBh+nS1lf92Qatj3Hk6
pSfl8b4zMxSPaQU29Fc/3ca5JDM93OmkqUhrJb02KfUFNkN/TKeC2Lk/kQoFVj9KKnC7Jz5fBXTM
s//xDFNLqOCikjsSsZ3ds05LVvjqtanELcclyGeXZh5wtYwxxnYhwfNpY3oq/BIjU+4Oy9x4XxsO
SdULfWlzbeXfXLufIKgJNLTqnn8ia/wKuob7jJsBX25dweQBZHMMqbNggTDji/YHTbzOlp9FbGfw
iSt/4cqUH3wKkxvxwwxgqlE8wtjZCCBb1Gh9MkNLWt4KIqjOuY2ZPnTjvI4XqwEspE98QyrzFXmM
3d6xXxvJORjiIsIQzB8iIdbn+Z8CP+SUf8uPOfiq5HaCI4uu17gkZlvYWAs3X1dHLWKNWAb/0BhF
ptOdwqcdVuW5BqEFVcV9+F60vbHPncETMfIzs5zEFPgcLvH7ERDA3JD1R6yR2W+Dhh1uxIp/Y4CB
agXC5Q5TrC3a4kqFmILYooGLENCwwj4mKcnLNemLAnubpzooEeIZQCmMTNI/7Ar1M5mxTkosUWSP
4EzFLrO4rDHV8gqXUomQ8fBzuiiyxPI3GGLKJ+w/o0utLRADNeQ8HYcKMh+KYR8IXiMT8Fg8AMM9
DG8ohNkE/jGtRmkCgWy6U7oKGTZEdBVCME3dTDIXx/niLdEuuBnjQDNr3IubNH/e3j1XvfSgtKpv
EZPNQOotgZkRbl/Hb/SpCKxqwICKHiGcYfqCqPatGFRlNRIgnxH0bVV4/c9pMVwZwtApb2saOCbI
rGkArQvOtXmFsA8DAiUPQ1IUNXj6zyCvbKXoPpLxxB6h3plQ0Vl6xyk051KnKIGpDKqQQWWNG4H1
EZh40RQKUXzFDpBl97OvoJdP/vAIshuO+tBGN9WNvmoPMzVArpuZO39Og1CirrbX26YKJaayLjv0
RbnRKDRcl0zJu2s/D3SVc8MAgkfnAu7EupssmvDtORiB6NRdWOIp3UtziGPINvpBINb/iWFQ+vrO
1hxMpoLd8zBdClV7s6pydtCWV+AHrjS7HbufNNMfeY7NYpY4S6ptBKNMP0EWrckvbnjRqGuUwKHO
Y831I0cjPeiyu0f3Pq6u6XrSkNPhCHGBO7DJQXLw0rXf6myTqYQU2qgazWIM6Is4juff2FLzip4W
vHug6EcXEIzXoXz3jQmdZNbxyli0TAe9kX3m97fqiIZb7jB9MMXDU411UpfT+QDpXTjQadz85S8G
AxlUszbtmsRx240TwZKrU7I3slUWTW2cSkOKfnP29ArrljWThD3Kd3Gi6yhUwhdBG7brPaGRkco+
UPITemdsQ8GmQ6gy7iPU9O9jk5ud/5HwshDJUKEcekLK7cMMMQp1BvQUqOgGOTdZ6/rORIHJmy1y
MLj5z+IW3S0ilU+UFEOk2TBC52j+eDXRwF1+LQ5wKTRT59mAz+V7TGXXGA9vjZ0d57pMOREQofJw
tXueHaG4uYw5Al2YjoEXqA4wTazjP63j6cJm1YEAE9kvIrtWu6gd/8onsoZKOI/fzeFpdtlKaPoK
Sx61JRk4FcDgv9erM0CQoVrNfqTW5gBex4VYd1S4mdQ25r4B/mDtKItDMx/HAb3+V6l9AGLUBkB8
wGRPetRYCFHehfyqoWT9nAQEDlXlhAoVUE27jRhBhlIjDmB9hjM/cAHJC6DUZIK+9ErRD5b27Kvp
3G26yhvKEuqyEyLCIKNGCoMeOR72hDQCoy/AN7a4tPTvaZ+PT9OxqId+hK16V4XxFfEoCVA7mVbU
MQSMA8iVPXgaxk08qZkaUrz65OKccW4454/KikZRcjMq9gsi11LoHoRfYusp7lV1x/LfmBhjyCyI
4ENUQQ/pdi7IOh+6jvjedjHXxWItajvTCZjPCsIO3+dakHVmpXeUvbiJs61Roc99KhtZu+1L89gf
kZVU2gWF4/jaHpko4DnwcXlqxAbSAJafQ+DWyIQ/kGnZ/YD/6m/F89IbKZ7i5saCePj1EP4lih0a
GiSoyL5TS/PNrn5L1DAjIyUCM03mVpHNtKaLtNlBnUOUzN8PgxCN5XwVNZ43cM0tZ4HIizic5TYU
jSM/mofvDZ7SH/9nF/Z/h5EzdF/ZsfssX8n+JVT6/twXPs3SkoRnquqaeiPB7nJhV/RfjLysTAGp
Okhy7qk4/cn/5i36zfvSmsd/Hy1rp29It12f9ywQ09Gaj1xlkYWjzCGBS4Pc3aPZB4iS1nBkD4PH
+Manj759jyWHXvCJOEvG3Il5yDrui9KyPw78cvT6RdQkpuVBGB6wW64AUoZ4d2XuEiBUou26Fuo8
W+5tuZjLTnLRjaldPPikCIG1uvuHuInvmdVpU0aW42zEXICv4+SFau6hJY1Bj1VCbZHUhvAqP+bZ
XaG7fxVtE/DC+3WtT+GzSdk1OA97904mRSxsrP2DyUnR8mV+e78TftFi6W8u+4d6+llgUE2iPn6W
3iu3LUV55rr7UMz29mQFBmozeSiw795ke5uE9G5rOEhqCVr44m2tlQ1DrGqb5zivcLCchlvXage7
/eVPxiUfmDr2n5Q2uJDH9T8is5H4/vA+wrl9RmW5z+zokxomIvXvK+N8TedtSoqK3qtZiqPN2/XL
O5AaPhwT9Lt7lcaCW0HrOE8fdeQC7AL0WWnHrNv8FuchBJffQsrM9oZMQ3Dq1U9kuS7yHZnvgrGP
C5AJTPcYx0WL1+7whe8MXePxpqMycNfdE0YjzEoLOyEF5NvGQxqcn7qa2Quw15pgd3ax8K6FMaX1
cFPqbS9WBVdBkiCYpDHxQVTNZpFm607ref4YGWRAgzDL6m4EnBcaFPSNGdxpTHedTb5OAAWMrGMg
UGuXhgqZY0lvhiLVjJjRbiCCi9sxXYSPGd7WcBXSxRr61QJSAAk6cLyzRQTsLjcU4hxGjAicfPKw
mzUvNNMwl6gpbuSpPsk4TH+UGqZRv5LREy4e/2RCN6i2IgUmWAKis7wu3yXq/vgXXs3QkdCnh+fs
IQ4l8rA/iL87sHPR/cxhzu8eTarkom5/gheJbJE1Bw2EGomyK3PrS1Um0oUYJH5cpytfxw36ExMC
jtQj4YOeHGOqloW0GSMn/M/1JhsYxEuO1ipHcGYaqoFx4S20LyqQzCutx39F3nc37siSyChrEdNZ
dWu97RWhipuWjGTcCYWdF1wsuxlCjJ17k52wJZJKePAUSqHqBjqjBSoc86bsB1fhdvszMltf9Cp3
lK0BMF4PfVfhWBzdICWstKl61kUpGGI430fXM4b+0UBRTeFBBqepC/YoToMTKeT73BjRgqYEX4Cg
NxsYoQb4ARykmmAh6SsV1L5vbZpmLqGPsSXauXxOBVD7Vsa6yUbUb1m+xCO7LoeymUi/nDlnP0xD
l7QPEe9d63e4N3PR0+TZuTHoET5RABcrhApYw4BU8V+67n1P+cdrrKL2A/TmSrTh/bbMp9b0DxMY
nB6x227SPj7Odqxakk/P13IynSbkz732sJuMq8jxxmd5CYLu41lBXJ9E1FRlUpL+wbrKZ5n4GQGD
eR+fi3DIfKiFVFr/Is2X/JhOgkm2Sd+f2HeSEDeJwvtzM0mCdymvupRmJMrkj4NKnlbpC9Sn5Yed
UsDztkf0xo9NpYOCfpJ0xBWjNAtFOFhZdqNi74dTBK9rlpUUvGC3VAczSwAe/1fQrfrx1VlcwGyt
L4VcngF/kifWjvLwPtjCUqfiJSdQtJ0H7R8RKyNypaZmCzGQPT0rztunSgsLtYC3HicnD//AJ8SQ
g9dd8MD7dGM1PP2jx9T53z9EFDIJeQN1XpFqMr83QnUvZGL5lPUvocjvUbbstTr917WWVbLQMDN1
CVLFTE1UsgqVUF/2LWlZQ1lqAxqLhnisTvhrVTASIz5fbbbuFqO0m4HDeAon8y5t3NQnp6+8rc1e
21lYMuURLXQynhSJG3kx6bwb4pqN3g7LxVpPzGiodA5VlkBq88vI0+Sw60K8iRMJlYje+2tt0jVD
u39hVMoigqMrUdTTPhs7OrSvIgq5lKGaOqivDT34ULE1o2pR2me87t/oQ1GEywd0op/IsJwmFUQa
HCRIZUGzaqBmDA/YSPSMlrmu7cMgwsfv7FLtbBQFxStCOP/DEYaW+s1EI9JGYhs0aXmjI/UPsw0G
twlkxO1feeHXG227uWTuyFVTHmPgj0yFasi+Qf5Lg7Za5DyBfD7UApIXTfG7dCMQLwLCjTWosZVU
hEA2sxLZCcIKraq17nxCPPpNQWmOVkqpieZ92mCaplX/aRRWZfyx0A0KMU9jOL9n2RJhOJL4/Au8
kSlkyaWTjnqrlcOqCiT4+iwJ8q3Lg0YczKBLvmFq6IZ2NMbrTZPoexR36z+ZGkeGhbBC5KPUCTXR
iwv0Iy/kIfbb8MzaPa8oBvAgJfzuHUDb4/JLsMyn9AH+mUX3ld3V4hH3b7TlmQaXI0gdlqDe2RaC
m/ReX+N+IwUWdhvVH/gWuutLcH1Cfhj3aMWCgNSVdbmS+nKamS2dvUR922OsOUIoS2FKCiUurlQ1
1IKqnAFyZQsbQkm++udIO6hW5AjnzbN8nvg/dKXX1STCMWHwBCInPwpDetQ8m4l5o+a/dYck6xDQ
ZMmrySFgwzL5oU7dD1s87dwRnRDcOw7UAhKyE9YlWOTBw8aYYLH8W68f9Bo5qh/CP8Ze+L5MGvP6
I0b56g9R+WU7kOQNRoJytrYR+WihBTx9zoMCer4o1qspy2MNIQGCkdwfW4sRbsx9tyD5VntuetHs
bHxW/Wgj5BxcM/Dhbl5kVfq1JWL9EsGfCm5QeTH9g6pwgk98yC1CJ6HTfG0rB/sf+YA/P92ZbxxA
hAKFtqoOteqpBTkTvbCBFJRimHaJFCiB/Qcp4WenehinWnq7K4VCATZ1YvkH/r9GAG/VnX1092Hj
llPE6n+Ieb2siTVXT65E4PGn3YIUqKg81qfmsaZUqIX5OXj+uNxG1ccxauX9CwyVX3FuhDLGK9rv
L7vB3p+A87KIEKaZ29OZ4l2CDMfXosFH3EAXV5WXTKc9W6DhVk2mcQ3YG7e8vW+rlGVt4E7GWdTY
sRR/J3VZ3isqij+f5wPgABeLAhwGTSzUiS8fdeYcuQl8/hcUMMxxm7k2vvQCOAmq4l86PSOvWWYd
ok+vxLlBgLBGQEOwLIXz2ccFMe01Pn302kgLMRNu5IEA3Dm/XIXmYHZgz5pG+fl2yk52KH1nGpWb
r0a9fW3WbpXKZj14Vt5AoA2ESRjsgvSBU07yRJPv0tUGUApfmgQgGh8VSHHl2dHIiwQvq3434W6u
iWRdpfaMIC6ApbfxzMOFlyRLJhGEXk+7vvLD9l2duShV/EBvpXTz6p4NF3WFkBcDt2z8VIAoowkr
Kyhjn2iae4bhjZAaiMCy6s1Dowqa7osPVm3aDDSuUjgXtt9F1OmaJTImCpCaIPUtvudAAu/7wNkX
I3M1IbiAj2fdwqqKJBAtKrfRq6bB7c6xtMRoQJ9WUXjrUAgzGMz/5+OHI1xwz2OWIQXo5v/aAAIL
UxH3gnnCbJYYdwjVMAT2TF5lAk38lxMhRHhDvlYQGCepouENBuF2mYqqXk317xZo0XaFD2OviuLr
VwWs+7CYeAQw9NweMLCX8g11YpJZMXKRQmvTpF1y1P11hxD6xaO1vIN0mRCVhciqbeLKo1TpeVxF
1rmhuL77Hbv8II7BFK9oNWnhicYzn/QLWPNPrjJFrUJQluQFNIwtBYf2iwwJHO+aOZYsPPE0TDnB
vfccSGX3aEO+4tmnmw53xj9AI/74YwPh/SiMDCLAmN1lLaAI/WI11QqCpTpSEilWMUx3SEIIovMM
//F6xWxAeO7izUXNOthpY75zKVAqQsVfaQ2h1qqDRwWRkFO9kFQ9NxfPaVqfYXLYwLgrfxylYVcN
v8HLex5k4Uy7Wys9ZZT8c1Sg2yrc+6n1UNg0IVQPuLcabK5j1uOOZ0Mwl/9Zj1ojhx8cftnIRkpH
gTcoL1jOGQ71CJP6R69eI0SBVDli2s9QLEQtHeg2bfIMImbOyUZpDF7FkdStfTmXzcfMvbBUDokn
pXxpE85UdkRcfVKFecBs3uD0WUEFV219uMroaHdaGeXwTjmSSftJOWceEUTMUtluFSG/g19Y2U9C
SPMHKOdtVHsO/sm2l5xCAdrY1iRSLI3bqO0IZo4Jbmf1QnmHfCU+t+IAtRbgXRt4OBJT8EfPDVNY
8o1PuKkXTLbeScbzGnkEDE3+HoAsezymU3DKhsArxTEtV7xFfE0IXYWlAChPBSkCHhe44Mf62Nih
NgG4JHvac98kjVn5VXGarOgclaBWFBszdu7hYLGy+Ure1NiFzDfNrJhVA9VondqRaXoYjvn/ggmO
4D64dyd75yctL79HIJeIwGP4rpiaXgIVcwhHcd6PHt8h2hOAf/oM0NmHJ7tsdjNVyFZWifJ7PFJC
33nyaV0WTci8+WzK1ipuxe3u1LSHUCU8ibD0FcY3jNak/xFKgHnr1eQwhi8eElT31FQw5lTEDoVy
RIoa/qoYNdUjB3ooeh1sGk/robytU6pOl5M1t0FcN68NVxWkm+a4v3aCsZ4UpJl4v9myFLJnzf5c
VMjqhIxZXN0HEHIc3ab9MwvMijn6gR3KU/4AmLB11Oc/LFoVUQO/f8Pwc+fdzBRX97Hik0Kw7Rtt
VwAmy2fli5EUkLATeuWVp6GwXoqJEQRw3yS0Amk4p2eCki1Us025DK10lc3Z2CyPikd/gWVJ/3Yr
+l5Fu9fF8zvHj1KY6fFhjRwEOA+lgadfqkNABlMrfFDic+JZqU40ze1g1p0fjR1qliObY8Ry7Ykp
mkixS3bm/DdYNdHr0rj3OtarLBmsuhb1gVOxKsMfITuMkWiC4LeMIq9/esj5eB+5Oc1Aiun+qzo4
kfnN3BSDQIRtA/1bUmpRqtRaqSmmCmx/LsEbuA9t5rTKV+Rp9n/Go/y/3N7yUoYkIUjBTt58boDn
cfpUpvDvC/5mrouHmICLHD2bq5YqeaAZwIc+wqzdziFCRpdcbidSXGXDsO69obl7QQ6bd+1KI/Mc
JR0zfmGTbmPI2+ZqG1oDIp6LXr8VIIs6vXiXSVthM94+bmwPb5sKqz5XSpTNN2NnMFP73aNQpYGT
XJCNfhpmNIidJFanKQKWKJM6ukzoMoXh0GNY0CL2zfRmCs4JlwGaw2PeNllsJLF2fuTYE0Kk+Bav
yg25yha/nINcTVSBYKH7dVfV8hjw6NOwch7fZ/XdUEUJRjNr8b+Uz2zfmX3kmgzTkDZ1GOYCJr4n
J8DmfHHOBpR/MmxexAQYjt+dLE+PWlIpGvJ+bNyZhaALyBsYvX7p8aFImaZyCWcqEgZWso7piOLZ
ON8SQFAWb451t6XlJo+OPqqTjd/RPbAIOc727h+P7mgLSKGkKleEFNcPf1O9nnzh9EGwBMfBUcVh
OjCtgsAg9GgTJptl8DryGvdWDuacJaXwBah6zTpUn2hLli4WZNS4wvWVfvIOaYk7Qyz28BQmSbwg
zITxyH0TPSimGwgCOX+QRaqGZxZAofY0Owa0sAC3kMAJ2EOiE2dxZWdoUAdPrdzRGuyIQgMnTAOh
ChU5MHe8qrNuKfyhnmHxY5UeXOaW5SaDMw4sm8IAbBbEB57jKdarIqBj7+1Fv4Uj8v0sKn4Jx5xO
ryTJbvK4aPSvBsJgzCCYA1BQ9oXm9/hV149966B8qQ9DhQm0GK9dnWRe8bPqOdxEL3W2PxjYLlAM
Dio848JoRdNrug01JxYyeuk+G2xrCNFeTyue5ltOhabunGptyRN7kWZOpKWtJ8Ym/JvUoAcad6Pd
Ge5Vpaqj6dF1z78N5ZR1sjuXaBdVwNaytMPKBN/5jfNzisS9Mqzw2sZthRbdpI4JKKKjG6lpddT1
5hYXhpg9CLMbYkaIJ72bXNtRpf3G1e5CkvBzvBskifSG6K1XAuH2B++p7TT63BBJLUGMeO90geYD
GY4m1m6hfDD0wej6tsEt0QMCM3OedgV5BWP2XqvMkxij1IJQOFP6iU0FcWarWJhVV/aqk8J4rZ/Q
+So30jCpWgyGhQ7XtB6KwLIpPjSdQ3SIYAZUSMnkTzUFf+pL+Po8vLUnqi2fR4j2LDG3Kz2zwynA
ABQEtWcyNLwh1DH6Hnv3xHShNnfOhfA/NDXHlhAyoq+MARxdBQiBgrVhFldVC6elyzToWCbYsUUq
nKDWTHBUx/f3fW7nZbsQU9tH61m9xRPg3LzjUBHqZ3lcD6CZiMnRDul6hxM2wfi+J+yugvGgMwnC
8p0MsBzYvrVWNmv/3TeMIQUYWAx2DCTycUzhXvLgCaDFuoqMxGFL6faOsWPR57fjBYDOjunWm+EM
CXwtTnWozBR8QF2gF0/Bujyx/yCgvYbcaeynBQlxiOwR1YBZ+JWVbobtNYJGAttS99z8uJ1vtvFc
UPsVG+h8aNyngVPR5lPW8LqIDegknjQY902JAHHaScdH7uoHSoeE0BlUDLREwxZEE0L2vHXh5U/c
RqefVoNP3+sHK2PTQkstbVBW6Xi4usleLgcQCYa6kaIWsx5AN065/9M7UBqtoiahKy5USjrRINpI
deJfSnxcxbPKTBtPyLaVAVbSMTvxBgm/YtOGHIBxfv6Mgj1ba474WJXS6K94wZygrNKdblp4Q68+
kkEygNTk+toUFh1K1uB/KvROTh1yNbl59iJd56yAlcHpct0Yh14YIsfAQX5U0vw6xy2HjQ1FflXZ
toheycLKLvtJL3xq0Bgm1IWRZWNyNv99nGXVpZoaRJWjExFM/1l9AYmMafaF1wrEwjfo9LLWPBSJ
DfU+B4spSiK0C5ZZ9GfvmjmBtN+2De1rc7fpvwq6oNlTl5UnoXBC/C9EzMEoS1nOxH6NPM7/ZwvB
9rF+LukRZhx3eAjJAzMwSh+29GtazhDCOBvDLN8ozzw9vNwgLvjAF2Lce+uRDYy8t8Xmgdkpt5ye
aI2nI9aUKE3mqvWOagGCKa+LbEs4jpXg9hUQcKmsSBihHjyjTH7JgLreupKTP3Rz+IfuAjkRrCwg
SYJM+A7pgDw8mWHobLLl3ndhb2OysjIa1IfsmBgU8AbE1aTbbskziMs397wz3KvRi3Y0qVEylDvS
BVLSHps2w40c2xE1waC1H2anb+o4fZMQYq8wpc/vr0VweYwJIN1t2d/RQ/6KefftytSov0vMgF8u
pAPpEguZFz6ly9lH/24BAN3LaP4mKsTVotHZnyoOYiISFQbYEtQilGeOmMVzSEfpz7zn2gfUb2Tb
E/GG7hieG7xn8LakrIaEHqI9zEBu3avK10hvJn9WuKCCOVz5ZWAA2MJ7xkBnk13jO8wiRfJI8/s9
oj1hpdNJBmiQhC7EfJtPipMiMqKimxhjutQ8GybgrHE862JBxW2TuWC9T4mb29LcHSpFLJPGbF44
1mYqO2unbPFdzcJfNetEcF4tZ15hMmq8t+XfddYnd1o1ZU0oseNtNqGVvos9JcBduoBdYXElOqWY
u8vHPxIkxkdeDn3+tlJrdOgJ6j43algqc8HyB7sPCV5fk04UwfLBpKiH44eh6vY91kgwSg5hyGhK
Xyjj2URKtLZN6cOBzIafAwdOGldp5VcUZu7zQ7iP1TDoDh8oQGoSFzXvN9mO8fQ60jRI0DTN488a
EwH0I7falyg/6yfc0n1BEHt3kpFQgAD7INZhx+5HFk7kXCu4KuS5NuepphGA513wgnVLx3JS6A/U
Hnzg698CjWauAl0lWmnPfHGAheAlsTWjQ5iu0Ws5giJcEZvn28zyG6yodL4yB6/ISZjJdcIRaX3R
9FqL7w6wDtx3/9rxjEFjJqht7+Pqt7yMkvlvjBTrdVxsmUOorDjCKD4W8HNcWo0jgsZYVDjVPn/7
qOdfXKteFvPssL0C1g14SFgOU20rqkaC3HpmCgxfsgZNuDwrpiVwazIKZf9RR7/tUZLnMhPwhUrt
i0ADDSrnZbvp4vrKG7/MyG2q0SA44EPWr8f1RgQW1dZcp62Jxr9W3C+AfYRG2I33eNYthFQzOvsO
SfxDtQUh1OkGpTW8lkWJbiIUdyJLogqIonW5CE1wmbh2YtkMqmQRfhi0npR4+1YAQUPepZSWYCfD
ulWFKPxVg+hyJuvRQYek/mSBxtZdAtwlwz6knxHF7Cm00H9ENOxKnnOk1qHa/feCWUoNcm173bgt
PgMX3gV2hkbvN/53ONzyc/7d7NXcFEuI/Q9dBunVtOrj2IzhRZV4dxcFuSmge1vFBZUhY2eFffDK
aAJXs8JxTB0Oet7dNou+ZAkcH2zmg7Y2DaIQ3SpQvpzVNRDAn5ZWuuPXZ7HwyIEsBwGURtw+y1jP
32jX4PrgtGra+mfZcPlIH4L6MIHlk4UxmdS0+uYVty0AJmNKcsJOPh1xV0uFA+6oseOY+93gsgH7
RbsCiRH2mHavzYM/e6a47YRjI21JcG1v6TVNynWBGQKO4ktMxpVEMqSWQsJcTPDN+pA4oymf328E
CKquifTKgpFlLQFaTmxEzQfuuPoxrD5IBmPo1bXb3NGdSexgrtOkv0PVUY8K3302Fb05DbfTinz/
Pusz3FHGJQhj04JdrrNDKYHK07MhkZRhhjHVii57K8EJjkGnlFh/1VJesj/9y6BqCnrwoIJdvay7
nNgZNI4rrEHyJwEZBwgVl2LqYxRd+iBWTinE4Dx9iYEI0u9hkY2k60QZh0fi0oL52z0SISyFegRb
Dewe+fr4EYu05SxFUAxOiEGiSdp5tAZZkXcg4ZKofUJnI3Yhs1dZgG+HmScLQnSKe6uZ64aLL4ru
8NIXRahIJsN4GFhMU/O5n4VNP7qKO+sxfz7AAeHfxmmwDUG0STYMrhMxHwnZyFYkhEq5Lbj2c9za
xr2bVj9SEL7fP4b5spOe0xWdK5lAvlrssQIbxfy6tF2oF+aLpTB1mtNR8zPYO6lonQ9l9g9DvcQr
wl7xD57wMQmalGrZtpqbHQCvesg6paNm+jdm18DkDm86olGiuMHsXUI9ODQq6KFHYqtUyV+xTL1E
Sc9Qh+EvOfktdTerXHXPCs9fFRzBRfMudT/N9qlFKb4Kmx9FjWeaEEyooEoqmp0aEn+aw9FwDo5d
hKuiKFIasHflm2ncL4lBURl482QxkYmKt+dcRiOGgLzHXUbb/788ydhpws3ws+lCy3BYayqe5kz9
4debbBEmcISvbBqg9xxJ4EAPpUpzqX65ia+Z0WPG1iBd7JayxbtXMwhMN2KyH5zuckN+6SKP3Oxm
Vf8z55gXzPjaTZRPTdA3L22Ca/4ZZxN/ex5+j/zd8DDYTn+SKnx3/gj64d6F98lxMmNtbpRa15nm
/mk8xx78u6ATD2KgUw8kB8qHOPkLO0DP1/1PJtusnPF1XibUjEMqXo2xtiIvewGNn1O8Zuo9M4WG
2MjoDNbHEqfhDI3oQWl3v+lKedEle+mOGBCeVgoFBflkv8//eXzmY70vGlXe9CGNhKY0U2JF/RbU
Kya6k12vwj3c7zaHKA1/gNeqA8chSZ5oJJikZAEUSJJbJ0tup6LeSLSZ1WX5WkYz7FQWev0m3/qJ
FHdUrEqhs56zPgxWHetx/T4C6qiK1WnEGxBAjf5/2GSYgFSfSTZqI1qLzcEwS9ztFe8mw7LTTuub
Cy5XZyZ/MTnBSbzR1eGw4wLjr6UIr/WvBY2Tiz+kiBxFSxPRVNOHlCu4qHFodFa7/yH34bFQWHeW
wrzZzZ/L7cKUv9cg3MnHdvEIJmDYuRNHkQgkdZAxOz5FgBd3mzka88GUfB18euBnMR7Xulgedesf
tJY0vyzoJi/plMiGxm6qDaYBvHkhPUYvxCORPzb6wmFOKeV3U48n1lB0pTO7WoTXpFXFl6Pl1FC+
jo8w2bUUyIaPFqU0ZoxOsJtEJf1wQIAxdLp8klhnywcmxfXX421v+wyyCvxEvFMIDvXuDiGHilJB
7mnba9bBUQD/Z1Wy0lk9bB1AKqCVVb2/2W+e12jFyg3TrREf/T5kXAFt72RzSbQ59bEXO0XbX6Q+
gn9WuWvlQDgVScqhSqvUZm9cGovZj6vyP1aVAHOaYCf7DVCBqVAkW7BiiAILkqKtxOYhQWLwlswt
Jk4E1+mZgO5Fk2K8wPSeM6yL8P7JYAlHr2YAywmmSB4KIwYqNr7N5D8fL/oI50DMCCAToicFUwBP
8QBNiysTYNAaGZKZwrmjHChFlgg1NqKdjF5AW0HZ54dhLiLwVLdbCGyLM8Odia3DKYXhfK7G7Znu
aTHIC11izcigZx4zDr5+uC0qzHzLw6cqAZcYwFbGNI3wmfV8GKprOxq8ZVEzl+6mWHNHGvbTxJ6k
0V7Cj9b5pg8ICDXkJFJQi7ngLOp7lGawW13138du4ijobc+n8AtjF3BN3oLtwx4X9VekR3cvmYvQ
jvz2GnKPif5+uXKbaU3F5s5M/Q1Y/vo4TS4cjYCAdK+Q3bymvIBZtSjXemrkXLg0LbaqETe4w6E7
GZ+P2sioYgBRX0RsCv8iyw6TYE7e74+TsCpwBjsS9i6JLChpeP2cE6ccrOeONbNs4Q9sCNOdY/xF
JmvjC7JC45ZHmQM2u3ZSfhmhz9kRnCjvXar/6qaUQJY12h33YioCzPkREI6vykp0SpILEXqZSQAs
Emk7ATaUzSbwtohZ3gbPph681tnKWcU2PYZfrPTWl1uFbxnX7gVOZtStBKwQrfZs01myEvxTMX3i
nsyWVKUXaCbH63ydjC90fSTRAM4ACt00vO/NAB14JFr3AIoVnRYML6bSGr6t5xObeHsYEyoreyMv
l/W64ovBq0pT/jgs9RJ8t24L5dhTHJEkthZUj980Jc3wSMERSMYUieyjCtAmE5os8S6r7pOAKvvA
uASiw1Ec2koTAhr0rlIuAs7C5GvyCiy/nWQIMrglMWErn9KfjG025PrMNdwAorEZLset0mYkDZd0
Tg6c+IlfzAJIUkY/cWqkyDPDqTT5sOd6GBeQdO+0xp/tRCz/9s0wdduYIrAS/dBQ40/dRM25zJHr
QOAUB0iBwC6cCPwS95CK6NMXp4j/haX9ikFDfKiF5qzBx2TOoLadtjnXNEMAZ04xc8yBKS4JLGx9
WIZfLVMJjB8h9iBdZBxggAD9F2XTgV8ZfztHeIa2rSvKc0KDVeW+ZoWSMvca+91sXQkBiqgNftb2
Yze275AHe1VkHYN5DUr0KcZZr16cHnmBsQ7IeSmETeJaqiR3Hu0KXnZe++HL9BP6gUPGu1XfDz2g
gwgrxgHBKMnQs1aRd8fpSBHAOwZjQ9V9gH/F9SRXS5HgOfaTpMsF0xaBRD21QsdGugDzaeZ9heYe
Oyxu5Gf95ePx+JC1oCFBMNo1M5tUfd/pYk072QjUv9KduG94ADCBZZ9EGF9Gv19cRrt+yR5c+E1L
HGm0FmFG1e5xOL/vqclp3aVuG3wuHUVuHpaaZKyDS5+xkXX84iBD5+/2vxX8sf+ZM4OAgkf0QHy2
nr4q6qL3xzv1YJZEkdL3VdPafVy0yx+9lBKIW7DtPuPpJm46KFp9J7QgZRGNbox/U3tSZ/UPJ0Ao
07sTlQDd0yGPlNLxeSBLq4fP6C7mx/RVxu+ZUC4qYQBlE9iAuhqgQWCruN+5seUbSFaL34GxoOVb
z9p4sTTacu3snqzPjPqlGqNroumdoxAqgaS4V6ZWbX+l4zAmaQg3c2IUYx82Bez1PlaT1kfH/OJI
FZH07M6prE3QZfHMuiJpJ8Bbx0VeALFbsFz2SbktOqNHlBxN3Ddl/dmFwd6LoaHX+y07xJZeNp3E
qAsHJK84BwJMkJJqxtoo+7auPhbrjdFzOqp9/C931YPxnqlsLHGIbXfIYysdB/5WOZMfT6SkVH3+
WCnAaLz1FApk/+bcYRNWiR0L1510Kos9pjdBU5mkAZgkVrCTFXzT199+eSXV8uvWsn5lZ1mWmX22
J1almOFWyuB/hnoG+wBZua/U40Xo5BsHNK1BCb2E2zqjtp6isvmtPxaBDYv7hdq2nu2Pv/0gerWZ
vDf1BLdf/TMa5d7J63fQUEqH3BgxkzWUCVuO5WSJGDcbl4F8KaLb5ScgzugU3P2d2T39zBzQb2bw
pLI3MV+S3EVekWMctR0H/5tatqyy3yB/7zlezZsRTzSYj+Sea52KK0dJMLTnBXqt1h0lap/rYY3X
SNXmvr9x4QHc3vFS9SOj6+TetXKR6Aq6k1o4kx0Nc6IqCyMO3G5ymVvGhgus0Qk6jizniY0KmOPg
I7wBdWMdromyL2YEfZZ6ALwqdD71DY9XLybAidLXhfP3hnWdPmWdEUqibxsOGmxY9P/Td0x0n3n1
zTWnavhNWzB07ZNAoanIs56aPmxVrF4NNO8KnxXNwGlhZVc1cvoRGOu0+RoaLj+9pRKyRpZcUgOK
Zt4EaDJoGgb6ILZnrjkqN2kW7FFLoRmyXWAWNLLuGwhfoP9nyiwiblrJ8fOY498I51yZBrReoJc2
jIB6kV43x+8w3iHeEU2DFd8zhmY+f3aeWH+K7fpQ3sjW/e4ofhjUvAsARcouAU+JAB1hnNXviaxB
YPntTnvv1MBA+vw8n6fiIH1a/lmTfqpdFCvNo70VCSsSIVwT3ohEl0KoMFvd863IxrWrQo+HiFK0
5gne/XJvnC9WHQZSeAsUGONqRX3gEmPbqawv0UgJcHx68mImkrAByczmkTH/Cewxa3HCHQsTqYFi
QhB5ClewYYcKOnR7oDptjTskfy+oxGRqe8KlfUcncKLI4Yh+DJwp3CuL/lWJTRuoIinAbNbY2kv/
vu97imkbYXX05Rac9GHG5lP7/NTmalYIZUPeWDrOrEjyvDD1fPNveqFmefFF9di33sGvnMEFo3o0
APLu6MXEUtK7qU4M6nPzusKuW11rSvbWoN2E4shHBZqwHM/4BIT/qud7R7Ui3J/JVilUf19HeUhC
8EMbse8Xq19Zo4xKIqEGKI69PDW3NSyf/PYMpCfoVCTnTqI2VhExuslG87dA46S5HHgTSRZJuTF4
GZiDQ4Zh43vmOfAAIbpOlOiE+ROGnmnqoc4lNLO/mG2awHrPfCTaoUZaSAX273qcFnc14gWSg93p
oolR+TzGEK3mmmt9654TXofJNNRM+L1RvdRnUznYJUiPC6f2pIZcCBe91BDp76E+fiH3AVVEKClA
ByfNbgVf3Jc9bkiCVUB+F/7mIYrgk2SDXqki+1jA6QLJcNjEv5bVsdeeyX9SVHx5gtCQnuECzLnv
vWWh5/9favLitgQzAxxvRPNK5RR5y4D3EIKEVktAlyKs5oEGaltnyfT0BuLT4Skx8C9Qg3a0YX9x
lDfnMiCvAbEvzFMRDbJV+xnQi+vN7jtwHflGzvfR+dRY4QeXAFucNiYsoVFVSY1nyLsMnHSyhn69
tYF3lIXTT2iIGjHpvq7oi+pENOsbhvWSwq3EHt+yL4bzxGI9HVIHNjIPM+g/uD9mknE0xh0AlwdX
ANTsB5wXuM4pHE0xiSq1ERJZ9ALLLGKBoLNOZXERZBwr2+KGa7hYzF4aK2Sjllw35Fj0C5OJzk4J
vZYTHSy3oJ3vZL8yajFiaDlN6qy5U6G+tsHgupODIS0l21lJnxQLwendzT30y/dN1L075TlvCsqA
sgBAnKaNr0Orx5FWLSQN6z/dnGzkBFLFTBXSVx/srJ+Qv1dDqL0CUHny48QvF7Z7vSjp4cFTe2w/
047CU3zgEmHY9AihezBiaE9FA1533V6ImIJ3l1DRlD5ydLC/UXH0U0Or+AF17h0kXhHADn0oKkhc
FwvpZ49mcQBRgYi7r9vx8V55M+dfDUA81F1yVFVfsnKzm6IgZ3mJZr9+jCQvvkQitAIY7Fb8jGDd
CmBx6seg2PtFnVD6xPqhUuHbyy0GQTlt878aUKXE3Z/TN5srcGhaN7BTs+2O8754VuUpamiPNQs3
SwQHk8LrMlWNqlLI71WLB8w/jdaXwsXrnUswPCiWdjFGKp1K3twHRcJ16TTMmmOPiorLigsfYgiE
OZRhaV17w9G6/5p3MtCs/ML9/0i+gaVkIXM00KVOm2VHd8p6kBqZydQ+EWKzT+xKQjz8asSY5+JW
ly2UHr6iXIDZqg6WV1CgdiATYOk7i2oehtUXdmYC6Dd7O7v+99quTy7zqbVkMXiySSr/3sbbkEsP
7hYpUCZpxbKFj4Iy5sLklQKnIWt3CqyWAtS3xi5BnXtGbHA1Icfi89UJB8pYwbO9TiaarqeZbgD2
Phs2Gmcfs3xR5eqTuOzIgpY/UAhBZ+X0lGPujxSjNwHyswcqE7lYsq+uKNLhGZ5BwunvNY3ItKz4
C69xtoQyBXLRNN66wZVWHGP1uJYim9EdfN+RWz4qF1vlYYo7niWtxcKO78EB0seVFfD+DLRlhyw1
N0HOsKFTS61RdbVOLhTuGRMLLgpCrGvc3gh4DbYhUs785Oy7fqNVSP9a+3+7RJ3QAmIw+/IgLWfM
VbflNZV1hl8MAOMPwJt80WtrkLfhRAX9Qu0R32zSRysTp+gM/hWnyz7fIYlCk9MdyGgwyb0nBv6O
jE7lhg+N6uHWonNtjNnGAgSV4jCFMIX7nuFlUi2ZCwmtTB7stOigInC6bUa+tBtGBPIc8NqTOPix
dK6JXYNP0Y9otgfcdZBD9di5IfrWP2wnsLRAa64LMXXX8Q3QBGCBjn689MxCW/Rq5GkMVeJkw+i2
NwfEbBD4dPUOSz4zySYgljC8eRRZzjHOFY13cbYAOexzCxnbdsMFjioY1n+ETRfrBhAJLsDpenXk
Uyg1NZ2HFJtGvQcVoO6Z0xGLnzgVECyTl4ipCvbhtdDOnJ2CUHfu2wk4xSqlCt1jbuX4Aj1PfcON
CNbnJpTZZb0u/55bNj9QYrOy7llntMAH52U0NFnaGAA69/wOMY1a4aJfY2XBwkgrhfqH3+CEd5il
SO99V7UdxoyejvoRbm/Wl1tsp1TYpq+g/n52rs1iSwhoK39EzEnAnPaqwK4pwUjb78ysFFN8wkh5
simR0jlFcRr0dvNVLujTU6iXguY60VaJi7iYalgv3nKN2Q06Ct6lZea3aK8Ynz4G83vooeNtl1Dd
c/oNF5/iMY5tG6Bw6t72aB0UzexC5ZZZFZ1Wqg3Vqedklq2+TmdFwywVMfoICgD5emizqUnUtOgg
i8ufGx5WEfWjk/PF/eBzqg9on3EPYkH806OR4jvmhG7M7qsm/WyBh5n0nik8EdiuXHd+Ty7pnkV4
/3FANoFoFMiMz3mvc77XVzIZmYTJhSNow42XRuVFiHQjpuFpvS1mRYrAU6DzXUMNymW3vx+dzO90
CZWK5OOAOfPI+aXu7QPHfdS0+mc6nT/txtKw1fD+HQYxsrjw80QYjZsUe13ggQhSM/BB0XD38Ix/
Yt6X9C9a8se1Meh0Ny6sISpw9FGxhhqiX4KP8cAJ3l5whW4tgzwNIOAoZLVwJYKnx09s6Y3khMBT
xSH0GLVdqRMGG/O+Rx8e0UO2lpJ2HP3kAE7GOyRWPqNXiJciz5culyKW9zS1Y1MC5h0v7jvOeP2V
44+ukxpsWoa71wodzaMCO2308Kf4bWAqfa8oREO5dMj68Yogszwwe98nrdntNHGJ16jsqJ9NhFHU
ke3mM7AX21Kp5PeTlyazMG4EJm7dhxb4/nwQp31ViqHLyvhLy+tIuR7zAZT/etcZWP/gan9mXZqb
c3ofzQdCgH18ffv5S8VbAASWR8K0DytgbRszvswmJZdFCyWi8zi6R47JiX87UD62MOHSo90YMkhi
o44yZaMs0r68xBbO+fKRXkDIslCbvwbwtX8PHPYAuijqbA8+9ZHrFnIeaN8kE2IMFQFnFickWW8O
+BpxRdFa3baKfDu1l1C93kdzPyX+tEIDpYcZx1bFEXs9higKfyTaEEyvBsidggZgw+t8n19yRIf6
g4AYca9NTQq655ABC+pcBYrzLLXm4fwj7jT/rSpLKL27bL1aAwODotuLaig4SPOQMVp6rU17zj2x
6TUt1Tl2XSUnaMzi8ADYUQedVYKc4DtLzmeFaJmmCj4F+yXoy8bne7WnyijyLQyxsN9EXspeop7K
4jWj20sJGQu5aQtgfZDri3Ikw/pCFka6bnULQnm7aOkMr5gWKzrLcp4hFPwyKpAsD+xcLZncwJCR
APAWXV8+CUKgiLU+UtNiMc0ZbCoKSV75fh13xJ3o3dzNw0wAkxSyRxdbPlwcq6HUKh4xh4i1rFqI
/nvmpG31cnkLap7ppw1KtTsai7JCktqawDPCf1aiYJBlfJjRonF2vmlk2JTLFFiusq1NOZPNX+k3
Z75Cj76DPrRRnEFB8s8RuI+Hs7KMWxXmH3Xc5bg9SE42oRvqivFjU55lYHNSzHqtnnsPcMKzdqif
Kbh7/FOR1rXpJ0ZguoWmffFed0AaMrb+XnAgZ+Ji302ZeGCYae0Z6abi1Tr5aDq38CTpmXIbmAMV
kma7unXdqDvxqDI7KpIro/s/AWqDGzyNHYnrUyc+3AhKUaaGf/rwhKfQdq3QUWAUohZWIzAJCO+n
JaT+HnLCDR/1zFq5oBKpH1riR4UyIODXI3uuIJ6knFBBLFwdUhmRgWOXKcHmvwarrWi/WbfSSQ10
3vbnD+3HfAYmPIXxVfTE+BseBVVU8VrgBqWjf62GfZdGDtWOFWgiUPd36AZ/swcmWUL5aIdDFYrv
oWzGvJL2U2cFKbb0F1Jap7160LCY+9qVXDdSx1uUv0C9KQyP1XYyTrK88untQNRipwl1KmvWnE+L
E20SabeNAnG10aGFvGr9o6sm97nOMyAEUpHCm2d4+cmo8voPRezQiZRfTz039fR0R10tHbjPvId/
/SjsmW1rJE7J5QoFOObZSTDFLCTEXQzI3D/DjdNL3515NGPmtdD+JuE7wNlGVZ5t3PABKUupvTf/
Pc3PNv2Fa/6LcdJ2dTWgqzn2R+DIqMyQENZpPge9qiE1XeNWEqL84Jv+h66TyiFYotQxEiW9RYna
IbKw7gcT/tak2lLc4ssDuQ99TkyC0sb9rE1pP+d4sWrEQGetZ8VUSvqJ3bJD0y2xYOSRGzLmt95e
/kGizP3F+30tbrWg1FbenODTeXEn90CFOunSwbOLnec4HGY04qo05YQFAq0flidh8OcVmg9bhvQN
qiSE3XFCfZYr4InSm1R5jbSKHQs3etCXTNtynZIjTsQwm+m7Hf29OXnJQk+VaEs1dPTS5VoeygWi
veXJifMhXlWpP88JYYTbBbU8ceJGDnl82CJxku7eiGAkG5dBlv03YettTaG5zuoofMFTYbLHoJye
2achIVZtAiqiqX/qLBs1uHRmXJXfgvOMy0zn37kcXYK6x+WMqFFel45Vh4MEPuApgWYXSWb9KNvh
gxi0HIEt9vq7Kajj89izbSeAvBW7xJ2fIC7KbUcxHq1LKURyWDge1W6fq+Cu6fvM7f8AtXPufpcF
S92kioJmCUZ+77oE9qmBjWEtcP7oBc9AAL1thn6fV120mxzFevhcom1woCoJlO6jT3krdVvkDdy9
Bm3cmLmnpU2fZX618wr65/YItb+7to5bAcx59ri7mfmPQhaYn3ASM395xRkHoOrysh+QVSK/xXZK
WXoqdJVeNVN7M89whdE5ycHz0p9S8ZXyknmeQAnhThKjlCBt6pyZd/U8bT4zr1giAWs+KcOq7A6e
ppSQwS1y7oX30V/1VsxIVlhZjlpT7J/XQ2gtA+Fx3m18MRio0a+/2q9IDFMaJ6sSRXB4pe1sJNiL
i7VBC4MIC0fjnx2XFTTQyHY2upQJMnFxcQ7FclM9eaX7Lg0T2ULxNH2EKaPhMpSzOZnlRLzAQ9wj
q3gS3qU1jIgeZ/clAE4DYZMpsuzNi9p4Qa1SFTgoYcE3zGDTA0VFmCbtXcz2MSKhtP9+p19kWJOe
chIptCjn3Q3JhDeArKLGrVQJYVfeNTcGtjYT+L5Ae6hHHgnuR9neiHWLvnbyIujSzW7nm8eLcWyR
z/Pmt1pV31HAjeymnj1Hw+TY3TFdrKLbyY49cE0bsY+CSyozzl9FoIkBLUcNTiJK8muKofaI8zWI
zYdHJE6yebY27jyi0V+rvaGrQ6WA9nP4GRoVBdKQCaC1X0c/CZj7QmnfVDdj5DWqreyIA7qBnWiC
IiZSVfJj/6MMMDMhOGuAcagS69lkwnUWKBpCJqNr7wCmbvEubNN0NmUdtdsqClbpO0px05gUuhHK
JmVXiWUa7INVRnGu7ZRUzPw+Z2se7a0w0qGPdkUSzAC5Q4EP+Ij6vpVzFvWNT3BeI45VjN5wNndO
Zv1Yj4Ua49zYo6I35LwFru/g5pioJw1SY0+K2EqLUYREOGREwvnWCoo6/n7FRCWTQUxMkF7WNF+9
vIfwbzQc0r1ZqDSOXSenBxMOuEvMgEOgl9yHRdMk/VSnjknZIFG7IEszCM9l4pxZsIlKuSSJJk80
xtBTZ9pWJNiKZCVuxhZS+Bjs4LaDj7nL9/PjO1skHNEFX0wV9ns9orLffLzX11UDMYTidBneo9FD
l9QIQ+SkLLDrpQfMjZ6I41VKr1Y7zMjaZPtP4b1O9j0lyqyt1kPPXNvGrqF3Obp4AMvVIZrurhUc
LwiQy9MOdZ8vLnoFweoEs0csoZiSl3vGBSo154iLNmnWutPEhJfpTDmw87hlJX5qClQ84q1uaokp
V7oyshkIG/O+/ADHoocfrthlRt9xByfy90hkhqv9BypKZbd0rCX03aJVIRiYpZjS6AWJQAz2r7jO
WPri1V8NfDVoun7nXP9NmgKFyttct3E/cu/Mb9Q/xGWmhSbgZmzT6tqv7md2ehJFQZfY1HnCK8oe
ZNO7GbUFXad8XpnZPUIeQEcN6fQLT88AinipdiG/8JdiMS7nWnA1Ll+OSMAms7gXYy7mycFIZPuf
2GmH21TOL9f2d1jSHUeochBwRQafC+2TmdWyK/gnvw6fblUpqSmlyKsLFAXqXdivMgzV5R+ruHko
DHRTPe5shcFvwjB7icqjPRQzcMAczpjsJOKJkqmRKNjKrGSfaMRF6W/GkDdxVC9hEyJ+6OLHJhP1
R51N5ieWsozof73I6OVoNDGD9bWx9MH7vKaz1s3Qnc78AD+kr1bc39/AqkMsAqRaWjYPpmJP0gR4
G0OoX/TXVKCatKD4SkgKxqcI1JUFW14f1CiVxjc9636lKeGnTSGvsAbQ+9mBK9UCNUfQPBg2uZ98
BptzLHp2z//aZ3ASQxw9fiGLXBKjoocXwgaMFVvwT71RsiLLUwnKgUcrAJB8aqEppZaY1pOgi9+P
z3Tf4enj1KIrBTT6NFaCPVvYizrKlRMCIXClGgpHQrcq0yH+5eMvDB3/7oVPHJE4ZM7ABow3ESZV
3U5UsVnXj2hxZ9jp9vDkxWh0juj0tdESJUlOMDfoT0/rUhmXoBtH03h3zlT1jXr+yx52Qoaxq0IQ
ca9QcgtDbEo/t42MZvEDbbbRJrqeghNKbFfs58I0uranpUrDDGeIsGt9QnpcXaGQMRjJ4HCD3bwC
abBPEIbRJsrZL65oOYIUCFz1JSIRp4RM4n3zI5otECVl1vSV6FFIQDp9ct1hHZkaZq9r4VJXNqzF
eYbIXu5e7FWGFGTpmFjKClX5GUZ5Ctx+nUqRh6qhfpLk3d6zmO4WOwGuPAPZH+xBVd8v75j556IX
pVDA6KD8UJ5Uz8dz25cTSYSmk1aaimugkZaWZrnpVZHY07Vg1CuNUi8hktcB9P+HIjo+/tkQEHYz
Yhcm+NFmPuvjtgQzrvAwb9zl1IgW23KgHoVQMVuaXwqEd2c3o2KWT5GJ/LMtzckVaBW/pC3wlPBM
Zw6jyD/ZVTPdE58ywH4iIJ/0xGZdCHhxVTnt4sJKbY0Cy2en5HrMK35zT/LM1O284xViUtM6Rhbt
ZXmlGaNAWhZimk5TM3d1jq36YGgzL0iEpCiBy2F2Kjx2RI3569YmLBYk5GoklSISVCUFrwO/UeK+
nUeBbofDHF6xQFnhCPkoEsLoFNM0Nxytdq9tG2x+OGIwm530vMSoW8bNJtVrMlOn4JpYMRpxlon/
vG4zZFhGnVk6mLdBeBDmrHqkHrUDJBRjvbbKJzkj2jpmXUUHjPFERNiHyKiAensPL58PvG9bNlQP
DtMdvBvgwVDtmGuRjsVJcnDGKJXtLbsUMJQKfMYJwzTJHcdkvwqYrrPETeVtU2t0Dye1UAN8zMjw
sEv950hb4FC8iB0THpoegDpg1ZDAU8GTwfvo3QLXCDTNxNEqintOaSnnmd1StEgLeOPJ6wlxQeBX
SOjtTxrD7HEOstdkfJcqRI6xDHPiXXOo5G6AEQahTDsjKfDw3G/J4SGg4C2hoUSuNjmjjCzXoUq8
Xt6LSSFHr46H5DLUtWz7yQlkDt4uzcjFdWKzvQbavBk90Bx+x0TOZdJuB3d8gRlW0bxt4BLW1Q4M
f/c2mCnz4xvnKQK5QHXwIcEQDkvI1FNOqZYngYtcnvc6qxKMmwW56NiojH76wHMCqcVCQKie6i0H
jrRE5oDFYryp51yc6C2BNlov4dz2jjpofmYx0bmxJOjhpl5mAToWe2FhYvMTuulGMKeBRimzZ36O
+ELaDPvnhy9YaRos+N+Ogb6QAns31ooH52mTj8L75YHa5t5IhqHRov3dZhkcrlyuc4Hg1mQj8LWf
DEIqP+/CHUQebH9a4S0GMfsDfjHTCXjTR/jfL2I/lMfmLFPEeYELWPxKhUy1C7AA0Di7+q1zm21k
J8ebOQpC/+oPS1BqbCy8bSItlo86JmxC7dHFiT+WaYpxPvjrDwUG7gsHG7OE3KqnWr+VE9bnAgEQ
3OnsA1tpGklr5hBwdoW0R7+KQkeFoxgflMO8IGfwX5MlVkY4cASC8Ti0xg4KVvjEsdt1YSZCwoPN
QhvOMRAuxKx16Xeq3P0yynC/lVFYVPOS97EO5eM07lk1U/WPw16gvoYtywBj4GFAwN8fbbpRyGeC
SInvEjzvjmdhkQxAaZwsKYaml/YN7lRlniCxlzCAFDflCnGiKhPQt4M5jLKRV8xLq2ZuqBGsSvNn
5CbLqAssOsuX8H49hAXxTQxu07oTkl5kvX2i3TMcdIUd/ETvl11afshKqBckoCRfQIHHDmGX85+9
xPmOlav4R7ZNUfF6WvY82BtefUyV+PG9nR6qEdEk46BkeYsE3Ry2S4+9LKpogiJa+Afdsmpz6ABG
Scs2fPWt+8BzNzwfLrkj0tUx4OxRbnPkuAQZAIhgfat3/haF7C4gGs6XaaYDC75hXC5KifD8hmkQ
dzkjRJhCjjU7dGiuKt536ZSCczI6upHp4az1XvR8O92XX05Pxv7OM8oxz+1UF/1cGWK+GqXCATZH
XIbObT3sPZcexjBIed3kERC4qrpzpwwObgQKC7BYhEqsMWdnQeXXvgysuJYEX3y+dIYm/Eiulk8S
ZvhGR9eCxnzLfaphdsXKjNlYqR2q8thXdXLF61CBr608kNRRWYsl18LipchRLCGCaj1xdFLsRW1+
V5lKQKx6F18lwgLif82cSg6Vg3PP0eG4qvoxLiOGfv8wSnfbDr//FQOsd3WJQEBVqkUeGf6MWrY4
OKIp7WchAby6jevedeYptRUcoMRa5UbECWSphfeO12CsZzsOVP2BE1GSnOjgqruGMLHcrsJ26deD
OSYSjj3JLDjBZuNfFRkUnrZgwIMdxYH4f2yt6qy1FDvOTB4aTbtZQVcSjWbmu5586fr6HzeWa1/m
koyha8+0oyLyPoz6VEKi4nU73yHfgGv91w83e3vviK8hJDjahtKQIyf1fgdeaIrewvYO87GqklHI
3saAerKAZWu27ow/jOZ5NEJnAfEHzV5UDvX3vtwMGd6sxYQxp4VW8RBe75ibzszKNRzUVjCT0ivl
vwlLHD2Vk2l5omYvJrdlnT3eUroM6hqIr+EySZdvvv3s1I2UCEz5xztNkrM1+te0TO0i5dozflp8
88KSWa21bulUYjMGw+tajFq5K9SbUfnj02r00CpAmC3G7VFR9tQtPW61ZdB7KDZWPF3dTdtl8LOP
ikSVUU89pOHoC9KTBIzAxIcaDQvYrcs4jWgNisBpMmcdfO2ivC8i2X16xqP3dZ53DZf/QMIa7/3u
ImdPxN9XwGD54cJPjNwWbWR236KZQWuS9UEirNurlXGCAItFxViNqQoegEsJbrH6ETMm7uXd2tQh
Z6+Oqt4zWhoLv8VQ3RxaAFdQV2DurHWzuoeiCn5/UUOmErzRMuDl3cpZWzcoG5UbTSW4FChj3ZlK
7sa1ac7+1d9KfN7wrpfflH8LBk+EzIjw73unrbwoihjNTkMHl2oiGdOmJa70gOjvXa40E0P8YW6X
1vUEhkuN9aKSn3PugjAErX2GDGOpHtEFy3MpD3iXKGC/yJjEVWdtU3EI7fQiTM9Y3HlyskmgEopM
Fcl8OswDCgRxot/svCmAUvAPL5HJ7ZsWpI39z1kfogE71bEo3EYwKrdiw588uWVA36nXlQree1j6
Q//tHs/FLSIRKNN6bJ9KspG8uAjRe9qN0QDW8su0E/VjLGJQFKRajikc5bgBup8/1zKbMfs+pJAN
oPLOdBR/9GIPLsieDvlZtjRJdyX7zFzgHXONJ0SUSQAdNLe/vHW03mEfbJARdjTuRZT5UftxQxD8
benVWaYPCj5aqARFAMG8aMXiJ+QLg6Jl0wclrq2JsEPhlBK8i9tniZqH7wy/Ng/6SbPDJfhUb35t
k7bSGI548bFRu3/4W7yQIn6JtyO4CHuI0IXWxexLsHU77xqe5z4Se3oP+j6I5HrSbPT4X84i8zm7
eTrCi11bx3QgkkFT+Q8LeTJT7o0d2IIJxZwWMakDSrijAUDYlt+HNu1Z6drUqeG6H25xjd1n8NMx
8eN/fdTpeoC+jtCroEEZySwBYQFmP9q/8056T/2HTB9C9uU+sj7e7xY0awjvgtL+IOhI7YzDuVKn
FLsUWqBl5jcFCzg4SLGwAJ8IfL/LiSV6rFQ7OZavI/9Aakq8dev/wBS6ifModsq2/BcE5DnUw+Uw
DazsWtjAdYqv6iuknlzOoa/B/DUsLV4FIh+1uMMrLyDSvXiEuNGIRko6OnKJ3jPia0ED93OGIctt
JQSGbMF5c/7ZUY5ncpkY1C4NA+N98f5Ul+bMvp1qpOlG7f0wwWRa90f2LY0CIiUbcSFDyGispav1
9NXigAA848+EDucOGamKEjr0oiaWHraMMxH6ENpv0cqbSeEMzJkLQihFrj26gsFBa6ZbN1BHC4+r
Uj0GxOIl7qaMs6ksXZrqqsmpu7wpslOGA8Urd9dJEgUtwGDvdTVnVYKdePXnNiiFFAUaM7LhqneD
L1t4p13oxKEr+kAJUyG8HeFPuce8H1ez8P9bzZEawkLL6C70cyFe138Dc0uP0tfTUi/lErnUhKvZ
xldkiA4WaZSiU9xChcIClNQo1CIBWmWaW9eY7TOnxrW7Ul2oWI2kZThXaKnxomlwj/knCWbLGVoI
e5xJ4J6rMKg3rldGqdfii4Z/GdGBQ0MPXHzZND59JMWPcBj8JZNalJeXE57vfQoL4L3mvk97qYXW
Ed0acMWSXCWYoYbVQCIfrxTH4Ce6fyTBbOTu93YrlN76hjLMFzSKHEKPuPUwxabc2AHf0hzWw0D1
Cc6cv4sOO+o/cAsm5ElYuftGZj790oYl1/zyKr4nyLigX/R1Fotas9fV5zRNMnsqExC4Gbw8BphO
qYaF8foGr0jsaOtHVA3oQk9nnbh7xyf8wNNmnW8V7/go+kEl11vzVkQ+Zp+jyrdpbER6XrBSVEU6
Q0TLaCr8zvLKuD18LhzpEbs17SwTi53x8tq3M+C0g1NkLonikWyZ5pu0/pmfUMktacIknLtdjPji
pFrPYWe5LbXVmUx6URDVDX4K5JFijXnbIeY6VSxYX8f/GcYbIxBmAKbAWCU3fnpP1wPr6QLcmAHY
8nydProPdhH+svAfIvBGds8HeXA+hHLut3yW2tdt7DuEQi7GVlvwW1uHGfXBqqHsqQv8Nx97Ym/g
uQN9wCVinQ3QiJWVWFUIWxkXx9vwsD05+qYU6mA25r7R+R4/6x6ZK7cb6qEDU7cTt+127s1QrscH
jJdJbR3/ymu21tJkzgPsWQaGIr/AdggIYcsCEN3gR+9/m9/tiO5elAc7UncbboMxDn+uhZVcie6d
nGDrN0+SxWO/UV2bu38rPolSwHw3ytoL/Q0Q3CIFMP93Qqti3n1JZudSG0H/jqlJw2OjvDRMhptT
tad8Gx8CVDXoIzZHIz9MGE5Jjv/sv7Of1kwgxBSoHYiYhZX3+4uK4JyG7vUfLEGFVxnOCsHmjYAV
3mrvbjJax9ja7b57pm66s9V15a+OYOffJJgYOD5bWkZKarAk9QZuSoQf0BmyNL++05NZm9laEXLH
4j+fyyA/Pdvp3Sq40AhAvmbbqtJRd0NdGMx78Mq5uNqCrH6FKUUXlGVduHN1jp3NzX7EZ+skY6YF
ZQRayUHf9jwakRi2ywEH8YENigDhOCR90zbgpvt1utOL5KV1iz1Gcm3JimhaHfsZYt4e9gpvLdNd
OPnUBk5z13wei7luG4DPfcbLvcWhrEf+soNcaVI1Cxwiaye2nnIyvVtcmMXmyL3OSIaEZ2bRk4HS
Th0J+29O6UHlmWVAeRTeoWBdbmnrjjKoB7eh9X/OESqGmo0POH2aEar+PtkQzrL/rVAbwAhnxX57
VrxSCYTgRhMQC+i8nvIEff/hv5HXS0L6BZsQEgaaVTC0OoV8SNoZK/3n3m/qJ5500Fckm9r8vS5D
6rUddMgI5Z3OlWeAZYhTQ4ufVKT1NTrGdDNjHzwKf51QpUUdpGM6yJnvRf1L5+4IrXF4h7jafP8Z
ClGAtNMNX1NgCZmTJXoqdhFCQVFeXm+Ex9cHl2wocIbVyIjkkvDGfz5DmIpN8n+ztdgfF3yJpj88
Sxlo7bBPuLAGZfeheKKvxmgpjZ+yRZAaqv7ZE/oINfWEr+uSSlLELDcrHn+cOZcCK4pV3ceqqIWb
Kf1duGkAxUat+xM5SF2hIvAtqzQmGSpJCZ6U0i2sgHDmjezg169gJiNyxryTMMTAIfajk1O4DqWm
k/Hq2cNn5lq8xlcRsvXGfLIGlUq297zNrQJx2oxqeS5bugLyrx7eoAR8LJHpd67Q+98GU3D5N0Nf
lNNo6PuTtgpGeIcw823xQ+mqw1PR4RGbM+RkAf/kCaD27ByRbLEZf2YOz2JT4x+btnYoCrCKMTLU
IHnXkcpmh8sOa0CmyT4cL4vMa39hWGx6PWKW1ieIxRjsKwJ+pRPkm7g6sEbXRddBABfTnEjjAGaA
ssWVoW/eIZFWmnk2BDVX2pmB4tUMUmNxh7+/qkAumBGqSjRFLxgJcZ1FnUISi0rNi2gLJUM+BCyW
XbpL2AUvQlJy7YSrxDNaSGQMwaLCJRFDls/hI1h52Js6sOkXaOIDMTHEosOqi6WBNPJs5Pcq7Avb
fA54bfZiOEl5jKRPyhUajxNf5Kh92uTRIDTnGjBy2o4o+99I/7sw/RTJW2HZbTbHPEi9fLmQJbSN
AEz1sydh8LPLY7kH46qzFGvJiE8f7+fof/GfDF3+BG3FtDmQ1BXNZUMTNl7xzxDV8OZvMtpJKCTa
xRzLL0v/YGKOPsQPwnlCzHHS/5+fL7nQzLxwcqmxxnfLVZPgk/XQqgQvfBE3McKHlCMhZfVeeTzU
jPfpXw9y1OpM/+d8EPqfAgndKwB5SLWoZDtButti9i4IMfbJZIRrdjWdiAKAxTB9P8izl1m42fVt
VUSH5TF2yBmUQFJZ7eeHdQlk7pB8/bZDGc8jV6JmK8ofNj/2jBt+3qZhxu+ul25NdQkqqGMXY9x7
9BsAa5vSLuM4Wi49fisno8U7nLch2y2WyeigvLjgLq3XsoiQ+FDsvWE0d/jH9qH8EcO2pVB2CsZf
j1g18tsoddaq01kS/irW9M9lzscAqPbAYR+lGX8LJNwURYvT/bgSp4QkYcP6+5xdYVSxvuQuybzW
lWNdc+4OAAR/T91pJ8VhMHsudkA3z0H5btIiQpB3a1GBI862YVFKxQtgiFrAFO0Oz0o5OeZWp44T
nIbuX+kuhZ0ABjdCylVAlHHqAx1bpHXJFZhGR4A2hqqalYQZh2L3BoPaSGiF8DVSE+n2YcAaUh1o
AboPy9W3Flh2UzyyzGAU5MMfJxlvtm018/Xwun3x1r2E8FHx8T2A1T623RP3xl+Jywq9x7yIHY6X
xJzpwze/ajz8kpL3nfHuwq17jQOmCWb9mRdYMVXnStk2Bz6LX315UXtSYknS+vXhoSCy1aeyw4dJ
WxvbkAEwIN43xFhCN8aUxGdnnKObkPhyEzMCW9jCeGlQ1OZ74+RfRt0AsWIoxMIjez2Y1zlmCef+
2UifzlRnNg3+dSEF0jeyQDNWTmxCmibR0c3FlfuAejROCfL9hLAwyyu1vkf7SRqIKZhsqVA9/ZvW
R/1mOoopDt7be/NJjKUT231zMBZpkvtPZ+n5gDqbURR+tCiPD7zdrs6QTXkXQEXyG9G5t88glrsy
a6ZVXh8m2AoGjzRttOlsDSg7Z7nShCpWUwweeiR6YsnflTDd5OjzWPkNUSD36H2CcMOd8GgeBp6j
GC+vuQ2ANt+sWjzgu17BT3+r6gP9ExmZrN3DNnNmF2KtP2IwRMtbHEKQuhsCZ+5F39d9SowRzkbJ
lG+Davs6Cbij4Wypra0jOfumT4PIalQqSMml6Fog8Qka+cGvZ3eIbQ0VvpLHSspvplb4e2twM4AP
IROqGwFWgx9wKlOw3UYZYE/5hgqgdXnq8qIwDCwd/L7DHnYaCf1xhEb8ztGkGNWfmOChFqy/Fauu
vnYCqORrVuY0DyYTcXw91NZTXTZOmo+30nE8rtvBDxPoyAWJZwl2907pFqmWAvsAtFxNZWfLVEHp
vxsCZQVmwBzb7ut/3ief335DAG3C//yzmi3e9hoWfheUJfbFVYPb1h+ZCFpnYtxL/PwDRtH+6qHb
F4TRoSNMrv6f5gKQwPwoNSBcoTsBtL3CvubJxTJ5KhLIoWf2Av5oyiUr2J4gFrbF6GdIYkrJI3PR
SipGUl8ylyUiCgJTNpL4yGrWfPIocQmAYBx9etJalf0KHunFLB6/hDqGijG3syRzT4Lsyoj6j/Vy
m3BEI16K1oM/IfHRUHCnUKl600tbG9TYvKkXR9BZsXIOnuyYsknA32brOQ0CJ3bSydXivLwuIu8J
driL6FAb0846/ZS7x0Bi7nFZpdS38KlLUCKKPxRqdk98tx0lF46TqAE7OWa7Gg8nnQVm/2U3FLLc
8SD8bj1yUc4DHA+1d8jb/qQVz9rdOpJW0BaBbmA9BDXuLuHy87/a8kEURhCkbA7yEs3fs782IRAq
V8nZLndNz8uwB0IzPHRAawuhfSZbGdMdgWH97E+ly2Q8N5332JD2jOwZBUxFItFuF7uRbY90LDWn
jBJItNBgSRpZSOyamNsSOrwNfnXFZyr/rD/cBtuG/hDik0fCAV2bDBxGFcn0XoYPvhMImiFNsEq4
66iZIdDgTDnkXNDkP7/VJp1SBHiFgHSDYDtu9zrYd2JfZiHDck2gHtlv7UiU6ZdoyhY3PDTW0pNS
9Of/75aLb8pI1DSnAQNrc9E1BNPzhGq/J5gzgFVB9D30CA6JfRKWRlablZVmPkXkZlWoEbANDGwF
rTSoMeSf1WUJsl11q/hh+NPTU6NCFkdDEwgk/JwoExCGilg5m0Q/ZoTcDipi/8USymFctMjXfYJF
2b4yMd5gj8ebKEXWduXrp0ztQr+6Tm9hD0fpbVA5Rten8YpbyFp9yClAoyeGhqzg04FFD1nKmegH
TRL4dZI1fIsVer08S1WTt6Cb7A0ihvaNQtdgUid4zVqiHGDJlQqTKbuTMEI4cK7cNZc9v/wK9Vkz
KGbL2z7v5owcG8OmPms+zOlldKyr5YTWGu23NLrYff56BNH8hVW3rnbuSgSHuN9337Top94HcOaL
5T1Gi4Nk3BJnQ6tyKOVKgM6DgUqwKcad5TCH9zTbSj6gAor7lqgIiHB0IWz9zZ8yBfJmSZqLHOpA
QQ2qHbfaekAcLDZsgxxnmreJCTkhzR14SENDqSaob30rfSa7s6qXfWuK0Af6iusssCkRaWH5+pmb
wTieG6HTAsXpWhjfg8VkMrLPuXsUhXQpTLlejHYdc7rpcRHOAdSjH4xF5chHzR5DuHeWa8dRIbSY
FatO6Hff/6/u7ffuxxzGLnPlLfwAC1y+l1DUAnTKVVjq4rrifV6PE8wiEFe43lq1mjLCQos9Tjy3
uOHp8v25+K6AmtNoeMC4TgguqGm7axOskwp2u/tKYm2jqvf0gPzxGCudTdyvvn9UolMZKJske0v2
QVjWhMbE0lkIBweCixLvRCpEZlNVXEuNN8Gl0NRlPMn/BUS9CzPwY3Pflxv61YWTeVlHs+T+HYYb
k2W44HnEPEheEg+jbm+v/SpUX2cPu3s6coWULmLJoY8jwH1c915jXi4N3p+QHAa2esOhEAesiJV9
VLL3hEO+OaQZrEkxhyG2BqkXG/b1isgrxBIoiSdaeceTHpxcXofxKesjANsvCqft0n8pkYN1HOX+
1jSCySfIz2s55xl+Kh8Ac3Sfer6OSkN7vJM73Qm5+JMYcUPHZAU+Jmhshvj9WQFT5WlOcYPFg05f
VOiRe5ZLb53/DWFnNxXQAr6CGo0mIYYG9Uyy69Ge8O/ModN9adPiZDoZCWebOW/Rg6snwtRdCHIX
PMxwPOUdcMIsBEG6Ve+lAMALhX4Y0DGKaLQseFa4mxIcFBjrlPaOazkFumM/md6yGV/3LvPQM8QE
9FDO4kFdAlukCDiK/9+K0hnRShn079V3Sem5nP+QPgq4KUTU/hpmgp50Cfr50EKE4nSiS88O5xnb
HsmOEIIwIbIuv7oojv65TYTUWLtvvlNHP/w5HpPM1Yd9/YN5c85rMizjY1KKdpA35afG8CAiSi4f
rJoHx+882azZPrdQPZ88m21e0sxd+Ii5WOH7u4lbLKacAo5lYoPYjQ2XrP4rs3SMxIvaLw9fy3OQ
AY3QIcllwpPP2KBLvmmDIfgg/jsOw2cgkQ8xhz5MKULlb+USWdgFRY4pOeWCLLYxwHTWTmmX8XzF
u3k4hrFl6eTi1LufuruKxycc0xB2C6F5qAS6t5XdFtLnm5d4nZD1zVLLxucujYWnavCnWxLAo4rj
/CFeI9ziToT1PyitBCdbc0nATX71p1qMI2s1Ags0eHzs9wBAgEspoLTZDYvonyurkLRTK3ePV2k6
u/ZjuExB68ferAmjDHRNfoE23VQxcpsQJ+onmd0qrIXoSGf9yaU/R4lSTwmZZZ1adZorzx04AQWt
N7m4YAdPe4rZVbvC9qnEIYn/mpw78rxZzeBlonGe4BatE4D9pVp9sFcvkrQ61prds+5zjzRWaKl6
h3S3Cwm/JZBDfwwo+K+whlCWoe6S9bGrUDh9qDDLzTNR8Ai+HLuOjMkDJHGH272rQxtJBNn2GhQ5
3B1I6TfxdZvpdY5AqIkLMx4X9wYAdApCFoUXbrNHMfkmbqrDd+ZLNFI8TYCg1nGsFRE+OElJJtv9
22hDJ7Vdofv5SvJ1GqM4Hg6lsKwDfYi42lSNvMKBwCAxD63VGBh56DBvd5g8Z8I1cuk79LqTrmdz
c81E5TFbPGz3lEDtcBgW8q9gT52v008z03365qwOrgY+4xeiM7QaZCXd+oR7D9aNqRHva7YV3xTW
MYaeqGaD1DZ5k8ULzt6+k2ZQ1BKY3SP3ahKc0DSt5amd0ZkG5k76W5oQqRxqyM6x66LjDJv89S3U
iHFDile0Z/9gYWQeZQyTxzir1XiJN8jZIQBNh9ln2AUFSZTxZpXTiMIrJ5eAfAsDUA0EssMVNLMa
bkbkT/dQ/MmYR1Hkk97EQrtjeuAx1PQci71tzUiN3pCao/725vL8eSjofvaRyGgBQdYhWXeSfW1l
22k4UUNP3q517VBaZTnVlugkHFX+ewq3rajoMyBSStDNl8ywpfZ0GZ98i5u1FIdfWU3MblVDZlMO
YeeVp6DxvE93A06BrGoY9RJL46IxBKEoE9IwECdSeXPA18KccowGH1+AmxEMHWBcftR8DJFoPvtI
MG3IQ09kqfsYIFufYy4ngkYH4LYyJISBizQAu+KNrAZAWHAFJd7jlo8FSJKbK/yTvH9DV+Jg+b9q
mkOex8rGPQ03HTJQhcjoN4sS9bILZpsVcJw0ymLKAOLRIP9Py39jOaMDkJrG9mfSJZIyENKNjtD9
XDMhv8cdr+xsAPKFcYyih1kf/es8uIWjaiDQep7UtSnFQLbjcnrUwPxuXwzFE6HbieV7tdpjhRqB
CQyFTrpjPIwkQNE4NpC6X1aLNQi3SyZRo/1vkRwU/6IkA/hANiYo9g+Qg7Lm2OsV3ZuGWzAsreQr
peSLYiypjbco5Ay1XrT8Ns8iSoaQQ6rel7q8ExfYAAolgvGn81voTULPK96ZCWOWCImPUa5rVrBh
CQSHkfPD6tXDWljyqw0XfgkAVPzKe48el9fZZnt8jj875FSUspX/K8GqNX2GWZF8X1IO0lxl1W/y
zl+eYQ3SVjaVa02r+a+CpvJSvR4Q5joB0JIIA0GK5z10KrjcudG+ppVwx5KimGlemC334YJciP3+
id068gUu11K0sCg4Rp82uI1vlYedcSQyFmIp94L2L1GoDoTUtSi4Uk3evga1c4SHawcpX/gEvtgD
6kJGFeSRhZIUgJ80c1ljKbIYj8IKTKwEXmW2ijwHf+Z8YN19IVB5ttBqWY/yogu1oLu52dJs05YT
NwRS25tkKg5vdJD0lODIUj2vN0pDM0dn3NJvTDA81gdc0tI7hUupZIarbja8xq0+BQ++IUFJqE/+
Yk+7fK8f382uJ1MsoFAE4Nmvt/nykRC/WiUV4d17EI2ra2R25+UKx6G9BlSCO+vdsD6btL2Gseu3
jOYmjr8buo5L8+CQ7PzfqxCgvlDZCw7ZUVn3ONmZiWQHeq8agNPtF1mJTCTc3LNF0SN2urli7ZJ5
o09b8F7wp3QiCxzUx/XGnnO/z3F6Lmh4sh5y2dhsTeqoFa/Z8vt/nyoW3lGp2/H4tPLA8oE//uqJ
A9UjyTl4/B18WTtqnj2X7QqfiFyCBeWVpZTkd7JwusGsnML2fr+tqGAGrqqhNGa61Nv3ncSoJ97Q
F3FEThxzFqWaakzlCiCpyQFc3qaP8HcNYKhrxQvXMkvQ0j38D6tW0XWQ8nb3VfEUr4UdUORUJp0h
K6L3mG4NyUakp4dCVEFg7tgm2rDTHRj+BjJ79du8HYbXaTR5e1dueIgwCtAiwSGj1RYortdREX4V
ZvJOuEC6uwvn6mViqvhQQ2yaFtHs3fxiroU+6QVLtPuSljWCPU99LzFlhy/cz2cy7MXCtGJ9lw+U
xYPj1ZCJZIiV1tw9ApPzyhLj44M/hd6xCKz4YQqCq6LL/wj+e0i94g5SWdaku7EmQRpLfjkbjtwz
chbGbCjriiklPU0qMxOHXhgq4O/c8OdFGbytUWMmY9MqPcSJeB7OaVAvzOga7+sv0DTP/FBnbO5R
bi4M2jbvz0sNjc2Y9D31T4d3CgW9sJxxVV28DpIXCaXFtHLwhN8BrwVAZOjovtYZSJ5gb/YhmhIk
Xz9IPWffv1RO/4YGujkjhkwLGTHXkmjDA56QORwWsKVY96PF84bRmQPehwF8Pv4SyhngL+MHpg5c
NE41iepoMMifDAMEeDJ2abmXh1tYLRQrWKfSPn5zA4mp6EkORdR59MqkgCD3oeVK7P/fWApiiiHc
IdNbl40kzRJsxymI9oeAcO+Mqf4p55yP/ZhPaBpRez9Xq2C19V8eyg9ZU34c5P3x02PS1dxzBgUv
0XJcawY1uF8wnp3sq1JyIiAPZMQaLzc4huGxWaIBlxDTXVzINoesNibQCG2HX5t6XMnuB6rTf62Y
CRQcmfzSi6KoZVEWHzgLxQEVOKVcclXcKoB+lCbls1WRryHlT2v0Hr3emn37cJ6Xlh4f23Gouj16
djjtdT1+Y5aQ2029kkTV0gKkNJo/lck4TSgeiwrMh4TtqI7c4pNFoMWo0wngxAvIgcchKx2rEBbA
JNIidtdftshSQJnJz7NGq1eIXyzG510PISl8dBSsP3aEYTqtmL/cu8QWi+5knL9PcW1t3CH+QcOx
vdMGUBQ4jvLndxRdiIuijdVGlZIHijCSbXywnX0v7zBisMe//cs1GNShTSNrabYfrUzR0pHoPtHZ
FRO2l0zgI1/gmLBrVVFhQBnlxTwgG+uTBEN06uUky2vQdKcCN6XOmvMIwntW18+9VASWm31KAEPs
qJ4V2m8aOb41K1kSYNjKvP+GTXtF7WMyW+kivMZeV++Muwl0suGKiG0iQjRghtUtVpiSVevyDsnC
P87fQHrbaPAE9VG++H6JavAT9J0pimZI1ImJhQpPJFIviiDt/IapexMp1ISAligmcM+Q+4vu4QFU
XzGeVsiLHbQ0vudG6sH4VNX4V0CJ77fHIp1tLU8e32Chnx8UcgPexB39ZcewymiEpDGgHTBdhcNo
8ug0/X+dxb4rEb76orMhu92Ctiiy2QLFz/zmrUuajoCTIRZOO59/yWTdS0LOSLjiqu0i3yeRX+bj
+pJxQZEDcLYXaJDqGFPoHVCFpHexlDD+r97VyUOTFPquzdmPpGPBPcrMTXOO1L5a4ndwD+JRyjDO
dviYR+6EzG8Tq4ASTSUYYSrPWJ9Zd8mztSW5Ah8zVOleWFwWNp/gM1XXWTUWwKP5g3P3noDadtDM
25MIfYow5l3HlgqTBaIycwbt7vG5MCzkruJFHzURc20UR0krLqVog7SMvgNyzjL1Ipd4fb2P5g1M
r/S4ElU8Jzbg254u5crVOdiqRFJfujdouUhXi+w3d4QL8RX1l5Rbo6QZsRknis2axRSP28qbauuy
y7tP8LsauUr9OqP+0f9XYoyyRJFY9V6i6YtLkq2LSULEs/VRTbRBnHS5uUPoE7k6+H3EcU6J03tF
7Oul5dXAtRsWjr7HU8gVdU/4R6GWkIu/QTkgFDlVq9w6Z3RCszHIYWJ3VLQ9Mhx3Ao0K8ON0NjJC
xVtVoWTlBol/cLij0VtnPH3lMuohA8km/mxmPaBV+MK9TP+33Rl313Gqv7SgnlK0p0l7xapvEW6O
ueMjIQQGNzDeipibkjMCJxO7sw++I27SJs9g7vBe0/PuzAS/4HhccWDQheCny2WOTqs4mtQ2eXrJ
1SoKgjbJyN6JqJcZIOJaicxGjrlXaWl+UbGwqfwSfwozNyJu3BHxibCynSFY3uYn7t52SUZVdpjV
6rTUvhDXzUg6IdTlHG90J9NugBQXMUNIMOMgL710IqbPIBX5AgAIm3X/TNfro6dm67LH/tdC5UX0
MxviwzASU8VNpH0AX8TEshIZ6ysg/NFuTDmAQqixXEvzhSx+r/erZ6TfUPqhAvgdANBclUQuhw1B
Lwv83OAUVS5NXz4LWTU5eyz+emYNIjmv/9/Cemqag3g2PLm/aKUiwduYompM8tpgq6iHbwKxBCRV
apCWrjkiUTDmfvNvmTiQl5a0OZcCrwfrkrZBHWrEhLAJIPZZwipI5xdxOZZJ/1G5W7RhRvrIcImT
Vbv6OX4t+rmuwc4yRMWuqdRGIwqssfGeFBmXTh9vPyyvLeCqvj4fOWVTdOCUFDmUKymXkrMZBu7v
dnCDouy7u9nWFkasmuVnCdGfdOBAxw0+mLY2sqQ9ItgNkH8mjS+4cdUbh6fiO+IIByBd2NiidXG+
Wa3T6TvDz3BTQWf4qR9aiHLtJHfB+KVdlS/6LtNLo6/w2lACYX/kdKXlacW6Z1E4LjarGESlUpjV
t6X/oCAmyInc8j04dDN81zTM4a1srDRxWyfKnBoMfrUeqNAS9YFtwUxzdgva85N234blZilHQpYK
r9DtVRDUMMSwrPJiMrb6Jw3BAjPtRB1KUNa7ogD+dmaIM0k01ye/nbbvulcE04oyreowj/C1CP/o
FiVVhkfvSbrS8KWh7LdI+EBUVd0Mq1iSyLcGA0H1NadN4RVVgzYemmpKnNx2NmwHOAeWctwVlpfz
mkB9B6waRdjKT9vgH5+1X1kvKDBi8s9UPsis7XBCQQE0kjXSrxtNJOsymtpIzd8coSTFIdnoCci+
H+jbLuLd+up6YxHRpFkhZeLjK5yXS9MJuKuO9SWh8tFr9UUjGIxZwFX3JUemcHzth+xDONVHDxAt
SjEPpTNP3wS18Ffvi1Ie4kePHaN11NCN8VbACBFvh2Rxx7DJmn6mdJpsoXhXTzXD16PylB4GuRCo
Q34IdBWMeam2/Cp0WoMkcy7j1Q90XZVJjnflSPqNhyheSde+phGmqfZCZtSh1rTO7Bgm9r6ywhmg
PIfpVZuFBYgsHDBaLmp09PFJss2PwgTiAfm59ELXXrLIdlV2CdFS0wIRCgNhFP7vxSneIJbV6X4m
ruPZP3b1p9a8avuapHVYcd99UYW61c3a+dUVILu+KGIOgxrc+DfDdf2NgnTV1qDBlg+idVXCUcsg
OzuGsrRwlwMsUXkwfy31sjLy6latMXCqXcfS6D9GSzE0Y3REtF9mXw1N7jru6ZgWLyO/S/LbfQcZ
glbaziMOwMSFgPage42tI+jV3UL4HgmHJ87OF/7ALAYSjrVVDet/EWcqY9AvC3/1fkhFW8/R8yFC
jWPKWD+xIHHnaV5Tl3D6ei/7xQR0S3QBw8LnvkleW9Iy+0mFNg52cfDMFfVx2Ak4xyfIdA8txR+M
/bXBU2HEKPHAimS0Lk3PVT4m/ccktAZumC4VtR7637skKtHeyaG6AicpWkU5gDbb6FR4J3naEsbC
RsI1ixDfKCmqgpcOp+ZVtLdDM2mzORLZu126dkuL5G2TYpjpY95YrQZvivSOg2XNIxHrY+0x0wAC
GZQECnF2rDD9JuGE1Jvo8JOaP6yHtwbHuiYep4XBfS3WMiISI9eSclISClMPTXMq90BXc6UUGoBs
sk9Y2XGMjHt2f7Nj+Q73pNnaCZMiFVnVk6TI+MTUbWvYPc5vmdTD/gRrnCkTRp46JJiSLHAcgHMb
GDq7Ig0yyQ0k/z9DAlmZ/gsWcvljRsGrJROhhINsG2xFFZNipqoaGaXatgmp69DBpVqTWdnlTHk4
9KAjPQlpimu0tdJCWXdTrdcMtVUJnSJ3jCWOg1PA4qvtHlDIq73GpWti8LjNNa6kaLIbfpPbQOJO
8tdCgQmQOhTIi8GKF2dD3HoXk1vd7Dj+QJSsJoRAtBYmfKMUoRFomOejFh/NyyaoOxH2SinxOP19
8zyWEkSg+Ax7IvzwVVjU8HA4t8KxsFptAhYElbQXPS9cDSKsQOeyTyAqUloY2KFhpEeZigntQ20r
+hogbEeGxWZYwlqYCIEHvi9ZHkqVRxPSN6e6kqy4h4oKLhtVlgMhC9TebkUQ0tBNDTjBj9qmX6qX
ZJ2HIIlWLF45O5w9OH8O759IAhxypdTGhzueWsTTax6EhNW9psu6pkLt+ZYLwWBC53x/Y7gMq+bM
u0NFkm8VzaRLytLJ1m67pbe9sFDAgxEfoI3PSooGiaQsrVAZ725VDg9nY1uUV5eFWuTM2B3raVFp
nTjEg3/qSaKmWBHzjW35MPbhKoHWfR8D0tXmoJBw5TlojR8MbbGD5D9MKUarotub9evRObz04UY2
PACu91Rim5ex0BiRK/jHS7qIFvEW/uQ7J7FKq5JR05E4ZSIOwUFuRQMnt56vV3h5hnSYy32WWL13
D7ExdAVcJAuVjPRTwDyXSkSp5x0uGg9NB2iu/y4s9hsC47ahYmjb9FeVsh12MWgwxx9HAmsCqfXw
UxNjMBdKf1ogZ9gpt/TmPpelGxh+F4aUskci8pxjaU1ZpBsn0D1/AxZMPHGwJUYSm3UsP35DGx4j
TGnaLix7TxWSaqt38eA3xzmjarGjxgH+PlaHzLMhgOVFL4BP47EAqgjVqXJFSm6shdY4nkRV9IX1
3ZKzB8FRbw/WKAkQct5Piy6bAIJ300Mv8keUuUuPQx9dJZSoyML8GWcPKrYtOiFipJLhyY6WFNnM
vkD9T5iQ1cUHJJKxx7YUX2HqO9vbwRmB8OW1BPeXsrGsNE4JVk9neiYNGZ/1odSgy9EzR0/qWA3C
ZNfy2gPw/hMIx3tWjPx2D5AJ4sSpWwwQ1J7PsMmDHc6vAtc7ibtPtPAUrHBEoUR4BoRPvzcqAKdz
Dqbtti3Ud5rmGOy4kwyvJ9ME6Oh0pgC3nlZLPmxwdonpX1hj7XNxoVM6sD2qH1aFlGqse0wEpUOP
zQf9Z6SXQuQBQV7sH1NLxb11eH5ny6POWCKWaFkAMefEuqgPARFBO12nTVa/4vHMohNuEabVnrzb
x1jK8F6Su/SuG5m1yEC9GpONxKgzW8uigdL7HWvU9CwkhJFEQdJrBCBmA2tF+vn57c8HtsSSXVzz
0Yesv+YDENJ3KZrkDMwJS/Y/gwnMsSjeSq6buAEUKpo90TC3udTQSk1f7qnUCw1iIVzm7GevUD83
9ZmiwCydczgYyWvXOxrZ4TkIgVav1RvHVk3PRgZ+N0QgCIJFLGN6l5bMvQQljqE11d36aAnwmm1x
WOuARCdc/ntUdHXxuGS5+i4ZQp6QR37GzWaV+OTGO6LqhV4chOviGmb9UifyikPlNLhyUKcU9zV8
jp5v7idIYjUuTbsU+TtI4RyBt8KYbttz2AmOqsGk2IDJAUvm8X4ESS0aTIgyYiyU+DubcWa+tBmD
lSuX87r9ZvMFaydW3J+G4CanWmgPtrBrwaVUmtqHvoLige++lHwUox5DqRkoDnd8F/NTFrsAqGfO
87oKkm7IVFa+h1xKEiyIwq/NvvhSbYSXSmReO4u1tO1C8brI/J6aPWqsSRQo+yT1eooxN5w0N3Yq
YxyOq0NZCdU75RZAzE2Px11QSJsvsxCWEMU7aD0EVaAn/6T+nrS7aKPVubJgud0j3mNjzxgBID+P
eY1kF/WM89+H/DuDL5154HbLcSKKWqjEPfKjLUo+XFa4WpZLhWsrUO5yu/nxxrryGGhvGTLP+YLy
afRBK63NvrvfLsLGAZWDzicKNK6cYXFQJjMQTyOOPbBB6vvQqwUmYFnm7cInIWjmCaqe0sOUEpoB
fHWc7UEc5aC+icO+a9XZJCqdzy6ZhQNFh6D3KrduZO43i3d3g36+xTyQxflRKa2IfxDeVl2/B0mk
eZSqLXJvaVysjIKHNquN3ZrNIv4iLf3RBuG+Y4b0BIAJfpJvhpN7D5JiEF1+81gpQvV16bzle6mq
PoTS30ge4+YSFERST63Us1asokds6KAvt660LdnGuqoUZKuXfb/toEWzm10Owqyp1Uj0Tq4DXJ11
N4HyIxayyTZPE0phgG1mjvMmFDrGU2+5yA4qiRYig8hzF5btM3WRPOh+5RTg4+clU1knDeOYpET3
WlLay882CUvfoJWddod4dT0zKRLBllQhx5JmIeZyIkdKbSCWEavFJkvOimadcrzgaI5NtMk1o4b3
ZUxcUf0ovDIMhzqN6DJpgd9tkYaY9ZQQLLRsQz2tkeKKilUGqAHmlCZgz8WEnskA1K0RU1BHLulD
gMPZxhP6XwHDULlCbd8sST2oYdoq256YBZgLDnWQ+6gBeX2Quo637lyWk7yAK/gOdW0x2T9UNXU0
PqdGFjkghysmdJKg+3rKt0GrK/QexaWnYUDZAwi6FfEK30gPvexFBMq2sHREjbb/RjD8LClhL3rj
4LCdfJBSw5jEd6gah9ZayPB6orXKzozFOKgx8oAQnIx4lZiEZK9N7K0JMVoJhgZ2ap4gF3K8+ho1
oLGVCuK+AWa676ymeug4sf6EpgHGaURKYoE/+koK53UtMnYNLea8w+ZgeCifscp2FkYfxZ5uPX1l
auHTiTQZwER9+0v59D1Lmg8i3ijNUYTLrBvY+Si5LRqAkl9jK+RtRor1/RZcHQPDadE+v3zwWE3H
RkNA7XF+GsI4Uo4Co/VnfXq0BJy8xizyD+UBAnuqBGELx2FAOnBnRCMra1xpbhv/VR/tqJ2fcRlz
IxaTjkc78iks7ZyhSvhW/Jf33waUeslryrhuUfrvnMh0HgG9TuIpml4eLbBXnoETOtt79Bv2sq4V
9Pu3Ol27Tyg7xDyCtvucWxpwogC2JkyxjlGZemwZd7A+px8/FObDbeRsCSfas90xqQeWThiW2qe5
xItN6hueB1ZzTScYj6YcmAlkJ63VjYBkPf+FybWzJ2ZxQccrjovWqygNW+R+gzXfluSljnYBYWI4
tsrRkFIgMYkczFSydqdf/I3IkSdmHGGQM7ngKsSlekyTaMCod1ggZoOZ3NnXFRCmwlcDdfGLoYyC
McWvusCSlhUfR5qrUtgSvgW/T8Mw62Y0H6t8AFDfOkGyQKadBeia/xlKPpbOJvByeAVOonf7v2t6
MeoxULB3x0tJO/mb+e3huxFQUtToF61ViWScmg+re0gjtRHxNoIswWRy3+tbvtr8cQghgKnDSXF1
HgvEDdEk6hebEuH3AH9t7XhYBqlO4hgeNvqgSoU9at0vfIRokDxfMkVf4VUAvJr+aMaxtjYr0l3c
hcLqzwYXkocC+3ZJB8bDZOZhLbXcKbYttWTE4UcqSXOT3AG0dK1h7cIEaSNbaswIPdKlRqwUtM7X
2YjyVdNtOfnHX/JIGSfOYwlVcN1I2lHtAuvhw2l3jZy2tEHtjA/rp/w2Sxl0nTK3c2pPy1aPAPs0
EfTBGv6T1FBcbxaw2gBNGj/bRNtd5YIwlqKWh8JJEcWdYzP77xRq5AbWNnILb9eXji/OyAaSPcW2
5fPq29w5m4wNleJlfqtbNjKt3ZM+rujhLULwcFNZGvxFHYp8nmvAu2MiyiL3MAD8t6R2LCy4ipP9
IFMZt+IBBPogdOH1NbNGj9QtPHB2RrzUD5x3RQV/yKm6f1UQRbfkV4cK4ptMSoP7o4PcRM1gcY0V
s5DJDgntDOpKvsbss0rCDd+eDnHhYiTNcBWtGG0mj32BCCMx3oZ5hOCVSXBHbOmGtd8fHGKO1gWO
vG8/z8uUetoLEYk0XbgOLEmfmWdZ6TOAgXa3A4TJG9ZWDefmY/1EmKHqBXozoqlnGkoYZ1q6F8qH
ev0/z1qqLIhbkJNQeum8gd99oRcnQzLE2cywGO4vXproscUfSFcyP7VE17caIJZWv40VbO2GVn0Q
0I5QfaeFyU5NeMAcoelRdzd9l6NJRZT9crj/O15mvnGr5QbHOhntgEnk7qt7NzC8v9Sid7E/4Q8Y
Rhje2xnAPdAK1WSV0vIT3I0D7iIZJn8XHy+id64Wnl97RYKMIIMWAnKnK2mvtJY3Hg++X1H2Mljk
FvdYHAN2EuuRt19J5gHwAnIeyA4hv8c5QsoPCWad2QBl72U2VCwRcdfoWaO26elmwMhjygkFYZHf
r7PFbLkoEaamcomCjLuUaOGB6TOzLARgOCcX81pQvE4+2VmnjHaqqr5NlY4UvFJ4D3qZiLifGKbZ
Xi1MnActbp03WizOFS+VesuI3GO2quEOnk2xrmmRtvwg9S+4yy35mJNArVVuZse1cuoqZkiPmqDa
W5SB3F2Sm86dGMy8FcC4WQoq4I4pgnvcHtqJCROZ4/4TvuiDtrXG85ealjnaREac98WfQCIJYh87
U7AsTDM7xy7exzgMctvBVaRgpXrCs7zl9W/5rZuX1q/VHUE7b4aYFujv95NyNlcxY/XaBYukcK7k
afp8kttd7mUJzjnjm+m+seziy/Yf287OYghOgzmF9o100DqTjyVUHILkIkgJKpszx9YP0bbjIzXE
VhlhuUCW0M8mB4uRQmRfI+1P4QNw2I+tmAxIKhfbcVGZVnO6lLdQsMsa+SO7i2fTx6wKOixZ6WGe
ZIfzTZITkUEKtvB6s+JGrb8dkhMQ3ngAf4w700QtDsT20lz+AHouP4BG0h/NhpZwDcYUO0AX4zKC
Wn3JL8onRTpJ18fNCWWCRh3WNmvfPL/VqXOA33VywwAiT3aiOksmbA2vWKuWuewFf0M85XK2dEq2
Vep9Xi+7f/WVgCgx9vV/zkWZUJAjcEp5F8vfBiQdqqtJZ2lGyu030m5UPbdzuN6IIuSqYfBNgXXN
x0Awag8+ceYuREl0DuAvNTvad4RggtGLwO9h3npu15eA/To7vh1TFHBzDh//H4qTbN0nukPm2lDs
k9Zu4u7usxuqwfz2p0LX17GiHSQGT1Q2cW4AorMQ1ga8HEv+BkEaFjBEaZAPTtCpMokPm605k6ng
aR+shZsDHAWsx/x/TpDN0IAtLy5bnJr6wLtQQDgO/cVTH2GjjfMtYuTbjsl1ezoOLKCyv3Qhw1PA
6LphqQsf5BSw9FZ23fYHmvTPUzzh9TKVcvPAqdrDKy28KE71AkQCnTcQD1782HYC9BfbdfLKU8vz
NrxGbHouhjVgHPiUtRtg4MJAFUn0eoql6CVjxt88QcGh0Ii+hHe6v+taoKE1V55V8DIehIOX6AEV
Bqeaiu7FYJBB5vwG2CtU4f7qmW+Tbu/BRqbc9IMZeYm6cnBY5dkz3wXaz1lemm58/6ABLc55uqDK
AqXe7uqCkfFAWJFCbfuQOYextQfCacjMq67ZeLgoaAoJ1wxtd5Kli7cLXyZ8Ee8bt06/+OpEiUrV
ZAhxbbXvsbrmuvKEl4fEjlvSh5MhINcNzJVZIsTIULBF+Zaf6351/OYkBpRA6QlJfH4+PS14umaP
DOZQ+L41QHX/f4IBuuK0PLAXUcE7Xzfm0R3STqsiOF3wpEgsxSnS8l776ZNmjBD9eMaAcoooHUaS
gjOaFW5QNkxQZEwR5otp8PSuHcBbIECSZ6X2R6mQhI60CY0LXCfMBWevZ6o6KGMRRAT01ZqotnDQ
mqlnF4wX07r6pGf1Db8n2cR6M2pxLg3bjxObdNO0z6Np934rBRxd0EJt5+aWNNzj4DVr0C2GflWe
PhS6O3i5LNXjvZKtdr5imc5abQsj71BX9gMXrRt7Gdv7UWSGy2j7D2teS/yXxk0BcKB2k+nFykFp
shsKecyF9Hp0+e7NHSTTHCDZXf51xRVKz2o95IxA4kRkzYF+2+b2UoR8iYY8Q+IGFFbpYXtBtKaU
ympUlbNzZT1ANsWLjlH0O7UwIjL8n2ZB92U9CvaTZ6nxKx3zvaFYRDrBOKDSxImlRgg6yk3/e3TU
4X1WHa2mO6new9+uRO8/dmOIdIZW3ZA0mN05OoYRJCaRUHy8G3sJxdSA3cshomYsjbiyz3Mdr6CG
joYzirx3Xb0mBUr3H+kK98jmkahmeeckUM+BDaNKntFR9a1D3qtbWFb3ByINokq/M9W+UVyH2Vdi
YuubabzmSiPxhIMv0/uRMDrU/cULCsx6+5yePZyham95l8SqPKoGFTIXO+d29PTj/CuHGWHV2YhR
3IEihIOO5jNSRJWaRb0ZHmpmOSo9atYIWwKUBCZ5mdCzA6FLy12PzPw781n+RFK4pEe5crlX0u5k
2M13uZXJnODLwvFa1yZoqHItYwGdjvw0MU0UmTdu8gGllsfDZ83Srls3fbP7gsqW3Y7H36Dw8OAH
kBWy1CfJV8ViI/VfmTuK+jD/l2hPAwaFGsyfk2h7z6nDGz076ymM96gtkDRdYlAST0UGE/4hFHMw
p9yGnBxgKwmfypEtK4dTxVoDmpgTfMH/ZzljKYUNzl+lQqWLRZxk44hUUEk6ST7PVk8SuGj+9p4D
OnPDn84ws9eVVxC2Gbkg2DO0JXDexg6ggsaYQUb1ZjshxCRf7JyDYRv+Cq9bYf/ciXJ09Ay8GMig
lRdIFONRWWnanZ9OFlqQ7qoxjZPEt44e4TZUKHzguAfEYp905BJ/QiWht8KVzI/mzhBVT+dA9Ook
xmJNYmgXX3xp2rOJSuggz9+wwD5jguQ6/ug0xOs1bo3kz2rSQOAo2DCxU8dfyQPwEbW2PJBPYF1k
sOu7nvFmJ6gRzWcwfd5iBy5kBJ0Q/Pd4CClVSuyz7NKGZpX1Sao1YXfd0TVjkfttn14URzfILWhd
e4Qv9gg8fxMG2tyDXf0NXwRx+I97xdkmEdHbd5o6nLrYKasDvtdJv/sFgP1GdzwY/9ssdvRhpN5m
JvTo0wAuNWi7EU7/qm0V7lOvQDYlMk31VhvnQM0ECCGKU4ZESAOy6xeAZiivLbfPKX6K9Pi88icQ
bIBmzpC4xdBfLqJXgFmgxLSHYDjMlj0igcJKIzM7VaDY5tMsJ8LR8kTxZtpgEefEfh5Rxv/NSQOO
/Dz4sDdV+rHhB5TAlL6dcPvA00LnjeaAyxjP4omWHaP5Lb//zaTnwjo4HiJGkuc0lw8YPFzy6eQi
rNsiZNPYi4KbckBNm2Zx9EPu/9eE2O/7NmVlEnUeSSzNhq26c08jlOkd3Of7QZH3sQTsXuYeMpc/
EcrY2taswoV1kfy5XixB8J32sN70c0OHjwN8ziQ64C5tzJJnpQ+5S7nHisgr4GAUN8XK2STt5MZs
bDXYCkxAt/sPXqJ1NRc4x/lbFghDe+iZz4y3A70FXkIuwj2XziQra9+QRyoXPVb7oGqcjGEE2bNO
JPcInnc76yiUt87uYnGuYMBN3vyU5SbQOqgN/ldcW64fHYKSqzWGUXzPLiAof0J6YqdBjPFb6PG/
bOgliPtHFbieNWYBXg19PM7SOBC0lnkyXiKd8Ctlqhz+VKuRo/AeSuAjQ4PiisPsBBvwbo27ygCw
GJyzPSSFe5GCIJj6jX43fL+aJtHRl/0mh0GWqRZuF4zIKoRqvaIl9JzJLP8CjbRJuTQUBJgPBgTO
3U4PFmuDOITxpPVh91ZWZI2IJgLBh6GhExRSWmZAy7Ixjktn11hIGp7OPou0eK1jDSjkj6z2pz7Y
7jHehy55qes7HCek190V5lChct8DBTM1YP5VVhyeAgaTZPJbQBBU2bnA95eVk0VbQq8kVFWPpN/o
e3pt9OhNig1qIIAF5z7MR0GOsgYTEHVlW9dUS+GKXEVvHxthmYNahXqy8V6q00UhPANGcCBcz2y4
N+HHmNzsXT8bNETgWwA20uvGpd6JjTsQXjVgVUlYYymRB1OyAX7OTkNcUaxjzEn7mg6jqhtfgZ4f
9NuIvHnb550+xhV0XjGzs24Rt26bLOSm9xav64Ws+9zUjQFuQ1ldTrABkFbPgNjUjiDIbfHiIsWp
6XtdTHtTO1wFzMYtNa6Wk/vavXbhF8ZwGr+ltc4YfnJo4G8RU7QqqgSkLhKRduOrpqFffzEgJHFR
G+jH6qGpZ8XjUf4Pn35Ckr0UMtvueGZESqsYZzKUINnJmUdNfNvExzemwtyTL5nYLtG+BUIBt7Ul
DHbPRMgtsBe+g8QNDVfqsmlPbeixRSK7CN2fwGMs+BF1ZTV7m1VhKZpy8j4ve4TqN5+hPxK/Zv7I
gqU6IyaCRsEfeS3rK9eti27l9t0uatB9GqowuCuA7+wGShzRgsHkp8BdjmBpsPYYNrjWuHKJOFO7
IdHCcXWlPqC9CprbuUXMRxes/HxSPdchjdCcOAmRM9NOJKPok/Yqe5a6h9Ryl7zJR/8oxTpbovE7
q2jvx/VDBMreeeKyayJh2qEV8BmjP+G+PyUujcCWfcOkdcD9+4C8eHBXosVBL80iptMXgJq3eHTo
9CvZPS3mRRKZEIBZLpS+hJTRCWfd7Q3tf8FZfbVBShLIF5xDtZzkSIJUHq9CCcB+Pa4dzKC7pXUQ
FpCbpw9mRBy9yaVOtlDZ9SOX/YAmNxjlVI9X8mL9MO1w5KCE95tLW/xe/MlwUEPWdZk+O831fu4s
JTnaP9QfcvVuYEHvhDawo/Wjc9nEgSdHvdZo5H4lcEG3VPk9zdYVZhErqhB1CHV+HVA9zTz9fKdH
i7RJ3rPjmcYtBEtXV+FI3BVds2yW/+qo2qopuPlzp/3fzEqrG2vyyYD9HJKm0cOMECvLfLiJzdcu
f3NzbSPXeYd8AWcqs2WBv5g3Rh9OC+geZ5na0YG9OMTGV9fBGPh0Ibrv/BJEobh4iiZzYlsi8F9y
khw22LwpPvnFHAmGJKyLFY4Uf3/bUrRJtETccyBdawx+IECIlx8KE5d6E4dTdxxwVVNhx8i0/M2S
13ImqBwkUmTVQHGNRMvlvPfRsIVN0SWNWha5Eo4ST22Mcdn2SeCkfO5Xtb1yQ4OZxAjclj1JUOKU
t8rYmajlgOjcHG674oxWpq8bSZYSqUlrEjgMrmz0VuBRMaSCjVnok07zejtAqm67NwK8Ub6XP5Lg
TcMnr1VkIt/CFEQf0+kgEfVyhMhLnX8fo61NVM5lYUggkBEP8ONYuyrSOk/7aD0uaSq+Ru6erYEX
R6xaUhqSSq2cZpkChAku5DBCgoua9yEkTdyQovWjQ7Gx0CUKGATMsE//XONZwPAwyj6o7bdrh6P+
uBLFUoZsEyv1rkG7M921UsRB4PV+SxS1u72qZuTQXebohtPr6zJqJcI8hN00K0XmXn43xXl/fEI7
vrUCBV0EMEI65KcI0sJ9GNI0fqLzAPfhbhJvTyIl1edjaHEYX28Fc0jEjGANyTko9fVs9NbRQBEq
unaurVdheTGuH6xamm5vCmSVBch8EWilO/7JWRWRKXYUb6urHlrH7ftWn/0LMRqiC+dxNN1HZGwF
MPfGGkMY6QYYg9s1GL7tW22wsLnArqLh+/jUBxINWH1hh1FEhpNrOyGfWG47Y5mWY0uDeRgvTeQm
3VSsfJmNJt9mIxfd9YBfVr+eBjNTeas8RHb9Lzsjhvj+RNc5D6xs9arCp4bEOCiaDrW22S2LDP8V
OI6QLB4uP0ddSK9sxkK/LCilcy0w+w6hGD8xyVGbtaZTdFAjOcAczhDNOxrnwphu5ryGyxUB7t7Q
51jRbSXgMv5AZFUxHXeNqnCL6c4qw1RkIdFXyVQlZsrLvFro18rufb5sC4gNQ3pGoXUsAYQOz03r
0YPWX/OJmBRoQdM6PtOut+SI3CY3RTPTpVFEwbVj9lmmrShrSjwaUn1g1zsAyeBOwdsg/OlGSpqb
xhaq4G5YEfIMRumFePW4Uk7LQ/5kZnw4I8g1heDr6Y1DBFmeX8JFODI3Jov0e80+4K2ShDZiJ0fN
ClAjQ8XVbS9z/tviYGmlwLHCWPZis06HzoKrmB0LFp+if9FYUrZ5NnT+DlIhmEKxxXItMri5Yccs
sLJUhZS0ZConyD96NDdP3s6YqSu5zHgIiyvTuGsoVkidZd42Vwj6rLqRmCcUUTZTr+sj0ZY/HNm6
IcZoOKWRWUE83YHHjZmmUMiRaCeFMLZPL0zffglOjKyrYwf7RLhQQv8DXF9tLT9/Q2nFHOf5HtWg
5bgBDyimcf0zTsVIzjIzm65YPLHThPnp+bUSihNWliBAlgJC2GR4PK99Lcm6yggYC27yqIyXVAof
gtD5G6toyP+QzpZ9wpRDfcsRMlaw6UVEoOxN441f/surP4J8CU75nwQfVp9UuvbXHr8fxH9ZOXiu
eIPrfTuLwZwmj4nzY7qC1eyCbKRnYuqaIpBHvb1/INRDel9KaCiCsZkaOFOx71MWY7+Vw9yGSx/n
GpQ52k+Zb4JOoYwDlRCq6Vy9tvsHOIO0zX1jTVsU2+6yDjg091kpLvf6OrMuuHpNtu2zzTrty8Yt
B7nrgGGR3+6EjkCRziuXewDpxAfaevbbdY3ZatwUgb4lJIMf3fqxItAGj+klbOilz7mAdLKLw/sN
BNrT7rzNfBxeaR2QbbKR/JYOqFr3ePJMky7UaiL9XkyEfIQoYq+TRfZ0+XRWDFsOg5PiHXTzAlAC
J2Geos/0dRad3iNVPh5tVHLW6Y4WwiogFw8B8zzA5/Di8nkKM/m4R8CKZkZRy49FJtvMIxMsp6Bc
EWmJdx/D5cQd9ZVSZJtA2/qOkTXVqZMoDGxtBZsCHI/DjfJ5//n7NWQg3Jlx7uPEinEpECReRDlv
/Ya1HgVp5ePQVw4dOR6ZGR6ECd294qfg1lySPKT1qJRWzahkP8cNgKKOepaFpT4iLwpM3IyCr93c
TcwLyw72ZAI0Uck9vUASxhuo9eGzf964GT2tk5EhLEjtnTgpi+670T61Mq+bLflJaXkQoGvwBIUn
2j1UE8iVdp+YjxoIlugf6DgeCWriowYoJOWefdZA/PoKULe8mf5CJlqzEJquhuvBS+DVqy+PyEdL
tiqh3t/TNNnve8IGp1FSeLDrE9Zh1ZOWtEuhTZIECkuqXhSKzXKKBPbvF7xHNa0ITgKLuiSdZ6V+
O/5bGSgZlY5pd5AqTdki6Pz9u7YxAxVbfZmij643XjD94iCTCgbYgm9CSvUJUV0J8m3lubrutDj0
asxYHiGx4CWZBNUOyQjEZMJ8TeWOAJNBfBnOMLB+qzLpoJeLDqqeVxWL0xQjLCWwunFFpJoGCgvY
nUbChWvIesWIwPaITd4JOV1B7VQECAls6qPZQ7DfcLNydBVrdP6lfRyLOJtJQE/zakU60nH+MFgH
UwWiig3aXxv3pHjUFCgKMdfowtYRAwFunifOVwfvX/73MhTYK1EnBjNDbUb4dAbXIoiaMauBBf/L
jNhvirk64LEY1xNPrY0v2gT4ldUL5csM4rKPQ8D6TtMKTxtBJ66TV/h8H2eyP36UOYGcQbdChO0L
8fmbMa8W0xgoTl4QKcn4rAWV6vkdBgyQLo3Qw0hfyhOHx66gA8CwnvBxhc0O6Ylb5L9I22mvOFul
lj6L1obebL8uVoGMfX0/eqWccTs9rGYkUU54tl33oT1IuxLrWE+oA2SENISrjrcYqBLSWj2Zc7nl
9j4zQksCsBOW2RxdhjiQV0jEGn3XxS2D5oGqKElS2CgGruukaozGqRY5XC7v6LvbaPm4QMaZdy51
35SxG9NSLqN7uGaimnNeoW0zMQF+oG0H9gKY1lTIlQhoqzynhKtKyV3J1yDUEQOd0fwI1u68xEAX
nOlhGCnrPA64qSGzNLCVFwpI++YOqeArRO0k7r83/kp20CeLRoeURpynU4ET1ZE2ntaKXOLq8Ua7
j+/sJbp6+G2zTyIiTBpsWuVXAwe/xcTWQYGb0YrFhgBHgzoEZyK/epi6TYydDNWn/omVo9vVke2y
NMeoglqeGR2dQmxikq+uj5GqU9pF+PbnQusG1Fs9DCg93B7TbA2WISGe6GyznAGOD2dEEKWYgxFD
ZlYwISzDSN3naBdWZPxS39CN8wjBwVIdrIEYizFPxpJqVJbzjEuqQ3HbGOBffDaVjyg34FCaI981
M0lgvqFX8Yiw6aAcffRRQfOulnrNBfROG5EC/w1/3yYDNnHgL6xrnvg7ggpK26MZbWhDfPiuRv90
3+5Sfzc93ZXyjFPKj/+Rp1ns4ruNDZLv/HtRDP8i2CxH3swElyEsyNzwF0eMGnhh0QpLLT3oKQUv
yeL5yv5Ga00rbxIfa63lrHF28ZQ0A2Qa8LWI4afV6+bta2uCPjkkX7P701CCm27pE31Zz94hHFoZ
Fc1rB/ySuOIfqIZEaUmvIFw/hqK7qyDOhwVMON8EuprUnC5tIKnIoDcvmeJr0pDqWBH4vBYboruH
oUXnexy+G1rDi8BvW/n6xEqGmozLnthCRwdMtEQAgsaDdlrUOH6AfCK0NdoWngM7RRn7ZYoxdo15
a6cAaTXcfe/eFOfjcbCEn4yKZX8aygh4DF0Wx0C2rIwF6iWmiJHktzQ2dWWp5GV+PgtIu+ahrw4O
4xE8Om4f374QuzDL8q0R97VxFrNdszZni1FNKZd3WhOCtIYdh4TQTo9aN1b/KCPjADL0MB+qQyYm
70U/X9YD7Jt87KlKbr2HkQ89ePPhRBB6FJTSoaBsWjG8x2BSzWvuqjUgzoJED/uplIUcVYNPt7rH
+k/QEu8ClB3byAyT9Je2LZviK6liztXVAJ/7ztjiK01Edp173iNztzztuTF25rvtOyDOEytiYtOO
AajVQEJjobV1VHzW73OEIkeJQuGObzvuhubh6vTlg42WPxz2W9x89fhn1l2eXYFoywEapL5z+cJU
Khj46AlAWYLy/OpoJeWHAargwdbJ3QOLtq+rCw43OcpFeQG9IhsJ3E/4iqmVgGVjZXGF+Rug4kTY
EIupf3hERYd/rUJ5Lcgfw7Y5/IcnAqiYodQZo4g4TClOs7IJeXgNBDg7HoXX3IODXje7kYXFdEqX
XLLQy0Asmo+mUoKClCWOwE5TFkSdg+xD90URwMDT3CPOScoMbLt0T0XwyCmf9TdZecbyJsJjVIXl
oZBVsxiaeaDZRio/f3jVq6kMnPnmUfylosLEpbdjpZx/BtXPDkwf9Ly4kezYxpMP2bKUZ4prfym1
sdBCGXmWP6HhbSzv7HFPRVjFxc6IqTQ76sm0IE3GxYgDxIAbgbfdqBbJGCmYZDpCPPu+OnxK1hWH
M4iUM66u97T8ku8TQRHxLnuZhZJaF9ujKMEn7/oDrCoQXhqEwxggU8AKuEzQilG+IS+WL6fbptF/
JawBZ8ipWcaUVeuwk7SiHIumoMWCo2MmVTDlQmFXF5iXNVfmn6v0RlYqF/NrXZ5SucrEzi1FDsVH
pyZKQB8ZLn4ZJpEWL+7X/VkhzV1sndrTz4V7K8bBMzCyKnQLz0lOL5Yp3bEDvHlGxp6YxDNY2a6e
hmJCXPZxQJq+18U95FZSng+R7Zb0N7NxjB3HFthZmQlN5xrJbp6hoUQmX8Os3gtzmGi4HrMbaVd1
A6qSpu7D8fvC/loM8xtVHrLp9j8B1YZL6pDLm62VzxIdVcbn9WxthjgW3H+llCVjZ2Y8mrKk2zby
B+3iCWIhDM9u++iHdsgqWXCrA6L3/ygr00JidBrzuSCAdTedEL6TKxgHUxYbKhTOEpDj+qvaeoxu
u8JytcDesyeZ1mrVYnDRG3jHoyFB83Dq+szYniQYL4ytby10w4EQcC0IQB469mzmIFowv0ksEwLq
dEsbSRfNpZJfrvydij3UCxGvjHAhbrLpcqQF7HEykHTk6izABYvd090vMWruz3PH6LwufZKD53F5
JXxYro6Yx1wWPLjSlmfIJs7jrDIHeUVw75nm28pCrkDD/dc2YXZ44+jikfScWD/VnHyEEO7VQqYk
0FFrR8slCWOzCiCKaKdFvsDfJC235rWoHQl28JeFTS/mOb1w2ls37sh8K9M/7Byuy5xdTP9NKgBA
2QXlvpAHbsXHUvjLx/rZXFHbeYs2uXBbm6N1w3vh50nyVWAzrMznWe0NTdls7aZxVTOe/KczYTYJ
WIHm0eosQVn+uSS9If2cFz3FE4ZCDSZh7I3GIXwDsd8WGFblEBnjhKHpkyN5RNT3GGU10gmsBPpg
ToGvAkzDLtUD5oF8sxGwMzSKUxPXTzr3JQNT2QrDCz8jG89zgahqwirA6OddddPZPeGWUXnTscq2
AdvQiDH1crZg3Oc2Xnu1JOT/R8QPxAY35Di8GNz1ggYuxT0OGfscjqFCehwFVhDPYS2jLwpoXZoy
YTyBmFif9ZFIAgpMk4ZQM50PR95FSym4hvQKB5aMbLX7ci7QXHvukOi5O6brdk0wGIPxDMvzPRfz
VEIB3aMjh16T1495/qPWXjl4iYzh2PY0vR7Xay/2J0A9NTC1hcyhEil7nO8ZX0UWbx6huB1Dax73
3op3kUihy3hGsN/AaT/nZyNHKslpZtqWPD9gBNNKXeU0s/f1SxFYxJxrZwtEc7Q3yTJP0HSZv8Cd
tTZhs+rnKbVQMx41A8CWZOatJ9v4qiQRFSuy7O/RNcCdvrkjI0w413/XOQf1mK1HRwWVL+j63i4t
tI6jj/fWf04Z+/s2qOr6b1h4qfojRD/er+aoVHHugyuMwx7MfYgNz2DuqMdvK5Ijy/WFp8Vx67b9
OPk3Guox73BGyEvGEGJMEQXTEwpJLgioyCqAksqFp3baX22S2c8RiWlpcabMcR+ODPaSuAP0XAZL
PAGHIvBLX+cJ5Lo4OwN3uhi3jW6ys0jfnfh/wNr4oICEtg0/LApK7J/4H4Awq/CeuLs9EqyJP6wn
s+5qOR6W48NG8L/k/G9PqPGy75ahZUHh/LDvPU1A9vmbV/bbStdfHp1q6LAbkVIYc1LGhbetBiDX
Q9EIqyTT8TkrIrg/pmQLUiplNriO5GVpaqp0JMDdljWSLYBBYe0YeuE2TrJTcj3hpReu/ZMx5Mmq
E1mvLMs6xS/BIeWc7DrYGc+gBafcPA6y39l9INiEgVKhEnpqiyZCGkbF5uzpWYjbwM10O4OwlOlC
mukldWriFti9E3eQGLA0mBmewNCJ1pYV9bGfu3ziZIdGLknUx8m/Rgr4WT/2ENb4QYcK9rO20a4q
I5FxX//CzxFeOXWbAhdI4yBTNhwwoeR0coqgStGNJkNTKqhyLlAk6V9392xM52eFbs6PAKoDc9T4
UoZJkGt3R5wEX1Y2WqntmIIizlfXi+03TuHPapXP68A0t2Nlt1WVcbpDfXgrZkxRH0yjz9W5f/ZG
cZELdxsHA6TSyicHR7oeGLKm+sKePvS0o55kPm/rh3iVNPiA5fyx0UCCNoQA8kf1KAFkpmvuWmMa
6edxkmxujHPleTnL5X/cXBWcByoRiNna8h/AHNEoO71jwy5GkCQx2bZYU+61htj1fqGR+eF1CGal
fWWHvwyq7RG/Ky2o2D1YluIdA5AyiS5MGZAhCCXIUW0A043XVFh/EI37PcT3widOt1dNdM8wcsyS
+EbeyNBWGgLBX4Oo4a1YD48yxe0thbgKOWqdLV+1yu6mAGgeW/bB6+Nw9RAb5TB3/jOh0ARRvRl4
Bc5lVA0ooJ7IZTmZ9mLIcvoQlNs+KVf7yglTF8dqbzby/O+heLxvSCm3JSY8XqF0lqlXm3sRb/y6
hEYfR6AWuUj8Y/b1+6YjJTtgnrnMF8UMl7U8gY3/04ANdRP4pqN7qXUp5qJERwGvIq1dXc29Ha83
d6mUyip5qrFX8fhjXBJkfQ23PPEpG1kUjC0rxXw175V3CeBQaZJyMoAhTVywniBLOakKqdxnaKeq
id8oDd63BEh1zyZd1wHIz+L9SfslRdAyBQK+355ruFRojUUzlcBCvCJoNEXEYCLN3Dq4W7b8dW2x
/u+48Mk8FU57OXnM1r2hyBqEchb//zLdOxeTIf99R6AFdiowiUTI05GwuDkbawdveuizVFqj20vB
z3nzEKo6GTv4gRkvVy3rPoWJitjQKwLRT0IPjVkoCAK1Wb26f8co70jDGULGoYr5d6ywTFP2TNUq
4JiUDgCLll4PXoNI0OBx+fSk310J72bfew3V9vwLDB/rgin8aCes+gfzhXQjL+/WB5PoPGx60wZV
Ico5K+py/l3RbDGq8GR+MBC+7r1mSz1YTuTVus5713njh5DbnxKnuPwYw/sjjnyauejBWznMBLof
LIfl965bPy6zH0LJXjJnkH2CDqyjXV7szWF/n5FFFphO2a8UYXPs388LOYDAg4Em9+o5e4Ihuhdh
kWwXp2wTtgx+AEXPN6gQPntLgje2w+Js2d4oWleVRSiK+CuBcEq1s9yRQsuDQxR+cRPJB+dhd72S
Ib/ZKGiowOu2Tnypej/YjpiAwPI2W0xiQyvi6AVF8ssCrj34pH76Mn35iAGrCh0axs3wmT3wgmom
7r8s/QR63Tj6gegQUZdvs4o+biof9KR4hmK3EznkpwntqX/WfaYE8UXPpvISHKhGH5nhIvZdSlI0
u1ZZGpWs4FdTEnnVEspxjJz3yEIwy2lsFc7Vk+D0pRGvX8pkqOOvVfRAK/krZ3M8NtRfbBXvD/73
OfllqjRH5+d56PT8My0C7ala8EsiNFmZyGaVkCLTZMiLm1Fk+/RMVvuCYQ6vBYvwndLjp+gzr+xj
/BA+ygfqBkYkUEXGpatNoInXytPawx5G7eq3O4gXuW9PF5Z4chyCC97SAmz+wEajSSEuzXNJuV2b
oPe8rkDJCpjFvrrdAiNmFhxFbxGrGnN+e/RefGk3Awk2z6gZnEXsErCV+yvLzEk/jwk0q5oyjKah
GTOL837kZaW031L2LMYBCRhVjxqINXF32zMrzqyGF+JSZSkUrkGJdREA06Koipm63K7sKxm5p3GI
gsHVTuZ6T0m+3UaSmHktShliCd6Wi/yha3ruCKGMTOSKPI7K2c540h0Lo6Dtma+2+NTqMMjU4Pd7
y6+QrXN9K/1GXWoRhvgl18A0ItRtOCfHNkCSKffkBvcAMNFila4906tb0uexri8Z4R2Y6X03uvwP
MFaWE6yPz/tDlwMzf3dQ/k2fQEd8KKcXtXBFzHbhnV5cY+W1Y3e28TaP0A9SUh5U974Pum5ReU1u
Uw/AQIsJ/p7by+2ds2fH/UVQtb1pCCBAjeSMA8shs0G9REsAjIE2qmiq2Xr0bnKNVxzSp+cTODOT
o2rtFzWwTxjEqbPRhIfXJt4I/pWxfk43mCLPhTtaMkIThioCRdSyfPHJodKwuqjKtDggpncDDncS
RppGjGYYZBy+bt+FtkhkBia8sLDwqdnd3k5Rag5Ncc+xAfH2YCxoGWsF1KXA22U5AkKdztQBf1+J
gOxQlQo/idifGQuOy+/Dk9C8g6rHtv56rb4Urwse8ndcRTY4x4BkCenfo+JcCUau3lbq3Bs3Nse7
9El2HeN2OyPQS3cvV65lRRqCZL1EWSbVjP+VLpQSHY3BYNBtJeSHfNn1sNWjboXpoeTb65Mj0Seo
Fz1KCf/JVc3/Krf2wF5ghrOg+2mGw3hRAM02EUVKu9NvaAHXwdNMISkoX4Fj18RmDuGtIWE5SOlN
J9w2PUsNOc2qKiAZf1KR3bR0scw/PAEIO9ezql6LrcZG5B3ynatwJ/QNi73jqiA9I6N9v9Q+7JFg
h7mNOMK2S+i7u9A0cP6z8noUWXVUpRr8x+uTkPD7CVw0/rnHyNBXezaki2VBRQ+pz0LKAd4YfTQ/
UMPJlPOAiFr+OJrRD/pTrkahbw8dyFrsmBzWupxTV2SIN67J+Q7swTnGFCBJrNXKEDNjA6V6plZf
8mNidbRXoQrFYpVPciDLPwbSbmLAqBAZkcGiwvqUrLJR0TDHJI2fluZLCjv64ALHcI9p59yRO6li
iv+gpVu7bJIBj5QJmMkBk+KlR7ebFZYf2m9SsxP4XT9c/hOhlF39XomGYvfnpkYx+VF5WrhtgQq6
INl9kxDAibHexVINfk5T+2H6LiwJSsmzcUPrW8DTf3I4iGp4cW3DhoScWoWc0HDy+1im9wP9Knou
Ykqi6dAqLuUplOBY9Y+h7UAyEFUnS8/MMz9bH4Px49GvvfcUB2n7rstis8iWPYzbNtf+LnSw5yzR
MpfP7k9IZV7wuTj6Oy069JlVk47mdchSsHKVblGKQzHmNiyGczqiR9NLCoBwkP591vL4HrfRGEaN
X43cR+PDZIzhtXHvoh+mNUQGL8mgKvvsZ9oEz8AC1hjlMJfiZc4Wrv+xomiIrESTJUxWjx4/robj
Ui5sqQ8J1eEPtFpjhRKhgB8120X3mkfYIoRWGNqX56JknDFS5/hfOprabm7YCXWG5tXvG70pbH3q
NfuZgoPt0S0rFsouMxyaXc2ND76iWdm7y6q1CThp+LETDfN09549Oufso17sQxM8QUCSXxuIuFLV
pRbW9iiuz4CkiP3y1JGIMctCK9xieAvv99SNs+ihIl07W/oDnaEOIZpVS0YpRgpyfZG/CqzpIJuv
Ao6eGGL2ug0+ROsnfnuxMcQb29LKrHUcGumpbwhQOOj6M/n6dZFDlrgYuIVWVjwkOxGfXMUJ/Nxi
0H3UrsYvcKizPfbpob8GGXqL4Bv3jXoqKxpbeuV58jr25aGTPh3hxYw/4v8hTB9qd6uYRn6kH9LE
UURux6N5sea8AuswrKK/TRs4Hs8ds2dTyUKhyXW/ZEJf7ZwjKtYeFPbi9pDWJGUL6LtBdU9ztfWY
d+T8ZA6lVaLauQqy4NiwsXqK7qO/HGS4JxQObIpfk11Iyi6v8hN7yJOT/E72jZtee8KVNkgDPLro
xXT7i4ASqh7y0IaNBwAkgRh6MTZmSztImY/4a7sAli067FDpZ9zFY08kFBRtkKP1y9Isl5RKK1bb
CtxYoRlpiMaLWD3WuMRKTaidrm7gOWyE5/s5SbB8sunHMFLqfAy68fMa3qyhdsiyOljUrKIwik8B
GTJuadTklV54TseVdnz3IpOLbtc11iBkcIWZLALjK45Wt0syUVtXA8PhHMJgIP5gMaKgO/wIVF44
RDNrAgtBglZw3io0qeObwAgQS0xbOfRWxROq03RqZg91NJkfuU9BLqHIr+y7BSoQ7xzpUBcKPVVP
OWqv9K1LS0L2o7atDwTP2Hf4cfvLs6mAjtUIyGgN6iG3FW5nk4ZaBTTRMreBjl+R8aTae+1GawaA
omHStafEDsbbobSSQH0EEArvbzjFdZr+QV0JGPxPmD9V/wPytUH1lY0yOF4Ha3pAPKuL5p86/TGa
dEAJZLoiM3ZiJp7y124UsPbquwIobISuOJe3gNYqzHm+7A2sTcRLYbDNBvN124La67tzH5xAtnBc
GT6cThwKiVTzV2YCfzDN5dWZXs7kXdu/FJPuFm9Lo+UsdgPQSCXpobb2roFE9/u8oLatuhm9cpzW
LnFaYW0+O6uBh7U089q7kSoK/KTJMtJbsFY6PuGimC1BZ4RTNe6QA1UADA9rifFAghLAMAb2mdOM
ALrOWLrWQy6gWG8tqxupWTUaO+HGRA3J2+/yVc0oY3KtJ6nWgEQ0WYv029zRte86M3xN9lU0fnGM
HupTBB/uUHGXNxHRb1tg7uL5dqMz9aFVfA1Uysn1HSZ9X/tpSS6Gcsi63L35RcAg5DSH3DQBClNU
+h8ngzrUzs+muhGB2jX0BlpsslG+3d03uSdktyYvDNavA6ryBP4F128TEp5WVUhIvze2RoydcoPf
iT+XGf4g4Vv2r4hCnPQuc+C+DMPRx/oSeh6jPQxo8GfS9Y/1MxHlIKIuXYEmp1+U7yLN+SKzqSDn
fjj6RvvGKS+AWLhJVmQtszToMaTnJdlgzmxn9HZN69uh6CTlJj6X9qQzHkhve3Cunk/N0ibbINA1
YkMZAGk1kb+eCXPE6SheVe3DyG3MzTUINoZcSNGpzU34Xiw6TUQRmOKt3toYHykrVQInrZj+6h9g
biUmbJm5PKSadeDtaPC7+vglWEJJloOH8Z93F1Xh0eihonIzp+iilSEpNxd40cVbbxUPiXMP8VFz
wm8zUB7aRTsrCAssr5BC6mxhTdLJE0fnBckvpLLpJRCs1X5HksKlBivmboTDLErxaakx7kAEi5tl
F+6iS8IuoEwlysK5xcboB8X2pCAcXNcc8W873re/wB2TmmfgkM0h7yJtmQHGz3r+m7lrOg+vt/rg
DauDVJQm1Krf1w9JkIDTqX3TuNqRJ98FaBAOW/lOFgtbnGzP5kU6D/+2dbAvEuI1GSFdTcoUnD6v
z84JuXziudUJchFpK0+dhuuYKcsuN59nr3vKCaQ0rYfneeVJOkRBm7m8SP0bUTV0pfwRvbXQTcAc
FvcV/ucRb7xn4YNneHQ4iyxwbuioGXfoJ+wAEirmXfiLxsWCIM8y7en8FQQHMg8GkzN+ZpqM+FDV
tv1KivCZXqRqiXxSJcbVlKYON71+Kx5tULlQLeENdXYtYWyiqzSfydkKGf5ST7gfhx1aQ3Xg/hWi
yTxqEBR2yWPGfV1VeoACeOpvi/EM0PDM/6emlNfQwtHQO5AMI+6N2ZkIyP6oAkbwS4F1rW8nml3W
ZSt8dE8dot+40wKXIX6pjOsIUalTI4w9kB9G9lLnCILxdLVt0IGdQIf/ln/RWvGxML3k1GQR2wqV
t3dSiHiAdBELCPkeQUM83BZYcryZk4VLgNN1GSvJejovcRYulPCL/WDCMUqMLZnbTZQSryi8oQOw
cXHaEQHjVf3jC5VMm9o2Ku3NW/I6V6etnFmNRL4j9MIJNGyRoyXJSmXqFX1wNRyFMDj6dt1ttjCe
H9ou5wh9dPlJeyiil/JlZ81Gtt1TIh+vdB0kAybrEAhMc7RMcB8/Hwoauem19WEtvWkP0FhAlxuI
HLT+r3Ou9cPGkWBgiMdaqprrHH3A1tV1B/2KgY2h3IpshAY9onhG9FWQVKFrYgbyZrIalJuRRtML
VdfuxzqIQyMgMCnIVI+hzWBLydqDcP8IRyPNPMF8zu5YbilXoC7hfQoR5OEKP91EnEQwS+xHuy3D
qfogMhkaItLmQS6UGmqbwJccttyowKWBuOFKePSHYptkW6XGMSk2Y0MDW0cy/APRByZKz0tp/UBO
YQW7mQ2kecTgPoKOvcQY3Nu9qDG7kCS5Wv4UXUy8ap9cSShgXUYC/bWAiEujXD6mdnLG+Ca5COMk
LBqhJaB2sLzLVKoxqYyfvZiRFkIVm52gg/HuTBuOFPffdRaCc6z9PPSDLPVDH/566JRMR/G+HNBU
9Mk4vpGYwP+T4cmCS+Zxms1w0eTPIXr2hYDXxRiX4rEo5cu8G/xXMelAdxdwh901vIme3XoGXRHu
vRDtrb7UKN3CdWLMR5gdPbaX6t0qw+3qjILl3nnAg6K/EGuYS7YtwkSiES77LoMw0crVShu1ODYp
+J6MQGDRwqGEAfYF4+IsF52vblKxrfVQLrbuYqsyNaflE3sua4WP8ORBQUTMKOegw6S29BdAdRRT
RlKWzyGRn6y+qs4U/cMSvSlW2pUQNvNz5ZCRNkE3ZOshKHx/A2KJIJU3Hcmqn8/UJ6wyIIBM4J+v
njwS8iK6qJdOaux56pMg4RLQYlUn7kyWREVXx56fmWmCkaRzSsuno3IjiqjTQssjPkqCzqwKfpQJ
NBSBv61+Za/foL8PsiIZH3qkzIY8JBH1N4rH2bv1JsK+qxbaa8xtSOMUktmTje53gej6qL4xn4eW
alHg8psE2f6RkTNaQdwn0GxLwDQw1jtSiWkAeJ3sT2bnKc4RtODiMgVvuQHMClsA4pBMrkJ0fhCT
g5iBNahfH8p1NnGgvu7R0sqPLCUaoLm2+7a6J0Dp26dVYMr5PUx9owSKPFTPP7RvmnZGqZBQBz0P
fbkqOA9Z5mvqH15uKGrP/YOeeKzF34bJnjpTZ8Wa03Do0dwtA9+Ru1NnLax61R1D7HvpTRCjw0fu
pNEMb28v0W1UiwfFGyQZebn+3SHVYWg0yW1SixgA5tVCf65HRqyxgVuyHRZibvRCP1iX/FxzO4Qf
bTer2n5cEjrPW2S6SCvEIdIHBHibPnHqAqj6Vy3/8SB30/Cg0jsL/xD3XrCzhTvAylEK7W3CytFb
v9y+LuzDtd+5jouhOvUbC47SEue9DC68vygISk1QQi1yUYBYslsIkxh0RD44QfR02uen1BvPySFy
gn5uA88U53ovbeaaU7bOF0xMy55DEFVbN1FALT3WRAiugVWlHdEvdw4FVD92Q+sCpcOcPtX3zQx6
tm5p6nWeiRy4RpB2U1cGyL6Pcm/uF//6v1qN9GQy55WdyHkTQURnQ4Mc6HmLw4LIVh4W5Ie3tpQg
HhW7Wlnr7mHNQvko7dV6IhiP8FWjz1PSPxividwB0Lyxh/ZgJzZqMBx2vft7rpM+Fv5jNcKDaKlU
5xz3M2qAU/N5WEnmQG35yJhWbUu3dcSmY7QTYDeNuJh5AmYzblDqKkSLLWX5dfXPi6VX+mAgAPVb
T4q1gYORepwbCA1oQTyodlNPg7G3iw8cOmTsTBnZbshrZzCWruCtVnc+hbbHVKKG2CjRIm7lvI05
AuWn4G6nQwxBEoPYRzmRYLZHbcCtuj5YG7SYUzVuHY+UtoIR96IyHoO7eJtAN5BI/d++vKKE1+5F
nxkQFCfqs3It8aGl7f8sTe0MyAJum38kamEz3OBof/sCE7I6QkLDtY7ZR1zvOBSN5zadYQmm6xpB
TeSG9C+kKx4Her8UxN9VQ+D9xMH8/JhFQZWtTvXYxJibhkBMKvwDLSxjh+nuxMFWnArexkCHOOwy
3UfCu8HHtS0324DgmemdH2XdO6KnYvnszm2c3LHh5vompGJyFqOiVtMS3EqugjvXa1coJZAszuOg
DpvSE3PhjisL22FOYgPAo5aWF1qcXAb2mTEJFACXmQ+r3H0AzM/zs4IJ7GxkG7iIGYb3lvCkvYdn
zNS7lMguB93ZLqzV34N05UJDjQhZEAqkzlUgGQSkv4COnDEaAzXYLIHvGOY1xHPIHyDlMtwNGNsV
lCGadxPToDvH1eTx2kqZgZ+aLAsUijq2jR5/raUmBtpD6a2V83aa2MyGIL2UUegeoMwNwc4Xs1dV
ibAJPvf3w+cHhqkyc3JVKlyqEeZ5317akPO6MoDfvI3smdKNBVybUCJFvdNcCQjsJvOQKMtqH6Ho
as1AEKO+TB0C/00QDuyYm3w7223SUUIYS5+ibHjwHn6uxOJoIk0fv0l68vnrZ7MYAfIjY9QMri4Y
2uOw7NTSRxzYHO8VbTQY2W3O4vCaEtE8CXxToz7KYH87zL8AhG4cHmDSWhIL68KgSbTkmYu4w82m
gx43yqhh3xeRJRDvq+0cAQZKYc0q2WQf743jDDRQFdfFQAkphJM96P8f+NreNDHLUr/lez4n8cq+
DYyd5XalehwbLH6I8E0dIL6Ayv6+hCgKJ2PP2c94PD5wBexSML5f2b392eEdLm9yXnr6F5z93dYk
EBh8cyTCbppZrPjhx0SMAg3WEDxKpPgqknvKT6q5tpQaYb0tCrw4yxoK2BEy4M+wzTX/yQWqrpso
HMuxgm9hm0kFUmArtLpCZjGDwvmqhUckEhhtUsvbWSCy3FMic0eKmadn52t+hzCBb2fjGg7/rSDO
K64BtSKcrRpEia+y88MKg/KD8SKNAf29GWSyf6lp2oVQv5uXjaCCuLOUamP2KmtF54cu4IJA3tOo
awdmdvriPDi1pMw7c1oXef6T5G75OYO+Tw1e/f5uzWV2toXNEpnlI8ACXuGwNT3fLnENZUjem0wj
CehErv0qL+RSZ3etbtIFBvznSPbxFQLVzOAMnGFaU5tMNc85x9xyljWMA+RHpmL+Rchrb/yD8xkt
T5YEuadBiLghZ9AhI3hyK6ZV1ncgwbBwezhPk+Jz/nbAKT9vW9OA/i+d4PyaZ1xzxWUPYG5oIjq9
FuVrr4MTNiIofBSlE+Di/SvLmsqnDaHjcJt+9KE6w8FkcUvisQ2Sew31j0FjXsP/kbiAdFvZhk0x
lJ9ucWIWRSwssUuhJ+ov+HbvBOqvWmiU+0ZGh8jcoaf7qw8aw3PfiRPbrWJ0hlizrEkxra7dBoQs
NF9k9x0Z1+PN6VIZezKhGRJ8TXGKuPb0fHWMmMtFAqWIRNpJwqDExF2rdLZvda0tWzKDlx8fY+I2
ZC+Z77pdrZyv1vmWoz4Mi4by8dIe+n0jus+CVxKCN7WuY3Sp7E9yGDgPb0Dfd0nNksLJLbZqvFss
eStIfRd14LIsFRK3BtbsTGK7wRs+IubGHHiJ/gvlSGke+iTAvFdZbVPVzwRFswzze1KTU8GyO0UE
ACa8tmYVR8Az1Z4NzefGbJ3Qw2tRJpAxAtD7azqEba7bq/qv6/tzIYVgbmWWuWN/KFw4ifrUoj+p
oOP9Bh03hoZKyItWhyFUgRRaxOiUaXOdiZV1WNlaoGSKnapaNsX2DKhRlClhZMB1Po2Oh453dACh
ywvZwzux7Akx0lcgYw/DILhaSIKzR4h9e+0q5R+E3zcBCxEA8EJagQSsmaLfsB3gSxeVEGUQFLKN
PuqvNOJ4roFMiq+aFBkMoZ4LOYpR7UVHwp9zUMETA9zcL//MTCXMy4pqYsy8WZDF4ceMRaqbavxC
fskZPbE2T/NE9Lf3L4L+lxtT4LYhx4qa8f0ebxPMisWJoTYAW/g4kreI3ma3oljcSkRPx8dTBIvM
rqx+LXEsbpagrt/Ea4vSt9FSBuhBSYjS7sY0z1TE78D9pKkEYDOUgta4eGKarD5b2zWDSGJfyNIJ
g80EvrFPwFVAFyohOnM/jheVLXB2hia+73Wm+tIZDJ8asZ1qm26D583rs+yCoTmIa17010Xye3I2
mHQm75hp7NR9vRcxURVs3x4PpAWdDYvnsiL/JoGlgw4FScSQvrcB4bDjK20IXplKyfRXGtzR7PfB
bt52k5cChE0XLboUN8qqmAuGchiJonbiUqCtWQg8XjNNhHjBjyhSPH/OpOtH6QFldFhWKZ0YBcO6
kH0r9QJk167BCPQW2SnGNkwpkoLp4UGRZw5seHYyJOiEK7CbEjQknZAOnphtzC88FC0pMzkeVnch
oOrD781JxucEU21ARjR5ZndCUIEIfXogmQqQu8jZZhxfU8q5ibmX+KhdNJhPTG3qxnI9n3BeUhke
HRCq/E1Lekezp3EDQkmMic2FstanwOtBpp8c5tQdSqZJpmpLmCm76+lEMPCkGiB6C5fLUY7qhGUE
kw0Z4S4k9IFzBNxB+3A1OkfC27nsi7rZFgYZOFvJM3a13+7rbVEmunCZzHwkBTahLWulMymSNHXA
kGsfDVs4q3lZ0Da+wnhYNzWvxKNzErIJI7JZFjDHrz6biemzG7FsxfYRAim/PT3RuwA34S+jj3zY
8DzLMpr2xlZ+wO0oJwJCTSHeK5pNQb2EMVf0N/f3NWwhIcc/lQyL7xZI+fmBmg3bVU9CSkFUu4n4
joc3ps9D0L8ZbrTvbMrGmacBrPrf9vNTI05aCki/vIkizW/MGjyoU1PA5ozVHzt+vCwFwKuD8uh6
FS6ec7aUmjraJe582WvVN6a2/Hyzf/nH7cpFgfiWlv90XgVT9K6hEa9oXwHTQds/Awyd0goCpiRP
+IVOf2jFZFqlmOhkiBL1YutW1vy7yJHX2/TFcQop18HKo9xRTYMRtC2M5thKX4snbUE4MyRuHO7A
54DBBOvyemxYaXHFrPvqSru55sJCxf8clES6ndoGk1c81+K65pJZDI0UXXj8ZzeleoqqGggQa0yL
Y7rbB7gZ3YxNfNjNK9f1zEUVor3l8OTVofdr6JgNMsPcPVC/noZjkrpOMpViAmNm2lQNXTLmfrap
OtfYF93+kqK3S1+NLWUT1dSpVdto6myQ91P7QUTkHPJhe4DzChnqniHj5cYvQ/bN+J5A9WkmXmFM
3/TXOvv41a/98h1tWpKSzWeapVA2UssPLcwO6dJmOyxiTvpxktTfxAHv9njrRUUlJf9CsgqAgkwT
W2gG1nL2xtSJiF9ovKI/jrDpUjwYk4ClNIWpvkwfkcnNSMiJ76H1B33AxjNl2EP9rhewSASCc2pW
BWN2OxIPVP/lGmNhMR/pREOt2sTe8OElKINLaFOfuZMCtAXJLyLNAGDNF+x7rncquH0V668MHjF3
ju2Yyon8Vu1ZKauCEXDWMr1wbDo/LIxo55Am6KdFXdVEyKlolIbaYRUnsZ+30JJfnWt2B42uRi0G
c7AB2XP8+VSwKg42QMjY5vJXfF3EyeTMujATxpGsuYCVvyBzvdA20StWzEdyMu42V1MQJ367ayQN
3VIJVA81yTAFlvz2pMUNPoPazlmnWQVVZ874N9yzCqBod/RnOhH65+PkQAmzLTjWmpORDVikXni+
NC9wheGKWcWgmOvHazNZeUBe0ND1cXxPQxeObmglpHkVLgk6e8S5cNg4r95s2FLcEp8eXxriBHaa
BUErWpTwHB9wNacI6h+Bb4Q3s/weyqoFVbBCZmOA2DIDJJHbstsucy7uvDRl0d12txHs054BhUUY
tb/ubKP3kJF1eerEyX15j0gGn6d1Ygvg6es1aOyzsSjgZDQ1KspVy1gsKOHiU6nUs9Rd/ztDeb4A
hLXjN0GtqaxrH+Vqf/EKRPNhd9OJxamgvKCU5Qk5A9ceiuVkyu0SeU8o02nXybZpKzNX4M0VcdX4
70lVNPCqQwvxWn1s754wZW6QhOlxf7tmwodsQJRYXsSZbf5YV86OzEVBcDe5uB4S2lEN8Tfzgwac
Rpx664rJbPmQX3/9Tu/htVJJ/KgNOxFzCfpzyWjvFuVchSCt6LFTt9hkaRaVClqH5xhBjRGa8hhV
IqznIdsKRRyxhKgVaUjnam0wTQcZSDH1MLtmixK+CuO2xa7yqkAs5QhDoosKPn29ezMFaLfpeds5
R7g5xl9sN2++/cl//tDa8G0UyXiN3UlOkns+cjuyY7Udl3PrCMEK20zL+bD3sK7p13xXl5OyPWgs
RreUwDUwD+jyc+PpkhVvh8sQDKKZfmr5TJCvU2f9bQy2hVfpa2+L7poGiSzMVSDRWqcZ7T59/Sgj
OG/VXqPUHd2k1nwZFEl8XZZ3YzZC2MjqjHvNMD7lpLofGaXu43l0u7gyjqgmTsP/RRuk5AI0GtzE
S9ZTTwCkxGwF/ZBp7OlSYJOeWbUrTmXktBDDlz2iX4vLjqJtWmSWsw9uULhLANWFkKyN1hw1riZn
TMR02u3QMphnsdWXaKgIGaM2ujOldtcLWHlQ3GJD/xhJy1u/fH4PJER3ySZGPO8IOrsVeur2gvat
syiQRgxgAek9MEefT+8JHY3W4pj/yWTlVR2X57aiId5j9KLmjV3yRhcZ8eSyBy2c/8a4VHXAQ/Rb
cOys/wuCvpiBJuEBX9tBwUVXT0/8EVvjy0hDJKjKHXO9wTHh9lHwOcaNP5dOoQzBruVTDs1z58Uc
JQFm2oTeXxOjaCParGwjkbMCapG4fEY1q1rQv7Gs1aITXH5OSItGgQpi2helBLJtCP/PoJx08oiJ
YYcIa+twhSWiwZiYEntWOlHaDMcqVXLlqd7fX3KUH/p0o2iaaXnTbFwVOfsMha16PKMz9qnUFH0r
+2KboBZE1YRY5gJns2vio3nVNTA/XqLT/kMurny3yjY1rGgVkLMYmu8BnAq8428FFOSGQXfdxDGv
VB4F0xQGBJPvXIxhSyMn83T5Q2id/7oi0JqtZjc7qxcHe97PmUBxejag4dTcbWhhSOU0d1PyuqN4
BWxnHGmlhgzV7k3uPA7haZyAQNoEKRwTNlollaUEFdj6eBYcZv8tDmR5kiCSimfuwgwE8DcEyYYj
N06Zp9eq5Kr48upJKC/MODjSpmDofGqrs36Jq/P9ksZEa1RIHelUTXclme8NhPkhQIKT574dYCBt
ZPzPQroNxohI8YaTtvQNOd1qh5PvwQN4SW+68lEFNHbRve9Q4bWMUNnD7ur9NTRVakHiFLdU/Ayx
U//Cc+pIz9XAYrUVKm+NS4x7x4GywN9US80yg4B4OFz/tSYhKraekFvqnZBuC+cN7/OrBSORCyJd
Nw+WVHv5ehg4usIZFPH9h74GomwjYgyK0832twLixKZQCpg1sNGBiqAApw+65jmBXyDazaBkaeSG
kXdOhOoJCX9bGM2k/QX8pIkdVxlM/K9thLg53qKU575QCgTkKvECaL7II3aRzziBQK3eh/aQPELS
xjt3Shc5F4DG5hyhxgs2TIc2llWAK3lz/J4Z23ou6kgY8hr8KpugqLzM0c9cFf+HKxUAf5DVJnfJ
vnCPt5QV0Bi0IprrD7+kScchpiXgAcVkGr7kVXCPVd6vEXWMDX9s2HmD4ohz6gaFsTIGm1r2poSq
S8yduda929ao7j4fdLIIE5WZYfx52h1F+xSy6Tw4OJnueRWSEbkabTUEVAHx1orsq2fbIgxuQlSj
0xxefHXZX316HEP1oXZSUe5Gy2CV9BNAY2qcify2XCRbzi3rCIk+ggjdam3/OnCdq1j25SsKaUML
8gSicxApZAFEVC2F8BPKMrL8yh6redIK4FaWh5eaT8KARXBULCaKMRl8YMSxnpFDmuFCLdl7VoxL
bfrC1FFL4TCKVrO25s+9Rk0QAembeYOJ70KNQW22S2jFo8fmZdpnr2wKB+3fxnqojjk4eD69PifV
XBeyDXY0i7XqjyT1/g3z4J5rUD2AqHAqrRJiUyWYva6uW/9VsTkGY7aMkV/5YdjFSnu3pa4m16wI
iZspSh2hw2/Y+NlypoiT4BkqL/0zKk2cphhbX3LjpsruR0WXeC02yAOqHDFV7D6h0vuJaqQpTQfA
J0VqZT125A0peZjB0rF2wxFI2IV+RClZRhPhf8OL9qXbBhgvQtN1rYCSjZS3t/hCULM3I/Le3dqD
fak01y8WENRO+PLeIZr1KOq7zlvuP64Hho9s6DBCdxIv5fZDFPV9vVwc6sa+sbChsGsE4u3o91GY
1NRqjZQeyIuyDi3Ey/h+wChAqqma8Y7KhuVGxTyrEBXmqsWLiULKPQI3rOuImGp3aX/ZkXE2Gca6
jaCAg3Y/XQY15lD5/2i+EWoe6/9vaHwKr9qKBjNNZLQcX9uOQKQyTqntngHhHbE+wZ6xI49g/6FB
/pcm9dhLfiaaLj0rRAoAYSd6usTrj7SP1jxTa4TnItXn+Av/lRA/W5FJ/3FDdcqrNlH8T5Bj6HO9
Ln/Rs+7UdpOvf9gMkwVrL9D7mj0l+XayYTRoWMZgjVDnU82uX1uXTs3Kla3ME/z26O8YKvbAP6vQ
+koLfi0CD2oXvmlAfojXM2NhFSs/dBvGdsO9qChLaLVKp8IkdVd3vJU0+4LCADw6JiixlMfQns7p
VNhbKq4SOBvCig/zuRoOPUf4cklRwjrnaO1Y/v2yuPe+cdHs/+ynermHy1Sca3xxidwZby98bIu5
vrTM/62GRCAmpCbe43jEkrZTuFCwTnUuldera6M4vgKnX/Jm0HklooCUMwVA5HPwkL+emu72DhLQ
VKy5NWHSVpX4JLEsaezUnG3/ykFpfLKlu5ru8BxO9RTEp2QHOFOC+4rdr9NIccXpJGdjqozxcVSP
jb9R2j2A5heCubATKnpohSXtTCtbKMCSzdetmD3eeFlfPrN/YxQEMELWocKYNRp/F3ZF1xPsPUOd
vRgfmcKU9PNV1qT0eGtLtTsyDKhnYMc9XSBuJoVt+uVianzVuV6tvWa0JeYsHhRkBYG+dWdcfbt/
l25yhokwxnT1Do/1hng0kI3c9ANTjaonui0ZVbpG19WXKfwyntaNIInYEWSrA1w5u1AScwLKPjwS
2bFkSE38idDUsWvmnCyeGErFKIQNPPhUSfH9aKdFrQnQo3ktKVcxoEKjaPuD81eb+fAFO5OI1ebt
CA2iXq10hccS16LZUVVgQ0SPbJr8BIsRP/xYmVIkLDWJxLhfrp27K04DEEEnUdmrfLXDV3tu7WSu
bdo7swqb9MbXvd6rIPvJFjmHCpBVhOUMPrTjIdiUzfQqPUB6P/kAfhJgz8tsaYSqkMPrE5mu/zT4
1mHdWK9fMSJY1U6RUlWaC89purESSRTesVjzhAGaXXz3yeQqYTB8b1SqazHKJBHSCuzp9Ns1kuhI
Wl0j029hSP+lLmWcB3jq06xXQiM1zx+SpEPoDu4sbiVzIIVatVp1LuyvrYPDgBVAB898PvTB6iCX
DoxOi9C8bypDxhluI3ezftKC92m5sOZ0hfH+oqPsBkl8bOL3Q0dW5uGjXMOZwiBWNt529+JeBGOz
YF7rV6o5Z3Ly7nYvyzZkREt7Ktof61/6IKsnuHC5DxU3NVvb+fZeQ2bR4uQ5+ED+9oFvtW4EwdgV
LZv3BPhsdXxncmS0U95sXGEWHMemEDtyYjWypnhuSAeP3kMG0QLuMvkx3uNMd38ZCstIS3Dlmst3
zy40ebo7taWOMl9Zua4RtbbusdgetAbD4CzMPadOi6YUeOmHTBJDZwvWgUwkcMYnkzbCUaq47WqL
5iYij6U6sTez3RggzF2ZYpQx91klTs35FpW71RaN6smE6eehubu/kKIO+cPr2YlP0HgW+hQLF82h
hNk9hJJMysy+WXRGaXENxB3F8x241qbII+/7UzUpbDWpeeUnIhmwAhxhUpZUknW0X18hD7cYP6Vv
uklQEhEZwDsj+bfGqEk+i43cF9ZK9mDXu7cIEp1rAq6tzR8FqYbkCcNXxZEaXVZsCSdabE4UmA2Y
UqJg0GcFQWg3/+ys/2aGzlGcA7hiEi4scK5Zpyye38AKy681IZ5zuBzRmR99LOsz4a6MQnqYNBY/
3RIhDfx9H+sQmhFQRxAw2qRAHrE1iXrbzQ5s9quix1tFRLI6XQ3ymsoTA/CDnxSlMFhgPMMuS9wC
EFG2/xK4J7wW27JG0ufQyZw4PJ/LGTjlTLOIGXyf/EFe1yNwnIzwGxU09gBETr9/nCHKPI+ZA776
UL7T35r5/e2IwN5QRjEAccb11as2MnZM7wtXkHhz39Wq3U6tDrPrirQv5ib9fLBxqqUGSyCkDVYu
HW9pa8voizpt6Gkrcktf65K2jv4fHGKK3wzmgdzCpDwdxA4n3MQ3Vx4zbb9Tz6x15K8WnB780Z/W
sRZVrQ5GegaK/ZqB0zKS6aogCFBK6rG4mOEFbDUu2BDREJKwAeUO5e9lI+RWTBUSejpSO6WCfZJb
6vwtO/Xaqy9mHEn6ZD8ZVzGY+/9fjRi8AINZ+5uO9DK/diUJ5VjKhKLnR5SHxMBJcrvvlnRqMXA+
7P3b4McHz9m8FLU28PoIGXPhU6bZljteda6CFzqWV/GHRWghJohm+ejwhxv9bc5BvXFukCYLO6tP
Ucb/xWNWs0VVVPMdZPxneAsRgw9Iea2M5NsyvldjAaY8tqbbBblPsHxkrbZvH4c1rXFTbp/RBBWi
9jeg3elyQHWc8gYoAvgIFLx3eC8RbRw17APg9iErhDfx7Lm9A8dbFslnC4DMvMItZPSHEe27aekK
3zOb5zuWnlH9mn1M1qRDaYVmH/AnvLVOqdk/J9D5Eccmk2LEqgGUxM/oh4VTTnKcVahyv74TA2Yd
dUD1NrYcd1fcdi8t6UUR8L2r6jrPI+ZI794ddgLtOgE6BGp5Bhr/hDbXGkM0CO1qicvzTl90WXBq
kP7GiNkRTs64sodNhLe8bcMcttuy6QTJe5M5Q+AkVqvsE+rB1owgrhFSp0sylbSv5CKJRWyRpA7I
a4QiSVeACVesIiAohHJvKoSACT3DJykXlm5AxbdkFhCkh3BikCsk7iMvpj++YEtmrADuG/xwOkPq
0rEjmpstfqNAKrZCdB9J4bAjht75K/q3qvoZNPlTLiBNXrz7aWnbODK/rOz14amkIv3JveC0EapW
1r/s28AaNONfuwz5mejIBNJXfILmJjD3izFpsmWwFypmYPGgrzcmX02T34t3jTCuNhr1fRZSLK/q
OfvbCW5Bby2MUWe49in8w/CTgZCjYxzUy5Nf5HcUK6IUUMzn1nGUNxAq3BRKStPYMdJ5PxLD+ijl
u58j6rm+vrVU8uDpvyREFP0ztC+GKsbAoy/SucKqyRvbRi+NDzIsYPELpcSbX+iamOM9HLi5UUpC
cVVRY/Mjz1e94lfTapMYhIY+wHGL92SqKgWmjC/yj2LsH4yLxr7Ickowq+b0jsWWaemlx0eJv5C/
4H4tjeJb2KtNaXI4kRiZhvsxqMl3DYN+umpJVUO2+0pdXNH0i3gO30iO318EsOhHfXB6GVUBbGe7
Ls7/PxIftc5eXCvOqbLldbzT5S1MMX3fKpFAEZWjCbpq1CppsIqBj5ZCJ79tFZ8KErFoj4dLYe9G
pgPRKjNHrzhy1yqD8W3ZwcVjgXHW9pG77ccebnxaK3oBEi289NsXJQcFXpcN0mRjiS+4EVMe5PlY
2P3BGvuDbYEH2d9G+ShsJNL/jGBcimxD6BpM9CfOnfqdb9OUNkGwEo3cJsN/Ctzs360QGEtd+MXu
q88r+L8jUASmpH2z8WaPKGIceUvcfHHXMU44vzC5vUMarKZkTq3iISDoafncnepQReE0VjDJSdsK
ecG3Pi2hluOlEyNySU4WGEzapUR7fZH6UH48Tia4ZRTRifn5AEJsiLyo4mYEVfol3iNiX19GsTlL
H+TR1U4w54LutBfsdQbOq1x0U1H5eovsfkz7588bDBaA9fMeKi0zresosDr3PmLxBgUG9FKf0HVi
ERGY4jBMEXDUj7KvDY0VV7/O95Wh4UQZimYOBYngb0cXG9G2uh5ondBgz77MfzY4v+NRHcGLj1YU
WNeDJeXV8GqSX02uCZ8uOyMngAeVRmtcoHnVbWi2+Ox2yqh0WIV8Rdje5zOenwZBL1eOQkz1iG3N
QGUj4bu2cLTK+sH4rak5qwJs0y6gXNlxQyQ4b+vlVjSvxBTSCUn41xpi1TKT8n9tptrn0vNVf3m5
LTsdQon++jO207Wl+GfnHY4q6rV35QcEtl8Rdlq3xG0M5dqmEb8L3lBc2eDn59JqPplfxsSqLU4t
2SjFgA9rNztUve1e6tT6LxM+CdyDkC2R3jfECZ1L4y6bZ0ZZCHWNByKpV/AX3t0ywnodlUixMmp+
E1LysZVQsPac0v+dR30f0qQBvu6P3roaNsCzHmIzNLAE030GmJM7bHmjjxIdtaY3j9n68do0zshC
sx3xPAEH7+K6a1v7c407I9Nf7OJTELbcrRAqvmJKbrfUVPL9uNhqYNU4QIG00+tnJLywTUWDTIgm
FNhbT7uhiWhYBfUichLyZGwPoSUdz9n8/ARmkoMisUnyAf4p1T68mScsSXuFtpfe/a1MznLVwD64
0v7KNw4Tl5iuFf9i/faPC8h6tgS1+uroGWpfpeNKPNNN2BxaZbGpbQjy78YTrR1hJ3o6djiSk1Ln
RxCPYpW+eqasNYp4R/aa5sOHo89uSEvazwJSqV6AYAGAdPEw0XMYU35tnGt55gLJjZjR1lkp6miL
b6/Xe4vYZk1mXf+QCNKLHbo4H66Bdpm+QwkBO0Wn7x5BiIX+g2UjHJCMDhI/O3jQUORjnzXWJ6QP
Pt2LBGqV5Vp2hqmperf0c0vnta2PKWdR8mN7meZAM32Wxs+RxLpe0IhYvsYX9HnaKpWlFW/1EQYc
uDIblxEnWBAS1DP1aFgVxCj9G6yQp0kvBoetNoefFKt1MBbbUfaUFg7fpANRpz33wq4+SXH5fHD5
nrEa8niayXbrw0emb70zsXqezVLRGhe1rPN5u4CjByHCjP9oNSptuUFonNCyU8cxKfQEgO+CqvAa
XcjtT+L2Btk9arJehwIoamhw9QkdWbnVB7JH/450ppLmYU5uhmJIQe9nSt1KJhGcLv67xl2O1vh0
ws5dpB+QvKTnAfmSiwBKZFzuQfTSqC+WI3347Qce6I3UXTvUV2EMsq59rfA4l42zVEdK2gIPROQI
IkN966XciVcXTTbrCfHmch0dlKTYd2J6AWFmX0IdOXRmXSUqvcWOa51yCC9Zve0C6Zxcwm1EYFl3
8wYXQSp4R5OU/KXge8qV69Gn/vtFCyDBj7xejDKvRoDw9yJaDyaBIAIBmuilPOy705U+CkX9Cv4k
6naqfzoqAmOdTR/esFOlPXYPYKH3X9fkJZKpUDJJTxmknhBA9TGPpBXaFAYVQqJr3egOtobRKLRy
bxEmJB9K6Cy2PDkhjTdK7OjCVa7GD86h294u+JGEgy67XugSH5fS10zulg/o0ZTaZrzgFZ66OwMJ
dEbw/3yDJV/vLI//m06uLuIEaVlWjJB9ieoIxHO0MRwcIEcL5ok54QcgdThFrR9asea+DJvfzJbA
Ht/zy3OvE6RuJBn++nbLenYk9nftX9TQo7bIEKyBC8Kb8vOb3ZPHy8jXctzZUCJU/BIL0XKypGLG
6G8dmu/LpJ/pNdCpuPma7rhPR803de7vjCI2d6Ge8CBt/NTruxLNL1HwrKgH01cMZQ1nw88ehHhc
YUznjGm0q30M+w1zGpJ0HIGBcy6IyPBywvAIav3J7AhH8r7ppz2Ty3bdqGsjqyZ1PnaNPAeu6v4K
NlZFrn0HqSr4jd2l4JNORKzLOj/kaL5wtzpRSoG14Y7Sl3o0ok34ikLb8hs0UdnI0DFQwF47QQCm
ExO4C7mA8IfFiSVM/OBWUwnJvFFK8e2FwMBb5uAUE2Fuzx989zH+2ZnSwGTRlSyuX8PwtWEcU+KR
2fk/vwVX8PRhm+ThmgROfSYDxTRITngDwAHBXfPaKJXrXtTaGbWkjmSVFWIorIIstkx2EpDyR75e
oxc0Nahp5K1NmpdBrfnzX26BUvmdmrMUUQh9rHq8OrEEelbrXGEm6R8/WAT4hLC6ORVxZxExUR2H
Fy/LxPSH8eSUk5sl8ZQQ3RT4wWhUlh/JD57w1mH6hK6li0usdHMEll6azw4HByyjJ8uVej7G4rej
49xsWg8/aBjzCRyR2IOt/PonPSn8bzjpLITtkAQFIRU+qUFCpt6Zh6T8Itm7Z6dKHQC4cvSWOtOg
mHcay3bsca2MMun4+BVveacRE4+YKtuxIkTmlMTzmTQjF31Vuc8eBxZYFFC8zV33MO1x8kzldeRH
HalDSl59aU5TI27LnskrsWoWqEPQawFkl2ACCJCax1+Ij5Me/CFqCfhZg25b316OthZ5lJpn8Fgg
AIXUKDRoIIjQkrsnejxLF1aN5lbksB4bksy0PiSeubOsjB6XatjCQfxhovjfSI3MCxZ6LbBBLHWt
dGxabCRDM6FMrlwLdtlanWzejBsMX/kWcdiyVR5Ezgq3wbBt7Ycp3tn67+Ri6noRJk5VSbTr3GQX
NlC2DbFFAx9znYJ6jyvxkxW5C9q2zXp5fripiys2ITCEdvJtJ76GL8KCYYq1kLNAj1vb3Vj9bTd8
B5ZdTc6bL6NN1FJ2X6figLWfS2OFXAgFcWX3E/Hu2w+hO2IKjFEjByChEFdptb2mAW5Ndtna0XWs
3GhAZm4FL6kMykIriINQxry4WbfsSPGUeus/Musp5hc8oWDPLOK43uPzYZP0K/kGWecX4pzUT72X
quCmw6l7yVq4YjXXfYSY/xvEyTm6h4oggTfQ0jgqXZ4bXjz5OIZxyN+4cfyl5aU1StAchfConCFF
G3bCyDvnPb/WN1RKUKcyqdVb1Z1Th1KotKxmb+EVcSxf9xS+2MXJ5dzyBUijXnjHaL58iY3rRb4p
uIQ2xV/ZfIVS8ZCvltXmb8UWWkq2TIXj4IV1xzea6VbRvC1xgWBS6PD71qSThgfai9N0sA2qKXh0
RSzgCKTkDTy88zyE3DvXafg1kjom70EKkP/O+/yOAgbDxNj7vFLgc9IKfsPU2ebB3Eev09wK3Om8
jpN18aPIvd8ldaqw2CuoBEmLHQw3jbIYkaD/yCb85cWzLKEHJ+d5QSgiBenOKtc4VOd9qixHnuUK
PoNIdGd2LH/kqPl0z6weQcNqKufzqFU5qCukvcg53KN/zmQ2vJ+AM0O6BhqorE99Hk8kkunOFMzY
B/yWdbuiz0QEHod88bo+MMWJdSXdutfhIAT9PqSB11+NeiVaL6wKv/Ms13xfKbu5dlik+mkVjAzb
t54aJQmcxFyOP1BNTaIYSCx82R8sXoC1wwzMugo67LVjRkeG02eRDFZO2ZI+loMPa/M4GotH0XtM
U28XJvQ4cHrv6VRxhLwMGCPChuAYWtPgYzTGrqIg/0qGo7f1k2wkUP2++H3qLx8D74dvxGH34JzI
WAyc6lLJyk8ktlJOJij/F6af4CGm17S63c9ZNX6rPbKsMOuoa35vA4y46zJkm5t8ZJ0/zAOJWVD9
pK0is4K5wbVq48XDdGaQxX04rnVe2Avh/jBX5sg34j/hkuZ2ZKudzKkuzaqeHc5LK2EWOyHD8TsA
ftTgV0CEs8oV6g/Hw2sZf5nCjQilEn9Wwb+DjzuDdfkBIDuDUbWOzfsDlOtcD0zE0i8vOqKL4ECU
/B1ovbbxqrEfH/E4tKEleOsZyJ6pO9uHf95o1G6iQfe/CR5/CL+CI6UyG9vKONaWh+3GQprxU6H9
v/c3lpKBbziVDDM/B5WNJBfLEAKP5Ixo3bs0H4pxRZdmm79+k2XxAlA4AN3qBIhBw9CD1nFcfRrK
C4z5eIx+ZmyDODmPrXUZSQLDaXIofOB4/vNqhx92/Ac2Ko4QixyGZ9/8tBIQQvMXmC22PNfoKSMn
CAbp7PaXVt/eAzAXyjtGt541WbSZvRCS+CypOn069HlV+TQuZSS580iPjfs9Z87a1yoTRpQEUJ1w
qlHC1Yb9nOYAcKDAD1RvYh0HIQHQh/vF/uxlOqjrzJkWlA+r+aPoZgzSevUeKE3A6BESP92641FA
VgBN/YTMCB99AnAre97MGkpF6ixIZ0YD5G5abYbAEka5IOcoXfN8+Af6UMjMyRIBM4uVrPnNJPnx
fcyHpWJPmCIGJlNaMXyE5YDLhNX4N5X6ia3b8gISnurMOZQ/iyLzppQqpHpujYSoL0Q62gSU31E6
iQ2q5MxgB9t+ES8mKmdkF4B6K33FbJKpX0YoMJRJtweYhULPW1FynaHyXrwoqmKCm0hjdQxpmNk7
2ielpylqB46G2IrNEnBPa0Sgs0eLlnMoYrbr1Bv8Ex+cR1eMJgk+bJdjGOmj8EIHii/CcAMQb5T6
eocujg9kgV0pUJ5rzAUa6QA+lBaNZJMn0SoWxlYIRNMybUvYM98E5bznGwwEXh5KOxWlJKN4k8FE
y2a93VoCMEoyyZ5h0KTBe4hGPWYOH9stCx1vimmF2IXjsx+h5gMmUgp+rtmuv+leGVi0bX99KmcJ
r5DCFp7fP0TXoELkf6MR5xwr/eoZJbAeLcjmYqoPtFTedv2CfSGfu4+jNFMAzQiiSfQKw6NX2MGG
Rr5Zzq4C8BGay6x/WMaiXuZT1RN1Jvb5stpq5LhyA07+gBHGhxPCT+XUptOgGtNJvU14Bs9Nun99
ZX4XMalOX2IK24oovl6ZRk1uqseRBhXF0qKC2SHT59xrIGuDlY8nRKuqq3oD70QkHEFQkymYegEo
thNJSpvG3Im7KeO2dxdDDzd7Hih4QKy/R4h9KdPb7znUtws951afSjz+xIbj86O2nQM9VNcWZnlP
VZAIOz2YGogW+KMmjDB7pq6eCYg1R5eo1cdLud4Ntb0UpP52KtBiMkpTFD0QmnNpq3eLmXj4JcBP
eg/oqDkzncSX68rp7/MN98Rp76XF/F4NYq42WmBpQE3lsn3ryJF4Wj/pcYV94QLdsWZnRPHCDu5V
+e9j9QTknQCBjmIrmGA/MacqlWfs//IT5OmSl/e6xAe3za1IGtj/dMWn/IDf8kxxm+4j+Zptv9QE
GWQWe8xeQxbFzeAogH0NKa6WX/QLRZNF2EtqhUyWkpce8OFLgXWYi62DFZCzINSMO+HykQYz0YI2
dobIHdgufHU+IbAwuR2I/zchVIUC14Yl544nL7ZiyWBp+cBJBJ13ad8OzPi2iSJV/IO+1PwYTkln
0yH2IWRnqJTom3d3xTaGXylM6PU+k0NeFDjdk0GMGuBIWnZ/42M1jMAJuw/0rCseBQg/G4VXNsT3
g5MjXAgInC7XKF08+FDE6HKnIwYdwUKIqUIU9WomShrHyvViZ6oqv95JeRs2PzTXA69KhV/G6V2o
ZadJ0KHigb/ITrmkxz10X9/CuxN2uspT0AHUiTGF0UzM25m7+MDrgmJcU3d4QNISw04F8HP1I1HF
TWDqbSw5ZT+ELPi7LIJ56ZFQxfZsGwnASgARvp2Sb+8jznCkJTb/TfPyXv636/0rYlBOwP8MrLaC
wGs0l5ATBsbJW7/0/In8W4JH32CPwzgTXn5tepoKHvY29OktUL8Uvw6o9sBuQA8JdPhocztcz4AC
M9+7602BKYQCm5FZRzRwfVxDOYY9/jHgYzkTBI2k9lRaHW5B/ktKUJn7qceC0ohaL6FzM1bJJ4qt
CbR9a3JofV5CR8dp0CtiZGGeGRSf2/5H89TuJgTF8GbsneLu7+x8g+8rl7aojd5AkN2MlnpSdDQy
5Pn5aKShgyBnRc0teXd5/8NWX/tGDNouATy6XHHabu/tcWp4VfjiTqipS3gtZRQ5WR+/xC0RIPSz
jJ3Gb7bu9w+1ENWCKh5GSinmLjEXqOZO+Drv0RsMFkem72K88r4q/trJX7EgkkZqMSk4s9AFl3oA
hCSUcqZpn5thajxgKZCySMNqSrmURBMfXeKd9W8mivuy4H1my/574ztQWBfWuHrRwFPR81cI/G2g
xIE37pxZCIb/Ji1Ura2XYKyRzJ3x34y3AqAtxXz0nVNjhzbWYRvqlhU2n/Bg9m/KBYwCc18jMe4n
RmFdUlfJNY5IXJi1TJG1fP40qtBuHztB1crkOsNTQek0pG6m9cZb/nDWvfdY8/Ek+VfRNIDuqVCq
Mw8a0GHKOSlQ2OybSmInVoj91Ub+Q2Pml2lx5byHgTgaup+Kgo83/hyFuTKdu1mmvskVtZnxyoUa
bMZZECrhB7Hj5WTwLni9+MhqyRkdeR9vlbusPRRHF9w2E4InJrwlnOahpUF9ZbAUkem91schvQEC
APByJ2L6QcSERU0KmBVgwma9l2V/jI01qtaGNoBU5EnvlP/+ZI1ULILWLsUtNm/UqzEaDCChC4Wu
2tn5pP/mKFYbNgkf09jxaCKjDFlXfsEIxrWrca/yElgtHSM6R0TPwnVU9gyeyHh63ZMC4KcVffTW
uoRhcnvzlvDA6s39cOhn17vqNrqAlx8UDLoafXuWhqYtCyMxvsImktjNO0QMJbegTrkCKq8inupa
KOs+RYUTW0HoABCCo4qDksJGPKkoDvatQdc5IFX3V+ahvEvSlPfH70ESe70W5wZatUwzynNEWvys
pCBdqaS5T5twg4sRgzS/Q8qzTpcb3SIQJ1UHc2rIFkXJRxEGlsJFY5E+pxGcreiJMhFa9gdjHCJ1
kvYFLQxFZCHVuPR7oY05nBg94NfY+GdKYbJTq5BKOGRdg/1Jx+qKTaq0fUGHX2SXZp4Z/s0KKg/W
9gkrR+YUtq9TIyEahY+WBALbdHlR1rQGRGkb9XBukJ1gAbLNsZ0+K+Lpkc0gDwtU/Oq9zpmhkv70
bRLwvZgtNkoN1urBgqA26ai+ckA34sz6SXpSlxMXY9doY3RSBBSZdbGSpHwH9JVO3Pw4flenwNsv
EK2QB5SrhhRWx9YLWz6rymAdNAJtz9Zx6TQpAO1f32LBmWWIcK6zHngJFKc8wjp8PcbKSEGZghpI
veChJuknH1dQ3uFEipilo17itXrbOeFj+bs1nidJUp1xM1nWXLVQ9atIwsQUxcMMLLWEgkKWtqwM
p10phh7DSl17X92d5qca/8wlYyWpUARSKE6cDbAevpngUYc9MmnEalb0qujVE0HTqQfP7VWhT0KB
bMH4o5G2W2k3AGdng3CsDPdhpFk+hM0n1gQsmRoIrVzmgmU9T+RIeaRugMufwE710l21nnm8A7S1
yvYdZapLNqvkkEHxcmMTJKBvyHHiq79RIT2eSPQ49v1pv8mbcmOSUWlck5YlBWOsSmaTQBXcuSbG
SHKHqcKH4tu7Emd8c4lJCU174LvesSm7Sa4kfVqU19tWOw/5wRC6Y+olb/WVmaJHPkk3A82IKRNT
CWvmqk6Fj63+ndYh6wOTlAqW/hCDSs87cOW8MJYH7JvN4eYOZUFZrGlZnKAC/gHhyf1nuXlEPZIq
SQL9vG9SsD60RPJoIj5QWWOsarUS1Q5w5IFd3KgWrFnVVIHD9ZsaYov6Gdo8uE98MH8xuoQ5KieQ
A+dsJeuUBehQ2R7EC8asJA6lva+MWMSkvx5xmsqvgmuhH9Jp/EySPXqulGS4uyuQ5CmzyRkVJyie
78PBllSBpj4oUULI77WBcKQMs7tJhzbaIi8rAOpMQgWKEvhku2oR0VXGMVgi39GTsVF7aK5lbkuf
kq1U39ZUFqzV35uFGZY9l2QuyuN6wsX1aOeAYxc9iI0xAa0NAzbciu+n0QX64pIVXjJWh8i3Az0O
GqgaMcKxez7wh19vcuAv05iljqMyfCysu3mVyd/KCRZQRd/8TK630SvemiSuv/NIAjPZK35jNmD+
ysD2OEm/sqHRymUU575c9trONGp6Eqaz/LxQVDAMO0SLfGfOp/c0uYiaU/IaC/Hc6p1/4Ja7pKeN
zONxCaLJasg4t+K9QxJ2jrYGipdWVsLz/rHHb9XawI76CHWMy6nRFTBaHIglnwTNr9J1a0Jbs+CB
sj4hZ/1KcJJZorREbC13un0oKjSvz+TmM2Fm2jX8HyNZTEeLa+efAms7fYQ8KKdy/Tuv9SAW9wuR
HEeTebx3tbJg8sNjkrEL8a8pGe8nWM9LoLMr998mmPpdeZSxaYX3jNz0WgGTTKFJopGMsdtZLx1T
QD8zmg/9NYOrwwbG7erteNUvLVdyLP2zPaoT+WW75cCsOP2pxfPQlNInhpB+bdVph0T3MIqnKf1X
lLUKHPRpGKBJsajy95NjXIAaI8SOU5KL1Kvw5R3MDBZMMBtJifVfm4f7UH/dB3UB+q87XcttEbU6
Nt3XOt+Fl6u9ouK82OoboUSCRe2zL+/XGHAonwV0dLmeBPYe5s/qhvp8/oTORFitMGdgFhcJE30S
zzdUYUPdt5B2H1MVqOGx5YWThAgdx0e9wepsZXp5a8rv4+/p+qzdlV88bmzM8P6365l/rpYS/u1c
zeAm1NfGZbj8+3Sk9nCdYQNPMqVMoLtYxX8z7cnRbekap2RCr12VcUQr0iZFGeQmzz0aFYret2+I
3F+HK3ZPt6/MFMktr9Vfz8A6Nr2LTo4qiRxNpx0zj92G3xXd4sDVQqKMDZh1eHEYWZ90X6tCiVsu
Wo0ruW63/gMbtROPOYyAOPHNJ6WMtyUFCTZ9Q5gSuLDI4zd1x6dfX9xymutAqFVz0IW2pPLm6KAX
FKq9PcZJNB/lJV0UUTLa3Baw7DDxrRjPQooBI67994xNwJf56ap/IHylFtBmWgrXnMqwmw+f9Bmg
8gt9f1IZwxGD+kmMPSlwND/NpgFJQClAXNnn37basLUyWjqPrbTQFjjR5DtHRc9Fl7eFz9fDbbyS
qIFYCHHgYKx3CyTdefKm+ATrRbFeXcbWECyd2ZTK+qxUbQX8uNMTZ3oeuomQDiHJmF7CczrJEYgC
g5NzjnpLlf0ys0RrGNfEcx2HiYYOEJJZB9riUPpYPtYAmQSOPkNwwnMSCkF8MHhC4W8Ejsps1lV3
GYtFkhIUlHPybvcuvTZ/K/pTNzr9y1DEV0oCLUdhdZRTJS/QH4RrcybOoYJs0ggNBRKHEPw+7aJy
0+HPy4ySfQXjFwDDVcp2RTV7aWPSWShrad0lP2qFYsN1DgLtv7HhlyKaCtbDWCJL/Dgabx8L0Bx+
TtfLsP1GXFeHA/3RT6QQW+lXT+vRId0ZHsEDIXm/z11Vm7xqM98LdM02Ubrt59bK5SBJXzrwYxZ1
u0BdKVWvQeDJ1zdKn7rWX9WqSbfV4Gk1GkZPs4PPMGKnSRUlLUDhALf15Zv30cXOGiHLZptkLkOE
VpInvJAQfCgJd0PssoOJ3Oh9C4SzDsJZq5VsrfIMmjtDTM5yormh2an3vhLjdABdb+SGN6nvZP9/
7SH53CBH/zJ8vTtVQEFkjPqBYRBwY7Bq6eAHkawOsaG+Ja9rVmJ7ng/T2frr7JDb+1xXAKesoLiM
8PESfcs7x2QX5Ijd6BoVIPhpC20SyfDA/zaCBY1RCf1sq/AjznnGmXlPKxP/+Yb33wUKy+Lp5tpp
U9AGH58+3s9AjaAgpiS1C3p27/OHhqJpp7wqRzMPLUj08ge7IAEItYPr/HCs05vU1JSrYxWhWXve
3NufRCdKgc3Lyn2CDYQzGIBVG1H/6G5xq+Smx/e7pcEuVqYdZlsES18VivxsOC1FoQBGx2HjQ5Uf
wDiBnLp/cMb5lmMcGluN8g8pID0b7dW5qvFcqGQyv/NDjc2r8X0Y8jm2t6DMhyMghH8UuLqjrUjb
cFeV2fnpPAtriuGu1X2ltM+aId60hAn5VsnbqJ2XpF49MZyFuiSZb3QDHNPAZouAA99Hj5RHQZH2
FDWLzZa1nAKkGixLmFYM82hFJFG8mh3Fi5sFqXnvZr2pZQdZlpqcp0XgMNR/qWErE+n1paRV4YFa
NKOPEuMc5z3zo0OG5oAGv9w3VFt8IJC/3MojgpVqGOkn/S1YHwWdhlu4cmetsQBJZkMANZUA3CTC
IF6MspUO1VFYBeOzH78UDlqjnilrFQylXA7g6/WN3PAVRO3yVemQOY/f82RDDpHcARWQpfdOp6lv
jNdav7R8Utox7J8Bh7tItGMKHgNaVIIrikLJtJDV7NFW7HwPt1kJqYsuqntQmjLxXiR352/L/EqB
V6htsaqpKDUurtPAxnSLD69l0p6IOd324lUQMm521Pub8WqxuqfSMhxODZ7sInzFH1AKaqf+6hYt
ok1XJ8cWlWxqrF7566JdP/+XpHfM8xnVR/P2H10J65hYn7gHbFwLie1Ej+fWkamRKjcQNWXS7gFY
tuAKO0i7M2rWM8NtbAUg/8ROcCd7hM1u+auBQ5yNbCyYNBAqVU9PsMPse6SdWnPpZ6HzzKoE3uSa
wdSjWGpSnQDk/oADNr0Jef6bmdtdwRWWwMKeK3m8AgHBIzflKrkkwcKT22xkJMb11WvfT85uYUeI
C0qEosOYpcvnNuzotXgfaO+T5zIL6XvqsZUk0h1QjkQfLuVVByKOqQUcP+JtV22ZENfFs4vf1os6
zeQZYfwxipmVzfp3NhyQWIZTww06UasHKjkz4jsIkBglVco5LE3iCp0TQP7Fu+BAzXfjLUeDXVmX
8GjXOj8g0ve5VOm4yzjAr2N/bYYNsb50zHt8PCKxOoTXRIh7ojm4vJlX6Vq1ns4iTihpzC8r1THJ
amsIpQ8z0CeSpVh0IJkrFwsKWPU8TIT6dWDKrBi22Gov7h7atbnXkElciXY6wYg27S/k32FPZDZc
VEooSOGmSw7tc24J6RAOUN4wsJpasZKdjTDgyzLmxz5A0oa3HlMvqwcZXlV3FEw+zz+L5vlZt/3Z
tamobVGrw3ydaRiHGptPl1NRIECXsP1OosizJnpIAJMC+UIP5ekNfq1MO9gQDDkhNT7CBBzMMHDm
W9mlKOi/qMvured/4fzVoOV+D8t/AOyHfruJmEVuLbCwfPyPCmPjjmVTLX5Z3yWbEcdMQNDS8cZR
rCgf4QKNguxQ45pVDnYavv+INFo5bU3xzxxcRREqsLzl/IUjqZTmgku6Pq1ZVO2eBa8KDZaABubP
nn5aaYNR8rpUEgweZ4tLcyjgrIOWDm04Yy/N5/wwtu2BTijDl6cO0kd/4z+YUbvgqcV4N3++zS1D
+CgwblbHMKzO03ZHZIkOD7Q17UZ0J5tPAgKmfPw8P9Ipqc3NHzWRZDT9ajD2EJvNl9sZkntsgZ0l
gvv53jTuqqOJTsFx1NnSw0PgQJh/Wsf/JX16nEZBPrN2lOyUNqGoNdtoCNVCr33lg9CxCnbBAPCO
yiNGFnMZSBz7cv/3bwZ6lqvdUPia+4U7zdvqjg1/fQhPmjtcg83+iXaxTFmxFNrmpo6vl//swDjt
6gkm7T9wKlOaO7xUkurAughnePt0CcJ3fZ5OTFjN42MoTKj2EKxA3eIcGY6VKE5IxI9P3huaHr4a
TDgxJBQGwpp248hxWQicGHXq7uWNSLLMj7w0it/YujS07Y4XZWqtsMqaAZtNX6rsfB5SKvJb61Jk
CSfmD6mkgknoeOu5vVTlguFaReCiCrJFjHlbyDx096h/epYGuA3UoHKfSyj+Pfen/kJXtkcc3rQO
3gvhNS871J7odvDBhqf/Wc3FsmUZtnX3l0MXKRt5foBvLAzH1MQh7fWAx9Jx99qPrtl1pzzEuaX9
59tYb903YHXoBeONemI2rsaw9/9va0AbDOah4XvLvhs4IyZ/uj66maKnsS77/vMpr8G+aY+hnqN7
WP2F5GcMD+Bxm9QPsBJ6sxYkhjIJz3odym+9Ipa5OYmJC47DDV/OcWwY++ROegAg2IeMPJRtqZZS
iKovYs4UEKTA670Tv4ya23DSHpGBvGy48LDTGJKPkp4wYZoIW+ytbZ7p2KIOrV2fAoimMzdIMyeN
N3HL3A89J2ZfgyE0ssE0BNWS753T4yl2m9dj3975aO83HsdXiwuMPnY4D4Edfa89TVJo/gUjtSoQ
9HyYG3Vy/FRzaWpSp3s9ImR4XXtnlllDcu1pHKaE0LlXTPqL9MiXw4pYPXH5X5sWCg9A7fyaPt8G
BZ2cb0g1ZsB4RP5n+zHs/DXFZYb2iYCELYayFe8p8qRESiHi/+GYVNO8D3PyJFab9a74NPkK+LAQ
x2otsv4eveZrRbXuyBxqHMSRUXYtjZXWOKRxeYqnTMfkPFrEGajSVn9L9sLR5n7oSLAN7kpcTVRn
0FSryMc0ALRhZ9HIWZZBdagGYZ+1sM6FDr/13eNVccFAo79gUzCZ0MrBTYmnKhMzHgPLObISzfXu
d0jHhFSR2h3kvJ/nAhBYEX4Q4Qg672oKA9+3GbmKk3cDO+0Ibj9i2oS8LaESykIchsUMjTmoRq/d
Kv0YJ4c77tNo4cw5dNddKKkxQI7jAE2VfrU5tt7cHXfDiBZ240kUBqE7Wyne3kp9hQRarMcMHVIV
abF/huqKZ4dXJQkm4eymCJBT0AD5pS6G80bCF6pFqotiOT2zzDcNuhS5L9H7kNPfaa+3Zt3l+DC0
kb0XkUbw5FZUz/c/hiCYfXMLy7XnJxTw0sC15aQT8q2K1nCD6K+lmc2UKbS7Hl9LMUiY3LRdwU8s
be0W8bhG8xcL3tBWRE2/gVY1E84QdQ+2NlNiwnfYh1t0sdBEduHLUKelPHMMbYs/UfHPXcmY+EjZ
mlVYYf8sTFNLUDVgO11MDEZqcaXktC3iV0MTq6m/Xu4fE1KqUZ5acBcQsxfoQnYCeeQHTVykd0ZM
t+gqcd6yx18l5sQ8ow0K2mwFRj6Ncd2DKsKHo4K2hc902rClIa2+vBst3iLf11cQXWm7oKhcnvMl
YkyyqXfd0639083vQ4Ltrt5Bwx+TuA9j6KJnHm+BAIX5ymHOHJFAYWuFd81iplvtGVzL/E+ermYJ
nVoI9FHugcsWDG/Vn+hs0CgsepYw+c/TbnPCVULYAnbPaHvVwiqwlVh8wS7Tiv8gjY0f7HPIeHUy
Xl4Aa87BBKUiFBGT9ks0TW2vffahcdDQuJf6HHOwtsDmTPvZRONDUvcexrdiQlmvAE43Z5fEu/W5
BCFN6elVP0z1Gptbw3v6mRyjz53Up+gF74L0+pvQz1mdig1EFJQTNZpTGbN75BNjNMCuX6NEUKlu
9S9Ar/nI/usN1wLgaiTR+Vq1WROxx6kZFEOSOA/ZRcW+HND0d7u1wkm8ihQ6il9DSIQJTD4RKYpW
qdsLtzDygJqYbKEgDFE7FzA1j5F36h2zmCnaKjfjsOSYaYeihXYz/m3B8PpFj68tWsXHHedKqJCq
vnf9lT5dc6Yb5RqCoEn5fBLWuRYIIYn96qMPBoqpE7DEQ4ugEH5/ueScxrDG2kqwi8MLVszwthsP
LNx7us7tdl95QETq6247z64nQzzJyWcapxqcUvkeAabzVx8mO4Q0s2r+h7zYI5B8qFNS2MwAAbbt
UXCyCu6BK16GQciAfjXeVu/TzZs8/CoqWug/kuc/9LmDhcNjVozUaMlW4mCGcyYbGr9buCvei4dP
6iB0Lh3ynqmi02upisWW+xIi6E2oGPKBKKFDWdzNsJp/xOC0OPgwJq7Ie60oMpH2GmEHZhcjHXe+
1DTfZ5wvNIcaU/2QLRlmD+OC8o77Yi6roHY6hoswB3d94I1MbF+rEr1YKDEdIjLuyOD5UztEqkJ1
NjNOZSyfQRaXHSlyvHMCg5kAcCoDNORHq0WBzgE2pQztlT+jsjYDnMT07QIdzpPdRhTfqQY6cegL
pg/LthHKRqLleKS5lJ5kGfqeFyzAacF+u0Vt1Kmtm8xVjYCmKerjOd2yuEgrT+/oATXvWU/jbhkk
gHh2ClAdGW17GH+qtbWsgGd5m2BhyPOSubs2SH8+4mL/6yV2Hrru1Avno6FlkGj95MenlenAtn+C
NwVVuNhynjEB+tEm1JtMD5f/eov+1Kevl8wRDAAsIhHnrqJnf0VnZqemXwtiH7ziT3/As5RNhTjt
Fam2LdrQgJ3xAzR+WrHMagYZcTT2/65vohXO1LDTZqEROJurPNZgkSKgw6pRpF3M8RN7kG0lIF89
jm/L3MnyiC073jRRvQpzQ/OBgJ5Zfz+CfxRcCoSsPVQjd40wsMbC+CJ3992mpKUYv1wtpPr9O58o
HsHwZQ/xg3FMtJgZJ2RvAZN353gwTVE+Pde3PYzIO9gN3sOVuD3O3kJkZ11lFjEqkNuclXzfbKc0
L+scVZadB5Uq4RG1eYtYWGpMXiNy5thx1kLnCJUdo7DU4Fp8Uw0FNQaj6pJBC9gjcgxlplC2/3xD
kbIN/NfWbWV/5lJGZElc6NeUUDCPnftg1PzLFg4tgQzgE+BPR+MrjkszVbsqSVqm8S28O6lQddq4
Mhb9avaCldkTFv0JHEQOSgif2aBsN8J6vnJaF9OAHl1eZTPhl1AHHZYY1JCmgU2gcraieYvQZhHz
R+JPxNT9WJ1ZvBDz4Ith2dMS9ZFjIpLVhXExI8jnkGArMwXWPWlSWc+x1CpDaR46kEqYuYPkRTLX
FAz8yQvDb45qqObsCC6o/FpyVYUuuYj+5mEZMMtUcpfLI4YpAMuMUPgRh24CwMeCyydomiTIEqw7
7Y+jkrruwX334uMj4ZhvpEbsvXk9TbYpVFCr8vmJldviYLHBUmUy/WoAF9Qc6sekoOojj7A8vv60
G8QxOw8n9qQm/6Tbh5fIlzq2vfENDZj4CiiDpCtkbRNKQjb0uyspD4X/hM/5AoPJlw6mCQ1N7VBW
rfb7/t5ynFEkJM0z88jQ4gku1fUiYse8kWnvCUlZVhTHaOcs7HcC1E6abeckGClXM3/NTk4X3qG8
pPPza99VoJ3n6oaYukwpV5t+DvTVp8N8r+z8a9DyrNCxZpP87wUGVOFCJQlbSiQa1zJuSPeGDehE
NFMAnReqt7MQ+cw6g7QncizTc6ZadHP10ACFv0ZyTeE9jNiS1jlW66a2FogEkBsOzdxdPP6AD73Y
OZmNnx/dts6PhY6cNBOhW4CyO1H2T7yrmgQDpWKppTfYEsdCH/lkpe3sOHuTPPwWzHyB+tTn3ZzI
ejLp6HTMjtR/EsfBWJea27lklb9qQZBlTa9nliZY3kgRwb+8udAMh/SUsvEQLK0z4bhn8ui6p1mK
f6CI+crrEvPxqIREl3ZO2YMX1tbco0DTnUaSvW21zqi0ua77DCSJ9iFTtmgFo3BAto1TV4oSYMzJ
LgEwevMqAhjpFqUrxKMtoqpxgLcw4M2kgjrOVWoMF9He3SCr/IFAe31nqmsQrLQ/qTpiGgirnbqZ
ZFiVMrTcbDFcge9hNRwDTMOTrU1FCEwjle6Mxc5zz6pY7SvlgY08UOD8VJpBULpoPIOhs5OU3Uyo
SVVKDpo/kmaTDdzuPq96kblwTYicvjuBkk8Sdw/aZ5+a83pOp1UwNjLkGkrqJzmMp545cWTXWPdu
+SszcHtz8taacFb7mzW/l4oLXQu84BYCO4lyNnAK+cxywNVVH5nfE9ToJwXmxSwu/esIqu3x5GHr
grVQAIRg+sKuwJF/Nrod8v83x18G7KaLvwZ8uh2qNfENFTWVWTyc/trfx0n7o8FqRbS9GOxoIgWe
wOcdJ9QKLpdXvpQUZ4QFnt8fDP3xbYmOO6Nstj1o3jZWjO0OxVb47Gw2eEsApG8AMzjpmNxxlaYS
+8RfYmTN7CrEAddohezHyNX3tOOXiFmIga/VBYHYkGV7guhHPiLYIJ/tUB3gM7cndK1Gxhkeb7rh
yfAXjsMOPgvVHf3UDmqvy73zFB3ba8uhTSLnwUBo6Dl9gv/Zwc7G/Wzd5qQtZserosxoSsjFX18a
83hf0IRP4zJqqCblP9/rfWejW0/br0OerHhSeJhu/qpqD5XaTr7bc7tfdN5jtADx2YdCvd8oEkQ4
ydXYX57sunYD4w3l46ze6AKYZ6GdyG+MJjVk9agw/Ku/GlKzy8AF85RPEIy1+qG2ke+rL/VxmlR1
DI300pT/qdRE5XBR2G7OW8IlrCY/zQqy7koxxrTS1CJwK5hGS6AujzwwY47qJq5TrvWBunr+hLdX
Pi2HDfMiJQSnK3GEwdJhxI5qvklqQOPy1+U5hQ1biSKrtLmqKcNXqhwM8eE/KoFOkR43utZf1uI6
3w7wZpIMMncSxBy8CHZwmHijGSZ6WBXzXeFuU7Z8Jq9oC5nrfwgQSS2cQ/jSvybU3kXITTp7HBeJ
5sMSylWfl18J9S+sXXJO0EtcNoMlnfOzHrfZVKlPIDdXIuvXVqjs78lNwzU32RMDJbcnzAFlNU5W
2ad8HtZqIHfd4HlbvjIyqF40iWea1r0tpZkK82YMmR7KgJcAoYbUj65zyqpRfsNIib4w0D4tA5uM
wW3goL7cEu2YOl7ux+50VHLNEzkOkrTaooce4UXpGXpe2gJTOPtjXBRlpdCW6+/7YseHqkOK0wDc
PYqJIwzgVfVkrQ0X509raON9ec8afUvMOATkS3M50Z0HwyyGZ5V5jOi0B5kNd7xBAks72y4adZWW
f/QkzXusHcSxUVq24a3vLKYcQGHEkP1wFrMQtpRhE0KxcRbSgd+BLp2VZPpxpeuhkkVctSZTgNdJ
T9paB6VcAt0XIqzKajbo+4zHjXECvZU4CdssvcyIspeW0b4lJc7iH4Ldxiw9MNRCLNOKrP6KQSzV
A3j3asMJBc5ZIaVCBq+mG44fwWBknBaKlnhgDXe3HFtP7IUNzDTLa5bLdyX130cJfXgiGDNqEXLq
PR//59nBy8IssTHrC2w1tLUbZnfVyT12f1cSmDTpuCkOMN+vV8vonokmyTHqM/ywOHKg4inSw9v2
dooZhc8xEs7ciWVJtd5yz4QzAwqKeulTVmiCkLqVcU8yYsyW+pN4WRN+b1S5V6he6sLGeFoAXQzZ
pcox/yLDm2rsp19m4AoaTV5qWFUCkcjW22dGvhj6hCU8HCTqXZwS4zStTZe6+szwshS0+d8IlFQ9
2/402OrxSQVgErg9lLeOg5xgdU9l+Fqg9dn5LCR6AOV2yruc8eMRkOJcIQjzf5UR/fDJIUoYSa0o
z3b19hBrJi2RrMR450LcCBaZ345tfE1lEFNAwLnCdfacTN9BvtIQPHsSJL1GhYvY6nP9F+S/Mfvm
NYfAsvhxveIGV6x8WlButSa/UDkCpKcsnHu+2iA6bq6aLG2PgIJI2uilS8KMLiOb8w1vraLfakTS
Ly/+jxTydOIVVIjZDSgzIbiq4ALBwNzX/dRctddsEXdjAMe6b9E8yEQozs/rPP8S3wSzIfST7H0i
OWZvPjj/w2DKIWSCJjBZxosWqx7SHw92q9725X9GG/WawC2ok1Bt1BnhdlZWeu7J6eOkVJ+oGEfS
Z0m2YfukC7Ulh+zoJ4LMVMPa3jWaFIhUTE9L+vssChZwf0KwmGHdD3Fa9dtbp/wdF58F/jUx5hIj
6IhOalRQHFtRr9JIndWoPfUI9KFeG/vLsScze1isvNFNZVEY0BjUcNrFbUMMWIrzeodhgBFUC35s
6wa2Ge1BgEfA3pcTM5V5FkyvW8UqY2JGfvVGJNHdT2sXkJffz9hJuOBzmQtsUZOdKMzhbeaLHChn
KcyAyAB5X68PKa8gl5pKBh8C2OUO8JIci6vCU4v1NYrQRXVlpjiiBh6Pa6i22SDIVs9druEOMJrQ
jKm6HqgIe+w3VeVoGVaKtqm867oMM1R88CseWwkcNNXlhq/nTLCt4a/CVwlW+ah6G6Av5W+Dc81V
VSxI1ThurhI4PVfJpUk3FDmcf5E1Nv2hjmaGawgr4nMYz0ZTZHyLsFKKZ2u0zlGy3K03hhfOgs10
4GJR0h7Vmv0gNxVg7FpHiN60krugSieTKHqEnoz5fjR3geQTaMruRyhafeklgpArb0kzCAOQeusf
jwFNiTjgQWNL/xWUn+bAQBpKafh9+ScSFmmSGG0crUr2BY9GTFmFMQ6dfiIxIJcFOtgYG4s6SNit
hDeAT5rQjtCFXZ3lvn486iNIB48JuX8DW20Uxlz3/8i5eew6iG/3fAQjhQejbCjEzbkGt8c0F86S
8OR/zXR6qpcr4Z8nxf/Cq22EQcSK0B6haO+YRwflcQIn11IOZe/7TaCKVtv+zHri0t/wDzFYeeYZ
zB01I8CvpLK5bAfpc3I0YRdBzx6vdxzWU+NziFyzZRJ+2t7Js3C78ulpxu7k3v41Rvmw3TAL+Y4I
pnrT4E1JXKScbEGzyaUdF8+pTbW3pXK8a7z73ckDZz7bxlreDUOok9vaKiH3hjOUt+X0LzyIv60W
YYmtPy8YIbxfjjJ0LLhzgBiG+IeB3m74LJqaKTLiwg4voICo78H0NkiXX9NAHehZtjzG/+a7HTgf
q8AOn1G31AXNvRz4Ba7Tk01TJpXtvbSV6viuux1k04I8cXQ3JQPefTSXaLvRjunGdlFjDdawk4OU
QBlTw5wIMoAV0JUVJsh+mOk+EzC+h91dvo3Y2HB9QfVGyZisBO1WS0B69iAdShL9fHhm00T/LTPH
8gdusqypBODjReExWwiWDdGhi3Pk1Ityt4tr7u8fRf0yfGWtB6l202HCpvDmDhkcRmzO3Ldt4fys
MG4BQ8Le9MQNgxO4qIW4gYNOHpc0FiRyf1+NEjRTg3NY+gl/0AsaVav/eFXWHsy7i4aqfBCz6ZDw
ad/um+F36SBzaE+G4m6WFi86CdbZcgga9KPALDLLmIz5E51Y6glNZzsEJdC+PDJaBVWLstGFMErA
wilkUoR6WVHKys9bIgWbMNuRntJobkRi0IT4xcle7PE/ws2z6XrRuttTPlkcbYl4XmJy/NEh1W7n
k/slE5lazdAAjbvwdEL5TbJaIrNoLyuvt3LlT4lC3oUXZtZEpsxNUzYZWCLkvX+FyMEV+2ZP1wQJ
9J/3qekawr/kyBX5cp3ODOifJfmOkMo+hm8pmYe/JmqDhWdG+MrHDiQRITOOOLaYBG+v2gONVIWU
MDAQAmeced8NyyYSv87uzoFX0gRbQq2Hbw0mf7YTueJBYtDnwyOg4dniwYNK1qjFMrO6koImjIBX
Nf2M4Vat0lizFkF4OaTH6dzJzwsx/v6vkAwDxTJk19j+Bd2F/8soFyhN9mGD234Zgqrg6bDlpmTt
OdC0FPT3S1vzoSm9116m6s4mUCw4LViXcf7s/nwg+sgJ0D/OMsw1ik3OeHZMW3rBdCITG7PQzQeU
j/LxplS/XEAB5E6T6UmX+hllypaZDvIv/khB5TVMKZI6Lj/sfzTNZWfnP2dwxMcqSjRIl13kFUrA
P7WX2Y+3AtxOEH8lcaP/NR7WlCwc6o+mngiVBwhRipEVD4SEJ585ohmOUTky+BBJUvm6ZiaEB8aj
lQqduRMKKH+Zpnw+BIa8LdnVLdS70+qogbj+SwcxII1iSscZKijoHIkVyTSxx/fXnUOc/oc6RZP4
NYW0Xy0mVUpfVu3TbGYixRxb8+O5Bvml7dErJim9ugDyBGfc5ScGNGhbrNrpjHaBrTXZdzCboqFD
yLSZ059mMayeqZCVYcwhASJoLbJdTvkvPHJ1luVuA5fV3EpSoR2v3JN+vUolUGHhAO2Wpyg1SlPQ
1iVntohGMlMXIG8P+dnWzY3dftrExUNd8y9Sa/AetSv8PvbUTWoYiDT/oG+/DcMxYKKUukH8nPjE
Pzl1LP1IHd+FrfKLtovrYeWHG5WyQPtiJNJAkcIInUPa1GyYcA9+gEY9s8dbG2xe+QDwHF8kC6v1
uk3iukNNY3RIlJJuWkZDqL86hfvYgqH8iiNNuK1n5F0pYS3/sIgJsqz/Tk1jK4IlVZwzwYb2wQxm
Ou3T3YCAmaSpO0Yqs4sNcVPGktLeElKiFqOaIulkXQdUoOiw4vNqTQpdic4KhQX+Yq+8aYMVK0B3
OkBthA8y7ljeqSP82ZxfNlKRfDj7kKs7ZeIyF1HRJDJ0388/7SsdJLR4NwLo3A52VqUOIIDcrgQ9
IuZ83qQo/AbsNa4l2CovFANmi2sF1THTdFLAtJHO4FlFoj99HSRVvCHER+EtYzPb3nx1UxAatUED
RZ2N/MnCPljJOBmGceN7M82pj7kLw9rnFZTJfHWXZ+bzkocSI+0oBRmDD8XQVkh1bqVwQbS14ZNW
V61EeUzXeJw9KkZOceDdBOaEn0K7D3+ScHDmIOR/6BfLmrMyW3zk2RzLDVouuqi1/s1balvSQMfG
P4yyIPu8VhghURuqUf6OcteptUu5CPvNXa+pfB+3ERm+WPwKkXp+Su5hD7vazH5mV/62Rm4LaNCk
sSoxIUKqwahV2nlAmdkpLhRFqjSQYmk5w/Y2KRKMQFsRjmfHH8zS2MTVNTFcAYymeaallqtAdXdm
UkctqOALKtkK3Y/O4KMp9t5/k8IM0dZtaLQ/fQLlwyUZpL8oqWlf71dXhtOjb3E+G9bhA7uqNabR
irXDknTlzuZa7xDS0pkh0g0QPrJZR+uHTB93PiJImL1iXgQpg+/E6UumomlXrOpbfCzEkx5DeMUG
ldcKM0vxn7j+EtHbcnDeMXn+4wlPSiO4c86o6Z3YBFG5QHGCcD23ZUflTQRbGBmcrFpYgDA0PpAM
V+ywpZ0txCDW7fe/oLCZyN1J5BPgFiD4uLOtaImQHZXn0UDQCoacpCsPlx/dSrZjNHl4GLWuS4Bd
uWsXUr3xVRnTBHedHh4xwIMDnuQmt7ZK6NYvNWrLVp/GZY4psewTzvsqHI9+Smnm1XJ7+ZQySijW
FmyS0zD2+kOCuZtnavV5oh2UksxjPALONv0PxpXwhnKJDCyDVB1UOdgDNNJtfVEwYfv0IlDzTtRU
NHDm/zr6n+oLLgViF1Y1lwiwpgCy5dNgvoECQ31wEXK1HLbmREzpTR29k5C+P7U1gkHSI0RdxURw
CpcV6dgn0Pg66KvsvCWoBTywTwMYhR9ISMU1xHktIY3lSLaBc0nbgq8eGpKyttWOZ+P81wZIQ1jc
emmXAac/naxJBo0sETQ/gxpPHmGaPNh50UBU3C8CXiRwVNwF388QUhPC0HBw4+ln0XRraQZGy/2n
mKbVY3uIM7SdMpu9iMxBrxHyvEmAHtyqbTMnpByJ12eVKdNGiWIgRqgQDa5CFrXYz5miGojwYQ8j
VeKZrgpuiKq6pZtMlj3mmuNLcrMZB5skDbTUd5Z8DjmAGr6I4WbiEJdfJ8mx3ATmVWtfcRSQnKY8
n1m8g5s/V+QCdW20KCk4dywzXMPvTedkOZQt1XtmhZa+gU7KvDu6ApKNN46IXKc8eklEDXfCdlar
dOE/N4Lg/BAfNtcSdZgcrQWqoGwM6f81ebaNeh3/IOJLHX/n+pnHm8dKe75fkFfTgXNHYFjiv3Ff
WnSU7Plr3DSaGoj/SWA/RpGi6wHMD0Ni0gqcZJ8jjcYbF2C2WKDD03SDLxEGbBoVgOOq0pgGGiGj
IZ7QH4FaKgfiDnYTNi/d9kgCpOlVU+vROD19j7r8tmADSj0niHqDhmUv3H6Dys2Hw4QQ6ZmG3MH0
NdT5Vwtqj4tRBloznQZeLqNjwvYX7AvtrjZTdVCNWnZIb/FhH/uBH43l2e1XTPwTzGkyh2oBILzX
xhFLamGvPr8AEOit+aEekq9Mgp2YCNtltE0fPVcwYMLRyENT88D1/OVcTIsdfqiQtvTNYFmvhpNR
c3W4VKi+UafAh3FNdowSzfPgmdY58SwH+5VHb2HELcgHJa1vEhCA3rfneVTdf2yckiu0MsPtPDPp
uwEnPyQ8SK9MdDoMcWcGIuzpAr2oRaGHeQIVilpqTbesFmd+tZJynDWJkF/vGDtApshdk0hbwhsX
sOI3TdyIQMnA/QKlH9kmjkMfathYvkWEa70K8mZxdu4UaPb7hKmr7ebKNAePK4zoxjDKSWrdODvu
eHgI7Wair/HxgXRf2YA4LGdtw5yW6Fud4zH0pefqIdtldEg06QRRNCqyWzz24+DmpgXVaZFI51sP
kndq/EniekWjUgiy971yHOOQsTYbdeh0CuoLiEeGa/Z/J637rRy1gCG6ox34feaSdPIb1iOLtyrb
rWUcLO7GfosaPoKxICuCsir6FMQg7scb4lCvHWc2Hu3b+0EOhKMfFzRQtT38q6aE4vgIbP7bFswo
cyVcsLIHvEDkGieS0uc9kwTdhS7fH84XmmS4AVUN/wSlGihhIgykIsgemWmFwK18tMruyRKUqOzu
HpwL3uL/8XYYMNhcukJt/5FU92aLQj+c7nsCaDsRzD3XwGPJVrb5D2R/1+mjUGVDzOMXavqnmrFK
bEjpXUK1xGEx0GXL7qw2McsXz276L0Zs+51T6htzP/YrnMOHetMZ7duIptub3NTAQNx1PkMH6B6b
faWMOFRK7TC5MGyKULOpsqwenLoMtWiBfexaObKGkFUF/ErjpLiQTERvM0GsRm+nsciICr22g1Ei
AQnZN6j7hsbbWahfJm9irBndIQqdIM6Q0HGDE3liSGfWRe8RcjOmSMn/h1eZ07hjb0AAPhV6sPWT
g73Etk8q6fkDsXOsEFwfMUmlZ4oCmBr3b7ywCLpnCdnIPEGSKJ1/PomHTv7w2IUqVFd4GD5k3ZBo
/PCaMkb9Hn7uYQCyy0cZ2N+BLCrX3eHovd3frAj/mtRVrmBk3D1LyIn9HuDonVF1u6Q55shEoQ7V
JJQkdZSa/egNLB2gE2pSLYZCfXihSGBKIboXcsl5VRUk29cfkqzh1hwcUa/2DedEDJ17Q9PsuMYH
iFKoztdTHc+t3erPieZGC22+qrJZ9kQoEUdEHO2O5A9BN8HJ2dMfFACgdki1vQH63mZL382vqeWZ
RTH3wLqi9NEpZDbM6cecey6vq1U/NsldfY4Sf/FI4t7xqPmiCel8xbjhXhK97u5Qz7uLCSp2gQ+l
4nzMINQlAcEV+Zasrrh+eu96+kXNqhvJjyhsp0nFv2Kt8GE528Uw/ilCN7Wjtc4LwtlCTx3qXK+F
WJppFg2pAMrwzLCVyr3t256JQE9dhTLcI3tcWkNBDYzjqg870QCtJjFPMx9YJpEusAUF9Sv00Isd
/swElmQTDifoaznMsYvYDq/PfXtnDvF+uRWl7t79xXFUOnn1y276pBxudvggn1KyPBiWVUexeL3i
5Q/Pc0taDlgXMzjJT4UY33O8PKj08eLEs6EVii5FJjVWE/0uyjgziKcZv3R54/Ir9TEXWZyntwSJ
sMZpnS/nlRJZeJWvaIa1qBSImZa0zJoouMSMoA49lAKcgCuWDJDKq1MBp5FA25bdu1BimivEbXTs
/WNYKm6QgfcRk/alh+P4OpN9F6S3PqZgr1io+6J8lWiGFW5x31cSfdHfNSH60yx6iqYf2x/c2ad5
1QJCyxwoeM8Wc3FIEQueBhENh7Q5Txya4IfArL/b4rYLV/u7IQW4Ytm4+/Cd3Esbc4j9wCsacO4R
dMsALxcGBuon7gWrLzGf+0ahC/TstNidIAlWtxcFxMcMILXQsirUmgT/tZ0QqHC0XvNUkgC+W0Sb
pM6tNpkBVk3e/lNvcNmWkUtxIGDRSszxQuUCubMPTnMaZCayKHeOBJ3cKq8pooJGASM3GP7OfpYZ
Kt7DNCjykxUBWSv3Cttk5mEZdrSYhgTfnauXgYsRNkLeDKsBXhzCGq1bWdmFPTIKG916fMQRRSiD
koEXeXGrnPIunjVLZca7EAKYRgR6/7x83MZVy3oEN2DSE2IO8Fq3W9QLQNitpS+y/RMkOq6N9Lw7
Jj2y5sVrcvwgVP2euZATN8KlGIAI59f8kkYvKr7NvHAcLhz7gvTK3/fz0uCc/RouCY40+TaHx9Rj
cRu/X/gQkFwZPMX5gE9jyYeo9eO0tq1ZN2SRtTAmKQ2koKwCFkX5mGCtDrYd6aJtkAYxwD6/QzAz
j9cmuxjWZfOt2GYb673O9OHHjPj6eeQSXMs0zeoVYWrhMtgl8sX99DI2yDtPNL2hzqAWtLYcOpHM
464DRnPAQd/1xiQ0DDSZrU/XPzQ5NFIbxbnCXE+d2KfUp6muakyIQ68c8qdn5QUtXoEkif27vaMu
qjLKnIrJlPYRcUuS6uuD/mtlnE4BGPtrD5eLW4ZT7x4riuPlmNEn/ooE5BH4GWjTFkl3WGLNH9yT
rSsXdENpIYsWNz8iioKdSBPkcsuZH9yv3UVatZlc/WuPDnstgDQ40avt21/QobsY2Nh+lAviMomM
ecrTKm2qRYzcuFRRNODXV0UfxoT0/ph+Gly/Mjuwulf6G/ieCQi8uBRI3sKrUlL6nrqZ4QpHV0fb
PxcS616zGFitO5RMvN9f3DPIlfm3tolefEUG+QwJzaMNH88Zt/64KH6lLOBOQHKq5LpgtyllwjJj
2/PyPhFoy+GzV5/VYHjEBR+m3A8cYE9+tbQGX88TJgGG/vmaMWQOqtKmlCRs6we5mlTOPKaugZ2I
YEM9QnHOTtTnHL+kz2EdoJpifdEokMMArf2mOL+vRzfTvJ+Xz2vhacmZNiFeaL5+/f3QA9fZSDhz
JAOpBNiaPX81dPVKpMRBaqWcam8+LZCF13ivWFRYUXDsErVuEiBdB48cVQckCzaRkr1xnVhszOyV
Iq+Ong7odb1pmu9rIj0/CkLEFQ24uaQrLs4G6aSBwYIR9JST3s5ap65EM6ji8TmctrqCtzpBSC+4
bmz0obbyBT+7et8vWS8/AkQTn0XJqZhQDn4z1Oq4wtTMSfxPYmmiMuA95yTNqcFkofgAQCygbe/r
n9z6AvSIqDmaV6zvYWAzqKUPWETHIXUT4CTj1Th4isWG7w9HtsOie5kD9RxyNSa7js3ypfX13MuO
ETeicR80qyXIBt5uKcw3Or8EMvzQkhblW4dEtUaNYkRZsBRjaWielDARgh0bMPecnaeh/jMnFGn+
eWzdKuHd2DbuTv/bTGSGwkuvM9bBal4NfwJdRVWzuGvJ2txFQNEt+CqrPHMz2HXmNjvGyw0Nsnd7
t3HiLLGoZpnYSHOQwaB05Tb08InFoCKkBqH1uyWyGfYek9vt2XRH92q4ZvXjlNAC9BGNo6E94PTH
6iNY02KULh2/YZfg8YmBF5YHuSgXqte3/C+EoF6wZ1ZgPQCfK9uWacsUdaIsY4HRMsxE7zJf/TYK
aSxBaPKV0uRavukrQoeApu0vs2KWmuNe32eqbxGejm3bKpuf9wOYu/YvmpJc41KmMGWf9IO9o2qF
W9LD45oaO6OWg0ZrT5brGeHJEqHhuhaZrYywU6+NNLepru6R8VfxbBLHdIVOwP9fF5w12QtnHTWN
GTKFaBBaheUFlqJWV2EDq7AThQYlrHMC3++PIsVX6YlcCmh4uyiAH+p4OJqu3a/4GSSudnn4ILq0
Gnzd/zrHK7ewcCuZqm6HU9o4EOpr31fJLh1C0RtfUCwPXnHERp9YeXOT2ip0C6660r/RQWARGDmX
rKLwVJDtFJvl5T3AQL/V9T0g76E92r16lprKK5U2Fo5qYdAQknw3fHanYn2uP20NcdZSU8kezns4
QShRYwmsHrJlYEKueDVQE3MXJztiD5KW/Fk+Hfj45BxTl07hjuMSkWrwA0oZLThCEEAc/GaRA4J6
cjKECfuBxAvpP47rHRNT4wbJSLiLExyn2NvLtkG29Tc8Ds7XEMqJmGLzSUnk4ZRw3XrjbS/c6EgR
wj4P+DpGrEc7T13wQW7iIaH14JUwOFNEY2zqrP0GaOUD6tWalK8iSfcKEdN73ju65m30ofYgETm9
s5Zr7mcgpTqiFPXzQ1cxISxEwnHLWrSK7vbpyNTCzx9B9f3dBEt+0IkZ8eNy58e9ZoR2l0ADuSuL
sK63JJWasRJxMFwMGNuoySuoXC1v2aML16lRt+NRZXlONcWMYIWKtiSSqyHXQcfksoFKmXWKSRRM
WRtvrsQWMR1xin+bWkLZe6zqrOjTv32DTaTz+l9cbwmRXPDCWrySZX+VK9hsxWTfu4jx1uB9d3bn
odTEnV3MHD3OayAkzZsO2HjkOIa3JNUHX45T9RMTH2hz4zFzeWL84JPcL2D/499do3Vv4HpLGiY+
BkQ+bwPEBii2TqfjO/qESd0oMKh2cv73b5f1ueJZUVBXGq/V60/eXSCSJgCmV5DZU8Z8rrjDd9lz
JyF51KXfd+ubemvOJJxwaNEeJqbDbmiAm48aX1bhd52FS4dNVqD8eEzaFRkOk5DqYA916v071FGo
ZQb+/KA3+xPeAeGgXq9BIib4HJgRWCj3BaGfTyFmWNSvdENSgjSwHZjWEjmV0SdN7FLmbNOtgRlG
paijve16nCyjV9AjEwVMn3O8d+yJjNzKz+rj8hVWIT4afBk2AhfOZkgLMWd4z1Jz0gX7b6l+D6uc
+Yw8ypzIu8gQG1v7TTE2Jrs36A8BRA7FHiinoV3mqdJmKjb2qdTeU4bOdO5Adh2dhfZn6fS5Gohz
LPcE6gkEpbJ9dMaRQJM0DQf11O201xNiLMmTYfq+svc0adcKVajM7APQcCx2Z9wQgC+l//d/oOzv
R3yOyzx5vRzna4YJNrRhhnjXvIps6W1N3tR2DMq0aqbtCFweANYa0C2lQ4+KECV13LND/7pOxxEm
zXqeKI4shIpYNCM4u0xig9VCyxvcYjj9A4F+iVP+0H1WxS1RfCYHhgJ1YbjBT3M0GsN4pCEIKTfp
9qpPH/XyYBjDk9trsgsCzJC3IzKAEiI7guNbmLO9DHkYQinkOpxgF7MvJBRRKHwyqeQvpRqc6R0p
zpgTLhLdxvO4UeUYVRw9LImLWQ7xVwnKEBmWsZPuiKW64y86i4mFsS1f72Xe0FI3iSXUINWa7PGz
94VnDeeoO1IPZTe9YCWAqldeUOymZuabg+qVgyt45ktyEPY2Yqxj2pMMZoU7vP+5PeKQQ0A7T4GB
yyl/JlrflqlMIz9oonteqyIICvFj+893UN/5aQ4Pyuxq+2FQCtPLzQu/iv54n+Jzw+ss7iWKaTdI
I6BmJPG/VYCCLYHWl/Qio73mgbEqfQ2tGhVFE8gZ4wu69JslN1VlX7mvpZwczNv2rxwdeLhTRqfi
yvCNIcd7kzf+YAVZlS+1iYYkMaC8Mv5672yadOczmPFMJMnIawJBrcV44skzQmR6xhjFsijjNePs
muAer4HnGLY1syOZ/6BKd4rzomhZ1jwjNCVTbskpPKBMCBc3JWrAwiLmOEpfBecRSEbEJJ1WGJ/l
70AQ/XgexVbsFwNdL6mBm1jdpRQdphxHE3lXQGMi/UEC7iTrP9T/iJAPwqgMLWwqux71cy7l+ezQ
tjwqCnTi1nyKLE/LGazYdb8uyMWbLwuKjKdGkgLII5HiwDwwxT0tmMJIcPQgySV1k4tIXRG9OoPV
2yj9KIFUcmYMgq3Y0E5V+TDAKn+eoJzmpbrrDI6Uxk2scL3Q5sF6gw9YV23uX+zP55y9BrIr0CiV
uObey8PGjSW50MPQ8Oh0P0/olM/um+V58noHUzdoSURwHyI6znGYa2UsLoYu7HxNqaLmt7tqIZOG
lsEd+uq0Y5mLqUAiXRs9ktCTCSi44+Ru2wK5K4kMOwdV72OrYfNnbfDJV7KoNQovpgsuIADZPXB5
sHX6zQx8DSSFtozPt6eVXP/+JK3IqIxMCLE4SW1BHz+I00KJO6pCzCXQMJsUw+hq81lLprNw0F01
8x0BEpR2W3VRaxUqSmfj3bAzi7QJPXzarawfnR2ut95PSiLtjvommtqr4sLZ1Mu+4bfeVy8kg4+5
nuPnSNTEZeq6QqqFL0J94hgA3faC256lZEK+/ZwPYQcrp42e6RUDahbjeNP0vo5lrFC/M6AwJ76w
fAxF1zT7Ya3yAq/SHsDYZ0qp/KaYBGG+qbzELnUAllCFLMBSuzDGN2nWLn8mIJ3fiHccl0VX5YSo
NnQ/v19AaxX81odn5Xig26gZAB7lCsyofXWI0Kn9e/kXdAOgLebo03XJxjtTA4nvqoD4nqjFizdY
vwC1BHGUWIw7bPddmTXN6bYItHR1h60NSsPDNreMbztUmVGxEBor6W771iJBlunxObKPGy0wSPK/
WQhyCbQnR3kcx0RzR8DEQypoP5sGlPJ6yRNl/A+2DTzSKo2uLY5BM7emS8ABzw0O8748ccHF9xSe
XxIlZ9EIAUXi4sTislNTSDWgEHVMGkbHGYy/TRaELd78tKVvFyqZpvvDcOP96FOpiC3XUAX3UL+t
a1jvlZPKhRk1KftBYjU5KDnZeGj8XHX011cSDMrK+GnSGLSR2j910OTrkuEI1YHwxR93jPegvrF3
vw0xc/6EcbDNXky08s9Lbwsp0qxa/liUz5yTzzKk+j/qm7XSrT16jI8H1U++Yg5y8/9lxL70fryE
LGUcpeqd87+kqTwMw8kNCT7CVzMbUqmso/EXw9fUOw6maYCC9JqCPngO9YpDcm4cl27VnMjlbFSF
7t6GZjl3KE/Bnep9Q2w1cqJLoSgJdc9Kt7B8PrHlcFxQeQwPYbZbdFzLCXcSRjldWY/wwCVfbAiY
oGcOl6K9MAFJz2+glACfBkbM8PcZt6Wrsk0IuWX1l1x+Puu65sELxPiFnszldPP/Ttb+LJgEqWII
HtcO3Q0sIlVBin5XbZXjDkakqE9rAqTecpIKZ3Q31Eq67KBPsxivMwxfhZFDA0Jsy81+qr3AcKMA
e6AfsCXXNrkbB4HK38Sgl4mHr4hewfU1rNpHR/g1ABDM+V0oNjWZU44u6oA2mgkXt3C4jJWDJ1Ky
/1/5IcfP+EjNZMH0eTPMxTY09vH2M1avQdJI1penyxsHXH2V9GT7HAoy7gp+xkBXwnoGIRR0JwRO
itVARqAJIAjuc5e3MYhfBubyFjSeszkQ/HpuGaKOZJqQNuEJ0eHUAJFXOJFzj4hMhhEFuabA4d/c
YGRRbUi0NVjTy8WZuUy2vm0r+USRhCFLhAamo6nK5ZHtkd52Fx7cv0yYFm5t90fgVe7+bckP34Xl
4EXvCLcB0F1+7ItRC5+D6Wxo5VvzuGjgQLhyefQUmgMjYPoFtYLZLLdYS7erczoLHVJ7nDPiKf3A
oS/X/UGBt139Lua/AbqsmwxnbYTtBcI5L+32ZnF5XzPVteFpRhREQB6UphU1IIoaSfXhoWGzPoLZ
6Pzi06DgJpwMxP/HRebIaiogqLYnGMxvND2jTcQE75BUKASEPkdhb+RoKkX83+Eez2dtLVbbLrW7
DEev8RImFBVvZNMorGBruWu+Lc7Y5q5c67pLT4u463eoLX5OX4U0e5fpVUmajuLtke3mgPh/Ri1Y
WK0L5tjjBJIz0Jf3knZcTfFhhCpPQyJyPQ6wbA1TNh/j/l5FLtO94WLvrCI6//RMi78giXI3+UCw
QX1PREeQNBv2sc2t9OLQLOhQivNp/MCTcWIZp4GsJ6zeF5wyGMbXzgaZ9e4fL/8Od1akngRweSRV
xZ9FzA+UXM/7ZuuTCakqlv3G0Ctxd2M0mBK/XxY0OWoQJtroJ42ULfRx2jk8BihNxSGYJJu762eo
ClD/fZcJTAxGny4ojO2qxVROsEoNdIsDaycbRqTIi06F6hMX6D5x4g7bpl5+BIR+eAGoTWl4Jxsw
/g8hPP3n4em2W4eVJBY4b2YrAshr4tmYPlr5NBxpWeMtFvgTizz9F6kUi13kBsKZ5Db6pforjVf1
Nm9ZOWvxSOxsvu3yzQwMEKfhY0DHPKJJPKaLOefjO4fVoLvnUrl7eVJhEkRI8SEn10y1Os+oOj2y
SaJFCaftt15VRrPiEgiiFinf4erGa3UZ4h0Ric1OLtLNddjvDLl8+YuJXlh7I+BfzPgWSQiMLKEh
3ESMVqaV8sGYQIw5AUSffaJFOtwWE4vAJx3xNNSkMxaAma/KXsu9AqqfaHQZz7HCGUCgz1KMOmC8
/ePdKkIawxo0qAZJEkothaTFPzKLNJ0YhieXA5FS9hLNgvh/2krf2IldasFkYneqCF7ZxHn0m8TU
S69HB25Y/FuQ+EefFBqLeUHYDj3SUrc92XUs9uEcC0IsPXxVhswKO1nuT7Rjip9TkDCVAJkcGJFW
U6mQD2MfSX1Z1fxwHovuGEHYl36D6q1s4SweQ+uRlnoqb3sZ4wiSMojWCrpxDr3sGJpZu11ZlBFp
Utsx/PJMvLauzBGzkbbVmj2LKm/vz244vuCuhwcqaYsMBy3N6ZAQXfsRGP5Vncu3Fgqz54yZfwDp
D13PZTHqAi1RHSkd0y2lLYwLWagf0H4H9N4ntW5xDpbXeTlfVBpfDf43H0Nf3RqHxgAkHqWGYsir
ARqc8Dz9cqMK7h8sw+I1CFRpquM0KEWb+5uplxeqKjU+k2KtQifxJkOBnH9Qqfcu2957KkTFfNVZ
0Zgm+o0euFsdx9DXgXalIdzjNvvb0P+xKs2jrRHcRcywICv1t/XMaij5wYylh2O8d6BnLLB5xVCI
kWs28Z2O8+LLHwWtHnF/aJTWszPiJr9R3Lr3g3OW6R2AgsmXshHWi2U7Ffmd6xGI+g1/mKmFxy1s
VwHGKOOR2mCVnmzagon4YwuzYEZfksUWqF3aCHlXo6jNblkjnLgGx/HB+GX6HqEf9YZQC7LF104P
e6xAnAYx8jnisAXGfcAnRPuFQrxo+K2UNXuPAO1FrncuSGPQsO1yj6f2YjkRXecVVzRBWoDyg8p8
NsBDlV768vZfs/CijMinIIyKY0FRTMGh7TPl4joXqSa2o0X+NSs8xiakz7GnpJgH1iyDKQTsu4kQ
NFDsuKHFac+XohM7b4lWqy4HkIDQ+CoKRZwK672HFFb2aYeKvOvyz9uCzz9NlVNpdK3HlK2E3P+j
1LqT2LUmxgEzB0LxLXfZL3VWo3c/VmdFzGAsUe1YQUoSFaf31ogL+yq7jy9ckF2rIBE66wNWRf3t
083HBjh5KcOIt3C4lCSxFv6aUhwkcQBRUC+Sm0rGyodlufcex1ntbbTs8SJfS5nIQSVNq8zdqc4M
yrmNqwivgmanZgFWHGN3i151qrHCY8CVHGg3uN1wn0/iNEx0d+Iy65WFFWWOgLZ5NQw9KxyLiAnI
Y4dwmPCokUvm+afXoqcNYONuFSX7EpyIM008IGf66XhrXwfhZ9YgbPaVplq9sw50BmQbjpATsR7A
KIPuTQcrc0hX0HMsMNu8DCfZWB3sYLGB6VRwTBThj29sGdMJBFbtVUZLmXeEK7jlBT6UpgESwJd7
iWs/uajQOn9vr1eRQlfU1QJahB/Q+pQ+4xWDB9jWE3ELXvIECIx1v3DWKb9TiXad1tb8p0TKlttu
dnxNg3Kzbl6ey7rYej14d2KoFCyiu3fv0IPP8WALCiqZWUtgr/O012XosVZMH/bdSbnADC1W7eXt
IYByQ2PepRcKpNuJac4HLR8eLEG/7+ItWEEMp9RjD9XqgiCbY3AXJK9nfcpMVZ0UCrJaDyVOI05X
50Uy7M4NuU+2iUne7Be5Nemvq7Z8TlucRu9qnmILFT0mEI31kJnCpLyg+Y3p2/8/hqnyiWT2CxO2
cjI9QVlbX23Pdyb2oFNe1nfdaJs0p4WQszyjsuCqCO1YWIWJjjY1OTt5FPhc5yrVxitOndWar1/U
2It/kYtLeSQViu7MXIIJN/L4dSNZsOeR8iZxSBFTdH8Zni3a4/mZLCStFcLn4Nf5+mNh0O4JwwCP
wRixtf1fYQIYnNg2MmT+MV/hgHn/80icfu8c3kJCw3hcIAWuLQWSE+hjK9rRGOg/aeD5Pev7d8/0
ZLvwES+CHIRZXm00KN4Obh6M+e9QIR47x1T80qHYr2tmDe6hV6vks+x9Md/sehyfP6Io1AA1KGw3
rehmfUcUoG/pLfmd3MhMZhy39gdEIIJhVRMNcxOVv2iufW7zA6Yv00a/XSbI7YSrEkZGT/m2fvJu
tdRR0bBaCxVX3VcTuQZs+m0i8KJRtlGqz8b7nhIFyoe9TEopLeMtisTccXYcmdLAF2vZ/DoZBLtQ
iq6PePlOf1ClXynixLQKIhokdqHhJfO0mmjxgh6SX+nBL/+j17W8n0ePbqSClqJvDDKSdorF9jOn
gnwL7B2S1JiK5co+dNAHI4yuYbO2jGK6eAMjXei65KAVl/WOdHRZvr2zsQAbHecVdVGrMhEDBHWs
r3JQGdvTlTFA2M5tU4iKL3X4k+qT/CwsRykuCqVlKTsNmSHW0wwcWcXJEFyGws/bZBSjcW5Gu2X3
mealnEDnhiNFWEu+wtTi5J/pFf+gu155sAqMYZ3PdGBJew36F/AluO2M8heBzasAv/tJpQWzD13Z
2SEdiibq92LpqfqGgZ9/wuaeQMzsNcNzBFYf54FQ+HXwz3GoYxlbvjtt35uGKFjhC5jkUOLDENUn
fUIz23n/HXQ1GoBWD1mH6Vxtu5gFi6XdDq+pTBfBun7tyTUF2OCnnFEjvfxBkJgJPjvc/ouGb5Jw
M283aD3V7IYXsY50L7vUWwmDYqiaiGK2AUhHus6wQ+FOWxW//xsPUdorn+4YrexqEzUABDo57qsT
QdsCgh2UDGRrq+SbIyJS3uJ+oJOUoK16Ilgpg5zLMg74w1Q56gtfzifzsEGbfJFboCbWpEbV04OY
Us9bDa82AXywi917lvhmR5n3NNfMASPvpeYqLrTqYdaHRUz1FppKb9CIDBtr/Rh5h1wAgzIi8hez
+2/NoY4VACb5PZ63j7Quxr2G8yi+614M6Y3TA75SMWk/CI7Nz4gkzFIYWdrFL/kkT3subTGJas2h
5Rlbh4KP2pw5Dq3+lDrGm08c5l8JScJdGdjbhQNZzJParDzwsXvy+rSJcZw2ZHOKnmAlAvtCHQIx
le26f+m/bVAtPmkmgB+PvVBLX00z1nACdYBlxKIMEkGdD/7RAH7nUqR6Wis89U40ynA+yWpTiMcs
P1ncqhYzlxfhVhGtjJX6vQWUbco48EHOkE88TRUVoefmG6lC7yaDquBm3Da/qXcJcQEcw4OCSs+a
a0dSqYud59BRNWU8HZJwxR8Xpmh7WolUjAa9BFBls8J5zGGUPyJqkanXf6rmaj/cX6ejSu0Ht8dd
gnI45azjYNiZjhPrypLq44SJ66fNdQzYX1Tsbp1EG8BUUamwOdA5F9ogHV+FFIVePbAW9VcpLMDo
9g9Vsmlg4X8roAP3XCU/8o3lFblpPwCG3wNVkNz55Kx8wnwGk7RnSza5b48Yy556iWd/fc3N0X1i
Zvf7vqRfFF34LpimTtg6WmEJMq4nUi0IIscaKUFyQZgkVYqHyFiB3NK+lKDAgCv6BkUdJaFflQJE
lbq+yL9/Ly3SDPbIHL0WbJT6Z7cP30ABBwkJWMcAa7bsu+KXPNj/wmn5SJjnJbbDKJ/TaNw2FzpV
22C5m0atLR5f7KDX3c3WrZE3XUTFRVjKuTB3p1qyLgVmdtv8gsGuRAsTLbUq2QCJ70t3/7/z7e4E
hc5V9ZmqoIATIdk54SMO3zx3teuKX6XeyaPJ9qSZJvN7Rh3hKwqkRqX3817lB5QYDKuLAQ5ADG1L
9oJUuMKrEg0sQRvOz/QR5Qh2ZX4C+Zcf6QFi10Gqj3tqtpiFOVQTEm8dSbuB0qQNY5mLUinV0jaU
rh7tBsDxK91i7fdQkdY/Plij4Flgd+Egt+4XnhEf05yCMxp+tOMzawSVFtJ8vOeg0rJiYvSjX9SA
8Om92atdqiLBNat8VIwaIDwxVpdONPlKI1LO2Jd5mzGwgfUIpKKk2CGJE/nYggAdJRKiYalXHuXm
B0+IJP9qE1xu9OBj1kPq40grXfDbpTsngokOfp4Nu+YRZQj8PFVaYPrqih3dJWOmlf89hTojXfNf
PtFXIHMf6rucNWsQ0AM7ZHFoqHOx64Q7GJjvUsOzGGTze5wDVD5TJVa2V8T6mTrSt8pZ0p05L9af
KVA6/sSK8uz17F4asAsxdfex+5O7i+yWHZ2DhL92D6+UxXznfc1V09+9duA0Q7E8e6Jc4yzA5zOG
N73HPC1eijr+zrIw1Y0l0cRnmEJHd2R9bcXQiob/1FuBXd9A3IkF0I6cxbV2uQ53lk5mqNGkFBqF
NcaYT9CCUi7PVNnaXgkaAAPHNhPBBwVOF8bcXqSB26+wZBHxBy04Xych6m1a49hejDUfpLxODTv6
tIIGeWoxAVJQzBqaG7ZrACyMi2f0wH18a9MsLWrTygVxH4+3A04MMmtbnm7+qmPd1tjhgnrJri+4
OZnmBO1LIMlCiaN732FEPDm31T4JOWLYep8fvZvoh63E6YiPhwW7iUNZeOFcXNOF3lYsF6dL7ylz
04mHqGVJbUmv2kGSPqhSkWyIV3gPN8c/M/ZQDpGVO6z0mNRLfpRaScbj4jspNcFVKaz4wpt6/ZUo
0hh+LMV1s3Y2VFQDIqAvj6CaelEVS9wS5SyI0DT57ustXwvL1yqVGT2SWhKImVqQ7VfpRuvaKrIi
/uQnImpTXvnHiyFkbfIQXZzPhlKKK4Q6Qy6vyzwkRgKwN69o+PdHrXmw/3EuODbXAhHMwulzhq3C
mc+pwanDqCPJNW6B8uJWCkGAtRzMnk3L3yxTEQADujB1y1/KS0M4Vs325OyiBAEQMzjvOHZniwf5
pawCTDHyUY26y1NrwafA++PjQVnxcUQSAw8Zd8hM/2zNsvm8k52pVSaNtgqPQ7Wkxk8Rf7CzDLrj
t7GOY+Fbtz39qEOXIy5L898bzsg/3gTg90wEm7Lr6t7ZC74C6qFj/ehsvPAaeLjr5j+z7AOacFW0
IFOxCQ1dWVdpnkeD1SQ+LDS9b9rk6WvOI2U1+zt9MbJ4hmd8s5g2bEImTuGwD+qnD7bNg+ZXtnWL
GOOIIAsItpGTuJNiNw79vsCoUny8VHxg45mM0XrI78qdBC/wO3gKt0xQBY3x31XryJqfZGqyUAA7
jE5ogowLoPh2zEviu5Wa6LbzroHunV5ak7E8h/UxUUllBK0EbMvRLiZOsXJ2pfXvk524gxIWsUQR
yhUy8MUVcndnd5AoSBGpNACWy1O1LNmQiCw0iqDk+V+vx+EiFIL45/M9WsfKESli+eUASZx2nolD
elArv2BosOvEKBhyq9/RSXZdf/B8BiSM/6Fbq5LLzPyfvlFlOrTxki5NxQm5rfkrm2bv66eMGPao
dtBilKOHmlM3GSGNNhqXRGzrkPnJ0qnHOs6+h2qaVqIJYuqpOZmZf1cjHptGkpEGhpiNGTdyABI8
blA6aC56Z7w2+UnCs4SSCDWOE7NzsiddLCN0riqgMjFIVxBy+DdpzIodkmgxpbVCD7hjkMXdHUpl
RVOeSXHfpUS6BQVE0B91XVPsbJ9t1xwDjheE4VMw5eIieygDIYIVS6KHChaw482FmK9k1Aw7FxQG
bQj0FGAVD/xPAlyIgBbU/HVbdjNYWowjS9isMyc=
`protect end_protected
