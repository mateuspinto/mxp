��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���բ˄Ɗ%D���+5�p��w�A�v" ����ģ��y?���]����o=cGnR�pˤ�=V[0�����$d�J;ْˣ��in���ʤ�R�ͥ��+'�������{�X���4�:����ۍ��3g���w�s6Ҕ��5���6�U]���3�pf�h�w���ٞ���	��u!�j�*�r���ja4���L���퉥��쌡ji&�v}�VK<�^�N����[�PԮDL���ߞL_�D�_�E{#�/++�
��ȼ 5�t'4 ku����7��8Z�|��G��{���!늯��G�լ�L���*N��@HaI��$a�S�������g���L�c�?W��e�$lk+����#G�_j*+�mb|� ���((��=���'/�%R�N"�5K�I��0�P[�vDN�v&nW.������A fm��!��ځ�*���W�.����[/<4��7x���)�4���3�Ҹ�#GI���3���	�V;��%�-'	[<;���w��t�	q�L�_��biJ�'��d�v��\���{&���nq~���EP�B@��(Tò��̔��{(�S�s�Ud=h�~}}�vQz~�$6*"����X�1��g�L�k��L��ٺD��*�cD�����O��^Ru� ��8&�'�k�@�0��A�:�v�Y�Z0u�)d�l���L�Y@��#�c��
k��F��I�v���^�`�ى�$��1M4�7G��
������/�k��w�d矄=����]O��P��tb��f\��G���k�!�������$'%�ӵQ�
T�ºo�}��j�j� F
�)q�����CB&�
�V|�!8��+�Bf�3.��J��
ծ�t/�c�^5>�¦����I0�{$��s0N�[��E���P�F���)�#t33`����� ������Y?L𽶀Vڲ�J�3I
O^�cs��`ux���$$��T��ҳc�����o��K���@�&lwOB��e��]u�u"&l�� M�&���n�,@>���a�+(�B��Y���}���Zї1JC��I�R1&Y����w�w
&�p�>$�UPd�|Q��!JJ��� ���@jaHFS����eS��%�\g!�8)��=������>(�%$q����`��6=K��u6�[�6��pϘ>'�a�O���_;���e/���h�0kh��,/a����G���Xyn,�e���V)��`8��;��]�UN>��y#ݑ�q�ˆ/7p�\������CUY��۲��d��吔�D��1�B�}��jk��׶,\$%M��D��@5�3]�L4^�"W�<v��C1|�~�0�M���쿱b��鲳�3g�"egрUO%᡼�h�@�y�j���;���me"���S��IJ�?�p�I�0��Q{d��8y�@/΋�a[ڙѽY�ʑ�	����6w�mK.�7����jL�'�dγfU1U��>��r⅐aQ$������[�,�m��@���mV�����w�����Vb�>�<fa�ϙ�^ ��%`e� w/	��r�� �:s"�%��t�ʅk�GH��kjgY����rG0�N���¡@�EV���Ո��ۻn�\ӛM��m'�4�Vܧ�Uk�kӭ�����^�ʭ��և���d.2}vMq���ı��,>ɽ��~�(����IS�	��clK��ҳ'�$t?�Y�r����|�k#�F�)$�I��se�q��U_�=f|	�{$�v*�%�-ZL� �
��f�/qL�=?�9��fQ�.���2��eT� �u'M.��������R��9������KʴV�:6�;�/��[Le�r��c=i ���Q�L]�?l �ph���aZT���#�7N�c�=&�H9PFH�T�]4���!C��s�io{��p�r-�u7~�4�R����7��y_;Lը�:q�~H�񩤈���E�G�B�~&���#W�rҬ�9v���<� �	Û��ŝ�M���0���'mNd�!�?��>�6�.��p*��O8EQl�}��ж�l���yFPh���Iߢ����q8�}����u|'�tV^��h���V��X��h���{�X�k[�(��WO�92Y�Ṭ��)4~,���	�ʕG/�R"�W��_�����(T�`���0(��&�Qc��Ŏ�����3u��d��Q�#.������5惡��Θ^��\���	z��:qa�b�3���l���B���Mc��K��?D	��G��|����H���r��62QCzg���7Y4>�3�Bߚ��9i�9 ��N�	� �/�f#|��8X(��鹣]����l��.)J��-_���亳��B��VDK��j��]�2��Q�*������6
K��͖�WA�@�)`��<�ռ�(�%n���uJzRS;}�Ŧ-~���Ƣ<�Qg��VU�
�/���=�pہw
\>��&ܘ��ЪX����b�K8�-8r��#�4��R_�-������7��NU֗2ZR�_��[ǜ4�� �EUG����R։dƔ��HU���'�O<k(��-?�����G���,ZzGh�t{Z�q����0�:h~8q�t���)Edк�P��;�'؃^:��nݾ�2�q24�9���3��:=�H����IlEW���j��R���E�Bpw����N��F�S����ri�L�
�����b���V8aӑ� ����*H�p�K)�ԩ���o�W�:-.�ʙ�ݍ���JRQ�!�h��@��W��/(1�����uM���D���\P��5��N��Z���a5[M3p��Q�t:m������B�f���Bj��'?W�;FxST�T�+�s"Mf���޸:��q,��x�o�I�M�D[�~�h�Rn�~�z�(?�G��pUq�b���l��4�&��L9��/���>�� s5b��MM� f�b����e!_�U���)�Sv�;O����&�?������`�^_��ܷ��$%����Ӣ>�W��B�y��/�m�=!�&]�BH�af�Ja�ѨӤ��GVW��<;0͟s|�>]�ZY�w{�ҍ��ޝj0��^�B#4�*LS{V�hJ�k���>$��d�H���8�{�)j?p��b�~��N
��c�|���:Nwh/��ޮ���V�o�Fq(Q�����i੸��7Dk�	����4R�۬�+H�у�g��}J�hm_\����E��{���	o,�(Z
ֲ3ky@�;�;ϊ->���Y�kxG	j�n� �Ｂ\����n��'Nׂ�"���Ȩ'Y��!�΍gۈ/��1��i �!]B�i5�l3׀0�I%vԹ�)[���܃�hx�~�A˥}#�Y]��m�%Eg���3�&o`������?XLT�Aف��׻"6�c�-6|Q�Zn/�66�ȳ�.���,Ό�~b���cҲ�]J�˒�C>g��D7Z�bڢ���L����EN]5jkN�����ugi~g8���{��.�W*�uJ3�Jb�)liNkl:Q�3!p�����(~|���a�;�M���k���ڸ�4Ji	}�i}�T�Sϣz�U�0�V�M2�F����6v��RT��!��cuH�XلՈf,�2I$9�W8��e�|�7O]�EGeF���<��Ρ%l�-�,�8��;�<���漩�[���,:��ٹ��8Ŋ�L��>\d����m��2i�6����O�z�ed��Z���/h3@ghp
d�dO��#!K�ɇ��G����Ʒ@	;l�ڤ!��K�N;��_�b�������[zU�4� ���%�F�^_�N�S>Q9v�� v_"��΀��9�eDHvN��4�:��~�[��� bNK7�ﻁ��<w�L�+���A�l͹NvzmR���p��ÿ�،Y��7���Z���Va��M�P�3O�xN8�Cm��vRg�G(�*��d�g���QngJw�.�^���]� �,���Jb�}��+�r����&,��V��Sў$��K����0"���X^V0|���ཞAD��R◐_|�7��� �T��#��Y�D�k���dF@�����V<�J~^�4�o�7�_;��o̜��<i*!M��Bx��}vh)ǪU��(AH 
�=4t��/�m�Z'�`�P{���C7���la���࿆47"L[�0c#k��w�f]J�O��[����:�,	-�T
�+�j�_7�����iOI~���='v���e����_��/���G��Yԧl�� �"ܮ3/�T�_��u�P���X:�F䵢�,S^�B:��C7�3�!rO��;R=���,\�s
x�V�8
����<E.�e�'��i��._�]����0]�
.���,g���0ݬ1<!�.��)q#F� �b1K�Ҕ��ĕ}����ՙ��V}C�*UT-뢉�w:������3�F�ն?���Oo�nz�r�>���_.����B{l'GN���OZ���zK�3�z�_xƤ*~���<��KyG�N�����|H�R�i�G!���57z~h�E���SH�q�H�",���F|i
���y����Ӽu�{���
�˿��4f�����-�	�>^�2��꛴����,E(����:$����]�#0N�'/�d5��b	�S��e�R�p��IP���c����W���S>自{��r*���V耪���{� �g]Y/��[��@%>>āq.H���Ɲ��HuV|W�}1�c�)
l9ƕ�J���\2ğ9Y���a:SY]�G�
�Wg�Ю<���C��D8�Y�&R�y�^t��Vۋ6+ri�X��]ܫ��U�@�@h��<�&�ʐz���@9r��O�7_7}���⢠h��ⱍ�3x-�F!)ǾՌĦ"�S�̫�=͜+�B�&D�R/>�iY��4�3��ߓL^���Ķ����p�v���VK;B�5C^z��U�xK��{+i��B��
�u���5��V~�$ݻ�7u��}Pg�?��Q2��;�঳�Qh-��^���y�9v�3���qP3��7�1�~n�j�0=�܏f��B�_Ć.l����]�,U:U�E|u*Zy��wl�����H��y�Κrm&�,���G��呻z�����Į&$ciƤF������?���~��䝃�$C|�!���$UY�.m/�n0��ѕ7�S��A�e=,�A ½������Z���KL�C��Q:���E�[�J�l�?��Q���x�|?���z�H�����U��H���Ses�э��TR��Z
��|�Fny��5����,���#��EF�2��9�LI	�|3[�G���,�q:U87"T�y�S� {��X�jP�K��קNz�*7����e��E.�{���=�(�t�[q��ќOu�1�,���� %��y;�D�*\���'����{�n��ۛ�v{��M����~���}��\������/�l_�l��.�O��Iv�uN8h���sZx�������i�x���$gE�[;Z�J�aix.*xkx�Ii;#H�B����R�e�n��>�!	���;]�3/d#b4X	c�&R�@p1\��ȼ�S�+��U;	�ta��[���:���~�d:R���U$K�`���m�7��)���T�?�f����[Q���d	���Q��.��4i��p_�n|����!�k	k9a<�����.�*�Dq��(�OiEٜ",���k�BX�jl[YA�܋l�4��R@�nZ���s�XCߐ��tp��G�+��L�"ǁ��7մ�Fr�����([�.)�ɽ��4��`du�ɝ�)Qꌚ�	�c����;��+�) �2��tب���:~ ��i��V"��F�������nh���[��R��{Y\���@�WtQWR��/����ryS m���|��閔O�2�K-�u �1�5
v��5F\��sX$jO��(צDW46 �:Mēsu0T;�{}ͫx���M~�7��>�@ A�A��Z���x�D�����s_�3�A���Ʊ;_-�޹�t�$���5���5�褒9,��t���a:&7��6o��r �O!{����u�I��Cuш,�;�8M��]�
�Ǳ>��.vG�� Ǥ�a
��P��Q�9XOo.��(M����GSM�ߪϳ����"Z�2�>�?Eo#ij9��Y���J��f���5T��-��b����ks���<Z��2C	ޠ��(bB�Z�x��;�	���y�$�7�:'C;Oͼ�E�N�bQ�0S�}�A�LOxܝ6��=��\�ִ��`�'�X@��Lc87HF�n[}��,���ܔ�"1u#394�Ť���مa?m�,�B�����Ս��tl#0S,���%����9{�%��ךI��^��[{�/������W�\��,������.M�3�זּ�j�P��0�p�q7(ݺH�J��AgI�92�@��Eʠ��[�f@���~o꒪"�㰓��A��^�]
���py�.m����ꅿ��w�L�Dy�H�gr�n#��2r��ve��ݥbڱ�TR�N�_1v�Щ�`}\wV7)uU��.�z�$KX)YvS'Vs Nle�kP�	�5Y�я�.�C�e�X�c���v�5"A,���<w:�qu>����|Z���zh<6i8�2�����/0p[bW�w<W���"�����V������5����,rK�k��_�r�K�̓�z�D�o�9��y�d��;~�8%
+Y���>&|�,�K���vc�C���x�c|s3�BV>�2Ngx_��n�����K��V�_���6�c� �X��~묣����u!�ww�S�T�zx1�撈d�������}ۑ+���� 愾��%��
��FΈ&��[�H�|���%�s��v!��Wh��3��izIo�\?T���f4G����]��u�]�XW:[(six��v}��ҽ2��X?u��c�����_s`���G@_]!�|xL9��(��c����q6}�2�I���k����nWj�H�\�Χo��$MƦ�:4f�B�?���R+砱N���s�ks�y�����^>�H5*۫�bv9\�Fg���Ԋ_"�s��L�Ϣ�@�r$�r������g� �=\^SZ� ;\МJ�&���m�d�.�"x�t	6EmHs`�p%�J�h@��F�o�_�*�).(�0X��k�^��jW݀[����ԡA��"���si���������N���<c����`{�����Y�����#ԩ|�&��`��q��G��~�6VS?b�{��['�d�Q�#�(��uk����X4;\��n)�ɴWr����Y���Q��(l1W�����
9�2�������XL^���+��E4u�g��VԦ�������P���p?ɓ/���&B�N�nA�@=�wG�u^e5<��{3MK/yfns�,Ć�D�A30�|�K0�n����@t�ŷ8�z�f~���\^b�x9�n�Ja��؂`���/H��.kE����U��a�G ���ϧx���|�L�4>?Wq�}�3Z`�Hj�IL��s{[�V���4Xe?ػ�O���{��SH��*J���GX��z��&���켼�i�Q��{��K^�:#-ߵ	R��$9�7��bE�1�n�ߨ?T>���1�l��P	���!�fRK���q�Y2��WK��Cޖ�s���}8�\Iّ2ٌ��[~�l�z\����]}	�>�IX�<�.�{���0h�e�o��(�gh�U�`&k�!��`�ٷ�A����7=D�-	�$\���8:�r<�K�ЭŲN�ބF���`�t+4����M
���pֶ X�YC���`���w<�+��僆�~&֪���b�:V����b�s������T�k��-�#�y�5�wՂ*BK�R|���	E	i���>˅v�HK�M��vH�G���^$q��6��]?蛯�9��)�YH+Mg_KF�o�����?� '��DS�5(Ã&��Oho�=zw
%}�X|�����[F'���
�0eA�r����H�,u��Png0r�&����a]������%\�	�j���b��bQ�����,�@��3�ȃl\{�!-��D����;]�!C��~�D �R�?�b7+�$m�wdrƔo��tB����%IH��#����q��473�{V�s�d�)��j�v6wXI ��8�_C��̭�o����)��ƚ�ݓ��,���l�����-*j�|�3_Y� ig�5;<�u66��BR�%�)�$�ԺhQG��5��'|�U=|��I�;2A�g���V�P��=�y&*�T7������3��V7���Z��?�e�:e�()�p�E:�.�蝀 ø+�[�j<;��F��s.�M�jq�)=*o3E����P��jN�d"/>��I���T_|d8f�3Bv����62�Y"� ,4��^��l�Q�D�4��:���:`���ǥ��mD�R��[�u��>������f����]
^�]�^р��!��q(b�n�4�?O�xl���F�g��%�ı{���YO�A:�߳cNU�-Z�/2�nӠ��
d��[�\~��~{"�\aKLu�{�˟U�#؅C��d����`����e�fnFV4|V�.��nC�ր`���U��em?���ss�ʫ��o�7"�e��g|�[T��Y�G���󞃈�D����D9�&u�Ğ
hU] �W�*<�qV�:�fH{8�}��U�Kŗ�`a�'��6���Ġti�Ŵ�B��r�{� y[4nwU�7g!,!���OOȘ�{A�|�50C*g�B��� Q��V�@��&�_���Y[	�}:��RR%<8[��R"��%��P^k;���1��0�O��A�{�����g)d�q@N�i�v�K�T��f쐑�:1���a����>�i�J�cO���|�M^�9n��uw�=1����nn��Za���z�rBe2΅�>�0ٞT~�ʺ���k�+�{G��L����m�
n�_`Z,��������8V��R �\� �%��\�|q�HW��"�#s��j@����4���������[�oq�����y�xKם=t����N�ش8h5ҥ9��V	���NL�q$��h�pv�JC'�`"?�S���"
:ne}�L����7'Ȃ(@��d����@���k��Y�{۴�&�!�&�y�E6��}v�Ea=K��d�h�p9e���'��<��H�Q�\mX�0�ttQ'�9�x0�^c6d�k|�[4�)�[�E �\
�!yJ����J�%��*"���� ��x!�^�>�*򒤑��d	��= �+��R��A?�%bA�;MS:N��!-
�$�#/�e=�� ��(�w`���z�Ox⨿ā^*�A��~�.H	�f���Yj��le+pK���hs��	��](��q�N��`� �`C�̴U���ʵ�W���h'��Ϥa���U�u�k(�r�;��^��q%�~n3!�ҵ3���wʼ�YT_$kPf��[<}�h����ܣP���Z��蒈v(Y5vh�Բ���qI�R	�it �����,��R�<�4������?Һt����(���B�z��*׳�*;&=�������UqC�G���}��:Þ~�F2w�BxgA-Rچ�ҭ�\�4H?o��F��eK�5քS_�=R���2��/ϴ#M���[����,0�� �|��^�A��e>59��o<�5�Mf;X�fT�׷�2�����IFs��ĳ{���W�N���Գ_�*�	��3��'��D0m���P��%o�b�A�j��v0� �P �:gӵPh�S��$�`��+20E��[��$��M �2·�8�j#b|�-�6&b�g�^��0���,\����Ȥ�/�s������2�J��W��}p�І����^w���M:J�d��"y�A�p(4s��i�ua�{���r�蚇\��4���DF�L�-j�n���t��޶��J�	�PƧ+��#����.ó�7o�c���DF�,��A����(*��D	%o���\���w����V�_JN��jW���Dč���ˡ��ޡ��Uy*z���V:���M�~>�Z�3��_S)�<�gz�%Q�rT�󩈬�q$a騏��}+�à�1!�{�D`���z6���*�Dx�
��%��!�ą�E��@�>z�<NІbnaU4��<6ZJImem4�=� Vݡ�`��m�ʐ��(
8P��Bݚ����2�
�a��[{����yI���7آ@�ך�pc�txL�U�� 5���ʎ�1]
Ł+���LV9x�ٵ�,*UA� �-�`�y��Y����v3�F�W�j��[n,W��{��[����ı��-@U���bi�JDj`'����Z"��灤 ��p�u������I�Yؒ�,^�cD���z)Iv@-���\�xa�1�"D��ƈ�P�˲J���)CMS�E��ef���
k�/�;者*�cx]e3���	���sG��ò���E��Ws����n���>[�B�����^N��|��#�\vgu�����j��2&6���a.A�u��n9s��+�wss��0lqF�>J�b�
���k� ���@[	m��\3h+s�_��D�l�˳Z��葤�NsJ�:bM�a��e�,��:py󼾀k7���.ݘ&�����S��,�<5�����x�dzB�q�Њ"8O&oe���Y	��E.wU�^����%&�uUXئn�z?yمa/����Q�ɹإW\O��\((��[\vT��c����=z�.3G��ƾ�<͉����Ͷ�ǯ��=QO���]_h�[[Q��%9k�.e���'�T4!I\q�;� d��5sq�	���N�F�������ά��8�*ƀ�u�
b�	Wi �a��	O�
;e<�/��$�����I81�x^^6Q'�\�0����1��EpK�0�j�lL���*Ӳ�����*�:�o;}D��5����=�<j�`�b𞜹F2sY�b�x5ږZ|�h��ao�hA%"6r<' �xM%`N��[��@�U��}���$�[rͤ����6�N¹O���K��B���Eф���5HWM�{�����R���J�*�����vѠ���9�e[T!(�+V�JZ�=]\�EK��`5�u���Y��G��g`A�k
���S��(�z�_�	ĉ���:̍b�rJ��vb$�b�i��������Oj�{��:/��1��&��ûB�7Bך~Ɛ�(�'�-ԣ �5s�s��͸$�4�}���8�����!�qu(�Rm���ӑ�2���
Ɠ��X�f���Z�|JE�1w���F��Scǆ����-S�_*�p���ꬌJ�Cd�#5��=���sĈ���Q�ij�U~&/;�M���%D	�������ԫ��v*��st��؇.q��//�$��  ��̵2_�_���`��Q6�nY/ ռk+���/�����vV�yx���������C���U�CGЇFv�����ĭ&�.�W=�X+��ۥ�M�Qاl�c�
	�l�ۣ�[ԊK�G=��t"�"�K:S.�t�)+�s�az)GD��$�C6U�sUe.�8� �at�Aś�1Xv�����Hԫ�ݟ۟Z��_p$Q���^�j���AF�7�ŋ&[��d;2��G��̀���?(��>����q��ԭ�&�o��"�
+��[��}��m�H��9~*����1"�� ���|ꞵ�p��	�z���5S�Q��O�0�Ӹ�s�H����Gx|����?C��z�u����:Y��
�R	q�cy*��y�?Gi�y]8Zo "v,E��lY�c�E����?�/�)��T��@� u0��Y�,���W�5V�&P>��!P8�' ܖfv�.M�~���v5�4�J��(sa�Z�<Kҽ�r�~ݾu�	����}4h�fޘ5@��I��yj!4츓׹'�Sw��� ��u�h)9Z�v�9�|xݴ�=W�q�,�����tj�SE�A���c!�ˈ�����C�=�^�z�r0��������n�)| ���Q��~4[�����/S4e�[���A����e"�RCa�I��;sK!T. wm�����Ά�$�m�Q�
c�=�#�,)�Ei����Eڱz�������&�G�N擣�=�H՛-��_1O,�c$lL +��P���)ѻ�t�����h$�(�97�9�8��B9�+n2d���'�I���/T�r�4�bV@��'�������
����S_�x޾��8z�Vҥ��
��U�����4mR5���m��<g7`���GTB�WwU����۷�9�eI���\�B!�j[ؖ��=w��[6n k���i{�ּ��q�
�g����d�X�N<�o���q�ʻ�~�2iiqkG�hM��6���ԂV����2�9X���?|�rڹ�Y�?���O,N�UBӨ�yŶ!��2Wx0P]��h��t��%����D�N^�L;Yi�����������DE>/v��M_�:�l�¥������|>ѱ)���)��
�_�>���LL�"���q$��3N����t���F���Q�Pʨ��"�Ў��F-�e�K)5��#f�^��9����&v7~D|N�y�;U-���*W�5*b�g�7`��E�GM/�٭�6/��S9mK� E����VB~.<��M��G�`t;��XɣL3���Kds.�+�H��y������X��[m���-UzU�s.p�]���OȦ�����<� aq�S.���<o����6j���o¶�av����V&��H3L`����!�3�A{�lVID��9�7��m���T���5�"����T���d�����-�qu���1�T$i��판r_�0�'[�pM�P�ʅ��_&�]ߛ�"�.h~�c�T$�.Ŕ�^U�*�!ZyP���0��&�Ά/I���2ˍ�'r�T;��2Ӌ���:~�q������Sh�h����:�OM�ob� MCh�&��^d��ʎ���՞|�bR���YCPz��wud��AEk悰�G���׆��HGB��*�1�M�h�&���y���H���?�%��ϧ�%��<��/�Zb��+�UNC�Ԝ���Yi}� �{s�_��	�;C��6�2apaY3�z���B��l��p�l����|	�	����7�����B|�sN����JXp��	\s|x2��i�K�۴�e��;m�0>�I;�pK4Ÿ��7�*���暌�&SG��a�O��#m��DG���F�	 ��M�z�ȿ�*d:&z����I�qw��S]�5��~�A{?ktR
m�mUSǯ�Jc^ ܀v��q%ؕ1�ӿ�2[�nNF��4D�܋R�u�sGLu����Uٔj���BK����9|�IBX�5�ӣ����
�����o���u�`�ja���9�3�^wM�Y�O�Qovw�-ڱ.j�d��p���}��x�c�H�@�����g|5��Ը2�}
��C�ݻ�ݩ�V]���tM�@T��#-�mf��#4©����_�{U��pٛ�� �K��Z s�`}��Z�s:
\P|�,l*��QU�\CNA=n����)Kө`"-��e<\K���J]���71�=�%FfG�P��c�f�N�>Vv�{*#v~)�@���ϭ���T��p��N�!��Rf
����jꬿ����dR� �u�FpJ���2���ln��԰����)��&p�Ђ��WΌ>�Lcr������A}�9Z=;��Q�;��f�E3U�����č��$PZ�lv�)�_Gs����7��	{9Tg�٪�|�mW��&����U����&o=�O�ۙ�t�	,e6Oy~����X�z0��f�Sr���i�̐GxV 5�^]�
�ؐF�������y�Z~����W��@n�V��@� ˥C#���"��X�T�ٟ�I���wR����0,��]vȢ���|D�R�N���z��K����f�Z��4�$��yH⍞�m��)8�2��_y=t-<��� ��2�5�?@��n'�IW�����Gc k��o����9��Aj���^3%!��9E��D����_Z���h��C��p��\��m�K7D+���x�Zs��L��c�uX����ą`��0�	�Hۡ��6egl��s4��M �*�.8Fw�_�kE{����i7n���"���D'�G��fB�H�/��*c��oGymj
IL���&"t�o�&c��s���7�z���Þ0�����kqf�9��gT0n;�G��4���~4�)�����<{̢�ü�PCE1���C�N��uf������X��85���&�(��w`U��l��U��&󭈶>������S��\*��W�<޽/Y���3�����2�r��E���x�������ou� ly��?5�� ~=۫���G��+����}#���g+�4�`J�0���`���̰/�~.d�&8ȸh%m���vtY�t�(<�D�x�qh��w�@���$��,<'�gZm<s�5Et�o�#1��(G.f�H�.�}BO��mGO��^xQA��[�ۣ �*�O�h��ķU�dxe��k� �n� ܒ�E�������q`x�!�{���߇���[��BU A����oB��Ɩ�ҭ��	Vڿt8J�Ul#�2���^	z\5�j�l�&E�]�'���T�o��9?�n� �磴���0-�ۈ}6i�RЮ�.�h��VP�o���nz���qw-m�~����$l4LF'{,]�������@���,��zX��!��#U�J��J�.��F�f��''�|��=�� ֙3����_s*9�Αn������]>��vRD��Z�(\��l��p��U��x7ò����׶���W��u!j%s7����f��'?���e�ߣy�{�^�s-�3R�[����M 
li,��hƆ�8��)����HS}���3��fnƪt �3������O$�x(�rC��C��$7��Q�_
�W���]��ϵ�f�@�iڔ5h���f�<�����	vމ����y�[�I�zjl�Ĭ�[���Yβ����Cf�a�i��(Z*�k 7;Z�K�8�A�o�׼ b@�lC�n��f���\�����͝�BR4��B4�v7��k}4\�ˆA�ˮ*�M����y�7jA�}6~�ѕ\�G� ���\�+
�����˨�dE���VI|�[sH��J��J�cHv��v޾L�qMj�N����Y@���̈́���3��y���M��Nʓ���^��|_K}�����i<��u �����h��4P *A����div �{�D@Z(H��K��Ǡ��Gw߯��⣪^k��@�ip������?�d��@P}S6	�n�!���_:s��H�vWpŅ�VJE�K�$9�+)�׾3�D��5�_o{�=����Z�Kbk�X���!�$��[i@��T��r�j�_�rjuY:�K!j��h,�"XG�r0��kTi�V8N
-�+���K�/�q���4'��� >I�V������W�������h���P̲4�Ҙ�֫�Uo���g�9���q���@;P��_٘��h�KMr�a�)���e���T`���p�Z���|��l$�O��Ĥ_��IQ��aVO��2ʵ{Յp�p�	� sK��J�<�"��sޜ4�o�$D����p|*F�`���F��w�l�!��}����l�X���:���J��d�b�n���-l��gE��%�Qca��U?s"�!�R�#�����v�]�ꟃ���<��Y}6w��/pY��ؙ����DR�
�N�	��JvJϚ!��{�����P�����"3j�;��D�w5UD�wK��]�9Ko������h#�l��������<3����#�������2(*����YhX�2���!��+x1=
]1��L���iiD�|P��P}{�3lس�_}�������e�}��$-�| e%�"��Ɲ$����P#���-[(���8��=���pQMf��5�p��:�X<�1t�=�@�1��[�Qh�<����6�>�OU|���os�Z����lOf