XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������ĦƗ����:<� �2U6�B(��Ӳ��$^�;y�Z��m��zI�\H���M�� TM��B�r6�n�Y�^E��4u���ѣkLS�ޟ���N�	�!�~
k����z��:��S�;�����z��Z��i ^pZv��ˤ��Py�.̥�pz�ӂ��W� z�
A����8��pGO�������`����j�!���`�T�A�Z}Dy�tt�p�Gyw���QCv�2��[ʽT�<����#i�Ax�6o}�V�������Ne�pà"�y0t_3�M㵽sp o��(EFJ�sE~��G@�pC��c�4�J�T���}����y�H�)#[���U�v�����7��6/�t<�m���7Ovu5I&=܀���b�0#GMȭ5��iȼ�(dh�D��ȩ��c�
_3�,�H�A��+�ޥ�f���������n�TL�e1����Es�JU�	G1���aqH/��x���,H�������;\<e ��`��h�P�qA�;��o�3{��/rd�֧_^ًع�iݯ�K�0��{'�%�7+y�Yjp�a��X�! XH�j"�O
�˿� PVr���X/���q�| 3�_|@�"�?kO�z��8�A �����8Gx	�},;��E����ab[(k���!Y����JO��Uc�R>�跡bz�_'� � �*@��#`S6�%EbN�?�V�A7+g��9H�9p{g~o)̜U7[�2�����D��Z���&[Y�BXlxVHYEB     400     1d0=��^kS"�e�r�cwu�c�j��<��(�f5W��{�y|ʧz�����͒	��=�NGw�M��Z�9��0R!��v��E�
��S�Cl�2%���f�m�_�?<9�8������LO�ߘǫS8�$;)�7/���k�ƾ���h�o��l����}�v�����:�Sz(���F>��	�� ]J���\}?"�9S��2&��1�
�c��P�-�8��'���a�wi]�v*J|�"�R���8V��G�J��n�4"������Ri���k:
Տ֖��cC��!�_&|�mX��ݠ�,[�s�j�����u����Z�:�Ѫ�~-���tK��:G�G��@-B������Q�~Z+!TX�@�q�׻f�����(����a��}o�#�iP��28Y��	\���m�o.��gu@��(�J��2_�o�7G��Ҿ�)���i5��0�XlxVHYEB     400     130������� �NW��U.����ͥ!94�/^w���eш��rg�2To|y3�D�뇃Ff]l~ַ��^�����O�_��>�QL���w�	��ݳ����1"���z_����ί�k��i�#��F����)�A�� ơ4��o��vҕ9�v� `�bP���3-Nhp��4�R&sE���xh�B� H�����o�M�3#�r�-�f�_�-�'+�����v5�U��9[k:P��oأA?�q���I�P ���@ގ^�ܸu�r�SMT5jI��cx �A��:\)��t>�S�XlxVHYEB     121      90^ژ��TX��&}c6<�:�)yȒ������a�L�BM��I�ܙ������w[�⩶(�l�3C��L��-��T�È#���1�)�1�{C4y�浹�q�j�5_w�^�h3|p�Ŕ�E��ƥ�SV�{y�
�~W