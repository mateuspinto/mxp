XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��^{"Jr@�R*�G�,tٮ)�Q�n������6ؤiy7ԑX,�a��y�є��͏{�U�\�J�>��x �@2���[�i.�cj����g޲.��t�U��Fh	Y��Du] 1���2�۩��͊��g��U�t������(|����� �>�s�cԬhS�Ʒ$�kS̵=x�9v��.�{�*�8�k�$+���v��:E�^1��n�?Z:�سOHɆ%N�Y��(���"p�c?��(;T~9k���h���e<�i��n��z+�y�I�;�9�!v�Bh�Y4lՈ�?/�������i��'f���	�/]2U����v�z����/��������Tϐ�����Zʎ_��I)�JX?�l�Gn1b�v��h5:kZ�Y�A���y+�3�9H�����h�X+�݉0x��h �e�~�TS6�_e�C��B�V-4Գ���S�:�ǒ�<���,�#�ނa�.���J���T5L�͍��讲�'a��S��rhn�X�CH�S�edj��G3]a�w�=���A�C������nw,a������N6Cc--Y�����"\�S��<_����5��c��B�-)y�%��&o��ʋW����%}��Y&���P��M6	�W�<h���W`/6���W82@�ڕ�S#��)"�C����`_�B�(��3�n�+=��Q���!Y#����U�`�u�a\rs�X+죭�t,���~B�gFGCQ�9ӈ\����/R*�=Avu  RK��QXlxVHYEB     400     1909�h�E�82�^��M(����Y��]�.���������R,����X)�q�ȵ�=�o��;�I�W(Hq��-�L������I�jީ��ꊬ�	��r�����d��b�D���H��Vȼ]W�s>�I��lk�hL3U/k0H$��z�X�u`��栏�\{�Ll	VJ�F�����E�$��@lG4=�9m�zG���j��*<�=��_�V6����ɵ0��*ߗhX���D>�`�s6>��av�VK��>]��j��â�9�M�
��*��4�@櫌�SMG��M,Ek-W�v��`�Tw�Nk8zu���9�<���y=S�����DU&��u?l�N�>��T�i�"���@�s'����x��݀�~��C"�ŤC\x����Mʒ.<!~XlxVHYEB     400     1a0�~^�. ic�<5
�3sI2��4dW�DL�),/��`��P�$LusT���zC7B�Kw���;���1p
RG�,a*������1�-�׉ٸ�1U�X?Q��^�M�:�i���5{u:o��EF3)��:�1�p,�9'o��܎J3��6A���S$n��^
w���	�jahz��^W����.ī�{b֖����i�+�ޞ��Ӗ����I�U�p`z�NO��>���W���;�S��2_���# ��7�k�$%��?1	��6c����]�]z��cD��E1eM�Y�П��[�E���)b~Q-�4�垣��s�JIyY'��	2?AIV����JIʄ��Aш<k� vx�e�:_|Vr�Q��YR����TЊZ�9��\����	�叁��l�XlxVHYEB     400     130��z�NUύh��p��׽�� �Ĝ���F<�0VP�!���w����Ĳ�F�Ң#��/m�2��k��z`gV����;h`�@�q�D#)��u��ن6T���W���Z!.�5�g;@�r�tB��f�RujS�
7{�I��,��=������-Y�W&�A���V�I�u��o���`�g����Bf���<���n�_�ڭ�Z�Hµ������P��=i��d�H��$���C,���@c�9ĉ�Kn�º��ґ���\<��Ld�"��\��֥ry��L�=]��x��.:�_\��XlxVHYEB     400     160y����!��u�g���ĴmTM�����/��8��j�J���9E���{v~f�:Ĥd����>�
D!l��A��+���U��txe�N�)��P��gb��i�BC�TUҮ�J�z�1�XK)����K����X3G��"8��Đ_�$P�=��B��!�����X�խ���vv92|Z�	�]ew{��(~�d��;pǿ՟��xN�_u�m�K���T�W�ˌE�s�DdkK�;ѯݚ%l;u5y�E��l1d�~���*V�ևM� P�p���q������2k?�` ���� �眫��
��PL��N�(W��p[bg�]�tJ���?��eYi�M�j�XlxVHYEB      3a      40`#���tڦ�td��Ȼ/��4W�e�S�\R��i#z=��xs�*b��SYK`�u'��5x͠