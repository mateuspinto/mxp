`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7472)
`protect data_block
G/KYpSBAd79GEzV0q5GPFwtU4R7SVzFGB+21nugi/XZAoqgMXXfZRzh+mvfN6jOfRdMb2rLztfVA
2L8wKk3ua9SM5iV2Fw958EJ5qm0w4DAwKrIL/8KzdH9TXqpFwHV4BvZMBXoYdrRIM5UcjkMb2dMj
O6Zlg+ILt3ekBMUM8z0zB2B7Hx7vMK1cNwAdWC4h3JuOhZadXwxaFgCerP+VU7tGeEgR248jXtBV
KAgdYw8rMtIAVqolUpXeb/t6cBYESRkrP3dwL8XOCu3ZVceZ2cDqK48O4lMv6AD417/17cDOVGv4
R74E32y3VxfGI8TUBHFg8zWrw3ANx3tt2McScRZ9laK99e5U2Ciu0ut3DBF9TSAlGZF12+3TxGiP
/mOln3m+TALtY2JbLY0vEeFMMG50f31OBeGzSkRY2U6FdclH0hedcIUDJDstWBv2NpVHwn00cL/6
uj4sEUJCZxMeasEgcp0dP51I2Umd68iXfaF3bOz+E7eFMBusifTRDQcp/sG8LemOjIe4+M+WzX8D
WZeMHydAdw/6O8lDmr0WM3GBq2sZWwUipALzSF2yptYWfubbl0XW5l1ejdeqfQa9jicvIRz2g5au
IdH4NeThbXKv27EHtP6iRKcp7o0oVPNc3nOfr0bD6GlTqBhPeRpQ9KEmy/1CAKmVYWOjLc9Arc36
KzLz9JfFf+L/cuuXvw+6tkFz1/6K3B/VjlUR8K95FBO5C5Em51w2w5OFhYgXlxfE7ubp7pPeoOqS
aQcMoOmqMmf9ZhlIoFBMDGcfGQoSm4rKaeRvAe0EfoRW4gpUZUv8kEfVYIftyXpAWZ6mUsTw4AyI
WZE0JzgBwD8okV0mpF/j9nuJBP/Aklx6wj8TISmfDbmg5LXSZ0lRtjXdjrV3ZiYJgQj3Y3Me6I3C
Cic+j59nkKWSwDB4FY7xSImi2no7vIbvL337DZUgU/JjHHnfXx9NCI/IA/WiaCUSQ43BYoW1E+Om
FPcm69bqLgR5prZYagoM9AlCz94oYK4bkXL8M2xG+6gJgns25jciyg71C2A8wcXlq9O4c8dQeTEU
5rM+/INgj1EkB1a9IfBWtEEBXKPOaWzwbO3qMyeevIW1OSekUfXgNu4BHouuc2cGz8O5EqYhD/Va
23kTYjeaY5fuo1/m9NO3Y2mPUoFP72Y2O2Dxovs2Qiv795ZnTiSg7ZNJDODKYJFuAwZmq/kmNyDM
jWvoxfG4Z93zmbHkV2QIfG/3lDwIi1MFsc1xNgjVM2KIBbTMQKS5uckgf7Ltd5Vv9IGV+ANQWyak
SeoRs0dnNRi7gsv65PlsHI39LTc/bDOALGgNDmlZGD1pTBBY/VE3Nj92tds49/J1IoTw2eTuR5bA
3QmT5eHn8C3V9MqjM7u0cDdIyR7pFp6odt0/px9SyFMY2OhMvs/agVR4dL0CDio6OmIXanZw2yjw
EAjb1J7iBT5IKXnpOiMbgDK5ZEUDBe8PbPNPDtt0qQbECYxnPd/u1kca2XC0lnUinaDOmeKG2SgM
wXnnczrvTTwGaqQFvvj0ofO99HeBk9zbfhg7Bh7+xeW1/ywxP/u4ufSsSwHzVDWpOzyaEKMdvfNL
GoD7ehKeHCE31rxuPN/rKp+LFk8zpgiW0rWf7JK5MKQC/7OW9+tURLGO6sLvngjhqBkI+SNm3DdX
17KfJmGFs2+G47gnvBvTbuH6Hpbg0+Xmdd4ceQtZcrZKhcWzxxp+77r2RXPeWXiXkjRDe0xFEmyj
zG39cl3KyIuoXJkv/IfY3iyMM/lrX9CFP1v33J52AJ135+GoPdGwcRQ++GxDZgTb2QSf9GLp92V5
dwHYPmMHqMsfgFJjHvT2PdfLcppLBpNsZ3SqDsK4T5TevWizBC5RKZXAp6jhG7NdI/8+cYSxmNjz
j2UkPhyCrvaidCwUAAto105fySjz07FlwYfR7Lay83oi40DTuviU62vEZbF4duQ0KOXLo0DEmCNW
fhtOu+EfXmMb8AGPbQABuckdp4UzNh8TkZdRHWjNAPRsnomY98oxtfiQi5wnn2BpqVCixfa6kT8+
ohQsD5nOti0D2claggEaOkPcZVWfKuO3eYjSO1lFahulgWmP/CcDc7h0uQQaCK/RBTfMB6tuWP08
/P4hdGKZX/sSeRcO0Qi0lUIV2sK19FtUZwLrGg+MIwRPEZW4hpiseEyG+wofEEoGc7RUcr5rtvDg
qoMXrrSFMaSJ34bK9wXNOkEwt0tenWewZPiLvtZs36NFJPIlcKfIxYCbofbQdl5sj5y/zxVG/aFf
MQME/WeC0M8oCTVd+T8PYfpgfSE1bSHdkRaSDOp3pDLPL+DvKojSiQ9OXJ+3VpMuunA3PLofBtNO
zDi3iviyCth8FS0GabFOfyOZU1T6A+26ANWJKLl0IJ1WNXBRTJaA9TeSUyV6Fv1TrYWPCLbXogUP
BSVVgztdyfyljHN61GnT4gOmugMmzB/XQbNk2G1U93L1TgeoAkJCOjGNP++uHKliRdKfdQg3gEWZ
opUzc06jADPLEb5mmffwhjk+Zs/9ahRupBb0d8VdGZ1fGQJr9m4WvKOg+EX5VEY9gmBPT0s2hGv2
UHHfpM3sJt9BFhlOWBOB8NNhtCrLzTYvqTYf+xKw4m1gq1UBxhTPOMC6rYYTelCuGwwbda3e+ED/
xudQncboX1i4GKX/oeL32ssb090mqhvKR9vCczXyaYcQc5ATwJtvC1/KGZ8NDPFZDg41eyBZUXB2
Ho3p+hnrWQrEZIB7tfJO9YqWpCqOf8SYdbkqudyjKfzS8A8wqONnFsIz9sBk7DA2VwBccUtul7Sj
c1s2g2hFEPqHe221mOKGyJeZ26ctvdOmalPdnJqfVGCZW2HvW4kOWEbT4Wv4rGeNBSk2m8CmSz4d
NTCYpwZ1J9d2tt2wBR0o97cXrxywcu8lJj3/+NGWBGQBAkZ2VTHVpSzFa2h+XuLmKT18PlLYpIy8
9b1VKhNRSTWXWNq/1qdvahzZZNmg1jKeHfqSDLe5XEgYgk9xfYzRvjLt3DKtsa6Z5rGAjwQz19DJ
p63xvzvQfu6K0BMWX3dsxJDN478/bzKcwyLL7HSSWz55EoQhrXU/Pro295IffpdbkUlubkSIlFI3
5e6I9qcSpt4XVEJ3Bui9hpD6jtV82I6w18XXJf31Ywd6aNdb6ASLQmA0pJ+rk0uCgVaNsmYEQer7
0dPBn00xr8y5i+LvZd7soFJXl1oWvqoR6472WU8+RnYuV002DCa9Opflsn9uFHzlF2zdd/PiUeKO
sY74Cyy8J7eU8Zp0dRFRW/aK25W4hv1QNJ2Dx/+BWFZIobAqHr8UXyhGmBkZsxn4N1+3G00JV1zr
zhuR2rxGDWTKsquUIFA6ZdKTTHhdzfSXmkr2yDYT+6u7mxJLgmu+kCgGemL8230F7E+Giu9+bGnr
PqEh6Hd4sj3uhWh3k4gewgCMhETINAefQ8Hicav+KpVJyk4iit3RjSPYBEC7BHSU/OvItnhCW/yx
uf00/hIWaaegya5/3cqJDdwzS1AgZZISTFSD4XS0Ca/OH6K8DSxZku9Wab4Re0UTTJ0BIDaahIuZ
IHhqJSOU16srrQ1YgHv6mAUeb6HGElRr0VYPXXajTAoPpQVKg4LUZqZ8q0ZpQYWuhGPi6ZUz7Bnx
q6Jql/YPPVthSbDWUmLBHwCPzPFGXV1XhoWYQfiYvpQ0DkOewUPj+diD3I3rqZ6uCbQlux5LPA2l
rlv1GuBHConUnNe0sThYEb2Cj+mLGQUHvteMEC2q1cdunY8DCdPcOjbETvP6P/Y/FPVBvvo2lkDl
ZKF0tbZBmzWh7W6qFR7lM6O3TpkGo48h0oqDzVbze/GLz2+y2f1rrA05upr0sDrd2XtqFBcUi6JG
at3yHdwTfxX3zsbmzSjhrZoK9eBgo310pK7Kj+4X6y8FItvwxIU5Fmska9xrfXvJbdjccM4D23Wd
9WiEmWldRG6WtqROqSGh7NVUbyMMbDH1M+d6ssex05qwmZmcEarcmZRledTJdHbQP2bf7eD/yqMB
+itZHWG3HEMgyMjTEW4TPpusLCTmDvLR12PEDH/MchKcqmWq/yYEQXZ9BsSxpv8bt1w8F2K70PJw
CdcXuMLOF75WbdMZGJYughcW9Uy1Eo4nEbFOIeFNxTZQO4ajdPxTwK2uIqc2yygtPpVC4DsVis6z
A4tFCiAfCmseZ8XqerMce/pVDuRw6H6RIoJljgxCYDfdt2K9fE45lIPqQhx/6wL9Z2mTqD+Zlz6C
FIHMejt1hxX+/cgL7lbzUPB5z+RYOLylkVMdq05qG9F4qtC8CLSTPbU1nU3qJ1qH8qnpip9Q6MCo
ObrJXgVfOk/aEfYBdVtnkCsr7wk7CrkQCtWyxwkZIJwkPj2eZj5xcOYQ8duzQincsBoIGEsqNhax
HfJIFA83LT3X1uynu67Q5b0l2PXX8QAa+nbzRnsjSJJmrBupHgYj/uTYodjKt23r8LfsWsAJ9EEt
uOAezQgBMX0J248wHh62UZ8zSD0JCZL8f4/35Cy1nUCTG7yDA6zxmWgBUwIpDs/SalyHI6xgl4b3
MLmfRWC8LhDdlY3TtXwK0tkVvKXNKFYqsgBZSqdsLBn2N/K1EMKnK86Ya/kr8Ewc96v+PtprCDxd
/xZHK9XxddRE7V4wyLX8+XxJE2MXmnYqEzN1jXSZsWQPAw1ssAVAPbQ5TZN64SGKqbAXiHRZlT/0
QKyrt1LH7vEjpanDEBBDOsw7/HQxZpV7xDWSzM4fwD8uYxboxU07qCxqZzF8UkeJOUat4uN9VR7k
g628Y4ZfdN8gRO7zOb4DqsRiL1lQ5ZHaDxIKOo9rMZogezNfS/ddiS7rXA+BvwbzFLRXeMFhcdoq
+7V2vTfxd8t28RB+YaDmGB8gICYT+3wuS6PnXjgc8BkhJHJpU0LWEEeDG45vXRWZFKyzV4cEhXjB
BELCQNhI7VLM8jDv2oIOpyx3/KW8GsFvblIzcunFi4Sq8n5VYjVhtpbrjGu5sxriMmEFL6fAlF+d
TNoX8kyYEzJhfnCy3n7rjk+r1XzaMjTgbAmD/eMsYfwHMY1SF+e9nZJiPowPUCjA2zE3wc+ZQbDC
VKtAnK0aHUiFKMngy77/Mnxl5VXIG8o0tsvp1KM3iEUj9uh4hq/C0zl5J+k+euoPQlGilhb/mCzI
ULKxhijJ4Ey7bb1D0PscE6VwX9b0SZa3YaqnQcuYnzrKgiY81HTXBWGLjBWrMWiBLiOpQ3IeThZH
s8xat4i0EgpKl+Q1tMFa3wOm9OSg+tERf3sxjjmIG94ShnJUUMZvyxguPtDCknK7hA3mavQhnDS6
zEAGlBrKrGsNtaOPy0cdt/p1ThrfYCI033S2oP6peIyQm60SwFINRrU8prIQHZ+IE1J52HdTB6BI
F7cbKIDrWC7inw4HyGZDLrBgGxwcaZ+ziHzKzysOk28xCcraDrnbuOfbRLPTPOH8xzyIVnJ8S4Dc
b2wbEaGSf2p6ZNf5PhDtc+G9LBoiVYkOg3iNyYxdnzxWTshtcALcRVBJgJWqVL0VSUXimCtp68wi
sMG15xqgz7KxyvSpDNRRtS50gE/+KrFJH/nKaAY4yW5+pQ+72+JdoflgdiD2T9HUauiQ+qDjN/NI
owIiR2h1x6lb1NrM4mTUCxz53qrZuyIbW5eppwUCe5tGovWmm8Q3nrJzvosOt7N5IGOvWaEAq858
TDfeENCGA9Cw2HBQBC67hrzuQiavju5zoUdUtWLciukh8xvck2wwVoBW7MgVpZRhKKGMUz2GYj0t
pUslZx3d1AMYozBw3LcYYSLDOV/+yirWSyQD6akxHOjEpgR/o+Yesjic82HiqCIpoXm1qVLBsdwa
WdA4r5wbFnop3s6sQMtvHbKE4Vu8XA3QfgLMyoFwJ6dtajBN1WHtIQ4n8HA8ft8GF/OR1sE1AynP
Sz3LPRopY9KsEmQL6YoNn68tc1ot/R5wL+Qma7RKUV6he1VMPp91kS0kmNhg+NVRTtc083FK0VY6
zytYbDDQDyruXMnfnjX3wNXJFyZjabeNYFHjDzm8A3c3CUvn0Fl2AR0O1G/mEIolFm5j9GrLwEa4
kFSiHvBP3nzdTeU1xuYBP74qyZvHhZxLOZd5isEuSCvFe1iJK+JQI0DRE9UZP6KozQfQnF4dJslD
mfSc1SIXMvazr6+O8PQ60fo8i8wteimOp3Xzxtw0in6cpRahl4NFCQTaktBvb2Z0TZjE/tbfiZIn
LwxPZl4EZ9EL801syqbdCDG0hWNA7wewHsOyxKcIqyqbWxi6YQ+588QdRwpXH0DZXuWCG1pgKuot
cO/awZchkq2s6bLSl13/WPsFh1xTMCaaIIQFi+V8hR1QU/KtUGjkDp6pCqeYhM2HeQzRgL+a+hpD
Cehriy+PXmjLJxHBwPeKgm6Z9Sh+PNs3W9ChlADbfm+90dpF6y95XUOL1j+L7u+h5nD+XIvkhZRP
OQoO4HRGfU79KUxgp+RpfZA7i1urSVqB0gL00HQL7/xXbbnepIuhrgUgsTkTkXHSFLf4YFW4sXGo
MI1lcFprjUvp7J8Hy7k/hS0mqdo9UPVkln2nCX56LwkWYJ4XGMS7beHc36PjJkHNWBtElK2sEuWF
6lBM9tf88Pt1j9v7jMTM1Vtz7X54nnX1oVHqkOeDLgZK/XntITETXSipSdC3qrRFk5nXerD9QDr8
nISklXzBr7BKdbqHDS/vIWCqkNRu24lQ4W/BfLZWU6PxFtVSMssT2I1OAxOBXjqr5+oP0Pq+MdZ8
uH5tbqtGavxJEADOHkJUQIb2WFIm87adQrbH8ll1iRFTuCxWxuQS2MD8BBa/dTOevM9bEzoSNE/W
/BHuao9wc/U539hSH75/jVrV268CtGrfvQAUXXEMTURSL++YJ67TXD8SywXZq7MkUw01AX/+hJM+
e0l5cvN6VfY1RYRkTb4rRN1UiSZzJDbLbS3NtkNbntr0EbKU/xofuaMNcIUWqeojBPwpiP6dymjj
UuOrNNQZDie93pSPPVGwZxiBMscrIuj6k+KtXPlySBmZZdke/RkJ1iNFAFS2YlmUK1DE0i5eSwXn
xMMuCK1caz8YIj2MlUlD8YvMERkxfJXALgtzEyY6jM0QbuK91RXQo8/Qsl5uzy+n5FEfncd29PJM
wHF1wDvj0cRwRpUXc4boOTm5Mq5mDgeLeUO4g0RvAQRhmqzCXHI1Xq2Q5PEnfyL8pBQJ1WgOu44W
JBH5mgWrPhuytjps+kKtCZqRE5XHzvzQFR9fMFkioIQNgzGcEmCtZJFCS5xPu07zkone+KxyK6og
ytTOVT404LzPY167zo5ZiOSfePSxJv1UrrrTlWFAnvVPHCYDkhNOdKAVirlHXw39IaKpteHNqZwp
Su1+C3pHW5OtWPkUd2AI0sGJCp2M7R7geCIJun4b+YuYEXznNpwcXCqULK3khBxMC8b1r6fb94yt
RXPSbGgV9jddUIldUgx+K0sa8iy1K6MdS0HoP/KSmeF2lr+pTVbaHiiiZd7JqHjszeb2LqE1jGna
5b1PARcuQUr0mc2HbJRv5YtXNQEJdlMP679oWADUUn28Vr5HOWV7VSl8FtVjGO4XHpFvMbY6CU2B
ccv6mrI8I50vm3il2dT6z3BekvsIqYHN8D5JVD06t6v82XIcvKIZYF13K/iMdOWOyL7XFAyofnR4
DunSsHY8AalncER0sUw3x22NYZ3lr807w1Q+lcODjLlruVKsTY63aCOCVmCvd8kVW/qmVRS47Izd
CVvIHcsa2a3cUbzaWOZASr+u9fh/ObQdCG74MPorkfGhm/5bTbQ3PtWW1vdL585Jx60tZ4aQNAFf
JaUxff1xDHiNVG9LF2Zl55oxxqwgimxWtoBhnygYqiG0dSAWqX3oDhTCzvXyZpE/eT3QSOQvMCY6
0xSWY5hj431yxctNTVzRgMLRRS/2fmMV5uRUfK8NYkXigjn4jD0axPoS3U/znuU3pC44uj0xHbOI
+fgFlLBSI+/De68dPrYxyIW8a6ajgKL3vXdz6iAysDf1t2/nqxzVdkA8vnHIBshyeMeRLHlvexMF
Zch+uUlXniRn40MjQ4aheY75jkwYQIGbzzElLJ8P0ZtGB/+1IAWdQONw9n4Kdg9X00+GhJwRlS5w
swG+d16AbJoBrc4Qv8MXBxfkPVwKWo7hH833YOp4/KdRFoHa1dcGmBIRxzRvMe536fSQ6EbROPLH
6wVc1bdnbLmcYEH33L6I8o/8StKSrRC8MWIKCcZ9L7sLV1QeI9ybJXeapLjPLt/H8+EXLf7vCAwT
nrDkNq+inQO4WP4NO/0YGMo4U47qHn5EiYLisQWEmDhcdUDTUYbHsNSTLkrAjCZ3OQgqeukQDc3D
WV/4Q8oe6IRaF2mspn3U9/Qs2yCthm7y0fcQXZoS8Nbexwpz5fHRHku1io+9aG/M46s9z0EftGAh
ahRkBZzv5BPEWulA4QFk4afddZOIgMIf/YhdbeoN20UJvDvzZmdTlNEoJlPIk6P5p5D194Ni62HJ
6Yw+GPWzH6o3X6jU1AtD2fdYg+fdP0SwW9KD1LkEGcbga5hEZx/5VkiWfnwjicWPa8MwDY8jD4Tt
H1PXkJZxXP2EYOWqnr+40G7lwltzWALeqgvpcbbzFw6cl7TFj/0uSlNBuhbC4A9FsW4sjOduPz+8
WMPEiFl3icMZzUXcL1ZDeA15VN+kA6ArplaDUgXBlDxrWYeyfNGnfJb0nwQxEgfTTFTJ5vLEaRbp
Eufpq9TV9RIKqIvJ3J5X2KnhDEiUTkb4Eg60VO4xOsDjcvrE1MWfR3RpOneKcpGbsKMQUH5CO5aM
PX/2dzwj7YkFzvhsqHVdqb3MtlkXIGAjLKuRnv0ZL/zLjrj9bplcu8cb9oj3kPZYG1b1ZaanZ+pV
ws9bTEn+/whfOOWn5cV7RZFvjLOpJbq9+JkTN9RUqp2tJ1tSXvDvUxz9Q85prtWRRO63cV+MeG83
C2WGWKAYZhILm7vKzlqIZvEgPJk0/OHOtoARnBF/yI6WCQc2iMLwiHis2DK515t8t6ZshBDi0XBx
QUP+4h/yq1NGjTEaW9Oc6TjWyg1w20FxnKNezlW9Pn7laKh/kxfchewQmgp1tRiPPHeaT4Wxdbsg
PNAP98DEPGEzPTEtvlUjDH7dEAAOW8oVy0pUY6FOpw6TaHf00WdfxTzjIJ0pKFSw1QeokW85XLU5
OToVzyTQP7w0Gctbdczg+ZtrmGrs41yddpuHf5+xsmPefLkuoKNDtYik/wksaIfxmEo4j+yogbBC
uceDdw9sGumGvupevigPLjb2Tr7firXLG4ent/QLm1ncgEw9PYBEsKS+F71OU09dUCW4pyAyzkqb
O7olcAP2g+ow/24QbQB9HLfvc1Kchh6/EnTdISNQ8mInWb4x6agK0RxAugwkF6qZ69sJmQ8FAOj5
gnnAzJvH1LLubDooosjFLkydolBTT2Gd9a0XKlvq3cpZxr0pN7WSJVd4MTJsBr0LHnWIXfBIQOF0
Oh4BAJa1q8o00+rzH159nUXImHN12APD9CgQKWPf0Y9tT/1VAidrW03b0kof2wv0QHIdJx38MtO4
/gMX8Y1+Pl/wz60G9otuXvz20mtwOyrDogGEus51bNEEwSGiuZRFdxJF2z8cmUC+5lf8r+TK98RW
s0njUI4xQX2F/v0JN4PeNZmqzH8oUX96tpoDYoIoS61/F3YekQfjazhVE28a1pNq6JE3IU07RKbL
SduS3dzEXW9C+8hspyTkg3uLRXy8Lg6LgglyqsORVsfTXbDdAXND1w//idwNnyO0hAzpoKNykcLb
SgwHS6W8kQcL4azUjPLPoT5RQoN3erL6FuNhNdGfDW4PefQ6wm+CC0gdO4RMp3VZ7PoigMya25CH
JBdNUm8eVbqvLLILEyTCe8N8+VC4Lt5T94diDYjTkVZU0/KrhREhLnB8brN3+CKzwlZBrqBb6k0r
sW6hSnA=
`protect end_protected
