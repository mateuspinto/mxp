`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`protect data_block
BlUj2nxF9o0THS2Raey2UpNZXXFYex/vuZzG0jSnlEhdJW2QezEnyT+2ZvMYIXzDqTzU4dGgdKM3
OjmBKLiMal9gQUHlCfh0sTURDNXIOq1JTeyM1Pp0lXhjmyJx0LVEye51bOxyoFaOUh5aEElciAes
Ze7VIwPr59L+r0J1Nsjes1bfTB48uey55MfGh/kKV2+IGnDls0amElRFBNhW9Gihkjp9QvICdaEL
JqQ/wD/pw68TJIso4mcm8zrnZaO5Zoo5P9S7vu6OtFSzHELNnIOFAwhw4z7oWdmaWYpPMT5mOs80
qmvp9//uqYbg/NlWR81vU7oP5GxqbzwWbGYFoBQOAk4SJ2WWAC7Och2km/8I76F5FBTx4if3EEAN
mjGCmzta++l4whrWd/A1ylsRGsQ8OPB/bToYxUG/Hw4cZ6qrDm/XtAdUJDUWtpGaA4Q3XmpOFe0x
ekwHJrH3LTYCRDV+chG+H2pBiBKfSVM+SBnziDv5GDv/VqBz88XEpd3wi3f6fmMTjHi7SlmgSapW
/7cpRLtCnhHiCtHeGA1nGtnOr2UQpSvWG5VC7YMU5bpypt1fqZ2nek3JdAk1xHsoJU+QhZZCc8aR
7TMkV9E540CrKbYKezj262ZZKHGIi2mwvpDizlvA93L98yQ4hZWMH9c9ing17arBbDR30PCJylwH
KOLRmzgyxigvcItiulTFxHxoZVjpNwtBijYetZILa/P6+t+ksrW8Emh6dz/sHNkA5TmetZsuT8jV
RHXpV0Lg4rjFRkaDze5BEvkCEeMt+MXrEMJyKLjRtUuoVZxDsI2iN612AIXVX20ogdHMHvS7b72r
Lqm519WGhoyNmukH994pN48de5Bcvm6Z95nOlXnVMZPc4kLGdMZDQX8xRGv/QUuMIrbEQC96f0jn
74hqb9dTL3dFJtWEPynRiyBS1a1gRiI2Pu2qGsSQZj3db+uPISnPZQEBmn1jgHqB9OFmTCe6HisT
sPKVhASoJTpoWSyrHIibjQf3FLNRJjX0IV46+3BtGsHuszQ7zlVDvH1sZR6yWvN5Qy14Y/Sy6qUu
00hEH7llE/eYlooSyfRsXClgKi1x+gLDch2mxvX0B3ioe1Ggwkn5vW9ZEd/wMk9Mzv3VmDKa0+cN
5rTyZBodhhcnwz93E0bZzIWDmtdvkOsG4Yo4bwYNDn2PiFSdUIkG4USoJ0Gc1Jcj+uK8Km+FBLy9
A0sKGUuju1Jrh6WneAr0ezKMmcHJvxikxLBKb07Ugz5DWg1fqIafSgc4/SXOFIv2KZj/gfl4CN2E
+NA8SokyqUSqrxrHpQXXMZEgWWadWVmfFgQooa+GsyQDBJWSay7FhvQuWY+0zKIWzm+enov3WyIa
E+leZkUeQCLItisoivCtb2gsvsrSqPJhiwIDxXwCJcd+DNaqDQ2oWeYVgUjMxZn/4CT7APzuhCZD
y+kWfWDrHh0OAJisDGTgSzsSzK6pJ/bg15MQ15n48rpGmV2/m5IOzMCo8zjVTRo8EsWsyyhayqdT
yR/0hhCxyaoTABr+LhtTrKZX+PcvX/VFqx2zSLu6w4hQ8h4eQ2xodQbX31vWy5H1qr1cgyRnCSwl
tVCby3Bnwc8yNqacBSW1E8mPnVsTNZGicBHVlWJ1Jk/MmB2SAAi5jiFMOP0AUHASee08AccozDzt
QDpnyAdShwLYrN2VZmvsi3wWsN0e+Bl2iV2C83s5FM7d5lm7j0V0D9EqvQ41Sipr8md32x7ffPsd
GmDIFAQ+WxO9nObqiSvsJeQ4yXQ8QuvVHFQBR2YxOHGVTaeEuavN0EYq9cIol0SP7KiLya9+x9c2
Y6bx9bVraPKqtG829jRKUbXOILf9RCvn3icrvQVfr8j1e61JUNvs4d98WoFvz4oGD5EX+ZgzpB7N
FZfpBiP+mAP7GJRWuZ5CvdEd4pXk7zgbD7j8DRNeRXXkahGhq8u4Tu737/wH530rbyiu03zak0Z2
+n+fy4mdndNKCvmKGLA41m152/0SrY2di5QIAw4yl1SMoxM8uekHpyftt36VVQCEHgrRo6dXTD/W
j3EcJHKsQfOszV8qAOr+eVJQ/x51wfYr7pZabUelEKCIZ2MAXorkdJPNUj23psvlK9fKERMaRyqq
3odfa9fLjDPE+NsUq8Y8ua+HeyLVWhXdWcoPxsf+bMXyhvhchJwONLXD1OOgAdpdsBRpvH+HcQeX
MsNoqmfxHvjtihh0hf7lkTuaRv3SY3uGJzw7wsGmXIsdvBkx9Do6mURAytWFg1JpaBfs/o7MVlkY
tIOlDPfNcKClpDTqYBANZHkQmM3/sX5ZeeYkuJjSJDtrUZTcBcjADiEZC4Z2sM3xP5d+NzwRhaNM
1gWn0eEMowvM29noaLvTnsOiKKIEaoKlAWuYWPCt0XCsAlM2rArn8dmibYAKmzTZmCZfWH/Fne1f
6MwXBUJZFRxxoShTqJKQR5pLocYwls9mxEsPnrjXcSS3+/qyC3USJwXv4R92Yb1ldgqff80F0Lga
1eKrU2z4UW/hIw2yn0W9HEyabUKfeBWkFIiWwzR3wg7qOV+DXTzHVj29NqhfnP7pXbGQjDnrg3Cw
xza9PzN6b7jjs8WdGZp7u5nRWACn5ccdCpFBz/G+xqib/dXNg1gAoAyssbd8TnfLJiw76S8UQ5CB
qw149xXZVFgIVSzgNZwqPxvc+794Gk/sz22Q1yKvMTodvClrZhk0B6lgFVbew2B3lAMWdRamxSNY
q0U9ZM4I8eVYT72wJa1YqpFqye1CZrTH4+fGRedjgHB4S2GC271+6GHRQAdvCn8u5sMiE3yWJ2At
ntCer+wC7iCWqnFWcQDJ+LBpGyzC5ZJahvF/d9LCIYbWMG0y20+DOC6LLPSGw9ScSLLFBhizPIxC
1hC7EQw2bcuzll6cQ2ixIy9ci+BNoej8Vi6npxR7UlZqsYluFPEGTsUQSYpM+tW/3vKp0sVu8uVy
CZS4N1varyJWcdDfsnixF0OsoostJt9gb9hHBT/zB7oszBGVCx3w4dhR36ohtVDHudpjTTtGRsnM
1FviUAVG2Oc9sB6m01UsbxkOdwGqXk/TIj1wJP7bt4cWz67P6RF2lu5xWzOjrhCjkd3spn6ssbEF
fUPUDoFFBXXs1w5zvxM1pus9Hqj8uT2RVPBh3rGbSV/IMLDsR6vzqdkJJqRTjRqMLKjKzEX1fqjM
QKnN2IJwuoUjNG/z00D2neQgPTMY3TEg1BVc+9h0mCe78NZSl7GAgKU4oTsyM91hvh7ZMQOFOyhe
PqCkrRF+il7njh4ZtF4sN3Mo8thoWHVC5+WnK6a66o0oh8RSMicxVmzjwn9DSywUHltwA5JMXQ1Y
z5J1bQXtFkdOHiWQJe3iyfwNdzHUpRpAEfkmeLL6smzrwZ0vOZFFpY+hbcWOvFLFwhupwPjnhjOa
82qyKOTOPgvGH07m9Zf5ND/5NmMzF9xsYCyqqazvWCTelz8+FLbZBzkBF3SiuI/Zcdh3EfYscAEI
nIE9d02ex2KCRlJXdiC3g+tXHDYc3l+LIhh8cbTratlXzMc0MCCvbO1FTTkWRWZsKF7ivmLBVSNF
O7aLtd4y2fgBFqcLBnKrSkm94NW+nPnEmMz90okcNmHG1BPTyppKXPdhaaxNAJCtudLX8J5DqwC+
z+Jay+pa7udbOBT+thNmdD9Nlvbk1nFtpJsh/SgMCwMw71dTuvw+JLzkPS3GHAUdUHm/bFzuJyeL
g5pzkANrshUCDP2wCJIIRjlXtILE4kPc67IAlT9JzeRQ9Lbs0s+0tTA/PjZL3AVcoBtoOB0e3yQa
KZej+ELgCqW52QzlduZ2X+N4hFU7zeA1JwfkhKnnTONH3fOUnpL2rKe7ZguFlf9XRm/wmzRSo+45
mf06iXHTzyyUx+BfZkW5w4mtVO9yFNPHdC497YcqcDhLKegjYkzu3WYV4ges+l1EGbbDAM2W/sSn
Pz7jtbRoa3h7j5aZs96jDVmE0gFEFL8d1bTWMfQpFavFxZ6HxwdjaoZsSi+9gn4++7SsKRkvQHor
CtXylTOF/bKDmZ86TJo7DHUB0Oto6NKTOcVmL7uBGtCAzCurnwq9KFckYF93D5G9H09NIS31Qj9S
gVBbAyiUpguOWW16ao09MruEiueOGddqv81ueqCi3U7ZuwiWHoHGSEGzVvOjNLGf5rrgMzotdb9i
pft6/RMaFF2ENYtlv3qf9bKK/wCzXiJgpvpZKk8yJ95qwR4FGVQDlEaJpKfXkjlOcdVdXzj6UF0d
w8m/1O7k43rcZM8CduTqDbbt4V6WET3sSB71b7EhSWuVPkSlZy/Mt9p37zyuh3ShnRHAIzNQbp5N
27iQqxfpIZfiDrL+qSdpdE5ZXf8YYQ83gKHf0Ol9xUQ7ibPU/zdUptGWmqW46fpmTkyvPrzoGlaa
6O1J/M03zCOGJlyy543gg/oXKGQ4lecwMaJ6Cbcam62E9ITtZyjGA0LfhZUnEnYZt8IyUpB+b80b
tMFGWpPcZQxa0EBaLHz4fyxkNcDUeCFLTVMsCBbCQ4wtTzyc4B18o3FnLdROg0VExbFu4P3rS8Ym
kOAqpONrnUwaCxrWZdyteUON/BPABRIrMLf5e1bjFdTS79UsYfLyuj6YLpFb3qfsm4x+vXCPLOiO
ymgpMdljACW6zWFkWwqG4qYr5JbHRQ6Stheq
`protect end_protected
