XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����J*K ޸����ʅ�UR�`B�v��`��R�d��� ��fr��pM>C^�4�E�֬o ,�ʉ���Ⱪ ��L��N��C?��)�<��o^}d<���aK�=Q�%Li�D�4�ѷ$��O��
{u:�q�!��s���ꠘ\Ÿ�qFV&:b=��[GK`G�|qYЇ"^W��N^0��Zb=��9+X���	�M2����4��h�b�p�Y=#�z�0�o6J���b c�.KBA>��g\eƊ�O��K;M}}7 �N�m�M�m�c�ی��5���㷳�
�>\$��6w;%{ EY�8n7�R��{`<~�;K�v������.���%%4���H�1<�4��veb!6.�=�ֻ�bhN-���@����)�trin��\��T�-q�M���IB0�[�j���T�L����O9�s$�"� s��c�3B��.���P:�b���W.��w��uW��9��>e��(��tY1侱,5�!���K�{Dk���߿��ű��o���_W�"qfY���^�1�.~s6���{��qqj��8����o�'�M�[�V�k�>%.�ݔ�n��|^^�7���b���hj}��n6��4������Ϳ�D7Q��N�`n�7r�̀g��6������Z��}�����T��*��6Xǌ�0�,�hz�݀�	*7���pʳ�H⃉���X�)��f?0pJ3�l���%+���&0�$A�UwD��h�b��a/�f=XlxVHYEB     400     1d0Ė�� �-�o�K��)l��q���p^��i9h����ޫwJ^?8=�:��m^�� `���r��%��C�r~�IUe�?5A��)0�::Y~�`3d50~��5 G!�#���8d�uQ���"RX�ekΗ$.<U�*��*��w]|:ع��_��,���TW�X:9R>�j��B�;� �`�_�۽����JP�N U�o���j�XV��q�N�B�"�~�J�kϊ-j}�༹�
�U�w��{���w���}�����Q����t<V�#Kx����ݐ8���E�����U"F:�!Q)Ҡ;�����!�����!f0��� A�1pq<�v�A�*��"�䞳����9����>]B7^4��S�@������̸z�#� )�T"ڮ���y_�-�*�:�����ʋ1ض�/rX�����6�6RVv����I�HdJXfT	\X+��dX����K�4�XlxVHYEB     400     160�(#$,,nU"���dfN]�0�������-\G����i�3JC��{��Pÿ�～��0 wW|�S:)�6]Fj�z<%�2������X�|�{�w���3���:�춥9BwW+�� 6E	&)�	p^qxҖJ*+ F��
��b�>ʿ�	��_k@ �#Ks���YeG��]v�1�4�@�E�r��ksy)���镸��,Z[�T�w<\�r�	r���Z�Kr��9��>���J^�vё�����ע׽����bڴ����@�N��3:��T�B�iV8��Л�4��k�Жj����5����eU��x���xJ�J;eZ��nl�f}�2������1KXlxVHYEB     400     110��݅w~�����������2��	��\E;�H�i��nG�5�П��B����� ���,�f�����So���W��&�q"��]8oм����u�ل�JA��I���5r/0�����R�zW �� �I.�"��[Š����9`�Ź(4�K����	#x�[~�q��j��ݵ!���d�Vj=��T������|�aw��b[�_ȿ_)7>�h1G���c	r7�Z|��T�g⚯[�	���	��P��w�pݱ�����\i}�˅��XlxVHYEB     400     110��Zg�?nx)_\�Juey�A=���p#܍ �F3��]����-��	��J����'�a �`�	��B��D	�-:��Z�ƻU�^hvU�?��tI���ҭuW�6+q��u�#Z�U��`���N�I�����p�3�b_�����4���������/��.��[��񤒰R�#�tąG3��AV}\`|�3~�+�1J���#E��4X;���U^��=��%�q</jD��a�~=0/�n��􍎨bmEMi?�}����GHd�XlxVHYEB     400     150�m�Ր2�;U��\&A\���!R����(��e/�K�qgZ2�T#��xTj�������)��$ԃ�>Z�@��#*�O�� Jѷa���2?b��;Ww��r�K��R���ɉ�7 j���z	��L�W�R2	���K9<2E��_=^_I�$'���ǰ�6I(BTB�TF�F�̱'����fG�Urf��cL����ʕJG� ��4Z�|h߳�I� K�ĴA_�����E���m)L$ֳ��}/�ܰU�5��8Czv�|�d�k[X^S�E�8 �ى{U�{"|��D�x��4�?��}��-0�0Qް��v��+f�6�_'�lܷ#�XlxVHYEB     400     190�8OsI�Qz �hR?��p.w.�zY֒�?��aV��EhA ���/5s3 	rr��$%-�̣|��B��v�Q���RkY�m��v~2�s+���M�y@���P,������2��dE�QG��_���}�\���t�5X��W�F��$��p3�$�n�A��J;��p��&� ����<��3���F��B��d���ˍA/��|�P�sy����p��� &�ي�p�&��^�� ��a͸�O�_C�#aiq���v���P�-&g���B3�y�E��1Q+g�b}�$��2�I�@uT���pԈV{}�3D�?7��`��]!�.gI��G�zRn4҉���Nچr��L��f���!i1$1(~�:�x�Fk�^�PT�u&&�W,�8$�H�������XlxVHYEB     400     150�n�'0Lgf?Z)g5�ggᓩ٦�A�5o��5Rp"�GS�h�d ��^+J?=S����^K>�#*�b�I��g��<9;�%~(���'箌�#xz42�>s�����Qq|(Z*9��	�u�+Z���g�o'$u�윈&ֵ0ރ��b�==���pB��m����.�%��1��|��-m� �����kWF/�GL7s����gy��z����A��WȘϗ��]
�9�O�8V�bX	Z:�	��N��,��"�7g��m�l}�ڗu��V� U@���g;}is�!@�ɧ���!z�f7N%��]���o�H�^������K9�b��O⎍�XlxVHYEB     400     160�A���{$u�סb*q��P��2�9�-fɵ�����Ҿ�fZ��x��p?�";n�z�51c|�Qsw���#q�q��m��/�g�+�t�=L+� ��A9�B�Ʒ���)�d� � k:j1X�=EM�.x�:](k�����r;!�i04���Ȇ���ޘ�-��Q�3z��~�R2���������`�5ߔA���I;���Iފ���ؗllF_yU\��3�%��'��0ղ�B�Q:d�%��x݃�.�0͞�Ft�k�g��^'ֲ���!8&?�����b�#�-��җ��q��EG"�p�4ލo��n��F��`����ԑ\~�v�����\�u��\XlxVHYEB     400     120�|3��=�N��h�����t��6v;�KE6����9j�hL{���N7���%y���Akv�li�u�PE!�(f�WM��^(�I
(�|����È�$�D-��>�ү~t�\!\�}��~)��n-� M��RL�uu���i�"6���"���g���P���c�ѻbV������'��rM筴�MxOc�/��a��D�'wt[��1��I����m�������^�ǧQ�z��!��ފ�w�w��ߕO�.1S�Gk����� ��t�oz�L�TAg���9XlxVHYEB     400     1b0{̕fED���Ȟ����t#�e6��w2��q�ǺԿ��&��u� �\�jdZG���}���ꑤ�c1���]��΅~a@����}���� �U��g�m0mN�P�����7�H������S�I�y�'�c������kH	!:TN�`Z�����*U�=B�g�r"��0`�h]�q��\
�Df-��1�)K`|߂����cN��́N�Y{D3��}���}��C���5B>��D�hĵ�������Zǈ	���ʟ��NU��7 ���ǪO�s�yٜ�\�|�ܷ/��@U��3E���Ėt9���%i��Z�i�Ҫ�Fzc�!kOV��Sj$L�7�-��8���� .���[[V5Ds�@>ѻZ�8���G�@7�z������r	H���Тg�gِo��rp��W��3j��XlxVHYEB     400     1b0��ΦB�'���geiF�V�� ��n~s�I���'m�2 �&�1˹�6l�DE��c:�<�ܣ�to#�I�`�[ӻuD�s{�]f?���x�� ��%?@N�ex�*�sܖ��E���yȊ�Ԛ���-X�d�(#��5����
'���n����3���Ļ�9�y1򂓾�(�w�-�$���,'9!�K�-� �EeF_�,Q�p�sp_��VV��̄�Pc0���"❩���<YE�;��US�A��T��3�_�K�Uf��e����?U�ڠ?t��o�Y F�f��!�-X�A@.���*}���u�'�k����;��vl����9�U��@�ηH�K#!C��&Hq����_���#-��ڋ�5{[P)�o>�
ҋ�
^����x�w�Rf[۝i�D��:����̈́���{�21�U�m2S톢��g 6XlxVHYEB     400     180"`b��/U1(N�g�+��mI������O��@����c<Mjڧ��IFS�itT$�{t�?�X���?�H�/�.6JnAW��u�+��� �'����M�`�b����~#���pS4�M���I������-���-~�ǉ�P��������"
�]픷%�*�E�UV��\v��o���}'��u<��t���9%�?B2	K���v�	
�ј-%[� ;꫿�R�����T�>�;�������0�o��`��[�Ҷ��2�?Z¯">�+¦��u���G{,ej�]b��w�ߝ32�N�O2�!�-��f%�	��@�
w�gC�/5l�!Z��Z"X2{ٰ���������m�X���h�^�)_�ݣ_/S��XlxVHYEB     400     170��d Oa	�ռv��x���y���#5;g�ՠ�?O:�[�y�^��f{���!�
�!������zR���VH������S|FP��C)�|�\�uB�0��qR���B��N(;ܙ�M��'��������j˥W^�O����Q
�dHL�V��*"�bs���gS��I�A�Ӓm�l-�71{��>�c� ۋ 3GvI��J]�U^Ǔ�6H�ZbӲ�z
��%�o���
sH�n�V�*|�ٮ�K�f\-8��#ռ�H6��a?y��G�(�|
��r�tj:�A?����0��2��Ƒ�F�7�xX�w'K7��؊��x���W����1�� �N��#F�&>`����Z�XlxVHYEB     243     100;዁����\��������[���x� \$�7��Y2��tz�}���S25:��G��>�KD�B���-��}���
�\D���c��T����E'�b��X��ɾ��*?7� �c�p`=e��*�Zc�WX)ĭ��$0�f͑SR���P�y+ٖ� �)���`1��op[~Z�,N��f�{�����ql�$�B����R�N��&��V�A�(�[?������
6ϨJF�����f��U$d��ד��