`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
kmXk7fi/6yZ07IomIcZWu7ChLSyxleYzty0HUR65P5gJdqb//Cv1DbjemQ9Oe6q3dPBeVy0KFAPv
z4dupCf9HTXPYlOKsls3Es/jJtJqILVl3EHSDzTkHg0kuzDSX6dtPjwBiM2Niyw7KYOC/QfK1ZjR
hIw1ziQgbUeRvvloiC2Y7SUaJOt5SjepNnWnHglaa4ziUF9FHJHiHcy1b26qrCqQjIdNOhITlYq4
mH1Vpuh7LZD+0NOA29o1PxCKnko1ED3/oQlCqyk3LvNWBu0QH0b95wF315E7n0iL+oxz529PsJKX
/9n8yrd74Kpn4Zy+HB1G2DGfRLqltnZycnoC3Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="VjMrts+G36mlfVSAFDdFA3haKyvYORdai/Lh4ezvS+w="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3840)
`protect data_block
Or2tI5XeJ+didi3rhxT4S5rRxfuyjDAaba64seo+vPg8VXi+Fw17nMCTClD0Oqsra6TZ1Pr4sicD
yTTUF6rYrVyUu6CFAWrMHf2TeRUS4IOPS0fuXA1Rz4ePbRJ4qYTKEBItB19hb0nPDstYFmZIExbR
HO1k4z/F/3FF0tv+sZ6AjreLm1YseVOQbD77dSV8vdeKZa8ZsDo8/bSwSgEHYBkSoi1axkLaq2EL
6EbnhNGV4OHv+YTbkGlTDB53EQXQhc9KZ4zlaRkeFc382REGkj0L7B2CkNHK3uZvQ/IUTq4AvNe/
TJ6G4ZPewwimN+4NxYOKFb8IU7igYJuKMPKAV7K0x+1bDCIzoqbkdCXt8GN5Yf/4f/odpe158DGt
IqIN1jMWmqUFVh0mxv4ezCCQ1G/0WIX8mGjJNvCIvLj8Y+RLd+vVDYvqUD7UC9eI1M6keo8CpZAJ
9CbjJzK1GvNIOyOnwL2xIELAzxocd/b86kCGkUbu3RQimzMq/B3RHaCv6kxnSdDU5P6wAROWD7fX
bclimexCdutsy8cY2huJblMH/08CAgqSCVhQm7tew6xSbIVie20vFssHC2iSC5MvryhQl6Ymwa69
htbdjhsuiT4NzjZPMXuqbmwLDmovxaTeEoGldjJFNn6XENyYqy425ZuQL6C45mQbm2rF/2DhnbNB
eCsDvrALeFWH+MEGjB2q1Di1Qf18SviI6bh3wBw4e/UboYCGRvoWpLG8snZItAgAHi7e4bo7OCs0
+exRX4AQNINJk1Q+n4iX8sASI+f4bhYhLIkYL2PksyRS+HEdSI5u7nvYkzzkiB65eGQWon+smw0u
0xTtlExsbDBaFpuqsHZqj17bEW4oT3OMUdoShKdw1azDZ1oNHK3GeWgaEMZ3MNx5iAfv1ffbxT3v
kMyEvvtfwI6Q7US4EPGHapXluR/wJRjmdKqZTTQ4L0YmuxIvPZTN0iOr3CDFZi5OznGKy69yKxxG
3zFvOC5nBU7JZs8iC2QoTVUw/sNNrsGKZN+2x3ynfHRvV6Zoj2bLjdPr1pIHA+TxadkrJl9PKum+
6XYEe+9PTLyZkIHpxyweu2hWb2NTd0FvKz6olfbX/TfbTjCnmdvsBiStuGUxhmSqLjIHDzBRE8NT
uuYz2xUSCjwzD2JiTvIZ2QYBFWGfF422uJAWStPgF2BWblVf2KpTIEKK0ycLuTxEZrpq0m5o/BR0
Sud6SMN2rkew7pxk49ugUjTT5czrM8C/3s+FVmqcoT60zvCdkw19fo69kAMrWxyaGIZ3a09modgE
R02/rfwcr2DdbZK+Du9nFRQOUN15LVabOsViDroz3P/3+6tQQPSfKP+wj3HUsmjv7Ez+EE8UPu/z
caGtvZbT/9MhrdnBfR2BWMNb+r5Rc9cR7MTpy9E1FIriAFX6d1+vvI7vHpv/MmXXYolpwxGGT68B
+uUINjWCUAkp18wecdPS5hRJNyvomEXVvHLSK133UYqb13sWwXXGzcsfy+rY2p2W9RDrwj8OgDWX
6nRuqHUDi9gS6ypKGKi4ZmmdJAH7cP0i0CjNSOwEZy4Q6r3hfPRXb9t6RTH2IVmEAe0gaMGsYx0Q
tACrVf1u/lTsT+9bpBqgHHQN0ddEMGuk2mKt5+eys4i1NXR/XJKH7eVkdc2Uk8WYSX+EVZV7kgwI
GC3TJGP01ISsf6Asybu5t9caYHECTk3pWixBFeIP7rJuhgggpEoy+V+xKCD45wJpP+VbjR3jOiUf
TjaHHxvQJeecHaCXhtZubtaOTK6dr5j+gvcoe82lQ6hhdtIkCdyzCwI9WmqaPGttuavS2YkSx0OV
B5vL0XRG3ITRS05e6psA1CvcGdJ9JfGwhy3shMKL39U4SUxEifvCUKIvpFBFRytC7o5eRoy+ehu1
a5aPIuogZTNQjxrjtaXRgIiUOzAo1tzvCz+3ygSKDh1m7U+eK0CxT3rx83qzBhk3r80NYHYwvdyt
2xPaTFcRZxVXcz3cNwJ4B74ciNUJ1gsYNC0FqKPy2d7vqUv3vbn2jO5bwBMFSxa0ynVcWx/JtWBN
WDHHcnP1Vg78mhyWNIEI8QnCk/Q/npwCt/HfwsEyrvxTPl00fArhYPGsgN1WE4qXZJaybw8ocOKn
My/ruRsbloPdchlNPdoP9nWd4CoIpR00+93JMHL/7q9uGs5/KWsbk/XD0FQAHXHEF1sFMiujA3y/
lmcv/5Md+7fxW4o+Sy8BMxmd7m+d0QCgtl3gnNyANRSEFdhKm/gd8fQqwvVPkmWnBfwr7/Jcwyb9
vKoQIPNqHnUQZW2BrbsSzarKlFkZpPzS94INvY6KEJJyzcytVUgm/TiLwpcFA+sWyKCCzugLV1Y/
MZOqOXHy1IRBjcbOQ+tJJqOXpW8qM0RUW8LWt2aGJ2lApowL2Ln9YLcFWDgg4oNKo29fXORmixXw
CZ/OrLdFudrszg373K89vaSvvYPG18QxzBl4zGAyhAi5XIw0MVtXlCmr2PryHbE9uGp4YK6R5cUS
k/p+egi6ikR+YBWjZ5rf+88jvYnhGx5J81W/GMZJDpcJ3OB3EwkzZ5dk/PiVVWeCTgQ7WcgJX+Tr
G0aCBtKzp8rbvl8OsnMcXYeeIhIzrum3m6shCgpX+O4SjpmW9p0lT1SDimCCyXthin+rzBRhGbNT
UEiCrTa76UZbJSzsDR5axSmv07d4yjJPj5nRnr0c6BYfIzf4FpjxuG57/81LSLra06YT0kmyZJZB
BSxA88N1FGMlKWbu724eRJHsQKn+PKqdt+GocR1va2Q6pii2Hp/cxdebg1eC+t35YAZZSWQHuXkZ
9s/gFHeeewMmo/l1Z0p5d0xJQYgEqAwE9R5hS6wmYZ96CFw3JZHF+Br6hQq9/4iF9YXgTeZ7Qx25
8NDql+KtAb+ilVcUqmW00WiJ+zbM1uao4LsI6TUGo92Y13HbW0xfECDbCx0EnTiFEK7cU4upBiC0
Wf4a6cQBcXIbF5Q3NsC+KRTBWplm+93TjFToY2zia9tGGPxZ9K1MWu978wd5YuqfCrfoVQ40x1us
/TKjxDCY+9omA8vrX6aVtY69rcRz93U5DqvNeJLUr6Edsp3kJrr1NZDqpOgfOzPDBboT5kh93S9S
NKo7pJ1qsGMj7GHlZK9EI+bVk3beAPatULrf057rw7Z/q40mS7+sI86tBvnxGuHqXPGDYjrwpviW
ffEie5NVkWbOVjO1tcpaTlKtPoVZLk5VKY0WxO6y8TfzaBQnilwWRUqfx3O6biuAi+eEnv3op54a
ZesXQXUzXMntwCfvZLIfVkiHPKd0UbDdq7DlWk1+YOHk1IQ+VoDFafArydEi5N37JkXv0dSpJlMZ
uHQOqFOeS5MPe7IO2OuF351+lsEISNG9bRo5GNaHoDLx9CRlN22DZWbI4I2obXbU00GrIUw/94+Y
XayEApjuSBufSyQHWbtfaosYVrVoKOgSORC9PUKELyo4d3MFcDcOSFE1bAsxSo1Wb3R/+R1e2vok
/7JcPW2ogEQotD1MrgUHwFH6HgnUlOoKyNysCfNIAlW6IiqdPLRP+1r5Qa0Jqy861B0bUrhxFclj
ptjVMRM3MclaMEsb/jBixoHPhOnEhJbW/byAPmyBG69h4d6ySKiAqMct8GvXjP08sv7XYpV1zJD1
6TifWArWKl+f1m9pg0UUEbUQ+F23wh1+Wq55NFVnbqbJO1GdRJEAxQAtAdxt0ri/5WKY4uBkzDii
5ChOt/vvkXFXNBvQvHKw+p/oXM9uudZs8SHN+hvacHxSegIIqTlsdmVHSdEuk9ZZmzEl8EQ2yp1G
KbqweKO26RZ3bM8IK3r8Ha8IgObqr2NKOjH5CFDq7MhaQku80ARZ0dfop35RqkuFBk41NAow3+m6
c32x/Y7iCEuPe82NE4o9kj8+3heIT9lA0X6ZgU1fRcQmT+yPC8+hHFIaR7fpy4s0uV3hREjqLHim
musPK4DXL6AyB9+dmlO5DgufHcEo2i4MpQllvWCHtLCSYuGmsZuxj11rUSpEYGfJIlvVk2MsQij6
3a4B2cerh0iEI+H8JKIGbYiL/xXQS5Q7z4/18encLYH8qrEG17C1rOglmBHdG/ZF/1pcVgK5gbtz
FWFDzcX4p/YaMCuJTV2zMQeRwC1Km2hQ/WMreJwIh9/QJWzKLi1eHgle51MeW1lQdLXzBTa8tryq
72Ug0+rkez4vh5F164tdIyQo7Z7tHVkBeCYvBt0A59jsfMnHPOZGkH/uMkEXzyanauwWmJh3akDg
9sYUwsIflgkKELNJrqwdjeMtQNK37RhMCAEohxut5AiNU0pHzeB33Sq/NAKRpCn7GLWQJuLb27Fg
FGGvnqfkjjAzNGYWMfTqm97r2evT8ZitoKjp3ovKQNHH+68t05EAJjoCEPrnNZ3R5NCAq+PzZ9Gj
EfV7T9L54HT6G+bHoVEmdBudmoiqIYO2ILYYff3zJIeZ5brG2aVSM9H5djuqQEcbVH9Ap0IpKHDB
cvqm9fijzEXtC2tjEnVdfBjTPa97RhuYGxmf3SzWqyJhkjgecXIPA8dScFZQISuJ4rB3UIa1nIDN
ZZ6o4XBVn0nT8PEPvHo9NkP/co85H55ySfcseUlezXR8awmtYO2//pm5Pl9uQFSJTo5/EGzAyJSz
EN6wWYIUtleOtn5dDE6Zx5UakiVh6HTsg4yN5+ekFSBnrVL7g7qM0SJUblgxPx3vO6olkoLV45Rb
Vfz05pdoLF7TSmuUt2OHOxnvz/0/lk5WddIkKFX2Qai9nwohLM5DVr9dQsxqHYTc9ODRQW3NaiQb
EJBSOK1cA5oQFB4rTGFLl/xQXrasJfvmrPbyXZlt2QMqZszP0A4IUWy0qKt1OKwNCL0/IMFzTqbP
PoO80/ZGvK98qiFLWA1N61hIr8+RlafFtfBxPFckAh4aC+0FBGBBoY0M5JP0ZtBQ+SXcS2NX56qU
WCa0O4d14lx1OKa5cziOvM391YeEc9CYuHaJdsdsQCwL29t63rW0g7S6lnmYWGYSD/BaPpXUmdr7
MnsQaNio7ft8gYOY/KnCpPqHK2QWMNfkYV5NPfVTawhytqjuUfz4JSU8l5ebzvkJrPDyLiazff76
Y4ClYqnEYp1HYKDhxIjS3i5SFKUZ
`protect end_protected
