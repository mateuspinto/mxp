`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
ezYt6Ulls7c61KVpglIvAVe/MWz/LofW+TuFy1PW91k5ipP4bLQsyEatzsNOzRRv5r//TbMakFUI
WBw0erklNiFIKHsRND+Nib1+FkypUNBrfUP3/OI/Os/tluGb8UHDyWk6cZRWrwmEI+3csdp5l820
CD+AU7kjC0naJESaJkIVPw30wrYxgK+/JlK2ulGZbETRKI1gI3QrtifA2Ki8OdWeEkS46mtbt5Yd
3TW9rC3rfmb/+j/lQb9JMH1aK+VAAnuUc11oT0VVQceVLxSUHCKZPDKiUg9eKmXC+woxUh+8XC2x
iTV2K3GV64aJ1ECIjH/n8DGkWy8Z9Vq34dfD+g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="NF+/uasdHVUfaQGpIE46n9fn4hZFcw/gvubT3/G3/84="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2800)
`protect data_block
3SxgX/k3Yt//mXABdl9sZaLua/Ef5mTNbfEZJO4TcAESdvHVDVxx/Tn2Ol3V5brVouzmRf/fahqd
tsAn3L+U+YHas4Dscy2NipUfw3iaxpfFBc5RUzP2d8q9JUnT2bVeWIvtxlcN+O5syLHeRY+fVUpP
4opdtBegQxqqlSXRmIhpVFxZaOKUescJsBjW1Rj4aN+Y2Y5n8yHjwbb2koh6g+rESP+k8iqjUnSV
UOCH5nJJnb4v+h3bxP/4GxlFu+eJ5haqGec9n4nyTe4DUZFrfyeC4tOFK1Y6eXTAmceSthSVqqfN
2aoMLXZxx1q17F0qL7mfK3lEf5ZZTLI2KG2tdDiHEsBkJFhS0ijQl3GuFUPwWj7mYrQnHhjrpNTb
c18yKRASy4AkWL/Tge29XP0jlj+oORB98XcDisb9YS7HjQS54h+K5FUaCS5RFQZlaLZ4t3OJx1v9
QecAP2d1kVNl/8c+7Dkfrs4uJEKD24AL+j+07dD622V3gvCgOr6Kth0KDCLfJ4OagyhSeGfbR37C
soXqCJrhewl8dQbhjeNsrImf6ZXHpgrci/IztK0QvL641wyDLdk8SmiZnpnHUcmX4hCgw0h4YhwC
atuK9Bx/LIwAe4IJT4kvHGQNLaRxzbEDAFuXU/jXJQUvfNKuuailPePIRgkkfWl+PVm9xhPp0DAR
Gu9Bda0Wt8bq4g5kJ2SgekuYJUdmQx7aPkEfFoaDotttbyWZ2BhyglOytnbZG5+96q0S0u7RHtcW
v/WxchTkUs7WpB+BmKKXNUYYGlcf9a4+57Okf15pnuToGW1hw/uZZIY9rTss37muGFN5DbRTUm6B
W+wNmvAzQkD7ZXORi+dZ/Ud9lmMWW8TUVHCEx/OiF1KjhEqPfUAhMWnArmFOuxXbwrhnChBPBAOC
CF4HScFezwUD2hmWaKgmQe0+W8cAFvRcCO93lwgpKAWHgsKcjDegnbZ3CMxExeMWcpxO44YLP85n
E6gVdi2yj23QsAIxSpwnPq+Z1vgXy2PlnDOaBY/Iwtb4Y7c1qMAj2+Qo2SyimiSnZMk6r6hrwxH3
H4kCPC0iP9xew0iQ0S9G4HW/KtaetRkZT2STQapA92bgG1smC8a796psk3GXU5+z7WMSGkrHQ+s9
aNmEwLerUxwbLQkYMwzJth5cdZVyBMHKNs57JDqeTtrQnjp7Y8YgU0kXP8qiPP9rvJ3rr+bkDb8F
37CvlttY+tgL1PW4fUBn1l7hcDyW95lEiU9YNo00/T03AxZ4e1CJ4p5iSjn+4OI9xIkg/bQKxIMG
Wgj5OYZRD8FjJa9E+l0Gt7tUfCK7aiM+OoEU5QUyVubhdkygDZ3Y1Fa89kHPcT0CJJTsflS4g8ZN
NBs1u0HI/H5lzLep2U6uZXTYZUxkumWJweSRU63PX6n8llU8ZsoLPzjD9qBS0zqJIeqPGOD+9UgS
l1WRlmkTL+cW2d9y+eg7KHCBquc+NImabV7TMdNY8Bn4xIFelygHKia2awdx1Nv4LJZIaN+MtACn
PWeMmhQKLOBjvanIdwzF2vIfeJ0zL1EIVtcp4bkzEzfEtkyIfmUIl0LW9w503y3YOuyQJzzFgMDJ
Sfbm4cOFL9kH4Sd0jX2uSqWQ7v5pElL0AmZ4U7jw8n8JBF6uAGL7zXAiOfad7At0Zq62mlnONk6q
Kx6VPXOSOTovSz4j1mFBxBSYk5vj0gPTytduS2QmO2JLOoHcow9KyB0GdVBBp7Vf6ghDrSgfFwqM
+PoCf5J1ey3agDz92kt8mPGWml6qxkvv7TI/NQaVrrLoMe1CFX0by5JzHjs75fYIITbRuF1eNvaQ
CMd356GC9liaRJSXCnj0t8KK/U8kglKz7Lf/449RWbvUPWfdLWimV4XSRo6GOEwq7o83N9T7+d/M
l6aikUewYKRFG6NyJQW7SHnmAFExdUJ82hj/5A0d8RnRFE2sQggKWSyUVt61EwwRIebwap6/Rjgr
gv0DtDAdzhQQIi95q3aHwNts2+7WSUID8ZoGQYMUIjvHm5SpQTjjBseLl5pF8oNfej+sPBg61Y72
MiuKHFSqW2tPi4mk4a+/+qKBwkHXqhSqGmL/wp9XBbbPBrnE3XTlp3KkfKBLFSoZl3hQG1aXFTVS
q1/bZ/QtTLsPxgSausgPpjNfEWDVL9b5aGgqT6Xwxaiw5KfYUMb4RkNiBdG9To3oCsvXzpvdTLHI
oQcXf2u9F+O70W/p5iVpfe7dg4P7fGdBcHYrf/JtDR2fw46DoiNZxrzNIEY1DKD1aaN2SpAvHfBi
BVvuv6gYIV9Ssw6AjSHZ9Hictqx1iUo+qTNc/9nuK9Cn075e8aUe2hivwtJ4Rk9qRym1TjdkNCx8
KGj36+Yz3cDaDKlSJU3t8c6wq3XXLY5OxpxYo3VdcWLWcNxAU1f/rA7m6yDwWGcFSSRM2rDA8YQJ
rAJfqHjO3KPMgOlUGpQlpkSXVFtFxs9q0s3bWES+nY65NXSlRHOK9ZAHu7RWs2TbleJGsGya17yW
PrPp3ocAVigLtB1eDFmH4K7zkgHZbgyIFRt5P0gP9b4GAF/D3T+yY/wGoAi8xFHR3AnNT4fGQag4
IjvAEs8PSdp10Gekr5j4q1IjxpGt4yOd7+ABUl0uCyb7cWhjxTDO8gRIl95uUBkNBcOzLSDUb72B
jR/PiqSG5PKJdZOiUTsjYHNdlw9Vfa4dvdwn8x6736OJUqO9p4QgJm53XAHbFlZd2EJoPZftFx07
Ik6JwBacXj7TeH2tQWBLn87aDQxv9F84nXAX5j8gWT6fdAnuPSWO9UZ3tiTMp5n3UNEMJ4hGhda/
TrlvNj7i0TaFXXQM7Dnpk6drEUuhkelqX65pPESxiTn5SxOOBOACPKgE/Hi5zpBOe14MpDcBuhIp
RWvFIAU83MH3dCbIWZkwTKR1ZXWnAOb6F8xpxr6uXWwyBBuNy8flZtS+tTlxlrf8gdQzgkTPGTnE
AN77kudrUshGwpZICXo0dheNTLGb7MgElPu0ld7ASrQSeshICcn/MKnRfvegzCLvBpK08Og9oRho
AOfBK5QtdWhtBQUBoJPqpJDqGcqio5mhTlv+aagtKaZUgYXQV1xr4+NqHRlutu/e6dBfY0Q9CBgS
unwciFJ+yNb1v+QCgdWTNalL1sgdPCsyTUYG69ng5yZ7MVdhZxvZgHo8ztQ1LVdqxN6lLWYP1A40
pwKhJjrfCfDyo9zea3MQUiZUTaH22q7yGugefV3vsPIAr3OBjV9UL3PqX7eUj3Pv7yP+aD4iR84v
2wRoTlm8ihMVV3dHuVdIfsNCoapK0L4qpc28ff3zPVXaWQUZpokTLGR8N0qx8qRXclqEuvauDTsh
5ustQGNW5jEsQQuOqtXBy2qUPTIhhhhQS7Aui0W7XZjCN1yACq+hRXpOawUwQD3UufkLyn+u2kkg
TTnE7z8dEXVSMNeCZgrIuW78nSXQ7B//vJeiZpWI5NQliyl7O79eQZmRBfsM5fb0cXJOLVstk4Td
ECJf+NY6HBQWS+8lgYUAmOhTtPKhR+tMIOrsY0BBuVnzHHa1gw0t9vfJFUtMWA73IrvpyT+HbXxp
2zhO6VJfU0pQQe1nF78RqajhizhAqMnAyrecKiVVzcwd1AJ/adxGtVNorVkohdyLnqbyqNIKupH+
xglNYGfcRhQZKGpP0IKEoPR7kH9xkp8o0BZvZqnRa45OrNCeIPrkWzhdlyZA9qu4/ih5YjNJ1R9Q
lKWkb0zGFw==
`protect end_protected
