XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��+8PT�<d��'�o��zkF�S]5b�!�w\�S�E��������?�5�J�=�� 0��ʌB`����<�&����ɵ���xV�`�t�����Ƙ���~L�08�e }w�$���ѥ	�9��m�XU����8�SU�V��mOڀ���3����p]-\Փ�3�í���ؽ����fp��>vA:m��I�'< t�~� �
�dƋ9�®-�k+��b�Sp�����=0.y�������ɋ�Kz7��_��+��u���Nt��
�e;]l5�a������gc�|SSioM**���j����;Zӗ�ϰ����8�����E��\�,�JZ�;=�_�A-���էp켪�����>0|L�L Rg+��=��AE�51V1������a�qx薷>|���{�*���/�T{�����忙���x���h6Y�b<�4�� v�����f%�8��0�F�ʀ��n��xu�+�����2��?�IɄ�S4��񍁡�ӡPU���^��am����rL��A2����Y��&6�.�W;���s#<Y	��) F���?�$��#H��e�t����d��
W&�S����'���	��Ѹq^"���̕�6��w�)B��6	k@�c�л��:?%6B��������WP��'uO��Ϩ�(E��G��6��#����	�t�e���6���s9f�阀��}�R&��5 ��r�4��#Nkʳg}��XlxVHYEB     400     210Z�-Ue��7a��^Zm=���\���Ҹ�S	=3���j�������iAA`��#<m�����Dh��<�;ŀx��{^�`m<Q!q��h��Ո�#���� ���YNX�72�5w��H�u��7����?F��j�]I��1Q�2�Eu�Q�}�� ���TL:�u8��^ix
h2��y��Q!�)e��A�4���F��z$�f�k�}>&s��1�%���x��T#�β�\����L��GmF܈	x�!J��
A�Q��ʀ�9�tl: �q\�:
�5[�=\/ ��/
�7p�y���T�6Z%.gGظ���FE�X�q.N�"�D$S�ߗ���J$�k]~j�Q2��ּ&@���'K�<nSbZ���Tt�xi�Q�.F����>��S� $ÑCd�'j���x�8빖uM�0������u�(B� �*��ӅF���d����d�x"��G����;���x�b7K�U��;q}�S(�⑅��Zҧ��&���hM ��	:�8E������E
�#�?��`�.y���XlxVHYEB     400     100�*1�p2J����r�K;79��D��0�K�����dF��B�����MO�f�K�;�>�Y���h8�HNS

 	��5ן3��u��P��S����Ě�%��jir�3����|vF���{�������y�b�~΄��vl��b��XЋ���8��[�D+mLe�&�h��$�{�"`�x�A�C��(�fg�\\:S`R7 up��W�%�X���>Ѝ���|���x�ʹ�ީ�d5XlxVHYEB     400     1f0$`�E'ӗ ���!�ڙD4H?�BR:O�XG�����CH�˦�Tb�b��]��xxh��4���BA�.���Ϸ)]4=�tx�
�\�=�l�a�5&��(�2"륞Xo*p�?������@Jq&�id��]q��S��TGfq��C��R���p���\B. b��XC��{Y��Է��MyO`{�U#�C��(V�%�����Z�\�}����?k�"
K;�}G�Ԥg��T
#�B�j�дI�g�)�<0�Q�́�$[�����[����V-۱R7� ��~Bql��l�;@�s�-��rC"�J�!VJ:N�l�#���`"��� �FO�P��k�������,����b������AC� r `7%TL�Qh�[&0Hn0��c��?�аv�����3 n�s8�?2e8��\��GJ	�4d�E�7�B0kL��~�lɀ�d��2XIH#�'�j��n���_�\��L(XlxVHYEB     400     230�P�>ӰŒ�^&�?����3)G���+ٗ�����D$E�\�������C+53���u4��[x�9���4߸ک�̂�!�����cS��K�cƶ�Kh����&����g�N/'�z��V��7�>��B��HJ�XF������HhH�f��dt ��,��S2)9顑�8�C���fp24��l?�Iq��'����6>���/�O|U�@�Kl�n�*0��<�i�RM�!�y��׉f����� ^a���ҵMv%P'�g�)�1�^)Y�@�jY��ƍR��鶖�2ڝ�k����-�F9(�Hm[Z�#�ƶ���xM'I�4!�"B�W�3iP�t_��D�v����+`';�g���dk�g�D��1�%���b6w�.��+b��	�k�+�=�V���M���3)r}�FwNȃ�Jc�0D�%n~:P�$=��q���f!թ5�k\��b���Ҳk�[��%��}�߼9�4=���NU@��O,�>d��&	<���a�{*[�%��:���/��u>N���Y~qT�&_�d�~j�k��3��.��3�XlxVHYEB     400     1a0��T��Ey1�>bQ1m. �*+���n��"U�D
�Pu�A�M/�I����[) i�%ܤeֶ�G����D8!����@�A�>`v8K
�eφ\cPEY�S�eyc�av<�@ޝ���
�%0��t�%���1�;�^��7;εXVp� .�c V��.��z5�E��6d2׻����"����!�L�l��z���$�fd�y\|�oF]Y/��<�IvHz�P�F�/�+��C,X<���;�0�j
 ^�,�!		(+/Y�󄆺ă�cuY���Ty��zm!�Qh�Ƥ�ޯ��{����gX�:HZ�B�D�$m-h�n���=o��4`������`p��@���E�u�G`���b���^▋q��Az#iN\���u���͌[\Iٗ�e�6�$�-���^�����)XlxVHYEB     400     1a0Pㆨim4�f�@D���ncۨ�ic�W��.��� 0bm����ZW9����]w��Ƶ$�0�Q������7��̃n�n�����S��8'l*�9:3YF��)<��wr��Qwgw_���eU������&r#�����@���b[�kBa��Y���(�Y��84��w��4�����v@���Gm\�w�j��y��FBž��rf=	�z�v�dN��9<єn��MK�%���}4��4��L$c2MH��a����]���yU��W%���bg
��Z��L�]�8#�z�8�X�H "��rN�ݎLozX�WB��S
��o���'���3M�A{b�eJB2���bg���Q�u�r�1%�b�g���.������ĳ;�Nc�����:�Ў�c3�b\�XlxVHYEB     400     1d0p������7��}��R�[��o�b���_@t8���KL��:���
`���R䝮Į5�D�t�W
 �B��Ȭŀ����tn�y
ά��[��U˖��l�mR>}����QJ��~8�Z�e��\���P�z����ʢ��Lw<V�2������|��?f�V�Ȩ�_����������>�opx�xi&�ca��QN�U�|&T�~0�~i�����.�"��n�"�|����f����8k:
})�umi׊Z�t��!��1~������ƕ`�)�|�M#t��d�Gi���Ӫ*+�������#��c�eV���Ǣ��@��9�N��Rŝ��O΅m������Q������⹼u��--�Ƭ��,��(���gMX�CB�\-/��a}���? ������Ee[�+/]p�?\�*˅HK-[W{Ӧ�i�Y�NUqJN*�XlxVHYEB     400     170-�EɈ��pi�&.>�����V���W�|Y�;�M�������w��K;
���d��ΏP�'�R����Gzɀ����Z'�T�<\�CD�I΢���K����f퐛V�ML!�Yn�p���|:�6�Hd��#%�Ƒ�6����>���ٗ�Pץǁ�c�"L`���y��󂪮�J^��}C�WMN���/1boE.ҏ�'��ڈnB���3�j=��V,���R�l��BE5��v�����]Z0jm`W�����/���i�����LK��5��h]�9��m^���&`ڝ��e+�|���`��>â�ʇ腿\��f��E݊��Ql��^K�L�0�55l毴V^�Ł�H���)[���A�VXlxVHYEB     400     1c0"K&�����z|Z����e�}z}7���!}����i/I$<�g
ZK����'��9���NiYܔ���YL&�'Eb[�_ɛ�PO��ⱂ�o
d��PS�C����D�I�?�n �m�K���ڏtnp��r�N[���Dx�r��ݚ?>a�Kaou��FK?�(-r��Z�G/&�I�M\`$�sG��f
��>�C�w+�Y����B^q���Pjs�r������
�O�t2	�-�	]�f�Bg�"%��W1&�ylM�x�z 2@n)d�
���6�$4z���/&L�	&�I�
*���w6K<��q���V|ӹ�f������+M���>�l�1ӈ�5�-��_��q��V���z�N>�w�z��`&��)���ё�ᄰ��z�,׌j?"��[��y@��<�U���0�^��6`��D�����:f-XlxVHYEB     400     1a0i��42y���8n��6��;�t#K3�k����ϵi��*px.V�2C)���ͳ�X��w+�K�㘝K����C<��W�*�Ud��dk'�AA�?5�P�*p�~�;���:#��B[-`�sD4z�'�ǉj-��	Z{���`����Lp�k��Q�����d���ي��~�� $��}GިM,̻�9 2���>��u�;iPg>a�m-��^���lQ�Q�A��P��4"�#�L�"�a�EX�?a�#��E٤���q�ag����[�
��z�g~J�B�YBt�cߎaD�L���)�H��?q�{�Kj����غ"���u�M�Q!Gd��T���1['�,���>�Y���4p��vU\b���^��oͶ1ܘ�h˓a�1]0� �J��XE6��a�W^1��(���0�XlxVHYEB     400     140�d�p8��o/�M7�Mz_�����T�
� �֜�Us#�����ɨR>�p'F��7Hļ��Ngq~�"�G�A���ҧ�_!D�(��0���'��ܱ	��_�6���v�J���%]i����s���T2p�X%�S��`�,������\�3�О�u_{��e���B�����)`@�-i�hv��W���ځ�������,2�ڮ�D���[����1�G�H����������gNqm9�Y�oQL/�*��G���L˟����OS�dٯ:�-r��2|�d����5Eh�����	/P0b�:rmn�74��)��L#A:k��XlxVHYEB     38a     180���Bz5�����}�T'�r��ظOEv�F_��#�G!Ŵ��J��丁�t-nIQ���}zָi��.[�,��Q|��V1Ƚ��9��/t��O8��-ɯ�%ڤ�&�<�/�r�_lE�皏�R ���jldʩ���a���!f���Ƞ 8Z��nߏ�T����5����5�4�J�����:]	��c�w��B4,B��+����3��gK,�&��CK3}Ӕqx�G�L��Js�G��}>�J��EyJ�xX��e����8AW��Q^D���P`k�	eK ޵*����*◼��'�R�!ǚ��zV��fK�kcC.k퍐8C���c��r�=5<)1�I>�����m���S`J���