��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��Ї@+����:"�� �g*�j����$zqB��`}��F;: ��N�m��v����~��ɝ�}��吻?W��y�\��4�,��� :8a&a�"d�����KA׆Q���\�W�U"�h�<�@<���-uĺ�oZ7N󝈺�����xnU��������5��g�$�Õ�����ϫ���dP�����</���G���"Ca1oM��t��t�6y��Dƫ�vO��"1aڅ������Bʀٹ���=� B.��֘\��;�3���!V�1���BB��e��c+�\=���lgƎ��*τIGSYK�ԶҠ�9T� @6��U{I�r�7��_���M�-�������$r�Sx ���"Ul(��J�+O�"��+õgJʅ )�����A;� �%S�^I� �4���}�3M! � �.Z3%�ղk�XR"�ʦ�B譼�>׶H��]z�o��Cu:�ñ���؇��ǆc��j7��S�o4u���,im#�cP<<��@Bx�U�r���>#)�n ����X��#܏̣ � x|�B��U;��!�)����Kݵ�{7A$)���kB�����l�Wq+yV��ż�	�~����iA$'��uG�
��3���_S��Þ*JR �ǟ�h֊��ax�@��x�-����1�q���4&nC�}Vu��5���|ӄ��H�I(�̓���C�0��5�90#<P�%8�6��+����[���������`j8��E����Sx(���AY�I �����a˴H�"�e���m\�R7�������2�)cE����|J�-ج8���:��v����@��\���$�e*O�P��"�S��c,R��l�H�AjL��K&5 v��M�`�W�L.����������/��M��j�P ��$g8�v-���?�<'�����/�X�SJ#��$55�V�3�Φs9��"��l�ҽq�^��"�/�*hL��m1w�ഀ-_o$�`�/%[2k��*�.d�� f���Hg�RKMj��R��4U�O����BM���:$}��t|1�[�g�R�*%N��I���TI^ܗ�d!;�7����җ�T�[�w7FU���q���X�G�a�ڼ�>g9YpG��>Ǳj���5%�I?�G��j?�MN3��3{p\>�X_�����9YܟE7=����3A��q��\,��3^7����ٽ����}@�<|[}fX��2��5'�4���ؠPW+� + E?�G����|/��$�����8g+����,f�_ǰ�ϳ��ij����Dea����V;�]6�l��a�p!�+�?�
�KTS�K�fߚ�!.�޷Jo�?*���)C4��v�@6��ѵ��Ӷa�ǣ_rI7�<Ţ1�(�/i�Vu�i�a��+��j(%ǽ&"U���հ��.R�K؟����DE�)KFgR�B�iw�*v�Vva����2���Ƙs�ī22��QQ��կWa���B�DO�})���1�sL����I꣊)����/q��ؗ�-+�)�{\~���g6d�h�>=��U�\k��^�(�8V2�_���~�U�E<	w���9�i��e�������g���v*������ޣm��g�Z�7����σ��e!�@��$7�:g\=���r�{�;� 1��kʛ�~:;�`Ȟ6�+7���g�ί(��7v�r ���H:�=����ɽUp�%��� ��P`?t�f�O)�\�|魘�^��#aܻ�Z���K4�w
���#a���@Ep܊�"X��ܲ縐�GƉ�~(�EBئ@Bx�2v�)����H�S�}U4�`~r�ʽ	�v'=G�v0�foi��̳0�#_]1 ��0o����ÂJ�l�mF�][	I��)�aR��t�����,���f���g,Q���D(�a#%�=�V,������'04y���	'��'�!���9��t�9��.^Ê+��q#( qUhؼ���,�Ġ�;�Q��ԫv�v��A�pY����XZt�ǒ ��ղ��T�~�at�;X�p���~ښ�I3�Ǐ˩zo��Ǳ��	RZݷ����3�V��Ήq�H��14���Mam%jɷ���C2�};�	�e�6�d���Ų�d�WM�B�,��4�w�VQj=6~M�=��׀|v��g�?�5%�=/]!�4э���{T�°WA��
Y�,ZyU��$_�2�dv���}@A<����o��IdXI��T��x�#���^��5e$@����_nFI�e���Ţ"���_��}��w���B�uX`�$��l	��Bm��|�|�gXrW9$��X��sI�=�!n��
`<���H=�ܬP��+(qg���Z�]�l�w��0�티����t�>@W�W�J@�t rtqPJP�m�\_�b��M]O:?C��7=Jϭ���x������Q�22S)W�*^7�҈E�1��-���1	4U����c���O�*�- =��OZ��ha-V��-Gp>��%/� Ň��8K�wIt�3]Qc`*C�+?�l��>E�f93B�\r����&�hv�lXY��ٌ�~�8ɩ7�~@t<7����c��{�و�4G����.n��,$
n�d����3��g�t�W{x���B����(��')�0�nn%Xa�v���{�����=o��ixM�Wܔ&gP��o��]i��H���+?�����,�/
ό����$M��s�l��'n& )��A؜<����Ϟ��Qf�Kaއw�����])��MAr��R��{4��a�hn+&��nE1����ű�z��a���k�����v	`�7�!E��t��OT��е����w��q+�I9���i��W��Zb��i�g�r-�������}���@
N�����Θi?x��(��6��OyBV��P�3o�������?
�]�e{&^D���4�
�1��r��^�m�aW�-N��� �w�k�K/Ȩ]���9-�5"��fWs�-���7�Xl3���G*�H���Y�c
��z_f��Y���(X�D1�����'6�|�v�_���;x����d��6z�=�(n�M�1)0�J�z3��@!��O��^o����d��,5�����Mu���a!����kp���6��ֹ���b�lӗ���X4t�I4{�[���'���Y�X��z�Gr�/Z+�b�E?}k�a񒗖���Zh�!���yN� ͐��SU����7v�`�����J%"��/����� �N,�8��H �o{F�ŝ���^�/�(*��3���i��9�rˆ��Iy�LY/A����9��aV��yN(j�CK���v�Bf�����B*QRz�����m+�h ��=�_i��i���"�Y�+S�a��Qp4Z��c��VN�1i�4�?!���y�.@����-.
~b �����;J�����n5�cX��:O�[A��a �)���KӖ�W$^Y4a8uA�6Y�L�F\# ���*�<=��z�=�5v���m�~����(Hq�rK��6����AZ�Hk����ؤh��ެqO� ���P.���z>F۪�ޓ�L4�ě*��x�)-l��9��V�K����Q>����q�z#p�j[�zM8M̈o�r)% �-1�ʁ@O�`S풖C����x@#[yť!�npڶ�"L���%A�n`uþxGf�B�h8�4�Nfw�X�� ������%�����G*�*(@11�U�xQp�w)61*W�<�u���ؗ�5���9/����[����
�БVfV�V����/���q��|���\��"*K�<t�? ?�	Ɠ~�Ƞ!���X(|�� i2��u;�6�C�/+"*�(kx<EZҎ!`b���]�A�us7p�n�3QK�M��{?�73�v�q��ҷ!���#�}���F�J�_�"��3�3k���33�����?'�]h)�u��U��m�iK8p�[��MC���,��a0 ]p<7"o1N�G��ܲj��ު����o�}`�A�9���(��$���OL��U7�&<��iP�wf��X�9��
ޒ�0@�x_�����1mz�d&][@�a0]���S��Ԇ�:11(��`q܅ZnQ��/!Ƿ��B��߹�7{�ч�x&�����f��8�h��ޓ�#B��/�,���5E�<p�cP���wXF�w�y��cR������խ]P"��-Kk�N�Q��v���\���A����-���c�Cz��.��KXx�U��E�f�H>�(�i��|A��A���x�����3f��Y�@�Nh�XW�L�'>�h8�O�ު�}P�M��N��o�� e���qv*��'X��L+3��mĞa��|�5h>)I{��2�+���p�VE7�t��}�ls�g��騙:p�˨N��#J��l���K��[ёk�P������n^��>���r3 �P�7�%����UQ�-Yh83j>�k�-w�.�\s���>	Х�u��~_e?P�D_z�䍖��G�DT-&Dqo|q(�J�T��/I0�Yq���d2Y����5k
��sG�_K��Ӡ���ښ�Fm��Z����A��5�N;u4����͔�3W��:�2���Ң7�`B���h���h݁�!Q�V�����Ͳw�Xf �
�L��$h��.=�x��N^%P�[/��3�g�S�C]�)�y��Z�ȋ����Ժ.剁j�ޖ}�pm�q����9�x�3�U-{�L>*�&��D.����Ľ����ģd��S��~q��w�V�()f�3�:��9��W��5hz�	$�����U9ϢP���=��2�|�D$30�sf�J���'���6�ƣc�s��5�}�[<���󎿫�@	�
������b�M�c��p?�W}�b�^�d�m(樉A,���� n,�x*������)������@�������%j�zKA
7��tY�� l�f�H�6�~�������V^:7ks�ah#��m'ϓ*(�:_������n�=�}� �b	�"Au�o|�oHP���o�J �,�q�����u�P�qQ�*�*!���u��_!�vJ������C��EX'�C���j���+�R���æN���@`�p�n�DJ����!���~������EU7��tߘ>�yd����P	()_��{g]`���}�6`���Qlr��t���p�����f�c�2:o6� ��ic�,�t#

~����q`�_������)�|��K��Ľ�����i�)o��uVX���[�����s���&X�$�u�?M�
n'Ａ���YOu�iBZ܍&��*���d��DO�Tѵ��ۯ"�No"eѳ��B&+9�-���UA�Uh���Z�J�P� ��� t<�1�b!�(_����&\��I�	d>5m�Ku1�Rbio�H!H�."4�o\�H�h�}��n�����3�H����f�,���C�����<VD%N�1��-B���	M�����Op�h�)�*�%c����vjZ:߷�����6-QU}s�C�����v�\^?Y@h�$���"�C�c�j0��HL�ԉ�tvl���/<���NI��2���]7/���s��Ŀ]lP^��)P�������vS�����L���`�:<�T����/`t�g���Uҽ��H�ԯ�Í� ���\١C@���ΉÂ��D(��W~�K�>0��1��J�/� -Kѻ�R�@�樊��b�j.��i����N�3����`7eK0,5V��l�r��d^'p��K��Fp+򄝓ٌ�	v!B�خF�����G�r�ՖM��h�Ԫ��(z���3F��]l��af �0U�"K�&5�������m��A{i�7i����������FN�}O���Q�ű���`��}�/�:1��\���������8�C�>�ᔍ?@/.���xC�J��|�9z�w��e��6D^�b�핼<�u�O=�T��i�:�%��]�S٦�\�� �ӄ菸*	:#��8�c��J�qa��^�7@l��lM#a]zZ9�5
��5���˹�ς�����ѯ#u� ��a��A^�4zG{���AY�%A�̓���'�V�t�t�|�������Ois v.Aч�,4�.a�RrV�dq(�Fd\�����mʚ����-2Bf��)V%[���7|W��#G���+숨p�B>R���?����Y��'O�ձ�%y@�O�r@�dm��/l��*NA!N`D�'`��N_m����Yd_�&Q�ٵ��8W���Z�ݎdAb�Y��dӽW�f-��=c�R�[+�{bkv2_��a�qݿ��OM� $�iQ�I��R����}I�2���������e�D����{��R�2��:��r0]�04='�p�=?�Ѯ_jWGWٌ`����W��2��]vw�aWzo��#�J����"���0��L
�]r�[�	[�- �L�Q�b�+q�Z����tNP�UQ#e�����"���ΨE����q. ��ATslJ�$b&��Pr��&]���L��;\��9=>�pb�8	��)���

7��ã�\��V�T>��s��0]�!c��' Y��x���9~��͠G	a�6��Mal-Ũ"�R�q�'c�s�%��a �t%[�b��cdT+`��`��%�`�\	�<���s�
��i]�۪����1B���f�jx���5D�Axڛ��Gr�ƚ�@�%/X߶�o���r�"����W�z~�ue&�Rs���_�F���+h��$�h���N��e&����T��Ѯ>Δa2(aa=w��fI��e�m��蛺���u�!;S_.�g.�,?�f�e�Y۞�dR{���H�B�\����pcM����UT��l<�IE���|N&�/#_��
-[����6���3+�7WUC�r��):�lGT��Q���z��)!,��w �����Kd<���K<��oʈ��:\y/�ls�y����.-�^������,�2n�8�?��s�Z���eC�9;���)\���� *���<��N���c��&�g��Ǵk�a��Ax��^1��}]����$�j��#���`��K���v
۶ڌ�A�� �[�ύ����B����
�tp����j1�u?ӡ��0(���o�V����޳+%���	W�M��\�<}f���W5�ΕiZAT-Z��a�X�G��L4�<))#� �(���iVA.��{��	tz�������Z�P���| IuF�Q��E��Nu�>N\򰔚�4������]�ǰ8X�#���x:��z&HnTM�k�;�ɔZdC<���%�E,1��X����[E�4���}?q�Oزi�sgTN�&eo��i�0��1q�����5C�nõ #q���V)����{�����#j���|��tuϴ��m����zu�V�����$ �ag�� N���Կ\QӓRvC�R�2p� ��AC;���ۅ̫�s'��심������d�,t�����qXp��$�o�u��e��G_�ੰ}՞�v�����>��^!􄉭y��o��R�P���B���B���z'"b�o��8�L�~ ����(}�;.��:`��m�A�pϰ)f�Ɉz�;�Gކ�D.�x@!�"�EB�ґM����%��ߣ~�r��rw�)�6��2�������/!��_�
�"���oi�{�#=j]�xuw����d��	N�Mp��ŔBi�ؘ���¼O����wH�R�h�9���:����kI9x_���4w��,>��D����ES&0>������#�[��9R�Ӿ�Ju�o�|��PF�ά�nʯ降]��f�f�
.�R��
��^LKYT�����dEO �5Z��?Y����b:2w�����P�f�����"��B��;�FΈu�n �CE(�Tb=D�J�U	dP��	*>ؽɹs�xFMFǬ+�RC��]E�&�j&dH{�e��y��B2�o����S��Ӣ����8���
;�h%��+��ね&񙠟??�#]�D}���;�����iM�Ůla�h��"���z�w�xՕ`0�������.� J�|�����~~:<=����Y�!X%� ٮ
u�ͻ-Wް���9�y���R�(IpCػF �k䲫�#�P�#o��3�<4ao�5/�om��\,�v�4?m���]ԯ�^�C�t�Յys�e�W�5:�.��F"�˶��]t�n�!*f+�� p+������١$"J*G|�:LO)�@�TR�H�w��!M��
�6��V��rҋ^F7�	�Mcܔ�J	k!f�����Z��}�=pာF O�jt�N:��Y�>�1j��0Yf��,�h�b�(\�1ʲ>��ΚB���1�ԁ�����F��{a�L��R��ޱ�dNn�뺩�g��$��ߦ���Ӟ�sc�,'e�d�^G�Ӷ>���S�z�FG��
LyR�,���R�G�~�k��07�Q��S��l�����(<��o݉Z̘�nN%[��Ű���;?�6
~�볕Z_0,gK�Di�MD�A�on�|����T�9�JDU�@�f�����~�\��[^F���ウ�������>�V��ҴM�Tȯ  ܜ��ďȠ*b��3��N�F@z��Ϧy�T�_4+�yls��5��o�x����P)
"�0}�-<�� ��E��_
SpCuR�A���j�jBT+�^� ���	�b |D�\K'W�FT�^	�3�h�^��ݬ:.Ŋ�j	R���|�b-����'o��`m|��C TѶ+�g1+�,#ωjkxqLЌ��ji�ۡ������^�>�`��Bns<�!ʐ�|ʇ2jn=�2TO�57j�n���f0��%t���[�����(����'�9�D^%��M;y��FZ��U�	�󍎽PE6�]U;�&R��u�\i�EJGKVe ����^>�.������58I��<F��U��ڈoM�����g��ͅXǍ)�&*u�&��ׄ��K�1{� �7�c��nոX����.�������xEl�-6S84���wx�!"Mem%%�U�nbc�Ӑ������`�1���?\��H�%k�`@�d�D_�N��v��g=�!)�Ůd
�'��������j��>�a�r���ȯW��(i&r��y�!;z[�̫��ҳ�"���-i��&��2�Ŵ�)u��DM�QJ��b�Lv����)7��X SL�����&߈?I.�A��q\1%�M��q6�H^	��ધ�;���+�"�K��[�<��@M��7�+,��)y�A�B*(���o߿(�G<-��~Ջ�P���_�h"ǜ���W
�J�k`����#}����y�3�D�ϵw�=r)l�"�>C�+ ����N�N�5\R` E�����_��Hi�]l���+��g��ꜘ�T���y]���I���F�S�"��:gyȇiXEؚ��
��9��Լ��Z�s,:���</#�}�R�R
�3��N��A��q�� ��)����%2���G�yG�f���� �X���]g���UYDxB�ڭ޴#ĊAԫػ�|Y�&q�)�'#����:��H�:�t7<��:v��G�)�������=ĺ��#�T��Y D*?��Ŭ��:ǩ��dD��ʄ��g;�D{E����H��XAJ������J�v �a��I*+�?os��T;P��P�N����v���!"�ҝ@sT����5U;%�;���/E�%��
'Qgw������ӷ�����/���#}1W��_'���j4<��[���0���h�@��2��|�^���#X�t�ᒠ���D������f�xL�@P,���(̸>\e�m���q��NnFcF	��&��fK�)��}��p7��P�bMZ�:��l&rd0��~_ͮ�!�M�v_���|�З�o�|��v���)���2��w�V`�l�Z�4���0$�P���4�c���TAѧ�	�u2��=�z5��+��i�i 9�|�#^������
�uS[�Z[Ud�둮���[p���:/e��闫��m�k'���xA䙢漟����@����N�;�Na�E!^f�&_��&��q]Ǎ���(�i�O~�MT��A�:c!M�9���c���W���j��j	jVc�����P�)�U=3��޺F�W��P��"�K���!k���[���;Dr�P�Ǹe>6�����A\"�_�r�b��x���&��dO�W��#~�� *xw�C:3��@���P�,Ȍ�_^��!�R�M�%CP���h�<��'q7y+�D� �@(##�ZS��?�4��a���J���ʬ�'�NkA�[,/%�g����FӴ��Z5���yd�����܌���v���#�Ҽ��o�d����/���׻���c��,�%X{��e3�!����e���@�/�F���;�T#n�r�l�_���5�׌x0�Ad�%4>zU
4NV�����(f�����ji����^�2ڛ����D�{e�{�o*�)o�bᩆ !��o"�[�f�BQ|Z.[��a�/v�$��J�u3�|�=�wDxes&�ZV6�Ƨ����<7O�ь%M
���\DyQ:���\XyjRe+I	�3"�e�@L��b,���U;����zW_' ����o�W`��n�� ^մh��F̆�O����QQ��o�`1��`?*�"F�C�/��T�/p�p�6��J1�V���I�Q�e��-���/ӷԙ�v�zNU ug
-�8����e~�1�%�����]��W�z��-�����P���C������CL�ݞ�om/��&�P��>��:SB���I��H"[E���wP�K�'���T"�X����:���h��:�MP���#���}�mL���_,�uӿ��#���:a��Q��7\���fF7I:�(B�*Ğ�/7;�=�|��& �TL����?����f.���;����4  �ͼb(x����Q\���`wKx������$u,؃�����d����B�?�rK1X+���1�e�q":�m��G��d�A�
�xӈt�d��N��4��E&Y�tm�E>gc����w��`mǤ>�V��l���ɓɷ[��!�֋�z���w���u_��6�M+,�D��?����w����ŉ�pG��ٹ��)��zi�]�ی��y�ŗN�s��
�Q�$��=hu�5�ۗH�~���z��e%�Tޟ��Q(���#Z��sD��7x��2E��0 �����[��֡���[�Ծ��d)�!2>}z(Ed�؄�������א��H���#	��3��[Vp��wl��x��o��߈�`5�|d�`�Q_���ͧ�vA��m�1�U�t��>���#��lr�ά�G���\��-!Z��Y`3��X��U�$}(>��Vshg<*���rt)��Ɍ��}v�U�-т��qB(��.���to�[��*8�Js0q��-	��%OȚ�܌������(�Ikݭ�� �K���S/S�_��Q��i���x}x��S����z>
�c�zo�BC�|*c�̇w���9�U�b�E��y�1�?��{��;Х6��K]N *t=��a��7����)b5+.��C�GFO��/ʇ�1�~.�Y����ى�C*ig{�{#+7s��ο�x��|�ɶ�U���f�[R/�{$*b��+{ֻE�����TX'�OI/�)]3�{���<$�[w{$��1,U{l^@��U��,���3dc9��ػ\�o�8$�����Z_>��?�7$�[*j	��t�xfM,)�fS;�*t��<s�(���h4c���+�D���� ��4�\��P��id"J^�.�`�Fb-��hL��t���H ����A"+ �E� ����O�Zau�]��tG Pʹ8�)��ώ>��6��~���X��nj��L9��6@��G���Ž����:,��&f#�c�s��7�b��2?�BH0����;;
�@\���!�٤�_d��(,��۴���l�3�Z�#V������R��])i�Є[(_Rj�@K�>���R1�H��L�.���\B�~�\��ѣ�pz�$]ÑTؒ�A>+��t��fO�pZ�����`�QV�v��TN��?�-�p+�˾��ҋ�<a��@oE�����&��W�y�x�D���6��t'2�p#���d�z׭�F�жl��)&�a��RS&8��ѽ��C=m���L�pb�یc���(�T=�
�%��_���C6�.>lU�Sk|����y�1��x�/��-�]�_y���i��p%G�N��^O��15��x�8:�yQ��X��T-�����ݯ'2�	���<�'��1�8���ZS���ӗ8q����	pD,(C����A��@�.��J���a��[&"���? +����i�Γ��n5�eہX��0�x�
�D�<� (��&u�UpΒ�!��=gZELDx�Y�`ڤҰ�c���W�HXxh:�ޭ~�[|���&�XBG1׏։��0,U.`A��'l�ud�v�*a�K�)|�g��FH��?Uo�?K��qG~?��:�8�v�u�d�漶�=:R�y`Uosx-�_��0��~�D�+�]p�@� ̘Ek�yIS.����S�'�o��Ǳ��i
��|�k6v������"G�爽0R��W3c7��"���8)��YM���4י����]�Ңx�޳�_D�r�[MB残,�,��C
��fY�mt�E[�63]�� x!�3����gf�)g�C��<b}��ɫ��e���������v6�Z�;8��^�X������@	h-ER�"�	y����\;3�}*/��	�v��4Hb�Ty!:��ut�4I
9fI1�
i�N?(��-�������]v$�\9�i�?�q_r�����[[�K��L
i�h�k�a�r����-�Ӟ)�ϰ2tsU0�ҳuG�&�;��]�c;�c��rSsf3Բ�T��+���D �0E �E6���n�X�t�<�|e�� �6����S��7��+1��s��?��0���8�)��Qȣ�!Y���\4��в�u�T�jfw�K1A���yw�z|�j���֨Q��F��{�f�)�*H�|��
nt�j'�!{UN��Dʢ�TM!o��%�w�(I&�IB$b�j����^P��4�w��K�懄�L��쁚Zov��J��'�dj�J�7Q m������;{H��[z֑�E���w&�{���&i%�kC�	�q/	�J�����_�$�G�l`o� �?%�PP��5�1��$8�7X��ˁz̖��|FU��	����:;&6�
l����P�����[�(��b� ڐq�LɢzOC|9��%I�۷�+;y�νS���5������'@�3 �)g��oqx��s+�n��,��3�6��KԸ�B{zʙ�d'.�}Ȋ:A�����������M��-��ϭ|n��  �}���V	ڗ�Ěv*���aM�{���!�E�� �(v��QEKx®��E��^�e�A�pύ�U�X�zZM�����xUj���L}��W�ڣ�f��b�<��W�q��:�z焠��uu�]	���ޏLm	W?��E�'�U(8�	XW�6u���08#�F�x��-IIm���#�t:��Zs\�7�g(�Ïʄ��ْ�xp@��c
�`�;lz�/`��jX�����N��̩�(`��=I�����L������񬌴!<X�{Dc&vb�M�CӮr�;��P"��p�3��t�~��Rʍ��i>	����}���/���O܁�]V(o֐2/���dQh��R�k"H�D������1�� �q^�ʛPy���=7k��V����f*���*�l,u����`�|�N�q���}Ǭ	4�Q4�H+4`�biz>O}�
�:�3m��4���N��g�o���F}w�$R��%�\�Ö{���y4�&3ll��TX�ҝ v�<���ɵ	6���(�BG����a��� {�쉰�\*� ��4�,�w)ł�j~���tnn ߹=�Gi�U�wU��I�M�!S��e��D=�Л�hvW�m�a�;��u�$1o�Q�|7{���<�3��7�m�y�*�y&���e�Q:�_�7��}�&���/b��6w�n���M�
����'��d��4�h�����$�Yǭf�j���(ƚڣր�~آ�Rx�9�(uR,7�9	@�暈K��p�42ZT�B8ώ��VЮ�Z
xI)5nçh����9ym�oK���X.wyRw�!p��0�[��Y�^�M=רR`E�����%�Y�*C��g(�%֬&t"zѭQ���]H����љ ��Y�Ɇ���k�.��y��oo6R���궢�mZ���|&�x���D��O?��r%��9��*�����]Yfڑ��(� 9\�p�p�c���]��	���&�AQUx�N�e�8�䐜������@7\3�$�d���L�9W���Q�q��tm����꡷A��h����=�ǯ�0�P�-ˤ��~Z�e��.�(��R~�?�3� �e��!����~�P�>��8�g}�Q�ɔC�k���A��)+ ևG:��7܆[.�%�d�W��<�Љ�pI����;r�W
��Ay�z��v�0nk�Pv�?B`�#�\gT"[юL�QN_׻�e��2�1%��;�`�Cy�#�&&�/���K�F�m�J��;�O�Z�����҃`�����X�|�d���ŀ��g޺�T���;Q*�WY��U�t r�Y�&�N�$l���T'�ˊ^����g�?�)I8+�(h�Iƫ���8��k��u���U5���`�����{�O���Mޮ�J/�G+����ɽF���"��s��ԛ=��7V��'��K>b��q�kCM�,�/���h:�jm5��K-?+�/}O���>�XU=��G�30�K���jE��y~�
ڞtD���琉�o����_@[��H4|����#tQ�pT>5�� Q��)��l���iEX�_d���J��O$�yO�v_�(����O�� ���[�'R*H��S�Ƈ\5��:���� �����޺��T�u��S�� �tw�d�a�ո�$��P
�b������h�>���;��n��vlkSP��������~�Њ�0D��ߌ9Y"n�6�j��_�^���dH�g	3��"2UR�c(� ���om>H�	���mqpH7����qL��̓˱C��rQ�{��6!��;��ܐHlN���QԼ�X��䩴���*�Ȓ�ق��(NIыϢX�l��'`�O�V�l�����|�c�#?�/&���iݿ�3Ö`���f�:E)SCSG���"�4!��Nmbٸo��ޥx��8ĸg0<h��8���J��X{x[/��H�n�����-�����V��	���J������	��y>Lʫ�����Pm�)�&���c��p�ƭ� ���DQ�'��S?��+�C#\K�>�z"�%Zʗ��`)��)���,����4�x���'�s��d4���H�Oap�K���5v�s�*7
zV�j�4^�D�+*����uf����#:�-�U���	q6�}+7>_}Z2&�6�mD8C��@��~��o��y�&[4��2?,�-.Y����Jl����8g�g=�?ɶ�q�`�C�!�:��	�%L�ߣ�C�Jp%�\�d���װ F������1��#�̮�Y;��#oZ�(�]|�Uh�'��(f�o|}�Q=��1�����B%![�����x-��gx��l��e���k��;�^FF��!��L�h��/*��UZqĦ �[O�)���i�9����yԨL���z<�����s�@�~��#H� dq&vd[X����J��J~�iIW�:��N��߼�Tb��ў}@�֚o,A�7�7�c��+����KP������v���ְ�;���^�u�o���V���x�B�]��l�r�|v���*IG��B�I�%�Љ����#Z8U�?g/�pǋi�H/�iXJ��"���T�����@��x�����>��6I?L8e�K|��<ZՆ�s���d����իz�*47>��24ŕE��`3�����(�b��աI�
wʝ��|!z��\��Շ�>� �a#�ɦ#跎�4�Qt�G&����4�&��� ���;�sc�|S�t�1������I�_�%a�8�*f�"���7%#��x̀zYf��1��.��	V\�Z���!��&�R�B��*WkKC�ώ�'�}��[��j�:y�@�X�N�0���-�8��n��!F��j�����=7�&�E'K�>��t���:�Dy������TJ�E��qC����`�@�.;�1��}��={�(��n��{ ��|LT�'�
��Ɗ�<"MAQ�ۥjs:LF�X������!�d�EI�m�~�]v��Lt�5I��K���U�z=J)������<)��Y\lÜ��%�Q�҆�������'��]g,\8r1~�*$̫n�[�)�%��*2R�@�z�
ن�f@
��iww�P :�S�gB��p�`�kku{�ޞ5�7��ȲW�efC)�o1�fӛ�c��hfkE$