XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��&!���؆��������p��Q�	JU���C��BpX�����_�u]���ߓS�O��Պ��h��{� �H\Un�������Ǟ�]_O�[<Y���pdn��V�C�������i�H�or8�2�6.��!�O�D�U�Syt+��nǻ��	`�v��>臒q�h�xgm�R_t�Cc}(�6�?���z �� ��d���aEm_���/Sb�Ri��Z���14���hkp�\-u�[8`����@0���H�����5$=�B���h���,X�EVoP��KL�@����RCT�[���[���O0�o�kAR� ���mQ��iv��V�Y6�����bU1 }�hvsW�M����p�T��>��ֱ8��uU���}vɋJ�@u"-�xpM_��Ak��t�-�E�P�FIX��أ6����b;P[���ƅ���ʺ1�Ѥ+Dht�פ����Y�Z�ߕK��qձ�T�`C���\�/��;G�っ�β�n[!�H�J��~B�=����|!�Sf�MT���
e ͩ�Շ،�ed��j�l�!��(��߇[�3'ȏ�����?;-V��4����t���y|"rRP����Oe
��wK���.�z*l�{o��'�CS��+w{��v�#�F'�=M}G�{�S�>E�jB�"�B�8��A:��m��X���s�F��҈
3����P���G�^)$;�w]���I��4{�#Q��&N���c2�A r���S���z�Ӝ��?%��OXlxVHYEB     400     190������(�Gq����:
N�f��q	�=sf?��	v�A�J�Ŧ�<e!��bB՝�/R�rFL���բ:�L�����rB�U9 �\1gj�)'��z��ǽ��h��j)��;���I!o�B���)ݸz��xΈH�_(��0���ׂ��t�]G�Y���&j��)m��=�(�] T�@۔�gA46��V$����--���f�'�q��u�/M��aP-O�5o��8d�(G�	ð�%	�����q��W�T^�V>	ݬ؀�U�'s9�#;��R������oդ��\�v��#�F��@f�،��8������>�@�<k��! at�q�dmʺ�'��T^$GC������Tf�ĭ߾�H�@B��ǔr��5&�s4�k_5K����a��f,u�~�XlxVHYEB     400     180v�0~IAW�0�}w3��%Rpf�QO�!W ��
,���Db�C��T��
��$�H���1��yu�����i$�*�Kg��U��tQՂέf8���=���_���F��tb����f��* =�Uy0�v�7� �ׯF,m鑱�T�8�)����ÿE�ٮ�֫����f�v߷�i)�<R�K��N�-�8�^D��bt��:ڧѺ8�A��ݸ�_g,�N���@o6��'���ӯ��\]@P�\z�ظR_�!,��(�pڌef��a�-���P\��"���e���M�.��bܰJ�@2���uA�)���X�dO����|���wPR/�)�2f�
�@<��b�}/�������t�m�'C�u�;F~"XlxVHYEB     400      b0K��i`n�v8^�M���D��A����"@%�A8���}KAsۙAH�ڽ�+����T��(��F�������X�~������7�s�:����y��!'Eb�r��k�Xv̟T\���8r��
~>[��$�X�Mb�	>>�j}�G\���^_[S��0�MU�17�q{d�Q�Ky�����y�XlxVHYEB     400     170�G?��6���.�Z:��D�lP��k(�+��_�;�jf;�\�ra����mܢq6�f)0 ���U�/�M�*�6>����;յ?�k�
���-O�W5�=0���eP~�b-E����R��'W��Pn�y�g��rP$4������.���Ϙ�٨�İ'~�����7���G�qV����8lnɳ�#�2p�m��h�O���["���)�Cu����em�*Pe���r��,�7C4ӊ!�c����f���B�V��I�(s{n}|i�C&��Ρ�l��t���X��OwuCj�Y�-��B\���_S�ğD7?����:���4n�W�rX0az��.�y����E��Ö�GIXlxVHYEB     400      90F�{�����0%K���A3�R(
F�!8c�?��ޕA]�q�wA6�?l���L�hc!����g�aI��M�-�t	������b���f'��z�<��3�}��胐 ���`Lx`�o¸�ۍ$)��_s��D���S��d��:����XlxVHYEB     400      90�����-%>��T���\�3�lME�.7?�EB����J���"�W�����������5�u|��5t��+۱b�PV�*~huԦ���඙�ͅ���o�$�ـ����ޫo���		�u����t��K"ת����W�XlxVHYEB     400      90
.x�P���m7i�PdH$����g�Y�=3�U�;:�=C�Oof��[�z�84p��Ej\f�K��Lp�(�¾Yr����ȱ��!�j���y^v�$�F�+e�n���.�E��0:o�������O 7P��$ҥ����XlxVHYEB     11d      50i;�+RtmfaP$7d�Lm��3��W��7�ـ9���I�]R1A	���B24en��y^�s��A�Mv?*םe ��