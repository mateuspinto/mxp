`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
qzofvjN+wCxS5IVf5WvuvoBjjYfagLUAwn0jb64/dw1F830oCjKb61Wfum66wI9an+SifDgr/JOc
2sRxk8te9h/EB4QT2H+hrWRUx2feeY50PCY+Ya9TvMfnsOQX80gtlO1LfV9465esrba8yA6H79Ws
JxzFBlwTcZF1idmWiXmP0qE1Dw+E4AOP6MWkp9ppUGpXI/0M8zkHFs3/loaOCx+rSk6kJ6ISY0O2
MMmILZ0sPabQuAWWbth8OF0FJMWQgq7b/mpUltYrdH2ZFEaSBx8bvM8i6NTLp/zqr+VyzKxqcjEx
dDQKqu0L4ZnTknNDG/NG3w/qzBR0me08lBw33g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="2QQ6iFWJI+Go5EZX3RuhrsMaPu7v7T2luzk5XFEeMnA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 54480)
`protect data_block
Bes4xR4cDdEcsiV0tjMsw31OK25Sn/74Ew8ZlWWtxZLjnMIvKPcWwtdqh0cZLJ8E0POGi8oHw8eR
kWuo/QvZ5080elXa5RSIHjaAMFslwID+s0Oc90U2bdy+okb+1fxMy8B1QlO6ZQFsLsfyQNWztuIN
QKJ+CAD0Yg0sVWybu/TjW5yAzmHtczss/sommV62IA0r/0Q0+v5iAxx0Xvy1PZwuc7V+y/xRcURF
/i7HUqf8VP0oYj1k/2fFpqNOgQbErkyThHkMA31apn7ZVglzdPkf2rx9GOLWveSHfk8k8US4T8bi
QDmiKbsYKmnNSqsKb+Q3jb1T9pEqgCC+F5Bjx4+VqzOAgp8zXLqLV2iq7h4+XeBmdP67vRhogypR
UeJUM3dSCCvSSGOFoykMIMkQ5Zb2Ysyz2o8w3I55DCswFlNbMKmXuTwE/fDz4dkhUriMk6YLJrYK
pbs05OfxBxOatEp8Jpyu6nnVfEn3kqXB4kcz030LBFcdjtQp2BROniPTvMRI5PHZXPMAXYuyQwgY
QDmXVpMvSmHoJK1vHgMDq4kQ6yG7cjz//FD5UNBqkos3V4wOnxvXJ+d1/RTaIdFJj3OHsZthY6Ni
et/A+RAsUHHaRWmgbu6010NWNGOhHxVBtU2uLC/rEjoRCxoRxa569a/OEYPZZ7kwwuQhUfJZg6FZ
J1XUqiUJCD5AqpBXvTOEz13FsEuoN26LO3K9dVcrnv5tIhUCrp6kbDcadU7vx2xvfgnhbPSyicew
mTfNaqp1D7fZRnE6ZQuqmnZ12KJXYRnygBCET2gDijoPI+k1Xe7yTEqH91mC3vBGP9Bc2N7MKGIN
myUl13IXut/w39fQkmtuw4PJmBC8ry1EX9Mhcn7rhFzqsDdSDQY/5+fA3u1l3/UT6SfJoVEmaROM
TRCoIbTI4Tw05acNyb9m7Iv7wn4CpugNcjZ8Nxa1ezvJRrRjREgBXxN9FFhVrs+gKi5k58w8BURf
nhe8o4WIRunwy6JFzE2kATJpPt64TInPRBiEgTyudh2/cOf0u4sCNIQhJhKBo1gR+GgWksAxCqC5
5yoafZKKVnHOor79u3MykEa6gW7C8tYUdKr/GedmAtMs6WKxbN+O/fyDDLDErctE+9ySy+lPse58
XsOcoksNeHU1nW29khzo9JWYw1EwKrs9+GCt6lYTvbmhf9TKHiyOD6tpDd9JJJVUplCAosZ+vNOJ
GPvvsM3UXPMipBo/h73z0+HMkhmaVPcDrU/nOYR5zAIR5uZaMHf7UtQbTbWDMvLz/HHSrGX2wE27
mvfWxwXGSePtQwH3M7Dp7thzmL6wk9S0I4h3+CTssaDZPgHXrnkdODtJBwdtcvENARvlKLUdlTB+
LU+AanFBSAMMBPOLGeOrMKWh25yRuOYCV/fAUX1w0WwMI0PJF6HLymR0hjG3L+ziUeoJdyDS5tLL
dvsgPbUGNNmdJy1upaJw3vF8DPkpQ+kmsortQ6x1e2WXhPZgIgUzPRvpQfyZLWO+9ZiiBFC6QE1j
D6zJWWlqws/3cBt4lR8KUoVW/v4St5Jb0VSJ2fcrwh2N993cj1ZshEudFMhb/nLBncFQfKMKZPE5
m7FJBdyAiP4RJedtdQDBBoTvnVzYL0+223jP88awLieVKVnKADTsowpwDgJGsdHUFqHs5mMT4gZ+
3ucGRFCP/Obcg3IzzHQzGbrE939Wj7EgsPPOSQ8RAmqu9xguOryefYtek28FSX1beUL0u9nW0OLY
JQHuY6xlZJzgxeq6xxsTGiqXSfKt6XONOweJhMrzvo2hhoqU53YYrEi/M2P4y4r1l0jmunMW/AEi
ZEJnUcCHhZrObsP9FWmgwiCe88nZejtRzBx+ONS/9kv+HQIbxTwXfHuzxjq6c/+kyZ5+UFEigrbF
f6u2FDSg1qId2rz/UboaQ9pEDsfgQsKADPO42JjLHoQxv9wWG20UR260fWt+FL59o25C1U6tVYDv
tXGf+m0ry5Y7uYAtJlul0xxewCImycOpPEKEoR5RLE+6X47HF6R5trzsPFTJHuEtE4TmxyYah/D6
ZEo03se55k4bylswnBzE33JkBzDPBYdhwrRyrmFsCL8g/lKAx8RCRTrg4mJRuumDYYSHLjxDMRSi
UBfEEsoseIBwd5mGxpu8dhw16LnVgKy0+uiiVvYJXMwVPp5FN1A8ZgoBDR2sNmbru/zuDcRgOZTg
+XAADujZ4zhT6BCdkeekC8x9+y6B3aweeuW4ePyRWBetvv3Z/E95t3C6qpLQEFj92L8G0oMn6p9i
jFR4u9hoSoU8iH1/xEgNflz9Yxr/lkF3MddT32CyHKzFaLhrHNZ6zbzjymkIUbGhAkSP66VP8tuJ
IVv0wepFFFQqKTG7Ks29vwA/HCNTkYk/L3Nuzhe1ElNLcqPIIK5svRp/J5Vyek5Sm8lb64dGPJNR
LXPI2slxqMMtW7qAH1DwLXtAYhufjJRqaklpZuAzaKbMOqKUHiAM/g5aOXVH2mvxJXJSOU10Tbp1
/jKVI89b+zYpAkyROuCr3OEvb0xQruJqaRuH8Uj0wvinZXGwgDoUoS4j342w3EouR8/5Cb+LZvP6
ReX2lF+7u4qQQpdopp2eH2dsm1yzsT3cPM4S/tJfUCLpdKdOoUDd7EYDHRLgMrHcqP8vru1NvFTs
0Hvpi+C7KhC7ShdAMekKOTqdN+qJebtTZA5Byp1ifMOIq17hrk/CcbI67p1jLpLAv16BBlUZm5ts
TGkWKja4gqnVqZFefeBRRMMmOd12KCK0jR7ImAnjlRza1C3crDApvrlpzozDGQBmijcocXufZrH2
D6zFtvlpww/OPladDd32p80czYhVoJ7THuICCGl9R7N46sGhDlV76Liox0vjwzxAHOGNrSKZFK9o
kWRK6nO07kr5jCOwjGGZ6Pb9vR8PHzfntsc20VLSAaoMhK4RJtbs87VRgC5hFXH3Lflc7rHmeb+2
vIAYIh91+NJh2ZCjGcfudGg8zZMTjwQnpv+4+SEqf5BDNeD1CEhguYTbwGFkrSFC9fUeyCbe/GAt
YVVwjXwbR4fEDIQ/O+9YHVOWuMaP542p4LDE70TDBi0mu+YRQDjU9dBA3rty+vhNAtRBdzPZX/qs
Lz3KmISfksklDrrvEPiXyTQa6SW49kT2Xw7CcYi3Yrhk/uvnxQ9ut8X+aGfoezO5VXHIBM3CJT8m
PeoVW8heWLLRnXi9opITBao+GIf6qeJ6py5vTFsUznkaqcAQ2UOugLmowt+BZQnT167QgbLqQX25
VDld2xeqqop06Mkd93LUEYExeVjE95hYYhq0mmDIbKlXVaihzJQ0TLEig6JgX65HoHOEBsT5Txqn
rRnpmTPqlwpjuFgXKDxmQC6QUR3JWHi9SDlX8NkTt8Ql74QTX/uQHlyVUFevOvEiOE4aWQ8jcm/J
r6jeyXGVxcNO4avC7OOF1iuPiaBLKyd3Qh1JR8TixJTxuiDzfdEulXZSRf2mFGrapTY6zJmgGZW0
AOPhv7yOqzYCKKC6UMlNuOy2lswaM2bmaZr3hIbFEUS3sheNQnLzxMu5GaZuD5qEkNyGdsy51Pwl
aHdRizZ9ctGO4aQK34sgmp+p0UItSgptgkEaL+jX82LgIJEWepTzKs+dMZyrdEYx68Oy63sV9BIW
UgZCO+De5VHNJrvsZ4euitb58yhzCct31kxK3Njr7EHOpHVgKNhLtCeRkDgD3yLJHCxEw2wl8SXd
H9YkKztVrHn/ZaD0ItR5YVTw0J1d8cz+fZJJB/Mly1M9JU6toDtPduCN4qokQE8HA/kcsltQVY64
aqrBvuzzJb7pr+FaOIE4lJYLGpTpvJB8pEHym29b5iHeTtC0SEBgMdUwJVKyzNYw7yTO0NlhqfUo
glj5gG+DnDxK3SDZ3fu3SJgXbaaGwINdTv8lJi6Yb82QTngnfolVfS39x6KZApcbNt41fXtA6u+9
8WzbJjJZf5xGl3CcP+jnir2Akr3o1bqoIBtnuAJ7WrtRG23kOxNevUrq0VunbCLd0W8ROzfE6Psa
w86Chx/W4OYcWzBhjrvk/+yy3osmwI3mr1jFZ9Mb/E96y/FKRJdu7PAZ+nVga6OZgiUeGwrkj2zp
aRv+OdLJLgu5sX359TMTcU/OzUNA5+qeVbD+TjNRCFOWBcKoifpv5j2mjcWyuVMHILoDyldx7S+H
FeVm2MTAG9vilDOpHuiQQyeyU+S/2AodcRfTm3xX892ufI8fesimiNRJfTrWiEZWJCIuykHza81U
9Jn/BkBEHYfypwTvz7OJJqF7d1veda9Z7QdVsDJir1k6MmuydilmXPCRYBvFkEWhTr0F2YxWUZ8m
tWqKd4avP2VEm8SbZUExceEJiVyfPC6a5mdC0E/0VeauromCvBTpM40RNye7O8bDMeFy9b72jd88
XGApbvzeKAlobRWVIelER95HmTbf5XDWVdFp4fUi1u+5Qc+slRhLink4aXvwh3m02P7tTXcnHWEx
DStfbqWyRxGcfVFwprSZWLH6hosvgE8fSNE8cMY5thDhMlPCRc/4RLgCuI02c0JgfaQw7sE0Q06u
6sld9ndJQF3p0I+Zk0vRjmUyMm9jCqDq2GQc648YBa18g3mIPqkPaP0WhmUsLWip0YdzRgCh7dIV
BGsIPmFvD4SnSHofuMgYybbgy9JkQtNV28xsbLt+4bsYoONLrbtuMgXNbj1ZmvTiCK/N1HlOMCi+
hT+9tJW7QpRQ8OuzAgOgtjBINUxhGsZ92pwfoUC03/iyIGxRcvwneWA3VNMac53TA4/vJ5SqIUYx
/PavBimsjMBHz7WIUAh5eCe34TNPUIgXde/bt3IiJC1WGZ/NrpLv2Yt4c0++riQ2HfYs23Mnjx1M
hZ9FUFFCHasUikYe312JZwkXwH27Il9flhw/oHbNSRcRc6CDz38FNyxW1SIKoNwmUEeBQCsWvjXI
NgHIr2xLiwAGpKw+pzMVPvqMeG2Cr/4oQAS0XeCE+WVCnm7Slm2seatd2uCKzfnlL1//+RPP3Z68
ZFAi+sXHE7qcpPSLmH1pR6wIH2Q7sD3+6jZAupt0dzv4aqN/Poy3ndf4cuY4FVARtZ4TlVmbfmvv
GGR350r8I/lUX19FVRtvkB4nIUtCk77tCav+jH+yPOC1ekfn8y+Y1SaZEX8Or48uvXpTYMZxajgd
tJi+EYwCDdZfsLiUJ0Wo8l5Hz2/ZFMxXYKkv2yG9v3iGOB5vh5w0g2UVlomRUEBm0aV506pGgiqe
47a7Z+9QGgvvRr04RONx2RDap0ggOuKQYL/Vq9oQDrFmd0seOwBtQZjQcpq7Q7nSezjekWfUiLS7
q77BQ3kZhlSx6z4wQi39y3NDEmLs2kJ0cUe7H5fvU591NgRIE++T29iLa3KSJ0edGkeDap9KPJ6U
lznEk4sYOu2LnQPH4tqNgOcy8c8FpxYPQv1FHrOUnvpndB/0Qr2o7EcK5hxCHUyxF2bwKRloSqko
2/hrZebfl//rLV9PZNKz3gKaSiZCoy9zx5J9uZCArhXuIzoiNJuhQpYCZFlSGN5JK0DC4YdNF39C
Dft21USeZwsbpEAFDiePpLZTvUNiKKPG8O+vDa2WJxLdrUqLpgJYGJKSTb33zDfufNtLXIPkCuiX
A+zfG/AI0NQqEScczU7FBUe0eA8Z9uYAHqCVf+P1Y0JiMBiB6tx7xTmEVbuyKCrqtl6ejSHBCbib
iJf8q97bsGhNLGcdlM+LXMiqxe85PL63VVhu8OHFIpfbuijd45cKP+ZrAtZB/hfLEX1GBoqsLK8U
7ZzUpAnTrlk6yX3O2wN4MRiFZyFffqrit5qVxZmhkglA34QJuqVaxJWTNJvlLOiD1xa0oYep7UYO
8iNVfZ6NuRgxDwxuEpTfObWvywgH0IcT9h+M+6T4M5sMJwFhuu9pRSSeP6/MPKnDerD4rmVOa2Zg
t6ds8pr6EwtiT3SeqEO67Kok7ee098zwlqfrhooIUbCntTopoBfplUnReRduqBW8Diqf2st8DKVs
pYx2F4aUiIEox2paoAYBNmCvrHVJUtMXkfVbkdoMzCmI8YLx+6Z/OG4zAI6OhrECtMLQtFmpwKPJ
VP7DBKhw/0orrxlM1B9iRKslvHUCdAsndi3ohj8he1L0PjsUod1lbV+BdH48ItpE6fRae85KFxbi
W9/iege41/MC5xjL9A2lnVGSuK22D+85vKHqFs7g2FlMid3CK7nwhczxkWVgaS8xWJETkPIGd9P7
TCntKswOQHopmriLjRNO+4oz3NjQst3sOlKcxG17yPHgCF2SpDd1YZVfVheMv0RJyMpA0SikHeyW
V6u9KCkRh+SvFNgGvIPuCJtw/S4FYju8P4iooznoT69i4sN5waIUYix1FJQNZOlA+BB21+lNqOIR
fddO/ScWcY+KiGGLZlZ+t2zLc+D8zvGUrOxJL839cWCX8pyyvK+V2xbB/PsicYCEQKQ7kNvz65tO
f2Xtu3yMn7QpBBdwjoUk10yMCerjpS//tB+xBSOce8eM8VhRQTLw8gbsFSx9o6YMywmmeXKcnJPh
mUxboP14vG0aH0QPJuINXIYQn6c3pCGnpMpHeeZ/9hHKnvfrNU63dqEN8mcpFqD4ffUnimiMzfwv
gCJVb5Kqs4otU9i0ZNMqg2LkJYj3ICKFCPMTpsqqSTDkcUbtqm5MoVGYKMwxJROqfG1NxV31tShQ
7cshrvzGM1gXGlNXqVgMQywAhKfX3PjCroLa827l6qxwkOjgvQKp5hBljE6dLGg1PFhs16iUKj2z
MTWm5oMkKckJ7Fo8k+ouhcn1djDY+f78P10XWQHITj3jxCvFJu4Xr47/1I7/rFOE1uvGbv0h4Qh3
pICUdcja9SYkfME3UFmV7tCDgh10zqDjO2+y1sveCaBMYaWBE3MO+Zc7Azq27DI7x+QOTumfZ3kg
khicRdhNy2XZnF36A8F3LdIF00A0+v7A1G7i5AsbRQTBIPKTUgGLmw0akuhwelnTo6uYf0zPy2Cn
/DElIW4C4oMepikWukHPgVXDTOdlQe+cmAp2kgRl8NPRySz9XNWEmlQotOJwH6YJDEiTbzqIspnY
IAsVv4jz5WzDDbbPQygHWGsQwtlWHmkeq/mncuNS4DU2j7sWlzjA+/ZKg0pze+cLd6l/v+SWpCHZ
z8nH67IYWOdvFyZq5Tw7jBuROepZrwVOMDtXr2rhC+NzMlsjUi7dd/gCgNOUkBNaRwQMGSJqdP6v
FLutalFzLREQmrHLw/YgboAGUzZ7yLtTBNRr7S3TUKwMVZSqM6BTJq2Y38BjK1Nh8K8e6S/o14WD
CM5mzYjnalSWqlm8xT2sAwNxvPMu60V1EVAxSNR+YNocjzy4eLzFS/MoTIQVvSU3NOyrhydDsxWv
3xGZJ1jrxidwVR5elbupLZKuSp8vd7g/JbreeNmegU3M7/gWOyQVmiFqdk4IzFt9MzLlccUR5d4D
xhu2t62l/k8D/pSSbjRQFMX3oADjH6KEgwpUMLAjEFDUiPOAGjagr/GxczrgzLjiW9EIuIu/G4fT
W9I8pK4To3Q+euUdLHQZqUErk3+91gnYSQM1CLnBD8W4NSIVX/xoLS1MnEeYJk2X9xe2GEWNQyXd
pWJianQS2x1DkWFWnqtbQtqPYymAETQ63/KyivEJB83yuzvDQzb+EGWyTsbA5dnOB2f2/nLAsJ8z
QzwtFSHFwHR1Xe38z+kcjJxk3YpPFUm9BSYW7cRN6Nwt30UH+LzAiRm3f8XaFPhQSJUC4nFCAdfQ
S6XNRGzRQmVGO1qELQQnbskxh766IE1dK/A4oztRY9V4h1WPJXZWwazQPqhxYuota3mcRdrYlG3x
mdPElEGc5yTxfLqseBnP/Ysh5B8StXswmRgbSHe35BepVESLR1fthjJ9k6zsLUHYD7+kzz8f+uej
RLFAMzsiiQ7ldfqVSQWeQEmNwDS2+0ubmTDr6GUgGxxc5fM/hBk79Fji8kpYX12WyawcR/Rjjewo
3X1Lq54Xu0qc9M1n6y8JgbR0bhy5IE9Zq3TNs26pNJFQTdFI2w+FuTR2+dLfY2XOsJ58Nj0asTvW
Y/IEn5MSOAPnWUEFZ2gd07zGuX8Xo0H6XTtfuG78kLwPstH4jFEIXAFoUoHN0yMbws+IxTrGH3OH
xyyRzZZoUFFuYvg6oD/xJHF1aQtfl8UkD5MsBqRIlOCiYZLrcJNxbxAoGl934KBJ9RxkttySNFTK
hh6rprsD5pNPdXqjLthgv2jMjhY00ivJj4uzxoxRUwSKlC6MGjwo/6l86heIAhCRTFj/Lyt0yNCp
HAxT7VAcoumJHm2xWFvQ6AAlYfmQXUQOMSL8X9u2duzlSBhSf4EQILceDP72KkC+pBA8uxlkk6e3
PrMApoi4fKn5dX35pzlVUrsmdDt4swsjj3oz4LhANOJFp47RKiILFmboGd2dLxn/t/2tWe/bS/RT
k4/lnNFbuHfTenwRoRUUaXJRNvfLQ7MOaEVeObaqyNthCgglRSTAJIj/0NphXszMj6dLIuCxazBf
1ALo0FL6eRmRilN6AuD8yP+FTr/0gVjfF6dV67kzqXd1vWzUJESKDKUuyLMfBSZV0xpPmtOV++Aq
//K1FHcW39yAu9e2AO0RrODkGolItn4e7IIOcB1uhynuPyYUDHfQstkHOvXza5D56eN0dSZQR0/x
RKrodSThCQii72dhel2eQ0VflfxCatgI+YWybY+Eq3ZuLuMB1V1sSUbGeUr2CdWK6MnNr6S7JPSl
PNMxab1xiMXaX20VvF4e8mA9RDYjAd/rKu7Dw6woLtWkos8dGngFqJHVpRL1XHXoInw9hGmOLPrK
2taSsT7PNor/E9bmrWByvrVB03443Y6J5hSr/YLd1yzipi5JLt13hbD8xB3USaAPeYo4IlKCq7An
hl6zs+ja+0tLomUYnDh5JK24LZ6VjH0PcFneB48X1HfR91u11nOKEBVKkYUxUILGLsxvIXl+Q/MX
8lhava9htbYXnIX97Z9CZVfTgeJmOg/acMshhlV/6buah7HvRNN0oSUgA68YhlvhOUEVAXmh1FGO
RNzVgYDkLnYIQ4ferrnam4oZusnlDOGj9fcXgXPaZNbpj0OEWIkKYSiKSlelccicwuYIZMTbZv7j
+k3/dcnhP1a7zI08ZRozrETodxT6vZmykS3H23d4bIZsQDynBRxFwDTQIqER0JJL8k2bv0qsWZah
vJdQmZOtdZD3G/9PwX9h3x0ZV3Z7vw+yE81qqkdn2NY09MbbrrjdcN+SO0ioPxf0EzD1m8gl4Tk5
mIUIZ//yJ2QFT6+fpbHWCM/9louRlymroKpsVnGiTJAUK0Ew1nMejWa6SPv7qaqGRY8gQLzBztMq
chmNmrmo9DW29rWOmbboATlHeLuIdPrUOZfj/0WYOyaAAiq3UOVLMBY5yN+kkLudyI4U+rPRVoBT
z6BPc9JsDwQ5NDEvbqmabNLXkawWGi8w9p7ZWvDGFdhUF6mB6Q2ijMFgcH7fu3UrqkTNWY2lFHHo
IuWRHhRluP3OawpA2uQP5/hhj7F0tqA67esA4zuPEMwcJltmIIg8ENkgJ42/g4Z30llXBRazejuX
8XPmT5cfZ/C2lO9bEbzAinOGEmhlr7ZjgWv8FhIdH7w3VmWZhofQYc6vrtetzDNGHgosgYVRl6ZT
3iBGd0EQFBbGCWZeMf5pUHMNRv3qXKzFckxxuqDi/pGVmMf8vd3JWtd58Mhnr0wfLkMOj7Apkuk9
e2q6OGSwmoALtmLJYPnZ2FQ9WhZIElltIABJiNtcvhYoiYGoFOXlC9OEsOSKPXpQkI4Qigtk4BCc
4w3ccAXQB45XQjzXBfgv+AJ3l2yrW8j3O2Q0Px6m+OQszXHKZi5yhrJQwjdUXdEzLUZsA3wAKb2I
9xCRQ6ilIvt/s/rrevIGSvfOhk8v+Gpa93G0o2MHodEstjj9ZUVRPWAya7Rr+wLVgN1PLtA5wF/w
B0dBFRK5bjadTuX+jro38CK3V1s5Da9JHy9zbBUfHTkV+07WCY1PBwIXgQllj6lnKF/TYCZwEsyS
lGIlSwJ+3S3PXmTmv/PKp2GOEq1yDtVYy9BFHI5psGxd5aGim+7IkZlhCGTQ6eYBKDD1lR+NR0P0
L6vCLuUU+pupw8jJj4o/vipFQhPPIUPOVIKEDTg+GULCQHO8KGlrcFFCHmeNu3M8T/RqyZAzz1ad
G+59yHLkCa7x4WM1eb1WpYWMsZfIAj/N0gOxIqkN1y6cuZ5CxZyQX9CHAE/z9R5Laho/HCzdbOU5
vjRt0xDzkLF+7G8St7z9wAMj4RCXybA91sLES0aMQWQ4ebBhVnLPiBq6SB6ArpoQQGm6Nkk/h0WG
tO5uLljURuFZmHfqMPwt1cv+95Wv/a9hr/N9412kUVB9m1j4jWXTyiV5wfdocAl1rMhYW+DvEzhl
oYpkXEmJej+BlyUeQ/pR9kuf6SP/CKr7TaDWpv4gHIQuhrvr/dn/mxc5o/xvAk5Ot7IZ6MYO+kzN
vlL9dv89d16qh0h05JNRtrf7BQDFGg67A/biZuF+6Z/W5u8SxMmMXNsjExIm6vXxw5zpaCDAkmRc
S1uwGNy57cBXNmhBDp/hBNlATAIVrPKXYkKdw7a8vzvoGs2GFDHboo/24IB+Fv4ShqTEiVVILG/M
k4UHhB5San6hcqQA/U6EgiZy4GS953tO2jom2E+Zw8SVOrziR9UFeOJycX7vL3OyqyZUKvWF+Mrx
DWR4qr0SKfD9IRvfTpw4wCAb2IoPW3WV23feoFQhvLtRFWFboVYq3LyJToPDc5zO9Fi9+3gnZmdx
tkMac19O6VcEDcVsTYP4omBsj4XYt5ugzAPW5loXTve1nlieky9bVqoENgGqc00aShA5YGtw2uLD
iaQKayni3pGA045xEECImhhWrbM9ErO1PqeXRAz29NRJDLq1gh477yrCekrZ4ILcJsIhIInGbA+U
rbIOSmJxPrb1zZTE+HvMdgVmmKeaWds/yetSrLmzcPgmV3o6iobK4ySbrgDlcpgMhVpm7rmd49Oe
FtxwMNzq3JMxe7GtN/D79sAFW3MAgWaTfMKiaRDYC4sfsXwjcljQ/S9Sa+FURuv2bt6M8H507N+v
wBgM0rQEDkgm6I+ui42uHFVRxmeCNjGJgr1nAisklq4YkWamA5qfOaaYIKBtqcjsqjxv8QXxNzaq
0eO3Bh8i6pLT4wIwn4j+lWKppMK4wpFPSTBS3dmg5T3qnmzmZNxRyZ4KtqGxdBESQc2a85Y/pA6K
xIhCBiHj+ULl+bbhG0F+Y8Ryry87VXtdNaPz8ndbYmOp+FayC4m/96es2Og9YucPFS8ywRUGXUxo
Fxotw52nlszGAW1SPOUZq6JDYpeSv/LFwC1LFm0GfHocEQLS/fgcPAZFq60OaiCP8Bd7q4VBmafJ
NfUcoojn5fZqCHuzNjJJoQzMXHOxiLw+N3QlMI9U0bIrouAzlwqtwQcGnjvc+S+6+5AtJkshuZi9
/1SH4ockcdaRQXwp5bNCdS1QjhYO3lRLYhTTv42hORJbu1oLoJpdTGdr/w42Vvxg9I0o3bKD3oY5
DMjKV6EBtlZsCH3YlIkhV8dmX43WluNuNE4RA9FhhR9JCh0tVm9n3vadKW2kAsciopvulfW1bvd3
tkes6Iv9jaKcPaKnGFFncmKzGFmWsrGqKLEmqu0FbxECrtaO+nBPFvgxccuBn2QOu4KRP88O7xdf
Pxp6TEYWIapJPAyxJgRPH6MSdqJxegEV6hU/33tAC4uWIQMYtfy/d3VquRqhoVmSBp940WeLXfzv
2q0DMU1//zmNYVYEbMBRu+7HgjLP0WaHuspcd2SF2+dNcnwjhK8QpF59pwzCVk2EDatBZhKFU3UC
4SLvxZdigaNB+FG4p5fuHOWLrj9IHBXdkyvdLIltPeW/ULzUf0ctXkQ+7ueE1cEPlY3KreILtFq7
o6jOrBSNez5+O7oBwtmwB6ro3DIa0svnel3dhP2txmP7OMGNRxG0H+LZZSipKqfYmZ0wL5KxKhmD
Pj0Znzr7gOyaSRhwTPLlWzq9YOHagzYVBP5+4VhITHphDuEylYqYn7dqEK2eFwcnk1fyKlOynHn7
/BBuKE33xaf3TwjAy67hcEjsU5Q1lVZ1vioc7X+kdZ6Y9pHXPguevAnaURts+dLbeToIPfINgSVw
gWc319v0wGBEhOYk51w8MmezxDCqPxBLB0s6/t2cziXrcv6NIW9G2EYUHYgvhV9UBOM+vk8KN6dM
ybhUQV9xUjooFAW5OxrBGkPJv8sPfS12p0aNyOsJgmP19EQunTZaD+LuP3vGz6kZUhuDPN/evaV3
SkHBVSx8VMb6KIkeMr8nd1fIl2OY/wUdiYzV3IrTL5WfovHmG4d0RP81cI5hJRwFWN1zbyQ4HBuw
rHA8f6+YtlbCMDn7dcLwh2yLqZe5pn1mHrJkQwk70q6i/ZpXMei83vOUgNcH3oY7q4I8lFdFl4mT
E1EG1lWmzirTWd15tOlevrRuF4KrzKkc7+JupmSZWFL9t7VugLjDsponCxnD70ppU20WZRz8xDMH
8WRxSKOwieRfVzggcrMv4OuHgp+j3JsxcY1GASHQM338fxXPpVbt3heAwMnkbYh26TduYMhBEdYJ
aOsip/jSkrgqgRd/Ga2FLC+G3grWE+oGEEq1Xi4hfeq0cvP+JtjlUAq9BiXzGGIcPSQ/bXNYRwr4
++xEXBEaDcb2xbxBIQhnRi9DA7lEOb5YR61wthGZL4AtlJu7wFZWeMot6FtrT2O6DUXd97pW2fE8
/XgUo3yJ6hjL4rDPf3G9ECBj4zA/TMZwics1u0qAHvqDKGxr8bVw1rsPU+IUErxMRsHit72si7Mp
bWwBHdj7dEPZ4Ie4E2/c/KvtJRymh2zzwniBquvbzNcGgRV5gkFDbSFJRTe+XfzYav5QonvNwioG
Wf4gwVdh2NndjO9/kaZKjsjWwCmAvNKtfU7WQGR5kilcg3zN3nY0zvO0oJ2DZvuDLlzsS2+lnoKS
qdcTIQLGqRgkdUAL+V+I9B1nKtOdSCPGxRJgLmuAja0axEQ5DLr+I8i1XKWj0PDbtemlmhmvOern
ZkvFacMGpqw9N1cvQyBDJg/L6m6dLZUAZEQJG1KIkTPql3tsCDyzq0eSVDd0Z+6wn9EgkhZQ2b+E
FfperEP/qgwwlYxoGDQTZzQJ8Z+aUTlSCQBKf7Sk40QPBlwCBO5EpBFkdQIwGZp1YAOevI3yNzIx
PwVd9HLiIgIR5xosyMb1mt8Es6V1wnuh5HWpBAnOk/7qMaYb4Xw9tNkWOyfr8FB1ioUpntZYxASB
jjZ7i3Luixxl8EdFXPnkA2Li04exLJhPtot/SYld7CaziRtxkRdIxzfvw6/aMmgUTsMcI+ESHRJL
UFQCPUWhASbmI9GkJx+gW5S+8+QPufUeoUOTa4RQTeBMtWWC2n5DQHDEpLbZ8IRcBoVGQHu8e5+m
2XbiaOwtBZ7Z7TPDX+tQAhhXpzdOxnvwPblliK2kwc/PfcnQ/344G4roGOjazjqjJhHskyYyOkKp
A/5SlLVlpuL9cGPRiZTwBJQNg8+STTRpcWHKOmFkd0XQ1919eLBzRi5L9ji+VHOxmBe9+XJUKqEE
QPE1tZZgZ2KDrYJWz5l63CZVB9E3osMyz2Gin9OK+Tw4KGVdtcdp2kq8vWIfhX9MBHnoWw/alNDT
oiXgVX8hjCqsAiC2at2Sos1jhkWYj6TXFudqFWszCL9M/RbEc7McwB1Efo1CpKVKgKNYW0SuZSx7
MWSVZdSSSWM1SZN6GjSFFexf7n71v+LKnJ8uEIbE5wWLj5xGLq+GvYB80WmvK1KXH7d6rP91sk81
pmwrl57p5WHGellGhDXfKfOssrod2riqzdpLGJNBtmXbwDO+tP2GWgne9zqsNXQXQ/rqNuTSyRrZ
Kqk4T36m1i+UoRB0UbTF7s7uPDVpi4Z2PDRSOwM5SzujkC+fiQSz3iDuQ/jT4Qv6GgB1kOpaBZ4V
l9lRsL5aNL70BJqJXWi23E9HMsDYa+v4q/TREu7sR1v6E/F32QKPXPyYoDGwJJwkk7YdaBG02teK
r5jFB/sfDlfsTszo57vLjEK6FlAFmU8QhwwKh/Dg+YIjS4kzsBk4KZVKtUvbcFQPfstGsG6XIqbv
SatRRussdPG239/wMcVxfjVJBkua6C4vp8pnrAZNWswPuuuj3EOv5w6X0D4YY9fW10Yxl7ePibiv
3MBs2S62nwRS5gQ1mHIgUjDkFBrtFvnzwC7aUJhp8XH5LXlkJ36SP9ynMf07wYS4BuIFOA3sDmxd
IdTaWUO7IevVsCM3DXRRSvtouh5D64FsYVakiPRLvBEzNCQqec4LwSHopwMnLne0MOcTovdnhujF
AzzYjAJW+Xtc6vOg9yFjGnXkcpzhWB6hhaJx8jkZGYIRqeymxhkpTjbWQR8K6051hM6oTOTcAwHw
K/etw+IoALCFtQ8zMeVZbwUcmK06Y9PMExzXci9fJ4EN9cpK+L1l5G/rWz4D52OHXvWgGGkfkyjj
2/vfZ/dDxcw3wA8h5bXWVgIBAiimHl7bVGQdTUb4AyjgXoWW/HuC8dWb2FiuHhPXGlGKLx6hsTrs
Z010RRxHbAy0LiRqkCKf/DfciJg8vpFv0IYLbBjdBK0CvAyllaAv3lTGMRsi32wfkAUIZso9i2xO
nvJFiS6C2fsIcogRbDzR9r+LMGh3xXHRYjieMe29RSP3uq4Vk68XotyQhqURBNMWKjU3wARpHSvK
8j86BYsNjp0c2yo3n5ns6/ARinhXROudGFkSSXKI5XZWAmaSf8Alemj6I3NC09S4TnVoWfC6/LfJ
Q0Q14OBv6lrFsUJzAsH0cKPJ+0cpDvtYg0MCpmEbGIP5h1KwlTmE0E/b0IBbU9VnOVPoAV2Hm4kN
hnZJjz+gH1P1tUBToqFRphMv/dKtkP2KuKnKnn3l9scTMp9o5gEBVwuD3Uf8vBGba+d1/fcyrbmx
xsJbz1nQXZTxoOq8eg75gSDqynyF+HFI6WnDi8thUVzRbp32y1tuceuJld3kvpTmYIA0zkcxvTzQ
gZHSHI6fh+gOk4oZfLN+sBU+MUP/MoCyIiHE6mCKngTLwvTQy4ribplwTgW4PscQdmF8Rzvbsu7d
1MnyRnuzqmFaDcRGCzWfCspu7W2DYBKwuiG0yyYFzj0wRJu4DKCjkRhVanVU3FE1OCNxQAvutkWh
Iv/lL7gPNYn4dIXW6m6wRmfmDJsTlzYUW3rAbvxsLQD/7LymLgHOG3acrf/u28BjgfUa9EePLo4T
Av593aPfL0I6VnXm6iBVnSQtXxHCnGP656h4YGDhVkhmSDY6r3FDOXbBSFYN1iQpiyC1i9RXJcuP
hGPjO3iS5DB35zS4WiWUdyImtIJt68lUX4r8kAyjl47103sDIbL6JdYJXB+WCs5mJU9mZyRbOeNE
XH1fXDYtw3ghaWqvj4LU7bzcIskckt7/3pphP1N3+JSs8BjL+QOtKyV+s27KDkvsEkQj9lCZBv5f
oIc9hRSD+Jm/uyxtge/kqqh6mFW+hJ6Es+VF4e7q4O4zKznp/lSxP/9I1MK0hMZ6U3yZbHu36Jw/
FBoOu9g/ffkM8JyfGeyiE+DdoSzBazXRNGlurMMP/9vbw39k36gAMR16M3WOga2qFw6vbsaViFa0
Np+ST7lecUn03hYJ7xLa0yfaXfdtKC096qRSBTXJ0vDW2ZaWkvHPnTjEOh0wsKvjDXO+748B+dHM
eTOD6IiIjwFeAkUVfamaSps4Sdt9dbTD/SpVJJt/unip6AwQJflyS5OybQfahzFivoxEjqgcRgkK
PK5o6hifa7OW4xRl7U0TwEO7QsjOr5D6oqoWee/2Jw1yqljAfo9qfxKyMeQ4WRYVT66I0o5Oth1H
uaZZeDtbXvSFoZr7+xthbbAc2+XJUmLRUwOrvOn470Lt6pAQ9XBAqTsDxeM1156CWTClwcpUeKg0
VR95oK/Z8kX7SpQO5yh10y9GVjBRU8hF870h7BqG+SNzDDVEtsP7NaHVSmNGUSsOkk/YJZScZ/nY
9j3FdHXpzHCroRKRiUtAw4txzFNQbJmP2pbD9bpgePhmdec01+GIq29GDVM3rLl98x9VWc+t3BKE
aBFcmh+XrefS61tkyvz3Sn/f/oCVr98MAGAW30LQW0v0KocR/R7B3nsfvXj8o/ucRbY7NUn9FXL0
8MWCxbRQcZA/Bn41vc1QSDIDNXI4IQ/NS8gbea3r7/gJEBJ1qmsihGDUbHnxsiU0txPCFcBtwZr3
JMxxtlSl2lyPidV3ROVDKQqHgKEh2JF+Lh/YiQeTMHkaIs58fsD+s5jE9q5r5xZzwLVxVjTXX9gT
uAth9YVzXIUgoDmn3e5mdz02HIlPO20cjdzF+6nNLuNv9dRDg07ZFdKg7s9BTnzgFgvryoHIMbpy
39VMoTSYA/TytEFW06qiQh4zipq03lQVMbmjnIJmwhK8oXp752SY6oWEit0SP9CopZ+NtuqJbSE6
SmvpT4Cs4qZGM1muNqmoLWacOBz3dT16FEb6fy2Nrn2kYQm+I5TJhshEaAfwPXIRlZAB07FI+8bJ
9rRTnk8el6LWs261kfXrrFo/vhe9hlYbCK2df+s3mSBvrKo+3sYngwkzIcw60lz4NZJQgfZNpiZs
RIbuEm4+jSSs7c7m5Tdv0r3E3rAKCk7BqyIZGcPtjw2IGLyHEJL8h21E//hw/bv5+781zgK10WqQ
3fMuwhr00W3q7giaEjvIZgRL7V270j0QSWAwo5gfeOGT1QUoxYgkYAbnL86sFqOFx3go7GjpMnVk
5wmDsXDmlbTaYB8zG2Yu4Ta/JFk+OqLlPxTS/bQothT9QETfbNdnbQe64Zo7RZqW1+rJ5PbXST/V
ST/c0FsCYYVN3ARZA/L7V0xGdJDOVpMEDwXMBcd1DJB6wA6Uulf+M7A+dLAOVzU0OvvU7pC/AXtY
oeM75Ue/CFKzRON1g7bPb2ERmNsPsuT423NUcaVwWnz8Z4hoNbTcmHJjaIXMZhVyBM+E5V4be3Ga
63Fix6219L3BixPipnov71bf08BAHDIua8exx0c4B73oodKdUQNkHxxRio0nZnM7lGmNeoZ4yWQP
v9VBpKGYi/pm/BOBZzv/fvKfhaH3c153Bz3W40Q/EhfZv8MZCkIGRHEYnW6JDwcoouoQ+7dYuu3L
Lh2t5Agl/4GsC4lmouiTiGeQG2o7RsmRKT2AVJkS5wXyppeam4/ZqYpRMMNbsf7iOhqa71xOL92v
9Z0S12GEuB932jvZvvJB5NyfkrZmhraIKxausoxLrH0ODhTZnEbksBuZFnBSQ4DgoPCk/H8ENJRS
gR4O/ft34H2ZM0ehrMaATu1hkpRjMikrejCEHjGLPmeGFlja6aha6W703ym5g5Va+o9G04OxhQnJ
hfuTLzX+p+TbxfHZ5OKlpZaotOpIs54DRFELwKv17u8p6/ddy60JhwMKZVUT7aIWhv+T1t6TO6dR
EwpIgrDv1/i9urj7XCE9wWpMiyKqm9e41ZOq/xpFczVQW4O7J2c8zflRk46Jj7n+m0mIh2ETu4xD
KXUtubX6q7TFuVxizOvbfPOY8lYV+uN0rbo6LheUeFdm1OhIR8anfaLpxFxd8kR2W4fRw94TkXQT
h4m+lvhOajqWAutQrW1N5J7xtYjjTsREU6BByxV7LrafR19rqtQQpCgzoRBw2c47NBbTCKZJ6doW
5WgaOspytxmAJi/GYBzVdVeHBdjEYGUD5vkqkSBQKluYVskqSdgLlmdOaxX33GpjGsYPXvn/WEyg
VcVObeJ5tKw+E/gVYukNtVm6rYOpYzLttxlUgu+OzHU6yj6KAobtKBXW8aXbpb96RFiw6Eupjetr
UsL70R7ClwM6bwgJCDUZsARcKVMIcNjJMGfVkorKI6txhNTKxY3Ms85A7F0b0xEid2JqGIAeZUsn
KSMjS0YJqrhxlITGuqwUri/sK6Bwf0RM84/hG5vjqvH+ej+6+7cTlwxq7YXzQt1T3XF+8pFnr32/
lgvJerP0Pyg9npDB/pnoJ1PIDNOpQ57soUMYrMylOTuY0AnBo+qDlqoPhEQoJJ2H2RiSquVzOJb8
TlH5c5GBQI5dY4/UQYuM+VivxC21e3LpMb42V5WYl4MD3zVsO0p5VcRKZyG97Wk0OzlxtG/7lhdt
SSDuyA4/oa5ieuuDV/Un3rrLDONJ2jNIXHTK0pn5Hg437ud0Gl2fssgnVwANfKXwFP6p5OMm8PXI
JqX+b7svYl6Q5oYeORTKxMLDehHXX8XQFGrQ6WVlnsQ0deaL0eqwYjabCNXFJnqo833nu0YDb/n6
sEA7QYnJ6Fu5gU6FsBQPp91el3Qo9m/EH5C+kVOSZHuiq/+atbJyyR3pN2sx9iBDWWNg4nqUQmzQ
txdkSJKJKVnLeiORDBF45zAXunKtbGgjLP2tZsLS+LB8LF48FTYsLD7I8IeSE5j6hhLB7tbDEBpI
+bdberGD+POkNlsqmKcK5ZgtDdVddHplIyp8CpRklXgzke1rOs5twGgtGdSi1YWri3kiGeV7xVw1
E2LDo2a51o5t9ziZBVatUG64dXskOhtwjhAoZeM42K3loXJxehH9cKe5ymA4l3hCINwtWIwVtxlA
PKEI63Cbh19EPW7M+lq8iJAx7fZkDpH6eDAyjlVcMPg9dhDmVYRtFyK7TOX/fnQwTLYyRiFX12jy
I6yJdCGFginPz9jSXlpVkWkRSukxtDCpllauwrM6ZraO5mhetpU+x2WBQ9xAQfPHMkys3mdVocYO
AA98WqGh92BtQAlLPAiCHaaRW5kNXHNyqEeZLdzwXz9+jKgr6CxFn674lwP6l1wdn+RvKZh0Xyc5
9VrRI9E0mQ8bawhZGlv7W2/49VGE1o8h1Sr1aKRGfGPZ6WsD+k4eujAL2Kpz1lakb/Wefy+zdK4X
MwCyJZ6TCi4MOLc+LiIb0235nlykTSGCNicxuahm9xRt5U6rDDjXib7OEy7fLm1omvuB9/qcOJZy
WjiGnI2/Ar7fvzIW87HgAg+h6c8bGX2279YNzTAJDWTAB+Y2abIeFuKqHmYZm1eZQLRLoVQTeXx0
QsJODKU5z2ropk8KpsXcPBavQtM0zL/+jySWiUaVumnulpSj5HFjuBQSahAoylf7ltkzTXC5/bw1
dTi+zw91cM7qrMcdxApY+E9UT28Z58nNnm+3DX9K5yALNXvTsTDSHPVPZ57QV8r8eO5VQ+VsaDa9
gaYUb5X6XONsMpa8qPXU1CuZ8udEdSqZxHQbxP1PDvj83/Xs+pnpYUl26f8bhgwluUvjRGflnwmM
9tl0A/GnH37uijtLvmaujKfyHU8D61SrRZ8sEVsVbNYUayIOJEEOIKto9fvO+Cavg57U9XpLa4rq
tvYzy/+w/Al+CuN5MNRZdzXg+49PjqirtxkMbg9XALhd8QIEyNuue8duNTgpVQ287tn78LZGQMJm
YsIMizb8LPkAHQDpozM5UX4JBo3i1IQv7lsFDZhELBQLOanfwXS74EiIznefiY9Kva95AcS7Qj1G
PPsj8P1I/qwcrkXoIkIMAYUZcb2YChao8LrKSz0X98lx5Jow6nRljQqgP7+WVtMY57px7SDbFORD
MrAo6Nw+GQlqC4lnsk/HKadvQ+ssT7+HB/RW/CB+gV7bR/Ve9+eTsNin+ldRGz33Gyi937Blk7Ck
4/zW+KTFTyeM2cNgHdGcHe3l263DZCC5WXdU1TJ9Vbk2xS//EeUC1rcaClgbaMd1wTaE6IBRX877
8Kw6YmF0Nc/tG2ERwPrX3EwAJfDfDowNATqiz4a8zraktjm4Z2LhyZzv4Hivx+Jw4B62eXRDprKg
L99RiRKnv6rc0ynNNX+0omRkYxbvbQf12F7pFtL/Kj4DFtYLlX4yF6l0uZQvxnT/OdRAdMiFun5b
COqoRd3D8YhO6DcHxRowMDxrl1TFtbuNhO+8AkJp6+Dex5KN9X9Sq2cCD0LbA0sUeTKoFe68vqQ7
fF/f0QtI6J73QEGiJCQk7buxfnadwstyY3UPisH88JKZ2lx7oBaTIqelNspFypf+7duRscXaenrn
3YjsyvML/1zVl6f2ZtBuuBQWlp+BNHGTo/r818MIYk15ADYSx6SMws4rw4t2+86X3I4qjCveWeEC
GvzSI6fRpLaFaKZoM60felXfm1VOt8ESj81xDNibt9qd4zTtmVSYEbNilONf/ay6DOv6gKeXJLgq
3k6s1mKPjxlEidfpy9F6W9ag2+rwfAmtiX/Hb+P5PhINf/70ekw/ByGSBdmRRbDKCGjF5NUp/3jM
rlERVv5kRoQG8kW5Khdn0zmxBopGCZFM6Z75bi1PzmeZuIAjkxAkKHAA+FDnQZIPZI2myzXiGdun
/ktmOxl+/WrpmYYnKfqE4TYfKGRDZINMltJF5Xm80FhlkoufVdq5i+AiQKXrCn0ZzqMRFW0z33Sn
MTsSbp4XgR7QbpE142kgmjf0VxKqK5EJwmKYPGdH32Z8ccodpugPlQdT0cNy6NKNtiXI4MhmT3gI
KVvx8I1iXZbGbohAo+WAKUBXPem3VIKtGvYVOUh+5h99GxoGsNA8xeHNO2FkAeRpLIdJMTbmAXGK
JNK2JzfsfWas9z7MCuj68IE1mR6B1fBGvvzyvkdXDH9dzZsZT/GahXNXFODglhqpUVcXCFKCaRTi
HnHTxvh3EGjXO2ZrH+D8DrEi+2kUkl+CK1dKL4QvR9qWlpaF6VVMQApoHgxf3IMunbI+uD6rFDct
OuHOJmAhrCzhIXhNgfFGigSNafEVUhij11y+qKhPz8PwB9jzBTwq9zU6UYI4i9IhAmZB0adx2j4d
X3XRl1/qEsgAmdZMp93YYVcG5Is8WIe/ce3XF3DqaCIgUBXXGlz6nwULYp+HyoSykCDw6aOVzKKf
p5/jSIC0XtnMboOOnVfs2BclNtFAFnEkywzDJbAV2hgwBL1sLFg/OyUx7ZuyinPWdoa4pHJawm49
BfWudMdpl8bzfvMVX/oG8c+niGmGOGyajlQXehJpJp8RCRY9dqRCJVe9jGrx+gn2/SJpZkp93KhZ
OEnYs4xR3WsU9lxIV9A+ouwJcogSFjjD628sMmm7LY9w4mnkZ8ghl1FXvgV/Kf22mIdX6ru2x9/I
8q+VmlaW8732QJ36DojdB2ol4arkEOZptcQUKrbj0ciMSEV6PiJxRCGxLe2FK053V2YBGv88aBa9
Ee2EYt/07p+J65I7dw6KjRRGDqfQaGE0QcvGbVrcWLb1QmNmDKjURON6OH384OhcSbILqjO0DBpQ
zjDWR4+67B46YtKC0wcgxIouKNKVx6oZAjg6j5lGQrKyqbmNZjV7TBYFfKvAFzOxtu5gwNwoSsug
8HWjGcLuxWyijgia3++66xHjs6gEvBAyTJ3kfELAL5cjgthJlUCEQJp46+VTThDvsao00c99xDP2
5M/jnbbWBfr9/VPB9oX+jBmRE3DiR9wd7dYF7Cj0Q0zWEcDTm72r/Y7XvEXXi6RywaynUjk7HOBj
zLsuOqqqrnsyTx4u/8RNgnuPSHZIljiPYZaBY7l+4bF6Q+BPyY/1KbVxhXzsJWfUXBIbFj6uLWXT
5hKhyvdYbvrVLQCmEE4kE9GqoJYMrPv4VpsvuJHV4Dmi3WQD4ta8UW8jyCW1BoifO2gPg7y4sKIE
5vghn6JCKZOF2zP3uXf3DtfNDGMU/CYtNV5ExTU+kqfOh2tn4mzBJYBRA5oLDjaQgd8lUHL6q8wI
buHHYA30AwD0ueQLV6fakyUgEbOlLWFmT2B2w+UjtHGzvxVU20/z5UN10OG3NU5zqCa951qEpk4d
u5OrtixUVJyXpESkpRHOt5Ublb2gwkjXsUpqDxSem2sdf5n0Oqe+VhZucL7B035A449QIN8ieezU
zM4IADNene20dYcayGdtDkaOJI3F0ouL3XVorJOCx5DR5FimkpS8UUVGWltcm5xDoBQ+h1lS4igI
/oXaZzOxMRk80TzcQUC6+N0se4Arw7SD0Olc5ySMP7ut4IHyKy7HIp/GCLDGmJDuVcvDnSa+KDnH
tAq+34LrXcucNOo9ZDC4zci3DTPum/4EJ7Rdor7sJ4gU3Ji+M85rhhiCFeOwrMG5BkhjNIRHSSfC
C+Q9bdSpzxUtegh3XXqZgGLgN+uQvppj2kz4URRgUwdPCc6E7t6kcraKujupyWMDc4rxyWiuTOo8
NYskJ0yhKddU5pRXPa4CHxDr0/4LkucFVnH0foDJ3lQQO2Z86LZxXkwz2zLAaoWEnRviIsvBLrvL
R51gvJ0xin3vjsn/BREehK4SiO1Jafxq1yMdf3y+Wq/Igcl95i3aZYuWvbCnK8+DFy34T9mYWMNO
GKgLa5BUCq5lcnXQDWrBeERZK8WCzgfOIZ9jSd2r661wsumZgJZgg1oHLqPxZDzdeb3+pTVu+T8J
ODA2fvBXJvY6dFEaJv+TASaE61NuHbDNzdSBN89/yEKkfPF2i+uEbqH5/cQNy07yuJlLzxiGzW+e
DAm9LHvE91gFoNpYKBuA96Sw1GUm+Qo+A3eTCiZqH6t/zRx8awOvfdIj7tfqtkb7ONxeFNygNo9q
hE3ShEvtHcJqiVxHLvWEsRynL9oU5kop36hA/COUbK5DsiXhMyi7TNf2CKCgDc6x/TXyfe4W/WL5
yk6DMZY5Mlqk8vLHU0Wgck7a+b521wt8D4dNwRAQfVHXbFEZAa3MtDr1uUNGMVLw7h1CaQrLL58r
uFm7SmYUL9hgWVgWeFkf8YHTuVR82x4uL8SDK6dB7YdW8TdCGgp6fZuzf2yutAnqp5WgAeMID0J9
9XjF2UT9R7N0dd4c1kfkvTdISfsA5OVggK/e23IDKILz4g2kTPCBPVinDtZtm1cub1zQCIm51OtU
MAkvr+WGTHT1jSSrOCQZy+s0MdHUFXcXZPYUFkPX3PrcJbgCTqkzwlhz8IFp8O8FOrcW7/F01LSb
twzT6GN416peS7NpMepdKNi/T8/xb6woj4G8CNdOSFNZB3ZNjzrAELCnX7XD5X5jd6OlxzQ2t+2X
Xbfw8Os2u7ifj0MpxoYZbSZgjNv29IvOGvljsUtINM6nVyhpujepra07sOTpHqZ8I++nqyidcOQJ
ReCC5PYwpd54hs+0eRoKYH61BflhGLsmS/7+GEbbWQkwlIt3p9RIiZny2AA/HqEgtoUi6LBw5UMT
0MmIagAoaXt5puFIuXqGAqFOU8s37sAWA8iCFkIWmktB3EsOfrayn9UEJEcp1GrNs6bN+EfderNP
7ekTM3k0mq5HmA3x/p3iapN7bV5bl8E9DzMM3H0w2x5H4VOKIsaZyzf8EjniSDT9RpK8hALZxyzP
O4gVl6fDJfclWYs9cYdQ5z51Dhfocltmhcx/dNdrO95vHyJqRVulbBVPkVYaWjxpLh5r4Yid3rJ0
V1MB+4bJ2Ht7V7M7nXOdCE1km5yx6fjfn3krhw6FMt+f/WyRqcwYbMSkjYqCrK6+DpnmEweDeOMY
o6VqAJE/rVieneH4uGgLwaOZLkQzb+XuruDNEC9qIqsJ0jvSNTnoc7Uz4Jbreew3Oq1KGtpUQp0Y
09nU+a0CMCOr4rj2DeX1e/WgamFolxD2TkYzZu9hq6+bqCvAU0Dn4ftTjp1coxIFrlYgOYE/yFxV
rDA29PdvwO0QnsRqq0YygbzaQKeuH1Jk68wuXRMc3nH0n3Z0yUInanOCf2R5Ig+q31OnHl7cw5My
tAOFL7TULcj5jpepkAPA8AhEeFjZkemwCFKgee4+dvASD9Izl0Jp5ZvQ2pOKBzw3tLyXXew/OzIe
kBDDDScuF0vVWFN8stGX/M93JSqc1abkczgkQUDOE16/CEcg8EDPbcXQGA+cjoowcDPGP0XUy8xb
4JcjCtbSPZfmH4vAn9q7X3ySBVSZxOduykAOXh5hDXPWu3+t5en5V2lad+Qg+KWLgyZ3Y+SjkuOJ
ch45uqBJ7qi4YmLsvjFN09R10AyPPkCDYy7SGojUC05qUR+FlxIty7Ox5ZolskH9b94ayMzA8k9/
cYuiXP0TE6bHPBUiZYbBSSrIS3E/3Pb/RgY5ynD5I4Kumyen/pjlTnGErj9f4RS6obPHnOmyuu/k
xkAy/NNls0RSy9x2VrbXlgR8/gVXa3cKRp9lBKXg9G5djiitBHUiUrx+WjpgWs/cmDzMIcRngeve
Ga4BIHOr2tb1rxMJTd1TOctO6oygSDECFxGMtRqdrz8aZZc8boQEu4i+EH3Dd0VUTN/agh/wn7k0
WfARJLcGltrfwNtAtkQ5Kib/jX536pFizJRK60kHgslSajRJOjwFf6JW21vWv5BkXgZAY7xWPfZh
kxFpYVojIdTyM+XoreaGn101jMq8g/ou5hTfKr736dbAj/45WomaGt289pLxK1Me7W9lrLrAHnpQ
yOkemMMjdg1cAdvii+vSU3yZyNceH8jduBv+ELyhi7vChc18yxj173QUlzv1D2Rx8aWCelMCBmwE
DMs6o9bRgGm5r4kVYLNiVtLm78Zuh7mzYHDJMMvI/JtR3qSDkodfYPcqlXNGc2gokq1LJ9jbgsuW
4+QgcssMq+h3W4f4jlrVs3pbjXhFQPMo/s2UzcX6EE17hcDiLCth7HfiefKt24AjbUZ3drF5nVur
TsCWIQ17u8Gn/J6uuenbi/4vJcxG2fdgY++odPfgFoAw0Dzxdgg6gi5he/GFL2bgk3UoONqKhMU+
PbPp/1zS/bSvq4T9oRnT39OJ/VFhPFsDZoExYBNq9C8H/P6e2/5aYveYMud7GCn0alUUJp9q7ck+
eynonrtmLItU6YmAcbJPMLgXOFLd/Brj0UGnrk4YLCT5+rOYA62pucG3HrOOEmwQhzP6hmK5/I7h
HMpzOQ5Ck4X+5ulbj26sinltd3RT/FYpUoSdQlQf22QTNGdnY35siivOxRSnjokqXmN/2i7pf1hL
0Qrq18woDdBVSouEMI9B4YUr+H3+ezbSuy6D8rYmcm3+q9ba0Wz3LwqAHIl33bXVN1/pRUqDLwj4
ZURshTSYAPmIlu/RTPtgpUOd1+4Kr9mv9nk4cinlC+B4i3Vqfqdz+lDsKnUUK03lfzl5qkfsavGR
68OHMKeIrmfG0khf1UCBWTcpGQCBA2Et86/wsCn2zjH+reORrHzz6Zhz85J0DkntgXvP1ktAS8CS
e0wtNnrVHV24szWpdw2rz3i9r2KjpnBgqHqF6A44sc6Lrm7X57Nh8haqrRrR2XzM78lHw8rER3vO
VoJTJA02GTMtJ5LS0hI+6xHzMvzeGwD6dj8nBgULVFJlXukN/YOtHlV9y2iIMBR0UV+Agx7IlbSR
KRD48ZkGt7yQMcuweSD5/Ib5J7LyXHHfiTVClhZVBg/rOf2JMNCFTR18Pn6rBxsn4gnOAAlFgMh4
Z3ugP96nMmeQIbUxM00RKrYrx0HXBuYhA7aQlaaDe+lqjI79eem9KgLJg2o9vXJvcDY6rtRP1APd
Q5hhVrsslO5WeFjnnunL3IrhkLr3QiDsUoN0G/QOoH/RvbndYNORGO+kTT2vEA5t8DLJX6Ro+Foz
fdd2SYau5yrUScsYoM/ABqgD7VvrXwIPHAzAxlaX0JNEr4xro/30i1u2eq9bXi0KzQDqnlCdvOy+
Dy3iLsmASHngC+C2liS01dkelAzeuxsVL0cbO1R4M8mZ2n2eEtrG4zQkEpDJ1XtEwUu51U/XrEJ7
+C5usbKaK9eKj2pnzkyyFH4a8xABcJzSHj3YMDzdPhoIuYv0nQWQC+u2RX2gopfZZPeUDY33Xo56
JJ/uNXwVAlQFic0P170P0cHLY7YM2qgxHq+hXsfI9L3uzNTEGTOMSPZy+SFTMs5cf+4q5Z2iAovt
/svj/nJOY41H8PWD2vfJZdOp+ClQ49V5s6KAHsrv0RuqB4EJ3Gjo0iQU6lpFscl4ees6VXaDazr3
+AUIGdp8cc/GTtorWw+VpvSBLsVBCZn+by1UMQghkvfEFczxY/MM0oaesSLmVwmZOghxAob1IQK2
EtCejkfjsz8KhwUyttXpTBJFUKL0aTd+Pu+nGNrHZNLzBqONf09sTWQXr0eoYsUbNykEQcvg+RDU
BMkXmka9XL7BkSAEjciPeV00US6I0zy4M1OWqHvaiuc2kdPw7w2oZSiQNtVkNyi2pRh2kOD+VseJ
itz/2rpY34vNqN1XK6oawVx9KibnbvMIETUnPN7njNcYMnW40glfXuKd6M2l5+gFhxWDXkbs+24C
3q+POjy8cNFWQcoLNJMpQV7SFk/PDOyVZRCBXVP3gSFSkgM17jVPr2L/UkOTEYgjOAOE2ki2d1SF
Bw+/K99WIQGWCc5vSHvsiDCZTNJAFAOs4H2yMqeK8SJJoyaJC6enICoLVrACAub4CYgadORq1zAv
ZQQ1RVlzhb/IghQ9LAHcWGykDxUPC8oFbE1/KuYx/LTlXwvVp+FaypCZzMzYp+rfDfi8OquGCrwi
f8lLaX1i4EsFAln7je9V/IPlf/rVQO+r0K0RG8+r1KkLnKNMQ5wp3Gh7fvdk4dixE2NTqgtarpzL
zOFZb5DZhEt2SwnbWfBBIxoV+O1763/maayUn/n7TTSULQYJ2oL2B6K9V0OR1T+2FhqScUTGczeo
ND4rrboU5aPoE7nLk5OEpNTBrybX8/sxjQnJrpLToz+wWcbFVTyAeMqiWINu5Vxn8noEa6SHBT74
SLW5kN8PV4UmoFtGOSTxEje5oD88hHOYZa/2K33+pUpWbV7MlGUUK+kiFGN5vctA7dbSJxuZnHhp
g4hBAQdevWxv2HBL0jwpf46ykXQpSvtTxHs3bOD2zuiM/91XIfOY0G0cgvODGnRngTZ8D6cKy7Q5
X3Um7D4c9HSSGFcaUCyph7/+y8gxjhsbsYh154CvH7BVlvMeu+BdyrV8dEFk8zQjf6p5dEzvE9GF
EDse/CXBxChT/M4TCONqo5bJnxokAtC0A3dpKTnv2H6nXoGj/Xk16qsownDimOX6N+DZF/jGY2Pg
iPSW8vf0H1YyCuNfD53ydB9zfs1likzVdGRDKqWZCiFaYg3phdtTpQPz+rHbqvp5fufiOcKDTb23
RAA9ONnyShfbP0yCSINEpiDs+AGrke0Y5tis+STBMpyot2MZZkDstrEw/Xy3Gku5xFifaE7N0vVY
buzv9JPLwPkzlv9ZractFglvsJyKEQS02JBXrzEMfnVOfMkoATxkDwZHjV2Fd8Xsecf+t6mnTe9E
eVYxmEpjNhnflPwiaozJjyZ//o+7Ys7OBIpyB0JNbJVbj07kx8pM/SM0MWH++/QpaX0AJFp/VgMQ
QVEl6fPamG7x3LcGhUqrd98iFDUYS7Y+GMtT5oadSn5aPpiAt8c9Vlnj8hLJQZzo2GMIc0GU6RV6
i8nvf0TSxb+4iGAXG9u8Fo5ezwGawpCXCqoLEbtFZqwvUdgvyCDqRvAZV9oSdAuL0bAKkrvO0nts
Wniq5Oc1gGBKxnmPlUcPnx8s3rE3cjUtDMSwlFJV56DUB/JrS1cwnzGiMaNW/fFoH7JMXGvlH8an
oisIORwYmZZblrqxyE3P69hTRQNUHFkiNOPDCsNwJEE4mhEVnynBYDV2HUeSE0/vgqYOC4KK/tCl
wyqOBEdVVEmfTO3uCr9vCpfL87d6N95k+WIqBmTFBRRKLMLABtBiCvQgWFAxXhP7vYcgSCHqHbl/
tQ310rVbw614ETU1ZJmG3S1rcqeYfoMKYHOz5XHpWm4RBCOeWH3I6Ov9z7aZM0bCRh3a+MoZFW2i
wk1arprRzOmGL29avHm1Bb3UT/PSqOIYAgkoNj2kcpPkvAeVaQrRe0NON13jTKJ7Ohjkv4NMJWhc
eRLp/XiOGtI+3+eqsO/sYb1KDItQi62Yt2pnYBbYndDP4CY1J5Fd2NZon/wEg/hSdriRk0RXpJli
tkSx2rK/7lO+MalSNnNdIvoeMyaoKT0r3hAlVBiM2Hobdx5yzz5+FOmatrqOQoVb7jjLD5Mish7U
yEU4TPfWip4PdOaGZygx+b3+/QbupSL9YAR4O0AuJUjwxyeyHH3EjlMjH0vz69mnSA9PCxjSglX0
h9Jv6wFIk8Qgwdun8Sk6SAG9pBTlBSQ90+7ZU7UEFCxTiUSwwUF8+1wqjV3FOWaTv43+NOBjPyd6
m0UkyUd3Cvz/D/fXXTijc2PMTMKzWxGA997TMoQ4kCVUgF3ibGxzEnvnVSgQHPs3Q+ubF2SnsO4W
taj5dXq/FVZbst2DZnWwhZcvKhQnHpw8SwYPmwv+4jcDK35yBojgBwvQYA11mycRJDnd4MThIKUo
/3LWXrX0WTr0k0pBWeGRmZwIRREhw4PLVBla5n447gd0uvh/814FuiDnLDSXBVKAyrK+fPNh9JKE
7jQRZmKOgrSliRFpuhzXQ/BW72Bi58+Poxe6f5XU6cMSIypJHfn88Q6LTqSjwSr7jZ9VCz+YqZPD
gLzO+kfr0gsFp/5D1i0yhs8DOrDesOVAzUayzf5hcfG80t77w+oCLulNcZTaJKQJGYmL7v0mC+2g
L5BaU1HM7WUFTyOsCSo8hWA/JrjRraAd7eAg+6tDeZ7KeRlA8wFnnH0uAAKo5Ru7ayMhpw59PKmY
pkArx0W7j9B+K+sK8vnI1ZaVdEvluEvjoS721+jwmueHKW+vXRWNrTN5xQVEPgiP+/h38vXbWC2C
HgPpJe4nf/tVBpJ5qGVpsHBhIi6a7c2l0LOW8eGqxAJkiZmkxmAhsbjZd2wNt+8MNmXDYn72Hy8n
9zNQfAApYlASH0JGoVWmzrFsFTgPzv/47zM3Oc9U0aAJZI+VUthRKeLkMS6DKD6CLuE7EL3a6zeD
HggCOBk82iBmDLTHPxX74wwSZ+49uGyYXZrdEffkvjvtS4ZfFlUrjV/a9LlWk5A16/th4e/ubGDe
67qOpFg6dfJRuj6Rdy9eedVxBSwbOdui1Jte/bGd5UX47KaAp+lGjSucU/k4hQHIucfRgZjllSUn
sWisZKtU+ptpvu1YrOL48X/eq3y2yMkiZQSViljQn8Mzhhk0bh4ADOpdkXQN5r+97I/iEh7lYrnT
aZVD9KRHUzwbchrXwbMVFEqtUa4yHb5ZEoX8GIzqXo70Met6XaAePXwAR9sZOVoqzLEKq0CYLfap
yO6Q1d03O+DqE+Pdz8n2A8rVrxppNYG4MAHDzOzLoDqU0iv+qMMxZKQ8hKXQO3IfzzakWYVMXK5Q
Wtr7px5aAo1CkfjyBgK/NXeg0pImqVgG6AHhTjuSON+/PJf5V0G9J/LxrMWduMfdFYQtp27SH4Zc
QPZvq/GJa81DpTXabWq5W2hgYAv51eTZXPN4zhxF7rNHuFFtFPTrGHwEXe/J62ZFEwBeySdr1KAi
p8dUwb9bD4L3w5/e0Pdx7/d5HRsdMwlusq9XTlgIuelcYVbO4sD46UwF341ghJWsHJIF2gpHW3mV
R602A9I1TTkYaE8z9TK2q3dsoyFzBo8OYudQNMd22R5SYmqxV46X/NTIMtWhNEC4hYTBVX+NHppY
/vxCDGwKUYOUEkHA0kzRXyZlmu9/4gjLCDeYMaU+YvoZZxPKLcoM2Il6ubJIqFsIxkaltvK/lyJX
TxhjLEfrvzWkswFSNhUG+wwp5njL5P0yOnk38kaVeL0F0HJAjqU1/mr1vusHBo79akLTPyHwm1H9
Cr867E/L9HYKkUs8m68zLr7Xed8Le4vdKhaVJLFjWWFufy3LE8MXEaoA8j621Byj6PSZS11Ztdgh
A+dy/5+crnmHKFm6IyXkFmkZmV0RR5i89sJGpnpMzl7nWk8oOUEqCOFmGLSCW5Sbc+PTtDs3sEwF
GpzpD8KzokckTsfbEY4zIEUZ6rl9qDbxh50XixxyEhUdjd4uap2XVd1s76IFmjBgelFMV2xL1ZLR
FrF3LPrIVLKLA+QHvjfrSOnnJfx0BnVSdw+7jTiJNXKSU3nigjf0hlxekda70coZiFojl0YLOD/y
Z28nxI3y2UF3Ge/LokvuN1ZlVNXNwsyH7FjMMMfKfGm8pRSclBC01U7O/C4MDkU2BoWQ8GsSCNPB
/s6kZ1/gJGDdWT5q0vWDxOEONFtvoYdioZBNKrdHLyKVHRyg3RxkrTiTEPXZTwbrKb+kkcywa6pB
EMlL/iK7KoK1/2dOQgfm9nezz087wbc1caJQDKUb8zhP07pSG7zkE4Rg24d5Y+jw2YXDIeJuY2sP
+CAJm3v1jYBxnhB72GV9wzhg4yfBCzMwWck2JZWjSlFVKGmsVNUGxlMVb3SSkKLV+M9x35txY8He
uY/+YZtS2gV5fUO8mVG4/QJpJh66WOlnlg6MPySMsFt5j5mmG9E1ioj3rS9WUcrQEu2seb+0+K7t
ru7CxuklMmCqbEZKCU2FnADu1IyT3vcvdn6E4Ixm0GER9FxX5OiCR6y4yxQHYBTd2tonhVS36Pri
NW+vgAF+J4kJGoXyFwP2zYCMS1BMlNhc5bKMCr8PgmoAp6uMdVNYHOvo1mu5vADDySgQksqcD0Zv
vRoeteLG8cdYH1I7JWsLsFGV/68RbFpwWtnx23ZNUfuHUaVh01deV4oNhfQVbar5cOy+eDt3eY1c
+Dcp9kQU55Lf7tjUBehMkw7yQE+P3q/AGBoNLXBK9bA5TZ0YpOt0e+LVuqeD3yF91XZRBA9nujCH
90Q52CFMImUKqxlkMXheJ84mKFKp5cQP0clQ+kddX7n/pUJzmtoKhkLxehbsovqjFPA8T4okp0cY
YaD3s5wt0RstAQeCwuwVc7iCqZhzeHpcOO7W3sepxOdGD/b82OFFdEPy+LH8Ag6CyAq42S2YM7V6
hzFYYm/eXSPM/JAxi4mccKG57DH22JOJRDZIAparAuA76j2XYzv1w9qClazsyh+gxEAe/dlFpSCr
ikOVg8t9qAvsoDqjlhRxRiMDQOZ5FGwhsYFSdmZrU7bhfpWoW0ADlLUBzKg5liIsn0AiP89Ykj02
wZHY1xoqhDBEBHU9go7QTfKZCZXN9IQeo0LjstG+xHpZ3XLTS4/p7yo1wo+gwXO/6BKS3jnh35AD
yN54V05fegzDkO2l50Ya447k+DJYJz1nU4Nv7vwmi4AkQmAGu4mGyQeb7pLdi1QOr/ytCpX128Gj
x8bAL4t/FQF1OeFFCqlQJebLvKvL7oUiCV36pQyJjXxDY10VY7T3wPDSak6zZSrDt2JoCDSaVEK3
mj4GzGVHajBlmneimDLhJrioCG5ItIPULJ85jROP5SksrqEB13hiORaP2HdpbYl+mzkFWt/ohpxx
J07WIbyqeVZJx84VTkncZAk8iFQN34lxAkomKe1Uj/PL/gxX8WJZ8xMYUTrLrZnH7+6juPZWqLas
NsLizxag6cUOlzNT1IyGps6phF9Aut7YkVB/qYu6K5SyL0Vvu93p890XBMp1SUBT01GwFSv9GMV1
+DY8kDF/ZVYhhQ3p5x1yRSeVwMtuDfDGVgk7CLKalX692iOYtGTWrTUmrqdGm/QPuyGSuxWgqzJx
nbkwN+BH33Jt3JEMGUdrPmi+G5f850qCtCGLMVQme60r8mIpdxFHQ7+kdwXCusqTTf30Im5lOe+r
vzWTogZWEzvAnaE6NirK0jYwkJgM2b4LKVGa2VwxHbKwAB1t3MiRtRmm0UebQbfX77myVZTMai0i
/R6BeWSfU6fPHJy/So9yWaszBQJRX0N9TE5/zwqyMM18koxiWmcMbtBnuvutZ23z27bB+fF6xhlB
BtQowU+8iqenuUNA+d6pXaEZemMxRjT4ZZtjblRebG2KwW9VNrjEscDnMAQZ4OpN/zk+xLtc3wpK
whmyEYlWJf3gzc5YtpPWm5Srdf8RIxveyt3YLQmoWtEecaiftPBBA5ubDnzWDgGI94tVfoDt3+wJ
hZuslgMwPIVRBcJHJWMI8uzJXhPRiigxOBQcWbN+6dpRMA6Dxh7AumDuYcvC0pro1exdyKDfZMZ2
pq0J4HtJn1OpuYYhxdwvNMXPCZkMiYGAxwhXdC9ogDXXuXYJ7tkyGG2+ZrztwWmus2gfQryGneK0
MItSNuS8l58Ez3ZDq3LDbhw2sl3+xz859dee8QZU146ZzGn/dY+q7A4UjRk/B5KCFFvBhXAVnzAH
y9brx9++tzGYt2c01NCKCZ/erpRXbpzKyybxQp7sxC76zrlLml9C5I2oUB0wQ1Ny/JclRpfZRqb/
qDSZzQXn4t6nlhc4S2kF7ZYCHcjkcsrWA+0NbddDo9CMtUwgpdVBtKAPwcKII9UI906R9C/gFFZq
U79RFt1/copP//0/D8fCKMIJMKU9N3uYWEZJufjueb4SgvL+QKViA/qdHfNEpupU1aGBQVngqgVr
TZy90klHxMWlOXuGIUTVV5nR3t10NS1v+balR2qLKA2jVaCneoNVdcpJNW9c9nWGtSUJhN54hYG9
hLV16esZ77kOwTS1LDxQq+BBrPtIkF6wECIL0lstNBIPcpNaL9oy9J1IIla//KAKShfvi68enUiF
k1caMeM4euytCFCi3XrE2SS7g443Ty3WqUC5BLlccGeBGlofrA1ClHxa11JL81knnBr7k+o0oBAM
sLscn7oNaERM8JZcBfWCwEJQjVDkcA9T7t6fLuvxmA1beR5m4x4H+0O7K/KzYzX6B7umQmo8IjSu
X9rh+DvKGolshHv5qnrIBAutovf9rNu7vZ9nCvEyfetsYSu096Zas6LeKKWIzjggBsiouszOfzJ0
GhqNKATd1X5DBMKdFelLH8c+k2WV3pN//nmuM4jkzcdCI/mj9KSlqBFtRCgrvzNHnw68bIAzNMs2
vXHVXAuzMncqsKt8IFd4P6aYvQoaEkl6PwPrEqq8uQ5kQP83E6hqZMOKIcEi4RWczAFTkncRPZxo
rbPsW59MIholrsUAhN47mk0HPEpwKLHFpR/J5DJXUeS9HH+MFY9KTQH+9JKfoB4xO47GN9A07DtA
5BAPu2A7b1KTA9p3tvbXSjb9BcOaR/06GEzv4FY9Xn9FrWIblAxYCHQnHZhoUleR2n0UymHjuXEm
AU651plKwgcJdcXJ7Z1Nui+O6ulSQ2pBswQNft7xlrVNV/oeK0+H/vsjc/aSNbmVmqD4RkofCM8k
pILr8fN/+KrN5XSvNdLrhA2RLdfn+k9mEq/h8yxlIBGABpF7P7uceOKQ+cOpkybqqCS9BI4MhTHA
CPRi+515Rb5bXlXHyR2/++3OHezPNBq3uRQ3c9PgFg9+IQDfYwrKMcxIOhvLUJzcugUbj77X112l
3y6njbgiI76Fg7dS+4qullaCsbLN7nm89kumpSDdrnujCa2sTAsVyZwZbMp3YciNpzgjNtl5Z6F4
QzqtNa9kOc1+OlIcN/j4+r6zqeVQsMCYrm5dUjLEQfDEzFVX0IuUWcPtWAZHNELiYMJnRuxgporp
rONc5t3RCoeat+GFP01jfs8d5l7a/K/9D5JIYjdA3N811yRGJmOTl3j/vOaKp+kTsOkvdlJj6qXU
kOspUoCUKJ/gtqBkUKh0wyCqpRjePT4WKeVzRuh9ihVAYfXhnq9sioUHJw1IdQWB1KsAOh776FfM
mpT4Q44qFg/I28Tk9oN8R/OYvv0BSEEeCcpM5601nwPEBYBLzsQ5cQVvw2v9Xu9UVP/4cwt7t4ae
ixVjMwLjCsIOCaraVKVmuTS95YUp4oym2So07i43oNlMzTtNCoD49dp+3eLRWnH2KBAUP3HUtW81
mEdQSzsLhuDacF2fLp3Usu+8E5MIoXIFK8VRa+hRq3gjMe4bhYR3IziI6891PoDDc0dOvuK/sFCm
OKR+xJeiYarKNJMO5HZWU28qGbPbia06SBRWa1Lc5/1q5q0B1TbroaubQQ1B5ajSgJWtZLKtqlxI
v7fDVbF5YnewEfXdp6PgTCErmDNi6vK6KQQhS6XwJF1pWqvoUnBJxsZSy3bJXIEBhiKZ7zFfjiRS
PcwIZ1/cZVYn08bf4xKCb/yIN/otfHXNSip1n6e6ObEa1DGtdzxrYzLTU7c9RRFqG9ITWKsJeWB/
k5KiEG3KqICFjdO9Gd6itxGCLuUGzeTPs3+qvjKM02OSJKlTlfrxjvIb6fLYlZNgXOvtA9xGvQi3
4YWkobvnvKQzwlPGF3SyUtOSNsnNoA/Rre8RCniI6Y78pYiGNJ5yuyUP8jLJSbgC5zCw1cmk42Rw
NFpeNTWvz01FbLZWm+UEFBREVUXCeajRu4mjXS5l/l7hd7U4SHDg9QRdMft7EYCAAl3gnJtBWwU2
hoOQUww2E5n5OxMpFeg+nVxZT9lc6F+0TyNVmBYENe9vIizWpm6Gmk5WtJgxeXe3QXxQpZYIOFX9
JXwwhqO0wrVzNPbgu6REqwoANAIQ26T/es+K7W1X3aUgga9t+I+dfYbejpmp3tDD7RYmk7u33jKz
o7XNtReqtmrigLFImKAPe4hu1MmAazEYGNQxSoEmwYQn8k7OI6QzhHxh+QD4Ve+qO3A8wLl0q6Lc
P8/aUZ6r/l4fu5HxuWOtVQGXoWCUl88VPl4wotSl94wysI6/VgY1o4Bfsz65s4rLH3/InjqBY+Cz
zSTu9tkXN70YTw28xvMt8n7GvCHd0KIoL5mSh0NReXa5IDJcj5FNI3FGIMdx14TJq2S08cg/Whli
T2acdqCdDluejyQDRua7otldWvXXxkC//sgrRDSvGRSMzQTnJfrxOPFocGLg1v64mWVKoTG7gnYp
k+m8EWGAfzO3Lvh4ahq7jTR6ajQ02ZNzn2cXo3vrjXbAyqtbKs437TSTCg1MICbzXeKrjwkwjKTn
CuieviBuc/tCaqIpXrDxcdkVkTaLcX3R6zOMfvpUN6LfQl/LQIXasr7HOqP4mKDPPB1DHMMzESGK
n/fDS8beaxJX51JFNPkLtjeS5oZ2eJ0Z/7K5EWLPA23QGJybIeqebXgwROybi5rb5O7IKV/mBGWR
fq/O8lgMYZ5MEmst9K61cAs9atXt/i7OWYAugf6kPD96IB+9z6m985TMWOGIOkPoqMYRbxeUtNWE
0UfEFuihnYOSvgzYJeE2hYf4qfhRZKK+jae0ys3L0lq15RJEx3nPInZnvO1uGpgy9cq9FkHFT2L1
sRAss4nhxe0MLVqYo6hiin8opYvJLaqEpr3yTxWT94/jAqYdW5Q4W0WK7P3w2us7gYgh/TUYdiKC
rzrgdm7PRTV5wH8pc1aoghLyemZwuPdF9MOw0KlJs8qY9CFBVesKagoOS9voSXjcNuUYx9ORXH/W
DTBUXyTr46Bg5R+DQmT7z7fn7rFQhjSPwDZBB4XW+859RVZE1j8lrGWmpPvutM5ypsUYG/XNz1YD
feHG1bynL0aqTkxtlu5iv+XWLwp5VA1+DIWlMnU7J21MuQr8J2ptMgHpe/Wu9tWQzUvB/MvPCyTB
KmQpARRLwRmr/nSIqcjXC9DFy7/MWFc84cvGBeYQV921XtjfELdG0V5sEyfDHzsy2tzwVENYze6O
/RP5XQ3kH8t9GBvKys8nbEF1EtZpx2A4z+/eYTnNtrHztlnjh+Bpl0ej1K7V3ePxO4p/odg7JltS
iNkdR0GDs4wmfTINU5FqXlxOSRK8mszIsj99BqadoTVy5NTRBfYFDE0NfHZxGA31ExaXhsOhfuo8
YpdVQRc560C5/1LtFhT6Rqu0lQyJ0SnGH3HkSGAXZzivSR8iyz7oX178IY57/CPRdW2W3p9uT5Tt
ATe+n63pojjzZ5pAsB5d7xrrEnKas0QzY1bJwItQTyqdYi272bfSTTmx+IN4WB5QdWNSvL9pJpEE
ad52TZmoWh0OFUTSsfGjdFrQ6Ng+trudGx2DY5LOtNZ+90fHIrBwVzeZPwS/jwv2XnTChCwJn/iB
oKVIPnVPepiDZ3gILlqEhjyaCUhbA5LDtqom3jzfrDttclUcrW2rNuyUhsUCCA74HKj0oMsQdL4i
tAQcSE1eR6wFDGJlnO7duhmb2LqCj/v8hFoWkWvvhRamy9jqyr7nDuIJT695E6EIAd1p8vauqLVk
5xojJnK1eRPHoJEsFZJZjo0cbzrZPriQLbEMLw94cWNt0kqmDZ1sbAg6ZWs+2Xkb9+rfNwAhGHnG
xzGp7kEltVmaLdunIKo0COm33ZClYNERtKsebwCpz4/q3kGdKIgsUXi3jXewQdiVagpcnkm2jUPp
S/ibtK4ZKbigF76eOnSmrMfH8k3f9cLgX9gzzxDPGm/Q323nf2oE/aNgoHlAg9iVlPNrJa03wWiJ
SbdbVjNayR1Dy3V20duwDAM/bGfKYwnXs6IhGocia17T1VOyvXgdEYXLGlOv3U7K8FFjU/JO4HDI
CgT5TAuR9o9Ohv0GH6x4Oye3siZ2ryfy72/H6sdFTjgkEFYVDNNdsEvz/nlBMDAoLps7AjxqT3Lc
P5EtEHW2n4b0Z25yLHSZZ1L6dqBfKVXg/H8Ui4fvNYXzRUE26FpeeV5kB+zw1EwDLkZJpVGI3zIR
9sUGDYoZurDhJXdNV8H2CpmIV6jjugkyCD7JaURccJnNGJ4pw1KAypxYGFz+S2HTS/0oj5jfkBR6
7vpBsig2B9wioBeaHAAwJN4RF5l15jx1SOk1HCnghAg3sNUwC+rvQRUYkCc6Qfm/BmS5XyYEDIWb
Z97s9yCA9IrHeVu+Z7IgA7iJnSbZsZgQ85uwrCxpIJGntWtc3cBEb3nph3iuo7n24UWOXbtkcLn5
muKY3a9FWlGgL2dY0jOzC7jx9qPs2rVLYOu5NHz6WE3yQywyAF6uHGZALO9SSceQAKv+GLOkKknJ
+6DMg6sReERFkbR4Ya5kbbOnUBBFW2v+2yxdXVE3murR1SqW/5l5aLHXd17nz8sFh2gES40NwCsT
W41FFaRryyvj7UCTVwKJYu8yypojSReb46GEBahTFV7ehQ5WHqUQMaqOGO50K/m2MQHF4BIyfRGx
lfJoiVXISlQCTtwW91oOTJg0u5fVQWRDgUe7xGunR8RxSEIWKCLE2+vX8sN7ODkMVgXCZoZrA7Oe
HCTO4LExP1c6k8JTHypmgSknmx1ppc9Bkiix2CTS1m2EccIDlJmnyXYp2FGzz/w0DDiqP6bDXSdf
pSnHuLkVnRfLo/r19b01RLWvXgY/17MFbfG7VyPWUbS9WTAm/6g8Z/QvlG3Wvx0RVEPgDetS75PS
ZU0azXkoitRa4uCcE7H15NNdgUMf0fXrOR/MpWa3aRWbUxxh8mK7efWU54yQYVldJ+3dv8BiaRPG
spKWN/6Rm7q6rGu/DlBSWdl9nxXi1xyVtAOMWd3U5lGt5xQl8tjtkARr3kHOUiHNaJp/4K6TIz4f
aS41djuI6hGgunOb4/XunPYYi1Ui6rmCnPbm0x85TGFnTM5z2t7R+iB9+m3RZKgkhAP0RHjw4RrV
3Oyzh1kgx6qS48zpfrVJunOYPjjeJQ+6e3aXZzFuwspkGf5mPZvg4GnX3XFDiGl20B75VMhwxERG
sUOwHjs8JKZmK5sHkchalDqeXUihDGtcV2JwDuii8AZ3TLFD3qlZ5fiad9A+GOHulC9nHdzFrhhT
QqEXXAfsjV9d0z2BM+TWRXMPH263dwAOlloIE17YmGw8RwiKRZO8Jo3XoiKoTsKG9RVKIVCre4NS
PXRI3aKeiIF+3VzUXV9cQuP1B5INUVitF6AQKUwGWBvyTkyw3X2CK8BXz3mcBBfYNssplteEPaH3
Y8MxgG7CKcphVGOcr/wbnICba7lzbeOe1+HWC0slB5vLRQKGLJVkUfs2EfuXdyRKYVSOGB2xcFEU
ja5kYnv7RsWxri0WQVGeBo5wCfdC3lejcSXZ6hCnIjqIOY2wVFRpDQ8TfZm+d0o0FS8CQpxF88Rz
PDY89A3M55l/O9/eOdulKNhP7X00lJlgAM6z4C0BiIKEJHOVadTYdS7YarFinN6zuXuTkiM3M+lj
2KhSPs83ANK6UJt59Zb1KMMOtW9cwD+FvjExKci42DwbcnelYCB+2r9hfWTdIOISrVZD0Ei/33ew
g/qczNrZDZzC/soNUe2O7ZVZMWPrbyGXnSfoidzRP3+lyP7rIW5lGBORvcl9KdLCM8QHQbS91beu
+8QrWDEwsDYMXb6zhHNPurcvHkk8D2GZgdVEr9Cth7vhhfvzQt/75rTgVNSMmuhbkvvulcZGKb7V
/6fEJY2FT2AqIqn4Ki2uAn1gEsjeeYji3bXwhAMlb6/rQgdCkClaHSqAN+kD1XzJmbZ1BTNivHlp
CEbN9WFnbt8/hS/qYudbLZa+QCw6Tg2YC/iJe4CdjpGI+d/lkw4fvAkW58gwPakwHXy+twrZvr8J
9VuqfJOxWbhRKF3W7r9Roy/XSSVmtCsUWUKY0A/lfR9bZwPRTtE3ytoiU2NTli6PKHn5ThwsgLfK
HMU63zaS6g7K96fUT9Ij/dJGj/t0vSWOkaJLC/V5/ScR06KFP38vVyM8zelSYS3/NLLNOXsRwlKX
lXvOlwlfFAnqAl75R1y/JzsAmWhW0kVqx7BOmUdwEEK2KwoNVDF/R+BE8DyY2MU7NSUyk6nkxnOA
okEmPJV/m6rzpXUu8/zs/r4309jyPykIznuZuo8OamdOx/psMs0FTxOBxZ401OrxC9fVaJjS7tEK
19vgJ16XNO0QCwt9u4EEVuC+ERMouATwDnJ2rOFVFw8s9bsVUBafn0+mVPyrm8udLcMuNdCqMnET
qTSPBKk28pfR6SS035grcu6VxZTYTbbs8D+rASUTptsZ3DRDjRYahuZx6cLcdLrQPAAxbvyS0ceC
0AR9qSNioQF00f5rMtOlX7UbqEv33AECDQjpxA0rYWSIff6ZT/dTtaw+8khEVDrEkLykcGT0dQ0C
kLJqK6YsWrfw42JFdR9rrb1iZk7MptOQmGUYiLQmiVDK2jZUK99Lm6vFv9LnZHFr0eYpb5EckDmd
JGzdlNw4/u76vi4Oip7xiRTMvVDJJSCQV0utaf23QvNeMp1/bY1EK5OMl9n4jxWEu9352sQ6Dqox
ZJzVXpMb7k4I8A8eQhTfaW7cxf28uepsKaknHkE1JjDUvZKIdd4PtPohmt6wqFYS/NwuQ+dldJyM
unhxz+dMqVeUsnDwqsBC8X3xVrVrx1SQIF5+Zc2G8us+Duqmo6fFpFEXlnXoF2Bu/xeTLvdLf1Jw
2NPyqTTzYQA/dFzZKEmcJRL9LDOk+GZ+Yufgf3KPjec383p7IgbEjuh0OyK7IWS0hsvqaUFXsbPm
m1UoIO/vtw8Ool712pyGfQ/CVbWfs6Hb2lmIHtyHut2HHUw7tUraDnZLul5DlcgnDTx1pESVr260
/kFICyw+QAA+7z1GkpqWf2RdxCYRXKeNKjA/MHMJEJuPzRN4tPNw6A6jRS1+4iVUJpgsxrz+2d0v
PRvp0zfX5AL+fnPOWU7IC7/LtURQJcZJy3Ly3heTPTskcGnFl6KHkR/lYeM8+Kn6rSHX0rOBfPZ9
YTSrosSKuIn+h7aMP7P4lfqpAzVGScgmbBEjK5rzIU79bcDyZE0X2meP+1V8kxnPHNwbf3Fw7mul
QtKJb+h6UZ1PFbIdixevVxHqG4plCdBGZ3krcXfuZORTL4E9iYMbX9oVHbZqIui3c+tdSedlJIKR
iw25ij3WF13ehrkmAvu920wq1CdEhEWtfk02B7LPSOSPC700yEsTnsu3Idl0Q//Yk95b/9f9xVXQ
OD262OsbLcZL73SyA+Db4mMf/Ne+ay9IjJ2WoInMZlfa/qD1Ip9iTR9MXT7QmBCodADVDpDfHPAP
QkVtmPI3ctdaXspzTqPQa3NHf7iQ75H8XK4k7ZFRf3J3GD2TsElu6P7fz0QAqhpXOJ4g57WWTaO2
DzCNM9Dv8ckS/LLYQ4TGXcpE4lJhO3oQW/WtmSnQqxCfU4N20e5bRYrlIE1v0C6V01sG3yX3iDK7
oJ0VmnQv7rFa+qSo7JmvKFWrnyyKdBLMq35GrXkRaBO2iGveWQ4VHdkimUI4PZi0GJVcW32T44t9
ZjzzXzVkAIYkyOj+tstyUdCZuUwgXQmzh6Mtl/aPfZqQp8IuE4dmpKvc/xZ8fngUvM4/0RFchK9E
30laSTpCCm8IKUshlImutub03eDFi2fZDUornYOqFeglmRd7gJgk9C7YG2u3aqvd2/TbZd2oKe57
kgQJghBhoFxcSu5hdJrpreme4Mhnlqen1HcSfew1bqi2EQnEZlHib26b6vCQj/vA4rppH+dLYWuX
GTe0w5OWr5HrqN3M+3+kBhUuTB8KA2vRv69gVoAnbYBGC1jmxthfkvmaVqsVxJrnUBq43pBCf5j0
ZBFw6pGE9uTlxGQB6o9D7pgzJneJhTRYnEikB/juEQW0LY5SLRHXk7i6TeOaxSQvJ9ap2TUIZWQJ
ENWIXcwSRATrVF/pqVr0Jn67X7/1LzopjyOfyFbHSL3Ne860eL7DZsDZFVo7PSONzCeVxYZPIYyH
dD7nKovHD7gK35opKcanstiPy1Nv8qHoYW17eU6aqNUHraRSSrDTX66mK5aN0Ym4AG7gkjxj4Llr
Kn/paR+CuyJMsT0KZm1EY7T9C+rCm1Bo6/+VFVZAC4sYHYdJLkc/Tj0mtZ17vTRFQS0FHmxxka+B
Zqnsl2TLFiHXHGJGSxvdv8+HZ1CJYMImkZczeWZvDH7AtkG2Dm1FnogQM0njTGSkn2XodVGa28cb
NenrqmpN8MGUW1Jk+JA/UEG8dthh8a6RK3kN3gzLHcay0cKq8Aoc26VztDO7fowmdJWYXgzmwj1E
7UPt+c/uYq9tnRQCSEdGG0ruQf6ZC2sJ5L+SnGvPl6iGGZBTRpFqca8EeNZ5yrfuLaVuG6M/gWJW
B7mydh0Dxsa4MqsV9/IxjDuvxNU6UWDhsnIMix/YniLdowhJPNmPYJ5/fuMjSnt8mAmO6rs9xKdn
CkpJJ+ZroL5Hk99K3EcqeLCXA99IBtUhwtBH1Dg0nw0+A7HCaN1k8BRsZjvid5hroL4j3DgDVUbK
bSjnS96ScgKJZSMJ+uPwQ5abW643VuLx4BSUG4HF36/rfBtnnrkYXf0yE8z9LTdcBi6jhHx6YI+m
F/b1u8e8tcEEf1xNKJT3j/LZE1OlqbZwzULiH598VPlhCAcW1YSPBfc19aQHamnNFP41xXR37nbo
oIANuIe1vIo2Jr5kuiB+KNwibaIv206ip0cQbqI/n8vqPIva/l7GeccaU8nm1Wi8C9UFZLB+cXxW
OXmoM4Kr5z0XS4kWp6hg48EZtn7qEvAncD5CsUGiaE01wJts8sAhwEuHmhjDP5qy5TmaTskYt8oe
RgBPpswZvSZBIkA8j9Cp5tQcRi6y0pdTeufhdISrHX7Fryhs1VnZyGRXmzspNtt3AarTHPQQMf3u
XktcZcrT3HuQB3sZdr+EY6huL/gEEg9CiL/zP9F9KpPAMdHU/WxfTcVFQU+HtZtLgAef2So+ZVml
HXUaUfsEJ9/Bu2j4KgWV70rZUg6+ct2RfwvTgS6AtKaxo0315tg6oS5XIeZu9daeAHOtdmgba56K
qKmpdExw0fD4/zFgBsHGKhJc4/rQ/cjy2VyQaMb1ITdN2yY9panVAAPF1WrY7kaWp3K0g5IYZl3/
sMpdvafXGeqNIkQVeMz6V9l4UFw+7vhlKRnmc/2wU4hMAnjItJxO5ql4U+vpORyG9R5IMoIz2VkW
ocHmTOAZs4H8PdPbpseIUosmdsdpAd6qn9mCAKbn2bETZlAn3x2D/0W/P2Kv+13lZ/K2QjEv+5rc
oqxrXt41vqXb6dbgVqoDyZFEVH/9D3FbhPWb1RAxfRpZTM/X+yUPEGcK8oIt0s29meHFIVWuGiqB
rnwpCGQqkrtmbML6uGhmg2qMs0hZ8MZFFmN4uSoQQHEEXYCWIrIxNZZ4r9ZR7mq8vbQllKNCgjPl
bHT9FjUFtTOxrTQtIKnIrouIdQkDJ67c9I5LxsGQW92CqHLRrefgSCPH/QUFnmjqF2kZV+yDMqUm
4Jh7sJLtVJZc10gRFYC7wbEN+aTbTTyqBop59NRoGL0xJ3+EgC4Y4RXuF3wTpxJu2KtqGDuDHIDi
fP3swt5qGhcLHitD/nU+9zpMAqKJ6535vlk/52omSBNjWOCtLlO19n1svBTfxrtlBbopisBaJQz1
MY/84X62gn8lVSqGMgCZGihCIHPXacDPEZhp4JOfpmDiCSY8xnHI0KYIzRL26o2tPe/hjbkJs5OK
mjUdVX1Yyn+52Ejqj1G1IdTmq91N2DwJA3gltthjZXmd7AmpGp1dfaO9AZ1of7aN2nFiu6ippw2Z
wD/k3cOSNdmRHU5gy/iXsIyBZJqnDIMp7t7VEqHOu+po2CLGyvaQoIJuILLWuZXodiQvkl4wYGoC
OH7bM2AaVta0Vh+YfTZwT/tgycA71adgyvTv+oIzxfj93LUsUzglcBP70pMv+rClDFwP7hgMBp6s
bpD9pezu26k3DSFBH5liFIFe7DcMqiHmiORMFwiClWbMtendSUi5MoOTrJmSRY00N8XVwimbO+s6
fGSitWDEglRHNKMaHPQeGzbhcY5WPQR+HEjfIFwq76XIwqJ5uevdTvcvg1kYEAuqOKrJQDG2bbde
o5srDC1S0c4WPHiDzo1rlRYMytICLk3I5GNoS2FAErkoQuGuh6pn8VRPjb4vltVNSh3y1j+L/Plu
+xp1VmZVr284aJZneCIIQBplMgHTt0Vyl4vvs7l8VCNdOAo18rXVPLCJSqC9YOLIhlg6ZdmOhpcC
duFhCHnyD6VBH8rhRPLjzWH3neA5ndrhm2xRIj2gyHpFbrrUzLIdWnFySep2vo4GGeVvMOs6FsqS
TsRz1/8L2IB3d2gmGvSi1fwZhYKYOR+NCCyJ4TD+42PIFwQ8SVSUxFgNt+JzBL+1xsb1X8xv9L7k
BB/QTkpRS/oGMkZ+kBUxDnZftKH769Oi5eZ4vtMmIQKvX+SeLxdbJ3y8zFuHkkVe0NRoIEc5jFKG
dXzIKyyiDIFHe6X8TYUT4YG5ZHJlnaovWS+QG2RO1ZU/k1wqcfRONmW/Up1LvrPeVEy75E8iGPu9
3fMzFSQsEsTDri2gAojaYsTWCQvhqwbZ+uhq2P/kabH6Vl7xuBywUpy9XWJXrXfs3lXnuYMgnk2S
Qc3MIMKAA2OtYVhrF0OrnRb//NIpE0lxDHibYxtoR69SYiu3eP2CgLSNxLXdUcKc1cJ3YjKml97P
wpLlqh27/1jHXYjLKOlaKpTZyFnTHaorLv3qE4/pOvi1z9YhIJoUm9eNig84Q9LEmAyCDxSq7jj8
Ck0UUSkrm0vXkCnEe7h1sQ3cJMES/w8NrFQVYOGNcAePUNxWkUC2V8dCV9lc6viquIa1LdPvQ2xu
z67rcirvDCflp9svEprpGTKQsHVxeO2qCzNaHGNli7rLeAh/CGcnSkXJyFHJXj5M7xHTuuEosvgj
7Q8hQHLt59MaCC11+0dj4pCLbMfQWRCox+vWmmh/PJPn0/JdUtqnLnut30jNciw3hJdgeqEn83qx
UZOi1WtRHxZ8VTOjMpS8PUj/eqChsq8TLo9GB0Pdzprpk/YKRtTvJdwtfhirrJKF6T4/yMICnl02
09n+OIL3cmc0awOSy7Ht3djHRVEehJ6FpnE9ByY6GmqiCyL7bC9ZB9w/4v92Akm9bwm6w+1E7DSr
NO7PCCBLkVlwK0t0daXXMOhaxslaaccqYUHblVqjzahOvXSD/WEvzPaBEy6/zpdPxKbkHO7NWgCc
DdZDLIHMcymlPrhoMzTFtfxbmyd1ULhRtWRFk8tm1PZW82k1MKtdpF8zt3TXx7mMvumF3CtIis0U
DOm8hrswc9WC6CMgVY6J1lJqjgdyNIXOq0+7lYbiiylyM5WyItqG74RvUxp+yvb5REmbJp56TrTK
Plg2JQj4nJnmSD3MiqGVsTIvqGSxgavQQQnm207EJPiSy2YdJyMHj6qTTBfd9yMzUgJJc9Qv3Pcr
T1xArjArHeZTssLcA8U38j+9sh3AzH4ZHE8MAKNb2C7d0V7c94HI1rKIiN9iw6cRu+o5GwDng1kL
5L7+TTf+hNPEkA9nXhUHZFvdQRWo/pnYL3TRvwVtdNrI//ZPe1ffyTw5gFZAetVoBcFh77qtCMxj
5tlSWVBUvE3VjfJ11exFtB7f+V6KFc1yNde1/KjtPnG/yM2ZsMcUFiO2bvW49toOmJhHaDvrv/hr
+S5WhWLvQCxc+TBMQ04CzUP8tzdcDqzvAf1YlQ8W/EpB0QZsVPxNd/I5sUHKEkC/Rv/e14Wj4Trh
Djv3IC6N+JpFncVD6OfaUY4OTvZH0gmIodjKQzR7gsdcniA6qVUsSZUoHDbLroxcassom+CTbXv6
h/7mxCwTZHustsQyYOAuZT/RV/VIqFdUrLRLusadFjnTBz7ufdKkEOUXaIXFT+sBeIbhuNhGzjjf
dr/rfXvnGVojMr0suZc5YfcyIyltMoCaWdpNV3HK9t88CGE0fh9n4Zfcusg35wF2KP+NbbcHaqO0
WikH31pF5K9Gk+MYXbwlZY+Ay9vOtb1czFzaTcZbV0BZDIda/bcN0lqnAN5xZhB4xFOIDoIBlPGr
/mj1wXw0MT99cne2vd+y2XXtJHClmE0zbol5whO8S8o0BF9rgAMLwxMDboQBmJbd6hdsNTDaI9EM
cZecQv2LamLl9RWeWVvWNSHdxj+PInr7sWR87KT7L57wVEqvSGkXr+aQg88bHr8cp6KqwpZ/+GuU
KtIK0WYw+gSbPaJ1cnnImcapi6ElDtFM+fCG9dYop34QojmYtYDsHbfwdJc1zpQ+/vX+MnHR96fz
NciFk3jJ78Q9UkJhdN6fLp9aLHLUcq2UdBm4VuJvZIysGnvgsNvyeCzv7aJgrr75OZuSgjPhCmh7
loNICYHP3oJbugh8e0oVNjvuO/ano9MAIHOjTxEgfSXjBIUrm8RDIFXrbCRhGefRBHTo6TKvtGqM
6LLe5d4J+DkOi7DuTJUd2+w6c47NNuNcgpOv8yNl87Bt5pVTG2UKoCY6CYQ1orkZUe1AOK5mUys9
0ocVQVT8HZ4tdTX5nkhyUUdiImXtvT3XGpkWS5hS2ag2q1GfnfzFCy5WRfGkhTz/UrbhUGZSJlc+
E4KJcL7lHwBpY6uh7+fTtdyTKeF3/TxL+iHudAqJ7UUp+eEl1IVadbygmedb/7dAeoTFFRdWhjHx
e/e6vZ9Uu73RiwjSsOzrbS2XoD35sdUiYeZe1KyMfxtkRrtWbNpIT+VT2nO79LgpsQRG1At8g+Sv
8N6rM6klFEow5XvyaC6oLeBD08WqYykvgT2w15ENXA+axCDP/4pC+DmoqPXtoNNXiMFHlx2kaTnl
jvGxqwmr+gGevwvYBwEh/36DDQdjzlNCHR9+Vu3z4sDJE5JXpZ9ZLIW8eEN6rF0gi5V5jJ0pqZSg
Lom2InQERgXzWvitDebEuGzJxWMSwqWtKYwKvT8A7N8jCPPkN1Hh6syK0ITJGlTl/Zx3qng6Qq8U
hharbkxsrTSmg6xOy8E6trF8sX3yY1ogXy5WYhX7bITOkw+PR7K6t2twbVM+L2cPihEDWTqXDfU1
BHZXWEiXHIJtL+jbPyd5ttiFE4wX+pIC2Vk2CAysf3DLymc2IhM0jWxawgvR/dXbUzJF1iIV6swd
JfouqCZv4/tBaluvaC/yXGClurAaBTX4YCvGqMRuitZsNbeqDiOlxB9ajS29i7hdQ/Ibd2bPwRnk
hoPjvPa+B8QdQPLAzagw3rkJXuERPJvbcIxvHTU/jqF6u1sL3pc3Ofee04f7Unqiglm0a6ZMNVcq
113CC/xKpBHQs4So9VVFlz4LnmmUAvP15twSxtDt+UN9lfKXzjx56PVfCDcnfSNaWlpoz9WWNdR/
gUgLDCUzER42EqawXmXDQXEF8OzLIWcd8KNaeCzh/HxvogcPZpoiAAc88wZ/vXl8THw7GWtg3cAV
TVStytIrEz3IEpHm45I0b3AI3l1Rg3YGWqbpPxENIgK51vZRsOdeTvQBqQg9Tb6hsr8N4w4fXKDz
7uztsRL7213LodNutpxrEsHJL/AZ9ORiiKTr6Qea9ralixjVtknT6TeJ4jTW4l4EsuLEUIbgmE9j
nB0oL1EG/IvBKMWKlsnJQMCktbMH1on4jWEax1vXNjApn/RD8vJQGgUHxHyrZIbFykzvSQvL+vKW
CZgv1rTqnRwqzOVQdWWnYxM67dp1++ORwIVAWLpTcgTtSFrR7VcLNEBSjryWypj0vLXSwP+HYy6n
9IQ8K557imwQytkl04qT2LUu+aNvuJ8GSl/zn2vPFZ1Ai9jP5axXVKlVEY3IqO6WHSFH19eNfI9P
si0KBqT045/JDztKmhiCRtRDxmqwFsX7cObEUaMjnm1fAoNK0btooG6kd43Ay9yma8mrrwd8ogV8
vM3nHglttJGVT7rzrMO/xSh2BYAIEt1nAZrkjQQEihJ3jdB6nLhnGOv6vBoUFODPJXlBekV2UpmL
fiNko0FD/8JFYjYq4Wb7ygugFJPsmysSTLx4/7yjYLvlJxZwK1MJ2z1gJ4Qp9DCXuImIuN285T55
u53U5KRRFzDPYR1i2PgCjxWn/h8om5pMoHpf7nN/FX4cuv26bcMIgVI4E6PXy59sREYD6nYtn1C6
RZuaVe3rPal+JNoqRQCqJ++4xiVZPn1k0GYUfZBUaLKs4Kq6ysIsCozGZArWC5rxg01p2Mqbk8Ql
6uqAlYpgLEc4l52nfToyTzKfRk77mdC2rFnoKg5JNEmDNcyZ4iwWLc62TmxSfwrUlB4Xs1qegUwB
mfyjPlMytzZ3idgC0gupgPAmBT7EdUjVrjMAP7/YJB05CNjsJw6WoPYEhOd1RC+W0VliJfqw+sW/
sjro8HySwwuPq2kkVJ+BmoVzSOQhFjY9VwV45nfNjIQUGK+u1sdjJXwpATllgIYA/CAoFIg2Z9OI
Xh/Jbtr7R6cGEX4LnyuNkZHcQ27ERcQGufGZJPLwRZpvZ4TDYbvE03sPfbiMdaxFRgC/3zZ8qNBq
S1aptl7h5Rm35/Y+okR7jZe6tBCekbxp37ip0bi76Hg5Ib791b+AQv2OgXY0bH3HSlWoIFfhhqeO
dBdUd6t+E0F41FTBGX8I8Jf0UP0xgP9Ou3uTGknb/ALq2JDf4DaXRhluv/32CGagT1Nz1ScpwGSm
JXu5qJQaCHk72e2HjE9rL1TlwXEf3UIMuMrF9jJvb93U/9XFcLUVUdflBtxAtblP2EFpoft1T/dn
TnhBHm0aI6eQL9+/hRdEjcsClJmrVuGhvhwXxg0moz5uqrO6omLVjUIN15Qu7ufCoGQa3GDQui4Q
wTeoan3z6iyMwrTZldCAgfjHqQzfsAauN1rjpX0ZJLHBQtZ2BjCq8NeUQfbSFomf3/MCrEdr7H+W
3tTmoows8gOEVXPAV6A92Zt3qkjHpzkpTcePMYOqUIjD5W++5OKNCQgNsC43Hm2hoDn0D6grVWvC
co6NmxjP3oBSmOyUILsFIs7vW29AXT1RaQNi9C145GtBVHkA5Oe0Qhh0W4HWzbJ7cYgJHvvvtGZp
R2DrB5IUb1lk30BbcgrwgrPUe6RUxIowq2gXJBc+DkjhDLne+rn9v/HKo9I50dvH5L0K74iECy19
hIHDstCLORleh0b+G2/2Aj4XwO1Nrq/71gIAFwVSHN5CzfoF3VyuIhxEUXJJJhor3bWLxQNk3Z1N
+P5e5/3vovU3kRjQioxgwMxuduvsT86njoMurgRLoMtMuWpuCiCubyXglcD5zVyVHyH3nFUKA/Q+
/Vl9b+9PoExV/T6MOAMqhy+KzjfO2mTmGbA+2mPCmlgXjBo49bi/8NEOFIGbWFVLg/p5/BfDC5WU
rzC2zXJFnsiXc94XBW+fbzsvYaDOhBF58uYl0DtyZUU4s7nV3IJ6Kg28kv6LvP/c6YvMJfJMFkuw
mOfn+0qHe/77ot8Iyk6IPWVmOD0DpjlPnSVOLSWeq8h9DDPQ7u3LHyoyMgS9AAp1ddRciPJmCecm
5ifCiCQu6XMMbqAueWe5uDDu+NqC1XCviEa6e6aqwtlf1ISg03papmT6eyH06Kbe38APzwQon165
g8bDalmDcNiWK2GPPCN2Re4SY9FDV6lKL/QLsETqv1PQVm871K/BPfD2/CtZbWMOjCJ3dZvHAyb6
lXPmwaLVVFSM87NYeqlqN98+0ftKGbyyPfsUBtt061lU/bM3i3FW/61tpgy9Hc9x5eKC6++Q7qud
j1lLedlqRItwcwDeEP4gU11bZ0eCV4HTAVYkwEBChuTrSp8YpxnwT3wv3Irwi73M0rOM8c6LXSPV
bLhX9Sy1zhVFJwm7aEhAqbh/oNCTIR5J76GM9FkfyWG5OxGO9z6l+kgMLUEN5PXBSLB88/TjWXOc
kCNJ15DYz4jvs8kVL482KU36/ZHmnwJe0wtiJ342laHFXTcv2iiJFuvaopP4ijMiQqhCMiIwwJE2
AHS6QPh7n1iO0gnwDTTSAStbX8RIHwd5863sMSti1Bb/+7b5tLdw7In/ZlJDn/Zc4S0fEgPjiuQD
94epQePlPRq2tPtOC57kAe6QPRw1cR1wJGu6zAewucnEAZVNIeSDUFwwzLUs7a8Yu+L2UpZ5TelN
fWF713HstpkOobz1giDNerzATD7oL11RJg8QI1evqFrzrCdzOQaSQbU1ohvfvIKKOiwoRXPoBe8P
iEbZm9Y+weGb451HwBSujgqDnUAOmsf4kE3Gx7N+Y7EhipHem1fcPmpOzLz5YCAQ9x5XQijajCgn
eokiDQUuZmpvedPpBHAGoXLi6bPuelzzY7b7p/QUL2VoIyYo4UZf923bgD3WbZhWNPb6yySyRw8D
KG3XXkSKPo4dUtJnI66uivcXQfUpiCGzo6RGDFoR/PHQi1BezaIWBFf8elveaB3fCXMJUmRTQfdj
wXnaFZDhiXS3D6w6Owfy5yEioD6pfjcHapq93YN47mxkkdExsM1pTLdJPtGDXCfjJWNZReO0ndrg
IpbMkNCajFZfL+iXDNcE/OPuZenbgHLIOIgg9MW7M8kzkF6bPdO0X1MPeTlXBcjpZ5FDWN15ID7O
2xs0q9IPIrn1P3DAkAnsXsU1EPr33A9i6sUN7IxHkhOYThGaQ5GUkQJHKeaM8Fvq26k+xb0LZlKn
HDuSv9Wfxp8N+f286eOJWpWCBErPMo0IaCTvOJ/jd/VgE2x4C5Y7oOChn0/m6bY302nB9EjJ9Qee
Sb8H4jRV4rBKbL5oDTkvV+D498teEYupO1oxKxXmVaxNGSfhaW+5KEh1QhgXa5wYqR+XN3RHt4zj
BZbWsUBTOH3/ZLGQMNwuJ/XqJhV2l+9rvBlWT2IGOWbm9PlJtmV5tZ5DMluHDNWcaq0vFTPYShDL
l+1itbF/a2bvz2ce+aEaqd36l+Q5LRu6JEp9j3hVNFEQp/uYzodDMyrRpHFKiwjMIBwomQGhNaG6
oMBhnyaBpiCg//KiyDTeCr/xs1jXZyQzfDwUZwW9J5hCPvb7+ZKKgyRPabw98Vtn7JHCQ1FEUnfy
cdWqTUySAgVa1Z/3ipgYB6YMK+yugD9K76l/SP248pcudlgQXLX6s7zlFeV4UHUUHd60mqowmQhC
/FEwYRDoFEhP+ZWmidjJgNsYua/QChdumsy1VZ5NqJ9u3djqzbDJNRlgVeYJFjvpmuPtHynPYosp
dXW/T7mqc1emVTZc03cDpk260/6V12cKFizW3ZJjYwwOmuHk1LFnHV17aXqO5nytDGR4hN/2rXia
pdv/Bht9l9j44m8v9pvVPLG1eXNcuEEZnZSKtR+QLZJm9VsxXe4t+v1PYHmC85V8NvGLOpDoH/Qm
gWlC9u3OASyxQ2P8LWPQ7TxMemJYjz1/RGu3Qvppa0yaWqVqwechOIKM4KBjo69m24xcHz2d7xGt
ucD1hvH25ucv3HXIEgAV9CBy8oZ1Gp62Mg5MfkRZnXBItW82pbHWgfrDK3UMc3XOjk/GPAFdOSzG
S0hIhojK3G38dmi3o8hbRDte+movn/0MVPqrJuoZl638Kh4bY8s93sEVzt958JTK0AXJ0UVIYFvp
QVbrRiJIEdP2T6MH66laCV9nUIvcp8T6qaOAq6vNoRm3EUJ/WOgUh+5PO+VQIJI1NgP9yQQN+PJM
6ICPQXPH1cMiabuy9JftCDY3S/e+1+kJ0bG/flKA4fqy2mXc7vL88hAMma6u90aJbKjT7MAfZVbe
y9ZoCicxTZhaIHsEoPfG4JEjhCvtKSfD5cP0O3Y04zD8kcf9n35JDjsulwDo18uAjJ28K3kt3p7G
P6qbS85JiNrUNEOu0fnAyA+AOxdGc/T2hCAbeCwTSVDSt4UDIQOg+GvxK6WvrUzRqotQcmJcan40
pfgiPhCuEvbmidBIw1eTPtUOQkfb52+UVCyLOWie4dTHYAnSQw9T34754ixbuVjcv5W58niJjzwq
31WiKmaAa8LAYwBBSGbT8Zyui31QSdLUdCbqg5rpwsLaKwFhjlLoztSU45qxtzlR5hYA8eORV1/r
RQrGQdH7TA+pooDgNWPAHaP8SUPvO46R7KhIX4kYta3+4q7NOkZg/jZmy24N82xh0PfygmprjXl4
4qWVcKCU4yA3QZpfrtZqYWBwoOB1jpcsdhqSEUsnoKTQ528DU9I7yZt2vrdf4PC+Bxu+ZnI/mtBK
cC/5xqlcJjcs4sx9Uf8Em286ffFJcWmZGXFdmUFd0FZWAcoO04SS+Sow9c4CUC3/eyARItFTOiVi
ad4gCIKiyjt4s3Ivgtk0ZYSrpW2wXKxCpDKqS9MPaT6NbYxmephLHvDLG9fQla101igjI8L0udjU
AKu51dLSqKvoNv7Md9V1TWAZsmuZz3APjljRMyuxNRkvw2er66cv3wvDloi3IP0LDZzD34YZHPdE
QJ4Cz7pQOsB2QykYn30um0yPK7OGuwVqGb+wR1jwRXZiTYTFdMP7eQBypDqkf0PWE2SwIpxXpmUN
jcbZf2vQ+J1xZcdBg/neGDLowjV8QgawIA3blOa5j9pHFylf5lAjhAgRezuR/vQAL2yUF+jgfX0Q
JzXoZpXcHyvzuCcXr1nSSv2Q+Or/8sJu29wOfS0J+pQI2KcrtexgHU/Qo3j+LV0GagpPqY2cMiX9
Lh3Vlbm3p7pKmIXJx+dHOpYxOk2ERS+rwsqjnjqIxSNuvQg272PAPtvlQGHoSOwjNmp1HTheJ0q7
/qAYaselGDSPBAfCReVX/bXDuIXfk6aTOfhV63EGHxQZRnjYf1uYMxLoLO/KeGVfXTlYH0edd/W9
EV1v4xb2fHcs3dQl4oR75lWBPpiSeFAoKJJDxNBN/M3o376PlZzbpRkGX0iSSFoxcywmcbooSYTm
7QMuvC1WwAKlmfX5vW7QPh9qULUsQkGjZpC0BWP2C1N7PiUiBDPvU4JQ1gmeXkX5kAPVnbO9H+sl
YESU786xQxvyDmNAIADs6zd3AyDa5r/3X4S5sgYmzdCy7GjEhET1SfF1Lf+vve0mi5OCsix1AMws
mRXXAHTtjYIQj9C/eCriqvzt6zinWqZkHREprAR1OJ3p194hTRa3LZcNFyhDMMkkQPW5+0J1LssO
hU3dAJWwv1IX7vQdnzPV8YSPxRTK9xurC6yZG1xUVfzwLKkNXmsP7omqcbAHHToKo5zlfhmr4rkY
aCyrqC2AGtjgWessFRanaX7qnrH+RGABdMtywIpyb834NL8MnVAc8zr+Q01V7VHduvQYqRv9Bes7
1ZpeGax4iCdXhkGMdn3jJaJAqQ9HWPkugqf2/rlWHqX2EVDKZE1c/5vRgvmvzD0KU53x9f5NcXZA
0Lk7khsN+ikXNeIfwrpjHczRm4KsSHEJYmeWQie4g7v6xWT9c4jDEQYNQJdkss3zUgVLoN9uqjg6
kRb+6XGiM3Lpzo3TvQ+dARx7tQJNGMDupGpemVNNM4CRqKgWtwwP1blwBLD+lBBil9843H9MvURG
svyazsZdzqxXXk2ZV9s73Gsk0ZEh0UbvfXX9Do0Jerbqc0QxwCeUHJWvC08zqgo7F1xKiRyzJziZ
uiFyiooYE2v9nAswGdBcTJciH/PnPyZ0KuslVl8alcWvuMzT3kQXJ3/ICSnALxVcOLU2TuZNW//b
Dq9tRHJghDmlz8lvW4zKpQPkDz4Nb7tRI3w4P3c1FUwfVDrrS6V/7VlVNT4K9GI4v9TYZDyVl4Kn
0zLj1Umzn/XerSYufGr8X13e6P5HxiveKuMN4XeSoH6uqetFujmdj9zzYIQuOoLqwkbevHwneYtV
8oAL8N89SvyNU8bAqXJ7jaXy7IpxAQbMqIulrasQsO2C2YH+JQ4aaOaE1QL9ZD15/meRgmo8rdjL
e1npBAXVTdMpWRJk/1kfVoAyNdm8HHmR+EZgWBO/MbXTUuhpXzdrannBQ6ig2Uca5p/veWQEpgF0
fIb7nyVQjNFaiWuAkV3qEWBptnJ5xdiZhkiHZ3fT7NK2vmEYee3sklApyGLY/3XE1EmAEFpLv5QA
0tgoWvpURbXM5d8IKj/MtcvGYcefbro0v5qEccqu64DPpw/RnPKqo7HfmA68GTj7qOJCcBx7IdCm
5qWd0tCPckIo/P9qihNDU0dcCnWA/SJYpXai6vxtPUGgYS9MsB0lcMC6Tfeecz0EzTbpMqwF/RZR
kdhMXi8DEMmr7tgihvc+wvHj03ickvhnVrcZpw4Hei25yq+p0AYXacz3VgZL4uZ3lWtArNMfPnTa
HfJaz/oaOBa2WH6hsZMJLQB35pYzsTJFKptJufiyPd9DSvM4D9z3Uh/kDX/bNKAbPKqJpAv7/VFn
3+yyO/CYDksEmfCe4LwIWIb/iKteWOSnx7MFeoJ1qsq50vhxe7j/NBE28V7fmHc9ibH1VcW4eHrv
WTK+ae8PX8NkkHQ5pVaJOGCYOtvShp5G6o7BDH3H3PkTPizUIX1+Z09DoXnmRhVt7qJdPB6ZFTdU
NfPJnG3PjQoDgvGFf9Osip5pmGjvucuDbAnOypQLIQbfIrACp3yk0QzkE1fMgFO6Kidlqs2m8eAo
dDXng1+9pX2CjofkBMmStIvegGE2GbiRf3we7ou7/2JY1AbarumAVZ7p3WBo4r0EJebHHxDGt8CP
rXAZ7kQbtUZo2XUeBCjLxQ8u6PnATlU4uKtjIL9vNGRmShNu0fjRsaIQ0l/vmc2DWNCfdlAaNAQ6
sIcZepzHeKQMFQmEXpXWLsoSTK2DgeV6FsZNAuLvqp6p4nF49G6262zhzspBWZEoLpCcnzDMVOu7
KAAJizCeXTWKMTm8JnSgusEg7X9cnca9nNzeK9I/tMMSi+5+LwdNF52vfwGg1rYdVADB68Y7SOdn
hEzFVYFtfSl+BSsHjqu+W6rHViVXi4vvdXJ0g+op/8uXPcecSsOsGDNReQGcuxrA+8K3s9Zs7HOk
3yYXZpZqOl9bMSH2zzBb2h0/Qa6Cysb8r0x1GjYBM5QiXAq6vVNJYy79xjR/Ui+JhTEMX+1snkm1
JCoNoAjEusigCfaabv5dkjerAKFpbiuqrgMUGWHfbhnB3QZtLjZCE0xUfof2uCTKlu3MXW47wR8b
oi9cTAb7JoOcejlKl9aL8n5t/KarQX94YM+fh78Z7GCY5vMXzxs8qKgyStriUlQtJiv/2DxzTOfl
BcfRvDLOP1t6EpXjM40deDD/raEs+HaEvXmXzuFv1U9W5ewOqqv/9oSxuh+zlezY43gkN5feWF2u
+lGNgdez+Rk1dtRp4aAc7gNnJrcCJY161ansyTLnnAi7DjPxNE5QKWMdlWs8ymVFvhqsQfvSbB4+
iDr1EEOT91onN9oMGf9t0+SQ8ewVU1zMksegwmQP5NpL6+hUyPYzIFruBdY+zk/zF3yVATxPEcvh
ROkVirRTP+ZiEcGf2/Dc9js4AmicZnTgAw3ozcXlGOyG808JVUUdKKgFRSWoQhI5ZwWwRD0xgBiO
lYkWKnYNnL2rRNRyujQr/LmCjOq8K0/H3oP0lcOysmQ9z1kDHrg/31uwrGR4PQgLy1y9qK4yY/sp
NsDvejDcmkwGX7ie1b4Bf/0AwB0Wm67lNph5sy0cF6fB2zpToplYVkcXQOltnl9PyznNCD+a1Qra
Da0wTpW9SlIkjSjacJb92lVDN6OAjqiJOPVM/maODKa1LSxke1JPaH/rrdieOhn+Cz/JqMp364lO
s6taXNPNbSe5bI8NYS2F/Xr88M5e28ibGKY0hHAtrIaRpudWinBDd5FEZNQES5XeQqJIMmJXhFZF
nv5V3gwGQ/BZ0WFTuxbzdnTquck78YYoXLKo3n8YBjszBBJb9yP4BPH2E8/y95HWFkvTzzyuMuB9
mjsZHmPkQsFoT+o0DKC3euT3qPcfXRNOLVpy+HcIYO7Q3Nagmj1Z9Ga+dyAafEiwxHo8FYUSNRZR
VqM+1ufCWRmd3Y67C2M8ol8iHGJEAi0g6o2C7nZlC5OD4OkElMMUvezDnfsxgprYpAN/zGG4y83a
YqHk33+GBjK8Cbozoso93BzYWsdJNNsLw46g6cKF4I2D2gK13Xua890BWLWWJ2/Ki+oY/IxEDtpF
kvc4cKK3u4RbJJ9hknYc+mjulW1yINFtDOIRB/YCNH66vh3CzZGeQe0WBfsQkwItR0zvdy1hyB3M
zeEVtFuoT2VGcmBRV2L8C2PAjXE6MXY1bHbJ679xsXQpevwOSxzsScQ0+pVryySZ+46oaRbac3AI
2qNFXbXcTS4bnjG+WESBgtrlwivKv1ahVidW4bjeJry+KcXj23xZamd1zI5DWr8yflsYONTaM2Ma
0szsf+xFGfmUx9mU26nTq8V6VNubz1e6ND6zBevR1KsfN2VlFpJfRCZreGLrmFFfQ4jeqlxCANF5
NqdRsdZ2T9/RkoAryzNxteR3L4ZgYAN1ZUyxHdXriuNG+ChTiFHJ/syhFDRXkn4M12YdhvUD1Saj
UVRA+6gILQ+4kJ1vYaZ4XlvSvk9Ux76L9bhEANqWtDYlohbpfAU3ml4b1Rb8xrscGs2Vs9Pqns93
LsxtHXP+PUKdUzZmS5b5AD/fDYPCMj1Mu+3Ns1gsS45Ohq62VIc632bw+x7V2mDjJckJWMLHRpve
M9IQvir7BLIiscGpguTZHHDrVs+7o2r6SMLORAbmCGkwbPqrkX302TmS1Jr7L4/TJGOQ0Lf63+Hh
qpWlA8Nadl3zuO4HAMg8ZRxf3w0Aac0WNHQUeAMf3A2x+o1+1uTaoofG8wV/HjpPxxcDzLSapsIH
gfL2j//aebBfFRGthsmyzvUl8SdXDjI8ic9elEe3HyP+4/MOSPAYexIyCz69z4B6ad6hQe8kY2AC
AqkI99Kl8hxesOXq2WtfRHwTMsS+XaCJinurdFEmuq864McfCHHambMB4CGsHe/e0abHLQ9ObXyy
FWka1bN3xWUExAfmF1UF8dy+R57WicIBsx0iRKoDuHEjhbQX94OOMvr4JkmYDeSnYvcRUrPqiniq
111H6FHoWCoIxbQ2mcmYhShnToWPMBY37ITWev79W0Ll81Dt2LQhF34ZOYAlKWRJX2y9dg3m0jzM
o+ikbbvvTSutyXJcmdxyVRTHrn3g2ouuIMpaE1PiIhZBECtLKeMaSsNDseF9on9FxxxK5t/TjkBq
KeSF4AnwT7mlA1qCn9Zo2+k3FqXwuHz2eFtLfIcdRrd7Xt1uTlBE96mJnQSUy/sTWWdKVcOTpXL1
d+wFeh/V95FR8jiLXdxoxaKTXPGJfRqqBe4hAtPlYs6KTjsz6rZiHaPwTObIRQ5f6pJPxGQLr29w
GIy+RyhYieT7xsENM4aM8LB4G6hrS3mOcI539Jfdf+RN3DwfvyVlvxWn8ARpyz7RskAPH6he72PZ
16oULDzEfrg6wbufEUSkwMFiDBUEY8IkUeKEShdLq1NaMg3ojk49y4k94VojKw1IyxsCY7Meiwu8
yZxpNY4luf6QAS1N51lsDeicMPxl4lzqNewEMWnvcxun64U8JYw5rvGUpFueqzpoaCCxb+peQxjm
PwP5ycPvVlJZGOQc79JOtHMc6hHjSXj7T7FCu2UbigkBZLAokfPqORjP77WLIh+F1Ir2I4sSY/+0
HNjFphoJM1aIGT2zUFSckbLf25H8UDyI0/N7RfTCePeyTTCY3cxXpORfhZqwsUss7Ipa0kWrfeBM
fc2LagXKtaUuYJkGLEl2m0p1kU9tDfJDXC0mPNwFDhEThBkJSAXTTUynDsmvolbJDQ68w+3Uv1S0
1iVC6sS1xUaq30X7OmVVh1sIFVVlANPAmAgUoANpmdlOaiXDAGr9k4NjGaHX6tYoqT/ARQ6n4/XF
ZL8F46yl5bEtNjNLqLYsKRxvlwRJbAxeJRpVXmGy8a2pBNNEhSzzATsgzUXvJAfhSX6MZroWrh7s
X+A0ZHwv+IDz5MelW4u1iaZeSbVIV+Jc5XBQX4aBbIP3D0y/p/mAsjU3okyeB3QWcFhW1R1E8mwL
ZNBsSs3yQr/jCoEAabrRTzGz3oY9FWIs6Lx9kDD1jRr72R7QlgJiEwY12cIYAOPt9OAOoGyX31Ze
md9+tGP4G0nd8zt++1rmi6TFRyAP9wzf8r4glIUcuxjJSWJL5qMMllF3YV/koqAQig68LckqO9Qc
Zg/mQByLhgremo19Tq5f/DfLI3jGN5DI0zEwqKj7Y7BSv6rDLjRr7ZxNxP2HSiN0E4CYp0ZJJ3CN
BMWvDT7OF+NoFQC2SqRh6neShHP7qBpVjpXyNQk3alkKbIQCTK8SGZ4s2fiX7R5QsRXuNJvWHR1H
Hu8oP1lsz3sVDSqkePOHW9wx1X+UUAgal6CTgDBNiOe8avTR5Ij09p2mKGKjgGPsp5LLmJzAqOkM
Zfe9P4+SWE7iSHuDtCLE2gYqO3D0G49lSCI8ZjUIjNXPC7rScQeUHHnPMJlyAMDbK0smofMBLOoJ
DDuy+0tu/DvKylTVg2oD/z1YeZ1y2tkUCuXA7pkp54SY6sgukqBdVGMpE54j5dKQKgmZnte6Mnta
iuBTQ2krj09t58hu4n/eWt5ZLMqKAIcaQ/JuF1E20Fa3QjuivhrixA6fqyF9ZgXeefIRoy3oiM4C
uz+8NdD+nfWDOvhRx1avFgfSYGMO/uHTUTFXmURr3lFOYa6akjnw+XDPnI1z7W3S52AV78quhfxE
mnQr8c0GvXxcvR7gVIgLV0SSDOxgIHbP+CvQaRyhTTZLTkCHl1tV4gDIbDXJyd7kUEY4CDGs3Ymz
OSb2/HP2kBzLvQjqHb0K6bLNXZASkRT0EDHAkBFAqvD7ynRqOXdR+gEOBoNNIobGWJ4O9NK6gq8C
YNEDK4uN5So9T0MhOruNDXtWdPZ0mwBhpQl7YiEG7vjxTLtYcQ6yxSLtl+yAx29yO64wBXcmUnSk
/2MCwxDwYdDWaBQESwyDRoSdX/mQ86BYgqK04EA/xbbcIvtJqOgSvFWy3/1Qx8Q4kNV9kmv8z9MY
ldHp96QSVV+6fO9naH1V7CuDCSlVH6Q2IbCBLMzsjaYR50p5a4E9ipW6unu0Qf76eH1Tu2bw/pbq
6T4tE+M46VEE+N2k9TzYfJO8D/BqCgQ/VEI2HSaShS0ymae6RscBJpNEzPyM3s9YoLfxELF3md7u
AdexdHwxpOGfVGHGE0o+bW8xsjxPZ6SHzy1k2umYPQPzdTjO2xmhkdQHmyL+W2gUL+J2eMCJbW6P
2gpz+7BAiJ6zNRZpsKoQXRrSBdSzYCXqIlLz4Sidvm+JHWmsweuMkSz0vLsNBqrg4Ntj5YY/YP/A
JlhNJW8hccLdUr6PUq9WXoNDl6dFaOB2D3k5qts4pqNE2i286l5sp7pna+fngEKS7EWC757YmF2D
aeK64Vs63fFkVEuuv2api5KBEcPApW0FpuTu6xoEbcme5tCV1w5Ke0jmxXCTCizp7KbbfHfYpomW
BacjmOmI7bfE07otd2XoXgH5FQcT3bf6uS/gkGgsXCom6X/2giZkeoMjfbcNMdJJIKAWqvZaAc3N
9qYNmMtlSw8L2VtputNyBXjV46TtJqxwxwnjE9o1XOr7iAdm4oIJprrSmP7/FBztBwRBRPPfM665
2x1LyIYxNpiafPpx0DCiGzda8v2vj327NblhBdVxyZH59LNh2a3bjk0CN1LPp0mZxXI91/F0UQ3H
VT2kvU28PGAmOuS/Ay8optLZLB4PsWr3TBqGcStBvHiNdzQFK75/7ToJArUAswg2Rb/GpZT8CZSL
Ec1d/SAfbYOwvPS0QGjLpRVpA9UZt7kR+9or0oQKywQ5phGrB79lrwv+LEgXcJRerZ9KpmktIdd+
66Il717Swqwn3Be4RzDDrs1XfqIi0gSKWdxyPBqdI3nSy1AfP2Rj3Er5l/eXvEsgucrQe7scDDvo
BThym3Nedjhox+WyQcr2p+/qR72aHePyjPejRRpATbUekfIJKpBwobzJKWBh6ddDuw649AbJ/1UE
nvxrnTqfuRgXFjQzBsFr6ntL4SXz1tDKV8ztaLlP29ahBtYKMuk6yoeem1wLWQA6kPP5kJUg5Tcd
Lp7Wg7n964+WPATmzvojl4oALkpRaDscbv/D3+CH9p8IaLJeN8lxFaXB2Gnl8yEvtTRVkz9inX7z
4SpyZzpju2OWHyDfcfevP5eTE0cEQZGEQRhglLYfUAj+mfMZrNsQ4hbxxvfzHM6RBHeo6n7kt+lw
cA6azKCaVVwdZquL/JEpdRgqE+vqv3lqR6wihLTElnmJgeGQtqWClNcxzRTYB9utywZh+xhlQ/VW
QE7qO0lOHL83gid+EXesdsMQ5mNVTSH/lbiFropyXWgtFmEswe99GkfaLK+JxPYu0c+1FY9hb1Kq
yameEa71nydgc8ebCtW9D1JS1JDTN7yFwo9K1Zx1ZUAET8bFLjJuPZm1/rvEs4PV5F1dvVU765V3
GA9QJOHBOG/vVRbj5cW1uKUM87XUqL42eRFaSPwVY1xpIszpJfuTWjCz/an/XrQRdbyfPALB3aNN
aFp7WT7AbklL82C8ilvcArkEyUBxvMA+KJHX5vx1aIi3bFl2u1AlBk7FLaLYzZf+Gnc61egFXGpx
l1XeNYD72y9Wcj4AKobvl8Y0gMG0WKsn3shcD07D+PS8t0gwCWkgVXe0W8+qQFrWvldeelcAGkT2
N654QHwwAiU22eMCtRQNC4x/c3t/3tQokooXiff6yZmEfVxJ9J2C2BtfuaAGgEwcpECazVvupdVS
7cnDE9ypGKJZnQ6UQhiuRUp6HJC/t/tsVASQo/MlBiGeTlrMW3roWz7lc04EWveqHI9mlv1Tq84W
Hjq+K7KJiEb3ZU4AHWNp53xwYXsLamVImgXkNdgA6Zghkfye2HkQntWQ+JQKEPZPfhZbEx+bEJ0M
hUgQhkwW+/qN2XpufMzCmLAQSNar7egl5AoWDn3ULz0XrqgS0cwZKR485X/RHelcBiqvyq/7Tfbf
Yq9VgYLblRx/XDXbhNkTdLzDoe0teH7Lt89iKjur5WKsALwgojB5nOO079etgZNIMrAVuPQh7t1i
XlYAGKSpp4hVhYJAygFf+p3z6hKbWDjqUFcLrpHTJQ9dX5lB19i2cnpVj68KrChJUiG0DAu3icJ+
7AFTGIsmYYDlE7kOG2lty1iiLLzJCRnJEfw8mpBtdCYkbxhYA2jNLZczNULRzqfx6DBdfOmmsBgw
ydvg9Pu0oEyV+TH6u56aU99OJgduI4VwyWwML747UPIsADqe42ITN9NnRNjdEImTmN6wyMwBk5jm
vrzULnecpkbX8KOZISNfI6Obd+4bNfx9Wx3c9x+1iPYKpMrpQtjiWH7k8tiIlzq6UnRmCMgoDZH3
k+ZSDAgw3M21cXS6bIiaAaVk2duKw+0nBz7fokzeIqdlTCtcJo1jQkqvBJLQd3wV7e034hzKDF4y
ANYld/VLHUF+DR0lKwyq2qWxcU2D6DANKNip9smPjWeWsYUxbk1qUMv2s7OLAtsic+asH7yTwoEz
L/gh9LLdZg4sBIIXa6KSSxNd1nAkx1W5qptvCx6SJfr3y9EsazUstmRyMH4K8UbP6UI34CJQa46w
0mDAWOR2gatTJGTyQRyN6atboAtfvPiAbtN9MZfzZJGH1jH1AIHvA641kuOYrJzimmOZwFhykXef
5VP3NqyxhQB6bOWOwV9OKbLvDCOpuFuigAYKA4V4R+PrpUdtclk2sT06QTcWAdGgp0L+Eu+q5R0o
61qQ2slQZUNj6+DI9KmfTuQCRGZNB36Hccrtf9UpiRYYqDAK3QAkaIaUN6qQrRyZbY4Ro38ptn7P
KWeScjmYP776QQ0ki+ytJWcHnf+7h69GgbnTDcF9GtxfqeZhl049QyNE3PmhrVvorTfwQD2GIkqM
oS7Wqf9tcGNVwmfXNZgrjdMoWGhMO/2LmzJYFS4Uq8CLJ+r5IvomOsBPQw9MmJzPQmZfp6nADZG3
/FwutHRmFJY/kub72CboIUBj69IQiELBQBHA+s9c9IUnK9eZCQKKfuhDPURrAiI+a5DkchJXARsz
zOXPFmJ63TK7VlRZHpWPUm5i+VZPLT+QIuE7YpsdGvvfP2roVDz2+sJ1LQNEGiO+rKU/S+MNdnZy
mjS4ERnVJ0uifH/5Enrt6KNhnXKXRGJGcz9Km5/FYCriIyQUMZldscn3FjS6uV4cAsm/p5pmIX38
9GOVycNyerwQ0/+KGFOFgwcr3HfLBkb1wMzDdtw68muiowv60ynOmae+8wTsonaFvk3NXsrkpdEe
JHFGkKNEb11FUhoKYtfvk31d8/6XHq//YxcSCq7PkOHbIEJ5qc4lwRSfGzJDAADO33EMiP/IBoil
X/hV3PkhpsRfiOe0VlDHipATuDP4DU6Ncmtcu6NW09vRU4CHPIbXRsCjcY2J6ujxZWWtjB+KtiMV
xGonbK8/O8pLPyZwuVqDR9tt8BtBYr5hv0RHU+65xgTwUcir2NAmXkyATXLYCQk/gTAziCkgAuGQ
s7PFKz7dbB6hvOoWdw4fc29sUmEmnWoC/BwMRyhDAoKB2gh7sH5htC4jRK8l2yx03wWH/5nVOdXx
PI1MF826mJB/lbLcamrfuzAUo+1JGWwCAQAMU21HUgcZa/AYoockbGcpROHuf18BJ4WiGlZGB8lP
gWwV25/LKv/LDDZwqdx4vNvIMeonhhkYCx4JIn2dljVs+np64tl69ddMq/UR8h106DM9amMu8f3U
+TzoYgWJ8iaegGjvBE2jiBFpQ32a4v0zhY8A0S1EXLr+Am15lna6PswoBavSRADYg2TJf1g1f/rM
35p5i3M3lTxOrce28gDnjXoI8JWAb32ZUbj7jbQwWORFPmUycTJPT8EiwmfLdGecC/ChkzIcMjyq
L5LywOY/DRcPYYnFaF31iLJDQb4ctI1KGn12uMawkEIc0Q/A4KFsmYCYjv0n5QXNoh8DpgCEm3z2
d0N5beWcBWHK8msEjsNnDQ+9TO8p1jcGoPT6rGFR3R0PJ3792vzKjXTbWpXtaJ12L39Q5OupooE+
4ci0gqgujm46L5h6EEpeakC18VXsmkTWeE5kyyPsOhF70vWFc0iSdBwxoG2YiuVWXEV5Dx6VCHs4
3SthDIb6h+n5dOJXqfns6AVviUozsuMuvEpsbtECO5hll2EDP/YNPl9i4BaOFjm0Rd0GE0qnu9Sr
WLz6bNJeZ8dEoux9BoJ7tGsg37W2E0iRaBHCsmSpEf7cCgyQi/Wv7E7R2nh5QBALOss6+dFtEB5X
/tBDB4HBQybgdWCsu18X5jqnpoFM65jcq+17U9mDEGHS9Qs7PBJE6GcBBuRPY6ZjOdTNdGXI9Wpv
wwvpyVFkbuxWgjA0UIbUKwHwO/WDHVwbddpppgnMJbOdH6g92lJZ4tC09xe38cQT8xey9nEaKL5o
dh6+IjlHKb8EHU1TIROutjddLo87mUqb2OMjcZA5QYCCb07dt/hlQ+m0iwjVuOua2ULFMxgXa2zB
o9J9cgHka1AIUvBNQLAQaCBd4gstuuZTIV5JBTu3cu/Ev+iWcuI1KNsAGh4BFbBCp576nq+jRPwE
r2ztiS5dL4BP9Mc6mcKb5lxVGBer7R3+lPaJ4hg5YkugVnlkc8kDBGnzlORVfyjnBCMwDPyUo+op
fNihKp/tqHABgib1Vs2FvqG8q89LmhpKTYilOR9g1ffnK0YJCiDPWZFoOLAH95JeId/Sm3aBcIy5
BfCZwc8qfNglUTa/O+hjziVMnkvWe9CHngXKLIlsDQ4MhvSX2GmL3bc2+0gy7lhvJ9/7XjsPTHcq
6+q79GslrjCm5o4HDDICHnWfa7+iPS3ggk52GydoNu38Zc3VHQnsrrghT1XcKyBe+5OjWeSvNGNX
lR7CpN77doBYwX48DkPOe45jFNlv3XW/IsyQsUT8EHxiqDVvBM+sYbywSuoTwNoluDIOPgt87z8H
hSGjH+y6qwKfZR7Ohrn9jrlQG2z6VzjdMVWbPIz4Qeious9hMdl5TMVt9jlngl1MMVDr7zqtjxEx
TsnyQ/yxV+Wd935FzU/FIGPEJ/jOgTdp64vqAsjJZaslfDY464ZnQI5Gyplg3Z1Wy9FHDAi1Ei4S
9HR9OtvIlE/mZrPj6bUL0B4plWb0n6rO2VdooG2TgwfM5/CWGuQln1I38Sj5HAvbD0r+Y3IqakyC
n2mm+DBWKtXovQyk5f6dmTrgletNnXjPepPEfoZ7QrB8IqOuIvKSxvcEGThJ6bUl8B4w71BWzcDs
FlEZslOUa9RlgkAZHlIfbTIOHtLSQPR8zEDrDfGX8UmvhygFbJb9T+FVi44b7d1Fdy/EHYzvzFwu
RsiNiDsrSC6OKVDYGxk2GniBl8kWy7a+fK8wkpdJxjfBTwGtj1k2k8fQ2izHyIp81j6BEfckLMtv
wpxEQFTG9v1cXAJ6e2lr0lgy/P0dSByPlfLMjyg4u5UMMLLVrjsnvuxaUYqVRxlhMw496YlJHbuj
BUYGUsZM2+5CBj0O/cMqxGfiQe1f5+iqwYam0cTTN6kap9zukDlesWRkYbY7/lF+nfRlWeOz1pe+
Pqrmjvh/roWy3bHar2Jj9PaHppD9blj2Y3tg20VIqSHkrJyN2gJ8IUV+EXVGKemAGQ0DWoyrLp5c
BzaxXeNy8hMwC10jU8qVHg9grBVnjaZjZrKrw1oeO4yots5Zf7Ve+57LO9pSosOHCJWXyGAO6ekK
xeEPTqLbgorKkhL6lnMhZqUeTDL5j4IIvBiDDUOYO1DL6eyNBydCea2rNiKbLIKKlGxM011Y+I4s
1O7ZjbJrHVCGlimZwd0wBqH7My8JmAA0lYUC5SOouwHZrRBz6+6md7ReHb3s5HU6fooHEjoQ9LhQ
xLSniPq52P1HIq4FVvN264Rv2+oMzx2Nm3gdoQu/nQfsBLqG+T2NJf9s5ga+JRsBHueRTt9G05GI
vL/L+cPUP9WP8oVwmQHWYzsr+IbhXoZv6tiPhmFbNj6U4hN+ss2GyPifZFFpAq4mPPh2UJZO0+mX
AT+yEXMI4Czy5D98r8lQRzfnw788hRmxfIq35O0XXpCv0kIhDqGO7x4+4sCk6TPiH8votmG/GcT8
M8AWFwubtducMSwSKfvRn3ElZ5XjFGhIiKnb0+1omAKqLC1YnoNRHITCtibrCMuasJ6VqMUhmRRI
rJJt25zkSlz6uptbrd9XOJtJ/sDzm6t+qzfBUYqMeD09vXVaWEo7/Pw7KDMtDtxv8yHQ4RiW0sIs
38cWt//cfTKIGfwUziLV76EVLFUYa45V2E93IVZdDzrRZ2E6ZG3p17zX6C2FqaM5PTRODR/nA8GG
IMuDC5EAw/9x8Qus1vx+ilXgOrI4XbPY6Z0+B+LXz+ks0R2CWLUrPgfuQXOum0Kbg951n9VvVvOd
WIazkoUR5GHT7Kl9v+oWnPBjP1ib7hengNNZPP0ISfaeeY1gEJ6ixVL024xEdjR3oXT6LYnNga2f
+DKutvYvJInCrvlo3XAu7YFyH2qfHJyvezAzTpcHYf1bhD5fpqLaD7f4loQrgqKaWG8lWuLxgTDu
IPpY1H5LwfbgSWOSSxU/T368+pUkoTQVPluUYzdioniusx9OaTUf1HcZgGsPlHQYfIVg9ZfMXAWf
bdzICYIym/WRGiD0NR+w5n2N4qmBoHFvX6CBxn89xD66EHhmS6AlDpeVycYBdbLJdZdqTgqNTIz2
rOHsfKpnS/X+H6cgjiPYxcKMisZSa4Sl47eSWgkiGGdVY+R3diVY34uLVTtSPslSVawyrz5joNeY
IWPVYXeDQl4zBr+olQJz1IcyIWNbA3ODGIg5+wBZCrhiIDVOoojEWFRgrdsO+FruhqzVSdWfeqCt
PIBAie67BRmL/GzbUba4MSA0sDpM6D1mpGPOJCtP/bVbO1j17XrQFEtsf4uTOiX3foMnQ+uk4kjb
0eOOD0IERNQsVc7aMoh2MgHQBE2X0rG7tfv8JC/nbEwkPJCkK24b6JqmUY7K+l50VqGvmpERqtgI
CEWXGhQUdDra5TWfeZM1PHjuZAFMkk4bwA0w7jYtjRSTTIJhtw3x0C6lYyw1nbyjovSAu7kpjyJV
1udIkWVbViQb8bHs8zavfQhBKh+BBk52GGceSp3vsYmk/YNx02Fpq/8A7Uhizxk7G0EIsz619ONV
rfkB9ynIGXxdz72DXi6Nl+XxUaMJiCNj4Vk/K/TA4HSt/1Dy4xfJQblL2IZO9cfd28PGRFf7gs1T
Nd/l06ySVrpD+J5fLFNkAZI0JxZhdztGiXbHVujo0JDvs0T7vK+ZZG1/EsjgNrjm5E3fQwuukGg1
uZFxlSCtg/9IkzcXrlt930ZatEZyVFzJeobcvwKWhzHZItpMq4+VcmpXvtXX4pADi/VNKFTLwoQM
McrbTCsa4OICOK8f5U83UwbgQ4oczQ0w4OwyqT1N27VBwsaH87orVJdUhOWKLH7AcCVVpE6WaA1S
rvmy9/WhOxl722Gim5pOtBrdMzitEM1yjRJ2VXw+7uE/hgByErFLi+obpvojLhMJBWLrcVLDgOKe
QOLHJ+A0sI+dewCtBXZmLpFUft3vpeZOVATXsHq7GKKEZVnew8ezCHUIbrFoiPvpdYA3i4/W8RFS
WP3Tco+u8hGFZK0xzKmLFqNzpWbcP2DyAaUQC60J7OZjSyWkDvaxe2VH3CZ02bbk3o8Q5OXaq5zx
TSze4Bv/cduluW2MDhxBAj1HwqeNG+igLs2vHN2vJfxSdNjOu5uNjtSOyfPpWUdbAR0R8IvQ0nOZ
5t54Ytvhof/bkhUhm8koo/sCINgCcWo7puu0QAJ2EoE+CY1zwZEG/pCCfipmISqDSPODuUlxk9iI
RmY/uU3bOb6ag8xm0Gqa0sR3U0V9fRIEDQ/HvWjczB4EQLYQYnh6hOlHclkfxScWkrK0zpNpCZgm
0z405jr27J1HEuN3aFzKwsJPvD5VRvZVSbFnzPnkw2+BvuKunSpASFQfJPbggL45I5QnGWvjvbBG
8jDDYFqUfBRTE8DiW3GT82+iObaNmIRXFKzzxFK45oxqI5SGMU/JW9xavCLDZjXK7rhGlO+S2RLy
Hdsz32rZOBOvf9/RlfHRGUk81LvG4//niuiZme6eUzsouyAtl6o6SrfTzdiIt10oL6Mddvw63MiR
CR0sEQlNlJ0MHIQm57I7L+kiLPk93c68Jnth5C/mo6QUh09tD5LfHtJJd+OHeDmAqw67P3OnsREp
yZIA5wktz5NcoLwVge2O2+UC5Qg7lU5vBf5dn0uIhKyIKtMusaCRHdu0clWTwWn6iSrqzN9MJjjN
xu3CBhIwNN4clTQepjGi/8edDOqWiqm8d+NgN0fw0RPxbDZizkCeL/NyJH8K+go6vjVNl0M+jsLT
YKEfIu7XpkEh+zV9jCCYJvyYEeT7ru0HGpPKA+xTmXKySpVUPvlM+dxRAm0O2ohxywHo9sPi4Exf
GJ+4/drjzyVP9SSZDBpz+X/NvLo3ibPbIfrqspxNFApRl43WK8G0wF5/vs1O/AU0vMt67YYxhMfl
IbykGbOtp1f/6AF8EyvzSFlWPVFlrcNfc46zC21xlRKqY+lWfuywxc/3cjVZEP4mq2wYta0YQomV
hcojG4oQC9kK1F7G07IV0vQRExcemBx+cVau5BFvcSX3h0H8ekx2zYHaTT3e/jqOhdFilZ+Fv3lx
bvJZE9UKWjEWCBIpKBvre3Etd7kNRWmBHlc2yFYbfAiTvpoDlTTqFq3ILaQPZNnTdL7al3DLAxzT
PskqSmu8s94LPME3QcOa1EAel4yz2aQd7hsA8MBEnWdUrHqF4EaWIw5aO6ANJLrgJI9y7OOe5MjI
5JGjj/lae7YQ24sh2kGduo17CfkisloRxufenoP0DvU6E3CG4hpDPpNrXatcp0MRRxu8MPDbQhsm
SqSazcrzsBPb78eKNUkHHIGscQv6mgsXz2M+mWV+9Ji9D9mETaXO/NZ304Lt1Ui03H5Hx7Go9WWu
1pYMFvOynOIo3nySFNVktFW/8hCtnlxlUQXNBFeG+KVHuJxNg+7yi+lpIYXcAX9Lskc7W+bF6HjF
HoTiVocd/0kMbTyIrR9Y4cl6LE9U4PIp936EJ1XT7zUeH9cuuCBbfyHMJoRkdqUwEItGGEkgwCVp
rcA6Tmy0zK4L9fsSKMOLlyNRm+7+94N4XSjIhhvTMOxtZVEvWfHaDguqtUPoEhF00BefoNXXEEc2
Dfo+I31c8Yk5THNKvkqXO1HgvL6TfqkcnSeYQnj91PZozEaedmgb+MLlUMuLLN2SOD4HIJJ4yAXc
VWzOWtsPn5dyeV5nr+VHQeGA/TRDsGC7n7e0LNP0+FhdhsJzs5tMs3MiuCJs2aMSAON5GjrsLikv
crXLufCpzTQDnMhiGWYq73E1G4Jlc1b7LZZkZ/iiNOF4AKqIP/PTUhWgWRDoeXiGQdfBf3R9fp60
02ZLtZ/W42ULOwNw4mAzpv3pA8xBTRxO/zEkqu4vLSDST+o28LqLcnQVE7OPyk7R5y1th+M54y5e
AwzQMdKkKUaGdK7RYOVpNog2X6uW45BRmTpMSXBw/WIma6qm2ozs9kFRnoVC+xZqv4dFMjotGLMS
PyfHlUN97/N4tMEWsjHhqJipBsr9mYK/OdZv5Q7ABfti0FSovK1dRnIPx35CDsuVSpobuTfZ9ibk
CaXLi7/lYxMv7xj9AYlYzLVJgUxGeTJHlN8cPFq6oaofYveMYItKymOG3RzoYZ5a9yCLPRTTdwg7
9QsJMilNy1bq7uYcXNdcA/igx/RDAKuVMQMILW80jKpPOKDebGYpt1TuSdOyqwYsx3+7pvh2G6Rv
xiyf3xsQhF9+/ccDtyyiN27UNpY/M0jJKv11iCPQHKdzpO2lQxvm4p7CXzV3MNOilFT5kcoI93Qu
hWKEVnyYZldBmGesdebd1PDB1uIEfgHA72E91R2VR8PfDeww7+V2wxpG1+EKhWFdVcYyulYA+Loa
A5UKLHMaRtQOEvpWtVkWKNm3HGnHOtBL3ICHH0Ljk6fi/F9pUryI2cCyrMagMlOLXmvRDCCzhZGh
lBBDV6L5RBH+0yhr+NyLsZQ1IN2UJX+OICEtlZ7cejJFFdTVKCrLOCaUT6eBrHhK7Q4TxFLBGqCP
HXbUxUy8Ck0mLNXfPB9xQqBnQfL0+DR6sZKBhu1oUWtF86PB5mORQkaa3Es/eF+PPXRXPubDPXk/
bbTWTez6XF45Nl6G5phyT33JRUkKte3usT4pFY+mNFw2lX2URcEdoh1U+CKbBjmFjHuRXVkgtPEr
Yk0Lni+HPB0jSXuPMAKW4C7+OEDtdyqxAaAYPt437bbGp4Pf13YrtLLOvKU7GXhDYwKGInhRavxK
HKzCt38yX1A5/GkvnwxBvhwqYx8A5MaQCpvsl6OhV2Yh+J9hmeaKcHYKcjFDetlKaTjPSG0SRKJV
ut0gPqK+2/tWXa00xLAwMeWJKoX6XoN3PvhidZ/5NE+CoQLgDrY2x6J8KMz/oygUGuXAMJVBFuux
4RFcYwpgzpJnB0ReXSlIah5udLkw3sC9qkbcKPkCP1X3tna6tEqhudZsJQPAJ0WlfwMe0NDJKOX9
mv8+u9f1ekoXv73YYgNZtnHfyhE84wujscLEEwXT/fYXBhVI/2DEGYgUObrM1vbyBHQN//uVoCdI
AdgwV5fcSrQdfv/aT8mMMPq+n8UBPFuuAsP2Bq2YwPGYEUfgexYP9pMmTcuNcxDx3wPFdzcCjIpV
MSUTVRDuRgWH+QTw8B68Tt0Ab1xbqyTXBCwAMjQf6EDB7a1WN+rV4bgWcK4OyOPNnZoW+DUvt4ns
ct5YP6LfVKqmPuQT6C6xw28aj8NDTlLuutPJv1b5aU4ADF4Ny3yyMAwLuHhvXpQf1A5cLalK8pFa
hnUJ5yPNkp24q3iSP1WSVIIr7IatPuPcH9lh4CYeLrfDebWaiMOpL5PrhXrOV+WRVZcCaO9bkGR6
C78lCJsyiogLeglBxWPuWBLRcHFrnhJ2J+92eJjHocEHrLuY2AYF8ADKE1BRVAISOSuIbpJ54RmY
rNmr+xcUN4YqHuc/nyNTeKqDiGK6y67/oj0UE8WZ68qTxhgekCbeXoFhXNEza5MtygPOnzUW/v1r
yYi1Bs+DOYxFKwaG7Dc8alK0c5VsvTLJ8VAWvtEs+Bivt0y+TziFClynrUwpTz0+QDd3AKbz+v/R
7BdN10w4ST+tTndbjESuYXhWh2FudRtVD9qSwL2QxPwRmT5PT/Kh0KgtGlD3awbLH+AlcLPtoa27
px1v4FQ1+0YiuMq7I+jQE5t9ahu18tzU3wHF3I2T0ap1gfN1Dvn8qvZ0RtqCj9NBMCJB53vLkiUw
AE+nTaSksngYQJr0NJmFAdX8xG1PtwBGLQCpgLW6g4szCLT7BY/fzjvxdX6WPdAw0VkWbQBozkn4
Yhn/6+uLWqK1o79cPshmdby6YusOR04rcHqO9nSfWF6hGigmtIIKpP0pvEsdlvmi+mJAxjl1J35o
sX0KhRgdlEgGpMFzOsL1bUoy54cYSngLmUXwdCI/xtU3jI+h/ZKP8/1Tu5yHfPX4QZh6qedNw2KG
B1k7Mt5D61k4LQzleVzIOQXNxlJa29sij9AMH9+0isUTiCb62R2H7pUaOA/yf+dXD17vvrQOwA0l
gUnWT6eFRZ8qhQjgChlLpTFZiXiRmBPw29y9cNnKnVAVDlRAKeyNKWyuY/8NcHmyBBnufXejHxAs
4oLWx9zkWXs7J0DfZhhoJJeVp+3XX5g8pFxKgDx0s4dQSd8WXzGketXP/aY5/jYqCR0nqmoHwv8z
UUYjRvILn2bA5m8zLeh+KvDCyc09/c2UxrHI6dXd386ij+2ihE2sh5eZ1xpjfwZ1EESd0lWsYCiP
RKFEoWueZjMlI7NmrwYTmGrQnAivT1UyoLMRla1A5KpVwI1MBTruZgJ08QVD9KQQRDhx51XMu9VN
rtmkEG92AsTSFiRgPRi/abKT02MigDBGuN4VitVJLbFV/QVVjNXfD5atA8hfJ/B2fF/Nfi8tvIZ9
Asf8Yn+GcHpHyqDdvViKD1vlZeTWzFztCdZ+M1pbs4zSID0wUadud6737QzE3cL8ZxhYOW8KyiD1
8mED8GhpijCFjbF2kj5MVMGP+8lXNbAsh/YBUIKe/uJPBXGPd70Up08nbTMbQsNY/hD0oGLK8rtd
I7D8z3asd7Ic02nD09WpDmM2qRLJ3YwmjTqV7WNgkH5R5rDJYHk2yG3Mshi1s9U7EdvzQ/hsWXDE
MIeUdQXxRMVEzquB52+P47ET1M7G6Urkn93TfrUTZqAqeEXpiUICi6Ie2VlltXQKdS/OrIUT9olD
K3b5kzg9zMOq5FTiKT/ltEMS8VCBXHpY+ARGMjo99Hu7q5Kd+nY0p131O35UIel5Wih/lAfkIW2A
dFUn0z5TklXp6D06fok5s6ySRzym9sTGxj8DDaBL9j5x2TbXvHveGY7OFDrGxUxlil0A8HqnxBvS
Yct3FDDwn+IsxXzSIgurYtoeM1ytsit1EdyUfNbbgQwkECQCnlSgiwaHuBqRIPhtmpjb1ad7zwHt
CwIt/A1ey+41xQBoETx2UnpkjL1xqTFAzRTosAnD5QBHRduXz7aBmuT14/rd04kz0Cq/9iuE1NT/
VTKjqRqeL6dHJCo8yZzSRBk385h5nuhVcgxhiEM8YI0btlNGrMckeAgDT/4mV4ow8JF9abys805G
7DxAt9LsrimCOtQTpQ7jc9WNHUOcpt1a2Eknst7Wjt94Ne7qdhLxjUpUKDDN7msDyNdcUO51BD0P
sYsfdCti3cPGGXdBlDkxF01wKIQXu/HF7iBIOaalSzFhJc1O01QAbt81eff5q7HWg3Pkm5/MKTFd
9JEs/6TLtGxHei4hXSvaAvU1Zm8qc0SJZnS7PbSZ4KfcPQ3HpG7Jcfmt3KYeUWUWCnPgnMOhgmL+
3Dvb6/Aio82xnCYgKuhW8yKk7v0m82AawRzXvvNaKP23BIC6++wzbXLS2X+/v+lixkTnrmoFCp52
3nJ4/P5Ce9nQtrxW+42JL3TuOE8bh8AwBEE3G7ldSqg46BLkTsXz11xAAKF1wCK8jlaDfl6ptdpc
OB7qsZIKiqDQuWLhWw8TBhRzO+oRl4VPT0I1L9UnPf2pt3KU7nFlES6Hb1dTV0k4SbjYhuJlRLVj
g0i61VRz0RywrnABINh5I121PULPR42ZoefMBCiQxBL7DRQO+2Npqule1QFJKDG9I6C7hRvF6I2Z
euN6OP3gh9bgywT11Ttr55agvV8UWz9oxwxq2S/rpmW6GuBew6LLUwWfTnNb50hldynWuHBQZAyV
4GigU3zUBRzQFvwjlekv8vMeYUFLHHdAPzax4SDrVdszgfg33Lv04hgDuR1A21Yr8XAj7QXLN16x
0Noyge1aFRR8mfQ3l7ynWOzRZ1My4qNNigAZllHYvh6WXK+G+e5v6bC+R4W1Y/o3nd32/MIZkXBs
4Zm0W1SSOBER+gpbmkFkYbQLbjfNAyABlBrHbaivT3p+MmOuK/Ck4PpctfcRVq00OrYggRhPJoaS
YgA2rfqijn7XT3NB0yYLQ0v6u09V3wkf86i1Qbc9F8IlqSTBKx6nNK8R6b/GDGk5FkMSvpUHX9Wo
ZDmhNVaDePPbqKuWUFhf+ai5vh3jujNcyAiVdkW7E441RGRh1RvUS8FYooIxc1sqI5Mz1h6FxWnV
Jcvqyw5zF+kTqVZh3tlo8RJV8h6Oij7oqX03mdFY8XWux8iOay87ZBSFiXncX9iFQs6rDbVkEc5S
BAqaanjWWyyAcGcXw4Yp6ZMF0BL9Aq751qL3AD+8eJQJ+rnKxcCzBFiMKFac5efGdl17cDfLhP5j
Bes3fTUt3A44T40batKJ8H0ARWjMvGerZOARh17Pmd3IM0gZ2We+JIN4+8ukgJ7aB9RDLbOM3KwR
msZpFS9+IckYPB85/VEW1y2KnvGulB7V4d0WHjdDrmnmnTeclBNi/mZlfzZ/nolrWVw/p7Z4UnZ5
d6mVz3c7b+li5sJREcksAGjuOy5/o2NBqrvdFppxwJawFYjHyw5SGsa43gmwiVdrikaGlBGN3eHP
P6uO218WEJYurW45LlmgE+l2vbiXu/ccDRdlagyJeq4fmCoXpEYU9BkxTCkEMu4u2e5wVZUZtVA7
EEhMQlaUw8gJSYPizKjKTXkn/LGyt6uNCK2jqEvmuM+V5xW72SPjFDaPi8Z5JgfbvTQdmMV+381L
344eHAWSzI1R3uJnSkqq7Dsj9TMPn/Z0ilYmLU/CCXEJVowtUnhsftfKilHoYe2lnMmVcJbLuXw/
p4j4OjJMhqR9/nwEPSv47yTQxiiEcTYDwzW00HHDsx8oka8gnJlLTaeFCPPxN9wlLMkZQbwG2gff
gWdjPuGPQY/N0ID4n+vGbcTgi/nPkiFeC9otlwBqEelXHyx/cOzXqCmvVoF3ovfYjfSD3sEpJPBG
FmxdzhJkOGsmNyiQ3NMApptGfY6UKF92hn8Zke6DvQn3B4VYbDzu1A3drdWlxwn5eMeCIPA1ctNf
RpYIQtRScCMJSMUS5ZreyYgWJxISUf9ba7yWBVDhGUbmD1MoXffJQ5OAoOJGmPpgj2HUT2csazdw
Sx2jpthVYdptt+EgmCPuYFfLaxUB4IuPO38IxbovHRSsRMUDN6DuudbVz6Mqx/tyAhcIpFwGvi7N
WhRLVtURHCniegehw3Ci3NvVu87ykAuix3eaCmkV+hLBmmKTxzRG0rL2PpyIeuW1CYt6wOaCqBGL
xwh2ofGDRvibXbn/6bT5DHq9gxuRjHymaoFnr98I8rUQV6+pU+ep78bvHz7AIsGYWLx2fBzZ4DDX
OZyoIvsxcSDb1bg5SJ1umVd7gYou85VqTS5+nrUHxv/6ADi9+d+1axj2KTXIya3IVeUyz/kUoQ98
pBRYi9Ey59smYUJ61fG91ocTVm7CU90I7EWv+eBXMIWS7GutGa+E3wwE+sHfR4CFiL9XnV0RF3FG
zkqW2IbnA9kaFccEvbH7Ik8g/B6PNwDBgxVfEyHOyRjcZnrbekCwoV3ba2OcgrsWz/VSA4RdAPq2
NqexIEHUzf/I6ZFQ7gaWAyx9k2v3IRK6JbYOEDhckwFV6KFV9PKib6kDBmVI0BZIJAGxiq+Kh6Vx
r/ReP6KudrIknGbxDMAjzxWZDzmweBQHshVP0OXEFGdukCFBAYRu0hdq/KRPeatgSt9+jnvlaAGD
HaZhpjSvbPhOLqdRwyVjgn5G3x21EawcjaVASxHdFi1RmwDE/CkaWCQJmACdiPdSARAaO5lfHejT
KMUqEv52CVCbxSFynOyv00VIQFh4NhcwMGnHrWBPHmDxOjbr+L4wQ3kIZ67p
`protect end_protected
