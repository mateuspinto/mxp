`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17056)
`protect data_block
mVGmH/fT33JfQ/QFIr/LgbPDSgCoi25NPPte3CaUWPHfP0B5qwqwYTjmeCpOw2tjBnCzAxEWJ38u
JNgzMO4VmA1LZKfG3RQZJjquJjBdmkEa4sPg/4uHfLZ5m5F8R1/o2ycV0m3Xb2DmPQEaq1FprAEt
f4MjtMjl3jrYMHEY/zENr8vLGfZGqLCUz0PHJDL9SZQ7kdnEjBKrK+dKsajQUTjSDiez7z79Fd7h
ENWNyHoaksJ5iYVzfMWUINeYHiB2OzdiaQegYsma+Yfojz3wzzC4trfx2jWv2cqHYgCawfYOHlZa
It77E6Nw1+3Z7V06oWZcWeyzDN8b/D/+hjFkctu0jKJ7hVO0FIKzv1YGi7QMU2oo/dEOXIx8Ivm4
DPOAdGnK4cEjWYueXPz/2oYcK8EDxdvGlJLwASVJBHAeU0M7xXSgA0sZTdYPZSlOFetpRQbitgcX
DQnfFnCA+K/cPYGg2O96HtNBL7s7VQO9H5/ncpdXeV6R1PBz+xeam0RFF2YMlGtT2x/GEd5eKP61
UISg0fVxWGryaQjtNQZzEVRCu0/ydllN1hLrMDjuZuPieO8+YIETTKcH3IrP0FTyVxRf+fb8yH4L
s/r2kqq0SlkiN3/SxFx5fOPXtbpzkw/LD02sh7Sa2sBq3C8pcnU1MPnA8VCBQgSdNaYgGvsrNOkw
eH2PifyErMjWfQO9Zuep+RhAkUYbhcZuim4ILhjWdKJ6p/P+iX7v9gUekuWBkJrEyGjJ/tgHtQlb
6hWgnBrgLU+3kYIv9YCmBUO9LHnkvAOJ2iJDBOu5ja4NIqkNufvODHPKNh4w3G9Lsl5dIvmDq1pe
DiGPazzfUn/B3rfzoVIivPd08kJpSQM+miOOd2Mo/zaEYwa458xkeBhXqptAVwd6ra/jpwCbk3vt
6YBnxVNIp+S57w7XVIjGp7kqKreKGlYrk1DbD4uKBG5IxmMPtkNhrnuhVtFB5gmgHvQXwPrBZkiF
J7Kwqars6lENXat9H9Ue3xyF/njgSaHmuyy4bFUqnQ4IxubkFDGVvsRhW895Y9dFXLjHiT59wMMw
BSHMyAzPH8yT3ImL6dffyQT9BvQsIukQJIa9WVozbdaTVbFuwKyue/q3ppZPRlxOzuNcNZxw9VEr
MRa3KdWgstbpmNjWyawQWqE3NoFPnRkJAA8t5HpHRx/hKHOPTYEMe5WetGlBUimrSyXSZheU98LT
bngie6sfthegy9/imFbrgpIUtnvaKS48z9G00UfG7LvcPiEq5vk8qT28YNiiYDjURXYgIvp93xt0
prJF/s6Z6g1clHgLdFtnBbAK6TGjcVluf+gql7zXZ6y//i6Hsx7LJmB0W8/2DPYp43ZfYtUfGtG9
fW5gO/hARsCzN1cnXqTkPP6f7AR+PxOlhf4OLrthoJ/IRbrRFgCk2itRqPKC4vzHolLef4Y9f62c
8DSA1gyJf2P8TED7IUwcNNDtProAq+NcnfuBf3cXie2fxUspcfknL/G7VrLHN4dk7EnkX2hM9SI+
4YcusbFbHADSMHzsNmVCw7FwQdybz/J4WC8Vzu98DfNMI1CbCrakeU2noSuldsdOJqjdlzwzBQwI
f0O/+tTCmWQ5AlGWZ3wCYlB7JsfTvrg9DNkyv/5Pw4pATrh6PfA+SFX3u0OiR6O379rYtHg/2NIF
6Wy3IsvAaT7UKd7hhgPHSmz9d/RdeDWF8szbWZLvoLe1pTS6puw/qJSjsFFtRRrNE/kTkXrVCf6H
TFmL+atwieybotbEe8lor9GaeEVeY4+OepPy23mJiZuEZfoyHF7sj58GL8TY1PCL2U8vC3i91tsr
V8e5lylTuRsKaJ9x2GCHC4BsjWeDnkyexYL9XJN+tUaesSv7wEWslCmiYGUk2URYHPixQFSj3Ag7
ioImGBRF9D+fBHb56glE6NvrTyu9ZS/SYtgTKjw50yN24VJA7kPjqLue2RWzC9yKGbtrvG5NJ83f
JpK7s3WYDEyHf4FzD9+vJPM3Uduf93tuf5aCsdcwLFeVtZSVtznKLG+yGtFsIcRFauUfwlk71zPs
l8bLuwFJgzN5gMfZebayR4pnimj0tV3KGgk0kijQsfBSEjyh9x+iOABCPkVqcwhxesjCGLwnJLfm
WvUKgnyqAxhCGeBgdqoxr2l4TZekX1gIdLTbWExgseJubwXQnZp7F6gN0+z5wfdabCvFOd5v8tFQ
N5WDvFLkD9fdtnUDD4aOXdZRNEo/eMchCxpYfUCzppcjxpuBTqvvl5h012IEvZUryaiNFZiq8J4S
9prAi8Kezyhb/WJjUxQbaQQsyxgSPSfHBmxYayvfUi/Y1pQL3dIB4NWQKqE1xf89X1K1WOddTuot
XS0vnDPRSW6J9bIiovZf89Q6+fpWV3YXvv5cGrjcav9uOhB58oy9WLop06kUYSaqmRYQJQYbjAm3
38X04ECSrJpb7cgW6CYxE65zZV/t4pSNEETWDo/26CU14Opa3tQ6za9Fw233QlTunWW+erFbqQTD
3Lw2l0DsXl42KreMK8FmeN5mnDR2jHBj9SKFKKE83hTOM+SA/QfRrInb/fhXD4I8+VB7sK/ka+7M
mc+YB59GzjLp1SbHBKBOjBvxqm3SElBReTS2+2fWnkzFWxAbhEvG7z9WKJgipeduMdV8zo0X59lk
AFhdISQm1gyQDsNt4SY8+KOJKwMgBQMbgr4N92cUcuHOcY5hbyFa94GohWNHmTiCvAdeqJlQiXCR
PniBmZQNrBYSUHAiRky4K78SIyu6L9EPX6RIPzscbMSMj6Jx+lTFv87LxfaRtEAJJEPKEFdf+O2S
f+varMLCIDAKo/KnoaPBZQ7xMSs/nf+6N+1o/vamGIUJaUGDWXJH0KZ391YjJf+xUwOQpLePf0YD
dBvSj3XnzQHXVNpS5jsf5FNCvBkCSEZ3/Sqj45M07L6p/+TxbdVRmT+CFqdtFQ9H9NoRDRhj/eG+
S/T6TajhfzYohUmOv7UJOZnBEFu6H9Edg6vXnP/Aaf3hTkTwJVO/jYVO62+QlEL0+9EM4dnVc/bI
OEjbZbEzUGZEvGY9XyAlADyQm+zdHqTgX839KQdKet0ZArG5P45nuIZckFgl6TWQTy+clrA0IstG
eViRYpLQS5W4zX/E+9sxJeR/SOOYB8Qn3ZiKmSoxoJzorSHGOZXMY7yifN2MPxB+f8kZDF+z+Fxo
l/gER16vIS0p+ghlbW8uVlv99zzhtAhgqmtxqxAXI4JLh2OLXDbE4pPqBiBA+Cdv8z7z/5jQqb50
PSVlkO5QdHDHUtgrCbR29gm6cISqGiW1mslA00YzaXYKjQnFWziYjg3zTTlqxorZJ7acKXGANkru
LPYmogNm9gEQvIqgasUgAENMjev2yPZp+sD6fC+P7/hWgwy7X4evnfAfxP5yFM6kKyfevH9LZsxo
sOI10Wwcxy32bQBMKsDDrs6e+lph3EvLtR6dbOYyjYVcZr+LHauY1OWS6PrGrS9Ah3DmOmwiikR1
KjLI6fIjTnNb+Lv9TrmWqSjvRjZBZNZ/cbqoUwF433RNXyJqlKeXlIzf3tO7O4CABWG5uc6e1/gu
qSZAfppmsGREHEYYBNCANS2trlsM89ZFGvW0GmNQOqYLDTOWvvDX7yyEjLlGTyxTBe/0Usgn0bN7
bia0aVWPkjsfIiDAY6s+jn/7gnCNkb5wx8a1gOLyeih56zgt3LQide3naqfCItaM7WAPuB2wIR6e
X1cV/bSBdYHObyAtSwhfwC+oO9eafo+G8lL5P8tKszf0derufRrOcHAD/p2CK88OlodcaqsQFA5n
bzVIQNot4l+dUTchskyKxUhl1uiS+Kw59+CTdATZZihs6UyDvSGT7h4JxKDXqyGLewPwH16mw/2y
n+8ym8sbKrssdKCwW3z+VcfdufQOiiLl+IFxmRsFokdVmgoT+AIZMoSA6zHFPxIDALPphAnWsa7O
FFpa/PUq/pnxrY03CkSPdOcJoivH5vfN8PmMcvypxvgXDSCObKP4F7L3VJbm9iW6f9X8r2oVNLlZ
DtKGX04hjFPM2K88UwK/a5l1fC1g8XlqW8On/s9Z5DQ1J3aUQIoa6DA1beFO5ems5WMEtx13DrvR
tg8e2p3UkvxqbxJWH1l3TfYVB6xboNSPITb5z/ZTNJVgo4Xn3MLawJK5fA/3ciBrSj5pkY3F/lhL
VU0YTIUhdlZYwITinDX9mKG7omB78elFkK8Bg2JtVYXEWUiszZhEXiGFYjPdaiQ4fk7M0A/fQZHU
nMcOd/XRO/kYb1sZA84SAbko/bsSzLhuLJV1Gc8S7RRk3uw3j1xdBetH9SfG2p/ehfWhqyqC0N0m
Mzjt+jENpc9v96l2qapRPSqf52ZSnpOrNwupB5kvyxmM2YwRPto+sbfkTVv+8135NN9K2pJFSUW+
0sv+iLjsLIatKEhGAoudZvZA82+4Jt0QnO3b3+85spDXIrBSZetPoQmh8+pXT6ylJuaAKpcZ5e4A
KTLTI6NME7iDJgdgf84GYqUfmTUbEwlJEr6aLSs67891JXnhgEAsrloBOuO4wOjieFT+BCDUtJxS
JYe2w4ONyb5qL4+sZnt+xcMMiFeoHf1lyFMYXgZLddr0gyYgBuT3vkcT2AS50giF+EHQcZWBH5+E
zMtcDawQqwy+0nhppguu5roesrFy8KgI0t0WJ7YoOr5CPqEsb0MDZDGCKiumAWkwcrDBUaUjv7m3
uVJgOuvHi7UYmUBcKMRaMK52vV4A1ts3iGfB/s93UrpVvnYs+458BQm8AhJsUV6T2bWErODA8jBq
CO2uMZxtsr7b6iNq0Js05Nqmg/CBYLhWanIl85eBCr+cL7GeNyXJTjvNNmMEUDo7wpPdQSA9AvH2
jIzjOwEzpKxUWyYJY1zZUypxdPr4AwbHmnQq7mXA9iEYULR9fY5UOhweknl3nrqnYre/4HYI9gIb
SgqlGdf6p3sdQTSdfzZudIcvinwLLHmifIrih4lRcS5H6qPpMT9Kx19D5rVIucHN4DFlyohZUG1P
wA+yLPgjIAU+no/LFfEtUgXpgCcu3F5c96zfLcmUHfS4Mcw6i0MarjjVyshHJqlfIKKVqIY7dmkS
X/hcfIzDtqERqopo9RypBDTaCRPqGS7xDSyz/xuyMhKimaKGbNUaFfJNlqKJ+tas8jp8jCVyAezE
BjDDv5fbaKKWGtn3+8B6ErNLMH/pD4KW0+I1BmxfYbccpmzXglvRUX0nNZMCkDe6oDL2jWrOOJo4
3VG/dZkFe+MmDTdFSW3wi5CZyDvmiSCp0NPO9JlSHqVF9wCrZyvb3bjwqcFz0bQ+v7VkTwi5n+66
QRrWI/ersR0rfLdoFtq4qO8Ut0uBFz1XsmQs/XgdR9KeEuyiAwpQ/R8UENZrUZjDjJP8hRTBwwE5
h8zn/wU/00M1qGq5ly0vh6TxVHf3GRtsAauWCOkaFW7+ZyW8uKen3C3FGcr3uDFYrKNhOEAlieCr
BMQO8CsX0jIZGdCNsJa34If9rJoaXIMucrv/iiR/HunfcmM+q82XNAfBrsvZFs5mMTEM1eRxMgu8
X/VB4unb0jAXBx/lni4JYG/4jIRJBLmPxRDpaV91QPGa5yMY4DOZ2az6IhSDol8Oob7UTCEUJ8ge
0807udEw+/ogx6sCo73oJwkxzjQNTIgEy6yIilXYM+pg5kJDVqwV23vcz2TSyYjXQmjNcLeqEjP0
tnKUAXhywYrWkT6mjDhmkyM2J44rBhxUe6NfyB9xvHRUt4co7dazVSskyVJ3KgOJ3bZXCJ44UWZR
4v80Ck+EqLkqanpi323X/wcqYm6vPoUXKt/OcmrH4MpUQCuOESZkNNi6Sx7FxdltX8BmMpj9iDDu
zspEr1EFtLDoUkC/134QGpmE7MRew60BBxHE679CBBQTxIpJk6YAcP0p6+JitYvUW5/+I1M5VuHw
z0bW4q2JwV4nYIIoW4Uby+qojpKJ/v/gqLPndUJ9v7lmHC8LSxXt6MI0hfoKCNmjKdpHwp1gt8+Y
PLG10SRgUP7jdQ8Xu06guGHwtPaIeGcxm/rgNj+bk8JrcLDRN7S+TmORzXeds5Ji5EQjaO6t6W3s
h1jU0gtWMH4o80CTYifAUcA2PohcJ9t+FOQH4CZ6UT97rAZGEgOiILcmoNjsLDu+04Nwq/p4ajTT
UEq6ZRHoyeWMKNOPd96oaNhxMuKObUXlECYEjS3RdgozYEG5iP61AJ//DQBDCXXZHYUG7gw+R2Hc
yRS+v8X/U+3so/pUnhrx7Xa3KJZuQTP02+Ma4b21CTdcEynK87sqyoZnanpwrUufWkHAt/e5PaKf
B/cgbhY/OUwQfGr7L/8K4JT7QE1zTbEYeKyflMV6nH2SBHNeqk5R0wuJlCFPQxu2VDG7oJEx9ISl
0dOQ1Ks/vb4GhK5wLrNpKGVWib7FkWlOZBNVcUo8an1lxhAewUPtKvacrbMFhfLPjONkPP1Jed7F
b7GDztTbWWMCY9BwqMAi7QCKTdVtFH/RRGVG+Im9EN4nvVzsYIJuHq7inIhDnDZ8gjTkE2tNIX36
5Qww5crBuKsyZYI73AqDKra/HJazHCGupUIB0hsDpy6aYMV66NEb4BQqPwTF4aNDg+i0k9psR/On
zOItTXy55VMC6+I1gRVU4BN8h0FImjG1WsKMR5t7lOpoJQlBYaRChcg92zKp4j48p75XGmQthfBw
3b5Xzpze98e7vFEa6il4EaMM5ST7Qbjv/Z9G1rbAa1jfDPhLZgYln+vLE289km7b403JAbHO7MQY
dyi0ouToLeuV855d/FTCTPNOcSnAeLgpalpSuojVEfcDyiJUId1Pajj/BTmQcZz8duriCiQIvgQI
U7Gj+5byXp4NeU/ktas24mhDf76QVSMedQRN7WLu4nJGsc4x4T48Vnr6VBAXAbno0VG49sQjijcD
Kk1t0EkyLqKNr4S4uAujO/6ZGxg9MuZeQz+AMfW6LoE+FLStd+8QbTzSmjAusF33p897vI4fSQZD
lydwhDkPNNj3F9iTMKdSZiPxXliQpw4pIuZT1/sbJ7tv4Ve19nmBleXnTocGMLTO24RnjTYZ9ZAC
uzfbwyL+hlJZp51L8U6/MRj0jESP2BNVov8GQeyAwERnbSJCpxb88oVI+eJh9WmbgebrlmHULlXz
UhkAO6J8fF5XT9obUAlanqCte8kJ0PyFHESqdtqctbD2Ne/JtV3pPkpZIPtchgRtd/3UmPJ4JV69
Sd7b5SeYmDdGjPuHx536W80/b1UM6NOytcVllisan6Txp1+zVSL0JPUEVOe9xfF+pvNXvA2Ix5Y7
8wqEmf7b+a3vdcg6bgiaEkkS5vCOa1DUSqjX9ipSQSgeTiRNGQ3gIDC5Ob+MyX9WntyLU8GQdeYm
8xLl1oA/e7wq7v5smef1VatPnV+bJ+UIz+C1Lmcd5ZL99PhC6jKHg0qB3BxRmPFfqP3wMyKIgLdI
dXYoyCmAFDnRFyKE/BwclaNEjwYjQED5TAHwHw10sYDae8Ddqa/VGukATLjGKnIn0d7OxLcPdBOL
srzYfUkvxBHpuoEGo1++dGKN/mhNHMb2InQm9WrpZKGTcurQesfzreXT9H2JLnnRqt14g5Zu1qAO
eERfho0wisVgejfvfpMmbCt+9rahNkbWv5BmUKdiytEODzEUm+yO0aTs8eZGWtiWtkapqM+4z7Xl
/59XRFPGGQIGF9NXyEUG5LeCNBpQuYsL1ikAqtfo2DNtJcyz4eA1z6min4UZrykmCXOTL7p+kTka
ZbN5vtDJ9UnX7cxmfOVbnih/LLn8ggXL45FQ6AFJXFMo/iLMcia3CavJSsmoLlmJPx484cc/q0kO
8aWObzz7huynTmqP50NYX23BhaD+aR0zZWV4OZmfrDYtqyIAOg1dkwhObcSgUqv7y6CPqhRfOPPn
9okmAZehyIgC7iSNDfmjFOjKHn93qldRLZu/vaAjPqxcg8V79WHY0kmrcsWsESqabKLxyX8mX97R
iMpuv0Xl/PdGwfiXHnxhkuYPRRRJekX+UyKlWHAJMXZ01mkCLtx8x3SSdPHal9ndQv35D+GPk1f4
JLjSX6urEbOipN2L50wR769zsZ2ueKBvZbyE4ffxYPtj+7zc+EWzk5s8U7M2T1mhj9luo+ocJ66y
k0CBYUYE53EmjJ9uMwvGcC1bdwOD5DWBuh0UYJ9pqNgdXo41pLCBZu74zIaH46TDe+WyMUCEwblv
q20sFTC5FMgwX1+fnpznGPYpj26XHpqC4DCtl9hyacty8eKn1KDj5DBKxnawxdllfmPNGCJVUDit
GYAtFxD2k9N0hZ+UCXohrxTPPso/GGgKGfvcy2vpOz/8PWWnTo/tPLl2hwylCZLsNRyXW/PnirsT
la0nzCCvay42qjDFltZzNbYBH7suCN7rbr4+L8sgu3hhkKUo1b5A0RQIQTiqrE7ffvvbG8a90/0g
OzsE9uXTbXE8LGRgj5L+L10NQFgV1zQ+0b3sknrLUuxFti7uEGGYBhR0NnBcUWA1xfXeVl3Cs9n6
u8mEZBUU0EXoJfSWMJl9YR74luxBYZ2KbT5fPM6sD0CSJAOcmFn0c3tgfMmYIE9QH7zW1VyTXtL/
OliMuhFomByOQE/TmeguYetdPIuUPK63K3htxTnsmngmfb+N1/15Cc3OPGX0VZEEiu5LU1N6lmuP
3JYpxLo4G7q0+8f8ib2TCTPd+6tsZXOYaPEz4QQZWets+//TFq22Ru5E7FoFN3+SJ2ywF9f5lZ1C
4YJ60ElNJgVtav0KJ2oPU2ArrkrF9vAZZEQ+d3TDmj1gYN6im5RdZfS3zIgSaghcuuRLGlASrKEQ
Kaa6ba8zll0bIxA4H/hooBKy3W56aPXRfOZnzVLGK+SdhkzfWYEDbCON3Q3NMQHfAcqBB/hvHHQC
gVX4pGSjrelc75Ro+fmv681KQisNFjEWeKaAe413p2kZzhKmUplIuovlIcvUGtUOJBxAETKSIs6+
VDtw7H/bObGi/nx2poDomD2lHwHyXWyt553tez+3HnEWNAMs6YxmIoOkZR3brlCMfMfWw1azLp/E
HIFz1t7Mzc8zDmhMkQuIuu5ZwRx9CZYLUEEb3+mR0OqzKVM8gKcWu1k0Thjs6l5EcO357ItgaXvI
rfsWwLTkboizky/A4zSBNyHR2JITGc9nRtiBRcsupsOg4lLEo6IbLYLm9Q6o5EWgjukHbTBGPu6G
UL25DsCXvmXObwOo9LAy0WcvTBMr+IBj9Tr/0U07yKF1hmUBahWLBVJqteGLD0a6ccZS0HdRcCkI
0ew5ho22wOlFPChuEsUByXQGU3hKA/tei+8dG/a7KghtGhrzMM7+QZdWUDPsMMvAukFE8ZNmN2kN
R38COZGPTlC3pNIOEFyS+P9Ei8KHAU3lsLhkAqsZH7odGfXvBgud7ClwmEplhgcMRk2lhh4eKNLZ
ISTVZivQpNrZdDdBs2//J3EdCBkGJzxYginRhuEeRvq+JNANAVF7Y4XPKmEXIXqy/Ij8RDl9a0yV
oucbs7K5n5p+3nuW49HNCpPi07WchFe+Odcdb8/DVs90VA3vTShNgWczDilX6vtHxR2smFBL6MwM
Z1q580hzTPVlZqVAFDpu85y1hg6igp+j8ujoeE2cweRW1vdvrSCyFn+AYr5D00PyjteLmcPAS6tn
amTmuKWqh2BHQSAgJWINo5afHDOMUE9qmVD4a9jKNBJwqrUO2VmH177piFYnPVHSIEmV+5+L9oG2
HKvdak+PfTkuqmvrG1N31reMgc1u5gW/vNt3QwcX4BOIckHUxDLqrmvXjDWCafREZkqGBwqyj0ew
o64TfurOAnVoke091cK1PVRRvfbLbdBhEyVwUKXDcCA81RuI9ic9D7EhRIbWS/liZK2/A9hesHbm
2QJO3BMrdruDjGLkDN/scl7Q/UaSm65iKivW5HRrPXwNBj2Fzo9UOabDh13WM+VEsq5yJtEi4P8t
PV7nggRk0o5FcxJ7tlijU0EWj2YF/R0GANxFjPo+tdHqdtV+k69RMXNTjC2XE/7q+pecpcX+dxgf
mlEaiAW++SjdzvBHe8APbWDLAvGIPch0FCF4vPseVa6AnjwnIpdjHfWz4dUqyrix8SWtLW/P3fpU
OCh12Jzc9mN7zUX36kySLhx8ZpGzsbPZf3sFpna3unTjSDPXEylGyr1gsZrB23mrJChMIu+7e1V/
Ido+ofXKfWXF+jS4YJqxpSMmHzMND8r5NuS2iWIpaxziBQ21yb1xIyEU5DRgZi6lUmcRe/M4vUj+
AMiXfVSD5S77PGoariRhu1kln7tjEELg5oq+nN3DoF5Azcg4+sjH+gUxS702b9fpVR5gcrC6ZG/d
x0X2hhxwt+LSh7wLcVOmycyllhFh0FnPzBbrYukeSSEAO+fBIgpuLHXAm+XNQL4e+xST1TRvCJRC
TaLZw2wcg0Kye034Voi6hEfmQ8igxnYjxyOt+6h36Y6iMQ8ISuFKJsW1PRjEiF8sjmzOSPsZp3tG
vtWPndX27Icn51W6/sXRQipGW3kGyfEyHSI9WDZ6ckPdVt0BVBpe9aqUlDKy/aLjo6QA3jDKqIHw
Ni41HkmtgOQbCbB1flaKTMSzTsJO8XPbvixuqU3UpIDgjMpLKOke8iz27Y6hzI3aBz3ascwjipH9
ClnuxyWCcr6NeW02ZdPnUCAfOFOC9V4moLPUJzDH/C0WG1h+t4pttqe1HD41dVEbNeZMZgW24BGt
TsfdbAtNXSdd9hLitG2uJEFw5GzZH+Mag8frkrEjJECh0kOIbdIydT/oGX2yDpB2/JqO5b8szdCY
q7Cc9c+nojJULOPLYIL3sHgvCnoSXMSf7DFSpQXFA6VF5x5Zs/ksi2hdOkXIR2/5+eZebxm9DuCG
45xOZKvJFwx88htQDnX92G5M/llvy1iOzqFrlbXRe/q/A3VVyO3umKMzh+Lw9o0mh6o5fYUgLrpn
aLqNYmCcf0hahak9N+30KNbh7YM2O3LS9BVuyhDXLLXqgaHuOAF7BBe1TeB2WDD9lUj4kqg1hmYk
jzYT169UDI1iSeIXJPP1lUUVbpilG+XzfEkpvogcz7AzRt6y8d46nHtKsXGZCtmWXZIB2YoBEvQk
ifxRaWVQ1QS8nfDExQ7aRUIeNT7EZqu58eBuYmg7PoYN9wdehRygn8VHsC9451VXU1vfTART04d4
emjDW9irtVph2V9GTUWSB4bLUFbqi35bhOV8q0hiHePmSfaPz7xrKv7HqRuXL4kJPhfsd8GnUz0c
42NUH4Q3Ne3dp3Gc1jrz588QeK9Ej0LbnJrkJymJ/aHrQ6mMPct4Ikq1A8NszvUIKygaIqrTNTS2
At3aZM8Qt9Sg0G77r3TarG2fmDUlWVxcDe77uVna944OFNO20lGEhbK04fNTuXORvnfiOWeoDhK/
memXk71liePUjVE9Q1/fyWIH+ydi9IdoRtmumUBSRHHqaY+0dHFSUnGnw3K2Zby35C4nfe1Vequa
XpHPb8p4KN8OZyQyJDQjZqx4lrx1oep9qaAW+wEUSQ/1//isvkUQtJ6uxv0yMS/+TmL+lNZ83MRb
aiiLd34UtrmxGmtClNs4mnC/mscGFAQZUQwnZ4rP8ZCEuLKpx5f2bHelNBRdPalAPBEhkUvwB4to
wYOLPqsJgZIpZsUWWNgic3I+3a5rBbXHpXUMELjRY0Z0qIvdUhc/D6+VAAuNkswlC7QBkagaxppd
b+Coa5O3YOLImDx0ifUJYouFZ8XSxBK5wGwgt0fdZTxUfAzlLz0/jZzOVCcLp2SoRYHjxSMmnn+L
gLHP9UzC6+u1efTg/At7Qcsd/tYDt3UDauRZ+j3LLpsmJLwubUvkxIEgUbfSrx3v+tram21oWGZh
tZL1WsmOhA8wB/UJmYQWdt1ag8FwN+6+oPcfPI/+xgiRK1xh/BKxNc2b4/f1gZ0UNy/8ar4PU6sc
unrzJHOxFvzcwL50nI8n2FkcXOlGLhstFUssuJ0rXYwViPdxZn3FsQGg4RWbMTwsoKfPRWmIBnyj
SRwoteqRgDuoJI0QHzfkOVXKaSSvZBtTeW5E071OpESSI5A8h2lkhdTKNi/jqmtgSCfPGTtAf6oO
cd6BaaqIXsKyZXxiKTfZxqPkapEzfvharRvp6MgVIADGa9oVmaR/EGnATJA4IgByeAaJSYv0Ln3k
T8g3JQKB+3qdOeuNyXIgeQrmelHAk9EendXlAdMMWHCH8dHYPogMBHFlD3drEpwGfnO3f0VWMzRX
MTWtRUAKJKUzLKmDXb8FgyneC9PrlXihEzo7xZOVeOHxKKnVT9ocMVxCHhqoGHlaBD/0wVWDOy5b
KwEfvwI6Rbiztxy3tpdPnj/zrmhUsPylI85P+aS88w8FQgPynpWiPjwYgKmjMhhNX00/5zaIoLd3
4crdCLkmaXU7ptfBefVLR3xPCHZvzNi+hf66Zm5+pZu/8GlbhI9ThdEzuPqIfscEAMwcvp7GCfJ5
82TBZzJ0NMUNsf7nSKjjl5ITR9XgCEGxCziC4ahU0VBJ6pdhNjUacKuqkdRITpM8SpHBpTtQ2Mhy
+6HtTkh7QKvpbODtAZXmUud1OnXObiEry9IKLni0vdL48J6YQ5/eeJk3bep3INSu+mC35C0K/PKi
K9jfMqgsZWOuM6UUYQzoQ8ud7qzKlH5ZlrQu4EuhhcsDOR1WNkhefUw3NFDt9M8yj1ydUXV97atC
PdRQmmQqugORXC8owjteoamezreVSacnoA5lsiNiLtZ1z/Ei5gbVYTollDA58vvSvjzmGNtM9chF
MSy/kOCDzaigCaxSJ3fCSjBtE1HtW9I6cppFI2GlX8+MH1rnqrkQeKnmBms36A3FWkLZGsbYspnl
I8gdCnghmP30Hxsi0AZp9fi6HTaYCzSSWF910HEKmCS+lDfey4j7wiFQAQ2TabA7XUu1ltCn+hYL
JndO5Nz2uABzzSJbYGtCyE3DtHPkiTtU72dmwN6/bR13ZUGPcA9SU4uq+Vwl/PwhrswT6v0FMxlk
SIVoi7g2G/ESy2CaWaYgyvllLY/xknG2YMYAlreNeLSkVaJHhgOMoznMxdUoCqZ/H4oFltUfiYAd
9LBA1cIj2jlWsRIPCwPmeYIjivWcNYvdRfCbn2WCl6qsPz4GXMrawBRYJwC5KDQlf6v6S6wU1BfK
WiJyFbNfDNK4El15pY7N9tHL1q0ZZMvr/PTiZI3VewYObQN/Pqfdw1N54prf0OtCxgZH3ZS48a/9
9Vd7I/6mo1x/fiAi/JMxkNqiC2MjH5F/9ugViaWkNDuFUgGUz8XhYvyrQeK2AgcccE+zJu5c6c+c
FG2DgFN855W/1fzweVz418C2pZ2QGXSP++JKv2GiYrjtzaeGD3/mftPn6UL5iP6xwJ+wEAlhgV+r
PLUV+08nD5CaPzAA5aIXrV8H4isfft8myR8fUqpWUuN2ntw4h9ADKpkLr1s6rTMJBtVCuVd2x7oI
AIjatLL5a0gxqC0CwJVJW6ck0Wqz4r7xDnQLYNIcpr6T5PQfi3hbsuImwCrYJ5b0WFbDS8/mP6PU
V+G91xIfYSfLluBEPfm/VwPA4RpLv+KDo+Whum+s2V0SnqAgL/2Cbuefl7RcNnCKZu8ZfgDCmzWL
aDz4GyNBRlqcFOiD5+JFOLtDyc3vkW0DUTN+8ON9RyDUkx3crxFHVXsWAFVLyKr1KzJjprbkchX6
ZutnNc9XY2C7lyjTrA/e3GxnHaBNzNTX8gfgm1j1D+IPTfQPwxwrIa6c+R1likLE5enDRwsoZEW7
74A8BGoAfaR5k1R4MFE7gikOh21KVnJxWshXFDiUZ1UFZ/Wvn5rCswA+8JlcAvswZkZN3tmO4BTU
V/nlzxlSQbFG2HYaBWi8ML4/sQhAxurIBjhbHcSGRfPvUpip1riEJZgVFghS0kcfN+1Ega1TD7ye
k4lymlizDNXiRI4OqR3Sp4F0umK9MsQKB+LdyuGgS7LuJYPrJEXDVuXjMbmJmiQKBQUuifxU21rQ
3r65DjE6g+gkdpJ+BemlhRzinaybMBs5cTHo/utkl7M4s5ZY1AZEexgtQT/cMD3m3fOfFrigupqw
5df7FzfacvHq4BVwC4OujA/6LNiY2GJ9UJH+q+ThOCNPnP30AoK7tkeYbW9+41GVj1EW28XKN7kf
epTwKc3yOjU12BFy95YeeDHiYU8ABu3v42Wb5JEGvOb8g+yrAMF+McQlvnHjZ6WmO8WEtXyJb5F1
3GkVUeBNn4+xK64TsUBg0pnkSTFq6P+iN62D4CqxNvpBrtsyFhfbrwr7c4/7z69YF2OZTB5NH71i
QZIA3QC8AANlKOg7DW71K46mp5XDP8y7atDGpWGA7wi5ILa+hzYL0Q71Gs7szCFVsKouObZ8zms3
rfHV7qSfI0/88g5pGe4CbEzj8LzTYZ+OGSx1HToJbsPnNxlasaIue3OSPM/OCnQnw2vy/ZBQId/w
e68vByazerCM5fzZD1R6lGfDrGQriULG0DSZUQCFcwKQgx8M0cfLt2h2FlpiPuuac6AjT8cK/6TW
tuMR4/gouH8W2igHa0FLxAr/Nd/s2kKYUyF+vaP1UlB6JthE0CdnRujrl99j7JHqQlSL0sM6jDrF
Q4PMVhZt1p+RLfI87eclJQIXZvW1vPz2fb2/npqAWNdMvvvEPHLPTaLnGc0Gwd3yn8HSpjTHBTrt
13SefHImL2jDjvrDYmpsqw6TBxnv1Wysl1n9eu9NNK9YcojSlKpEwKi1RMM9t2zUiLqaK7jw7PPj
ghd8dvG41g18/dd8O90l7DfKQu9kc/efDcBPOi0BhQu/BILTUC2lOKM577+fNCHRQ3RpQpk/p5Jt
E/P3BXaRl3iv8ls2TJ32lLIovOBdHNoLwwFTK8O6wPhkva1//2mAKx1bl52YXySZmdYGpHnfNczk
gfAZJAPHXv4nM9d4oczn3lSxqag4An4xpuJDjMUMKg/H257lPJXfHB+08zgZCtRFClkx6qaThDjb
uvisC0I9Loa+aVImyBVJxH5FnUj4waVkUnWcG2R49E2E23NksqMwgYN63hE9A3V6//Gnmfmx6dLc
eV6EyHbvTjtWh3x523S5yKSB/1nazF/usO8c0n+AP2rfLtcN7rETDrUVhDxPYK27UzDAuCKiEm/8
DZrOzdcYzHnDJyQLXngSv1HW0DocVJTHRINbqZTZrbcuah+fDYHY6zhJscXmS3IdkcNzolOXwzh3
lZU04mX5tSzUma2O3FGRZ4BmANUvg+9DVdyFtI08lh0/2V9/Oxe4/CzIS/Dv0qF4DLDIkvSSTlfq
GhGhHpPPdDJsG09LWp8KWqooU+dJtjgoBu4BDsRGwzA0QvIOR92/rw+3jU0wFoZy5JknZVO9PFap
YgtgVlt59YChPXQ72luTQBonCjj+jeXqgHl8qHSw87V3/DbuFLRRBZt/zApHyeRYMuwx1dGAVKTv
lH9BZqoXKGjKBUeDEGOiRFUnDTKKBfhs+VNSeVCchQJu7g2CTAJVeYz+3vJt5qSVqxr03ogITsZT
pszqMGNoJ4cJu1tC2uif4b9Ye8r2+MTwvr0tbcJQNrbPVV7YCloRYUTS6ZGtdTJmuS4FY3lUP0B6
jwl1CgAuuWF2dfcN70xBJrncKTpU5qKqeE9if6tBdhoD4vAVy9tCJDcKFlE/vmLyAkcSy0qZRiPZ
gueQxSGaAeg6PjPuANPvp9Ci8JfHSXZqZ1O89yNcNSJJEEDNow2nY2da6+dp1tegUPFsWfAFKRlD
wquu2g16PFk3hbHVi3JcBEIUurbBZSe9L9LpXU8dLjthD/yNCU2Kzo2jdMD2Ujq6kAoWRlW/e8Kl
RSo/0UT6Q32PZZzew9ZgarkKfC84LtRd7HDoOLPDULGuO/nVK4ZEJnAnl0Ao44//7Ws1t0Nh6sUN
cI4/6fvVsyQmYJrfNlAyloevz3wN0O+kNAZ8GjEPGx/eA7IBCuJKe9q3B5i6qmGtCkOMrEDUaJe0
vKNTHK0lMt4yT4VTyDvn5BnVuU00i3YyNggIW+Zt3PgCobdIilF7QF7tkaFljeXok3YoyVaTBIYV
mXhSBd+AwjEBioSQz4/Utr9Vndi19Jv3vY/H5Nda5JfHl8BpjNaCQdLftUqeGCx+JP46d1qYz9Nf
PNxpjUxck+uIWoyV1AcOUdlQrFfh7qWVpuO0A7bTJiiqTwJgET8//OtgkUM2Ez0reNySu86AUbY+
9HJ8BXIW5PSfAz9gvSnAQfDnhYgbllKPHwszmmywS6Oa2M+U/XPQGyEzZiVGvRH1kHzuY4Q7koh7
W2FUYvb9miLUaNr2PtkN7Naj5iYk+UhF+CIL4dukxBDFG4fs4dplK5sScHAIQCmmOkbilGp1rDgt
tdt0cKPrvXOc1bx8Wr8gx7rKFtumv9V2eUvFYFFEZDelFGQUKco7sn4yIvX0uaLrT8czAN86iH7O
nOUNZv/jlbadOgvK9o2YUQOJOzHKX6xiBIoG19qOowEV0ZRM6eQqOOusQjUHoKfdoGDxEkIW0wV1
yfotSye8crPFUBMrIXdUgnv9et/pU8EGBr/0a+7ziFJzpjJKi9yRM3mJPLg6UOwj/JG4idhyAfVR
lYoZVmPsHe6Ok7H06xgHAxYIKi75VaT2uj979NZ/khSrm9Fsj4WUJR11LMN0LiReoLAwlPSm7jHN
9FbdvxjnwD07nBlRnvM2ixJvE7S8gB6GSrHGecok5JgXY39xyuq23MzesQ/GHepLvAdOXvHbd43L
rQJ9/Kcz6c/6zbX2fB5ddnRb+zTZV0CmCPqJWL6AnHcxrCJLIZydslFUYgIuVdqqrZTKXHAmBsOb
B92SgHiiRF3OKKPko8/8qsRxrLKZY+A7lB3maLVKh+jAAjEADgpOkSHRx1s65h13B7D2CuRQz+MC
d40tpaY564Iw05bu8INU62Om1eyCMf8712DVCYLkyFDxK2kSc374NDnSjhcmc8t4z2jSP6+CUuH+
CSRHDoK02gWnOsS3xHbwbHOZMurlArUy18NSCxc4+FUoF1jKAv/9JLG52rR9gARHRek+HDnXN37v
u9z1lRQ7OBjJpKNFKmtoEph2lkrjabVqY+rc7VIzrnt6BPE1ZUr9M+TMP7OJm1bqz1sfaiRAQmT3
Gaa6zxu8bC+MsymMysSIjfFpWWXC/nBm6T2qYiNJa4FfRy2AnAPkOA6zKc5co7w6bZS2rr3S/BMT
/CRJrnHjAzRx3EGSAN85Zzp2IyGOf8R6BXxcUrsEwvayRupqTl8xRUi3LNHZmk2qObiI7o8jdlGr
jnlYC0T0nxDNYaqiRuVKNG9pNCREE9l/lxvl2x3AI2r/lqeWER+4hkubntwYF6lCunvOzxk5/S7P
i+Vi6Fd6s4AP8BQ9HLJfjs0IahFne2AMPTafu+k2Rl3RJZdodyEJXQZmrEjWLo577COlJ+npxBss
E75AJsYUXbZHCmuUVd7QZLVOnRPmdigfn2iBzGhmbQKkljqZMJIahAtdbMUb1SDAGCb1dKWS1KcP
kKSWKsd7czVWwFzxpr2a+SOZO230wFdApcMHq8VKBG+GquFU4l4hT0y6Vq5CJKKCxGxkZynzH0w2
awG5/2MCnN8ngaFJlmIsCtI1cu4G9r/hh+j+vTWjGpwbaMKbruqcTSsx7pY2Mm460atrS2MsUJyU
sgodM/+SD50NBzhkunUHTn2ERnvFWKmDDIStSAbph1qbYdZo1iJkXCfzdm+VlB/WE/E+fCNsq6mF
x1cfgR/gBySjilgALVjqGOywifbNlkD1G0+piMJTCw36Yb3b0eRwKq+V73CXN/KcWtTBqdiODyGb
s5kgO5aZxAUjBJzXW8M1VlZMB/HHtjCWzh46QwkHkb7fYJjQxkN9L0n1pzOACbfqMmK53r4vZooW
mS36uIRSaG0J8tXrFKFo8woliVyq7BakYcZWuD5y1/6TYUQGS0zJujsBXoNyeYF0HmM804gvBntk
EXFstKELd0Z2aRRZLETIiNBGqHs1i/c7DBL1KGM43d3F4usL8t5xNkaWTovieEo6zngROLJtX23v
8D+hV3mFeVz6cpZzEjRsGlmJmcKOFyqbWunc8scxqOUuJFOAM4g/yW3vKRD7GtW6SrU6ZxeRgJ2E
pBzeuVLzHMdc6vr40Elr2CakYBlL2Vk/z/1oFhIV7Pj84v8X4LAFk3GNeV4CZfK6CYtW1D5wFeOX
l2h5JIvYm6c9N1UEBoXOteIl/rYw/PIoJpRmefxiWX+5s3hA20qil9ZUMBtkN8GmT02VNhOBNg4P
AQCOTrnGpOBJYlPnCMp1AXxuyiuoQT54HRWrvMB8RGZY8/hBRsrHCUMo3UuoHJcDRQqiOG7N2+GJ
9/IPVy/pL8+P3tsNEYDecUFxBxuVr2ilB4QtA+TIyFpaIH7Ppe12w1Z+/QoOw1SYoX8yEsbnHLx6
LLj1otnJxqR6Yy9deo7Sy6f8eiqEZJIaaHLqMYfdM+UPSPTa2HxxTZdvGFaiLlwzqC7oDYpec0aR
e4UH0rlN7MYDUQOAVjRE3DORVuIIpsHDX6ykw29RHpzldKcH4Mo5JWc4mZUcRkobn9lQhhpc09bL
+P5TROBmLaVRPLaEEaBIx/PVKfoqwPIRTcuVNBJ9zQAo+gEHzP40uL7GpgSibBk0rNhtQOOPc/xS
JGWIE881TVToVUyZEmcOxofJsBJG6NOnGS6rS+IcSXlAgFeY5a3OgkaszucZlDsDQbBQT6EXar25
CpRTeyDG+bv71S+7lQqnKS3DwtR96wSMfScmjNi80TMG4JK4KuuY2F6VLWSsdgvvX6iLFp+B8mKy
W9Y5PCRCDYXZ1NGy6+yfyvDCHsKPLdAPhtyNwYCuAVPbbSpgW6acmOkht7pBJ/GAggJmh1Uz6qR4
Tt4wF71DQ+ZO68kwRcIjyRYWLLOGTWTZECW7oUhEGMBqZEHHDWQeNkka1ZnXU6o7FlpSWIJADRPW
x43nFAN0ZQ5wIKhjLC8+lQd7HNo20auzVPTzSMUsNufn0su3le+Uyz0G2rQ4mTBJmo8DUXxfrqlV
kQBoyG/uWp4N1iFXq7Skgn1bU0AQbNDyfpx3j/vbzRuIBSasK6UgDgGdY0I99qc05Lkbr70aG/kG
X88+rf76y+0mAXtP2JfYZQZiepDg+5lRVop6tb0dwjamC59G+4KexJeoydHkMRp8OTHYeGncKRxU
l8xGqlg6YzSGCUQN0Q17xANCrpVbZbH4OTpfARd1E+QhulIcbMTclQmI2IGjlXSSX2Bf1H93jhEo
xQBGSERtfm8SqJBt3M7jkNWiyTbQabKPyQLg7IBXNGWM23J6fP6lDiYK6U1bRoM0TKhqaP3/49X7
DQZSR0onHQzPbBu7JAESWQnbm8vIaE5C3M8kWGuaW+jIqrY7vAAuozjloHxT7DYqRcWAMRy727oj
RujkRgQoghQwLGirUDyqklN3ZslMtnHe/FRUXoq3o23vVuxUPUdeYOXiMQvWSyrb533nTtNQNC9/
ozzXzESWAmO0/FLCSeThViEtNZ/508JL9c3uZwrjeOT1MDs6HXfVetYRE9ZM6C2X3HdFSsUHvgCi
I0AYIckMsmJdnoKUHCdzFK6Yxk3Z7Hr1GvT5x/6QctyfJVQs81D6VfRagBVQ3LXfe74td7LfFPGx
P60Ahib0z5d8bqJ5VSsBXBMiEzbEmAJyyBYpxWsiEcK79017HGqXy+v4hb02d8QGLOsCX0dAGXDP
dLhMgXQ9klmZxdppkvCmGFBERitNmIzpvxGQ6gkbsgUPY7fVMBiuXMFNoxUJMfQ8VUARWUBDYhOl
KODA8kjk8j8cLUu4DZEfT6l4p8soMVLXOIF5fdPNdMjqM3wXiBFXh2UIfG2hb9YOrH22tpkG4dS4
katcT68x9FyxqXI6veWlVKazR/mPvKXC9cf7GpMjp+3DYXPhZwsIa5xG8b02QTOBbEzeFql8AESI
q50Ij9nfFitBJGi1RpJgE1Rk+5gCtdJrqKMAhzeBxiCH7XcyX+HtCiCG+VjfcOHuuLzDqn+D90J2
CVdSu5Ar8J4I0OhahFTMun4Rh6DOzcUcMs0201jg43ksgkuaafK3MfPTMwWlZAqjHHCLUGYo2Dwv
J0ppMqrNMXs8tZdgTdIyy97ntVTF4b2eB1VdOPdw3IEn9CN1zKoYAy13iviUV0eDfA2KHx+VmQ+/
ZbF2HYRP1ubi/UrKg3zZecZ6IYGEMkyMkkjiYv0H3X1cOb0w4cJfHzXuKKM7KVg/PfD9AYOoj8Cc
Qw8Q0jMiNiJ5QQzopaV8acKucR4Uty2s9CCTx8dxcjn+0geZe42ILg9f9Qo1VFz3ui1hPaB5MBGH
bknSpVcsDuE7y06NyNh6iarZn+YTNLHLbhkt4BRQ6v3EMcNXsUJPrgEsJU4m1jyYKDeleossjbXF
QOv2YVmelj1TvBzE65N8TFiPLubpOn3ShKCp0h3j6/lutqhiKUXGlaRtjaZdfssTfVWhH6VM1eIY
7bnZKRJ4ZZ3CXkFDKx5Y5vkGDEu9zCbgkuadAdwu45NyBE10A1nel39h31QKBFwmyyN/4lvsO74l
mb/79OE779V4t1FSTYBSbIMDaJxKffuJMS5gUCbPrlrClQLgkKXrUxw3RY86D/uzGM2OGDPk4GuD
pgfsNaOtig1PU1BDfgkdz5XkCZP2F38bOxuMBeTdkOclRoPG4zKWl7rNabxghSk6PHmoKn4t0Y7s
G+69UYftsT/XCUZOq0ksRMj+1mRcc/chQCo7d0CgX6VayE2USOdHe8hnvKBXQCTRB3ZSequ8KDTH
fWtEw9h5o+AJZqHKfFheus2NHLCL6PTNYUFH0V5E/+r2SQoBFSWC2NmyQPeDfLIkMNatzRVMAUYs
WEgp4Q3ovu6nO+vDAcSkKNR1GN86ZthAWHbkboAkGRcOgRVk+/pv3TsNe5OH5fFO8KKRX99on9g0
RQK/AiSqpKU18Fqx7RSj5H5K2YBBWHYPReiQISWF+98cDHf7urI5Shs/YpHXo5F3sqpbEXE5bJBi
JS/bCGHBjPazwpds/q720yRbCBpx+By8DP8ZdtMDB+rPPYWiIX8wcLT7QGOngmY8TUYQezu14Zjh
HRj+NSZdhohiGS8wNrU1vQ7u0GIecJQBcluONbs02ZpAkW77Es95mYiBIstaQQhD3zlAkD9HhLsx
ImIUwkjOIF3ab1okFg3pHr3GzxvifnlbecrfuAz92eBdeMux+h8zlobf/cDRUff4dBF6X7oKsEQv
jOMZflLRgYYZJ6q29VEV4BjVmgxU58P6JYAHvJe3909mValdKa4ymO5+HtIzDluQJwUJ5IdWXVT2
8WOX5vnbRoX7Kz2smjW9b3zBqeA6QWBATq+RYXAZrYJnGjLnSlmEJgi4Hm0j7oZG11mhUB2jTZcU
lYghKkY7IIucy+dpDxI+zyTfjRXiN23iyIk7nIj8FXfzl6K6bH95+bksG/dnWdegWaJrxYdomEfy
hW084LVBZs0nGFw0i8615IaGa+jgi6ytvARCeEq46oAKArKlmVhKtzzOqwxEGIL+JkLRfjE+Nlfv
CWarrY6YROMnDEQHY/QAXLG7lBzZxPtVmkl1hQQXF610C7MBWPpW9LrPlN99Zav5wuwVwfm5Gcen
FYDE1Xc7RN8A72CT5KGwX4l9u1ScAa+jxjXGaaJM8V8g+thKJvI7bu2cnXGDbmD9Rcf8HQOvDIqt
SkEWSRSQslcJPzcitazY5tMrPhaXVA4UdmMIRSHUAx/adVXgL3lgcMwYS+dGCOpgW25i4B5yOrt1
FNy6HIjrbBqe90Q+gix63MSH3FVuqq1dj0IWrHMMAgiZIaVvgIPyB0D3ekZN2jtS+Scd6WW2DAZq
f0522nhVqp0u/i3jigcc5oitaqDFajveuqqYqWM3dI3oAZs1wwimOxTKh4+HorwqmbSeqnkZ3M5h
H7VjsWUh3NP3yJD96GZwvoHu8JCMqnoY3vJu+1LMFPyC4yO6gu9iL0jnqepoZOn7GIkqllhlAidN
3L7LTvQXORvC89LMNN34ycMpmvczEiYBjqaXGak9YYfOqwAGQtfvU+gQeQquynf9+cFH4IZYDLg/
YLKbUCSm9VszlPLXgfOHvgbmbog3yhfd1q182ltHjM8xEhQJS/cBVYgtKXTIWhe87DIIbL5Vx8+l
C4Gn10umkZSP/s7Zn/gRTobN6V1PBueAWyN6rovFrErB/g+MlZ+1gEY72L6Ts7M42bes2Gt2jZI9
NMmkAP1JdDsgvW+gsArS20/i6crWdEP/c261LXkIuonBKPtW315+0g0PITSgdIon0b2HPMLiEzI9
J+1nVG3poBSoQrQH1DNl0nnKvclvb+w/EIKEJ5cZay3JEWACp9UXBSUi7uSXhkunzvewy3o4NHR+
8O7fJ4qjrg5Tl4HAmFmFcLYuSoiSs2NGndkZgeNBMlP67wCkWhiKm/qvafUTlvuEbbRZhgt8nLxM
StuvbeGqLCwT6d2ClBiYIfFyLzSNT1n6DogOI2WNi0q8k2WRHG80aFjOJh6wgxs4LTt+avwTfCaR
YUSDH10zAucaW+g43KVupIhDtt8yYckrcBqczMORB+8Zw8F1YmNzGpTXCNSP+pqazumVuWQTVSh0
BpULRLvcd6iPLi5EZRprqLj5INXinCmbVMo0ogqXRFhH3LN6nVTvrg7GsVwiRJpNcobZKD40MiV6
JJt2OsuaUmFMOeeO6p3mJQL2qZWfFvCNE6aV06xh3C1M9qvS3gjDyw1zbdMkIB8t0xW7XI+QzejY
x0gdVsU2ma/PJRLP6w==
`protect end_protected
