XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��yT�P�L�{I��Y)X���j���K���r�f���>Q 6�:�ϊl^a�R�B �W�M��a�6]Ô��q���ƿ�}�]�d^~���q�0�����m�x�Z�g�E#t�wʤ���b�� ^-1B"sD�uO(��
�O��H8���KR�嫛-4\�����4$t���)�s��?�3��4�cд�c3P�e�;�]6��L�:���q�y��}#D�����ʮ��v��g������P�6�u�o�x���'K�L��f3�Ϝ��Tg�3�Wk�}�o!#E�^��W զ���rAA�8t׋2S�N���`��0(�
�KѠ��|���e���U���C7j�3�,Nl�U�c� ,���������ɚ'�)9���;��<���n�(�{�(�^tD�v�5���&%2������j�A1��A$�r��h*E����n~����1 �
�0/���ϭ5�~��3粷<CY �SV%�(1���
�߮a�c�W�I�NB!^�[���l�i��䝣�,�F�3X��#_�����LZ�p�cO���D�|>Ԧ/4J!�m��۬��׳��� �X'0���j�w2� �šۂV�cA
�����T��+���	X2n���eK���6��L��o7Q!�PC���G@������=
���WO��ΪPUŒص�d(�S�t��s���J�?�P��VFE�+����~f��4����wN�����~��>�\��2Y+a��qԴ��o'��̀��XlxVHYEB     400     220XK�i�P{.���RϷ;�q���$C�����QXҲ]�D�7�>������W�ʻ�y��%l>�<��Ԏjm�t���! F����z�-��n��S'/W��
�+��/������Yvђ�XWL�gP̓�8�h(O��,�QU�:,��J��f,��j�c�n�	gO�Wbl	����h.���qimS]@^�93�H����p� ��6�Z���<��c�W��¸%,ۧ�y�h?s�x�ӧ/�y��D6}De�����ƅ@>-�%�5ޚS���S���W �$�g#TC!�X�Eb�`g�n�d�wJ���4@���[r�iU�rGlu~�2,k@�TU��[D�>���S���]������@�U�a�[� �����p��C�8���[�0Ҷ@�I�9ߡ���;8��Rg��^�	��!��b���&����<M��I��<�P�$TO��r��}�������C^#9IB�c�h�i��n��4�p�c��с.^�]?��
�����k��鐵m���%L)sfi����XlxVHYEB     400     220D������¦�l�b��C��_Ƨ����eⷾ3�V��M�AUu{ń�J��a=�k�\�rw�G�y�\F�T,��50a���g��r�)(M86�B/�7���F)D1_��TD1�l�'FX�\d絍3c0�$S�N��J�	^A�
���Ē~"�a�Pֈ��r*p;��������"����?I��5���~z@��N�f��u� h��X���*.�{/׫�����F�dO�nw/� �}�����/E��F��X�2&��'k�Ƅ:ȸ�H�d�iГP����Y4J�l|	C~����`�jv>�щd�wQW]�=���T��9�E�,�},�+���OQ���fT�2��i���<R�)4�n�eSؾ��q������ܮ�S@��[*�254��T|	�i��w�o�R�������%��+b��D�&%�;CV���숋��A,iW� ��d*�[x�PW�s�ޛ��Q��0��$Db��,	�Ĕ��_�[�`a0�n[r%%?�)��o_�P�.:�d����]XlxVHYEB     400     1a0��Ѵ	��x<������*�;n掳WI��X��9l�7���!=�P����Òb�����Wz�/��)��FW���<Y��ꗽ�-������L��=�����<DsW�ˍ��E>� �]�,�9H��5|�Ջ7����7�V��F�~n������WD�Q5�1m��m�܇�,s�G��l7�I6���Q m�{�F=�ɬ,�nr�b�7�c�B�J�m
�}�I�*h���_�SA.�A�L ��i4�͎)��ㅫ�X߫�|�C�H�ֈJ4�v�V
��H�\s�a����n��&��f�[��ViJ�jA�TC�w��BH��;�:F�ܑt��/�U��C�lP���K�IJq��0+�_��c��PɂbH�|�ā};�!��͝Ê�=�R�ЈZg��p�����XlxVHYEB     400     130�	=<w�6�� ��!U�@}~�����я����T���������(y��,��g�Q�$.�����v�ϥF_f�������o�vw;��k-W�o(A¾>�7cʘw��&;����u�ga���{^A�K�Zfi�~�e��0��<��wm;��	�e-�l��D�Mk~.Nx�Ћ���퇔f+m[ȾFs��J{����3߷̥xQ�m_տ�I��H��^�������cC�0��kV����ڷ�Bh�xQ�"��,�Q$t�Z�K��Q����4)�����tz��k�� ��C�6XlxVHYEB     400     140<<��Z,��>R�k�J%���K����wa�5��鿽tL���gG�V�������w��� ���&�7���4`k�T�N�ǂ���/�s�%�I��g-���u|��ua����'B����qܨj����� N-�u��4�ܕּ���2Y��X����֠�+��ꭧvl��Ͻf��y�Xt�R6�T|���JC��s�3c87!�c�9v@z5z�e�ߪ\s�*�ջG'���D� �}W��R�������~&`�sj�#���n�ҧ��c�d�k�޶A�B������:�W����_�3�]E�j��(n��;�XlxVHYEB     400     1c0�b��N�G�[����!��v�xm�u�N��3\�a��a*�0�/��}���(&�(��|A��
-S�!+�r jv��j��|]L9>��C[����~�ɮe��ކ�C���!75�4s>�A_�R�{�e�ؔJ�nW;�L�����ԣ`��C@�e��}�d���H��Q��r���$i{����5�}���^����GD�Y�Q����Q}���j)�Z	����:Z�	i�T�cd��$X*n�;m)ݡ��Λ\��J���@��y��������F�N�4��
�C�R4�8��D�E|���]N';�m5�G|�q+����q����6�U�ܲo�ΤN�:e�9r�,~F�K]�I�.ߥ+�#�Z�����*N�f�u+�bܐ������>0H�HǗJ���0�Z�]�v�5������m�}�-z"�x �6s[��J��n���ߢXlxVHYEB     400     200��H0���)��ޙeTMK��OŇO#�L�EF)�HZ��4���2fGpR�����MΤ���d��DVgG֗���SW�=�6���U�qՖ*Iΐ����ν
��M�q@%��d��$�K����;&~�T��#�+� �U��z��w�a���j���3[�Z��]�3Q?���C�ئ��u��i<vi��w��*��><��d�),�b��F!ʦ w} %��k[��7�k.��L�w��$��d�Ϭ��a��c�mO�B��B�GC6�ӷ^ ���2o[��&a�Y�P��1�aT\RY|c�	3��6ۅ�K)�Y�CW?��ͼj���j���s�;�M{�͟�;���yF��� ߕ�x:�j
R���Q��WC7JO8�̉U}˞Cy�(��N��l�
�Qq��۪l�G����/{S%�4^$l53��E���Ng�1;։,�$�[�F�=�����l(]��O�:ZwO�p ��f��A�XlxVHYEB     400     1f0nBt�%���m��
���G~�_��
m͡Y�Ǌz�L�P���y��n�2.��BB���}���7��\"�m�|@Ƚ�fÝ-�N��6��Zlq�g �눼�k	��%?��r�(��ʎ��.�d��w͟��]RK���wANm���P�����|�;l����:P�wCA|�� �,���Rn���*�N4R�k�	����&�6[HA��5
�i�u����X�/&���]�ް���E�u��q)��c�A�.f�4O��Ο8���#�V��[��hR����%snlrGZ�m����s� !�.��=��f�����7�{-���U�`�\���Z����{ )��DS�ǧ�*�K?�ut���z|c�L6�:"X2�0*�B��q��	�����pQ-��<�$g(=j�Jh��Շ��@P��=<xEÓ���D+c9F�nQ����o���<-^���\d|8�b�����f����]Ѐ{��؜�����XlxVHYEB     400     1e0q�k�^v�K��5s}!!D�r ����$v����=Y[o�iݼ?�CHc�e���UX�7�[��[RB�R�¥�%�Gη����Q5�1Օ�%��Q�o�Z�H~��qQ4��e	���^C��Q�R� P��>&��-�e�����<��w��S��v~�������fԻԖ�,�_���H:��/�#鞝��4� u�j�4蘭Z��9��\䃙q*M�`R��_Я�u���ǻ9��=ŉ)#X(Cd�޲��ĿWj�ֲ��e��Ub��3�\/��Y��-�Q;�3��$_�X܎�'�X��� �@��� (lR%�jbp&��X��-�46Ҟw���[X؀{� }9:/�3o���*3z�%�*e�����]~��߽e���?q�7�,jsy�/����,��~��|�/0��}��=1������s^���R��f �5Aw]m�u0O�Ռ�mǵ���^�P�A�XlxVHYEB     400     1c0�Yͬ�N�M��/�5�s�}��m9��:)���_��֑���ht����z��A+����+<�j���ܸ���5�kNV��n���"�}Ũ����?[�M{=	�ʒ�;������	�G݁(���)�%X{��B72/��OTT�qH1�&(@Ǣ�z,6�s�"�v���If�� ����݃G��N�O���g�\� �"���^`c��E��*��x���L6�As5{Kpe���ٝ�w�!B2��i�n��u�pI���-����i�C�0�T��J�QS]��̆=���z��R1��8a~.!vJ*O)R Id�n�B=Z��%�i ��h��CG�-_}�����H������{r`����dԬe؎7MM���<���X͔|�0���׽T:��j +kĺW�))>(@��u�g��а��ߦ����z������73;�vl]XlxVHYEB     400     130�AS7=���4���U���]T͈�C��ӗ���R�_���gl��_�Ę�⹷vS�.w�)~%�+����D���=�e}��0,��[ʪB���v�*f�vt���\d�����DOQ6tb%g���B�����]H���$�q� w�T�{k9��a	e�_�q�`d3���t�J<w��f��*��Pao�< �D��=~��IgL�Gd�g��li&�{Ĺ�|Q5�@��H��-X�fG.�@�^�q쇩W�y.~QM������M�r�V )�3����<���_H"+�i�e:��2���XlxVHYEB     400     170�:Ռ�q�3���Q�j����'<�&L�#C�6ú����� �zn<�I�rT��س���M�Z���WYK�o⌲�ؓ���c�dn}X�Q��V�~<�*.`��.�rXGGo����?�ʿ?��	�ٚ�[��H�����[w@Q��_����#����7��e'�tV�!R�&�����Bt���b5��b�J��d+�7[2�VG?�k8��&�|��؇�AU����1h}�PD��ula#M��<ӯD�D`��
�-r��1(H�Ρ~lƪ��9e ���X,,�g�vJ�v{Ҡǎ�!�cS*}��=� ���<�Q�.mX�Yd��{-��׀+7�EW�{��XlxVHYEB     400     110���D"���HS��\]����ZFlߌ%�'�����#��N*��G�/�H����g�3,46����lK�fx�a1T_�����`W�J�Bغ��#�>�GNgP� ���!�i|]�k��8Rn	�+�b��9�T|V*su).ٹ��@���{|�80_/���g���8�a�2�W�l��B�=P��Ȱ�U�e$[��ʖ��t��}�NXK�Cb6��P�6h8�I"E�ΡG�Q\�z�m��L��Mc5/�|���ɓ^.0����������m�XlxVHYEB     400     140�n���q��GoHE�#��H_����y�L��wP7ohb��{�Rxw���-*�y3�!u�<:�%�3[�A"ERy�WK�C��F�f���M�&�����q4n(��}q{���򹯻B��E �p��mKh쟟��b��HFr_o
I@� ��⚞Hp�ϞG+�ވ����l'��o��s�<-yU�D:����0��/�ue�;���%����j���R�*\jw,X�D�2��F��T�>���U�lOG#¶��)=��.���Q�N�-ф]%��/mm�K��O�WA��ގ�
�@���XlxVHYEB     400     130�^�+��o�lW�u�Z�T�Yb�*Y�� \T�E��Y� -���Ss�
�Wj�?q��!m�T��lQ*�X����Jݾ+o���_"�#ܡ�j���������Yq��3��Mu ڶ>N�*`4�@��uE����.���l�	=pڂ)sD֧��h� �?8��k^��m�&M����N�&`=�""�4�3h��|��^$[�ħX$,TֳH�$���2�K��F �>�`�y���$<�4!��Z�`���H,j�j� �
�����&�<n�$���s�B�֏��*>P�(��2	���|�c	XlxVHYEB     400     130'����,!cQ�����E�a�br��0��9W~�����-�N��&n����-�L�ݚ�Fj-T��L#�\_�H�������jO�2�(A�R�Rl*�lr�=S��	TԯP8���լA�k�B|#C�F���(ߡ~#\��r5�}1�~��oK�kk_r:$&���G����1�D,���
�+s��8���Wc���J&7]�u�^���r�˺���[��ц��i�QH��HW*�z|)_7n�v�i���~�p>i��%�>������:��$��k�Bz[[��}��^����XlxVHYEB     400     150�z���n֬��g�c�A��߈4Q}�����{�i�њ�It��T���A��i��_�$���'����"�?́�!��G�}Pqn�L�kCs��F�����F�J��FP�������I}d��2��?�]N�Bw`0H�-�����\o���^�6�n��]B��Sɳ{Pފ7��̾�|ı�*�&s`U���D`���8t4��ink���;~����4S��_M6.���+о��M��}��2��b�-ܥ<�3%9p��3i�8�-�q��Y�mpuf�(40�#@���!�h������a��#���)EI�2�q��>s}%3ޯ/t��XlxVHYEB     400     180!�I/�����Y��kם�t�|]�J�?O{����ؾ�pj�O��Z�6�],��Y�\��DO����G:���R0ɇ�����9��mp|Ȟ��C��q��rG��k�����=�m��
�*���H����{���=�X�Am�{̓�r��R=�,���6=@4MST���������$�S��)PM�o�q0ܬ�V�5=fT���j�~��cf� =�O�E���������X��YH$J-@����V�{L�bu��\oo	#�2%�q@���֔F���ę	6r��,LP��Q�aA��Cn�
q��2O`b����Q9)�[��O��Ǣ+��T��6vF�u2d!����*L���`]�FA���XlxVHYEB     400     1d0�i���0$��Р���	?/�2#ѵ������@Z�r7�y�P�K����!�L7�]6��k/��Lz��u[��(���Ip�=�CRMA�ݸ�ϛ������w	�3�����v��I��H�����e�$�p�e��IK��)B&�N�#7yޥ��'��a��M�)ڭ��-9��oF1�� l?����R�rz�`&'�ſ)�as���?[�Bl��-�3������D\�J��m܋�J3	�Z���5!Y3Gf!j�H�P�¡h��K%�8�#�!�pc���nuB5G����㚷��?������::@ɨx����D3A�Xo�+`.z�.�x��<�B�U{�4f�&���/�~H�Ft]�h�F/z�,���������Ӧ^P��#�u��������tvFJɂҶ;�`͊;����p��S*���d�uR���P뀶�~�j,ɰ��)���0�6�G�l�XlxVHYEB     400     180+�*_Sjd����V��,Pm�R�p�Ȃ~�wS1�y�l(&�pp�b����ǟJ�;8:�Lg*N�$����$O��
�w���U��q;�l6���� ���6M�ul����`�NI<��d����:"�
�ߠqp*K���>:^Y���Y����v���{���xr��%�h�~���[P-���Йi�Cg-q�ވ \�V(��n��ށd�5��������)��D&��u�u*�gJf��tڝ�� �}�G�p��;]~H>�S�F��'�q0����VN�����&ԼfD!��ދ쌋��_��H����'���iyM��&���Y�5���k���8�x�{�02� �> *(��Jb?�f�0:�a~�7��r���l�-XlxVHYEB     400     150հ鑫��i���M)ś<rOV�=��~U�R��3�N%���2d�[�捕�G#�`�
ۑ�'G�}]([���;�^\q�,�K�
b �9`�By��.�l���-��}��f��a������(�C�[�{#Z����Q��~��(Zv��$'nf�t��~M�X�7#=@ol)P����|"�\H��j���ů�}J��	1=O�A��i�n���GJ��Q;6�q���Ek''�~k���B�RN9/�l'8�
M8�Qe�g���Կ�~w�&�mʶ���`���M�����y��������X����s)˥�]��
 �1I��hϏ��C��_��>XlxVHYEB     400     1f0��5�b,.#�G�%`&
ۚ�~I5_��,����owf���;"�e����~���J��6@�K�/��t�D���2����ȿ�gZdr�n�zMK��(vq>D����]ٌ|�ۼe)M�;���)?Ю���dE�iǅ�8!� V��+|�� l���b��  ���S& tc23g�v����8 ��3I�x�&��:�]3@^O#UM�y��p���Av^ڤ���+�^u�^���!���bg�/��/	�I#`v���!���Uƙ��G	0�<s��h_��M�������i����}����Qi�y3f_��)�2.���j�3P�E��L&��r��lt�?�F�e�H���p�rwt!@�d�Ձ@<|� �/Fu3;o3f�!�e0���i/jd�g�3���H5�ki��؇,��M�;}�F�Y��
yN�릱���e'\k� ��bDU�_,����բ�$rԽ@b�l"+��P�%sw񙟃XlxVHYEB     400     190���cfh���JH�Oa�/�'\�������,�\Â Ԇi�t�w[\fS�f>�${����<=�QmvX�1-;���dW@]�Ţ@��[np�1�@�L��/4$1su����8��n�aMQ�j�ΓUA��,_�� ����>;=�E����$��������T_���٥�p�8iq館^O�)���!�#��AW3W��'U��HZv��s�kښ����-�b�#�	6����ݶt�7����$�>����OvT_�F�}rHTV�����O��4�� K5�w{u�=�C��qP9���	S���o2�eG�V[���s���d��(W^����'�'.{I���ጚ	��N��oB؋~@	����I��=��ڞ��'v	���v�XlxVHYEB     400     170�.C��U�,c���4>�O�TN����ӄ�B1'����\�D�1Z�p��C��W�чj
v�^�kLn-��s��{�3X�#���goҼK!`%��V�����ԃ(���A��#�Hf�0M��px'���
���h�f����-*�5Ə-��e�s�R�����0r[�3ϻ��2�֬�	I�h���|�Q�u�y)�"�F�_�A�o���dt����2��U%�ZШ,���|�4)�7�-̖]U�8tܷ�GϘ(��기�z^�O�R�����6�_M���Eg�,!(=�7�vՀ�I|V��V>ӏP�7��lȦ�^	��o�-�$ʗ��;Y�r��m� 1�P8��%�P�b<�XlxVHYEB     400     170�g�H���.%�1\�=�F�j���įnȂ��f�9B֤|�~D�:���������=��4+W�5�<�*yq���5�>��� L$"*%�OZÃ���%��c��J]��O�K~<�'o���^�����+��`,�u*�Ips�zB#k*�U	��&����dS4�9��.�H���0���!�x�.Q��)��9��{��kK+/���+&R���䘓�?���ә���j(���S=��J�/�Ʒ�����������Aj�Ha5e��":4J]kC� �0,��kc��%wU�u,�|p���3��=P;��
�F��m��~�}x�!���R�F��\.��2�ߖ� f���@� ��j��G(XlxVHYEB     400     110�G���������$����V,CTIIdyރ�or��֮<VGK����;CQupVY$^R'��	&���q�o�~�|�����}i���6I\������5 #-�߰��B�Bח���G�ꔺ�m��B����?�<��Z�."ʦ�XW ����,]Җ��������b���ё���t����"�e��	n���,#C47-%�i~4�u���V���� W.�p�ڒϚ気(� #���B��Λ|;��ZGG�`D���3�IXlxVHYEB     400     120�0y�f���$���8�8�3�N]q2�,<��~�M{<a{���Eeؼ�~��P�� Sh�� D��v�R�T��-{����9�s���g!4��?	����a��.OC
��$��D�l\!N��v�@K�U �Ȭ�|eE��_��+٘��~�����O(�{��~��q��!s��.�Z����~��}\�^l���Bʓ��	�ɧY�͵7��Z�{%�'ػ�h�Fh;��EE�Ʀ:��Y�t,�����+�*�w ��g~8sf?m_����┫^��j�v��m�h� XlxVHYEB     400      d0��w<����↑��4�g����N�>xM�/I�����+�M=�"B�r$����p܃M*���D�!�#�"��Po�e|1���P����-�E��a>�,�sw�	��Mc������ ���a �~�<������c��ן����V]g
��x�q�7J_B��χ�7��R:�@w�������M�Sҿ�A6�4ql�y����XlxVHYEB     400     140��	�#�.�j��I�8iŦH=ť����b�ݠ2�K\/D��Đ��_kE�O��Zq$�ҝ[>l{��蛍	���P�MFL��C�n��:�O����S��L(㈑�V u��?>�\��5A�H����:�7�|�q��]F�e������P��6U���W��^'�B�=�߄:�9�#h���y�7�������_e_��0:���ں:��rɟ+K܌h�9X��J��{��n�*	ݔ��ٲ���,�x��C]�w�d�T��11�J���>"�	8����~��P:Nh�������D��ߎ��k)
Cd�G����OXlxVHYEB     400     140hW!���(�Z��J����j�j�����Dqa,�g2�gc(�Mp�V(��M�c��ѭ��\~�,��Wr�3w�p}X�Kx�'��� ���/D��?��z��O�i��_=���^�z]�R���F��#A��[�q��%����!�HEoCȸ�I��ŵ6�M
��|���b�h\���׿��XbϊM&מ:�	�(X�[��]U��X��=�t�a/�i�����b>Q�Wʍz-��x]�$� ��*�_t����>f��z=lZ5�=����^m�  ���L��LDW���1��ꘪ{�l }�0�9����p}��XlxVHYEB     400     120�XWV� 5"���S2��&�Gw�z��齯��lp��Z�Ǘp�+��\(�M��������9Xo�e�Jio����R�>��P� �~<��M���2�8W,�v�7o�@P1����������Y	��/���j5qxJQ�N{.��g�e,}��Te�J�w�w=y%��t�S������2�[�Q�d�N�A#h�&I{�d ��	�Sv�3Ի�hv6���Q8Jëe7����@��%���&��[�[D�ט�Yx�R{m�SV=����pZ�
�P3,XlxVHYEB     400     1a0_��uq�9�����cԶ�F'��+��� !v�D>��97�!x�}�7bY�[�y{��+L����/�{	Z4/y�2hW����Q͕���D� �L$���A�[���d�Է� s��@��B���%�Wʃ��i����Fa���D�2�=�@s��r�_�J�A�����<Rg�^x�����H��{��jX�� �5zDY���$���-��X�K%����ٝڹ����^/3�����Qg�qn'v����Pv0��ɬcMu|�/u �C=�:W�n�ڹ�}G����&����ܡ��8�?뜔P)�����,���ź]C���N������1���@E�Щ����pw+��	[܊b��v�+�߳�mw���u���{�|D7XD0��v���T��=�XlxVHYEB     400     120O>B?�����*}ܴ�1B�3�bN�y���\�jo�ia�O�3<��$�J)����� .��v	�~%�Z�ռ�ҫxܓ��ݤ(�cl&����,}�U�~���喈��"2c�銳a���gH�U��3͋iD��?BP��jX���ɜ劃�a��l=b0���J�fI��,��^��]������v����d�h�[;����D���557x�g�225~��Ԍ��������ٓ��7)=QT-Ȑ#��̈��F�w� E��-0m�3�d{����J�i<��9XlxVHYEB     400     180��A-�`�6ꇖԵ{�v�5�P5��_<.a4ؼks��O�c��X�Ok\���W啗�0oJ'g��+̣�m0���tWܝ�w�:{וƇ�O]��:�/�!��(�C�{�=r��ƫ�BZ?d*7��\���M�(B
�bqV55C���~z����Ȟ�#�E�����n0�����%U���g7w�t����K�z� ��v��ƾ�*I��`sM���5-�+�=0�L�d�`�^w�ơy�f%���3fj˻W�����-�u��!8�gʄ���s�;�6�sNFۛ�Z��DzK�B�jSҁs��dbr;W��������e]db7@1=�G]�0cA���Q_d@��I����;�)XlxVHYEB     400     170�cUS�
�:��AZeF8e�#�3-,���c\����Q�*��&t(B��!���b�p����b�z�~�i?{ͦ1�D]UKi��G89:�57p���ٵH�
��(�,}����#QԡfJ��U��#U����H�V��a}�n[I�	��b��'?�Z����ԛ��~6с��a����'�m5d�b��*c�7�T#���]`�
Pe�}阎�ep�}��m��Ӓ7i����F�7:
tb��f�Ë�io󋍗�o��.ޣ��&,���SwV+8.8�9깒w!�@"�-��>�S�ݯ�_M�  ��  _:���DS=P��X2Z�}���"po�v��98�+X�8(��\�I���XlxVHYEB     400     1c0l����	�&i�4u�	��w�������O<�W�,�Ol�܄?���9�8���q������rxy�OB�E�8m�R���?��e���@��F�q�86����l^�c��M֝�ӿ�Z��q����H��X�8^6F#8��[U{߽�.�|���!�U6��w	���ba�����w�x�Jpm������W*��[��+J�o�m���#%sX����������r`Y�G͔{�>I�#,�x�L1� #x �0B,qF�^8�+�$�P��4�&��Lc=��I�.�
��.��(��&���Hk1�>�4s6�D`�jz$�^�~A�]��33��{�ƾz��U7 �����s*�}?�����eu�b�FV�~�!Fq#�����B�$P�� X�!N�������P]slZEv�,r��+)5� VϐXlxVHYEB     400     110B�I�B�F�U�]��Ơ�dk:��Jd�a���3�'�y�`�4��g$2 ^�����G`���=������E�ʈ�sJbid�� "�.g#��5q`���*��Êf���+`�\$�w������g>��c���^9��MHK�xY���r�j�<�[s�K�D�b�Y=�:k��^��<��1�<H�f+tҚ!3ގuM�x�3�z�vێ�f�àn��sW��2��g�f8B��V�OJ�t
"A?lht�]�ʷ�@v~k[Z���$&�e��~XlxVHYEB     400     170r��.�׾��v*^~���-��- �k�?����8>��aJ�dlD}'�eH4r���3E���L� .y#�%��CZ�e�&\�/GKD��L��������-�G:�&b&I��A�VVhI�5��V�a	Io���E�����+M��6��ﰫ����l��3=Ac; I�-����c��q��ԯ��3#��� xM��=�_�B"���r���	��+|�(�X&�w	[Y+&+j4l�0�,����|v3]�C��H�Q[R�][���~�s?�J��/�ش����~Q��jQ��o3�<����K�.���g�u?D_ �Z�{0�B�zNa3û�(йKm7e�i��I��9�>1��VXlxVHYEB     400     170W��J�Ay"&����+���_�S�N/n��c����o�l�)$���(??�=��ӌ1�"���C��qB�Ј�<�%)�LM7��ڽ'��(@�2n,�^(+z�������7v�UCn6���_�ӆ�;��S���(�;~TX�86]���IP�:���9y��z���&�N�i�{�>5@���_�G��5� &��+u]9H7�u2tQ�{�]����m����K�vM�{y�8 �K���:����V@/5�OɁ��r�~�" }��u�iT�e��W{0 ��P1�z6��$��@��NĘmUF���M���O�$��9�I��E��wd�u^�m��U�!	�-Z�)a��㛇��}�0�XlxVHYEB     400     190���n|'�I��x�����UG	ְn���h��pv"j���E���������h<ά75|2��OvB�Z�,k���=��������3�\�%=��쇛y�n��==��V+n�
��8���nP�T����w��y�|���S'�d����KX��	|�8g,vF�1|���_0�]]�h����rr|��\�tA��B�[̝�}��W�29�D�9G��a��#�*ĘksԬQ=|�}�B(%;S���jb�m=�p�d/��#5p4�N@���FE�M��}xCa�V^�M�g���vC�*�Da�;�]�"�2y��*��ϱ ���]���-n����Z��KS��?�,2b�d�vS!��P�q��d��8y��ۍ|�ǫyA�JЪ�XlxVHYEB     400     1b0���M��DD�!�����F��s�M��;�Õ�e��C�HsA��M&I$֮��\� ��n�RAn�,m�$�1�i�qts)�!�Bm�n�c�)0.��~�-"�/���pV��Z�fh�3[f/�HxKU��֓�p`��@#z�if����&]1�XM�ػy�-;�/�~*}��M||�E��Mrk�m��U�L޶-��C�u5/��H�'k\��!u�d���罥�r~���$���"�@L�֢H��\��(7>�u�6]3�޾L<��GA��x�� �.��/���D�8� �}�Ѝ�S��H+�Z�b��]��>�*���5���0�����S������@y�c̳h��;�?Ps�b���[��S����v\7�m�
��0��P���٪�P�I����m�eGXXlxVHYEB     400     1b0y?�s��2$�k"і����^� J�o�;�M��I��06�>g�J��;��d+{q��۾#̪مC뀖Gڷt���Co8�B١a[>w#9�̮���GC�Vz��o���Y��'��Ö.�yG�k���c�b�hKU��}�0q�>��T���v��+v��f9�Ep�B7u��:?�*�y#����r�WJ�˿$6f�
 �js:79b]�К�tg�S�e�餈�'"�ȘX�X9 |���]�#me��YI� �,�D¡�-�7���d���߼c_��@�)��hf8���͛��Yy�}�����҆x���D�e!��V�1�"-g�� �Ҡ�)���99uh������kO(�vCB%N�uy9��)��y�8T4�� ��ʛA�.�aI ו�%0B`6'RH����-/�P-1t�m	}a�XlxVHYEB     400     1c0D +Mj���v�n���>�" ;��/�#O�~��|��A�2|o@�M���,Z�x$��"b�4�p����5�pը�bvC�v-�q����;��J�6���$I��¾�\�Ҹl5��ܖtmkχ����@�ؚ"F��<���6i�e��vAC-��
F�nnL� �	��%;�1C���;1
�,&�Ӻ���;��@�8e^� �����Z��$j"z��H�Y2p�v�jզ��}�uſ��u��1y����/vR�-zgE����_�M�~.ZX�oV6��=Q��5��2�Z���4�����#g��� _^�m�M,�鶰<H��M�r�A�6et���� �Z����#j�Iڅ�j���^̰�~(��Cm�;B�\P��dؾ�5/��BH��͗q�E,�2T�:7,y��M$��q�8l}��XlxVHYEB     400     140~>e�ґ?�ŉ��Zx��1~��~:�ϓAIeь�X���8M4#���.�jv�龲_=�~U�c��7��aƅ��Gy��Go��f���䐧���Y�?�rЯ5w���:��RĐO���@1�G.�u+GO��qs�-�5��(�3y��òp��JmI,8�G�F�0�}��y2��	��$��Vc]R�h�E����QZ�3�4B��7_ޙ�B��u\	����VA�=�X�@'�d@�&��* �t`��ɓ��&���f^NŠ6�\Ւ����*��*·x9W��Y _�7-�=���,� ��}H�vXlxVHYEB     400     190�d�q/+Gx۳{W��1�o����`�q��u~��0��I|��y��G��6�,@a�6�Bp����8�̗��a���������Hi��@��U�7`�7��$Wt��)ܶ d��PИ��|�T�U�qs�\\0vN�,���۠����K�j��Kk�v5��J�OkYr���2'�C��Vi׿c��� |s$�z�=�hS�nV<����ϟ}
IQ�G*ȇ����ًB.��l��aCPY��≴]���ou�zۥ̡����d��*�(Ë��|��
v`�r�n��cA"��dT��t���JJ+�r�t*�koWLBON!�fڭM�zkB��O#��w��E��5����^�
����p,�Z��ԭR
^�9�Ԇ�����*��Bi��=��PsXlxVHYEB     400     130�f�V%Xy�D���(�)�p�Ԏ��头��r!��s=b9�a�t�Źΰ=��Y+Ms�_ʹ�SU�at��`j�U�����"|�F�D��I���Р��=<�ӈzUHH�@�(8E��t�
hՁ*�qd:���l >��#.�����I9HM}t�Bؙ|0p�9p�
�����I�c��;��6{�wBn�
�S�
��31��r�N���ߴ��K�J>R�G֩N��z+W���c���{���QiW��@ʤs5W��sl��4�#B���8������Y����N8��9�l7�KJ�yic?xgi߃&�|XlxVHYEB     400     150��c�C��sGj?Vm�,�W_��Hj&*e��� Ί��C%֟n���gG�gRuf���������$%�d��Q�Z+�
"�ii��/E��	20Vk�؄V�����(�z�(q�$]��&h� `��x��<��h��(��������#�+�)���I�Й/
�XN4�d~e����HAj"z���-�����n�z���̣2_�9CZáJE?���wG���IF܌f���������n��*
ܵ=��h��W(a����>� H�Y�$��fRPy9��#�}�Sz�?�j-��De�M%$�<	�	����<��H��y��8�&nW�XlxVHYEB     400     190��(���$?�n������,T��%nb����d�G����[fv��o���uv��p-6�x)uͳH��I�+{�՞��H\�	��`63�/}=��>F�
J:�)��\�z�s��S,e$&����j �(��">D��,v?���ߢ8f��o(�^Տ)HL���Z�
��li�L�}����VE.{��BN6���>�m�`Wsh�[%�ݸZg��TD�H%ٹ�K�H1Bj��(�%�s�g�sԦBV-@Q�/w�p�'��e,�Z��`�33�T&�%(4�hi���Kʾ����4b4
��XVu��T���f4��`=�et�IK����t����Ӎ E�s�}�j%��?"�OC0*�ȧ�2a���K0gKE����4�*2V9��XlxVHYEB     400     130�$��w�L����6��A;]B���6׺��hSK���\�JݨA��T l_G$����M�e_�sj�"w3I�|;�*��?R�:�T!�4r&قP(�Ȑ|.���!��dt!�Ԙ&�
��7�M��-�<�Ҳu���\�Xd({ l�7��ҚF���v���9���>���$e�7�Ч) F�#J~:�H�0_q���5-Ӊ�z��F���N�w���{����$����F^M�(�3��z%X{xkP#�����Y�2���ݩ,��D93CYX�gR�L��p���LǣS��:���"TB�p�XlxVHYEB     400     150<��!��� b"�����`^1�kgtw���ҋ1���NB{�㏫�	�zq��߰��1�\��s,S�>��v$�u�Ǫg��_��F��^����NbDS��UP�m������8�=�k��k�Yb��e�'=�fyF/��D��Jb�N�'�hS��*�b�Ѣ8X;���p���W+>5���?�䚡n�~3�`��G�I���18�[�)-��T[��tZ)B��ͬ%������P�ul�ńcjv�k���ZE��(���]:�2� �v�v���9Eu��+�5�O�ˆ���#��$������T���\�[pR����B�͠�(��e���&�Z�XlxVHYEB     400     1b0����MtDH�z/˙-�N��%h?X��zɜ�+�% ?b�ײ��K��<BJ5�=�J���
�m;�iDq���x�Lϴf�#Ң�pj:����Y�m��	��a�{�>e�W�I�H ���{�4��=w�{��]p�Eq�4p��OWE]����4l���80S��m)	��L������0�� �5'���vFS�mٔ���mٍF�p���Ԉ���Qw���T�C�E�)�_�i��J���/�wq�H�0��OV]`}r� /_Q���.�T��_�� ��g��9�X����0�[�N�C�w�mb��x:#U�6[ ������T�Y�"������Ґb��L�1�eK�UVl�ks6��s�/��]����g��u�(�ł��b�џ{%��hh�ۥ�@)�����=c���q�xz�j���XlxVHYEB     400     1b0ѭ�x�#�#X�p���+������x����:��w%,��7�j�'ݶ�I�V��b�a�d�(|�c)����m���q�g���n�w%��7����8ܴ�6��q:ކ�Ȯ̓�1�Le��ű�G�ٴV^�^�9o ������{_��N���a����Ҩ7�%�4�;�H��G�~��۠DBm0�e$��\��1�ρ���-ܭ�{���Z��VW�e�7)��滼'��R�W!�Ȟ��!0�IvxӰ��a��O�A{���&3]��VV1L(P��1��mJy�Z3cN��������KU~�.�����hj�s��t�&��o�n~N'Q�q�۟��"��Zjiƙ�{s��*
���f�s[ �w���{g��^~�;3V#�5Yz�\;F��Ps��q�����@h���S�{fn\6����rX�����M�L��XlxVHYEB     400     170���w��lk`K�CW�[�&��c��S�ϑ5�w���A�|�X�a�Y�u�����v�]a^�>��ad�9ȍs�[ �_f�B3�W�ϻ�mA3hV�+��^y�翮cR�y��
y��ݙ����B
�)��14:A�L�pIv�nZ,%�P��M#0��l�%H��-Q[^��'mr����
��+��95q���ƍ�`��(P�x4ڈnFҹ�-�3YX�������:��W�"d������
F�w ���G�n���/���Z�[���=SZ�?�Hpeh�,��K�t�������>؅su�&��7"b�`u4[�)E���_~ܿ-g���
�X�,ǂ����dT=��4XlxVHYEB     400     1f0�	ѷn3�L_�Ӗ$8(�sm��9�ؒ�*���#�*�X�Ty�k�:2����\w
�JǪ[�~�q�s���3�8<gJ��՗)��!��-���v̶,��W� <��>W��{[�E{�T��i$��F���}���I�4�kAhu�Q�C�=���V�ɃG���ɋ.U�iK*�v�:Lh%��i����}]!���Un�Hv��F���)̬Q/��_�{���sx/�֙��X${��]�o����qI!�
^��lCy����xC/���jI�;AC	�2N�t�K����Pq�D4��S
�B��;b�'D��ƻ����a,�'�[�N�k�7v���3X�p��0vw�Ɔ��6-ȥ�<��Sm0�J=3�`�ϱ1�˴vC�/f��u�뗦���r݌ާ�x�J�=Vt+[cWgvm� �h�\\����H1S�8���U�Nd��˴�Es��D'�����ͷ������
��A;]XlxVHYEB     400     130�t�jƦס�"C�Bn��3�|�i��e5�Q2f���<u��m�߆����"��*���Q�$]:AUF��n�C�^����h�x ���C��B�C4f�x��7%]]��ї���ś����>��|M��}�&�׵l�d��J��\P���5��7�~D�S��MĈ� �U3r��{�o��u��"zr8�Y��]q��nK`Z%;KJ_��XIP�GX����y�J�zvJMh���y;��L��M��y`�3���ӡ�=L����3���{g��,�Xȥ���j/����=��*���u=Ě>HXlxVHYEB     400     190�NHY�@�:�/Y��~�� Uѽ�v6�l�gϱF�9���8�&�u~�B���7��vW%-e���	ߡ�%�)'�)|k|䖅�rr����=h�Y�ݯ䰇��4R��ݹ��o�����['�>E����J��,%ａ���r����vڮ�w����>����LQ"1��vb�Rg/)���V�T,hu˅ǌ&��*K	��tA��v������C�!�R����o0�k\q*Ŗ���F'��6�y�g����uėG)�P!<�vQ����L���jt��]�wњ�>�E����U�|����g��U�J�N�ٵ1w�v#jU�'ܵ}497=�%F~7	��<yHh����tg��6r�@�߫���Ydl�?��ss�k��XlxVHYEB     400     190��O
z��p {���yx���'��"�v���3|bo�P����W��{{=��%o~LWz�T�d��2�`�P�\/�y�\BHT��vj���	�5yd}Gw�0p.�Y���@_~WW�L"�Nm�<�L�^�z��ųE�3q�fx#�,}�©�m��^�46�3��'��Kޖ%�o�d]��φ�:@@��*��!����a`�*Z8C��	�En(�M ���8��)I��bu���U�4�
5�G�K��P	1�9�m���}!%� ��S����3"�{�x]�x�X�	L���j��5D=rz��.�4��9��6HU'��byF�;�D��됻�۴d���������$��san.�x�<��z��i�`g$(���qv�ya����]G ��9����3XlxVHYEB     400     120z ��QځCj����<s�ݚYq��"���1�Xw��1�G�5$�XYWC�"�R�}Zp�DB6����t<��N�F�Dقe��a�U�~
Hлrzf9���j�|kuW~��>����Ӷ��{ou�}A�`:DW�Q�2TN�v7��bNE��1�-.����2c�_�,8#1���q{���/A�2�vF6��jl^�]	[� �t��f^�9�K16f��a^fː�R�۶n=|Ur�꿗sQ���;�J� "�Uj3L�� �S��(�Cm�Lf3Ď�;Q�u�A:XlxVHYEB     400     170���o��`Rm��C�q��6��.o�Z5�IU��V�OrV�t�U/_
�����ı���+Y�!�������+�&��P}�����]a:�c��!QH�_4do�|��b�_V_i����k�H���ݟ�����\�� ��@�GL��U���d-�M�-��R��x˴��Q�#?�K(��PĚx��Ȋ@��oe.5p��8me����)���I�IP�4v1�0�P�_�O+Ĉ.��.?m���2��G����iˀ��o����P�_�)�ԟ���k��tM�8x� ~>)l�K��<�Y���ͭ��C����1������,�!9]is��2�7tg>\`E�V���_ʜ13i<���v��P�XlxVHYEB     400     170��Y2��E��ߏ�m�/o�� T��Þys�%�ɳ��X��`2��`�9�_`G����s�I�1�ȝ���� �@�L5P�/v��т��䒏BpN
c��P��T=zW��&;m�u�=��3JTf�&/�Ms�|IB�+5p��O�X���
�S�m�1h���|��$��,1lb��).���=w�A`G!�m����?,�w��l���Zt+��E%���%GVS�~����Ӥ��{(��>�˲��~��R^�4��#�xq��wB#�/����.���:��`�&ղY�l*��Ci����8b���_��awS"H��҉[c��\4�}�l�s�F�����s�R�ǿ�bЂ��/o~���XlxVHYEB     400     180��߲g����Ui���.��+I��t3gɌ��p}C��1�h8ft�G�~����v���ʋ������u.��P}xT*�ծ{�.i�+S�ƼF��@�[V�G�Zq��-�"��X�T	]K�>�K����5��3�)�&d�sewi�8��ƛ� 4���@���h�i�d�z��r���9��S]��ɕ��w���y(�b�fV��DE�_�L�ZC;z��b-?���۴S��R�^���&L�Cr��2r�4�:c��"&[�셤���z�4S��Fl���о���-l�>���b;�̲q����[����������'��1K�#�Y�|�\�p���uu7ej�,/7�V ��^ah��9t24�ʼ�XlxVHYEB     400     100�&��"LBF$CL�\�k1ߋ�,�ȪLG�� ��G���L����W��RCAH~A�e��$lY��z�X	c��%	q�;b���=��q���*�PD�t�ھ:��,���G��οZ���ۃ�Zĩ>x��k�����ln˼���B��KS m���X�~w�8˹��-���P�xUu���2�N\	B�r_���3βz�Ϧ;��N+��;9K\u���������f�b��&��Q��P��o[�S�Q��XlxVHYEB     400     150\��^��,ҿ;
���5h+��t��ʶS���	K�`�zn���$��d �0��=f�'YH�M~��DE�:�!�͆-�MG�M�.����Y<�$���������7[��k�tʾ�Y��H{]�:�vm��H �E�9"��	�4��#�ox��)�����|J�t��=-Y�����h����oO�ׂ%��$����Oۡ�u����&��s�<����k��"�DjZ�?�zZ�]���6�{9�n��(fl!g�E&vX��pz�#� �ɍ�E�(�w�e���W�KϝO�4��)3Z��Z�cJ9$�t� �O��R~��B�XlxVHYEB     400     150�ۏ��3v^����^�f�������D�,N18х/4�����z?����͏cT5o�J�/�4Ωb��)a�g�5kP�_���(�F,Ŝ�(8�d
sA)�͂TU��jN�����H?�_���喘(R�%���H#"�砺�����4���ȴ���	�.y),��e��9�I2tf	Lӡ��;�St�@��o.2���Z�.��]��z̧Ьv��"--�I$Z��;��\�e�7���K�U~�j��Ȑ:��&��#9𛺇'���yxܕ�7T���4Ft�?s��Y~h������Y����j�k���س�lm�v��of�Z]��/mXlxVHYEB     400     150��&K���}Q%2�K/i���D��!�N%�=�F�)F��"�4X/�&3�RU�_�i��]�����0���c���O�[��zA�Ś�#>�q-��Y�]��{�ދ}yä��i�;d�5S�`�e�?���W=�I,��OȐ�iY��TwSڽX��<OfVnI��4��t�.Vm��ӓvG�\������UsDh�UJ��r]X�BǈJm��zr��j�=�6��&r9�`��D�[LH%e�rO0���f-���c�D��[n�����M�Ey�@t������MaM�b�`ޅOVCx�wOl�k�W?��w��[���$���ƽ��C�il�\({���a��5WXlxVHYEB     400     180R�����d�;Q�iT�S��D���M=mr
�D���jY�D��.��x�rf��U������, ���]�fˎ�����5����ͽ�Z��j뗉�)�K�M^S���.�I��U��S{ј"�������J��#��X�R�Ҹ�4��]�iv�G[%���>w��Q�z'�B�>�	�����ʀ�ё���c�
�+�9�z3k#�&���O=}�*��}�q���o�?�P\�(������k�&3��on�k��:���vW6�v뛈�o�+��'׾O�����_K+>����0;�r�)�%p�}���C'�v4���}�X��m�F�5�;��T�&�=�\�OIy>�b\�^�C�3o�Uo�+�n�#K��H��Hu�m�2�7 XlxVHYEB     400     1602�w%!yoIh�����vU䂙S^_�a�)��!�M�j��sb�m���D}�fE�O8�d�]�!�����~�y@?���4�T�G"�*�r?IlT�O+����@�J�&	)�B;ɰ��:��Mv�?
�����.����G�#��Pt��25���إ�n2L��ގ�-�S� >9�z,jP�)��t�zE����ݝ�͸76���IT�Y��,�'6a��m1j���l�ʿ������#t̥��� 	2��[z���) *I��e" �f�����	M<����cpn�~��.A?e�t�E�`j����Pd�8�I���E��:u���q��XlxVHYEB     400     1a0���'�=ގ�>!ҧ��\�L����>���k�㪼h0��Fv�cHg{������A@#èM�_/�}I����J�����P�������65�4A�<�ävE��#�4��<�@/�����f��d�`��Nv�#��T��̆���4AP���];��`�2��D��R k"��"ߎ%J�95�GR����ݚ��XE��M�]�h�+��]<��б��z�a}X.���}?��2�������]~!��O�u,hX��ɑ�ČgD���{�s\�������劲�egb��M�+�����Iwjusr�L�`6�lv.�NO�pؙ��ơ��(���Na��<D5^ �ϰ�D���0��5+�������u��9���e��Hy��A]O�[��)���N��t������f�Hb��"���XlxVHYEB     400     1f0��gaޠ�:���\�Hp��$ޱ�\��'+���sP�1p�lf��"�1ѣO�[�VV��P9d���[]�V��5������xA���Nf_��	�+�{=Ne�������3	SJ�Wَ�<n�*��-��T=��x�%�#��H��)�& �Vk�]N��r�k;�+�ut_�Y��j=���������@�A�SJf��x<% ;������k�)���_w��+ע�l�����h�����zS��A�˲ O~�t��g_��fR3+Y /*z�S��q�ք�C�����\�H�6�Jt��������k���C�d'[i�tۏd��q�(0A�&|�֒\�R֒AB?��n�?�i�WN4B��!��i���Y�6sK!�f��H/&]ϳ�0(BE��&�&ân~�6x���(�K���7����)f��_eT��O��ȜĦU3Yj����P�ߎ8���+N���!�#���ۓ�k�XlxVHYEB     400     140U���K����P�=s
����=TJ&���e�K�9���׬�p50�:�O�+����:�OJ� ml�4��D�.QI|͚�v�4V�B���yAۇuCM�j?� ��T�Y�׸�p�����9o���-��jq��dј�J�nto��FcA��$� ���]��a���.��9||M=���yVY_�;�G&�C�ܙ���x���Eg��[�<��=nAa����f����Ʀ!�oO����Ar������ǏS���Գ��U�6>S���|x����2�����өm}�{��rV�2|��A"7��2ځf� ��GӬ�HDXlxVHYEB     400     140xK��Ѯ� �����)a�k�c�&�TZ��l�h����%=uip���%�~�=
���ć5�zL=���V�~�m��0���Ժ�xΊ�)�_�?X���6!�E�]D�)6��Vc�X�M���v�Ȫ�:gਅ�[����������V[,F��m��'�|c9����L��WwH����bԌTZX�,��V�cN�R�\a�z�~���B��X�R>�q�T-���⁖��ׄbq�lH�WL<�N2�ʕ%���1��9�5!7���tV%�����E �ڏ�밺O�hΩ|)R�����q�m�
�Z9XlxVHYEB     400     1e0�Ӄ���^��SIibs4���'�f��q`�qL����S��=K��8oJyȓ`np���w� �ssU}�+��q6�b�c��_���j�!����=��]�j�D�G�f�U2� ~2u��q�mQ����r6ά��_-D����]�L��JV~#�+��������j��dxl?��'9��$a=�,�(0��k��nj�"��S���_!·�Y�^��yZ�%���g84f��e���&�(i�����\��X5��k��+^:8"J.U�9���������K��Q�]뤻�en�kz���l]t��t��O�j�b�������0e�C�����5Sb��rzv��6�Z$�^����p��\_�TE�g��	��dU�ʌ̰6�Gm2��kM�1a;��b]iR��џ�F���j�\st�v��ۂ�XO����7�oSq�s�NʌyAQC��x��L��5�ǚ{20u�7�XlxVHYEB      90      90/���.��~rЌ�W�0�c��*��@�y=W�5�!������*�ǐ^J�� �G��\�Jr!�st�vz��]}�L#�݃0{Q�%`�X�?��3��C�hp�����I�R�F
_x�h�ߊ��y^�ϔ�W��Lҟ�3