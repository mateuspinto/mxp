��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l����&C�o����@X�;��}�)Vųp�mb]4�3�^�#��_��P�;�nA����Q�+�\&9��&����'i�%9��̦Ld�y��3��a#�G7��wnH��f�����>�2
�ZK�Jc�ff���t؝�>F$�b��Ո� q�G����M���D�ܜW��vS�# �����m�'4Ԁ�ϝ��9t��1fP�ʄ��Ϳ�̛�g�F J�L��;�8�Y�/֓`�B���k����D�ϋLzj���%7N+�u�ٕ�9�P�)6�c	MAv�D}��F:���{]�����F-@�<b�7[�Ur�����Q3[µ��|�÷��;��&�X�Y��d��z�t�mW��: �%S��J|�r�+��P!j|��93|]F֥p�O~98uH:���E���'8�ԏ)�OJ[����,RX�,��Ji�X��q�K���ȗ�>Mg2O��t�V���1y^�&;I�!R^e�͏��_�$�6xM�����c�SO���ō�͛w�t0���������C�G:PW!c	��l�Y '�=�2		�N�t{)"��}��#�F���O#�&���/z{�q$��|���V�T��,��Om�W�1\\Cenj��ȉAk�@t�v�|�ʾ+�Ĉ[���`���p����|U���4���4h���̬uKfWQ���*Ӣ�k~�<�:l����ܰ$��.T��r����)w�$�G� -݆�籑�μ7qR�������5�X����>P�Ǿ�5[�-��}O�<�-�B��Y�U|�X{]z�	YS��d�c��@<�W�\[t�����U�Fц�9����σ�����'	�C�҇b�L��X�I�g����ë��'��"��@�q1q�$[9��F��1��7�M/	X!�5��<S���,�a4j�Eي�������~m�a�NsD��4"/�	��C���D���v�yy��C����6)Zө��߹�CxM�Тi{�Uy�U���!�v�<b$B.h͚�M��PN��anP��
��	��?��63Zr��W��!/����o?�A�������(�i^���u��e׬�n����>�!Ӌ:Z�Ӕ�"��Q�l�zi�uU/Í�L��;�J4�.߮/Z�kOXi3�Z���'>$S'j��qJ��Ww��u����MUJF����į�m�Ui;K��'(��t�ơ�%��M��V�9�oϺ=uj�xy;�/��d�
��.g�@�!��[�,q����nA��1*\^rSs���γ�%��	칶μ���h�(Nxw�&�P�%��(L4�H��mIQ�z�}��8����*N

��^"�Ib`m�w�&�/��5�&.��l}��F��U�6��`T��&{	�����n9�*�ځp'Sg��K�W��x��ȃA�u����i� �p$��{I�Uk�U�@`�\F�͘�A���[�@�2鏃Ȍ�zmzb8�z�e��!�>瀡.w��c��b&�V%FG��łjX�I3�U��r���ĽpN	p<t�.:�7q�ƾ�r�dZ���l�f