`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
Lv6bfjcDPLCCqWZLpw5dVFBcij4d8Ovi7xax8ZaUMNlPa4ukPhvlrC4e/71ILQ8gV6EhgYtZ7r7V
1yzhdbJK55i2w1LZGztFEQCazQzVDMysjFQwxDshO46qGRBoFpSXAt3JlcUPojAEGHFuxe2vD9RL
Jzm0qHSakI3g0anJq6E8nWRWXAkQVIKfS7N0VFGYKbpJEhGIEAL4qzXBJsObC1Gh4SAOnf7/fjeA
XdrFBWkWTIKSamkN6i5FY4rQTzQsCzvmdw2nINZO8Jwbu3WoasGmRR6AiZE4ymn6Z3bYex1oZ2Vw
+0onpT1KI+ARdMcAUU6fykHyTQwGj/+LyQr1jg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="iaHN3eidZPIZpodG2/84AqPvu5TkcOMTeR4A9MmBeCc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1744)
`protect data_block
Mu4kfh0gd0AsEeO6cKyH7k0km3wDKByU91Jot9e61QKhvcJu7LfhnQgoNBQqMmD1grKkIm8ULGt8
O0xfPo1HSjo9K12N4epmn8Dg4FHJvQqJxqfGa4fZPmk2rtJqRL0W/ifhN3GY8UXmgG7WdFQT0mCx
/jupXkA3YWpBWYQX2dKc4SR/tSIxugGgHrLI/v+5fBWz/Ei0OLDbOR/9WjdKOyBe0aReK6Xl3dHC
fZS89Ju9n7it8M3rWPi7wPPPozZsuI75wBJqQHyuz0dPWiwN4RNCn9zRd+47Rj8Eow79VBf7tyXM
Owmsu5ordcrvn4pOZ+UTjhYYz89SxIKw4+OLrLy+pIaH/97KI7fTyYSMHW6NIhYhMqnpkucueYor
eX8RrcGilWhK0ADIUKc9FEkUQkZDOhn61JkeZvJJIWNUewGx+cruvCuXWxOAZVMk6GbUNOS9tXkD
8nU1kctmVW92hT2ewtQsLnb95sI3la9rif/oZsXB5jvfys0+YXwX8d+3pEGJWlNi8jwx2r02pKCs
STbm8QmaVQDRRnoepNx50DRZAhyEfpfBl9TZe8IAFMoj9xuE03r0UtlAh2mxpSYKQXUw9OOzyJKu
xtx+wK6Kxd+EBdcMDkDcuCg0Js2sx04hWLzpkuYJk5hyunYRGHdbF1fDxifGXHPokK801G6jhV34
9wrfTTKZnVrhoYU7UdVPxprgjRCoOtMEo9vt5gOU5AjGhectYp71UWsKeViBHyEshZK9m09Oix5s
k9jkShZnAADQ0JkeG0S6XvPXQLmqh9urT9WPmfg1IsoYcqw6S1e2iCWakFTIabCU6i1z2bddJbBh
fx9iRX3ff9t+pArTg8R5VdHrqnTGxztL3NoiGUxDqKedkZ8N/JITcTd6f8A8+v0AItrLKSgPB7fv
hoxqV7WDQoskyjdiLZYvaMFySF+OcR/gAUMu8qRxp/poibTxvgDE+U9LUZn9syJAWkx6kl0FRI/S
zuWhNjr/6ayPSDk8cUuX8gFzpQuYfUYeq2SATLCD437yzbD8APF8OXDEoGVLQEYXMeAUSEECBYuM
xYynMh7+Bj+mXijL627MYp7ANWZqGo2YxZspabF5ENPqbKTjOOJY8AGFKCgnBUO5F6nopBBec2/S
bma2SkBIXL8eQ6dN8I4vlH0HQjQ+90bjrwkNid0gMnMkvN5CkTMYAmWa3tt2NpRXmhZJnoBRq0Ig
SoM9L57X5JT8W1RRNyQGJMllV5Ir68aNhQddNn3hc6pQ+Y/qjrY0prfoaKoN7qLkPiY3hw2aNmJ2
ZmljUZvGaGrEo6DHu9iXqywvYxLEic9zCkD0/KdpdDc/FDnkydDUeCGhRke6NNfdhfr5aRNv1j3e
UOTOcEm6mT/jIZH5wjn0zaVriSNjgZ0xCDhSJ7HRgx+8jFXbjed5Aa8ETOEIXbJ9dByubxpGJCPD
q/o1C4dFhI42dqzntrz1q/U2MMyYBpXXYnbzAIJpSgsYjhNhKN9UIGMf9FJbwtgmXL978C9CHHyb
GIioNvT/8isZb1FTrV4/6WJ5oe1w/1JmdBjrPxqaJqHDylAwLIneVAsqWra/hPXSSVT+xHGPBnqL
cs0MasiOdhrlExVPEqV2v5F9wbAn8IqcKJrTjb98Ads7K45krXE0JEAlnnP+8dbLac/IB14N3tNk
F1FxAz7qMooZN3lyawlI6c1QoInF6dv+RD43b2+0C1Wok3eYYF4DiOD/VcJyEaBsHZ2YEpXfkrt1
9FajoupLvTGHyEEKg3byqLJZ4UYn2WBzWaF/KhiqPBJ+3Y3U6kYfsfdc7hZyrgVfPDDV8D4G4Hqu
doRLhGhas9WTKnmRaUV7B/JQiFhiK/YTf01XdNjLkvUE986eVaYSsjBbqkrMem/Tqccl2YA0z+U7
OaeHq4WoBhCJf3xTgaT16fLeFpLRm3L5nwMky9NichtirfMAvCdHhSoXnuiXzHD0WC65LGW+67Sb
+KGKj1T6nJpSH27jn4QqADn+l5+OHQzbjtOsEoNxOLFnXUbT8IakeZ5elgMTwAQ63vUYoQsMilsK
lAEG8TzJqbdEv11F08Ft89dUwSsur/8EenzwkNX+nI1lVlGVEXEgluz8N9FpadwJqAXMINYkUNEi
1LSrmHdxMg1zBit9XCcsEbXe7hxDONQGI74e7sDzqcxprjpT+peiJmfYnK68RQENknhMEPekmQr0
xELESjpt3ZOgvsFw6H+8GszuiaOcVoiAmMevwSkcZkppz70i2HTX5KHh6SYL01bAfF2XeYSN+Na4
8pzw0GxRpJBUt85QliKC6MlcEW4rtVdoLJs9OLCKDSkHxw==
`protect end_protected
