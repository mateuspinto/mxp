`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3088)
`protect data_block
H4LYIzB/V8Caf00yoV/zfDjzMWaQY4RVGqGLW2V4c2+PFK0k1UACs61ScC4H6K/JGGLJNC8KUJzw
WmPGnE9MLrncpvRs8BTFQ8khCNG06ZWqPQUIMqGNO0znEy5KBylEge5dJkxxX42OsZjfp7+TNfnJ
HpY6NHlRj4p5Iy7yUDsB6Fj6hlbtk0t2AGUvQTI60XULmdV19xLMVB6NU2JFp/0bD5yR0vPDWjg7
/9R6wg9MG13vTJlCDE+w/0PaOA80N0DXJyi8RZEcFY0775zTC4Itb/6AEGJ7iOb2D2vVECmL2YAo
RTtvjjXbMU/cGAl0qWAv0irQSf9SXv3pAqJxSz6GC46ybJC0HGHNR4Y4yEYrqB5QF5QTgzP0mTfe
h7FaOLqCGAqybtkOvc3IgfCXlTcm8YPCdiakNlsuQqG232NUzXI+SZKoV6R6WTtdkFYLlyCijgHP
fq6iQHM3DCGWSDbMVRu9ZVDWVeRTNW95jDi2nZGCY5/m22rM4Clc0pnyqBK4H9RXunDWNSigyngT
sKitjRHPq2LypzA7eIiDsn71m2VbHYjek/sjfr/fng2Y+DPbEFt7rhTdASjMvIhsf6j5lANigxU9
b19T1v8WNmGlpcJDQyeSDSnrbP2hlFWOGeysESIXtyaNE1THv1UGrgdygnyELv5ja9mNd8TC9K/r
9uJTDnQaGqCg/bla4qBkFF9XD+VorT6/l+PJfxAOQsS9VCXOZh+ZDe6dMijS7ck42RbK6tNojl4A
AKLV8H/4Mq3bQLrtzLU5obTQmVaHUfeOEfOH84wCLsOvSQ+7CeWP3YY92E1+xDsIxW3OkyetyS9Y
09Xmxu4wn9avhDu622q615lxYmzt6ESNThnNRO5c7M1xtxUW7+cd1vHphMCzqywXBJwBOF+6via7
7777ifqleoRJZs3XCByU6OY/rOPQeF+oVM+dTzRHLU3ZrSXp0phgmL0PQaiR/DbtyuVIgm45wUf2
s6V2oVY7aE3pD0Xc+qBeVHxUsWvdEWLYRQcWOq9Gu1c3WIM1bzDPqtsNzypLFEd88nAc7YPn0Ydl
6V5dqiM5WdX68PuaT8Fqc8BI2g049t7UY6e7W2yG8doSXB2GoTM1TwN5bRDCYJDS3HldiPieb5pr
zU4AAzxvTqDyBhjO0pdzAX/gyaTuThnkVUd/2SkqTPWhKxo5WsvXvanWYpqasoh7kiqJsYHyRUk9
n3pkychMh2bbT2oOrF1ml7cuQbdkt3CS8IuBvdcJ+3wReZGCEmlKrE5UWcPOqHBysE3YHH1pCQIi
O8Ev+MV4Uf7BzHDB1MwvHCbczimdVRITln1Wm/77UrsTU7+XdClw2UQmSixxqZzV6EWHgiNup5Ie
syFSylpsAoeqm8zK5GzMaRHjkJ4SJS69cpyJR59jIhciifwifu8Y0FWtKEzDSfUjFvuTzgb5tZOc
Lh/S+YF7io+rMgBDhT12r7HmAaxIUa0AI+gnArDG7B/TwD35jniRyXXCENbipEWs7T4GwedpVVRf
zHFW8hEYr6Egjs+2lu9BwerJPl6OTe2GRJB+bVFCLlYM64wmFn2QggWcUs0bStGdm2QKNi6AQZ6T
AI+UeH+jco/esteFjQW+qdTLG96J7OxjubKWGev9KeUlH6p/MsaTlOBmcatNnObntonBL45yITDj
4vyjTmSnx4paY3rrzHpCDsiIYsGCarPczAWF6EYApJGCfnlr2N1ZZi6oIynUDtF9eTSI7sfPS8eM
pN03oxXiotu6W0yJhuN/Gx25dzxoirBz8mpsk4YpP8wa69GqnhrQjFk4/cKaxnJXG44T7xfOfIyu
E2TVz+UQzjTmbdUQxaStfuIoukJBZhWJD1w12fggHT3EWMJAMlU3LurNSs1pfxuYA3bom2cGdi95
q6+chN4ILXE7PznCYtLk5VNVPgUw6mtgfK7m4fvuzHT+m+0MUYS6VSUESVoexmi0fQwGjeCGF5+k
xlbwPXGJ/PqBKdk5NmbEXRqmS7w0/5EDA7BZzIPdbvp9UB6jwLVr3cUs4dhd5NbHl4OSyFwXn0di
r92CjmF2cV31TCgT4/8Mrx/rE8lahHLcvGvUQhu9dUppFswqGYVm22clcm/502t8Ik+ZZyd6JgUa
3SCw8Y8c8OVnSQOoltTAPJiREe+oiElKSaYSseSFAU61FUEgxtayKG8aoRd5kG5w8MYBgkezFwho
0uPj7oVa05V1sFN1cCbNcOie/knq75ckJhPF+hRejLnLtkyXptEspFV0gObLrdq0xap9ghPA62qa
wrRsxDHLsvLboW55R8TsXti85fzZXQRcl8CWdqf/bm4PSit7RMaB0XifON7f7up5pJq0cInvH0R0
uK4R49SbzNzV5Jnk+pAv/rGvMtxdz84+zAcealS2Y9tt/zMn4PTococZZBEbluyWLeAmt8sfWtVJ
4LTEL7k9g/6aCN/QHLRQ9iyIQv/JjrqYhj0npO7l/pAhqO9GREOim9Mo7RI60iHssX2qZeWXKpIu
VQB1LikBOjoD7XrU2yrNaL4MUiZYDRQMyEQ2gnDAWkfF5H2vgubH3nAmjY8SlQJv31AFYWuiCG72
Umgy5diSTOFpOlF4pVQi5uBdsY8G+ji5tKiskZ0HicIp+pzmP2G36o9NBK3jc2quAk/V8alf7mLA
GkFwwycA0aWf+/8zfpN8FOqlw08LKbDLTkTAmYoo78Lh0+istJ9gkYl8ewAktg+FIB9LgeiTIGiR
PkoZZDwCqMEnWPUnh8GHNavf22/I1AjpbQMIQV1XYMtBYPtWojPqJ5JMHbmnniNMDTNicvbTPCBA
8rEqoZEMIbASjRpubZ+3rpNG8i99Yh+bMV4e7FCH9FuiulYQq1lQn/uAF7iQxfLNUWQ9LLsaF3P9
baXA1wsDSMgXYbXfQcLvTkUd0xR1SKmKhMHdfwk3chfXnrREKxcxoE9qEhjuqB2X1fQ5/Z3nPxoB
jsIJVRXH3xow7H0YM2H+/Vun/2rIIkilTXkLIWyP1WR6L64VTX889FuWqEmR7O+vVoZEfV74P0IU
/WWgTh0wcPbsZ2w0hJV37f9FcqQyy6kWtU1exLVFr7Ey21Kn9sFscGViUn3tCcdsuff1506ysEvU
WBSYpExNyFG8utEBr7oEVWRdDHbia6KaXcglU1ZG+/dHXsWTQrU74CNyNolMu2pmRu/oLpcxLWPU
+4vCyOJPbqs8kKRdCx2ekinGdm5MF/uF+b3SdAHXkAoJmx35vSzb+aKYtzPV/kXFzc56lIWyC+nB
i1FOGaBRlbmc5qT+h7AZ395/43hrz4WJMEGo+yp24FZJUHe2DFfRc6wpjFvhftHwSmUEZoV/cLTu
zzaXs0iSjcjoqWRQXz7JZPivfnJE70V+JdLxsuYIylscRIuqGKnnnvVLFmB0R3/Kk4Q0GE8WILi2
AEMZXphKc+XOZ5FNRKzU/qGmYJ8jI3JbBgF39TIXBGGhq5AAwdkjoyO/vxPZr8fYt14uX3G9TrVf
wWoa7SOjpYT18xU8fTgPTJNmLo09sVkwL89pwTBHRM8xKFy1mPQJYzFzlhbjk9mL2NJjHVImrgKy
qVDV3AG8LmUSevgIVnLxmz/XBoulqkT0VNjMUkdFFWYmc005ORyxwUoI+JDxG2gKiokPzKHZO01A
230CTCpNjdjz5P3IIhoGLuesmh0fEuXY26WY7SEqMycKN+E8OpaKa2mHD012NtbH7j9tzqJAgQtv
2Vs+X2xY5r5fbpPIiYsJLrF7bR8V2VKUhvpVZL26VWdsSdUlW3L8yEUn5bx4EVMdDqMoxWNlGxvi
jGbrKdYNtEXsqj6ud8hObHJ6A2FXbDZD7v+AyS8rF4gySw6p/VuGe66xz5lESejAkI8Jh8Ty0VKO
Z5jER64JeeAlAPk/xAptW8e+eODoPnZ8IrBm3CNpUMa64zk1gb1c460S7gpuV8tXs+JndI1LICk4
chH0LLl1KPiWszOM2xERUVTkc0VV4CMPzAZ172TX04jtFkemD6H8mReblB0KhRhKOfx4YrJ4x9cU
EFoDok64w68bUA7dr0cW3ZvZhMbksd0D64M/6rFjUiIVDYaNCfH7+RbgefHWkYrP2hCRqVDOofxA
bmpppfojvkaUNg==
`protect end_protected
