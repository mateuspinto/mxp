`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
NuhkYqA3F+plgc8vHxA3WfBX6jWMK+5NMDSJ/VV5AXS9NkxUBMssLVL9pZ8u6TaAuJtpoxt3uEka
4NbT2j4WxDd7v2Wy5Vtj19wllcmjcjjbY8iLY2XVAYHi1EwHnuYe7OPU+LhP9mNuLYjw8H842dZO
qlHUWV5sko1N9zBKxZvMIez4Z2/TXJS1fqcByzkdcdLqfFLskZmKwhpwZcfIRs1UX8O/CMc865UF
WNYE4RaWMIUjfNVlrGn3gyBdf8akkizCF2jqUtlXTYEdkGaSz/1FCBjBCtyMDdK9oqXDGwIHrlxT
Wmo5Lra4FAVsa5uFIjfYlN6g0lc4+kkDS3PPfg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="nAtTK/PoqGZZJivJppOdDqLHLl0ZPImzWpSlorpGl8o="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20112)
`protect data_block
0MkcgvgmOTyhEU6+0KRGHaA43HZ4Vc/nezbwbvjVWMo3yhv4ZGBYBB/ojDD29Q/mEeYqqOtWqovL
F+CqC7DGZ56+1nZTYs+Qj0eZqwtFB8EKQjis3eOWHW5rvumeqDfUspeyXXe3WwGlM0M3xswj7uep
k7ex0s5EFwnd1Vg2BzOVRaGc83UdBH6qc04K63a8VG9OLKpvT66OpY/+eG6qt+VT7rVO73IrJx6T
B3hQ7204Zwl/37tFPXfO/LJAJKvujp/GGqUdivlTPjf5mFDl+bXTUJwG3Iy58mhPl3yN6V2Ck8B5
MiuaZYMzucP3KriKlRKurZFURe/iRGHqDwQYBQlcu47eXc2Mx+glzGzE/sfA3020nZcnQxy+lOpu
Bo0024T4GLvRZX+8NGiC5pKA15yW/EZRWentSXf9Sge8G1TrnLSH7vUBiy1sxoPFGCQrhtLshZuz
1g+hviRoo3X9trgincMG3G2k5jRr5tjV3nZEzzieWBHrhsBbyf788Kq7uvFr5ZLb1q2dxKvRqF7g
Ko/OQ/OpwTsHxBhfKcCUF2eOuXGlV+K1vyAVtLjFGZIF/gjSU/Uw2fAbsk+BXNvqZRyDh5VvkxWq
Hlm/zKO1c6PHSNdGiHud5CBRR0ybDzeRH/q5hnfd3IaVp+hxxQYQ8S9JMk/8GkZlZtk1iLlQPTS8
rj3zrcUqRJnovVg6lE6lUk8h4AIMkEGU991Gsc3+tbLLDvyUxlHYqlyXXgu/FQ8dRPvsZuYE0zYk
5+cbExGWHo9FEAKe3yQNAg6JT9HgihGjHl5VdkjZOWpVcvMv5qPG1JLDtb5L39ffEbNnHaDcwxM4
vEnFmOf7Vuojo9GcXsF4xM8aN+HI/abf7WlNKUTEevkNEGXkp7pfu3eMNM2ajDlejqKEqiaEWfnN
V3dpNYsIRFCFNQ38nlkMooD0envktmN0ZVd8TNMY11N7Vy2MVad1t45N5Qgl3nDyMpk2Itxw6X+9
atvdnEFGDuE0IuztNXozypkryLDU0Ym7B+YOzD+GMZngK4ey6myOO3Gr5yNnhVZVDIDUYf/wND0m
SIiMfP9SdIYyb8ZnSDMAk/50dX6Vr6ue80byN6R/PV/+h9afNdcsMbwwMwUuklLJKDrchoTHHqgY
Z+cav6F9kq30zGQxmtR/Joca02BFwMo+hXDXGYWHYhFW16nBRc0pxQc1WW6SfHtViY9CpHzemV16
4zjhpfu8SuvvlMPtk7L3uFMtLtjqz2sZfAC7MWnoV3OBkEWnbY1R9OP9vVyAzu2fueiJzA+Mb1mP
6NlXyB/XkS3UaHHb1g1swR/96k9ujrJDRC0pPc8QK/u+v+exwwYWRp98pDSBgHb1/Pba+VdlvgzB
kpm9hsjcajfvmkdyzF3+U/4XXROQ8SayBrQrAtht1bYZj7BmPPupzCQAFnC/jNo7MLBGbMDxFNGk
3Lg8pUGmM3KzeVLCe+hKqf4A2idL9UYBV9E4jmtjm0NfeKzgUCsXty/PUC2ogv5hCC20LbxMTtIm
caq4jyz9hzItWYmTHSiYdgGqlTaxkpVUMTeoxawauEgPdmt+ekflhoC0zbWEJYhgYVPN8zr5piVw
8unlgl44/YnlHuOy0ngVZ3EvHsZImE5YGP8H/pw8Tn8kUk3UN4DUm32D6kSyUSdRJ39vgURdx3qX
kCA21b4/RDcQYXMrHUXtRXHRVPLpuHWduzjDpl8CdbLUu3t2FtG5ydlD2DHMF+M1/A2Gq/MakZUk
dFvJYbNjnR0ZGOuQc9i6T1mH+8/fdFRrxwOXUfn18o13dxoxU3zz0YHY+LB3ucWi07EeLk9Gl7a1
Z0U897Tq5NZPZeXmkCGgD6arXddL3wSbaYNpVJeQdbP/wP4xBOyb7WSx7UW5KY9KFn1y3pffmhPq
6/QfsIocC3LKh5extb5+Tf+92lpIaIj/KCeg0mG//YxLjDGynk/9IEGkYXlh6lJi29IMgcC2Get8
oNQ3JdVVrtZw7xRyQGQ9H0/KvFkykeizeEKlwe9E6Ad6jqzuqR2p8YpG4CWt1jc/dd4w+5Z5Yzdx
WiuF8dytxciyJB7AY4Xe8DPnfrGfu8UKdOyfTrHQ4Ji4lQwAlOoL45OzsjQl8FszCWuyKLf/cBhc
YDk+xVl/0+vchF0cU0HIs5GMHIMiDEU1rjOR6GDj2jcmLKePRho1GmPyoot/wKXnBwl9uknXJjMe
2rHSzT3MasBlbVlHVPKmGWz+YSsGeWuKhvNYdD12zWvpjc+8nSWpPEis+NOHmSgf08y1tC7CQyxh
5Jfbl7pe8qvcs8LCMyJigHy5hioki6kA/guuDwOrK/E+rEJuDR0woFRdOoFk1kQ1ortj3dQp9hCY
EebNh7VUUEdKieVtqAqGQphAUMDPkaxfdCTT9pWrWXAD8nl8x8rWoux5F8NGDKN5iuUCqhlgW2TI
ivpiSNFjM//aBdUE36Co7oFQQ1jfOItew/gIIsWEgrM1/PKpv8YujKKdCEyh1mMDYiMDlZYSeHLt
HtggWrwu7IGAFSkad8ZdGFiS5H5PDsMUrHXWp3AayNg96el4aQzyeJ62nNnvLHUsyfNdCz4yFmXY
wr1JBY4Dufdoj9ciNv65ToJf/kVMrLcfH0z7VKFU0nrWhEFPzGhfwBpPyTEWn0tpKOMC2OxKRJ7n
MstIl0kq+U1AQpsxm+TrMqn7qLTx03LGnEshimi2zhBRA8sjeaLHM1ONOE4RvnHQe+OqOTD1z/Ub
CzU6C237CiHPn5sZlF0CeUW3yYSeFbZacezi+RfgEqORq2NpDv0QbDfTmEbmhVK9dVOafEocCDyl
22ebeGr6FPWOql6Nbj1bIrV/WbRww/eH0Hrp08j2HMuD/rEver7+mEdpUI0mTC0bUKtZiwmjVzck
8vvJvB+uTW9rlP8V1hoS50eY3iPvvFwLNrcGDWPyPC75GHUPSw0q0VMQLp5ZpJbwe8d7UNBFI97Y
FIiAQ+2UYZmjdp8hMDZVWPWXjoy/ndYv/y9Qo3jFQjbL8s5508hzXBCS9Bklf8sNVKV1xyw5aXq3
qGtWb9vLbs+L/EvhpTUyv4IUMG/sXxk+yg18Bymplk7TZxVDX73ROSOFQvaUJELH4PXJVvJ2WV7F
+bSZ99hvWLuDrY9npwcI7PhqTH9VwR9+S0sNMbjAvGzJHiKzvG6z9BYHOEF8loN5QcfUmh6f/pGM
JiqcYTIOyh31bGTuKXn2YUUxx/3RvH3ka6vZppowzv+Q9xmdLwn9vAUdmdjSwoe417dpYHjjJfcG
j6EMBEH+l2IovXjPuzTIK4UcsWhHcJS0YVQeWKuGchSIk1CrqM2DoKoBhV8K8q7fMglDaxhnc77D
NuKFFPmMeoxDoKMkBArf5gWNFK7KVuHDn2iDt4RGwFEUoallkA70pF0qe90A3W6ztNnjB1w6bStl
fNU97oK2IP/RO3LU8Ft61x54kuvQBJQ95oroPbZMXPs29s0NbeNXM/0LiE5bz1BWeJ+1P/7OSSW8
TTIw65G9O6KCLJsnNkZykZoiXfM4L8ifPQdZY89Ep0/8PO4dxtKh9Q7QXn8XDjtBQBFAHoWZYWJA
itutHMpWrP8KmHqa/z71R9ZygMPa8bguO8bJeEPHuiglI4j4ahoJYUBOpNQefITr+erjjyLGVPRy
SdZeMSWX3ZlbGcJN0zaZyVP/HJuUhJc7ZLk0L63oqiY5XiYNnwg1K/T6QmFgTL7WKan2YI551Mix
ePYOPBw1NRShiok9WWoqW3t1lohBP9cqpA/Jlpt2Wu9q4xd/3xTLyEZ6ahVK4ayJuV3+PIKe2bAU
bPCPeqkrPGmsLAsds6lH+Nl3tHXwt4X2MmZOpZ/KcV9FRONuG+kYiJyyPNUesUUhslmepyPolcvQ
iB6DLCZR+zRKgGQCm6Ll0aSNL6oeVyUSzWhzqUGK7On9j/wc41KGxxMtvkzkRoBSjjCrKOzMi8+B
QztGrMdfzPV1+jdJYonSo8DNJ0S7n0ldsoiOFFx4DLOlRrjn/NsMvrtnIktrHmCNMszAvn9qep0h
9rb/jyihfuEYzdO6fM8uRuN541Q0iMWWm6JrdSYe+jHRKsn2Gq4p/hQZ/K8P1Sm82Oktjcpf6aLm
3FhsWBLFu7cVrfCP84SXIIz0axs8UDnYP8pCeQ99RRHh8ySaH2lZuUPitASwBI9ieTl46g5aRbMm
Ai1Ax71fnZyqbqTWUxfZNOIN3k3Z7/0FEu6trprJ2pK4q8ZYdOndUxmNPNjZN25ZeTGgCWyeOB5G
hy30CYTXfANw+is6NnnpKlJdeVhFk7/MhrJmpxhCLVgmfo0LkzvT+CaKywhU2QVRm1STXBXJFsjG
YKUiT5sr4kAfuG2RZop+lb3Anz7jWQJy4DefANzljpbDsIicVBzYyWawWOiVoacUNnG8YdmTGJRu
zfHVTINDbfUnnqDDJkh10TX4NV9xxS5xpb93CftQPbfAaSR5+tr3Pa8vHUnX52WhhrqhEGMwXRP6
nHMUx8PItFK4RctDHoyzqqSpMXHB0KHqDZ26Qp1Cgw0KMnTzZVVNK/t2QPucvU+U9o6CpDpVtKbz
HNzmMF5f206Nlr+uc2r1lMaFPwUp+f28zygDUKatN8gF3uPDFNr29bEyMkkqNYFk50Vnuz+fO+Zi
5Vn0hDroc1Z2Jz7gjSqDZ4FuovVILCcwSjbmHbUPADAjKZCm/Sif7y4RoC083D+3VtHxU9eMLtfS
NQUpI7SyfVxyxMDbkE1JjPq2Hc4VMn+hyJYU9NLSwZLCGn4fOM4zvye98jLiv4HN6XPKUQJuFgsp
p0wS7CRLP3xJsMZGfmxI9x7uWury/N58vPgAvV0KDSEXO+IfwWgBASTT4vY7TLBOdc6aOrD3LWr4
yeedV648Gc1ZjJlFMbwq88xB91d00+5P/NvMyerNQs16rPnKGFWomJo0dJgjk8rXPhGEct1VKJzX
1Ktk/t3vDF7Rvac+faS+DtSMIvgBpnpPFPx52sweqWQVNa+UUNFciEvgX5yPupCZ3fmbvyQUwqCI
uuqXA0XVuoFi+UngnApX0ixylNHWAvHQUUcyEapf/et3zKWzo5BNRVeABT+7yPW7Tbff04pyGJHE
kgejrCEmGhP5SsEFZSmp4YyKK4xtFqb2S7NuznQJRoNZbvayU2Gns2QEos1zIkh9NF03PR4EdHQZ
yWfPacl2cjuirhg/lqfIgutk4SqEitut8A6JFp23YoCxBQtuT22+cKiIhtPif5FEtwEAhS9wdZ5W
N3PgI4mm/Ha+XLJkZjGQ9E3t7oiYArr0uUGCUIKTgafQrWu2MJGXFtgiJGCCfmzy8PIVW4SH/Axr
C569k2XlQ6BU6NORKyBxahtxo7iy30csG7ceJ7hM0zbR5IByt9w15ltdNsy4j/VZ4htibsM9/3i3
Xg0Y9LSkTZ0cTQZ11T2f5HIuhzwnzleTlkqSqWQrmi6Zilspx1ndTbou91iKadVq+eda0SDBI2RR
iZyn/QWxRybww/MRkfjD954k4LO6zw0JEmslpgHWpJ1uyK+5fXETl1t8q3PR0ddyECx5gu9JjBUk
LZk//8P+g5fm828C+tJeAlFyYiCJ2DMeF6hGpf+74U7PQm6QUgOX5mtLroOwPi6uaoCAJZddSUSw
UBB3ydlFmWJM+wP6iuuSwvDSKP9NlwL1kT+bop2Vyy35k/zdPmdcHZgGyjI+yKDWfdvKApXvfISc
D6RI/XQX2Bdc0qhmOsV7olTYAjjzEjGuNaoMiLvyd8qSj4DfaZwslcrSF9iNmBbfG8qt/UKpkQVV
9SXYS86XQiAKgUTWPjS68L/LNikk4mOucM6trBVMYIt6QhnOsnWfWSEBrY49K0RUNcyjVWAzYQGe
3hJP/v/m4khNiShh+MUsq6YzO8IfKcHdlYyj0lgyNnOVEkxovahhm7QAhr7V0xMfEaCrvcAafWoV
cbv3lp76vfV6xtW3ClFOLVudf4xpCpENgQMJg30DTJkKX5GyoppLvNf1HCbY+hcUFZNWtUe267sL
cOhLo5HKCBbXfQaNfL4ds0+BRYgCDu2FEMy+Bf+LGIxUHrI7steFhdaF/BufbB8MdogABTV6Bb6X
k7cBNkZAgXA6E5k1TbCQP+XFz/NUFJS2D4deDQsRYCdT7sh6Kf31SjlL7qcbZNvFhFGg0JH4b5pR
vK/Nmo9nRw9/13TZy+amy4F+IWwMm0Rmx6WpggJjq6YAK9RlqKLHpFwYxIFh1oq0wYfd2mnzxyOV
0QvyW2Xzp7bT8aWx2I2nAijtlWSmPJsFGp+Ud/EUmUYpP91QCw+vvlWRCK7J91vP+AkVIRr4l8fg
rcHpDLtge2jb2pt+S8jcSgOWBhKYto2bMEaigbQpNiVAZ8wH3aDnNapNyDScxMq3bCbEMRirMv/1
+SD1AD/pD6KVwEx8pdEBkSyzrfTk/VZZN9jGdm4/PAkBYfQcGQF7Yo8gSPt0TjUJECcrBnnNcegg
CpfMmbDRh/A6r24kWhPy5y/BaZatvCKY7FQX5UJY7Pdt5yL18d/ntunXUqJBU+QmMT1gc6Adld5p
OIjDXQHBvO0YDvaG8nALs5mP/3i5pwf6k+TTPvzeKISD5rlbkOhrie1U7odT6WyBSs/hnoiR4BZ5
8NEfdwU9x4U9ug0yd0pNjtpWcRhh4yNPfTxDHSujkH0GNojTw21usUG6GYKnJwBEBEZWY7IQUs8y
n4UK3d8AL3mCcQ8F3xM3/iRtVqX9+l94/J2xEZ2rVNRmslQNDkmel99kZ71x3Di067knqYQVvJhQ
CY1N3Jz0h0m+PKD0esp95mpOS+NIRl8BiTeXL7xricNP9CWJFsQg3m1VtakCz3iyT9kGGlffypjt
4HwMA5xDkckMZ9dupRAhGVyHgHkNK3Xn4ZYY3OqBZmCN/oiVK53kTxRzo5h3GG3R5TQX56d4KAIi
I8YBkbXCQ7fJ58AdBE/ktwmy7px4jSSs9fkQeIGgMtdM3XZkhD7IBjLV6XHk7JLxx4i3w9yF0E2m
qpaN1eUqXYKwTr/YsHhVs6zX+DXT6m63X5hoXhwwjgfiCvtTJP2g3xnqRHgxni+Y0Wgp0jTbVMXi
Hi64izpQMJQCUrIsmLIHu8//IUohILBrX0GkTpC7WjpFzhZnCsSVAYo5Fru3pbpauXq0tFtF1k2e
5vJt0dpKo8xoDhdbAeD4DD/NTuu6cRDXLnCeRtq0MFdVuCvg7Dv6XkuTBehcby0uxJ/5gA9q1Pk7
G1m9kfc1yOJz1agllGpNoMJ+qg1FsFjSldjMrouNHfIxu5AxS7QnBKzkiyUrmaRuyHXUA/cPmHZC
0Z44HcHZsipZRHLyDHc3g9MuZXfEOgqRvhO0e1UXg5yDwDz1F2BqIUxdPQWHXQ2bUIKauwznkUWd
e2qG6zgzia6RdMIStO9jUZQNNCbHWE+p5x0ILS0D62aMze4WSNZGwR5o+nlWFKq6uUTGnNskauKz
69WcpuJoB0bNxfl+VQTUGFt0DWROc07v5MbURdviLaUHD1AsRixhceAOGPeYG8WHB6hhuz2/lMIa
yrH2S2nwxJfSUIxQxVX86rfOIAvEmGMOZHluDqzGF1UTlOm/r/Ytc2mtsErxpj5VerRMSFgZzVvt
dRguJJOTtMoW/ZxAqXLIga6ZTpdCErd9P7Id8tpHZcjbzpi9kyzP6LkQ5lfRZzsbyNAr+q0BEg16
JGKw3U6IvwS7gMm3U2G9yQgeCWgDs9Bf2d6Y0SlMoaVOBqs2xwGRKeN86ixqp+EgvcHUVpOoDchY
fsy0im89Z1IdFtjlDnjabMSZJIggvAN487eogkU1Sas8ZXLypQ+PGSFVrzCOu4pepyzF+WlwOrS0
9gJ2uNYUqkA4z9jXYBEpbqUIcbPBXK5M7ZalIUY/1r7PXTPm4RX/ehlypKsre+k3Jw5OE4YgHNNu
i6bRwVkQzQyS8aJpk33y2zDY9IgFyPP1oAQ/woost1RXtct8PjNh5QMi9+XGOo2LhaeiCQHlGVcN
zSSmGO45rTBzy/+N9ScQvw2UFcj0TzTXmD+PdsHk6IO8yzK4XCdqC5gh5RK7EGaD/F8jIRrfGYg5
aleiwI7bUfbLJfoTKef7nSirEzK/RoUtVnw/GRe+0Bl3wbP95SqYUk2GvfwgBzoqlTFJbI9me7Ko
gNkOXcXq2uNiqVAvX6mfiEREKGDfV4pXAdgwzmze73NBLCt6ETUFdYCD/Tb+lC/A3/u1vcMh6+Sq
zc4JBjtwSbWxCAfm/pHNcdinw/Rv4MD5qfl72UlCeXtFqBEwVGpi5puIXHjXyKNPjQDTgE5+Qc+g
q1AKW77ykvxYOe/xoKoY9gINTrf1/Oi+fa3VPxIMSrtSUSnBt8HR8QCSrA+2JIhhlsr07rZqLybM
XsPTbXkU6Ddlb5cZoxP2dJrsr+/+4+W6iy3+d6LeXwScxoSSHHI2nSUeRAHMCwTvg151E3FnLUXQ
bSsAxx8iORbZ8kXDnqYwdTNM/M6scOai9EWY0g6pKkQrYQEaLHBmul71+/MZBQ/iw5rjOWRfbpPM
RqzDx+R/1uDxMqt2czkKmzuPSljihqPOcgo+Ccd6YYu7LYhA9xqkz/fBop2nlXhmJZiM5A0r8/MZ
IPUyQnbUfWTulYqvt2jwXXcMYhiis61DjYJcKZMGk0W8ge3ijEsqlWvwkNTVKFgvi9pXuvXTkiMJ
08+zMfjvAZtB/1OPL5IXBTzJK8akFTB6MMn3O8BaSlnIgRBwWSLnVs7qZFDk/MZRgi4x5RYvjHK0
b+xgzVrrVrFIfQRXmjHGnZ4AByGFyYs0LmkJOlXKiTzBIQuXSb6iNBj7rqjZYGu3lE1ZPdSihIFM
/D5DUBy5nGZHv0SjlT/X+BfFpMo+/GYGcCVzqDw6BPF60dA3GakhEsS9NBADi+M9sgzTNKLmltE4
Y1Sbo2Obw4VyD4fb+/kgKGBCCl9Q5/s13N5kCkzJqoPOWaDWFcFKeIyRdop7yLCaSa5WRYkrwtjV
lqIJZ78prD6jiT+Mmb8uMlyKAuySSy8LkoerJntWEZlQo4SX8kmagbA6RZUuZLePT+5bTppGX72F
FL3QXGFCTpnoxB3wAihKWDFJDUjeZ/yKFquef8f2jTm1x1cGfzxp0MW8WPVNOlEXozkkRFPxcsMA
pBtOsywZa+7G2qDKdvfVQ9RSU7RK+2Xb3VzoZhd3N2wXZeLkfVXxCJeu4puHnOEeqfCc6BVh6lDf
QvWazgVirl+jzFkDh2wjNoMg7wrz8G0ZPSB4t6KmQDPTb243aM23kwZ1BD05LZItsNReHVdHdA8y
+8WMcxAKERnPKMWjOtJ6wCdiV/gl+PQS2ZAqqOdTFtTF003s4YYfVMOQ+183wezRJ7asz85srUQg
b3NpaQLrG7moqOkb4sXxqiJ/1T4I36voW4p9FN/j1fOUb6X0tg+sjpnK3kiVgFmEvxycONvJ44B/
MlHQ78Frtm8cyYuWb/JCbwC4v43SaS9AHDLNVGzHNhg0+SrfVOnaKdfuSOTTYnL0XxWTMwD9yjOg
Om853LmbxbmIbqYz5B2eYUha8q6vGpxA/LKWTF4yhKsr8WrVk0l6B0MVwfwuGDSwLUlu8cbxZTQl
QcfBOv7vjxc5UU3V2TgYoLpx7gOLCIIX8uvTevtKEHLfrahO55MjrGxCzYNBPVnKTE8BYWsFWe8x
MompvRuavAZZqd79GnttrSpEFMHoPcE58uSOkK7q05uVGG4stWI00koPjAsGSxVXQxIBn1BYoAEz
pHmA0rU3Goqgl5cGiOuzs8a+ETRln6vh+Ku66KWiiqiJhyTCxksbch+hopPXoUIeLWKRG5OD+bg3
cllQGPEX9Cu2qUj/25lr7+Ak9UhVVEkukKOkHT8JSrnhv1R2Qc2jsurE5KwjmBfMrRJpCwv5zEdz
BP+LNwAspNYOnkjELlSzYKVH7zbsXNBCZrbuGaONEtXbiVNnBIHrEteTdbT7WmpqMXQWfKKzPWCc
QoFbabk98bnVJzf+cAsMgwJ6H6tFJDNZ13/QJDpd+K08rdG632VZYgIJlluPyjtWpqaCMZfB32WG
g6p5U+vZRq6lQue3M44rgHZBj8hb2uep/PtmWYvKjjm8T9+qFBmZPzPS3ad4U2XxtxOmVhUgTxhh
33lM72NNdx+6S8NcB9MvW/paVp2SU+mT7mKxfZKeGKxobwbCN4vkgVgPzoltTZuuweGYrGCmB7ty
gAs6wdwh2DXVoM/nmtS1r1EGEZ2C96XM95SsovEMOe0VlWUF4NoR2ubXnV0O/2CVrss0PqHjG7rx
DV3o7MqCUbhHCR19Naaj7HMSIgjbd0XTygIquHdxblw+0pN0YSas60UnQYxhd7jkYWY5B4XG68T0
JFMnTDOJ+4gI72UI0y+1RS6cNcVNFMdd17rwE9ETirxwpI9BVwt7Pr2t1vumDGLmQq5dXl9e+vAX
4pLAdExhKkNRSCvs8as8mtvqjLokdt169BGqwH3ZOROG5gy35iQRRYy3RDNfwtMPbAeCBOWJeIxR
yLEtZhF9E6yPcYVMUiKa6NhIGbt+/h9H1yH1s7G2z7bFbsp0EQ7pdYotqCIX8/S+IsA6I68umgkQ
kxkefiYSMAe4acKybC25scd9WftioO6zv/9TB2yhlB+YghLvRcYIDlV121wgaM5P/qfdMrH7/V/E
KYAt/w58MVILJPYHUT2pwy1WG8CuUYlife/9EhQWYrSCq7eMCcm2RXA85ZFezF7rjITZJ7uooXxK
qKiz8BycV0Y8dqA3rCWtg+P0+mMszoD5LYJuFqRp7X6EmKJWEjQ9y5UffGt7c4bVoM/5NAHlmk+L
0X2w25NXL4uGM/zAyUcFK4qwmY8MUg74f+k5sbxIp2kVjqRoWHMGnpwxDVz9HkuQF/Kq/imj7tkd
FAw61rTUdagLNs2uil42HD//xRMn3N2phOMV/CE++AtGuiDk4j4Jr6UMMJ1Qeat4RKQJwUeCDC3+
kqvz7r+SyCzzha3wrvuzyATSVKV8+Ap7rT+MBdsdBLgumc9ZNXMAL0PfGcPOPNdF0CfTercsC/Y/
1YbyJ3PW8XXuh9zaFwo+zeNkxQIeyBYmNW54W9WO51+NsggTuM0+FdTRFXHmgsA/MT5+BRUJyV/v
96gCXO9FBGH2RbJlcxt5CShYIeqa31h8LppKN76lG/SXce7N378OXBDrenPcf0POrxGwB2LOh3FN
BPFZDVNnd+Tv6WjKoFCizTKVre6e97KSUb1vGsLLyvGdvv6qYGbdaMDbAXzzoSJGePptGFmnBGHt
znRNPJB/0ccH7g3VQ/arewa1cCiuhdQ6Xf8TkVq9f99kaGaxJ7q2n7fiIcaXWZV9HuRc9RYdbdaf
fR7palnz36F28OMGyT1ujbyXaCfJcbLU3MLSopjqaz7XvhucBe6N+wmPdvc5eCSEo23PhzxKiLfq
XQlI6FanPdaIsogtoCpytnMhOjhP3li+RWClDlvLu/zWL+KlcOk/EoW6JNXiybha6mpz5OwcrA5r
Gke0oRbg3jHevzTfrVTUq7Lwaz3N78qN0rgrydRCpTBmSsLw3byIB8ClktaAkNBD27Syw647D9WD
F3qg5mS4Uhc9sZcZ5HCvM/Wr/+6/x9y1Syv+Urzp1mhViXGFEK32eSXJzOfjIObRSechNMN8q+s5
RJGcho4+VOoDTjGjNYRi0t6hRyldRPaWbJnwhZeSTw16uDTUiy2lUgW21B1rG/LI27UoT5VNGNJX
n4XGXPddf6lE3145c+UleJLldb36pvocP8Qy5TIOJXzUGH3nxvCmx3mTmMiYfYzcAkV6vZYIQVuB
SYprpgD017/H2FDDkAOOxEWx+hMYRSvCAHkG4dDE07bv4rEfI72y0rrhpSSbHKuAtDio38wKdNzh
quZT4DwazcLnykr/bFSSw3eqlHRet/upmn2PVoC70eDxTnd6HJ7icT77KeqbQb4JHH79CRuasi5D
h3Y42BWv5Wpv4wmikTAYYclm/j98cuE42GbChT+exKbiE/qXR0m25oLpINhU7QPKXEAKOLv0APaO
YkXxEsGJKX8l5fhUn8PqnOqfU2x+Yc0aLjCdSlyOruaG7hr2790ObURU/mHbc6hQYSBnMCF5pBr+
7Ho5WrByjiJUANkGVn+xqD2mGh1rqZl6LeYHSQdguHORbdPTj+yN9KKL5mRJLigpviOI7iywpbh/
7nd5IItmTZdvHfq862leqyi3vPjrogN3iLLAS7uMqz0bSedPRvuC1pSTbT+S1pBM183a6eYPn4og
AI5Vb3uY+i6hX9jgItKOSC1lczuaU3gfj873R8KUZOEU+gOFJz7xeRM6xpgaYSzMxFrqNkvnhDKY
ZZIsKsZuFbNRtssRtVvr8L7sf3SfmmTWT9m04a7bRS7MQ5piISduCSpviBB1uOXfuFGDhsd+ZKVP
nNFFCR2cE60x6alluSxO0SXi/qcOUKhHDdvJ1fdmKjYUYgNU3MtY8KYLHfJzIUd9x1HfMFHBQcQw
kWqqTiMy0ow0E1tLm4K7v8lYQBW/1lefbs8Z2cPgSMVMvO5tlvoULi9hZlxSaohwuzmEpDMhSPiF
nSI2MA27aytBFK1VxVq7sNdPdE+K9F4XQkZIptvkK7WiLjWuQXFCkqcqLp9twgaAn2jiFBfGJi43
r3gs6EkvHSnM75Bm6BQ45O1tlHT5i6aA9Wz6gy6RGvBzJfTYVunfZmZasiEAVUt2oMt2D93VVeYB
afb39re45edpoDhNotoky6G92//9ejpIIwAsflk8yxvrfiim4kfz/mAoCivk3nIOlLJiCr7hi/z2
iIFatQFW8m0INuYutuDUkyIz4OhN7aQ4UtDRSDfPSK9WRueHrCzKMJI1Nwgur5x2mJXcsaAJymKo
h1D5Trf5DKc8EA06KATW0lPtac4XrSF8KIE1CvA/o5LsYemmQveI8x/MFKlZs+ggFgs2bllaqZ+i
OG1Uv2myw1o8Ysrw0gSt5Irk1UIOrC4cxGGNRzlNH74LC4FwEJlouPM4NtkRYis2M017ocWcStjf
sMc9ZoS0yVlE+l+kY+ayL/SgwvxfRjZ4+UGASit1/GD1Url2zQoQpFesyjqB/ASiRvaEpXaKe+ZC
b+91FwBlGUzf3CPDCwV+tMNZLmDGj/KNihrD4awhSmFNa1A3FeODRNLWipreJUf46AQ824mIOXSw
8vmLA2w5pz61/bTAJNiXw/aH+QDfWygWWIXyzwpRfJEwRTyWAR0/LP11LvqAce/czqKs56SIGOvm
8Ret2aN9gwzw9TDtvd12zRO+yF8CzfOQcLgDEeQuma6GdCIZKcNQldMi9R3LVkN2JDjn3wocerWU
6SkOVFJ3ciE1If8z4bmqqd4kSsaTCEpZSnPJAW7vTjE/H6zwv1oN15MxbTMW9MAnEqZQxwxSD9Jq
2/5RES8SuVUWAZnjpeDFpRMdCYBd7yLO7dmPGor/q9GOl5EFlzFNx/zGntE/w89i8YZbFXUtq1Av
ATNJvm3QidosnRqNkmRnkyeAPd80b9LUuXRz5HbFHYGBZrZ5VXr/5sIa7PTapC7bvX8dOwpmkwPh
rHqgyMDlfWHC/vHpRAQVxj9rfLlwnI+jeJr3rPyDpkwr1D10F5HYF3tMnQB0qdd+qgw7mrnhZd44
rMQlBKIsa7mCAOotAY/G7xML0/Ha/FwklYkj+ajAWKvMkolRkdlGNRUAgq2d3TpGlknUka7C8ghY
itpmkmfz/2rFOHbE2X8UlBPVuVB7jX1s1vX65msGkw2oJvWTBiNOqN9yUCJOqNUxAr4pKB4Nj6xP
EOF2JrqZcpIKxyPIsRae+yvrFA13NGXFaZddYss+egaCBxOWHUBY7QMVHoBM3rn+rmGCwe4H3aMn
y49aXR2sCTTkf0dY7bmc4NbXf8GWYiJh81L/cH6UgcREcH6cEvFkD6jVrfXMAlHQSSdvBuHAtXqg
0J7ZE4mDJD9rkKcwe7Lzz6Pc7Dfo4LoGvIC0MJ4MxKkGbG8afICIGaukAOIdNcfrGrmt+kgoHS3a
Wh+ruj5XoTfJf07E4nEFI7dlKbiIkSSF+GnuCO/Qm8kNzr89r2TczCoC675kIIIkefkucN2V9K6N
EZVSOc0WE4vhNegmu8+5YpFe74phBAXvT/ksLZJeV3V76zKo/CNyv+U7ca4vmzGmBirbMY6UyKSe
i0sKzsReEmpg24q2SubF9RymRHyfK3/+afWNGD88en23QEpmaqq/8rQ7e6Paf3ZLfQSUxZqdPvI1
WA8zwF6Xk4LmzbDodvXRzRCZVt8YvWm1jQFFHcoGr5gam7DyuLhL1eecpN+DELp3eZk5XgT0Bbdt
h+pgiULzhPfUAIRe99E9Fe8+bvGvHqTYeaUy7D4Dr5oX3DoBA+yKHAy5nNNjHaLBGyzxR18a1yzV
K8ZUoMY3LkasFwrdNCiH3/slhxqV4XH17fVSdGZgfvrE1VxwgpT/ImHWwXWY2ZU8pozRtV4WXq0x
2prWtY3eOc0iHfAv5RT0ZMUFqXAbFCE/8SMoP6MSZjVu3RidNWZkM6vc2HMbzP7xW0PsBqw3Upjt
Q2muTGXEUDLT4mlHCyvBzRDitjwY9ECWMFEVr5fyXcw9T1upzfALR/Kq2cGI+oISML506A5RyqT/
1Vg9fHg607+pfjHc/8BGJIKNflrByHcfSIEB1jOobmFj5QS5Flckrg5yWYMz+mhs3gTZDg0tS2IP
CzLD/ncyplhUqgVsvn75LdfLS2O4xPxl0X749247wlX+tNxHxpvDg4vspIYpHIsCjx5aHnMc0yFJ
YuHOv5i4XXPbmv4J9K32cvg8hCbmrkAm0BYHpQXBs1br/QaUGsv6sEO7vPzlWrplSFzWRWR8VBLs
lSjZsaSdkT5F9riDRSz0XS8e8wLuACt/6Nza6yNuOu0e2TZQCxqNE3GwMl48YrQGYuc8rBB7PZf9
2y75t0Xpg0RMgDVzl3kZpFeeHqOsWKdF24QN/qsNdg1KPN14OADC2Uz5g/vYAjINo91U4mpfd0DM
W7rC+fdQ1h0MxuTMbv0dkng9I+t6x6fAyziA7Bpxq5aDZZpD7Lti3Sk2YkAXG0p4TdlYrr5tlnbt
OO5x0/fJBSk8hN441maODAlba4ulwn7+sgok+3avTtVoV5heaJYCAjGG+f17klzZh+E3i1V+zbuu
fz+BfeTjBE8iOslWTWm3Zm94vl7D0KRhcJzQdJYj/f5RuYHdB4Xx7xClpzmM0SowcqanIbgmCCjl
+3S0jvY+dpiH2dWduTUcIAuJTirFMf03uIYbbg4h+eMKR31vkjAY8WkIg8p3pjzr5g5UyPKtApJS
k9MG/VEx1SKmcgDHgIIyXnOULKgrIDNmuil83O6DSENgI6zxByEBg4Qkft8ZM4yXA3lAID4rWvwn
C/T0ItNZXztrf/32/hxvd4P8zmQozvetpEPAh589f9K9TvRO/7jk7WN1oron143fyRVhmQLoS3bg
iIdMcuqenxwgi6cK80/HzC5GVbuPaLztvtPIj1lgMxFFwd7Y48TTz4/ZJ0ojIN51wL9ufV/xEpXh
Sn/eg2NGEc21sTaqCw8Jx3V8ilsIZBf7YFm9rkMERLY4fRxG4jMgqfW+aBKZO2yRbr42iYh2ReyR
RkyrXKgaaXYEEiioALyaBpg9VpI07MHNVNCnD+8NyYQUfrFjby7w3wTlulyMIn54oTpRFmcqneZr
YcKQjhi0tR+w2k8J+4U+Q1J8K4Q9aCKOqVa4D3FX6R8Xn/154y85ytPF6Gxj0Xif9qTkCNmJdRPY
oc1elj4M3dO4QnljCVOZJC3p55R5aQVNHVtR6WZZyl3bdsvyruIZsxJt4xdmO9R2lI/IV1bWpIxy
n4gi7t4lgzzuTs/zKST7HsC2eNFLPRFKCEUVcjaIkmDWSX59QqLWaPCiz7/9WG3AOpTsUA+cBIKa
8bwA/K5+0xGmWtCrJ6pTS1OK9DwEOXBBrfJslnibgXN30JmhyLbjnUDwIVFM/4Ic+AShPjnkeujc
w5/VAy01UXyZCTpoaze4tkoc97Cbzkaa8Pk86KSV1vMcshYnItM7Ywx+cu247z5LXWXfDEHSz8fu
Iogj7RA4aEBOUNSMHfSnX+udun25t1QhoboJHct1hdeiSF29lq0HrqaryEaekHlaR7F0jNY5QxbS
LJM4CfR+CfYbZJMUNI2x/ct8kljCnDbKc2rvi7j7IerfwcD/pwxEGZ/xGf29ucBAnCup3VPaUs5S
jeySFT1DKi7X1mNPZiIAysJTCE/EIy8fVnt+1ubdpdB8GWiypj/aEHIZdc3FXcwWfDJLzKW6o20W
aLsB5yHjcH5MZ4eKHguN6EvKj5DqdFVZR6doLYwZCYAwuFMPjuYSkVm6rN2qOf4unggV0vDHGsnb
SVv2TSEI7zwoF6xgMj35j6v9CptogZSFSNYJc24oYvVk7M06MBWQmS7mSrcD3RB36rvBT32T8rUE
aRsKjR473ldZ6nonpJAgsvaMv58pkg5UfHRvj+/UgUKSDgmAneElQ4PBloMgOaZ5eKO3wMSWXXTc
JkcN09nq486xgJt1yc7QT5JnD8QwnPs18bUH2606pPgGhSkl0zGX0/xGduFSQB+qv/u2qBtMVb2q
xNXZ070gY4Zqw6vNT4Hilh5P65n6sEcM/Qqk2lSJfchKlKJpnUXKhenJcl6ciGIALnhl2dk0oUgd
d8vpwN2WFCxKC5eQ1ikvpWW8CPNm5MCtbbmmLtKvpR47/mdGZGD10eaBygen2VedKCaiaqQaIRk4
ay5+veizYPQ2ptFzsaY/wPgj+kLiNjpDWxX9HLurSVkGqpxmsjvycglhBxf++ngNLszl4JQFFQF9
Rl3s4qudBW3icv4V/IMCR2f0lKL6OaC/PmF124CZMv4eIis81KXugGfMQaF2GoISmWySpVmIsnjt
gxYZEFb3JgvenIwa/wVqhxISaO/ANO0aiss++eXrkwi26svqVW44i4oUAyFLZMald0APMTa6b+r2
g+o19a0m9En2u97CM7X0OZuao9eTXCWHqPJ47VfJHOCRvbqYZuO4j3ZJFAasnlZIkm9KX2+7KUvA
GwDfUZkFmjWPE2kuLLk7r7CBw6vdNG0WcYBPjiguF29TR+0DvTEWxcoynkjwJktCkWvj/74yZApB
NbWSehHqkXNjZlgOn+iHlCH1ql1+76cMrQZ9uvQcskSABDykZKe5bwiOytsBNkFzTkEBXf4voDwv
ylfcYOweEqODDA9j3J5YJ2Mx5BxDxbC23zgs0roJqn1TaVwIa/2/7HUdkU8yyt9dxfsJmBY/2ZoC
UvBRjRRdtyYcM5CgD/Sk96csF44zLHbGXg4pIaeneKJb0NHpkYOzPsgeWSCZJHKwjIqEFglTfoFA
Hx9S+1CDLj0TKapRH4s+worWJ5X57NQ+9eTbuf9+0DKe63KVntHfQUxTk06QZn+mAVvH7RKt1yoG
nS/T4KKOExuemHxg4kBzu7IY0/FhXLn9V8GjwyGUFd+X6TO3SXIh+xVs3NHTfjikH1kSZcsVlsBd
kUwwj6Va42ywHnbMjCP6ccsBDHdGSDDzxjlHT/U2M9ZBqQGdFcuJfhYCUryTR9Kwxl1r+e3i0qpr
VueHiRF/6f4nVu4M3y/BtTw4zP1FhTBF8R+xccjY30ndQ+acMjPTXzQ6z9SainWbgJJNbl/9iw4D
dqt3t7ujwMxoQ2brtGRpnGJR9OaNKXrzJhsgKh9cR+zFX0OJCnHtbmrcB4QY8ojB7lPa7/PuZhhh
OXjJnBHJav4O29UnPCZYsgmFUjJtv0Tk/imP18H/xH+O2dRs053O169rf7zqMrU3Ti+g4hJSfkXp
7agnA0E85/couhxFATBHM+bHOHIktoH3TPcjZ+DmaCSxEOEm9oOYxp1WNLquSpKnY8PKavBr8ciW
dyK6mwS3Mv90fCihGCby76DLb46DouItGNl8lt8Dg1qLOkUfZ3X3wCWS6e1ApctwOZDR8Pf63m8t
PgAnPcLSG7D9YbCQ3mW5LH6+ZT736TFz/9AAJ0ZLr0WTC7I10IZzZdBKgs2ou8AF1AJEmByM7wH3
wkH3KnD3EvBvX2hu0ossd1VcE84QZ9n37V+dSX2u9rpulj2F/DM6oFFpiq8rB0js2vZvqsJaLLbA
uS7qMAMQNXkA7/DoByho0q//l9yA7HSoZlXW9Tch/ZNlezh8Yoh4upI1Ce4Q4gWiW7Hghv9H/Zob
N+LkwU2aTUd4hvgYOnzti3od4aVFxOZefAonAQmgFdfZwhAD237GpnNOswZaiTiAEVPoZHtoYQGO
GOLSSq9UsP5VEZVlRwLxdzGdYpPI0tclgE73c7KG/MO1fnsxGki7aSKTd/ArtXe18gwN+SG297nM
EszPrW6+bJjxugwkLB8utOuAxfTwG+0o+tQzR9+qQ2H4sSBnrNlKTQ4jdx/j4eJ3AHz8HT/aPP1w
OKfi+R4rwp7thZsRVzsOn/CbB73Mq6U85ok2HLWfsFY1bqLShPXGXGKWvYXTcGgQ/mVJAGZylMIn
VuQwAu2/Jnyei7Q/ZnWVP7S3KWxscadNgacOjc72VcdSuCJbC9leff08sDktkVMjLeJYQgyl1FkQ
4NfMFW3UkQxOwKbQCqHR8QfBhLyzz6HMZDJg4TxNdFrY/AN6YFZgcA4KR9Ps0jwVaBpGuwxHyCDH
24F4xfXtfBYpoCTEi8cq2/Y5sZUkforlT+AB0orpJPxtFJeIGCepwdIPCpCwvvWH2S4uYsZUh8hK
kd6RtCImgpYUxC2vVrKW/+lxMsGVWaDfQ+4alzBQ0QGeB3c0qup0TKY6cLMH0Do4YU8CrfzsNYQv
cYBPIHbeGIIManwID52KwHVzsBubz7ZMzgdsWYCup8WT4yI9ZaA5FiNWFQcIwNuQsz2E0qp6CAk6
WsncXbU5sh8XkJph55yTYerGhldBTMzHcqqPukIHpaWKUqF75q+GwuMiBOAsNVGLltWBpsYTxETY
r8K2s0QGxblCUndo7ipi07ngCYJf141Je94VwiBNjsn0T0tmqZzmdmRQBICbN/bXfwIf6EiJVwyp
WwxCSI1NjF/pz1ay14jzJlSgEaJtVhi70rM+HU3dmgrnSgSxWhqXzNvzrYKWSbl+wE3eMvnHwwyW
6889v9vq040Fd7lyLJRpStM3HpTHFpOygVp0CSLX7xcaZpenySSE2xk2653RblF7FG+IJge9eySL
NUlXzis+Efq99no8yjfY/0DxyMmerJvB2KMlx6iy3be5yMysnstHv1O2xfFShQEdHTj1nhuEjZ9d
FL7+PUiyuKawjRsmGVldn9dnCwEZifOts+X1UuPsaarU5xRAfahXcrwMI4Y/+sm7PLWvOTrhHvik
+UOjk2iqm/tSJb950KoJmr/z2Xuq89T0eYYYO+pMNP3djM3g/vZnsTaluS/CMFawmEAoMt/6ibio
zj0bDXN7YlBkZjtxEcYpVN5N+OEK+/MamO89BDJItwipc9aL3vX+zy3dILPNNhLiBVEzzw5OVzbj
/CeRdos6eb99bKxM02Mx65CpwmL918qgoZ4dez0WfzrVcjROROI27/l6LL1QSXLzs/zlOJ9eZMn7
JeCJRVBeAaFw6hCk0FaoUKsA6Wu/DyTJIHiPP4ufnGJsUUMJb5Rhb06N0HDhr92LqYxGZfi0M4zW
G8wztvhhBvwrZY3X0Yy4eQl3S7fQsqbtuTojkHWe7HGjVo56EzTyGLV8M0lqtJG9HPpHzHaiOUod
aaueVXne125iII4nFjO8jjpp1NuWY1QibpZmy33fcXTw1AX/Y+3yOiSruK69ndmi8rnAuZ4V+5bu
j+2mK4svKLdp7JUoo1Jj+ARMj7yXBNyR26AWML+bysH2uKceBZ/m2y0r4yUrXWljlkTyWQ+DWyCO
EaJNTvJPgeiXnoDufGKCvjF56KRKve2+8NJB8aW68MhVbmC9/90gRZzgIjbi30yOVPWUa67AiOHF
klbozYQlUljAefCjx4L7CqrEQfh/TV9yNYdvwLnF2TRl45iKhKHlEjNVIaRLEB6jXsE7XXxoU0EQ
dQsQ6JJWERg5nndYAsUDfAr2+jYXie44BQkmVi9kQGVskV6mpn3x9qjskSHcBKaUk7DAH+p8PHwd
VMBSSJrWlCKzTHOjYWCJ7zBxzbFolaxowLK0D1RMTkDLjZtYLvZnGNUk2rEzgKYZ74Y6XWwk30rY
PxxVTSiGNpFxulfkmZ/WKzp27lVEQDzGd/atJBJa48UF6nrYHAomsYJJaDx4ehUfKR25Zi10G8Bu
u5IK01Z9U6nwEtgRkfa0f+Pp8jcxFExDhhKMAqh6TvJkZtQEkEdPXlD8ayBLn4zpW1aVeu9WNcfs
EeWopHTZu7HpjsjxZCa1Nd3zIQz4uIRCsLguo7HKu46/zk3NM1AmFbr50RHfKAgHegdiXQBMbUKs
YU7VJGL1l0tpHvxwcSZHxHjkqesByE0vMCP648RIrLm7qKdggHmCPTiNEVeoSnZ3Zc/AwmE2qFuv
QF3QxGhogFmRnb01IXOM9Jpz3PMTwDoItBkK3QpYoqZYmbqUAyYU7O2c8guA/6VZN4AXn9MRTHwj
CERShQ9LiHIpZKFjclLF+7yl/V9gHQ5YRhXIJ1lT95B5zd8sSdHBDBPIrIcdB3+opdfuz6t/mpO1
FXj5TZrSn7TMDr2RWt4VT8RnVv6X4MjthTU4lH4FTnAX+RNF9VesQvy4OaS2BWtTminGRNpM2T9K
1CFhpcM2f3L7LPPboqeM0+XYgHOhQvlbFUmuV+rqcz8W3jIqhz7hiEO1uCvKVtM351qOeqg7WR1G
Lr3kWPgjtSisNtCHpuJSySbYD0f1gjzTkdkEn6TDgS5hoEhYq1/XILpwZLZyMmg+zXyyq2kLu6jF
KFtR6UVdItPiRHTaLQj1cKMZ0EP8IUcinKbx2TIamKrlSkyPkrljBJT1fagARbN95OLAf6jZ/sAU
U7NSWlpmtm2RSd/wIQT1VMra5yUCoIzFymtxvoKEcsFbRZZFtE8y8ekvvA3a0TIC2y6RE1wpgKMw
71t0Gyift9oILO0YB/jAvaKSYROwvhrPGLCJJtinjciz2ylH9dYTcb9vnP2TOycuFSXqfrsHDHxT
6PBo5Vf1Q3C9WDkp3Hnb24T91mxRM+8zqV6oYqVXyI0gWp6qmcY48aUO7WgyI3+4YaVNtrcl+dj7
ZMlu/KsGqffa35bytQYIEOufUNXgIAuaS4HMSwE/9i0pD7nzbliUvpydHRrybt3fsReAcV7ONCWL
+AVrnBkDyZmpSpnrTwPo8XrzTPiFhaYH+boGwXivvMjX8fJP/dfWQ/ZIAo8i6yUId9fOpGOZGLtA
0VfixnwfAI5HJMYNY96ltfDw7st4bWGvN/YGxdOGg9BX7oPFEMlo3oL+q5Iao2dsbCF5Mn9I7Bc1
qQvP2D8bXOQNQuuNRKc4Ofapk3KXj4IZJWMuFDHa0UYGT4aTOajRhmhR3tIxHeFDIR0gE9IGTEBM
WC/LOnx9lcS60q2X+RVNQMk1cYhk/+1+st7EZhiI9YNOrWAh/kZUjG2fKcG4/DuwVwpBACnvnBpu
Wy9KXA4+DtJoPk2wQyV7gCK1N6wi7NnR7DErzd1PAhy+hmsJKNfBYRfvgq+ys1YmUiYw/KawRTXx
HsPeoVOCOlkm+B7cI/Q+FS3bmtPL863sgab7TpS1sBSaLW4YDf6WJ+gdI7IXNN5bOgtKGm4HUWC0
C+dwpfJoDaf5Tk9VEoWHWjRc2yQK2xvPqUJ8GrOJjUwBBHo8SMScDnCFepHVIbXZVnq+j/YIe1Lu
DMr4smAVynJMuyuP8QctgXdI5QJh5p+xrnhtiQAkH5RHE0NAPCG2hlhVQIBfW79Hnnbu2HG1a/Va
oZHL+IkZl8Drh7pUYtr0Zx7OXADJj82ATzQCgfB+ZE5UXHlUFCcOiZSiP97i9nM6Zmvigg7fMQDk
QIs1aTWSZFJi8g9zM/SI9yVE7pL9QHvvYHjeN2GXNJEX/sftBeTm2k2fBbmADahuG4NbY7Dz8cmN
itV3KlNEd9574aZkvXw7BW8ifthpAbZaKtRwQsgVBnuwtOkvWlv6lzn+JnPLBuHXUMkr3ewWW2zE
iEo0O7rzMUiBu5p0dc9jT7hMNI/ZXbwvPf69u4PD5hvEXitTQVV4qPru/73N+Aqg/4oztPdq5Pam
Bf2WBr4parVx1+LS4l3IugC9iRmGvCEPhYIpIYEGsjKj/pNyXgEtZmRysqL0e5yLeEGFemi+9dgi
xtKyeZb6/kbS0MjSzV/InNPAM0yvVAYmUaFc/pdQcZ1XV+cSJVNbS+t6cf3OVWFrafSYQhM7Y678
IqPmhmMoKsUTqSBzDKt8beqikMAJ3NYDQqyWLVTxUKkGsPcYjD5gpPO2avyIRFFI3UjBb8M5xhbI
S4dXw3JVvioNRiT8PMK59YAZ2XpzxMeKPEnu5cQ5DuXckizPXfwgEg5pXz9gFtbGeSe8607IIb2k
VV+dRf9TEgFr4r1pv+lzjfyhVuEkv3rxpE1JQz+w7bowf95qE8nTknSLyqxPToIjbiCZdw9ULajX
dglbIsRQ6eJnpTrqPUnOQNcwP1YmHfEeCBouj61GNLub7rMzapg1GXcgzEtZsRPqXmM5xM+iebn8
RaDTylL4xEBJB9baxwJO6I7bJmv/whGAO2PWzcGKPYel0sVp5J3W3ylJolw7an745JhUUT8qNtpo
fPL0ZkijIiaFXVnTKbDzS1gtEBEQ4U0rvLTe/S9UFthRrpMx481kvQyXtMPzLJGYhoKaRoe8Smf9
VWiN5HGKV4ESu/uhyrFy+peji6YVjf5JoGQpFKMI2jaaaTXZjQjHGBiGZ8r9U/Vfb3HPavh1vDrz
7/EEPRRHGx8EeXNoEoupBLaunPSNXYzO6zDmfvp4soeGUHIQ5CDL6byU/eI4aqpMvWlQfHxhoaDM
b9z6YbyV3cOJ7+iMX0o2uvnqaqOFYDiGkGft7+dJGj91aKMTcj/l57MUNKsTyqjnho9YQbqos47n
lG3/EMtJ/no5zC5WYkKrX/3z+NvKoZdeMs05UxCAcVtP6A0Itk4fNZoJhIsfK2OfVe7zEJU0rwPK
EP11JVIj6bStw4lnqEgkQ0RpK4N96W1jwBxHcmX4aHayGkn3plSk/h4O1dT8sVmR8YVjHT7IoHcg
Tc0Kn63TP+ixCx9XzBlPVzbF7AO9Xfez+m0TRDiXb3/1RpdK1YGZKZkiOQt2JFW8qUmwxyTqAzGL
PERmjPPGpL1Vp690hctDGWwjOzVi70y97hS9k1UzIZefpCZgPHPyNTozH/CmScJhhaKPmW69l+Ye
v5ZH50V9p105F8wrC9kJXHG/7at9QPqK42tpa8Qq1jQDtLFvbFieqQWw/l1aRhe9a6Mg+HnDXC6g
7L6nS4esOvAhdegZhHnTyg2izcd+jyGi4S0NPHX1EEhMkEqt5fMDmJI4R/nuEXFmAlM9mTLv90GT
NbcFZC/95pUKn0a6vX00LruW0toqeQQNfy7Qizk66DqU+ZwHMIM5Upi4dWPo+svH0q/z3GEeGz4G
+qsJgm/jK1AdMMaJIxXocuVl3YW9is8/EcXoRCJGj6WlfFd7X5UqJuN4/CbWnYtHj3XLzIUocKZK
U2cjHf3sXCTE5gv9OhN/g0bzQUjgXL5tf3SK4RJWvkkTcWi2gtiiFamQpSvoQeU5Y70EyQZ4Emd+
6seFsBbe6nZvm51ifb3XJ0MbCdVPYJyqIGcruOSVJEfix3/d1i8kS1DmuIU0ssk4PqwpkNWvffTf
SO7CC+6PEPzfKJu+YU/8KGv3dbLOjLi+E2Lz6vKmX/Jvaf00V9FS/bgjbbOqyD+5RBIxIvRBPpvg
XtUmsmxNKVRneuKcnf11DCy0f4U7H2wPKukGkq0QDRWfV4qI7Labz62pc6wFQQx0ZUAgTqWCRTpR
HWL56oQ66/lbNVJ0UDExh8KE0Mg1pUOpGwhXAAcTRYByVTpL7j0fwIjQQL6tLGtipbxoxkxzg1iR
QzuwHcxZntPjM3rjanTaD2Nm/RLy9h92hLRIKo+2441LVLJrKtweKmDE2RC+sG8UzB66UkCQ/0p9
Wci6vIyp607CajCoOV0Wgwx7WUtXbdgPElQzjsZBGJqOTrl1X7WUGdnDB3VyRMx9PUlBcmV/w0g5
RFi90yaM8UAhAfN//+E04AY7+SXjyooZG6qLASkrDqmlpTNlHwDiQ+vzlQKQ5fWYkfszfhrP4LPR
GqKVOovFTHYXVUe0nxvEklJCt7Ch7Hr/oVOFOghj1BX01G80fD94HXgLzvoNJEm9uMQxR7F/t78i
QeF4aShp1Nj8EsaJq4fM6rYt5+wJoLdkbrpZPFebJy8O+q0hIMLgy6sRokCpiP959zmrGAlS1YMn
1erhAn2ZcLLm/1OHJhr3PocCzKyDi2GE5R8QgDunQ+cX1DNKMZWa3pF0ex+b4iL9PJAbgVAv2PcF
WnFku7C3+jIMw0RONYsoNWDIcOU4s4jUQCH2ro7m/IMuxJ4fBjAoblRg/+GE8xB9WkJG79CqN0Uf
nmSTBVVwAwVY17X3bOKswTVNHer+9sgChx4KpKt58i0cr2ZfsT9x2PXNR+VO2FUXZIdRf+I7MNy9
puBYiy495qK+Nj/1Xi8DogbyPnn/Vsk0PfK5nk04OrUIdorCMeE6zmE9g7q27+h8hddplD4AIE91
UhKueiqVEZl+3GCq/vveoM77rrrggQ6Sf56eZ39LZ0ypmihIZ97vav3/d+sYrmvPHu8CgmtreJAv
pG3/XPFpJUIN6F5AZIIi2f8X4KMU02KLSdvcosfTwVRUbAivJUKhPLPNXSjOiOyUINJjScaSsMyC
BOc7CZ9hf0YAFZ+3joQUb71PpXdawYbQlTDAgjvNNIit+U+u0A5+XoY+AYyF7Hw+UZcpWo6sXoBH
NIfRpelIlblzbg3kdkq4lPv/CDGUnpyz/BLfwmaTHJ3Y3oIdSt5gY0V8Jwm/P/JGk5REtciqU0K2
x3bed+9r5Bu1BKQlMYVLeIKigoYdIFVTg47pwjDB9LgoSCrow2nAlE9J3wukajABeI2dtOXVxtsk
uhRq8mNSwjPvnh6IXxVCniXaOMU1ODShMx/3O/m0v1ARuTCXPlWF6zh4GXbFASOLUAh8eHcZuqBH
S/I+z3MVfWXaiJ673P92onWnDycxAEU5PgHE0Mdw579ga8GP2pGcQs6HGmqSfJr0AHYmUN7T22gr
rAGUYctlLkMyxwD3nFqGjkBfdnptkPsNPyEY5uRCBoMOKQckAb/WLSXFn9M4qgLYV5CiCePMt+KN
Ov+xI3PC0TQ5D1igl5oYxy6GxWIVOH+Py4vdLGjducQthY205P8vR5mZb5nYn0kGzyP9RutUhwHR
qCKS7fod3GGyR1tfFq3uGHeqxhfdwYlvdvFXnh5Ed8n43h0+BlTbDQvMZ77aw3WEQV1+G3t+E+eT
5b3rhQc8S3ENcQYvu7AFwVMJI8HSTIItXJ8ar7fjsWsLGeqXF56gNJ3ath/9rlT8h1VH4/lZQjGH
oco60Uz0AQxBgh4noAu0Bi6kmYY+ThmY2K8T2nbo6WRMk36jdNndc6OPiNtU3flfGrj1W/Nonidw
YbW9WA6/axhOi5eFxvsiig4+ynUEjPaCSjRb5BOg7E+5hU/CEXwyRw31+QLgN/BtkkQH35ozcrCt
2rW+1Y4or2G2JZNlXZtaeKXKA564CIxRiCgJYPM2e4hh5RkK90XAt4NG27qnPyGf8bENyo4NKYD6
fizxIz4a0MW5ACrIRuBHt3C8lw0TZR3mdQjPOIyIqcg+D7uwKUrjUKUKeBp2bq3kp4yN/X7ou8EU
c9G4ux/bwSt09vkHKqs28Z8R6nHOjPPmHnbg+v4s/dpv342ks6XMN5Y3cvw8mJ/fOQ0ZAltUNbyd
6U719Bd3pFNpTJ8fn9kUaDS2Mjdz+Qr92V7FxYwNGdjg0RbPxuQ8b6bTYztwEVPUfO9EFJCFW62y
FUnvI9I9vClwhcHCG5N1kvVsDt1ZBY7RzjPeX3M3zMBL9F+n3/50yeqnVTKlUqMqfXas/Kzq1/a3
YHZbZkov3vOwuE6KN+n/6l1Hq0znRZ5KiaWcN/7n1hoHs77QJlWpx33JbxKhA+rohH+mVhX7tzL0
5AE+O2VGAY3RP9VVzlO36qP3fuVHALiGKrHYPWN9BLT9LZJqL8iEELY9wBXaXDnNYuiCvgOPjXoK
kDjeXLpCevX27wRVH7SZnT0g/rsW2OQiV8UWIQn1uZNT6oFgVPCXQuHCxSZwYTnvHKdPCwdI3+hy
CPmC46t3tyGkBvTOxIc0gfO5tYMDwbeLEUv8nz1zI6aqAipKkHWuYlcXLnoJ2I4dM1dnVwxvxL3w
MpSud104Ov+cOtQApJww1aqD40eTVzY8BgU/upTGXt816PPCddDItQLQaLTCx7VFpnyxCrcbvsfZ
5H/ODFXSmz5qsycQemkQSE4O0TobuFpCRmSjPYG3EeK038zCtrPQtb3Y9KjirAAMxP3h5YRjFhl1
x/Le8yv6PIIHHNnz6jfKLmApiwqY2+swM8jETxQlH9jLLg5p4zQKUjLk43Apse+HYeNHRiH96chq
MNgl4+Yv8QBZyJhHtJsU+dXkPWxSsxGeXxaZQdr1LFBM7BTab8SV/4aJHi0oMDw+dawlEgiZD8k9
EgdgWZDb5jSCopcU/MvBA9dnGWsVpv/I7y77ghcOeDzzMHFeUNy0egLNoSNdEKrrkEMQ8HCbmlah
rlOD2mDCk+H/YbnX1/aIvxgHlp9B/o/VzpgAkSCUfJ2EmMkp4iZ6qvIbVIF/JTQgMGH8oxlRw3P3
PqrpWFhB6Y5/vMmKBCJnbqe+VvpmDiVSAROaJngdqU1jwfEYP/f9WlaHqra8eL62
`protect end_protected
