`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
kb94pcV1knhKexJRl/9sy7SM3McJjMsiJ5a3JxJ4PLlIpxbL5nAX98FfIlFxXF7MhWwPxxHTBdz5
IE6tGVn3oEsTZt14ouUNlYI4cMcdv3tXGS+2iAc4YwcOXlIs7ny0z+e90mzRgmDwopccW49bX+WA
6F2fLKAObn4983ji2Ww+ufPD0OmDQNFoUi3zYtY123yUecsOBFvEd/vafqOcEZw6OwSVyQ6gJ/NP
1DE/Um1hhNmx3pWcy0kOnlknvomr8NmDUv+a/F6mXNswxEn9IjqM4RvvegylJUpRToNRsxJKTa7E
v//urRWZY/85HvGQBvd4+A33dlBt7NBn2YPTQw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="QTPeGIV+NGLcZh9sLNfinXWa7KfxVpvzzztMTySwPBI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6544)
`protect data_block
xGtRmKzVDi9wkm7ixa5r2o7u9OVFw+HuCoRxRspdj7O1dkGlnjFCZUPn5fkQ6K1hc4rVfntRcevC
tC9Zpb674//jp2YCT4aU0pLgboTuJpAsVICqJbYUpZEGNTrihIHlPYe5a4ZEBTeJn8W2KqRbg/n6
+MJC0k1+g7eDiJuv5rNZhv9s38blZorLF8cSVKLiq5ccPnu4QQRVvWrMn74NMLVYy/pyP55JQx+t
3yrBQvKQ52Vgk+FcQKtitlsmA60N62xm4tw2WK2s2XpOk9rWC82xTtccFqH0K6thpTmnXgeybz02
Iag9gxx4ct6NsX9PcbsIc17nUAlH1DnxKcqHgfs9AxJUZEUHTHNE7RmG6QYaQudRr9iMxLwQ28gV
gcxYGS3fCYD2OganyA5GQQbr9orqj/3/kcwa6sROtljGbTemYki/MZpopB6z+y1Lp161oAnXMNi0
kVvLeLeS4g/Gh+ZiXGTd5VKBllvV0bXrLXzTBdSIcChuhkV6C7yvgruSSXnwjClwOb3Lvv8OpwAJ
dqiJyUuUCh40a470VHh/KiaalDE59LRZbSU+tatJLm8nvrVolS7qtp82MHiYfhCbDcwNWBtY/Hf5
4H9Zfz0MUqvgamrba35tsPPj5OPwIyUOGHilvumYKdnYxz48TfyhItEsCnReBvnAlL76fO6ao7gR
9KvlEXUfAbVbHtrrg+McNDn9vk9toWyo/YyGtKXTOrbfyuVttv7fs50ZzEUfjWiBT5Me1CWCY4wO
AAlmLSk4/gOGWuya8HclS7gzoGv6w2E0t2/GPCo5leredvb2fP6wRnXPRkYfKvzchLEm9fd6WSs3
IpTTsEl4Ul3TdTBVFnmqsU4lFqR50E+1Hg8t6enazH42d4EHO6UkLj7QB+N8/to+hWO4UYtxFpBk
vkWyv0CX8hpUbI2nwQaiqO+TQybLjsMVI8so1bMViRXAygCLaBzWGgA9M8hiC4amdpjFvnmrK5r/
4q3SnxmFpVP8SbDXrOfVUgz8ve+OMX+H7Eix0FDTD6XWjlmcqpYrD6xfPl4vf6ImMUHyRa3egcez
26H3oStYlUujtu1Ttm/GHlSXsSZM+pzEhznS08FHuFA3UHeReW2dqiE5OU9MkrH+UY8jk86XiExb
gzs/d27qI2jVJy0b/zZC6CERLLGftUnEU5ng7GF9cdwoOU/rZAMWgpFPEuxWb5Wp+W5MEbkQi+vt
5R2NoRlKAYTxPDsHThLuDfTW/E0HTBcyx8yS9MBpVLR13Gyyg61vrXEgCCspm8OtQOWw3RayVPZs
+NvfbwUCsGtpcc72UGNgrIsebcvXYPLVz8wOFAX/JOZOtP4Xa/JbdizVTtyJ/ouQdLowvchZC3Te
mjbLVjIzxvg/mIiqIye15Iez1VCzDdyxvYSPoVOxHvSJuRA8FZVtKwqUqZZ9tYtnXWKabXYiwXc+
xZ1GE9RFqPFqHpTr6JgMT8gQmiAPsWCebMEmxRK36Q4gs8hs2T+vHVOdYjAbHdN5N437ZjVXnTw3
3nHI/jIrtsJYNz0+X1Ug0jGF2HwkW6W0i+LRXon1EPMGgd5rNwR+FDpRcyjTJ2sYp5FoeCCHU8az
RB4ew5HUknrPbCzEtAyoJ2W8B1QXlIB9I/LNyZeZWczpqYY4vCnBH+LKixeLjsgWeIELqvKddQ6D
TC6sI6eWPRe4JUX0VdR4b6yqwfrlSQq5k4d5qjMeZJaerkjnnIhKDH9sOTGmHUPjBCtXJoGYhgdR
H/smpICpZuOQFbF46Fdmz8mtes/cMJMr1hgwvCMkrOSrwNwt46MBs/OMhWTkRFPtFJ8+vCrHwDMA
FWv21jsDAlG9cZkQ/TXjbZPLRDkhtXrACE2IKzp7E1AqRtvmiuYyq6BZR6Q1gpKY/rOUIUyMh1RR
SstfQcF/cS1FWiasqiW33OH+37g+R72DmPwaqyjYP0o7r6gOf5EPQPBFN8cTTls8sU3gajfRiLjk
QjvX7t6DmCbXb+mnG1nk2q4kCGCHu6rJAT8nTJi2vh4A9rF8IPbi/1IUzCVCSaZRfL+eUkusbhy8
nZZTAn3/z7Zshpc+/pL20owxNXbtWnt3xSB8Wkb9+a9/bv7N07cwHryOYc3bMZb6YJxsbT5xVXfj
FBmzCEyxxT/ho24CbXIQA5Enx4CBiZT2kWH9aPxGLsk7bp5WwFtb7Q4h0tkAsfeCE61Zm93ZZGI/
wTIAgb22hwoljbommE0KLRVhyOgAw5P1Lv0Q2f6ygFPP5kfYp3+Wtu5elQQTl3XAUe90ktEEq+My
ZzNOlpOZaRs99m9Fn7Q4uNvQYi6jVL1G5qV3ZD8rLXXWjpfZrVP5G2hJ/rtFFszn1hbwT3kYpO7+
nWrk9hRPkcZ7dUEytbyQW2TABkIgUwS1xBHYMciqfpgRfcHbmpd/VBj4SKpU3haCQoH6KEs5e8Td
Q6eCGvyrsi6LuwU2YKUoeC9lLDw1+xl1keSsQ+v/kUlPDXQ6ayG3pHrC8IFEU8efSTW+NBBpXqNw
xTpqhd4JR4ioxd+eYFcZCohx1Z3s27XYyGlZo7cnx/ilYkw+lx7RLGNb5wkdd02fiN4rXBMKIAb5
yRJxuiPKtKhARCn2BNi690/qCqe7Q/x6NzE/9dX5PAcPuQCNXizIWqR18eukV6fasNYdA+jJgki0
T32J+weNK4fnKKfjymdbTGXuJMfvNA5yekOV5ZIodiIA9PuTtmRhbIK0SHZNyme1hB2cOmGldtBC
UzVZ3Ks+r7rKirwuqsCzOuVx3QRV6I7eyMSUJxSmDlhPTeqrVTWgLGUK7wZQ9ZG9ZdMizZwaXtkX
7fowJ+zjfIpGWaKFCE8yBaM9Yjo9S8bwNcIQP2XnItJfskOdoDR3JM6kLDAo5aMuTIqMYpk/z621
/bBLMPydzar6A3qK+Ecg/o1/EcUFGtpGCXG6E/UtFBVom98h0EehASrM/4Qw61WPw5YodJE07gjv
9i1RGBJOuU0iUG0NBN2oWVJDF58YDLFLxMS0CaI3kQPUzYEWSb/5iD3OIIeI1OBFv7gWkwXMv+kt
f4yOJDcUjLmHzgUU3OGXZVArsYF7+7YS+IQXyrSr/AlFmbnGAbExSBL4qWJ82h5xu2sqURNmqnze
dE+fOftPJFAYwoIWVP1PVNdr0ivL6PyUxRvmwQBczNO7ntaXaFZkkRp9XVBRV7JnE2Sp73VHSX9w
YJUItO2CmjxWk1PhID4ZdUIRqCEigJdlSddwhWFoUx6OBSZwKKCaUh113av0YSxPS1vIGfbMjtSf
3UIieEjRoN9fw7XUVjBxCnQdhz4L3ujC7plQngIDGzCrrZ0PWX6SOgds43ehbjPxjovyRbKvfm70
aXAfs8TW1dKZe8EZHOYm6PzdpotICIVyIE/DnvNO0CH9NHXy/lWe+LF+vQQBM6UfwyIQOk6aZT19
ougTpTKcT5jMbmkGq0cyjTeZ+HgsBb03bKbkKUGhUjl3t9zETnYI0LvgZHFcBMGnS0X7HWfjFfAq
5wXMRCyVBhJFrwo4+GDlr3NED6Jtwgug87C9Z0hRvm9g7yHQ/sxZDrNlDjkv4RxNGyxoC1KcHuZn
CjTEYhSv9q3/7NywPZPElwOOjpyrqMNI2fL7dY1GeDDaSN0MzgCa7HXw0F7jSXf4gCUGh1HXV2+8
I7T4r4x6iPXxenXSSff6wQodkHlpe6XFiuLWRltGAx6R/cVQaDJRkCPByLh24UsP0UhFiIMBEgMo
R61IlWdvKG452hZY5Nb74K7ZTwUxJ8+Bxv61WaNSeoqUBCXCKxr/5IQw2oV5zsNDOWOlV0mA43hE
g6iP+L4VxItiT50ecwGTT6Kys8OJ0sXS4wXHvMnb2MExpY0A/5kPX1CKxuyk4AgxrsXKjozU/CyA
nLmTisnYnQJRgdOvZVn5+FmPMM/9VKXyBnri84RjQuDMKZfwmSLBESsf4bW9eDlXCdBLgdELcE44
QlgEqdg5y0w4S4KEN+bxkvQYKHaX5MoJEs67KLNZL63EVuLzrmfiUeKVujgKTJGlDzaAP69AVduJ
+opfOMohR/UoEJ6NWTkMDdnBxF1BWfbpfuyidkxjzftjZqHFwhFveGQl7hnLayyF8fsY1lHDYui9
uwcCIR5jVjmLgSQxLPAgIK+PqduHc2a5gs/DzUV9CBg8upttkkAscVeP6vShAyQXl7VcGzI7eJjY
YL5wrILygjHjgVX9Kp+FiBEi0s6Giq7nGE6onlKMlg0c1/MR7wii/wuPFzyDJZrd3T1gxRY7pebS
x6WPdbSTNCOxSxrUBnXINbxConnGW1lLudbQ7dJbFUpKgSPZrFlZdl8T92cty0y4zZe12qtV5jtJ
6AJBjayL7Kd5Kn+9Bs+BRzi8yxdspJmXSFyxJJKcKrU6jmSSE7yjijfLuzOuvHI1a3YFyw0+uODZ
goiEX/0T1agy7P7FYjU1KwXZGcgmg+SGjLpQ1OOfh0cRcKDEoRqHgO8BUar+4ed/B5sNDuBk5Cpg
suAGM6k4j6F3+Imtb/Yr1e+VS0YWll0NkCGJBup9146JiwHVDwLUVcljZKBA4sa5HvVBFnOe/B+I
KhivpO5cT6c1sWucYqHmyGvdyTMsIVVq12qmpv8uf+i6SMD5Aqjjc1gzE42W86EJKpwgUP/Q/t70
HFjMCvzdtpnH4MN50iDtR1UE0Sj9C8NGs7eerEBV6eQBo+o2PssjeB7e+5gfO/iKextu8Pwwrf5h
BHWapjKU/hnKBUYPIhRlLBlBFaJuC01Ts1h8naxDRynoQSv5NeO4V16sH3V+zLYL3vmvyHzNVgmB
/Q0k8zgHKivHNL5Moi/FJn9gKlDqWb7iMrq78PmFVtVVwqiUUR8edRta45WmLzXJQZpNmxYsYOvO
JJXp7R2qsWaZK9+ESp7GbfjTxC7aQxxCNCsT1tfbFh50G5gpO/zxEuQGWZMPCK62U9s5jLApKCzG
vUKEuRk6tjcc5InxbHosnEvFLOk9tKg+aMo9Lsqb0awBESFhyfYsGjaXn9cArBuxep+B3Z8ixyd8
tWB/Z0VHQKaJbniDF3panZZX00c3Uz/6zXWcpcnlfwffmks7g6Z6q+vFTABcpxfhVTeE77T857QJ
83zKzjaVZooDI/20bv6BtAHGXYwsCc5lO/rm0195MD0o20p+GxIe6cWnD/Pfof0LuPXlMG1kw/9s
+NJ/IbfO++yJlj5GvvlUw9xtFuUAaUpYy5iZCxFzsVsg3La9Dj7i3TDhxltdKq4MHRf2RLZAB78U
D0pUkyjVPWQePTiL5jWMKHal00oNdl+/dpTYhDUmbyCytWlXp+4dldmoqNe9J5DqeZMbIjGwQeBN
2n2Rv/iIYeDb1pu4h5CQHMLXQikaPGczB/5WfC61Guuy0J29SQRmfHlamKPUlkIhOdYEemz+6/mk
+pdmiESOjbGth8bUZJE4zzGDVxt/hY+HJywqWZwEX4VHjU5dgSlL934mKnAhvE1RrNWndPR+iCCE
R+NVanQv+4nUhiG9fvV8rk+wGP2WM4dL9xnn5e0Ht5MlvUp36LKbKqTjhD9y+n9aVG4Spt6nxC3L
xwiZuMjmt/Xy3KJT/R0G5S4agej0hXnfl+ZiTaBxuquQuKpiiXcs2ZtuOhATxvRbgVFioa5/YZdC
6rBa9HP8hxTR3tytdKe+SenvVGTY+RpSIzNEh2feEb875AjeRp6RKL33ETf0BVPJStPxWXykenIv
Jjm77Zlox2FgLQYUZdsEGQejkRUnV2ZFVoFrgIrIwhdNcf4wIFXgLI389XREaEeWlkvg1MpsTrNd
K8jtNVPTnM7gK+UFamq9ybMuwJqJihjWIz7nNOo1+bUtlg2r3jctMbSNmQQMZu/UHIppvejlfn3S
6n2ycOzvvkbnABE+LgAvyDNMU57jVwBup0CXado3xmEuFGJMgCuTVa5rr7wqp5zI7QBN2elH+pp8
9i/wLLDv6V1KrxIa05L6Xk4+BOp8IKx5WLDHYxXTY+t5h/sgZdCcLBv+4SBPldrfCjDHSKXoVuZJ
JP7KzfJkakaDZOt8+jCRu2Sj99GUZCXEk1ag9ayKZIH91MygpRZ2i1MCgBNDv5iwagmxT5zEULvF
iJMMUHGfgRST+PElDj10v90ybfRA908kKk/xngJDganYsT4mTLAjRwTQc8bqTOf91rgsA0iFAKcE
1iwXKGNmoDrEw57MaYpzA8mMswoFEMnwgfd6JnMPJXlgKFoKvA0hUe9AOOaxOHDYT4/Xg81HazJn
5+Lm1prja/Kh1SF+oYLUUvUZ1pdcLay2Lvko6hm2ewUP24Qq0NyKeDvk5Bifvn3GyuMudcUTcQBZ
37nUu/1A2aMM549CcF7VxFalzHftR5ChcB0/BB7CWvmy/bSXq1WaQ5vYqSUhC376b0y1vdOwDbDB
cq/eFS436pkRnxZ5/uJjjDTHhTPfkoWjQpwc8GdvgRV3cvCIOXHxgUQ0pSmDRLHrBvNPlrjWKAtI
cI3s+nwoZLABOckqIe5Jerw6zyvRNljUbN3t8wPEjPSQ2J6WrKb1791k5XIj/QEpBUN1RWFXpZ9x
MImhmQUgpABH2S7WnEsbXo+3B1udYuNmmDKmqthVSeY/oEhUjSz3X5Vyy3Lu/MxwGzRWss2RxuJP
XFOFwCVIw5ojczXHIOToDh8eL1BTzxBHe7xJFxSodkq9O4PC7v+lqJZybJeawQEAHbgcPZwhyD2f
gVDNvVmBiHWiuoicXWs9Gb0pBxX391rm7UPX2DhZvaOxrMMkp0g4+Jm07N0tjDzg4wqrCiXY4poV
YuAWufNbyWWSTYN7UuZv8oPxucYuOQ7a8N+qCVHUkMefDHO1fcS0VQCM+ky7po3w3eUPi4xrFRRg
vNHZ4KXRvqFySTGCFPFty/+YMOdEEVHHu6lgO8Aiu0KJMwRyjMG2zX/ZgXyKYwgOtz6XHL6GDbxI
DmsbNJv4Z7e548MW641IR2f6B2j9wwVeSe3m1I1GPiFyBEXJmRecztD/YwsVOvL5c2LWWK38V8pg
P7aO8f9KiRLDsie3dd/UsP99tY2dA5KTXpRNA6rDXYDXrRpbBUb0pXKrc76+i+OO0Ajx2/AhKHcj
IZkLrfm5KPVJOzda8CDcexAHhQP6KKB0oqffjMS+gVj4+yWNQgSkaHcJ6LOlNho468EHYDZR1aqz
H/Y7tXov7B8++TMxJnIUw+LSVc9Ki6E2AjD+NvGdPcyE7zilYRcaMltx+5fjcvN2SnWMOKDu0kEk
9Oxf0NjqSipFfxjMfpYG8LIhmBUBeEI1vTA243c+Igbadr9L82QXfd5Wo4+LFK0g4ReL4WqS6s6Y
3RgEMbZHY5Xk8xsWV7w5yGGKm3gbe+tiWFBVR/sO8Htx82WZGF9HO1qwLPZCdUAhB6yheKEGBdgG
0QmJq2Pz3iO1bAlsVOfmozVyEqHRak2WHGIA3y+POmQH0H2GxshfNVh7DeW6eVy2ksmhVofLvbar
769SfjRS7oUUWSWa1rNNwNx88auw52G14EwMUlAzcu3a+u2htGRObKER9JSbcXPI0XY2DHD3N3Vt
oML0sfxn+OznrlA7PK2kKmSpbBbZw1oc+fwLkyLDbl47rt8KMz0hDPm1N91gIrM0Y3nz6H9tCAm8
TYMlbmsHdJRIJJAdqT8W83FT5wY8k8i7R1CsRpbAO7dVfeywuC69EBHKPj4Dxc2VAtb/AfhCPDiA
als2jfntbhZ96PpKdbFzEZnu78Y85eLmnIYRxojld3RWDZB2cqoHh5rW+xF14I2u5RhN+X7tZPGY
nZkfqWbCaTUgOFirj5jUESJHvkJSyYG1ARf15IQJbx6Fp335D8peFWOx33ot+vKkAcgKcZWru4wf
2Foxuw/dcmYjoTpPnj6f2DaIqlX+6LWxQsVsg+/IxwZF1skh8nU5PuLgDPttcFCZZWFBPVxCfk6Z
fo5Z/1jlQbpcLDh/VePafdFoZeXpdMzARmnrnwqbZj3DQDJB6WRGPJezF1eui77qBbV3+Ml1xuBK
v55N2G30zhHV2ipYg9MrVaWN15h9G8bbsf+LczEiCD+zy1M4zU/Q031h9B+zniMgQizK1Vpyd65k
E3MYDEMD1h2uSf+1lUjGoMXG5ouB1t/ZCPo/LszaRMgKMmKAYdbrbzfyQEhaZYPYTwdV1MsUVo3v
/AB76HJqW+Oesq350Yimnwxwm4eYwQtFEAJeTKSDGy7YcK1/QUnopMnt266OJCrZMuiz74eGcqeY
4zl5zO9lxa4u8zQEmkDRMVb76Sm/5HoklWqv5ShuRcErg3g7P83Mi4IqHxTVN8X0sx6L8iE7cA+7
uLBVp/Bz3JLJCki1CnhdSoS6Xvmj5LiRfrNXZagXDVILIB7s2O2feLBgXYJssUqBcw45c08fmoN2
suKsORURHwkcKGC8jSACzjdU6YREis8JmQAoWnIUrEoccGitJbVL3SbXLqS1s1Dee5D+usVk1W2T
qmmb9tvPPyHQXQipW/u6BSHDUsVjgyOwknWVyuli9xfupuY2VpLC3IvhjO+mLByjNkr94dTMEq3L
xKPjsZkpP5jCGvf+AiDjCa43PT2METw+VApkE2JSMhfswxfqugo5ENv2YmjSPSh0Hi0daWDxWcHi
zUzd8TTQ3mnzDR+qBnJna59RJbP8SaGNqb+TMK3UNhq2NE4Pk3HQ8kYMStawWtNExG0M85C02X82
0Jfq7VJhK5Yk967vtk9j9fxEB6/fpCQzgCiCRseSempgUaVG/+UmKVEk32dzbQ==
`protect end_protected
