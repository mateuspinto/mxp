`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25184)
`protect data_block
RNlzJorl3CMVohidZY8veno0KEIgj/jHTb0/Jn1w1/cMUasPC00l3VmVfZh0eYbkK2aD5iHgmU52
thIhbfDk0yWv6/XvnIX6KKMLWud6h2dSMWjVtVVTXZ5iRxfut/B4dvZOwDL3yGezM17Z2n9BMRFd
t8ZPlld4SdMMcCMLFO+DelrmCuHraFVGRK5Y7S+/bJOAJYFtEFzNyKky1UazwWNuTvA4nyZWNyiL
Ey6RijKXMnhKMwnnX1T08nm3SyI0omkFk4p5DKqZ/H2ewUWbCD5/K/QG+YbvBvYjzxfFoyIw3rAi
mVyLoPFit3a2+XyZnBV9kybk+bs/AXDPPqLn5Z7apgeuZdOFGpAGlUq6UZGNQ52pa4kG1jSAqVwb
QG+U8TRW1cMNOQ9zg0jeClN9Y6jyLP/Oa6+wB9JiwS7M4lbI8bwqodiUj1k4+ic/u1ENvO64beCe
Tup5T4GZopAMyrhlyv9bdoTMaFzgAKUOjSjdVnk7ZbhvqwiCvMAUVmCNrqx+IufLOB8DMOI8kFgy
t5KN6i/eM6EE0Lfu8Ve+fs0EnA8iJgItJZJr0N7OAWNqLHLChDAK/58dbArB2dOG2k0DUoBwlTji
wcdn+YJP8F56qfKdJYmJDib5G0Rbtn3oB8+Onl2LSeNnC9Kq17pAcMVZKSYd/ibqokBl7lA1wTd0
Lah98TJ7yo+fWdPms3RumGzhGaFHYRF6ZhIR4vvL723YIf9dS3tbxz2XtNWjpKvexqhlDGPxJ5g2
40GLCiuSy2YAF7Uyw3n2UaHAs/jwnhygl5L3E7iJzI68y7eKw4FHdfnLqIFZp926FzfVQQGQX8OJ
LZJQsWXmb5KAVaVIepjp6fV/5GRKK9BAlObGgysL3AV0v45PMJ5LE/goIq6t9da50qA/KQ/Ndd6I
5mEQ0/tBwBqlUNGMgHe+izvqt6xgTX2F0iOMgZCgIZ60T4Cf56n2EC3Ay7OIBZRoLhV6AF7n9w9i
Vc0jZXbR3e51nwl4rW1JQXGyaHgOnMyH/4ZFLUMoW4TeG5ZrBG66oh5nwsBrLj1xc0nCRcaV15iR
cZoh9ixeTpq16wqY2vWPq7Fl5djuqvRF1z5J8o76aPGY8poWUurGhynhFffZEIafHC+gU9u0bPch
WuoC0TeO6Vz6atcfo+qznb+0NMJg+Nt75AaM6X5VuRfplGrAZ2NnaF0NPm37KKitdyrArdED86mG
wSJn8LAge93SrSMjv06PTwa5umWBbOzJyfiKWMCrgONcRY7Feu0O8wOFkyowQtv9M9+ioqTazS3d
QfCMl8ReVlCz+00dJWlBvkFYSaWCCfw6Y+OrtyNn6JH1GDMlXELsQM60VuXxYDPSxuQqesgjtdjM
W2JNv5Dv6VRCUPNL/HEd+umWQY+wV2CQaA4DUEDKLC+gQEEbzB0U6UA8b9Uy4C5WiRPN+GKozSVs
V0tWu6Jc3kGvKZuxR4jsrd6ymNWP1j1s5VZvKAdHDfmoLKhWw187KvDePXdWQKRONk6UVoyhgvE5
YZ58tgKYmX6OoJJ0NoXulLFU7gFTRpa4BOQ32jgsK9EYiFDPsSMSCCm7Dp19esfBo2PCcbbrEUCU
+eZinc6LT2HGbrPyXvVdSATnkXiw9dEDfrGTkC6E1w2gtc6pQgdpMfwK0fvwTY8cIDBz3egskLpP
DttuCg0cSAIeCASAaY379Fyu7mcxfnellGfg055APSGFUJIdw1IhJJ0bLL/ILxP0tROds/0lliF8
uTvAyq0d0msoeox1s238w5JGulHOS0EIO1ldHLb5z10sRNinzApvx82NJMhu+WrSSEufZhLXpVET
myZK2ExyWAa2c2NPojVRuY1G078hQgNtBI+OB2xvYnZDBzpi9u9ngEkPTzymypg7ZDh1tr8nVPyZ
rircNRdSxXxvwiOROuclGMdYV12BWFsNVoPFPyYaPsSG9LB8HlwJAezruw4DrOs9Z1GwfP6o/aXi
mX1tYpvZvH+4ZN2gyBIUZKevY07EyX2bIk6aj3I5wlwXM9k9FuscLQr1+zubsbupGc/NDQkCE64V
d+Fd94KK34USsMJwW/fmFKruui98xO+ThkXFFsaM1qZ2ot5lELr9j5Utcq8tgysEUgOWJpszUfmX
JjonV88pljSqUnbJx4OrHbG24PlJSLZUS45Nvkl0Z9Uuh+lN7FYvrMkUWVbVcQD3iUKwCU/4YWh3
syS6p0swjdScwEOWdRmFGlgh/Oxl2EcYzAkXEGNARSjdlatFcyQ/dfloplXQFgSNlGqNqSpVIEIl
OMa9ufhbltEEVuZWUe0NfvaCPAv64jFjn7P8RwYhOYZ4Ra/XDDow2Rzeys9v8wTMBbB22+dL7qRE
3gz6hcHY2xU9F4GcXXzWG3OX4iI5nUM1IDgydGN6hlCkyU3M/4da7NWz9c266szfZHUmD+nQNic5
K4hOz9do9Kcw7tjOk7QakRtsVS+GugHJWTmn343rLT3S/vUqD4fB5khS+M3PEJn2K6MWatq1a9zG
YVrN+F/1R2xWAD/5e+KI/E+qkWElTB7SCSfLVYdjWTT0XNG/5VSEAg8M/DvzYJl6Lx26IzRHsWoU
o/hqcNSLPXmupQ5LCkd2WuSye7dmccfPNukiqN7/07UreCU86HaZaLiNhSzqyyM9SLBo958oOpZg
rcw4bTP42Ez6Cmq4c8vASzXsWQksclIthRSjhBA65WATlaoY2erW3rAEr2bNVjmV9KIveRmvM4sM
vrjG0tQ26n88HasNQp9WNm1vKXHlkGaxE1CNSHfSHy88FG9bYgLlTxsbc1n0BOE3Ckixa63l+9xP
Kr/IsO9Iy74o17nBggX40McADLTQOYqGdCapJzmOUIeBfRLUZhO3DhUKlkcEDMJOZdU+LXJCjWqC
CtwXEZzIs7qXwkE0qJunPZAPJSlisiF+fUrVTy9kFg0HAnimoXYzsz03fpBb96kgrbZoZE8F0qE3
1mx+0bsOAx/cbGLLTb1nMSgKCuF0oOi+6XctYAxCKGqihDtnRifR7X3YasF2qdj6FCJFMOyMfvMi
ZjgVd0wBN2MPBWQK06aRG4zoEqMhywb8C9xcuw61D+gob7JF7gLX2xz1KTOcIuRLK89yqHBJR8KS
g42hKKKMK5XJP05YTTfjIYbJtYq/WD203862IIiVzkljJKjZpuqiUdu9ziTNwlK0GroKfoGaccu8
cJDYPkK+3r+1ynRFmc4jCp8ccsfSg0dLfMvSvvVmNuCH6J51rqtEkmAM/gEabJMN1hP5R99DQiyC
2rgstcb+Te3DksniIM+NO3KogSd1lpEJZgtjYOaBkVwTpLZue4BfBmTBuowb1wh7/9/WNDyvbN+a
ngxPIwcTT2DwlLBySx/KVHEDREDFThHNXKX/8Gx4+od468+BjbKbkGYweCq0siFadfzmmmHRT1UN
lQEm/9MkPG4W/UySbQzxH/lbJ3oGtBJypp2ZjAjR59gD1I4/ZGjOPPQVVDVsamTILPZXfpy5eWiw
FlbYPUaZLbYSgEo5mKOZ7MOPDYENRhA4F9EYsJGvvQhhlfO4RlGsqIuvqm1ko4FbdPMyh6pJnGgF
1LLQwv0MSzsumfWwctf+ax21LjX54seRa3eEQl7lN0V+lHVNT1SWR0VZjL4mSCet7NgLnbBjqCay
X12XGRai0AhRRhU+CVR+h1tZNRlSIXOMezupDfgYgRofdvetiVrWTW7Xig7Fw8Zue6XI6WbN+sh1
RIBfZSZyCDpzQ2B3Vke6rkoCekemTeDrPk2L3qOkgW9yyo29r7LuWksimdt7Jj/5IATihz32KE/q
othQpn9WZr02P4JG+mfbKg1I2krcX2rCjDvQwlO32Mhi8TD2u9U7nHCSAxhnWc/iFDQfBxkBSjGv
Aj6a+XiT6bbQIBt8bsCEOjpkKEIIfC8GSC8lYh58vkoyRoftHXPRImQ6CY0Xm6xYi1Wp8TxA5cLQ
4LIywGW2IYIC2m8+gUH60ycz7LLfpYfU/mQIptSdjwbKucLfxeg0AMMOMBid/kRycov1IbbmV44X
M2QLLHtEdhPNqSL7HPRpi9MA4Gd3dAdI3uBlBxfXpjM0dtq6io1VgQpIpiFt+cIxXcVvS6pxyzFJ
e7QbGBC9r4gq4fUhWefrodr/MHtxtcjUCh9WeHBe+aa5qRFMGAJ0yp7RB0WcS6dopxthnMQg92ST
zpdYRyxZH7+6sNZHtqC3gRWBnPv/ErvcX/vNXUVDt8zhncTce8LkFvGJ4P0qliaCoT8T3+8KuTmA
CcpK23z/sPjGP5+fnuXUEXz+cvwnCiYvQ6+hTNPAJTpFD26thq1lACUpWBVYy5Zu32TyJOCWXq1v
Eo+95Jc0ih312X6p2mgH9lbKcfzpnhr6/+X0SRBllKSgIncira3CSF3IQdCaENWScr9IdWTxiywW
3plvciLkBYBvj5pkLDxp6bQRL9pkoWLrzss4EDlSGVD99eD0DuvVJG1FQXvBrIhzjDYnGy2J8cAi
Oa782+W8D2PWdlcFuQQaqQietwEFL0c5VKjJ86ZoV3g2NV9/gm+rR3eLFHdhDkHBWWGs9Us+zo7V
lsTQKsSS7bG68eJuAMyFZbbDVdR2rxorV7d9xwZng8CKJn2zMXOiSYNKvnG3JgaOHr8YPBuflSlO
DeHLC+Uyn6FGLDemQsdbO67OzVg/D+nptzF2dYJfrSAlVxv9HQsc/7rrmqOg9+3NYuA45tke7ukY
v3XUs4jAgZD0RuY+uvbHNVo8mx1bPmedO9VrbPfY/kRj3qXvwqsjLrJIcAIzhbRjNi3Cb6//ep6Z
T7H/j1rYf+vpbOd55cbBhlJI+MOvlKWdwCdkXa9O/WkyJn0eg8cfogMxhA9ggE++84ULfcn2oXb2
Rf9SSg07un6rYlop0gO+U+Jy5H7YWuGjYdKBc9gRDCeQOTSnHQjlwGpaDwOhNjMBcuJc7eFqNrnC
eBdFkq6csRE8IbSw0oQQMiYwQ5yhRxpavBrW+kM6JWC9V12QMvkwoJe20KtTwF9vKyoc/zTA/SyH
3yC0bNnrhCdxz4UP0JvpH+ECcfEnw2ZPK204I1zQhAsIz8nW/QHmyCY769dghjV9QB6jUS7u8rkP
HUmsLReh++plHgD8YVYbKPSh+X4261yRe2zsQ56Wu6Q3qxfZZ06HvTG5qLJd1RRLDw/kr8lModxT
M8OlSexLG11BJuWFuqIQwAvos1Fv1YqCVt6CCybx8kNI86b56ZGK8iSWSvbRlEJ05UEfNtAYYXN1
lfunr5Y3MLfFk/XixaI4lhF20RMOcjvEXIJx1Yr0x9VERLzSTtgfeJn8h3q6YMc/nqrhcdmIPHnz
SWfrOs/+NXPBqfPeZEICaI6fXbxs700TCa6UaBFOqkFi33DZ+yh7kIFRfcWxozbyqNnBgENb3Mt5
/IeV02TIBDmVxPZalMAxeH2hqZxsBnWZjU1x5DydzK+Cu7+RFEGdb+0upTqYz8IKIePAsORGx9v/
c7EeEXw4ueRFKl2n7WximZdLyPePNPqaz5auKEKfRaPDAw6pWnXnqMswatTP/BTrEL7ALEMJpbaW
kpXiP3tej9P2hpdPBvmc8fJnb7zVPPI5yP504Kefmzgvw91e887oEugXpeLd1kyE830SNin/GnVJ
hnU7PR0H/g+37iAYoQwVsFLXcqaMZvcT+hknp57Ral2MQyIjitmTf5OFjpAWDco1luw5MKCLAsDK
bCLZaZS898xVbkZYdiCxW6LC0UXOK8j5+0eFoMUJ/lNWG7bmn3MNDtyhlg9VSl2QVVvhxYJ+5mac
vqAwdcqAmR/X94FKhOVKekh9d1xDLRx3ekOt1wGmAg7rI9lh+Le7b6XDwejiltL+tgGwJaKsjKDj
cK9a3w93Lgl7wdUxH+buF0Y5nqKb04JLROo1iRZpTgYRWMERiJY0yF9tL1G7S0wu5wZ2AYVjTyVs
BtAEuqaytjoD+6GbgXqiyyd6WylH1wkjgmgonBP9SFJXRy1nJnrEgSuXZyXdx+aMZgrVDX+Z09BV
55YGn4ZRN71m5MaMKC5tM+DsGo2VUfH09cyDT4vdV+QFyEi5BuLgB9qKiCyC/2ylCwcNqIvtaXk+
7s3+v+lg+nTv/+6Po0GvMeVqTV+VilFsA9bjZCA8+UqFPBk26l0BbO07dQo0Jav73N0aS+vo0w/6
qon9/piGwkbMIF+fA2HVLmrgDKcIIMWiz0JTg/JqsHBatzHLio8PtPc+wK7dXRRslRZoQQB2QNNw
oofwREwCrpZXfb7MkcF37NYhWc5PzIq/KeS7kWJXn5pJo7wakILhK+7Mnb6z3Jkb9JEOtOTfVB+g
QxEO6ys4H6ZC9tkK4Mn/XD80pcN7dWV+fjngGJu4qgS5sIsmnUte9vlNYEfJAylBtO+PZEB9Bqgo
eN01N7MNcdRTXWurGPMyTVyXtNu4CPcEp0oe+Yyo8esfHwfoBPCCqalEUNMQPlU8N3rRXeWYlWhP
kL4N+5oQ9/84Gm0CcTqffkbM5W9Xfv2rWwA7ni13KKjMxhFXd0bHYAVYrMQe9SJknugC+f++zW4f
xXCaTP+TDF6mIYQxEW8b9SkwYdl/qHun44O1ufhfRPV9xLHzpK17XnFBQtmVYeFx1RI4GrbxRK1D
znQeheh8YItSfcl7Dq6DqQywETF9KbvKlITE1+JgWYzzUMPpDE11xJ0iBLSZCJEFxm2zk1YLDAi2
G3Icb2lALi8lX61BShxoZCt8mHHJTgwQt7XOQ5cmNWHd43M2KgKMD2eLbY77N8+w/RyowpC+Fgp7
9t3x7ZQaCfpVPkt9MKajgMO2KLtKbReU1xgx75ySDLcTrhwYevQBuMxTim6Ni1wkrhbiQJ/b+rwv
2mnbm63UqUH7Uv60Gz9CDGzcg+0jgxw3NUywFCmZXrKhQB6MlzHJ3gKjo5j1L90pIv9UHSS0Scoo
CnskotwgPO+49X1X3JvDuF+U1IUbrARdT5diB2+BhhXfz3zwwgMBglAK10s5piP45/6k7VMaOtot
2S9B7C2tmFt+UoekaDaqveyGABKKXcv9e5KH6OiJv0aT8aRQ55T58pRyOVx6DZ+sXBLvB2yL24kg
Ma7kCZCFNBBimy6Uligcbi81H6GC6Y69ViedsoibzODpOsjbURRNhlLFMCOiHSzkL+3rSbIiev8E
SyiwrG4SjpK2SOT25J3S9nDfAlE8hRrB8D+MdRu3BO9WjCuHezwg52krXK9LA34C4Jvo2PSDZonw
W/mVh3bNi2pX44KFHnZ6VKPdV+JcdI2WP26Tehmk2EzUYFidFRa1wOqkU4k3hhM1FKYaXjb4KLH2
5CJ9AJFpo8OPNuQObgWgFHJla+kdbV4sbe2aZCn3oCwpAGowwGUSglHEQQeaCuRKbHkf0Gjukxp4
A7m/PmtMxgaU9eB5cd8+X+PCctc03xiJzHXkTmUpXINByBZhDQ03PD/q4Xnd/Zvmhx7bV8jEIX8h
r7SIRkfEOiqFSJVmWzZc/vyBnUCf7T6KtvReY/4QoHhgSDNs7DQY1s1WmUACjC4X3wFkHNSGQVSW
j1D5nu2uT31gRBndaGqZJsVGVze2sHpuLi2+GyWFxaNKBLWPPIuvykDTCJfgwdl90GBbgI40BnuO
aG7YYkZhTdZXHLZsgqYV2qmO+B28C3lHfx27yLnWbmBqF3NyFyx3Ysd2WNV1V3Aq+DQDw0KY9xlE
uilu7ruAD2uwEl4hZAmB8AoAzVPFzpk1mPRA3hBvpB15h2pCveCLbTJG+5tlgXoCPWq1EUyqqbOn
P6vDEzgc9PlRLG6ZOty6wD+7mNsgnMXa0FdKttd4aXjOtp+2cqWJK0e3JrSSJqMx4X7/Y+n19zcB
wcwwX7POPaf4JTE5uLMQ2WjIPzwUthLt8Jswb05hO6EO+U6k2Zh++3ONYbW5SebbWjvUKbRqC90/
YWeibUy1pbkQckrx4teGHuaSay12CnQM94kwSgbF4g91xKTXpFyUvmnrZq5p3LjqSr79djTCYWFU
yM6ANuicIkGJM546oAkkSNFfMyu63jbVoKUdoY+2hbAg41dCD33jkOgBS38R37kRgnqHVn6c+ahy
jNU9OFICvRruVf8nVrVfQVuphhyzkzdePjJU0kPHApxYa0Q+iNbs26GtBB9W6TZTU9YVei7Udidv
elzUUxSyLL1o4UPfVbbIJEJJqYJ0xnaY25PmR/4L97Ra1WYvmaeH7oJOngopS0r3++JPA7rd3mao
n5PI7SAQVFY50Yx0/c0OKEy7g6/IUcrKTdX7cv89S8LE5XKwUfiGLN77HbGglRyDlCQQrq6wMuc7
CKrM1kRdqHMmp9wBbozFpIOkwjBo0jr9YDvO1DBRJUinWBAmfUXitqoDvfuR6X8McFtqTtco6tvT
Ci+N7DG7GJTmx1/PKW77qKlirvcaM1wLnhD03Ds8HFxQIy8+N/YU4tmoJDn54mbNn5OMyuYXcXgl
ze1pceJV6LlkvWSULpVtR8kjZfd3lGryLl3XY6rcJK+1MtDokZSUUfmQNFYfskzNV5gjgRaTIdJt
TzXvGt7I5/pf6h+hxN3swgBXMTxtzcq6HbdHvMi2c4b5gyTS6ivseIIcCVtRLekQYj599YooZ971
bwuKPbRTYY7eQHtdCslfbdKo8bAsQZbPj6eTQ0TVsMMWH/9PKQjiDGSZrcmMTs0mUCNhqtyC9xQV
zXA1zsIr59XX2JhVLoj/SxA+YWqV33k6we3nEqwssfjgsNZOyeGPc5Zk0Ywy/tiBT8fAx+Uw40aE
QbCDGwB5GptbUR+1u5yfQiZVHb9mvANzsUCcCkEX5pbNzejCJEZNPlEnGL4PFMRvuP3C63tNzv7z
Vw0Xr4+7kPyKwa2C+9uipi5kW7sZFtcHeMzqHFNUuLZdKDtIP0j/8k1FcWpKoty1sosAhXbqz0ac
OPAi0Yj9uAviUaNV7w9y4Oi9c0qAL1psHvgnUIa0+SdOU/lrT/gsNyRdwOgNdpg6PujUq+bREah2
CRxgrnQhMgP1jtY83Rwvvtgta4en3UplkmGQs3z82lkMYuG/qQU5hh35U376ZHiGaBbQm3deo3Wv
h0jzhZksGuN5/u4BON3YOqeBmkgSwsE9kKVZF8PwR7Za3cHVB7iGCpEAqlNv/R05EzcPKw3fPDfe
OAmuNu/hu7M/m1OCo5eEplkFBKsFonCrUCS3sU6UH2JrwU+QqLlTJjwBXmlvZJIEEoWPrAb2MZrA
jtRBl3CFCvKRonWlmQ74OK+FCaH/WvstVaTOY1liCytFCBvpfz5Gf7y2LU7PIvkBbgSbW17xFsXQ
qa3pYEkOI0p/FdN6CZxNU895yACdiHcIN7fCaUhs/lpoGTS7GjacXOx3hDbgY7At63SfRf43Eqdi
cU4Jj1Cb7RnE7AlHQUS1Lar649cX5PU0nviZQdiylJ9k4zp25VrUZaL5fy/MPYVcbNUiNBUVWbAV
NlNIWmSIukd9pq/Tyg6C2oWkK4BBjjHob6m44PoZVn7VMngUqwxeSa02j3Rbusu48anTT3TG7p1K
6pEvzk1knyniTeZExSFLdCnesNudwQ4H9XWDVLYI0Dw41zR9GEPPifBTRz+1+s1AWmwzxOMF/esH
sxrqXyMlexGWqnfFPSUFC5lc1RHE9kM/53YwgnBNCJO/zBVg5V/61JDYoQVAwh/eHNX3JzqNUe2M
XtacrV3B2pbNd889itL/TkHdMWUY7kv8mEeJXGyV9EfjpUyLjwXS0MgykCX35eOfS0ePdqUnkX2w
Gl4xXoz4LbLNuzZSxJrlW5zL8MwRDOOZS0sWnjlOe4wa2PiroBgV1YgBGQk+4JqHcB1i5+OoN2NP
mfhO4iIGRUYdd4vfD9CfHuQkDmTrB2jdcZ14SEZ+extZthDBdZnL93YvX1x+H5KABTXxdzqFAGCC
BCEYCKMqwokQXyWbFvNtavbhG7cqKLeNMDChlmODz9dk+mQ2NuIUFYa+laQay5GXAWCDUeQfFQIp
fqaQNr5BAMLLK+XjjfLLxqTAooY07kXN1MZK7+vBEFoFnt1lUG8x0Atf/Hh51b5WrGBrYRxECZzD
pGmis7PTdNtoJhC5zA6ySlCCBEgr0B9OG4yHSW21ONlk+C63LG6papodTAx/K2Ar4fp/OH1Ffn1t
MDG+yILJ+I+Eb/sLl0G+GDh063JfRf91X2xRwk/KbZg56p9KBmFJH2Fa6ApEQcXJR4Fj5xkT7WJA
JjPHMy2q3AztajrqvvnAYT4HX308neUH8NjpdTuhak/ER73mCQnhci94g/lc6RLn5XrQjhMUO2ts
8M90Otk32otRIvoJnyoNSYDtmCXdrH4eQMuLSnK7cDw93iCHTvkD7WyjOMYvNnA7jLYy/eOPKtBZ
22cPMQmRD/LZAloHuMhjbkdRQZxPuNKXw78ZWP7LrIEHefZ78Oc71axiop4O3IIKviLoyk8UsUSc
ykdhfh9q0CUXq4/ZM6HIJGTqTFYahABdrqwoag7+4XV7qSzI+/v9CUiTXCfhyVW5n0AeNakAmxZF
UC8DOA7T9pRMfiq22y6se/7+OFmebRy4+VD20kSe1Mc1t0rhT0KcW4ET87TzGojPFuA4bLbHAhSw
VE2L5n7jtyTkJNHA/jDNOiqYB7B8M4jtvzFhbQgKlxXXWuHGlpi6Rxc+gNZCS70drjdcNdE3/XTM
0DjatS2RQxZ8RFvNMV/XOFrve+wkQ/iAJVnbB3SQ9PPA9G+NaEJsxDbfqa4XRMp+8sezQ9dopF6a
S2cF4YJ3BoTt3uo9pflhhzKpcSzl3YzGhieOjsfePYOsqmcTeMtqAQdkgC4HKkdhJ+6yWOt0gQfe
XDLibYXvy3s+g6ClqHCOo/KpsZv1+SZq8UIHPwkIMb+gnIl1KLCm2r+UFdN6DpsW3j7R002XVtuf
MQ/M5OgSuEIHyPnl3nhu/FCElmTtx4akQKfHL2zaQktoY0fPYwrRFIaWhT98jdD4LVfv/yTx8sds
HNgkSq05FfEOJls2ERDeipK4QC7EzoHiGFHMvzFcwfQzNfFATQztkwiIhgdlW+1pugdJlVvuQgZQ
Ni8NZ9vArTPOpgwAZ8m5U8HZU/DltdwG5LF/Y4S6YcpKxL+TsJVGEyJxrfil0lDjqdWANnTNt9yK
U7FmJQ8hW8KcRgqBJveoQ9EmAAoeMo6LWXOy88E08hhtbFBy9rqn05+YVl0aCkgCG01hUVF6DI9i
6hWmGf6qy7q+2ri4vXnMGibuGYuWfiVLXu/X9AQPRigGBIV2c2JB7e10fkDYFrsr2P5zddV8uvQe
tdddYcoFJd7gORFZmQ6+PhwkUV/P9Aha6rYSTnYJKEvOhxnD4JBBK4+6RZVoTOPhoTHA3EPV3QH9
aegAkVh4lew3RJQIAEx4zG90V6JuEwqJpA6uMw4O5h5fXsxprCviPRd7FSqYlZrbXKUh0BGIPPDL
N6ifizK+EJQ4eZ9k/WZt5arp35ZziApT7eH36cjNwQ32ltx9dCu367tdieVeYtj5OWRJwyHyHFXr
wErm1HObyFd4/V6Fj1r1AC1ZceM6cIyKodloD0DDOHY2suAdhIT1QuEIIzuZHMccYCNffdtcFSOa
GP+T6Qn9n8+tiVk63CsM92WfHtWu/ajdT9Y6fFGwu0lzUg8eZcYevfWJCfe4lMNVG6VdoO7i53Lm
5daBIwoyznvBeRWgNYC4Xpbkf+TpqV4R8MdGMDhvBpVOEl0ax52jsSJSDzwVLtaqKtW7jbv/MsHi
trXeAXSzcChORt4CPapfukOpI6djcxzguIqhmAh7cJy5bkrQpMmGJ2b4jUFFPKF9eQ94ci5kjYIE
4e7I53xQztYFBAozdoEyynJDxr+an9n9vrlhAEOD0kK0FHQVIXoUfQ9qtUHMBbAQj5wGQPM7S/6b
wCexzCJnfqpJaDt8hNDhxumrzdfux0cGk7FGCzSblxjuqLuRlrZQtWnMe1kzTm66dllkcg2RW4jR
guP1bl1fD3u1M2GAyWpgPK4QsGrYeRPi4FME3QGLggquSqksTIS372nk2OTDY3Y95bU9hsmBZxt8
gBGjb0rOgwH7gihvuOFAzxUOkt90Q3wWgXSVDqGVEr6NgBMQvPA0UoV3nNGi9uuTMF+waMG+6veB
lVk6vpyhArVo9VYceCSliRN50GykzrBcqzXmF4zUBhADMKXF6d6PuIvB3y/wMjWURGXhPVxV3BdB
/Uhb0W8/k3daE6tV2RuZm+7eDd9oYrI62NGryKeTqQm4b5kmOFKT+jsTYrJ1uilMJOkpey8cD6hb
vV1hqK2W5nxxlONvqBch3zqrUPMwdfyoC13ggmVm/ikhzGDkIm3B1/cZJOvqewTc7ogFDcVNl71k
MsTcmWkoUclzABH559g4gcNAqRyOo0oti/n07sdv1H+45YiEyRmlF+2aZgcR5T97RUoYSrMPGmxG
OcSYUX9ZvUNJdBNGwYJO3FblVB4B0JbofThfd1F72XcEucq4NIC3hfT2P9HN2WVOPD2VEiORAlI/
ITNw+kL9iyFWxA7/WEbjoXwh3c2KuDEfHiYs04Md4tuiBHG/LV585jrOGGG7mkmS7VVTGGyZZMum
N0/99fouK8k48oicAeWkEnU9BpYuaeT3qbjqjJhV8bBLzdijObT9W56dshAy4Z4G/0SZjOGq7l81
g1/eMkhZoH0TXkag8Zb/7y/Fcx18+BcRYu8fFkosMD7COQmPsb5ZpXZ0Y+9tfyRdX9pcIgoo4mfk
Q4jeBe6qLZWQQcZMWknYnOJ88uSx7vM9yalJ6X2JLIb5/5CLPCyFH4YX/gnVpdRLHdLE1LkhfPqx
8WzhtKx8YsV9ipQ/LFRzHT+/HnddB+kKPgUJoKIVvG6SG+X1wi9pCX94PzGv/fRDNzHU6+VTx3VE
8NBHzGiHnL+gKY2WFxn2u6CZhiYfNP8KK3STsHYajn3RZ2H73z02C7NL8kjKbwFuMGwpgVR1YAmF
JbxcXTlAJ6pd27Z4Xqx7vG0Stj1wEcNdXrC4HYJ4/zbK0Ppprp4MlsYfpHVUWmLhZ0KsUZGfPPwS
Ii5wQDPnVVPKfl/OFpd5AGD50npn4fFprfjKdb3ICvsW5I4iJFqD+jAiGzHjcgyazh53KzVQ20LP
3jBQpD7fDL0VpmRbDumzaMQxMiTvrkyCx+wzRi6l7/czjCGE+VyzTFmXEXbh5OifIZJdJDZEpYqu
bWYTmsLnWatO/mdNHB3162etbyU983YxWVnFg0JmrgRoyTZnw52AwtJsueyd3lMghF9FXiWoHqx8
Qy3+Hvw6I/HYnqdLOFtAFOakTuH0vU+azOvYuCQzGQbY5vCy4JG8/YBDi82QdEwKOWZL2sQIP5wn
MeQVMeNiozy1RaaVwkJp27nc0GcTgqHwPbIPCcuLz2gYIIqtmsP6vhu9bVdYs0SHNUhcM+DR0mkt
NC+TZZoI4VOdLjBcCpZJD7nB2WQbBZSTScshqodAg6SJJAshg5VNxxRzu/0VjtXMSmPQbiNFTWNi
OYAz2SGXysFMd4cWUhxoaRe6R7CnB3LjnxgfejoUp36umkb6aF+ZQWF60uuMQjWw0V1C7+QMPeWI
KskaMsZS2zAzb1GI/aKpJDBTj4QB3SPVFVfk/hKe3IIUHtDCMx4pqSe6BcynbXGKFMTj2X67LHdb
wBRsbyVcA0mFy2HLn2hlM3Pg4If9IpIWoNI67MtMJ+TNBfRqWlR1kr99cDsmiITKguuHJgKrZRQ2
lvzH4q1EFw2A9X6YAJ2/4dOtCq2MGreyRnLQenRSiitvXsBG6jCq8Js3ZiMXLFNVhStYBRPM07DT
9hgHy7kFX9faSUiAMm+FjtMoeKr5BdUNThEO+yGD/bF/lm2q09puY4BRVfCoizSdG6OXpIdF2xRA
MQ7RZghH/+ZqM3MkkPYlIsRTNx2t7X0QkCWoU/vdO3sCvEooCDFkGcwiaUo8CZOGCFPBY2Q4xDOK
Mev4r+gd7Qu4FfrS/nw7cNUQF1PwyFwleHmy4wY0iOW6Eggm7z+r4dBPaS56iRwNeGgGkrwecq/h
ygAmxjCKxY3X5eanD99iBAEUmdvHq0xYf0bQAnVLZPRbPhmO+qsVNZeTztseasHhNZ03bvrIO+GT
/hqrqxaDdjFUKtQQ6iiT+MCa9HF2bC57x6fKIcEB4sHrCZc2yv7TxzH6kEj3mO9Gfl1B3dFVrIk7
clQRmqoV8aO8N7oMvDm3PN0VuzKZURsrGgyHoeiAGIwfD79jskrNDmHP80bqrSrNTTzdsq6Tc47r
2nDikpzrZEYc78XUl4RuxGpZOV/njdtOKZwO2dDBipDy3/mOcWhpzZs5UVxqS1Bc/PTC11E40oEw
3SHBIY8D/CWDaI8OjOaE7x8y3rUx679bCh3Z5z4JOyDkJdkvEcz1X8+a3wo1acepQ213T98EvMam
xdRxddWZi52TeSgmuUh2OOgfW+zo3uP9rpC4vmAQ2CcIpwolOSFjL9m99MvKT3cQ3Hsg8fcPmS1g
nzC6w/5TXHm9MAZsYZaJSj276DA5ujplWF5bRbfqwWSprfG1HBI3ke0JbMFBrBRbHJfSIjIaWkyd
lUQS54OoN4HRUQpyk2RlS8p76eBbAkxztT414cL75PpBYI2OviN0KCbfIIKYigshImex+sB2MO/l
N6YpYcQus8RjR4a/1BhLgp3til1n4FHuMO/k/EPBKMNXZM9Q9OaiD/ExA91++VSHfzm+bjUTQkON
c+6vwydn0uLolFtnBQzLFmrLFSWTmFmf3ClksLc6OBcZ7GixSA7tCvRfmk+UcjjLkH92TSJ5qG8n
tNZD4l0sfK3RW50QTgVgsXNcxRWfOX/nYNE8+/HRsCH8Ge5PXFV5nixNaBTIIolOISLpD59XZBCR
yGCgB1/agIbUK9vMm/FF3OvK3SWHN3Kay3gVIWK6Gxz1cndgNnXqWpbt72HtutkviWKuPkQai/qm
Ha0y3LxVuC/zaLVeOhHi0+MpG2aqyMYu1a4vxnokBZGXGRE/xYZx9pAdDdpxXe+WAoEXCaCh8/5V
WKF6hZbAvbaZBcSz22DGiS6QXyXUhASqVfLb3kUBUdkfpNZyA/BaQbwHDgbIk+SWQfwBX0OulkCX
2DmZVZ6HikuILYsgTEQpfpP9E4eRoCQ7iZM02vwRA7f0COjI2HAks12StQvcZPquGvVeeslNsIL+
VGSleIQr/ipnbvzMkmrz9Ui40GIdf8E/KVU2sEprWnwjXUwgF2bbxFdzbQqTvQvmr1nsJiyPwX6X
/v1IgNKUlb3RROegpsROtlBQNAggS2XcEJ6qHiYy9tGShtkSq3HYVxYKDBJzFgDTiiSwrSZzng/X
2tMwTP6Mro4aZZxRIQjbx0w3KaNHJ4lc4oYQziD1IALODhtvcSiBOM4YyUeNMl6D1L+N7xkZk9QO
F3By5VGBaHvjRtFg5FpS3u2kf9Gz4rq/+yWSjkJ6KcgVu2+VXfGgDX5i5BXsP3z6B46v7R0aPCbD
0tTZhg7guZxNs/ucEsfdfsZVflSU/oZmGgtZ0vp0LynyyuGZAu8z4WEbonW/KvEPninPPiciv0Hl
aH8aZzKofhznbCVW1hWuOEO7mZnFCAjggyRXBNpYAqii5IkpNjnFv4H5ztg83jAhMwLkOyxZFlKJ
m4RyWFT+Mo/chRwrX7GXNFADOFmOLgNGRABj+Qp4OPix8MG1Qacm+oHpQKvj5xYnedSJYtvjebwm
X0dUpuE0sKVgd/U1yD1l9GmCfwgt3EBIlBDzu2F42K7fu+yp3Qp3gSnvKDiJgMnmbdXYbVlNm76a
btX5thQnhURxhSrcFNBeC3fSD1BzwTsl/cpIjAVsurenq1CFKEaDm5UESsnZ5kivgpKIqAM3FgPT
S3lbrRhr9FqeOPJm2piPZBzHcMnRfKug5HfJbUHTbpiiA/jpZCB0qOXgd9QidoZdZysNPEdz7AK6
adz0kIvVMexNzUzS03uvmBhMKGYSwgPSznDuAECR8Tmte5WQl/W6ESXlc3HOEi5HV3gPoi0+cVby
WuNWIkms3kRXDeHcS0xp17WV62K0X4OQlKhjpMHZ3sWnpJArSgGoQ1yLaZjdtq+DuyaoYbYUVWGp
q+Odo5YQDWhUpu3Lm5MEiw4wM32LBB2P9fQvChdfS0lAfY1BmCEe148sJvNLKq9bCd+X2qPyVe+a
nMKwpQGIGngwufvVl0r1fxC3pxyiSEClL4vRdhA9XqDz28ojFsm+G8g6uc9cAwuzagUkVDF1CUv4
EAjlGywWjQHmNVBvHvmm1+Eu8c79TPsyrJxU3/dVisCsbufO8cNUCfDhnZesPI3IFvGz/eL1PgqM
Y9PTmFCn3gcdBBCBe6tseIbbLWvlQjXiTsouSnA+o605itKppNFHWg5K+H52RS/xK0h+Yf4J3sWE
qNszWmU15daLVl2WzYVak2FKJDg4tTus9fl2zFtxsExgvF68L+WWmWeuVCinOSiwI7cPBgTrPyiQ
QknoxS6Qz9nbBqPMsqhfzRTg84ML6CHyWfvn2xW2H3jY+o1KQn407O6lFwm4AMy1KxUwF9zxJB+r
OuFwHz5D+j+PYqKLFs9xNDsUz6JBiChN/HyOT0QBqVS23v5he7rOZvctP+7HXdEmd37Dw2Jt8hYt
1qZyHXwrF1FkKWZ5/QIEKa3hjCPpsLLg/3/gaOXu+CSd9G1igwtfmMEHDv1dlL0r5CFA3ZJws8mz
aUyucU6+2GP6aJg+6z3SUbKycp22f+3HkrHlGOCwR++6bBoPofuzCJDujL8TItfl7gNF+5b+I7fr
dIMGUPNgjF6v8zEYR0kZ90Wi3GU3LbpZIivKcc0xSIdE3ieOAbsFTK3TaGFBbH36XSrGi2MKbYiD
nt3wfbpXXXsKzeZypdQuJGuOunQ3cFDq5JmWaSRh+dfdUv67SkQ9XCiN5lAjb7FxU1LmnuGjOVsb
7X3xn4HjJ3NWt8ubjh9q1reTsBzOnhMXOyGVHEKfBQac+8OrhWZEcdvA6X8qPJ4icLaQ9cmT3VgE
ptRArE5ahp9jT776Qo+GkhWkc3vK2pK9MRV9Ez2wP+tHAanNQccr8H9jA367eD9UFI+gWYVkDDo6
+o/80ofTXoEH9M7nyn1U25RVmN6xIOuV1aZDXsTdZbCNTgS3z7g3iK+g8IoQxDZfHJ5Feyl7awen
wdFY1VY3Lz9/qV4pMxv4FiIdwPs4Kowh09EFQKK8Towt6FDfhMzxTIDDBZi31fEUKK5fpzZ1ksPc
LpM0sb1Jvzo5VynWeN+l+WyWUuc91KFj+5obUnCtoFtSaZHmihyC6SwLJBkRnFWDc/95BBnArFSr
bn44tUP0JR1npepRxiXx4K9nd5KnlFW+Suj75lUWNdkp1cVJacTUE19QaEoPKO7czIxY7j3RX/ge
TagSq6of3/IaLN/1kFmoY1ZGS7zqB3rl9Lll+gHsGHUZb84RpsPC18qOH8TDmBV6DWuYv5dE9z/o
SYECWSXHx/S7hgr84xwLa++/tfK1JU2OxEg59ja1UjWbIqLmEh91LrRxjUyJG9E/fntse7OfNUBv
3xkT1lmL5oprdooO5vBew+FZUHuDHo9q55l04kyOTpkIjEmBOzE5x3rkLK9sqFA3a/oCNfdqi1Wn
Z4YwnxExKxbP1sj3l/+GnJ4MnAgwhL4pM4C5VWQf8tvl12YfKMiZ5zwjyOkJGvQEa/1hfyk7Gs0+
d0gc2wqHOnkHQepjf2FdlKjDYcxF8wnIMYDvTZTYxIyqhcCSGaZBkZg4Z+A2kWKBoBPFYsIWqhsJ
9o2aHjM+s3m+e9IjmksnH3Pm9QrP6S3IBkkhGsg0b6HxbRvsBM+RTK9OLr1zC/NQxTtVoqU65MRp
J10fAKqboIRIhP7r4ysS4dn6XMA09DAAstbFG8qUu6xXPeHSLDWFRd4jCktwUl94EU/5prwIJfeq
eS/loT/78KS2frAStMQc/lXiPr/DFVIvqKhe/SP4tLNfU/sJBRHTQ4JEAkuPa3lvg8tfeA4n/pDw
85HSximMcnqROzMVG1YnRpenBKvSvzSJonBMIccraERyDpCnBM1YNZQkabJ4aWXZ8U3e6pYnYDtj
ALUTASwHeZ2cM01dHGfGW35aniWMJGX/7N2HhhTsrbKr7fiyx1ItZFxcUZSvZD0PIH5j5llgNaEg
FJSDyoTjaXFK2nywHtvTYEeMa4VzdPhJ2qm5nlNtu4EwzZ19ZK2veeiSediazJucwhgrSkJA7GdD
2CnvG5VuZB2AdaD9+n9B6SvWG92Lp+R7yL2XDurmCW1Ql9H0bO68+6nzDcE6CPEPbfer6ZY5uZtI
hxKgk9SL+sVch9YcX19o2DpTKnSG84AguPTQ82BmmrVG7Uiy3i3F7/TmOm/nqhUccHikQHnAov58
lPXFMDYr+aXuHSYL03JP1ufgsTpq9ZIahXqCtQgERMWyQmoqBJ4AhI3FfuxWlo1YkCbDMHNvYFws
jd32isjroJWuPxi3T5VJIZKcxFpdQlGhXmUj9nbp6LfQWalORVMO95t7whf3D2PRCfpU3AiOlpam
VWtfYHe7fR18Scp+EkLL1s2enEHI92QIk5lcGfv//qi+0pJmf7x2+8TZxouHrAO7mqJiUcEpahJk
FGjVjRYaJo/2NKQnouWQz2hmAE6XeptIznhQYabvMy2Zgi1bsl6fLwWQX0YpJM2ctVqk6pX/Thes
Morl/kM4Ch8i9xLFsdxOzAQk+w1g2oYpB7NkBb9XncuTdEUUYx/YIXFe13HzZ7L95RLZGOtsHhBB
5A4S+O8lCwefKCiPW8ETF2LsuIWpai6nayUZdW2sPjEVqwRGImFyzkDCprbhaT0MU3z6IM+h0I0h
Nc2FQnZRF9tHgl2pqYTHnxGiVniGmYAL6MFyG5TfgvQYXE8OtUGYOk9ydtjlB1hlkZdnRLeh7hiT
MNg5CRWwyP8NWRxtLGx5fHfPaedbNE2CJAtXwoQHemMljSFFE6wIWfx3fXF8O5URDHaP4JBxIMlW
LtVxe1VSfH4FDIfnIrO3NAbF/jW7L/2XCnZtyaUu1voeNucERAa5JPrLRbX7r4/jCHT/Qkd9b2k5
3qnLu3rfzTJ+elsDVvYnEp9jIXRYclhbqPmuYnr5v/zeVlCtsZwfl5SL9Wf6d5gmPc2anl8eMth1
m65CZRRZu/umZ3X0iFTXjux1r/fVSeo2k0BOIb5Y9o/f0tx0soBG/7OwFkL/N5jmHucaPzAbDQLA
W/iUXAKLbvW8RKWKxPRLSfSnA++hRrHv/4LGqckhZ2Twt4/y5G4o6uX4pxqjhPEdgjl4uegfOzWA
2WKj8UpbVkCdhawS4ZBT7gfAsQACiR6oMtvB1XguxCK3JPpupAm9rOeNYo5QQX0u9t1PGBz31CxR
y3h5GV9HeiD3HZ9Vx+hl2qO4XuQHY4hCSMf0ebp8DDORpy2/+O5ZeDRifTcNDtkJar+Uj6pXowRY
pJjX1wDLShZ7VoURF6cI66a4KsUVBUrky++jniwhLQeOWgMtR5/N+QX9zwTIo7b2IpXdV+V18WdH
elj46iEQvlYxMFByO7yE1uwqaDpXRd5B2LnL0kJu4xsi4cEIwSTbCe3XO/FfP33zvLhCaeHlZhQs
7UVXohR1WQmraB0C1tgHzUQVUuXRo9Wq+URkD1+iKXcPzJMBQIs9xqMw+MRQWvmk6mJHM3rrvjGj
QbmFkgj0A8t2si+XVXpNEYGbAcaIrVWdDBdttJTC9dzvYMNyaqDOVofV+9ONEXaqmGAzL94Y/Irc
OkNaobVQtk0ticGxDmEWaJDU+bnL0o6cRprYlHRE4Wivh9NG6/8/to8GDMpUwgZJKRdS0mBa/mrA
C1mcrs4f9H+eAMXlg3xNv9gsS4s95OO+Bg3wugSBnUjgDWq0erwOnBuQJPf4gVUZuN4hM0+k1+3u
iWOAEJ09b/K+SbgShjEBiScTCj4AXzdK1ePOS9gBoZ0rCEzoF+w8IIVI/UGqCSFiX14bdkhpO+6D
SohsW7GSbfAeEaHXlwugJYvTjPOTr6zkJIYavusGqsCPJ0VH1PeUhzfHlCkKoCvJ18TViQ6D5ekD
A/86a99OIolepnW6KlFnPoqmYy+m0B5X+Z0+mqhnbVPza/KMggHMPlVW3lnuebLx59oMpSwvCBgf
zM8jNMuMmOTQcuZGbf3dGLWeuLT19VpB3zxO/4dSQR3UJR81A981u9OhLc3x/MBXKIx0/V4FWxjB
0PGjB9Ku5h/q/Y5wxs9C42u3PTwWaGDe/jDTfx0O/efWklZ6Qwe1Q/y8YUd10p1BrGYGMlJs35WF
8KVJRwXEW8kEpxzWlpIYJ4y2GaEbivjZDH77BEa1nI+oYMj/zbMB0fD2hqQTiSBhYkz1W22rzQVQ
nKPM+ciKDhVvzwL5Q8rZS+0uMQVZ92rlfRJ1YnrQiwFaNucITrbtB+qaExgQvpsqC8YJapbYSS/P
le03GHW9Bib5AjtTFUrdYJ6+TfQHB9YOxvljcG9rqTEgBZGjG3Dtf91QJEp5R3nUKAYJF8qYzUgA
44Gcjgtm2EUh+dp6RGrdK7CFEc1CplITu+CYn1huKK4PHjhApneiyW9ROxd6AtT+ZgahY6kzdG/s
paWsmlXJerOIsErwG+kaVpgPJMVxeMvNo8JaiAKk8KG1xSg4Wk0huPjj1mKON9TuADOMHbGqjOa9
zAZzt307z3W76BeOoS6sWmI6qo/67HJFumxybmmu+lBnDQ+72G9F+a5b4yrhwVxpRJIoY2k23ozU
mJ/v+lKA0OSmc+JwzB0iK53rUQjEsWnfV2S5UHF4sQ04qoD1fTe5FVjeHZJGN0NI/w5ufPMXsvK2
wZtiCeSanp4b9JI3jKOLGuXDyH1RhlXcmaAjHqLMgJdB7JUGY876CoysM/ILFlabS489aXoE/1RA
mi4kijCRKoWj3MJbPY3LgkiEmvq9Qn4jtlEQdYTDlFIttRO+5OyAdbYg6sbXQUNeX9R5dovju3iI
Ng5itYJqiVlKIsgSwHVIQigp2vEm2xDDIpryu1utz2SA4SspmvQT+9zAXHzQofy17TPtVTDiFXPy
BR3XBl9Ta3xL6C5LUORSM/X0Ey2vybkOfwLzuB4+J/WLcsHYLRD0xTBFn7tRN6bS0JyPpV7bYRfs
zTqxCROhMlxhgX9RamIgIivbxeD3TkoX3u2qjOvHEe9/ZrSHQY7fTnRngDRMhzSvBwJIJemyJKEr
BIqyhvkF8PLsL0XPYiUWz5BhW2yHNvZ/PkFG1ZhkA+7A6muuOvA1zvOj9E5lzgtKWmjpH4VfyzCY
xRwWb+JS4lch0dq3+xwjgKdDGpR/Wl7muuWAHm5fFM2l3ZOtNwZfu28QIxQ5HUJGmLTz3kqRKftW
9uPK4pI8scL9rI78uYpIT8cbuwogZsZ7daQgMJQqacFRnJvhKzgrawfus8uY1zVNcL46RtXp0HA0
OuINm1eDlOQg63RQcEqCXL14GJpu+cZpdZHGpU9Nem9aXJVtHObKjemDcCOnNh8FFDnGsdH9eBlQ
OsXrI9ZIBV0OV2SRAle9WrNckZ2QNvpLlwEA/WH1kLB5njUVp/I9+GNufOfdppw5HGfTnHg9kNFS
Bu0lsuQwDRbZUWn1QNW1Vi07w/udwVvz0AzbCKcA5im1UmAwZfxUxJhVb5r0x+IXLLHdHEaeNxF+
fPjsHauelV73oc2/RlCZPoJGXb1/RrZsCOOpHbQdr4YdkF0nwJSqcl/E+S0IB4kceWDpTlYs0bxV
dVLzCX/GmxL9FXcKPktwXbIxPzewAEVkheqfBqzPLQf4j5Xre9RbG1a2upR4HG/eDeHu64wkXP8A
UA/DVskwUQ6jikyNZjs1HVIk8M9uOiYHhquyiQBbHJhYYuO9OREzBA9sS89rxHflvvGsUUdbkdUJ
qJuZcZ6Oov9XJQkWf2RH+FYfVmNm+YfvdopMzKth1Y4yvUbjV5s5ftEt6qWmi2YONoRqjxtTfx+K
/0PCYZTvQFYx3T/UVcXzF+yTN7Ee/m6RG66At8Z6hm4PYtAGJ4m5YXUw0W5O0gOfKpIgekXKuG7e
aMSX0qxGGZNWCruKKaYav1kWlUR4asVzNOQ7KypCdGBEs2XOFuNyRmicQpJdPHnybUPjikU7PsPX
N0xhSU0Ws+QnWdecjZP46NNtUl21VDk3Y0UR7CQK/yYnfKmy19jOI0gtPgGZRNYa9HdzryEgHd1U
Srxx5wDlnBsBHEXOVMjTK64/wWp+2L+idedK1DI3ybW+/e5FjsbNkXT7HB1Oi7RJPMEAPkAoFZww
UN6Pzz72RUUiEYUxmSKsCY+5BsyOaheypO7Rhya1ISewFVfNYb9XjkpykbKbatNq5htMKyWeuj2N
25J4IE3qOXvTnic6nfjuqfhASxyYs60k7EshPeTS1H5zpTVn4Kl+pzkI6/o4+FdBmsEOyLG+Oqni
oeFyizEUT898sSDYaIcPLo5MxJlZKUrLb3a/noN9yknlcGosO2tSXGHGu+TeH/2xqRavI/Rrkoeo
ZEY9t60uh5H3NJbX9VUKCM237e4/GXGkJGlN9r8SCDiORUmpznIIoVZCUzgypAPdZ35lWC8ntLkh
9UbXGUn2CkmwVkh5DanQTME+f6eRYtf9FEAZnAh+c3TZvKcWVYEoKxU0GaofOI0v6lcrW+OBEFcY
R5rYMpvUliBUxDw+QmM9A3uMGUhvK1SpsWpDcCPiBrHXibyIgKVlrIsOs+UJfiNoLw+9wAzSvnp2
MaVHSq2+uhx15Bi2DZz1SphU1QGmj/+3y+dK3MGYPcYClewsjcYcluoPPNtdqJuCiEggZMGt2V0X
BkuTT8WNpU+Epp2V0rLP/mBVOa4GwWQKPQV3vWQdvaO7A5wuYWWx0Fc5PL2u2LptgW/mW3xAXiG7
5WM4vXH/kngrg3uZDJNASojRTpjSBSWFjgQPrZlzPCY51Cc1yN5MS8dB0+xKW4d6D5r8N7mrAwPJ
X+XtLciaxB0sPDMvNOXu023Nf0ros23ORkyWcbYQsmS7TwIMBl2cXsmygwG3Op+X60l4wMKsyNHo
OkNOsHryTqdu482wZQNlVAJediGdf3itS/Cl59F+uYv1O4XuTlgtKqNo5zKB+e/ZDSa33CzfNBY5
9Mxsn1flBZ3zomjGtVKifoIkEMoDbzgBMtjM+ctVXGCUCsNaWKuIZwWXJncCTdvriv88yp87+dN3
qwmEn6b523W/U2CwD0Oo6byjDW95dnm/cnmwIYkAtSltQpbJhh2qUCfZ7ntWZ8FOGLuhFU/HqORz
75M0zmvZzoep79mKvI/aNiOCc06nK9xDwTsSlp/jmTjASdaAUaGGlQgpx3leBHSOfmD1Et4eQ++x
cuY+EjCUTl4FS0U/PmvS6e8eyx+PrZcuNcGSyMvnNSIIuv+rrWH2GzpudJIKrbIUNSDSTjWStGde
RlQ53cKghZdw5kkzYovBzDGSUHpyE7Wmr8yn4Zv6BRYN+iw+tjPUIUTVvVIrVimXuunRhJDQBVVq
h+nkoaiZIFMFBf7jlvyD4gndVtcmO5wslAbefSPEPejpIJ7k5zRPyLhq8vNOP1E+lCOa0sak5vAZ
TNiSjyggL6TBJZ7paxngH8Z5xZLqmw5k7KUrqcpa0yZ7R0QCqb2LxUtYoxT8yr+pHrgvpr4IQzH9
iEs8yR/GOKiAiVm4vFS22WmHdhOKGNFUePNAJ1RPadmg6aMiW1sUjUd4WZgut8FrEyIBLNjvEYmJ
q1+ppTfZ5GLnToggiPKSTw3kSWm5h4k0jLhZcNZNZVUC8+3U4bX/0GWd9G1b9r2mHB5KmBZHbYPv
4gCKf8aWcQfpUt4HdfgnkL/RrFyXwaZCH3QbkgdM+1mGnS1fpC6x+kWwzOk1YUN3FwEaW2WjZ5nj
pWm93u8IPfsJ6eAmpD7ovL0W9mGF5uoD5z3Nndw1MWn63QREVi90oabdCaG7H+PhCgIR5se5cZNZ
8jpZB8hY/oLa0RGok3CxVIYLvf3R0Vv/ZLd5dIolMl1iOZO7xQvzbTFm2QdqyJOVUE/WsKX7RqD+
j43Ia+dpIaP3tMgGRrehEwfAmmfRuBWxICGT3ypXnfc1gLdaLcfuZ7JQ8UzmFeV3RkT9fcrPsPl1
hDMwMfF8bGTyweDaMFckMnZkvRXcXBAejyVBOTiPN7HzeWTYj6Wqb608nHS/bTqCw8+aSlBi5umu
/MgoLDFLcK9hZMMhT2WMrUaV6BKiJm3ndDQDz8p3Y+Q0WhhU+9mcxtb9vDKYOZ4S27P29Rzr1s18
pbdHY6DjzvtSp4Jn8iTGTrBEawRBllUqvaYAC+QEblwieFShZEMzM6k6rrak/9LQqD0UlNt11iKY
7xZRHWi0VtG5TiZScHcgYkr+qfokbazeHWfSXzbCLD3WJhRtid2tfwJ+DaogJdUwFrxM9oTwIUDI
0xyB5qbGdjpraHr4ZZx1btjQZJ+ddeLoenpR0Fx3O2tXK3H7VzjJh+2U8jFdCSxjIbTYheHEQp9T
GH/s8N02KNWfEhLWduU2oi94sRgSTiqkAfV0jbKhpXVZNbjCN0ZEa42bdDpKwGkBMXEcgedE0oaT
NjT5sF8291hYXEJKrT7fuaRn3SCeg5gmBLPfcivpPttBAety+4s8vMStoP4yjmacarKeaszrt9Cj
94wWc312VRqjqDFUi2Q3l8YamDclOK2tbk+K2PgVx9PM/4rjaDdOvEJV6pbiUQoRGH89g4mnYa50
bR6C1J5WzS68WFgrcSJW7IJnLRcWX98j+A5pcHy5A4YPDB6x5/SEtG4XlM0fAdZV+OcFMWCuplX3
S0T48ycQ/3JJ2p85zbvXbpzgmyc8xKftMaeooEuXjGCeyNzrJTv21lyfGgXxDd12HqXjXmleu9D4
ufmvHQPz4W/dkluvS4fig6G54v8oNuJWVsw5QUIF9gNliBMP01I/cr535YI7yQIbl9hAIPVJdD6J
fpXznhfEGvmpfo4E644J1ob+9DH/IiFnrBT0+dinKIDuIwEvPM/fuCKaRz1C60uzMQAUPOMGp2dJ
cccDMU//45F5RMnzVvOANVpxfyRZwu1hbaee7EC0mB7gioNR2i/JOAOj6R3uUzAP+gpg/vCYvoWY
sogKswUI1viRK/lnqYseY2fRsanE9K0GFYFcG7JDtXnkIAnYYxhu49IKmvH1XUtOgzF6dzZsdSfp
/ySf38+y1tEggYxgo+5Mvl/Vfi5jC2d9g8AxcL1il8swTC1qE7tZcxHDq9a2CLqhdKfMsarUbUiY
J5g78uVQkra8lVKpdteC9XiVqly/bn/EAk1vTXStIadMTjJ5pHxZbROhyfvF8sYTEWeYtSc24paf
Smnf0O3yt0CVffxrt7TQBgUdtOT7jm3gqBVQjT5xySOLuML5785a9dZzin6kIo9i6ZlAX6faLbTh
s2DhIqsLWGIPivnz1PQqULhAH/X+demx9OKFVMVQXm2AeVwXTO7sPsh/1IceK/LXq0s18OGLl9eH
pSUCuVL9j6S6XxhmhABeCiyY/7lmdNUtMeavatXGvtH9rkffT8jC5uWhdcUpt3H2YQATIr6cDrdv
YTOuFD4if3Tmfp70waIVZ0OTfkn/y9fxp5nnEwvplOGBgaGxidcrlcQrGYYkA9rh4QYDcmbUgZP8
i1vK1gGkrDtg77j9jkVzTifWjPdG0f9kKgC9JXagTqyWb/m2HZNbfAcJikA4isPXTz9KrE1aci0Y
lLElnYY4dWyWu3VA08YZ0tebsQKw2583nkEnWXFYnUOg330r4rCsjFUJn9/Q1bxFI/SMNuA5bUZF
GXXHwC+NJvcO/1neiyOpOQhzn0JTy3JmirUjGmjrryu4SZw9L3JqsOMSv7k3zKtYgLVVMOOQVjz4
F3CWusyb7sQrC+9gFNdlNEgeZY4r5FtSOBIVwfBc0QuV8fci73ipLLCNNazSW88PzojtORbR8y89
KaUOsWW1gfm7fvaAbdtxmt82z8vYGp/g5/VDGktWUJ66BNoZoPX1lVpdjXm6EYZE8NzeGDnOGLor
JHA5dg97095omXO0BIaJnJOrnDrDBJAxicS0W6pDSxV76mbj2UreUDDkAw392C5K0DysTEU5nXxr
LZPxhhgfIkvaiY4JJu3aXri6n2WMBnvp6blPmQD1HexMstaYxx94xz+ARgSU8BrD39wSHLbiYggD
e7fapDRP1N8EDKpuqroeq1JmrtKdHpfbyIo+6/9dp0OmqCUcVK4g4/MdIjT1kV3UbiKhBTVGZh9G
Y6/6FoWy2w+GTyExLhTcNohJrkLYrcpovKAtrxDiRjZ1TvIjZnm1JLIvViR1UHPfJ4QwTVoJAMRW
XJUDfc7UOMOyKopvvQcUXJQMQvF9x2STsqBZjLJOHzqWYz+z9A52DzoA4D1lybTfhFKtB8DE+axs
NwkU1aJ8UM7K4fZYnUa+5cDK9rThGynhd78afRcs0PAubAjT8aP4/8uBjACAsLNUAvgWhM8zO7fS
EHN+gRq6UCQEmrZ+L1UxOqGbgq+59/TcyVHWfNZV6Jl6ge/tkPAZIg4OFeMDUKMkQix43Q2kTOuf
FaoHzfZZS4g0tXiyN9/Cp5bb+Ar/T6foH1GDBfn+g+Dn+WqaGB268V3rvuoVSSCv0CF3y+093paH
tLon9GXowoCzydZ23+W7MTHLaf2xPm7QnszJsy0EhVR7fHcrXymYCOB48w2wC/19T13EI4OjvCeC
+Ya8FdPMBwN+EeXTJxW7BXvL6OT/WBeILKsEP/6Uv/Z22ww4Ol7M8oQUrNnoeBbHt6D8CpKc7NpU
cImbnTBvy/+LWojPqGEC3lEebUr87Yb+beNO3Sr+Ao69Vhivuf2LlHbLgm+P7fc9k13p3Ye9om2b
+AKG0f6sfxuqLDpY9DcaYtwMUiKu5CV8duW94whNWKlS0MwH1PP9Dw7b1eUQrptzRNyca0PRK7Wf
wI8voVdiFyaTEdbMDEZr6gassmailvKbxaUuk8C8LsP+1XeqPoUIwPkB/9jxMpf6+c29EKZAxMS3
Nc+YLvBZAabH05UzN5cpRMXVVWfT2QYvnUOUhRppIVxlrHd82O19kOstkrQ3k59YjmrVHnryfNnb
1yuAgfCaB/faPtk/E1JCxic4jqS1KzVoXAVzVuc+CoRKmFGdlZHtfNc6LVv5S50cMtInF+KQfeHe
QmMF12/g928jWdwIlkgji5uvs9iiLjEVJCDuyQydsysWLJJ/ZOx/7j1YkyeaB3SGqaHrw7B4+TFK
70wmwNwn4R2IYWa+f0doR1VpjKDUtDhwuTxPFjuNHquFCuK4l6udxmczSWkEJtlmW/a7EKOMGsBy
ydkGkMcWaroF6eBf/ogqgz8VIlL4T+G/Fywqq9Z4wdd5xqDm+J5w2Sfn9LVuR2jM1i6T3krGYQ0W
1bvOIAtrUjPFw+UseUhXDumBtG1IpjTDnQGnL5MOyQfeXU/K73pygQyMm+al5GZH67yp5xjX//u2
4dJJqxyoRxe4sdrfcFua4Zk0rqxeAvnFmmwsligXQHnfXGD99OLhQKWggf0iDeWvWBlWP3Jb7WiK
bdjD2Fg40NGHmRavjz0cEnDQi1StzUaRb7RgL6pxNBLAEpiwEdojo6sjjqEDT3ZbJA2X0V+cq01s
hppw98I2z5UgAgFJqgnF5RmCYVZJni1ZWvW+tXwX4WmuxCxJ66oxbqYH7X992KuWWKcjfw439C+v
Pjmj0Ko+AUUQTRpo4DOehKF9tv60Q7JCuy3upyCVCYhC3ywyJWlTJltzOv+Q1XHWHXsyOZc7jEX1
Ea76ylAo2JruyxKv3yAsK9yAya8ubfA5xvbM0VP7dtoBnwu0iH0p1WklReYk81yEsFWdoAeTxcxm
SPpvQTOhwynI5Sw8Rbumcm/3uhG85UjoOHTRfq+oDXdpIueimhJ3h4I98lSBwmQIlCbeBD6VmGps
Hx0SpM/AGGQFNVVEBdB1A4Ce81cPc0GnVRIGBHPkSPQ+6lTLjlf4ef1ZIxLPZGc6l6LkvaUkGlcN
9Akfw7pYCXs9zlqRW5PJh7yXJ7NTSWVE0IyQdFPIM7nYXuBoe5sFpbjXUQ0Ivos2vIN1tCx7Ye67
69xdzsU4axXckRAGRplkdgODZVtpHob2zgYLqdnM5AJWhVsBHR40iTscxXU79FChCLf9TaXSrAyv
1O4NhpFu6wYpNXQ+QCYpfFCCFOywgIASljj/CCp5rh+Ml7936IW2WQxnVwre+rHxHxZtiKN9G7vt
cFuSa44rLTJ+xlOezsXu9n6S2czHCsRDRCXjVCw++uJ2gSIQBNjwnrAMMQUxxjgrn/KalV1c8Io9
6onfqZmVw/BUge9wRePclYar205X7dBXLrmk6fvazbVphPAjdbw+D6fmAlTpCe2FAaCYabdIKZN9
MJItUWeFvOrXRdKtoW+tyYK98yjBM1zuN22T5ygn5ZMAYFvPc1OJLryHryWHj/p9tahIFyE4tial
3NnQ/sF6aiAF3VVJDEOBLVmR+UFea0CnTBX06UCneEEzg0/fNCKE6SdGPd9MEs0UNONj5vsJSlot
fogd9H2M+WJPKiWx3E+td1PXc5QGCBQE997zMpWyJ0ARVe6zkzHNgIn13+atf3fMqlXhMCpO8RFA
yLpxQ5iu5NAGwmL2d76vLXv+U5+mtAfIJuYm+V28lE82Kv92+XgB6T0OJLT/kGk4pp0/6SsBtB29
N55eFA+HFXG2T6e3ixCTzDWy0qNmA6BfM1rD7XNnWDwhyhS6X5nNVp/oC+osowWxnAJs43Hg/4ZA
f6XYVTBTQZbM/kr8irMJLkajZc2Wk3Hyo8/lm1LtP912QL4Eug3Im6ZQDJlWjn4iBcZISmyGZjos
7lIW3EpssUv24oViv26VpO/75mdnPQ/fE/lUmiQZd6NB34SD52Bs/bj4T78XbrSu9w5895aJywcm
kmlTALNy+6qAJrqXZQbAB25MeBEVyP3TIjKXQWGsugyqbJ3YrB1eS5WGYVdyeZwpo0iV0WP9Dyux
fvMB8knJbM76FAzWOxD2KVZqDkOCn9Qj0mwYv2bJrrRTqWDF2XXO+6jFlTL85KLu4qhVK5qIIw9s
DNjfvvwKGDIiF1AmY9RTKNDvNu5rKfa3TUqXHZfxd+wVrJwuBd6vJFz/zga/Dij1zmgjYPt6UleR
QsG3fQqSRMN1gr0cdpqMcl6D8dN/TgSncycGAqXRt7ls7UL49OHmvz4B/p2oQle0grQyDXbzfZcG
SJso3C8KyC+XV2RMpSXslzDqxxYlf/Mnq5J910UEDLS7yMv95OSBIozoOW8JymJ4TUtdx5YQ8PIh
5gWPl5m8R6jLmGO40R576J3OkqGiitoZb9Vo85cJuIq/x5H2xJyLPfyz6G0zmCDiwDMsrP7jyGP1
L/d2l0p1JrZkMSlo3BCJf/XKBmLkrBIsUC4AfyhKIxBImLVBy9Hm8quTFpJZmDcSTLQr3I3hQwKm
uqz6vkMcBrC8uUCCjwimmOv9i8GGhD6jXZhzhq/2zQkHUPffe9bXLxuNsmhlkjphQzKObfKKOC/J
HACglmDiEaKra0AjS+h6oFFJ/vuVn6zyXQhg0oHDHLRbb51mKYdqVpCvANxAh1ONckuzTayxE9J0
t+coof2UEvz6sTtkxqfMSGsDH72BoUninUzW2RFhBZIsw4FmkkaiWWUhnYC2k0o8cXfQ4JGHSZER
Ww1/aNOx/KENpj0fcKbjs+f/O5oZDUIMgcBg7xpKKXuGrjVaFQx9StDC0jxxgiZj82d1D/vQus5O
WVsK1115rSmZi0+qF13eZGfZ1XArO0p7uItd0fecz7nctorUut+nNIj7DxCZEf0TWptFrNvcSZkG
4vJ8XrrbM2Cc8XPWzgS4FuAX9ekTkUpsL0jeLQHFf6wL9W5m4KpBmpsAYpFtkQ3vbdo8zUI1KCvo
fd4j8wbO/DcElF06I8RZfYxQI/AFoUImvRXAhndwAPa5eCFvYQ4XoafpSqL96V6o9Uuifiw2Cjba
vGm+NIGFjt7BckQTw/gjeqBjxGMM2KkH/bndRiTXT8GCKgqHkHCNARNie112+Ub+Kv8IuHpV3gzW
uW0X8XR7wq6VINe5DiNnMZHREsrZDwkcuCSO3KIfD/0SA3AkTkxAkd7H+Gr8fqygEshvYx9po0z1
3E//RhNelTgtXWhCpOBwKYOWKwsN9xzXWkYfYESoTnwj1+pbQm1P28bkE/e4oaZzW8lot6WuTPbQ
54gGKUr87FwAwq9BgVkuRhUCERJyuf1a1XGWBQZI3tCnn6e1ZIiSOv/5WPoYKNkmZcli9vW9nLJ7
MsCriUpB7guGQhvXDCM0th3zoxyfo/4nlCm8WcXPsuibuaQIO8iWpl6RNxWASJCS5s8ZAgHKI5DL
/YurrPGm7k3BvdQc/8AIS+XkBXw3otTCfoK7AEcD8BhQU4k3lm5oioBV7G9P7kxe3uy4N/tTbg3k
SlYKDS5z7ZNvK+yk5L2tUAS+5lJ47w4/QAgZ24DvhiPSZqAVS2RPs70LNasuy/SA04N9PvYq5DKo
9fo9EKv1fOCSPvHjKUwB7KGFfwwhsePV7zgg2sY/yqsFXbtm9ZLxQroUR5EP0/h7JLwFJChyV3gA
hHITZ3zJtxlinvaSuVIzHnXUzwEKkifWNIVLxW5Htzz7BJoqGe8uG/4EJ7/vtOj6c0UcIXHC6pK/
KogAS2V/XGJTn4QFsTmZYGJvGDmtYnQtOAGVP9Q5aKIgDIav6lhOYEhOY2aLM9N2QAGauExtf2/f
JCEqHa/mgMxzKiqZJCa+Y5sc095unFeWMdj5lFBC0C3620cXMGAqUeRBVh4LfcubhJzrqGk6mJyj
8qljMH7i2txjOsIYLNR8a4YQOoF26PTyjLcLrkAg+sVqYZva2cbUkuJrMXvKqwM06M3gCCsIrnAI
gX/hpo07IVwuuQc3ieoLSKI/rT9ixXyJt2TINeyy5u8QbCfqD05mE9810EsViyl3HLnL3o/D3ZjW
3qLfagcgDgf7waofRgiEPSLHhEp3LelQquriqeD85/QEX3s20pVUJ1fBkQ72kZJZDMGwKFdCu8PD
JvdBdAf9opmVeUslF+ipdGyCzsQqzXz/fMTk4VEEXuZ4pyYabf3jyjcxK6/4YatMTFT7x8dF952h
ZMItEHxAj1FjvHGHz2e5chEH47LYOB7XpHdY9gYPHKNgqoXNP5PKAzcG3eRP+r+dgqsS4uMOa7qc
+DY2zevRyRQgQQGrz+/WRKrudGe2gPIWw3uS7/gOD0V/DUU8elPGFV+P6UAfMEe6fAMddGlFE175
SV8qR0KcFfDo3laRg/uBW1O6ff5RQf8x1PkBmZ0M4uqv2P+H+q4ThttV3JoYwwvltTbVlRVwirXC
krvCzX1cxF89bsen81QmVBNV0sHAQAl9YruEl6LyYP4nPv2IWfmiozlzN3GWb53H5zxcMLm/TiGe
SC/iluUTOYT5FvBFEn8u09/zswYGzSo/aDMtHH8bYoigzUDHn0G705lGeO4OwRtFKryduXb5+t6F
2iaUx7oRJbOYfXJDqbAHacvHwv5t+ScDMBhIdQOCYPHKb9R6JpLh509q3NOatd+ksQL4NrVra8HG
y5mVz48sV5wwJJeWsMQsPqseeIVICj12JmVEWd1+UqKHzSremSpRFyM5aqq1OMZN9giuQTyR8f2P
zqZL3Gwg2EbdFrkygS9npo2oUzA+2XsR7aydUxFvPX6ILJhhPmS34Dfcuziu3fpoRwx7vbsuD3/5
/xdfhTtcAUOndLMM/560VYWLyXfhq+GcrKvF/c8EgSBqJRhKiNhmL4uzz5/X87eTRZZck9UAEdBs
yZJdu716Qke9+o6ZdpolvsB+s9OkKk54RO6l/6RdY4dFz04vPVyxtqOl2iUbAGFnsUk1AjG3SLz0
/IzV1OQAT+qyqWw69Lp1KEjciGw+2Cbe7kyKO3WakchlWIWWVLX+Qf2g0R3zvSHT7KqptsoCvINy
95nHN+yPD7VD/Dcpt8br4PBdmd1MSur6vHxkmANQH4bqvR5odIMvulPnayXYYlOFW3we8sbSrmZo
fJ/Awg1rzXHLQF/gP9TOteD9+0LWfoKo4CeqxBehA6NvA0UIs1w+h5WSs6Sus/Q6Jngk0q12RfSI
fkV13pN3P6xigK1QlRVbHfesIGaN2/WNhAFS7MK8zUGYQUG/3PND1GrFjVQUgXoR3r7ZHqmqNnsU
+/bN96EcKMandGx7XT7LjEnFw0D1psR6Wx+sfCzP2y8sK639c5Kg4VBYW0j7o0EsYJ8PEgrQd/PB
/NvivRaeCZrwRvvYkclRInBgAJrJDMs92xA3xAMv6L9QljgcNu+4ouXuCONiul333xIAtr980Tvj
KQ0Z2eBU8RdI5wh30MiqFpBfJG5b+SBPq+cvBv5LyJ7DAXNtGiG8IRRR4Wr8Mi12aIRCcuVgkzIs
48L6NEQ7FILjnORaII5CIhAUXmFSdF957sVJxkOCEj2d0K7wuco/Mt+XZXTBbcvW4GVDLfiqN7Ua
7JQSOC7nOof0LM7fB73NJeCYccWO0tLaGfWnJwRPzr/hxMK9EzOJE/azy9yA+7IliXz1n2sLDhQf
BKl83ngMzMuu9WEfVk23SUmHhKteLG7hlswFG8h64lARsLj4+8ad2VXdqIOkV3iJjmIMXsiG0mHj
j8HGCJnkQtOuufr7t/CZv/vlFIvUgBDfJDpXflK5Z9nf6me53nKYSqAx5JP2eeciXQQmBuzT64w/
0aObtDHTTeeEWWU1dvRaN0Y7ep5BusSE2tu64p1CPj25wkuwF1tMSyV+YoZeKiHk35JgLdgqZJCH
F7gRYEppx2c45aLeRGGVcwuhljnUatt/D/6jFCvVFFdeGl1VeurnwwgiuA0Ir+xJPYJ6X0Rf3++d
ig9nN0f3WfCUUUgf4/6W/Y4Bmkmkq7Wck6gHTOrmxGioFEhmVJnos0grzGGP6b2BUosbFvk0/05k
V5WM3NMRGQWFi+KqYlWmHjqklDWQhSmTIz/Ugo+27YYDWDV4JIRtHyeX/Dq0cJaaVIy3ftoVCbyT
v+CWo41YapUagnS4T/mlKVrbiEFSE530LL7fYZL2QreAaSONcs3shtFxa6HgQa+FGb7C0f9fEYPD
34RwnQKWtWRtYcbgvD0Rbz4qQNb5W4LS8EkNt6EEaJuoSElfSJFr+feo+kKtxcZwRp8d/MUXrfBv
PeDn0sqDHqfdGa/UDMCKR2zUUHw2Zrl6ONSAZqeuvq7tl/92dW5+FtJEQY1hTD1jrW+16xhKkUVj
xP0RZVcm/rlmESAbKw5B3YIMp16qvE5B/gavlkImKoBihkma8YK6pID4r6q9foqLqsHWFMskz9IS
c+LZVQx6sGs/esJziZPaY1VJpVIewo0XF4Y291UCAlum1vWKnq7vwLXv9hjpYVB1A3vsKQaiff+6
DAvFU69T940fxKksHB0TlJk9e2ZBb0GaJCTzSfcANd2r1qwMU+dMqG9oNJkPiNYZjFFAoJkIGcTH
aYZjyzBqqy5njkxGrBxKU6+jqBGI6bH2+iR+WsIkCexBD1x/Xdji9PycSZLeWfLBlSi/bpH/HwSN
D11krEW7577Li8g9Dd18omkYqVQHlCjWXP5JfLg+NH4t1HN98kDMhrkTjUwlhWR516VYkDXDcq+s
G33iP3eh+YFd7eqRKLtPb7irOktxJlXGDAu4QHUrX8xXjF4RCLPtAgJvVDn8Z2s=
`protect end_protected
