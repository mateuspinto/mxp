XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��%��T�A�9��H+$Hll+6c�U؀��A�T�1�_[;W���	5����?����t�Jc��3IH���˦}�z�8r�Œ��E��\_`|�g5x�i�xD��{�F6jz ��� o�5h^%��L��MM��-d�u��
w��ߜ,�^C%���JbH�B0���U������T��&Wr��1�������k1Rb����l̝�|�� Y�Wp
�j�����܃q*>%`�\�6xdĈ�Z�"�~����Goxn�cd�T��`�����c_*#�D��X�n:�mv�4
~&+2 �J�b�%�A��J��8�_�)�ZwT�z�s;"��Ik�o�=�-�D�<ښ�%���搳s(���x�,��w\��:nW���v�)�i.������?��T^�� �����^�������ٞW8�{����^L�`��R���h�oϙ��?�{M���'��7Y��^����@��� !ĺ�I����5YA�ϟ7l6)���>>.��bē[�'L�>2���A'��.�]�\�ഗ����j#�m��W*z�P�ʿ��W�	�P�Vv\C�3��:;C��-�G���`�&�XvX��+��`z �۝bf"q�(���cǰfL�V7�=���Dٞ�>��ٹ�-�!#)2����w6(9�~|�b�#^O�TGB����
�;�ZPx�R�ʃr����.ZKGlB�S�M�t>���۔��EȐA�nD��UEo�aP�|��2К(��=��v�I�æX���$FXlxVHYEB     400     190)�5p
�Z����0��F)��ѓ��R�_� �ԓ��]v�$ƪy=�]70�9��Ou³$7Ѕ�5�vkk:{g����4����ϸ`yu��jFM9#�r��ؼ��ao{0�%��sB;�i��+��ā��rv�y^�wx�N�2�XX���$ޔ�^w]竤j6ck]cВ���*Ĝ����,�[�j��n��C�+�=�a��9�x(+�Ƿ��������dQ�b�)�ǽO�=�]I���C��H՚ĥ��1
PBnw� )�_*���(����=r������*̒�OE4�e4���}��2�	X�R�~A�#!�%��I�G�s�<��o�O`y|n���Et_Z���e�W�[I�P+W0��Gy���iK{i��g�W�h4��?��FXlxVHYEB     400     1807�d��ZM�Z� ±,�(*\�>�ڍ�-���I���-�5�&FvS�2������
O���>���Spnj�_M�=���Yym��2|c�����g�'�o�/�P�?��-�"�m�=�L��ˮ�a�6@\��g\J���v� 1��,�DM���|��[�}V��m[Y]�8'-�R�cI't��J!������P@\������?�VUG�P��9êC�-;}5��iT#�
�&����"�M66��*yE��ofȕ|���-6�ߕE���#Z�Qz��JTn�e�H�V,���A<W�gv���m�j:*aG�0D���+ k��ѿ�A_bU���C�?#O{m�� ~�q	&��&������S�+ΑbЩ��l�D%��4�p6�XlxVHYEB     400      b0B�>�������x������8���Ԣ��7S]�kK���S�*�o������	@��E�8d-N�/PY��E2M
�&_J�� _��rq��Z��ƛv/�:�Aټ��K[K�?c��򄜎��su8���Ui.֬�S_����[��z� !�k/�5��lM��ۥ�t��<EY{XlxVHYEB     400     170��a?(�J��}/N`�'�zyA\u^�+�n¥\�~M��d��ha���#b/�",I����2�.K<�~�U�;��ř(�?�c+�b逛�������8���M�_J��+%�>3���}��U�`�/��4�c�ͼИ�]ć/��'�:Q�gM�Ȯ�U�4�MTe�{��_� _&�z��c�5�4J8��4��"� �����C0����Fq���G��������[p=�
�U}��M�7�j�P�#9j��x�v�䦍���x�yJ������Iz-r8'h�յ�7h�����2:X�% 4-XQёJ8�{�k�:t������.���75`O5\�/�!��uj��XlxVHYEB     400      90�����=�?#�iƩ��ӢS��"�XY9�c;#I�&�TB��
��6񖶈�Ntj8���^z��ذcK���k�9�ZrD�oA�W�F
�=���T{�K!yrL�#���X̭�!KM�B�d�[f��w��W�,8��1��*�XlxVHYEB     400      90
��P���Κ��_��'��[��(B��g�Rlhw\�(ָ7ԞS_C%��ĆxR��d�`��o�_y� ���.a6��Zc�"�ö�7
�׏o��}��J���&�8����XLc"��@���4l"���M>B�umqOj�YXlxVHYEB     400      90��"�.q
S�>��bP��-�F�N�?ĹRǋȰ�+�UC)W<P��?�`�L����8�9N��A�+�$Lv�1Ͻ��b6�@�n��Xmw� ����`F�q0d�Uv���J*����d<A�q�q,�i�=�O��<��4XlxVHYEB     11d      50�f��NZ|}�w�r"��o6��_b��0k����?h~6q�Aۇ�aq�(q���߉��d@��`3B�Vv
{��8�0