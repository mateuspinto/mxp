XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��M�ת	�=�>��,"c�E���{�-[���N(Y��v0r�jÂ�*t�|�ǹ-n͟�/:t�k� ��G��%�0|}��d��>����몡7hO-%�}��`4#�8�!f�ԃ�1ȋU�(㙆+�����2v�x��ZͥÏF��6bE����?�uϽ���h���B���v�f+x���G\m*��u�@TP�InU�������+�k{;rt�ɣ�U�C1;��
��HDU:��S
���q+���mp�~��!��e�7�"�������KJtb��+K;q�,P���H�d��ǼE5���}Ƿ�ޱ���񲛀����V�ٛ�Ǡ�3B���*�ܴ�k�F��7f.RԲOb�LtW�U�d9/�M����{� zRow'���}��Kn��� c���S�f3�����U���"��)��E��N?*�Jw��Jy|�D	`��Up,Q�ds���;�h}�5:$�����P͋=��޹%A�߸̞���04�S��1�'�8���3H�)�|��ob�����"��sl��th�K�-��v�s�L)��Ͷ�ML�JKQ���>�}
�j]�s��s�%Q�-�@z���w$>B�D?�bq����/�Nv���D�%q{'+_���.j��j�k]�e���G�.�*S�R�9ƚ�W����� ���K'�t5�ܹ��>l����G�t"C�9�oX��/&y���W��q$�ը������]*#�_�|�59%�iRA���h�_��s�P��OsM�$E�1qXlxVHYEB     400     1e0<���r��2n׺�4���9�i饼1��jڼ����~�A!��,��(�5Յ�Z��	���ˢ�}�h�1��Nd�𞦒�/��U�xZ2N�F�{`�@�`�F�.��
_��4�|���{� ��3���쯣H4�1AQ-v3�
����"�o1������jHo� � R8���S�����FKY۱-co��25�����V�?��a�#���t�-~Nݯ������b[\�}	5��V�C3{�:��y_L�SS"�n-�4��J�c}Ux�Z��T'��O!N(��F�!��1,���3�99��F��H4�H�ht��n��f��A۩-���
K�۝{k#�iH:O,��ȁEY���`	l��]aK���dc*D�"/��m|�B$�e��HUB�E�������30h�w؟���"o���!*U���=8����X��D �'в���{�-nZ{{bֈ]�����y���}XlxVHYEB     400     1f0$:MT�f���PG��1����b$�3���Q� MY��Y5��!]�Ai2����@�}�'��3b����ol�Z6r�JZۇ��� �jii�=�������c'�k���@ٹ���F�`ۿ[*ⶊ?��Ӈ�Ŷ�\�R�`|��6S��H�SqɆ���q�]�0 �~��A�ر[7zJ��Em�P�r̈́c��Ix��n�\o6V�Q�Xfev �}E��6f�2�$�Iks�܅���ȗ��;X�r���9�Z���
���.�P��dp����	�T6���Qn0�(_����P���j�C�-�W̗���đ�i��vc��xj��N��G��,�Y�OD�:�fƫy�ϐ��6��A(��.[�D�!y��rF���֭G�>���M1���U~yҴȓ��Sf�[3�ڝ�ø�:�U�Y����1U����9�!���"�?�:�ő��9��붗��b~�	����3������U�(�
�{�h�gXlxVHYEB     400     1c0h�Rm�0��&��]U�}Kq�"i�j�!���O�r7���}�K�DMR���5�F5"�DIw_�ޠ��r�*���Ϩ�%c"�[�C�Z�ř|�2o}	�vʉ�˳�ළS4=�U~�.�*�e�_�))vrZ85�i&��<g���g�������UL�������B�N�u�f���H��;���i=�T*�����Z�	/c�e�쉂�Z�|��V�$Rb��3>���B5��o������8*C1-ˁ�C�`�{���d�Ѧ��H�݉���GlV��S_	�:;^2�݊5-�b6���Hn��:��|��I����H�i��Y��Jj��ă���\1g�����D��%G����'<|��pv	��s��g�|� ~�jK�M���pz�DA�Ӿ�6��u��)?3)!R_?����33�@h�N��߹�lj��̴����
)[�XlxVHYEB     400     1d0����2+S�2"��j��]]�r>4zW_HW��.,�M��ԗj�uR�jK`RC��"z�D�B�̫v_„� ��h�r�&�$u��;l���o�/�Do|a�雕�3���*���YPީl�0� ��k�	=�����zw���Y��P�K�D�t���^H�^��v��ćh�M�Z �k����OM��Ċ�)�Y��[� �l,nn��eU�7�r���X�&8E�3O�X�*Og��Ƒ��<��0n�����X��m�n�!ZX�:Q�t�)7�V���Wi:�����o��	�����z!�ue9�����ۇ�3�h�w����:��w�R)�ϭ]�p��hS�%sϏ�E�/�� ՘'p�K��4eJĩ�׭4n!p��(_�.nF"ki����Em�f�%Ru��S	��M� ��&�4�����4E�"���	G9^�i�|����C��yC2]t"XlxVHYEB     400     200���l�>�����0qI�G���V.�&�C�&��텙&����W;���Þ�g�OU�2r�߯[�A��,y͔j{�;�p�H:"�Y�0v�Z�_�����琲���LFф��-��V���W�P\���P�B�ӗ\V ��ۆ����Y�>-�D�ӒQ�+��>�^���oNE��ՃLS�+k��
�(���+��=�v^�kj'UC������
����y��+����@R��X:� �B�'�jlXv^.y.�GU8�#"�ܧ������4 �d��+�w��� 
���2�,j:دp��R��Z%�bw�/N'J"�`���.����g���;��Umf��Bԑ8�������\o�Z�;���
��U�Μ��nޒd#�����=U�*d
�[�I���S0;�`c�`��x��&�z�Lζ���tF�*�2�.5D�X�n�ubY�,�E�i��5F��X&0����1g�6e�l!k~ڏgXlxVHYEB     400     150��|Qr��P5����?���<�~���~P�耨�u5���@Ӈ��� 2��eo��qU��+ax!8l�g��G-��Π��ȃ�,B�"�.���M�D14��E�i�y�l�'��vΝ�����2+�/[rf؇��i�h���3���pAMi�?f.��y�ST�����ʿ�k#���72�l���F��2���IUGR��Y�v�1j��ć!TE������}4En�yJ�e��v��`
_�ZI�F�G2̉w�3�ŭ�k}�F���h\MOF�i����`GqF4��we����z���S���ŏ��\�J�ޚq$�V��"5\_R�XlxVHYEB     400     170J��׎�#��~�U2���Q�OC4j��꽵V4<�X"����Nq�)칛m� �1KT3s�����4�ٙ��{ˆ����z�������")�+�K� 
*��Ə�E��~G����VΜ���q>��y���^'��W�E�b�L�4Ŀx�?ꦧC��:�^dΥJ����pC���1Ŵ�V^����m�w����~����HheSjv�@?iÚ���=�Y>�Y)j�Ϊ�s[��1�rXO%�L�p2�L1���-�d��w�:t@`�@V��\x�/K�4#�X�hT��-H�E�c���en�gM@t�A`-���fϞBPM_�ɐ�tY5W�=㿽�2;-�W��E�L`JP�#�b{�XlxVHYEB     400     1d0��6�;J��9����py�=��$_r(�����	}�i�b�����!t!nCU�+�~A���F������0�V�o��V���n}�K`tɠ{�+5����9�I�b�KM.�oLخb6��ts7	�֬.=�
��9�,���H��=��_��P-��n�+� �Pf.2�����+�v�;w Nu�W�܆��h�d/2�K� �����'��:F�YMD����3��k���
�4"�K�cB����`��ޥ{��(aRZ#�p�E��CXr�!]3b���x;���4|q��ko�h5G(�O���7�P�?���^�J�bK�e@��IB��A!v�W��%uq(*4�G1�&�Q�,"�B��0Vtmk��V�(�:�@.nn��y3ɄO!�q<��4��uu?rϫ6;r	~)0'�Fra�2�&�?�����#�KQ�[F�s.{w���,`]XlxVHYEB     400     190�;�+6�/�})K�H�@�<=���	�ęjn/0ovׇ�I����մr�.�(�~���S�����@���N;,��Ҥa�C�0�d����qrQ�m�4�̮3�Ե�pKHtw����J��v.�o�+�u9�Nv����z,uE��H[�e+�!.�Y��@��t`���Ǜ֕�Q3�2jS��ڱ"^���E��3����6��5k���.��ǰa2rʶ�:���^8��:��1rwq�/U���pOw�P�]���z$�[��G&2�?����w��~�5m����%�{�+��ay��Lf�P}�6!2H�!�f�_UDj���[nc)�z��DsP�X�NvV޸��u9�D)rt����0�O����*?7⥊H�������f�/'�XlxVHYEB     400     190��p8t��	�6m��0a�I��Hwt٦���*��ݒ�;=�:�4x��R+5��",�+T#��p�ؙ*��P���8�	?�������G~D��s�FٛT�#��`E/s�Z�BL�[�앞�
�: E�9я����]���ދ��*ʖpwZ=*4b�Ĺttl7�\.(����t㍄9����v��z�lS6�rSk����EJ�ŵ����*.��#ݲP)����Kd��hj�E�R+=^�t[)tBџ$���A��ʮ�u
�-_��� ���X�km'�	�uV_ ���H���E7��X�K�j$�?-V`]A�u�Zy����V������dED">5�����\�Xh|6��$?qe��e�ÍL�������-��Y�XlxVHYEB     400     150���P�^�o���Px'B#�_������06]����y��δ�@����Q�wnN��0R�;`k�n<54����T��S-^��ݶ��S�˓1���<��OǓ����=�6�حV�7�p��l�������5�U	u�|�n鷝�D���A4;��j�#/�r��j��
�3�V�P�ʹ�r/����3��q�q�(�_V<J��d��%����?���H��/���GR yQ����ȧua(!㝘%	4�����-d�Έы67���E�_������?>�6��g���ZD��uLyK#����U�ڒ��IV���r����}���������XlxVHYEB     400     150-�`�Eo�{���j��e�kOQiH@NS����D��w|�s��J��
 �X�)����o�r{ݝ�s�Mm���)�	5��/� 
Z���O���GR��wh���Ce�6!�஖W���v�M�<�g�:P\eΨ���ͯ��< ����R�r��ؘ"rv���m�ƳΙ*�Nr�馳��ZH5���=f1�������葤<-D5]���E�_�}�O�o������}�^��92��K�B�=��=��ʅ�*v(z�Y�g*�t�@� {ݪz�_p0�sq����	�d^8�@wBD�\>�e
�2�Y���l�m���hXlxVHYEB     400     1c0�"Cj�E@����3�4|�M�|��9,g�*�x���Ccܝ1��g�(����ې7�d�?v�Eu\%\9���o�Ig�)�^�j����ߊ?x*�^�^� W͉b$d��b�'��>B8� 5��8���ޒv�!�1��}���_nM�����nP�Ф�?�~�6k��N��#��iR�u��$�R��ڋRޫ#+�s��߸�9\�$d~�&�@]&\��-t�3��/"<��{o��-+9�y�g�h�����dpv��������bwk$2�U&�s��0�U7�� FAUQ��N�����N����Z��v�DS��bC�y/�\C�v�i8������i�$A��@���h*��Vᔁt�GS;�k ��0��^�����=��p��e�Fvv���s�
����\�?����4S��*�ԯ�������T�02qXlxVHYEB     400     1c0��5�6W�a0����?9.]������`pG��sR	�K¥�_�`��+�Njx�r����o�s�M�2)��D-N�vV�����|,k"6zu����CO����^�=�=q7`5�����,�{P��qq��'>���#����݈�����*�83���
���ŧ�5TM>�� 5�Ң�Ɉ[�t:�+@	Jv�"Yŭ��&�}i���F}�g�A9n�6�Z|��`����b�ϲ�<#a�ݔ	�;B�(���0�ۏ/z�w;� ߳��[�����E��?tG�?h���L�jA<�R.?�a*���aǛD�7��I��gŢ����Z�����/"�0tJ�^�YQ�ye-w�����
<��X�t=� ��vӫӱ�9g����r��E҉���WM�1C�ɚ�/��K�ȭI��' <��:>�ڿ�I�O��XlxVHYEB     400     170<)��=��jNaj�vG�z��K��5��*G0En���9
���8 ñ�����Z��ձ���t��yH� �L\G�("q�
�5�
���e#���*�]#0>iA��M~�����)L�c�[*���)B�}��_�3�,۪���	�®�At�W1-!²�����Nn{`����!׹�ԿxCԎ�|�dt�ŋ���ú�����2�*�fo�W��
nq̌\l:sD�I�J\E�ɪ�\��c���/�t=� E6�ю2nra'ir�xp��ͪ��T@�0�6m*����/I&��+��z�͏e@�c?�NT5�@e|5"�����w��{̍A}���
>��u�9%䒶��W���1oZ���XlxVHYEB     400     200��fk}?Զ�pH,f���u���l�Ɨ��PO�ZN�!l�O'�r*Փ�ݒ�T ��.x.q�����&񗑤����:����<s��c�H.x�G�xbȃ��Fe�,��f�:�5���%aU�v���٧�w�����E�C��W�>�x�C|d��氢,��yQx� sӷ�JR�"sW<%� ���Jr�"��x5�=0"��F�U�cPk��'1���7hо�UCJ�t|��x�_ �A����y%��'ǩS���eK�n�֖�0�F�8��~��#ȇ�c\~q���Z]h�-_V.��S(������i�N͞��A�B4��^�� �qYb|�s�zD�4�rU�K7�Sӌ��Y]�5d�����Q(��E��!���P�Š^����y�fb?r�m	u��>^�A:�)Y�zF0g�q)�I���H�R8�%w�G�B�l�l��Մ~ቩ7#����[y߱~���j���!	��Ug�����>.��k��#�PA�`����!�,XlxVHYEB     400     210k��S��1�LEO1qCV�t�חxf�6�qXL�D�����:�[a��T8�C�����P�gu��H�'E�A��Ljg^�$L/�|'6GUjrl�ʋa���V�gӞS��z����������I����Q �_��P�Ú���^�'�ܸ.�ho��~/��<��rͬ]$�ƈ+���������\����c��w��!*?sN�<�=����xC��j�y��L�g�6�kU��d�z��`����j��X;3�ǅ�1|G^+�U?�O���ELҤ<�M���0+�@e�5����.�Bm��!��*��"f$p~d~6��%�nZ�2b��jp;��Mx�S_���@䟕�0�������k��87奚�e�k0���_�$l]"�(�MWp���,5�� �f�p����--鴺R������{��x�*B��O��
ydoᰥ,!/Z&��^hn+��j8/v�75��5;�t�m�}�]����Rm -�rN�����;�׻�XlxVHYEB     400     1c0��
���s+��a2"V��>w���|��m�=�����/�'��B��?ly�?�vf�f9�=���pǡ��m!�=s
M�AJ��*K�5��r�F︬B �_��9�$���>���jO�ƪ������С��L������?�)��w�>��L�P��jbJ�8j���,ۅ�粔���,�$��z2�^�f�.�cИht���p����+��z�1�y�;�4��ml�%�lD9뽊�T;�� X�l5�N~�����-O㮷f]���O��.��ǔ:�ʴ�JW�c�i�%����_��x
C?U�v��������Y���+qw�6s�.?�pՠ�ˆ޿gj�cD�De�%�!<:�r����/o��D����hej-�y�EyU�:�{���C��!���I����K6:�B67�1����ploɃ�G��9X��ȈMne��{ֈ�[�wDB4XlxVHYEB     400     160����BCFm�#Ak�\͔�@q���Y�v=5���] �?�R_灙��L�|�(}����B�q�j����{8Yj6�2�p��OP���7��������f&�Wq�&Ё'��/��Rs̝��=�M]t�X��I�l�}�&*�5���lzUh�Sxu�@��h��@��F�H��]���w9T�^FRvr��!+2�M7����� ���v��]��زH)�2���J�l�XD��	P6�Z�u7蟬�a����o�����p���z<A��*���!�}�d`�;CM^s�#eXx�Vs�9 �揯�[/�L����0�φ��\)�R��Yex��>O�mXlxVHYEB     400     120��V����RW<Dy�R���я����3[Y{���N
DA-��I>X�~�%�<p:��+a��1� �F�����݈jGer�ș�:��,9p!T��ղ-ט���c�|����=yhlU����*k��}S� g�ko�pc֓�q�!��0�ҽ.��M�O�a�0�2"Ұ-�%a��WF9/�9ɮX�n�$S���EԊ�z~����)c+M����(��Pn��@�dfu-0ݕ�J�U�/�]=\LZxo����of�A�E��W�5���J���~r
XlxVHYEB     400     1605�ZF�v/"��6�9���F�}�u�$�X'��	&5��L����ly
����*	�fO/Ho�I�A��@��W����jrj�>j�X�n���S�A�3Ѡ�G㖵���H֌vR��pR)@�d�`>�B�oDK��;����̲��t�N���O�5��	h���;������r��~ME�sm�7��y�czɐ�i}	O�&��!/̐P��p��!�U�,2��ph�0nT�^-�	�'�ζ�ᬖ����q!L	Ҟ�ܰ�%#��[5�mH�;��R��(W��Rb؊D�U\|,6}n�R��A}�#^ˉUn(�+��+cf���z�F��=l��x�O�,aXlxVHYEB     400     160݁i����,W�T=;���������9����c�vX̩�����	�d0�\>�Qvk';&~�W���(�?�W����6P�!\���Au��Ĭc=�D(i����%��{H(��ma ��������V_AIaE��h�(�{�2r�*�>�%�'k)�"������U9զ�8�|{G���^��$�*�L�ȶ  ~�Z[?�s��%��fO��d9d=m�~��$W8k��&����Pmz�qE9c�"h��H�؉%1��JVlM�Q���]�v���/�V[��?�^�pQ%��6n?�|��>S��M=G�U�j՜(	�������i����XlxVHYEB     400     200�����D���z�$�������Ey=��/����Uw��ZV�+��<�͒M��<CՖ�҉}���pH�]�}��-\y��u��"��i�h��^��7i/Ͻc�י���^n�0A>�����S���3���H��������!�aR�������	��i��R�u�'&��qL�1q7܀�m����>�
!$p�Ew&��������s�^iӲ��$��/�P�]:�ƫ��4�i3},(�86��!"�ڞD�J��;bkǔÁ����-�o㣕
6y�����s���4�{�5�?/�Ҹ��u�#w���T��#�}�s�Դ�{4n�=�D:����ZH�UV6���L��$ioQ�H]^�)J�O#)���T!�\��}�ޭ��g���l�vSSeeEE��v͐������7�W�5|Z��W�]���l
Qc��-k	y�g��Nc�o��i��82م�}�����<�|��0B����xQ'<�-�J���Q��D�-L2c�qXlxVHYEB     400     1d0��$.����2�D�̌�.�鞣�lr�No�xs�~Ի'cs������;��}�/���a�+fn�
޶[���՗����d�Z��fח�KL?Us�UTb�2zm�<'"x�7�n�a�+^��dlPD<�e#�U;Й�T���l;�p�ST��
�m�LQR�maY�2�������_�[��?Z��2��l�y�͜�L�jO&@H���J���aJ	�P�K*\ؽ�r�]�W���>ػ��i!�z�<\�Ş�[�5p+E�;F`H2�~��@�y�L�����
r�I19�4p��K��n�Z�8dr_�_d)�A��U�T|$9�U�Nc�EH�7*=�!v��S��敫��F�#$�A�4̐�8�e�_�����
bͣ��UZ{@�6I�>vG@h�v�� �=�ۈ��Y��e���Mb��T1؄��HF���c�\�p�.;������N��H�� ~
���XlxVHYEB     400     1c0",�	j���{)��s�گ'�(Q�v6�laU�$Jmy'�q������{�y���x}54��[��1�b�
��E������\�e�YbN�i�n���H��g���mʤOn���hL�~����]\q��`��w��P �S�?�Lo�=s��0�e$������^z���}��+�Y�:�����h��E6
�.�FxУ����`�i��H��e���2@�z�3��(P��#�=/��*�k��0]��mvឪ-�*���E#̶y�z�戮Gk�I��u0�I6��9��S�?��*�_=�խ\bd~�*��*��z��zAְÏGX��js0\��k�X��PEJ$5��ˈ���%�ک��!7������q�����.�u,��_��8�#����o*A��r&�ZP�s4�~H^��f ��L;�XlxVHYEB      42      50�抶Ҋ�X�[��>@�!�*�?z�c�FBG5����<n�8'�D[k�{�v��ca֡�����q�f�s���+��