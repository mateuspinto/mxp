XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����#]������3|���<oq��	���.�\�k<i��ڦ��P���"�!�z��9��q�����O��u�i��ָ�����!���r*^��ب%O�w>�gq���e��7��˕[\��V��~����p�^t���`F=ۜ	$@`��'Ey$���9��W$#a�v���{k��U��ǨeSf��a�uC3�i�S���D*�&X"���3�4��h�^�d�ej�n��e�&����}���ß#?^�̥�K}�%���q�����"wx�g��o��Ւuq�Y^�u8s͠����^�/4�
`.�9/�uE�uHhbb|�W�q��
V�je�,a�w6�d�Tͼ�q��������n�锺p����Au�*��3�{�xD͐o����� @!xVB@�ߘ$F���YB]vKsD�"�4FV�'^ګ��݂���
�u�O|_%KI?��>x�6%�6���?�ڶ4bO��$�]���"C�^�rtU�nJ���6�w���i��I~��J+r�||?�}l�%,�'O�'p����Vr��!j,
6Ϋ>��6ń� t�-�6Ɋ� ~T���z~C�W���f#�|T�(��8Ӹ��<l%<�XȚ�܏�9�:���(���㘓&��M#��;�mk��ҡ�B��}���:Rt�Z߻��w�}�c�4/������uT����Ս���
1�c}����h��FCQ ��ܼŧ��=XnOy��b��Ev�F���^��Z�a�<�Q�Z�v� k�>�XlxVHYEB     400     1b0�>}��:E��)��ho;,�	�L(*7_X��d���$dZ���2�>� /������c�����'�����"���qCw?���Â)��VM���g�D�,����_�����|2��4�x܅�i�p�s9ƦV$���T����K��3�9Ǘ͏�����3|뽍�^�kz�꾔:9��7����.��������f�-H�uL�j.\�o7 �BZ����+�m�Q]o��Z��q��Ape>x�
i��lu�v�k�R�����[���1�$n�J��Gy��soΡ�����gP(�r�Xu�J���s}tR����oRz#x�Gu`�uv.ގ��qc5�ޗ���y���hn�Yw�}k5���|�a�f�4�n�Y�u����=�/�yg5yB!kd.��
��R�d˖�gXlxVHYEB     400     160 r�=㍏v�0�xW$�c�����KmJf[P��4��T�d)lR@,Gs�*���rX?+�ަ�Ѱ�2�����fSA���,{���x_J�s��P*k�k+�;O�BA��/,� �o&��X)��))<����pAc�`$:��Ω��W4M��~MT�+u�b�?{ _D�٢�h|s���5��T���u��l�wav��~�ol�e��Pժ���?�ٻ�P���~�0M"u�!���"����4�5�ӌ�W=�kg2���J9D���j�Lܣ�\͸$��0���]ΤGC܀)��S�ЪdU����i~A��g1�Lxz��F��e�6Wy�$��-�qd8�XlxVHYEB     400     110�lS�CO�?�� ԙ��M��@� �F�s����U�;>#���|@�C~oH�<j�m8�U6KcrgJ�t|O���1x�^����.�^6��0W�m�<��R9�m��>�5D�*�:�c��[�����DnS�gQU���.�䄅�7O�i��N#�Ǒ���m���[�YM}��2H<+�N1p,
F��h��6��$V= ˦b�U�����έ�6�3�J�f�`yB�e�5����M>����ӼKGDŷ+^��3�>�OXlxVHYEB      42      50*�j7C���v?����{p$�6�&��B����P8	�,\�z�K"��?>���k�a3�5f~ �+"��5vd�Iz�