��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���]X�FwC^�n*�Kkd馅]AƵ�Cw�Z��0�|Q.�;�.ڊo�Z��ixM��q�1�y�6�Ӭ4���'~�i���i�M���J�yF.b�?�]�U�s�p��s���POK���%��7>�S�����C�A�տ�׹u=6��5�J9WGh(#`�P�H�v)��K)��A0�	qJ��\�����L?x
#I���r3�3��b��-\/� (}��}|�&pʬ�0MW�
iI	҃��4Q	��Rӧ�`���F�m�?E{#�.��wP�޽ѝ�k��I'�����p�Y9�R� �x��~�3:�̻���&�"�_ۃ�
x����N>҅}�RTFr�����Qg��q��T5�Z�w�K�Zg*��Q����sq�jC.T���g0F	g����4(l��Y�24�L?-�|��Ⱥ�Uiz�ݓ���?�V ���8�Vg|o.�4cJtt6�uԼ��ž��Hi�X7��t{��c�L� 0@k��Se��t��#�I�
�B�3��	Z�~B�t��.�y��#��uA8��"|��[1���#=�kLt;��[�G �.�%�~���;��,��zhp<��T4:������\T��q��6��W���3�L9Z�x�';p֫k;�F-�#����X�~)��Q�_�T�<E7䄗����?:G�Y
��ݗIx���HR�6/­c<���>O�-�+����3g^�65�^ Dl����֙�"��Z\��W�����<�4�0
py��zw�% 1v��tV��$��5���⚑J�JЅD���"{��?&Jnk�N����f�?\�L!�02�\U��P���M�bL3��a�L���-�i�֤����O�u�v?���E��������dJ�e��y���4ȫE�ۼ{,���ͣ	%�^"T�M�������"k���T|Q���ٵ�A�H�y�l��fю/�}�Z�Bjf�{ܕ�q�U�8�dM�`i�Sr�/�:�����|1h�7O>"����:�HZF�@����>�W+�L�"��-�/�{o.�^�;7�"��-
�{=m.`i��JE!����$��/�㸁U=OUe@~-�Ѿ�1�k�O=�?�.��>���Mkͨ����ZF���C\����kg���i���]��:e��G�-�i�u/�mG���P>ų�\�Y��0c�eK �&��1�R�yZ�l{��V�G,*�/6����v��-�S�j�TlX��#m7���������/�t���:t�'���:Q�qZ_\��I�&�6�<P��R�95��Gv���yE`���{s�|��h�Q�o:����t� ԁ��S������Ԣzx|)�@�q� p~8%����:����Kn�ю{�N**�F�is���-iGɣanŰ����k������>���c��GT�����Kd�9�F���B���U�g��}����[O̘M�ׁ�1���/��=.�$��A(�n�!d'���m�/5)��g�x"Ȧ,��W���9�l�1�Q�jne��4��+&ߔ���3�,�ʉDZ�'��y�n�m�
�	���
�_�C�R���2'烱���
���K&?�Cx�?O)a��)������z�yid�" ́�~�����F�T��*�g,
<oC��(���v�W4����D,#�K����S��
I-���ܴt���$])M��e˔�X��eZ�p���:�L<�O�z�Z���(��7	���S.���kK�����w�l̡ RY@ m���..[�	��:�zw0?o�\OҤN#E;�F�� LP�lA��o[Ԙ�ݷ��X2y�����sqt{��5h��L��^�]U���y ��s��������ʘI?��Z�S�1T_hz�K;�
k�	�3��G��&1�����Hɯ��}cn:�Q������k@M%ҹ��B͔֪\�a���)�0�ǒlsMw�y�	�	g�l���l�@��m&�W`gP�6׶�A�dټ�k礣(Q+m��x���i6��N]U	�<�:��b�%[p�2�������I-�spr���у�u�0�8O�6���
�؃}�,�s'�_F�r1��mH��2Wl��e'���"�(��&I�x@/W���k���!�@� PC�{+z�));���0.����Տ���B��']�ߡ�	�i��ZE��5���/m$���ޓ�K��Ma��n��#X�TT������Q#;��b?5h!�  �w�y�ه�l�����
�ߗq�e�����VA�
9,���mA�E@��ʍ��fXp��{V���g�Ǉ��f]�j����x땖��(S6vuwaDRj�K�	�	X��ߨ�R⡮F���7��1��=8?��Jz�H����p���������8o?S[ʙ9�&tn�E�H����k��7o00k����xm�#�R�#pmΠ�m����+�,� �߯ف=�x���ٰ���*��dKIk�ci��N��v��ګѲ$R��v�+�'#ȃd"{�н,��S�����FJ4(@e�$����ʰs�?��D���,V�C�9�#a�{��u�o���9)�L@`����ϵ\P����f�������)Ewj0Yz?�;��	�lʐ\t�+�1:or�	<S$*~'�ghwAu4���E�������^�J'a��D^4$FG����WG�I�?�&4�CBw��eu�Vs�\V�~dn�j@3qԭ �tI2�!��tY$��� ua"f�� q���ɳ������_H$���3GIb����E5s�Y�Ƃ66$�Oe�i�/l.!����JL?m�L���O=%��[��n(�=�0�ֳ�%~R䵀>jm�k]37
�Ti�L�>9�<R����q`B%Έ�N7�P��R]n�S�EG>��1�N��G8�%��������?j{٫�m�XH��P7��j�b�I��@�?��K</��Ēߎ%��Z�jjM?��S����W��z���$��f;ab�P�$%h��i���au["��SŤ˟\�q�pP�#vx���&�Vc]���*��\�n�ͤC�t�t�A��z�э̰x�Fb�{]O��)�s�ڀ.r����*'Yo��@�'��L���?X`0Զ؟�XpJ�T�ˌ��F�j�������� 	�����%�^��]�|���ck¤f���#ic����/�kw�dT���uX��N���S���d����#VBS� l�� ���<%2>X��d��V�kI\F�2*!5A#	�٭N-��P������2z]M̓\!}��Շ���B�'t���o�4�XΟvѡ�r�,�=�@h���W�dr����p�e�}<?Y��0����.x�k*��Q�|�l��Tg��^�Q�
&B?�,���O���I����Ǌ;p\̎��wo �G��B���1>�	�4d�!,5����PLT��]iU�~��]�!��t	��o���1^���`l`K��_���mI{���G�f@��5c9�'��e��*�u�h�V$�=�w/8�kch"����L AX����*�W�pPQ@����Ȱ�w鹯���)4mqY�>���W.�-���\s��
�U˺�_�Ȗ/�=�B�o\�a�M� *�_O����۱�5/�����.Y.���b�.�SD���!}r@��q4�O4?	�~��[�M$�Z|�~�2����aA��S��c����Ku���P7��G�r�A9p�j���"J��������.��/b%�W�E\ǖ��c�p��Å�YA�mI�8ɵ�,ET����M�c^*������0?�W&7m�����>��]����
�WT��\��7,'�ꠊܿ�����ܞ����o��Ɠ@�w����^���-��q~E~�[�z^2�Pr�*ë�y��R��~a�I�E������}�ր� �^����,���0��iXHh�fǞ#8���X:�j���Z���o��"��� ���4�]����X� ��=�Q��e�Bo(��ˍ{�����<�k��lxU���jq�᪠��"��Vq�9<4h��-�_uA�.��P��'ɲi�x���M簜Ѥl!u�4����c�����)��'�s��fQ���������|�Q�Q�DX�U푿IV�{dl�P#���T���)	�?��yj�6G�r����M���'��Lɍ��r������3K������Rv�P�.ETC���v���GH�8��3��"�6>�,'�5��Ϻ�	�Q����+���	�6�M���w�%��x�3(ޛ�J^��s[�[V%�l-`�#Q�����!ƾ+�1�	\��Z�J�u׸�vZ���8
2%�u\�K(�'
�G;�������k�RR������̛��m*ĭ��zL��_)�f(���(-��8�	5+�Q�X5���.���f�JF�By%�(3ѱ���W[�i�1���goZ圠�u�úH�YzC
�C��!�U��_Q�E:诜.�3�wVZ��ؑU������)�F���b�I�Vb�E�hu�J������.{�U���lñΏ� OM�/��]�����rT��������'���k��i9,�E��P�se�5`2k֋�,ta,��ש�8�Q@�t���*�Ā�T���Rj΂,�Sp
h�u���Z*(���?�V��b�E~��9��� ��Y}��\�_,�&�K!W�(C!�{���ߝ1Ù�J+�.u��8A������h�q�i��W?+WZ0vI��{;�,8������q�@�0d��y3�R\z;fF��l�M����vU�%��:P+Ey{P+�X�}��
f����.�- �T5��6���H�y���w�?>�_t�=p\�}�K�
>����_Ɗ
��`��ߢ�t��K��Nt�����qN�_g*?�MDq�kx_�d�B��i�(�a�������{�Fa�j��g!d�0�Zaա�6��j��M���v�� �~�^����ǻ�U��:OX�T ,���7�i�?�MM��t�&�g��/�����@p�I�i؏����3�s��bs�u-�^*��s +�h���o-���х+i�lbG�f���,t4>�W�6V�+H�2@+tL�1@/��+�A4��l��䈯S0�<�wc�d�~h��>;��(0�|'��h�z`UAΡ��6��RP����Ҙ:w��j��<Z���?�ηa�E�/>'y�ebޞZї�=5�Fc�>�� ^#��3H�>J`� �T�ݬ�+��uy�ac1�ɍi�z���pM�,���Pi��í�ʲn1�!͡Gkp���A����A���HY��\��V��� ��['�d�@/��d���~!�ZGC1�Q�ͯ��CK�G���II���$�������I���-�5�[+���R^ęd�Rd����N�s2��a�D<à3�o
4���(��Y��9��_OϏl�^DK�ZuX���ozP�U�\=܀�=	�yy��I�0'�Br���V�FI�s�ʓnl�i6�q�M5Θ&w߱�,�R���&W�lI	Q �jxe��Hh�a�^����I�s��\Ws(��I��c�N/��$�!�Y�p�M����p�p ����_I��f��`��R�sE0y^ԡ�b#3\����22�a>�
�ف~^��U�ݚ��Yogh��PL8=u��\�hw�����<�3��քO��	�Ǘ������s��J�@d㾒�?��.��W��g$)�Tʟx���s��n��%�&���q�M��{�ܽ嶒�����Tn�Z�]'s���.���S*�/�h98nTA���L)0ǀ9��޸�"^�X���<��VG���%f�~��W�q�ǅpFeAܲ��#�N��f!���P-"�΀��u1���ćЫ<��=oRlgj{ �v��\Vc�;c��g�4C�i/�&(9n{����mu�o�{s�&�l_�d ����x{�3��T �h���%-�A�J�;��H�&;g.�t�	�r4�����6�RjTX�D�D�lbkl�/vc~����p�{��È�Z�v����,*�dG�OwH��d�ǔ��$�y���!?��}�����f�9k����z�'�*����Cthh]��p�<� ��M�����m߆�b�nU���F�u㑈�Am�u�j/�R"�k�#K� ���:I��H�ַ<����ޗv�-ɆŖ�Ԧ�q�7���Ҝҩ�������մsB�z��e�A����8�!�t�K���������~�.H1��`\A���ى�96XWNv�H���@	�)cŗ*{l��'�vbm*�^f�(�j��@Y-p�h���S���q�v0+kD:�@,c^��X�5	�����2L�_"k��^%�i4^�íU����x�e�BP�"{�7�n�'*�e"��n}U$11�������D<��S�U(+���Oy� �ߪ��1�ZjE�/���냣h�O�>�iă�V�60����?Ov��DY#�L}�� �ɑ�2s(��GP��L�X��T���-���j0`-$m詵C�B�^�����DW�vd9#��b��H�QaDhl�Ab�Ё	o�ag�� #gs�>�,�,;&�u�O��ʰ���ɽpOHb���8/?2�g�y�VS%�Q����]@%9*/=��Nz�$��"\x����c����$FT*j�\��d����Zo᭠��Wý��4E �z��FTp-��gH1ꀻ>}cm`I2$I�s����;�կ�����7�PUbv��QN�a�\6�q̃\��~��@��bKo�����:>�Whk@/W��)4��(C��m�T�6�+�X�:<?����3d���é��.�����x<�Lb	��.��鄞�ob39/��3Z���K����W����kY� �$�(�1�d�ۛe���h���N&E�C%��f3��✤V��pw=�o�N\*0g��"JPҘ˶wDЀ��f���&̖n2� �U���bZ+�ƺr��~q�C,�����]�_w���5��G�/�Ҷ`�D0_�_(����\R��M(�C�Q�E���Eo�s������4�C>�&OdE���K��텚����E� �̓E9(��0�=-_�siO��㴿ߜR«E03Ԛl�=���Xg�������C|£M�=�캌[�Q"aFf����t�?�A="m� ��--��M:�Hߎ�w�W�KB�ڇ���ߚq�����H� k$�.��N�xv���i���r]v�N�ϻ��3n���N�E�������W~-�qd�c.��@��L�0�>��;G�=A[_��������͟����hG�~ �o������t"q����X�g�p���{�{��,��*�b7[�%�>
�1�-��rɛc���,LQ�<�.�=���[����ʋ���58���]7�X߂��FL#]����X-L���߳�I8�g`;��Mf���.7�K�l�չ�^�E����#[`��x��ٔ����`�D<�v�0���sZ�U��yG��j����9atE�J	IT);5[����-k�����&���$n��. Q �(��c�e=�ֹ����a��%���%ĩErʑ�^k_OPA����L7^�?G��E�$0�y����sbă�D2���J%,��>�&o��5�4���Y�L;�/ƞ��%|��ӲeU�֎�w:��?�RL!��.J�� ��F�A�8�`kt���)�pqK3!���J��  �X7�;��`��|��'�%�E�@XyZ�vB��GS���oӓ�����f����,�V�Q�#���+TL�q�6+�H��)�Z���WMzr�NOk�m�z#�+�*|,Fw퍏��3��:y��c�ln�tzn��ЈI2���$�=��1M�>��'/�EO���l-Q[E[�0�r�ǖ�sP���<�t�x�ّ�#,U��_Yş�Q:��@��j�3�>�p�"ɶy����Æ�ӱn��I=��aٳ����)P�K2�5�-+6A@��2R�emXn���b�T�k�ݲM:6�М戯˿��:��:7�UG��V+�>"�B��3+���7a�Z������?�� (u`J����r�r 4�ϭKa!�tQ��yo �e��d�OV�s���P!CQ�#�P���Ö�u]�xW65�M�Vjv��PA�vﳅ��8,)A^w��Q��e$����+��Tyǂ���*�i#�G���������,ʱltX�ڜ��3�!�d�K���n27�H�Py�m���
av6F��;�4�Y��S%��h���ҳ���ڔ! 5t�ϊH2�����S=�R4'���w���P�݆���r
�����0�Oq(vՅ�����ȳ��c�"3�$���\���[��	����$�,�=Gʍ�(8��#2��:5�-
I�'(���z�=���J�}�,�e	����R����C?Ao�A�2���aVw�lI����dj�_��ZoR�;���&&!���p1��(=�~h#��,S���q�S"yX+�f"sKZҏ�ʁgS�%��湥�8�2]N��2R.j�{�Yg?�K�y�$��c�����uy�ß�ClX�$܌��� 1}<	��𔶒���߈G���E���?�l#�y(��$+fx5́F�2�2t�Qɩ/�U���i]�,{�`�W�b)��p�i�Q�8/�k~����af�Q5K�thؔaٟ Q������~~MV��f��1grτ��U����-	�i�ɢ�{�doA���:�mE/M���)ĵD�a��A�}[�8�7.�qF���;���3[�5��=;�Փ�*�	�x���}�'��'�0���*�E���7��ci݄ap���i1n���9����'��9�S�.Cv�����T��)��0aa���ϸl�Q��6��{�1�\���⽴�؞c5�� =���;R���O3��A�����Vq9�F��ȃ=|��q����}Ŷ�"5�[Ϲ��0�����j�Y7�_��5�z�	�e��~���cݐH�l�6�ި��dдg�0~��j77����o+�J�0��uv8L��\1�x�s�H����e�����ݿ��J��@���@:�M:0�*0��gY�I|�ж%@U���4��C?�FQ�2�����-�*�K��r�	5��(o�؁���ί��c � f�	];�`cߠ^%�!����Y���7֝I�D,	�P�X�U�������ة�S��>C�ҙ�4����r�P]�0X[2-�3\: s�/�����V�6�P�U(bN����� �}(�mv��=O{��p�PI�]���b;�_����L��J3�ٛ���]�60^�ni�ŻHx����3��|\.ai��I 2�tA�`M,aJ"����XZ�����Y�f\�S5�<怱� ���Ħм�=��&|���b�9�����\�����7�/���#���-JH�gݝ��s�Z�6]��ud|�/UHC�>8�MSg�8Xm1%��� *���V[��-A%�Xw�K��vJ(e��KJ��O�5�b7�0�o&7M�M�{Z��N�W�P?��b��&sW�LF�<�M3�/v���r(�ւ&�^���tz;u��.Y��5c�u��~W�����.d'����d#�<����	��p~?�a.T6-���G�FKU�����[�����#�����-����n��n)�V4B�_~G�[z���	������C�9$\�L��g�VY�=4�?/$�]��F���L��Foڋ��E�[�b�Ae�Zq��#�`m�y���������q��<1�I�ߨAp�ρ�{Ff&�
�����o0�վ�v��`����_�M���D5��$�<�/����@Z~- �-~�_�� y}�1GgF=ã�� k��0����������3�6���1I`�&�2%J�(��uX/RyAQ��̼�o?�D} �x�K��g<z��5�2KE|��Cg���j��������qvJizXQ#U%�i�'��;x�����v�}G�\D��dP��
��k�z�F�o��>����͟/��"�a�Ykr���-������(��ZRö��������ֵF�3͒S�}m~�^:+��W�
�#T�.O	����s4(����MH���}끤}�|B��\��>�Q ��y��t�~�a:R��@�	��<n�h��PX͜��T?�m�)�R����C@��>������������)!|���m���X&m{���{��)�3n�Y�56� �_sX������b�g�䏤���a�,a%Œoh�n��6�'�mao����Oz�y��N۸�&Z�2��]�i��EM@��5���̚��r�[���+����JP5&��]���d�{�8݆}�H����܆'�|�Z��ۃ�~�L# ���C7�[t���2ƊO)y���kn�����x�qm��'����bW���-��]&H��ϼ�ƭ�9�\� ,�u�mp��@�l]1j���Fpݑ%���@�`U�9*�
۪�[�9=�-�?o�-�S2�vdx�7:DW��c�e��B� ֜A���1&���B a�5�On�KQ�bHꤸĔ�#�� ֵ4}q��R�ak����/1{��a�[�-�ݖ��I��9�RIX��$��	L����wE3Yy�웄�OҚS��OYD9�d�-���c�*�h�0�w�Q����J��U�3�G���_c�6CC��MS�� ~v\Ȫ4��)����j�a�9,�.�M|���H)c�1�`��=֎Ѓ�=���j��ϫ��9�`Ms�1�Eg\g�4��['1�{IV�
 �D�_��r[o$�����1��Ƥ�)�t5K2}T���G��tRJ�����UҾ�F��⪒�i�)N
`�_�A��Z)�F��V��n�*7�KoK�!l�g;0���C�9����9��F���s�O!�A�$�B�#���^\_����F*%�P ���t0�� le�����#��-����?7u2�1���Ju�*]�^W<��8�D2Z|E���wѡG��J����a-�3hsw�5u'N��/���RH�����oɥ��2bI���(���)�1��I3� �86T��V��%��S��?ţo܇\D2	�"����z�^��/ĤO�NX�*T���e�Z�Ou�{<&���Ļ��MI�4�<o��;���7޾�#�nǆ��2�io��}�}�������l)�U8So�R���O���Os�q��� x8[̦ȿ$�,b¸�;O�g���u<W@O4����Q������I�0��E��`���䋪V��3ٌ��d��Ei ��=j�d��o��u1'��[�b�F�)`ฉ>_�	�Y����@,���(���2=�Y��:��t�!��f��!C�C\�:Ky��W����ns���\�X��09�Ĝ:l@�����W2�-���!�g�H%�QIwW��<�r��gn����Y{�,9E�L����=�%BbR�*�1շ�����LV�g@(8�"T�}4MW���;�,:���tzK:K�=��� �a����_7���Xw�*�QKs)�πR�Gz�$��Ŋ�Zk���|aU�\�޷���"6�ÒY��8��Q�}�����CE��Sr�[B��e����V�*3���M�{!J���c������1�Yv1��A<�6�<Qo�D!��ߔ�o���"�6(�D����2�Gr�B���|�t"����|JSr���s��:���)	��Mx6�ۄ&��Oo�H��Vq��x9�#�x��&?o_N<��(��`f��WÕ���v�$Mt�F5 -�(��,@CA�L�g�.K�')8��o�T�{ ؋l	�&�R�vGo�j��n���eU8��wC���::V̒
 ���?t������>��3������Q|fԋNy/���'zz���;�B�0�.ބ� k�ձHo�@;r[0��ǫ?�H�LcV��G`������KM@x\r�5l1�\��.o�Cr�=�žDsC�;�`����\�� ����`��	�XT�2D�=�=G6�-��&l0�ge+�`�����C�SW�PT�*6���NT��
��'1�&�	�C�V��u�?�����w}H-�O^(w{T"��pn1.�F�#��A��{��6MMp��	�ĂZ��#��'�x���$_�ą!�\)Aؓb�W�S=��G"����1/�`�c�h����2��=8�QbO�5���Ç7{ ���%r���q�:�jh3��ɼ""$B��=�Hxۚ-�bO!��w�I��1!ޥ�E���S����m���i���Ci��Y�Y�Z�@"�N �ZѐhC����T����2�S�t*�,�ݯ��+�׵�n즌ܶ+�d_�v�-a���h��g!~�7zƫ����= �BWn����<ր��3�^CZ0��*��G��(JH�}p�g"������c�e��{�2=�����'@���m�wΜGx<�������5�-��r�5�����sDm�`��y-���R˰��~��&�n=�&��F�̟����U����^�R$kMv��^ 'v��LF�����Y|���#�`����a�@��	F$O6 �E� ����!���1�*�k�u��l]C�O���Y<�B���o��ä���a]���g�V�	�ۚ��6(�R>����,�][x��Iy}�f�adrb�z��W��vN���BG�]�L��?z.�͆�m��m9׆\�wUa��K`��u�M���ǃ���.�=u$��$�����7"��k@;���9O|S@$���>�7̦bk���x揜�Y���Z|�h�1(g"�go�{c���:����7V@��ۆ��;L.���|B~]v����_:��fqE+�����Ҥ�<��;(*%���=���V�D�fO�uuAgK�G-��D����a:Knl��b�A�A#U+3	{)�e�jI��0������u±Tʥ�^n� xxّz��OL��������,�w��i�.]q+�	�n���>>,v���r^�<����\��vн\l��y[{�>����M8,k%�^��.��H�"������9��?Ԋ�h0N��كI;��dx��M%/p���ҫ�v�z˛��J!�/�,��'��b���
�OJ�q.I6@�x��1F�z^ 7oXq||��JA"�����`���)�ڀR���Ѯ�Sat6��,0P1��1��?es�q�qS8K��A�`����X�V;YP�����p ��A��a2 �E�g���v���<�WaW���KBl(��8©�)
�/�B��@�fώ*����:��%���,�P��Ġm��1xצS�F������4��XgK(OaiJ�
��n�D�z��~��>�Fd��ϳAu{��(���P���d��Z@f%RnL���?KE�_`����-�U�tĊi�b��x*�0D���Q�r<֓H3�<�g4�&�qVj��*w۴O���L���9ɧp�x���q����z̓Ҳ!}�QsI�\�[}���_���/��i�<&de�iM�
ѐ��W�݊��zM�q�ƶN�>}�^�G�vʑ{�;0�D�r�B�=t�<�u���Q`uW/�����E�f���rQP�GO�Y�-	��1<K��``$�>?���o��Ⴑf`��*��oc��R0��k��֯N \E�M�Y�-�����	�Gt��g!ue�υY]��.22���x/r,��Q�&v�ć�8-�v���!2y�L�Iд�y*c�K@�?i,)I k�_�,�u��T�/�!c��`$R���,����C L.���-��N@7C+.����b����*!���::��c�h��8���Ƙ�(�ZGV�^���K��~�(�E�'�}���m��0��V��B�#}�/��n,�l8�	`)�O	��/Nf��_�kKF���<��2���a���8�%c�G�t]C���Q�/mE��e�N�a֜L�,��<|v,n{X�d�(���l�w��2S��}S�f����J�)�ҩ�r��̈́�g�����E
J�	�tʭ� hm�DÀ�3A��*B�k� CZ�Y�[vz�qʗ7��ͤ$#�P#2Ax�h8�"��
a̓RM�o@�[Z�ݑ���c�ܬ�A��˯=�ک�HI?����J=O��F�5RTu�9Qe7�SN�yИLK�&[;B�:���QǵbJ� k�r��3hn�-�L
z���@�� �z�C��)�s���^��p՘��o��0� xP��+%*C��nla^&^���#(B�<����36h�ݪ���rx@͎Ě9��_W��:����7���F�G}���e��˫���-ݖ�	Y���A��<砆�#8��(�9q���=�{pZ�o�Kh��Z�����an	LÆ��j�4Zb[�YY]�/}�2z;FtѶ1]���a��+`��x��b�PF)�*՞!�T�v��
(섳�vr�,��!6e��0φ?K��[+������/tgw\n�/Lp���[��'���7�zª� C_!\�g���?R�&�/�S��p�$DM�ɭ<\Ëi������U��3`5�)]���*?6Cf���KDi�Rn�F��?��;�*߸fe/�S8���Ɍxby���K���Kػ���!.
���y����b +�v�N�t��Ïu�1���ǟ%��<�9�)�"�eQZp�W�w��i7����=\y�˜&���q��:`��d�F��! i�=b�3����'X���P"`c|��L�:��K������z�����2�e��c�1�ܷ�sE�/�u����2>�����W2B�$jԧ����E\鲣��yY��ɨ-k���	xO̠{X6����]Fq�MZ���X��K��tļ���9�ۃY"�
�$����%w��5~�7v�AeyC45_���=ev�?�@�1�$�+����-�<TJ�f�f��%��x��S�5�v��N��(�%�`mu��b�m�"S!rꯀ���n0���Q�S��h�n̿�/u˘��QF�|�3:�[��9G�VP*]�N` ���=Hf-�U����-2��M��9u���_�D��[k�q.���j�ʯ'�٩��M�g�%�OU�O� ���S��V��3x�2ۥ� �`��Eȧg���>�	-���'�D!�f�h�E������C�T%�I��E|Q��O���4 �*<1rI���I�[՗*z]48���u���^��W�v����ƺ���ЩH�������������.�(S�(���3o۴t�2���re�<$�p$��]LeN�mÄE�ܜQ�/�4��m!W�����8�0u>��q#Q��mriC�7��s�p�g܁Õ����.Z�Hg�	�����\���q��N��Ƥ5�,��yz-�c�	��ZT�����cʒh�.a�r2�h+���H
�&2�uo)8��Xʂ�����?6o���2�o�Hգ�TT%�킁�\�~�M� O;|��2IY}��|��j>�R�k	�w�/��oK�bڕ]mʭ�r��Xr�az���g¤��:��\*A�[~UW.,o��%�s�c��"�w	��`W�Fpp�J����J��~�xidF=�ǈ5d�aC��s�Z�=�R�R�D#�'��l6���g������QY�M�!��3�t&�'s!8*�W���Ϟ�J�ة��g���j5<�ϰ��K����n1��(Ê�t�P/cʒ������$P��'��ȅ�i.B�Y�/hz+�Z��(��{D�q�]+�d7|z0)=��D*�S���i�������F���a���Q��F��R��Ȟ[2�*�ПM�7]�6���h �t7�%�'�"�w/����@۫�&�,�&{46�U8n�ы������3�E�G���~��=�t�9O_���7>Q�n�.��Ǩ��%��z�^"Ў�|�s5ό#Opa�$��Į�#(��B{�7��ڧ{=ҷ�.3+��T�|H�
�.6��?�j��ư�� ��ɝP;�kn8���䪫j��^$���x0P&L��*�wO�?�/���'FV��q���^hgL�_1[���"ٗ���$�h�%r���r��{?4�{�v	q���z7A�j=y����F1����_�����|I�Ҧȕo�2�?�	��Zh��s�b	��t����>{�M�{��&QN�j ~�zd�H���j�6�b���('''�\hM�t-U>X�ɭ	�H���r���8!Ug����1��Q���޶�۝�	5��T��'�:A
T��=	d�m���<p
-0HV5�(�+�y,��כL����G'����u,��E���F=Yܬ��(��@�2�Q���z�� 6q��)��4]h"�^���)_I�^r�Lq�#�����ó�B���o(_[G�f5Ю��VҔ{�(�)�Ls#���6�͟���6��{�'���э}i1��Y�֨�v��C�^�������&��K�aH�Gr�}[���5�������4E��}8�'��1{F\�+��`k8�#o�����f"����o�4��t:�M�2Km�U[����KT����yj�!+�B���ގ��#�s>w�?1��������Y��ѕ�)`�#(\��X��"�PD!hz��M��t&
�/���+�3�
{&&�o��yfM�� HLB	��j�������TqD��:|�)#��f���� �{Ͱ�R�W	��a{W�6%O��Q�6��ڷ��4���˩ �,����3O  	<�i8Q��jX�I��o��N�g��Z�xWfda�=�I�4���8jP�lI�5~����ǉXkє��$���I���,�F-��)Tn� ?Z�anQ���@����n�?�`wف]�PJ�]BW[_go��9��_p]-ĉ�z6^�K=POՋ�'�0e�H���*/1K��Gr3Ҩ��-��"�I���P;�Q��}X�8�����.�CU�;��k�#��[fV{}��s��]�#�B�Ϊ�f���`h��e�fE.�4�v��2�aeW�ȧ,u�,<>���W��H�sm�~ <��n�0*!�� �ϔ:2I1#pf�����t��G���XVDU�^P<�g���6R��&�K����yc���B��v�w�F�y0o�)sm�Y�
W��L�aD%�+|`�t�Ѻ���	�A�E�zx����eQ�6gx.G���*�Sړ�dqۙ�>u
�$Z��H�Z9��V��I��/�c
-�Z��ۇ ��%<ч�@��\TG<C՝.��lub�����'9#0}�����9n����_�\G��8��'���PP)���Ü�w���>DQ[�C5#��3=թ{a��d�]�k�,�`a�@c�İ0&��v~O�"֠������i��.'G�V�|Z�Eҟ�޻���=h+�#Y��O���]�W����|�r-�B®r���0#ԗ�6�")��Mt?�v�yُ�uB�%�_��3Rf��C?�c$d����U��e��7N+�LpO�0�X2GLV��M7C����-�j�X��KL!��L����j��ۿ�\���"+*��%��T���rqzt9���b15UW^�(�j�pu�8�ꂿ�H"u�o�Q�O�ŅZ�R�1�ia�+iXl�">�ٺ�)Բ�����&����k�!�� ��b-�-�D�n"~'[������k[�|�&y�Q�aSD��>H�[���9O�d�nA_٢�e�F\����.dF�T�ɾ�8-�D�OK.+��+ �����}�� ��^��h�-�y��ӻf����(�DX]���(�lX�sm�	'q72�y�}��gIRwm��=���Y����Gx!ds^q�J��@ ���HZP�ե@�ԋ���25��i�E#kn�I�Z!ܱe��c�������.�-6@jj��fW�\�KSt��yu!N5�,?��"��o����
 ���<e�(�\0��ߎ�m���צ��T��Ld4$����-3�jPm}��-��UW��k$0'e���(���(Ia�. ��k���D��l�X���&<t��%��%���a�$�s�p����֕�糣!�ݬkYy��nFW<��yӰ�/X�rw��L��)�P�B�10�EU�}��v�t�Q�Ə]VL�B�<y�~����D bv��9(n��"O��PO͢�j5A�Ťm�6��*�9ؒXm�d9��=	��#$+�oDE��<����D;��	1���	�d�&%%5���"1��oBќts��O�c��h������̝a�If�-�z�V�
v�2i��D���}�N�zz�(���z׀=Ec|s2h�W��ՉIY�5���2�;��l�����%zo^!�w�Է>a�]��O%V�7��M�_����y��?�Y0>Rr�h���A�.�Ī�eL��s�N���{��^��H��9�����ˡ��L��O�?��>6�3HoՒ	�ꝂM8m]�?���"?��	�=���U'���՚@bJ�CR��_�$rUܣ��2y�\]��o��g5��f�g��Q�A����~���,�_��ȣ�t� �-{}�,�uڬ؅�Zc�2�"I��4E=
����h� ҅�����%V\��ɺ��%hܕ�s�2��T��r"�Ӥ����lm�ڮS�KAբ�I�x�1��\h*�{>�ـk8LmQ-�I��������2�enٕ�4 ��,�X4o�P��2Q+[V{P��]�|`��Q�c*4egݐ��T�� ;i��+��NgB�r!]F���z�DH���/"ݗ��B�SK�wKo^=uT":���0��%[ҹ����"�C�a�B����qp�uWx ^ӯ��P�E�/H	i8�#�v�QL�~	M�B��_A,w���$�� a�I�X�>������=�4�����{Kn������f�TL�9"��&H\X(��)��%&�|E������(Z�E�-�K��h;�Х�=��c��Z�4��H)ҿ�7��cȵ���/\ ��l���ױ�蜩H����Ł��n�C�1��$��e��S�yz���)ߥ���`Yl>���CvDf�$�T<�`�����䆒qj43�-��!�q�t6=LaFZ���_������->Cadv�05x^VP �,Mۉ��4=����V��΁e��($�K^*2���r���Վ��v-п��-�� ��L��m�n��PM����߃�2Xn�N�h�C����������;�*�ܔ8I;��%���G�6J�L"�K��i!#���"i�n-8ˏ��X_��f���;d;ŵrS�(΋4=�Fԁ�yj$`�A(��s�zxA�6K�:%V;I���W����+��;-X�w+;Vx�H��[O$\^KzS��	}}��,�ԗt�;���T$x2Q8(�%P�:�U'��˨yЩ�E�L0�:m���>�Qv��/�! %fe�
�70�������8w��sekς9?�O�Q�~�uW�G��� ��i��C�Yu��^8R���O�QBЎ�v䨈$]��eD�g�7y����tf`I���X�b J-Zl��yS"�-����L�s-!��bʘ�I�BA>�N*��):?��J��s�p4VO�;z�6/埜m�'���~�[zJ V����߿��Y֋Ӡ�t9?��+XW�rv,v�\�%dD��U������*2��!�,ޞ~����ltް���|//�AOEO���e�YR���vbL��*�^�v����k�u�	2�����n;kEn�O0"Ř���lW��9�K��6V;��f�I2I����V����ݟ��AO��GH0���Ug#����V�O���t�l|�h[����٘䓧0���A+�{�3��jV�+N缝5#��d�2`x�@�p�,T�B$�l�]EM�'�nfXĘ��JIΎһ��� ���o�:]8���NS���
�J-��ѝ�Ӈ����ZjU�Ѱa\5\s����P�~�'� &`�2��8w�79&xe�f�L��
{N��Mb� ����j�2��J�Ї\N��edmk��u����8�sp@üRgK�i��,m2��F���:����n�ݜQ��VZ�Su;��B���(��~H7����+�D�
f��=_�3��)b�o�c쑢����V`А����Q[��.�����[u�s�֍�0Z�㋑��,�`�94���H��p�����V6>�F�v�@3�'��_�k"�?VY>fp�lr�]��H�v,@�eKjR���'O/����>ά<#��qX�A`�F�?g]�;�T�61-ȷ7�\\�C_�huP�3Br���gl#h(O3~�L�1-�E�"��l}h�?.�0�1��5�Z�J��9N�)U\R��2�EL���x �(ʶV��y��Cz�:��H��?�އ2]��QB4��O�Lo�Pt:��:�5vJd� 7H<��Ό��&��Y�M��Ń��4j_3:��]�=�f�B�xLu�f�$fI^OH?�9��MlϤk�� �v���#�Q�� '3��7&�]�qB�e��2��Z#F��r��5o�]��H�R��N�ٸ�Zw�$�r���Y6�,�y%1r�|�Xt+ú�y�9��(��o]m�~�P���hλ6x��v�QUˉ�����wI�W�I.A�|f�1��H|2)t�T����ė��]����Z�����՜���p�g^S��Z§;�n��V�k5׺���Z�
���K�4"�j��~`�ҩ`���z&+,��m_HQ��!O<�#�R@���&��HV߯��a�eʛdrw\X�ư��e����f�"jy�s�VK��팾��KL���Z�ʲ��K�7�\���0��
�<Πڪ/Mϳ8��Du���%�dwݳ_�����͔L\�E�r�ҰD������dX�_�-�����{�]+h�<fGF6�3�L�IP�o�8�kp�2n��0n�"!wʚh2���{�1I�"Q��]Y���O�(OR�/��;[������Y7���8%H�c5�!V��R�9�as��踮��� Vv���e�+�I8Ed�V������a�~AQ�dq���`z��H���CG^ҷie�a��3i��ZtG�S�[%��߻Wd�Y;p�9�
�
ճ�:J��:td\'`&u&E�8@R-2J�(l��v��1L'q��ӛ��6��?���{4�TZ>2@i�j;{�{.�,x��z�*Ԯ;N�=Nw ���~e�&��I왈�O���8&~,:mu��T�5>�'b+��pnN'X6�%Ӽv�OOX}�F��M5��kǅ�����+���YCa+�H{����rTɱl� ⩱����]J8�[�E���}s�	bM���YQ��:��L8�υ�=Bq#��l?��Ё	SǾ��;u�5��LZ� W�H�\k��[�u����P��!i�����∘	����,����8Ф�ŕ�8��[���W��>����WΒ� ����UZ\�C\��y��{'e:Z8��Q]^���L�2�����[�2~�p�3���yr�I7-ŸB�������5�1�{�����k}�8١9Ay��Ц(��Ǫ~�!C����F���|h~���(�8���/�t�O0KQ��trz6��\���WZ�$)\n�bRn�������O�t)=&��>���{��нv
Dx�A��`, e8�#m���$�Z/s��6Ǻ�rg"t��$�G��w�'�[��z��@���=+�j�@챗;!���B��t��W�	��m�\==�l�$�������]DM�I��s�mK1�~.0:cw���8�4�|HH{�6Ȩ��P�����`���$1
 SKէI$e�Yo��~�t�B�hQ����-i�E��1�o^sU3��ￒ�d�G��u�X��f�#�*=�BRn�M_X���,����{-x���&*� ���NMj���3m�N4��ϡsmbzC<d���G�;��q�&E�e�yտ3��	�����E;>ji������Ad)�@T(��-��î��x��#_%�7���+!$�792G���� �-j�v".@r圕�/��r���V�t��L�����.�T�ixo�� �����]�SO!Cv���^G��h&�����c�ө���L�l 8�o�Hp�|�sY��Q�W3҉��j[|o�ᤐ�t�q��jNW����Q/3f.4C��x�a�&�?�_��z�މg\����f�>�[�7������:�	5�w�1�S .,tAu�u�X�uF�.��)��KY� _�-�_2;��џ����B��G	b��?c/����+*�s�@Ѭ<x$AxC�kM&�չ�'�a�0�"	K� ��CX�?'��AB�'91�	�6V�Q�A��W�;���k�s�����\�Yp�/�&�_*>��|6�9b.��pe��x9��P���,������6�LR���?����|�tX���1���!9�ł�6��?�����#ɼ}�M��e���bnK!";iPX��4��)طJ��r�[Rn�� 
�xq��n�NK����]/I�y�WN=�3d�U��b�\X�6�φ"�9�q����t���%/"Xc?���r�[��^����Ĭ��7,sd�겫�b�M%Ȳ�}9�n;*�W2f4���
�U3�&�԰Q�-`u�02�
�[P'F�8����n���q�Ei:b�&;�(�@�R<0e�l$?e`�lѴ�/�#ژ^(�2m���EU[D�����*?�F�����+�J!(���U�v����I`�@tj�?v���� �Zi[8��Rr�o%`L�[�AH��'3lt��U�������l�xT�"���!���B�#F�4`�l���=��z�欐�Z���]����=�����Z�6�5�V�|-�"�a���{,�|�?��l����rL*�>I�Sb�6?�Fn��:J$����K���׫�QWK�$� ��mh�U�͚/o#6���DU���1u��5[wͳ��C�Ws/��<`�9GQ�l;֥ңdk/_�	y���p�
�$dq����3�s��Gn��2[�����Q��zЯ/�����"��#V�o-��qK�'q��%U$��b����G�Z��nu%������P���q������X*��r����������w���,;4�Ɖr��ad��D>�(���_��J���׼�@v�y������b�>�����Vr��wS����?r �-"@Ğ��-��!A߮���܇�.���8�'^gX��EʫN=� G��ux��d�ن���g�rP�9h����1�����>�#�N���)�x_�]�����{�)���ם~�ۍ�h'��Ư�垵A�M��4�΅�Y����,v�A��`g�ԃ�1L��ӅD����2�\�l�ڀ3�BZ�w�*���ѕ
��2��7 y��B��'�[R�YT10
9�Blz5�!��U�3�(q���^=���<A3i6��Q��vO�<ח����u�0{&�i�R�ly�+'2����Y��M��Ç�X%֙r�ᖔ�k���1c��Z�po�(��q�\�q�M|C.o���0C���u�t���� H�-^���# ��[�`Q�W�/���pA�ȡ��}("�a��4y�:|p���P����y�1)�\͑��y�JIєsVr��e�~�:��k9k����Nr��NY�E�0n#oGPP� p��h��p#1͊T(��qE���Mn����4�T��܀��5�oC�xs�,�(0�H��8�Y��!~zl��L���Z��~+"���,:�^+[h&5��W��GV��^8������P�l���[S�E�������R�b��޺��A�?1&#%W�c��EwP��3.$�h����n[(�68��ܞ�8C��6Ԩ�2L�a�ȟ�Id��'����g�i�f��I�w��ZV��F.+*�9���"@�7�ѽ_pj�OuQh����Aaخ'��0�TY���3�5�u���0���C!��/���5�<ى3Ƴ"�u8zY�6}�X��M�n��e����������ϣH��2z;i��<(h��#r(zQ�;g�O�����A89��9����g5��M��F���VAk�|�lU(�|������]��ғ�[�L�O��n�k�����t���64m�l&K��v�w��)�G+&�p�v��5�
���z���(�Zџ�\� f����g�����"��A��2Zq�l1o+1RF�T�4{=wDyȒI�0�.�+�f
���c��Ֆ>~���7>���+�c:ב�z8y��������$���n��ܲ�
����� =���kd��o$��
�����w }u�W�-K���h]�\�-ۘ��h������o��C}�Gy#R*�u��d�GϮJ�C�$��!a4帪�qָ��d"�1<<5�M�8��,�"����߈��D[w�q���{�N;Q����,�������