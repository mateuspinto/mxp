`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10640)
`protect data_block
dlD1umHVTHLMwy4/5i0ZhZkzyxyFRIZbiFAHkXul+FfI/+LWVTaKFzTH9qnGEi4ASAxuQY76s1Hi
308WEv6KZnxzumzHJRTjtZZp3D1DxUbefgh0sJ71d9MRZLziWc5DhdC8FGujAaqijE207lvik4b3
C3V4PACLv0AFDsAu0bB8XAdUmgRg9cJuZlZeLOx1qbhIqhhBaV0DDJUJN1t1GO6nB9BzztaiR8jv
bXpn4huPjwOFqYHXIeajX1LiU162cBrEBocJQ76cERyWmWZDG9eChGta8l0OvcchaNwYtAPNDBz3
oC5B42AWu/b5sVkR6lpBFJwA4OXD48pe7GYbVQqXW5eNi2nuOZsRhlHc+ReqMMphmV9uawu0Bno5
2j6jN0yjMr5G4Xje5jp0RWeobD5lgcvi5fqjsvOAi0ka3QvnUcjVO3j8icDcQiHxwE/WvxePwlS9
ZQYJnyfdxuuL8ltR2grP+AbG4EmBuALz259umcy3tGetQ3c9jPgLKN9KZ1bFx1ZDVbrVRiq0JhuA
Zg+mvDh6kFxk2y7ijo4JXn1phRDlkScFNLUsAcsGms2arv48wREXSG9MDntD7msnGPnyg2suRzkH
NSrpfKNiChtGd6w7cL6zgikM8r3FfIioNeQapHhu2TXjl80PZlzslicna71lW1vg/XTpvqZWn6UA
eb9dmtq9uLo4qNXYKRiu7f8uDtykvNTB6TDD558grlTZn/N/LZMPwMxxow5zYt9J5IKm+4i6dYKa
sMB+O6cJL3xZCvS2bcwHTfZSkK7KHGWUfIWTbWlaf9PsaMPDauPX93xIjB+mzs4sg9vMyZ5EHgDf
De8WScZJHm0DkpHm3vwM0AHN8S4fOGUKtPjEVN+4dtjBcUgPGQ4qrwcPQCDB0YfUb+NhbN72qCes
044NpndfbEUd0U4O/vAazHEwXJalCVZ8cZvgE78GFUILZZdQWszTX446B7n9+WB1W4NKjC5RE5ls
96g2YPy95SsbTbbXm136BIBW68D944TU3grJKb7xeuGNZH03Xsd1nXUNXg2/0mSHok/cHjdvmVIy
lBbUIRpIJYb7CsxvugaoTaPfkaXEe5O/IAWVihQptT1YWTSh6P30GJtTHMl5x/hoie2A4WptBGgA
+s8TCwbDBtzV8A+i6WrzW0k3N6vsKaOcuncmE4KHrKIjrZEuX4+/a1PLcSa4K0B7bszfJ1Jyd6U8
S6ai9nbAm/uTTjKwXH+F+dmoU9OFS/U0D3HGvuYQeTVYGyVg+WpkGqnAFWjYzgeubIh40Od/JkyN
Jouyowyem7+FdSTfIuQwWzmsvAisi05YAKKB2kHMwbWH68tlegg1HWFe8skfEmVs3eYjkF9fmQGF
hfl3Wq6aCjAZ1B7g7c0GUaA8SZK7dj5FR1fI6G4UNLMsuCG88Iku8czGvrNYfEdGrFYI8SCO4iJy
l+2hI4UKVqK0ahIkufwFviNAvPo04VB7C6PkpbWQMf5mv8U0GZyPZNQ9oxhBH8tOolPP1N5QkO7s
SIrlkdI9cidZhu1pBPstyD4d06av84D/Ew73czj3s7YyZuGtzH5cpEQVpoZkqjuXNwZaZOoXNoxB
eDl3kYRDhd2wwseb6fJ2dsTV0kUT14eY6eNKl91qj9Z9qGFos0Ti8YA3660uGv7n1aTHFHYUskvE
JXtfltZKmSF/cZ5/58Ebxjxuu52Kjq4f0ipe8tJWVdfZJvJbpXOVdoa4ePgK2ZJUOWVpdlMttytl
f9Bbx9QhNzx1bLK239YEW1yMiWw9Khp0IP/QoUR+vvyPQ9e/MQU3ZqQ+Yt9AJE0m1GTJ4eN5tnzz
gbIs7sj+8ZBk0tXlWWX5pzbTgAgNAR2RAY3sZUbZyTaahRDEN7Nk9S4hXD12XoGifsSRmGzDlRr1
a0xM3Rpa+ao1jGA4BKMSNK09rpeFzm+gQ/HiwE2WisNjQaDlCgdSbJbb23Z1nCHFKROsLk3QQzi/
Tw9d3CJWfu+C6ceMjB8PCOJlsSmY970aMNicQcSUOhXHeXSy+EAcI+HdWaVbWFVx43trfLYAr/pN
7yAwfraQVelAgxwwsR0ZQD0Rfo7KcsyOqPqeptbzIiCqUuUEbSj55ocvUFDT8fEA6nt3TmOxhsFU
aHcFoaQ6otfTyZKT7esRfgUXDEjVUO/gK7bggBepxXA3CjKgP3fEEVrQWtSwGCnexXoUFZDM77xW
jEaKqcIeN2mpYRmJjf69MWeakZf10dNjlx6lKs7D/6h87R6RJJ7885edRlASi+FEz339jhsnBABN
E74GgYiFfeb/lT2r3R3AKsQZFxWSCw4oqhD8Foky/QkAQDByIVzm1wGgk0mS8F/OB1GV0u5N/ehQ
T0bME0UIFl6oDnVL/pW02QrolES4rcAxVegwGrREWJ+zZwWalaxokyamoEtsCepP4ZqVYKJ1sqEZ
dln3o7Iz2rdKl0XAtFPeXSBSSFfyNP8K6s7Yw09CxO2V0aEcxA/R4IxLAOhtUmKc4KsdgzyVdbgx
GAnNaoNjVlLlaxR6lFE3x2c399WMO84nym/Nv3iCC8qXjwBJZT69XIl6DgKVAgXSGL5ptvFwgN2k
2ueIorG8SklUi6IymO7y1CKSqLb+IWNLCYYnwsX0p5PQbROh21yI2q8e0YLTuI3UJcFzjT1PpTHX
fTnFKX+5/chJUcw0bateOEnhOxLgBgTdOrmGS4YEbA6Mc/cvYmhGOhLLT33nf2em2GgSYoKWwEgu
7oLW9xVM7YFAOVQMLWb3urk/RCHQkq2u8K+UzEaQkO10XKxn5/8a86tLD42QBQyCaZFWYs2fyufW
Smf5UliAvAF0aT3KfUbLQ4nQT+ZRhL3H2u8uxn6zkbdu9IXLZ7fQesTUnnwMY9FM4N+JV46iV+8Y
owOF/vViuFbbgHuTZr9DeKeW9GC5ZYMKdXS3c1gfGOg+2p9LqDLFGKpeo8Gz6lf8PQCnZDaM1rUC
1wQRp1gdDoKfqUZjv4jqqXzsXVEN7ldKjMivCv4+pOul+SyyP3VRdVZP32dGuSqe1qoRhI66G12x
JSP6jJHzR3hjoCkYh9+T4RT9A5TA6oxCUkUC3slAuUoxoZxmc7rMkgs48LUvgxYpYdXmiaH/KQwG
5nv9U0KT4E+aSDMPC873PXmCI6nNHkxeVt8+ezMPcvlaBu+fgMVUAqBUkGC1iWbLpD37M8LB/Jq5
OxxHeznjx95/KlL66gkEw/vI8XtbCv2H9wcStp6UZdpZge8YtrNJcBNqTdizyzIPXY7VlyfxJHh9
u1/0ySQu53UU3cWRuARC8cO/UmuwoiBtwDDSt/xx7SEJz3pQxR3WTyk4DnJ+NSKeuIllS5mJ3VBR
he7EhleI8/AZo9eexUb2E09rpJOMuaaUnDucrTw28WWR8eYaEW+vjQD0WMxyN9JOD8Yvee2ccLI+
pwXRyoRkTPQ+1y+0ouhBQWU9yH+OP71yZdTYFjZ/r5GCKA5ZbtY5VvUReG7HHCWNIdMXJZILTHZ1
6Xu62IK+V91QlOzMPSgBCotl3j0wmF4RwS6P11zMhUFvXyFLD/kZavoTc6kFhv+OTJ57qHbHJ33R
CwX6+3DcdUqDCRp0gU6oZEzKlcbNxN3f9VUEJ27rDqLeyyEQl85hNmp6KL60P5o0VC1rdj+k/UgQ
f3s6VhDTTCIFi4010Uz42nU8eFtq2mN2UUZHwnw/mjFsJL4PowYGQIJxtjr7OYQ0H7NJaT2nFjq8
FQsy014dMV1AtMcu9sOezx65SfEU1a1Z26Ax7Dk2mhCadiHmV23/25wPFiWFgw++JBr0e/IdgKEk
adwDw+Dw47Q2dnapLhjOmmZoyRbrrbPu/KPcx/E5dAhIA7aOAJQshaVuVjNtKRzPz8IKZd+5lFBE
PGWJOE/a47g3eSHA0iYcFsZUAwNAMhBQ+Qcyd48cAAvWoD7OpXvg4giQUXFfY8JUwaYZEDn47/7c
1G3mqNC5oc6WubnBnJw7qxU4MPxxm6PAvZT61oAX6rVX5/USKJ0GpgiA6uttCfO68GfQcRUGL5Xv
V0AmBjgXPibTP38Ua9YGw4EIYqMe56HPIPHid4dmOXVyydVuaZNvmktLsMQ8SIPTQrGtLmSAS5Vk
WChqByRmFoMJLAmAkGdkRR+1P9eWhyCIodM71Xqv0N2oKwrOvgEhQpINrV/PFEzmhhtZ+oknoirh
PeYMS2Qbkwg8j/oZkuwBguvXOrAbKBk0yFpa7gUUmbxhfMo9mzCOv27xGYU3mzEH7P0rW1XFH+bh
voiTtZ0fdXSBqdPmHTeeiVC9Cdr66ww4F+OZi/2Z+6rBri8BfJeCH9uFbdmWJvgoMjhld14rILi/
GQDDniRrCXpdaLBzmDDEqCRsO79FtPyFBZv9UxJ/AbK853CRhRzME8H3gWMhN6L3NRv34TdR3hLt
Wg3mtPknaa/gIQjDCdKCHZ2VtOFfBeJb/GuKchCUsrRDi0O/SccVr4uefZDOw/2251QQiuR9CBK1
Gked53JAJvWTOBHGRJUoHN3LNM9QxpHV/phRAn3/G4pKyh32wyjg0qVcatk4z12+iXOeZnTAbgbD
KGCXhJM1t9ryxUmT1iAWY94tL7cP7zIftUHLY6qJq35mAkPsifydDtddIBlpcRfnKjGHWz1k5iG5
Q27g+gtmPVM1hsnbwt5VqQWjBacMI9gklgZYh4hw07mLOnwSUpdcUS+QRDyJZjVILy/+d5OquNZ8
Zm75zD/9JtOLSTk4AuK4eL/kAIdSRoMstLeJ0J1suz48HlzqU9cAy5dmEMNhJf0M5AU8y8qHekLN
F7OBQf+4BuQEuuNlPbpVelW7jO0QnJ/VJsu2oeU9BtOivFdrLjwwAk7rIBcD9nTh2xSHPd4xGlVQ
7OhnXLfv+jWAyKIaOYh7m2xE9N5b7mm5U/URtYYwSnGjQqdyEoCjfJw2HY1TX+4fFEPF9HtEzQ7b
6mw/nCX0yy3ogGEjyyvhtV8/2jxm3a4wsgwye/h1UT6O+uKfvpkjoCJnq9v3yicKd+gPlNh1R7tD
rqUqnwJ1Eb7ZTDuezfyOJ0OaaMZ4MZ/0UGNIly5vsmlzyn019DZAfOVRam6OtipMlj33g3ollSfg
ZBfTK+iJi5t+WLcap4e6v9P/myyfiQkkuiQ5BJqyJ3kMOTYxmG0jrro2T0u5nmhow1ga3Zzjinmd
rIQygTpBmpMkHyJFK6iaM0E1Ais6jZB/co8Z7aEs8HNSRq/s8yCkeOs8G2e5hjeWC+aUhXfe2CZH
BUMNg0YgrsW1IfVuDHJwqXzNf1eepo4xuN6s6Is66ulpBgQp+JGZrqgdwNYFNmX8T1WEPOCmmtDJ
r6azX0/NCKg6jcUDYIQEpvS7IYdHPSQMYn6Y2zP1WHkgAvQYrJnxlqxc2HrIYISFKMP4T5fEsBqQ
zCQ0bjlDwv9ouYOJDaseSbc+2ZjAFf8rCue3wu407B1OGB+0snoxBaih9IWlPM+QokKNTZiswZ3Z
OBOgyQpYtfH+zo+2IVKIPExL2PV/AZc90fgVu6bCHgrYBgI/oP/rxWejQDEse52+rvooYkJbWK90
ULC8jFrz3cOmtF8qcaIzMhDS4tPFn2jwPRBeTrKztl4o5yvOytM8tIEYr+ALW+zPrVbBnBnbqYFD
/geTdgg5qwhZI0hECXauHDdEbN/VaGcGFIDCmptNalql+/WXaOZFj1YJpUCCjGKiGFcy7ic8ABKj
9UuN7OWqfQIwEaEPT0wQqGJaYWNBfV+VhbErOre1MIbvopwmi41yjjGKHjQnFt2S9ON88/fVTz+9
eVZEnVwrkKZ98pkWlJbh6lw4MQcrhRo0pMJP8Gtg7P5MR+JRN/zJmAhwHj0VhnIGQ/AzsFFzJxSf
oVVOuoqOCi0HOVn29gbQvWeJaljNO0IwtS8UHLepfO0RN823TURKwKiDczWsiRQxOv0j9Y/bP9e9
hfwr+tltqiTbqGRUVpS5SWMMmNVcLECmrHyB2HVYxp1u1bbcYfguRE8QePm/mgalzXrX2aCagVhK
caWGcn233IVfTMiNSnyfBCyUsYGYrBdOhOlyc9S2nom9wnvIoxyJ4S+Ispe3F+2WMBbYOIFJXa3w
F0+SG2TGdpEFJ9TAAnHdd9ch5L4liikMjMyQY5TqyxK5Xxt0QAwojExwlQ1AoyFPn41HbHoHiWuv
Kd478Qj6emzRZfKRDFED6XmCK7Pc4QUCtXdKn2BopSRS4bTuh5SROWd2r1HsHHEMrQ/5cFbajzCH
TSiS277NtsQYv+xpWPDbxF90Io0hl/504Y4rhcRKdEUC4rWsASHZZvE13c6R0Lkp/tTbGQTZFAR+
d+mjdAFJfdLKlRIHwVFZWDYlg0j0C/SoE2zz4ZaBcYVGQzWLUnegbYMyEutnEmaiW3iuLDNG0Q1u
236dYF+86jVeC7kfy1Co+bjNwMhzmTZOH/4QpN0meNnEtfpAGFfEH7OoKL2tONM/99p+IaFMUdKc
q7brAXn+OQ2R0PjaFfuw2wuzgv6iezSs5J7tm/DTC+DvOThO3r3vyGg6wr7SVts2g9ZjodGDewCW
VNweXUue2Cn49910yZRsTSRWRZ/vOqfxs/sJwQ8RbIF7VQVMJPlAGbIrZU0CPB1ejeProTws8fci
cOwkbr9FvXeWhozbz7NA06Y0L3eaEQC4g9lyLTybcUb4PGSuBqqvV6U7FuxUCLC4HKoyZTT8NiEF
Rkl6t1NcMq+SGuo/hmqE+2624/WU+/zeTz6OsH2TEGpDPluS9HgS0gUvQgANH6pg8XOHv3EqR+dP
zwXYep8HQmvQGBIVvRFK8BuZF3Pw/WrjqgKO0sBOorIrcNvyruJMlr1SZHGlWQuyFKFskQqHavHZ
66B+Fa7ENRMBqCWQ2OzQReVFYF7xkKldF47IKbOewN6vRANnxdPO8jL3Uwf3ZabkOAFBTn4hsPR3
gSpKtpr4O5x69wsi5FYY/u5vliZlMksaB3Vncfp+AmLRwMum4sCzTkYQ5C83HPM849mVLFG9xvsq
JbzoYFo/XV6mGiRRIxeV0e0mwHwUiaOEHGSe9Fuwfzpc+AH16ckJqOQPcLc4QZzG9+n4KivHyAts
LS0+QpPjIxpGY+0FW6rngBrF2osawRxI8e00Kaj4okDJt8pwrSdAb36myBuwONqYyP8ELf8cGu7I
ImcRj/nfal50p9E01F0ga/SQnZNwJZyVOF+e2B2WD7VUenFi3DMaUbJIQdJGeN0pKaXBIIakP3Cm
biurgNf7DDyFIiGla65855xEHQIEABl+zabq/6pg1R5ewMrujGx6hPaAfj+x9xwi81oFSkxZhOxx
fMF2bKNO2Uvlnoydrwzd9zTBT3oF6PjFngsvqxdmL/UZVcDzgA308K0ZnYeus6I1fx1giFfMxTWT
HGXgRBqJSKT0GQnir4bhaY5thYYb/DQLBgZxzd/iesnLOpHDtRI9Aqz4MFAklNhrkrhuZHQf1TUH
iccvojKHSEx03zON9uBzB2k8HUGYutu6Qs0tgPRYK2a0pkdDjdHaOLvAC9leLyXzVtVL1/Xl9Q6B
VRZobURyrbXtYkj/OjGtuBkr9ygEzOSJ6LWJKPp9PcQeQHZx9VH6KxGFLcMtGJd29dDoU6p6vk2f
J4vX+tbctkbrlVU9NtyDMc2TUIl6USWBAUwv49xSE8IwfPYBL/HoJZE6raQlaUCAOyp50FZNAu3c
UggHm3DXl6/a1cZxfDxvrUjJxHCLoy98z8DzuERuTkdacxh1j6VtMMYCis2ajxRFsHbjmBZQAO9i
laY6BoEHzpDl+MT3nPZ62zXuVIvtc7Wmmv4Ne2YDnQzC7sb/Y8gaOisB2hhWamFKyVLN3EKCgfV5
h57K+cU2FIfrboZOQkycSksGWfAaRFtOhLruCWS8kcMS376rS6MIotVwamscU+cK7AVWYRR9u4IT
CV1KAc/fcFLPF0vyr0RGpURTukbuYKzaDLWTZWuvPTLEQc5CiktQjt2OGx0mkSx7SK00U4mqu6C/
r225XpvXeEvcJVTHYwxmtDImsZhtBpi8RFpZmlqx2eB2anRDS8M1p8UFde62+U0Hw7eJiBCdkwv6
5Uuh2nbpzEpma2yxVS8VL6zyxh1+331AFbGsn+GVluwZrfStjhOfELVWPpEcSQOjZ4EA46g2/ml2
12vjFr+MDa2+hxW1WfdcPUvjrCiQjzRMaLYP5j6gtU5ltRhvQiwEyij/SYLDg1Wy+MLhKCZSnF2L
nbl2kBjUiAzGrKdAMiX0pUpwDLiWZgg/VqtS/8IPhJ9VkdhN5sCe8j+OuZiVcUbDA+MjK4sOrT+S
xE65LH3IfE7wdv8vhPkc1B1/0+RPmlAZJF1+5Xdt0Fo9iJHS+p6FGyANvLRIKUOMmYp8Zf6QCWbr
5dQ7AM2+ErkV8Hfe1+8vQ7BaQwKx0/znjX0bCtO0Tx3CI/osHtJ46EtH46UD2WjFaviRzwPouQsI
omhPgi2fyCydt09Lzfb0fIMJnK29fkZwGa2PAECV92INEYBQ75rsevtVqzhDyl14QTIZa6aRTvJU
ptEPA6aIntQJ5KzE7xfj+cTDKDt4DDqAQSGOG8w+ZfWEnf46hIz4RWPDXVy9GOGF+KGmaGpDINWv
GS9ovn8F4Ba8hCNGFp1yKmqKER3MKhrJgNxe1fLoADBVCrZoCbf2QX4tt4oPaHenTbICytAJSaFD
g5e58BsfQzBa+4XtYn7mBZAev326nt3FUf6I/x5xGabwCtI/CHqTIt4y9DABcy/qtV4K/wDFCBYx
b3L7SwWfQWdEw7YPXFsZe9ix70MNf1IjNHl9lnI1+2Db6te7wluj+O4dsoxHsUHaOb9jSOzAbIoA
CjRarXeVxq5YmjgNHwO123DZN0jYCFj3rVUTjHPA/cuo3rpr8aC3U/WsUrHcVoKYc+kKQg4WRp8x
z34HqBl5LLcpTJ+nj07bUKpZoEzm0qyw3ioprlZjFOgij7RUJ0tO20fuAm/axV/jUYC9F1pTOuOf
14nYGxjAiyAheQSG5LLIlB0eBPNa6X/zSKKZBZmRDQHDPwB30FIXyduTPh+9h/zOCrif15Bh7jw8
eO86gJ7wNZwYwxMyCh0h+ViCsvRXurJbQElQ879j1XQ9cFkPk3qCv8y0fYPe0G8n+SD3iObzjvoO
vXasmzs8rnYDZ7aSFHjEzYWI1g96bXOgjYUzV0FEkrJcd2pyv54AadFKcj3Ml24yphaLOL/ZlD9J
u/VuAHcKHnrTE0iV5qPDNhwkQRosckg3GXO91lLM+eOtN51Bo71TrEcSsALRsBZyZMNNkYZGKZSz
i0HZ/MzrQ0g7ptjU9o21BXJznioq15/3eDM3HdJIm+ZhRG66QaZ9qv8PeQgunrYd/Xf6uMrVyIwI
0TBh2OjLQn7O1jJllCnFLA7249J72AW4VcP+J19y63CfCBR/Xes5k/vcEfyGmRn8AI4/WFRsGaq3
osquPDwPPYsmCy6jvPqDNCcRd8jAITfNoCRJj7CTg3Iz3IxlsGVg//cUW/pC4IZox8FMe4rvr/1e
FD2KVfof4NAbA2L4DH5kQPsgnaBbtxrygt4M2tu4EbHZXkY6FXxxO6Z8T2yoOur6HFbbWYoo3bQa
QwzjHQiqutd01+DmPXCmi+CgSJi61HeoI/lUQNQasG2IixxB070GR3NMiqKgWpgHcVjmK8h6uWLp
L4KcZBTZfGviLBcYhrePXK2S+bdyZaGR3ggvVlTS2g6bW/To5y8XiCFtfZzgDZgpl1gYqnlcLckv
UhdZ4cTbD+jRtafhls2ZWgNr/2NBGPwqB4q8hLzJiKHuztlgMLEUsoiirpa0Z8PX8u0+dUyoYW1H
7uiCJru1WGgQOWPQ2HE7Y8WohkSJrtvtU6Jr/p7/7hcnnG350xTY6OilEVgSMkdFoHeo8nAqQf08
P57oT5kGjli6fpmMh/lWE4UEpUbRONQZUDAPdvmTolonHrM0a3M5SeIdSGp1p5YjEOQru/k9U4wr
afSRrxPU1nxr+FnMyfQ9BoTVdx31UhKPJEh5yQAUsdCHXWurQPVAitJtas+FEave2Bm9Q9tMvMCr
prbd88rWjmwjGeea804ch86olrJuQ43ApBlZq2CUi1hzPSHzp/DNTdyhwou5VKcf7HNRuKWMbASx
hjqRxFftEAEhoA1VGHhhJzpyaYIUsmljCAiYOcrojqwGnEYupQvTNGekhEH+tlQW2grAWtzsuG4x
0b8cUsfvu/q/4XT4VYrtRWYOlyM2ABAZA+XWnm9QIoDxDkzTpUIAX9RQQRjAWMn2ItKzBIPUD5nj
3/TJU8mxuIv3yRYWQK/NldrIzAHJQhEpVVJfXCXp2P+EuOUPAcyNHVgPAv/nN9WpEhMGRWnMZZTg
b95/TQ1YqQuCxSbJw3vb2YjiuF6VJU7ZCucndiHlnC3UtvPU/nhu21FUzrwGDAK4FIJAJtidWqk+
lnDh99G706GB7/EwV4I4qwToE3cDhVscqHoH1t4Nn7911lXqaQ67DQWIKZj09SJ8ffAVF+Y5WsJM
6hLF+ccl0zdXHrf4XpdbxXS0ut8RXlC1SwnsK7py6PxjPdoHwnoJfE/rmtwBBsar9YXf7wI8dAmq
iJXAJnEo7krv8LajWO6djhKOA8+PjElxFOzhbGlGO4IrAu0bMNCY4mTd8Tcpm415cLV+QXkg/WTq
N0+4MLbEVm1DFGFLHZ36tlF3ZtTsONb7xzUa/8hVu7F2hmWH+CDXFjYEaPWpUdk2B0ZKiZm6ngO3
/dkPMlIcehQRK6I3Klym0HX4hfNVQm1zvUqmEILgQx03uH+rSChjHQ6H2kBJTRxQjC2eo5e+hi6l
cuA0X9tpV0SosmZMty8lczx9lwuT0nMxq4dWnNJtyPTOnYtsXtMyjKRmtYHxNDwRjdXGoGF6IbNc
DibaMQ/5bjlaWujHvgt+gyt2TUouMGLpycJJ1wMnuA/hd0WRjR68PjTjrIRlxo3EXrVJkYvemlAQ
FFOz3dvZmLv2dVO4ZQcXySnqZaUvy2fjoocUnmU8RwZuMo3c1VtQzbif5PbLddTrX9ABk+31/WTQ
uMb3A01vz1wLNvDjxC53ZNF7JuiziPSgM1M8uI2ZYe1q0pLoxEdXK2vM7taHEonKfcTwK6YQe1kx
vYexm35jsTWoAz1iNYlSHVWEqpHLuPEWlQeLIPEmJXSkLoG00eZfbuXLANQ9vvf9PWagtZwNe5XA
hV7RuYqVwrMFrQLxQLSTFPzBpdBHL5ad1Ptu58s+dQ+76A/8E2vbLko+iYk/S8sEmbVZPYcQwc3j
yb0u6siHFLrdt95ZVTYug1wV8t9CWNBa6jjOpporL6M7zvYvkph1vEVb0RmNkjHRHF/SFsrMkOMk
ckLRBQCjjeu8NHXtjBhjQqE2FBg2Wzud0ev2R2dJeC0s4r0MXVfrgnjgVZ0diuN6dYyehWgCmHnl
oyi0Inb6G7Ntxb+wTtpcLVXaM0yAv9jjZ0HvG8FpFlaVNE3zwOZwQl+k63wV0cyJJm0bCvTTwwQ0
eurv0J/htNI23YUDmDzdm6pMIhPxE2PpRx7WwVcdzAjSYCVg4REbtF1nigPfuXU5aySA8HvGSAaO
0Lwfq68Da5aAoEUN2T3WlkX2gLUsNhU7QcCybuevN4dw4iA1JD7y/aDbOiIzQGyBXpEjRaHHhWj8
EKI3g5zo491zK44c47ck4uxQlmvgB266Zper5T9xfy/Okc1FvyTjxaZeBc0SuFPJqmRJTIbT51h/
wR5oy/rWaXCVv6F/uef8aVs4vbtZm7jRjf61p58jdVlLILuOSDTEpsyWH+mFAM+UKag59y7iwD69
oOeVkSqqnjfg5X8okS3JlYwJVt3NN7VQrOsaSfP3qmlj2WM4RS959EZtYjuvtzBJEa4DH0QyGt91
Jj3q+Z4pI9bUlCZuJHSa7UsFrfNtQVEZ55ICQ+5LCB0kRK0Q39UG41fyTUkG3DIbA60vWRaPm8XN
hrBPQYndj/2VGgY8Pm153kRqU/LOGJj22a8usec6RPyptxayN6UkSRhzD1nv3dfBfiM8lwi8CNHX
teMeccObbxDdQXUlFfF0pYztoY6CZ6m9S5NjoyUCCFteQ5MQ6gQSv7OXtvP99+fuyHA4lm+MdAx7
bJjB3eRCLQEXQ2QiZJIMZUZKRaESpcv+BB/WVpvf2kK+9ekXVkFj8hQEFUzn6zQ/mI+nTzGiFXvP
qLwebBjMy3rBhSl2aWckjXcNFGzJmBB/nVWk+XKOrLX57t6AHa127N70BC7toN2mMxsM1mZaSebY
Bg+Gx+Vz3w3OGbFew7D+303s2VOHOKi+aPJbzDp6xT8eDQzpBW0H3Ny7ZmINzi5fSr0CRn1ZFS3Q
LlN5MuBPHo1drGfRK/r1G42i6eGE3/PQN/XQoYqlO1tmDxL20xJlmyKgjpanzDkVUE8/kW+XqV4T
98HE1OlCjrCvyA38CQEW47+jTpoul6c17akG4/661W0qcBOMLbbQyHDJPvysp/6wHhfFdIxBPzoH
QOeMXJLowF7s/+Ae8MABOQ114hAFs0Dova8tVuwkpBuA52Mz8MGP7Hnmqzyaxxk86UHC/LEP4MkK
RLFTPc18D20mTD+fuMJJRlOMZsEWy/8gnWCmxyvBcyzo9F+RLF1Obxj74i6wvjPK4z9By1aJalAg
gzMzxmb+mZ8HGSmGhGWf5c9tTOPAXUElM/Ja1K4tneg/A8HDWKTgoq4TuAR8F/pfhLd43xGQus4W
81TuGGB9u/4fcmtfXMHfMLm9GdwCcMYmQ+JDtuK4wwFja8ae8xAn1QqqiW++8Cd8GscyAemmP171
Lu1eNGYxeOqKeUzYsUs1YaRsacbc9jxn8Gb+ytoEYgPe0aCDhpW2Atp7BrXjlxrkYat5PA6jX4yP
7OFSsAlpH7w7MP+8XiOgax9wWn2vWVzwF3GF7iYGJEwPXJYPeiRhGhSfgkLkLfWOGm2FbwTOw0jM
NT+3Hb61hfFqlB5xd3hwSGGsOEUGuOl7XkR8RBFtxmAiHDhPtYyjMKYPDvzZ/C2N4IAeMbHj3ViA
auG7l8/9rW4dRuQMDYKK44bL1+UFhhO19M/i6EvrbMxS6fAuKJv7le/0ThzSy6ZytbhKSontEW6H
fRqthmKAJ9gxfU6VvFjSQUpwUz7FXBZXBbA4ODssa7ho6o79gaTBzcTT5BTGO56KdmgXbOVD5BQX
BaLCkuYrNRHSc5+tRnmrN2e3moiiqzjNZqamKijhCtXKwx5y2GPLiUqf7anTSC2L3eZQMlk8nBLH
Nrp7ob4iiVpQ4nlyupqgjSF8b/DQIfQOas6n+k/sWe8q9KljuKsRd6RFo78+EFe1phYhRp5kpeq+
p3MqiiyD/GX16WksdKlE19J/RsYUZMidVLhCEj1/JPLYFyDenM31qKlGbcOdJqYocg8P72ZYoDQQ
Oa7B23AhakIYOPWZI1n7H0PW7z1Bz5F57Tq5IacrwYsbnjoL6A2A1KDlYGkVeAV8M0AkSWXOj88c
VhJNpFTXtGMKYS7B90EXMvA3XK5KWs0i+Q7ttFYp6mSb+mQiKufKR0VjQlm2LtdnBpPXX9OmHPoj
zYc5G6PNt5Dfg4Po2ENfe8QS3ChozW+iFsrMGK/Wd6VDFFMfGdaW34zrKVUV81SBx3u5g6DTqp4W
YP1rsy7k8LRSRJG/1J2sa60yczMui8IRNwedxqLVizbicP0y+50WyISTZAqnkUcIEBhNHW1HmI+8
CR58dJ0TGXZF1a8FDz0LdQ4XXZpJqhtMqxsJ7IH9IwIRM+KEz+Pr7Tz06Ut+ZICMCPrPx1B0TCmx
PH4yz+dvisv2p6ADRWMEhnelEg/JQTVf519avVwyMVKT07+lzs7+uLiZY32exUDreOLAE1QUanh1
NvFV6UXU3qR04TuxRHN1I6FVxRhWR5JRSFi0mBm5VP5P7rV0zkOFkH9gSs+C+VLtbRjN6qpURBfD
m4h2Wel41G3fCcdIcREC6ZMcrHnqVJ/93HnRYJSHngDISNH4KJFGUdpxh/q0H3Fs2BZenpIiStuO
7SeW2ckTLa4iYI2UIudQglx5zn26FvwRVrh6lLG6K80K9ikFEC9d3zQApjOTYIO/exJhCNM/3fxn
CZHVbHpYsBFZtUNd55R/ZjtRk1PbEKm8QvcW+D/5PqtvtuIiUlLi5Bo5iZABGkjVDkZxfodfGzzE
1m9urzlE+5Ttm75DcBQfQw405X7EOsau4XE+luKhpuY4F9DWefk=
`protect end_protected
