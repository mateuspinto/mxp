XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Og^�������T�/��7�0|�dx��<�M����	�if��q�����6k]�E��{��9��uJ���7�E@�	�7���S�C���m�&�"\�	=�ey#�=/s*⹂K�|X;���k'
�醃1a1��L0�r���Z�Y����4]����cƟ5�����Lé�"��^`|u��w杬k�H&EŬI!�p��K����8��^3��@��D�턘Q ¸4�0��A����j}~8�<2�8'}��Rq�|Zq��u�6���eP�+�?:�����*?>�J�S].H��~��ൗf�[�z��v�W3��G�����2���y�P*����P�Qb����0n˪JV4���0h���8�k����(r^{����K)��	צmߘ�ŭ��	/̓��I��YK����vw��^:�#&ɥ�b^��cB11���i�rzˤ#苙đQ	��m����2H��7���ο*ܖ<�Gy�fQg_U�ym��B��f�\S|�P�!�Y/X������-eov��d|��:��ϋm�N􇸏J���_C,h�@m��О�����6M��\��:�����Cӂ�m4�����CNR3��K߅�⯂�o�k�L�	�=���I2�6`00m\�s�Z���~��}v%-��Y�w�bڍU�x�`\]H6��-�M�CPL_\���0U'�l���=#�����E�����^�g-T��
����s/�s��|D�Ü�����~�����t\$XlxVHYEB     400     190�R"<�
�*���wV�4wT��!O��<�e~e@���.�+�k�Io��9v%U��ɾs�.(3�'"�B�;$'vh�xx�Z��.kfp���@��/��5��he�=��AY9"�/p"h��a0���,H�Xl�M|���p��y��x$R�[6�������b�y��M�5z������pLk+mX�L~�+NL��Ih�`��o�1;����K���	|�瓨�����ID�J�0��E�����Y0Hi�L�
k�b���0��k^�ś޸T0�����#��@ܢ�}�ur$�*2α���i���9�ɺu������aF�|������
���=�h��{��zWa�M���6&��`�v�i/&���Zv�"]جW��/���XlxVHYEB     400     140��0��5����&�E*I��a��ҥ1@��D5��FXX�Z�_�m�:�֔���<u��@����@�܏�L��хO!�����o�܏V-o��L��R��taxlt\{i�1m^�&=NA��@-{!��	U���g�v**"��*�*AZ�����h�O}k�*�P��ai��s?6��Ҿ���/qZF2k�q,D)"���*6�tӆ����oQt�Dx{�oQ:�����I�K_�&
`�/j���7��#�Na����3��*@��^�G�<��;�/L��h�<��P���n�r�s������&Q�ʶ��I���XlxVHYEB     400     170�� n!+��ǐ&^��e�n��+}<i��6a�E]jX�7�1�%�/�Ķ$��a%� {�(r��O��K����9�>mb�Q"�����_�Zi#o`ҟ>b^j�O�~�<�1�ߪ�%�Js3��tB!jbpw֬�UmpFï�E�����tX�CO�#`Y.��ê}mC$��0l�U~�z���ʛtW����]�(��e�ݫ���0T��:�����vYR�r4� 5�"��<��q�M�s���`��p�|s��)�D0Z{>	xn�����g������A�8B��ڞW��$NY,�&��r�AE�>r�� �4����zG��|���������V���� �,9l�J`�	���w�XlxVHYEB     400     130�3O��D	Q�1L?t��F�}����v�U�m^�#���F��k���k�uB�l�Y�80�������F�׸G��3^_�uT1��T
5���A���̶QS���Sr@V�F�zѬ(�,"�!��U���(�և�;ꦄ�հ�R��(�C��뫈���>�Yb |h��¶�$�e��Q��#5^��$��B�=q��(�G	%������&#�K�/��bxX�|��
�O��.,��珙�Uu흉GPN�]�z�Ui���,|!N��ț˷
��C����]3�r�G5
>#�XlxVHYEB     400      d0恪4��8N%�Zg���pxG�U��j��c���f:��Q��ZEXl&�wLR�ʹ�F��7�&�+�}����y���\P���k��ֆ���Qm�1R�q�7.���������a�XQ�)����KX��4V� pK�?i�E�'dnjDh���'��%g��\:��R']W�39B^����������� �����T���O���[�"��D��XlxVHYEB     400     130��`c�CD�u��i^�cA�1D	��ʌ'��e[P6��E�롕	�i�)(��/8�[��,z���s�U��ϓ�e��(�_�P;:�`�`̽w�G����*�@�|)���p}@vzpk��t���]�) ��%W1�����^s��Ӕ6k��1E��k��ڑW�U�vA����e(��kU��W�#��u��=dڙR_η�v.�hT������K|�
;ah��o�� ��v�V����?D ċ(��w冂	eЍ��$L�c��+��ʐ�d0¸��Kdӌ�:��=���#���XlxVHYEB     400      e0�2��v[S�t.��bµ��N��+
�'e�R�s�&o����[�W��r#���������0�7�-�<�;Y��q[��2!��L����B��0C$B\\$K��ci��E���3rW$�q�m�zP�z_*�*a��V�����.����cu��Tm!50ƥ�6s3�3����
�̴x~t�N������r�k��S�����/� ~VXB�f܆բ&XlxVHYEB     400     140�~�֚�|R��׏�3��8���)��ӧ��(S�}^�<�I��*���A��� ~�ͽ.���+[�SfÞuo`^cc�[����s�z�v[t�:K�0�>xRj��z�@��*��j�ڑ��re����MK-3]����A��B�#/d�藼X�?8$�=��?-u���t�S����Z�Q+��rR[��1S�sԇ��V:�6�O	���8�~ۯ���?��䵴�>���k���M�s��*bO�ϣ�2_�:��Q�Ihg����? ����V ��j#䇘�9NP���RB�D}���I7�.I�W%�m׸6�KXlxVHYEB     400     180]2h9�����մ��H2�I(|��=��,A��Zw�v�����9�*�x��f��-x&�Ԍ������UQ���K��h���f�R����a"�p!A���%����7-C��BYC����h����5��UHdYA�8�<VF��=�����
;i<m���g� »���v��P���� �>,��S�E��m|�h��Kcc_�Qv�����U�E�Ǧg��"L�^o�a�FWM*�p�@琘�{'q`|�g����-��j��H�����d��E7�P<���~9�ׂZ
>��Ĕ"�X�paH*7i�ʈ��@U��U�1����e�@�&���0������79�8�N����OO�wY[��a����%@�n�U�߾���cXlxVHYEB     400     150�4*�ـ��!}�q�x�P	���J���!��X����nm#��T!����U���J\�d��s]��e��R�\���Z,r��oYD�?	�l/��̎}�$D|����7�tw.�j�ns�wc*��7	�r�0������aL���� ��kA�~Q�@a�iq8�:<*������O�4�&��u�'�d��! �����E��@w���6H'�:�k�oqޠ�?�+���2amb�rJP6��)
S����&��wF�yak���.��9(��JjZ.�6H鵻�HE��qu�pk��(�t�Oښ�F��N�:'m��G	�e�s6��H�K+��XlxVHYEB     400     160fؾ�E(%�c�%�L�a 8g��]�]qA�����&���8
bw2��>W�|�񇄹�g��.~п]'��?�����ߎq� ���4���`��͌{��k��W�>l��w��y��5�Rپ��4���W0ȨoU�Az�������Q>�y,�:�]٨�OY��c�m�.7`l�0��v�||�� <4Vn�L�OCg9qM���Ax|�EH\ȭ�l�f�J��_A`��#i�3�1;M�];�l�o���(b1�Iz��G(㙻˻z���WoGo�t	�V!�ek��8��P7�ܮ�C�J �q��Lgp�a畖 Q!�LV$�o<43������)�f	���z��������XlxVHYEB     400     130Ǘʔ����S�j=/��Lȟ�h���F�Pz�#�T���T��o.#�p�����ڃ����Ko�R�������f�E�aף?X$\=��w<�h��.�KV�`��熱����i�������A�Q�� ��� ���
���HG=�2#�3��,��1_�#�r�y-��}�m�д�����2v[Ks��/��)�P���;�^8�h�/�|�\4��o��d�H	q�(��B�|�`54�e��<%Qϑ�&��^�DrV=q
��79=�D�����z:)�[�յTXE��RI:�XlxVHYEB     400     140�	�����}Q�����L��.���Ʃ�{/lP�����;���g��r��}�����&�>����~�Ĝ�Qg�\��;42;�J�z�y|=m���o?���R6x�� /+�[m�#ήU�{����w�⨔���7ٜU����r@\����^�s���鸇����c�޸R�z����po!I�y�L^_0�6�w�ָ�������'������߬~E�󇑹�:cm�R.�+j�.b�)E]��N޹2!�kW�E3,�CW�-���O�\=�J,�Ξ�����}�B3�A����$�%��XlxVHYEB     400     1a0D^��h@�.�d��ߌgϹ�@°�}�㿶�0KOe�H6��إ� Nџ!��?,�,].�T�n6�;cxw��c}�z�8#8 ���r�F��NP�Ԅ���`��U{և�w/_K�^s>�5����tZ׺�z�0O@��?��u��K�y����k{���/���%�L=��"�R�)��IJ�e�a��pO�Y;���A�*���3'�j�T��`�G		'�BvY@��L$!�uӐ�G�=Q��:��}Eƨ\9m]�iͻ�<n����"�0Ջ�P��K[�.�*�ܲ�P=$���+6H��JnE�2Wk2W��c��z�[�لAE�I>�Cv7N�~�|�S(�# �F-|*������țChҖ���%��)%�幎�y�y���X:�8��Q׆k���ʥ��$XlxVHYEB     400     1203�a�s��.3��e�N�����rhV���w�w6ֲWտ�"����A�L2�
J�Ҳ�j�O�*��NPn,����Zh�w5V3�d�	5磺}��v?{�a�S �h)��F����)U3Rn5Kx�L,�A��d�(�fAκe-�]^����d|�((��Ʉ��NH�<��������{1��xZfї,{��Eo��l����K����ѱ�2>j	q�͠L@,�������t�Vg�;�$����a���iLF�	6��vG5`�m�R�)�
_����XlxVHYEB     400     180SP̣z6�T���v���k#��gD:��$�׬�}^���`��[7���ם�-)6[�'
" ��=�"��x���R��_�������e}��t����M	�B�Aa^:�=��Ӌ���G�˴7����Bk-����'�H�Lo�&����.�+��ZH�?��T|~�{�)�U�I}���������<��у�F�UŞ��ϲ��2o�Dlna߾��'l�{}��� =.��q���'�P	��Z�H�(q�M�&�i��&qn Lq	e����a	S��o fZ�]v�,�H(@P���3�)��~EpX��.��	�S�Ce��4?��h�MI�� o��S^d�um�@1�+����x���#�O�����s���H�#&��A�J�XlxVHYEB     400     160�Ҽ_{���s�.~�ƚK�Ŗd4�ԏ���g=�/-�ԓoX�0!D/�)Ε��t+_�q'�p���;�e-�%_I��9T�|�uhv�8�y�u�K<�ͻ����ń�M���r����G�n���|.v����	��؛�􂅜��Q��6�+�L�Q	-@V���$:�c�:��D$^r2�����*��4���ǐ@y��`<k<Ń�3�]�ǜNT�e�jD8��90X��y�Kn�*��ثS�j'(~!���
�Pa����v�0u 4��M�[�7�`�jA���C�C6�#����o���C�g��Q�|�?q"��K*�:�,���w�d����t�^́bZ*RXlxVHYEB     400     1b0������8�{��7��TK���=2!-tV\T�mp����iDVw#A;s�����@t����&jF�w8�E���R�9Q���E,�x����իc����.��j1���s�*μ�eOy��6�mL��ºIB1��m}�.����dL��%Lb�Y����G��x1&�����)���Wu����h���� I�������_u����e-�CJoO����*બ�N	_�x?�����}����-�*�E�.����6	�%����K�?}(�u���/��2�~N�\����'�'R��ۄ��B�0U�ӼN5�(��%�k^)��Jw��4Rc$��e�<�t�a��M�\��z��a�v*μZӅ�U������QVTʟ�{M�|ܕ7@�	q�|Wr��pCA(L���~����NkRȂ]?�XlxVHYEB     400     16008U�� ��?�NE?�)I�!�zO5�t������4�ut7d#p�MMO=��C�6f'�Io��T�de;�e���6�*��F�\$y�O2�`��bZf�����|�XiT����İu�)?<qιT{��R0�$��=Ւ�����]�c�F���6[:n��y�R���酌����	*(�ŎL�c�N�o/8���XrI��.ٲ\�4oHŀ��G���?+��������IBO���)�I�x>�0�#i��8}��g(�r�4�e��g;�+5������ɀ �%��E�y^M�/�eM�Ѭܕ�5
d�,�[�mV�m�Z+Gj܂�9 ���>�՛���ʸC3�h?XlxVHYEB     400     130TPT�^�i"ǮIw������v�L�c�6�P� ��<��M�l\{�� +���84��:���J����;{����㺬�WLHw앍�� ��g�gw%�#�p=+��.^w�,{�=t���Ԧ�>��	�
�_�˥��{�s�]�l �5�Yc�>i�|�*�2|�"�C4-�szG��
������tY=J_ߓGS��Ȫ��\�� O�	f@Q
�
���S2������-Q��6顥HL�}�uq��o�I���d�9�6��,�k��#������,u�Hjِ����Ed�%��I�x4�݁���d;�XlxVHYEB     400     140B�-��;o^0.AZZ]�L�F�V���S]��0M�����j��������ӼY������ͤ�Zo;��6�L~�o�!��}.� J�Ҏ*���-'���-?�(}�ԝ#Z��;\�`�E�#��v_%�����U��p�;�<���'j�ۍs%Z(Y�$H�.*R;�v�1E���H�w�������WP)2EQ���;[l��v��]� �Eڧ��w�����.�P���F#�*Ђ��z��m�����SD�v���T��cy��p��W:Ѻ�i-ԱJ(�4�ٱ��dG�KX�^m��ڍ[����"1�|8��|̚y�SXlxVHYEB     400     130?q����7�w.V�	]he+e�ǆ�z�
8�49rg�<�!�+�bl-�x�����.zbJ�L	��:�̇���`���[\~\��G�t6��l��R�ޑL���L��=��E��Yf�0�t����+:���
�w�T�e�]�]B�&z�Z���5�j��lM��=�?��)��F���/��.21����,�1Mf �V��,˓x�_.��Ѓ
	�����Q�O5�:�ݺ�k��d�%=C�o�f��ߋL�b�r?%�DA_$D�	CC�/��i,�F��F�8}ւ<�(1c�j�R	]18�}��XlxVHYEB     400     140��m��AEﶚO	A��hG��
6NG��wT�*6���s���Y܉l�r{`�H�U��㖸~=4�.%�R��<�<�ư�s N��r��,��?�v�RaU@�=?�̵fFidWџH�5����L�#��2Hw���ޭ�܄[z�E�w*��}Dx��U�j�u����bb0j��w�7!�ȁ�,.� mP kk��(���kO�m����	e���1C��G��?9�Ef��?��z�[�]v�)���v����Wc����3�0�/2G�wLki�1SL�4�%"��R�(�a�~�U��CN4^����XlxVHYEB     400      d0�`&�|�X��s����:�n5�1����CH9��Jk�V>�)��"j�XA�T2n�6-�y͊T�ok�3�<�D� 0��i��0�"R�ٱ�g%0N�eu���T��EQE�a}l:*�(���g�\��;l�]RC��6�zK`>EFߐ
��o����3%�� ;�)6���]�&Z/��e簴�~����@�a��M�iS0���(�XlxVHYEB     247      b0q�d��7`{�;��ʼ����i��X��C��m�<J��%uu�rb(�L�V�ٔr�˜�6��6�A��u.�����Ti�ۿ-����e�
�{���f���� ۥ�^�H|��8B�X��^2��o�9���w����fQQ���8�4�������[/�{���&ʈ��B��h�u1