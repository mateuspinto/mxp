`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 53104)
`protect data_block
4r+u2+4iHQ4ph9hKpJJtgkgnMCGX+vyBE8b3HswnDRvS9u6IRZN4AR8+htTDAtP5wqU40G23IVEE
VJ5yY5iD3jfJ8xMqBQy8d7DBRD8ViGxx/cIPbpf0zxXU1/zmb0bdV8WegU4/9e1Z4FQYTsYkC7II
vNX4TinKlv19rtTnh/j23I5Fd1iW0iQvPLRpiTgw32zS4EiDGrl+A+9evIqufCiq6dUtI4dDZKSa
qeeB9RtfzwMCyh2NqMG/sRRRrOQ72CVznDJX7z8+dDBqcF+/i++0QVdrRaDqgPQFZhhyLVqwMmbu
XxJtgrGOOjIkIhWChGkGtGTQmxPD5IpauGDzx9ov+PWWzQYWHuNF5vSJGqyHaq/CooNDbBvx5JJy
i/Gi1WmajLRTefY1AMR0m2soJHRgkfG4JaHHl9nchoN4RJGYTi9eD7TZct443j8v3Jdbl4tQV1rq
TiPTecwcoFbXrWQlyTpQqGA661SFyZuFaaWcCL9kiKWIu9E0OpeatJa2g7s5MOuVXp1k8xYfrLFw
q2f1TkqIBMg9JSUSESUBhEIduTzIzbhgA6//vxBKDRI+qBoHVfrTehhGO1CHxejRm+dLl0u89dtY
kPRn9DcEvh6w+9YKwyEKcMwmZmLRBJa8H8rtEwU9SQQzwWm0BKPXfHQgY5LmCrwZui/AXS6dXVe8
/diMSwqM3WY5ySPbJX+Yl7Wd2gvVUwrZdVPbgHCR/rYGdNHHGNBJov/xC7yVrGDGp/oeMXYVJuFm
9FXq0eaEgrwQPQTtXoH8IcVSlKRrHp294/Wbt4U/Vs28DbnqBQ7O6Tiib2HVzgQEC7pZxrVcAc/2
0IUdv3iSOpAgbOmY95fnrw7JvAx8nZag9z48nBnyOPgblru3iG4isWcCXap7NNgSixJWD/2doT+F
LRQ+iZqb8w3PX11+IOeba+P1OJYZtgPfPyjTD3++wIJ/qTbajUfc5Q9NzQpS+N7teuih0gy38nN3
3AT3fbIxX4SwmWmphACGF0KSMus2mVqj/Vc99MeHiAS5OrNNS/1xNnpXaYLYlFyw1QgeGCyw+Elo
GsxiXRnM+gCqJuBWiOyb8SLKsd9J8K/XiXMMd+s/vVllzrF9KF4XXJPymQ7CPgwo55voG50FIHQz
7w8tOlbyNeuIVS3U7IsuJ2wwVbY9VGdgv9zkofY8fDu6IzM31zXxdmSyOdiUCOmHHv6oci3rUd+H
GRj4cyFozDTIug2sYsJiHFAvfJnauKpN8LG+qLJqib5fvPe0QcbOw3LZD/Vyqgs4AhhyZMyWrdFM
CKUzSwyta1OCc284QZ68gzPx45jPpq0ElEQm7tMwV4djoT2wWsnzNMxR8eAnKwh4bEWvOYNwpS8p
Ddhaml0ub6URIB6DXl0abrx4MUjgEBvFHJi6wxm5UBgS5xmZJTUr+rw77FSrRNqAN9RH4LBmgvUM
yXwVjIsTD1xE/ow+y11gWJG8dip3xv3V6vN7N7tQA6DMMsicb5IA762p+Z2utBcNLE3jDsaD/KDT
l7s2bMdlXnETRIuXmpx+O7TGY8HzJ5HiSem8+HDw5qyO18Tl+ofG9okXFB/2Ne6gHYPx9nUp5TWl
nMJlmHVNdAreuFUkauNdlFImQ5VOW9OBpS5sTekHlztwqd67nKtSsUkGsrl206NXm3fTeypDJSNE
eO58tfAEn6XU86RkL0qBJqz28DjFtnPIhonSwNJPTmdKqophdUGvPwCAGldaCUJuTwzKBESvsg7t
Jjhk6NggclXUqrBllLQVN+pBrqufAxGoQly2+WhzrCXQAC0gwz5NPoI0FnNOKRu3UQdhwzaLkFPX
axLnCDFSt/y07A20q85yqIfR1FPyHQL/FmmIneIge/nyDFnlntkVJMM2pT+GAQj/BwYHPfUsAopN
Anfnbe0MThlwQilJGJyJU9912Zb2twAdhp19KSr8XNrA+hf1yC3hvnk5v5Pxrp0/ryP6d9hg1XH1
xPUOs41nEuGpjfr9HIQm9HHH0F3aVZ299LV/b94XY64+isc+4oqPd+7oLIf3MwDyp6L4aUi4e1io
0ttJfbwO6Dp1owBYrW83aNejM8CzBAeAe7q6Q6PCG253ZkaNCIl827PzlmC4S6/e/7cslUdsVXaZ
bPyPrkkrL2gtASyiXMCUNCZU3NoNS7D7bilMj328b3ux7+aGeF2Bu19y1DAGsLsouyssvmoS/WPg
hjgFBhqQrfrL4pcNQ/UpO4Bw1u2z0MR4aaZQ+L9SjqjOlMYz5N0s0B4EbMtizkB7maoxJ768k+hS
H3Eb6t4i6U/gIfA1bJuoU6QiOyF7qjNrLkQ7KLF/6hmVuo7HHmcKt9rR8oIDfPU9UTVipCj5aSN5
Np7gWLZmUbQY0dBuGQiEF5QXBALRIs++0AmMxlmPiB6muLQEgTejFIAG9pIW9iN0xS9lCXbMLCKE
dPO2domS8JxuzpMNxuLvAunfhl5sQ+jS5jnx2rQ2DlUPCPUq3/roMsiWDoySHUdzEjPbCPujpJBp
Na7QZ0VZif/IiMBlBFFxiekUSRUGBf1BrhkFiGRMYzsU1QDI/YRqoORzeSP2U39coXqo+z9uA5no
3mB1MnmXmWbLkrppir4ScKM4JKALeS3TREG8sLc7ZTUyJ/zQM3iM3McVzwsJF+W73rDV8GFeHW6k
wZaARaWPT3qydmokJz+dS0y2i5ooQ7zaBO3hPfR2TNkUKS4/oWMKv8WsSjz/l5R2coKltgWSqKLb
zbUGRMSyvR+YUPtBM4olmZVG1fKmyZCUL2TO5X+Ie4AJl4wCORoAfdLcY2+PX9+HmDI4b7jtJZrv
Mk3fmLdGVPuy4A9Z7EXWjmyFeIte0e8NsAehl1DXy7V9zBmbSAGhDnfENEQANfVK464UbEo4JXcq
fd613ZOnR5Ilcnas4+ZvILFl6zsRzrKiaVRQf95sciYr1MIhTiGpCaG88IC1PJRlYoHpO3d4vHpc
7a1qTdEM70NRyOyDK6onJx8tU3+a4gELXh7CFHhTASZJGLdMYTtuyFV/R2dvdFXrwZ5bQwTGMnR0
mw3nP1NYCPZZZR5v3sn0VWd488LkYug6FOYw3in7q7rJCeYaOoTwhBedV7v+hEMY1xuKTDe9R3Hi
0MO33GQAL2RHtsUiBDKyVNx2HXvtSo3OWCLxVT37bZueg4BRBHZOVRFFJrPJYbtc8xfeXG6CyS6R
xLodL1wCXe3Z8fwudAkOQ4DrkHOH2vMMlacV6+8qY/eI470Pl8BdFGhx0omVEIDmoywxkFBdt9CT
kDA2qCjANltbr/nT1flSyLKOvrgY5VRpWifCNhZQoSfc02Ln+s4mAeHa0UAL1oEH41DbcG4zPlgR
NgOIfLlOrc95WRaXnVEnhtIdmCl71YkkLqE+NSUhF67LyyBxs/sXwzFeROdvAiqrMV3+qDWDgKkK
Tseu0kf/nmEHbvQV4rZ5a6OkD8Zde4QsyVR2Qwdp3kKj8oonY/7jS/Wqh7ctD5SrFVV7pfVkFXVg
gE/Kh1axaYihYjon2Zy+M6rZDErDg02Y8DhuIjrrqEUYOf9GcCpT0LcDzivOAdH4PHmVM1FoXSk4
Sxbv14XZk5Y3AeVux2rqeNbTSqCM6/Y2XE7AsFZo5/KRX77EgRgzvHZczEK8FSwoHVh7ei1iBwPS
A2/3gU7hKS2ahgg8LyptmhkW6a+E7J48Br1XDwS5cvo0lVslj9Y5434meoVhYiRtX+MfqOzlA3jy
rF3ND0f+WtqUL6ejS9yh9k19u+OuEEaWTaz2d6cQ2z6OGoCl6Y1zlqMqH4UQ+f2dL9C/Jq33Q8Og
6WyoLGG7GhqkFek8TpQ561WYAzmys/0fMQHHja3aYSV6rXkSct107ht3u3vENeCUASfYNqk2wHL/
mSbSHVMFfKRjlV5RXCD2GP2W+Y6nRwdu28A9hEmh0CjkeOOLpGbIlhe+zRK2P9QhNt1FwTZ891EO
X+H7QO7bVoFcVwUkgFZfWBKDEq8aAMqbRMbGr2sRbMEAzEkOn0yQQS2EmycpIPchH05aQNq/CZ5D
cRwyDPjoSlpjepuj+NJRD2lNbAv/Z8wg9AfGYaBslR3QilO6KsIUW6l+vnVZAqpmak4dnyIOdyd0
mv1w03bbVHhYxwZLnRE3PE4P7XK6j3YiTqr7hwHhkmHXy8IyKwHpfYx0OpaDlVRG+5KGv80pmyOW
pAysFi5/Hgj6dbksdiuCfNVZNFdFMGiZO3fBc4SxVvM/PRjkSTF10rK5LecZFGV4q/75cia+0tgT
/ucvz0OKzR/CAiuQTemufe8a3oYNTX29a8ZcmGpAqYt3kDe9LMieEQOqX7cB+ZM/AvgxezlCHJy0
mUgSlBrub9Gmk3MAk4XvyUBPKs/cTbKxCclZ/m2iOjXpUHiI0xxiSNOATM48gIXjxYe5mya4nAJD
rHib/VQ9QoWqaRq77EffaKK4K6aJlqjQF77Qpg1+xpV/7Px315kTRtrONyLuai+K8/cMfrpCU+lS
ZI4EbOYO9xxJI3phpkF5YGm6isAMZMd8yG1VpwZ3R9lEP1BFCt78IIqFyw3Nk7e60a9ey4wn13x0
02hQV4XyXB0uVoQeqdkMU1ILnlPM4wkRDZ6M7ZFfJU7wzxREXx2bqhyFvv6+raubhcrBf3vlo2Rl
+TNugJzxRb2CS345m8W53OuzddG8JWCHlei3Zk0a5GNrSAhiCzpJTXClqvAvw/jpj+Fe+YuQAT7f
I7A/u62n6jBEoha78+MT3elax8tY0CnYOZCxL/MYK3M28A25pBt9NCZ6x1F01efjQanwCNuMD0Dp
ZXXYf7IGVAal0QITcJmNqMQ+ZmjrCLtnr7ZidsRuv/vuyPl7fYtZbuOW7iUkohACEMPRbm8ne8zi
rewtyrepc2PLDR38mpTw4OSqdkjw8ken0BXJwMNYv4f0qZB3zcsLLOrCO8/dPSgscE3+YMtGjC0X
+zmmPB+dEnFfGjPBzrlYJXL3Yl0Izpkas/UZ4lguw0TeY7UqYayRnqaKIbFu8YVe+GffDu11CTJD
levlGVHekHGGUuOr2G6YRoPzKjBrdKid3+6lGIEYR7Jhrn4btscULiEPbAgGe/40CXQsklnhukwj
tRzUNXB2QJ1ERD4ypCLa1uTYsOxkqMGo3zYzNEGSlQUqRMRNhMzIPXpOeno6oqfl/ezdwxd1K5e+
5qK1ZbcxFnOIOm5QBmX9+GaIpqVXxjv70E6eqxa9V1Ik3h7oHuNCAip/L03pri3vVNcjTbmaF50F
MI+pt+bEmw77rylJSKbKnG3znbopah8+NNRc+G+BHdh6L1KJ/VKwS59u+kgxdzap5hsKspgBFutu
j4RJtsNtrHf4S8mu0K26UhW40fccILQ2orB8Vl0578Pz5saIzSbhmd+RsI9XKbx9kGjGGEHpvcXt
1wlIyIiihQk+iuCQ3mh/DcBf4r0IYWiOg7U5XLYJ1OWynR+dfP3sGqi++QN0wleEIej6M3MVDSm/
bzOopySfN+z6mGCbIH87lDWtdkyb7QhYdCFhDMI7M5eAqM39us7zpko2q4HE3v6kDTjvFDW47wG5
L8pRKnlm0wYvkBtkaAJiTpVZduDvo8nHNfYgdvb8w6oPYVhzr4aHwphAxVMKeEVg47iovJ3WwGeW
Ninlymd2+b/vtRYV6ayGT2TDxLjUfhU/ysEyW1q+DyJlWKGo5OnOCUjoTRE0qPXYthj70A16sf8B
iISwIOuTdp4DE8gBVoXhxSv2/I6TGQYrhuAnRxaoajo9eQdQwKZ552MvcexhOeI13vYeFol8XozM
+BoeeW+lm4i5bwBHspoimobA5BfvqTisBE4iHOHP69Y8Ty9zLGZjr40gN0JUVZV2c4qdqXvk+yb8
chS6Z4IInzyJaUKxDmXIYXfZAGEPGR51SHy1CayBwbCEd0m/GfVQEIRgUe8viROQXYZqySQgUz0F
TXaYKfnFbNTBz/2dsiGXE5uYYbu4Ann64vtV73C6Ne+5bRxCpE6cJoj3t3SjSLRjQIjLRfIynn3i
Z88prpfeDa5zO+p7ku795fYUGedzNB2jqn4TTelSu08YgwWMIqDTsuljcIVpd8HdofwMdZLOTGrX
WnwNmi9QcDfP+JPwpVo4gPlC+pQme6WwrhJnfnwEpxCFuJX+MXuWf0m4sN/+4eTz32hRHsYpRVTl
I1c3Q/WOtg871Go3urwuzrPaY3sKo+ZfwLNYMbl6UvVuNgfWPH5RPnGlM8G7BKxhTHUALLWbp1q0
g62T4HIJ0VWxGnHydIiccSc7ketO6OYdqm7GsOSfuHMNPPFe6SR/QGOGAAxjd9gJb8fEG+OIWbs4
UMPGtJvwlRCO+D0dg6I1AaiROekz23lr/JuYjzUW3jKvFynRP5BJG/EhNvqloGsK4LKk++M8L2FA
9OTl9k+HGVxOTdqNOvnhawt7xWqT3onVXMLaE1oF5vZThPRBkhIJhsxI+gmYc1H60VfI4WyXZB+Y
FitcxuSxS9M27TS+zLBNN+GjmrfjIIDLKi9b+ai/Oox31fwA93jlcQq7gEsc3gNTR49foERS06q6
QqWBciaRB8Vs114+9RgM3ADiTB2AnLliJN5J8mjZrTBFyvQB3DEbsfzGfCMyFaUGwV7dHfhwbxD1
KhL0SVNFya+fo7WjXrSiVmPIRaO7pSha7FE2bq6k9uoiT9Iw1BzrlS8CW+QjNSNuZ/WyVk7v5vq/
zvVKgYigZBKDBmldBI48jSHaeISUQYUFH47kbHJmdAiS+YZytW0Ab7+/t/bmV4ufXJS8VDGYC1fa
YsmYrWleb5fJb1VenSvHOg/HuRRIPfMbb4hcNXuB4Slwqn8R78wuXySO02yR72o/hxcScDVYL2v5
cSOwD8mQhyMHviHXGXbqsVAw71ESGEby36cJDWX+RU/jDjPUqFKqAvof8X8GUlbGllqTMSZO5qEm
kz91GWsxExkYm9IX99bgZPMb0WXZszMT8c7MJSyTMwgXlfEMauVTMblPk1wL+SPznwkcS9EJwUCr
ElwUxftf03epqC7qjANrzEv6bOszY3IfTi5sJ468Tbj249WMdOU7NrzPOoDHjXx0IZuC4s66wDc4
fVzEhfmDYwew2akpx7GpUifvP0hCHQlIbhz5+cijGZdOinJse322pCxNdxeobUuXhOr4D8HKg+Sm
6Ozi6Ihcro7ydOc2BJYEiDLmZWyWSRpGDAvPw/DAsLevnNYP/58uINbY6uNZP1jzmLTcocWkzIrg
FTqEdsT1g2sLS6o29zF1l7C2W4Aup8/NJAm7TGyIMdkTH2Ada6ZNqG76q4XPPpq8OhUB+WkSsxcf
talkiCA4dFNxcprYfbFeLEVMT7MB//zFFfMjun6xNqdAayugzLZUZSZ4AtQ8PYTf47ef1DOsROPs
6Ydlekj45GdhyWP3bOkbzYGu2qdd+Rq/aHqPWKHPbrOqHiJ37XbJL2OxF1pgqET1svCWNIa5HZUO
dWFkDyAxST0qArGHMtbV7Kab6xSbJV4pijh/kLkDnENgdE56UVhcq9lJ8ACRZKVhyoyoTEU2SMyK
IbYazNI7J+1D2Ldk6kF+AEJN2iAwvaRkiP8Poyd7P7OGt2BZUDs1dDxBvZ+so0nqPImIJQ9U3Raw
WoichpWd/yozx1Ygawrb1v9pr4JzOnTaaHzCxfInYHdAmg2WEZeND2pz5Z8NY/4e4ZsHCXFFzpFP
NOhgDcGmdiD6IHmx2bMST1SdJ5Xcs8/t3gy7ZMsie8Cr7pREc/R1siMrevLMM4ntgVyn4MOXarIr
TvL+FmQpQo1BIPEjFIzc+ZCI5oMqw1jSJHCKt4O23zqFjfNwiVOdLKIFTBBdG5XGDpsrLwSbC/lr
X5auu//B8ZPevEriEVGSfmX0qsKxhauuAojvsPT6vokBf/Nh7/EmouLFwKwGzt1g2n5swfD+m6n0
MneWfvPUPWI5+QlnOPkplYlUZxmIaeY9gw//hQsF1VkQY797s/492nw0SHfDmDDbMIWRLJoImfZM
6nq19RkLFDtMgY7D1Jjj4YHLV3FC86aufWIpnOeauNWcSCHkUSMJLlEqYZxyTiB/OmTNTHU1NVrK
ywO7VjzuTzQ8Kh+CqMU6IPK6XC4e4XQACWPTGNETGSiG6ZCIh4Z4SsaOZTSBgbygQQ3vD1sZVOEG
rozc0oOSzEPTNqB1tkE1DXrAin1ZyBP1rC05p/uYuZL9R6vnRTw8FDQ5p3bKPmh0yXJkOWOlb9jx
OK8t4Wx5Sdh9q0TYDVHR+omSsXfKgVyKZqFh50yWdM86IWESRB/H07suUy5kYrHHNCrogS6wiJ44
SBc5xo9oerj2Gb88N/9vKFTun7VFJ7uCzIikRgwiyYUe1dxWG6ZyCVG8N8kKDV80Rey2vcT7NrfC
CVFfWrS4en2VyRXJ6r4AOzKvIPbh2z/oPmwVtViFExDXTvVLYTLKWZrRqqigcPGZMi2I5dQaR8wj
jjd77TcevktB4Il//LAa5PqJXMnU3MMHlfIGRKbnLeCkpBF3bs9PAQmpspqw/P0qMnHnGQcTaluz
qDwXIGBDBV1cEvEzqhbDyBiG/CmPqpf+gNNJ0piyJNeg62t1d7Tc/bwUiFXctFFn7l1Pd3reNJ16
4K7WeJQuuLdeeObMG6xCLjtyPiMnLbakTa16U+vWCTR3+zpOzCDRCqva1//o/weV1vlG6m+iQq5c
/njjSVODOIKTzWG99gGpSp+CjY5L+yuRcyFEeSyCVNnqvQ1Rql8pepaCesNSqUJP1Mb0x+LcbCpx
6qwi9+zYuBFGfdq2jeupVCtis+mvw7pTwGtjQwFCOXijccfU6duvghqU2Et/BmHPdleZWR0McV8Y
lU6IWGbR2AdjyVH8ogebCWr+V8W0GjyBgPlJxsyBYtNHPwrVdPj8XdOtkSeFxiuWajY1SHLcDjpf
H6QI+I8y2eVZ2W4J0Kd6CeMbc+HsxCc+8pj/MElSLMsWehq322qzhJ3sUS5/kRMJOICUX1PuU3qn
JTStvibhx8MdxB/GSAOhW46JAFL1EiOUmyrPv0/ZIo0d6v4FHj5jj0UQ771lUyLLmIUVuePrulRd
UUBRaSoWfglc6EZzdZtlT+Jm0g4hL0RKoF41lGXuGLupsB1pg5yWaIdK87bTtTTWC4tcTeYauxby
gBLWXFYC7hzNQeVBg0f+9yq/NSqVJQq0jjrTmjPFjEodDk0hkyybWVN5zBNkIZMMiEp4YmWCoTkc
wvOl7WlV9+15NSkxI18UZtQvb6mpjxd1EfXQDe/AjNNQLq5JCPSh9BYaIBrBd2euEPCMFmxCrhLA
YUDI/7E3L+QEWiM8/NvPgT22yQWkUbS5DH09k8HXtiRBfhlJnt5uNcGbrgUBmE2mRVY7NvJAMKBn
MrLEGB6MCYYp8tQXoSZkNUTBlOLmbPDKjPV+2HkDk+o82eonivfnSWI0Q9938m75gV8LEVayQlGA
VZ/hlIYQsJBa8pU1CElKlrUdjsL342hm8Ubmhxg6rl9ahXhvZ8c+GPDB86/1TdKNzBW3rhpug2hc
V0jTLd8jzKy7Io4M8bZDTNg6jJjiLEoQC63SWRn1es9jPtmwcUS631foq1UtALp1lWFuz9Pl4Pe9
GmWIvNVQorXnUpXbN8hkDFypX3eXYPcFiWwuDegHd+qsFYXK5Wa38tQW00iAYx/vCO5HXKJ2uGCi
uEbamCKZl9WsSm9+RhebBzPVqjG29f73EVlyKROkA0Q0BXnIgqC7nq8Z/ufmWzIY4piP78qF5Zv1
3u4S2fZgO3UgRc3thDG1MCGcLSbFFdQobXZ6l9lzuGb5am0/IG+on+vGuoyarzL5uiTb2F4Tu39e
CNGL8HQHvLAPDVmBm0Pvw51s19826ha90CZLRHxJA4JVNuxAiafy2fetsL9Rp3s8M0HgqblskPBz
kteeJERCyJk84ZSQ6R8iYiYPl63RQbQUCe2DfR+rFXhG0HuuBhW5ezAhjfp5ejSSBDO+MCobvBgU
B/afeSqKDG0m8EJOWuSxkAGTL1C2BjyIbBpa4pdLSB/a5QGp5yFDJW/a0J+cW4Ge+O5hzqx3GWYr
w/LOS7cogJ9pwpB/wLCFmnOtZZGGhy0zUC38LhNHyj8gQQkZL002l3KqD3lkoUuQxi2PaVMnfXP1
odBAxdMPcyxLevXPcjQuxdICL+AqPs1fwpG8ahIRVlOFt4hY5CVVt4tTuyr2fTIvI7U1Aa2YB14b
fJ+jCYVEju6CUoTd7G7C6w6SuLSJRobUlivo9H9EZtasdYme3crROSc5y4UiQK/cYqvPvnWrHv9n
Soc0jlUufZcEVXSijNJWnZO4053Nbd/8C9rPUVVkDIm8iRqWzXnzNBJH0g51QcslIN1xm/EekL6S
zOK+8yfWb9LG2fIX73+EXdk7a6qzOxaBRcC8K0+U6YsRGDAexFCDrJ1+HjI7F6aQx3WWsSEwkBDh
00KGJckbOmB4jVR2tXALYLDQyFIPz9f6xYk+3ZoHmh69fb3UANyARe/A1W5Y7Uahjfu2FkFByRJJ
1jYB4Maf260bMb3XPHKhQQo+qt/qxcfesU0FJ3UP72/lp/UQTwNcp+VMvLRBJyCeCUUBybGuBkXJ
AJ1ZxeIAgUkkuRGZzAip3A7ANHQ4+1vDlfqK7iAMv8HGe5wPkqYc0bfRHNl0gjg2Tdl22TiuqJAG
otoRf0yaxAqoSoDPU/E9VUknFM3P7oHVF9B0bv9V0xEVb/rrerKnN06lC9aLDgZHocwJWONIvXTM
ap9My4oI49ceKtrxAflkBlceVEq3B4VQrj4nDNhN7jmvua46yHtDrmxcc2vUaGeMwmr8U6BzOxVu
k7X38GjQdOETy4H84+KFVNdRjj2DQsGdFZuDMPiV5jz66eepWqR8+plY9ghftDL070yanWADEEKN
2jxP2dz5DE2ujnmy7OtrAIgrtnX0TPdsdlljYuHUv4WTO6TzGMyZMWoVkSJ7mvb1/IVK5paE8ib+
3+jUw2HOZwdEw+U5L4iwt3qYEVeyLPwZJ/lPWormzLOVfddEHEFYIpuOC/LkEhjzB8YqKFaI9JtW
j4mYFmYppWAgWpyIUXrX7xJhm2dXJ/iU2nPvs9DYe/BhRjcLYdTK2l7pY0r2eGyk4ksBRNK1ej4+
vQFnph+ZLZDepPpV2ftx+DXcKdrHBqZhCcIgRnPKF7XIs+sRYXImx2mzY+AYj7N9LHGxrc6fn0eA
2+OuGgxIBaojC6RDGZA3enwDqeMAv56TT5UTfllBYiy9lz0SlB/HQVcLODac3c2FX6Cmh5dS8z2r
it0I2Nx9XXm1prBStH6emmmVx4ZMqgtgDUx5aPkKIpLZhnkZSjUl1N9xYl93QKsB0pq7w/M3MSUQ
AlO8kzjnm4ZZdqj5L7PUBOLIdXHkZUbrMLebI59l8oPdLyVti6UYY5u0Gkgxmvq29eBgQv53tk/M
TBWa+iGvZzd/0q3JV4kCN6xAltzQg7lXSjovFOnLooDfugHgvOoOCTByy05z7IsejXetO6Arc/ji
ur7zAGiYK/noW4b6cRaebctlurfKoNWi9taHjmN3feEeub48a4+7bLGOmDuXbNE3KOs/PXFqNT6W
xhkcN2s58nN0L2Lhoa8VZBFXgQlyhqp0pJ/wDdLXGqUPG0jOFksTtQzf4CEoW+2jGxhuK75Y2Vga
wpLXMcaRx3M6dBMt+04eP2djcUjL82K83CynPL7tzNTtRDto7vFzbLzSgbfXvttw37ujE0an1A/W
fpw1NFCHaXU6Vc/fWT8pf5CEBqZw2QhQVQpZ9Ld8mQzj4nEIB/OqTXr2EZbMpGcKveRnUZQa+qgL
c2+BaIBIiC4bVIvPQr00/ZVuVJJPTpmBgu4ZAd5cJFk2frr1AqSz6/llmgNDvjg4GVZa+eGPnS/x
rFdnuz4yw08WDjP7zIb4uARL9gGKT/b2YDZPhKP1PGQPHd98E2UZhZ2NmVKqrT5haXospmsbxaqL
W6oV3nyfc0LZVP7oQpN21GU+Fx3gh0j+O5mdVOINh2nB2IF0iitFFk45UBm/1WeIe8ITHbP/UJJQ
Lo4RUQwhCcVvcMehR7Hy0vRNUUTmWXjcRKrC3g0T+4iHzh4fLppoxILrK0bSNa31TjQ3auILs/Q3
6yGRcnY9oBeXhCEOeEaCaM2YtQl8a6CzbPzeNtzFJev/V7lRwxRooYeIRdry1Pfyxezg0LADbFCe
/5D/yQladisBRi6zhzPYYYDzLCb2ZIUHOz3VpyzU43kYyi35L5BmyDRJWvHJAwwywOTh8HTTwkJi
/0lqDBZG1hF0wxx+UVrs2pTGcSSaUkfjA3upbcqacEr5+ayeHbwIWg5Xrm0jm3R75B7h4KSXYqtB
5C2X3QImkctlNH3sjbDnZY83ebG/Rhz9a0ryx9O1N28vxDFnlZYvhZmpdD0YOTx0vYxWLYAImUHp
o40mxcI/PRjQt04ypzY9w+vmE3qgMFLoiv33q+P/Dk2bm0PJQxTuRG1wln2MgkDHlu6YCmfln1OY
oG8ctOl+ooAiQrtyaC4OBZW7j8ukXGn5fuorxhSSoFGxWy045BJyYqTQl6gau1ems+0GMnFXK8sI
5ArgHe7mp8YpsqcY58+uy2bb+LAySAQndLGJmKRp2vGHeBlVfgUH/JzO04rQOwYuZaZxbjJg/eff
M6dxDpxlMkTPNZhzQ87PIyIHRm09gSLCdWoyuYJd32tKu3tShqaUwA2SIX4TEZ2lBud6gNu5bsjq
vUSAPw44l9SVEkzG/eKeHc2X53sPKLLSEJuZDyaoFiaac+wV8Zaj0W5OQJY1ZlThhAFQkEg07WGE
DX1ORfX3GvSmNs+EEV+NmOVk3Qf1XZf+fh5e3xKebDFky+hwMEyzMwqu391jAcKB0oOnF4XMYZ//
VV1W+RalZY2ZgWAyMhHFjyZZdZqOT1KGipWWwgT6qGCufcMl56WacGpCpRb9qvqCG/okq6+rSEhc
5hkDD6owNNlpfoBQBXH0jTqr+TqTsZBjd2bedRl9FvBLA6LSe9ED9RVDM6Vt8G4ylSdsJFIHYRID
ITtDHTG6C04VT1vX26YTw47oXkBp0Nq2G0WoQebonSrpaRZoGzn4fmMPojDMm2qXafJui0vsvCjS
GXUcqcXVBSJIrFPiY51iVNiAzHLXSefj6uLhWOP+NGgYBfl7SV4N6rUQ0TPJgbxoJwFeWXT9yrEr
sq/iXgNMNXYtGdqHhMAb/+vYau+tYKak7G//QquQh7lyEPMPJ3Ee+4BUHZxXQkq2gvVi9K2qz/zQ
eLUkU9o19e7cjhOyPxr2oImtm099qz67oYd2UXv9tG5yDRPXK/SxPNdPQCXj20hKPVzMWcu/iAM0
MarUksKva4Ma6njSh5gisuK20x6+uys3EL38foapM5HJRa+L8MsTNLKMsewt+Xyau4impSX61BsF
xCu2nq6QP1se1o9Wjux7R3wSdtTX/r6m6UwMvw4CgGGUi51xCkf5zGhP/VlBWdXB+JTs8vMoyrMK
90iMUv/wIja5JMU3Vng/7EQ0jrZ2FSM8M4GMH829C5bN+W9ELgc322xPOT/hI7pYo5QL8T5CRbkO
NWNaOJs2/k5KGSILe/jY7qiUtwutWb7fztJlwwDT8Ov79D3KzfpLym8EPbQx/nMukyne+T9rHlF+
y9qydO6FuzVti2NEhtsiB7ii0iOgAOmEIkOWI+pOq7qpUNqihu8WTtcLq/RbPyBCK4VBEZceDf+8
vg6ashLyUvwDFG80Lta/VyUeTYo9W8z4ug2RPB5CzQ5nLhlMGJcEu8ImiNoX7OqKs03JOMhh6h0r
AMnHwj5b+iLBAhBOgdB1tEqkciq2o5lnmlX8abO1NJROdktDcgmWwoZaOqpwwzfxQUuT0j7VKc7J
PJySPGhhC1NgGlc/fXqCTOTZScZfdeb7O8rlKXWYx6IdfKuDyM1AhbXAN1YWASboOR1kOzQF2PUh
39yJbVtoHUoO9NOvwC1VK3iAcHWJdLHAoh859+MtmTCL4q0tpIPICNGQlWOOlOGgmVWOF/bQvsb4
vI73HFM2knc2zyl1d0+rwnptiwi2SRJzgADNJNGeSKX3IJDCoTQBmmZ7oEPw1w+au6lKDIi57mLp
iISOA5ymy5MdxcKuJ/VOcmQN1vaNzMz1c+/n3FM2TKH+NiN9pnsjmkxjNGTG7UoYK68pIt1A5Dli
6r4z3JV/zRjmVzL05W1KtChhWpSqPj9CELR25ckTTnqK8n2iD2bJ9v8Gg9cSet8U+uBBXhF7NOSo
VRUwyFTJiqg9wNIYscP/AZWQWedevgIkTx4vBn2LkB4+AzHH0UgW/XBL9RRJGZbbCmFavOCRne8s
pKqklLz5OQk9YBKkJNv5eBpSSsYuwWlrfjqhVCyktJAg8tTxivuDTSTnImDrJoXRFUoJ6uPxG6tn
yIcdFikSnuIwVx0P1QHnx4QU8OQzkamsYTuGs9VjQBtcCGpHlkD4A8y7i7OfVr88P/6aUx2ePSUB
wKnitHVKvxLrwMjRjw1IlaPOMtkrCj/eUmTr1qWmcD2/aAGR8L4cmw0NMnnm1GRN5DSZlpxsCnAk
WHvBSoaVW3F/BsZI74yDnNT/I1Cvrer9sUEq8ZYgy5MQ75FxntUjY2uinKt4qAh7duxta5ANvgrK
nKQCpgsdg81CoT8D+0wJuEewmaHhxykSnn+cb1Exap5OU2O2xvq4Jdb5FC8iJ5dcGxCWw9NbcWm7
ooNC1dDM7zOBhpb3Ulb1ulesFAojnbH1hA3sPGIDQivuh6kVpokixZkDz/1WtGa85YdcyLvS5H/i
ger0866Czu3hqPG5lqpwwr5EZ8DMQKE/pBnfEv4IaWsexZmjvCccIwX3E3F68arlPvEXkQFWfCHO
9xb6RQI/PlXuejZyYP/cy4MzLIooFYpg13fe94Fr44COHIW0Hma1nwbS6+PduVF+qf8dFU+4EoDh
aZxeujEiJWIQ/ZmqYMQYJdom5Y+HaZAJzANG91tiIjuaIzGbUiH4eRVlMIrfSDyNClrRvoB4atYJ
lYvdglipQORdHBY7hEcc+lovSr6xw8pDXFxEMVK7swczpIY3DY5BBoZbbbINgLARS5TvQIJzpxVE
V8EZsjmKVw0ea5fnq0b/eEvIRGljWYQLZaOdkCocuety1sC9YOi4QF1ADbcNrBrLkVFgAxR15sEg
x7W5ziEDmvjcbc4Q/iHD+qit5+oeoDohykpNclZL0Qd3dUnJMejpJWcZ2MX6aneF+bJ6LAc0xP6H
WVALMtouiDFYzqvrftXiswoBcqonZR7lC8uHaYaemeC74MNDYLxJd2Ff+ZKVxrskOah53pmGQxw0
HB0CA49XVeZ44eqDVJdmhudImsDBFdHcvPdE2lezxOhIqYBlWJxpXMBkhg3qSX0rU0OqXQApH/fW
irzocWTwyBgJtQqrMuvWUhE8/YSqkEWIu7ViTyrRYS9YiHKcXbei70sC/zMOxTHDE0aQMcuyLp5K
T1SnJK9gXuG7WPLoRumXkauuq++/LBo4Tx8p/v98IRs99h86klw2iioLHBvuiS589O6YqpbZbBAp
/LHrkIziePNRSL6NRUwYTXPO8Sl8RsScsIFHmMQyGcemPdi5e9elPX/y2+DSMIpu8qXNGKRRY3k/
LpHUYT5I0z2j/TjpTe9Skw+elKQLaYoJYSrLc4w6U65B1Qj0zpzbdMWXJbBkWnyt1mXqFvIrggyT
LrG3MWcxvbIZdzeepalCNPt2oDOyNP9dfxhKA6cBLbDhTa4yiX9pHXDlHScf4L/PfE2dBxYOevLW
UaRZ1XyuGniRPx+SLRas1k0aaKvM+wGo/7S7mcpbkRCGP9iBrYT8Zj1lDsh6Bu/VGDPJ+cQ1hGkm
+nL5of7VPJerNdBl6KOk+C2J89z2QWkK7eMQlPOsZnEleuir6SguWgtPEZTWQxTYHoR/xZL6dXlJ
/rDD8LT9rTSwSGKW63hmem2Z1h3s5TyjhqMcwi/i7yc3y9ifVa0wS5PKNgbgWFFiMxKFdpdJ4OO/
To1ds+OaY9Gv2CO122TCgySpVojFd9fCcOlW/npb8cyKpytMqqbfVFZ05Gtg5k8Q/u0xT/O3CEDS
63Wu7DLTRVaSLJh0KhVj8VlPrvqLFsR3ov7kzqkB0r0R8I/StF9/hgUe33W+8GS2rzLuS7fI9FWA
xw7zXn+gR32ShhQsM/3UzhU4YPi7zw9S5P6XFCW2mlfVpceYly9sITc8W7GQ6xsFFayAujvabz4G
jT4ndC0ZRG/KXnrHLsslBQEvA1EDQEc0Y+0aokp3q9GWzzAQqghFYETO/SWW+xFig4wU2KUdA1eW
tgl7CfrWbF4DImFIEGI/Sz0VD6FK54hs0pXB10tvMRYJHnlCMDGGEda1MaFclTYQLBzm3v8DwPsD
4JUu9NAZ41RxjjZ/Al1c40D3qATtAIX5zmtOS3zL6EdCQrQNK1H8SzAyUIKNQQ6kV1VE6XKH+kbC
7h7ihQhLJzGFYnEJUa2fH2UCBm2omkU7CTLxz75/MQ3ybo1CpbJHr0KYGbh3cZvvu9C1Hxt8bRaw
OA1I6P3DjaboTJjFTuCdPWRhph1cPovJVrPTdVhZbg6Pwp3FIM9GO6hfSTlubKk8omgnsoRRKZkF
ZFvuqDM1V4/C1+xJQ4YMVgG+lh6RNYkwAalln/YwW64qlWTuZhlzrQ21L1rAeix3pzT0iUYLg7af
KHGEIw4em1zUDWtaIqj4TEMgD3hE91COQ8M6rMjq4dVJ0jGAFgIizgkEZigXnbsGjHzCwYa36UJ7
PMvbzv5rP6z/RMQKnSDspETrhARx0QT+0J7R0ZvFbNrV9EzJHidikc/JqnBAbhrJeCJGrhHvmCZk
RtoecIRVVDfxa7Oc2NTy7YDlUlCAEBpsRjrGWA9flEUm4Z763ZvgTJ0hTNxXIITVmPNBUcVTa4wa
rWAZLpWGQw2W6xQFMSfqvU474CVIJ09moUDqFVTdbbGpXIs3Nosfwj/zg9udjDCANnBkJc3ZA+3I
ETtAH4uvS0XDR0oYycal3wrQC5gInMUlZoVA7hIeglb+TfRjMqboE30ebEJ83DolxUdz2vhUxtmt
AGWH7wTMhlI4r9tBeUsoqKt5x4CBM0hQaC8M30yAa0lTPXHb/ja5vO4cdpbmjn9yaAP5k0ReC7jR
Y6JvAj0JbDGgrg52Oe61xS4zYDrP0cchmd6tg3VVW7CNtzOhXX6EwZBAON/PKxMBa8SREQm0IUhT
vaa4g1MOD47Npe99GSckzG4Irt65on+UEofseK2Ql9ESMTeTzJy+uNwgS1hdKOORuykQ3INwVEby
2dRHQWb7tGFtjHtUPMcjDYxzPb8J8IPyq7IuUzOSTZvPnfQgArSnDsO7/HyJfFyJTKFW9AyB9uI/
C2n3yuBOTVFSLG5wdDohyMQvahu1Cwwha06vwlehEufunbhOCpHBE+nzlYvbv09nzQ3Ext97kS24
V7eQ3IW28JREpQOKDVzGXMEHyHOZOczCYbyW5JCUNE7X4olCvuaWvyx8fd+dIQiwYDrda60djWPb
+lt8Ixe9qGAJIfhnNlzjx8NxO3S2BMhBTcE4czrd3yyW99orBtAgaPpop4pyVsu6okKpziVXeTpb
yRHcokXwTODX4FOT4X1s1CdOFwdmzaZ+9R5Pn49cWjU+F7UBqPh7T01V4qDWMHC+gtsm12EPGzh6
qoo1M4v+PLpfyHLOxElTrl5zGbXqT0bgKipWeq/qpCV0gxpJ/ZpU7yTFt7TRAu9rfAUtUoGnCQ+u
ZJx1RyYuczlH1uPfaDFJqBCGCXJIy+aD3xQBuLQdvYPI43Qbi9GYQRaS+a2zMF27+7JC3748ZTJs
G0/dpQ/tbFRkyq7d3kOry+49yntpOREcGqHTuyUotIvCtdwTOJFCEHUIr/1QbGRLNolEUTqpsCdT
qMoI9QkAo4TG/r413cqMMvQONoME/F55AQNTzRJAwNAeTK16n+22pAIRqjM7VDmBWh712Jlx1ptO
wamPzbzgf7l2qBhOxFyv26g4+NysN29EWWi1hIfalitc6XTOihOuCUOqsBmMMoBVhy5Oqpqyqiy6
i04pCcEQR2zOZdxhSyDwxQ2Q1PdsThEWYs7PvkdGe2EMr8KPTsNNcat5+VJZFerk9wFOCMmrhcOq
rsvEmopCaGvP+uE5IzGRDCEgYeg7xbOBeQMqKtywinOn3Igg5uGl90dx+YvFoF0fwfNH9rQA3yOc
HojhyLBdeGdJABruJ8ZN+3Frpv1n1htzJpWzEkGMNQ5NxeItZPH0FXFkiC1BYdwGAGwxjJQM+1L6
BQYZ2ve2B+MZ9elE8/RYLTMhTQblYZEKU4V36JFTUFvgxTVmayZNEjVGF1Ix9xCpGV8zhgdZS0Yh
P3BM4mQ7xWk2Xi5XUX/B0YKoWG5gl87JT5+cmhpf7yMvi2oPfFIROnO5wCEo1ivtqvZkHfwt9dg2
nqLnUBM7gGqGz5Jxmi9xNAwyF079IDIZqz+linqYk577jaY7EjEkaJ+rpkxk5ixVfAVxvu1Fe28T
zDv5GMlE3WubXrQFNdlilNmXdjjwwux73cdE+Ku9QV98sU80hvxVzTONzrvNUQ3QmQWA9AmJkfTW
HkVaf0VRN5MhkvAKUGUl0nTKbhSqV8jJ9cCyoYnMoPL6WkGr21zI0JZF/XJ71J4w687M/4+5/90C
m7FR7DEN0rMbziCFzKVn7fL9T2LW4OEZbQ0A7M6l2xgncf+MhiQCyRFUei0oZHRmWIsy2VDJwW6I
DuwCQegKXfbrlqIVtM4BgIlPEhYlUkAeriLGmwvdv5eyWLTafh2h4KD5gqe5E8Hh8mc2Q2wEy+lG
o3cXSMSP/LZ8TgtGczv0srF46wHaLIWTJDbtMr2zrjX+E47mTsNymqZEQqhj/xs94Un61SVTPL8B
HJzI4Ac7iQRKdCILNUiC/3WE9863Xbmc17nRgMaFQ3AyCX86k/epT57/0t7E6PTGhc3OC/9o7qZM
2Ss0TfYZ7rS4G7YlHZu3etKbHZanN/ZiE6b6Ro6oZj6TC5GGq5BbPm3Bc5unEamMnq+wCM/OebCs
s5h6+zs01MnjAq7KTzDIIjcD+p0cVvzqXu0T2YNNYyZrPOHhz9S92+DeeYOPOXp0kCsdi9Ukm6SL
KLxnlrYeXUGpOJQqmEU0jD6cb+xp22TpkhkdyCaleeunuVKw783CcvqM+mWUvK5qHsDMcvj2F9fx
He3/PcW5AQUpjPSozOidoD96VgqzEOvkwB0/VZxfBvD9SjNbec1qLU5Mgtv+KB+bd54x5e5Chj6A
H8RUlkvIMJ2kTWOJXod3X4M12vgTR0zFgjUUAjKaO6Td73uxXhhW5JbeCBPk+KhCFEzA3Q1r6w9q
ZshOxnyRghnYCzZhatLMa7olHSevKnyA1XD93b1Yh1654BjwcRc1VFEMDIs2Ro1CUSt5We7ZabbR
v+y/pGTUSwTHI02eQu87hLlg+ZZvFqBzqRwp0Ldso39WcO/vUdBNfzmPX3wNHjyPjFBLTjSK22ll
QRKSkK15CT6e66/nK0/A+f38/9o9dr1jubj6dbHRKgQ8k5h0vKkEffub7UyvN0iMbxS7g5LobwSF
hbcogkCdA2HC2rlMWTAd5WyEPXJ/mYNfk9bfKgwXwguGsoJqaoBIw6eRVOIGvmpi5gIVbEy3K+FY
JVHrMxrWAq5J8Ckw2hrVep72wbdACFcisF5iW/vR+dwNjgld1PqkjJfGLUfinm9nUYPsneP0GTJh
O5ERRdPzkn8Ww1hVr+uwH3OCI222IY58upTkOZ6j6aRqpYPp5gc3pe8m08lFlyPExSIw0YEm4bkY
P9JVYBWsscmqxLnIe9WRbtXX0E1EjnMoBQJ9fv+zmQ5XzeMGbeYtCZUn/2rkXSrnJuaDv5sy3OHA
XnoMzR/M4GGYw11qcKxC6FAvuTeBANS80qh0kXCuAXTgKYXfZWsiQftP4/U5elm396EwwoPaw35J
ZL3xbcDRc+ch3FOT+SZvYSuFVp9iUc0j1T6ChOjBI/2TXBv4xLQSvJ4TBW/QfXDlxOIa1eClpBoL
bPTiX6+g+OCxMnNr+ajU5keoLjiQI971nlCDK2NHdmeZ5XwyHvAn5kYpg6gVhvKM3K+lrCa7Optg
KXawX3/HupLFWfOB8DJXInzNHXPTSSyuFfFUdbar7DRy+KqviUT5DzxWM0oqugwXX8HlJmScymdb
GGZj5kJsxnJ7RITRmzJcXZRfvx0dFicHjzo+0MRFMpQ2G05J42yu0AWWQgfxXDo8UrISvx+C7vw5
eNXm51V+AaWC8VGBSxq+pBofUA7gh0fNjNF6QjR8koDUt0MJOC4z+ovI0v8I/jaycGjJj0fkZUFf
oGzjoRH7bDi/svEdmATaMsX1ML16WeZxLKqLSKMA2PkRw3fa+S/uJIQI6WYCCPD/dLQ7bzl2Rr1Y
9yK8DuoMrUFVLjYQkF9FlpAFcG79fwjM6s+SHLiotnrxUKDIH8WA0lg1mIQI62pFoZtemFakl3wo
Vb1dM95TpVmrvB+N6izAvUedTYuAs9qHgvCSV8THLuvUheHbvPPInzgp0Hpf38rOVVwhXBhC8lB+
sBIL4TQfTK+uUvSaV0ErKBKbkaQeR7ROj0H3dNbY0ox7OWzvcFvLMAz4mby7iTg/yGLk41ShAvHb
rW18EClFVH6bnA/J76C/Iy/EuhHyzFwen7zpTZgynxf4Be13ddB74FstHSX8YnAIaegqCqJ83ey3
o/sBLHZQS7iX/aEIrjA2jC+OUCFh6ddbAm1jzSWAvV7qK79njbjaep36ATMlZkIr9+gZfGwj3zVD
4jgt6qZI4xs+9wFaTt3xz7ijL1IXsKw8Czlg1MB2UZDTbojPe/YbmDGB6EQuaBjFHcmtz/JD2Qh4
+1N4LvkUDymVrmcoMS0KnKiwUH0P7Y3WnRekcRSRpFo8sqUQyST99KmOhEzREU0+2n1UloR/a2L1
LdepIzQP8MM4q3JKyzFUZnzK96mpIkgZjI4eBFMdYSYK+T8pE3Gk9ToRZQBs1dL7yL/3aVYwDMRk
gQpDBm1Xgg9BkWMTGmEQVHaUGBXx/6kF885KdW+qV2VDBWOrRXoOxjC2DQmZN6S51tSginJ1hCMy
/drJBrAbK704dYUFWroRXFZTQ4GYdT7z9ecg+GHfhAGpCmJADZWuzdXdFEXRXIZ6vMS2EoCZ0eWB
mUvrAXOhvJBQPN1qDFgyvnanC8T2ubEThbZVxxNvSGVrfJjxtFcEscXqI4fs7cqnoe2GHSO+Shrc
F2jJPW4T4eI/X0j3qo50fGEU6epLlFDL09zSLsxOuhv44PN7wXf73P0CrpLK81iZzFbs/J24uIVz
DONbhACbmbi/l+EEZMWq1K2pbhh35gZ3fOL5oQxQNBMhngDl1ym6doBMRaR1+TQy9ahJmIiA2wT+
wTEYn1NfPUSmzj+HD1AJRVSvvDvoDhvhtAWnB0WFbJFmYIB1pIMj7iJImTNT56Oogjyp47fI7WRf
O03D7xYAnsMxn8oqRPcw5OqmVNZrffFP3IK8fCKe+LA8OGb1pP/Xl7byprotJMlEAV/JJD/Lmwiq
ttGgQ5FOOiSjeL0N98Udn738Dq1OSCFkJ77LiIWEIY4MuW7z2c6A/MQ/LLQV09hAReT1Kjw2rAzz
afvIvTWp1jxdJbFVb3PWOw/3qx9ddzT3mce/TY3aBWwHGf1RL5BFlqGE5HTP2asJdZtBYc3a72Cz
a/e8/EeoYYwRV8cz0pM0QBln4bFkwsOHTZCl5b7eJ3s7LRl02GXejLMBhYcqqV1VZ33HnziIJY5B
s4LqUS4g60TFNo/I/FofTJUNTXswACpx6wKI+iYpoCxV4KWyEltyeMjHs00oIiYJc6i0Xnei+LL4
Q2jvyol4RH2nM8+leViy1+KOycztr98PhvJpnn48zr4pKMm6g9uYs0EYGUI817Q5zQdHXXyfcZvo
P3nuIlWzfBphGtJO51H0mPhlTiGoXdqOFt/BT5vp34rtVn+dFclAbrlXK683Ub5kPMvPQWXjWDYk
zIMD5cfNK2wHR4usSNqZkV6N8vPuxhgk86BXLqDo/MVkKx5ZwW1mgWVItbuOZXEB8HDh1cz9unYw
BOTmWcUvHDlrn5WsyXSLZZA6r82kVBFCFYCBH/f8SgTZ+1yrdwmSkB6KjkwPUOd+E+ufpyO5zsQM
SvqKy96GBOKzLqVFRBNEKqXCEVsfMoImnxV2JRtW9+gQ+eYfwaoTOIKvYKTlEloVvWtzvW3m4flZ
Y+xf2bkeNSg1U7z4hLsqnkOjcmRixhhFoAA1P709MJUPtbNhGqfmZE7umVMWb0ZmEywlP+pgZXx/
My4qfSFTvt7xA2D6Iuj9Ma33ZJEnKkQ8f4W0x0M7H6eNCb2eny+9Mg9eNz/8RomzyeVOMcbhZSwA
lx/0mjFVavqyrQ9C7FG4yLGUIQyvocxGh+iJp3NB1BT0iBxz77jmY6oJz+WXvWJxRTvdPvBJQ2Gg
FE2xwhVH6j45yal5BHxpAoNV8aT21XBMr/C03BgBKRqXPpRW68Cedlykxgo6cClirTi2sOukIEZk
DAXB0GcTfxWMB36kYmH/MJ74uYlYP+EnJA1Nw67Yde8ZU2lRu/PT9o+MzRuolF2VM3t4ucfeRj0U
u2v69Z8pNqJwKHZ8jAl3a4NtXvq0IiBvHHXvRAqtNNjQckLtHDEWwYIS0g+Y98aPaifLW4P9s1pv
HatHSwp+dU+DYGrT5z9cv3PmFxDwvTdT2SsfKt1yyCkFgJC2v37Lp8djz5hK6YidNjQiICjLoDoj
vLYfItJBehCQ+2xEc3Uy8pPG/3n9VzkK2diXA6xTHll4/9Gc70QIEq0V2Pgb40mbkfDKlP6ecMM9
CvyiUwKKhppmdfaK/FG31Wdv0X8BoP4rzFQuutLr3tULTXRst5Vdb6MV6JVMH+FCE3gZExKWVtvD
HCaXNZqtwCJHEWNLwCF8JSAsi9HcfDLsHZlCa3ExSq9UltOmK4xbdlQq0jNcaLCxr5yw9+g0tYCJ
7BI+YBuNNAOwEDFdbcClu651ogS5vaS1ANEP/ikAo/5PCOGvtQLPvI/gDs2RKyXg5T267im02Uaw
/Csit6KuTpMZ5N/Oro67UoIpV4GEQ7AQ3643ybJmy/05ZsihplkI5vxZdeRiQ8Yb/VC3LQwDD6fQ
hc8Gza52y96k6gF/dZjwKPnl4XAJBvNvEr+T6nmE4iUiYeLvAZmaIc0j2Rb9KZfyZ7vQjmgy89st
3Gpyr9L7M8NbgN34VqCpCAoy1o5BdBmhupNJb4sIi3bVk0pCk+Z4Hwcr4Ovy2uIww7KRMsao1YjU
jyJHeqkgkKc7Ev1Ezia7qnGAxdcWKPURPIdepmccHNfYjgEYoaZlv3iro5jag/Hr4tmbDfO8l0XZ
fCdtBlb1SGekYY30kINi3ZXZ4CgcN9myT6SMVyCF1WgB6oKsS6jtNFXy2lWjVh2rNVSy6TY5E1uz
2kv1ZMsl7F0tVmfym6gu/1GqA0v/2sVpIr2betUhSSc3R/hi6t6rluTt6XLN2NDIvs51+HsU/P17
sRs5u3xDou6moX49ZyIhzMpEr8xBWwgFS7hqy7YdRskWzadDgzGFEDoXLuYqeu8JBJNK/wDZIwul
dyR7bHPdu1Sud5LDAP5Xmedb08wTMREBvspSs36e8JfcnzM/da99gocK1FAEnjvz4L/MbgS0ArMF
AmX/AGEBxkpVdWgZavFHKytuR19ILQpi4Mgf6QCgLzFzgK4Wc1PAHO+TjQtB8OocPOux4JHkhLZk
50Rl0D6VhWB4xOCMXNSMWTvs4aHhnPhdpqzGi0+whLK5IofNm4Q85/DXmBc6Hmmn/NyqhSAxqMfk
AFtgeUWmeFnL96KI8txuEpUUkQ+qmF2V+cs73oxNulM0ptsJJH4J6g1Ti7U0pBIBapxus7jW2TRc
3X3TF+54z11t7GkhdOQ2iE4wnq1agBrGGbP6rjE4YAY2n220rDBl9YiMwCeD1CTof6qDTUN8XfEh
pjcLZMEEfijic0K4IZPyJqzLDox2yM02+X9imME9Mf5ofWdmjbK86cCwkNhygQ4C06vpgEidPCir
DCKU8Q7A7MgTebYREhdDJoiNIaEIm6sspzXKEi6q6HKeTUSkOhQG3qhsvlYhh9N/N0fa21fOV20Q
VdZ6YAlnEU6M2y6HJzupxJi1sI6WiOuf0z0zPmSkbo6kHRruDHFQ44FNmQ3GOOX4oaSPqF0udPYu
E590FvbFnvhkHnQ6R31SFuMc3yMED6TH8G7lQNBs7gGzFL5AorvX8Pz9AT+ebm9Ks7w62DXUZVF3
5t9tPXWakFq/xQoX+axkGRgZgenPQW5jiiXvu7XRZCqJe1VvTdtOpqnmi7vFNS+WC+XWaajL+8wG
t4GopDQyivjOFlpAWwXmIYDGz+3ijmTZ15X1mka8bUf3jhsgX1V95lpr1MplzK9GChJQDvi3cVgi
M6BU4JHPKFPo8rPMXEjWNMMkfzWwApm0tSQAFy3ZgtFZeVU8CyIUrUcg2cjpnxgzxTp+qNJgmvBK
Df0aSSC8VU7jLBBiXOt+y9/RlM3XwPfCXzMfvOKLylPu2cxTVwAqRf6i5hsVr6rIDDeKYUHRk/W9
mnYWKEGF9rMb1lB/WlEGr9hi4fj5TrdGmMQVJNkqYtDusQVlpmkmwZRM2nw0YlPsHeA5dnGBE1GM
LSRfSpHy4iP+rFAJYqKuo+YWDtZpJ7GmT1DAzsuV32+Aztj0FroffnRlamcPPnzs2buqn0uMhFcb
SEn0xvzDy9VkB3jtnZRQyWpEqE63BcpvN+lmr70fASZJhjP+JDGapvjZdu8fxhJ1MW6CnBEk0quT
WieMmu8OlDN2cK9g4V+wTuIqMjKhZnIjEB2EM9brMqssGtW2svEJgvOHb67rtLfIyYS1vm/W0SGj
u+RLZvv9uvnYV4IzHEnUa4MmOXIlqwwoAml5qmvCBtsrV1Hwrmil/dTyAiGsDixV16j1GkhiRoL4
167+mUbXU79nuoQw4MhQPIwAVI+4MvzYY2OfHBBRTnqRUuQPB+LVcz455XEDyn6OqR7udFtA/R4V
/gzPLWHxkNPFlyL5NwRv8LEplglLshvqSKnn0IcHym3tmRrKK7pGzGwMTwa2BbqMs8HlCL5GGNex
ce8FaXHib0MWeqYGFUkga0Ni0BUaQhEhaS712fdJxaeUvAqrf2FFKX7XMYR+nKB9MZ3mleJPaT72
mbZ65yKpNfo+OkKSypgAh7sS6rmBes9Gkzk7p9dQVH2c7ODzlis5ffRirzgBqYtGxmzpN2xni5cL
bY941SpAy/NNuk+O9NU3EIkXRPmBHvyWwjUBoc6FAAGluNXMrt1xZAp93VQiSB4VPubkFVxe3i+T
yeVtJmpOAfhnQ3S5atapJdj8hfzA1pJBsXkM7PBnEmR7+fhGDzmxS1vTky8WSueMelJ+Z/zuekRF
LfCT5o4uD7oxG96Rv9sNQqCsBltWSu2+OI/+8erutcWtXCr3a36EBkz10Yu7jZI4gktpCm4qKERL
spV2Dgiw+zXt7Bv2mCxqiJ2JAdTJ/nROacQBNKTF8DI6nMhe/R1McDFXTSwUEX1+J91Cdvq0B9QT
wtsqEtHwR9Uj3+Hg/Z2k6j0Huj0haoBjJYNfwq4s885dHELzx+LcAfIlIV3IcKaHRd8sUcklXjqV
0MXBpzoS0RWo5ZTUqsWTAfAwMg6oQkNupM8evddjDP+3GXBQxzCUL2P7GnrJYaQqU393laiMz3cE
a4CX5mla7tZGgewRzLaURSlQV0t6sG2NtbAMWElCQJpwHW2QTwiaZYFROZAF4mFCb7UXwj74r4CE
33yz7ldvJEyf37R/sWvMw3Iib9HFG6SecysPFZPcP78bJTmWI8PzkpBHXw+6rR7MNG0J5qrf8kTN
NAB1OqXzAOTIwYQY96WMZUH17tOLS89o/YsDrgjeRecLVgdO8AQ639Cr1yK1gcw/fmJCXgHre/fR
sMTYajcUHe1nK9fakspI9WW9NM/DC2sXWCGMFegf5dZUMXRlWRCNLcq3KeVUbzaWcS+YXvx74kY1
oZK5hd+/h/kAZ7LbSTkq+cW/doOf+LsBam3jaKiS5hsMq3+J9D7hYFyHvpj9crbLutCLn5h/ubp/
4Jf50vhVll0yd8Nn3XlxPntvGjRUd4AW9C5e6g+q9clRkBsg+vZY3Thv844NkR/SQaWtaOfzszLT
P/nOVBkuREfxEJCIU0LcioWEeToCEdrvUDsKzl/SPDmQBmgcT7PPdqoc5MITF9bLAtWFVizd8aU9
DyxTcp5IoGqmf9P7NhqmBfm/RDRNCCyBvrVHTB8H/Fdvprm8IWdzp5tsJxfl6BhAPQMfL4XE+h3u
trKTsoR6n00L2yHYHBNJ8S+elRMuqKUh7PQjPFh5m2v5oi4eRqlfSJ1KQOnsTPpXAwCz0OHUZyqt
mZA5yOJ38i30Wbwm4Agp7ZveCnI6m8eDyyMAUb/wFTJN9NJEtJSY3kYE+6yOX6vJe8/uohZWrK3X
CxLeGP+k9dDSWdKWcrsMAoc6KXc82er3WqEJtjqm/ACSsyH2KQT0r81viLF+iFdJbColHnig/IIN
hm4Lv2pmn44TFJWaOa+GkIBLqDTck8AQ4wu4uwovtLb2guBoeFkh6k45MdBeaXNiVLUkH1oHxROC
WqXx+KqYid46+4u42ZTbnqh/+l7DVtVWWnHdxRISELTdraUSZInKqjBFNcZgD8HlelxfKGcx+mkq
mO22tlhwfgvBQNApOSJTV39Q5a8pPR3gpn25B6ns6EIGYDTEnRvvB/tnTUm16y4rYdXoqcv52Qqp
1U9Kb3FsewSt8+KdNYsfsWAq70sAxMChDvwBilD0jrGSns7uazNrDKfA5reKRtmqkmhxWG0+7JNC
kcQMSy+kFX0fli1LEYd9mfzBAoYp9LN403M1TfX9ltwwubLAtOBkE7ivybuCr5R+sZtuH+vweit5
jUj+gQFBbQ+nre5qgm/HLPdnFMAHBM0RQDTRgGP8wlUtjrlnQovIin4fcz0OT3aeLP9epATKuHbd
cG6HdtYCTLLKZutDhZXIEJ/rVGkQyNRmLU1y8cJ68Z9CkjdLW3fV+WfNhFDcyebKhTtr1xUYe7/5
9bXZ/WrwYnfUGib8LEVBht6Va37vkHgL2SeSc3nRvTSiE0szVut+yjHbmwVwiwaKQLkD+5D36yvm
37waQm+E+VsSB6Jp0EHDYHnmrOUqyBlNjVwX2FkP1+6IWuAlNdbtdfMq3eTXCntllh7ToYfoCjnv
WihfCcwu/HztTfCLHTkFu/eWJD0xdtv/lr4umC6oqUmBUH+kDO5dp0nk6A9lt9T7T2B1GXqz7hDb
fHL1j8aYl00wRfWMWbruAvJRk8G+i8ocSweCYblatxhCUI9NMaR5l41SFF5c8BF/g08+ic+7Tfoj
Rfwtgn61W8ZVO3OH9RAuCdqst03LcWacLLj+VQ7RXTpOJYJ9mAZt8IEsjbT3HH3M8/B8IlVEAShU
hCpNGbAnH1lqgzwtmT0ngT+Wm6TwsfHgxFOUjVtaADPBttGFTcR+n0SBtFJsFguFQOfkUIddARim
IQhB0V0eSuiYlJC1OGPYutu10YADXPVyPhZBKzeLocZqdd07N0YzptHsJHa9zk9xlc4SZEdNmypZ
379LV4UXszD4WnTVK5ZzjsvUaaG5r0E+j6d6avDNm8DQ7fYw1kx+LQQhrl4iTwBjYpLKpw4GNYCi
J7vuhr9TB4VQEPARG4U2yEjDYUwkZdPwqSgqUKExzFQ+bdYbPrjsjyb4xWWGG24ixT7HEbfK5ZbV
OIYwIaC3Ivu9iDGuP8BbDC4ijKSxgUDd4NLTN2SIM/ajnGWUNGzP7CzZQJDZa5sIh9giEhJ1HCX4
GxFnRu3BT8HJIWyz/b6akMtKLZJKLrKEg4hECBghZhfiYwVmdW3WOLJntZu1QCpfFpmIg0K5KUcP
F74D5ydrBonTejn0qy0QojopnltSVnq3QYw8pXgiHupcyj+Gy8Z1xONLrrPXrzjMenrroVvaUcnN
HX0I8Y5JExUv39Dls/YujltEULAP5m8LswV+FsDSibPgIM4BbYQMDVJItz/kNaAjnKh8bjUHFSbw
ixDkEF+Q1j0u/fhvQMtneqE5wcRWQ8bx7dNUQe3z86pnuLhYmdPnsomZ1GePb+Kz1c+2cysb3yym
E+cWeX4SjaQ8a10rCeWlwQIajT/Tv9CWZgDb/oIxz/gp6X7g5a5L2Nc2SAsbpf+rJofuTkODc/lR
JAheUkxFGD74Bik1YH1JhD90JoFud9Vg3oJuqvw47hK5JSWsf4gUwGz919gj/EgUtQ3heab7MZ5p
oy3fCljPKCK/3PUi/oFi1/GdLP1VZb4/qZZRKstNWs2JrIfN3uW0inO8V3pwgp4wX6LgLO37BLHp
L02qO5RuMmPyoOkQ/16YiC5AtmxWXOzlxBiMtjdza8dg/qDpSUscB719+6ohwOb8ylGjfjsgOhNy
uzZkKKR3XzTTJR9uyHqMGzZN0LABzSLAKzYhsdlkh3RUO/Ni2zyae/XjRiCYawj8is2UELHwr6c/
sU9Dj+pnTXOAAjtIeBsyh7D8sUKNvte6wGD7aNBwAHBoDxOwvy6mPX2riuHjXzrWn/YnQuNGfxgE
wDhe5+rcCe8gxk7YfcVcfu9Oja7P1Fr9+0EMbkyuCZd56w9fhm1izbXLvGDHTFHA2Ti6bPn9EtiK
4i0c562bbjaSbgztcrtoDzyWnMnpZpAaT/A0XuaZHt3n+GwbSuYjFgqvATqFB8IlznV8FIXCDp9M
6IA9TzRYDHDiyORt/w7GuQJFI7T6nj4MtCW5MRRYIhIxkl+13RYZDcigoD9+JWBsAw5HdB+j2711
x1QVJqTyX1ESWs5STiYp4lq5oIlKPtWJzvUPui2vgHQNx9STil/XvKItSaWqxwGmQ38RxK84ADdm
J6xybYZXXQs2OfwL4nlWNm/fje70pw46TxGmRYZiP9MSWE8UkPrchTIcqJ2eA74nGwEuK7grqutX
R3qp6MXVq3JaFd/QjUh+axhwvDmSFYInSEOrTABK5EfN6mtS/ctDSz2WotvyfgN2zflc6w43l0M0
AWLOyq/qC+02FrlNxBT6q0HFerl2wkpRzo1jOWTZSfAQzPgl6B9G+3t4LNhKYJLhJQY6RNm7DCEi
BBd1B8/FVi3hloXVYINuG3lGzd3XggSh40U61u0m3Jkrnzc5T/JPWEDEAJTMi+k5gP9Thn2D/kLj
ZtKKzTuqZt9eyLoXr3I6qcWuQxWcHPFPOK5Qr5Zwr/z99hPbpCfW9d4nyv+OjzKPTHWD4TK/veMo
sOvvK0VLTuDBwcG//XHkEiUQpugRrln8xVMmIcOtXKe0jv70zKd8E3DD/p4MJ3CltX4s+XKi7RfC
8GoroyA7nFGmIpVM+G8PipOyYAPmmMMvTsq0XqfohwQytsBZNPDqTUkaXgY4AxDieFMHOelmXajW
VSyzYEfJrx8caZYMCKTQz2YcZ9+9NR0sHiIJdNBln3RAl4G+ZYByUIJnzgYGQl43tOq4nJ8ESleg
FnyJd//tHRKEJox2P94iVxZP+rddLshEDSlNaisIKGzhXAqKA5/fQ2JkZ0d+0CGz8KGDEFSxkzCJ
9ZQILZr9s+67MrKRDh2FVd0BE89A6Eb4CsGjDg9QZ9Y4Jz+qDbS8msddAEM/B/xg92/KWK5CMiGb
5AFVpg4xQVsJAYyN/HfFvpKlNWYMrp+eQ8IjiuIJh0k9q93+RlDS+eQOYvtXurFP1tnobtoBxIVw
OT+A9A0vfhvphmiUR3olNn5SG4c5uJFSrF1xAoVqusSv4Wb1dkXmBNlSGFRGNMjj1Rc/vPcqYp/F
zMM/BLblmPBYXJIx9oFfYXkgK4+qb1ddShNWMwRc7anA8TfOC+no7+0B70jslnfQBmnF8FKw84VN
S5X0+w+yQrPd/e7uGIfNLsW2yo917cAasIr8ABlMysrFC0duOPVnm8hmP/vdYfglMHnpUCwYfHjn
bgKivMRVKocZmlq1t+z+8alqI7RjMfJuWf4QmJnRKI4SN4I/44Aa0MI27R112FQdsoeAs3XaqM6f
YmhNSze6a0FHz8thLpALgcFjWlT6zett2IjyZSS4/zyiHWcsIJBIYlzJUQ7xkCGQTN+vfEGn2r9I
k21UY/XMcCkrolpEgIkdV8xQfhK5NeHw0vw6ZXh1AmiffQiow60Jambts4LQ5WAyz4ozwvFtLOeF
HZS7yjpdo/W1POn/vkHcVXVt3fGxhvWDw1TDGq9zl9Rr0+9IdSh4c7jkpMa8opfYoc7H23IX4N7z
57XncNniMRiVJL/AuituVDWAnSIag4qCnhEh23foYBZlV0qxlRfuht9uXobwcCo8BkPwCfv+yd0B
mJHpTXfuhlBaBa4EVu9pxUFDeqWQbYq2rkAy2VSZKaKvXW5d7Yj51ZutWJqRRLJGOfQLXYZPWgXC
b1RZfsNEhZQtYUImFVuL8KHmQWJ4COy0FiWLUZdMaYJW1eZKje4FK/2SCLzSfOqu2VkbcPHKAIQS
Nu0rjdvJWwD1V+kDLuCrcqLGPMTCrGhKcjSm2y248kf0NOH00KBzpoCwIRmHrbj3U5sADBArTKw1
L9n/9XKSSood9dTNvja/a1R+1JVWMyrKjkGaydZjY0hIMhjnbN5QXwfd2ZdGzwD2xwDXnI9/HbZ/
b03vitWj+Wx13Olk2K+b2iH3oVNUCzS1RwkFRSDBnfSfYV3fD+lW9HmSptORGM1G+l4Std/S3FhS
JXIpg3K0Yk7fzN1C60ZmPM8e163lb9JYCXfSFBRzjNhxpc839uVX9xH6MVZX5rUtmjQGkc5MiOwn
3te+5gZp6tBwuAo8kV/drwsjyovxq60FMMxSL4I/nxliO9gsck6rb8+PimZ72PDhEGdIxfSO74WR
AONqvbtDlo1q5yUIofZJxlCP+ccJ3NPkw5Do90t3rnwUGk/2+cEB6CH4+mQRyKALE1IGPZrHsV6f
BwFTRsJdOjXlNXbBqnCTJqqgBjC+8qsTm015iPhHE0hrsVbQlGylcc8CNNmmDnPkAtXlaydzqT/F
vU9IoQlfinZyPu7g3F4CttQ2g5UcyUO6nZNRtpoXPrr30vETNTYQE997CJwWTNCwMwAkU6IgkZg2
0y/hRQZmS1UuCMWjOdL1jp5Huj+tLEUa0vEB6uvRCbaYZ1Ki4n+bDmzprbrzZ90scM9p/ZH1YhPM
+q7ALAw9rbiuJdVi1itFAIVP08UIX3UBEKsUiRxVx1RuuOCaEBSEjZt9Emh4f+2jcTW0j62/5LlX
1oiOIBpQiyZ7kaKBwJCr6aLyGoGnVAK1HNTUOqBMetZC32sYhAP0mNjDP6U8KSUSbBlwloHOYh++
zUXfg02vIMJCT+jPmOe+cSlmv2GN7AaVGZKBNF20uHIflZ+o7Tznfa5fMp6gILmcywRbtcOJV2vj
9mbsI6MHBjWvGIxJYb0HgBzUFCURPQK9nFpBope8iMr02wVDPHml+tpsTOzqa3mOHhrxpMD3V1Oa
sKDShhAxfcR1QLYZ+U9Ba3Kg5bokX5j29PrQX5crSa7rvHD6ICGDfBq+9cprKlDFKs34TKnqBOI+
MX2+sYWNoGEQPzU7uniUg0FhLgzpwqKCyzfYDbHNqJ7K9RJTqaoi28acTwLYoOFQuNo8M70u5Gtz
GE6/giK08xekkoBtlkqt/rynkEBzZa9aIymnWHcxq6o+6AuUB/lktv7h+8Tzd1NQovXPPAt91/tN
utjoiy2HGvUmL+bF32zA/ZdhQQq2/4Cxp+NP1g78RumnuPAi+nw/1MJVVU7Ih6oF6FSfedoP3HIY
VT8+pAajl14vIIE+q1CbCWGa4I1nskf+OlXs9MyjKlsTyV6/Nm9v5+13EZbUMva3eTmRGcdcmG7z
1O+ryyoBvgUvMDm7N+qHdVurKw2f2HKByN1ICz1lWeImN9MJLXKopkVxl6srfB/KJG+b+WBnDR0h
l1Y0cFlItumM51STt4ne1KnvcdKGmQUbfw4pHF+g/LXEIRAb9hOD9wNUnqQ08ePP1HS6nYj1GZir
HdMIjeonQVEaKJET63ckZQh5CyMuALqMDj+i5XG/U+3Az5kY5/HtIaHAv4uCFsw7k/XHYFVfGp5O
5t2y19cRVzeZqqHOxb8Q48W/YI2poEXvsf6lFxs47bTRdEFzJ9lWD3SqcJl3nTIgBmfIiN1N3KYA
Ej48yfXNFeVX64SDZ8yAJ3ZR8YAnpFUcZfayWBWz7X9ajbKR0sQSUqZ17Icw5+wkycZG0pCfnpHR
YxleA1yIaNue0qIKB7cIGzkuTjCkjrPucwvKBMMOS0ZtyjeR/+TUkJ9c0ZZkp2zEwZveqRfoKE9h
8b7tvW1vGsymjOgE40CeerPYjhhUtkMlswx5g3vSmZzuzGl0i2c2zJDkxGrQFa6UCXF8c3tJ1aAq
fFvaz2ym+ivTZL0qrSFcSq46YftOY4D3qSNfihc9wEERiE6Ck7NIme3zCBOiU4yGplPvdkmbsW94
T/z2WO3tvTRL0Hdekxuzu49RtDsFt5f8ufXck1TVlnrllydyniA/B/Y24oBen5D9t5EleE8tk3Jd
QLdd9gKkpk8oXsfIwpvCnU3/ZLHLzuRFX14CagQIVYGsfH2fLLSBogzp/KPPtQYM+OfId4C2EXas
NgMpAqKRuw24mE9op4c6gVS1ekcdpn5bAJNmvReSvPqAsyVBJLdgN+dawv0KtyJyRhSu8ikId+uc
Xh9ufKR5Q1U27i/ZtzojB3pjgRnITgE30IBraEh6Um7sMFTJOWcADsvRch/lLSsRQioDWKJlzlIN
v1r9GyloGJO4eglyAi8uPuEw9sy8pK0g9KX8goljGzChhgfGzxMMpTCKyYkDIZs9aivq1mDsXUc3
UAGw2b1AiHb03a/iQxwfQ+5/vZsnQ8m6gEscHkAfVO+wQlnjj9U/jiNXxWAn1Cx970zeBCmDWqpS
3Ry+tLG+GgCpFdlmtdMP5fmPkYLDwto6WMQxG6dHJR7onj2MnrB3b+mHK0SPGM8MOPtcxxKVQrva
oDlIt5OZqQ9kzrHtngu6nc9nulU9exNtFKaemX1WYM3Msho18qXtH+XopJYOVKl2/+CVehMBFERR
I5MYkye2+pay9iWdyvJ5JsmF/7vour8DxTcY5CbXkD7XKmkeoCQ/5abO7qsBCgr57WaTVQVpc0eo
8MRyYi3XGxPyU2r0ReOWZY4LQcyPgQnu34+gnO4uwzyPvGaZ+DIG/n197dp3xQqcsLka5UdVeGVl
BMcniBVd3ttdpq6ml99wIVXaCVVarEMwgs0uac3QikTZXNwETanVwE5FUzDJvHc9ZqxXWgi4IwaF
o5zMxEtavebyp1ETZZd3YUG6NEODecmS4UQryeoswrqXphnLi9xHEe7K463Imd9RA53d7XRi6/fy
5johRgVue839PPH52Xou1l4TeLgB0yV5AiFzoq+oiBTIAknMmkZ5cbrhookVjoJ20vO8OJqcdjd6
uf2My0QMBzJdZUdaz+LE4xcKiQkj7YzQ+7RdOL8bYjfsQfbrGfmenGc3VImWDrw5j4pSm/6zpDST
PnMnMAOkA+pdw7wJcEXkyiyFcgoIAdb/tfz1AJQO/tfYZHYAA6vMA/QaPtPVR7ry/W4WpI03IYxz
hQf+INaXTqbOop5aWbo2OJKxwmo4vtmgDciL7/fv/N2anSwMDqcQd7YoqFRJUcypxkLVuLs36o01
Q9nOtVe/+TtulJGCQb9qUFW5rxZ7DOECUQwlnExjHrNv8immUeQrgLT5YKRciAtexbQoysmwSWxJ
RUO3rRs9iXua45kFod88FyOGVZPJCEqB43ttHIBPt5OAkbHlX3XJMjAF6eIj7DuHYCw3TT/2/Zjf
1wYZ7YUXria/vTeEi3hwkziqKlrWUEeo35v+LeXPXoh7wspoLl3Iuruajfg+Ej2B/IO5J4gzOX8i
pjTFYs8wEICDLxRuGNg5cv+g4RCIEkzX4bg1gPNmlzcv0RCuzIaT9StYz6Sm7OGZrmLxk6skLFMQ
Qpi2qVhds6MUt4+zjKV4kg28f8Kl+SJRiAg77q9GgaVdFYh2lXjCEtLYPzgcB/abryiY6Z5TLYhC
ZEhDQeOXY+kS0tRbbfVv7EQL4Ubo+/5bMDZLKBZUmP1vGc7Y47SMFkspHsiVUZiNrTdU11Ra91op
6Q5oCRhbQwlO+Yfyr9C3s/GY86b/6eYKf15xpz3P87+4JKSsm1pEBaTTZUPFRHj7wNN14dFocK75
QTJtqBwcHiPvD0nw9I4OpcLj+qe5qFhmQDbFCaqJWbmgYCIICW7ewizj5zzHyiqZk+f2UwPBrhqk
VrvxgSqNRhn4bNVp9nK4yB+kKVFm5NkEB+2oeDIn9rLG9sPPv8NMiQHj4mObwgMB8ZSbUKqVapks
id4zuBgghiEGktLYlb0mBzRDFdDuBmF8shFptoFN1RtWMMacUj31DUizw4Ssn+iUC8rnfWPE52qk
BkF+Bl4MoJZFHVeIksnxSv+HRiqidB3R/opFZeSUG9rO1FjbD2c9PAzf6bu6Qejd7URyPBceE6yM
uT3Y7Df70xItFaDis21arA5Rw0u1AFW5WwLRSupjdDtV0t9jQiwm47bz5hyroc7FyYQTt2zeLLHz
eZev0l/jIIl+oU4C8aRWLFDSNMoTSL/6lB1232+dVgIPGBLkJuq+Hol2kZnEOgZJsUl1XX/CsiHv
aymgUdLHjyW4ZvQN7sSqEyzbLNi5CV0H6n32Kb0s8r++InS6eecDwnSCzSfvpM8Vv4wrmuV+AKmv
Zsl8Y6lrMZ7jODAl/VU9cGcCs5n8RLIGCFO/nY/MMuGitt4IbZ98Yzm6SxUTob315M6KsR8nmgL9
iRbBJM678Q75D/PpchyxWQ0jtx1vHOwXMmxYV4Mti7HcnPM3v7OSwSONr7z+IcY8iRX/pRdd0UY/
TcuDjmkFrxgTLEeERK/U2h0Vywli/vxs91gBwEHnkmx8V3+cBEi53I0qx++HewSCkWA8kSS3JDu1
hgq/qPKXWgVhMlNAhgKtTA40y1KVfnl28WPjML0hU5zJ125nAFfrUX9I2weDj7mETwb1chIrem4g
20ueGRBTvZuL03h9cGrxHEFnLyfPcFZAUN+xrVWCN0k4htkXZfdigIvM3L3kgO2T0CU9X6j1SG6S
1dHQbmOYKIVfF6uDtg6/jRajOGcu3aDzaoH0DNqnK+CwzxeoFhkWBpV4sPJIpKzh/EcjH4Xkk7uN
mB3nAFZQHRhoy6wbpDIkZPMJV+bpAlKp0mNZTUfmFQ74VDxroK3VjpnAsTPJ7GS0E6U7Js8Bwnyg
EJT6bcRwdgCRi4wBPe5ApAY989eoa/Ur8l5BYIMi51DVpbWB/tEas+Pbcs9Y3tRVye8beXLgPwAr
4BKgwKqyRBFSFRxeY8KZqvyEBCEtYzgZZdQ5fclnbOAw/U+HmBQYjVWrY6AZUxeIISvCHQbg04aM
yOABXFA6Yjyc9mUy0p6/xruEoQj2uT+UTgjjANq3OSL6bzL0/WYs07RJsec0gRFX3BacMNp3Nl23
hq0VIyQ8voWW9e6312l5bgwwLFJbIzgl90apD8E9T5Uxvsyp9Mll7a9kI8U1sUsYSdwuId+UAYUY
RD9F/938bnM2unV1JJ4AtaFj5Ldag0P4kimn14xBxvsCULPcRwgvSxLYhMuOfUbOHVQLgRBZRW8i
UeyhLL9m29RxtKofyN/C4IWF23WURsTnJcH09pKaOZ3z+ugZEFevnYZg8aW5o2Js9XOGgplS5khT
ZasLormTKfvjRdybEmwd7tKOqOzeMUlghM0J6qErI+DCXBXT0IX+HBjhL7Aa/1SgowLa0bXQ1KRw
wNWJnpRvHCIurt2X8xI97tnSdVs8Xn8oXUBhyJMDQzFfqrBQOCdfUCY19slAMJ/uVCiBC4XRfcg/
e1muyfEfZj3esbQzZznP/bMDtlCqRK3rTA6cp+lBspyKPzjdPVIuNcHIlfI8055iaxQk5UtFIDAR
ACx2hCORLaUWvAG+J8ZyUTVu4qn8sEasJOfayIUza8YM5QoajEB/VfmisE4HTWkjf/xCgbQD/wLr
F76Kpiez553FRRc1V8Nm/xUHa5f16AJBRMpWjvitbiN+SK8h+QkU03nG+6qJM9QVpI04R/ACyR01
PFSTqSh/aWrfmqceOysADjnXgc14B6oGXum1Zqg2It0jijmnej6pLD644ktnfQSkH6xE52o8HTN+
CIYgC69ztlJbHydedQcvpITmAFmKKwpOPVVSBCvwhcATNF/DqrTToIWs3BMvNbSbiN/UaMA373gl
V5q6al6DCra2PcTGcXRsQE1CN8LvroLA+TK1jM3wxI/Oz7kFSCUdOt80ulc6jOaIacAV8WCf+KJN
NHBV0v1Awkt8sDj2LaQ6X7Sa105s5zIwkNMGpADM6zAYeZ3PSasB7knVh6fTwDqpGTmM7ILqKqSd
HhLy77PgQyNE5KQNj7CxS8MlUozz6L0WQ06JC4gTl1pz43mdi8BRpFH5jNKsH3a1CB3rt1mZjFp5
UCGhWZHffL3SwiWe9a/OdhBY8jma7t6oFGTRuDUOHyRRd/UhoS/TyPzrMRmn3XoQwLt/hZw7VBu0
2pgE2Vw2/hFG+XT2pdtXZakcjTv0uSTNoXNAGClCH7mQGmJoIj4CcsBSpzJnupot7VSXSclvj+28
91uNqdcrAWWOONu2xr2h9Pasbds2XuNjJ/eo/v9cBP7+gI2Gw8haR79zG+rG5dytsUDyb9a8uFiW
wtcI/Caknp4ddsqDVLJ6mbs3wbBJ9h5FriYnzENQ1JGBNp6PeibHVWbymO0VgRM8XP4jGr4BBq6C
oOed2pKPcZBn1YU9EfLI/DzU9u1/Zl5tQYv1+cKZoA8dnfjid7r0A/oi5505hOkREr+bBtv7JBvb
MfXSbJpzvQyuIJYwivz17lLFEbcF/Zo8gz0/BjsRNq/kH+b9U+k5Vwqsag+3I99O4fRqltHF6aBH
AoXyaJywkGR3fa7C3U5htQbERS7lM4HysldUDmJkfWKW+YU7RwVXApEjMx+/2llG7i1uItsPuba+
87QjfvKtlWuu3Ja5RYeCiORaK4SP5awWU8ejF0cUmSPcR97mcI99VF4JGE36XDaSHg8sTdJe65Iz
9aHkaJ1/7F9UbX9l/7J0JzvIr3O1+LBGUlEWn8cF/nSBcYc01layA4bPvN+zd5G5SE1D1DNsZxMn
IgULLG3IaSw79dtl3g6LaYg7/TKT6NCuIm8NtmuN8ftOEBDRY/Pl8izsILCxjdALYnFy/DGzehzm
qyKhHqMBTxcNihZbmy9ocbV02NsPfFBcI0Op1mrXtjc4FGYgvmr0m1a5E8XcqcV3lMJyeEUktOSo
GwAM1yqp2FIaQaHUbAZbiTzo0BxrcADxD9SciVSVFNy4sWA8iqVIRfSmfAWfScpL63DLAN42R/Me
LTcKvML35nwrmJjbQEWeonPGsiu5si7MqJDYncuq4Cy8SPYp64SOolMi+RvZ4MbofqTCTyJGCRKC
iD2BJ0pmlReq6s2Y5Z4Ey9fCR8CBBlsYgvud9+/IvlsN4uBIw67WH93Q4HhvAwgk6Hhyono/e4Vh
fb+cqFTP9dPxxZCva6l5vMf/HgOJ4pAArBBuzJfjFUq1ovPSP4brWry34LlpI/Mfatdp/zf5O7Lv
EPfYB9+nZKJefElUzg5fdhTmALe4+u9KQoabrt9iATvg+zYan4Xdw8lY3sMS0HEy9r+Is+PdG8i7
DDnmB2EJ3vta/dtQmp2ew2TtR6HrG5p3nn/W29D8zL7Owx323g1e6jpdCXbiiMWtbQ8JLbsOag18
ibwjsGSxd7FGBbiBYkNlMZ9q+dKnLSrD99XUHNnhS/pF0JEdstJuloMJdq3F0GSPA51O0slzQAE6
c8b7Vs42uiULVYS3E1DKTwtWdZpluYrRKyhz4q5aGEcFU9hqIEuCESvUSMq4p/TeDaXEm60zsUmg
S0qplUQDxkfnbDLDVS2y9Rbst4zcwSt31sob761wqyG4DNvUm27VK1yeRdV8q1nVUunQsxGZawsq
Noaqs/jSEmKBz4UiiK2SdKFcT7w4bZ+VhaPivkg7LyCruGgLF1xmM9p9XPgA9rfQ7v2B/nIDhDon
BD4IQ/0rlID2lKla3nl2SIRLTL9TLfnZ+focSf7xeYEAjh2362vR3U85/zLGXP0FHFfg0zBnVIRj
FYvmRhYCUaWJJ4kVSDrF2xzojNsj/HZ3rTHRfhfqGN/le9g3z+68uRu0n08z2Z8I+8PFvOMqsTBy
AXMhXdW6Q8smBlWMWaGzqJ42jvucfz+TczpwprazYd3P/n3DLXBK3CVfLZjnJ/ftUbuNlbDrZcJA
E5Lr3hOcJsuLwUlvAZrJ1u8PZDow9ljOj9MMklxRTwkhaWxdSlkAr0tkmiO7Wi7VzboCFvSl15Y/
5+Sc/Uj5PhG0pc8rth9RhKf1+8hJxmaddccpV2/h5H2tbytCnWtJcCOPWuQuTSjbujIq/nqNugKO
63I+g1ZmL2AmcGqvGNf0dFM6YOFb6yp19xlhTqFExu5NxlSV2N5qnbTzjFWXcHHqR0Y86JHnQEmz
RWXbANzcFxYt8drr8fEiXHhip+OQqOkyaNBlN8LGgXHqoR7sYuFw495PIeudzI+0gv/eRi2X/Oqg
IF304qjCirTTSHaG1Z4X9mOxvjzDRDYErjpkwZJThevviryrtuRDGaIaBscNeqqSqWHl4ggKCQRR
olqYJN6f3KJSVPOGgXlm/6bRp727JJl4EB7suBl/BlNroRsX78W+3VH8uBu6nWbCq8EvjlZjJq3H
PnwCHyEj4mj/3Yhcrj+9txQLuAvJVNaT5DIa53+cj+bu2dnuopqLIjTAzBkCmgp6+lMxAoI+dSi/
SdvzLVkdGHCkG4UNBGIrdlIJ0bLAJfUWz4Ly47ESlRwLB6RpvKal4Y1LPIYbTg8Xzp/Z+1WIStOM
P3TFsyfX4DG6cZmz3aO/lWYPa3sDBQtnFX0VFkrqYa1SWeUfQZW2hq6oUkgUNKkipMIcgDPnyh/D
2gatmjtBbeEdZWT502Zhbjg56ogXj2ZdNTiInxLGxk1GPZYfrR7AFLD19JYGCa99LQtoeevZnRDF
KDBbNWMCKqwbRMUP6KD8TbhESWGbF9h41OXhSX/b8Is74eXYkXp+RtzMF31V7B174c8lPwvLTsuG
nvI1u6/3NYYHwuUuWxhi9VpeCJZjEGt6WhX3qSSB1afPML6e8vBEolb8meJNdtoA1b+P820ZmiSq
wn1BtK6srrnl9zI4H028tx5C6eyno7Zmpv1GXWygUS02oIuv8zpJ22sYu0q8dAVS7UuAyrxWp1x2
IUaJka/hpSGN4Q9860S5Qb9GMqGcInCCyzE072d61GUZguwtURGCsqL9HStq+C58gmOUYb/FVqS4
yxIIjKiBOdCmVCS7txWWalaEUMHl/WKpfPnCeLAYcZ839W9YexpBmzmogllwN3f3txqZz6Vhie2i
5wPxjyaB2josTvLZYnuIgPMN1/14UsMTbfK9E9heFeB9ghavCoLRk/FMK5OPTpdmxiOL+adZur3P
ym2BvNdcAWv6L84ry60F7ZlN+TYOcs9/iZckYtbfObVtidp7juqJ6FLB5njEh3HaZyMUQvhMUqbO
YWvoXci+EnALD3JiaIc/jocDIVajPJTYwDwC2mXLnjXkCNEIMCPs93xXntA9VjAUZvUoXC2lPpwO
WsU09vRv7jU7CxxUpyHP7YEGv0xYKXSZd0BOVLd3717xUi1JJiT0dhQ3wnTBgkVX9clFlO4CeBDG
b/dl4/D4h7yFA86NdM0yHSs2DLhMlXeE5in+z7VgGxkoiGMYHLuYsl37IKrA1Kc7yZcOlDnHg5iI
d6OtZ1LWrSa04GgTjWcq8JcV9G07f/px8DxeUq15ljzTP8VLtz2KPBruVyM+P1ZC+Ajmk2+0ukiA
2Rs7H8FtLvZT6yDHc22MDbNni04h1qFqfzvhTtrThUEuXoh7K5nxhnYvNH1j80CKuh1FyuSuWV8b
BK4lRxoKG6e5kZY0gsR6qUL5JrMiqtfKUjjUzCFsYqv4XELqu+NLl5LBspwwQ31Fh1oXr5Z+9tiG
ITP2LLo/6S0SOipBKYuubq5E5xwJFP7WAFRPHW4vO8LHIHDm60asugX3bH+Mb5O4emrf1Pyt+N0a
VsJ40VQLgNatnMDy4dMAogMiENml5VlJ3mtU3iaAYIS3YjVNggH5/7oZkKPbSdnp01eo6gRz0d0X
ILBkNgCgERNEXKruAtR7caVwHtIc67sqarA6WmcK3BFHekgfw+kxHk404P9ZpHlRjcXUrIb0NUjK
hC+W7JtX3bE94XwPptTvfwDRAg7Thxey9lJNxJVW2FOZ+TqqWU521iNiniMYWmmzV4+E84P61DCj
czNc94I+TmgEhos4ESIYqgNntmIJ5ZipbzSmnaCMXYF92YCULgQWPyWXnOn/VuUjCxNalM7eNnKF
klE0iH7ulK67ZZWHA6nJKzRKIFEFBxdjqpnx3aU24CWYW4AKLeB5FgJIr3+VWG/lO+axLOT0JLkT
skaSVW6VoiANfcuFhjAxZKEOCOPxm6k9rSS958J9ZgUp6Rrjt+6bJWdaoFskB92ZfO9PGOX8+YWB
B08KZs/pb/QO3hFBdkfyHf8wrvJ6ow//E6BKT5gf3nVjmZyaifb/jS9r+4+yn2893E9SRJ8FI3zP
BgTufAJFn+d3WAKxi85RUFKeZrgUxhVP1nwmgMCHJ+ZRTJkgmv75L3gYUiWyHwXKTlbtcEsH2DwQ
NEO1nNmXuyCpTHcEkwk4t0Jp5zYWe/19GeOdt6tnSdB5dJntf5bO92Sd4aydv33aPsKNG1I8lfpS
4sfQHXSHz1Go0vBgPq3e0hvdu1ReCEFGan5Ma2ybLoojn9sIjs1NJYf4Ob0k4ohkljY3BwPa0+qv
tHcgWEzxF1yan11jgDX3Ut2qchhm2PtiMAuEXKwe3p5FHO3AM6YWgWSysZUDlVj4nr1qSBUSC0Sy
fztK7XtVDaTa55RpnFALBfabJmRc69C5SxGIm+E6VkgR5P/oxbClDx41ayt8PYxpefcoFBAXNPoT
M+ptxnmbz3KIOKg1akblDHJw9opRZehLZUb5ltg5j1enxlNhB+7vn4Ol+wiwrGzelg6ESbNNefjl
tWDiHdyuTr6mHvhUxXpcEDCJkNAHBYlh8EYEAor943bGb49JW2ZXhVlxSA+7Zv9lDwzrdWS6eZC5
r1SCa/6/0Zozss/fHXq8HPPJWAXePbQBnUQhqh1JLwOjl0XPFA4+gRV9aJJGEtiRpm0uyIgYaf+P
qBmNcNKHpcAZn5H4jqXoqfSz5qePieDO4daw4+LYbSWzrw2H39I8dlG733AJHXkHcG6STn6QIZ87
SNX1juOw0PTAt/pdKrk5LtTwXiVC04Jfobj4mZ+/+DpE4sfddEIWULMgKvMirqdRQWlMQ8TUSJ3I
wWVVl/x95L0EMXkowNM013QqD7kDMwsNdH2CJDrpkDhJHRFmHBW/3v35k0OPtX9VjiLpJDXW/O67
VSN4y5OU8P829ZMveKhicHGi0/HeqfOA/RvtxgfzfypCfn89MWKdGNFAMMbtwyrQ3XSoGhz2Hl/q
JAKe94o9bE4iR8OvVWQWLwGIcR3t1U3q1piLJKw9yLuuD3uvKmRz94qgflHURQu6y5sFwyDksXGN
656MXBW1FjhTOd0qEDIs67A0loXnKNSWascn0RfmMTcAjKrn+GEQZNWy6TUpeP3bcM/sqQKCPee0
Vc/YMTFoyJpnDbBGUUc9tRpCV7DvGVaDC0qFp90I3aVjGminXEe3GlA+OBW898zRFppT+VW0YLEB
zpu7G4MWeDWF5W6fOkAqdLYdKwGlhjEtIzKucncPNXn4jxuYGYUh0f9t3jRDi2mtrz53xZjDuLZT
uOSKE29FoAw+H5NbP1Iz89fvzCIFIdYvdCcQYk+PBsE4EN40uW1N3FhxIrMwhPTck3QCrYwpr1Rw
0+oqz8LYwPUewyxpxAonGlLbYyqT2Pxxk/ZL5HlmY5T9Jt38KN9VEg3CmuSNIA2NpxAYkmXQkKYO
lXR+mfpMRPf3548OEEg91t5erWE0JLTP8h2mKKBABYyHYipTX3PqjrvEANnsXDC0GAsAeSQLe5yT
Ptl/M4Whd3gVTpaSEVH5wU3K2ES+cyXP6RxCa3hvDzA2y6aZPJvLRRFgFyjXdF8JBjd9K+sNyE5A
O00ORg9gjAQ1jR2t4TSDECupS7CqwtKJXcv9fesKc8s9fA45zv8E+Mj0hUVHHe6GEct1vptvRIbj
Z02pDMrHz+jxa5eUT9e6laDGSzIvQqR/cQq1ycFob3AL3k46og/DfjuCyEd8qP+vukp6HynDhVwU
SJ5bcQRvBKIToxFmbtW5MR3yYfodQHh3FvT1T/nXMlBW0m+E3eFajPN5Eu+K32/L2yKxrEuY+/uv
2X63DhAd9Tyu/3uTPe7k2L1vgu+zFlR6enEP/uidxzU/I6DIpUIBRy2kiEaMz5X8x8/tjuO3bLeb
SrYz7iy8HiIQVzkvNdNs2KsWeVYsMUy1HkjCHP3DgLbClgiPNhF4ZWhogB/jwysMKGOCdjr+0Z6O
4j8vaV8b4wBaaJxbR9cNRWC43AoF+ytJA6A8WM7E+g4C3YN4DKacwMT+4X2NlJtTTPCwUCgXZAUW
IHI4AJd2aR7r6ypXAG+x8CJexizcnRRe40OlRIqFlJ4dvIojl97NMNABqU3KtDiNXjrXx1Tp7NVF
V37F9JcLuaRwfwE+CPVoCKbZog1CZJjha+R2DIs+0nbpkf1VQJJoet2WrLb79nT1JHjcJ/CH1sbW
Tp4HKsDK7kTZLIVn6ACuIkScmLdHb1oCwSQOMFOr+ivNdvZVeKmcTa+kqMlIUs/QLZtaGUg4mtH9
YyxqrAMUI/kEIcdlvOBUkjQ/mMFN8xuNxuVW63o4RpX12I2R8GnVLgg1+Al1zYb5t3sk6BphJO1k
d3xqXoKzupGcEFTiUOKjhReZFSz1Krx/eVwQkvwSo4Kzkt5jr2N7TCa7HuDOlRumn1ZwYa+jX4lB
GmUVEUxFW4I03mF4PtiqKg0zmBpOj+8VL/TttSGD+1dSJGF9KfwCNzcWmeKBZdEguZywy7YK1HJa
g5Uy0xMftStPUX65Ah6lu3SPbMH7VVIVOvJF2a6Mmbb9TtLETJrIQEp3g/RclV8xA2bniTUOONKq
W1FqY7royfNkqLmQhjNsfZAjq0HEy/c6qIwm5Te/JVEB9ZEul95xUJs1t+UnMHhDJRPVF33Tj/kA
e7N81X8rfFvwXbr0jVI13Pk2mnehnbaF4duCq2dRgiohS9roIjnDkIBKR24twOZJBjg+sPqsO9W/
VSBH1QSL2geVuVU5R0kyxz0IMawcgxMVawDzrWLkR+aTgn5FY3r/p2I6b1R98niQxN3ASxhyuJHx
E+KjW/VWhJSclYcNCVSlHk6GhGKv870gmdwyGiSswIjf6NwVDTW74BpUa+upyEHOvbYOoHgGUE7A
XLveu49vXC1x5/7lHqqGNusw/E/gieHkmWpj5+0QOUUVkkdPHzuAkywwbDBDRE9HwdtIDFbxltbf
kjtxV/e+Jbj3OnvL7CtKSVccO82K94xxAlvuyOkHB9twj1uAm2o5sEW6vQZn7x9h2eSeigd4YYAC
m6/glYaZR0dLBEqWOQhwJXmtCLfQLYy1PhzqPwpnJbberYCd8w9SLg663PIstK/HYxrASbKRf/00
0s7CIoIk39YVdSiUvx1HBQstblsaqQuiQeFlksKpDIUye92j/vzAu9RtZ/95xZsjAGEoeUoEz2JF
Oqi8kC5Ilr+/8mWKJPi/+dd2OrfY9dK7pRxA/NzhSaDpUurjHFfAYM8CJCeJmYRZEyyu4mECVWc3
w0LVRWOvFbzt/wv4jZpNmng3mIzgMEwOIO3ZItlp2PWOTk0DFbb4lqIx+UW4Itgt7mWbi5R8kSxt
kRE2QIqShQm0Lqep32VfJ+N27wyEraJUUlwsmp+6N0YB38iTyaEiQvVA70Be7kLs3N+D/mvGu5oH
ZfA0/IitSYMRd1arIAQBYvODYPyVDD4gG5JfxGWtqfVd3XsNcbJOeG0Ye2Wn1eN/KHNhEsebg3b7
+0cL9OhY1jAKrqOBDaWUSe8CKjqs6vYMFqPCSoftDsz2qbFjoXr264ulMOQpk3T3Fkb/CadHZfA6
3+yE8KoDKlo0vbAUjOY1bL0VoD7fvS5ENpxx4zzoYU8Fta9F7ccKvvHu+z7jTCJTkI0VDKaGC+tr
L/Ai24jl+RykmfRZumSsnhrGj5Tb5tI0yKjQVbpUtZ1+jzTtEwG/eJS/YMXkmLg8KP2TU32Zc+ju
uYkRx/u7sz+b5QjwxYZrhvowB5oqFUaf1j21ReeOU9oXyG+Xn20sfKcqzd2ZZ8EqRJEPWPzvW042
ITdWAxGmfuWfr+zR7nT2CKDG5oi2u7MzcKxu0bt83ocSWRljduxN6I/4YqYzS+OB3aBbd7XxuR2N
wvAUTeRIUCB7PZx/9YNsb104rVAfiImUeHITIynTTG93cr0FjlxMXTLnHar/wtyRaEs9GF0vYIA7
GfgKe2C9HF5pM0Wv3Q16aXqeRPhsH5cFGGA0bSXFu0Q2iTZhbTwFIO4yGo6M86UJXTzU1HRuVpLC
JLk86IfJT+7E16XU/mcEp3k2odeqLqTgsFhW/Rdym0xrwxVr8FnyL8Zwt5Xt4GmkAFGOyLldY8GF
+KbLCAgA/wMb2HOfl9n3B+0IcvEaysxkgasFw6z1Wx2dgIik2eMw61xIQOti6Q6jGcNsWOJJn2Aw
VQJxOmZapRLVIIMxk9cOZfTOHsQlSlyPs9GN98fTHEUWNV0Ws98524lz/wJumVMvTqmzy0RyVqkm
OheifeY8ycS6tJP1W910iFf3+Osy09SwuDvX/Bo8fFIiKJOfo6OWcrzF7ht0U6OAS8kOq3t9ibSZ
mGKjx2NNRi7drKcwWU+OvvwnLPE7tTZDge90N7pQUR5ycgNLXlj6l3EcCnsc/5IwyONpYF9vbOaZ
N8aNTMEflHREz3b/S6YcruY+HK7iBSYKOrBTDvaMvbWbd6y5oa438Oh8OmYkxlWqqjW5jf8hnI4O
Om33hqHKJoqSuTJuqI8zxLnWytq26ZPq1FqBMiezavK+jMYW45ddvgpXjPacJUwMu6k4yJjAM7jN
Y6q+EpvQMHOOV0tF+umeMtXcFhAZ/iymfqtZnoA/9rFoCzbcZFy+pFIRYXRyopV/emxGPF6GWS2p
+Ea6agL/ojMmVhqfKL0PhGCsQh1Z+r6/xGhss9lVFSJMy4GwXDw/e1XTvOhaFDN+sIFbKg6LrZyL
gKJKtxDgKOK2P1wg85RFslmupY31C/qn6PP6AzmNj2OZdnxHkRjCLf2XYFN1L21FehF9CM55jjFU
xeZbelXWwJFCOjqIhtdVe2Nc/rbaz255EhMfpt7IdB+SHtJN+cIKhj1V9om+0gNzvqdNHv/EB2je
+eUAnk2YHAQoVimR+DyGh6WMSaVnSbqHZR9Q16MU5vnlwQ8qmCz6tNu34pHdlCRg2dQ93teI2V29
L/8FDZPQXVeWrSQQF5ChbJAGtNibcP1h7KsdjsQ632Vm/C5KfD8mXMa1Vn7G0i4iygJk980cso8d
XTypW/ggc7qPGxH4GFH1ENIxZJrxw4md9wajOzoy31iBO2WKNCkuRP+Xd3k8MPKxa6rI9wbTMreQ
u57Xk1XFmTK30cUsQN4niQunH8CbtW+XTV7BeWaynjQ37dn8GXDPdv0yZEuVeQUHj++++e7sT5ND
lN50HKdhB3JgbuujoZXIQDVA/6e15J/jJFvU0Z65Y9vB068TN3FbFJLEXL5KOa13a7b1BcdT32in
YRHt/3hlSAMG4UGWdHMKWqZuy3HleQewrULcyqzcRKu721qXKSNYHH6SxGZXZJNlD5xYleaDtREE
nVnWQvUjsBCMVpqWE/zsmwcryDDr6j5vrMjfwU5esCSE8Ju17X5cf/6wo/w1M8428jjaEJPo4yO+
RAoAVNDhFHwvDNzQQ0r8HxlKRtW/KleZkFHaUoJ1pt71WyPXFXwGcmttpBeeHmnTep8jCf/IcO2H
O5u3r/FZd5FUvJiH+pSq9D3IXhb9q0oxUYeQPQ+NrMC+5/OtUoCK3BQ28WCObPcXBUU7dp70DH3S
YkzWLSzed6RWJhKPpbjETKbqSkTwS4jRfUW3NHmL3P12ECAzjJt5+jEPFpwBNtMOHFpXKIk5zpy4
OhSSW4hfqqBy8duSMIBSeGwZhEqK4KZNZUDIVoYxjymUEUHOjbOoDkdt9rNJaNKa9uIfUYpWnEmo
a/Rit7i2tVkisqCCoVM5x420IwNqxp+wfkAg7jv2/j6OgZXSj6Cw/HUBJN7MhcswDJhRPqZL4SCZ
Py44QB3euCIExMiFk8Gm5gbSKSI3oU8CjRESvCvsw8xFmgy5aP9osLkE3VQ6tnez7c9w+g32Q77/
e0jz22hklMVoV8LfAlJAm6/3jl9bOa/60N2qwpH5cGkJ2+3OhgxTJkE6Ljb1s9iu/rX1+76P1346
teZZeQGihqfjrB4p7kQxTMFD3flcq6wbkYvaE4ruF/iCwYaspQar3CmYMjKSpvBgg+6RO4SYy1U0
HmeBM69zgHKl9ZLjTbQT76Kn9refh6EJujoJTY+OUvMEhSw+EyF4sxuD9xn/i1/U+BXY0tAn1swm
nNbEWMiBfKeweQKvB3grgTY5JcRIkUJKQdYV6E2EXRKI/ZmUO2piGXwgWvjEt2kcX9rkB/4cerCT
EseaqTgm+q9bCOsal4QwR+8PMgXvJ5cF0+sLoIQBELYSaG+I5UQNriMQjqWVJ1tNWws1CJUE+R0b
H9qnihMFpH/RY2wl978jqs8ASRxjPIPlU4bTljBLBq84VEYMksBgX9Q4DP6zrDb/3sxn5LQcdfKo
3/T8qsDAQiuQRlu7LGu8HsBl599HzGdp8rUeBuYZR/r9kIQmAxK5/lTrfwTc5W0Rm3JTfLVs1o3t
iRUgqe4WPLsDw4w3wNsC9yRNV+12FT2jlwhT6W3fjJg2xYCtwb6oyKb1HO7pnTdg2Vg4kIHxrdtx
DJecBmGaEJqQzP+mDmEgQ5tSfQ6pHqhTlsET/38vtR2Xg9TP9BTdB9qr0JpdtFfAmM4dLXeK4M0L
i2kBMcnis/BD1VuggE/MG5pUvfLw7YrFE6WeMCygMyX9vdVT0uS0fi0nOz4vYTP6g45YoaYCp8Nh
cR0jgBJcyr7Hza8o8WK38XmbvsogYP0iXo5RliYf4OWkU+SxW+VJRjDTF10+eRgP0m+KycaqHNuz
aveSvUbBcnbK+I1isdFgAelTizF7izMee6aZ6wumQhZdk65I1N0FLPxSz//OLCOFA/f2g/C29l68
0GZ+3RtW6yu6Pas07IuyJ7FO2gxQ6z4yMxJYRoGyPVMtfiT8QEvpwkPg6sJXn20vzTcPfezwcPNm
toTRdG9zGthbm2+Hv3LptQvfWCNy6urJfrVjP00rgLr11rc7zxhGhgXix33HDHUFwvpflGgEmoAv
0WxgX3LXX9EHqeBm0K2V+7zSXcmOfiSpYdfhRQMNz7SXvZqHZEihL4xV+Yb0pToEanDvcBSYgxnC
VMeKTaxSUwSAtQeqY9Qpi01wWpEJV+oLLvnDmY4/aytx9TQZw8oXjwjuTxsk6WFFbZFaDzVDb4Q1
OWvzQ3qw7zdMRnHWbEgpU3oG6uwUvahwDqzCYsbKxNLpVugqxmHeR23+fm9ZHGE/a0n6lD1VqS8J
mj7m7XADO1GvU+XIzy+Fz3kBZHB1zZE+RXi1K6RuucG+fhExfEfIK2kzu1HNB5qM584hjhEi+2Ny
Q5MIZshMXgK7VV7DVLlGyxv51NE3bWRogf3yUmM6WM8Xtf9DVL4gO+ucdxTDBiFket9JEhXn6dWY
XwSvwzDEBe2hfNGFqPhJH8KYcHQ5e811qUgCiUNUcVs7/Tdrok4EwSmO7tqvSv2M3JI/y/kVRJaN
uMHgjgpWh5xzFYLQCzm+pmQBy/+758amRZR0r9jGh3PP0tXDtbJSUmfb23z4tzdnLaL0AFV4eJ0J
ZkthEatd/JfFvWNUfVK4UbVMuERMofb4b4QtZuk5y5TyP2HG+GBSyNK6Xm1GgPp6NmDhWulClRdu
7VE3peiWbu6jE33QsOv+anJgG94z64NxRSfCTh29b3wK5sJ0TN3g+nKpII5fdozdqiUPLjljIeDE
9l3FwgcaguexCxsCtA77igtNpYt1fjLCCrsN1wovbiotirDlwpcu3RGjGRvCVpap0Zsxtcsxk2sP
pdA7x5zu224afPig+/gc+4dAmT0cCqN0uk1BWgs09iunL0eeLB8iSeKup0FIKR52Hwdfyj9aEYQn
9crEmuWZns53elQ3+WIup1MUQqxchBn6eYLj2D3GbxaYw4opK4t4SVcnPjcTBQ9lAORRKUCGK4zO
JEC3uVLiD7b4Sk+9OnXJHc6FR5Ygxm4VCm9DxdlWDv10oxUTkni3HYgdvA5JUGB+BciQVNJrDZML
DlPbeiF8FCj/LIybHWLu2Q1b1cZB89O799GSFom8AesQZXrbUlaOydFW6R0G/cDDA832bwJKpDCE
qIPP5f/himQCQSEgla9HcUHeUu+WuQdYb8dAxuVADO4C0KELHrFyB/+jkgnmygqDQoHpIH6+qbks
xwIe5nCZ+4agSsCnGJg5UFNHcJjqiRkyWK66CuLds2pIefIypjYlqvCtjdqE4MOqdAjGli8yOdch
oC6fs3NrbA/QBfQd8wQpw/x/QXvBAh/NXFnqs3zrTwAUDt5lAQTQwHFOrmw+c+vl6p+bsU1C4NpG
d4Oa3VgSQC+7BcUrNUIoW0W48D5ZqarfUPTGj8YrIUgtZun73D0A8dw6zaVn8BTm0XR/HJZ2fD8f
xWpGjwD8sXPO5uCjRcMkPSHJx+B/KsKHHNEdQp5afdoS6ELCRMoHwR/zvVgIxOIYwi8MDqBMY7Ia
7H1GRd1zKeIzW5uRcbvag9xw5TzJ5SDR941m3gGsKEQOEd1EG/S3zjxWHRFkcxcfwTpoQBT09wBq
T4F/zSRZxgeFx+b/5HUhjBtzVq3mtJt3QoB9szAUho+7beaHI/dFJZ/g/TBa90hsCRMn0jp+lKLN
iYoWPUrgyNVJfFBUZ5hvGFawl1BF2Os44Xc0f/77wcDjWsRIMcaoQKM1qqtkk9jS7z4Qxo6oFoYU
uGbNLtwokbJqdTYeoZE/Jd3GawRyl2h8fK1GFBFx16E3M95WUzqzhI60tJLiwNYXVQvT/VlQrwaK
rQrXWOpB4hjpZPXMY6lZWtzc+zeDRxy/zGJnzRKrI/yMWg7uZuteTsNdJ7oyOM0FulIQnG4l52zk
XjcVNIWWosaA8rHo0sXcMyeMQNHQLVWkPRyNioo9k/JKMD7gmQ2CKnggQK44+dU4ktV+L68CIzoj
Z6wVAtg/m+WKbdfH2W6wSf7hrXp+4fU93Tv45/MgZIMImpCAytPH4djYdlelGLf8W6ke+Dy3+DhI
TRJj/2tODlu+rowBFNaPHzhfHwc/Yki8f22/IBtxi6IW92TbbeVqT1Z/Jkd+62EWQaLV5TALYVrT
DnAQT/yx22AVv8MumfKRi8nRBgUdHo3gHpiEdGyo9FkpYkMSXdAf7ruUvuD46ZiAzo+IalDvrkNz
Sm3nuwj0i3QGCO8lh1wUFIn2vvZX2frvQ9SYLlrT3/Q9tJnAdXdAyybLrNhNXpCpEGS7Cn9NzsWa
IToMG9T0aDWskajPslvWpyu573eZmalmA+MCs8MTciY5b7iBYwfn7iqc6bwt5gy0GirA0ssZIg4m
QECQyTFcl7cdP0v56CnzYSdseI7+hU3m/pCEgNAngVWH1as/PBx4IEkw4IgQSGyOklDcBYn16Vx/
GXedrafZ3+VzzTn/NiMxYkarXSnLprcf56txOb1JBX3EIpH44l44QMVP0jTu9ri0O1dEVco/NPyM
JKe5zpz54RKfyeNDsXeeeGa+jGqx55ON8Dai90lv5B2QXFDRaaXN7fI5Sy+TpXzKQBhMQuVho37j
jpfEN0bu49nUupvEZvcrF9R5Xu0ONsH0Ue0yuGs1CKK7vtqiRKrnhyTCcMoBrsXZf25nuaMaF+sI
8u5xxEWo8vPxBt/InM7z97wbXwDSeQ2x3Rw6tCvMYJp0dgqiY1qLMZDq8X5S0c1m4QSJ98Wiz+Il
wUUuS2s6STIhqjpFyFTy3DoOqoiIVyDJHqMv9fZQSA+Ehs8cfnsb5GmYv+seLpL8tKyvvDq912Ky
pYKEvYCJLEBet8tLjxke28mPcp6V180Cd3f8cOzU2TMS2mcq+Pai7jIw/P2GIrRrQ8cjua7H3e9l
c/P6mT2tXCRySbHh87NFIUj0N522PMdoEdu0vt2/1usMzCXQwu038UAfQIRI8HK4NXp09nw8TUPw
37Q3k24wrj51wiTJaBGUVxq6ocG3TV9vlJTamcMkVraG2uB1fGnOuO3CAIB1lNeA97q8eV/1phA8
Ls3j04lsS78HBQ57WZktpY6tpat0AMWn/kfqVGTagY0PZCRiVZ1+OKBicY8x4nMKc3S3Bm9tjYBL
H4OFqvK94OPZeUNtZeu/XtZQryTQ0WxkeZX7tV0bZVzfaT7aL/ox7DbbgmLrChRDR+ZFUyQcmYYU
HIKi4lhNE56vD57mP4gRXPSSUPglz3BUZ+z/c7vo4UVfq59wpW2o/VJRW2nSN9br3pS2eE3e0W2/
Qq75LM9NN3adz5+95+KDzGbw0Qd/M8NajWxpMyyVqZH3FHAAOA3busEJHMvqljxLv6ocxv2SKNgL
3ZgLTz+Wxsr7Fbic9jERyp+UHLYdaF2i1DATZDoRbd+xA6lmQtUyXqrTOsZYjxu8xhKv5Dtut8YG
Z2wJyfDvseNDvAIJLhvklDTLl5mZacF2kXSw/7Wi7xUSB/9kBM1wHcxLGgqwFkmyUmx/ERWKQ22/
hHryBGrSOqiNWjy3hK/4JDaXnzwS0Iz1w8I4GrAwl19Ji85e9XFAZOh0qGwjvXUjqYXlC7RTQBgL
Ihv/FFjNA0v1Yy3Nr2cUPxO7avGWwNaxqYyshCJLIKtN0rO/03Pes0FAuzbY5DU4zMYrXaB4i971
fBlX1UoXYtZJnxerr7Z5rK47wyc30UO1808dBbOHuqY8Fxhp9F3vFT+FuNeBdcIsnYGbnY1rUQ5g
Mtg2owT+VC3QmqUnYpabO1bKpaEPVX+vWYas8Nk9AXKHOztRrvpHuGvp3fNcjmP9SSLP3CoB+3IY
g05udEi7xcJwR2Xoy6PQb3vL4mAqEkMmrD5mVY/m00Ah8xg88MTTlCBrNMYluvMJtYuuwnrYz81Y
DoL0jYcfLdB/LVQjRot2vmGIcOwQrdybj9SrQmul5VHU7GKdrPUDmn4GLG8z4bKXrGODgLZ82PGE
AsRyaK8xnXmK1rQ3kf1g6GIN7OJ/hfuh364AR+5GSg5Os98E3Q2MWm9O+JAwTMT7DJzPmHNYiPPt
2EQlYnJY7ale+phnHcBUSXayw805enfAiq2O0qAnXQfOUJbF76TOABJiDmffnqjG/1B8gqhfADS4
7lQRnXOSDr4HPFqKn1hZHmJBEUc+iKDworbhjOIG61jXujIeBjmZ9R9Nzux9n1KpnpeAPRoOYZ3K
hTff7grsz4Z3oTBGOVcuEnvu7lkpbNQi8feQDbj5OHfa+FlbO/F7ivWoUYJaWKivnF1TczUar7D1
FUxT4XX6ZhYq/woEsCCaf9URIRDtxCl/Q7HI/+FLVZLvkUBS9uJgRfqdqLRlLSJXm0yCNazhFKoG
wEofJMWXkY2poBAbWVPwWBlOVuQ1v1ZCnJsP6yHCtuBqjZXrBU6EgETtDGOAYqTt82W8HnAsRKKY
WRiB/BqTTlpXM5MJ6lc2C5+BLXFEC2k4tz+uw2j//7gys6K39MwaAQ+G7e2Eo6gC8bziDi3twV1o
QbrbsHuZSkWg0rrG/8NKQXDl36QoxnENz64lTUcLoAhBluD64AniND1L2/25mW3SzchCthNWUrwN
RdgIHcR3haZmSpX0Nq8rRpeWnZOepoPUh1krHgUHB2vNRo9u4ZuIfatiH0Ng380zlxIWBz4JxbjT
td3plS3RcNeck1ZuHPFk2V2Fgu0a8DPuRjjWGePf9iU6s3sZCUap9ltsp/9AVH6JObywGkl3EnJe
StdCujjpIT0Eh6XKCAmfwmGS0x6zLs8o0baEKToggbFSVcZM80uFCP5LX3VrlJN1xr6XV6fasFfX
HGF+/6eYt+BodkzyN+TzP3SOY0rBoWpk8UAgfVDQHkFIS8wcuWQah7C3NMW4A0858jL8g79rqEMs
pvKdZheq07TOx0v+NqJtx2uW6gTP3zL1HlxMaPPeJaNNFw3s/RftvPqVYKn5Pz9KVLt4ZCH4XFW6
6S22NiBJPQkBvvOh9nMLkaNxkL1kjBhgYeyXWYvW8JsIdZ1yAV7fNk/KpLA0FyRxT3JaaUT5r/4R
3pMYZw97ZA2owqzkOrBzIVwmgTRYuce1w0RHmgeRfV/OJE6jlbOconienGn6r55bzhAy+UgyAs6b
S8a7vKk8TWej88ap5X29oOFb3f8i6ZGxLeql26oVLeej4VAxtPLlV4bUXcLFzHLfiHUuyxam2Og/
VPFSGe2G5CgwY+MezYf0ZChWfH4Rq/xkBuaOMvQlbFrgDL3mAmiNqeh8pz56bgRcRvlqXT9Ly9PZ
Gti0UkzU0avVxwTIsZ/PzYdauLNm0ocQ0cSQn+X66Gb3pTH3ZkAAPHSvej2dmJLoPVPASddYY+/e
fpDnrEvA2uri3+XM63ZSsqcjlqlJCchC5APZ3eN6pfCu4TevTbUMsbELRCr08GsckTGyYWIEFAZO
f/O+T/b9so4KPuB1a+M7T954wpHas8xc48Wiuh6TtaK4SrYVVRgJqi4kKebg2CnjQVt5yEI0dIP7
QKLQN4XPCXWE38/tq+WhQSZB5KgFi6Tdsu1aPotpos8bxpduobitIvDK75L1XVv7svzZ65nMke4s
rNzx4RoGSQSlNq622WkptO3qMHm6VVy3ZhG7vjEsn8C2PEwm7z+ywhuS3mpaZQok+A6ZkAm4Vu01
b5Y8MDfwiuUNIpJ8rBvutnRIqrN3b4FnFEnPKsdW9j2PCNdgDR8EdrDv/1MxFFyqRoqArJjoLlEN
IMmVmKtPMCK4v6OL7euSKVJmH2+nrLD5ZakgMu7130FlpEVWOkyu+DoTMLJilQdVHcFBrbXi7EKH
yQLEXn2VRc4ghdi9DnyHTSOgfnarJzYASHj3W4UwhdlFvPUSXpli1kO/3P+3JdDhRIQ5YQGhSfRz
P/Frssvn/rbsMhwHM01tDKbc1E+bLGVlJkHAf32YvHZitMcE08fJ1MjmHRYB+oEHe2WTv/Tgt4JC
7H0Z4lWCiXzfderWWzEvTvnXjlfavnaa++w3HrdEBfQfHEds0tV/8uugm3xzEGuViopKwzK2kqk9
a1TTaOg9JtttZGcZAc2PUGEfdp2t23lgEC/eNlcKNM3UFPEIb97oZ1DQzswFDSaTjskJivBsoSm7
8FT3IgU39/OWC1TL4Atrw+W5crCJYxSYCwCndlswQxDH4HQgjAognoVjW5X9MLyy2MsoaXI2pdiE
UEzC5HDUhC9ygkpdlOwZNBDPXq0JRATQk+xBc+CBASpsyOvN7Tl+g+EIOaxjvGUStq5gJew6z7jz
A5GuAhqdZjTcdi/LbDiBPpJ4kdg7hIrDVl9bwmmZpJXxzqV9sZifUqzRmsjjH7GJYkk1SSSsodJM
G4W31IFkxsf1UIjgKRNEofqWSoRVGnUHQZDAxVMcV9oI3kBTMjKx9fcJMAePgrNZwJnyemDSbOhV
bhZl1i5fhYwPBiSag5oIeEdaeBcs9unaoyFOHDI19uVTh+ajfTcgHnw1oM2BGkRa2ZjrEX8gvAiI
T9dphCcv/5FDA4t9udZoTKpbd7CgPdD4HhExbV6srube3fSBRL4mthUjJjf9Rifejl2kHkgtJSHQ
hoDXoftMhvVDG9xltB4pM9a+YbCQZX5slDR2s+6SVvm4HE8ZIciEBVaIJzouyzr8wl+z4A1TAhbB
JcVNzx4a8A19bLYcr54qmSgbKI8pKPOqGVgLE3dYVmZ+vm29cx5mQXQmiNcsYeENqGH3Iz0Fqh7c
q9K+aABeGgaqzwQOWEgjjNi/W7byNeNZEWbDjloIstJsGNRuiMjtkHkUV8E0qQj+Cm9/LJa9hRdn
qFN2QGBMBHnMIQCOzkffKnG1VacDwoVhLWKfq/qgSpXEl7doK79B/dM/cypy9wfBQY8V34BGtB5p
/COMwetz4YC0wgnfcJ1/NXIeO3ktCr0T6yNObNsXvvlzoyEwkOTtETWFW9M7iwHoe+u5Pahho3Jp
hnZ7woPQoPBJ17wAQH/UfnZ0Z30Q1Ugm0K2wUKJyza5sg7yh3pDnmGnLtvOdu4Ws2XI/NtoiyTxu
7IeUF2DEo4S9ng9EWfxFivO9mS+ZPIhQSrhV9OfrvsvK44EQ/u4PZH14/psyYX4n055CityZhkCf
P0hlY/VEOYUeMznFCPoOmZjk3n6ZzP/KvkvQ+pG9iJkA5gA5dHPzASLC0D/f9A1TjE7AI42jPV3J
yCXa77vJBsmP6K/CND/GgcoqnTIzmcXk9OYudw71dx8dXPXlgeCCrU6+g+XgKr1m8kR6pg9QNvZj
vVAfClzMWyYZfl2twKGrEFc7vDbj+Ll6Fcp3Wf0Wjc7bUZt249BW1NxFH/UvxkgvNcUXb1F2wp6a
Es2zDzGCIkV3XZy1XEUOB1iYxf1krIZHo9bVCfGOcw4OuZfk8W2LJhvshy7vg1olyAEF/U4YB4Yy
s/oFb4w/uZ3G0bdFNc7v+SnuZSaBZT20kLfVFarc65Kdyp4BgrSlaAE3oAQw7Ns357k5d5+cQe2J
rnikk6L1ZflS7idgmK4gcCDgdXdZCMsP1k41E74ux8rc7wLPwJ5VbuBhAPJJ5xEoEwv90X1DaJKY
JG6WY/DQj6Kd/I2W83IwEVF1dqJyP89tSYL64mhY/cTaK6IyntuFfD8GZZURMazsSsAQbUyrxMP9
bH+6/UJtmvJre6wdMISkCViYNtHfEoLiw/SsFhILPCe8y6uJ8RnWqRy2ZbWgBcdYxttS3iDlgwl7
UZLByArFVo/mB96JY2WuJoxr3GzOnoTKVRWG1flnKoxFoom7FZeosBKiizsTSCLKNZKNsxJNXqSj
KRjX+a9miJu0CWJCaV9g7J8UcDm8DvjVjaERWgXy8sSX3QqdLeBu2AieIPCeINRvlMAowdPcYP1v
ZRubSp6jjRZa9BxCAxQRtLeNSeSoi1+FD3zFlKRuA1/+H+j07iLeLUlNNULBz59AL6kK6t/AZhmA
hxRRzHoC8rRbbl0TqZgH5Js43GIYw+WKdl2fo+dv5Jia5OXT1R/0IeCve+mOAws2nw3JOwIX41UG
Py5NriISK9wQh507rnMF+b2d7SIdt7yVz94p+slHhwjPDTGXBiZvWmSwlJLVuRj4240Rm+VfdkwH
Gl4Q+ZoKlCxeCLaFH7FK4neTUjc9vUcMOdzy+M46LI8UaHLsM1uLrdY+U5Pyw7p7J+O8YE1GqmpO
qmjLExmfp2CrIToDo3NZkfsfwYtPJSVqx9IJPP44Amtn1dD/OLNDW95zo7ViB0eqNljiJB0QsIl8
B1qh1tFmt64WTdw/1GPev0FF0Icc+PpNhDU/1MN2NgjRVKTqM19EpSWXoblOQZCIdjFZ9WJMNfI4
LGNLiFJnzETmm0VSnZLTdudaKrCfzktfl11IsYa6haAM7keoHye0CfSetvPppp9WkqzvembrB9Ri
66eLBg3pyfpXjYJDM8Ly22CxTsaQ4dcK0l3dgObwG5P2Q4NbmAtSIGCW6KLnpQHefyD/415cAM4J
309x/AAbJiKxNaCdvh4nEkW99ZOW4jt2nhWlqEpI6KEo9L+OgNOkkWufxb2Gl0yOmVyiJpf3TwVc
mu0sHc2NBFMvvbuPMOFIi5Rb6mP3zn1LnqRC9lpy74oSVMPqrHq6xxu/meuSIhu/O98HtLDCh7Ps
dDLW39uvvNCxm5rTmpMW1KeEakAct12qPcQiM7QvmU7OUT9OBQgbKnF2JNBsae/TEq+M7HZcKSMj
CjbFoeY7NeqjjMlNiz+dVOSD9tKovX7OZg0uB2XTsM+tADmvLMZu6C0vLjMHTXR6ky4U9/QRJCRe
DOAZSQjgoyoXrxfFW77PyeSGCQeLEKtMS0qTsSLnticb9GMMvK5in1AKAo16MJulIZxBiP/sYI3K
HI0GpZ0O9G3g77tQswhZN6KIv0ydyWhLqXtB1vdTaQzPS9kY/SKjRxlDWJXSLwaU9mq+H9nHAzNi
0tdunwX7YqL0ywl+luUZ6nuYztsLayuwDAj7ft1ZWp1TNAv2E8kO4NUFkMTyqi5Z/PqFhKdILalQ
OTLqtzni60W21UpEmBrwaz4rzCndxrLObQPeTpeOx5M/3+u6/TygpoKvdM9rzsFyAEsxyAmFS44A
YIA0PlJ0S0qfKehgufjpNk32DcenSrpHcpOgI2TQShFJsNHe4jdnS21PD7kBgy0XtIetM6eeX0Pg
0j9jTY9VjBKr0hnANsedSd1zuEoBRyVnnZL8EGsjyAVCGG0yWqCaYPWjB6zq5/ymGrmo+CBkwzpH
UacgjGMPRXXN9wK9xQXeG73eaUMLHzo79mUwcV1L8uyms9JAKEc5wN4FUBSkvNFT2pOt8VT2n7VH
BDbNTKIUjBzBblXEj2/L8pF3yjjyOlqrJyyMT3ReiR1pI5hJgOPgftfKmSedbVByI+kshSarXZGx
FOTtlqCEJN7bQMZ6M6Ev+5a/XjUOH06kUmthIIOpfgwjpQ3dIoN8cKiFPeWwyprnT5afBCZxSVbQ
tp8fka+ZtDaKNFLGE/K2076ImE2qM8FvDB0kLqOrH9oFTRFPvDwOI802fzVEEycSlDLlCaUb9TSD
twUjrfKnQ2q/ysAm5jk+PyxJHRC1B41kTqd83sEzEwEfXFlEsWh4qCUXNMzGWjF3H6MFRaEc6S6R
Wfby9Xj2g2WWy2+FnKoSSXME0XaMjbURbykql6AcXzo+OGnTa8DHKjIVqqFJYvEMgBJ4Fk75SicI
VL1z88010Uzgrncm4Wx6YhjcNRctSpyzsTTkBm6b7ZnbE21E/fUAxOtm7vSvQa+tLJlrOGp4MD9u
0lKZGvlJNa2kqWPUmNl1/KdE85oYXu3bYlv/AgQvn80ZeD92AP1pOf8j/qPN6LdCtQG3+Fw8OiGv
jb+Sn+7S1/EbOmeaXTtePsHeyO4GljsCP3mgTEtS58757AhJZsrQorFlovl50AAxg474hCESdon/
JR6jZOA1s+7GVY+IFbwlNy2MwseA4b9zUOGQevy6XG5ogTKWzEKNty8ikoz4UjviSFpv1JSDfW6a
Dm6HwpAHc/YIZfPA7/RHxajtM76LeeOIf5CJTT1DiSz9mmSmSrk4MMEO6s5kLya366kQbg9iuqH+
HzckqQGykrIyOlQQsjERtDcL/i6U21G1zFwqtHxUCt4gKq6j7TtLUW1hmNuYzsdlL4ISzUw3rTi4
ENw35kIRIgjqbwbDYzOiySKdjWm5GtQpKr2qJFmwSP/DZosIYcMT7RyHlqxYT+zwdtgipk9r5u/V
pbZwtlNP73bTAyfVVa4yOWL9CqHBPkTjwkLZBOLo1Hv+1tZIdvNn+JrXvLVyg/KOsbzoi8QgB3wU
FxyfNeMDcgQzqbXaulsBO8aafgMXXI+0hoAStHVS0XV6tpHGpvwIMtr3vYO7GZa4W1MBIqWImSCF
UP4fhPgLAwj0r0B33vOxsrNNKJtlYLRX4aFPm3rT2XEkW5CojpNkBhXGup1nZ5DmAdmDVesBWpHQ
4/LZ2zYXWiGRQJlqVjPlc/yAtDeuWXtWA6Jc0Y1tBN6/8SeakvVGK0Ig07oBRBCoCTApQf0OweAy
giUQcTmQWjhqJsvkZFeGGpp4JkDJbFDtOVTqUf8X7NJisuT04gmjB9NJqYP5g37TnBtK4NSQnRxq
o6S0YO9l0xOeQp2ppGeMTcuoN2Mq0uNz4HUysHhFxus2BrjvZI5JCyVba1JthIhmsqdA2IBHQoX/
vIv8rTi56Uj8LQUz33Lx9tKNW1sjXaYeP8Neq88yr0ZcgCL59isFqP7OuElOCjsg+Chh1PjFftFm
Q1Iwqz4n5NZwbPP4HtBJCohZVViNMUabnBkoDrtptcrhv1N8O166d+t/eTevLHk4RxllOFfepAdc
ut7SZaoCUgqV4PKGmMw6ZA2ZCKF4PdMT5xEY8ifBEN1JkVMWNHkEhZE3EbHZObxu6g5iDXx4Qmtl
/9HfVIftyG1okXmWZQ2yZqKJIHjusyU6sXWMvZh7kTbLZrhbCop5lk0hsjb9yEG7yK+lWVxJe+9I
2yMLJWtT/6s6+7QyBT8WcM8hMtEiNx1uFePJoIrYRgJN/sNb5YI9k+FJQ1jvgg8PqrdAviQkjJ5i
+xzQsO22rwNlD2zEp3FUp0KjzdBfqkacATVcURxGFHyjG9xWb7eOPAZ5VsMku7z6V0TtFh25+tZy
iT0+DocIwFqtNmfuBAw0tquyl92UuL1XaS3krjws4tt/HY3eW+n5aeb3f/h3nizUI8j0fSEEUrTI
+Xj2Qj0xi7M06xTiFsiyvV5frc5ziXQNB/d89pP6aztA61tVsDtihJOTirvIFulbex80J1w6NlzI
oKPs2SPTlhPSDa3r0rN00iSFpZrkQL3A1wWKCuAuI/dA6s6zywd4STHujU+7sSna0UO4T3upgBgl
CZHGNNsfIidngiZoF5rUTyoLTnP0AXOj6/nt7gQuvHBtVVzxOkjkbuADsAO1AGUi0AS+kuz9liXo
wnkN52OTrp0kYoF7d52qe9csUhSneL+3e0cRg8KwEJwTHXOUSoBEzLz0lbB2NefOKs9prpFLMBHq
YdhuYyhhRdoo+QIIPIIITS42AjQtnJcYF1g26okgKB5WgWnoAwcLaJ7jMlsHQUnq9CtJ5nQR/M/Q
hCBXAzr3CNEy/FZVmIMrwFFIOjLIcbRPNWJZcWtbE9R+x95MeBHtkse+3kzmnRaY9gJPOqkGxuFs
Dm88L95pWJdRD0S35fJW/APauljWxkY5pXBrrpIbntQkk4J9bqyjFNxB55M8ytIxbTt9oNa/3Uka
xsEQ884+bLrO1/oBCkKZJ4ImCp7DuUcdF9+pVCexkYBUNOZKway8oWRHuSoRofH4/i3C3a+kJYYL
dAb0s13en/P0PVJpOAyLCLVjTQPdiop76n6LZAMbG4GIxH+2vkRVJPbxHDGe0nYB+p7wYurFGdJP
cBgbhXDydHP72MNqZ5GxGVjICSa4ST3BklcNfxUi3LqO1n3ntenfOEOn+EDINjD6LdL3ZYRIQdpM
kiplMgqgzAzJ3Py0JSyt2nEkvmt5eh2bEXexscbbdumR3eDfY8f6/zl7EXb5kDKLg/AfuS2wyrRL
g6M64lE8wGe7VzPxRRPP/hRDziZxjZKkTKtuHbTFC0eriUXzqEI3dFoGEaYoS5fDgVe5Xu25ZLip
H1GtyYXJQ9zIWPHRvMTB0kbKCQAbovJ7+yHSTAvKqdzgvM2RE36+olDDey6QdLJzYbYtaLkymkLo
ayXP0/EqN45k7MLpz5EYBBQzcXBogVrGqNuqlqXnlxzi+PxhdNRA0zNCgmcX/jA7aDoImB6ep2LQ
ATewsMPD9GG+vDhQ4sozk09qS6y/YUk5Qs0bG9KKBwzoHq1nXWJWt9MTa4k3rSaGtto4zLI9eSCP
ufa7/wZpV1R8iIy36VAHpUN8pqXVd7eQ/fiHGhf2rULVIzkjh0o6w8mHAC1x/38vrxoWUukxBJh2
CPTIanQAan6DROHuueH5CQSbQT5dhcJK/+bhiBpUvsu6c1SB4O45k67pgWmFq4m7HxgG7GzMF9xk
4zyML7MMs78z7TTilJL7+wNGopyO0inqjQKnvD+F3TDe8cD0JOGEnPaMSn08q7VBMlx4rWO5agpL
lJ9tyCS1w0jBG4SB/7BP/1ffxDzMSElzJl96I8tiGtk6VI/F1ZWQQRsdWDdE4x7MADiOh+ChA4Vt
KEgr0PhSikMLeIF6SkRxmIzOiJUufQpKo+PDZkFw6Md8tVBBL5k8AvdSqXUxyjCLfQaeWGwRn/AU
t+e44vMs88yffCzDlNhZScrNH/F0HUS0T+e1PJrfqoj7Ibl47yWePk/HAZI6hxsYrp0Ju/9NUUVd
pguvmK8V1IEFhqsl3mpMO+Nk4+XKwJgPjeVWcF1JucUhSlTcugzbdDtVK8+04vM5xIviqagBnmVH
wgjRCB/ZfF8wOTHb2JkPA6R/ctoptGSVuVVxJsap+QosKidk+aobcytu/5irXRoYoAfkO1Fmn9zk
cZdJaGXmsEGsFMnBVOQE3RUES+I7zMDx7aMAee3wgMs8Cel4UUfPhqRx6MUinS+uhYEhlShsfrgf
R/1EZTws+u6Qk5+dL3eKZqTnZlBK23b5gLDER8dddvBFWrGxqo3UfVendVPH8zn+0j0+Yzcb70VP
7utTtBN8URGjfufTIeDuFdOsYKmCkfrUD1fPzT4lorsv4Lhg+BI1K77y39E5vd9AzfzB1lHXTEnl
EHqnl5iHjpOMq4HoKUm5CCZZ+Lqt+s8/YBZMamWHcC/VqwzqEvmPR1EBRcG6U7zfLaNtH1PniW3k
p3fb+dR06suLcBinMD/KByam3Sfn2SMljhrlGEN1/3dlb3S+1GRg3HtT00UP+czG2Kic+igvkZX9
m6tIDOSa8KsIIGoF84Yvw7Fp+siqtrAmLb/M8PQhwnh6O6svYH5ifcr56Lui6qKGCJK8Pz3FlO5f
nMgPCme7tyWzN0d79hfogxMjgPcXfCO2v7i2uVyPh1csFwwcgUnAuGbx9CU5FMReyQ1HzN7C1iBc
3XX4bonrBREw5q4lDio1ep6g8IPeVeAqEX8e9D3VgGxDgE5zW575H/Zroz/EDfwqvRq6+luSCPGr
lF+cgQgz4GI2TGNCyLI+1F7HMAprzL9sr9GXcsY+tDTGY+8sqFhCPB1t6PMNAKd9LYipRjpNDdSs
deWMvKcm+NJG+Q/3EnTHVsv1safzdi8PgjrYH+YfCHlidfFztCkmOcRPjAaUei/6x0yLy+m2oMQT
bPpcaJqWkEEJNff9eU1QWgNnJKdiWrkFY0h2ccRvgk9LjRxunyER4NjW8T2LVN9hbkD1AfxMtwyJ
pF0zO2d2ACqtYC+nScsslvtdg4b11GCrldVmsQHThHDPdS3H0XT9DDXGXhP8OgJ5g58qACFGqRA1
vxA08pU2UUFCv7A13/tmN21N0QCi/Bs5Q/oDWDcm42ibYXkD/lbQsI7U788QQSvnApR0LaPj0jUn
xAWbQYamdSh/iGwT/C9dAWNR1npuf6lQFgXkjw/tAHKvMkqAD85/ZmUYatSos530g/LAjK2+ATX7
XJ25mFw5ZRQV2EcRQagJZOWHtlluJGicvqFULQswwLu033tbnKk/fzEoVqpcSJb3b1e5fnAfzXxd
W+AiWWKiGlrmk6Ul35trKMdQ7LDOOiut9TQuYubJLb7n+Cm2oIrtigOUnTrFTGj1KQGnnfEOgO82
UIPd4aGQbxdBYwR15IjcBVSUF8lNKyi0jpL7S4iLk+U/ZpvykilnkcdV5BZ8m8NO4+KFjOeyHcC/
SDn2uEMUBCsSXdzVncCtflZpF1cLn1lPl0+2pYxRSyZ5QaxLbJCmi9m7ni785rY3spaqjNGA+FpE
LQ0oD+1UNAyuwUmhSO/bjNmCwp0c54waEvonThKtvsLRI1gdu+q0S/CR0I4JXr8WliFsoW1RvzHa
2IdWe3/YO/Tkxbmm1AR8QaOTfR4ESptiZLbsY1sIqf4Ifyf5CHLLUbeJ1NF+LbuNr7mn9cd5qZTa
PUK6q5eEKlAPKS49CK+V38oz1miuVBCJDlUwRgAc3lts0MVRsqDEJy62hZKDEmcen6OGCozOIUG+
r/2yAeuVBfp1onXWiADNuZCliLOVPDdKRXt7PtCpkz+HcTDpHi+JtMREajTJvXyqrzeNePt4YMBs
J/15XXmS1PidBgGadmnxa2M6B1Z1Yp3fI35nWHo60OIA+kNGR7XdhlDL2dJps8gqpNqaH8if4Qh6
rGCVsEE+NAQDogIVc1l6BenmB742e8SVzbxCPJnySd6Ll7gETwB5MDTaq2bVI2Bs+JR5xZEO6ubq
G9AaHz3Fx2SzSCjfmdjwkB2vR4ryvl5ZN9ihl7BxIiyQQKnvAWOaMMP9WJ4DI8xAPOE1AEdixbo3
TZQHGmkacJ8CMMj1LYGTgfmOE4FrZRkL7jkE0HyuQ1qbOIOvFxYEfFQ32pMoYVCU+ogzAtY7PNeG
ONxh+7EM2XBvdLTn0PpWwp0bIhcR3POd3932oTzsITVAV8BaYMhNqI/mWUWoE/JNiPcdVCFnAySA
k5rriqpRGhyFZl+xCLzgKksZTH2JUF1T3j/tBfsbctQG2UCZ2VUFrQVbj/7fqjYPkJ4WThcaTyGo
AgD2udO9GM5u+Mk+OApnbw3wk/i6L+n5Q+PBVT/VV9FC3yrp14ikSvnZlwoDic+8AONMMTcuHZoo
+Zcq49+AWZZQRcPXy9hF/4MhOAJbtq2LLgxdwuo+fY2py1QmdfiHS2eTRPm9JDd06yDmboDeT7hc
I4V1MtEoFOk7XJ99KPK8/tICxwWMHmwivvk4CsjUh3UsoxRlX9FcIZPfTT9x6q3t3Crww7LN1w7E
BoquQYMVXNQzDzgs4TZfLbwqKbh1q588YA7qZWYmV/P2VpfMK0LGvrCeUre+SPiG/UJ/Bm3hH2qG
tKrhvWAoec6ndwKBlXdIn1SzwhguPiDm2oDVoz2iEzlor7c37PtseJ2mQDYe116h9v4KV0/+HJ+M
aBOUmU+twqnd44XGICIr/hHhP6gIWe05WIO/UE1isoF3JnAQYwvMUd7oVDuuRjAWqqrG2shgtc3W
au+kPVvTDqbttsUZwDeQ+JDOqIAwjX3YoflB+GE9VMW7lPtFQfDlmGN/X3vegGmzPN9MFMkKjfM/
VDJSXp3++ln6C/38CG1fkTEJoVaLcqSKUjfB1re+CESl5g6utoRDjk8wZ235ZT4ehB451cz7CmX9
NZ/th6PfLnJ9KyJAujWaGdt+xq0Fhl8/Yds79k39ick10Nq7oCIpCjV+9gNYb1uT+YI99uNnZSST
vvrsXbzcYKCv+JH+8lsuNAdZpMjuDxqhyL5gt+sB5vSKy08IUKuSba/tKyry+RAjchgRYmbVUdbV
19NvNiJkCsrvBjAwqJicYGWm79Fu1sohB2GWRyxmxzDe39CDOLtwZOT9bMvETMObmrxMRyTN+7kE
8ZT2htE4G1SXRw/8O4Mivr7YiC5JJwX+M4eUaMxdScrH0MmWN7aTDPqnCpFS8ccCDXjA8Iw+T7lK
La1kMeFwaiDbLhbOVbhQXHKmfm7VauZjXGahEDLyNLMXtfNugxVxl5/k1iUYFGIuvrpnzBUbjbZa
uyeJPzCNYxGvCLfuw/A18nzhOUihFMNj2lxS0JgpgfkZJHzJCnXTSjwGcvBxU7nK7WdMt5xa1uYt
MXZsmY6eNnAWX6NfehBHWp9cPcqPZiyPYc6QhQrCBYtJv1ODAajC2JvhqCfbP6FEBHl3qXHDOcAw
FXYqLXShuU12dYoOpMUIocNdA14tZz73V0yY0M4LMYDhGKtHRk99IOpJKi0DsfiVkBY+CufhxWyY
sCAlB1oy91flI+mhHOdV3++/MiEZZE1QO9+w+IxHfpmSQpfYxehuyFyMcBmAiTwjaDp7+8ii2SyS
tMh56SONf/2IS+wTkHVY+Xa1c9TiIArQExns+1j6mxuaHanjNje6SONIEE8Gxe+Sp0rP/CyglCAb
aUIT2650KetTScUucje1CTFsbdMjHE2yCDwKRR35tzU95ow6rb5zz4IUK9h5R1a2w63FecPmqdFL
7CAo/2TzecughCyfy9x0KntMhqPtI5ajyQuJuwsV/kaha9V7fjy5nigFu96GUH4gMIBwiKrvZOs1
T7pJ95/u6XN0IGFMy/eQLShbhPdJia5abHuckXblWwMtC2SZWVEkXZGRu8I2YbJTNQhz4QnV8gvy
QWfnnYdg2tzpmslMHzjonZtmOwvzK+SbLFMlPC6s7bFtJhltXb0GI3/jAm1E4PF6lfvg2SPzxe4F
UZGKZv1rVzEGYv45oztGS9Qayn7jfhNPOJv5FLU5B+4K6a/PqeNOAE7V8g4zMUpYN+PT4RaFzSrY
x82g/0D9SXYYT7F2sVV1eHLAP+1yWdl6UvadQYAGXA9o+bv9vkdbMKiG4s/MAlW23n/4/lWoZfj5
ARug1kDck0uz0VQrYVP3kKerrmVmlhv25Rr2Tcb5NtoH1pm96nzYv9yvjL3FEl1BDSjYlH6yxoiw
SNzdLq6c3mB42XUV9pYQHNOZnoQDcSc49lAabw7ooTFAEVn4T+aHXJsn69lHzTSpXU76A8wNpTW+
HnLO2gQQ+2dBOXVmMjP9Fg+LP5DHrqtO4OkiSRIgnvS+z2QGEsQ0LzmaLck8un+PYKIlsl9o13r0
XuuxD1+TwCf4RX53tGgGnulo5G+ZkajP+UwWJyBqq8Pi6OOz4sUxY52OULlpslLYtPvQmSiUGKNJ
Lhfx3xKwEmOeLrHFq/DegC86HwaxbiFZsFof9LPFiayKpBKuOaxox11ML2CySNYA6j134vTzPqmK
rPhpdfPlfx1wC9obPwmuSPF7L/0/F3SRYlpOLQIlVn1cFDdc1O6XOf5CG2sj1nZ2C5uM/nbgPczd
qzrZo8XFsVr/ckeI5TA+fSUrPmQwgaJTlzOeJ5Kgc2vAvoYsmsuWhvQyokz7bD1nVttBtP5lFsUV
s5zFFmRiBxjnm1B1Dw/1XYl3qKkO6Cv9fxXPKFt8GH1XI4Ca5t0ubCHfQZnH01+K1DWno67k3R0h
1Ps5wQgKR5X5BKDRxvrUFZtGR/NjaeXsoTsBNi379iN13o8K9Y2EcNJ3UXRnyr5LuC40z3+8UsFr
CE0r1AXJJsNM5RjX0e2CBxco0ddVfAL3qG0wgVOx1ccYcYEL9Ep2yDNLIOtNOXh0G6q4aUxJKnI1
tw85ko0skKL1YUTH1Sa6DYJ+QI+cyor7xBBUlzY2Co+f2UUOMLZbPDW237yf71VRzSzpssK2wcE/
WWxiHv/hNRhqFEmhuCb21n+KdxG5W1xITaOU/rY4q5GibW2ngz2bqroPhHJL0NJlqRY5BDHbnxNJ
13bu4H2tiIzf2NVlLqevCCnkKsF6v0sfS2w+c4en5pzYWB9/8ZVVLpiaePh70WGa4Pez9s7WaVb+
gq14YjSFNDTs2GD03DMqMslCx0DIjS/tAcl10oWMLYkPJE79+DetpXR3e+VE/NqNbk1Wh2F6Wqqy
s8AgHzaFcVMWA9y1jC9jamMcWfJHh0vEbL8lm3fGmZfi7PjwLIRbcWTiSQHBdJuAd4RmVkzrgAjL
hRaKMHuvzFifzrFr1TVBD73IBJYv2+pocNPWt1QBQLyTlssQ0I8iiPf4pXtC1YTEx3Mg0BC257/5
a/uz3qdSi1PXQw2RCv/kkXyFPnhQvvXkWnX+0wUruLfEmcpjQ35m9D2i6+C09hyXnNqA0P3Sas19
1HUyxzEDpfW4RIstG0pkoL4uuHQxcDgZD7hTzELANl7javvZHi59APfoRdhwkMs2r2WjfeQhGI6M
tfw7jVI4Pugmv8ei+B2CfgxKFtSSdg23WpxHdSZm/lubHyl0ZKQgJapqFNMPK8iUtoDwL/9Tqp3V
9Xnwpgu+IN2q+604O5Xa/vJFooLrzvK8x0ec+lmI8szauloVtsOlcdi0nNrq4+wlg8uOHJv9BW+J
vq5ukiLAx4bV8buBhRKq3A/G3Y+N46uSuYBQZwZQjXtwggcOgoeP887GyxI1Asqy7EbUNpzmDH13
ka+76QaAZ4m7Tor+P5f6Xo0TGRcE+/1lRc3Bg79tpMPlSOMcUblQhZQzeEWlH9BOU8H9QVG1BZcJ
cR0SmRi9gp9Z9fF3azotmvLcHblhGFhBuVLQ1EYFpsQZBXrCavnbdmXip5M57Yp5M0nRu6rHENgj
YYJdSBNiA2Mbte8LW16kcpfcwO7PTDAtX6L/+8o+biWtzI+4fXD1nBny+0lQYsO8XRK9ODMwOnaE
AH6UmR4pyHJBAH4VywCrYMYlnzfwhpMLItZxMiek5uL/pTW6Cwqj08SeXwgQKP6RH1lD8ZVwLl14
0ua1hGSGN0uNV8YRCuewvudyu1COfWc9eCZfN0nq/DBY2kRJ2bVLkqaK3YW/WwseaUsUXMbFdqW2
txF1+nsRJwusmxMhxlWVqKGt2mUbt9jwSKXOZiG950VsmYU2Enty1MuIhMjkQo/A8OQRID/6E5Zl
SwzPkki2D3tSu2nj+9HoKgnsAwbVr3HTl56Ysx8qNpYVtwcfGWXs2y5HbR9yJee2n+Ek7Adb1K3W
qhV4fPR2x7iwspyoTzJDvu+Qsi2prVJOya2gPMiezUeWvfKEvaKtGoqUjR/ZkjtyxzxwQoV4G9Vq
2bIuIZc17cmi55NRSL8x6FWTApc1jrVqMvGzo7/g49zsXXny2cLQOU2uw+/fydt0Hx5z8+a3Yvu7
o3UWba0mmeJNiLInvQyD6xu+HADxie6xSu+b3SH+TaUqwRwb9fomW/TlkE+CTrabLaQ4zBFtjwan
e6XQ3sQotsY2IeSBeCGU0kwq5etm7tyC0eF1Lcypc54Ns5KjDLt+fQl3L1S+IzQyChT4Io2nDHCR
WTtHp5bxbYv6y3yfWhYZcdte7IfyTeXs4w9rCQi7Jbb4dQQaNuvxbMLljGvvK85nOq17cmIUpI2/
CcdSXUoCtNHg9uBgNnVZkHHwfwMTxy6us4GXRI/WHhhXN2wyj3TremaxSIdlogATRTblByzCW5w6
HlfIR4VNiN6KljHmmtMdBkpnvPNqevSBXuZByNG7gp9Q/GkSdGj5Mv/POYAWts93rwu+8rF4+68P
lNsSyYEjPIWTrVDSYATLrsEc8UWFklpZ2KuBH8P5kaF/obaeRR4VmegqBuUlDjqTvWDNOBcNmF4X
KEvy75uFClayPd5KXHGZf4LGBYLZ/trRB5bQaJiSxAcKGZzfgwDqLr4BGYfu8i+VDzWiZs+tHkfC
TwaRE8+ZYTec58eSV8zSeVx6w/SY60ZnD/iOd0YjQE9pMUGTwMy2IYvh6BUVEbRSc7LuDkxHkRRf
x480ue/A0LJffBQLqeNslT1UooWjWry+cIhy3VcQJtQ4dTYOEwr5fuft+77jkJKSTEZ7dBfCDx6u
uo+9oUm+i0pxMRESDEYsYxECQguXDpseqBRzVJzbwjG3Cqj1LbepbBVYC8so1b6OIEtk8XSMWPVJ
uvByjs9QuYGTY1DH8VNZMSO19gnq/vqTmhdFRlip6H3GWFu24oPlMyQmT1RjQ/hhQ2vNnbT9CGks
FQcaQIaFQvjvassC6KtltjDOcmHZsPw4wayN3sBPBskpNG3OaEw6IWv/gOHactDi4B7zxdH/Y41n
5tkf5bz1jyEEDyaA0Mo2AhWOKNacTdNfXybbHAnhRTz2hjAFOkyZpgm+tD6PYA688wPkO1kfOin9
8GccGxdRbbjQPV08OxOOqUKnJ08RShyWXP5MdSnA4OsCkmAxoZ+IT+ohIc18vDpKE1cIg9eFUys8
giAiNaJs9Yvafj4JRN6jA9RhQ0ijdapVpf4QKzHx5dJ7XucycoDg7S5uLft45POIreVw4/bWSM+U
I0Y4Bz3b3fAZkxNZNOqOeesiyADG9HhMtwkknPtzWezXLAUQgENrqLVGE5/0oFFT3dRDVrSHQp2K
zMpwsHTfCZ1QMtIH9Cq8NEBV8sBvcW4zgeFZmqGzAevVlzDxIFWe1nDFbTo1OjaazJQdCAbDDSfX
2iEs3MKVpIpL4zR++uFFl5WQnRBjhvj/MUm/UbfF3wdgwkNyf0czu0lA1u802IsDF4CmiRnC49aQ
GDL5j1uZuTutvYdSA6FpROmruDxPBeDHvIu56Csnc/kdD9dILmN5rb4rV212e8P8gs/eXU3cvSrk
CaGV5v8K7po8aXSrvEsHy9JVZWzG1efuhivSWpDNH1nAcXHFrNVJjX+vCxxgP5z+EZ2c3BfVQvfP
7Ly08IVkwW8uAZhPp+dUe4MFCLmFQlg5YaswJDYzzctGbwjl/0PrdsnM5xDzFjeXJNINgG6ZbLXt
HhwGCw1VxkusOSUfsM1Lk/fLqYMwp+sZIc5R9lOAUwhF4XPEjz5hADFhjazVBW+JXHDXI3RRlVtQ
7JnoNDOUywkrpIeZ5MPX7XbrLOs6G22nze5cbjwowJtZ26/rDfojoI707/IeAQrhJvWsnveHa7+h
mg1lx0Gwv/02mUjdLapFU6GK4/v/jqQAjup0hGERVfeuHYV9h7TWRJWuhwX24H/NnLo/XwFkzlAd
tymlx2iqCmOtWrwqJISuq4mjZy58O4CTtPnFAVmdFawyTRedoTwHZhn87bDnkh5QHQ/as0XN5pQL
AibTpH6EmuiDiQR4rCgIhGghoCtPXYwXj/TscD9XPz5W6bEQ8+jV2blY27k1jpHvBqCNG2l7Obti
RZnAwVIje7CgYf0bWxj4V75YsTVhXfB/eDyY+8zN71CWA0SMjLA+1oGsUwHFnJg40RYDa04l6npU
+k4yiBjPe4xcGrDthDD9WZL4AV7uTSpR4DvZkdVVrRa1ngXwrwyqztT012Yjw8C2gr3F7VEt/VC6
EGEg45nCtHsAUV59l0T3zTYw7rJ9ZzbchoqNsJGx8BOYpauaYcToSeDTjs7OFXm13azMKcWLPxlt
iggQukdfXh/3V2wM3PdpAuWxn5+By6juwrW1ES1F2D7xgx2NSRXbcmxe2JldYWIhggI/J/XxwZ1d
V7gMYaIDqT8T0q1k7AKLj/5hxmXIlVLF5mF5NkM3UQSOoLzD/ioBAg+V/mNrB+v3cUYMSx23VunF
/h4AFPBOlXgP08CbLnPtT0dHZ9QxrmbcS6+05ByIOWO++9sW6nJgknffydBjEbtC04edTOgjUzLS
nh5TmSwCrs90DTRT3TBvUQ6kYRyDpyqfWGPPR9frSvBpbBB+OSbTjMyBXhXbhbZU6qdAymVpwUHv
rObdA3qBmHySusD9h0Rcuz/scoP+nOwLCZdEmuOp2oJ4Z4BoQLPxfqkgT0JrM8MX6isqAw1b3j8H
0qjokwvcloe+2m+9WsoRgT8mdL9/UdDiZiuNG7Pbal+EkDpM+N54oeD8BPWgdOZQ7oeQHJv0E6EK
H/+BhwED0BbyJmKmtcLzmt3eSbV1nk+sQxGJXL1swx3N+/pXoaWenTi19Ro+ijrsqWJsl/oxEUma
Q1Mb7o9iqKNYaqik7cQFA8RmiE9C7wIdtmosS8PYX6xIpGC4UD8t3fKUv/n5Dno3mKZdRzVFjk4W
pgcq6IK9rK2tvrZYpgq6ubEY3XdVqHeGNOaPMr/6ksedVO0jzUthBM7N7e8ykZVIuEclDroum44P
8GEG5mQcMaIQRjQ8ILEi/P6tkS4EkjCfar1VmEgnzAvC03UrAHIZzD3Lj1gH58lzpITZJdyxCvm3
IGzz5AwAruNo7xcsrJtZM2iOJfLHe/5JeKSguIODwkWobK8Xt8aVNFqoog260X9tRZ4mmo0aczXl
7oJ5RnzTfn2c033zzRPnxVcmn23b4DhdzwdSkpGLlO/kmaJwgaipiKMposAIxycsP2a6BIUVV0Gc
vfusLDh6GNmKF3vUQPnaC/adnMvjzJV9eHYSv7IznY+TbdDDnWM4vJB68xUIhrPSZPhIsjU4HhXR
jtGvWGL68BEMROsrJHfO+NfSr0v956AjoQ6NW7KKFIbRBkXy8DrgSiEhd2VnTilEss0eoZk/S3nK
E56wYU6nmJRJh51n/nzZvgMJt6JpP70WzDUC15/kgAp3OaiCKzteKLJR471qEGiX13u+S4E5PFIV
D6UtXVO0GWpdjibQoimBn0kK9x2204fDFYF4PAaIGhSoH16Mgfw40ndq2jdIquyOTuoagV8KUozB
CrvxNxIHQKDgCcKtmAY74CttNNjY8j61nCA0OVnTCDAu0neBsldl3uXzdGXHyIp/BXo9sUUlRJGX
sDj/jCOw7e8JSCoj7fCcv/kZErcp6SMDrrE9JarEY+6EqqpbKslczRMvXx+Nr/ho/MkcOTnbv0UW
FzWYW40xgoN7VXHGJN6x8zaQP0mtGHVwD/9xDoMWBzXU1WpVQmzTZyxNBHaizzxmtCMIBpBaVcBG
GIQbWFoo+WyavQT4Z+M9XNpXdoY+72eb+DMbpXFNQ9FXnM2dIPnezjNlIu5nXNdZe5WoQ/mvWajz
oALq6XGNHhtFZoPgt+KmxvVhMUwpArrbHWfxUbClFwF4McqwDbwHtblvKRncRGk+nKomJpmNqbBV
sm4ooXkO9ZPAXFidrgz4fg/C6XttrPVMuxyIIEaT2FaD0RrFXBNiQ8Jw2jLU8jvDtrLJ8w9UaZzH
H3aWYQ4rva5OiK7Bo3atuscohumOSV6E+R1dnsF8Bg49IsRFIIbOugQrAYvIQ8D44Jxe/8Ps4pBE
UwI8remLr1USSshV//aH0Ed5NzYAA9zqCan+aQ04gthapMAX/xZuospB1G6c1SvqIKRQAja/zsrF
TfHB1waZYutugXJg4m2YAjVuoByXzfV8C/5NKb05gQ5DlPQ8yBXuADSAovs7+WmQCHV6YEGWC59z
s/idI9DwrL00NM3oh89PdHfUy8QTKBKlCIpSJVCkIWgErvjFFAUD903gFhuTTOx+UoPza8kEoXIC
5FxiR8yx0s11TS1yd6ERohEGfMA6gMFkFLERzikUEx959zjm1w==
`protect end_protected
