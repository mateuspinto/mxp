`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
0USWSUGxovGsyBJteYpEoQ7nuWc4VDtTv9gqYi420dyTlnSIxQuWoAxJIaL1FgHxekuf+0TlsNBz
vyJJgqc5dMY+yXJ+5Icns9kLEJ0zHIyJtFMSnuG9hSfhpSm//DktgOozmGi44mBHZGO01jHpZqhm
oZ2eUefKSEcuI83TMmH7PLe3Ph+Hfa+NRv/Y9f8uhZyl8CvzU64wIY5mLhCzS+aVR+7ch9v30aeb
HTj7eNp1sAb6LP+xWJPg7fB14qnYyu4zKAZtkwj18N/HZXtlV2xGekY9rxPtmY0SZE70vwNYdjK4
1wIZ4dr47SG0ZxnMH0+QTmukQQG4CTARsuNfRmgxd0AW3/0u7gQB8qP6ZgU7HQVyGHw4y5doTtHU
IxK5thZTrYOuYp6nkVuadTQayZAs8D4cTzi60Q6t4mc47qMh65YS7CgVcYmr9iJBDQ9DWFQKrogk
uFtdbqpUNNHGEW2lW7S7Gmt6hdxw1f+NM78UHcZ4Otrh/799R0+d/bg5jn/DVGhW+y9/JGecV1Gz
HuFi8d9RuHrfyFe71r85RR5tQxHZPVGAZlUVLUPmQfDq3lkdofWuJJuOouQj648S9fucJbbshNVv
o6B5af5KvxXvBUyJefYVQHLI6hCfZZ7ytGM5y6G9vDdCpNuOS/m7rH0/OYsk/dnvn0syUPf0E30Z
sENdWOk5o/EH9g4FtT0oTj4A5JI2olV4vI48fOczVK0YdtyJzhiFkyNHLP4ZLqulXplhoIiNHPwK
Gr2eQwC+kIHJJN4i1UuBYN76KZby39nXQNhSsv7EfYV+bw0Gc8EsIizZWFn1cSJSVk9TK6+4Himy
W0U3nmZjORdjdlEOEX0FDGU5oaF5bU+OcQwd6DqDFlKcRUN43cYRhO2BrF5rHAZb5Fkdwu3hLt8I
YiuTKoiuhcV0JfURDjjHalA6eawS4i371Q0ac5vnOSyuTztoVKPvFf72B7nRSagAXp/AOaRiH0ms
pjkuCSwAtoZt7tIaPZNtscHygUHHGvoMgK3VHb8z/yK4Hol/YcwsjSx2MvJqauhjjdD6SGvvsW9G
N20pipEdFCk49sUcAhTXmN+sLh8A6oLf8ojhL+KJ9N8uYUmY2tTKsYl6dGsoEHe5b659z/8dNq3w
2md0/uXCehhWlDtBIh2LouVAl4QAPx/UKpMZMouyPtBixLRFvo9wZYiUMCuFM2FDkkeentv0p3EX
QRMQ5rmF2cygM1Wq/DCEU68ylRTPZ0jdAstTCI1VI2/5nyNGVS9ZY2t4yzsij0bwaUoEVpXFo2ug
8C/KeWwnLC8VuBclp9iHwt0fx6w4xodzhMf3cTTioRPK5ygVJi66nHp3C5Vfu9UY8hC040NqSUdd
c7uC6WeZAL3QmqWuN813FJ0jNhRRez/M3HqYrwRIuTfUD1dSNZC1Rke/kAV33fBUjxlWrnEBEqPL
u0tEAd/lIFbcT9XS3hyyEuzG1I+gnBHVm2my+UOburJCvd0pGPK1u/x/tyihjWxca/4xRtP7Decf
M10r1zCcTO8cC+Ekghwz9EMyzcAd8k4X9iF6NC8PW7SJStESZdaGh9cAPrNpcflTOgA5GOGw34Bi
GHg6by38ZbnS6YO179UyWt19iciCynFSyqBw3EY+l4LlF+K0V3nnOO1GatRlSao5mzQhbJPeyZPe
8XGKoqfVtA4b9uzTyDRW+7h59Dxj87MgSk1o5q9VTh73erEi9vjK3eqzIm6WBTSgtk/oR5tkUDZJ
otgtrEdXTFhOkD7XHvES/kHI59BR0lekkTAcuVgpatOTVPe/e6HliX3/jyqPXG7jbT8dXGJ2541i
REDe3wc7U9yVHbLwlZFOH6wZfbrVHJhKnDLfkV1M1FC8PG1vlefH4yCXv9pCzBDw2oedGLm/jn+3
gRZtcXpG1EwyGwvzphiBOAIg9vI+lD8acR7TMqpPr7GiJTN0Tnkh7Dxctpf7cKsskjYwlg4FVx5Y
u3Th8EjHkSgsNlUv2d/CMCV53itIrqsI91fG444+r7mDRon/AtqGLaQnXTT9ENTlsLdW9Bozv5it
ZJHLdMQrTbJTXmJOqNIPqsv23YL2WLejnyHiPcz5K6x60RP33erJ3iABMWeK
`protect end_protected
