`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
oLZRe52EIDUmWFgloP0nSEDfAFhj3dP77eiCDDoDaYzW/YPc2Q4aKa3cK2c3YNKAtXWlmO0yDz3C
BRHQZAzH39zqdE7Zc++F5eSQjJOj8dU1gIRrZqcS+5lBIzCJl5UVBhWYs89mujaRFF9Pc8xRkYdY
iiuet3cCBdHOBXN5+bDuF0IsaFx/fsIa++BEBjm3Q2ldCLAlNwUPsstuMbCGww+Slk+P+rPXS3wd
kZc1dbhZDxzVUHO+2kNfeE53SKeR25vgab588AROb1ZzLhTq1i4M5tT6+KH5dvYUNBVS6BGZ4gAG
5RE3IdYX/ROEIbCOp/R+M3MdvhLkD7BlT2dutQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="C49YPskNBHacWpxdU0ezhofbvHl8gc+4ck92dUPI+no="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13856)
`protect data_block
eQB/MiKJ54p4q5Vl23kUBmm114qaftkm7FH7qhehRtR4anGkD/4OipBEjIuPWD4dX0wpwf8KnliJ
Fn0jUOAQZDuYzgvNfX5dLRdEl1U2MmuQOT4+0+IVpF8aTFFNQMMnb6hMnEt+Up+k3ZyuIsjNFTq/
lpJ8cijQw9RS6iy7ufvkZPxRKTGWGC6DaSUsE6W+PxdFr4RoV9/NzXPqAx35kRBeDK2jYJXGGHSA
P6eOtldQIsJywGP2wdMjNvnmFK486tacF2YCPWqWgtH0DCsX3p/r0hTxhaNICT2AvmWnmqvg1DPt
f9mFjl57tShJ+aSE+sfImMNs41ezat0qcV2fRXyld4TdzlxExD22eXtQjrR8vcBNqsbqX4iilnC6
HGYX/1UXgYgWXlGB1yMc/kk9XIUtxuATfCD5pPDSNm54EZaSm/MlXUQsK/o1SCHsljD6dOPcJ1zP
L335YoI7Io54yAEwQXdukh4cjJV8+O8tcWkH33Uk9QgUsC70fjHSJWTd4a7QNOheVwwY2onaMdtv
Khp5xDJJMVKoKhtUG38glmBgvehH8TUcFSIHyyc3XRru0d634iSR0gh6BiZ3v9U4DlRwi7XDA4Aj
88xC9V2NWR3MQvkSFcee/IgdPrHP9j3Sub4cHjwNVWePwLkQYeY7Iq89fEAk8c/pSOKbKT+7c9kh
pKcnKseJpwgGE9Tejxs33ovtJUkYrWwTUiUiuELbwR0O6tjS31Cq8qCC4IJL3unXZekE48zyB3Hl
Le+OOK1atA3/PGw60O7OfrOFz6XS3vl6w1MPDrDdznL0pesU5gruDJsbdbAoS4hZrwwYSPXKT49L
w4bGVnqiXWguXlyKzwga848mEpvtzCgXXbg0a2Gx1LJBsOGQiXhIHDxcPezGj9YV07o4kvmfgfo8
Fq9rGwXxfYL9HtxHQcRSFcmMP1S6+zufunwbK+x69xhVNqkh97Xk1v+IRVxQ1VxQJztGtgkXGH/j
8yzYZ9YtNY4N/uZE4+mARVqBxQv8BJwwVm3z4FeTIeWHmOCWpAhXkwlyJ4HfjDv+lW4plXaqG0CI
weFz6gNTN4AaWqTRlMrI2q5bROh1qkVo4CYb9FhXiZtqib+dyLpWPtjYAdQYMRCOLy4i2Gu0K9Ij
b4u5Fm4mQMkMwGb8qGHI7izGVbR1t+VcQcNfXtmInLQw8xLZzLJFg+3vb73a0rdb17oGMC0HEkl4
j3S65j3kKY4M9sqx9JnTNqRjZuzeD1M7OxX5CwOckbq8SmvGiw1OjUMme9LCoB7i5X8Vf/EOMKFQ
Hr8QwtKq7QjrZ2fWd5Vctrg2U5JebZ7fvgzi8G98kTm52ax8P57QwfLkG3NrLjWia6ucF+aq0XRz
bRiZv/tx+LFYpipHVlEjigUZ8xhggT4oEWqSwePS6a1sUk9qNfn2LynxaD+PsRJJvCeGs4nOnlgL
jiXLWG4a77toalO5hQwX/zOU5aBHcr+W1mDNsxxIztxKRDnh/T0KHmldbaN7mzLYIEY93+peGHbZ
9L6gN7aPmZ+x27WvPRlgiyt8T6/MdEJ6dqXv9CJ8W47SCL4nu0uktXn76vSmfH9wgCzvvUV/m4gm
zjheQ6/voJ1nPNdha9XN1vN5CW8/ZYeiyuAyWUVYSBmqEiOjxssMoTD57PqZPrCqfkL3cXv9hEOs
efVOlGPgaFMtUQbVKqSZfkg2/AWjHLuY59oYSiAXU81Eei3qREeiEz+q+6FEdrvGvttwTAx+G8Bb
mVMFoamQuo3ruHJ8Xy1CLH0unJFQhOe5lcUkwLLOy5linMfom5eFwZK91kVCDiVMPAFLe4B5dqzx
J6ExKmyBsEbgZJ0WKmyaicQpUEhpDyKG2kBfLCdjGubjTLJGrQYDsdr+XZElsai6TkoeVceX5hQ+
kiVQsAR20pfF4f3qgsHLLQ6OqFgk/lHXrlgN9+23Rlf88vftPsSyinALiC7Yl3ihJ3r2M4Cgo1QL
F7dUdvxKOFLyfnqelmrAynFxsxVBFv/IVSqBC8hzfgyOpaoXbOFmDEUJ56Z9WCi8zgky+jU8mVTw
8RckJBMIJVHU7fsamKLpV93xnQKBe1D4008SlSwqPVgr9fdPQtFykH6pOh7USNoXk+rD1i2u2XPS
V+B93kXHbS4HJn8Ycb4qwCVYhRQpuuGl1w1ZLuUj2JN9k05b/6cxxDc5kynraQuLVx/Ae7+ZH6Ay
wwyj5sc8sBgyfSWKxtZfw6UqYBvjSHt+tv9YZamQo/6+jKHzvFlaDu4wV9kgWBB4clyYlf7zZYcp
+EXH0wNENpoD6dUxlZf3NLOWhe9N7llBfyiHRCvT0umOzxKOANUfTN+/OJrUskqaRHfHmHOdt9WZ
u/qo0BsHAkY3KaGpwwtuc83GRHamktBCcHThqrYmRj0Ou5zOmECpCiChGrxcgXJB65qO1i7qdnPX
sLAOAK16/hp875wJhLXjb6VB9q2XtNlrztXBLuqXW2Jexdz5IlHkF3T2nDaZIsV1SkAKOQ1N0vQs
4cmOYH+ccN+ejsg5PmaQA/kTmQTyRhXs5zqf2qPE+nNaLBNNaH9XBYVPFAhEoPFINvaYJ0xmxlGE
YP/M5HSLs5e981CDIISsk8MD9QEgy+ne6B6hST1D6gfG8/hioByt40x12jKIINBaifVOf2OZsl3D
0ghr1Brcz2Csf22XQ0pOkVRpbPo/Oj+As9GiEKlFPKZZMR7ZoZ4Ik/Rg4lSTl68ctx90sUXBz3ot
brrWSzq5P/5IpkK4KR7j9r0lBLQNAQoSKfmiKLtQF2FhtCn/M4efASP+PQuP7VlmgJpy/i9I1dIk
O2Avz2qnxtAe+kxyzClTB7oTUwaqDDKUL1hKzhyn/MP9Fp1HCTFcaNs+UUTG/dS6uawqwsMydag3
MAYaP735PSSJxmXTpsxdRSTWMPotmvBOi5BrEKpZPXJnSHt8vtu48GnJuJ7NYW78Lqba1BPgtwPi
2d4maLDve5KDQ7sqV8vlIhmw+oOXpM79dmPxnWKKOiopOTL4yMA7P70CkkCwMrnA2IW0ujsF4irD
b0lUzy36Z/P0nNc8S1I5Um9sq+guJ+kjtDkLTA/1wKo13eNYK4qhC9F6ngF+c25RAizuoj+iV6+F
qFD4wQqEZvliV301yuuIoEWuATPTeW355nkgzmyd/nOVc3jMwlafh6jucVgm/6PCtwqUuR9Cvike
YiBDZoa/C3byuz+KCJqOAgD8RxqPgn3+MlYn4zBTqUTEzQPizclkEKoRQb8WSBncxvPQu0w9R6qu
IdpkXvEEem0g0FLQMj3vtDA1vHc5lyL7nx2hihOQFMn8+45caoflmEayeEsvqNJ5e1zSatUrlvmr
l+5oDTgZed67bQhR3LGnjwBNCu6HEIQZ9E/mf6sWmidsC1mZn7m23nUexNBuiqpxURqzqO6B5EPK
1PLasOsNrmO8eoVQe/Ksw2H/m8r3lQYVKPTpc1LQgIsNQVAmrc2AsJXukb1l9sXxe/FaCfecp+hw
bseBWYe+IeYzlE12SnoxpGi5HJgEHwLbS0h0TcdnBAhE7pPSjVZjOALi/yyjml11Wzswi0Z/UumA
oaTZihTgpbGo2LCnrJFf7cs1xD5vJuVWR+Ia0bq0Izl5Mip2lfDxLQ2YfnbC/nrJa2FQKQLJV5Vv
JCePRC2ta5p986o6wh6x7p2L2l8iayVTXDbj0anhpRFG9Ew+d/g2X/u0R1rp7jfeZ69BetW+JZrN
wClQH+izVBrAyal6HlckpDCT4dSqxXFsBO+F4tQuD0gV/PShVFnRFzZxnZV7k52d5UjluOJH54tW
mlMiSXAFxwB9AFWS7liSnsqE06XfokwUKZIJn7/ggmearRZ/kZPDTW5fcLQpeivmCUL93VVVdn4A
z4H8Q52gyfL3HwJ4KBXw4vvJoowYEkJlJysFcKtBGMlt1KuITPdRM/OJhFe8X04VT1nY0X1lJtew
Nr94di6sAYHXefSJq7tcsx5aj0f4THdZdSayqdDGXBg+K5da+e5ViwCv1H46/3YqSQZGdMwmImhB
D6u3OJj4s49AcgsT81Q0jyyd9MuLVCFnhEAob1fhztwX/W45ZmoeDYEXjJeKSUuG0qKkHxvuJ+Ro
OaYaxjinBEH8ELK2Vv22WfkV+N3l8me+kqcX2x43YboLx2WZL4L+5qHFDAuzOXltenpWudJtQ0aW
N09OqhNAjA6ZAqfF5Lb/N75wNN96l7lii+/EFgm3M8s6404TgFV0toANeRu3okSc/qBGZr4ahYQV
ceYWLGKNPZJAxAjlW2F2/0Xz65TI+9ZrAjafB6PiMsRAoyvatWIegJnnAXqLx3U/NaJs4NoATdry
a0PFvIyfTOD3Agw3406Qvylam/G7w/NiHh/jmxl3XMxK/8JKQhLe30LUq7mKRvpOp5Fo5aalfsUu
N4t6W2qOHVECwm6Rz2q7btEtdnRcM5mJjvjNwdbC37UOB6KtPsK7Jndm6J4MqYnN5wjKGZ2OU/WG
C/Z+OfPgqWUr6I4wXcDVMnRHtxoFmkkVtdxCd8n3tweV4PjbkgeKhzbczY+RFyPkyk5f6ti6ESMx
WTKeG2ENnG5z5YtzRP9M037GGnO2ZDXxwZjZku1lE4ITWCxwNzVyu1rn91x7lIr/sgJyZdc8qxPc
QUDBJ82w9DhvdOiiiQO/OfrCRCI/XesMDSsL7JUiHSvZRl+wU2W/ZXG0AAYx00h5X4pVhM7qwimi
7XTvZz73yZLCspDVQMCHS9Yx1Sbk8ExaOk6u3IxMR9ilHnaOeFv2YP2Tk7gkN7sm1q/ivfOEA3UT
dx0/4YloDU4NpiVA3nDfh1tex684U5v3bffw+20lO8Fd7H7sMzzOxMTFvOOfHaUl3IL2WDacdFb3
Y7O/mVif4/uyRI99T4LLAh/4l8cwKlSfJ0VhHBcRR0MUJe9aS+wKWdw9Yxlh7cTv7WlwXpD59a2K
+K7SJh0Kw/S514Lx/PLJeGdipO86Hpn+BT7eDORkex3s12ubfFteVI6zqY1fx4NvwAZQGbujIt7T
DOT1CncibBWghYvXL52O4x+X7hdbsyLtRaIPL6Go/6PPovwYi0Nt8Y5esHFsj8HP8uioNKf8joe2
d4HSa5gs3oy6rKkr5jKUIgagddNSuWTYCkJrItiqKF6SF+LBj3f1I9il5w983Dsa4tLBPo1z2b4/
82L9S4Xep6qMgXToRYwSk9hVudt9DNYfSZeF+n8xyMX+LnncSyeX1DdkxiLhbKBJjVXOCaUyv9w6
rBMPvL2rujZdzIK4hedW2vxxSH64XbqpnIwDFwYF0eV98FKl+teZHlI5jmMVDul3iuz2fRQCAuJc
mtlmfW08oys/XCBra1eznSsHgdR48R+6Ogm8g4gqvl8VQNa9xaNhTaen3VVr8D58BMk5NyeZwlUm
5/nFL/7+P1frIw7LrKrwuinW4Rf3d5tgp6HotTExXk4bbqWte6Vkws8NJUcAXnWsxBwNvFR0d/a7
WGUIjGsVjIrkQ7KTL95GUhDxGiRPH8cMobz2aHfApUVACbft5pyB4czxH2xrjJ7FC2zFtPk/bZeK
QwnrH1ODnJ1xVglCWzP/2nvlXTOZDxiiz1HUglmuxsAxedl/GWg8Z78HNnOUkX+z9PjGUbY/phC4
4bfStiMdla2YNbDxWuMQ8BMbhfcSh9EhLWv9Zt4jH4+1SQiRDHGf/PG4VhqGhpt5C80emHS+BnLH
019V43HE1nQRYARQH5262Ln4ssa74QYho+EUqn6ewaiLbb9ek0gvXPkzGvJpXUo9zQY90RsW9sA0
PlzMnrE8WuHmd0ShuChAo6mnbo8FKFjWaOVNzP2WSJ0KOyVxQBVOv4afB3GcYXYB+/XJXTNDt92w
InriIBFHdg9yyqi84gZO0lhzp3ylqQl+1/LuQwZodj9hKDu6vLhPXyRS8hpnC8LmcYR96T8rqRRi
YXJ1Il6fjkCGVn0YOV7N2Z0cn7DuyRKLFLNg+zlsNoUnJuxAVWuOOMsvmQkIT7CxfJsTAW0lyT1b
vL91+39Tml4CVDwOzHk+AXn+nVYegD7SmTVYwAKNCi/Z5kJ19E+l2+8s2YEd6k6F532R+fBrF60m
TCfyQjlPMutS8zqHpD4f7e5vUXet+vutZB15U/L5/PNxvODsSFTXK+WyxvD6qFlL/1ruABkIbRJ0
Uwd+lYFT24UZOudUtIATRvefMlW4OpvRbytNgOTg783K1mhQrA0DK1vYk7z99KaI315BEVBrWf2T
l6V4ahr3NwE921d9mdaBFNi3V22ay3pSwMQpJdhBVs4X3ZKfbi9oN7UpcqRrtsuGPLqpVYLMQQpZ
Z+19aC5NqWMXBnLCbNCI8R8J4X3e9RvTQ1eJSCdqM+KwrFyJ78ApBCFrQCexJKdrjqzfli63Hum1
usPMe6yLhFlQ5tg4z+KqdgoS5iwwmsNf4vHAO9ZBW6AwQfp3UMD8GY/JLd40SPIqF9OJydXqnETp
VfbViga+Q5dy8qhhZsWcJpT9XLM15ixvYHRkRL5ueenDlSP0bRwpIhyoxawRxA172a74hSQcaF+G
dBWMPLJqbaZrQmV0ByXTo/eKhd3L2nvFe47WKYYhokm6jJez4dZj6fI2+HMqnrdKFPFEQYSrzdF0
gAtYTBHKhOC0spNnSiR4aDK6LSOwtF5rT69Y6TsLgLewCWHUJFA7Dyp5cOHWS+uVPl9au+qcnOIL
NSblKSMaUq1EYSXN11K9nt5cFb9tOSixbJ0LMm/b8rrvGFc3Yqpd9W/dEsALjV0jfDiF2VMme19Y
czIkfYtKi2wyeHSLcZrKLMx8CIOrkcO3yEKY43gVN0/R64291bT/+ce3vSM4qpyPcAwd0W7S1dvv
1CWBZ5/Sb4CTEDUJoY99vb3qwWXm0CFYshS7vmc+lQ9YaTsRopYusx9Z9quQQX2VAaBPdS05Phvs
+DPoya0AFup7wvbnHV5Bi+QsIhiIznhBbIAjcqUo+lf82wb/HMhMiTtLxCC9g/Q45aFzaW4Tae0n
zTY7ONZtfsWu4WuCMbzvenaB8GytkqyW/NfUnpOCy5vJa+/B3zWgouSjuBxtLo2lw+fLb0WRpsaO
pXu6oIAgT5mQZa6QH58eHqlTaiThq+6PsoEHS9vpk8hyCbOzaFjjulnDAoN7G3NNGUXRF9fF9yGo
QBRgzwLA5uX4zCICNjUdIVInxXKDVQcrZHarJJnfSO0JjQYBHyAOK5L71F1B5JhiX0364LMfLX52
jRGCJA9H6Xt0R9TEotjjGRg6i2POkKoEWfXBFpDWLLt7foR/N6VPaGLLl0jk7K1yDUpE8gwH74jr
gH921uU8927yzKDai3Ov6glPPe9ESzukAyqzJoCU3twiudR7oIHOhfLtQtGBve1UUkd+38wdu2Yf
na+QNFiadisqcuKzbyh+xCfjvKAUiVrl/gXbKe6yGgSI1xa+J/9OFwlCme8W/9lwGSMdQzAK4Dzc
ia/vB2vWaxqeUyb568z5jJNsvz49qj/SESubV4+ynmiB/GSdipjycKtJlhTOI3sETf1QnJ+yalvS
r10sESz8KiN6ywQWz/0TwD704dfgAjcR3GZaCysmS+bnZ0mO9CzXGX8SNIzlUeqTlCStL9YUs3ET
n22CsxsXKBuZSKZV/PKNpehBfFAoI6OG7h2uNX5Itt5yBx6lCjFbc36LA40IojVFQTTFlLqnOMHZ
RQyD/Bvv5/QIGkuGxIDGfOwapfYQJYLZZHuijDG7txEGjea0cMQquDsjsT6Y0q+UTcty917YHqFL
CpIo4AlE1v+BfEk1+dLJSbfGm7igIOOEbP8ZjbAFX8ewvAzgAp3UvV49zaYvkKrQ4m48TcWDI3qM
VT9Tx8wKWRuBpQMOnVi9LzMzz2+kHTSYwJnOtgiZwFiVnyiv3DvuGjBDc/f9TZ3PAOEPgV8wFXZs
IoVreCLYsM3gIQIAHKoV9Ay1Y6RNQdhAlOxh+ns60db0QywZ4TpBjUVMdXR9gFcpSu9JdTqPSC9c
0jdwJlLnjEUDdCkOnefdKjhHRgwq6DkK5UO8FD3L3pFWBTy2qeSIRnBz02XlcnFSY4ObEJfkizue
0zLjfXXUVJGF/cziWFEznaj30nlneBYQxeRX/Jx35w35zemsdTo7FZqW11WUiDmZ8zi9ACoNExWU
3/IoANlYh12g6/nmA4r6/6nNBRbBxXizwWABFZd47FPXKcaGqVFQffAD9ut67eecr4WBc74Gz1WN
Tdfc+U+hByVYia1TlQ941TCLiPm+PF6uyWlOa7wW9/LFZAbo/f817b21gmBjmZuDBlRo5NFO28uQ
Y8XxfX25c/RfLI5JUvi0XKFnSgf8lZF2G6v45UYAFrdGLARb6dv7sc9Zw64bq4DEBjeIROD/puXX
tLFRJUyvCDqCaJf6p1oUrnVO9voQk8ifHt8BQEh8gYkf+A15FPHQ18ehl7gswrnNdfPmVb/2LcDh
aWlwIiqSHo1Qhmp5p1a8sTvn1SZXsqvrE8EE5wY8k/8WeQVbASHDkaudA+1sPBECu7/Ith82SrqS
CZ99B9EwRy0Au9K25c7WyyneEaQikamEka3DNsR/SJQsuceLvdEENAhH2/WGMzugFyR9H3kY19zZ
wkE3j8EliJfAOizwOL2CoFd8TwuhHeP1+eOvyDYb+5UgwUXpTQL916Xnet3A6AQCkX2ds+U35hNJ
Mg7GOJmJ7ersviWkUwo+LmepZBbVlD/zR/EEkf/HZ7WPtztna37CNAvpoAWwb5AvOunULrqLesRV
IUAEGMmHcXl/P9vADWj58OLuTIzWZahPEBQKHOpWVOSoDRnbHyEUGj16sFqUQd5/75a6ITC8rvMy
DXtUpAfHXYtuWqz8IuINMC40KOY9CI+iM7NhWatV5cQ1+IcT9AvRD6cJbQNWEXEWPw4U2ugweuDj
F3YdQWMNvrs6STRvpnxGVmGY4MAqV4PW3thQt07sgeffiHEGct2mr/siVViBmMrrWF6hSgcLvLQb
KRE/YbbeSi9s0gt/1FFTrXubmv+NWqWFLsDlxFOBPfqFGO8UHfvzsvevggTT9ijQLJ3UqYIzzoqp
F6BG35YqoKBdgfkdvjt2x2ZtVH6W/QDGSi6QI8Qs1TouHtFqmzVD5kuT8HshIX9/sCW4xLTPlTPt
6mlOegM3fA59u0yYiuqak3Cs2f4szFsisDorbFRqXkYfpzLqitxUCh91WdDWB0i8t0543uZJ0ojG
wEWIoDCA594oXqSQho9EyZV1BFCAf5tWp36IZ5+DVE+sMOUHIuQgo+iSTCtEWNjFYypt2deJXAU9
Hcv6T21yQJwjU6ZdPvT7HEg0bDhNDb0tRU/Dxa4QQgspLrUrFHG+iPzis4tYlIcGnJc0SB8ioiuu
7Brx8wPvghFgIRg0mJhVj16xpxbXImUCLWhQaVslMiD76XhmZKbD7ZunPib62OoCTspVRdYEF7TF
k6N9VSwzW55l55BskE314p3Tn3fCbw9RxKDplmxF3oQx2+SssVGtP9hoKhxCOOxVHizBZ1LWUDj6
1EImORBQeOsv6UG+LAXfrTfw49FJ6stWi62WyhO+obRajBXw+evhg6ZCKxcndRsFuY/6Wsrfs0bz
MdOE5/LAHH7yCCBRfg3ggzoKXfQ4ZRZDLzaLVSXTjpiMogf/vW/IfwczOQUBKfPIt7wygN2Lk5lj
WQ29kdqgu7NwxUWUBKHuDcw+i35DC5KZx95D62jISOjtruLUWYtSmrVPpmIcraj/O7jbkkZXvTYi
NxnAE3MzxQWRiUXtjRtoeXafEiPAcknusEXGD0bfgivOp1BP3K2a8FluZs1iLiUWfOtYYQEMtBFQ
KdOKPifs1R7CH8Jk8ra0idBRr1TC4kBhHI24CmoKnBOXUKdEr4kiU5bb5W7PBqwKLzatEzgx3mlZ
2jmDfN1Tl+z6gFUxWYCjbmNKD8AYQ0cQ2FxEred8Zq73KEFVWIs9lPoKn5Nvan8zGGm1Gck/Xsjp
rwlZyczoAo04H0SSvTV1r03T8BKhJI69uexEmOVrgYhbSaRIgJ2WBbxi4S4SyE+8/D9r8DwpUT/H
XUCN0t1womVbk6b6XbfsDhcT0UvwH6cy7rWl0mzsNbm+9mOxfXLqi6CCx/qU3INzcUzjxp/Bl2I9
x7zF5JiLOPPP6OTzDQ24AFmtfJ/DTIG3xwxbMOH5tBRXtI0CFhnygCsC069p59pj4kDb0fuPGrB6
bCYhrIgtnn2/nSLBC0Rv5ZOJPwuGd3QRBELLiHephiRDa0rZMWEaMQbT1dB24FZjqPqoIo3ILrJx
IRIoN6o00h5Djeq41Hn6DcrRoRywOZLHBPocvQdfUGzahRnO1yDNaDEY/RpG/tiCI0pTbOXi5u7K
ODnnS5b4ViCqGwf0bk0u6Mvk+syRUjCruhBh+Nyopht1L6XDCY7FH68Lxddx9VbnSqAtygQm3OEP
jrb9FsjlvHUDqwwMVyciZI3DzaXDr1rqN2ojngwl5RWBaBNB1XgJUgvlfucyFxk0ySWLOyvACZvf
CU6ypIi0u42zY1sOf2elRnzi7BRjAsULmojOq0OtIUSgxupD6ddHtXeBXy9M6F+bPmgNn0ESjFzB
nO/E4QiIjWByzufPYH7hgT+7S+6/FtO0pZzGqImC95QdyZuhbObKIKIvR6LZ0pZDzD+Lm+1IWZFo
ZB8JkQEKux77OoxbVxbGQ5QDdI/9D5P0fFGnBo9I5El9wiiZDPf5wqHWKE/wVzZCRNfpAMnM5HRX
nQ24K98c2sV1ZjT9dj3hb/+SGWI6oUhUdhd7LAnQJL9sXc5HfsHT3PzcDDsWCkJCRTWURqlLb79D
QmIZ875hBxKe5Py5vvR/4fAd+f3JRCsHX94zbn2JYEG/5bLqK3yNAWUBd3k0+fID+7HNfum+MA0h
Whzuu4tPijd1QaDqvVrI0orPTL1h4AyGP7lIQCNbtZuPiAlxteEn8FMHFE0k+dpELbPLsBAkMrlf
yRPtYI67KVVllFV7bP89mUw7CJ2dVVShC2B4j3n+7UQbPXmZOtaJ8sn1FJQhIC2aMxu5+PzTos65
8Uv3I8er80Ag5Hco3dMPcJZTFifpn1DQ7rdOVf11yFAyHbcgc21aInuFLYQaksRR745fJxNxcA68
9/FGZBI8Ho5iLpZhX5k9CYAI+2Fx/K3MduSuGjGWyi8F2lNkwcgz2WYcH9B72uoMCQeCRuuI9gZM
2nuif2fqavnlIRc8cqS+fYwPUFqtDq6Ph0IxMr2/uaZQkQFg+kmcdCiWIX4/Ci+sxCAzcqNJtCtm
PjSfJhDHzpE23iqTEN85C7rHpbuX4m6Q7N4kSu2TT5HtLLuNPDft+JZ88+H6xFTQMLBKtcf4K4jp
o80jfF0fWf2TTASU0u2UETC/a3E9sr/FinD9HYrHx26wyEeewH8aeK5JLiBikfS3vIOHw0N7meWd
e/s1JXeJep0W9veoYdo0jeLzJFXzTJoIDkJFXyT5zWGO86ia6inkzVvu56CoLukEro75rMa79Cv9
+pKwX5hQhWeXydGqwaab2J+46iuB4geFH+EeIe2aaZU9AlGl/n+eYxsbVsBfenRAZ1n4iBsDvgSy
GWyvWKWdyVnuNJnGsj/rtcDBkWq+n7GIsf6O7r08c/h5PwgKilYkeb9AP7OdbzJncOwqHtfSEpMu
/YLy31Lhwjawc2bbu3Ei8G3C2egaYwxaWqp8hPizYaEgVPkflGi0eSKaXXWPqw7wVVApjJmX7Fwr
N4QsSVs8zy8uXWnmY8Gw0MuoMK6aNobLYnagYOMHlgvhoPKDYFn+ZF+TPGe2jy2oErsokeJnTEb/
/MtaHHYYpsuEVrKmovZNp9XjhdGJACuvhfp9tm6kMqgQVLL3RJG12MI8GpFM4p35l87TpgJ1CURB
oRW5Lh3jNjOJvIhzxe+Xao+7sD/8XKrXFjlFVBhna5C3KSSjqilzWcLFdSiStNnNZcq2m2C5osa9
q4F/GuY6o5IL6DQFoMunvOsHelCmRm2SLn6a3C7d51uc+NJOEOmGy0nu8EVYuGpKYuXFGcNscRbO
3RYVgLAxTNb1y7vl2nrjW8OLY6/yVhDNfdVU34/WyoYsz+DKBQE7UaESQ5Yj6XoxbTIAMjX0g6+k
IvtkpoKFo03uhRVon22V/m+aXlrnCmko9UOfi+6Ugx+rJCAYtcFEShPhpaEWFR/gDFUAhXvNtkLE
oA1/Ukzes4ovGzqkq5j6fqV8BCcxuwrj3B+g0l6rfSH8xiq92A4WLP0M13YKad0worhC8oS2jUUP
xujIDomAN3YfWC3/GRoqu4avUko4QnTORMw8oMsBTPlCvNcYAxx9pc8mW0kn41PHIq2vF+hnkuz7
CK7obONaeG6AoJ7E+q/MLS4G4OjD1GDVBDbir7vJD+jnwxy7rqViwjyvNobNrBDCmSqceGigO75q
oU6Zb+yqX2WVVAvUZv3nYZhi5CSvuorgL2I3ZYN6DjkFEACTWGwBlLFCRyOk5n+C3387I9bIIn3M
N2yOwISDKN6fKk6zMxGm5rvmGQTPcpxsRCCqfuuOQ0d6ue3JJONdC2+sW/FoN9931K9ryTN24Gfo
QduKTYTIgtHnuZFhVjy1d6GyC14r93HfGdqo4FjaFX4033kI5Ikk3HOIglrZy3GH8kenwO1P1wFj
CfM/jhJRZQKJzM7jqfEMYAJ0f+Qz21n8QFVG+ArlSS9frc8yp2DkxNmwWBsm5rh8AvKAa3caY/s/
+30T1xdRUImB9lSvyrMYj/H5Ql9Mk7fGyF009F+OhozdkPOz9OktiC3heki6T1DGhBq/fRq459uv
kEdwIe0K2OcTWjR+m+IJmeKOGrG5yPZgngxRoImMKSsHXddiBTe5yt0/ESqZD0oqUSSSGKUQXMLt
lYjzpDqkwczGee1Ky92wBtDZpQA4lv4J/kKpxMjmqq7Znh81rZ3FPtO+FnfScxB5W0FR+RnKEw2m
4KpL0OcsPqNsQjf5RXC4n6ULBy6p3AdxTRdp1MOimcWrBrHZEcSNtv82g5/E/2I3rncc+ZGiBt0l
EPcWaaT0DP3K5hcxpKBn3rVpB4zhT/TK3TF0jvmS/yUjHX2Q5QL+vrrmB6cJOW7thoUSBvF3xOOp
EtFmpHb/Zg58m0toH4C9AEMOwhCvyK+bLAimnfOTrGvG90Vwz4NbCtR751iLCAft3YWfbwmQU92t
BPtmemVjqRyeMQi9dfS8FrD+P8Un9hh6xlyygQhazwjl2BokhQoeiWcWgPV5PISg+UzdT0h/lwh2
Xy/2AJbrGFipPm2Op5VQ6TAXyxFZycgEr8upsO7jtSo8DIRiQgOTFduLkh2NfaBC2HUTa/MKrnG3
sNo5W28KPlWc2Qwz4fG/DWGs0eWJqEVSH3+H5FWQ8QSuV9LskBHvkzBmACWwuLrgesZhA8fl9Ra3
04/mM+25l8DyvdKTROpnmefNt1RHbQfFz78Nr5dfnNJdV7gMd4OCHKN2UqNssaBvbBc2rj7bdbdW
maQ8djhRg33Zm0AcSQ0Yf6t7aSvgVloNX+a2A8rVJGHvaR1yP80zKidAQ2BruznXkMPqoHfh0MgL
JaVf0LDZheoiY0jbji6eU8V7KqfpLYi/MNDxQjjlvpBs+t5mD8vFisfnVrXayVs8pMNXjQUBIuu/
tftMyKhRanZ79uUITPYF1BVaxfhIhGiAGMjCweo8g/4gc0IcDkCtt6Zwa2DULPVBDPx6TnuLAdiU
cG/7zT1PUfs/cz/79bLuJ8vGol+QSkKYO95yeuU2TVK7C6p//zlJ9QHnl0RJ/XDsnPfSmu8FvX6a
fCSYP88EPvQ/TzAZzOhMRovWeov9JTzjtIRoxar2qEU1VFuJ30zNyqPJ7nmub9oCKCsYYJ8mMQak
MVCWVwvkU8p40XxjRAOHoVZ/iBWKnV6FdBqJkY+rD5udMgV0B0LLU3mojWaJciqkh/e8nfg0L8V5
QrHjkrkzBzT6U8UVXj6IJasF6FSAtBVoFSepXzx9hFt2qmfppdJqFOy8sAL3U1sHjWR8mDRVttku
nPCkdqv/OUOkJ5dgzAqVgtYkTNIRQsaqMC4619FO1+trHESHDyUu2hlleeNIACR7jAzyHUhxFS4F
IfeNcQPxUNTfvSucIFw/SEaL5ch0bT6vdNosh8FukG8srS0NQ4ODdC93xPsDh/1DhI4nO/UeBl7t
lgWLVYdnj3Iv28OoeDdOJ8s8rqe8qCZn/pS8UoYTFeHsnrNAvtc6tyNhFxAr5Zg+52i7VI/R3PwU
pMA4ycRaFgggwxIeHL8l+Gm46w5iW3ytIXpLaXOmnT0J89aYMOGt2sU+pJIAgIlh7yf3SE9kpmuI
6ugy5ZXHyQF7yOBF7gscTw3qvsW3jiDGb/tY438IlEERXn6nxq8rBSN0uJ6sbPAWebIZk1sOW1TM
/IfVlm7aWfnBYw7dmtHOeeMAXfkMCd6BYAkHgOO0v2JJIhuvfGm6GBr7sdrJmPhwbLlBfdqXB7AY
uC5mANXSb/3WxRu6tsivML9ZNi88YR9wYvUX2NOF+5UKv+a2dzIR6FCKqGgbDvxbjdPVKrNt2npo
QI2jYwkPCsHSrj2HFRqlNWrqWvA417+RA1o4hirrhgXyX/kTyuhuNni5dP8U51acCDCGdK5jqz2M
KehL899M8diFfcnsJ2/Ok2AiVNofe1MsNTfU+ZkdcBNLyPUNuW0a/sNwiK/y3Cz7tHh4JpkCiYb+
XlAAQW5NMeLm+FUkbXL+BBqhKHbzLgOHhEolwNTcN1PW+5SiFYBkjFnLM2vtrWbB4LEXkhG+ZSED
VtZbwmORJLeg4+mk06tZLdhuslXupTym7yzW+cMrDoitI1+puhKPaPQ1D4LbIax4VpwmJ3EfhMr8
di8ufrPPtspxbonDlvIGlj62pecmDrQM11B384GvvlNTAE2kXhFzrSLkRywmmSt5D92rhmHff5fm
JM7/yo9VWym46af/lvNJXWdz97TT66pequ35mmJvnpSTE1dTf4DLW3BoRz5FOuXtdNNH2HN675Mp
rNHuhC/cvLBDODNlbvJI98wph1bNBPNs4MZb7DugWmxTuCL0aHqfg7Pt6JYFyCkcuuilCbeOopO3
tZGLsNdMJvgu0IVxazpUjAPR2QZTdz/i9C6+kQaD8/49+IwHEvdLUyODjDDLJfDZQ4z5OeOtg9hF
yKAH//LtpCrH9bkZKc21vIqdtz4Rh/KyxH7rlTCrGQUjJn4zmo4rxDTLgjlDITkDMYMmvBd2Ki2B
26atd3+Sfub3K01Hu+UA69qS05LyvJPU6WZBkHQBWKvhwzndDq+J8Ajucfg+H3TwtrCwXZM1fQ4c
13xiT4nYuCgBMBFdyxn83S4LNcDt8uFCA1J8nsnu2dWdrpx5akqbScv00csAFS0yZaoPwu8ZTjQM
1eE9Okj7vfMDgSjmOZ6lSDPkFgLOyhJ5s9OlWQ1UWI166V1594/kCgp1UzOJ06FyhYjIJBAq20r8
dO75aMxB+/hicfkgKU0Yvh+Aozadv5m3TqYjfMIZzK0TsujCGkjDYdNsBezRXxiaMFxM/ZW8YYaU
s2Zqp5DsNyRz6ynWHnVz0GlPj2zZH9FZ928vz9fuths8TjSyBnuQ06JUdRWyBKI30o7xghBbQdcd
IvVK7UoFxM1/wWKdEgIY5V7n6xLKiSpSdDsZ9uYrn/+eED2MISZYMY8/C4RgnMgcvOnWENJGckaU
965PPUUX3G038m53Hvv43QraBZ03kGs4FXcsjEiDZ5pCkkUvsdYmOGOhmBL/WKU+sEJVgShM10jm
tcsV9TBCsH13VjxjXpnkaxw6i4ac/zrgusycXCGlCqWasT0yZIUG+h5ng58Ox1xq+Km5I7w9aPfA
ohGBIfvDHFiPxkC9gHHCnbXFAaRX45icB37UdorL6tsZt9YfbCI7tx+wrm/TMBWn1aBd/fInxNVp
DFnjs2do+BrpJHV7Fi7f4NBt/JQ3mJjqXJgY7XX+nmxgYGFdJQtztbVYhEN96FwhLUn5ZPi6KTzU
FyjmWCxcJUAi4+RBotIeAiGiWM6rIydRMRrOaxXFVCcYHIvH8GahNOuyKKUt2Rc82PrajAnGW3XL
lg6/4D+8shd/msh7mesN8QzsFmj2U+Yg9bjEk9DeF+B/FDxwAw58deKazNbAwGi7iyuVKDBBWWNS
AJqzy8o7WdrP5aFllvb25fFnfFJFX6w1z2kcbDmldFo4xb5+bHv598MnoFUIO6V/D64HdijC+2Ex
bi0y/QDUj4gdk3FX+LzaSLrLx94U09Gpq7zvtPRg6uHZkdqx08jUYX+PGmIPLe55Co0u/QMfkeEn
PvJt9JmbrXRa9gsmAxWPBG5Z4aDMJRV4ANVr9ktMfznyR2wFqpgbLWETvYkCCdIMRxk9kPkX/u4g
3QnDidTG+K3gFikn0+DsPrS9ouuXutOz47HlNN8PT5QYcrp/zs1FtioIs2rPPQMfIx9NMuO60/k+
Oq6eVf4N0vaSqDMRd103cpa66K/P48iWTc5ftG6PtsXY7nvPQDcQWYrD2NTSJLjj16YddDraM/bW
XU1YWrInbtymtLFAzkKvFg+oP7wZ6v22lS3Hzb0zjUbqqGmGA1mtaYXMgJPr5XK5BhXsYLS6FJ6q
KEvMoEpR8fvovwEb/AzSBy5qw7J39S+TdufPfmKveytzNDH5FWO5kuiJ+wgR7cL3+Tyd8t3hWtw5
PENELDXqMutOoh+fOQXnucPocl+0b2FYJWAhjZ6Hwe1nV3qdyN3Y6DlZqDaJXT+DJeZ1MnJp0dgV
a0UVICFhgvrI/iIGgXY82OPZUuF9loMCSIFsTOfeMh4Df5kFqYrEfe7JoV4fCXrhZt6GWPyiksM6
wNLtuzFUrt1oDME1rh+sU7Ilq3kmC2aE9NrdkGaFLnlMH5urFZMYqjVATxU2nEviM5tM/ARykWkO
XCeBcwIAKbSNoak7xD4v2rM3cf8GIRpzSe0Q0pZZsIfHqzm83W9DCa2IGcUkAsHDAzEJWf5124+g
HWYftMOAueL0HE2BNBj0Xn37hhkEVudhJvtCeQqxT/VLJbRsD/jp/vQ3LyiuAfU2EBvKsW8gYMso
gaLSfQQPXZW5q3t0OmlnI3J8YDrOZkDBV+Bv6fFV5eSM9ueSUHDw5sRHiliHTdrR2+a+FHP+aXS1
Ga+P2DqANIwAUMtMxcNJxB3TxZcRCep401yLIFDonY/qxTZLtaFRufR+ROUox43thcRqKIQzW/fc
aFHqnkZQzF6Vr2ItCF1iCH32r/nLrgFU3goWqei1M1cOPE2rAwlTUdD3Kem5+gMU2aLa+8hldhML
iW7w8FS1QrYI7Fj5vLR3cmZjvkCzSeSk1pftpKDS+iVX4DhElO3qGwUzP5qKRrMBeAt++DyKaeJO
mmFg9XEYLDgG3FAo10TVBpwQUs/LJkteOZ5GruGqgUJsb9meGsTxY243rIE58/JoeWWACSGDc7rp
W4eoIt9WLVNV/OjY3pxY5fqZH50x7zewb6lI5xYqNDnRlkCcQcT+87WLCKdkKbnyc1zQy1Vrm4q2
07FsEeWidSDuinbi6VmGM+KEUG6smnyaApTjl3oGkTUdFpfFyAg85caAta/eqXajINj5BB4RQG0g
1sQEZFgFrce74qlAWGyoMhl0ahHDpYBvwmkRKEf/SF7+m2ZV5dmmNZUBjDEgFzPxHSkiVXqV2SVa
gW4kxez0t6ccCfrQcxvLRrv58qRSLDldecUqqedlbGulix/iUv6L/05/9bPYE4zoZii2foVx+mh3
BGlYmhonhbzOQvbCzDH4xRvtEmBorNl2wRCq6NWmlaMSPRzQyiVsM4YZL2Ys+Smlm2/G6x2e0vIx
Kj5daKqKYBZTqu5GuObILBFrxafgOLMp/H2IZ4gnbt+ovDORmyfZhqDTlnWObcjOqfcyJ97KBkt3
18Bj3FLO0vkKb5anDw5uFxTa/3LG2faL2WSEXHRXqKGmqEflN8Djq4xAo/s/SQAps7xD1vL9JYMn
UbucEMl/XiSVQvPwZ6DSMx+H7etdgxBMzlNSJgO2jStiBvB751+AOztpchEVrlsss0UgdmnKuPFU
+ZRJyILNsjXvyV2m/hRxNyxzHj87f2hXzQ2J+y5Ah6jRSt4fUv8Rc88XjYdIzarsrGWKAirX82vX
ehzZM7lCol1MqUU22+7chmSwWErDE2yVuBeiAEya0NaRpuReAy01pbZoXaOKxB6UK58iGO47QaaX
jsX4y77+hHC1Mgf/tkS2SLEb8gigsCEZ9yDV4B/kpJLYSWTsvU5jUKG7ZgGeF82gQKgQ+OPJxPYD
FpR6su9Puv7ObN6iBppDL5A+YP/UyHDaCr1oJvHon9VpBNetZzHe/0rZxsjOrfWM0GdtP5zemwUg
+F3GOysgVXdjXvf4lcz8JzWSr6qKFYI5bk5iCtwhoUlPnUQVZpLJhtswseTNqIEfdrfG/nX+GqYi
zN+c0VcNkgRIv9hJ8ynwV+rpRJbD5NJzjjrdjqaCbZ5doJXFmQtRZpo3H6Fq5QvvuZBTVsXfTAue
MQDT1D0=
`protect end_protected
