`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 53104)
`protect data_block
j3UiMTf/XPtN5LkCBE93AhLn+7QX8egVNO1uCqd26rPYevw2oen50sJI0o/zrZVPmjfks64vrSfL
vyZfbso7EZagCbkULWoSu8/qRv6Vkvr817+4anIPvUsmnc2RsxAg94QUenaIpQFFi8Bqk41qh4zM
tjtCMiIkkaxsAHXnMEYnNGjZcXh3khTT/fTRDtQQx8JsuSINNrD66120Gg5XTXoFO7O4JAkKD6f/
CbJ1ZEb+QgHzwO7A7CHma3CuUMMQHjvzdUg6K4JBULRCgnTRofEN8qpFPwszRJB6kz2fayoVmRlg
s61lzr3Ox80iboJfAbi9eWvWQrNAlsJMFbqxixq45xaCQb860usTmgezV/Nf96YNxjmXZ300+Mok
nPhGGkMurBCH1zBZGfk/Lq3jG68lE68k67M+kILIuY2OwO6TVBRk6+MqEnLW2k1+zYhJZjFrfY4L
yXUuDXkg0RTLjj7emP18P33bBB5tWg8L6Ff2LRSRIf3tEecVDGLBgZLu4uqDwUIFGNP2qZZtqvax
m9MdtB79l8W+BgrAfg7ZRNygkzT33QKdAaIwuiToDMgbsw6MKs6czy4NPk8Arbb5hfGH1t/b3Uax
u88apT33E6dnKaYZBZB3rBGpdNU9KpT1uw7Mep+LYwwRx0iHpSfLfkmpfnVzCsgGmYjlYz2dMxE5
Kjg5vA4reogNWyVBOcLlwhONfCjvnfMal3UE21K7jWWK5nr4arcfIw05zVx5YYqFEOKdBA7USIYJ
uknO/LMZLtDA8Vx8JESOhMwifb9cdaw1E4IuK6srSd1HdydcTp4FfyVgAS/MS9zjPJhkrfuitOIn
c2Ifqss+aCCFF56am/iQC904YYg5NlzMYRO02FwCDiajW/pPzOPu9wxXpO/FssUB8kLgAanvxHQR
AdRiYM/73CpNKGtKj3pNGtr0io/bXV5vGfh1SMWB9PxKhDkkva+Pmn+b3sY6ZF4o055w17M00PiM
80h5vIpZi3K5z4Oq6X3LF2JaxQZsj+taC/YbKaPOkY5Z6Zl1fV1C9XAz5fHSP+P33ewW5veUiaOi
U6/suFIDSktOEC8kQ2uzPakurKmiye8N9R9kTPQx981+vdWcCBs2KAJqvB1qgCYsFFIc/rKKD1fi
jUO0Ch8frb56UtMxRHy8CfrFQkwbn1dunqMWWv/kWSXdTf0R4TUbdHloRoJrmunHToGS8Bu+wnZH
l2Wuo6O0RhuxJfSMEWtpQoslS+Feo8yqNNPk0iYubvS4e0l5fB2HjeAYPteZp2OpGS+1AlxhH92B
bgaC+YOi95PhHbVKrJGx7ldrM2SFQF2KM2XGJg0H99O9TDcQ0qD1ByK7BuiATxIelKOXBLVafF1s
Yaws/AN3BOSladO4YO1eGsrHKdfPptP3nZi6fb5RRuW2Q2UyMZ9RdPE7HZALbwWPWH73ypWh61kW
8+EjFD44XGEyLOyCZZa2HGJpc5eZoA7Hd+N4tdN6hKjusQGZv4YIkZu8dzCherOskFKZz2l1M5bb
oN7IRmBaJRd7QizCTZjTDdBu7W0LGhxJyKSSQHN+P+iJeCP+hQiSW/4kfXhzVfO14baMtV+7+2rn
UDlBcCKoxjopaqobGCqQyivHkvCToJpjqRAK7UYF8iUAsFiG5l4tXAsJ3C6BtHKF+uD2+ndpq9Z2
6u05r0tYpd7abwHkvp/sS9gbl+GN72Kq9foEniDE35EKwyjflmknueMPt5t50WeQ2Qn88VNjAEHX
YRSjgWIkI6eIA1adCpLbSfbBOd9IEoFxzCZ8gdMJezMJn+oaEatDK9pOHIthIhNy+3YJ5bz2u9H4
9sESVFkb4nUh3OILYdrrfSBhLs5awNd0O1d4I1rW6NDkkaH04GYablM2ICbaxzk9qBm8l9pdvZxE
W8u7PbfNWJFWuzLkpEPVruNl6SDn9E7mq2BV6QP16ONSumXQ0RGQRs2Oa+QSbIKIfWntbN+K1K4p
zkSTZh3h3qwPwFocr8tkjFjYiRMwg/02kaQdr9F8enX5Wa5Kqj27jpaiAsd1Eml60l4LtOmuwnlo
ff+4pTQnPYqddFP8xfTKrafQJlB0JsglRE5zFk5+GljVHOiW4X0syvHyujCRqOfSFPuGcBeEAOfi
XkwJjoj9xf7VcPMRx/fLAgsOke+8Xo67FbflEVlIrdA9QUVVjOjrBqlOf/LskpjRDcsD20Mfl8Jm
C5bXj26gf1d2OOOK51ztcnTHukFcRBjJ6e4xOPRBMvhBL2DeHzJ+QCPrxu38kP/ZV7PBMWh26kdk
y+jNwxzLUmnm/AB1aDHFcfo1uvbkics20aj14UOVFL87uhxL/1xO2VEql9/T5y4KQFYF3g3rpL7b
+WyH4YJ5HW1EK+VV6jms8cCapiFjXfB4aS9IFgAdz1lmgu+Vle+ZG+cP1cJI+suFsuNaPLo6gxpM
0dsyST5omBEW4BNAkABMMSk6r19BR1IrX/4NAqOXnFu1g3Cx7iSGwYcN5kM51b9XoIRzgXW6IY2B
+m2FhgHAN0YdWYC1Kv2EOnd0l/d7/FWGnxQ/aPvcGtQavurImfDmf5OHtKaBGlimK1Gr4uRhm3ch
YPEc7TRBqLbJD6NN6fs8CsKsviJVKC29lr0tjofbDqpNMP6nyKRLSAslDh3U3WWVsnCGjMI2EZTD
L7S1/L48L+xg13jSMkGYkDfFnKwCo2sFUQHv+aPTnjlObUpNbz1haJrbqD/cjSu4Lf+U2mF3DkHG
koJ7XcgoC3ybgzlU68Vby9VLMq5QJOo0aKylLSv0ij8J4B86qVMBOfzZGR54ZLue2lh0ynZfvHN2
EKZ33/unwzaABcU4Vhow8hYn0deNQLLjLtSLYKRJJVZHwhGOapxxYKRRDZFfS5gdC0pOnZhN/SBs
mczfPLksclCsHlFU3JYybVbClgKN5l2Rk4tX7dWa9mY8HaTROVrUlMsUxCuoTl8gVPg8nKRSbzGr
TM4QCViTdnXnaT8oJMCpwHHj9MYa+Oy7xNc6FzdUrtYjrRzyREHfRp75Q9JbIAAz5Vtx0ED3gejI
IqK3hm/AUZbAx/aIZChTNqLq/2nsOw2iUIJSGCE6tW5DQqkEglyXJPPc2J9k7zr7hEURU/xzO9zG
99eLZorEMs8f9TIGQXyCyHuEK6GIirCiy06DYW/w4PE06pHfa9EbzkKLUgARZJhgWdnjZnfVw/Ct
VI5jihOi6G6eFIFFGP+d57ic7J1ZpjTEFZ6PxF0JB5LMyIjaEAoak8B2QmIqOcoupWcqvMnA8Zwm
ajH9t9m3tEc7KkYd5swktHGcnd97klL0EiZGeIBtcNIQLzZMUKZmzCVgLdyknw+TlqwnrVAdKaZ5
6furNyZsWlq8uW4h+AL1p2lDyeKXS1aOQIr/yS8mjyQiyQ5WY0XwLzwbY1DccqvHHSmWbjM6tWri
VrYTbr1fq+JPMOUwyio4X8kCgzpEHj4K1ZO3w9Zek8gDJy5yZh2tHPlJoF9iVQ+LjvldQk9tepgQ
0zFKjA2D5M4wZMekVMpydjuxYo5aPYHUVZkh/FNmTmMQ6E2tSTXq1Pq3iVc3wd6MV1G3V8oQMQIS
e/hhYvbSzdB2onQNBZVGaUs/1kYG1LfbQu7T6vkNT2Y2ptiWppWdtZ1sKgT+/WXqcdtbSwSxrmh0
0AtlxYhounegkVtDDWQDxuH3cNkC2f6qVt0oT5UneXca70lzPXoKCu6Rq3E2v2KJPgP/C8DbbrAM
PWLZmnx4Zd/INQYXcRW60460jSw/INgebE7COeSwDngRPoMX24IDUBYvVzGkxwite9/qWM3TAfmn
18I7oxXa+KYGBQcGyVdytnDiCc+Lz4svBlGBLPgOR4zbTgRnSnnIuQ3ZibRhTV8MVoHe2kXRmiVm
mVuhOQtHbbwwzkNiainEVMiQwG91MgrPQEDhAnMqrsy8Z/1TStDryQn3lDQ2MyrO9jBz5pVX/IDV
dJ53SGqW/2q6WxROcAfnTGqzI/frufDnfCS4115RvChv4yAuOjfcsOZHilxs23FIP1HFu7Q/0BeL
TkD9Zx1kCPdp6KTa67aevT/6vnEcky259qY8i5XQPOutHsttNFFifnG9cHzXgB9sZSaxqa8fe62V
O5Dj9tJZs8Xge6LUvks4mxeZ3s9YkUWPUNSZ5JUsfSwGfyLugdqVLyc/HvfOe7dBXgJNXdlgNXSg
ckFdqGaV4uCJ8gToVmPoimTs1h9xBmUtoUb3uON1Yp+wL8c9wzeCh1LvEsvDdPIcTn462JR7OGh2
CRGlnzdI3tj+BzwqWfhSpiulvZ+jmRoWir5O2H25JFJWb0yshKBaszhl6cqADtar+hMcf3BIPC7z
Lw61lNacAQ1u0pAEAXdc+RA5jSe5A3ZmMv23M6tZnw4RtI0m23GqgWLgMtV0QeVrPIIQ0ki4zrjT
m9NGbeubWXjYmbTtJ0fDP17W334zKZWCUHsV1JCVO7SHzymE2r2Z8tixeFCbY6eteEi1F3+QONzq
Zf56AP7o/Sy9eyCIePVlZ5GeSuFDKmq/PB2h9QTXrLL8In+BiQj6pWnu/hl4cwPP3frVsF8U3U/p
oLwUgikIpUA7FDC4Tssx6HVIApHgQ7WOZsgoySYPFVHtxvwVEDVWXn7jj3lhdmwvuSnIwErkL8Qy
8RtixGt5IPi8gXbqlpE4gnR3Oshn2Ym+O1ZaomCmfL1VrPrEwrXq+2yw1hTgpzI1IA+ZzdoQskLc
RrXEAIwMdeQ7OX/HUEeUwaICACL5n9qmgfozrrZqlKnkXM9ntKAnH/IDbBwYYYvzCS/a6jnDEK09
o4B82gSuBAcx5vJztnnV277S8DXfqGuQYpm1j6W7XSH0MDVJlzjr72hTUSTQe8cwXuKnS1QgFwLL
aBjK+VoBYFomJ2TE6Pq3nF65p+SiEV+ge7k7fBNozk8XuZRQt7FW1R9m/OS/YYGQngKd4k5NdJ66
q0hYixF3fag2WmjLP8l9fakxvtGN2tGpZykltpGCbgDBsMSIJByWCVQTToz55atigqwXK7+7c9xk
egOHBdRgj1v4Vaw+Qnm1rWnuob9UiIkfYtmIattUe4DqjIHBVsOekrBjKmYVwydG1EgfDdQ8d+yd
xdmeGkCMAZdAutI6MQjCzd23mH84fooGD70RcrrXN/pOCK8S3ugMf/U0RBA0uQcUt5rhQk3WXvsf
OlBaIWcr565ln22A3ltOgL0oMAkQsfy/RlofrYDH9ZfC5IK8kncaQF0Y8kGuMHoRy8Xkh7LuaBfj
vXMAeYJz5QE5Qil+pl1EsZxukL2ZIGmsmX22X53kc3F00lC5UmCQ9kNqo3Fc1AA//fKn+NzemEW8
kKsu2FoNxLR0lldFPOi+aBrikrcqn3Kr5843heME/obB1O4oOKYvEtTEIksFU3mArYf2yZfCgCAA
8d3HHci0cRIGvxx3/hAb6FYYJLpUZZR/yB6cpn6//oCKD5yQ0Yt9tONoB7L7k3fpSO6JeFx0D59Z
Vf29Z8fYY7GwdH50NZ4u3rQc3cshtlJoDMIB+Nbq7+2fz9+2Uqw9KSllS7bYamrB8OTMq/Jnba6f
/aY8/EDbZivCasfKR5oMkCb8tQJ7SCYtm8mRsBdYXbQ42mjwKIf4jB9+KDz6A+2RSEo6ULnxEimh
TPV0sDSNX+n1m2kpDgY9wzEXYO3d+sMxUuXCwywYUe4XjigfrqNmqYmmtPUwW3tXByi9bqHJBcoW
iNSMqgScMLgo13KGoDsYwQhdzGw3uQxSqtL1HAMMBB3k86VXnZOvEtKNQnF5u+GjassaRAUcwEAt
8PJGQNGnhVqs/ZZgiv3Me8khc4toygZ7ytyFNZ6hij9gIQNBr3xRqbHGExMUZyKmGeI3lenj0UP1
OsFPklRgHvLbCjHrHZHkg4WfJ7X/H59Jp2NgkjOCemZVWIChtKK/Oqgqoa38bHZg4CQ8eGrsjbot
QfXxpYYunFr/Ns5uY1H+wxLqouf10MwPayanlTo423ELrHKYgq29TvvpCK4jkq8i19/ovDOaqts1
3uvulrY2HEmCIhHS7uUCoJffZ8VE/TnboGGKtpOewAh1APCyzzs+WdFhw+zMMojN/I3EgUWNxLX3
1iK1ih9x327tpp56Fn/mLw5lz4ohth4Y+fuJ3AUeZSjCOPEMq+ZNicqKap6Fs0Ugj5flnnGInas2
6L9cO2why/wWArC6oUw2KJMa8ztXK/Q2gaGTyxI4zgzn8qB9Tzci/RWipdIt5LD5UGNi3WMenyji
bNCZfmDbshmV05RfQWAmhCjxrUiOMfRsC7GN9j5otIJIWn05rxd+ZgVMr38zNbMuITe6/8KBEN1S
uVc0MW/OGsYJgQDLl3tZYaBMHpxYChDCVSJHH0882aR9xfjP8KtkHZbUxduU/C58vodf0u2s+PKJ
t820WZEwaqDTF6Nyq7XGrxHf1r3TSjvCcASEfWB3E25NCraaTzMZJm13J1/d35l+aZT6VezgUItk
01h7Jvab0+YdSLHKTo/FupReAkKKLrO24xQPRSHbg0fAVK/q9e0HC4oGEuAjDaDAY+u1ZdvWh7BU
EJhuAA7B9N0h7ro7FRvrikmFtaHrnOHnvxYpoJNVJq8kcCtUQHZXznQiKCquplnkly3MTl7PDomJ
8/z5LEWJ8GfJhBloQ8zPcFzAiYCRpY/4T4/3XxiZeJUTn+my189GkfcO1PyF72Q9oxD9c5/HVxQL
bVHpBeSjkWRtYobjeUst02RaigwJirbT4TeFs4wq0VmjgjYSg3l+GHs4s0PCQQSvEjqHOzwicAsi
W1No+nVobDtSeyYpO6IuAImiUneZUhqahYXUJFC1m9Gou/Gv25gUqqqIG9aOCRVhz6CFdK/wEmA4
2XTkQ6He7OOYgLyxQ9EXJDOZg1I9Q8XkgNmRCV9UR5E4Q4oehoTOIM8ihNinMB4DNOLhLcPPRfhN
l9mxnL4pWP13apBSTt5H5aVlSw2u2xBsTWa0rfhPIHWWVzmIm3gmOFgMWC7+ExHAodyLIEtmqiLC
cB9Xu3VXC198X1r3gv3Hd+fAVQWMl1TPq1kzEoowatK3ecsIQiDAU3HB1RSqdTOolMKpZu9Ysaap
rymErolI19tkk9tg/f3UCO/3ZyfTnxsl+mZQhEzI9gwzM/v+6Jk5U3lSrUxEo8ZuAuShgoypf0sR
rIXUlZJrl178CkbEuAL+iqVGD0QTCerfIFrrfcPZ3FwdzRbg0p2OwxCfPB9MjjPqfF5hTZxbnSZw
dQxkwiEjcN59WYYQZkLUuxfjJLAFzCzuSoPUJJtGqoMxlC+oSbMuuNIQzWBdIdO8oIAuQVT52Zys
tfCA+VUnntz6z5wKolRGDqUgKsRxbv1JiP6RQg1PXnIlIJcKD+ySdFf1No7RVoOWkNceArWT/zlK
6DL5f4jSwuYpOlx2GDINM/sCeW8Kx2hh7lMXtoRECVcfAIgLgzPyaDM0QJ74ALY6ShQxnDP/cTz1
+8zimO7JDLmY3lBCZ9u7uafyscFGw/2eTCBHjF5BrJnYgMNfoYXjGUGL8sNfGQWN8F6Hl2gw9RYR
3X/sHrzn3/lX8ss0pmiF1jO229f+XwOt34ZxEVfcM27drktG/w/ZG/cUWSch3DWkZagnBgja8/GA
Z1gJLhGmWm8ERMToNi2z+nKrcTtjru22AiChUze7ejzq4kMoYpyQKkrsAKLx2hmeUcBk4nhOoFUj
VAwZcrswHC3LaNsMLksZHfjxv8MZ5frFnCeR1Tg3LSUb7IKEKTDjVSe/YKWCRytL/gOdGfkyuess
fQ3V4pWw6ZbjrNZTWmLq75khgbrMNlESgS3q8wQzFo14shv53r32LMMfpaTYCTyD4TQO6XUwZjdz
F8c8ybjunh9CLiednT6yhaUB3E99n1t31wQbu5C6CixzRzvnd+vi6JKK7ZG72dhbmgzm6yVF60q0
s+ebG94Jx+q4WAjsPYft7XZhGfvETm59TphxK0MhrkgiZq+mXZ8UQXka+8JzOan3c3hY6nqSqf18
CcEKwnypd/S82GAbR0mQ/EcGGIhpMonNh9A62tUrl5jlUA95/PCCuPVTvutHViZmtme00UwLH03C
no0dH4saEaCDQf+jATUFYOHlP3IVXE/G6kaRXJRvkeVekM0wE4vrRnU/qgmI28f25ZZzf6Nj+5H/
lCnd560r/RzyKc/zU3iY8YSruxCQCwBVU3dQRD0GuIYd/4W++lqHXMh70lWm1nWhuER3NSD7ONVB
DJi7BmrXLYNVhK0T7eCVQqVXWTAmqBZldTHOqWSvt5jiYCYmg9VjzhFuDqTKb5eCDij7/cBoAK1X
QuexuZSnMrTJaN/0weQRPtzFq1r4ykUla6u03VcpKTcCLXFk7vwHUUU7izd1jlfPs/0ALN8drmRH
GXwDqcZM1fIUkh/H/ttEWnP1IE+QoSL3vIG2F/wDs+BneXe7/kFKaYLM4EW6hHRFzomKGnFdnnGU
ZpzZH2jmus2iNcyzDLuUQF7A2Sf9KpxC3+FHXD0P82sr+Z6hIPObJFqYDmraREMxTzVMuqAhc10l
1MsA7FwM5Xa+QxUKvmDHm+m7/iqMZhXHp1Qp5NECo5nCAWo/PnmFT29kDqi7doGtHYsBzv2p+QKF
uOU/8HJcczFCgcLXd0N2Kq+hi3SfqzeLDN3Om4PO+vj/itmIFhhgQH4vk0fKJG9XscerJiQ4X4j3
+9WJ4JGMrzrH/dB30TLG1J629VmUt0IRynagPUWPpt7HCWM8CL68/xLpkz6VOlTkrsTyXODyoYVG
7b5oAiZ5NAQrZ/J6kLqYVa/IaTkG+nyWTg3TLOmydOQ+cQYy9M8uBnBiu0SDZs6IEZxpBTYqmbcd
oaenQS1Z8qIhFkSA4KHOhBy1M4CUvLwDQ4hYdCTo0VlsUjPaLuClZqVSiCfCWlE8UIrkq21FyA6M
1q+ScdbRLOHfGtT/sbdQ60Q4XZzQna3VE2plIomi4XFp5h4jS3qq05+BI8t4CZMHRR223ojvTHuc
2HySJ3fEn/3R3PlRVhwlck2L+R36x53NnkVRTHTWVTDUXpuwQth5ri+5PoM4a3K3qKxwrMyOjNoP
q+q2uxraEF46ryKyixxKJG0J0QwFDVFZFTdY9g4hrzdbSJ5KIfptTaJGS1GpXAm/FMBk+hS/puNv
cZCMne5Jm+E2FEENqpU47SYbwqgiGy+6uQIf+joVMJrcsAPAl/sVrX+Tptif5xkESGw3LB9LgRuB
0r1Lg0c1f1MW4zOMPsQIWoVPQjQbL8oTFgCj3MQQMOIO5Nd2/EVa7TcnWwhNgc3IGUX9j6z9PQv6
3VbJyim2Qq3I136nnKei/8eFZqJbJlnanhlG74zfjIejjW1+vej1RQRDQRUzKFo5aCYnkQhAS21c
o+f/TTlosF3DWKGbwUxGWOlOqvqn8cMkDaH4mtF3Pvoja96Ntts3RYWs3pTSUY4CKLStw83+EOl3
mWOKg9GnRbKjJH+Gzjs4tMJjHvfulBUJDu6KC4iPPjGnCTzf1MMiFIkyVsWCFGOi50zymC1hU+26
BDpFhh8CGJvF2GWaFlUe2lpBNZY5F/2tWhZaloD+vh1X/GvrykBd2IdogXUlzRY/Pc8tw/+CLa8I
yHaHFNG/n0DEZmxP4YNB4cW6APl0ZH2Qng5x4uxA++aYG01CQBQH5zYKhAqTvVHo2Md9TF5p2w1T
XWdN4CkrXPaD72k/jcoEIEe6lE5/qJXechDDRPe0yA9+SccBYIuWlIAIxzGtb01nq6mt1vtnmSLs
fYwlTUWQbIrdpeWEVqKj8/lonxMKuOYIqygyMyz4flf840VqIA7FfnXFFf4+gfVV6VemZLgecvDr
Mii21xoKrUFsWJllpQtBFJMuBweVCTIvFJrjOnBfWOWeFjrFM6gT3WZ9uBXR+6QOlDIWf2tHLJ70
AkyJOZt3AnbdLhz4HjhXO5CsoHiRDJ1RdzfG6JA+Vw50WPG/w/YW1LHY/yOQvik828rtEpqBe9OI
lHY2AmrwuAyDfTsfhaRqcuIbaIC7B5Ciwf+DtIGRMp98ujGFGvQRT+1SigaYiB2aC+hFyd9XOscl
OxI8BNPDxaR6QVy9op+aAAaj+VU6SfiQDTpbfd17/WWHDN4vhKnmX+/NoO02TA5Xz3z33dQHvUUq
9eTX44ZKX1kdyhdSSpw+1GsdF8rhI65osDEM7XVoH8neKOfX853odmEGy+X8+oCkD8kbxBTM0SYG
gpAIV4PnVfcSbg1MlJbpyaFW6z2vs+6Mwp0Xlbpbt1z3MOiRDXoyK5EwGkI18Jn5x3ufBfaEWEHW
/YIe4uuEJ7wTxtXooe5EHkGNL5AOUm0eXT8tDC16wQI8IMh6we+hpc3yfnwAghENs9+xKT51Lmsv
UYsvzZ2O3SNp5WsQBQjY4bzDL7iKjp8O7nmSQVEi3pJ80+xv3VnjBtoxMwyh7tCoXuXOE1H0W3Ed
hQlbl8EuNq4FL7a4EEcy1qi5+43YoJvRF+NvKCOoWiq8dnviK52+qObNqjFDbdp4+BHwVrrINuYc
epCb502sDmRdT1+6RHc4uLZg5/z7JSYREVAPE5qhzt1RRnL5MDP+nqovTO2qOwAb93W8AVqMZ79N
savCI0/xat7mgsGpOxcI1xuBltbn3K/u6WhrI9yClbEjdsF/nuNc5/ppYNu9Uw+D5VjFq/cv+IOj
8FM33aZA0snGiY97fw3fgwRk01dJ+vVNBbuHFAOeOIZZXbGIVJq3HZ4IIYfBQqO3QsIkvHQ8f7Az
QlB81l78qaEYKWklg168k5RkxxxuVZcWQaH442nZ3FLsc0deKLrtq0HtnmC40OET5p4DgzwkGOhf
UyKlGdW0tMoVWLGQ1Kqq3Flm0WmmDfsD+u01l7oGcOI8J+XvNyVd2zq7cHNLcaiTeAB4imnpcHW9
1g1wMN1F5vqhEndfJiXzatZXOCoXocA88pF86v4icNXCKSqxgC3/3X4E0tmbWawzSDbUxSW3rxNT
o+ct1eEdV6yYNAIELeCGxdEg1gLYF8oCc5KnqvQ9Ai1jNAMeR0iWTwEyjj55/YszBtHi3LC9pPFb
ztk3fqNgM5JGNt2lTDm6L+n39WizeWfEIWMV1jPL32AwSQ9l5hzFjbHI21V/ohnHjCiHXRITrEyY
cwChvc0Q3cz+Iyyy9ocThFawjwaFVjR+xKl/Pw/U8GWlJ6M3kfoPeZoE0pytuz7XeolW/mMvvSfv
jEs2jDUuL+rvwgUwGen+53oJWqmOtEHHOXPfo1pmZ6o6pG1ty7V4+RXXN3p/72dRw99im5uOAa+i
io9iXfAezo0xgTjR06wW6Cfd8YKXXK2VrfV5tdaH6fITlunTF57avGhe8Z2H7TSPN8qdxQQSHcJ9
PiXo4h8jHqoOmezypvJVX5LjnA4R5ef1A5LGNlkpiqyVTg81OcH9cERyQShjp0wvbm/+BoILYNX7
R/NwaMOwLkSQzQCooD5GvHXX4fSRPusJO4ECyIXS4TyJ0fnv9LgNQegtTjfMIEPBWYia4iEPTlzG
Gt4iJDCPKYQcup9WBvau9l/45gM0IFfBXhjK7CqG4E2WwNtmVnPpWe113taRGBjO41xxKOLN0/0P
M/srD0ou840+EkUTHI/UKei3X9gte5/5oEfftbVkSB7i9/xvvzz1cfSJ5cwBA4/F9hZz1g8PltCp
XzW4KsXsCyoL1X+jpO8+HPdQhdyhj1tyGBLaTHVUL7bgfiGNq/spMPsVdEN8U6ktQ4F+qSkWJrGA
+6dENmYD4UvjMqjjG9tmnPqJWU0UKGnFI2G+rKAvCRjVgFMapTOdHB82yJVlQcsBz3oly5DvJkPK
hJTVEZQTKMrsW2LK7cq89QJmzx3NCGPxK2H0TplXrf7oGjs4o0xiwI47R1qvu5YO+1JqtGqCpMpJ
iHvAK2Qae3igXkqCWgAw+E2BmC9xzo0aPi4vow9u4AaPMZzfD8DACenfW9vOi3i/tmLdtA555Fr/
xkmCLhgyBOFBAZQahkeag157wv6FZclhmXn7t8UBjwUvQCJroVmDbambrz/VgrsyZxQsQWrHpXia
vasbo2C5J5E/sCaTjDkNFu0IRTGTrRhDabYcpwxyWilNmsZY//1sJnwJ1js53SHzOSN3V1gLbeMq
kta0xFmcYve80m3L6qy44bguKITwarDluSOoHeUYSORtNUS74kweFLTN++D9lYF+8tLktbCnETvp
F8G8QFOMnXpqVLAHv+yFZoURMotSEaPKD+VqPoa7zgCED6MMMd67u/Di32w6QJPD946RlBTuhBxr
R//gN9KQkLsrW+hvTOcTTIdxGfOk4pfQ2ze3L4nKQ/glJxlulg39S9NdDALeYdALdJWUDoovHchy
dy2FYsmBEEBwwDjKtXk2WanOcywFjbCbeQEBXT2REWtYCfgbSmRrkZoWnzNt7BLR5dMs9TfSpje1
ZHJ/paS7XWYBRqrj+GMlKffhTbzvKqYZrhQ8TtGNVtf15Ha2MpHryc/rYcaTcgMMm8+j7GzJF2Z/
YBdljTMPqpIGpon2N38j4l/wwCgMzkwmKtoyWS8pA5azMXvapcZSSxgcyCC6EwhvCjYCYs9gU0iE
XD+yhGqW384gbPIyk+X8oqOVhbEP7UosrUexDZkM3SzOLhg6YUmN/7soeKcd/IH24KBF7yBSap4u
WClcq7kibso1oiBcgMkCdRBMb/65wTuuQ6t9B7l3VM4OLkFjQSrdp8eAQzZWpmnKynJD3nOgXMBo
ECZB8OnCxTpRlGjndRhV2GfzbI4xIciCmxpEgJ9BdFTsjaDqw7XDaVV43xoffitlA0RIzrU1xBoq
94QfUSthAfGTmrMU0OITKxZZsXzR5+6JLOeu9jjoK/iExCELQIcF3aQt7xWnYqd12Vi/1ZLCCl0h
Plxbf37/MFixIGl1Kz7MPz3umNT+wOASDa20HoJffazEpGwjN9mAb2IF1VonZ3wFITeWwsRVZxl9
1oR0RWIx8xeJERerZbQomMaoxRAdPyg00VGPwhiAApaJbaG1PT+dfeqZwK2DISGGDxKxR08OhbDG
5dPhNBFh1kqY5FvMDZAPcw0xJ288grxjTJMY2wP4HuHxx2js29LBhh8RwMtT3GNe50qJ7b9SrKpW
TIJmHofH7x1euH7iI8144wZ38H0Y5xQ2ZEkRsJkzGGh8nV47uDEIf1oHhgRIaZkjJWDXq3c/eYlo
xMFZU5HeR8qBWY7Dh3kH4e1QjHOWhl3ZJM0PH3gW2b+tyTA7E84EgvBMf1it670YDPRi0Ygh7MLe
cuF6PvNeGUcVedBbwtI82mpLB/Xbw0Yx1EZ4pV0jipw93HqWBUVAAmoJ767hlpQbWFojSxtVZ3Ye
pgvFOKwU2Ca0P0G12DxX2dZrF+59IcZ3FCake/G4Croplmf0P/pyOzvatmCnn3DYL/Yp81e+dNXd
fmpgqjz2HOZ+xjNFMRE8ZhPIGzb82T7XlOLxgs+58ieaBUJ5T+OwUsvqOhb6dYdGp3tj8dI0aCSU
DJR97w4rRCRxwxnHzf9PGzwqD6l1DrshBB7TA2V383VOfUWBsbfwP2tZfqL4DuZThSQa7fRjkDL1
FEcIf6QTa7X4AzJbNSGrXI4ZfYVcH5GuQdIc7jUDIsxIwxHdJTH6l9YjOWXVMN3Qz0G+I6gI1IS1
VWQGErJ1bfl+GLhCRt3LhUttJMI+tRCV+oV6uYxhswZ29rPFiMcnDLnmoHtbFAKL7xioQeYgVI5E
V1ZvE1XekQkSTd3qpIfAKsPhIQPV5zXW5LSQgSbGmQpPtvVqu17zDD+20n/su/XU0Ybj8Yhl6GEr
p5RSeS+9MwHNT2pnjOk55KIVM+MPuq+8V2wVYLO/53laDAX2PF1yGqBmlifqKmt/v+32MSTaJ6mT
BoduKNjrgL5n3YzP4zDDs16c/vQCec9984iC7raYULmczQhpOtryE1dUILznhcLHHT7gJGmHLpWa
utPOxCjkndBL4yRgwAI0aR8gkWxmyqUMKGiW36kJnyEWjPCSxwF85vH6GSa0LnPizrm52iWgjk0A
BVc53EcVM/q/BNStTLchhQWN43OvDM0SY5EtzQVMxAHaO8QmLwOu2KC771bMCJdN4m1MryrPBduR
v5AhCHnxK0zACGcezvGGvgI1xp0sDM9p6tLKnVpP8my3pDJrMtnWRDwtxvdkbEjmrvbYed7ndaRb
hTM2PvgCtB5P07cmbLCXfbkoj2zYhxZWtztIOwbV+SitzwrVODuK7RSJ+VccLMz3zQed2aOntU/5
5DyrPT1BWQs6yM8xFz2Bk6ucin00LhOsYztz1y4Fz1ab0BltVTITWbYs1I14nhVwwQV++50z/2Vo
VFN1+txNXeGx+XN2rJtYE60Lqoyy6PTdW7QSoBhxTbIj7wRK9TWUXqMa7FFqqgbDk+NSFKEW/YRm
vDF6nh921G6LusUT1JxfMhTqY81w42Yn8xG2F0Pr11Jx3Nkb1jJy6bGINs9kQfep7TBwOKA4ps6E
Q8ZbH6JS1nl/N1zFM1OWrmsMUIErDj4PUQZH1x9RlUDqURFzBfnvlNLXbG6Lh+YteqsgNYi/0bxz
kSnkxzubaCVMUvj/CemlUwlGrTaVNOVA7MmfIv87F2vNu8xXTk1Xj4UKT8hWxZOhchZ3PtnPWeIA
LnKrQ+dAJcCEpDIJ9YW54stnKlHsOPNidoCjKTq+ntrzwhWP9iTpB4jA3H+Z+/epB0qrfX/+dexI
Vtrrw0KrcRD9SU35SMeBt+Q6liy9qG6NWcIyISPG9brypRSFrgP5H0QJYFPgMx7HVO/9XQ/wJP39
4XURgzJzK3nt9bf7qO7MDc0J0vvKJOlJbTIyklCHQ05AqZidRWxBIX91dNRI5w3sjtB7UkRwsv78
ugFZczfdLYWxPV7CknAyF6NJmi+82zEtSffz6UZAougUFS8h96LR8tqb2N6yp5m+zCKS4wBbId1n
O1wxIP/3ITrSeM4fWSlmmVbij5aZ6sU64oDW6IjtF93IrD2I6oAnciLIRU/L+j/xalZb9N/Trezy
RlDy6V9CwC2pqddup/1/Im68KbpJqs1joiVH4nWZQRKWjX0p5EyeWfZ0uCw3HaXnW5g0r62QwL44
3F62nq4PIRpIF4GjdbniNKVdG1qDMMrmX5YZgrNzewNRnzNG/B/d++P05LSy6u/bPgmoJ0kJPYUB
P3vTd9qxhWmPq7GKUc8HofGvugAqOgJpGuWWGR86Erk90N89l0fZp11ZcN+x2XQpuCWVQe7pzuNY
B0y+7Txcs9w7carLCVeve+HJwRDO1rBqqrObsD5r7hg2lqSEkXi61+LUrscVfY37Rq2e2y6qEfNu
Fb19b4H+TrjJuxQKAOVHyompYsfs4DEjCLKXDFwoYCQTPLJv0sfT0nXp7N9/yPohShjErtjeCssC
XFcpNb+YGZM1L0/6XUGreyiY8GuC3yd/huuDXhkd3h3aIlMhu13mGFK39rkaz87n8i9uPDQdX1AO
akfvvjEcQ8SMyqI80g2Pavt5KFrrVPjyGL9MZNdILDExXw3DHmrSmx8ivCVetyW/jJT4vb94HuJh
bVOrhnjqLmSpSWDnnX5DrYKW1Z7/Qz6BjkQCEoIwg5pSOIsWajD5LKM7pRZehv59+q6S/5qhkQFg
exMkEG2unUTU5/VcVJqGUA/v3Nt4KsSTHbu7NyMyNK1NrMRnC+Ijil29U1ki3f8pFULyEzbvjSUy
KrlZc89ufTt9WMGrIMyBh+qe9jG+/3vOiiBZVOYOCmFQbZ/vXxtutDRUzHPBCA45BkB5AoY7USQn
Ptit8iSkCGOCyCx6eFQhFG6mFfagsbaeUh5aAfsZ59fpQqkOPYhBTuwVAdkUoZtjnq8Spx/4w85b
dyzkMLDGN0U23JWXOe4EDW9WrRzbNNEBzXyZ586ufp2JYg0JurKEitwphFY+N1KjCQAhXO2gWRKL
Z1HLIQwrQirdZy6On78SwfiVquWCHlOE8ey8SAF1Ub1ibQJSYpNAaXPtj/Hhu7g6e1DFza55Rly9
IUs0qU1ieegfIMLImyULerylLkRaulz0DyF8geYuTSTF6Am1RpmNaThB8zvNzE5Hz2d68Dn+/cWl
EZ2pnWgw/zC9V+bVt/k+9dOjOB1ScvW4SlWcU6SwkMQ51yxZnlSkQ7dNcD07EwnkKzhw1Xv+g2XW
GntXGWOag7xdEwxgfskCzVH5vj619hGc0XLWT9jzN7WyTa4Dj9lbePkZ4Jr7szxHPdNrH6aZQyVR
bebWuXsHb3F08ax7PXonhoQpIJZB2s5Tu0OJ2lLHgljs0TFGWvsZDFelLJnG5oK1NVHDWsZK9Ts9
5g8HPYvKHBobc64twVXoe1sTeKQF5ih0zzoBM/g8PTAExiHROGYuGB+iWMb+TOINAP8kldy0jnA5
vCv9wXHHx/5M66xYjGvxfPb9Zpo0OPbAk4h27iDjEV7eDicXd7DmHAy1/toZrLwiliO8J06OdY0q
xmr83CR8LLBviA8zxr0TxmyYMTUg0GykglzNTC5DEyBqrISfup0TX8bag+BVTUmaR6JvNyxa1M2L
zi1ib2upOHthrPmO9hVLeVWlORuFN27vstmGlS//3rXdKO15GFrvgePj8MD8QEYKKOIuVK3WYXVU
K3qjypSO3Bb/pxKYWg9kBJq4kb4iFJUy8uFqYqxCNHP/KccnR8eUbh1Sl60iHOK1LRSW6300Brix
4LOu+ZnXM7x39IUwG/EOEPxx0vFJvEiBgQMErefSmSKx82H1QBr5ZnU3oQkPZzXt2cb8fITdd3Gd
2ZEZSuFXo0MA/FYoZSbXfHOzxsCSi2oDoYSeJXvHFf/ioT4Ce4G2oqe9vA/K+l6Ko+WWODj/h8ig
RoMfLWVhSiARD7UpPdDsCk6zV/71gikBnvQMoRlV35IkrV7YMCavVHxwzrXENm+6csJWSBy8WRL9
IgzRc+iXs3u/b/LE5I8aDgtmgzODIEZOsilzOJUv/EMRxtiVoDUR6267vJmVJXrIsKh85OxKH4rG
1A+RQljFL1z5HzTJkYTCEgZdSKllXCmvN6FNUn3ZGlv0Mqb8YXcFy3lkXUZqCzHIxv0YuxkNdKXr
HWHZecehHmny+regMN5wPbVcNwzORL0Agsh6E86a9ydVAonysbX2GevmpgSWKhCSCROoFYiMxvo2
Iwn3hk4BNeUUWb5G6zCGK9Q44MHz1oG/j5uhs0j+66OnrKz4+2gceVJvLT1+Hq1KIi848EM/vAef
cw81LgpKHcSCKvPHwc5aCdVLaOgjAVvN/ZrvLv4YxrsmCVERwxIF11lDDKAMGLflzxotWljZW2KH
dg2VQUz2p0K1HbdOpDLMpTrhPoItmBnnZs86LlTy9iDVFXBf0XWYE32G048b4XjFnnNcguj/jURC
7TvRmJotNHc4VsLJrWLdO5iCqvdFaBn5czjJKXPpiVo71/vtUe7hRPCcvo175HH8Ht1HLGxGZdUK
aPtnHhEDMxB2exB7Is38EP6J/4dyvcYgIdTCHNtsmcHCto8s9qYD+l+zw0NtU6US3Ghirsd1Kpwl
jo+qOci7olynJwlFGCIQ5Dw/elR+Z7fCNbROhKsF+BqI9a9X7YHaTjn4r7NmHnIzAp/EQUGx0kpF
BaPhvyyT85O8jaec64PVeRz2vHJvEzsoJ4XX7nGn5lJRDwmmOM9yueKshIqcjyX79aDosvOfH6ls
RqTdarJBR+6zGSzaYYsnN6n2Wv0BHbLoTyEBV65kXPjsuGEYLX+TpMjdNo7qwDyLRtYIczbLOQVB
djdGjIfz7g0euXGRhbmxw+0EhIaFcNVcEpiu0WRoMOkFZgQ4SVIUvaFZ4rgxUo69Q2vmqyHMzU30
3LT7noshqiXLPHChz/YClPo5gtBw7jbj9Qc803YO5zeNMSIhjoNoUsUSaal9Ut6r5GtIK1rJvs4E
nCxJQC+NJ1zwzcoqe3XcTzKe/EETJmdgdHlU7HeLNLzedAZBW6MKBXDszMeVPDLG1TrmpBts+Lrl
v9WWSF2QYA8WJAD6DttybZBb919kH5RkB+c/9kalZW2xtiGVQrT+mBOSrWRYEi1wbXfrP9Q3e9Us
MnxRyLG5aqv5prUcm1vhEXwVAN1pd0JDrmAOhnY2Xv4P9j9a2aqUOAIuAmFYE84j5YNEvCBgTWyT
M84ZgBCU8SeLEvgkQDIelUpYIA5ghNjB63TrvMmbLCugp6ronGZd8SiMXmseLWr70m1z3c0CcI22
VQQoJBGaYqUTyAA0drUPQEpjCAb40pJKcG82yuVVuQGmoF6QyzgMDapicVeEeyTX5YBOqz14QeOU
UcXVNAIpikYa0FNnt0AIGR74J20A4aOgOVtm9+25NeGg5io6XJLUG26pF4DqWL2qUhCUAbvO5VRc
V+TqNjFaDuEGyYv+tRe7KJFFoaLupBPxf5hWmvFBRlFahNxs4CaJSfnzj64WBH9Ifamejt7GzEgc
Bl/UNIHRTEaOy+JyZo2NQYFtZepC/e7blKWetZXJ2L3z17mXFzvL8wR+JM2KjY8uD+tmu9NujKoK
fwjSknGCtAU2Bqzwy+ALJGxUeE/xRcSWb0C/TGgDzhw8gy5kejZIps+Sh9lR612nv/k38phXQgeX
IK7VivTRSaEWNRv3vrez08R6suy1hz/PVFfZZ5ecaQt/6KtlTgKoGyfw9rvrcVa+n4tOVrMcP9bX
O6rC9fAELJ526nQE7meQyCDp+4Zu8nTbqb+R1fuTOUGZuqm8xfdxgb6vdznF7C6ni3zpN+chdrpJ
hU0aiNhHFBj8H95o8PO63Xvvu8EiFwDZm+0+hiBObPpA06ioeAnKLpcaHzxaola/6iuQyGRI5+PF
hMZlILCm42c0eGTXBTe6FmgrUNmMGQ/AY7xdtA1L/6cyw6ruXJD8o2Fqwb80xwJO9Oc0hnRS4NWQ
E5zaMC4dy7nL8vEpuH8xv9wub6waRxLOU8wrVR57LHE7Al85Pg1fzK5NyVMHboYxs6Fba8vhIvB/
R24Gs+/Bz2Lk56s7Va1oMw44WWQje4mfuW38NfUB/byKB4VlukSZS1AtHAyZIsFNvzFDFCBsN3rn
0d1ailgE3fzFYVWny/NFcXHe3MOEl2NgVD+3Jt1yLPl7N6YO1mXE/7aFeOnjB/waxSWzqhgAkFId
k+Jh6yJ3+Oxp0cb4HS9wJaT8pR3f0EwinVFC3/m976Q/XuSQQFx+BCJnIDRnTn45dfQL8Io6UVQa
s7rPk+Ki06m7CNQacWyK7VpLkP8tXy59GAZKFuVC0Kpkk2+G0PlQZJT+Tx2oWjZ/i6lkehnkNfSa
D3KHw8de4Oo98tHRwy57a4oQjERawkoie6+2OzT5c2JgpFFxmYMEzLa9Ki0zHKYy3sRrRJ0Xy2BV
lQR8cdgavvv98MKQ6fsZTaT6kHlM6zCNknMa4ck1IEIxzkAbBZ9eP/EPhUGq+n+30WzVfKrebFnc
FanMqedzckjmloVI16qRCH9m5a3Uvv3MpWH9TcYgaqJqVQQaL59J2JG4TdQe5L96/SAfj94wBj0o
OgwA7bNoi8KYVeqBzO3e3Gk85tgoMEnnRTvpxFWohU/fCF/GGVrAImdgls9SPq0r4lPP4S+NW7IE
RBjIKe7X2gGmddqiYPn/zFEnwiwq+JXkya0YIOnPiXaaxzi/SF0kFn4st2cik7GuUCeJnqkIuhQy
Guci1IcvY9XwtJf9fRFutWl6kMmP6om7qMtZSQSfd+sHlVI62S7NlyeG3KlVibd6gEiC2UZvJp0r
nfrHtgSDpH+zOL4oy+z2Qt7IuRw0lFbFSYy6W/SYKM8XfTmi3+BQBB6e2JjRtaMoBTfiNR2bxbba
BmPAu8++YirSEer5tewNQckr3mFniPJQzND/V4EdGz0Pj7b60SAobhVg8I52wiaXH1PwWCL9qZgy
uIM+DTOOh4dXwbNqQkTR83z3IqLedVMslldwpeo7a35jNv2TEJMTDr/71badgqsiBbfcJSZu8EUo
WoA9D3EKc3HMigQHUnwxMx8NuiNFWeQ+0wbxAT7wZ3NGx5sQy94U2GjoDhma3pLKBujaBISlLPxI
zKN5QbpsfTH2jmErts7yIHgs5Bx4ufxKNMrk3gXiZsdCQPpA5DtwS/8uj/P0I09lQPxPls3fV6XP
/MfJly6ERj6JBZqo6Vg3pvezs1FmFtgYo+9oc5NkVDLj3dGqdSqP6XUZ+HAJcHvYopLEZUPYzEOB
/03RSErUg0sdh8JLsai3VQ84mntr5ngsyNkXFXs/WZE/tHGWWzMXSi442PgtGlbUGMy9h0PSVb1b
+dNIanXhCPiF3hTI7A+F+lCAnhT9ha59rYIP2qgewzWChS6puVbKEN0xy1g9BElQwchFQC0yi0Tk
aCziT/qCfropEF5LCI1psYNsdexvoOXf2q+l+n4NNDNou9ZK+VoDnfiC9/TkahznQU4/j0S83X5o
tqTPXv9JE8afHUOC8uznk28y/YzStZxW67hiM5UfKj+4lzmjRaIVjUB7o0dXiJr042aLjt0uniau
4ANLb4LK6kwhXXZfrnUT4ZwN/hNTIXcfyZMPmnLzN5PLfhV90sASKJxGtsRyNB2Nay5qbcZp5sdq
AH0Ucj6OAjuI4IrSLRfaO3O1w1y1CWMpR4zigrJxFvKIgc3LZcZ857BIU54ngs8lwa3+t7zYM9Jl
CUhNFkiZWQnw9zmEy2Quf5xnVb0QRW7SKrCCft7TPZ8g/jJjZ5xtMbme4b5QestlHbsJfKdSjvBT
yFrKMco3miHpXaxBV5JB//t1iXYS1dF9J5GDnqpAw6QqADZGNBdu0pI4aKdjtV6Z3Tml7ANCYm62
0coblYomhleBRrsrMs+FiAJSznhKaNXZalRJLJnoHiGlPSkr8FMIV1DfgsrAkUixFv3pequMP9AU
X3/w7p58CnMcCICCvS0lpHmdfABjhgc91wzQ4NtvLRalJTrtsfejMQxBlZg83XOcH5EVtr05Uydi
PFdHQ6JxRLJxcTq/kC8y4nW3kMhhTgBpdcV5ZVdFtxtAejCGoXzktWSPZyENxt0/VOl1tHhFKRb+
m9WyNQjXZx9IpqMBTOjO9w8Lf1o1Tq153ph4vNREP/eS+yXdjMbH2EatdVzor/2/22ZMrGZOOoZm
lUMc3ifA8IENz8I2iRKQknWxPasr5reJERudVxF3rXOeY8GDmp6PkD4OOb8ecAU3tTPfdEzhi3gE
y9fGmAq5zCzKrMPFEAyDmE97ZDi/h5ErOAaEI0ELG76uR2WxPOqWdwPv5dkjtKUFjMFeV37O3sjc
Ufi8KXEtK6D1jOgLvExFb+JvFzAOKga3/NXECUw7FxDBAyMA+KGF3htGdRwnhBdqRfq/B6czlaIu
fuhMSDrxcln+tM1K7IwuNCpK3ZPiIEdwVhoApPagpXkJnU/3RS5VbyMDhn3vkPS92Z3q8iG6oftB
qYa4sZwhl9lbpO4mEvS4S6oad+QXSQlBtnXs38I/uThEDGDCszeki5uwkwDLRT4U5IaCRFdqdGx9
gNCw1MO2JrThf1KeGGQLhYYrx5QLfiewz5apsSbgBI901p7oSs/aEaAaUUDqGXvzMJ1tjwLVvSBx
F/Ol3UKBLNmIxT78ru12Z8BS1Kxivy4PnTZ9q9EAZpYgGlTgKQObPs9mk1qcdrLk4lIXRQ2vzbe3
PcWEhbIvgA7gOfE4yhVuS4MIuDcJuwMUxJCUYryfXPvydVCcgDha/zMr8Im1sSTF/UxS3wqSnApf
TUlawkm3xARkCbbopfW++0tyQO4ijr8mBlvFDqWew55LAbvDdtFghNX/ZzKoQnL3dP5CSGr36mkG
pDyW8F3MUqvh68FcTG0YyX4rKxuXNsgm6ahsziXrcXeezd8vSVJQfE8Iq7KgzffjG8D1BJhrruYK
dGjlnolsY7K0ZIZAFjkNhKQRbi9DrmwR+D2bq+uGS9GKkjpWDDHUlce6TsqIKQDKad43paENZszd
XSjNsN8sxCj839Dky6FJZOILOulmoTmC0F8bqLS9r4IwXJ/hBunsaWnfOv+idBYsk5aexH7h/Ejf
HHEadOqdRwxWANc4xtEJ8ncsw1x2OjjUpu6v4q0BuJrPI2OQYU5uIajtrti8QzUL/ckcdDecb4FE
kVBkekzFxufSI0l+MsMwzMLbfeg7xqb0QkQYMWu0o2R/REtREhFHk9y7fgIo5bgNazZDAM0Cin3c
cjbQKovkFKpJFGZjP+d8/2fveq3DvFqkyAnpRlIHPptWNp4LbJ08yPO3ORvgTyvGJcsCsQZMf1ev
aRIB3pZ3FBKhNerH8tABsNYOJUUvk9SgftUfJQAHBpwzRPHGH5PzZa+vD3O5SRB1w22v/UFEyPDW
iIl95JgczyqGD0J/yO+XsKT7VPyPj5VPdXp4nNUCKoabGJsxN8q5iVvi9Umnv+VbAaYBhbRXAy9y
WnYMnXJ3j+U9QFmU8uhRGg3sFYkb73HHYJpRA1gE11sW0+aMFODLkqwDD/f8xw+Gkyvb/zfzDjAo
SSMQaOy3YPlhET9ZgsR8n53T3WlcmFPjhwWuZFFoY64/ms/9BnxV/KsTUT5/h2BZNXQ84CECowBX
Yj9+JXLGbmnV+ur9UlnDtAbULei0lfAF7aOMy5UKmvcfn36ya6fXwtZuzPPaqNpUwUrrdPTArDGM
56J279ZvRMh8hKz2zhCdP4ojn4X3Pxbg6UGuQ5NSLWkOsebiOjJK8yeLMz+68V9tAuVI3i11k1QQ
D2CJ2w2NH8Ym0gQGdfiHLpOomylrU10KFYyFyB9ziXSVx8x58SmhR9f3jlNKAzLzGF46nJ9Xwb6b
wYcRt+xbRJdOX0erofbql+ARnOfYK5fYTqmomvIkSqEaeLl/9D9Mtkfauhk9mY1j630/EeumuZmV
YB3izGdFEXeyavCnyUMQyOcHnPmCsyY2cy+NB0NpC22F4nWSghN02me/dbHcMo0gPcF+jCo99Yrf
H/+NVPvGug3R7QxPjNHJkQ9sTw41I8wpAXKmrJ3bZ7UlBpQppEyXfVcE2qEBFX2A9uXEvFma9zjK
DHeWzHrbDX2775cScaPBGlq27M+suFHnPWFXRjz7dps/22kkRWlrRXOTJ4EZdJjrVQWjD5zZKozX
lqQezh2+X2v5X00zW5+X5SQXzKlfoZdJrwiN9u2bq+WJmadqOCU6oXwTMRDHc9ZkqUtZegx3Yahh
gaVuB6RnPLehztDzpi8fYJ70PwHrAU3+wO8gcZWqRzTPBbFaVwBVhGeRMHZy+rchiyz88nwR3fuP
Ge9LmKPa7jier8Vc5w/1gomb6eqUul+eHAQPxOYPbMGnMXKxl8VK2pyLPJyjGYkkFckWcYxjhe7L
jef29O2gIH0Koxw7WZXnGj2F9dR5yVoOLuNUVQ65wbGcyY2U2NbPkmuLBm0/vhfotpeVNfombCA3
DtHbCHAE7SS0+z7o7V3IcwqnUSrXqmobrtRN3Ct4miPTcL8Mvjm5fW7pfhA4Iy/YsWKTzDNTdnb7
f82MHDyNSol5k9gNneIMdAFsU6P5UMl8f5Q7ZWWSeEVzr26nOqrFBnRqb8B7nZ60//TjzcJedn6x
hHsfm1dkUjZQY4Qc+c+3+Ol/0IOvfFZ6k0KqUpB9qABpHOzDrcdw2wIFpf6mudDq/P1Noz5OLiz2
lkyQy+p86llU4CIjeSrDMv7Zy2ESHryTm4IRSE2iNWLE/aRwNo6V2ZHajDfysn3Ft9KuO5vyiGNc
lrC8gjwV+jnS1icTeKkqGlu+nnId+OdEQDFIzVHMyMlq/6o/Uqn8osf6O+0XUJzOP/JgzpJRHQYK
vTrwy3O87RDKWtgnSpfDS7xslN9+LEtfjNZTRel/1hxDqZdEIusnijRV6/2X4j8meLJ9zAx20FBl
//S1wGTpbCCVJAEhm89yCsBynAYZmLUmrdyLXa2zJw9Sb1ri5QGtybhjv8A2nJ+scAzpT4yn+Ph8
iJqRXJOCwKcmaG80QYB9fGIqhitKsauXpmglkzDIfQi2w0ZMxF+3WBGPv0uxLh35Q40JYC3c3Y1M
7FRJnxjv4vLrRGgNXd3MBJXFCd5vlArc0x0LM/lR1DyKlSOdReuqqHJvcpJHUrsytMxKgol9gd3k
6R0FJcMNEn2x0fRfq2Tqdd1WwahZSnmfJQxTiILqp2tL3FdeygnBia19wDRz2jDBEDi4Um51JKKI
ru62O2SXzDydqWtREIm0cvGaCmHbT517T+6ZgjWWu0Lz07+o5BLjFPTI4UtPR7yX90G6NgCxIDLZ
EjQBKhtQ2ucEHvtpQjsKlTyqmvauqKgzBW+OvraoL8PZG9p5rOa7MEzVrCvIiUyjpWKdeevsKPze
nIHfLWAAFNl6vk2h7PUnDK6CtQgUTkGLzcgxx8AiUfNNmj1bJpN7rx0FChEDNNrdeKLk/88TgC9s
oXgH5EInxsmcxZCZxSUHoU+NqCNhRodTqD/rSsy+VxvK5ifk9P2dxLdtMcwVmFzV76wT9bCx1Net
QBXD9/J2xkBgRvSbX2r7o3r6wNJ8w6spBx1qdM2xYtjdW6OU1MVp/EXthLxLDkYIDwpi/i68j0jp
cNq+7Rs9DpSkm8Rkk1uAIG+uQw09B2F/mdNRbnwieqJnY2gAJh3W0Ak1VrqIIZognhbu3q5Mnn9/
eVKOXVGx9GPOrDJk1f5tz2r8fPeIAVfGNBckABVhCU0vGSS8HLtqVcQn98OmfnuPnZk/M9slwgtJ
5c1GoMce6s4YqaQP7Bm839DUnc8M1lNDP7rBqdFo3GiKtb3w0eyTYcOl5oVatvu3L8uiWV0EfuXf
sjkeQoSGMV/tujj+H1rntZX66Inl99y1DPrvBSMHxeEGcbJHAvMlhYPiWcP/xryib8rPfg/YjuC7
4CNltlRQhu+qyJ4SD9Uy3rOsBzzk9eBS5o2OSkHEyk1DZGJ6fp2xMPGXBDkgPO8vAO9ifMozrtm2
d5l5sj6Lbk7Wf2smQIQoPXaDAVoXL/uKuW85qtKuK2ezvGbEl9gXK3crXCDYdY8+onhVNZcUQ3dh
gjaiXEKQDR91p6Ac2jX4NPy/Hs3jQmtpWrx09EdJ3FbBEN8F81sc9lSxzqNcOYYdtTRWZoo6HCJ4
kFRctVP9Z982QJBTijkeehnIJk/yJc560ecdfCqbh1zLsS4bzsUbGNFi6g9Gqr/apN4P7ycNOG+s
bj9AyFzRKx0lq4UDADHmJ3d28uqdakVyKD/UoRePyB1rcjipcvAdFEbj1Cio6UbXfqLb5KYJ40kl
jpo0WmuXuE3UpuahKfen2Mtrr3ApLsCdZGEFetI3AkfJrD1InATCe815m1A1JLG/WNiq00BU2Bi2
8Bb/PocLYIoo7x80h3+17dUZa0uw1Vi5ofaw4rx7IatFrs7GdmDBoCyB86iOKJdqIPMbtn5lBhP1
uhp1K8UFyPokJlnxadT/Kkap/ZaaZa7O6Ij0+96iU/Ce10SywYSqCyvdDF0SjEaFYjWd0T1Vq3Yd
JvLzwoe323QZ/p4ncSWZrxY6IjVnwTb1OAsKVkV3b8FJRuxzP8BUSPU/XvWNt4o2bzxEkuLeJsAL
uUXn/7kcMObOar89RssfBMcMr0p5ebuqtcw/uUs5X/Z+rTG9XhOpv1DNsncgogz/9oJbwg6U9Q0l
3/i9uhvUPYOyoCbCPVkCJhgm4DzS91rJF6xVLkNyzt5UANRnLzpDlJ7fVzUNPx2CMiXqsXxhxfQt
qLmQcE8xhcD/uN+KA9TNE6S4NOj/YGnAAqRlbZImS3RyZBlfMSX6NfJbwrYtGldxhNcrVmSSuCey
Ad6N55oe2kVuF+kbDXddNNRwOQUIp9igLyhibCX0BFDuEnAcMjetX8QNe3DvrUdMtjK7jLKYMiwe
B3h70RhJt8fNpnUM7doZVy/USnGVvQuNu2p1YJRTFVsPvQGqj+3A07N1CsW+4lekBhlZPU9vI0AW
T327BdKxuwgteMWNC2x4t4QWYbfPKZg9BpjkAp9ghfiK7eVtEIcIg/AT5jLlc3M8+0emN94w6lp9
t+HQJf5Ull7GkETSMI7t2PSvysIwIqETQSgQctP/6LFkADlkp10Kq0uq66wZ99O3QelfPoiJNvnI
sTPZleWYOOwBO++iRSiNwqx85mZrc3KN2G3K9pDDkS21bQHx1BBPMgOsXtrm/5gR4s+/yNBVeypx
KQwf6S2+S/65DdQeSUQ8yiMEQkn3HgwF+alzateqbJtf32St7Nk6yuHcdXWyVqFJhCMy897iqQLs
67UDj3qhalSI9kkt0JfdTulfN1AKVTp08ECpojR07vWByVa1H2+CP/25zZo4AHaJ6lrjOfMMJxlk
2z9zLI5hieYqcLbGsjyVWieQLmMRQHgbGbzDqfHlL44uY6d/U6JRKC++fyEcA2ZXuqwrUkiDcDPG
v9H0T6g8Scs/RAMPOlx/KT0IXQ4JIZqPM4oQgT3lDq7miDdbGmL5RJIh7HNEYw+S7dhSnbulBl5d
B4f4YAQfeKCnsV+rB0Iw0uyHJdMKjw6WSA+wydgz7jl7IwLdmB2GUHkPHWQMzW236IO2/B2OAnIU
dnNFsZWF1aC5yyulPP4w1JCkalLKaN8OywY0HXlzbyoEOSLZdXkbGq/XlXhFnEgKtJTfv4TC8VwL
XpME8TnjBjBfawXGJDZRXwdyR7nlCR2Ladd+LQKsvNm0qbKeHZcz+qbjbYDvx0AGEvLezBmxwRk7
jdgWcILNRz/cGtSTQxE9qyYb/248aSitgZfCds/K36GKkItoica5XvsaE4oCTTnnhNyovHQjKoI7
FWq/o9aCXdWGXod+OqUi6Pb8b9+jPBPTk31cwwyYNuqy1wEzVr+rRt8z8ByaXFxTNepARJ0EBNwY
pA1aF1ge5SrweZxBr0cBKcx52xvoRFaztFJ0/HoyGory+2zQJvAr1MGb/xusN33F031vAUhHKfW/
pTtCW7UbC4yXqO6lXqBdhxGefmUjcUU2VzvQdPF0Ie7mJFO7iNlxHtfJEBKIsn08YaNAx+7jVAYz
V1PEvYoo3cf5wBj2TcoUcA5u2vnOrk3NeKxPArNEVkVmFNkWLgSQxpL+XS9vxPTQICpGdHfu+cT9
IlOJqOY8cd6noxhAquesDIVK0+g+DbWrvxblPXB8XACOcOcp5yLdQduJpgnc+VMREUrcvf6IoQB/
Fgod7yAglPiRsRuzUQ+6HJzCOuXWHv/5FEPIu41lYamfvf4eDPieYdYRLDnuUn49+ta1Io833Sua
42tkhWuLXoh0OZpGLkU7SJUiNVGooHF6q0FtMLGVuCzxZWC0f72svMg7Enb/BXRBTMWgyJEBRKmZ
+uHnU5fUBTDYQnZvSKkl7KbKMmwCAxXgP4lNZlzG58gPDwefEWY2cbzrnmGhxZVf6SzXZcC/TPaV
ETe3Kn5lM4sjfI+64qS2aiwpMCsnNxrvRPYhkSZdPip3jiaW4Oi1JMp+EyLTm0ZvVrUPXmDafWem
P2AWPYVrufP3BhRIfGWWszN5Ey8ZquvUrEXQga8NMjc6Uo8mVQiW1HMAmQumYshTS27DIjI4Spuq
ALimZgqzAYnh138tbVgqtmwWMybNNDMX5Pa2k5JtNnccI/cOn2LlcI8q4S+bFN+NQc88ZjdI+6SU
ic3Dkrb0UE6bPFz06Tssrk7A+DXl68HzqH140ge/9xy65HGJ2zgODgvxl1mvwz1jyYL/NLc3TFsG
chA6b9LDHJDtRA+W0zIxcpbDUJOoz2bXWJXUIkrOTuRyM3BwUFLRx2vFUvqRWDaR34tYoq32UiNw
wkVaqpBs5tmu6gbAp3EmZaXTS4IVQ6rEbfwqJKa+WEXm9cP707crNrnAhI/8UQvmYNoG/LTU4VQC
S81B7KhoEIlND3M12wCc1Og451G/nmO+5RGYHxuHN8UwlmEitR3kQqL4B2RDMle/iTvsRJ0zIYq1
4HTPpYgjQhyglhPEIkoJY/2xKy1udg0E9ucPhbcl8X2vsWqGcs4HhSFSNkB+aQvZQW3/paJayVF6
yJQtl+xbGfm+qtfFEmrPO9HAYIY3gvWCYyhUvpgqeqXUVCPe5Ye2r7uGxZEdsXUSjiVWDDGKBh9b
ddwt7phvgaeSMeqLxmKjgbP0Y78+YYeiGK+XpNCX9GzA+USO+yvwIGco7MmGGvKY2xXwRNBpYkf1
RYxg+O6XdMApxAlaGn75O88Plea9VXf57xF95gauicudDKtI5Q7dsbHm34g6eZNIMGZK15EQhpeb
13yteT3CMVCFFNXE0D2Bi3yg72T3mHpNBecfe3xw4qx7ebjg0Be8zyfTuVyj4hq2VyWmx81XmSsE
bgMesrteoS7SSYpya2oXa/yssLUVaNv9Y0ooB59635rSaRshfih7eRILvjz4xeV5R7X9axHQdMXd
QnhL66LBeo611O0uD5lbVqdsp8MQN5pLsUNEyCQCkJ+ec7Tq+662XCL1iHMS81hasqSPoMT2agBM
BWwiPOEOHK6ucWL/fRN7lRqcms5XgAX9akVPmE/JqzKzCh+QRcpB2iE5wiVwR5SyKZH1Du1IMBlL
u2yEmCGrot5Y8phr4MgW4hTDE2ZjyP1rlVe+Fg2TfWADDMDOTWsRQy48VS5IBwpZ12ci7D0EbsmK
couGwd14zA6hWGAiPixiuBEDo6k2L22PnSY3+sydgyKfveYLFe/4RIVmnE14Yjfkyd45BQWQOgHr
5iOZj333/j1RcURgE/PAQONBRwlFCh5ngdqjOsPspSHnR+9J/Tj3sZsf4lFPUPBuHtAy6AZJ+1PN
K0tDlrY2fQnsXdz6REcWIt2h9+7LggG8g/9pSk794ALcRU3UQOnRR5dxeOV7NdNCiiGfjRk1vVuB
gyLCwU69NQ+Zkpt7r8lJgFlh7sD8376eq3CnghAFxYpQAKpCFacHhIO/GS8cVU/3Lt9deEVusztO
aJ5pDDqVWYSPX5cwqx+2uyMA7IvAHJBXEjNb+C6qDsSh12GUOCGaTpJa/ACZoMjJZ9xcQw9ig9Mh
/xA4FmUKGfor/fw8R5TdL5WM/AavEi6I6PDa87XAnsGGpPboenm4lKH4KTs/XOa9VbbKsUvIyIO2
trlzwXmyv95Fu0r1LBw+H95QiT+m7iyBhVEvLasrkaDF+DueEp36i4cnOqJQM33VCOMTB0RZoojB
AiH2jDdZIKcqtootKgwZDuNN5Yk1gQ/nyBjT2HScNJI3sI6ljIvp6GQ9s+XUA1N1XIur9bhLD39g
smal0hfbsNl6XcMrjBGMyjJ+E2uNuDw45fY7jnp018ZHHbd0ICH+xjR22D6PGqMN0Isu7syoKzbT
Lzz3jeKDPcl5/AgNI75iifIn73pwFKYFEl1EiM9iUVNFqCO44fY99uSO8x5RXjKvNIp+QCXO5trM
bKH1e3rsLuiLPoGCGqRn0pUlRCz48RER6CZ0/d8KSXcs9v4IUd8Z2KZlgeBa+PQvxxJGBuKOMK2T
aujFj80js6MUsadt+wh2J90Jbe3mzbD+0jk+dSJikTROoHYG1t2oTWnIcQafib1B4dMdl/rYubGr
JY5dk0GK36UkP5OyW2UmHKuxED5J8b7pjVUR7dXV4A60Rc1QjEMwk8c7CGf7sgr3y7bM4wwbG2vf
cqW9F6LuNEF8swzvS7ZEmZSO4zTju8tyAYcQ2/UszWIgjjC0KnWT0TrXpkfKGzVfQUpgjxc1IUrc
SG9f0B9T5w+nhVgtxprnNhz3HFY6ChlTmciyEh67yUBBrxQVhWPkW9jcEwt3loHunrgsQQgA3nhv
PedcRPqIRyP4MUq1Y5qCpqpRZz1CB+xxdNH6f8/xO1oFvpdtna/Tw+SvcxE6AGEBHEpqvSiiTSCe
wZRMiNihrfus5nYkPVbHiExElkTc29Xpky9uP7f21pxi5ZcsJU/8wjVhieX4oT8wfQNLqtbTyQWz
gTyxWZBJhGTPwi+Axrd5I2D3Of26BccckzMEXh8VIz2cYKtRlJnlEyuk6yBJcEd8nJLaf9Ds6F8u
rTaRQiAsmtiJ1DO8SyVp4CxKXOy0NdgEDkJI5wAqyiZUJiq4bZpjjqYMwkplchOeWlYuWfVMQRsY
hzshcK6trKUv+LfY9lPs9TVl1Mt62PlGPbIegGTGhBYmJvLPjDYWNgi1XyIdMhlpWIVklB/fEuVP
7F/Mp55rlV6UjTeP/r+LxpGF8/BNOGxKQBwBbm1h/gh/Qix4zoUXF9QqCmrv10IrpMA+bBMbApMQ
2DIub8lLRIARes9gVaAoeDF44SzTuRJU2fxRLdNATnvkBp9vnb2r/Yl62D/XC5yXocvAsIoH9n4q
kFDMkx8RCeIOHi4Z3aA434uW6Si7+09wq1Hj2GLCUVTwTItN7hSMMWbKo0IHw4uIwhYG6rZrtfPp
V0DFrNncHI5QkGZd5WxWR8n/XxP/Lj8vYDzaEsCSVFxSvBvBAkvx9mYDr1tQrsIKWp5Kg2JM6ZQN
OOD+N77VUsbfX11+rSi4z73js7ABHWk1YtuZpEbIEIzEqcKvNc+VK8I7b5b2y8fnuiWRTh1rsFAR
InOSg8wctZgyTnWfu0scfqw9a1PGxt7iXwqPZlUTJQRmu9cPLRtcu+zJy98jqkOZfcK1XTNHVmbe
wxHnssGWTrztKTAw6MYSthy+apR56DURdq5aMyDUPPtRm03ZQoL8Ytm56OBK3R1DYNZhrLawzCeP
hSDG0yROIkjIxhIBZtrksGuY9kx3mAhcnSuFKPMNE5WbXFhOP9j4OjclAwXe6jasp9GgLbpGjBRh
TpDR9yjyYQ96Q4BvgxbLS7jntOwJ94Wadqags40MdUJ42KnCXgEZRUUCPqTBfG0Wpc8VnZCSuLXI
7ipMxi72OO1HqG64f0fCzdK4TSB3RxyW6vzPKmulbPcSjA7SJbD+jg82GwU9A7ep71tFMWn2Gt2r
orvO4skG+8Sw1t2NtF07WnHMsZUg/QtJ4iEFFnlcqwCrJzrQk26kHi5ZwwQ1VdgtpN0xhs9az/AN
kXLUbK2g1MjWEmEWJGbLPnGQpapBgXmdbb6598OrbJsdAczqPk+b0dNjtz9VzYJZdOFLndCNT5DI
ylytYEFTaWJIzozBKXXNKKmKZbTPCZGZkKbIMTZ9gn3mG/DWLePtwRA7DGE/b4cmqn14Y0INmKTB
EKo1P4FmHfucwaZYyqFZAlUWlCDKG59ofyUjgbYT0LhgJwZtvAxjS3YUfi1UuryBGkdrleke2xjO
oZ1IgtkxutPMATyK0Bu1KFO5BxqJAUgbTr7ockP63LMpXgor/srauHLzDQLCE4aEDbFgeud/k/YJ
jWhzMPBVi/JFekr1adfFWe9srL2EY47qlbYQQ3/w3GFxJvV9S38/hBQUNTtp0+1gZn1nMIpRW7Jy
YmDlL+We6CqyrDEhq7VQdadUgVamTFbdsRkoYOfrfYkfa5NrWnYuDP/V6MPxLTmakl2cMotz6Bzu
039ipgPGo5s/a/YSdD/F+EV0HGuCQKZDYSfQFaI6DLFYoNvQcy3JMdtanhy1+ydg+rwRPmcFf9/r
oWJzfRqibpWnI7EjX69ZUJCDAyQpcTE3oW0nryzpiZW2Ic3eDGqUShkm8GhGsniSX6+Z7W/D8Iqb
/JT1Sp2uHZvMg6G+x0UfnEM4TH16/xtTB7cAadKYsw9RV8Xwqi2cc4D7CFHJwrLbO+kj+vCZ4mX/
WPDITScNNAgEW4Qr3g0iFb2zZm6GGKbjxoju17r1Ng9HCUVws23wujcTbxmTDJfuYAXMy3iEZi9H
UxX+XT4chZecLLOtotY7B8iD/awdG8p4RHqHvArlFkDvwb2igRTuvELw6D8XcwZU2FbIXZiTUSRJ
xABSRO8UFRm3SpyUh94Qo31OnFmcGaeR0RXzbaoaVZJoHml4NFSvRtwk1q90QiQOfDS5DcHfEF6i
CamsIYlzRe3HKTfQ0LR1Xy0G+8Wp9ERVXcLSQQaEAWtIK54u5BRdbZaluAGsZG9lhZsC3vLSZ0HJ
ttb0Nzmj94VNMe+SXniaA7jSnhmXrukJfcvgDsjif6UJZiiSwbgjtLfcONSm60zE8R4+cvz/wpNf
mPKF1UXL+igOeWVYXcPYaftDOTetCpcpusDw5uewoguUCc2/z16zIg7wcBTppVj1MNqjd4tdjs4n
7ezrHHCL8QNvQ+uZCBsg8uapYGnAMM3mdUFV3sM5cPk9+qDLsE/t8eJf9pzeCbG8wGr9pP3oBjSg
N5irIzdohC7F3scQgT+g9YOrjwzoY7RjPCbDqc35/KwR+QBd1IQ4Q8P9SrgMA46lynYOcTMSGFOT
WkOmgIUJwANPxAtgPXCK8NvPilWfV6WFYF8WMs40GV1Ui5fACp6oFd5hSJ8eXRj4RvZeqYqIO3pn
B4N8qE3vb4Prepy8YDBqf005QFrpQDV8PoGP7FJhfhNst7hjWOb9gfD5sYW1zbMm3B1K7Q0xQ1x5
FCMR0ddLDntnXc6hCpt4YWA9pwKJhYRn5E1w8IZ/p8aElaL3jxBKGZWsa4cLS/TqjDYiAzYRRbxI
S2DJ7JdOIdiVsYjUKzVGW6QXCyi6fpHZMhQBxL0ixzlVnrE2FX6XYkTiYLap45bYHEESWsUro5qV
iu+XGkvzteK9MVHZxX2BGaH21OHMObTx9bj8/G8ILk/DrBxmo5NN8PetnIyJo+tqt7GPd4Fw7Rc9
jl/zjLPKQe6yikKvo0J976qpNrJPH43622IsXpiz2c08zIQZJu4erLG7vOAYZ7qW8P0An0GDKi7r
AcaF+u8yD+FjvBInmoj0JpTz9mAoq8QgifQf7qPdE4KiyppMBbDrH9pHPxlqC/e1IfVlvJoQAsOd
jzqrZ00drbYIwDTKwChDoIhbXAOZ+r6+pQ25BT4LC13IfsHN5BiXZtxNBMzvUHYN3SGzKP29aGDd
ReJ9wSpiNbAWJAP2flWXyFT2Xk1+UzweQUkW9BtbOkOYRdM50Sm3kuCgtruyliTiktmwOLvdQQYN
CLNVOMSFnPqujmHeSYV2KbiuLQVmHid9z8fGvrwCH0F0tN2u9Uqyx96fo4qa85mJbO7yLmcsQsvM
eySmG99tZZyUI6edZdb1vuaCG83uED8Z92ks08ReQnY9CaeEOAw4B0i5Yp33C57kqqkm3IiNeQ5E
Bocd70Xx9F9K4Xnppq8hvwkJxF9OwMT6ufWcemKrscfNuMftZlNzLdS8MvhXLgmFvC1xfgKjxg6d
b7Vp25zruRsr4ld/q+msEkaSpQD7DtFu0PJpaE70WU2ekxJbHeWDd+zRSnBwXHCsfSdK7NordqB1
OWYpAsTdyDH0JxfZzvRsnk6dO/w1WLeXWa25bkRsqlBNoz+yCWrM2XKvO3NXNCXUF6k9w/1RQlKW
/ckXlFTGDMS3/LENS7QU7nWe2lhtGIBqErC+9T+sgQPed5Zri0fSAFY+YgqapmOnS4EImJiRs8dw
p6J/9nJepb4TegWKDszP5JHL2V7h5OQwGIlWyZRiN7MDmVUHMOTBRdErsLs1lOfgnzWlFRf57tHL
612N4gsBdjzKXvF65tF8iz/KdtMNBWO3lp84ziWdSaPlH0ArpdMgfO68VxXzEq1oFqyOxYyibnwq
tJPBzFCZ5NCCmfnAYJotQd98Qgx3HtjVKvi97espZtGWqXziHOOwqfO03nhsuXZFTZjIZzYRBJJy
+jsZFeY8zr/14ac8na2sjxvNusMxv3hMArjza70R8x5CxTFxoDUcajwsBqrN2F1OSadlmZD98bBP
PlgCuQtDBNyGOTc7JhzYUibpVA0Uswkd7MlBMcH2C7uE5tVKgeQhtYDK6k9SVf5zjC3C0gDfYkdG
g9yaRkXgegoG5q4j+Tsnt3+25jBDguSOHLD8r9ae7LejuZREV1jHNMBUXo+wa0+NXX8AVNhUwwWA
Au5Lq/HinfTGK7oHC6+NMKLwh5CODzFWd7wtDkJNKXvhSveA018LeB3iMO+fu2iqAW1Ir10GMXW4
Jy6coZQ9gqfV7WMJIqmYitE6ySZAlus8wlNDetKHvz3GQr3f/CcN6lGQbCSzloUApSrzFvNW8VYG
MnWowgSqCft1Gn4Lch7hQHi/2hiMUaFjRUWjQefZr1AGKk0ADREcSHkTlUbIPTJz+3x5PvziVUb3
bk+Gl1SCYq7oqKk+xRUw4yt845sYFMN32C2trb4aUpDH9whCFxivPzNg5x4pWfMbXDUWYGtpEUzL
p7DMKCjxLzwqlE8zxuvwFP8pBzGL0KOPWFJa5D6LVX6BeMWlKHPaJSy4WM93XjH2rNCaSaZLIPze
vR/fW5rmTJJ4ql9xbOwzjEOQseOVLxhrpwX86bc8jOnJtMoIZQroMKjEIKbbZtWcp1sN2cWoo3AD
FO+1b8vERv9XxhW2E0EJRI4+rSVAPMNM6LR0VUdOTZmEg7Z2ixh+YbfEDNh1a/7qceKhVI5i76TE
9IxMSw5xZj9S75QXbVnUrNu/6by4pjzq6lAVeh/XDvCnSsnJSXfu/XCf42XzHGhggWvR2nIbGCJE
LwCMRABzpJS//7fagk0UCOsyITSDIQ5my84l/Abg2ZHI0bcsKuG+yxt+GSSPNXLJFyxIXGGf6WlD
1qKjUgfBZDIDxAONmV9g/NlYp/O81YGaddECEdkBX1ns8QhnwZZBi7mnqI4uSU5xyu77J0xRSmYR
jAP3XZZgs9KX/iB3j5Jxt9ibZgH4CPYaIdz2Sg86bPREJ+Lrcek3m+cL4W8VjCc4pRlAWRO8hhfL
4HfxC/71ByiXrRg8igTYgdSW14rBYjLIz/hh0Icjpd3us/CwNX0KLK2QyXeO4oTFlXOCN5y9F4Wh
aVc0WGzGBvRf4n/t7TupXPrFbZlVRj3cTJ9b1Qhhpqdql6nyr+WxDqG3r9jASP3ik7AirbShhv2P
VlkEzLdi3rg0aLwDDFFsbOQF8+tJDeejMA0x0uJFJ/avraAF4hzg05Sz4+BLF/5tN/ZAUPsNIy5w
Snyheku0ZAhRupEfgTlZi27AUQrGqtNbvEquuMB0KaJ988kPz9N1I+1FadvIHuLseaD9AQQ2+9tw
GfSwiI+vm45x/D3ufMHgTtgnuZ8loT3odMFrlhQuKvI3nKuyyZ8SDzoCu+tvVu+QgdJspSB/Nisn
7BcIFQ1V/eZfDcEuhZYUQ7vmMZlEdVTr/0eqPaMG/RHMNRYA2BTgh0pWiNb81XN0ijReuLWDySd/
DOqFAG4AOgdZlt1BLS+a45sisl7/opgzk3N+BeZhHTLe2QZNIF0yvivl/QZGP4JJAWbgpVqsO+qR
9e/WzaVUsYjlv7xOP1k5M6gmXHNmLBQrkvQ5z5L4sDD5QDjHZmcxZbjcogGWBKOvc/kUAoi4OjmQ
5QFx9QAFTBxMVAoUCzc6esUfqj44lZPBJ5Q4DXodEZdwBIoFdyGMHWQOry3sx5Rx8IOe6YLj9Z2e
YxNyAP/pDq9Dp0TBCX2Ob7umXtbN746u9aaIX5e+zj5WzTiWb5L6sjXAsP1DKplQO9JoVtxy3Iih
9+XNsGkS8oLHINyXJj34B8zg04S/Nsw457Go20m6V/ky9YsYKQAgU8w7l8KzUpaN1tUfRA4/aoth
Di1i2iqq2jc8/c1WJ6DcqXGAunawTbBPBEdlihK706BXHKSWD7CGxA5NAyciLzr54608Z5i0dIy1
Zgfa6zegTc3KTkbqLbZF6I2xaGDR9FTu04eZXhCd3kbpiK6VXark6k0FypsgU2pq7UBGjpaDdjWR
iHEW+4p+w0FxD094O03M3vWA2rNvyhLp3Tuyc/5oxCADKKJL7DuUP7Yct12avF7O0R4cYwrD/1n4
MxVrdFZpuofA5EE0rIQNQKNDSzXSzxLMXjoEjGLYIgDJRc0F05NVDjkKn76tS2U1XlXxDkOX9EVc
foUdggnztUJ0aJTdxiuOAdnM80fkIBEc36yfTqLAVnqaqvvOUOYBkcEA+aeNC8CmTaDml5tN5sjQ
JYKbsVSHoMJY1B9DK0WW3n8+li52eEWU/jIaAcSavLujAE6/c5KOSAIchzAh6l1MGt0DgAWhIpWL
uzVMSab7Y2+Uim6d+RHG1Dl2oTdL64N+9Mzdxdc80w6diuHRYjvH4o6C0DxcWRw1qtjQrQxfZ3jw
kIgyjSKUNZpGZVlctqH80ARUOy1rOYr1Vmv2TX4TgzMrpoP4GzywBiL75ywUAqqs1ItzBS95k0zN
9plvhQGw2jcoJYASSYdtcR/m/DAMxLoOeTe7La8ZuhsuFVJ4rMzuglSF6DhCrmpjNM8a+zdHuwOx
7CW9/19uMwbZ/LEnOL9UAIG+QrRUL6cAoPwefChK2HmiZBMCL7VErVS3t+TXkRZis4TKMTDMsd55
oYWFIYSgO9C0KsLNJK7n0Nk50NctNAjCS8dKUnmRtRb/if8N+mVZ792L3wOhq7gsUG9vuP8RngyX
ijYZnnOSCYurYYYIFARghmo22QrOc7NgVbkVMhzQgJqpfLNVQRXOwybFZ7dqIg6xsb3Ke2Jx6qkr
tGJrpL5tCcd7i024wjFBGk+p47CmdfQ7ois1NPdcSXmBiH8kofln3SscdlYnZXHXvAqSCcnH6KZQ
qZ86O8gI3IgYHKyNrg860+ZsBHDhK/Lzzj2PuFXYdQqLXUvImeZ3h5HWGzgnNo/nyxUBaEQ+WuRP
rtFL7KP89F/jaoqX8Njlgfp8l0S+aT+Tgxr4iOGRp5rt2fQo8eaPWSNR7yzKqy38Se38HfSuAN/x
TMA+PnwnRp8vErMKbnTjwIB/4sgKGNdTluILptWwYyMXE7ZuMjE2NBHgtNmv9+hUbz4WZF7nJBsg
qgmc/2E2Hph92boDeEa5v+sIAbQ84Z1zjavM8uBnd8BBk900J/vY17AU0zSATARNIgHYlzqFRTzy
rnc2iImHzOH2180J0fM9nvAfO5Y6fucHn9DLkdnjS00JNiMKiTDM60vU4oewbVAnjukX5lehFQTN
v+QTOfzXJ32wWKkmc/52o60XsqhdNigliTQk17L1zFdKugItrowipfosVZS8NQMcuoXCtnsxjOcS
jvGZtKJ7Sdcvyfpk9GCSeXAa7G+P4EaGbIggCXBMYDZKP+6nQ0tOoJzkjaMs+YqOqzVaR65LHz1G
jblcwgsz2iCRzEb9L+CohfsO+NIIqAfM7IJjseVYe/ZSHDh/NQLLDp+ctKUaFqv5xRSqVtTWTTJk
AURavQkDh3X/IPRYjvT7I5y3ItqzpwFvZLkS+9Cqq72cDB8egwaVztzoWyXhjb/1dvjavv0Pia13
XprVWqHCB1WyB8b9pcIKpl+fln6yZ3YC+6Zf4bpSxsQCqr0jR29LQrpttbNX2dtIHbTvk88G37QL
mAclnnN14t+EBrqyPXitTy2KMFG0MDToMal2qnX5lF/5AZ+jUybGy4SguGFCtmJSp+XAdzQeXCcA
OZsIAvxIm8TgvIsGqTnu8UzmpRiGHXeZVwImvaDqaR0O30STe4TZv2bCYcd6Mw6cnP9P+pz+tSsv
V3ob6Jm9SdaSA/urMksGTVlT2Gk4x7bZdYU6C4vzTvYHWJKtjFYgZXTgYq6Bwb2GkEjs7PLNnhCZ
1frZIT8W3vA1QJw/hB7rpDS0gEZidNZdzdRmiiLXXlWRl5hiqGSBTgYuXoEzUz0q8hQlYUEmI48i
sYCxMEGUCHy7W37wgKeDj9shZWPWxvw3gJ7xMZCYvacGgZu1CfPAoUUVKtj9EX0He63vg9NOWFKr
aZT8OTJ7kfDOAMK7CZ0iiYgn8IFA2Zuc0zP/JylP8YYFq6qLiO1rOQnu1CsWlf0k7l0XYGpzpNjd
hVQGpTd3lAodHxLcjlWIc4kjMcBarjwqzW76cf6rgWYQxEN52vYqsOJAgloXQb/BRKC2mDPq33a7
KJYEABwBOdZvNhF0qU65kndy5kcYwy9VYg/WYFjhaKJka8/Vo+XGU1JET3OBj1TojlFJ+7JCJ3UU
SOI4mCByFtrV/bgpOD9MISmiaqDE6zW4f6PfgVBG988JFQJ+PZtGRULdDhd0TqtWVGNEyw9Kkn2I
jmSvGWu69LgMbU4AZlNfP0bfrg6DXnp76VFxaPVA+lPoG70O+Ff6nxQw+SLdlkYXQfbVE7GmXIS3
4YlcSQXca4rno0eLRhShoQRLzHAheKoUSEX1M8yTbfKfo9kToMWkxV/sqVkA9lLU44dQ5qPJWcxn
dyIryjqAKqy29XB0Nk3xtzWkLuhEgN+yHgTL7NQULqFRvV6vyyWMR1wz7JxpK/CetkTkPASAjiuV
Vk/Q4fJa8gC4ZJtbLeaAZx/nH8vCPjCezC2nGViaDlbzKcrJ2q16/WgOdAK/DbYXGo/vzh9Hoo5l
kdgVHA+/5HKZCnFSvAZyon1SFEIwb+zyxi3xL7PAx4bKvT0eD+o4sx7pbQegbzUCDcO+We+2CPgs
VlkbvUJSFFAYiTC0vTgiMsmGx1+VTMVdDBezRHLlvv1+H3UTsORDMTrHh23bC5EoYXoqCiEpD0U7
dgE1CwLUGea0loLyt2+j1s+u6WS3TMul0MdkwG+xnvVrRxpjFDo7IR6/GhBP2kjIOMlGI8XVTn2D
4Vqm3cjn+Nivyo1rCDNQqlQst4lo2wwdiOedsyeDrItdB1D46qmCEjDjKV/gnQIYbJpeyB+Qluaw
VqCOzBErHmRdCqnu67usw4p6+mepkWgIHih5zO6F0+yg8zV2sKUt4Gj3O6vDJjJ0ALwDkTBZCuE0
0AbDa0DxPsI2/fg9fjGr7upRRRLKnsyelJer+K+obm49aM/uwtBSZ86EFIwoZ4iTSF0SoNw2dElC
KTRmmUUy4/QGKuCGgBy4X4GHFRG29iK6znt/CcOYyF22x/XtAP8PHLDtVr8AV3ZDhs/M4oTfr+XE
vnIlwQhINOuVn/8hgeF70fSWTxY6UFUzCFSVq9qv9zUc/V27m6+CUT+ynuroteSa7+oG28oMYkoq
Kt7AscOux7w5dwUkK99fl+mxHBkOLNAsINFfy4kusrQQDKfXxfhC4vsFHqz1hANjlTSGL7YlxSN3
VZbzOKYiH/sZWToLCc/F3CpVSq60z1PGKgz1it4fwEP6iYj7PlYuRGqXOGxAEeqLVAUPB6wXSlvj
DcbtbnJLH2hbcB4QoQWDOwUEm98wdspPc3SKas/V12chm/lcum9lZGx7IvLJreSaTbo33HzXJG46
uGx3cxyRLxcS8DBYLETmisOpDiVC1aEPtaedAEBE4jlcI1aTXQPLkx2NYII2Fb+/+zgkYziEzS+L
Kr2ovTIAKNU+McKHgbdSYCSyq6hRpdaXvBOsWgymOiPU20f+/M7TvUG9sWxhxBNqAhfO7HhfZ3ag
F/y4a8xVjADSvwDZp7/Ud77NXFiNNgVamgNEqlwidgD3iggXQGolsQOu10EBbWr4nTaI2nAQEx7f
R/nRUaBa+XImgn8CNA8lve4kHs9jxVOXxl9g51hlz89au/HuTiW71k9o8t0COFm0/GvxFjATcWyB
dFyLHgCEsL4VTjRzO/DRikWgIggQcgPATbq+PbfJm25lNFEyLfqmQQRI+2qr6XYw7VURF41+4rFg
MLrm3gKvwR8Q2sh1+4i0NNvpjhQHNpEpUbNoNtUu7yAF37L7Kf9wIR/Aa8ZWFS+RQEEPuCbZAvE6
vdamSI3t+PXoCsKl4RmSJXA0u+NM20yKHdpPHfwl/rDbbpnpebJ5cwnor3dCsya8azVOhnOD9eG/
z00oIiSj+qzcIPCsqiGGI8RBW8ijOt1jbvz7R1/3fVA3M5IEb7MEpLATZ7K+w/a7EnnHcmygk65F
kFmr48VzkymMWeKIuKc/G6GDfCBMwKAGtz97h9owDh6oymKn3AVgXJjdbU35DkuRWecNkCB5iizr
MXOiCuXRVdfcuZYfNGu4zjS2sdr1QxeUW+1zmkYA+nNGeydGqNKHCT67zb+DnwvmWXGpkWaZCusf
8gm2Kq0DZ5YZqHddyOd8i1F4zFyAa+NvQsEJJSfyzA9trRVGYo13AOIVV1TIMplESJLUHjooKuL2
Knx3VAHEJrxkSRANxordxktIl15xeukehgctJZkjggcZUtzM5Tt1oz/gesxLsCPvOzS7yTGFRqIt
MWMzf/6t41pD+nLuTUS7jcyYjEr4BxussUIORtvjTdyqgFqBPe2NXUHKb+/EoHAckGj1NprObu67
xbFD8t//LemAYTz/GmiLLAVWeb+iR1t55lxomKjf108i5/Xo5zGlNTOJJK9fCQ4ARWpX4hFAv7KH
zoeDnlKDgpuHeIDpQTMCCOFGRxoiluROGkuQKH6ViJ3zWe0i/cxWXsnyotLg18nzdFC3qdFfU6a5
tYFfOE5STFTqcW5/3KPnKNK+1XCrzFQ3qKNvV9r6ibB1uWg6JubI8oiLUp5TfH/luBxlmRArCsKA
1MzrmlId8pbIP0cnF8n0sThVo+6rnVu+zuAFwto0aRYllPw+2+KGun6w2kTFAEotTNWmU+fUkdP1
Ng88KLXiNR6a13NH9ycb2aPhGsPQFnXIX3kfk2upFf5CeUC2rhwPgkOqREpSH0nier7qvtMJRZ09
dAjQ0z2rMqkXVcVDGGTW8/8oh6CKCojTZn7XrQEGABxZFHkoqwnRsIlEYnQL2xqHtlZg6J88Pa9a
wv/jJ52UQzG4o+wJyOVPj0jaHerBfs7GFYpArJzOteAU9GOlgYyCOw1bm1tOp5npFmpdwNpIfTRy
3/CMWP3ZTO0tQr/9n3bfcw9LDk2bgZwdm59ep5TOx/+XeXAJUvrEi8B7zITntmF0blMV87NSFhTe
+RyqlOKihsMD8M6iuPTRe16mlJL7BeACB4hvDXKfAH3xr5OZlIL8DSNHIbTOZhpH52wVKHxYSPjx
BHNd6RJWtMN0sgatWdDsxIxvoSUVc2GBIIVZHDykBIT09yol+HM97V96NY/tCMqSQwbNOvFexqSx
3q0AoTaQgbruu8qqyCKo/ZMiawmSyvmlONl7pp5Nhcx6VaH7iyWdLwyczZr/UTRURcLFGuBG2nsu
Rl5w53501t4ZbJwoZZnU7z8pECFigb3ZdgJBcHmoId7g+KIbZsfr+bWmeKeEEjMV7BYjZJxHdup6
h1s4xe5NuZR97XHrWXPCzlk1U0rPD/YCKxYYFukNqNyKCE3zzh9tgbpmsKGeVfxAgyKgiooTW6TT
fFV+QzjdC9vrajC2+qr1ffbhIlaxbuiKG0xywqV9K3FvqF5jESpQWyzbymnsNyD+rlirSB0UAMY8
mDsxMEzD8QZoxPcQjqP5a9EY6eE3rHOGwCRlIU3EaOGizrsj/oD8qyzQRRBw9K6iq+bgVK/x6kfW
rmQp9IaniQvFRVKnubEFn31qxHiJ2VQ0qtWjej6rYvU1ZV2qYvEDo/PVLBbN2y6cNTI6i8/eUMBs
PRD9puTuT0Mb4udw5almYcp856frpvVREgtG0qqGqJqM380CzU9x2f6yHgZGqRbpnLt5x7Zkh8Du
y0RM8SKt4+Q3Snyp//iGObMhOJN3Ifg2NZAVFmUwu3SM5HV4fKn/6hBSmeY6CfFTRvJcmYg1nVNo
UdtihCfcmi7MyVwDatqHs/6uDn3/CWMULaGMfChc6QR8yyiOQ+G1JOMkN7xgR0lLLmkhDYJCqRPq
k+uDOrFxmzKOdF/ptz7Jwv2WU5Z3O3hidne6qpOpa9/9BPjTmYKWMgXq3BNcaR3pdOqp+TD8hXke
8j35PUzgT2Y/7nleVHChDhbNocSrcRZwso0yl93S3HUt2chxldbHRZYZlajnyIMjVzQ1SZ4lutwt
trSwUEMgNu3BVqV43iksvT3kbVGqs7peTXm3eQCR5MK6jibiakIY8HZ+i+Q9qpvyDWNQdHszQorv
7meqwwqcqRYUmAX9V4DtELmujHP/IWNAiU9dmm3Tl6a2wBQ3mrlzpSSvRbW7RSXcrtjKQo2CybG/
IowpED0ksEan0+qhvXwJOaE2nDto/IX3jE8SgM9/K7IyAyaudCstA80KPMdyNgsQZupmfKb2BIeA
vfGQ0XZhUi8AoXOis+ufRbtZZBgqMpRiL5upN8d2voRX3/U/Y9k0mAmQmjmv5rGIOOAqNjMmNNdx
QkVIyLjtevF/pTfLhQIPsARpkcuam1tpot0PPxBLhNfEiMBXGcKM0AcbNWVtS4sC3/6Rh7LPWQoF
TqPEMNdr+h3u2Nck3S60EK79sRyCFlsJ3lZ6avIX9q4ZcOSR8o4VoiC75uNQ3ws7hNb1wt0eP1on
eGEMk98jMVHPm6PiMQVI6AEah6qK6c3qmW0A5wBxKT9LEPs2e6QMvo+i1hUlgmcXfLPC/0gZbZDR
ZD16uY7cir1q2f5QrF1NhfCPmUxrlyMqe3VDHnpAMw3QpXysOpUQYqwJvomukOu8VpPj/7fie/H1
EoCq7QuEW6tUM+2K6sIDAJMyyNbtAnJoS2ylOSiQ5GJfvZvYU97nnOdJjiQa5CZphCL7FAR8xQiJ
7LOOxqPz+sGj+dYx8cJYt1kojowiaq5r7ZiPOG7EXb9EKiDgCPsMUOBjvNIXcR2dFVWTl+/m/lkq
mOzqFnla2lKBLZdPnKp7oNl1x7LDheE7tcG747RfMHcyHxKLABvkpNTgjkk1rL+51CdyNKU/Q9Hl
yAocTR5T/wL3dfD1GW2pDBnGKlHUhVONIzb/PArIP+JHKRMi0PdfwucrgseNeGrpHEyOgm7EcNiX
A1EO92pnxYoLFWungSDQhAT3G8oTqYv6dEEWSTcVoY0OQ6TKfQdXMXD0JdPoQDU9C85SoyyKba7I
FA8S2UtbYZkOblH/rOFIwKgLHGkgA2s6ri6cQpcltCi71YOQ0oeA4XliJPOszW4Zbs0wmFERgdXB
IXKmCCF+Iiy2B8a7i77o7Mm1X3f/pJFmYUKqLE1TmVYBjT/vtTJhalIEKkAELZf1obpYBEOVfK52
O16PGt6zBT9g4YTBsi/9AX/DTBgGcHMkdZ4iIzFDps3djF34CM++CqsJFKIwM5bG8AN1Fedn9I0G
1iGQBkbT0jOvTFpd4AZc55X16HeICSwCKWi7dQ5aCftJHI3plbpAxbI6GbeZ9BHNmfi05gIreMgp
S2A6qMCUg+uV6CKS/9FfWEj8Z7K5jjuXSd8WyIUiheIKS8dg1qeQo4kkn+l8lu468pF6FS9XHGuB
cbFcZGYOhUlDY+31snjqme7WntYcH46IUhL6XrndoBaQe4ZVB1anwaX7Vb+gFK6NQDyb3l6ojp8x
pNwxxYHMtZ8IRgonBxTENj5Nsyi54pAg+DYpSN/qM1AN6fPwpIrzfsaXBVc3QjUD+T97StJA0Jd7
e0rLNEbSgm74o8833/jteNP1Gh5AHQQ/1UWJfxmRWxQgi/IKagM51YDL8rGTBOS9g99CVyWAhVzZ
bIrf4HzBzVblnN8JvqmsVX1eNTqFYoKTKGAFBmNdYGpGPYd6NWUWvjG8lfJgW/D32SP5McYwYi40
AhJ7bGkWh0wP7BXtNOk9dNUPdg7l0IunH7I0IS+M3pxQosZSJHX7tQ4yV2UAV2jF54jm1YifzU7J
TRCticVYig4HtDYKVjVIY+G5IhK3FqV3AcZ4rNmAPUTZsMLY75dK+uvmKzCKaXicjB9jEgCIvj8k
GHuU7wXmtYw2cB0tNY8JuodcGsmHCvte8Ek9kH7k4+n3CABABXTboqhHZKfuPeNGT4CkTvtT43GI
CzjhX8/oS7HmOPKuXGPevsibzd8HZnRIHH2UmMrniFt+N4P8LMrS/jrZphRkjtNXoJVs/tUktihz
4PmMQWNBNaRMXDdgPtuiKR0h0AwQv68xpLLHe1XQivZJ5Dkw92owh1oH/qrAFslVa32twqVLxzov
c8mgGyAKulsF9VsgqT55M4mlyJRzFz4IN1VszixDUKxR/YVZ9Vk+Sqh23WhCqVJRU6Bnm59kxS7n
+xwX2YHSis6cFE0/eC/w4iG4YeVDtxYdoA6O/WHKcxhWzO7aU/9NnaQJMrpIXZYSa56KuCH3vlB4
ygx0MjPnKv5YdXs1y1Xq/CK5qXAK//h09iIrdLc0YLx9gfqIXqPNqavTXDMzl16KpKFMvYWblE08
6N7gATtBMVkC9EVVhi6BMEgQIOEBZ+0qQidY+F1WOaDP69YCCPFxPoULIJSKZSgABEyp6DQMl/FB
2WgezPRBRm6ODuPZojUbLKLYuLcZT5uzbI/Ezq+8o0kOsElsnFeWTKUV5QuLPJhVvKG8qGZW7s30
z9CeJC0On14fIEEN4cDzSTbuS7BzI3POomBuXR9gZonI1H/X/ub1UC/U3s372O1vzsqNXt3PAvmd
Vne0E4Ytbqwnast32xsyuO0SXxaSSuXPJ5FrI7IPmgTaBcNyDD4ftcr4agwYG89FsNgS2kyCIRkQ
iDmjNGPJqMJfd56Jj/gKUen+SLle/r6jomccR4XfnBhJA6uwWVWkeVHXoD9tzi+c5PTqQxQDr0LB
89mMU0SkzKoep8BOcqOt+6B54QwaabZG54LLVJF+x7Qoo3goEKamkidlJHTzszIJdkUwdrHfKKvv
scmNFdcDLQz5eircbxP5KYwNGht7GfEmIg43QVUO0RuBI/OTTn4k4qt6YJySI6UXoBzttXEWOu6V
Pefyhi4haRfRqSZjzkU+v3jKfVI/TwkaO5znqDPK7d936ACZYceVChYZmywsA/eGfXzJ7R+PCHAV
umSpenuzQk7lwfVwxU2FzUCWeRs1lgbV7AdtyQ2XCQ7ov9voOy/KZF5ojTJ6/873MXHFqrtEFVUc
YkPnlwPSa1fdpxWveUBwI07SXTgflID0ISuOoqB3dBvZCSp8oaF7qFwmJoHMj8mvfeCS0gCGyU9W
+Dbm4bAoxw+A8nh0/bglJAU04+ZPlpkkbOkePw8G/Hd+3bMOMAHiLmrhHPKVu7L7AJ5qzItq2Aow
m6G8aclBwvU7VZTb1tEsBoLUUXpFLFjpmidXCt17JXkazrn3eRvY0gBexP1NcfllgNmlYW5SSd6S
dPWQromtzphQwnJIhuphhZh9GVvjfAIwjZFzjbM3Q9YILjaXxPTu4QVZSsdxI3rrnLNfIFO4eaL9
/4WjQioYJql4dXFYiuLukEXWI0EfW0tmVkd6qGmdJGq/tINCHEvZ3b9DGmPnhykZb9rYJbsCs+2S
MCiILupdZU1ACM4NNJInPDC72k126IQHx9gRxjyQ25i9IG14/xBrk0czXDLUBVD/jw576v06HaMH
ek1q+P06oPjBFh8ka9HiUtaMFQp797G5pYOlaEp1PBCS+1YBNmVxtp11JpclL+3FwLP+b25PmjMK
SFtxWj3q8rBbnLuC4guOdRZGa3++kXcVzHpcwzs9HDi2AjEPK3qTcif7TgIqQe9siBnMwXsnBWL8
j4DInCPOSQngmsEq3ZXRXqDIYGcShBLpTRRhF1/mb0ywX7z3bEspcU0/Vo98YQLaY6UAGQ7lH7QK
eQoWBTqYHs2wb9iAnIUsmLUPjZcEhtDlYm0ua0F0H4/WpHRU2a0jWHz7ZejnR6kmHBX7uyoSTeqE
MCCPhpayCxsF6YzKEtyQI0ZIgw4Ef4JU2RG51t+GJ7v8jsQDyk01VhhBiZRjPXltwZO8pM6R1tSX
4QoGajFut1UObKx5JD5RFGua858ura1eG5ClgLLDG41+N1EP2YURaulMGWP+Kk/hGhLhtpSmS0jC
VG/Le4trLX5Zq4GtZOYxeycUmpgovbQeTca/V7/1vPA0Qw4l/AMWgWvL8Ph1/2Qo1UdozUK8v6ej
b18s/w3HS+1X68bbIkR0C19dThImt89Rhkb6XzvU62kZLOAYiwtg4lQrbC7/JTAos8FBG4GrHlr+
RhZdzZ7dPzwVuuYn597pvb54dvvCturuzjKcUME5n6R4llexK+ua1yauHcAtoULzhuX8H4qXnILt
VYdZBCViDV7M8XgFdik6OVsc+FSceP2Cfo/4rZshkXQT8kkfFBGvE50UQfHlx1mO4em46inn50Yu
Fu/oL2RcSs6qRAzejO6svHT4giasKoJkI1PDTdzyuQeVORGcXGoEkNwM2J5ZitTDM7Fayk69qoEY
0qtQqXiAf9I+dzxIpRbRVgUd7aZQAhmPfXJJxCsyIBJ81thJ9/7KJdE899V5wmlQ8Caz1ed69aVV
aE7Ve+UKposIQBp/aHZ/O2ywtM8HP7oMmr7+rUjtjfLgEDz1soL7F/ebSlqhhLj94yAsYi+iJtoD
eTlL6aOuOElSkO7B3M5HuOvabC+qAx8vbJGuD5J47io5eJ9/Wi/MHoa0GuECtWso6jGQkYg8IAil
GVt1M6DyKWF4dft7tVkFRss797fSzUOnag7WVmr0YUlCsNQg35KUvikVgEpF8BrmjugxVnUOJSUT
2xJYuwmZ2soKThWzvDN1iXTukDe43myVH98+K1S3gBZ+7ErQ9gTmXKG9nNrF+PVrHioOQhRoglL+
X6TthlkVsxOaOGxqvtvtZ2KDDkZsXucw9gu3F/BrXGIBiRPG+t5B3jW9Az4CJ73w43ZwAJpIDJO/
iUsTysZbedy5yE6m4JUOu2rbzgUbJE43t7cbaZhXadWUym2M0lo4mBRjwwbgB+au608I+s5uJ3MR
gCfK6WF9z2LYGhx4TGrPw5/w5uKOntcFPpp234bq1g/9kJXk9qLt3q22EGJ0OqJIDrcjTpCwxiAb
KNLipAfQqlhoUiaMMEcZSfAeoHkymUk9bsKsqhMWQ2skwSHzsLel4BMMhwm+nRBSRsIx20BBS34m
H8kne0j02iKkiX95DartUUXhj+vqqj0pHXzLr/GN4E/ne4ra6DcnI1pz9hUhkVPjMBme+l/K6znn
U55fOHIN+vM6dzYsF6B9djMcPdu9TQj3q1m9n27nyPndpns/rjILSKreoEtpnlTSunQABbJtcM02
OQajXOYYXt4MKlxFAKsMI0HkwCVkDdv8Jy728Oqew+xMpxeHBUd3v9hqngi3sT4McXds+1jdH/63
iDKwkBEoE2IGlJIBhGCQQvvwb37NqsdATDHMdvbfoeZw6TEFs4C08Lx82jf94Hi6d8Tm7i95aHgd
dvA0kOn0iKP10fsEhQl+bIIgcdpzffEqsAM3OZmUrHsHIywnw9FaEEFLQQa8CEXa5dkzrLl4jEcg
BZTo6kKtSzbh86nb58+vcaiv33qbNIDPNAGdVApsk6BRoHDD+1ccnqWSy4kEiydFzUVCzo03UZgF
91b+VdkHdBM2hbEV2duYcjoU9nhJ2Ae65IAr3Hm3UGdpvlvrYjVCEhi357CEPWRCn3wNBH6BgVo6
89RBlRO1C8QH1wmsF2uM7zud2nL6ZLP02Tq2pFDALxIgSXJehYplPk72S7+uhWD7lyavDa9il6LU
GBqEN9UR9U1zjeCsVT86k8LBlKK3pmtdzQ1+OzZQ1LH5+VHbDORELFJDMQaSC+9vkeNp0eV6vLz8
HgyGws1pnVF9x4VTL/U3/PMG7/km3poF4d9uD4h4ZuUSrQ5iuUr1jVfDMEV5CF+lM85sVgdAgEnd
q2UnrI8z2QaETVE+ouosByteSWpUGLi44uWMFNlwqFhVQBHT7/tkExtp0kNXq5NZL5QLo3ePf2dD
YgBYGfh34OsHzra9olQN7n8LmRQtcjbbcQDMnH1BkaM3MFlGgqdx7hqErYg/YF/6i+No6YFtypwy
P3cEwgEYnY6Fxpr/z1W31dGSa0PjaKTxVKBBm+3/Rj8tm8uuu0gskEWCpXmUvltNXWbdCuH15rKL
qb7MecETETO5p6Bx3/VG5ZqjLfGA54tLJAUVcALEa24nBLdBOYkqvvmXSMpAt0FGOiA70+uOH7Ia
KAqQnuy8+Alm3pfTXj/oyjVQbjWyHrRnB3zgUYAJbpPoycpzz2YqTUZ8XOxJMXILw1KQMMpC7E3Z
UVHSsbZT4RC46kmw5o78Ffpj1h7FDCtH9A4YLt26d8X9MLSi9/SHVkZPyXTOrXh2ccHTS7BQG42K
3bQPcPG1tpLz+91Dps9zQfPMtrwm8wD2hFkzDlnVxokzvDO7vaox3852O1YBpdHbV55wmwah0kyc
US3Wjqqixh6U7NELKQGofEzqVg/L1bADN2eZvhb0kKqV9y1GituJhwmZXqNM+uy9rTA8h9s8dB56
z59QclQhIj5Y21nCgER9wao0vRSf2d7ntjwMQhV7fPV18nC/+AwnGTtuEkiiMYqfaFFkZaCDp/Rn
+KdG07BCjDu+RKbMAANjXRMXdLn95lISOJw49snpEq/FwXsvPKCt7QS97IHNIQdIfbAc1EsdSNw4
d1IwSxmtA1XmWcuHVfgSSifpYDHJeKyZUdGHHo6bBU6Z49MU9xZITwPj6I3n76GMMrdixWL7hE0u
1wGYAfuOXbe2fn3bHBNtGevbxafmMsWMrKte2f/H/Y/K0OjtM+nGHEaZ6nZ8N51eSplfFO98TLov
G5uLsnyj8S9zX9bzj65QlYKXY4ztA7WRvt6++qhcNRH9hUsmpInfHQxV56gBopxVqYKZpikLRn6K
C4jK9duBtpHLmzdcpjAsOoMcVBBpxZLF3UwY/2ogpBE0V00mNsoQrw9IBJh036Baxz1jv1NJIh9d
2CAGDCUFVrT9e15MGDcBfmPVQWGZYXEURkDuOvZEpFVClc5IwkK5ZwF6ZndU4U650iomkv+ulYcz
OYRi0k6rfyRQAAt2EXv0r+ZdmiA9aqwnctX4kbC/90xx4xDuA4cl+vTmPVJWvlG3lCeX5dmo+92p
gMHfLgDqyfssFoaH4G6l4KcTgJnPyYVm7Z7S8WYMUIfn7dPYWJ2w2eLtsNlnstfKbJbqv5eHjZ/G
/qDzmkudjDmTlND5h59CtLnHEt9QC+iMeOlkDaRdnSbM7QuMx2QAk44hLIk2XYKVLdRu6QZXbW98
qhBRw7NKm96B1pjvW+6blm95/tW3yfLzhc+efzPyOHaws6I6Drd2nvplUFHpKIn1G/xHPPQ9XIMK
eGCDIrdzIE188x5yDKGRZeJO4S14cHzAyo7CANAc/JT0YjmieWfxWD1YAxg6ylX40F1m1tAas/6R
MYcI6vYJpe2xkBO+6EE1d4/ilSqK+r0o+R/iYugB6N24Ab+Lwjo3VgfNNT897+D1IeBuvI8x0HFC
lk+tLIx4ipTdx63Vhn6V2BwRj/jKUxzhzAgpePJ4ltjfDW7zUE+TxNQwx0UObECzaU0LdcNcFSEc
7q+ZdMSL6eHi/eNvFtsqUg0KLIf6jtGBlMsjF+/JCCqC7QZeoPteQcm4hJnR8UJfwKUUiHOjAsey
h6Y67cc9pIArhA8mJSD56h2C/iKyN5SDzM+B+LeGA4jcj4d5fQX0pebbRwyJBb2QHltejS1n0h2p
P8dt3lLLr22b195rBbqmSpauA2VYN942kHywtRu40+rciLxGHJcHq+GwC6A9h6nScrobFbjmx09W
Zm7/DNetO5ClOhB4tEOZ91BWWJnAy3a+8dtDPLpWdc4E8uIXjMkI5l7JVDObcg7uWrBEPZE5L4iw
gIfLxmpXzdCWC8z6O5Pr7iEmnnDXBfSjQJpLIiwUKJAFTXRSlUcGLPC5NqPjjY5SRzVWP5/cK6DM
kAlo43h4R23tYqQWGw6wrOF/qauj2u3c+FzT6FbGhQDxikJUZcwwCdR+5ElFCKVkecXp8pEwaBCd
tbjhSnlTHQ7zgVo/dxZWZy1g/2S1MCfEIPQqfalS6jcy+cPWWgj640eGXkfPpOKeGAH6I96+GeG3
dKoJuHGa/nqWPchQi6wgq3yUB+jaVObCzGezzsnrZbhBaX1I3O5Q36cNyRMrt+24IshOyI0qIBDb
YRptzEYnCDMA91Q9ejK0nujS1lLIAGUB5lBNdEQXs9NFfC2A0OSoEKkEUPrmEoNP5yu43cMS7w9L
k4XEsUUp3xqWPc7swVGo8vwQWbgiUCrw0w0cohO4wKRyqNFPWvy9JEkN0jmiHxfc7CR4QDt8/YNQ
K3OUbIfomqpBuv/h79+S6jd/Db1AkP7SYLGl21mBCBZQDWSBQEPiETSjZt86QPS2TN1M8ENgvrdh
mjIAXboSEVhj2td2C/E2Hz95XL99GlrKMYLca2beYph11U+R4k9yx9dFZ80C9T2l250gjX9d5wuP
VsDFAo03yaj0YTvuPdK/5SrnbnM0kUkmo4dxskuBCP/WYiz3XKH+MNOtng+8QnegwPOBfVOc3v+0
hQVSGYkS3GXf7JivRhlhaeJYXzeJ4CA6+VBFZXg0FOagnwmxtuLUXMRBlLrVb8FGaXBnFq5/64ex
IV+l0RqjTE058AETLpaJ9SiegMeroa0dxuYHFbqp3O64AZw42VYDlwhhCA0GeCjLnRM4i1KCMYz3
6ADqxgO2t/14HP3xxj3VIXE4Vf7XgKUG6k9qOtQXW3yUGHu3RQXGla/eur+FRSuCtrqE5SeRZNX3
+Ao/hGsIjEkLFGN3qeKLodH+BpnlJGrjHWT+t++LHHvWW9WRD/oi0//F0caLJrgCvoyspAhjKU3l
8bc91HpILuxUi+0uyhB3N1YIMSkr8bpZghxpjG91hUE9GBGmU5zwHkGsuGchIc+rr6Av9DTwJrGy
zmScAEqyc9J3dKLYteWuhjXuQ0fk7wXYThpwb4bdTnh22lzKrsp5P6C29pqHjYvqNCXGg7rxHa2l
NLYCBY5vDMdbxKw7lIWqp6UffDAQZqivWlCL4KRZwdapYRYg5btWYxuYZ+XEX3G03wqdsRQ5d4wK
6SDizbIwq+JcYPd+YXkmvEgf7Oa4alAY8Urouwl2STuDkHMpIBT9LoFtbCoPo0p+T0P/Q4al0GdY
JgfByWD7TzS0mcWvrGdm/Llk51Kzlnm0gNG0XlfQYgbB5cN7kKTkwiExm5xd+w4eE2NUkNq8rSkE
UxAyQyd8dDr6Z1fXB/W6g3NllokQNuDzVQLkNuXpmHpy6gvygy5E6ZmpSO0agjUa/SheetqpwNk0
eQsDkNmsAzyzN1Fb6Amh1zCXGMQMtp7CtDt0d+6KceANab4BTFMFkN5p1lPcG0VKzGqnsV9YPiNo
XW15CBYEbUPVXphi/AGk3jz9+SbOHoNNhYbLCoolGQHnUDZHHVTT3z+qhzSdL0CjCK04HThDD85Z
o1vaL1xMDHUb6rYW4Uuhj/Th3694/olQ0/f2SDij48MP66FkSB5Afjj8AfuV6hwHn7GCYPIBdkUv
S2Xjtl+N1jvjD+3Z+xsPTcT5DWzP07adQIfZltUUuPvzPLAxRSl0AYc02ptVc5A4riktGDNsDjrl
M3eB9hBoa+0o/k4mUdvLCjzzW0OFySMVXaiAWO4UXKtQy8eutasE1G3GhHm/acM40u6HpuDJHslb
AQPfhKqyIwmr4W0hsXYObQ0WKvaYy0PSyYfmDnsqfe9fMyYbqQIHHoMwMbF2TQ1Iuq2PFJAIrsMN
48yslKu3AaYLHlL5EGO3dyqoNAE0OA5II0sAz56cuWaBady7SjuE9txhWyfc63ESk4ad887nQGxw
ac8w6eldGEkJYOdUQx4JKPydbmHzwxYitL7kWTfrhhRujrebBklDi66iR89PsKxy3x/mW6hiwiCt
pAeOKQWxAVtA6Fg4QbW/57YrgWeZaGhCDE1gTw+7sWBFzjDCWJsP0M7ufiVSBflf2L42/DCLd9zo
vJ0TNsR/yZb319eTlytoQSOfXGMuiu2g7r9oJMxTihVa562jN41pCPSGLYTaO3uAA56oN+sCJTCc
XA9NhfZ1RL4A5LZjixqONkBxxdFhy/ls+JfBNyRY61QV4ZkeavEDjw1KyEDfLVaT8Oyhsnu4PWbL
FURN7KQDrBafR0EEKL2xurrPm3yYfhYlOCOT4QfCvH+1WlJQ5bqg6BYFDLNXT62xtBzCfFLLS52S
YWQAWxBPeNGlBSrQXcjvqmxhgS0gUdbVZ3M0qWCdG5PGoaPHr+xtqwPWeEQRqv+4UhMMBzLMECtJ
iEiTWwjL/h4t1OMYMS42zC4/GkWw4rH4A8ntuw4jwlJuLcU1cEItdp+WpFW+OulOK9rwYMAPAgCY
OP3XzNekSVVSecz/g9qk5x+eAC8eMx/k79feE2U/J5fgTztnix0gfh7HNtqTOWT7QBHsNMP1fyGf
6gzTRTNhi6IQRMOENVfqOBJLkwIlK1AZDCmqeTUu4L64WFH97Z7dHi0f9cLGLHyw0KvuP5cxViLN
/Vl9DKUBVJgTAnjSXXGHQJ8ldPKRM25cA6K0XimKCUy4CCSQHq47RHvMUnPCEFSh8U+FMKHqp03l
kEbjULNoa+OrfgOq0ZIF3Xe7n9HaEZdk6/2xlWh2rLhOE70COJ6VqfQ4S+Dz6MXEd2Nq2j91XD6m
58IgMJKvZnW10IqlSBErJUaQ/yidGd2noxfFGHAVMONGmhezmJVdAugeof4ot2sI3fODASk2kCeU
LFMQf/7K+KaqYB7EEorXltUim8FUMW2OfmVDLmmhzrNGIZcWD0G2tfdfw7qsxQYrHrIo3RzQej5K
Hb5+Pp+3M2T1UMlZnmxBE85PBKO5z4GybuHRdgYEDPHmpiq0Nux7eTstnktPXfgfZ/fQx6RYpjjr
k8C0g3MLeY8R/ZwNEoeZ41BWCh1h10I23YZcWmHjqt/zuyS0iPYLrl1v+vgfw31uK7G2/kZqRVN7
mHQyWz82dYzDTkWPxbxACUzZJbfMmsZKLASpQJK6TeMiPQKvjmxvzjehDb2PrRJRF07Te/gIdxo+
X+3KorwEGqLvHffwXt98UM/mf9ynce8qCjamWMPFN743XB0LSSxgImOTgqMyT0lpH7q14e7PGbq7
4z0vEmLKoewzGk7Civcyy4KWn4mcAvPS9l0Vh3ZaaNH+YRZq1QyAKOHp97Z9wP6Ny+2TvNxQjcYl
8rPXJabhrRU6ObBdl+3F4BfIv1mhXpviYjTdFefkJqT/n0TnvmuT0zxFCQs5Ln6Gyt7VERJSPudg
gqhH4iC+EaH1iiN4eiPlE+LikFAnuSXqajXW6XeTE/B8BH8nG9zQJ9xAJ1Lq7lDs4yq1TbZepNu9
p+TmIYFmyDBfnka0b6Vvop90s1BYANMPDo0yohVhtBUXcLw/mtAblt9quK/mFaKYieMsDDSEtlJW
3cQ066a0nnv17laAVqGjtckB1pvtgXLF3R19jevfNeDkOSXOaOM1Id+cm1CeMYkHm5q8x+gRb4XF
g51TXvNSlGRkrYmxeI+UJEBFMEVtStzcIFb5pAzxs1l/KKFQUOo4vxCNdRWkTdfX6B4iCOCYhstg
jeiZ7b4UhxmJfw5l/6HfAcCbOEcopc343Ld0hiLT7cdxQ1V2C8A5vSiafa3hw88hv7e9tE7exyS5
77zSfLuP3Bx8hVp/sFFkGrMQoNlo8ZqM3CmsmooO0KkGclHBAdjV75QbsTtqj5s0V5eFqsdeIUGx
pU9V/mtmVZC/eNz7GoENb9W8YPQS+RYNwDg60qU6bTqwFoq7uVlhxPbVYoBjjwvUOEFHwgIpfwOO
vfYIW5qLe7LBAm0pUu6+BB6rlEWjR1goHDgDKX06Uv078M9dlmF88hGN3veD2kAqigyCVpljb1wR
MYO4RZPwOksDIQxZd4EDd4CIuQQIK3rezzEstwZpJI/mpYnXT5us/cto3IcHaTaoGREIra4hdKHe
CSYzw+8MRj+Y3wmvrHpCbAsVO4Vkekm1S3Z//rEalNxLeTUN4Ch8gUF6+z1r3uVpSYJl/E00aixx
WVOTbOwGab6ClxgBrnUAlsqMS7W8g6NEE6/gKFqvESRdlOidyHsMjqstJaTXLBNkHCVJ2ejOe/s6
jqB+BJwfVw28VtWmR9R1z1eXpHvGGFJiwdl/36qWWnUboejTOLxjkkA0FN3xd6CZNtsKUf1vQmQD
gEry9dyxvaDDfpwnai6maCWeynenVZTwUAKv3bvNSRZyIojSN87Z0MIvOzof5tFSZw06eXoGlB17
n72m5mrgGBDEfRBXKNLb26mKb4On+s5vpiM4rRImv98scv5HLo6KBk9BQx0O+jkdmVyMSKsYtaGU
J0lKmgoBCzn0oJJie3RhtKMmxeg1BMBrL0pDn5eCLRmdsm8nkv5MVcymgaC7CkmN8SJzYNT/DNZV
rv+6tj62xC/1y5pkL93GKaplWCOeiTTLWpN/R0JqR0Nww0sk/T/hSw11gho4yFFJGLNyfyaQrXic
DpGSfJ4Ni13CbQSs0Z40PdXHlw/jQVCLxjvEjSw9nW5BfFh0lHnAY/eR7u+SqCQWB8+VhDKBVMsr
hsPQ+0nU5l7rTFO93YOpYAlWid8XSGnKG70mJL+gM5ssg+uOqAHb6gqgnlPsWSDMqjmofFZ2luGU
RMTSfStrhWsjiDMSNNBSCdEgaXCv5/n1CSUdLa1bbbJGU2rhwTIRnBPqHmGRQHPT5ONtPVp1q+B5
LtDS7B78b8XuQnsDC2Vj96tuk/4zFnctiN2M5NSDEBF0PlAS+rw8arfv1Y7WjNiiHQuxGGsBydCL
tKQEn2rtFoKXaCCzL3ya1QJF80iUOljXROsd4K104q4O3egXtEAab26jSXolGNfFP3nH9UrvtRTJ
qH+dDxyfQBb714VtRXA4WCNK6iu92D46hWexofQvnZw/VmPDA6VUi8kedH/lWQk8OwAUaKHM/+va
+ndU/+rbCft0IUQM0e7ZHB/w3fIGkTZzJzea2ZaKNxF3XszU8ObNSC9p9Mib6qrnL44hHZsVIhcz
w+6MTWEm5zHL6tsCQy+rWwTmCE5TsMxKChVL3g3F+tXCfzGlN+zh33hyMNfQ7Yw+4v+NOrAYf+cR
gsTCnPZL6sl0xyM9ZdKr7bjuxa3JE0gpklKGWA0EAtJVB2Ekott8XRGOAbLkC39g67gnbxDyWfhU
mEW2eXelB/FeWASozQ73t9zXqZIwXMlh9BfypuZNHMvXWf/MqV0fDOgSavFrDaXpFNv4xvOPVIfB
7bf7wZuWoMOGbebCf1ciDbUvc3me2dufSUwRaJsnqzVC0F6WPrz6rkl2qe5Zr2HB5EeEeg/VoU49
RcgdkegGxpKzdb4XJuY4a5Zjh0Se5B2spRjd4Oj25hsuAuj8TbpHpeFSG71Kxokyry0vOzdJtbcl
RzLchd0r8L/bO/zKTM8p6LeZj/T/iQtukwAxRzM1nMXiiMqwbksMUQr5FSQAg8/X4QOqcfgcik+Q
GJkeXojJ1SO0XcW34ZGySEth1xyvYki1FO12fZSp3kmvaQcdWNpwtDIP4L4nYwK3pslfpm4eNbXM
PURP1jtvcMAgEUXykDT9PbZgdhsKPjWLoe8QgGJfS2JMIOWlBni/KUJuR7VbwUOeHO4U7+Bezx2m
qZ/KFiF/F2BLUe8ZlUEtWJeNhA1D+cKUwkOVp911XJ3YneFdfhLvHyKFcH4I23/LJp4uTREiwLVd
e42VEUlff2lNQvaasze/l2KMT68oSQj1FocT1Fm+AlQGZIXopiWQRF6Aoo9PZWsWq2TUn6J6Ar85
TF2w0scZjq+kdmaNbdEd0mkCKhBdnXnMBeTEMIZCaKtuc2f06b7uNm/E2cHszvijp5vsYtoG8Xso
OQWE8HOc6fslw7qy3BI9qiJFs1Dl9+Kv7ptpYWLyucm7qgzpazHphQoZE2XlXddmxwodZB34W6Wx
rCRoiYHZ7gWz+rd84PYRnk/atBqyO5mJVprMZGSjKyDaBfTgIu3iYXjMp8CjZuWvOYK+1rdu7Czr
ONKW9GvU1uvIveTluieFdEtPYr1V9SYmCFhiuFbR6TAQKA8h2dztKDr3WuRap+JjAtfU5ul6+4NQ
kh8514PdCbvipdmxRDBYstkd0ckcjkw60pF/YFvoUTrxgUKKjlow2jI5fVOCoP3y1E4wHWcZtORw
PBW8qQ/hwAbWdwJIn98+G1hTalpBMsUYrBlT2jXnCDtT5geImoDmuq4Gbw1tV2/Gb6HpYmumYZlC
pADhWfEaeWgVPU2Wl/PJWiSt5EEDBo8IR8/Bb+xhOgkSYT4iKL1lD8R/KstFanHnLRQieHFCTSeQ
w0Y0uyj5rurEyGfE6Jm8f8r7AlmahA9BpH0rOO+qUH2531uGFyNnJiky77mOTkHas/SRwxTgf2po
lNCKwZPRojTsrXNmOaVYU2capUq0wW5bEUyxqOgeX0RkLz+gZJ1UhCs+bWrjMBQymomUTdPZaIs2
glPZKXRW6awnDOjPHIFAW+pv4QsfKLTX+igJ0XCHaImH3Vsujjl5rlRQJEBBDS+vBO5DLM9yQb9D
piqTuz4VGMCxmwEtUrqgpHosMYn4zXQtugsjqHNOao+p4bJRNR53nq+NIwfE6HRMFf0bG7jqMeSp
JiEmDE9bgKMspKHN4ZdJLZl/E+OKy7v9TuERcKhxkjGLoGjV2WP9gUhfYzUWYzSrGCJI7uqfUZpS
rDBW04SuIIMHKVwaeQXAdw8ZzaOWdgCf294hFYm+CkaRD0bvdKDYSjwzlNUSJm7pXymoj5mddoCb
Iu6A5cQxySBdFH8qmdv+CN4pxfEMjlajJzSDTOtWSisJToBb3EQ1ictajPkqUdjMfeZLVNe/xmKV
DWiBDMYFST/r55FdjB8XPaqvUThFr7sULMrO3zhaXbXHv9B/5ZqcO8REL+3kD83fNfURlrzpkoJi
QHOeZvm9XQ79cmD7P0ORiag28cdFpIJp+/7/uGJerJxdmOSOdnOAYRqPkZKrKNorJWmgao09fyAn
J9d2ti/sOr6b2K635BhZnsnoWDyexGQi+bavsAVkmjXuBa5e0u7C4+mxRGTB8bSfSwjjCM8AwglT
xGNhNZ63ImrNYLeCO01sTHEY6YEuImEBILzKlhNeXXXIn7vLg1T+f/2XRiIzB0ouZDW4NuhCZ4Eq
nNFFTfMpJ8Gp9xAv56ZIWvtlVqPGD+KkmI2/243YwGe3QU8snDumwIY4RLIhmxKadWDIbhlfZPD9
kkerUR3MJarhoCogOKF3qm8hy2yEGIS36rmGw230p0ix5HuRw3Fcoy8S1psaBtjQ7By5cP8k2TPt
IEfDwJvlqF9tffohZeq3eXXl6T1iVNyDjReV2sv2zdG03zLi2LVSCL7+svaWU3XxzVukbE+hMxDd
7g64XUtW1xugP4EVNJxzliQkLFnNdJYxsb3cg2pmj/ndhQTM8bbUBiLb8uN2jRglD7f+d4kwzTHq
MtChA9TUR6DEgQV4BncUgAQnacpIqUXOA6x2v+GJ1VPv+YnLwvzjSPzPRjjbnfzfgAIpXUolMDev
E5/UylJ8ZsW6Jf4tl4x9U3vZUKqj2P6Fgz0E1Hjy5QT03pTrVCqD4gKqGNr1BYj18c3HDqeyw3Xx
SePkkBcQHs3r6KqJHgEM2BAOvFs9ORJF5kOY4TSIVYXpRBDhl7gxDzZOoO7XxOjhC1Swf0nY+Sew
dI6S2t+yQw3OJlt1beYHQXXX0wrMBBebEbz6FVkPkNtpYTVGqoRhY8cXejYNj91vqT2v0OAJah99
LNOFJPJu/E/prfJSIqONA5R5t1fGr7QsVn99qvzFIFMiScimQY/BR2flDQ3UueFL2zejTBh1ZeU2
UqxeZVDENfTfHg0+Jb7CpkN84XObFmxdLwO+FysVyM7t2VH4YUBWqdKLiplGBzEGBdt2Bw5v21HZ
JenDn6bwD6zCxnUZQKSmAyvl03/fNiGSddTUz+ifF89yc4Cmh3RL6Xxg/KqbUBrJmMpZph7y+jp/
uMmmQIMD95cSvVXAURepWGYdVkxI4Ev2BMj4sHroSZozPOak+jHrn8ergq3AKjCTRTt7L0rZMDjB
PSk/UR9SAC4TWDwHi5KOdcvPlaHsr2KCnxPPoA+u1AljN6ze9A4JgDJP9o1NZPzGvZsfAGO5E1eK
f01oSxUkb4tsL6d2nTxaGcO4R/MFaVM4WnzL3qODkZlsEdu0kXE4R6p2ia7pmBjMRjRIP5DjxQeh
wlfcf/93Sn68xVe0TrbTyta8NFUOVW0xpcbN2nC9Lrs07C+ApDpBowBdO7Hpve5XxLqh51I6OLnf
dcaQ8u5V31SvZ1RipvkofiGezCPLGU/uj7h22fqeAfxmVaZ0bCdm3CyBuWNnk2cpAI00Fcn1hLTX
B+FDpVA7GaxEK0mJYQzQOyD+gzmR2LhSGfWQazseFIwMgbXf3L6UcBA49t1NhMiC7ZF+qhlTuZXE
Qy8nyWMVjHmObrxXbapsRR12BbJqifLhZp7ONrSUF/JRQdeb3EijyekuOznCEz+/XL6KemfE+8uf
CaPjcXcwNu+JXZQ/1+XIy+2dG16CYsv0HF42dJ6TDivSS0e5XVZy8sXpt6EJantws/2pGc1u+bfv
dBx/PgMWDCnKdA5cMcEv1HIEozPTMj4HWII0LG2dOT2AsvPoirGWSLzdqt7xwQ95Z7Wgrtf281LR
ouOtxGmSYo8uMcfRahC4ochN+ZTKk5DMnLKA0XcozOf/7nQH3ENZDBtfIEBl0xWHUIU5ZTxb497o
5UO1WBLVknGGOwRZOcNMKPE0kQOb4LDDo2zHqqnbVMAEKQwUsKN92rnE1zri417zSi3Sqah/CHXN
PAVMfy8MsrmUamJiHD3TXUq2nqWYtlmcXYvr9Ok4UE2ROa7OfT9gt1z1NmkFG+nuoSFiNrP67ZAW
DGY3wtcdCAgB0vYmxqpFK5irivo2MHt+06Lo6vLahoOqNn44erstYF2eA4CvUYJ2YSluwHS+w2SP
ovqYU4U2U68e2OtvS7FRLdELghsJS+kmrVO7hGS4+OZnRdlmgDDRkSa2qCoATkeCwjWkjIOXT8VM
3YbyLFxHayqXbbwjuy6eJc7fo98T1IGQ3hYCb9e93ldogbcspwMEvWoe+JPdG5l+1W5TatW/9Vc+
K0QF9gV5eQUkZMOXuaPkCLVCo9Gfu9VyqvsONmO3Bn8sjKmgE2vlwZaThBKu7k5ZsJPhT8EJLICq
WHUYPVj2wdtGszy4/hUEiEV9jcOkAr2HF3ogR/lLOmQceTrtgxO5xwC3TVQSiJg+X8aU+kpHGIVg
fvPgFoDDwwaQHBmJALuq0IaO0Wn3/1VwR5VatwwxTqBX3Tv9wzsdbiJExSGA6FSWzS4BCPKvtHFd
LcLhRPa0e9PRuAJqNPDtdiME212OENj9qqS515j6EGdsT4oLbpxavoGyzYRGaRMffZpybpUZQ8zy
q9NQfftGnJD8TbkP8SAA0YssqJ6KA5rC+gYVFR7RDgaYMertQkHyHC7/MP0Flyc7Ym+wdNBfkTtd
j04l6rKma6klXejYHWw3CYkc4B8cO6OnKzv9bueWph2Pi5BGrJ8nUOOvjj24R3NJvdW62kz3+S4W
MWMZrxZC6/0cr8sbbP0+ZUuA39zvSRgzia/Js1ZQd91dfExjUm62zAu0g7oc5I6sTPhfccdvWsck
LHN9X7XlkTltp6RP1+wJoOP/f/3jnJn7WL0ZG1XWMgXYLvMCIlrpWbUg+lRZzZaiLzXo/+fF3oiG
snBPJ43gsraRHrvSWi/UTgu0edE/zWMdOMKEtY3XES5a6SnP5YbhqsJk+FaY9h5YRc6+TzCMt9D4
Hyls+C7GsxwvFz5H7IdQVDrUdL292Akb3P3gjnamPdj45TvIx9Sgf4vjTmV9Ev9QHizsttEMtr4o
jg6YScoK2MaC208ScnqDYpd+nK94xrqaAGerUAWWUrq9XlvRODoltdot5bfP8WtGqnBfLsmhxaqm
Nh9dNkHWeixAKiEdBN1CtX0smB0DAKu3vVWyLFOSCnrkS3lUXekPpaArgASybJvB29Qy1NeL6IkG
q0Rapz/N+n3+8Ndw6RIayWjpPz+Dp1K2U2nZDC1dZcP5dXBGMUdMjk22ls4nUuMEjCNT1D9p8nNw
3FGp6sHisNymhnTYYC9t+oAtfGTtHb+pG6mXcRGgA6Q4W0v53SQzq70qQ7z2TxVHlpdOJCAKEGCI
14kVbntqi0L8+wKTgxRTb9vOSSyMrGGtZqkOVob+DDLhNLKwHlxuJbAngndPcId4ptnkt0Hq4Trd
paESIlhscHAV4k0x2DtvzLgTIjc1OBFcUSbpT46c9zADLebli9k8Ztvh9eeoyPzT/QDXtv9WAeSS
ZBEZoiOd7NBxQ8KQNi9uhx4lBYmbVs3l0BBSFpenTzRqt9ORQC08WqzYp4t41l9pBHv9HdRQXeaA
egscp7779yf0Z6+ZmlyA8Uqnx8jdbxzKjjQVsqoDIy8h2uV9+EySj3p3GMFj0gsnvHjhLNpvszVG
w4466b4VYOvLhUOlzghRghrbu/hdu61Rge4l0pS37cUWN0F6LXsK5KDyjAllqX10hywWh/Bo4GRv
iFMdLcBYjMClYDMVFW0ZgtpX0fTKxbdjYec6jf8/u5bSMS389h0MZSW3LCbGzu1q4fF6styeuUaQ
77KuWmzIQieL50bh1u2JW5LEgHsgYkUYveETi4bwxGvtO5VBdmc0TNooZ12qpSdQmWca/HVGWl14
F4+ohLSnH+esVcwb0ddly1wSHGWZLorxploXKG9WdYsKW9WkvWKQYLAq/Fsr+5lWEXxCbDd5+sA1
LXeSOrhTx4Ltqp8qLfx4cHgXFhHRabryftIhkefTZ4oJxD006pxRjJZGJQjyZok93ICD70D5cxnJ
hEFHOCmE6hkyl/ZuT+NHn3An6um40ZLiHnRkltIdYGq2FefHv/vG5N84r+J6EsXsJTSZnc2XK9JE
IfQnHYcj59IJGhrVe/jm4kdVdvDu8hMdCPMBAp26ogA9DxjOF7dNxtIkLT3eSthUSkQ0H5TxS12m
6UbVlTzklx1s9wS6hRk4/UzDoyT5XYmR1evYOVUI4PTQwzknDq5MType6GvvbOTIm5HISLhcsJ+v
H/B29ikWly0G+PCEKnTkw9jVrzaK1odh1Viq6JDREcpiCHjCw8OIKycwYpALkySK5CfgSebQqmSU
KsfHPmXz3xvVhvj3kkl1QCMw4cafz9uXOdl0jWP4SbFcCrAGprBJ3Nppe7BDxVItrlZfpBwnKwQ3
+GBYEpBVeiT6A7XMAmPyN9BPhcC0fV3rpqSCjz1cwzylm6o091vSijzycuj/1FqujqLTSCuB/qo/
pgyoVGhnem+eehhWiIAvHqESKgjqQXZCX1sHk8S+/mHGP8CM6T0/mYqfYoW5x29OZ++2vRgZwrjK
UuOfyiilNlw8cJ8WMAeMpGOKRmGdrBsxMASN1/vp/q38DKaL/DSYrYpfZ4Zhlfg7tM0dy5/3xMtG
OCE3huCFwHw+c9ryVeaqsSPy1syTqmDoY+OjdG7+tXqVj855oaSYg3oaTywp/jXboifFEOovFQMg
c4zhnlC3Vp5c9FptyXRkHIIDCVu2enqb5bV+zDu+daUoZDT1obRa8bBGEHfC0vL5XX0CJ3x8jvl2
S+c6uKL/oh0ZnVYaBcb5GmbVwPMTyv/8uZUmuMEFhhXSamBl4Jti/hBAW7KF511jcmpt1WuPg7UW
Yw7qCP1S0qO17MMUy0SSu60WgeGsssmZ9ZxcxsaX61OccmoZ01reYEy6XCoosK4Dfl10i6qhroVk
GbolBJt87t/+g64YPOSOH11m+fQFS8gikvHaFFHOuWyYmgUeUqVwgs313dINZ9S2Bat2jEEV+tZr
OMdE1BqV73v3AQ3eS39W6z9iGEnYa6PafrmycD1fYwcVKS7ztOMteGK/FWtH5yZgvSHN3U7jcJ4O
KtorG3i0PzmfM1PDZ0kSVbb+t/g4wYYS+NrCNUi/+JKcgNodh3ua0R0Ic5Ja5WyRtj0c+DamFA6G
ex1Ita7mNxve3ALn4GDXBblkvw8TeN/kDwqOm3hsCHebegwu8FE93FnJCCoMnVmAs0s6OYkCQ6nN
fOph8r3gTgb/rFvR0FU+hbSduOfhGggPz3NJp5o1/IObwQ2TmWnBeYHdQy5yqMcTZlcEMdIwa4qF
uqQY8KkFPX0oBhByfctb/sXM/94dDLLlm1hd6j3uddy4pxNS6mTnDgEgq9yMiGZzmMVVOD+DtTW0
cqqRQqstyd/71UXxw3sISS4/6Zlz1lr2PmayopGGKvfS5if2Z/DcB3LhZSxEqrITWaVPEXWRdx+U
I3ZWjYUL8skHzvkf2taoThVmo44CLQ6M+PoORDU9FasKq4P1+GBhK02cZPnxROIPmkTZHWG1fpuv
N22iHAEtRN0kSPtBrSeCUYYE/vaB8JMC1afjpnGmrCEq1F4Pd0+/ngLMl8Ey6IDZj/34P8/was+U
c7QswNEsgw7qXQxUMnoa1MmDw3vY+c9cacaG2kIZA9DC7ysGW9mX/zR68RHzdnIsYPxx6TLZg99n
glItLKEptork2Ca37/Wlyk6gnI8SfQci4Nkv3un/ZZn1LDOM8aobZN95r4eEuwii9KDjdoFRtDYH
dtw7phuQEaY9Rgok1X1SBa2IrWPoddlvPUiW+OGAD9qah8G6I0F6N6Cb6PmsLGze+CKOL4e14bAq
OAmeKbHkVEyed2aw98Dc/QU2AR/CmtzbvpiJm4YF+XQ7gOhSK0x8kk+CF5iE1UP6p2ndzw4V/uSp
UMG1vV/AABQKmKzhV40su/XDjnRMPUtbajrGASHMOKCaPnGCUhbmaoRmeRtW2s5vcSNo7Y6DA/86
qLJ5xD2X++YZu3zwK9kfXrAK2jHrxE1f9IcbCiMim0HQSe2PhFVGA7JELpQA+ttAMZ37LERLt459
2QqIEqJP13ijOt/8wNoUTV5+qbav+0FSe+4NRvYtT77+tV+ke8wOcJckMo06gTAFbR1LLcQZb4WY
nwli21Dn2h1EfYCZzyxuK7t6tbXh+4i0cwcwSlgWwIzQD+R816dIGVMeYuT0OJUJa6wNuHLDydmu
8Xfad8l+X9mMFPr7mxRZTvinBBMS5fHOYnCt3AFj5WxRoyB3XDyEqd2NwUN8dLgD/3bHyf8NA/UM
+01RqRmLEt0+MOqKLGOJvIFYOC4UT4P0FAubij/jLiCW+aMWLhuPvHqRvKUNGTpr236gBeGb8br2
VYtohxbLAg4N2oao4ZkS08QExDn3a6aMoQ2rLhCqfcLvoRlZ28ANyy/XmJJkIw3r7DiHbAIxsG45
iid1AULsD84idmyturFZOyXuyrWf5Q7yXBFw0OvXLs9/yi05z2j8gcAFh0uwA4gS7ozpfrGFCDIL
vBczFZyizLyD3ORrTdWle7fsomrL9ZEKzxYlZcka3IlWP2kI9V3luQcV0Q1mXnW0L+l65Ui0irLV
h1Zd4UO1VQg/iBQ9ZDfcNhzI0q/lJ4MpOCLV7ZZfgZrpufxri7bSfYjmsuCwXLb7SoX/8+2TRT1l
a7uO+nWo+AA2M3LwizfNGpNCRWu5waY9Ce7EUpWHq0gkgsldw1Fu0jbdRCTJQzMD5VL9MLNQ2lQR
f2RWVd6iSmrAp3K4e1L82+0i7x/670QNJPtdi6ZDkINKHmns62u3TbNH0QbgJf6m75/Hdy+/HuiI
ZnUX5Nfkwt7mJNt32181q3SDf0/mykAYNcjQlduWJFEy4L76yKK6H1mCsyLmSgmz2Hu/P2OTcqot
Vr3fZu4gglgqcmQae4t0geS3k6YeLM0DZACSdq3G2LeqRqhQF6wA0Kp+aJkTIUtWXg2d/97/L7q1
WCUmaI374M8j5vVyTKqruds2IINaW1RZpdnHQ3p2XJCHW5ousXpe3JiXLeo2odS1nYL9TedrA5gy
FxVK65GTJ+vWY14s2Hpex5ArXtVRRKcAqGnR6dMEEtM9HMZQzmum4KIfw60z+dlgbIzZ4OiyFODi
n9cVLv2XFOQaqbl0uaM0pAZ9qojOBJxF84U7ewNS+/MgjxJuXtb+lRueM3wOz408gWnSO31NXIKr
BYsx42PI1hmXOToqHUZFxDSbzV3RUTJW71/kvqiaaMGhRNU1aaq9oZrGvkoT29qhnzyg/ZeE00rZ
1X2Ux5zvaCpAy3KD7/RV4JtZYErxbZvDMJNUPwRONSoAfx1+tCaMTwLqnk7D4YYIks0gIDlLMSh1
NhL0z7BedWydg73HllDSBUMgSRkUnFoDp3YsBlFkOyjOOrCiR9Nli0PFr+T3JfhUu20D2vmXakeV
Ic8l+E3jqnBECAncanR6YFdVeFE1CPNcp1nNtuRvx+uHmSZouJpQ2If0YyximR1PVEGzT5LzGLzu
0+CFz/NLH1qYOe8FZN4Mt03QHybZ1WR/GNziEAmU4/j9SmyILwm4/G9mOcAOb4yAK1BBnOYBFA8s
R85fiZPvxsw6iht/x3ByYCkYjuncytm2hgqUCZwbfV9NLKFjIHlvzFWNlV6h/TjydV3k7fU4JQwW
eEDvAJIlUf2njyo++Grf7d6yZWgLfQQIOPHQwlXc6lqmaNkbQuY11nsW4cGQ1bJ3pYUs1cakX39E
W9j9lFTHHj3g/Kq4bfN/QOdHo/PyXCDZ6tEP0zpQiiD1mr4QvW3oKVi/0saLCP415LJ6C+FVrDeQ
UR1de3xeLADAreqbGolSiln2XiB0IzyvmQao7CujNOsZ7rEORz+USGwQ1LcD7iKymWY4DnPQC2R3
d/WLaK7vz8aQYDpQJqzqfIMu7nzS07h6y/MDN9HekVUwwCN3dBHY1QSJBLi3RgbwstT8l7r2nr9y
kFcFnzIQ1+Nncxk5/7p6c0Trar2ExUJUgQ8oLUEHLO7LvtIk+HcPgtse1gWGO65mEB3g9pwlYXUY
6JYkTBwlMmXFfnloEkYvb8lqAvIld5mZJT2Tyecyz+CefkGUimGgLc+d8e5zQpr3SFo08Gu5aJ/N
FXIsTgzYRFSPyMgUDTQB3mspHdcXZRHndwMjA/FrB0RT/nSrE6uY21A8p2A2QuGlUc4l0PmJxmFc
Gp6m+IhpcH+0xkGxSNSe2Yn9Au0xMw5ta4BBR1qK9YrIq+rJ0l53coXnHVkqe9aqkLhDhxAbaiSG
KtzFpgJUjgzA8Z+Gt3tnIxWOdsgq6tYkVfAFiSgNfgY2zHKAjucTz97BiYS8vytCJygUd0SUTrQC
uY3d3bv0lNR1eeOD/rhEIWDm8HIDXKLpx6itAVqBBZ+N2PCrjrFhQb7GemhT4v/3gsCYX2wRJLzt
+k1SFaLCZnvlZTBx4MJjWilxt/1HP9r4k5BwC++I3FXvtJvewu5MdXN7CpFqNSmdhZj37QM96afD
9GWfnp7N/4i/7eGvgMWY2rR05X+Ak0z7mA6bNPH2b9Lv+n8azfKZK9cz7SJcLgTkI1hJBm1LJVkw
z66/2nC1Yq/WDo89m35fpY26OlfMBMcYkptItVT+c5ImI7nARFK9BM7BQmghKvlbe+qvTM7N9Rpr
zijKvtpprV1ufXF5le7rDoPxjE/TcNYzqCOJhFLK0xftI4u8QXGxaDr0IM8XBT2VUHypzqOsqEur
i0Kg4yh8jhWp033sAs9t0rKS2T2z+NApyuRUHCtr2ZrFHqWxz82tL7DFUchuozPUfmDplufTHgkr
jKNZlr7A2j1wcloUMKtwMyBvbLAcCkejiuut6lqQEZ+0ZIN4cFT68TLJ3PxhD796SsHa7aClY7DI
6dBkdU/oejHz4oXEyb6PjUHKI8atDCqmNtxgRfea1hyWHYTUGF22KkXpQ0J50xNF+GLULws3KWlZ
QE0tSlJhBm3PaLBFaBEcvq65n+Sl0Djw3MixXiaIDSnAZVSH11sDAf3vpY4BiUmGqgrZ2mFB508h
V0jKWcMLHMLptm72vu3ti1lriglhalys2aixEFx12VN2jm3Nlm7lsoDqD9FBOgoYeP//krjd4Rw/
V13mwyDEo9kYgOXBUGcFfAXoyseaKgM/FKWndSWsR0Sv7DT8GyMyeKmupH37eWlSjtCyVLSxkA/m
yi01zEH/rHN5dFlXcKZe1RKF6Q8X8wUEj8BQU6uTIqsHjJWqlfLCNhoL056FtQNO3K4UmJF68TE6
6ZyhULBhz9etKG64yty/CHLggkZ18FkL727r9flYGvJNpRtcFAP0rZKfxzkXg+C22/VkjcuVdiyh
ZWWSpGWynnnErPHbRM/IHLXsMbqadsvA6Zy7/8WSdLWOEKNXMWHWIZxZg9W09kAo+lGSLfSkFpYb
6r6lBmbcs2xDLMlbdeCzt2TOUdO9hNzTzqygCGQdEG03ufykKLfUdV+bP7Qg1lgZE2JWCA+1UsZ5
YUMhNzv6M6oZmQ9G4t7hA6vXGN4vr62F1n/vtjGkywClDvhAFa5jUPDvZiDXApmYeILZZfClmJRS
6AIbJB/KAnarCkKuapMDH9XOKMtOsrLiJYDLD8GI1lnffafaCjdFs+WWZraHqd0igdzmwFTMCYEz
4g27CDBzP39Mm11fgeCC/W71P7qmi6iaWCmqQ//9JBzo3fogMUacTltoZ3p0/O9/ZFMGby/2Y1UY
kjx/DaFT5RJ/K1X6d/XwVu3vpnDsL7CwfejZEPm2e/9d14uQH2Y1WxigMnvfIhuodLF395oC7WDl
td993F2g00f5hDT6+WmOzQ47k4g+JismkHK+QQh7ndYO4e7tg0BqfS8SxyfSggMS+Y/16Ey1M8ce
RuO5oT09BeCZVrNhWopAdjdGqkw5nIKDfMF06x2es0oqkOND1rd7Po8YtjvTcwioLIjYNmDYXdVd
o8Me3ABoYmCHPt5DJO5UcfzsAYeGiXXKfub0eUwStUi/7+OtK03Ee8yxjvheliBF7ArnpIXka3zR
M+VFd+yCyxJIxZ4/BZ40qnnXLAbwPheHfZEchrgJMrffv1gnoCYfh+rgyxAy5pFd6LzOb/6yhgMJ
3RHwJI9Jxxb6w56NXKvKh/FYSUmlFzgcOd5FW602xvg4XVRjpC0oRPb2WpsDCqdeEW2gFKnXQrzX
LPkhIH7rzAcjFKRveP0oyfdFIPJUw5bG4F92jOPd32D7SI9Beil+++gQp/Rr8IyIaQVZmtHWS5dN
Z3ks9RU7Ta5fqJHia96OboBWFeb99DIHagABNsVmSRjSdmPGJgv+RWZa+iE3Y3Uj7zsP4WVHHM0n
SKka5Drae55RoRVwUx7ePSpbdlrECDa+W/B9LIxK2esDzcTqRoSmgyK4sddjLyn2+SxUjkR7rMyk
83JFez8SQs2ahi+H1q/l7mlwaoS9BE4hGPLoEyBfW1Lck9djjUZw8gjiiUZYnvdL4yoioKjDz/9k
NCoY62Jx+TD22kN2On30vxYQRPZQfBIx9J20o/r0nvJkaFYphwGfzzK3+5er6a+5p0A0TVUrDa7A
2XWv2nHPMVngFa+yYY+rmBODfFQRV21kcCXlnF5Kp8U/KCp75U4QEp7iXfYAel/+nc6uTtTu+0nk
u2GBowThk2lTw5qVWTxOtqtyoslTDy+n32DWAEjoPWfQN00w7Rs0IQO9c4VVsLkyPRyjDo6p538z
sc5HjjeUFXnpSyaqw4UzmH6HFeWMfFBg0fMGLcijb16snT1rh2ywQMsfv6uaN8HKKkamOxVdF+1B
E6kf5ThW5qZ8086lDnMIveVdbJtr8hheyoiivD0ZfI/lzIYWb9mQ9+vBvP/8gdzcdy/0ZFQB47Cy
Q9Gf2zKbrZ1ue1Kyiy8HwpJ3+n6E3XdCgHsuav4PLuiiW5/5CESuNbEa6UoPUDz0fOgk8Gllv1j+
p1eXMa8QEFre8ljKeCl8h0r821CAzgaLEJaaWPu70WdzRemZ8nMv3LMSbJ7FaQEeEwMNACyTehGD
lqY7Wz32BP8h8uJfqiZ2PfXRAynliCxt2zNJcHV6m+rVfMy9k6OlEhd6ZesFNWIECAw7kqBDW8pt
B6D+yygv6rgDKe9V4C6ugEe6xPFiBmFEkdxsQBmVsQkr83makQAzTVMNacDsGdDQTkKGT86l/a5M
AuiZlkezI3R58teY8cXjORJnVIbCoLG76SQLQLTTlknkVJhjc103xxPtEc87eb2x8E3KMYGn7gIV
8rI+QWvJh9ULP2ntSClF3HeBN/Oa3Mgqt5mDtqUq1x1msDA3XfjRpO7/OF0ELzDIfTKKifbaMalJ
2QW0g8LLSGW+rJPI35pobCJc+XZAwdyKS7f9d4uzVpgatZchxGY76Up/dQk3roUZORAMP4mKrkb5
znAYJRaP20ahG+sPmqaK4UMzkJuOPqd4DL65uhvDQmzztLpU4MropJn+9dji5GxbJ+c/NS2ppYuF
WTHTX7y7/pEFY38aubh5InT6kw8XImuRoCL4huvlYd7UZfi711oyj+02B679XRpmDteKQUriTTPh
pQ7BzrP6n7cAFywhpxNw9iIKa2hAqx87ZQDS9FJDXqCIxWOVHY4VhRyvpRbYf3i6NQAxP+58ylz+
pGBJAiwUiRYLj2xjRqoyfIkau3srBOVATyuP8Alr+6u5uFHfAR5xQyYCnYc5Ml1WZOx/GJTgxWhb
538I/g1umK48zX8WCAUqKsKsFpijoslc3ayWtQ7BkCn/kYsctJr+ux7mUirlsvZ5QJEAHWaLgY0r
p++A5I36HMYbTjvf4oALpLIzRCT00rD6Y6dTky1KvWaz9Tbb/jU47VItg4bNw7Zl0aXv4r8VSqmp
llvy9tR9uyI+2gkYylOTfGtTii15j5/HqVtZ+mKGzb3YalYeAM1DuPBDqHhfvxbh0ThOsD+D165N
qgq823HsKLWqvFAsUNmmAuXL7a7eE592o2ksHGia5CpW0MRjLaQ+fSz7qd9CXHSX8qq/X5hzjxzP
YctztgdIiqtPAV2jlEbaGVWIgt8F/ljWRIUTcTvpvit0MHLiCN01vm9SoUHWqI2sH/0OoyjhX8y3
+f0D5QQHJoniT2yJDfYGfLDET66grlH3GXgROd+42A3MfmCQkXZXt97lP02Q0RjyR8IUzr/7+7P0
nB9Z7R0lE71H8HHKwyBNlWEEcgLuA1afplt8LEZj+6FKmVVP3M5N2kZm7pZ/tUq+oDoO9nbq25eN
HPMfkm6P2d80qy5x1xLjTMmDg5MKiy6QIt6Xaa7lW7xDaQgu94D/qoS93w5T668BgAmSue7JJVFX
kGEbT5cswA6A+i5TUmdJg3UGF2puMXpCV9e5QNzGAJm5obXdof4Oy6AA6DQipXGbDwnGPiytF0Vq
HwEXTbq5mETkMOAUOrYU8q4xmqNkqVsIIL5EwPIbhdEI0qN3ChA426aKl+KcBUZWPmmb45o2kkQj
aQMMIvmSp4g6WUgzeVNu5YTcs7F/aV5kh3zCE3FfmLcIESWFh1g8qdHpjChCATjVutUpyQPyKE0V
JvqnkGzrAqT26ttmaiyBmwKh7iyOrLDPj3R4SqXjIIZJ8qtCEc3a41ew1vwG4PGVOcWwnYEpwryi
RNoHOzWV19gI3ZStJESOTnWW/C7iDg94p0cvsrRAErl2sgdvvaaAknsibygbV0XjSFJbjkiMig7S
gw4RqXmCi5glAHtlPQ8HCFYRMcrSXd1+qXSj9COJ87kPfQScNL9mp1JHHb874jQkYXEFplrxAZEC
s9bypqlE8hWBUtrEKzKbqVa4yZNtHLEfGvQv2UuqkxKzreaNkVFZeJhbGa21xn9vZMs1kLWhRjHj
ylHY1tEnf5c0jXEfXRNLqenMlHB7D4XwyJ5RBFSGrzh75Km9vgirwH8z6u09PQHU+rKBC/7ITD9p
mwHNmY5YnRTgAwzbO5SUjbXGxFGpB4qrXD6MqqfukgHGo9FnIDQHCuhZpj4dVByzuhvHtsqCzWnn
IemqYMfdVyaIOtUMZ/1ePesrOWxhFOjxVU3C0XoRQpMDqA+CbQCOJI+7zaUd0wZWTeTCxCU5SCBl
wuh7ji8HjUJw5WRl2qeeLuGrSzDCUXfX+OWnYMomQv3Jcyj4dc7Dmau6wJ18hw7kqmnBbGcpgOQK
iRNJyTdie2NzyqC/+v7Lk7NTj/wjwK/ymPG3+hCLlPhuWRKbbfDx1y5WXbl0I5MHLC1JoASbgh6W
8F2Bt1clCvMvqVqFp20rZZIcU/OclyxQoj4FWDXhtknyDiYlWFJM0OqGJnVgIe8R9j2REkq6ZN8r
hTeHCO1/K07fvPpIoBwCyhPQDH8QSnc3yn+ZwDeizIxfFijs+eGTNBgUibpUyX49kqdeWmbQVlLb
JNQef1jFcO5VTCROpRLP6j72Hf17frJLSNxc4Ixhb489Ec52rxb6aULTBc1fXq8V3wZ/O5MRG9uA
R9VBgAaaea1tX3ARsrDctvuW5/lDNsBlyx0igchEuaZ12wTPDjnnmYzXHUvzR4350f0SBPkmDU3w
/zCyYSrg6kpVHrOZmCaNuhAPzuZIsnf3itHYJ20SM78+af6lU92jh99yovo3D7Qe+49HpJuMdGWE
DooOGaDAuiE1W2oaLEPA1lI/8wjzB7j7rGv4OtgW84ON2m4FpdBhA4GVBy2rDPLUog/ucdByLqWZ
+sJtBY3yM5MZx8W8MvEvSg7dP66ZMAH4pVUbYL7Ozov6ZZ6vBiXH1Bjj/BCiq+6jhkqT8A9o0e6d
Vs2ElV5duvLomlglONHgW0I+1xB3dL/Cr1VKdFD/RQiZKWVtH0WEYTLgQ88wEsak18V1GpS5P+ee
cghwjuTA0Io3ATktBEVASuDhbtcbKapHHwsGc+VMAwQKqsb/JuYYJLvOrFhjcgpKJ4sZX5AuOLET
5g61gII8fl4ywwX9e2PUKd7ZGKqFoy1PlmLtBNtWVUNUsKEFDl5Tihhxaj+LMGrpfh3/VAMV2Rpp
yX1T1ZHCWK2T3K1QQods3U5Lc+VTt6CZ+Kp/kc+NKnvFFF3vQk7jMv07xWGUca6NDncms36T8Tgj
2AZfjlLdrp+xjuxginzT42og5/beoGq06KWTfcON3MpOyg/FUkaseXZBeegY2t+pi/uw251LNazv
T/HrwapDW1W32pRnpertd1FC9NnRae14Cgb7naQBg/GKZDkJcwFBzCBHp35RAmq+UaHxXDJiblYg
VYBjgQ+00BbmNV8a3+pitYSwGTu9A5HpJ9swKUJtDk1NC/Z63KgQvwcHYalsTvEwQAoNWHTXbE5P
9G6iFbwLs3OzlWEFPcd8kfD7n8x4X5ftLB2CqQ9aVHVsBgNaOkoKcpHnmFJCsN5Pa0hALitEZakg
smnL3iq7jMNNTsgHRW/su25VwHKfk4rjvnKgNsaKDWHlWPHTZr3PAe2PG57G+TWq/t4benhEABRB
Vx+9ldfOY06PqceXxU1wMdRgbNKgiDL1DqL2SpWjQ+RirA4/lZXmSu9ebXje14PbMTizXKqabeHz
KuMqz3Zr6OHewUBxVOHEAzmW2/x4iaDszWYZK03RAFkiLLKdUg==
`protect end_protected
