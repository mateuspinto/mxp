XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� �&)ƠB�$e��z���>����^WQ�ʪ��͞Ӯ�{�d�I
�
��`z�ǒ���b�4C��`P�ouhB���&o%Į����p�@��`���#���y��8OQ_=Pط��������!��AF��J��������ww�U ���+��2�0&=Ӻf�e�����`�o�6\f.1��l���84�� q@�k��/6�j��R��T7V0��1�J�绀q�-P�SGI�nP:!�9���g��V-��FA(�N��[#x�1kWʣ��:�ƭ8����VV�(`K���)�J�QSWƴ縇�$��苉������*>|������6�|yf�7&��hp5^Y�ewO%.�	�`V
ʂ�wL|m���h����f�Fɯw��˰;���W�Pm��Mt�Sl��6�������?.�p����X����A�+p���j�禤���4lh���k̅��䆴�D_�����O^�kx��ug�K�aC��������������X��Jk.�зV��s�쑑���72�9�:�:uV����By�bX�&nH��WH�+�������["�a��\<�h����.��BR���8ӎ��Xe�7wt�{a�^��Lt֒%���ܽ�]M�8呶xJ�=���vدs�p�X؂4�hmXw��%F�Ѫ���p�j�`7�6��Y������p[���)�x�=��[���+�1���%ӟa����h>S*��|F�f��B��1�
�[sXlxVHYEB     400     190���H�Pѱ!���J��"���B�&����4~OQBsEY�$LL+�`�UB��5#^
�F�Aq��BW�!\6����ٷC�]-Il4z?&ԯ/�vj{�M]~�z���CK�@0���ugֳ��獆��d@i�y���5q�u6�Jb�>��������.���/!RȄ�y��t
�f�;�`�̰��$�UP�K�})�q~4TB@62f�Rz1 
�(�	�"X*���<�f��ۧ�.��7�0��W��tx�b#HZo�|�;5΂m�Ůy=�>V�̕m��M9P���B?ʁ�P���C��/�I.� 9��#�e��K�i�#
��$227N#�C�1}�gh�gl���r{��/t�h���-��#Sf����<��`-W�|�� ���L�TvyXlxVHYEB     400     140��L�����`F}����%ej�y��͑ҩ����m{`���M����FӍI/3�؇�+�G�M�.-�p���=\��c��([7�W+W���az��ɂv4������r�9��NC��-�|�� � �%{�.����74�����w]l��;��᜜��]�b3qؗ�G@[�t�i�?xjN���9������cX'D'��#	��
��$?���ӍB{�At�_#,�^	.���6s�����
%$��`��ɵ��۫R3����Q�u�f��PLT_|�8HK%9�� ����4�,���2t�c�(�O!e1n�?XlxVHYEB     400     170H���`ɫ�ס�h�����{9�8���$,F����!˺��Y�~�]�m�e��(�zi X�
4�9pY�8ځM6i"��WV�p����\؋�T���7��e�v�KPtAV`�˹��D���(�Dgu�]�2��q#��,6c�&�_����Ńx�ͪ�Qx�?z�	��*�����܎c�y�c���-~���������zy=	7~D�f��/���vaC>�n���Qp�g���O�(��z⴬b���5-�`�q����Ԕ����x��%
5.<>ӳ���`������l!'g��[�w���vJ;~{����{zz��]�[����U%��aS���fu�tS�.����2�1�XlxVHYEB     400     130�|�#_��u˲��̑Sa1���)��/�7�	"���&�ɵ�6�z���N��/�<[�uᬰ|H�x޿�������ĥ��˦��{^%!�k��sV����T0:vM�U��.�/Q`��Ī�̢P_� ��u��YI�X�Ee�g�x����w�(��AI@�n���p�5��"��ye�E"S�XDu'�sl�[c�+.�1�����AJ8�n��<�X!c~T��i:k�QxrNbT(���CAkO�������@��&Ic��M7�EXt_���M����XlxVHYEB     400      d0ד)�/��l�J�0/1"l�'�K�b�"bvS�.`݂Ʊ�p�\�`�2�|�f��-hF�v4����8ǥ�΍�wx;�����U		��މe�����8\�������=_��5�\Sz�*S+k�07�w�򟮥��&�ӷ-��Ź�"�y�B���Hڶ������+����8���ĥk39 ��Lt,˟��5�Ɯ�/[0���*-�XlxVHYEB     400     130Wi��ϫ�@+���h��Q$?:�Ӏ5��JK�zZ��yd�2yQ��3[ʕ���"�H<��Yu��d�e�\$|T��÷���<�4�!���m/�D�ܫ���>&4;vxΗ8Z�4���.�m�H��x,��m�ƌ""���.��P��]��9�R��
7S�ݞ�����K�����vmmV��X@��>���_�
$e;������/�}����Í�#�8��4Cj��tsZP�	./�G�3�G!��י`����lSշ@��Ȱ���e��ڣ�(�
�9:�<�XlxVHYEB     400      e0�$m���X�,Z�(�pKd��
���+��c6�s���� i��hi�{7�bNCcWp%�;D�
M1ee�*&��%-܅�{�L����ę��������qY� �d��z���B��NXZH:D]�p�K����&։� �1����c��nR��Z���e�u�A'0���XT�>�o���W�7��>�o���)�'&�/}�C�j$H

_��)�,ֈXlxVHYEB     400     140�O�c#�5��iN����(���_��B 
%C�e2L�k��pe�Kd���f�\[�P#�e�v�6��:�|�u��nvc��Q�.�R�������|H�ߓGK���7p0�4ۨ�RĜE�ʾMP�gp]�y���̹�b���p����ə���+pN�J��"�I�
D��O���7d�6�iüf<��ޓk+B�+os�~��
%�N�sy@�ć5�ʺ��d�<,�(�����Ј�d��vp~���?E��*���/���9�_XɍM���+	J�FA��v ���s�^�V��aջ;��i�N�̨�W8XlxVHYEB     400     180t�P���g�:�0�MR1�P��5$f�<`�T�����&$ٴ���
��Y��;�Wxn�:������0��
��nR���!��!��:Zf�f*�XV�������3��d������7��f���G�h"=����r���vv�u����Tw�x�\L��/}�T��<���M��_� �Eؑa�x�xU�Kw.�X4J�[� � y��]O��g��&OR�vC] ��������z��c��n�8%GZ�%ρ!��>g�l���P#d������g'J8A6��,��ݻ�})�T�$��,�SQqU��#K��l9����I��??	�L4��TI0����ܐ�vh+�K�����yaMdb�C��"�mt]���i�XlxVHYEB     400     150's�V��%<*+��-��:!��w[MH�D�j�� �6/��[��|� _
}��a�������� �mRק��~��%��_iH���؎�~?�����V��|����Om�]`�S3ܳRi��O��eeW�`ˤ���gk7>�}XΊ��2�;�XI@?��	�V8�)'���z����y��|Y��U)�w��?��s����{'�"Mu���D�?��o"�=�~�oK�G⫡,��PjSNyjj�N��"W�ݠ�IV�|T�	�ptOP�6�(�	#E�[}:�&�ט�մ�d���`B<�L��5�}�級kS_R=�,��nz���XlxVHYEB     400     1603� ?��ɑ�}��ꥉ@k�2п��AgU�A�-�H�#n�[�c@֘w������f���l����Fʇ�f��u
A�~D_?�#"��qUм��7��&m��Q�׾���k��p.~�^$�?uӥ$F�aԖ"���>x�w@�F@��w���� �O~M�;E����c|�x�z��O$��I�OP�:rm�OND
S�H�PK��r�B־|��L�hƲ�S7||E&��b<ݙڎ⸦}(�dU_1�k������w��7�����+��O�{g�ƋG�\ ζ�u�.Ǟp����7����rƽF�,�!�ަ8�t
I	/� ��#���a�oZ�Z��"����XlxVHYEB     400     130��<��b'L�k�������>�-��*-��^ W��e�M��,�ô<rWi�݊3��/��<m�¯ay�o8����}���&��f����0��S��ڝ��[G��5��ex4�7�x�ѐ��jP;��g�}2�i��"�$�U�W���6Y��C��}�@��K$�[��y:`uU��2�p�>�K��@�=s�~�)�F��'F=�YX�!z�2��Y�.��S�C�C2<R�V	J���=H��}�٫_(I #)��}�$M����I�V�w}�0.ww�S��9��d�����7UX�I�XlxVHYEB     400     140�Z�ܖߢ��ݣW��	��֥�G���tqD�R��4`�wi��"op;�	�)��mG���� �t�OX�.�th=xt����u1����2c�ם��b!̧���Wѯ}��tb���RKI��Wh>��D�Й��C���!�V�vf��(��6�+�3�h�8�UK�j�U�o� �D���{S��U���#���uPÁ��C�{,��]dJ��C��|�� -�&n:�2��iDɭ��|ޕ��&�_�����a�;s=�}�e?����#�����t�^�/3�ٌ(ojiE�CO�9$V`a՟q݇/"NI�μXlxVHYEB     400     1a0��0�dZ|�خˋk�j�F�v;���7zs+JB݆1<6'��3v����'����W1��@ύŃ�6��8�
����ʁu�bl΃�.��sS�&�G�D�2e��W�=����+_��T4(�+f5NS�m�����1���\T ~���yra�H��Yc��gp�`R/�#xā�:�XQs�[�jI˞��s�,�񏽽ӟY�>B�����Y(�(���{9̮��cs��9�ٵ4���md�����V'�y��+��ɶ#�yκ�~Q��oq�p������1���O:NEt�fQ�$�
��TU�夣*�پh��"����H�%$�$H*��ݘK�� �/<N-�{I~�}y�Յj`��ھ��T4�f$~M8��n��:rE+�M������2���������� ���N:ċ��XlxVHYEB     400     120�n���>g ,��M�?1�V��^�6��}�X������S��I>l�6����m��F��zɋ7y��_1��~7��M�Q"hv�����ap? ��{�3�Og�����U�^l�W�֝���}툤�E��6Ea�K�Z��D�����-��e��SѬ���GAp���I[+R���M�b�f�|S�8
 �IA������܍S�9�4*�7�𤺱��XQ����<C�[�L{Z���Q���o�C�����Ve��/�U�����Y����D[��ҧ⻳��XlxVHYEB     400     180��v�����jd�,N��M���̲L�oH��(L�/����顐�D�����#�,��ֶ��@�Z��	2��[���T�g��J�v�`�Q�#�V�L���p�b�V�������&Sޓ��!ׂ�9���ė�w�F'`�4k���a�%<�l��)�:�/�ܥP��`x�ayI�YB���,�:RHs��i-'C<2ܡd�}���;�s��p,j'e�;=k�YQ�Z���a5&mR��5Kk�M,p6�k�9Q���@�?e��Q ��S���=�-��RP��<��D�M�Zs��xx���Z!�3"b_��ˠ�us�Z���*��'q���]|F߀� �2��w��ѐ�
;6YJ�P���"�XlxVHYEB     400     160TGA����-�;�nT��&�G��wi����%�ѝ��
�:��2x[��bk K2�߬>�|�k�3&h\;��ۅN�}fD��I�.�Xԙ��d���Tj������l��Y ���(i�%���K�2A�"���Ax�����j��z��D����K������#���B!�0ݑ�Y���p�Ⱥ�S0!\�EL�Y:��EW�,� ����w��3�KT}.�d���>"u�đǟu��	�����	\5�һ�]+��HfM�6�h�� �&(�-z��	����(i�]m����:(�yCw��d��L��J2������w�;�/@��O�ŀ�O���ep;,ꄎ��XlxVHYEB     400     1b0���$0U��q�I�g�V�V��	�4���r�C�n*�O�j/$�Ha�u��)�ц���l(�oD6��*V�;��E�A�A��m|�����T��;6$�_�n<v�*�2/Ɉ�~7�rۑ��f9���@(�@�9Y��09��$|#�M#K�� �[1�+�G��0.���1�Y��G�fw�K�U�U�u`�JT4XZ4���(e�g.����&�����Oi�ý��� �'�p0	;�j��	<�z��)�r����wִܵ�~'�@��o�(�ZJ���!(7<�(,zLL�:��y6#��v��D\���86��9^.<��_!�u	|����p����-
�˒D�Dǃ�Lp��Q�����ѥU�ўu?�(�׆"ͬ_^)���H#�����X�@�U|4�.&J/ŖѴ�+9D%�XlxVHYEB     400     160�0���"�>��B�KL8� >�v:dL�0���?&z1�l�)YJ�E�(=8��� t_�H�u����x�*0q�GQ��"�u$�p=7�@Jg�k�j͂�?�E �����&��[�|Q�f�o�U���&��w0�UL�wh�TxX���ƽn25��<�_�;�E@͹=4 m���=��/&����@z�d��`Z����I�3���2Ӫ�������W+9��I����A;�)'��m��
K����*��\i�����)���m�������<�Ql�4����]Dv�Oovs�@?�r��`LX�G
�@�Չ��,���$җW���-l��ĭ�����I�"Z�hM `*XlxVHYEB     400     130���PV�\'Sw��G���1g�@��kh�Ꞛ=v}�T�L����E�ж��
+Y����h��r�tW��Ʀ}JA9	+2�^�7 ᑕ�i�P�S|���O��h�/�N}�J�0$�����c 7�)�Q��a��V��25�)�Ρ. ��ǚ���K��O͐~��:����i&6��*rZra��@�BdƦcمә�+`m����R�䏤�3x^��Q��٩�I%"�o�hJ&��k� X �P��!Ͱ�Yw[r���on�(0̊�K��۴��������m�����6wXlxVHYEB     400     140y�~�e'Z�%���*��
Z�m��J%�;X9�mq��sS�����U�l�G�^�ȅ?E���~O߼���ƕӝ�T�`h��*�^:%�`�-��	�)&���E7־�����|�ם촼�h�;��T��,4�~���os��h鵘����Y1*����L��ἦ��^YK��q�R������f��гr1��P�;�.b��n�|�,>�퐂�=�u%Q�H�Y���fg"l���ky� �V��zjj
{�gEA�e���˵A�<'�.��fi~�^�N�4���==@Q���&�d�H*���2/��c��@g�ۜ����ٚ'��XlxVHYEB     400     130�^�Q���.�m�� j�_�82y�pY}I�T?VZ�V�ȂyM�g�DH���E� ���_����/X���z�g~��:�[���П�nVޖ�s���1�5�0� ER׻�{Աo��N`�{F(��l��S���ټ�˷Fw1�,���Z�gJƄ�"�Oڢ��7�+���7����_����x���)V�2�K�t�Z ���%w���+r���C�\�f��gVG���H����d4��˷�/M
�!,d�J�Q=6�YV����i�Mw���C!q�D����X��Jd������4q��<�3vװXlxVHYEB     400     140<(��$k7+פ�h�Є@�MA� ��f'x�I�#�6?��f�����c�nNn�c���K�v�&=�<���X*Wj<(M����-Ί`���s�5��Mf��l7Dk{DsO)�簔Jqi'؇�han�w�`J\Y��;���V��F@�W��}��L�@���{ܙ�̓��ĭu�:�JS���{@Rw�
� �Ai��Ї)��/�}�(�:s����ϵJ�u�N���������oP�Q8@�L�Df�\kC0�e��rrq������������C�6��v�?�W;q0�o[7v�<��ΑSЌ�XlxVHYEB     400      d0,}�`+����v;�|��}�3�i>��5K�9��7~#�)~O��W,L�s�w������`.�A�KD�]'�HJξk��#���Y� ]�`�t�8��Bz-�۪�Nf�^[7��MP�RXv<� �C�3��FS��"�(�5��9OX�v��z�*���Ӫ9�HIjQ��Od����n��$��2h�x�w|<x J�\j|�o�o��XlxVHYEB     247      b0�p��x�i5���:�����[���̖^��ngŢ	���@E_�鼴6�_j�0=�3iG����m��t64�Z/��]�8,���,ݏ��ݤT���<PG^ �+!��#�q�'B1�Iv�:/�����^��:{'�Z��Ԃ %����]�g���v��^��~ L92M{��Q�I