`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
P2j6CIhXQQoOzFx9MAmDpYYCu5nHMgDZHQVn+offo88nIEqthSXttdbUpWFZ9zteGxA67aIbdCG7
yIIfQsD6SpjUmOCJX4PiQjojx+B6q9LqD2GZA+OP4zrWmP0RCbSkqPHaUhhrOD66zkmseNhwqUH0
6ovpkip7fH2wmDSSWenHIUph9XgJG8GuqplbFqUHNhUKPuvIGJoSeUv4+JAcVlu6m5ftAZ+L5EHI
a80JJdg/6mk5MspLJoNuPdYsdgmbaIq7VGjvOQzyOvNzhmemP1Qu6elRu2n2mFeTkGVMvkNZxhTI
2z3mK4k9DAsO0Hy16UwTkbL9sfHDDAf69fkGDQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="dvoT6dLfiqtRHnaed74zWjcV0xvSjerpfEPZWq3fgKA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13856)
`protect data_block
CwGF4ZgBDvSusD9Pda8P03k6eWdsmmQfT/XFlmktazSnZieYZrqLptP1B8HxEIlbPp8P/+St/Q9P
sAjxm++vULQ3fzGv9GUKR5FgMsKxNeeiNX9E0HQxHtmrCPls9gTecTsSNCF0dF6czkfXDFQ0Hytc
/B+gR+f85O+jNuy4T7Ozni7TbeJ+ECRMvfSxq+LIFup1Xk74e/olNftdq8lFECmAY2UvvI3K/tjR
B/mRbF/7gzI37o0SysOhELRVGFXD+UACPO5/mJB72enKOR5oWgGZ+mNbr2ZSQJMnr7UYzQW0DDed
d8VSbK43Mw/KMmZcfPwZgflOL5vTnsGZeok7VCxyJrJ373wmpLR0ncdVWFsWSoJk3xrBJ8GB/txB
Eh2rIh01srAIf71pRqI/OsBeeN0Z4qfFsGMp3UGi5UZzX1zCqkIBkVWkIaG9M0D359YckUXsLpGY
oNdxbQtGCFi61dJxSgY0dWQ8FGnt8a4gwDRrRtkAWPI/2l+mzhE94fGz44q1OZQJToYx2NIHfvVv
QolSevYzfi2GbmeEW1bOQqSkwO8/2NkUBS7aw2jzTkO/+wwdWg1CLPxy10Bi5cOKTSUIDckuPq2E
C8FJUVTtuXznFmTXJpQteVGAzESrSQT7q+Rtc2muRxq/JEeSc2J4Fz6y/EPPtM9IWWhtut5fZdoE
vMT40qvuch1hlLhdOkTyWPLluXJnk1f03EKk+ftzTi6CvO/bckLveyqdvKiAq4nvYDPhDlKIfZsL
tEoxSh0jEIjd6UefJidAoqtyjM7Ki57nTeSaXL/u/K8QV5qnl35zKlIY/C/lUE12R4aAXjlbQT0a
036LuSjq2wFJIh6a8IhsJdswix6DrN49reD4EbgGVd7wsaUOGFSFvIGdmAG66K/ZiXLRrm8X+iGQ
8SN2VyqjGiW1tjaFTO799Uo3UYbGZYBJnzq8VdkYrxfTiaVRWmtYxsAaWqR6oxzBl53HTSUEXdfS
u1aTolozBP+YfZQNaSup4p+U6VpYQTomNK6qFwh0CeFAD6UG3zfw2K9muL/mt6KsFGHIbWEIrFj3
/H52wAKOsngt9r6iV0vQxc5WdjFX0csOYzeY9acubOtIx5/1/PqtlkUcTkEDkh3qiGUYaIRdK/ep
GPU3MvYJTa15AF6m+d68E58nCcN7bOPL+wo0j/k0TnbFY9rpvMCpw5FPfC7SxTsMmLJl6HQ4aZSt
/zieUqL2jPLE8BeMdUZ4J/0oXMO+1stcC2Lcp21l4pLWr+s0lDG3puJmykfBctXvqsslntMUqben
oIZGOJn73YXUqI8FEWIjOsZZ2/LXW0tCbGv8ZUOwwHGn/uhZ+vhjBAymaPpuW6mGlv3+oc/EzH/w
QZvhfSPMplt3uNWMnwEKYFPT30GkIsXKaossl8a0/LGvIUdEPVA3iumxLsoFdremCsm/giqqPkMi
NBisWT6hnKKiF6ixbZYOQHRwyNRimE6KEjZO0bLQPrv9vJ0yCs2vUWL9DzJfWudipfEVtbrq9ZIa
q9asZu1S7iCiV39KqJIk9mcUEE5vBqjo9qkJggies3AEg/otONTrr21M3Flyg0+1kJ8tZnuOGsY3
VxpIlquin4RM2rFV9wOlzOLc90G4/Y4470OOiQ2SYuHgVuo1EVfmtHFeBffn2dQCPMRxGr5k9cRx
j8k4HcW5c4CF1wB94qp5s8N6EJtnIZEpgogkiig+xDA7bgkn8Y5FoWGX1MnKHGtkMU/pdNQLLNoH
ovy5R3wE2DydWN8avTSEbg4SOxN6Z3NQAMC/H8hIddylNuhdJ+hd5GJDsEBMupK2sJCzXF1SDc1p
5eKtHP3KxnfeKJ1E0zFWzPRt0BI1jlGm3lfgy0eQMLW+z9F0mDqcwApxyKJ5KJrdVQcn6aIv/RNm
5DenYOlDxbpsldfvjM6DCaCe+7sK6PYYa676fRM+Y83QutqcgucmmIBIEvhagNPxW+gZpunGEVn1
5OVHy3VtQ1PJN8plZP3juoO39hKrYxghYO/SmfG+G/dKG3HE8KDIJL2i1PstclX5MRf1v6EG6Y8X
advrlyUcjs5t1GFwAcC7SjI3h+dpNoeL3j38TfBIgc2KA3w79oXAEiCkxVotqVc3znP73fzcA3AE
rAryKMx/WwBoLIATI74UR0HlxbuvRYOfoRcBITO34A/u+inADomskdq/4mpJ/CSQa/3sIJvsR+wT
H5R8G2wpZhAwEJmGY0XKu827YhD4/ldI6n3s1EeIwS9ZgaAXefWFeTMzcLToDMFwvblaWBFEK0Ne
jLiJisRH7QWJERopwTXqqC717khEb9gv0/+pICVcXnnncOF8+HW3iGN/0JHAiRPOqzNaOf1Q8xUd
Q/HfesEw73vS4XkSGp7X5/kKTnkIo+ROFZlJHYpHr/ji9z9Un5xDSWIWcGeXkC9iZG8ESYF1AhGq
CUy2x/5TqkQSKZD52mu9UUzXO6MxpbW8Z9RubBHNaUziFTMJdxu6KO/nFzk7mDIem5vS/C7pOM5H
0iGZgvPmR8cX02ETDMZh3c2PESz+RxgN9vB7mTjeQCWyWb8CqidcRu8cRYme7W/GnOTGc/IiKpE9
Q7ig2UH2GXQ3TCElsHz0DrYHLc3clcUVmi8wheWyCthN1Xlj3Lt9Mbbb8kUJMKpgCaMa8ca3bLN2
6s/NJXP1p2ZVUdvgPJpGy+0IU+nagj72ADQ4joyozDyOrutN5FyMjnIySvtGdKETLjOvub4yjzkS
FH8uu1EhFMs+fikaKC6hx49lFasD3/eznxAfX3UWP9jzxd3uXJg8vuKQXyTzM+9l2m5xVbY2StQG
/0+GGFtKQ1RnuiC/BsJQcQHOqlkg1F8KsMQfIP+7hAq7553ATIKDQEPDFrFaWceB22Y6BJG1b9vs
klyH+GBlsifuiUpfDWvO/R/cdzfrxJTDjZ20VDbMN2ecuabJxKYmvT6URG1UeyBM2nZQ+XzQUyA/
BQHkcJUs7/Z7txiqDjwYlK2L50ya+5ei6HQ4vZPjkEBe+u2/ehD8W+3FrV1WxVPXxQGpaQsT0jDk
ZbeZTDXyRHSTIUlgV6Ifq2WoIlq3c5+S4RcDyXKVxiwm+Hh4aGTHNwnlWjQ+yl/htCuLiM+Y8UCh
FcussDcIeCWY/A4zGLZUWFgZ41kHAeOSJ4Kj6bGV3urtyLCchJdwk3MpAfZOEPjaHw//tSpSezC2
h8nf07k9I9DLggerF9q1JQy6JurO28ovKPHLmk2OGfK02tJWfPnBFXQtuOGW00UX6Ixrk0XnE4ni
5u2zn4nbngpLFG6upu+PbNRGVyJnVjpGV7AKvQAV/Sxu78qkFJvUucalikFEtR98506mR5NUQdIh
bnykXY5G4prVN3Lk4Gy2TJ7RGrQ9NCn3kUHamUfzKve/9CkVVWDfko2fF6fFGsdDc/mt0Ss1gMge
tw9zfFuy6XCNz5nqwSRXdefIc1Ta2yzIZjY4Zw7GCWvzh3eYLAVS8bUm1S7XdS5Ps2hg9Tx8Qa8b
drbEFSdVG51yo0GqvD9sB924xpKAYcEoU62t3qguFW1654DYkv2muuya005xrhKTMc7DdZOZbPVe
x8VR0S+sz5NlMLSluPM6bzawqdtzKzDjUt5M4/izlrX2y9zymd/hCEW7Z1KqW8HokSm0JxDUxf1S
+wacOZcNJJ0nHY7oVqciEww4cFzC9zJOppaswRgPWgEitSAwbXDlpoaY1SDYkhA6sAL/xNO7gMx3
xsPXKI9ghcnlZggY7A3gyGxsJRh9uyMnLOjuWUKXNlXKNKi5wGQ99KuBioU/CkiSS5hCf1lTGV1Q
OPEbiy4juv9CllcrykknlWy/Xd1WU2vF/xSxdtHG+9EnDqDdhd8q7HDh1zvLD0Fto8OHp4OlDsuC
nrH5WTMaUP51ioWLPkN+DFIsbdExjVpdnoneK4bbBgnuWJi9ChMN3W72vj8TBLecPmmMeOud+iK2
bdc8WTitq63w9JxWypcDB/pcxXN0oJC3WTNnv88h0n7fvHrJkyID7ni29Na01y8iHMrWkMj/F7Tc
HDhv/9ZKtgp17UsMrfSHFChZ6aqjighVEkSi5bgegkPAIxOsSLg3TulGngadgzidi/V3QwJGInVX
AeeytK9D3iIwPIJi+19IRD/J0g+UKd+KPEmj19UatVuD+D51WFT5/ZyLi3ut5TFPd202ZEma/7fA
YKG1OKbMPE8SVI12ogANX/eOE9pEAC3LzI+LmN6a9nUSAffAGlI3LIi4xk7oWG0IjN36qRKxu7qH
ycuETqf8rlafDUTCvHz5uVZDRNZQ7sDnoAKfhuGT1X4xd4LPe5v8QdwTgm+t0pblZj6AIwWSf+Ib
Kh1TfJC2ecJv6Db2+XplcX0qtqBPwY7hYMPfPONs4kDTRwM3yOmFJe2bjPnPT5JqxNYA0KEbXkWK
m5iHlzL6BIlNNxLCkl1FIl9zIMv4pXOBfct/SUbi7grZZyialUYxTxFmT6sfiusH6Z6W5Lmo1fpD
AHipHZy44x5zDzGR1m3mlXnTpM3c1Mi29Pz//JtqfRzuGw5TcEPDubbUouVlOtssmEExbArK9LC2
GwhtjC1pYWzSdN94sBxlIWOWlJ+MVpGSMQfgNYkkJu1tvEnt1st/P6fcpSW27Z9Cn9i43xW/HZp/
ZtCXEls2q5g42eWSA+kbf3cW0rQcebQXJRYak5xta8kDFnqw5b74VpyNd0YJvz1XYvE2vRDHalag
V1H5CZAeoe1QbGurAI2wOSs/HTWkzzeRZLj0D4Zkq1VzygPHgkWAujvxxfCJC1joPWkGdtwSp7qx
LbAyuVziT/F/ejb0RAVVuJtLAWWhM3yjhpZRgMY0UDTDWe3KMmY3OKq6N+Z8UfBctuZstoXOJsrl
n8s4Qtr/1kSBVBKRu3ys2iCfeYnfMKBxMh1vDvKL4PhRtkohb3JZ2QEIQqQXv1/olsqdUHwXxfXG
1zfR0shQ72kdIwmidqWRxIl75eSSV6vF+YO0i/xCKaVkCTY6N2F5RZ5x2DHu41AaQ4Ha3ROGy/1t
+qzAXTDGZf3nQqRoO0blts9NVZw94adzEV3y0UJNoWZ6fKuUegHPiX/R1PZFOPaS1npC3DhR8XLX
Q9sgcFL+TYwSwc8vDUP+dnYeWEfjERsoxRaYVwxSJYxDvmhMEpALsGJsu4/R5CovunDw6x6tEAoO
FT1Pe2QOeWCJvekcDEmezpCnMbGFGb/C94ZudbRAOARg7Rsi7BYghs7MWNwq4r1PZ0JRj1FSnlG0
8qRacN1eOFOAstuaIaf9D/5O9gXlJ45uYQKpugpjLIjvxDLA/khRBiWRWrwGck0Wl4JEVLLSqkdD
jG98ByxwOvirh31kAe2EdP5pCNd22AMLfGOOGdc32dGpRBhPJE367QCz4Vi6Aqn2V2Sol/dTszG7
w6qAMSUMhd5eHB4L8wzaSLk3wvWzstiCh6lx4X0uOny7z/LQhg1YIWuARMJUen8U6UUuGIOz6Ljh
UyDoUKA5Hd/UC8EJM+Sr+76J8QkMDwkL05Uz6zm43K8Is7kbDskfOuTIcRLSXPR90BqO50pCJ/k5
h+LpzSnyQBpY+KDHzXdtkvfE3KJsfc6GN7WdV8Y1SNZrcf6ed9UJv7Z0bAUxnyjyk/nDaWiwDegK
b/rNb3jI+jNCekpnwiTIL5ad0C8fNctR3DLCtWkjDrg7nUNw+gVXy/MBOX11acTKyUJAMfZWqPeg
iDJCFcsxXz0D6Qt9wxVzu8kFJmVXnekLg6Lrk2yQDtetTJw0tTYyinRGS4Znw+i5dGbeiZ2M5HEi
pokDPFF8Vq9U56OW95t9BqZVhbE23Ubq4i7nOWnJh4tL0CEznLvtQGurj38Wafip5IjR5cUT4eMQ
CUlnVW/4fh+crEipTY8CqmIGXIqhla9WZOpGAUBqUmvKd86b8u7JoNtqxnAv2OtK6h3kf7rCW/un
jAopV6Vk/MdBpedGt2KTQXiyY3nJNcSZv5knHuC4rHBlMfrkAZS2Iuus7Uls6Zq8EYwCROkwzQWP
m9GK/BHUNlEIUiHdbMwlndNnWpU0uaHz8tpGoDzYhOBucx8P9tS/uz7lH8Wat+Jegvqj4AhVTnp/
JjHS/aiZOxI2v1wI0JKZ7owMMWJcRhnapGzqVmjndrD5smM9Xk1IAGawmvPQuad8wOf/f/HWZ4Nk
67znveEENEjR9pFFC29PLSv+YR7sAgRuSOpoIjX221XWe84q39dkBRo7x9HQv288lTei1ZiJrIHV
nBSxWW6p4JlEq0d4zuhWTzniKA1WQslzV023bhgSghJ2GW4nTZekz+FQsVmVDDKcevSqKvzGHxLo
Es6P/FkuQrFbDy5QhPI48O1wKqVkqebrT7tknFaMcENJmRv+dcSF7sniuLL4C08BptpdRvKe2/FX
yQzURdG18LDruIfZoFb1D2ZGuiHe5GlPnV63cy27aqFNwMqAY5yOEjhhHeOCsr+rHsN5G2gdle8b
OJgG7Uc4HkRiCAxQjji9PcsDScqCo0q2FyjZiMDV7H66E7fWMnvJXQfBhhYy98s38iNPVKsZM9lL
P/wapwYP5m8XK9lqIdO2D0US1xvw6xpY1LVoJMSSAhkMV3hFeqJFRZJkIwr7aMkcJjbOl7WoWSMg
52YGqrGYSdJrN7r5rjV0XxRHnIUEozncSZlKvewj3Cj5J+uya7XxrBXgcIUyS9Hzih5FxqlNFILf
2c49wafo1zuycpj17EAKxUMgEuDJBYHSC/UJyiISxQHE+fht7OKukqtPyji1NU3DjgemWd2oxmA+
xZNEOwKnAY14WzDGL2FyMiKVoR9WFvUvQ49zXrDHr1ZxWj62R0EiDZOBm+59t8sIlPan1WaZSolF
WyHSOGBwYGxmpi8TDTMXfMZrvmF2ObnP08oS7nXdtCLajhT9joOwylaG+k085jXC5BWrcQvZlish
I2HnMx4zHVho8CSWWFniOcnM3xWIxrOjHK4OlLGGJPfdoDeL+ctZGNFdv2GHAdu5mqjxez5xsElM
OKNrG3wfUxNR3OaLNPnU7zDCP0y4eflOJ3o3zOeVYE/TjtMt/1EGyEigX9pLN4GKcuK94hPfNfdJ
IO6VsUEPk66aC9bJHliaJBPngMbZoMk5B7Cy/rO+FQIARFffuGW6I8WzSKGpC68oPzmDc1sovdgl
QmHrl9aP8L5yWVAZkHLMo53vAi7sWMNSueZ609E75KY6l7z5rHt17jNSchn1LlnhX3GiTcjMDj5h
nhH5cepC/KufUlh9B6OvmEErz9kJopTwAd//UIigeRZlqLwwo8O8l9OdkgxuqayAg4Y9KHEeemZ8
256qPzuPa+ltCHWvN621lp7Y+NV1PeI6JB/qvQmZIt1ENaoSllGq8DjpTkznQOQFWjBG9mA/LfXi
CULk/p8CenzPZKnTpXTRcQDV9yKFlqM3OeJaLCF7hgiUbPr89RQc0dSrCk4gPSjdPlZYlkGvcApJ
KuM/6Scu5ywrMbIxn0V0FxwVyCtjRDiEzGKq7R9jbL0BU/LkgiegYGDFZzeeBOHO3nvORdVSULJ4
4kKA9bsZ0p28R8ojWoovMpKfs+91uQB5tP3khtMLdmk4KQA7cDOanPSFm17c7UaKxs1hLtc+Z/2U
jFN5AoM6e5mdM/Iwi3Mr0PNIoi1fjkTHYAHQZ1GN4GHZj8tnsAWh1TkYP1mFjSP58YDDDwNPqxac
KNUQ1ZE4X5ioXGvkIJYJaTrrkMW54QMELwwq84gXg4oRj81zIWmg/Be5dfQVqNAuom8X3XqMS6C+
rYXzaDnOvfN8QB6uYwGOpVcayUpwrFHLMNAXP5eB/hMQlnIydc1stGNVwKkwhc6zN4N/LcnijTiY
rj4g1pmoMK0wP55RyHHCCjveOchWUqpbfr4//NnVovAySntuAOFLZGO8cyOoCgVzmADFG+6nvWEy
k0R8F5PG+yy7wAXEuiLr5prMFMx8yWblz/WBLMg910Pe4fSYnGCo0wyM3twm7STdvyQ43fDbcC6q
r0fMnjVFKiOs1d/Gr9OzSycYTCHx0PARrx7/Ulv2ZkZ8KXCuPGsqMw8D9kmcOVOOq4D6psILbPiU
qLmhdZcT49DygaKh4GythS3YGDReQpDAcINYQ18tKX9r0sgy6+ljUvtHX+IsuGS5IwV+Aqwh+Dys
n+pVbyFVrhqATUtdVfGiMpKBBH6Hz/eAWwuFRRyuH/t14MGSXVUl8I1GbBi9tv6I35ao3EI0yS39
SwGtttDDWL840nm6c8QfUhOABNp5Qll6xdaFzzOXXgXacBP+BD/4ePJf5OVX7wwkkrUCt8FXEJD1
7KCFaDvcl9fAC+zOoNdJF174mpoOCLQlkKhLr0nJxBeomqAlpO/KxMjzH3J9M8BwMgAW8nrSQFv8
LmagGbkXna7Wmg+S5uZMNxmPpk0c0UvWjcYgjSSwXFTm4UCeROsQ96C23ikhoyxeCIsoMyj7vclF
PLcOCMddOlnZNlADHGL/vKtlNDa89ohO0l4r69pw0j+eeLAIC4KYYIUgTuC1G8EDuatY4Yq6XZYb
9Ecx93hdTD7cdlwMFj+Ag8h9uLe8kHeyDO4hh0J7Nu0Ybwr2kCD0OuVxh9pegLnEEF2Xou2GzTTQ
9Pb0gdxvCrczy5Sou4djHftAtfseh30CvTQaww/hFnxq1ZvDH2KSMcm1/BYHV1Z2sJmhCq3hXskH
zetAnVBsZNiafCvBDrrJ2SKS9OU8IS7xMT9TcJeXETaIIXnvxsdkO4lVwDBHNgYOOSVil32C8k6g
aArS7p18ZD9XAB9OTK2js1Fh5uwFfplD+ZmFraKl/srtHPbBXAjG714jJ/XKkk47R0jxX8M5KE4y
nDENAB1/5GVFj8HA8yxDGohLdgSMTSHLqd5IFGB/xC2Mh60mowdfCjo+BKvBDS+wC1ejPWp+aDR0
mRfMxSkP/aeq3Hccm7CEdUiZubc5xyfMF0z6OGNg9+g+MgSfLQiX9lj40R6DmyH+T1yZUP/myQ/4
rYP4z1k2sF7auF+63GJO+No8XKbB3xd49uOQE5q7TLNZs0G/6ulMC8lvFEZ3TMEl7aD4b/HkubQf
OY1ImDx8e+tOpXwBkJ/e38V3cA74jaM25isbFkSuKQt3lR774IGiFFJwMyscZFZ3GrjfBUtr4sFf
0l1A1T8NJ/YWwK3kPNt/ck/V/FWlmXOJhO04fIBvo6osJ3JWUpJ11ghHhHUCJ5nb8mMJSBeMNjBr
HoiOrqZW9Ox6m6tO8fMDh+gM9aiEtd1N+kTCxA0j5QZdLrMvL9m6t5AUzotmAJqzBpqtS7Pek8GH
nOFSwifvntuhQrXNTspPvd5YoGEmmy2XBD1ygsXWhoHondf2hYRP1raIv63dypDwOpRZ8NfdSNYN
tS5eXMC/HrivTNAjQ02H6V3iA+XN5WsSumse8gN6cfd1q/mA3Z+AXaBdhYl7x14B61kKirojTqzg
LChNk7eDccXTjpE88y0Ipkp0CNGR9mMQw+Tw0kgbkjDKJNdWNjVT8qBzzLWcJpDIzxu26G9r0z0z
Y3ivSU5eb0tpvTElJ4XpT3WFKsqLJBmS7VdTYXi7o8FKPrdpoQLh1MrVvlb+FHGO5YvWwAYRKrhh
PWS9s0qWqHFQkhXt/zIw1UjUDAAt1UZqhs47QUcpHoRoDHv5GJcQ/hrQsd7wRV97D59Lk0kAYYm/
7aQceAjNWTkM579nww1Ea8OCLQiOUzFQIe4uHq/Ochdsna9JYy109o5wCB/5WTX+BQpn91Q/WB4E
43qbfOexGTn2BzUsWBDMLIeB1TbEWzVkQbAxIfjoCecsgniFyGmJJlHU33MOF9kbTG9Oz1/+kO45
2ySKsHMaTr22VKWHmh0gVBHBJPe+P3HLvRPQQuG/DV2hVz7g6VP+Otd69fOVzIoV6xoI292ZOVAV
Qll1w9cnj72XeiBGasudrTBpBKiAMFF9Svhg9HSVs5hrHQT28W7Zohr8rQzF0e7KeLcKSfl6bPid
RTdpPWZgu173b8hH+w4gTPGpPoIk7KNl6mGrPNbq9MD2K0yN0SAF3OUePhA9ZIzvEmSYFSgAu/cM
IvGcJZHrJsMK2myr0fvYQGTZ0U/5x1kQZ53DRmHRgh6TnxbQdOvq4bIHmIir3hc5K9EZLR1sKBe8
B5n5MDPBwGEFmU2omZIKZK+W8RKGEr4QL9Z3gSIwAT6EZcUl4Q7lVjnEAUOV5FIcEhYiMyvH5x7+
VggAXqe26vijvC/GBY9unHfJiLeuhqC1stv4nOfy17bBATafF7ocPkygvIrW1d+BUsHh80FGLVK2
ULnmb/8dwWx+2oj/jdmZfSdKFeuxr4IeTHvzVSDefORcNraJ8BgfYbv123APSveqaPP3pYiOU7d3
NTFc/JBsY0fRlshvF357Ani41zsjFGOI5UYxn5RvyHZ60RU+OhFuSAzxkjPYNJwVBqeMCh7QmIAR
khD2/+QZW2QciLxcz/DWvP7Fmz4XWz+w3qqdqk8IQr6LkR16uLDmWByFCPVf3uUW3PccNnW4hkdB
kd9bRmAVNPVdyr3v3GOnA5V0F0+bh221OLhftD412MpR9RVrnea5Shhf+6vgqfd5Lb3k7/dyYRDw
JM5lHQUbVJ2VMRbk/trzyJRJgcVXxLS1OSiraLmt/f7sspDDwxA18u9DWIy53eQwaHHb8grVyXRo
w3t48ssCVZSk8FNocuVHwQwII1wZFhJlPg7gMwKUvauGAV1/aw7gXK1KAu9HTTeLpAImsrDswopn
AFM00oGT4cZbAKoocNvKpWdzkUR2bi074ShmYJ++oeeTsHApIbMlrTPI8q6cL+F33oXazMwWHXUD
37LyZT193MygbqP/MbT4XuLHl26+sYGPiSgIegKTokZBEE7OondZqOyQtAvLq/8DV++udwzqfl7k
yeruTXvTbZwuLX7hPKEui7WKYCoB9GycBqvEofwkZFClrScqNJLQmnKHkMEymQIycLbwIp2Hcr/Q
BKyapYrOch+tuMFkynIGi3L4k/7UIXZYQtosJpMUDstr1vJtWyV+7dRpREqeLNdX4TAxOt7ofdhM
ebAMMmM+AAOZVHr957wZAvfzBAFcI3vTeEmu8AKt31EK2JuRfCApyRs28VNIzyH+2+2JFjC+I7g7
hGh3FG+ffOKDDMBw+eF9lreYUHCJK1id9LLsa7BgqRre19Qnepi+Ci5okkxhCNtaNGIQfdhj7mUu
V5XXiAj6cIAZyDdrBzJ/ZLutPkAP6HFW7PomLNCRBFGI1gZVw6pnfJEJe+S7j8iOpwJuTtb/PQJG
bbSF8Nw3RMaYJOauIkBUhY5bOfjcHnsb4UBp8ZyW7WZHzWwtxN5EdK6iV4FkWjP34x17GINyg8na
bFsg8+UDv7Yq4h6ErOMBQJNGx5/jX7WInZLAwR1skVQtFswXY8o2eHzQinXIIr1sFzQXWsKano0q
VpV/MAnZiqUUjIZHGbetgfUOWl7eHdBJrrabmCfXe7VliRLbB2xh2FhaGoZeQDb5ax4fu8fRv5Yl
EFNPN+VyjMRlqrXqArMdyBHurRlZJgJ3v229gbMa+7Q3M0858KfdEq5qcxBbVTfB/1ulOsoPk64Z
d7zmNZDRzM8PG42eGobecehI2Xb99WtD1dDNZNmHBJwC/QoWicCcNXJZDZwtMdIsX8nFlM99i12R
E6rQBnV8tDfxo868OrsShsEF7lZ+ApCloha6uk4vbYnHdB68yhNNn7ckbEZFoBTkS6wYvYRPbB13
gvreNSpr/j9YUavWZCWHl2+k0d/trzuA9ywj5rvnmdn7NGvXgF19EckC5ewN+a2GNZL2AW7q5gtI
o62mVkT2LEZr2ZEqnksWLWubs7lZXyDZ0/rYikFVrvmWv38eb8mcGzg/rY497Wh7/bfHqopdHPmC
uSiKSiVgfCczKNAOdYElprKV2XdIhgtw4TVCNUOHoK3Ms3QIAnnuDdh08Mwm+m/takJCtn/Cbb3o
MpibporrSDHHgGimJvEQZX5iyDl0lo5y3lGcMKwxvBjN5PrLVsZIFKqKu5a8q09QgdoBg53HesnH
7lD2xXH9OZVy4Ba3v5WLjemswVLDsSWqY2ElPpOveTOLymQZJtSdTV1pv857GCzSS1qmBB+psNY5
12l5pXJqAQJVh6yZl/FREuZZl+mAo261KcxfmwMo8TOzmGPyCh4G4LFHwyun8zNNnCKYh/f8JFoT
YIlEDgPW/TydQr6uaWedusXN8oVRuYl1NFxs6InjIgY3nzxcj6DsHnLtKbY6PydzFRBoV5G0wB5W
ETfr6CWHjc7nOy3EAlDeeEEoA7FATe1R+q6i2mR3Zc57Hi66pq22g0+XEtyhQBXLuLeigpx67TE0
b18i2Bm0j2heMleLF1RFi1v5bX2A+tcobORBBJyga04ag3PtoCj02gLU2tPEHqgLGaGA/skF1bfi
sQoXtWKkPEcP2v6idP3OjePhwNrg8JsCg0gW6ajo3l6t0Yk84G29ht+TFDw4Z4IsBtD5YIDorxY7
J2c6KTMqc8Uo5BX7qR0S4cmjAMffIGSKkpDIQorTNhShhg7fOUKjbin/ok8lQTbS+d2VzAJq1nmM
sSBNFysebtwbAbAcx3xFSz7Zm4sMY7PRyoLJ+IstNY3/pfDnN1VZ0HwWEv/i/5n1hlpP+raiEoOr
i5qhJdXmhVQhPyoPpg7mvIZBL/0k1lONs7F29g7kH5+wm0hBgmagqbEMVaGrn5ZstMadeUJI1U6g
M8ro2BdE0hH4jYUFTFsVlCyamCEIN2EjMiv0/nHvmZfKPwQG30NieHgEE0EcxvAqkVSCYaA6lJ+g
NvWr6Wl/hUk7eJKk1x/jwEcrlk/+34L3DZ1mpv5dF+SV0WJ4aagb7nXIGiqf+TbSjg3DwSYmLqr0
LtQp6kDSXBIOot8Our2WE6x94eqcwFOtyWbonNs2zO/7Khv6tRU5iRb0n192sEpXFuspno/7lEcy
9yfS257BeK8HGUA2ld+7jldOfmPNvvoDJbfZrnwPlxGuX1dVmQNxew/B/xLbHIogdaQ9KzhzHPZw
1JEjmUsw2uY+XwXM0s8QQfQ5sGsX4wp4a456bv/QlNWQmQurjOt8ykZsEkUVwwaYqGbSWUBSVod1
Vt6jib6NDI8UE5yXY/fIwONQh5LIwpQABNS/o2m7qHeSFysh61FjoEFy9RQpbt51IKX/NQ0VC+11
EiVN7WpRz31KeWAJCibPYPobOrfrRpz1PHhwOl7MeqmlhJOUUEjSqVJjnuFkvahUNkndZJ8tcMYr
/opncPeQ2L9bFydXPRutSxkuHlD/gE9rvwTUOK7QDmnVQ87cUVPTXhcNn52YEncVjWU7LFRPIbDD
9PhbR+t2Tkjgw7Oh3yZ00c/UESctmS4omyZQOyluJDpo93m0KTnm/6W9FqT37+DLOj73ps0lgrrG
bSgEeajN20VBokM7PlHcbIY2tPAae5Hb9GaaCfLsGfpTD21hBF9Qc1RNNEbSc/eMj9x9xlONIRRa
dKjnyh2Bf87nZCNIRfuHu2ekOKlnaDtzJxj9QxfLVpp1AhHz4PI1kdmij1j7AWg7GwUQexDI5DDL
x01D0zW5tdi/Bvs/NE0CQPlctvRbMcfzGhCQR4Nfc3OoS/uyynDnWEfOGc+FfuCZ6yZV4OkmrNYV
kSkBraZIY1th+jHbfGSyIP1R6vGNXDbhOIVwtUFULIbEdQe/WaMlS70EBqlVQT5R9cqtFVhlS+9y
xnINaRiD2Dya16Tpp3SOeBdta0lOuGSYz69CCvwK/xRNusoIse4yCevLpCj/V/xQsRT/Nu+FjVF5
K1KATJHqQwQp1btU+d9nz3hxmA0dzUFCnbCiY6+qb/7FXaZp0rc168NqzSONNSNKrXHXqU0uJ9er
bqMvb4/NhCDLlV0rfHiGg9ENi8xWvuRVwAHYoj1x+HYRvm3KsIqw/sjSQgzlkiHfgEmj5OU72abc
O4tXAELMP6W4WDYMX+9T9lH6Xroug6slh3Iw8lqIsS1Tgl7ZaskyjRCadKpYSN4yyqgmrXYi7mNJ
edqpS4ByGNFLBzMzKjaM8KhBf1JJUWDUUId1Z0gSZPD6YpWS9R/AxdYMNMPG7Sii9qA2hrEnZVGq
d4qH+Nhq/HCwSMukNi3b8MvvEtxBJC5KvF4qQjCl7aGPhuxl8ZHBrtSSPXuMocIB7Udn6sbKOvu8
lv+QFhs4CAXNlzoFYd2ggn1RWVcwNwLf2P4tlrG0kvh6b7ClF1kNEv6cytUiKY3gX2jnxk6nlkN9
aA/Pfe+VqVHicQemED7bQUAhmzexEp6zxDM+ZCKSZZ07zDQ6XLLOF1qoJHc72RHl0ODeLwV6CxvY
SxI+Ny/t9iHFqk2Po84p6LJHT0WKrymTnpuvaYrNjpfXEvdv6jUL+62vmiqP0hhHwAAcR2yasGTN
rODno2Hl1bMztmhNZXIjP9hYCHO8r6twITS/tl26ajCYhVpS6+9J16XpTsJe+jxYHXbA6pHhCtM2
wy0t7EfRhbHYDHnHyNhnU9uji8VLxZHGKElcEDUTdaTZegS/Qma1X+6MI1maRZlqUmiOEq8zWpQh
95Ybl8kEKzv5cAMaSf5eXm4hzRRY9MD8GYU86sLvYlJ3x+CAgrPnmXhVX8WPJUgX7wZjqOcJK8We
81o0b4vIBBjArQsswUAfGd+xh5HgJZErw8O7/pD2EkWbcw3l5SOEfCQNaUoU1NLMOkStjhhDCYnD
Cs6uAb/PK3CQBS2vw2VXxsSLrgzRBJLI0ayPEXary/SOZ/YHJ1S2vP7nKTCgde9+eBTgkbyxf280
7mgIdmyLhlGhfqWX4zJF4oc55WTcLkpFuSR70ed+vnclIBQOppSXNzLq+OLOFJ3Ocx1o9B4+T53H
v0DHpt7niI5JBOqp5I725Ex1D3VkiCOPTJPUHio1z8jwn1ls4SYl9dmDT9tl6zsaZn9BvMeNWHog
pDj15zyvvp5rCAFR/2Q62NnZFn0vlRbe5PJO+PLTN6LS1kG3JZSaGj+jsJc1UEZJvVpXsqw4HqXG
+ca42dPpOdM8/ldasuKYKWJg/J9V9HEM7hClBf7tnd0bXDcG7a85LbCUhjbkRRVp1jijO0fRLQgi
1EFltr1WkTOvTHA0nbWeZArwsYXgxtJuQkK77ic1b5daST2ajotzDr0egjVvbVrDUMcyzwl1ILfB
y9NgAEv+9grgnk3uKH+Vb3DvgWvabzS+EbqTlSKSpGE194yotb+HkIm2p34QVWwvsqTIqMqD+fNm
EuLkE9gJg7qXMK2WA3wUC55i9sXVFqm13MeHtxZ7W1ZncjDQGxx8K7nub40eQ2kPjmHWkvrOG4BC
J/XjFv6DPY14s7Lm57pLETCfkm8lLWtT5iymXZUOIuCpIkR1Uh+kaM0SlxtnQNMyVBg9FANrOkqX
BeBVaGjX5d36nLNWEiSNXJHDCk+1H9i5GxKm9ZVk9h0VXwaOwtQpiHXzFs7P5eUuEegncnRk91Ka
S4Z/++WxAso2Do4Aa7dOFRMaTh62fQaPkIK5lOszyHD6wUHGE/d8T2OTcQem0HUKIZLQPfd/IV21
hGxe78BOHZKsv3e/96wseP6WfaOTsNgEpDBS8nhUm6cwNC+Ygod6XQvwe9l5c7bbq//7qjQ86Rgd
YaoJCao+C+nEyhJPN2NMVNmEQKINWz9DBO79VhJPCwjhAwReMIMrXd6zQt93tg+tiwe+OzYE5CF/
fz6Y9W0n5nVDIqwIC8KPzB6Ee9y7oG2Gfox+vlVKmPeLRCeYpj9VhtnT1Ln9OdZaQ9GkZiM4qH1E
9IddUeMQDJe0iR52kMHv0FQEhWb3V9fNuJBzmX377IAxYYWGmm0jaVK1mxgct0KtGkXZfaLiaQ5Z
2NV7HRNwlh9ZchA1xMc8XaIM3VqrsqzVSWB42fdcmWtIzXD09fd0pv/BwIZQy8tqjw99IeUFeVlG
TKhMlvN3EqdJ9se2BdyeMgBReOTmT13vL9TpfE54E2ov34eUHJcfeUbQ6Nj4rCnfioLkO2Jb2YOX
nNQa6dYTECecKe+0EmtxncEj1MjGK2KMgRVi/rlO4582JsFa7Gq4ot3qglpHC3AIvNmsYh2Afntv
55IfHUup8dTSj98zHdHM1hdG2xs/Hc6I9iqWg/koVaA40EpLMdmrFIGZc6UFRQWcytoiHTq4AMU5
bnprrKynzozEL9Mr/oOvDzMi1WvMSWv9wgewXcdUD7241VuVxwzHJ+6hyJCFXBw0VFsCjiiQoQEV
ozUsjtyITaO4Ufkk956S3mS7moM6LwAumy4VPc0QDVWWgisaRIaSXB56H1CSl6a4+wjq6m/9Hu0C
dBN6QGBEW5dMk8mGGuukVTBLbSQ61IBhCOdyN5jFgloFbIzkC3del1PTlyCt0Z3vDuuvTVnS3IoG
GpNDTBooxd8pjnH0w/XKlAfi3Harb3P+u9RUpLOFYlxKBrD7lgaS5Zvrqfv/yBSc5kabCmQ9+mFe
teu69uQQnRVshyHCyBYp5H1NCVZGPfj5KT2O8j83OfWxA/ftlqYgtmpHBRbmVCu9VqrIZ5t9GGWp
P3/5viIDtv9+oSV/tJMlyDftGiLSWnG2G9DgOzRbjMwSEdPmhMdseHh0IVA2+SNNv0iQUHXPAlqG
HpqB2mOGw8uMjgOSAqc0iXA9HUQXfgVZVb1ib69FlVGulbMiBqQcz+SH/wFh//zaoq36GCdQQwtR
jVsXwcF8TjaI3sYe/Yw8D8fJOA9KFQu2xYRbhtQ52h86IbAHjO6+8rdExpOiJk9IXe4OiDbTW+qJ
c4kzVpdxQJutHDyR9nLpsAHs93Fu54wjGoUCvegGyJfw+3cRJIn7Q9na7D5I4nOtDw8T81dKEo1H
j/VMYI/ZVDDJSTTtJjq4b6LQs92s1LXpNWXpASA3OYbBPSEqvt4t+U7MwFa3a5XV5z25JXT65F2i
yOOpvBCbv0uVqvrIOKFIMFlzBNtLzK2b94rC7dfp9M2ug0RF6JOjj1t80eI7WpzR8fUcrSxeGHtu
XzpeGCQnmNk9Pz7U6xunT+jzd7R56DvyEZG6GLOzRP5XIHlU8g3PEP3sJeYiXv/aZtO1iUQA0OWa
1cwGq5YmYeSyajNzX42HwwOEf2bEwzmQur557fGIlbVgcDI/Gl6c2uzQjCwBToFl42aPfBIYHImH
jSfYUyoczLWr+g8axZ3cVzlx/eDuKl1O3vriuWJms1bSU7PtPNG0oN1oRQzv8YOcBNEy69XDaHCL
RYjBzsh3y6Se9gHFCPdmATBn1YpEtMmVNbMz/FCnSoxmhfW9H+wolpLr3nqzgDgcc6BV3qyY/xlX
vumfC4f+SxNdEox0Q0CHLc9tYVMJw4krWvMdFyp4fttt8QdciwQXpSO4H2/Mx3c5P6g1wgyydDCi
Lc+ZCOxjQYR4A+0yHXfC1csPx5EIXefKKD46IQLG/2gaOxGXn18h9j7wMlCABMPq4ElzvHRCV9Di
LzFXUFOjx//MCfejOa/slFUN07mnjSihS8WFCZFPn23PQn10hVmxRUyKX3SijE4vzMQG/7NVwzAo
Q8w9C+rlqUkW0TW+Pkn5BAxsLNIJtYIkXLgYLE1yUoJTgpTgtqrFDvO54lpzKlX/iy3WracfdYgB
fuhHjY/FrCW685SS1YMTnRcbaVigbqp4ibtfC8trApOpOxIpMb4xiEN3A89bUXwIhCd/hkikKgIe
J3m9hJEIRQ1+EKJe5R436KPW32LQs/Pmc7ncpbfVwdhZPS/6qMprBeK6+dD1IRUdRWOZiEvERa/8
LOdh57KRo2tKLcuDg+dpf136dnMuq1WOlf9PsKxn6xEr8j6tHH8CcGMz1OZFjf16xU+UOHUZTAKy
T0MWjQvHOdsa1GbNi8UMtxIn8Iio8FxkW86nvzAMKMYJc0QnaU6vA+zl9iIVyt+NyfXQoih2Hs9F
EM70UefCug20H8waTM6TQ4OHdXXmQJZrAhA+tBGqpvkSJFJmFWyfEuTqbA5Vb3UCM+O102mLCw+i
eSFzdevgk2hG/3+/Mt2DslII3ssEtQaWDO12WMw2o7Iu4VChGRJXvY97Rnix+i0Bcq5YjBo6HalC
lelQKPExHkcn75yK23J2NI1CcfmSo+dCnY/Pt0DBNtxr4a3lOXUE8TVkd7CHen/ipwgaU88yqTCy
gLSRwRnxRoRy6Xcv3oGX+XXiGbaEO4aMcycwj0vYOdTDSDw3BwSppXU/KOiOOQqTua/R33vFIVb4
wjnpKvRmzZ4KwaLT6+GTKD3m2V5sBLMo/l8QwSx28j4dicklG8Dvvm4VjN9pM7g7MfgVuXUYSlSP
Vi+5cR4wiVjGKanosa3pJu7/beWFKFCiVqo3/jNPVvNR/Z7y/PdO/wCAym5RK/PfmXVEuY8AfGQn
+iX/Vhr207b5OuK34RlJGXm+rhvVf+wjzmBZO+aPk7jTxNYRGk9g4eyjK9THR+Gqz4JYJkjtcFwj
zBc6LDwu6qROf/+7j70tybHh54gQBiJ5Dsfnpyvul2JUgJTyNUDlsptI2jCQPWOcbIsn3klYBrCc
MDABhVs=
`protect end_protected
