`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
hF7ZiJ3r1waHilLRTNFq3T2WhAu5WNAm3ByOne8Ilp4L778VMS60B87k1QX2GJvRI+n6NECP6ilA
MBPaN8cWD/wyv3cNEsIvuuIzb4gDG4u2ES12yA6I1vl5wKm5AP5mpF9OcduMFyFUgPk9o+OeFOe5
6Fvj5QLRTUa7eljhid9VEuGmViVMYB3DH6wEh3YLHLGP/m/6s8IKZxVyZRyGjVweYQxzS0wDRK5u
bLxEUMf+/wO18RZfzV3XysLCn6i1I9+aSNmJpVkRy/vD4wSO3xrX5OW1S2YDGHneC613O//dEKYH
eNeA3c9kUeDnAcX9Mz4ffoa+QqWWXdhWQej2rw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="jKYWQcnnKAUYdxoFCpF1vsqVazTfiXOyxVN+fp0P0X4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3264)
`protect data_block
Vvyo4nByjH8oRMIuocnijuqod1xhKJDvk28YAU8XWqkDxUNQQb3yXvD698RuTO/tvnAseZ4s4M5R
5yl4Jk4eTviHFj8KwjKWw5jzgK4aiDZ6temnYHTPEYoWIvK+usEPEdjGuZpODdQSMNTmYqrZTdE2
4sUsM0XBVUnczZzFGzywvW6h+gVpflYKUEs1Q9be6g80VbqQGXcP357LU3YuGWUZO4nXZ6YpXOQ2
u2tSPQ/y9lfsFc7AvW4kzFHZbtgV1mArtApyPzpGFK3FANfPCyXafKnXKYaHvN7WveO3GQcAo99b
1L7Js9OdZ8JhaWCezAw3zFFpJaDVYHRtPg2OnLlBoB9+ZBu+QUde3fp/7PjAKo4Yn7tNqqNtBAkN
bNSkmp55z1b1yvYvuZwDffsqLd1mTyDAhK+0csxhOuHN5EUTT2DdrC5EgFO2myR7JDxEcz3CpcFf
ecpQoW6BZjwYul8SUmm3bEKI5TIbKzErDLZWZvq6nfD89efaFFnowoMQINO3ff4jvFAT+YClCyyg
9ItvyBh+Q59ArlXKKJCVg9u8Ud4HmT43UvpIec+WZcwebHVqg2czGEA0br7j/Yuzja+j3s3yIqV8
PQkwwBT2gW7+dgE5seJMjZOOwlOttZJDa84GKi7Yb90qaHBGJmDYRqDk/zYSmKOsfC1cwUL3r9I8
VtSTmpsLtO6lqv7qzZk6m0tbGKG/UwSoaYykOhy5h2jS46zzUB4d5+gO0B7IUMGoVjTx0NsFEi5C
YBT6wMo4ReUNvCuuzpziiiTNUbl0+MCoHVq4wIphpCTdusM89+/Nn0SSsuTbEqFPeB0t/OhzniWo
Ebwv80PEycaifLwYNELAAy59mzhPTyiv9giBGdCyiFekO8PNVpHCla57rx6vKr2UpvOW1QQsJ2j4
l7jOGd7YCwME6AhlFsgZPq3ATb17JkCGycEaBChj5hftwCSQChj30ok54/dOkaioWulCws3MVIHi
Xa5BPNZqlcy4uYkyr4DOSSmggM7sxo5FjDgiG5Gpf3P8JLSo1uUpPAn1q9iZlyWtpMhFpYU+FnOO
yB+EHsccrQxRWgzM9a2gkjiohZWhEgBAzCrcSzeSRJ7B5TbO3WV+OFeDyqK8ZGarB1JrtzMLQ+m4
UFAdOfZsB3ZRAJT0QsDF8xt44R2V9SnT3uGI/Ebwg1sHsL+kPxybbmDlj6KxVLgg+T35MDMfIWiy
v+nbctkp+nsd2psFMFOkW+BMwIeCIu5pTdL7zRZgSMmET7tyeRGMyN2A+ljj0vx5L4b1/xZ9me40
mwOcfIyqwz6zUckcaJ+/ktKa7e8KwBzZyHfYvbrXJPr3XpT00fBc9cV9xFgjP9jqOF17mB4JBvNm
OHpsjr3fzNkZxrTSiFus129wEtMNaysBBQL6r2gQb0eBzl20TTiIAN+nUt42mQ/E5t1J+X/27bPg
zrGEyISDj1QohTOqRJW4DBorDVTGF+hW/1I9F93QGfSz6uqCye1qSvFBZT5Joomtvo8eL2PmNTzv
++08Vc3kCLmowkvS6bi2OYS/T9VrU+FXCfKT3d/6Mx2KzijgmmU2dZTWGknf18aowBuO4OopzZiO
5gw4AJwG2L/l0oMxa7G1CDMczVeDl19XpQo3pgJkOUYJgs418ZWj9Pl20tjZEwbiCY+JZvt52zLj
O3pxLpaOiMbuuKG4IyHUsb4LLy58qiZCK2DEL+ukV72dXFhcbb9/rgQGRejoMtX4TImc1rGAgI1y
mYVsmBmK1W0MvIk4h+Wxld1pcCTH8fUG5vfu/v2tmZLkg3FYw3emE0dmkwKlm5DQBTruGq7NO4bv
sRMx4xyuAkj/hpSOi0vkuhlMIJ3Si6kqrQolPA6uvPDVIUPOVbra6MibyLRcmdvnlOW2xE37fcmg
D2rhWR2AbsPkaxCOkPMQ01zeCSmGfMKf+DUtcxVteYXnP988Bqs+J/bp9UrE2wkqwMAt4jrhDP7N
dAUHR/X34w+556ncyGZ7Vb59pHSswh218TP0v0ij1OBB/vJkr3scWwbT1Jbl1rPHVybxalijXbog
LvpY3dz4H1E4/5KOylJFqdcnqDW0IZ7rQnian15n9PVP1NsZVn0mQI2CTyxaDLs4vSKQvFns+uA/
AKJpwTeBclvVvc1Naf+Ggf50r2KudzcV0igN5AS7x6eVfreP8jFnq0iRTO4VNOtwCvzxF5D89a37
K7yIscyUaAKXZ3peXCrmDCB5dYP1mNarLDStN9/NEDldPhj2XGfaW45bdCjx5Gsy9gz3ChlLzxM0
AjMNOtK2axFgIaJ/TnGKb5JRmlRTtLLpQAmx/Jo1EB7Q9cAQaEDMaTs03jRdCN/hEhUlLbCPQnkm
dpuSCoNg0YydzABW+lB/AaTdBm558S1q0H3KYXv3CAlIavKZVemupIlNsKXB3m5l1sv5rPsbQgp7
3C3lx0VwOBCP/mfqH7bccaiGmXksRFrPy0jA4K6SNS8d4rXFyEu3Z6QIwuMsKLF9+WL1BBzI9AxZ
pZD097WNlCXrJnz8XPh/1NdpB2goPhScXaYtguwvd+TOwHQImgzQIx4NOo+lm5FK2zbshBexamlR
VdOthMWoGLotgeFgCp5TbVpWZD6z7Mdh7a0an7nwiuBY1Q7YiU3SIpv96mv/PHBR/iGxP/kTp9mG
S199GkN5qhvm8gLB5uwpRT9xldSD2TV2twOvJJU9I1SBRVybENeBbAIo0+Hdiu6Y/wEbxzZ3vrXR
T6ey2x8pwxukG4MjHIEXhcZdl0WMb2mjtIh7Fn9KS1GwoFAMQ3JfdKJvo8k4lFBFlN+vaCC5iww8
IwAVc6n3FXCCt+J9Q1O6BxZwwu7iNfyJ7mgxqrF5HZEhey+msuIvFJnFkFwQTqKd1QJsN0TyuPtK
yNEt7MkDfNrBOchC32D9+ERERTneWObRBP/6fDWCc7SjgcYgCzVTgCGJQ3IsOWhGLY3Oz2083bxV
SV6S94odD4LdnsRdPJeiONdbDz8tsYZuW8bb/DsCn0ravT6eoJozaWiLqFSXE+/j6O6odh1WzRUp
j4fo2Lvi3eOCYtlJ9xLOkPo2j7ZcA3ZZT9mpvnTVIrVUfl+FemHo1/BMQzwmv/mxjXxNYpE+DZ0d
yJizsVeQiAoFqo1NbJ52HcPbD6L7191uY3sL9LYe/tAmb2CPW6fYHiQ/aquxr58mLKqLMUNiN8OJ
3ojatcKmBQ/ifK/AfWSB4MX8SouGopoHSlFnmzO4OQoPog/5ZAywJCoj6ae/9kClpsp4VRnU2dJD
kFGylY2btqfOGaK7hEw2qX4IZgCFBBSSc2ZbWVBa0dq5EMRSbh65Ph65VBfz3U9/8xBj+Vu8EiAv
i7yYsVGQDf9MbTWPfXinJ3NGZLhNFhfLr4rjWv22s+cOSD6JwKJgiZUdtjA6AlKWpdnugJ4aPI2S
/TZqxgngvgG19xxfHTV9iUJs1THcu7YxRR4ILwtjdropMwQhK22Y1pebKxrvZcqtaMV/X+N2XHMk
/7Opnhqg58bUSQonuT7tFWX1JEchwTHff3x1XImQtkdEf2FSSiT7eGVI99wVXaNJqR25Fzi3gUju
9JtsASDfRFGi/eaHe+17NSKUEypbe//tXDRGSpZbu3hVFB+QMFpyPC/J2VMbVTTsW58CKmKi1QXm
OF3dMF1VAIpsBghyjV/5T2+WzEAqK1iMxnMS1GlXk78YDEm5CMEbXCrejIdHD1r1Xi264EmtNrBr
uOdb4BYjqo13+R6Rqcr4oyCw5SlLNTVe3pNxqKqXFi+mg/TUJlzl9DRN8ED4J61CQYw8aUkuBF8d
qwXu3S9/oMEi6WNwU7ZLqWtfn+bkeiekUO6I4jrgEh2RbmlZPZRgWhttONw+WtERaRibwmkxOc5L
vA2dyZMTyEJBOeI48QvxBPB/UKyqwDtdMVdzjNLjv/YNDPeXkrIKbO4LNPmFZO/4as07G3UhXpqI
7kdZP5DtMbl1bfDJDobyQTtBVTCVYj2zeSqoLmOUK+u8XMvCslr9/NqRza/hHVHGwwxHP0Uw1esm
7moPKyeszyMCBLtCd34B5wpr3MiuWRKUr+Wq661+nEIgv3kZUnTSFGqcsR6696ohMYYlZg23Tqbs
xHirsfeSvqGIxJXpd0U2ugiRfi+aGhxtOObYXMufj5lji7bv6lwwGFog1gci9r/r0D+EK8p5pMb7
wb9+1RK4sa2OqCSb55EYQnE8wgiBUdA5x+vY4iT+enFoglPzAmy4b0GIoHjcXBnAdUzeTSQVpH/l
0Av+ks9g8TIICKUXSbul21TTnbjaIdO+tOi6b2uE1l4ZhgTl4jV5n4o0+L9XwxciaMx7nh+i1Ib7
6ApS9oD1m/JrihppQr/D
`protect end_protected
