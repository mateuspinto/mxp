XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��AiN��Q���'�A�qȦ��#H���[�Q����Y��"Z	MBq&�f�H6J�9x�C=��%��(�V�k`s_������ Ԇ��r�K�c��ԭ����f2IqXDܺm�,� TLe�<w�3炑��*|���I6��}[Ѣ��h���_�Tw�^C��93c�ؔ�GmSbr��j�Mt��l8�?�6��i?�~Vuo���F��>����x4y#����<Pq0�>^�"�������o�o��d��Ӏe��70���f*�sa�i�L��!��4O��@s���Wc5��!�y��=-�B���D�zØO�0�\���c_��C��x*�e�={�C nDI'[0�bj{��L�#�}�ή�ٱ_���[���߈(p>0<�1f����@\����_,�V�T��=;����x�^�r�'�������K��U�h&�C5%�'w���S޳�~�EzD����L�@��4e�V�d.EC���/��ю�����l�R��=�c�qH������q=�v ��w�)�w1���X�{����n�>���c[�oq��ߵa�5������}�=��+Px�����Y�%j3��n�[��>h�#�"������<�޾�g�5Q(mi7�c�i�6��1��[�,v�M��^(/�$7b���J�a�mQQi�!�hy�{TըX;Ny
]�	�vxQYz��<&e��T�ދ�U�e~&�&��s�s�L8;�ke�fL��HI�1��Q6Z�h���A��XlxVHYEB     400     1c0�����jވ0��]/w:�����g�,[P�+`��Xav��	B����.#j_s>��{;!���7x���}&X��C�P�x�o��-��f
Z+,G�nW���!�-���8i�
���O�r�����Ή��bM���|�IH������ܛ��~����ڎ�m1������p)*C%w����o��im������Iޠp�=��+cE@,c��OW"!��;�9�c%��  �3�/��oe�%�r W�6`�Z�A v�dQ�������U����Z�KG^��/���\|%�	;_Q�E���q5� b� �%���.&�֏�{J��$��>1��.Q��f���upo!��K�T,��:�M������|��� T ԿF��R�@xJ�WG�<]y�u��U�0�U�4��%�\���l��x%���1���n�7�XlxVHYEB     212      d0��sJs�%;�I����W~��-�Nu�����X�~�?��-��ρo��W���8��n�Y��F�Kl�8��?O�A �G���=�C����+K*�����RGU��$1k�w���G�7�#�3�o��_������da;n7٪�m��r����������d+���j�x���>ͦ��N�(3��n��\���@2D���UB�0ǩ�~