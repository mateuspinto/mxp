`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
MYeFQ0ERWIf0ERg4dWnXebyQ8deRdk8Bx9PsR/qhSjX2jyS8s6r6IufbUOszztf/fpA3tQmvqQOF
ZTZtVDYAVWM10pQDZitiZXgMu0MPNTrZH6GZf9QjTzwFQ/D27Vso1NivVSwYSnhGvxCWxnnZf/iC
Ts+Fl2P7kM+tKgBGekp1ZBoXQXLICHfxdi7QhO6jTINCAoNNRNGEiZ82F/tad88DOn/cT2JMMMdl
hNIIqsVaU/3rtJulztgZ9NCpdGRGf53zJCwdyajUCYgL7basND+O1+vDGxkJYlqA1F3rQseUGtBY
tatFBoFAXjC5DEcyvSq00fBkXsiiK8DJ0CRfsA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="Bf0Z/vzwQoGBk93N/lT2FwdixbsGzWEsD0m/NfZVZbM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18688)
`protect data_block
YVgrJWFZ2t1lXuuo83rXybY1yMbSRiytN3E3At6XR9bs+eYhLafqqJyNYcGMkSTVagDnLhT9Wuke
yYBJaSB4hqprBFnH/tXN6NPmAl8maEpGJmyMYsqJXrBMr9VVF+ycPNd0LUB4SaREX6mRaL76aHl1
yz8FndwWvMAHauCyGnFEMhcnIMRU/spSvi1pVdRyrr3D4+5aFMBB4pgYaX48cQ76S3Dogp0lHS0n
4SWntI6ZW60eYIZX3GkNO4YUrKXtDWWFyBg26QqViPqt+VgJnBtitLS/t6Nf73shrWR0p5sXLFOd
3FXEGAOyVUzCiOgNK1IyUvfl8y2jtQCbBqGglMAcCUHqYhJfmwDK4P0jZJzaOTG2kYuEaGgWSk9q
p3oXvOgCSqXHUFJg7e5N+s7q76eU1jB4kQvfNnNFV2VuWrx5LGKFZdW0aE4qp1lJWhaRPhgIly3z
0asBFoGu3wNozdXAuqJEycD6NazA13oK/4Md+V5Uga1v9/ACUupWhK/i5n8Wc08QewY2N8kkhRT6
6M5iFzK0Ssgk7PLA/JVxYCauu0yo6SoySVm6CwNCh4So1v08EKw1Lvye5l4Eu/gnikBIL/J66Usf
vL0Fz6iV7ZtBdSXdjHmarUrQo/iz/0mI+Mui5cN6Q6t8VOopJhCYNN7G8fFMqzNgkV1aq7eg30hB
r4hS8Xy+lKTBPY04qrDuhNY4Q4dWcAgZ+w5pEo7sPSgmGUT79EBbAvsM6RhWsM1T/+hXCWru1vbf
bsiLN2vOQcBy20/ae2U+ASHlLCBwjlj3F2JaFPWLuz0VtfcegapOgtxL4jQP3QF0JB8lFiVm3P1T
vAgKoUe/o+s7bEquHSuO+QixHin2CYA/uTOw1sAY3lD0iGqHSR7/v+5eGrboGBzft6qg9GyIfLIN
lfAO1Q7ptpD2aEQwQD6Su2hReIdUYQmLduHvlpvk4fInDlBG1HM/XgYlnL/LeN8sl7BngUZg1G30
Z4S3heBh/EU8plwtDzDmWjhpf6U3gR45pL0Qv2Ju+wulfQkpgB6M9k0LzVKK/FtJQbfREkMBObS5
FZIRYxnups/HX6Ga5WugLb0/27VK7n7/brTT7cdLDj0sZ1P1pEURv3kdP2T4jPMqvdZVKVv/C8iT
s8qCbpfRFbeG+ZPWJgZBOHFxk49c13CWrH4CHoKn3PnmTW77IqQNKGsylK6IlStJKicJdQNHLV+N
akI2Rs2cfY1qEbXZ1iWG9ysEbhSumn8drCx6+AlCzzrc1HW7MtQ3Gu0yXsRZcEnuvr34hulh+jPH
P5NAFKRvZxstlkOhl2f1qZ1hlVtoZZrvUWLfH9Q5y0WNcC49j2AmHlIVz17O6MXeIg8+TFJlUz93
Lt3BDEHGtxj+VhIWnYGIWRsEa/UIXEnqnRtUKXWXzzFhDe4Qn7HlYVGenNftROoY7LW9s/Rj2hA2
L+gvQe9BDqHA+1VEMEMyALA9IFj1mOEiaxWcNcdnhNVOI2XDbjPB70pWeVHT6kbdqRyum8E0pMYS
QhiCXITeH6hhRSsDRA+ZvgeTKMRJWWl6bP8hiRFJzdUZyVFPqSKEZ4xr/k5oThPM/jOdVTiXQ2PK
V48y+XMlfyWj5VUqqgpXLgdGvkryNuyP9RQtVgO0bbV9RWCz+2O6xgRGte+GfI3s/42apEuz9yp6
QDKiJ0nT1Ap0VPg78n84AF7S+qDAehJpQJ7var3+sK89Y0U8R7kDlD04nunFJQcKlQfVW/lYa8EV
5F0/3NHpmyenXy/2Q80cRE9Ts979eW6xPT/USz6AVEv9eOyRyXApUeX9gkYbAMxqUzvCt7rZxwWm
Yw2qgU6u+LpWckCWtA1wkeXoAudO7TNRH1Dweihom7fGkhrRvmmcARjgOI+/bTtuMEFLXv5/7ENe
I8Vo6YnYoIDJQCebHz/SwscjmTVKEduHgSmMA5VX/114nlEa1RND+G5au8o+83+TEGRelxDo95fI
i3qaqSKt2d8WE6D08mtZx82pPrVv2XoEjRwQNuRUb7khIqYnOKPCG6v8f8K5MwVVPCDcN3jjXazM
GAvqrF5FiAmzPnZ7Qw8/Opl6zs/gdyPFcSUhdSeHRMsuTZrCqEIi4RSx4VkdOuCCLgnbEx9idcZT
Ejj2ttwWLqa0zthkjN3UWZR1PcxwFpyct599Wk0ngtSjpse0e2xz1hM5ffYHkBp595TLJmAuadcQ
ya9VRXhf/hJ4gYGACYtAmn2rROC0HqY4j1moejLo6GPUWsMkHNY5ODgXG64AcKvJwD/aC6ELh3n2
0Mx3STMZKLTXx7Kv6VzU7zivUJkCKIeIqvtz5sbX1E9NZVDoBCIN0Tq/nph6s5C/7bwnBpbMVkWf
XjGFWwiCUH5si8s0Y5YlY2ppI3ZEWhC50TJRVlU+lBntE5m/uYlzNaKKVotqvxgUWhnp/f2iCwNb
zVM/ijMCpeW7hnvZLBn8pMckTxZW+akJoM2uHJB58DHKUM1LPTLWt3CyCLu+o4dTGmqzGRN7mvSn
zkXqjkgGCetvaRn+WWHRppC22Ry5tSCcdFxHphsUiC6wfW5G0NO/l1nqe0kHv4aY9e0kjxYzv7U6
EreHtEyJ2AtUNAhMbZUp1vFprr1K8KIfQsF0ego9ehNd677+0DUWIRYRCGHxKxe0VB//bkZ5ssCK
rlfuvxTqHAoF1Mg0NBEr4JmUoLOZXcHBZqNhmBb+1Wx9FJe4HfJn73Ptyu4AXA5EFQwu4dHgsTQF
kpyj7qMX0BzMohBAeZmToWxf15yPgqYgOlDtnrYUoTz2klbGJPGt97SgOvghpeYHOAPkcSJUjfCU
D8OKh30PzHebAq62r+EppQLhqsRcaclN057RjaoCPYW32TufHX/XMhF1C6B05UWkfIwBGoR6VWKR
kjx3JjkmcacARC1Xd1WfdtU6pENMs3xjejtQilNjHKNoNNJTj1CDYeccwW1XhBWSNKoJknw9GQpw
agneOQ8uyyHTNQYsOhm6ILwyzo/1a6T8nIje2lvzvAOrWpRBlIQX0jqftl9SySNWnoEX5kRxNUYA
zWBYgC29O2D05diXhRaN8gFqSDd6RXTUoYeNVblR4rj0+/NIcfV5APlfs2OHAW2TT70H1NDDLxri
9oRchyyCz4+3OFIIInT3enOS0KpRAUuH721CW+s5EQHC00ozd/Fd02ci+e2Cp7kOO42chLNlKEiv
bFkdk9mXAsstUx5KUWTdonlKVh0yFi3UWkHE8Piy8rP1QCKr23mNNKvdvY0pgMMFD4oUU4f02VLg
qMupQyTFoCtn3yCIl9+DfmMfJeOOYTRkLu1CUsYED0TESY/doRaD5QWAhyBJFR1bCMasJYcc5loK
LGlPP9xpqVXxilNao5Hpe5alrYzR+PTyJcCy+QKYM+Xdmaw6vsbhR6KzJ0oA1QFZqgnQ+qz+ddAh
j5TgwP0kBx/zEkrLle1Q8SL76A5eolvV8Nu/lWoRKQK1CE8nImxFwDnwTcUYkuV88sFCpvXJaKLN
+dQk9yGNRZpP0Avvwe2i+IaDu6GD+FQKeAFLtRdZB3Pbf0LAGtyRpRmvyDzHT3uxWz6o1iqGMhip
d6NPwhaFtjel1Sb6cOd68UHkiloiEOccZAuM0gk2hUYuhnQVna/2i49rY7DomI+fQhru2SN4e3kN
qWaoNufQhdB+3Fcjgpf0H9cW3suhIUFCiLQtBCm0GgOTalIRWmjKm5naQVqQWOnF/EkIp7X3Q3zI
aLN5u8/c55BtiIuG9hJ3gR21n+ggXvKM0p/DHN0HYcQI8aDFfxL9P0kXSSabygZOl7GCo7BkCnLK
0e2EDTlkdbBWn1UeSIGJhwoWsGJh16nsf0/Q2azBZETWXZ/hy+7wbDq0ru4jZV8hhLYunF70KG4I
0xSx0aFgZ86EgnObqzF3SgKdGwaUAxebzvL9UeC4vIenwk6qtlZoW0z4Hoxcho1gKnxaD+DfMFUd
gTBR1HlihXCj+yFvppeWnZpsFJw89NhRO+m4gyS0HPn9Hqglqo9pINEqUWZbzImXRzIMBM5nbrC6
/Y1nxT+bxAaWY0FJtxfvMd4PLEFPBdmRqyJmEQEwqJggi7WRWwJfKFbdMuDybvxGC5F529cv0pkT
dID20Xq/YkpDnjCHjB13bIjeIhj3anfONM8F3YKBACHn9wPr4Pmtlyh0dVeBLdctQEsc9MZ+1hdf
5k8SWcE9TQScSb7EvlCCtQqBli5+YX4WOvHB0fP0K4tBaP5QxtKoqfPvN/5p2z6hyNwVed4zRmg4
pjfFG7uH83Bc8ErMfjxkfE+pnwixfXQSg9bgyo9GKNcLOkIb3apEER7DzS22CJw9WcN/tSs1coZg
+0C2l7SR2hbz5NFAD+0twwRlzq7dlSziAZldT1DKZUItCB6VX514jR50YjUSf9PDukBp9nHNXvCx
nVUD8tM53f42yKY6G6Lpqj9+iB/vAMNv23EicVmkOBkrSYu0BvtpnoGIZiJkxoYUV6EAGRXMnyTd
Ob3LjMczSZYygzH+ASVjH+zT8CWmrgoo0gQkowCVZDxxy/oJ9xYM1kKnDGB+igf7r9WyAhhnN1zj
GfEmyLcWfnFzgJhKC/2VmwB2t5I5D08wDYigomBt/rzocgNDSsRID/OzKMKqKbzwRJt489gMVQZq
9UxLnJsuZv8KQdG+1gQ96ISfN6/WL9j/wAeHPlkn/7YFhD4goRRTpu3P6mprhlZsbNu8XlflSqvh
ghzHmuNDVSpHAp1ExIdsn44019L5EJo+A/4Ht0OxMpouHfnx36edcFPIEyWu9WXvBrGQD6407Wsm
glV7qY4rv8VkyS9YnCcb/LVh53pq8DXoBbWcgRCIu30kNQ8oeImDQoBRsL7vdteiNy43PLTDRJuj
DS8AS9iksv/T3lQf37aptapaq8rmNnNxIbG1t8aMOOhD849lUcR2nbK0oiLkyekwGA70ulCe5kaK
Zh279zCdWF/4l0itPChz5py8/L21F2/H5iROrjcbRCerdEJHeswotMPZwHVanucWMqn3cXUojE+3
9cSHsf0Hht5dRzdw1cbtTfb181kU6zicoNkDXBtdHZjEjPW9qsTFi/OSej47DMckpOZ3QQJX2uIF
UPBJtJuccke00rQxVnHB6eIJvABgJWUR1vlsQOa3yVVh9InRUSpKJzgFAmlYxyNXkMP2ReykvPEy
j6mkN4KHiwPc6HZZXVLSvCnoQlo496brDYg4BnJxBRb0SlbLo3ScvwnhP/iAkvuoH1hFMAPUQFWG
fZOzBzSDvgzJ3K/Oe1HZI5I6tC6WyXwbyGg8VeNtfvJuRIlkSSIERkaCd7nvAl3eLFw5ntLTLHfU
QP4PdLQL9d+sn+e2xUXUNihiAEDnNQlhhW8a1aknGC7EFV0yVScaDR/t0/O7BZjjNI94+O7cScTw
TSvdcwMFRnnTOJv4I4AzqoSEIKbrNQTWH1JKe3uDaejzpaHrXBIoYzJmAYDzNATgUyMgTkS7P+1k
aW6oDXzqYWqs5o5rPw+NnDwBtHxv7vsL5Egcc7UkdXQ06NiPtWphgYgS2MYY7Ur+ptI0fEWzYNd8
mpPima+m+vaXMiSeSTgyWgi6jaqekjTDu0MFaebp5KF19PJCGlbxX4NobPNODcVQTV7u2HjfGYGM
QKcbiqqw/Vm2oHFxqDGt+927r0oir8QYRFnS9t6iGUdhv63e0oMOAd1UgulIX/tGn7X0Yqg9Wdzn
Xu2oLnSmhtjKYsIVN3yDODmONWux+lz/eK2+eZRE1Tt2wfxUeEPa6Kj4HiWqEWrR2IOhWnn2uY0z
d6PXT54FhcPhUDcJo3nxXZmFfR5EUjEjuBOZxLZwCqmettj2+IKeySKl6SSImHtKDVJNuT76Q8MB
XB7YS03t/JeFzgDqTygm82nKIWqkotch3g2OUOQWq116q/7SIAHM8O7p+Ilxwu5vGCVQlHBuvJyR
URffX66M3+1kAm7eK/Px+Y/3+m/bWM/iNBrAp2x3beI6hsTGeEzPvzXMBOMZtqg5sn+imnVSTvkn
U0kGHDmBDo5unYEgTgtrvDuK+gyu1hQRnafidprI91DZw7TJkf3qBLlT4lOsLPrRaWIiTFNdQd0g
B+WheMc/Bw4aOtuy7kKAgYF5sSIdfcKj14qscFLXua6F4c2zk9FGwed2mC70tSDeJPMWzYSLAwzE
ca+h8DGPMHpZdV0U5LI7ZCWaCu3ECGFh9b1uyg2sKBf2e/oeg+X5YWoyQFQKHMGqi72XK8aR31kB
/VSMAhh/lFXS/h9VdfTHr9OrBJi2GP0Yqnl+dH7hMUZvpjSpcSb9ZvSobpw3Ue8NlPc/Sm0/MYo7
Y3pdCPtKg5ojpbvUT7X/ZtJaIheF139mIHJej8IiQtbyXbuuDLHdzyWxcy7u7teaO3ViAwxaA+Gt
RYC2cphSYsiyqbo9yoMmyEQJo1gbZr15KhSOFWlKPezrwgALFclAeEb+MP+JQNM/P4yTymIVL3sE
oovjNReHaHM8ftuwTr9YnSuUCA1rRTF77+ABfcZy0D//6IuDjUdKuOlBVMUgp51uCLHTDoeIp743
Ea2mMJfmxGNbXBCpCaJR9UXTZT1XiTbgWNPZND4fpQKoIb7jNB2mH0TQsay+czEL6uKwoBU0aF77
jqh8Pk228tneVBy13LjOPgepr++/OvDwlS2ftNoUOK+qOnsgvBz/FrUc8V5m8JBN2yUvqZDb8BPm
3XdbxBGRzYp2fzMmTX8+2GN4IrqGElRNH5TM2YLHE+1r5P8ATIcFLEK2luhmLPFJBllzMMC+IQ0D
rfkBKmRPoyIIK9XHaynUan2kCCUVCXIzPPyviTCCXlk8OQ0wadO3FragGqIsR9qg3SqM96BdWmdw
5nRpGcEvHZkwHMfQh2ZM+1CrBLUiYFC0t+AGx9r/4m48xvey5n0dzThDe50YEAv5Fpi7Tdc8zXT2
7GFgj1vnz9hkUHyy0YXu0pMRddsrfWvL2XlYWUsoPOUkHBPXhb1wMORhQMoiqBEqgiZTmEfdlxxe
LIY8Ka+K9A4gPZ540fe3YUZeCCMO3PObRvrr7aNRynHwqIeAyxgrlTfvZwjA9SecoKOjNCWBOvp9
mA9seJIwS0qVgSIQNB/nhbIOZEC5Azx5dlhNsC8O47H845FcYj0q8Xzp+t6MWbg9qnmN77D+gFxd
XNC/pixsRx6KKWLFxk2Y867GKfMjV6n3ljRqS/xeoORQcGN0QdpfEib47baAbiTzW+pJznR1/Z23
NXfeEkAWu9cVCfTV1Xu9n0GOglbF5lvpXgRyIWBc4harRcMFygRjBosyTSEd+pF1jiv5TkzxAUpB
yI1aGGQ3LicJSMUkvej01twDoeD0c/WCG42WRBC2Um+l0eL5avRQVKJZhL29nWB1D7IZ3mvxXoH/
5cwwVjR3t30+MtyMIDtKz+WdLySF3MvT9manMlDHfsIQx0AEvJ1qlTn3s6N102JGzkVMJcMglcrq
J61YY+/HgBrtWc4OjvYmsXfY1JP2J2F+vTPcIh6wQefFCVmIxLcKG555dqPQBZbw5YQA7jpIwH6f
8+opG/W48IpBo86Y2rQznFvvM2m4EB4/6d8JPU1DYJzHpdKQGDLdBWMOfLRg0EsyxtAbvr2owvhr
uu9mVkCMMbcM/WySwCF3wjVgfpEPVQoUCLQXn8ypawl7mtIDsbFVnlTzBqKzqhrmuCC174pwezyX
XxkZ8dyfOxjAvtuDC8oyk9juDFMB+hAg2bIuRC3+PLPX30+R+yMMU+vLOUQdF3pqn4qOf7e34OUc
/0whT82kX0NasZE+tH03bxyL3YnlhaLb+TuucLVyzRD9JbIsUPgFNMA2doDTj9OQoKfHDNDc4dpm
bhZOPBUAdwIVZ2x/9rT/tWO929ABbCOLNql8JTlr3JT1owopj36Ta6H1K6ZJrxt8+MZFRgeojHCH
947fc2NirwFy5iK9HEvV1LYUTpq1K73ZdPb9uVZZbb/brctwJ5WvFzJjedZK81nra1h3ZoxvWs5k
KTHilFHboQWQMBTR0W1xCCSwQHRnLao70IiBmoVTgyqssJmkbko3Pfft1rw7ibmcjujzpoohZJvD
h9x8uJmUeroFde8uvvFxVkaR4Ahztry1viaKpPmw+V7I2Kp0U3jQtKHmXad+D0yoPYOx5WI5Zgun
NiDYEEW3YexwmWA8UeagvkxGW3+om4IUnYgYdPy7xOq4oYWBWxOgfcsyGY3UkKsVm+lGx/q5GGUQ
LUjFJyqZmcoukXm2Os8dc8HK63bSdl6QsvlVtpqcE7rqh7e+AZGx4y76dKYqT4DfMcOyt8pymxmC
FHj10sQvFgvKS2sPjvC8f4pVkoKi6Psnm5n1yvuS3LLfOez0BSY1YoyVdcwihjpLMtUGa1XCu98L
639QDKEwa8ffZ8u3rOS0CjDqfcgtNl/wqVJeTTkmpdZeFi9ejnlFICHRx9WP9Q+f5iy0hi1lTXlq
f8FiGacIzFVJpmtA7YXxwVSm7ONGIdfeCoh2l/RAEm8IC1GsPRPBFXkktkLX2yipwZPzQD+E7Im3
mtwP3EkmdxNEoCH3C7WSX4p77DHzMOlr8Dp/Qjhyd864SnXreRGBWQC/vV0mBURkbze6KMb7qFn9
5NCcsHit3sa1ud5lPOSTse1wHX4+59ym5+4K6RPTiG/VS5IFWELeJpQbOsE1meSlBeByOuFXynN0
S2D5PcB2XWcqGPo5r/VpVcVVuyq4FLVBYKs5hg12CqbLcVYV931heX+1kKCqpLrZuKhxIlH40eLu
wjhoViftC7IILIyyTHRpmfd4PVFyp2dbqd7Lh1gMO4GeTZ7fUNZqmHfxJg2Wx4pMy1wo4tLI3Al4
kvJQVwmoPbniCuqxPb+o/AD+voplROsGLDGThwd+DxxtoRTNEGnFwuL9LYRCP03CA56nXFEyISQR
WrP78/fLDiuKdSTzsnaWT17eS2lRp1myi+KSJwQNJpj11sc3e9A2CwKH2WuOmbly9eJLoTNhBa5a
B1QcRLn07K87lCTz9dBTEX+VnNDl/pXl6FADivFPGhFvf4pFuKDpMgrKveqJuKjc+yNy+l+xm51E
ofOhdTn0wBQLeTfCZy4SUWF4ofqOleZoc1ZyzdWQ2XYtY+5KMuUBnHhjz1RPDzd3rQrQl0VWOv7q
5mi2O/ihynvqmXic8/masGLdIR/1bCgd3lPjGJ6aa+YSDJru/diiFq8dWjSOCtmu/pKZ85I2USSR
xn9LaUJHhqNXRsA7rC9E1zlJYtizNgBMn+Wy9rcX3mJuq4cK9J2wQNt9VRfO6M3Qei/RrLtqZ3xC
Omps032AwQ4jSL5jB1gsQwIE5fUhJ2Nm29+cEFl+DbqayFUJW8llyqy95TD1AxqL9BSWh54Bo4tT
t7lPtB3XEcOaBPa3A5uFF8UciAiLMwWTwseOfC5V+JcYMGDi6zInHHk8Zcz5UdCYGpjyljWdSVa8
bs4/pDDeHS0SILbkxFSegZHcdx+seh4TRzRrFPpAWdRS3lqs+SmhrC7OXCgAKsZF3KMRxsZsh8g9
LZbNX+IFAlngM3JlMNbFRhqnc9WtLuz0+ubQQ4Xk5Ocv7Hl9SPoP5f0r6tAAH1fMVRUO0vBgIusx
p54xKfXkfotGmwMxMsUlJ1f3vkw+a2tFnqiVr2H8r+wkFQFtu6sjO+ro4vt4tqR1IcjY7oAPukQx
Ef384wsq2HAOXkvSTJ2Hg9fMyw7s7ak1QXkxQPUq/v+/mLTqzYJoYDmbxqAeJxiQ+Zlhcr/0/2sC
IJCEEPFpmua2FYUYKQG4iGF0VOwuXHzPMOYUZ9yMqLLz2IchTRUF/lshHBGz5eKOEGJHWlgzSyKW
+R9sgc8Ui/FRUcmeRJLMPAHfO4IJcBxvOGfA5Z6Jog9QPuhRKNNtAHLVQ7udXT9ki0sGlb6jLfVT
2w6DorX6yczW924aaniyxzkYLKP1MjZu2rtYLkNCoUpbrht8TfxG1Z4g91gHWmtl3fW+JEKH9hFS
6FpaFnfj0k74NH20TX+P4UBVatCqckU+JG8Kvw5Xrcf/Yqwn3iyHMCC043Q7lSKwrt9sp9LUmyXU
MD1q4z7SxHu/6NNQMEnm1ouMb72KX7/dWvCo+xaMuNfP7ZtHpGdR/6n6t4H396ZDqx3/RdbvPGCl
wC2rukYmw2mDop4r7YoD13bOdAHhGZSnf0SKnE3QCa65F3+nXoSK1T/Mor8kkoc8G041fLs0bssC
N7VX4BYP0LDenPNwrUROOtEb+N+NRds3bcVvuytZ4fB24ZbNduQRZekPiqMqEFnZj5VBa7D1Fth+
wm42Pe2YrSZfSfl5fQrJ4NumrM9y6zU4BIgOra17wfybwrv6ZDRJZZECaOyfzloyRljE9Txi6XmC
jl/o2rjF64Z8t+HbjXTVeSn6Ul4pkJ5NRNuF+xeW8ZpbkIVFZ9IZbwRC/zrndvhC6HVYNYssDseW
1bQcWuRBfc9RvNVV341aKk4DzFRfiJTGFgcjaXts4sBW5VigrvYJhf2ytE8IlR1ocZlPZHM4wbfr
qOfR4GjlgiWOZBE0WeMMlFJ7B20LDinVz2ZtGPyFxe2xuairIUc85JKu9sJnfWnpUlNhCtzxHEd2
WmZByJY6fMlv0Dmt8Ef+60yBnoJSEjf81SQdbbNc3VwH3VB7UBfukomKiM/kjz/0oASZylJFvByA
/bSlKoqg1c3Cg0/XaiONkc/zLyk/BR/wk9OKNPEFEvKOiQwD83k1LG7dHkWlDuAzJGAvywIWc6NB
UJSzvyOhCja4A4XVRLWPoPvBUGTqUCZWX+j0QsqMzyjSvxpCKyzfkIEGR3pgAafMBRH5HQcLYLLi
G8kYPAVVBD3NMi39Ux8Q1W1tj7clNobYYD1qyOitjczmxH1/O8Nk7cGYozWuHIMiJUPw84o2dvaJ
Bhy3/3WGHqMlCwoZIZ67capB4vxnQacw5u6pigC6aHYGe9T5/c0hBlZw0RWpHGPS/HQtTvtG9/Ly
QRU06DKJdvyOtBwaUuGq2TonTyiC5jPPt93kwgmOb06mahpTI/vdBi9/wIckpd4ZLflXE+JT7qbd
YcZzC6Qs7Z1Lov9PlFoPnHSmin2yoNr3Xbcm9k97LORty9unKzgj8cBdIXvfMXqL/jDyUQj1beSi
c/myBoK+MEZccPBaV/UzR5Q5S+iU8Aa+LJoTr7sv7YpI1L8m5SkJ0jbc0V+wfT29zPHUz0onbnJC
Sb33PCFKUoUGJ0VJa6Y2sAJLaCAHMnIqEc3hmXoDsLtlJMjJBvLNu/1QFl9g3ygGfAXWpBTtWRvj
3XClNtLkSWe5/w28adti4csqnYxe7GQYsTmxuGLn+Iop++c3zrz822qOnGLXpL2SoJkkYDXr4unL
O4l8rMUSMozIXH2abGbwOAH3pEfQMWTk27kVjMa/JmVmmnoMmCpzeKwCR2lqXhbOYjHskC6qBqRU
MrIXyVorIntUDK3hrWSVI8w0VZd3OcKDiia1rx+6rLfAikiw2cElEVjzgLa35RtIR/3xdIB/npo6
hSv2+20kQrW55u2SxzZHPnmml3ndSc4tgMvuYfMdV2gkQzkd8pFgnoyVJayVwwHRlv8U6FU36dEB
B8z6gycK12rX5qP9WHEW3CYWlu/tgb4bQyb8xsEwRHg3aP7LQbyM0wNnu33Gtnzq9dd37tCEI9JR
0PzVbKhw8DP6TRRbty0FRIbn5OHoqdbpo4EqQ91Y20spEzlTYUHfuiGvhLDBkPtjf+5r9Q4MAOEL
tq1929rlnkouVh6VWMQhsyKBfc4MrRV45ch9L4UCoCueck3hbIC8VIzIYHGIvNlvUlYV1bO2VRN7
kJu87rWf+iDQLO5J3saLIPJ3+zkpBIdN5Y9+VQDFCHpy4VDZVkRcRnKY5p9mYkE02DuS+la2rsLR
ThsBmwBM/cEBSoI7UZIGS95KclVmEUYsP0TImKDxA5yGpFEXoMvahuKQ/qWjLx6RGsih17VsnS1w
F2WAMJClqAOaSUXb8I366j63iOIxOgsJuy3LsLrOHchBPVPrKa/DFQDrHJuh+DU2j6BP6yE36PCl
CleYb+OUZZeoSXkyN2zalWkLsiRI+BjVrnIAcZK20K98PPC221Uiq6GKcmR/ta7XU5XUKN9qXnKY
WPR/8flOSJZcSNCD88TKuehHkI2L8/IdLh3bPcC3gFB3WzuqGqD0fup8KTYT4q4jZ6DuRdlILgzN
DLVqGjXXOtwAEu8YAuAA3oAUzyyIn4koRXtbDivJpfitAQgzSyXpcudCp/+2FiuuG59zom1Mayoz
VnYJPSVBfQZSuL6vzQtGKlFwunstGW5a9gGOrl+ijMwr2+L84X79Nagm5lcP0C230ILSDslF+G/a
8f3CnHpGYagggJYaAu+dSLog359xJLNzjyIN7UbvvE/hRbkbBRDRY9QMCPuB047Sw6S2hTvLFizL
nqkmc1S5yqsLIHGi3cNaZAl6k6nRySm2vPfsePUgP74cTLEEEPxnPVks2nQSVgXkuawm6KNMJBep
2xlvGNtnLzuXD/8XXjl7H0DKeBsPlUD9x0l8fvOBAIlHfB6QjpkMnR54MaaLATq3+NdiZ+vpiO5U
s2E9Q+ok8Wkht6WF7YBVGh9moItVjhzEyvb0Mjxx6U0Ehvcnkvtqz+wzI2GHM+AVhAcXk7/ZjEKe
7TVTvPEDyRaOat9JXT0fSCZREMXIVSyt271VI4iSx0XK35ep7AePeHQ66EyasuPXOTMAy3rDpANF
/a2L+KsYSuqZwXRqOy0o+Ly7VAv/VbqGIiIUIpfEH63qT9icLPGs5uNCBo0QaYjPjocOaO1r0+9b
6zc+XVMSL+Ycc1i9n8A6T2Yc3vNIpL9tPxTenZjhwSb4MulknM+5uc1KouoWTS1E88h4Vtdh8Jq1
MUjGDKMhexPtxUkveFHEjRMhnzY6PdqkYrUMJGULdkZLg7/JVgtL2wSKUAfTe/efDjwtNBRV19+Z
qLgbVbguKM6f2lXhAy7b8j8fX3fr/xRO8mKUZLZBuSh2wKRQfV2yqzWciPv2mMyDOHIOHM7ptAx8
fSGjcZ4FyoVCEVyyRq7rUjI+LUIeqVH/io2/pOOW9SUvLxYychFkE9qzbXOKOuWI6Aec+BbErAEh
cfj2Ey5wxMkbAUH9QUmeVE/MwzvjeW928gpLKavVOrgkXOwqac2lrXI3Bnolvs5/4S5O8cV5Xsw/
XhbDSGuuTEOrBs6DiDkDxLSMuKtWp9V2mUxcZbM3YtAJDcrKTE1X80zZKVhYNqLP4dJtC/vUzihg
Cpd+4bMjIthHJTIx6HUZ9pZDFtFPEKfJf/8Kb3Hv9HoUFbSTZcT2ptVA8ixrKSrXICYpBW6C2jlf
R/Ialqd05EMnxEzhGbCKrWb1AbkHUQkdp/JvoK8lSeG2VJwCPxOfWmLwA4BbLVkuxTOfsrGT9C9G
7ch3i3MQZ9DvUhFNhWtvsv3+iDpatkLJG+blQR64dqSi7I535Is1dsY2BmXnO5gYp3xsHpcd9bk5
rVOBxCzQK9xTcDpsiXiPHES+hmAD9GSuQRQq9w102ee+L6Nx8a7OHP2pYzUwT19RBaOMhxfail/Z
mHqMr1fwFmp8K/6F2zaPN4awIRPZtd1yoe2iuaIEwZNHfI+9I+hi8sSIBxk+SrbDPfprO/BJqBLi
U1ZOwhir/EOIOVqMuzY8KEXyGbmrda22LLoW168IH8FtzBK/96kevGs1oZCn+FaXi1nWjme9WcgD
AY6kmSHa+c8x4Zgm0cfJUf1pobKfp+3e0KacKCK//PYiOwJZMwLxftQTG6mMP9ExRBNep/uoAjAi
9LTKQX1dcqfyvjDcND2wL/Nt6aObRLyi5/Xzls2Yl6DWH9lj1ZcTenc67ZatZLQtSboiti4NQFu6
lBGsMrI17ZcZIPbGbmrJ17sWrV9vAQxsolOhv7MvCUBIkc3PcPZePFxJswznr8btztfXWtZvDFvB
6kpaNwABqS7hwhsJSsOzQuwCA/2sSZMh1jvCU6VGp+BNWsUbelM51a1cYy6X8v4FEWgQjEgabUWP
fw4mKYx4YAwGHh0N/FiQFYiNSabGyYLVzWPazSqrxZdMvH9oyvKMweOMGb6RdkR+0rEdH74XoNm7
+cTZJ1ClIWIB1xIY6MZDhf0eg0YvuxkJ4rbQ5YUGgVw8RZSXpfFa5+90mG6DuTnbEP+9Ut3c+bIs
EaFTaHxoftFN8VlMRsZSRMp1RaefYyvemABX+RxEcuFMlspL97Dj0C71CYQhxVswspAquO0Th75o
0WWOTvwBkFQFILqiznFBcvItWCiFAodlYz4Pq8wXFhENrzKjAWzl+iMywrOtCS5ykFvyqYEBKILb
Xs1UFPRDBGMSrkpmiQw611RonUKAt2XuAaXie2EQhkyx8GMnGUGxht57+IiHhg1oECIDX18JYcmL
oa+zhyWjLyqRwZkwq10Jxuf3lcJB8jA48Y4LHa8TWVJ4E7K+fxI2O6kkNubejEDQhOMNhD2ShWMU
XxuqJCS788/L3PM4tmnUQ39QSdwvimK4JNh3d1+bjiQOhZqpMpqkWX94DgZCXZnTUBllHPNsyJni
iRsz0yRc0fr4AENgSNWdDRK+PaSR3AVpwRzfl8pkAbaEyhWN0xZWj+Cs7e9owDcEA9i5FRhonWhK
zg9JQelKjlLL3YG16tFRyRC8yb52CRjdG/vZJ5VjNAAVUEiXZt4Hccq7Oq+2Oy8ZJHxqO5+eYodm
sQnEODjOAvEklVeUscxECbcWpQDlOimL1cPn2NIJVK4qF5u4IgQFZa6K6P4Z85e6wo4f3cUgkycR
FiaJcMTFD3TjdpQOyvvFmeOjON+TdHSM7FKLVFiL9P+HGPimeR/cVbBPS6QG32hwIrr73X9V/kTZ
ISm5xnuktwD63BvlAjG3CCt1+3wem7t0atz+Peixua91Jw5Qwv2s92nrUvsdW4dN/ampy8QhA7NP
wmI/5VbuaLlBEdhk6OqYZCGfujuRpAxJug4oAeBKgz+3sToFQXuT8sbHKPI4ZcAyHFnviyCBIKsn
5u+NY7jrfrHO12nDdwDmo3ils0YOhcFXbJtlumkFmyXNSqdjaacjadGe+3RC6t2OvAjXt8qLPm+w
YiHwv3eN9j4OHpUWhWS/uDyZLL2KBoIo5XSGobg9VjMw2etSP2n7f12eZAqhnQHzdIxfbdBTahid
SUwqxvXeddCIb3qtzN01QiWLoqvMMt6Us6nB+EQjMXPSCF+pnbZlu72ZHcoQyybL/xN6GLvreMlc
bAsavQ8F5FLs+JCMJuKn5jIRIwdIzlbCsrCHiXXTSTnZoyLi9JuGuKFNzXH3F2/K8lBknWMHJK10
W4vVKKlc8lOwep2NVnapfzmsIF39tmDYtUcKthVkLdfoXjL0jXpkUwIRHZI83JWDddx4EL4z8cI0
b+4PHqz2a67IQy6vACDPkahieJbHLjq4uVcmYTjEwOSyVTVgeTBtsrEXviyBhMX4Ddf82Fwq2JsU
XTNfKGCwmjrMTSfoTqofHTKaeybGQB3VSHy8EWYHgtCEg3SjK97JkTdkdARcJRS3Hf3Gtn2uOFm9
m9Ky6vAsVSa6UBFXnJLrtoJUGPXDhodi7K9nzFtbV1Ifw+VHVEvRkGGjY4hTRL3whUnxg7GlzaRL
/3N+b/BLfv9edf3ITpYAK3pktbRGt8/+6pJy53/VaoISUuwVR10BMxCykUhCzfQdCvU1apAmCXDZ
ycUaRG3oVa5iFuUV8F+zmwMdsQa7i9D1bY+TUyRLrE+V+OYuIh4UvWl1+K8tXrZpcguI/e5MmWAl
HsQqGeP0FKKXv7wLo8DtLbG8dU0AF7hB4mrY/D37i3HtPv5zPtSiKybsc0R88kTbw3Ub6xhhvr4a
+HhaBkG+5RgYeWBQ22rA/ZGKIml1JwOsmKklGcCSWP4c5H2CkGjL2YsTWW9tDsQ+2vIuz1NGKd5C
SiWaxQZgT3lE9Kb7QuhNt9cIdQk0WBPdeImjFV+Qj6mZvZ92XxB6DbyWDhS32L3Y24fxawKVjMdR
6IuJ6i+MJPcGH+JDpEUEOE1glOBwCCKeqdVbsUVkoLpyRSA9OXegnUWPjYY8cWod5hFiX2p1P0q8
djlH4cqrDxtHl7/E2jJSKlC4YYOmtJKkRfoWxWUEVSVxxlfe7tMrcIYzGn/PV4z2wcygV4w8k8Kk
ZOUmAvguIle1QsUZd/XNE9VM71Uw4gfO7ocxdPsk7PwckhCfJ1CMGuimubpyvzmAToVH1jVOI9hT
Je2NZabwHnRmhMoB31qBn0NRDROgG5f8QM6mQNGxSjxWp4LGTr8k2Q/U6Lv2zI9N+kamdV3LNZti
Iq3CTaFhVsttWbmyuf2L91jR53uBm6F/2lkDNaV1MIJv+1qAzfiPkDTlYqLg6eRji03raovIsFwK
881wabYdrczLlXZrV/qFsIIxizl2OR3QaX24uH/w6c19jQGhBkL6k51mBtx9lg1YUfIR5vZhmFP8
vr1iKIfdocnKS03inHXJQpTB3CSCYjWzdlb6aOdUUP1zn/538tteDk6Qqol69ciPDhYeK3Ve88ow
Z1G6bL2QgP0ZYzdZY7LwXJ0DRI2fOo9MLRkPRvFQBsvu4sxr66VtrisO0gqudTf9ievtBQdQPn5e
cwV77DyCVUNKaeC0M07OB+p+7ji6taFdwshzEmuAEfDrUuZi54x0boW7qrSKlvUKYL77sEf183GP
TZtGx18k6NaW7Y6Q/FfdzyImzjEHLEeA55kqQRYqOatE1KZHSC+kAv70Txncf2DxbKGtDHDHB30t
IbPXJJ8xnLoK4DtlhywX9f5jbdSgZb2lSITD/+RlRM3c/u/TRekN5/gp3Wt9MeB1T1LLB5bLmku4
EGecXRML7Fq0EVEA0lJyub1Uyh8dmfIruorm219elu1IBgB33IcW60lMuTg6JmrOwVO9X22T6cJ1
nEe+hmtn1mXOKrsZX53gyNy2xgzP6W6NqaYR7qygjqHCgPUjrD4v0NjpmEHbHuBoNVmt2A0cs5ja
aA/2y7HJNXs1kiz5hV98Sbv5Ij3oefsyxGuM7Q8HdT39iCUnSskjWz+PhkuvJOm+RQmjbJA4XPwu
UgyTb2i73LSrgsvjOK0HdVCBfLH3LA+OwAOq/8vStYnXfQZXG7SFt7ylpCfbIwmAgsg/JsErPdve
f7QHHQLkLtGauCG/xUyhiE+GtSwuyEOdN4/9Jii7giVNoB36KgWkWJ12PQWuStF9eXCwxbME8JGR
0L5OOSL/6VdxCWK7fa/otjnybhKBYKD7o0T7GDS01og4P17P4H43TUqRGTDPE9GB7NkFMSo0W954
DD9Cpx0yT4wi5RUSScTx8u/KdAY3M4n2g2ascTaQ3UFbU5GZjzcKOjGjHCOp1QtIQPFekW0GBEEA
vxHzX7u0rSoemeip0zMHPFJGoph3kAd3qnQyYgJPqg71ieupmHUYf88/wzFQPGf/FaNNNKfRg/++
mF8l+7kCsKTNecFk989QGrT6NVQfaSWosfZ1RDMW9BPqZyHQbRDPQLnqAgrecn3b6CodPUiN0urx
eOjwBQmrp4urNrg7QJ2CojfF2b+zLd3dFw2GGqPTTNYdmIS50kR48+wRJ6e4cZcsg+FNqmDobVN7
bNGPNIlVw3+9Oosyc3NxRCBvuLNz8MfEwmbJagI70Luc7JF/eVpzu3GHnug0KiG6I9Zcb0Jb2r52
sni2bV5rzWntgeCjXwuhfpJp57clnIXhK+NoUqyNppmlBCmZDVveHXwJPhF/DXg3mXistiAsjQ2m
0IjZMyqvKEPkHCLbWiraROU0GhcbvJHErweRWsTg3WR/RnqVF8qfkC1+kQHrp4YIAlOnHYhA4SSz
V7T5VcsRUZABlNX4mUq7+hClznV+T47dRkSy428A9ow4xW8kZmnkCKFatWqXke4bLi6Mi0urdDeH
7wQ2hOrMokD7YtSU6+bQaGZJJRMT5Dhgh0oWZPZ4bRJyg9gPhafxLQkcsj1sVnz5zXjVOb3SWvWX
cHcjauAtntNynxYgrf1cY/9g4uu3wAHZxeruQtpAPHTwfNSclvBBcmR4HCEJWMUFt7DRGFfCsr7+
zZ7s82GN/EcFK45MGGQjpfAjH1pZJ8u2HlHtsHkMqozw8T/VY9HZzD6KfuX01gQWwEVafDVa22QH
UfskLFMOjll0utyXofWttNGhK3TtOvsDUl6ODYeBanTpCQRmPhEO1EDUJm2lb5bWCCSBRMeMwfzy
6ta3GIjoqvz0uB0qWaDSAtuGC2fsK8lDTQIbU1T/iKnTxn/fJ4giOAWtAWYxIZd14g/Jr7US2Uri
tuVfry5D/ALR/aWy0v7eysnTJMMdIBGaRRRWj3dcsf/gtmxzbeeZWfE8W2UJPGTtMoDJoaswkKWe
nlsnWFRKArL3wql+a37vRqyIAJ/a7L2RnGhFI/aR6FBCt9EHD4INrOKvPSrK6fZ0ctK08WX6gI2N
TJjVy+ZdpRbRE9NBp3wh1IQCU9+wf7x7lYXZb4Q/sYAMORDzfOMwiB+HIxkqZ0LfnosP3PdRygZz
28yLy5j9h3iq5GAOPig744RSDhbweGvvFSyP5kiuMkptSshII3eB2mzwFhLARpeEk/RRiy8VXWuL
Hz5nkcVGi26u4zcb60/1sOCc7/jTWj5ZDol/++mjHmzLQPq8Lb24f2S6UwLA0juCEvhRgqCvwaj9
wmESjNE5TrGCmxhAdAawOSxizpxhgZ/B+C0WSpt+ASED0aFzpPFh/Bvi8LM+4rPcAGycJmRJM44c
at+wSaVGKKeGsRYDAxltFlYD7ftSTeCC7MCr0tm24f96xK9XAdB0F2bwZ7fIJupgsA60vrM0wM2O
WQ6zB6TideSiYyWJUS4eG3BILT4RNcYnZbaT2bPg2QHsRGLC0hEm3wjW4hKKM2E8IBZbtgCf/kLC
ub834ZgR+bQvJkf8lPgOdo0vLW6vqKCEwCkgzyEX4hfxZi3gjnEGiR3bK9E3WX0MsCXt+89TzlJb
htZ66swuwtIYrNqfWuzNOj1jtRmYRTOQrDdvane1w3J01sqT04kkNl41dhMRJpzMlAXJ+cRzLcHm
2KySl6995TQS66I87K+om6poUey9vqLNDwG5t10tlAt9kF6m8BJXvi2WJ0EyXCXB0vRI4AgBM9V1
CyDnKMd8CsYt+tCWqk3eAyFNWjL0PmRJNvMfHE+oZchRVVHAFQo3doErr8fFRnQ14u/qiYQbgU/I
emPGAmmoMlYXYC6DQe/ST21Py1R1kQ5nrF2TTH8uc/o4tiRM06m21/2gVDyVwwQ26qdCBd+PPo7f
NYJHwoLenCwEnIiJHH6vhl4Qb6kkaMmVDoEaXjUiyJA4TU4jxNW+VtyqgRvxbSbt7c0pAp4fRwxi
QNdP4Ezb3ciQbEKwSfzGLCQ13PSmdDYNjOVb2Rz6NXc+U+x0dH7e8vkeBf6XZDXSty8dxjbvUsAR
tgAi4y4i/01sOsnOIFm9H9maCPsOamo7LixUN6rwn3clITYDfBk4YtH7isu51YUOD2pvZ80KtDVd
zIPQhpw/dixaWi27jlpbioewSt/3YD1ANLnaSYWZeN5dx2Nrz1IJZFTiFAVgbRZLuDeYujrTh0Sy
WsMFKvPxFwALejIKV2QKaLKoZz0HANRMZDzcq9VFZ+XMYVVDliGzOQ2BjgEvJpUt79kCH/aJoOgH
D4c5DLIbu9wxdmHWIf2dHmyAERgTrSZHXEJ94sDj/LlJXzoNK1L4424NzmfyleUua37ZaHfW4aZN
AlPb+Qo2MoIozy5TW/eGbZNtqa8LJqucm/31adB5Oj2/M/FYLfRG7WKXaEC2P/LLTT9PLpy7XCSW
EOswVgnogUELPW0ywkmS/F1jaYcTsMxWXmSeDOV3+1rBcRLYSLvklqQGjDyioJaKJnpRd3MeL1H6
Tf7o6U0gdI9/EaiC9b/Xhj8HkNZK/iYoVYKywnr66twQ3d8cyevqpS7eAvSsHVptLm38EpDzBs3p
/AIveZjvGyl0J4Gobubqowkicq1lJ6sC8cJsR7waZJcNwGtqPuaz4u/ZHx26iMVX74h+P62Xz93q
XB8rwd2IKCQqhWjFtBYNu4ou7EwRNN9/9X6RSZGeGw4bn0QdB9rH/q+qAmbMd99UEYub4so/xYWX
lMXiiCrGNZQgy/lr3Y6iPmELjQws6/nPuYSkcvWY1vz2fyzRhXWE8wzZ54XJG/IID/8r7IyW3Qzm
uVt+7B3FDotsKIMDZB1QLDDTQNoMZmee3TfcVbgZcR6hvMj6qrW3GuY6zYJJKEnZLBQb0uTCfKgj
K9h4yzXbQgKZNhgSBWvQL4T1exF6we06G4vn2pct89KOSRVOut4oQL6DGYTjpwk7peOMA5tRTJBv
OiLZud8ikiVaynvA1Y9oOyX5yNmp3eYr7ZoSSJIyoVs7zlShv71cLwdcVV0crCmQPElEBtJJjRJR
1F4AAgaapxim8Q1eIl6F1REGc9R8TqnjgjcCXbQ6luaiwCrvTGN6N6P0D9iqXiSuboHDcD3cMSTa
jBjNGlSh4InEEoQ+kO7EfZ3iiNuZCDg+GCOe1kW2kOg7Tl+x069FkBetsLUua5o9Qlz3lTIS9AZA
Slx3nP6emVOE3TupRGSYjEd1nwFqLuI3os1yd2FNT8GYpOFCgVM1DUwHh0OcniWhwDTApEicrYJR
3eoE2mAXiBZOpWrK9cg/WkQKoJuhLXk4WTjpKdh+x1N2V2squkOBcLuufAcnGmbE5v1Zso9YPEnT
XeYVix0upCjOm7R3B2ZKhJJflhcOcvZWAGWDoZpIOYd437a1+s7WZ685Emz6NnCYdODwwD3FMCbv
JHSIU0HOHuu2ahZOUvxkmIVe67Yng2ONWeOrLELjiN3VhF9olgZpMLW9piFea0p2m7HDf+/FuT05
DGwilmOMpr9LEOg9e3Ap99UDYLZ95Sl6uZ9q+Gf44EAJT5EVrq0JHn2IWZIBr5hftfWR5hZOXynN
qMH6Hm9fkPp0pB8jJrAlr3XhkGXwmzPXOr4O568KhjrBkgIS34Ujc6lcoo2qAS7gM5zc/ZR7qlWd
/his14lHd5sOlk2QcApMErcremYU/4Kb7jZwlhZxNqorcTv/Pn6seb9u7Z77escHVstWELacwG53
fLwguUeLr4iTza5op9zvRXrjLg8cWKx5Czh1eZqSmTX76wLkp8CS7WER5jsQWzLhKLsVQKVQt1Oy
M5px/Lk/aSdDOPIAYJdxPHOUIl+8+zCyiHqWwXlYgtCls6bxFQLZUK/17n2cxN22eHzptU25ANQm
QqrRAavBaE6+gEOUOn77G6NVRd/5l20eNilII23xkYvL7Xih20/v0ulMhSJ/9lwhNSgQw1xzalM0
smOQtutSjapo9BNj/xLM4UlkVLz6iwbntwAOUQQ8M2TmNkNsfHYfC+txDWlyq15Rmeo6wdS18E4e
GrL39YsiAtyX4PTANbYd4Cd22VBLsZYPr/qYzq1jSodStVSiNCkCCM98P+F+1BdneVG+LLVpRdnh
fV0HtQSdnXjSw1UJAC9XZ823KcMMN+zDil8Dk1IAwVHAU6fCGEiHIjYE27JSZmPXtNxu0i4KhWY9
uiSSJSYC9F2X6imHhltsitQ1+rRR5MemzL2PBPE9vTPAGZ4XNckgFT139+/HGhXE+eQTNnOu7DUQ
fNl4Pme4BPL6fGpSothuhs313CBgL9P/jF5UGJb4j/uBUMtBixJbiskiElMcumgNnBc6p7eMMiN2
7SVZski8MwiPJqAJ21aYmWQcZkYMfuF12GtuOw3Nlt8qeDHrlaaykEVnAVSuPSSr+r2F/770Q9VX
07gPmZH4SoBkwqHQnxrPsjHn+cLpvxhaVVVzbhAmWgxji9UVKJfZtC+EIXfu5QG+2iE0FKDbjTNm
WorynQzaZT5UriCTG+aqHIVYgTnDwyrQMIa0EJt8XlWM4c6il79JJNHlOI8/f/rK/bxPkIKKj0VX
GwH2CX2i9+bqsx5bNQgv9yTxPnt/pj78HWMyWkRyAPW0g968Eqe5qyh2OijVDD4gQukNp81QHf7z
AIbhK4DZQQw1A4nE21V5Pmy5c4Ly/Gl5EnSyPNLqkRz4lVy1WLhfr4l0zMKROBeZJBaZ7Ikt1HoB
ROO9BNo0tIPGvyPu4b2VQHJfjxpikNGisJBlE9VDK3cxIXiTLZI6BYh1mYRz4sfrXX5Nxvt1gmHu
tMEzD9Cn+A0qSpeTnDQ5QTDuCrR+faBzyxFzMFoAaLaEhm9kzsx2rEP2YbSf8AB4+BLMQhoVd/CQ
qwmd1I+mw9FPOAuDiCUPLUAUKig6TwVIk94KtpeyvrS6W7drnE9zEYFi8ES9nj9tVsmNEigUqvLB
L/PIYsnEXaW2reD3Ny2ZtP7N1nDm+Tsz0fBHJ3rAG0i5RyUGP51TaPgk8FEFDoQLJJzo582PsK9T
Hp3JTwrvMpSw4bI9+rFjaOj1JXoHd2mmzJ5z3LtNJCxS+nAXa2mBc6C5NpTEu10k6pZSaAXQ7oRk
oipziLdWtC28TLkSZfp7l1fS0yu5C2iQAUvLuVM+JCq9z1o92Pgyqv9XiYv9XD/IBx6A97RwgEIY
B3iSHjyubtCiV+kfbdbS/jne302Pg8zCsKJR1q9txiNLc1ft+Ob+NGRQfxGpJiAXYviE0tL+BSl9
Qr8GQfSbRZ1t37Y5Lep+WMzYfMnyr1FMmSRVdMjzSK8brddxFLbKssXRbICwewDj86mrL5T4eTWU
2s86OnAyrP8+Umc0JU20cEU1xr9Q4ob7jJcE3icF2VvRSXWFSfY0LjxgfxDEfToBwMafgc2zmOVM
EMVqKyqzf/I4WbTmykxF2zDRBCkLsLc4mWKsXhe+sCLEyPeOAnYQCVjhQEroim3Yme0RvL+prC7c
QLhopU/HS/vEoWrazdX3B6KqhtiK90qmooZXfCD3eHVq9r/pKbT416fMZ1UYVPl6cmDUa0r+s0u3
WaiiUvO0WkrXRCV0UZL+GRxSpCoSV86fUJuV9DmAbcKeoUBlqDN+Hd6F7aExJDHIBPHMJt9xdbNi
FM82rRgfeQobTA4+7Djicfkre6JvYGlh5bJFmpIDUpvgr621yMEHBMcldir5RDdlpG/l+Fsr0Fxd
qQoer3XRdSVcY4BBrOS8k482r//SZ93XwoUNVPr30J9G+wTKZaDDX8UP+pUzsOVIFMD23w48MhlU
zmXj72GPX7iLmFCsVmb6xBADU9pSD5PYbGLFp4sqX4utmC9cymXGbJKIpJavqxOWIgHVzyy0zeMg
bbHd8/Jf1OfQKgcrgjTW/owPnn2i4CcwPs40x2uj24mbk0ZBeukVYUp/FG+K1v4i+3QKrkTlACok
O2yGv/SfjO1+LmXjzfowR27iTlPh/XO0VCZA2Ki6AZCT5znEs6+ZD8TxdzldXr/RAtN0a45RWV5H
d5CdTlEkS9tgZY0u9N9wW6OO98PsbFAL8oxji6QSX3OvYTEBF8x2PaqPpzMrzi1ZUeWBIB9LrHkM
luoPH3yJDBDtNKsNfWGFTRnAVfVKEprwzIjWkuQwcGSKg+HRKs4WYdzqlZ9ikFMe+T96mg/Bd1hu
7rY1OhS0Sjv2YeRerw3zbu7Rw5WKclPSM4qK0aJSrmY9oH0FbcgStvPL8+GZT+lgQ9yi+BiIaggS
dcjBehf0kdz3r5tZHJacalGl5hJ7gvG3F1Gy+PmShrILQ4HUYzd3IkynFJxHTSFARaWTc2XXqEYD
jTkM+sZtu0uivALWWoAFyyDMPPhFvOp483xAMgULyukUiR4RXAnppt/X/TdGdDkKPAPDylDgGtXE
0knRDMqd/oYnDIntZcZhx2NzB12RsmEru3iVmVz5l1I+rkuNLm7a7igvS705adSy3PmFUEX5XDe/
WfNKiFQIdeyjhhgXkAZZIihqtICyHnDEk0FugLO+3+z/0ZzEo+qhso90zOpfa+G0+TFhOXBJ9dFe
SIIWt+upgxNzruAcdn6QkiC5LsTTfyHN4TB1fGlzLMfNi/TAoUHo21Lnk5oRCn3a47i0lSYdRZjh
KADr8TTcthlQYlBAyB/e3uFP6K5pHk1kfm8sVkPrCqLML47zTFbc4GXm/lw35uhwSdAR602YkkJE
cMkYglwRRkezeHXrQjhJ0n/jCDQii3x4+PIQ8u6Lmxy4XR/3T5GZmww9+zoTXGehmZJV2YUb3NVq
BTX6EDEBsURz0mpZjIDYhu5Z3bU+HJqj8OcJElGUpGaGZXrFhoigUMJ8LOV1l/gArQcVopt5KWQE
Mk5BhzNb87R29zhdW/ir2uQ2bHowesH60Vflq94X/k3c1CWEgqx7HYVEGcLpxRgUdvFYfFwtI8Rv
0BGfsTZ4S5H66Qk224lIQXOjSu/BXLnGOyJcRWUH6+Z3KXYR7JKEc7bClFNPMyHuR3F67tovbSEo
4RokevcxOxeeOhaI4wULBDssciEZ7HRbl5kDtsjywFocjDLMMGFLMbf/IJy51ZIkmNFYWRemA5Us
9IBfk94rVLHnro7ahSlKB7At6a6vexCaOdVcy4UE3gLTzzniekeBDqImw7gMCHfsKml5KRBPAE/L
zKNGGh72oJpHzKxgeys5Aq1yoZWcq2SMolHASypM++Pv7BUa6256bw8H0hMXfDWBRjuGuKJObl1d
+K/KiHw+3ad7+V02gUA10rpVdzSXKkG/tfm/8FhclA+4tanZHLPCy1FsPifsq47o5qF7Zex7g8G0
Q9jH1m/yve/ebICOC7geuqFOy5cJ5niR7ANKSfp738giY2eVjA3H5YqWt9vP6MhiYKUg9F2gOi8U
KNOR3MGp66CZ7agTClzfmMSWuPMLPoE8JSEt1QZ1YOwA6bng8M9SnJT4lmLQ6MEMGXSiWFfghlk/
Oxo6QnI2sbSiFCjy2uwptIfhxVaFudOZTIYpaV+SPErBPy7aqeZpH//F8aA6u+SsNqJ8qDPF571q
rzoWPCfk72cgKbCbZsdB9SU9kb+CK+s3hgjuJpHB8PW/sGr2XwRI0AdeZEg3kUkWBg==
`protect end_protected
