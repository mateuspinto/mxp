XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����qȮմ��2�!�h)��+�����DcƺIJq��o��f}��Sg'�:��٦;��Zh�xH��X��j�B�P���X!a�<�S��dxNc�.���'��H��%�c��D����Q%(�s��؛��-��:K�u�[�$��b�$��jBo�dhT�x,ť�`����͹���ʖ��*���w|�Y��hR;q�˜�)�`0�`1F_�A�2���tD8�<C!*[���3&��zU�*o�=��+ͪz�.`�r�Ͷ��q�Iq?��9���~kB�=� ���ș��粼aQG����fzf��g��ó{��Pb��qvx-�4��+fy���_lq*R牜?6����;2�m0�!�b�	���io�4���)�p�!�=���ێhɒ�z�X�m�e;A�M� VF�Y|�ꁻ�M)��}��1��HN&��搓s�/20��wG��`�*�r.z�Z��`�t�bݮ�B�X�^��j��]�GӘ�w�B����J������J�$3�X�Q]Rm���3��p,{ǵ�_�RM��AD7�:.l��[W�����7Z�A��5�q�^�����}������zj
��� 
^C��lDl3�U���єs�w8���G������	��#�t?�P��g��\h��d���}�73���pa�N9T8�T��#oR J�zL�J��F�h�"&`�>͢��_����3>���|&M3�-G�o�B����}j�G>�?�cuS�[Ω���\lXlxVHYEB     400     1d0u�)n�����^��%�l��x��[�_['^�T�ń�<w敛��Kg��7n<P��@.�Nr6��A]4�4�Ӳ�-�9	vJ�o-6�+V8%�cSq���ߊْE�����N|����>^W?�������^Z1���T�g8rs�@�=��G��f1dR��NA�2s
B�Cځ�E��7�C%��G��8IYw��d��i�Ѯ�DV�6�ߍn�<d&[J#�FW(,�(E�x�g�����`N����$ZGCV�j������H:���w���K��	T��|Y�3���|f�m'd����{�m`V?8�s��5�Mf��dWk�clD�ix��0�c� �&w�|�h�;����XnZ\�F��$\��r�`�Z�b�n��4\ ���%�I�9�A��rS�)���P�x=��_W�S*TC^T�\ς���<1(zpv�ޡ*�e��XlxVHYEB     400     140l�	rs�f�p�c:e3�K�P<[��h(f��+\T���8��/܏�K󍁯���V��#��P煕�\�����Ū�3s����Mo�����?��rނ�{U
k˅ZR$���8��U��h��N�@�P��CmĖ�8�.z��&C��6��8�G��4�TFC�����+O���I�������Nc`���),� ��[��7���3�1}�'
����)ڄ	R� {s�ߟ�A�r���&��',� �$q�eS)��i�T�j��iՌ>��hWծ �R	��%�u>�}���Iϒ�ΙFT�g�e��n��MH�XlxVHYEB     400     120�Z�7�&S���w)�S�ܧa�;&ax��	�5���qȾ��!%�4b$ �'A�j���?/	(
����8�p6��E����S�N�*p��})7��$��z��
���E\O�,��!UM�ޖj ��>0��)F�*'��74`���<�&�ǽ?���F^_�\Vӆ-\��7r���)�8DSf�q�pƌ[��ݔ�~��F�ZQ ����2;�����6U��O��R�N&�p!��=F¤lsU
�j�`r���ݫ�p�A`(W�Wm�V�I�L ��������

�[�XlxVHYEB     400     180�s�_�%o�]^硈�/\��Ϊ^�d��.<k�l}�tb]z�dUW �(�_�����.l�(�Խp0�]e�]2o-e� W�ɺi"ç������+�U
��@2��4gK�.�Y�k�^��G�_������JgV�
)5��b�OU��|yg�o��4��to��+P��F�1� ���&g&����s)����ۜY������x���ۜ?�>����������:G*��n�KJE�8�Q�4���Y�c���"77�x��U�o�E@w������9ql��&���@�Ԩ�}�A�H6���=e+@O��,'ź�s��k��+C�.�> ��|jm��w�dW�U�Z<��牼d#]���Kv��XlxVHYEB     400     1b0�%�yܗ*D�BY��+5��{�@Q��c�� ���b���`�9+>�-�-l8��ͬ�S1?�zA�C���O1N�=s6���*+�!)?e7�J̘���bO���a�$v��b���܊"I�>J�*����m�q��u;�Vg(��&}"��r%�l�Y|C�$#RvXz�pdt��a�I�~k�AXA�
�����q�oܣ�H.�N�M����Y�T�dR�ɤR��6&�gÄ8��3���^�Tϰ#���c.����Ϝ��+��U6�[T�j��r��2�$𐔅T%*/0QB'�~���`�0�0)M6tt��2��Yj+J|��%3����*�������g�Mɦ�Q�����9*ܙ�A��'�;�7�3�w!(i�Q���?�|#��.C)��X�	�.�U����('�#S�YS0*Z��XlxVHYEB     400     170��G����N߮,;W�5 ��&�03z��8~�e�c�xF�V\}0����M�l �(� N��s&�S}F.����$P= �+�ߴs�Y�n`�z-�(�)x��-�!��|~�R[��׽Ai�3m�T0��j Sɲb8�v܀�t���=���̺᫉��^J&� l�� ����4ι��C�YkX
k{���ga��-�\��{��NU~��h��y\�q4��$!������9����ɬd^q�ׅ�����?>MQ��w�ࣖ�J�+=P;��"���X���������x�	���9e�*iL��uq������fff��Ǜ��q�����V*�A�'���-G|�l]ƌ���ΣMXlxVHYEB      d5      803C˟&J�3�,]���F��h$��q��e~u�2�*b��d�х�b|�N�b�)ĩ^C�dQ�3�
���r��2��K?R�팋6�3�Ռ��=&�|� q�=)�gEQ���+J	�q�a`Uq�5#