XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��C1&�T%�j1O�~oXY�S�*��XZ�7+׭Pt͟cU
�o"c,���3���Ơz��0��E��:�|�Zп�O���^G_Lii�s!���S剀�O�u���ajq��:�IEμ2U(٘9�ߩ�ҔM�5k��&�ǝ,��~
�f��<�0@/�j��
�g�Fl<�U��,->��e�xEPU�"j��"sz���T�����X���qg��P��$�M�H8�8r���1S��J6U�b�+t[�|�
<X���x}t(��sC�!Ox1��+�xT�����u�����
���0��S��F݋JWC/�n�>k�U�i_�PWޅ��S)�h�ݧc|�ˋj$�}�#?Y5i��p$D�ٟT!� ` q�I�̷�d�`j�n �?�A�|)!mѣZ؝�=.���b����-�E�0jrp��0h��GB��{\C���"�h�%c�o��ziv<��5������P��]LqJ�z��Џ!f��/�=C���W�	s�^�:�:%E�z���Rդ�ْ�
i4a�~-V�u
V0�;�Q�(���*�l�2�(��ك�|��6+�{�˱�{F����6��o��x�:
��]�>3��H&x�mc�o)_���v����nV�N��tp��Ϡ���(���	tX��Y�`��"���u: �jEu�ؕ��]k����_Ǝ	��¡k�sYF�| �����z�tF@�>�/!�]"��ǆ�Β��z�y�Qr}rw���ZrhEl ���Vl�XlxVHYEB     400     240��2�	h;x)��(_/sV��AU=��7X�=I�]�u6N+�)�����4�g�E��BC</�������D�%q&�������V�!j̮j�4��jL�;��𦕗F�M|O�o�+ ����? g	WK���)Cv�b|�K`N)1iYe���3��ל'S���p#6n�!���W��.��$	�XK��,J(j��E�@�'S�y��V%�A�t�IE�SF3�ڊ��MM��W�;zǶ{It�>B� fJ�*H�o ��T��+l"u������Wf�@F��F���'�����NӼ�V\t�d͝U���0����8����X�d����d�	2V�j3�3�'���4_��3��C1���xK��4^"_��UC�� ���;ɴ��w�.	{	�5�]��(|!Y9M.e�?s��0�E�G:���Y#����@�S2(�HvM߳X��Е
�`rÔ'U.�A�i�ggq���o�-TVz�[����y��ޛd8�a)0q��﬐�n%�R�eӄ�5CR�;� ����
v���F���k��:��+�̴�MXlxVHYEB     400     210]���]�z�8N��uS�U��
,s��v�'�������=���Lj��[�]~?�,�(@��1b\�x����=Q�vBi��3�<3?�!�F�\���Hr��qA�v
�.;���c����9�i�3Cr�W�]���@���X���P:?���p�$���f�����E\p�jA�Z�o����=�7�M�r��TPG~8����{Nՙui4.�f?�g����}�]$s�3u%����0TT��"h2`Y��$��M>�x3Ϭ��a�]�Ӭ��Nz������ap�ۖj��"2��3t�;�Ў����K�L ���Շ�d��8���6�iN��ٖv����{1ɣ���B7</���w�Ĉ2z�{w Л�R�������u��.:��C@i.0�Ԗݛ���#ZQ���#kfS��4��&N\uo�e�J��V�.9B�����&���1���\��U���)D�]�҅�����s���|&�}yīKh�U�����;�M>���V<H�%9�,25r�hP~XlxVHYEB     400     1f0�>L��P�W����79Z�Y-����YԌdu�+��[�܄�G��Z��E0�I����r����u'9I��g����;"�,��̉QL��Lx��:7���0�f=��o\�+6ݚ�`��<, �k1[��%�w�-]��s>��$�N������.�����2�d��	�2k����׎����-D,2�%7C�\&���d�y���Ά����1�*V��A7�����;{'k&Jbj�@z\��~�A?���B��W��;�\2K�Z�#�i��=aÂ����ݙ=�:Ėc"�7tw�ڎ}EEWp�h�QZB;�����edr`�/�V�	c�W�N�dBz��:�>�lO��eZK��,Iw�Yk��H�RM	O��x��l
J�҄�8z��BP#���l���l�R���#o�cʞ�[1]9����N�bI��&B�Z{����F3�,b��N/�н�?�h9E�eW�}+�ca�ȼ_��Jc��`"���XlxVHYEB     400     1c0�ycO�4���؆�A��u�V2Ԛ���m1�!� -#q�r�kB�e�n���cDI�ԕ���@ų»��ӯ��j�[dF��>'-�*9��:\9�2Z�a�y�Iܚ��r����a��so��G�מ��N\+*�������#��m��9ڸ�� �Oh�0�Bΰ�����!�$����0u!kWޚ��f��k���;Q���_�-��:m4`�uaɶ���lgO��gz,�:&f���VϚ[������[:B��@!����:l�$�N-��j�r�Fd�1�=6��L���"C|�Khc��|����r�|	=_�j_5���a`!vW)ԙggw�P4��:d�[.���v2ȑ��'����[+��@2����X6:����(�D��8#�]>G9�v��x�C/M�cPf���6��xۙ����c� .�G���U�XlxVHYEB     400     200�G���AW�� Jf�s�k����H�#oK��?drb|l��ͼj�q�v��x;�Y�b�;����g�����1E�x��_�uR,����J�j�:��O�[]��(
Q*��s*��{��.�G��_c�,͒���)M}Q)���޲�u\�Cu�=,:[��xZX����}��0�&�:�=@��W���o���uc��Eћ��U��F���.�b'��6Z|UQ`N5��>���� ��:�1��I&=�S�R>v'�}�"��8�1�E4��ll@���	`���� ��Mx�Y���O�F!�r5�"��Ɩ��^OI�n(xo	��z�9Ij��Z3P����b_�7�&����\N�����쥧H�0�"K�>Ue��P%v��|V��F�πR	�a���ۆ�փ.�l�>�Ϩїh^�`監�
�H�վ��aWO��`����n���bX�8$���cS�P��.A-�I�� ��u�b� � ������~ߐ1��AJ=�A�tqXlxVHYEB     400     120��\��n����a��A�>;���jR�]��`��@P�)'r���S�42�qn+������δ�-:���8C^�}��^+�"����kG�,�.B�,U������.�e�@�ռ\̖~O��w/[�x5�䧤q�0m�A�؊�Z�8ہ~)g�t�g��5�V!c3w�-��'fU�Q��SF�)�d�'Z����՜Wn.� u�޵����~�w�\��8��f�᫑�m#�6gN@���N����Yݖ25��H���_3h�6�_��q��!D+*+kՈF�J��	�XlxVHYEB     400     1a0�}��fs����O�X-z��F���[��u�x/�{���
��[��������,��}�k�h����S͛F��^=[�����SHEÆ�N�	�iX�9T�@
�/�'�9�n�Z���d㝩���xs_����_��c�ә:���^�Lp���H;5#Nz���^3�e6P��wS�0�� �V䋮�M�/G`4C��?�f��Թ�R�*GJ������Kj[į霱��L1�3�ӰW"mj�Zd�������-͜��?ľ|aH��= oK
�K�4�F��Q��5qDτ1�?�`p7�[� �`v�ᱍnd"8��Έ	}��jZ�A�1���Rq3�2���b[R{:ϲ\x��N%�K	���j1�5���Y`����� ֮��f�ZD��XlxVHYEB     400     110�5��
�}��S���<O��vB��#?ʅ�� ������Fqα����h�M��^�q��(ȧ����|��Q���6��������q͂Qb��-�L�*�5����dX��wn��߷ׯ������i��Kdp�ߨ%��!������Q��3���N ũ�s>R��%{�6ـl�[�0G�R�q��:�N�Bo�u�$(PmV��3ў%	�"령<���`����XX?Z���p�.�҈J�$�վ����* �P���:��/XlxVHYEB     400      f0Q�^�ޅ���+��1�g8Pʹ�gMexG@�g�R�觉�����ȭ"���X��+�?��DiA�^�!f����X�9���O�T�z���M��^d(���i �G���fa�|���K���Gj��"�ѻ�������
땏Ɔ9�j
s��z���Ϡr��>��O�e��pv����h,q�ƣ6��1h�ny�b>�r5�X��J���U�������/����6ꆇ� ~%ⷌ-XE��XlxVHYEB     400     130�,�<��<bx�+��s6yE��M�d���Us��g!.t��]���e�!H��U38��9��M�ux#���8���\�7�;ŉ�'�bt�>��.^,Z��5^�sv��(a�1if���c@ ތ݄7x���q�L�SaU�lK��[}~���=�;���<��];�~�J-�a���Ǟi��B�L[�xV=���9��M�>Cm��Nf?��\:FZF�w�1N�7������'���1,S��+U�mI5I�ڛWW<K�Ol�u����vJ�>��[;�V8%����\{��p'?'ďXlxVHYEB     400     130�?���n�xH�AS6)=�?,5��h����v�3�RxA�����TO)x���~�JK��!����zq�(�༛��Trѯ�4���,�y^B� m����N��J�q]���d�S�Iw������s�����qˢe���4���Z<;�^a��]7��⿄�%a 6.�ٝ@���jl�� ����[8 ?R�.G���'f�SP@D]�]�F�4Rܸ�$ w�CN�>zJJxKv��G/md�WD�ν=6Uup!Ӧ��J@����hC��W%���>cYG�m?y@;�x'�p(:��H�S�&� ��XlxVHYEB     400     130��rG6fyk�҃�>Q#�Ғ�*&i�mAo/ҭ��AlD�h
��������N��>�0 rd��?�)���F��T?�dBx��A���M�;��%]4�C��g���wJu��ſ�[)At��(o��_���ђѧx	D���L\P�{�I2�UAխ5ݹ\[�M:6��'�	�e?�eMC����y��x� +?�\�n.2������QT�*���E���J�]I���1آ���r��eޡLiy}R���t��d��-�k�YD��ke Sk-sR-]��\����f��r�XlxVHYEB     400     190t�W�]�	�e�wM����{�^��P�&Lr|5u,�f�5��E�z��>���I�Z���+�f���i3�X�����(��������-y��V<��i$Ln������U�n�02eʜ(����N��/x���O�(VR|�n}+ˊ5�F`m!�,�ˑ��Ccx����cS�롲C���f�,�ukZc��Yl
��)<��s%ϭ{��xb�}%?�	E��y>��V*T����KQ��k�'������K�2D���M��]l5�3��>������HE����5{�|0�Ky�%�24#\i:~4Ӆ�w��B��3<!����k ��N������b���(��WȺquG��(�d�)3N�4�dT��� �ϖ6YG���XlxVHYEB     400     110��Q����*����3G �q��-��w��l}o�2h� DJW�
��ͷ��A�$�$����Fq��5A��97�	B.)>]Q{� �^�����[j��I�E��1E%�J".zp=��a;��Ս
�W� ����`�\|�/~���#��ީ���y,R�%�d�Dĩ�S���M�[uB��.�p%-�a���}�2C׳L�v�r\9�F��I!�NB�Ҙ۰B�����ʾN�r�����WÚ��z�2�m�F|���@}l���:uXlxVHYEB     400     1b0t�EMy�W�d� ��湙b�����7�bEG���Z�4�w.��s�1�\i�n���t���<;���4���A_�@
�U�-�fCq�w����MpT���p]��%� �̳�=W�Q.���=�~���)����VI�+J,�IJ��-�
5pj�Pg�n(ڜ*���d_ș1No��A�cD:�O�3X��h���vD�?����@����߮9n��R��أ���C�#��|v�{D�쯙�6�>!��1�O�b.}�jd��% ��l退TX�sI`VA�j�Ob��4#i�O^�:�)@L�4���]�4�C�Kݓ��-���ǭ~F�:I�FZ�����9]�Ve�r��۲��a����N�3l��u�s�ц�e!��3�DjO�xk%�xo|��S��S~U�vq�XlxVHYEB     400     190���"�=�����%'z��K�D�:�r̒1)�g��9�P����?��RyF� 
�*��1A:S\c��[��=w��p�e��`8����}�>�=a}$f[8KM��_�u�.D�L��Uԯ�τY�3r}�7�_Zғ"� Ɣ��֠	3j��[���i�/{P��K�A���>���V��  �`��UEjjRU=m�c�X���;pƜ�=���>��㵚-mrH�4&9���s��FtŪ��`4?�<��#F�&���bF%�+�
��a%f兣<vT�����7 �NA1���_��e.�kr}��%�e`$/Fl�mS�ҏ���3ޘƺT/�7Xb'�Z�
Sҷ��^$�S�O&�
�=��f�~�j�q�w�#A9��O�2O�]
���kO�FK�XlxVHYEB     400     120��
YQ���LCP�C�����d�\vD���m�ae@	4Z�A�e�
��*�f�r����5���"��
��<��3��N�[[Ν��(����x�T���l������zEpK��kJ��f�tq�h�"x��_\6���/l�D�Z�H9�`��!*9��z�JYV<Y�t� ��aB��v}%��i�P�G�����!10`��x擱$�ï3�)i�"M]:�W`�����S��8�}�[��I�	�NN2�� A"�bG0�pH��J���'���ϥ��QXlxVHYEB     400     120�j�yg��v��20���Ɇ�/�������HQ��-X��wJ�6��a7/��+צ?l@	�:����WJ��#�y���~��zlݧ��f��fܫwGۥ1�F7">N	��]�t����)���xx{�E-�@�i/7��(��$�.`��bd� ��M�z���������Ǆ߱2�8pZɿ�@����]{���=ڗ,�%VQ�c�M�4v�5��O/�	a���	O
r�ӥ� 5�d@L���k���S"�����4w+�L�e�V@�.�*P�}����4 XlxVHYEB     400     160�9�|<6j�3�h�|p�i�e��9{n��^����|����#����'\T�0��s��7'�ZO�����S��@ɤ��2���N�9��l�c16������qQ����^#�t��6�3k�cyQ2�Y�iN����k�8���=�jy-��g���;�"��B�?��3].o�P7�!��ג�z�+t�7x�
ц����c��l���Ҁ%�N��
�����,0�4PO�%΀���[�J�C��޽�)�X*����i��c�@����x�,r��[�P�ą��<�C9��7b�"�����&�<��Kn^�a��A�+�IKNc���R!
O���Q�0�di��s��XlxVHYEB     400     150���Q����<>�RΓ@�v��,��k�|��I�P](I7��k�3lr��J@ݶ0�s�5���0���P�ǒ̹�\D���IWW�:q�So�B���e"���n�:�~P���G���8n��w�9ip^���_�`�ܢW���")�!,�9#�q�Ç����D��f�N�/�z�sCI���� 5L]��aLF��h�Нz\nP�dPb,yV���ѯ�Ө�=����ۯ�1���C߅4��˕r����f[H���O�	���^�\�%m�"����ڀ��àT����Y�/S�K�bk�O�mc7�������V��>z�!!��N�^XlxVHYEB     400      e0J�'�p�沬�<�M���r��w;��V�!:��[_�WI��k�E�S\�<;���_CB��_�|���g7��'x��i�Xk������	��"p��ܶM�K@�6}|a� 5ؓ���rdC��s*�c(�Y Q=~�Ӥ��Ἧ�q*H�� �j�0\�W�R�\�7�;�:��0��$p�רw�kij�;f��U�>i�VM�3����XlxVHYEB     400     130��%8��N)��.�f�Zit������N��n� w���T��U�&K�&f��Z���\�Q
}c$��~iG���%��Ca�	�;e��%[���U��4È���d'"�Z2�?�k�	_�����?��:���/�O�ǡ�Q��4�������4u9c�r�k��hٓ_;��OM��EB'���R��܏ �VMX���^�^��
�H��Lj����Ց4T���Pc�~ү)�7K ��q�6������5�ռK/<R�H27H0��ݩ�U���,T1"oH0�[����&!���XlxVHYEB     400     140ʶPݮ���&�������,�t-.i�{2yc��]��־��r' k�䆓�¼��m��<�n�p�8:�H���f`�a��V3k�~�@�6��5?���]�N��M�L\�����I՛���Z�r�:���#(C	��_��7G�?���iU���NFS���G�@=b���iE��-��$��8���>u����Б�]��nÈ�h/RQ��	y�T��%%"P�Ь��
���hD�BG�����;ZG�X9�j1���d��/X���
�vuf���+}�N�h=�x(���m�(��y���K{G�7�tn\�4XlxVHYEB     400     150����k��������n� L��J�L7�5�'�}���7���G␔3?��C��57f�Mi�p�f3m~C�MB.��`�u�E����}�6a�Ŭ�>��ؤ0w�ԛ�E�������{���l�l���&T�AC;�����؂1��j˶�XjW��z�Qyэ��l�Ա�|5�	r��G���w[YC�x�W�L%��3�J@�I�j�_����_o7�9�)j��T�Q	&SǞCّ�V�C":]�pf�l	Z���Z.�T&�c��Y�x�C�#M��{Vl	P�O!ۓ�/��Q��x�X�����c��-p�H�6n,��T�>��XlxVHYEB     400     150K�(�{.�Y� e�g1&ѳ���#�%��j���.7N�zt�y9�w�R�x��Yn���.C�T���CXWu��jޝW氙�����R-���LL3Q|a��.���o^*
�Y�Tx_{���� g�PAu��U�7�n�C�����d�D�)�c)լV�aQ!qJ�p���7^�C��e��x��[֊��7��l0�L��i�ߧh[#!Q&�G-a�@��,i�S/=�` ��n��|��̤'w
W�>?�4wNk�x��U��$B���$jS���~Lx\8~�^=��*jux=T�FG���;��xN�w	v�+i��Х�۱�S\pCs��Zn�'>�XlxVHYEB     400     120��6XƦn=�B�Vn	�gM�����z"�f��{Q�$!��-Jsu`LD��YpM[��j!����Jtor����:��-M-��{��[6��)��&<�t���zd���r2���{���J�UNUw�i.��H؝���x�0��sV�o��@(`�9�F��f5�1� ��i����������1�i�N��_�=��bI8C	O��\g	�\��t�G����Z�;�p�[�#Й�;RXNFR�	<��t�S�F���)�A�'��0I�:(2N�98�7;$�x�k��е75�XlxVHYEB     400     130w�ܣ�Y�$�%��1�7���|�kGSC� ��/A�B��p6Ϭ"	R�zMD�*Hd����
;k�Ͽ�N�qd
�/��
��<��At?SXSJMx�!�ߍ{���Y���ʷ\$��qW�j]�V����|��v_M�7���e�scb�oC�a~C�HN���6��gn��Y)Y���$g~C�Z\���5�T�=�XH?R���'�Z�m2�*-� ��e'���� ����<�����\I,�V���8K���8q�"�Ec��D��B�M�<q<�vr�m�+-��1��D��H�c���$�AZY�XlxVHYEB     400     140�X��8�=��]�a��A	�K�H��
�(�ⅴCġ��W\�t/�W�r�%�^���
ֵ�1��W����!O�ֻ k�s΋�bށ��\��D�\PExE�YV�!W��3�g����/�$�E:ݼ�n1�sk?�/���A�����MD�*}X9�;�WM|j���Q]��D$���+��傽�=̓}�d1����� �]��ѭS����Nƹx�OVҸ�ȯj�z<��S�v�����(������/O�:���<&@�Q��?l�6��U�A�����\�=�.V���'8zViu�{[���^ v ~�XlxVHYEB     400     120WQx?�G��Ч��h�y=���P��C��Bj��~+j�`�q~���Ѿ�Y�����畨(��^l�9r
�=j�r�bQ&n�y,B���D�xS�u)c0����j�#�˾< ��q���@�l�u�g�� �)D_�&���	��Y����K���d�D�m3�Z:$�T����B���3�Y����������5:�-uW���I>L(�C���]�4p���f��d� �$����v~.д���[���i\�˺`l=v�Pz�*A�ܜ��@����XlxVHYEB     400     150��F�C��ʊ����_������&�&4��%jbiџ�$L�3�՛
:����k$QHa�Y!dNO9�6(����a�ŵ��
��B�xO�Jܐ��2H�
����t~�x�M��9� -�gh/ַ���@�ׂ�3⑋��h^�P�^L�DK����žG���)�/�
�[��<D�2bJ�|H�3�W%���-ބG��H���hs��,��X��I�o���a�ʠ�2�x�5K�������c%_��h�anu0|Ѳ�M�&V�m���T}R)3la<�M��! �!�%v�PS0V����+�Bn�h�qB�>��,v{�^���]XlxVHYEB     400     150[��
=h�8nF�þ�&#��o���qh���;��������j�W��"��Y\F[��4;N���@�C��V*)�
Z$�pW�R������Y�w�6ω�<�QrVk;�Ng�2��j��)�@�w��B���U��(ym�X9�K7il�ƍ�wU1��6���
�e.5�Kk���,�ljw�.!����h͏�C~�m<$E��{��G����Vm��'�o37��KV�f���8r�GZA��iX-6������4>���x{Q5���-i�:��7��W ���Ub��Q?��d<}.#�<A��v��
C���I�N$E/����0'|XlxVHYEB     400      c0�@z��{|v2�`v��P]g��g��Ւn6�ߎP�����0{�Lޗ�9��5������cS4�qIw�2U0e��CG�\2�0����(n<|���Q-ҪI����I��`�U���ix�H5��+H�-B����Vw��R�7����ZwS濉� S������|d2��#��(b���J�֨���y_'�ؔXlxVHYEB     400      c0.�9���WPj�s�C�01�B�u�$��7�	����i��r F�w�������ra�&1�^��GCXN�@�;م��L�ט̟���
�
Ζjm#���t[�X�
!����ֱn8?���+$P��߁�5���_���9ך.e�9��{��%�ٜ��r����E����(�2&o�;�T	�XlxVHYEB     400     130���'Oo��UПo7�;o�2�Y-�Q�-���XiŃ�M@@�#k�?�x��qb�tJ)x?���3�H%�|2�$ֵ������[��;m�Ēڂ�'y�"wx��P`��p��jZB��r���ip��T{}��1$#�g�Pkűꕲ��b�ܹj���߬��9�\���g{?�"���/�8Ǌ���~���{7� <�k��JU��-�k�:��tyaІ:�T}'�c�^��lX3x����|׎����\(�;)�-li�?��R�kk��*N\���ޝQ�5��:n񳪐��YXlxVHYEB     400     120�l�Me�x��4k�֤2,0�Ak�5���W��L<Q�Y��\0mس[�u;)k�:O�+�WA���@ԦU���1�ya�7�j�8�KҘ�pH�v����Xхu� �Z�G�e��ݶ?�39b�GQ.����k	�[����$�����'��m�y�fwG�/�m���#�;�BBש,:��kh��S0�k�,��*7��sE�W��u�FE��٪�FS5$0A�����-�٭g� 0�ωlZ/�$*p��6�U��<�6۞���i�[)�3�d��x�6)LҁL$сXlxVHYEB     400     100��ي֦�h�^*�v����Ӿ��������UCT����
��~���#�@��cj��}I�4�����0���|��Ka�Q9+Q�d�7�V��
A$�yf�k���´�����@���bK�G��u���㺽CѮ	�RLxQ�]�J�W����m~xkn<��N�;�T��ZEC��ٲͪ����}���J߿�0<��7`Ϩ\+�v!��9h��,�����&��@y�X���s
�����^���EM�)��숒XlxVHYEB     400     160�����0)�T�q�:d�&�t8 �b�J��V�x�,t��婑X�s��N'+x��LtѢ�.�❋�K
���@O�w�x<k|?qC�PU8�s���@!���b^�5v-]V�||��o�5EV�)�G���_��f��8/�F����M�/�9�z���Q;��&&�m�H�n����Qͭs�����<L?��0a��WK`3��'��������޻˩�����:���u��{��j�#'���"^����s����;�ق���O��,�s���	>�=�y	8�\|�Y��@�ҝ�6/(2��V����=�|�7`׾�'���޻Y�6I�0�PXlxVHYEB     400     1c0�󂲝�)|���= h7#������rQIe&u���@r�T�F���_�jq��A�J��R�ž�TG���L��}���#w���>�g�k��4Ui�vR@���u`��x��������RY̖���K�FF;�TD;��b��f�)&��� �w1����$����`�[��ѢS�i�Eİ�����R�A��"�h�WVd�'��Xjϯ�c�&�J8�����C���bB3��.x�bF7���=K��,�vD?�j�+�4��@TG"�����g���໖���u�i7�n��FP|E�Aԟ20'�"/Jr� {8�NhT.Q��	+f�}��f�>\�1T�6�%�/�?��V���FkfI��GQ����y����J�<�ە��4.&�� ����>���F`�(�LZbum�iyb��T���G����� �]~x\�0�c�WߙZI�bl�XlxVHYEB     400     1d0*S�ߴ��]���Ժ"�&q�D5��b �'�S3׹ 0
Z��Z�O69]k�����U�$k.-�1AZ�0����4�T���`T��` �Y���2��)�ķD�kJI�L}�Hx�2��P^�b,Z��Xݢk "�q���S�֩&�n�-�Ae����?^m���j�emw������;˓��۽s_�����
=�4�n��vO��ПT$��p�2�'���$�B���0������E>�9��%7�S&�aX�7p.�B	�v�S��@O����������wh��$^���"��l��a�%�k)�ă�1������f0�B�CMk��t�k������<r�͢%���JmI����eoG}�իo�]%4p�4�A��5�ҪT4'ܾ�,K��Rܗ}��9�Ɲ�������X��0� ���w9�J�cb"ôb�ʠ	*[XlxVHYEB     400     1b0��$Ư�IG�^t�b���$�xL@@�����T�8ҭ
Y�3KZCy���������X8
����h��'%�B����1݇%i�XP���F�fk� �^Б71<Tj��QG�����'
LU|fZ���s����3�y�nN?ڤ�^��\L+�j�3�k�F؛ZVYDp���E�g=V ���	��2J���E��3B��
+�Qv�[��c�7����6p���Qd:=��nNs��4<�*�Mh�s��y�Xa��5-�9�čO�6��)-���&����Й������u;2�o]=��1�?��/�ϟe(=&�3=�++p��[�g��vֆ?���������ˎ6}/�`Cg�|�zh�gaX���3\�`#���Ejo/l��R�gxy�G^�Yv�'�j�_F�Fego��ч��<�ؾP|/X��XlxVHYEB     400     1a0�#�EgxT���-sΣ�g)H�!v�Av�a��3�?�א]��f���A�$V7�?;B��5���Xh}oo�Z�)�S�J��9�Z̳o7=p��!�����s8ё*�/��Em-2���&���uF�7�{��)q�::��ycp��gj~.������Z$��o?�\^V�/�뎺��?7:v|�Q�g�H~��?�?���!<��vL��� ��{m`�B�t���d�	óy9h���K=$�{=�U-}�����Jb`�&.�A(��8f���j6���1�V���~��6������l��!bA�b� I?����~
{��t��x��=)�+"���J玘���nw��薾�Ѱ�l'����A��J�����1�Gh���]���
Y���^�HN��Gq�+��XlxVHYEB     400     160���R'!�Yݰ��T[��5�����B=�3l�J]0Rm*�,��`�ܼ��)�@dB�L|+�2�yťGp�/2�w[�x�<��^�vW<{�hc���rZ�ܴJ<��V���7�Xi����bq��=E��>ˍ��K��ҶS#b�L]��j3��S'f���&F�����$A��fr��x���w��JQd*$�$*�hqb��v�[(�x�{�g��݌W��A�Cy�\Gb���g��4N�-Z6_GW�AP�v]���L���x� r�y��m�v�K!�~<��m(-�&�;�c~h��	����T��X$a���BO���^k׌�L-A5���t�r4XlxVHYEB     400     160r��P@����������_
�a�pЧ6��!aZ8��_��rT,�q�h�o��q�4<�	,�@#���|��#��w�/"팁��,_����� :������K!#l�^h���Y�A��0 T�����XCo}�T���hTsn����
�(^q�Q`����M]��XO����M��5���|Jj�?�%�9Ǘ�R[�?8Ju�G���xd��.s��]`38�h�
wJNhG���K՚��?�:�7ؿ{�Bvs��\�� ��#��|o�m�ϓ����>Y����o�i��E��Q�Ϝ���}%藜ɻ*�B)\Ƹ��YT�K�if�vĖ]SB�~<dwmed�pQvXlxVHYEB     400     180WB����㒭fGc�G��Dw�m�ez�	#}l��fH��� �,����%�q�z��t�(���"��0����"i�M֟(�gj:�?�Ѳ�\;�bq7JL>�X_J�J�g�ő���7����?~�H��aR�ꊩ�t��+>e��έ�w���7��i�d�uF�m_g>����1���
=&1��r핻��Ĉ]�_���%�wv,!�3�z��,p����
���Tһ?���.i~��@E6�������0�uU��5�[S���[9�����C��T�5
�E��.�Ϗ��F����:�b����6S3|y��w�cR�Y]I��@�!�Sf��ev�����j`Q�i�Z�v�:��.F��E$�J�:���C7 �W��@�[~XlxVHYEB     2ed     130?f�3tu,P�|Hm���G3JØ� N\��}��&pL0<�;y��{�JI��k�LO�ߊm8�h���6�;S� �(�>�������Kta�H��9��{P��9ޚ�A�E�Vt�4��)�~�gH�{�a��WO�m#�Wў/�K-���o����&����^b
�Oˀ��ڇ���A��j�>�sĎm��L�a�ѣ;y�s]9��JK��x^�$A���=$<��a)��-�v.j�Vg�Y#S��`���E>6Ϥ�Ε���&Hޡ��G��������f�h����[T�,���-��.�