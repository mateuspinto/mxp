`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 100176)
`protect data_block
1iWuifXuyVGIP6VgMqj/Gnx0WXeSB0EoLwv9mZ2AgIO+PvPczfCMVQVA621iPjzAFaX4jkHR0KsJ
uaAk14dJJDvnsJsZkOlKgMfan5jcOTXY/o3bXM4DpYwYz5n7AIZIQPaaiYGUeGQ2TlyE0ZuK52bZ
wwAqP4liBtjgE7U+i3H8WjF/THQtJyzs+ger3Xo8Er7NHEIZCD89iZZkfCdwBi0ewsb+R2J6bmVm
ABmLQa4YSZJgEvdyV0cWxblcw1Sm4+NPVrmjQn4CbVqP3ku9x4aoFv++Xb+w2RqQWIBZMUY/cJxc
xftz6dEcgm3SxBwynJrTwR/LQo2z2bRo1XImwUCgDYGaxOBqKWs3uH5dH8dfv997lAgMOOngUuSt
pJe5ZPW/vj4788fPBY1hyohXaI4QizYCqW/FXDsOU5lTEFqA1VYUYjPW4Unewszk4KTMJADsVB2K
PGDfLxfRDvD1kZezXdhVq1PvIwQtqhwR155m4rD53zfG6VOmOJ4wdnaYXyU5SdKWn3xOrqDY33Ze
4sDe28mQOK+B3px03cZwmHcpi7SYlGTcTV28IuS0kj8yqpDdBHGgmUs6oH1BwizEWj5Pfw/Qnuq7
AfBQXbiAcsT9K2U/SANThOKlX70NpNhw44e5kiRfXOtzuJ2nI7UDGSQVSaxl+dRy6YIK5tO6uZyU
1hGYV/WfhMAxYP+APBDt1xdiTYXu7BMCOSrATIBq2hd1YR2QnD2k6I24JIGCS8q2mHzXEoL1GMhD
fjJZerzFE10cnLAcm68/Rb9SXHGN9gmcqgRx9Q3V8/k9fSZhwGahMpHDTtw0E3M2SL5rMvAkVzB+
cL47DDqVMwXZ8Yx6p8XEU6n30fVLshDy3R+8EF0Y4NqnKBRzfAC3CwCW0AM/jMRk7vTWRBqOb5F4
Vq4rTG4RzaeSU6tQrOWT2CmOuShGIBQc3dfc8rSVwLlP3JwcqgmyQYLnJ4sB7mXl3Y9Rg2VSeiJW
xw5ahbwToiVEtvYptpbTgHr747byzVla25X5yl5Ghc32OttERNvHsb9mSMc1M7i9BCUEskzULisb
vW6w2lh3ReN37BzLuWJkdqzFdFFCfHwm3ElcUGyiKbYdcQlt7WuHk25NXoxOwPUjdswMnC98jXfb
LdoE3F32XQoX8tUi1gRoOfMdWaKb66MQKozfXvjEnJ14l+gyFpGtqU+7rMqME7poLfSMrKenil+Q
G7rfT/czcEQybWD7lJZ+B+CG1PuQSidtb07hhaM5TTgdvAwfjcZEgONA8TdWb2EaGhLNrtiZtXad
6b6sqvxMdx16y/iHy0TDO/mNjhn2z+iMF+UlaLi7BCr4aVydNNeW35EdMHeV0Lbytp4e3CYb2SUe
lWy7H5hau3ZifLH8dz1ooyArkAEELvYZSUEdSSw+ZBXqIuZOEl1PHfYFbRVT68o4sJqZhKBPctDf
wqN5RcD2GkSQggDvh7bFqFZi91obi8lshLrgQa7U4Taf3Y6xK/iL/yXnvHrPqLmdi+nr2ztcD28x
MQJM/7TE61g123dmlw0F5ICamy9qz+8KHl68XIoWDXq0ZP2u/gGvWK8u52ZtCV6PFnGCFNF+0ZYh
m+LCRlINRIJHT6D1t6CC/ixN2qaDmvMjkw5khes6rqxFDgffN2bapdIv22aQ7twO8Lz2LVV8gAQh
gbIZYTQTDHBhFuFa9BcxSCWcWB1CkhilQqMXsgFQ2tsw5pYnFJ/BZmGoerOXf5U5U0zdQqTUg6Xu
M4ImAi0mYm1X+TOcYU8ziyEoHtjRCHlQg1BrFo5n4kIHfhpR7VtxNpPEHo0h1INXgfZoL6ZNTrPc
0A7jfYf8KdUwDJgTcxrKEwjOLPyZ5Fh65jpHPI4y34WhCBpWGW64p6J82cCMrFLEBTeAQSes6LLe
g67ga+8TNh+8IS4BorW29o/KRzmEWUMH7W6/vyeHXebaGrzCzikulQU0ktdZnaLSM3lX1zFkfyr2
/BETfeuQ3Hu6IZspZxa2odcU2Nymnc2gOW1BAgac8n3i9YcXMpfeG8cB+Sya3m7WYSDfNC3yyMjw
cKyByh4mHIdO0gHdjq4dtng7F4zIEbecFKn7MrM4Nd2K0MKlhm6hVdV86xRa0njWHpbtZfNx/eK+
fqDOl0hTws9RzH8NHSXwV4JtLhoWkh9pmbCoCMwpqIcxCRUIaT3cnYz6aysw8/d/sQh0HXhHC4mB
Dd11wBYzpTMM8Xmvx5OaoGkEa/mA3DEh4qLoSVc2to/Eeupnj+7+kNL90tNuDjczvm4Kfm1R2pr+
9pMbrK6RzBZYl/03cDjg5Qt/YnR8ckiNxz4OCoSsVCYcP1VyT/9xnYGx7NcvoKDpoVM9Pg2bmWdb
+lKuwIpicrlpqd9rHc+BQ+7X15v6wqFNvr0QSy1PCfzWoXJo+CLsLu2GaCc/RngFcCo2gga3CSNK
px2PPoSEid8IFcHOqICcaq9B5xl/KsZNx0R1zIJPhUj8QS1/eX1cKYMDSkHm31YacaOsdzEMjJqd
5rOUanQm87vunqkuNaG7LxCdukLU79jrT9bi5vRtcPw/+iW8RqGbMC4MSdYSDgVWmA+G81HVUuE5
kL4IW65yxQ+lcssOV+QJFGxbCRpSUdhFEX+AzibBSxK55mK4wN9FtIZcP58AAZStkyWUJ1dIgIFz
4urTheCZEqqK+rSa6kvWjckpY5ja0QZX0TCb8Z4aMd84VResa951Q0dgcru0G2mkBXa+ciPpYEwO
LqsXSe2v/LdfUBXfC2ITjBPgZfv9iXqFLeyTMBZzw1eOyGW34kA1apFCYI5S/OnAYnRFR1WRs1ei
ySjsUEbLyiq8kogUbVmk0rlaFmLAPMTUYyjXcSGyFwLKVxUTq3FWToNfpB8AQ4lxdhmnX3ZA5nmi
SHq0cA4XxOFVSZX4k4QjU1Yj7ArJlKvW9339fItwK9kjYvT9f84z5EMr+AzUxMR4A9eGGdirTaL/
lj5EKo7AWp1hcM4Rs4mOSvGbL4qAv3HhI1IIkYDC+SMgoKrdwZ5X1cQUsCNmIDuqXU0PSi0Z2jiY
oDio63Nv4IFPk+MiXiBgHAoMv0kIulJXdSl6rYL3MybZ5gkrroC7dZVefH211JJdD7Ab7IyMpGHA
oEivNGpjzroeY+wTXZM/WW1ZM7Uw+LNUCfSxJpAXdL1CJMbtVxLLuemGCQrRx89X5cb1BnoilaJu
vOt8YAwPtSsLvvVwAzwldmdnE3+tpMTlmlvzjKph0jzq2W+4dgJPPCsQuKVefVGg3nkaPKZDYZhp
lQ3ZcDLYLYFGpFOo2k/XtxnxjiO/lfny26OK3QAF3aZCSxz2+kPAQN8fQStzQuHch6PDGyrigyuX
Xsg89NUtdg6imnKpvOMbKx+52a/nWOKLQS7S5iNXWhruZ15TBJpLqqDBAw8PlkPjGINEmLIwdZ07
L+JRyjQZDAH8Xw//JOFkjY92M8pzZ7NfJAX6lZLFUTkfy65UgSKNBF4KMOWGG/TFp8N6sY1j3XGb
jS2258uaQNbFdvOch8abBZPOW0RbC7PGHgDPoAAaHmXcXaRjr2OH0xV1yXwSSBT0yN/SSnN0Slwy
V+UXYvd/BNwa1P1Rqmi60p9voC48HBw/VSiQmO3wmB5BtHh7PBtprPEIDj+JLnCJv7HmN+wsX3yn
jsvrtQm4xdvtC5R+NjFyheEPxGqEG4U3ZlZ7ekQEz6SBYVE+3jLY4bRt5gztH0pVpU5Dz0iHne2d
0IaQoQoo4p/v7mVGL/09NuWBKntBDbOt3Wg/js65kEFS6e9f2MxL8M78gJ0WeArl1EtdNMKEFBPT
LXzcTeH/1ZjmRviDl3bRXKA72x9GFTPLrk+Bm5Zk+zmwCTjIYXXt8QeKzDxz9+eKu3LZP02QPGbs
RJSS8siGcoNb+GQ5rif2DBSGqB/xcnGZkIuH1tryc28f+uJv09dFtH9RYGgGCR08tRseSlDMUrm2
clYh2Tn3eUN1BqtJ1efJT9Jtfzs8R3ZyLE8O0jwix26DyUBZu0xqnBmo8k+k07B3BILd50OsWcmA
y/8T3qtGT4lD8RTRfsS7LTGkaqHK9wbcmOIPO3hUm5fokYV09TxTHKkkGCw5A7DysGG4rGKGwoYM
14zyksiNbbFeJIvMktuqKZyvMtVrJ6UHFYLd3z4VUeObtDGumK5XBE7hq6wAo+HzNyI0oiCUUlry
dILVRdBurKXrtgfjmiPQDpIC7Y8PHW1UM4JFisASGi1H6HnxR2Or4RuC8x/zLmxUAsL/F58VZYFV
XRvnSqDVqmaaSrIicKnEONaZ7usWx0AG/6ojwj4nKqtGl5pnkXf6BZ3MjKq/PBg83OwOGtHXbtZc
BrG9CIERKj4cmqx9mfQ1VmGIKUj5S4I6q5cQ6hqvTIJJf4zv+Q/Y/0Rrjq0uviY4kuIBi7zxfGqh
rvlWNrJYdtQ+h+WuCEsIapK9jfts9xOg5Jp1NVjNMI8VhpEcL0lfb+pG5fD6WViRtGXpLzF3PquU
gQG35Saa/cIAjkhLb8CWgpJtlkcDz2pq+/yaWdAU8a0gwHYJJElGCLp7wchy4wSYFXgGNAYvwaSt
EZSwbXdxs4zrNfmDwap0UDiMWfif+b7rCXJpNjAfByRQgGtc2osZ5CGjHazCT8LsW/IGmTma0jVT
OPzDS3etmsv4lZbq3MRL1QicvRU5LIRV4T0A6UyM7PiPxMU7HToFf1TqDIJu42vX/fNGliqYk9pD
kLMH+emZRN9NTFv9qo8ukrLDOTzrtuQ1AoiUg8slYWNOvZhfobBxfsk2XiJoub6UHSrk2eG8aZ5o
uT/6YD9DT5cclbzIBbsEKajB/QEVdI3B6XIpuHjwd6NVimiKwHM0Z3g6R2MH6BTyENRWEbnJ4ice
o0XE2PcpX9oOc2lxYDpaC/GoyJpBafL4fg/GoK+owHt6g06rkqS4WHCl1xMLJ9P6d9zemjdPZLSr
mmkrmafCB3bjxYZN6UtYVySW45UVSINVHG9NtgbhXZc7SAnb6cfSWDtFUNdU4uaX0yztl3i6ErsI
es8BhLB1pL2tWvmGCgtxfXb6hU2oXMHIv+cbrdxhsOS2HFEZ88HY5S9Gz5BqkAMCunen77J/H9eX
lTV7em7kgTwx0cMdevwOxRoydwkrUj+JsN9zqMt8silD57/OFMasjOWX1LI1QBWk62KZ4UDiBQLM
obRof27mYm8WId1mUTPEkVKmMJMqw2GQ8UIPEeBj0b9WDdGIzUriY7rq8ByCvjQYRXn+2AisQ3bw
9f4zjRLxCLq+OI2oyf6QQC21HP9vBKV3R2v+JC/GgZz1Dra1Ddzky0Pp/W2NoWC7bHw9D7vb+2Ic
pyF6Phm6XbcCUFcxB8NC0AIF6VgiawYcnq8n8I0RCC1DXWtMV5LOff1qqf+2MsH1ezKHy6l8h6It
BKje9DTUz2apDXFUCPnCMxrpszN6XHYP/kH5OWEr6UNjOr7tuHsv/2xkPy0085pIgrng7mjrZqJG
RfciG98/8TC7YtXdZuwYhCZBij3/wA99bamRplHMKwMmrs/6gf5eXN+oA3Wn/6zIaz8BoDShCe2p
uYes+aTaqXr6GIyc/BFXUuMSodssI9bFkdezYCF4N97h1VBSM83uBolubdWiNHLEcZloF0t7I07+
M+FuLRp3kDSZ3AD0cFMXgKg7oJ5pBigfQ+XZrVNjTEqACSD26K5+hG8VPKBwAuBGHaFHJTiolDs1
M9LiSlWRHENtt7AocGwyExzl7F9zwXRKLzmZACazdYtSqCEOwiNdG98Zh+DrvQdriTcU08X4uV1B
Yj5TY8KhulA3ZxlMHK7lw65rPT0djhUGvCTGTU+U6X+CC8dtCCXNKko6G81yg8bMfumEvo1LcCpj
TTfRZGQ3NVRU4VshgqzspX5hqVSR1mNvEZaTt/NSVlqyti+wwi7qBCankEsQ07zCsLX1Wo/rBCfu
71spBCUvwzln+3LuIeNTx8ygMp+LhvH2v7Q4tFN1byKiWYEzosY4DYzPg686JUq0gdyzy634nGtj
6rNHsVfhongLidpQLzPyl92XpO14Z3xlEBcpx6KI0Cmh1mRSdb27yP7uTkj/rttrXHlL97R8TocT
cxHxGW0cMyPGVS1CA8VPc9CZKm7I8iGqdy2XQztGqc4hSJzmoO7T4lChlzSyFz0RJE0IUCajMif3
H4YDd+BSllc3hwOeiVPlQ1eIAtxtabkagymK/p51FFPJb6qx5JKN0JMoFZbord6pNweuIBRIW5PO
RtTtblfo1Mu30ASip65oz1udsGsl3OFnfjK86C6V+MlU6xa5HSF0FnYNPGX78rv/wQjUzi/lIqxA
3zdeX9qCa4NRioAqy7lMu5DSBx5YebzQGiEzUurvc45dT7H23bnGPMDvStmI09nBnXuWs236Ckx6
46Evf2Ctz72s1CvOkl83bEAX8UGAf3Bn0tyObZvfRbj3QbEouOEAa+zdm+2Dy0rdTcTmRnIsKCPx
pUheM+WCbtzini4md+25Cz5198qHOyChWLReavGQCVRUk6ltVOkUcp5Ty8kM6Gkl6ew3MR2eBDZk
yoHr/WdaBjOkMeQiKL7HOfOIsPNRTQcszMdII9AyGh5p71CpaxSNj0QwW6+eJcwCZBidekWBf+qI
//lh14PDqpbUoilI5wI6cySD1VPemo/rrySB3J3CbTPGv7zM6+p0YG4DCrnRluaOhNugxkE/NC0k
nVA0xK3XLEmZTRPOUdvRMmg6JZRlcS4fvH2hO6ljTFKWC+U1K5GWx7l5JK1VYOeK6VGTWoVL11ax
W3KxrqaK8m2tC1YX+8JVbYOZ7/XA8d9wpdEcMl6wvlnGzwJqitJ/xNQEuPy2ciiZkY7kdqTLN2K9
1expMmkkGf1I8F2fQH6xIRVce+xkGPC7qizBjOlGnoA73SNGQZ4jSIhQzprEt4+NMjWd+Lc8BEMV
6Es+Qylz6/SOp/l24Ifr7+OVR81je0+CPrjZgOKhvzssXEBRAoGj09JB/k5qiXkKkKA4vieuW/2w
p3NoNjMmevuqU7WaGZW1A5BHcxKPOr5Mm6oIzVMLnH9uvczS2GERuatAbfeGO41dlM1StNQDOlJa
MZbZX6F+44ase/BnqwcGvTSsQCMlJlcp5/zDtyBRK3hn1yWKk+i0GwLLrfNSCMwMhZ5JCG0oERM4
KcaM+AeB5fjiZzGNFzb+Xm6hbUNJAIMN+H8iH56s5AFuQHg0liNWtb6LXIWPx70wAKTl7HpGCmqc
mRspDzTih4V9ln2h3gwaVwzNAwzMe39kPCYOg7lvJDQPf56tjl+2GoAXRwb/dHFjtIJp41ALzQOO
EYGRt+Hg6p6H4mRAWeIa4GtsVph0N15eiKDEL328UJm4ri8VBao4Ul4CA0m31fI2nVrHw+blO3h2
LyG3PtDO21qrifZwVtIdoKWzqWOEy6czG9QEl4Ii5+sQChMKkiAZ/4M4XIYC62oI2WKMD4JV/T6X
LAFBFolxTEMT28wRwWfFR5U7teWDXNc9svRychEm0tyJp8ZvZpkKM2oTAUCC/HCl4KDL5xh+ZqNQ
kwsAyw81mFMzPHuga6eT6Lzz55AfuniVJLXXH7qDC3AnbDdGsCupbPQKAsVXE4cKRdWsIsz/lpFA
soIgHxQopZTVG+ouWfHbBq+pAjISswiSK/FmMO5lBf55fKKRX6IAMT4eBGW7v7xRlH43NPDQEXqO
5K0IRD5SFqxzGCaOJxHToTcQ5FASIFAlWBmCzCrB5uM4WLGm/nQnpb4YV0vVbDfyDzNUa7Or1yGO
haYzeatv2Kk2RaK2iPdnvFEFtGMMpalFIOppECRTC9uiY5q5dMweL45A5oF+87jB3wmWtz2BHFBx
hNBg9SlRVn0vdTJNXFoi5F6F9VU3gyC9x5XIXon9ytoruX22bhlmz25+jC4siYN8tL7x7V8eiHy8
uwm10a/Q7TVfjqfiEihmwaoo2NzikqEyoPjdHdwGGhGqQa7JRClqk/YCDUh1fFp36HZDN8ZSJ5kT
Xnluoylnwv5n0Og+Xkh7kTii4NEneIqk3YCNyijRAxSW23twA8n1Efv/drROHcCtRN0gQcoCXR+L
77UiwYoQVXa+AR2WYQPm8Sq+c0+cdfojBcKmWtkx/ixnndawWxPycaCSFuLDII1VYizvZjABJZRP
D50vkps9WGvz5lW2tiiBc+avxz+z5iKPrbehz54JIgS9kcPNDCudb9NIVJheC2gadGBr8BwCwVVG
SpolHWof36Co9qjaESQaQb0ORqHm2PyCvTLEfRt2GLJKJ6NarXUDIiVkYqOoQLnZsNc3zGLmHFpo
4SUOy8K/o9bmn7YW7CjwC4RtGKNZQOMlLG9yIVP3PTxSw7z/oQKhqQTtdDVm5RoZk0L2VzWbO2ZD
QLiVw1KL1Z1jmKplhTzcMLoHlW6qujnCVl1OhNwtedOhUqFz4t4ERcD5zJMuwrjD5yVB+Yb561Am
R8cPFXHpVrmwgLhOcukAjE4eg/fWfDjJMS6dchMjqgKstf23TkMURkpkQA+0SoWPZ5WqVSs1PAnY
SWDge280/P9FhoPBjvcgu4G5WF5p+YIp48AYJ0tH2CKGuXDmnVXNaejLLuHtTraBdDXOiTbXNfYV
NksK8T5cKUXLmyjjwnPWqHCTjkLvewbQU553Snd0vfISzem/GTR8PINjdYy8e7T0YL0OkTCPHbtO
ID7F3dC23gzcxrBt2iu62UclSVKFJ0jXbR5GnsJJaW9mXUqOX7pg9aL/MD/zWx2rrHPzCKv4dtVi
G6vaBReqirf6Su+UsBQBH/PYtacOaVBVE/TtIz7n8NdDjRPGaxtR8JKZXhAcmEwcx7ZAtZWSXrMd
kmVWSkc4H1Ot/NLVDq8NprgDBNcOHIa4QC6npf8J6Q9cCHhnivVM2tKrqLQ3b4SI5GKAks3o/Ew0
uixUtY8l7Ly8h+DVPRyn+ThKuVFTKgy3h8C7/tGcpexMw0CS7rqfSqC9viDOLRKAdS/s2Z3SSmdB
PP7KGCXmE3vBeBSgzSPiIuMgTUWVpzmR41BLPfqJHOUYNyumjB50bXAdYxyjGhUqrGHnI39/3xxo
QMbrSSN+AHk/iPMRRe3p/cPuZX/h8nNLa08PpuD4jal9dnR6okSc/l8LwR8fKt6BzPmApdhAIqwj
WjzMN5amVzP7H71BQhKkN+kiYcpDsRe/G8xHhtzQObgtUZpR/Il468dJGpkLG1IEfklMh//TDygb
us2TUbzG+j6XiiHV9CsGA67DhuWZspEDrmcsXMDQgVzbm5/rT+zhIbOvPxZpeFqolGr3+Mn2wceE
8ReThFtF0HwZe7V3ymclgc/q0XSoK/qRzI+outdonLM0YtnjuQCu6Qs8vcUQLvwSOyr/bjVUlGUz
B1KweATfidhdgM1xOHQcPldaO4lyFzDUvmhgRBh7abntvzxmlKxAPIIgfl35CJK3MqDlrgPsmyjK
nBRWQfG9BCgVYvENsadgWgGXMf0atCqy5SAQai+2i8fmR8BFPrvZ+orIr2DBQS0TpGDI4SMmk0Dl
Io8g2sRFO6JGjXYR2GylL+ZJiZ3MUVlqmH+wV86qtnxLebevSRXrSIsMX4qhf4Gh2pR2EkhUY27q
4QIj3thQe+iLwI+vSLAaDm6kM0lO9CKgk3p/D57LVj9XapHCRfNUSuaE5eU5ZuU3f7+pJqhKvMhx
6NFCp0uN73St4XDYBGAv2fG8G5iYAFwcu6SykK9faJiU5DyeWV2+35tsviCG6h8Amvtm47DIvi/X
ADkPWSvb9wtXy4YhOoBnL7N83jjnLpwlKO6w18mSNWaO0eyXA2kRnZ33VJvozaLi+Z8JHF3+OS6M
a2zesomScR5UZoEwNVcvNvBUKisgfoBQk4e2Bn1RkWFXR8DEUhwAiRLJmRMDY7lka3XoCg8xg4cG
a2yd1H6L8ST2GnxEzvRG9gTR/V9KNFv2G5GVvS5ZzE0MVbXgo6dUm1S93M029OexzSaDxLiQFtlL
A1l7BiIbSRPRE9Yt66uiDnAzG8wuRPjitXrVfA0DklGSeHfiQHNq4F9BHjcVdeDBA2oufvlG2q/4
HiN082t6wz+FZ3N1JggVX7lv4hJXTUtJUVpEM+pnil9QYduCP55EPg4NJu2sSS510q22oj6/hLYN
NeixyeNtWn7AJlda8YzrvfXsEVsGQ0GarnaCJUCwpr02TJR88SNQiYsgjmK6MJ+5T3lvQyUcjYbe
Z8hjH3mG7AEwAw0C2k0DOuZzKwKOJP/7kI+bHFhCyMBiDPypgpd3hWKlhy2618xsIr0+sRC7Gj2t
IgMNmncBK03djgyDWDO/Ug+9zmHwddjkZu05NFLtgAMqkpcasSPyeB+06Mj8KgbHu96+C15/j7jo
mt15NykJ8uByAqASk/r5jabzyQ3pLCULqQ9h99sv0lpUVOGcsAFwh6v2/6cS7B7jP1RawN+OmC1c
+Tu3ePXgSiuzMc/GPx8UQIEzqgK0p7j1zbwhR8IiR3fXmGsPLP0RewRTbzY2urpRdgPWMBHx4BzP
8RtruQ7e+DAR7D6FMWEM/AwCXOEG4b9iFf+qKnbS1XTkfnJ+iMKPJWk3a1an0MK4D6vlpSFMwJ/j
ng6TjUPP+Q1+Q4AXW4H+qLYLYym9RLIZ1zJCjCkvJs90eXmlefBr4+dxYUTzIrc2Ms1baWjlK2T0
LPSPglq0IBUDAeDo7moJb+bSLQq2MWcMXa7Qr5LsndQpoJ4jF7wLtOL7FeR1PeI7JfxdIr/4Kv1i
BhYkm2DTY945WvFbcQ/Oi+cwmYI3HFJmygXYpCJojNYWlszrHQSRvsjrQci9LDpjtr4GISUbbRcu
SwX7R8UGXhG80LaVEDJS+Sc1iBSI5TrwoWfa3s4T8JAxpZFi4351jMrP40hTbopRfa8yB+jEDlOT
z4fghFlEpnNrayalwL6icQC5t8mpKGihh6Qhokupqw78Ihm1NXPv2SLw16w2lLUtBy9gxWMrh2lt
KZ33TThksDkNbP9jTjkrTMwXhQqxhDXeieIryEB85UQPv7T5Dsjm3lOpyJgxmpoVvlQl9TSe4K7C
7j5VKGNlxP+g7CQVVDdaOpEz7WvucCkKvmncC4YsElmbNMsPVsJHRWe9HLCeNkVyKh7O0pfcnScd
I6k5laqY9oy3OSIElveA7lvWuKziGctc3a3KkGVotgqoiYvsVT7o+gKMuBsgN+zxlmY2qf6EbIhK
QF5pzIkP79miVsRUDIJ77vggfBEWLc2rlSaB+h1rFvHHDOuoj6EELKYwFXG1n/wERrJnJIOGxGlw
dGmhiVOE1zxj7tLEdPbRX/+K1S1dhUk4jusjfZm0zEqrQ73mwn3RVTlL/AizMsNY9LbyRa0N2FSZ
g32ogw0h0tq1h3ybMQUSQLnZRhCK8tViCBMajx89LMjTQksDogkjC9gLKtD/0VoC1+M3LX7gZlkm
MwT/I5Php6hzxfAnxrYotfhHofLSXvLhA1RPoA3YdISG0BpKkH1HWdvZbpsAgWjquLdk3g/3mFRU
Xe7dpE4o4vVmoxlWvK1jR31iJ/FWfvAGdXk1qJMkRTdsFHtQFwtoM63gPhEoIbIy4WuUKuA+Fzkc
8qX5+P3plJwM3HBk3kbgxvWVAcbh3FDzzUPme6PV9nODeWafHWAc1zcSQwi8lQ+GBCp059/hnlMW
Uimjr9T318SUVkSYX43qONCR9r3I+Zc7urriATa2cASYFJg0SI33D6CKWYmc/TU3T8y/LgpkFdTN
y69fKc2u4kG3LdrskycACNQ/uBNO67sttUHS3BjtSD/qJk/CPVCsohtC6ju/SiuWHDM/TAyqYKIE
/xhKghokz1aX6zkuGU+9V/fwG72SLzKt6xMzLodeCuFYDrNrlLHaFp/23uKn0jE1nmbnX6SDqa5u
Y5E3jrnc70JLp8zQ74yGyHKU+re/Qx44ET+TBGzB5hbTSYRK/IgA5yljrG2gQdHIWjdyruB9OloI
794gqym0O+7A8HUwnhUxF5rK3B3+CxE62fIGWzVbIHcSM5p95oO68r5S0UZH6Nv+xVCvGExq/t3s
eDYJwkPl4QBYTSOiAw2xuNHsjG2xGKEdLEH5rbQa2jWMFzfREU1HRS6jw9nzEzA/3+jlZhTwBDSv
BbZ2h5pkH6EeWpOFbXbcu+o7I8G9yEoVmV/dyz1nssDCyDF+mO1wEmT52QLkyXxxsR6qz/sVE4mz
N0g07qyvlGPnjVF6Pz8m0X1hbu8GZz3eMRBfKp4X3DQ2QoBpZyYH4MhAAiSILXEiJueD1OaOzuo8
ANza5FINRy4895u0MBcn+kKN+D5hhwQQ1D486d9ZmXWcbTQC33Mp776IKO0XMiE8mEKxmYaHau5p
eGhiOD9mu8xgepd71dgH7MFMh8NS84r67ihEXkt06bDF1JjVkKOMNVqpbYzz8gJdRSTBoXvlN1YE
h8lLx3nPhrrUcV/fZOY2FOI04YfdMq5tt5SDTU51rh/jNiX471vJNnq1nnuXCzkDj29NF7K7bQ3y
h16FE2EpTH0KziU0+R2WSo9EjZ9B3hya7FzmxNtrUSpZ5gWxpoq8sbeZq+YUv81mGKiTvNDyg3Yt
rFAS6Bn/PCAKmMuBCJJ5saczDWwQdcTfe7gkbLh8BptUlV8pBYVTqKQI8exTVB8OAkXnjaKWuzoo
HU7VBDw7Dwv/jMrH6fZYxs1R2EQ9pU8PNYx5Np1tbWMupOLe7IOA0ZDjpH4ZpHh8WP9HHRtMBUE5
pGQjdu76ykTXQacoI4X2WxaITBhTLBQJXME3ZHa+TNXuEkos2vntqn9mGnCZfoE1pSnv9W9mpokA
Z+/MO+/4+QSL2HrMAVwCXEb7DAu5Ff1l1AtNcoOpfAyWGtrF0QeGiidARXpc0dyz/RbxJtB1xePn
7EKhCUO/wRVFoIfoHUuPk7AYpVcEz+aquwy/iZ8ZLOOCbgAlOerIDh0GhyKqEdy+PVpSpmebSk9x
j9AM5ClUvJZ0Qr7CowAtbxtUOSWlW7p9WnU5lrIirsOn/eqak7QNrEKRRW/NAvgSRl76/OrlH3y9
9UETAyuMhFmZIHP+aYOxGB7GZlrryPAM28GywAD/KKdQZRF4tmms/0xDrEE4EW0AUm4YbcMhZb8O
qH8Ra5THgSpvXEAJXuzEb3IPJJhV/g1ooKZsddCr+uj53L4vOcsg6lFnqzbWZ+kTDhQZ0ccXHaqa
+GpMN8OOMokjtLweQbRU/SxBHoEhLqJu3rQ5BoJ6Kn6yuv87BYSrQh1S5wL9wLqtQ1CqzRIeI9rR
Ugnr6JTfkl2k7Evrl1Shwh2895C59h3ecHqg3dakIxlVWDVWNFWdW3mSsL335uiaRGFuDvW5c7cR
bh28IbCCK0daZdiKV3qsDahSpekVc1eHrAAbjdH3Pvw/o62yDj5dI/IHEkO/pYqLnMl+cEBSJOoe
wEknzg5bPadrrDeD6XF4bKpcKC/5SVjlJFrC1BfhBTQzJPvBe9fVTWyp+kvVSKkDb0fE8ZZ46Qoj
2iBKdjoIaF8Y0Hn7Xoatb5iwisafW00aKfFMCNntyOdJUr3M65+luMXUujUQPCC6I0ybpq0fND5V
VN6JnocuJhSEWLKaA1Zw/5axNr4NsZrQonGNLW3xzBHIOLYrVr2t+XcV4FqBxowZgM00j+EnRT2u
j2AeNe5gnATMQXw4cTk/W0v2xZLKJUi0ArviMBtyg4T1hFWz4mvdQtzbDitoZe99CeG55yQhJMo0
OFINsTTw7UhXDR7HidlwFXL+OGYNQoAdB7lDAbxx04usF+F48+QX0Neeh42DK94L+YWDflcUtZ1f
I7nNVMwUYOrij8w5qINFDEv1fQM4VlVRpEElpMiRw6tWMueW5NU96jfb6ydU9gkfd/mzw1e2EuI5
+uGCAP1E+jyiE/n6F1g6WXGDq5Fus5Scw7w/NHj+rUlhe0XBv8u97Ba0goHSIX0zhPjPX8gGF0G1
eaG0FQ6R74u6ySG0hezHbp3k6KcV7z1cXbkc96j7nZxR9i1Yq4oki32+V4XHYfYaXHe5fDo4soZw
sOqe6mtERVKmZqIx9XXVvhvlzQAvrdboPkbR6P7wc5mjAO9rx6U8DRnl7kfpnl7xWAiQPOVRPbeK
Zr3K2vpzWWDZkJI3/3tr7yGWbDbci+cw8K6DZcWsjIZt9e1LikVQJYRa6kwOz5Zrd7fgzd/8d+2z
8VSjLSESnKv+IQ3OnTRbvS4cTwGm7+MCfok1blCZSmYBiDBPz3OIF7wnKd03+IFtHC0fhu6VxZtC
gpbdK8Eqpe+32zAyLdm7YgRgKq5FW5ovDnzbCbWCO7DyBXncBFE66lNK7y7FnSzet6M7C009XI3v
pV6EVv/jv0+e5Php68ZiRoyxkv9T/RyOBX3GhLaWyP3Bq22J7RSHfc4af/gbRbb5UxZEnseanZ36
bW/Zrf15pft2Mb+87MpwGoMwXECxNi2w51GRudODgklx+xXOJc3MsiVDvn2ySQXfvv+qhafCdgjI
8Wm8dCaGprWdA4GMgBkQh2yw2OMnNWKdZiLd6G5CRg0nTgL/k+KH0/V/Afv6R/MXI0dMycgpEkc5
EvMZuzh0fqj18XialqyTnRGkivjmwX25UkxobjzlsX7PpI3V5zyfXhCW+9hRmGlB72yDFhLCIHhi
BQc8LwPbQIGrESq423R6ostU8hwRyLSBohO5pevjGfd3/J4x9/l6cqUi5SEGD3tFPKrrrRD8a917
GY0L6JQC+PC5clnA7rLtXozn8AEWF908+PgBoXWFW+wKEeOE2xskekGdNpHc9ok4A2Fv0+3+umCe
+HhFYU8VYYxyrYvx06FeQWJCg2WLL/kwEmLONeZxq/PPxI+xnJ1stbuZx6hr2kT/+JdXQS4+MeTI
hVi7CLFLHcwDiKRQHCJeFRhkBa19Av1jWhUAVckRqL6u0gERlR1bpsr6EqB+rILMFyN1L0qA0vhr
ACcxzOyGmn80lr7VHO72Ng5i8cgDxHgcLnVqgxjxRDJ7yte7Gv1SgVWdWJPBbjvdp/eK31aQZ3gD
LgMRbVwTqZGDQpxKMeYDiMiLc8fhe08StjAoHOaVizs4rEIx2b+rhIqGONkXyQVb8nAQXVKwDOUC
rvf8dbKDbeTgg9/B1lu8zay5ArsxzWPCl+GM6bTXsCsps+2rpMHE1i+ro+DdKe9Z3fZgVIC5ZMF5
LlwAlG3k4g4z/YV5rE4paPng210dER+T421XXCK1UKZRw8x3Azc9QPHSYGKz/S64juvxJ7fpMi2Q
ZiZa5SWsaSfS2Sq6fs0lgA0q7VI0Lr1qxnAPsOhm1p3/OucNKD7JQP24GDFhfIXEjeaRQ1Dd/oj6
Kg7d2HNEqC1I9zlgXLbVBBRLouhwAMnbuBNfejpWKmt2lo8OQnfA96z6yJcQqxn/WH8d2mnJCJGC
WegQnWY0REjma3JmWLRT0J3A3qT53UNxhF5ZcxccMvRm+DQkCyo4W9v1hWanY6RALYG8m0g3BXlb
n+xKyyscJPcy+oqxKZAgzV2sy4uGVNUBZ2HE8iKEsTSOCQ58SLc0jPAzmJIzILXTn0PGIlr2zVWZ
h5lv+Gk3a06VC1HT2EAD3eoIh3lb0LDtAlL+Q0RSvZO8KOEd2WoD/cJ+C0oPJtbuvCevTCQ0/AyM
bTE0nl0ELte1VJgPOZa/Nk2IQVgfTOhEVtwDcFsOre2YRUWtAbIoecWMBuFjCJvPM1vNWQ5D3H4l
jY+LsdjCMIBMFVDNs6uhaZ3bU66Q+hDL+es8EamzYSX03LL8R2dIe3nW59/t0lnJvMLPG/d5ybGN
OHV5ydu72zskZQ+w2GVC6ipWY6ZJo80Ehp1Qd6U2gR5wRvU1EAYVEe3BhfnYSCyTPUbI+Q8nq09a
goRMjHCihMHpOw0zdRJrQbCowoSjH1fkZjnYzcTLUV3JXwpS0xVlFTZMXtmvPuxl5iE8NP+3yM7F
sTwdYEE8MFdsKL0SzhDjFy3S+SVQ7KeNq1SHXN0+H5x8KqRr7FCtsXVCx129po3YahSxnVg7KgTN
Af5zrQQ5oTEt2hks7cXuBgBUAocBBQT7Py/b0EZAw2tW4OYnGw0DL/U6Gn9qT241YBBVw1QEDrh0
O6TyLvdHEbboCHaobhpfewfMV+LPaRoAy85kbZSmCnOn62oi6vaZkdF4W1GOTpNt0pWYa9yqRVsh
jSPWYgcZR9QFSxJWtCVC3dWVZgqTEQPJpmVBdC4w1sQ6ISnkvnuMI9M3x6rpnHxzPRCuJimQFFti
Zdp3kG/8vGXiZR03kT2uCsdTXHd6+Qy2jVsPACJpDf1TQe2fGlC4Bt8JEBKaV01WlBtcVMxuTrXN
8Q4zGF8cMS2H7h3DKjrMwfgwIabifgwbiEKuIK+9UXsiqarGA7GozG7q2TgNtPdX3WP6DoenLeSB
tBi6cRPR4Cd7LaQuWD91oIvR6llwYn5Kx8sBtTp/LKtZr/j3IjBaiTcOue83XVqlhoQqCWAdZMfW
XE6wDufLc9SmQakQCzfeuPhcdH5oVbjVpQ4tfleaRWJWPdpO/q8Rb3xVyjBylcnm0vDTB0slV8FJ
7z9WyqjYF08qEbUp2maNLOMOIOtoUmCb73L5rJAFRyfTPMhuufQYdhwAOSDyghNxYC2ruBnak4N7
L20yifNCMAf66p7YkGUZrj7MqYNsZGrqQMXhwJGkyK40jYgohlI+ywhisncz1wJbjbH9c5GYSfj6
QUIn66xgYCe1UoRIpnmog/0CPjRQ6b9Rl4Pq7OmlPEqfkIxXpHbTP97+a/ep6EU0W0U+tr6IW1Lr
5WrOBGgpAqJ9nnPY8JgASvWM6BrcpWB7pYzzy2Act8UulDBmOt7xIiU0bMObbEpcEMMrYMlIF0O2
TL2vL1W1lH309DsU1hNay9tONlcdYDoj4LndKfubLaltz0PhNQjXlI8hBLl4cRAsL3fSQv+Qmp+J
ZU8bQlusAmJSc0+D+zf//UAFSvtiATkTgaU11Nnr1bAJyWh+Oy+Pov0Mta/vt0v2CyoMU4KPTj0/
G+nnFR/sMfv5rE0bKLvtpkHClrTMumDus0vrtVPKrnRnlL//MIJpI8qgOm5CQpNPfHcostb4lE/l
pPZ+kORl6HhmPFQKAs7wTUZo5WfinLUMJHYacnl4llJ+5xKxGCQ0ssb3OLEBSD6qv1Cx4WpEGRG5
Z7JmAUJZviPoQNUJ4PPdPh2UvmwIe/RF4UI17PyEhG519sxLi03lNuefK0qw4gtrYoC73lWB2hgA
BxsFTT3ob46urWmbhOmCBYmvzcarn3H8pSaeksYuD2WeJmHScKtReibWaPIZbrDtZ4k0nHJHPMyD
feUvHmLD1/9BEKpk+UyDHWF8r+T25nXol2ITy592BnfEh4ptJ+Uwv2ovUZZEcEq9fI4py4quh3MP
/mk/Fqku/hb5OyE/lK2nbDB/9i7XaVc9k9SWfSFRrOlk/1NziNeKq8xJXi4iOmw2SNStG1CfsZ+s
VnZfd24M0bRPkL99qRAZGiK8Q+M401zZLF2WdnTa/4f+lNvJhJsdJhXAaVOhuOckvUuKn3hGyxDQ
slERKJ8+fQE4RJ3JotUR/ENOEq3DsKKOcgfRIGP9FyZJ/E19vSI6IP6VxHk9E3E0spMg5sb8VKUJ
doJrBEzaLHy5N+ShkqurZP+55HC0OKGnuViDlEcrYjWlbfQSJlpJgazYgB0rf4Y6LubENDSfWQtA
VikkbfcoctLXSrSCIvx4JHRVej5jnIHlIYyPSjWQ5E2PxVFOVXTzc2MjzXF6mRUd2vXGYAX7oC5n
XdBCRsYFF0Hm0hZBNf7n26/F1xzwmWpurVIdUOETixt4zwcZaKDZmvxgSr1Hgb/29J7ju4hl678N
4ddVydwMya54g7gWytQH5ySzR5h5cX711mYzmwUGJTh3l3awTPp79LLDVWGBDfGY3bopO+xlYz/W
ig+N9ZgN013LlE09+e0VtiFZ5sKVF0ORBvuZcTBBnR2a8SjIexnYICr8k8d4uG2V20+oYQy1sWLr
WK25WuxDGLRQWWgkTef5bKb6hNeE6k6DTiGPBBj96nmrqueaGV/8HEJINPYfN3OJJT5IaVN44NuH
6U2y8+mfG+XO29pluumfdqbhe57HIZYdAohid6ln5VXcIKAFO4YodKxFIl38RPtLry38Uw1R5+qJ
OWJ1Lf9DvSS85VI6Z5Uuks9QEo0SA6/+ecmXSRy2JORTqxIU1GlbXoi8mIi1kxx20/OhVQZCY0aN
DmTUCI7P1+Blv/C+H0+N4/1XDOsQ3NC8BTKVV0SwdaOgA90EevTBIKoylk2jiwdcAxm26dh0a7j7
Z95Nl7Yef7W30z/c8U4TLFOOFYATXDEQizJ0E7j1pO2OdTsG2QzcaYqzKyulkIaGtfvPB9j9Da7c
IAhHYh64nL8WzWkBBxCSF983/WboHFj9o1Oic91pFNVEaHryNQFIcRFR6QfgArcb+P046G6hpTzk
CMzY4b97GunHSAwlKlV6A+HGk4TU1IKu7s/wQmY1veMF+ytnGhwwuE/UMxxKS2ISporfzLva5KsC
BOz68bQoYuMDwNn+6d2jG1ZOaEz0I9Xmw/UAUiWoe+wBcsIf5SP8GXnjrcMzana1mBeqY6777aLV
ucc3GBnvm+EpGNGrw7imK0ubEhBHR08hUNg0wvYUVfm0pr1+SCKJPVEcaBPACAqoRcurvSNXPbNk
rZbGmMk4sd0X4v80JzIIhkHCrz1lmdFb5NfSqboqHR7ovSm9WzWnCoBGXREJwPgwpcGfBTLAzcio
aw3I2za+FeA1sAZL12bMMv1x5vY9lddt7ff/qpM2NzQMQkajN8A7XRl/fmyVZ6sv/std6wLuZMdr
1wwUQfiM0Q2z37ioweSz1JJ0z6HKCjA3X77rVJJjVYeHLBZFT/1g/UMw4+RQ29ECX9Kp67hy4DrR
Z6VI6EkrIe4zVhrKwqD5zVDlx7esUmJ2cSmvLNEGEdZsD9sVm+2SvLqfYOim2OrtIoJgIweFGoYC
8ndheg7NUkNWSmTYqj9/r+c3p0jotdnKBop6/viuPcUcABLAD9XBtRhbinr8jlzZjSlmnT+DS3qO
FjXCMZ91keeI55E9wWxdHXjV/aO61+qXtrELb+9d9LSrXHkzIHQ94M9w/u7bsBBxZoBfi4Bn17R/
ut16dAm2fW/Ml1gxtlvuW2JugmTKhDPHhRiGgHdLKea/fWjM1RCmlZHqdy6B05Otbz8mDYg0MTpI
o+3wGKmJs3X1vc6n+dFuqKyc2EK2TtchJISpKIyl5q/3DudpE3opQWHshCqHHtnmXHGjS1Q8wlcD
oSjhbMjWkCDg5LeVdbDoQ7hCgQ31EQnzMV+Nqksrj05W4K2yjGLJLd7u+69lYlWCG8/183xAMbg4
WOb/HZ5SOaG4dlsFNNJZ2QjmhP6ep8Y5xFFcbCDoQJKLVnqEZJgZ4q+5AYLs07k3s7hM5ElTxS2e
iTfmxe2YBZus0X8AZfY4r6nLI8ZUaWD5d5shXVAcyBIwEXtOJ7MBR/dFCluexKVgSKh3tKRhjF02
B3wGYhDEP2mKMA9dkhYdxA+9+NXk9FpDt6jl73+RgePSlMDPCk/P8aF02qR8XgKaqPDLwjZJvifR
Yjia3MgEMarw/7NjUa2b0LWenl0iYcfXteeuzeoRRsSvF8o1cZkUBiBatfXUUMAdfLOj8OUr5tqq
k7i6aqz0+7APwzvf1zrdDv5HiRWFo2HDPiOCYtPbRZXdgl37bEKGyl+X4CbA8KoSTpByK+IoQym0
a1uWSM5Qn2pjttBGxIkJVqzyaB2OGp61kjwGAW6W3V1Bk34BHj6DayFsvISaPpk0CdCdPk/9diiZ
jm/g10OLHbRKj3I572cNl3OJvijLj8Dbpnno0PxxYX6v27cKPGNa7bEsw6Cr02vpwVqSkkCpAI1l
QlOtUteusifr6EBGrEWWGQRpSxXO4pxJdcKQSJWueijXVDb1RULPlhG9qsdjNHaGUHEj36PIkvCO
3S7GRoInSPtB1DlCHWfo67F+aTevl6VeVB6Jj27QpgjGefD2rXS7tuaX+j8O53uUCjP03Hz3Tdx7
dHw1JRRR7Gks723AbR60OByg/05fVEpFLJ8mLSSveKSqEgDNU234dV85r6nNAI/p7XVFWqMM+BHz
a9bEoIBEDflBlNdgucL/9euwWYtVHgmb2roQZetNYQeg7AwqZ4pB+q2e2WIihQLTveTGiO0uhZpR
VmjIcKbg9VyS6UN9XMkcB84d6RP0bN6KXoMCOITyBr4WB+Z3yP4Ml7P2heSkRjf1bDYMborvv09g
3F+jbcIGxfNNVZKTC2AHWUnStZ/DffZZB2UjtpAXpgdfGbyiCy5yjjUmZuRrjDLVI9lJXuoLHanM
BIwvr/koUa2TLPIIHLEeekKeeMW8L8SzvCJnKmo7N5XrQhyveEnkItQIkqH9s8l+TxxsanPXcxQP
xOFaBa8er4VUHfmZmCwYrl1qtLrNR2/zbMXiRJdO3pyNrh5mj3nXXx+/HRM+F4KbZki/8fqc+AfR
VmwRPObQVG49YL34F3LqvZ6c6fRHr4eYcinBPEKwwiMWXUhS8PzYy3w8cSGgGDVO6XW5Ohocv8tj
Pk74+Cdj+3+vOoUKqFzwo6fMqHdW9ztJx0Wp3YMSCOeELGN4RciXMsyMNpE/E4XYLTfQPPk3S2aH
zWhp/C41VQ5BfMi6rDEgKoA3e0d28UFaN54jBITNE3eZ7zHaRRqM0CACxS/E5o5Cpg1Mw3RyeBsk
CMGTAg/5YRf0T3iZN1o1n5Y4EQI/AmGmR5PMn4/ewi6/BsEVSWObAdkBlQ7fPLqxbmvsGG7sOc7m
EbH8qd39awyvLjSMe3RgjdP/zakpQfuPdab2gvB+rjN3S/e7Hm1dThJutuFbstddeKyoYRbfR/tR
gsENSZ1/UhQH5LmCex9MfH3NKz0D7wYU7XyYsiJScRhICwh5ovtuXxrZ7M14kxWc67rhSyHozWwB
59HoSiS97YNb8wXJMiCumrs7RkGxiiR249WZN0yG33G8LBhO9vzQttzSJ2Iue5lr4MAZX6f6try4
HBLQyX8iDrAQJOuGwiwFLuhhdTbevBssDziPz0SEIkbPrGUyFI6oOV5Ryx9vb/T3ryMnUKg/ZClc
yv/dycwmOlGbEAnnAWiy+p58oElgyJ1xCSB3BvV5lDwzkCy/Kd7pxAft5npFO5fSci/TyAu70D26
nduqTZAv9sb8NTLt7UW12DgP1JkCPoWZ7rORTV96frXDxyP1JM+2OaABwenAINYcp2SSDi9z9ALB
H/prFrXBCgZQw933AmLDW+vquH1KI6xFk+Gxd6Gt94nFinkdNz1ksLniwGfVM0FgerqXd7t3LK+2
jSgZVwZyiBX4sZfEqMkiaO3W79Vins26P4tvMZjZ1TNouaqVbzcfIfZk0Yzoghi/F59ARHhyBULT
vgujc2tXLrfHYpPxVoJYpJDxUNVr9nyUk03rAFNh1f6CascZEOeYbkV4mEZL3f5L0yiC7qTZhz2x
qgTnZofHdQ+9ttTr+XlSjg1/u/cnIEyW6hVU8N1Ay17C0wov0jfKNH+Z8TsJpWYWCVkgnQHC5Es5
nD1scTKq1gPvDYqOFqoQkN0Is0TWIRcw0i/RVKwN6qufHj4jVzz0dEjcNbVpSFpi5YUtGV1GWKER
0SHA9CR60ouk4mv7SXngaAS2dxeQxBZaJJ4Tb7wC17mg031KNCZD+Lt23aU+7QhhnfHnLYOh34qa
8flyQ+62vrDWWbWaPAi3oUFa8N9LdFd3raPaopY3M3J7p9hVCA634cu+Y2MfW9bspOHmRVQNNjeJ
y9cZ8x3DEAEFkZ0D1QnkGERw7D5qauypmcoYHy06XgyVXw8XqpdUSx1W8aP6WTK7usDi9gxwq8EE
T9CiWIdY8Os5FbIWKG0bEHu8iO+hlm451gMiIMKzB9ebwgUd7+EWC/4kDgfAhN+GNjVfcgmlhxBP
TjeY+A8JNUjpnsIkFBCuNFjcTFouhR5tEgS0tFQL8S4NjZntU+0v0SptRKAc/jtItFfXeuuF6yEG
Or9bf7GKz59vE9ZxXwudn4xzxjCtR+WijxZmQf8SdlziSnrlTMPUZBYsllnixla1boZuHE9E+HT8
gQVEVbb/ZUi0QINj+d76Kr5c8J1UIDYnzFzJmJDc5YKD1doN6PhfpPthRPjbPKM1buB6St257zwl
imwZyP/p3epNB8u9OCZT9R2IR+GxcjsKI93U3UUOeByGEvOFkDXBM/cUiz9kr0OcjVg1i5/2WToL
3eaNyIErQwOI3CebnR/WN+2Dvgqw5mGLYWaBr58LNY80rtlf2fgwa3w3t5NI+HmY1yLJJEN6pruX
Lzi6Kmd189eyeXsRUEynLd1tVXFxSQyKlOxcFbbroL4zDCW2YSXw3l6GeFdWAO10owuiuwS3eh2d
87Gk9LwJmHWT1tMMQJ7mB/wD05LwQsfT8wmajnJqPsR9dTQXtNVKbriTihKYK6audVFaAnEBIt3n
qXFUXFDsMlLbZ14gXKW3ZmMbJ/eZm3JQTaoPYC8Wv/BbOlVBJ9p97aeS+mnTxMHTZgoWyfOHo+Pq
gqR7lQyVjffQo5zgAnpg49dIxOIHIVu3OmwZqIEKVggygG+bRW7Qa7m45awGh8sL7QX0wwbre5aE
Z4hRXd8/42577LqxK/sHPfDVISFvNdjMG7+ACHWoso2EPb5/hQ1Z4v9WYRn73AbWWyuS9b5vE9eY
fP/iq0HwP9yR5vitr8YHqPfvUiC6dzw3nx9ANuDN53yKIh0NwsqoQ0KjPeBy4w9cfw9At67RJkIJ
nqfHkqazL8LxPbMJWYihwCSTECTc01FzudZ13g8WHK/6s4wvvedU97lX+1XvAE84rRykzLPXbwWk
S3/A3zeLBT0SqbuYKZzTR9feMJQe8ir273x75ak14fECmp/0TMHDwuhRJN5dRGG9m0VFvWmS+NBJ
tXEilXSMCIQ5ntcdzvS5QuAF8iVXEmDLjBlcGEE/kMeexoag0dVzq62NTN/em+zsTB7W0eKMlXAw
zwOM2s5r4u12vOQNaGQwnoEP8EAspbciB7H8QLojjtl3idLhc0/cNn/vi0Nci6Nex7fA4mSbm0Ze
zItcowGJ8gZbFZnQpO5uB4E/46V51gXjv0xYHc8+5FZF/5nc6A+WW2WhJqZ1yQKtgPTPPQ3aYlED
QrB1KmKYVzDop0DfiWy8LnZJsr1qwJGwFz5FfGtMrwYI8PPlEO0MlhM0aswWRPkAFn1/ON0ooLdC
TCdEQBTL2mdNdrnaXr5VVyiMZux5wiGygrQ7WE4C6n52TGLTV9zIJA4ahVpYO3QjrdQO0QEHMBfn
xqDml6ga3qFMUzobstv3367cVoeiJ4PWbnLsnqRRaZU0DHQo1LNJzT08SJheL+Eb8DTmd379cYhv
5D8ZlUyWI6DYpqSIeT21M9JKa2gpA0xFwidLmZzbU9RLoATnsNh6Pur1PU/2PAZGBWF/vpaXiYBv
FNGL4xzPgVEwSqHSsskYXe8hg6SmIkstVa1n9Tb0Y/U63KLp8zejLDi4OHroDCPCx4KlcLQ3QYgy
8dnMvQSmZZWumzLGozmVo8eYhQd/PLPP5kb22NTDkAot2B0/qjPyx85cMtO7cJg1f8qLQRQ7jQPP
+ZD/UpVVepk5+30mvLqqXOW+E/AyUO0+K35uUPMvdbTCkHEvhgQjeiyKKLc8J7eJbMIwso65UeSM
yDZlojoXrCpPlRdqOrXsfW5R0UJecHp/F40bnb5yCONIY1cjY+hjWXKwh/pK5nhaRVJKjgSgdzHs
mxXi8PKdyzTTNP9wzdSOorgZIuD9XYpL8VyoQNpSd6SlDtCagLTJsFl1KkZQ/wPrPvNN/5+6Qkwo
anIeKKA8w47kI93zpDktVuXKDHjeVd/thjMU4MQQQ2XIDmf/bnAyj9F8cIw3vjy47Y40buWzETOz
1GGkfG7eEhYEI/7QoUFIiXCAayVBChWhp/4P63VL0PpCVj5+GGTD0De6g4eK1tXE/qdDtBuvVpKF
KuvgttVdVQALOeHbYA5IjlBCfPa7BqDMK/Ssl41uaJnrXaQcgy8D2tgJ/TnuJhtYCMgBdmUHgU8+
cMSMMaBzdz9RMph4u9zwf0Vqoprn2e4Bwb/xxBDjlmf2bmPFwTED6raJ/UPiuxDyOtz45bmX2LMX
O+z92Su3h+GksFhfJA1Kt0Xc3lv+lrinRm0juvKlb7oL9aE263a38TYrs3AvSDZujBJSi3xXsMsR
r4JC5RvBESkQoNMancu7wdClPiLgSCdT3N90W7hM/nvVZcwTDIHkX9ZNPCmNisXv5l2BAAhsMouN
lb4wI7TA3OgOeSrztYx1GYC6GA8zOo/X0xStkEyEFQQjmveaHye/6ZmcOwTz5G28035ckXkIC/nW
IavjnfYMtn1C0q8hbfCxpcu4xgH3jfPAMh7EPKqAVIlRtZgcMo1ldweeMFal10gQrYOHuQxqXrRw
OsZVNELXKhBh2YYzrIhCVje8Pn8YYKIX32Kfk6MRHBSUQk0zz/gJ42w0XNPEAC1a8ZIzhhqk8D7m
KpRFQZksUXFF0youEWFpV1a2nX421M56lt4knRBuBs+D8XNveqcHeqvWW8M3Pn1oxX96R93rLPZ7
4XWKBWLwGsKvqUoK50HWQDLOT4gcT9TtqCR9MATAlM3gVz8pSeS3N8bnc+uhtvbX7nT0uXGtpNCL
NZvjkiR3lPlgxyxJdNf3DnpF2J6Tt/kXMtd/LxroKSYvJ1bQ7r/Brl/CjuA+VvoqokzwHXo02IHU
YLx2nB8KvTbzMvzxWK4/f3jOOfbZKAJ43ufrv9nHEfbWjFAtxzoAqoCX9DlGacT68PILw9d268zh
GblBsDwZj2K4JNV04YqLu69AdYM9CycS/czbPMalzqJXIwkYEUpLprVbfMMlbfL6CH8pMvhXhhkW
c/hfEPB+2faNR4ulv16ErVvNuTrHDcTpfhJ/jR9G2SqP0EznRtI/TZl3YZBsbkzIi6M12zYv1wkc
M+1BEdHifjYEq3JN2ZTFy8hS9oZ9sfMrVKFSy67Ry4N+LGLzzuV0aS+/spOI27U0fgjMjyhLABUl
bb7MMFrQlvLoDDqXsHy59Aoi3QC4GndUMnsGKt0taP2STOCOsfTWlTO2NSez6MCoVT3lkMl2lLHL
rtAE9HNqeAri8/VqZcrp9XOBZWSXehhzl2Ey8grcrKMnm7DTGpuaCH+tfdw/eoyyfZDjkxQK6n0x
MS6y7OFqFHzsjQ8TC0oJmsoL2QnXYjbB0F6MzMx3YBIduIf7My6fFCfYxSb4BBkrxT7FMFMTpizh
efHZyvWjW6P1gz3NAIiZjLWi0dvKjW2M72zomfMO5+E9J4RkqLzp/PW0JYmjm6tDZxT0r8FBPJLy
77AANYyuozuDmCRR8TvjT9Va/Ew2QXb54kr1VgYX3nICfs7Hwj7sfKMWcvwgnbKJ764fIjqzCppS
wtcS4jrtjeauY3bdhCnuCP6AI/Sk5I+vfXzdhZuR9N0PrwgiqllXdT/uvvu66npHwxad/750TmzA
Zejw+982RNBbZzUGB9w13KhMPFf8RqvllAKTsDWmALW5bNUaZ1Pq/ydDc6xzTaGmymh2sl8N2Gxq
T8ARmldRorM3CeULbxOf2/daTyOcdo2glEUurJah9sdu3r30n8jkQ5gOHQRbpIwRpaYeeG2k402/
H+ucsQv5XdRs59DmhnQShlKKgoDWEixAkoQbJyVE7T7Z0A4JZpZ2eqUjnNw6neSvi+9utDZSwZcx
4hf55DG9gg/OST6F2OhjOsXN2gRGxX9TizDMEJ/mFEEx9dp6b0ciEmOI1H+eOHlY439vW7Gj9TQ/
38F/faGDBvS0H7eXUx/sYA91sGTEVybVR+fA04zpwnN4fDXQ5zvg82rlgICGcum/P13tcvNZ93at
HQncAw+wojKps/eqr8FCZHigYRmV6dUct1+tG6Vg28t4nj+pfRO8Sr1DY5G3VM8yM51S9QZQ2hDU
mBG4/7zCVildQdN+DOQP2ljQgjtnJeV3YkzSZ/qLRvtc30yWjAoSLEaLpPmLA6OKO4fNfeJ824aM
Zr9ra4+EhpoHE6IzABacn+NicIBHsorpodDH91quFIXu1uO6pqrtxevoCMGEPmNtlTh0MeyHT8KY
42mERmvOUmVyugQ23Pl66eN8B6JRtXIo4KPUw+X35OucFCsgLHict/+mBuB5HFHVmWgPG70pzwLY
Wgdh+BU/2dV7jAZ+7afDY+6gm3Q+WajoWpUaU9uWoyD9HxJZacXR/+pUUAg8Qi/+yiaTOxIDaJuH
MvhCxN/iiAF/cTMWY1vh3lNA14mQawbrLl0XUUYjvMPFCksmE6UBppIkz5IRRI4Xj6tbTrbWK0WR
6iMoTNbM/C9FIiSpHlABN9LAtya/cM8WkGwy0nmSpLujCbxC/qIxsHf9ibfimpr4sRK+DR6Kc4o5
L467FiQe9M44D68rDSUoqH0Vvrv5CcuNGTjgzZN9bqlGd/HAxMHp+vOVTLMRXa8SxbSo+lN08vZa
v1RV9kn4hovo0VD3OCO6kbvmiu7LGHQbM4Vo+jyuEuRK4A0Bfp06lSZasH1kjqtLpROYaWJwC7JT
yKaw/4wCCjg3aO64+W2UG6SE8zu0C8bBll6gBtdsCOaF5UO5sMzlQoAiJhRNAit4nwUfvBGbHsOI
2T8WG05gmWwOK5/qQvohnrQrMCmjCuNDrk6HDwsqV1wXeYHG8cIkMttQOQhQ5Wa8OiTa9ygeWitc
igZE9nqa7UdIRE5HKnERnmLP+7csokGZuiAPyR0shdqHQhqjphSgc+NNI4ZAXZSvCv1LxTyTum6B
V8DHNaVUyi0erm8lKQa+8egA8J9SvRJfFqvPWUoHQ3tIepty48oxt/HVbyOO5bxGli4VenZt9YFn
JESCj/lfsJD7vnzjTKzdBdWay+f9maeYkxZFsIXD3Wc/z0W/XkCmJCDGxQuR2YtPw1s+owEQyVZU
KPB2kI37WcTroXp1Ic8ojW1XnAFo1SjogZZNCihm1q9uSFWhVtg9fWwzD0Q2vwp/JetFPCtg0mnj
tpPTcA7TZaVfoaY7FfEXB3Ml5dwqQ7WtA9B+B7F6fy7VF4jvAEGbDlkkEMxzknymr4BbKEoJh728
/6y20EyPqw2Cf4AoPcevstoQMkMpZBL0LMSDa7AxNNgTJEGEJ0X+Xpii2+FyH30J0m9gn5jFQGKg
79KgcwTnXKNQWanI6ZIE5ETvZVJ3K83FEdWlLWO5Xm/n7dZCeRS+351FH9zE9fpGFsD1C1+4ujwd
dSyWjueNyVraTKnV1m2tRbSLCtcZYhDhhYpVrik/rg/+52Rb+fYKm9fsBrN2PGKUx3lZ3xZApSps
hQJA5dOJ5ipy2TAkz+j1KTlQxpplr3dRdkhFM74ElMeevyoEZJudIvjdrcvr3CUeCq8w7XdiszxM
D+cM5mE/koPbFRoJdfNrXgOukVWrXEM2iJEJMJAi0AvSGu4NNIGnaELvjrjRSGwHMK4hUMbeaRcF
Mjy6EM4qNrN1c64/qRxfGzEnrqObV3mS0ttmfVOoVF5ljoLAW3kghyuKcXHnk1KrDQFFOVgyE0Gd
+DVVxbSmfim6SYaolxSyWKvK2vaLiZS7pBdkL3uK/Q8BVbalvozRYPIPIxejNDabV2vWIJLZPZt4
O7bJXpxq9YfDfuvTQm1zfYFLRF51V/Jl8aISFf/LJnSVqkNv9SfCJibpTk6CHjOXPx2NNJxxnvSb
qQ7hoysgxOF4Ya1pdQsLHRqn6hHZt/3xILnN/s3WHvUshJWUrPVKKdmXY1v2zNLdIXygFT1AZxPv
kzsX0wQpQcLF56N/cXWxwWIVJKRAjmAVYU3lI0JmBwRs7x+WCTxd/qUhdKRgtTNBOl45JYIsh0ji
PGwgMQXhJPckO/T17HS6nWlrtx+vaW0hceOniSSEEGPDSqEaqH1myJ3uOVHEvoOiAiAnNV8y+ZeR
nCqfx+9iMWMSpyruqy+GJLT9BLENxlS3lMCn/CcUsrKC+5TFCTcIdxp+a8wqrxrpFEricMzuNond
RPCqvzA+vdXvgdfm3HzNR6oM23yb3G6GI9RFLhwWdj/edxlNvRB5O0pkw1Cg4iMYvsausFtdQKba
x2pL9Lz8CsI0hlXMSOoHi+UJtU3RIdCkONuSM7bWFW/NDtaGN5FPw1kH7YsLmYW14lBNXgp3YzFA
ON/yWhcN4vDYoL/QynJu11pwraVqdaDFifv7VrjewsdeeKmDw/slsAG26cPZqPh61Df05Ulj5SnM
+uZ5g2HKRZY5CrychgD9y7iukEBVrov8LwrkJZE5Yq/m+5mUkuqpQo9jObUnY/4MPX8nUe9zE6s7
kIkeP9qgQGBJELOkXAQ0pwwp1c+18lWo+NGdzC3RyFsKiQArE3/FaJkS+X+Cf8ioC5IUV5tzqIDH
ArOiBAok8ChtZZctZ1Qeq49IitPd10UQbm25vcQa6fPJS0TbtLrDesfL6+QZbg8wGRzu3SdXlnM6
tZnZ8KeJUk5CTovFUSXiQ2QSLzeI166V9pyB4oGxU3NHDO7qcC84hdbTTsuIvdX5OLBansaHrHID
hF8xERG4unV9P8Kiqa95pfdbbCbGJOGGa8VbDUlwUUHthsloRTiekN3AuGA9xZrsW7CbxCAtSsQj
uy1XatzyNuVfZToPSp6ZCJu8Zka2PU7uM4U70LZ6exzsp08D7SbYkeGXzQ2BguoqsE5BO38JSwrc
7Qcm108hyjMH2iOcar2apzI/CXTZRvJrQ+V8GXKZuj5CmzuJyDWN5CDKEwSKuw7mj7wd/ItdEv5a
VCAYdbc370WU2z+ugYMuxMBpSlD7fOtV/bVbbPRbQMgqonvrp1ABx610CXDOF13KMWNCcz3l/MTZ
lN1TA5TJ5HTheOpe/A0TLkFKBUoOvTeqpuRQSB7XC7asD8xyVAubYqb1vas1g5RJT8/mw+4Wa6RZ
rvg8MZEmoh/1k1LpU+KYytcCepiCrG/7jEf3WZ7WcK2t3YZTCNkkbUHdK4j5qKhaznRd8p2gE3k7
0x5LEOQ2IDKwJoUUz/sPLv3wCT8VHv4CZfttNKr43h9CtNk0GD0Gt1CJsJvQADt4lLOhv+8KEUZY
qHU2h/128LcLDPd0oOI42hZ2iFkmvv7vH62dJ0imKm1SVPDbLH1L/wr/Ur10f+45leMp0ZtWZHPx
JKIz7nApG8vHrtK0P+qlICYw86qmxe5JE52XAc+j9DXmggDq1y8NKDfpmMJpc6rkCSuoAZ6Otb+4
uYnYXAhaGT/UdF4BuZG35nXurdDnU8yFbHnARSMpz6rxz/S7dE2uSYrtXWK2OBZu4hKgo/72gt0u
PwoK9Gx0vT7IhMylh5jtNRbaox4GasEdA7VUBZrHjzPGqPJK7lfIzBHnJQYv25DYNqddBEEXBTPJ
8mE2g8UHNIZkwrS/VRTZxze8Nk+ZU9LIuTEMTCcEOF6f91FVfJrtLIjDgEkwVWa5ZzFtBnXqHl0J
PgqcEmGT61CW44X4Qy9Dh7TpEvKCbJYTZN2wG5tKF5n+YMvz91Z2DqaKmSJG1U2aHBwBFOcPMX6N
xI5Bxifift40ETep6z/l/At2rfnPr4qeoPCPPh8BSEw5msPJRVQwiftAbZQq/1AXfMritAibJFf/
wyWY+DMrTKRSNrjuBqSb3sWmXOlTd7nZixgkZKe20QMXSCGlr4XbFt2tjyE+ZqrECqjip/WEZNDU
AQ1jePuNfG3kyrLQmHhxEbK990erjwRpnIuHYWiL6rL6/PRTlR+WzLFrwZtx48/ov7Co1ALKEeu9
NCixEB7qE2xscXem6fGVOY5kdpRG07se/yqJypwms51W44wogxrQgF9n0sflkirR19OMgsJzpM5m
yqBqo37NBmy1QchJ4rqt4Gj1FC5DmMOZN44qMJMTY9m7BdYH4zW+KYx15NHIYRJrF7+poXtG3KqC
Zn4E4fYCmtdmf1f+aS3+oH+rYdheI+T6QR9mJ85X2TMt5oM1s+JHilBVCbPvRGLTm+gd9DGET4go
w+v/7eOE/797ImaWiXfXHzGUHFBZlt/HljMUssY6xhc32pzXmnx4oyRCUTOD1SkObk0zv5JPVd26
WktrDX6LJp6PZAclu/OdiYRsf0HrvCF968zYrWs/fxavvJGn2+kvWO0UafmM8ux/V9BSHb/6FZ8r
sM3unCNr6I0ckpdWNtlKPjGFvvn3vq70a/gmRwbo7mO8A6fIZ6v3FkG+XATgqcdiMS7aVBXX22Ur
QeM67CEZkuQa2FEWnQOj+VVGn2xKL58ZybthilmkOwSNOyLapmWUHW929uRRseOc/klFmiAtxEk7
sB9zgLDctAFHUL/6vGhqQq7R6NZuZ6Lk6urSRnyRK3CJ/4kNViKfJERS3r+e5G6ou7KQ0aauiTDZ
mrbRRthm6CS2xlkDj2YNa+uF86YTNmSTD2s9oDk4EZsGUJxb6cR8NrYsq1R81XbSRANPibQ7a84W
FYQarxjU1Rermkl39A7y3Q6gRFcqjca5Kuhd2tvB09aTE/HSHw1HTuWcezi3tZoive8w/WaFSWlW
fnQtr7me8y7ghOPzN4y8c7MBZRd9RMW2u6o2CLv8D61pYSvPiWVOuI1l9Xl6/GUM5QFGFP1xy2Jb
XgEsN+wwDYYE4bBl1Q6+wBNtXqO8llxAhTvyD2/IW9PEvTkjdh/7dzvve3zzMtuKwv0RvEig5n1T
oYOG/kcMVty30CVPLfjwOw39My8u2BE0pFxHl0RAr/IKdT/iwsI9J4cLPhmf5Xw6nCsQn45ipwsG
+A9DLUrQxPQEYj6CJy/FF7ZBIK+JOc1jkQcPwaYW2xemTjYHw+spqX9pzmyfZfwMP3QF29baZACo
xh1SoKZ79Ap7c3xciVAS4QjWkQq9rsX7XPViCX+FzSREXvxevGlc0Q33OCh28rf/3wxqXdHQ7SjD
NZUPHJadLQljjyCWQilO6pk3J0MBGtPQmAQJBHuxNfsa6V8HYR7LlQLpMtgO4hbSLVrYPphQ5FtQ
m73j8qU+HG7KuhytsvvVA2wvVO+QFeFNtu35jOjWL1GIlH/dvRQK3xpfDCH6bsXiZlAWx6OABQdN
WmACmxVrkqlgueZ7umSylvPAwilHc0ltT8VdBHKP6p1qgAHgEosprKkFpcuONsElt2mcSj0dO1tH
ulSJ3R6L6puk59ILaDVo7KoXSyiHk0HAMAN4bKDzM9ilfp2cdf6y2+97f3Gk/s/coOGcvZxP8UUX
sy/XeYkIfbxeIhYn8/cCrxCKcXp9MWVLOFbOIKXA4xJAiR6NbGf7HwqlkOPNj10e6CsLFB/5UsvM
7lBzl2gsQxqFcrKvy2+QvQ78C3iPzgsQSR5hIF/GpppBxNGUDaRNHnLFWRqdB3vlQTZ2wS5tUys6
hYZ77L261QPDdqZ1AeMJN5blSvNrknQw3J9PPEy4ouot40nPJrZLgjS7NLGj7ZCmdwPXUWVOcGgT
TYDxG/JrmrlB4fQnciyYx0JYMbr4AK4Ey6DZ317qCaVWk6X1JTuAAalxhHh8EiHhpL2fNo2ZrGMb
l5VRfSz78Tp0rS8CJWTVbjQFYS9oJ5o/mZ1UBarP09ZJ5Lj6o34mgdeRNAUCtT0EoPfQfviYWrZD
bF+scUc+cZz/k6rb1At645lcuruQPjoEU76bwuD0nOW7s0fIfRwoF+S4lUrvagPWsJ9MLRm6tnv5
nJ9T7y+KtUjz2VFY+Mw1rtOO48wpwkSR0BlkiIRbwaMBlyrg0NvGgyLbCnlsZD18MRWJcJyeIJdW
BjEcvcJU9SFASE/tgdediHkCnOgSmhKMf8YV9+Md9DaOEOWue0kcLOm0qo1d6/m5jriUDOLKiRty
O9L/6V7XbH/JP2YExZzTHTA+n4RkAKVRrB5RcyqpQxryfh1f+sNM5h7HTDdS0oAS6ibRWYjzd5TB
79/e2MeI5qF3dqSzUfn6TFz9Uhelk7KBJKA3Q8EZ1mDNx0ASZ8plDv2ug6n+CNPF9Uq5K/PLOsq2
aqhkTbozzDax+qlv3d+YX/JMpm2T84RJjQTSLfxg3a0z6FsnG0BU4SH5v8+7kawliYincRMSRLE6
FNfo9bUHgmsZJZ8htJqrPAb94DDanEgkzfO4limUhAdNuoKclhwOMLG0ZsjUr2L0D07NoWNe/KQn
hlWhMQNfwsdbtVpE3oF2tEkAMUtplvtxvivujDUZBmadIcVa/mRj8ErIVKBhnTvCPly+fOd0pzQm
4dsgGvgQJSLcBvH6dyLvohhWy8phgjgc8drKlLDV2QVYROlh+xhx3/i4W2K/yfz26C4vgbSWkmNa
4WoleJq8dHEnF5SDytMCclxgD5WVp6EcVGzkfRW04KPNes+v3fPUcHbNNmVzR9dI+m1TibsMnMEy
toIT6B6FaPW8oIxBDIuhrbGgQOsfrEH7IAyrDeEPcw9xl4SY9+T9UUWglcIe8RLVSNNGyrZjblvs
MRZCC9JwxJEAkTqpfaQRAUKC21xCwn4y83PTJ0bj8vho4XhkB1IyGPhgICFgRtWyajitIIbewMwh
aBNiHCzJCx6CWzprCeEZjYHaV37rrQ0hh+DnL5CW2vWuj5aju3zHfROd1bQnxe+o+DMyR6X0y5fO
4DEElTMGn/lS3i/ujlwI2YEAM0Pszmd9D7oPLdGiTwrqagbFcN6UmL1p7dGx0VPqyAqnVdjdTXNH
8xG2RqxhHoApki08p7EMHWaD7lhY4uv6DkqVGKLaOGPPj1EQP2pSfwVhEF31U7bYYJY6AO+vwMjx
Edlyw3kUnms8xSSYkMxDeAjABf+Y/BxqSUXBDm1D7/KzQNtziWB/2OYDcleCkQfNdj8PbemvRr7m
IKn5bIksljqxLyz51FAIhc0clzfAJx5OfGCX39rgoxEyb4vDgScsOZ9Flh0gBq8Z8Khtfe25kTpU
uWexYgP/3AkSeDlUNwW4/oKGpSiHjj2EQ1itUo0RCPIXRDLxP4jDScZVyMVRvfzKjsQKm2BE9nIc
ebQnT9A/FV8N05/rGAGOgwVtw0eV4SV2vKdCokhYaIbf2+lXAeFYsgIVjof9ue39sZtsmDxQEif4
P27pMI7I9U5NagziNVuBYSVNWeiUY47ZcTA6IyvLMNrLpEPO7YMYvTk4zFUrYyzkhvYhmKZy9Y+c
DGBZ2wOipXV9UYLnrzxjY5ZFj3DPp3n4cs8U1UWQ+WpL4vZEppVv0UJ6Ae+OmpelOKMRtI74Irv4
bc12AmCrQywBWx1cDRQNxIckZQJXkt27vemIAJsB72ku7YpZ2puDmcoL9dS36XcNl74WV2nZhjnJ
aKr6Ab+H+P5lUzG79yVVYBpYTuHxkoBXJsd78EhgPujD2h8RxKKCfAJ2tZkSRFew1fLKKQ58Vg5y
3QqDRnobslcBp4GzTzQUC9mVmMTMb6gnlO9q1lyfyRPNRuRSAI9/jFaWdYIkDtg7uqANKCweeJnL
yp9EbTV5rL3vs95+XYDULciVwLiBswJGKcc/hbzorbdML3mM39R2XqaPkrJBUye1wX+vmu/Gf4fW
Q8hwVeWkX6HLs8BiSMsbzqrWuT00TrDSsWcO1ZKnAqbT2t+kQA1r1E8h+xru2nbUCKgMKgkrzI++
izY7fwMOryOqrZYQiRiV9HtHTqmCh6rtoeA+8Ou1gfS4eX0gHYirNeRBbDisNh3ZLht4JQWbZYOz
lg3FE7UpcA1+9lQ3UtqxOLwvHdwrsqVxg+ad2VNdAagSNUh4GAoHZpaw2GgDioBirBhcBOE97VpN
s7HkGTm3ksZrH7cHZtrLPdGNRxMrQcn63uJjO/rsiqRk1uMrnrK2G4uWNcxH749rKUj5J6r1ru9Z
eHR1W1QOkskLZAFU9RNlna8rCv0KKkGR0R/ie3fW2olKUHipFt6BVRAl7yJeBMSPJRiAmD47LscO
tqnguV7jkseQsLDE5Ex7OEMR1+vOZao+k+vpPv+PHCrl29Mk9cal/8sEep8CKds2dWmSrApRu0QW
bWlDz7LZyAQtXBATSMzY+B/bOWuT3AC9eMvSkkDW45GeBRPfEh82OuqI/3GgeEnIlQMLzdKhje/r
30tjz8pA9H2AsevocmJMkZWc+vB7rXAzoUkuanFQWhlek4pZrqnnhjkujLkDhDis8JfAyIJHhopl
IUGjupPXif6AbjkidZsDuPIRuiSW11y5x9+S+sTqRrLffdcAgmiKN+AXkuv6GSkMNHrOPPpMoKBi
hc1lTXv0Qe3TYEEylYy0T+Duk+uBVouk/bCr4wPexSjuVWgZYpwLgiODKh5YzPSvDWu4UGcM+JWx
duyt35LP47YyKOGI5mT/oEVDCgapDwd7lG5WbgOclLwVGN/A40QgtoI6rlevPLF4nKWc7TUKa/Hz
J3XUvcIjWs2KyrBC7t+NWEMN5IFGqAfEm9539FR8hOQ/HfVSux/RST8DQQlaicuBP7otuknSzQDS
mlkj5nBDs4mJI4NRXxw4ajQSiZ8UppClp70vLR8ZQzCF4zol10ugxEvwTkfpgCV8vi111MTtJZQ1
9FK7twkRw6/JOGjb8y3kGJ/C+4+0qwW8CGc9OqBhnnQF5mOFReJOO6rxoOQxq5U+2QTsLZU2nrC/
7Tzsvnc5dG7LI8hMHyiSgkEYBoHjxMpF6KRBzaj5UPPU2c4go/tdWx8aE0Bah31+zEoaYQTPh9Qt
PVwy0txh91Svy9YjEWgNqlNLMcLtxxaSbD4aCq3lH+XRxgdnLPRDc7BRAH6TmxgFQGzdAFHeMtqC
K843OHwW5mxBa23BhOtXVc0taSViN7OLHeYJ0Y3SCl/HSKhLKJY3CIwFz6cYcNG12K8liUYcLGRd
DbCOhWCYtj01Vc3ybOh8rPMFHvk4ONoXkxmUeNNrVS8167v8dXw0n5ST7v/ZIp1pqC6YfGhA8dKL
Cnh3nhYLxyXIL/FF6ddYXoD6xwK6y6kTyEGry89WTOqSXpzWSAEd0sXN6bbv12O1IwJO5jxVWGEw
uz41Y0zOXxcGMX3zuhFjMVxczAdV9MuDDZdlKKIzchPnmadFvrjfcnmtBkH7ntxr6QfPR5p6WKn4
G1xjUOfsSBtve+2nnz06wS9778nEYZTPOWsXfJiC3juiG3M6z75XEAJP186G7PSZ5f//WL+61zoS
Zp+mf/7xsePpoqTwabdw+Dg2PXkvM4LUFwDdUZPYBiWaHx0s++0qQSk4YPfbAQHyndzjnie7YWvY
ysXnuiulWrZWbkLqa2xuLhdbXTX9HqJsM34e2CGD6Fr40+dIWz/CdYWpF13qWtRGHwMNlMRFNlIv
p/+LhzrRvRgk8kLx4hlmubPhAZ9+ynk38AIJAkcRZJd5iC8XNV0IPdjIA0htXXh53vDlmYPB0PIo
sOq8ZurKegMsAtVlM/0TDReammMRdwTHMG83eG6wpVLwImh00ksXDDxWFo7cduiFB7wd48HbMDXC
+uhjJXu23+Bbe+9ZQGv+9iZ94IpVLBUxXp/erydfHHQA+RaHIeorOzlQixslQDoIYfYB80ux554i
1+I+4jZYVGoAQpELIGgaiK7VWCUIjUOE7D736/LyjU+1xHkMWlCK20y11pFbNBs21OMx3ze8vXO1
JxIbdtu6Uaj6KIALYQZKHPpvbnQfaZLzWZhkS1UygaX5jxQW1q2sAqreatyfNLUVoGkLRQyYd5+p
0bust7OxH7WujsGzeZXD4kHG4a+WeWrlyIIM0oopXVvGRtv0aEg0dIF3G8QO3cbpEbWiAaXGCYUG
wtr9tasI0HaV8dkytwQp3yUVPjz/dxpi04DarHrGeRRoFWxDhvs3UYo8fxa8dl5RaQiG1bwxAY4B
lvGhuG8mqVi+jBwPoD0UW38FDiUsj6b0ZRPXj/i42/x4szOftcuelQ6vFRQUy0p65p0GUldW+5cb
c72fkp3xF3ifyreyYNPpxgNmc1BA4XW+AqX4Zw19GQUVqi6ztXkhhd6I6BHLIz7IUSWUQdFPf0i8
3M9aNNAUqUscD+9Up9MYg1o8+GLQk+7vW1FuxMJSczW5Lqsw7gz9hcdWNbSBzZwKcE2dCfHFPY64
r+GKOUzHJricCsCzmOFF6mhU/BWwH+k7lPvaC9Qc8WgdHbYJTI/edSSPhgH0UJo3pNvBgaHaTAqe
wfJaHe+ClH2b5bGoLGfdVHaoiIpIxYpaG28Bkpc38hwrSaPqQC9MsPc42NPhHFaSykVzMKvyY6dd
JMFrkon7EbDGTCZ5XSPXOHge+lJoZZWLL3rK2DgI/jcytHdtwmzwSUYj3E+n4/1sSKr2Cvmik99u
4feACeGiqE5fc34j/8TN1UC1rl/kylrCUlzii6VO33xP5oVH/8MmbwCQ1cWGhRhC80He3xwibx14
+juA346X6g7USzcVbXaT22pK9MVirZ74sipK8g7Xxbx9bb16/a+6iTaW0J7CaUCJRgT5DNHWfjV2
lxZ8MnshY65Kf0rYnqozcMSd5XrqO05wves37OJ+4rD4lOquDXPmoxihTXrLjxpvLHr4nz/rE8y/
/lJMh8Mgw+rUZZGsA5G57HF6ehUmaG3OvH4cmhAHEMYAiM5qdIBcRNf68m0hqFIHVdSH+bruzQOZ
/Nmkcdcvv8tj76JAY8yl15lSRl0tCI0IBcKGFYovCBAQCJ2Fr7QxyLiYhE/UaibRj1g89H/Ho1cK
m37tfTsYrRoVJ3Txy3TmCOe60R4ETl0asBOqa5xaVEe6eR4Lk8AzlrM1YQdnT/WxLF9VsK4c1Qmr
JkUSNzIPV6QZR+SmtT/bTXaQiOEBw/c+8mDiI76ZJo+iiZ5T84K/FZqhcTPW2GvfnaL7xbcY8Yer
oe3GcEFZBQ2BUt3fKfdEuYNZWmsZCEaD8MTgSVuHqy5hZV9Fst6pOZyeUSCTAhvsaU8VPNtZTS1j
0wFLD6CArtNHS3veSlkMfi3Ly4Io8F4JZ2u64h3byZvRbB2RnnIun6K6SMkQPwIYkqYY7DJa0Sf7
+WGcKEqNkT9c+Cm8SVF7zA9E0iiZm2/VhBLAAshV4Kdc7ti9CzI/PkIpPNKYF2UWhtd+w5b2/gpm
ZwqBEgMJAtxGaKgdkwePd0G2Xrw2GW2q9xlwntkpKXIygqdnJo5SLKG3B1hCG2wOLh8JvIV/nKI4
hqDVYLLsWUJ40d0cZgCGCIFGkLO/ATVO12zQinJf1EQjW0nLVD1gYzu++NQmC+rVcKsWT6R8Xj8h
o/k5SQx7IYGaFsT83EQ9KNtARmgXVHaPDnGVy3/MBO2yDeaU8TLKPfHuzw+JBBm/xZlDcsDbrBRS
QYjUTQEngctEep0gJ96gHlnZwg1FM/8jmfGxbssaKlAJpyR3FlQnMzwZ0fo2Kgdel71GnloQrk87
R3kQ4/ZDaCKj0gFPFhxHZMAC2jJYgbMoJuuHcmsWL1PDMOEV7cD/gOCc8lHp+x7hhJsEhcb4V90K
APp53V9eqolGp7QG5+VTuVXdA6TPChnBygJl/tY6H/l1tOEQS/XGnSOfARk5qumraItb0oQXAaPN
xL9RMBkFURsafK5EhqggKqc1RbUnhd+NyJ2Ht7G6ob0iCWZr6PRgffTNsY1Ib0i78I8GwDeDj9GF
4IXrEOfkvdeXBRaSbcR6t0hP+0wkZX/w87LL71zx0irqrmotOiW6EwvtD8akTjpXhiI8hZktsFy1
g8jDAS5Cbqy7UdpImbDoml8xqZ1g3ZeGIaOl9RM4tXW6qW/BsdT/GhlyR1ydwIPmgNlYupmasf36
8qU5MwOEg2WOFVJxYHOQYKcw4iGGnjV7UvhBn8sl5oMw4btxV566giFVlfnJvUsnaPrMp4DQdDIO
R0YiGcyDuJr3yJUxaX6VBi7E/jbjMnrnWe78EOzb1FELaBXcmJFT6TYak2UpRV9VoOWjlN+hnC4C
MAv4FjNLeOAA4AEW6wRrviJut7fyYkZ9MIPAk4UUDgjeo78/5JshVR/I9QthOVjGBUHZqpbYC8SX
0LcBijZ3DmmHCSY6wrfeU5NoozxBJva0ivdut+KibQMyX7x0pTi4TQK4aeG34+Qfd7OiomwbK3wI
BjZml/kSa1I1IF5Cq1aiIkx27DhX4qm+O58SAJIUyGyrOFmfl2QW/DvNCOlnRzv8fI19Eqbb9RIR
mkCb8oG8/afwUFX8SRLMTs0Rh5+sKz3SsZjxeWTb0sK09Mdy7mpmGW9KnEfL3uJ9L1hQur3q7DgE
PM8SPcr/0i2OCDoh5XNjHuBod34nxs66ZkJDL1rwXsDnj5lHsYEPEQI8NifaDP+sP3dRQpkDOqYE
FNIkJLzzSnC+qyuxYZInpVN2CAxtHWIvB3FkCuigLL87YA80tD+bJqhVs7WphOF/nKhB8y2++2Es
4OJ1yHUa3dqtj6XuJa4N55I/2n7Em15+NZILwmlDqnN1KuWSjHbPWpr6NSEgOpLNj1PwpGX0e9YP
dM1jaHvgY6bSEN6fNxbkYPQ2XbXUbf559fzYd7oouHEfIFK929eZX6Kpbsh+uOSu1M2EauaR+h8D
2L5AgN+JL9WM3VL1hY1Qls65c+grTFOo0+xNFrrVnd0HBJNWzoZGsGb889wC1BLreoSeN+cmPLmp
QWw2LfD7MbKk5byW6qyl/RQMVFhPyn4cgxYxW8v6oBysGNN+hk4XyDx1U3UWQ29LxMIQO7c4MFOn
99MBr3efxHAX7lgg9g56XHLXiyFEtmax6ztZOhG5dFWiPdzLdIEZptqFTGQHJSgWTiRcenAbvNJ/
ZeojefSBpGOO6Ez2ZBI70uoSonf0yl8Oxq+QKUnxLtrplXYiJfVzb3D+UonpgvsnbXiEdo7O4UbW
3KZjUq6VEHaKnrSrmQd9UJnG5vVwF6UbGOqjfVT6IJkRbQH3sMoEvlzMpmJ0G1ZcgwexNFPy8/rG
lZV84P0YqAJVxSnsHZ0RiUx+NwgNGja9vU9hFyaIlvCRmBYdWccl3Sywk9ZG38mj9EfZfWUUW7iA
veRsKwcRxk8Kg1GRV2KQViYfhTOROlS98p3GJK7u2rn7RtdVcRQQxe+cgg2OfHftesRS1kQKMXKR
RTo+NeW8lcHcqiXhtE+PW3jzV9wrvFDDS+Zr2hdszThnwtIy0UrbOQD5InDRd/FRmbc79rRpAvWe
jEMVc9GX+t++S2yP1+BfgcLbc/BKLxYwXrxJeMazyOTXQMUwXfn2I6jWAPk0F1+Vk9AyyVk4sua2
+FiHnxdQKD3/94BgRG1Aybf+OV4iKqt+S8A0ddj3fERuY37IfvGwoGx7x4eqEL09LB/wGD6ajw+S
2iQZ0vDd3NiUmddR86lmizOA67wg2zKtpvq1I9XNCAaVshfEVfdZ9cK/fWZE/7+6q5I+Nqbed/qf
gD0bHPbjn1EXIiRQGQ3l3O2fBiOgQPmy+IYj4WQbOL0CguJD/EMUYKvVC1TsAIbQj4PZTLboDeub
TtGIbt2vOMNT8Fp+sgFhLIHWdwSmof/cMUfwIY4StBEU4ZYmFphfxzL+rjJJppNafLnykRSGDk5m
XaQIVQAMev9zDLjymw0JCsfiDTbXhTYIS2426l0vSHXlC/MeV/o3Cz2cIiGHIGfTErVzTBse98qs
AgY+l27bKyF9FmJIXOB83x5vzfkPBO9LdjX1LOXoPUIBEur8eEz4fstUGR5Ub08Fld9kIllM5JCY
C/UdYIr+RBK381NgeWhIyyj4Nj96NqhqkdfAdF9CmYia6mfvoc/Q/46MxlvT5ZnqtrU4KUDF2Er6
xCAfazlMUth5nglW6mT2VVPAD5/QlGcz+0VrG/2tZ9HWaLZ5YTcSjls6ZUssaZOCTYZ4e6bKgqzJ
RjUox318v+CeM47vkfJwJX9A/F4imuNF/T/E1f4khCtauD8RJ3Ivc2gONthMBaLxY4OvZU7nacAN
/eJ9RgSF33cR4GNefUBKqw7mLTg1xeHoGgw0451Ns/nzrUapRMg6NLoWx/d/uWZcbXTdZx4o/t2K
DzAEpIbyE0Uz36/Ovf5WtCyPR4qeDOXlgKW1s7hRIMq8XnGD8uBchE8K/eetQSxYK36Q0T6ps0Fa
gPr1bw+xfax8AzaXTxz665FasMdJTE49fpPYxeGPT/1o2mX8n3aqXu0K0bn0Afmh6j7FGKZ6H7/5
d/UEy2eMry8ZqYt367fsA/lgmSSXkPypONAz7aqWx6unqtxOhyLNc+uTMKwyNgr60Uha4I+FDEUL
uszi+/Qyba2vaXlf3ODsV9f5lcnM6YJwrD9zdtFdwV226VdOCxqBvbi+/JaPk3HyqNBQQ2+D0/Nu
6qtZJe8iW+cKNfqANAf50WvfrZDBV55ZWE6CcTAZpJ+OO7DCunbddP8v3csBuuhBVku7rQf9sfWf
zPBUZkIn744QNPQ56ROM9fdmCEDCLkzdAKJ+Mb5b5lls+8hIqPI/pXdmBsZYBgnmqIh5yQe9I8WQ
A74g/4NLfTKalxjH2cAgqJwvduWNOh8Kaby9dzIys10iVgHgDY2fsxPaAYjFCEVUBVpZlRAyDxJf
pxg6p8uXtUB1b8zQliTtCBLZGiILnOc9F/aUXXHVvef4sbtOSquNG5PYcAjv0tdFKWbv3cVlkTnE
0AQZLVmLlWG0SIfhsNteEPWVmFyQI1pzkpPy7/BFIHVkaKnn1eM9tK6zFHknOISDJTCnCKuYn3Zj
VVwFa1Zthp+D1Jiq4sY4NWMFr4+XqWj/qm90MNW1fwfyH8YkiGxcuOMRZvTxjdGXGJ04stE27r3c
LkeqGsVk1aQzwwQYlHJ6s9U24Ymf8EWNi+Vy80jEIdpNABxl8qRL/pWej4anR2s2VoIE0PCDKvu/
wTT+4LH3L5EGxiDUyJeR/TN8YKApvokcBCJlzvPTOB5fy+PFp2Pe4VdTMFXrXTWOuHhXG6L1oxYk
ut1dmcaspL3wKDXgL4TKBr7YanAIsh3tGCyQl0KI6NvlAWCvb839HsEBWQ3n1OfUwvtDi29VXRbG
nkBp7PS/L5YUrGH4GBJ1l84Cd0nNJZpMM8jG+nA39H+6ZNgwMnxuXYMlmMPbEhbQbAzER7hCc3su
wkrm+BhYBNZFHMEQMY4MZ5Y+3y1A0q8nC/kOvhWOfMMpfk6/N9cuzSUtZaSSqLuTxWQruEDRRy7i
1A1hEeIgsggvA6aUXvkh1Z1m24HiQ0GiUOiNUwES+R6wKxaWTEfx/fhbZiuaiPHoHxApGXgGEWL4
sHC7o9VaWDqIsf201Xb5mgJBAdoExtGBMzI0e1O8dJ8rBSUV9zNnxb9wk6BIHc6ObDb04Zuvoz6f
QJ4pyqKQysITvYMaV4+h3Z3qPfpbDiq1XHAW5uDvbHNGDPmpH3/hHtpakBcJjt5r9OUTLftj6q0A
/DepeDYoNEec/K1JgSxlWg+kZtZ9PnlcdZ6ZbaeQ0ffrjcbTLvDdGU2Lw7vROc8mmKz1aijJAj+u
/O6lYlbFMYZzFRETaqSHIzWSHNqW2ombVMwKyrCYSKVF+ML8icVJUXgs4HEozW/rVc/HMpbkltWF
j2lmWkL1Z/CuH/+aiqy6k+NUzZVBLHEJ3FND+MqZYIvHsqjWQ+aLhHfDafBZU3YRVFpvqEEl0SJF
pCKcPGr1Qz8Z98wq3fJX9D31HpLJHsnJK9s2uk+08qX5a5utwaeDfingNg/G/7HAMHnlfYa2nsSY
tSP8MFy0Gi9ng8PpEI/l9qNi71OM9PCcPXYsSQw5LWOCJ4Xk7kVtEn8kby9jKqAyzhYm8XRRPSUH
16F/XxubBQ2yByhRnz+9rwQyksd5KkTLhA+fE9u7b3MKj3xYsCScsdHJ7dQ8nBC3gfHEKD6SMdkA
Be0vixqpSJn5b1DWZre6UCKyVFEzUlUg+df5LHLHZxS/kp9akbHoa91yJ8gNno78Hv/pK5m5AkX7
ELT4EkOs8U242O2pQHFy7ph1Sts7Nnks70cIROvXEtvJv45a8cRlSbpyO8lyXm/1iteDjqfwpYEg
Xi82TjDW/gUmIJC9cMfsjL+yq2xtFb4r66CT56Mfb+bn2MCaLQ9ObF19gCGEBmVm32ENgaMzomHt
fmvLFhBEMyrRvGGPvncjwcwbz8DCpQLSE6Je7n5aaPa5Bd+YyjlNNkLNudbSMxqzjerFY+n4H5QL
s8IN6ujKZlv6hUNPOMBTGQuyV2v8U1qaZmvFQlYfRCrBnO0LCSjNY/qZeI+QkMYOo5viHnzWzpuc
R4vBUtn5WyNb9lho/ILZApY3+9iieaVMcJB74bo11Z9/gP7wCNHhiVBC4q3lQxKnoRs351Aw4AHa
35J7FGmoRiFxwhpnxz24+2FFeyvlIa+YadLyPH/VepaKKTpIqQdO8j9IMfEbONpbZWoHQJxAzuZT
ZqCUJZkuaa2l/X1ePj29TMxWAG+SrfHJto/LeKWPffhFJp+cV/HggOPuEPQzsipAvULFYXYjCPUy
tw7RrhMKT2Vs8bxqzyiRblPyOmIPRo+FkmWR49ZMzMNcPIlU5EvCu5TEQsQyXl+w94tdNfQmHak7
V0QSuiTZAunAnu4mOS8rBU/me2NncWclhtOEbAubwaBWMaQWAr/6dt7AmAgklkTg8a93KG7FPHQp
wY0WhZMHPPAGSJnffgLciCxN5YB2AbgpI1870FFoSX09WdoRlyWj8pQagPnQrpE7SKAJduOZvmnl
eEBVbi9vxrOnTHMsPyci8vaFgZJXPhWX7o3/iOAFro4Mp+dVlBgpaDxV14RiC8+ynzWSnTw8v9PX
RwUwgZued4kPIIXIrh2uBWp/CQLjCzLqJWQPjljf5ZAME8viUpfSy9odC3PZGKBUj5gkgzQ19/rX
cnjehsfzp6PIthEUKri75KoNQyy6GhR0pfBX3gPs3+AgY+Hn1c/Dtx8rJc27VpXaikXsUJqw2OM3
DUmKLOkUoqOotqdAQLoAy6/CwKwvKemuGDdPyySRqoWwIcG3yisCrtK2Mr9Zs9K9x2jpbzL282rF
/GopVkBGWI/ZnJiXQJlFqjJQDrCfR2rOKlKEclADNaV0WbfVQn/W7/GJBryZdbiUR8fkpaTv8sFw
Fpt8im8o+hJn3DWlGCuA9WoqapdOSTPYJsMC7g6mZx+XXRg59qEl/MQ4UUs0uW1KZTvJPH80tmjb
04Ff5pRyL4h67+s2lfbYgG/gbRIeYiPe5cGO62gjSsk1LHe7pG2Hr2SFStSzyhwVmIjRbRteIBLj
vvoYUHCPqzpyoj4Wy/kOfcUu7eIrcGIxnF8mgBZgZIdDG1rm6rDkbct0hw9DeivKUClfYDg7bfAb
T1+EnwNPZ+o+U47Lr3gqYMV+LSk7GmfxFnN+B5PEuGikWsMcQPtm/pNPW140/foX6Wt70wSZmnkO
49w9kZhpm94cLhVk0g/SQYhiD73DZ/GhqFZY6w4AyY/k/SfKBAxhenhAH64hHSaH8RIWuQyhHCVC
EtM8A5HPOop0A4FSxQu9y6sn3fiqzOD9hUZxDfwvBtdd36sTfLI/+In7h8xcCwkOIVhM5utzx+3h
0ht3RaZ+RPphUNOs/rqh7gtenybKnE2z8UKhmTHjWZwA2CLcRl7lDp+lHFAM6fPXSUkVz4eV9uvS
XbLrhgVZourNikhNyHMSlmx0qJSvUOravoSe9deEatR1/tIltqpLfZWK4lSX04lT9lWuR1YDvyS7
+U+KNOyh++5t5k95Prs5T3puJBF4KY9Ijn5hsYgwZiAvG4fBqiQAOtw8opn6bGYN8pBT44Bcs+XS
lIuA6CES5tYQx0XeQU4xB5h9HKJnL4dnt0iAv+5l5A2+oeoX38ajUXGI1rEe3Hz0IXgzlFL1TQ9x
kXo+LEYpwedMqwsDP/fU+3kNcvDmLNuYSwoDOCbsHoYkplYwx2l2drQhqgVJVUaw6BXNo9pZ4n1a
VaiTh+l00V8Y5vFfXJlkxjfS+0kvm7Xx/GYkrY26uNls2reaTWg5vBUiQ6hBJ9fetD9UfkfT2+qx
hTAH/m8kquQ52jBV+H7UFyGqJ58K/xfH8T48c56VY19Riq0GZXBcv/JCI40dgM1dhSZE+1kWm5+Z
I+7LZe1sjuOhfjCO/jwB4xTjCYbxfdEJcjQGJjp13xI1UHRV5krvlSUoiXOE2cnwtreoq55xkADw
3qkGNBAtQCP8yLcPukaVwuWh5x+LeNKzSaYXhr1KCF8iwvuxC3KsMOclxs+I2keNh0jewKRwPomd
SSil3A9eKYG1jAGlyeSZ/MqSew03qR7VEKsH3qEwQH/KntOhMq8vt1zJjK9nRS24pX8auvr+sonE
TDcKPj9MeSnmrnQIGrhrJyMi+4+2Q+ZYKKeU1QV7nKJ1YxohIaXfFBh+EGNEoIq2QNjEwZREJqgb
NUuRYeuwkefEWUyFwQDcY/OLMuLT9yfEscsVOIM4Uzvu4Farxbdm9p8OH9nFNu5bh1v3O5C2zGBn
7sXpPUH+k+RB1EiJkqOdMBXbg7xqkKX6Fecv5ksmYVsQFKNY/9j57euguCOvN5yeqq8/jnU8HNFD
E3beGjAncApT9Y63g/BjlacpD//f0RV9BIEXh72LbguYcfHlXNhQ8GsZqMSw9X6sRHI56P3LQZe/
yo9cinBcVR+ZLATvsPx5Iri+AhLAwEvh6WzAO6gm4Xid86HOdgsuifszeuMwpsnhDXTIA1m3Qomp
+Ufx2qDGj6EVZeD9UUCVqpi5A5fmxvzZjUdxcF85Qpbx7B5EMzfeZThz/K+GjjRCy5W6xdWWs80Q
upX260kk4xIhJ0C+0cNqGmHqBy0cfwi721I8S9FBXAw+EJF8q/pDahu4p03N8AM7gqbJWtXla74s
11JxZ3Khn9wSZpWbYrVbBtu32xr3bFjGHFIGYIKMSyzIPPTKdOrnghiAWWpNa8nxdRvk2etUVzNu
OPnM31DxgQEjqfmGzGFo8zg1lavOWf4MjQdGSmOEtNW30DE9M9B4aBXEH195vonRyVY3pZentEIC
SxK5vLrIg5eiPynVkR6lswUKurovRIQRdUafmBj9v1Q8KvVJ5swraeVynwuOC8fxdkRYxHhXnljN
IibslhkaMRsiM5vjAmMDKzNt3k1+40qFuoeskuH2f9zpX0JW2vxRctDOyydRUssgwjtxuYAJ+9YZ
4xliIGs6odeueLt0wEGSUEODBcpdOmbME1QGAABqI+LNklInJ6f+swgfw3sZ0AFOjcrupRxR2F/g
YWRyEXmLvptJxXdQcbZjIagCMVgzLRl5CRKfgi5siNvSLR85UhR7MIbVGfV1Pw51/2fMXM/Qnjm7
6LfSzM9ZGK4urYHfoDfgSvGK3DzfZjt8R0LooDYXacROW2667G5qYex1Ajk6oBJ44OocS0T6SKuk
rWyzkHNuQ1LCa4JOiNtYKSw1adtPl5PmBaExC66mUY81wgLzb9lhqJNq4sT512V7bychRHH70pZC
edNO4M2GRNt8N6le9o7aAhAy58OYAetLuGVqeK/ap0V4emyps02Hd5mtBanNXJKnlb0dVmActVRH
Maaj1mhpTjy6n7BNSgGQJrGjDHd/rgABietZ7KSDC9PQjDVcUchLAIow6aSbptjmHgaip7HZWpf2
t8Q0wEo/hF5oAdi8MV+jT43bX9oh/8k2x+N4fuYl/DMT49oNXJAcz4XKrriJ/1r32kkpVZzubvFb
wpcLXRCf1fRI0TlOCUQpuvXco+R1lkU1OGQKj4HqKsByN4t5JfoOrSOl3/GYnyeN9Rs5bE6bNHRY
hsJsQ85DGGpGxQ+H3Yi+6SSeah76s05fP+7KponwNw9y/07vafNXphiwKJ94AnSflo8EEWQKDZbZ
xsTqSHlPjJtZNPWgFwZ5LytupFXlbzxvJl5OYTnE66yfbY1X4S+KPUyDMK5n9M7CGIV1aUFdtcY3
HLIXnHafxFnrLlRynbQj075tNbfI1gcS8NjbR4BAgAupd1YPcAHZcJXXqazNIZa/G3LdR7HP0Qfc
8jysmVnOPfr11cetW35T+pH2SGZFjW6sgOUk8WA50ZpWp02HyngqZywyKIVi/Ut6ft9/B9Gmwfka
xE3kGVBTxY5JWd/y+3LLfUBAcG3Hpvpq8I15oLY5WLGhHyCKQj7+hn0C2yyYYG1dMUOVXwFIw8W9
9eP1ffVDfCucjsYLy2iIgR9W1jl3w/6SSrq6s7Msv5XbH39pV5o8T7R7l8fFTWKBg4fRjnaEQ5Z2
tgSE7kIU5+BorrJzBU1UOFkALzAC5zhQiZe5xw9YO4ZNwCWbw+0lx42yFBFXvmuihO1WxTmfcE7j
Rs0py2L0c54nwfOEv2bnpy6tz6N67veQvi9nzkndCJMAY9sue6LkIH//0UDNDrhAc+bpWknBgYee
IEf4elYBB5FcYZ9c9q34SMOHMNpz83pH7o5i8CUKWS2Uc5h4XtDiTP9LrjP9BAftJWtYE2GmSWBe
HDDGgMfQrfMKh//VtA18DIqrj5K+8MPp4Yv4J6fMafHUaCuDiF4nieNQMCMT6mmiGhKUsFi3vVoi
CWObpovY+Tudn52qc9sASqQHKHEEfN7Qn6ybLo9RZ9IL0BEHsNBqojojpEQUi48umwhkHgXxPMLG
GkAuvD0RQ2ZKFsj5VHFSLQXNsq/e12ULF8BIzFAPm5RWvsEzhzBRBGT31Besje2FgNUy0XHZ3Jlc
Ev6BeoeYx7e7IuFhQ403rbF5B8kid9iISYYPsZ0nbi8syG/QBge/B2P4YKtV3Si/NCsde3DVbLro
YZDfOBWcW2BiZ/OnCPlCLNeFuM/IRsEDRt3fOG6DQxgDZ6FJmqaKasJLeQccMWpFxJFg3Ar+1FWL
635OO2bOtl/+bLav4ryCfkoQcELHipEOmxy9jepGTIIYD5ze3ZiOPqreUPtRco1P+IocHJsMrBZz
/6olE//uykC6vMzErIz7Cqd4N0QP0FatdZq9YjC9WvEUlkF7Dpk0zFPY/8fAJ4RgAUW8gatnL8Jj
LfTQGfmqJ0+fds7BblR58F7Fo57vMMh2nSAdiULeSjwW+kaYYTYI9bANTSO8WL2MqoO3/wuA6+QA
Foj/ezkWm1I6Ju1nZxr4orhg21TmM7zEgXo+YoG0gJuSTO41VzFr45gmCiXCfqy4qoE05etdnI8o
y96JaEwQbQ+m5gTn/ZrcOiAXiR6xcxYOdRLWVCyBq80BMWGcGfULQRQ1MiTCnomvmW6t98/SfQPI
7XBK2PfKvPEVc3I1VHyIlOua6jlUEsqHpnynUa9xgVt3bukyfmDjGsTPremAHbPOOHa/7u2eovdd
v7P2jDo/0yx540BPqUqwzlI8gzLF8SznVT+pbY0KoYbWIe5kvfZXCpI3dK2tiEuxO7fMXbctngtw
e6UAykF/MnE2eWy7D0wv8hsQ935RHpyY4gBfOqqRAdn89y0bggkV2GpzG4WWMpg1ZOhFenC6qqle
vMNbDNYqttuPPkl/gr/xSirWMroHVvzcoh7id1CNFLpRGR46+xRwPgqe6T8BfMPwYVdD/CQA7JMZ
KH0XOJcpz73vz0zNEZW7jAWyXZrcpHetAPEgOhipA3PoaEiEpJ8OURf29f96fDZvwaQdbs+saLTi
gZfV+Q8vlkJ+v1aK7Ay5wv+UBTqK9/hMSqs+4HLzxhwziOiy9pAZHCamET+/Z0lxHGvnVmr5lV5z
5Pj3ReaP3vO7ONaws3iIxFoI68aqpx3pDkWwlIFQmsq1k+XIGKuasTFUHlFMd9Ud3BpMcra0qKin
W9YYRlvBVXsucJFS67f0SBtKCHbR1E1PnSnXLeXx20uk62Ywphuo7lEBVkNmwMzZ/pcXQuEobNXA
BHA6BjA1MQOIkTTrfCp6yDWYz/3rtk21Cba9ZiNYB4fvUZQt5myNry40Q1jc2DLyZpfOE/uaH083
tBw4XW0ozjLN2deY70bjRi1FeMK2fl4jJTS+AUGQZ3AbbT0Nq4nTb+W6cIoS9t9kA5RF90ZeG02c
Rg6200tr/3OD14FkyYK2X7AyHssL4FeeNoq3YN0N6J4k4MTZ61N2o3+mJoXipUuj90SKdX0rKrCl
FRwVOfjS05GUT5DupjrLPUCz5wXJDNkxnSrEHmBnE6iLp5YmshSXiPyW27tqcj47ZqY98ADw9bDs
H3ieyzeHpiOj28RXaeW7TYv1iFqhaet4bpazM3cDdJSoYC9Kde/zHEzZKDleCxZ/cOmgtJowC5aV
/GH+eobWbD1h53Bkxn7ffdnO1/1eSKsDR9jDrodpFNumVj77It2Iy2DDw31amc7RNZCeNwjdp57c
kvlgAsEcN2Pm1n3SML3g46SLMWk8odSb7E2ATu/WAYe0M19JGHbq8H+ynBYcjiHAnViWQBORbSVp
P3//QNBGmCBEmyt2idY/DKOGWur52cUKZp5UsXGHNiQfBhrG2RyVfDMoFo5dmeHJxg+i0X9BerGw
gSgY4FZ10Y7F3T5sSwMzuWsEcN8Pz26nY7nHjQp8gT3O1Rg4u5dJAh0eK9+j2sCJjF+M96SMaJcF
lpKi8ZIbqKmgKVu+gTjnGI7R5HtTjLfr4tPZ52LdqCau6A2s6HJ5jG4qkJPGPBtuOYkV0yy0Accu
UCs7F0NEZO/9YRVIVPPZXOMEVUNBZShuJIi/ouOjJsiuzjGSlvnr9yTOXomGOYL+vnNjAtK7Qu6N
tuK4RgYA27Mr3sCUoPeR/iLOB/Ty4yj+kPNQ1IVeENHkQmuGpaq8+ZmVWb9mAZraMm+0O4mKPwkM
+TCR+5fyx656AIgU89EDpg/aF9Up3Wh8w3O8BSksBjqJiLuI3vTew0QObmGCIWjVm1mFd6oSwFdy
9n7LxZ0+JmtvtFfzeqfROuYVU4MVpKDzNbFk8+z1/+ymHkRXl5hu2iWTPr4297g3Q1H0NNxnQRDi
wo9UCCE/uKWNwIC93HJxDjrodR1aOOiG/Wyk/SKPX3KJBFT860ZuMy/PphFYE0OcMxk2zbbukTLa
mpNdIvVGmmWe4o1g0ZTxMN9WU1EHWooG8HRrPIwtphQsLH5XFjWrlq0yVAy7VfyEYzsT4smB9UQB
8Qw5krni0kR4gYj6d2nXbEywk4YoxoosRF1pkeBL5dSF2xMVVE7dQ1B0q75uHRuEBSOcx28FaYav
H4On6TyM9YXO3PQHfJ7KbMFB6sUUWFjMIcjWX7RjeyeRqpM8XcYxLUjUF5+NIDn1tF+d96f1m5NH
/hM0yyXeLlmEZev3+Ak8i/yDT49K6JM2cgL31Exzc3uLOc5m5Xr+6FUqJcO/kBl4m7jpQ++J/JIe
I1ZXgvC6dzhMuo23z3reGg+DEX7g9dSCQ/vmgv0sNA91V4Nj6HaqopzzjDTBHQtqdwQAUxSMND37
ix+sRZOrcqhIqpnFYtNm0tC1+FET23v2SOonm8ywzNo4XzI62SxFLqHm1+Fk0sYLTKDfYFT0V8Bb
ysuYLSGknqC2keLODS28l7iWrEG6z1bIhdi/hgBAyVCWr+Cjj3gVOEceaAWmvPR9Z9yysUe4K8eX
JyKbdcqg0VI7Fi14pdXEDJSIgwBkSneGZzt9LAoFVhcU7aAZlk/PRXRz0DjaD8HguI7RXvTOWzEE
nfDMSqffoYfdqlcW2SWswhHRK8aHhN0rhptQSy2v4lyufAi3q+nregd/I8UCaDdR0laLeIguBPHS
c9znrYfKhoyOZ8+d9dDRqquvLe5favjiGZiuZUtWyivSzoCH0nqefMnf4R4yNbm8hTca+m178uvF
3LjAC+ssUc77Z+w0yXODuLMfMpFDOM8Iyw8lTBSyXmhLwll+1xEaZX8DgQmtp3812hOcgQZ0WS5n
u47vfbNFi7dnwAwz8Yf5bVTFe1dCIN44PWDAr6UgapKaG7w1Zcc/YeRQHqkIL7VxTEyfNLmyecBd
cCNhluXjPGIrKKvM1uB1u5EBlusjN8IT2MwxX2FexfdwzHatkTyd1MKAvPuGChCQoC3sr0t9noDE
RZ2gRAnLPXFjdWGEvDBzGLgZO3njlp4H01gCtPhCoIqgTVfdqRripcCJpYvLn0dR2bVfhjyRg0Kj
sjqVxSWLJeyB6M5tH2Lv0m/lfW1NFYqKtVZyXHhMHphZWdsIPQ2or3F9DgPENoAzZqbvuKaZKwUU
gk5Lere+Y/QY6HnaaVB6hUEQq6MVs9qdgnWYQeS1hVb+wG0CZStyEER6//hT95+qzdqGd0s8JLpq
UFKzQOJ9jwWTjYie8FWp3GCEpVdXucZsTWNED0nFWSrg4HpovtH/qmHOCvmXfJhWFcFL7kVwXZbj
t+0ifycX6HNhUpd0+MLg0+gaaKYj0w0XCQEXd9kuiz38eMomLjW4P/E/j9rhLvkI0ORZCm1sKGqF
E/NM7yKAWvRN9BCH4l4eZnzU+0Tmuo1mmGg4QyIguhqZDUznw4ZSODIR1TcNTM7AS71nmjZFZKEL
JDf2x5Uo/2YL1Fflj8j5Bd+Wko0IVZZLq7PgGOgsSnQgv1XNMyu+reFfzx9KWmBXOkAHFsZSC68B
re6aadDK0mjHY/MhCSIQMF/vP8UMjNP3y69eBLV4qKeTVG6ufVfNaLk11jJw3h5eIyrBJglwINd0
ieKCFIo1I5ld85yRhQDl+gZ7kyOkKbAB1jkqdw5L4I40ffQDXsBp8SPVYCg0REoV0Ulkwea7CL3a
19U9nx7pJ/QB2OSek3RafxEWeMP0yHkLNHomoEobVFAP7Sq1QYooo3PS0SURRX00i2zU6wCav2HY
dCq4Hyg+D5pOxENT2ZzWeqB21RDn9jWzWpQcUMCr/KIS+J0mcqn1KOXiYZJuWfsPlr1fMXL3Mfrg
ivhcYSa9DHddiuuCKUIU0hZGCTXSb9FVyGJkH0vgMZ0JeNFN8gVSgMKU0YXGEwOf2PZ/PmiKvQLi
th8Pta7lzrh8kf9Kc17pKMuUHWbZBA9fz+49WrSHk6sYWVle+CHu3ic2UfWc+DqYlOXajSKQeu2a
zlAmURpnlGB28MdzZJiM/n1V4s66hdy3IYolVnqWIBntUwZYr514BfZ8VuRB9C6mjGEfYtmLAcZE
d1+G60GmX+Og0ZOWUu+Kd15yTNkVBkjRJysKM9lphw7rLqSQd7ZxHDXJS3Td9eYaGJW5XtuNXn+1
QYYCjls6rNefGCa5IPgHVW7sRmvYwHCRXjjgw6Q6pK9PWWVlJyQzjIwanJJwpHMuH074m1o+7JZy
bQkSmfPHHL7FmeN8fEqGiUF8XUSuq2dbD0Ixi46GRpJUx+OezqBJyCLLSw/nmwO/CoaVTwJxwKwe
04aqjTDeSjeHoJRwlzdJ0dtmt6zTMF55XjW4YySgW6Z2GJPgnF/0HXJOEVAM13Q0HW/d687wcyS+
LlLAVZr+fd1Tt4D12wJVlwhI4/W6nCcXf8p1hEC35pqHymHSary/Z3BPUzMK0vQbTv/afo2vdzwM
n3fhlV/kf7Ohbvi9YU1XeclDiTaIOzir9kNsYdG5BevJY3iCEcaw5Y8OX4eCJ3BJfVAbz1pwbD9z
AFgHF2u6QoMbTohQ/ORY/eWNCGrkO5tBBy5gQmnZS6CzjEGVmpnEtEuhYLmte+7+sP6W09EImgkn
XxBNgDV7oZSuT6icAvUtZdKr/pwB+soGvdvGwLCRMH6XHW85LTjmNYnhVRsCdfa7VWBqbcadlhNZ
+li3R3nGyjxlatF9ZCyrl94WmtSp2Scrux848Tkh/Y/mchd5RflkmTXD4CDa0h87w5FetLoUOyRz
vvctSGBnbfmUEoXKP5jsXV2PsP31IrHcmFbBICYq1ZcPpQna623R7TTpEhmUvoam+c10/N5S6h5C
nnIMiDg+E3prYzjlx0SzXKTykcSHcuSTirk5QMqzhhEFATyBPMLoGBG94Fx5NbpHVkyt3d+2El/+
1I+2PmKghm5JuQSdCiRzk6lTLdaNiwKuMJ+OzV4PYf7VJNqUyg1CNtv9ZFaY0t1/l0wKPNSjbzhy
8jiCpbkHMLKz6zU/2AJF1pczvkgS0349+28Lde0WS2ZUmp9M3zhD9THWCdFgw30qezd3/fR/WIou
0pEKzhr/98DvG/lcHeJTgrG5DQE2K0zep9uMN6tdnFcZ6u2uL3NqKel3FfGr8TIH4eFJ/amlyskG
Pe/Qnhjm6zRd7dkIitV1m1bitBNLwWUKCN2eL/mHaceqh7ds1GzU5klCJEdBKqxb+Yg2syjWnema
DaGaf7dvAjGU43hI+vzyhTdmGaM6iWOrbYDmN7qNlVfC/Z52H9JpedOpMCzAOm2hGDCPgPEos+yU
fPbO5e0zpAw2AGjynNrZRasMWB4BAZ5gPPSIAim+YvjAO46cASrDm2XtnPyWF4EdQeDzOHctnSUR
spBVZ8+s45UtnaNfM1s+AA1dnBS233WJ4fVJ9bTPS/xgf6v4b2ZniqUedd5AVNzqKxrj25Z4rXYN
G3UR9ZsmSRi3hQjWtCE+mCr4GGKMZdKwYw+L8iulmGZPlJHZz9Ku48vYA/Nkxodmfs87ibJG4GdP
YITpDX+EDa4Idy8yHdP2Jk4JhyfEyVl+Ue+r8GxFEeaQ6fg5HqMUFUC3gUEZ0N0C2uqpF/X5sXBF
wzuPcpCIg5lCczZdW/FD1M/00o2d6qiKE/soPnxdYzj7FsQaDnLZzsUKi0xh+Ivi7VQQUAaeMU+h
ldzNFTAg3bmJgi5jKcOgzPE1T1xXu1W80N0Fs0ljytHas311fWIG6j8L0MgijD0Y1qJiVfc7v/O3
pQIYzQ6fB2Odg1LTocSAIhDLX3gojOO7MhVctPPbkGG14JOm3SU/x5W2Br+sGHEC7C3Mh6D52k3R
WEqsR21oExyYTOCjkjMY8OXyxy3n4DecL1sGG+2qHmMl0X+AFIp35Z3/PMX6KKwev0t5CW6NloV6
1MmQk6ICojzRA14NcVWD3lGwm0Vh9y3kxPVpmvWnPuVle9E/bnsZXe0yKYGzPCcNlmcragzoi7sU
/YOgiRUBfxMWhbxHXFhtMyL2mnGDR1Z/qKuWYOvcaIKiwftp1ECaE9t5uBpdGi1tTsJJkEjKIDCf
ihCtDwnnyUYM7vKnQBPMy8mrDUbIWGcBVsRCIzGPo2xPqt3s0Cg4M36Be0SXV1gGBjOOHsL2y3eu
0cmq1cjIIYoRu0sWUHQG12WsSqGkdq1eYzdjT60oktmRoi+ZyLxlBgt9z1G3wy6vL+joTLt9h8U+
56M4xF39A7pm5DYSS7m+6b+bGZaNiemFm9anrLCzR4Uko8GU/ZV4/YZymy9O4k8c1+iFry0o4C9R
HN7YlS9/9wr11lpxlz1EUNmVIBebdD9HGUlvXioknDPMcQOwxDcxs7aoqDS+lZGF5SZIcNnCIQWY
mqgGC25YpGsOtNG7VuM06+FqFSVGMqeXZ7HyBzZePw+ZEy7Wceaj/atVECmSQZYNjTb47UPF6Aaz
1tOHPdrJMLZ3G+nhRu5F2WP00EOBgTrH2CoXgu8RH+WQqfZbdzHKHfzu8ApOgNebjCay42vTT94c
Y6/nny9h+WL9Twz6j6rBYYto7mebOQJHHKEQMFEgvqb1k+UxQhkFcb80HRa1Ho+AMZFOKQSYGa7v
8Ur7k9v/9og0VzoBBp7uFql6YI01LwrgY/wjPqmNi8H4aYw7zXEUxXVX/jk8wE7oW+dpjR0gKwN9
OTeKQpNP3amJl39o0W9FGaOo8+7tdCflEdY0AqPdx8WF1Ue8YJ7prItfA0RC+PSb0CeGMj9UucLR
hUkUPRueRfOS0wUPFp9CsGB8PyIaW7bomryjIKczQqpOvbpTei6rXRehvsl9g7KoVri/4vEohxH5
kYtD1bPY2duoUYQl+eDMj8fl5ZoPg8w0BqK6llKYDeZA6rIpidJ4ctssKUxL8MA8S8Uja5xPYoFX
sKZCN3IPGhKNcLmmGDGyNZU2ZPQG6UGwtP/buPMVwJdrdw7iHNpUbRHwDfRcVMlyfrztt4zR4DrX
58CqqWx1hGkPBemhM6dhQMGZup5dTTy6qo2qJpHyI0Uw7sYklqCNiJkwXVp5JBm5xUHzq9+mHzoi
8XHAZ3Po3C5CJoq7bWjFqNiGWKbSqP0FL/3COk+XatxyWe3OaSKrGPnnAtgF1mZ6FzXAMBQgeanr
FEB5mpnBdHazdenchxZ8uuLP9i3ABhlGcdLRSWU7mhS+pFy6hCPtx99EP33hckfeTUp0mJyZs0iu
Dd3OXBl9+rwk2Y0vG5gQvCGuiWEpTilu/D2x0CQSHw2+dI8va75HYQVbMJuAqLOdwwdXhwBamuE7
dWZlYNvIGcp32s3RCqDuO7sL0wWEm3XXSrxlrK+zRCz1bi27Z5dx8gqbJdTCfaALVVsiQhvBEG+p
+okqKkaZbThFPZ5wwzsliJ0wGR91VMNFHEcsDE1dAvuvc3zW5EzjCIMrz5w930Ex1JQIyaprJeUe
ed9nq8At6vVc6kvicnPDBhoi0WXzNwn5rjPBU6/6pDdM5O54QjcCDfe7wYGHnNl/Z8QuVh9mp5M/
ZTl5HkVvojnjzfGnHq8u/49wGl95pujCYbKPbm6cCWtbs7bJt36eUDjzno2ZbpxxRJRrWf5MsBM3
oSxwTjCbWwOG+5JnDvANaC9441LL3rD5z6N0uUrh2ynojvozpAjL9s2LK6Rec8ZG4qR7IjvjSCa7
YJul9Nfh9U3B5MnOtZc58FnbXFEVS90cHn1AHbUrdbiZ6n9roCiFoZCkgxIKxaT4DCk8nwB1aBqG
xUjW4qDP+4PYuIM2lYzlvfN7U7Ux2ynNqyZ9j/JGqQDgqp22lOsbCnaReVXQCfKX9M1hvIRTtjDL
FvUTC5LYTmOC56HJyk7pRFj9YwKtuNB12fxJikiYWpyjUWd89PEgRmURQVERd7FXuOEiFHqnFvjW
MJ0RuxckxTKAgpLDsKH99a4evDRJcA38NUEDBUwOvezBk9KsffNnZYU3a+byghTT6Xv/yH7DN8FI
y3ET+IUJPA80xDIQVz6PWEklGjpA7ZwtasejEUSJdVSiatrY+/8UBj3YVX4dqy6nYQKmaDDSpfh0
6shxPum5Rc6JnHbHUcc9C0tt21fuvw4LCCMdcErpUqOJDuPeK4LBXLwqxTwJFFkUquwV4AyNqDp7
rVbtcCdY/kPRkz6Qs12P/rsYXH1l1prNuXiaotSDMzNq+/JORkK2otwChoUOZ73sG4MuRqneoCTL
28ZGfHVDj0a22hy2jma/O1WePAiERjfknQLzVsYbAUsHjSSocdtZJ8SPj+0onc3UAT/hnH0GlzHk
MFwPRzqp8wIb1fpBbfMfc9dNQz3IO+aOC5YAlrNoty82Rd8U6ON3LXv6kTM6p294naJjljHO5pom
VZW/dhaPs/w2XnS0GEyRnYnmi/IE6q3+WR14aJdqn1XgJpGDj/V/b70riBZTfaRRZDVl8Zr8KeGe
ub+sPYsyo2QtX1GICnpBby4DIvsyf1Ye+OnU2k+IslKN7j8DyxD4NTPAlKe/5qiVnh/NX4MwYlOb
L5kErx7dbZt7e9fy/HKOJ9tPDogMmcMhlmSBe+5WoKz5Kk/DDUzs7yGFuohuBeCQXiAfGJ3lzXXj
SkPd2OW1I+SrnOoNrYpYeqf5UbHr2c+Ahd9NDg0aVkUbSkXO4BaMA0jGUdogkPo1ehO3q+Ll19r2
wKT5P0iP2oKZh32G9hldHxYAWKc3NLBnogrX6y0424qD9USnhstzdQWQkafzbgr9Fs0hNHwfao3q
flxGEeZi2JKKn9XCcCWBv6WypctqA6qQiLlYxmvtuFcwuad9u8Wum3typdNLtfvVqVHLt+Dnu+Wr
Al5/aGR0FmjJrzRjm0lLoQCwaSgAs4TCXai7B3vDbF3ol5FO7XfQLj7mqKxPCtKqJ1GD7ARPxrjl
HDPxSZutEKNOteAS9nS65XFlFB/ib2UeSCTQTqISEeFDe46jcwkWpvy4YMfycuwE77Tqt8zMHOJT
5TTjpGX17oAgjlfUyMJcR+A3JPFBJ0u9wA/VHJt9WoFXMcTQN7EwoXuOnhMchcq5bykkd8uqIzGH
PxEfzZYFIg/ujIFy7cesi4AWpsa9Vl3LhF5YQqTO1wL/5S3e/njyrAnlVFKe/8shJP6w+WOo5TVa
kEtUuQi5XOdXRozn4fItAAY43mPgYmdL84gb3xhKB2X6toovWNO6URdRA0VFl0AV+i+AusEa2/CD
D4atACse9LWP1h3tftiAsZTmrX7VkYdTrmpDoYtAx4ZGh/IAGVXE4efztKvqHpYYTcdXRGGW71k5
HZnzAWarYTRyCNYT87PmbZZQFTQpWwQohQhpHmvhvGjLL4BglcY8D+8+VoY9GWwrRYcLcrHC9CCj
SkjA8u8xG+Ef+FHftmwlb7YiCt3IXhiLrPaBq4dt9TKnWNlySg+PumstxcM+eG3hx8ausyIVIpwS
KbS/yCWWTjh7E8xcUT5YrvsrNu8uqNdx81kCbIjCqoqhk52alC+Vq05r1BIPIgtj0FCWpOTrtc0e
DnoSa42ObIJTtqVEfmyJf1ioLFDUs+6LTk43Bz8DkG70B1NxyuaUIdf/uKth7d5P9PsHnXx5Zpjn
6AW6V6JtgLYlU0rJGE34o2wlgSQwaPV8ddDopmZv/bNhtGGnSCN271XJ1O+QCfcHDZufnEKmRNXA
mru5dZ1XLQsKTwDp1uhwfeeaqQLMyWWEdAXt6Mp4Y7BP00FAvy9mguA9ED0CRQCyC2pzoV3zOyWr
sPbXyhmxCHx266b9TgmYSqi/l143OD0R2s8W9JcFY6CBSvCLN96GuuswkK87rhGekvSqn35BjQFF
C8kuJ9eY6/IdbgxEU+dg3Rve0YZJIJKIhonqUDM0GaTnmyo3VCU5G+8ZiYFO4N+Vwo6MMQDR4n+E
b20kVwsfD/IVp53EOGxgxkUukoxd8IWWyBXPjK2p+E/harIHEzC6mp6ZKvn981d9AY9jYCI/dQJc
X8ra8kAhFadBcjjRTidj5FZeT818MZr1V8Pu2xWY+VsGH9zxGVqaz3mrRJ3tCKnCj8S6XbnAaVs+
5jgIospXpDaXW7aqSTeQu7/ycArx3EqoJxcqvm1lp3RG/1efm589oiSf06Htt61Xp7rTZlvuGYWH
13crjs7rAMSUBCp8fARumCjANQqVypSYGu91DVLSLWnGpIecp2TaoWYHEk2kiwD5fizFuuXPhlIi
viqVDtv5Ohuv+AgZY9YINA+aV3Ag88FaDd0Xgc5EFCYKab6OeP9dEvmDl4g0IcS1VozQCms0lMGg
r/4v20XkXZhPc3M0aWvFzRWKFfHfqumOZYMEVO+X0tV7HJ0rSYT4HLjcqeMDWxXw/KeKoVpxSKKH
Wg27f7kOqSY8uLHjYt9AwGu9clmIG0pDfsene/TzZb2SxU0iV8WFt2Spnxi2BTUBrRQQ2FT0yudl
jFdW2cqSxj2cClh1skf28GhxGGHkqaTf+hhigVGjco4Z1PhucXzvXAeaR5Ff2eEo1ccbR1deX2u5
/TpykiZmxXi/ekkDEDb5K2D/MmDwMAvNhGNyQo/xAdJtNrZLgmqsouMEm0uEJTvITV/b2kY1CJSK
US7IMEvSekHxhM3xeKrNgvEtEuzMfoD+8wmQYCGERkkxU4rruj52/imBipwX2S2+OCLb1JMz3ZDp
P8NPNpohpsWZbqQaQXsJ9C6yJ3yHQ8XB8Cs74AbpzjVjkIjqpGNZhRVkNiYNz3nIEcG+MQntox78
Z0t9sWbt5HK6rh2vHFygRYz6lferuBpN/M7taUN60yrqE2nfik8UsVB4n7jiaHwTXmSrtOXe05lo
27/2IcV72SKe+zMdSdB0Dk0qm4euSQ0fmWGfFZrftmGKuDBAxnX+BXyqqv2w2vhhlnEo2w+2r5ez
QPGrWbS8+vdjrvFqWhUKshVRWTkkRhd+XY9Ohg6JHAIkos5zg23/cKoCX8bVQmkq/0qWoVt7Xru5
P3O5ddAS9/9svOqdQZ8HJstgHLi7H0cfmj7eaQyTj1jiFEUxtt/GLbt4hiDYUzuf5xCHNKFLa235
TIBT3dw0ywdNGUaHBb3d1gq6P/tmcYTg8H6gZWSn0loDquyNTbhFuTtRPoIcxKJRLsA9aYEhQXEh
SBh8ZQdfyDO6UMVIHBpXtBGI0zVAIzh4JHHrVXvxakB2B+vnsbJBuImIad+amlOS6b2M1uEq88iu
jUZ1c7l4iXa01TvAd0ilOvArjEkOWbmzpgnUxvoYa0gY8VbuOmGiPO8Ji5XDuOVOEM3nr3tSrLKh
D9pFagHohkrGBwq6aT9ySqlyN7eTYN9X0PB1MTTcJDt3x0JGd94TifeRkFaIT80wNBtc61Q4VwFb
fj7NfgIcrIx3jlgLRvrrBMU1q9Utr28a1MsKGYTC0jUlxjF4VS/JwBX8pT9W3ev+kBhzAOuW/Tmx
xMaI66Ek4P9kHBoAUgwFnikMs7IyqEGqdjLdW2OMw1/XkDgb9F/OajhH2kyCNFmjqZaRMtxaKrG6
P3Jm4t1oRd43rRdh0LOp3pMxmyv8hgHLu7N7R0Q/cYplgt+1lZpR9Z+2ZhU7DAOPqoib5ITSCYcJ
KKZei9OzL7VOdGJBNg/RHB8CU5BtbBHD05Y/aXxNigiGkMc4IWRnZ5r8U6oFseFXzg1hHrnwUnSr
xQ3luIAH2RyBkhh4VcV7BA9QTZhyvs5ubMLQBtMo1n2ouRLkGEgLu+eOIx6R0tm5NAqgWcymA8bv
6y5nrD2yebBoaLCcwKqOjYxgncf26lcWDS/M5aScZzl8r8DsmZLCKfMZA3krtDfjpAKJGVO1pGGK
5v4e9HnCgwzF2CG76DpSWUPqNZmAGnvBE199PydkAS9D4rcyuOiKbu38WSiwBX8rzdWAS+OzR4tH
D9+uzlKjxeZqw9gipo5LxksS4ZA6PG52Q6Cu8M3LSKd63ryeQw8JoUvzI2yjF2LwyBB9qJiLnnf1
zVALc5kjmOsE4rhzdhRspJ9FVr2/M1DVtG/krabeMEEOrG2hH8veTKWiU88QLFvzEmZgXJjSh1WZ
/i04ivFrl/XsbDWGV5CG0OzPbU52RIEBhHbL1HW1l2Hce3FLBU24C0XtOQxmVeS33Tyvc50kn6wW
JdETY6Xliv4LcLbRBhvwJpMgRelMr1ljzkVL6LJj/3nN4Tcyxk92rqGYlJxh5iwmCdE4Hel+h6+S
uXvdwzS+1zvGh+XCtCVQAQRR8b1fiNbsiGGFHQYjLeWiuKjoV+rwbIbsvG/3DirOBX4TsoZL5xI6
j6FEqDumMqZJNgWHKn3FBZFS2bl0O77wC7y0zpw/GMyx3W9myw3eqOfazpULlouSJQilJQuDFpPl
zPfUmouEtdDaycIQCmenowe5KWT/ithqKbD61YJ7W4s6Ml4Kefu8duH+z63sSBtkvmbIekvutzlB
9usMwL9scPMahc8wILc74oI6JJJqghYS6ff4vV0G49Gtu2f4iwfRQZOKPvVN/V9xPbE9B6fAAOAL
hC6Q/C0ogqcGOaktNgZNWeJJ9wGhbTbAyDvt1gYuRGBxniba12YChTYAioN2asNI77y/naJLzVxM
w3eX3l+zzeRVkVsyXuc3HunWgb8jTGdTiSYsiAzLR84lVBALyXN3V3P6MlrgYsf0MSgrzf5dXutR
8AkxIempv3nbR3GB2vZzvSHOtZqHdJByhgrsVeITi2jucT377ajqCQr6w6oKqe7c3EG3P0KBvOyc
8a+ISHfxsK/nfyRfmaO/pF8dn5HZ3R5QR3U7g2QEQKWGzFtD9L3cAlKqV6ogEzv7ufWmGDwQnIwW
aur3VEORk2qiWQBmpuv0TQNpHdFHgu26lt0hJAlXVy/3VXndtr6UdO+zN5Rau36KLxQpOTQ1ABIk
X96GpfxB6BSc+a+SOPdEgDi8ek3cIYedED1u8baj1XNMSjNjivDCoxi7LkRx//sLAIVD3qgZgVF2
bozF6FvLPsBA8pT3z1LwMMtJTV5FTcgeDr7HMFUSu5ry1NkBRQM4t8Q+57SyoNdUncGRSEpsisGU
2ZXRHXli97OlD6ejYQgVufzKikQb7W1Je5UWXltWPn+2MmJkS5oHjc5EtR9FU6Qg9byRIlj6yVUx
LujPBckxN84p46aMsR3PWNkWJfer3XDFIDNIgurbbECcZ1SxLnEdZvR4x1tT7ytCtBXDE8jCNnQi
xtX6630mD29GAiwIGNGJquXTywX+b3IajscxXiJuyHOaA17+zKllDI0/eR3/zeON1MANDNsDq8vW
G/B5R3SV9WDa/MQ5A4IZv7IeP3E+9a2i34H+BnElcsLt5emQHo1k9tVW5TPjmG5/1VmNdPRfa7Ue
UxL7ftqhkEtD0iEyzLb4zVtLJH76mKTksa7ctvjjTOj/qIJT3w9XPNwHm9t776xAfADeWPM9Lxst
KZwDKGESqloVRMeK9NvbPt6NC/DRtufoVcJ8oxcRCStyvoqissORa/onHul5xc985szWoZy/stsa
FAfvBJ4agQd1OPzJ99GusMuz+BudJYxScQ4V4xK8RJljnq5yMvq1+Hb9l31PY+hvBe6PtpSqeLm0
hJKSoQbql/A7EYOsasX/xCuB7UL9t2Shhmfu3JgU+IVuqFo12LA4U3UP/8B8GWP0CVDzG+yMK6eM
ekUnq8n46Y7O0v1/njDPxrvp3yhMBkFhdTpaGcof2KyQWENtanwm6MMUTAdPLmUbp7G8Bhm3LeDS
oJNJbszM2SyyIQtEHJMJUSguaouKJlcvCVHfmvKIz49bequ91Chx6F1cWqu5RL3fDlZANaos8Y2k
YZJRfAU+DZ5UMJIH6KGpHFxNtH8sxSuHV6OT9ROmA5o0gxwUbIzcwTX4P4aMc0SZj2OMEtAh7Ip6
2zh7+tMdG/+G9DCvYMcYVMNj+MBB/HAiAJliam8Yb0LQCGkLuRTJ2cWMmdsT4a9NIhTeL6aaLZh0
gP6Ln3LK2MTNQvVrEc8HB8iJI+MI/m4GpUpmMy4kG2lH15MS8JvhPCZ6xTFz1/nNlwGP6Q9ykfvI
qAk7gQZ1x+u+lxAJIIUkjnBv6nsWqlF0vu837Y/knKw2Uy6zyVNssJlOMPUiMGoaOzyxUv0vDQII
mG+i/X+zRTkMtFnEcmM69MMZ98ptldpKjJ4QSquwpgLba51QHDOBg8RoLzjP2JYbqNydEu39zHuz
Dha9Y3Oz3913ynLsgsdvzWvOjQn7SFGmSJQRtmHuGUHYEIwEFGNCOG3nUJaA3irxpFkpo5hPHiRP
N1pvslv65GXs16/yEWbb5zyM/L+nRZTxpO7ggt/RK2E0IJ0hEIfjKWu4xOSvdCj1Pfogb8uT/7Qi
x3HF6b4ElZzQ5IKjmF13PjELZCjuanmI29uo4YZIxM8nMMhhS/gM3hDryqEYk2ARMJ9StbFO74+e
HlGyzlqA/DjueLWqgWvRnD68Aw+6Ua3lEXz7LjahPuMhb0Drh04YtMCAxAkf+euoVtNKAC8qiIek
b5fai/XYMzjXMbxGGQsdnHxh2mzeSkbfrZ+tvGcAs5DVe/1UlUN0p9TO3/CHlEk16H5cITmVhrVi
FaiaIQUYaGq/SIzrj4BZv0uWPj7xIgVsLg2fOIN/onAq71KhKqZp4gJsqXAek3XwYgTsMKkAVdA8
9jALezW7fxcTMFiwZJuI5DDhYGmGjftF23Q/iVU7f7geOGRm+I32RNicy7QdXhkrX59cP89oP2qH
fmCMxkE4Xph0Njv8bNCKb6ychDsGgqmxApNttfidkYk3Db3vrmCGsZJsPZ6NPuutQm7C7Q6HZm/5
M3zKUv0xWcdT2n9ya4LobXQRPzRIomJipUh2zv2s3Il/pq5Slne0eA5oHCmM9txVbYrPsC5qgr0F
/cwCTppZ4g2rc3Sv1yg8vbfH1IJdG7nf93UfKVNUHdJ3bTS1p77boWK/5XY+q/k7ax/45mqdM+Fc
9xBD2phVDp15hi/VosEusH/p82Q753FGtOgut7BpapQt3cKFApEnwcQy61rrj6XnzkSZfIZ4Ob5r
zyAP+KC74AuDm/U+CE4zWc+5v3Bw7LKYrbdxmz+GGyT3JtkScShgHqO5P0ciOn4/Rdeq+CFShn5e
hi8fxCYeImFcjcjkyl1OHqdZRJwUKAqkdx6At/Upo3ThnDNUI+5YRvG27lE3DNm3dH9MQcSvZOAc
Pn58SA8zfYvDe/p4B+NENHWVJbZqrW9nLT1m6qrGOqFRx7Bg2u7igL7YQ7v9QfNu7rPMXipQ756J
qJNb43DOt0DjInGt0Y9bOfrz0mTpjjDN0ULzSP3Ir82cOD4QiRAiJS/xVstDUmKvtHfOEsBEPXSq
8Zw1jPCx/MwTahxJw7kzt1cjLAHu9hbRyQ/U34JDm0PPNX2eg6Ifr3Vbn+WgDFyjWks7zpXwxCzR
+I4ukH0DzvjVR2gZ62YBF2qCyfE9kBpEyhUGo5I05uk3gv21DFdL0eC5Cr2t2PQsqEXIcTXA+CHT
sF3fbVVRM5t5qO/AfT8TyL3IpP2YdHkJpOHrzs3iCVXUzYGKrbMwAq1CP1e6Gbsq4RMNWCvBsNDl
dcmdzZLzRAEhlvq37dRcX6U3OuMMOiuCA7Ql4Qqe0yYQ9iXrBq/e27a3Z3gsp+Uu8cRe/WBsBwul
dcRybhft6t2zYn6BU4NEBbS6T9604zPnJC6Lg9Pxma7axjoHrhiQLGyWEpCpPYyEvUFAobQ3dmZ2
uIT0PBvIMOshSPvrRbKfB6NuVmSD0IMmiyXEWGyjP2gp9Ne78FGQiTCF0I04p5kuhtFDj+sM90EH
E0RykxJW8RbOqX56OHLwUQ/aYO/calY9NfBm7W5KrDUCN7uuzEM8tmCiAi8ULXEbXcb6mJ0Ry5Sr
vNoCXUWg92yaGpcCj0V/nKTHACieTw7tuzKt7XAwpxyVdVw2FMQ2IE1bZyJ0fjU3e+xdDQL4KzDY
8JHOSkAzLKdXN5pMh+OMg+z/xFrB1B3DG9QFCs43p2gz9Q+nmZl4gvYSC5eAnA8l56xi5lRWiiQk
Wg13lzTDs0fdVxNPzhqg3WEmhLLk+fsjt/S2x7aflL2KCKbkceMN89xN53QNJakBU5aGNRvbW1Vo
bd+csDtd6AgVmtO3PXm41x6KTuLKy6EDy+kqkNEyBjypCr7iAi+/1Qo9Rx8DJaKPdqOaMgCLK1jz
PPqXbO7Q24Tmt/axWn1Iojf/EfPqdNCqnYq2nx43LSSQfi6DPM+gQHgPs4TP2Ws5mp+P8zFsIYWj
I4NZmX0kPgEbLYQKjfe0lgwoiyUoDM7+RHfbuTzvaiQuQI+cBrRHCTUpU1uP5tuMootU7Eul3YVt
HqONDMxhdR8NiSZzY0zfO8XCbdSmKayXdcK3CBIgWol3vIFzSzmmseljXO2UjrWjXpUaAKlJj9/r
ajRTHPOjtqTmgqjaI6j1Sw9f/m26yoLt0NbFXCpmMbCsz/NTsW2bIS0aN+elRwtRBYQhIrsi5UJY
ribs2tAyuKJcBUJ9nNuOBoS3HDyewvDr95dYHKvOp69gnbQP4dguQverG3g6TTFF2JtUK8JZ+gb5
zo2mCrUsLWxP20WaGO2mym33V6kysIl4+NSYgw/YgyJsQTjA4GTNKJOU4LTWdlSvxOlEEc3YwXxh
sI+C5/LNOOzTNNsym/t4FvqdY0XxpcO4tvQZxtcpJ/2yZctyFL388UmtEsOcX2N3cJzeE4vitg/G
QiZ00rLlBXjeg6H1B2zPg3pEfce2BNr0YAOglyUf/67MUCB5qvdjjAr/p4NQ+fUl6fSPGpe0ebU5
7ga+uyujp+hZLOjS3E42OnSVCD6Krik97AJxJ8V6iYp+5fhlzEjz+gq1EKxJbONr55w/TUpECr0j
GoujULmRbHSeqPO4uxGfk8lDHQLRCflFIxdLJTlz34cqyycmPaMm41PGWmFatYLmI3tFbbm02Ks0
sGJvppg1vUlt3EK0CqRL/izbVb664CsznZbq67aZad1/fZpmwGhpFK0fzBwjczyILfrx0aRUfVgM
nW667i70LjeI0zZkFgXncwyWyPRLFgk74oXydtiCjh1AHbcojIpMlZwT3+iq6WuFYvM1t3yZRf8u
il9Lsy9deQthQ3XH8TlJCLiHBHvnNi1q08Osdzt3lwvz1iKSumLA5RJWwHf1KRtqu5DQLrythQzB
pYr/HrQChEmuYY4srIdyvwC6IU2fTOpjHjLqMlamU0qzG4mrUMC5r96sKOxKiNA3CoUNhq282r9R
P+BTAm3uovDeWeUioetJVLUWr4KxSU9SxFhItmFKhwTqVYv0XntllrbubB5YMTiNyV3BymVSqY8P
BJghuy8uHh7r8yAa5UbZW740PFViVOg3HnIx5a8/wAVLgznRVOx5WFWjCKL7ep3731Kb3+ppE0Yy
2l5DFQ1g5tavadg1PDQ1+erMG8GoMSbQ58BoxgvnRpdWNzAxcbNfS0oqPJhkQP7+AFoi+xyOwyHz
BwWVyjUEC8y8QfSk+QXLc0xZ+uZIFwzVyJEPco5h+MquRBDjmvEcrngeeuTcZmbgIF7ZrSZQcaVV
ND76cfzqUQMZZxXUAn5Ydu/Oxfrmwm9ho/axpCWqr34uY6i4FlOwG6mVTNz3EpYZx9S1rVZvDA+t
o7OR5O8wc5gHTZiS33uIzgXZiy8r829/kttmTWIKYXQ7vl5GiEEQqmcvpGHktpUSrDxtT7gNyme2
UZGnlE0B+g83W4pRBW39DPzBcXSJwK59jLtxAOk+m4RTfZVyBa/FzGAjPub369p39Gh+6+85Gohs
G0K5nU9y0sSrLdGozgl6Xbmg+zzQEBz/C//nG3GKB1A2TkR3xg3NbSXPl/9GNFEVXJbQBOSsAqZz
jOJ1EAGkXkX9DZmWcG8n7JL8KQ7zk5XpW05lndkLVDSWamP5nkhBsd9jnL8dvUOXI/LI+kzpUTLJ
JeGJpVGCdTb9oV1XOr2ce8/5vExRV6fKRfg6flUBEHIJVUF9EcY+I5VIOQAnHi3vpP5ID/k4TPVQ
BO6MfTymBOieFHs/JZJEad+UmdWo6hrARd6gevwN7Fms0XGlEsOswpdPpnOZS0ZhShhI1fLsFm2Y
yIjTFjemHMP7fVdKTH8f1V4JuvIcOVMu/+cGFyb+RCTl3jbNICOqiQXmrBJrQ+oapr7GDhPsjI2k
m2m1mxiEw7tRqGKX0VFlXIALiPnk5U0z3KSlraPHrOY6YeJFOOrR//jP02KMXpV5DncbFuGO7lE9
Opw983UfvbH2aHHVIG6vF9szkhWYAfRxCSDCHZIaUNnEDdPcAQPVoNMYNRL4DWR3bxlQoOk96Nhs
79AR9l8QdtiXoLDqUSu94AHLUo2Edqj6zBgmppmfRUDVuX6cXt/dtIsgCjaF8yX4wff7XU6Ys8+5
C43Jj5JPZ47tGDBHkr1D4GJuf4OJ1/YqZG2eS9sChKJo3Extw+DtScND/6QZVNowM2JWG2GaoXGj
IWKQWKI24Qw6mTEzcNXmBUxGJQkCxeyXLlMma9mnSNu07PyKO3tCT6AlJc6mz/HWue7ggNVnJUa7
cuXCLQNI4h3GwULs9RrXg1b3yFQV8VbcZ8SheDTDx+9kFjzdeQE0x7S5Tq42WkOIZtA0KQvT/m45
niGB/1DooQsmRncIxQC1HxsoMlqf57Z3RXf2WvSMuqbVQnS+1BPMtodOy2S/jiGXfnOYBDNlPKCD
hH9zbX1d+Ai0iSfVHgZsg9RkAfwgi9flH3A07fiDqKCQGpzW4cWd/2JQXJfT5CNHQAjGH33dhXgi
rmIJ2EI8T6v5P8t+g4FMBehxFl83YpI5q5DoPfq6HKGS1GcA7s2y3CMj71yeKXL9RAaBTIIc/LxV
2VwDZgFTuDHt8Sqa2eSsa3eOw3hPm2aCmxlKYFt/xrr/kOk6U0grp3rxhfXVE2rbi1pHT8MOevi0
AG85CQtFPNotq+jTCf1Khq+3EUYLFlO6ZOvACzck+eflyhTf2ZegJShagXOBoeZWhL4IDdvB2qLE
X3UUrwhduwHFGz0K/rzue0AHdBETvMAPeGI6rh13JAcUZ6aHe425uJPd7FZSyWgj88CbwkUKPyyy
sZQi/XxSLaP1JemLJQ0ZQP046+neXuVPp9rD3+5OnGcQ9fey9jMCVsNef5WvcifzjNUxQB/JE5kM
9mUNkJq9WCVkoNEqrqYWiQirUmBwnnA9gQL3L76+LJymtshS6edVw3uuCrtMwsF3D89UH+1YmGZD
YbN3HhX47RkPs6rxGGeCeD+5pUFNnmfyVwYRm37qcp4PjsboRbEDFeV+hqkQpUcuYfQ4ybNtoVyN
bvxEhpXXFrtKeaftr06D4c7R4YQ9dn68GlOhBymOot9eQSZLJuGm9AiE0ZFlmLEgwOhnlONd6L0y
FvwLsBQ1vn+Za7bqbkYDYmcEujtZNVaYIQIA2xStCmz4tsPn5Cx2+DUXZyGQUOax+pwFail3yxte
nWXcIOQGfv+yaSjpa9i1LM5ozAmwQjflUpDJFuD/R6LxLkqH/UKSqvI9BJxsZ/OONSJ+58As94Tl
2zck9MIaZXR/zO07SDPUWVhR6smILXn94gPfxypAK5tvTDyiwHscWgGcTtP8d5OarcWpdxrjS09f
mT+i3C5l/+VHKqp7wRY7OZgLLiZDo4Vcbbv474m608t/AnXlbVqVhnwPpyusbmQ330Cvjkl53qh+
W6pIdMnAxnSZ8jBcrcpybwbAk08aViV/jFVB0YxDS+T7KINriYCT/P9iRV5mLDEdB/9Hw0/6eOJ1
J5pNjL9MDQIeFdF/QrN+OrQeSyDKBGOMwI6mZBMlGEzFE5Z0zUhLwN3qpUKtMa+YAro5z7dPMOSB
Co90drFBroty1cr+t3GjTP7bTjkbCq5vREWt6QWA6ruKmeIcjFltbOBVqZyVKfvJPcvNPYJb/uHf
I3xNe2vr4ze/68DoPj3lD2T5xhpXjyvkAG0mkcbdNQroS6gbiVi5eIhy2hTkGRMSQ1IOt4dCn1We
nlFo9qgNvEX19nqLMJ+gE3udybYCX0xG7TebMFpAtPrBfLH0ohpheSmn53TVkwT5Fmgyas+5kDs4
S7b668eIPSNmHquS7IF0AFhBXPZVdjL6GqeDpH5BFnLzfK0EoAoOi4tnIldWz3ddHTj46zA2u6fB
ZPgNVUofplgL8Om+f9Zb7pvsAgqztr9ytsiKQTYOpIFw5pAY4P5aixMbZ52wAidczO9GVBWuyMpO
nh6JLrwbKuPjSGvO1f0rSYglmH6wTObbtVc2pvaQItKeEKWZ6M9POPq6hCHobdQ/jHQg63nKJWin
c/i6gvYouRB2r6uISjVWaEtxnX/ZlTeU2AxrlQtpC5YntfgbYXCfokaC8R9Yq8elp00nl9vaZHUJ
assIok/KTRV6FMr9OOaMjL8Jv9/9D8+MVd/6xtsTMWjYgIdL8raY7L5cOumgq6FqAr+ih9KtuXxa
fITe4M5JfgMarxEnAL6goa8Uux4IO2Xq4HWt+xjnTz/VoQhMK9571zEeKuUlEWITKSAkaY9WUcU9
ot/jj4p1102pCrBSa6wR00ugNcoPStYpBr5jqmATp3yWFPy8vI/e59xdQ9auqql2R3yBkVAHUo+l
S4NjAgAA6DRgr0/BAYE2asDwIvmFO9gQovvwfNwL3pvrT8vYSU2KGmiu1QH2+GVNsMH1yA0CzHua
TslvGEd5Ep+54p+0ux3IWXP/5O4xlXHeXNQtx3PVpVWiAnK3PnmDMwAa6yvCExA7E5PSTO3j9Zfo
jpTFofmzlLbE8PDpGZ/bE2uOLYHTZuPDgVeEOtjxIdkFnEqaUwFe+PM8duTHrQT7kIba69POnThe
bAutcIdTPpk9GWlVqCQ4yIu4xoTWficXwDZLrPVOtc7kusic35GXDts0eD9N6dsP/VfCFoVQBZ6o
eNDTcXBtCP8Of/SRilCc2S36HeHhw4MYsIHtx21X0CetVB7M6IgHJrhsGS0qw+WI12wUJGBD+3Ru
BPbH/K9d3lapGs4qXZbmfybt+qj4BeSs4vqcQlfOLOWNQQmWXH6KVSStRrWRsG8NvihE2CCjIqVJ
6caP2Ilv+zyiKMgPoAvYNovO1oGYAdeI+pRlgf0rwQSQDtgCpAYrXTG1xFIMCFKcM4tW5PTn+zSM
LcfqfawuTBXzgr0hUxsNwXfgp7R+dLT4rw5Q80N3K9mdIgGUiatnPxeL3dMyCGfLFkRlCZEx8u67
ictcUJ31eErUhtP/wxH7Tp+BvnolM4e2DPbJUeyepM5vEX3ubJc2oGecBOwEnbFfDGCI5nxhTDnr
F9gItLsWegMKq6Ut+nl4IvHhl6Oc88T5fbfs8XDQzUxOaWkClADeKw2ZyglCdtb9fNr1zEd+Wk7z
q5zL6qfcrRVSfY1CIvNW+m1GlALkgtigO4Ku2qdnImgWlCbDb0o37d11Lcd8OwIBJ90sPfuGXHwV
yNZdSa9baRU5lQaj8EdrVN9AjPzI9+AxuZnmVwFCDvr4XLKvIRN0SVW7Bpw8wHIaxZRdUYFXaXX1
r9Wm3gF00chsiRFj81s+4rp4C1gw4jhIbqFCcM9ZSm9RGwY/fUyw74S8CsoJ1mY1nckRWB6MD+mU
eOtPp3CRqhTKZE5M4HEixnqEDFmzXf5+v11PdrqTgV7Gk3NfTrp8DKkCP4PWmmQS/ptyRhdlc7zx
HnsUzqxx6DgwkpPgGuOsJ6NvReVtVOUbPe2IMZ4HaB3bkmKJE8oGcVGuPKAONUOJe9bKpmEC7bWi
VlKnQdu6WS8n6guEAWGdO6UxluJr2bP7m+t/93HGxBBPvwS7O35YE4JaJ63tYNeHdHeBeE6pNX+q
jfro4uhgtJI1M6ucduicuv14CZZg+oqxSOuGIy2ZygpBRei48mWFyPZ2GD6zoeMjLcEsqaNQYM7l
MLGrzl2fVejs7hIcAaaJl2k5jfQVAJb/rK43y7gri5xXlQd4mi9MXHM3pgXnbZ6Pmgqvb6agJWat
aQoJw7qsZqN2KSMwC9Yf0RP83FK0UGly55pVPZ92nwJr+uu0NMA3bWuJrFa/3sQxCV7YT0VHELGF
VySpZk6jfEOU6zU49fVi5O216fBVZdSuZD/J7hEPRweNqKAirfSG+DsYC6UPFEGS7v9PGEcdXkcl
D5Ps/edKBttDT6nbVymsRViNGKU75uMN1mvevAOOA77GqTFYPipj56zmPtAuf6Dpyt95ryyDDy6q
rWS1bDjK/OYgYV4ohMgolnR9fzwe/t20GF7wNiaBGtdiySXjajpR4xIuopw0pImUOeKfCJ7sy8bk
ytru7gOn/4dRZ4XEgZbpRnFBu3vbBkgLJOyekKsvWwb8zl6WFH0C+VMXVYTC5/NGeKN4jUYN5AX/
UX91BWY3SM1lWODzCoAvoIqxCS6DBm8oEpcYJ5nWd0C4ao7LqKTvjOSJpOjmiv8fptH9N+43+Zvt
F/IsNog4pZsE2s/St/WECOe3zdOg6TVJLe+JRRHiaTOa/pLWIg1PL/XhbRaP2vKljTy7zbrZo3Wq
ZggOTfQRbbB6Ba1YpAP1Ix3/KqALWp0xA1R1tIa6AQan841ZbmWo+rF/eaeLoWNzDxkPk2SxiAJD
4VARloAZ+O07jUtx7yHoltIEFS3yOtMuw8pd7o8mUKV32XVnH2O3fcrP8NdlOqbQAZhWQUmRWsGx
IX8y6TT4yvbH7Q0bDG7WszcGMzjjd5QrHswqTcSB2PwZL6r0vkIS90a2Wznkqutd1MuZnmPfD4C1
iZ7XfAhf3KXG1SBk7GWTp6yKTWYg5uBV+WQ9MfShg/muCoyC69Y8xg2TLLgxV3Ku8LxjKx1Xuqcv
4XUjS7cFenkPk1CDnDPzPNsyI97VqRW9s5caw6BRCoS9yzKLIcrWFqTgqn7qz3VK5puNC7VkBdaP
ugfVBqBzOduMy0IyMmn6nrw2GImXlDZKQTYALdXTnO/G/WgmlikwGuHvHL4qk8HOF+E80L2WmWcu
3rjdfPzZ7jQAwl9r3txNkba81pAAVWy3SGlyC44K8RLuPlAMHuUFcAHqz0fZwT9uhdSIn0LeFLfl
apF0gDbrvBnZYdf9yS2hHeQ6vJ+k1fD7Mql8uRvea0/7G87s7iLjLsq27i7UuIwdQCdTr8zFDoJr
HxEvS4np0uLUH0ZjPq7HGWw02gIKb6GSM0qX1KTAKGWvDNS7KHHiBYiN8cSS/FGs7WYyhhSz+FdR
LQtBRCLiFz4kNNRaqpRPFXS2gOKwlVN8EHl6eq1LU5dVIpveWF50Frrs+DjAMdQAc//3xSSvuncu
o9oDWIxAALsf9IURSpostzsy+Uoiz2lJZEt0x8F3+pXXkVdoTGttDUo2p6GBon5lbu9aBhvpQoya
QJYDHLYcVFanha7l7XCeMf5hsvVP6npcsdcz0ORvmEEkJWJkRANGIaG5ebpZiGZNRnErxiXctFiN
p8N+17lhNZl3JmXIp5G0PldM7Na5rJfLYFa4P4/kePlMBtEDSBiHSOzbDKXhujMN01UqkRR82huD
m3JC7iJbCA5f0hMS6cBabBPJ81PIjHUNEnX+uvYlBG8xr9rVvRVEngS/iKdLSWetHYHkk7w7sEUM
Yr4LXgeEgr8ATlBudUkOEleWjClCPXlmYpsVdrg0wFhCZMz5j2RO4qa8Hjf+n5CQ7WBukmrX149v
sJtM5GZKrMpQIEEZTzGzQmWdwGv6+ft+pvs9JWLEkrdNLysk2q88YPOQrB6hKoYD7O8YsuIdtQog
fGAvHSpbB6GAzLyUCpimi8TcxfMCWO0oN6PFYWM+9qB6f+E+t92t8HOQoiZALHi6ODkkmrDIdpLX
3xwPfHrnpfrgTkeuBvZ/ZixvIhtEJf8CasQw3UPvosUIUhGnp5awAKYWuLEV8rQ47XEKZrdHyvgy
8tMbOmJ4hx5/nRQq1mSySkcSWqG/3+j5HTvObi+vP4Irhz73eIYRdRt9nPszyZKRJ4/89UtTgrP7
O7iDMcIeuzGbd2mpbSZ0gy3VLQcoBD42s7tGH6v11FIVBr3m0u3agzoWkhqRqNxHAqKGqs3uQ5N3
NwRQ3/WF1eaxA4BtLn/EjeQ+tXSRMW2n2M8p08bjnwsWBH7OoJaNvLZdXQ3B0bvW4fV6z77fYL0o
m9pKbGKvZiwDP/svfx5Etmy3sSz+1hwu3axQN/PjvuJR7LO6K0x+y41R4ZRUrLCdT68PGISDTp/1
LrFI89e2G5yPIY3JZR/WHzlEjH6FuVr2V2NNy5hZplUT8H4OuKoaoNoUvyPkxeQ7KcK3kRRXuLwD
OD5M5MvopR7M7KmfSQDDE8tdJS9kkzYQnuZUrM8zfZ16ZGU8AB0IHRPwQYLXuWxE4eUYWyc7sFGe
vGW8J4T2pLNsPyB/1zO4w3mCaZrLqDS/mGOH57JMQ3So6CUz+bSnuU/4yS4rFx8izqgZbSiB+hYW
79AqFt3PHxeouWHjCN1+rNKEb8KyT/u9/H8g+ufrbrNTd+Dfiui5H2iehHRtqiGUANF53MAE56Uj
SvpMIJBhw9dfG/ea71j6wUGI1gd+QRUTETpJHWp/hlouDWPlHjkTSVhUiKExrc21dvalKvt4cic4
xqKffQS35uHpeVjfUyx+Mh/ccy+RnJPmE8tfl61JMDOhJwMC0pl8HoYygtmLW+vD9j6aMRnxkcCR
kwDYRPTJV2/Bg4UZ/UUDqFPYI+PCJnkR4ZFA0oa8/Me+FHGFj2ICANnpvj9/rAdhr+anlABPQqSS
iqlEmmnOvlmvmzzJhr2nx+pzwrzfnRu1WLymbqmu4QVSzZC2XnjvmUUdD58+PZiIt+LD32TmB3Ng
+yAYqdBCwvfBccOagSixorWyvE7rEjjqkPAFdOzXWTpevlNbOxCT5w0jEO2xj32rty45i7xA+tND
5tAGTcHdO1l00gn1B2k1QMP56RowWA5w218PUckDqf/qIerM3i2QGRby4VG9dlkmLGoqivu1wXro
aURNMUTBvzt5FZwoqjgof5VjbPyNcm34WmK1HY4cpl+ol+NMvBPGizMtcp+0wcAxKgnAcrDLkTAJ
3vbHSgMKydHE6ooADUdfshquG/u8O57v2Kkd+dUPxNS7DYgKDi0GfLoE2x1UeyPDZk/d7ZnS81F6
K9sRSc2/knwNk6w6yZoaW961Wl1SZIsLJfQyUgzsM9k/8Qu9+YVUuewTgOfu97M6ww+qNe7E/ams
FQbUur/J7FCBaCVn0WF6htjOF3dpO6vyB1C6JADijCUB+JMrn7bI8jI8kH4tBJ8YY4kdljNNt2FF
1LlhcpkdK07CJ6zI9NWUiFqLGiSvXliIgUd7j3D5YfukIMgY1nMLiCNrpxQqR/aPLmyrAATeTAbw
v2lr2ellCiUyUHOJ7GHTYYlR+6WwfmLFosNpsH4I3CG0eSZ1IWPg6eOW+X2m9OdOMt5F36RLt3+5
bCkaj/aan4PUz1AI7T5i3IetPUwCufC0iiOXDtm9WP85gjZrMxX1PqBkAtF4V1fCGTTmDWFzRhB8
YZB2jl0aq9ZPX4yBtJW5TLOoGQiacMSot8nN6RkRRNyLYebGqqaiS53kZAm2N9foNFjtzKZo97Hm
02wfEGDt/ZqbrPW2fv8slis4PzNXu0762cgvz0UMCx5/zaixnvxjJgDonAEWOdge6qPdQ4nt9MEh
uIGSNfNf2y5LZA3izh5qrHUrh1iUngKMcT95BUyWtQgSQWtvEjBIsx9cllIHELLZfNHEp9nXnNu1
3R770xIfNW6Ws/ZjkyQq121rnwkh/oNM7OPVDzpq+pNy0WMWhd+ndk6nHj0LGFgKNHkR7Ilgt5NW
u9ekm9IA5vabHa+37Zr50unDfxLSOrfMvLl/tevwMHMdyoH60mrLGKRSqKJIecLZlt5qHR4FuO6k
VK+ZLx+WDVxyd1c77yKpVOnpyShub7cT4lhfCy2J/Ogp13iUZXeskePJAIxDYlVbIQ7qW2hAEAt/
a0nFK4kpi0PlT4q28qIS8ZF3leuz3Dsg26y9tNUvOqppGKTSBe6ot7eSW1YAst/IdjrKUiIi9shQ
JIoiMIIdMCFbxaWwog1PQ0eMEvXysRbGSgefXYs3RCTwt5AHc0FVBnlFHTG+/kjsEQp2biImimO2
+qtmVO9yXsrFkTmlMtxsUKKZUASpb1oM+rDGYgi+JgGbstOt1+q+XVE0IUrNuL5pi2E3SUN1rqrz
cLlzHjCoy60GHGWL/8FBsj4pEEaKkNPUchy6x8k5kXoyvxgnxLszEzXXn/wBKFRGYJ+LZxjZGkfJ
GXC3gir5cmyT+PkCy1u66jhOxGT1I/EyoyNd56aexS3vV5eKJcNEequ/c7aTt7Fvs3nULyF5UkCZ
uyYWaFov02Bx3wtj0rDmjhQQ/manwRS0Hoegx3f1K+rMopuEmkZnn8zMLE1E29pF1YM+uimAWHz2
Fv049/fmuSM/z2tUsHBlRRTy/1cVw4rZ/YpzVHm3+iWkZ5UoB8QXve2nKWlLQ41U8z2XjcI2Vk6E
46cDvA3K2YPWA0LmR43GkUerwuw1aK//x314q/0j3kg/nVF3NF4xUzFjS+TvNHV0PmmmdYvSGUZe
XC/ykZB5FLEoXeKIyxjW41DVPp4w/mWHdAZ/bW5SRNnARGKTUkqmqXXziBa66xhd961D4Qs2o8Gh
Pn+dukm1pVSxt+zTp6EZWTCmbfdFA3LAZ0pkfhv074mUjcfs8bbjA3ERqEhwbeuNW4lGgk5ZB153
Cbb9iAL4H9Qs+3IG0gYXTnmQYSVLw8t++S5Rmb8VIkFx2jrWxm/WwPQ2YuNfTaBFFpWmh+grg7dx
2QdvO9xHC/ykOZvwkzy0m5DYlJWdb3yXrRqVpenYluH5rppJ50i3lmm/l1y73ItJr420fdlObNC1
pz1dcOxN+zxTMp6El4pfsaz2yofeN9nAmb5iL+hWg+F/GxUPgaqzpxT95bAQ2ioly4Hd8tXL8KWW
6mhArOVT4Mav1DRUFf2WPMZPLnKcLolCJrS0/y3DLiMJPsua0KEM6OaxEevadjnd55/ilwKzl2at
dY5YLxPfKshWwCOdAw7efko9CL096b2quZDOny/1d1dKyVVo2oKHYqYQmEWRW1hGEIw5X6UHgj5F
fjNhndz9dFrYlu7F76gixufQAIZ0qEb73jq0tM3bkcOviQLG4URlrEGaTRkBF4VL0taApNIM9h3B
d5MuqVigkHguNwd6ej6BvWj7buxtaYreFcwi8ypVeXKYcGs8S6t0cSKXPIoYMNzSqeE9DU6lZGUE
Y1uaEwbPa1tm62OGbnvO9cFh7QzOIQjv70a4kTmRmO3TRPyxYS4bKq2WbsJ9ZBxRwLnvF/YT10ay
iBRnm5JyHETGvMnROS2aJLbr+Ci4whfKlHG1cLP0N/H8KrNVMdXmSBAamtlEG1DCDipSuWpIfApC
Tu8YYsAwn/CxXDXyFmJk9laD8WOsKQE3QdJ/JJhwQcKQNOEqNlwibMheGA73PUNA4FOJRlH90Ddq
t8uqYyjcQigpTsVyXPwTb9lBQ0w48wcUo9u2dvVn5GgHfnK7HVtsTB4uvmp9sik8XHMA2GgEwm92
aITPvMZHEtRqgcvAZqVm2Az9ZKWSZfYdEd4SoY2rDYjlIKzhZYwVD54PCDrGt45W8a3gDg+xcaX+
c2qywtTrl8eJok7IAt5Qk1VIsgxhTL8uiZchzfxKWiAbU+PL3R6+FY5IIs5Bt6g3vtRIDx5eBkyr
nj6l48+irWWsrbXF9ebWvRCD3wN4SWNUvkmRGHvlyAFgUxywbmzIzhIyOyJec4F63gs09QXL3p5v
niymMG8wsM9486n0FKYSVR2HjmYqkqxT64asVTGBqpl9e2P2fhPqyUihxg7IBirCLo8LiJwpynLV
2gCnd+RGwfEJGkeGpWH8YLKr+kN1souD+Mad8I02hK52oYizQgenyy79kpR5KeotKzYnWovuzFEd
0R/Gn4Og5uYyU1ppvlljlRNaTCvULoYcCWCF9/LmCkGUjp61tOpYGC+5qgX7PVzmYfOvMmQUQgBi
Vg1Ho//9HM0iT9EQoONqcntg8Yth5UiThhZ152bF/6+UDrlCXGAtiMG6eP8tII3bLjtWWG6LnEC0
gftxD7YcnTh4xsXLM0U/vW5ifFOwnXpKgscAXubqGd8JyxNKN1ewnzXpC/GH6/IN/+JJB17Lp5V5
o1Vbao+/bjFIZVSjjYQSiWz2ScETi0F4mmcmQfQOytMfRKeT6kf+pnjqFzW7RQVBFIPOrKIlM5Et
58jFz7FYvMnNUc4yUfTLAHfIhdqxi8duwqvQgIj+gKOHd2t6gom9xPNSb0Sma3RsfA4gHnB/o6yy
u/f3e3+SnIDEQKr951J0smVmTWuP6StVV2zpWpGPAAn6Kcf4o3pAEawvGWerWME6THuJWE5/xZSU
gusLxVPIHqydwL9su/ai5xF8fkIkpTQBYOO66VB1nwpchIbR5kZLXtyOhPLtnZLykr2/zyJoVsLm
1D/I7u1fcQsGy/h3btx3QIzJ5fYh6X6It87ObfdT1d7mb5CelnYosUX1kF5+9ww8UBT0oZmm4RlI
5zPzWd9maxtLNwKUZXnDQv5LU+uJ9e70KQM93Cnu6XWZRLdgKkKl/Yn1hdkOVfn2+iuqQ0mQx/qy
L7V3M5zglb58EJlBqxa5GwPRkJ6bJDeL1KM+gDZEhG3E0y7hndbvCNhiP+GMqP7bbRa3Cv5yoyjF
0NCdAUWg9KJmc7Q+WF61odEUtS48l/qxN2uyErS6jFVwiyC1G6PLfoGN04Qhi0gKD8ElZvEjSAOH
Cben+Cz79UvxCo5gu7lrOqhnI1ySWKXvhWIw3H/ufheE08YQsZycMcsL5jhCOcBMUERSNzaNQDC9
xEIEtpEym6vJ0a0e6KrTjymwJzweTmwXj8WwgB8Fc4oN9O/k9IhJI2YW5jHCiVxjZ+Yga4lVzHaz
f7J3qUweuo5hr2buXIFqYFE5GLmPPNu18kzS6xqQUbHFJvSZfmYWynMRmExLtz1yY8AQamune4Jj
6WUTcFMT/8KUHZyrnBgG+Dmgm+aJO/8kzkQz//fRQ6tH4lESKGaWttIAOSoCVJUxfNx8eDrydH17
b1pDHLgty0Dxb6Yoy4QpluzlOwvR4OnVLUgJaciRCiIOgFZd7gYEM6HSsyhMzR4zInwjoAaXrm7B
riyZZ0KcMJ0gvZnIHR2AOiw6+Kj4Ea8SMV5jO+M89TDEG2Dku1flCeaLGLkwtVSoUJjrU1I2uMon
AZ1WFVZ4X51moS5M318zwqmL46PMUGNxHCEojbT+t9oBfcCqxrp5sQCCOgOd0glvh7Oc1MnwfQXu
VCup8n75Y96QSUyOHJ/rD18l0sjYQnCvTT3A4dkjk3YQ7b3FU4H5V9nDLi885NbssolIeUeMhGi9
+HI18fwMWbCjhtT/5y0DR0hR2VsF8wP10x8IiTA25/lKMyiECze4xvhhfWKmT6qDwm2bYhlHC3AG
p7cJ+eGcz8bw2PA8XopWHXfZO4/GQsU2eCEzckv1UxtUwwbkTs2ymbKoNi1gQKe35WHqu+WEDZP8
j3GLskGtwc7yXaw1TO7tv2Kmt2Kcx/Mf6LdfhgyLpIaaz/V6BvGYfGEs9SCyZLDdELTfduTzDA6V
RRcjFpRlJlWqPEKf2aIUSLcMyzq8ZLnhawvErRhaSLwJvmoKZue+EZqmKmfT3BzS18lpFLrAFnZi
/kq43IfCGJK08RFGb2EFBYWHQl9P2yW+DIWXk/2CMrGBsSK0LZyHgtYVx4Rz438NWR1yda/53u0n
3WmURagPjcCudEd3X+38fLAu5eQcVSCd+nIOw5WJHF6tNuGClRkQrZ1gG/6YIqa2mTCF6UqUiJMq
gBQlUaT8GTLgCFZzV1ckBQpSwL4QOB1VK/CimVGmVwOg8Wy+z+SO6OJZAGC6pCPkfUMV2TvKD5jK
rXiYfyadBsghfk2f7NcT7E1RvwNxpI8IjLQ9uxPlHnutQEC5QdIXPEdLfXvxfMOopjVM1EwOTFSv
3gKf+go8BD1G2xqz1rG7VcYMEEZUL6Iau7g487FzBMkSEbh4Tr6U9/PzviFVbu7j0ACqJjhI/zGa
TUIE5OMfSRHNiC05JLAx/3/Vw66PeISkUwv1aq9Q/yr6YP7QBVWr2p7fHPUkfrPrTDRuXCxo/CHl
SYENZOEUXHQQ9GuEplfCeqBqF3kvRUFeN4r00bzKiFaR9pWwo5NkVzAY0bf3gwa0Ad2nsaa7W5MN
2EpVRJOyV2sA/Hg6BgJ1YtUX+CKhq4tmwvTj9XtiVhR+SIySFmCGSdKSMT6xMttzUCLyb8xxrTro
5A2Snb1FaVRSPDcRS9BPf8c66rsMX4+nr4FUXNtkpOfAQP+TAHNvI+bXw6XFZtMUF1ueeivPMGlU
xFADVHDwwnubHpX/sxPG3ykJybgQVn74Alrx7wfLjdjJdSHcIYxGzV6SMeHBKwAWFfZdmglx1fnX
C7mT+VpDRo6HcsfBfC+ZqVFUe5UasqlLw+/CDoKzLqqw/PdGnhbir4w4UxKP+T+gUxBC42NRil7Q
6gVGOqMIvwoJPibSLrIHj55NBWVYg/Gt2Tm+D7hYE9odQfoZmeqrNzU+8ZUu/pB3U9ajqy2AmtZD
VOg44KNkHACLxt4R8uJLVMZqF7cUQoBQyD6JMGAJ+gR/sBWDaiwqFJwhqGI9DeHG6Mrbk6ekVFt1
w2zdfaFNiiG//fwfhQP6DgR3tqsZRDeZuhHqi35+4tvuuM+GuQ9E2MaVf+mDJ1mU3gEfWMuxzcm+
/5WGLvngKlx7xCKil0W/Qn+U78Gy++/OBZzfQ/m7RSvj0P0uB+aVdWwNd3ftaVVj9cy3c8e2tFRY
qTpv6HjVfb8ilfGtBaq/rtuY6+WUX2ziUHDz/KoeZ3deWEL35FcLle84/ihRyS+Gob1UKo+QPWe2
owi8Nrq6QQlQ5GDjWb1ml8Ah+AouPOmtNvYrw4zLCbvJcoUsOJlRp1szziQ4nQua4YhF6VmrBdNy
FOx//rd/ZasZaN8wygg4hSEzgP305CKwtO1V8m+a11x48TiM4BHJpiG5KgO5D/RoK5dInrkWblUv
jKepJtCbSobkN1Gn0YPJy2/9ame6Xxmyg+9ujC/JvbqiB8Kj8uhg0nbuSCY4nXbEQc8rNsqosDOq
XJdhyJyLZhMF+NEsD7pL7S6L9ox6PbbWDH7q9zpPev7vKXKu9KanFUjEewdJ2VV18Rlg9pqInjQJ
6qPak1HYLLRBMV6bgqQRqiNM+vy7ULujl/K3/dBzEDfGte12w6Z8K51J0HW/Drnj9wGEfk5Y8dn+
QTrTpAdYxRTtmuoh4vrr4KiH+C0qbK30TPLwQ8RQUoKQaCbE4pQei5kVdelgXpX50e54Uio6vRJL
PGOVLzJuddOAsDlJIvdoSZPp0Nc3NCc0qJ4x2f3MV75qf97EQYEjYv4xJQjOlT8VyQr2ZqGq56OG
DtZo/Eoc6ujNYcROB1B6LQnMBnns9XS+eUqY3+8IzmWuy9BtSJ+QcLUxBrvsBUZoZyTwwj1bUcYN
NN8mnKiBqyHgrlxZ+srEmdFh9rGe5FKj5UvTixRbkRvfqjsYrYx8RdhESOVMlFHJrRkQndzY7ewY
1ixiPkDx9dWVeApA6NqFMgABAOczglwj+cRJMlODPpWy2rMueVIpajo9MXk2MsU3EyPHXMcjukN7
yPILFLRApIaXpOyaJzmWbOKB6PlLNusQkRbfBHi3e5IPZ9VLUK7vcavb/z0EX0b1QPgrF5tC4cee
rJXxi+iYlEOrsNWNQUNrRDwhL4lZ7vAGwVtPZJxsvrurld1HyqTV6A1QP/+vW52liOpuPKe0rSsI
xp7bvpcre695eJ3zXpihKoXfXJSjgMfVDkjDHHN9DPhl8K9brxvH2218p+LAdkXES7LhGWaOb+Gb
jY49iZ2EETpV2edaVShYbzSgDLOdOb7CkfSLd9BpWZsI31KuOCzr4XCOjKiyc9CHy9I/K1HCUhr9
ABa90zm7TmuJNlb+JVoxcqm+GESqsU2xnOOYPK85hQE7fjKBq5Pvi7IglUQQG+hEh7B2ycQlp+GJ
1Z0rMbmzhAhUxq/gRnhLpl2crcbwJHHaWtI1IN8PZL7TzQtCjRi4VXiI9EUtumKp5PXQD12RsNBd
4SEQh9+sumiLkKbBAIJV7fuB2cOaIdVgPTinI/OBd7b9fXbNcrXgOTv2qfmJqEjFTDFe8TFNml0w
FDLUow+zXk2KpCsXmJ+XksAK6bujnjK1I/xPHCzofm6Fezc532A5gHJ6X3LtDtySDAQBIrKkTpXN
MNUwltnnoP/122WEwcMm4roIzhOpG/eR4zsV4bnr5pHGOEyX2KEXLwKgURIaPAUQKX8eA7KS/Nsn
5Q4Sd+RdflOvbzcLIBwiQqNU3AksH5TdUe9MJY3amVtI5xzLyJpehPn92bkIqKN9Q45mQ8F4d/ul
FU8CcuBZMqNZEbouuqbGPwyuAO/KzpO++8c7EB0EJAJ2RNQltQHXh0E4tKaqBE0JOX2Rdj+rJ6Qk
btM5VzsS3F2FupPWCxMp15nX2nnfKssanKo1ktCnyf604AKVIEmHyZN2+X1okRd/RKZ5o27cs+bI
wAu79aIceOlvJqrzmwkdTpBMeV7/ehTsP55o62v0u3mXKOPs2fw///TZZmekGWeS46w2CnwDqXAI
5dhqRygEQrlQhOE5TUxEwAV92G0UHEZ+DSxfO8NLtflrU+oqyAPSeXTuWbCpG/SZgS2dzgqknZ/j
SAOJ2m1CbQVGk4h2O1NOKd4WX0/ZJuJFClFHKvhWk9ySYMXa1+5pfeOiz07BV0jh1QM7r1fh48xH
wKpakOHsTSaGrZ8fXTQoiW+Hr58uZudUcn08AgXt3cLndwmNKGo285tCKZJ79zZOkos+n6EYnuVR
7jNZdspTHbQmfOXPSXzqDYL+e2Q1xKojADER106hccrOunBxdPHTDBkkhlZ+EgXYbsxqp6P49ZcI
4880Wv0k222B6bXqRXbKb15rkdsW2f0CgUpykluLB9aOp2+W3KHfi6MpW15rUjMmCM/wRBBEqJb5
llTdhyoXgspUVx4qpQxXEIgt8L4jnQTXK53eUHRbdFhJarBLQnceUiZsczKrneQYplYi9nG4qRCS
FscEmVdMdZteveisnJnnNd/gueseS4jPybzVrDJRoVeacYSHF7YWHZnZs0bx1zYB1qnIr9FHijdN
RRIvzu5ENlYV3lLvIUuuTNtsck19NG023CIMJHkYUWYHZC8cLBLodu/oNfPxu9cj29oy8dpayPUr
BSS5qkr3/1Y3A3ogLls6Tqi5ZE0YC8OLz1DC3ROD71yWk+YNy1OFmg98n4tZJ1LevAmNqeceHEpH
MjPCDy/sNn75/yAiGlJpVEnIxzMli2D0BluX0R2Jb3ZyaPVZiOJLG/1s2MJMSZzFzDITNcHH1ALl
gZ75h09BZW2yyOTAGNbWPBhkxGiPRKWllodgF2FSTMoLTSS66OoL0iggG8PYX5Z4jRq7c2bnyxh4
94XMG5VjNbD15nbEj/6AQYEYC7YI4QOPA1baSUcX38p64SuAOvCU2TqdqCRg0Xa/67KfMr2xf1PE
MAagZeXAQZpqdqLf2wjC2YUdmr3eW2A/LbShEy9rfyuvms1jlKptTUF7nesOh20p8WKV5BlsWb4G
m/ZG5Z82EH/x0zZf6/sJNsFyf0Q4Oir05+z3qOGf0D/w1Cid0twlL/gnzyiEya73Rd9pRGa4jtDB
uX/iqvcVgaMa4aVc6mpJbPCgtTgb3rYIJVN5ptxj4Ull4PxZwc4ArGI+4pxwFTla9LBmpQ1x3cVw
+i42N/dNYlXl3CCeG0NI6T9GG41Hij035b3iBseMkrc/b/393Vf85U7iPNBumSnixY0Z2bD/HXyp
GueCAyTUxftw+rBuh8jaTRl0NN/eExTUHqTLCH1qlTBxzppGiE/b5Zq87nYhjJPSL4xY6S/0LNDv
TPNV4nito/uhsfLyV+80JNQUrnJH2yeQD4hEbsdOmNx+zEnLOtsvbykPJiojHVjZpXNJ5Mg6SF1T
0Iq6qjZYgTuNvLuDLB38m75K4lQyVL1VN7RuVkt6T18OIV2w0HSWIlsBAErdLrTM5lU3lpn0OhC6
MkFOGAFXj/v0lbQ6LJ2M3O0XCV7CDrX0zjNuD8OTxXyVSS2Inr2m0uXVtjK48jl2PLMDCFqlhbdK
wjUpQ1cwBHJF+Q7SmoGoiKq8z7fKmk7mP2MuRNepqNh+NHQdJDkRdWJcgD4ZL9qAD/mJ26I7KePZ
BIJcnEm1gCY+ZSXz/5h24aqpRf9Dcgq+ypt8+L1jF0kpRE2QJletxqKIXEu6YAaSH3BJCPHNLyHQ
NcbHu9L4JQ5MKOLglO7hntmGI1T/kOz8qHgU1jWz+IA5BDQbei7Dw9VqnYRHLVJGRlb3J7u33hra
kW5+VV3ZLS+jLrczrzIQYusZR99+1m8rp31aLrvM+RS42djT5bHmesyH8PF2WpG86LJIdCg0VDel
/ke7KFgYAWbgA0JxZHGXzsr0ziFNslPQSgJ1G9I0OyMr4U8RPFIAsZuXwuI2ZnZwPgHlFddnBZ3p
P72/cIeE/NeP0ebyqtza9pd2Faarqif/r9dFpOPyBnI8Re9a3FkYAGMTBW/kC1Dp/UQA4SqVwnJS
kscZFAkGwrCIZ/noLcU1pHJcGaM1KCLGaLIg7YySE0oytQyTqQ2qdmm9v6dPTQL7o+tiZ0ZLjc5T
YVT9AiTQF4yCYoz44gizIoDPTJ9mtfvUrRStE4Sr01GD6SfJwCGe8JAUVpbvQj27rjF1KA2DSLmD
kKdZ7JAbpi6w5SjGbdUb4floQPCUjmGtf2x3G43lJUglDoRDD7fey22UhUlkgXooEwtXuo80YHB2
aofP2Wvp/7Jb/7ufgPtq8qj6Qe7z6egt7EFzr1lQbPUil9jiaLIuV8A/IVDiQcIW+4NwGff9pTPo
EfioCg0KdSJndt9PHx9U1xG9qtG/Z/9kj/a1YObc+jCwyHksinzRLGLzmJrr9ETcr0QPvv1SJ3wp
dzrJ5pGZkLN2UO70kgOqjw1aioBkJRK2nT56cHzMIcJZRHrWepUSQesLo3cJwG7cMzW8BTGcalSd
5kw/6rk2IHRS5tePVL+pUHNHnZ2cDKEOiBtCKlmfVctVag5ZcAwumXbaDHXXe1JoldIwt4gDmW7P
3bJJq/pifnNb+vQM/Q+Q2kvH/OenpLOiQ5fZTl3inE1b1IgTYXnKqif7MKH36kmHzI7mAu46WyZ+
klOa3xKpKmPKfg+ct+ECOmn4tSBfHrrmXe4pEtG1aNWNNAfjv1lUIKTYuyNJTGoEEg5MUmOdCuKE
/g9UyiVK9618ra1D4k3kjr4YLVlNVV0T7rQ8qTI5kK5uYMiyAeGDhobxjrVx0wi5Fkg4oMCENzu9
pZq9jIyCkDHTtqY0hY595jm0FfGRJL9PPUEpzqah6GUTmpRAmMcyq7VMbV4gxXg5juxGCA4AgEXD
cWV7svMr/BItou4rGm/zCeKgTkHWl8/Rd3h6ngz3JdP1rNZnxwRHyFi5hxgJhx960PMOyq8cU81N
RUI1BhN2z/amMjQJxqGUWSLexXDB28dk3swNmn0CSaM+X/GnK++Hk3lo0KERl0q2nLuF5KW7yoeX
mJrnPx9Qs660iH86Q28kIqAHT5THqsSh30ckz5CPzO9RDHqoTPSd9mzb9c6KrRULYfnQQ5zyWPpB
3RwoGx4Wzepfnrh8u0Mvvl8qYxlcvA8Em6+IIBKvsuMRubioOdNSez30ayh/1TkX6xK1ctqnuToD
N0ECPBSK7ArQZh2a2dj0joUTBXx1VMSlllEIYL7FMVtNQshmyJDZt2+DaSN6f5nSJp/tdkStmx7f
0KYtsQnqg09pTM77y2JJ7jXneJOegk2zb508qVjY15XOa/gHvogakgKSkG0Iw+C9XEUnaMGl+R/u
/pGELEfhKrqmzLZmsBUEHMH09y6YJE8OvuEennK/H4PMDWBZcCIMN9wq7LzPZ6nU8+QA5XLRXqf8
LHGjEFv1TCti4bwwvLiarkO4SAYvQa2aoEkiAHoZbUN25b5noVqwATGEJhY3Us4U/XgjzbzIhXau
+YuKjY/WDWFEVgz4tyiQ4P18b8APknKmbvzR1d0ND9j4vtDlAjt/95oTrG6GMZJJoUStZYUFRdqE
8xaFKeYaGeTlor4CEDUPNVqIz7ftEF6WeYY31EbQYz1OhnOQVdk5C9avcv5m+9KO8OXfolxg4Wz3
mmO1obDUnBI5XhqDVB7qx5lbbeEpEY7gb3l9gZJZhApi1be3ziNPSbmqU2V0jiVji2YlOZ01yQ1R
nclmgh1LWlEpJB0zI3ZjcBbgdddizha+e/7P8zSgx4Wd825VDQbttNGrXoYzDzV2EaabNl6HYOOc
MFB7PocfkxmjFlia/Be2Yjgis5MWUItSf6pc6Ldia/F0x0ke3c0ONNnf3d4rTOdXSr2oVIdOgm0Q
mI0FzwVuOI1EqoZp/iiaynfAyCe2NtVUpyyQRPFS4bUSYzXPc0BsLuVe5+xU8b2okke8W+jmWOkO
n779CWENA2lM8OuuZwScbAiCHKkjslQf+ssNriwKX+TdkftVgB5CXtWaHVqXJAE75hEepA8/9aqE
IJotVy7HXt7DFu9wBLQln3dOEUlWzhq0L+sJ1ZI0KqI08mOFEAQXEdXedqCL9uRE7Y54TR1Sg1LP
7f0UeNgJlowPSl7aZ8OyFdD9Ptvgjkv8n+l3ieaIT/Pv2R38VNaFdawAldDEqjDyEN2NYPNJ/VgK
iYtDMWOveqsncZ3jT2TUjSfOg7VwgY0AbsWz9P4pv/7TKX5cxXGFcUug/OAaOuEgD82Dxt04InBd
gNVvAtauDDhWl8nSqZxKoJuow2ubpZy41HEsXW2MJAD+UNB95Ze3kL5pw9nX0xmjDxNzbl41wJCh
rxEOHrey7VYI6RfWu9zCDWu/JlYFWC7Bl7UMhFnPu2RCjgzEYAMw8wvLXT7SuEy4PZaS/7nc9g6b
o00MTh9N88Jr3JvXgNRoPRrZKYVlPeP0pdL1jT4jKDPRYv/XyeljnRhuKmHWFhf5W8v19mAAMMu3
2eNn7eSM2Cr1Wq/KPfY0e0J90Br9uAZts/1ChotAj4gray9YFuz+EuxH2pu8Bb3r16sFh83mDsGu
tilw1hBZntigDZ9gjp70cD0R1WO9Jba1iwx17fAEL7fIFkDdeSw80aYp09+AG6o5qlbleVdCRIgY
2627F5zMEp4NVBRovmTQQdFSScdlu1UKab7oBx18hnO4pwxXiwlolArdwMy2ZWVaFSdhi1m4Eyk7
9zC1vj1EcaDVStKWUuAJoYpGuC/ubeXGsoWRa2ic67KvD7jir7gRicJezDoYGXoKDiclSVFesAOk
I1K8+YDQG44BlAKNaxt9mXfhZliah2RhCVcebWqMaMmikpzifU7IXW6DyvG8+aQh7L2Eh2P1QSMv
ddoeuyeq/sXw/1L3Rg6rO7SCt69/sBZ9NGS4Dgolmvo4xi93p79i1M6ZJjIoOs/RDpqb0hM2ic53
9WnhaOkstApumaPx8EWtQd3y2Y68Fw9JdhEUIiuJmVufd2KnbkbrNlJzFPZxZvRh8vI5JenAtEaE
Ei57G3a9wcKqoEppbeV66BUI5C9mzSpXhDZ2R6IUpfsuRUjDjc6nDQPEFzEBlchYRMAj8w/3hkD/
L/e2DhOU/AkZ8UUQgDkhm4+ubpLTo5nqvkoNX7Ezy3nfxBPBHFQueg6xAB9TU1PmCQM6bydUvMT6
fDDN1cRXFkj5di1SH5LgJnHhUcArtd7L10vng15uTcyesNgCX/Yw17zvkXz+jxYyVeUek9KkaQSF
432VClpl9v4csasJrKcga7JXmmiTxyOQwaY6tqzFYOpB/7MxLprvPEpdvzykALQ/2S7Pl9ym84HB
Y2thZU6hRzKvsokcM+iRrq9MGg6iYcX+Xux7cSHD8vx5E43n+L21tX4mZ0iWvYsDXZ/t8O3MHXFK
5P7j63qEH1xQ8oYf/De1y52JpswGsl3tj9feUpP1anJ28r1H8gyNS+35syqL5UToM7Z2sm1cMQib
dyNRTFMIKYOdRYBcx7uWZUqoYnBA46hOoyy6R1x1kpqyyobzkiPe6gunK7HH/To5p5TLnab4qbf/
7af5DjxC0sJ9Ao++SkkDDShC8BaJkj25a/J6nKdQTIJyZet0kPL/q22tOU9iDG2hS2o0Y3LTKAuH
Sk9iHPYUfbTCyflwtB7FU7SDEEIrId1kz4nzSHYUAXILK0xUi4e30ynubL9uZuxAn1EHra1GaG3O
J+ejdxEGjs9mDPAje0GcjV07+c48jPSLQVAD2poqnhokZ5hkVYyL837MA9TfHcpjIqitsBcYCr87
BdmMk7UoiRH93zocjaHxRUxHNIjOXBVcKPOnHW81gTF3xJlD55IB8xJhErXQ7ItaSKDMvKQ4Ofmh
QJKg+GoCy9V+28KvR5xyjanLsEoWPwYOZW6vQROU8Z+vzjtsHLRVw0bpUNbkbWhBbUeEJG2laI9r
dSRMiRdC2qJ1a5ayYVDyW2dDDPqvtQ59AY61zQXuEnFyhtQ0ObmhFu3yf5TTMapZjdIRTtuyDuwa
F065yfxenVNB5zJHsG4Acll1ruHHJqyzj/Lx/EwkW9mttw2qCxmeldef587zUZzwpYHJlESJyShp
FPTSnJ+ZJZLwMx0IixD6iA330Z9kxEbra46CrnEPOIMv7PL7uUxmuoYgu18KfRr0A9CjtNh+HLWY
hLxdREKx40Nc2ZUwFp77aJnYrRoH6MjesLXwRelOfaA7hJCbOaC6WtqBmN7LwrC2JUBzEQLDusx2
wz0Z+C2y9tT5LlA2l2wbx4VjdvBFYo4MgxIp5JazwST7+bYwnfbQLAxsDtYnVNY0kqS04eNY+7m7
lGanNsBJ6xx+kX3rt2AtJqyRTs4FlEtmSjgGIMAmpCmfufRFx0Xwstn3x4vrswx3OyuIzaxpClKj
761YD09LqSCuDQqQ6zLLqTLA5VgxQH3M/bFfudwFsygsqYMqnxRvIpUg3iKGoZ1Q17jFe0QEWwZU
Bz5TDPHxWs9s11rKSqOc2PZVFmTjx0USHmNEy6AepBW+xRhdNGTDGAswdJNDJXsrHJhdaUwgU6zv
gBfqooJTA96azhjKgmeku31oMNGmdDJuaMNQDW7QUkQHIqduBzCZ4gGnULMOVQtjYfZup5wap++A
H2jklkHaJn96Ce8EkUjtJNEH/1wMOmAYsuF5ahIFTItGN54zen7sLxNrloGKibz2OLjZNUpsuiyW
RUiOyRz8w9iOiiXlJ60gPlpeWRAQQwY3MlXT4qB83j+m+RcjyAcQwzGgLSn9nDomRzmoIXq1FeNf
9kLUopzDQlZVUVYDwqyTeikP+Rnrw5y9GI0BL0FewV6L3ko4I3XA307cR8In+kV1vETHrm5fM2q+
llhZo9Q7+8mRXxN3qIJ3K2pO7Vn4oUy5sf7QPOSHpHipEKv8z9Cof/y36V8noSk1M/gFv31Y+x8l
/EWzvuAJWiR0BDZiJ4X7Aa8pbglMElILjUhyy/Bx9bywMM5lI0ZJn2A9uoTordx0Jzv9u+CaUiIg
c3cCBiyR6w5IxvCGmwxlGU2QRCgZw63OfBCpJQXSIL5wqM7tRM5SjitksiJ4HpHAGVKaqPdbAFNH
OPDUo/YihnkVUBJM6M1f9DEd1NdN6fcKQp6eot5QB93vp6gdRxBkZSJp/UtCtb973MSBGBMBvR1F
KM46CZsfLAhnix5ixoZXGQHBLuysQyUFZJy/zFSCs4jpuOQabblp3ftN93gtvoDiUaRUcxkgYyAq
5s8zdQrVQJTMdQ0c+SlLlMAGPeZ8btLrqkUEcpklGyGCjf/cdJumQeZZ1P0pcYsbIrMZj/QwIIf3
ydbktJs95s+aenlUTdupUcFQBnUkB4IFqfCB5H3AwkKU92qa5bvJxC6AR5aOLmpkL5nWlyVH+FZk
vLCNfMQ2cC+3UX8cwflNffdfh2NI+EaNqEUFjuFjsoRZeZXVW5006Ax8LKq3edv/r+hre+mgQriw
LTy5qFHDhclM/YmXA9vWy3ilDPYW3DtUbfGV1L1HKiUc21SOCvODxNMNErU8UuTD2HvZFexItzVv
8FYMXnUHfwiCxmbUPECdgMvR6hw2Um+KXE0qFv/8Nkm9KIHy1FtMbYeIuZDQZ1A36jJfR0HMAFoL
WFhmY3roDh6soy0An9PkuNtxNYcDC+PXZciQrFJ4WY9bKa6Z5fd8uOZZG30Efra0Ttp8p1/0Tyh3
MUZZnnyyV9mGugOvAO+cZEt60y0Q/QPuxzXEgmdqFDwWJUfwYe/w8yOqAfxGBZxRq3KmXlvhW++q
Om8CZpZbeGsVLIvtIMlIPCJtsaU2mhqWtlkkwOs9gkls1HcekSURniwCupCxdWbKxyuywjpwSweg
0NYEQnyHwtIvwkagWvxNaaA9qyclbchZKw8Ibt+s+TttvA5/SA4V77Xmo/2GeyhS6OzG8I1FWPfY
3Pg2bsAtwRlJa+K8fnyH9OPGUmglnGWJIdKdq4RP0K5/ykJAFq/GyAdAhBXokQ5DeuYnM8133Ues
5uJIWwuPtDppZlkfuxkl9IMFziaRb6FZKRXZeuuG+rgoDHDVzq9WP6Y7XgMkJFp0gIIn97mGVVzb
LwHWkGMIZ+G2fUaXW3w36DSmc5mopgwTHgjAIsKyfsD+/UAO3eI6MZaJPNoDkS78GOG4izju9z2g
+yM3XxPpeIJIIXn46Xxc3gpRynWPWSnB4TZcc0ypsz0ASyEyF+QDIrvxbjiDVNMcjFo6lPrRIsxQ
5S2dVmzbI3DOg7cSt9wPwwtN9Ps159tIskqUasigQnpDy8wGZnTOxr4eFOxzsQQsgC6kIubMU+aK
NvxTfelCEJUkAI18UPrqGZ0l1/GvFY2C0bGfZTA9QeuOBn21CkRpjTBql4mZ+HbKg2YE/D6y5om2
g0fHIC1ITSQ6ZYMM7/Xzp4Dqi/5CE9mI4Lzdgw+vTjro9vIZtxGA976CFtPmhegiD/tfDumbk7YR
Cy98m1AvHsrplm8V8R5meEPyjAcyBwx18BWUyPec0VTD6orQQK8KFh9eLbgyfPAPanbNYbl342Fr
BUcse6YDM74KPGnKr/i+BKPtBQKEiIV9Bal96qhyy+CpHvHe/TmcSaQ6xG2E2Mq0KcLX0ySkNhhv
TBX2P9co3WWDldlH5Qbj4saVEcEssuOgmMkCtxf7s2Rm9D1TpWcRBQfWYHPZFoNKFmPgymj/Hu9c
WPejQN89B9AlrP3Kkgy4TNBHPCgolNI+qVi24148WPzRW4ODqieCJhKOPgtaqwc4w1sSQn1kEXSf
4OAyQcFYDxc9CLMQGO6D5FUKVsaN0js3knykkzLF8c0EZNbDMTEJC2Tl2/atoYp3BwoJysE6NZGt
X4kE5NhzeS9IvkT37knuIW5LgERtV/xwrDrdq5uRmMeSAhic0+QSXcjO898dDY74o4/LDGy6OBt9
B3/1kOmGnHFTmIdSqL+DGALqVNj5Irgy3Z7BJGGzmXtFRQRptDi7+YKYeHE2e1u3GgJ/PNMoyev6
EWHENYgflg42JVRQetRhNkozPnxlcjktHbemTBwY/13vFb6ftlA523rPNw5j1iRYwsEGWO04EZZY
faIP+CjbnpKo5HNDsBg4S43CwTXEBOUR1wWqeOG4ba5GplJFgUYKHG+BwUNmSjbcqWxsF6bm8SZu
WrDywA0vGGi29mj02UmAeG/gqyPg/5xC2atUCxIdMT53X55/UUBwT2mrH61tjQK7pR+ZLqTeQdF8
Fl74O0fkYgm21WC4WlkerqQYIMFWDOUnEnCZrg1POm6Nk0p2eUFZgqIlZQC02BVOqIjXQzKlgZBk
TjiFeVdPkGHwhmYisnz1PT86uYiDK6KUtreZndKWnepx9tskczxSGgSQwus6bRRH6bVuU3Hd8Ykc
WyaOMJhl4+0MYGSeLHYMiaYW/Cu3yPH0FTuSmZ9Ya+d1+kfR84FeYaGyCBj6hSNCMatNEZ7/0JD+
OOgMHys6wW+h1OQYVwxMFaUb5oiJoTG7pwVkbrhEjOQKhAPqbm1EKdht1EEyw6Dh0DTIHrJpS8q7
DlP44tHrW1zJTXB5wxWFt3fnPn98Kf2knsM1SkWiJj76AaRsHR0CY5rYL9zAzoMIkSb1PINhnyMB
guV723afAeM26mtLc8ryXB5KAwmp+f1TvNSDThhkGbCNTjCEUcgAupZau4JG5TndcrPnfLFoUhCY
UjDOtiI+QgOnZNHgUHQUBZqc81S3LtXIbC7D0vROxlnbuDXVLHjGnMzTRYT74as0DuVVYECWfYqq
BhTf3fsZvZg0I8/oBSinl11/K5wgR2bPwOVs0ICe/VSfBTtn2Al6cxPSo78jtxemA1pUwv0PkE4H
3diHW67lLYfSMIs2IaVrtxWCV4AdtptK71qzlbcqQPG7To4FZJUea+FEdpiocRl89MELpfb87+Du
vC5h7WstgUBuha6wSctLQFysHW5rR1KoxzxPz5kvJRfVZsDv9WU/RQjnc7iVbRYm1pkT2EAMVF2W
Xbhp/SQApL6nHeqokBAIMVJqKTLff3sAzoc1NEg5v2Vr8OMrNPEgTZHdTqQmjwtfRh1eayhFV4JR
OxReaQv7IU4jha6qkWpSE2Cr8LLkqWVXfRLkR+f7Gwpvc1NHhMv9TEC2sfc/rb05kNedzAv9SKDZ
8zz7kpJP6Nl1MT6mQNvtYmC7Ym0yjEy2LE9TPfZbOkAhWsETCwTW9ECfAe8anEvebiz1gR2Bw6PL
+ZbkS+7DIPJrkMOJP5sdAzdmD0ed+gtNZD+Q2le41LJBuBK1CsHhKZNwGsPIAH2dc9OjSmDEN4nC
W6arXl/566Cqt72JoelxHfI6yRL9PNtzJlP3r6x6obFxy5Q/ky85LoaQ4U35hMmgtL2WvscoQWIo
GBKpVylwTvHqndXn/oQOFWz51yQyYFsPQki+bJRUcq1ID8JBkyQVu4omL7HQpWDUHrPCYC0etYqr
wa45TkHEkTuP3W2luoupUAWAOx9hQW3Fj9D181/2SaLeTJPxoiaFsfCjzM+1qVG9kWZz7bqAZcMa
N8vZJFcVE6iVG3OQl7wDHtDdTIW07yHOVtA7OnBjzc9ZJ22znBUkDSq43f0wD0/o2OLw9PXmWHKd
F5Q26G+aw6+dcrsb5TtEFaFr2KeeSxrKmbqDUjklrnnF7rSjlLFdeCu3cMAV0HsacvbycpAa6nZi
m5EnrSyXr4aboSOLjWKa4eWpsz1DBBHSbSShXJGS9pPIdCx5lASnQHszfa4sV9gqyI7nP8WDYW5m
Oaxliq0UIoqXK3P8sIRbqofp7r+ouXuaJ0TJd1MoC6Mi0InhfSaDQC5e1BUmsc3+idkoIDSOSoZX
+Z0GRis3Dll9I0hl19v9MndLO34NHni4lswg+86lJZ2uhNPEM4EHhMSbIiVuG5/RyJ47OK7DS571
ElIyPN8v3nOmhASEeCb+dNC7VQOheO/aLxXhuIR3AE9alfaIBpyemfgmYolBH6196JvoTRwUqEIr
2G7N+jzHeEIArAD6oxs52cQFLv6vIox6KTUBcpRyf1KYcr1+ftK74EzgGo2WipcaBJEyhCOr44lz
KXrZwHtifkPB3d+Abm+g6+011XONjd9xpfUGf1fU+8i14aZ2zpXHLsJJWOkcvZ2mTNqsym7FKeZC
Onq5gQqiRVgs+VdK+wLpFPccWfqZ2M2FDt9sUvkVapvEYWEHfLnNKL5LuC/hXQ2dBprMzZqBNGhG
sVnwF5ktPWLx/+D4uHW22Iz/Kt8qp1TruwKWuFyBmvqgwVuLAtf3KqoIfp0UqTr9F3ocPpxOIh3M
lZl+y27LrP5nlRe3EhcKEgNnL1UKWozbBnrNBOndR0gBk+iayvxDO5tojGdl2jVY6veU6McXUxcw
OBv5vC9/qREAZZOus/YO2oTvkXBC9G/l7No0Ni0okgDDscvYAoOn+AQ9iKWGvXF6fD7X0i5QBvqv
cO4PAe9TgFeOkfBj9TMYwLYrylF9A45qfFE/jrqyVEFouGixsmB3UTTHO3zuwCrcGIqeuFXdwgLg
u36ZMnj43HTOxiE1fIw0p3W9vq6WUaJ3+mfvCZb1kO9hhj7vGD27LCgCLv5RPsCzG2kHKiUVevpf
uFiyYgjubzf+26vrosOn7x+fdeGOuXZRutPOPQXGTq82hg3pIFXRAFmv7Rzw5IKmiykPad0mz16x
HHdouf/kqIqDjLBzVSaK66FkIjLR97+m/NBjkuSjaemiDQD6T0Z3DKHhcoVY4JmWCG1kK+cHJzXu
G/DJ4Lj8tReweBdUbsii3BloRML8gKfESgw2JUt6jXW9r5+VMYE2+0Y72EVj/BrXdNAE5iVDGHA6
5N/Ygm8nAkR6JyxYuWnPAptuTxVn+cS+0V+9csOJmfUL+bGnahkUi9jXu2XAZmAgufmtrwhQ0mBM
EqiJgptgjNl83+/NClKu2C85yBzmxiXdu7ph2SwRCpezSrABPlb4wn2lLmRspTWBldmgqKQQd8iZ
n/2ZRqvxoQXtwo4muSk6OJ/SOIX1k5OJnANvecTYKcJn5kOocwbtYziF78qPBGsbPczc7FZHmTSx
oDvr8s7rOePLLfNbJcUHeljnqCwIw+wWSRlTPDpVW99PEpfIyh/1iJnxdpwMwnIZmgswhziGlZHw
4FoJL4ia7IDlBB1SHYzPgZhHqxQXlzFf0vFmiuHXXV0t6UgWTq5yhNtMep09wpfQGYB+mgI72j0F
lbwOqSTPc5Gvf0z9ciGsYBRQ11dSkELOm+cy+0ghpX+zi2HvMFZdcJTt3VF+xZstGIvyFtnuX+My
3+5+C9pWoGcLsk5MiW5GCSPSoOhBbT3xCcYCGwrPqLYNkvDD4KLMYl33z9gMrQmiK8deNTd0Sf+u
YgRWrDvccSCmHKYL74O17MB4avmMIyBjQ6sVeP7v581wGlGJavHT1GGUj2G/wHVHES6PkzV97ghg
nzaPPo4kInsJIpvyU1R05g5AAUVNhTs2M0qWA49jFyCElvEe+3ShPNX8miOG1lSlm7CyhjAdadGQ
7Yn3HMNk4r1UjTWV4M++7ynOBpywe9p3eZ48SRwukDjsxG0QBPOa80nUgnBU0TbyGJwbiXvJPeng
7LSYQJigtQ2qQwmVCEKrMZGaST+iolst/KKyWx8A4IrwnA9udGAvHeTzSfdpQ1OLH1M/Qxl8XdUc
fQYamvonfCX5pc/+eSCwbxvGiBq+2mB1gGGUXA2phcv4lBLEdFfGMHwFwe8gYNVzfbLoFSBDwYuM
tkPIaixA9P6VPjH5iMBiLhV0sqvRQKA2bs7bC9Yy7cR1GQJ3O1kAUJxiOO1B8ijaPnlis+o800UJ
hPys+3d7uT0rSC4VjXKZH7iblcExAIjR9FeiWSmzFok7ZKChg0ylfcS0JRIJQE4g2ccWgIoMQ4nv
5ze/CV76jbBRyyvz7vD0lK/41x3H54tsf2jR2mtw0P4V57ULsLlUP575bOjiwEL9ADhXzatLPtBN
zCfQx6860Cxr2PTWSFUXJ7Wrv/T4oD8YmVW7z5EosYxZ0IiJGRzroUN5iRxlRfXMHDquO2mZX01Z
WTg17Hb8NZxzj5vsn38JkPPmg2GR6fKOTqt+pvrOB4i1LbOzJ3AZ3m+JC0OvIMFHgHasZkVRDo5M
GcitBaOpT31kQCXxRD2bYkArPacDsTQEHIkfP+xcj6Y9lYcODV3T+a/0VYJg255CNhfEk/cT2jzq
XNFUTe8DMpC5eMwjp1IrCyGHTt2775A1Cb3VFu8WmOPKc3TetxGLg5f8AmtupUKjfIk5ndRCd+le
VoRgjifEmx4wku+dLh/fP67kNHweKazF8waW0gnhlUSd7GGcuKP1l/Q9svz5Imdee9zQKaUJHjYO
yRdrzeyGndzj30Qufm5LXwUsT4Q+jgFpUtTQHDbHW/0bbkhSnTBGERkht7Yba4QWVW/rtU1FhK+R
A2FY3hnLswIS7yso1aUax7kZEjNIW43ZypB2sWtASUJhcmQ6dIfmtEM2riu/WqxpIIWcTW55KJ0/
QA2tXY202XfcwHzwJD4llC9Q3r0C5jBJhLIZuMJkkncmknODTWY+wIQpdLONL4hbBr7hSVzxkPCb
y7unzAXGVbwpPDfLyNC4vYMxl03jih9ke+OZ62P7sWCn0mdHR0Tn6wrmrO1KWNB2rKawufCONDfP
iV0gMRCpmQD3PNPbJxBBxrWyjHdCT4HmhK9Qgz586bc/1Vx2lMXWP/NIkWJtWcqDD2d1eQm+MgJt
69JTTQHZGDzxDas5elYDqtLe+WwP3QhjxRDQ2zh+tJPGrJVftGFLPY1kXY2ED1r7ZPlrPmUbY0Tz
CbAOw5wHwpKepbAyj9dF8R42ucaANVsdgFeoA0Lf/egd/KfgFDBS5yG1BQCxMtfApmIGIV/kY31S
EDkIQDYVDDaoK9lWmZckKCTRWCq5Cc7O23YHA/Dcqq6FHZDjbZ4Ut+P1hwQnirNwadqgk2UwfZde
IeUzXjvztSAxNB7TUGHj3Ll9rRCL6Wm/8mutRI8W1pPpZNLHzrsN11Y0UGw+RE7wy5gsl1jg7oNg
CUCUCqko/hccpBtLlhZNXB8HiN9ITN+BNSDlUsanUjuMkKUIYws6OmQRN0BD7uzsSnQmZo07vHWC
Yf8NLPXiyHi6LQFadYX1pnMh5Z7wFYh9X3JRBEghEaL5ig8lHWwH7b/GaeXjPlOaAiJoTMC00/hk
eQSKXHwpnAFWjYCx3DmzY28AqHw+CMhl12pQxzI2IyknKFbX2YJ1TMNrG/jobAEPJ3iub7OTX1Ne
erjfG4CbGx8ZtplKNT/3fTY9zpjtrREC5Maxu71ug+l3zia8mlyzvuLEn40DG7mGsoUHAbIhAOV7
TAzhk9Qbg/+Sp1wEZ1cOh8x9aTAjYzGhNujaH8VVs8+DseVpimzIux8SsO/PIuadS4cQEaLXolPE
QKXQhVqYGjwWt/iwjj7nmWIBAbohINvDVHgbE6m4hRsnRv72tFeqBWUwou2hLrod8xOQAZ5TXTlM
ZXYwiruLtX4w00aECydhAShsB5bFtbxnzslQHLjVtQAb9CwILQnLvQvmZZ/aZ4xO1v0xeoQE/daJ
jFkQC6qipfRPxCaqNYC+h5/ErlmZkUOigsEI708lJy0Lusoydc1YF0nu4HiaUEVd1pqxCepz9sjt
tUnrps+SXOxvT/Z4AmExjlNn2EoQkp4XaXLf6fQcpHKusXSqbNbb09jYMsCuKjXeoJN3h/w0BNTV
IzD0qKKH0/9KjmmWuV+r0St4DHeFEkf4eQdciSLXcaqqL9WHc2XaLGxMm59sL6SFjp1aCdGU5431
hfx28XlwjuOMuHaxEeL2dnI+ROYfJebNtEZKAk9LtCL1HCOsR+IT8JnQG8oTKTmgaHYpLBeGYZqM
UkxJipC34COgzhuxgPm7fbQqVf6zShjVQHkb0csmZ/weUu24vY7VJBdFpA+bcY8SaH0Ruo6RhgNS
CkS2IkdZvitcR96V5xiAPDNiodFQ9kGUKgtc5WI2vSeKWtG6WcIhxLeolA8jC7YZbgqTCEcf5qkH
1sUc1NOClBuXhlYS74bL9s6/rVnpeRbo0QgFvhanfaGpsWOs3qRvomvdMsmqRTU8fIeFO1vqSZwS
WSqMrPyyIkXsOG8QnUOIq9aBZah7JuWU746u2cjRZfb43VZ5fVareuw6p4gcUdHVDRdJuuMYpsVr
rPwKt0DXpfatA8DNabspZ1BXNcOgwcckqThTYS63ZkbOJuYWhn1qL7A9BTkPhBQAE3L6Tu2TR6w5
Gl29VNZy4zE0vv5EvbBibDHWuRew45WObGOy3Jnnld5uZ8B0uF6DqhdB/FhOT91ZLIhfyP3hzoea
eJCCDfKWyLD0GD2gqh4qXW1a6Wqsc4wPJFVmAkp53KxlP1N9Vs0ExMiG5JRRl5AOydbqiO6dPhDP
sGG8xRUQe3YCf6LpLR6Y2NTGRGbWjRWGVkkyA5ew8YzSF0rVwzVWbA5R2nizbHVz1aY6pbmf9AQK
4q9WY3QLm/eQtQqehW13wZ8Ye+aQ3TkHIyQ0ac6YFm1sTVNVZ0UEW/IOtgS79Sg1K9uGOan7JpQw
dMfxT+GkFYdQDBZFfkD+wlSEZzxF/g/mS81GWeG5RDCjK+LFQJlqz7b04NqvZDNUfeSpAcRJlkg+
naksn7Akbb3KcYist6QBgkYnJHi09BJSBL7cqWUGyVipiSR1ZEl0Dsl7c/Xg5rI8cUotRLqPoURZ
jfj3Eiwe52RbklG9bsR+i/UtopOOEB2nKza3tYEcQo8Hw5Ta4kMR4WPglRa0BqehBWAHOFfOkYRR
WWDWxHjjmEwAg76gS1hoCz/u0lrjM0DC+EwBzKM+4On+2chyMtHu1qyed6ZCNsVIBEAXADVJlHnA
mrzsHGmQiBmJ+2k/031SMhY5jAauYSJgD4NORUQFHiHpyg9/cnb+IH63GNcfauP/tdnjVIavctXq
JxvxlHsgNItmPbgv/6MvVKuPr2O0s0UBIRRx36+Msra+7oJMPUI9hUGUOBymw8d9mUzTIr16qn2O
leyjv0Bk96xQ5yy/dIfCBAQ5mWWzWHAT4Vxxjb6LFSK/y5bA13M+PORkbvx2ijD/ChI9ldCdSJoR
RQwVKd/2X42yuTTtrcistme1+PgttcU1HxLT/cAW9rTSBK938jnsQqTOOIuVZh0aHBMTZ6zeWPJi
uTLOSAb2kD4dq02yhs4taLodMciy7jgahih8h6NiKVmzIKkmSLyEcLrQkJUWak0tCn2cAxgGKGgs
NYIoffZq+qMY9ZaCJl/u+GaYTBmUV4PD2WeYa/HqQXNm21guz14IA7W5uFsDDjvQ7hR3UoPfabnu
yI5yLumAga2fGFroNbcJvYSnsZiLH/5ai+z8DmvolLIVQnMSRdatFR5o/T5MK8CvMEa3c/bIs5wo
KKRrvXro8T8X+qGnuHXoS4lLizu1PQzJYPAKk+VBIyfSS0IRKpgYBo9iJtX/IHk8sY7xod/onoAG
yIjdw9TskpbOR0kvOSqOkSwqKqJs42uEbTMgdCrRSNSkFkPdWBWZlX1Sfc3xrs62b+X7V4vM02WZ
yCODDI5lWs9/Tma/TBbkEDvPz4JG9luO5rqNoICZH5W6Lp+5mMLaiOyIFjXYilgGB3UgVu2gy+YR
S1DTHaPLZ414prdSNVYOpns5OqInBkxvSE2BjlVzHSPluMhaDKMyyOYe+ud43cyV3ysuhUfSIEem
IKB400FWhnPnZmBmupcx7JZnCk0iX2rLQ9w30szzABPZAVKIU2pzUkKu1PBRUyipkkqMnPuX9pKS
ArFWH7Vmcsh1jKDafEATn4BW8bhPihahFMXX3r/e6F8eGeloHEvjzZRGQ5Y+6wsaAWhlAH6Ty0S0
awolFiXYlvkGYsiY4oBJuLKn8v71bZLGdfLYcjjzGjZXWpPyzdv+0J2CyRfa//MJJ3seHS3Fqr1J
q02mYxmeQFlqPPMCsBkXoci6CGRPkdCcIpCu3ebf8BfDRf1s6T9Rwl1Xdug+Zu1nFKVQ64psTqyi
1DoxUhYMScGa3SXIDB9/MUjqhUYXogr23OFoLXwkDSRCLVdkYnLVisKu48c0CBrHTGKb32sW335O
nEtUl1DdU5TaGNTUchhoweRI1msiAQFlQSu6HXKMECX1O2liv5KlaadXCsDMvjhANPWO4oLEAtfL
yk1uCrnEx6rvz2oVRCdST6BaAP75yJZyZgjkk4vNae9/5mftHoEZgF1xR3ylgmWJ9+GI2g2Xc2uQ
2Y0DLyFpJOnLp0nFBWHALwjEu/eeIdUZJcvKy4xu3E0l6THcgZUp1GeDG5HsC8/Mi+3zhmCAKefr
d5L4HFpC1C1qBtjx71E7LCnQI/U09fPgujh7HJjaNI5ZwFH7grGlhdYLyd6AO/+b0f1kKbWHjOFy
+jskoNKnYO3Kq87l9qTypadM3Q8SRA1MCQenESOJwZuCPKPNbme5kmpjsSYADf6xllYgiNkp8QlF
MZ10T9Ryrcpmi8AI2VY1Z0mgTgCbtF7p42G/Uusa3wRJwPNitVWO/7H3nfMOZ98ZJE0/q8Yr4DKM
cXt9j1WuEk+hfMB2PdOAQcYEtU23rkKjHD+X+snCLUpZccarKgkCjRjKUZAlLT9K7A7OrZBH0RsN
rsH0A3l1ImOKKCHaq3K9Y1y9gtuCb0lbCYaA68dxVqwwVrxxgFAzpq40hMMPdkc8V5gTexUC1Owb
N8Ad9VGtoMfSarPK/HaaNgWkqx23cQ5G+2FQEwihOeMgTN0qItBr2Wx268Comlnx2Mr2HtMLB0OD
6Uity4qSIxasGS1URP6tKiSGutLYeQLV0FTGD86Ry0UXGvQJb0r68UrflGqqH4ldIOf0WWj09cxq
G/U+8X43LUFF/+LHDl2HOQ2MwC13Tz+DdTil2JyCl9tp5jSgq2+u8jFTx0xna617lDmIBZ7BvYSH
70cSbD+X0Tx0YoXtCrjDvhoifjG0WvnPmsJBbZ4ll56lN+iEOiBfM6BAeI+mp2ffqOn6p54pI68D
DBHTWJQbvSKWH8dR5KN3gImNlMMud1kabKU7HGg9B15/YyO8+jQdiilnF8NI6JORyLFnFx0hlitY
nQqsNIVIw3fVZQcxtiF99XVrRaVtL8PMKt/5tC4mu8w4nFV46M1vAMVgUiBSOuXF7xflnEcQJgN1
RnUFp0OX6PPvKjCLnw1+JhPhp02PP1IQeQJ13uHzKcc83v8dHlQZCLglmBDvkBZWHJ4FgucBISn9
oStOGkD2r7u/i8f8X4GxD+xVWdbOCgzjAOgEF4m2zN/ARN+7VI6BeDsJ83cy67xLqk60JPtk9hiY
ypPdXOslWPu0x0Dsk54Mpc9VBluYFieNX5RBV5aLHvVEPN4oeevWbRaJk0Eiq5To8Ib8SUFwVzLa
ZLfShmIa2kHeLQWhBuYQOYBiQX76dWDYRz4v8TXODzGKzpjogpryw6sc9jJL8Wg+4l993tVigp6t
IqUEbDmxM4+23fHoUKQqFIhOPvID4bEUO/XVPpQW91faDzhxYB5kSSMNgOxssXc+9KJNWy8KgK/8
Qj/5q6uHf+XictVwgWGlsp7wpDg+Xj39ArHSDZW+X41G52tL0CSW9zNANusgHsMN500FHXPdUK61
ilDRB7TDeIb2dN7xcp6cF4ZOWuhuxhm84eQ9q3XOcBiR+95pg/yXC4RINbGGPmzqCsOxEgAuQg12
sK/6SsX2AeVDutyno+WaxqVU5SBc8V2eIiJ94tLe+Iy4BWetU8iwcsYPeW555cF8OpACBxgFwBof
QPYAKvPYbZ5sWCeOmF63uS/eMmt0MIq8avoZ9PABxSgYHNpQYtiNIFmCDWwXontXU1x+x1xhOYQq
x2jMYXZNXR3LEOEWUldwA7AhytItRf04QuIxgXumR2FLB/flK35QttwanWeQtz3WMOx3lhdXskWX
/Fy3KZZ4mYmhXQ3JgCVCLJsmgEpRTasmEBwy8FrlaXIpXYOaqbb4EBc+ElwgERcDDBGVw123yDYt
sHh9F3HvE9NznrPNnM0G4yVLB62hAz3cpicJuavBYhTzgmWhq8ffaoayAB6wG1dZTV6HQL8nadfp
+NDxGcHdjfYJfD5pMBDaDJHdha4ck6gZfrtus+GmNFNTOrvm4gkD/q2eKMxEkt5Ple3PmTh+8EcN
Vryw3x7knJPSTOlt3ECygeR2Ldb3Da4uWd7UxtNFYPWa5HygBdfnnX4B5uDzB7dbm2tvWRw4ZEL4
7qt0sIzaqwlnT+8sKTVvF9YPIeQ7y+kV2wUr0Huoo1/1VfooG+s5TeKDDfOoagthMxJCBd/e6o6O
hxcf6wYxqQv6LK+3tOelUo9pYSx7oJhw5lNoOQUkuETi0F1L9vOEwbFZ3MuAxLlGAzQHIMr6cmN5
EUNM+UktwFsa14m6oDcZbvRT0waG2cvGDAf18eNtmHlWVoikwzJj/amk6iMrIZ4LbXr/rXtKWJgW
6dRexnhrc2boCYjpCKR25sF4TqiJrGk01zWqK36x/Ak9zMNrKS7egEhRiySpjwybjIESza1ynb7B
wlVWHlRG7tt7I6UzEe34mq+2G18Za7wiojOM/eMQre1Ekx+dR6UWrhdKHwCJsFug4/RzYCYoMxxN
EDYeOAUJnnmWeXAVQecmn10eZOQVUZVorOYy91GH6uVFYi1gOoXss+9UCQJ/fy5yssA98zH9OnIj
5u5/8uNojo/YXLazelC5iIiGthU0SlOXVDRNLDjzM9lG1dJer2mzlTVvR8GqNw9wAE9asGOZ7cCS
ZKhpntFf0/agURMf38cqUWYJbScXbUJRiATnMD2DONqg5iqlmC1gsOhB1tgMNJY2qZyWL18txh9l
1BUuVnE5K40dYb83QFw83MWVS+FXLf3U6mMEXrOfZnaF6ZeNXtDtpRaTMHJs/2pAIpiRFAmhudus
HqYz/eEaytked3oYnHPfbFrAGXFbSuvliopbJoFlUcJ72WlpRy4m7ASQY3oeiU6dxCNbTakZrLXV
dTYO5AXiaK3rWmg9J8/n60d5Jyye6eLYyEoFb1ptKnAdbETLSVI4DP0XQifIdUZPa3yN5ekmFILn
obsadEWSYFMyYy2cfL4ZTnTaiY7KpwPFr3Yzu9tGQabDO2CVzzK60d2NcBzIvVHpyG9XZsfZuFwM
UbCf9cXVk/gliLhJPHLd87WSw9SKlCtJD5QiLeAmiEcVitXFnrQLbwty9kTGixGWqgJws7e7uG6e
RAva5AQgUY5WYCUolAVXgC0OHo2dqrNeQ+Av54h6FJlcqIpFPG/74q4FjpKlOd4yFtmr+Pyms55d
RF6498fgyzqA9BYah78B4B9K7V12rv4Pqoa8GbI+U03O+A+T5+LvB/LRGvrISNUpBYMcHsnaKthm
UsWUhHwoTgAWkwgFSQLWHdmrWeK/DxGhs3sgJ/G/dILSrtjNg/A7QhDACN9zJaPwoyTQy5+SAsdF
c8DUOkfKNyQdMcq5QZEj50DJXi2sE45tLignhXr1soWBKxzMUNjlt/TuHkY7qTsTcfUWnMBastpx
mfK1E1rynxxDRLI4f99SOUkU8MwTXWSAsbai/dx3Yq5hskYYkXcUzkrt/ptybq7+bQUeIjgCFHxq
5VZKA/OFUE90lXpX8RR1hIET9jHmUcw23eJkEP38ySGIAFgBRiV6iQtIllyux9C1TLqHAYahH1aU
oyhw2tSvIxtmZz7Dj1HnFb66mL/WCQvixjlTeQ5kGn2NxVqWpwvsQCltwx7CcUi0XrP7aeAudqij
P8NKMC2VC/0mxWLZIzvJPUGvEYd9Uf8H5HOr9+HRE4GGMZW8q41NBId7YdnpuMUcdxmlr8h3PByi
o6PGIhNlGtDdhJVo52gIXjktuiMnGYIO75ghxrj+g0Dc6CvdEO52Re8dvyjIfUpiIbSSJfvhGwJ1
whyhSpTL80qCJP4Zp6djit1vM1NnanwzHgqCv7dL+ArsuK5lAQT7sjSZm7rGySVMpD544lO26IKP
4USjyF0Qlrxu/4FjUuwNCIL2Blt7NXTvktLsmyLkBudOmREnUkRrtOad1VFjmxg/5y5YcydObv5H
CrUctC37LSfN2ONsd3w9o5XOJA29GjfgztL7GEfPzKFjuhKIzriOSDeLdcSKQQikQm7sm0ONhthM
VR9phILDbwUEJD/1GZXBmQTsUmVCKbvRDC7/IeJqL0Y033ol0TcvDPhV4HCW0itCEZXq/iodLJvT
Q1bQFtvSAzCFpXN7vuahMvwIDXuvouNtKmpWrQr4Yfn7ZmPbzkTzMbeX9MnlSVMR+igrsneKodXg
w953h2ItlPnQeCcUK1FUKfL3z2yUwr9PIfS9pnaCItakS67COkiUWFvzCahzRlE2xUrblzWoAzZl
jzMZ+PTHj4ea7clLicWq6xs+Kw3nJAEQ//Ih8+RQM8fivy1doP2fLOmUnxUYO9MgzJHKSQYx/cZR
LZux5aA1FdQhD4zQxJ7WDM8XXlMQK+FUIZ9yp578VLRsTyFFKiWAf0Rh4VP5X7ssD158gnmltDdu
SpTXOS2DqKnJlDhj/W5xVVVYVQI87bgF1S4QbR+a/3+JM8FRBwOx2cqXlF5GRqKOav+8+vDc6IEN
Ewvq3r+WYzZg06gaBF5gYhqaKC7PPRFr+cN2zyzh9Q1hsPxH/BzC8uurNt9oDFYjllwvM+X+E7Ne
F8djeDH1xBhmM6ZK3Aa48qethcP5L7QFLqDcjICHSNgk77Acruc1D4Eu4VSvBRRj0J0OEuhoblP1
8A8xtVlm4IGBq5u6XCAI0g9joChA27qS9+tRCN8GzKguToAc6p1atuX4/Y40JE8r5XunuLZAmVCI
FRQ6t+d9dIJRoPKAhXhm0vg1oef4GoDN5lZ5gHpS4tZvAtt7CiGmiA/C2JB9QFR+kzfq20yXh5FW
syYWBQisbxVnPB66JBxq5uOOWen1H0IRasfYKrZWBvrrFx0RV13Kh/aGr1sad8MLXKhrFfeDerem
MO1iiosCt5B+gxnx2ds3nSIaA0at6rGs5DhjuvFIWWtF/puVzgzxyFddB3OO/Ci92VKbQohtkFoR
+tfpQvT6KsK7kiPHwEnWy6zmF5FBFnH/oRu5NqPhYFNd35pJa4KVbHS9EChoyzaYinIsZelJvD0u
JhM2f41/nO9BpJOuJSsm+kKtVYrkG/imWIBUKiLGjYEgg2qPrcMxOOrPloMaNgAkDqlQ57Q5y7Vq
W3DNvnKccdKsQOGc4qRDld3zf29yLtbY7hPq7XdLXAorjI5mc5Wk0BwrJoFrXchKRzn7O5puDl/2
gyluPdV1BTJvt4xo65Wp6IbJrnErPCa+zubPSbf3ENEgL2KWX0S1L3cx1lcGAH/tamqtnNa4S8Nc
+e/izOmw1l4ClWbq+Hv72MHiyc/6h0pBPttUiJK15L2m3fS3mIHfVwuEGTep1WIUjtql/WVNeJ+M
k7w20Ad4faQo50etiSZznjZ5COwsDPNHt48J0VM9DYag0mCo2kOPNgxrbPdNVoEcoW8qucV+LCtk
BObhzzByNLS3YD4vrOrwTk3SsEyDERXePVvVnRQsZR6B7AHLFdZnDOOrwlsGkoEY0du8Zi2kk3ky
P3gYUogD2TSmcOmpAzQOIvhZfSXDUvbK6rwkxb7YePTT+TS0ELk0b/n1KJu+U5X543hKordi+vG6
kv5iYx4QNAnjfkHHkKSAY0Wu30SacPX/AkJYg6wDTg2qbtzE/+OPVNwj9DF+Ev9c6StlDaFYFJEb
PbDV2EGkh64S3doBMM3U6Y0eK7KILu0I+Lba28resbD6KmYdQ60xRQg5LcUvoVZg4EJ4RMHbYZIB
C/iWXxE8e9tQIFfMWHAu3mpYNo58cgqo9yDeVwj5Xp8b1/WYWg9wh5S8e6ddIHCiS1K8ZFntK+Ag
YKoeVShx8RES/2RBbCP9/T27NCzjYH20E6yiiudA3WWVIteDgCY3vKlMeqwhrkHh5tsGTwM9PSNq
Z69/wFDbVaBZBp+kd5rmDbaGV82A9i7acaFPyjjUhyTp7h5k9iGH7h2REizcY3plLwfm38V87+le
wvvlQOsd/tTqrNkLjAN/e/i2tDzaZbXAy8fK1abSN2p9gH3jDlrdADOysCkygWethUh2Sx19WaAS
tj3chkIbGSDIpuhg4ruRZytsm+jhXks/l6QDOxlZ9W/mHRg5e+wUUVZePIIX67kmpVC98vpb5RbC
KkXJPs/x8XmtAo65XUwt64gNpUd0gLY6SkOXn3o3RNoZTHdpm9Rkx1SwTIoxcNEoGxnbQidbMOQB
vx5+4/r8FcXnCx2/HaFW/8yVfzBOfAi5MxvDB5+LCK3HE3AEl89qgK0I416kt4T5n5ZachPG5+9l
lAHDQI2oUhX/EgRN7j3mLmsHFnIr3XIQQbbsDda9ewBDfq/lmU7ZMqHY2AvtvHLt8/vMpJxNDUSc
4mcNWggzoQeDKb2olnU9K3tHrx5Q6A+oEj+1MEAflPr4tVu2ZRHUUkhOrDQJSSVjaB3abLrOmBnA
5YGNNSQkzuEEOMXZJCTkuqEIRQU74rrKFQG5a8udsAcvLbIm2sRDrVll80vuEZT4uYTSog+UMyc+
dsIMSYWts9oZkhiOfZOwDM66EIjbfv3GItvDkhv4PPx97jcciPipNbqXO+NcZrGLbcdKkf51vlNb
0ageszxhaYd/02G1mBJjRPqX3rWTLbizsZL4W0EVET2YaFPbs5V5jPR7EpCQ78xQyep4VA2ZFZix
zDN+BVSQj6TT1gel72BiNyihCOWk6UbH6bzrpSt3eXMXfLNmpLNoOpwttoLEfXHJcsBCdQ3MxaJ6
AMm7dhKVgldSfzeMztTVlkfPauPOzK3k8EExPAg2ndghRwsYip+PiXYOV9eF9dYJkE2hMzoVQY2r
PSzD/mQ4YUxx8+kVrlU1r0qr4ZR5xTK6lL+bK/VYRrE047GEQ5/3Vn8U/ewMFQuOek30ZaLOgOtV
ORGEbYZBOCDT6SGPytj9Jnd6Fn07NLjFbMjTFpF0G32poBJ7NFKZkEHa4y1Z4jNjSIoumSIdWnu1
LXiNM/0p+uIMPw2UcPy6C0KNb0PkvWOVJ1nQtmLU7Q2AiKNgYYBbjcyawMvSl9DplNTITRTWBt2X
U9a6BBm2bsYbaUoLu3gYAFuitLGF+z04V9Iao51D4V7LYAZSppTVHElHlcXacKIla2onE7lqjbCo
AljJODMsNaY0A2GzgvKGkCTWsfEB4vaSCs7A91cnGKRjlGNORR/7gDju3fntf1RfwLzABftvhYa1
M7XycK+PKiQhCMMOACgSZtlJDrQ8WG388nsT9kj6rhdFzVTfPcJZgGcAOkKHiD3Q2gdfMQxcIlHT
dG29/kNvYI4aqrZmFasJ4a/W655CC3miLtdapjpKjQK5JR6LqrWmFf1zRcc9Y6N/uM1CPGs/f/Yz
xZUsw+VNUWdhFLo5FpSkpmuyV+9vez4NeBIWIVyvb/oAs2pHBqzXZvNfwPWgJMxmudiuXJfOa7RG
akMvbwmCrjVGCFvgjD0hWI2nzCit5Za05IG5GtWzSIvoWoApwHkJdIcizviVzb9sKaqf00qGg4ob
+hA11P+B76rPmLC2KJOMW8ecHAxVIfe2i3n7eM1Uh6GeeHAse+tomuyINYbBV/tKogRw6EKtutxG
uX5DgFYLrnGHoI+AFCJ70xY5wkqm0SDw3dj2mVyzqkvzE7wnco6ZtkoN6kokljUpR4UdKDTJtN4Q
HjHy3oKiQOOthzRVWkVUluqAiJK0gcr+UxVjwvPfNnRdC1Bj+r5YfsGEQHprvHorJHJg0vtR0Dgm
77CxCTPhegQ+yBaA/tWWRFREAhxr/qMVh0v8TRzgSUCnwpNevB1OHHNHssyHCXVtEdnb9MlHNWny
XzaOzw6qoqp3vAWWxtuFlwezb6YjvhLr8YmedoTABRjb8cKNcXH4y7KVQ7MVFc+79WFLr++8DIUf
nK4hqNe77z9Eou1ZJ3KyL5JbRafbasyubpkLGCjM9a68duuk4g1LJFP5BqgdPLdsw2+BXtYqifLI
8JtbBQ5wOvVMmRvY/ESUTJ4jcT4bZII95/Z50TJkx/aP72yy+9hCu5N9hzYWs3npwdEuv6qlX6Vc
usLkPXoewimz9aiWRxdZuG0OFDAAxIk0VybjoF8Vk8+E3IO83JTOEwh8SBRodZOrtxIJWGQADPQb
kh7SS3A99gHSmRsXbhDqRJbJIYtpKyLXmPCNm9KAbBfxQMMT9D21lZfUs/3+lLEgefh0j6Yv1AEw
Her8klF2shrR5COEv6aihgn5owbCuRYhhf0PlTjj+gLZftOM21zqZ6HJeyC3aF9Xr7Umx02H02NJ
duY+1mvLbcmAcv1tArgnGCCqw8otIWgNVUM2uBmozfnZFaSnetwBCaV770MYkTvO6UPyJOD/NUME
rvI+IofKibj2PWMRjqNHt2f/kOjJc6+dsoXmfOWVBaDujJIQfyLW0tdVoIHnSrHXZl5efflTE7tM
kWhk1lDUxLl4gHzHx7+owIg2gbp470Pj16xRC1pfsKxsEF7+Hv575JZ7wtBHv2EQZvMmiRbZ7Hk0
+9fXQ4V0QPuadqibqQ2SF7uWMx3+RUj9I/XW6NKPvw0cdlYGHpKjsZw56nlwwZ1pkJOHfhz80rLm
LZS8Tep9gT/39xDHOlj8p0bAer6bdgJHG6KI5kJJfKChFWlyO3gTyg3oJmC/xBV4SYTGv1rP7Wk2
Jdmqxk+hE5sVEiXq6Pyce8FGfNFVPfc2lKBKH4JYYFWTqIOQ/6LMyabr6eqK0+Vkjf19WvZUNgq2
ywzL5DG7agn7MyRVkY4d1qqbI/It/aWNAknTt+uWxsB/c6KOnqCer7H8Vl37ryFwd8gxARdiZPxi
YZR032VOn+kdwi+8dCTUEHBQ6CpEhHP4UxGzUSpyg6hZ1BjaM+ABIOl70IhcwQ/Sh6lyXZQDZlF6
KkdMizgYDqZe/TkN57xGdMCyeDewIOHhjvct3tIVjgKipCCXycPvgNhX1XEfz68KcEFuEQr1sExy
8c/lXMKNZtwqQdkaMdqciYo3QjK3azGsM5xBHoQ+F8ANkeiM7dfH634IPvlydNRsCzPklEuWAkYu
cfjLJlPsoQuDDtF3Ww0PBfsGRRMy6j1S9LvUzQRxuuPr5rbMIY3CdGF3eJV1PNCQy1ldxf1WA5hz
xd9hcevuo5xY5tWdyrFv3MZQ5zNpViAC5vl2WFZb/jgZLF0Qg7Add9/++4ZRt1kznkxKU1uTc1nE
l/lXT70J7jiKJf4YYrteLazpRRlfn1SNSdeHmBE5srXNyi3gLg4BDCwFrFTRYuG0Dh3OfZ/VF7w3
wHgLhOw3Pd1+ZgOe8VnZexm1krRc0E7VaKx17Ctt0twuYHZN/rE/KEeeGO3qmmRHIfrKBy9r0R0/
se0wb9K3kaxSlbGQJkWmtzTX6ur8BPoETv6CZUfuL1SwpxvYDhTAlqbnDGsuZhgm+C4dLVTyI39A
ooiljHprhFtO4az7eVgu7MOvhvW3g3OpLy0+dJNd3Pf1fdRN9obQ2hIUrsPQ8DDDLQWkdBCNX4AX
12ThB4Ooi5xFqnp7mrDhZx1T2+IsVfmloLrFooqz0NHAgHMM/6ocoJ30QgF4QfLDFF0+vjZhk2Xa
a4ZvSqdCcYqda07rUXcBXAVtqBfv2MrW6EfMPXpbh1ZH+IPlSv9n3meq9SOXE6pgS+aT9FRpK9c8
9s7Vtgh6F0GLi65iiu6EyYWnsrPexN0nATO5kjpKjP5SrvSdftBS/MUL3Zf5PmVBWiJ113s9pHG9
jPvVptBjuOMAXIaaGsRcz/TdoX1RHCFO+QfQOKOwf71+WqwCVpiXjVhK3lmWkbBZr3f+VStF9D2g
vOF34hU+jc6DADEu91vRXYxdUTPAM3HQkWDB5+WQOeuLbsxowJX3GIR6qBj6FOKr/NnYicbwBamY
cb46REZZmlDygrJRNqaMCezJ9vH1uKqD3jziarHxoHukFMfUbrt5sg7UHDROU5DIdJp61p/9dnbZ
Wr9OTK6EtRO6T+tbwapiQNZtwGI9ivsfbwSef3kyUrDMBAsbzdFu4p9HMa0k9eOSSSyT1xYfzp0+
ZYa/1iuDbXIIYAasEYCx+P9Q+jv+PzNLWpA/SDewcfrW0178MwxX0jp6mx+3L+C+Ah9BhrK8OAWp
3vG+/gyUhm1FhDZcjm7wWoonmO2fnfu9hF+b522EF/N8zGQstiIOxCgWPee5zWnPeO24CTImwpwb
JCGio0IJ19zhFe+2GdnZALYMGPeYgQETGorZWbCYR0++fbLqZVoWwzWzGGNOcUXFtM58KuSpRsv9
wsTNlkqNB6Pv37gAoTNb58YeWtqbRT8TtknMBVC3qaIsUzuyehBDu9hN18TgPGdz+HvX4Uh+LqXp
oIh4bRW0EbrI80wcjWXj41gkyrY2FjDQ2tXdC6cuVOWtKgt7IVVzIzAy3MvaH2MY02rIQb9/Iffa
qN3c1xBU3hLXirlg21GSWoHqPc+ZGHpj+VxNn21TQOMb5i/HnkM6t/jIMtw2MMQYQkuR70KDm+ps
sxJlSnMdMKjV4aSP8FXbmV3ZyqO8XZ5wq4BSGalyqSR5eOjCz/CjSO5Tj+hngCYO3E5YSTL1UnBo
8KTUh6bgwGPkJMSmtnHyBivb6L+jsS61yt4y5DdmA1XX+44NL9nPUlAsbNknurjs2XwSWWiF8k14
SetbBWxNDdSZU0qqXLs+jL4U+UdOPf9w6Fh1Da5OJBpTs++3yiTa1Ib2Co4h0CLAhiOlB1Edpwwy
l+hSJFz3Qza3B0W2xHFIAsMwrOy8ct4mPtXrAac/HDRPWqCgDhppUZ/61fQxG+YQXClO6r0kxzbP
pw34ZL3BppQWdEpbdIDua7pUm1+y7nSPcc7Rqje5FRwHcyb9d3UP5uMGQpclhZ2YpcEZx4U1xKjP
Ng8ayeUhYGRGi4ChFrcdqXH07ixGqA8KL0dzWhkCgb2FtX5J15tomwqARTajs3ahLKAuOlDb40MQ
GnkyIVHQFCZ72bAeOP4CGUsz3LVUmdisw+ruBPgb0tn6iGcMqceA3+9/rX544kpPVPsoBIxkPato
B9kDP1w8Uc/wSaGFDJNX46b1ogiqGFaGc157gAUiSq6mAd3hc5fCPHd4yrDetAMuZRxIC7MPlM1p
FR0Ks+0s79p65Vw9pwRtBgCkjXdkecflc9kJ0Ff8nDZ2QP/LQbo/0ytmsU1CTEZLxqHzwYGnLQ3a
dAdcaQtGj6L941o+aiFeqxT8mPwKSFMxX3DjPrBNn/7/tjg2F6gNZ+c5ZTdW+r/6hr8RQ1e5Qh+A
ZeZ0ek9Lw3OkgnWIU+MEa6d5oVeEDjYNuOhoiC/zsSibpPkM5deb3/gNQISBOJJkKI+8/o6UYDu/
UpXQc48JeWirphD2SCZsk+re5rH6S3s6lKR0uGZyIgrwlzNVULKCHCOFtsvR0lwAjcF88B+uyh9W
vv6nEVp97DFCjWUM7tEcfIWjKJ9PeJIh+4yiELWFshy5vvKQk75Ld2dAlIX3uxlsboqmI8iVExnh
yKbG9SQ7pN3u3000bAHk09nwqpUIejr1glFsJoFNEqIhjqdmDMSELJv9SL3FI1ksMqZJKH+KWd5M
Lrexl6Yd4QvqE68wsYVk03AyGEltyM0TddZif9EUcHruYx9pdz59lZzM9Xb2SQPsvP2rsmyhEIVQ
LKiDCQhQjjWkSI6ohF1ZbrEijkD4sb1aN6Rjp4okabEzpSuujGuak3CGlN102e7w0USC9ArhNTsY
opQFhFivKCUsRUJy5AwRvVffg1qrlzJxh3Lknb9DbC47D/keTWrfp1X3oHEyjY9Zso/QkxRP1IWT
fqDyG/VnsSB2awJ+AO8k9G9UWwHwDvAycc0/c2q/owfk6z2PMKc8NVNHfQ6RK8FOuZIsXrC/vdRj
iW8NAzP6G4XF51J/eT99SaagP1SzpXZBOMkhSEHDClqT+AoIuLEclr33stSLeKKaXNZ/bKSZ2MmV
Do4BpxL47wwC8aP6c4PPz7XqAyLsT42UxlAqxLSJZeJF96ydcFQT398KI9igcBucJq2jQXQv/9Lr
ocna3wWp2m2VgdTWMWX28w8dtOV0/qMWYXvo6wWx77egDOI6xLNy+yvcsOt/MKzz8HjvZckVL3J0
q/dUHBM/8ovUjvAeuyMqsL0PBR0oQDPsxMaRBwzypcx9On4K6ckdmuFIHtJZzmxtBbPtTHJ4i+G2
EW7Dxx4PYiP+ubZ2/rArAkqrDYUKSFBmazLpmhzIXERJIiRUbf/QY4eT0n18laJQiPd2nrQndGwf
ok6OGfvvZIyfMk1kOiJhKFdL/V1dW7R6iHtHD+jH5zUdHOh4NCocevumN/p8ha0La4PR57jLYi20
uFO3H9TP8hzsFo5MYqK6WgFszy1aPwK6GrWekYej8qMlNH2Wqp1N6DwDpDS7Y2ms5rrYEdagGa7M
FK5GKlWyIojTeeAv3P3J9KXtbwFIBFN9PK9CG+GL3FS7f3O+u7v2zINde4s55zB41ZC9aO/5BzdP
lueGllJhNxUaSKUrEwMtL11XVh81XNZTl5VbPqsrefMn6BwAARSvYHs0d97MKEtJLdlwZZ+jmWLK
H6/vlz7/4mIKVkVSGhpC/0BymTP2qLfPdrcIsahxSQ9LVzYei32VHpv6a0WXrx5SWen64ynjRVuS
b/4DQzpgceshW+Cn8cE8cmX7NoVYNz62cw0L986OSlbewViE7SnYcJlqAnxeRdSC0FNeMph2rZEU
gLDBRRDpS3pWgsshVjsFDvOV8/dCEkHSETOaZ3U/njciIztPWMNPfjb1/uAOlqOK+8bMaSk+dIdi
GA8bSxcAT+CjeL3S+rzmYmssZ1J6DUuFPUskmnVixwaCYmtt73b3CVMG/s50Cmm6VHH2QMl34Bi+
zFML708/kWIrlpXCJ9XdSbW4cBFSBuz3Oiq2F2eQ+aJ0ajKYYHNvIH8nO+J6IvFz+azSCu351aX7
CtHhp5MKKO6AVBU/drsVRtPjtY4smiHOviZddCSnkkmJ3JgaLolKlImkduwvo1NZ4LuzEiKwxu7S
U5w05N0alELgCqR7Acv7k0tKFtM61Xt6DJFhZbYKMzl75mMYxhvaHPKO4CXIvcH1SiTOrJvVHDy4
XgOy122vkIdQbWM79uOYR9z2XPcTXsCvD6a8eznTyvXGGaBKppkRS3US22pvy/tHw5BhQWJraMWD
e3E287h8KBiXug435gFeQMOzIF5zYtLKJrAInDNuvJ/y0U3bbgOJ1C3a+bSjiTnq5y3jyapPOlyj
Pmhz2ApcnP1DrEzBcgh+POmli0QM6IToU2p1xF0H6Uo4/XFqSj72YFdycq1cxBbZ1AbTvZhhSbun
pSe1jWM+N0+UNaTu1SZBgD0bEtL2EPudA+NrT6gXrC3NPtJSB5I/G+TVZbBxBwvNpfyeFhA+uJKQ
DfBYlezIrbwSpQ84x+QiaC8U1gGM6zYUeZchz7YXBANEdOyXwq9qEM/0x0EAC1enkInUeQohVlxp
BbHACRKaM+zGkpOMiAND+1MmoI0I3lzD/kC3fV01157BQ3rUIM5kxTOcfXoCf9IFypgDe0lArqIW
RPAXbx6c69aw/7JHc9dX7NYlzxx/y03rQUn0osJ4DvGDFfYlmU7azPOaZ5WPwx0x3qNp4nhMSFID
5LoU4oKYyn6Af9rYQtza3lH81Xr08IpwTjzID2r/W2Ync8o2SBQ1Tq5FVDBa+xeOf0jkkZblOMzQ
TtZjqwHJZiQ2eZqTIjtO5B4sh1avOa/NkDhB8isdlud+J2D2R2lcCM2V/bopFQZlsjxt7Khsl1Ob
U+i2SIKfF4dkQKf0AGwe5n5FlJgGZsDT/+Ecu+vDS7gJtbS40pwDn0KfMawLjpNWZs/XYU4IZQTc
UjIhmMWcJFZMj48R0+4lmbg6Jy2NJPb2+Udxsd2OdrHtfz+lPUSTZif3T1n2dLSa3vMEXrkm9/He
SBJTBiIid+7a80giYjPSmowvxpL7zwNHtKcHzXuNPS8i6VSiEgyR6GkrmuxA5VBEkYgWhiZWf3NT
og/gpKLdDo6+cGkxMlnbU282YKRN33eXE3Kz4uwqW8WYHbkfpFZruoj56+jT8uhVLOwJAYMIEqqQ
Vj7tOXhIq9pu4cSyusn6nhkXJhbuX5uJWlbQ6v+S6IJssJIQuBO7Mrhbu+WkWlVPJcM6rshxdssN
12f+OawMGCkUfKaJt0X9vQ6PMl+4h0rvpxeNejWn4dxoU6GhgURVAn3ApA9hN88neK9dDWZFo/nB
h0z9WXb3lvclrfpXQ2XwP0AWpGS36BgqXErwEwpBoqBKawNf9Ij4PfQQF9H+wPYQyK3kYmK8uQQG
/6dVlvGtKOUTsFHpruiozhnacJrcUls0xOxOeL69LXDK3QBXhaRE1TsThLwIpuEM5ALTEj+jXrg6
5Il9SAFf8sSd35JqWI9+TacQXFFuD/dTyVax+UR6ZtLg8Cs9IzHGs9Axc4pqk/gMoY0isWpmPXLw
wP2lB3jWb8lREE5tYOwDjwEs5uJ2ybyqvxnom0AitALLxObPCC9zqM+GueKZoRsLSX/Oe9oEk3AT
mt8Lqh7/fvBrMxwO8zO13Vot8xsAB43G+ZQpT0X9hqI/se8O7lDjmv4GWWO41oiLwItkTW7CEJPp
XvBOdc0mzxC8MwwNOllYILMDjP3faHuMP15SEPECRSkWGL1hZ3KEG8f7lZVuyDFzYNMmaf31FZb7
E+Ki6N3V1M/YlxqD30l8z31nVFsz0Si3vwfS3tD7u4WHmJjbotudvWwmg0Ea2YTordJOYZtN7muT
8XRwo0AL+5ZQYQ2IvMnGm95iD4AIuVKo0Xw5sd2J2EzcGfcaj3nErIzAYQwkpGJ/Lk4mwgSTqHDS
9ouyJ9FFh3nnJRLI/aeBpWldNwD2kICYNahV4Ho7n1pd5rTANQk51A9flTaH8+blBzAaIw99BbwW
TmSacsYTwyO0qnTmH3+fzlHljgqrAAUxj6j6QkozCxM/78rkLWa93Yai+GLhZpojJVYaU2HKHvgp
wWr+5ZSUk5k7CSmCD0wvIay9SreAqrOGEHV+xNjA0+xhFufCrb8/U5s6H6KYL9gwZPooMrtDIXvx
dmxA8JDUV/80Vl0XMaFChTLEnyAVdB80guMSGZEPMkOUl4YRrZX3P3ngKFesX1mnJpoYn6ySa069
l5HHymLZ4xef2N2WrNxQ+37bsO8FQhKJPDIHVSSiqFTMoC8G8RbrRuQasD6GTVXl97yLg84p0yHp
OqC5qV3i+zV7OJrQXazt4YuEntLnOK/gHeQJV5VHs/bmLYB3Y8v6F7D75cQr18ZYOGemaenQ8+O1
ioiCHBcVH51WMOAKpaY0hetu2EnldMDUqKXrS+5hu8WLsNXIgRiBHAiLiTUljWlgYN1Yn6f6Dk9Q
DaJdXjMpVQqYtCisVuRoR5Dk1n9oghNN8sBg9d/LcyeqS6J/w/XWJo8l74O8rGkiaXrZczMTv9gz
gxTgpRN0hTbnWc0EErd3nknNRtQL41tGPE3sl94FMsdL5qjpMRRyYh2PX7PKRuLdxXkh3Gsn/DMZ
Dlc0Kp+5wRxZmKKjTEFb5IYBsAOdGFIcLtLOBjtU2AZOrNP4xDZbjn7GWTcqWYkZwUd2Y10bnCxu
+nM7CjNsqlylwExnOtLe5onPVKxhMExFe185Rnk1LpdlvOUPf0ZiIs3f47fzl0mxHUT1ZmpNJW7C
/ppTIz0DNY+qN5S4Xtd/J1hgSRzlbcvjZZ14gtyfEJWK4FUrw/rFxgduDSfn2Yr4sm+JCxx+PuFn
DvqCbF2lvbq0jcoiJ0xMU5RmisKetLxbUg/vLuW5WQhilfLtJAYAettwNNkwFzcATG8HOWOgzP4Y
klA7WxDDlv3e3CBuiOKa6b5f5uB7RobcfDwUUCDE3AHQKkpjmoFzw69y8pO+71cLUQtZAITcXo99
HMe36YmGl0m/E69EIkkJnQcUAavAywbm9tDSFkjzocJQexH6mk24iHlzj0muOHFxCqcnr1Ayi9M2
sW/9SxZcL8YGbZ1H278LXz/0gfjlBkbW4Xzr+bE7ptRwBRxnmXPrvaU71cRn+k2ztntWBUmkeCZl
D1fjoewZfCR/KjE22FTfknFmezYp0l1TGBsSId4T81rqKkEd0QW/QaFyQ6vnGPSoFk4mDQg/q/sY
KH0vImP61WMzgCHPJpBUMM43HU2AaOt8hvhs6QYRPwp8Hb0HH1m6t9sBb7BZJD6OquVQss8T1IGp
FnKHlPCDFiVyo4w+10eeKlpILvPU+za3BCYQWZsgx1P14X//PgmDo6AKtHFkte7fkfIJ5IrHmGzr
mM1yO+O/qBdQ9mU5w3SnS1kKRz86pkE+7gljtbwhvFVJvrhj5oDxvMiZlXgRyjLihSjb3UByg0Uu
Zk0EvVSmCuHtxXqwwGy2V6G0Ckn3ei9dh+BzSUXgz1tgSWy3j08Ti5T16NZrh5CNQBYsu+yB4zsp
KWl/Ub3PswO2LxVkaFFe9omccFOXg9DVmYWPiTnE6cPbip1rH0b/VhE2S0MnQAh0+4fCmm0R9soV
oI2IbsEvjyOqoTK0aJKsn0tLjnABzy+zlhDC3rA/BnrZqKYnOi99xv80Sl+THzTG0O/WObuKu3PC
tEWQ0zEe9XMeJGfFrVFsrE+HTV/ia4jE6L4C8P4L4gwMH7gRMsLtciI6ye3ajfL6uc6yOeuGUpEX
fc7Mo3zgCzptTxtjAzSaAvuevGRiulNU6RiVM7b/A4W2noFtXEIfANfhhi4sZR5p9M8zBeQ5325q
oQaTBAjmc/of5qVj1MEr2rDuy4WGkPgLepfMutMgMZgtwNuPZ+L1H7qv7+8pS08HYkofJ7topUPD
zO2aoL6V1gAwZNzkXvlLz43L401Uc0KdXKNPfUV0/AiYqKzZlSYQ0Xq+a9WEWPy2Rm3w4ZKlFzEX
WtpqEtXA62Z6KPCtAvBolEV/XBYYLTE6J0zsQbMKAOrDzjfNQNBn20ycGC66eKy4d5fNvq/r4nmO
a7o5xQmwEKAb+QNY+Dkg9bQd+TUNKrDByTLVfI55a6Y7LDqfYjrc1OZ0UQFuGTxNXoKSLCOb4SRd
CTPW+DAafaHJTfc/OFapXOw491njkRYZxXBp0gojIdjcf1ZDKEyhJ4Pcei72JUYIaSnD3kfkDCkY
R4pOW2ZSYhe2nnAwD6HwbM0F/hVD6udpTljWoVTIl+ThTfK9yA2puJR0Pi+Rlo3wPwLySJqs3UWJ
9Wzmw6sRXRHw7xhk1Yyjot9tosKue1/ZltU7KXlYQ33JjJ1yhRemT4BlQSfQH23qIJkGRrYwbBM2
AOMf6qXxHXQd4AsDU9fSKnasQMvujgU6BRGTSR5fKrLBg9D8NLZ+Lv+fOFm+HpQxJPyyb7Dmxr7f
4enkxjtn2jC7jxn18uBoHhu+PUDKlz6Q32nLmxcX75xcRbLrltNjUQbgceFrGxUHIYMqn4mmlmxh
+3pnWudxB9cQHicHxLSbIQRt+kuDje8JiObj3MkjAmk+jvwkwviP0Xum01qZk9CfLEOgaSPNVd3n
1rYjlo9WaT4N7hYXTnwlyboSDb8OrQ1ixD8Auvr2GOOr+CZKwfAx0+tf5AonHiNHgCbkCpO3hVYO
RgeRN5dsc6SkpVKGCHK7d1ktogIuGDbdDQ6kndYNCXMdZBXdQSO3izJuDbvIVLg6t1Y7zaNLrY9o
R1hToTjby9z1dkmxqkabFEXsf7s2ds0MJTbedaiswqeSF67yJaaBQKfnmeDRNU+1KEm5/dM/30kn
f/aWlwZcl8C1f5zAr3lOf8zwvl+drW4WJb9azphCph0SOeTZOkEQbg3BPfl4Nb6SpkNMIcwQQXyD
DBsAt6XpiKJAa3YsUC49hkan9mHUW050MLgSiYPTjsPxMX8Mqu12vlZRKtuPCXbDXHAb8qhxK5tD
uDkbC4YBFn5SaqT2z3WSRXUDkC7s7aq6fcTqSMrw/KdXX0jVm4xWWt0iVvplFtTAK6UubmIhD4bV
KE2MwVrejjW/HakwG9Dck3N223VJ/p9oh3/LnrgeUuhB0dj9pWj7gdXmWzdhOZ7lBCCgSWIPs794
47Bg95e6LbEg2y8eqzY9gI4GzsYpXz4agRO7+a57pB8jeQKbavChv4I4c7XuBzYJh0g+yTKXCjit
rkNTbiskcgl04oWGoqjnAQckUzLg3AHtXUT1iiecAYXbIf6RvYEZWVFzY/Dxo1KWmtTYEn01qEQu
rYmYi5GNYLyccwoGgxeQ5aSPP4CYR7i+6kqZL3IiUe+qFCui8qzTgrdXFHneAAvzJ6k1DO19loO7
ZkUtCppckeco5XdS0KL92JpBcmO6sGm3YNpXJPiibGA+7mc775CVGn6cEr5lzXetet8FxRG7jwrx
wBsFI5KXyuI3Iw2Gs+IofSOCZKUOFApUaL0srb6kp+6yG5KMAkTqr5ByX7zTPuuXt3sXh+yW+RrG
WC+4uqLW/SskevqJZQce4X8zZO1Rj5cWKyxPsfQiBw5jdyPEkrf5tpvS9b1U3n8WIoLK1D2GaM4/
D04j2MCw4mRdBVAIAZpvZMOCaQBFkZHUvROoqpceqJDuna9nvvqQTO1Uq4Fd+i/H8GMc4WoHAa/A
4rb4ywws2h2eX8M4bbZrY5HE4UgL2Ugh1gv7mgc0MRKKcF0GdRwtJjefnLHJIp2Zi7TCJf99ZiAI
2o2n4qkLE3XDSK9E0CWaMnUbjY26ltXpUsi54GSdEShqUD76JqBrK4ogZhsITVXbujPjpZEgP6EP
dITuxLHK7njXYWztHhTCpvnA4wgA7pJHw8PGKrwzY7zHOX2KkXgWDqg4prvzsT/s//DgcNhA006x
vD2y8jXbaqveACAJxQ6QbbMPftyHtQfW9xpP+0Tkmb1X1pw5ubprkU/fneD7tHN2Sbyr2ih64Xo1
fC6Sc2o6mbzM1LnpjuxCwOvSJN1HncANLcM1Rr9c2nCswBfxhi3H/nJevTOvytxLx6eTr8BwDwby
cuT++406zxyBq7auYNafbH/pkOSHVamor/LVz4OxpXeaNGPlDOWVA2DawbBy/ieFvbTHgUQD+PYQ
F133NtvL3Y3XAeHdDbZw/zdp1rfe6EMq+Hc6NHaqTD8ubtyViIYrCGI2HJurw7r1AJEcG34KyUME
ch7AqKJJ4eez87G76MhBZzgB472FgDdN6sQR/HednpFydJyo6nf0nEUATO1NUqj+s+soyS9e0O+7
ZhQWE4KWJ8PaQjxkfSB2v/UaCvOYvcfe9tSHk99nhRlEOwikf4iYQQl/lTWXR7smxaCP4RrGDbHu
WgpF9JgIrAZgVy23OdJ0OKL44qECiJ2YOIik+3EqwnMpdEJRcL16OJNjU7bGnm2r6EyA5kMX0u+O
aLaIsqiLrOnnFbIPyJKoENw9zearjLT5FQsLrT7EY44uHlBVoMuH2Iw+zpiX3gujpdhP2W+fUTIG
M8i2zncN0d9JefZsOVzyubUO+F3ZAvUXt3CrQ+IXO9ty4vRQILNNBU2HoylSJsgiKSvqwq4keZK1
O5gQua8lWWX4472O3mekZeE4XJXOhGW7fLmMCvdnbFNbPacb6G8OAECre/Gpzw2khG9moe2AbzXR
8h9stuxcloVmZeoA8acriYyFhzpd3JJXjkMIJ+/H8dm4rY8s51sKd8q9kAu3E0a05e7Q2V/VbbGX
cSHZeLgOVucnwELqiAtMcNDqNRpDSND00gA1168K3ZeuNQdMkzM4JcpFLDjSlgZexU1AYDSvGRCY
zBLutISrrsjSTka85t4BwfUC3B0tdTQd4XSOYxEXAJlAsHYBmh0ZJhJb/52FXY3lNf0upNGoLTpQ
Ehmim1OGnK3kvsXZ79FkGGCHeklftd+h6YhsTYL9xSQUBlth2LqOO1YOjGId+Fhu3uBE8MqvZccx
xGuoy6r1GGH+ghZJoJi00tOnqQYiADmNHMfxDc1Zvd31DvYCBI2Lk8vcWcyLfZDSx1NMTpmaMtqK
0m71EW+qSZtYC6gCHOq0oE0npzDYuo18YYuqDhjFvgY020O4jZ/szaUF9/QfJroCCvWio1SAecI2
5gS4BIfpQ0DZsgEVvrDUzV8iXYE4pZxwd9AULqsYmU27yKjsoRAZTUQrw6Jywznq7B5EKspkKjXc
c9I7Df1GX89eIsJKgX+akuqgzOhXec9FEU3NxQSh3MiFiaYYvz1v6dG58hFwakT+/sXwQqDLTzTV
WzEB8KeaBBdAk0OTzxhYNIEhLESrbKowp1YRcF6B2NmA/RIMqRuiQ4W20ihEhchnxtMQo28KTudH
l7kG9phZ3uNBfVidkMEEHae9bMk8pHYzMjAXpUnhX+vw07v5bdwhJkzl6VefGzgbfmk7uyuuR222
A0qsa3ZZV9VT6jz0D/8QnlfuY93li1A70eC82YTMEsItoPqoGRgXu/gICZMhCavTqFZczlYZNnp+
TxG12QD7ODsMyhCbX3IMopu/7sR3DGRq0pYYTr/vujFAu8MpN2VRMB4ybCzU19oMd4xSD1U8z25X
oz208k2BxAYQSHA91hZmN1Ta1h3tLO5nDr4kSvCe27aMrmlVT6Y6yIyxtRtykPPJSPKqbo/fPS7t
j4gtf/YPjM6BkuvCB0tYXiuuIAveDAvaB+ur9jOx2HhDjLbJ3PhvSkB+syjGVRqY7lennRaSuwkw
1UHkduOhzwtw7F4h7KqAqq/Z0VtLWDBYzqv9bF+vd66cNj/TPlRkbVGIb+YNmrGGCZJ8gULARn8k
BMN9WY20zt3op9rc0xQXYyRZ34MRzCF9bo9h/8tVBtQ+cuIJyV5zuiSerbFuDbd8jWekzrTInGuN
/PddutW7bWcbmD0auIPoTW0mW/ja8UzhwsUTMKnxzOcUgERXNQp33hHpHS1wNSs6OWgkLBX9RRtO
nEdTHkbMGHh59Sx9gEm5Jf589++as/P7RiktcmIYPsBgBAPCQuOTeu7JMBqvmE+qAIUKZlZvM+7g
Q3gUafyOk5QsIg8h9FOAHiGF0l0Z6L59mX15Y5tLBOt64+gycq37i4oULsHdMOi0GMXrQnmYRxjb
j/N5XP57HiCnd4BgsOqU4gUQQsF/o7EZL8G0P17Ee/Si0Z5I4Inu2+NFr0pnJU15KT5I/1pIqF+p
IXV1plEyl4Heg+LHzJU6NMJT08B1psFtC7V2nBmlYr/2Y+Uhqy7YGAuY6deqd5VOa/8lzw0kIc2C
yG9E/VVqP+zRzd+X8cbXTkqEuegACovRngdq1Xm63/oXjXlPBujkIlxBvRIW9H+eC9mq9IOawHNe
GMHYugWQxKCCw3zttXVFY61lJ6pO88nFHIn1tk1UgZ1iCJ1NBZcZ3sATfaVecq/gGt2ckpQskPBt
xyK/FzLNNs21HzgWk9VDCZoYtHfQuW4qCZ/Vdkj0opzWBvb57objBotg7RbKWE+4U9ODMGXBWYpY
PCmguXO9P7k/b3bMrzsfl+mbiLpkfTwq1yfLNsUewwdZjYELD8LwYpTd3WuIlk5RyDDIzsFhopEv
3lo6tiNWiZUwDQlSuWcq5I5dYBOqbkT07lS9BP45CYoAqtubTXeg99znUB3BzrI3fQwK/O9/USUL
f010ubkxW2xjWPXHNglpKgVsdqb0aP8nZIWmcEHE/VfMcCGcbZ6Pq0jzOKjr51wxUc+HS6TN/3Y/
aS1OIKDrMdz8GPFV75bUkyZmKqkCumc8ghKYRlk3dMcizjMeTl1h81tTDjd7I1eviK6seUpYvyD5
s0IpPu3nNCRvMvAc0Avq7l5U6unSXnL41jbFubIL4zeufGFRy6SPFPer63NauMhivkVU4z+zUf7E
TJ2d+Na0+eSWQlRRzIUeHilHQbNcxW1V/JXrsIM6JpPBnZMfv/eJQ4HwxQHcBEDHbk3CiEpkAu5+
W7EqBSDSCa0Xg0FxK5IMXmL+E+cM6k8XK+VdHagt5WFCB8dOEj8yquxpZduTrfT0OO4tNzgYVGeL
LUCi4F2NKEdlJ6Q6I21cVPnqikUOs2tLO7ZlkuzFg2dqyE3C5XiQWJ7kjcHeNLWXJPv9tDaqjLwf
7GM//AqvsQZKu8xnGnhgMB98miQh36teXYVXUjz/sF1/hiuvKvxpyKscW5wjclnqVal7vR3YKthW
iwNhmTQ1tqGcFbdPvWskDg95jxQW8DhnH1JSz6y9nNUAw9J5LGYF2ItwcJBuRMDW5rh+ljubtV37
OjdZwUQGKUgs2bsqB3VAhpnsVh3C4zj+5hfA6uPzkRoUw0Zi4hlqaEjTmdNoKi08Pulbf0VDE8yq
zk2MuIaxxqidEemeh3xl2XGTQzxTG9PJrZP6P8UmUZ7PLqoBapccgFpOpG5P9+PAdxlJmfscx8vK
NRCHk8PGwSv8dW7Xth8F8DmBGRVpdy3nXMErmGnNptNoBbsjdFpCUAp9783TVH/leLPSPP+y8Zcp
UgFITWbLBQQlKx7fS6PFXRtbUJhB9J9RhlKJ9Chs92yYigUlPY4c56JEqknsv28lIbaXHDOHDHoc
ELe6q4o8yR0b895zj8YXkNXpP3Yttc1BFcl76RCse3xT040zUQLTmpW1XNF1ahdUlG6CazecqQJr
2xPzW7qL/7UIeMUq42gRx7FU+onrGMv/sZiBzaN35l8yOE7ksyt62Kiwm7wR3z/9/LGnJYBtbDa+
VRHt0lndGM8Hq96FfFq74ZhzCEQdQRuY3rlRxV5hVVx5tOxTNRzWkQXK3zP/gl93Do5zwtC4//hF
nYhdirAF/q09dizne4s/iD9hsTihU4prT0SBssZIsPKX0xu8W/grPxNJmy0/q/sbQEuABqr3lpUp
Zft1FF9kd1hY4DP2tSKVzwN7AMS/CIsoKKplPGG4J9bYwD3txlKWSwDrbYuVExl6eUcOhjnsrOex
jhLKox0DoT9YxbHe1IrBMjgd2H7qc62AundxI59Y8oidMlT833obWHEzq+tT9lFh5fyeyIVtAHHT
KB/AycdV9hj36kFsVXgvxjBeGAYgK3p/suXX03VUO+xBwIgbeTCFUiMqXlBzqQHD9qwALqfJtBC6
2jto7xSe50Qy/j/f2YZpdA8uRjS+pcMDam26R8C+R+HKgFEDD6KLeaRTY6bhSRxtx0twO/T+OfRC
wq/KiAtX3dQp5eIN8CQxLIPVIzykdzbOho7hZ2HICw4tsd0Q/InyxBg25+VxxizHMOSwNr3W/gaE
INAvyTIZr6qNAPpvBX++0rF4raR6efZV79ltADOtLZH1Ya8dkG7ZTupSI/j5OfJ2yoFe8H1FFjPT
xKxRoURaG69zrOJPJis9h33exJqrI+DYcuJOnCUBTYEPkdd9DWGY+VIkXtQqhP1yrp0r0roRpq7I
SnJKScMhsSDKPSygBEJPwxqcBuxzQvcIbEDfKEWebjszr3h2j3+RJ/FOPxrdcQ+T6/7UEsk/L/iK
Yvzw9oC25OTQ93PRbWeaimFhpZeOBzRlwvQJDrlB7RSHRbusvlkMtQmDzzcyaYFHqg0yI2muT8tG
+cdSR/ymv13L+bukEM01os09Q85nWWTf4mW3GXzzK1MBeohdy/YvuSLR/QeYoQ5++NDmqhuO5smz
SJ0oyidUcmHQg8X16tPRdm5AftVdL6rQtS/Pjzbl8aYkTRimaoUApbn06RlR4Le1QNai0Ruty6yO
E56Xo525sZjGBeKnICHHHfutBnasr2ro+F5Ixsc7fh5g20H6jhEafF361SutviHTzUW3zQInJiPU
6UDyzrB1OLTiPLkPws9DheRAkSMg3hcu2uvvZXbugUeFEEiJ9LbdO9gZqWIdsq+u8w3lhdXw6GHP
4vB8pL/vdJV+EWcenyt7cI4TkYUArraDtuFvgECkkN9Z3+/ooSe/yZP3snvYjnZ+faKHsJi5Ao5g
f7MXssHQODeGtvRh16snHlVLY2w5jGS+0dhotsid3//rYJA71GlTFOw3C8ldE/pycf5IUV7oarxc
i1grcnk/X4n38+5xdelV0w5s0bG/XwvksTZ8FaRuZnoaBKFm+Cyd/Uypk8FpnJRhfVIDQ3e7bMB/
pZXGPYMbzStg6hvSV19CMYf+pQbHmeSY/O5aZHI6t+xKTWLLXG594ba8Xh3ziUqbkwlbdsfIrbD0
L9rBiyRrDWKwiEYnmpyjM1VuLhO4mPUsdxIpBNh4U/tWNPDRrVdnQvU30bGLIQPOS6L6Ng26sEEY
04ZL1VPFh3AuizM+KK8Lp+Rarw8F4gvfxQUttJpVwPs8zODCDsMq6gJSEWpV4pj7Pw3V8KSe6QGA
gC8n4UhaCXCd9LD3XoTeEy21CvJqQykVHgcxOXd0EEy+FvRU7+XgH3K91ClPDorThHMqp+IRkx37
QdjQleDLNy9u87wWHDf6jHogFV5Z6pM424LD6lZFs6lwtQwQXyd9tsPxTtnlDVE1e8Sk+bqVibKX
pnneoF+KAYGqPZOplMhmccfnXdW4DLdqK6ArWkv+y73GXUUabnDUU6dwLdsIcA+p3bliGuIlLFmJ
DJXSyICIiUAXni1o3Iau5/LwxNKKocMSaM3Esm0/mW1eazAcsmuQTvIwIh7VWTgS5UUL+OB9cVLn
ms+yNQ0Ur3UBUiuQhg9Es6mvi6xsWWVjoFZOXxS9kKgo1za8z9+Stua+57+FDqIFOPcPE+W9LKQ6
OO0yq3VYt5gNQFi1tU6txSymKjK8SfZz0DbXxpsRdjcBMo2R2DC5nmT/oM3xNEfI/eX6hWTIbvH/
qLVUX2WHV/KD7Z43Jl54B0fUVIE8v0oADNpdM+ZJQ1M2w/j8VI5MDjvfEpTNU4Pu9jLSo7HXhtQM
/KG2DqSXksSjXe7Xi+pAqBMSjlgUkKGQRvwX4hK2bXjjrfWqdSYPyjgFLqh5yUwGbxWG4BDMFJrt
abYfGpK7UrcKBwriYbeepwgVFo8enD8CNODmD3xQuJK8TTMiu+4aIV2U72Qe/kjUTHEVGIBASZ1J
iraaBQOcbhL1WzL1CRQsm6km9JBJ8kArB3d2U8ijp/Gx0/1IQqiuoqEJqfQWZ4jNPCTMrmmJviAp
n3rJ2zJf7D1TTMaOwDkS6XXh1OWkMeHCtfBguDimyVTfzidW3Mu2bX9Mdn80QGbEDrbYuHeqmQS+
B1NI1KF6bDhPGpLm1YJWC/zUoWsJrEO4gzUw2tvYWgZKTROKpeDUKHdsh2Uc8HUOFuadI55csdsw
MKE0C05m0ITWJG0GdnFzabxiBEHcRZTcT6nohTQPpUu5STT2qanGjZ17ARoGW1BQZL+rMhooDm3k
sQi+GXiy1IEFnurlz4FSSrxt9qJhM57zMH3fFURWDR27BbeUxh3VEDQ0g3G+i3WbDeBQSGuK4veX
UitvN2oFp9wEscUbgguegk8Sa4IccYalIEEgpgPleAnGJdT69Tv+Wdw4KDrkGM2+0d1P3niIT9Gb
yH1Is7iLg+YAS9iRidtmAe+jCMfavYBYbEcpq2iegIh7Gidu7nM6UllRDnKUDFnQ+eVUoB2L+JHl
JSWHt6GCaz17gUn/LjCRp444D8cpP3/f3oZ0wcLJXvkpcn/VEuO58hyh5N3TxK9IZhU/BhhNBveV
jrq1srf78yJQSgZ2sfP1S+Tnqbau7qt4yuxWRQxStJJIk+QMVkQSs+HfaL9s+MU1kpoDXUhtFnh8
x0cAuPHjJc5jai2esiH74zSNbh22FqdxwG+mAvoeHF+oWzAiwVsoMP7GId8bs16aQ2R09dug+mzF
EyRflP3TRT2XEfdif/KddHAclbWBPIdvy7SqW7NW5E5OZidU76YkvIq9J+wmuzbTwGw3T6G+b4sd
m515h0TEX5uQ847tcGED3HEfdFUcZ3clRluaJdS/O/KQeqwBiRAiK6Y+Bco42CAOql6Og6E1fMKv
DqSOWZcwTBzgl4azTllsOQAAlkeCDYOR44CoG7jJq4gV6Mvm5Q/e+sc/Gj3pPVpObvuTI6ohmT5B
jHW7ATeyejzKfWIQYzuoPbf0erKneczvKTTvtojcSjGZMps7Qy4OOKWRsh4d0HiSeVdB+IwMccjC
Z9OcuayvZ8BV5K0WzIlam9YKs6YuizMReW17D9ICfu7gIOoTdhtNhl0taE4K87d/ylVF790r24OR
Me5n3HxIecDPP3GTZu9aZBSQo6zqeaL4T7tplcTJKE90pz6c09tPAuybqBr+O7pJQ9Ndw3io8Lqq
GkDGTTX22iO9+Z9k9T4VoxCzW97vMIobzVMQ/fvmssnqX41j9JdlaD54ueCAqJEVoPlpgVzvKKyy
9hM6kJYuxy1VT/Biz3lCVSG7c5FJFmS6S2u/M0kWpCwZ2sL0UKMbnjjYMe/7Nzcvz+KeXq8KcpNZ
IEWDlzabDdGC62L6cDDeOlbHUVNpEm4oSrZ6oHg9Wen0AnxlMabW7vXixmYoVYXnxQqAMpP3NwiW
HHSWM4pGpHKT6MVc897WIFDe9HJ9Afb5fRE/uB0ZrhW0KgEqG7xVHljxPKBGlmafibcW8nhojkLR
O3O55EcNw2aTKqs6oxxKNCd9bg8mmOI+dFaOk2PWA8wwEHjJnfTdMtisfy2eiWlQFLfAgHJCuCVQ
h9odR+kelKsUOve0ygtF1PrDujYn9s2mcickEQJga+pK3EO9AfdVBW+3531yPfa6WMl6oDKsvsfF
+nTbaNLpcziMhhoPIZVv66X6Pd+UBZfVSocGLj7EFc0R7ghitd1LYt8npj5wqL2dysiTClUb+jbf
1PRRl0KEcER+5EgjZ8w3Va7nFPGE4imGIuBXk6nI09znuuJMBLf8/7ZqEc+FFdY/42K8CQAiUM4t
Oz4Y+mBA4gvP90cDAthyz9wvo4Ci1oxK2OrGnSfeTxZtNTJdXBZsh/YYfVZPfJi5Rh1JxDkmTMPA
OoYBBE++EPU5X31MQCIpP8zMVnh/AwfNAZ71wYouZKXGmTiLkz9AsbnAB0LXvufOK71vw70JT/Ke
sDE3a9GIv+7Qe8qEIyf3VKoV64XUK6/Q+Ii7ozxgaIzYhmU7nlw1FK1KTW+JGeSiDpsRC2T/+95X
1YnjW3mdCrgJ5Dibatn5OVPU2LQeBc8NebXqg1wpJt4nxy8OOOzRHcaJG9w8XpZDHVEMmQ61gnQw
eRX2CNor+UnDwpbyY+weF6tXD7eF1miyMs8VC6qGEcjBDTMAKHpsH10JcvHcNgYXYHsvqxMXw5Ij
l53rbqAcb4UJQMi3i6g5srQkwGQ1V3m9gXzjqjm7ytLumC0eyDLox6RlaAR/7rO0kD2XWy6wSrvs
EN/uTqhgnNN2troCwGjXOzxamkPeWXPtIgtPd14sHQEFawKEdqY7rG+VIDWNDVoBvV6jTykZGC3W
Lbkaj5JT7TPIo0wq5HpvUYU9ov1E4md3NySpsEFi2rHUahg/i/wLMS/m+QIT5oW29O6TAWFWbWZf
LFzYXjnIikSzLjpI7BvoBNDtd1CHG5TDxgk3bxJVJZo8xZ+ANzP0KvQTtgchgXuGcPX1Qp7TSeMa
ATXH5MJ1OyfpwAOWpZMB74LD30goWrb6gWHtMckozpfdtAVNmgDK8dvG6QWE2jLnbNlS7GuVLYL5
AW7kV2QOx9MujMr2d8p03PPXFvYdk8ilx1A31L4EqTVa4D80v/nLqHhBVr2Lp01cbtTcFm5erdFX
yhhy4T/8ZzVjUzwXRPluZqrb1q7P7RhOLUdi3HDfuDOzEdstAwiS8Az7ULKw+Ktm+eOJjCIjNDiq
OwRLN9D9IbOrGSEpOmY+y9Qg2IxDWahh5pJNQ+kXyPHpt+QQ90WXQknAZMns/oulQeZpdnluLa8w
5TvzIpbjnkkc0VnddrRmmqmBNZal51Z3/yqezZFy/Yc11tmcjbM4iq2xIsuYq38sda18YUvjInqj
zH+HQE3R1Pzgn684UfzBUrcRd77B0P9QJvkM1GtB6KL6T+X68NKas6gOUx05OJI6arASDZIIkLLj
pUO4hWBNGfgaVCCqa+bus54iTNd9A88fZLWU9FMiCJKcMEh+dL/DNcAoJMRbbZK5pMIcQNN8vSfZ
ZXPU9mgUMybKH3527KzK84oC2feb7Jr20es2muo+XGUsBbgN2iehRkCdrxg8L6gmIqCaqNKjvz4R
faDsfYf6uRe80KtZabOv5WkIGiWWzuSqN8Mo2+gWeW2/h0QZcTtswPzqBdtEB4zrbA1N7uFjdSWh
GCbDwu8vb0QXqG2NvUmqb+xUt3Kk5X6aiMGn3DmayhJixv4lU1ATWA5OoKahBuTzUcxE6lkGrvFi
1d5NfKqZmRSwVSsWr/NRKhBE4Z5gpMGIiyreDvT3EYqs45Uy+j/tQuiPjkc2762imSF+HuuU5TNo
lKb11It+rUG1HJt/KllwBaCSpMHRDHfxTYMlC6CPeQs+TVXZfMxmexu1Q222jbDMSR1xttzPDlTO
xw0CjSTSq6/F+sx5ayBtcrRL3HTDicdbUM6b/ixsTL4YYvCz6PJXt/uIVhkQqaCX2hjHdWQAXyY3
qTvwEJYO3Q0dHZW4SZ7Vm4G5pb0gnax3PqBCQj63ez4SMkuNChsXoml8d24c1I0eRLOnGPwfkcsj
kPdvw+lz69KfSDLz62lxY1xxf/iicvtnO1TRbTAEncCxywS3f0db8azz5yItPFAKico/mP8+Q73D
NuOwn38Cd85k5tMQPL+F62ThmOdUUe4GZNg+KZFEYSC0Te0lmEhCXOUnq5Pg4To3mp2gLWQNP71j
e/pBWfNe10D9ZOsS1OPQJ8ioKuUTjRyGxzXzPr35EVy7Qr00yooU6hL8AF9hDxCr7kBdGXI9pT2z
YYMFCzpBB6btu1IQ2X63zv185QMp0JZ/6r27OnQlfdrECnszOFuyUbhvPhkJOQkRGAIR2iGzGjOd
Tc+TrarjSN2+r4RIvnjaHdt2bxew1Nr14mUfh+VH/nhnx/6wYKmlkylTQjcHK88wXrZHxYRLUQzp
6O9VQLsQUeF6ycfFcjmo5Dasgo3DtW+dPNYfyoyqubcn5+qAWzL7zjKaPBLb+9Lm5XXrNe8zJ796
iOApxn2oDKdKTnr3/7eJbV6vca+yz1uCtwsg5v2ocmmPk2FfVhvGgKhiDVxgtR269v+xXaEhyzrq
FDZh27vMQLECoAZZfaKtXxjoPc83dmNG6NeOONjjNVSbeLHG0HzPsRLTIPn1VdC5UMwnPZbGdXEm
LDBClZ7AeyI6nQH8pFDWoHv7XrDudwfyvl/09mLuMagMMlZg9N2f28RGp+z2gtIyPJybx33A/LQV
18pYHTwpPbh0F46/aTmi5yKEBWsVQYHUxCtxH8DigorsJ28FmFR8lCj7X1T4r9jTkOITmD2j5kAU
f2A0KmH+K8JgCJujCPcaDSsn84aJPyoAct50mqAbG8oFEuwhjAX9VmHn59PhKys4wn67KIVezV3P
d+5JBum/63Fhrq8WAl0LLFFqgvmXFMJTxfWsDDZ9CvYBd2wowxx8Xs6JtPz1NmArezC3/iYNdqjB
BHKR1BPqEqrrB4bNJKovyUzywdwnbeXsMHu7KXvds4ceo3x83KkG1t/fwiF0A+n8GT5/sYGIL9Aa
pou6EUJD+pgXebaTIMS7Jk3nbgK1Dnl2BTt9w+W9VImw1r4vFc7sjZE5fkj7ZLNyVn8PCYb3QzST
HBOAx9h9MYSz89DMl44Vu1x+W/HzEcnOOkQCpCUNay8UTKGhVY/dGm1lfkL0NQzLup+nQAywU17X
hKhoSXTP4SB5XaUmh2mYtAmNvYyBAUxbShJEL0HUlZXztGB6p2ENcS/GEf8i9rkKC7gfs+5tn1fH
OaQBdoRuArbZpYnvc0WmwDvFnuMhnCCehaLkHzqTrK22UeCeIbHVEvC4KSrEqWh4WBwq4xR68mcL
iCugxwk0qMEl/dSxGYSaw21qNcdpSRO4BMXsM4fMvqv8OF1du3ZF7Up6f2rKgiMnbGswd3h/hOTj
YtyQW1eMEWcyLlgLRHktx5V11w0J5Az7ewRO+FGQ5ZtmGRPaKsd/lXUyW94pvu/KAjZy2cdyQYgJ
wARjz6Hb6YMzpYFHAQx64wiFqbWpabgR8L+4377ME+HbkmlGkN7M0iVDTjKCeZD8AZk37ox5qmkS
tMk+k5n+cYoq9YsNfbHRMscIhqFw4xiAveZlS+ca744O8sL+mj5hcF5Tn9F6WHQtYnh6ANaIMp+u
cBJM1LYS3JU/rJZFgGfz5ZV8JQjPpzbHuIX3dq7k7RqTU3ghEwrkCoLB5u+jMF7TwNsUceeaBVgz
Da+DLtbJSVDjgZ0pyIm11ad6IDD0peu8grmmrhjFY/7y0aoEBK8Vgt/Kwi+mKuaE7JKnJ67PUlMk
4daqRet2n3kE+iNgAMH6UY7GjlZ1T4kmpeNCCHa8rxinEpINHq56eWbXUmN1d19BmxPmTwdh5wKp
wYNxCY0wKjYXrklRPD/4bXOf8O8Q4XGusTBMH5JogqcnEEK+rGF+A6loMoWBvGUkf0nw3xCAxa6y
YC87mucY0u4xn3KrmD1lLk7rdiMuYRekRTgeyHZVGF401EhrumWBAMyagoA+OCJJ2w/X+KB9Z9Zn
fTbqXouMBaE0gxu+8DmN1Rt8Uq902Opo+T+ridm4rHlp5CgxkmCR49fHhTSXNhROvv/z1PwrmNG2
xBIeDyAgLwQrca8fnMsFvC/XFUmPLrMhPUx+f8Z8JrLCAcYr31w4+Y9vE/h7zCrx6e5kO3XoCWJr
lPy1ThbeBvji9hcG63a88ZDQaxs9KDfZsoDxh3rfuAwEHU2+PFg9LGHLmVF8oXXLg+SeNoU9Rg+R
7isK2t6YTrfFWW7fbZ+XrlOZKDrrRg8KNRP0IfkODgKEw7gfnDAGuMVflHGMv0S7IO9ZbQn487lY
YQa1OyLqn+UJbKBZHeX9SGH37RIS0ZEuPST7d2YR7p9u2tX8NbiG4PbWKyWMN63Gw3qdlnfhc8op
VchFhzdKQbHAc8qh+jE2x31EjxKbhheVh++pfBkYcQK0qq4lzjolk/zVxeoZpszud5DNGjhkRFNo
OFEn5R3lWpJ9SKJf9xIpB30VmF4JegoE36cpVElWtjqpyic0pC37hpiNlakkb22oAZWJB6PnY0br
jrZpzrwj+ouwW/cp3un4PfHFdvtsXKfqTfS7fipaPgzOYwgYcwcGWN0oPhTwshFfpMI0G9/4b7v/
3Uqc25UZnQruWu1ncCDF+MESHc8PKpURmQOy3s8/oviwO4jN8g+ZAlnicy0iCVd1sPLmcz3UtbQ6
KMZbqlncomHczvMjGOpY0dEddaXTSvzGt7CzrrrtiEdkne1XxDK30cnEjv6LDX1acmz2A8RZAwwC
J2aPweNCgPIos9Jz8npga3ChrGkm4eZOoksJhlgGC4hBYJkKqsYsytLkqAXq4cT3RaUI8XmPzPiq
TWP6qXsCWq6Y8dMlPCjPRIbt+8uiVJvHncs9pnVpop9SSxwnf3/cDtUjSisgF49uql8NHo/oajwg
FFvwbxWpaQi4ZQW8TQ7QjC8J5w2/re9CAiI+yButSCqYaemKYKkmjrfAYT5KIi8th7ZTq5dJ/Q7A
GM2YSDUvKzyMHDQH2CKjUoq82D5fqLi3jUDEqpGzcYLqwAZIOd+dfb4guymd9aYHXdo4ohRR3wnO
cqxzET80Mph6EkIDRcGsqzn0Dkx5d0c1wnab0CSYHfdS/bgwWP6edWoCtRjSyxxxrYdiYGEqWSZM
jIREO7CFZ5U0b/7bKAVs3ez7hhSoLRHgEaEaVEPqQQAO87e/GCxoekOf9L7I6p7z7c5Rr7HG/DHy
Zh9BjSC7i/c6zPd2Apg0/fzK+NHkaOpFhD2vtBY+4jjN+l6CEUSqVmHeRk/kSYRDucbInbuG9tgh
yF+IQWx7awOTrg5baiU6SGBWuDXMrBiFIQ1dUr1tvlEk/tidElbg018JQw+LGcIp5DVISd/w6s8W
LMJ6bf6RK6xYesXMz5pukOjUijfR6cWTGPxFq26/vHyL+Y8cX9kxDU/kTn/OCXDnyYniT2yIrdZL
aU6Yr4SgNWDOeRMcVwGEU4DuA1EsCX2A5HTPJTirQZMOXLJZ2uOfRCeKq48iIpVj5HGW7lYOJ7xs
NqKKJQ21vub5Y9WtOi/ydgIi207jydzHZwIypeHM5YHQuTupdw+ZjfXlqlc2mxLQtkm5Wrqz42t6
QL8CRnxyO8dpvgkkShSu7wk4++5TrMwKYEK0eIlo4cYin0ISFQRBTaVdSnha1aR6RzFSWnPIHnD3
pBlYpzE6nt2PFxAId9s1+UzyNr8xCD/FOJI2/K8BQQBrvEmGoBCfTW44mY1LhiApO6vNO+mCP8nj
AK1fQDTrARF+YWx9KmcWbMdomT/cgiP3nW/ZMympmxzQ8dz8WW42Zwty2lv8B/glKyXZ+I9MLoEH
pyfh4M4RaGovn+9V18LDLoTvkxnslVqIO8imzWUNtzQymU1HHILqqwzhrjwDLA0tzIYvpsFqE0Ux
uYE5GDWyLdMYSKLUfZEjMo3o7NEGzB3H98dPtzHepy7ZueW+V4ZcW+H7VXBRfncVLv97qX9RS3F8
gc3Wn/jcqRtEFkJGsLacPQ9SidKuvW8r8iiY7MJBqiEq1K4dloiy3dbtbuT9xntWJ+ey5VJAIurf
UPh/8ZNFhMUvIwHz0bkpa0n5Y7iBSpB/iDTBzCv4HbZbUU6oiiRogCndiBOF5xCiV5WqtCCHiwJU
mZ5r09hZ9rHt+36r5elkV1nMlQSm1/g1KU6Au0eNxwqUie0x3yWUa6fDxB7/fYY7MSpTVjBsXRnj
szh87BJ2/VFSxyiMHzOdwGMl72dqux1YJd+j3UJ+plmnAtgfk3eNu9Ol6g8BhietL1cGs/xMCgp0
z19VL2TgRORcmzYK8tb/NV5ku9nkif4Y0JiZnWNL1bhlGizqytlxLpv7QQ2Fcyas9g3VGMeYllbG
6QHt7u9/pbwtDeQtLo6gmwUpC8Q815GPIbGzq4QdsvHQnWXs5Yvj9XEyaxleEVahPVu4hW3ttuak
qQ1DR0ZTZOGRrtDgA0Ak5R01jo6NdX/o/vQkyUg6jf01b6BoTjUE5si+cin04znYw5I1G+usD6YU
EkhRgwXI8Wg/dVOneYOE4uz7e8uImnOxVgXyvm5aQLwKppp3MV7WmEh+9+p2gQQ2VpYcQ92NkBvc
Df2ej2mlBwES1NlFB80dF/LGprwUuwmMY/FeZT9MZ+C67wcCTl48xZiILSYmZlF7BM2s6Q8o20Fc
1dgYFuAf6mU+PB9O8ricVJwcbPZg/bAdAlF5mOeeBu1lkN/GucRZthoGlQ7funo337nLkZQDZwVn
LXi66EpaZ7M6E/cwPCR7lcjEdpO6qg8MsbFokMNMYne1+PnWso6A3QBR+x1GLsANzKZF7bC16dGJ
Ztn/R2dJr5Z/CO24ChdZqdWgTfp2ulu2+M3u73AqoAqBKhkemrpT56Xg06WkotoAxDEoMfpfqo+/
CakKU1zdo4p8avklSbybdV8aq0U3+NoMibOXcqq4/yoNUoZegsq5JIjxG1pxfiqWvBabLk/nCaW7
vHxGUTOfpKXbMi5oSMSXVsRe3FJ+GkW3nslRS+bYeKzwY9U7rtvlyg41gv4dsUh1ZwxohWdHHmRz
kuKKNTEMqWKRndxzIq82XGIBo7fRih5Q94T6NWdnovPBqoMjASntCJaJ9spclIyEBsv+lXRIIyus
Ct1rkxG/pROCzFs6IbafRcvscKAuyluhWUFSmKladZPInj7kB3uFplUYg9M/PPyFsOfaiYq3xLBj
cMy7TWMd/T//Sg9ZxSHRzcsPqTONbsuEf85DOybuIc7dS8n09eTEpAcgye6gIv8Hno+zlNFLQKVh
qc3mKKED10/32+1NegRMViHuiWtRUZ2rkjIu7iqy6enmVtMoi+MFLdtxlFDRo9pB9Syh2nwR2p6B
bT0OFJ/5IcinQQNhldQyD/QWXXOyNfBPv7H9u8SBEJ3cLa4cQVQstPkLigAG7tqGI5IWpF/knTzT
Uavbriljo/devWDOO3WSugLUyQq0NtR6uE+OAJiw/HuuJ2+tFCVFYcZTOD5BXAbUIy3DMTzLgc4e
hcJHJOLhOeIrakB7OC8Eu8OU9RRyP19+l96D4ip10+wW0JsfEjqMORPKk2JYfHxA+DrZ1/zIlLd3
Bkt+C+4hKZRnfE/Ne5WHzFDMSC6wIU6ZjZ86zeAjhOQfgXiS3qEtrQRQhPaGKSQTj0VwbAfj974H
bp5bVw0R6TnEsZbTwXz3GlBWPvbp7S3+bpTatndlPONpS93LoF8RXrxwE8sVneSdAVh/s/i0eIy/
qrk25zY3HSqLGyjb82VROL0QTaN4NyPpHrAMwnFZqX/mTDwGwJPR5xUos6EVpB1N6XhVIOn+E1L+
x7vjVIXKb9cHqIc12Zx1c6VvYx/rNtbfOD4RUxSJXH2XxDF0nqpsOLfs2bpbCcgHmb1zWYVW8ps8
hXZ2/Vd2LbjQVFZX1xN8oZgE8eN23viOBVF0moVpekFNwjpitSf+ynTEcegP8rN4IWvBzdj5RuR3
ZViZ+Zp3YG+2M/nZVvZM64/I3SGhWmjTDF9RGrkOVst0cj8+65S9uaIaT4o2SB5+/+I7fcy3t5td
FCBZKBNVSGHalnhOB0i4bQoAjUmdyH/TEQkgkFCWRnkMGDTFWLolqocihIIBp7tIc4sgpWiQf9+N
gWH9Y15Too8hkSuqAtmLshYSG0L5pQ9ndz/jOW3KXN6sxD411V+6Sws+isSEWEcYCqVN1RYiuNGb
5zz79Cb0o/8Purf3uyn7d73Q61xUtLWck7Nmqo4Q02GiPq7Nzi+9iLTmEdEeV4bXjOLWarH4U0Cu
AWKCRCftNNDQ2F/WB86lNJnnFRkp1RCR8Eaw9/SwG6Ojfq0les3F8+kkCoWC9rIaOF3FrdtO8zMM
9DtM1xF2KZ+W3kIvgRMbemrQSATCFrQK9gXA3uBFw6SXcTQwM8Fw1KxxQrw6vIuc9hLHVKKIobPa
uWGJeYJM9Qj0rmgPG+SjwcQBXa/TYXK0N7DADNwEA6L06lRVF6u2cLBr+xhflX582d3K4nfMa5Y7
qg/2CIKJo2NLsYHMuvvrDqrLk8Ih907KYeNA0a3hrEZUalRjMnMQRWxDT3GfjQO8U5uQYZp9GNkm
bcYy+THB7P1r/LHzvKMDv/o3Et0IYKg2JKL4vctTL6+SdNtoOfzBqzylc5qkfhlged1JTugRjYnm
R3k9+bHk75KCqB3uVvk0EfsiciOw+VQT5QXiAZV8Z5GOCdFidBvd1OyKMGzFQywlun9s0wm1MWYy
1CxlM2D5EaJHOmci1Glf1wvkf5t3C8XcvGzS7TjNLV6v9zOhZ+AEr3R8LKryE2bHQpMXT3hFLJ25
atjUUAx5oj4toFuytI93J8phjKfToxTicJPoOXZg7V4q16aX95pfNluTvYgdH+KAOEfIFLT/oI7v
Yw24n1Yh34L6zV4RctD8e3uFbGDtA2qO+XE1ohfHD6dz0TSxUSPWot2zVcrQPUvr483l5yh6UwxR
jz8SjhNOTlw4XH2r9FuKefoSvF9i3ujfGE3aPHNZuEZDK6XkSrlkWT8oJWEi9DkQS0lLM3Zm58Il
QjD+LuQmn60T7p6vag4R0qV9tFq2LrXBdXbFKtKUnYr087lVLT63YzivuwV6/fsDIy/3b7/2K9U9
Q9NZe0ffC32EpAnBxPTl3M/W+s+WT7re6nggNNAxBN/+4IS84U3t2I5XiEMdtINr6c8wcUE4tvOz
eORhkmR0Av8J/0SsdhaewmMa949DGjaJ/8oPFEu686pMX1lNAg+l1IWePIt4LGMvow3QfufwXIV/
w4VXxKgqt8R5sIf5eewSFX+PZZ3W3+3ogV2h2jkqEfn09yBlIrkWIg53AVMG3/6Zpiq6q4CtlPLL
MyQLQ/THnisySnZcpYh5fpCKx7LXdCj/S10pWxTxdC+0V5SNTWGFqutq69n+wpDHnBbOjUCA7JpY
1uG3udFZXxDqw4h6MwZqqtqAtsSK/hBJGa+W0P/HmH5yHWn1xXwnfONT2+u+luqAKU5gEsEB5TVV
qvNzkIFTJBBXpluOCHnlO6fHBKjjP5aJ8+1mKmhMkQNHOdLucyKx0W1iGtrYobIwLb0i3jsLbZoZ
UyITun21nMby8/rHR+CgCbMEQzNV8xJvMDgeBzEH5EHH5A0ydh6GuaSausR+jr2x0gIkZPW9XBdu
AJuXZxizIVJfE3zZYGuhiweElsZ4fXYOF6U60K3oce7ElF4/EkHzIvGzy7aGA7MmpLlf6+yn/iOM
8XDwlbNq7RfmLJDojk2akNCVJA0zXgc71YDp2wKBLXNwTTvS56fYRK88NX+MOGqmt39fGvcjpFVI
ywZYBnPnk+HwY6MAT1KWFglzV8aulTNjSaWqHKBDRFOMpz8xTF3wicbxagDSRM2WaIIztQe6LCT1
E9gA1sIoaJue4Hq2fouLELDVZejM9D+g9QQfGMKWOSpakWe10GRWc3BpBf2ewXD0dKuOGUbZqeYO
YVPblVw8SbVKX3uWzWuaHIzuwMy+4X/7x0UdzixoOAHyACBWKjaeGTAZmC1cawvmK+Y4o10UCzhr
cv66aEsQyi6bvqczIjYSBkdK4jDvxj6e0ircYO+F0HnWZKPh9L2PjKk3RhBjc0dys7A5Pg0AYKZZ
/ETFKeB+xQQVPZ2beUPoCPH82bKbvUu8BfLpEi1sDUMQWr441oZ4QIzd8MIdUuwBTfNAHPAiz8Ge
21LbYljeurLDnhqlyboi7E5oojABAXsau78aBs+WkKYzUgnFhwnNd8u7/XnoFxH/FDYDX8OGxYA5
aZjgJ2juHaLquSoQDmHB+L/uLTfgeiC7Bfu5fX52sZdCgKxkzQs6+46DPoiP7rN62upPW0BThXJp
Yut5KE2CuWV56L3E9/caf29e40CJ9wqbSFheCCquAqUW3W7208ghWczU3dqfYsii7Mgbz2IGwzl7
jaABOwVlcs5b3pXdlPOzDiLkyBO1nWwik5hW40iZMWM4p/3gKkWOpiwJ64PqpoqoqWJUc1L4KIqc
yPcEjxpzt/dK2P4Zp93IUB+W5HmQ2/oxnIzeP3hVf4ak+CJjazAx1h42nXUCfZ/8FfHAgaibJ4aY
WgtlOInBYO8cZtBln7qiZQZrD6MPwo0VJ4FT5L1sNiDt7GvlYT2Ed7yK715J0C+mcWDhEfYiZP4+
OFI7Q5HkQwaOW7TgMOJpVZkjmtP+o8jPiOeWSeElvvGrYwbCxy1QhGsJPWOSOlTQ4GWGTbskjtau
OtAsrgwsGEIN5WbPaVtczRi0M3alDaUmqcAlovcF+Hm+zKstbZxzBPF7VwTLFUTcr2qCCYqA5gJ9
ARToRNDqkfGxCM/lVRDw7ItG6vDuEP66p50njS5isnL5xVc4/5jle2vWtbrAaJXuwF/HXT2zDcwe
2mVidMCfuipdbKXE9dUWEv4v8gTAHpC/3h7b3WcuGLZD/WFWX/eGeJCyqmUo/MoRn149cV+R5euo
icBabWYHtj1YDecnrx1i3GitmTm3pZUAm4nZ9MX6xcaUxrjpkwkne9EFUIGt30bNHlHx7MfBNa4x
GJMsesNfAp1U/0wregKZPnGV9QC37mou5oAWFbfYEH0uCjUzSDrxoMJ3QqHFHP2K+NeJR4Mizaio
cEFMRACMU4buNCyNme04i2lhv6+HlstQLvS3
`protect end_protected
