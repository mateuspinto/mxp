XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��K�-�d��8�<W��4W�7���P���R���M���N-5A��p�~E X�!��}��*��R]5>rULG�[��>�/�$I=�(|h�A1
�׼��>Ry[�j?�����B_s����F���WCm�޵�e��τ���e������Ҍ������q_ܟo�u��6"Ҥ�Ui?T��2��z4�ҁ<D�ǻ3�!�ӗ�o��н���'�[�f�a��J�~R�3+��Ǒ�o�L�x�n1=F���m��Pj�U/��W�^
ec���l�!Ǥ����܁{�g[QB}�H1~ȗ�Z�t�W�8^���>�s=iP+��B�OWϧ�+��uAah}�
�^��$\�q�]�� �Y����>z��V�v^�p#]�-���RG���x?#Y�R�R�Q�R����L���L���H����� �+�߇�o�Z�e�I���;ER����n��v�&WY��CGK��A��R7NlN�2��������yZ�Y��ߊ��K,x���V���6=�O_�	E�/E�G%���nq6P�����y���G�ox�A!*ˡ`&��Ն�L�w,GD��\�8�	]/ӝ-�@|��8���'6��*� �{�og5����PGB}�W����:��%T+�{�D�Dt��d���= ��5z	��q�vҔ����]x������Q|�S,��X�����5��Os����+_�-t��b�%C��rUw\�����()��d�e�6�������MF ��b�uXlxVHYEB     400     1b0O5q�ɘZ�Jml�Z�r����b�t��������ن��<;Ӓ`ήi
I]�1,1#7v=a��y0�TTx�"t��j��F S��]Ѕ�Mc7J̎lA�ҽX��X�'8;�k(���-�=A�i&R?AA�!1L$ ��k�')�nH͵$�uݮ��`̮2�G+�6+��ȡ`%�33��^DZ-���	`�C��F±Q�`��i�M�������.��߯<{��T�BK���:R<N��H��)C�&.x+L��ӸI��9���.J5�f���r��:;~H��y�����Z}�ظ{x�4��|��P�b+�*`�N@_������
�+;|d��H=���03���wX��u�jPN��R6�?^I��������)|z��4���jU�P�d��됣i/:�Yq�a��B}�m�����ϭ�t���XlxVHYEB     400     1b0C�D@Ff�%��	�xv��{t#�|'zM�ћ-�`�jn�*-�g)eHt�O�^�='ҭO+)����:�c0��n��P�PW�Uˑ���S��{<�]I���]Șο��b��]��*I>q��%q���,�B�l0��I/��y��p��Epj��!��5�"mm6��b.6�$��ˡ���+� ~ȓ:r�.�yZh�|u��1�n�/���`/��'���K�e�G���#�<!��X���6+�r:ɞ"�M���fk@2�W���S}Ճz�gDQ�w���WM��e(��b�)�^�'��0��ۀ$��I+���0߆ړE��WB��U#艰旃�/��+vEl��^���J���͉�����4wA� gg��;߿!<����ZR_�N���w���E�#rs�	��$�e�槑�<�XlxVHYEB     400     130����[^�o<��Mb�s�7���ϫ�<�@��gF���D��oZ�BK�~�q��6AD�q�rXd�������?r����P1:����$?^G.�Q�4�x�[ �埸|9��6\��Z�#]$�_�i߰'�Fr��P2���GERM+}]�d
-�4
|t�g	|����F��]��WGa~�w$�b3�i�q���'�T˭�j�)+����Ua�.{mC([3t1�A\����j9���W�E)�+�A�CfߗUKz�LbĘ!u�T�
��}��o���y��B�w�J�	��XlxVHYEB     400     190[�#u�φ!m�ȷ�
�]X��P�,�a��jƕ�����ve�"����3̚�%�=h5�H��udh��0�(w}��������A��u��茐���#6�q�������.R�� l����ȃY=����
y/ޜ"�/���%cO�[v�uYը����U�BoFq�l�;o>*gWOFSs��8(;���.�A��wt��N��-sJH��L���|�9�0��{�[%�rז>�R_����%��pŊ�t�3H9'0En|8|���s;���n�L�u�J��  �@��LJ�S�4�`�f�G%-
��Ŏ�H�xC��r\�?+$|�SD��tǌjc�N���Tȭ�'���P�<x7k����V�*�����kJ�-�dz0�n�Nb���XlxVHYEB     400     160
���C�LR!dW�A
Tq�j8nl�}�I�A��(
6?Ϙl�]���̯�pHER
{a����* ᱕'��K�(��G��Zzmi8_�'D��h�4 ���*�j]"��1�tF�!��֚mp�?��o��pȕY3"��b}Anƪ�HO��,���~���7eS)�6�06�թ���$�UG(�@��A4�M�܌0ho�9�z�֝�,#|���ѧ�֌��X�DC_D��{���s��y����j�B���t�"5�
7=m�fZ���ߒC�.�z߉TZb�#�.2Ho�_��B���Ӛ2hB�& z�-1��~���	��p�������Fj��|A���1�7XlxVHYEB     400     1b0�͇�&��Q*������QK+�y�s���X��դ\��ߵ�@�['�4�bSz ��9-��n�c@`�T����s�-˫���a2�|��zU�<5}'��[ɉ���*��`4�4(�O��m�ؘl��.-7�a�l���Jhp��%�Y��0ly���)��#��(|�9�t��a� L�~{
����%�{�Y���d5���@�g���$;�+P$�՘��?+��)�����&����m3�|��w!o++
���"�+��v1�׌6�3�������;��v�"\3e�C4as��A�����,B�I�C�@u��5�P�g<Z�;��bhsnv��-�JH��[�к�d���	�ws���x��o�Ȑ��{�
}�h�Sm�������Ve��zf������,�:��ERXlxVHYEB     400     160��_nUgE��7�}�`�h.�I|`*z���W��!�F,�>�R� z�S�jk����OT:�w>k�,T��"k\`�Q�*���Y)�=z�z�Q��%������ȍ�p��ߟ�d���L���d|tDsC��"���tYb6Hz�RƑ��]�1J2;1U+F����J��L��[�T	]M(q �[O�s$t���H�����9�Jr�m���J:"����1���7ɼZ}����M_TX 	��"�~i׼�:�JG�4�<V��pP3&�����K�}��e^��� ��R�$��#,�~%�֍:FJM���NL˜3��t�ӳ������G
Ħ�
ƜXlxVHYEB     400     120zwh���>f����k^���ӹ"�����(�Y �5"y����N��9�U-'��Ղ�.�F\��.�VsC֘���VwH!Ӭ0�0fd?��D�����[�B���:�NGNڧW�I򘁬��u��e����$U�@�M;�ٱ�;�j�Mu��!Jx�?�*OU��S��9���ˑ��4���b�B���{��M�[�v,�ӠV�8xc+ٯ�]2�7��J)�@H&L]<���n5eL6�d��Q�ܲ���u2ܓ����@q.�qmt5��N5:XlxVHYEB     400     1901�	8)8)r�r �C-����,zҽ�Z�<�8=*��`��/�t0��JH<��q�JScuQw���m-����6���A��J�%����7Pu��������EgiɎ�F��Ƴ��,k�Q�}*�D�,������(��������n���r�
��&/B��aݧq|�32�Lo 9�̆�jH@B/�%�k��{�A�<IG���yun�zg{������F�t%j����{T��.8J�˱�S���8�/���G�79����E�`f�!��܎�D��C��^,�J����s����K��x���;�����k;YM4$���q����xcN��y	�=�;�T:�G�n�Jm���1}�0�'�mB4��(��-K	�l z��-r�t�r�XlxVHYEB     400     140K<�p������ia�	�P"�ĕtQ�@e٨L.�Y�=>�C��ڂ~�휙�>�Y�eNf��.��˪�6@A���fC�Lqo
`���Yo]k��n�{�ٱ%i,n�-��P�u�cQ������L*ā_�|Y\�W�蓽�K���S]oԆv���`.�!R����C1<�H�l�T�,�ֶt�y�Ǣ&�=�gw���<�E��=���{tR��jP�˧��kŒ����C�)�U�?�Q#�,�`:�ղ�N�46�\4k9�i���$"�"�*�g��WILe�WKnjA����H�O��oH�)A�6>Yk>�XlxVHYEB     400     160���&���\�(��Hz��܋l*��3A�]� ֋���ǧ�"<����Ԭ�l����/g@�'l����_�i��A�̑C���c���!�TV�p�Z�Z�?��\!�v���j{l|��Z0Ř�p)
W̻���
�D����u��B�!7D_hPpW|��wYk�����r�s�Ȗq�eһOc@����}�^!�G�9�Id��Ʒ�u'����m.~�9��C�8���K��f±ϣ�ы���_[��3z��A>
v2R������U̓5�7C($خ5a�r�#!�,�]�^���}������p,��[PenZk^5�7���Z�������N乙���e�PsXlxVHYEB     21a     100G��;�sC��5���ω���3OtAn���x�~��O�h���-���a��&��iଆ���5>���,3x�0�H�t'6�f�/�ևG,�.�13o]�vWUE�+�����b�&o�q��V}��8���zFj��9	(��+6�h�G��+?\-��E������h�J��,�d�	u�`��ES!+(��R^|����wB[E�0Ĺ�@����j�H̐��i���1�7�+z�T�S�;~��َ� �