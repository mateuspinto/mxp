`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11824)
`protect data_block
sdDuCbgtu7Zr5rdXNPbHG+W3J2J12o0nkQREwTu0ZbItEsLuuHahsOiLYURxqOCiU5mmNNUcdwO3
THkPBgybf8cOfwfxgItQvuRz/1JjTsAOY8YkCgLOqgwC8pRyoXJPkpdXWEsbYz47OHMFXd62DLLe
0eUq0bKQO3YU6aCA3sbg88FUu4BYEHeu8H5ZlPdvZbPpEk6Ju36M8wR7s2FTBxw9ROFse3W/Oum6
GyY8k5nDqr3xeTTYXEaHIdEjcenT03XSoBP4rCmQFzORObt0d2pSpvNnPuXs0OQwi1papWFlUccl
+U2V2vThWwCJrQoZrrxPI6mvRaU/ltP9Hfl8n3cDWaSUIShd5ntAY86bAwUbYG750WjhgPN+8VC5
DfbojrM4KPPEb9x1mq38hWecTDX5/Tbpj5E+9CMNHvM30TEPwlq6gHj0Vg5javhr+gMRjvr6KLyE
xlIGyWMB3QrfQcK1ltRU9aczvx96hst35LXneB9+Krsd9YwWZGC4YI3XTvSB0NXC95NOk8aBKxy+
9pZzoa/AaDcz4c3tL2MitIp+paBAfVWRu8wm2WHJNvNnVJoCSTV72Pj89vvnIZX61BtVafm+kg1w
CTwntafouxaQV/iPyWxk8h0WvC6Nr+Jbcp9gRxtZ1soBOt9Ud14WZhSr+u+EnT/4TxHrSASX7rcC
BYXTx7TiMvPtbYFw4Enr5MXHkRJQypXdP0WL5j+clOuY6iY6RU7KldQ1Q2PLW1xdJ+FI9DX8fJCy
JBWVkWqLRmoU1OXyDLMR1TsmIM2X3GdN/o21LwMnaNlYxybCeeAQZMC2CQuhXjmKYyUvZots2CVP
qGKNzefGOf7EEIGYgDbQacio6VRz+80Y9UNSZFzP9ZWIzGj4fD/Bq9gtQlEKYFHpy8XDRqBPdYw4
fdyj11H/F1PDbYXjdWWnsHYUtcD7oklPBs7eh3TH4qrPCStmxJm6updOgYSgzCHs6NVX2HRwWufA
rPc5hobE7Flo1EATYKF8qmVtS8qBMyBDbZ+F8yo55r8xfnpqhf9pWTr9jz4fbnHRC1ch0xyBQoFU
8JGAWyxjLWWOVcv2qWGWm52dOUOygOEplByVwqOzFCY8D/316DNYat5OggL6SC0o5dxTz+L+nCnG
HgQOJsImooecHFRMQdFLoZQVdWyGxnmXNvAgBqRcLQopmNmyM/S9ZwiG5zGMWhidKaVdBXvFvOyH
sMlJzVGqvZQmeewNrUHb6GM85XiW7QQ8nnbM5xd1FGwibwNiIktGH7hZpgBOR/2CKonyIiM29FIN
Dkruk2lh7Iz7SJJFWvO+IeLF7hynyXjMNzp8qCobQy68rh9BGkynHB/Rj/D5c7XZKKF3JtEiBEHd
fsVYY0Q8mr9E91vPYVFEO19cr5n5lFzRbiHR7DTPMhWG7Z5PCl3/UeoIjei6gn3TZbodzlog3kYA
ZLJf58l/LI4qkAsTpr8EUVb8cUezveQam9r23aMHOtZyQNkCpaAk3KAcuOo6XiKuMUaYF6XNVM4w
VSYOYV18uyJLamG8PdjUUISGnK28ZuCqf4Pv9EjD73UvDIHlzJ+MVwascMumBkWnM5Vkisdixzgw
DwbTE/MeZ/psKEydKuj0IWw3ZhdGyRjEgDnaGncPSu+k122rsLqByi/0NUCbtq303ratT9p+fTGW
kC92KlV8q/NiBFcjjySEAHktYVYOi0WdFqlovPptgEqMo87iH+qR2wjFO5mCijZkfbWjAtyMs2yK
n81p8/8bw23dZrqXnfG5slW0jWMmnXcqH+qzs92g/Uti3OQww+3QTjROg6jRUniyNbPHK6LbPr8U
UgIl+8+Wa/cFat2UbscAWOQghL+XymPvrCoxVwZUqWgZIaQMLd4XKRsTNsvKyTgjEwz2iSdkCmoL
y80LP81dRQLkWcJ4bwikVDOxZAPyP3b5T0xCFvhVRLGoabC0ZkmHQvIgPa+A41ZGBoBhyHFtmhcE
CeQUc66wmPO+Y67mP97oaIEzS3AQZFRRR0a4VhRBLKo6RguIs8PI5zEca10AdJtIAxcZbD8cOmlJ
1Uwi4XkIBc68oSuMPurn5IKIPGBuK1IIeL6k7PtFWazUVFtH0wO77aaRSfLjpLLV6T7QjP0WBq0c
ddEfa7DjvnRSh3I82eBZBPvdrq/c3Wx9WZiVYSIv10DYhGXnq60ScPxQ3slHdk4XlOuel7RU2w/i
FjSkYiMh4cMFDP4CKWxJUT6NBrZJOopEmpmpWnPO91GKdUj9woNdsRGwxq8nSTjyWBo4Q507/t/L
yCwJ+cZgI8wqgjcwVr7sBoJUL9NJRBQyUQfwMhCTy0X74hCyDyv2YgF96GFSumOUgTKMw/OS/aLQ
gC4LrIoVWjFce2Xr1VZgzqBdLLS0TzvOebWRwZLY1GsaVyBCHOqw30lnbJDvWI88VxRDvcRSfSxt
hXX4eblOGMstsMCQDemEj2FaaM2IOiR7nLOFp1nMdUdIGo5A9a4ALpX/UcFWsuegRZvQnzgJea1L
xzKFHTCGj1L8WFH4AgKjr32bFwQkxsdtIEgNqnAII27ncJsQP1dT0yhngitALpK6DhovY6kG/zBO
sHjro2VqKFUoiaJ134+d2Ji73Rlowyq1ZqHXTYuP7fChP4ng1kdmAuCKQPn5DE/jSNwe+n720bUT
kCjYoj1s5Ozskc7CA2yfhiW1yyaLENbMPxoGVq8VMQoQNv0o45DCmwC2wf4jzFFuohqHFMztDdPb
iwhds7kMH28GMZAYnq75bcHXQ2zQByaFhu/KK16vl81NyiuDBaVOLakqiDWEKusZF0CjZQDMSHhV
KYZ8pQQNsNdkL8EiZnJIY69dDFDpILR833JZ/TVglVRyrTvCFeB2mf0MXBkdH1iuhJYFY/OYAJDN
0L8lp9KHURg/n3Ci4traZT2ZIw6docOO68KWXp4p9UK2mnGe8Je0gen68cEX/zbS5OMpn/ENeWuQ
/W+uozKa0DgGK05kfz+9kqGbTfckFwaY1zyyKRTHZJ4Lq1IXGYxS+hEBs3uh3GTU05+fIDVQ44si
KrBLrD8PrW7PRdQX1uvEr6qO7G6arDxsN7AT8s5DDXk7Iuc0EXZBbBM6Y7X/j8po7l7bC2gfGN5D
4TXGtHKk3Pi08XOf8u3o6qwSzYqtJDLicIAOITUH6Q8yj+VEslRQ4Eop3+GJPMs6wDgdat7bKsvk
3smyETVlDVB7XBO28hFnBeQLLmOUybKW0c1BOZZMt+z28eQIpH5C+HLRClj35qy+nmvT6NWdc6+B
xDkZ7CKx8/omLfUJS8u4BUkIXWvtSi+IxHigxuSIwcrxNn7eH+D2FsGMswalzN8CPgOGKm1NNpb+
reV+lastV3Ok0NwUJPLKzPOD+5X+WV6/9/WAhAneykArA0Lh46pfeZQKMYFSnJsN73Yuh5TByvP4
I8wLufZdVYXO12ys/1/MpIvpvWhZcVMHGOVhfHd8M7vGO2iCy9HbANO1n+bHMfXn5+RmcvB46KNW
0kDSw2IP5YvGHVrL1DYYhL8SqgCEQd+NNQTbETSsl9IHHrAb2aUbua6FavbeosUelK/Rj5EDdchd
hGXJTHbX3S2q9TGNYz7ADmBXD7yquEVoWMDphVw3c489hbxj0MKMRpYglXwZhhlqswZqHjS6h/LY
dVIhQxzksCZAX+ykTtN9tTbBZ4oGCVaHPfvWcz/iz/BDQdG1PmR9EQkR8YACR4S+qdp7UeKua2Wt
Gz8ULmvVxZbjEE1JeX+wSd9HwE5Y6ilM4ot1dQ+4s+nQIQZWUUNgUH4s3KfcSqs1RIeEAzAKI3pp
SbV6alF9/SJRvfwiu5O1OfoHDEW5Kvasm6U3ZAsq1H01h5PrU9MS5uVCMKNkKSVSV3G2FP4W4VkV
lhfYFTKVtnmVLHH2SE913aJnDk3MvPjEgkTXDh39ovavifim/3zh55mq9HxZSItEUIjVX98lSvBq
HvT9OKXxAtAt539jnKOaMlBTMZBLiZimdAG0OFfekBxEV4kZ/cQp6+rlqOxhVjNmrOqhbmPkbOXe
E2rJDhlV+3exqi29V8E33eqHNIqkpvoGzl2JAOJedsTdGuWoDHkJ/7IAdsigVCIorFJrwlzqRXEu
f6OLMTfxtSKAAV5+kvaIbeUBYmtUq689gmDVRL4wX+RB/IKdhX1CbQCGUrH8cekpw7BqDiL0DPAj
MrnU1N7ooWx05qIESDAqcoaHJHMKSmE4e7ZVIxXMPzqRCpDZy92qHRvZ2oKLokpi/Cr4qZXbC2VU
Iny7zUrrrs/5I6pwaoOoCvWWBattcrLWt1uYaVF0tE9PUOvPDq3Rbj0mQTosVKwYpDkgWWETfH2R
w+ArWCaMyP43AwV8bs81qhm04daRJLyw9vMobImDtlSumBeRyHa9URofge5OuQGQQMWb2U27vAiz
1PjXM1gt7ethqK2yHe2muBUaRaxiDYaYcLqXPDLCrzfD5a3F0AXwOY/BUxySBwqfP4I10X9qNvDt
BKjuLM1Vy6sUI3DbvnLmzxXOgZbBntJrJ5NgftR8x9sQhXcQ1IzVEDwbls3uBRd9MgZ1+gv0zQq9
RMkpT8Dxp/DhS2D2kY/bYbTi0hWPorgJGUvlrVyEhKzeAIofmGeTEYczkODc6yTHBWj95tQUhpHu
otxQXNxfQ0YSi4jQzUqe54riDSZeTKFZtT8qOMUsXNy9uzFKoUxXwSw4b2pL1XxjXxYe45GMd0oF
bAc0+zBFy6kwXj6eVc6nsCRaWERZ8Itj8ttPWnWVYTExaUHNz+1L/R1UyRXSuUS/gWYJA/VQimzZ
r9gwBsqCE7ov0f7MHrS9tkIUdHptSwWk2YmTHxQcVMhcZWql1tC8Vywf2vkCGxUMiUZhUa7c7E/o
u2TxvRXHeCjRB9wT3qeoyYoQ6rLWhK12QRhSqiFRfGoiZlNMQBDve9W+3vqRarnkL6v8v4GonTkk
xD+KcrUM6EwNMXTbVrV+WHdC/Wmzzt3+CUlRsb8A77uQmEKeA0GM9DYsmoOmwEvq3Hj/sGmj0Ms3
WDGfsrBlnObTWwIVhMvFAPuBcsTmn0XL+D7Y3dm/sQJ+pOg+Hl0W3TuG4GPc24fyyiF3vXbejMNC
BEiDGBTpA/786Mq1+eNryuYbcqFRIRxXzO6oQ6ijyJOMUPaBXCJoNqW1yr1zhGmZ8f8cvKQB7bF0
Gqt6WM2c8cAlZC7xsUd/vRe9Wd/iU7tYdroxAVkyGnpW4CM5xmlwRcgO0zMYKEDDyzohkljbIC6Z
9EG3GY7SJLZHvbT+0P/50IpscV/RvPbwYEa+DDvmR8C4ec2k0G+IAxj6gFUUKdtiwKzZG4t7RzEq
KRpApyLL7xk4zcSWfQKLeIQxcpHaS3+8uxaMK0egCxrQrdU2AYJw+WGtazr72r+7wE01MsAmqnVn
dzAaS0LEZIqLKQcAIt0N4s9m+eB1ObtX6YqCusYYvk+lMyJ0rxgLHftt1c/ERyNFUqZlLZ6lnlD1
NOjrdL68n3rjtGUZIIbBRtNqNhWj8r+vOM2BYojrO9v5/8vXfjGou8vci/a0K7CvIj3FoNEfvmmq
zGYrnSJ+VscuwddzGzVs8Z6IZsm7YL5lM3G1b6qfbFNDVhQszovim9vCtahzb5XfKoPj4cRKw9QI
9NvlYtimjfS8yZ0xacbE9mUAlIvkYrqO20fFM8ERmeDfIroYLsmKm3LnGnvUGnJpUhE9R4KkGr5n
cmsj5BNW7KzhUpkx2bu+PG6wv0DfTkHL2djLO6UfHyatrp5jDKbujjGNuDTvxVSwMNrXh0CUsocY
aYGiyOJYqN0VU2u1l4JE8sFpzsXdvaFouPphha1vAjBOItQjz3THkTXIIDC5jg5Ocs+fYX/NEBGJ
10NZcB1BlwmNpYccazH9bPdl+g2U6aGnk/4ghjNJzwxkUVioW6kog9CJ/GDAF/okH8hwp8uXm7pM
dgAklWVY+cQ8AALlWOKamkhbiF57dCD1UTMWEcJ6L79L0irDFgYMpfMM9SubPY3B5JdUtCNR1U9T
4Fa6pgj94DVJOlDRm5WblqFALp5A7kcxYF8KrGF3O1OH9YjF039LyWOYF2ocNt/uvQISJTGxqyZ7
LKpO0QaB6nmiBt4Azb6UC/IUxIjdMV0Vcq0uTOJul5wqWSdxaOjmEu37bFPOcYLCDkYomz2IBs3i
gM6FYZzdWLQ2147lkG1ZLwq+ez23Q3o7CzN6WjImocO52dlYmE3CYAhcsFKjENrvIVfwcDvQwM5M
HkPyGmjMeIDUVw6WBP8ezSUUCfV9/ClEQblD8LOgtEMn7ql5qWpXzGbRZPKkHcJXKG+axI1cdjRO
IxWWQsZ5WghHskxXc1Eixxgw+wzsg9rVIzdG9FS83vCiQ8N1bQohsyGi7LwpEEym2AfnGlsfcm1Y
g7/uJFLbEhz02+lmByNlrlLq2vG3+xfma1rFtEkLhzLTzvq5hKQZmH4acdMsjeVA4W38ZVjF4Fia
pQn9AsaVUH3WQsK0SFZIEDDi9iI534+tMtu1WSdHZwFPX2c9W8VkG7q+Qzo9zZ+7ypojiQ59TJh1
Y5nCoKGCUi1UoX+v+UwzBpBR4UPSQMBtNNvf2bzSLaI38URspfoLmlvy2PephQLsMuDlSg4kp938
+XfpVSVspH/47MSF/ne3sGnQbuft7cfBNrYjgQk0KhzeDbBzkckwAj1PS6VE4biavjaGyFm50pPM
yLMsfkDyjmjOvgs+VHN35qSpu88v7rjmoLRXp66Pmo1DSfMlhatE8OpaGXSKPecIwcX6WPu4qZvM
nY5RmhLw/7OXvQoz/p4+JpEjVcjcdnDzFfum0/QjPCiKgxUXd3PdBtS/6lJ7zjVUhYcSWkL59aqx
jHJHP6D129HCosuLEy8crHs2d1h4eNqP9dg7Q5tM+nkTqeuPxfv9Mvr5FLO4thMZL6rL82vasWqx
0Z0897rC6ROsxV6vJiXgSdQ0kT+4Xa8Jc1h5DwlixeYEFgX2kFPr7SQcULDX1HLsvTBI9vQDDwbL
VKPaNRlIEv7Hn0jb3+mXMFwZUUaJeORmsBENFgat0SCbq6eAQg6chDvoYgYlfjSDqXqKLkOrviGD
Ud0q7vmDyXsGmuvOJBefjp9d54UjqS4pLrItrnGQModP9nI/l8wurMKftJcon+0vZ36Enk7+yRJv
xvfrKN2LYW/1yXXngjK989/a8Z3cNIo4/d7eoNyF75rDfUTKgnXB7g+fVUUsCKv/DK57cloKPiE3
93OXTYu52EwznI5q4XZCZ0r/+J5PMnadjsBuOfuVu3ER3CF+sq1yhlaYoffzFj7EH/gDqX9iI8nG
jMCGfZcL9JSSLvoL74TMcJFRVfwm3iscEVEM4XvCEC706XsscBizLFCX69PignDFjqZqHAOB4Nze
hj8jPaDIdStQKSdbUagdoM/VIU3Hsh2JfQu6LgWXpYJ5lm5TuG4RvFc/2xKJE6Jp6W+Yrsh/taT/
FE1pTLO4c/ZwpZM1lB8dRC5l8BbXTQzepZfYpvtjS10kK9RFlMz0xcZFmUh6K4NFilLd53Ih8cWa
8U5JholqECPl+Dpfv8G3cXTW2wIRflermXUetDmMOndW6e7KP92yCRl6MOmxM1hV2s8iv1xIawHe
DEMZ2k4f5bqCGezIDLn0h4wR18oeJNJ3kOjQ4aWr7MJyo0Gu8bDZYhi+pEizVDB8sLjIpureiQlX
Fd7AZXiuCBvsOfLkGy7K88WRSSe4CYkL5WPm+QrX1P6R++qToqgZvz34fLDx+6CZaa/gzBpPLqox
cI1iDLei3NLKwN8FDJTHgPVS6Z9COsY5AyOmNBoScoRHVpr8y4BqjWiGzaBBDqJOOFEMsLUmIvAL
gao8xw9ndcJNdMxedVkHNTVM6VqY2ScZAxTth1OhYtMSHgPMYLUkoNleEbLpDpnIDo0DlIfgr/De
jQ468F6B4w34zT+lfYOQSaak0LcuF3WMJCWX21I+aqfqRS3Q9MRfvUdz1Lt+gpI3UJ73eRAP7IZU
TO4HwM6QyH+YIT3/j4foxsQSXsIAXbOYB4vBJjyt4hxPd3Ok/XtqxlR5L4Oez99wowgwVTGi7iDW
11EoN5zusJ4Ta2BQu/loyH54uHZSCRIC7JTes8444yD6P3NumWdvRVwngR/d0O/NmU4+RyE3Khae
FowRWjmvPWuxxGSgz4bFHMpjhhlOUgAWgYnlOgAomYC1wBKwjcEKpJi/qQrjy69p0sKt4piln+un
c60Ym0fKgKNRHtG6tGyrkezb9PQRwyRV74AJJ8fH3aeSQA8LwvpghYcqkM/IPEexyuELWUl2ERvT
qhoJUknHjI71PtwsOKxwMqqvAF8xcjsQ4zWU02wvmh7zzZaRCF1HmA4C5BxW1Pmsri2sGwOKWY9b
YxFAoQenFCkgECmkkN9byfJ2CsMYEwTZPEEXnTQoAxkdvimWMq61BzUJa8W88R91r8CGyapVwK9Q
Ps0lIRwP16tRfHlF64zWBRK+/h4RQBXDEYNriGYat3NIBr/drGIksQ7zc4CO7BZLbCjHxFldT5Mq
rLlBhh/nmos0KO5APs3ZA9u/Ux9lSVHqHoYPewWf7DaGUsraqNYrs5oxbXWflyff0IPH38h4MIO8
ePaxbLiH0cvhfFJ1VLgREoYQeTjiJ8d/OcdYiA0pzMM1O5L196qzovai7DQRo997OCiQHJlB/tP0
2rmK85ULGVdVbbb+FJc7KxGWX+eG7lo3abVprclY0eZVHPt7L5i3FWQX0KpVVq5d4qGFh05ur79O
btoADAca54RhznK/Sg7CD4bc0IHeHGMvL8Y6WjwMDYORvFVpJWBDkHDhBnjqxP4ldY7yCELTF1Ov
eTXNo+qGLamRE50lCc+Srn6pxcS8PX+g3C+nMNu7CqzbyLXxtsY/MN/q4B/eoOtfn4Uih6kqZfGV
i57KTGEd7sFxSrSOrAUXziA8lE9jcH851jKdgMGOAyDyOVsNwnMNb/zaz5eCZSO+IfvBtIaYtriU
2Zx/V1jLuQ1z2cd5IrpCumIy9/UVx11hpB78LFlZ3pvLpI+TcZaDke13ly+ZcvGOop/UyZ3ZfQ07
rjB9qbscrjg2R2JftJHCyJP/PSB5gmbDDNxRNilY89B+bObPsqjLFhdAX2tBaKm9R0CMmLKF/sbr
lcXAOlccE3ucrmiZXW98bGre6/oAkmB6E7HlGborNxgTnhVbQ1EyKXcJDQiHgxOof8TEFQuDZtH6
yQXc+3v9er3Y2fgkjL7mdN5Rigiq6Ct9GEwLnjBl/AqHTAHIzNoyoYG6MkoUdO4BMhYcL4g84VZd
ILAoUdjvasz3d9om5e8NbWb5V+3feSWmsUZNyfuUlcHMVLyCRwkP/3g5FNVPIBS5dZo+a5wCjLu1
6v3BKON3UhMWk+qjkRwoAdUhK5088dGWaLRe3LmpoW8Iuvf5vJaLHzKqMFeV1E0ZgjGoREVipBtr
ZdZXj8SqPJ5LnzRbzWvigXVn122igYhHa3n93bLmHaMXjPSXQiM52iNLTPjssmbasE9QUg4SVxl0
U4LQwHO4TUVnWZmvEE0KDR8xCGt2u1N1iOg7vEBcXa+P4VGA5dB01d4Zg9EoQMIybNki116Flz1R
2a5npT08Ndcr0/MLi+MmVkfg+N3eMYTtgOyn7Ca9EqWM9kpixwkgaCO6Ot5dhzbm+ikncp118XdG
rDMmqVDLFKFtx4pJlD77sqEuwBh4qQkKzKEMHn4zIldaXs7VZYeo8sXmPcrbNaEDWBeFCZEnoGLM
ozAvYT9eh858zpB3+hcL0ZkaCoLbDFy4bRJMoL0dmrusons/i7SBRY4t/kMlFiL58nfY86nZL6nr
fkwbITMy3QVqhVVkudxGkAuWecchvSv7Co4kLpRoiJ2gFMbmT9sj1b2emdwIWXTtbU4NQ42ML1hi
CSfcU3A43XRgyzZ1ywzUe90d7ke6kOt/ksel9RptqGRtpDwrQIroYsM95rDcKpo0AYY+JnDsxcAM
cezBJ2kMLgz0kPeM2e5t0bn3t/sxC8RxMaJUGD+mv7pon+ii14omUul3IpY9TFlFvjShfYioqABO
pCdfgO4Bh6GYrOmXxdDGDYSp5Rt9lJTqIOw2gpGgpu6IrqfxnztI1zGrNihUHfp91CrKoO+07pfG
qKmIPE7cX286vPRte+MNJrqmiWO0J3SIjGBcp3A0gy3HKpqFmsKoApipiCRwD+grGzdIR3unOMxL
mhKA/Ry1kGVK8ctYXKM4RQG3xftSvKklAN46KoTm4igZo80avqRBi19Gtxgx+TgzCfERUk2HCYhm
6tH05hK57rRrpQRva1RUOyhEI43wdRGUqXnfL+lELQOiK27g5Yf2et5xoCBR6QJRCAVeyw+7pnny
CL6OfNZ0vbS92YK2XqrrpN5VEkL8dwVPGSeSP8v4tZOAIOM970+eTvwQ4shulDiKSISGf8yjL/9k
OXypaC03TFizNxMc/rxge5NowI0Z8QnT1oZEVgVr97eRRrO7771vxnpTpTOtTe1tI6z+DziR5AJY
EZyo/KRG/NXY3JvXsWGU41FBcDV+wjlpHRRRlX5PsGCdI46Xa2fwtfzJNJadssQbRmr9WTQaokDX
HB0z7r7uQwjllipsFyD/xBb0fes9fVf5PgyHKiprah7mYWQp3NloOuL3lgXKHdCjZe0vc84GJaDG
RebZ8m4MogzLhvxDkRnHc4BlKHScfoziAhZjT3uUt9x76vSyPY/bC4npyVsmx7vY6KBX9LRJhuuT
R4ZB1UarwAv57h/pM1OLOgmIwOB8f+TrpYB3tx1+uSN5RQxNOehLQrGfmkHdy/E2N7+JL9CG40Sr
jFmOvXmidY6WsgUshxHyH47Q45ZNZz/K1HTT5Zo+3SxUqsPW70aVrWFYOZR2x0YTt2Hkyx2UQMVG
4Wy/R+aBB2tICzCfC1Z42K5sVs/XUo29BngSgqYVudwk43vRxPzcRzwHRHadn4T6tRLs4C9D6xAT
Y18JJ6zJp3+7vZEvCJEABBR00nsWCc1SjVbatMgWgxpYD5xeqOPZcFpRnZsRaSmThtqx3bU6eII3
+4AhkWZYZ4kJdIhQEDeDQHTH6XCx19HMp7MMpqNdIA1fH/Au1An3QmWKuD6Xs5+zAlmDY3yHnSej
6KtyjB+I/Kfs2TmOIk+sUohjiqtESiD2jleloRnhrIfUgjsnanuoSu4rzts9caOe8++nXzQT5x8l
NMxllpzQxGl2onfy4r9hTw8a5k69RSo2xFWHFuleQ/nQnDWex12w1cACIL00y+YnqyL5b6WHZ45d
Tb9ihryRm/vfh8c3SUj8FzWSnVCClO7artKHjGK6ZultmVHGg8g1FuXlcIRS/+FkCbDimurGpeYE
S6dONJ1x+uuPURLHj3fLZS5+P5DE+7gEsSOcTkbYCMCDDpUDBVkl14t853djAsPHKZG/DqklB0O8
g8mh84TjnBdy9SKkswvSikqAjT6IefnD5Z8UvJCrLrvJZeNhCFfIeTb694k41Q8xVCfsc0VqfhSD
P1+YssEBWLSNUm4H+h6RYrrXi3f4T+oxJuNrJrLAsMdSU25y8ohsJsgG/ZwA++zyFZyujoB9F7Xu
55xpWX3eu67z1Ru4zCCZf7o/5tV5G1aMiFEJQsAb9dXF8lxpzCK+/Mhj02r5iB/FyrPbYt0mh6BK
EMk3wEN6Z+1Baxoki9aZAsutSVVDA+/3K3pLeIQbonsPiEZ2MS0WE1EMG8p5acvjHLg5z+rcZqMP
SpFxZgjeDE1mn3DtTCzseoqpSBQmvzDnuIdGr8cFjkdB25LcboC0Or3lakPFTLeBq9GzXCG+XGR6
eSwXCxcx3jmW9mr74XwzFVWEFJHUfyqBPpcZeA/mcmOh4LyEGNecL59PQLOo1BAdpQTSPMtcg2xi
rbGFUrh2lcuOHYBGRVfqs4eVtAg0NLiAtQK9ZFWbByTQ3/w/TYtol23fH5VGiVLxdjEWMjwFPFZO
gfSLixM+u1WWfShjEg8ZDhM1T7hudvLvJ31vgw75PfAehoDSk1ezzUiqC2tniUhsGooNRF+/nS9x
AB/at93U2axXqbAlcUIfyGPLaWOy74tKXd0GfFjX+wjAkP7MBODV6uHJdkd7c4voJAeow5d0nUP2
ujlvW2YmlgFDtAbnEJpAGCAqpNf33ZDMMuQrat9UqYUf5dG097JHAHyo7rsU4rRKzfsuhiAR7tsy
uAhMlH19kIz0XZcf/B+WYaV8BMMUnmpdNiF4DGckSi+XSY+8ljUMp4IxkukA+9hXAwte0OfwL6t6
em0WpPzc4Psc8jjNuGMOkJaB9g9Wtm+Fn4LeyaGwiktdXxUJ6TR4JPGADD+HJzSnq/DSMji8Pytz
BnwXSvA20AaIdYBFLzc4TonIfcx1iYbI2Oc3BUmhDpDQTBhUDYnpCst4AvDDlaXMk0K0CPABn6zk
uoWwDFkfrN/qi/QQWUcSH3GHCvu/jP4S19fauxIVv0MDzKS5dFayO996mWhOGPuoMkh7xaBvCaYT
QyXH2PsTAyjAK1qaVSOkte/Dq7ynAU8qu4T5nX8U3xw+Qic6S5r8QMRrEWSaZ3HEoYYB7Rw5Iult
C8Aq38L/RPxj4Loydv8PBG4McVMbRRXXp5X3mGcSvdbXsnFs40PLt63dzof7Y+TNNkolWLbaBYHP
hRuVzV8X01HsjKVAj6YmMpp/kmIvgy2oxWVHu1IiB8/dqgBBgPPCr891WbXGHrhHM2hk0okOCI+M
USc/nYRfFQK/FqFNOo7+F/KlYTdRr5/fHb/d+BbB0hstinU1EjH0VGhI6M4WaUhVR5ayvzX5a1V6
W1MUdlDbMj7x8zxzMwFJvhcBtM/WM3Yq4laEzKth/42agCHlYkFmOszokZqR0eqhn9qAmqMfJgA7
KWcBCBWU1eAyMHZakqCZ/iebWEP5hGiUg2FdcoLrJeC2y62cwzFrxPA16Dt2iEnHN6ued3Y5B79Z
uZZPL4BSOQAH3iwwz/vYe2sd32bxz7eWDV+ZLsrcM1FlG8FT4H0nFK0Alr0psnn6NhepKV9gkBEz
Uc039y2ghdRWaQ2nP0UzdYz41f5VGT/I2zMoOGZ+HfKSpb5ZNEzoBixYJPDIpOpNuCoV8O94BoYf
IbRABkvWtEZ/F+rJXxDDno6ZtOuS35i7Gs2RECvj31TTBCSWct2GmgbHRc4VGyedN8sX8RWE1Xyb
9IUPYS6IjrOP/f3wb8tsiwZp5BAhtsiFh0Vh3bZ/Yjm++WKgw0a9BJd5H28YBJq7WTPIWeGLsNMX
LxLHDlLiUW9+ShbBMjDHBTEGj/HupfNOMnyZeSvGa2er5VVrZXcB3F2b/dOhJo+PdRv4zR+7nPAE
SQRaXD9K/aCbWZm/ANkoS2MeEeM0xHAWte4NWrsVGPy5PK6gmsMWpwoDyQ0nXN/26tXNL/EpYlXB
KvSLWIS6m1gFGr3cUMFt+oED90PZC1VodTMm+smZoywAxLrX6x2H2SjjOl94sMCRpiNnhtnBlRgw
1XgdmzhjG/bprDcCPx62fjy0FOnrFIJ57STJV4X6AjSCMe8Iwe1pD5XKFcOiW8uyAx1Mb1wTdVjc
hf/obfUpqVNewJ2rKZRHvE467y/3eABvGc9Y9lav5TbTknR1tZUd4jlAWzX/svuvegRkY90i0BOf
CRdkgMqeD7GqkzcimS4pyHCI/7tJSqskyFwzj/tw4GQ5IbiH9nWYQxuj4CXsigbTCXlSwlVph17k
TjgjVh73a+hC5xN+48xTv4yuf2C7awLydlmeMXFjtiCLS35dcewQKwJzo+LqTn5FTIdW3e7j33cD
bZuMKpucagUK/Of9Pb2Mpg9Bo03mdkXiO2zpKei/631VKVsjQVeGFw0b+tl8akUWqf+L3pzMEk/J
ylJx+JExevEMm1rWpbK52oHO3VoYfuFTt9bqEbxu9F1g035xCg+RzS0rnpeBaGVpBKkYzoH/uafD
P1v6Wp/k96C1v2qInW0M39ZyQu5beSDlPeCLNLdiY6xFNyuFKpAAXckcpl0F5jLrblX93t26ZUCu
uQBrwzfiui5nIn1DxSkk8qN7uxvebJax0/mESZMUxNJQi6RRWyO8VF5n9fGO2ieEIPGrkdZIY/1b
FvlUjiIGDD5xhqp8OlVN5OAx7K0pClOl/SmsUepAEQFSmTj2dsSUm8SpcEqY3Tag5/bS6synpZM9
u2AkygcoALEMjHmq4uCb5vqPan8iXML75TDKPeRuxygZGC8q/ryQs5yZSuX4stfwdgOgQ+4UNomn
6uiDojMpdmkXJG0yLwbo6ECqDbFfi7lipK72Mb3Bun/dFTI7j9J8pM/Z/9a96nzhKp6OP6Njv/RI
YNlbwKSp2lul9jt+grPSgm9iG3KAGKcd4yosy1ugUrJJtG2ecMj4GyZFAb1bHtr/nDyyZRbGQkQT
XLIUDZjZ7ImGbMWAWvou6Q7LRzwYrSlfFmUCzHfnr8yvB5zErcomTrubRZPnpuLyTEqqQLfNl8pn
SytrdEm/3iyjNJNcNarR58DGKVCj+cT53/M6tJ2GZt8p872dw+caZfpn2PEYtA5azy/A62t6aur0
56BV4+iBXjtmSyju2MYSEG7wHWhNDxMXle4XXdKGIILepHEa6MImsxv0UQq9mFfwJEqGzVvqukMN
nZFbmF3PNzpemex4xvUiBxz5vTEZVeFPaSFZ+94H1APYRKkOB/SN1djQ0iw6x6BFKsbF88+9eq3O
BctWLS7s+lf/cZtT3WjxC+b5iQoGvpr5WRiM2dEQIxGM7xl1I7Nm+x1Uj5HYxaM1PkWVNIo41cvv
Eo8EcLBvRilc66taoiNeo7YwdXmj20l4LZY8P5fMsx/w1w8zedyuMUBEIVDhHRKVjh8B0xL8N77l
AUwTUkUsX8/ZA2i5McsBPF5G/ZnY8kD8XwjCGwIeWuddQt9yUyOEyN6MZnV1fDPgJhWL+8NWV8cC
XHzVXoQfTBOB9qaCLKt1ifoeTymj99iCblTCkzNwMpPcbyHlmWS5JNhg9ezHyzb8hlIgCLFaAV2t
J3HzSmKSiAe0XnysNQtION48nyDUGTNUJbPzJA8V+RozdNRsxkGbxQKQI0Mv5noA0p0iome8pvJb
QaMc1ehzSuV0MwyLg/fZvBG5H+IVxY2zPXmLDN4ariyWFdwhUmnyyY7b9HUVeManV0DBi2kRUvqb
S6CUNxHzXFXqU3hWFAvfptGaGGLGXmrKlhujv/MORriNKEtQYZdBYQ9AXUELdIk6+QWkZrYulL5a
3wAJ3uwYdWaQ0VfiXxyJqd3r5V+iMArO7+SFh8a/cqXNj36ONG5HhC8wxi/UlSvVD+b3X66xQx0z
uxtDuD5/qSPvJ09YOwwnHP1tJ5Aslip0XsGSktWD3osAx6EVWg6TZFuB9IS3T9mLVOu+1CW+FpR8
ry4uVOmj1B2hfP9BHOsfZK4CaHN892swA0+5ULJTnPNggduG2w1gt/3umPkc6gAQ6vpArTUm4DJy
D1aYhzFGH0yJWUYwwEK7DP8m1M3gHJ0QmAYCEJRnSiqYIqBwZlHDT1X0XM2agUaDYNNp622BR+ne
Oq1nyBx7R79NMCmAnOzig3xoqoIxHg627bgtZ1tbJ1q1qq1I94yGQUICA3NLrtFZSaQEy9a+W5IP
9GDewBmxlXQxSWytPELbjP8LjQdKswzW/w74L86CN5bFbuwTrvzc6XcQV1i1vSkWGLJ9IS0N+Egq
1f7c/URNrjjk/9w0Mw+Qy+lLKsEkFGBGwsFWE7+Ka88BZzv2f6cbYjeNXpnXYB4SDbnVbfBPJnr4
e+o/qU6BHlHwEKghYI2c8aDiuINbcWdWZw==
`protect end_protected
