`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
PGRRSgf06dCHp1JlPLtIX9Q2swIFF5gAt78gddFbuXC/t0ROFuoAucmNbGIyTgIpB3IxX0DNsC1H
77UqznaJ/JKOHgzwjNaMzhFGIJQe5LTx8JXti9X8IncAa26B6latDDn83rWmX/QvSc485VOXptzZ
3btVVSS0tbCQ7l9AmRF5s1foesKFUj0GeIyoStn/YJbi9cQrpkPb+RtyqAkyYeBZCTojCmC7cA7e
W/jDTyY7mZpwxo3975r8O8gOP+uyRI6nXbBlx+N7xMroizLL5U533nDDzqSD2pDv3ptXYsV8f5+Q
7h2ChXbfwkj1y9rCVdTz00y0nWhTNKD3/nDZhg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="gHGq/Gdek4X7kG+9JW3CbyBeQY9BeWUQZ91UUTmpAP8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9984)
`protect data_block
wvQK+c7O158c35iaJIHhMRNI9tJDVNYjx0RtWRt5+ClgTcbPe+GT9Vdp+nmC8A5cjOR0kB/ryqtp
l72t0EB6uvIdvgLANIN29p5DKRIIzhxpqoOuH04uvto25v45Atzh10D/UGbzE0sIoa7vPk7XzB5O
Bpy4ZVVxY5vB4sPf7rGxWdbZpj0MBSwfles7FajvWs0YrpoV8xmbRMveGlHy0cS8j3mAOpTvODd0
85d4L4QntnGdpYWjimQv5gqmtGwk/6pI5FGE9eJ/wCBhNzpItQ5HijdhcNXct6KUuHCGwHZOdTQp
tFOhV3YpvY+wk0phTbi/kH7CReTA7NlGnHhqSg5PNosA5Hen8UuBdIDLr+v6jD/VegV2Sz4y9htS
iyHVaYLPq1m5I825cKzi8h1+GrnuSXqlxDELcBqIRm4CVK/19o32qSXLcM5gdelb4UHQHRgrkd0/
q5b6GpOlG6oou5VypmOGUAzTHrZ6xdeBWbf85jPSr2LA9z/M/jqNq7sR0NVwCQzi9sQBItkS2Rpm
neRQfsEEDAAbaFqiLsCkmSEoqlnnNeW6tVJ1R9cz1q6oX3q8NJMOiUyIvFAfCA6RdaDzIioZSvhf
sLjmwXBKLqb7RJNnwR7Up+PHuRtXt+Caf6NULLfF1OCjqrQYJuIppZcgyQ9xbVg5V3SZJ4wzrl/Q
XRqq8qlk0YSOGgKZwxdCchvoMKGWD4ozSC5WCdK0DvRPsG3Q6iErlz/WW5Fw5f0uT1ravpkAAFei
b1qUKFYtI2hrweDOdY4guEmZxkqBGxrScJnM5TVh1Wmwjowxwa3xZk64eXdVHAF+3d0JxW/63KiC
hyOoGtQv9H8cj2pUB6Em6SxiB/WalB6IHnq+wAWjwkt+ZIR3zH8m0hUk0ueYKa5/eyHL3nha+HOh
FbAlUNgbuuYftoXQu+QlBlWcSUwAZ2YMUGJlyIQIbH2GEUwlHo5/lITnG/B2YE0tMsZObj2VLp7p
lls4FgYqHQS9shPIFZD+lKdaBsi2Xu88xNw1EJM9v9ffyJcA6HTdmIPWt6Dn7glBDKLIIfKYlNaX
lhnWqYTh+nRX2YqYtHefY4NuosYvRu0BGu7eo7mdQKxWDb+CSaAE6kYZJCboq6gQXjYZEwYoVFew
5KnBwy8AeT1uSxzMUh4riamqOKc3MK0vWKmln8Qta5M0YxIQQFO0Lh3HyPITIM0aRcDGFk80HxEX
4UlYZ3nx/w4qG+fbU9jf5yh10/twIVZKyf8RxlMuzBtWukze6CBOEnyljrLo4N1xxA8Ar3pZSk79
VvPHMkHF90u6kmtHzTdjNmARnBLvqycUSx4DX9MiZxzPhTyFDuEKH7KHxoB85wCA9eDr0u7yQOzl
N+On3T2yvrnd15GhpV1s89iI5kt5PZh5VB0mg20S36RMq/t8G4yz0ddQ8T+o5QSG3L2I+JEnyXAJ
SRnHhBF/EanXqYyzuBtKIMx2L1jL2kMSSN59VYJHUnjRdJzUFXhAvwOg+D38JZ4O1koXlms2m4/g
hfpSAaYwswJPq8/2RazLB+RKrpkfbV4EhNNuae9UNng0kO99jQCjlihRA1ybF3PstxlrLafPoTYk
iQ/UBNaPQhE73LCTgdqWBDFA5tzkpE7+JWPOMTG/AFOAco4zaJW7QVTlhMR5Yq/2KApb8AKsa8Bi
QNDy40W0tX/ASiLpsCawAVWaO6nPdEZ8bd/5nq6hgLAzBuTiuIDjELvE5AzFNFy12A6xJaIU8sRD
tWJrCf7lu4MwM+DkMJGMVVABdVnDY3eSnSy/mREMNmM6Fk8KU1HxRRWlM8G8Yfp2/euDCf0xk47l
nqh5adQLqzPSNNgCMwL+rGT28rHQB8JPcnpYPgdoGIZP4DkuDYjawxE+SSROdz4gmscDYKFKIZq4
zbOsSCtIbwMCIWtQ8tvlOewW4mZjcFKAD/VGU48Ger5fUg1nAr76+UerZqMS/xRHmzrOb7K8bz2L
zaWj0pxNyQ4ZTSjhVQOBkcnJRvtlZ4YLoxbUK4Qq2WrKAN412FLRYrrBROyOAvseTu5fzUdbjQwk
yKiEhzve/htPRfsuIO/bUJWWSXIeKxPrkSmesx4dXvEjVHNSPpDwwrsywcndRia0m8X7BkSi2Kgq
4GTc+6CrD8B7lAVBMYMjexWQVxDMu4yHtqHP8gYmE+f5c4o28yiNuZUQ75O20YUXJ2uDhatMTd2B
XuLo4c8R6e/zvb0tPmxwXXpsXV9RxL3b1neE4W6m231gFgnx/2ZJGfrJlhd8WGpjVjJGGRTjc8qb
5zYipAtEITPb5++Ar1sHPOGoE1aOdNLKpbyp3lnKoUPjlKlOW0foT0baZTy+4yEJ1ImzexanZAum
unQEc8Mf0GBionSehbyfJ9Sh3EPrAXEK1dSieJQ0UxJE10QzsBx4wwud/Ovn8e4pRUODQYKWASsr
R8PmCYZuuOqdyZ4qQ9WtTNO+x7rKSE+DsylrdY7ThYW1mH+vxpUWSHHM22Tt0xA3/uHY6eJfn0d/
ehTViExaYF0efxqYpI5032Y0yrR9zAJQjVGQQlKYRPzEgx3PjzXzyW3Aqt2kIaOVj3FPZEhIp+Xn
8/9SCIwUpXCEX0iGHhDYXUCiunuqojyMyjL568JuBDC5r7gpG8zv7qlBHWSj74lWqNAqjWY9lzH4
kWk8G0K0USNkm7hzpeVPd+5Aoy5rM66X82emcRwUacbkfAEoc+mOWkjqZYb7TLnv0n2cmcxXj3Y7
yqAbP7KjaiEh9URG/PEwu4usZPXQZ2tDeNSqDrW2LNvIMxoDXC3OWElfXuyaWChMvKUJhPbytSaS
owJEAcV3Vsd6qNMYlnMKRwZpZVgOCMqBDXrCN3MtgOi9M267u4b+rTJyrl/lGvf9waLWhNo1hBAI
fbVr5WZX+EjalKrjX4tcmEllDUAPkArUG45uvq2iAiriTPCG7dbVheysYKG0bzUFI48EUovvtqKq
+mgYfSwtdOjSPqM09b4nHt/Ht7aGBDeASaB/KIQRBJuOtOxGFqZ7hIRVFBvlEueteDzqKk0dk58k
bXhBJ0giwRyFRp5qVymUCCF2YdvluI5kyzlppEeHb4SoTOzdG69bEp382VdvnqtitsrNoLyURHgY
Za09UJRp1Rnm639DszeQTryfRwALrzMz52e2XctjMfvlgWIoNv4/Y2+mLn3gi6kMiASFsV07IQe+
u/tW4foBbvBrRZnXiQaqtaPGx1Vv/jyVaic1YxZysoZ4wknnQJaNv+PIHoMckMk9rcvcwnr/gSkG
7kfxhsl2+rrLFlJDo2X0afc6MOHp5oPsodo2oHNyke8Z33zwYzC7uidG6//BNxHiC837FJ+7vkBn
dPcFfAeH3MXyRMKRrnNctr1XfuLJASmKL4V+f6BhBDrUzNeZcvglZ8GmxdyP1G52uvWqnG7oigVf
UOh4jtgrASf394Z1m/e3zxbuOJxR+Rk1MspkPjDFOEdVz8cgI1D8QsPW1RWqKKg441F/2Q6qTGRV
kRAj8bDWusbkdhJ9R6jW8J2dbZXDuBH2BT/cVScsri7erAzxp6zz8IzkQ1f2ObOcObbbJiOBpqNA
ZczKbn0PXUAWtyk4xwEU6zZu7kMv7dY+lA0gE4dm13Z/3Un5ohFyv5/NpnNMqrJAuiZq6hORjWib
5rTvkkZWZ0KLQZpxq1wHfn2aMh5jgtL1QzpyYszkujK4GgSjIVywq+Ur86XTlbNQPUoCO3XMj+9Y
Wo6weYJtWw9Cpt3qH31Bz8KR4LhxZpu9DaGhHKQeV2Es4jeitQ0Id6kAy8xOXxRpz+wKDLLRcs0t
TjST9higeYkjm66rm2X5hjnBAK1FMveMjaMqffhRW6hBFqID4pSyRJQbIt0HaYO2ZpayRE9ZiIn8
O4ni4S++UtDZs079ZcJwOEEjV0v62b/7kMz+9tTN1Z2pGXV8OmBNTy6qoYLQXJKk78SQsSlXYhyA
kTjRXqKnflrqGGx5glLVUKAPCM/naMXgdagTUhiAMaQNcPwYMbTR/ymavJcPsWwsdUX0u7y/UYJn
yf2RzdLRBfUV1Y7M23tnRRLGQtnMRdBJIBmK3HBXye8izol7i8HC0KJoxjVxkBnlPJ2Fqzweyun4
AMkaAv7t2Nmu1BbYyPJAT3ml452JaEFkabKPmFJWLKsdwHMOILQ9bi/y4ptCYPn1/GoTR/mN9Cq+
ProqJKzw+Jqmp8f626FOp/LDP2fzYZVJ8SS54geUt7k2+c+07LKX/6Qw1DplmTeknEgsAYjWX53j
SFB8YsfC4vsU/iLmt5V/GO+ylgbiWGMMENmYOGMy1IfZs+fcXi4elZttS/caB9P59WuuqcVTemvA
sV2LvC2/1BjHnTx2d2Do822L7KKGiIDAY7uP6GydgL8btbmVen7LTtbCCtm3KVjQxHbt7X8AMlNO
2wsz9eBROL1N6Y7D1IAZlMObOlfOJFo5IVy9eYi1EkYScKgLMf6kDlCUb1pc6FiAr96ulteq40hF
24WAJmcmCMhNdG+UTeDhtZSfCzioGvHxxVsnZKz006E51hIvb4JLru2H+yXYUdLRS4rOTLNuzXSK
v63SRm/ddRSXZDD03PFVb/Hur3heSnWmMrDLUT318JdBuvG2KnA6P0StBHbdSUGDwSY3fMOfK/X8
o7Kakq2LazgORFFt1xUwImOBeFZa7gW9yfVJl/AKGTjE/jLFyYcRirAaQ9gwCBJ15zxaaE6j/VRf
TqH3Y3vljvI158sMjTcWrNOwrCsliC0KyKChhvYacvKmP1gMfEYfJGWP9FYtSs4iFkRSlI9lHv4E
jddLyja9LjKIFe8EJqQVvAKsuf3bCxi4vejYnX9K1UKVT7VSx5W4kjtmRHuvlbxl/UcM6i0W4D3y
n0bJdON87niaqe5XNBsDIo+wzoAsDCao/3BHu0O8It3kcc/PRutIF16fMg+P6I9rxME5+whIa3ZK
6DVvOr1HlSTewCUwTdb1ZiHHgL1x4/gz3FqGu8+qNVoFNeDxmil/KUc2YaDWtEa63p6zOc7mtuja
UkT3Wtka4JtUVKxwLlB229obSyRBLhWsGNQvro9mQYARgq2Pg3589KKIfm17z5Va47wknbF95KcK
QZL1HtiMAk1XEwYTYzXSws3C2byVnTPcwbt/DcT2vCu51i8ZDAqq4vzkl4tcKqcntw3Fag/nQu//
gf0UxTy/eQf89aji33Y28DXYC1wbAqbQTIMmNlP+gTgRhiED5Qs3ZyRKTT5keKyatWqddVAsK3l+
NZaYuT7fAILch5pKDUPBI48d/bgqDXmfRnojtGa//xyUMXk1uau7wFTy3nQ33uCYmRKxC6rzPhtl
ZTJyxJ+1IBwPVND/ySzPxXGO8gy4J2rdGufQCc304Y0ZJOPkB0xSpKhYEo+xc/nZozXXXRXEWGE1
mr6LFsKCuXPOk1czEgUHefrv1na90VoF1948LcgZGHKWcNwylVwvWelS9SkAn8UNTdpsOFmfruK/
QMBsEzz7qHiVs4H6r8qKbOBl0fzKvtLROkyGpKLadgq169qbriGwhnIt+ZExVO9+6SdGrxZLTyL1
hwLlXeLH83pYYQcUJiWsRm4oN2/oUw7RB0XjbKC1jFmgqFJ5Pf6VbSti06mlAjxVVlUNZpzsAEQZ
Ch5jucWPI7Zc2gYXjX+KfC/yAggYALJwITgpgtmSDOkSvrDEAj7O6cHVulMR3EZZ2jh8Row1+v0R
JIq/mlTJ7C4eKzsq+foojUKJpCj0BlSSdx2LVOlJNC/Tdp9K7zmOXiJOdfKHWxnmJZ2Be4aGxsY3
jUZAg9I4t7uGyq1rxlPbKb77LaAr+obqTnn+iFqC3wNjZG+Z5Y3fJUuepkMg6pL/MhYCSX3DWD3f
ABkUy74sPj3sAAyhBel2hFnMBWDjPJ8vcpD0ENibsUIeWhNmyofo5xVkzPTj6MHiLVn1wRtTY2jK
Z1b1+qVyoUfeaA3ijjd6rc0RKiTzOEAR8rAwtINq32ceVkGysqM2Asg3SMrexUycOXaxZQSMuAF9
QtExSflXxqx2eI5k532pa71judBc19L2HtjeoTtAEpA19oCs+7eCcBv4zEo/H5jqgSG/iFqUclcx
yluDT8xFfsjd1fPwjGl2rovOMEDOfiwjLlHJiP737jv36FamAEtUs7GbhNuin/jjso3y4iQp+iLB
M9S+xOStQ8HjJi3ERI1fZi0yBMn0XpNuwKuuU3JQrwvyYwfYyCqUKIro4jfDnuoZNMY0yFUiNJX/
QHaObryhgfrr7GtThmW6LGKr0FArLFch2r+jG5tJ3EymJjjj0+JyWN7KEGPBL7oLMfym6hK2MGyO
BS8S946XFRglF/ercu0BY5Yx4wX6bZPDUQT9Z/GxGyHjy9P3kTxC9w+40llrB8Li33ZHWYxorrZd
mORODOZoW+6xFcdaWff74Nj53RTYCzGEy1evT27Jw2kLoCXhTce9MZidyM9Z4GMSYAeq8Z34NrDy
QUcmXQjmlOUiVYE15jUBj0wyLddUs8QIkBzPT+Sndqiv4p7doRCLGIggQjREI2p8Gbn0iCRM5I3z
JNmBojWl2qOUHNOOHjw8AaVacij+7iEKM7rmMlj6Zg1SKYyjIIqcEyVF8ftr4l2bemwCsZAUEEzh
7TfTTOsGlk9zJNolsnlwX+wPRsB0ZxN+7SCBUbBc5O38CxK5u71Lvgqw+dLKwrh2XrtR2Sf+1xIs
tFnAJ6szImxKiiUSpiTYL+k+pXP0mv8XVghSxxNoDRTM/SYgm10dHVN00TBuLW3ZrhBtmc+L/heS
2AAJrstb6dUZqLUJDwhrIGNUn3/1tzZDTTR37KFOP5cubvbdSHDVOBre/FOy6DgxFW5anEc4Zb0P
om/Nh1xpBUPccaMnbTtrvHSex9+X2vqgQ+Tn2B/I9cn/SVGDgO/NSjpW91gjX8dGMKMmE2CqPNir
+caDjK2H2wwRzcQCmjfq17cKAjs5TEELG2df9BeXrRTyAL3tNZa4cnKvtCxsr+JwcztjzlHZ5zLC
RWCvaQNEeHWr0/1cWbm3osYgJ6sF/t2pf3WLpVgHoVzNyAJtsi4qfMWkNeG27PA7YmQLZqHuNcOj
/wpzS+aINvjHXjHldOZz2IweUoLBCcsM4TZG/sKTuu+FRo0zpDSLzVhe1VcTQO+cXMu3yQwmzUZ2
DPfYnbfLH2lnWtVQ1TRPVwHCz1OX49RB6mHRwTJ4W1pFKvED7Jr6C75i0ELu3/q9a+3nEbgejDoL
7YcFgnlojSnh2/1rCJjYWJINBu8SvBt/JXHAQYEptEar0MbaSCmZGTxbysPGa6vioyORZQVQyD7M
KxH7ZWySmwi3VmBSAI/zbd5fCN/IUH/ckHhTW/SZTJnJ1ErU3KVm7nKPnBUqDG7w2919Scg5KbYn
LHzA1wFJDLdd8bmeds6BmzS1foihKKm1vaqAEL+nGDX11xKQCDQhWrOiKta0cBOmapiv284QxTUC
gvFW84kvZXArGolpjf3OpdcjJSeQE82ReoiuzFmU1y4oKUyODCHlrLa+2Nt/TfO4C3JUQW7EKMxg
qqIy1wG5UEfOk3Y0N3KgsaRzaiiQkLDvUr5CmELhDfO1RnJbmjeSZPJXiaj+0vBghff/wuL7HUUl
dODLacZhEY0RADxVVVcOpS66++z6ZShnXZgXoOcRYWD+rnhkbzRQOvOy86Xof56btUy1DeTxOosO
CDUHVCdETxBlvFo8tWgdXDxeT8JOuSHsDOL706QDNvinrhllxTdsFGx1vGbzDbo+rqWgXZ/zIPFf
JoAiS9+e5uTPSSa6vtrzWqlAiVVLEBI5k/y1qQgOuUVWT7mmzGZtitDRFCNzVd8ZGi+Y1oOIoSnn
85a6vEGQt8mwBU0WdS6MZEdhNvMnorRYVbTyqcY2lHTJnz3hhWbB5pfrICm/0yzbIa+Krr/aV6ms
9bVVOtBglNTMdxdyGtlg0efEJF2JYi1o2HNVj0lQs2ylvNgJviWqqANdobJvSnXSdrBifklI/bUD
tEdEEmNsVHWH4bn8HvOHW53myCGKWS1yS3dw7h+ft+F1eEgCRuJ1VE8JV6tIVP1AJmrcqGTfz0hc
LTLUuKma1r0vCwDuoaj1otA8IrMSsyz3jz6T40bToB91CBBKY9AS9jF1KwWnnjHw5qLSzViLdPRK
QOOzhYmF0f9ThZQz691Z0IOnKa19GUr7xOkPO785jQxBnjPqh+Y+lY9fnwP1bg61AAq0lpZfvl5Q
EPC4ixvbndh+lOjyWuvwWJgxf9zlqWiSypUjnOPdmn8EjuoZ1d5nGhNUyPNZfcl2Os2+o3VZrafm
6+3onukq5bH7AcIi5w+HiX4FHwfps2rZowoTAzAk1z2S8nph6ML1QJx1O7AnUL+VNerKMTe/xtPr
5A9aLJ9brKePEHl/wwTELXvYo7zPjHIKVrrq4Cj3cifEB83ejeq52TY7ewviq5UzeVhPiZ9Tn/ky
z5fxVFFySV8/sZSc/KjH6lb9am20gXcwnaeKFp8Ynmf91Z7jTzk1mzWc2ZbS7Iijb4acDtTz9+Tc
gNe/ZaP7sunfhoEv+fued/YQVVFVrUz9m8h5Aa2ixhXAGGhItgGFhHEWfbs9rYYo7L4jTJYStZql
erlm22jWzRHx9uvbki8uW81OgSylhMnTv1XslosduRY7kieZ+vAaClOGQ84gF2c1X6bS6N7dAuk0
QiPKeWDH0s3AcCSue7khJN6Vw7G/NlcBh+DA1L5UZba3ugXh2av0ImFbV5lw9fnBRQpFfasNPTXE
wMC+1GiT659hoBEwExd0SN2+1EP8F53VaZ0u4pNYE1tTUW2si6E4rEuP1bUVBRYiOu4StHIrznoY
JETIXdtPhXvXulrLwRSPMi6Q70TML70OTbpcfjzr5ue3M01FKsF0XwbWjPf8mEoXA+R/nFQq91JZ
ziqsPPVYl3cpFvkMsr1TsZEr8+VROOq4j6Md4zuhX4bL5rCp7FOQscmHHmiLoqLRxxQ/fC6SXItu
m0mr+72xuhdEOKIGl+ira4IGQ4t2H67DYklucE4isvixiNg4NM0PRFMXC9+gHANy5vIeDzGMUz9O
IXHirzbHL2FMyvQ0nJ7jRusTOj2M1otRZZGzFVlBmQtZve7nrYDC/j4Ynosk+SsB45rWqe0ttWzA
U00a1gEQ8z/OpgTb10eYatk9DmbFuYPt/ygx+Z5sotNlTn7FU3kIE5+XJcjz3Dvmn9/23WG2w2kY
z6/FK8UrRvc8RphGpTbOGpoQB3XF07CJwv0ouOzhMQktfFB8FaHZAtddWbcm/kmYIEIcIbT7e6FH
I7gHUXzB6v1DPKLONVD2fQwkiAEeHXH6MPWSz4BOSIJaIpkepRFoAc3qtjs6mMGIOhZcKY1ShiLk
InqG5PghQ2Dp8pGaR8aqYT93QxUnnKpg6FCony+c47Ek/xZCdCfQYZSIW6IpTgeHaozzoaDAVpuq
HhbyRsL3GmhoydfLHZ/i/Yxfkpn1VL4G/vL6ENCH2QLZQXiaEI/IuecLfdvoC5uTySRfehiwthHX
N+uD8+wPypoxViEvUaxGL7EDRgVNI3znPazkQyFtrn8ArES5QgiWyymz+6Yyga8SaTGSvrayv17B
RpZx7cZXc/7M+A4NxQlj/SMTSC1lZxmBZevsaYClA86uRjoFVwRf7HB1Ab9OLOHjulbKT1ml9icS
BMXrRPdM12kZOV0OQxXYIJXyXvQv6F49gi5frawxIy7sH3hYJ8OO1XZ5zCDRa5I36r0xPFBnrZKZ
/pwGN98EjEnXGj0eP/q2sbAnvsRpE+PS99bKgN9Z+PYoDY+l3+NJ4p4qznXcKZu54zfh3jkLOqGg
/cVYm0Jmk2ztRxB2pjYag1ILb2eaRJiYsYFfWRVyX13jahABVP3YzzRzhwPxlSG/BKeDfi5bTbTs
aLW/wt9hxuvNSU8gPzQfx7K9j9fwrPGGKRrC3NmEc7LS/KailAQPEqM5MvfELMIfSJvYd06Up3oc
lS7CsILQ8ofii+N2l0fBQDT9+ah3noGl+3xsK8yHHR7GociEYbcAHeIMKFiMWNX0gdktzXHVFt/L
IixstzrUbrLzff60gyiF1WeE+kB9OTxb+toQ4fe4zwxVcY19ad5ykoxsMLexbkic5SdtqR+ErZ8W
uiWp7ZY7XEAe1ZARDEeLyN+TsGLeTMe1Q3QU8sUIJKtmU/OzGCz0HVMPjhgfdIo95Pl4x73TwJoQ
RM824oDWjGlFLLSsYlkTshG4o8BUdEinHMDDLY0ezzwuc3/rXVln0pbDy+FHPnUBbD2+kpZZXOeo
EdnRnGs0SkIyUxqrX/PUxRhAh9uexZbtu7UbgEWlKoOvJ7+KFSYHO3LK6NUFimROTLk9HtpG4JFs
jG4jaFJXZsBcKAFnF/tVdHYsKPRNt/+6w0SSptJVOf/PEMe/mtEZeGN+h4GEGtfudi5lVeO3vmuE
c3lgfOF1rUBw8eibUhmIcUZzOmqa/wSWho0OSAFFrlqGYFIqhIWSh63H/KcDWFKALCxPY2BjX9Pm
ICIz9X5ZixzVhr+QFB7eVZKzJv0c9tQQ88KmrNkr8x9RqFbhs/Tp4ejI3u+FZid+77u+LqC0dkrk
om16dzxZKb07EW+lNNrYJdy6bba56QtQGnUXyKkX98lw+zAXioF6PkDLFNAgK3pw3/OG0Fbdp7yg
6pB5yaL7ZXq+eDZjNv3tLJbwH/LEW+jUCD6tlcCTHx/AttCgRVrJ5smEejmJukkyoxNsvSPYX6ym
FiUVpzphQ82Wv2nsfwXDXiVeWQATjjQaXmywOnYuCSxUuM6ccxKRIJ76VHgA9pmJM9qVfeoXj16a
tYcLgBPhDxaEB1fmb8adxlZvmOWlzIXBAEHcHcY//OByNbpVl9LOdj8EPF9FzKfJiS/FM8N7jLro
byGF8XEm1le9nUbIf3fHLSkxxi71ieCTT+JPEqzS5KLQcdJsyiYgccBqZuSdxsVifBS1BxtUerQr
KRWsTWfxq6WnoquNG3DHaGyNCfcb/XldVTQSEPZEDz+viaTJhUDhAe2G9prBB/kcNMutsNDM1x/G
SKIVK2db7cv7IAX9BhbXMwA2IgE/paHBZTrZPanfOOZ7y+03WDvvTmhtm65KgP6EzynRgqzHjSNk
TOPgbMM4SsapGMRQClIN8fId3uoeRMfHHe3K+95rriXECOYCXfBvBqp3CDKTQFd2pJc2P5zFaL4x
uxpMVdnDDiy42H+DUkU7EftuAlrJH4DpN3a5uucn4lDxzOPQ/FWLSimZFOKx+zzCeVi2H8Ku4mDa
RJP/h5lK7ljp7zTiP0oiom7o50Aga+QvkPI6kyDYz+pANh0ycgkhAtUlZFJJxfLidH9xZfAOQ1fr
eupE4w8/b/786DmJix5ZAkwLGHrEkruLOYCQoF0uNKQua0TioIhdUSdaoxYiHIvsiHZ6D26blOTb
+xUpKZrtxDj62TA0aN4+vTIKwoQDxXbfIYxXKUWc9i3h3zwT+kLAPwBjPsgIoepIWvffUlHqGR9u
G1QBlmTJ5jMRGPoGroxoEjDTvQcwo6vhGUF3A585YpnfUZU+79Sv5FwjiHGY/IDTvPrsoSGM4Js+
PtJ/BpKHD1gdKq0ISK1Vu0GMJvw3rWtJdLEERXA7891s9LJ5QgDO6ZZmqIGncXXSr5Bkdgkm6mnP
1oErkFeHBTP3rwMw1vCqVPl6n7OcV9vga98Gtsdy5eRMJGvaTY3oVrmmJnpGBq1Jh6GucJfR3YZt
nnNGpHM8vUtmUv4pA2hTLsAPN2hk7/dbu1JnjCtQtPPa06n6b4YQDWCeO13WTqBXRpivx2vGKD2G
Hplxa3FL2ZGea5t+vQpdhGVOvGHl2kauyQWMmLrckJ9zIklC3l7qB11S25YczGUz8ZfAimFzEvu9
MaSkDWXUchlTPY8hA2g5sfIAJqkTUDtuYTFxUVVL4nlrgsqfJjETHyAAkQxw8USnmBs05gSAwE6a
JDRmL/ajePK4OJPKCyGlpXjAb/oBHRp80kDEH4zY+Rvur4nd0iPSHfEPexPoaoU0gquCk2iSH6pP
IC1/45fJLLE9gO7vptj+8CC7lsS3JLIrSdxp9L4HL3hrZlxXNuGW6FgEbTBa/XXL9eIFTC0LSKgu
XYKni4IF4sQ8GxLPnLPq3Bvtla5jANXukPe4PaaKtaOgJe0gqc6eUjVvjCZDT5RuMWKXzisWAjmz
jJJI4Z3zheVQr+LBvy4LJ2T/dar1sbkEvsI5EqL2dWRzFCrvlTdzNZT/TabQEfEczbcvl2qaf7XD
wB9Z7sbkNDvy2Ic1P4xa6YEn1+Uw9YHp6Wcn4brP8t4IxFfk2AibYy4iJnZkes+MolodUs4UDffg
785TXdrUtUDvcP/dAmyQ7Od2+ibabgB210iY/NzZHUFshYSPHo/pT94NiRhZnod2qHsTXHAxAcX2
0rCPCebwnlXe4T7h7YKmY/LmYtTARZ8JcwBrNFFf/FJIDUFAJMR+JvLCECfAvKMUO1/ha69vpOmH
LFqRVsNHNRNDQmv8Q2kHfs2dZYf8g3X5RlJty22hqVCgF9OffjOWnrcBsD0XElRRVQa2jXvxXUUG
7JLDTodDxaJpGOClSxroOwxyS+5eQf512Gi9SrO+oOObJwIM9mqptQepvxWD2Lg385D5tmaZTWTb
MYWmry3CG++3goDY4uMruZMFllJ0bp0IjwVis/US8TuiHMkS/pZ3F7s+zPhD7GvlzNK0MeJDbzUX
ydvO6VgbsQ8kspIkzCAaBdmu3CDi/4bN67Qc9n4aT+VwFjcpevStxK8QPwyF1WXg2toAcQqmFP68
7zAagQqfJHRUEpelvzbjMGyMBDc+6t6++O6la2VVHPkYnGtMpxKU7W2BdNJY9W37sMTPLpv0ItRN
n94nrcDx1Pqep7HA+P3j0/G1ejOvED7KIgLDN3rK+nyLtCqls5SeCWyAa7PmH01dOtehKSz21F4l
8C+QVvep1hP0CTMQrF0mVZn10b6ePO9i8WXHeDe6cgZUSKninaP8PIDIWONktJef0Lv6qzL/b6TJ
QsBhovAftd07P0Zakw+9C/MeShBz5JdwEDNALiWzWHfz9Rm89Ka5nu5jNVjWLJ9sinMA65dxH8SJ
yBJt+H0sW9iYZ5J60H8ZwG2UrrLgTlz3bOfWFt3LmjRGc32TOINJBWmXiDIj7sOmaeGfiSpezeu8
LDHxsDeL9ww+PlSqNAxUxUQAOAAghmTRWNcpJJUmgyPjTbHrI5bZxxFl3/t2gHYXyRYe2PQ8gH5Y
P38hFvRI0t6Lndh9FyiS29HIFzlDBqmgkBWipkcyFg0Q8tc5U6D3vdlstObhED4neyiNx0d9o251
Xod94XI1AOKF
`protect end_protected
