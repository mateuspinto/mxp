`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3840)
`protect data_block
lsxDSd8ReD7iGzGMCotiLDxvpdoayiPVS/kpJHhtgMCaNSRXW3aHbQ3vsVs4BZdCcB23TvIp760M
HSFHDpPgV3ivn2RK0pS7SqGrcxl64+yX03da3iQqxz77NENJ99VyANkoZ3ghz01yDOMh5ynmJZIL
OlV2htaG3LzKc05hndCMHh6bdQ7g722KjOHKLc5OlD7dlqVqFJ8Xkao+yH48fQRttCxIv8PsQHqX
FgLYpE97dLHLtHyAT8NDZF9kqgKIoErU5z4pPx9ufbEo9xfngTeJ8bC/Z/DPxS5tYYu+mDQ174jK
mu65twNkdhnY3f1Hy4+cyES8cnmcaZLboYbGV6HReXagC7HTb2Pb+oem3f3qzbTY4jGuFcXSiAcl
O71Xmd/RkD5cxi62PeyJmUG1nQU54Pm6plQA419FLWy2yQdFVCtznsdl242MjKMs9mKp0bQ/DU6b
8iM940g5AFzdd0YY8M+EIBOJjX5LuNPvO+4/DOofJlTN5tJxdW9i1r5qYhsQQpUzoF+oozYQlV8L
sr11rwrLFbHPp3qRyGS7eNRILAq9X8dqbY9VZoxnEr7cayu/KenP/Opm7jIn1EfVldSzgLBzI5Hi
Wzz0XcT7ufAZpsdb+tBAsZF94/Z2ygV9uRUM1ilfM+lkzETIB5G0A/5X7hn6CDce+gzhQOuUOOl8
N0RGC4idkzkBnV5NSW7ss+BfPyhqw+4ZDeaMXXWap0Lk5ZH+Uy7krT7qNSBZzi+j2ufrlSFdaWaJ
Z936kccm7XGu6OxpIsljZqoGMZHNTpb6zgeXdW9xY87euiqP2fhqBBbklRVz8O3L1eORGP1I9une
9MH2N0w8MvU2K9J26CTmRE3pDY+rEM+nMX+5+in3WUautLp2mmAQHOYh3LYwoL7P+cm25WhVHhIL
fGm+XJvky7CZa7SR5a8cYZa3zrqhDQ+n0JCj6d840sHtIpzgttNfbYJSclSDmMazmqA9vwCAVSMn
PkGPk78T8lqCDz9JEo7Zb05+3K0nwoO6jgHDfvEkqgyOhOaahuIR8yybyhgXdd+KNZQdQZV5GpIE
1xvnN0/bU6u3jQV9OCPdMXZc93C3nIYxwV1dPR6PXpM+ZaWDxmuT1H4ZDvWw9/XJvaY7t5m6MjOq
DpPYftE5ySzhzATnpxs6MV6CpIcxdY8kU/MCdZCLhj32JEKVcC+sJES5gJw2DO0XQbG9etBqIycn
h9DCOJqEe33DfwfUYAJfXdJ52nEA+jnCZ3KpwLDi94C5PtSWyhVcQ3ol93u9TFKBEVjUyP60JvIQ
0MRiisOd05pVtBZJcZHXnaLWHBk8sTnT4W3+mW03LjmoB/b+J+btlPS4iq12QJGFK89cqO90T9qW
/nTR0g9aBQ0iU3J41X3Xkh8NxQv1cnYDZSAtzFJD+pbqHYNAdeos6cAE50CFf0WQzlcsuwksQrHd
IQAfc2cWetEpaUzHAWcq/9rVh2KD3SSAfHZvPSefW5k7dlQLTNhCJDQEYlBcIlLNgcbCHy3Dp0HN
MuBGVyUNI7f0uAAna40nsXU5okly8Fw9TxHQFSRn1uqI2Cts5KCJ4OqCqNcJmafvvu20ZMWt3rB2
gZwW+7fYiJKB+J/YQAo7gYRuVW8HZuP74TJ+JsiVMXFE+hWDqWi89Z6cPqSScPLoz8BUwBkBDI4X
L/RsaCrydWv2df9vW5c4i/XtTixdGHsqjfdOlXMjstqXCDEyGPcOM8fUSfowd0fRrWaUxXEfHWpx
T+YnnZAQQ7+lKUeuQ/a5BKxgPMpoMrFva3SF5narMv0e4hGELVOKB+jFhKEo+qvKnu+ZtWVCFuNr
SJww/FiPLRDXSSaFMxs3yxPBfdQyo+rmS6jKzfx8tGufQUiYnL4iAOPAuthjCTUsLZ57dKOBd89W
tGy2yW+FpafN0qQiQAQfrqcAIP8GodxkHZX36JZosU8j4H+tt3ANALRjoBf49IhSOkpFhx5MPX4C
CSzOo0WK2aRkSBdcQzmTJDSbb1RrqqSAMILTRLF9Da8yo5uYDbkyHiJCCZ1yn2R0oegjbHFb0/si
opjRGxJ9QSUxsSLiKqn3J5OoTlfnc/0piaf4Q/M+G++GTuSeokp40gkEsmJDPsbEyGNY2neYqIRo
ZFHfXPWS1KFWPClBLCMKLELg7qYfLPLW0BM31p1Pf/rHSOxALfCb+OzNqOPPAZlK6mSCOhFC7nSF
NRJkjiWWCbLwCQSejueUXK2dI6BbpD9DB3luMuwapnBcOffaNnuhFR397SorN+Ie8mI2feqPqdKn
vjXrd4FqMpepy3jOyZagm6YNVR8E6vFbxUXBta7xwAxCPROW/f/irkrsZjBMeTQx4G0BzZskYGLB
VMkS0PVRXvyUatwM04DqoNXKCefO68y9RNw9NaMkrwGbCIwHseJMhkJLX8sNokT6O7aky/RFmFQu
jTl12JrunVK/HEb1CPiEBZ1pt8N6rn69ax+KSd19lHvXO4NaHT6Q+1nSbj4bBDGR51EhWJdnrqkn
RiNakHrIyemZTh7nc5Y8JVRJ/UD9Vd/dr8Qlb57OYNrwVf20y0cU/+nr/oOLaiSqsv/WIxMv2T0m
sO9oimVBr5qF+9wAwHigCH7Ad/472yCKfNffKVW59FJity5ZASmef2FOCKGs364/taPrDfjrUuyp
FOwa7By0KpOxzonFbyt764k0Rr5x2J6/0wmVV2b32p0vL4LrL2M7fIZ2f4hoPkhVLWJxMlLCJTh8
1sIzH9ZTpxWwGceUNSEHkKd/feJy/baxBsfF1iaPQ3XFwxAeOZngLPacWikymAvi8wBIzka7Tobt
CDgSHxF5+rriVT+/QA0SJanA1P//V8oU1N+MI+tRCEmOQhbV6bwmBW3BQm6JWUxEJn2/aTbKAvkY
7/jkPTRvnsWBIn7tq8WB9ShZfm+x42VHKO4AtxcZmoqPxH2jcU4m5xnT4zffzUAse1tPz9JVj7zH
l5fcGa1xaU29H1D/8LLz+LyKMSwei493D6WwRUf2aJhHEmRWBN54kwjW+jXWyyzmUtNvch5RoUid
4n4WYEoPY8zY0KqDeG1PVtvoWM0BBAKmxh9cXoHSYZg4YaShGA4cz0awFXk1XSMpQOlb+xxtSIsE
2Mv6W6cFYDJTrMOuY/NYF2jbEbmfQJfoQutGyYt5karYNVPpuuRHtggfyQNnZyDCWt7LfxVB3mM6
EU+5YglhlyLRmH7X6jebGOxUoSaZ4pNtlu4HC9MRYaISJPfyDBFQ5qDE699QcOcn6xpVEHoHeFHS
bDHp5/h2eoW8Q6kUonqFTKrpyBvlu77ywComsC32zG3d9GgyVCc5nf955AbqbNLaGsxtotKby4uK
vxMulx88/MJdWaJZcfWRxsRHpepu5W69femB6oXod1BIXwWgjiBUrdf0gDpMMNQMLNYoongi7nk4
VJhhpJjwc/5jyckdVu+4fqRwbTLgbQyMVBdMOWYRfon4fwXMu9Nwl2JjhZ6ymgQpzIauRsAtxxr6
ivaeWmaXqsdHHKNPqmIFPf2m5xiDx4Fusvb7buCVWeSODRr1MH7i34Twq31WPRt68zqjf3Cpp15E
OAi/jtfEoxQa6ujbAV2rbN7uZq716/YP4y2V1Wzh44YMyxU0nca/Mn0lAxGf+aCReeTfU0fW973C
CSrcs+nM3Rp2NNfEtEJQVZds757vQjUKp1/CLak9WC4oSTYJrB7oDKlqH5KpAkRZWOuPabJ67lTG
zattguOvC+DGvJupHJCxPbIPimIBDeJ+PGe/62OUrqz9o5J8pd8UO26/frfJco9Ie5QRhecxuJP0
ckZsqLTXXWeV9gj2EP7uwFJibY9oZ0g64/RpL6O6scec+aICHB0YAH16qdoC4SUXg0hpIMSzymoy
iaB+QtOhKbVGxJZ7zqclwgodC1kYQSzJjpZEdBnlWfwE4zezZKEQ/e/W43IY3bvma4XmdDVF5C0z
Rlj0iNWjqOMLJGj7iWepM3C1V7EqrpcEtm/6RSr7pd8boKubMOkAQwJtLvcOdcUK4ac11SjuAHPh
JydbcbXzseR9E8ICUQ3SdtEn9T2azKbkLgL40mwEV1uj43zu4V6J0mXyBl9MBqhvxCVl61cg0RQQ
jUPNY9F8uUbN2oa71ZJlyT5PS4DUoswT5syX0PrnmutukAb3SUeL//rPwTBso2rqslqPghivqyZx
6UdT4GDcZDlBM2jH5mbYxevyytjNpscVDqlbn2bexsfztPmpFeDOR/3T196jnavsbn/hM6fg6gyW
cM8DxEOS++2Mm/iuR/pajItQLnn8UzM/L+TlkalME/uRGnOKXr9yYHTO97qosAAatICCjXwo8e9N
PQVgVG9Oha03Pb8VJmYw5QmSRb6u80IGF+AVkEYx+uvodkeZhqA2N/WHEjfSNpEZDFXh3yPlkl5m
RGUdzEa6k5nME6hAgi/hxxI4HWeDGk8E0ETU7Ft32hVsoaCWysj0hGlcnoEDg7S2JkX/08TctD+L
pA3ENsshKyOoin9r6F1p8byRhINtiSPBn8ZehZ2ojCVZERIHiqw4UR1ruARZNkEVjCaDGM2FFFaX
nHW8EkJYwKenbLDXx9t7u67gnvsXSDvWfrKNFKUQTh7F9tofxsmuq8ocFGxgEe8n0v5lieZcExuv
H2bhZvxfr1CkjqTFvz0kAySRRLDXwkgVo5AyLgOjg9ych1OSpDImSNJ9XYlDO2mzqu1B9/qgIyj7
CogkDFFGYLYBQZyn4OaWHrzsdl6Q3XioQoMJzvPO7xLRmZGZqemdJvjEjDCFB0LF+8yzsgYXniva
OsC6+wZzX2Iz3ECiMCjs/xw6tCIhfxufYXsKbeW+Ten+EYVUbCirW4bvYD1PvHXbigSf4Vx//57j
jnV7s8aEzYIvIM1mIF4vnvBjbTTzQcYnVgvy/RVliSSZBeq20i++/Fvbj1/7YfUZ4OBoUqEzVkBH
yhIHfIfdtETaUa5XwPuHxF9ebO1c6pzSanOmu/8vIsHqcHa3NMM9V9vd1kZEJrHWjeFoaTvPkLQo
iGW3YqfSdwL96uoRUWRqdmEL+1y6XEz5ehbLRN5SBp4eWS13kIIf3D/slbblIoBTzgB4qBL0gBuV
8L+AsouFAkC9k1QQoRFodBBbyHkV
`protect end_protected
