`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17472)
`protect data_block
PEXZ2V/xJuFTLFCLfDR0NzmxlRc5vxeey/Wig90xMBNdjimPXG/BAj6R8vW5kRzW3SOuzf5B3Btb
eQfkdw6PRGlOraA0VjhBgDeyTYgGg6eGhbcxfcH8qnWEL/EzBQj2wm5c4jVPKjzTbJjIYaHcbE1z
GsFxL5GldPF/nqGzkQmVKKRYta2zSVAoy2v5DB0q3Nl6fDNwxm2lhUKmhDaU2ZuthmyI4jfNUrR2
aLCS2icmeLgPPscJq3pN8Q95j6rCnbq8Gx7jwBVzdyhGQbHNMcY9QGlDEYXgtbhNQ1Rj4A3gI8Sh
6h7iXgvRAhXDitcnvT5qnvaio5OURLIVVHQw02om5nGBiIIkbMYfoavy6lNGw5b9pRCvRB85KdKz
GzAMA09Dyd3iX7r3MYH4vZU9dMxgDUFY1k3p4XAMFDJ7SyLOy0cXmxVd1f+bO3NxDLiS3OQQ3fZ7
YkXMaKMfE5r0V/CtsMtTI/hrWU8sVHuuwBc0aeYci9YNIpw3jDafSPh+O17t8ZGrD+oFHDSs/dG0
na24QArm0Bnb3iRWqAWBCNavH1ptR7LaS4D0qOsqD0Fgp2dHELpJq5ppK0jic57nX/NL4c4cIyhF
VDsrvKpZY/7AGljJxqcnSizJlg/ho03kfPH/d7t1DhTqdszkf7lKVE8PJfgcLcXcFs3pCvYAFNR/
hdTQvlDHwfmUmmVJG0yqXW953zdJtK6HFMOlrauPYMpGP/acFw52rJ84FZnVk9vPatFg4z/X+n8l
n66Xuj6wprpGNVejy2+VEKDQowYuYzszq0biCTalae4zpwu0brPakvc1JGbUjhP31z9BGhXiYMp/
bpCH9iamxmDiXeAHCgzkrq+p6TF625nMMcBpX1RGAF9GzYs4B1k9gbxe7QPD0eRWKDnG/BRy39Iz
M7BKRgehLDAqd3L9EJydw0E60GC/buwq9rDcwEfJMOK1LxXcEFGf4hhfJCj/idd88TfQxm/vhVzw
RFCADFzOE13MKJqQojPiQ5wDTPptMeoXv/IyfRaFNgeMILNPDZ/yeo3IHmA3335GVc8wmxY4vNli
gxME8lnloSNA9ywa0noFbjCXQ7ymzJO4DL1LAytkklsPc/w8gPfRt2ebq8aP19HecEIu7wsfJS65
kU2SJrx1UOwi1lN82l7zW7IWCinUYwJvFNr8PRe6xEyZBHJsfOVWWWor8hlVGlzhJ7WHoQxwfCmk
XYmNaXPcS1JGkpe/+HM6+hOmZv6S4HQKThT3TDNeddpKNstdlJJnbtURS+szw8+8tsqXXhOH0YHZ
lzr8NUNcuFgLxmmkgRwHNRKqbxiKEDrWLImSA0rJQ3NpfUcEHV2AVugN3cYgIbW/bpB+QDmljU5k
w7A3K+Z/RbyBYWPtzNtPf13JsTzVI05mjq+6LUwnL2zUjqJvzp6pL127//fQ2vHiQGVxIL4GkfM+
CPd8XLmKfEPi61F/ZUhtTaarqM2rzhzXSiqtY5oaxPt784zO7+8qqBLE/9Xyz4aNBprgpbRSsaeJ
9tUUKBGanFIQm6LUSPSWh3+uKZ643TfnTIKMOWdv23hjpoufSd5nVr/MLUDuzVibfo09azhQokfA
iUTSN6csYyO9pGf3099VglAszjSxUF3He/DrPaVK40ysc1mF8+ZMw2CsXdFFyua+m0yUZNMJd6ec
xXqiL1T06JE0Tf5Nf4mOWW1dmSYx1RH57Iae5/9vjk8vS/EfOidBN5UylqzkM0ba8MTlVWQW7iz9
yOFzhkteVeMGpvO345oT6rdfKG3I9FgG4oEvYbM+doFkK/VQPNTT181cPcPlXMe7iH3i7rA2Jknj
oKURkddTAOQfA3eVynb9ouHmgN9HL/T6/S8XkGaTfQPbbwjDRgK71F+Z85R+lMcCpKM8zfABR866
u52hY3GFhH/ScW4rTaROM7NnX2X2QDgG3lCtH9lF+sjVFGNFCmlIhbYkSpbhgE1ZSuvfguhDcyOh
rWe4pM0OC1EmVPsJaw2aM79OsFbA5Jpj6HSpbN9sraQbqg+p1uMBxGQzz4M04EJdURmZ3hxGI6sP
yk9+tg40lb3QdmPAGmXE3EBKBMKzaMrwALkMAhvuqwOdKReo3j65WIP8g0bGp21nvPVcOx1qyIm5
1XPxp05VuQ+SGsjHYvr1voZCtcUwMxOATBKAWuqURAvCR2xVKiv23Bn+triVJwXWir7R4Ak8JvQv
Pdoh/Qea0pIuI7fWTKRb2hTKFbcjjlZcRp/+lCDC8S9keif6C4NTWZpUrqWV86PX9hSYdOb2Bm/K
mhMKpzl65e+7y0eqXnLLKd4hB0eLwEHp67j6tbR5JkFHML1l4qXgZO7IkUvfcwT/GNFASDO7fR5v
8mO0Ka+9X93mINLMVoSS30XPLuHP5rJG9AR5gTih1SKj6uQ0V5rC8E2zo8/gSWQ3xjLZ3Zn7Rsk3
EsNtPsHLuUdSU/mrfOSU1r1ltcGN2vWtq82t7v24l2CXFu4Fbc0WRxvon5CxmgTX7Qhg9rxF+r9t
yUS50Ns3TIOp9bdxUpOPXtJxRAWH7bIPykdvEWz5YJbX2RFMnMj5O5wbJY3nxQToKMxqYz1tQE5A
2/S60BJHP6UPS3UJWwZttcLaKNWW6hwuA0xx9cuLWWumLJsSTKsWDH0hOQvl3JNxcZoT+ILxVPcs
jeMOXgvvZmUyS8RxigDfTBmLM3wmukq/PdRB/+K064qvTQIKsFU5YfZO60N+GrLrU7CsRV+hB42/
BseIq5654Ag1Gs0y5bxPdHzs8q90ZXmwmeQdK+3ej5cE8UitVDnHcSJtTJXlLPuShlfrnz3vKjv9
NPfq9wC3++G8ng4m4vvVDlkZAQivlQkxg91QSggYvfd9mU6smS24aWmt8IGK6tnyzJTJepvXf8w1
AcrfHlfBg1IlnVU1uvgjgb1PZpDNYobYpFT5eXsSecHeeVEo/cQbKEijfJ3MB0jFlSs70COzjEib
OlR+l5pZr7SQDreYDQhgKxKn1572LDGRkBBJvSi15AU4/142S6dWfN+sEC4mnBzsR8hLYg0riDHN
LkIWccrnYAxo7C/SlTmhpbgQM7TIhZMQ6Y0ZYa/RUtOh72gbtPpR73wxeqBcH8E0thOVo/jHk5XG
m6yN3nmvvWGEkPyRvZkqMMft26zXkoEDExw7eWBRpbB/WTkbWDIAOigN3cmkiGBj4IQHZoUoymZ6
o0y5Z2H+2JguEjh1PLNEpAiVfAqmSYiEwBKOfoH76xdFf+CKKQPUzxllUk4GY5IFR0sdb3Q7q+HP
dbc2Ab5r/byyg8taho8yYKYbrjJFigBr/QawvHyy/bS3Rz+cuysAca8JNbhdwYGEKvPhUNkob54K
ZydJsF3FV/7+SimmiuBMfLeEnkROORSq42l2fhTDX1VHIZFxzL6dbTRUWLcRxPpv86cZEXoJ1Oza
woU3gzxU3g4PI2q5y4HvP8xwjhTW3WC6IK5zDS5dwmARhUCr/KcZaP8ybOYqsKWxUib8wK2plckl
irHZH0Ai04zNyS9rMy+GvDVnvaHuiZK0DbJEthc9hx5IR0sJNK1HsnTH/kPeeE7ijEYJNDyrJoae
T+gPbikztEJRBHkUL1SxL7VqRi09ny2pUdaBUClSrBwRUgaQWYy3krg3GHWWd1ohTD/3OFxsdvAs
oM3R2Uz3TdB+rDWpj4VrzgAPK7YsQ1xkbjbpCZc7KZEMdisT56TrRmq09LRrHZU/TjWGsB4zGQD9
7dVRGZQ1ibR5QgZse/4UC8ZjL0NsgFfYIHbHRWsVRgBIVypwTIteshCZmEqf3jEqO3gg1/AEuOfM
Ny/2WJi7cfzvdrPJE6jpiA5R1VwbW/sEEYexfyZi2TpzIalwmjNq29VbmuwWIAj7SV53EWh9PeXk
wP6SRwNbJXkd++JqVaRkFeawzcBlKC+nTIpJsLP7E5W7EiiHl/SzJP10otva7wRh7o027qHp9XPf
bPrirM4U3LT/w9WyvLCbrqDzNeIyeiqjZ6iu1GtJtTo7maEwQ6hjQ3qVeEPMCO+X4vnoMCJALINq
o1fRVj4Zuh1OZ8Q1P5QXM0aiaF3SfWN8+9YJUI3LIdvPxxIjpcpySbWR5W62CxeUcmQP/FYirnLt
z9veKw6bZWlWxTP+/i2Bm5iiiCXSzIJDGYHTZbs9rAg8dedm8xYboAN/NziBmDGn9AaQG9bY2Lq8
RVMFaXeyVD5Sa+oigzZh/nGTVH8mdI8HgX0aNch190kitNkyaB0SxZgYEKnkH3HOXnqtl1wgQUgx
oR8s75ux4sUTJq2v81dZLDQ/bXOtTk0ZNiE/LrlZ4iSXq7HHpw9ogZT4f+6yV8l368CQkJhoSncZ
mlJm1iDg257zioywy5pAP3HDttscH3xMIu31A3fLQU0L4iKk2PEgtMRYq/+BmpyD4lIaHDrvmulh
XUx5t3s50103rLY+nAN1qpxhzJLXYKrkoYeDa/rCXrqCXb6N9qp5PdDpu/PG8y+CU6LRanHn1IwL
6HEj/nOuTfCdYWISkdSUM+6i5Ftgp2U/cGOVb0TKdh8A7/+3hb3OhGFhaQmvGHEuBkcHybkGXrkn
jBb5Tq+9fP8F95eV1nQl4HUeWAXyaVeNWsz8odsCgyjKuFpDJiWWVqwUuJ57n1XuLQ+J73cE9elp
oBqcdTTgd8xRMtkKgeQGSIKHdxnuRnob6lr11nNhF/ThAgpMfHomGuulJI1d7/7fomY9sjEAu8ch
qiDmX7cbAfoK4JTD3UvHw5JrFlfczWFZqhRQGf16zLft8q64mKX1jQg0DjiffKkpSWpZGZqNUzQI
+M5GXnqkw+kLCXnB7u8yGT9LKVdpa5BotRnkrZPr1YEa9D3uGKnnH08pgGR6jzDlAydKyf2CRXWk
BJATDyQxho8SDoxHOzIq64HJGHmV6uqjDv8Htw5M8BAL2WRV22rXAlo/d7qilnJKcwGAEBCCuznT
twnc0wdgJNa9hCWFpHguvOysRi4bWZs9i6rYctT0jE2Oh7BTPE2Tio4hkfsbpcBp/XHTcJvKUh2j
nIxS/zkA7wGOX2oTziSs2aDwlMjgb3MJmJ5qBjsnCV2YzZ/vQFWYVq51HXyHZ9nTnJT+0U/iP9JP
IUbTtOW4vGD8H5rShq0R620OWUQfS0GB1fFHzvE3a7T5DasWyLAY7vX+xkQZZQ181oERWEB18IdU
Yc2zKVmR2ZxE1orxz4LyP6ILqaCbYltHMACLZzqkMCmYm3JCYZDQv7TgZTakZTzwLIvQbJQQ/gUQ
zBP82imCbNqfwZhN1n8rhO77AwL9GOmCJ9hj5BjF35/7P12V5MnVzUEjTbxOZekIhE0RkJB6qa43
lhIF6I5xWNuPD0tSFTYR5WtBJodFz2xqDTgYKlr2VRuioKae6tkILTyOQjxodpMhvmsaFvIwIsHH
Y1aPxw1QnvmOjdC/Rb4/AisKQ3kfwkkZz87V1je0dkO7Vts/OWowePHTDG5aTJr3QiNLPlP/RxTL
y1hjldzfYCXb9tCMZBpXYFrevz738bjg+yuuFyjO8/UqMkH/LwwLGMEJaiytLVpM4GZHPVa5hXnP
hfylJnd4P2fEcTfcJS2aWMB9bwooL0nitx2oioqvgLhmt+iGqo7kEQ4dAqlyCRUUUA0CFiPqe/0R
jO0nngXOGd8ZhI9smRr3NTNgQoSt4LFKM7pG5v6Ey20ZjE754Qnsl9BvVokM74Wa8+sESQeI4l4B
vcB4e9PKktbUf9dvYD6xDmj0Z07RP81RVMxc2O0etTDuHmxeCtJiKmu+1yo8WhVvA19FjTKwGNd4
SKWmBmvKl25QlJNhRE83S96EirNmbWSjyy5e5VjPO0Hs+WMwLBMQSQlmXr0lwws95dQGQ9jtW3+d
RTa4wVg8UhI2CXwTjePvzoK2E480Oh1qBoNdXODwUwJIGPRy4d1TtKzM7utEnp8C264lG8x8Vgao
3HhyiXAs2NsEtmfrOoo7aQeieTJGX1Psv5VLRr4Sl/xNrDIxz4BX/pEoVkweXW4lLaMABYl/3A9i
aGxpWpmgQGNbdBI86L3/gaSFaG+knfL0Yy8tLmiY7RuFA3GP0DP2VcUoR4UmXX0LMNqqc6Kjwlsb
McRY9efgsRe8m/jDcitODkJnIDaM8DlmEQ/8DRnUasgfrr5qgwGLREuK4ulCrK9zD7MU33aKg8b0
y96Bek4tu8I8TlLj1U8h4cAl1rSXWtMKi6NhGqN1/kU1oGN9HDxdzfmdB81q5Ky8n/YiHrLyliDY
TnT9j4TzNo8rVA/QTZRPCWO1KNlPFZ0nU9ny002v5sIxFB8TE8Km+MgIFBgUm+p+pm9Mv0gWbwTu
tvDr4IqIDOwEyu8pdLRQJAjjcuvC7pqLwlyFJRr4y1p/bEMYBpeh+KNHjUsPE2ZX86JLcHWTS51z
r9ih5xgCasaXzobY+d1qyQE+9O15bciNDjE+DWlOtyluh3x1DwT1MtWZnWr+44Amd6xxc10ZXB82
Tby4UblcmtUiE1rhIRGdTA7ZAMqpB2yFemV1IG9Bkau5srdbMcrB3Qo1THJFlqtPwInn+SIdlqRy
+NVx6buE1W+ncYB49tw9GV4+qMMZqY6tb7ryXGHaIty8NEVcAyXIOd4lJM4yfyuvs4Qm4o53somz
uKif9W5kzjao0HYTtWsB7O23YRXaE+LvnGvmbqN/Qo+0080X6tZT/yzTfmwL21mOoX1wxQxOtoJ/
Y0UpgolFPM8cicqfnsyckBjJQoJV/b8dvfIOgQz582g3lasujk5+0rczwzCl7B44C2JBrtdS4AGI
Uoc1H0jkpAHLz9f2jub6VHPY1x3Tggz7wHk/z0BElbmdb/jwvzFAHzIujwq7ShUiswqwBxKka1+Z
mbE9KiCfW5f/GS5ZTmDHQSwtM4yswLLIAUfSNwD8Qhg8K1S/zcQwILHnZBEXDAJsouh6F2ZRHmdx
gBCwIbFquTKIUQPAQ4JXXa0xgeAQ7adcQ928/PJFIDUE0s595HUlQ7XzR6sUy0egLpBc70Ecp6EJ
mtniu8n+V4X5sUHFhyh0A21srIsLYGTJ1Pb34ltNV7/88/dMYYJlTvT4E3MvIYfQYTpSaudGDPcg
BWv22w7sJy2i3fNva9Aaat9mh0+rNyWE1HTYV5i9JHoNVIgdXt0Q5ViUq2hmQW0FvKm7icXFy9Xa
xEn9p/eafrJ5AxYN1bSZhmTJQFHe96xW5g/TKPciPh+PAcI7po0e6N+2/4IJPiOQ+6Qbc/vs1x92
P4lxH980bTjSj+MfmoMXLKcolRwE8OOqHu4vvqJ41raAehbpF8d7D0gaiB3NVWSP3tveslvoT9H8
R9riZPv60DHZUn/MdRxlM2guS81wZUNllwzrEFIuKJEW686fRUWoN2eGEcx6vDJhpOeKLF0vtqcw
ITR1cIc7ZAjz8YLkkJiYILhTdGEpydwm0LR5rYL3iBChVBouyUiQRr+ZFj5j8gt/gj5rmrG88svE
OFY6MHBT5slzFiRwbat9cEAR+f2i6v5U+c9s76hFUJxSduaNBFo7wHVVieHsF+JubBLBZyNRk0mz
BfiLDgOVWbLLplvXPv+qGS/7CGotjbTLiNJloNgYNCMaMLFhXHpFgrZG4auJw+n/cFqjGkEPwsH3
IGjwjdCpjFd6uEsiXmY4mLX3pgJpSl0ZvJ8JKquy5nnEi4o0GjOKdNy85qMVca1CzYC0yHlsnVgA
ka7hII034rFuhZ9B5OSa5HVCZ/gZl4PN8XWHfONwdufMhJAMmdi5wCHlslotv/XxefCx8waQVEWZ
9vNvlFbqk+ZtyOKjbof+/lWzu+y5K5jBzuLuQFFWqV1G9pUMgUQk49TOl5mYUEEvv3Kt0HN3gIp3
1igxMIBKCNYTnUc7ajv8sTof0qthXa9V4bJ6ZxbQEcwCF6WqlBDmwqK2zlN23UHFrMQrUd42Ty8g
OC0GPRutkYz0AIBonVuJvhrPNxBFPIgl0JpecdmDTL8fhuL+JY33V6T6PdEVhl/dbF3R7seMfl4X
sE28dQXcKosMdle2IprR6qcXEZyubxGeRDexu9Kb40BKTUKCZjuwMeDSJ+4bjWGkhh0jGKXjf8W3
sC/WNJ+aVPh2X7txuN+RVv1V/sOxgIyEhpEQHirNrhYzHUHUm1isJe9jqRykz2KqfT9zCAQFqCjB
8Ud3wyRBz6e0G+JJ/2MuE7V2NVxa0jfVA22jHEQrgnU80FUNPfwe1JjiNJVtM8tOBTz1GIXw/0yq
rUhFU3fFJBFoLKpMfW/aI+dea+RjlAwL7zvc8/OfdWd8yrvR8aiKMtWFVpaH/noOSVlN5QdTrg+0
Z8JGOj6LN5MaP8C3vgOyBJKWR3dc4PO5yWKV2AwucIcdNOT+RCpmeOndZFXCeDUYPHozYceu5gPw
OUxe3MCSMRZJuzBcuqE5SmybHbWQ8gXhvaNi4koA6cSI04sjS5oQbi9bOM2czbdrvM2ZR1BjLfiU
LZVXRr59tNiCwB2poTqfi8ciSJk8JEm4GkFmGJndZywv5PBJGhgir9RB3JMnLvgBmm1AUdWuAox7
Q6wAzWNE9/ae93VgSTgegaFhKo/NdE6duTOYAzK+HHdi4w4kvyw5RxKReRfzXlogXA4HfQxDH051
SmCv1TxtmLsx0ToF1cXA4sRtSRh7KbDciESMe+OZW2TYsst7d5c2XrwrBgIpFEFkXGRIOhdXa023
WSfJwKTDay6p5kilR+NVr72T+VuWjZnjyja/D6gzjpPMv8YpwTJ1zYmPCcLtyWKo+KEg280NyF1m
OROEfpPV0knGUpVBoP8HmRvUPIxywuvkb+zXN/mJ8VgLtTR2bmSQtGsxYvxm6jZyX9EcAvAx02xx
s9M6ww+LXjsqFn1QVgbi8kVBQRzyllHohub1b5Fpg+LIlZxO9UR+dtvS6oMharRPYvY8g27rsXs4
+sneypmqnWWP73hmqmYQAzWl0hybX213fLuOwT12+KPwmeuZSIUg84sqzaosIZNVM/worVDtg8H0
J07jbr3gVgMz9vwDfTy0Vpoeaks1z6L9Q9W518/gLIrJGWc9qnyRyWZpKbzMLy1OqS/6Ll59xQ7M
lBVaQ2FxsmOEkRqdGK0zgJsZNOf/uma1kbrA4InLgXq827CJcikZA3bzBWcvjEwblZU2szIqUNb8
5I7eLvISJr0W6qgta3toNY2p7zF/xJW+YBqCZJ2qLJGTcE9z6P6i8qm+MetAZSuM4gn3XtYO/ZbV
PqtX2l+IPKZsHHuUDBbkPzKO7kOwkqfKD96OgF9vXrCWTig+ek2PXVKbAzfEt26+KYv3RYpxVhe3
FXVzj/yTyV+NwhvOIh9BvDdgdgoanJCFUevcynE2ToMY4upsAsIuecSiZHHeLOg0MxhRAZNBS2Vr
oNeBSbjBQhPLeBt7zIUH+r/FCb76Wgf6eL3pE9lmmj5TA+LaeNzuxzrRwDcTf5DhymROSQdf+esf
QVjLQ1ZSez2zutz9lPWcoz5YLRUL6ZPbPBRtXGGATEaDdDVpSs8Oxwov1AuNwlChPOLF7xeVjhLm
V+yZ80OOuL0ZWIA2r5DndOL5T1Oj4fb0yzKEUB0d06KxszMSmmiYhFscJm5UkrCpai20kCwZHj33
v4GDl/iSw974CwWiKD+QRVRGqTZ3hjXhZoQRwGA/x6bKcS/91vKWSpi1+c/gCHaylgJ63iLjCHju
7QHwgKnrb2lBrGQYu8Tei8M/Ulcvum3WoZ6jEPmE2J+QQqA4Hfffy03wTxxmZKCX10ebM0OgQrX6
twIsnuEy8ciF6/94+bWQgQcapOnqvKp07b2zbmxHbwD2tFcVxStghxRHsOyAX8vFYK+W7AdQEfcs
4AVHgz45ALBogyLI222A1kWRxPWoKg9iJM4Zc9B2EvoSFhghH81uLx5HPg8RWfPGXk/neDr4xnJe
QMUX6iDtMvhY0DmZRCtmsYGJCKeVIqI3SQZoB8YxfLfh+ISkcbRQWZeR9rWIKEacDeOYkkAQLk6U
TSVYZdVu2aBlXZ/kwDyQS2q0KFM2djn6uo6hF21oUCKtf1FPYgmDiUQOhkhIc3GlyyqGR+gy4HSm
TttB+kBtqoVDYqMcJLcHECGHZWxZIRRmy+YIzqOyVdUgHC6FftgyW88WS+PIWyd2/1ObYpfO3Yrn
BV2A4JemMbUngSxXu9kuhl4Q+6CYFeUWai0ThYuKPAXXxOAzdYX17753DZKrbbm8XvCzPdru5fVI
cOGLMu+22Oz9zYeqVjtWeMvAW0lvSyRmyKrQ1TQvmMttRaq4H5m06qI/s0w6kByR03kO+4ZXcZsB
oeABEB948NmsEjC00l2LUCfqRjR4rX6JLYRHiOcWS2DYBtykMngFK8UNQj42vTezMxaup5HIIsOG
3i05KeexBnwsDXsJPngOgGLI0uZH/zJulBveJDsLbi8YFyOd7kxy3Z6RXmiYv7YCuZAiP9vd0LZA
3cOxDv8DlnmLTKmoVnUrrjIEULxHYb0wZIUmS8EgPUZHRqdvid0HRDMx78nuib5v+S+keLfy388P
rmBvS/fQE6o418KLBZa3gmJZNDPlTCjb8KXg6ivnvki+XzF7NC3k3HVmb0Ldo4UsSYNw8kFXYEbV
lip2QlHnV4JO+SZJrQBL7ZbI5g+bKvsdYBE7ijBzTJtLh0nkLseM6p3lHuDReeFDYiaV5Ad+BG7a
bMerukt63w45eU7ZflgndsygfwRAQpGY7p1uW5lakFGJBSikyOn1iu1T6VUv/D3dXtNcq9ApsmZK
IaYXOvvDBendSWa3GV115kFbBNrM2g8yk7kJDdm4w8Wku/8e6CoADxLai0L33hpD4UamjeKJtWv8
2sMdpG9ZBoNbEo1VfZSuCJqOnzqDqZMC2qhdiFxnwP42oa240PcwqzHPD+YvRnzOsysXG43e9Veb
76GIXXFsxtDjijgvCPuVNon/tDe+hlHOIJP7LJDCfnclmXqyXnNjujUeTY/yotSEeqLEFWBvrXSW
tXE2pfEcx3Dy+FAj6Ll54UBp4mFh/tsfrr2PugHM34hVSPNxTAAc5p5h9KW6cQSeqKgRrpqTI78G
y+FFfTzOZBx1F7DvSmKG92D1R6dJmXo10QTdjK7oaiwB7yfgUH6dszmO3eJItWsxApeFQtYhIVOV
XI0ky32fOBfu03PSTwFL7/2xDm9M8SBeEbJLTkvvW2UgxLEGknFNfdKgVcsSif/E+JP+9bpU+8Pn
wCvtugQhNVVK3I/TpK8RoTcqZA8mTzFY18a0849nAIJHfZmi+PtEFzOmqMCXxieElix2DGXdf9tz
0BfmLeI/JH0jnlQJkdYH4/LyyOfp7KWkaEC2j9MDzNAJDejXIkXPYcTsyPFHU/+c0E97r4Sg4A7L
Z08PSQVus/LsLKpOWTK2fOTGRxr9zMq6qkparKfJE5aqIkd4vJwcboBSYQ2gKQ0jKwpvCY8JQi3s
0lIHbkHAXl9mzBS0tqVygFNOWMj4kG+yPR+UuPTjsPGH/bMHv1ofYdd+i7OTwaMFJQkMS8zgh29E
0TrbCPZZZzAczjf5o5mp88MHWRcYu8UngdGKt6om3S34lQsa/JWzo+Sedl+sglNDVYWtLWF2D4V+
97fZhyUsmO7/v8ycjDpmLIP59KxCMKaYFEUHed7fmMKBea6CFoFEd4nEXXYSIgknrzsIHx/RsEbz
jp6iuD5uMCyuDKzNucwgcQZtB4Md0FvZTl/JVFxXVZW1kcUSfH3rvL2iZdMp3NEJKoPhZdKgmS+F
pephST+J0Yhn4ggto6M8FvbJCliVMEuwjhnoSkmDNXN5vcGaQ6CW8jRvQsdPLrRYthNsSUPrhOLz
4oI7EiXofjI0baiZ7O1XtFI5TDVhUyyA/eFZDlh9mRzjBYcygHGMHFZ7MaF8BDnaXq5HmDAw/QBD
wpsV5ifNqm/dV833WXJqwWWxFeVtbyF1Uboegjy31ksFinrMQxSKHRaPP2PFca08tMVVD2FSZYf5
mv2iLO5Pkyps3gV9Ih3QR49EB5JkIeQoPKTVCSoN5gKOfAzAaBEzaoRmAkTgGncjwS7j/2jmUZ2I
Kz4EPc8wbLIJXToGsNeKERbc7rNJdwV2E/iU7eDHV9lLv8OjP7HyQRlV8gXT3Kv5QvEkih0+wsvT
oMSOq0f/TuHnbjqpGQV4GDGNIu9kyPL66sSf5Vgkp0krbiBlcQAjIoAgZX47wukx17HaTIADhHQW
3QGG50MQuCCwqn0V8NeTsK649W1bzafmdnO3Ts+hmmxhACw1tvuCbkN0dPmmTS+HeaNXCEW5cSAH
WlDok5VnqTXBwxY4Nv0/Xcl6dnuP9Qk2H/H6ePwlP+QD9+EG1M/nbql095lOEOLD/nyMIa2SCCKx
Dpxcp7v5d5wMgKIjvIjUo5ErvTI8k/aZ2Wahl9MhB8rGKLpleI1Gn7yTgZdM0ONjeS432O2Lf2sq
egJz2HkPG2XxrXXYteDN/6QU6W+JKsJUmq84q/yloh/U+3o4GzHcsr7xAL20g3GCkjuGbJULrKPO
8yrGXeZWisDMZFq6otTG+psnQcZeLVvD4qsavWX7CV4L7lv1BQrmfuAiT7ifNgGRQUqXkCfOOytE
E3WoRKctgTIFvE1/0P6NRJlQc1wTAZ1jvtw6H1vvGp4Bd0dMSzZqswrWrrc+llUykZyl2YGzfcOU
PQV5ZyYg+ET1TIb0EVHJLVyy9J6t4rt1LXXkrZtQmSIjOuQrHNGRKfkF+lcOW7IObVKTti9jBqNh
nkE49k+ab7qrwZwaE4I/w993WNOtIYbfMt9ueajUaGLaOfuOnodlDpB9T9N3M/v8dEEmwDnxvjtW
Ivtu/MVfPyqilPMcANIUS4OymwNpHQbaQt7Jfl+SxgHrLNVWtZjMHAuicWGVDnOQ9tXgEsAxzn1d
OWlsrMbHmwgc7FBP/kV+4S9DGLoKmzT3k5IOUQgzOQ6yll6lsbqGn7e9urZ42IVAueC8EIgx8gsw
KntcSPdcYpP8ifZ0oMcZ2Q8p3G/l4HwX5WdnGh5Ia/iYpUGnjsBNTL28quW5JLX5IzQiNrsFR0oT
uAVNP8Qt23y3TAIodNqQc/GdtUD1depNZpbjH+O0WFCQrunw/K3odc8NLMpzcTyGREEkbHSA8ZT5
PGlcs/yX2eEYUC6sbnBOZQCbweaFtHW1wvOCX6UDZvblBkCFxqX6GPu9tGa51fwF4npO4RJFQna4
OgdHQJXOOr4E/OUs4ymZsPgAGniC6+xInKvuFkBJdjyFIiDLHh/fC34S2/7NK6++WyeSjYXQ2Bt8
GC0zu0uV/d0x4WGnEfFJP4nXom9gcVeGWCUR3cSct5QDEt2ExxpUCeSJawml++hHdnFQkOv9mI/0
2VZB1/omk7qGcJa6RVi5b6fe/+U6uZut4/Qw7HrBdlrJmpXERXDuW77hd+dXBJQsdztt+pIgbgM5
r24b2YQYm+Xc4We9OTIafq432UTqEfJdhpNmPVGvnaaxcbnIHMemHbGni+YW+BU4P7bNtXPM/nT3
BO6mrhXpaVM67O4BASBNz+fY+EYq8oJlWec2FK37okknh3QdwI5t99BCbfqpmcuFzGqiBTnmew/v
YDHp/1VlVleb8gSBPgPiRLA5DueicehmmW/csQ5YDUepsjBW6Y9qKziCZlKy0jdqbRVLBP3P+gsJ
U5p1WaV2qnG90zaXIyuJLqRC9f6BsIPqB3IL4FS7JePmeFnQGOFAK3GkkoUDQ9iJRonP9xljIwnw
r77o7uDi5QMchHzOjbZJa7sphKXsaLPk8PmIbeMxOK8nYnALcKtGj5T80oMKRWwK0frPLavjD5+N
3j1GhYf5UlrY40HwLYKWNaw/geACRWLu0BGkgTQhN+AkczOUTacfXysB7HufDTDtKG936hMJglrg
U8h+kD037hOenesOvUaR72emsp3TqlsDSXrRpIeQm0Zhm1fTgsZBKSFUf2Lle0GujZzAyckNgfQa
3OJE15BTZQeVSkBPLCCimz/n61ZCbNYKvuSN2fjVspe0d5nGWS11NZMjhABorpL3N+vdlwMlyMIK
+atahmLFL44LFufWbyOKVl+W1yP5Aq3XIIdpM3H26+FCEQr4LaFIAvNCdO31/vJwerrvwE8nQqtI
lwVOhaEXTHKHVY5eoJfEyTQx3BvCKA6yPdb2KDGF54RDgG+gt4/a8qaGIFWDmBu02JQh85V9rGqt
M3IW5KuWTrpwiiypsqy/eCYPUCdc/TEzKPTD0icpP8lk/zh4NxjfXoFeqRLL1O8vSMQky6e56Wfu
/uFoPmgeXO72lNetSWqPaRZ1DH6wrwwVP9PB/v1BZh/yJTQ1ct85UsvOBFnUiaG05MwuzWwA672/
PsDiO5YC7W7QW3/dHeHb7nTorpUnVCVoWpmcvHZsIic6ALACRRci4h3AMq7RiWYgopjskzLiXq5J
gAT/2FIqUrncHaAdZDSIiTfvqbe0DY5BNXe5HxUrhyXqlA29A9Sro6EUfzGjRkbfazyVz6vHSEqj
ZC+XXwDFV+zQbff0GbpzsLb30zm33U7dCDQEpr/0vFAuJrLUbAwKeetsuPLMtRTADHH1YJidvTlb
rrC0bQwaPCmTKwDLq8VqP7VggJsNPc6UVBvKfOUOh3Uau9aI+CAKWy1E8pd1LddbpZ+XO8PXDzvv
3Kb2LneqDSNDhXowE+zNxcKOJeqGo3Ifsp/0OlZRBbzLgAtLpL2PIuZDU3xjOvyiytqXK6HMKTaR
TFMu1RZ8Wy1UTwXge5u4bWWG2ZqBAb36Telq3yCoizhbd5R9Bg4TQxCXgmmZR6+WiDKU85opcUiD
HZqwYhS0slz5SWvPNEDbUv3NiCyepUvHA8NSqjUTZ/KEBGTekylNGui8HCRw8FlYinGihC7vYlXX
0gJ+bv1151u0PZTEMXMuSeZFryAFVVGFvo15t+otXE35wEljFjrUDCJ1249PXdTFI4hQ0wGfNM26
PfR5EqsqlkO+PIS5CsDGjYWfdiOWM8Eb6P45AO8yJzMR8FQQL0ZT3FZzcuqZknjSyAN601SoCQrd
P8xCmdemVuDzN4VSe/doK1WgN4aypv8+KUgEAnLicAz5eymY6WGRiJJsdu1XR2VX6RjUZkw/N3FS
Oe1SMAJmhcjWT/99J69yCyiAu+hkjEzImwbqIU06VYm8x1UpExG0V7s2sqXHRg2eHqcXGAP8k2YI
GZ5b3+CA19DGVAq+bcjBtaXpD/9cYHtuVSPI2un2zq/ShtChjHv1ZdJlOW7E+R5K4Z0ZI7d0KU+Z
Is8o0xGPn14UcJUKTxqWH2VoijggLQemezkUPRx2pUn6WQMkNWd6mDHNOkZJt6Hy6lZg1rDZeAAw
XYN0IknGXBtz0qhq71aVxFzmIZnOBSgg0Gkdu7brdq74T5z7BnteNW70LMbnK86LakjDlBwg8SjS
Pml3t8Vn/kP/XO31Ezi1IBsnxl+7h8tT1lsE1KAOu2mDy53vVLfbby/3Zy1/UfUli1usXge8yqKv
MWnLmoeSoLPEtYntNZB+XfNPUOcfUYFtNL67UbHYVgD9+2rOtB/j75kqllEyY1GxJhodIL0p6J6P
8i/xXJrFEqNQBijcSAlDAxzBzBp3QqKFxvriKBdbuFETFM4OUXQcesKkxaWtOGyO8wYGeaA8ICmD
FHrXvnROib1YQrji9OjCqzCbVD5y3b6pmGQv//+RGbb+qBNhG6EJ+5du/fhz5Ipz3AdiilqzDlT6
xy9BSxwjPy8w/b0TRj14A2eTjyAEad+PQ8GCi6lpcA4rhXxAj5rKL10MAtvYLSoBwuq/ZpUfsg8H
eBT4bKbBtDyHacJsnsmVONJTAaExvegx7TnGtdY4uhwkSsO/n5pvzYT1XIyT05ueR0v8336g+qmi
r9YT+kxnXL4LtgQP3DllK81x2CLbLHD5CF2kuVcqDD7L7QA3KYszSp3l+r1K3HuOTa3zMv+lmrU2
jbleefjNhH8LyrngFh/SyqNaY3qVk3P+Y4QQv3xwjPz6FejsdnXaTMhkt0KUv4hkipbqQf2xTM2C
M8toSAsgYNQkShiFBY8G3PJ6nkHgfbB/1g9/KvLPdVA4sz/fd0Fg2aaBIYjqoPLerz+q+RfJdr4V
P09Hjic1M5vKSlS5S9bqm5HHyEqO8pFXne90aUwDIaQdWPFkn2ZiHdhaKouEjox0psOgGsH07s3E
7eZq9+PVpApA4K5DBg7KNh8lX7vwB0oVjkIDnj3B+2o9hop+JqW0grzBCQ3/HahD4Wxh8eU0TfzM
EcAIKOYF3Z4O7BezlY/ZAW/x0qQR31LPObYMv35KrRGOwdqu6BcDffe+7cE44wSvCenTMbhwpXzB
cz0dt8EQ7ZEJfJG8i2hJ52zQzSLMP4apHL5qFnbsUsDG3JslqzRKCoY22JnSME3gtZQwY1KK4eOJ
IvIPTbVHxi2dICYzyXvRBV/B1kCGzX4TaAexoTZJ2kvGX5Uaib8conulRGNpXAZuknE3PbiW3t3l
crrpZdVVG2YeVXOQ36IQxLESauAcmMVPYmSPnv6S9pFKDarLC03EBsfXVUTMB4TpmhWLDHgX1GL0
nB5qO3QbMhJvxfxNS4GAai8uZKWx1yHO6SMNyoSFwEdeU3Jjw4WDN9QL/7kDGEUYT856o/imCxFt
7O0FQ+J4JFw2DRLuGv4K0uyxMYp0KA5tttm0VqWYguBHsKIoXQUaTx6nRUbgbbULkQPrpu/UkJfz
Xr5bAJDNwsoNdmXV1i/gpUcT1kCGjhc+3TGfcS7z9hqyFy0AYnzZjOshnA39TgSSjsTg544a7aUW
pzUaXnjQ7SlXJOakFnBOWo2HArjymQAKx+fbOJrq4ygob+qyLH15LEfXYAeCSwpOdKu0FKodGWzx
+aE/Stn4lFhfbSFHZALrIXdCOLlgzEFHRF55Jv7gC75iSGR+CrETdc2RQ7f/20pvxbJDPJ7hycah
JcNbMy+jMYTr7j8Za/0sj9bs0siiB5hn8lFT+kd1k2PpMS1GNJsG0Ee2WR26hZMPpV5hJxXasLpO
yw+MWiteMArkoQ5Q47OAZficeU3g0wmjNgSX4kPQSw7Nkdu2MRhtU3+ml0CVxzobM7EGjthlcyBN
KviMMDZ9osHnZTMX607mzQHCF1D637WAbpwNhQ08Be2kKiypFziYlNzOdbdQa6VBq8hZg660fBLC
K/8uSj0VGTB5oZtCNDBA++GEJoKzSxN+6bhGAbcT7FoqnaM1QG0YPxW3bzXoNwm3xVu+k0guAiez
cY92uAYgahtjNT4rWqExLuv0sVhwJkGDkh251FExEtkMEB3JLY9sO1/tJ6RBtocXJaJIom4PV3pe
isGWS8mhxyhRQjfWjvJqityhZqb5XzQ/ccG2pSO0PmKXwNmSms+kf2LccBOipsxMCF9xrpsYGCMA
YPtYTMihlrzPmy/gGCa6sjoGJjx5oCjVgzNrGNjQpmsah3ZsW/dNmSPcPeGoGy5LaF26zPU+Bi6x
6PWZBfwcuQ3hl+jqDavJ74uav374g7Pa1oQzMJpMER3vlh7xnj93mEon70vjVHnUqAGAYKKVKmYV
2TDNOYGvAlhq3YNRnc5Yyy+SY8f1fPeG/M/F2kSgWzal5YElQ7wAjvHoWUr7Le0zcjXpR/BdUX4w
5QJvNLlJpjidPDaB3pDR++WABN44MW8Su1aV9xzmUsL28WqnBXOC4Q2X7LCJp3xHoNNcv0UMQqB8
dxzi4rcf6nW1YITlgiBKODEnK5RVx1x915LdehfBaxw1zVPO/c6jGz2RKiSaaKugQKVepZgzkRth
sTc9x/4baeXv2o/zqD2BPuNOLAzzkRdCDiqtqRyxvrobASCmqaq/bNDNIYroJb0yPgZLKuTWjU2M
appHm6bZ4lLRsblotoXZOtUrcvIB1U1/rJhLbdtnQlQaFdefJSW9QnZ314D6/kgAPBrlisMHtfpY
3kBK1kDPImecAKBlAajJGfLQDMtbZKMFtk2sg0Be00citmqfLvhS84O+1uyqDc878rkeOh7L/6up
bekW3UTkvYee0Mn/lN51H64V9mgQRHvhOo68DBk4gBGBcJC9V1x43ERoYuHWmjyOoY8d7vMJ+pPD
LapDWIRonyKR4eGOkKn+8s3WS3/jBuHUfiLepCVfEbei99CQOYGxnM+veHybvjZiyIjh/tVFi77u
BVt7j+codO6KyLM9CllbXCw98UCBbqWqEWTdG8YPrygEOZEsck7MG5BQLqZRgoP/yKjgp2+KXAnt
j0EmGrB9paCmMriIcZ52gFDoE3uTMus2D9RKqeUwQcvCwnBQBn3mENoUmoU00yXVognkWLyrrmHm
CbhoCh4SMuIkG/2baETk/gvTFA6WwTzf/L3d/9w1BcOW++oDSbymmytLFRgGmhPbjC7Wt8eOZHcX
D+m/EpbFnrivqIdviLphXL77n/2KgUwMkMnTg9dKmcRUggAYxCM5wHYNDsTdTGeMKY5cN9iGbw1j
88sfZ5IE4O4rcsLiA8b4ygl/aV362GJa3ktvEsgQpRSZshB7FFpoe3PUvvFUaol7t1DYXzDLNFOR
o5UZ7pNWohBZvShRF3aC373JisI9pipVZiHUmfqg2sTWOT6y6iDvCVscngEDHQAkIivtpYQjlEMD
tztrqlWxbW7ttZ9TqAxkLV6yHi6KqB29vEcr3w2vMotsd+jUQ9AZ9K1d0mQXNJeyEVO1ba59FyKJ
NmY+1IExG0NzV5BR+209gSqC7rfs3reMjht6cRP/xaW9067NN9X4gdHCMitUQNUaaoq0RrlU5tGW
1AyC6/vEnKpS9aFIW+WvspW4OvLjyoAaD/wgS7jlXWU1wuaydRB9qc1R4jGQLgWfi210qLXdH0oE
x1YQSwoqf6pQay6SfF5dfNkvJc9fGlkCufn6CDbk8t9soP7bnsFbNUj8aZRspVLxxwhtdfJYwmrV
OcnqlDM32NSOwBCBQF0yuy4dHIhWfNYozKjPvFstsr6+RpC3xjuIHVSn2xl4A+lzuH+YhRqmpOQN
lDKlovg50fp4pWgFArkPp8PY1zNaMK9XAHanWTCqrvNWsbyPEcQjyo+9Ebjl8zwJyyLJqewvOi6b
xU0yRdj3+s3p6oU/PDKO+PvGPCzKNmjFNN9KRiWAdX7EI3pB/3vrtkqI0gqvW0pn3U8YY+eFXqRf
LeW5oQqH9a8yJaxLq1whDYVUV4aPeq2xPRx+ITRTa0Ly8H33gM/6rdQ9W7lbrWWWPv++W9EidKUZ
J7akcQTAnm+J0oz1AiCMKxmIqa+0t7W8pvAKPVXMkkuDRwSfT2pbGmZXA94adKwKrppFtoSRaLP1
1Pu3+DdQHkfE1iuPXAwS6pO+7Ksnfrl3yg9VjodFSZodZ6MAbgTPwgM67GdhkDVugGul6tzWzUil
4kHHo9xL/2azRYlr2OId52GWuN9Xl3j5YnNJdgQqTrkYSL/278ze6+pA2d5pBbQeZLX8/zJEbWbh
7g9gnDKVbldpwiluFxElhMyQ2i1bjrPbwN4/ufGFVZAjpA7aYWBk42Uoxf8LKTDl8QrtIOZNl1NW
w1d5Pcak90C0026mPcffSOHqTDMc9enx762X1O0IxmSM7/EdW+8EWoSw65tZFfdChv//2YujYaVT
VQr+uTmdsiZg56l6AFFNsvH0qQcYWFJX+kDidfhDlIR6zknXEvuvbCDLwGF/+trNA6oLjRMMzRzj
tJrElILtPvIGj65Y2rmt6nvBxwys6N2cc8JMc7F2v2s6mpimPOm3aImQrBUnxpEvBj/Qaa2oJcMa
3J6f88x0Dj9tUy1HOcrEqY96ZLiojtWGPr/YKtEB83IBtsM3RS9O4Rmw6Lw61VqyaWGoWgAW+L4+
dFQqgU3BHDLrh8EYpKIPNarnmPEibHh3cfg6POg7OVYto5B4aFdpujlpi49I1sKs4tcx8gCRxkYc
bZ5HVwALCzflOegeqipLqESmmLhdnNS9aubUyo8B0yYlfO1nZx3L5+vLIBrxfJynZzNSLXgqObIe
0IaSofhswM++w07Y6uqcroHPAqIcK5e92tIZPGjEd/Dhan8j1EZf0PME5FWIkrhHfB60rW9v5FUN
L0/g+SndVQ9MAsBAtP4vHk0auqPpJ5jb4SbAFoa3qOLk1UjtKHfIIhNJVIbRqDJt+9q5BOYBtGL8
JJVR+DJmTspaixTFumaT9lByj3xhhtfefl4Gkr7n9hFLzLR9GTGfDmeHqJIAl59itOdAu58zqtyX
87RvImR4TJ/GrQMtr7ciO7uFMzHTEDJ2xDQwRb7LTF86tdbgQ2uFIzskj7G2gLa+HpQIY3F8MbqD
elqFeoSASLLO2NCveazp8w6e8LME217fturCsM1kB1m+ShUZ9216NIE4sFadNTIIGmCdEmZAzHmY
6Hc6eLaDMp13PFHKXgXfmOc4F+8Erxxzaz7UHw6N+sddbdFlS0Te4tKNU52ajChWWbIId+0ZRjIQ
5GWJYvGGXplqpCCnDpBBpbT2Z2E84hxzEz5CwkGrBPcQyS8F8XnyIMQQifk66y8pLPnKGurlRtrc
rybRRqnpK6RRcAWIGfmTnlU80sIam80hwYfqw6S7qXrN68LHe+R/qMC4s5J5h589mrFHZcq7J+Kl
wpSRYnp7PurLojmGEem0rQpsLEF+3cwW2m1/4pys0bnrPTJ98U4yf4JvrbikuOJr6QW0MzLPceb7
NDU9eZmhRCZPYQm0H2q6ViFwC0rijXh+6xZvBvEpooAkHMdEhUOSITRp4yZmDTgIUnv/lFn1p/Y+
FqjYo7ZDOJZVdc5e3VO7/Vfd779tyjH+dqM+uXqQS1ra5iO7lz/4t9ryUFIVZ0Idqd7LXQu5hO6N
zk2I3N3CYn2QZtxuz7qKbVyBygexGoXqJJLLjvIkvTbKLiZj9G0R2Ke/rONAlnQoIqCUPj4/DXkJ
2h1Zkxqd2C/M4IN+t7yVcnQ1X3UbRbzv4rsnrJAxwaFsgvNPidzHuY40tQ6mZMlca3ntfMEv7FSL
JGAH2pLDe73INiflc3fSl6MCGpxKQmQhlthkMqtx4zxL/br46M5i0S/994qQzqbk9dtmBHWfh5Kw
A/o5JRCQRwZbsQgHEQkGI7n5+V8n7l/4hoO4QejtBP19Vs6pAhEQRHUrhO5S/PxOjqx6t7EL3lOy
C0WHmamQJjXt6qkVgLWW4b5U8lpnSZtKDbMt1tnpgyH7NMzL2dkSznZBVcaTt6KWeAURLRCLEtFE
qfC/osnabeasUO9gDs3ShyQPXU45/BUWzlvJe8bfhFuWuhjQ2796vSm/NqaltLRXfo8NOVh/YB8T
MtUZAqGHEViQTpeOrAOznEzH66wLZWC9KYxkPE9JjAw3BUe+5ahM/uGOnKe3HEmA1+RqxBR3cvIL
Hpnfh3pzat0qUVR6r38YXGvIaD1Lul/99wHyxmozFQ7+tNuKpXasvJdjc7kB0aoUaFhKgY/JrV7g
qOv7FjbBK8xhEvD6XgTjj8BGP4upB9Gd/I1+4Efot9ejHJy8tG337Xgnw5Mv42ujx41odfSC2Hb8
ETOaCMqw1Nea1xrg31L9ZlwGQY7dt0JLEg9CbQ4qmOXfOgws7mae53uonU1OiJtfpPplN9ei08c5
5Fb2eker+eTkWyhPLcCMnJGhCoTD23UYzFG4OWk3hAfTd/wWQCwt0oYPsW5JhTbkSpcLCypXxViK
rO1TBH2GqM0HQbTfz+SjOl0Ekiwih8WEAnw7O1/vnomkN1fKDEljkk8GzxnX4D0smX9o/E/R1O97
AIkyg4zBj2BSGT6Cy1Lq15sCZ055kXYbGeF5/WNR587v1fNTvPakKPEVngGUJxLLjH78DNv9kPPc
3/EL6Sm2cVP+JFa5IX/6wLGIyRvFoDuM7APLCk6H62nYYuzMIPXh6Uds67UzH051y2Uto/fhd58t
kCBXfM7qIolDeEVavH6L6TOc4Gv4KE6J6LPPP+IzEUQcf9w/BpcaqAohRpnljzZl3GEK7VLjccLt
szUH5XyUGUScugWIbUWvsMZ63/Tq+W8rMhy+fmZwLiys3qFNgJeivIHYJvuf1TrvVnzO4a3f0NPy
1uN4jS4NWkyPZBm2Q+O3x3kS80SF0iJWFFau+uTHOxy2ogbg9nuTK09awmCYwa86T42Cpoq/Ob3U
ZboDN+sY82/FgfxkAgXdvB2/BNbU4s5m4J560eMTJN3w5G6c5jrQXamyJHI7foAOQyhGafEOWwnV
cssFq2Q/hAtbh1kIthfVKk2+BgY9oo7wHAIeRdIDQYVcboJnpufGiLarD2a8mCHbunRmMkul3ytK
FtT6YkvOOp3ispETdh8Sml3rZQrPJlFGhp+7VWKyidvnYpsZUN7ZzW9gipgnH059lviYKaGEmHjc
4Z+YnFyFs2CMLL1M4vnp6s8PzNM2NRyudsDV1v3PnloU57WlvM6W4/pgP6qxUwbWzuV46o49D4hI
xPo/44DeVPKeO8qRSmlLwMWw7WoLN0VIUPTtXSmjdU4fNoEZ4D4UbWSi+8D57wsXzBuN9dJQcsFB
q4v7VXAmDYtCtVPFhTiIdEy92EfOMrw7i2vQ7vX9VhU6FWRqezF5JFnYUrgCwc5laS0+8cCQ6iT+
9l+rPaXnx5I2UtwB7awOzoOqUw1Dk44ELVJZ0w7uGshrd0K3SEqXDp+iWSdum+lqj481lI5aKoeT
ukuVjOTUwyP6ENNMFgjqIqzq/rdGHXwjulhcRhawQrskOJCGCepNOolplw4RhrfsHkz3qZNbPmQU
UJ4qbezm5KtWrPUeOsHud9oOvGY7XBx07+3Lb/Ojq67iBV2S9pKY2IBSHgYVVDO+8Ph95wKMNFka
u1cwQJl8CnrVSDU5nXV/68PaRJDbdZPCSvC1fjd4f0rY7jK4ScP/SxChpT1NnjVmWbzhQGdt1vW1
LE/fBP34+wCz2R2Nv4oD6rneBPt/4LOjRmPKP9Las7WWsz3uFkDV62O3clbJI3sEEDAb9XDhjR/p
iinMmhZtHyecYJ0qWMBpgZ9QVblzzKcU4JANnO6ZQAToKeMy9f0+wve34VfVDu6b9NjvTVRE2jmi
0Edmw4BXyA9Qnh/yhYHEWIxmCMY7I22QdOyrHasEX0rqyGzM75hH+rKhuMvxT46z9De8JHwSy9SW
G2CMPUdQTLsFCcuoFnGiyi6XAPoc2UICLxzP0fe/nfIQ87jkf96JhcCWpH2rad4kIityeYzpYLFL
ZKhHm1FXmFqBT8zWu1zwAYOHMYm5PYOplh5bgldwOSlieolF7hTeJqhPA5Y7JCP5myBBZq5xlEgE
8GdbiVlsJkRhx1sYy10dSETGaJ7JPFOVxWkww0rW009DrJQCDIOuViiRil41Nm/2sDAQxC/aujaB
jhJsaRhcLgCTVq1plQHMW3etR+fWRXxFWPHyi1Ev
`protect end_protected
