`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2368)
`protect data_block
JN1BO+1BH02pw6Sx5Kj1B893pV+oLB1le3+uKrXI7Q1i2REkFqWmtRwLC0+K9piDGep4zjdgr4Ue
DAXARTkVxBT/mWdBQipeywYqkXkxERXSsr46exbRsrb/Huh1sPqMeiJgLCjMaGUZBtzghUomqUnc
y8UBbcsywkuUjfY628GgvcKMrj9BFaCj4fH5GdIonOTRyT3JdQ6v/M8Bz1/1UVrCn1wmRr6rTsR8
d3I+WpTs1AFiNJCnjusju//L6hqL/bZuVJXnU2Usafnv+r4gj3kgqrXPDLncSyvp0Lqufx4vrYI2
7ZAeK8DYgOfukPTTWB1gumFGRUbtQ34AdR6IQAcTN5AWBVMRxdrZSVstNFDr7iGQYSc8cFg2y1f3
0oh0V4HLd6aZZhm8onVsVOfat6rmg2VNCAP/F7VwLgtvcqIjNVqgutbT3eZPgRsZVpo+LIJP66F5
zWwSmlNGWJfWpk8c1LdvuSC5/BY5uH7gC91c6AnSZ4j5hnxzslALpDONVAkLOx1yBr3WDsfKpDoU
ItmfBSBXe3/+m8r9iQu2fK4LYpTW2inNF2H1aUbk/79mVXEfnkuCgYx/hva+ZLuWHnEEq2Oww12V
ZPEgjAVX7uxpE9GsG/DoZtcMS6QT2Tclrnh8GI72u3GH9FR4WQtVs0o6oPgFhD28gmhEtl8wOTU2
4I5/SfK9mnIBtKr7Nq3+uxij6MlIQezHtFgM0PXxe9gCmR39W7yezhqPIGHfPro3gA5fn//+5oFD
K4LWRw8ffJ5umSguoquK32Ao+gtgPm692gepb/ZZCqtnFZ4qO5756v6sGkzwQlicRiTFwr6CDQN5
PcLm15rOgVOhM06IGeQmCpHBcow/Yn+Wk1NxVif8q0EljYjrWXDZoQ18UodH+UhvyHpCOlmNz60r
Y26HPFIFFgf/9ry/ynluZhXhwFkWdHHHCka9D164wl7BbuItlKBqoEtlr4CLkn06dl+lIDruJSe7
3zT80lanRJ3TxgENYR9gNHVvcT9TCgTbYZN6tZV9JEOWmi2cnFTmE87YCZ/Q1EpbT++N3A04PpZo
AscpQ6F0UOr98GxjZNWr2bsJGSmAgZdnToqjJaN1JgZa9iPdqCVlKww0NHXIitg01Sz8iEMfNFOy
i05X6Avh5LNrRoCtsXuW834B6bsiaXO7p1SQRTzgC019V0GF6FbrE5E6xfNuaJKmr5C4FlA0CX9w
HLH2tkEMyXjDLogvuVB7rrlGsOaoSi9khlMqFjODSscIXEkbB2gnK9A3MX0nH0XSOrKtVPMwl1KN
x3Jv8jBJI2DCmrNgdhbM3a3u6IGK1W1EAxl7E/fWAWnBtp4n5QgD8EfSiJ5SRb1FZs4ImbQ72q9P
YscXy343kQpbt2AMKIPeD73OjcgmdRm88INveS9Uj59naTza7AvrARGDDuZRbG31e1axHZARQi4M
wVm/1HVMt/H/I9FZdGtOmE9Iw1AJrGfA2oOfqrWo7cKYR4VXkHKF8IivCYJFLUD1vdhYiIzHmrWR
SO58mDNQl+tNuiHHYHEY2+g1Sg2EASs0X/Gi9uc+T9fj+QD0lh3fT7IfoRp2q+DDDvjBuikZjhsi
h+WnIk3jKjvK0k4RhWmH7ghNCNrkTarzrmO8yypNl180fYQmV3haRSEdQU8QTdL00NPLgLjVEdXp
iJZB6JJnO8AwhcLWS9a2s8j8zj4tbUPolwjTV6LDqbWdqZ8NqYsBQ7RjREyYg7rfu1LMWjL1sdpN
raSlsqcIV22qGJ3j8on9ue59OQlaoblaXwuIchEGmVoz3kGxcwaqEwcFggMmpXp6vr/MP+wJATui
ctbQJYzIk7iK9lXZywPYawz17EZiKwPtP8MENjxQ+D5jB/O9cVS+FoZZlbJhiPAhMtDgLNdN8azv
Vo4+zafSf984vhnb7xOtRvV/gfMtz2ldd7D9LpFZpvTq4hTpyyFtv9Px1EAIo6JXasml498a8kiD
8LhUCMjuLsVDecOs+1e8Aa7MKiNRYW2VFg9m8zZA7+4kDRAwwvLXFZPTWwtQ//FhHBNno8diJGa8
zzObNmvdg5lKDRLz+h6UZgOhql04pgzvAXTwlQKxvcm7y2Y2Clg1RurO4BtQg2QMoWKp4WBeGmca
lqKQ+NtzjKSeBC96HNwqAfluI8+HWfwy/hDb2ndqZt9okA7BOMs9xQGcgBb/ZVkNJHWNgeFtFS+r
HR0n1P7LoBFWTkfsgw6SaWoNwPyBgjeaHb4OtZ01R2MgFzp55fw2oe7dJ0y3aTEQo71Dnsy9pJrX
bvFU/gOUf7fOOv7fKYPlZUo1TsvVHTbQHTT61PxZ/1gh1UGvwul+kzjkLjRvrtMWxraNo7WQTkSm
cKCa7Qjk4GnaSaCw+BtFDIbDmJs8vr8J0Y+W/HpQZAhQwmOVzStw8Vz/2LEbLMAtcIbbg6KVp9Li
iZGPCYK8iYonzzQj/KiCLlRracicJxfVo7pcwYXHjo9jGRMP6DqP61gyVZWfrP4CessWZd1VqcA/
hG9XyNs4FctQEqXNiCXXvRnucoK806mQghnRxrgOWmpZj4G6xTHtDnTKTXQAco4ZApmFzO1BSnhT
VxB5n0OPizlM2VM9aPjqSgmdxKN1dXprbT31DyW0f0B4Adrrko1ztX3pD+Ys82lyKSY0lrjk4Uxi
SLqkIqk4cKyXoTLdQ4pibTDy+u+dHtS3lzzoNAT+oXlDUx/1Zq65lpuXnSEDklwNqymUEq9JxJiv
xr68oQJFZkVJ4P+mDMcFE4P1XRm7wO2RqN0jRDZAXUF+YXXShDDq/ke5szMSSpZPHxOwxOKcGtO9
kVnYsUvvD+7261XLyDAmDdXTfvn/qx2p9UHQc0nRHaYnJnPLMDtKaBQLgOh2cQju63RmJhrcVhNk
0gGX7sugKeuHi7Ruu7DIbRJA1/QmSsiqt0+XnUFvJzDvvHUlAhZDZw+B2Y/vgZ+gOOmx/Pc41VnM
5XAH25UDmKP1005Gfzr9TQuMd45Qt8bjgN2sUjFAznbegI9id1oKsHQB5s/t/TbWqvT3Sk5UhBj7
qlrbuM7e5x5Xqe7nqEjZb2t0vd4OM7c2kXkFK44520DOP/Y1Km0CLBUJ3/Jpnt6utVnWYr0O1/CL
lA7fQeXmhHP3mXrQJgFAcW8vX3J//29qfGV9X9e3tg==
`protect end_protected
