XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���M��W'	�U�7+�m�ȇ�n���I�g��a���?O���R��4a�Z���p�Bڶ����	` �ݓU�dg4v�i塧�X��#����߰�}#�SAۓU@��s�Ą}�M�#�����]��B�Jj2j��	`��\^���I��$h���@����V ��(O��n]8=�����>i�1����E��ǯ�A����0�p�0#�FJ~�&�Qp�'���2�̪/�\��DR衁����[US"L|,�4û�t��R�pT�s�!�rӎ���LL#���{���w!	']�'�̒�ouq������wI��kc$<�M��2
�XE�y2�mb�_?�)8P����>�ڼOV���I �b,�
�T�����~n.1&G�w���-��N���׸��(�o(��¤����"�1�r�<�]f!;�������p�Đ�:/Ԡ�'�n����@���yWBf��u�1�u<�l�}@|�7�E�K���bY���J6ڹ���x�@u�1,��M�F�I)��H�������$B.�F�3N�e�mX ��	�Rl�[�#�p��Ӕ�Ɉ%�T�,�zg�"�f���uȒ�Ł�����twlxO� ��D�X�K�[�_!p��G�=� t��㯵F�Ij�}*������%�l>�ur]��wأ�w'�)��v���N��
��/0Js >��e��taK�q�*�rN:��mN�fߩ/�D?���y��x��~8�y�e�w�|R�l\��{Wj_��+p��.XlxVHYEB     400     190���Qa�b?<���Ե�KP��L0Gf腊�H4�6���`r��j��nO3����Q���,�����kC�?=l���8�H�`T�'ڮ�M�Fb����_���)�����	���?�"{Q@u�0����d�`���G̿�H�!�/��Q���u�w+��1{�Q��	K_~�&�	���&`z�:�JPh3�E-�G�h��݌���A�^Xt��r��A�����M����1)��1���훬ͣC�C�g�`k�IW�[��W�F�Ѹ���QO�LU�Z	�:.�R� �I.;�Ƞ�e�K����|e��@e�y4m�\q�F�J��Ā�	�+Tx�v?rT]2f*X�Y��t��WU�b+����t��-91��Pd�(�*�~�4���}XlxVHYEB     400     170�T��������י2�Ƀ�3�ԥ��Fi�����K�mRq�.{\�q��0G���t�_��hj�a��@t�y1�4Z�y�g�V?m����pIc��	9|�@�c�ޛء��Ţ�PJ��쒭���2�uT��v:��x�9@x�ۚ���VK�y4�󸻫A_�{������Z���bAe�>\_>��ڼ�C���Ѭ��nG�כ��M,����S��k�#T�vr6pC5>j�b/C�n�mk	UZ\�������4-0���w��������	���KbIP������ծh� ��P����#@׍w_�ɡ��tb�Q��^Y�_���7�����d�i1]�UL�q�)XlxVHYEB     400     180"��b@: ��)��'�}�ۥ#]a�_^odu"�q��/���t[lHsT �ٮ��F?G�υ�\��ë�߫*�k@7�*ݬ�W��R��n��g� b>�[]m�(y�9޲�"�EL�+�認�XYzJ������ˊ�l0`+Ccxl�~�|Zķ0����)"�(N��4/�C�(�����FD��S�b� 0g��*rV|���n�6~��?y�i�����5�a
�]�iI�u0�n�͸��1�{i냘l�o��s&+��l��-���A_�J��}Ww	�W�0�l�0�ѩA���4����H��+GRp�a+ʈA�����<)jY�ӈ͠z�'�G�xn6D�C;�Λy������R���cB�\�+XlxVHYEB     400     150���g!��j�W(NZ��^�F:S���TfB� �\���}�&�>�&���0�<�-��fi�[��,3
~]LЮ>zѭ����X�LZ�f���9+?Ҹl��i�C����o����;\�O��*~�CЭ�|��3���j�1�s_�!�
�>�)��4W�[-���,�3�b�J�����]�\�b�42񴢃�*����As�Hڵƀ��|��}ne���<�V���K�scv��:��O=�;^D�M��DG���2�f�2,�(�t�K�8ȃ�6e]�6a`���Z��P��kpH�{�9br��������x���;2{��%�9�<¦��XlxVHYEB     400     170\3,C��{؈��Ǭ�X�� �#�
(�)������m�u�n��0�*/\5��%�� ��O�+F��T���#߽ ��.ˮ��( ��.�D����m�Z�őC�!�!���(����v�2?
��m��Fk�S����I�b�}��I�-�=@$�y|�Ą��7�fE�*�T���Z#Gr�5��3��/��~	@��ƹ��h1)��� n����3Ͳ���RDh`��N�h�ɼ&/ߦ!��S�`n���K�a�<��:�o��#�c@q�����ڣ	��a��C�yW��P�k��:�Ռ��E��j��[o�WJji˦�������KK�ҫ�pvN�R�(����!����	O��XlxVHYEB     400     1b0�,M��8Ǳ��ET�(t,�5���EV�!��������_i�&ĭ^��S��m�#`( $j<�+�´�]�r��è�ŉJOiZ7�e6��wƇ�γ
m>y�t�h�;��G���#��ȅϡ����>A cAR7���zx���<�h͒��P�ʅ��1W;��f�}K�Lwǡ�}�#���n�؈v�[v(��]��^6�碝����J'�9
TȨJ��c�/O��2�.@W�i`ɮk^/��,�9\����)�ך�F���o��v��k���xf|��.KϜs�^��:�1@>.FK���Wf�$s�Z��i�R��X�	�$6`F	�y����)Cf6�;�9�y������c�v3�y˨��;T�8�l����&���=���2ѫ��ut��ٔ�x�
�^o[�9� �e��^�jbXlxVHYEB      e0      a0��P�ɠ�̜�FRH�������e��y�a��-^�.��M}'}�n7hY�F�����Y�离�R���5o��.o���l���*�����Q��o�L���l^���KH�n@�{�w#�gjW%OPq���>p���~*�u/T�m�8�_M��\w�K