`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
VFkWCsf9AtbDCWngJZW8amj/w/bDCfpeRMieWgejuMOzOi+P4RApZ0vdHvAmJgPdl/pWAPF4Em52
ku5Y/A7ZJD48twBqx3UexkYMlKldKivFtE4Is/fWilAHJ6x/ItDL+iVju6Y7A5dfZukK9yCLudjF
NkvsbySSLvnIyxj0nTgFGt38hi1Hm08Qi3zbhqqC1bA+H+zwJvCHgoobnibmFyeSUK3z2c+YyO//
YheqbZ9Uee1S+xbQKVs1bSgr1jLG0zLrAiNd7AJfB/9vBiFOiiXLkOBtx3CZCNGJXw7CAfV1RAFG
8q1DNJtsTthOD4pNpIN8ygxzQZrlQgp6qZrTjw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="+FFB1V9vO103rMIaQSU4H3/KNEbLjeSnNkrTAvGZogk="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14000)
`protect data_block
olePeugB1hfL8YH1zXAVsEaOfwNV5luV/XnixeWuxavBY5fIIhWe2E7nPd6EIB29KyXjhYDwD5H+
negc5OqqgLdedTr6fKP8AXxarmEhqd3UVmPcbKlJYHC9XwnFZrcQFmytbS+m6QOHZDOR8GI7U+WT
M2dflGlXMD5Pw2vzIpLQC7US6skwP7sfrtGu46M9vWZohp+JcrjsVWXiFOQrN2yvNRQRJ8kJjcki
qE7ATPiH6v3krbfo9h99eM810knl8DauTVskWQ0SfdYoE3daLDKxbDxumqoR5OewhOrNh8YjO2Ix
mvIDpRgcRcmD2QuBTVDzF6Gipas63/yyjPq2EZRc2JbpP9sNQuFay1wWKdCrpjluKar+WPW19YZX
TxU5YsJLunH5bsKaEMLHvLwIU0f140QpSWjkS6PzQOc6ZJKCKsN1XpM83JAZ+aGzLPlFPdj6e1T6
cUfDQcYpfSucjtI45gtuPnvtOWYqJp5sjwl2A+5Wv7+qZpQuxwzLZ7vOc3T3jVfr1ampVGyHMgwX
Kbh7gKSPbaB1Gfrxv+W4JTJUcC1X0ehWW1Uw4Rt44D5NIzUFyjX/nGvGksDsAwGdQuhI0P37W/Zz
LpL9PtCPKeTSIXa6bOweic9LV3MujlQXNvpjmLbWA8WJrRuhh22MG7FldKN1mcpo+eItX89820by
pHUDQ8Iwj2mvJK+Yn++wRXYhSBMCKnNLQRxw4aPHs+xcWPWmW1/ENLw2BbrsUpcdDGkMA3REN18D
te1UlGG3snRUsbvsv3q4WWGs9mVpPW5sV8rlzHPiJsHqhKUpsIqKgZP6pl35bqyQTe6MTNkPGMOJ
zKe2lnkSMJ3s095LeKMDHzwEo34jhGFnUwYh6Ip7+HGcMG05MIGRdi87pTRzhd4DBgkU2kUWY/Li
LlksInpry38Jz0rGscDqhyF0kGxs3Uypmey7QaKcrdsXXNAzPfvsfVU3USXuMDAvSPN1ODogHSZA
OrZXoEaCF9EkNXuWAJxqW332BO+zO/5qPUbcOcbm5xNZ3aLvbCyNN2rggUCrrvVVyWX1yy8W1AO7
/CZzuiTGZlXcaJgv0IPb5NYD0SmmViME8iONqPR9/SOoT9aPz4VToDkCX1KUYVzRNSCmUyyYIF6o
w6qhmvOmwDG/3Sqr9iy+XAjyX0PWyRpHqkr2Wl6NXAkGJaWUxNn124286zF3CYX7q+NjDqQ+ToNm
dQG4QySw2FqJXhQm1uoqavnR7eu8huVvoRLHtG3VKywzGwMeg5u7bzpmNGDcFj6ObXuhQ8x+OPCL
t2vZDrLKFvvFSmVO3XgR+KlsThasvjQNExCIJc1WqRPSWqofJOOZ5bt/tDQyjGJJCMuuQx9WE+zl
Pr1erW7A+8zw6zHcZ3XzlFgxp5elfXLFYJQnjDHsUJy5H8wr9oxioI2c9OGXacWI/+m8U86P25CY
zXStC+e9m+WZAtrNuJ6m/5BgGiTmdlmyXx/bwOxGlQI1qwF82u+pxow5Aa1oizIAA2ogUFxS5aFq
rqAAyxhjpHK/f0hZsRtXImfVRjG55pM2jvGbCjhtlJ9wXgsY5U60O2d3gBkcy3/gTWwzFOUPErKT
eY2/V4BjcTvNBKjLVXKiK/3QxXt9Ns6deKFW6TN5Wi8Ys266rL1BKdcVj7efhlz9HSKuT7JJBnwS
kHd8u/vJRZgSQg22YMNETGhuFFeGKGcb4L0J/o0BIvmf5chvANzb2m3C2QanqAOiwtjMBpj+CTGE
y7/DiA7F3AaRlsWhBOhofyKXxRunZc2sPMJpeOK5sbipixm/SUl7ygUgpAkdN4Popff3ZZbFD4nv
kSBM/utCrU11tbc4sZt+BAQjka9+9pEkh/XwIwgo1qEr9ZTnQhCxah0+FFiV6iZZ54/azA5As2lB
xGPFIRD4NEwDXXgkL0h+WNx+AsGuHzjq/nIl/1VN8N8eQVFGGsFLMMfFSi0kvttFnz9jH/xlaDRi
TLPHud06E7Os7WO7o16xHQiGSD6bDiMcmiEd6yR+Qn0TgpXCp1RjJXmzfpCkaaBhK+h2LoLz4r3J
8mRou2LpKQiTTxLH+DWXMa7d5/bhBeO7cmlXXk8m3IhUUhww9hisWYAv4MIyhE8oMXwYlWgIzpsS
YbhFxHpEM6E9L1Kkrs7hrnD2GexmiPSAwa0f3G5HRUh8zynikbkuQ3T7aqdRdEwGBHatvd1nKXku
m7ve/wDzkGboWHTl+NzR+DA/3dKQJOIBoTLAumTFbsLBN8m205AHfN1tq+FDEw0rU3zmuzAPBiXl
S2uZlG6aGlOpIg+YnueqLRTd6QDxAcfZ4NlH3R2BL/UJslxR5oEKUvLD3SmDIyJwJeL1wO/VJDqu
3FuTInF3wI88/eds4chOCoiXA3ExQZMF8BuKEFbSZDpid2ENBYPuvhq/X0laVXcvrRjf2IB1u4re
JyOvSh3QNRiLitvIXo2vzy8rFXHWsUqHVAw0DvVA9lhX2O9cHiegTntvAgzKyHqxXfFIGOfDExkH
tf3/V3kGbrUKbN+g4+2yOlDL+HfWyGoa+yEwQ2pfbmNcF3HYE7cFLLI7JTCI0bcv7u9d2FpjpAmB
r7lFEpiaczDHWpVlY6GyqjT85ViX1uut3HoEud78Bi5knD32i9nVfxYyVdUoY9h2pTL7o/5hHwU4
i2ZiMDcjxhV0YTARYxboOQKi/ECoCDFoDs8h/dO/BRNAuNzv+8L9TJ6s4irk62QUrruxYNyZi4NK
v4hQHW1qHITU5j10Q6IFzMY68kG8bBQJo2UMJtAfHlrF43OJ3uBMMn/1KpPFzUxqyqm1kG7SZckk
kT50GtN2vG3CEfNaW/Aoh3lroo8cyceyVOmQdfmo1uPLfCewiHuc3tkKLILjEF8A07mrnXyyoUyF
Wyujb+m4dcWJfFNXrreOH7CEljKBb1ZkI0AQkXOMvajLncjkGVHU8JK4ZhcTKYYJQrbESLugL10N
fQWJGtaF3eL3V5naU9mvjaA7Pidz2F0gg148+rIa9K56rmzKU7qHg6nNTOpGdviHVW6n9+sRv60Z
L9/pltIYbHoqvFS2Zo44rve0xTY3hNJP0Q+99ITvhbXhY4S0Yy+xoE5kY6FbsdBsJtXeBMoEystd
DpVVL0C0JqKVlZdNka/HKnjDa9SXhMZ311m22hYsIOAwuGBbLclGY7QkQIbFva5pRaGy5m02Kmaf
fhTrZWUltjI5PcMO9ErmQa3C7yLCz4MnrUjybXcm4/t88wDmxOjgunwuRLNkesZ3rN0l7hFfAx8c
YTN3JqZkfDskvMIdp6jyDK/OjXMbGGGuIO6BMb6cFoAoTfn3F3+W6TOQdmjt/okwIzIPSMUlOjX9
Lfge4ATdxhgRlsNY3x4RibifyETcnioz0rS7Lwp3SAD1mt/2iElY0cnTcCRMVxiM3SGe5Qu+Csn7
TCVnQDmRMUCSthMupru+BD5CbpC951+ZnOuNT+u0NSi/zBSF6OmXHj//bsbnxtE9xzrSjKJ8J+Mm
sc4RINtj4KsRiewKLqKjOMsNhIoHFiLZuiTAFOYzhse3HC1dX1Z2XZ5vtKDW0CtPKphg6BBggEnc
rwAgkzw6+A0O6rl80578FCeqpio4CaNTYK36HjskwvrZZE9M0RjULNWumcfB5a/6hukKqkB0osoX
AQDtKvTlXWFBIO1cXyPTaXfB07y6PhYpWjVW1rcSkzz1dLHfEaJSTAFjSIBtK0JNSdDquZHDf3TX
1wYMMpscnp+qZI1PbIVU7+apQFWKq8WGBTMJS02FkDvpOEVUQuxh5FysTNIoYBqV3LVHt1EocaKn
pqx/CG/I12SLSawllxkrS8jyLZ0FR4vZfx0ZuOfMdw8KZAM87S3t8mj/LGD+Ois2NqBPXCOCB/ZA
6xQm9+qrt9uf0goKsQjk3HI9skahMyy44DeQBh9YnZc2rKlTgWU23BMprx47NxOsWAiSsUVbeYSO
t1ocA8c2cv+LjYfVROU3vetZLFLyXk/rcFJFEAYYI6n08udybyUQ0lY8vxPWcQDuhPBCf1lTzaLF
R6Za1Nd3jeQjPfqPgqFNMhjfSbo4S34sQBzjq6Oo/w3wXQUMD8n0/8TSEoo9gJt+Wa5IXNeExgba
xHNfVTsG/3pADB+64N9HqI71obK8tRpKIJvWcFYz7RQ6qAkshbJhpbZHCj0E9cRjTHcC6m/gkQdS
JLTqu8KfwiJB2NLHlkErCYzic7c67KsrS+X+XUDyb5FQsugWEAWxcvRYVXoLGO3l9312ygRoVJAy
PJNzMiG8t9zC3wqfvF/w3ods+E5Ru3S7qAf0nbPmB3v+mMhHEhIgewv7Un9UqHcU7+w1Yool3uRC
8Qxr15mkFHA/aMgtuvAyqHuMliu440Mp1E/Z5NMYGUczloJzc+6RQ8te+hk8Y2wYUELitl7x72o6
xgFm8oMW5uqa6Yy81mjDjNwLI4xgErl6ck54VQg3TuIE/H9xpWnhudVT5kFnB/XgPzjLkg+MDraz
HYm5pfWGFgal0SafSoH9ih7g6Z9Wt88AcLD+F8wF5RQ1WyYFaen8X1AkvpdDSJUtpGNk6KQHNw7j
JusPC3NJPdfWF3hNYWqgDPOuHrBJDXcbihk7QKQp+F+zXqRRS9aCK8FBSidjnefIPQ0yKy6EnRg3
UDGGo8kRqJGhRz+hJYY55nVFS8eC/L2qZbxAl844WOvfrhsY2WujrIYwMpanBoRb0CgdFQdNTNJB
gB4LCtmDCITA2J+ckiw1BU8j2wTwRqbbUH5s1dOx7678kP1u0DUNDvVQxOth4YxPM2T7okAzpQTU
wp5+sIPILQpcSbX6DURpcprJRBhZ1QHD4o8/bH4YMZpjO0StvRQYb8o8aW4d1glDH4++UfPVC67j
aEuOOg5m/XtDhxESDcyyqOYF3dJ6fLEbd6S5fdULNJWlVF/akvmj5AkniFnKjG5fm0y8BCwUHIxg
Tbm6uV0OfSR5CyeIgOCf0Divm+S8zSDc0qxALOKBnK3Q/Vqad4D0PgUnc8LKCm9MVeJYPV1gvhRo
DK+sT9QpO06C8xohKdnCn2lrPa1Oh0spipwL2v58q8vdW/HVNoIF5gCSBn4OKa+GfSLNaN7hHONX
mBCCycfVzvjiE34YtK79U2NEP9gTT+0Ra1J4PCS52z3JWf9dLD6jiRC9qa1MhnsIS2uLSFmDdD/s
1Ckb6WpOAtflHPOoeWQAN2JboR+Y6mzwdUjZZ4OTwt3mMMsgoKye0RwCJdidQM5nggRXV+fUwvlj
z8OYAPDnDNpFzSCTHqn0zwCHBz6PW11L58UV/rXZ5L79m8H246pZlCatQiUm9tqxtNBmPHF7ocEN
V0PLjm2X8ZN4hS22xQiJyNSRPTpI934Lt+GrEAPzQwmD8blrrChGiDImYKLsDLHprcQmwAuSB6pg
J8TbqPHR8q4Nj8c94stGib6yD/58NMfr/AlylhHW0VbTPt1tqxJ4mxY9nCFLLpwyC2W1eWSOophD
86ynWS2LsJeEGJUCAsNM0zN853qv3psNttTNyUhvuGtjnuQEv9G4JljIDDrW36Stprsm8+SUDrXi
OIFYqNTYZ34BRgPDksuX/NZT6OVBRJNVPINzCEdcJ0yooeQQ0Q1Hj2SHKd4M9gvAqiJ5oGbYV1h9
b9dqXjUcQKTjwTE1bYvMm36mCDmGr8jfQ2bzHo4zuhYMX6cAisDzsjSghsViodRzjFxqQb6YSYit
z6bBaXn9T6MxN/t5V6gj/vyAsWvaLmMDd4HWEM3QfQdpITDWl2vXy4Sy+5+E37zIF/q8NPE7BwDn
CebgO6I7GEHvhfbe1ELVdl5JlHn35Yfay8zdCF4nI0lDNtS+makEIviI+2K71D7nGx0jhTVEp5KR
w61j7TeXsBwM+jHz1cs2CE7GTTGqgTR1gG30OiY6kNlYvSL2ip6AlNV1GkXnc71nIHx/uqkZRtFi
pVlAAPCAYlxGD3Q1dtb8JZyG9fza4x/tH9aL3tr7ADzSgRHtQh8GEdItoWkULO+ojhk4efcokg3x
lGVzMzuS9S19P1NqImJ0GW80kPBHtg77YbHXIwVLD/4dKGysiF0EN7ryPZgQZ1DOTjpPoFUjfNof
KNhv7ZOrxLGB7VPc7aheVxi2vNiDeU1R9pWldw/mRiyRa30Q3CnwoxZIy3SS51lKz2TnX/Yx7xeN
geGSBpbfUIYFy7K6lCxuUJ1B4ite4G6wLWPZEA+Y9P5OOfMik1stBRFYlFrFn0LmHaNXp+5G7UU2
Hy2Vk5axgtnroGdqcWIdTwB2XSWHx8Y7WoU9/C491Eo9Ulso3sQ5DDY9XGqZsU5VbRbS9m1ZBN5C
9BsCMnEd/JVBd4ox6bslshIvy34tIxx02N9U7XMfz1Qu7fpzaD0GdVwjNed4wEBc5GAwQ+MLMX35
Q5H6QHPFNnevSmCOJENfuIKeN1TneaChov1UHS84mVXC+dVUHW1L0uax6Y+w+d48cxe973Q2a9M1
O83RZdh9xAfyurWsq643pKot1y/F0S+BKj1ZxgOrKkEPBLZ/3tjx16V7KNxHRb+RcrCLjyC+wKk6
LoJA7Q6cGt3ZeC4ssYx54NgfL01gVBQWLA2xmGd03HSCH59dpbTD39HeQHl9Ibh431fPUwuUrT0I
1Lare9DKzwPqZtUe25MjsQHf2cIAkwz+c0VnFq7llWup714dGYf2e3mHEXCj0TD4p7R7TDBmqSMv
cSUEd+j1GwgBKV+IxewDQLnnRnaKbPlvX/1uLsk6KfStvlM868w2FBkmMBhsm/GrXlBbxXfzpxto
/wTzxczLb/z3oRi31FOjonVvPedHuIa17szdVfsm8iy8JkVYf6/TH5uXB9D4yHsDg+HREzXg5hD5
fMSRZQwB7/b191uiLCpq93x44ABhYXljNElG+vg2capPaIPe02C4liuCzuY/Iwnaf2ESbOWBh2MP
4ePyTMyjpE22dzudrOEg66bgBEhNPIrAmFrQspqSHzYFMIzc1ilAlDDb26x6rATOuCt5z7wFv4AD
6+Cqn14P5UZvHZ8U7ylDMIGyqfvbBVhfOg+prevBQ4p5O2XCWLJvFe4S+H3P9SDTW9/NyBXViT5S
0CN+Q087GDXobuhKzlMKXOvNEB55svXA0w3P19ScjJcvV8eWVjfF3Khkb87BqdAFJSIyVZs9jA9q
9fPttlYxPJBya64uI5AZSQdah3YYQ0aJ+Da99rhMq7nMuaNL/lZWqJnTaQpmZOSssLB8LJGdfnjl
U6DvPGGD0T5AOfMVDL+b82Tla8/vgW7JJZjC2T9tnBRdtEOWKoojv0t6eT3MGur+Cxu8AsEkltSA
Bm6aSTtTVIVPbk4/H4xMRjt67h6EEBnGqFjCL3r+hm2jByQKTIoyGApqXDhFVijUT6mQxVu44O58
d5+LtqDpC7BQV/BrXdC44RgbXeEP3IgdhNbaFxAy5z0AVeaxNHvreFXaKalbOvNCgRRJGM4GqOEU
3i/yeAAjbr9vMKY0BilTBT7z/Qi/XZtI/qSvEEfc0zSb4e9ZUbD699PFkZ2YNh0M5yjWAcuDR5EC
SOUiZE3r8Y0wQS+ZkiGLZD803Uo+lhmsXD52JHApCZ5WPfRwm3aCmxo1wTtNEXNjVhZKV2Aze9zZ
UofUbaC8LiD53Cr+ReeprS7EsM2hV0VDnlM9QuQnjUgcgRBH4ZNZgTQN9pdw6phK0EDXN1tDuRgb
K+/uAHGaLIG/Hvvjs0dFsfwqAfO3DZVGnFfylQ7RLZPVo1BbyzJdiyXcTxUpGwPHa4fxFiRX7Xfk
naJUe7lqYK1ctixGp4OPHbw4tcpyLy/NwJ+a3bPVrD1cycMbEsWEmxeEdAvdafYs4dFx+EEcJlJR
dMa750mY2i1f3DIh5vkNoi1KMiuFDaSrCfJ9s6Z6jmOWWEX1uQe8ttLnC1NRugTzxMc6FtHGBMHm
jshbcvAKsiCvvDp8P0yigFGXCNLJp/H9q/eIU5PfDI3vHnlUphfVHCREljfZ+e5o1Gubcs2fWT0L
Xuy8klDKlz1FwGTFCwscjUCTbG732y5zmOpjpr1y6ngp2NZdBBGusQlojVkUd0l89x0EqcH1jKb5
aSHoPaYSf8W2ak+jAOjIRaB0RvELH+jxVJq2D3O91MxpEBiK7y1taVGRxYPBmbzJ1daR1jAPaZIE
ID+u1tyfE3OOHolQ8pSAaFMGs8tlzenGJ8hcP1u3oDC9XdozzpjfGtxqk2GXvn3YvzrxxlXXYIs6
1151hJlvQ8CQb0tu+ESNC99HwApM9rz/KJ25Tw9IW1shnFU58ZCo+82dIROEe0ExhQjQTZ3SpM96
qhRRPfeRd67A/X0mHz7qR6MxSZOPgQdOklZ24HMJGb7WmJ8wp/Um5V1DoBLxEoKe3VCrA2X5AFlL
/5chkNvXT3EJIO9DMljneJcWBHeDjcVWBjNwCSJl+3f/xTRpsnHuFAHAZlQCLhcjgLiYbCVq3BAG
6nO1ULZoTLfBBOgZ1oUpT9XFeBMLk8ZT4gIvhWADNqmOQpATiYJBlXYcgAFQydIqromuDC4hxSyC
XRMBhRJo3wXT/Pbc990M+RWnnKuZEv7ub9lcAAk3rsV4tHyySiQANTgeWe0ssaTqdsTiogjIpYjM
G28ON1wUEhCsoZitVwAImW4ndiQF69ATggaFO0IKOwtrpWe5GkNYY6gGq05z/6p1SprvFUSNbyGG
vamVGLAiVvW6/8wZu17IH8mRsul1OM8pnbqJJ+jjuL2UXF1H0vJUAkmvJZmuCUQwkjamWIhQ9Rcy
1KDQh9N2IbUYoubIvbw+staXN19Kdkx52J6A8WeAeI0jnQW5+1yavi7L1RnEVTZ1qtzigtDwTghr
BrNWAJsD7CWjZTWx2MK8+V3hI/2MC0QmFogOPuEOoIf+47mhDCQ4ua3wwphK6iP16BtvHDRGEoRN
EjDpL2okblyuLuH3kV/PcGAoOs92cq5dnkEzt1sIODHwg6ADPWn5ULpoNn0NMLs+TCtWfW+JX2gX
mYAxFaWOJAnfQAdVHZDlwbjvnyhR91YwL8W0MVqyW42gP8dNB1Cl/2OKfWA+yEjAc7qDwkywQyYh
FMO9uO0+3xYJhSIqAC9zujju/cvoGU1mue9+O/ZP5zNO4EglghkWEUG4AfTuK/rWvJ85wPBtyhzv
7WO6uVKgCenFUDgYvtlMObETxLWLkkQDM/a/HuwETPKb6b3b+o2UJxdB8vlP9wiEDGZu3qbuwWc6
n1icrB4oCat/DB3rYT0t5ffRMQmE8PzNkcm/kUAEnQAy8I3S4fI+ZSScRRfFTpmYYkpmHhUjtcjz
E3A6oikIdCGnPmabB4sJXxyohnJuvF/k4KKmWpYXubbJJZX4jYGWebDq+P9ZuTBivUMuQE25F12F
eKujgoQRN/9fI7LA1CVCTXHrB88iRhTo88tb7NNypBqCfA4ILW7IC7w97C/Hr8XJaB54qS6Rjio+
PU6abz+o0LyXPWS9CkGrhrFg1sNJce86j57s/WX3Mh7ItJKereWLwphbtsG0VDRdwq6TBmfdZ/e+
KDvJxOOhD9QcoNnrM/+zFf6YuBG7CjW1hdKkF2x8o/dbpqeDoYoxgYZcxh2t2/Tw63EEiCJESub1
1HCxGBf24Kg8q4fqgJCiKNvKyCRy8cZXUIYs2fgKEfyAzRRhLTXBTFpsD9mrGkBaXtPujPH154/2
YLHKs5wlrntOWQsm6mrLaSrJuQCow1wFANaJOcbZzNS1JsBakFXW4hrv596mRy5flSVwvG6+7eUi
9itC5tpjDOhgmzEtE1oHSwSYL1lumUyb3oUZx4Hug9WDNT+/bBWuB5msmOfuTy6T3PxMfJ2lC1Nv
wxIt1anlKTqj9QpGv5YZNeXwGSUTzyjTCp8x4QaSJat24FfNJH0NIAypFlgNQWnoczGFOOCJfOsM
nTHLtdwU6/Clbzl3vdITqRw38l8zlyNkyxMSnfQksrchPCh8At1un7UPnKM6Vp/9/fLJN34izV3n
Azaic5JCem3ZHX46TBZ71+nDSulHaam7qAAYNyz/rqx1qIC9ldy76UhzycgUPAhnkn8iJwiiIALf
UzaOSWo0FMcL0oQ0yx5WNZDnoeTChKh+txBt47R0c5PzH4jh0dKHkZDVHMkxL8pRoi1ViNG7xS/C
Pf15//GUHWhIhrWc86WWJN/qd4NtiQ4RqWUAPTx9Ll32FReEQdSfOw2xNqSWUZzCvMwcm0g7Rkur
gjIymlPN6cwsO6AfLd94GoXP6uAcTM/Qh9Vm4SX53yel6h9k270JWXjE8HAWiRaH83Z3Do82JJRj
PRgac+yVZSzuYGA2eVkAaRVIPTxel7Rjg0xH98+vAMrxChdGhIl26B9p3hyD+RWMIRwWjE+S2VEA
VOnGyMi4R+EL2yP1darsBj6V84O+bRYhnRnRF/9QI8uaqmw/fDpQbHvBl4FwUZvIyCR87E/+y2rg
1CXRCuJXdulCjPY1goCRx9/syT51aMLMl+cXbyycGwLfT0iswquios52RGzIfhkdoerRAsmJByfb
CDixFzKj+x6H29JtxknKybieTZrn9Re5LuBqGh5bSzTsUtenfuoDYmbndX9OHZ1BGGL1YobpLk/I
v4EIrHkjUk4SaxxKvTnmrpE7Tx5W7dJs4FeegJzYRv9Y6nMj2pfZWguuA04VLMbb2EvnCfUZcsxB
dU3xlfzmga8I22ORE5+W3Ye8bHtw+vCk8v3ZNNaLYFRj8DCBB8L4w/9E7Ea4PX4TLLMsqrAUvheh
iCIwuGInkmldXYxEJjtjH5nO5Ke7MJI87upLN49/4g1Twz2lJE25lHC8StsUYCnXwgrJOn2Xsh8Z
mypjfNUKiAG79RRYry7e3QTN3hZ/LLa4qGh3GVn4EAHQGzTzb0TZ0lBb0CTLgSmjxuz+Hrf2HTeX
8SnuIxfSWRG8N3XWjB1O5orteo7jVrzDGjXPtnZgCmIDzzH53zBL8nSiGsl4aAGBZYQNQfnrWkMu
VDYPpjwCefym2eJHtEObpLMtfm1Ah46mf57WozEJ7F2i3KQSV9sM57kZYj7Gcyhdqun5ZHxmmidt
OjQSiDxlGp+Qmjr/DlzOq7evmKYM4VK6S+DymFTk1yyEI7Cw3eJTmxkbrsGDEbaDU/41nC+suSHM
sQ9d38UKEO4NAJ5yAviQEEkrSfS5kXn/O0nA6+10hJfuaSng0vl/eQtTqlmkAqH8gyNcwcXUw46R
u5To8hBBhG/xwV1VadglF+MyBkqjMkOCHtEAN3DuEH/H+xtsODdDP6QavFvT7hIkpaIcSzvEPrYo
dy+EJombeNHWMiQeBvc7giN9Wn31qxOM6Iv4D1Lq+5Fb/nm8cwxuRZjPlAiDpYDQKt/FUv6IlWPe
hQLYD3GfxWH6W3kfrAam0wYnvid1t4O2wnRwgrIJzjI37F2XvyWSHWJ/KTCWn3hrn9rJPcZng3/Q
2dmPZQgBfB6uzuz3THcFki2AQYOAd+o66ywB6xde2o//wgr0+0Cvpwwohwl+bmbbWNowkgWaO+Gt
Gf23I90Hj8ORw4NLKP1AJNLIbdOXWovxCdeUbaWfzdpR61AUL3tLPaHyyK5GQzWY6cg7/CVHjXnN
+A6Q/SX+Pi0nILYtEXMsAZUtSxVzUUORyBY/OldH93kM+r10sLZdIoIf4ai3o4fXwueUEiTDwxg5
n6pMN9+YuRmmQcWOE4cyTjuOLWMXAvoQKLgQHq0eftgVOOs43PRpvSikwvK3Ck3FtPXz4PJUzvUR
Zof5wdWwT5BDDlS3RJapFNVtpC7/PUhUJiXmZGwdAMXHJRC6/pMJYfUaSYauLJ17XGqT6clyPjYU
nS+s7qjdp83fxKBN7qbPS1ufW121dXJV+yk7+srx2rPcAP196WWyk/F5DzhTtYZ1NCZjLaEeyncs
N883xBz7OpplKMMzuhIcEoEbc92GUOu5O9Mu21sSl8tMwidNTKpyvj/crFbbiS0QazneCUrENdmb
HxRjouSR8yMbNlcCsYQX6Un0SjQCb1jgTYEwcdhWdswcNi2+PWtFe9+ta/BMpGK4c8BPA+PrMChe
rmcb/yMJdZRsJLjQ/QxSYGWC35NVZ2oVzhnwWcB7DR28nRhZkJPz7bsRU8Fhm0P87bikldCu5vi7
IkAuJvNlku3WSb/ltD+jB/QZQuZuGpEDfKog2l5iGoaq6+4Tn/zJPyRB8EcK0nslvLq+ijs6H1zc
K4UIy9qOqNhbtg4EHtr2Vl7R1YBPjlmH4sg677LwdRkxd+iNrc1IYzQdDc405E2u9uwN/ucc/m6W
op8VPSEOE6Nmv9l+oiW+1BZ2xJFgapQtSacUl/HTs/MVVYLM3I5UILSHxbD0ToF2PElYXdvBXZ9A
CfgO4ujcFHzEe/bO8t4GhK5VPByjFvf1FOqtvLQWL8OfeZpCTGVpaI8i6RGmfVW3J12yjeNsAdXm
Xn6FRUu+VapW1Dafxbb9SmBNYrYV+Uw8PFBGHjYbqIkYUO+2k7bhASL/M8OGv0+glt5x1sxE837l
n+g0Ponvn6jxVhijgVG7sxKTHnMgb+roPioUFd3PKsEZxMpqNlurLKy/VP45Ns+wkCXGC8eKyOR0
efCKEhtx6YM6Z2rjh24pV1RTwSTCpGuR9LSp64KMvf3LGZ6cyeUA/SEJOR0fuSfeEHwNc4G54cs5
+7+bAGOdCy73nEvHahlnYHIaTi3Ezud1Eo+Dilbc3uzlQ06hNjIpHQHkQBeD9kUAyegMnH5IQ45V
/PWCvDEqWV5S0UtjYOKcr4frU9k33THh91YJBk985AkmlAl/RJkqYfcf7msV4xwkz0uWQovQ/tq5
9ouZEOkCS5P+E0tfydaR710E+J4XIM9oXuKb8DEV1tz8ApGtm0QttQrcotRQXmjl8kS8f9rkkFkl
dDvIhiVBjA3Vmls7OjV+LF4BAO/nONEEqnb64WuAdK5C9tawQI5jDaMYCUQGgGvUrDNho2xkn1Lp
5suwg9aV1Vo3gVqZNiEstLgUoVjOkjX6CYqriI6vd/2FEZAsGHHSyevZqTJId7GysI+wzR6WTNfO
28DpE5WQLhxFv5KS76dBcsGqwbCQzyLPwalAvV1a9WdRRLo+t9MNa61H+AYw1Dcf63lzI3s4XMR5
8dWV1mMCH/M2SvonMPmU++8U+LJIGGon7nsasPHkQDOXX6k+4BOUDlH7SQbvXlsiFp3tvauiqtFT
e9DsIO6qXtmp9csH0ZypKH/GCc1EZEdMwJ5657YpnzwWuA9rHZK69m3G0hsNTbcijHCgYNp1cM7m
aMUcjfy/OKRE/sDwIXj5/erf8GGGRq9DykgnE0eh0E5cyTPqnxdMrCmxkRlEgIAZwSPhRO3peKfg
KSBtAgJIs5/n9lz1WcVa+RMuQF2KUhHNRHB8yYuoXeqR1+y+/UKreM4yaMJJsYErDKZrXhiFhjcW
/y7/ynRKgE1nB2HG5kZ+rxe6tM6uYw496sb71MWHePNb6hUt11hoPWrqur4fFUqTNroa5TyU8YDS
kQJkFJoIzB1NVoTifoSdT/yq85M9aA3VA0rklUpePbCnGVXYginFKejPIB4WKMuivwofBAKQ8WCM
A36R5R2qftmm4KBwY1YeWsIkLXw/rd9775sOCxUTIXhzN+6znFdnZZLGhYsMIuRzjsoAaz4rFrPW
9m6pgQhV3xHNgmJnCngCw6Cd/ln/TjFGpjxnZqQ8gDS+uXjGGp3FjP6oDlK0spE6Js9M1uTge4wN
QlV6Rdfp4Wq0Zw5mAYz2RJVC3BOHwFadmFj3LSL28wB7N5IHLZvta/j5xPcQAZ91Yq8DUZfsO4AF
Uncd+0sKc7z5EVtUUcaMUemEd3qhYfy8Lix4USU6ZtW8Zn9sVC3FCcSq4x6FVYCd2ZmZyma1E/j5
UZU7XjFPhyRGiY15v4S6H6IoJ5soV7aipowx7hQIlVe5+OYAOCwCrIPoPFJeFzdU/B0tw+vsuF9H
k59iLCrq2kZsxddQOkzokH/uAqV04Vnj3cT78kpHII5O5nZNN6qTe0zXgSZf87GCh0RK5WmBG6DL
sswHQXCXtToOWFDjsOqIAG/bxtgLM2LkJMk0n+68x7pTH+CtvDzSHheg6zCq1DQMm8SOCcbxMzhk
7wMAPTNYjTzPXGfDRzuGe6nOK0byZLtPQnLlWq6Wk3cdcIzG0J9jSpXMDzE2bEfjAJ33PNrVRork
J6bjN1/AYH4vLFV28HxSaD+3A4z0RzS4O2BXoQ8QYypICEl/DVjxvcLqpE83AgPg0o4FAMsheBUg
xdLB98glnmxNO3FkmxGD3RQ6fjKeQTSQ4nOKd94QZJi/R/zaxeiPILPlze0k/kavwQSVoR8CGZ/1
3760O7i/O63/82CM9YUoi29VpfXh6RV+I7X36uov19iZpes18FyE/oirQTVrpJRRta+DhcEhrE/J
HiPtjkfq5V+QpBWJWO6VKDta43vLWEw7V6bx6Hz66CTxjFWfptxQuTBJOB8Zdi8NrEdtiKwQ0E5t
xOr/noMCxVaqCO/3t21GROqMS9QU7z8LkZvi4K8HaR86GELVRJzzNCItYnfW91LDMAKuU8RFyD2/
kFrgK5/3FAmgB80x6+Dz7VBZXJIImJXNk8/3Y1g4nMIZzL0gk9wGMoHNFBZgIJcg2Wx3hBVVAGJD
jfAXSZynrPp+LZB3P8AYkAIOi6MIvb1HzX3XXXl+tFS6drA2Y9BGjPIcee9zFkDiuD9eGPPnlRPF
RWGc6fTTgWxGl1RoFBN2e2ezwKUcUzZppWnpO1/tZHBjtWcykrkClKWS7bW/4YUtpK5XCCVzCVwo
VGvCQOB1gvvkLTklcHrMzTQBIFyQxE52VIo5/RIiah+Cmh3tqElMFe4yoyCkXFXdgZT7KYzO9z/h
WqbOJhVpzAZCmRBU3ACszEnFNxy9PLNRTfBOYi8HYX7WCziXxVQcWezNNVJEvOZAJ8c5r34xPhUi
wnWp3Ktzd09BTcn/wwZgER7BLZBQxA8B4MozGo8NvbFD5pfx6Rw8cRjgBNlvJ8w4aJOcZ85MltEx
0rYQcZ77aOJVIW2l/MarVEclkmq8BibEOe8bv8TLcIxznbG72W3oAu0I/gUWszkBeMnVsocIiL9h
CXAFGYJt7jpsp9bvE+/8KYOpXAzj3Qc4OT4/bOMkQieOPzYRmKcgUuJk14j7XtQsVZBJrzBH0o0S
nfM7tgcETIrsvR4RTtEbMQCZ7utIz4cqa3BpwGCvmB5+v5kFB8T7ZKDRPbwaS4lwaF0yKdUdhLqy
nbG1TcejB/ax2+RUPu3Y5UIda1R60nvOU7vUxwEg0mNlK8PI1u7rZztIiv3NtjYmnFrH48GfsIKy
3p86O6+Y9hJfhwkdquEQ0zD8gX7FhAoL0IiBJFAx1Ez5aFNmbZqytGvZ5AgsmswAVNYtWJEVSpbS
lGbQe75ayiHvnpdhdo5G+Jt2WJBtb9NB66bq9Ui/bUdZD1i59cWNC4H2bICJ7lO2ISMxOBInsVUn
LVxCLJUDNNyq9UdnDyTLRMVdRjDpBnRJW8imdj2XNYOEfFwoOe3X4FcFYI67Cb4G3Ikpaacr8XmY
qecNtgoYfxEq63b/g61EkY/nohJoToYsgTRe9HNh0fdFX01xYQmQ0+Qa6J2n2k13TtIoflt7TIFA
TYA0Fc5uooIZXvPYukFuWEmililzryCxJyv+rmc8StBulsiyaF0+1LTMuyC1UPHtEMqQyJdxDdph
6Tx2HxvAqSkNvoZRTiq0WuzA6W1OJxc1zJk86pnWg+Dl2Q3QEra423AOH+rCv/39LdcQQH12uxAy
st+GwaN/7CUslB15ncAQXOVJka/FVcZkTzRjigAwR5gfEbkTGen3LuCs3x4w7OlFMuS+GA4pGA6T
+wtH5BW48D3WaT6gRgdx0Aepis00gNXtBWkYr+yLRJwyFYzQe2RH5lGpLlc1UVYRPlcGWVOEne3M
2pfT87svYA09Axq9KiYxWdeJHeBRnGZKCvoP478ZWUXhu3I+mWVfrYuJXzmi7zInwp2L+oOJvsl5
GckHYmmhlnSmBemgr/2gZiQKKpiLzpihAjmlYDJSJiEYqTdjVsuSvnNevKRf/3FmCsOpQz5V2W8o
cJuGpfRc20YvzOslmX7Ox1IlLGnCx/jlf2kOsmCo8/RMIcElrE5YbQa8jD9C7cntcvbfZZEzacqz
3ksX16aJnzKpiJdmf2pibm/mZkwriR1qoLnhLTAUSs6SYIkvZa3DTVPYepJl8I1lenmvduE4ytB0
Wifa7d8oD6xehLxeSKaGeqdR83Vfnh1ULPz8dmNKxed7DgRpObD0ddwHU9guw5c4N+eYPP0rpGa5
5RSl8i42KCuNVeRGW3BcnxN4IOy5QLUrykGNslMlzgb5E7t5u83fXuQPCQnhqiUn8M5pfyklxnkp
Pb12Ad7tqQJzKOUqSqTBf8QuM8V/qw62hzwFvrJpJ5at1tm3TQQhMnVmXyfCzivt+0HuV96GdUs5
Uuyd2ko+3uWYapt/ZtPYBxSMKrfMe7EhHIiE29ZriVokVi2rIxwBTooZGIegFhUTVi+9Dj9IMUhn
vSz7NCu6EEoVCTkpPObXD8GSCll8+0KfVtd//eO/0ABviuZSNICM77bHjxGB7NlS3r5QIQPwpXKA
wK9WRPM9o/E+TyfrXG5C43BjvEKQuV9d08JwaM1uj3qOVMfHvEJqcxF2wtaGrZM3nHPE1vOcf5kZ
KvuORLEc6Kkz/BXCCISpJp9grUinhLmTmyw9uaG6KHxJi64fCfCNel7/dBOzqm5KA5Rn6hbbIFcn
Zd57zgktiRND0+W2BbrEN70L6cjk7hAE3+GkBx0mQFipZgwQwTmOp7T3vbGJuF8LQM5tBqps/TQj
hzQiuotMMEy4lO3Ifa+uycSLAWuD3J7dYrxv69oVtWqygny3NnsrvG8mdk/tYvkcWaK0rT6TFCKy
ij7WbsJuIFEo8UJPWHPXYyapIPDzn86FVAFle85ZptxqngSRsGd28u3pavQ+84OozA8edRO3oLH3
6r69z43oTwp/0IFyh25sCESSLtEeDvlAESJXybIQky0sXMka12U20FCyDRBeUg0wkqNGZ2ZR7d2r
+R7+kXNpBZMqT9s4zPexHVarKDg1Qyse5XXfNjpQ9mtWjF6XX0TGlO1V5clX/NNiCbB9SOrdajXG
0URwAnRi9LXR3U4IYQEHG+pupthU++xtZRPwn8saS5K6OCy11AfxOARQkaV17/L+p24euoYRQ3fE
XmPQb6iRLL9J3MIbhCNdy9KxIZ2XU+fk9NxjsFUIjFXP3Vtz5mV6msUDHbSWrrROGnKEfgEUgecU
nzeYmu/Xg+943q9Lp3maX9UQfghpFHLtpMYF0Wh9i0yGv9JD4aBZnyeS2r4GyJ2Tc/ci0bFc9Rss
fQ/2oe9hpI85aDsFDruq72863I9srEgWWlIPzbrDwcFbzKW8OJYbJ2TfPl/SHSI4YoC663VT7in8
Xnkz2UQc+JVm8K4fMUGiOKRTeke1/w6BdaavQ3cSPo63RrJMFoMuzxcpu8M9+F6Nj5ifNjTNaOGO
azRKn6O6Ax9x4qDspicqsVV+wS5+6/i1g54gWIPuMcfKgen/so4WzuE5GmmyaZw3YHzFKj71qOiG
dKPIppUKXd/a/OB/RRIwix2VbYrwckhgUwkq4i0XyNeWfbQW7iSSZZ5xguPJS4n5vFJaP4LBXKvf
Pd2vYEwGc186GI/JNg7dlhZTjWnnLQLTbX42xvjm4MKEXuPPQMEZpKS47wbMhn1bJ+/whicK2y0D
nEhW3LIaV1Ghz8dzif77UrffemJOZnyyWmVrVYQDu6JQMhwsoh1DbU916QdRrcajT8qYnyTdzj/E
SHHrwRHBsjYZALZjMp+Qe+EXxgGgxmK65go0rau7estLVF9+0vRSsWDuleZH5S10gjYtogB9nnBY
2h2PJxFpwCS7/tJpIaPTnxA4vR5k00KWJ/7sacranfD/RoP3f1h78qBOrEtpXEYFNU/5EwlzGi31
lDLL6+g8hqwrtaOUQVC4gBdPePN0eCaEo5nNiqULVhQTzG6DDJ3bn/JaL1+j2KCkgTah3o0/llT+
oTfrHa2yQ9M9k7cYEpvyGN3RqjYc6xnhRTx1RccAnUCDmJLivANKtujwT+4PKBgUgnDcSuYha14N
XarlG+aWP9qmR/dJlLSVmH9DSAi4X21lv1QzL/U5PV8On382UHGC/56rsyvlhH2oqBVbRtIh53pG
ULWZ+rXffQIhCq5owyRExVIBxSSuzyP32Y7GXXW7kUBSuZVIqW0zXuiQtFuR3EAOJaKMgxDqQ0Na
2E2xzTnxqr23hQSB/DN7Wkljj5Np1H8m0AeuapCO7O0qJEUsT66UWhTIHqBKICMQLA5Vy33FF1As
oeQ8LMba/FuTETCS/IUQck3aWz3gih7IDhbp8teHr7i0ifQBufcAaklWFHxx9baxGnqQd9oxRQPj
CkTWoccsSA8KlU1URjLrRzvT1v26pKINNpFww0FSIjdRXUXDjyGHYmk1NUZg/rVwCt0EEaXUItLF
sRA2327f9jFT6E6pwrK83zD6QXQ8QeqlFpbhjOx3yszZ1fltjJKGGar+iNwukhTrhCeo4xE16vdk
/hiL8qssUI5mdOaniW480xRGaOqBDRxLBb27tSo3xFkTWV1u0ih3ixeU+wOf9EyqjcxzhTTCD176
+V23tPgtudJ8DOn6fysARnPQf321gFt7ZeNTCqkYVGYmrdA=
`protect end_protected
