`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3840)
`protect data_block
ovAvGiXpawidI+nRnPMSjfoGO8D+bkbJmSdZbjixgQ0FP50+kV70+BtDghRceNNrIIHKrDes4qeC
eGGE4mnz8qau405Covgo9KGXmYO7S1IW3ibgsvOW36cgxYQ4/69dw+Ru1D/CY11TpQm0kn8uvY77
25jG+4UtcgzOdaWnbZosSI/6WG3S9Qw0+nJ+w0DchKKdVEUZoFMU9AC9c8TXGxKOAJTPVzIroeCv
9HyiIzkrMb7/rThAC92jO7fW8rg1rexnNIwYDY9GXRCOEm3Z8OZ29z57TF/HI2i2PWXufNrNFqcJ
Mnzt6G3TSWID4etS0t/BnTM0WI9YRL8fb13FxjA0/DCAxRMM1GCsXEGp4DaNm1wtKVALr3egsw5a
eGVfmpzZ6mnmuvWSj8WMrKQVhSPhZ70v1eOWjHFCPuDCBkUMkU53eOP1jZUJJrgURVOjZv3ehFjD
NK5yELXAfoQS2mPlaWVcPOj7aipPdAm55uWBYzqnq0HWwxndvgS6YYU3QZhoGOlUt82HE2uUJ1hq
SDPioO8bhsev2oHQc24uQTeRjLfybCh5rRXK632ZvFRQGINiEaZxjLbDv0oMYAiZqaFugu9BQ4oV
5pHY9KCTvRnhabErDQXzfNMkzaLez2gzEj0ej8l7MrbLY8ZjYy0k3RlqP2VLmRzrVFsd4n/RiTcW
K6driQUusoky+MvALGAjFU5g/0X1ISvPa36vqnn4z16uGA1+ZvzmKvUa0wgDMYWI/aivGqBMGitQ
7g0IIy6LP41cMPxw/S73llkax4vHxw0kHJIVBnal75MFQTVSWxy/XTJOVzaCzWwYF6qC3B4vXpc6
C8ehBD9acscdEM2OFB5A8GrtC/UH8/1lv/ilrTYoAnP5JNY+qq74bp7i1U6Cv+6f5a5CxPD4sAE7
9fop9DKAPR5Dqx0E6OSW6fOsUkureNvBzcHp29Sx7eBZAamIe0LD2WK8i2ydEdtNWKjOiOq7WHSi
D3yFoCAm/L4OhvZRyD15H1dU3UZeb2i+x7km2+QPpObT+LyN+jnq2BcU3D5nZude7Co0703xTbRw
5gF4lPhWflLkuxh6koVUT07H9GUvFshUak6XTj7XJVSbje5iBd5BFb7sH6QDMuicYQxTeJj9naCJ
ZktomVDS63/1zygsBRr/mbEXLR5UNaeZ+3W8hpnu/0mirPMgmGAEvMaFf0gfUKi32FchCZK5D06v
+cGpc0juhjBsPVoDo1qQysv3pJbwgzpWv9xtfzo2shINlp+tzJiIj0E56cbbB5KMwcvWQU9M30jT
wNiGhFjsLKEcRk34FzdK2E9TP2jvZmmhMLHieuh2gh+beqhB7B+piuj/oO6vECvzrsUztaqTsS/G
+06dBbHfMDD83P/jIeyXpM94nH3k5P4jnlCRujE2YCwC4d6DWUSccXmV9bwXC4E2VSYfgeScfINK
e7YU/rS1q+/82KtTqZjUROSKRAXV68Mq8t3AxmZCua0r8xcX5731qKSdx9hNRlRvxEQUnHPgynrc
m3qwSRpl0IKzU0ky8bKqtJ6+Vu5lundeLj2kZbwayJdhidzggytx/Y4sdGzflnKdTvjkWJQGvNwq
bH6uub0pS3Sdcr4UAzldQ5mxjzVtih+SI9+XfCN+SAHgBDVEGYMYwmdwbNrt16KXTAWweDlsfnW+
1ife1eob1ku6icLr18oB4GlOW95lsjdr2y/1gbhwPuoT5o9eNlz8LwmoRxlX1kta2Pm9LYiW8REY
WWiIcH1TzwLKb7RqPUe1sk09HSf9aVyiBNkKuAjtmKHioG29bTYZLzpYdpQM9QUDV2yA/GfPOZ+K
oSMyr6HuAGJ0uE1nXjuDkNdbCLQKwtvuY4cFAGag+1QtmAyuwjTOn4eMTWa09kC2HldL8t1DmVv7
X0vmDK2Cy/bbURuJxAmd2dNfJ0z+4U+fAM55o7064Be+Z+7GBVcBVBnHU0KwIod8yKEQbcPAS3zX
Zy4Im8w2iBpaAqD69IRmILkiFyVXLvKemtwkvUkvamXGzlOxy9MJRCQYqPaANetN0evXQt2U9ONu
96Z/Yng6pta9uH7VvSL8CKd11GGxRatQjU3yDCtckfS3pplKtJB0oFC5T7DVLiuQ9i7y1vrKGUZf
G9WxPjQrW444by7A2P1EHdHuqS3FuUWWqYgFh3kOPs7Ig9cjUTDJLVhqziBECqHniKJI25f02ail
eaVW00ybkRmHUWNbgBMiEqeWt3iwsgbE629kQFpHeazc+ju50+jGjMRBKA6RlmzsnJMMVan6+h/B
+Ylt3ALUOFvCF+7ISBP31AzCkUd7n6165sHRWrfy42lMGSmLqq2gYRVTnIoUD227jDxsVnuudHAE
MZBxQP5BG+u/dV5jDM5wRhNmMdXS3qKU3/RDuAIXnCMBJ+/G1Yfe03A3BdLPromZ30MH3h6xVO5v
kaMUWSa+IOYL4VcWJtS5Crvr/3eMcwt2NrvfY1dyf0B5cs4p1LDMDrfqzovUk4d1NgbPzNkPtfqF
a3kBKEcgk6IW7OvZmF38tdU0TNcU6+rTKAWfR4Zzr0wqlPcaJAhgmS2RB2287p+ddH/k+H3Sqswq
AnmMzsjGQ3YkGM8f7OwxE//hE0XyACUvCFPDe+gZRnmhce2tMXzCK2xKEs5G7QNjBjOifgH+j9es
AaxVDv0g5wCHohf6D6PGso2dDHn1pEsqUbZmu38UNF5vsinBzdRvrP3TIwfD5FzdUypz3gr30FN1
tXafvz4/rqIrSxMmefBo2DTkmxcBlDJXCtTmdUizHtJ5X/7B3eK+gtKV9CNXE4Q9z9wXGlBVptT/
JE72jup83JhU65ApsJYs4Wx+JLYshGS6meh9AFKorYDUn3f6sR/1ISgqP1DYz/bSrSCkiUIHadXo
PGHTOYZn2rzdXH3twDfaXLSUir5e2iNGAcqXxss1A9mNSymozJmeTsM9cvmRtP/bWV0Sp2kHPVNn
ndjGcW5/7mrkzNFP2fu5UfIkWh0YQe3jtjDz0D3XeNxm9FOI4ZENXtA+aDFd7y/YXgIck6RPs4xm
2s7FakxvhskcBYOOQUQhoND+xzw6TBx1AH+RxXGLVpu2vh5dpQ3rmAqAElyRcHrOtsUcFr59EzoR
yl/QscpMdd8R09U8Eg/EiQ9rv20RsRwxKhYfQRxPATo7v+r+Ia/DP0P6IN/mkHR2EZRvDtcobhva
uttYzhNcPap3vQoHuh2JJ4EU6SJ/n72EvqMrraRGRiKJDNFHf/FZ95xtH3FzUEsyW0iqXhcmDar/
n6Sl2842HzD4vZCheFZ97UVs2m/PQGWoIHnHALfgRVqOy6u/8+MVl7T7y7yVg1YbkT4t5LK/VtzE
HJF61AoFGL2By+dq3nuB6Kr3un8S/9GnU6q6xMcRBt/kkpYjH+yEnTprBxG598TKnyF/Mm7JHdCV
x/Ok5LdSOhFMM4fTfw8Ku2jaUa+jRtdukhzCPTAhXoc+3nh1idipo+LdaUYNYY3K9U/8V+mcHeRM
Fbeh+UhNTiPvkPe+OqwA5PJ+1pwgQQtpc/st3lfkyCLJL7nREx2fl1Hd66bfZCr8FYP42EN9y1LJ
WTFVUoKBWPcPig2JCm3Zc2JFT6/MF2SCdCRWJnMqm6eh0OI+ALiSqD/oeeNN6EZEE1nc/DESUnWc
m+/lI7FsUlj4+cnmwo4mhOyFUguQZ+qEdSFU84+1hUHg0XzMll4gFhMKCaJ6PUIKyM3ecT5Evm0M
KempYBcvqygXzTJ0s4/y/QP5ZxmEh9iwjVzC51vJ/rLO3WwFLV6sJqk5CYMumBj0jk8MhkQWRGLl
F5DlilokfD9fTVX+OPVQeIFm1P5Ldc7dXAZSO2dUaxOoy1mA1uZWzM/c6W3hKAWDp6ytbGlMPuyt
nudSEdwV2DHHP+JbYnf4d38/MM+c/O91sj0GuxsL/Qy98C9JqYfWbNxjsw10BTPcevHiJosFUNUa
4pUirsPSlAJCGLWk/uxblwxSTNV2tg+P4hJvp2vuWibe++U2wjdyj5kGUaa8j/yn60ePQSJ95/5R
7wCTTrMHaZ3cNtkNksEoBrsLw1pyYCF8YSJuvXB01Np3h7xNuL3wi/P058jIm3eQ2OX3OKkW63dA
eglMmWJmI0gJ6+W/VPbGFIQTGWWKELRtBD+ReVPuDt077O+F6wuiaQYK6CLPeKEXAvKjs1Xe8Rli
/wzr9veE53DEX/Ty73bfkrY2nQuSQ0+yIXcngQuQzeBzhdVS3Hc1oJJLbI0YeE0cBnTqpulyxX7m
GK7m2YMPOsRSBCq5Q8/u64eM1IE+a691sGtYVePChpjvJmLhHK4jBI48G/wPWQUQWhf79K1GGoxc
nkCnCFewVLzAV8OsuXo2gicjMy3uUuvwlBjgbSaTb0bF2jlAR5RPL+jnyXt914BcuHxFlR3xhqyT
at59wmzPTyv8pJYDTiO5CmeGUzduXQPZSXwhbY6E+XlVkHyzYVtWx+XPowQNIIwloUhExBID0Grb
Ld2shxdaNDzG4gxVbnkrsVZj90qEah9BoMjw+fhUfQiEKUx0a67sq9EKlqIkHNevKEArta4Q2Bcp
wUCq8FmBe8fPgV8ONhPfguGc5jD/dMncp2V18meO0IDe3WJtRsPv8K+jdtcu2+x/OaCiahtPp+4T
4oR6YX5jL00P+s6CW4HN30PLeo6udlSaw5/SRrb7InJj63KNqSWLokBTCdVau59vlRyrxsniQZKx
uxBXWIneCLpePrrBZYMugwTkdcWCvGtYuCDX1dIKxNE8P8XQ0jqwQgD6JbZvA+uR5aTNdgxnVgSa
QSCumV7mLQI4lEJLRHou/ZrnRqvnTo0AQggwwU8feyRu35+A/plFA6uXvCF2+lw6V1d1UD7oMOJT
9WVkLJN9mBfE0mQEuRLnTbkeUsiPSQjXPVo9M923jwzXlzr5AzFVUwGCJZ37rOnXMtGsBOU70AKo
1jU7QgEvI64E9LzmBSlYJgtAddLLWv5dTg3oRfHa8pj8dVv7UPvofc8ObLjyGk+gkkCArXJZJaZN
Udlfht/KUqp9B1JjRGG/Kkgm7PGoZC/5NLaC4LIf+UgYegZYK/e7tgkRkIoMSDQdqGJxgseO0EGl
JdtYN8CIx18Blr4Yy7IFt7FzyEcS
`protect end_protected
