`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25216)
`protect data_block
0USWSUGxovGsyBJteYpEoW8W02FbNrJXo9hkt3JsuKpm7ILQ+HgaYr9HqI/0RRMAsAKoMjbRuVsG
6yRqnXuFpMLLudu/ukrTS5X1Vb3snZO4Yrj4IJprdvzh1HKPqH8GQKZ+u+P6tG8Z7pDX/BpYVU24
NeZ4PVvjTeiCowSXfRqUsYefLW7nr83nDgpcgT+dIMii9iYXs95/1j8UYj10F0gnWaCN7OnsJeCX
9ThIBfxmDmWdoVyTgLxMZarAetNfbUexqq2e4qoP33AL4ayyDW20C3o6ybfK6rSreWDEIeFyAaMN
BSXfGIZkPa72c4h0a0PlwRV4zJ33iUkzqmf3Oso5RCkK5SLxTU5tW9xQKPBiCFDtnVBWe59bqkaY
qQODNywbw/oI07FTFSTlHdzq2yaTHmpv0zA75H52nshReNtYXXdPY5jb5145W5s8KPPudSCfmt0Q
m/eeQqzrAhyC4d4fgDW91kKA52afiQi4lENbguYn75r1PQ4sDeEpjE5TC1aFddZHLfKRYAPUpobX
kG8SSDstd+LxDmnlrtpbNQ3vdF0I4I8pbrb8evejP9tnsSK4xb/MYkrII1rFjayp8ci1JQ0gsLTR
LBmfeWC32EyaYomNG4dsZOMMVyiFFPHQtOICqxzQa3Fh/kXKFX/DKuB8TYJejJqaF66lXp0r1BZ0
etAJ0KesykgF3suqOZWuuYHgbMB8T3UZIY0uvu1eacaPEGwZIkHQCD/DnFZsPhe0/bha+3kCO7lb
LR2XWA5twP+lK2wvUgAefA/FXbx6WPXMiDI0gggBWaJXq/5gB2ENRimcmdBtMXF86Ntj4NcVsoEx
ZK6hOM94ZQrc/sRcqUzmDKfQCUXhe2XAaLSJCAXe7m38zv45EsuBj4iRyGahn5YEOFxVCK54K54i
iPbBrqV4Fgv68NAlFFQA4D05Y7QctWK9jlIYcEmJgFVSfCRZpqB5+qsMEeHuIjVkkHHBAluEOO+X
+OEl115oMuW/jX+86xZGmNRgKwedofwHsSvAAP1OyGyMbCT2jAZ7T/0iCauCKLqJKrHHCG57Uru+
Gj0vgDr4HxYmEMOdOvJlEY4YNiZ3MaV1Lb4HBde/x9oQ/AcFrT9EO+YvzuqZn1MoHrluAyFRLqiy
FqNGqx/pBBkbWP1ntpe3M5JSry12LkvzQ8TMSt3uEIgem5fayFDVLT2ITHdgOKTIU2EPQPlTEpIa
zd7KSSUV0pZNRz+9ivwiF8ItqgQvNkJfcriNQdmojfZH1MJbyTn2ZD6RDiNR+qekq4+E+4BRlLbf
FFcOlFqEQ31Cj+u6p5jxK8OWGADmf5bBgigC/f1eh0Dhk0IjzH731fgQmYvxn3d4d1l0T4Ueldq7
WFj918ML9XneFqCr7KeyWmx1u6zV+Gp89/nobVs26IaGHxhS/k4bnTFbrNeEqX9Qz4g0yWGsfk2r
Ry0Nmuc6kId4qYeQrPmwuFz1jK32eDOLByHhJNvmra6esx4LKHGcNOCAO5KGT35U6mWs3wGCeS67
TyzYiMO0kPDsPNR7no1zEj6ZXJBhN2pQg4YN5Kgu/ejcFwupZPxecBibb9YS8XJh6oTGMTyEh2nW
kl/Erv6RvtdYbfnG2QHdbrlu2sRpdA9AS+2teGcy9b5VgKjx1GaUnL+rIeWdEoVQvdQ5wjVvi0Dn
4hBsi5K1quDoygkQhIjL3UP4aH4XyFQ2gtT3TbT7UtjibejFGgLPBsGD03hAVX0f+6YSUTZ5gXzy
cpQfGB7x5zlTNK3Qg/SI7E2nKciAHvnZY3ksUXxMAgfo8XGw2o5uIuR1/Dh+r72CvQAnZeonzam0
LnkSk5kIZP1/+DyUKK3Mw5ybQON73G5Rg3iiorGJ5FjeJRkLZLUytU2iXtarr98tP2i5YcOTXcSR
1HvpK8qqGN140gc0er0vO1Li6kYUpsvON7BpxEtMtA7MH0+5so2lXVJQ5lFuOWisAD+aSMnIRGX1
yCARc0jaHM5LqConEqqIasgnRHegvzHZb8VwlJQ6wviGiEX7OjnYLWNvZXClb6RgXrY1MMTsuYz5
AqiO/1r8jwFjZJD57u1v4N+NE9dZuuTm+s1VP9qQVz68q+5EDtO/xp0yEBr3K8JVZNkXfJZJyAxm
XCP+3kR9aGJbPkvUgNRTY+HlUIQQGCdNrjiASDuBTiaYE5DukefDIEBLthBWa5PwNpNktnN1kTrJ
ystYEB809Dnk3ZBGllzV/++v9TTiRkisTRSKz1CAFG9WXf0wOB4gbLIXAVmVc1xgDCkTQ34z6pST
pWIIEfWLWOsV1Z/6cXMownEHYSFKaX3tyZO0YQSTlllPB4uepaWje/T2EWMuEmqT2hqHkqbbIU0u
bbbMoF6H38viY7sMKnPVETdsot9oRmlO5BkIy49EbW37WWtV1T1CK7NuJWKhNyTTeql3WZ4J2Dvy
F3oArMTk1lFRxmJTjz31+0C2Dr3ItwP1Q+d3QIKCZsB6e0eWa/IGpO81Ag+NnRHDOFVg4QcGmwvW
UNlGAZ9LTqJyH7CZ36eu1TLW9WKEAqXkJvf671dqfUgg3bxklRTyAIt8g1yQ3GcqrtjrPuLungw0
0qqq7aCXHuvBE0lgFo/EOfvh0EtA8xnTcMD2loVUmZ0AcUp4hCeVnEHK/I2D3r3PLlaCvDB3znou
1NpfrwPy4FVT8cMYLdJpzrPvvmpooe8fHYxJO49XV4Yvqmk4OyAn6MDF0ZHOxSE3SLvEyINka1/p
t4+i/ndOfh8MtNgO1QU7EyUJhobAeXYEwsJTfR6oaAnHjW9vfag/uTm83jp1d+i+nhad7Xi2x9g9
GD81Kol4fB2C2qqHx3tO7zvzLnnPEy+QX1Tdi8EdvOtTtFdxxl9Z1bp+hPhq1CeZeLiRgsP1kGRB
IH8kaY6jVM4SLskRBln9C9Lt7HOj2qiotYAW8km0P7DHPEJ50LYgEfAiI8lDaYaaeIM7DGOZ93FE
PSeq1nksYrzR3F3J5GNFx0F3DfRt18NKbxarVmCH4yc4gJPP/ZZHLzTPyH9Udw5I0nGfUHkSimwZ
YSkHd1Btp6wXmuKSRiZqDjJkULN/okMKv9vKDYtHDGTAa3mCtafPBMXi+o5Rc8gpUeNG/K0sAnpo
Aqn4lCFVh1lt4pLrpzwXR+SIUCoJZdlVjQm8DdiTX9wPx3mhLIl6aiUYPH2F2sbB0JW2DgAoUTot
c4HhVZPGUrttfKb9YNKo2m8igvXdYEK+PbupFH8L2Sc8puj8wBOXgmhbVUCEkppB2qDBzDi84Nbq
J9XK0tMzWbj8aB+sqwI8BL9h8M4GZJ1Kxu7Ah5rj9VNgUCVFggVVmFRNttgLIitb1NFznk8MlQQd
GDLSn1ooaEntLZXA8L5lT+0Ce6aBowUu+Ebe2bw/IvcT3cLCz/pLu8VGTBtQcfyIzEIlKpuQs5mU
/azw7lLpwoRpuGoW1kUdmXXRXRze+ttA9V9BHV3CEbZveUa8dnjfTfPrijlnHUUoQqXSKWP5Hq4M
ECgij3MyD5u/7ocSFOgyBFnFlpTO5+yZ9+jJjNIPEng0jCAhpjQ5Ps6X0CjxZOktfGji6BT+CDIK
cZHEFsyW6uX3GiczuDcflOqL9oxuG7XDef1oneIUSzMo3PWfRfuJ/Fflsgkd0hjlycuBhfGwOrMd
Qk2USyKBft1aCbIzYDE7dv7iU5tNs1u1/kHSrkER5dCzWHHBJDeicK1uJ2/fC40XEaYhVBoL1i5m
jwWXjnbg9X0S7WAeYvcig4fi5JQ0gkZtBgwQQuMMyVBpCdD9LeMPVuuF2CC7m5xYLXphlaLlcIPk
3k7Q6RUU+fTfUTSv8apq6Ka3WG09OL40+uq2V8P5vHClHCxjkBXTMrxS7Et1FNYTrXCigp/hvBqM
yyVrpQfcJayQN36YYfo17O7x3fYBEYN6KrqNJrXKWZNpjL5BFkcUzE4QRE1vVFcf/uKnTe9YhJeu
i7fheajGouC7Z2ENYZ1rgVBLOGkCpk6VcNTYHDWempp+rfl4MdKC2LTjIAUQa29X8IL5yO5/Xi7W
mFt6bGXPvUuapMPNm0mv9WIGTmb70C+vrVUiAbrvFJlloJMGyIehV6MkQK8A3+j2diCTtVdR0vdO
+u7i+GwSaGXIFOhwUvLw6z1OuL7J69kqGhL+RE06v1NPAbOZ6pxBJi6FcBQWwb4rWEJjdBa4rdn3
8qTJww0j1KpzG75sR0O/odyQuzm23rj/LTi7AB85tBXzLa7AYw9km2R+wvG4y9p/4HGGbvCGCIQK
dLDq4h7vuyRpbxs7NyOJi8kARYWNll8O3b9H6uJJkmnGp9r8oR3Msr16uV7DkdMaR3u2s8Elqmb5
U2he2X/WtUMut99Q55gBfQ7/mtYLJVMbaVDbI7rcRMd4cuatU9/g0wHGur4XiDJxtOb+U73wRCiu
WYWPGJPpi2lKgAKwaAwpwKWEMbm/JiNFj+M1LVEStFw1Vm2zkCXhA5dDHEx6AsIgcM5K+NG1/ffy
kqD4IdMpFQvliE+aUNYwTVExtC2AF5giZ5M+Ox3tytLTmTfuV+A0vPd/TezJrj0M4am+4KEUhW0U
259ByE6K8R+AXtysO1ApgBBXZI8xJYwrlnaqnkDwhPPAh0mQn1zOL5MuQ9E4DwBPjC7ZP3vvl9pi
Wz/80Ixo23mVo0ifjzgpvwO0BX/FExqc3kelqlHXCMSx7iI82xVCSZPT2PzZuDAUx1xqsr+Z2vN5
5AmddUGc5emC8vgode5NlGGGlhszsHJ18vQ/s7Q2jh6maG8+BwXed0WDduR3VVt/1JzalnlvkiVs
hwEhRwTyjSCujGZ9K7qPYKHo4ck7XYhu09lrk+KmH7xp7lhWJ3H6g9D5NYT7moHFt4ej43dfui3B
4Mmt0a/KJyyvoUttZ88kHo4kjA8NCq5PpCUGUhzAqRgaFejTjz1vBCGqcoWpdykYNTvrqK36+Qk3
Occ5owJARjaWzBjkwOBQ4lp3o3DkTeKhfspIaQk632DBQdJKm22vqhMQ03p1TxgaNTaOqvv2uwTM
xnrIfLAv7d+VjlGpfv17VUfV4Y52XdoJmjCA7yFVrKfEEF3FFc4a8RoOMPCKyCqvwUmXvIg8ZAi8
OvlgV/w2suIMHdDJV0ls1wybkmbaRXdW0MUlF88rmxcAT7eCNdv77ooHrzgRtPhZeJGK2Gkxjn3p
lEnSdWLSrfddcUeDa+/c2QRHagVKbWCNyEen+rq8ZB46z+L3+KgR3rcjMcMTID3tBBUKhh/xMq4k
jSYVfCjvWLal+jZzKkSylU4r2mhRY+zXJkOeiDO7DOCXTBGSE+LiAAB5mCcSL4lEb3lLXYvburgl
/1//Y/Jp03qvhe+sv/iHSwBY0K1BdtoydzJCvOi/KYs8t5xM3UXWuKbxa+HaTtTmDm2cgEr6MokJ
kg8ApM/pFiCHdno7gsGOSCkVYD0GPuSgczASJ6P+3ZmF7PQPODZ7lUBg+NRTVkh3QlrfvDNwKwpX
Jx9900SO9/X5Ew/xfO4ur+b2Vk5+Xm8hDjvCPwT6FbckHy8US74aiGcbrKx3tWA6bhLX901lG3ZL
gyw8qhW5YJjPaUuZ08DsdspSy5qd85gvvMFh5rRGFgIoXsRsdAUfmaaHyDaTYaS/6lmSBts982RW
dRhC29MO0BdZCZcd31QNztS5IMwhFrrkTEBJ9G+Wk7OqnD3X4GKjVmsJqubG847X0c5XSdVepKE5
U2NYYIwOMXM1rh2N3ZEkehlTyUbCvsK3vx2LDU6WDsb+ao80ipIfL0+4lKz+R+JJgv4tOw5kUgn1
nAbty+c33gUHdX8JOQtv/rMJ4+I2g5jCsA10L4QmlpZR1jqQD37u1zb50SNkwJfYwjCEVSJyA5nL
jr2hKsIPT2q2uu3o1//yFhJHkb4NReUPe+lRmtQM2EP0NWILpTxQtmH5h1zBiOZh8EQLzTXwKxcq
pmzBdkGhvldpQbyLj/3APXEdDVFuAnCYpT5dZkjCuuYDF0emJSyjUw7hJLTkmLiN9UkvazGjU2MS
usz00cJ53wVXzNGZZrg33TP2bBkWGLALhotudqMA3q/s9ZsnVOFW7THhJgNvQjRs99C7GG9YrO7B
qYQX2vnUivve/7THj1eskTi2l6z3/LIkMpr+AV62gEXbHgE7Bdbuprx1b3FKXH+dODZtZucCmJxs
OquxeVzqskE35koatb1CX9g2yF5RSnL7ebyRsi2kkPwLLrvKmYCgOireUmzyKYAIrevyyE5avR9C
7UiIl6jR9GyGDRzjJSFuSY31evRW6s8vBnehw2ABMR8v0H5VR5maBrxBlovqDzihPPU/sXmtRquk
dS6G7tgk2olgQ79Lhep9UI97XhjLsvclA+lXbmhUr0i9VjrVZ+brS/fYvDaxZPwmJKbmrEe6Tz/O
0SgMCTZuBHsIxK16LyujiUGvrL1ajUH+ixzmK7Z+mMgEQaj27Uy9u7rkqN+M6xiv/mwyxY1QdMPZ
mxgRMFotaECAlba9bK3ykXOnDA891LoFk2X6TJbNzsz+Crr83Tsv8XPTZ2GSD/DicfVxCitA9RZH
tZHfi0jw/FXTA+YvmGzA3m+mmoya5jzqskx8R2XV3Q4GeBqx+4okCWiFyW60laKiQVFNflif1LNg
BDrA+gWxgsQfaRF8CIDLr/cXkZhrKUahhRQbbGGGikfgecVVtPQM2EcsEbT8qVEhvg0Nr4xPucy+
SrbwMrp3xv8x0q9cc6swy4YNQtZaU/MV2umSU/H5SZXzzczDlxAg9jSNIpSediNMxtc6GYdEIIbX
/GdGoufNcAcngJAvjQWorVrWrlLNzFqZeKhivy+yznNZ5CfSZkxFczjN1wRQAsyHdygeYyeOqm0c
/aVqIf8w+c5ih2STpWMCqsduk1odYbTp+8/41XrPdruQ0ayhIoASr7u6riUiWJPCs4r4xm7M/ead
R7o5TKJ0Rane4GkgVtWfaAASC/bKYofuJvsadlOYDQFP+ZDOLteSDKSswoCs2V+ux+6Ia84PUoJi
S4b6gBr2lycHkg5g1MCwx6RSy1IEsme8AUSy+nxi04HnkZGlTxMBqk4pK9jtwrhEbhXxRlGSolbp
fRBDIacOJS0mQT0gGXOdhGQZvaVpFbw5WE1SNVUSB9lxTbH+13iHfJIU5EMsQ6ecxI4JPZnoHTAr
i5b94Xbe6mKcVvXp+8GMZFjgs4DYcgCwNUDZ9QgZSIzXKBKM3yJArUUu4hmsYcDuhquRsWhUI205
vNS8PGiTJAAXSpL4d2NWBJBaOaQzPCzIqgvYYa+gyY57rgM2r4pUfxZqwfC9waxRaS+90c2C0ZUD
wwBp6djd5N+e6yy7804kNuxEOfbXE12J7CI9gUIOPyavC7SLaYI9TrtWnjFmdOJTX4ICyVB1qAWv
1CU4GM5YDz5NhV/JnilNJWP2Ax6DzRTEwn70prvcW3dLKvuUPFF2aHB0jQI/Qpuy/G8LE7CTS4YY
EHVnIFv86uUZ3LslRo6SGM8LLtWEHMb1YKU1ZY8NFrzOwciHasX9GdK401L5vkyze6k4aJ4cwzua
YpEXkYOVJTx0B1NP2K2Oc2pp8sK45UhvD4OT4C6TWqN715SOdYgCg5JnOMtwxun18x9jDdS6vfq4
ofPQdOPR/p73kDkKI2lDSZ3y1S4syYSjBGilxTiTQJU5LYEPBclqVravVj9q08ULKHgHKFpetvLE
JZN6cXqHCM0/Y5FzASzTAndBeKVp8P/sf1NmE6s26/3jZXUHl+i1M2UnDCTyKH3OGVnsdKuToFzE
5jDfUHUgl0O+tsUP+gl9yvouC1tYecZ5Opq+nYi6e2XPZVtOCHGxWT39375cGTiq4uwyiD/fARWt
HawHf9vJtri3i6SFoyXBF+08EhWXrxTmtmixo6vvqH/X4tj0uWJhAQBwGlZTLwiSe9Gq66/NVDjX
VOiDIS4xF5JveRhlyoJEo+evxKxJDebjnwsFqKsaJ0Ryj7LFHpCRtYFsOB+pURP6Smg8BDhhgOqS
/kFfqEUkLc8KSNVLkfRN4a3sO9+Iu7Qn0oVQ8bQfFacO29nbAUUaPnqfDEADrT3hWZPy3Boq/HFB
ZNo4AO106DXHMmz7IuejeyZm05oW2vav8/x4DVZH7jll9DQzrh3IOIhkA901ndbl+Y7qMHFo9IwT
Sxj6EM/2y1FaE+pLQVU/WEaPePFAam2Wa1Aw/QQ21mbhkrG/Y6C5G6s6fJ+rVeoAtGTWFcgGL9Kb
oHqDgA2z01rg14MNXa9u7eK8wt1mjx6G8ZsF4NiyJIFehpSzy1gOgiLHuy+HAzYA2NyzFPnVPesh
c0vm0gzjM2x8mlc56q41Y2g6ag7zBX3eb63H9mCk6tEi3SQlIuRDNPHglSWUFnb+5lRSrpiUygUE
CPswIxaTqX1xmJnzlznydYMYnYKzxeYqWQZYtGarsiP3IeoJIhCf5twmhFJoZCYNe5XPD201d5PU
VoLlOU8Q0kbfNk7Y/aL4gnkS5GDAYw2ZkTVB/8yBFjQNrZQSnE4OVb/J2OWJTqc8X8eVJP3tSp31
Qa79yzsIMnjwP90t+1UvzfMYAbKJ9qXmRH/4sFdDxOrLZG9QryU6S6aMe6HtHqTZ22IcLQDDRvDE
oBUp+B1cOiSNznyBelmkF27Lscgz/LzVoNqrDxXV1VHUAz0edp7l8rcNwpqisgwxVFX8UtoQETJ/
e3L/X+ByaiG0slHDQ+1DcuTGgSBtwxWLW/yMZb9e/yt81GKbCeYCT95e6bkl+JHYexNn/sMnJcsr
gp+Sn3KLKqKClG+DiiKE9jpmV3juaVtYzn3Q172SMpkIXPz2xwRK4798o3EcrH8tvEBRC9hgscTT
XGf9utQ7Gwmu6ucyOW+epG1xKVzLiLVltR3wXW41gLCD3gmj/z8TMv5V60Z/LKqWufudbm8uFlyV
vR8z/MU1CdWoD/g38H31LAE2Mbreq4o3dYb/YA6pZCwSsPCjmkRcDfnEEZXG/NE+Zoft0g6Nmzms
88l03sxYgX3G8THHyES85fFg8Qm8knBp85fNVw/66dx4oumV7yEcW9jU8c1Q1Uq8RjxorgYlfPsP
F1b2jJ8iPaQMhLWtl6K7vkQhcXaeyOH5Cu0qpFn1I7Z/Ns2IX+34VEP4j33CzacO6emv2UfGoMCs
FANcunxfj2aIdyNuxQcO4I+LzXm5zUVWfNl9ghqb9nW1lojH1rEFGlpq70g4HOAleuBMWwPFTuBx
hX8XrQYv06wbWaYVfUrrJ9ZFmfM0+vp49fu5uLrBUMsh170wQ5VQfyQFqmYzKBXbstLBng3gaxDb
GlYvHh12glhA2TqN00AhenzNjTgN5uqiYugMp5SAFSLgywnlEQ4sllcuivK3joNH3KFE5LyiP4Cw
Y9B+vz4YgsPeUokePmg8+v/tq/sZ0+y3OMyGF3IlwSwaNK065VLZEjvHhzkvetMqasJxxwWI+E9k
S9PL+sTyTzfn1Wkhb8tw5o1hNlKYaqfBdFHA2mYsYEqHpJc2qTyShMpRt8tWfyH323BgfQWG/ANq
YEnSDUFwsKlAKbXeishjDPEQWWnsQM2apD7ZTwjrxgfP5p7dUS08D/UqW0+LsEtsH5jkXs0W8ThS
al4zqNzjG7A5oyJ2HvQrq0dwSQeCHIeXkFtS/q+Bh4HdhnePCmylpJgRC8U4LhY6ZWQL1aXmtudG
yFPh54TXRlqxmqOXkQgD7DCnZE+Mmpl/P6QEl8iGVIJ7qzdi0jL7cjZGxUshS8FCJ/Lr0Vwzx3gg
nqKVldRqgoRr4hhZ6bK/xzmXgu6dRNnTPADViC42Rbnz8TRh/eRWLtMpwB5T+8dTrZSyEUrp1Tic
ZCJ8w2uAjSPEU3kBbc/8MHAo0BUrv+mwCfFPAFvr6g3XkOJogj5/mYY9S8DNHIZZmKb7QAVsFD1Q
FPttCQHsz+YglfV+TybQsIw4v/5zW88u0O2lJhOIjzpN8B5Mky4TmOeF4JfTZLAcMtsYf9kPEX2K
L2DGahjbxrFrvMenLWeVB8b7GUyMcknKywB3S9l584bivJTVuGN6c10MHqjZfMl2enLjoh1i2eyf
3USe4pSQQjn9sjgjQVAh7Stb9nt+Y0+Ywfjg4Ctxky4p74HnEr1oMMwkB4YnSFtMsOlWf0DA6eSZ
IODp96rMVuU5YqORlAQjw9sHZu1+CEyor/Y9OxID4yipSufh0v13SMAJJxBVsbl0qPPrNj2Fml9O
+NuWJ5caIj7/BUNNTMWkbxbCB2Ri+Grcpp61X4j/RRzbrCKZqCZs3STl77lK2ClMGgD6/Gqz1BGm
IGfrPHZ9YJsObmgeyX/wLyu2AJKis+Y4vzqqHEb7ZrUyGn4E3wU538GQ07TCadGK2O9zbiU+boOY
b42mNbx0y1JOWAx3EFheBdHTlR2GiR9/7AS7kEcwL3go+e+kWKX9gE0mz7M+bD7WbgEX1YIc78+A
jFoFjRrHxUaHkDhZfSEjKAmsb+Vz0bsh+nU2+ldYCFDuAUw6RolIDc1+ebF5BC/F0VJRM0oe+HMg
IYDMzxQI8floAoAwSDVVH3Do+OY4lDniGgpC5Kq37V3v/LYshaVoaLolHoTHMx/s6+9vuIt5V2zC
Dn27mj+mmLF3ibCC4+BjGwVKJSMJobZReltAXR1wj5j7j35opLlVI+lAzd/B1nQyZwRYyaWzsFX2
kokRR4spfghmTjVaJhg6/YanlNZSW9JBiPvO24UBHnw581lXxUEYfR8nXMG64UUwgRuYHycFXfbC
78miGVLONMw55t+/3I8rU9EoXfdAZqB0twMecNLlEWw/yGh0Ihr6sXbf8Ge0Q0UNnfVhHXMtwUnH
Qkk/aAmSxfVCJcI3jJANrZr+4eyE4/Lf6W89DN6WqOeqhO4tze9cbEJJahHzE+5Z0FL7znt+Tk2Z
8104jmP/opFC4iMCKrtnW5qFFeCxgeNjxQmXFNE7GuFuOMQqqpqKProbsnQuzl2tJM+kKC+V5jsI
dHYSUK1PiLQL4prD72Fa2hyA406riuOw8GKr2qDziU06iY+MgZKkBKfkuCZDzt+HddNlIed3HRr+
QT0iTLNkvJ9+zI/bLAIODxqgo+A3PiKW+5rB7LJ+8UMoDQlLpMN7F8uB4oZthxlTvRN2aKVQA0jy
qPt72OK0RXMnPGm46PdEiNx/fSeCAfye82vvon5gH0KTjYCG/rtahRK6stobChjXNoxm+N59mlHf
3jb37sfHz9LG5DAadCSawDbQhsVPk5rLV1ZblglU8snz6IheNY2cH2CJ5irqhDcL20mNLLpAvsOn
InoEEOXby5Z1U35LRcykZvzdixEle6R5EozI/MydSH9seOLfd/vb5zS4pc3B9V76T264dfQ7835R
cTaa57STQrQP9maDcqMk7MrvD1vIg3eiXJq/1G3dL0HqBRxthOSrEm24kZKxoNaiK7/6Fmk0YxqL
QXsPf08JQlykXYWanUUZ65zuDwseJlYyQqXl9NKdjYRtTjg/mi6VS74IAkLCx4ssBYDL+abd8ODd
Y22nhio96d7fRZ1FviuYRRytBhTnrbziA5ZlI9VRFdQch/BLrvkzh3VWpIMA1RKfev2dwiMWubVe
Ga9g9IlFNCfnVfOGJjKtu4lYHuzzVTVvZ7WnzXTPbhvDcJBBU4MVPuRvCsvLkP8/zQCnT9GgjAXf
iMNildj3fu71W0I4kg44y+r4Ba8q/TF/MNF0GiBzKR37Z81dIVDc0uHTpIadwn5qo50WcIN3ZraF
Q/nGfklyT0EW2/3EFDE+CrL6xLCSHwt8ebIwLhgzGehpojq8OEGMGZqH3K+QXFurIOgOYoRsPk5Z
ew/IHGDJHzOTiWX81NbI6/I4DLJRcpOLHjVBT0kQaJMyS8f2Mgu8H657CggUoxTShPdvDkkBFbR4
KVpzzno1TY+W0lqRhzRRXY6wBrL9d4vDWieHy1mhZ2dSIuHDb+iJWKkyW10sp+94igkW/6jtMDAn
mRQMdpK37wqa9P+/GbRMQPFTHu+HMgfUkUpw7HBYxaPID9jvbcHTIGAQjRWK41ggyqia8isJfXMi
C1BLsJmBX9MXckYYWwdutyJCErkUGOnmayfufZpTSbRu/sF8R6J5cT4R2sArxnoJVJQQ6so34P3i
Qsu8w+OxV8Xe4Qi7doFppBnBYlsSHZxCDIkpLDIEpAmbz57whXSRlrBuGJZLDacNouVRamMJMvrK
hSXRQdS2pDgTKtTa4ds8zc5JN/mn/hrzSD9ohIoCiFp8wChU54Wo/OWsIWK125OcEVF86wjWXNNU
ECjNCGQYqCwpS46NrEMIVlpcHrXXCZDQPjmHcbxAky2uddH3h11Jq2itHjs6XBIrl1lbWmvns4yz
kvldfsWQ4UbxBGyisBzEvKUtwEFdSYA9g1qk0+i9+UrOokTEEa83LxVDshBa0wiByykuPx/fdPle
/QmpGM2S0MZPcu5cfOxRP4OYcRmB1biEWup2VB3ZSiaKFsUOXE/PpGZFN5B+t+t4TTHzDWibidje
AABzKcew7L3l6Qy4Nipz17T1+KMFqfeZXlu2NqD3MhDSIRr/L5ns4misloRMf3nR0UUlS7KmgWSb
pO3Poq/XbJ26/LDoqCfgMw5lT3vfWHEdao40mj3BqUEYgRT/UfTBQct2fUCcZR73pdxHJXGUWwGw
DF934EJf0utl0XAkmtxZ0k8o0qpYpdxa5w/Ju34eHwAOlmBhIwJsg4NsHxQeJKzwYlGwJFrFOUKg
a71ROfdb7UkZSEMxPhrawUjMRT+VmK4Cq7F5zG4Wyebzma/2yoHHrOav2pjCMccWy5FU1NBR1HTg
AcKXJXpaTxvk8g+gKHjt3OsjaGbaqsLmZrPLLaeYVhgPK7mlQSW4TyWS4HK1XcthOScL8nnFhfTG
7BTbLhBkiiiJK4MHG99ZnD0efa/KCFJnO9iNTd2GOJFM9MIEf5ie4t1Uy5AT/mm1tAFnzrIxRAsQ
w+N6JbvQlQWx1rVi9HhOCzpGxUfD5B0wXRdfl46fEaymS6ngNIDlKKqFENBRUayG/87t7gg1+C2Q
BKkQUOg9A2Y4VRfIZwfsoLFoli+JDIeqGEXLO0uSGpsx021DL+rB/u5AeDG79RGv0sbbKr4uctjF
5eFf3EOvfJIGRJVNESrl4xbuFsT0qx8gRkkVg/O7B//cHjJxpRKrY/Ud7n9ygfJL8R8ky7mklo0U
rNNdQQvaLKYWMNoakOQB4lwphsXcSthbOKcuBTKXUi4q9sQL8wPoy+doYMoPu1I5FNxVhKebkiMD
8ohMSfXXKyRtdfuJnaOwErOTyvmwr6+j9txSDa1GSGB5MfiOQIgHjLAbc9hgxdt9JleJHDyMUtF7
CfJsp6IK/Pn+30Yth2e4tegb5pMS3q4jW0vDOISYH5sEzpNqdihXrOFGeMBDIOWEaakLYBMePVmk
8i5xAPyhFGtFsR6FYTtGwDDwQVACGxrnHyHqn5VdZF4IFHBdxvw2fuov3lW8yBfnaqRzE7zlYhtI
J7fCdVkIGDkV/FyFDv/MI4QNjUTJ0x3F9m7QdutDo3E74bDfNcSXyeC9uv9DbofXnkmhvgpjT8W1
ukiLDqJYOkpw2wxSM3jAzD4RGGzg9pzfO76yoHGq6lNU4ggG0Bq3RpyRauiRjXFmeB1H3+jyVaWW
zcPglPBCNghAlA9GoLYovy7w0ZNGQeR+XwZORaFOoI4KCqyKf4VCk6HuxNBjbgAC8L5sYmjOiUda
k5wsMKRHwCtsjf+W26pzEVCDBSZfLa6eeyxlpYp/F51Gg08hqZhb9OXqANUXCE1VKghw0J6ru3kn
x6pvekfu/QcGsMUsPUTnyiPS2uyziDfMnl1862A3D74TkX/OQKno19US08maZuxyIJd0j97hHUX+
T89DAyf9bnP5D9+/rf07ovC5jtkyNWLtlgnmlAOcGBn09bI5XHT7NTqQH9nn0fG0s1Ue0uTmveXk
KtCXCGsKbJNYITNxQuunGC7IMzi96v4bJoyuUYygyJBU62cQgZEzyoLrB3YdCMJCNtXw0TEB3rnS
9MAdGDrtXCmYD3L0rMz6XaQUfpkoqZzsChXdfkAMmL/Os6IFXWtK43Yko+G+61yA4gIDneRROzt6
3FUykKy9zsja5I/hXo2vu4H2UQyLWD59q9b5IkhxCTam0bt947gZECvUaBqhV8EmFOkPJQW7OyDC
zpuUBZi3LC2jXJXmr6vbsQargTGGKWDtTgvFgl5hgNjHjCC7VZNFUZYHkApATFEAHIF1tnEMqHBP
POR0Y0H+jn9R/mhb3zg5fRBW7vrLtDHp8RfE3E/oFD1t13+Y+KE2g0i7a+ehwTnNh1GgeEzNGyhx
+mtheEyGuzbtUV4WuiFZ6v7f8h/pCYN5bWvEzuWW1SikIiCc7AESsgI1Uz34vr3DmZl+cuKDlwHC
ITuiTQl1J0VMSUEiZqEBsR5bMaeVOiTctFXk4XG3uo8eIuAsgYvSw5mnptfJst/TlqOqTycJvmBF
+uQS5KVGIAlHCufsr2OKKzm0iR6ugj95CTRmvcazNiZPuCWhcnYbu4Vzp855IZuj7eRMbR7QBEzm
KCVr9ieb3FR5iEc9rFs28kJz2OCVHTkuMV69KIRk3GuXWl6R3jZn+ocpMZjhZyH2+/LgbRH4Wrae
ltswiDy25I2rZO5pG/GhTj6t65cyoKTjcd4NxYIGdQnj12wczxWRW/XVrVWfYHtI7JB62cTnJqDi
LRPxjEImAgr0y5rL8TwjOB5DtQZ/xA7mqz7YgkZlmmkyY65K2piwMUXH0oM2HFAVlFuul7JfOgGq
7rZdeG37/H6MWOO3RHtLmWkJWLTewaw3xQxKvDtTjfr5ahlvK/C+APyaIsOZVRtDHIMPyT3oX8Cv
1ZcP/THWiIKANvLowtasK4co7kOL3pCXDDQJfSIQR1/fGkLgYlr5VpObDkm6StJJxfuMhzdWDsd6
I+q1xXJ23enoEalldG2TTu9uw+jlZUlcuN45L9wbi6aVkJnOlNv5lGXx9fxAr3YgPBu0ejltor2t
n57wBGFCAXjWeWOPWVXEJXjKOmRqDTbC/lPwruxWHbNNbDAy2rhjmqjXPdfcPxs5a6vDvNJcMol2
N0XZoTyg5ocwImxLDmFWfHEMoatsngSULAHTypIltREWfi+31HOvSXo6C7qKPG/tZJtrX63MMeRI
bm3LaetHl1kTI+1ZisqegfybB4nnghmH/ozpQehB6Zp8Wkhg3kQIWhbQOGbg1lBwpav5Aw3nB5Aj
Pjd+1JXh/dXNb1wx4CJOdnx6S1aYqzQvp/sliwKjEtjVnoikhmu/Ng6wzVXBOKzNurnfnkMFYWRI
FnJxKb73inuXBMLQMfzT0h452eaHuNSmlvIqnHFyTVKXQPa+Z84idCEjstsOz28LM8O74nsh0lUv
lpnsXcqy6rGnYbWUbeyzu8t4JMgvZZOFBevdtbw1MFrknwfItfnlOFM5StkX1D6tVrwVDN0M2zvM
uXyW15O3APXOpslgeDdUHTpuyiEWbE4BYN4rA67EShz7ME0HtPViw3DqLPicWhqAmPYI0X9QjLa7
OqrUiX8nKKIdAo78ePkcI9rwLUdKYPhfCs5q7ZQ322DoidrKRZTCvTRU3Js9TgRsjztDOo1HazYi
vlnydqC3GGOMDgRdCmlgSedpy1FS6rPK5PBwh7AS86kIXpUztx42XIto8auDRqWuK+XOIvn+CXhC
QEmEwjbcuJxYDyEIdIMRXai5afK/kwfIg7TPOj2I44pn9eF5ur6ZOl6FV9IjniMZHsjbg/XZvsLs
6mnlDCfefKvTMU9VWjckeh2+NXaGSi5ezOv4s5mUSrXvExHMDxZSPTWOTUamvxxdOnBvWUfLPfES
OPKBhUQJmygNbwQLRAFpW6Payn7GFcAyDo6IO4Eq16REK4+mnulYXTc4dI7kHaR/XtLsBattTUDV
41O1wPDGsg7FjwTE1gJUY3Ri1vjHCQTZhj2cULmdizydZmHS6p1mghfOdaHsUGFkS3yl9Kq0WSVc
klLaoVLciQqXeM5XL6pefcdVCI5bkXjdGUabvetMTWSgg+RVd6g6Aqy9iVX/n688My8qvlmEU86i
op9PTU69lYIiIF+4RMhYBAbsNir9GwdZP+Of+PlQB/JwzHMdNYwt86/9dmS01PBzZvKsB673U+SN
L2mh+AePaNMY9PYXkhk0PWTgRrVELXAr3RJTY5sAKzl0mTv37Z+cFww1XwsLlkDGq93OiXNBJiiN
Ie6m8B7K68BXgGk6L5wlLIrE7EzuPEipBxJPfBdUrNENInyFl2eCoQYzngS6ymbWQGakCWgDK4I/
jg3BpmGs7YVxU/8lSGXTlSRW6FBF1GVEia1GHHhDaueGVqBnz6K1j5uCSPpUFcvKiFbSTJetZcx1
jfAkT+s6mD6vAZ97IS6G0GYBINtUyq97DK7PYTzCuZr3D8p++Ek6iVLghS/tjVeJq3vbJKCrMgOk
U8715vlrIs4SsZL0z8QIyWXF9eKz10k9qVJL1KADD2XK1GxTub8Y3GbTh2eiWPo4aXAgJPk643ab
CACtmfp2gtlCWycGelnaR/qjyYXCt+eOXTfhMJ4e7tusdN6+FidoYIYau/uurr/+TgCHHYIc1PFD
imGTdNvuqSiIN5JkLy6gIKJGceJgA4WQ/iEP2+3ZwhhRDxw3LFZVXKatfXRjM2yX283jBUOtjsTJ
bLIlyAxTzmUNxoXUDA28mO4qUgZPPbbT2trnL3GHR/oaNMCIXTvLpyaGt6TxRlhhZa8vgujvu6IT
39b6cvXei/hzwoHZ8kh2X7T4c+4cyt/9Aqk6rFjvcu5LxZB7UvfWBSdncGTqUIiFmxaGP2Gqw7h/
Dc5ukZfFMIo2NPLZ9C1/wEuUCAoMno/2hXa9c4KU62DSWte+g6UXMGI9isiZ1doMb5Z+lsHAQnZX
qGQFNTnz8LlPmZbm5PS5jPkOHHIA0Le3dWeultTackpiL1n0d2E8stuaWYmiMGqQ5E4qM9/b2DsZ
YLU8ZL6if+D3w9RkV5Pn+ggQme0v2kJyyyiFDh3fTXVU/xVKf9qdVxSssl7tXIIB4ibAKNpfWIn/
5c6NgrxNA7cXn20S7A6Y6aWKLkLtNsSVkE+kI8JSokKnTJA5tpYFJIOjxc/vzOCh6WoSDNjNuh2h
aUjoC+r6lOFH+CcyJ4zNFO0PVYt+RQrc3I6sEinuUi33yFX105NLqZkDBgJdQnD+3fF7kIWXzAJp
vBrSaY6BVc9sUvwnIKazxO4PzOo+8Gf0vzkclyITOx5++2X1gxIoNjozdJHkzrbQ1Gv1rx9QBPrG
+29JZ+I5dEAof/ca+7Hl2guCpLJ5qY/vVL+/Ua49c/Rqk7hBFpOMZghv6BPy8Atq9Tqrr/A7ce0J
XFvrCm2cnipneFAOqRZivQtKr8ennRJjDBU73i2bC6H9BcTZy5wod3vlawxkBqJDzocES8F22otr
PSN656b3e7/a0+UyfDMVnu4svyJvDv9KwOi62cnZ/QBqjqIOPRxd/MFpDX4S7aBMboUZloL+6g+b
6ENwvQPTbbzhW6MLD3f0AddMqT3Pm0cPvtIOfWHPC/vN4CQnOWf5UmCbAAfPtO2yd43Sjv+cpzRt
iCsaaDq2HBJ06Utrcq8E1HaM3clFrmTnKIwxWOd0FWTLwCVnsWxn+7L/YQhPZ9UcxdwulYVGim10
XGDB/kCiHmLk46rErS24qoEaG0okXlpy9k7qJFHBn3o20wcl3wmWcCGofTyJKUBZatX4eVJPKfnc
5sj231Ec5oByZsZAg3OGXTf5D8MVfyTDq78d6/hnFXioFM/m1slqa7vNyQYxQfrnbvuJMqlMOWdk
y1zbLwNSP+tPstunMCz78g7nwuSebh/j/NMnlzqARRJFXLETO+JuWrFaO9anACJ8JHi7LP4fnaQj
yz3Jhv5Ma5zTvUZHdNQ+G/smxuWRr8yuHUsnywfqfCrMVkYmBc/0Nt37VKIDQ5bWVMZ5kMCRNZcI
XvtrrnAiQo20aMsBqdrN9KyGeQs2nYJlA3kkqDA/oybWBc1/QrtT82fspIVNlpUsNdZkfEHspEEz
WX4z9b32w2A+M64eIq1UPNLgrJGAVMkmWTNXLC0P8oioepW/ChbAEUq7rRPVRdS+7/NK7skQSyZD
hxwA5SRb2Z2GbLEjhzcgmpYcBwbTC9SLPrFqXCtkB+kUaf6aQzOY+1Kz1/afFrhutIZ1M5ibOEOI
Sx+caR2qvB+l8ArMgFUYCjK5aBM76yd4uNajJIg/UqbXYgyza5T2ELCJ8Hshpk+JidUv1F2tm4tj
6IA4gN7vLV1NeGQtXqhnoG2xj1o+RR5MDXIa3M+0Gs+I2n6Hhcv5FIb6TRBhsJwmuDE12/+o2qtY
MfjYwsrYcWhVJ5Gzpd7AowWNzZq2RZAM9RP5w+Or54MZiQtsoS9lXA/n4dtMeKPznI8oc7U9+Hsg
cYxY9Gb0bZcwBWgjjBvZLi+6D3TrNE+LpigZ9WCIdHwd2rgZfdgGWbD5L/jxSM0p2yLWxr0TrH2k
+A6lwyomNMHI2lycKsn0C9T/a6V/l4MW1KWB7NGMzZjeUxRoUJvDdBwnUWOHstyydI8fUMoPQfXv
qZZCvkkpSSQmDMbJR2XxexDttXhwpnrZx3RS0+u9nB8RYoareTIfUeRcpgOhM9i1S0BunNJC9ML1
St1m/vw/xL3jA/JV2hCQgukdTnMqVgc7mljDNeJJ2HBuv3r6SlBVTbSpDii9fQwTajLrAKx8SvCe
ZwYSuFLiow8q4A81IB4lcVXdrNdaU6+dfZAsQSCJCn/JHvpgxLSh26Fq9iVQsqxibRe5qp/KS3Jl
w/PdLpLIALdT6/QT3ByINYDGYBQFmRdwaU2rIptv6gT+lNX3YK5KVp2n5z9Yv7H2AzIPLpv/Oq5F
T0WlHBjIXcBrvNHZp9eAKoqJB7y4J0e4VKyJZFBcJQY8VTw666bgultg7YfTzWwD/+AIYRykmS6T
3iWeYUl9myixapwetNBV5ngpz+6LNWPGsXnz02Dcl8lEWMB3kFYZmzOhgtBFn2twYMoCDtf2gH++
L7RA0ckiVs7782BK5QVEMmA0GgWGEtDL8MgVhDQzdCzznxLBKxUmymrlduBJJ1SVbgkmkOZ+raXv
oUh7JY7kupIInAQeewyqsZjYkAx3nE8ujhUztE1enX3YbqKTTMF8P8+9G7AH8jX8Vf5NVXuBH0Ts
bLoJh9zrT6ztbUi1ZK8w66VVbyQtwlrYm16v0fDgzkLoCJtywYfRkLz9+KRVC7Kh8PvhuCCmbpNe
b75bbg2B6aKAryJIkU4UV9OyWuqdeb3rTat7koSsWYJ74lNpzATshrS9bzQnUSDjbXkJ1IciqyMR
t+fG6/EACZFU7C9cDsudPOsNGBACLAab7LFRPHqXniPTUFMz09R1y35EteTvQrUvj1AuTxZpu7nv
qVHRgU3tShRFvU5BZ7Gcendra+TlI/OBwPA7Ej/DuKGz4r+nyOGjo7yHoAfSQ1TUJaNCuty3Hmxr
OD6pcHvzBHffyHl4W6GDKQzu43Em4U0M+ky6HtS03eeec/SSXLFXGNFeO1qoueR1QELGS2NeQ0DF
pUtDIY9ZSrfIdh91UMJ/t8hLb0u41fIo1uKNqyhqbuoR7AUQJaRKaPHBonEEpiGpOqweeG2AFfow
23xBJ0cOuBrEWfJD2S0+wWqEj5Gw8r+j+mSHjVz4MwsH2+f/7K3BH1NxaCIoiSjlxr+NVtBfFRwU
/gA/2VPsb4YbjvCj0yWMIJtc65Z5rSehLcNIYYTwO6s20oQhcRGxnxsJtG904t8QpWsf74PFVVua
vH54Wqz6ybEKCEb28rrMZMzPdMIchGj9XORgAJNKtQfGiF1Wixveiu2I9oblu5vbw4r1lvSnMtJD
H6AYI56d43oU7PkDf9ypjkLtzYQE2dy8JA5eaJ7opQe81I3oZTp0enp9yWOvt+Tis31d+Q2C4DBB
6DLA02iwQ5i5SFxBavHG/lOFRkAXfSRscbKcUIYnOkfDYJYTmRFaOdKqPvmnYIFHoYa7K8YAnB2E
0XfhKIlA1i/bajE9i6MRX1Klt/UV4rEWXhAmRP5IbUGo53RZIJ68lgdmSn6Hu6+cHYCfcv+BDKoo
mYrBo+odsf650nbSvsicmw5/tYt3hxdViD+OdMENXme7NjoYgPf8pTiIcIHj5OhSGCuyOeM8lonN
zc5PUTdvQyx69QyXTnJGY/l3MENyungn/0+9kdK4e7VM+/J1UdA+y1BnJTQqLRSg/jDfUuMWS5n2
8GC6cArcstejxouPCv3YudIebNYiB7XO3/ZYlzuby7AsnHeQBPMxgEWVHUf0hdBq1WORC5NiZZTB
r8u2qu1wNxmqe4ebbWVQCS8wxSDh/T4CUajYrN8wNYn47dc4d3ndJalG1k2m/wJDp29nVCc/daDL
9hsw76HopTxltKG2EcojvGZmldjJwu4HiCovpAX+0aJjh+++D0UZxjDyNbjPl9WUdEWpTstRb6aL
DTYJe1aGQhOQEHAWNr2uQdbKpmHWGo1T5/WD3CUSyQy5jdEY/h9g7vdvR4Szcn780vdiNP/6e5QK
IUNFBCxupZ/zEm4L4JeNixB4gUiwklUwC4a12nNXINe9HEJXviNHak7+9djpUtG2KnNE5lqA/rp+
7aaRDrsFQGXzTTtX0FgmlYmvFw/s+9f+UxtyhpYqz/ZnyvqMe5cNg0BAowF4ii8+2eTVpR2uudAx
b7aoE0EAJT/zyf6WgrgBjAsWoooEJtdxWXfO9VihtaNO5ZbG8IcAg8qKlwr5yTcBTMMGpsN17hDz
vv0QdApKgUIqzTxYZaD37CLg35kA0M3H0xbkuL6BQjbXzbKq4xCIr0oDEnpTnVfGSDrZEI46U2wt
a23RH2oXENqpzvNEO4SHRvG8v2HWsFX995eZLCdw5GLQ31YhdAwIUC6unahiLzLrGj7Oq0zW6H6o
azWuCRF0sy9HFlV+IwRUCbHbewCcT3pltV64DwB6F76Elw7g8eZx+Vp2h2SwR7ZRPa7iukGS68gb
jsrtJ607l/wHFDk3zB63yTddsEKCdSYnt38V0r9yTaGIvtspR89wLcKio048YZEEFH67bWtWs+ha
iBjFo18M6jMny91Cfe/XVmjYKTvf0nZDk0AswLEuOmWAeE0yMP3rv21x6wGG+RkbHQ9xI8w+yYcs
LbZdTzGG4TxzznPqZVdUGUCvBlSfCgXbu/rWJLFaGQnlB5PENTKYyI69p0zCV6Dos2u0nngseAtI
XHF1iFrIP0sry2fDiM3QjBP7/059d3AVBmKZQ+FCE3V6TLKb4ZB3ZVpVZHGtPgiq8KKmLH4VjHnf
K2sQ0FeZweNNhrypgcilhxwgI0V04bIg+W3iXJ8/RpybaHVWzu1+Aa4uU7PW9CcEFLd49A2/cf2t
2lNSuczpXT5F1GVleVIKklEgj6DktI69B+pNejiVkhOop6VN1IPGp43sDbqGx/TVHe0NkWJsJd0b
Blnl5gVg+iGXsxqLQoiDezOUFHGT8ITHD9YaMeTdRjkB/437rIR50I1BqtstNJ/PPTCGlRQUeXyK
1mOYHNZWQacfO1tosYvs7rDm+K2N4Gugeqt4N/UPT37vVyDr+Hx5612SwZGsvFrV+iDLuuX0sQfT
JzWMqcusoRvRujzPCtJNVC1pfTnRc+NOB5uHsMOJXsL4aJrVoxNkZAHqHFrkmvLWvD2VHcm1iTpi
QgBsbcOL4MjqeF8Tdp8N6gl+sCJmxJIXlS9283Zc/inzZFk5BRXJDxTMNSYRjCTvdoH8YbHqGDNL
wAAMR91QpVr3VOvrWTuYbi6IYZ/kuVCui7ma78L0tcWVuyG4KS8dXDIU907YIC95ZVyM/qmfFDM/
gWlrHLBK2QIfBcxO+FM7EBKctX8FM+qhH8sGrWWfmbvg91Cqv8gUYT7zSghDfkD+yaHumpMcpvkH
UzokENR4nL0RFEfT4pRnpLL6CFX/oPqV1IKlhBj5qv4JyoYOJFQiev1Y9gNpY7NORHDkBIEqFm6K
6VQnDtV0k1NpKfkGsr6SQOMC0oOtnOX4IZ+NCzVaXFmrmLxmG2EoOABB5V3fvYoJYryaTKtqY8Hx
Snsmkj+X78lIqyF2KYcNIgzuj2/dX+XZKWaRqEQY2s6O52BxS0HO6En0wzXHfuToCj9KEAbpyGLT
PT6NmC9IWsDPpV1QKNPdamdlqNRS1W4NjlFnSSuTgl+6syOOcIy+3Xh+cRNVwmXC0IHxjwSUrV13
QJCKge+8xp+cVojVXBD2WwFc7k6+tACi+BHY2TousYHaFLkeADSoxnjt+M4Tua6XNaBB2cLMsNe+
fy1U5RgzYEy0pAW10hpBq3xBcVWIbAhvVOpynCXBbWiYsWoQlnVFXmwLohrPm0RUfo7KPu5tt7IA
Kix8Vg3x24W/FrimdYlOnuUU7s5wh0BjrycSjy9b0OfD6Veg67LSstY6ckLUlFarw0THzpe4DjB8
SVsmWhqhNFqtCPm29ym41Okn1SIo+plfbLs9W6rB09kjW1MeXTwYtBqXVUMcgFJ/0KF5ZXbBAtfh
CN/BPNcn14EMuNLaLWxKQjfRqUyfkxDMY9mmgNUbM6thwCyk1M8fOO5XLg4Vft/wGwU6pBtB07Ia
6Es71XitU880gfeixU9umy7DYngMVWqpRYvXLUDu+k5E099oWiGWod69ynaF7qk6mBETN/QHcL5m
q6Zk+Pgnjecp1KPKfm199E3ATqQnPxXWyZjBqdumfj2QPW7pY4utQ4WJrVC/RGeLuXeCyCaRZvAP
KchyU0MLrFQUkup7xXKkBwgNebsOUHTNYowQ5XXGl2d+tLeLdA4Zfw9tD9idZx4RHOpuaQBVIm1R
MXg0aNpto40b0c4Tj0NIHPVfY4RxAN23akv2ZRENWEZN0DUS4Pg/+Hn07RvWmLaVMHMS+DcfFzrF
J6+Qn5ksT761Bg766tsnJ8VZMfRFXHZklF818S2y3j9mgc8UDYyD50HkEdSojAdzb7wOjuENpiMN
eiWLroPV2yml1bVla7ZmwCZciDXW68zpNp1ecEuu16aoyS0bBQNOmJYfhVhDCmRk6+wWWrYg+Sgo
BPneRhWrnXE3Klw1u40KNY0g0GzhCaeC0hP3bO2ZkESV3/idlZDSEYzyYchrXREhHt2wrFjUNQpM
xXxpdclRwQGI2Ri6kwOhgi3puCC/jefPz9gkmpLTcHlTqkb2ZplbpG7hTlLFv0qOPwKY2M9VqW6G
vQK6ledASk+fyVkcd5ym8HKZ6Hn9kwxSXqFxyO6J9Qhkzg4wPBjdRdriz01cAKBHRVF0ZvN1xg01
gyl9ANowKHK+4T3kz2vLYJjMm7MR4Z6FRLneT5jSnxNjs4Ef4DhpsIi03tW05BRwNLz+4ufbYlfn
LVJHxumLr/BF+hFhuhEyMIHWEZcWzEpBQCfi1Oj4XnqaGqnEWRKEyt8nOqR3UHzUL2C8NzIpnSlW
a7xIlKSH7KkaCK41ko4zts3UCNdTQHKeCFWRlJdfx67W5vr+SqIQfaHyyXAQPBTwTht7u/qASDXN
ulhLi7XxcEmVLnQ1iu50Lh/75J2ouUV7Izeo5ugRmMi5frjwHWAGc/EIkQK0byj/h0GP2By/JSFM
MiEJUsjzvVwDID+oEoTGTbYzRzzcvEQ2AUlMyj6SpZpb90dmWoU2Bthv4Q2E4J7chGCdwB0p9McW
l+zYWIsUF1hD+jNq+xlym+QGusu6+XpCxakG/ihTnVLBAcPVQm2hqbDO4GUyZMh0Kmpy6op1/WoQ
6H0uzCYfsjo0KjH++NuwW2cYC3S7d4a2zL2RPmhSxMGaDLN058JejpUMDtrS4MIZCFRiKCR5EzmO
4KYwlO+6C8r+np6QeZzspomKRp5veMbqeLfKSL4nGbVsaX/nnlAP+5hGPJKCoP/1kWHiGoCNqnnd
mUt4Oe0+NOz+E2VTI2SaTNPWN6F3yXR7iggVVZ42Yj9wberRSb8HJXJWjl3JQT6nESoR9pQuI1j+
xwDZ0uwNSwmPfcB3ZLtvpYPg0sCc6qEeODyDYgb0MHhEfrnrKQ4ZGkg8gYUefc2UB6motKvC9syY
23QTyH4AH1/sLES2hFhEy6eIV8+xMXqpF+p76ageO1Tn7yHxsWznOpyEQ+wnMiQD8EAtUR2eWSVe
J5brRbVgFl3vj+gHuRL5FKhDjlYauytvR2f32YDrhCdXqvgRiddYGJ0SGstoYfKP94Qg3Ymnim4G
BRaVHS120JoSfNxT2APep9zc9wzoAgGaVoobXs5IrZ3O914E+UExRSj0FHn6pNyZTjDgOv9G1HQH
RsbeOPRI1e5qIrVVdDbvFihJSCxmcBfn2redrZCmT8CCxZufsi4jQVhwu44N+TDGEgbrypxCm5nZ
n8xrDPV0MrFjjVT5EKkXwit55CwWWjr7HPtq6O9Mo4mB9vJE4bzq4Sx6sIStDoRXE/UN11k966FR
MNWnNuZ3FhLHy0elBVkBcNeFUqw5Cm0niaUiTztiYAwopVuZpWcRI418KIaddGcPUzIQh6pNwchx
/YwSYdY8zIXLRXq5FuLUTputyp5R15PwIooMsNCFqdVEsJG2QZF9mx1C55uw4g2VkGtCnMdifg9c
bn60n/qj9dRtuYSvmVTMqEcUC5yqdfjWdCiOjO2OCOeP+uTMbjBH5S9UWnqr4yM1ZugDQJ6CKL4k
JFz7FRFQNUqe8C8QkRQVrMaaVvyP+hdEioivA8Xj//iXHcBe5vEqPSqMi6Jt/29kCS7suJa5NLSu
7hXDFKJZCo1iARcTgDGajbz0XcX/eH9YLP76RhUeOo30EdXuv+XAxoj7ou9MFhReDDsBYZ/QyV/v
EMKshmz5+hTQ6mtgmL3a7hTdMse0/vFxkV/kNwUupC4eJTvgEMknQKWlrs83rL86iC0ktBrXTUmz
VaQgwNCGNYrQ4zjJp1HzwjivtyxBd1ULTH/jpCQwwB/QAw1PW8oFV3gis25Br0WhzJl/+tUbeBYx
WXQ+FhlwHE7z8y5lYjrSBRnfOAmGgm7Aubb2HNueLgf9m8VURPD6dHixRq8H0DWWOPhsk5yQ764Y
tAcjdp8ydLSfDqH3qc9P0M4r2MV4Z7QIvOVgNTiom1BOPGIfKQarZx0yES5VH20ce+b3WRRz6ZOl
KX73HJRYb4kH9ekJ7NP7zeuy09N1mj0ebM+h1n6ikratijCkdyxo1hoRyZi4SmVkZ4d+pDbdrtVx
cyGrVqHA2WQjz1fxaivAsuD0bVRtTUFiqVSylQtbKW3s9WaBbH1v2GPdeuO0hf1mWLH5o2gKdAdt
tm6vKF5lOVeFQmgrevuSi99HvadVu8/Y3DsxxV6fgVH5bYBZnz47dHTASpMhSFHgSturoSx9uZmt
1VaazJl6/JhwspWFkO8eJbOkMb+YHlDPaKGOVHAl+nuUh5QqyxRNAQc3EjoO87ZvLhtfEqMQ2gwB
GjYNhycu0C2BHBZO3jhoze6kuDCtuwy19mS/7k9Ekj3eu+kTceyEIIxQplMgdIbOgRlUwrOquZfk
C8NxxEk02E7/B/NQJ9IueeTzVKVOk1pwC6v/R0fQId1u1JPIkkn4NFrN3GOAfIV19X488oDOwLrh
eXVj9HgCemwVfzsDm4RlmIxgN3BNwbj/Sc70/CKPKCxw3iSamM1rw8HpXbNc4caltCDWEH0XbHmX
3jFjXDcBLpuM9TaomQRoWIKE8z1F+WDalTotmC4fR2KFLPGxWlOxgWxnWem22+QwkAtefBBP3iPH
GIUUhn+OkLat/kIdWx47/PS2m0X718tw1VQQLxFuTLpiRDxWeQmYMI4aAzPgYeqlPPHpbpR4U5ik
T/Aw+9hnClS3wLAYDO9PSylTk6u166b+vwb9WprubYdudHQI7EIaAgPoeSZWe6WMN4sv/ARDh3+V
d6OSE6nGr+ihUS3azsLTqOmnFTM3QOIs1n/fVifdLKclt1gUEjM4kZyq28MfHZipTxB3NCa2hK1u
hLtZI6re0KKQOp/QFQQhcrd2PCTfIY48ueiVriqbm/H/fsQqOMEYQUtQox617XAFtGVR5ISzRW/m
lJwJg12xjiq8sueLkhnR4iJCerUMzVXt46dYKqaFl+Kkf1QXPA3cb4QR0BBUejMvG0T13vYncKWg
0GmXLFTNuj/n/tFh04/SDzboflxrYguF4pG6TqJEW1BQVa4vTktPt+rOWGLrZuXf4FQgpxcVXCAW
P7KWGLOSXZAl4Wia/ZSKTf7bdbcDFymA881LSDpEPG1wpsX02jjP6MjlOm51D00VGIpcULR/kQPL
Fw1fDjaM0qSkHBXmfqzB42OLgNHURHZ1llaNqpS8mZcjE064uB1bII9oTkU7Z0dJIBg7Tx7gF5XB
ABJW7nJtbDiUEOupi4PlXtmhMKpOa4Ph3Vut4+1916vDh7hvKP2ndGycNke7gkHj4sMtTrPAr+aG
xdffXfUIyeJcZN+vQQazHVcy16VJktsvxolTypmLWFaZ8cm2sNuUKAioxbuqnN34u+K0Zb9z4Qdz
tV55i2+/SFmrdgYkDeNmM28au3nJhwP4yCaADD0qvGXjVoToRQww6SbjqZPpjsjiACYzSiWUFtH3
iG41WjdUPoRHKfFl4DvtHNIvBkYriGJ4dmfWMmaWkXJkHdMpQv8GZtEvyyeSkuk7vKkj9wJN4y3J
HMuFC6Pmz8aAQCQCx2qckp0ribrV+wSRYwqSHd242fNywFT+EGbncIQUJkEb5zY0dyWqh71pHSuF
SyHJGEHp8M9DbkKAg8eRYUYN2mrgl+HzbCPTjc6stovUHNHMEcVWYHNPzEolMh/m2b9+hg0bEXMd
WBNaCe0Z+/U3U7m1oBsRbMKaj0Z3pSm5vV9A2IaVUT33pjs5BlEYw4SDRojphegDf3ZEVNtU/iMI
5qwu7XjSCLUJCVLa9kg/5tVQosaYRo5l+yMggPEz07Eus8LkK3nJferGbCZtorpa8K1noNsKaqRK
aW9YUiL2n4qK2IlJRuRxCxrzO8iZNNYQIGB4oRWZ+eHreG+7VJ574LOHXxZ0sYDmCJ3BuHa1lKTJ
Rl7E2wDs3XrRZ8Lqow0f9Zc6Da5qHIEefw78TBOs9A3SXvCTg8g9qWOUUm4BB1zk5Ip+63NFAcc6
4Zt7qw2bR7CdylrRZFjBI3RZDptvcu5YUStnNkzD7qJ8kx4cnGxFMj7OqLP64B4YVpnq+XPR6sPW
9RXuXYWYKPrGhgF0YwNP7ia8nfHs8+gGnSNES4zjWHrmSWk++mEn3EznTdOwidubiEN6ik6FI0xP
9DchQEL+5FZYmPq8DFNRrlQTwmy96xaJ/YlsIGTTvwM1Xq2K5tuZurR+j6bB8pexnrkPpR4MMQ7i
lgcduTVWW8yeFj7Aw2jwTAROMiZLpS7by1CSTIFN/b0exf7eWNhP4J6eVwL9MtRssiNyFylAja7Q
oErOyo3s2hDnC6b9bnCfEJY+YeXs5pBeZ1i76GX7XAf02dSl+zuPTzyRPcs3gh68RQXDO86Xo38d
r85gkanwr64gXQfhAms5wO1sWY+li/PHnAjRoBiJ7AxYcfp/btBKv1j4uGgB8cQdvkMoFKW9cL/f
VFIloahle2T46Idj5smhOeMri3Q10fbBkCx/yThwDurEB4JItAfQQjmA2JzS7UvIPVEZ5AZPNwOC
WZkdjgLz91uzAtVIIOnu6Y0uqBWRe3fSWo35ShsVcYYb/bRviG+TDOA+tHxuolzjmD6PNwweMopY
gS28CNsNVmM61E1IQfJN7h336ctNVFDXdm43h8H85vzEbI5M02PIBW+Ggq7r50XdftNfwA3HOqga
xHCRmoKPbh3aubPeVe6yy/Qr1sNPf/gjoB5C3178wuxCwdpruMQMBuEUdPS5V1Y/QCJQeDJsebMu
KSQChUJ8MSaACdoV13kHESrh0LDejBCghM1oUIVaGZzCVY/z0T6SqkA53wuN2CWfT4YIT0vx9Fd+
zcqKDawO01NkpZMdrZhvczncZ944IRXOTRMP3DORy6n53IMfSuaOn8PaEGI4O7BixEPeM1RYAkOa
9TlkZWn3mnCNZwLatgejCKVLoFLgLC5ThHEnfA2geJ3KOjYd3eQ5pXtXKLQxClZsqTL0/ZRAr5wa
Z/w2kEy/Fy4vnMWqZ2z7NooY67WjPCkhv1YbrTXwZL5Gcf1uPMAiXaPsgvHWYQgSZDSigyEXdCVH
iOR44qWJhCk00kYpjj9824kBWre7PJRN54fEgppC6o4YdfuxBvYoLB9DFTFx3k0MuRwwpoRuo8MT
cJtLKxIO6VLGcLNYp3KrTHJPqIV5wbxpeQSRQUgrT2fUfYGtEvActtXtshA6HWqenuvQXyvIKlbP
8W8+kUUtomPpHzGa3BKUy2SrGwYW+gtBC70KMlTzVpvOxFmoSFA7DBJOq0vCK41KqYBu56Aj9aqC
GizLY2XOyPQONTKcRAIqiSSifeReKl8EnSrZb3/gPVocxVM7GPpzZQgj7S5t+sPl/XUxvxGG4Duz
Wa1NfzPkZzgse0ZyFJG60MHUGJmtRXtCaU1Xy4olaqxFFk+TxWI7OQKDZZa8tGVzBjwvvj6Ennyq
cGPriX/bIE4fecHkm5/pnr3IrjuIAmK8sxW7t7XXgwohKcjddZb9R6/pfW+3g5BrUigX3MTWqbbK
r8aAwKNH8df1aug7ic00bv6bKygJ+EJLpvSdxkFwIxBKoNoCnf5hko8wz9bK6bG+oJJp1S09Ujwy
LDmzYU84ut01kvPid0mQEb1Z+U3OJhxnmjm9VwaO8wV2seD2yyC2Ch/DOJ5trb6Zc6SrXyTZdHbc
z2Yr84Rll+zEXMSx8aUVQWRVRbChBh4Sz9kEtT8LrCAOYN4P0Rt33KZ+OQhbm0H3/FkIf/SP1nSm
9FMhlPX6JCqG7Hl/dfBq5gQSnhL7/1u29THRCVkKKLJUNKnatzrTYLrDOWNEWosv/RC+QsGtVdbg
P++DrdJrEzBq09a3TnEYyTYO0untnb/Irt6KYBEnJW3oWv7KkhdtUNantA+E5b2olWHYTj58+0Ja
LpZSpSIh5SmwUzSLc2zrHdSpwhww++17JhxEg2d5N1pwdPOiV5u3bU4b1Bq9WORhzrekbc8iBJEG
/KdQOwLQKGAfi6zlHKObgq0dMOEMPn+7PnqAUW2nWkLjhi/C/h4Lliz/dgRiHC5GKMCOVYQ6GWo2
j7hqUOW+8Q8oF3vUEZaZfkQfIkUBLAiimzP/NKmEskJPN/h0/COZtAvgqi9EKakKnY3PbuBzYxVC
ShSzwXPzKgfIHmMT7H8Yb4mAJcqL8xtqTjT0uvfPVQCj3I0P/1DyCF0qznHuaHKzo4OqlNafemg0
pLhzf6nKdkuJWd4VJv5MPlA/76jBOOqDepsmvnLPRB/vE6xh0DBDDUhePGDLxx59c4EHCEYPyv23
BifyDCduzk8MLZw+YelmjpeEzvlFjn+heje9Vp1Lcp5BnHs2IAlfSIK4uB9BzjCnF0CwGBmnREZf
TsgJ8iGqZT6YIMZAovG91lT5QjKbMKrQIAfiv18W/susvOzWH69le1pp10ffDS1EZPx4AL2iuI1b
EN4y92Rf4BVQiRefF7djpjsbB/t4XOXrtbvXwDyDZvloQDrlxPDuX38O4CbqrEZUXtqq0mGwrtFS
zYmttGlqVJ/WvDTCiRlWKBv/08lwMPHmn60gNGffigwfxgzyyHQLLO8nEk/qfU+gJoBNJuk2PrPL
PW8yfUlT+mxPl32z6qixcoBv3iI6XaLO1KCIgdKvTMVios/wxBNP2fubxGyb6izR81FnRHXqY4gG
Z8/Ge9u8/kUTnHIX03jWZE7dDl7IcVRbtpL8Aw7Uvv/wTbHqi1sBK8Pql1/kPar58Gsnb3tuvjQO
Fq82p3YDYGbh1CvsCrI94IANNvCsYqKkfWPr2mZc1WTo1MH2tAlz1/FC9zZineXilt+bRwcXHybi
jlAS6Wl6UcdRjNHF2nG46gjk8E3Xh+sYmJW9TJbqPtuDsmWOQ+DNmzYAuxgGde+4i63k61B8GQZn
h+wZ65jNooxG5jAvXxT9p0fgDhzSRSry0qRlScMlVVJ93D9ZBqX+nwjsQnnBukr1QKfpxDbu5egC
Mf5fVpzmu1icl4QMiWkJLuine/oOm8Z7/dd2lsWCeOtQRCCOf06kXmzME/+sr+p8Oe4ypjq6vK2f
Ny/9iurtxzwehpxc/M+lTCXfBsz4lKVVCnJpxwtGa1Ut31Y3AsCLS9Nzd0hKgDkG1NhDNR82FtjO
rxJg/4oTIeO/SIaNhuBZXiV6jVGfHs9CtIZGUPXrh3onxI9cXQXRkmdWArbz9F+htKteNQDVvtbf
+WjbRj7l0tokxe7hWL2w/iu1Gnk9/o4HHcXXZfEc+vgAWWcLWKcmApg03r+SRr+FOSBiYM26Sz2L
GhvE6OGcjGwnIPWb6pCvPE2q2dl7raGDYHWDeVcFDmCgdCQ6Ah9cgBXS4dgbDJGhrLrLMBaJDKqz
FkQVIVbUXUafVHKjMLqjaIS2q5LqZKkmOLYHlP4gXcuaIXw5kFU+NMMbTOI6/uyhjA7kFbWhfXnD
PXUPVNjbgIpL2u0bp6S65YkEfFozJ0w+KUZi5QUlr956qlTXr5ZRhuZ9e2hBWw5xYhOFmEbRvp7k
ERuqBXARk/HJXee0iBoUEwl1dJ74Dyy+0OPVMj7dptqoqmHufXLLZP0PCNgKkGuXvWfeaXo9W5xc
AV1pd5T/w+i+QCacEwLmrweH8e02K4kBOsMYnzxjYMIZ8sFwq+I7N0X92kOP04eizMVdWWEfMdxp
Nztxpp1lGSagjuQsaHHbKefkVTFAyy+Q4f2uczpGeAi1zo+ZeDdfCYeYRo11XFqjgcLWeTcUu3YW
NhRW5PnmwnxStipJw8c60hNCgtIl1AQ3Eu2knp4bv7aVaijJVy/WLjEwROrQZREz60qEcs28L4Hw
0qYjgTgUp0GFSpWLKcw6ZdlbmMJkrXXVQysotlP7cweL3tHkkwek9WNookQK8zNliFJ4q8NiBlU+
4/JN0eJnXoZfqUW3sXqFcLwsZpsV5Jg0pxomPeW14P/yOvraw5B8BNikI1Sn8XMJ1HTvsV22S+yw
0BCL3bJc3CwWCaqqiTE4SLooChA1Gt/m8gWvO+MOgFuC2SDv7rXhW6ZEJ/LeibyMNQ3sPB57gg3I
7d2MZCEXShnGIi/Qy+26sTq0FlvP7N11RHWDP9f8K+TsWMTprNGcpk0vBHB6Fu9ym9tdDaxn5Nwq
bp29MCkROJXHTPitCubPWuJSVNTK0yd6hKY4i7vPOkamYHX4RA4CxjvUVGHmPU9NMSgJX3UYT+51
rML8oUSD+ZQIdeDvNfSQjxPQ1+xSY0XmKg4xI4OFehXlMK+w086zeQC4pMGrw4RVlvAKxE8w96Ce
KHJHu/zHrgKPJCaE2rUOTWMaG9k2D8VACvhMtUCu3EeEcaOAUkV90tmq5zCB1naErO5qyiyASsbp
H07/IicvEnus+1eMPgksGL8uzMPV+PVHycXeM99fwxJaJOIV7IpQkuVICqGGNfsu3vFXJZK0N6Kp
RAVGnp7kdsVv5uslnx90aX56jxaZoEvONcvHFzsS0A//boaywlgYeQ8i9qCVO9fOe+4lzRKEy5jD
3aNgFkjl6nG/8lGBuaNe4gdsUgFkxHXXhQSH0qzNFeBI2fe0aDmhxVvAnvRxGX11iVN4nVb/nn05
w0myQJQ1OO0fWPMODTcNDAqA02OHOu2PiwTAAUAEhiBTqqB+lI44YgPlIMdRk8b9ZrLKIevWhQMW
DLi7BOykIaaPze2OyU+kTFQ2mdbklBanFI1MFjKYQR4FZHrJk2rTU8pC9MLXriDrn/d5qZsyDd1R
bSpdJNTugDeTLYiUVUkrs6D4JMN/PTtkPbUEJ+vDZbo6n0B6iZhMKOHJlXbRhxgIW9udLpS/WvLe
QEy071zUxfrj2ECYv84HhYinZDFDuvsCU17OfTSYK72N9WEZI/NJfBis0Glm27Ubyp7f7cpeb0um
WDqxC4iYPwP0drRJnhPopOnJ3UfinIGhoeGo93Yp7zCYkHz+pYf+bDWqojNbbMoymZ0sYfRl2onh
wseID/V55XODYF7Vl3nKOSgfiNICpRySaiCgQP3LjkO1wcXebEkTJp4ZnUb/fYi/z4umt2pNOEDW
B+jq1Ua6n0veM1x9drDwngmQq+FHqpjBGuef/FSitQdzfcVjdMJLr8X8sKNJcl1jZe2RfK7wsU7K
Jms+fCQ252HVD3gyfKXh1eQmmArIyWZOaii67HNLsC2NKkRNZJ2M55zUAxN8rgcpyR573pDZIGLC
GLwFmwek16w0zS6buZeTO6+rtsdPXcs8pWoKb1NPhv7NFusVhG8Fo9lkx1Xt1lu2YqMLCKvx/HhD
fB+2EG1VaijhiAiocWu8/p6tz8qpMORBdNSyBT4760K9BWarwBAxgUj7M3YABaqFi438391XHqpf
VtVzgwiSQwEPrCM7T/CZ4IeQMZFfoMIUgMgy09eqfg6jkAoW/K35saGJ3bxmpK80LHRhUyt110i0
0gdSx5iqn+v/vwBY7sBB6agcKkj3e+GmUMQnR9XRwoMtKQu4UIuHm77n4XcMViKgOt8lNodQC7HW
FzZ/iUjwKqFcgb8M1DNHP2YnTsjcjoWPWAyuxEr0Ns+oY3MlglBf1ouGMq+0QNm0l3yjkdMOJ2CF
cRzHZ7/+Go2Bg9U5VrL5zNl6F14f4u4eNDRZckVgCutiayjdA8vNt1BUNGgKvTvwRgNIUPle9y5n
p62ovEj10XyQsF9hbUsFh9g0B2A4eDttw7SJ+Q6v0QdG/0t7pQ8E2viJR43ABZDy3EeosPVuJlbm
F1vEEen5Hxp+iJeimVjXqAa9NtPp7aGwlxQ2DNnxdyqURC1yCjT+bSq5gxvq9wCsC8h7ziiRcuYU
9E8bCswoBHQjvPzXwuj0PUaDWz+kVviLHqAJOr3cWdA0VchBbWgsjLWBbtCCphe58v0tny0UoSVR
HFqWqcLiWs/Zc66ZmrTI221lOQd6qcS+TtjTGdYh958NyNJeuGVKI71tua1Vb0VXZlw1Wvmq+Dyi
Ftx6Vl4AuBiQugW5pDH7N+5jtqpwAvjtTIkIQV4Mv3aMm417/Ql84yo2iHkTKImC+wjJa2azp/Sf
6OVNXD72f3elVqFZ+AQleraxkNzB7OFbEOWHmZ3TDIGc6l7pf2ANUDsKJOvx/t08iSb61roZa/k1
ThvcBCFeSXfeZ/ZZUMZvDvNP27MWxpmyU3U4hLBzjq8qLeO37lmZmHLbjA3dIM5FWa0Ghvnyjz34
ERZGTqIVNBFBubz45ckYro4bjiymXm4QF+niyfmMSrkf/+BonZuBGO1On3lootAJCbMTrwYPXOHM
EHpfxuDSyCo03VST9XbBhkZF679rmRq80jytAVXXfwRGx7A6gpvrVwx361FnHAC5odM3klent30D
FerYN0fofQmHQyE9XlePaQcbXYXl3niYywICgyb2Qx7Rceg9z/M/FMm1oJyQ4q1wnWifZHPDptai
VrFJ+r1zijkTrZrE64YHP60JnjB5f6TvbUvBjiy0fNtVPWNE1xfsoxybaoaLR9ZVKeQ1qREZr5Q7
l7JHoEaZ9qdRMXjtnuDwXmB4CjcDtnBWMqoRluqcM71Pq7onwXekED7ifMKOGn2WJ84yWWNJf1XH
E068WaLNZMbVLqf1rljkvBYrrmzsug==
`protect end_protected
