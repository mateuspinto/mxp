`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3664)
`protect data_block
E9Spru0vpRWNQIP+j5vGVmXraX8L41q77Xv4VH/i3ywa1I8ZRu3c+9t3srPEg4jd0tu7RyR3iSNB
dilmRnVZVpuQjaj2FukX0jlYujYIFNMh+qH0tbCVwD0pidxw4wsUVsBdefw7LTARD0ou0eLKKZEk
zF7CcLg6y/iAopbGj7AmCRYleZB5609J6H+RSBWw7bJNEfxs3kPO/ee6vKeHnCS/uyL2HbmWen4w
Fvc1EKev/0jvk0zjxchIUGSnlWIrgglcSgztLsOhdP2NRQVzFBI4MLaF32FllBnoLRoWirS921W2
Xkf4j9xfuoEwE6hwV8K324Nb5zbnIA5vSxDZw2YquUIY+LLJgcd68WOelkRRgi556/mCvRviAYIH
oTmdAdDoEj/Q6R7LIowpQhZMd+mVYK8mkPhMMtl14T1onPLepB10gHlMU+hlpCBiB1m9NrYayWM1
j9gGG+Z0FqbYpXqSdkUKVLdUxXADUPZtMRtNqkHkxa6s9wx7ttp54g+wtEHsysbpmyGHeO3ME8GL
ljqHctYddmvO7T3Gt8E1/kldg7/YRETkYW72zAsCxPDgbFuEnTDL+hapW2GZXtCscZQAgPqmKwk5
CwSvcTRvqcErRLiRnr14BP28xTLWLw90J129U6Ok/tsinYmIexN3jyIKwELkdRiQSvKx9FUnmDqK
vpBTO/CgJ0zmIyw5jeBW2sc+SIwZRM5rOnxW5aZNcyQm0D+kvICyuTrxCPpCbemWuVFh8oy6yV3E
hFTizqAiweFE52U5mExlM+Wvo39By9tv7ceQVLb1WUySR6qIMfO1snosUeb+8Ox5lU0gNmOp2D/k
jo1oQXY/TCQli3KFUjgGbciy1Vlb38eMN4Z2zeUwGcdUhJhjpJtTWpJGdilDuUoESbFCJIFUZNgH
f5VuFAoe6A92LunjhnHxgMcaRpp87/ee+8W5gaQkg3Rnf2KMODXSlhOTkumbzGCX6R6a4j6l/ZA8
Qkm4hYLjczv3cgoO49mZTC1+j0JL3Dh5pB6zakAh5e9lJWhCvIojbXnj0ALlwJ2OS+e0XOTLAtsu
31Jdn9xAXZmySTqlIzrcifpgfGK91jGNdtVTcTRAQUZfPGagR0g8fXjwscya2QyfFsGQ6+RqsJr0
wCOXPepqM+IspPaHb5O4IAdg6kktYxV3v6FMsa1cMJGLMxWnBfFu5hP3NKMk7aC6iRcAqWc2aj6l
wljts9+31dvZipRn+kL+C7Yo0crlZV7XiRsYnorKhfJChtD9gVrDN60b3PvgAW27eHjKrYWGBqRy
WegAm+OR3VZa8TY/Ga93Duhlpdlt1m0VwV7PWg65zVe7p9Se/XW6OTghGX/cqslKxPQgEcvfVtEj
FmThZQxW0B6vRPmg8zgu/ZfpSgcIjDQMlKav2Fj52kqd78sSJ1BpctmxtpF7fZehsgK5Oh3VUQAL
rdaRlVMLlCcr1BkhfSXfJ0FZ3imWayBMDR3UCiozFsT6yEnhz++aPKaag77KM+wEZiDY+7LXhgKh
Lw80wEWhPhLaJj57vk+N+9+Yq4F1Qu5S1fG/BGwSr7UjzVR3kEz2WaUGYUKyKRKzG4HemdUGjXVn
ZkLkHS4g1CucvJ0YfQND1mJa5rZvpBcCrE0aA6N9iqHuZHQiYgqrR/hMzC0ujWCcrh6Pr+0oKsvk
ik7zv0kBcTQFg2f4HlOWrTHZWxUw7kP2F0T5l4ZLxqRLHKJNg9meSX5x3m5I18QnUylY7eOI94G2
DKa0EG0TsemAVQCPP2jMnfWUDqeV6KbMU4nEFo9aF1YE7II+49p+G0NC5iYBixV8Hb8g2zDrwKpH
NQNdEeNZ45IRu26h/jRtsdZgM4e88fOwsgvOvPOdSmNn5g18X4fWjTynWuFizoxNcmCsbClMIHHS
zpR7r6jwTEFAze4trkqUsgRmEFSliaqTeqjpUeiFZm4R+R/O87asR8P8NT+wKJeIX6gRjpSsYIFR
b1lUHnmDLkRpu3vmG8sUq6Fn9+eoKPRtwVW9jzXSsu02fJ85a6IadL8mMXYzgtGCn82fxsVIetZp
NN6JzQFKEOXwn3JOGVGO7JN/8JvUqgBzw3QWyhhoH/IaRIVKkSgKba3vL1I9z4Kq5QwXH9Xn+aYS
UfpF5oun7QmMfjxcL3jaGraSaeSIWWcfHHZbHpaRi/JTGcSToxv0mxy957Xo2ytEX3Yy+FCMrlLd
gp1wGL/3E1awqsx+zHbacLp5SE5SbD5k08f69V4AnZjRn0IIAirdv18kPXAjMEeeUfg4OKoTWlVP
jPy1/KD4Ke9OQf/QV3Di2eCXKC6LhUQ556Wf5r8VjjT/AHvud4KlDjhFhu+2/aQy3Ma3WnXcYQ6x
r6LsTP0M8M08iwJ9hniYL2wSxOvs2KG2VVNG8nkFSO1T/Beorb+tRwUKcv8yjKUEtdWc8P50HE7u
nr6Zq8I69LF+OGW7f325EYqTgcpYLQwznt1lK+gfYsZxm8LIwFhll8y019/zDl3quM3awxYSbRqV
fTpsyyEdGBRK5EjixpVvgLdIJsIZGOt4E7Ll0Yzi7Arc/5+FCyHkYDLVOoKZCG0xx420vz5RdVBg
iWxoz+6gXEkC/hF7aKZ8njK8hkBL9szY95vd/3N9BKhf+XqLao9RIzvn2VGoEIhz+huRNKr8qzSM
BJXJNPyRddoBJOWhgwHwETFqoZPHC9FjYybVJAyp4TyVkiCglBafYtDNaePfWS068q1zUlQn+5Pe
jcL7a7HAc1OkVWkF8+dfEF9MMvAgbf7UPlOfdZ/PqWX8OtMpUYQct+xXraayPCSJMZKrG8mSjnzW
mF+QdMAmrvACBKdPqMzkYNx5SaUdOpq2ULOBb6GXMz1c4xbu/lp0EYdQAsK2j3xd9dtEP5Smq86/
FndS5tt4FFZD3IEgTiNcaWj9gzWdb63duRHzMrXd4Y6QxTnZaEOCBE6xmTG3fssG7Em0kFPw9AhD
UlJL949ycdy3/B5oFbO2wSLSPGXwwWu8xYYmEkDFnRwuxdf4SzLWSOynBAJ+kA3P6rWH0oB67gXq
+4Ctbr2MUHHJU5YevNgBhIwQRWdgHyrJBwcWD3y2vfVbTveDrGaLmXlXqPjwYQtKAdxlveEVWDiB
RNj9hw8JH9DEOJ7NbJG9Q65jEgD4jpIulLn1utuNvyHaNkKofZ2rDNNSnhwhtPOL/bOmselamdLI
C0K23EsvjdKuUV53IZiK5Agu/xhCfX3NTLL41QeNsSahbS0iJdJUT7thB96WulrXwVp7pbl/yggE
NcCXQ0OMTB0pAfaePvIfa0rqZIOPedWKKeiNSPTnnNQQK+g14rktTPzJHFX826WNHq9cQDvkmD9I
epB9jMg7EFTPu9H5U3FCgVHlvdwvlYVBSPtD3uYKTmOZp0T6YQyU+UYFyLItHhpMyDMPnlXkG/tW
Jb1QEpGrSeeL9EGSDpCaGVeQOX/yVVeBv9eOTE29Gztnn1jIcze3px0W2+iip6Oe9h486BHrZ1QK
AWX1G4oxW2aHZqzXE618neXXsEoYwebJ2grYETDJYLm838TOYW0W9KZKtbwMtsTFX7Hc9AxnhYvf
MYN8hZOHZ0jtxv1sN4FSc6Qbz9YDSPW0Cqa93Xvm+q4uEPoNzHRgpCdX99SecmbiWgxhj80Fb1Nk
tOQKvcrhNDultJvP1rYDkkPG3Gh3Eq6leQ8RkDcxYQsWy6nCZZOMgMoTPbSFSvUg3090vMoiedqy
icZrCge0gdYh9zekhHI4yEmLWq/d1N1LwVjd9aICFqBg7ilWVVKO4caGwQnv/kciSatEjpr0RkBV
XHz6LZN21FNs07GQA5moIj2P3Os4nde0fmqvvT70wh9Irw/6rA82I0ijxV7G43oU5fDXj0vQXHdv
epzibyA3YlqE68A5DBB4e3EPFvtM6JQo9Xw4mhx7984nv1J0Mca71dZNnxXRM5ikUP/wLiISTMmK
TPJuu1EyrVRWBY9mYoR+cMe2zMq38W4D5nmDuAHAM2FENVgl+5jLXvSWObWQnbgGORz4PyxAoDV4
LiBlJ1urYDXPICldXy805jDrxdvaHrI9xVUvrop8VbVPnw7FWTUtDbY1+hlLoIWEvG4Ool6pN6uI
yKQcvKDSnmy5CApCn1Lcr4KglBhT3QJ9P7AerCdfXNYhc7GivPn0piPSTTV4VEX33b5wC0k1q7An
W9K6gRsgvZci0Q1iI04rixVrfiMHrNVIm+Ch+2G+l8nW1ibHTHQ21iMtY3bwtN3sshf6UAbye1F+
wt2tq9StlUXqbopJRTQOUAD36pfaaaeHtcj5prFol0givYi97r1bbUkElm6PR/0w9CtZN5C7toBy
y0M95hS4KjJBXbAkCZzVcmei1KGUXKjcc3yLZHY7cSiu6AJQIyJtV1msUXBxW30O4rvnlBpY9wCO
aMn1yVOJnzXQ6fk4AzVoI4k3/jRmZGShvcKZ+CgUYUqTRk9pvppZ6/vbRdmepd9MLtDK4PJjJqsg
OiwyyzgFhDDkcr2NZ77NnyXXLchYzRtBM1OIkOei/li4X8gjccwDI0PRXAghepBT2SGZiz76ep1E
hHBjDKEz3khIhq7cgVnYar0vc0VPUuJnL20KD4JKksk6zsTmRBTvB/YX+RozSBoQ0TfWuzmAKTht
f5g33YcPitCV6cvb05o3P82MEd6j6IEYBUCqiPa6AyuXJesy+1QF6VZMYhfjaclx/oIEiNocW0R7
H7VJouUphexyYeBnowA6PaAgz3R4ute5hqgJ3ART9XoBGgIejWU9izJDI9GQvBXURvff5Zt6fHPv
uq09KHUfRTh8L8EUMPJ4Moh11GqKcFfwGqK+ky0YOR7a7jfb93IMBfd1I3+oD3ha+N1kc4EuG/rS
i4HGkt2VtsmDBHxjBHxYIA==
`protect end_protected
