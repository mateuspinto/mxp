`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12192)
`protect data_block
oTwF5P2olxkYKdFn9aTOPmJVA3SVvGXSiUGyJ4AvkRQeelME4kdmkQaLnqMq5zIQlyH0kYAtQfId
UHNjV9CPri/12YEthTnLQslQyG7EOYDqz9eTznjnVVLcnCcH1UvjhMwWcwMeVuzTTH1rFGN6vpfF
8o/mFnrq4zsoD2r+H0iC8aitmtvyF9cU9LOotE41LCaJlFFnEhOzrBfLlHq5L7DTVdke56/JTpWm
z8+EAZpg9f1qHQZ43tCBMnl9czLATevOPmZT65qmfkiiCSZK5OwL+rNp/h/x49xQ7vKw0pXvfn+6
ZvjlNLHZ2lPWH/yDWhBvHsc6iMXXObp/eD7qfGL5J36BjYoi/a63gupIrDW38zNO+v0ux4xMEDaa
b1nMwjd3pqP7BJQOFJHeCKFKeAhXa0QUUUamyTbE6Zq8WhLc/ery80dSlHhVj5n8wz3eE9PwwMp8
7+xTYvCxZLNRX7fpcveUECpD7RyEfQXh6CV0+d9Hvna/CzlWhNiOwXhNx5xmyAkPg3jtJCDhjhM9
9yOpfvFr+I3BiCiVA63rJrpUShdzaoYxRIwEVARg/E7CscO/etGv/3vmvD3KCZpnlqD9lPPh9GxR
Iq1qVNmR9d1k2g1v3/3i3IsRLR+2F4UYZUUX4MrgdMDv/DYftZ5iUvf72WfcYQmGqzmiNf+E8l2/
D7NF6AMgw3Key9YWmg2qD4SyjIFtgmkTb5vFudz50FdJDKu+z+5ZNLAGLriKSlYTNoFadpxs4LCp
5/lxbSc15usCxMVRfYo/7SjpCiXX4KRxdbv2rUlyPiTZ7Y6D4k5G0UYcjotMjdOlSKgXCeh/9bZ6
YOqDiNHxBKk4fbp6PrAjijHCp3wPWxqb66PTEfZy2QzFt9Cg3KnH0aZwtaBAU7aua4EOoA1KsWkC
Xfl8XLLxEZwAByN6y22iYsgGto+n2HcboiHq7wSVnCWJw9D/lMx+T44Rh2GtFCVUAa9M7m0VouGg
wjON32lXPXCPuKfgon+fSW3yom4NsaEO7hUh6ALoCtHtxhxYJH/2zZBrokdvCfZ6+mmQnTXZW43z
Z3sYBbXPAF5VkbfQYmzQcbemcCyrViPTM0GoeJze65Rn8XLMxQMs75uxiMsqcjg/gfjqvtpkmA2g
feYiwrMXsMhtyqEXP4HMJIHFKmE/NaUKlSptDdkqtX3GL2sJYoteMT7pPG8jnFqv4BEx62uEb5LV
n1k5Tp660zLFQkM4gH1KsyR5XZ1Op4FlnQoup0WRguTX+f74/uO1i5M8AgKKbnzEm1a/Hv/UQSsW
w6MNAUlM9PNuF204SIDwq2gebANQYlmCvm+3maCckn+CjOkKPIHCvTgWAbROmUFMPeAd94i08XOr
pW+pjpqr1WY4i5AueZBPkE4aTHAZtZ19vO4o5jvkNF+WG6tRD3xZ9la/Nqs2OCCpGHHBu7bCmjvi
hjlkQyKt4WRn82psj9Ta+KU1iPD28lnVMW0OjPBKC/WuYwVoRKfPiWYpwRny/V4I5WzEKP/pMtc2
hHwAjbrn/G+ebRV1ANRz4zHA77ZZ0L7J1GOYYkmBpFQau3f9bp83xnll0GGyQJ40cwCP8S38UMLQ
toooWWEkfAzGv+gt44d7RyLSPZgy2br0JMv2xE/VZ/YPT6J/D9q+9vBtMpGm2wK8zvoR6v57ot6B
1NX5Z8QfGjZ+7LJnKIdkXZuLi3ndoWDiDgokE86jbB74oJTy+wuAxJAJcWcj2NblLO17aXHvXqrS
mzYfy8JDqrc+zpg4W6W+UaZ5pQrWBqOuttbf72juy+0ML/cGffmo4V0mLHJe3xtEIKjF9TYC2bzl
YhPQt+9C+H15FapWl6Xngm1kPyCRKn91uZAKDWRGd3vYtGVTqbnTd6ofGHC5La3msRLP1MXJ6cb1
FHqOgGmGe8zcQEgIf04vQq+UljqKQsxv4QgfBbyxezshe8OpRHBMGh5AzucwdoWQ0EwrrDzj6Gp7
Ss9WDhLVvNHWPTsUf/4uFyixamIg+xnOAPxSTgv1ol6qqD4kQq9nMrnKR1dXhrHyzt9hpJcTddBc
PDuF8V0CdF6T3ixCnHQE98q1hBu2oHhPrK/Y2QEO43f5urjDbU6zsCspEsntnsM7L5vwvL892emQ
ltpzrryWs+j15nz+xMzwF6CZ/g+wKdtfAa/q8gu0APqMIFoDH2rjrViVOYshgEF3hmM2KObYUNjh
HQhWqZooYJG2XY8I2hvdmO5credOqZKzduTW8pL11pQUWD5jH9XZzpWAWx8pEGW8RnkyBQGN4ArX
ah1/urjNonO4a8cv6xtL7krBUI2aYM5ekx8bzFj2FIwOPjP3B92wkSPDPdBVnOJpIZkTaemRYCxd
hewka26ImsVaLTcdZdB3a8XvOkMv5aXrotL9iPAzJeVsDpYfrICub2yDYLdY0BV0SAiDnrLwnigz
uYgrqR1FcfXkboXFSu9GpBkaLAy20aCePI6ZHCxUuPsY2Q76OBA38BVoPoTsceHjSUxq2lYNSdTL
3WTuA83IxuEc0IP985RxaynRA+VR87xrG8XNBsUiuOOPGyF3Vk6EzQLSGwn3krU1ThPNjzs3ZLZc
2TDoGELFcdtDdjC7TazOulJPJ+jMyEPbYL9uT6yzhdFSmnvEUUAb07hVfOI7gmeD25/E6HzduAmM
h5dz4NJCkNttbqdyuNl4q42HqsZ8G8HHzo5BgccPYLJjjeyE4CxHx81EOb1mQhxa1+NYQTrQWvfR
nO4w4WiWxv61Z/hBnSo4aL2eXZmYlPcs0xUyNHC4B2UZqcuEgv1ojM3Zhia0oNGoL3ZyDZFtjmVa
ZWzCSQLChalEuN7CAv2GJudYvgvoqaZuEn5AKSSQxnqX9AVVhERSOciyQqFjE+j7I3EwwPaZeRyd
cEnzKH39LaFzSaJlNm6Rcs8ReYwFSb9DiU3IUhjLk8ZfG7Q04znY5Ifo6+bn9DO6t98gKF8sxaKl
ipB9HIl6153SQOkVCkSgaRHWLTtQDFy6nHnd2CtHDFGL1qFShOv+dB9Gl6E3ys3sBI7nWvaFXjQz
LNGbD8ewspDlB3+y9gb8XrLfYuDTFEm/1+Vz7dA5cXimDZ4VOEWk/nFl84KD4hNceoDKFedYgbyy
9MkIOV9FMWzmdS/zIMDpxPykLzRNU2aZDITlTy9IRqUfwo09EiGdcMicIRSe9gFRWQH5YeJoFQN3
ngF7jQr+SAdjgmJySA10Ea+j12ZeG9kJbtXR9DE0msHkvWDst4ymwofI+mFouUh1J6eljc14Qh2w
N0jA44WdXxRJ5vXVEBI6eOvvb6r9tdbxntpzEwwjstnVRSHIdxyqFPqhV2xW/wkY/48z72txtg/8
ZeF611F7PUWEgvoaAb+q9BOQM2K1SiyCWqh1zAYIFdiPUOxNNG1C7S+MTm69yYT6YdBQT2HIlFAd
d7IenSc5WZWRBsmWMF/QvEO8Tx59q8o3S3VWTAwSA7BbJzUJznksOxFiurnYDudsNLXzqiZU66pq
ELoFkDqtsJuWP18UZLl+7Qkp/SfITPc5uYouXcucZwRNt8bV7gfiEYVScbNTwgCQIAQU5iSVY2Pp
IMMeoJDRWZ/4xsfeye0I8rV50ad5fBCCZ5ZgvaJhu4yLdRThOkqNw+z3zTM4IgrroVs4nOJwH3gR
7jUATVT+YdJ98PA1c/VpJ3D0yIhC3/8SUXHalgVU6NWXc//UIVy7Rdt6lOwAfBj4xeb0mbV97aMQ
CaTr7JTzTZC5PuiA5/iKU3+LZAE2FfGiMST/sTky5ihuAi82ul9OurrFKKNkY8ku2a52LJFSAENG
tOfdylPvdona8YSx18XWjgPwPvzU8m8NHrykwsXzfCoHNfbfrD48cB0jGyy5K2YkmN6zrBXrJNF/
7QNRow8nf0/ymrVI8cpRCJX2BOp3LD2FeNJJOGPuIl6iNta4Ai3KtBnALVppE2d4GraMAhuzi9fV
9GoU00iymftDvk/v1KyNuozXx9eAoGtBB3dTbzMSCUPV6bgbesTOhaouzdrVME61smsCu83K6FM7
EqDUMtnnhDDica4liIachbSveCNzOUQof1FxKFLeRtKuH3vjsg234HtllF4bfWOLXDYlTXqU+/I8
+RU0vZADPBsBixIJ7bblimgy3Zop+Wvorf53E1f57XLes9v8Mrng0aXXf25+rqb45xQK4Vwsj/JA
fDmHpFVXSHBBrRtoEQmdV1ERxbC9mqbNvRHxI7agD3n/drNwj/aoO8YV+WmXn4W6aMM75TKui7Sj
Tm9SBepFbCmWYsPzkQyBgQR2ZgwWYAKwsaK07YxM7Ge/SiQBmrN1TPDWiDorbTXrfHbBJd86WRVd
5Ci+JEDwV8LlBVpxf0V71hXInN45//EN5gJRv3Ax3oGtx5uRqQhLRNXIPK64dhw8Tx9XqODup88M
NuIoOyzjs0LNPaVwmz9Ufdy43XbrRK1WL4w2EKzhLun+wSfBVyFEK1ybhr5eTDut7yjIbgs5qzNK
1lGekeAT+LdI+9ADZThGp0QThe9w3cQZui67LPeCMce53fYg091DOwFlcuTYQGtBUo05Y/kTXfzV
X7XPAmvssAeKnTIoqgmfBgb0ovbgfeFMSjHEYNJH2Jngwbt+C3cyzi4yI6Oab5pmhphMtRQ02t3O
i1o62NpvKlyVon0Dba0ANDHY0i4pW74fe0gUt/+lH5Ivmd2ZgkomVXs4rBVEPaMWhIO6/HHmVsW9
8exg/FhVM7kB8PNa9LPhSXbv41rS1X3Dj1ARH4U8YEv+zFMCJ5yJumKt75eX4RQmZ6tv3fmYd4S3
6nELq1cPHDGSmASTO0toB571XGJDcYMVTWHYNFCPPMtrqoiqFplvXyixvRI4aHJa354Uk/WHoNxQ
aGrTGGZOrPFWlPVQXnwxcMPtOdOfkA5Bmpj30iEJ1DZnA3X9ZyWTSkpHewPLLeRnqRxIrEPUHacx
Co8NQyBL9ljWLJh9RaTFbh6jOM+66WRvMqK9dI8d9+qJHQJUi/MN5yI3WxL47eIrCPSv7NoWy8Bx
uh3bA/zDIMdClDq9NTU8TodWAAMqOdea6ZNzi1DFyekKHHffcSM6Oq3t58fUl5wue6pUKIyYto2Z
+WsA9sNIhrbhADaqOe/6KjPxcC5GVoV4S+ichPRLYNjOCuCo9uiuyWKbdS/tCEkBSRM5Cupj3aKw
JrIoErCrNusH2cnhiXnCVRAIESJr24S+15JJnT6DSMMu7Eyze/Xh0J0z0QQiGgOiB35cZcn8UsSX
3tXDmEleDjq4vYOyPhhZudAlDdn9r4+sshk9t96QvgIafm9vksFvreq0Gut4EUqaLoMrfj6mISR+
8v6xAM80WFHzNNHq8oBUjSLCJfkeMZRjhUUEe3Rr0QkJidHWXI6XpAh+xpFoIl5HvDbQ7XM3b11J
yyvW194dzsLHVlpSqWAqvv+2ZEr3sC+pSFRpoSy6c5/yDb5ltAKCP7oLH14fh1/8w6SP40lhTRtl
6BnsCxMU7VEQyKN49RAth5o3sOSg/QaYGtosufVhJ/fPie0xup85vPCrcn7yZQhyZwivlyT0vT+E
78Ef7ccFzw2IBYEyM0ZfOCfeFnIhB8/es/2l6BwCT+OdfNTiiBtIuB7MvI2MB6BE1g00m6MbpVwI
0Em+yyqoyVrDesuhUDavwba4arLw9KePpBkOuB+S7cohzvHdSq7yNkO+U5iDTRL9qPDJAMP/m6KZ
dLYUdfx14ISlDnpw6/YwQ+L6HBmJoeOCJWvD/MZKuxZSzv+kylREhJawS1RMOug3pnAp1X7Ki/NH
pd4VMF8Ro5yQPaDV9JwJwU7AM3cqXIIJwNO7eVeo70hbf3C6T7EAUwH34KBpqfowkF3cCOHobNaf
4eATCERrHeb8taBDDYzVJ55oLweibEpeYIJ+68tslw4e7OZuQxwa69hix1/dWdWlQqhnvhHml3zY
jq7cYP4wgYyUaTvqo+6pI198I0XmfCEOSYrYd/D5X2dZCJvrt8odmxSZimqLm7rHdHtlWgv/ECMZ
IEX4AkBktdplqo+aBVbWe4LDo8bo7IGJjyHuxcpl6ZdTlVMX6id8IxmR5wk7etuYxyhASTauuClN
cZcapFcQh8/7vwh5Vp4RvujdbeTbt6ZvYy4NgiNNN9ccoq+oER3HzICGoah0ght9UE++cSF45L2P
Ob1xJzSPTr/711Pu7VhOny/O1liojYOMTtKjXVaOJBM/JUDkCEGkGKzsNcc7KfZcJ1WaV7TX0dm0
Ut1VzdfTf+Ar4XzbxRoy/HJQUUFVN0qthOFZLV7qRZzG9vGpDkuzmu6vZ7qQlQTjRSMRVCcGUoZM
DmjFF+kOIg63wyXEvTywCuEPIl1qIMLu/eMJKbxPpzHwwhUqrOWhHzLEAQ7N3eHWGE9tgDfW65pX
V+YfILU8Abc6FpjQ9oibsj8Nu11kZmYAxMGE3C6i17MHL7XOCmOOggBrfokyj3TV4Qz0qjWO2piF
vRtl/+N4qOvRTRDZiphdZG93RUwFbqQRZjeIMYqNMOkZJDHKb3Lp8I7Soi263pfulzQ02qr0/afA
CaOZzTV6gDhQRKofVQ7H6JO4OoeYHWcW2z7P2IJoTkJXr1HRXVvAN9vhGyymmVG+eFPOyh0XkenW
h4rN2pJ+HPgZAkPpqH1lIuj5rvGv5KQvsyaxTup61VNVcIDYDbM7dF1bktNAawA6uaAv8dhcarDM
LCOgoObGNWAqQJlPyN01QwauYPtf3gLk4fw4HKKYv7V5niYPWx6KctaQLkaytUdLJoNfGwjunFMJ
JwFg9ZpElIxa7qk5zPU0Zm57jB0fY+sNKfJC4g8cHwj/FvcDKUaswebBNq1Q0m7q7mNNogLpn/0t
4KFfGMVUmiXR+Ke0B1/Ba9yu4G5IcLLVuQWuD/pUp/lAfj5c7zaogaQc758Hf09XvRTNRu0UMk4/
ur/bhRWYftvQYkaxvaD93sqmqUKEdFmlmFDvHoPaqI87bHaYJ0e2WQ2DjnSW4K4/vKcid73/qhc+
AK7zfOCUZAkpQmXvIn71IcGs5AQBfHTUTjX1a1VlkafuKfhdUp66FTMZ2Wylr2DWr+CY+nvyBXsI
rjwsiIsLMZJ2aVzlbikR4Wa2ZOC6rWWG1rUkSb1PzsXQYboDO3yRNzYr+ry/d4JCgoIxLFsrUHlk
Jt1EcQc58O81T8+dQeb1qqPi36JLAb2Ep4WkH3MMHGyxho5jqMsch/x2f3vEpwarqxlro07KIk6n
s//g8WSUvhI+XdQz/NH7hvAj4DiEFb2TmlJ/C8RNqUaxKGMHMOiaD1WRgv3mfnuVVl1oulOkYeY9
YXpAgja2UKINsMrzjo1hdZ2YVQJgNCN63ys4eZIdDheG5jBXEJq2rpLNtu0wZH8b5O5HihBOtXte
ItC7G4fJ5Opdh/Gj6t6qR7cwt8E2thGsTSDrrlMRRqcT4v+5HgZHMJqv8cAOCb3cY2ymP2zI+LLh
qAO0gAXMO+xAxyzF5o81WiUii9WtOTVRZ9DT82w+NaGNjIWBMAeqb5hN37i+uA1NTsH4Q+ZVjIRn
NpD2buJF4WBtecJEVMxiisakyRiI6LC8sOhLnPKlD4UNunOErzxm4+3fXT/jQV4y49/nY4+7mB7B
viYW/cBy6EfLacS7QDJOUB4sm8pzw/ODb57nlhmI8Ln3zTtHwq89ry5Zh8LgxDDs9SyE4hprgfIL
OuWU7SosQR3zBEkkhvnTbDR6pn/l8kJ30VmPn+Nlt/xAIejbwYjvpkxSwbhO8xvzDJ9g3klE8D6s
CFDnhp6QTzas99rYqdCenVqyI3Gg8oBMF5hOv+Z8dytZnQQythYSVreUOlP1rNQ0Lm70+56U5jzQ
slCUl83iquYIgPAeL7B52rcsfCGhBbxRRbgIYkvcJeTjJ30VNI2Q3xUFeHDhvEwAD/Pqm1gpSnuZ
rkeCUixz42jI7qhIafSxIAXCfr9GuSBNq52YCmFXXxPwt5fcH4G6lN0YH9n28QAEztfJikaMafQh
Nxe32tK/FBbQHloBzSalLU+ECsGqCDKvRqjbPKv8TcycXgY4yicXOUhrLG+d664MuTnk1L+q2kR2
LbWbObs8Gk6Yc0eLOZrM2HUtqxYTetrop/RgZtt5aZXhx5m/DkXYFIic2AJhE2kPNJ0nbagAmUPY
XPjCE0Fq6B6ZKFxGuxRgHUNCttJTpFfGOZSmHRK6htQ8iGVERip8/a76iuxLnz6ST+mlQPze36Gt
cl5+7Gj+lkBaGtcjhUk4gjuW0pH4T+IYQYUHESzlztcPrOTNvNwW/7XpC7423B7+/fZzrj6zvL/q
QxjH2WP7+VRQAXDyExB9lDKEl+JsLlU5mV9F4oYbfigBmwAYdmtHYzJWk2Zxbj7fOmjdhkf2PaZc
dBEWYR9Dvab4zXhLicF27l9dkLZPdsTeeTMErho1nGImeC9gVUjUOOQBkeNVfp/X9ct0B/J6ek8W
NKMir82/eMxuEThmbWz6om1tDbOSC5+KcsKym79bbKvXKx/KFm1qh2GJkFD1Onar742lJXzEWPkC
2t1uXw52Rk9Tytdxo10CrYj3qlMwws66NcDg8YUHFjCfq/1IUVeQiNvlSEiN1RdLNP3pTns8vdpl
sLGyHOvb8QohD68ppbgWjpW0fKl7rrJo55YOBMId06HDoVX7UEH4n+vDXdzYBCtJB3C9ADlQB1Hg
IgidbuHbI2LLJgcL3nTEDKsQ+oTQGd6P8EtnVc4kXI6lWmfpCJJl1jCqtqgRuuztGeC6/GsQdi4S
3T+iarItVNNcGBJ9yU4xaCKhOur6QH7HlBO+gyuAWvMsWIx17JCy0+i2O/D0X4FYQpqa5062el+Y
jcH+q9ITxWmrB4PKwbG21s9gKLV+tYzgFqGgOvsoHnB82OZcYZ+kkdIziqlhstfjX/92lecKPXvw
Rsq6cfivRRlVkeJ6+kFZ2bY2kyZ8RBA32CN1FEU05QnYKlC+wySjxdQH6pVkSOFUFM5QkzszdEXF
GLdBORE113WUqMsI4SfnMi7u/7+FX7884swlKjao5fdY2MNirAkPF5YJ2Tyf9keQZe5ncocRNELY
9e8GNr09A5fXjhwLYmTsczeyCxvwtuEOqjJqjZUIFbmrjD2xpVmEfgmBQn/sZ3y/Si3121yQLTXs
R87za/wdfh0nFa1FHuXrty220aSGjdfbJPRItRYavXTsypaa0NPtqFbQVBmEcJ2pSw+dX2rK5hTI
mTsfbEMpVxXKJV3p2gpkp1A86KVe6AIdW3LE3vEXfoQyVZvZI+r0frbFZNV2sTCHbDkxHg/I+l8q
uUz7d1HNY4jfX18iEOHBISZ0rHIQvhrHYyrZQwY9lmzEcgzdbLpCs7vSlJmrJjxWup2I1Qkhw9oT
if72Rz+hpScAn7iUO+T4NOMGUaszQ2s+6aEu0HZkI+O40Giq5D/uB/vfg02gffqfzbpVCih27+ya
Il9WoGpai1tPJxbQm9Qe8gpz37tns+P/iuN816W4IiNWG1wr/QJwzquXIuRBv7L9PrNdEm8TRHa9
vqSPeLhe+cPyerBzaoh9YaP4uFQwMNaBsE0ENF7Q7XpHfZzbInbCn5HaqciE7zSlL08ede2TMAKg
N4mc75mCeqleRoKsjbSwtf7fuda0BZGhnPwJhTRNyD4zp6Cyhg1IA8AnPkRxzugbQlz3VcySZ3/d
+hGsANYv0fHQAWWS+3orYsk3rtGCDRtXsjb0agWYv8lxSorpy1zHfJJan+w8eu6b4XDcBnyKcx/5
MYUrtDenkNorLx8iwD/PIk968xBPudCMng/2lE3mfYJAHzeEZaIAtx4fNCXBDmVNfNuzmKpdIM9T
1JkaF8lYUad7YphZF9yRsBIppZRWXGc9b9AQEXNa19E7xeHFcux5dwpP8BLiVPTSVq8yJ4B9ah+z
0llaB7rdpbFGhdi2NoDuzVpk0If9+c2NSJbgFnjvoFYUDMjO8o9S7r/U63qQn9Ko/ppw7b2tewjv
OEBaPgUMqA4cVWk+aVx76mUdH339/dvs3fhbYq2X18R9W5uaAYRcBFMwIVb/RuLI/1CivuzPZcGW
wSGzVxNtup8318L2saOchmzinHhWjTR/IWwyJjEPunNZhREI7EqJamOYsbWLhqgtZcrWOQiCBAIn
RsjntWuD3F82DJ9LHidQBZS4haPn1XDv2f0IvwTJfIoiDzrsnxc0/P394ezcfaGJO6HTpmMGYuYS
d6OjvG3q2hxPfweXkgWlTymyCljaUrMDK3UminBgoyLaqikFlQ5D55wRy7l1+d0IBxZrL7MrkSze
Iz6KsiYX0rpFV8ccUX01l5Z/C5o+A1R16H3jLFe/F2aZ2MqNVBONNftX4GpgH/eE9nJCK2gK5BFo
9pM7CjB8AtX8n+m/H65s+9Jo4D//6m3xYjubvQ3gxUivJt7mAQBifmLKkjBQTwYZ6/U2L+Gx1wls
rex6tNtxj4kC79pCtS/UUowdQsUiHEsCJXEKOggpk0/SPhWi8HdBqC7vmMOEXQ26/tLtKiumcjAN
8GB1VWR1cMXlPXptYS1OZ/WjzCmJw8bgsDRA14kayQpjHJXeLVKgEh4TCWLWNQjwqsuinki6uMmt
Ak8i1zqKGmWkJaQQoJvh3XLa4UNU3bg52bQf5W8hYG2BStMEI24+JhcBjh3Z3+vMnwlSkAMha7oq
cLQbGS4YMqTyp6GYZqxf1z2k1/4z3b7T9ImNsNobL+lsWORBbIX5c0JKdGKZpAMIBPKxZdN5ERZa
N49R7XKOQGp6hldqs8tazDc1MTJcdZS9IXf+jx43qxEj2rU6YtqufEUT/MvDuBC17UQMhmzLZQnx
If6q8+tFPwUnXmbB7BWZeTv2P+dk+rAuq5ll8q42GH7UXLF+OjOIKDkkeiiaP+I+gBTnM/m7fQDZ
jAAgmYjzkqn6kO3O+MBmGGMluuu5Y3c0d/tVEtR/NcNSfXv5SYwvr+rIRVjG9TEXVL5iomKVE2r3
L49QKRKbgopNpUuOENnPWJYlU4PuxQ0XPdAqP0qQMp/mJmF6hYE9iEBzOt80UjDbCqxeqRHFGhzs
OLs4pnlDiCTADk+3Tn5Gc59j8Hw5U2nnJaf3r266kFuobnBuN+F5YZPsvLhI7Vzx9oNc3YgigHnZ
NchGweOL/djF4zBbrczJW3Mgglpfp3wwkuGlhoshGlBBRqHm090QbrywZve8TbOXRxrK2NAaCwut
WBIglv6IAB7I2K3sTHZetAFOQchi9oo7fHvZd3Hinj4RpT/jwU1ohvjbSAWzcW4NKV6JO90K2udc
6pml0cXwWDtlTJ8RCGNI8+zIiaHONXXUxf9hpTjUDoUZpi1r7TqVhUyfAqaORAU+0slRFWO3hFfO
uiygiVn4zZzUb987MIuLdIJLFdNoEMGf5Qg4pEYIptdtqmQQWEN7f23PshfxyMpbjznRBhXPvLoa
QFR2D/cVYtKzYcNjFT81XEhpv5iNQIP15wEL9OitLJJOgLw4upQC9gVuEOrue/DxWEPdzSqoTr+k
F1liw+HxooMz3YJkSWidolsfoX+fUKQj+0yFPKywQzdrYjUq49Nx01rOoNzCLApzJWClDayKsJY+
CqXHG/CTwxRs0UfC4GvI9DYJUXlUP15ytyTBCW/9yN5WiNNxXVHVOnbYDp2sTZqhjWxMYEbBIKFS
GcoWGNkjaY1UpH5yPC783JdDS+lewTa4uRDlrO1KrcmHfpNzyP9vpEtlxs9iLrOZq3wZ7bdmfKBa
BioVINrv8uOqe8G2nOz218gVlIEN2VnNLYecM6S1nckqgMJ+gqPM2KWv/DweQROb5cCOV5kkt7mS
aUcW3ElolQQEffBf6sTFb8hu25oOO+aDVRDgpiBUy7E0pfg9CR2GWjTIp1RLng1LImO2PAaAwtjD
efLE8qliY2lvg7icFTwuyPi2+UQEmLmEhJsrDVn0cD/rlJwxP4t7fe5nVv+9d44vIv8Sh0TsB9w5
JNuNt2GBkSQIVZE4l28bTT0k+iYjgGvjXCr60CcQo/bYpxa3ZWaWkMXISOX/A5iNlOJAUvDKbOds
A/FUzyljLeFBWbfyYpD/vf7/1zceZzfazy21+MvtV7h6Q/D3JzJ7tSow0yoDT4Er27MlMHmcY52f
IaGlU0SwoNmloSKN8WdLqYncj+tmDWYQVifMn7Sysqzme13Mr0okcLZhp6K/HXMlf62YqQPuehFx
Gd1rYcLKqp//OQ7c7drPZj6jp/nC1BGBexHMoqf3eNMZIFW1GgEkMcSWqVCtCj95a+Ctugbc9wRn
HDFmIb+TBB+8XdSV2sg/Dfen8npijpLe33BBY3FuKRyOTrJpfLOUm7dh/o9tjjW7tjLiNS7+r0fa
6iIIIqlc21oOhBBRk2r25Rm+e1L3MpE59Uipd0pVdfBMMhoalpfFKsRo3BQYskZYu/1wboZPnMw7
csHyX9edpVq/YXQ9EcNO7g8yuk09FDiJBP+LMoD37K68BYfe1IDFcPZHhwj2RwQEzzK2z8gS5sHi
PYdj+HXTCTQ+PYJVrLpiLqwpL28KzeksqRzzvPDexWVnbDkJlk2Kgh7xVtj9kzv2NpVTt4HMGagW
B8TRnS1yTzvxtZ0k1aRU1f2e2fFJPW4W6xA08P6bmPX52hzaSK0me4EEFcYbS2GH9O42mCqcsF/p
Pok8WzqtjnD9uhjotrD4LnbqbsWX9Jyc15ubOt4CQFxDMwSBsqHgYghcqJaffzdTvm4vO18AJ/rV
ob9zVHi+cZaB4ucViL9Xo9VqsYOc15SpFJbvz/o7HDqn/PwuIgvzzCWeBAu7Sz1gIVs/9vYtBM8U
Z1b8K4UL1rhqOwAEM8aVxSNylENIDc5vMEIwq7zX7jCdqxAqK8MJHC0E1iuSYXzhxq4bzEjU5VK8
WU5jIeMP8MzKC7iAcpDLClVUPJHmrcFkDDAB8yiXo7wu0fOs4vcmeREkrp+Qt1KMZ7efKaBa3P5T
JLClENVDLuEmmIEuHnAesjpVvcc2ib2L0krUjXJV9X14iqw5MJSgYuWIql8D89DsGxG8QpAUXtHI
YoXOuMtV4m7NxNv6rm1a6abXL+sp1lMsujD2pJuvW+MvtIhZX0RkWIuaBVIg6iBybRcDe3j+hrHg
HA49gktuWPoFWIMDeibx16QoayB7zEZV70nbgaip+50RY25zllnEBqcE1FDMrv12ARy23mXnc72Y
LfYg7A1EvuV9SFpJQ4LaqEqgsbytSHVyZjRZvP0KrxnREe+p+2UkEpQhVC+amjQFxhcmq9P8fXHl
HxrcPGRq7kuRP8UYmxO5NSI+ByeLqpuLfKkrd6mQJt5fgm0ryhboKAGggRSCWw3iBnpITkT9dVd7
dF3NoNcuS7kpbuPFqsJz//38jJ2VYwApuuE4Rq6QtiQjMTRuiBZiHiFRK+FbZ9hfn+GFbFWMUZLx
ofVLne//CWCdMWV/qrUTSYSa+0AXX6+/byty8Lf36hYbi1XRfFmyJwApENaTaz6eLjVnbT3ZA6uc
w2DJ619zLqD/ungbgTTb1TGY8+GW0JgRyILj8mY17AtcMOZ19yawJZws+j7JHBR7x1mWt44reIZp
vxtRpbo1HcLKGOT5Idy1ucXkLeEILfpRz7HD3PK6WyAj3VlgT/NRCbbFpOq0OOc6d6aIiejILdFi
K0htwo7wIL9wEts5dhhaO2wytKLV4RBTDo0bRBozXZIw4AW9mukEWw9KBFng90L0KNXVlE5/4HJe
Tnp6mnpz7qbYvo2JDe2Pqk1o0nTxW0yDLrnhJRTI2ZAYerYvX7IssB49hWoNjcQpdqSS/IMHHIex
VfiUnliZxifSlIBSbVs3l1c6En0ylZv6yi4S3yj+mSwxBUVjoAQ9CN0XxE4ME40vznWjpOdrEfHQ
lE3GvmZJ8OrB6UNtURqZx4MhBNj6Z1hbBql7gdKXUhAyDCVS7M7LVlb1tPg4v2Z/Q0PkNj1MbZYN
VzSy4IBo9hTXFkTAeuNM/hY//z4PGId/yhIhAAuM/9nwd0HvwDqYbOmOKcNYtNRpPtqT86yZEMgn
jWm3siQSxAzlea9wZi2nIkjrDA/3Yy8fY6Qj6Tdj9FbNRohJom4P+xhFiBPfU/Pq5eUXiSbTXcs3
Mua8lmwLbgKeZRV55vuUHuNA5LN/t8+2XX2YW2bOy3q+OBI8dCj2fzm+85OmMHANEgliu9CK1DAO
ya2vJ2H3FyrUjCNQSrFrQh6oWO81z/HbOVT8N9HP0X5ymGql5UGtOitWVA6iPnvfwY3Oy3Z2q6LC
4UHOLzIuDDl42mkrv7OvSYKYt51eMIOyp71GD3jh5mrzldFOO2lU1XOrmTjXcO0sYg3g2jnnfhkK
4Gn10x5k/PLIORUg41uxNKe6pagOA0GSLZCR5tjqwtQejibzZqO3O0kbrEMarFOl+l/8AucxI1R7
8uiIQrY+sVZTtOJwfMfu9hyJjBiWXWYCPIpRNkTRi5RqB3J94w6IkU1oNG7C/uj0caEBwVul7jm1
98W3KrT7blk71QfaHNfRG8uHhO3G9iMe6TYAcCW0hh7QjMIjDRUytw5Gg9EQ7/AG3gz52T7D3SmN
SSDSDBhSNMnziPEbLGkjVOgVp8zLtGpDJsl4T8iIiT5doxif2Xi+ukVOxP3/wlAHlmaYcldP4tOi
xSIqsFtH17w3lHomsm1VpWwCO70bQ57qYGW5eld959JhowfYgT7235cZlF70bG783tOHSyK85e+w
LXP5DKrEGGYE5YQLk24DtqI5QxopW7g34tawEozR+4/5jqMRqIsduj+9rBsizqFa0EkQi4uk+Wfy
j0oUkwi94BuGMLTmN7f8UncR4q0Oa5AcwFgRJRY9P5feipI9hTKFxtOb2q82EzgMQVbaGNXTswtz
g6VKI/pDDWuKfX9v8/tMTXWwqm5PUKf1jh+hozflLOLywp+8+MgZuJaZuYpJmdO2VXtf2usGtQ9x
e7IgEAra2bZCoA6393GvqSMlezNKAlQ1nrXF0B1QTPXPfeLktunsH1ZfruBw5Np6TUgKpJ5DXEZB
GzQG8DkQHeftGS5EN+Aevp4uR8vd7PT7L7OxBTIa88jul93GceF6B2YgvFjrFB0ks6GB7LAZg860
s8ZU3+yVr+aYi+UsQK3gBN8rMd/yWQiHnwUAMd/Cq1iOSJQr38fB6BD+6rsJzHwGp2xSi/Jcc6Aq
3VU9rsMoHUXbNs5jxIWVpdEXDvNFST4uJSjj3iv8BTzParGE/HwuSkgGIpjbS7P7cmtR3KZbvuA5
BdNUzSd8Dpezt6SqzlfTLZlyHP0ZgiuJbYFiUW5CjYGb71SVHmiq7dNzkjo2GjAFm8Ah8guyOa52
G0owML8zT6TfKOHnWXes8ixaxAG5va3Hm1dlbWKtCGdXRXjYXX1L8jBxd+BL+1VKXn2SEs+U7p51
d0RA4SND1I6vzcIz/7mNjIrvmmmU+aDs6fw5xntkiTHgF7BY0BLvQzZMuA2s1p1OwQlsUXpiT+GS
A1OBPx0aTpISxJPudTsKtdiuG8u8HxLsLqraG05pPgNG8vkEz7um26KHMJj87ADuJJ6JFqmhHFFB
Swzc+c7GTs/P0ZXWicsrZYYvkC2Zg2y7z8/6twFsAAOKaUb+j8l2zQgynAXrjImuKakHnzY+FQ2C
lH07QSFePZnzRUC1RJY6UU1nhAdP1LmcPHrv8T43RSA3ZL22mztUTtQe5xRp+SdcnZxtwiIADeN3
2mNtbwvZaKou2O1QymKyDZYYH5qbpFzseQ7ypHYw+eKPJzZ6aONWfmxA2JatjlTfcN5cyYyCgw3v
rSn7QxfiD0zZ1CdQTJw8H5XIUjcf81Vv9egEF0HdU11T2w0J280ujrxvlpEhRg9eQcSoZ/W2IqpC
NyoxbY2PD4tBalkn6+d0AHnXz26A9bow/R6nSa+pXrh6TL5pd3cbgon4aOrxTifgLRID3gBuGvdy
Ak0Olmu17T8IuZYOBXkXRxJIH9K3KboqYPI7mRAqilhIgKT9PlsqWkP4FZ9wYEcPq5/P0B5KEqqD
yZqYh84W2y4gYw9kElwB30gCduzWfbjIXvjsNhaTMoWQkcdP6YprZkn6UN/znLsJVHSbxNrtkbs8
7w/+Ol5MhdY438UIU1dKiDzzmzRJnKfF3H/esuld7EbUg4c7Bk8hWdCbFwS0+pSNFuxlsR8ea9oG
cJNObuQGTCWRn/RzB7KJc/8ruiabkXnDT4uqz9Mi2W8WVSoW4Zxew0W2VKShX6PsVPnfkGiksYQq
SeUpOjToOiFvgi8F/2+XLsJgHLEKJsdqGzktwG5FgPOZZnygmnnd7ZYokLM/p1Kgp8VY
`protect end_protected
