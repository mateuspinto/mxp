XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����+D����"HpUb����z�KV�N���nJ��[�j�	��`���]��Q_��x_�۷��R=x� ل����>I�w���#[[��pLr4Fmi�g�6�����A�L�����;'����QmE"�J��W�2(j?�U̰�T�
�#,��^%t����tTR�mP��$��H�
u��-��u�և����o [���8�s���4|�t��3�4��#��jݵ��9�7CƔ(L�a#g��ƁM�%��C,�;xLvOJElx��i��9}Zhkv}��s�4D:���w�p�,�L���o�>�-��+ aW�?�l�ª�MF����d���Z�i ������m�0��rS^S�Z7�:h�.N�# O����p+De��s�Ib�:�#w�ň��,�
�H�˫����X6��P_U�7��u��pҍ�klq,� d��;�d��`��tb�F%��Ntr�+X����ٸl`�]�.=J�h�W��n;�+i�ϕ^g�o�����F!w�� ��TO�z�Y������Uz�wJ)��j"P+'�Ε�懠��+(��!*ʧ���h�A��sx���]���&-n_�&�7�󏤝�U9?@�nў,���*��e��4�,N�����=	U:�O!n�J��rF���4����wVۍ{���R��T�T��l�Ĉs���%J����1��a��Z���y����+rՉ���0.(ʸ��O��QC�V��XlxVHYEB     400     1c01���8�t�c�l����m�?��P!�|)�R𓧩+��,��o��C����'�{]���LTsg�L"��D�+/��9��*6S���z�Z�:�j�?D�>;Uq�U��$�P����ϡ����T���ƕ���d3,�W�O��s�cuCw�GDM��v�X�����t�C�2=٘������Q��^�I��08��&��ONH�gw�C>yU�:�A,z�r��1:f�J�;j�Qm�%p��kP)�Wz�)��xF�+�fݲA�:�O�S�S�i�!L�U2��^YR릐K����[��4 �
���+2Y�^�~�ʉ'��-
�DVc�qW��"#b�;ݼ�@2@�&�D����g������S�D.�K��ʥ���8Äй|�.�u�A�J��z�{Dg��X����1и(T�`��o�hC]*�'���ظx���XlxVHYEB     400     180�̥qt�� :�$�r�Z�a+�_��Ðt�.���k�bm-.6%�ϔw�@$�7��'UE�#��z���åMY�<b�\E{欄�ye��y���&j��T%�K3a�Ln_��b�a|a�����5xm��ҽ�Ǫ�5�ݮ|��M����Wb8f�� mW!�&d�OL�^h ����_�*���2�쾣f�M�&�M�����ݮÏ����W5��H�H���� &s�7�;�B��0K
BM]P��!�v���ȱz�ݱT;�7��\mH�̈���8�k��UF0~-��� U@���N ƉB́��A��c)��
�x��z�y��C�=�Y4�^�AS��~�j.���,�
�@��:�N��բbCb�XlxVHYEB     400     150�2$˞k.�\�!᜵�b���X�7v�%�M�w�W��������Ziղ����J�#8^FK��Ì�����b��K��͛M1��;��7re%�q�9��C8ؕ�"u|�P�Z)8[bqi�������ih56d[��M��ez7�0}��
N�#@�w��U(�� @n,on���B�t|a�0�(�Ң�v-�4�]�2�MkA�ӞS2�_�y�u:�$2��ƐmU�E-/�U!����՛nJ+"vP���j-�Gm!!h��޸��Ԩ�OW�����Đp�U��6��t-�' �@�"~�����@�҅��\���X�0�׭؞����)�XlxVHYEB     400     1b0	� b%J����p�o5�@�����ǝk�;�߈����=����]ql�MKz�ka|]2]��՛N��!}�r<=o�Xu�����	������Z{� �h9���b�5�UX��� �y�A7�Y��)K5<�J$��]6z??��3컻�O
sTvw�5���B�3^ �XQ(�1�~��F(�[���9��<g(���ȋ|� �*V��+��V��M]�"iNK�b*e�;� ���7�)��	��/�o�+��4]�?�,�J����ӳ�Q.�dJi��%U]�a�"P(�!6�%��~H�H��Jf���ZV�_��?;R-�=��7������@Q%���YI3��^,�M'rB�J������x����8��(�FS������1I���D�C�F��N�����5Tė�U�=XlxVHYEB     400     100-����`̧�`mb{;�l}�Q�P�3 ���n8���"�@M���z�P��X7��n�����b!�y�=.)O�n8���� &rH����*ȱ�k�7>���wo���
�Q���ݦ���3Y�pG>e�*m����'r����d�WtP������+k54rs%���<C��Z���t��	������yM�6����L3W^¤#b��rO��>kuVo�2A+���c+��s7��	u���VJ{�XlxVHYEB     400     120Ჺ��/˂+X9�C2GG����fT�	�O�|��F#y̱7W
��x���
�LW�"���z� 3���֜	�hw����]�|Y0�"�!O�s��$r��7���O�T	���#�J^���]�4W�~a���|�����F&B�%Y��b���/ )��x�\yi;t-khSO�m���W���J5��w���r�2�4I��:$zA��|��(��Wm�5gT�r�`�&FcA*���٪H�y�S�3��g�´����[v���R&=R.Ky�����aJuC��kXlxVHYEB     400     160��������bCK�gA2?�M�[��[n����tL��Xݦ�̲<	Jϡ��l�E�}�淪��D�Ì���Wzs)��``�tg�$VmE�L��	1�i:Z��f������	]������[��I�6-;�g�xl�c�9yr�m���$}��Q�;An�1�*bC�����z*��௓�����|�C��,�9gr�I�����l6�ޓ~��ԺA�z|�	��ݹ�F1�FC,u{����L������3��e��'K� ��p��(��謭˧�	�k��z�=9g�p5��K���[�x�ܩ�f�����Q��W<�P�<
���6xi�Oǚ=�����w1�LXlxVHYEB     400     110i���J�����:�ƝF����fF@�P��eC�N$
-�t�M)F�:k��ë1��� ht^�e�S��³���D��qe����xtg.�24ؕ��e|�(%�e{،�+��ȡ\k6s2~c0Hf��^m��e�[�?��XF�x�JRz�ͅ˩��h�[RxPM�=B�A}v\�����,��N�m�C�������?��t� ~�+�!B1��%+ sR�#��m����.�!�,�g����>� �[5�t')ӌD򆨎m�U���C�XlxVHYEB     400     100�ۉq6{\ws}�A�F*^�kt�\�7q7C%<���:��{�ʃ�+�@�q%�SL$���� �j��6�g�P�%?Z!�s��'�gzXW��V�fB��XI4'#qI
 )1��]����aRR�N��4z;!Oz$�A����'U <
R*��m4FJ@�t\��s8��H]���N�4�;���֧�M���ˡ�*�6�Ϋ��@d��D�c,^K%��{y�H�H{��r�D�����K�uI���Y]����Gċ�XlxVHYEB     400      d0��H�w�2z�uYq�ж��o:z�d����X���V$j|�'�kބܰ�����G�c7��A��;.���+��i�[����,��nX���6��<Z�:߱��lr�rR� �}?���k`��E��>|۽/ҡ�b�i�ܓ��k�P�w��x���I�46��I�9����}�Эg��^��aRuk��t�KŜf-�2�XlxVHYEB     400      d0?5:�@������3��|� �]��ɢ�����@s<�l��޴����n�u�L��1��;j=#�l��\��ͭr��V�g�I�BK�KS��^��`���BF}����&�f}aس;+X��h"�s�@B+�	�τb���8?k��X���ʧ�o���B7eO�k����"��5?u�=Ed�7��8\���w���c#"!q��U4XlxVHYEB     400     130f\�8a�����QB-���*�Ьͥ87�Ơ��R��� �3�#�ɻ�S�-py�U~�WWw�#>a'��r��d_j�����7
�B����8$���8�0�r���f<]��S!��^x>9�#��1�����Xi}�)�����m������Z��;&ҳ�H������c�4�w�IlB����|+�	�H�k�|4}�9V$�94B�s�CZs3���q���y�3��۪���m����2=��X.a����qR�SIf����S�h�O7:�qk"ʤH�\|�V�4��_N�k��uXlxVHYEB     400     150�sK窊.̲��yv�Qq�9��gXA����ojP��jdYFXv��IW���DG���	�ԐK`Y�<�g��?��scp��5k=vε�n=���Y��I.����k��H"�j��"�<V=��T~f��X�`a�|"ESO`�"��#��@�q�k�zpv�a)h���T����%����L����u��z��%}�����!ׇ�U �6�K-���j��k��u$t	1�f����k����������/�R<Z�8N��11���]�&�u[u�G��tL�"HE0l}��?�=i�J�2�
���+.)1Gć����F��x$���4|3f"[[XlxVHYEB     400     170��<.]��xo��Ɣ����y�>�@1�K���KV�e��#Ĵ|�����?�����
���i��=�GE��/����[qmΣ��(�x,�[f��[� ���1�L�X>�;�j�����jҵ��'��~H��p�d�����Bő�IM?�Z��ߢ�~M��{&�X�����Rz��|����mOe<��A#�Ƴ��}�G7rU�s�I>Q��gtb��u�O_^smUU.k:�ZD�{k� _ՉIڗ�C�F�����f �*KR����W|��Y�GA�\k���VfK����Z�E>Vu<�ڎ��$ͫ��V$ؙ�g�0{�)�������"dB�8;p�sv;y]��>�u�ʪ���XlxVHYEB     400     190���S��}�9v-�E3����o��k�u��� !e��e��+r8������
�/L�,�������O<O_��OC�Lb&k���6��d��ݹ����9齂�x� �N��i�Ħ)o�����y]O����@,6���n�x[�T�Yؤ<q �2�����P��~-Z�0����X{��4Fo(�����#o���k�A��'I�'~"�v������
y�&ӎ����ld+<�ɛe�	��6�Va�����Z`y�?꫻�Z~��%��!���
��q���t��M��vٲ>��}��1�s����L�q��R��<v�En����^��H�������%��5���ap��U(Q4�j��"L��F�h
�5t0��}�i/[lp�v2OW'%4��E���3�nx���XlxVHYEB     400     180�|b��Lի�G��0u�����!@mSx�6��U��ұb��4��1���t�����; 1+V..�Ϥ3��&������ql]ڣ��FY��a{���ǭ���g��҅,_e�ŧ��H�[���q������Z�X�j���C���c���;)�Ek�vQ�U�La����ՌbS����F5u��`�ӌ%����"��l:֝�L+�3{�_(�?y$u#c�M���=+χo�qj������K;]==��F��װ`�,��c��؄��v��0�sX�}z]X�H�K}DE:.ӂ|���b��wS(A������?�C����U���F���n�o�k7#2�|y�񍛁�iyV`tĀW��|YҲ�tǢ�XlxVHYEB     400     140fՎv�l�'����J��I�}d8�8�3���Y;��W}.�1��5ꖻ��܈�p6j�ze-��j�LnL^��:��)I�L$�]|��\��!�[��@�|�S ����~��o�A��>	羺J�ZI�N�]o��B�b䷺����	.
ЏC>_��v.��OJ�%o���FƋS$`�\�t����D �eY�Y�g���0�y�nPZW5�_Rq�0̦�_nj;�
g~E�b%q��u�ۉ�����}��i���3�Ū�p��͝4 ��#���nl?%����a��A4�sY�,*��
ߩh�77%��3ҼB�XlxVHYEB     400     130P��%��CtX���$�V������؄Aok�2%�҂������_a����l�5�3~|Ϣ~4�vz!��������U��k�0��X���&�+r�p�=
�i����z��l��U�dp�D�D�ٽ0]��������b5��Q��B��r'�;E5�\���Z�}P+1��g�<������v�����#M�ǥ���ö�%��Pr��`�}���'?6�6�JJ�uyP��U���U�J����L��h�A��m�o�Ck�ݨgO4��tz|���B\0�4L��/d��-�Op�x�KXlxVHYEB     400     170�"�he�db���f�N�=������{|)�HUȬ�k���b�@�,�
������\���q��ڼ�)6-�}�LR�I�*�1(�a�+��ݛ�:�dot Ȏr	Ÿ�QHV&��+������/~tlRW5&j����C+�"+&��Q6�� �u��ǐ�CA�_n���q�%C��e�f��:�~T��`n�R���ɓ�Z]����@"����3������n�D�	}�Tn!YD�|ɘ��DqO��
��RТ���촿�TogҘ@�������-6+�M�Z^�f��Km]�+���˚��#��{�Jߦ�����%�n�^c�U4'�\���w�64=��d��J:XlxVHYEB     400     120Ԏ����Z�
.�'®M��3�����}��w�	<�Q�@��Y��t�*m�<z��/
��o(/E�k�KA�7x����L��s�&��g��8:2��)C"�C״`c� S5�F�(&��N�OQ��!�"��Z
���*Wœj���̢c�*"�ge�3��1`�a�dFw�6/Z�6��<	HB��/��\wM<+�ˌ7h�P�-/F�o%X���8v䬍(B@`����,���i&\�Y���BÙ7�e��M/�[E� ���k|�k\,<��T8���b��XlxVHYEB     400     130#�-3�^�ǀ�EKZ����%�*ArzkƇ��s����|N"~<�����nl:�,�<�0cV�c�i������E��<~䪧���K|P?���|��C�/���-�ǡC��K�e4�Jl��A����0��M$E��Ja�Ј��*������Y{ɘ�p7'�M�1�8��B��k��v2����+O���T���.���nԔ��%js�J�Џ.n����r�=�f>�B/w��|�wP�#�_q4�*�j�~��05�B|q�i�!�Yy�����iط��]�gLj�'XlxVHYEB     400     140!�ŝ��Hܑ�_��/� ��M��Ӄ$#!;� ������H��Ī~)~�j��� ;��Vr�qC[�=D�/�nه���[������3aD{N1=r��8��M��w�u��"�M����p\�I��1=� 1�����*�v�������`Ǳ���Ȕ�{��#߫��8=6��ڕ �$�+pmG��	��-J\*=F`XK>\�9EQ9$/{��*�S^C6,�zb�]�m^�a�DY���݋���qa�¦�՞[?qAB�e�~��k3v&H_�:��D
H�',��I	wo
̃5�j}�?�1H"Xa��kFXlxVHYEB     400     1a0�	f�ZQ �Jذc9�Ӗ�Z��������[��cY̦ �7ڙWd�:U"��Y0�ڏ�n��'[��ǆx�)(i�O��'R�.��AsuHeh��"�V��\��sO�׾)ٞ�(�$y�k��h����N���ߜ��b��w!��.]�̐�Ē�nq����޽�1.':�5�  ���9Ķ{��LD�t�`*+�5bN�ԏ�����K�Y:�g#�)C�is&<�
����\|e��\ʿ�}�%�L;�32�Ͷ��!��*�Lsy���]�� ��ǳM�Y��id�v�� dW���;�s����Ǻ�`ب��-��]�8�pSu�JOa�}>�%��1Sd��#�.��Mx=..h�`O���|<��V��$+��ތ�g<uV63%�R�Βʀ!��쐳���AB7�8)�gXlxVHYEB     400     180I
x�m���E ~f2���ě��*��C��vdh~�C��gb%�� Q&*�JJ���8.DEk�M�s����N��k}�*���ÀY�6b�$�:��e��UE8KkD:{�� �����������$��T&�.O��E'���]0��ߵ;�M�5�=�]aSw湎ȥˉa�0��+d�y��`ԩN�#2[��/���v)hF�-��,�Vo9r�8���)H�UD���0w��'�4��0���?��ӡ#޼s
80IC�S���Oh�(=������ �G����.b�p�s�т��1���,`���%<31�0����؛��Zrh���ɻJ>���b1M������8/����j3�����y��F s��j'j`��hIXlxVHYEB     400     170�����8$Y��b��g��(�)���$�
8����j]���7�Ez�1�2Q����!Qfb�=�DWn�N��!Y�4������)�)�3��X���6����wu6�-���h9kaK��x�]!��P�57�y�h�W�Y�0�U���տb��^L�v�
0����#p��E7&QG�r=W��J�b�QZ�y����>`1��0�ŸQ1��W��a��#Ξ���~���n�fvǹ-��n6�=����F���(���2G�.~f�m�����:�?��w������C/�2OO�AW�z���� ���&�E�5�b��y���jp�I�Ò�K/n�=[���܏�`�!@�$!ґ��z��q.u_XlxVHYEB     400     1e0�b�D@�h�x��
]n�R='��p�P<�����gԋ�#���bJ#TW������6PR�� ��!�+ޤj�ᴕ�1\))p���#v�ѹ���rf��y�,��L���-�jB�b��yE��
�?Q���/���� �Ӽ�q�"K4��|�)�S3a�Ѐ��J��s�3	�[c
�RԳ�g�mء9��tc|�s��5����?Ҋ�d��'�uW׊?I,���j�S�Y���E���+�:Uo>��R7��>W;f�@�F����?���d�����3o�ۉsK��8�W�ȴ >푒�;@b���<Q�R���n$���`O�3����CD(��"Sð��P��fjZo-z�����U`�>�:0?|�O�B��p��}��
��Œ�7�QPi��y���h�˕A�5'/ s�l4�1D��9���w��
^�j��	`�f-k���kp
/�}����N�u�0!k�=�ʇXlxVHYEB     400     1b0�Ľ��9��t�Б'�O�[��|�w�g�)V����z�ߜ
~�c�q�$<Һ�+�<0J��tٻ�G�H9�f�f%u�+���|�)Axw��[�PŎwK���ʁqb	�Qn7��ȗyɈ�����5ƃ�#���:`����f_J������N.����:��R���$�Ӻ�ƃu"�w�?~٢��T�RA*�	;��f7Tt����ǢT��kإ������U�ݗ�S�g[���h��>�C�����;���fX��U�]�T�*�\Bu���ﾯ)�����"6,a��8����`	����R�(���0�w��덯����B�1���^K$D��M���I��nh�c_kC��x�/8=L�'
F�Z���Y��Eށ{`s�ۼ>n�ț$�	.R1�6��s���K#dvb��}h�UXlxVHYEB     400     160 �5#tսHs�y}����%蕜1Ӂ`�k�{=6���B�����8#��Ņ�� �J`F��h���]�cj?��B�.��p߅A��l��X�l���Wk[9��b&o���F�s�~+^sz�M:{��] �.�D�RT�^�٬c�QN��#{3s��l����1�;�)�Ib,z�(��쪓Й;��3�"[�Ǳ�&M���R�����I�����@`)��эd�'D�S`�BW�l��1jO�#xe^�Ļ�#�.^еD��>7Tb!��=�D�bY Ȯ�AX�J�p��Fލ��\I5�̏��<�o*L��:d�ľ _ӥl�U�[�9�����C��%�XlxVHYEB     400     150�]�%�0�Ԗ�Ĺ�=j5�҉�m\�u��,w�I�����+������;D��
�q�.9��\��N ��yy���8�(�n���)w�mw����U_��sRM����)�|7���2����|�絗��rE$��Dx"X���淪�݀�K�?���h���>��!�]�,d\S#_%��#��>�k��LB�oB��L��P�0`�PYgS�����i����{za���A������ui|�gwJ�M����\01?aj�IĜ{q��@[PF�Xrƨё�濻�8ڱ��i��[�7{\+�D�3�>����"Ec�-}�\�籶[�{�V���?X�	XlxVHYEB     400     1a0�Ě?���(����s$C������8d1�>pfOc[t|b���D��0)� 9zT5���[�`�����)�w��m�u��y��Z���H@�!�Ee����w�Bd�8Ө������.�<������P�69�@N�l�)�=���K��~�3J��i$���+'�L�����G�%�C�6��1�����%Kh��~VEk��b�]V�M�^�d��I��~�h7|���=�ښ;��Z�S�X�T�Q��tO��)/��)ֱ�d�=����F�)�t����dm�(�-P[΋/Ȳ`�۔_Y%K�a��)����J��{g�n$O ��<�H���&r4M0�6"�0��Y��)'h̊��ٓk�@�>Ň�ힿ-�NW��~n�R�>���ʝA�'k$�XlxVHYEB     400     150rc%�eƷߨt���L�~{oy�Mb�Xja�Bnyw+P���;3  0��n��dC�&�^R��n�����?`��<���q�� �0D�ee�������t���Fr�8�gώ�7>է�3D����u�(��G ��9YJ	p���>�;�}ٓ�h�l=����p�	�,�_�>V{�bK���l��� ����F虾X%���~K���Y��������n0>�`K}8F���byQ�S�+�2cmX���q��fƠ!�ۘ� >������J�]���i��;�z��p�\V��$'��a�a2�i����R��Q�,���?��D�XlxVHYEB     400      e0|ڧ��5]}Deޱ�U�P]Mi��R!p�Y�*m,��g/[F����#�8���Ъ�JĐ�T�آǆ ,������;4�U|�R�ᢀ�n.��"u�������{#�K�<�n��$vL�R�u�؞.[)`TW���|�QO� k��6��_�X�R<t�1_~�\'�*�.�rM<��;��6�q/�a(� ���l�iI+L����h]���5�B>XlxVHYEB     400      e0�FjL��B��9�kz)ً��&���������� �w���T�`()P�j���������hE/�=�{v+@|��'c!�*پ�UL�v���s��{����T�0��O_D���(�����B� ���B7��Rݘ��>����>oZ܋�R�_B�]�b��7YQ�3� Z�syh��ꙧl��w���H{��8����ʠ���i��G��QvB1K��&<�=��r�GXlxVHYEB     400      f0�W�6a���/��r�a�؀�к��l$^��r����F[��ݚ��6�J�	,3��q���j�;B{+
��k��p�W��J����2 ����\g�oO'��-0�R�-hpam~��	��(z-Hg��ˢ�w�/Rd���eF�A�R��܄9�}�~Uh�8S��=ݻ��N����_#7QUu��i���W�K���D�D��Ɉ��7��\}|c7�p�]�,�Ch��4C�Ƈ��.u��XlxVHYEB     400      f0��6���ѩ*�84��E�;�U�ێ�����5���ܫ���\�C.��<�|���l�]\2��&�����ݐW:.�;!����G�EE�^���%&�% ��1ae���C������0bt^��]�#�G�s^10�]�i�-�nsf�첛
'�"i2"2������C��/t�&�贀]�xp�!p�,����USL�r"�<�p�|]���I���ѝfq�D��A5�Hh��XlxVHYEB     400     110|Y�^�|Q[��Q�_�]������u��v	�4��s�r�o���e|��V�M��w�)^�1ģ���9���Ǜ�9@���;oX� �n�}1�����/�鰃�O��˫q}h��1�4��b~��7�:ĸPtr��ٓb�p �i����^_a���� ��R�@����w7Mp���7:)���c�n�O�0Fz��7^М?�!�αf�IfS3��.��}�l�&�*��k��Y�!��[%�#gL�j��)����� P�zp�u2o�XlxVHYEB     400     1b0<��2��&�r�KQ�R���'h���ͽt�N}���bE+�����7�4��CI�'��z���ᒽN�Q���QPzy/�m��(�����8���OD>��%�:ѼAB���JI2	?���΍` �����mXu�Īq�
�K�~XX�I]a���Wյ���,�ҋv��fA�	
��t~`��+1�dZ�w2~�f˳C�RuRb>��VI:z������ߧ��y�t-����<+��� �ڴbM��� -p��_.�s荭Ի��2���?J5�a�(M	
��1lFh�(f�ii/��I�x�q�NoUs/jL,E�X3�	���
��W��'_����Rڋ���s�`�Q�)A[w4Y��6�W�-�흮-ۥ>F��/�l�hE��Ӏ0Dә�"3�<b<�߹��y$�C7A�.�x��gH�XlxVHYEB     400     140̰��gf6���.jV���%Bˌ���Y��Tw�!%�X^q������E�]�����ho(+Uy�e�o���-�Z��Z���̠ �������zǔ�Ё�����)%>K�iV��B��6Ŭ��n��Ol�na��bg#��u�m��C�d��Qz�m��4o��\�!�m��i���Z�G﹛�.xs��	��A.e�J[��rɏ�74=JnK4�h���JZ����\��yU���?Z�Bb{G0c�H�}]B0�e>*��=����P	ו�T�[~��y
�ɮ�C�˗_T����h,��ͱq�S��.[��k�<XlxVHYEB     400     160n��pj��:���iJ��.]��fi
����=��K�^����IJ��0�6K������2�>?`TxLh۪�
x\YkM�v%^�=��� ����z��o��K�|ae�]��}H�&^�fΕ�F���1�n"����b��G����X�Mra�qCm,X�\s�gӖ#�Z���S�����>���o�p��X���F;��O�Z���nAA�����LRƈu�O$/�j��2p_�c��B:1�M��N֖H�t��{�X�v�D��)���e3`�Ѿ�7���i� &���e��6�.g�S��N2�7�6�߬��~��!rض��l@�WB��Ȝ�cXlxVHYEB     400     140��r0h%¿�7�)����쐡�^�1�]&�)9�2a��E�c��zR�U�;����9ۼ+�VN�?8}zUR��D���� �?��j�C���b���r��c$>\��Z� .$h�v:�ɪؚ�ެ&�{~�8��N�p@��Kuix:9i{����	��b<M~p���h�)3�Ba���v��$
QqB>��6^[29/��wO��>�`?c"v��r]m������W	�@c�5�i��r/=Dᥝ���9�SM��J��@'w��t#2p��/��v��$�%�毗ϥ��!����o@��[Ŝ>���fA5�XlxVHYEB     400     180���]A���wkH\�#%wF\ҭ�CI�
qΙFC�m�4�O�C���ZK�O�/�2Y�3��S���H)��L�\:���s�� &���aͧ��̓�B�<�&�_u�h�fت
��iZ�\�7�{����'#+R�[	ÛP@^�U�H�+�v/FC �8�'��2�.kjWs..�t�߁����o�H� -Gs�S»�A̴�������J�\��N�T���Y	 Y� ��7����c�J˕(�:"V�B�{>��p�o��9<�.u��/�q(2��KwF��_)�H�:�ʿ�[�y���_\z��h�S^��`F&ݨ�#�VM,=;N���"ʒ�G�^�����ͭ'�Z\/����X6��j�9����P���XlxVHYEB     400     190hp{��V�7��2�h҉u�Qmo>{��F����fȜ{ �����r�}8� I��O��TA'����{�I)�V��X)b�?���'����ܑV;������-�����<n�
.��Z���=^�}�-��u��`�5fj�r��LUX���+X��^����!��n����$Z���=)�c˘���
��q[kuAD�������oR��g#�ר�ݙޝ�����o����l��ᔾ+]�A-<���x��0��7hL]������\(����i3����5��I��a@�"@-N�mn�쨔��ˌ�g����Ŋ��Tl�|#V��5LL����,Cu7ܘ�<��	�U�������������y�Ɛ%#�Z��*-Nܮ׶�*PFXlxVHYEB     400     150u�H�Ù��Y����1 s�/�R���v�.��{H�$��@\
�H�FW��܈M�h�h�ŭ6+2s�J�l�{ӓC3�;��Lҗ�F�}/C�� _�BVǢ�1dEԥ^��ު�N�jKL+�)'�Jy/�]�LA���d��:�=K�E�Z����C1��Z�����v��(t���L~SUy����$�����(e~�����I�A���&���g�~�=�nC���I�<�y�P�)���^�˻Ҟ�	��8�#҆�d���\�IMW���GC}��.����3꘸���Z�}�:��	]eDE�����ѦL��"<|Av�Ԟ�����d�Y�D���O׻XlxVHYEB     400     1a0>oe�O��9��G� ]F��(P6���������R-�$�C� �����|M�þ�%�\?nmm�k�3�4��k4ͤ)�'�<�2����M�姯��3�vr��$!��ؼ�Uh�����0j`�����b�]��[|�
��{�d��
�}�ƫ�,�?Yo���#���T�)?��n3� W����̲�*a���J{�v�_F��M=P�R�QI��$� Upl�B�ޘ�PpK&��o������k�u���<�	7n��g��t����ϫ�.�h�xz�e�IOZ�V`p��be�\acwXj���f� `BT�V�u���AՖ�H`����K)��r&;Λ��*�p;�LQ%T�Z71�i�@�?��vQ����	�[��־��;XlxVHYEB     400      f0����-[躜@S�B\U9C��!���(.g]�vHď�b=�Λoc�|1\��\�J7YX�=�plm&��!R���Y'"���t ���s��ČX9�G��˼�����	��t�C-�=k �}Z��Sб$��_��r��Q]�N�KaJ�j~�(9�����o������^+	f�+Hv�W�1J=^ 1O�EqB�y�1����� �t���e�_A�T��{1*|j��xP�C����t_��k�XlxVHYEB     400     100<�����-��@>K�tϧi�|�H�|�^㨾�жD$�qM#Df7 ��O�#���..�D�h)��6��M#dMo�v҅�s� siQ��ߞu�BƮ�v�n�&H���3��X[8���� �69��t,!�����*�_��� #�V;��� ��lxsޮ_� Eʒ�;�����j2�K�F 1�r���dw�!s��48^.Q�S�w�8xa�ϼ�c�幨�{|��Wu��A�������}B
@�`���XlxVHYEB     400      f0<�=�˯�Y~��?
�j0;���bCZ�^��*�ȇT���j3kt噊#��鹝G[��|�������߲�t��k3H����v�"y*�w`y�l�<%F际O����uL�Z�d���6�F��객TR�R�3�S}��&��'�9���E��Ԉ�[�4�IM:�6����������n:}�n�~O�'��"W�r���*/�{�cW����&��F��꤆�e����0
sXlxVHYEB     400     120:-��ֹ�{�$�?�]Iҟ��z'�Ud�m����D&(!�_��1Q�8q�6���N�N��*�VZ)�T�0�%`���ڳ��6 i��P�Z�� �F~�.1��{�0�ٍ:�y�Ը�q�E�Hҫ�zcG����u\�����+��iVN��(w>ޅ��	��p!�ZYT����}�����[�<�-�o�TÐ넦�m����'��/����� ��������?h�7��b/��vsY�N�N���`�&��!����1�v�DOZ'Ę����}�'�\XlxVHYEB     400      c01%�vo��,������I��i�r�_�gޒ0P�KmI�3�mB��"�y5wۋ�{�;*YӶ���l� �N@GC6@��7�R6�U2�z�c�3�+�_q�n}F4[�|1��Mu�W�^���(�A�R�����,�"Z���n�Q�|y�ڣ9k�F��5�[P�N*ܠ!*t�ں��^�K��=��XlxVHYEB     400     150\L�FϚl��������l�x�0�'��z��������@�9ǎ����k���l�!��9=�N&W�1��:#�Ӈa��*���уl\
uC1\>�:�Ԙ@���+,��F5�@���K����UE"1��;ǘ�d�Cі�Ǧd]�}����%�O�.�I��N�p�?�}l�,	mi�<�ÕR��F��$�W�i_=����B��4���BhA��s�AZ�
9��Y^�93!�^D~�t�P�u9�������gq��VM�
�4/ �fr�uq�|UXiJ�U�
<F�Q�����9�y�ׄY����?%��^��
� �K�*]���Rxv�k�pXlxVHYEB     400     130���)�uq���FƇD�.�ϋop�Fp���ь��
��H�.	�S#��}#��D�ϱ(f����_"����p�ق�.�=̹���+��=wyLt9g� 0a.�i��Z:�6C��]w��{��S���4�UX�� |��N�Y����3�SK8������?е y�[��=5S�cR'n����n}C߀IS��v�9�#���	�瓍�=aB_�1�MK5��]�w*�e����"�б~��(��d,WeA���)��0�U�����������E%�J�P�z���S$8����lE��XlxVHYEB     353     160@�WB���1i�G��@(�V���6<�d��EYBS�O�y�|�G"���M�(��*�g@5��x� �r;�!��D����!{�?���!A'w%�������'�Ħ�Å���r0I��2��^��{ќ��}r��C8J���� <U��k��� �5&�)=���bt/r;�Q;α�
��z��T҇EtM.d-�<���=����~�Bmz��k'�w����I�HҔ��i@�A�y��½p�,����ew(�L������u�/�E�:���?�nXY祯݋��$�Q���r��r2V9k�F�2c*�����/W���/w������(~�n0�A��4"�쒃P�