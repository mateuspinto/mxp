`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9152)
`protect data_block
dfFNtpuI8NmyHa5RCJYNsAZfgdneduGvl53PXXyUeW5AeDP/9QHxjX33PfG3wJ4/pLrdpxzqVsjH
MuA8YfdkR4WLLF8JEJq4xqvnpspKvJa2R0oKA3A26w3qL/JpV617CTiuFi3ZbUBvCZstVwGKbQeh
CzxmVZ1iBURQeEJmUSePMV2RZbKHZy+N3AzAptPflPmys1/KMyijwAxVmMyxmL907E74qtFdsg9S
oOf9XgW779KQyCROyysnRR5t8Gkv3yjhB7Cs0rGoY5HcqF+uPamCSjNDJFt/LvizuW7ztZ/OoMd+
+FBg5JUEKnLgTvXfTSV++/2BZn0v9koDeCdXyK0TYbGcpIgfXlSteDIUNcQg4oHzANAxQcy+j4XR
BxNF2W/98j0W8sRvjlI0rycfnuuwpGE76+eS9po97taNMspZ2LP3e1X6PVAxeZcYlJyrHlRY1A+C
T2GCpzJWpTnwIF6weW0AyExWLQSkK7G5WkOJ2FWrelnMXm0bACrbmcaKrNTo/H1pvbzs/XoFl12V
MUWzVq4qAu/VlIWBg9R69xharmraT2ii3ST6Mf83QjA2x1OCmfH5n/R1BbFViDc4P72W5tGtxbEn
DkFBOpaictBESYXUC8zWhaila6r53uTh12un7pTwortL7TNu/FiP3GVbZ9sSrK5VCLvjsZuasQAW
DCmkuFwG7GxpZWflluvmHy+vZhCbyhoSfcWtSDDiit2sf3EaW/jmoM7fTyre0LQ9iIUQAyLS3uDd
ny/TMWATdAO6ZLAoqrFLkSpA/MxM5qDtvGLxeBTqn2bsmBIxemO79uzIFXeaOIKsHZ91pTsGbSYx
L8Q5BxNC0EAdWrKZImcyTIj3jL6Z+RLR4sRQraYExXuKUIi5cFw3DMYA2lUQOvQHyM6hABSwPLfK
FX5tXwp+e02/vKYurPvcb8Y2r4lbAx5k5SH5/Rh/QV9HTeE2YWpWWvHrAxx+HEs0Ef8PuBRrQm1g
QAbdySoFOGy/arlJCihaPQj83Iuvmkue0M0vLJR+boTeKWzKqFl75yGVo8cspMYiukzP9Y85yqif
k0fTSjib8QAcBMuvFaOSgBGxIrBg0XjpBjIjnwfrFl+rwK6gn/pFJkNLneMDFhVcfPq03eefWqFv
Nu40qhmgY4oT70jIZaLSksyXugjcmvcSLcEntvo8xRBnNLAKpu/DI528m6S6eYzOKO1dQ2y1DaR7
ukPIqineUwVuYMfnIH3VH70EC7cKMLb7uPrE7IPrsZPsCVth9P97sRBSyz0+fn/L3hQwlqGsapqC
hW+igE6ZtOa6+5yhM9Bl+J6KwUeRFPrn60MzNzl9jH+XM03plWcGHvvv2d6ZECBlzaLo6LFazItd
yxKzwHOBDDJtIxANKJSaAqxhQEf1kUgJtbvxPQOcOG+GTsSMY0Ir3RjiBhQBit1msir0gJXgP/1g
Q58MRvtPmhN7wdn4snIHQsVDFkP4bT1ROHpyhU0yom4f/ggT6e2IEyGFDT26k5w8RNANqwddikfg
Hxv30LowWpZ6TlJ/lrXTzMf/l2YpIsvG1couJIbN6rkrbDTxLOPd3UYWX7ykWSvvouWL2YBmFNTI
4geU60O9FqPV98scFVE4f5xwa9oxLA1iAcoimLsE+DRccffsfNKVIJoAKktPFkN9VmHeZCoUs02U
ULk7itA+pP3k8MyfwiMz4ShSwlnSCTfb8n9pFoD7evEIPMaWXMeHAhU6zKAmBI4+19zswGYiNlH4
rmN2//O8QP7q1Bwi3owV2JasYAkM0uBurV1NlMh0TNT17CDQPHP1mQCWpbMCvSN7XNNhdcGpKueH
PD6mifB6ITE67PdRDKUlxqkB1dtv4Vyppc/37LnBOlbBYd/3CHOsk6omRmuVBmPmiZMtrbG12uqf
uhduALHfJDOw+5y1m+sI1LmRitqd8r2B9o6qGhA1+zZiJtiq/zYwhyh90kjem6uDIcUsLmOQYJ7W
xQV86psPXCWCoxqldE1UMi8Rb6rvkWwhfk0OwS5yQ+GCIIABVtbd0J3a5crGXbCHVWWfVufDqu3W
+L8MDKg9iP9WQCpuVr3TXDV1+iJwWm7Siw9vvlVgOl2T1jpdNy2oYrMnZPc0uLDsWrApK8vTcqoU
Hm9XcfVEfkdMCc45oVZrwaUBK//Ra+ZtMneqwxeZXmAkfPjq0mHYj6HP8d6JIu3YrdgDJbVAImsG
5OrQSYTNWx5NKtOn6S2ZB35TV6mIGqLrauv3evHrAcfUkO526eZAbEen9HgDqk+1t3dUI5iV4kOk
dgniou/H/Lh5qFgohfduxKKjgnGZgOMcOvIEclFGAZUFOUu4ZvoLerFXvZpd784qDCiPntPKPdXu
sHjxazYedU2r9lXMXTsbiSTOgEWrT8+pSYr9s5/DTmskVvo7WdXuaNt65E0Gn1HZyV4whyTOX4I/
tk66xpNwocYRSWGihtr36NqR+Nec4bq1lFJuzsB1YQdXeDqSfeUM9Avg1IPB6EbU6cuOLZ3A85KA
f3ZjF+wcPSlAsPVXW1o11qCdXCTTTdqpLMpWlnFcrnre/klqmW3Rj5kCxynVC5UurquRy7axPyeN
fFU95WlVkVHHujacVBh0231yZUPbWQbfPfT6aYA0YkdgMvhGzbUmSbZfzqscAJFVZJG6mi2HpL3O
Z75gEvoh0Uxi9bysNqJeAD1v0nkuw19sG0DhahM2cdqymWJfDpF0bmKvYOKLvw5o/t4SEIUPV+gK
uSa/MS4H9D+ZWAw2swJzlq1m/TY6mn3Lg2VgmF1Cjzq47l9RaScICcMZoUpjPFMixrln+EkFg/ip
xoKcBLp3K+BhoQFiwMY8IAHKNOTAklbma+cxfHtCPYBWLdWfbDioeetX4gaf/UFzIQzS2J/y6W60
2nV2H432b1puoo9pu7ZeJ4Y2UGqUf6DshsUveQmL6f+QgQCKRQEtHFgAeOxFSQLizcdcXXXjGU0H
vVq3ODJClsAUHZP0w/UYUcR+7xoTovg6elNcGfcrGQ0kCSyYT1xm9mBfloL9YzAIWKic4dxlcnG2
PMISegRYIOPliyphdiwuCmf+5v1gj1WvXxhZlUNg5Ccoh0m3TEJp+RBHNC/ktEquko6rtH6K4Ir/
kc8VeVhf58Yk9T67XGkn1YZj5EfWZFFkPR/ZeuyxdN3g3RdqvVeQSrD/5zpK7u6C6gxLKOq/DcW8
g2dv18/BGkAXBsKbbHmSbTmojPqUd52XcguFwsa6U0bu4VMMJemAZexT9zPSFe323RH7Xd47jPFi
w+H9GgkXoNi5tWgLxH8ETvK5edLvoKk7LE3bXNJ1X/Ook9JPea+UFcRD6sD+IObuwiT1j52lRABu
Wskp2z39KKTQn/CQzg6E6b7uC6AX/ESdp17xNEfAj2Kqajk/2sthJQeVdw7zAFtlqQvUQVrKkPP5
02HVj5oB1jcDNyfcecijL1aarfpIG8eLNWiM+FK6KTALW3HjVQggVbm5AJQsSc7Q0RPdxhjWOwsm
zIIIeIPyPe/8WsoWG8jdTzOheBKsdTJVBbbbj350nl2odw/OTQ5Z/ksAsKBedrcRuZ5MXXlfemXk
a8aL6QiOu0FfQ1qFYdEGp1nKjYNKLGOxuq/4Am1ckrp9iuxLZkFTMjeX9RI5h1f7GY9qqgmM5Ugx
Hj4g6Yz5LrpEsEW04YS44/p46JHRGih8+iQ2UV2OB8+mAEWKyalFjrG/dsdK7iyJPW6blnWf68P2
avJPwB/RS4SYOqmM9QF8WsabO/e6EuBr/RnFIXG9ZDtnC8IZ/beHRr575Pyx/1FmLGYLw3VyYeKS
/tw5rKalC824c6X8mxozX968+7cuJ8Cq5K5Qru5/p4Ih2Vcfa3j5pfFRa0DrC8hpuCEuPcVFxgza
MQtp622RxL7qf2bJSs/JZOvz3Xn+EXhWARIQNo9H49pXPci1gY5ssWQGP/wdwNvtfVknlhQTyhhu
ZgJef6uBXRniEeup/uDFulAl89FooojNhJLSRDwLus84suStekawm6NYyPGfVbXmvMdOcdt3Vpk/
CtlvCZPVq1ZwNgq8CUjvSuygLEQj6kw+mKyXpHLk+IieTwAkE78rIc1bR4O62/HfZGPjCBXXVTVK
/a5GRXY+L7QDhUcrr7MRsMpFCKVCx53pIEh8e8PGJSdnFgvvevxPxp2KJr+0CdzSCarqDRBLwBzI
1cA6epOgWRGoAEBBGccg9R/+wHASx4gFzxjvgHB9VPewcggGfX4h4sKBjw/oPUjDkwHREQPp30mg
z4caPOq9XUHUi2TjKPPiNiDPv/OUNs2BIBdyVis43zoh/S8apyHSi6GVJ0RwUbF3CqQ8XIM8i1db
A8yPh+UKXXLyfKMqQIEsq1sIv9Vt9+r+AVAnQ2semsQGttqcjLmF1PPJuxp3++z/yabxFIpLPXEz
KGok4WWLmTCfE8Jxz4bG4/OxsNWwzZxFbXr2cO3jwScc6AhLyTgKaQoOxekeXzWzUvRgLuako7TE
7nuhRpeSgp3yRlslsVAtwLMM9tpyGkylpB8j+j8sHdulR3GU702oV8tE2TnzIp9V9UofCmcJwSYW
Qd0iiRaiw1pW9EBrCK3WK663Ql8eG0UulK2ImgReBMQqBXNHqK5rKEjkIkbem86R8EyJbsy41ipq
B9Lm6FiYX2BJzmh6p1lHSMx0WkANoMG1Ygg1xlU4gvZNidkFoV+d/21sAAOYnRucqYAxmkmBDQUR
HQyfRYVr0Mn+rLRe6CwsZ9wSnspDRXasMUd/sZEQZ7BLdAMgqjtZwLM9B76EmW/d7plpH/f0qs68
am0ITsc+YRXtFaEyFPXuGul/tn46CHjlxD8tONPTEDoyB4XCGnxv3JQcwJE72X+J1V017hDtON/g
AtYgHO0seP8Smlk0lxsj3YlL6GmEps6UzuEY68JieCTaacu40l6yaxEXFSC58RQce8lgPEiSDL8k
bprvSzEwpYTI+WNGNAY0CtXCVW5A22Y8ZnPUqIoOkx5N1MPosnPhegv2Nt4ytmmkOZnHbCVzvFUs
XRo1n8sso6StoEOUEmHRcowcXR8/jidwPSBqQcn3ZJshyq472IacRdwLLRFIpcEddOtbboy1TtlD
orPA4i+Ek1y6C6vKgWLMuXC6SRUqkH/gZF23/18fDYt4fP3yKGC0v7Kc9ZHsmZ1617AzQRlCsmv5
+DKVHAeuZaRRt22UVdkgLwJ1WfPnzOovYoGiMlLJ3pOhx72oxcWVVY/EAGZw2XiykZVlpbu7EMhA
8FLpTNjalmC8TvFIEfrDFA+lqkwxZknSntiaaXO3VNN9q2XGc50tIxQOYkhNkiLP7jxBPmJLS48S
1UKQKLnO9b86PZBzD4CbZRozNi0p0HwtqfjTdxHDURi6YVCkMB5+Zlh2QMQKNPm/o0wUKtfxSV6l
lJlh2E9iENSWHAGikKo0gQhMqSttvGr+nuVdVqCeTpmjD6LuJaDyBSHqTdbgciSbSOEbvA1wJiwy
VQqM6EwnUNkYMBmm5QcQ8XGvEo7zv2c7WcJm+mQfo38z8GgnJKwz5uzbA3YuGMrRy7nLNqhu/HMK
LcqYDg1UIAD7TLA8b1WrM3DMMp7lL2mmruzoqqFEARWYEXidEuVI5b09dFT26zYB6F5NuGTUpydZ
6d068KpBmg/+HsJKVMpKn9DEXYORs31VdK3lWijyIRP5XkFGeIAjJ+PrZVDe5zGzS21EQH+Jrcwn
cQQxgNX29cpYPYtngfLTt5BMja3s87B+HLPpQodIyuIwgcS5U/D7PSvGPNn/xrZcAGPoupjR45SK
Zp+g3YrDuHcph+Z13tvRE0ABIheBdwfP4lomz2r3oH+d840RlpkddjxcrYHOWZay/gfhW0ZBZ3nW
2UYPnYhM6Lxz8w1zsnTcqNT7VE/5++KfGd0228I1Ql38kHuYqlPODMVR/K2G92gVEU3/tHekCmQY
EEL1l/5Z4SklnjNk8l9guMOj+GzJXhdIufZWZh5F5ATNEtJ8LN7SRz54s0SMfP3GjkRlQfKP1bRw
w9GWHWpeRN/RqUazvN2ru6Rv8v4vGZiPzyzWa8qyuqQUKyYvCEp211Uvjnw6KxDylqC8+dO1J9L6
IYE/XOLSNqz04YBb9Qn3r3r5PSZzaA8UkY9whgiWs7VJ66423Q8L3/qVdVd+EzHzfwK7JcnAAEW0
wjkhuMm9PES94NLEVqjH/eHB1zWCIV6oWGj4yB9wH0bBJJEolLBpFG7wck1dH6GBHSv8mWPM+M7+
acZEeBtELx32Yb08YZtepgC6DzoppSeo08n+UIoOFdjrLOQcdO/6txPeUyWQaq0OgiwkAqfi7jXX
Xv6BzdMqEMC9d3u5pu9rm+QE99RCSXWgrUtHR0HRabm6kTH6iU1kzrB/2qEqmB7hpzc56Lovs8as
/raMUV4Xrp1n26gLJQj4M1qgmih0jmRZLBQt3lYrl7LGHavtMg0F9nT+rB/o2RHkQ1/LrqMSLbXV
HOD1gayfAYjIFzJgk9gzdQR5D/ADfOydCkaim4K8Z9L+iOm7o3fQUn50Xkz0ZxGt9jCOEcbp/nsJ
SsCzsrtJ3ZJFV0it0MxM7IOHkrtv8w4I5fmEfDhAhVux8tZ6If4yYRGAcwOU/o13zpWyESepLKST
HiddCPlyzNaJp3eELkcn42xjYFuElhyZGg78ML2jS5vtfKR4MUl2RIlCLstmiuOGeA8mr8zT2JZu
r9oMLCjHHmZGZY2KTjXrfR5jmKrGX8zhuptZILHIvBnPZ5nwyItm19xdKNgPHpHRiINe3rLJt0AI
104pl9e3LBT8pZmuOsnrmmkEmvYqukM0GSTs7kZyyneL3s50zHlmpa8MyopOX7y7oGKdQp5ZpgHm
MT9kjU+5KDrLdH05BM3lGdnH/UaP0B7K6byhPJZe5sg4ifuPyQE+r+FualMAAzsuJA1IXuvpavCQ
UdYCrxlLoq8ivUR3AQJYejzYCAdmntopPwLPKCIHzedvBI+6mPLvnzSaf8y5WvGVkU4poxh8fQlq
KsmFi33JutUtCgAjuizD5f7Yt+eTyxwZ9Vc0EUmKkOyuaDcrFP4ZnHDF3wuTbT1wkiCnftiLnH1k
xayJpc1CVP7r8x9dLtkvLAPdw5iDC1Q9cF1hFDixcQfETO915vIg9++jM+ynnOBeUIn7TYIdT6cW
qEEp9f4dR/pLOMuqXWQqy084UhmZfgYnseIX5yhHoJzPnb7eYzcd4gI5+l6kUa0mEGPNLS4A1MH/
cCp8AiUAFrPOd8BjQd8zt/S+6stidMUe1b1vm3oIeqLT+axJCUYYqfLHUnbmMeiMH3daNoRpGFx8
TFxnZLPVtfX8r5bkLVn5RbBk8OErwc70dCZNtAp6hE8m1wzqIKJnM9fojzw15Xz7JjVMf8HTfaFL
hzptZSXn95dCNm3tobbLxm8ycvPvEu6L7NvqrYAciIbuTXe85IDXi0jts8HW1hrCvjUEmX0hncvS
soSPcH7DwhBFWKuYhjW5Ty0a3Q8Wq7ebLfsavP25E/mc2SXjkaor4KmTbmWUMeKVQMUnnbp0i3J2
ou04SaHFOzQmGZES9Vgsywpfq1PtWKOAgdGM3AYOObNG8dp1JPexhJlZFNc1lU6lvEDBc8cyIfRG
kANECB/KpQlFlTFLohpO2TE7HlOSstWrlarYCDDmPwzkIAPmjy20hx1O+ywylIii1Ve2Nvlsxguj
bMuCvMF1g3kwadI0o8in9HHhSl3mG9gpHZ3HVUQ+mwii20cyQvs6oD2vItZy1hBFTBAZkqOS1c2C
hLNLioeG7Epaxh5jjXl9oTBH2AWcW3N/h5deQyptOM7eD9VwwKxZWq1ZU5FWVUYEF93eHEP8ceJr
ym0LUu0nmcU0fB8rr+Ybjac/uh54sdfXN2KprC2TpXkK8ZaKNjb+MXjPpuNvBux91CAkiLyoEzet
HDqwfrubVdQeYEsCJp0LU7jgh3cWNqyGGH24NIY2IPakBrePrlOaaRK8+UFDNjKpCphSpvBCUYn8
6hR3PJ3KDDMl34JGPNXdJkAyBkwvqUQrLnmWJBpEeni3IrnALEPspe89wdlJnXyTSnHCv599tJu+
qdp4gwBV2afrM1ZuMTeLONk0b7bdZQwkfyn94W9jyAopQYW2SiaZGyTT73VSO6tDvP72bdjmTnY2
7IUm2ikNQsqxsunVYvdV5hELldYtVcaZBYQB9f1DogzG5DDGbKjpZ64aQE/JuEGnGzmw/FJBqnNC
5q3wVD9OqKkP8RdRAat0cv7mfEXYxMiR8neTNB6+Sx9f7CC7yLA/gdnbh5kF/ErAQE9qf7Zwg05t
ZYhUIXMXpGtVs4A/6A4max1MIWRoK0GdOQ2aQtgsjTyMwm2c+NB0kodH6WZlSkmGwwm+EAkbT0Er
L0B2vkLAxgw8DWX4+uJBolDGcnTWSZDeei6IILdIV2Z+bK7cGUuALvItDIvuW01xQL0U7I81zzpF
71C+/BT7ybEe0F8e2SF7SioCtz7uj3G7MjHg0Q798uSKDD6OkB4MHXzkVyQigUx0Jez8g8Cgr7Ht
3zQIHYTy38h5hg1bLjzsMLX0D2RCJDyTHK+QNW8h2jQM8rWAkYY/hLXYVR8LSCqh3XL4Q8Xc+kdy
1zAOY5AYzJMJfsyJBQ6Qi64DSu5LVT8waEdSX4SbET9UDJr06/1S3JOND7Ffus3l+XMe6Pp8KNp0
cuZ3TZIOuDu+AARr3Y0rktIps7Nz96x+5/VkOwCNS0C7J9Qm5NzNnbaGVvqgf9ZzOascbXPt6qS5
lH8zq4ynsb5awpiViFwEdDmvm5fKaV9t6Enj8e91tPHFQGO1a8GlGA2od1RRVUpqEcEaJBzpNd0a
eHhYVZdfCrJB13p7oQ2zEbFyiJXptDRfdwaByuAQzU2J2n0uec26+D6QzaUrY1Jq6rHmWuFFPSnA
PlF+RfyOeN+6uOeTAUkUN6mnZN+EuYylYstrUEIG6gKeXeHOSlkgQeW5UcRr1r8ceV2LdzURlpiY
/yMH+SRMOqgiI44NeENvanEQ/ND2NL5tnwY+1xia7ukYZGMJYIMrmr5Cg5pHb7R3rmq/p0aRrxuV
/mGuwGrtonSTFU96iAWRflhH2yQ6avx8j8IO5gXenH5KPRq/tGtfuqtqj3d7OcsnzXG5BeB5cl2S
E7REv6WwGzV96L6TRE0zOlDbXdRL2mNhnrIUHMSJQJhrdmrsbcNTYBQKGcSWe3l0i/d+W41CBCwI
Tubo6QrT9wSi4GXXtO0XCFO6pjuaaGvoLP4bEzhosjUGSnswdAe7Lz3bdPZCsgxApf6tTzU018nc
pOmsvkjg5eUW57JH4kSSKXD73VNWTMOr5Q3pq2eLeLYsA9nRwgvn2msAE6jDRcTL9+LyyrkNdlRq
7crvfwMyLU3vYryxco6vk1cu4fyDHvCB0ziS7Mxs/gliEYUmCwpvuMNwXir10bFx5UwM51+b4kTy
4Y/6EoNpNPlu3RQnPaCgvChuEz4JmX6f6pJT8VkvSI07By2v0bJvNU+y29yzOqszv7dBgcnnVsJC
jnXKsm+9ntvoRwZJ2XN7EEnKOTgBIlU1+dzagG1GUdS07/8MfAFaRYrNkCrfXaMjm+6q0L9g93/d
gPg6c66icsj3sw56IVr7CY2yabfOEs8m/7DBgKnibQSrHtNdPX2JGGmOqmDrQmJdnThuSp2VX7C9
6NWgodTgcItv5EK5ivmfTrK9MfZwTt4JADUfWnKazx1b4jU8yEy0DehO79mdFg4juhnI2zdlewkU
bmogwRXOjHz64/2hQPUWefjiyXnqql0crEdmpNBUEpeMSvO7TpzsC9ayvH84sapc0foMML2nJ0I0
k77EsBh+ICLuFniaUMoo/7DOSa5j5JP8T0yE1znDtkbJ6ddekHFDUTW3LECWkZ8+xir2IzTFN96/
Itu1vnW1U4HruPU9AjmlIn9fRG6uqQYu6fp3XD54ujiJHQMQXBszHzKeff2Ud7267R0kK38P9kOk
3Jio03cZ9cUyrm0kSFFDAh9oX1rpMfr3eveXmbCz2KDNSboAv5sc6Uwkm/WF1ENhVznol4bjyACx
osp+ExUsFybcRTJnQSC/oDOdoudqePr06HwRVdOAJ5FYTShhZ2pqguHQove0wGEoaA8zF/7PTt/P
hJ/yB/ajsTazWXwBFXdtM2GxAZaqhPoB67dyQ6LwCKD1iWiOiHGARGK4zTUDt544suAaileKHA/x
ilmlAuyTgHbHllML9rkHywZQ3YQUOhB80RqJi74xTcpc8UxHBQ+MDBfBx4Sc01qG8t5VQYhZ+bjL
DmwFoguwOHtC3Zg4JsgrQ3dAPzLvVnf+kmcFr6qblMoUtjW2Z7I3QOiv4MJQJXaxN0YCkTF3W0vA
ft3lY+NSjgGdZ3BYxQ6XfwEnUdUVCd+v56iSdVTFXTfJ3RSwJZZ8jBYQgnPc/7VA3hkOWk62iHe0
Z33q1JYomSUTJZMxpggRTaRinT9hW+ucAc1O7Dgtg4g7pn6aTeQySA64u81vit8NKvYbNNOiki0j
oWBHeN6RG7FQiQThmAieepHfu4y3DMXp/Oncx5ut9fnVfdreO2vwZkR3VtxuwODs+vqy9FGGgocD
prN+zEtWGd3gjK+SNZVHoaXxGHvVgxeufCO9plwDC9Puv1cSKNUtzSRKBb6TDEwWiqRqoxVgOI+t
faghwyoGFV166eItwGEXvq+2xGHDdjrsUH2+W7cLYLXXIN4LRo3/0d6+uEIUIBuuqBwfMDd1JIX1
nDOgYslGWXIhgAEORse0VeT9Q1N30wpZ+MufBht7CwsgstEaNPImPyj8+OM/4axtXhIv9lcuBTPr
VA2gWxvQfTn7bH5BsPY3O2F4g8rac48ee/Viq0YcNagPqq6JXKTJUgojWFPmj+1svCYxMGC9O29a
6YX8nZ/eel3opsXXZUM3BiUshvQ5sKNZnly4Yko6M8JqA92qfTMTLWNurckInhAB9mygDW6gv3NY
YqtWgPqqO6qFkElE7KS69HT57nKjoxrc65FHCmq8DUD32R0TF5Ka6lHI9d6pbY8dzDQa3LYQ1fLu
S5aZCx9eKMUfgYaAK/eaCZ+LgRsGPLE5aeLoDucwbnVBAFpTmWxMFtTxTMNje84Cy0Sk+WOiz6KJ
Vc/R0e0l993wblngeUzZ+1M6Tjspznz9qpx7AjdE+8kkgk1w890DPKi+iDRYUwqoPAjI08mufP6+
wShQR4hQR7pagnTRA5Fi4lPupEXKzMTSGJqW/RbJjD6vHS8rrUakvrmm4b0Q6wVhM6gSfNz/5YaI
TXBkU3w7XVdwjiFAY40Lnp6Mq/ESDloDRN3k1fZ6fT4Ejg9IPmNvkGr4wZzsXfNYeDPvDq3AfN53
4SwfCcHecB7btUtmCYyoeodVg8WDFG/wzzkEsrhAqMlzX3xLLZ3+muaDXcbVmOszX/Pr/KHYiNAa
CIwCh7LFe3oRCfiJc2ijSKmCVwtEk/Ubdnw4o5nwRlLAlOwAsOw18y8PRmnKMOfzfT4D9gkUpNox
T+dQDlqww7hLYf0vlQo7eNfQj58FFw9VbBBKa34794ePUMryJDEzI3trnVUGeirSncwbOkIzqAHU
1Lk23PNDC3PgLxzsQ9ik/BUgv+qUzPw0fd7YYbGPUoeU2sOB8yrhuLHsTrUXEiTcoud47/2i3lDU
hPCo3jVn2ZNBnh3eEyKz9Sh1alMELYTNTSsj+bQhOvPPQ3U9aJ8FSRAnxizOjlRH+WssH5qUJYA8
6ZC0jEhXvkAkwJyfZmoD7dP7Y2EyxV3SpVjs6I66prva7vmczbUwTWkK0DCy83Q22DWxlhV0wXQ7
Rg5UvrJ9odaXgz012qk8eJM6bNT3xX7Szdj3VayVJvG779koI0mxBSU/QFEL34Zp0f8oQefu9YoJ
XaltDtnSEiMJB40a3sgfEsUtFlHsMlkmx+9f9wADuT0cBIp3CvqSzhjkSCca3SM3GnyV9a56fqGr
2mmNiqvtN7D0DSRs/G0d/E26TXmU2PZodF2iTV7KzqCimItQEc2OtDF7IVlLXzXfJm1xNb6UZvFY
fWribdlzKl/TF9WuEVKrTG98/bBDAJA7G6sEaJY2XbbFd5gFRoFoFLeO8r/2sx3cGqD2f75gkF3e
+tEcZO6OPiw1zlwQrziaGBo3rGwxG93z8rZs9xh+y99bkIEX8BmrkQTdjP/THWfIizCKro9HE82F
3mKvXDb4U8mv4NcpqCemgQoQpJT8f1nlTnQ+noVXY/0=
`protect end_protected
