��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���Z]�� �+J�?�ɲ~}��R��C��֢��=����7�(Y� �|̵�[�Ԕ����;t*�3��s܀��Q+��*��b�H`w�i�~1s�$)s��.o �#	�3�	��s����:�t�9�W;R�-{���[.��!�SK8�c9 �>�v�������$��pQ�w7�a`�������W$�f.����^7��Y��b%���Fq���-��.�SE�GQ~�a[DI����&b���(DD񗢤��t��F�� 3H�U�
�v烤k�=v�+J�Q!�"��Mj�o�L��b_th��&��"s�g��^�y���E���<�����%��Ȣ`�������U \"'�
����"aw��vZ��?=G��Ȝ��G�U�� 8�=>��|�D��4���%>2 �+��!�,�0�6�P�YX����l���s�)��;�>�c�'�<�`I�kE2��t��i��|���D��4G,4��
�|#���%��ڠ�bWjg�I����i���r6Q̄Q%2�S����2� 5���9Ve���7;�Yk��+����d����Z�����I�Xއ���m�6Sإ���Ȑ]��Ŧ�<35 m;�ߊ��/?�Ãv	y"݂���~������/��U���H\ԅ�U�+��~,_i���~Ԥ��C=��Ǿri��CP1��;�LS]�o�탛-Ox�����]#�⫔c"&>_v)3�U���A/�FV�>��/.{ֵ�q���R�Y�!9Nq�oT���&Y���V�աHn���h�$�yMf'��֝߫���6ϛv�o>xv��g��\����6Q^>|
{����7�H�[��eF��SțPj��&�z���oxA�@ Q�Jߖ�u8���<s�6���6`-F)/�^�(	�U	$bݔ�!$�o�y���6�F@6i0fCbT�tws^�{���|� �v��_*�M��7�:1822��%��xPB��[���U}-�8i ����U�q��ԎT<6���z6������>��#� ��Mf�>��-d&�1��\50�,l� 3?W�
%/v�0~?�N�k�ܚ5����k������ŏ��r�������E�|z��-c� P��7Ǵ(����@�R��P��5x��$qM��~���Ql�	aJ�Nh�&�ͅr��e��e!8��|`y�|w���k7j8d��_?k�הmn��xw/��W��e~
�LP��\��5u��H!�6	��ᕞ�š�����:�3��SD��	(��Od>�)��������P�~��6M��i�_�C���q���&��Cf�ҿK�I� ��,�h��-������ڠ>�̋�&�1>bڬ�Ƴ�������S��pOe�N U�P��Y��<����Hũ?V/�{sx��dx[`b��(�h�wi�wp'�B��=]<L�s<	����z�%�{(��(����F�=������t�n(gŹX�q�6{�(��0~�ǒ��e?3�o�ܤx�$5T`k��;#&�kS���
(�7D���F_ث|pϕA�N��})�/���G����a��i49S?4<w��t򮥛�І��| ���x�e��)�����Z�d��_E�v�7���8�L�b�<�HI�Źу�b��Խ��_By�Śs���/��u�mLl+�j �˱�r_��7��v��i1Fc,�{���vG�>���&d4 R7ͤ�Ɋ���)/~"p�r�������Z}3���sr�ar���8�)��ķ��Y�]/�Z_2��/�%ت�
{;�4�^OD�'R���ÒZ��`�xݗa_@Q��qG��l�5�i��Lѹ�ɿ6�#}:rIY(I���7��l{�X�C�ہ-
ig`ܴ`�hg��xR9�'L-�K��'�3F�H�R3�����O�z�|�)(��>�]�h'�bD锆g~�R�fo=�m�j��(X=��N@І�L��a@bl�)g�4�2cl�NQ�[���Cش��=M#-�hS�.�G���~��<�Ti��FI�N[X�r�ާ�����K�m�A�����t���Rxh|��R�!�n"����� �x|8�Pt��< �&�`��sc�N��H��`�y�Z�HHGݳ]�8_G�+���8�@��v-�(�+�i�?��Ē���q��"k�ȌC}���� ���X��9�A��l^���g�N*�����e��wz��k��d��`L|�l֫hh����8n;�vT��K]�x%�Vu��R�p�4Ǳ;@�u+-2���K*�d�v�qq=�Ws����kD�P$-[���M�oE�cb��/����M�m�e�"N~�T�.��#qn�|Z�m���*/�z%��}��TQ/k�v�A�;��W�)d�To�jښb	#���)��'��І��\�{���`�=�����:Pst�xo ������h'�9�[��N�>B4�-X�M�O�%R^��2���h��艹t��O�н֓2ߧ4��80S��.�|7���'i��b�>2�Al${萁�v_]:E_�2�8p�K�������+S����F���F�V�M 5�
�nsc�H��~D&�q7d����P�_}�'���v$;��	6�$W�����ēT�<��˃�B�>�*B��,|M�K���v_��%s�����u��^
+���f}���v&��33���?��:��=;���V��I�'�>�>7�װ��z 7/���-���9T� 4�A1�5|j����,\̆��#�vFJ�S�'+ןl65�Yq�ל�+(J��ƍ�������!�R
��v�
��I�B~x���<9?�!�!�9��M]q�/}��D�"��T�Yf!�g~)��&��t�yȗ�K�%���&�/�&�3�gT&p�q:�ʹ����Kud�N�L�US�3D����X��ST�.ڞ�@z��sp�V����w��Ԑ�BK�))���,?0���5ͅ aW �${�3O/$�M��n�r�5[i�V�u�2����w�~��E9/��'�_�̲�D�,��q<��V��*�-��|�ό��p�c�d_j�1��h�%U��\f��)����(c���������r��@bw�?���h��]��|Yp�<?����p�/{���=�Ko���
Ui�a�ǈ3��R�%v�^1iC4����]��ZmK(��h�<q�&�l�o�S��&n5��Z'�~f#K�qL�5���Q���>h(��H\̃W9�-j�y:BG	g+���Ꙩ��S�3��% �z^鷦�cO�ջ�'n�|�b�x" ��H��1�u����O