XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��T�8Z�J)Ԑ6n�$��N4�OI�Kcw��|�����"1M�e�T��C$u�{>{F��y�������a9qvß��˜�T�V��<jJhstK��a�䵺D��`^��1����g��.5��G,0�+��eq����^#N&�J����"Q�K�V0��2�<�HqT��V�M8j~1��~�Úga�>@�E�F�FX��VN�E�4�y=��}�`������R��^�����x�f;�;�f,7fQLAd:V�����yݝ����Vo�с�Q�OBvHf��-LO���J]5WC��0���+t�����e��Ht�%�7�B9|N�M��N&�z�-:�?	�:M���S�i�hWJ����~�S�܏��2�@�U���"f�1���f}�~Ͼ�����<?S���r�0@Q:�wn>{��vfP��F�{��/w�M��Џ!Ru�Hf��������B���Oe��<ϒ�?��"��4z���u��_�ܹC���*�C���1eU�������B�Rm�_F�j��5D��
�<s���rF�7�ۀ�Pi�Č)��\��&�(5�4Y������p��#r�:ڥ_ͮ�K����
�D�n��؛�&m�V���c��Ȅ�CW�-ՄWK�Q�lON�-XRP�����I���2(��L��,��[~�5.jg�����c�£J���5�ݸ/��E8����t���MF�5���k��s��윙73��3��@�	�=���w������XlxVHYEB     400     1d0/0���s�xM1��gj�M���v�Kq��\k֐|kH�U�����59�4KS��v)���
�R*������+(���<nk�Vj�L�����>�sR�%7����M�Ζ�L�{�tβ�-�QWo�~���R�0�7��/N�����	�U:/X��"ˣ):�Ř��4;��M2�2�c�^���Ja��UM�ot�F����f
9���&�����J�э]t��ρ��-��K��/6�*�<1V�xmB�K���{u�R5�*�W1=׸0«K�5�u� �,���f���g6�o�QS�6��"\�r��]���3�·�iC�<#�Ij�⺥�����9��|z�d��؍,̩7��#�Hm	\%š:	�Ђ�$�x��]r��@�ZY�4v��v@ѣU<��I��z)q �,��~�>{Nk�yk�\�	p�kB���e��Z�q�VbNXlxVHYEB     400     130p��
�)*3=��/�ir���]Qߏݑ@�0Ej^�A��dr쪟5���'Ŏ�X�D5z}���_����Gm]@|��~�*u�����)9����cj��"�@����� @y�#xk�T0=OT�b�1�FnV���B��㼲�@b�&�38b]�xc���i���p��B�v}�UVZl�zϯq�������/T�`��� �^�;�δ9W9.��p����P����b�b����/�
7D�ku�j�C�p,>��o׭ �F5�m�}�k�ۥ�j(�8�7�X.���ߖ�B�aXlxVHYEB     121      901���P��.�U�O��H-�=��k��g�m?����Kd+�-k�#��a��"L���$Jnm⊛���P�c�s���X�\`�[�ȷ� 3�E���7�e��̻N��������9��$d�E;��0o�^R��p���ѹO�_�ͽ