��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���x���h�v����Sh�-��E��ϕ�..͖Rh��_�����$�H�����#ڝ>�[5\WL%�no�a��/k�}��@��L�,(,���Z�c��3�!;�~�����\EŏL�	T '�?�	$ԷX#1B��`���Y����ݍ��
r�� [v��_�г�)ߛ���'���_�jȡK�b*���z&�l�#�Ð�M�g	*�������b��W?ݪ�ZK�J��WfaҸ*��t��|ʵ�Bm"�QU��vB�Ԛ%�z'�Z�'������^�}g*OzctdK�O�s�r�F��~3�Ј?"ʑ�,8B�C���M�i�7D�M��������t���@��MҖC�7k��X�tv�7PriS�r�z�u���g!���2
��^.� ���0zcF�����!K{�Fβ���͠xu��^��b7LB�aY�X���.�o��yy�^C+�v�����%rg��)����{"鱗�툙}9�j.,�Ly_�������q�&���hۤ,R�`G��@)o�9'�������^���m���?V�c�[>�դ�6�L�(ØN��\����۱z�x1M[� ~�x��=o����
��V!�Jp�-0͌��M��K�*8{�R�ML\l��T0!r3wz��JK��� ���*O��H�(�_��+.9O���X���(������s��?'�Y^�OR�:�ܶ�Z̄�E�5b�*w�Y] dNKO]�*������+X�e��b����^p�t�'"�)�+]p[�4_Fʭ���T>H0y���NUɲ�XU̘��|�>�}�GYQ���c8�tQ����C1���������ռ&��up@��a,K7���4tV�x�;���]۔{�li*.|ȁp��n���otv�K�����Z��?��Լ��8�\�W�M��L_�S=���e�����ۘ�᲎gf���͸ش�[A
:{�f�I:G�pݞ�ajX��Ns\��Xb����|��V⧕	�A��9Z�x�� ��+���|�L.4g���R�$:IK���TŨ�WPD�Fq�u�?�I����Uh>�炈�<+O��_�jl��M��*Om3]nj��ٸ+ha/���rØ��>�׉�G���\��=(b�ܝჀ���̗�w�w~�a�45����Bg���Bwnxl�{!�E{J�mx/gs��v�8���I})�>Wc��`�����d�VR��Vm�/Z�!�9�d,� ��3�,MOs�H[���j��ː��,������=�A�;�R�4�9Q���}-q���J�	I�H�.�����ڶH����������d�ߵ�����$Va����ac-Z潰��+��!A3��e<��ܺ7�38�X��~k���}*>���؁�b�ƿ!�S��!������@��?���&䮋 .��,t�J4�x��R+>��l��xB 8:9����*�{����Q�3Ǌ<v�ez|��ʎ'F�Mqm?x�/7��P�FF�=@0`4�{p����Hn2sϻ��>l���&W�W�lh�b���&0]z�2�]�*D�F��{��*�n�f�\�A�� t7uՒ����:�Nmav:��jɱ
�s�	b��5��~A�H��a9�q����O��ĔPM�U�'qH9]���ev�&��[n��(1���e͞���sl0}�w$"tM��MS`��N�l#xťZ��-1�6��US~=���͡�u�%�?d��x� ��`B���j�[�r+�K�B֫?H�\I���F�FY�v�$�Oy��g��%U�e�W��*	�']f���P�'����#(̶�Y(ϛ�h��ϴ�N^x�1��ܳ2i_���K�}�psm;��6J�Ү�&̱A�.��QTuh�����D�50�IÆ�X�SmM@�Y,j�1��F��j���	99,�R_���A�ɕY�U�#�R[9�p��Y�=�%=��@f�̿� K�P�v��������)V�xr|�����T�:X}�&�p=���Ǔr��ݷ�K���<>r�:����y��_���'
0N�=��xrs������]������!e�ћXO$���m�t7�R+5�!H�?��=�F*r�̯Ԫ��[2��<C;�TOMp)���~Z�n�G6�.��:\�p�������]d��^oT�}�BW�&�⁪����1i��;���N��gp���c�vR����+��r X�������U)��!�[p]�1�~[%_�l��G�T������rl���M�b�؆��8Z�ê6��ۨ��=p�.6���<�N�Q���Y��?�W�Ğ��{Ϡ(���hp�Ou� ����W.��I��#r�qe�����F����-ed����z�S���)At�<u��>����a
�x����8OqN��N�� �h�N \��#���3O\��C�j�Uа'�2 z��0�2��X��
��Βw�Q|\���O�"���=�������Y�O���W\���ؑ���LXD\��N�(�r��������x��>P�\�e��mv�8��S�%J�܉�
��E	���[X3Q%�jȡ���N��E�'�iU8N�Y�l�����8�3L@����C�Y�p�l�쪼�H!�p8�Y#�EB5̥�]H�M4v�� j��`.�.�+�(��>2,���E��(k; �� �r'H���l06=z��B2t >�����.�v;�P��+ח89wGv��'�� H]Ψ+��f*�mH��{~�S�<�
�~,_Kha������Q�W��GO��#��4���*	mU!u��(S� J��m��ik�]��M-P���J�e!���dM�)�����	��#\v�rܺ�Nvڗ_^|��S[�/	a���徊��<�9q��
l�O�W���׿	'A�gHgRvI�;Jq��'I
�!�6�/t
&D�yF:�Dg�K/�Dx�7�H-���e�Vu� J�g�}��|�����%����_F���@�C����]��<����]��fMn�99+�܃��6>��g3���Ǫ���q٫���c'�\�\�:��_�3=* �G�S�B��;l����\88/��i%X�+1oV�̔A���*��qc�Vw*�]?%��MԨ�����!$<�Y�![Һ\���	�{fJ��S��t��/������l�����$��e�
�I�I�.G�Z�>qo c��.hWf��!K�b{!�JX�G�Vtd2P�p��G�,�.�u#��������4������/�����4�3�+D��3L�t#t黨˦B]���&��2�ߘb���R;���բ&;4�a�SEBg�v�o�>sL��u��{�1J�e�I���Ճ��5��@O�s�,��Gz�܉�t3|����tt�wj��f����䨌H�v����������^|bv�@#	ry��A���9���1>Ą��{�֔��@.�sR����UxB��o`�������
j�j��۾�j�'G���ꠠ�N�ۋ�����ҿ>�D�M`����� ]fI�x����"����}����!n��֚c�>����#�)�A̋�l��9�H\z�쒃#|3)��@�R\�����|J���IGc�z��G�l���G�&�F��ESb.�5hU;���ޔ��@3�ּ�mrX��Ь�G�����~�Z�B)d���r3��&���p�����K���(ٚusY@ϗ�|�m�m��XS�Chm��=�14ɳ����{G��I�����}���*a�8>}�.���c�� �2|b��Hj��@�c���ٴ���Eh[�NC��fc񻭠���f��.��P��C�(�n�=��܀P��$�^N��zPM����3����du��G��/��m�+�M�o�����) l�9v�쀮��8X�W�_TZ�?�ݩK��%�7�hI/c|�\�	T��)�:���Dl�����H�+L���y�i�G������~�b��T�L�v�-8{�n�� o��"��$)�/�V|������'�/j �~;����$.�A����,7?j�o��~
B����MOM4@�-rm��	�G��o�I��IT`:�Nc!:Gi��fPۥ���*^B9��nTu9Io�����v�`��c�|�����
�a����w�΃����z��(i�zK�T�,�!���y6�7<��m7/A�c������>�ȭ�@�0�:W^uhՁ�3�D$��3n}'mv��/CR-a���e��(��s��ZrWX)^~����4��R���K��Ѱ��K��\
}p�'�
�YP���.Of3fR�U��w�&+��M�,��e8�N$k�wNBuY*�G~����xZ��O&%�\��*��mw!���z�T�"��gZ�j�JS~gI{ ]?���_�&_���Y����j��պ�]Er��mq9�r�n)?�1N��]�п�PWi�sV�K2��D�*�]$j����1Hi{��g+餏���F��Pp��s���I:�R
��m��d��$�M4P2�'w��|S&�'�,���L�v_��nZݬ�lu6��	5��{�(���nC������)���Ow�3`2�{�Ƣ�1�R9Oy���=�)�)�V��=��.č/5(��<�����Ϧ-��;`�c]�&Qw|s��ĩ���JLm�8�����%vE^���~&�2����@�ŎG�h�?�.�3�׉$;�ʾ��7���#�=}��#� bh���p)�����{5�����x�Ï��a7#s�!��~������r��;yl^����ׅ���h#��oR>�/n_��M�����ψ���L�L���A�����| 捪�,�ޫ����\ӻ�0��1�ÃB�]�P����bTU��*���(��)�6Ļ��j�^bp�s$[�W�1;4�ʥ	�lң���dH����3Y�߽Bul.�����^R����
����6��!iL�qT-q^��D�	+��1Gqlvm
�"o\Y��[� #��Iӱ*�c�����s��INٶF�i2]���]<2���n�xf����0@Rٜ���󗵹n|=�R���O�8]���$�O$3��_�NG���$߂2����M]��� �v��<�<S�]Ƨpi�`� �2��>�3�m�A������"�G�SPx1�`k:�Uˀ+o�w&�W[�����
�MS�s��� 8�B�!*�m�YR6R�B�xL*��ze�V&�-� p�՝�巖/}�܍��=mV���6��bP�ѯT�ƅnT����"���`x��ܺ��!���`��׸ATEI�4ؑ�r��1ܵ���]��5~n:�!=T<��ō�mf0,
�6��	ވ�*vhz���ô@dk���9�A_�*g��v��6�H�r��&��X��ץ&����n���\aA�]�o������f�3�ܘ2��!�c��2? �����Po�uUQ�X܅m�Kw�t�w�hu��0=)�M4��^�m�~T���X��[��UG�w{:�{�,�U3!�<���ř������P�"q-eO�'���/3E���X=����Q٘�yb������/?w1_�g��*
Z�g��S�����{�q�v�mM��1���9��Z�B���NH#�$��2v�W���1������ѓ������B�7��V����P�5�U� %���m�XAv<�%�a֏�_���z=���kd�P鯮����m����~�̄��x�,�����vJ1����dU�E�����p����\��{�$-"K��h��G-�WN�/���ī��e���!�X8\+��mq�.*�;{])C�śH�;z�}O�Rq�W�\�:M��ym���FAː�"�^C#����. ��)*��X��T��^���w�ȼ/@󴖘�tD_!�63è�8{$C�/�Ӣx8kK��88)F��3�E(%�rS��0^��\�q0�����L��K���dp��V�R�DhE&�lu���ㄑ��?�nSD�'6-JM+>ȟO�o+ �(awl�����3�B��W�_ ��������f΂�
I�+?��1��yw�(r�s�ާ<и�X$8�#n��������
)Z���AAi��̓�a�x�u��l��^�3�~�2Q�;w	0��vB���)���A�4��\�����غ����q���f���b<�/睡oB���"����C,�+�P��4�O�*���
=d�@�m�*��g ��{�#/����|��q����>l�2W�S��nl�f?j�I�'B�+���OӀ[�3����k���TlJi��`=m۔SQ�
/Ӛ.��՘x���mrFH��?����O<�GB���6�V��\�]�t%�M���S;˰�eG]#��