`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2368)
`protect data_block
0USWSUGxovGsyBJteYpEodqo/Ly3HSX186Lc4hUMZgb+BU5QFq3+qXara3XSdTasj79AiB4ISzEK
W/A6quPKaZWc8CzGGnm8029kblQnD0j8N5eFxTEwarDdvfDmKQ8DX77aYFyWZtrFK5EnAYeYbPfa
Czutv56s2ugbWQqStDgb+XYEkxUeL2UlJTKnR4OkRBzupiXNOGo8cP465xrUl/UBW/ebOJg9qR5o
g53hSZTB1iPeYB04vXncFmbAFqu/rp5Bt0//OH2SecE7qYAufIwENG7EYU2H//uvKo/F/gOmUrhs
2qYq8/vNnOgkhK+N+GOoZnpa37M9sXu9HGJBEGSz1uLo2EajhYyM0zlmTkGNg2ODyUPCoGsF+fgD
tGF4Dxs1E30XMqCYRJSI7xHoKHcink1qSXnnx28SOH89av53kof+X4ks2AVakuWTzpraK1O6fn9D
qFK5V3Q24xJYd9pmhhh2YbIbDQK5LOnavx7jQ6A2nkaErqdSuYfpDSTx47XLENtoOUn8SoHaCiFK
Hc8+cVW3pGnoVGPxEmEXGk2Yurxjk3wT8Lcf0QT8yzYz3fYJPgpMQ6aCyn51wyjBW3usYXMxIClt
jt9EqcZd+cyMI3AbrvdehJp/qajKHUdb6C/xiU2gXOaNYN1Lz68Wwj7cGuruwgHUH4ySVwNvodl3
ioQ37APMH1pZEioW7HsB5q2pHCBgmQShEC0FhMr3RIRPFEDS5jcyonP7NYmmJDaudrdmZiD8OtJN
rPKVcauNdU3EuhyBBH44fIvxvMfm2oim4bM6VXA5CNav06PpTpD3IuQ/hy8ua28fOBuyBY/41ccW
9sFKThjkrh1SrTpiYVAfZHXWn1DvYPCORQBC+P42gQTUCvrK+CjTIpb0B3qYKBfyAVQRFChMfvwj
8S3BMlb7/H5AiY9io7OLIh9AT30syx6cW6twQ+T41pdU4YYy+pPInYyN5pDmyjzqlcPZ9me5YTa9
CRA6fmR10MHtsc1HaD61EkjAH9vSGxjwZH28CA44EaHpQdD1bbl+s0BIxm37YmVI6lZLPXsVm1At
QxIfz7jyvPtehTLmlHfKyTatgGEbpjJww80lYsSiRC07bVjXgIkk2J6OQzL/tADq7fnInwL5Fcfd
YYc7xHo6+bO2BrP+hrD0eaHPfatSrF+eFwB2pKJUxS6b7B1C7rMQD7dVSPBy5bKHP0s+a18PLf2/
i9TkeZ5d6GZkvDlmHO2LEXDxL2dTFGzvhguC0JqTXYNjgQUHzOiNU/QOUF5IbrC730v0xTDy46Ot
Rb9y0DYQPZwlzVUz4GRfsA+1FlS+fgfLQhOONfRDOV5tdDpcUtxTIrxYPTITG2r6NrI293fMI6AK
ulYPhx1UzsoPZr3W7BVHsWrZbmZ10h9qOb8XvCFqN16mHvIkNvl90AK9ZA95WxYoGN4tRB4Ey2Jw
lpG4tmn5Iilhto4Yu4f8+c8Gr6w/wskN6WhYiiwQ0U8ye8iwRpG7zMvCMR0c8A9RvvZQxGX7c/xd
OolZoq1iId5nIj6ptKTDXOOTXwYO5I/0j9my2CPzfjRASCLtZD67f2dShGlQ7GuHqvSg7oCxN9zX
SLwVXAcFj5SMCI1qEKhBQSUop/2chjwdT2MdfX9AgUjkTj2uGU4MMQhEYqRXy/i8gTrOVGmYXKqm
+T2I5lAYaJ7mlrC05EE+BO0Fh4IVNuJs/fmw2x8q5gyF3K39i6rIGUG9konX6iKKKo8ey+jKQR2I
3R8M95FJaStjzE+kta660EKdSHe8enaZNyWsyNy2l5QxlvIIlKbvIQjHwrMl3FuCGsoH0HmL6C3L
2b/5fG1XHAxT/As3ql1UR5OBODzK5279+kyfrkhM1RTPycrXY2TNR3+e8/wg3DxGWasvWg/XkmHP
fMDWrcSm4bV04iS+dQNHrD9FP1oSzRQY2+iJ1lNeFQlfXfxhw4m0NxnpsWSxT9R4yfe9aqpeTsPC
3FJVY4m/xVk0hNNQi9nclRlUIszt8CR4RDkisV2Fhd90LruYcgtQJZqTidwIvui3W2x5UFqlROnO
q/DvtwsBBNOLVGhUHGUALNdZJXhP1vVMgGF3F8EzrrDumIUMXaoB/frRglkyfnWyvnPd4y0Mk44j
eGma+RDT5LJERl6lHUYKyLpu1145EMq0bEw7piMUVUvD6B3bsus3DhbCU40n7ASQqnpqEM8E3ko4
/qYU0fTvn0OD4wWIfEDAPue4JjIanzN53E9c1AeEj8w2NmkgsKYCc3ydsldxHNQ043pkkVLOH0EI
ZmpJyXc6cAsy6BNZQ0QOtpXPQVNKSCJE5TRMfsgTMt+7OmxqCrI3MVShJqLrj6OLTCrT6UokSLBE
WIZPJe+qF+fo2ifIRkZ40ZB+UBEXGpGNa9Ns3JU67N6a1hVVxP6F50B2Cv9fIFgWKWq12Q6Z7irs
Dt2GUIKUH1LQMTFYlouYgQI6Oakgq1PoLUCzAfavCeNQVkDJmJdxflENLmYsTo1u/bC2dC2upvcy
pOHAGqEQBwKsMisDPKUUAOJCRZlGvlL55+iG06CjJTTEcX2Md6b7PTrVik6zsIPHAhJxeA2N6miA
fOogy14LPiLZMqUDUUsIrihayeW5XeKBMF/8QXlibyBau5ArOlRWxo55QKtwM+H0hZKdHBWlRMPO
pE2Hj+R7jFCkdfiqRCdqPnQ5SC4k0zvC7Ck9jmouYCMyEtNyQtjOdJjA5OGuk040SAASwbn5jxcF
zYvQyvbu4olGfF9jOYQcuY3HKf4jZTJlr3cPqRrSnmcPcR1QbsWlq0IUeqkUewqoP+BplVr8bxWr
srYijZnnKJTJVznbtxSRyrO8uuLr6jeftWN33+iMA/EcDoSPbdOUsO5C0de/o8Zr4D9THDb0l32L
mH3kl+3Hqm9fHWgnhof9lB3b8sN9Y5AjMiapsKoyPY6zeWX9NtQt3sPqIla1Re8+rFXElbLZNbHf
33wblHv92E6l7dt792DWQBh3l3HDqAZ6j3BpAclhrzJetnxw+RgN2G16a/O9fVyWiK10bzRsi+is
iIhjItorYdOqNzP2h7IAdkXbswXkb1WCoCPN7tUxj2e4rQpatZ0r1KlXSKubIDy9Pu8RDymdMLfJ
+GwLLK5HCz4KB6vwAD5i0JILDE00cBk2uoSWx84tPw==
`protect end_protected
