`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3840)
`protect data_block
KNL7ve1Nx5eOyoElBAUwVHUDqSLbZrtAqIEknptf89vyhXz1WbEGvQ/ayxrGaPJB289sud7nBWon
sSmhCTdWWgbcoJAUhiOpp+GmT1CDrKYt6Vc110WfXtSYa19zfg70yG7dTB82NDoU24fsA5UB6NUv
8I+w9A19mBfUHJPhF8iY6DeTm2d+vuHeVuoWTa1lLyCibYC7HfWbAmBYwfiUG+OSZ3IJkAwQMHeD
rL8STHpHe6pHZG2cgW0xDBIWNS0by2RaLvEU6Kvlz2ZSZy4Bmw7/yZ8fAuGDxbFy0Q0l0TRFNHke
uFy89mZ4aWHRwdeGXND6AxfCTT5r9yEOCGL/bfwiGCn0Z8GAxDAr5uIWb715+wefo0ICWFwOiLgs
3kfPtWYk5B9idEuCL4ADwgl39/bwpnJmZwxLUZvu+snbQNWBLA5mhF4/rWZL0mRTsC8PJGFe+MBC
4JBvAKgY3I7qi0nuHkXxue3ZrKDL6uiHtZuzj/TfPdYRlff1XqIPtCvGIjdkMfvx6cx4EVcuAf7v
LsI4YO/07aBlaQ6ggPApWEb3fTjZDSOumfzUAvVmk9apsBKxDh6U1f1oAMhBfMhQ1jYcOMaqERPs
4avyOfSswf9ZLpE8cziA7fvU+uIrCXu7bqjYDaF4P58voD/pKzkrY/Fg73HROE7qP9gBhICVwl9+
Ljy7a15CLohrfjhA9E5z5VPk9g5OANbDkeCv+xKp1xcDJq4xwN8bsl6q2Z8PcbhIW+ARoldVItHO
YFoKrCRDyiLIte1I5mT7fhrcE4qUbs6oHmdefvjtQ8x/fo/sM8Z4NbJHtDJUvn6k+0OsphsPIxkI
1QGksjx4mSJXJpnL1PYO9SOTtpPHmZoEzh//XzGJ+JH8Lxpgso7XpLZPjNVeKYbOEBUo02xBH61s
sTbyLUVVD5EefRXS4P8z89eqifCMPwhs/O0N/0k9TzMPa3BSvsLA9LU0ft/pQqYLXLNKZKu9irNl
1I7Z0yksnEg45UNSvQJpmf0Qji2pAih7Uwv12WrAGyBfzPoBAXQwJsraHh9Nvv8MOkYD9hufuU/G
eyH6+Q1LVxDaeocWCvHPbYvD70cX8V3gAlEIsAcGAEiKMdoEvanBgY2HL/aT2g3OQFYZERDN7hyD
zYAIEhLec6iXD93dU+/2eC9y+F05hrq8sW+nj/ulBc47QBTUIOyYl83MdtlfbUdS4Z6zEqxnHb18
hy1gVzJr3LFF7qfeCUUBgFQlhuEKWxEEM0tz10IPJYsTPcu2uh+um70BRduU8vky3HifvHODS6zT
seLwX4LuT8mvA1GwR3aSSowKWcdsV/KwSizWOdjnwVmDlhjyVXv5+aeIBReupZIdizH23QLomEHC
WCvWK0uRg0v4DKR9vjVv4YWNEiiwW4wT1YkwlIHc2FZp9dpjHARvw1xdCvvqaYjztfNccD9eM1oH
NWsYUlXFYuzgDjeno8Pon/MiVPpKEpa4+P1vBYYP3vtcWAilxUDTl9vB86kWmBnU2VXyfvqDI84Z
FkC9hW8ETWkX93EUnSbdCREUAK0Cstka+z2a7rUtKXVEldJbRqnvffP+5QAbdXXAGljvCBDMIyeV
WwEpVkTGUlYyC0RgSfc9ZFEjWcefeUcAr0MXs/TD1+3fOSac0vcV5SLSk4GAvfaoazkPFo8yO8h2
J1oFGG3+dz3E5ojyGru79fY22sW7sEvk906F8pY9S7Ml4eiF1C2DkYddy18r3YzM4ubRUAuunMod
iuFVX6KSziEYNx4lfxaZx0AO1D1i0w6f9M+lMnHvoyb5P7496I4xX/Rql2FYjzYhGlEYj+bUeZp/
LEss/38D540Gyn17tOk+ESDEThVP4PzRHu8ciloyTk263v/fDpB2/umuh3bY5Yn0MrJ30C2oLWSy
wla2Rfx5aE9zCqdn/JvYEtCA95eT53w2PqUZnMMDcr4wfa0Suc/upHEevlZFnn2wlH8muV6CIl7Z
bTkP6KIRJaCEuHlLVlVWF54IWLFXAh7Jia8rR4Fu/y+RfOx6rqRQXb061gjK+uPPwpIepzNdiqC+
IKsVHp8ADJiY321TiRoNrGYqvGL6AO9eVqdaolYBC2OCzgDV+GC4eVwDjRQ/kp6x9iWYADG+9eQT
IsfQdbTI/nWCuWrUpls/UvvhOpXQZSR8k+VYuXw/u6EJcf/Bfld0xDNWfZLkwNocZ+lOM12LMXi9
f+AgTKGOWPV6jU07EkgIEzFgUKGOIfZTND5Tp+Eaf+R6JNrY2ZfCbZy0DTPvPlrEe16lCV28hk4M
ubOqOvg60pIuaTDBIQqGsW70g3sxLi2XOLzWsv4n6mmeNBh+18H6JdeLT7J5qXdLMAhP9tfRTlyu
xF+qtJNVjvSiQrwCuY+aWVu6cM9PxneYf4HWv2JRjDLgQSBi0s6fkLlFmu2WNu9oVu6VULv8wkk3
1bMd4aAFddOAFa3d+inzaAmeREtAd1H7VZlqny7lD2AYn8TVCigcx8xte/l41b0osWQ3UNyO9VbK
w1PYwRM2LXahJZADUrD2XIzo1cHASdHY892E8+NYfkjcZxpF58eQCVuKJDL9DmXUi4h3w27fu5NW
9ROJpD01tqfixxFlsbVDinn57LYdt+uhRHpzZ0UPB/GhKjN3FyZR5SKVt8TZ0FURvVTyQjZKujhJ
RmB/xxRHxTzHivzhVpeaTuJKrCBWPlsg43PDV/Fier/nePCBeQoOv5gkV7ZB1a1DY5dkV+w5zY+R
t+ZY/VN5Pgny0UnoImbi0iE6dRxSL+jB9v57iBY5i+E1gZYpOQuRxOXgTtXsKu9JN5EZJOrVsUKx
eV0x5F8GgXWHPfHzw3UzPrTOIWzcgGlha3a63LHBsPyK0ASTiVPiGriuCSVAk3FQDjdBm29oQrYh
3yCdb8RPLD06XR1GgV+U7B4OGNwE3qSijLE0HyRlSsI9c0zCK4rvdPRXgeeXThn0GBwAa3k/4G1n
B+NbnyZLCJblO2nEB6X1AkhiZJslqh8YExzz4T6EvvV4OiRFLQbMwFFJ7yGiJhxuNovatW3su6DB
kd3LumBJ32LuVRe4056xzlacVBJsGpM8O0UPljWQh0u6sCHHhxOYuD3Iq4LbiYmpqgUS93qU89ef
ihFjTZKHST5MiFt21E+f9m8+AEN57yde/TgNcvhrMOFeO8lhm+jVLz+vovjIZoeiioNSJEEb1+Gc
RKtPF3hw/nINClzGOorQ9q7hoYfKe+LoCBML1JUb94g3SidRfzhZX2DXnOzAd3HJe1L8gOz6iWrx
5uZTHGgJGLUhsIn1oMu0nMQ2N8TDa9Oc/UTk4tCWiouAQeEGL9mqGDbRbupjV1XmBoyipNxGEGzw
7zcFSY6cL0JkqMb39+OcI9zCsbF23I2MBR3xotdyM0HNOTDGoFcRH3+aQGV+uqAbvq/e0/Ljn089
aoZW6T8RxklW1qpXWNHiW7NwbHV0pxSmSVhOmM/ArSQM8HIME1upz4HXsIPiw/H6Hav6rpVOK38R
+8TckHAGuXpkzwZLXPW87TH6PQeZqWTkbuBbXenWrqMaMJWlGbPBSEgsF8e9DTZepCB/NDPsuF+r
OXWOv2Cz7pv9cPLHfl76gU+YZF24ncqUDhnJit0RKZQ5Mz3/5AP2Ijn9TNfa0n5EgH7dSD39l1AH
T6oh5jaiMshNvOhzxVAWbI03ZOxVhw1PN4vpp7G0+AgDvgVjYWhPZqdZVSM3pFpElYuDKMRFTwxM
iD+Mq++ndY/HP2lp3KxnlPCIfT8UKVcFe9WqRM9b9s363sa6rklM6UDOZGGD1NRTMW3P8h9iZJpA
3WErK/BQ+VxSC/0CmMYD1MosZ/rWdc/YvyFqoxxZP45uCXZXdv38oiEkzLzPdSaWGZtJQEhJZ4S+
mbDPCMk0+fj24x2xEcrjzaZB8A9zYtgzdMM/SL+aEJWxm/jcBuwpStmeiVlHGmHuBY/AM4i8siu/
JjgSmr20ApQhJS5U+8C8SINAMADO4pOFJbglviKgpzRW7/otUsqGlvTfSMDEpHs6rNr8TsZVym0a
1cdgqNpaReBeMQZuVD4HXrO2Trh9Aq051jzNfs5sW7DcFZ4YooFYTym1v0e3XNRl5xj6b+4+hP52
o1SkeHg04dVo5lwCTpvj9yXwzToIwHhmbdKRahtGKMyJpEGGR1lPQtEmezyaKt/5/PdjUrfXjLow
/msgBGksWWZg2NDrWrMSj2fLQkZyuZl3AmdHskfZMAxhTv/9lKbVWbo6zy8eP1X44zac3h/Ljbru
TaEHqoAZr8KDklFUDwP1QKQCP0v+YIW/ImphNKS16m7bLiPono5drxdfEO98ZbEmGJOY7bfrgEie
3mGNFIB+Pxso5Ku3d0/Q7ONKXKlUG0qBKe6eUDClz9XJWCWQu02tk3F+YRZCTsY9nURrCrS2GM+U
xL0LHFI5NbiCD93LfbFY65DNIpIoH+w+i0NYP1Cb20hRNMdBiGLm+wemto5q5svXDbFSSMoyjRZs
AEVT9MCIA6WHKGGod3V60glZDcMbMkfW2wDsjTS2ZsUf+urBuib0PaDMY+E64arGZ1nfM9RhDi+h
hDQAdh55ewnv/9Y396nRr0nBLTAtmDBR/soPb/2HXgEkMl+rF40vvJshuLI+LKXhCk7jlfOJJUO3
zMgnOx65rl19QNUi0KOprk27Zx9UJrkCaJ1pFqokhx5Ngk62O8F3eB/dG+s27ftfimXELDJqlR3L
/VrvSSRA3MD0oSN6YQ+UgepqivBUYPOeeNaii0yN1R8xRy6FVsbbEb8h0P8YJPJE4dztCyiyZ3g1
kWYuuXLOKd5rpqCEpu6mS00einwkODasxgMbvsGAYZc9FjnU4f62TzSFJl06tQA1o44xlTiTiTvn
2hpaaOwK2v3qM2AzwkIeB6mXLV4JfGYEmrBhxKQVDC2HeZIs/VAcOgk+nNrD8pheJo4xs4dEz4ew
aJtDh7S8+ts8YgErmj0G2MLJJBdVTJSqrdPfzBiGTQhjd8nMoOlUnafom7S/kxJIPT47KYJWsydy
g0FWzmF9nNWGwOqPNS34O1pY51hxMXacQSc/UzD8wlSpbMMlv+UX6liqkSz+KOkELuPW7fpeGl7y
UcyikAC/MPA5DV8Q2Uuit5cxUuWS
`protect end_protected
