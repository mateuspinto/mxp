`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
K366Lije/Xc9UdXJ21HwLZZqrTsGpZYsoaLjyaATHbfdr7d5zy4i3qLdrQaE+CQv9cdE95aT4Hq2
3CF5v/p29V++iYVE0AcT/OzJUFvGZZlGOBMPI4H8svcbv4DVYvn992BNn71jdR9J4SO6KJ+eSEcA
zTAeWSFTN3Dd6be6tm7iUIHiKeXXq0CSC/OOOBszE9Qg502QZ1Yq4gehCBAEyq0MglRkFxNxrimU
ZZ0lhLqU0JIx5SAou3cTYgY0/58plDJIXY0/pGQ3ipCtBR69Ha3CTXsOeHIfLuGpMh8YfbfpNCpV
DJr9oHp3xjJo/M1aJwVQ4DjomKZPR3TV5Y+VOg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="j3gNw56rYVn+0VLuDDX3TN/oA2sWsBuZnvpYW3xU5EA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9328)
`protect data_block
CBRdkTv4+h50VOFMl0r3uSt3BJmg05BKlO+kKeElAzZfQBoqZni5SUvgMu5uHafF1o0AV3S+dec0
cUVZ2/8uez6cv5uK99TNmB2fwjcQ5scuVfN35px2Wpte+49Z3DeCLlFR5JQJN9IH9drsK4uoz16G
IHC9ZesRUiOuyUOLr+WutW8YC7K18Uf6rx4L0JDjrQGJf4vlUk11oUfu6dY7cRNCytZN9z/kXr8h
+4w5DT5QpMH0FAaeVLJroLHQ8JFi/F173JdvIW3oX//qUnwLaN21CaXDl1JX6/5h5W15ihFqFddY
KxRVR+0XyzEs71VWvnEK7DjKdONp8+3T3iBNLasCUKtKF4DSnRT8dpsvbsAwUr+6M/o12SeA0AY0
ozfNKSO0tGx0JcVQdHyeNZThZK/NAXNv7SmbyNMvac6x60d03EMJUjbmwenc6p9JtIbRAQdyUAEH
WUNDv2aJ+QNCcUjTEK9AgxTcXPJuRd0JBTJyJXO31q2tjkSFcWw/Nz4QBKmdtQgERtkiIHinGIrx
ggrQkKgNWKQtVrqqWkHENBAUjIU+mrocfYEtjYDtbECLqNIu8xhj143TRpbwSzTYjjPrwXHPR+tr
XC/5rnCjSzW3/MlJYoCk6NNuKmbP1O1aO9xZsqWg8o4ByjlGHyen7SiiujiMzC2k1pCWB2eAfnll
H050nUTn1G2waL+z58pLs5aR87d0+Xvs13PQEJ+n5iL1jHEkhb3IqspOcPAD3bU7NkjAHQ9SaYFl
jeAwd4nvjQStzkmpcB7TRz+MZSqw4ZnJKVdREGyE6wjRTuSFmyMM8j+znHMcqONh3cJcotwuMh2/
tzgov97uFeykF6h8tFuErgPmxgKbYnlqOPPTsiFVTIhBJfckIipCp+AmgBrXUBU+RRMjpjKcp0Lt
4RfGR8/7bme0Mfhrs3sBSgqlj1qOdy6IZKUp2QuTD76dlKo+rCjManoHS40tYJUB3bXWKaGvVz6G
lw3fkYHTpf/pDeqFPqqNujpMl75fe4yAkJYs3mDV1tNpCsHaOJt15SHmTXB9f+61MOkbgAwqGYOV
cfDCX+CJC3rBw9BXVKCuCo9MZDijf4SpJ/0ZnWLfLxPVjVzZv70pXSuUwSa+NF60vcUqb5AOGZoy
CzHV1bO4Swx+P02c+yDlAgsZJKy+x5/QLX2YEPBZHnDgDfXMKAWsXZJetOivF9KiOqb6ft+S/j+x
LC+0lo4AKiM2i7W35FDGkvaORiBmMW2/PC8h7Jy9iqcdMjCoYyv1Gviu1LjmQCIgKQGvFlKLS2Iq
d1p5G3fYScBKLemR3pgUCU/QkJHhL+k299N9QbuikhAI2cxQEmnN5xfATz6bhD8/OQm0PmAjKCIH
UBjSiydhuQloA5lcmOb8paADoe3kRGitw1QfWarsH/59O6CQmV1ziQrIv9wcYGwa1mDJ1C0iuE5F
3GFHSxQSuBT17xrPecqQLhCd6pxsM8y2KHUJLkk+g2/73PUHkJRK2KSYM8BG5QgTXIWDzW6DuADA
QIwG+jP/FxUR3OPjzEKxru1qfegaFnusEdApetTigAmrNv8t0UsFQJbmvztimSWJrXX8kjclpa0E
hySiO5Pk5h5gGvboir1NQKzQ03BGw6G4HIGZtOPZAsyp+bSa9ogdC/ZAetRJ/GXJCJ/J9dGElwY0
lRy8VpyiM5PZ+sm2721KBncoHI9ao/5mY2RP1tGMdeqmjyWj/w21/8ZCTaY7Bk6lA3qM1Bwtbx1l
pHhM918bymTMDWc1ciul/g6+HloRfYYnXlLBUEaKwFynppasEV1EG7JZLrXeNBcc9tZAAc3oh3vR
QG+toasLqCAg2nvllYB0g7cHyDFOqkm0L6FPExOIxNif5aw2Yfler6t5CeKLD+WdD2OJHmVT1/7f
6sxt70g8bCjmNZmztxnONeYMS69HejEpsy9u0xW4XiwWSmvLPqPeOyAlWszAm/4Gd+6twwqD1hWi
CPOuDqBSTnpjfGXFaeMH1dHt/ZnSIGcz2an+jy5+UxwnosjNoYWAWQB6xLpqaK/LbWfM3RAg6aAD
Fi37u2ExYv8w+ukw6AlJsNWHteaAhky79kTSj++iwdKPpAC8of4Tm7AeLKfnt2Zn0p9ZzoAwnDIH
OsxGLYRPUQPNEq9IujUPgPU3NiidWWMVOVUFf8C5OSx4XucGYRSr0JfQISzCGg//8GfBmLWYC1qG
yFZL/FxM+GOWFC5Afd73bqhlGOV+duTPLbx8OVv3Y3qYfZLfmHQLibPk9PjkZx888WjtEBUgQfB4
UScfGFVlKRpjfxfcB6cX+/g3lrKoooAkV42qIjx1WOz6qylSy7EDe80OArMYTJvd17K6fV9jXxz5
5vsVcpZANWz/d9gMfw4dTfxnW6FD9fxUfWeIaGNO+V2XfykXMkLDAMBc5wvzJvr237diImhkggMs
wV1T+InJX7U1LJmyPVrmaD4WawCHrRgbwX6JUrZMsENSby0pLLo2oMP5anUkGYkEdXWHBlT+7q1N
6xLIWb1+VYBJQiC51O1vkhjdaw7iZRa/VE8oOVeLincO6c9Y2GAIWPrDhdMWmlQ0yP60UWkbxBMI
5vsZ1FDFRWnmNPIW/TEzE/9G/zLqGIKSql4xuOYBA6LQFD4i9l+cEg3vIs8BF1/5Dhbk+RhykUUO
qF/FUwbODAHHFC8XA89LPugs2tHddoXJO9F6bgYyzYYSiv8qDMMIYDvisTPBapurS0DxJKmtYZqe
mM69QD32PMBinDZVTnJW1prfLSSJ/1wkEsONPxlG/g4HpDFyqwDb1V7Iie4OoHZq71hfkOa2iP0y
hUOMKmu+dl/AEkROaubNfOZGEIprTlp/NwseUSG+xKANKyXpnpqfoDTgrP6P+WmBEDW4weGUhant
6G//z9XalYV+hgNzin/SlJuJ8L9/1/UrmldwekxjPVTItCBJiD1TDIsLXsUbVDAvaXqHqjXO1RlD
5cOcQfF2dt2OZIllKHiN1SROLZUnJja0jekuLpRTIVvGU4erN0AIVA0+5MEp3LcfonmwLOuEt7Q+
Iwi7uSamLBH5GfiWHHTsgDQZRIfPE4OUezs6pC0lDn10q3fBDi9GpZEqRI5n/Rnb4N4Hd05Ea4bZ
78EFFPB3ylS+QBMQ313AcruY9uLXiAs9wbGB3DcXFtX9gXzs87R1JU4+gyOSuFt+sVwPg7BEd76v
eG6WOt/JYUNujGGKZnkbf2kMdDAXdsRk66ddvpqY5HrhjUBnRz5GUyqE7F/FtZh6BGnnnmP2u6VZ
ji9gc7pBv3i1ciyIWSlg8W2gaRiR3JXTzB6R6H5RT9iOuXRDmf0JBtMmauDVUGY6OigBWDbGJ0sz
ESXp7MgzqKZdN+VmUTvYxvVGWK3QDBCVyHwI2sZyDqdimgu3G/3VWNErVjqOZreqHS60y8ZOtbzN
FIyBfaNyQLIg+vl9qbTBAACfSm0ihfIaDCWdlxnScWEwkBI/pFxXMMM1wTjo8Ap2giffuA8Lk9Hz
kkQb3pFDjc0Z44TPOI1C3wVeerl085OnQPkpki8qO19b6k2yNJO1OSCeVl4pgg5m0dO4hvxM8sJD
y6rxmkyzIpN76VCPxOkXLwkKCG/vOCImbfY3FarW7lSziE3SWvXbNcw4gzR8iev7xPEsHau8TAvG
Ngl3kMYfyxX+okzjLlvvkrwtBRRSA4YGSQsjeZY+MQd85WPaWz10HP+NTxsETm4ne5aMhlbE4iMD
+2NU9w/TshxDBG6H7b+yIdENpqny3sRYE1edsfio4fPG5L+MzpHCN06UgvOcM1g9qDNxDq6vaal9
HxFvuTAfnYm1yT9sXit8+S6LMWUJDjQgCQSbzVnzYMi/0P9YWaSFTGCBcon8Y3Fknnk6+N40aYrm
1iP3RBg36tgP/0fi0TGLTuyUsPJIyruwsFfdcZPKpyOnyvQW9O8wxvUIh66/3i+SfGsShmAcpDtC
2VOLaY5FM7EUq/Eh1hl0gFGircFp8jnycAzhJewVRVvlx78TOHmfgGdQDZvRqhpVYLXcPC77H1hP
nF7LS++CMJP2H7WkFhLGLZVdYWohSF6CT17+XLLMukGazX+tqUSMEY1nva0NQjJBQOHRwwoo9/6G
HTIJmc2yQicY2BAUulKMLomjWwTxcInfbqUyyHMBApHAt4QxCxrZOjcpW7y1ou6NbHSpLBKefNLi
/Qz6UlhMurCZwY2hlNcUBE8Yp7JqHslONbS/7rljLA0EOVDFFlmndugTC7RoRO5oOnaMWRXtOzqj
Zar9yZT4uQalhXvLatVZzWQ6xGbruLe+GAQ+By9/zWLrUrbAhEenwa02NDIanQlfX2YpWxQLwBjC
hTC4gRLZVNl+0UAc6n7/1/RzMoB4fdvIc3el3Qb1cgRbxnbj0QScKmz6TQMTvwKuovPMU4roym/b
sI8267ynshit95m1I/5qq4oLEEvX/C97B8wzYtC+J6NbtlbgfMZRWCRkjCJFYLmoym8Z58msO/EU
mVywK3IlgMp4zA/JTmHTaF+MttT801Ky49Bg0TBx0jvepYEDtoK7Aozx1wIJGuO6g1dOY9PwXnIc
hPIiwiPVKAKnJGnEP1pfCMQB6CHHcTZUuJ+EbTdFEPhv+RBqA6NDIYowaZ8Z7Da6QdTKHLBs/jZF
Q8jPNumDFFVRC5tt+fJuOIASDLLzQI/mj+kjyb8+tgSX/VEsT7+c7dQ5SLGjM3L3y/Z+RRayQt6v
Oqn4zSwXYf9S3EkBicQyG6g0CmVRyVnwAx4n2xgBIpdKkWwRTM9U0QZnqm+KE+PtFDx5oeqM4PDF
7AfUorWpCTximdMxyDu5X9FWGcErg2GPvtSAmDmnaSSGXupoasd/Uk8YZ4An3AzrwTGTuYqPcqft
Vj0uh6LDo+j0EyKxWVpVfYvG+ohE//ru5ezBq6IuWmeVhLa11YQFHxXhhQyZoloKZPISKRY5FWE2
B3iOP0q+TvX8AKj7kC2EaZ4lIlPYDiFCB8Iwz3Vu5HfCymtbp+lInHO5Wlol+AMi7wpJXah+XDl5
Gcb7gZCFVcw3K9TWJ6HyPE4iAYe4IWoDvXVo9t0WxRrPLU9Xbd36SR41rhyvO8Tu7GUw9n9kwtP1
Lb9RfIpCfRA28v7aQtSLCX0BrJ2YzSvnz/vChF6YFHImRVOcngDFfKp9GA4tTm9ilrDNUHmBT38i
uRdQhaX9ctvolTkyachxj3+FdWa5x1K/X8++SJ4scNS/8G3heM0wu4dn+k/GJGaXZ8fMznuqAeYg
+Gv/427qVZbu04T957oLDfO1w6ph/t9vg2WY4LPd/Rh+UDlpl6i0Y9hVFz3/cQ896WHwjZ9SdR2K
hnvYp5sjmrEiwq37GG/ISGbYjiutsH1rFinDhqan6UNKVS37qr4j/PJ0ZFQVb0W4SMwUo8h49KT6
GxKbm3fRp/mA35SeEQ7X8XxXBMi5cmyoYr5YrhQBV0yCR7VeRFFJWvrP/M9skHxY4N6f2Q248NNg
OV0xWyx/UzbJoAkRxSr6WZJJu0uhteGXU1ACuwfTm/GkM8LI6alvD2Nyi+LuW5BmoQCdJZ8sgIan
vz2tvKJpPNwRWDU36JpydfFAfEAtBTr59oidmBDDeu0htdB8w7pUyvErRJIiyiJwEBwCg1ffHpT6
7cM/Ql8VLvH+GEy52S3JOxuFcqdobFWkdUEjnYpj1o9LbzFovKl3DENIvSTz6KuMxbSatCf0krsI
K3F3pMT+zAnJmS6Zge1cN906eDuKLUNSnbsoYGioG+UwCJnJGFMeXkJgC29Z/UUZlyIOf/SesBWN
H+Rmp3M6TYnymSGuHg2e8WVXvxuJpam9TsO+3qhVVeD4AsSlrDM3sLw+JcW5w0GNBULIQ1BQgjTi
9Fq4j2HanwX4VnBBQGr+IZAFjAsj0XrJEi9MGNu0xwsR+81B/jjEQcLrBjSFtnMM1LVqVP+BrLgG
+r8U6fRDKENs86YR+zuHpRJODxLfWbaVI242rIeuBDsSVMeQFTJ/QC54k5tM1Nq9smRL3anBF1VW
hPkw8tTUzd6HL9D59ZuVPE5Ykwqnfc6mAXqJwKtIJjruji+Z4v1+Uis6/sMNU3VTicR3odIkvqYv
7ut+uOsXyTo7dfmIe4nW7xyF1IbcfZmJcPF/muPP6Po1n7JbGbNdEGPv1D3SCoVefD4WrG/JXevQ
oNeycU9BL89WOey6aXlD1/MhRK/Dy19TL2Iet7CHGEKHLyc7LZ0gM7XWSuvFabucXsM976SqkTwS
vO/bj10u7064yvwGygItNTE7DaAop8Z9NKCB0CskeBnM/b20HDixWKSYOkD7FtiEjhd7GccY6q4J
fZWpuupQKXMmbIYQQSji3SoUzi9r8mPZt2gA04545mN0Av32KcLH3ys8g23ypEcblx4hjb4w5fp7
9wDJlxdcwfH+NbEkI3Sqw/KhDEX8Y1AdOkhNkox/OtwpVoCDvB06loLpH++nDTrtgxayw8apTjJJ
PKX2RJv5o5OexbspK/lSKI8EvHJd2xSKPPiKEwmTSd5hBfT7mzQvfJbrG3WJnzCJ0/LenR/XZA3t
OMEY4EUBqugE5EvmExRKgPoiRypwNRjvAffBZRmPsl30ZH/T0vuo3gmGn8uG3eXtE/fH0pXtDxsM
6CoSoA3IoqUY2x4JqMue+tK4Z2q89opHfb74Ea5oIiNVDVFhTvG2NlCYsAAYhjSiVus20DMijSil
fzJWAj3LNanvZixnm0nqeGZyASKVtq8c9aBojXpoc82kxlAQyiYalV46gqHkkJ/1lgWFb841ui4B
04YoVJxOtJM4lfjEWRXA9+kh65N8dTC45VpNpBPteibLmHBPLy+S+65p9KqZYEf1E84BR9C9TV4S
TmZb0mx2gk/c2G0WdyIoXuf1yICNBdPq62LYbyMOo6S4q+5wiUVBMwA4vfNAplGw49WwbJ5TxFAZ
/4mJtciCqFtaaHiC7zAPOXMTOxMnIGcqtqlFyMFH7PV4rfgIMaocNDKSJgJ+xu6aA2HEp3GOBAhz
cyLh/+zRiYRJwWtxQv4mtFBFwnCSzXzAvGvgGlsWQD16Arb9a/PBa9aoftpmfU24TkkvGxKIL2bH
OsFjJBMpmtWPxhXL5caMa+gcjHE79cu97P2BZ6Ec2rdG4WZQik+1JQzC74PjU8oBhEYMJ54NBHtm
IZXzCu+CNt1goGdWdzGI5O4GjVx3rjaCDumx0gLM0IQkDSmfbpZwVsIXPkdoMBYoh9lgRbDLfmOZ
Tt0CPb6CK5rPNdZAsblM4Ko4jaV+y6z0Sd62vYy0lkEROHIDjaQVL/HejDHoFVCXFoPPstUhKMJp
3h8p60m5E6haU0okBPio0qDi8AhVosCtx/ahaem0D1UANie7ijGM+gal+AmU+CBPGEKJsI4G4fej
uuPVo2hmYbIIOKgkqp0gua0SHmxzCgD4GxT8PlGDR1iIw5VTm6Gfay8LU4cDUJq+5R8splIOvV4L
7YXgJHHGEiVGlq2YGV4yb7v59g1UtIqWjdfbA69dUXWxYBwk9sz3owsGLFsISr9pNnOqr/UuUBBd
z7sCKjXkkgWGeSf8NM8A5W+QqyelTAoCduOUW29BgQ3R9Df0IZu/pjcvUdGdJgTgULu/XjJvLWbS
3TYMD8uS4vDQPHjTPkC8LaQL8OJS48cXyLf1EbCHS5dWg6df4Ltj5A5WGfVGf8So333lDYtrgJAo
svX5HgKkC4s6woEXvt7WO3CPUuEtppjLWZaSiPZeN/q5HvucvMFbF2rOKJATq0ez36I1s1zkEwm7
rgqFjDGdhNMHvu7k7HNpPhrl4yXC1X65CNSiGjsBimqhiDMHAzRoxxKc4QHUr52053mXeKXEg1Yo
hXhyGpmrLUBibD0eLAblNje8pe3yNO4peTnuvSNI9Bc6iV3onISKGeqjgP9FcQjNtpj9K3gUQY3v
s3grfK6LR/QKAAY/gdrKsrkSQv3OOVOS/oYzLEHFLBfBT+rKjOsFEwgXmmzAxihEI1ZfU6B0shDu
ZRcjwl77LSJCYcUqHBCOxFfGOi2d2E9ewYU42qqWU7GPq+AvqoJPqFREG0Jxnzz7/mUYGF+e6+Jw
MaXy29zaMqBn1o3A/oxoD6F6Ee0nQx4aG+TpbFj3LEEctOBMdDEWXoAfflq9wqIw8y0PPqV+emqY
3IY+XEtcN8aKnE5Pq5A1I8IWG4yQ8TqlgOt+8SyBM+6omOZGHERFr30X1I3vztmZx2TheaRjnagh
VxzDwEzp5PGPtne55Rs3QDp4dce8+1CoZfO8uv4X0raNyOqOL5p6OkqNMvfqkz4uRCbUCCkvmZWz
XEmVBNNhptLbhOvAgTXmqfX0LJIoxEcqGlLHPgsVPVUTL6lMj//2SG5P94N0fO4PspEWZ1aIM7Ei
vWmGUQXLvTqm21GNUhKihlIo+9oFmBapCvxONVuxhsWRACJYVCe1DOHQSZAOeO5TWTJcxJQgPeWt
qOvA7Pchcqfi7P8Xko3IPiU13wM4mDaWZqzXN9T2ZPVcxe0+6tEFInJggXKLRqGGrGnLwd6m9H1+
BP55QVWSY+3Qgn6o6uYjicasZLyvdoWOqDQAi3R8d8VNeC+W5Wg2ZjtXvFq6KpD2jAsrGKoEZ/WV
Ah82F0xTU/FIp1x/631KMPddd/abLeMCE5QfWZNYCNvf0El4v1MJ33kE4UtxE+bZj0GFfUEMhLxc
GyIgVjUWgGJT2FA1+AosHp+nRzmBCN7aj9ZM78czx73x36DoLXN9aU1CTLw+aeUZ9mpfGjd1mVEx
yjJNCDI0gCcoutCcBWPZoqTDnmTWI/1W+B84711JqjwGH0J6i8fi0GLyx3cqqLGbD1GSry2rqGlh
XfQ/u5Yb0q4x4a7O5ymVv3KeofyMQw+A3nGxhQukSZRPZyRLTgZfZHklrIuCxXlN4fmDnaSH+emK
jKN8kQuRw/F/caqpF1cwKk03HuMaPnhzLA7ReaU+q3VGRDAm4spj+etldVdtT02gYHAbCZwVB2wQ
sgy1ib2J5pEvTZqjrW4GpdCcuzJ5hbtEx/vXDEX7P7PPiWEMLFqm26c8IoCGpoFyF5KTXd6RFp6T
YnqsuocEpVADhRT7+c8LejPey6ZT98AY/Kkp4WGHEewP6d1GrG7oVDrMp/CqUlOffxVKfJZAdvTV
jPLJVGGJShx8L24XPTaGceNF5UJIA11t9mS80GfW8KsU/+aJVb07pha+9OdHTAitPciwG1ze1lVm
frm/iU2iVZtX88S73TUS7vSFoDc3UyqYIUnJzpUT2+9FgOkUcWXo6WZXwlQnI1tKm0eX8prTAsOM
lcqOtf12z8s4zj7a/zLMyBIlmm1J7RxdVbZBjitb32i/ce4Xir6gao176yl4YUDviNzb+OL6HLSU
xD4npDcpZ85vMYbOdF9/Dv0nkN6uh7fbWH/hir+SwdBegm8qGvvWkxSIkovZJGCJCEh4H1qo46+k
3XaojsEuRVVKYB0+BD/r4N2tRuexdk3gA6lgLC8bgpmY79nW6oCdh4Xpx/ObUPA4204fyyHF4WE4
i0BvaL59bUbFE70R23eajDTKnTkiHNLqv3rmvMRIYBxz2x4/uWfBtu7kZ7DqZFX189ADsmi+nODj
bTezssHaR3bWLIAhmokt6kilajqBNkHrwtVboT4eh7m5NI0CfBXYOntMV5K6LfMpfh5JTwSBVy9I
DdZsDihFgej66TrL5Itnt0922kKJ0bhOW+abzky4++3QpluyrnAP0e+k4wc4W3pB9RtHaAIQ9fOq
cFN5JUIVP25G7OC5++mAraUEMugrvIqD1dXJKiEKfuvAvmvFYmXzf3sr8OHjwauK7hOAFqhiy4gP
YvugHiG7zpu5nrqLh0Tq1FeT/3GBU/nn7KA/oUnD6c0elV/PhZOM3JWQ0HNZFvhZ4e9IpH3HjaSx
bpmw4rX+ZwGFQo92eNPZ1Rjbq64uZXzSIRkIsY5EFI6UcGpjzTOFyz+jAFuC8lTnPj3cxSGTSjpe
oLBVRcAvP+FwfZENZ2wQS+/EMNUKRWzE7fk/brhMdLagh7yjzY4+NLZBJsYoX34yzko9Payp1XoS
I17NvSdrLUBQBXsTVlLvub5wVrrTXttil//NWzqzWqO/CqzPqV1l465EGZS2rdSw2C0gXDwbaPQu
2SYO0FEPQK7krExXtCKyRkFNwUbxTAZ34MvtayUPVfjsfjiOUQs50w4pgPMflusS2jqZkAbwDrXi
l+CdyljfOGKKgbfcPHU4erHvO4sSjkuW4i6QPBTetMHlwLeXG71CK4tDTJyg158moWMRV8Hrkzsb
u90Vu03taNOzfwLqpLTW6tIQmSc9IQCMVASRfoCf1/RQoixtZtVIAIDniQSIzGQDmubHwPw+rIdM
2eOlBcVwbPGErziwo3q08IP8bPc8qlggK3Xu01Q+X8g5JEiMo0VF/ewWfyqbV03nOcdgEBwb9qrF
7t84Go36P9Yv+dNJLUFrUa8ZFyRcV8I1SFd4Yk1911Kaqbe37z2wgqSR0DINLJhjoBsmCXHAQMVw
QwrrLGANMosDJFp4csi5uQK+U3ONEijBGrirqeqLYSVPwEXyKoOBsCpKGgGvgZqZHKiZjO7wxcHc
e9Fil5T8CAsULWH8Egns7jkkpdBKTSMLjT28PKbS93YM84D0ksso3aTMi3NDDeE25YuFNVHpv3jK
XkUIXQiicQIcb6RC4khV/thWvIpJxRk3JicZ6/aO2SCzr3V1nZ/bdM8dGZ+6WJds06P11Xbjc4KH
wNXZEsQdqB/gEAkeGNvPcDehUZjNnnLUqc+AejqKwqBtIdTlosKO3EmHjjbtCshgX8TlJIwO3bY+
RaCHEWwrWq2FdMUGSv0ZLGUgwXM1B+AIFGr+Snlehcufn0jI7nawx+8NNFPFK4ImkWV3JiVsnQhM
LoPrpy+5EfXIcN0mewxU5t/V9m8p1AkSlUV4AG0bjLCATL++yupIGPMvMjjxZJJKgmTRhwjC5Uk/
FmrkCgXTpxPQo5f/1jrNrO7DCUMV/4F5gR3v38VCbrmebUp/Sfbki4iZ/X3RioppcEn/58x2GnrI
0YA3pvxK+0IWGinMQs7EZ8rPb3TGDH2RqJaarNdEcE0oTm1gkSZ+X5kQ55NWpCM6Hw01YYCgI5F1
mkkYNM3yHe5wEz9PKSiY9x+Zd2RV6BX6QEj4ykN5QA5uuSXUq/4I8qT4ky7DYif9b9aVwxyJcamg
cRpf4iUuPJ7PrEA5i500WOFJK7OW0lsN+uR1aU4aBLK1V9r5yAAxMkqJNLv7mVIQ3A3mZQYLd/pR
eWnq6VyQp9GDjH1BiKMpk827ICnQ02zCOnKfrfsqEsE0Q2jAsj8P0r1VrEwbVjVln1n5TFfE7dyz
0HCvdaqyK6giDgMveKwSvvjfMRsbinHQxOggsMq0fi3UVto9C54t+UyUHJKGIKz/WtlJ2vETX7Go
usnMYku4WXJQSfKqxQZYV76tqHce2K9dvG3/kuCnCsVupZpa7iUF31T61ga9uhC3BUcQxvDwVPwR
N9anjTBX0xnDHg5xNa9t3yIGc+Cer/tm3oEWGemXYZD+62nGCa7O2W/+3ktZm/qcppGbfzTfV3/L
zEZygu9Lqh75ZG7wBzY/RRi5HLuExPeDDK4dVZ7yJFHuLD6xehV27sR/CcEQ+EiuDipFmMCChvrB
knPPDAGtvu4DmtVH7wiQfL/FMl0p0X+xduNENEBsEEDbXFNmTMmPAYrGsnW+YJPjSpp/cP+TaE/r
Js0DF6Y6oSZPoX8Hqx3idSvbd0oFjrLuCYxkUv0thqhQSXfD4wLcMVg7Ysdbzhio2RAJLVLU5b8O
6aptaV+RVX+CoEeExkhkO+KNcPyxgCUueOsXNPkk9TzydKgURJQHbQtg3PbPXSEtvTEgmAgngikh
kM14gxDSAktTnWkM5LNYz3cCau1DuNYR9EV6hm23FUcOQiYn2bJx6q6agbwVXCZ+fdY7d4XcONPI
OKZk/RfhyeJqfuTuy0jesPC27fLWXouxv2u7HEm6bac8iFBIJHrAlomH+2XXaYmryZlFppQYU26P
QcpGP3LazvGEeZL/LTc2ZcdvZC7RhsvOM1av1uhfRwb8AvKB/zTVqww4A+y4Rbjs8itet1mBKFv0
PaObv+5NP5TLAfp/VQS0JSJ8ZlynznoH7XYqJJuX/WAkVA4hTf8tV/Pqzt0OjhC+Yht/L1LHjvrv
4TEjlRRhEpDrKpCoGAZ5JQ7Az1X7N4HhlO+mQ2z2SsfbfAXSk8S0JHcBRbJoe441aLPs7dk+jtvw
Iq4EYyF3vpxwG1qxkOIIeTHPGZVVpuB4dI11IwTN0c7x2MmQYHKvUQRV35N8hF7FZNMpUOrwmcLa
ISVFVsZ7t6Q6nI/WBXI6tZ9KUPi8tMu8mS+i8DZSovwZ0yJVDFB+uwlvyDdBciuz6pnmftqGQROf
VpEv9SlHgMAr8ZbiZrW/6AYdWLDCVH6CVhMOHhff7NW6aHK73A==
`protect end_protected
