`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
J4nuplYbQ29eoqdS8+LDs/uD3yDRuXIdH6TC6E4yI3nGxHqRq7Gnlrav0VQFrxl3rfptLG71VSUW
fsWbtWDaLNaqYzF3oNFgAev4ztRBKrCMmi0gwZ+0Nu2mmNt8TuuBxHh3PaItIjfqC8Kb7w4P4j15
QuAfnsDWjGRuuL9/8yTyOonLiinxlSUuEdNnVGheej5GftkMJ/8tumdFp66mjDi1oN9Ay7ywX/hI
AoRlfHsI4HNZAGZPmeWEW4oCK99iLd/irQzrkfN/Rc8+YCR24QgREy0dUVcAVu2UWntkZgEX+9g+
LJ3dmLryxU9f91YwmnKckPkDOafxIjSacf3NCg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="F9wTcE5Oap0hwdE6aAkf73Qb3nUVXX2cHqnrReIQ6TY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3264)
`protect data_block
yFCYaRfEyuYwZqjGinYyiZ3EdsmEIdrtf/CluIt3NiUhhDT10zYfJzBkn819J/kayR3Sr2zRNCHQ
Xy0/WbY+iZ3BDlJCM67nkWung7W33z567ZwIPiY09H7bXJKSV9rKfgYpu9K68QLVazPaO4loTIJ8
JeAJP4PE8t2ZB0z43gpdlCQggyQkwRkGoMPMlvU30PXByxOsKSnWyMITFCVcyn4y8ENMtC3KPfri
cct7WkFjCC+FH8WEW/R4g1imkNBuIXCT+4DiPmwwWbfwiEnJqDjeMVk4Krrop5pxEaATvSGYec2+
RUJvWlUu8K7jKwCQAk9E5YM9dXCp+snGAM3NJLjGuor1EuMpbEa/xGvLdDJbGB2BDTntP39O+SDq
mJCu/zWWXqFb9cQdzyJRhQluuKk3WtbOPcOOvA08CFKTlYuNKIizmy/OgtS2UmL97H4BeLgcUvzZ
D0KGAcuZdmhcprdpS52w4KqBvArWunqRzugN6MZYmbOMbEDNFxWndTF0Qo/D0TzQ31ibhoqAPsxj
Te/TOdxPEPD/b7p9kFCbNqKt+h7IZcQoXVIDke4ZzeQqxx3zqi6SjYjJG13qbL15CWvZ2+0MlmGh
celLeQ/CzQSjHPg8Matm1n68vsQSTBGvgWADxwbSGnrxQY87OO8wqu0y/24cJJvYXdvSstx32zHT
UsieraD8SaIdMrtnfThnewtuBH4hnKW2Eznqgi9X1B9uAzNZowvtoOJK1mXtCak55C0VfIYWbsFT
advGnaI0U54Uc0nj/JcdyzmLKobY6qGQAHn6hdSapB5uLfz8r9XH7ENIWyJsOioJ6zYmobm3sOtz
cjMA4oxcU2p5FlVWJQK7nlXNxfZ9dGRT0Sf0FXjUSwMtYLi3Ryx1kGLcLRpQPFWwwJflPSbiTF/e
jT1aq9XjXwUZoV4nwNDRc6cLdPM7PbA1LpMWoFmFj+TGbfywvqNPU4kpHour6+Kxel18KIjxe2P6
7tl2NFzAgmJ+CSI2Gz/sv0azy3VuGoEBUS+QP/A6KrhDewkxWbRyjuIAHXwgDzewU+MqH6mEX3hR
HtlglxjoPglDO7ozerKVaKb+RYkUIHCLSg3r3aoFzdap05QTz3VdYGWPfcLyuhmMByUtPUJ7W10Y
qlTY+Cwq3okFmSfhf2tO9ysOlut36Yp7e+94P8vMrFcun62fqpYLbxvoA3PPbU3GWPRmmca6gtPU
3JG1xmgww8W8KU3cMbFihidGfX/G1Bb6S47CwgpPumdOV5lViIAFMFMWw8o2ZC4sG7/l/6znd/Kd
LT9T1bPc0bsFvFlYBDQUvq2ThKqpQfM2NOW2KTbAN+9BPSM6eVjecjYoYZnLzHYNguJO3EVTWbXe
va4c5XnsVHKXBEgTLf9rVI0/P+1B98DWA5edhm4CPsQ95t+sp/RqVr3zlj7PXBVArMQ71NLlS++h
TIEOY5RHQ+t2bXL4tEqWYLOn9PPOubaJqVRV8E2YdX1hl30oQCZ8ZDphHPhRCuPcqtjLyVV3poSC
eoQOnXoRtTpxjzIBmSZfjbq8teogQQ2QrRSmcQr89LWVpUrV1fkrXRnI5SzLW8Q0JWbIevDExebl
lDcirYy4AO5qoMY+OLWBaDZCQ13aoeSk+XMKySQGaZjO/tUxeL/oCXfcQBNdLIn0jH2/v0WJvryx
+YwFfKt3Op/k16uXkrtcAnhEm/tG3x4KJo8DcpNcF2rLSh9rS1nlWW6iika9eAgRBU/ekTp2a/9K
RLQ+tEHLNcGcxmt8u1gqGBtEzZtghv40hZ/TydCz7/+At9ks095oS9M2nqNvCg7/brVfXLZEHJl+
At+giO8PKtZUWeAoj6t2Sf9aUb0xR5U7d1aCEAyg6SacbMxDd0FLj8LKTLGjRQRaHSefzZqUUbnb
3lFIOQeZA0D72uBxeRmD3wQIvQZ0tiC/0A3Ay2s7LEv6WA0zgcuXXeziYbmfU8HXSJHm1YrUVp/B
E4FhNoCU/o3k9CyAnmPaa6j2gmsUfMnvUTjV90IMGzQa7mFrkXJc1Zy1ZgKaHON2umkLF8qk3YqX
Zary3tRc6DOeEU0eC1I8tJHJ/cQ2DtV7jbiojwvhMPO0JhVr35q7At32XG3yPysi4A+oNhYtXkf8
ygQKatl2FpPi0Fj5V1fe6z4Hbvttrnrd9J/3IL90pxKPQPsgmFNptfHMmzSFe3TgmwtQRi4oS52p
vMCuo1GIb315STvK8H25SyEWquOu/F9Rod2vmbZU0p+rro5Sx9tzehRtXO2ZNLYkpf0LcRs02weE
8Ikxpyeum+7VUT1LuCxwL/ZDM3oE69ZrvCCaNYeVUI0izFUY6Y8oXEBemEqaiPqTlZA6JEzbYA6k
CC9aFM5XtXrt1/VYJP1GqAsVA4O7GJepvsuIvOBpl1wbI1RFdJfAXqa5Qw4ZEXVZMAgtGkPFqJ5T
SI+ucxh1b1299h0TUSH/vCA0yjXLekoGlZTgln797uOnMOMdVsJSERHMtzWJSyiya/NwKd0+goy/
E17KBcly/+XC4p4doTd5dHbo8xcFW3xtJPouDbhNiNTOmAu+4T8eUFU/iVbsbdctgOtxCLjMInc0
2gLDCrUTU1ay+TtxPbHtDJZvUtWGg56eXeXAPc9ZszccnwccnZQ9zFSg7DCJoP06P0uNqwvrsFis
dNtySrDDEGce1jPUiAyeJRaGvqJK9U1fLw+iX7fxwwSJLEE4CJA4zQdrflbNwjCLfkI68vSIklkW
MiSH6IJ23y/qAkMpuLhNmRyeml/8L56UAsQuGJnL3AFDWHhOvrFDH4/bzCc/qbl15GNgB9tZQG7/
0A22FGH/yAtaQl95rdOu/R/gXZKddTtN93VXTqgjpDgEQbIC+b6rwU2aYiXBXIA/Dn/kJURmgPHZ
T4HkkeSVuSfjDfU9xicl2N0f84og2hJ8z5ggwI1bkun/KUqGxqGzTBZgy+Q2zsbAgApiSBjCK0oN
LVUlGqQY5UTjmkQMJux1tvg+fx/CPCKDA2GGkp/tWGB3nWnzJBIMmAlrCkU8oVgr7vHHAPz5GlmO
rbL3Nmx660jM1i1EVBReu5g/eLPA9yxf/ANHhk3T8btcZLwUMLrCIJS833iPlZpHWRDBMgEg2y7V
wOaQ1AuS1Iy9Wv5pSNFjxvCOkIU/3OVpjjBKd7FhvkwWmR+vYDNWNKuzhoMSZZV1PqHrKF58xr9L
WadNfnYUTxW5Ke/ACPzETpSyNi178UKgczm/QFlC940zxl75rCZ3d7XE4Bs4ZmkVPB2Asqw4U8OR
BJKJ9g2hBdc2v81TLELC64dZxIFoy1NIDrKu0mvocYCrDev8ZALW+Eql+Pnwju4CozgAK6yL09yo
2fUwvbWtBmeKvfVz0Ttr4wa+dZPR/L8g/r7F24iSzYL5itjZlZGTWeOjx7cyuvBim6+V33JwdE4B
6FfZdJI8Np1ojySqlydfPfd83qnMLfVsYrhOSIDu2RJmgN85KzLHAuQbcDxzQJD80DfCrmM9POPO
xsx+hsKq4n0B1pITF/MRvRMl+qGbgCfr4+cPMDZfj3ZK+DlXA5fMxMYU61TtAFnShSS1oKU0FPBg
c2EDhWGmt0Hquk47kTdbH8AmnhtwwyU+vXxycuNw+/a/7z2eFwLYNg+5dfY1Soz2ANPeVTpYDTiE
LY/S2UOM+rWerSrFuhpJsk0gMr4KAj3gpVAsBkC9r1WOE/bs80ZBWo2XtpFNFfFD+k2K6obrjqgE
vQAdpq3AC9cuAbvjiPN7bS8QYR7tzsUtCAXn2yT7QZfLl+HdsWORRsm7hCLubGbS+hVY+j0CPU61
P2EU6mYLHlzFC4MNmZAkBG10ZZvAkSunrmZhP9OmQ07cnGJ5NZhIiM56GMbwsgI/U4KIUWNh5iS0
OVWoWgFFBiJ5HcBO1KASoyfUzwljZ4yEIPN+JUaEqoIVxZW+Ih6r+myMpQ5BLWpWH9oj7LXDa/lw
stM+alRg3jBBc1TnAjjH4NzalR6taJ3bb+KwQHCLW78paDjOo/89LI/vpdC36BsGFuzO+UrzjydI
lUB1WKAqDHPwM1j/ugijokcmYItEp6fKaBrCSoyjoYLvJI11uxuiVw+seY7HROdsLcuS7kYnItrO
V9ZrKsgi1nZ+bFgJ9m8C+HKg9q5fag5+JUNUcdSK0TxdYNy/G97u8GfthgwN0hOtNOwaQ8AfbJCI
Gqf2JjQnLWjBE+ijgDlhdDKtPuGedoACe9mnbgCQEQKVEVe6TqQ11aexQpx6uO9jESvONkpzcy/Z
Qb//BQdDB/DH3gJka6x0pmMyGlEMdZNRDnp5rY2rK5/OL3LHsTYCWFqwQiuimhgXY+V+yNp4F72N
1gW8Lzr/aIJLFYpjoy7v
`protect end_protected
