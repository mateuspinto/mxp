`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16400)
`protect data_block
0USWSUGxovGsyBJteYpEoXBaIiwGMT+f2O0x5VEiYZu5TNO4CM9xNdaiIYAMdTMOuUuqUu7879kW
cA0ZZYSAsiTly40qXi6zFfDJh3QVD0872k36wdSV4h2WtGYhonYMBq0B6lnA24BHx9bixtna+tvY
VJtk6psk30Rh6EwHw5k0xvsxTUIMWmMjOw/XVKU29R0268DZxHVwL4ahsjtm/g23iME2ufDiQIxG
W0TVIQskWLLjULLB1lIDxgEznSpsqyt3dhDsEEDg/5ydLVnAaqPgP/b4/NgYuNGVHzzr9cy+K4HJ
Lkss3TjsMlIlGBA07elcfgYTE5+BwgMVaXQiMzSHa5TuIj24gHA09LHKg6ehju6x8NRm9TKrIvRt
ogoFUs59fqJmBfVKmPfDNN2lPmWYcELqJSslPBUhL/+UPRn7A2Uxs+OzNEKIVNUOfoOCPyujbIek
HG0GujzYYPAhZGZX4txO4PvC49YWzzeo+i6I6i56DXPRjzgn+HXEjG8MkcCIZinBwbfajqLcJ2KN
pji91ESDTi3n5qvqsbMFoH9vjeHomlmesSOFM2hTDTCfIKHDaHIhW36K54eenonAK7tja3+nCVsr
0NBoJHxycV4KwdIpBUVvqLcvG2lmInGcUzF6sK4uti43CL8g2CMAx9VI75ZEyHXUXsdpX01sdg5R
IttcNT7Ab07qtEQIPGN4jqjR3FPYtzsEKixgmto367Tztkmgk9f0foQWnsntTrPEkJT3uwJeT/Pf
a3d+YHTk/Ttt+T/gwcKGAWvrYE9KbOZNZmOoRfXX9SojK9eNzfCriYXckWk5JagIQHF3YeUqqvDa
KZdzRNqHhRTJy0JMspYahB+eWaEq2Tk4i7RdiHL7f5sdMJMAm/SYqRJ9RKrho1AFPZRADdWj6ayz
4xYiyipL1MZ2hKodytT1G+Ruy8mAw/EqiitdUijSoHieX018/tiv0b/Jn1NSXHfbKuAyAk5LOOZc
/c/2h/i2UjV7HN2ITomf98uEYuz9SeN9dIdxzlNruJh6vQkVu8gFk4T8We0IGsB9o34xq5WytBBX
mEJmtMkW6OHJpSFS2mNq3xZhrjPzrdcLpTiGY/d8x4F3sNhXZAkmnGaQ5aCPCx/wG3o58ZX3KUAl
bvN46sZYp0u6JovczoDoWt0/J82DHqaB+68XIJBDGQehSl3HtH+mrdtFfcv5aO/WfGFA22nic8vD
8nQBuV486cZl1V7fonrgFomUmOVA1HZFHXpxuiLOScluQBYBzqOlKWlKOr96Y+oXU3Q6W8Yuumi4
16TRS1DsH28eoy5wfZ6hsv2G3X8J9hf7BHC38ocvGhHrZrj6uq8oFl27UjZ/u59D0ZY8yxqVEDjx
Efyg8NZRm9i4eswWtMP08WpNN5fQR0y/mDxntphKd03JnkeAztbAYLkXdi+nddeTlZv3xJdIgQUO
dvhBxl4Ag+8p0es+Tcow1+qJkkO2WdEVpvTVFi615ha+ODGtbbQwTe/Pu48sG4H4YCKChwJ8062U
fXpl/Id9+yDhkCT9EB+ErMmmXju43muOd3Y5K8nt5JyYdKhCy8o1CVLNJNmmwOkkaMPApn3gikOP
J+TWD2At4aD0X0kyBwxOKCLl9NWhJrqnWFkc8KmwC3cI64+aCuEpSNyerFcnNxUvcyHxRNEleo/s
YDctVf1yTsBhh8s08UtkQw87MbNDuqfJI5yJNYFGk6YBdwQMRiNky+tKZqfva3RK+D61moKPBtR4
HSFCajfACEVu8Hf2d1NctzfTHuZpaC5bBWOqPcevRodlAchrE3NJ41G4yYbkx65xWsgBYmFtfMnb
srps46sSARa0XPVHaUYsXV53vOcegK8IHrMm9m5k3UarLvILJ4ogveb6RjiA+/DxESCi48ifIQYq
vfXrqJ2IzxoxvP0oNTw0y8Dct1nrPN+P9+v8FU1h17QEiTgyX68Qt3T6VkRtNXTGTkHQ0kJR3UMD
/dA1KSndzWhtdh6JjR4iRM4mCE54iKgviHohBpVG3iMbGujZwlgYpQcYhmVHxS9v10BMvw25EX/2
b/96Df2+1PicjTb++XrsbUBJrsEsz9dR31WwOGyn92U9wAVFcFIC1l5psMg6BnIPjKRY/jYQhq/F
dL3ZJwArS8Yw64nPvOhtJGwK5RhFT/eNodbbk7f7Z+6NYaCBqGLVqnmlzcaiQtrxhNNWJW1bgYqD
C+o1aghnVowqP/Fbw5Np2oIw5OpHY0+BucNQByfyniEdS4AMpHS1QHAhcJopTavw1zExkU+esWDe
uyU4IV2/f6LO5r6Ihz1eycNiMffoGVxzeIc9XMdKzJyrUOfvoe3sV3TdK3EPdZ1IpPOJOF9NLw93
mkAtwmylXqs+HaxKNCpz3IIw4oBeLSe2G3dEvuKVGNGkckr1Ly9ZNsLS+9c1neRtWNH94JT8+r0w
V3w0ot80+BIrZ3UBwPSoPvVcBqJYTIDErHn6oUN5L3EujwwXg695Js5odGQFwekIEPiK/Rd/Spfp
XyTFDRglDfq7+/F+SDBw6aY98pagMbB3qKZQ/yesFnGR3fbqWQu4+0iVhMXJ4vtWlbN0eR2yNw4M
c09lRNN/kYKq6qAsuCZbB7ZTnE5hqPF6kIglVbQYj1ZFB6T0dewIDtUdgg14OWd/d9whE11kDLH/
TYpNzU2vZZJm78xAzyKiuYou3p+V3sgEUZ7q7GY9Lz57b+yhjxQaT4R308wGL3DwUnveskDCKkM8
jOvA/gXutvzoelIwzdEJ6WGXOLnvryyAvJt2hYCwLmwt0oUQO/WS+9titR2GgAJRc8K99OOi/EdA
9WVYWY5VWqIipvyt+LSaQdV7P5kqIB7ng/Cxjorl5tBfjmvnqgaO3hJrlbAEa15UM+7fajBtFY/j
PyYs19Sok1G/Mcz58W+O2CBccjocRbjcreV45tzsxcvN33F31RBnST++Smi9U9dWDl0uxhhsgwIN
+ZD2VxsZXINovTaC82R0s7AqIoSrgbPb/mfqd0wxf9+XTwH6sl+TpEKz+r/2ZBhIHEklefgg+l84
MU4g9q55Jj2jvoWOTPx42IvI58Srfh5mM8IQPTMrnEm2RrVXcU6zxubtbAP4fIFNZh1snEJAsk7a
icHOTWSxQ0CZUhJd2Bkvoj/Ll82U2Nm+lS7JM+DZteZNddidTZkgdepoH8eJSHXyYiJzN6UosMAX
oaX5fVF0RJ4jyvZtSnj9nvGudjDx1l6nwIgqpRDeClYuUcBkYtv21E5S3vsDahmCjWL2xSa5dv/i
9tDAaLZLA72QSr4bsGxBk0deIfhy7myAdob23HH7c43dLhrtZ7rI2MvD1rokU8KjJ7FJ594ocx8y
zeUcD+tkFt2KvEkle0tQi+KtD7VEy27qeqhfHz1iO7feosiBkXSeZRR0idsBP09DK+pq4WsgaOi5
yvViFGjO2HmzezGDhZ1MkjfBB1xpSF0e+lU17/guSXMtUUY1oZBkVCuljcZK0e4xApD0l7rKV4ut
mfFSsuML5aiS6X1kxLwljJlGTe3WJaek1YPALxsxq3BFqmBthfkthZ/dMqf4PSPlwv4PZVY5eUkt
FlU8ASIZ8o4AVzbLdtlmbQXEBbY6btWrJEJOv0zD+Brn+fsscHj9jjboQqRvFV1sw/dHt4v8tdam
gBteJez7JLUrcCfzjv4C7xL54KX3VfysrsIE3HLMpAohdbkl6TQ5zy0j16RZTVVvJBsfLGrODhB9
r5Jc7qa8MjwiB/Ucwmr8/IzaLPDosT2QMT40MiI7x+yI//N2TEx+fTyPSb7cYQe2epEn89/Io+vf
W93k2OAijSWh9kF0kcCFHBDRh33voUjc3Nh87ChJE8Sjn5uJiVdkkvr3Wg7GtT77sHnu0gExk6sK
ugau3XuyuTECUd/5bQ9qmo469QOjkJtO4SglVlglGAxssX8NXz1C1o4m+sstQnlb5VO+U8eQ2bT0
Bt9mpFdSh2UMteINrECYKwKg8dV2KmmfDs+/ff2L6i4uLUbHYqTFS5M/sstTXuX2q22PNDyXGHCy
ztqQbS1DNNG78zCZ8CSQ4016DddZJhuKl+FAzLOQmDL9qqHqs5276s3IEllzp8IaeECyHrG7sYC+
W8WDw/EDpjcf74M34025xFydQwsQ9mKXBt1UIT5oDXSV/QR/NmR067OZMEl5oaRNOYeTxvQkH6+S
5IhwnO67szWl2fW1FQAMMHi2VtMTB9f7hrlTjmN+kRPRcN4sFDsD4TauCiO5tqfUBk05wefWT89J
xO2hs/hzr53btjgU/B+SOm0KbeCBNsetHKOpHTHL2gM4ZpYx/MTzhJaH0DgSZ93/UBVb2n1iJez5
IQ2KUb6mWphq/HSUnoX9EH91mNFrEGUqAKrJOET+iJT9rkN5k+mwYJWjN6suAGzVwTxYJV831yAH
HBUsa/5muhmmJcawf7dOrVNqT1FA0uYOBhREh1RoC1qh5Pk0zaE3rtaXmdeUUr56EwDKZRCcgdh0
Iglgsr2eY+RccbLUBb/3fltgT1kZJM1UMnZ4GZHAJ9j8dizLWQ5PIQmtsLUxrapFoV4O2wIjfu0r
R9VfLu7l0mcyvtikzOXN1Mrmdk9CaRr4Lj8NkPBuu6jrwMm+3JqdiQl8tgAEXT6fjml1/KIMMWCD
RDppvD25Kj3cFmwau954CPOVvMypY6FdKM/2PrnAhqIOX/GH/9pANycLsmLwt44u1MbgPtHhm6xd
nRcIlHVmyXEXE8NCyTSYtOpNp8nemINIAxhlGNdgbS1Wp+laim33umdO+OQlIgGhPOvcuik30lEv
3FCnEPny50BSAdPMVH2CrBgxQ5H0NMI91HBOGHDqpVGQNaCVOg7VJnqEMPItXr9b3my0uaLoZalv
6PCGHLHeQbe9p0Gz5osS/bXJzbAeFyGMReE9jBZx9krmZOECvz9XhyhVUfeu0wMckS4703t0IiIh
S1c+l9yizh94D4ku53XwuGBtmZAjbhrYI34JKGmNkowx6Vhwig86jNs6EFQ9AwKrWusNk/HdfG2r
U1nfhOG58NLGDm4ezzXswkh9E+Wf8Sv6RfzB7otBhtJ9MO1yAQ8WIb+K8N6wf2NUFJbI3sfrHQ3n
JA+Hw5rTvlWGrESlWzFZ/wtcBgvvBvrSmR2h4/koWaiZaYYdkipKq45VorD0KVOEL+G5kbP5Fi4j
6nDMcG9V3Qpi/ZpPda+4QoBsYHK6VnmjGrgFF7MbcTkZ7EUcq5XKC+b5vwDjIPJWBaNYYkt6OKgN
yfs1oKJ95xtXc9HXWqQ6fH0BJqdvZuz843V06tBfTr/p+tf7SqrtE64LNprrkm9v7hsKHW3DzpRd
9WbNWlxfnGrND9Jr/aooZjMUDo6JcM+CLmSwS4JvwZL2fCKzaMxtGwIPFOXMIHKC2Bj1r6uajAhT
1YO+ua4ry/hJTk8tqDRcV5jhKHG9VCWmJVWZ5U5HOxp+uukuGzMv5KMUVKl78DCZ/cr8370HGZyK
hxy+aeqkUHLNYti0gMWSYwHT5rwyVGzNUpETqm2B7gPToFVdoUTcUpZcdyl9WOeKCRd5TT1NG2FA
A7/ibw7qpbUFIZNO0ta4v7QuXJVPpCG0V/K0eWof+Iqn4439YoGnnSz31k5BNlxpFAdCIR/zLKRt
vMKxVOZEwJkuSF6HJtQYb2mGmp5BtZahmWoi0EiqXRV/XIXoE8xWGzoUmTjycIR9Ziq6JvzooTKa
Hh1FGbGynOHGMH7Jf5ttSbsa3y+spBCdM7QSnDI0rFFuXrr2xlFqbjHzT2MyZ4GUkGs6o67Rhb+F
E+1UhhHIA3IzleTlUZ/mGbiPTBT1urP1Wd7ahtr79ivKKlOz3uPphjQS/bOJm8tnSqw9m/GpaLcJ
SJgVfCY4joK2/NwwIsNMueUKltXBqd4X8qb+atnZkV9An2p0vJldbsseUvtmNno1BUkxTltQWUQm
VQJdzhd1CMArXw6mAGIpY8s5E3TXO9TMYlS6QsN+yihZk0FfYk0A8Hewp6MTik1S5XbzR7dYwpKY
ITwKQokSQCGspL/bMYE90MrooiFoi2pRo/9Cw1l16VzIpLDHIEH5ArGOpZ+ryaEOoZCtSk4O0w9s
CBPiNoRXyI0+fyQepe0npUElFWQWbOba28W/hYbHfZ+LEsOYRPxP6pNCgkSyEHySBqETSNu3B9d4
YoU6juHzC4belorE0mc8dB4MXqOBXYBTjxV8GdLYDnAAJsdBn3st62zbtUQIHbicT4jEyx5yT/oy
qJ0m9/JVfSA2jDFMDQ4BvETeSsHZWR+Df1rWz34ebNCpDKN8qPWgJCv+5OMtx7OZStap62j2fWfg
s9A2SHWdfA5Pyh+PJ9HPRKCOgv08kqbRbsOB3aM8LxXQBCRh+bhOw08pNp8o9yiLUPz1VF09w+3B
aoykQ5Ox5fmsTLciFsa/pAO2MkqlBKooUOwMmIVqDagdQfvepozi2Cm1deWA1BiMdiT+lHr0O5v7
ppe+WRc4Wpv7RNYaBOsiPOm1asrWDHIb0CWLOshBgckwr8oXSzVLTpD3OIlt19s13Nny1WDKqGhh
GACij/peauC8mrYXM+Em919z6ERwvn7fw8HBR4ekFIYFajHVJ9VoFt2qY8kJFi1kRxcsIlcZAom0
P1O2zsFXm2c6HH5lqYy50b5xrdO3fBQGICg7CjvOI+Ob2kL42U3skGWvuJiHdWXCu0F8UVkIkcAP
VTSFgszcLcuLYk1lvqhjzC0GDchxO56las8kpXPOB1LSTVhjtXZGoXDLkM/vLpPqCJyP2dR6g/4v
Vnc9jc4fDi+Ej60a+V5RtIs+IugW5GTp0JMOImTl8I47gi07dHywlsgtsjx4uvSdK3CzJT+UdQ+Q
vFhaXklTgAYlqa+4uW/+dBLZQitQmGwtv3BRBG1N3VSNPVeZwl0miF0SSZ2nSVLYa9tYMRZi+0/y
hVd1KSb40xxx3vYmvEE08etlUBY20pMabq1c8K6YAl4tQCByHiDyGqnPyroje0VqTBZ4b8iFh0xL
2+N8YmSLvh1/DcTE4B9EP8R/q3ZmBTkAw50VfhuKtxnesa8U0P4U9VAFJDabYWq8tOerhZOVoexA
Tv4o7VO+KSEDMBki7VPCEC93S73jjPescmTNIVpQ2Y+lHh+ytnT08qt0eFWqVTNoXTwQaGTxp/ik
IvDyd3qRCsyB6teQG94WCzn7sMLcKdBLe5JUq8lPCDMFEWxl7dp6aRO/slwCUtm/YOoupxgFEcVe
Q3t/iiEm48nDSB9r3ZHEDg6NMcDwfXVKcMcmN0nBwIHbX7m5N8OeiaV1Zp8whK3HeGcAPmMHquig
VYZvyFbMU7xTbwbTl9cmpb/HRr/xE6PCfaA/Ck/eCexgMfWPQK9Qd0MVePddphWDtMNf6QQTyj3c
T4cQvEoMyWmoPZzGumosslqpyCC2dI/9EKo2+QlwdgOBZAAPt7g9FF9eZm5CnNeXXfYAyAzzcBJC
ZmkSCN8E1Fdi24VDg7+SqKrHorTp5O0rs1hxiHj0eIjTJ5ckY7t2VoglB17+CsIV8/p42/fiWeE4
KQ6r1QBmuZKGFdeiGxUQop+6zEUxZNqzHNyJ9w0uuy0MijG04Qtuhq1+Iy0hyORUyYsKSSIHzxbf
u/48CJwgLrmeecnf/BenWk8bH/7XE2tGVayNqWNmYAixBVB4yXtRX+jBUi38uuKII0byCj0MUILA
Xo+rYScUx8MNz6N/xXbAOyJd3SvB7JV5cezadSjSHFLNwEJbmJHvmg+FeMZqsmbIm/mkLKv2UHWk
nIrR4Z289ZLYRGHychzdN/usPnKIbMIBgFz3xYx+AZkcUbXhEhVcc/Fa21fggsu4SezzikYSS0Ey
0QZ/wAEwMf6vNOT5icLHiqaRzb/dQIYBF5s8F4UR/HkmQpZXteYuLhdZhLVYeq3hdcsu8YJztg6Y
sNzwMThqu3d+yNyDkBcxT3+yJpReElRZ2pvdqa12QcKG1PUtgC21hMOSxl0cfEoN8yQrW8wx7s4Q
AOXHcdwgYLyLpnCF96GrjHWc+s/qTryBnOe3C3CbMFpwVza3ojb2FGG90KNsOATzNjasByB76GyF
d1dy/BAZ6UB7KsZkEop4c5xpCTaCO007q9Oip7k6dF9s23Qk+6Srw3N5iUUPj2Kv0Uh7/jOTZt7H
QE6hOri40FQuLXiNyNdY3P36UgfVKMmFV0n+pnFxymtRT+rwIPUu97eh9AhJM477PnrR0l2gR2Iy
GFezvMu37r/kFwmMtoCjDJ00b+6ItmWM/Oa/Acq5zIEwPIsESJsX3BYpO2aWzwjmMHGdWjam7gNd
nuJBfVDuB3ayme9XhxiwZv6Zsb7WgFQ2i8CkVQo5QgDLkwgJP1XDAlLQif4EvcZqU3ZucUB5WPTo
ik4K0LKB1dPTLFMgPN7Q4A/UppHtG+bvVXBi6Zx4Gt3clb9HJe4b4HC2BbD0/ocp3ijjS7xrKe+e
AL+tZAP/bNd0NxUFSryHV+oAw/3GPWxuAgxpHMNB0PgyYqCQeGiq8d4GTago+zlFxmZYqfIWBArs
wrvgmbDaPorq1shj23m5gDaOjeKuAUXwapPPmtM/uCnkPPgviMwwKeRPPhr8IJotvyzshwmnMr8j
Dm8FP2pv328C7tqSw82ltcWYB8vqtFPw7Y6y05Z8YBuJPsNlfnJ47tHn5ycQwPEWxA1zGqpEVTvL
8K2clJo73xWZelUqcmv3Lxxma/6PCV1pDjn0vwFiGeMRl038zs2R2f35BQiZJloPmb5SVpqPHSuh
ghmaGICE5sxOaeQ7lh2jxH8V8KsZy7km4ovHwdM1GPgO5+yVaB9DO2eJRrahe+pTy5G1aALHg6LI
7IoUSwfWeycdqP6pUc7HvsTmx5VNXLsrt8AWQiY0VZZrtf0aZKGEzXXdzjdOmXgufk1g7A4YZ/+/
J1depFaQiqbM1gcki9Xn0jnjndn5hoP+FL/8dOy1oH6XwkrzXc8DfpFcQeK6cSF2DN3fg3psCTiC
TUlB8RwQvqQLtMtukcEZDI/VNeoS9QMMFAPnalDraDh3b1SCIeiDAzU63j8k8zMAEWVSIBnNyVFk
krzcRnaQTmWLPkHywbNHpC6Ou3WO/vNVoHd+U5gRJ7cZH/oaP85mjhsBzDkh21DT/PiZHm96j/PL
IcR99vwy3nEd64bDTwXjJDqHNOKTmbtsF6Yxlyeag+89rb4Wg07XixOttMLYxvhqf0M4nM/FmIf8
zibRahUChXv5AGG4R5Q7RW5akHZKi3SCbQMrdVfVwBKkUpk2Thg3vpZPg2H8663o2h69pNGazRyf
OsQX0I8tRx1eS/dMDBQ4p5aM0WTn/ymHUSCoEj7vY20s0CnXSemKZs0ie9KhFcow6PVWR4fZ7DiN
/GOFNe00zB4sTXciWES4Yr0siu3kuG44mPjTNJyINrnJfNVDu0iRjTuXWEkAA01vlzRsBQLZ1bZi
Ck144wT2ZsLGdicVxJj+ErrIqXfHl+/FLkLsE6cODOTqqLMWW1Fs49L3Q+5GzvVc1um4N1G9tPTn
HrDNDd2P3JJk7IfihgKndl0iBczplklqt6p/S+yf3s/cylr/4ZWKoBthPlKwLodsyUwP4pD5fQiv
s8Gv+0NToCdryhv7Rg6VcQREEpBOEf7sbbO02BVJe+MpEX1yOLT8mJdDuufDLC4wHFQCR8JkQntc
91cvL2z3i09O18uyzg1UII+k/nsLw8UQuiul2U+XG8Ne+EUvHWklaicb42IhPSTwAO8ksDuUPgAn
AN53h2C5MLChqquVJyFkxBCcLyCnY/J5dC5pWv3TrRHkRwNndR+qNvO2YqZEJp9Bb60NqrLNdjsG
EcgKbD/2lN1kg7jR9RFkPahoN64qE6aiteF1gZ58KXIbTtvRYcOuGb6V1Igwhv+F3s24omCkpfk7
5JP2bUO5s6bAJ1ymtjQInIMBDYFJHxmAWDQYMnSymeZks5w4n+QGwiteNI+1DRdhVO+/Z5OGDi7k
SmkazlHcrDQOUWJAQVcvvvq1X5IySoZECe66A86rJYWwC72oUQDslqC0lfXXEdjfFNPWta89wCh+
/vacAR6wxJffCbJ38qjNLm3Yftj2kPdgYNsfiw/VfNH232x0Y0ZV+G3j7ePwV6aY/9hunk+uPgwM
QFRmv4vLZUUGnqFEUw82p5qfdkGi5drxsQlprEUCgghT/PHsgoMfuGUSBxufv3u2w7QixHRjnzLf
0jRF5bqmkVCw50QGS0zA8be+C2/Wv1PvbNWwbU7Xs5x/u+yL7JPmhoyQj0gPE/3xeUqE0+zG3iww
lcpeHEi7jQCXFwUudFz2KsQN6hcvtJyBGeE8mJeyGKcFZDmPe1jnOVnumz1uun1vzhXrQp/Czmnz
JFW92A6RAOXl4A8Vci6eCzWkwDf3v5VU4d1zbXadG3fVEBwhQLladU4ZwZbtKNXjLx9/TqP295Hc
BMVvudoqEXhQh8WRABCrC3s4HklQkXjMnS262Ic0gEDcxqfWo5zy+81fy1bibgw/9CRFWRiKV05g
Z9/03M0SBBLkiBXXHQC9zlSoGKlQ0jZx6uYXmc5ajvtj/s1svuSn3imC4+xucIVZmAjmh/yF78pu
lMuZnMizREYEzVpK5WFee3JVS6YuLyCKrxZNgkiYF2t8UiklNkTQFzl9TmzcjzZGkFeymShfJ4RB
67SJNx3zBTY5mEYx/R5IbqVjSN3q4gfMdW3nPiYvW44Vq5XoyDUB4VOuetsEYgg403GXuuORjeey
g/a8bIX6lWfDsBHRRS4UG30wzoUS3wtx1PzfKaldsGlBbfMAEiaF/Detnw/IlnGTbvqysUu/TSBx
2RGHwphn/gdfn01htzSCgJI8MwlbuweYO5Wjke/AWKexBY6rVX1elkdhoBHF2lcfIg9WtmR/G2FB
t7aQAMqF7byvzxnteuTE4TAeqWwNKpWsOn+Kl7E8SbH2FJJ/B6nQizdmHHCIvk8JtsFKUSTpPzfX
nXKCurHig855l85GDD+ewHFmxVFsGqWVqIkv/sgYsCascSGgGsczfjR1OJ1C2eChEPuHGty9IFej
olLvh0sK011d/DQZQGlVoOyA7gy92VfRqCw6cCjV/C7iu9eNAvWAJIK2Ue9L71uJP5vO1v1r3wf/
aRtWa2YyKa95yRiG8tuDgreROGQ+04JmKggIxIKlIKFYg+m4fgw5TA0Bu1Q2+54DRJ2i6mIxlL5p
deLCSmjCq1+e/SGM2nRv5WsEe79ctTJbCvZqAD7jj/QX7cutOP6H35BOkNKRb0DvBc+aOgNFe+1o
MqP6Gil8m6C180cPEqTHTE3tB7cXfAbPZe1x7FEyUuYkmaa0dMoTDewZl1X+v5gVAA1GNhp2I/ag
2Sqk7j8OTaNF/yrrlz/gvDRZDLooKBDb2It5UqEf3DPdtH2J7z088DzJF379rMOzHGMcP7VhbOx/
5OXaLZhdNP03JupydZhGAlm3LezOFmviBd0cDfwk4la0Q69HSge5Zst/PO4ZxX5by70UzB5C7/fD
SJAPJBJ4FXsiK2gnJ5YwsEbzy0mRZJtjFc9+TDyQ+DUcNE5BEjvqZnzNSE9zuEAdh6Ewn4meyPJi
lKYOsNLxlKbfL/GGrezCOWYVJA9XPR2f+atpDa229z7VQCP1APcCBQEpkewxxceC0K/W44VZPvrs
p3JDzWUj3AOkzxyYr7jUqo9UAZOisM8JvMHSaYu0b+fl0xtIVK8Hy/JI+v8hwj2Xp0UGgqn3+3Iw
dUCdFJ+iGF3N9dUYIsuTX33UkhEAOh4LnJWXatWcbMtrPYRVvzEqLDGb8woEx6VMLztXxbfJr42n
SPjwUZY+6qkdIVDXV6gGpZrV+pPfbSQ5TiC8kt1HyTxwZV4wu+CHwfBBX9qxGCF7Cix3TqFjA1ir
y+qJ1N3NM8+gMWdiM2JL3+0kraKVoYNW5DNzVCZwDb8boMskYF42fsNzkL6GZN/Sj5GyCbUGFEv8
ck++bVIbT+MjAV0OJwd/+qQqmZKCf140T3jQAoWDE7/4cODM2ZMEgCB/kxiNXqaNnblCZW3EisJ6
XBFxCfGk10ZW56jcdU1zQz9+REccr3X8wvA1kSADT+Ks2IeBuW8NVGKTmOwKsvdi3I+jlPBnWO0C
vHM4gsqkM75xz2hlulNbuXXUJxcUFQH3+K/8QH99WOZvDTM3V2BbhQIvT6sxMhwUEzRMlIvLARcr
JJweCQo5/ByTeSPPXGyuDRPmG7zatfVJ/MLrJ1j+8wbeHbmukBer+6VW6EUVsDFoqRd7qd/XnawM
VaS3RxowI0/dzwNuSWU0MsfYVQS7Wbp2jSCR71lhdg+b/a2GeofSbFDy8hSKYm4Ek5DSB4ImfsyN
J6/P/r/3fUMFLh54J/3wolrFyCaEYCD9qisHIEFyuoSid1Up0BuwGYGMmT9Kju7+bNl7is/7uE4b
8eRd3OcsboUiwoEfgd5twuLT2SfTQe3ziWxl8ovpNYezWV7pzl/LEvZRAH55kZNOeZM6zia4o7y0
yQajI+6Ade8IiVgT7jqlOY3B501mlP5vPrg+hkpw8M8Dj8LXj+GSYa9wRFo7FgTjARCm8AlHPAMO
Tjm/6IBCLU0h9ZQfZG28AyM/eIPYWNSsgoA7ZM9c/QGDCvGotuO7hDkZTgWlUhNnsJue1r8Detw9
idKjtQMwM9L7qeV9PZC1/S8aZ9nR2CSHo8NAwFMwDtlA+LD+97M2uUVoNi23jvUdrFUqDESLKDp3
D63WD1SCsm9bPikCFlD3xg9soLE650R4O0ICnJfZ4YxOul4xrxykQyydxT6wIPl9o9h+x4AT2Srn
8dp8vGt1OA7l0Iny6VuD++Uv/u4fBKVWVVi7nBHJ9GRifzqkQPUvWt+0dTmlExQAasLcqbrZOOr6
vgvMMmnBjUu9tV/1/QFbHvM6U93vnx9wxybl9z9zjt8duJ+NH3GK1XD9OSfjlAnhB8/92zIhKqt4
EIdjF4o7nuyDkWqjocnym2fLNMOQYK/iBzF9QsEAFP+8iR77lUjZSB6dcWnaJm4aB33L0j+Re7oH
FRYyKJqHcAqyGF5dz36xEwSoC1/xemZXGRlEMy6/mAPySIRaVDQf6oJUOQPl0Z/234DgQ13iovIf
SnjLnjRNH4vd6Z6fKqtmhwHpWIL+dhmWmzbEi1l/9yyzoBNLo3gUx5d6fRTvEknsObfNjZDq+cDK
oYtMq10fPsLS/RQkFTOj6PRw8ySZFsnteBS+2ONznfKK0991N2b1lsSzGQ58F8vlhHLg3MP5whvf
Rt0ws3Ipa0QHUyBP9VA4489/uj3s6D/cmBXxuyAWFGLsa4UyleSSpQqq0OdgOy/x/LL4ffrRQnY5
oiPpbOnH03LdZv4j3Vl8EYuDXsltknX1T5H/M32y09QedEydsYsGUYxWvOOs9IT3I/VIXBiI9g/M
mMFtZRYva6CspasQfz+BRHgeUKEl374en5ciCChtiGrG8raRHUDMbvYFILdg0Z4R8FhqlvFUia13
bg4+5MtCBBUYi7XegjsqLuEd/SCLhxIIbj9U9ZazursEv87Ns91SbQyF5hvytnB2pb6oJ9cOOhUO
LCH7CwG4DMbsi7La5oslSyHbuyr1tEM/qnvVxe7G/kwux1ZFHSFd1zK++pCCmE1heerZcBGTRKtH
qCTn4Y/aQBFaNPwtyK6twDdBZfJZaap28LD1GoCrHBtTU68vCmiNptyKSDIIBgYwvwHQA0CPZq6a
QzBgPe/Rdp6m9bcnvj2KhbjQAL8qHr4cP3ag7Unjrcwcjto28+eeS+1mDmNdOvuE9xhBk4ID27a/
4oaEt1ivob8SqlDXH6bvYbPBAPUuwS2fqeFEfGeJiW2nLjyb8eQW0tKLQ8i5cFAZ9x0fcjPjXztA
J3HwUFJ38rkWSq1d7siWKFGZQrtVLWu4o5KWKdlvlLnc7iALUFfMFMsEpfs+ouBDGAhR0IB6h+gT
v878+VkVjZgvysut0t4JjAHWtANsgwZi6/976bR1ywKLVTrJjb7o2hMTFq09/JxxRrLO6Xgpdya8
iaf+MB0l/F2bVxd3a9Yqxdx23OJC/m+5OECe3oLuX3tTTbErMQSXbblMnnj07M1Msxifg0OYoo/U
njihSPV2B8wvrfcX7OTSvQ2iQ1GGorS+zkKYHBnvibkkkArd5pHbTxpoM8+LVZO2ruYM/ehVJ+7+
ZWQj/rkvEFPMPlFGmBZOwSVnNt52tL7x5avHH/UBTBA/9X4WwhX4anBqWMOEOudB0xa3AQVQvB4w
ZL4o0mxeN0NJUB5XMV5QOnSooYDeEeAuuhJEDgP0Xp4fDK5eaeRH81eE0LZimpofWy8VdsowpwYO
82NKTJ3VJvgxMZNw4VmCrAiG/tvi0VpCKOJbrG+wlIHWvJvw16/gCfBaSFa9keoTE6GXB1fXxqqe
56rO5nzOHgYF3kQRxepv+nqliocVqYzgPwhsasdAoPaMWGwcWqIOkHIRcF1Hj7F+DyNZZi0Peups
Giy0o2f9MpvAXkARlUnwxNq4IMrHXaAjoUaMRumGmLsmn97bGNwucdZwmclvAY5T9nI/KbQJdhQ5
AchY47Eqd4mdewDH6+4fU+kaDptBS0eQzzPd0Al+AJLXKoMA6Om9hsaHyouK4r+HocemCvlhisGq
6iPZyRWrblcWMMpHQ1RSUAoUuyesEarv0dC2zuGKJI+Z2OdOOMDtdpFjnUxSnUP2sN9asL/wDD1y
1vkB7lwFnoHWbD+bZlndxCLlLUPiaT+Ks+LryKo0R/cL+T0xwBC8g48Sm89Fz+vOggAAhdPnAVIZ
2XWbx30vCKPJXsZJ2vW3NvcqmNhJGK9N4vPowOmpgbwNOQtLAxTcgHryvpoRDCzGJoWQIGWgxWGu
LhmXPSEN3Fa4YG2gh739a3Z96r2k9id+1VIBXt+6H2PfIOpVISeSZbC4rsYmIx1ULx2Vodxks/KJ
oodRen3aqxL0ZBmWI9uEMUn57HVXDF+8rX5pM0k1IexERLbpAiRzTkt+0g/IP43gVYt5ISUbvqUb
0ZtBndVddzJLQwpA1V6U3EKSlijGMHKwSyh6ZbnRwTZTjY2rtikLCPyE8FIULqEIlCPb8n5f1uq9
z8Lqsc88620V/xBC3pp1ZW0pgUZ0gONaGgj/MlukH9+nHBL7+tc8c5y+M2KQLr9wY8F9H34gbNYt
lIVa33/rGr4FZLQMK7V/9PIvwZLS8Y6SxzMlcLAPUYWUemuwcyr0nntSIVXVKdBssfwqSsTcT1z0
2Uytjw8SuvN74p29w2T+QEXuCvxNSheNhOBmZYx16myZOu5SosPm1Zn18ZS8B33jHAk/HEU0dgmo
jFj3eBBMmeARsEoDg8ViLp0CUXrNXvTtwHRdm2PsJLThldP5viFwvLiMlqhH4G7pGxbPfjnbATK6
qDEx0mxwIsTGbIzdmy7xZcOfwXVZJeTGDzs4uMhE7TxDHXfnA/5c4rbAyD+jg77uRpeNoXs+l0jI
2BrWjlnsM/DZ3w5KwiWWvNck49/DdrHhJlSzR1Dw76FjzF+NjzaJ/kOWasGYdStNEo2/gGnvdIMx
SYWxM3METyBTi043SEr5oDgwyCRwZCaAyo1p1sYP0qO9lYvAmcwqay7YGlvnPD3zAUdqIZ5UHJz6
8wTyadgueUeWGvzfShco7dc3NdmR200X6IjLP7fXdVno4Li2sdxgsOZyxjNXh1mD5bz5ASPdyklP
Fv9Tc/aneQB54T3a1aZ6fl7aBiN59lH1UDgBhMi4z4VE6apraAxOHbJN+i/onT5DuXre+urpIHea
qmiFWNZ7dcHBWTzTnCn238khQbx5jxS4I0De7gadfbFqsIWwfyIIAe18g+ooGgmBIzI3bMz3Pt+1
CWm5GAvokG9IiKrj0t1k6MVxqq831GSvZtq86pI86hBVjlvqpL63qlv2N/WWsmYBoT2Vlc2+xxo8
xdaIBZhbFz0Y4Ki5iLixB+Gpsgp/bfnZnZPE+EnYcfeqmj/BgZmN0HXxyd5dP6tcvq4Kwfgu1SWT
1/UMa3D/NEJWMZ5CAf2SZRGrE7+7udMy1hoKj8iTLcaCN2sPBnQq1HIheyfniXv6OLLLwInm5Gbs
BpvBvnskgBLm5SZ5Gh7zzPyPkWh78hE1+crREirxAJ2XYDyv/oA8boQhwhPgMqPSl2qNVYbaG/8P
/VL0CtwAVdYhiC0r+vkY699iLd7Ihs6nEczDiOX2sowfWg4aRZaZ3wilhRd/+pzLBBlgnDDWq/lW
ZWELrwAeZcvdinXwvHTc7xygGlwn6jNbUKIfpxIJOk6/TXwZZszWeOoZe7Txuij5VyNG5l0DH8RB
W32uCigVabsxsxazXnmv4QK8SDXuViZiob0gT6vIgMj80fJ2TKyaeF9xzb3C/6X6/+1MfsPDl+ua
jq5knuZ8uZCf1l0j7IZFeKIUPj/HCnjQR2yMn88Ps/bF2YZTfPPPfwz6M27Wi80c4vj+epH64Uvc
x7fEaCdRdkrlcFXx6LHxAZb4GjFQda5QT4zPj6s1O8wlCiUn3MLcSyeVAp8W2Is4WRA7CWRpuGsu
6zKno6DXeX/oK3oPDcQfR4CWE+5CtnZV/9TywCnY9s1co8zz6BuKPsZimFwbbgYWM96oXEKV6+27
BI+W5+3+bu87L12jgQ0XOq79yzqp6ydT32b+HBq+RdPhzAJmY17/DDXtpdNaMNPeizzkrcf707G8
W7ZnxZoKxrYWzRyv6D6W9Ad2xE6lBBnphJxzy98eXcRLsj5pRz9x5vBlNRr9g6WeCZo+jgEuXajk
PpHkbFvZgrh3RT+GirmQZOv+ZDVhub72P0Y8XnUgi7AnzRCw2AlWnHCSyRq7RTidpmqFzxedQMe2
0mlkD9XtvLRw7oEBPtgLAkpYRr7bCfiw+iDNFhqAafTrj9ppbJ5GQGUWzsSl1aQfBTb7u4yn8E9U
Ynu5I/IzOoI3c6LesdUcG+zODOPrwaHpKVSGOIAEhUa7SxWu97B8q7HTDkXBM4MFUBC3mAwXbbvn
g68b+H9Tq3JxEFRu2Dzq/UgWHRUw4+pUcmQGbVoGy5irFlKV0KJcG6uK/yRj7XlkcyGJ4X1xrONx
w/RehehVYmKZWOuZUxe8ufpA3o0Bx9NlCg1M0HBdkxxYS809tAKlpgxH9HbqGwISed3WmjAaPr/e
1LjUglmTFD2V32ntW5JYGr+nX+sR/NNJ5d1y8QSBn7UoYScjE084/XG2YNB9ateAr49gEwqhUW45
9mCzB86cAGZK34+hGXQW2lTHbtEdVOdHPrpRChZqvkVinQtT6NxJIHMdugf+v8AiOShTlkNK4MoC
i6f6uxIRnc2bDzlURVhL3xTSWH/0HTswYiF4JHKC1sAWHX6sdWxablviNaO8UU8cMtLeRoKJAhmS
ZPkL5u7r4Bwlnw7Y4pAkQtyohBAYAxGYsBku6VUxlAQ36i3pReaz2MDwj7N8FrTvafVdRmtg0ogh
1UtWWlDOu9caJoKr2ew6UAvw2RkTjx9NIE7oUn7ud8i+VsWJM2UYGfqayHFPKCkDCcVPJSYbDb5G
Zav80ak+K/FRYFGZjO7qR7V1U2aq6KYSmnP5Qo/VdyI9IJMgjQ1iJRYVPk+1VkS89NpJxEGqAmlp
Ir9+7LMTBFB02hQwQqUk5tXZWZk5jyqGGwW5M7dGDeZobZ6OiZZ0szGGGVvoIhLDSXCzqGbp484C
jq+unZEjK2NXHS7XUhxfMB4Ig2p7ODWN3h2W33VNNJ9jKfeVK5wVeoxKGVaEW98PUh8uaiQnR8Fk
c5opKDTtv9x2QN8disc86vWSNN51R4+aHBoyJ2ahdfe8sSNOwKg/sN6MUTuvQRJp7dAw3J1M5H3h
uEO1cBjPlYz/LpxKDyfyKBKhUQhstdOLJ5b5KLVXsLht0Ntcl5K/u4oh0kqNcXNQ13qHFhkevEJ1
WgtKqM5K/rCkE9LtNaO+sn/eP+dgeFHNWECDESwSfZBkzXATE+VggXWksjCO3XQN1Cxqh51lQscS
KvviuS7gVTxTbTR3dEaL0xUXPlsZ874mSbgmOrOSdODqEA50nkS0e/4u6I7eF/EbqiTP69px0jJu
4p9gHMwMyltznojOVAFu2vJzzd1vMKisc8kc83RigrBi/4F3hREEAWLGXQp+DoSKaJR/5KocHB6O
yk/l3B10nxGErbqHeHcaRrI/7isNbGYoXCr6u0NUWCTgMId2lu6Z3j1B63urkfciL2eCo9CRb2Lv
TN/GfflwEB0o5/Ct9YdNXmQgMp+FMJUnh1DDI+vGdnXu4ksTz+dzmkw5Ne/sZA+sIvSNkOQQLwVv
RTvpekfoyBiNxdx5+b2wVfqIRHDkcEVyzdIQKIdYGP32rqHwrPhENgRUFPLQFKRFkuAPUNevkHcY
C6of+Li3MU4SGSg1NZY9ia57GoAnwElxgmoOqb+lZVML4X8Vx83lciOwVXEacu8dKbvLRNvbjjG+
0WLjJk3GJ3gl1/0V7Mt4Uvm1ifT5v86SCLLkbNey216GS+X+v3k/fbRK1N8YL8MMfdWZoKw/YJg4
W7FQ0+y/DTw2Bdt/hIsYRZq1QnXaaFsLEdzZR6RX8c/1N3rGmam2hesrGP1KONjdY/kviGMFPjx9
tcfgqHbvfwjsGvkM8lIo/SGiQWmYfmS71Kn62ublLhP6hy+BFfY4EK+J6eF3FnzM/5q+XJy6P3OP
HngRjrZhJyVt8QarCupJzRJPJtldvO5uw+8vYq2d91mCFTJHbhfxAtoUL/hffQ1fMGwJ4ZxEOjBx
7l+zFYYWAo089dryLBqRSUc4eUp3BlE+Y0o5vEewSIz4SV+QHHKmoXGWWdJ0vjqJ6GuoF/d6pTcx
ZKCP69Q/tsJ77lvLZflVhimKRK7ADgLTU5p98FtlTCxcrLaFc59tINxRz1RiaKkflpmTDWGqIt7g
MCNO8I4Ef1gHihbySLtLFx7yvl7DP+qFqsPrv7W0uZyeAAZ7JfNLIVTlsSWt+9qCf4lwb6s6RRB+
sSmMfLyTEAW9c54glZTD87ih8W5uYu4CyO0K+JRgALj/cexEtXbUjzveqHjvkumKPif1I9tq6uiJ
bOh/TK85NFuK8VGJ2DZpOjLpMzRBz1yH9Pd59E29Jz8r310UTwe7Tlr6e2xb3A9xs9sPhSxPBmzo
3+nhNs0grFaIVOGAsLovo/PSgv52ZGr1NRNaA2xN+U3CBny2ARaH80Pb3406qt2XYjmS6RxZx2Ye
7cSOPW1YAQhIpF28o7ONfRlYm3sROuMlZAfXCO6ydy/X9A/x7eYfhT+phPCyJSWfvfo1BOsfeks4
AXlS616Hp7zAvpYTPqfygJ0U9Hhko2GO1W8q6c1c/xCcEFEQjRe4oFvf9hHp2aQAX5dn0rsf6/xj
W2uL2Cysg3V51AZH+HR2eGg6jSEHW1dbpY+c5BqezXAzk5hLH/LsLpNYf4SD69z1fC6JJmNpn4yK
2yvpLDiHZLVtfyngpPrFyC2RSJ/SR9/GXDe0l89c6Zevy2r7X1xGPeOKMyV4p7w4GL0Cbu7vimbC
d5I25uDpc/uVrsRS2NeEaub8UM5w30b9BdqWx/KU0NsjLt70fRhckSeM8o8ARCnh9T9c+B4hFby/
Hsrmvz+2jXRhXDm+a/VLmD2hRYlNUC4bcZVcNcRNuwnKQECilONtDDxbIcTlAFosD8bBZZUwHHLe
+xozorCgs7fdWGsyHvNpOc379XHzVgV0AF+XLCxTExAblZUiKzOlEh5LtL/fjqxkazC/XLOgqDj7
IETlRKZqQ6QzCAWXhxG+KA9b/FIvleQJOo1ODbRYCOEzn24/+xVKBLlD6cACVOlqVSftQuFiVCHs
72x6/J5uS9Qt6emUrXL/YE8FviHVGIYCHhH84WS4VZq4HL5KxcVXsDF116U8usEDz3y5k5QyvfiY
RAfU1RMD85jS5xPqQD0mLe6sg1RW6S2Bol795rl6sm8lm9sip6TXs4qcnqORrgF5F9/eFH+tjDBx
AlJL1/4DWV+Id/4sZ14I8nETJfZ31Pcpk86oHsDp5c7bCfLAiB8mP0Jd0ysCb+fd+CPYRwytMzEp
nzdnyTn+eq0Uh8Pamxycn8hxdUxnsbxOxh20wtOlRIp8lHki0YUl9X87gcqmVIv1l+dQlzRxCAdL
e0DeqEn9cM+c0f5xGROSL6sC360WyIoIzBge7OB1rTTjvZu9VCONeWLX+3ljQqfkcEequDNGWbF3
vUD2j1vr1x5iBzgcZgcfiSAKsy9zxEXInYTsnA4CYtQcgRK/j4NC2HKQtD5ttH2WeubGgv+sRKs+
N9MtsE+yOjiUtwmpf6rL9rgnzv2dJ5lIDKkL0iWbqrnoMuOvNBwEOEWUucJ/xwRJyCcxNIl5ZQbR
lwAfA9CfS41NHd6kzlYHjcLeEJV+bDmlac+ZUschyg0wjUUNlHzDs0LhB8/udjiW9Jutlz65aGkF
LutXFDWbuxDJ92mOD63XCU+nOWodXqy0MElTjU+kZxbCCDY6ubZ7E8r2pZyuhciODW9E/PRQ6Xa+
4uioKOMh/1AdnrVpSUVqIJkZ6gKuGd4SiYPkp8GNI11y08XGy90I1Wzh7fXbmR/ajUnaVNma4vvg
QOzLduU8dpT1wer/Gv0J7AulWUJCoYnjgGYZiIZAppx6agcr4MZMKmR1cSFSeBvNjhaGf/OJJgtm
Xrp96ITXx1c4S5tKcB7d0KFtggktQMexG3xbqxq5XSPQp9uf1Fx2RQJSTDh/rT/6vc1aur8dYWaD
6UPPAM3816js9WqP6Fxm3fBRIfH3TVUI4u/DQ63/xjbxbXx07k3YTYnCze+BksPxAHO4/kKTO7eI
Ud+mpS4BmGEatP+UBBvQceIDsmvC9iEV3iatV8wg/r80XiQBU3eJB7kwAgs1wcVhi5xp6yLDaqTE
+Xy1PpmNwBeHXzCY0iS/tkZBdCbXZXSeRvBzedRnYI0757bFtdNoDwaJ5/lrpkywn7WM24X1YnQo
6yAIO7H1j50O5h0qudNBBx0TGSreB2Myn9Xeu4oGtt5BRgMmC1p1hVZaPtMYN2rkH387lKqkKSRV
u+TuXIlDZ/+6+Z9yFx/YysEKeItH+PNwx/2Q8u+Icgwflnj3sg946/OIt6LmiRl6DPZtqDmvvVCG
1ygxmlRMyI1Et1yauUrBty4cXt13EMPisb6v1dV7ptPrL3hqMgbRCJtz7JNHyNmqW/uaiVbAUifL
GIYUk7YfINYNPv8BaoWaivBkm3sa+xvd2guYhiUGdxc640kaLbsXGDe/ZF57vuGPvCXQ5oN0JSb6
Yw46el8w6Nb0s6g8TJdFG+vrqVrbywH5jUZrH7mG13g+fyUPaxIOx/2L2hu7LtDfMp019O+yFgqC
ZXn8UNUAtbRFTpwqchsy+G2vdd8zwTWE2nxbxl9CeYZGbACLW7zi7yRzhpScyN09nnJMSZyv424F
OyPxuEo+S9mwJQjTIsbPdgMaJdsBpmvkFnE1jA3j8iq1PuPU3i+f70V5s9yBA+FFlY1K8sOyseRJ
eAamtJ80N3jYKU4xcqW1KBlOAS3Wj9QoA5y5003ButWGBDkSE8Utyb5fH3oxZxAOzjn9Z6WES3A1
Rgcr53U+gqO4e1QXpuUO87gC+G97i2QIJoyiq3rnaIURHRR3Ksx4VMbFpHvmLbPSaNTAhztUz/eh
dJTyt9tRu3zpQ9Dh/CdC9ZaIqP53yKMrPbyoOdG8MmNrcIWS6WoqOsos7vqoA+gzclsWiChWDIoW
TQTCokJwINUN7VDXD/Ycdee/G+RzlDcOunXz/NdzmNUcNxxNOrtB8UQq9warUqjMTH3OlZ7n26t+
Mr8p8jwVyBlblG2c3FvL4PyBgEJW3Be0HB/UQAwbvfWb1kNHVjVt0zbUv4vviAntotSXVOKscva2
/wDSJMAnnK4ECDsp+E324q2yu2Fhc3ejKXZadPjfJis6PRHS3qMU6qo=
`protect end_protected
