��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��а�z��+�_� ��#,n�x삢~��3�[��'�[\�g���n��P��u�L<Fr�->�-��s�Iz��ado��Lwe^a�e|pUI�.%��n��@��c��;��Lv�3�!�VT�_-�b|=j�V!��Of	�K�����Z;�3��_?e2��-K��ꍢ���O����h▜���c8k�g?�=0&V�Q�Y��#�913F�����:�Y�QS�0g���_��h
zs���Q�����܄m���K���&�,Q{O*yE!_��|����y/��Q��)�7.�l���/��0�+Bb,^Ml{fb,�h9ġ��c�X���'%���K��S�{8��~+��E@��B
�GxN�Z���ġ�W�a����3�D�tPN�&�������Z@��F�6�|��F���`IUT���7Is��R��Y��G�~�p�����_(����K��4й����#D�?�IR��K���<Y�'a�&����m���%>>r�v���̂��I�2MPjV�����3�I9tsre��s���dj�?��m�h����/��q�v-�;����Q�ׯ2ЬO�p���I�GHT�k�����!��!͡-B�Y؛	wp�n�!|�f��x&�~%�<�*��醕i�nkf�9J��%G;�y�J���&��4�0"K�|o���/���e1A6�/��W6%:шD>�Xu~DC횁�K�%�=�.�u����W�o9�����zƝ�Ћ�R���(��`��ch���!����x#��
��ʁ�1��gM�X���{B⁅�s���	14e�l�@��^͘a������d��T/�^�7=î�_����M�"H�A>fO�D3��
�՗��Sh#QǓc���`�&��,(��o�3�����W6o�	��HP��|fK�smm�Dc��m�'?ϴ��n�op��I��ᇙx�݂�~XU[N�����V}��z	{�r��-�w�$�@
zY���f���`�Oc���`��Lo�*�0�/�j�Q	��n;�2�d*��^U��@>��3C�Y/��wn/vs�s�(��`�T��;�o��E�C�qX-D�H�oe�$yhZE\y�{�M���	��E,-w��� "X��:�@�\#�L� �����ZtB����0MFN֓��!��-8Ï�Պ׬PH�[�K�.�}��,����7M~��:Og#D@R^"�d7�AǦ�	D"/`yAP(�22B��������6֯U����(�ͻ��ܞ���#|���z����,z�:�"�#Ŵ�40����w-��pZ��x�k��$�X1d≮~�pn#��S���"s��㑛X�@����v��L�]��ַ��f�l��ӂTR��.�]��c�p��&���.!��)j{`B�p����R*��O�F�>�����V�JD@$0��T]�CSd�<Pe8��ڱ��K�Q�N*�{L���Mh4�"8���ZKk�����<s�c8t��`�����Q��%�E�mȟ�e��F�oL	bx�P�b�A_�ǂK&�=��XVq��x�ko��n�B2�5S����@Ri���WY�q�#Jp2
�E.�p|��䁫o�"��Q,�h�Q���EJJ�L��t@�Nw��_S�˩	��o7�|M1OPi�WD��$X���Q)s]��I4���I4�[T���{rn9�VA��K~��u���Lv�S[z�U�f�L�0���̛f@�"䎎����i�}��-:u	*�Iu�iD���̃��+ck��')����+9�3~'�Bߘ?�态Q٬*mu�Ds�$�=�B�-	zc2
�a�-#:+��ڪ�\���!�/����4҇)^��.i�2��k��Ҩ}�C��f���\��6J`�	�D]O��}k�0N����id:�K,���,j�i%�h�q8Ո��MP��HDf��>
�&�tfC�n�^~���^ 3̤֮���Wv��;���Wl@����N�SҪ�_W���y��kOx��9�)�W`7ΰS}�(��Ëm�H���ק5V�e@),��II�V���'G[��i[	�0�j���+H^�Z}
M�zw�Ne~�g�8�[#i`d�sԫ�Vm���m����q��y����aT\VE/*W�}�pRɸ_�5'�Ѝ�\�f˅\I��}R���/�x��^�z�l�}��3���M:I�㚝W�J�����H2>��̽?���Ŭc�Sxg)��Q�cb�_����m2���m�v��j�+���Ga��O�ŵ�D�Y~����AsR֝e��s�^~�)e8~��N<���,��N�X�\���3���دh�������?o 5w�f@�,�)��h�H���ݝ��t�a��`�F�"�R�w$�V36I\��zk�ς�v�0�S��Hu9�o��Ƣ��n���k����yז*Ѩ��E8�u�_=��yu�"�����`w���Ō��T9���.r��jF��>n��H�N%�z>����T��8X*[��r�0�ل��&j<�Sh��G>�������S�^>�q����ͮ�,��I��0����JX��=�p�}�B����8�?z0��2���Q������_k��F�a��Ҫ��~Q�� �vN�$�H\����ܑ�y�6ゼe|{��h�xҢ��#��G�W��;�@wd���&$mEð>�&������y2;C��2
�����9n��J{s��D~���L�Gb�������p]����d�v��>F�������D%>UofN�rH ��~>`�����^�	[8{G��t���ֶ�5
~o��c]���^pqR*�J��`5H�L�Nxԉ(6yY~���-3����npCb�QY�{�O>:�tv����X����!�*0��*\��Bv/UI���Tb���Cv�@�V �s���fď�賹l��O>��+s�R;;�|�5ha��᥼S��iew�r���H?P�>�(V�奄)	�4_�ǋQ�!�]�Bk�9�>	��ҟ���k�	!�T�Aj�v3ȹ�����B��t�w/fq�z�!Q����'�dG�Y��ܙē�pH'�����!�Z���
K��'ׄԯ��	�XX�CڴP.$M�f�.��s,X���:�Vf�1�"��~F��G�Z��l��\8W�3��R1�#U��T�k��W��
��#g����Q�Gȭ�RTQ��LZ�et���B��!���]u�D���1�y�ޢFM��#׋�"ʲ���x� �H��<�.��[w�r���X�G��H�0��lJ�o�֊��ŧ�J��0��e�k�'�V����qͺ Ӷ��,��?wղ7JJ�b��Z��S�CG��|��1�Vyb�p�˝8>$-���_�.��@t:Q�[�:��z���N�Vzhf��,�SżNm؋L�`�uJys����:)o�I��%�7�^cD�[�L
�1���%Wu�f	tF�����s�M]�L��\T��ɫuk%�2	�J���7����w�f0�hq���j�W'ɓ­��6Q��%xlo�l�y^����S�H6�ϥ�P��DNrV>��|L�T��\�F�D3{t�i�T�%_$�������eJ��hʮa��u��<�����>�'��Vg�Ɋ�ɼ7�&^c��]W��ꔥ��z�/-�%����7X|FE3���r���w?TΆ/�*g��%��K�)�(���$���ƊO���=�����{J�ee��{�j��8�EZ ���8ч�cL�7�if����c���h�IN��xvZ��K2�س!�;�\��-�I�3�4���G�`Q|Њ槒��Ȥ���͋s� ���*C�
t�4�>���HF��C9�Ӹ��@^%�`}o���6�ЀT�;���t�q�i��=_=G,_�ӽ^�*���h��$��-ٿ�Ŀ����E�̲ˠ�Qs=��#�E�\N�Bh�2t2��ƻg�D*�2a�wQ 8|	c�����;h8wKG�ğ����M/: �C�}A� ��(���&�^��[��!�J\dw�3*�o���Q��������p��P�;W&VI�\`O[0я+4�2�yG��˙�{K� �?��L]����n����ե���-j��5���n,���蒜Ɇ���ܔ��j�Wc�B$C��u��@:�'�I�QM2u1`ʪ|4�i)�EB��
��1=P<8�y�4�W��<�v�?����g>6��V72�)�ARC�W�#�t�u���(5��-NͰǋ�^���4��z���R���U,�^D����2�'�f�0N���+b�'ב+���x�Kn�W�<��ᚫ���=�C����v�垶G;B},"���C�?��Z�j�v�ۋW!�kK{㋴�w�Ij�e��pS��)✝�F\?>y����z��ro�N��s1�b�u��(��Êܕ4~90^�>�����*��<w"���r����W�/J5�� ��j�_u���W�{�(�/����p�q���,j�|��ܖ'��?��$�,͡����+7�9T����(�I>�
O�|���#H0i��KDX(S/'�R��p�7�Sy�^�+	8�w;���œ�X��<�Z�,�>�٘x�n#� vH5�f�\������_�]��ǭ>�<v�_O�/C�g�(k��9�
%B�ӎ)�����ƹ��v�"�6ѵl�v�ٮ�(���
#��nPq�p����+�4�$
�2��D��5���ڨ�O6(W]m�(��a^.�J*w�21�yOw�)����U�����2��,*R����C��]M*5[���4��ƲUߤz�-�eM$/k!_��k����)�2���G��{�}P�0G�Al)���46�n5��A(���PH����B�3�[/�w�R���g���s������=�?����ݗd��*�=�:��D�r��?F>,u�Q�_%B()@R�vY��cpD�������`�LV�):���@:��k�Z�z�m����Q�a[9��G(s�Ua���+h7WE#)<NE���b�(ܐ�D�
G�(��
�\��&&נws�����G��r�?K	dż��+�@< xL��>�c����;�d�����`�(9�x=Ϥ�M���E�k>[�����ļ߲��^������D:�Fx��Ļ(�αZ�ҳI��r-���q*Qi�5S�2�"�P��ycof�}�/��<s�n�U�5f�r�.L3�\����]H��'d0��h�9���dK �w}�~>&�X_h3#����u3dA�]( �����E���]mo�?X�,8�����v.Ƿ�i'�Ls�+�g`R�>����1{�r��n���>2�d��o/��o�-Z�	X:$��㵁�H	;�Ѡq�t���;I1���Q�|�4�p��K�dp�F�='@N�-��J�J��b� ���/Hq?�\I����>�W�@�vp^�X\S�%��xk��l�TCz�a��1����O�$	4t�$ۡ��C���UX{��X���n>Z���i��x�'�/oa��=$��
\�����'u��7]�a^�~�R6��4D�W7I��r���ǩ��;R ���d��Yr=t��a�O�sz�>�<B2��j0)}�����r��?��~��d��,� �1����`�6K�=�S�	'sX�.\W'� [ƴ���ʝ�fǨo&v���C��Io�#'��UC3�f{����Y	�[���6*�2�4�v�o!�ND��rU�<($�{f����޲�dL�j��Ts��q��>��af�F��jꕩ0)&��3M%��.
����!�ivQYl0e<�Ib��HF%��t�����>'�����?�-�ᴂ|)�v����a���n�ߣ�����˚����-q�
7ȶ�i6��3ֱ�R��/?�2����f�-��ܔ��!KB��"��l����ۄ��a�	K��<�-'�Y�Ҫ����6�@-̲���}!Jh�!�J-��|�ŉ���	n�Z��â��D��XH�3o�pշ̰�_����� )�Rb�hP�jE�����*��q��Bڳ�74�,:rc[�}X�6�Ίc������0;�aL�UT�Ƙ����Gq4��*|�岹�+����P�'�]J��.��$�L(��@1�hnA�h�dM�d�έ�6z�������=��Y@�B{���Qx����SflKz��*	�֗�X ���~ō���c������uJ��V,'�ր�E�C� �b�[�{��^`uw;�`Мvl��T]	��/�� .��E�l�RIP�¥x�5k�����섬n|�d9�h�P}"�ځFo�v�y�Ӯ`2����T1y��̛ 3[�x�>J�͕��Uܫڊ�T��1�:�a�Y|I�~���C�	F�Hӣ��XUSu��	��Nu=;aw�ml;�N���CӘ5)i�b��ǂ��D*���}%_��i^}�x�h����L��Fsu��Fd�q� 訵�v�|��
����t�%��~�#�fN�.�JH4*|���,���E��vn�<F�D*)�r'-
n�F�����>iV�{Un�T�XJƈ��HcCh�]H!󋲖��?z�tEl޷,�V�%�B5O'��CP/甶������\��Y��V*w�#���fy��΢f�@�R|T�]����I�j���͈.�_�Ѓ���=B)�.�<���2��m�E����,����� ��h�w[v�	ǚkϖW�/���ʺ�F��r��� �Vi:�����"xW�4"�[���@�A �{��M?�>3PZv+����}�A��Jt����`'/�j�},J~���z��5�n�
�4~��Q�+Q��g��oUA�>I�T�L����v�]�[U��� `�OZ ��\B品qR�I����o��(h9�{�+���vo�W����{���)�N<�p �h�:�,[�2��M"x^hRipV�@��z=���-�<u�����4ׇ��J�m"�Y�'Y-�}-�U���fE@���Ό��VNe��g��T2�0O(Lۀ�hb�p�>X�m�oLJ��W\i����Ā��ճws��I�s�����!�"�caC������&�U��V�r ��Qn{��X��2�%,�Ji��vܚ�p�J��ER�p�����@����"���xH�:׿�c��D�M��M���,!�e���i@ ̗�:�ן� SA
P��=Z��iޓVc�"��L;�a��2���lA1:�Z@]��L3H�'�w�m�:��#e�+�Oo�݂����[�RFq�n�����Ύ{�<�~險EO�#�b>5n��4Kڈ�P�/��Es�n�MtҰ�w��h���P�bu�i�x�jj,�$#�[(��w.��]R�[�s�j��a�M�smJ�����27r�� ۾��FmLw�!�G�7��uW������__X�F�]d����G���d�,���(n`�����#���"�~��La߈�z��i���,`C`פ���˞V�Ɵ��BȌ��%�wGǍ��8���C{@�	�lS ^�~��n�g$Mۢ�8��-�K�A���	UCd���ȟ�|`+����*L������^=��㷏8�%����%Lx=��%��@ӽ����Ѓ���Ҽ�-( f`Qs��r�.���P;���2�b�"���*F�s&*�I�ft(�L�	/�3������������Z��R��Mޞ��G�H�Q�sT���AIdS��k�V.:���>���O��	�6�|j&�J},�K�5b�{��]��Diz(c	�����F��'h��*y1Q��G�k�snf\������X�G���'z��d��2�����Q�^�b��5����̵�j2c��~�78
X�!x�5]�n�ÑK>%E�=�"���-H|�cI��U�"��D�~�R	�v�(,�P��/�մ��m C
n��>3M^8�ǟ	m�f��M�TQ�>F �3��a��S������B�
�,����2�Em�OFv�d�½��NE�Nra��{��f�����]	���zJ������#���;�^CW�uؖ�r����
�3 <��+�3�zd?0+�ۇjo	�B7�+�����Wn�c��r�����D���.��s�����/�k��OE@�,k!���_y��
��D0�C�\����D���1[�[�HrA�իU�Լ.{.��%��z�y��-����y>{��m7C]K��P-��
�f�%��7is�=�궅fdFhy,�e����9�532�g��P�[po` ×�q��!q<K�DV{������p
Ywj����M�ļt܌���/�4�&y�H����-U���»eRX,ϳ9Q�����Y�A2�3������^�u�Z�w��g���ȑM49p���r�Z�`�S\y���<%�3����=���@��%Ք��7<��N
b���s�]1���#�T�-~@�k��c��+�g��/���Їb��=�gy���=���8N���<B�D!��`%���~�[�R4w �}��p<�`� O&�Z\����ϬX-�_ԥ�j�K�by�QD��t�7��e�es�3*��;B��HI���;~��N�z}pC�ȝ	0�r*����m�֥�(�F�����6����}R9u(EY<�Yl�͜��6J��2媺���P�]5N��!kق6��AD���(F���I勌�_ś�M$	�挀����xwt�7�rRx,O1��n�����O�Qm��ķPI�a@4���Ũ�>Ϛ[,�mvYD�)GƄ�".(se�r���y�	ǘ��?]�K;��}!��^0��R���z������'O,%L����ƛb��.�h>U�����q��8��a����$p����絡 <0vy�6䝒�ϳe[h�)&�l$���Q��,=��HB�ٽo+Sb��،�'ʃYv��C��H�����w��rvP�(C�4�����������ɐ׀�d����t;Kq�I�O߳w���5-�뼬��s}z|/;e��~$^��6_{r:�bwfO>M?�pa�@�xW�ڝ��7�%99TEԊ|3\�j�@���Fq<7]�^'��*8v���xRx�l&X4����Y?���ٻ��`�ē�`� �ᒳ_6��s���3GTZ��J�~}�"ur+v�F���dg�|!�YuG��"^�|O�y	�!W+RJ5@==����gC擟�:�ҢA�"C,�м�~�=�����Ycz�lˊ�F����i��c��5Q�
�n6?�-���y&��sN��x&����r-�24N�_6W�#0V��]�6���P�@�#cR!(��U�Z�	�8Q���Vl����҉�׽��ؘ�[@�C\$����	������t}�X��&P�x�����w*�%��M+��[�&IbW"��ZA�pp��1dP�pU��[�Z�����Ej�2��X|�n.ꚏ���u�/S�J��V�����p���j�bD峧�YF�F3m\)��2O0�>�ae~��D�L�	����G��!b�w^���%�#��Mr�D��2�bp��\@��.�D�|�M���{g*2�����#�̓�ݒ�f�U�
�D�����H��vG^��f�6�I>��<<���WߚD�mmY�GЉC�����Iz� �5s�+8M���#��񣺒bH���}c"��YgA����f총��UB��M�D���S�u�pfRX{%��'4r��U9ƚl��I��{�҄�Xv�Fr��Jf7Gz��x(;�X7���+6��D��b�t�� �/M��4
��\��f��x,������
�;o����L����2`֗�r�G��_Ɓ�)#HQ�m�̻�d���L't:ώ/�E��ގ��Rh)+2��a�~,�V3�}�m���3O�WUS�I3��ו�U%�	3f���k^���
I[�w�:7ɃK��ք�����p����|���:� l#I�I�TG��I�G��4.����u�PY���K 3MU���e��"�U��Дv�k�o�L�.dj��������Ɍ��d<�E,� ��;�G�6�4��T�}�a������%Ȏ����0���*�QK����D2`ڡ���.#�\�^���F����n�L"((��9vΪy��Q$�0��jk��-�2*{��=�~�7�Y��?�Z#�e��mV�USC��ȧwMơB|���Vqa�ܴz�@���n��b�����y$p����J� ��6��H��gӦ/^�!��P�>�K�D̚�<co0�rg�0�؂�^48��\��G�?�N�1}/��pa#,��#�o8�btwv�Kj�����i�FX�9�G��ݚ�E�ZL؟�>� x���り��yP���SLsXFBg�I����B&�+\�W�m!T������:z�/�f_�V�:�IZ�= ~/iھ����x��o��׌'��L�2�#%�7���8)B�BRG��q��e�-:�<�Ҕ�����YJ�^�1��ͦ��9kn�[�q<u�]#|bZ�]Mh�������M�|h��R|R��ȧ��]�!�XD�:����))=�H#v�w�a�)��˺�{J)R�M�)ʔ:�A��s����~�o��	Y_.�G���{O�9t���B�|��7�y]���"*�pg�a����}�*T�v}!�O���j��G���c'�MˆO�3��1��ѱ���LX$h����LHQI��.�8m��Q��?�KAݗ�A�)��Q�~��·q{���Z<{��r�����hLv�,��?�8R���?�Z�U��Nj�x�$4s).^�]�)�������n~6��]��}�rO�����0Ö(@�=�d�NQ9Sj
�Js��]6��{�xC����_���2yt?,}iY)�l��0��ɕ��L� �+5B��)�^�X��������P�s���v�6I��F]�ǩդ���q���t@2���I��$N$;�D!L�f�i�v�u�WI�%h	Bp]���nV�$=��v��tk�����F;r�1�yR�w�<47�""���#����Ex�b0�"�c�-�-Z�Ќ��N:)��mӴ��&6��a�){�/��5����"�g�����R��� 9Q'Bw�l��T�y��[��_�>�
�5喞 �i��)b2;ž���>�a��1���=��������ƪ��u�,"�a���Lا��DM����ǿܯ=�M8�nK���	F;s��!ܰ�E�(m��_�Y�ἥk�r�t
{@��&�7�&N��/G$�T"�d;����L!��3�٫ +��!ڕy�0.� A�l �H2�������K)M�WC�Z5���$�Bkl�9�b��w�-�EnW�g�b�K�����\Y��c�]1��ͷ��@kͶ�_ ���j'Hvߎ8R�ӝ�4t�c0��
���[,�h?H��&�*ԓ� ��èJ��G�0�Ι����績�(��z�>
0מ��#���[�-�y����jL4揿���>�H���8��ҵ��H�
�箰DM8��Td'�I!��ꛐ^�@Rd	���hIZ |��yg�G�+�1'ع�Q�}������5�"5�P��&N_!��v`���iu�`��:�˙7%���f�>Kp�(kw���O�̋�������)U:Դ-��%�U���'��±����`�={f�R?����6��5����=՜�o���P� �Vz`����������z��,^�,o���U>�>�̏�/Hu3(�q�O�\d�_�!l~GQ=3	"��g�7�ꄞ*����&ql�	��D闭<B_n��0I���j��ǔ`|�ҩ��<�;�+�{(���Y�{��
�ߋn�`��ūAaa5�3���H��/P��^��{a�>lDnj�i�p"��/8��^8�UT�Nw�Q��s2*_�܎��jސ�W�����+A�w�y�)	��j"�\�~w���h,�i��A�&�K���IRo(`�e��X�>	�8�	L)�j&l��uz����N�B�JnDZ
Gq-��-�?ƽ���メ�[��?���X�Գ,·�0��e*g�8�ܐox\m
D�O��'(n�������/�	����Y���c�}�-'k�e�W,u���
���M,_7o�E����5ڧƟ5`����I���M�T�t�	�aM��k[_�ޮ� ]�l�<@�����Υ-�h��Tx�~��6����0,_�7,�W#r����$�nh��R��t�nM,g���箲hO,s�֣@�T�#�B
C��F�ߥ���mСӆ͛;�oSbiׄ��AgÈ8����C_��.6�I��Zp��B��$���%e��x&�z�%��(��NI�b1����T)��{�!-Fj>�֝��cQ����F(f�;i��4|鉱�/�q�`��p�#eun� �_�[�P���ly�8�L�R�X�W���e�� ���"�:�6<l*?h��Z	.���2<y��6)���.�9��S���mԊzA�I���Bl��/@�)� ������������lh~0�j�B��|R/�}���p�6�k�c�L.Aw���R�F��*�t�!���������НlO~��^�����0�2MSt��Rt�H77�H�m�דyc��8�JƲ�'Χ�0�ܿVX���h��U�/�����w�7?ݠQ3P-i=w����A��K|�.��XbLuU��{�CgC�a$Ssi� M��[o���7@��3P/_�͢�7� �,�dA�,���6��b�K^i��Du��{BC��na�1�`A���*�@��B���8��C�ķ��{̼��_���Q,����%�w{��2��yW?��n,�� .4�\��X�=ˡ�wB�kkɈ��7ؒT'Ay����CV����1?�M� �sǄ�<<��)���'���Ö˼�`�q[�]�5�wwȴ�ODZa�a,a�O�ɽ�)r*e�tA�4��d�:�j}�F��U�p�}>��E�����W���� �g��
pN�W�A��K���\�B������0p�� �%ޭf)���B,��,�9E�E��h>��y����`��4T�{��#qY���_s��m� nU����F<�tk�Cb�s��)UaơC���#J�3E�gn3oU�:���17�/�����0�y�lH"�=�).�\g%�:����n�_+��2��O��P`��`�A�\�,�QE���)o��׾���:���Nl��M�� ���:R�9�՟�m�BVZ�Б�L��bͅȒ�f��ޏ��dN�L[u�ڨ���k� (	d㈟WrO�o��p��"�L�|4L����X��a��)�T�yڙ�v�A�l����zM��Q�����|;w��srFp�υ}Xb|���P(p���P,)��˦�"l٨����E��y�-�m%�_t\"$L��+0n/��z1w�2�^2x����7K9��<���Zݐ�(���f&��5��a�V�[.X�_n�=>u�:l��e��8�۫���U �D%�yZ��V ��rQ����r=.q慃sx!S���[
��F��R�Җ@�&�?ط��|&!=��ƙ`)c���j�Z��.(