`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8400)
`protect data_block
49gv4y+bQMqMtP+mNNuWHX8SR2+25oeygsJ18RwLg1wHQu31rNWcB1pyVgqOSPGsEPHwfiffZIpO
DUk7CaZjKJAIVcQPBae+yQgOWgBBkqHDbutOaKUy5nypfNX/dQxlMUESWjutFjaQKwoi5mDJGvxc
2oYUpG374x511uY0/mX1FZQEbN3npuok04Hu0Y71PLxU0RrQvrtq3WquPPWAIfN+jTOtDPWXWiMD
2tFxRIXlJz/OdgZ2KfBlM/7eERHY5+mTLqMT5UgNhVoPFfT7TjrVUU9pPuP7A+cmWyw+KIySl7Ji
xRm9mY6w0CLM6e1SdwivMxdFAyXiennr10uFmln0OJTqPocwA0I+2+iFIiN7PscYSN7SH7fVPrDT
kuqOabgleLhXPfB4xJqKv8ncuq/SBp7SebXFXboiWbR69zVsmPgSk571LRZLXyTCV+3ASfEF+ZU5
1uUBGJH2bHTH+6xZknqc8oEFDTvCTuwEfxHxBTaL2HPVvHP6mS7VNhlCsHCh241P/27GbWOlswKu
rULRIMuVXhlUgk/8Ffl5xnlIytocPiNQpTNhsFfgQxFc4baoqAWNU0hSQWr4pDJFzT1iWaVulGnm
p5f+gbWPzNyZ/3xSqIP+jkOBYXPg6GhiVcU111qOhGkN+bg58i5SCw274aHu8yeuU+r+naoD9iaj
NU1XEq+4X2+Z9O4CvlK/agA73KcjWGLLYLf6WJzTCXQDEcxpmT6v4aNaPOvoMG7IUQhhMBJnPEfq
wOTUVoRTWNmNf/gYojlNAmgh1WI/29Ke8Aks5tBMAV65PG8/IoS1lMLHOXexi2ic4NZ0noaSb81v
o2ymuYTES6gQ9XZXU8Jz6fhQIFkLEWwP+/GCF2QcnTAM4CV6+kBaugkh8UqqntJLlyDwkIJJHSFR
eiCs27w/HARpYFYWKsMRU54Oqr41C7q3P3PIbZqtE+WDdsF6/BzOeOJET+72dWgUHsKE/+lzD80E
yfikKb7zen+Iqx6TRFz9WC8tRJPJVe6EC/sGL1Lbo1p6KPbQQadmg1k8ZRoUjBqT9xgZArXTjwFk
ecSsfTOfSzF80cbTtxC7ZpGdkPzdtTFOuEimqS6hTR3FX07P4hj0JRqpUywAuK3fUPdKWM+FiFuH
7zUpndaNs3R78N5XpTvvNUguhAJv8LUEwwoaHs6WYjF1YAOLGwWHnnZjR8o1Wsnr+yyr8ggqsait
WgSnUWZZ1Gc2uPuDgfeRUmZF+aJy5q9H1vqEryequ+Ml+9W1ZqUWFSqOYwI825rEvxZYLOdwxYgv
vuGbYvZ+YUppJ4aalLRGej8CKxA9e4hXFVPyqp5rePk3pDPKal3E4+dO5SATxNyKeUAgtHFuTHfn
wLmNGfHMa2a1HKwVJAwZpF8Yw23Qk57OKkvwR8wFrMrL9vk/C1aoCCMPIHIpkkHucYgOU+LnBQFs
gpAZBjB6yBX9pW47kiTh7HP8VJX2dpO+msyNnk0X46rs3xpXFZ4C0+ghUFQJVhRfpKghidmvJ6Rf
89gOuHa+KmygQLxQP5mBBoGBiCD2YnPc0VN/E1BeU5Lrzgw4UGq7MOxoMEpb/foSUGJ7SxeD+ufD
nPxNbNItQs2/2mMYIa5pbzGuaFnqk9EacU00WELjhIPSFHsHoojy1e6WE4klOTwO1fdg41VHh4qk
Z5nQmWwKjwyUYN+BL6FLWRTy2XDhbhLHlU8+oaUCi4waVWcikKZHfU9S1tGPKH304ZlG6lOAoDbg
aG2v+VO5WC9nlKXWdYbC6j01XgzG2N6uNgsCIY8GgWZoVKq8ErdcOdm7XEf+On7cUHpfDAai78wx
MZstinjnktSjTw4DaMbrR4V1S47cwVVluG50lyvoUgGDh3ypWH27GGP7R2GYJFaXJjIh79mcRFBc
GbJpygRXZo8EHLiXNYf0DgMtZ7loCk4LLwgYSWxbQbDDqskt5aSWKHOBc2amd5ZzI09E255mGJ0F
favDCjAJVFOQ6HO5DfEAMRtM1eQzt2LNEWG/4tu1LcF71YelhBqrpjAeC8YRmgkXw2tHxixDkpxi
r268nOQQ2WgY4NJBjdUaMrAKeLC0x+KpnuxqUGDZWCfKGqkkbgM+3hdFpc5IbQqqjR/7gUOIz2OW
wLY+o9kgrnh1J4+fSAMWLASXoQ6lim5xUT8mEfCBJSjqN+U0upg8km9WeX4sSXrUGZ8Ji4Q4hRam
Tv9UkTcPApxAD0gidQptBTmwVtkk2NpBn5wYYAn8TAZhLDD6/Jt2ElCK3knHzpo/U1q5xil8jfEo
/iK+HUbBt+fpRXpxlrMFWeK8ALsDQEvYrI075ITOPdQ0xWb+ubXgiM01doRyhmNcHSNDJGLsAR5v
m2dfpnp2Qdm8s3QrU/+GlTuvM+7nSNgpL3ndcSL9ufjKMgoPZc4HRuTjuyS2f2glNhzXesEHICyB
wwBSx7MxY1xRMK38zVrCKZFsKbqCJNtuHjxqoX3O09W22Q4DfoOYDfoPWF97ZjPAOZfSCgRpU27g
OtJM2lRRUkSJLzCXbDF4ks5IK1o/0/4aLOLV66a5tlVFdSczWfD3E1wrWyaCgNakjNq5IbQbxaXq
J/hZTa0Wi1BUMFCq4+ytdVpOzE0FGWtwuyrtgwIzYBDnTrrBRkYXW/A/p/Tk/HEJLkXoLbp686dk
0obAF3o5czqjh6FQrXv5uAgtoXEezAWUJ0L7BBcpeeZL6hogXNx8P0eQRT5lknSJ5EgqANxExK9p
zW5WFg+0WiqARizfIcrr23xGwviCgjVqJU+xbrE8iDY2CQKGoaPLD33Cq12/quV1UUhgdoFCi14m
O5F0jngjJjhuvme7KyCraFV8t37yNSQ/w3m4KIrMW/UxduCcLmSJW2Xn6/0Dr/Ow35RTDsdGfZe7
ToYDEdTZX0prdyTxt48TLFjBSoEyT0C85vvU74f86qm4rediycXM7zhO/1zkrjK8w4ageFOaofbf
2hg0PWJMRIMh8EjrYudpuJ9p3IcaFjPN4f9cT7F3VS4MFtNeugM+g2F5nXGFO8p3ROAB8x8dP2w5
+HaxYbj/PRpv2mDDPyY2Ttrqj4AKvIxCy47p7IodS7Q6BID/FS8cxtWbkuulcVU0Awd17oDMYSl5
l+JL5Ce7pyRflyxKI1Xk019bVHHgO8JZFGwypy+ODLwPwPrk1sp13zur/o2bP46ELkGOatk50YJd
2B6ksq9fcwaI4in8ly/4q8kIC6sjn9kTOpTbNtbTaiWcGyY1UeQZEOGfEmVcLYMFX5zw7lZyPkOn
Jhfg6AjPgylScfF+mMA6RJz34lLglxG0wOTXVjhVraimHahyGIW9NNStuAgcGzkvpKt6KwmhvE/V
4Vb693cxvqiB8slw+wvbH2Npo3MZTAAWdzXPazuQEHN2xOBwvSOkvBMRDnWhSfAaQev0HywYOZ55
gJYDH/aF0UaSGXXaGGkVF9HeSSVpx4zWg/VLjvbRBsdtTuEiYwumhEQAG/3MnrZsj4cc0U73vu2k
sBpuClee84XbSakji638iM2tW4Vpmb9VDqHArcLi+P+CTB30YqLbLCZlpbGlEPSrvyLwoqe15bj5
p887bLzZMuXO5D5XlZbPAWRrWX22RrXKYDOMq+cYr5MCBmywbc67t+Q313ZFMwNbhsRv9KCpuesR
Sq4PlXMUNvdHEoRVsp/gTnx6Pc9FC64A7ccnNrMDuES7A/8aRfLMBVCcRxAL/eHM7o0cWZks+jLG
qHrrmfBau7ZwL4+GxM9fXlziXmysvtBGPC2Sr6DkQU3wYIJJRf7XybIrWmrMYVwRYmcqgiUAYcd3
emwZfpbw+VVfczDY4wyhGJNlfy6k8X3dYwqwPqAyBTcpgISXtU/ekBUlFG3beX2qsUdal1DDQQDW
zhYsO9Ij+HvRHVQUiW1W5bKy+tlUt/QlauDttog4AsHyRUGZe1WBLi9LiFAY8qE9m9+gCXPybaAr
g/QFHHyfTp4RD9L866AbUnNYVKsYxYetUTzcERcpUiiOudzpKu5gCB2T+HazmG7/D+jJWj8ItZXv
Z4YWmssIM2/2SbXbG/nkswZR3Zu1JF+fO165e/4uGuBmhr4xDSkWBspqynRwc+WNU2j9UCvUogVb
bxdaeyrprbIqgQ/JfVq+vjKDoj1wGfdRjcJJoCDtMdrsYAc1wW+1luikF3y1VeuJgr0OBnA05IRi
gTpUn8i5htKmwSvNXgFlBCwq9bn+HnizUBPQgupltSyGsIu8k6ugq8geJVQentWkWYPc9uzh6Bjf
cRcdtscpbBHJkQuM3fasDFzgCCHeUGrAfGu0t7DxvyOwn995hhnT/50B774uwXOszQ8z0ISs3BDp
bScZGvV8XpoKx5nhMCwzpuS+AHLV+x6DL7MIp8v2qEBFku2V5r+fl0Co6/c1ZfMTJKZ064unKI0i
4a1Abz6kHUhYbc/yvE4dqbmwAay8qSdVYUparse84AS+n3mUEM39qnKmwq0TnFEnmxSzxvFTHds/
0DxvEfTuTZz6ikMLyY6A2ILw1lvmie24gvAdKjebYYOW2f9H1IST2UliGzGm7+QI70RG62NAZrQq
6zpQz/bH/wrw7XPTpG53gb/9C7sL9ejBmiMt86+dqbqzOlj1oUOR9uqEB9ISclLHv1HXBPJtDeZU
NP2QQa/KBCDN0MLl/F9+Cu+MmwWp3EB43cu+ryErYIVeftxDSszFPzP2X+7eBnxC66eYVdQK7p9S
b6ruB4sl5U0+N2IFO2BmeftzNkpfuPCaBKlUc/F/d/zzoRQGNp9V6F5gVHvKdEJncy0mlEO3GfCH
sFQUSV7ecaxS4HVyqGfs3PKOVbjI2+jfPzaFt/P2G5v1OScyllI8vo95lliw86fCSrTeHRQJ0uRG
Wq+SJkFpuPSLWnVQGljgP0ziqcRGU7PtO9yN1e0kewu5VND1zdV4I0Bfd7Fw1BCqvHnSsY98A+69
2ws500D0sLXZjNL/6UBn62zgMhb/QUh8qKkD8GcjWuglAXcCo8/KCO5ju5NkcgVHfa1bunK6v65b
wzlYIJGdqOausjfA3O77gJhB7BG+D4LI9HFkhUCs7SSvmmWBPbQ3Vatwsbf7Np16L1IUgZefLnWr
PMToZQfExV2C85PXMU3+eFG+O5+AS3vCeJV8Wnu2XDDaa1eAfPROxOB+54dWhh9OiyfKOyglHIML
cbEOsCwnjVTqYk/r6wOYvPmaId0OT53+JrgEqtnFo9/st6a+fnCtTX2TP6ymsnMyTG2XZxvfys4F
E8aXNklU66pQXg0ZR+Xvycm96nImeOntxxNC8Ou+mF1/QR+dxQGu+sIPDx9GHLq00GpeIQajZrcS
DmY8zd9i28/dzP16TyEfYSGTw1SnKDFTYBfX0gMVwnm6eXiCmdjSSLJmFRsVYpYACwrJohOE3ltz
tQzoIiSgBTwNnodOs9czD4vNM8lS4nlR6qSyj44wWRe4EkCgSkRluoRat/VmPjhH0i/z33MhSkce
AogjyCI3SulfQPwp2OEB3XJqztp+jg85bDwGmO2TzCQAyKrsZPDNEBWeBBdJdTlwEbNIYgfUIC3g
CVcBUi9TPjngaSQ98UpOtcAUsaqOmu/KvPYZN7YxBDmTV18/rNL8j/qxLpB0ZflPqLaOYwMee6mR
T57X3ovvbRSmreHBtZ6iMypdgrpkIWEmxTUCsTKsXHBpkIsCXqZUB0R2ZFvgJxTinqD+nwtk+I5n
dBDNMW0lqbmgbX6Cu/F6L+yuuKypdDnFkw3z1+rVHO28PutuMjBx1YZBe5TE6a0JC+rgeRsh/3bg
Emp/AIre6X4p3vsgpIoYBcnBRzA5odOm4qU3o5yfuQxBmP9x775x+alvWBZPOpvyVXEmWNLn0Msn
VygyujD25v8K4UO35/vCfaeyy9L4y5SV/vlN/EgeFiCYQUbPwkJEyJGJhBmR+9Y0Ro/RwAa2ALtz
Fstw4qf6BCE9zJ3mzF2uXDzsEQjgH0Xm8KgBZYTioor6T11NY5zBzKmLqejS27HSxROoMziLwu/W
Rkr+gnUcnwkmtpVIQ1pCu5WIDmI/8FiDjvuLBzagsySS6f+sVSLu3kdG/cjj4w+PsqzIpKDbCSQe
9pdIhYeG77b4qxnqX61XAZhlnXnlBnpqBcJ5TQU4aEqbK1lyKTFsGNeJXVRsm81RNoZgB0hIi9gx
tD8HefafFuWkM1mwOdxKB5pxtjBzFZCvTvP0X9W20e07TOrbCHc3dJMWAsa1/Sp+diec1QHnJqxm
R0JEypLWdd53RFqaw2e+hz1l4diJRDEpEZwpllCl4dCHs/bF6n76SKvCyX++v9mwGs3uO69yfpSI
5U7BON72jZfSf9JofE5mzjO8+ZZ7gHxvGYkzV6CjXT01rev5l3lxOc7JQcOQ1Hu45BqV/h5SPdNv
izNdiiNsZnvBVcm4JC7glDx0mU3vaflh225cs6D2SPXQcfGrZFRKh0TtWIPx61M1+sO77hZhlnyB
qu8pAAf1dNoXGs5FUUv2dGUOCWb7zK6dnK2ekiT0pyZHEhM+sAY6+W1vtlXzFFbaNEOpH9ZCVzVy
vkqfwmlc70n4PF6VR1f1mj3IuW1lDRz/XXmgqC4EQVPVXbUHWUHaI1tKsMim1Wv8PFz/L62O78eu
sQ1eVxIbVfIMlIvXlxx5aFTLagl/7bhXf6xXQ84v40tVC7nHUXV0Yot8u/F6DD2MLgBBixK+458f
g0OAL4EcW1EDGH1UtJiEHciiuP9j2WeRzSZMrrGJ7fT1j62pWT2ytMV4cE4HChoVjv7AodgbNx6w
Oq1l2gmvRVk2Dz+LYaUdX1xuYKiDhILWlDV/GxHwB5/GQCs/F5nLzmrCgC4CPknas9S/d67M6Cdn
MfAJOBjMp+OouGygGZFPXqYJvuFoXZM+hbYg9mD1h2ruK2NfJr3Bi0DfBwECtRljUYpSJpFFwYMU
gHnd+bYskryFWOZkr0pKSOIKPM/BPErUtNsipelbyNYHEQ1iSgaTYnbnITd/w88FNhxkwEk8ljE8
/YKTXH61jXeXHYmz8gr7HRF9Y1Ftieg8oGivFCyzNR5ySi8+uUtFjib+LAK9HCH5hQuKg8jB6PgT
MTE5JjsXXlvUauXRzDepUw/aoG3775yBBJiHDnQOqeFtwhT+FdRJ0PVOPg5F/0nVqcM44NR78vlf
EpSE9QEZJuvuNzc5L8m0CBU+ex5Id8dbjlCKPNvendtzcCaw9isdWg+uDQdD+RJqLNabkaygXBOi
bqJgZKf53Ylld8Teo0HlGpkPStRUbQv6FD6FG+WfWpmaWSY5lXCv1puad4D4g6eHnJOsODlU7ppW
WrpD2ueVwybE3JPPET0dj6kyOYgvih5c1DhY9PouY/JyrMojo1vZE0dtOP/78n0ROa5Nei+Cf9eg
30/QdjGWGOBEgp5s/HKupNZiRp2WrCUdQX68FtX3lcp/FnlXXGAwfF54m1821OU6HZDPFbVIzlk0
3yHh9Mo9DJ8esY8T1G7SjcPllIZTPjUWTh0y6qp09TQ/sdVptl7/gNUwuh+CiGuMaeKdpErUvKqx
wmLWykYH5pTSvXjYfEbeIO/T0PCPGnTty9Y8vMbgCZ4BRXiE2QVAo4iVsdMsCbJI4BSLm0/BorYG
rJ5o9KREkaXfh7fXc7RqZB9T82ecYZpTNR4i2gxFzUpXCyZJBbgHFex35EcXL8MYdF0SnvK6kcS1
PhyAvdZZdnMENAnSMfjjcHTI1Lq2NtFaNC/P4xPoaf9p+pi1/cigrLpgGXrtwDW4WFgTgrlnDVL2
W8I+qoXP9x6Bkkd5T64I+L+rGQPubK12b4NjYaFuOnqo3vqh4P2HIjSi10PNe3jw0CqmNdNHbmm/
W1yAB7fNUsLyr9o3GofWY4hFD5dbZy5CLNE9Y9S1bpIfZqzW2zq+AzdQypY3z3Gbr1K1N8xrflpt
AMt2NLsoT1jg+jJWf8nfcfka6sMkc0W4KC7V3gknBchLhat2tcTJ+ZkDs+NSc3+XTOR1R8pFNbAL
5rJkmGEI0IUMv0wtQt5Dbp3+uG9iBIIgGjz+6cwBcWRBrmp6s01Mcz74qj9hL+0stJnVQmdnUnR0
y5uIQ93pH2gTXiZdvAo0ajnTyo6PDty6dF9DVzQ8NzHTpwhPzADGrjjxB7bcJfhUS04wp1CGnKEG
0FiCtc0nfTzZzrS7p4XHYmlYkcZR6BndoNBxJh7GtFy2E+rhOVpcwoB1f2wMGsuDmC17H38wqyzl
jKtpjphy2fuGWaHRWgyjUf9xla0vTJqJGtutT6p/ZXOQd+s8esgy7TmKOLjeBckuHeqhMHeyl5gD
Fr8GGioYipHpmYIWZg5HrduKZdJh8N9hxiZkEwkXziO+sSMJTY16bFRgS6jSyuNox+K/syJq8I7O
yvRBgGiCQvMgvI6kpNMvbOTh7C8WtV+2sVFBlzYr9HOLqNSM3OUqeTrAy08Rp3fx8TVxjPAXud/3
XM2g41JMzGs8kloq6m0Xwr1XGa0fc0qM/AapJNpCpfikAMoU6p4+bmrXFa7+uEoDt3WBX3ozbSp0
LNujargLIoP+K4RijpUwZ53t76U/PQ8mvszLs5LFyIgxG9rFZ3ZCR51xysnf6ai7Pz8HizJDScvz
h1rAk0lN/6wMtqTgEjCeB08Pm++Tw3IjcrwRVQOJK06eBsC7fjQFxNuuE2jOuGT1/JTHL+Oimtp+
hLahuIBt7Oti0cFZA1X/5dDQrgA83wObyG4Nj5VMzXfQAe9t3dfRybWy6bOzPQbjcnqvMFPSb6KE
wbXAvT2yr0IB9dxe/A1sgPaY9fVXzEdqX7DRppq04nVEDwb0saOCFw66FmRquZK2S0Fi3Z6Y6X7G
6p0O8MQuvlBTaaGR8ceAJgSq7Hfa29PbVe++9Z7PR3HBJ75I/RV/eXciBwifgxLCpOeoffdKEiNo
6x/Y9yiEoQeH9SmRScjlv9mfAcvu2XtBJqREDU20UPFgLZzo7Ij5QivOfgN3ceVzL1DvRK3Jw9S9
8vyfTr6T18iqMJM3Whf3mWIW4rPnkOftk18rn/kqffX7Ay+qtCMAa659Q6g3TTqMrTI6fPJr0N6i
VnDKKri9ag5gpl5yTbSKpRgolbuUQvMoWTpOksHQdNEi6zmuT42k0lCWWiUOPZ9s6POUgaAVfjew
JEs2oGtVlVCFy3sdankAJUNFGlTS1NIvFz8n1fT2s34qRGu6aFVqGUXxyKsKEdzcPk1kXXHbqr95
lPCYJPUfSFqfR/KQDvyRarmAe2mOg6wVbHYZqzgYSRSUoVyC4HbfCt/sNsy3fu2m1FaGOdtGVOx0
nOdUQKtz2voka0knzXYIcppelGbWO4AhoqDMRL7/4cHs/59QDFL3Gv6+GriXVSQL1S5LMTAgtIR8
N4w3Rt8hCM4GQEwQZMYWZQ2viKhqtVK1vc8nbs7eYNEl+hufpKEXQ4QzhIrarpCAsAseZpVt/vVG
v7cOzHZ++U7Nc6EoosIZp9K+PauiY+XWblcOX+NSJzTvtBWsOQXrWfu40G5HobYGHhQRNGzMx4+V
IZb7fjLtntWbTwHB2UKbHZkj2rjkIMFgEuoWl6YXT3+RvTSbVsjpCRyFAmRRpBy5YAcIoPmYthm9
GDu9pxEEgcKcOPEofb4lEoUQQRBfLevs8nxd5AcNApJZmK3Gr6671aUIvsFShrcJMKTOVSEJdnhv
K5q3yk0qmOK+How+RWDcDsUMfMrZ2HVMv07MkINjxRAhalG+NkIMPXzvEZ95OZVl9mnk5uDLKZkC
uw5VyZKL72AHXvEapxkgSj4hNSF5lWb4/7pVkCzdCXJKJMfZcnJUIfpAk6/Uclh5G73MJKe+ZxCa
O6C1N1N8Yz31PIEbPd6q7xNZWXvFM9pq+9kaIFxlQ/BZeI40u+UBPtBENL7lXqPdiyX/1k3D8XWI
ZZ8ZoPCSRLDhYI2fVYvU939F6yNSXL4/iwFFDOtsm8DB7QYcxYfWuSgwvJgkrew5V0WbcrfDRdAc
/5/fPqzo0WGvMyZItYYGTeqgQzNT3pODAp/izdaqRclT8ll55L8vJRoRi62k0aizf27gGT0TW5Sp
0IQJgBIHYT0vpYZEp8c9EaX/fUNVmEmPYoTg3U9W5sn8D1Szc5rzMAiXlg/b+yh630hfYR2oR6x2
MrKWjKlY372LtLvXi4XbiIKNTBysrNmntHqHJb2cEd5gEaWlX/nnNzIA0w7Jl42qbfBJbA46b74j
+GPht2qJFSqWNVEdCghVgIauXHhH4m0U++Zfqf1US/cXeOb57AmFygQSVbJzwpukrfZAdl+diWxZ
KZgg9ACmoLM7S/rf3AHlGK6wZ+i10U/Ovc38MWb/ho42MiJh6RCM64zQuW+XRuC6Qu3biW9CXZrz
FY384yxfqikT9HmP45jggNvayqZhm12Wohrj5hN0qEB0kas4oGlDwx2YlxWPGxg6tzDEzWn84Zhq
WLwzID6hxPvGEVw6RTurutywjTAHqyNGuS8CjUi9YoyiCwBgZBN4UeStp7brn+3zUElywPv5mTLi
jbTESHou317sWUmLpCXiewp7JY9m1kP7W2S/LiLs6YtwoP+WlWFmKzq+a9fyIzlb7H9iIeEICjGN
z86WPtw8BRPjqBWNbcJUQMHTw0UVhAz7XugJkWNDoK9nyk+Zbhh9GFmX2k6+1qEZ6rGpQMmq0tnR
85E9RZ4wQVLVz0C4KwQFGrtCuAuq29Z6189PAoa4fNhZFYsyAQYKyNLI/vAAk5HuMhx7ocTcVzx9
xMHtPpITMr/cRtU24iqefKVYeAxWFJYMnRTTbsDfxBavmi2KosiSlIjKc2JcMBiV7GF9nFkqNvN4
wv0OmU2nm8jgttYEDHKINseueSOSO37k0uKpxP276qiPQgklqackGhpILmVjjOFbwrP4ELnKP9FT
grByNowNspz4dLXN07jXVeMB9WFcHBcNwlf/yFKHdJKvzdZXqvxYpxrXi7F+c/WR5PUWbToo0Jwp
hrh9HD3mLM9XBp1Elryff6OZhVre1Lyr0QOumuwpyogfqcGNz37vuCk8490cOX8l6BK7ykWPEAjT
uMDaPBB6bNNRYyUjIrUW/Hz93bJ1JuXyr01fIx+eCmHTCIOuZsu07ZMNuVVjHqDzQ8YmdoknSe7i
WlOl2neCIa2yA69LaPsF9eqjzAmcB/COuoiXUO9xcuke7BBqfcceT+RgnFK2LrHJOhDfrSzzsnUb
SjtmkhGjG2fbgdL2nV3sgWeGpb60
`protect end_protected
