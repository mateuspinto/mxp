XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����F �VA�Ր ����3$��|�R.9G�ݳYbPe� �ﾗ�v�ȁu8�������zY�u�;o�UC�N:*�;�Zm���⍫g2��Lp�
�龕8���{II/����bZ���qC|�i]�N�Q�s�YX���ߏTY�������3���6��0�>���ǐa���6��[����nGB�(@vr�p\_:�0uq�e5�[����$ףi�3|El�#x�R�8�W�uD��8_B�&U�(��^�rZ���m:=GM�4lh���U�����(&{w-��#��Yafpo���YA�x�L92�ȿު�zR���.��"��^P�p�n�3z�\���e���[�EHx ��'�{�0q eq:D�	
[cAH����[�� �C]���]�����3ʺa�J�,�Y����Lx�]���l����z�CIʲ���"v�AVc�+ݖ�a��)g�ޒ"���Im�l[ )��K����񗜃 17\:������gn�z�+j#XE��cI(����ϋ�^�����BA�B��� S��y�`��G�ʔ~x꤫���+����=!��S�5�+q�2���b�2�@ˋtw�n��;Z�G�rH�9�a$*���47�^��Z�Ȍ��6S�w9���5y� ���^m��MZ��v�7��z<�3�N�eګS,�5<*zH"�\7��Fe7�=�:>� �|���F�T��X��ҵ� ^ wz�Y�cl�fqi�jl�[ms�6bŧ�U��yey��8�XlxVHYEB     400     1a0� �
���J_0�Z����צHj������m�K�m�`E�!ALt�k���t����f"�wT�)]�z�8D� �"�?�2h�ο�E��\�Lű�??j1ń��}���S�V�����i��M���؞�\��+��T�ox����<�س�2?k�E�J+��14��ߌldW��gۑ<�11V��v�*�����n�d�����PqIť 1EqMd8`J���{��@<����P&h3�:N�f�@UwZ��f�pD#��t]X�!ݴ!��r��\�����l��
/(Wy|I����k�&&�M`$�3җ�����v����yC]��(҇�;���n/��}����g�ɞN-).0L���g��j�?(g��r��X-��<t��>����v�a��lrW�XlxVHYEB     400      f0�.��i*1��0��X�)xg����C!�-@Y᫃��M�CA!�$~���~����߱��$W�Dm��Vj��KKE�6��3�֔��Vׄ���U[y,WN+9�M��c�$�^q$x[�x2,ݙ������%�&�Ŋ����Ez���~�M�-(k'J�<�WT��V	v�O{zoaȌ<�� �'���3A>m�1ؼ�A	̊����Il$MK/��~F�7�@���Oa���B�����}Eq�*.�bXlxVHYEB     400     180���j�>	�fp[��`��A��k��u��4�H��0��p$�/Ō`���z��=�܊�)�B�&��ξ�D�D�mx�l%��};E+ܾ;�f����bJ�r��
��Ϋ�%V��<TM;qr?�?u(`$?�n$	�7���s�(�g̫c�f��0?aސ8A,0*�t2�x�c��Z�Я�u��]5Bh��{�J
��,$�J�Y޸@>r?��pD}���y��{���^f]�vlY���T�m�����1Bأ��⪧��*d]�wߑ��
�-!ר_C�+��{%a��v�;l���p���i"\'܈ภ��R7	��G���q=�Э-�7�Fߗǧ�C N.���Pv�`!��{�?�RK)�M3�-��v\JXlxVHYEB     400     230�)����D¸��L����X����cȦ�!��5N����!qd/�A�Q��F�2D�m`㊑J�ud��*L�t��>�}d�ҷcѺ�Z��g���G�n�UW�3+�*,/���5b�(�w��W\9AQv�)f���$��+�j�&��<�>��p(��/���T\�۸�M����IC�7�"K7	e���@i������������Eq�m5�S������p�!�<��,/D܍��Cj�Tp��;������>���A������4��Y��CC�7�$"�����X��Ж�y���_����L�k"��7��*c�dޜ�� p�~#EG���g$F^X���(��,S�X��E����������|�6zK���W��L@Oň�;a<��e/m����E0��{PѕUR��l��S]�	,t�|��)�߹��P��Z��}"���VK���� �X�֜�`N8���	RA`�̛�I�e��vP�H�T�ag�BfP(O']&!\��G���a�҉��Ͳ��0��4�1!Vy#G>U�cXlxVHYEB     400     1c0qDZZ�`�wv���A]�j��kJ�>Ȧ_BÁ�Kk�����#����G��\����d�kY�:^W$AcE�E��m�h����*�M-�1C*��f$.�
�w���|Q���8���e�;q#_��;y[�[%`��7����s������O^,��B0���~Q,�?��@����^�m�zAx��������핾�ץүZ�{�os�;�C9��);D�!�U/G�%j�]���`!�I���M�e#���`��sJ,�#����К�>���߷�\qU}םղ��Y�`S8 A����d���pTl�"�_��y�Z6
@���Z3H��D�n<�����K��r��W���g����$��T�����|���R-pn�8'�+�~�Fd�tnwrL�#��K 1�o̓a�������Wqy�p�B����{̈́�s�N3���U��{XlxVHYEB     400     1a0�0��xK	 
]p�,q�VZ(�=De�ӀA�oR�������NO÷L�E��T�0��Iv��v��
4�eۙ��i'�6#�㻲�.jA/g�t�� �7ʰ�L�	���n ���SZ��\�@�É�;���������pAO���q�����ǠJ��S����*"�Y��j��t��9�m�qz�*�j`�	q�1�>� �v��zZ�����
�#����7��h��m�	N���-:�Wbsʹ3�N+){M���'&� y�A�c�a>��s5<B�4)�W@i�!�/1҂'o��Q�+� �1���vTE]�Lq���$i�$2�����Ro���v��B��T�9>�\�\�>��Txr����Bb�skX�Y�Y�C������I7tP���e=f���`@ڀj�@�U�V��XlxVHYEB     400     1a0$�=e4L<c�QW��u=e�Lf"�OS�� �=᥾@��%��:�C��2��4�4��2��G!hLrz#뛨���C�m��Z�=���Ս���O~�N��?��C�yF���6?ėF��T�����('�o����/�Mt �>LwLN�W gW�k��~w���C@��1ɪC�ulT�ݺ�}�-)ǍZ+vv�c��)�!�/4:���t�Z��bĤ�2�ֿ:�`h�������E@,������{��O��忽�Rh��>�FX��Ro�`$_x�ٻ�N���?Q)�2f�c�Z����aS�v;as�g�b���Qj2'���;W��:�n�7�������*ڬV���_� �*Z���U0�1aŇ�����%��T֠�ÕΎ��zt��#%8 ژ�π�X�XlxVHYEB     400     1b0Jm"�^.����7�)+O����2c���\�兡ro�~���z�ۿ�Q?�a�u�Z"�w�,���K��	�#d�MZ���J��X��W�m"��ǎ�n��OZNO�nl���+�X�d[|���)3(��?�	 :�����Y�K5��`x����%��a+��2K�1x铵�b��5��QV!qع����rT;�{����WS���?��칇��PJ�c&�=�@CRb]�;_���t��{xf�7e�m��;���{���2�׊[��%����0�����X�9	���:u?�G8�J`UϜ�:<^�6�����T���4
<����,{gGC�`���6Q��J�8"�j���\�3�͐c��'U]#���hV�����y5�L�C�V��K�Ն=+O��s7v[�8O��92�0XlxVHYEB     400     1e0Y���
6���>&0�!�p�E]�(]o���z��.f���Q�e��=z�c��ҏ�=�w1U� c/�b�����Ɇ[Tj�]�g �.��+[C� ��i���w���L>�҈�i�������^��2�~���%]N���B�(���bsB"~���O�;b����0~�T��x����#���ŜO\�����8�%Ȱ�C�Ä�tA�*�k��\(��M�u#����qi}>R%�
�+c�^�+����k��د#��ޥz^�x�%S{����@�@I0�y�vR,c�����ǱlT�s�k��+��^�쓹�4�7��?���V�j��t���� ��Nuq���`����՜��ZtZNBǱ���-I3Y�i}ڍ0Fz��w@�
>,]�צ�`%�l����j"]�E�I%�"�[�����:���Q�m��MO����g8�~�p�TɑH]yQ	��[�XlxVHYEB     400     170��$�P�S����q|�������Rσ��-e+��";�,�"�Ƕ���)IL�qu�q=��ՕO_/{���vs <�
���L��/�Lo��(=�S�_�e� ��T�53h��u(�ac��(���P�:������h\��]�x�cy�H�yn�#���'��X7�s8�"	e��Fm�Ι�)F���%�h��|E�P���rb���|u����#֠��aOB{��,�c�G���Ũ���ԥ��wk}�ɷ�� ���~;�]Ez�a���G��I�o���yO�m�j�U��/��|�2�/��-USŤC����ƲZ���Lnp�4��=��S���D�>�1�XS��X��������.��M7کXlxVHYEB     400     140�����U�/���=c��>�Y�\�Õ.��N.��h	�;���m�9镐���KW���V��F芹H�
�u��8a{=�22]jQCW~N��R�L�󖛂^6�o�ܩ��<!�&��b;���g�)΁��4Vʶ���]'*D��×�D��pBǾ��X���>�S鼷���#�h�3^)ޑ=݋�
:�,����>�ә)G�6��s������x�k��r9s�PR��-��XVW�����J��:��4Ck`ۧ���^4��_�d����W�s� F�4�\��/g.���bt7�{���!��s�u���XlxVHYEB     400     140i(Z�D;���B��j,G)�8&70��g�/ঙI�ʣ�Ks�9���&�X�}�F
���� q�I��tuZ���fC��j:y>`�H��(ي���s,���t���6
TҬd2�$%^yin��N�}�JCT���VZ���6�u4���ۗë[�qW����v˷�a��1m���o�=�R�Q�ˌ9V�|Ek|����XyB �@���8��̷!�Vr���ZQ�_��n��Ӑ�!�J�@�� �"!5�a>>���qˢ��G�֎QS����އ<����
a��o�\�A����q�Cؿ��F�㣅�XlxVHYEB     400     1803 ]�{�M�&��X���x��� �CK&6���|�����%�*��۽!֎[�	�\OF�tC�:Y
��:��byJ�m�.DU{7�u�p��#V�=��6;%W��̷��\g�W�������V�ؐ�s�vKd��?O�9��,�A�N��$�W��+?���1���1��$d��)�+�	�㑿��ӚT���f��Hb����n���{6���=�����d|��yg�"J�5�T�#��B"��t�~e	7O����"G�Ql^�ٍM�E}Y� ���eXw�Z�|m�/�M�*j��e�{�I�;A����~7#鵲9�<S�䪼�j�B}�gj<c�qSӆ�i��(��]�@�a�)呉���.�2�#eFIXlxVHYEB     400     180�N���P���}FiZFn�X�D��7JM�K~Eұ=�����\��C�~d�cƏ�cz�#�{�SX�2��#q�aal7�9Q1Vx�֐�koO{����-�yl2�������(�<�rR�B��K��m��C�yX�9	���t$0 1G����q�}yyG�P!�Z��s::Q��/�k��#,��_��?l�-�)=X�]Q�\-�׺b*�l��Q��g�){\�O'*�V�`H��#�B<�_5�6������>;�@`+����Y��\���(�sL�a�� ����v�S\j����9j��,�|RV�<������ھ���+%���÷�J�$�Y`�:f�o�	�k����q��H
����(`.H$�z���XlxVHYEB     400     180�ݘ�!D��::��5i��İ���,D8n*�+t����8�:�hcj�y2���%��	cu$vd5�1��E�z�����H�6��J��Fp��3%�}�C�����!	��+&�9"V����I�U��'@�8ʴPV�1.��h$�_or��x�>��~��6�K��)�)��I���b��qyA����6�v�ܧ���*6�l�-f:H�A��H��
�L�^�:�2��MU�6������({ٻ�OzB	%Ĩ�|K�����IZ�3�b�WM�[�q���T�TJ�P��Em��vԆN1U�Ć�o�@<v����;|�VL�M/�y�(��un����_�l�p�� �(�η���#���Kl�N���v�đ4�yo���Z�dK�XlxVHYEB     400     1a0zS 帻Z���6��b���Sφ�v_�����4侧d� ��D���f�yU4���?���S�1	�-{�����p�|>�.��\:2����o��Fj?�X�-}
�W����
�o�_��#ͬ'�}��[KL�X�ڂ���j�ƀ����y9�|�ƾPxdGb�I�����\�v&�!���*U��H)�`~�g&-��y$14����~ Q��;�Z��8{-ßkŦ��۟~�CV9���p���4Z��J��eV�7�?ˉ*������������Ks5$�Z�����)նQ��2��5&�m�A����ftA�y�^�+w��;RR�@�a���C��ye��hQCF���K��Lu�j��vAi��7�A2�͇���cr��H�g I_�ϟ�����Q����8ˋ�=:��%EXlxVHYEB     400     1a0��-�i��x��	z,�kDw'C�,>���������q��VA%�ǹ�U(V��^�ӯ/��%�2y"'�r|��w��B�c�*�j��n�AV,q8��������@Ҳ4��ْ�H����\x�U�P�������|���0 �5��Q������Ұ�hm�'`��{l��RA����Ʀ�xJ��Gl�p|��9����r���Zc����81�
�E��z����c��=[�3yvh?>E��m��$,du�bD�I�4 I�V�[7y�`����va�Ђ��[��{����Z���ף��;��P�~O���L��2һ�M�!�aTy#��S;K�F'����<��W�� ��¬�U@�)%�T�|]����?5�>t��_p������)�>���@q���h  2I3��1/��|65��� XlxVHYEB     22d     110�ߐ��}���=��G���X�QQR��T�9��ԛ��~��a`��?��j ��O	�2&�co�0oJ���
ù��u�A-�)�����|,�U��T�Q�T���~�0/w����(P���(�N����Ơ��\�C�����%X����\��
�/�ϧb����d�m��J��]F��H���,�)���@��`Dm�N�L<�P�\�F�%�+~�"׋(�ֳ��D��Zm�"��x�rAE�T��~0A)z8��;��['<l��؄��