`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12176)
`protect data_block
h1+jxv2mpx35U1DEDQ5W1w3QwSgyFYg5T7WR9rGy1vOZFZINlca2q2AfG/5M1GIRaUobV94pbrSR
rF0DZrZ0HIj6UOs8G3MCE9ntX1WPXS2G8pm2N722K5vHtfVZjpAvWXNeCBIpKidJRoQft8PNFEgU
mOQn0dhtDuLyu8F7eALj9gSNfQONAo6bSHOLmY/HpKbIYGZ/3YerdPPhOPLjXrfjvhLzBLHYYwPB
uJgdkpl8MyvuieQxtWG/CDevGRTY4m68OCjUduau8M5iX3/6KUpBCDkYFq+Jv7c5TGqwf+c5NiBV
bBuvh+Jy3p8SDc98Y4vUHr2kguvrpGTVzxGAS6HR2NIU8/eWMeUDiBav2BKuHoHrCvEWlyDf9KsV
/ullTnGY+AQzczrQJP7PlOmPq/+aA43zqSbY6njTiMdGDmLLOcSj3ItAtJB4X59fjYC9Su0cQTpp
JW/iGJvuzd8d6cZhHeWEv0jsX2L/OjV8cn+yS786BJWMSUTDGA44Ve8VTO88813GnOYy2F8TaO/6
RYMGg+EYlCnCA/z9YVoEWPV6b2HrVnp9FcgXCsEV0VNt3qTYkyYlxveoIu7XLMdvqhzPVchkuHXM
B5yKYcAwpBYExgzjxoERTGwDMHH0nSPbDuAVr3RVUw6KNmtdaXPn/nkehO4K5vP6KRMrWZAcMlH2
gSFRpBliApQJJCcxSBGSyLdDjtmoDW8xmK9kbi+fsI0zZhLOQsqY0BSIyDhgZ3lgDu5AkraDgqfk
mpFSkivJ1/Y4ENI0Wu+KJwZQVzGErJ6eDW3osyvVEkJGFxWxSRhw7KZ6XvDiTOfKzndaNF22EisU
I4NIzh9sCx3UYsyUIoK67YUVqAPd07mMjVnT9JDmU6PsEboQNmTkrYLZE/GM17hBFOZlApYiibP3
FbvfBOVfYkhy+18d7yqcmyMIPRm9I/7EN9GratwYa4ARSqRFYU3VqhEMaCqlpdEu1898UUMAYFGq
3a+YL1PqNcvBhtAFFwQ2ad7fDvtlANK/Y9xR9z1N5ogHhM4RII9p9WVVLc3i7PYd+TyhUlgrV/zn
r+m09XdDlkdxSU2E+yDsB3c6CrPmvfeWVwc+fT+GCybglMNxAasJbQE9rR0e6Ja7J9ZPA3X4ff/9
Ux1TQy41efvFzq4Kiw7oJ2OdLzCZ1Ps8j40wO/sDZp+ms+8HCn2aoSc6MHJLGtw5qJt2qPUBnt1k
o/lfmZdmqM1tFbZDmNubqm0rb4NnVKiI3wN0/7dcF+CAUDHdUIQEe81Kam7sg+U6qSw3sZd4UQZe
1Yb5rJD67VGjAip4pgLydEzqMQMWuQViyiPMf5XTZ7ovdSXgnlK+0niMgPeKH7i0gGzmfv8/8tQm
z/dpMn3N48uQxAbPuGJYtB1Zp96ORyqr2sHyc4aDmKf+pFnWVWVMHXmO9HDpoi4J5iefy9ZV8wo2
Y53Ip306ffe2EXDKpP2SUEEnzG79y3i2vP+qqc1cfcHXbc8cx/U6Ds3ZeBXPpMHnqeaAtLiH7HBw
T52n4fRmg5SsXA3/tTkzKuMMjQeXXuV0uGJuU9R7wHhEu+m4tJrfBrm9vWMgL1JaEyKyqp+Z1y8E
GQQI9C2p2FbU3ZXQchv3HNV3626NcJdvakI5d9A+Hs/4whT6gnwS48DV8OR0TiDshEt6IApmEgC5
8n/SESjf/ynahSxqMEOmynsfOtlb3QC5YDaScAYJs61AhKDeuVhEQKjtdTKzd3/4iRbpfyZ+3rHC
eZCs7C0SnOfQwCFIRuJDsIha48jeH1Kf/1Y8eoSoS1TMShwewyka2MoaV5dYSoo+zgVK03a6EGNz
P0Cir0PbDw+yarSRZkBGEWCzgi1Tb/dXtEhBJvp+X2dJG9PUAx2y0cDNAMhRf7Ji41Uqo57iXn3t
CA5C0qqIO4bDmBs/SdzyeEquPBGVmdLkKZL0xHYwoeqYC7WfG7pFh7ZZFBhvNLLtTUdgBE3ns0Bs
fmbkL1bQvOwqgVongpr+mVRFE7FhebyDSJYhr7nMa23WGPgbuzD/N+dGoyYF73XWIDqrtLi4YfoV
/lM5NxWJ1c7+REoa7g8YxhxRXavfWdXTAiggTV2R5kLISD+KFlFG+C3UW/LXERCtmsYZTCBaGJUX
kOBrLZ30a7MMBusnUgxLGaNMIwSBdfCskKJzRD0dQfrnYHLiumYx2+4oyEAzQsFRTcIgVzRnSTJ5
GDEoFLdCmTXsSzKEls1XyZBbs7KUP5UfaTqz4oPi7x3lXKqy4t+tXt1j7zHzee5zLLsWHqLxoTBl
n9Tn7Tol0zRJUMRz+xOdaEEdjiiosvSdz5yvZMxmWpNAt7rbxgK8anBkuUiGFp7iIdKcprlDeDQb
wAzvPfRecAvuUQVsUQeGOmh58O8wv2QF1RgHw2rTZ25mDS9shijOfkJnDcMkNa9q4M8cRWoeW8QW
ekB8nlIcwRzWEdpJfnGbzryt2nnungsf2SzKInmzmrPoaNYZ3IJu9KKKWDWmLds2EsvlsDW34c9r
bvTkc7MwccU9CIKdtlzDkhgkm+Vk0EIEiYSXqIYfoloJJa0gG3Rq5WYOEgm8TyX1Nt+PPGb8x1W2
d2sevhTYSb5kcKxBIhWBh4FjDgKJ1QeGPdT68Saw9JDica1EwqZIoXnN3ZLW9j7g5Bu6f/o3OL+D
S/bTWpq0LAS6vOvuGg/3KGkcXSwhqWCnzzBGSB9v15FoIiIaIGxYxWpzG8EhSIVLu+eobxGUjZ9C
ODV0fdTEaled+rfrl1yZY/dIpDkKik9mCQ4h2dg+9oznpBGOIiDqEDjK3EHjJTS7MckDCCpRMfaX
KTJ5zJiRaE4Qj2Jc34U1JdLu0ZKog9W4QxOySIRb3d0434zAsAbz6X3v7SZJHo48TD7R1wkPv4+h
YRVYmizhpMveRJ5GI7kSxzaCuBj6N8io4jcNXGOhvExFprjBX5xfyPj6SBjgcrzwPpgxNnA/c7q5
fpK1R0jU+/MAKaDY6e3ToX2thYvInUtIHeGSSjKnXEffwIp9l2PDS+r3qi1Wi6X0hR7cTx/iC+/F
zUhpJOtJX1QIVnrOh2WmFaMUsl4mB/UD6O/AtExwTq+tc4n4a8A4Acs/oOdKsDwshUpWcPRi/Gw0
pxj9Nrg4hfW4HiM7OOgccbmG1CrXmeCeCJuSlhBs7R3SZCE6A90NwQEU8/9VvGY/F72apR7L0LFh
mWRzs25CQoYPFUE6mVklVtrCQnsz1yKfc9yMBqN7QbzhKGrBgLsN/z7Rgvcb3IFKlMtu2f04XYBd
3XFGaCyDEcgkd1pAtX4ngNdGYHlk+JpHfbBygD3eOY0phTpNc0JewLV3EaUNC3tvTmeE+1+tqqzq
hb1ao0Ir53Q3J+uSa46wIZ1Fm/BNW54fx0WW27N8+PvN2LrrUvTUFbJpvDV/cQ/udy+Jc20xBinU
6AMI8aZSbY0SFkLreP/QaRU/4/YG4cdGw/zZjLXRNHr7+UfAms5GzuqeO6jevs0tbANide6aJG9X
OCMYv6+xcD+qyY1AauoluFIOM5lT4tOM3vdZa4flCxcqHfexOjWlrBwXRYaE0bH53mXGv7uoSQS/
vZWFfTh0Oii5MrMbIChQ9u9r1oH/ssI5Dd54UjVGVOBVg3nWKxfKaNAH+3etp4axj++rwbHW8ED9
z81DbC6krIQZaRyl6EllbM+5CGL3aDqwwepPn/MkDSZl8R1dhiy2I0K5aIFUZxUyzaDFtJ6HBwGv
mmoBrgAjp5NtxXqRLbjKfjPD3SW7xNGLL19svUz1TCqjKSdl8GdQXhgb2UFJJbzpaGReTdW8gOPU
rPoP0DjaazFIiDfVpR8cIhtQHXBu0QQSriS4ZgjoE6zulxZs8jPE/mu1pYzgxEQhHvXqu+FU43tZ
WtTK3IEVUWvM4L+KxXy538l5Dof2xBh2O04LsvyPVd7Y41iJVMnPlQlDo79w5zdmNXS1ylX29jRt
GCeS/l7xF/ls7KZpX+Qqtemi8AZ8FMhvDeWFmPWOix8/TFTr0/wJLUQd/ZO6FrlW4r077RbRqkGc
3bZ11wevnawrbIDQmanBajIEWIJGpWUXEYEDxz0M5beIlDef7gNus79FlGCo/dt2H4AiFiDpbOqZ
fnV42FW0SwrmOvF/UKiW6bxS//epTOKeNM0hBpwi0/N2Cf4qBKMvH+jCXYV6Kb66EUVd3E1ShTWi
4pO/PTbLQsOcJ7ha6QQQ01dpHG8D71gsf9on3TgNPAdj1N+B7ddkzdvV4H7wbOG4jwtO1Hc0wqP+
AMcBMAXfwJxkGigg7yboKCfs8a2Ivc2JH2XvCJkYc7AnvQva5kACzXEdpBgW+3V5ZNLHdexeL7/C
ACSoMnK9xilxv7D+spoE4OEeYJkPwVwtZCM5y8BwX1/DA8oi4dTP3pVv0AP1KCVRQXsushtYNB0z
eCke4reUAOYMHv9OIKCE93mHWKdzQoGu6LJbb0o1cyZ4l9J67LIhT/7bnUfW7hess0FnXQl3Eq6G
7gbxU88rqUqxkydx3xTT7BtTX38Zre/vGz5hdZ+iM5793EgITeGrU8mMHkBNl69PrRUMneZsKhd5
RhfDv2tYaPStFw+YSo7Ph6HOqU3IctThSwTHToFt/iV37dHZfxJedlRDhD6v4lta8QIJ4CycU8Uc
7FmeSRoqrnaWJdKaDT2VghuCgnzPNUVmnXLJJE/7VIALIuL0T5klZO2fCS3JQlyPF6wGar+9cPCT
ivo/6EHYjgIk6yjlLkyIB5OEPaZ1tQZ4jfHVVcs5VXTdme3t2DmHPxysjaYWJkwTOhSiiBMO1rgf
+XICfJwPgtCnB0ujXGLNWDd3ctNI50z5y942wkJIYA9ivSHTIVs5GRW5uGYkU65arH1G91DVFsV2
jyX/tv6bQGjMA24vQpjNHKeuYiOkIimLf28JrOBRaw9MOkXR/Djq/mVNAaDbocYIfM0a+R/PPRyQ
0VK0/ZiEG86K0AKcCcaqiRkoRc82yDxA8NJWJyXq/BC22dSfmE4OYLlsCP2KSSsC3Dcnd3FizC9u
t+8y6rlEyPHI2uJHY0tpg6zQ+vqfNVlrYwSUjozCUuxq/PqLGYbkYQ+InWp8mYBx4ay9E5R0lj8I
lLyQLpESmpvgsS3Xejv4VMURJMriw/KCtj9RLKtxnBkanv5MhR8LLls7Fk5ys+kCFQGFkWmSoX20
L7a6czn2wTaSf6cWLhXYIwsPV9uxD9B94qRyPw7vrS1DJ6RIGt+W19S7phYzmb82LKIwTBYZJ/dP
Yy5RpINoirIKe+X8zXRG7jwbwUIVzzQCI4ase8BSEajIf+DqzlPYkjIOi0P+dCT/GJk8MlMN+2SK
7Ucj7PH0i9oYs+8MK83bCxdla3DmxlNJBkFYp+cLO45wu3Iew4t+7yI0JYCY3DBZy1B9kAxqtQ65
9t845qn8zpXbMqPFVqqOfz/Y6XNDwQtYE8mhIwHfIlhNfsA7LkcZ5q3EzDzxuHd+t/tBACLpHRxX
4fNbn2AKdBYF6e2nSDpuV0/lt8yKmoXaWfRCzI0+zGCg0KmMpamPA1dct2CyxB5BVAwddfqvdieq
tTryDwdMxAIm5Z+f8JyHstuMpDs5uJpKawLeDQUR/ThPliaw0lt9aAQ6COLESLutCqra6abyxUz/
sKjzH9xPiOWKWBCW2ihLRNWC3jKxpIXMBbWqqj8HtvFFMYbCPUFIKG+b/IzN1+RPbxmDzcQbc2If
wG/T2b8RZhggl3x9Nxet+OjWntVqo3bAPc5M+BHOigqRx38Yu7uFu0ViKDJbwNA7qyq0kRI8WH5y
HZ27SRjvkeFodud5wcm35BzXaxD67lmBoykTeiXXCZklUX3PosknGet6OY64u9Run72Ep6LO71mW
D4CI4cFR99GgjoRs7gO6dni0osTA/aMjrZCESg7jlChdJNwUcyPJvtXAhxCbKkTTlYWyNCyFVU6G
bTCPYXMAGBg2LHhGu7QkYwZ8Y4N7q/kj6150MRPLoO2BreOvHUZVainRjV59ILgkxr1QFrJ5txCw
HO5sJfCIn58Be+r6j5JDVSX63dcFwrvvQAcG8gxv6UTN/ulma/rVsGFS5LfLarrhxFoJi2GQJyD3
1QSNY32lPgoefWRLNGQ7aRmZKupQq/66dU7g6Kmk8Z/MHqx9g4Wm1/0gXcoNIeJCW0IZ1Tafvd19
+W3PfbotsKz6ky0ugYK+ZGmsJeNuTk2SdKHIZFJnrakdPdOrEiK/Sp91EuZJKel0WwHyU/rk9U0i
eh6cop26e1X412BigJz5bt6ofqh/ipPY4KQDu0uTqU/DIONK9/sFcO1KLlUK+rVk4cdy3uD/Exbp
UagtUzJ9qJC3ZvXyjim6bVyVO8u2kOCRL8XOTzvmKrRtq21LHe86+kAJ5dVIE11jer53wt7+PfAJ
FtifgXp2UJJC+rOdSq0O/uxWAdxZKKUw9wsb098hmUwg3bK5uwalF64hjy1GflO1xoPlTCll5WFc
Qt4P3IJjtkQvCwXBm4D//Kzf1X+LvAL6w7F2JwQcpe9YXx3NiseYQ5CNOuK4cuIHh7Vfz/L1tC8w
wVOCxT6ausGkWJ6TMlwz8guzH64Zff9OXYEOiQWWXhMnSLJGGv48hLjjz01lZ2Nreg6Qc6igOtWC
0Erhep1rHyzmbNwdnookhaukEMDY7qNksL+3RChSEsEL1iyaS2hy0mH+vE9q8CjIQd1nE18+LQpx
V6tVe7+mmHXRUw5DzZZsexEuTDsp1BMbw6M9PiPWax/ZJd98lJri3XrJwVlbPGUj2k75GR0/u4w4
ZrHfOnYR7+5PGWlmgg7/L7Vo14Y10GnZG/labGsYNNstNNyOTb8rPF4lPDU+mc7kQ6dqAiEeyP60
GNxoJxh1ntjCNw0y1pDnlzlOdnBFMnEnPQFqHw/n25AliXDSPxZJFYESy28zRapc+fAYS1hMvo2a
DvoNHRdn5znAAmWFOcYUyf7KPoliSGEYcJQvljZgMp1Nigbb+HjUgs1e+TW43lheBwZiQHeyZ1/z
COCjM0IRt0LBQecE+2FMv2R9HW+RrVxxNvTSTZR5EeZDVW6bR2NEnQubnqdYsQSp6etIdrUFY+8X
s/iuCtWBLOOlsdKOQet581BFHY+V26zcHMawCdnaCUhpcmLADSd3PLxNYihRFntPsIeX69HLnRSt
atS/5/qked8ytKQLai0QMDMAYvFcRFmo97+TZk//1f0Fm6Ep+kqha51xa8Yh9H9WwI/mrevGNwO0
CPKEWrFAaCv+Eebd2ddUmj2nsZnuGt8JskuH0QFVH6pSUJAL5TSaE1xh5zJSEk3QxqyaxtXYIsFj
QDqxaO6xOFhBbn6rLEnWGd4mvwKgT3ED6tvnp2GF59VpJT8dXBRLP4aHR9O+TADaENs+Km4Dh/lF
EwYrZZQtYKZEw7K1Ax8ujFJnO2HcVkDJpbHGG1WL9xWm3eQoV3Bs9GBxE5HsDW1z80kKYUrSa0wB
bUAfO66Z3//fKp2h/CLQhBIP/IRmuktFURiW9G7bA46oS2CEQvGF/xRWWver6yE3umvsiYAtQAIL
HKao+nKOu6Xmw1FpQLj5ASFQfe4bby2pPXgTTfZOit1UKAp0d10WlOejuzP8dYoexS9Tgj+5IgZG
w6V5PSEGrhExNMzOwB3mTwWSvpBwHGzVnzuNwhtztQCDkmoVhrl8sJwBob5Vhx7WwHZXQhGcboVd
2ttDl3FU5+8lneT3XKjjDBaXIYeRix7lapjL+oWtv630tebmQCk7VGvha1gJXJ7MAENnqX3q1RtL
eVFSBoorX6whH0MnQXg5J2wXNrg4dyV/VrElw7MIvCAKQQGi8EbON23VY5y4QNXAZ7yEipFuwOUT
CRmtt7SEPF3BxmOI0HRv2I5EvbKsZTHsEGowngPbZZEXGBbteFy+sThFBEeyuUQtsrhq0bRFsgGe
adhpJ7FpjVN3aYZAyuSXY83hfypUFLIq2IuLkCI2i8kjsp2p9b7rl4rkS0vuxB/gN1DHlcbQpmRS
btkaKtErDbC475KTW/wl2l7A2vu1yyyqgqJjS6/JLNwL9VR0gW9Pc9/fi7rwIhB8n1FE5toSjnVl
7gint0Nv+uxtNkGAoaq0n/sXRZwoFKpjFGbpYjIH+R7aVSuEl2bz/2aCit32Pcvq0vxmmVdZf/PY
ytILxnPc7URWOE8QcZrrP7mcwg4t3/idpcy2MOW4HMkIOJrKt4cpc32BtFnOhEIUPYEhAl+5H1qi
bgma1oSQ5Ru1YcgLXNxI8n7V4zzvWgX7AsHeBDiJmhiHzUjtRAa4NgUfb/YPHP6h2sWcBvvoxFui
KJBdGu0XAHeERWDfgvJRon7FMIh9uN84ENEO5ohU1JTRhATV3oNHgr4GuAVBmxiJSxo6sLiBkxCg
DuVT+JveoId/6jsE5Xp7cKNCZsP+Hrn5w4H7DLQkbKLFDFAma/noHUzhV1Ia3pu7rgLAZYSqMO0o
hIYjSvI4rimR5f5M9+1EGi+OzBK7fcA+X4mi6xvE43S/f1XExC3NS3VO1BI9b5SLG+tP7g6IAdzN
lkF5XYZyG327a6hGBGXv10rt1Y6QIkR6WYXn782Lf8pUTfySDXVHG+Qlo3IiKo4WipO2a50Ilf6n
belgcFnLXA88RTRiDetSW2EDMfistkVYXKLKUs0+8ZkBFyIVVeUjK08aMwVG9W3hbELkLfMEcP3w
B8l99fzM5TCx3aKImIdqmdMBO2O+oZoEzB5ipMPGEoB1CxZ6SBd6VKB5KtlQfOQjkQm3k/+MK12Z
fb6N/aI5DBLhhqzRW1j9REZZLwI7EYlyjhSuL882p7Y/DZAd6egLmTvg5n6f3JRv0Xmqa3a8Bnvg
sY1ZP/jZV697oNH9cOQK8+dlB//XJjYBlHXjM1T2JZOKDezXDXkmNCVoEj6ltwYwMAJVNMCzxOEH
Y3hVciFo4xB84je+zzHbh2awGisPT7h0x6b1vhG0YYRsg7s9w2xsQrZNBRnXZEAvu01/i1qU248K
EdNUF+8LQd44+ioZKXOv4uD9vX56nWIql5drq1jo85nnOYF3bx7lhEbvVwKpK1eCsX2g3a6FcDy9
tPdNU07TZMuOB3C+LE96OQcSitJIhVxP0umWg8yPeLxEyk+ltXCtH3NJHZxtLJiZfNR9g0ebkMza
H1B7jZqvg3rGvYzk8lIxt9r4yrt6DliUwVhNpLAdL4SdVM7bGBKJITfveBtch5ADVMCU/PfE9qve
DR285MDDReU1f2OhcNaGAocyZMlZhucgZw9cCLpSsJA2D7cvLvuw4aQ7q1g1ngoFmkqe8QhbUE0q
faOLrA0x0bFnxtWOU6CvOqM9DKYWY6vHdvHaCZFoK5IVMC7g0XIDKstxML18uS4ByGBGPdLUTxdp
hMVumJURaIQYXs1Dj62qThVwJ0TRsF9xbdfdCvIJxwjWp3MGgYhvFrYbhcNYar65iLou9/COclc7
YfvRImQNlIkbSz4EdqkxEZILj8qgxHliBtyy+H0iAJyhXjepv7GdhZpz15NZ01bQo+wtEDrRi1q+
OjoCiseR2SEHF3eDzhG89l/lpdh1mOgEj/MqeXAfFpGEhszVC36tCGuK8UI4J7sj3KYjB01GrvCG
85mCulN51fpUSd9AT7H3QCDmMeFptCRfH6hCwnpg8vQOWmVBlirW7V0SA8Q2UrsHWg9r3dDFDPhT
79nFZOQ3/KI+aVXBWFNq+OlYBDicfUyvrCR7bR4xuMQxo0pHmeLE/0iCfATPg4nrwxUqznWq0ywr
WgaigbmpVOIukWQJGZafnFzWuZVzlI0VXYRRHUU4bpmmqWLxP190k1Vj/a3vH5e2WML70nyrui64
Np0QPjZt4IJXHuAebvyN6XM9DxiEpOrnrSPa8MF2qvVw9NNOfg/ZPczACmlGFYB08T+MgjZlzPhf
2+aA1UHQlN746w5mq1VENkoB4gNVln0ndC0SNmcw5LWurmG22tI1dDw6dnw3K5CcIk84jzAXZ/RY
fMgCbmCqPGXwe0WqhQ0SgS66MtIrQK0LgODNcS7lyta/725boAm4XPkxi4uwNIV4rUptkAK4zNqa
rNMCyIp48FjdQ1eo5vD8WBa9XcdvVcVtYKnyZUJJwTv7+D1tEhSfBXfQnljteKgoThS9EUk6R67g
cT0YHXvdsI8qhWoi8W0/jI5KaVkUSvcr5JaaojW40BJwEH4pnmiN1zc8nhILIq7f+dN/zjv0DinX
nQfYJ3ycYIVcm9iRf7VFXK7LfJlDDypRs2gGzVp4FUpY/CAJhgrtYzOq19cg1K6yt+L2nbtRgjmz
O57F4RCm5KS6dZGxS6a3h+Yg2kqzcrJVxMPP7/YD8igitXv9wSwj4chyrt9Pkr6muMSIJII+aVh1
W2C5Cs6IHaa5eFOrzgoAkBVAUMNTWFlbQWfGfxyB4/3peg1lWLHN3T+joSuN2PuKqxYPBBL3ynxg
Xev3qYOpuv+hbKa+UUrwOgFXBCwGYMdFBrwRBeQqGI8QQsS1/KNCAMrd1syhByHlRZmmtWmIH5NV
c2QZYi5l5LM27tjHhEFl8WPYiqaXZ7/K526UclxO0okeoZkG5WjuyhkSKy/TJgajDDv/lMpf9JzG
75Vzvt3tcqKqhJ+0kq9l0eYmVrHaoEo9v/dvDCvTE68OUd1ItA+8+FN1n2+3H8EIxe3biuPcHr/9
DlhSMRy/XfmMZ5+POQdUa78q7Si1Tsjk385adPuwTuWpQNQY1ULPvvHFty4uaEAUM2/65P3XM5Oh
AdzORE7wAhbhJLlpd/97R49e8AX9YPZTEZXF3yiYkbI8obZAxX46p6bukQCNpNO7RYvh2QGdTvDV
e2pS1ARq/ZFM1NKRPDeF0XR8ssn7czSzRHlY5AXpkBcdGsVhCE6Zqg5UZ9hXgYm7HkhaFkLALP/c
lgevjZjP3aY5TxwBVDFMbtmnn13ypytjLYx0hosOl9/BUZe2eEf45jWNpuz9U6uMtu0QCkttvrwe
mmxgKLXPEzO1iMmOXOq1BlrB3/2d9DXcXv1hsy8TrmB3GQ6ak9pvbImJTC3pGG1zb/N18lBieCNq
706OWU2W8SIyVTl0dztBMLdLXAFFRpgfZqG1y0PNCGfHDEIS+p8V7o/VBNo8z1FRTs9hOUbQ6iKF
j/7xqByKh/nVANinYg4ciStuwdJt1TpDaOcfW4QTYkDLP52ip6lgfeAYmOA/6SN6+JI5GtoFnGAa
zizDj1PRbf7QZ+DJMWZO9sLJip0+hX4NOKl1PTxZCoVemZR29CpzXDQjdv2qftPONCW0QKEqTz7r
hvHjO659rvZ+iLUiQ9/GJVBHTr5Bxfxg8cp/LBLjcwJzcsO/w4pAo3JajvuD3tBuh9vdQ7GWXtQt
xwyZJcrRKxDuNA9LyWdWOi6+YIUIMcyI5iRF+Qd5qLSSaq3ZeawqeUDbzVyqTaXnzCAqC9ANKDwz
7JWzHIztgpw5O6ifDe5hfJheh8Xort4ymkFyhipaQnN7pON17jJsP4Ju+jG3qLq1Fs2nLS/DN57z
+2dXhInEyx1bYadrPo7t/Q1BVrl/MpOnOAphtOq5EDA7v1B5A+sj8U5F9zmfll6HiArzNQsqPWuG
ghFX0Zqh+FyQ8K4YKwlEiXXeMWhjsJt9pP4P4Ec6y0c4H6DULNiqOIa38pormQOKZkL0jy+l8Q8g
ScUX4RfzCuLYWEQhE9t/5C+dKkOgvHXdudpWbfrZhnF/BYyZo4eFkkYuihIg5OOoGJvyFYNlY3OP
ir4Aru1ic7I13/1BsniQ3crKoHZ3ui9K+6jiu8m2OXLY6YLsRv7ZIHeoB8N6DZ2zCdlA39STGrOk
4qc0dTpFB86VqTp4kwK6VoqCGVbtT+xeqLe64U5UvD9VxFn6CL2z1HlAzxTsUyaP9vS0B4g2efX2
P1qz6YQW2hg3g4p0KjTtU53UtFMEPb2gVnnlK4hwCjdlqR8nqY33VB3sghJ7nE9ztAeqUJ5ZV4DP
G2X3iGy9O8ZJxHXHM1l64pLzZpzBQZR0807zDZLIwMwtSSZBWI0vsoSoUl4P9Ol0199Nosz4eepk
1naqBO/kC/ElGxYWvk9d6RNyWi1ljMbNy9KXdGLJPmjeCbk22tJWuqZqKRFDj73jnr5VaUSl0tBO
/ZT4kaHBSTtiX0QonOt/zjTw/29ST87aLN5Uf9lCDoYZmDsZKSIe0AECBvntbbVNe8q0B01qCdtB
MK9KvcULnsz22rpVM3hvOT/kyH0y9+TJ1qsdLqjU4AQZMHrxN+CddpnNe5fZTYIQu5MaA+jxhqH9
xYQYiQqVDTaUdFq+Lth5c6RqHxEF3N8A6aATOnNbibEgZxEpPM13kI7sKsPAZW/y+M19fMxhw5B/
V6y0wkd83mxXZShNsdihJAwTprMyKwYp+mNiHsUalpofXvZ2rnNg33CjKIimi5Fy6kF+6qBaFshp
+hfullwDdES3qk6zdnJDeadOKg/KF6Y70hLsUw+yhNvTyfpyHsrsAFGrVZoO4ivcNhqCa+ivNHcz
qQjIzUwfGbdaPn9cvQt3A1HZBTG8E32fNHZAEoEt6xALuUmyhLsq+3xUKn1PILlHbGhFoNhO3NAo
9VbdJUXKXbIP4Jqw0cRkMdeR84Yeya59mUW2cRYAXiK3AHrTppQTFH6wfFxqED+wTuG+jyKt/IEy
fMXN+CndkO8Rs7bVg/ILXXnKhz/RmKIvc+jA9UwHFeiChb/UOJkCWi00J6E455kxlSOLYTx0agFZ
JSzB13UYQLO8xdzEfxIMWgr0GGOuyxVF0bsAjFOmyhbuHsBhIWJLS7PfQ7B9lODIJuORrhycsCDv
ekd5pcM14wKNkJfmDzmUtaZy3YJwm45aXZoycbOljKKsGxHUlaJeZVt2tq56P6rqR26Cg0Os4Pnv
Wrw2FoVSYC14LmzZHQbn/OUScp0UQz1o9ENpe21s4ilDd3wITKqrjMGtfV67ddYR80qVoltTgpSf
AaIB15tDbe/568qSPups0rZTzbIVqmerXDP4jvd8ALx0yZ0Bj04LNF8KS25pmYecgLlGUQEYfSlM
5TM7PwVir0GOv9UZeBique7CWbRI8jF92d0yCxWmKLCeNQEB4QZxfy3GLYycgyB2Kde9A1+mGec2
6UcHlRnllZ4BQNW8co8858v2eTJHEEvBCuqdjnuO03cmlga1xreTlErSjsHGfx3p90G3wF59nXWX
f+nkpdkWuj/1IUlqXrJGifoBF5u8vho6hoLippMKpj/ImdFnz0ACSBryqAXz0Qe9Rk0SYPSroMfM
BRI87E6sIDm2Q4m1EaSgYsTBYBKS9uIMDMI/TW9t6+iepzDc09vi9TW3y+ZtiRldhTibRWnq+4Lk
ZG2pemV75H5btTm/id1BrnrV7Pglpv7ox81/ZUcMbgf3Q9JNWJOkhxh+LQCBKYerJK0dcdeHUij7
E7B9sstkfvyLLiqRA+npbwj/QbAnmz/8qYTgv0pnmSTbp/BxB1ZM+p/NkPcLzhy9Wfg3/6ykk11a
GHqv9aMJbU04+rN36iOKQUgYymvOEIO0lFHko10CmooxyYDPD4m+OfXqvboyliCxOKhun81heerE
uLTKTdR8sv1dXTyI+4PIX/qFVxvrBmCoe/ngDEFJwlddlx1yeqyiU2X3DCsgxgS4tn6rQe6Uuw7r
2TPHzYaS1y3533zqnaAgcFikrsGiRcXGkwyWr2C4Ye+0MJwmotHDJ0+yJRK38Y04T1+TZU/9Uk/M
zUdEFgVAApSmEdne2EHk+yJ3Zcd2N32uBdFs6GqpDkucvymPBPO+mCc5CR4epSSKQHwftILsz64V
naR0IVowrx44ZV97HFyfdSzkCrKGKUsrQt1a29zsEe27xv//kYQ6gAtqWSvtfN1Ady94dhFDywEQ
a5D/xqgCUVepgoriuGjk5lbEDRKvZUKYA7lNMi4e7r1Fmzp1r8Pding8PK2xvL5KEDmS11lVSwgE
MErB0oV4dhonW6USYzpqIJhru3vZ10Jt28i2LD9Nt440wsYhVjA6pQM6CaGKr2dOWZidriW4nziF
uvMn6n9EFQwcKDvhV4cBH7qSqKIf3N4ci7jQvJpQX5QYqbs8ZW1NLrTqziLEF84QeqiL56u5zis8
fJFPdleuARZKp1WaffxNNraURKUC8fU+5TxT6BYuQYnEL8xl4GDvhwcTp6IIacPTG56SPufPWzuu
YFPfvBX5aKfsBCuRvootkfDBUqwfKPIYocJT6zM7bbJSlYwRFiWFNeeYq8esse5tfihwAsu81/wF
xCm7USPSA9BKN3qS5Yf12EGTFmviZ/g8qzdslrGSjZoTyXS0D7YvMlTiV8NSRUpDamBaL6dxRGL4
DouYMteuGkPUvM4uNRuocz4F+1ec93bPY2UF++Xmrwu1W1U2yeyzhcSNGrkf117CPWtFuixchEks
wQvoGDyEzcUIyxA2L87tXWr1aL0O3Rj+yqELdk87MCbuKKCJ6us9neFvDcYJbIIm9J50fByitGzj
SObKaGJ0lYxeon42vw4eVX9dU8sNITx/BB7YZ8jUJzsVBlZxgLjq3qJtPCUMjgkgvzgcfGRJU7FW
YLUWqfET2w88VMZrYYueMQarBv0MYgKWv+tD1X2mYg6XMxRver4bRXPj44azeTuJm2byOZRFY3Ju
ruO4le41mhec6gKJmvOIRlQAaslI8IfS49MRMk/fkx/HU/YZwJllVa/8E3QMgkNSKv2EYPDOkJ7C
KaaSldrxp9xAAyeSqy9CL6rTub+jzTRESKLXsKwApJBG+5aRBPfMd4+0gBF4kpkOgMBbq3sMxjpj
HMMgX2qKdLfQR4sf7b9M/gD1dgnoQIK2SNJcnm04nYpVP1l70T9MePYRnSZ3VHlsxoHM9mhUbPcV
ShYopCCYLRXCgQ3WZDcTMCBQkOI1+5s7OLUBPChj+mJobExX6kjNCxmiU2OYCBcBb6imUfrEzNfk
gzZDL3laAQczkhPYXFThN5TNt3dVymljBKbGoOsS5ZIHUxmEeE94AYzmCMZVLxf2YiuG6ggV1Dn5
XmMgE/70++hJUspVb+ss/ch9sLif/wsxfEwwe7ZULc8zkD57RbYqo0KrjtYzymN5i1fm8omzwvLq
pUWxfJJZUTxVaRMJ3AqE/NZ09ksyiu3QOqm8vDNjA+9PtJqChMCXCCxrdg8maEX0rYGxiDOk6svv
o3mv4Qgr7tkl6bMajMtxli1K7kZnxZg4Z/jIvOvc4pF1/MH3ay5H4+Xssuc4aRuu8Gk8lvr5l0x0
9kAFsjFF7BLimh3K6HsIGVB9J/VM5vZO+eqm7fmdaa3x0WX23vAWbnifSAU0H6w0u4l72S4iFlYl
efiOUXfBl7aF9hAey2oksHhNysduzgS/k80p5pn1FVC+n0LuY2nhNS9HJ2V8A/1pyEoOKfOjMoMH
sIZ58/dTfH/FKWVFzkplv6NaClxRwgblF/w3DvbYAiquD++YMmWtDvQ5VjIeRox6QiSUAVFRTInV
RPrluoeHR2hCuEXfuvgsFQvgN6aCEX0XrxfAiXbhp0EGyf3VebFbEY6YetJn2asq9ZHi2IA6ZjK9
ZxCpnKgT448IuWUEDpG6NkRZtLmKxb+d0jF6p122SfPP7sAbm+A5QVgbTJLNsD2lyA6By81BEXe2
9R39Ho/IpMRuc1kTu0AkTTu5s94NzsC9ESyL4bD+ECb5L2D5BHH2JmnJiz0KnzTM4Q4W7ZjMiuJZ
rZoYqAxRSvguMWwDkU/X5EqDSeAp6R9NOdgCy8/q7P7NhJz+5icOBGJ5CL1sDUdYc2NXBeE/kQCV
oTEP2IjBy6cGnUGlLBPRFTXhAbbOSoWM5Xy75JuYyhN7dMrOIB/JuR41bk8OJyOCxsixPYsVECVK
v2x6fNCxMUm2/RBnp50JJfPTnTVhFf9Cx5LQPRLvZAR/C74BQMkAz6u0Z5n9UPLgMgGL7UQ5Tw4L
wSi9RfQ+9i9BuOYqqaB72+SGSoFWIEWMQQEiuv4PH2ciykd4e5abbIBGDofk6A53Hw0c6Qx1uN8n
doNCzxR73cPfNn73JVhLE3spwZRNJHG6R1p8XDcDzMyHLT5VBMRFSRKeMT0IhuqMvW51Mu9wI4ty
t0kA/JQAmh9rccWK06p6Q/QPjlODt6AkaPVh0oIf42u8HC1px3+Nyl/uQ05+iDYPu5EeSrHasWop
l3ySegYdX12iEU42gexqDjkdp3TtBKY+BLVL/+OBhuKLDJf6pD5GuTb8qnMbz4vAb6MmtZfoxwDt
0NaSdUW85uhtnWa+LUxgC2Gm6HEUsSBt7jhZlZKsPeI2+6I=
`protect end_protected
