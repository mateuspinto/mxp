XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����>�����C�s��ic�\H�[2�p�	�;�,F�f(�eC�&���B����8m?xʑId�+�v�IcQ�`��%޹b��&�	3 ���!�:���eKoR{�G��6s�����pc��Ř}��Ҭ�6��D� >���m?�VO8�y��Y_������4]Ƙ(�;��K3%셏��qY������`\��??8>(mR^6�?���K�����>BmW J���A���ɠ��&�@�p����/kN�phӫb����9Q��C<6K�,�h�-?dEHf=2�ȕsG��!t3��YwE_�:�_��ꬲ�[L6,R���%��/�9�zY�"��Q{�O���
ɢ��R�y@L>	�=����#���q���Ϫoj)Fb[>n$ܢ�'���q,��(f��(�NL����6��L�ӈn�nx��#y�W�+�H��iq�7_�my����1깠�ѡw�$G����e���TEw=�_E �.�"Ohx�,=O��g#��x�'��w�Е��=�'�F�۳��SX�C���R1�Cjզ3��	��4��(T��C��ۿ!Ɋ��L��K���^L��LW���5� ^����W��M�7����x{�V��<�C�G���K�?�����7c���-���:�������-��#3��$�w�pJ��M��i7q]��yB���sh��o�*��Ȃ2ǹDZ/ O��y��d<��	��:�D�n�w���@>������I-@�F���XlxVHYEB     400     1d0ޘ�����=�g`΍��l"�k8|\s�:����3��u![jݛ�ޔ�+6`�$b�Ԕ���FC"��I@��+�MkG@�Of�qވa�G�oz�T�*q�A��zVTYo��C5��+l����N�̡�	}���p�Zj��=�fM�r^����e[��oF�B^ǽ95�Y�.��B���÷�=%�"5�تg�u6|:o~m:��}8[������	���հz}nK���_SRv�4-��g�Ws�A�J<XԤ&d'P�'�A�ʠ�D�ïu�P��n9oYhC���yF�1�]3A�h�7�"&̝�>O)��I��ej�p���I�:>yL	�~�e��A��H�Ds�.��N��=q��:��pO�}\�B_�5�58Y�7��u�&�Lр��ұ�L$���
�o�ݣ���W���LV�c$d �$/�~x3 ����@�=?/��28�Dl\���3�N�d?�;hEXlxVHYEB     400     140*mpkd�ވX�a�V�6B�p��,��IG�(n�~؎�{e><�S�ՙ�N�T�Q"�c�	w�A'F�눕��x�}�^�lbFx�G����:&��VX�aj�
��ys.C���È�^��)������5+���b]��31n(��ijd����n�R/�_�K�vT���Mt�&������[qdX$�e1�wG�?�/�x9���P�����Rm��O�"�M�����!��;��g�D�
�WҎ	џHNrV���3$��&�[^�,l"0]���NyMAuiu{�_���/���D���z��w �ɍ��43�XlxVHYEB     400     180F!���ͬz��~����Zy�i�d��w��K�~����^��ڻ�;�¸Ų�|�}Zy�����rrLa�#�c������r>������j%��ڭѠ��eg\�"~��i� ���7L|�LQ*r~��DSLң^���bG�z�6w�E>�B���ΊX������9˵�߇*~ͥ\A��lCt��)gq2��xk�
*���hk�z�-�(�E��U-��2,���!_g�rFr6%�*��P�y�rd�XU	m�X�6E��[�[��&uy6��u
��JȬ���� ��C�dI#[�{���R�A�4�& 2W��
��ubqF��E|ϙL8���G���w�Ɓ��Y>�ˏ������ٽo�v�H�H&|4E0��aXlxVHYEB     400     130hҜL��]U��F�k�l�3=�2�5h�<�C�;� )1B#>����-��*��˟��`��1���;R������iqNs�#��y����H���t�Ұ�qs2�.��-��[L���Ϧa���^�����Py����H�c�	dK��c��
��D�Aa��꥛�������_��I��/j!���7�O
�����I�z˷lVziK̊&D9�����/����+"6tfse�\���g�}����||p<����g�a�%�ƌ$�	ڙ�c��>�a�Z���og��fw��dU�XlxVHYEB     400     120@�y��#:��l�*���tҨu׍�8ruԺ�2��ᷧgSbޜc�	G����T���c�U~��8�|�Zƾ�p�@�cxn>ϴf�E�J���¸���e��A�׋n�����f��g�"!�x���H�p�<��{��f�`��mFs�ZG	1:�}�å�%��D��K�a:9S$��ؘi�H`���aiR� ���7�V��B
]����ja�0�QU|�x,��P3M#?���ɺ���R�g\&y���#9�՛��if?S�gm��u�.��^�}"/\wr'�i�M8�o��XlxVHYEB     400     100���sB�%�ﭻ,M�H�	�"��3���6!��k�#���H��w�_W�J�ݔ>�q`�߯*������Í���zx����w�b@2<Lv��;�+� 
�o�1���E
�^�e�:p��r��z�,�,X���cp� �:��i�u�H/��l��Nf`�?��hk��v�(i��Z�i*$~�����_i��gM���1/�kB��<�>���uZ�@D��S���������DT1P�H�����9`U���e�����Ҩ�B��XlxVHYEB     400     150�
KXڝ���_5�̾�l	W(y��%��?��"��w�-��4�'rQ6�_B�[\;��f�%��9s�s�-�gȞI~��� a P
C(�dQLP��4�������*��^�tg~nC����2��$��.M}��M���F�4'��)$@�t*�K.�E���9ֱ#��z��4�����D�nhj�a�8}8�T�;��䵺��aۿO��V�UQ�nA��|��.�y�2;_4ׯl��}c�1�;CÏKeU�W����]&��wM�\`�d
1�-�.�wW�[&s��bb�e����Y)Wud��2e�+2��^~���ݾ�;[��љ�-4�a��F�XlxVHYEB     400     130N�0���ד6��	�����E�耾��h��I2bF�^2M����;�u+#�_��O���2x�����P}�	s*� ^�|��IL�|���hh1H��B�'�)_!����|+ �#�o���5{@x^�2��L��Ν?��/�$#?�XM��<1��lAy��o�${B堹�%�����J�ǩ�uN$��C&`'0>�5�'
ϴҌ�Tm8��"��m~��0��}�FHH���O��y�����b�=7����o#����#�E��u^B9?Νn^�G�M������XlxVHYEB     400     150�i1Lty^�(�_B�����U�T��O˝��������Ya��^y˳V�]�<�>��'HMJLr��Ή�	�qm�\��O�j��,�/�7�9?���g4Ht-Y���dP:H���4�����>Y���*�'�&�D�TG��xs]9׭�/kq�mu��7���R3iǹ`�Q���;�ڝ������Y7�}�"����I|w�Ov_JP�} �8ys����[-�0��~	Z�h� ��Js%�)����#	a��d��3�&�pgS+s�R1��P�D�#5٫��,���d���Ʈk�RМ���g�̖5�],�
��v��1s��^��XlxVHYEB     400     120K�]u�8ø���\����ü)�v���>��W��[�ڄ�\��C�((���ЏB �6�����ȗW"�-�OR��q�:x2W�`H��W�Z�)|�}y�Z��������7�%��Ƴ�G�$��Ax�.Y�vY~�����U�p�^�� @�Ж=�?�r*[XZlS��5]k�zo�VQi[�"�B��"���>�G�.�7NŎ�֙���tZżN�{�P�h>˸��|&&�*��B�=2��`x-9��%��/��ԝ��fg�?�u^@�zKmI��X�elIXlxVHYEB     400      e0@�=\r�E�̉b���$ ����d��!?p3:��Џb�?xFBc��\P�F���>�}���&� �ҵE|+�^�/�I'�<�7�Ǥ��R��v4���(�[�(ziZmͦT��K��w�03��|��|S"Sm^�4}'� YFk8ہ3�f_�Kj}SWC�O4����X]�%�G�tU���	���i�	���+I@z�Z8����r@�r��Va۝ES�XlxVHYEB     400      e0�4��������CYȲU�#��M4{v��^���e=.�L�{���X
;x�p	kO9B�w��'��vF/U���(\n��}��%#� �'��r/�]>�i0��ԉ���zJ>�凇��c�+p���&{&���x1�.�%=1��]�G�A;�_L���Cp����������Ri�H &���i���EY�V���m�����z�^�v���KVQ�� qq�XlxVHYEB     400      e0�2��a�'\L�+����L�H^m��8�OT,1�Ӈe^���;;Z#��=W��A����j�n�.!�a�/�[�(y��t��5[2�z&� ��ټ�u��]�e�Z���%�ܷ�;���׾���Jl��{����u$��/��@� O��ɅU��y���/~��1�C�W:���� �)&^�vaW����'``�]�̌Q�B}�Gowo��7���h'Hk���XlxVHYEB     400      e0�y|H(�\�س�v=����~�0�y	���:m��<LC���dT�э�p4����/���CrpT$�Z�<&[,�o'��8b�/Mհ|�ڲ%����h��$w�V����W��m��o:k���@�m\� �y��a�0�,TX�(�3)>_������|ZR �8����і���_�uxR5~�	Z�L O�W�|̅ZB���8�'V�5�F<]�rO�XlxVHYEB     400      e05�7���g_�d8;��Y?F�����a�:AG��\KZ�����C^s_[Ϟ)��+s/.����YGm0+f�0�&�#(� {��'����/����n�Ggj�R�`���n��"a��!@�!1z�{�־����������㻁O�YdOm�,��t�Ȕgs�}�R����t���}�%����'�`�.�� Oۧ��m��K�3�G���}�`�XlxVHYEB     400      e0�%�s/X�E��lm'G��d��g$4�Q������N
��T�<���r�
� �`�Qd
��Qtnĳ>5��#����m�:�r��K.�ܯ�w�p�,�T��)�|�r��}�g����&B�U�+���h&���O��8��z
IQ,���h�r&����q	*�t�R�Cb
H���S��	k�9mn�7�M��6����P!�v�����ኚW{.��:q���zj� �XlxVHYEB     400     1b0pD�pz�g y���(	��>��x�����[�@������ף䀋�Yصpǘ�?�ʟ05%�EGEo��*v溿d��#�Y���А��%7k()�tu�~�ORv�m���zu<�����%�N��`�*9ASYi�<QV'���	���T�~H�:bsWYٵWe���p;����C�	Y	�׿4�m _�@z#�⠚7S<d���J�S��������V�L��ܯ����j�$rQJ�WHI&�C���Ed���ca);7��7%e��9�-W�?��'���q�f����s[�D� W�����t+ŦXXb.ė�b^ﶳY�m���%�Z'�y��#I3L#R)�(ܕ�;uc��,�����G��~��)Rt2���tF����c � B�7׵�O^�<�ׁ�G���R��ҪF:XlxVHYEB     400     170l�x%�eNA_�C������
i��,�V�6�N8�j�W�����{�Q_v�]���N)���zh�wߌX��J���2A�/h�j��J�q�G� �[j�$���ʹ<L$<��Y�(v�zH�&�ۧ�r��w��p4��it����/����ĉ4A�Z��ЁRUt�)�y��M�EZ�i���/�-��E.��TU��&�D�̃6�n0��<�6hjJ��6�Ƨ�@�s�&׊�u@�)��xeE�}���E�
��*��裉�������0����/J��X��ϣr=�cΰ<~���Y�h���~�Z\d�qn<"��q��h��LZ����,��xS"[p�tB.�gH���(���XlxVHYEB     400     140�*���7�80i'Qp�XL[y�aQ�8�(��(�V���Z�T�w؜�r�}��UU��Ջ��D(��t����%
�2Ð�V���l�+ޫ���l�p]�N{P�z,6�
���S������ꤘ�����VA�Ҙ;�� �@���-'�?]����3�6����>����j�Ŭ�6�]�>�x��K�U����p�jZ���2<�|�8�����\���D^�^���J{iÝ�o%�b�p3Ņ�/~�v�PӁ�2S�;Y��}����( .��{}�r[��%�k�:v����4PqF���:C�ZY��XlxVHYEB     400     120`���2l+�/�X��׵鍏�[m�� hD��`0c�a'�nhO���\�[����.mz���7{Z�ݡ����4PA�5���q��,�ʷT�u����4�V��<-���:,M����v���X�A��!�M��Y�@�`���K~���s��wܔBoD���Y���%�>�=v�R��M�;����;�`�8=���m��� ��<�st>�
'r[��ϥ��WL/�͉��G\���>��֥z�u-��7��?w�P�2�>8{����`���R/�����ٶ�i�XlxVHYEB     400     160U�����XJt>������a����fJ'��h�A��-W��+���b�T�)e�r�@CBv�8ia�_�l��)���G�(�o��^b���6�p��h;�!6�^�F#�~.Ce<N��fi�~t�qJw77�FK��X����h��,���w�fo�vcQ��~A���)ޟ0�>k�)��G�ʊټ��_�a�7d���2M��9k$N�+�����9����W�N�����$a���	dZ�j��(�x9
'�SF~F)�V0��7YQ	��q �g�`È^�]Ӛ��:C�}	���2u<��+$C �-�_�[�Ա� ��`�7[�������ZM$m./ج=� �,u��CXlxVHYEB     400     170��t����s�9����<nGhlH��"�w35@�դ�� �ƞ����<郖�,���i�U8���X�O���ޛ���*Y�&;��v;�UU�[��ͨ|�rQ�^�����:�W���(�����=T���9)�@
Ă}�:R9�E�fP5�lh�m��Y��N`�Iϯ�i��h�W�o��`�Bn	O��L{�q��I�R*g�F[�|�%���`�L��C�[px��gg�t��7w>���H<{��f��W���gɪ�n�5l��2dt��s���_D=AA��Y@f�<��8��QYdz���Eh�(���,Ȟv�$��_(p[eŰ�N�OD&5Nd�ҡ�r �}���!XlxVHYEB     400     110�C�x����β���x���,��XOd^�0D�����-i�7A�H��0OM�l���I"�]L��eut������ت�q,�KbE�� 8^˿lB�=4B�j�+���`{=��#0�~�� �}0U�3l�2��[@�Wd�O=�O� �s>�E ��uvד��~���OV�ԭ���jD�D�OG1���O�����!D_�ȹ_b�-g���^��}��4z��%l�4j�z�P��������6MwS�n�� @}t�ųXlxVHYEB     400     170dzy�(��#`��&�9}e��7��2�}T]ǧ 4B�\Zݗ�V����4k~cO���D^B�|XZԉ�3�����ق+�3VTr�a!�d�a��)�ј����u�j�>�w6�����]D$i��4��2�:�ݐ���Ğ���pI]��*��8�D�̙�\�[-(um@B�����$��5A, ��JK)1�:���ݙ�{{��]��w�W����&a0!���x�W���,�VF�C������PM�r�х�d�l�3��O���-�f%�,�hV?���q�^�~���h���*�C�T9~ �]ܥ2��5���SW^���9/b&����ޝ�bZ���o�x�
��z�?+l��j��Óo��T�aXlxVHYEB     400     180����w\�$Q�JuH�PL�� ?�e�x��S��u׭����%d�F��H��,�lV?ay��B	���S�U�x�v��d�e|iQ������u�����:�B�5z�)�/ܸ��t7$P_%�ǃ�3�Yz��40�m�)��౧1.�ޛsR�����p��3��6��zK:(�ρ~��!M�U���jB���í�JPҗ2 ؉� 8��]���#��K�Eg�!,{���_��v���3vk���e�� 2YW;��?�M�ئW1���.:A�GJd�d�cH�D�8*��fе�/zHh�Zit9�h;y��I
*�3ڰ�M߶Vo3�
��h�-�FTXR���w��>��|�ഝ���ݨ&C�Z'��rI�XlxVHYEB     400     130ƚ���_N�w837�X�{��3�|M_#DS?�|�?�%*6\31h��DP�ov�M�/y�T�gZ顱%˔#EL�p?�t,̹]ՐU���U8��mrq�G���Z�
�)m�&z$���z�Y~^�?���|�����wj]U���ָ���(�QZbo�v��D�Q�LN��θcC�Px�2`dm��G|\��@��
�ώ�9l}~�oe�$k�`4:Ivq�� Igb�"��/�����ϢI�J�6i���e�к��)���V���F;:0p��1;��v�"h��4��T$*"�XlxVHYEB     400     120�f�0÷����{.��Lp�&o@fK�W�S�Rӂ��䁡A�� TӄQ���ۉP*_�	�h}��V�`����;nWW0�]�-a� /�_~��E�yP����#4�h�I�%���f�Vlܥ�Gy��-*P����ka���c&�h�|��d��[��W�������؆��tj1�7��ɕ�9��Q1�~��y�����L-��\��rYғ7�r�n��h���e5�p|�p["(LrÓ�|�)B�J�Q(!݌��2�G:�:��a����%8XlxVHYEB     400     130V����ʭݖ��1'K��d�Y�DO��@�N�߂���E>�x��\�+�����i����k�@}�� ?�g0�}
Ɖ�ݙ���B"d�5ej\��n�;=r��g9E���\�*D������OO<I|����בx�r��~*W�=�$ƺ�E8`B]�0�߇p�9�.��z�=��%�̕i*�F}�9�b�� �k��({U&}ٿ�]�29f�+܇$�%'Eϟ�#K�M��%@(l�-��]��"A1����v��S�ASAh]	E�i��=��K�V)�I�<�3&@8��2Ԍ��9R�ǔXlxVHYEB     400     170Y��-U���Kq�M�M�t��}�aaMD>.��M�/'��g���WC\q.�����RS7�*���& ��]�ډ<j*$�Wy�4v�uh�+1ƒ���i>sT:{�^:�x~�:��8}©���s�qB�N%,���Q�f�"o,�ڝ�	�-ƨVˆtG����};XS����������7��|+Lh+`V��&x��+>�"&p3o崠Y�WXn<|�`��p
����HD�wޓ����.�l"����B(E�~lg�}�s��-�v�`���łί�~��K���Z Ԍt8��������q����J��I=��8)�U���12����^m �B����jE�p�������I��҂rzXlxVHYEB     400     180'p�EcC� Ű�zH���
󿣦aB�-��!�$��o�q��� �����B��[˦�<[�I�x���1���q��hMl�8�^�@�֙�3w�S}�ɗXD��nI)�pv��|q�m�(Y��� ���P��B"l=["� uđq���..p���F��$v���-�Ͷb��]*O0''�����[NJ�pU*���0=KvL��cU���Ͽ��f^:"��	 �g���p%�4�����̵��p��a��:�X+&��.�6��@�vH5�Ik�����tu���[$al�B�5{�ݫ�*'Զ�HsE�B+���A�
�-U��O�ʖV[$v����1?W�;경9��|d~��6�z��e�O<���B�"s��.�x�ܚ���;9uXlxVHYEB     400     140Un�(V��kE_���i 2��%��te835c���1�z���@)'q�|.>�щ�ٍց���.�c(ʺ����	|�pX|����u�?����m�Q���Z��biih�-%�e����yZ����Π\�g�[��+05�OT�4�
�ͣ?M����_u����{�a����m
���P�&F�$x�zz�ChJ�Ζ��J-|�/�{���+y4��$:����(�2  B*A�%�Pt�"�%�H�d�LL�YW�� �������_��[�-�1.n�G�v�����R�p�@����aE��y
XlxVHYEB     400     1002��'Z~��-�Ǥwd-J�8���&�|W(X���iKp;��"��?�j�]C�⅏<J�ǖh(��K(5I.<Cs��Tpu<�ln҈s�m�����[�.?	�S��gc{�)!=�Ƽߤ�t�N���b�MC��:�?g�KPꍠ�,uRJ�S�>u�;:�B��9�_g2r����v/?���������х�����Y�ԙd4ny���LWz^�� Nx^ؓ��b]g�G��1p9�#�1ϩ��u���\XlxVHYEB     400     150����`�͕d�$�.lJĉ8��>�a����n��d�N�#S�WF�l�(sy���B9�]��/����o<3~�#x�õJJ����c��?�	W�����:}CA��:���I�h�BZM���*eCᵏ{/,�c޻}-r5��/�Nr��$ ]'� up���v�J��jpG�&)x~	|��䶎� ���
�a���,��:_�+���� �5�4A���C�+�Վ:y�a59״G��Yר��.�3�S,DH�V<T�(x4|T܂K��@�s%ִP�%����zȶ���d����8564Zi���R���XlxVHYEB     400     140��(e<G}Y���H���V��=�;�_���d����H�h���E5�V����y���
ō}z����i�v:���pt������%���y�&U��m��jI�>���?ŧ��.B��<�n���`���"��>{��o?0(����m��e���&�:4���N��$<�xEG4�
���j�N��ȍ�V[%��ly�x�J���+��'Sb��B풓�����^���>��;�qq�����ўС�g�FvIb�Yk͞���O ��qAʩ^8������K���M��:�	x'Z:�/���j.�:FԀ�XlxVHYEB     400     170�)�4��J+�lYO<p�{  ��<��U�ea��|�"��b�Dja�8ֽL���v/0b{�/1K��<����h�!�˟O�-y�Ncz4���ӵaU��Wd^�'��$����?D�ζm,è>�9�����JX�xeh�����`U�@op.�K:�a6`�t�㕒����GY`��]E��?��M�[5:�ɮrv�'��m��>���~\�_��#�����'s���߰oE�'�@��L���4$�(Z�SP^,q����=�N�]UK=�הּ5���e�ˤ�! �הT�Lu�as��`w�XU�S?V�`�^�Qk�p�������Z��x���&�N;��1uWA4^AQ��%��J̯������XlxVHYEB     400     190�`��_�B)jPk]�vK��ʏ��;�+ҁ����@
G큈�d[;l�߭�� ����K"��}��iv�UЪ��[�z[�+X[v摴�h�7<�.)^�<4x��?h���߲�"�����G�8)j�k>�9$禕g�9Љ��9K��.��;e��:X�}�J)���L����X�b���5���^y��6�d�hqk�k�ciY��2��	=�#k":)P�ԸY�".�b��O]�,�SI.�ރD6,4���������A�~RǑ,%��9�6��g��߼�\Zswk9g���A�"6x�)�#����ViH�ӾT�x�BHb�o��(�@x���Œ/l�N�_���G�'� �$79�����ס�J�i��}�]�]���� y��w,�l�`�J��%,�XlxVHYEB     400     180���<���;G׬{���X �g�x㿻DRף�օf f�Gk�R�pc�vO�����8h���1�����?����.nl��
�C Q��S&�Vb7m#��.PZ7���wCEA������$"Y=W�5쬬#R�`���퀋K�x�Cĭs�FU�w��L?��A��4�'�j�h�e�ɥ/�o�>ZJ����������'�C�$wyhmC"��Ծ=A7����É��⩾����U���y2!v` YoI&;8��Ԣ���4e@�:��ܬ}�7�#x5k�)��L����f3��驈R�)�a�j��b��3ؤ<�'�:pi�~�CC�r�#��h�v��Eҿ.����A_ЖE�����w SEߍ�Ȍq]����W��XlxVHYEB     400     140����ْ#���}�%O�[ѭ���T5󰀫�zB������s?�}HZ�v��4�2n�����m�$�wC]�@ƒ�`H�ψ;z��<EF�Lz�H�%�����#/���
����quX4�H1�x��� K��ь쎰"�C�Ƙ�PXE�2����P��;�[�y,�f�n�&8�xși��v�=@g(����jy�}��d�u(-��'���E6�����;�yU�Qe!�\����҃QN��h�����L+�|R��I;:�}�����G�ؘ�X0�2��V��nf�Ō,<��5e8�������6m�����XlxVHYEB     400     160��kfv��q���^^%��+�|m�6pt8�Z.<�j��]�~�%V��1�(�1w�tc�f6$�d]�N��6��i��*|�"�s�0�ܭr?6���W}E��7��\N#��p�3G�)�:3US�I�J\��)����^u�K���df?���F��S����������:�)��T�ۜ�����*J�o��3W��	������6t� �����R"������?�;�j)�u	T�κ�����ޗ<���U��������	7W�h�G��'�"���6ݚqYަ��U@e���E=��ń��8Ƿ�9.���E8�gf���!�ER��� �`�:J�H"�w3���f��L��l��n�R�XlxVHYEB     400     150�� �J�1�
h��e���{͉��#KӉ�����B*)�>J����GG�ۿ^�y�1J�B~�\���o��e�ݷ�1��3�G2� 5� ��S1:%����*��d-="��핔��q0?��� �/��𛏞�L�����a#�/�V0��o�/�(6���I��qe����6�Wa��ù��\��9��<3ֽ�e�X�|*j��yJ���H�����"{�H�pC3�B&{o��
����\@s\R`��	�>��es&�{`���e,b��g۟�& [[��ꮢ�⟃3�@�]�G'G�h
���b R��mcdƊix���XlxVHYEB     400     180%F��q�MA��k~R}�/���"ʗ��j�t�'��_�g-�ʭfZ2eB���.�s#5we�[���S�b��?䄸u£r��"�n�z�(�e_9.B�� ��� o]C'Se��K@*�As=�����#k�q+�1<�8&��e�U����}#ع �1�/�����sz��1�]���!��x4e�^���P75X��*l�rl�tg�sYVŪ<�ΞB�ј������
Ð��"{�*o�s+h(�a}���	gh3�L-�
����zpn�q�1�w��^Ne(±��Y��$���Cz�h4��\N��4#P-8-n��]0��3[O�$lD�P����s�JG�R��C/����Z���Xqlc��*�.\c:c3�XlxVHYEB     400     110Gu�ht7
��͛�ܳh�42b{��HM��c�O7�,ajOzCL�o`6ʋ�p�6_o�A6��mu{�rv0n��k$�zt������:�F@���o:9)=IW�X��o%B�)|a��r��Т_�Տv0t7~m�gL��n�)HQS���5kb�t�(���'�l���Oŧ�Ύ2�vۏ�\�� �:��Av�@X�0�L��˘�H�n%��c"u6'��Qb�hw���j�
��W*	�]h�v{�q��9T���j�n�"%�),kE��XlxVHYEB     400     1a0RX[>����Y�U�Ր���ԕ���_���P���>��0�yx R�?ǡ��
����y����yh;v?W�G�$�!���!��tͷ.*�������!T#|��L_+�Pά��U{D@76��;�"��RY|F�t�f�f�7��
�� ��2!�g�f�?�_*# ���囗�wrd�fYD�'5���".G���ܔD鞚���4���$�:d���(��4������&q"��A�3o�w]�5d����N�m �eY�ԃ�}�j�q� 9� ���>k"귵Yc�_2/K0J.�8�Q�A������F�%
�~�,ex�lX�PZ���+]@�S�T��K���ͮ,i��1�F&[� ~�Ldl��rQ�ћt�=�k;d5N�R��~̍�3��Ύx�r XlxVHYEB     400     130������rw�f���������0���P����/8D
~z��_2��rh24�52Zu�8�^K!�[�������b����E�7����/��1���1	�C�@��?��7��ν��I3�mݸ��
��^����&.����:��E�
�(`�L$�k�@��������g&�O�������xq�+nΫ�Ml&��}m��
���_Zւæ;-ad����]e{��3�I�*��V%����y��p&;;+��q(�ڙE(�ʵV����G�s����B�h�ɲ�617*Qm�I�XlxVHYEB     400     170�
��w>�\�
=������A���n~臊�^��k<Aۃ3]͚��;?МTt�ޢ�G���P��IF	��Y<b�#f9�ED�\�gY�0S��j�8y��uKw�ݛ;
���hi��2� i{,�em��z)��eGj�&�Z;A�4�����u�t�t"��(�r�Z}�^/�ʾoL�F��M;uߐ"�ڊ,KӖj�ge�$o�I�jq�vd�=X^)F�t��@���/���a�VŘ`�YB9�^��;����XxdUK�k�ư�[6M���؟q��"/��H�;��?3��Ϟ�ɱs� �����m�ߧ���_VR�v>�j�:Ҝ2`�gb;�'��2� �����y���x
*�˔h�T�^`����XlxVHYEB     400     1c0.o�Pp�=z�%^VS�h�?E�g�%o�dI^Tv��E�$���zZ<�1N�����/�f,����K�f�6���w�'�pG�|۳�&o�t?���@�4�U�̒�2?e���.���>^b�F��ʢz+��SO7����Y>P),�Ì&�]VEx��f��d������٩Z a7 �x_Q�w��Ap/X!J���v$�\v����L�4�3Zl�l���!��|��{s����sOt��\a� �N��-�T�K���,?�����٧'�mC?��r}�=:1������K�}1�z���z�%]WgR�w�[ș�y�)t�.�&�!��0ؖ���h���h0���I�x�L>��v w.����)������PY6Dˁ(3N�2B53���pR���k��������,z<)t�x�e8��s����3{�w�*��JNc�XlxVHYEB     400     140����F;�YC��u��':X	*Ş����h���͎F���e��|�����o��@�U��?�?�RF�"��>P���<��S�����"z�s$6���0�1T�E�S����/ӊ�l^�T����k��?���;	�5Ýתc�0f�V��%�6\�o�'��n�_�ʰ)�ϻ��iY�������{�xV�l�J��JdE*������ﷀz���Mҭ!��P�
��C��=5����uBP-)����,h_����!:r���A�f�M�"��	��|�0���;+nI��O��ҥYgz�75��Ő�};.XlxVHYEB     400     120QTn�,����B7`�/�Y$�,0�0֞7gO+�s7��!�\������ݭ���<^^]�n<pasl,��
�q�ZmU.��?8K#8A]�̖�&8u���ɛA��j�ו*��:Bh[��G��z=ku���_�x��&�򠛰�}���I�tmsDF*����Te�i��q��޴;���+��WDeY���}��%K��:+����T�*������瞗�����$�7 �ĉ�������)
�_�v}�w v
��������f�/�s��9�\MXlxVHYEB     400     190&wy�p#�!�9V�Y�����ԃpO����ؿ�#�K6����g�~�Zs�Yy�w���tt���Sf�9�3�U�\����P�W�4�+����O
ޘ2��.��6�`����K��6�ح��1(��y��om�\����r���dԦ�C9��7&Ή���i���9O�9��Z���}9yI�L��$���#����ͷ|��|1�M��S�y!׺���*^��z�C�R�*_q\),[tȋĠAh�H�:��k൯I˗<�t5�JǬ�޽sCK��u�R�|md��zg����w��E�w��;c/�>(N�hϲIxp���' �Rp'2|.�!�۸zX=���6t���v��ON �g�`��ak����X���B��:pGb�Y��
=`?hj_vBfXlxVHYEB     400     170f�GZ�^Ή^�=���W��:$6:庇^���)Tc[D>1��zy��?	]� �GF�S��\���8.���΀#�.�8M%;�I�Q��IH(:��]���a� =c��k7b�!��⌞�D���M�ʓ��fn�սe��ߕe'Z����K�oD�ڑ�x��q�������������(x�z��M��e�Bs=���+�lv��Į��:���m@��d�	��d�Y���ū��rKu�h<d�x�|����������>�i6]�a
��с�:��.&:�Ì��WyS�{cJ�ãM��P��H�tи��5׳��-S�Qm�IlX�kmM=��:'l MW�(�j��pX�	IƟ�VXlxVHYEB     145      a0ꀅ7���g2 ����1��H���i�*_AT*��ڝ<�����o��%��b-���̌�p�����NsfA�O������9x�z�\��
G��)�A��#��@yaT9bUM��D9��WOL���P�Az�tX���d���k���h�|�7~�<m�