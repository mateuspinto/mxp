`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45824)
`protect data_block
qER4ahL7aM708zyYmc5Pbr0gjN4e8YaXYZUDHYdlugEhyGvCB65iRlPQ8wDp+7duKMUzkYdQE0XW
LzW7R9to39kjmjivCETu4ffdY/OHb8DcUXNpsp1Au8HVPkj8FJSA22uospdkHkNpNx6nY0rnaDF9
N2S1VBcOvUOeeyDo6QX90OBzQpb0K9OMF6CnFqY9YIwtZhzz2aCMAh8x9XitlHGkRQyXCpbkKmnE
lhOENTB0pOR0qzOk58En5lq9ckdDEH3JfeiwofPGu/uVJvUIpuZc2Io35hrNFoi6QQmRx0SUyXw+
AVZGrQ2CH7h034r6Dq7UJ/vsEdOrreHCrFpnBM4oGMNzHnwFye6GrD/cQZETUdfec7X5A6bLFht4
zx9k2NhAYEiABNcFOLdSqnK5J/EInAwCalLwscl/Bh5M8iNiE/F1IhCOqGfe/+692zcoaB6ON5/z
WI0DbzCfD7mcOqVSe3gAyLTonqAzQ4N4YF2ttGmih5j/FNq0if7VLh8PZvPGblQzprZ5Lb9U3wwp
oAvNdCHr3AQnb7/wm4z30BY5NJviNO323cGW7sPkhX4JnfJiOIXJ3q2o76sAWxZ+3M7apdlpJznv
NN0EY5agWqjGTEqT0VSPkN5y3kBGWM3L+ihEPWRbnahjOld+b9wFfmmp2fC6fi1acU6NxXVEnf6s
1bVqv+VeWlJywE9KcoDkm6zrUo2pRL1HmfLnZ4DeNLtVmY5xW0FfUtpUztyhQG0QWJfx6jH9t2/n
Safsb0BbVV9CsOzFioBs3E03HZ3dLBJYhna7aq0HLrsJMYzRanJQ6QsMExFZEQjPG2Mrq1jDktBh
jH8m5h6RD1ue4WNi4wJvPiOzW3RGNQoMZKWWmlx6uT3o8oCerhI0JYLi+dhbjbKuj/3a2G5JpMRU
j+AO4edYyAHCOklG2FgOeaDREORXPl9gy6LB0YEbkHEe6d5Shdw1tEXf1W7vqZiHNOQSW6rZDvYw
ULqrMrWYh8NiI69MZVHeAjcxMKac+euEPJEvKMMKEIbICGlEIBnFwbMEloYDKKDTA7JM4YaOtJDc
Dlh6MgltnilUdwBTW5Aej/HbD2ZgdKV63qJzKBY+9J/fnEVrdPGy+0SU9Kpr0AJnbEgxOtkR1Pdv
sWypTQeXkJVQG7Y0c2kPLQ7sPfWxY1o5WHt8lO8ehy4Y5an4LhB7K3eY3M9vsnEALHbk0Pj9yfUY
5AIhf3QZllZdbFA22D/GLP8/pzzr0AkN6qlnAodN3u1Qz7BzUHNK3N4UN8ZesGM6tgUqyUFki/Ql
d3j+4OR5YWzUHjLYv0YBm/1QD8Pxexyd41e3E8YpxIZIdkw3ZqBl+vIMHkouUXHWqMU8yoXEQ9Gr
4tviEGcoOgmA74CTNgaKGNlr47MyhLpfhe9yzsCkOSTUUBpSnsx50ZCKKVtF7CWabXqfyal4s9UN
kszT2GXqIXDj3ZtfbHKDVfLY9Q0hUDsj9LbpqAvv5b2tn3Zao2FSXTtwEqAT+6i65QsLiiUfi3M2
TfZ6s7wj3WdlRmL40KLR2oaKvP8X37UeLaP+p07+3QciFDl6PvS1f+g1a1pK+hqrwDaF/HeZIkrM
b2+2B3lCiih59ou0iJZAQg1XmccR7hqqkSlq2Ch0gNVHfQ8WqWb0VKWTHkYrBjFEt5+UOwk7vwtr
wgb4z2xb8HwX8B6sS9Ju17FMFYb4BwpFMYgBdodKl1QZ4ATWNrvytZ89+QfKzpD9d2HoyAPbRWni
IVkh36WIFEEcS+UuR2I/cctLTzmXZbT0Sv8p+wQqghWkJGs7G+OfZCxVElvP0r8FUezf+b3hhFlh
14Bb0uW2ZEf36qgVFf3x4lhwmTL+4k+PhdjIgJgpNMmE2xEcYi5X/SdoIJHaHUUZyVqlvbHfLp0Q
QShv4r0bG9a0mMxIwFT/IFbF8NYdwd44Q7dNzWmT+szzB3dR3iP0Ezpo438z63hbNMYdshjzykwP
OUsCyFTg36ypFJLx033c3NWoDitniVHElBy/5PeyLFuYmJSmG15wXZy+R2Iu3c0opTccyguR9NZP
iLOXKyI7dHXemcGDZjo501FYgPYJnzRz/V52X2vUCKQIH7fLqZavTcbVEW6/akYWThJow+k+cGQO
g6wF/qDsPppQ8mnYOFt6THI2prX9LPenBlmu7Zzi3jJUDRt9xI2AbBD8hv9wzlHd6LLsbvsO7FXv
HDKwdQ4wPIuXX6Mcn7EB2tjcI5+T7sRheZWajqxsJDHhZ7GQ5h5RSLY//ZzwZwszCPF8ZX3sE+z6
p24CuHLC2hzVRn9Z6KurrkC7QER07t+vNcLT6kesyAOOlUkgmOGGj3I/rCIZzu+MH4GYG4p4juUH
K7XDyzLVx6WSpbMsUTi506TqOa9YH+4BI8oE2NU7yJL7Fd8RWW2Yhc4J/7Xjdlj9ZzOxiPGfQ5LP
Cr7npEmIdfaVD8Qlkr5TIiSigWXSk1W6r7DqRBDKCNmgkty7PjxVsIHqwkDnz5CJDoOrvJTFh1He
IIEMJWHIwsOgSI0jhvWKptdb66ot9x8W3DnFquKQgkqBeaX6OQslDdFpOEInqbwfnkSQ3kqHSPyX
sOIe7QqU9QDnFvvhhL3Z+/CjDVk95bSm4dUEWSgSeVhXR35/gzDJpTD9WDtjho7A5my/UhXw3OmS
el8AWOBui5Z0wSUlQdqWpn6yC04R2afVssNF96uNKoPe3MjcaJgwU6Szrmt0g4tLv3WBjolc19UD
VRkteEdtKRRm7t8vYrIKO0XNv0xfrHX7Rq5Rq7fY63kwVvOgo0aKW7iUBFT6B3HeN1BdMhtXDuVp
yhEfBekxww4XoPM7JMyHSk5yu+WTV65hka0MGEFM4bAzLLxOk28oq0a1Y6QFjz5QMU2HM5dijrBZ
hcGTZv8TdkCT3Jenp7/bH91NsAVywbw3jPUnHQvdxFuWtrE9K/ONfyem06qqZBTI7Y9isOZkwAc/
bDi7gEb7A5Sg9at5v7F+Ar664QEBcFJFy1+cz32To1XkZZ7O0PaSSmUns+6RhE/IOIvAanDR9PuU
WMPZFc6fxzbkDa/WNvZuhCnQfoeMEFV+81jTzr4krESHPhtNMGeOF1/QoiJ8tpVPY4WiPIoRGRyX
5KHk+FOXGrmiXsJtCyS4UNDtHrNM9ArVL60F+tR/gyfzjxQq+XEYJ3/gf+KGQ81FgDI2fy9JRjkJ
Yw5egnlhbHNdmI8p18NmSeXts0wAk80rw8ajCdre7T/iqe7+JBfBOpRW2V7f/YTpOlGslMXJUsi5
5WX9i0HJ4dIiUURzK1hyRPsk+fZ63TQ/sHzuPOZ+3E/RRqO6h5Scz9pTE8kfdn/oMS1h7tJ7GKyd
XYKc8IjtWJC7dkOWaIzzvRVLJOVxFlk1ZLSD9m4647PBw5gzWF2MldMfWv89I1ghBESi99ViQ3FN
/ojpkk/tzdgWwE2QbN+LMO3d7gi9XW1fZw0l5VU3ADDOe2hG+4Tpk09ygWzJ5mEWF0w+5RQTXYtl
L2Blpp4QYMx05d1M8IeAk2P16GJXw0pVp0X8BrormAumEDKePRKHUrppDomexTyDAxEWGdMJBn4T
4TDx/Bu2y5Sx+GSKpCV8EqbUPyvBlgdFOPaCVh1pyBfwA6Q/b9+RTvjcS3M5itIsvc4efWDwFQYn
B1wSmX+kBxCa6sd9FaM1ShvG+yHcZqtzAzTu/SuwL6lBjKKpITs1aam5BANDSVPHGzxkJmof5jjq
d5taqloQUDUjTVf8NO3hkXTDPhFslKmtAzTW9B6mzSsi8VCz94LAZeweYZOVl2XKU9QnLRDSINve
OZGBPq8Ya2xCLvqD7bE71dzRbAjZlHx+xiPcBrJcetVmSrB/s8iFX74g9w1YxDLX01IlaQkA29BI
noxf3jkCYIolggOimDAVPFKa7vBRlqybAMGCKSN2XqfE5zf0jQrkbKHUQLDhFSQMfQ9oD3QvVyYs
ZpD7NHGx+AC9lZq6vKYentYi6jmzFbVDkbw60o3qi3xsZd7R2f0zF/JrYW1APb6YJAC131F83760
aKOlijaXV2YR/CqqvsX0Efc1TzM4eDuefiYaHSYmykdfftwEABndfuJrACsmZW6Ak54Do6ilhe8G
34icrV4k26kVkgf/nwkZxg/l3+5RGT2WMjOj2YBc0JpFFh5HhXt+ulQQpvfFn3+pGALDMVAbERmU
QcH25TKsTLHAwFrPr3qS2fouQ3U3TOW1gkwFEw96vDD5KjNz3XfLcvVDHRACZDw029YPDnl2xstS
943JUQJrsv9Mrgh+7D/9mMUsk6cPNPt2zNC1hT1WDn1JSaVQObvEpWp3PC/Z0X5KfG5gESr1lWV1
FWdkvv5o63iuZca0Ln5XcMqRZD9My1/4kJNt3hxpg3CdGOxXgJ6OZL8rDFenlPnZmVESFZGWBUc5
py+AXmppvSHSbhBIaZ1PReNtAFLYQRNGZ3E9d+aXMpPeE87iebujA7Hbi6xg3i5rLI2Kpwb2557I
BPFvH8qZ9d01N0ROJY8riPV5a1B0ftV+L+EKvzUiydlxq5+J+w0zSsdZ+7HnbdUQnOhMJ5QTU5EP
ses08muPXpgfv1b47A0C5JXdt6J5JPizQoMDAGwrWR34VnQGzRVDSnlCzhFYqakKgwDsR4/DEYj6
BLVmrykBIUdIvDjkhSlAmhcN2/N1AUvz5JM3CIbFGL5cJjAUJ6Xsi3ZGXx+AxkljdtbV+1HFBxHj
5LN/YWdUMBA/CLK9Nhr3TtRnHGQbesLKiFdzNAlcA4QIguGSTPT+DNAKRIv63Gm02XIMtS97GUWb
uMbkTfQNaH3NXifsHukU5y0DXONB5DFDA2J+fwj0GBXanZ46+FX7ywTP1iaJaIWigGDDYxzG2CQi
S5TNDmygmDBD/9XWAEnL9lTAD27e4xdg3GgpgTuIct8KwNq+ScyMp+sk1RSqYyPtjnCkqWPpL4ge
lpmhQ1GE5GUnxewzjH3nWgsOmR4NGjwywM47bMos/jYB0ejyrRbNycutyPQ45aTdk7GkI1ekBCUg
cxi9MIZjhelIh9H0/UqyFx2FH6oDN1USw2Sag2CMUUqW2uuQwODej3gVoHYQSU+wB//rDeC2J0eM
kjK3sEq4T4Hj/bLEiylZ5pp1pPKHIEsGD+XV2wG8r4Q8bF9HxPTB+rRLd19gecRRPNWKKJcIbusB
hXsDTXYYvN5eY6luOR/X69vmVD4rAE38x5LgJijHdQBCK6kRz/X9mrkk6t/aoHe3ZCdY6xg9BNKD
YxkKQI+aBh/7LTTOk/s/QeIVKN6fF1s3d3xqddEF2ziFG4Y3oWEf5wACyb2BSwZHp9go8ZwQrqDH
wCV7T3D6/2jt9RklM2yOmcndJPwaBPrLD96Mdw6vmlW9UJkg/AERC3VgY7k6JnfCR/c32DvDXa1e
DT6JGRn8v3O28zIrPlQB5wsErK9EUKpSYfQ2tw4+h/ONqHOADcc3bpCR1LO4kyXOl7VDoR7oMoDU
y5ReR6BDTgxLjimFDRhpOJYlPqeqykexNeXTjvS6h501PtXpwD13G97Rp3/vAYvjAt89tKTJTe+i
ZjE5iu0oOD0goiVcKOU0KS+gvVbTAdE8G8xFFYBKsR0ZAVzLKbBqoCqbwtZF9SBwm80hUxyhhcKx
loOEvNckVNjyFR84eejEtLmImlTcLOumPkhZTSnVa6R3kWJgvsfXn0inU/uxg0FZIIfxmNY67yRj
GJRvnd9DntkGYCygs+SrqD/riNiL/qDxcBZbm+fL+HxtYZr1uKb1texl4uin5WPpJ1u9WSE7bZL/
k7aLS7aP3OH82N40gLWcnfDBhTe5LdSYbiGNVZjMZIJH0kcGZ7YFryxCLEZFllUr0g+rmpl95jZR
ssLyZjzpNCkJUbTybZOV3VQJI8DaVn0kD1nlg/X1IbmJVz1EWcrDCio77/zweORB3G1vIJaRRlda
dXqPW05JPGEQXsFp0siA1SaLXSnoyNnkFAFkqYkKv9YzvvVrWcnQQXCprduFSaZwQm7X8W2o7jus
Obf4G0XzU8pk4oVTs6hTSyP8EoIeJpR7D5ElrmkZAoCxUraQrFoR+VMcxkibRivTxxBg3Bm1htXF
Q5fHcjJyvTOMYZfyRrGo0UCUSkNEfVIb36w4ixAV6Go+G5Eux+BRohfHQiBGCFMc06eTHzmiNFVC
qbaj0RWFg8fvsIKL+9qSmtDCM98io1hHMASFzqRiZg3WIykgNhCAvuUWSTr9BgneBJkZy3Ea7R++
Zj8OT0E4amnDNmPjwUXt8eC6A11On37wHb41itcZiPSsw9dVbiyRGESCZUNINuzVEw8VBqL4QsBW
zul9oAT7JRkupiOoEZXm3H/JS8VNc2V0oahxuGUl18uvVZcOE4dIk2jhuF3gTaDERFcFgNcoswCK
ZbfOzD4IB07/lmdnGBiijD9ON5unnExJ6x9+PfRQTntiZtDa3I91vyex7IBEkPDpLbawLYVdDq2d
R5ICI8TajvDOEe2dX9mUjv58TCJhLgcLNDCxI/JSNrVTz9e8n2eHtNkh0Dfbyj6cwCDytpjnkqdf
vfVeUqpLo7GgDKZkdEBkqEshUEfq9iCGvrvirmt1ADo+ZklQrlD5RZKwi0oPO7OFNenQk0jIqlpr
OxbTfwUBUvcZvn3r+esGSuOHSEgVp0nbqb3hX95Psz/PabLO1s7700quWCshxtJQiSy4qyCbISzM
rLpTLCckCznIP3MoitJvYBkJUeXstylNr0v6EXhyoQ16VWlQE3OTwMYunXJZ3ShUxWlA0WDpM6g6
UouT52sY+aJOvZ+j3i8dmO5X/vgukNJXDapzSadqVExrhCh2kzjZsERcTKaWm8JDu2Dyf6h89D/H
Wp6KgVdUgLc/9v5awKlDe2yq97Cv3cpD4Ch3DolzIgIghczGutnY8N97FIrNW9hHajV9P/PNhGaO
9Y6/z1it7oGI0xwIsBWZ5NrPwbfrLXY6B2HoxIo8hnvk55ppJPRj7XSFEJE9gDfllr/Vk7QeQ/5T
7G99yO/4LtVN/d8yUotiz+ZoYPVF6NKP1xyTGlOHFbAVcquL7u1AhH89q/DNp8h6Wy5N8oTsdBaf
5MECPkgMcW3vy4dvWnk3OcMZvP6kxSK88hc2E9Tsr7qApfwGSFiB6YKuehOcvSD05y8Vy9mjtPjp
w59/zjM4zw4IVpS1Rz/rJ6wc0D55Doby/+P1608zS5O0Z2gde1kfxKRZBsL/bs6dZEpwEhsdU22+
PHJHV1an7ZhR96HxJe9lSq7L8c/l8M7oDzXU5AQOlk8u46UOzVPQ8i25jJ3c3KDMUswyaEZYp5Qj
yAvRs8WXem+hL50COmGnIBm04mjC+2PGOnUaiecdcmjp6vce/jWCaTEfI/z0BcSDVCMtEO//U6JG
jnbZsFsTzigXXcuwPMUNdkQ6fFkgax+TbKG8BFaV1Ec/bgGuYQcjT9J4JKQDsL+h1jWkLiBdBJbk
giutJuk5ANEZRN+1R/3mrHrrtmqkpEms1If+ai5PKzaoDinDyZqmNRBnQ+kWLHa9/bvlEV1x+e4u
M7ibz3e3SoVEyaCUNiyBYzQj1kdJ03hyj4hDcq7b4aemF5gjrCikIjcbDjTvAVkK+LIw4TiQxhCq
LKcZbRLVj5RHZRWU0wfPmeo9KNtjKLU5jBDaNRX05TLQPcXptEvWD454gwrLcgJUqeY8sb1onW+f
wLkIrpTmHvvABFLecMIpQmD7uQn+ahbN8L27t9Ju9lve4BHm9VSkOdxspVhEv39aKh3/W3MCxgXx
czjGEDtIY07bGAc7cek4BJAoSHto3iWTfxAtALYqt8OKV+kfaqL8fREDY2fu0lMA7pNBQBpbwfUj
DH1MAdz73DEJIywQbGjVpN+klxAnTQRvUmcbN0oIUKeBdtT4PLGmwBQBfeeYe2qLs3fkTe/mQwTd
IzgJVLMI6K2Y74uGzA2o5gHXwWubAC5zc1TiLQf4GEjDu90pNO7Xqy/YhGx4sse9ddISt3WLLuxr
dY136jFRIoAJy6xcH26nKv5pYP2ZqVZobhCboUUgpYe02gUSqa26PHQKeVVrA74R/IaWVn4cU0mf
N2nZa2iTOoNCMQIruOeQ5GoKJyxs/E3uQbL+38FaYOehbJfqTgO2KncSP2LEJ8IvsY+OtiKD7Ncn
//P2xwU8Y4M5MFjtcXGEZlDusXE8WcqAw6tmwIBg2ZCRQMT4aCotwRgiekUB6iMEQQhnsFLmodIp
I+Wk+ecK2ePQ4NE7mc1ZgnfAcvkJlLwwa9+up6MTC0+LAwew4xc8Lu5ifjDPaJAkYythVI/sMAIl
h3TThZ+9bcEuy1GiDo5o1dvd+3tAbY3qOR7XKtCWefzQHym873Ha9nwFFYCMXNqmWIbNOOUzkMq8
EGQxPjBOD7Mdf6jR4YuM7sWpJZ++Gh8ht7SWsr0bp8qqHjY1v2LjDO84WutklhFsoMb5z5sVH1GI
/ae0MFp9aV1zFjSuYy7QtUoqLn9Ot4GW/O3RRWzRaDPZ+gJFMSSE4d893ojy7VPVVOkiS7K7Ftn3
J0pfg4xbvBA4k/HJYS6bJ4CU+AkYZaagtrLZTTF5iho4BTpYexvI7NeoQ3TgYAsGrnYXLAHvPPtV
9fxoUGtXbV16ejeaD7AKEAAFGJNzotz+hWsqWS4RbyIjIbt6ynBHm736vdwnrleleF4gNa0FfLsH
uBHoAOppm7xw2WV4XBU7VyEXMWocIqHjUGukbE6qGAMCNes8bGRfE23sPD41Cyr0xj9yuRHc/Pzg
GywynlBeqTaEGHw+Un5br2ulWpuyBqf7eiCCnLdKd8LXZ70d2fPJh8as1dKHdbNuMnPFi2rXkQYD
ugE4+EpKZPALtQe3TFXnJId9Ky4yzxZpW33g3hPhjlJDGDIrCLHoxmgGH6myxIPfJOs5+ZeYugwS
3avLbRaA8J7c8pOdVATjr9ap0J7ZqWY+NJ9vvsVXmg8HXviX/JvFtALuyzx0MxIIaacngW7a84m7
pSUtpdnt0lwLpGgpKMdMpQC3s5F2iZIvgE+OHu6V/hZVQEl1ICLFYry187OvL6kGDmeYv+pGRYRW
k2Dk0jcwtUhcuPDxjv6VcAMVwZQTvvDE36VEntRpa+QiplcDQVe/GdQjr4At4DUneJfeUA5f7qHr
wqzazxYfyUAltDIICoPEQvpJRDSSxsWQHcG5Z1N4Ym+bcFGqy7OgYqvHC3Dpy80T7fRvTEUOEDRM
GMbnSx6XWxs2KjMqACYDcHWjymS1yYxAGdQcokXqtsxyhEsluitQk2ELE125pM0a4oR9Mna6utvD
LWyfAaFfV7b+EhWpXnU5zCDRrcEJ6hNF6NHGFd8izktvcC4zOE4Tc4I1lo+ewZR1JCE+CGlRLojV
cOQ6teRhVt8L854azrc3B241cKmi6uodNtAnf3zz+xFKBvwb5+iOfciz9F+iDq00LgKecU4IrZPT
MeD314fcNTOvBOCVUqsMD5MKO5GQsyG5+acOvoeVqHZVFbOmXBzArS69nLJmmYq8jxQqzMSrapMK
P0nxJFHBeobe3kdf3nCvN45WQ1YFEt8+7ATjG9LegHZseCVTAYKR/21ji++WAGisGjWkO1z80HFo
cCLpdh4VJYmxJf7g9SMWM10CO8hL9vcguJ+1xrncOEVFkpoGlcFgX31Qku/j3qxIYPc4HCn4ADqI
nEy2ht8mprPh+jb29fk0pdh3d0Ggub1z+8K2r95WCBOt7JytUOsArEYlD0mLQwFJcRrJ+xnWtOFz
03mfIQihtiSqEvKUD0M996utnkOuHAyMgzHYPn/AWS1FcCeMUoe7WCB6USu/L6HyrR1VXwhmGnIY
z2Mq0RlgGyaqZRTSyxwnXRYHUj899M9PopVw/hWF4UdFPMPMsLhYSdnSRf0OynBzswPa7ggoE7Mx
q+VH9jZfRPT0hmTft3MaF9BNS4XFKn9m6XEjXBjaWigoNCml3YUbmD9aVkHHt9N0cibenVSHjNSl
oRpx2dXllzZTb3JaDrf8c9sTXecT/Ssz12cVqKl7gc+9IC7MbLI1OxsIp/WbR7PV3z/cI2IDRiza
krSEc19au2YIbzUTx3So1aeHiC9OPFki7oNPm5+tap/1gUjxRpeMZ6Zi2AapMDkKiBEQbmZAIMZW
ifchdvtOLKcqUoeUnagjrUFii0TXIDh+r9P9xT/KIGDGFUxJ/CzwwfE7SUdRcMoBoQ3FduM2YG7S
ciJfGrSGlHfy4KaXWMvEHXRgigaQvoQb7DAZ1qO85cpjeVBBkuBfnRkr7dRoWkypH42IalrKqDnl
C/hKlm9pDbV3B7Ybn45O7CPMY0TyVCZ4+QM4lOpd+Y3X1OkQCbbVbxdg0xsR8J4ZzzISuxaYazOB
mYeCA/gcB/jML4PvMha9+8UcFmLc69O+PGzLBa+Mp55eYqWDX+TuSjG4S4Pleme3Wpyq2yG9uV6f
xRUV9DVDfUzyi7wK2X65K3KfqQ5tkL3LfYEOyc0f1IFJkZUG38+EtT1n3ngMe+DScbF1oZzsaLBI
wAUlHuKEixgcygfkF7PCAhyWT6VKddIA2Y+Sm/0FzmdN0Yl7gTd+qGzdxIicO7ndNQoKGvQhALIm
GWNXC+K9uIF8LXW3afaQYUtl8IZjB3B3gfczO97KDspkU28UTNQEOGw3FTcWEuE9H6cg3XtxTJX4
Erl6jk9UXSgTerxwB9j8IeZtFdcoxx33IV8/SvVxBXJ3Ze4v9z3uRf/tPzbBC7QYQ2njPmrS4V4K
uHfhmkUsVseR7OiP/bjSAQlp6Amkg/ycoM3s6+jW1FA9bMuyJ6gLSl1eX0petw63OhapiMK8UtmB
fmOq2BhkHybfw9zgLesPF/YMaKoDDXxj/AWXCRhmgqYkJ0WAK6RauekdKE23fPcL8eFfhAcD0da5
gna0una9g/xrnoFa7gqQ1b7b3wcUjBlmUpacferabKVwSw53rJYMOiu21JeBPtmfkO/Ul/OfjtOI
ouiUNu6mKCcrAP+qNKuX0cthwd+3eLR7ugI5FVmGBmMVJmjy1z7qAFntVyutmBaxZ8o/QKdlTlG5
OWC/XPZCTUfWm2z8wDg73CJz1YQ8m8aiKUy5pXkFDDmVjMLY73Pfp0eoJs6mvDbYGtkKPbPbs5kW
qDQb24Q2JekwNCZRK5Pz1MeLYpZtBkp+yX9ET0BW6PpsvXpsW5UYQpf5hEw+V1gwWRvUczUaRdke
x9clToaM4od93pZPzDQoFoiEdbo1iczMZrRj22tUPgezHVICaKymMSOZgDVLgBDSizFrO3o2sZcS
iyuUA6aOm0XlT7hQKukzUBq5ovuKFZG+N/FDcog4rLqJpROwU/ExB0aybTRbK86r2CCYevVo9b2f
MVyrdTG7tEDkyh+j70y1zw/TF5cZ9u17oIqsNdAh0eiCvm2JPAWtv7CtgbSZgCcQuC3ifXwep4Tb
fUo/TXPy4tNMMGc3n/mUUZJYKGSomR8qVe16WA7n5teRpsldSlsbPtKmwYhd6s6lRlFP5MJZ79X1
nMltMsW6vgTwNZfA1QQP/ve0AEP94KHDjSDB6V1qKnyPNG++PS0v/mA7L0/viRyZsTFt2VPHKSl0
GhTEnZw0c2QzoegUMl1izskruwaKptS/kg51mnbOYmX5ygelLKwzImLVXAhH3cL1P5v8f5vE2wLW
PFE/JDGxwvLUP7qQqr8OaGt71GYYrhUrdfZmlIZMutPYazb3VCZ/5B3BJ6CHlqzKOSwPE6BGlqKq
+0EvVuddHGDMYal6uo4NxjA5HMJ14ttTyC7d9mdt5iqP3nKmYvBiMQvvay3vGQ+q9xhEk7AmOC9N
k7Blh5wfvffr9c02EJswAoUPgWOZgdQ6SfFP6oDfgjjvivJqBTh/d4INFmhHcpVVpVCe7KBMl7ts
AL//K/7tzbB+N2/fAeR4DvdlLo6jWeiImicDYqqEDT/2IruNwxXqgis7VAK+1vpyxb3y0WrT7i2i
rjA0AoLHuypsVul2Vo2L6BkBJqmQ2DDpH1ke6J5fZRo8Gt04tJBo06RQGlt8VS/RtPCv7tHTYqUz
pbzMSpWSVPyNLs6mm5fcRN0MmnjrAKbnwhYs+IVGxLev6zrrMKYnVzGSvFOpCT4onwCUQ6UbG7iP
4ZpcDyEaKVlQ1vrIKgz9ziZ0sEvkZ6xBjCLbjlyyGZdqRrVD515toC8IVXavkAl4IgmNXhnzCSZo
bCoZCnXILDFKoZ7hscNa/AlajO4LjOCe/gOqCxuubxn3MRiaQKQ30DDQ0YBpbTegAfsa84RZJO2e
58OYcKgu43HDIA0glAByY/igzLCfFYsxrXhb5d++hpP7Em+ioiedVfe3nKyQRGSgteGm0Wecd4VL
bE9FFNgU/FTAxLm6t5LwCAlRZfbRzDl7Eqr5lTgWAvAF2nn4fzKnkr3rBalPvr/HG3ZVbbeVAGeH
73cwwaLhL5ptrpL+ALGzpPBTdbTRTjEwo1Y60fKaZn6SqYE+o4+7UbaZYMYwC7bBbg/qnZUh8RlU
lQhBqGL2eVKdb5/ql0dixrCbkVhn3fk+ZULsDbdefOkg3Yhya75crBt/Zy1Op9sxlKJ6FRR5kjyU
RjyeavNy7RyVMBlPP4Hu64mkLhFwv1thxtx3XGLkx9UbUu4PDFxu6CBzHcftwKDlcTBmuf9wkV+u
BCGzErG8oErM18VGsS9z+sc6vX/+YB0vV2m0PThxLFTdc3zb8s3gJa4Z8hTJ+UJ5hkzPpzXiJ3T+
3RJA3LVz/uYWi5Xah7yLLW8sqmgFJrE6tHDjJKS6lsxUgMSJF1Delm8MBvMq54Qlz7V+S+RZNjnp
JID5MSg3HuVevQmnPVQu7htvLmHpqv1P0tW8FvNy+SvueX9Fp7XEKIzy0hVfyOw/ixEFex5um65a
ar7hnu7lVYWXQOxt9WaejTCJOPWeIi8+gVqOnESrkcntjcUoOERqauADHn+klTJN9pqc4cXmq/3m
6Wfh+0Dw6epDw2BURzHv3g1UPFfPPeji/UooVcYhvvXlK+bLzzfu6u4bYY0HxaFwmfJNQJVHr48A
NuFnirRAjYaDvkkomXY5HwKq6sQsR3cy5b8Gh+SmPMzXimKRaG27wwc05W/suAtFf/60R3JtoaAJ
V3SJOmVh5OKhmw1PLGhc9z0AvD2BFX8jd4HLjJ3jBlbkvX3splwJMl3wwd06A57CQv2zqZBwN9Am
bxdSRZohl38GtqL8KiTA7xsLUJz4SrxITQYTNgej1lVohQ3yjMrgHVqBXFvDS0cucIk96WbkLvVp
lMUtel4A91dxAA8vekI8YN2JLtsp9RLAYqhHL3ML55wUUy8pS8Say/SNM05hVzbtxLoGAeNkkDYI
FnXpYC8nyUA86iogNkr4kxx4KDPnULGSLSlEzsnPSPViCPhIYlEzl/+rG7UKM0n4hWgzSAeMbKzx
/MPQDqba8WNTXwrirHdH7u2GipulfqkSw7vpLj1GXUNGtFFFAuyR2NOsbZwAxi/inUWrUEAlWzRB
Mm5hQpIHLnOlXzbDuFVRcQCGMjXC7T6uqf4KX/8G6aBhfRo7x0M1+79Fhb6cfaQU1Lj+NzhRva+E
FBP83YUFCR0fksNPX+eeDlf5gQNp5TqLIe8cB9F+gkf4MCmlNfk/N0e6StnF2VctMLVBtUKkoLjh
/awtcsIkIHFuiCzRsFagGulRzND4rcIJP5pBlP9qmPPIbsfBFfh0/g2QWCc4q5KKtzmpO7qpZeR3
E5QSoVq7XYUaI1Lz/ScK/PNxby97gE6sNyV4FU+q7QY4jzfTBKtfwQ+2EyKsuCCosJesxpqyrCul
8K2bihT/gqgwVpWLzSsteHEzBeV1bLcG0cVcIqeEVtCxKKgF3UHPQJqsN6Caa3HvMPMfIkuMTv55
kkeBC0h7/EXxWeIVcYPDdPeuxlDyquNDT5ErsniflBMQvvC3HrGUwp02fH5+MZqQmZcaLI1Umkq4
ozGkc0q0oHRzU/g1XHix+gD3gdoQ/vufsHRgIogd2vWrMijzLN+tYyV686VfEV5JNlCGfBUPFJuN
NnDfMfIm8cv+jFDFHeDAczKwzOHsDEagy4wCpSyRqjwV3bx42gWyPefgkPt03+s49LID3aF5iPe5
y5gtxOopqCptYcwm5w0c6OZLGFyRgGxetQ7xEASHPUnjxabvOj6396q9m15X9d2aaMh/Dyb4SVYC
kbW7QJuVWBkG6kwgDx70ejGDMb0rGv4At8hvvyDpghXvaxxXmrBVvZvysTrmpseNLlcDzJoC3PcL
ju7czhGOTV216VNJLjbJsk+YYSnn2a5yYS1ZFsx6jVvRM6RP9fe703J9Pa31BgDc1xdfJM+Mno+X
yOMi0kz/fbAxLhHFTc4whLHnLqHFUwNHucpcMolHoUD69TTmpBHTF3QMEh8xHXHfy9DnS96EPYGp
LbdXpAeHZWrKJSHzP8ZGD+GQ4ptmRUejoWrCLFnENG5o920rgPeyedGWWguWTub+zufh+ZOPufjo
LBTUuzA+Y4QMFuIGgX70YIybZJ/UZQW5IE4CI3TwB672bZDN4bKF5eBOryAw6gn+Y9V1Nk5Wvse0
brb6igOas5/Lm2pRZBPlI5cPquxb+AMd6GlDxlt1OoUtYpV9Vc+rPaAfEDcOD0vEssqqxdnuUPHA
HL+s1iwHb9fkbeNFnQ3EN5hd83t27KgHx1NhKPLJ7zDUiIw3AMtdFMwLX+wIUrq8QSSl829vo98a
pFEBT95yjZ1JAdbfAUIoTLTfgTSGkA44Re6Ov6Jx+ATnhI0VUIU+3gSDgOjZwT/k0/4v6x30aDsO
rlut05DUOlthj/vuX6noOBm7HAUihZmrZh+6jOhBABxTk/JfWxXrIIuQRuv0jU0bwroNvbwhF8Hm
dO4Hm9o4VcSMfAHtEK76XsDuFrExjaJmEeWPi6O3FRIP4Q2qHsd0WRwrueRBWYZGCyE6mmJpIU71
FZXKonHqC3qVxx23sj93vBJcEjPN3CydGqPmCZQALuAwqsoDqa2F/nF9yqZlPN14fQONPk2eXAfb
cRVhEDqbUFw/aebWYmq2gY37SJGWXe22obbOxZyIsI/K3eMO/F1vn2RDuuw8KgnaGACXhiZJaswa
x0aJPpH3hRBdNs+e27QOE2zBiMD/9zMY5iY3p8uM81caGzOruAfR7GW52e+6U0cbAjmMTke6Bva2
OWgwIrYkxAKKxPDzHbFhtE1CYQjoGaXewWID0P3XWcV7ZMM9gEf4bzVAL4Aftdsmu4c5PV6irqO5
1kTndqDY7s212RGtBc/3U4i+WhBzyztVr7XLz3xMRejHSbd9Bkb4ODLQfzcmqTyYs04BM3oGe1jF
VlKRXmvCLDM7NX/Zl7VxgRDoHg4wVPFXZ2j0DxKVXmisZfXvC9uTVuH7et6jOYg/aDIdS3UrFmLM
mDBQC9Cq1JK0FSenVrgYvAWbyE5MXxLVitYWToXlyfc9Ri6OzmKO0pDlYrdwzeaw65wtvXJdHTfl
9Wgpb6ZbsKH1SCxvjMK3UDuimLCDnWisDYABW83N4YlBRtYIPy1kIBakozpjL8b9maiTHaMZbuqp
FEmVGWq0lp1XnAA6dPDwt4FtYjM73gvcAW7f/n4iUJt7gNkjWSnDhdt+WPuap5UirKtUcoUbNIQh
4HtkgscBHsdhU0Xly9KtQRJC0zA4zYTUGzrfqUpWtt7PqHdckGmpodpYkKoezkmIrhjraRIigQNc
rHMFJvqKpfYG6G2Jo78DC6xMIZsBXjzzwAiCGb1cIT7cGsnhD+YUD0lBVwAqpdiVb7slNOYnETmH
tUW9o4ME+iMnpSq8qUbIlCtPRdlExJvY5CbJ3hjlHitMZMD3FxwyL5uQsNO6lA7uo2x4ytzLfs4z
sFgD8KOGH1CJ3itOjZuea/Od8xm2BQvrebOVFcTzUnTFAlLPgSgwP/6PwhZwKR2cKcyBOMfIQfCJ
OuhgZObgDACOSpZZ3aJsfenywOIWN25P/d6oRxC1u+To5voApHmAamxolcGW7aMeliwrZkvcWha9
gRPOrnXnDU/o7GX/ykgEtJE6t0LjsCOhqSnJKMErAKXzT1oS8JwyHCUuCxrsebiWzxwoMHJZJhcG
AKrmBzS6TF+qatH45xFlvTAO+q+oFHV3Rn+yUiP88udChk7b4DpPA3uZ9GKCgBjyPTE2ovMUn+ts
3wwp/IKO7S87zqEItGQmajXiG/tPXPYU93PoeYYMG08vOD834/417LczqvBaEfzbNpkJvawwQw6A
dn1KtkcoVqdrcV1A1PzP/wjQ4sxDWdIVqnv2yiuATFNH4N/+WvOgQXZrC2KuvMnOKl2e6a+IuM9Q
hLIVVSyFBWoqyfQCDdrZxkRSvLDoVIWuKv2iDquLuz4MO82o3PIRjmzDgjkKdmXklJ8xI+vJAILo
e9oudIHcuUbNvb8OAtcSzKOQ2YqBuHe2zTumUvk3PMPFUTslK4Th5P859RrPSN99vnytDPjNmZow
BXXmxX6a913wPprt9/f94OD+lTAfKOeOxaPXvePtEFk+h4haAVLzLZ4F2pH1SOjctpISNvob2QJb
wgGoEZUfgzvTSQLo8enem/7lR81X4mqbUmykGfkI0p23c+FAg4LzYRV1P1mgOiqt1HBiZ5RSrb88
peTtjpFUUblaslPMN0Cebn2iE5bs01x30BB3zuuoT7HomF6WbvA08gBvG064SVm3yau8Ax3s7Fnu
Wb/dHD//ALBhaosIXDF5KtgrITtQclxc+czJU6Dazc06jm+FuhXAkJk2+GVhnipEU2IrX8gVz6xv
iu2IVjk1i2w7WMwaa1W2FboFkho7POFYuZO5ic1bTw8XGW/ZpV6U1XTxcH7oGPF1lFTNCr99IWQN
lGMmqgc9OP3AS+sWqd6BYRH1l7TyhUZX56YsIHb8yqTs5WJ2ezvLYLMQfljDxLHclkgjvbtQxQZW
ns89Uy3JFJhH7iuVicRSgIfCDdchtzYzplRkskikeEWOLev9MCxtKH98Nw5gwKRdZ1A01+kB5VKu
/7fAxTvEGDlrXGou8cNtZtmF6803OCHAFYsVjX46IO/4ps7iAT7AmSy+85icckIRdy6pd9TTRojO
fE4xVaaZZNcLle5qIPF7F3r67FmbdZB2UsUFMwodhAg1f55LKktgDI2DeR4brz5MKkrh2lOdPAXX
FN2JWegFO02MqnoxPsFo2k1+PATUFLYkz/usgdm8dNjwWQIA9qJwsM690QkxuR/dKqrzUSkUn8tv
gJjdfvvqgIQcdlvK1XOHA56W/NSPnbnGtFp7hdZDFRTF7h8cc57H2CWYNUochVHwog/ndwQ1iqAc
RAjnhwwksi8GO3PvNFtbDL8ybZOMpV3sGxYAt8SdkIh/AC3QDPOxqqSAsWBvXK32lEwim9h2j0Vn
txOxMoTBgnoRLAmJjKoncuxtRNzzkJRJZXDE50w1ZX+rLJVKJbRx5+m2SAeWI/iOQxETwCyCzCAC
/SG65cQBnKxrj8XG7+atruiA8kP1RruAzL5jabqsuzq4hcJBoFzIm3Y1Er25XRTQNgANjiNktwUX
CTki4LimcrTFJAz3xlT6wSOslzRDg66e+SnhvRDG6Bk2EiPv5YRI8KlRlGtpzXMufQjlL6cYep7Z
k6OddfIhvBcbafqfs43WdIg2g5cjsLbszR1R2I9WNRRJ57WVLQUVDMwNSke8jnii3O5uK5pDbu8T
5wccWS2zslqJ9ZuHgLAX2CRLLvyZVomWsx8F3G4N+DV2hd9ccfcwEfzt/qVP18fgs9wAsxuA4q9J
ohnI/uQYygJmfM+qNKfIJyAg3IMXxpTcel/+1otMZhSzYp2Zvtj9iF9UQAmeBCZAP3ZexTwHnIkP
RdjUQZPSZjgLYFUuKktDqKRpkph+134GTfMeToQeRfBllaMJPbTrTZyq1rQ1YekPDnwcFZVqfKJn
1G+SlA92l/m0P3fQ0U8aDO66U1NFXlzszu+Vvm57njfblKItQNtQtO9zq8QvXSfGgWkTrRIAxvuC
M1CMSF2uZ0E8ym2Flr+1dX60VLJGE87i0VgbEE7HE9eZu9PH7pRJ2kmvm9HPX5yFTAUnBtm+J1Lb
uGVsV53WRqRUnIJIZPD4C7esYucLiL/QGNt4SdiXdObzL/DxEUi2hmx1KkM5ElvB2vzRFowv6MOK
+cWPlqKVv0HcXbx6pc0CunoQ1Ad4LpPX2+8L+qqnvrnxhmLc6ZIAxftMsFG/xx5eP2d2zXX6PlBm
FxZyqR3Y8KHZLaqphEgfkTbfZx8ykv0p2NJss4DIvVD/HRALE+vF2ypjH1q/7XPU3Y2mSQjQDiem
pc9U3JlnI8Y4QwgnKIom7B2R8b6WH4yIM1yXuqOhoMAkSRpdIAmKLXxackfdsqGSnSKX6ENLQXff
VhyI9ejuXTqHUNrxFa+fV2WMa+LtEXL51jwxSc2iVnl8ECEXt+5YfYmk+64FRCrEzFnXjZdtGlet
PtGOwczluOKewgHGvQnE29iOJpDqUC9+oGBuIDRpOqiYuGDd48GBlZ8xluhR4LN7i+UHy1dSkF3/
1e+p8kUyitAnGL4DRn/4kPyNBWWmWopTnApt2mle1q4+WnEv/9bhivkMOP5zmCuk8cMDQE8HHyu6
Za5fVsODi3+obkQYUCqzXZE9mu83lNr3gIwa7GfR4ck58Ldaw+9PoeKeUjeX3O+1CajGlfmbk9YZ
29BcbSVZVIQGHR427lgtEroSz+xaQoNAduV2exuMJaHnX2+80iWEtBS5eNnp3nWBTnF20Is9JtW2
ouWJINGGbSvH8zpNwcjOwR3GIXi5RFPJq97pi8gZZw4nhEQr83z4EvOP+Oi5ZETCIagCKiLt/3RF
P9DGFMDNPJhydh2OC9vI0cVQAK2TPDz3zWRDWdmbQPfI3msL+LsF5XWsogB4A+i1LYdO+m2qzGPM
8iI7gon1LD8URWxDaLXzVBp4tsyRaK57oQe/eQnQ+tD6ksNj20tF1+nWf7T9sCFuXDtYO6i5N3Iy
avhJM8b3xz+S9/cEY0+pQY1rPL4z3G1lbSIFi0oLwCKxkans3Skn9mtNIvczaOP0t09nV6RcU16D
GKA4lhF2YuexgdhXNH2Fzhvb/eJrc7lNwF97ct7P0Motgxc0NRK9hQBz0biaC0gjwNI7CAhmFMkw
coPlyKyV9FsJW2CFgFA8ssICc/LESMS/Nv8As2czdhywyUf/NCJDjwCH6hWsaDs/fwPo1WI1d3WJ
msi0bE3WYtBEICcoNzTe3gGFwsTGhr/zVgqqgwcdzvyTle1jFhCzN0PnQpbycxVTgfPDjtHgOWS8
EWzHuBZ+plrUIFHiRYnam0aqPuC3BvnQ5DYHCy6ATqMDe+s6kVrwPao1DFYxEp0Rqvy+DLUQrLe6
4qeY4INjd7Wq9K+WIbDgjGjSP3d1n2UcGy+ynzikdnNCEUqyjPeEJfRh6UXuy8g9+TLbtvx4kshM
UWzVw7FZsrvDAPlAT4pfKwoOMpn83IT3U0p35Ii674rAylH5suAhOdOV5Xe9AhhS56BnOACL4xms
XeWDdbB33TKjrmTaG+IN7JnmfdONPTiNrMPlv1E00l0fD0DiYDjapi0b5yeS0EtGtXriKbdaxGP5
fmet4mhQto9m9YSmEJDCcg6COoEoE67aM0Vn8EpEx084mzp5pbt310rcorrBQwVRMVCZM81fIz0l
6rue0CmdAdosunilY+gz/lFCg5Ecn6oMuf4w0H4NvdbLEZJ2vpoL8MSoZevTsji3nB7vUICfbty0
gCqkO/DXrH84d2RD48l/ruANUiSp5ihGfQw6iEwS9w8Jo0fHMr+NqC61SYI/k/CZ+yvGqiajVcBL
Od6Ej1tI6VSl32IutQJYbg70BkG5nsip7GEC5d05BLme3gcMJWFAM3Vq9MeJHCJW9B/m4GK6d92X
/TLpoqDNSy2VscWlpPtt5rLYWhn/pXbyBTLL06B7pmjBxbdwIDmBMUpUCQPtHqJdPUxWCyhWGQBZ
OklGkPKy2vl/vdRenMs8d4o+qx7Lc9rJC8tkFPECfsfrMQ8Ai4XBpSv+IcjXzUF+AuRA3H0P2vAa
4/s1e3Oo9WGnWlPr9/BgNEkU7oRhll3Lt14qY7ST9BMc+xVINVyWIci4smIzTawqmxEAscJbCQz3
c7WD2VQXqeRIU1oI58//X+9L2jku+0e/O+5VrPzfn9eOgoGY8Da6A1ptvr5sfy5VvTTeYyuoYzMi
XVOSQ7dGrhTJqufdXZH8Ek8jhhJn42fK//6KVzj6nQAxzh/NgeWoxnM3nTWx1yUgvpbq64OWWfas
1v9Hax5/MMfo/E6LuuKNyY03z6Uu9Wkv67cfB+7NdIVzf+XIcuVxzxMgy5rofGb9Al60GHp6BXcw
m5alGcnBZrbyoaszPl1D5I1Yz7XcBecv5NV6arGfncQpTb86IKaUxkBw+4m4ZtmGldSG9eErj68K
iz2BjpnW1R3Om4R33/m3RrQOQkVqiqoFR++PRt0sQFEYFO9ZW+vWAz/tSFpQOI7XSCBJmDc6J+nA
KGKOjbunU3t9cwpdKHJl4U1itw0lyHRlMPqTdiwVUS+BA3wXAaUH+R8N7NQPbuOGj7W5/LJAGRje
AFy1D/CGLiDWfwK+SbfaKD+m4zGj3VkKgkLbJOl8gO/FtuPTdhyv3HOBtFBF5rdcHOjoDAGglnwX
cqWgXF3THw/BrBeVo4JPgAYp9A+CJ4krBl1ZF9dQDmDDuLLw7CZkhDyuYNptpOY9zhjPUXR7xY5d
+4pcK31e4vIYlCLjo2/91uh/D2Ts4lHeGYPOrvaMepKwl0WdOt4fLBwMhm1/CidSIqSaEgp6eeY6
QaT9MnugH+XfwUrBY73vq8/sxpMDy+Rfis8sspgXLCNakKdmWssmSRmHsWPvMrf62U4COO4TWVpN
ifYlHWCs6PXOll1lxEXV2i1SF9G2okGJrtnahiKBphiSeLAFA7QXCmqs291oysGYEclUEMeVQJag
ux4guIY+SRpSo4UNVnpmyulMEX/isYtmIcqEgTee8OtSDCnz5cKVqEBNU0XOApOkBYWfCVignj4V
th4daotJk4btYY6Y/4uYQeOtr1nNVT9GQXNYcWpzgoIQqE39hgbMjwq6ewsFLuJrOhMc5N6yqWsP
HmMtb1Jv++mFuKhCTD94zDiqc93Yg/1J54c1ZsU6vLms6/qhbTOFrC1+dMSxLJLRnOjJAAQn765k
9K6veNqwv0HC/GtWcLBl/dR91Ta1eTNcID6W7/h5Q6oTWv3KF4h6MH9x1GHPnHyQa3OhfRuPwsE8
3dyFQ3qKix88t6RGwbRkyuNS4Dk1IVzNQ9gMeELyAKL8ppv+0tMl/GzNpAcd9V+it4v+ngdmlOVN
P82NB3WDTPvKt5a6iExMDrzuu6Ndeocg7+8+eiNv3r+QxIkZ6++9olfCkUYRruQMTBHmNDQjlP6G
QFC6eHiVZ2B1e1ehtqkES2Wohxrogl5r+06vr3yvBHAAKk1ukHf6QQsE9LT05xLi5p2FBvT54Kdk
lcUSKckwdlOR2uK2Y1ErWGhUQstYoGyK4L+9ctCb1NCaCJtIkplF/gW2GudNKk2sBGiRBLF4wdTK
aI/IpVrl6C1x9DLLkmMZZp7pjRTqPq2Kr4D28c2OcoLQy8IRildLqRbqfLuueCce6zmAXf0Lb4VR
h04lVntPfXHQXmeB1lFHP32xgTWzSntp3ZjaVoZcwvYVjz7T0zBFnqS+njuzIvxS7tUn+NvTEXIP
1CZ0JbzWuwyeXZ6mXd+RCmyz1k31eUBUX8WoemOU522F4uhih7IUgHPD7SuujS68dQlTDfolj9AK
dcMsYmvcwTn6fo+e+fBMt04wwD1XKbNlkkSnmyKfvb/xnptViewlX+fAy2lijv+mvXuqqpkGRO5H
BP6r5Zs5n7yVGwfxGHpkzP0woT382VQ0qE0UjvQdUY6zEa8oKXBrIlUm+iXViMhxZ+fDR8xcpd8Z
jqFNdY+hAU3B0TguM4UKNKBXmY/AuRU3Pdc3JgyVjDmZeN2CykJ2wS+m/CApA+h5ybhDgavbpUHG
mpzbONW3IEFrErcKE8686oSb+u2f9CO9D9Z1adbv/BAtcd9NBUJzceylYJGBqNm9pAZTVmUULlZg
l85F8NYsdP1BddEeMcwxt8g7DM+O8x9LsiSSrTt/+m9TgWz1O9JsmYY4a/8bfAH85rLRyFd1KFac
8cpH5XRuPE970zIr5/ehA2ZMWMeZYmkQi3OHHdj4DyND3m2pM07sJWQLRK+40iTWTsukHD9mnekX
Su5Vi6MTOTuaotdO1/n2f/XOjBMBsoEfTva+PXsv5aT7Dkr7BacPLPvXKK895hwjaEtAUF/KEGlJ
NKFnu2J6c/E6j01kDeLNb6UhDoZLFSpr2WAvIhiZ+FXKARM/lhlJYCHZZO7kk4RzCsyZTwfXrwOn
p7tDwxuJ4SaODvrcl3CiMK4h1YnnVXg4js7Qak0V6xOHofidgWM2G+n5UlgpQxl9g8vqMH01fDVO
zda+LWukEMiGIgrLttP5srY33xDAg2UB7I3JwtB7LK32jS1xd6n3dzXDENsBUxe7qI8rorytfeOX
QKpt7usNIlDqhi4qDeEMArF48et19yWXfR1qUjru0TfE18h7s4sORXkeLiaNf5oAmzrFLlONWetI
y7BFmPWvQgJw66189GKzwtqn4m24g5By6VMlygUsLvQqwBecpMpE4QzfgeVDr9T8PJRZovmTL1KC
Y3R23yiZFJyJaDVzvtOoOiQFYX+OHXU8ekEnH07GMV/AjXxeAMPPObg+pRDP7JiOULZaAVr8vD0t
guxNpBUusILuaEzjKxk04jQw2fuhO1cmK+twJDkgCvwMz8nxuFCV/Kr6dJh3MLGYaTe1nlk+3scz
LxwwhOXLNGxUEwT9RSA8DHHXtgOAU1x2U1dfeooJVoQiPSmP1UyEmuRKD3bGsQktegIWLzMrkAJO
IHcQAz1b+yGgSP7sDXvphPcrIVCicegLEFcMkC4QAuEDphnNGVokUCBVEx6uSBBEhXT+rL34/8Sz
t9B2N30tzIQ086/ysgoKikgnyNwhz1afWlnPmbCeWyOK01L5xQKDKEQA8d1XsB4zLyPvx5nH0oc/
Xbo2Q/szN8zIIpXMFs1ztmPKoggaFBrGhyn8eEPQPTX7du3Vljx5kUeObYrkh9wWkIeZOHEE11b5
SDs4ryRKKDsK04E5y9CkYzKZfdOOqwIoipyv6ofS+ADvOHImMII8N273o8jV1VrS8dlj437sHJFI
6vdfWDgOGhMZyojiZEZsrnlzxt56y9oLFE3oxaJdutxEZZz+tbI4ZBw+P1LNWozCobVCXLjI+VFF
jZnMDxcSFvqPsI0BsMomgxfB6vpKsKvTjtNsqOwQb6iOwexIoIvQnr3Pv78gdB8phKLwxH/PX+9s
PFGwbP/NXvUHCoF8jC3pWxonArC7XEcNtm3m+9myoZhkrivWs7FhN+tnUPlq4MQvMUdXwUGrvdhk
eQbsD38WABDwzbEAGy/jZBYGKY6t3y1lAdkFhEBxV4SS+y7FwfE/1eKpVJYKyxDhLfT5eOYrVu5r
eyCPn2jTXB4vMoZp2gTdEGwOXyAvpcnYtmFZN6NtAHrldAVpkVF32XvOZMv4iInk4Pb+RtdBfB9R
bVYbLiw21lzf5Kut/o/GVEL1XqNH6RWDSPGE0myPrB1yz3ITx865+othW9cMxWEJga38QE3LFgZ+
kQEaj5alV8RkzuSQqe6rEoSxe1++ZGLmCj0G3/IbzIRe3f5BRKItqxvJbja7qeYljEIWivUMQG8O
9FoWg6Qqq0F+USqrzgRp8Z5CzJd5b9Ot1iFX8dzxk89OpcyoHmfo5IOD6FeynX89WC7hFSn8WJW7
9EQKzYGJyFEUCnlDPBb0iW9N2tRo5wFXUQ6rhtjuw4SXnseq92crP6uNk14vgRQax3+9BytiTmk1
xZ707zZ7Kz7s+mDA5V16gtl/Qlq/6gY5AvJPuYv/l5d5EowcXvFtfDIcAbNdFO/brtYSk+6VqwMa
POj0I/WzN5p1/ParXdkV4uCxlvmyWG7WaVs3C3SjC/a+Sb3o0XKvMhCMuTB/CguRIDoi0CLKf85p
s0aGia1eoR5XmrTxk8ryHHZkjEZObWCVQKOnTRaGZ+OuuswHLtUKwJSRwQwDbc/M+cENPjymdFc3
lBpGfxpS7yk6f3LthZLOFRG+ziq0R/tCn+tCCODskglj7gj3WrOHXe8bOy/boA92pbpVcxK0Bmdo
jvEzci7wHypyiz5QX1ld9KXuzKXo7VJTdgiSEHVOAcVcitHuP7Dxut8cEi1q51yEmWfNVJErCTQa
d5Gugby4X0PfQjgq5f7SnGraPcZzxGNnFBFMj47oQ5LslBxUOosko0PJWn9+gmJBFfh9qQGqIw2U
q+Krsy+OaIDP5WnbR6CozrZaSMa8ZewZKt6rszabejYvo6kfidMqMGmPi82++LzGEzwAPbh3EsWW
91QpTIsivNwR3gr5WFA5fwqEMWYgAbaZl34E1wRC4kknnqPppiQLBPONaNfcN/G3o57ELGYM7Sz7
CR74pl0dzqZpb6rzI2uWgB0RIw06J47/Ci6N919Ou8Mezdq9x+z5bpmi8uw0y6zS/FBRT6CI6mXR
xN4tv/bR8334w+ikEPrpbmGA3EXdU/F4qQm0FN8tx1RUUoGXgMSo7emqj5Dnjt0cJz1HjzQRR7bU
7IMGwxumyl4znnp9VjS1RbTEtNbdxusAXqquOxDOPSnGeyp/M+RfXHN8vJmA7L7a1RRtZ5WTWLDe
vX5yZtyqehbftQpZYcRnX9tdeufs7I0MEg/rGDEvwhIGiOIeoM75xhQri7wnismKGJDPMMY0CaNT
rys0GnzPuJufou1bqoJ0Eab7iHL+kgGPJhallercX2qEyR6AbU/ly/oaacRT64GPdJfWd50Ivfyo
9fJnUy6abv5TnuWtwknZfNoPY5ycsHDbw+fdpZ/MoipLg1gZpmLhPWyea/141u0/AmbtBMluOrHM
iy/nvkLekwXxjDOw9ex9yW7SG31ia6FtoItbM7dQqUm8j3OA7oXTlKAKHF6KZsvsYhMVaaPzxx4t
OUL6LFXW3HZHYKh9ECGl+pEl7LmKAlFJhQlwtqiKB5gthaZutePq1//ByULxNscul/Q81cDEYeJt
j73kxcWJL2MVQFwV1TMunweGBNPGDbI/IL/uCbPJqZJ2b16ASUwrVhc6wCeL18kaQJGLEhfvkRb3
vmJJ7hYQGNq5GcCb8+22vRtLThrtVuOVOmNBHsbLQoOzQlb3k9yGCPStJIxuSN/t9BKBIc3IJNXT
ogS1ypsHKZc52GQCCw6aMwwGNIERwuuCqJxeas9MhGz8/0eUuYV98Ybs5CvGjlmJv3JYJxhbSOna
oL0JDrYZgUpW72JH1w/m4ZEc3xDqm65nx7uPkijt+H/PMI0DuoZv3WzrGomLRo+YiCWUXpkIuevr
J6tdZvZZmnnqdg83f6i3bNAiet4GfND1aYDWEjzFaeQdUMQFc8Y4U6u3eqLoyLYUuDgnczErCu/7
kDGqwt4Pjpj20aCEGnlpu3++hPMAvBAwqxw/NwnyreZWPrsYwR+q2DR25EenbK8Og2ydBeqJhv7R
z9avDWFRC1BaPHThXyFzqXTEaF4fuFAaJgz4pQgrTC/O6F4NQ9aY+vlLYNs3yDBkPa7l+ZQNwH/L
6xwoTCEj3bAUQeYp3UYwABXV8OJ29dRt+D1y+ghKuzyMdqB7cuejgyoH97y5qd6doyJ4OIskvg+7
ElzEe7buvpZtsE5gfQjTr0oMkV1R/dfF3C8Ptdw0qDo08SxrRfxOB3XAJvXny1vgJRleAYqIO4fF
Xm6KIaeE3O9ebISpAMKj1qwTH5vlBGPROCz3KQc+vlX3MqIPbIuzJtRi/o5e1O/oJKuir57ufBWK
Q9R8BVAmDj6nWM/5SYXYVe9KiajEpZ413iB97jUWDTaq/mrHadE8/wJ7ctk2VIqoVcigQjIR0TAn
T5fvaDaJ2rBjnyySljUy0eYTplbCBcWLvFizk0+ENXiLs7LJuirRVsJDGWfqgnFcNmtIqcYbapiq
wpqB5yfEPS5fCS3bS/0MN0fMbT/TJ0lXH4FwFnMtP9lge782Aa6eSoFrX3ZLUpKkLpeEGU8LQHkT
5PwWT6nzly3Oeuj6qbdO0GCEtmTp3a359EYu416Ra1VamrXt+a1YcqS+0mOmHfZ5/iqJBHC+dQGU
ckGpnKIgh4It2+UMXNwsX0WZCYBC+e22g2PhJCUGjYq+kG5TNQorga/tZmEf+pdtjHEwExHvt3ka
lVM6Xy33O5FMHJ4hNYs3uTUDD4ZI4s1naO1VyIKds8ElbV2FvQyZWpFjaKkWOi4k9/i+HTTDvBNF
8e58Vcakb+UcgXtAkAsp+GqdNfOjvGIN3FBnUjEcrXE9OTmU1eI8uMc2rXwnhUqvnKVZO5djcsiY
Gnojvik+1Fb1PdOfdYIVCxhwHwtgNl289vUZaP7oGUT2p2NSVyDiOeBcuc3Zx4rkf8NrkIj/Xsep
Gvt3PuzTH6xE8Tqf65VVBBwvK9fv14bUaUqj0x0o2z3Hfb+3mCOsiucZCLHIZF+EEW1TSJeirybf
vmFC9GZ2lGxL5HPK9GNhwmd0Crg3p0Cj3FqJ+J+5gdb2IopX+ci3J4NjZLMnO3ipoUnkl6o2VRmx
YdVAoTVFrId+LYiSs62ZhgqItUaTa1wUwoVCaB957iPEo6ETwrCm5E1ozWzEP4AHPyUAajD4daqD
hlYvKCt+DXdoIhk8S7+pF1v7R8zJRvl3zAno3Yfv+fJ8NN7P6blifXoEbFlI7xxcr7RHSU0NgA78
nGF3/e+dRCvpjc+KQUaSCFGReNpia0bCFplHwAIDTCB7XaPThX/4UB0JyiLjtQ959Wdu6aWejSiK
bwkVxGgTg1CJ744CojlE/nI84ahI4G3092QYWrx9pgUDiFG4hQaxHi2kIsydt1/nMOP7MGML++rz
5fqrGCRcIQtohAXV2hQSZlJq+s4Sr6SVcnUOy+dIeDfimmilIN56XqdBGIH72y0sBykZTASOO9Vk
uAwnMR/K20fiHlx1bfAomG7cY1FCnNDAGdlEhfYiyOnZ7PBfdcUj/9xjlYnSSC40SX/n7sWr4sQ8
xSBEE+ogedrTAN7qzgmr9FQI6KiB8+djIKn2wYbJ26FimRhwifKAZVz3+gP9SxHa9si1TEjemzMZ
w/prUSRwIocWmhJgTwEJX0Hiwk3Z5g3U2Psdxc8SPNP2gxT9NsYUGTi/X0obj2d1sm1EL5le5fAT
6V5jVWxeZNP4hkY7BlcqqN7ltrPTBT8WCjBaERNLNMNdPwwOB+4BgHKFpiVdIhAAzLsiBL25wpFH
YAEQ8HhlxECOFv/KiPlPJILFJcdvMBlsZ/HVTaUs8k1OKRfohJwXXC9Ft2CQ3Gf+4TaiR9u4s1zV
XQtGzltC7Qyr8hol6AlaOk93PKIOM2/UGP5eVkzLm7iPKPbVIZtLkbfnV/n1WlJuoibfuzYA/zEw
Lis4oi7kcqtOj5Bco24gWc9mlGNrp9falZyOr7ZWQUFyqL84gQcBMkVNyk4s3kcRm6vhJIJLieek
rRG/85/eaPxEYLJsH+WvnmHfS5AXzh78Jzg+gwWC78Us4nZD3ClLFp7NYClmqphKsE0r8qepaght
zFer9Ysz5XPW7fHI0mBPNjDAkHYiE7AjRPKCDnmSW7Dm32gpk6bvkBek5S5gZ3BSS3CGMl8nvxbw
hHBc88+WtCja+ARBblmsoC9b+BenCgoqf4AOe+lfx8bevDvxpufQHuTFuIkk9emI9qeeg/cN5xcq
1v3bJ4abq5mH52KPYzvVS/95RqtUig8ZKPG5gphyYgOhp3+y5mO7d+6+IGcThsureOi7n8RRBeSQ
YC14jf4y4KhGijrz8/KJHZc6tMMTxAGUarIUyHO6JjSQg5s5pie6HDtrxGNFRTPLcHCAToLZpvHl
sYHHE6xOsNFIuvF91pmuIyOFs/91di2kfBRHDH5YTMwbWSCvU3mDSXQT1yc/lH+asUSNKwi3eWh6
FFxcrY+tl21/uw3dqU9YDnuiJIDIJ7lWqZuiiJXglnhBG3RiJ7cBnp7wz0wGUWYTkDgYTYmD7Up5
Wendp4b07VvI5W3Sv2sL76mFmKdKQWCavw0/mvRVJ7G+UGjgmtSnEBWz9WJZF2g6JsTZfDgRFwMl
qydsIo/2AlKwcHLu9R63GzTr0WsnHb3306ZTKPnIM8SpEwmOF5IIxBq778MKs5Hh0DavohmuH2Oq
QQ7Q5NzCOfyBiAZ9mvkbquhAFOf7LFN/roAelmD6QTh6yD51LyDTJYG8TDO9j8uW/eOMRNAXpZBM
sf1o6c1/MxcDoP10s2wrg+xIfTZLNtOyn+/1o24MSNbwhFb57p0kehrNJrNwxGW0rWLFhk9wxvnA
ssiShUpUl2ihBvtyk/xr7Xhtx6pD1ejGQxGnCu6PNQcOcz+8j9i2OZLxzMwMZx6c5Ayn4kJ4frvO
ftn3VpjxMHqYJvCpMiFgSCd2sLAxsIIA1DHv7JU3VSq3HIZt5Gen5CVru0JsHptoW39JTdZOMFQM
dBZRBGmJit2+FNIZJQKm4KKf6ju+e0/YeFrYu0N7aa7HdoKnb4jG9l3DVqDxxil8lqNASElDCdbu
pUQrXSjBIa2GwvXE/3cKa0+0MC6qBMQAhhrhlFJ7xvnEpHNYGt1vKRMrEhGNyOHeuSYI4DiDV5Lc
nWzLZT36nTL6nQNxNvmnZiJh4Ezjj4PEGrIJux0j6zej8t8mByd0+ZFxwFvsspgIx+p6FVafWYp+
bSvZgRGO08P2dM9CDcdaS6FuS0U1TXatBH7nM+7tITZ0MTVUSNyqDW02v3mNyCdGb7OUo+BtJHzm
+7H5YYeY2iah09aCd5hw8waGm2qYKzfSmsXzXJX1HE97Va02R+paVIZwu8/gQ9/RHvI+0gJu3+iR
K5tNDL/7xc2hRHENAmsfbKcGjd6T4+U/rTS47XBr4MalPnwY2bh+FtR/OT13vNRAMfg3qsXykQcW
c5HO7jGgugKyLgVS9XWFXIJRlXxMSrQQwCyrlFarjC42OshJJy2DZWpOaE/qH4REMjS21Cyyn6aX
TacUpAgzEUcCqb1JT9flA36GQH/SgdEJoIaqgi9xE4f6dtmwUHmLp0+mbwCzM0+TupQicFu9gLwT
Vlf3lyS+iz3ozEb/RCDWpasmkt+Z9iTva9Hq0zHW2Jmtx+2xhQxiUqs+QV0gdo33F00TiO9pZkbd
zW/w2utzIWmwM55WnIypBbi4mXxK5eziW2D8LHGNfiUc1E/t6LkjcucMBSCmLBxmljSoWV7I6Wuo
e0LtEUqQq94At6G6Br+dbf+dvM54PgpVWH+U4fGAHKE+L5JPBH/1ZyrhR5AGW7b51QdpnkVDk6RP
X51Q+PJCJAXoRQzaWj8g10Ff8T9MQhYwzTWtkKVC2LOiDLTNdERK6PW+E6HDcBOpxEdOgeFMeN8S
ojI/Xru38lEqclmpZpg833reLJOG1td8CY8NVrTSyacbL2hThSGlk8/yMrJkLQpL3pa+zNl05f/h
7SGmNqBGTSLMEGdWmxGT0T3VBuSz/O3MrctcecEMb2C5eYujnpUidxdUxlBSWakTHybKx8rVckGZ
7eCOJ3qUCm/Dst9HlxuUHjgikSoRNuqBjuWH72mNX2BWX53I/aLLH/qHT44+n8PKy5JmTGgvME+t
oDwjL5oCVXGOq/r29vq2cu+EemOcmBw+R/k275oloEOIx/DseKeHO4hfTEaQjJd8ak9Z00IQypw0
gp/X6aJdyKLNXrZUu34kGlTeNc3YPWdq8iynBVRISpg7O7iyUDZ7WX8IHjnr43o3tIbTi93bdP2v
H9+gz7Ufx/TEz2V4yd3/K4G8GcGEozDXQ7MbkVQTwPzt8t2XOf4WkXT9qleEOCyN5alsq+F5Oj5i
RBf2kT6JCd0PTLCsIOvpLHfMcVht7kaRg/2W656sCs/m2EgH29lJyjXwSyIxNHw65nq/aypKy43V
eSpF4YZmpONg0YBOqIqyClAoC6AAk7KATblnuuRE6aYcXSHmfJ0xJaYLVcxikPKvGZ5Ure7QMBJU
YEcKiPn/teqwe6vcGiHG0hNkhGz2yUiAXrSSQl95HC4CdSwcVvIi6rUqHAAZb8GkdaQtLbbtVdP4
DucaYNzfRxWLmW89GgphCEvHJL+/bJLdfw678zIC/SUj4QmyWrQxNx4R0H2aGEQmVkxFNqqIwzro
JcLEJ2IjjV+5el/05FtyLsaCdT2V88/zgw7Vx3HXHgXC8zNCt9TP6YjGpBwj+E8wSa4dxfL7zJd3
2xnMHQ/MfEE13ycLlCTELwfLYq1g6LHxkO5Sf+LRiA3tUPCl+J2+gRhJIS8cMkgEwXWWRjnHNP6s
d13xmgLVW7D2kNz5oSrMSZdum8l9yaCYKM7tyUKbATlN7IfoggOhEVV2SVUCeOpK9HCMGzMxj2Av
O8PF42YkLDFoHmpOGOzrEP7JZOpSrIVVWza2zt7RNlO9bgBDZ5gsSXd34IA53xw2iTDhTFtaHOp5
7bXTVZpBuiAxRZXP7S1a3zrvuU2qYYGNj0H3Huu9aT3gF7UmO6C9PcNhRPFiO3cnrbRihQebg7eo
X/d9DwdxRxvRnfOvp/R2L4/lqFrnSxhQOEBwJNsMp6AuAvnLII42xp9rXMAPscOqCIyecQrkSmZK
T4ooqn+aZ7Pe/NnG5amh251/4NJlqgZ3X6Kb6srhxBH8yOjR98kvQGhp723g3dJyKOiybDdMKMZC
I8IBRgeyCaOXZ5wsxq8dT70DtSqOHQRUcSF8S1pamNT1g661UkHh3VPdsa9YDxaDS8tU9QTgomWj
FQ7R0r/Ah26em48ShdwIyChfj8zzecxqA9dJIP2Ij9awDr9CYF5B2kgQC6UGposCBEutxHSSDKPE
K4wjmA53flp5RvSc66x+VDiv3dZoYbVAlBRyL+oeJBeqZba3X1GaylvKS9MlpUQGp6yWoEXjMHgM
qDUYbi+hEU+Djj8QqY2Z9Vw8ftPi3ib3CcFDJ9DR+1sNGoX3oij52uQTz9N3nAZjE1ePWwfsFkqo
HXGJpj5rLwFs2DnjlSPGNuUb4nnt3pP+ou+IQd/A7zFIPV77TRYuPv2xQ/OCrfp7XnUNagPP61aK
pp/IgV8N9wfU5r6lx64NgKGCsXoU8OywLNMfCByKDk7+K4YDXVSjZE3IC+SG7zeK6tiXm5N6j3f2
OT/NqamL1y2W6mqWGU4ZagsL05zcyRurNKcTe1BIVAxrNdbjF+7n55bNPJ6ikK6qtiyYZBd7Z1PJ
VHpJfaWGF71Zs6vxx/ZhQuB8oL9Y0sNurMeSAqeVAvvHTBD40rSRPSvdC3UZ6FFU0r3Xoqj4Sdtk
q9oSnOOOHaEW6QcXQoezouqkoFQLcZ9qqjJOpAXf881dEnViBwvgWjmqoucWdeRoJpy3uHAhcbFT
X5yHUhGR4sMNTlst9R1pX90HzR7HDdGgsw81IWmko6Q1J0lq7JkEUNNZS0Os7mJQoAyzUNMX/sRF
p6TOXLE0ooMS5j2OUXDueOj9ccXTyzkDyU55ZA/PKHu8XZ6upp4OkJwDpH8i3Hxb80foJKP6VKwz
GlLVXG0edoVegDIewpwBK7eZrxIqPWEkxinEw5KMmZMSoZO39Lvfv1j8pasRStHK4POUYjkYQbt0
sr9H/Ezk63bEfA1C3Az0STaWP/TInzzMAiH8p754Z9WW8FuEdFWcE6nmeISDSY3J1qO50C7zPC69
91c7w0qL+e0udndzAvont8axJff4Zc4AQ3z8SWb2KvY9MYMl35hB7CmhTHWSY5THcAMxpv89qMzr
Oml+B5/OlGxuqsK2XeNKTXi3V4nDqKhIcRsrkrjxbjGTu5NNYtPAU1XpFFFnQtSSVigL3bNyycO+
sbgP89c/aXP4/cBYArW/RD/rRbldurkiPZO6d1F/YH4PJKoiqt9dhuP5ZTpy2kiaUwFHFDvhbdDM
gEfARz+mW5SJCBzC0+lziiIRj2gtwuZQC77y3yMFSwVOqojHCzm7gYD1oEhwA2PCxjZgTT6KaVFz
qDPuhZqTXyqqPF9rjNbe3/j7QhH6zoCaTUGchdOUO/fcH7410JkhwZyFiTG+tq9kQb37rGEnQm2C
tmJ+m8ZgDzuxKylSSKpxAFOQQs+O3ysmQFIEfaMnjHpM1BzlwIXTZ07qV2dWQBS7WNf7vzOl+s7V
GRrzpVhNc0nG/0enkdOoB2GCfhSdmED9txBtNUlFo8+4DogiUdVzeqnube6SzGx2jBjUOCGvkgNX
CwUHKmmsJYizZGgV0us0mgTjA9dtcUk68I1+HGoGNT6SCVoHdIGXqhfpU5WiDMWetRrFUGKYJLnG
5PT1DZjUCPZpbXwU/ze2d1GEkHHIhJ5aUzHVYxTOb4lj60T4qi15JzYoNWwg/cyuaSbqKb9OR6aI
0czyyOZRso5bOzwSkn2YT+/40YhdxA0iU5UuJrPilOVpfpfVtyDcKE3WlmHDD3KEZB4+ypqx8WLp
1ZnFnEyHksvc5TjV8NIkgBc8ZJi4RHVB+R/cOblTWxq87DUfpjBd5bmZ9jqqOFoyRHKG6mEiJY6i
fAKiXkAD99RAS91i//O2tR1utM3XYF6gW+WG5YMQ0QQbdOlvn5IaTFkyVv8oh39Qq5aduK7Um8Dx
DS7i8+MDVzlEtLGMdeKv1CulXs1/ipwmTZdp3LZ8+8igBqxooj6TWPszzdSnDMVl4IxK9r2fzRdy
7r5ZsdOJKATF4NC/aKvs2G9/Rvv2D38IvD9QXP7p6iZjSOb4DuaZtW1VGqsFy4FZ1LJzGWcCG1nc
pIpJJiJvUqGVZUEwZChPg7b0PB9ZdMmeyeE46gFuDGughEdAkPkRFslNa8i0NjYIKTGcl/S+vgt8
0VNUah3NhGqCOySAWfATWx/5PD1hLY1FqZcqezNG/ZXEjQhs+jXMONGiW8MIieqY1GAnRuW62p/W
LwkXZV+JlV1HFiYNSNBmiv48HT2td94rSVFiDBwLoX8P3gkRzdXhpugFmWdxir5k/0rGNGu/S3Wy
oMtQVoYFUikCCfo0AilR8aQ1ZR5iw0e1aw4K+Bxtdr6MSz1wmTX06xJli/8L+Bit0kHsIo7JdAkk
zdEdF2xhk9R8LKulWza552jjhxfDeLH06ff3Qch0KgyDpVmtiMYriQjiprDVrpxK30k7alQ2tk+H
0DtOpyqETZLgs65NRTfbZqAtOdEWt7jFXS3XCT7tVocDpwVT9RjcOiCW+roRKQLZd1uOru2Ix+UL
DBJP+Utx87YbgQ08DZqK0Qqj2nbWM6dv4ij8kAW9U4b+oarH+zC8pPakx+lb9oBxqhTTZbS1EbkD
55zwupvyY/HpZjcvd3b7Ot1S6gecqn6cp81n/LS1uyyOWQxlJhgU929faxM9ecFZoJPKIrImj05G
ydYdlus2t49zi0giJAkApanrb1AWOyLkxHwOHeA1TxRE0axM2VKTSRnne3bx6kBj9qjUf7KMWhe4
eOcJpachYkBMBeW1IqDM03PD8if/X7ZHlc4n5aycJL/3ZvjMK+H4MaATlhCedi35p3iClzhHlS+H
JjO78RtaxYPKLxf7YltSfQiMI4A7u1RUH3Q2bfwcMMVJLpJnFi8d7U/lebEcLn1OsYtbBPMkUoD6
siATPrh3jtmbZW+tr3B3xIvROrOGDBMrKNjhL9Q0szgRMMegw2KVFm+HlMWXQit6zBxhzNHjApcm
+kj2pIDeD5FSod0mgz9d1WouC5IFioJXFouCSHAiwMeppQTHRvT06nknrl5FAe1602XdEMRa86CU
+7Q3ZN1To7XfakKZkEEA1TeUzWLnyicL1UNZq2BM2GFBpVqoR7SpPrzgh8ssf6GBE/7KaY47sVfU
EouEqkNMpdMcvtk3h7b4Dop5qA9lbyNKxINI8rpSo/c8mn9AfWDzjyfFZrhFCGao0JwhcqZoAPTf
VLgg9xVd7LlW6la53VrKbHPvR/ocWQT6QVN24tl1jE1Er0Wf4yWQuDEahCLwBZaa3CIS5LRy+nWj
aAoDLr/jdUJ9FbNfXswriO1fSe11AmH/sjpU8jTD9uF0PfLj7y8XRNXt6zPqPBdBN3XtvCyDF7O1
wXKCqKb6x1vfeo1FsA66oi3k+oPb+9bUiB+e8GQwzu+n7M8rTjzOifRYUh2kP0k29u+jTPbJo3QM
50pslmSFrGLz6tspAOD4aPU0gZnOYAF541CmEhNtQtwOoYyRg8raycBdrY7A3W6jS924tPyad+wF
PSmClcNmt5vv7qR/F4XS5INC8KS6Sb5y8jylzlsbeahC0F9HrTHaCoaKDAoaBwIf1E6XlNQ6yMCZ
IyJ31gVsZLyPtCmla0CNBZsxoegsz55iv6keZ3C2cjPbtYGdNEOQG5vcYEicNiz5EyFM7nxeY7y1
itNvOfMBHpNdLIHjZs575fk8dgMW2fxM2gMxTlpq4rJp/z9jm6ykD9FkpXt/u5mQ8RfnqlDCXtxR
IGfv34x4i1RR30/4Q/B3MqsA4fb9sDM6F+bfn1JXzPRiFtFxXa1CY8sArmSi8bsLxW+/tLkmyH/2
oLe8/TPbNREsbyXMW0poA9R7P+Owz9YH61C/2AO7dmN9drYa5dk56KnajIKflxbvZquh2A/Pf2hW
P2s2K1rfR+dWNB7b4a8xWlyxmioomImjVvLtcAUrttGNDYl2GEyPH1i72+gXdniqrwR0nJR4+8nt
tOMlU5ECS4cErt/olS2L5Hao0CEAag/7p/25I0CeP6knmBv3Pe6YFgb0aJ2U1SQDcqlBDqJ5AuEe
3hA9CPQt/UdrMQ2Wl86jqocfms+yFpBBEZavhEm003+wW82dWernGktozrp/RJFN/8JbVczHL8zL
UzAh2Y/xQWaOF60RVoeQwMPf/B1pLYNRoWVHKQfLNtugIHCe8Oyfmb+pLL9ga/Ppcd+vP75m+q00
HWpHRL1TNOudgQpsdKSwbRPLxhY9mJYv1Z35awNR9IHSwby+WZWyudbFneleMElYHvWprVeAbjvT
fTQtDHp2QWxXIxV+DPyArfOdooO3sYecktgvu9ra6aeVZgfIm7CQvcsi//OhnoJ6q5VVBP8Tid5x
i4kDNYusvRjFvqtY5jxrsdgwJ9cvGq77DlylJnVxYJXclRPxpu4OF/izCl2Yh3GngfXIDn+0VGGb
0AcRogxmK2G6p7LCE5j4lJsw9+gW6vx82AMaJSBJZ4+ReKplRhCKRMTjV3dFoeAkSWlG/BcnKCmm
Sl2PuYiHOOkbgCgA4S/2Jhh6HUVzR7vWq2VbvYN817lQnVfLrO5bIWysZtqcyDFNLdOh0eoy5uMf
1xl2SNpiMjWzom0QReAGeGWrgALuy1gRExyPQ+Pwjyk2TK6SK4qippYbuTMb/H8s2PPN0qQoPgvx
V8ApPDqhxqYA6KEje/qrTV0ctM+qbs2H9QIFxYwFsWmYhZK9khPSUj1O0GyGzVnOMN7YoVOgubJX
cdRGC3fi3DK7Zaf2tMPb7+Ux6S99ViIKHNTohkAw6UVRSOelY/yXRjUjYeHGDtafSGW+S26wt3Qy
9k0YGdEFn90U6WgNk3HVOU+jQzWkwUE3qSvfxWvUSo6E3aXCwJvARrAOwZ9we8Jbn4ablLa6QZeL
8lXR5QiOAZg5je4HjbzF1NE6v+0+0pfPaCylCBiYDH1gKD9ql0O3TlU8ZssCPdOdxstkhaK1IqLX
pO83HxozBvyztvIn5Uz4AEOtFLEEE7nSxITrpcsPm5FMK4HLWMt2M5GnKO2vDSncB9HZlGihV8Mu
BunfOwHA6XEJq3QBvlrkTxA3bWHStvUdQJYUqVk83KLSRC4TFhWRWOpmBwDMvyJq75DfthI6+MTz
iqgEfmV3xoPvdzxN/PGDL5hjzB2oFxqqqU6fnexpWCO2yaw4NCLTfRpEnhk7xV56kk592vUcqJQD
wD5l7LNo70F7yarAc8OtcGYo/Z0V2wRegg7gD3Lj9P23E+dSTR9UXtEfpICGPu8UbgQaNevfUbMU
M97/Wc/SOaaXbQ7AZRpnrV68zjanL/aHWm8Z1/LWxM+LuD+sw1mYwEKyNlvWtwRBZuOi0xCb4iWG
0ZwCuP7AyKDzyRFR4bQwuenTBB0WPQx1PNYnUFA6L/ULJ3rqsO5ooJI0pBnjuDfhTFo5laDKrJdg
f4Lq5ylqD7/xWTFuMOMy8cei312R9GtbUfvoVbXyga25UG3sYCnEKY+d22d2oNgjy1743P0mCfpS
kb+fQhbQVJCp6p8eLsshrns5NZJjgD8kAC6ojDw9fgNUP4B7GI8VmBWsvFW22c+Jd7DPqWWo0NQB
dxLWxvCI3ZzrRYGZ0ygHvX+XtjXQFb7vojYYT5RTcUAZnoFsosWrPkOmkoX1a/zL+un5CAfCoGhH
flbJhV4IWDA6qu4136hY+oL+q1j1QIvz3X4AetbgbPCh5YVoMi5XH9V1CWdB6H+OZF9yvpygDLEg
XNKcIbzmyxjsOUxgOt5I4xduL7tAdSndAlTZjI64mioz2Q8QCl8x7yj7QruWlTeZ0kjusg4DEJZ3
K5JVk1n9pprZ6iHDD7dvrUQAOzqp6WCkasQrjrZoX13V4104ADPEemfJR5CvqvKvtGLRHvQ1Dtk4
3mQaK5MdsCN1fN9UfyIcSN3F8+Sw0MP8IFvSpluIuL7in58bJgCRUmO1hDT0jq4cymvhCDlNwVZU
RWy1Qbabk3nPJtYRt1M6AvyLt0wusPXAi6CZ3DXBaLnSPbMYUA4R0ScPf8AcoZ+eanG0380Gio2a
IYgDCfbHUEbd0y+vE8A5T0HKEkAI5GpS75MjF+TU+CyOUEdEZW2rWvKxRX7gCh+G5AJGATaleCaF
Hnv3TAeOs0Lp2GQrwvq7guY5osXN//iGgqv7cVPQdX+7AcDhHAfIzRGV/FnEN3INIrvKQs8J46nE
TRdVSPgTJvMBrYpxH4F7CIu+N2a3hbpwXMYV95r0vbFFhv+G13lTGvjqqjmTFG/p1MLDS3nPHqBP
X9q7fCTaJ/3VMGymEYOl7wadmFvugNWWYnW86aCFouVtPUx6nqw3kc/qU6EDlPi4ZVE6o678IDup
IX5rzN8M3hs27fHlOzRniJrG/IvSOwPDVSiWv+ChNxrrQuc4RiakARmSU2EGwXnft1VMMzdTz034
8Qe1Tsnld8R/bdMCsZyP+/Nc6T0EgkLPC/cGmFns/Nqc/6rdlLujB8+2fIH7vb9PBsU6Ks4qih4f
Nv1YDpt6lNkrdWSDJja7ubS2bgk+0PNY3Z2b7c7yahN838jEDebOjI28NSUXLKSVtaWRxGPMIJAT
cmFZCwajUw2KXPSbuGRqZk0ORgdFm5OCtSu7/ygSmiKc95yCiUPoL8DvR1uoF3nNrUePx5b2ACrn
VuNz8bGJRhcnzMrm80UPthX9nshrutFl/4x1hwfusJbPNLqRQC+1MGjGC1Ga8LK8tylEk9eP4pgO
AgcKDx0PGArGk4QkcHy4u9wkQKukisC8lkYDNWmiOxT6zRj7/m0XQ0I0oTakXDrKp5Bx2rN9wJ/c
o2w4U5INpPui+PIaw3CVg+YMBFLcOt+9mKHIIoC+KN0yzJ2UDoyahaCAmjtBS5uVBteDEwwKeNDR
ERUVyQyjHNbBmBhfCNoxV0NvIHogPGoIrHtx7GjV2oX3Y3l4WgNULB+1FbOMJAxie5OucFAstjAh
DEbau2rddPbFeFulxG518v88H/SkVYVJ4kZcjIZoVfIxTPTE4c65CfVq5erahIAI3qBC9vjg8GkP
epa06o852ezjpx0vtHmH8MVEGK0UMQg2V6hd56mfGP0EKinsEkDQ8eume3FavYFAll7WKrM+H40t
TmdctAAVLSpafP4nMypO77qh7lUH7Nxn4t9imLQPa87bEQdB+p7oan4FlaxBgVL8pnfTsK78/kkV
7xaB9kClRYui6zG+oWOk/1VvNtgogFo31lJfoczs9ycdhpujRBRV/hizEeNmoxYYplGfo629mjwM
78qwp1wKyO1aaMV+aIYa0xipT9QI8Hn0+j+STwREw2vDxSl8T/I+ouVNuBTPU1wnMCyqOeZ+8zHO
dNTlYpf/Pb1r/q4UWYRYARAL6xIuRLjxaNOtbi4hEgb0eWH4cl2528L/7oTgHqTUtECKMlaMqUMJ
aYf15zXAtgCjLiKCUiwBxS8D66fAvDEOCy6B8CuHtd0uoKaz95X6kGIVTOZH3o4qgZHZWbie+xjg
ewQOPe+abGrWbXXp5fU63hwfhTjfEcDi7Eh8DvHAtqa7RS7/LNOm9Nzz/HVXFrhxswh1tW1VARoL
6DiPe0WPbIej+DWW7sKaUtjogIL5ONbnLBdQ7LTYlv9GjApn4pMl5m2yt3qBmdFDCfnvwM6+4nMJ
zQAlYC2uMmmq9l6wqb7wP3fUXtDrKaG2ak1uoYeWzcUsoQGd6vjpVGGnSOQqdzBa/HpVDtkRiUHZ
7D9qM9nY0+y19hWNcfaQ5fbLvqtMofSWB+GixonStbgPkRUKO67dfGIQjvXriiOwT9Um1L6Llgea
eprVlQlnvaN0Wnsq6f7rRsDWEZjn/3kLpZGQSfXzM/shjeT+a568ZJp+8U1nIiNUkyCgQ4jFR8ph
9a2YANnARAtpBwkbZo3/LnPvvzefHNK0sa52uSx5+qVH0pZxEa7IgsjgixVmqmPLHEV37OLcER+W
wR7biJt7sxlIZXR5F7ME7rHYJeCwqHVI9ldfBG4VzERoYBseFm9T/E2lD24vtVpTydpgoHG8sNZk
osWrd/fp6JJ78e9f0SQ2HgVNmpYosxLG1n7fdT7TQ9QHzBBQDmXSXtSClkI1dStfHUK5t5HTXG4C
JpQ9Xx9CK7lkElfU1GiTj1kvNZF1ncmGww9grBtI0Y3W2L/7bEReGIpxeaeuQv5mpzt8mP+cnElM
7InuyR6n0o2tf7e+6C3J2EgwVPjwdfUCa2QLDJxg9lYyAunBxJCyELKNVM+yi+2oQ+Uf6qb5Xv0i
43Efft9uBL3SrcVTZKF9qPSItDlVLBIaQxNjAwSaLpMjsyJzTbH/r67g94t09g2DqVRQdjTZE8z4
PN8R+D0O5xhozOevF/DBXLCeyfiGUBxPsxx9CwTbWIg458X0j4O39S5rUgwy0fXxMs3AvfRRswuL
FG+7UpyGfYuxXPi+4AE7o9q+/XLy1NoJkjjZCYi1jmC/VKTzwEnoXSRcEAhjsW1hbMdoNPEg7VBr
D1YwuZqwwiOWZgaIDTtEjxN94Kx7LA47wUXOFeGFIQvrbBmNTDcvY4SxjpydcJizOL64AqtjkhYa
s2JQX0z4+WdtHNM3qCePToaWRcsIkQsru8ujMGGw+xhIr75hj7cZ3Nxz0pQo01q40okC6KpVpDZI
xgRrISinj86XZh/iWApYVsmfYyugIHAdpeKCYt6qrZu05ETI2HTNnUT8OZBSkA3c7BdF7kOdcH02
6vF+MLYJCHN7tqc8xwB7Aw16SiRDsbVq4v+PXEfQmZ9/GoHhUnzXBf435bPx2TZhWQ24eqozj2hl
/715oYxqDWUBSkJMNexevtmcvuWhLuK6BuWspZcG/xHO5Ncb45LDtFxQrMb4ch5IxjD423gUWpcG
gy3M2ukDzGG9s97MgVcXX/yAOEq5ndzDjVP2JshNC2u2Wly2LJDI+KRMyXayEAWTHNQxI3ohb0kg
BjaPApSaV+YiDFSO64Hd0ywgvO4nWRAcraiH/KjPXMTCl4lLhO/8zamHKURi64hr/uuVurC3WPT+
qzWcUPIbjBJ3RFYoGxanooKKZoFv14yPqSkIX2rbQb9vEIRlnrV7ziobBMAEmJWn8qZGMJPFWsHI
UB1z7aKCwKJ9F5CYkx3cilEdDyg0i9dGByy/hSB5WWIAgy1jxQRWe9nfyXWoPuQCsLRQvP9mu9lc
61xTCEMRlZ6Ix8zR0dfl8dAyqWzItWAYqJ0AeqgVwe4lTn4m+aiNLg6eUlTlIGAG/30v0IdwWaBS
+eInOKU+CPVtZvAQqewQ/CA1AVuKjrn9iRwFuYQ1Qx7hASFYsce9J1iX5NbxWbvlSROsEMBqup24
S/aycUgl+O0RxVdq3wpDVijLKTWv9wF0E16hQopBxv6oFQHvAaiwE7bfUACxx5UIf7WFzdvt8qhq
Y1bXVNyybULKcjhmG7Xxvik9WTed5IFWcY8gMifMFAxcVmOyFTM2LD6UXCFw/FfTbaBkffftjnbN
QwHJ2lpp15fISC+ZdZqLZygogyzE23YwkaWr5ERSoxLqO901FHB9XFHKpbaxVdBMLSWzgnxGxJ0h
6OfRlVP8aAs/UhsWlWjpFR+Fwv2dkz7pjTSwy6MpaCoc8sllHrlsgHm3vTRn9dS6q6IMxn9ADZ9+
30dAkq+vtO//bdVwEluiXo2P+Zu/s2xOi35v2/UBgobilCfB6rZknq3qaHPHmT1mZ+cUVIEfVgCv
OZ1eJabnoYe/cz7ShkNKYUMbHaXLxAXeFrWSYvmLaI6m5Mksdle3kFDU23Sv6uDwsizO0DqRwd3I
gbJ4SyjnK/BLpko/k0LsgfVR2xGc8klkK4zONvW1cEa2dAOuz8mr1dyEhgLIsKHgto4jBlD2hkBS
CKXiOImSF/zPN7lxkCK9nLFm1TbGOM93xdPlZOCK/8RgOEqRY4NS9NQDMGnRVJ7h660+oIXPfSH1
pDezIzVIlJmpnR7c6LBA0IcP2s6ZN8dDDw2RPe8rRlAJbUBjK6EPeTjHaOBfCgtLEZ0h4fkTPydm
8Fsqe+SdAm+Vb466DNsT/yY9Kh+PIQ+FvCfC81ifWaRs3Wbo3Szs9c+pBS+7YcZY22cf/n3X5mU0
xjAksb84vc/uyo+wScsZPj47lOrlKnVnTvzHldH0rfN/sVX0h24nJDfHisDO0jTf2CYE37G+Lpa4
zjF6Iz9+nC5uBcZ4YO9rg4zuLOux2ixhDpdFLNp6zj9lc63lGNjHXL/y+CX/wAxN71X6RVJkMVhO
7BCcBiURVF9/6GbfyUa7br4+FsTCWZphEJY5lhptbdF16VKd25Xc3t53c9+zEzMgCi6e0pP9+/sZ
cxBXs/bjaw5Wn4efDYYbv6ftfElvFK2J3PHfKqEHnb+wndh9ykF+VQmNIEWA1grYDGAtujVjwwE2
7OvYikWEWb7FygRIz3sxBXWMs2YOeFkswNFguDu34hJM5rscp6bSYezCwY+LnmfcA/OSlJjuNRf5
nYK1sFstz5N1tATdPRcjYW+VDEOkxR6zxuzFCMk3YTIzYLU4+c/k5lSlXcdptB6G314Pxg7v0PBh
KrP65SLCsOKWT+6JXhxtEBdH2ucioizGM8CDbpI7nMT4q8WKURcyFWsAgsLOwpjm2rfr6saJVEx+
wCJSeVpBWYb9IPpgcZS5eIDn6M753fa2wCACvZ2kVlVwpHc5niqOwWgNeS7dcpY9MpACjz6rFOXY
vpU9KQ1xKyCNpdqQ5gdxwUw5zj1sXQU3Dx11Q2sne0ItVSCDoIYPEVuqtbX+aZev9k3Sktm12PDP
L1FhIhRZ45pa0la6EZTRAOfsrgtnYylJgGkHN07o9kr8/TqclMmFVWqd7hIzbIlMx8/EPcuoaY1w
MXMVDZjtVl37EkuNt57vGgOBsvqIkQonBzi45xaxSNUYWWiVNI8B3jBfU5KmDLIxJHiqjLj6OVyv
JNAfvYv2O2WDLdbKF6oUy0IUiCoiGIovgzFLMiNki9q72dvWLjSolYaoprB2FXl4stzF1EweEBgJ
JyTUkGWfTs7laYMXo+xjp/G5x3/XjTmYt2hEoKZgNI/PXKYU6ayAMHLWd3oXOl+E2TRMho/3g1eT
L/8dFO1ZvnG5B0hYMfuUrHCHw8sJrT70V14zuF9DBJTACWdM7BC7TXeXv1xhRKlU96qpaUUr77/D
HzJ4tFFbPiUF8KU9UVWPT3q6+HfkOC4aVQXEYeiZUbeiadp6T8odf/xZa78woTQZuxg1QlCo16O8
2EGsOP3x8M0VP2Zf2auvu2UfA3b+DmccuO7LWMQzdA5wTyqHQuM7s7ElYkC74vx32SIKD9tyeo0T
futiHKgvaSXmdPf+i40dst1WxtNwS5KJIFZjREClcQjxnlL3SZfDEbDeNLAA10lsdeoqna18dJj+
SPWhh/P63FbYyHgIVb1PciMNsVFOxhA9bgVJMZYoO7o3TNwRo8T9XYUYatZGnqg/ziXiLuf4deqU
IySutMArn6csVK+M8pf8nW0EC305KBpJcGg3f+wrJvGTpGoDhYYP8suqx3oQfm4rDZZB69dLXyhV
3SazutoPbkUasxEnAr2VqudNvv/DCv+qjRxb5fRaDngge/KC1Bc3MAnAzkHdtwC725S8zibBwyJe
VhZ+42Po0lqT4zAS74p0NVX2m0zoUUglxlOiWZPI9rKW4VHHuOf2K7XhS/Ns3aPJeZlN8zvIWvU1
/K4PgVC9MLj4UfrKCgv6g+GCxtAV1PehV3Cwak0WjTiQmw9e7eTLviH6KRG4Fc1vIk3ZwhBc9l0X
QcaacEt8+cfxuoo0ICfA1lkbe0AUeXvG26AcdlHb6IsmFPvhvib+2PgtsaAp+K26ONnXhzU8BUVg
GhrF0ScNZ+o5TtY6FmySFP4JgLq1yoEdydeVeqNexmgf8yAfs9//6/imiNscA3yInr7e2Tqescsk
B32q2ObAfh1rGxSUZTp4jt1f35i61ExtERRZhysBZP351u0VxrHKGY+CAIR/YTy19mwdg7PkCDAH
VeFcbKhVkt3ce4QAERHr2oOjz9nXYd0g7q1Q/7oTzbvABXXq1VUQhxfzty4GWutCZiuMSOVapUdd
OXEFkR5+fDFHoTjRH9Xz3HchEU4GTX9TUUl/GLR7P6mm2tua2Ox244tRJIcKxEGwzqeWaXvuuDCP
Z7WvksS5EBecdHgT/8f6WmEHtczKWV9IBSwodiTitQw9oDAWHWfgkltSp9gfm3zsUro/iH5xd1Eq
LegkBhNdhJzoqmgL0yNosF5wtDwQUWXbmmhr2jlHXV/rh+Q69/DQRmQPvGZhsaiElO/MsPYXF0yY
Ldb5HU9SG7BnVkfsIueAqEth2bJYVsf15jRqmDzJ6E2P4crr1A2QrMqA2MVPF1yXYVaOk4Wz/UOg
in/hLXzKKtARErsOcPAEQSHrtYyTsnxZjY1s9cek/fj/bD9dwWJA+Bw0EWL7a7apZqyEAscyM/gL
ADu2zHQB/EHdk8uiDTEIqAG+yNwyNStiJY/kMghIYF7FNH5W6uNMzyt0FUhn+qG4L2F9BzKm1JHS
7flFGNKunZO9xi8q6i16zuaIpCgZFyyuohHBqrybemZcaLP9mWh3B2Ua5LJ1hgN+gamnAdAa74G8
1LlnpOV9piGz7b81rsisvQraBUE1LweSsSr+YZBvVx5g+Eg1TNIOlTvat+Hr3QEAmONDQhKSGUMj
NVVDyGhf3EiR6YCmBOv/cAZdnYD0MnZdJjAWurBgI0LPWC7MsNEjRwxhg4saM0yKs8dimlDxzB1Z
Tu++SsOhHwoBttH5nRoqG54jiX01KhrvMLduM3CNQXFKD3eaTVhTgYLOwaAWjH8wL0Lw8NiSDker
T6z/dweQwgSqqhUxxwECvH8fMp4Cj/QETpQ5TIHtMosXKSzFMp3xRvnz5oPMfgwX3/ZPKR/fWJy2
wf+wNazjLcvSD0m2BmBJPfs30ssEBJLzIir3aatL5Q+5IF0DzvcCio18KxPgGJJWZOaLFLUaKEGJ
7vYDYq1GY3LFaFx30dyJyVthgcdgP0QfL/oMcd5zCH+3WOucG7Se3b6rVXmXegLHXwUqooK13j98
u7iLsHzqB+DkYa7TI+Ve2xcYtW3RxzGrStF93/e7LMegkzJIPldhO440WZqMruMycKSERleM9D/r
wMbBT55NR41IkDYVu+UK14fhPlZoQ1dQB1+ifWK7QFrSM46GNZud4EuOSMpn+9PEy9i3U5lLO3gU
qOFfHpKmLbTlEdEU31et+d4PQ2lkyuIIHMFluasHyiEYbhe2Esd14gJBgT3uMQgEbJoWyAKxOgmn
GC65q8j8/fNLFI0If5UPmH46vRALLy7Hn3a/0XaX0uZxut2Gu6IhZ9pJ+V2KAdXmwhVvLLlMC861
ODMMyHt7A44QwyHLIiS9a7/Mkt4iJTDHIW+7ZvNyv2dIlqIjFU8qmG6eF//Kqcb3+ULef5vvR74q
d8WGx8wADyb+tVRnSmOKH5aARZVk3u2xQQ0xSJkkOuA8k/mPkU0HdIWnttHnyJDSFkVkAZ0GpQh5
yY6PaUiDT/dRCwXe5SJJs4155jnEFIVVnZgHnY8FORt7k0EUQaET5Pw8sJGVx4EmmPbpMkQjUSTz
uxMO0m1wgQBAc36nSpZfVqfSR0is7fyvEZMeBbZ/1996zn9Y9o249paqQN72JG7tjM2AIM9ZC2Im
SB5RHxyOn0uGrTHyNeMx8tuCdaJFNse0PWvhkJGoWNJ9t0oosCxL+1VYKWQ6L8umiOevD+s9zOve
X5DUd0a7E2ldhx8uZClXyYCuo0Clgc0ZXwJtmfPxA7E0yRYV0NTKbaJuo54fLGLjFPVbVFM5RAqC
p5b2w1DREktPD7wYGcZA2tlWRifGO+1/uxpt2ympJlfbDaE2qCoe/22HQTEwAlMiDCTadYPzUkpm
RpuoulM1XIv56GoNNvoMh7Wqeb2MkZRaVClxUL7BmcaQ57ncFt/c8yB8623cwxKM89TMslf6xZON
PzQnWS79KGbWvyd2fRJYeV2MvsGKkYVMeq7wAm0tCSSkIrzB+yaF6/m/Bq18EWSscvlpOtdIwxdI
UBpqCS15A6S9btKrA7yLHuqBTC3C+lIU352WNSnN0xN6a/9+NHdtv1Kcxj94uVVPT3dhHminr6Br
ghu6PcIE5K6ng7Jb3Cq3joYqUhYH8NWuDv6xJUbpBDGjvDYtp/vRlTLATTx9XlP4hloypMh5lFUb
V90ZkRBPXwGSDzGRSG0U1jz/mC0NmOuwMBPso4kjdVi40hqR6uvZkb511bkkOMQVozQ/iF8hb4th
mef+M4x9HyEshxgKW2oDX6o4dgEtricFQ9ATpX5f5LJhhOPcAc9H3Cvd5Qtn/BunHZgYbU+EfMAG
e+jqGWJ2aSDHLqF0ULzQ7DYJsswDFNGV4+37vgN2oXj2meiwWA8TSfNcoT7VnJ6zp29r3lf6Qi5w
jUaJzjamoXYFZVFa1DXZ6yApkao858E/JiaJy6FBYf9sbtT+moNtPbfUQCXeI69NLJA5m6EzizXs
BhBJCmy7dC6QEXC/qUoEyHsjedkkVshwqhvyaCSwXnjXPxmMvgMXpxZhYXF3V2/JuIQScsFzcNuB
i+JzXQufxPAYno8DgpzFESs6a8pS+wnoNyrgL/Kqgrj5r1JEvdWxNFG+rV4eBn5XWQsjAaeG+sxP
puAPDzC9/dh9OFdOdsvP2c4u9P6I4djwyIHuwlWUdtOrfY5Oi1AgZPuc3/VP0Zgx+XOqmhsKHx9p
Kv+o2+/jHA2mNB7sJbWyjzJXXqlex6Qosonb5OUtlOj+HmvTkG6QgbACZe+I/LK5PHVn8KsgXl6t
bORCSkaNv1ZQHtybbm1Qo2PVghdI4Bra3iOWLZWerZyXqr0f4VMLH6cyFNgi0RsMfFqP9KwEEuDB
4qWIDEoOml3FhK1D19ga+HIsIERxM5I2xqJbUgR1jbU77AdO1JmMzAp7ApwaEYFEJ7dI5bgxoRbW
IGb9IIerxXaMknBKawneuMg4HX9nIGSOhwXiGs0VDDVN/1gWPJNiYhx6RG8GOUAWJAhflYtC4HVS
MZM0nfV+ZOR30MGHyK9lmlqEa3aRxFUV4jHWJ5VGLIcNAofl9+NNI0lnO2u2Fr9yiFn6RtJNn1MD
CI9tFppyLRABO0muj4qeirzlb120lAenPNOZLYePdTWnWee775ZufQqad5dIwwI5anJ9yW5fa13t
XjSHjaTkl6ig9q/MqUz5LF4yG9+9Vz6qlC38TG+dzQPAT3wHk4FsxEvxEBBWpxiajDf5M9s4EJ9Q
vQyH069ZdN9VTAGJq4HrHrmDf7x+iKvXD8CKgwaYUbTS2OjFkGeLJtl8uYTWfLWa5E/4h+MCA6kb
rgGgJNcPa8un7WLF7Dnglj6mu5PcK6Y8QqYrdf2ANAPxsyGa2btIzTohXh/N2oPBMGhg4UxCMO96
kMfWi1KmUAtjM54T5Pt7qg/KGTjlU/bu4IDILrtg2H5eCCus5KREMx584HCuTuF6fL3SXaLHzT2i
3cIu3+Irgpz9L71tTXHxJJ31BXr2kVdu25YZFK8VGYrGJ4OcDCwgfcJcgCgqrqxtS2UvolgkS8cU
w79ZoLyEyD1funW9zVDvfBDCmOncooRstm6+Mn1Wlij7vrGm+I9lkLCOyjNLkGPOY8sYkqJog/xk
XWzo/9skfGXGB48MluYHrubuZ3c92TqXqw/BZbJ8LwdgCfc6LOfrz4L36PuxhCRGIWgCF/Na2eUm
0qU0gGS4rGDPAMnLSJaHG51CFagsPPDhuHfreGQ5qsG0jc0FXE9UeX7gUh8MnMM16aHy9wdBvf9M
qYptE2Vt7bq7feQbg8LLH6ZOJWYXcdtLgLzgYcNX5S6zmMjd+QLomlzP6lx/2kSdE2Z6Uz5JMxmL
urxJGUC1UKpHQIeFxGYEZNrwEgQjLDP6Gzfpo1AJLiGyVh8k/TSJVhGEMf/vax0oOKl13wtts6bu
lgIkivnyZnyQ+6W2yrZ1PUcxHEWhQ4om107YkIjf7brmqMGCM6nJfQMflrTlx+JKvDQa2yVOfeNI
5Uuia8EdcAVsyjt6xa0IC6khpe8WMOdyrnbi6HPGlFOX1TlbzppI+MbAginglOe80pJDFxst3+bS
/q5V/y6Nex1JUDpV0qaZHfEZ1N4KQZ68O9++EwAp6NnpOIFy6K01saLM2ljXBmElctRHZhwhm/Fu
eabH5e8rT04jzLf22Q287gN+eHZSPsSTNKtLL6wwojNYX/OMUORFiX1azBbJ2601Fuif4Dq24axl
ghbArl083P+2SUfyA2ezpB9LAhmAlI9K1t6Go3Th1KEPS+XhkO8y/7IG45RXwXiWgR9LlNv9idTe
KOzZKQECsIbk8hwFL3QbwAcCKne71EQOOvaBedtuYTWzHMNaGzaRNlnhTShmyZ1RQ16vcpj8IgOI
kVCSd/7GwqgYjbNZHQ6xVWwW8JEJUpKkUH56BXXBXF7WGN6IzGS1H0cBoDvso6XidWNvY3wuR7jy
48jNNvl4mvlKOcolgopvdD1wLGMUxh22Nzc6apZR0yTnywU9zy2wfCh0Q1i2Oj1ehGiXnB+6X3le
1Iy7ynY9PMgkLe/ED35tgWl+NyrEVBobs6e0LAj5udIzI5kbriPcHjshvsDAiHb1WXascfeAOfNz
JivvkLsgK0DnkqzHSYiboA5nnRZOD5cswlapr+Ip5ZwsF9redcJNrVWgFG4SlMeOl1QMl4PaFIGf
6WV1grEXhHjQHwRFMtUEoxfg85ZEEwW3QHbxNIpH2E/ZV4Bcl0ctB0hnORMi5WZoyhojoDehNeR6
9vtzz6R+VOXpMkU24Yizxroj9YvlnIAfacYo5lcTMSbNSkMZXOuVAZMC3K/1Ew0cP9cafp4Wr8Zh
ZtaSF7lYFjwDEq3qWMPST8Yyym6YSgDd1GLuDECPGMbWLS/9l8GyvazlkLPIetKO6JuULRNeLh4A
3ekbJsYgnAaw1pgacPHdcajceu64ZCbWniZ6/fvX00BSCAGAdshlCCF1VgcScAXhfQk/a3R+E/1F
dcfpKCT72CdjsuFWgbIbLXoYm/98m5DSwYwgeM71xJAyKcjiva445B3V4lLjJ2u+HhHdBLXd/51t
20WYyARBoNiPAt6SNKVHCnbFFgvscEk10n4S2lMwLarwLAT9sPWxMpUTgyzWBxFfmOM41T91zN1+
fdyNgSAcGtKYnblql/2cnKM90fiP45D6WHgFDcUYoJWeXFTXTig+B62I1gDXNX694lqP7eeH9fzt
UpFLR4KfKMy7xx2RIZbdNK6x6x3AppOGBi6MnpuVIpM/CPO2qPMKFDMIUTu5gSWrSAC98rJiauSc
GQQqq9YRpEBeN0r42zblK2+1XyiwWiyYtbU7QjaUYtBgKLlKZ58hvYfRP4Oa6Anv1fLk8HLij94m
XKhKozA9h3ZOkl9hlC/2p17+mJHieacWI8XQF85qt5mKSD2mBVedzkh6m4imiH34YBPgLE1yO7rf
cOBpsQi5oHgKSpm1uj+2u8TzYQ54FDm5KYKDGm89GB091UnViWQQA/ZQovwOLsoDR3FBEXpMkjw4
opk3Nh+WkvCekq9SBxT+Pl++L3pCfM63wVMPumKpBbrgPOBpqpLAnGFz+iysoPOAmptDd+EqYpRp
3x+C9ZbAU090S7ujhrOvbgfQri9mMZrtY9eQjcYVhpsWX5NzEXLhcEXkTntpWe4U1eMY+tkW/SrY
b3xMLEXSfabsbDuasnRP5ljCKJVwM9EImIT9rDGHfwJEAomQW6da3YEtKY7NiP+Y0o4R2h0ywoF0
gaH8Uko41D0DjPc5l+jtT+dqluXosIABRInYNySeZCHVS46Vs6E4bmhK3vnkndujGqqztui2z17+
JWEi1gFcLmhf3lEa5l7521ZQWsJltFWJrRKUJy0JiJb+HIIf8SJjyHmVZuNmzwztR+3RWL5C9KvH
w2ITe+dl/MoxKXmKZxSSixM2y6qXMdN6piwK51NPLA4jNZv/H0i+pAMlBfU1aSEyfVHyseGqEiRx
WT6wydvGtZF6NM+Ei+Ed8jCs3Dl9Nhy/Kp1AGyYvVw6Gv29zoSM+klKWKGvkb9/hzYlOjM/Uw1o2
EPF1GWjlLRJGwPTSrp+RYOAYoD/bVptM21+ULI9xWyS8ouB1CmgFME/TsWc4HhMeAmGpa2UY7eaR
/pjtv7V2gt8fMp4+5Bo4uluJmbFPkrpHE35TMMs4WERtdQst016xXgyqE3N/1mIVHNa8BjbdeD8X
bwR07JuVL48vNxiqULaIud0/Iw3ukTPx2SdQoGnYMlvcOFIIQrm6529MShDdM3AVXtxxZhqs6z16
fz2QPSPgxmwLawgbwiuUW9U6SseBajeLghz+mQ/8JULdgBLhlLTT6/DvQfy4WeN5paomH9t6QCbp
Hbd9Uuu0bBxrr8UMLPIzk+LGyAqUf+q9eAhTrU7/MeVgKWJubPBrSMbknyFCu6fI74drN0ktfDfo
BGo042PLKzoPAdE/Smmw84uzHh/Gbh+tp6x8Z16Q1/sP/RTNAWSbQQQ/o6avO+JLaZDEboapNhcy
pRhKVDgLVJ+cslA2d7DJpl0kvr63XEznM2Tl3o5PdjDYJOYkEDM8jpfQEuDg/VfUlvvTFJdCW2U8
ILFlTs7wDkj+D1tMWfGZr/yCNYgLBFOE2GNjcQsXtxS2AluETGan1tHJz0kgy8poUd1LryONkX09
J4oqrL0sQexbBnsGjb9TzeO0iCrvdDJd5MgF8qXyhjPAMQlbn3dT3GVJZt0RgnnSuKU4ua1/6Ims
mDdlD2EBrdVOKrcSVygpbEqba3VONfm1wDmNojKp2BR285jdWgOSOjV1iNNcSIy9gAZve/lVutwv
TZ0P66bXq9vgaftV+L2fr5/Bwnt6LM59sqkemiKcKFZLb0ctn3zjMMm+hFA+pbLj6/auDv9J6a/2
ufOJgQlNhGYqNWuFxxJmmSSAp1r5B9K9Z3N7W28tKh+uwFm/2AnIp1v3RCc8JVDVPL3JCPgY8UM2
2jpJHpDHUl/19JDfe/kgRrT5KjBoNnug76dtZVOMDlsfvIVZMM+nCjWVahoZGmCyBtI+f1mpqYce
u/TKIo3qRi6iE9EqXoI5rdWmQd80t5J74Gsknr6FMj+mDRR6UO+IeNfsZl7DAo7D80vrhJ3nO9MY
tvhRDS335qCzGI+35olTJ9k49F+Zsn4Llm/DokmM6AM9kwNgW3waqkUoSWQVhOWk7eHP+7rFviK5
kAGC1iHEG/9gCgMjXXv635ykKJQ89unlOrev8LmnY7gfWe6DfiChtWxNkexMqfI/e/T1FHNRrzxi
loGrh8CzWu+AFEVChrtIYGnOyVGbXaR21DjSHy7LE3udABTmnoUm6OUqfdR9U14ei3tD2mKcRG04
VUlltILmz4V2a7TdzafHT9IwB1Dz4g+vdj09HpjMkXTO85YFwWCN2ucfBvDK6D6fdEif1Sdy1MMh
8CVS/54E3BWlxcYGAvn50W5RF4L8a5tihwrhT8KfL6pdoTKvwQtlZ0uYnUP4J1qx8PqsMtQWHQdN
TEsPaUKfffn5Xok444iP6yVDbjuyGAXlsMOAPDN1aV4PKX8rkKiwXvYSSBzKPH9lY23HEOXhYdMh
iLu/hqvDsYj9Tb7vfl3oQvtC4elOEc1TmMTVczXMkdPbm0Vv9KFsPVbdtt77jG0KaGkeSNfN+Hfc
PYcoOgj2Wtg4BDIqY9FHYb2NSm7gYCDO6esM+15PtOY/wV2kh6RzVK9gN+1E2wIWuqDvjC6Ds7ly
78g78/uarNF1Ho7tgu2P5jCZFFz16wgBzYJWFS4DRSANnUJKK1cZwR2fLNxtwyUsz2pUt3DLeCxX
9ly6EXUTW9IafImBftugmlcuERwV93dsXWYPURuZVaOc8tJJSrqPkBomsoh5MIs18jY6UiyDZvhP
RjHnCAvth26Uf/XycHoD9Gsww4vuwD97jhEL/vtLiYHyK/ohDOwKVI0QA3X0j1RgcrskyNH5yXxY
b8xyQDFFDoS8w5PPgK6can6+FynRIkv56HfvlaVAVdghTX3WoIzP+PY9LmZGvAN/AYEFjwcGSaIW
Jcq7SqFttD1qSqH9ZV6ZFUePM+ncSMzsQqVVnYHDCe419xB1SR4mBMwGJaiAZaOxK/aXNPY9p7zB
jH/uvpK/h5VKVy2t8x6pG4Ilaq/ZJcI2JMWBQQHEe7xfWt3GnB/GpYusUAjpCBG0DVQrIwuA9kFk
1WVUMi6Ld7jHpCxkB9ZaalJrulMERNTXanHxgrhWE/rpFCdeCJKy081RnAftEgN89xZp+6R91Mmq
COkTCf1Ol/y1RFl4sFORi4RrFOf4YFN/H3ZzgSBdHcTwzGtLDjNLAXm40TnYp4uZVk9C74uO9e/4
477WVLlyuJwnxgkFPqsk6pQbgaR/wDSsitFqpswGmp4T9GFT0EUVVfdPCRrPeS+CIEycHVpBFUNm
MJurVMK+dlbYtlWsujZhk3M2tCr9O5CSihXTCZgdx2S8N0AuDayGF+cCFxEQWM+kfyi4m3eWZZ8v
Z5wIQsQ0kUkxDHaNnY/Yf1WqhOKxctobeQO7UzdD43hU3bThDxCw6qO6xxpHzsNgTzdvW5sDZ47R
wcQIAfO53iYiQ2cAii1Kl7ZH8PPGhZt7+dGxTK5K4MmHWKTfQseCcYbBeNxYKrCn8CDDxFY+MYqR
RMdzsmV618PWaYhH7/BP02ZlsMxbUTIJyvSbDjrjNFcTHEbCCcebbZBav25JU0pGZgaiNz6x0uTr
72Jhc11iTPUHpE4j6csZoDQGRrOy5sQy4ZDL3u08FgvQ2IYihCdeS13Cuo0DOux6cSkHYeHRdalo
kVhC52Wu4HQ1vBuWGbK2F88+QxyG4UGHW80nzY8p1R/Yw/7g+07dl07oCi7D+WAQdUgtb7fKhnxs
nXhK5gDD3MJ6iQY6gJvMJMNmRKhEUnn0XlQwatbRpFLY+0SmwoDEcL3okWwxvo52aYDKA6FGVI0N
I7BUdqqb2O+TsUijeVs50glm5N2KKo+9x65fWVtXg0V2P42zs7a3P/M0FkR3i87gc5C3YLLeHiJ+
MwPQ7cFuI1UqVuE897cnsrn+J3zbvQWKIwdjWo4MmZrcGvEvKgQJl9GBI+9SBEXlRwdw1j8wOT2v
lbw+UbPVnqoiDiUZDDjy2MFRaBwYhIBJKxKBJ6fMsh9UohW8RqsEFMbhEWreX8PzkV/r42EnZic5
6zzxpS6+iW1DRfvqTG7aPDpCZNC0nXDmNk9LbMTGjl53I+dqj1IH38OKIyEOxvBg5zac0zVPED7d
88oRK3nsas9ZtpPf03IGam44IVEBae4QPGY25CHsEqtHqnhbdNXDY2pIMPVl0FcslNg2MAcdJyD4
3nWTTMlcnIAnYISq9BhwdACVnR10sZnpWqMunj/6LJCdE4TCnDulPcZaejDBfJ0yNPljW5aq1jUO
EMF1oqePZ+4FHyxnplYkR1hJbah66/usr5x5K0kZlpwe25PQP77gVF77qanH0Akw+o7RFIh04yq7
ZxefvZdNLZ88hI+ojpqqppIWYV4Xem/uLA7dGCP4BynD0Gno7fGlwv+pW+w9LwrC1A3AIQLNC4y1
UIYQvcdToTu+bZP4Hdaa9jk9JopWDKmsZXJwAluNGNxYSZuoJYpTl+/2RvCnOD1kri6q9sGaHQx/
ekM1FNhgk8BRqUTUsYzCfHEbR5yZYDCmC8G1kNQ85JSEjnL++6ysEF9DgJDcyL+GMeaS+hyIqZJD
O5nktWUMknwWUJ7TdUAF7CpNkfk/6sTilUgCHTX8UTks8Im03pYFmSJKyHPSXLNspkzZ1WIQB6ec
sDesWE+xFzz6XNhfPqvLyxnK7uWa1z9uRVOfPzKUVoj8zwxikPeuWCoTE9dMFq7ypMl+ssl2OXDg
RruIcHQxCPwy4BoMjwei2FCu6/JUR5LDJaGmqj2kBi3tZypYcrpX2kLS4RyQ8vyo8c6JiBIB+4G1
9JPZLn1uePgq1XrHssls9KWaMFkJzvB/lIrEwEhnMvfGLxfnfQmvXDHhWQO+kyxOROzfqjeU4/Eo
TpyfkJuWE6cpkXd3eHTHinbCItPaBPtrLy0qYV/n4FnT4lnajbaI0rp6kL5/NsbF0/90IghauAW0
XlidKOReG9BUTESggyt4WbEG+VQE9OhANklctg5fmUl0VAH2PQ6eGLwBNB8GAs9mqH5D86L00mDX
KN38AK0FQapuBeCyPz7F/ngjIVer1BYPuMIh9HRKicG8LhqSK0fb48YTnJm6uU5RSq2y+FmhRa12
e7lU3BEJIiP5Hs3Y0v2x8MhJ4EobS+7JWvK3Pct+6YGCskrQvfnW89eWZP66h0JwD5jGDXXGmPzO
gFPJ8ScUOP0n42DX4i47/KipeAZa4Thb6nchHDGOdm9c4jBb9i2PwApd5A5bM/sbztAAEnj6cGwV
gr0nJTMUcMQybJVMVh7fW2Ij9N3xiGSXnKKFjx21yOUnlWU8EMBRuqT1oOXlpzR0WVcbclBYzQrW
ssmQGOoDBb450ngzoS70kgF1NUhuWZuPgXcYihigSNi1b3K96UFaj3vQ8YIuj0XJDfXY19cLi56Z
WoAiYVruzPbZkoJMz3ZiCFfaquATU6eUAuLjLH/xIOuSYcsEgE1aIx788U1Bbiak0mKhQTkB9wn7
YA4C4O837qqqirbRbKeDq5SjguwUX//Gdj6cGbKpQUiUteJ7speWQMNbYXUncxFMElQdeOlSVLaa
3ugcRAbA50kHYqhlvlWyeimQznoBQuJKJ3tRVp9w2ht6wiyseF0rlDYaS1d5K+zb8OIav0vl1Vz1
oqJRbRn9JoiMvvwaITcOZotIAAPDVbz9lseNt+IR9bn+jKFyP+vj21EUzhwKX1w3Cdl84fu8176S
y6ulxgr9blxv++c+ICOc/sh1/N+/W5WjyTKlRkqTYxcx7DsvfA3dqRYweGyXx7LNJzA492zynpeP
AzDOOovMuPS1fqty6e31DhQqWBH9PP7jXsYN0NbdSNN9pBAPI9/puGKeH8+hS7eSxZ8H/RejM/dY
VlbZBGDSe0G5giejCMvtUzqaaess7t1lQSy5NMT5iDzuS3yvCctxLwTFXujZDSc2qEcFfx+Lg6Nz
R2aica8o62hZ/7RyeSi5IbtpaKv9NZlkQCx4q3zALo5XYVjGBjLanYbomADLWFi5VWYgBpAFJQZN
JXVpILGJFj3r/7zPt8C8yK++q3h4wy9tE0QuwsR62UbztotTQUgl2WwmomS/QJU6VmmhBxnf3mDh
JXK5q6LHiYxNf65dwGFlW0j4s55lw1SX0WYiV+J8qOzlaFI+Xk1M/ttTboOFN7GyRQx5KbYCelPP
5x7FZ4qxDBCXzrQhu0GwlZLSEjdR25b/xqOEDZhOaetSZtGPqNyT3E1igzl1SSqxPV0i+MG5qSIH
MAlp1DThKjSwY03wHhMj5FOwNjc/oEEGbTC4/ozW3s04vq+mSzYB63GBNYJynhsTYdZZmbmxim/i
m3J7IW+iCP1AyVFXuJ/+W/UvOoB9BTHuaQZddJ/YNG2g/q3q/JoYRA1ZfTphZWAw2LqQymnYMZ2w
8lLF3FbuMIGrfqQzfc1gzn4WkW9QLaKO/JpjgV07dGvGF2FVPzKV3+hK7ybYfkoDJx9mKYxiImKA
Mc6ps0kmAh9RRw3w5aj4GZEXsOByuTjNe0ZExebN61FMt2BBTDiFSLwt3oYXUPS3a0SgmNPtuyeq
O3xOCNVdtbMqfOzBVRFyY2lzgpbd/6LM8CGApjxn56ZCAZ/8YAtPtXcNUab6Sidmd0LczRioaM57
UxMcULbde9RrwQgjPVb6ySK6UqyLtDMwIGZ8ucooJWg6Rtq25+cAQy5gNGN8rv9b6zvWuobgUC9h
HDC1PRqOcuS6f372+uaA9rBtVfld0iZs4Ku/sn1oLwRWlk8eGW31Etfth1Mm4p9ZkDGt7IV64xMb
+CqT9VhFvekoVHGSMNsFz4hiKQ+5FXEgzHcT7f7kVQhqResXpxyLvbGRAyDOdXl1Qn/HFgDD1REY
+WwfXseqJ6vQxah8/ySgJEVw78eq5+fZntXWZ32uW8QHeYWb5YoO1kMzmuNK8BtRHtyXC/I0tJF/
QEKCOyktLXfe4/yGpTNoGkDM2WdGuwIjZTrYB72qH3M0WONpkpk1nWx2SpyZvgxf6HPwDtRaJc+U
Aik8P4m84gt8RoVdc2y1NtHBi8Owkhhm/Ehvx/cboUeq6PiykA+S70WxPVkqt0wNgITOr/Z2yeby
V84xY4DkL/0iJcCtQp86D5UnLraSzFdaDAIY9xEfinEXL1tcyeT21RoGLWaQDBfFnS2j1DzqP7ez
TLjDQFwKSWlYZqHpa8qLMT1vqt3Bkd7EPUP5JO/TxjDvgcmiL9SZR6ymmJ1jcOs5H1oLWsG+pnAJ
A60Y5XcnQUn4CkGoUZzTVmn2/yk/q/T7M6DFTCHYKvDBw5GnP5LxOJfXyoMjdNUtd+USR44nXLP/
sZX/rDi7X2lsWfPhQ+SI6oHXj+jIQEfC39DOZt8AjD+FIZVy8oLx9TxAoH3l5spSktiHA/K9GCwY
VXBlIGk4HIj8GTQWITcOLujapmTWU0vwcKEDesrcjlVJ9J2xhrIbgZ209TbGsPUcD2cz4KHbJL/T
l8Mx14kyA7hKlwjy0lzqI0jOV7U02Tuc9IQJ71PVMQLWZBchygGqo0BKASXMxlXGXC9TyqYXJP62
K2+4zNxzEB9p6x7wo/2D61v7OFC+F45bbqVfQS8w2Cz/YOPzBxtgRRbPuxwk/PpuPLPtUwdwBabz
WGX4CZRbGdlRviGxa8sdLzRkSQCOTFIVgK5IvckTpFeKMptQbXpK7kUum7senn+tgu4f8B5WCdpY
h9D4cZ+gHgsHQP4vgNOIQGq4SIVKmvjOAC6sNT/5zVpbBWjm+JvSqWUtmFFEAvDxGr4VR4wmi0n6
nxKpUckjRzpXLEa+ApO+e1BND94rpcplfFYMBL9PPscLtppnF8/Fu8cnxOsCRi+3e9+qDA1zAGH4
ryVWhfmJ3TaJ+Z5mwQGjfZOp+c1V7BnZ4/t/2NAvMS+cRo4v+pBBxsoOsDKF/lDdJijAAxsrn3KD
ztHt/Or3IYjrCQQBgRC64nW31cTbMs1pBIoPJi+oCUcAel2Q8K9k3Nh7Ubjulb9yiBOC0QwNFKzI
+Ki3ymtBQAiH2hcMQQ9rR3ukHgxnXrJyouudxbbQL6bTHmha2y6WeODCAWPegy8JFRyfCI5xPRb4
pMHSWBg/C2AZPLOQuC+xtgBir5HOZNbs5mwWOvOa686RUFfYgOfiaSqWIpSnLISRFURYowRPgg3i
yE4IbCGrVj98pqoG/NLIfINIVTTF62jb7J1N2a2snCZBXbgmj7ApilSGBqVeSvOsKHsLmolW3C0g
LZeYMoLWUlo3/8bvvg+p6aDhbnWrGRvts8hTyRyomeIujxzvs29FeAv0f4sdxRiggwBh+E9sABKX
a49M+ICJ5BjzsWWz58d2I9O/1Rqtx74483WdYg1HceeUBaKemTYPacMqObF0+uNTADPvoTxLbnQK
qX9qvr0pjcs/869bHLaH/mBSIFarEk3AYWLZN44brXAtNrCo6MGyB8NGwUzwSfRrtkTKP15P4xPL
P34gu0Lajp7M1MVF1a8LCJIF/au6A/FCwZfTR5aTH+PLVTk6+qVpeyrrnp0RW9joBeICD6jRBFoh
wORC3Gby++1q2ecygoqNSsynEKqWG1PzzQ50Ic9+AFvHMITehWBZ57+TyzIMDRUDiBUKofQZn3xP
IkONzRZvigjKRK7h4819Ss+4D1HNDjzZDofZSncXLKiSyi9fqKWs2spBW0QC5gxubNc6GdOqs+xE
69m8Ap+24y9Omqyl+V4kUYZ9zovU12zA7V+Cjfn/LICNcC9xjLaoIR6tB7zH+eOlVv6ow8v23YXv
8HoYPMFen+gZhSd5hdmRs/aUqHXw38N26Ozfr/a8el2CtcWYzfZc/Sfd0EMYe+t1KjyOqPAUMmws
USqTa3GccWqSr0/WlyBtk0fWkcnN41R4YUwusRreZIB+n8NZkHxRqAbxfZ4qgytm99BIhG4x6IjK
AbMScjCiilhttoJ6U/NqZ3z7iEbBRwobd1iEWiBamfVgXWOG9XqU8LqL2TRlOVX5zaIXXtehPbpJ
737mwggfIh6pxxFr+bZJ3bbFbYWxzTFtOInYuYTEa3qb9jwUdkUWNkfuP1JZQVHrW9LNBbgLdO8t
9hS5+NFA9BVT57MEO84F0Sa/dPNaKLaUuiThA57HgZHYW1NV2K4csh6oVtG0AflSZ1OhB9yy80I0
9E5s3twLBj3abeMoNb/tQ5TC9G+Q1MPD5LQmt4sAv8ZzhwVqAd1xafb/u2wUZcqgNEzNhizXanvC
pkvVZmbxFeL+sowQnbphW1jpPG1OXrikaRWCT/8PTxog+0hZagte0KHPKf7Hnqn7vk7gjXNEcQMb
PEMRCc2fUPWiTprXNr2PGxk4xqks+YJhQq5nRviz/5Tt8pONUpURj8fUAvdhBHvH35lMNgL8lbzN
Tlb2azHi+XOCkTwjQ7S0OA0FBhUQMEd4yPi/MdgxWoIES3BwCOtyWdPd3OQbJHzlP2wc0WRTZd9g
HDsgxaU+fftxjpABpg7yvaosOAgbRFn+IQZyx2w+VZi3wZvF4N6G57VbRe8mItLwmXjp92B0TZTJ
1WGdYkHD5AzWV+EhklfEmKJU+mcRiyRgQKLjYuFaKS4qWZoShkd4IVtepaHGGj9QgkdpXKu551mL
XjiVdNCQBE/L+0t3YcM2rhBEamgvY3TaFPogclm4TmZLaQ/8TwDSHIA7AsVqSmiLIYGKRJlxSrHW
Kxca0LSPT51uEHByd3MBkIXZxmMw5hmtpu7SXdQv7dG4G3tI/1AygnJNW8dmJtVklmReCa+Ch8NU
9r7UYbq433msBQ74q0gbIkpIZruiuSTNGQ/LmciOX4Ow5zy7PTrBBypXLbZD5IDp7h3iN3oSWS+R
E0l8XoNH3O87NjZj97TEoJrOorlvHhg8BJqzyukqxB2qy+8O0y8VoUmBZw6Tm12wlN9WFjNfYv8Z
DkBRaeyKBLglpAD3/CnG9S7eUcPy5po4YLJ6Vzz0hQMYew46P0QqTP3+hFsZ0J0OZa3zV1CRsBCU
rvowwoFjquZ6G8yvYMwE1TYtdFmEvvPp/2GaeJ88cB+PRVZScEv5cYdPPKuxKwPBATZAQpXQl+kM
9sV8muZHqKrDCDu0U67hedkzTDjf4ROHAHCYZ9KRJiDUZx5Kr/IXG0YP2dzYrxkXHE2ZCoQ6tQM/
hsz8Gfgt7M+yHvlfZoVEFtNlIQDWjV3q91+5jKNl4U5AWJg/9p2ABQqHr1uu+bUMjz11LQHko+7X
0DcQEsxhm3uBGNCAXYqUvSqxHce9PVwH/4jlxe9IUsH0M3LppXg4y3fw56SFt+2qeiAEVaQWTnCU
l/DqFhvhOW/XgogrGaMXtQI3/AldLxKDKt9vJFGJaDuYrZynWiwDvnnwHFM28AL57fbfY6MfP8aU
b4JOEf8r0xunszmgp2yQE4FCJM2Rf/qqrvIeyaorFcXR0jHnWUIYKH2TVSKiLSB1wk/iJRl6d6jw
c0/PG7/dZZGBGZsVq18/lZD6pfHkUWQtncZonXvjW/4IJ3imS465GzOpb2DlByYcXwRt1J9DjHXk
qE6NVtbYl9/hSLR3sdsO6nK2EEVuu0eH1anUOlngsMCxJvs64C2Vsr5tIuJs2PkUkqFjnitPUrR3
aeLOtAu0cQNkfMhWy7hjwYZ1ImLgo3wG9SWFn8yv74nWm/oQFQW74qHyjdlPbcuEx+0tOmx/KnKG
F+Jr0flx3rlYpozEIJBAq/x/HFJb6CvMR2ppSgyWrpe05UQp+AUFWmReZn+vz0xWRDYdshXVBXOx
K7iD3RVpqs1HaAnYoM6fyxYH8LvNhoVum5k4mp+atD/4K9wSlLulSWu1wec+4RzU5mE5QpfbZ0qe
OjcYB3wqJmh68kY2SxJ6gR3XMTY2ztFDXQoRYCzfkS09lMcshbp1DrIOaadgL4yzo3nWbx3XT4Up
i98ai7ZBEDV1d6vqUCwcO9Q3GK/A/sBa4fqQZPRXjHkO+8chwdV9+jpr/1I6lqN3nRA28CKXZmSg
mXhINpAf3mRSBU+oEqNHAoo5hbpZni1KRfCG8w4MtN5diyIZOQwTmbA5WYJNA7DxQxBSsCPfto8f
eNa2cvnmIRSkMwkTPJrOxv4Sg/yGXHpZKgPutLDaycPvITCkGy0wuv0EKOchamrJvJKYk3zGTMPI
XofFw4TtIPho5aoYIbqHIq0DGGKuZRK3krTwKqGVtsnCEerhGZHSJ+LUlzF//SyQviqiCZnC/O9C
cA74A4+RH8EwaPJ5HwOMhbagQApbnhWEJjd+sBbrSAIsdOrTsS8wL/yT99sD1MxO6wbOe6Ht5JWO
GZkwSYqiU2Z3o6HLb0RNiy7s3nhgIuDblGQWVXwo4607k5ktc50QL+WgYWJoDa3jX/l2EARXwzMJ
yYaxS0OEFRUWnirWtHiezCebDZ96BlMRk1OGWR9kn2sUjAQOQft0tAge6aq95F5wqnUgRsLGzkO1
8nvLOLP6DsimfcrlpSWwxX6jPQbcb0w3jN1BQ36pzLLQCImh+j0fuJpipr9Koq1bVBfCtczXd4vl
u9hPwW6ejSUvKlqf3L/d0UyevT6vbFA0yPghgtcXvo3xvCk0WPEG9MJvQzDQnDOTIke2XHwgioYX
Qt9DY7desyEDj7UhQoDPURCQ9U58nDhlg3cbPKd5FrCtsST0Tu302xNsMzRuK1Mlk4InuEySEHJu
BSZ4uSl5hPITsNAcjLSMGbE3lJDpPTt+xx7ZUHf1VDGSnIzN799vzGIrck0uhdqiWMy9A9bw4VkY
zO5a+wyQG3VU0mGZ8Yg/8XAeC2kydLnbxriKcBqFulfiplL8zHsWSENGSHfTMN987GLwvOnp326e
+8SexKUoF7QT4Xk1KekDqFboUUB/y7/0sUEIUX5znthMnTQKmZNF3Zs2iLz66V4OWyBroizfuFVM
O48g2bdN6z8UuLlWPpR1+8i8Xgq1CuOWcZuiuoPsFdswQ+2kpNJxZfcgeDR2Zme2MKSns9rcXqEU
OEU0sQUo79Pyl5pVprx1FJX6YH2hDB1w46YvuywgbNcjTCJUqtxw+Zsgh1JO5lB9W1Ls44kpmMaM
GTIsdjSojJ/jKD+EzL6raDLcixYx0yhtbI8jPEMk0E/DrRyMl4FHE2HXflllXI8wnOJU8826QgXZ
7XYVYHZpFl/t+5NV+2gs/lM7QdkEuWC1J8owdjZtRjVnCTmCXQkrzPiFLL4+nDXuHyNo0nuKZ9T1
7IioQfOHAuZU4Ez6Cy9yiVzSkjnXLQHhPFqD6eNzK3dMcBcXeEk31Le0I3m0+E9ok7AiTMvSCrw5
RHJt0h5YGClBOmO75QLZdcUcZosoxe+eYfurxVOwjRh7IUs5GnBR0jZ4k9i08+gxNrJNYB3F73al
sHKjoU6q3HmgbZ/QvVUnvDrUEOQGvRWkVkVqN5oB40XotqdlEStIGErPufRXTaoHnHYblW1vMdRO
ccN5p0x6pY8vXKQwQ4OuFi/8jSDGbBXo0OPSZRqAAJozL2GAxuUed9It5yV7puA/od2YT/BVDTTi
g4D8wLV92V1m6BD3NwNngq/Bv1eGWHePMmjOJOnIAJICqzh3+4QTJnSe2UKzOoYkCg05YILSH4ln
LBe/g4Sbj0lYwFA0fjoau9kFGbA5ECPPHmEstIBI1ZU3mJ6+97ZUDBKty2tVuCMYCcfKQCs4gZFU
EBTl88+32bqVJCRW+xDkkUshPvyZ2eE3jKVGCQshrL8lhdt2rPdcjMMUUnXsrGuplad9gLBVUXIf
oUdEP0yj5Er0esbBSBMXAnxmZI6vns91ziO79RdixXpr7lSiSN7lU7oTkOPAkEM6E4FqPO0T0BWJ
aaEIhN9QDfkM8Cw4fyN0EQhSAc3v86KSxhigQDwjzAnN/o3vcE6hjtGjFxQ9kouwSpwwHuHxOxsq
+CkINw/eC7cEOcQRRo5Mu73+G2qWFmBuZw35K9OL24eL0KXoRKRDJkiRAeJRDyRSOplqAVLcGspv
ZpAX+Y+mU8ovEaUZRJr4fo8Caqb2UI5sbngi4EjSUBHXOJKG9q7zGKWyXRN1l9141gf2sNI7k8nd
gW6JuOhzvnrkiYKHI2nCzH0ERCOi8cLjwsyVs4whnCNr4vCTanU/8Hp6cubkt9GI0ljUaI3hXcLr
RdYh4pW0yfP8FcaiFkjMjRl09G06ZnkBlzHBVcEr2PFGAtgI9yzZUagGew4pWUl6OZLpHUiUQCYn
TG1YPqfb+5vL7r4tsBRKN8o7oilJsNjxZ1HYF5xyokQVzceLrebkVYQxNrujnjpLToPS/j7hsBkQ
uje6YRZcQ6PlDzjUPKJg1nTwxgdXcN9f5vSPsXD7/o1t0aMzRD4iz7fMqoyJPXSzMHQ2on0=
`protect end_protected
