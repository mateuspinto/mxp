XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���'m��̨@�S.����� 	P���ә5���'j��G5�v>��j
鰿�
C��2��h&����L+�}�90>�aC�����nA���bomѤ���Uu�&�M��NfKz�m �J��yf��=��B�)��@C�֜�Վ�)@N����U��"@E��Vb�ga���'9%�v�_��w	mTWi��$iĊi#to��C��Y�n�.E���hK�� ��w�U�zj�ܦՌ��� �Q��7��~�I�Xe���M�p�e�ZD�!��o��a�D��ĕF/,P$U2���ow���\�5 �ZU^I�-�d����Zf��}c}�ܲ�P�I,$sﯸ���d����Ħ���y��?���k�M�F�J��֤���x�Yx����x4a�JҪ���]W�N��#�_�6�Y�:���J0ǎ?<���/�Va���+�)��q��s�E�3�����O�4�'�F*².�����G�;���o����ΈbP,T�D.[|ſ1��#�V�Պ���6;���Q�gJf��zG!Tgֺ赱xc�ɲ�G�Gh�!ar����=`g�4�Ew5~#V�šёTe��S�Xi	&m�;�(���Ht���&�2K�P�)Plyc�0kQs�Y�W��ATA�M��!��2��D\�ƾF�a#�B�bK�%CV'���R7y�^�0^@����k��vl�5!�jW(eF�ΓHB"��Bb�*�c�xc1�݄���π���?W�֭��q���gVC�h�,,�/XlxVHYEB     400     180h���2�H��v@�4]��q��J��آB2~D�X�(����J�C<� �l�[kŘ��̰�6�?�s����isᯇ���t�S�+�i#���)���\���8p��G��_�nnr���N��N����Uz��5�E����AzBZ�J�{���+@s�v-�����W�i�"� ���Ӥ
S�_'jx uK�
z)��Ĵ��*/"`s���hi���G�A<�`@^��L��Z�h�3MF��
�n���`P��Û\,ЧF2��*/��� 1�6Cx.�]�uT=U^�A��_wUe��x�qR՚?&��cD7�6��"��X�%���(��v"{f�F�[�q�K�><\'
�n��	r/4
!7
I�9Xr >���XlxVHYEB     400     160�*��H�U֫?2~�ɶQ, �v�q�k��U�=��=��r��@�BL�aO�\�=��T�R�m���}j2<��ҁ��o�{�[E���7�˹�G!���H;������<�b�V*�s�H�Lnv�m���>r#oDG�x�r�J�h�*-����iiG�ݭ!� �J  ����|�/�l��]�è�	ԯ�\JI�J������ n���u=�U�x�&��RH����c�.>C��&��,>!��λC���[A�d�L�h���Wa��U��:Zok��9�0�?��u���U�y� /��8�)��?+ArH֩�L��
���DV��H��ťXlxVHYEB     400      a0�M
-��l㾯Ğ������Cؗ�>1�pKq�f+H��k�QV�f�x|�����V�����{�q�x�J'[������Dx��#I��I���.��7T�  8��#E3ț�/�8�S��V�`��\,ޘ�D���.9�Q`��v�N�2鳅�3֚�XlxVHYEB     400     120�W`�@nH�>��&������W�����D��yw/��3��b((F�� c �m�g�)��fF	iSZ������dnd��(s�%�����-���o����C��O����J��f����WINIX�E�%(��a��.�O�ǻ�Y���͞�����S�N�� C��>� QA�P�ƍ�(�=G��!�س\(�����-dk���s�gw�MS��&��H]E�IVr�E��ː����PQ���[3� z��� ⊵c_t�!�/��L�?�^0';��N)�eH�8XlxVHYEB     400     110��m��Bb^���B�e�����/���F%�z��H�<�-�s=U�s��+��UMkHE�q��m����͚9v%����2��u|�W@<��bH�]�W��ݔ�@;Q���B�Έݣ������I�)���������6UǑy�i*E�F'(}�	�eK�E��������D�GJ�i[�%)���q�4�2��uJp�g���:�k4� ���Y�bY]�ڐ<}��o��'g��f������\%<�7���vE��*�\���9����.���XlxVHYEB     400     130�gƝ��AN$	I��f�R�X���Ҵ� |>�탨�G'����2u�̿���<�Ζc]�ޮ�#3�w�u�L�*`���j�C}�J{ɰI�B���Еu*� �Y7>���-� N�5־2+�3�z��,:i�:~�1O��+���٬��js>W���)x���N�d~
�]3j�����ú�A���'��,kR-T\*�"�.�he��
oKS�?�,�N%Dq����s���3{+�mn�閈e����R��+Ą���L���*k*&)�h�vP�[����#)x҉M� YOXlxVHYEB     400     130�-�-�E�g���'AS�K,̘g�&�{���b�
A���"g�>�c���ra�9�3�󔯮i��uH��"|�%c�-?zA}��ӔjeӯED'+Cq�&�ǂC�7��E�;֞Av�O�K�cA��	~�S��F�fU t_!��빓��0�� `�N��;�n���%��VѯJC"Ŗ�CD����;`X�������?���9�:����� ��J�q�Zb�c�w�3�"W�'@zR����J	�D>"2�WS�X���Jk��˨��u2�""5�/�b��Y�;��ǒ�J_Ϊw��B�-}�W<�XlxVHYEB     400     120�2��, ���[
�� ����K0��r����e4Wc_����N��'��f�F֎%��W*s�z�]�8�c�� @����٦��]!�ns�kطK��ށ�%Y&�EA��ny��v���(���q}q��B� (��S��o��Ɉ�lc�\�^#�Qd�P�u�S?̉١�z���}5�۱��/-%?R#�8�N0��>�=�=����(�P�7hI)i*B�w�`�U���$����z8�?F��,��I�ĕ�sU���$P�����A5q�XlxVHYEB     3a6     180w�A�m<���ݮTy�H�/�=y��5 )�9�x0-��g���El֕,�z�(v��M��2+s!����g���6��u1G�����F�+���]�p�t�<�}S�l�jx��,E
��;���K������?���=(��\P!��J�l��q:���V��Ǹ����m@c,��I��wt	�FӰ���L�I�V��m����@��2�P���\��S�:4��3����\�F[��"�}�b^��sl�B�;���tw(���)�k5��N7�7����`�A�vC�SЇ��iY��r﵍����Q�ұ�\�'�4?ہ�&�Ҁ�<"�'����y�K�ɦ�N�4E�L�v_e��/흀�Iy�(+��T8�ՔaJ�