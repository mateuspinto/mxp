XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���S5q[�A ���6�����#=�:=u���/11M������ۉ�*r:b!�*����K���jw��y)��6_��\Ȗ�ğ���n�c/�<�{�q�|7�%��K�qW�Ip���Mg02�ֈ��k@+&p��[4�V�df��x� 2�?�V	��/�A!�|����|�!�BV%u4��0�̇�'Tpm֩�4�m7�t̜�cͻ��f���w�ַ�ߺ��|�@x�eBj�L��7����Y���+�};�h��k�yQ7S!��-�2]`"1��]��������8�n.&�3I1��ќ�C�#1AL=���ާU�*�z�*�=W������̃����M��>X�B�
4���W�Kb��A�B��иx��s�a��m�zL���R'<�==�f(�����F��h�Ĳ� �JW��.!���Tw&�z �����8<�j#������ߥ�&'�RL�
`,�K�,[��k�~��4V���'˞�Dۗ��?Wr���a��N~Y�>�����h-��x��{T��6�����a��\�QNRY���,͓?)��ν�(p�b�D���U���4�w�����Z(c�ą��$EM�X�DG�L\l (�L���$h�0���<_��U,��ږ	��z@�2!+4D�;���{z�6ϋ](�e�8?Ab��V�|Z�y�猍��lt�w6i�����b�<Fi��룚F�Xiju�]j���IދL(����ێOh?�$%��ɉ
 ���(�_&�XlxVHYEB     400     1d0nQ�k�wګ2ː�W9�ն�%��l��O�L6e���*͞���VC���w��
��C{�����SKظj�܏�͞�̫x�V����^�Jȥ�>T�0TU\;}���(��\g�L�'�
a�=:OX��� ����h��ܳ_���/I�0�H^'�$�FA��d�|
�=�#��&��uPh�  ?b�$�;�]��!|�ط�.��CU�W����I�:�'5�S�	�Iw]].2�K�;��y[��>Ԥ2vc�G�R-T�(ot��_'�'z�6K����'��w˃���J|�u�k�݋�k�5����/L�����u5�
 �����0Ѻ�,��Πm�
�y*�K0!/���Ե�f2���(*Tm�˙<MIE 8�χ?����e�}���!۫���ߨ�y����3�sF(䳬��o��;��lf�I������ȑ��l6s�
pϚ����XlxVHYEB     400     160DX���x��?�t��8�7����_���\l����>�(�G����i;��}��^La	���Q���sX ���
'�7�����ꁇ0Mb��[���υ�V۴$;�GxZ���0ߨwݗc���Q��P8��c�߀�����Q ��)
J}6�d�\��ܓ���g?	ڬ�C��hQDv-a\8�?霵e(�Z�[y�g-��[a��%��zn���,��J=܅� ��:����6���.^�8�{⏸��"�����27q�1�P��F �))=���cq �*¸=�&���ءM/	8�ab#�I��`"=��K��$g@��_���^$�:��6��{�*Z��l3���i�}T�XlxVHYEB     400     110T�?m���@L��"����I ��mbr_-b� m�ɑ�'��P�����w�Y-����Qw-��Nހ�k�S���w�Ļ}��[.��M;�b��ʱ��4�h�&{E��	Ճ/^�o��Z����ǒ�yf�PK}��l��P}�S�0�+,��!�2�~�eǯ0K�üb�����2xI����ş�u�yh�%�,Ѥ͕96�l��i\h����`{8Ab`!��-7>:����"��nD�x���ľ��Pv)u�?!!'����*[�XlxVHYEB     400     110N�W����'���v��� b��s�C��m�)|�g?ӻ&ǲ�o�7��EP�����`�U4/��t�2�7Ṡ�CWKΤ"�ɋr"s<A�'��F�[lE'!�m�$PX�<:�5�=������A���dE| ���f�hX�Ts�rFz;=�'mg�tl��GVP��AN��e(��f��l�y��� 	9��H|���u� m���ں����M�hi� A����NؤQ{^dF�T�E��²(���u�B1�=�n�È9�A5[��E���9�C)XlxVHYEB     400     150�u�L���1Б�Y��k��'*@�7?��w�樅����Qv���kb�� �5��[�ʧ��e�woƙ�NZ13k(2��z����+��,tK�ӟݿ�N.������8ETT9fޱ ���Z�-�;�J��ŉ�@�*�L9�bL�t�k�cl�T>�TUH�O$�W;�Tn@�^f���_L�B���3+|4��=il.���]�Ʊ�`�������
B`�K��J�BW��*'���?�J�nO �O�ȩ��U�-�P�7KU�A`�u=�����rw��1���D���l�9��D}4+z�m*���fF3�~�$&�`iXlxVHYEB     400     1903g�˃F�	�W� �޶�p�bk�I9)Ev{B���M�PdF��Z��A�(ӧ5�'����k��d����I�d���|��D^���x�����T�����ds�}��&Jk�;c0.&[4���.I|HKCO�vP�D�B�e<f,�����^Ji�i|6{�\��5��8��§�Di�
# �������嬨��O�po�*'Y�eY���8w��ԡ1OdQ�����_�\��z-�՞&OFEv��1b/�ݎT��I*�Z�(���F�`��9�6G��
'������.h��e��W��l�ʺ\�1�^<T #z�2>��
'���Yv��2����|���Z�q��k���^nf׋+�N��A��[��-�X��e@9/�XlxVHYEB     400     150BE�u� ��4��/gyMF�������~N��M��}�i���j$�O��_{�5M��V��:3�^PE�u0k�:�+�c�X1V$�h�׏�@���*x�mȪᓐ� �U$�R{�e��O�U��/�l�l���M��~=dF{/t���ip�a}e-���)B!�I�v,�+�ܖ���g#9��C�>���O�!���DGԋ�[��~Bl/�����>!�rMZ��"ŋ@[�}޾t>P��R�� ����C�>~��yk�f>�4�N��k)=�����K#�:CB�}no7U�k�o*'�*
��CO�SA(�ki��ֺ���O*8��]�߼�soMKV�l8�XlxVHYEB     400     160��i�멱�W���X�X�6��ӹ���5�ɹ/Ҕ'��S,�`s!x׫;p���P|6�(�Gc,��zט����j��#�7Z��l����=��Z��l��1���"�\Êq������	[��)L*"�.9{;������u��:�Z2_�7�7#�G���Ȋ�{����$�}�<��R}���ػ�3�p���mR��BEv�Xe6�l�!!�p�U�I��?&b����4�-4�Mt��gɯ[J�����A��%��)
�, ,'�DB�\o�뽜B�B�C�x������y�X������:�w�	�yf�z��w�}�²Z��)S�l{��!�rdm�*�1d�'�XlxVHYEB     400     120�y�g&V��'c�.��U���Y�J6��cٺ��'���6 [�/e�T��������缫1�3x�0�V	I�.��(�����"��J����� ��ҕ�6��1�)o`m�Y�Pl����E���i+e�Z��/��ʯ����VX���*	�#d��T��}��Ɍ�Jե#_�}�o��0��x��N�>�����"�M[y錪����(��{�ݚ,~n6��mF?�Or?���I�Ɓ�����[���R ��XPP���lK��O��?}�zHs[�G�tXlxVHYEB     400     1b0n��שׁo)ʾP��mw�@������$*x1XMWݬ����ʽ��)�ߝ�d����ֻ0��e����k��:%��X5E*hw�С�ZU�i�����Q01�Y�V���[�%�&�u~��0�=�sx����}u�7�lq*�zXHn�x���kp��D1!�/E�2!�ن+�iqA��4'�+lݿT��#Y��ޫm1����������~6���8~��%����j��	.��v@w��E�N����/�J`oPO��	�\�_?�V���im��Bw	CH{ET�Ӹ����D37܊Qߪh�.���`�ւ<���4A�6ڌ��Զ���������lf�]T�ٶ�	�ST	��~jP��F��q��w�5�/l���S�(E\֦W����^�]��
F����#�:��:��I�_S��eI9�XlxVHYEB     400     1b0���ߜ�J<8�S!Or�ڶ��9�����/�_��s	�Ci-��?[d�X���8m��-�����
S�P6&�1��Gף�l����FmE���g���6+�SPr�ǅ�u�;�-x1�϶��%`1Sr;Dx���ż���Bk�;"��)���y2�'�^��_TG?B���A?�|V�|�P9�g{�`���F�r�T�҂L�S�G����؆+�ܪK�r�hK���.C��b��72g�hd��̭嘒�d�ƱE�4����i�l9[��7
[w�q�}#L,�0Z�0l�i5sˈ����4x�l[�Wh�.@!���2r7�aJ86�]��'�]��AD���q��5p�u�g��@/�����w�����U��Hx>�s|�W��+Ќ�?7!h���ο(޿g�q��0��İHf���&�CCXlxVHYEB     400     180��{�k�!�e�|�1D�Zĥ����7ю$�Š[���K�0]D���A�,L�:�3k�A���ݸ�	�׷3�0�:4��+�n�(cmf!�j�D#�����_�TUJ��Ɇ�5��Ϳ�[Ο}7��r����Y �P$��P���H�kF*��f��sr��^E������^o#���OXߑ�be�������b���	lT��-&��K�Ѭ��M���4!Ƴ_~GE�^՝h�XJOɿ� �v-�1@��l7L�-�^tB�-Ԕ�D��~���L�î�g>��a�Rwݏ��A��}�r/�h����&��\��P���L�IzdU�KQ��P��E���(vrQ�5
}�l�a}@,)��D$�ReJLXlxVHYEB     400     170 �h��IQ0�&�m@PVlP����}b� $�������.i�r�6W���-X���+A������1>O�x>BWx%cw������|�UA`(�\��)��A!k`P���#Y/}9�sU\��Ww�P�>.�Uz���j�w;����u�|2	n	A��F�T����<���rBdu� *X�^l�[p��ߓ�~��'���S<�_zm����K��e�&n�}�./��#�Slz����d����)A{�G���H]R0���By[�>�39(�����?��xij���%�)Wڙ���Y��I�Yy���-X���ƞ�4~��^���FaA�̃�t�lS��yYr��@��s&��c�؍u*l��?G4�w*v��XlxVHYEB     243     100y;nU�x��J��ns���3���6},U���_6���j�Kq��>�m���0>�u�!.�[wڄ];cd���Y���}x��.�Szh��1+�$��A�d����߬�a��a�r �؈{]�Ss�Z��g������G�q����][G�<̽u�	�o�b��ãM�,��nBZ,�9���T&����i�ii�U׍� ?��l��,�=�R�:�$��@�����0�o-T��|	vn9��Q�.�H�X��G��