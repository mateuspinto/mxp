`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4176)
`protect data_block
aiZA0LITELmgudWjvWwGJyO7VVAh3ARKnbugcvj+3f8qXbCXsGHSMQgkrKP6B6ZXpm2xGXUPXX2S
q5BJ/I+fJNBrUg4DHDtl4JR6ZdeboOlU3TyMHuvJO/XaR2vydww1zNtkXJxnXJqxLDUqpfLoCzeT
FCI2y99GaF/8d9hTh5s9sr0xp73MMyDPiPrcvp+jfSkQtcoxgN/wQTyqDpYTGPLqtPYAo5YxaaLc
brKoXWfuwSUTminQZe/+tf3nFj23byg97CFm7ZbZJczbTNFEVIZCnYrBFMLMl7hMzYdMx+NxeIXj
a6pVdJugvgfHLLkM8Gqqr7BOI/NAX3ZUNdbIfLuJzypjMCJNfOwRSdpV7xMs+gBKAzlf3clEkSU1
KbLDe34x1kjfGQfR2gW8jWNXHgXA0RNl5+RX6jPr7GwGoCo732Lb8T+yhcgbgq7grrKlR6CbLpcR
CD2S3PoiZ5l0LHGkt+lY06lNZpHh5y+I1vE9D1maLJGeI/iatgQl9lLJ0RtKdOybdTRXuQxvNGnQ
4sjqwS0xrDbXPhoRy7FRCNt3dlOxTYHBIrrhhjGkQD7XoLk7LvUtpB/kNNfbw8NAYR8iIn4gkeXp
CkzQTyb+2zJdPE/d8bCx7PVu4hu3S/EykOXneCjdNQ3/1LrBh2k4rRdDmOGfhW2jYa8IrKURZoK4
X7poVUBt2GV2rTQWbpau3CgnLN+31K0o7eLL+Hj6FDLelcKNGS6D4TVtYtCeT6E2Ghcr7JKMFxfm
wS5tIk+qX3JmcsrqpDY/ctcvPTPQPSv83U1dNX5pT1iZc/AyPoSVMmIAadr2VfMUbVipy527zQBh
12I/sg28TdHbGyDGnCJsZ4ieJ8f8EakOS9gPSExBWU0VJSzVfvd7pc3sfaLkywfK81pMROZcFTeI
8HOvgqzYHGuHAU/RqpHF5DbF0KBjhxlGDf/55KUvdP6SDYnc5KokAxK11eMEnAyRW/GzJxOt4NoK
u9BauX76Q5xUn/sucZ8MmpnhzvuurLNeN4WYhRZcXgTIOfzqCi5C1V682WV4H8SSrleCM8xR0rOl
lPCJrjvejKzBtxGWXfhB4o5he5trbYULYbDDTb5Z4UCZuh2gbuF45RQfBRJOedW+pBlW+PicUkyx
EHT/d/hscKaFd7VckBtGRwx2sO+JvsyhPh7Kexfq1pyaSpxIfxDxcip5rp/OmUTxhDo+aSJdij8F
PvgmT5lYTTjR4jAhoYG38IGbgmKgqddxhM0WOnfEMhQzGqSGLjuvJgmuhCaRWMpU+CG46AnBAQ/N
s4NiKADw2yMQejW/RI/rMyKEvPejh+Av67elkkVakzOK9VXay4VUx4YC0WFHX72ZJ2556z6HrIHD
AX2QRAxsw4SzjLxfdl1Yn7Epg26n1J4I+E7oFCJWhM8gQ+ntIbAiY2P8lqy8v0hGmr1fPtheV1pD
YB+q+hgV6Yb7CphJg7S2Abqc51FClHtrHtdxxBGNxFCHLRmhRKUFLcgJJD8VoJv/Kek5eHqnb+LB
hw03WNRyhwvpbFVi0wWe/sc6flmyv4bEpczhT9hzMQTymSoU/F05SQ7CuHYddJGbslpLkMyV7qTv
K1no7T3WXDDhC8Pt8YARqWR8JDcI3rpv1JIJIMDCg2UV7WFvvNqJyrnQxZaERdkd1JbBmdrA+hy8
YpbYt3tbMTE8RGRujAOV+7z/npKzld8WYcOa7b/XvhrBtKN0++ZP9iEJpXp9dQRJX/rjcDKfCjkP
sAfru78rIHIwvLTVNz7ZZ6bZxAEgD8UrXWCLUCHxaa1JPaK4ASJ5JidvWtyMp3nZvWIvlU74kA2R
GcTgMI/gNCE4NDl2ECUt+3zU4ReM6NZWRmptGrjCbGWJeiLgQqSf8CaPhzcpSVHGqMacr6vBnqQL
zl6StzSmnlB8DT2AhQYRjNWsL6K4NuJXg/8IH5p2ZVHbSFBPoAxSMVacrUFIbtG2mm7eL/ibzfvf
68K7exoJr+xk1XeVxc+xrAMd70elpbsCK8ojnoitfS6oHFJvEH0idP25OJKogu+kZDEtsJH48ldo
/vuKOyHK/sGgMXtWdOh8zxTmtOkaMwlLDOvd+iifI2Di4JCGveAEKM8tAp1WRk8jgbkU0Un8ld/u
oHOQNhEKTOTXJdGDu5oErhSui0ysxGS0lN0Uz3D3EiljX5Ew5nW2KwVTmlFox9NfsqVdhhZcnT5J
F7PSrYzHJim+bMJbuX0hBYXvpIt8qv+qqqozxQ5pIQZfGOaXBNhdWniUz/Ib9TFORejSbY9E2Vfx
Wn7unhogzx0FVMLKQs8iERMrvz6emA42Sd52lC+eYbrpah/N/m7JHOtbrMMsYIIdo7o2bn1bsje6
OFvGQ9xhfgTFicMErKsnz1TYJ9caRywYYTtqAB6zA4NtAbvjVWhOm+I1ePQ2iAki1CyB1vBmI7Hc
hYPZ9CktRV9uBjWTm6BlSNW+9Wver/2bOlXORe2UYP3E3/9S0/h8zvYUKIn3l96q+ZaKJogzMVR0
Wb4G6AMZQR8kq68uMFGppFvn9YEKMA1GPB2KOpwCo9wxZ/m7oo13oif25Inrw5+Lg4Pex5yBToEC
VPv3WtZiQ/97/36NqtESorrSbU3hTFDskJtp0CTISkemksvE6vlLInrVYgG3RjvKZBKJGePR7Ee4
q2Y1YV7NCYnmk1Orzg7cn0H9xu+6Dt/ciHdcRudOwY137kqy+iIuPMqhXeWRNGVlcgS4QTG1gGzU
cIl9NkdS/Vqx+KbVlLSAzetZ9cZkxDP3wiMG4PsXKjSFZC03fuW6TrZ403SRWJiHzzkGNwyduHRg
GyOGbamLQsNJdiVpGK3xo+hvfN9zjgtY6cogkvbymBIYqYBoRbe2YBs38lC7xUak8kAXiWVtKqq8
yv/h4GfJw/s/5bZASwYlUyKT0moC4lkFjhVCK2oUxXDDzvclueMBO1vOhu50YazwDgO62dSfdROr
7tmsY6rWH34iKX5NCbCGxyAIu0z2L4bvsZCgnrwNgr2+kKb5WWaJivuMCpPqd7WNkdSomlhdIvhp
ul0jJZhtGhBvEPhedw4B1mjDWIqeZxC/Nzkg5fRH7UWpmN5BvTLmSdlkgJBbTSEtLrz7sYQGu+N0
1iEatW2uwLtXdiH3+1bHXXZjsOSjSPyyxuwPn4D71FkDv8VSFxY1yi8CGEy97J+bcTSre8+9FvzN
rNWlPwJVBWOpJ/d63wCL7WY7pLFLOnj9ekV2IA/8AeEPBPtKXO07WhimxbKh/PIhNkORpRHUy4HA
lbjL1i4JNfxwlrONVClXu2axrAjotShWSlQQhWGtQ8lkMttwKDJHDsBUVwkZZeYxyGArjgssEOOF
0HIP78k+vvZVzS8Gq6iA5gIJ3WxvqTu4Dwswl5qEI6NKGfVsiRenUMXd8CJCse8vRjrT9SBRz/tE
vFRj34CDOrJQgpXbshq1Yw4sowdEDQ/wlk65cuRTDeN5mEr45I/s2e0cDnqK3NAXbx1s4SDjNQFv
HokuRJc6C2gJsGiXvpxYYtiN47R/PmVRI9qrh62xso2zkIWQqRI+YA3M0PutotZCTlJrJaJzIipg
7tkW0aRH6FPILOG6dQoe6x1H6DTT+AM0PkJD1w9yZcSOba91eh+Nnl38G8nAxju/ikyTrerPsUVX
Sq0c540tvT+nj1K3nb7PgxC/x39zG0ZmT14yzYz4iBaZvG/YAhflbm0NnXL6tLfFvWqV9E5ComA1
FnmYr3051RByzjChW0NOaGocjV1yfpY1ZROEVTEuXFXbmCpzBHdx4zo49r53yCO+wtqwgmaGA1nR
mkg59aktagMyF1nrUGN5clzTEmkgf84IM0QbZevDEt5SlQaxTY4wIbnRTgbNCPweATzfCz6xo5cK
eL1dOQVO8RZTsk22t+fU2wrQfmJAV1ATkwY5Vh83t+6MwUIcYw91+lBf9cN/YdCw0h91Jhmgy7xL
P4NtimxWKjyPK1shf1ZetkyVo1Hw0jtSey+lijA188zQjBSuFQod+mZN+w2D5TUPz71ezFVXClnn
dcDwHBlHFkuRZjZO8fEOKJk2b2iAje0J4l+yfESBq6AO7ptuGgeq5uHf82BUsj80GyCMxQqbTbZp
nHqgoWkm9e1QYzNXwjcBgeLPdJkBhZlsmJOKvvhk09aPs7uQVC6M4wCpk/btqp0nEEEhiaRGDEVy
lcFcyy4Cbf28hICnPHVCIsEgptIWBUJEzTxGLfdHTC20++FSXCDOWOzutGE7VN27Rp/r97t+zRdG
R4dJNO/iWqmSkUPvV8bZcM9vk6uH9fzPozpIkBr5mo6s+k3QKUgNNa3mjPKJ0U+cbD6/01h47Mvr
eHLieDi0q630KmnWP+qP/vtINkwVhA4pDNHbWUtihgQ4J/ArwrAUmXLEfdEwQqnKcbhuRCcKyCuf
ibZ96/aN0ilLWryXYfDdXN/ZCcXL/bUSBGdXsPThVGJCAk9FdZf7I+v5cdPsPuEqq9Hffx8ECXXS
/H/foS7+0yZLU6PxRAHyJMYIzCIR3Ap0NjMhVhTFobZJKrc7rcrh9vBKzxbZQGCSneaY2YvbDjCM
rwig9iBQOmP7mfGZ0hbTA2nAM5qJQ3+dVPmI0iUkBmQbRQeXWd40ozYDa43jmi/eUx0LJ9ZLmLUd
ZOLAVRK/QY4os9Q5OLNLTpnDMoQ39JCQ670Uzolsjqxs4nRmhopOke0eTxudbr/o7LtOXHD7hMHM
Cs+xmzCGBmjq/gFuMTV9zdjHIgK44oinANur0rX0JJsR0aKZTt3QRpLnt/LVG+48aCIckl9lQ0jC
xWVcqn3fgJf48ht/l0Xi/na15X7Hr/QFnEGdAIrUyyEEGjnE+D+AzNLWyULRqPllRLIAkSkrn+b6
61CK9xMmAbFDkjpyq593QxaV3ToUSD0+m9PHK3bODYxlSA6cxSXREa+SyEfI8z6pZAqOEJgF3R7V
tAmtQ8e6g9SjVj3Eev3zWXjd7KnhkgV219YgVgSykmU2KFLh/GMWhykC7Yz7xol821ekHMEiM8sD
ZMnRFbnJEOTix54HnqaIsqUCfK/DI5ncvE5pXKAWGKej76++oxJfr+ddsqky1YhDMkxMI4FdlY2n
VMoGNluQixemj/QDtksOXcShh48PIUYJaqBDXz4SWv/if6VY+V/qjMN1xAgyjPypqgzebzYR4iig
hi9rEwmEkvXd6RXo7wTf73kZNKc4vV07/oL9uzWUi3UZi9YGKI5SBFferfiNfHZE7qtZEi35pSY2
DYulSVi1wyTLD1XGGT8QNurWrw2q4Tf+oj9jfdLzHBmLfXbDIU2KwZoVECOg3rp7AWJU6Y3WHQlb
eofecp2+mSpCCgkFA3Qc3RcAORDk7cSMRlb0Ap6RNLrJA+VrytYYBv+NKw0gnZGsMmHFP72S5KzC
qz0mvBWN5IjLfz/zqKX1LUurnY2m9WGI9gcmgA3nfdbC4BlM53zRdhUS0VE8Ho7YaxUFCz4v9PcJ
Ki16/JJrEhR4YghCenUuQy8L6eHNFr+Cs6dtSxIEcI8K6dXtRAh9fQY5LDa3wORpCmpJZ/8jCUI3
UTih8+RDFeFQlxpO+0nD
`protect end_protected
