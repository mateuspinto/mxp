��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���C�Qp&�ơc6wG� �����%Y��N��2'ਁ�O�`�ژ�͉�BtC=>�#os�7�kB �b>��_pd��&ی+�L��#H�C��*�j�ŭ�73�������+�KJ��}hC���-�����kX_���Њ��΢t�E����"��j(�]&r�P�,9�7����]�ݮ�nKˈų �L����Xh�[a	�Iѻ=)����o����w�o�@%�2eA����x'�5��߂<Ƥľ��a[�8�o�.;�`G��oGZA�ن�Y<1U��>��O��#�4!�`Tb�J���z��D@�.�0�Bȱ��n)�D��O������_�7��ϦuWď���}f_͂�K��0=vcЃ���#�G�2���4�)�a���w]9-�i�ߧ��^5��<K��Im�b���^�Ơ�=B�'l�b��s8@�a���°�Z>%I�+��c��QL?D�3w�@�qfú&!�[h�����G��_�q�$�v\q@�R[�	���v0�8 ��R�>\�
U�/�ȳ�ë��7C�6o2�X����]_@tΏS���r+�+���a��v��&Y�=��GګȒ�|���Dia�42q��C !����lTRL~9䀟�q�ǌ)Fc��|�[q�;�w�h��_�$P}	RD�6�=����`dc�ٵV���+�L���w��|�Mi[�l
bi��A�bp` ���5"#���L6�k}��#9��V9>O	b��u�x@`4µ� ��S�<}!���6����2H���I�v~y�NSI,�fXW��?�o3���L�%a�e�]B]"��	�)Z�^�T�t�*���{1п�#ɬEB�d/�v�\�L�S�uT�Z�.��yj��&�],�jʞ����Z?�a����䣈����u�sw�r����1a8	Sp��/  �`n�B�|(�������Q,�_�gz�g&|�Y`����i��� �3gT'�Ў�M������/�3�@u���.ڽ���kw��-z�#.s��Y�+�s�h0G�x��b�)j���A���&[�r6'hc��>T�5T[��,6?';�p���2��Η�9�`.��`\d޲���� }l��Ƨ(<V�����2z����@9W�tQM?;���Ky	�)nV���c*?�Үc��..(��k)����B���G�b�8q٘����)-}mWK���4�i�T��S��p�0*v�`L_R����K���{u��8���0
��Z�=M{�C#ܣ���S�J��-[��뮞d���"�/d�:��-����6w��;��9tq�[j��Z�Γ�
;h�յ�鳇����	Ia����=���А?�U_�k���4���d��h;�XS��'>�Cϥ=�����G�񧃵����%��G��{a�$F%!��Wl�����'���$5yԛܞv������u�����C���bD_�"�����yci&M}�M����@�����
�iV\��.o���&�6-ɦ�X�/��mY�Л�Q�4m^��Y��_���Kh�3W����+Rp�E��nBq���J�滘3�n��b<�~PN���@@�ߊcL��q؁*��="�a��$ǂKѤ�V7�V!�o�B�%�uV�AN-��mxCs�����u�nF� q�I�o���v^�u�� V#�PZ��/�קP��0���Z�s���Je�#dⳟ�S�{@����	��]����%�c3�ZB���y���y_M���Q7�@�Wo�N��G�����k(-	,�噟�Oo���e`��.@s�k;�p_ j�O��2�x���QO�Q�%�\�S��r�W4�h��^S4�G��u���w���i[Œw/é����p����޶�����EĀ6@Ƣ�th�[x����MQe� �3�8�r=���K<J����+��~���d��Դ���>��0��ʫx���d�%5�ǽ"��8�p��.��n�H�Cr�'cVk�P^.�a������hCeM V��^� =�!}�.����� �F i�I0 ������BJ+G2H��6%W4HUw��-Z)-,]�B"����;���h�1��$�����ш�9 �	� �n0X��i1��q�^��Ƶ��G�F4rXK������'l��1���-����݃�9�PF��8�;��{����
�G�d�&űne^I�J���6���������E�n>y�3��ǠD�)	F�8��EZy]���L���f�P�ԍ0��%�*���@��Ո\f��&�c��!��W����. %�s�^^{���D�Ku�D���"�h!�+= �Y�I�D)"��&O6p�V�	��%���u��s�>)�'���|d�ƚ�����mWm؝�-����ȵ�`U@L�[���\���](�7f!cu��+�>i�	��J蚩Z- ��<F[R�`�$�M�JJ}�۶���^��0��|���9�K�t�����-f�C�4ay���������o�D�����oH(TN;�8-�߮�2������ՄG�Q�V���HR�a�ў����g�"�xن��U�	�������jԒE<�݉�&���Nk�0��q~���������]�Fa(�Q�%���YT;hS��YM�T�s��m.�\o�Q�	���ަME"����` ���e���^K �=���� Ƈ�a4�J�b���~��)& �J�N5�1����`�|�� �0��|Z���Z�Q�|�aa,N�6��n��.��!8���=�����M���ұ)�����#Ӑ���/���u_��š8�B�ɝk[�<��k�U;�צ��"3�!�h�bP+�\�_�>X�@a�%=�J.<�&&�o��8-����y��W�T w�!'����ˣ�^��`-�x�6��7�P{vUDw�����)�奄�{�#b�i4jR:��7l5rY?"�.@�FJ�G�
�Ri��$~�Z��T�D��������Go�1�R �?��?�v��!p��e`d}��E*��ӻN��"�����n ���W'�0D�[Ko��!�^K�F�8�I��1Ӿ�����W��U㭈>��閼��8ӹZ�}�	2vl�&�E�3�7��ư��0��A�b�>�o�&�v��m���Ϥ.(F�5-��F�?��J�
8߃�~JSh���X��h�Uk�sy�ވ�N(Y��l%�p��K֭6���P���.��¼���R�;6.jn���=x3༺0��1�u4T5X�dt�m�=�[ʝ�µ�TY�����r��or���������+.x8\}qW��7��֗�o���#�ă�uq8��,F�*g4d3Դ��;�� %O].!����<%�IBaV~�Z2λ����%�i�ĕ�B;a�Y&��l\��H��?�C5���/:4x��08�1� ���=t����!�q�18"�wM$��)Tu�v����J<#����?vԄ�(��7�]�`TB�i�D�
Ͽ$� 6�Q��=��J�D�sU�Xe5otX,DH�iS�e*H��	׺3x��(Ȇ�߾��[Ob%��Yr����\�$r+|1�EQz�L�Ckz,�C�$�Y��#�L�#űP'�w���:E"��&vU�Ȅ�?9�%���iO
�������g
H/�UO��:�Vy#��c�É��C�o�C!z_�V���D|�a>��X�:y�`���.�m�uQ%ЧMz�H�*�6j�@)���%�w.�=��!OB���EO��%�_�Y�hE8,b��n�Q�~�'�NX�Y]_�4E�)�k��2W3�v��m�S���)#򡔄��w��p�'UhZ~�X�Xy��;=_�hNyL����k�<�)�󆠻��iW�a�	�����\�!<��^���a�#�'���?�PAU�3q�pV�"]q|�	X6���w8�k~�u�<�K;d������Vwx.F�Ă� �#���ӐjCMղu��2\?��	G)q`t�!�f��0������j��~q�����h��Ӑ�a��.Ǿr�c���&�}X�D�G��6�/�i�@�܂���3K� 3�FՊ��s��5����J
�v�`�;���I!�tm1#���wˣ�� Ni�L�bϧM��\<}����[el��[(��LZNp��<�G�k�QOC�B�_ˮ
�{a%�-��?�H�f���Pp>�$ȭ�Ȼ��iԤ��(�F�8��(zw��> �8l\y�[i��U0�v\(1����ș��^~:%���r'X�d��l�u����1�ju�w:t����ճ .�?�h*�|6��U�HyI7�*���� QW��3,<4��d��<�K�Dr*�*������TG���%M������#�����p���<�ڭ'��O[K������!����T���sd(љ";�)�H������vam؋���O�V�-f��e�=x��-��07�Fo�Zl{���5�0���$�xhLM���Cr�����~�א��Ke8P��c
˪ �x��LZ��73��Pɣڌe��RKo��	���n�h��D���e�Y�*~���� [�K�QZe�ǞbVV䒛X|@+r�v�"����-ٹ��6x�����@R͋:�Ɍ�BGA�`�9� ���6m#�g�T�z�S�pp��5�6�������d�/�3���yY	
([y��O�)ˆΟ���>�^��f�; ���
ې�_C:y_��6BΆ��`#=H�1��2x���s���EU��n���8weW���ɟ�$F�@˜���1"W!q�ؙ�D�3
���R�cL1/���-��д��U�a����EY��w���@l��T��c�	V�˝��|������$="��k�vB�I��^pk@`T�B���҄�@�w�AE��h��1�V�nj�d�ϼ��F�	�'�ԩ	a�~�P)>Vs_8�D�a�p�%��[b�I���/"���K���/ោ�/&�*�]i�ы>ZΞ+��s��a���$���-1�I���h��@7ϿO2�NC`e����9R�B��Ƈ��>@2��e=_��}��s�O�X)�r�6F�G�� j�xe��u�����]�P�RH_#x�շ(����T�;N����p$�`�vH6{���t��!q52�,�w�8��O�z�?�FzJg����5�rW�8e&�`��� ��c6m��E�s^�1�]���x����X�qa9L�J�ߴ�sS���2u\���sWK�`oధ�ti�7^��::4-��f֑{L� ��Kê��ND�ڨR�k����v1ڤlu�Ԅ8dX����(�?�4B]&`���p2au|�ߟ��Q�g���b�kS�p\��.��o�8����q�&�r�s��3���n�9>��4/�� �uN��\�m:<�ک'�i�8��{��&Q��>�_�c�����vQ"���j(�D����Q="�*h����!����B���X��JD��7+2��e&�H�k��ד�Y��茊g���f9��y���̸7
W���Wf�G`�������X\zգ�;-��<���voJ��Y|���W�NvQ������%�Q�<�A������J�5�l�-��b�.00�d(u�	e����J+�,�mr���}t��	>�V���$�l��2���=d���� lDMnUk�G��Dx�t��������O;�i��{MO��$r%�?�������KԘ��N7�6�BX.˪��=�x��Gz
;��s��DCs��4��[ZC��婙�:ђ3��bLa-γ�v��[r<�����h��W}t�%a�)�~�ֳ��RNkSx|�C�qQ�Ҧ�s�4������t���/���V"�5hb��BA<8��:���[f8ѫ�U����~�fI7���lP�����ڦ�6'1R��j��&{6�N�^���;����l�~`H?�D�W�$!��Brښwlr ��^Je2x����(x�s(��{��x��ҶN��⦾VA�9�r�v�TW^��>iS
���^sv^~�oh?�R4̿^I���ʲ��>��qX�"��z�䱃/S�z�)�N6oj��];�@���pf��(�^e@z��~�	g���j�Oԓ�,����^�4� �|�g��ߛ�E��W��w�:D�
��$;D�e�nt��*�h����99�q�xi�Ye