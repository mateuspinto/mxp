XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����A����3�!+A �*�m��!t���Ej}?=n��i�8c� ��>X)��2�a�!�!�tw�(�a�\�a8��MC�i!c�`�)=�4�r~����wa,L����?�|����ڑ��1��:�/���s����gN����PG�l4U9�*�qc

�C���,�(6r�d�`!��I��ֱ���θZ�۷�os,�%+("~�#<[]�r]���0��΂}�x�@K����C���]"����"O'Z0�?u��ۗU��H<��ܜk���7f������� ��h%������]D0̫���DM�?%����^1{hƕ<!ǦN4gOU�3��=������]G�=�$�1�B[Vy����L9�az�dhmB�wnV�
ǀb^�x��3kU��F�&���|G��m��A&�<$���\�4ǆ�B4�Z�0@��9��h�CK�p~�D�+ 6��%]����.� 4�@��v�0`\�ڣV/��ϭ�) �R�s�q�� �š�ʜ������|����|���j1�קl�G�7NԈ�
��(��� ��:tQ����z���Qҡ�{W��nZ�tk���w�^/^s%�C��8|E��.wHA�bmԫ��;\��)ұ��J
�� �;����K�ry8�d�����`�"L�#�M�^FJ.WeO=#=P�!����D��E� um��(�j�.�|)G*M�"�k4�I�8|d�M:Z^G�x�U"$Rs$���M�n��8�S1��֪u=�T�L��t�l�۩�XlxVHYEB     400     1d0�s3�^���B��������|�Z_��=:��z�*�{ExS�}Jۼ\�*�}���I�Ȗp9h�-�Y�/bEï�E��mǉ8��L�:�/�X�!k���<��J'�b@�5f �f)r���EG��@V�q�cu�c��3.������B��˞�;���wT�u�tb�����i���>�2�KR}��h{��_X�b�e�t���h�>t�V:�h(��5{��}��	��Wn��+�s[
?��%'��Y�˂1������V���q����V�PH_huk�.uۏ�TE(##������o>B�S�H�Ta��kR���:S��n�V�U$w1:�e!��o��<6@U�����������yo���1�x>u�d �>���æ��g��*r�M#"s�e���Z�ߣ�@�ي��>W�X�d�Ħ_���]Y62/d����	Z_�]X���o�XlxVHYEB     400     180<r�x�;�UF��E�3�2��!�w��1C4�٤���#4n[�"9A� `����͒� ./�q�΃���)w"%��U� 8�~�������S������f��1��Q{ y۠�l6+��a�ί����mV ���hro�������=�E�Q�����@�'7y��I�<}�-5�`�?s�������]�43�	�1�îla	a�(�R/�2�%���@��}�T��?I��͗Ҧ
�X|��{�F��Z�:�̴��n���r]f����	S��U���/�GI�uÅ�ʠ��G�3d��2��mp�-y���G�;c	��c p��r5��GVu,�ؽt�}5d�Ca?إ�����P������d��!!�XlxVHYEB     400     140E&��U�����"�[�` �g�T!l�ө��0�D����%�nxH����߹&�Pm�En�KBk�=��M�"@v�|9�=X�7i�lL���̄��ȹ��j�����ž%���X!Ӣ�m��d�U��<:Rw��&`�U��h�")�Ɉs�NH_dƹ���^��7h��<9�j�9��!�2�&kQB�$����Vg�k~Ëϟlk�of�����8�<�w���wߌ0&0��Ψ�M�L�zQ�e���`�V@��9Hz�9ĮghO���6-��+5(s�\�mhrVs��������p�)��^�"	XlxVHYEB     400     110uR=�J�|;�?0��y����0�f�V. g/����y��m|��!�����8\Fh����\��0��,KK������2� d��hw��<��Ẹ˫��V�s�2ZYZ�,!`X�Mۨ��Z#��纵lv�P��Kq��h�V�73W�6�� �������^��o��P��6��#Vᓬ+�|Y���=7܂��g���� q_3���<�+"g&"b��{���%B��R���{2�S���r���?]Vף�3S=�d���&����XlxVHYEB     400     130?b��=�a�l+5m�^oj�� �(�s�h&��._I�Y��~ƍ�_��x ��pyӛ�7��%�f�M�:�p��f������#�2�n��+��
ImI�ۅXs3����	fI|�������Is3h��nO�j�J���@昫�����ĭ�.�\ȶC�q�ch��WJ�d��AJ��M/�R�IJ���LW�ף�#�?�lzL:ed�QX��oԁ�]MD���7|�xƳ�n��ų�������tvc�E26�����M;\�����#��x�����Z������n��1?�ea|�<�2�b���XlxVHYEB     400     150�Z~��%j�wf�у�Ӯ�G�8ݚ���; �Åu�x$�ܟ7�!���DYl��9�^b�����3��NtJr7��	��)��ĔȂ�s[��/��E����bv|l��h��}y2�ʀ���(c��Ei���Y�Z���B�U=�+n��Ѷ���w�bI��Q�U$��i��߇�n��Di�̯�}p7��[�~���'�Lnl�<	���R����3�9���k�ַܢP1#�٣��=�V����F4�dm�����E�yT���6M�o��\L�[������~P�I���Rr�h�DP�Οz�pV����"i�	���i�W�hYW�1��)�"XlxVHYEB     400     110&�(ޓ��示�����<KX�G}���5�5� \0)� ���1�K@��j�ٹ̨z��Xl����eш:��X��hdktnȄ�=�sy���.��HE���V�,�}$ω�gT-_vI�Ȼ��wG�B�őYλ�.�7_9[Â��b�w���U��
��>�Wi[ކ<���&J���! ߌxeq����DQy��1�;��~�㧙ײ�U\���R��xᐲ~����Qe��-��gKW�ۄ�p��@4��_KU*�nXlxVHYEB     400     1c0�j�y��~�{���?UCbj�۵x��$�e�ӻRF��������3/>�֣���=l���ũޒ�>]��4�I�ofQ%����V���T?o��2?t�����ɳ�@�;���@�B-�g���+j����Vt�5���E<F��iq|�aUt! ���ʗ$�B�-�C#�(!��^�>�j��N2IR��S�㮮�j8ey��������]��W�����<'��5m7��d�<{5�ʳ��L���T���U�^���&�����'��7f�$-�?;6'i�e�ƪ�=.��h�g�,����>��^�54�9���e��<�Ye�.$��yd\M¯�?�m����L  �`%mZ&���
�*l���r�=�������0˻[t?��ct�C�UD�D(�b\�XةuXlxVHYEB     400     150
9�2�Ӌ�+R���.��E�wT屡���N�{�_�$�Je'/�%a��.` ��l�C�s����h��m�����)��ٱx�3�����5(�_��ȇqә�����E��bda����� ��-=f*��ˮ����yH���}��Gx���S�e�OIk{T��<X�B ����C[�n!ɀ�Mҫ�N����:V�=�M�C9�����M���df��qQW��'�7�C?_Q��Y>3��>~�!PzK]3����}'w�J_a��Jn���GMRΊ{�3D�Ȋ��d�����]�2%<�>��S���f�����E�vz�XlxVHYEB     400     170~9
�+�I��ڕ]c(kl�v�T���!����l<��F(�^-l���S6#���f��f��%��H.s߬Yk��;��:��|�����_����Z��CCmC	xPmL��Ę�SX� [�N!��BwK��M���P�ŗ��nG��zl����ЃU��
K��I���{n��%� b؎�SS�S"[BĬ�&@5`�Xkm�}�,�Xn�.�=4')���{4I��VZ�WS�=��9�ã��f�Ij���FX�Itw�F#�7#Hk�Q� ��7�O���d�Q4�9s�!�CfD�!bPH=g�KZX�,HU���Hs��S�Ս�-���l� ؊��3�[?�m�aK"ud}O7
4d�1�8�&��c�XlxVHYEB     400     170�`��H���aP��	ԧw��H�T|�0�=|��k���1d�nJ$ڪ������>U�d}+B� ��]����MO)��.��	Ps���<+|g#u0n�)��Kx5̡Ԕ���9�UL��&��v~xc�mF��ctq�æe�'f���������Z&��9ߨT�Zʇt�]J����s�ڸ��#xy�/�Fc����&����O�����߳N��H�ߋ�w�*AӃ�Gg�|��2y� r��	���������d5��V���蔲v���"�N9sH�h��j� i���r�]J��=��<����k*yF��e�
��҅C��g��|K_�*д�WŔ�ׯ������:L_>UԘAu�XlxVHYEB     400     1f0�x�1���+"�c�2PQ?H���3����Ȯ�2����ʐ�������y���6b�c���m�R�������L�"�QaB��}E��b��[�x�Jۣ8��5h>�5�p%8kA�ix�dae�Ɉն�&m�R�kuH�W��NG��>���I�����S@�W�
�4� f��+�=���:���?���-��kQ����5�>�`�J��J*�f����3�sĀD��c')GzT��Ju.���2��X1+ͩ�?6|��du�6N)\�޷����e�9۷Ş �8�3	"Ȕ�/�mW�.ͥS���#���b*�*x���A����9�JÌǪ��h&����}�r�e\)�	G��0��ǭd������f9ZD�5؆l�ޮi���4yK�<*$Q�/l��a����P8ZHn�t�Oʞb�oT��B��&Ų��h�5`Iğ�4<�ݸ�G<y�9L�sY='��Qp/��^5]��k�f�=���XlxVHYEB     400     170��ٲ.���{eR�q2�+��>�.$p��W��Q!̦��}���>���R�m(&Ō�p��.bF��;�ѡ��{�u��y��$�"�
���U[��m-#��R��y��Q��
X	�;��qi���i)�	 I ��|'��}Gk�
��-0(�s���Qu]���dh�JM{�3����$"��C�3I@rN{ᆜ�R�-�B��-��f��#��!QS�mmy�RJѕ�Y��m�n2[z�����G��|��aN��՛�J�������&'�R����
ИC��E�y�ҝzA��}�����	�j���C|5_�np~.ufzWc0�wR���� �ő�wr�^b(��咽@X��������~G��	X!�b)�XlxVHYEB     400     190f��%G��9����=��&��b�:�g�f�#�3�nYixV���a(�5ݛ)7'zb��/5���'gߖؑ��G_����G		v/RY��	%u �Ab
n��:�w�V���p���5p�q�%��ȎOR�;���P��v�?�R�z�$��]3,�"�}�����Hh�k��Sz��@z����z��Y
Ng��-�2���v�P0�=���qh��~L��������7;�"���Ș-� X��W�-pZ���E�)D2;��爅V����%v���Y�l�D�T��
��T��A�@/�N�C���a��iH���tAB.1�^ACtkY��A��3�^�%��E�F�§����(4C�'C�������w0�MD��⧥����)��m:�y�RXlxVHYEB     21f      e0����Ej�(�X#h����q ��]-@���٥��h1����)Aa[��R���l�&�#Ts=���u]��^�[���z:0�A����Y<��z��&��Z�%y��7���P�A�l�"�UĊ�(zcu$���ɞ���l��[\קV#��ݷ�O9K�:����'-K�$��R�a�S��gU��ک�}�n(����뺕9��V�a��5�F3JzC�
.