`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45824)
`protect data_block
aFtwKAssBpdc4Fvmke3rOcC6lmCuC0xT7Jht/6SlR9Zu2QzJzaKaQVRv+S8lCzuNr/RLttoaR+mJ
xQX3wAeIR50G336UzMtNOydOQww5OL6sATo1/TzcnW2/vDsZ49ec/KSEk0glG9v7lFUmMWOg8pmL
18fM1IsgxMWwmJLCGFmjMTLgUwX+X87t7HVjCy5lWMwqYcgv/1ZWgq5ncdwZlZBBHtjyWPTq4P59
KAOWOXwScq9I59t5o4+8RGjD3tTXmp0V3+XCfyW6KQqCLhVTSguDqHKurfByqKFnLzJNgIfTY4al
K2x5sii8kTVXF8AYZ5S8/M+GlQAf0H3Xn9iGv35YqrmOA5p49Xgc2M5WBJvAirOy6Pn8BeWjiVuw
YcN6wOWMYT7THWC1fQtepW6218Nf8oWD72n/mXQ6uIlr7asHzzmeWUCROFfkOIR+nyDCRsJLVOKz
XdII17FbAUO/GTAFCRPEv+clInhs3dCy2NF38JmiH6GK5Dyx0z8pAH6Ramo/+xMas5MCegMp4S7D
hG+M7Id3mTHrRBEULDNEg1P2B4H38iL57me2ICmpPRyryXmypHgTfUHgIb/ecgyo4WvUM86JLvLj
1O0F870bD+RCW7PjtYg6Chh0aizbELSk7WMk7c4mz8slcQVmNmJEoK0C/xU+KXqLQAhptxRjlE70
fhbrNTn0IoJlorBn55+WeU5ExUlThjtUMZx6y6XCtesuxjkWJMwvH1LujgAwWfSQzYPF9Pf/zefZ
d3ybsUTUqtKDqAfCFPkNYlKPE+BIt+x41j86TD9akOPiehiQiiTAHs5gd8RfdOCPRo1eGw0fj6KU
+MpvTPjaZokA6BKyeccf7P7cwgChumsc5ab1u1ORykM7qBO/8fQaC6sJWSDq/3ia8+lg2BlCJFZx
ENLSVgHFqfoGOnyr/XDPqlUyQI73bFiyf+7j5T8afFhhkbRpKpwcJD6GNcNxKENrEPZqimQs92Y8
4R8YGtbbxVB8JgpNmlauK+FfVUaIxi2wulr4OnMzExck53/ePU0ATcL3LG6oyOLjqfliDfnd/4GH
cWsokiobFwQcKzcQXxceY3YjIP2l7G7nB0/b9XkrFunjMjr2FPCbHoGIxUs2CUauN24vZATBLqav
6jubCnxpWuxKITMPxgKwHNwa84hJo0fWNIoYBrkZxOjFUMtAnjgd84odflN8LclehWPypPcwJxUW
4RDOJ62axt7bBj2fk+p31S3s79+r4lL/7W64e9exD4d2kPzP5xYf2s36iZocszpbVoliWK4ac43J
0nTKmMee9bGQ8YR11ckaU9RUtDLNsdjjzfqKk9gi12grOU5zGU3mK1fnn7uv0nVrGsaugr4cwrrp
x3hjOMLtCca9PCq0cf+09JtueBXaEL1jSdtEp6e37owJgzsH13dwzCxskJEgZIu0uTxKyNirWZoX
3fCeA/dEj7R0TtK1UP9C0otAbvllf7R/EoqG3Wg5M/I4Ak/RvIOKnMfd0++/kCt9xNVC7sl4ApqJ
1PIzqbngeaNu2SalC810EabSPZRheU7tJRhUSeg7dIO0zYlgyHNFvWiLHJnzNBOQSIvNrppAfMBC
nsl5lI9BXRw7fQ0DTDj9yUvxEEWfvTPIfNV3oMdo8tjxXaYPX96+qFdfzufL47n+pIutpf5cI+6E
k3nlju1JpGgUE/W0Ovou31Lo2/249cnwioqbBnBbHXnxeKN92eT/hYWp9vxlBLiXF0MeMSGNHPac
/8xrnns5JYWOcT0CHBmJuYLAea2BPVJMkvPsUR7gVQIjKnQE1G0xY7wiBWfot30SdLiZ2YRridzE
F/SbUjSFBYi5ui62gCCo+YOmriRvCu1ignxpueg1lNIiNfKMPf8zGay+UFXY7uvedTaw0fAQLhUU
S0I3KIQP7UwG7PuQvrVOvbabqDerxJyBbCcnX/MtRPE+P7rnZzUoHOm1AWiDMFfny2DllOa7JMQa
A98liUVA951giea18C1o1f2OykZ2aJZAUheJ6SHRNlYC4qBLVUehqtXy7X0vblnrfLZSekxDFdrJ
Ab1lbFHRRuSDfiaKsNKyguWLkvvuuwp0xQjsaWdFTTWqMiL9bditoz4fIGd+S3VnIiOrzcs266my
QT0S8mG9U5QOhHBw+VHFo9Dqb8tLAwF8Jxh9ESv799otPcx1h9MXHaSlKLtc53vPN0g8c2VcM+Gv
dbd5v9AVHbSBQKJg/W1AWt0dxm+OZGdKo/8owVBgzzNDKAOjC0MfE1gWW8kGOBotaRvtm5RasclZ
r7KwDvH5ucixe09yY7pPqId0iBvqkcQCfBuY3f8NKThiKS5F1PhJDJUd48ZTeWqDw2h3mXsQR6q6
uzAPtyyxdThw717gqgh8162NfWVUV77+nPhXT73St6bAFKfQKNafEoc8HyFiMdcUa0QrgfwP/X3k
f1IEZYbKGsooH0GPE79LcDPui132xp7vCOERbrdu73hwBT+utS2LCq8l9UsM5qzxKiRjTBxavY+v
WtaAiY2w834nQDRnBMMiYwm/P4omssu/munw6iYamQqvbAFGZ2vHp+JkgNkpvivH0z4proox/rtM
TUYo4wduPBYa7Be59W0hu9gTnV05LCqgBGO5g+MeTGBQOKL4QLczCFicVsh1vDGSbT0/nsjWjtJl
F6attBLeHBgGyRitHdGPgqejb/T+3GO70XSOfIG8/cei11tnzZ7lwH7e9m7vaFl5mTp47pSi41Ql
iYFXJGbRJ6ACq+5sQyji821rnhtfz4Vd9IEIrciBdvOJOYH55j1UVF3eCM+Me9PEVNXF4eiZzm8S
cOPTZlzmPNbUQXrLNmeplgEDqox7pHR5DgwI8D+mSVvInw3bSdatQcccfNXw+ERoYI88Z7vRTr7c
unYBbXLlAwV4PNOmWqRs1OchgHsd4ttLLqR39dR6dBPWW7j2G3PYjKUbu/n9nP23YQPPlOg5ub8N
JCblnDEOBDqjWhOafeHts1BBP9piZYM8Kzzu3tmRaqrbfGk38MGc+ZIHJA0ucLBUhUzuYi89rekx
98K/FRsXlO+N1qhYbpDYNOoC9WhZ8+gbQpJLkh1C5CGFdVgqrGLmQmesGUwU6NR5GHwUfY+E+T/J
le0jP5EyaHfX5z2S1o9DWG0Rp2WlTlFDkLXFpbPBVDIbbf7kUw5guhCiTnOy7dbC8O+g07TYjbC2
fxVg8pg5SsdC1JA/xdI3TSCECtXxwQ92dks6cPrqCxwk/xrXv2s+YBM8ZLUlJyytkqMlV79IoebL
50al7+LJ3vW/AJAnXy4Fu1dwN4GWFKXUxi8hn6HK+SdFKaobpTNpWUdTyAx9iyWVDwd3W3a8OF5A
p/wfjoXbluITLz4/bZMnrs3NzDaukcTGhg5XRbN+x7mVGLX9GnbAEmJufRBIedjIlH83q/chYNIJ
tIg15BrwngGnOr/CijIqjpae4EfhBLwuOPZuWvKA0syxoXsSokStGVwBuE8PSgOLn4m7orGt1PBK
qzg9XIFlP0QP5MMnVw3/FDxSIgzRBQSBuk9iJmWA8F8P01Oo1cnHsBKJip+NEw33T1qKySKLlivF
Ar4H12433FiTZWFceQyGWVJRieuVYo4votZKEYl2OMDxNizEDZkiplIxNQMIybNpiYDayROkMBos
omnD+akRJ53JpLqEtmfOOIrJ4eRMXDyUDdn+vgNHdeTK3vGGRr53pmJ0NVvLojO6q8S2ae9uSjPz
T8RDT4XbWknD4ZDFrszPWf5nTKeCOpocr0iZVZxHvKL+F0etTAQYupgnNtHIBSDyzRMejZJI2bKo
pGIzEAXCVl6boVdv8TBQnoaQ25Lx5w04XOjTEUXQG/eCgkzI2ktjHADgI00d5w1PS3CR+/gpMQT0
i8GSQWewGk5THljFDVxidOksfuAgqqzVH6KQHBCsbyXcciRgLV2Cqz+R7Hj/N+iO0h4ZlSdFSL23
XDQZAezk5sY5cuRXqpCCKkdeEWeGHWs3dTb3NNL3oJyl46MkZKjPW+YUBykS/BvhGU9WrwBcfghs
BoIu5CceN8VtbzARlAk7gX69/BojkLUUDyPuGPQhxsa148PSDVYRX4v2LGARj35JHucMydfaVVoJ
6tC9tlxS5iFEAIfR/JAfxeRganbq48RZU73wPfrKR6D+W2xlQZz54HMochIdyWVK11k1ihh0YlpZ
WuSayEwTUkjCPjPRG9n5A7wOc8WPbsI4VuzcQaz+a03FGN2wY8o1I215w3KjzqlP+7iIFKm/hPbT
5Abw6tQ7LAvQNh0D6CaJPaQLvDsX9BBDbTAJP71zjanCxB3/VbJXJdv09cfUxM8N1G9HXnrJABEZ
i2geoVNjtYRiMfHVq+vNRrNHbUGd7ZUwO0NW7q0bvzdB+DHPOsvYAwoXdVsVm53HzKD12mhesYgg
jv9sBcpMsTcaQdJ8QWUUlTP04NvYivnvBye9AKlrUBa2s1UuoM99xhmEeQqPPYwzbZcJddxaHvCp
6vusHpc9kgZwj55QRXTtHbUG+dsJOKhnIjTrzRXayXYSUnF/Y6SWrDQrsyPkoPiFs3XSAyGgxeOp
cUInaXR/FtFJ1ryIwl3A7oVRij79nPPWlT35Qn+6dA16koRzs9Sp9C8H3B3iSNnwnebbBDYFQzSI
cDWQH+G5JXgOCfW2+zG5UY27LMF3KvQzkskgwMBKywuCxkLMwzRNr83PxmBRp1TE4TQcwqIDm4IV
JU0GSV8jDq2Om9OmoaFQ2TnsxyVHlzNKp2yf6qvyEhIGLWiKc3jpAIxvycrGSo7tVsTpqPhcE82P
h9PQKKU/blp4RJOfWI60O4dg6W8ygX257ZwScDOCIaq8uSqAlQge3o89bh7+kBp32zchExnb3ciM
e6hodnCfNQ6suCGXi/uBZDUtb2m3dXJx9B2WVtYjPNot2B9AwphFoRfZX9oLIZdg1sXz9ChdCSfh
5hFe1BqDZvb2VBArt1lteKfEO1z0s0qRFq5W134WfECoA/g0E+72BKVzNDC3dCUPyxzyD+2ogJaD
HBwH0ojgq6rhn6si27XLMKm18vx5wKVNi9juPy0TYGeWX8eMV2my4EcOVjnnVSF4pVPrlo6z0Bwh
zz2xI8ZU1V8Gs+lkL50a/8McUR795oZfpOT7Q/H3iKLQfbg6F7YyMUxrtjLxz07O6k0Ut8vXqnlS
LT0IWpzWcJW3RlRVP+Hbvzam/LjF3O4bYg/kzSGVTRC77TiaUJdo07omZrp5CTlZfkwqhGbRl1tG
NwvvBQndwsOlaqxPpifRlgZ362sVXcdt5fXEYhrAPaVR4xlhMlnu2Iz5NuZwF03x0aterK7nWLkY
Q1g1ly6sWIwSW+StpXCzTEx3cqD8Smxg7GPritXPg4lwt2ExLmHubVzO/Qnx2ZW65+LmrjpGWn4l
C4hs4/+9SLrIoH9SRWOA7RhraHpoDqhi3XQb1+SFPq7BFv9jLWxfTFYvKsv/gvx+qB0R4/ZIeMHp
pwKVPHfAhv4CMW5Wj9gtK/n2LOSE4jJU86RY+nvbIq5RoXguCfvsCbp4kxeYFtQwVFDmJ4lpBHPn
m8oakToL3M3R1pasAu8DUX68HknCUBArRZ0qx5pBHXCCfoGo5TiVj1tVLj7X1BjiEN6jhm0RS4D3
SQ3dyRmzutZSnuVqmofxmJQph50W4sm4wMkuJ7INjKhYYMulo5U2PW9sn+s5USXGYPfjkR63fKyq
dJbjZuo5uXAEXKhaOUGwfT5RT6zd62VV+jYKqYNbff+HXdj6/V7U8k8cgp5jO9H0EV1U9NlAmuMu
Z/Pt1jUpJtF1h8Q/eQ9ssLKW1+vAuQzRJSXartIaxt9ye5K4yxuizLSzqDJ0oRbeNrApBdozoV5T
9I7bnuBsk0KfcbyHeJscKjNNrEK8s6tbBoBQN6AUDeFvJof+n1hO5dpeBrB/QZBn8uDCiYzCTGJ0
cmF36edBlE/sTIyUzdM0SVVejs96JnrPu3aWB5CI0DspTnEAxvmEJvPkLWkUiD6rRPsHpH7OhAne
wiYuQSQrDnFFo4Jjsq/sVx/2NS4mFgnKK1EiCwjq72v4uv55xCwoBsExNZxSIcaWReUPQ7+L7ntc
qPZkDR0UHzgFbYz96+nCwQ4WRlAomAPE+wL6UL7Tq/SDtUFcdsSzEzKeq/9a7cZiz1lb1ybdIFUw
tFYl/7iKvzgAjxqhdfvhMM6870CcYt9kVzUfpggjOca8z73KojE/C1KzsU7TTPVMnz1WRxkgj38P
LyJeflrqAeCLft0dkjns/Rrcln009obgBnIjdz7JuwooPuw9cTEv8N5/AcQKZK9FgaRMyAPxOhci
fcFfgcmsiim56p4m6dLJogj9OX+fPoyIqrICUFTu04BP9pB4D9Zd0BqsuQkZOIl2UzAmKOV9CvzL
PMLrAO2TpUxdlMUnAesfqljNG3144A0o6GoF2iD2EkYjnU9TLYpT8B1oq9OwCOGQr5W3MB+TbCON
+L1X8OYleEuZyKKRsLaLc0gfwewXMG1HhzvW3ThVOm3PO5VhVlgabEO6tudlXtIRrInu2zJro4Cn
ZWQhs/MxgOvPi7KRWbz6Tq4RQw2jWXLnjwIOLudd8yT+Yjp9VJZyDz2WkXCtqU5bxF+hSoVB7qnY
HcYXbtmGFF9YmwQr0rnQ3x8mTH9JzmwfcNhG1pruYXOxYeyD41jinU+2XBAn92P+1PMHlnDez7+g
+8XVxnJbBUlBOZvxoJ1haROx5LWjw/J2Wo16gMZyLPUDUUkn+wiPqR2kEz+OUI9smprlT8sqiGe1
EA49/bG5pu6BSzsxgrat9jEW057L6uiDH8I4oGjwzSzaFgQFjYx9blRnsWi+Rm1AOyf7+5OwZtZ7
QpROIqpCR5hgsPoGp6PqqC7WG6FSyJ2UBEYa6FXtSuDNPjc++K78N4Bq9bP24y5JWNszzjdx8Grm
dY7qyvplZEXMwEx3tD/o3DOL6zt/V5dfI2FXOdtSguk8r60jdGBTM6STSGExa5kemezC4XFnIimG
2+JJBrJ1yHnUxPQtC/4+8628oiQDS6l8J4qmJvOp9hfrOuI+99z87iWsZnqnBwbhGeXy/FhUNtmp
IM72bP7+SKKNwL1TMTOI8jeL4W3GOooi+pEm4v/RO1aTVD5gDOvE3yJiYjmVv5V4aOofR6l31n5p
AWOuP5JwZrm7dV0RBpSj973X+o+18/3I4fkChrEvxHGXQfpPkYQek6CgJqE49CHV1lDoyyoS+bju
EPBnGY7Yu2i1XHQR9Be5YSwptw1iiHjhKzI7U+o4ckiaKG2RTrdxZj0PuuMsbO38BqmD8+onM5HP
9H7gXKwG0tOCXh3hBX2nnbPL8EY4Y4MAsnhPaPyhZcuJITPaCblxOxeruFiB1hevXaHZgakfGf1R
+BkOgEkgvKB//B0NpzOQRgWWweWxJRVjgqI0t/2J97xkvWlFY+TJ0nWr30p+SsR4t+bbX9c4vttx
/WbmjvtbuyZdgWaPCdCnr92nWm5HStzkazn1xRcj9Wt9LkAth9g2wh1C6bbn2mNv/e/m8JlRBSfV
el05hEs6DlzDgaCBWQstfOfWelDRdETD19SDQpQ4ocitBRnluQW9lkBIlc36l8O/a5V/0v3THaX/
xLT25Sq2xzrDXXVs75CmT6SguwZUG23r7bTAK/493S/u6Zv8+JJjmB0kMrjeDKl3bBvTCFqwsw+J
n7olU7h621XTOS8smS9IzeahWoE9ikoo5RfeNtlT7hGo/4MwOHkVqY272r5ImFiBv+bJZFwI9lVV
xkQB24RcP/LKv176wboMsOLkcwLSNYlW8pEHIoA8AvmDPXouOjHLMkVPldgwN5YbLQIyd5Pv6LMG
qxaJltSlT0847NYV2CpwLPUrlbNU+yPQ9yPGoEzPrjNSJN9+S7N9ncleYtaVuZy4Y79d90tSGnKq
GJehAmlOqcgolDeQZtA9SYDWaV956qxo8w+s5caax35B6H37j3x0fjPCbKO98FyCwKzi4MmEEKAC
TEtXWxXPwskS9ZJhx1xIvAXatoMuA8CH40NNOIWHyghkOlCH9HE/Wfkldd5Ro1I35cysH5IF0mJ8
yv7TjBdDV7y2fa2SuY+pFm16xH9wcBAqeAszsvI9z226S+SjlUyLmmzDRnmJ5wJmI/3Iyboeljxd
MWnci1lncggv//u7cpJcj/y9emwG959uZFBX6Y2MMxCCwpWmofzkXdqHa8QFuK16Rwm+SwX+LcsS
OWsnoWupHQB9bcvwRri3Y2VYa+pUy42JPKT/Nf9RMSAtiBh7gp++ErImyPo83eenpsoab6vuk8yu
OnCKzWzURr3k060geJzolbJ5tZK4WxU6jyBasNOSQ1PC/AqNqgwBoHVt36hPwG4RKSJEH0AljNMP
uOfjPgIVqc838Ig0Wn/1xWHwzXVpKFCP5PHVcVCJl7J+o0Uo2ZmE5swRy6Gvl1QR9W3GtVr2Z9eB
YSfCelQRXTbH0KOeODjfvs1fslkleJWeDaRM1lpBbC0ROc0oSSFqP3t/TfFZzfWv0TwXXaA9V7Em
oVkH3gKYMvQy3mDIM/t+Z269d1oIDQvgpyAKl/xf4gJeF7zrKK+51/el7QwDCV3HgnjfVS4WIS6B
T3f7eEtYkZ3xcZlBOKPMpfRzAGRBh4U6pc58H9Oe6Mezw31v3qPut75/3QuE5kuMHt4rgcxxW5iH
ZcPd5Tf53u3+oQ7kJ9F/dUX9rZxjC3hDjRDfkL1TJad77GteYGq9L1tJqSs66Pe26mp2Fx67polf
dbDdu9DvyK6bSGbJGXFKOk3OcnUH532HDQUvIXdGpscNWWeONJTklNa6GbPQt4CC1AKw8k/dJ+fd
l/95KnCGA5OFLqhwtkQXDcLrETHEeJosd7Kd4KJJ5JlQI59RkSR3s6OrEWFRPLPWXqV193Dqbwu+
6n/AqNaaW8g47mVAK8MgOfpm81ivZG2NV/0RUFbNYQJeTTUgBUtVD/TlVGIRhgezM+bMzl8QGsCN
1oZpHRa+obKWSEhhUCwumNIfhGaVR/tN8JCYJEGm9I44WHBJdmWga4TlplzRNd7749YsiLPY9SvN
iTa1/HxXKEZZrbAAaV/MccjmLFdQw3WjMfo75TPLPdfwpN0Dd37/AL6fQP7qeUDhC+nOdwSi+pXG
FHzJ19kauY3Y3LDfb8/ESTB92oSGhBwpGvFIB7gsMscb4rpgfNaTBl9DxNJqncZ/Ngb4kzzJVzjC
7imj9m52DFRwZxzt2B133gkwUCBiDfMysazzBverFbLSZoNbYIMnApxitUT47hIt6Uv4lNos67+K
nzldbX+MPYMe3uith8xjzWXqmZWrVBzL0ikPzcyOtrS5/HXGyEH5qKLFR8aNNT5SIMt9CroN2LU3
sU36d5EV2rvV2Hkd9/bXutHc7gqcHgD+1hHK7PfdWOqXg810/XASTsXbIBClEd6qaKaQZvIISA8f
r1GZs+k52iKCChg90s+weaeq4bQ2t7NsuVAS6NjW1Q9oFobJnO+wqCsNVuBfZZVnp9LHKFIat3sl
gS+qOPXHHAOD9h7eifqZSHEToRhk+SKGpK8+okFFsfo+5vjs+JVn9GEEzSq4InFaH/c7oIpWTNcL
16gdErzW6r8WUxTGyuOBuQ6RIuamGnvKOee4BaSqF1jJI0rflkisl+/qDfTul5g4KLmKk/B5AbY6
/vNc556G2Jv7fF/6s/VBHjHtwtrKLDmwsvglmsMdFFVb8IR62CTCNgqddISnQGW17hhtaa8kAKmr
KoEFYOxg2cv9bPaFZED9QhxGBSyV+S7c3cX2NxN71IDwVyBJkZzXCzgUtI0eqwmodU1dLK0e879N
P9gESR3uI2m6MibX/4gL5ekOaEb3ek/fXRzXH75Z83wGKN6s9tMTk7u79rTs1baoIcwwYNPbwNca
3Tl+U1VBEcdsccBWXlgp5QMKK2Zq4kFD1mAoMoM30bBxQTR3zhJKVFevY7lizUEtzAuf5BfetDQQ
cm/DijnLgJXmUJYj06gtluENSHiq5nFidrw0zOobwgjCe4GDyDDXSWnn5DgEdJtE51YwAx3mZW4i
0XiyHt6b0367HnPlYlrxhZvPhPaylXwDshHgCvS7T8U0Y2U+wU0GtFlCUhSMSIpGZa7iyZIznXAN
/nInTTFVHIH+6zzT2hxO+X5t86MqNS45aUdqZSRoN/Bd2KbB8+sZAaz+LP0gN2341F3o1OvHnCMw
ZEDHyE7oZyDIMirOFxiy67TKnbSyAxjJ8yKmMU/esQNhlogd9/gM6mY4kzfjpzwi8YNqSxjRVJrL
86Blhjzva5Xw59RbJD2ee5ujL7z57P1gm0AM+LZ9VXnvBb3YYJvuQ73QeKeCynyb/NXIjt9yOGhj
6fwMgiXl9qGkKuTOOfC5MKVXaB7t5u2B/Cs/C6NSr+F8KWGkmgbljUR60SFQaTVS7DaEVTvtEb8O
OdVT+lKY+tkZVT6myFqFpFp8EBVG0nHx46kSdKkSlGAGsMvh0Ikun5c1MaLvCdqE0iawW9lEtsNj
0UBz1Npi1G9q6QLKcse534nZwsbcdCEHceV5reGDVbDOKsa6Om0y65nfWKJPuNDfInZmg9zALeEZ
E9/bjRMfNDSq6a4OxnzM++cNR8kkv8YhoMKfJAs5xbsWs1QiFnJuGIXfnvpQJ6zoEXV8jiYZIdec
8bGNrNa0RnUYYj1jn0yCwsauDFKsz+u/zWa82urcIjz1lCpiulaSyeTgII0rTLJad/iwnyo5cqJB
T2D3je8m44PcnJiK4NpzUVZM9xoUg4wEAD5cupKT5DE7xr9S65Vlgy9QX4fY5ZTPWimLZNeghcCU
NFyLuzSySjurZ7m4ssTmhXJ9YguntrVz+J7rzIRPdlB/lDIrBhsDaHc2ZF4CYX63oHyKqRF6Cdtl
9PC5X3zMUtsUhc/5LgsU9VLbRAb7mXQz+OD/fUlTPpTZs9cC0HpBulQnxppLgO7QgVCLeqD9HfJK
mguPSdluvscAa+w74DOuqDX3ototLhQhISGTS5FbrQGSAT99Wv+Tig4u0sfItWEMZHPDLNB6jhXW
9WEKU6FFO4h8sQDm0EXbvJKGZfvaZxoEtw73xGyjQ0qUV5uw7Njcc9U4TICJtBB4x6TJYlTEv0u6
niCRPH6fd6XIcou/9upDok1K7rUTZr71w11ODTOFXueJzaZoJHnPcH7PmxNtl6Ti5cTyH+8F7z+o
Q9Vxr1m95MPLExoq8pJijdOd2v3msL+bM4f3dDRp096Lg0eCOLOqJyUnXsAuJz13rwf5XWhYwGuD
ZrjLWCDR+UDvdQlrjO+q3UXleu36uDraOlfqc+iXFUH6S94g0R/9iki5QzJwetmqwtqkkxT4DBkN
gF8gcIJLcj6ePTOEQRfR2vVcJTaE2H1gTkAI/q1mFHt0DyNxvd4GqsKnqZCdV4j/Eab0BATuVeC3
iO/KqAmKwKPAx7u6Vie6qBQym5yopjdD3ZhXf78WmlagXBNItl5ZYTntI/Mmmcz5MNIQSoN5+i+n
Z+P0krIaEo58KV335VgzuOhHHHxae2yFtkuhjn51D0+CBB/Dtcpk43mdDbEmwzwcg21LS2RIFsev
GtALsOhBVU3Foh0UdKi/yRbtwgpg1TcDqideaJZNWrhi0pgi0IBSm00YOYunvQoaCD3MwiBJSWdK
J6ntj45/LGoTpnlhr6EVf1PDKZb9X02fViH7EfDQ2J1u9Fw7CYPxz5g288afoMV0lBlRWXAMxeqy
Zc0VRuH91wyaFQmNOqcujhE9qX8n9rRmO1BUPU6DiqOFi4xs2y4t6dmj724XVbIc/5aQjFiVofLD
IGrCF1NOSwS+R0jwyhNMq6VX9uIr+Tf7qjMuNbB1Rye3TkVDermEVD+BHthoqXpLRzb9xB/q90su
ZaSN6QJvIyhOaMrnRHWZdUkqUjqFRiaRri1ij9r0xzqDqHupARNFAE003RKq/BmuJtFgHbYss9+a
INNmNcUFBRvIBdYDdppyoyR22tlbYrNfV6El5bnezT5C6zXpMltjhzGGQFlb9BSMD1P0C7AHOumF
eIAzw17eg/WZiiXSAZ1vE21CPpL9yGha/+ERjZz2KwtkiZ5v6OKTT44/W2FlovmfKTRE5l2QI+Ej
/yicFK9o9PINAu39piJ5xD5rH4phr1RTickGkcFNK1eUPgZErEIXLkOPDrAp4DRCmgXatHNeQ7qu
BR/UQe8y8nywsFRBeMl3bzF5k+q8jMczJacZzBBgA1A4U26RB2ucfUgvu2jCMkGyusA+N0Hic0uB
oLFN82UdOCUGE7LwJJUJGZgrr/qT8unA2Fh1mSMEeCon6iuBTpNWZv7CEmMFUIpMHtJuXxPkjo66
q5AiOu310e9Tty5tdS9794yZ6qXYLOwT2fOuOfz+wnJnbKIJ5W6XRKVpfXX8Qb8h2bYxxrb5KmjG
uNZ9xLQEGyPh0GECUw6Mp4WXGGcSL48qpMoQA/L3F+quU/W9T/Gr+7aQhVsPalp/1AfVuI8qio60
HPcUltBNf7pKW6UJls6ERvg/Fwd0NOVzo2Lj3GnbsaLxO6UxIzxI4jTPJNkTOfEIKFsWY+tX98O5
IiB4adEFzWagkUDdj1DVi5l9lkZ3UfwFzZFUXTOZ8Op3gNLVV9VHJ/GbezNWRbEdz/xhJM0marQG
rkd6UcGmu3vVKYNkxOZksYkL81NNYsZSDRCbtM4hA3KoSSVzCYN06xhF4Mk7qhLcHs4vLfjxrpDN
irdcqqzxc7A3zbRBYqw7llMlQV0VcJw5FjH9oqKivyz7S28v3nMbNtnNudRiorROh6Yjut6SsAjn
EcpAdjwuehWruPzkBsldZN9Ir+ms8mu4BgSgJ9q3Iehdd+JQMLkzIXw4RMB/QBJAFhy6vB+oh5IA
k5RslxxOtE5ZEhu/RtQFRO2XdUGmHg1oQfB8iR0molJcnoy3CeO1lUVdVrBOvj+X+i6XnkDvtYQ5
7AXqDmmgADNq7Ul0kuyjv2rjdIijUWHC1DdOuKssf/54fHdVmg7yxaOWboaymuG32W4tnT708g/x
BVoDLtO/Txj8FVglmCJfDqrRo1sQpN8RZFVdytBAsMI7qoLrXh/WvJuwvgnLRiuz3WbpXAt5utOH
drT+1JysjstR2uibfEHfXcX6z28Ads8OePaTQit7wyqdvdSh169FVc6eMR8ZYFZTp5z38OiL4+fm
1kA+QBH27txZj58woVt3RaKtMnoCqzXWOIR0dWUoTDbsLfcJ2Rp0E+jAY3LZyfucIWMkzVi1udEy
vYEloy2PuSyT4z0ZpLgU+xC9QhXa/VxypCdQ+BB0D+PU7xP+4o1674QZNUnOdD9Q1dBx1Y+tZmDK
LrPixWWUNm7JxabZsjfm0VvHJD/U8tji/HgCPNpTWnDqLfFZV0RNMuTtE+6EIiCtYiS6wWliNJzB
nmmUNdk6Rvo8eFpxbUyC5uTNkP3yyPD0HTeyNpZ6vLwV31DbXTW7u/qbE2FkzFrllACdS4VGr6ZK
srey2FSWXe2mW5WctkyiyJ2yTWwPbc7ztDruAtim6R87nrYQkTIKxQzQDdTHTEv2wKFyqzXgX2DF
7zUA7ItyCJWe+UJNI4fyJy/xH/5//cubk/4UyKujPKx/bzANxDeApHhkt/IJNO702zmNc2gPguUL
eqWagsSE9QBICVFjvjJii4wlc3mKZHwZhrlF0pgLJkjZPHXO41Jo32i+9xZNyShYnWjoxtxDjeBz
DXNYEzVNQ1SEJQMH1s8Wu4cuLIpkCl3qpEnFJq8Nyy5FbRwX7vVG6nZtftzgZHHgb79f+X1+g0LF
lJP3AEHLzcS5vhT0Ww5Z5uRhICgudgq3T1oacgO+SWkBRQxpiCi8ioZyoCRX0DkOIfjI8zExHHYk
OvZL36KivVVxjvODKcVMJBz/JSOZCwqa4tlYKI8SXFceZmzIKCgkCiAvq5GfdUBjaqwqMKVEhU4I
V+1X+qalVhr/1p0+usWdOYDBRr4rIID1MSTCeyFUI7mudN+QVeNvmdQQ4SFG543zzsLli8nw+ZwG
B5cAG3Ih+xI6LfqWnwAH1dI/jrY/iGsS6RYztHAoZXjmsATnxDzob3CsG1MU2A7NxgLdFZO0rk2i
8tMT5MfJ9LPoW3JRbJY36Af/yoypvg5GMyDWyvrMzDIkNqg0g3nBJrcy3wHqCYHRwXdMG4NZdvtU
11aeAm4sPubzZGl1kX8F71uJUWR64R8mcCLHe2PQNyQ314lZftqiqwfCWHNKDHl1nGVnqDyhkpX4
7NH5jza+wIFKNmDc/0ySAsp1w7GXhk0dTVMIePViS6RU8HDgZ1FD0v1BMuvSQGOI5Hs6+4+NB45s
C99508qbLDJns53aPaTcVeN3ay4aLH54/qfkCAsVjSVnxrz7pVM1iRT924fcSfCy+58VXGMEQziJ
YnE0d9oi9V9yEVoVhfBYjgb1vITBgehWR1uzOSZFevIAAUUaT9xgLMMrwDNnAPibzCfkp313prLR
xwHLbZC6zj+lV8X2+Iyglx7qj/ecYWZYaNvD1ZRlaw5DVjlDFSfTV2XWyre8XOAfQAsWSn3hgwRi
P+qHdxna9CwTraC6fqblCcvcSg6S0qeJE1tZ8PQo04Ft7O+x+aXuq0ha9JSG5LFXTXg2ofDNUaqw
u/mOxgn+3DwtIgzzHlwnAKF0p9hfg73TZEzOnDoW0rvLPU57gKIG31RXKMIxwrA/fSUvwH1WrKE/
8i0mjka+l2QuyOM8+T38bvFIIEaXz6uwaiJE+dsJIWPeI9cVl4VlhQmOAvH/HXh/Mn3/YHd7vdfw
ZRk+fjc77SNqvGkwDCMMDqFOmgmRw3M3au5aVPMhP3DuT3mCeQNom1D9YFwinmVDlqRz7M6gdQg8
894fiZIA5YByYfMerkfXXASvcwddXetCHJfJ/1D4Kz5bWzVJL5L/X3rEmvi4C3ZWVIap+AM28Wis
FdQ8thqaSbFNMSBpKGQHsfroERupbUaMnt35fniDdTf3ZA1PXgFTzmwnjZtdAAd2jFaDgZU7on7Y
CENHvflzC1hrD1cRH0UjBLCuyj51GlNQZhciLu0crK79qJeFbSoObLP8cLXNAwvgLDttmAF30qCb
k/LMG66rhlQ30oXT5XRxk3ohwvzL0jeP4hv3jQwUM0Eyi+92KX3RoyYQLngR+qLaqrvJgFu9/XxC
nkR2dWGZjBTeUcIdraORvvs2i+Bqcm0RDpMVT5IbiEPEUEmXxv/nPkzxu+0PNO7YXU+B8Tf/Ye9t
rvAE8LhhonkgzkkqxUg0oMoq6NZlFkMKgPsp2ai1qtTDoAldMdVZksxR6a9zfcueaiT54qAqd5QO
qoNXbgQr1+AYs6/ObzeIGpzzgPT1+e+/mOhn09pikXpFvQyG6cWs2ionjPbDbfVRU+SoazqF87Tg
0D6GuseGI1PyNoli0/FZ+UcVor8Wa4xK9cPpW/r+jmNRYA83YRXBJvT1q78phM/AQuodKrVnO+DW
99cwiHpI4BkTSR/mtXeVn6Oh90Ao0o+qa3BspQdiju9oCLQ+X/jZ3LT10TwYNewvFq1B1DKCurU6
bsL4128rj/ky2iz4gqrjp/drU2hH/iShvHUi0/c0Dpn8OpvS7IRHa7W5WC4cp/jQd4Jp32JeHc3e
menaqeV3lzMzPEIx1JogytQNrukNo6W+1LuQRXLTM1ze2Xv+9WcV1GzLL+Dv2GrU2++ERRf0YSjT
+dVwYS1ywsnaeCSqbjx6Ksbrxt9ztF/jUk7WIz9dUKVL1XsfolxGlPwNXg8QvDIyspObuO7T5X8C
ijF5Yy6gdk8iMBHWwIQOFvF1rQQMH1yAerk4zHJ4sWa9uW0YkcOxKijwYhCfNbusOxN6vReGlRV2
4+gqvs8Tq3tR+OeF1Rf/D67aoqgT4gpTqqvZg9Xdhe9VwtU6PyTvwWyk2E5T3DFbHMcukAUcs3Nb
cydykP7C3SNSc3LV8Bvx+WimHMJT0CdgcJoRcMujbYPUz4vJ+v0qktG8x/Ix7zZpekV7SJIO4z/K
zze0jd9T/nOQRw2Y6Q5W4hav/MspSMi/VUz6drSTDsGToZQyRipXgyOsV3WdUIUpty8GkPCHiuVY
l3xCUuuCuxM4KSpqjoRbganX02WgTgZ8ZYsg6qjP9sGFDZq31wMNJkDk9ztPG1ZXQp9XzvoWOCOJ
Cz5QjnywFpcvvxxgiNFxzXU9pNVNYCulmGiobgWBHInF5CoqrUQHFEhcO2sAr10qZFr5LsjjOIjJ
y9BGgVRXd+M62l45lMsP1oJ5EZWUvFfSu2dQB7pgMvMRXORE9mAgMe1FeHVvP92fLjj0Vki6nlmg
a4AQEe/B8mptsUqrNzYbmPUOUFvirZ70O30Tt2VuVLjj04eOKU11dlRrRqyP6qxN8jBx4PWFSJ1x
yHvIKqWXq7aQgLvTnui+7g/iy3zjphE8Qk3BEKWvYERs/3a020ELsGeXgciBxY0x7weuXSywROin
vVAQWfbj2o5gEMGEo18DHKPb16K2LZmpDNBaaFGRyHEfarY/eCmwAWmTh4KSwmCf7Oom9ZXodOYr
sbqzzmMvx3+h+BTxmGV5iPhz2SqGskvmTvvkoDGyptMDaWL15kmQRbbcsvN3F3qSvwm3VmtxQe0F
vr2vUynKx/HZEvHvZiuWhnZPf/GAc8AO+uVW++Nt9BYrMX2+LaGP1pv7ricIWhVk0Ljn48fhOZPf
uLNEuOHgkWDFp5/OjBAwDl1jfbellJVi4CCxUiez6Zm3CZptyAeZpkWWSg2B3FSGzCxQ6ZwSi6UK
awVnVklejfkDo8BySd+T5j52Pa4QoeM0/oAKa48n9edP51lD1kDNWZfXcFuSnHrED23/iXE1IulC
FHUQwp1x9xopLDqW34HC6EUTpAph0dN8Dl3OsA1+5Ii7Uyqp1tQ+PdlxlXE0GOKpTnU9I+e64Ktv
K0u3IVI5s/rYFcdGvXkCdTr06RwwZapdfgBvyAs0P+DGWWCw4Jem+nAaCu+b+0ZtcQAudUnh69XB
Hk3NQSbEV2Ddh1kmAiaqTZBlfN2Ra3vMVy1jloSBZ8XZNmrCHjCoXeh3HX/i4dlcFVjb6kfFVn8l
xSw4v+ntsA7p2YxfRCxGlVf87P8D7V1DxWTMSXAQYLlRN/14M+sVrod3kUG+a44k8T9K7pequUTj
LexqA6JqB2lgZq3NkAl1wkBpEA9/7fnYn7z1ny6cB/d9r16vPNXG1It5DTUbSp030hmhyAqNU8Q3
VPT53vZnKW5U0eIjLo+S1IodzHY73rZfbseYUw1vetAp/tS0wkZL4IytFo46nmBi1AxiWTtKp8R/
gSYgJHG/DZg6JhQGvGlI4ggVLB5/XaIV3E1+AGKJuRBXCfMDsaofso4H6Fn6ko4HTnwPmnAbK/f5
FwKTfNhyqhGRetkDxPBByzOJF5K0mcTHUqUaIQsq2TIynzaU2IjRyT21DHdlBDRl+QcSbH520FAe
3VECA5aCmcd0jYhWwhiPPMOHHMIqSq/BwF6GrrDtzbFgfZUJFhXjt8sM9/MYSdoWsACYHgnIJrR1
ceGHMWBt2VWkmePbVED0Sjn8lgjyibAXeCiMHidy46WI/AWoBin8NJ7FYkP/83pMW4q0/ddDQUv/
Pk63LE2zAdTCjU1caAjjkNnQXo08zPcHQ8eeuXA9nmEOlHeAtLlNG0VMef1l7x21x9Myw+kKRO3Y
m9vM1nYznkMxsz3X0vrwxH8ut5ejMuvWADT3vo6gY9KOB6an0jA+4S7qkogSK5k8FdytywdlEH4R
EKwBwQ7QGfvfnQkQlzb/c4aZjdSmDMLkcOg06pN4NyBcGzMARZzNB4n8AtKGojY624IQ0YczBCsE
D9MJOmxCEA1p1CdG7Xz9oel1N+AD8mrDY9EEtcdMURrxkT1qnSMof5Lz1kCSS2FoHb5kYnhTXkv2
TB/8e+RliX5Gn+A9vt173iyljJ8Xr2b/5Q9TMrVVeknvWUOSPbfFK5/gqoeLyb+cxAAE6ZA4VlHw
jG1BjlqeNiwPR28yc1ta71zq5paPXwz4VSzsGrqCW4Td45i+dlRpkiCWgkEBz+oxOlK7f7l46yv8
wO6r0JNeKY2Qw94lz466xlBI0MmJwur2U2YuphK7nwDoAo4x4ucdsIUzKcFO1Pz/LkD/F0S+gqxi
HlvNxB0XKJbdh2GlYhLV2Az34ZuM5UMZ2cBXmMmBkf8HGnmk4b/hh/3yc46XwD7OKRnPV4FtSTnK
sptn/NzZNHCMw+FQrlnQRV52pxO34EO60XgVyZmzDniv15DxW6g03wUpwYUTZKE432PZWNmynVaa
QP8AIJ6++tyGbBfPf8pjd0t5wnkegMhI0vZbc+ga9k3z5OKW0yrA0F4XZcvDRaSc7ooeRJOXejD9
39zApaszOPpE9G5JtzVdeM59cpKDCrO8V+F4XSVMrQMrSwU98Q6hosC8wXIpgT/HHBv+iu4s7EH7
YnPr5AQNQWt2j6ISwXtHBsoBxXc1ExexlQ86Rh8IA4FJBVXidRPqHVtsEyzDLZubpNY6gztZZPFe
61MVN1w+5ZFZl15gs/R9b+53HwONvhfzezSxWvR4CZeLWTZ4JqBM+mhk+PWOBXjSLITzCP79lQwJ
lijZurNJQpeD49bxXFfrjSDmZPSYKL2xngUm9CgRuIsm6aSRWXbWOfgRt5aTLJpBEz0kTUtmvDfC
Q4RGGRSggV731RM0YzL0SWyY3vdueIyLDvPRekRVmyqGxr3h/Zsc0PLuU8isJ6H13Huibc3TteFS
+nEt2MOp12yVIzfsUHU0qjREgWnlCLAgDfjI/2ym7Qe4PI1KoW1WK7Pib0jOQ/Eo9dBFd5myCUHr
c5GcZ7Kkl9ixwgYsg/58uqKVVe1L+5YpAAutZVj+YNjX29jadq91ZahyJDNtv3zj2GgmaHODMVO7
Jw3dqfch/dMupR7wP7zaO4/FvgWIY/ghsBNHKLx6UFsiVllbFHiatoPjuydndvrnEpmXAzJ/tvot
F252Pz3/cAgElL48fivRVssCmFzIWMhtJzK1JDQU7EIjtooDQlzKfqCbs4Hh9UqocijfNF+Wlvua
Bn98NmKwXuCuOo1lKqa0otrmtLb+jpy90jQEYBQgetDF9mnXh4MwnQdBZ8BPECjSssFcb8RBcOH2
zNzxCbLPmhakwiXGK7migTw9LxYnEZGGXPW4XV+cEtC+dFKwwt35kZTuuIQwKpXTrvKwZgEqv3hK
135SoS/K9SwWC181s0Ctm3PqPhL0mjYZK9lv1WCi4Ny5hG7ac8U0QYYv1xZzpCF8zdG0Fu33y2ev
2MlG2Ae31MMzRVMqEBM4yXCHNAIk8e1b/l8H6yARccttChps0PjUUa8XkD4GeTWjZzfbKkzWmwDQ
4CZPLiYeh/q59n0N9jaYR4dFW0Q91QQahvsebTRTWiA6zPg066SowPokvJiBigVkEXRzPFgc/1db
yW+JIbLqH/g5h2QM9iLGg9GN8RWL8DHVgvDQKa3r9OSwHQ3tFbX3ebg5BrH4/D1kIem2kOMarPcc
5rN9tUubG222iWrpktEpGxeoPG4kxiIgy1fV444OE5cqq8wM4zvk+4v7U2tX6DygZ5MzlYtqkK/p
gJKKfD470iB7rRNeHo2BUNgY6C0sCYQmL/HRyjoL/yUc87rlwiqXqqGrfEQT+ck2hUR/7AwzV9eM
mCCwl38mLv6bx4jfhD7vz3Ey3F4RZAIGPRcWAp8qP/FezoTJ1zZfeQfKTNZUcs/J/ljD0chrx9fL
XsJnSGBxsa3etOYgCZKYQ3nR0F+qotH5h+GhlkUFhyzzqoscbprr/4+SkwlCrT0WQgNavmTLp77b
DA6+VNtQolIB0i5Avq3xuC0PQAu1xAzSVe9QzcDUg+PLH6S6h6ky8aGeeZUUr0jqTlAIigidAOMy
BiceANCWOeNWymRDWXbnKfOpp9eMlKe/vM9slCFPRokOfzGp7qyaS3lSlLRQEoYDRi0bqe1vPAv+
vBpuotxjCcXNQMpRmrhriU6kBR8py0DLDhFyj5Kc5+Lsirmu0Vi3JXwHIWjMks4D+1/59Kpqd3jA
ZhR+Y7pioBCgSrGWEfsyC94EgnLJmkqLSKB9BsjyysSUqz5P3mBc9WhsL2BATRj8UBNheVm2zYX6
B0dNkTaM9znbjQ8zPqPnSier2CEkA5oyGz0us5kkX0SqV4YDvalEc8eTL6yyzdBkkpNd626FJeQi
7BdIm7UmLeKEH4Uyr6eIRXOJWbg5RiB1+7H6tBhXBz/+VeRo3RtMCmUK1GCEsvGN3lViTV/dXvm7
uYC5KC4D45W/QHDmSZPaGWgzGXLHccNi5je0g2mvHKUlCXENDczASZaM7w2ny1okT0GDbjQZvn40
TWkfsOhTphfe/BnUCAAiojPeQdS+j0WK11gGTzxzC7bncQZNvBTBfPL2YayBQ2VXqSmugRBNpEpU
S+ZMZ25RHQi+4rHUpSC/8sQSmZvEM2d/xymTIArIi9B/k0VPmFNxjxxMK1KrjGMVDCSQMrGqr8Tq
VsQDxV8pN6IVhPgdGgS23/RdIMhTs+BFCGFRfnDE75WNtXkJsajBMBIjoXbzQBBJV1o9FJvBwU+7
MjKo/PLIiu6RybOVhKX+TAUOd3dYavDlOBm4vq2kNKN6IgFWEVRhEGW8J7TFU+GXGQZp2P4JKsEm
qHVsZe32M8QIzbtN9ZH+Xqc7I9PhE30T4WxDK7SyuZYgetIrsWOXbU98zPulA0ZOPXREGPBB4sHn
KDOS5g3sYo6bqe+2FV5Yp1xuW38NrQctF+2BYgRFGSpsnfByIh8OjXG2X9fuUg+uSbDCBxMazekG
qAcWlqQoJxMMNw/6SoyeSQODB+cI6jwPKFyCYKi8AomS+MIPdyKLBQxAnZH423hFgzu3JtIvlyqK
YxunN+UM0PwafMIDuEcSPzpMCColm7DdV+B+Mzxg2EzuGetR+xdB3WKXx1idMJSNYFQMB+zL0Z6T
ZGcmaYKzs+4neQkIrOWtZAHdazXf5XEPS++6l4yq/oo5OHoQqng0RgHWAiy8e8Ax7HlEX388c7+t
lYcdSqZa3+p/jPYUezUUHcBezV6TjbXQgEMAl0WPAHo3yqI6R215QQHYSjyJHaRPpLbvK8TQl/nk
chgx91xjJSY7I9DJZ0IxEEBytH+RhWT1OQh6f2wxZ3rXR5bTAPvPuYNxPF7wJE2MxDx8qNFUp1lr
4toDulFU8KbOfi39bja6m8xAhcvEQXqAbAXd+VgJtex3P0IPF1BmQ4z/XobOdLaJYW8qOU08LB5U
OtdtL7SUcPv10e5ugZ9l/xK+Bn6QEhg0fUL46jE0DPgMzpVibBFFlZdpvxbc6TfDIAppEhohQC+W
dpupKXYdbE4/bJh/tTUWd4vD3P785y7LXBEAtn8MWIsFMl5r5nDoXiStqNO8rbaJ9lD/lE+r/Pdd
oazypaNAYbLFAlw4J8zFwnFN2nZ+1tcz2vDVQ9KFWUzwJFe+F0IoIzLTFw2uu5VqZJ4GH+cXoKop
+ti4Rs9ACRsQP5a83LzCEEns2YTnp3yqNKVZkaSSfpf2SYqsC+ADITLdaBGY0UcUbGRXXTB42H4G
D5F+Jp/v9ZBVH27IusRv7BzshfbH36MofHgT184lFVFiG7YjfCT3zPE11uqllVVLWrYXDO1YzAr3
YM+QNneIzzi9ljm/OhbVGO/oqN1yqYFWu9ER8+4/rvwUQ13gWxiuDvmwMrarDAFmVwrlfx9TN7zC
WjhwTd8HX1EVmOaq5QoG9UcSU+kx557SpxPiGEvezAigAUMjUXzL2t2yqwGzAWq1QDGzqdBNwlu4
fNDS8eC1I2JzPljUvcbJ5aMLWuXBPoeeimxiQ5FbbFCt1IhKjWCdMyJqPXZ7UONhE4Pe0m1+pfID
SB77994KdRwipHhm+Kr0y1j7NW5rRG6zM4QUZnsnzCRjScp2S8PrL+N1l4fjrCFfz0XpPn2rnfYO
qCw8s8x5wphdbSNDZcsbkIWGbwrbyugdAloL5kpMyARG8BVIg4xjer0e3AxqKtQnvVdgh5LhYxx0
dV8rZTU9msZ8W4cwbmsoJTu1rw2wXgBiMiDp4OdQBuqiImx2oBCUOKvsFgrrNxUPre0N/NoBlGDy
ZDdzF5Qy144nP1aq02NLCo3WulMMaZvfuBb/8PRkjuhv9yHDRHllzlCJQ1S2xx+CoF8mAeiJ1dzs
uK9duB9BoAZ6ubPlr/tGjTEteQhz/cQ975fK7O5F/9J1YGpbpr+CNtLzBfrTADN0vN4Fag2pFUNB
/dV005hMCwmJWUPufyiJ+FJtWnlQ+yZwls7wZGZf/IrkPgnbAGVRe+2AXixCLUDnmNihdXfeFBBH
HDAHW9KINN+/b2uQjh2c/JBjW2yx1ttFg5IlRd2G3dP+CVA7GA+AAvz9vMinoYWGO6shA0NSRvAf
VRuHhgJyALxtNKTwqjSAbDgicXHuJ0VaoOf1Coen8hkBRv2N9q0n3n9Ei1DwOOSYYFkZg4uNCJ/e
xKg8E9ibjuaa+lsuV5hZAM0MRgpAR3YVzbeoao3TwIA59JAxD3Mm1bFrBeAQCMOT6fkV4qe8xOqi
YF2cLsh90RxI6WV1/72zwVZ0PuplgOFCY5UYraysQ+CTLNHEVtZa3KkkZOMlSVHYjZq/N75h17ix
Z+IxSUiYxIe9mAIepB6BOYhsg5/XCefzJbDW9At4+W5iQWnEpmsSWmwEOr9n9WHiPuux7DrHjynx
/6Y3gCsfl1hdT4aI1olJ70o7+MntrnOPpCd5Lyx+D8hFbD/IUw/3e8ZuhNUXq1x9xZo51he9Bv/k
XeWm0xE8fptln9K/XURkyvOxY9ENQGoDdzs72XXu7Atzg6Xt/t+GPpiU+n/gUOUIIiA5nrn/t8Wk
MjzteBSu+UFVczbnOw2v2O4uMPQXBbjpqune5kt32rwns2UCifMY7pxkpy3X2Y8GS6lkqmDMEEkn
pZz8m1KCnB/tp15eIj1RiinBzRzcg+dwVcvh872NfWVVF/r+rlYjGtx2bHiX/hCXoqF+tn6TWUqI
tZpfjrIeiHWan4SD8bZ8dVkwLpOY8wrcpRYvtX4HiB0bx8X7cXYq88Vry5eAEm2UfPp+VJUWLZ7G
VzyMvuJggRPBoFQ/mjOpMRAvFLYtjfVXpFrMdOk2ZQMawUFqbo1Tcm1UBLtPkp3Mpe1sApmD9jJ4
9uFPgt/cz07lM+oWqvNSHtbIY3vCGOawurduHBuaQUSLRFKbsybCifNZUTkD0dIvnwjzJXEjQZSR
1XSN64FgB3bLw4KYkH5P7s15zSTrlUe6GpwxFKdG6e9gJIhSkl4nygQ2OnFcsBrfgDVZk1+EVYBF
Ug0F8Rvt9NqdY/g2F8LNunIgd+tOoevVyCit2sGjtnV7vSvaOpHXAL1axGQgC1sRHDd53tptw5e6
TssXaYcKzengpSkNTLJWuc9pbRXjwxSg/EgcaEj9KXNPjgQjEODrSXVemfO4w3oGTvLqn9dxC5dk
+KxFT2mNhSL+BB+cPTA048irjrtue5hlvTcvjyPYzcekeUNEdGUV3sS8vT4dNvOoln/4sn1/Kjse
ZxliATp5uIOH9H9cw9bzJgPBWWMbz7Cvb2INkIceK7//njhLMl+5KjJ9HJgxTRu5nuvXh44t40jp
6TXNYuRr1Pd6NIAkJA1E3qrWS62hFHCxR22LW4hswT/tlQaFloYWy1c6cxKd161v7ySns46ucSlr
lsz6mHy+X70lOzzvbgyBT6GKh2BlAT0FUs5HdoNPJDsgu5zIQU9548jf3UoxWU69cdIj1a2+sMGp
q3Krlf5e4qeZIZ9d4jNtJ1xMjNxuezOL+jjlmBdZeQP+QbwgFuG3USjec4fV5KNs+UWWpQS+6wXL
IZ8CUIaw76Wxa+ohPj5Oc0mJySNUK8+0D8nFpaiEyYAPm4cF5lr1cM2EjRGRpwfXxY+dRVqfm8hC
yYjAqkufBp9oiRlg+c7Az79NZq3nIy121i5ewLUBv/WarkHgu/soNmbI7rvS4/xYg9ztz37aQI+M
jMKF6Ch7LJnSf8pVXMsTIE4J0YJy+F6qqyJWqSEDLsvT4eB2fZmITsBBgWjQYNvUMj884SMScGKA
zBIA88Ws6e2zF94WoT/G8V2yzHFnpGHY20ifSVPa/yXTG1Ljn0RrkMcfSN5zrSe42tJC3YkdrVnI
fO/jYO3AeX82SlamzVrtgzCV6HJEsBocoK+zw/VMdT5Bg0R9dFqZYk9vpB6Hx3AdHD9cWigIE35B
MTxe0tnlt6f7IzDz+ItJDq+mpYHpSMiXA9deAystT77my2KHEQqqcAj7/TZJzt4RTaogddVMhYRD
mBU/tbcOAjJ5ZvMrfB4xvj+h6l/QJkZ5NOyJ+6McXtCU9DfWRj6y7nbadI/5t06cDIuWwy6JMT5C
qysSpXm1J0I7/YHgqvd6s6fTBGaA+2Qzy3GOqN9jc6vJ/ToNkipW9W81mK0HySAf3CKJw9EHswrU
qWSWay2DTyBHIVC/KTkpRRdXfiLvSuoWWm/6kJiuRnaVi2CbLCFbskihuVoBj+YK32xeTRLpmhfQ
NIDB207grRO+38mxXAVJcP2TcsO7xuXKssa3cXQ2vpN9ZeOVYNJ5vS0TRqE06+qEIQlGN3IKyqHY
/MyYNQUEcJuRB3o4n890WslnKQdiuPrkGK/Dxknltk4MgGLZM8BacIMchy7G1AS9A8DxL8qUFHfo
7PG0lUkwA0ZnYXykqGsL9B1TXc20cJy+b8ZXiq0qWJzJmkOotI1P/nSEoFr4pXq8E54etZFJdb1O
XhCuZLi5dcLrbVg30mWvgtxIlW79pNB0rTKha6BYoki81XWchNwnGL74kWceApm5dwiSZgg8Psjs
4sNxSBMqe2uMLu7GC8w555/Jb9ofBqw4CBNU7XNnllBGqNgQWQfUqzbZiyvbGrIhq9ZwNJxRO6bF
QcjEEgg8YEMjzxlphy/9cEQGLo8ei5jvkjHk1zb4sPKa0KvpTNfgppongjCikVZXUpzN6q6MjsB+
0DC2cycZ2Tpy55uqCCef9vKvVOvo4xScExvpM9aGQX74xpnXtm2dHVaaHwJinGscYdSCzBmzVnVI
ZJwF82hXw+DkONbu5n6N9cVYEsiOkhigfysxcilzyVEqwjrFGLXFE4A0QYixO5Hxml0MRCWUNKGY
cmkbKueCvJwJSaoaXtq4b4g/qyzDMb3oeGneOGTq8dp0sZATmeShJaCfly5I29lQoLe5VhlItIIx
rkJRNnGhM6AbdthA8czGTkMtpktNzobN5r9dzKilCbkv2Q9aYiQXlGvKQFuE5ca/kYeOWRWeRINd
P9vYanV+Lm4pr3lv+KdaUPhxLfjaBb0S75FWimQUovLRDvyfS7xS2HJ1GZG58WhR7X8PZ9rUF3LI
UMD3ZATHhSJSPffNXmpX1zwQ5A4mfYiOSniPeBqQRL0Fv01c35RkzL/WL8nGSmlzGhhpRLLwXCS7
jhIr2tW1ImPPXZHuc3rkyJuT4izJHXpCWAyKDRxov0M+dsKZawE16DXuuy+4PSpQmETOI0eAV+NO
SeXiyA22ReRbqQwXm1gGJMDsz+EAIcsEiAUuEjOIT3V12kqLBSwKBWyK1ZC+a6g/JS2YV4oKzN3M
rXbYOW83Jpqq5NgitHmnFgBh2W5lE+IhMQ3uo4YkW6/LyquUQgH50siDMfOO/GJoo0n5bXgLPRA/
ewkec7pgnZ1JwmJMwzHH0JLoVOhiD9bi8Me+0ZglmdHlC2u/y0xC4EItTfxA8okOrE7uId7VCOB/
d+3zVsfrqCoWX4fuMCZN73ScF01cL7usMjfh1Uc6pBDkgDN80lHPVEtf1FZZ7HSk8nJWTbTF7u/y
5vFWyYp8a+h92WxP8y5DQPk/K8VUSDKA5eQ/GnkbsoQfxJlN4MW30Gge9uuOvdgGn5yscbycVLv5
kyZCTt4ARGJTQRcH5P3QIsc5pmHnW/6I70vuliBNdHeKFjMW1yZIy+D3dXLEeL3b5fnqLDX+RpM8
65NHW5e+H8sSAem6Bj028Rn4EJA71b41FNDy4Iq9oTLuHLkWQvYdL4PRtBUwKQI7khRIRmETBAT8
T8BwwMsLOoyJyKTkgx0awrzurbu3K9Sgmh4SdkFyAz10nZlap4+iwMOgtRXe9CY2FsWJ9wGNDXZm
mwYOA3zx0GTqqNrZ5ZgdDkG04VqCUitsxO5kSjK7b12FT8Bn7HFiqRwLFcDui0UiddHxGzWknb5L
jGwDajX+67l7h1GfA3Eqr9dZu8axxfe+dDCo0GQtOlmz9JCzzqribuNlHiGToWlIy+ZkXVKlzEPG
HXFoZLhQG3+LUzwpu05eMoIYxmVyeCXnutPw4zU2R1b3iIvg+bxeLx9DgPIl4ImhtW8gl0z8+t4P
yaNJL3mxS6ffY9IVt0OBM7jEj4gpYgqjngnmANdXVFa5ZgDC10/P51s7XYMFKyEytray4EyoWFdP
DbvNp++Me7ZY8TC+SOYnOyZzRRFc3rkC4/ZwSLxgVjSwIXK+k7bkMQv8CVPZvumJqmP1GPEz05+V
ql0ku/RluMQf6v8TNcM7umDF0EVfxmMvdr2gVVIoaHW7fqwUuzS01iRQgbBp6JaxXhQw/TcFtp4S
V6XumZpGYjPngIhlC2NBy2AX7uKncj1TY4arBsej4cnwy/rfEKZ8W+NGHbNq+xEWgC58/oRowQDD
2TOX9EqsSKCGfQwp+OH8E6jrCqA7E/6IeWjKGomzSeGN8wBTeV4xC0gldNNqegjvvr3mWJGKoRDS
nv+Nk5cRKpP4qAUQTBl2SAqQPRxrzZr6WmrS+k62HfdrUQqa83Z1AcrC6NhS8OnSqyz2n1WlveBa
qBkXZ7XXM+S/bI2RO9vMJBIDoBIsKYl5RHMJzsA9cO1QnE5o246UgsGEQ1Nv8Lu5PqGOzYhywcp0
A+JjhiWuHtZ7YH7hW2WqQhmYnXlUddqG+5PVOZlUuIWb4nebEJC5/hnMWrV0z6Qt3lTeJPtv2B4u
WjPV3DEmCtHeETtk0YQRggW8rNyddNIEbilvyrMpP5lp/V4tHdBaG95LgeeyzbvnM1Hanrw/IKIS
MkbfP4WuXkh0S8qZsOz+LIt8LCZDj+7ZwC1ktLNxCRiqZJkX89ldPxlwC/1HGO1Oem7J6MOSjlFI
xy5kRrPCzu8KJZXVAY1eth+/2kEdPHswZvY6g2qMk3AuDnT0cgj14Jvy0pbywF1fYzD/0YgaoO1P
hHbICIywiNUYmhgGGnM7OWsRZiiF5KGLR+ngr5QuA+ziiJ2IFPyKTWKgfyF0IOx3VqFABidTJMQt
iUcWyJm1HYyikB46WYTpVVS3mGdoMXuanxNAo8i/inF1Rrzx5jRGTbtbZ/ht0eOjajmVqa1k1nND
z/tJTb5Mp8yYiVw+nlZlEdlwWejfS5kGKzsoohIn3xF3bbnvtMsft822mnl4nHF7RxQCg4zXYloz
0WnFhkFVSckGynDxQCXhZdEAb5l24zPw3UH04yytkQPpj1/zSokubRlgODWEeY1uig6A5OuXOG5A
p+TMkFiun1v0P4KKvGeQMMOVNNGKl0gNhdrD1kTT9uhYxXa/LF/z/Ss/PYVpRd4S1DG4h72FVvBK
ujpHj3RdNxURlQJo7nZhRTeW2mqOgHZHoD8GkoASSSHBjhfRX88J80+OzGyQFeH+W06f7NAxXj4E
pHXpq/GREpV62Ziy69G2OigJ6gh+eERs8V//fRK7Lh30Zig77d/7MLqp7s/p3zIhT0hmq3X1aDtq
dn07dmYBJ+TJ0NRMCdFtd/7hxHKm2vlr86dZeGB3O6zGK+SovPIszgiOsTvy/9KZrLdv5FyEz5dH
uec8V+RSyuoEyKqIlm0jbstnbvfjkLEu+XUzibZftJPK54ltIoYDsgnzHQF2zdOfXddGg04RiQR0
jAJ0uFb9a15xoKbRoOzL3aRHW9Hry0UqRl03hlfRBI/aHtTl9cVjwkw6Wx+SMl/Zjpky8d2NkbFE
moz/z/uptDEpuLWwJ1pR9A1zqfHzufw9ZOTaeqd2CnSGqmW6WulyvbNAlDqGK7C6TBmb03Jl1WzB
9TcssEWpZd1zujDeUOM6gAXHInE1AXtqReIFcWR2w5eUWyFOwWNOykDg72TqKo9ITO1WekW5RS+c
Lmg8YjAjZbKQnTc2TvGF0Bmq4i51aSvyczx7wq1zhazCswGBgNwzYb8dWkBE/U1geeC99TJ6Wp85
295xwCk7hwpxH4O+CtocSJFxMM4rvYgWetWSP9+lJMlBoke0UbmMuc8c4H6j7kvNDudnsxJU6tj5
OtYkkPMEgjNIHVJ9ssuj43Grk7Lw+bb7a44CP3uyr4/s5KyGEaJi7Nny81lfPPePkJCHvww//yr0
e6ZH/iPyVOeaQFw7t60KFGYp2uNYfARVIgzWANmKFpZhVuc/6mFO/uM2JzEedO9ckRYJvp0FJp3+
XDd6eM00ZVPGMVAfS6DO3OwVFOZN16gfVjLT5Ct7Xo9L1e2Re1kxmswHj0uY24Eg/L3kDOYA2ORJ
9bGFuJw4JpEWOFUKZYLgwYDjYCk9TQeWP4LDt3lr+10R6Dw8Jk/qQHATDUNoUPPVaYcjQvjFjMJe
6uYjsIetdK5zhksm+rHgu2ZespGXB4NtA5ja8VGIb0rq/dMh7pwLu8oewdsspfTdMlBPxHDWbiUk
ptrQ5bUsMK366PM91WgwZtFopsEkBFUDjCtFnzAM6CJL4rJ8b2wPWKwjJlUnRti1phXLBMNVriYS
HVQy4FfD1iC2qznO69u2NBb5QnvnxjRV9TgEutn+18592mvft2lqt69s4a6SW1rP8S/qrEmTwvKG
U/RM1WngVfHxJVGF6fPLyS4KlGkJODpCX9OZXU2p89q8ObtfRhh2VlikSXfx0JgQqr/xTkqQvAc6
TEeFFao2EuqdZuymNpaXPPnnUNK/k81hhiWDLcs4ZkScSh/x6u2GPcchfL+D5xJgYY+raKhboVre
etCYyZuf+WzDITAmmzhpEr33ISacHn5ZZIf+IfKzJMlFQDc16xetklyBJvM/6QpY7qFKcJHa4za4
31hFrJ/3KIrNooAN+FdyaEkxmzBziLccJ/cEGzd00iJoNmMOyH+9YzO0dBkAYr34BwTjH0MUtvm3
IbSkiek20unk92dsg2DizD+XGmGs3nmDGD+AEq42qwfW1wwmKzt2h+yu75PrF4lnwmOjCPPoi3OM
JPZcwTPxCqtJff3MxuwoZMCsFjgBEkn/BPJQaAA9C9f7gH3nmpobjDB0cPna6vw+ZMWB1tBKV/lg
dF/VMkNXQ0Wd1+id4UHJdxs0/02JnBROzN6HP9Xpg7J6OR0zLTr/xDvx6iNheffJDULzf0qpa7fA
7LNTEm1Vc1EUFshBC2JHvHDOQek3Ocd5DSa3dmafoNnCBvAuCieI1IQ3+A0DS3mdi7JWQFdZgLi3
DOXRkOjOBXEGD/XULAzb8b8jCr3Lhz8TQCfEsptSMZ6VytIksEQO/FC3VsV0UIw+ssD+6B9FlR1B
W6PzHKS+gsVW0/KMuUfeE12whWAb9LV5RAurLi+zQ0WCc+OEEO4CTocHf46oCWLhy2c9ygtq3q3m
Df/JWiqjjE5O7nj8OgWlbQR7ME22mRjKxNncO35IP2nHCqs64NSQTGqqx/fZvLjGIV7elDGmDtmH
X+GDjOGhMVeD0NLguOl1gdrt//0fh2RdQaB3J22Mw7kI/Jq/NzhqQjsEuHmIv+kFDieNT3ExUZB6
Gxpa9cRjdVeRde5X60JU9mo3jHNjN1DHZPnVXkWAU2zoj5HUVV6EB3lHiIN1gVmx9eIxMH+sKSL5
XGEYhVPdIMghMiB1OpHX7S/TSu2af5pf22+A+OI5pHZgwgputzTFDsFmCC1RXkANL0hatTSXjlcg
a2KJ6BMDM/waD+lIggVZCpeFNvgQ91IIf7JaGr1FnvmgVHQBE5wW1rO5c79mNKjrytx0li9ozIkX
q+OJCAZ6UJyncaQAvztJ6+rvLGbpbM648AoItzbYB7O0jaPKQw64W3yPySh+46Gxj8+/1SJmh0Qx
6lK2tMP0pvoU0zdmCKEedmfQQyhuthWsMqqR+VFZTqsIvCRXbliL53wV0f5hq5CsiX6ppTTeMTnf
mfFVF+0Zbf1n4VIi6PYFDHDGak9ECgyvQIVgTw3RZZUlJ5gH1+uvu2qDGFMkDgbshTQ8jRD85n7+
XWPe0W6psPU9GXU3mLdnd4a4vg/3Y2TjdsDCEjj8500WZsj4uALcpM7l+0mbfMP2Mh+6nEQrZ2IK
pndX1t4PugWNyDvPxsKeAZMmW1906w2jsO5s5xn4jKkmaCCffVAU1orQ11XPequhcsUkfGxbS+4k
2gbLL2xhLW8AVBtevL7MljyWrj26zMI/IeiIWNQH6eVuKjciWJhRnaJ5VCyxHI9rJoHjuJ4Bz9Ru
LCWmWK9VjW7IfflF5P0qsV1GyV5R+LsziIwDbev4/RQABCnfzk8QFcP91PeHQHPX15gUUTequH2E
W1dFbhBLn/bxSj5qvvMp4EztntVYPI7B81aUIcZIBvb+ZuPBtYBweMvWdCRIdMz6Vm6iECHadZnv
I5V6eDsm+GCrAoF0uBAy/kkaz1388zK49ZH7hy3sfKG/YDeG2By/In7Bd7EWZzgH8faxDI7bUoeZ
ARblb2tYGRmiAwHO/fY6NqfRcc6cUs/Y0DXFq1e/fBNPfDpwGpaF3YeKF0mWV8ZDGY/i+O/Xbj8y
0Ap0Am1C8vwKY+NTvlWnxfQvN2Pm3GJYKW/RCg4xZCLBpIGDHy7iNz++RyOXVsN9y3/svuChGUXa
+Hix8EkCYxYcwyi2YL5y1xbxEKpZGC30G5JeYSUd8r9kbVhx3nRH1mDNdo3KQZGT9zb18PRefFG6
i0/7ruTyBlW3t7zlQimlSUvbVIT4RPLLddFFL+6TjMct8q8yr8rtx0LCk+aSWSRWSbY5ynPlHCc6
1lV+k8OgFEwuFQtZqoQ5ZDYZu2VLwKOg6Jkbxeoa7tnMnHJpcGe8Wr3Ga2vn1YckZF1pCdYsj8T7
N2VeYtgeN311HNx+H8TP+S4dRZ0EU/JzPm1J23AtWAAVcFCbMmtTtDCII68rJIZKiQ35CIEaFoXD
wWbWPvsVNMME3KJP7jx4zp/NB87opeEU6TsSFNMvVFndFXUjalfFkLcsLQJZyfg/lmNVouzR1WYy
St7UeOk1SBrvbNs02TNbibHFdRD8z4Ydn/I97zUwyWmDTNsUbLYsl5CH0Qe0iQokSXhmMZFV/OvX
rKSLZtSj0rRoumtH/6b3lnUIvPzqhb2omcwfQvhdAIx4qW8rU6OCdGPpaQ8U8bGwtMQ98WZYpddB
vMYlJLUVJtFhTOI+oWAV8vfBtcDi2vD9aw1kdWRMC2RxEcyq6nqxc4YfPkjwzQPfLrE3zor3j6er
7/hfmXwEZd5RbCPenoggVHtGihverVTATZNc7mroesgbB2tNnqj9xNvSvnd+5zo/IMFwd1ScfoSC
nJ3ezB4mZgHI0N6x58UTVNyxa9STX4TkHmcn8c4wxPKV69/+PP4FO5ipbBCxkxe2wUoCfFyH10AR
VEeOGTsTbO81DEOLyWmfOiWc6oLASaY4twf+8lQbrkUa9UAsaeiNPKxeVabV33Yd9U9UB/SrKFK7
sQHaS67Bx205uRGF1wR+asGr1lQm0W6LoX2NdqQ2wh99px2w/UUHUFjZHcSxZM3EJ0z3MblTwD3T
6bqXeCFF0txDn+cARqbjxaWessNTpAbqY7bsLKUlxIpZpbVR95xVC5UibrCoYr/jP/vroNv/RF1g
LQ4+MnYLEs251djCc8AHdlc1HRRpZ79rOLfda6P91Jfr+bvYDUJaA2XVeMvGAvPkqrU5PQDvANHo
N9GGf3R+/xQBY7KRevY4TBQo9ed8zgYu6m9Y5qRPcDt+rQqb8OsIr9QbFeZkKu92w31bVLJnDLJh
0GByIbSKHBn6KpBI3KvXNShni+4+pquC0qwlaE5+jD9fZpJEmZOIhuHaVHkL+/qn6j+YTgZCUAZ/
lgQYZJ6GoCF5aFEOsLNMDQ8lsa5TWoebF8hJoBoEjhir9aYyFNgTCButqUweSYP1aNmq3eirtyPG
mHRpeIhkbZ33HS0r96zeAGlyrmQy77YTmZmsYrahbtZPi61ZFV54L8YXkrx1NGY0BY2nGOENxyh+
c+jMAzh/jKMQL0EhRSvnz4ZIst2oEGyRor7eGxVhKRkIdKJSKR+dEbExYhAwSZrJcS2r92wUOkXJ
2EyEXsHs5UIq4gRrsPtVc8Lem478h6+cfsubKte5SjXfH78dXfCnwq1FVyvvpiZBmi+cNqf0r7vc
TvXOIkZPSTihT+iCEu5nwDpdwwNdVs+zLXVrP5BbRzWScdwzw6Hr1HoUfMwwH6ZpmWVkBzE9rqMQ
oMBdFAMOGDMJFl1WixIH9wThKUgcEWeQzVzh4SZN+NRevDxOpQ+kqh9Xtq9xs77SyJE+zPu5lUCe
EqnJ55JFfyBy0UDx6lwlWtZB2n9/fXKcX2K8GNba81soPrK5c1locLnrpFpFjcFt14W/dks8+7NK
wMx28NpLkpxqUvvTsHF3y/q6dgpCU7jk0NXtMLgm8gPygM6Y+BixogfnvszzhM0PuMiL2TQM/Phz
FbKFtgsj8/rHKXWARrPUZgkiQOo3JEgnX3CBb3LWBNooGWEsQxm8aNN4bJcvNkkn9Mxy7/zRthHZ
j70AdfTOA2ncQCdg8MvnWniqbMawSIWinyevG1gNUY7yMLeu1KVKz4QtFHGRLKwj20OueD+VGqML
MslmBgA8dnpdz0B/V9YCSXeAs0M2bdaGV7Gp6KWMe1KsjXvEfGuHjiKL/wcQ9wtyVaS7DRLk7ZyQ
YpCrIbg/E0HVZ18TS1xh6EL7hgA1DuBbOmR58DsfCep2ZXCjDGH8CuP47uXd0DrPphxkZksgs+IR
688FPuRRBCQzfqAlM8xaTZy7GCgNzbN6mFNOFg69XeKvP4CK4WhkvmqvDF9QO8Q4pQndF60Rogrp
vGVaNQtZXCS+xfI16DndnWZKTmylqKcTvYVeKNIusmKRjxMOPNZbjhhmTaJQeTpoCunGaYSue6D6
eAqfZVXTtiYEuGOJSUNAEGC+zuZbOh74DPjMEgaqW6xeau4XDBX/Q+mHAcqzDaeedp0e1UuU2Uu0
8TQmhb4iqAKZrKW9j1QbPka4TgKukKAHG4xNcnr2WK9JV9yh+H/pC/LiVV/M3iRYttOmHLqlzNA0
lRiSyeaNGQfPy/t44G2hdFvTTXmKGuewAR5D8stpeGTBb+oNrfJAKgqDvmJumUH7Rst5/2gflB7u
C5DYTyO+RyICX5foUlg1eIYuKVD+191oEy2/ZHyFc7bV+kUxg7MUDJIcqbxyLxB/SDl3My/ZHNLH
fTJSjFl0bEpqgzK0yeGbKto62cAQFxSPZNTnTVR2YO6n5T4u8BkFirlvOvej3zI+frteaFRZsfxI
R3UT8r8RJYb7oE/grqZTC+yujwqiXTz8ZPduMgoMgL5AAMzwIvMAo+sUwpQ6JqLoOlyhV8XgrtLU
zMlVDEtD+0kDU+2c8mD4R2OUpOsO6jxeBtC2vWxTnlnv/A/dmriSX6mc4FdrRILGjT8d/tvRLmb8
Ea4lRfxJBPqCMPseIhhVpnBnd6Qf56ZGi/gdFMx89y5+Em4lDdR4fKJjXZh+2z9GAhnzI4CUA+5n
ShHLSIvNYFV9NzZAf20yRTq9ChhyNHBt8hs3I5g0Hlg1c8nGhjreizJ2hoH0AaIH/4YiP+5zL9R2
mI5wNetMHStmC6s8ZkvhjqrtXCw1XLV5Kmxp5HHbNiyy+KaitA8Drtgj20z2glFkOXwLUSxvrWF1
gMw9Bm6q90rrOq/Nt2AnSQz+aAdE19moUp65pqg1h+1ZDDw80WNk5wRkGekNGkpejU/tNEN6r3aP
gKKjtpMdluS3MUrxge9PHRisMnhAnNM3wvPcl+esEQYwSaeq+yz+mZX1m2VltqefyL6CY5+6u1De
084fTXZWwY8SJubFpEIZVx3pGJthCRxVhBQZD2dVi+8jxrgxPHbnK+O1GxxYeqkNWH5ygstCkoZA
QE+xAI36/+6aHXzXXye8v/qdgrRvulSqDLaU/rQr/yvyVQ7HchlYrzuMqpcZoL1Ep44GBK5ygaK7
qqjA2xlWx8UcmgTleGe8aB8S1TwtOBZpF56AyAOiYsxr45j5uN1j9KNwkv/QTrSk905bwIP+LP8r
mBQ9czmUmUDl/dPBRf8tghf652f+OkW8phazEfd1TrFWKB/FwVMZ0DAU0HrgZFOYH5s/2r5bHLDD
JW/1U/5birlhghUQnM74HxaDI59l/l0vihradjmZ0DbNTYZZ3kE8SFZvSmDInSPvBVMq9BCkKFlS
VYOqeoY4Q4aQkBeGzPrNfmkAS/Yb+47MuyXPqH8eTE/Af/43HLvbWP+YgWtAz6Psy5iewL6OZcQo
hk1Ao8zNL1NkB/LkEZUJ/pwRPr/aTqd2AWEbnpJElBSmnU3dbEnJ17/8q1YEV0QS++q+cs+JeX4v
S+aKUKfLNG78B8chZal+YYg7L+HviwQl7GyMyQFFl8utWEIg2EDwL3t7aZfDXBZYHT0BtQ+6F98h
r2/d8/j7PZX6OZ8BCpF0Q3EQ2ME4tqxquWHuelZ9wp2iUPRaPoD3Q045hBopMhC0rmiX9N3kpzvK
0u+GY5RqSLNpzZVuowkQVpYVyGFabbGJGWtpso8LMh9Hfm/LQq6C5NX9OU5PSUSlbZL9pQ/M9uac
cyW9yqlqKjhmVvkFgWyCjnSMo3DpOXrHBuDcMJcOkhhCs20cj2/GAgRXwHOAAySJjtu8mOYmWyT8
L3NLPjJUnsRHRqQsqXDbTLEl09t4+XO5mLtZMyymmOrY4/+iJ3PTycSrjojgHElY5YCphJUYLHTQ
frLd4Km54C4LmBEaoB5dhCDgs2+lhTItyfhzeoQ7WmEQgDxezKiVa+9otHRXfqfTf13lLIqE6n49
+tZtu0/zeAJNpGGlZoChVQMaa4di4bJ4cSFAkNNje1uf/GmS6+kUfo/8f9gHo4WFcPjoDhdDzjtv
mMtRtw81vgX09/6p8gUh5mo3NS4loiOrFi7DGGsuhZeJYJFviUnq3SQewhQLWDk0JxQilIeGXJF1
wWXmEeUD7tIzmdFVnsPPr/STx+/O82HL3zI26/ptaIhSOEl6lBThG35KRAAl/31RTnPsQy3qAcOk
GK2cpewVYXMKz9TeVfADglC4/adZUB5fyybMa8aj6SmRCEjxi0qvkdnlEhNL0n0hG0aNBmmUMMcW
5X5cFZvpOpJjgoomOw/uQvwS5SV8rJd7+IHanLOTLbU4rUMnLSTkBKXkY7agmbljJJSE30iI/UYj
hrXN+sYfXTi7XISzRaEFqjfAebT0rYnX2d3mpfbTYjUuHew4e9hErbBtttHNqgATHg3jh6p6VwDv
I3bwuFf0YXSg4gxJ7tSlxZNCevb/PlcEt2T/85VC2SAnIUOUnJa4jF7UrVydQlIlG7aDha+vkiXJ
J4Sot1uTHlxmF7IbnPQ7NgcYI2RSBJ0DodDIhlckasycY9QJvKnHRtAvtAw8iAUmdfIvBDHPKVIx
NHj6ISd1NOT6944PcS1lxfJv5r/lGr9lojmgEiaC9Grww503OkT4SvR2M/3k4+uJh4kcAeNebaQS
1igRLf4ivMaWxntzPOfObcY9g5sXST9eIDdwNI72GzrN2eIxylxRu4y5AsyxoeeHg2mZv6EOWt3u
3h0oq9kdUCpsfNKWyvafbuM248ZmRdjG7jsBN+NmQ9cs5VEM0xCR8UuSPVS0qEKuXa279Fb6TwXZ
Yp3IdIxcb6wFd5fEs+L1qi5LUJJCNuaYWs78eptn2bi9lxrdbU/lSiFrf5TPAFA2vrrCsFF/i4Kd
sRXXnuYAmxdN5tp8MyuUybig13cew/0ypD5tIa3A1VKP/OrzzVXf2/ABTeuJ/FkRW7Cn94ElCk/R
Ieksv5LUyv29CkDlL6QnS93CIWV+dB0hUeWhP26d8UeO5nxtfeDDGL8cEV5uMWcEFhG/aHdxxblI
XrJiNDBqcpm3bFRpycIKdXJaOQ8fty6JdHJ193VLIpnjQn3VJSIsmF13FOLPkxwYXgZ1E6mIJ+VL
l4qSZ5E0lWfXl39sN5zWuKRWpVHzXI3hj4owoO029TxO1ohaRgnoh/sRywnGD0jjTjveVdyDDY1a
gI1zImlu3Q9eounIP9tx8/OFGzt6R7DTbxF6WxMwynIpNEzform8IZr4EO6pQHNJy7Mb7YO4qbAB
JYLdXPJCFyyRmEC/vA6fsFbfGTRKgWtbSfWK8bB5CZ0zygSynuO9nBaArUHDtP6+OofAJNyE4uIN
5wiwj5hOXL2XvD8E8lV7sZCaCAN9m5YpyGajzvUbrbW64U3gzKoqHBKERJrjk9gP8LrvthOUcVks
EJjTtPZ8zA5tGMvScxyB3TrHjaUOUtXnWeATThnDirfhE98PXB5SDAE0u9jHXAmdMTsbfkIfC5ML
L/NpLZ+Qe//ENZh4v0xJ2Alttj1dQvL7LyLWMKW4PISzDp4As8RfTlcU4k1YjLEYDkSC/JoYgYY2
TI7tAY6PZYeD2TAvg7oWa45jBwkHYF6nSb9M7nPZncHUZhNwtHsRoe4HUno41mIh8Y4KVdItWd6G
KIf/Bdg2neFzCxahfBte4c0gt3q+HKexQ17M50TQS9FXC1N/Eq3mcyyoGDPF3nKKObgvHgtXgpWG
swptrGYMb+wcsb8rSfKHRhEYsXIBOXM5+jMRBLH1ONHXYD7cENBAu1/86Z9Vt5KsvNFxaCVJsj3I
GapCdXrg7AhnG8ot6QXkrY1qDUvC06Czyg0626+9Klz8tIZy6ngPls7BBnEFD3cN2lpkIxh8pf0h
pnn0Faxmm0SJa/HigwqRdVt0jLzn/E4kj4E6ovuXFuNN3fQOU19+VuBSdOa5ai7ll+hBhz+6/Pbj
d5CP1rI01pcpYP7NMHsOOghMzBN6ffdZt3+BckYKbmnAGZa/IdTmLx3laBGzBPuwVzsuo4N4+/0r
+3IfjCDcEwOphFLJIvAbCQLM/JIWzKBE2fwOci0dS78XtKrhSyDPX/BqEC9FxXjr5MI1lRNcOf+L
kwhjOaqWHJMmXWnx+m337JaH+yqQsX6YPKRd3Z09bUZ2ElBD3B7PVLRheGSAQcRWT/3q3v4TuD8U
H5foaLEH/m6Si9J531+eYY6lIyrBpXrroCyiDh6JHv1j2XYgW15wdbV7U/uGcM7lxMbR1aWOd7Df
Pwk1TuIGGzoToKtdJ9td6a2YRQjItF4mgDVDgdlECFIqU70K7JcKlIfQzDG7r4UIvvQ0A0w6G/vO
islCvZ0bFqibfa6V0mn0wgaEyjtIYlMRGWM/AfJUA4ApRju1WbXiEPO4omfuFg33afzkg3tTY8XK
cj+2VLnDzs7HrAGZkLP8G2rIV4+eMwPpetyBk8p/Fg39pf0A2B28Y2+cr+VCOzKKdFTbfcxj9Xah
yS/wNS3jEJmoElx+V7l2+bdYN7LiI3mLtKw9qvIDBzYpYI1QsvZFnKJ16WoTtOmapEWyaJ1NikpG
hO9uMRpNpuVJCmP13683apYCri46DPt9Zu/3EXKq0WUnWfRarQps57qDM0E1deT2S5Hnq+5uXh0E
JeeEBwTMKg4j78jPd4aQqvzjXc2oizc/0xezoOKtHdNt2jRHHWmbkDOiUUG5eUZ5o19PtCtb21w4
znuXu5oEj/pXHmVwWwVYur/AtCSDxQy4HjKLlVEIQqwK+L9qTbc1+/K7WQztHIzL5na770w24qpp
8myTcTyF3gaLORLlIyiRAfnHoSJ3O9yHCFiFQp3uxNPCmVdj1ZHI2mrIpCqP/S0/WmlsJzgRB9hD
x8iJyy9LIX6v/GxipRSlZW+vaTLOpDBuldFjptGjeXbnOyO4fSooz1jzA9ZjDN0qDLSpqB25jvCB
ba1IgMNEaWd1iwDD/qCAf9DsZAx8M5RVJUKac/F5nVMD5LOXpqmixulE9zcEHMHiQJBa6cCnnatX
n1xghTZRcoFeUlAtbi5Sldi7l2mF2XOQmPlqGFV28TJSvh8iSchzK1u/rpz3WJpJzSPHBdlReIua
wP2sLc7ATKSuZ65D7MptHFMYF+Al9a9XQkuNrjBlNNUh0L5p1CXUk/sMHuh/8V/T56jpNvsgZq84
iY25nlgkHB2bJQhM7+FCndBv3Z3YfsVDocc1IT37TTdyFq+E9tX+AiDQgmwDawA2jNdLcPdLwNH9
2//ePW53lEHdQEqukJn5kfOwjjFCseN20KCF68QqEahB6cCYYZkHICF94XPbe3/3SaIrzY0ve/i9
z4Hw2cD1iVMKQqEs9SELEMwdpD7W+m4L6I+xh+ZKY1gLKFSmoVdZQscLeFyqA0gR1Sw0fPbw2Epb
y84ot7j3IxiQ8OARVeWNrspPENWprfliBAsKDRYshtmeWjXOP8QIVnYBfpQIxHMGC7FWsrSkwoSN
H+wB49N+haAD8z9SF8W3sNdw8I3w1/o3Ud0H2ka7M1rQAS8C+9phw1t2ndRzmvh0mPlGOhTt2uBY
PPK83q1NACN606tpbRpdD57OnuLJlpc3BrCLzpUam0Mn8tz2cWIywpmqTVhsjdcGa6lITywplTnq
p/QBBqVGWg/NBLR9W2pSyitD9CxQR/UFTbqK8VRMZKPscelPVpyxTRxG4OuDO0tV80FF4EwOy4qm
qV1rTIfip++79FoLVUEssc39WGwexBK54xPS0hYOx4DLwOw+blN6bOD3vwusicsnFar0AhGlo1vL
wS74GFjY3EJZBVjqmo2iNjQs87Bjw34WSnhmO1R3QHZVyOztfqbvwUbpbuDTkmNM74b6ehE+EEmH
8/fyAxFD+7DXEZPPmknpWGf/9D1O4yN3yJ3yR7ZLxVNHPJNFr3qT/Cg+H8I8nism9aQgrJ8g4Uai
lj5cRpCuhDeGCS8t0k6RS5QmkBXUXrEYoHMwLSaTYk4NM8Sqr0VgfSGuhVROZHkcsoknk93h3BX9
6dB4M8k3ZAPR+1VNPlVjs4MCh25Em3dubpo1eIEPvy9CtIXW3ZYT0NthOg/hrOAUi3B/9VRelTCX
xGnNl7uyc1bOVAgRmIBZqu0AEhNBbY68imltYyLS5SGoY0zDrx8fOi2WwyZFTFoSGzxKxbHFLERb
doI+MIVRI2HDMBcMGNw8CNtdnxfYISbsBVFc5BBI0G0C9946RxHp0tXGXgPp+QeApk6jC4M1rYSS
VjlrSbe8GhFYjCOoeBauleC7qd/XwiXH6t7Hatqh3uWnNO7MLUlWdiS53EqAxf7KmD7txIo879NL
FE5JFtnrkCwkHgTqEc8siE39mXYGijjx/8JNqbqjnUL6OuJU1LOTgSZ8Ck1RffuLjRV8DVMJ5lOk
iiD//YkE+D8dSaYgpFCFhogn86nSr1XPchXSUQYF0alNx1l5mw+xWfwDNe+n6q8juvEYiQMUx63H
QNb0UCyJUlQAwyyErgkj0ax41u9t3Xxuz5stcZXGDrmIhHJJ/Sy1oXanXdkN9YADyYoenXe70JQq
o5vHoEQlcwYLomksnODtakYBQnJM9zlGYybl/3K7D2Xbac1eEc3wJhYlzCVvq2AEgTbwIIB2S9iQ
FSpvSw6lhRkEcZbfG9vUTu4EkW62Nv3C2rLMD8fkqn6mo+m0iyoPdVz8UM5DrqyH22yn6t5fO6Za
d4lzBBgH3wv5KtDBom6ci+nsfaezmEJ0Wys59SjLO91Uq6MKfaxgHVSNAmgTjsMrvpDu5RZ7hE0c
SLgFBStRVg5L8bTcn+ukffak2GCpFI6/2qcNhMiBxY6kuYccTZwYvu7jouUovVs75Y5+5bXgHncY
sPOL0j4lAXaTMdKK6KR+BwdOQaNhR+x0nQBB9wp1eNTEr9n9aHKwzEIBY6us5HRZ5/ntnJVDCPVh
tEeTvXeKpSNJkU3mCgjEbbzB3bYWT/o46tuhF3J4IIKkkUtGQqtWPv+MhIw4DT35eWPgwipBzZBZ
Zt4kjrS5smHsZFedLj5usXtpntlwffLSOm1VHd4QhXRHCFLGPnkiSODR6V0TSYhBdk7goFzouk/8
HFPu2h8QaMeg4WUNdn5a5yLfuFbLiNxfCQ4v0iJeb3powqiypy70UVemsTGDKw1TyR0JUwjjtPIW
moqSiniJqFwABzr6ch08C04hKOMprYiMEK5ofxSevXGIvtwu8xBgo0GCjNCMxszzd7tyCUu8EW6y
ug1N8bMpYATcaoQxwh/yPpnEtLdrGrzsgtvtRFbpez6/fb6YVYO21AsGXsx2j307z2rhqgt0IgkL
uLDFPn7jqIlAG5hf0AUq45SgXdaiAE4PYxWcaLNS6PGlfWK8iiQUv5e0RIB+hcOg8GfiGDkl++mm
K4eueiCh97eg1g5UahX2ZMSGCGd53Vi/J/x6EBXSCwNmNEd9cCuDKZb2ALSxykLkdAGHeo04g7XJ
MN6MHXm4v35u34MbayuhB488JJTPgyRRfg1HzR+jxB2cSBvI9Mc0TZbAVpxDIdJtyz8Uq9cTpf33
TqLhLufJvOqgSa39h3/9Csn8peGQCOwn13MyKl1k7RyKAkKdxuNt8FsWhxLq1q56R7idp3vGi1iU
EwzyWAXahDl6IwFEq3Jaif7nBjUNYNKMhDdIoywy+Cu1HUFTc72OUXBRmc1CbeMqHeuGvsUepNji
k29+a1fkc1zRea/cmk1iEw+/b6QiO2K24T+ILfAPV8Zl4eIdFA7G6+CIUTnav1U4sq7l2DiEpbpQ
Hd9M/ibDZNcRrAXUfVGauYDNpCtxYidSQ/i93Zb8NmXmd0nF/ruP+C7Ck3DxCVcyxjqwmYkbWsle
xQRO3HXQJxOI0whDb64JuUgWGXdDInRJECBueIGx6YQXc/t9dRqDmbumF8fmwckP5tXcKQ4lXseQ
E7wjAZOR44W7Pnzaaw7JnLKeLrJ1cGz4fV1HZVNjQlVi4C5CWXjh/qp4pxvjSL9TOvMwHe0ROGwr
vUc6912eo/YyLDoQ+FMv5A5AZzmJXQLNgg/CvE5fsRW8OaHzK9iL1FRsC0eKID6Vsh2mDxizZiXm
z47bmhWhuOaME6ypJQJuy1Jkkzh8UPvt7odRsMlHaEeYSn4wp1KQZ6Q96hFPsN5WMJoA6wajwazg
fc4g6wXuNAGI0MSnRkSYstpA4xgtiHh2pZVofQwkc7wPXRsp0XpEdDrry53pCN2snb7IJiab7GHX
AV5k1p+jjV6GX91lzOTrLUFcgxLgKTzh/8sGjfzno355pywSG0aThyhWdAjwxGrV2XZqG1S+wXK1
5X+0tSRIXVjnn27CBAkfaXldzMt04ooA9CEK03bDWFyDO2OOTqvehgOQcl1MgQyT0wQtX/1CPjJk
J9q3qfpwTz+O/49kd1khZFtPEqvtWiMXb7+SmlolXypkCOy5tDORIx0/deNKP1Pdf4r06+s4h9jY
lj2hRC7USenDfQNLn2J6W1FlLV1vVLFGLGVRjXZQbOYXyZt/bWcKLdaklKFG8tt+HczS1bwiRgbK
bZfz4C5XvSW14PV5T+nVz8NIuCbdpKbYyWjfg7qC4Zg4Jzy42ZZAlYe8ZUkDR0TPbqqLoFwOWfGj
vnex+uPlpf8Ly63gPJq3/eCPARCvNvlWDJVJlI8X+D4Zd5dv370wvhjL16gPxCnHLhEyuT5KN7tG
N74y6oqC2hgFcK/CjFGVO+lbnA65Hqfd2qtYyK549wyFpp8rFFxBC74gO5BZTWCl81vujHSjno20
qr2v1VAEPYC4Faa0OwB9SV21zVIBmROZOrioU3kDN2ruSumS00PsG0//znfAVBO/0YOW0NiT8Z/s
fRrrw/tiEoL/NXdkxDD20fjItNZclcT7xAsoTQjcUhhhB29TrdukdwEDbll9liW0JRLXYEuFFolW
OoEFKVxRhU7HFHb8+Y+4HSA+LF4CA1OHKFyS7ozjkpcRdAWLJyIX3ByTR2HclnUVaZVvVgOb39Kw
7oBOVD8C+A1eo7C+Z6Wpvsqg61ceATVhK7fYPTQsboAexDwabbx+dDeqwuWqRXlsVFxYaOEAFZHo
avxoVxH2d0lVikI3VwwGMx12qRpz+JGqxkyl88G5lfgtC3CWHcXRsnH7q6rexwPLFe9cA8wZPNse
0L+4zU2wQuNbgxXOFewXLSh8haZHstJDk0KVOg6rc++kICPViYox5qyzsvEwzZY9XoYX/rJPauld
7mejQhjxHxlvHKsSr5GkhDYgeXissZYIlQp30xi2UuZAy/OfouGnUcVKVEmXEuNF0lFLt4txQdMs
+GCdTcdPgE9ZVKjfYJDMYwgl5hM5e9zWZ5mocv/aEEU5EZLf7OymrHRVYGC/bStlVaX70sFOvq07
ZHfHCKBvsH+NldSY09L0l3hWd/Aoy9W0PfjpAHXfHxOl3oOXqb6lgtSHvWBcMcn845d2NqAfdZIG
heURlmiImLyCebTdHwyORAHL1FCtI3WTi7oc2C6zdejbK1jrpwShua0ScTVRG6aBHRVcFHxc+hdU
1/beVXRRcKaH3qrLX5WQAogZT6/8+1yUAntq56jliMjnB8TeIqA3SXthBUiVwbgCbdSk7C0Ec6ez
b9M8SYka/vXCWbI+tCg5ei3WZj1HsZDDndyo6LFHLxNSfQnR+PB6dTMm/wGWaA3moPz1yHgvMnpP
JCghZNobH8/oyTiCL+8uOmwNd6+17L1FZNBfCQfwRotoi9v2ivNVvEciEvwKyW/VBdakDtLBv+sH
e9KRKdA2YX6qtIL1sT0NkN6D/QrnJjK1mKYJnnI1DE+hQJC5mN/ec8gmErU/KAU03MrTFNPGxzmu
4Z07E9nXvYZzR15BJIH7pUfjiEJx/xhPre9hZAMxGiI7yik5543FUl9qbdbUMcPCLkZz8JwBGDQC
O9m0r0HhZIHIn2KXUufLHyDn25jGQtLHZl/hh0Mkk6xz/KF6icdC3lustsD+k9yHYt2krzK8HJeU
R3dHOMGKggbH5DLc/p6QR98SVwXZxwz/4kEh8ILzEVaguJoIo/GH3hoMj19sKY+Rye47qsVDKWbt
AbzGwhsLf2hSRE1b5Ejn4OP3bx8/PvfK3oR5/4cEqfDWT+iNbKDgspAXjzzlAyQxqBbehlz2Goeu
m9wpGNlq9Pc28qw8pxwISGoeUGSCRQdGH2uXFxR6O/uAs/wkujhrx2liGWjiuYfHu+7cid5YB9wO
MVfiB+PLgX2jPEu4aFe8XH0HoluICYboY6IrcGy61bQEfKUfiojLKuxQCpBLK6V5ibHVeOJLtGrb
9mXHmLi1XguHFGntNZg0npOxE2MTSfj7zeAkCTO3yyOYDdY2QKx0tKhEGQUZskFU10YnJN4Rp+4w
ZbUyyT+aKBEWzUcFadptPDuXHVl93OMA3DjYerHV09rZIWwZI3xUQaS9i3HYerVoEFx/LLglWzRi
2VH+A3+7yHLRal4mLYBwJIneXInjaxml/g9ZJH3h8h0JGV9A75yEw+423p1wcEzm9LPyd5QGiYVL
UAt/eGMgv8UyAiuBvCJGOyE/yCWwIxdpoLojOPY83iPZkpsU6pwtNCQt/lfUj0IQDb+79ZTxrSCs
2UUxQxD7iEdZN0MbwdSGyJqnVxOgNzCvMQeD1iOvZ5OmZ6V7UcYXhA438OovrwBBlTbZD3IvsgcL
PebKrkSy6t52/p1zYmOK26XyLMllpy6oC/anzzxSyDAclKof+5JvJSohgjsrHfn//Zt+SfXZu3Dt
pQCF+veadfBf43tD/snEr2j65r3gxflp3MMxM8fKT2dZYqZ1WnzE/cFfRAQHxN0zyCCiwzCVgpgw
jxdb9Gl5de3S8gHwzfqZoMVLX3J3153kMN8/nN7WdE0u2bHhVLR3Jicb7kxsxNkBgYf4Khk0RfNa
7Z02dnAdBblgfT2k9GNgksM+UKWpB+zCSaaPsAz+V0gSH66/ITuDgMrVNmnLFhTznaD4f+WvEAvU
pE539noRN+qTW0sjv0JxAUKUNbPiBlWmmqdVZX5mJ2BvkalM6Aa2LXOO+KNR3+2CV0F6TE7yaHHK
1JBJbavXpVBY0THBk1wGaduEkZvQH/XZL8B5h7KW4106ngDLwgI2WW2+L1nx1h1GtkS5j4EVmSiE
47KSMZiq/9LnAUwidgAN544GbA06iGt+xYNEvf0m1BnCHdO9Sdr+BK/eBKF3nTldsA1B0UNEqc/n
ZwO+q/t/cRnhHMzkCUU4nZPdJMklCc774LOrN9Y9J5oPy1mC4okO09JPZU70r/WO123kfgSlOukA
eBidGEB6hmBROGqO7+iecBKJtzevbcSdObdzWf/jxcE2WtBPzORbM1B/5n4XgPTKBgFjyHjBoJ32
QD2Zd7YOc99pn+vdw1wJEsBOkWtxVWYCLaaC4A0vV4swImr3pBEyTZvV1pWI8isBg/9nH33ol5k2
fyI0YGVGxazJFlAoH7y1hmU+FmwMjJqh4a5Mgk69pzd6PnmJZ/MWvjnLt1nMXyniqoFwfzYqyY/H
SwvULW1WwBCG1EU1D+SAhcaLky+/84fbXlravutaJEaTa3/05OgPc2aTJ0luqDjmZakXVsw3dBCe
FpNd3LuqJ8LsY1L9Ebh3MzaSJeGuuzXV8sxyN7S2bYZr17+1BlHPjJ8jOSpmtk1QQuSVloRoT8Jr
hZCDNCX9HpoBel4MpoEqQ/hPThniGCkES+6lG7VsRQVceUXat5l34QcvQ9CgmKO/h5SKLlrtUpPR
TI7tU//BI3t7PwbwDB+JjmgHqExZ5JLi67/orjKBO/1O1iOjgDB5nldd1JVmk9WJ8ZmC2uc7WOux
OWKfDwJmsWwWs7AkmfCPMdJJLC/Lw9Wl6xms/JqJARELyY/bbNJwg1rmPgGr9ioMpjQvsKaJ3GFa
lBbgixmaYpxUty9m08R5bzYevKSKe6wG1v0TjpELmABWTfsBpjMxNN0DJpA0rYU2iT8twdhVKvYH
I8yKGySf41DVQj2OBnzGM4WXbDXlww07EnFMqBPz5g1IAA9M5SKgA0thjUJ+8HQwqrQGCgGoWhPC
GyKK/97U3u6ZXs6FGhKvoQyLBdqFrwJfhta66Tf8jKdA/z6J48S9n9TWcKPTE153hZvfKlodYMmV
C4H60Drv6UxE8yXlfwNmEAo1YYLuPhhPveEqd18k/dmNgQV07TXKij1EhK6VE3/cgGpmDdWUrC3k
qIA31cptZuMUytChUlINcypoYOHZzzJmkEKCdQWtql8geeIQGllP8tKw4vgtju/AxE9vh1clg/ME
97m7FfAHRF4F9iO0r3tA72ZoTIEGaHOVGdAtNmOxDSVYQ9bfuN1hqLIb8z3wxFJ7jSqqPYMXY932
UZ85W4LHWVU+Wy2Nss+SJuGhXAISEj4mOaCD+xGsIdRu3vJZo95jVnO4VvZS+2MN+tzq4bO8HfT/
YXOg0U+/ijeN+zUtORXlgDx2X/uFnshG2YSqVy7Q/DqMYXtjmM+U8MgcB9Ll5xv3TsElCEEoEXSq
0QTxr+fZ4u12j2/xTuO3vcFISlQXzWuWPPZAg0kosGYVDLv2ELaUjir5IIC/TwnfqihpuJ2Ma83N
N1xYGjIIF3QUsforsWtNPizewNcINtjFlg5J0uDG3A5nmbWyKp9tFcufvupx8XpEPyY+5E15fOXI
6LqycM3PAYxce68l4aXu2yA9US0fr8XeUidbuyT5VwCtgSEAQgua11bpayETCU1b3eJutTJ4ApwN
LQRIrognrunz7vStn8dMEVvilPuOG8cdC4MoGJb+/uVSSHE2X4d7g3cxr/A+uHioj+HmgkfJPVsp
vSE34WmnDWsKFWQBpYpjgDadXQy2b0pnB2yM3uP+Ch6yXeZRLJnTIYvWCMhKHLqcLF12SHXOTsET
SK8TV9yoIapX6kkeuMUJZhHN0clXCjQ3go7pjMyTa89LAA7ePYeVVQceceNGqJrU69sIkfIMgv3a
j0numT5H6A8iaZZ0/D8hsi1OaWKS1vskliIlQqZwaH5FWgg4Itt3ENaL30ZWXE8n0YA2PeBLGTbk
xNRGF3+xFdQUyBliyQjyU8rhemOg5x7ST6sjlJD2SH+ai0OpbB7Sh6xc/mBcWYHBFHr6h1lt6Fee
PbpO60fPNIXnofk5pTP6P4tU0Mn6BfW8ZKiGypTfZ/GVUIjozmEnQG2LxbFyWQVAENQY4sAlPocy
A5sCLvONHKh0QRcLu7H3aW3PuOL5zvxUDiQztM1oWewPaSbkrlgUiCyBnLgg7wlxVc6GxnebGr37
jC1mRRsIIW28ceUE43tXrWqYamxI6zz0lToc3HV66BQH8N9XaJ8il1BT2F86AEOmPHFI4MctjVQm
qD5vJ99wF+ignSuc11ct8gaVyNQl5OzFarWvTlM7I2y7Xht5y9rW76IaMFq68SmHvZu0v/qCv/7d
fE93/zoc63onchqBqKwapI43CaYWYVQZBMoMfw6IfrIllc7JpWpOP+bssgmLUMJBuiUStyPE3kn+
bmthYGk52ftlpqtxBxgSjdo9RHDb7aAOqJXZ+fN7Y8OzisEGMckc87ozH8W8wdokHtaW6m/0OS+7
aSijj15Ryagy9AyW1PXsJXv/CE9uHEMGyDNb/W0QWrrtjDfIocFSJK6ixU8ycZlS3qBqE3MXUN73
nTnLnEFpcQGHObhXu+N4LxthFrVTsWkNzZ4jt7VIfKOM6EM/dp2o7QbYzr14IEpDLwC1ZJoFF+jo
+yyTUx4DQAH9bv7pW+3+SvaIEecnGXmb+1PJBBtLqCk/ue4sk7LMCDO9cuXP92cTHId180Bi7ROh
irj3D7hyZ/z4HeggjxSQ2IK3XhWz8hFxgtlFawG7xb4NfvnfLE4JJpt0IhgXgMl2YoNzJCiua6LQ
UGYdwG45G91y2ha7uyxYyC8qpi5FkCSSpqPPK/dc2qDmERCI/KUCWFR/E3thTeNpnVScE+pB9WTP
4IQ59mO//ipyq6XkIG38PIFuktb4bO7QJfKgW/QiBOJZ6/EomUWdr1lJCN3X1mUBRLR96aIUuHL5
+xhxj8oR8+hnWYyHmc27nfOboG2TDXqzdlS52sjkapDMnO6FGTIW/rYHEbJ3MbA5QLOQoyrVB4Q5
nPKYnlUeK6nFfDJ+laPypEqMcVeHergtoIl3JoaZMuj0z9gojjRoY2Q4CZz7ZeV0g3tD0dfW36Bh
kbFOWUbpoRdYm8TGw7XRdUshBLmrMA6c/06EN8Ch1W2qtX1VDZgPIpEKG13tImRJYR4pgziJkUMX
hhrfwdwpLOU/JjTSNFPuG02S3HKpk9h431nyVm22zyKGaf/2qr+25EX5YqamFpasMcZd3DePZY+N
zoKa0unsFmtSp6t9qS3xOcvFP/QeT6o4Shkzb7nCF3lnrnk1S3tAW7WwYjoinUBp7rf/Qg52kSS6
bpz2g7KfKMA3q5+hv0jinuD1VxaBDmEm3bkmgIrFTqs6TMvYw1AbcevaNbVNfFPtyPXAWChvCv7J
kabfbY6SOg9/97lKmABC9mYYzn/4g5+q/M2ygrm+dib1Ss+CBd1LkuSKTzBQwmZCrW3xBRBq3Fvt
asLg52t2OCGxyHCc9lNFO9wM19hxVc5cEvPadPt+D3q4HMJBTzYS2tgOz7NlZNkbDvuV6Mc4iflw
FNNrZ6Waf88G6MV8g5N1+ztyxtt139QWgK/bhDeZzJzCO2NCoyKUfcw2hEpb+vxBmdgY4UqqqF5p
B/sGX2jH1OtIv2LLFl8ArPQnOXp1PxDCW3tUsKVeI7D9sViTsYXJv7Bm+b5ozjiANHL16CI4onQp
4qmbVCs9Lg9el6Q8C3rASwN5+MRhXMxKDCC895dTyCGqe8j1w2RCbu+qCAvyE+wMJx2Gq1S9z7dH
YDUKNh3iVacG7Futn/YjRDscwN/pN313vmUlTxt69E/feQqiI6z238SupHYC1TaRi9Pi2iCzi+lk
F1BTufrwLKVJ2h9f6EZ21rBrBw1R9UgFXhemELlxxY5Ovmnst27OuMmSuutEekIKqu7d3NgQ0Nvi
9g+dCuetCwi8vwdrZbe+2PgZ8NF1W39Oo25Ohc9ZP4oMeOSZUNwcKs0+y9u1B8Qt8s9I2MAxWv0S
3iSDToJgmIzx0R/EMhqKi9uNiSPXvIc2GfOjDObKFG9PIj6jl4SyfUTrpw1gxR0D4VutmPPAEPjE
r2sZCKpY01ARvPkqHNtaj6xvvdfojOTE/P+gHrNupIN7KZhTdNvNJmHETX1rj1yjLfwmWQM/L/Jz
ULX3JSBjeoCUp+4tNdmFbXZAt89gBjAA2UOBxRq43aEwyWOBu1/6BmNndG0MbJ4RRXclXogofpQZ
xUv73D++vWOz7+AjFbFZNTprwktZhgeAyNqDXdHaNCKD69FBwPKpWNPSW+trs2YpWKX8Wwea1TbP
ZCVEQ5cA+GcQEvf8+5+LjfiZenZ8I5kUp+lR3l47Ji6aeQ2abh2WAWRzaZ9fJe9FQ2IWyhUxjlEN
/Qvm7zHqrpwUDEOwQHF0d6UsgNi2Os+2kReT3+3sigCcwpkRIxKozSTDjhgC8UsV2ZOMPIc+05lr
TTqMrwDQ721v1WqK+1Gfna90UfqGP449R+0ZaZGplif8+SVgtodHqPEebFEewIyCn+i/jX1/DHuj
2XadRiDb3tQadWQVjILWsMXbFv319R7BwbyFFWS1NxtNferYf8WEJblRht5pXxxV9RoXSPmd4s7m
vFMW3eByaOaKRqQ+b4IidtL7j7zTirSLmeNR43uj4Z3WeW0z+bpKQSn2wveQZ8U8X1j7NdD0/7Wo
R6bz7I8ypgN2QMG7QJBueUL5JhCRmhh9L5HaxG65ukKyO5Zamd3dl4g91Xv0om6by0JWmE7gAikq
uaYw8MfWV9yVYCxC83f1nKPM+bW9QA7Cn8NgMcn/hsjCHoenC4sWRcjDtuvFXchhjJVy+4Cd5bDD
RLSZDsn2ke87EorVFsuNw5AXIPoNbtsLtUsjJHwDzv88JI/lJ9A/Qp9XN8zST9QqDVsoeKEdeHBl
nW1qH2X3JTTZtZXlsElk16EPaAST1eg2OgUXJJ5B9vKFWQ5dw8PF6kl32i3PhJgl1NMkvSl48OZk
IQdOCWbJh0tca2mUY1G/BcQzhRypT8rycOxbAsqq2McuGFxS5ITG7dIhiJmanYlEiNcugj9eu7/6
bZ4ksSZM5uwUIUwshvzt48fOWCSQ4GiJt8CVk8wj7Cmp98e/98eLMVMxeLu1ZB9ulf3fXwZZds4i
J+yRH+dzHvHubje2n/JhDvF3UvgUxlbAgeM8NTZduL1GzZewauQIUTVjEboWR8IAnKdhbmZqWtIL
Jfm14fCSFjljTED6Eaa0g93czeOADh8SRSGhn9EacsE1gLlZvf3ogfNYJwRhIHp6qi/qI1Opj20D
wu2aIF4XFBl9UTtv55TnGUxUDdskSx9yM03ODftgAClHvW7P0dVeQLLPLHFeb2IYTiZ/zHj8vqo0
QOHyjPhgt5gMavnUemIXREpzP33IbMk00AGv9cWo9ciuApc4GqqXoCBlIkCqrWxr2Xu/nP9Gb3Rj
AVYY8NfJr+vt4q8/9pLYUXGdeQGfz9Dp+H/x9o36BtAvD+DG/GyOk9s7tP9tJsc/uYmPl2PPCar1
UkGJXtBknqWTB98LiSovNQGKpo/laPREi4FX4c5QClK+TWRzdVgyw3Jt4n7FrHPLG9OKqgD3/ZF7
IxG/5QE1Dg3uZrSxA9NI7U2qSxQzBCcC2NiZYzUtKgkW9XxdlnlFBpYIkobaz83FqLskzpB/FD/5
Uv0vSgEhIsc65vodFMTvOxuUnu21uwd1bM7kUgsz/P2uzu6AWbSKuwxaOc1I+X1yrDUGHT3OxtCp
Ou2vYPvWv3pj9QvCXRclU+KNtlfMTotOGI0/FQW/wEm68irfp+9dUKo4+YKn04ZcUUiqynGIMcCW
0H6k7Cud+RnI1UkrO2/6MsPNSBjcB2sDd2t+C7vrjUueZX4grfyLzsbw8AWNlv/5V97IYU5iWHsb
AnlJt/FtnIFxtVUTCBDOrk0JKBkfV10Iy1WsAQ06RnavG5jrQbbzs8gEEyGvxAJi34YOQdKo+cM7
QWttsSuxJXhG2H+uOrq3epF22SigVBAdN4h6YRoOaeRfP7QAKJno2XUFoZNmu8EF6CXy26Ns1jF/
DnUq7tEcxPUtq7r/xQwOMN40OitTUdxWgSGy33CbmQq4C1gYQgkByniIHgsnkdGQU+XVwJqxsYMH
JjiuNc7xW6VhPxCLZf0lCnoa5yjXeVZUTQpHGgshAI6b1+/BOVUJgDWQeC9IdDGQaABgXaai8Yu/
zKCLvxyxOEJGvufd04l9DVA4p5qlG/WT1NsuCWxDCM+66MfgIkChI5KoPq8JJykWuhkg5P5m8CDV
USIKJKOZSHlwkySEO48ql6CSiHCtpvS0wGEddLWxmGr35SrBbIYd84K9XcizGiOpXv2l+xOc+I0W
X9cHXeat4UC2Ieru4R0XNGxP55GtoImSILoiHo/2yyZ8l1HEQ0b4HlWls3/ZVU9axJDSPXfhC7lf
uyKA7cAr0jJdMdgu2Zp7on+TkVsnakR3aPew2ghqxHFmn+j7QYnsnS2c4jAPsm6PiRE+vEpXL7pY
bbw7PFgXxtc0yKl2JhJL7Dn3K/+Lm+EP7vPhfz8qSEsRUKSeu8SQYgJa2FSk4alvpgjDWHiDZrhh
mkhx7XtEGj9VJ+awuDtX8krwUl5Adzwt9D9FRqiHCitdqgThxTUYfjgw8jkQPwB9O0Id3EUioWOJ
zCs/7dGRB2SBXTHsWvVHdX71MjA69uQvNt5+ol3TFlBh/W6/SAMXad/9fL0NVyDmhJ/FQhLynaOA
TmDgiuaR5PSvbJq3ILNrhuLc0Fsspr8s3xvT6BHG/6Y1Cr8YL2/WQQn1S7yu1OaLCKDutkgPgBvC
OyxV0x5QnM0BdGBws9T6YtZwz8FknojHtOSnm1MtEsnkZSGUrN02WM3pW9b7eNlAHZNiTV2LUZaU
bwMjIwSfwIwofYMOubeXR7ZjN0Km7l3IbzWZakvuzOgztv115I33uaL98hkbC+HLmgyv7iUiiK0p
4oC8bVT4TV3FvZAJWZCH7LnUNpbfQ+H+XuDiJOa9GISC/ZqpeAsjINyr0xRg9y+zp/w3FsvKTPmt
pJ9kBddhHQvhy7ulkRCksZez+VoCcJ3kXtkVmAJd2nnPAGkzbeIqPQxPpuNI7dssHuAKvP7eeNzN
RHAljElW13E7Osq2CVJ6yaDnJ1tA2W381BiRD3GC9TlzGzPRFnd1Sy3juV2O2B+2VVzk9VcnOYq6
rFkZKkY2peMS5IuqCLy64jX4xoHL9s/BEXCRh94iKFrxw/nHhCarpGM2km5jV1tXpkwLoamlpHCX
QOHWkW20ZuIEULcgCkRms1W/EsWcnilf69FpQ/dNYnWwZidxLlpkkM7mtWXdpwpho+laIjqPaf44
Ka5VdULLOjHLES+cnX5k3nWr3RpNMuTOlgItBytq6ua7gN0E56bTbJSWV/Yyb4PYPiZc2vXntKsQ
+XfdNLNxJT2sFKKc2OBV2Uj3D4ybpFKPBDGtPKjMFBbVqGJZ44CharpVEI9iTzAJAN2OaNXlD1Wb
RcsxFAwtuMT38GlYIqvteai2fqSlY++2DBbM+oIoFu1e1IfZMj40SbqiMNW/f/3Si+a4dE7jH55y
J913R7MjofgwYc2WfW6QpuyhJJ3ioor3vI6CsanKyuhS+aIZmoH/x7MbnIMR8BuXFOosVdebqt+f
yQn1fqGYxsXcfYoo5ekGoSQQtvRrKieb804EGzkEYUxc93o35tA76IS9xbyZUX4VK1ul1xFluAS7
dGHIqgWT9z4NanMUTMs1S523h5i+3l/L4sOlfcTLlMxrkl093Z8HW/9Mk5OC83L1B7rKUmd+1dEO
LMmFDLbyf58Cma0RjIMcESSa5awUqUWcHbdFXnjVolnZZwDq2mXm0Y0eNZNCCyFQDYL7/OwXJT38
aBehtypcjyqjTfNkOVFsbuR59s7HKmgOXlgrNRH49IP9RcbAElhnlkrxrzCEqoT32SCiU7mwCdlp
qKDb0bi8cKPIKHfmulOT4KJK3+dnYtcLhwKSLOPpfE0uSRoTjbBq1oib/D/yjTOp4vShaqKhyctS
MaBeYioZhOyAmVBQcIdte1GyiSPojjakt62qaBQdBEQCxydmMWYmvUU9q7A+aivj4zFztejFipV/
B3iRdhMXxpOffV8F1PZYVFkEDA0Ov2o96rbr8ioF2m3nwW6M9V32xlg4RvXuaiBnXv3ZZ570s1bO
MB6GcEiAdTyqGZ1eIC3SKIaPzp/vXZOwCM6RdRdoTOwp8XneDLzoVZO4CAlPW1VRee89R7jYVF2i
B1v1hqaILRK/3tD6+JAxIObkvmufeGwFkoOnn+s3t7WtYzhwfnqAn8TxwJzg0Eu6WSdVCkm8GYQY
cKa4Sh8nO7bGEale46qeMCNxuKI/JmGBS0l02lnu5VBoMvnzeIVDqiu7+fYG42cynA6/bnkxceg1
JTMS5I3UFYH09mf2JZkT5pPQB8iC6VwR0/vx/QNKGX/SeTZZgPbRGic6IqIkOYYOFj6Tk4oxfDUd
nVbj7CpgVVsXqclC0Y85BNc8A7JWz9812wWFy5914Pg4/DlhvlSE/+mtTEi0ciz9mS7D7nZYfR9J
Y2nrcYLBEhyDX1YxayBTkoO3p5BM46O5HLLV5cJanhkCgX8c6z7d71zWQHTcjNLIvbMJTAzIyujx
GKxWZy08MhxXzQh9LqdEMXWKD2QlF23dwuXB9EteMl2jjoJ36zT2O7eVyeCikJYa4ZkuQpXvKfCm
rV7+3KhHBP84D8DDvXQCw10he5kYCPV8OQMPvSqNndimRQyWciSz4vuaFUSeg9MfFj4F/ZJoSjNJ
y/iBlDgHyZ1RUiIejzuWw5YiMWYA9butPXfpcllHaYbCw3YyhaO3iNevelV2xzr6GpqQqc+TDaPE
du5GjZv8ln0G/0bmXHj5NPKwvuhJgwoM1QtAjacEBOx/2k97+e+0p9uM8QdncRosRZHAjpDiubVr
46BGbkHed8cg6cP61OJrbH1y4BA/5Tz4hmqnp497esXczsS2CdyzcebJfwRhlEAh1XF7DJpWGvXv
7KE9KbWtwpU+Qt/ue5m8JRmSXXoPBucBD4oSzqA4nrndfpJZusgbKpUDBgM92uhAAnhBqH9iNsVs
hQD5cqyf95+RR03FKcJ1ReUaBH3+u0yJPgX2NjVU301Xu4PIdbqYF33NE4jhu5as9uNtMIQu1ZU3
bUeqilnVG3BL1vUmDZSW6vQZjlRlfQaNKYg5V1Qe1qomHY7WnBZZDXhUifwgo+oLY9lAQfC+Tt6j
HOUnRpUYdPX9KyqaFoEjbaWoq3OPS01Mup7QtQ1rLIbcpxnPMy84oviuRVSvVAYrzZAAedX8nHt6
1ldagG13IUilEVLqR4QaqwgjXhUBhqplLaNyNYX4Her6QtwvS3bwopeIclfezdfc2yDn6rzxcN17
FvLzy4RrNt/SkIs4hwYbTQPoojHPFRrBqT/w7B0VDWpYAAsZBEAZtBWD+fKp+wiWp1REAIfHswU+
32ZmEcF2mW3wh5mAN+0i6hvM8Sb7TS25H+pglu18qYU9hz/9/2Z5cfPmN8HYTU1a9KNoxWpWGjff
zH/qtE1MHhfKydD8AqtxmCd2jIHbpbZNAQkXsFGdDQ6sNha08Op7irXxk4HBBJXcafEuQT7KY//v
iRAR2YZ5Vmj5Kfd0yzXahpwaE3Yphw6Ue+r2L5EoC4EowO53ycZzCFAsi5shFBbR3r7p/3H1Atkz
ecIgbNi+Y6takmzQeNyQaIh3TvdQFHQBWBKOGBkSzaBtdeHEHkMvpnGqSEYfXDecfsn/HSkV8+Tu
PxHrEV1t4xzqoLn7CYUGzQQoJrrjVetyUv9kYBCL+4zeQ1xUEldwTiUBPI55oD+MdAki3roTGsLi
c6mU0tS4cvcDSp44Wi3wSuAV+kYCKSotdXBe/+zxE/P2njOo/cpIBHRacuyAfCHcMLRkuRutelWp
wADq34JIRS5kv6Cp4/0KN11yunUqIPdxr21ppAh0HsEoCF8z17P9C8s+vzPs1TCB+lF0Do+VVn3X
lbVSReHA5yTTJQW3aUymw333tK0IMTT+Llp61wqb1Wxe5RMo3yIDHYrr+ammT5INIpxaTcBvcWEj
sbU2XzuA0fbIe5YgblxpvBc9N0jnfiy5+Djv2lV1fkvM8/vzGguw6RY4fbSvgPArVYHnfNhwZOum
gGfa9hVaQ0QM+fA4kKpZXWjohv9nn14nL+p2LaNXDgVEA4Tp46Ptb/2JKplfGnkYF4tbinLBg3YA
raeUmiZwnOsVqXARFxBIXkT9q+ENwu1hXZUFwYm02wxmztbm1+vkolVFkyDpzheGd+xC4TVEwzAK
gtPoIfu//IBh3u0aqjzvI8xTeFlU5WeH97LZ8DzySODcog5oEcMYYI6jx08odRubdS/R43jqQQvm
YFd+8dytUD7CU76OksljbaJKG56NPJPnXwK/Lq6mQso39pPPHwiHdNt54K32cRhGCKjDt9vISabN
XYu+URIQN4LnmnFZLAUVzCnxnwNAIEkkeEXC0QKh9QN9Cahfn9D/vVZymGMFNXLWizq4xFp9NvoK
uEWJ8EICMeEGcBPNoUxWBMybqVFsdoQXKNbOCplsrJ5zLZcF2nSsjkwKgeJGPnX3D2nVaFgNbPNz
uTOry7IoSQFG9CAHaz0Sp/pV6dt4J4a5QUsRtsiPMUo5OZwL9wtk/QHRJCs6iJ5EruZ0G58bbNHK
D5O/X4YULULe5Dj1eStpJ+d9adWDrgW11epNAlysaLK5HmFYrJkw7lcxmOmiD96SypLIfIVvZv7W
X3uqiovnPSbllZ6uQdzWOToo5Q2eypdXflbLdpSDwEWjrf3nFqtKefupeoMwyQXJg17q8suJsjXd
2FSN4J1XeS1PJuIbZCBByWPE0vlwpEiKqabrknhpb+KY/MJF9iNbZDeFzvvVbDp197JwQpSML2ME
g07ouB9C3Moc7Rq3m4X47Sfpv9vEDe56QnSkXOHY+62i3FcO99HIbpn7GU5GAHHzSHvWhWjeyF5p
CqvgS1J2RLVuN4kUIeuG2Su4pEzi+Pt58A0XFsa+L+q8ApogkDyunSQekAftO4BoFkzsmwk01Ki+
PWz9QpGYG/FxDkYk4xnq/E/iT/Mpz0EuDUdqL0K3rZFVIXw1mJOEGyMii7awg4jlwp6uNsyfldHX
d4uO3u4G9UmnV9PKBRuq3Te80zOkiCZuytteRMzspiIlx4PJgx7/Fe7bnkYKbD1MvvCL6r0fEICM
EIV/OYyyMYVpCsuX7xEow0CyA9AXQTAI1fPwx7jexXSNF6o1AveFv1pqO9kH4B9EIf4MI629yPg3
29MCGx+Cz9OKM9s21Rs9stb3XkvYVxJx0jYFA4kqsoJNCZo08DP9kutAragTKSfTNG0RV+aknD7q
UgFHlMHggR6/qRmx1LNjXocQe80pDf8shyJXhB7I1od6KT5DyutbBWo9o0dxxieiAhRhAAodGzZl
ZcVwspy3rzRx805wqMsdpjq3XBxiRxZnl+naQCof4F2ENqUFmW5SIJlexmrr3HDm8XxOsWx+HVBe
kQZs6oY5EirYcww/SbeY13P4fiDjkAbXXuIh1IctkUuKzodwBYCs/3UQ5xfTn3/s+rnrbBAeMbiD
MueVd5kBOQO1Pppqb2VvzwgOVAUSb88DfGbij4iIEjIGgMDRZ6IIYu74JYHxAYQhYcBx0k23lWDh
y7XTceSff04GyZHFf7UxE3oNMyIQ9HXbFgG+vsSBpS5IKGmhSOBS6K0ddl6s5yv2nXHrYk4CKiMV
7pgqp42ooRGR2+N0QLydcQtDYxk5/Czeda/yzDkT1m5AE+t1xYjVTdZjQPXfuLwYYc5QL9eGAjlN
8zQh1wS+nD3ErG6sMrG09e15/OBLla0dgjInntJqdA3oAZQdYT/OjmYbIL/9YO0EDw8vLBby+Yn3
NEL7rVE/3P+87FeHAdvaF7dA7mimSSWZstqTp82FalETPV5bx569/hB3sefjiE6424KxT6UogKc4
zVvoDqj8RMzyUyeh52gRB8ASN3jU5DiehiMTymikywuVaMWHw2q2ep80Po1otruW05sIxIMdSIwD
XD9WE1aSH1+qHi+B+4hWME3431vQuA1M2pPYuHRmIjjqRAwRr/tPDclaB+7DfTW0MBxHdEt/fwL0
Jx64qiyO59eNhPnHiB5VTXvHQuJp88yt/F1RTbPhixohygh2fxSZiUblxm34KBvuM9XI7vA+oohK
TpsUsBeF5RKZVAnsqbNdUzfBlVXoSI2J/D4rU9xD3IMZA5kOxiqz0Y1rwI3TkA1yTPu5lYKm6yzg
MiWoxKASwPSfk6vvz8x8po+ckZEBvRQwmrvmLj486Ym2bYJ2ndvrBrKMqdkdbGXNXWiNmQnpkmux
qQwffqTzx5QMCcun2gSOVIyaGs96biuYeg6DkMzTQOp/8H7GzdrzooKIciQsWbRPwYKsdWMSqOZK
zr/cXA/J1d+G582dKutNd4pJIApP0WfziLrvbZcLAGbTNwyt3RPdmG/K4ZpmwCf1VBGTa26X7vIX
KQHuEnNwncAGzf2QwHroj7nVzytIpHmbUD14cr+WqPjLb26LoqCT0EMqvvwYSPXYxsHnC7SQ5fJR
pMh0iVYSKAt3KlNVVCnipvqg8pZ47D377ZXvEigrC8C+ZL6luvobgJfVJM4AoBDBtYBDFSF8VsZB
ml16qO/z++OV8Hpb0h+nNlGNqP+NgV/x8gWEvMPM/iVneFSEeejCztWRd4zz3XNvqdbO5wjw1Ib5
hIKVy8d63SVw3bK9dW8SF8p5xoqplR+t0YiwB92PK7oIOUMCKhAH3JSon6eERbplwWaXdgGWh9b3
lqAEsjFf4yVMpmZ/NyeQMxO+suFRKD+j8RggIfkrktfX/OPxbIyzD3SE3CQ/w77Xbo4AYCF+eiQ5
N7rfVtcGNC8oYXy2hrBsoDKLDS19uxXxCFUynb6jKNDfG9cvq5uxBsR98SMmXWNWy0R3Q1FMwUV9
1oLIG70h88N8tPYT6hXjNMMb84gVKMAEtorMowmRwYcwfGt7F28M3+YsC5rxjf/Tmc5dNDU4Y3xP
H9whxUhd8KqVy6M2PnJptRWfHhMbkm/SdHKuynrSlABs4Okg5diqqcUDqDd1rsYgBr0J/nIyhYg4
iUVLIMZ5Pu+Qr1WEHwFYZFQsluWidF8GPQ9R/HqoQy6JWeI2GbzSHMCKpaUVbS8BeSx7Br/CWYPN
1Acic7bXuagPb0ETSRautfFVoLuLxCqb+Szp+EZuf4ft0OA8WM0OwyzpvtpQnBmBqJN6So25hOdG
Iyc5QIcFIp6rmyw5SCvScDnSS5dCVLl+lwVnduM+9hvr9sXY2wIy16Fsj4XL8ace3P2U5DPtsavC
SRqRMA4wFQmXXy29aO7KihlYzH33VN4SV21xj9JmC1syKNS5lAeKA9KKIHEwAC62/XypI7PmgnFx
y4VUvRlYKfnIZM7B9YYLQAwAdL+Y9gimdojZyXxRKqs/n7JPnWJise7ux0zH2e7N02f4yrSAo4i/
0yD6GCnEfE4QKCBO01QJ3ieIPIms4VjJztS0Ji5vLl8QQafUMH4OF2qzSFFk31Uaebd39JLO0Y6f
YWo457bATp8WCwp1lQbiXEbwoiq6HwFDYtEzbg013O0NJal2KGcXiblRrZMOEdXl7XqhiHyGhF3+
QMf66P1F6dooDRFWd7O5XpFFRgxF+Wus594O/m2wPF8RRuAaYfba2iTfezmiDcjyepL2bP6EMNCz
Ir7nzq/nq5NJMLmBg8f3d+Surxlj4gNTC+mXYnOxpjv/CTmYzgNghMFo6u+5TZAzK9J2645LXWwg
s4Lq15vfKQE34mY6/1uil08HUgPZAtMU6XecqLCop1HFSXJ10kcda+UM6r5EGJuOENLmxG3y3uF3
J8W9qZfvja1tWO21/N/Ysm93cnG155ptU9RFC/jxTMZLm8VJ1u7Cgg63nGXQZfXASoJrGNU6KPyr
41aiJ02hpOfLAInkU8AyIAbgxdllR9tm6ERcTDfRuR35hO2q/i42aWJ7lIwaPyMa8s+xSoCuwxd4
i6yBwnJ8M5MBK2baIp43BXcXzp6tixxVadMzeh4TPdd5NlpYVMA/mvfg8Eqrnyjoc4S6V/beJRGM
LfsccflJfXCfutcIO19YBa3svSySlCkU1AGZ8l0AwJ8mBTQmXV2Y/tE0dPIxP+Vv+q9kPa4jeciF
NfQ/tRWf3PSet019NkccPs6LSVdSGsSKKoEZjRWyDGdB08z9hX3ZsBEQSgdhEDxJgCp2m0KHH+ld
PtEbyQyiF48w9bFMOMKxjh0EvEcysCgOxv/EiKYW1o6A73urjUI88fSWNbKJyorSWltx+8xpk6Ef
0RMSRyel67JmH9GvErgwqgkBt0W8KHOw9nXn/lukXSXBMw/TGw84urxJ5BbuxclKzABKe4bve56V
PPAFfySTY0XCg+tQrjptXzWPJaaJlExybasarQexL8VVjqzbVcVbHFWpm/D0bXRnS3p9zJIcgruN
uGxVgEMVvYMtwzH8rq4ItMnPnHGvQI0VBtWMfBOwKnzDrzvvEimK6pGhHCrF/IPkwIXOLuavQbBr
G9nsKohMO6gXmu6dL147kMUIJ4ez5+951E8n0yzrx1rRWmTeSchw7LUztjzuyed9MFIERz+lzWOy
yCnEwqRT0HOcvQxO3t32S/LTWdqPBjTwzwdZaIcv6mlifRTU3rv+do3WA2tJATjeznw7JdA1uDQA
lGKDmTH31Sx1UF0lB6vInMG2JCe51EeI2ANuBnkKE9bAfdZHooIV5vG1uazOlQbyJR4q2OrKGryP
v4QvOTAMmzzi4pglz2wYJwbMGfHO9dUyNMml/aafR+Zzq1rpEGCZ7IfvKOVY+89CIskSN/sNlwut
FfZ1ANiCgyqNf/q0oiYKsFmNyB8zHy3rThHgqzLS/m69DhOioTD0f5H+/ax32m5JRVZkNEz68RVu
GqE1ZNNnX1KtiVLrAqann0PC/Jq+AcKqBXlMWOodvJ8iraqoC8EHUDq0ihQirXMXXuibQ11t6o7w
ATQCP/Zi+2Psf9XBHMNiUpAijRh2PQATtu5DDJqaSaimOj8dCAn8ZPdqyAyV7QITHGvXOioHbA84
SfT6PpW8TWmQvC6Xoz9QzpwL9zjci6bR1KsoNCuqIS+UvkrbUZ2REqH5YbB0uAw/33GQ/Es3fmZa
9stglVHdN758myUXV6HA9VC6cqGy6SNvo7DvLbgNAhmaLoLy2WVF1OmPb8n54womNRx22Ga3ZB0Y
onOwgelaJ5JqMprVdWRUGiHzcSRGcJMVjiQU3LrEeXxo9+PB266OPok3rqd1wCyOEmW/NqokolfD
2IPeriPEuT+piDyJXBgA96J96fmBGY2lvj1TUD22c5MFgO6echJwBqx5cbQMAsdFlejNnO1TXINx
Oiiip9ZeaUqWglrWpG4+7a5WF0jff7mccZisG+RHTFQxUM9eWdpjykI4YhKrwfb/SGhHQGb+57Q1
AyVVfcOBJlyEfwavc6GPUxFs8R06I9EgM7XEqnjGoNk1ymbMnk1o19qnEUrLighF3zvj1AN4k9uE
ol40Z1JSLM6j3GwaZt3zNQs40LEZZj3aypF/mlXYG0K/NMZhjdk80ZyFWyhfoCWL2tRSIPjzVMyx
UykYOUpnWiyL4M8tL9jW/FcwAnAyBjzWKLadD76R/qf3pWm8JZdGd+uzLGueUVPEMwWyVaofJIIF
B83NMdroDAG5bzrhlnPu5yTLZcXZbxPKnxrRy+87uuLw2sjlwaqh9WWf8ga4BISD/SYxEA0hbcP5
9NMaw3uoMe0SGIe78N1ydhhptN1tKqXQQJhLOAmtQ2eIGr3XfnuXOW5KsvDnlBPf/CgZJ7tkwSGn
5ceJg9UieUbTHsddC0aMmuCLCKiNkMp93F1h10/X7iZvdKgIRWe2Q04jHULVrugpLtL+CsJ8hXda
BdRzasVmUV+WtAcBbkIfbAMD2AcpgqhbsIPKYLFjnNX3m14j3rmU4G5u3h63Fnz9q9UFmupw0IYi
SSg0wSjlg2EADDKEYgSO4WlaLJMynUkE93Kn8ZUjPJWFyxOZXKoNqc7HxLwQq8DJL/fRdGxa8nVX
DVyLNdUDGJFrOuSeFwTj9FZjo7WQHTQwv1vp0q9e5XG3rUUjOpbioFdflI0rS3MCbTXLhhSwcY6q
t+9BqUjpGHD9Xebou8X2Y51dvgyK0TQuXSQQa+m6drfINU5Taf5oTxUAMLGZm1M1zY7yoMyJY6qx
mP4d5COcVBtSsq+zaryOsRC6pvhGYYVGCGf3tzIHs76WjOfkiSDr6DC4NFwytPgOYg2jO2IhEUIS
Mvgi22jYhoYKT/yoOicIdGhODfkTqIDkgX2jUIwwlhp/oX/JzC/w57TjRmL3yxJhqms2HnRzHVdr
dCzmVRws2VgGCRzfxQC0qeSio4pg84Q8K/VesFV9Ghda27T13hN45I0ebYfvl59T0gy+F8ZQzaq0
ZSPjU6GjGTK/HDP/j7An7yHx744ZMeqBQ6CKKdC09N78M9Po/ghrwjkGbG9fr9bSdsq07CNuhJpW
IPO+lrias6DUbiCf0JBOmGa4oUV3t0Mw2lbx4wtWB37Oyczbdu9jaIz8T/4HBlpFx/gwKgWnGjqr
vMx9qXYvXHVCCVg3YmgTgamV4irY/ruXCrbBkL38aTYTyheSfB/fdkgSmz/gTYfdqsbnOGqr/5xu
OykhAgtnPoM7c6WUaM5sIoW/56T7grf9SlqI0TaU70nAfiKkGHLnowvQpRef0jbg2XpsVxIup8lF
/OEo7do5a5uS/i8VMNDiwISC9AFhvVMVuIv2ORDID1eoPfAkdbyeUIYzqx4EylvyqRq9f3/EPyd2
yhCnzfaMQbt8BtRGvXcEJbFeWXBr3BpeSgHoaD8LP12p6wMA+nmBWmo46ZrQhKxe4x/cBk0qTJR/
FZscvG0esXIy8qWykX547nHF6YcLoUbqNFrSDok9T2yiUnlCrKhvuaH1UNCoSS8KQhhFmuzj+dtx
JkNYDzrXfFhI4yN20+ew5uVVpC786DE4Tvco4abeoLhRdp7qatcOlH8jgMGP25UtQmRqIm5aEqGP
RoAQTu9+PI1wqODmIBCOTvhg4xFfWytiOyFI0sJktH9olBaLUBTvkdLZbP0b+ZV+PXdueb0=
`protect end_protected
