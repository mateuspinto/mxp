`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2160)
`protect data_block
jEWNDSf86hwqtKqGxGzHWLIwUyQ8Mv2FDXbADKatwIxucWhtmrct5lGQd3vo3tPo9CIwLe3DAbWc
QOjh0SAMep1Ev80etFldVkamG++uyT3a/OsisHBqZA9JETk4nUxJaXnuPnp5sKdkfMP/f5gvlUNR
7vW5ck5NLjeGNuFoCwGt4suqadV/ozBQ4xQqXU80d20PAT/+FBrorGneYkkoS3rhiHgrtUvE26oK
S0622bfHdBHK9XKwODhcMChkEre3woF6Nzthj0yoo962V+m/ugj9MahzdG1U1hbahszBnv1HhJFP
NkGc7lkh7GkT1G6/CGnBYm/69vUypX6OsQTOJz6JuVYmaPmGyBsrgSh6JyyJ/BiFvjRWAoO03Otz
+L7RxQKfoPSZDCEihfozE09FwzgaljDMosEP1htIVo5zqWEUO0k0YwzcYhZifvawZwTpMcJC+Nd4
KONylu3ACWSP0nQWuqEka68/3i1f7C+GbaL+j+0JkXCEMfu12TLk4CuzloNZkWfWRwYt5xPTaIJp
4Ciowv/JG6rstNLLgAOajS6KVqtavElDugpZnZIbxJW6S1fgNLQU4RL1f+h61Vol2i2A++tCig67
qQLn5NOp9ZzgHa9kFB+jzOhkXZ5aPOiSX38tPZboke86me9fbU4WrX1WsHdED5jKvx5K6DmxUUMV
nT04xMbgG4mKWE0A+OJXwBzk+4poNqkR8EkejZxJsQHipHlSEfmHUXJ9nujup0zuTH7uGzYdWYij
ezHeFPSmB0USNLqxQYE9J4WKv7SNV2Fiogan0KRJrbhelHfgvp5Gz5eXVFS/Fa3D02Eqj5o/FmX4
6UmXjGwwAca4w0tkhJw8y6bfQKH3UgCMM2xjm1IeHIqM2Fz2KbiukXuG1MRWJ24WAPw2JPZtYhpz
1I/Hkk8GhbkFksiwcxhRCUAGwtwiHSocO86VUOZLWAOOAXtLvYMLB+w7AdCasIomhK8tK7jhu+yV
XHffQjLf1T4LBdpXCwY0yi31f1ekEKTGLfGG8uLes5nfoCbbZlVCCETLBmbSmINjhunGCr0xHl1U
JBIxb8CaSZm77Uey/CWGEhAZ7hrcDTh0XjFVH+UzKeKP85Sirmkz0kdZ1cumgipeUgk01BGIe+DG
R6Q+Wi8SlGg1tRD+ihM1uP1v7eKqldhkYGrtcYNyI02VzG1ZWDroHUXr/QdT8AflIDM1K5D86gF/
pubaB0wmPwWJz4whLL04RAQX+fMcvbXRYtHOeQqjk6thooDpBAnqr6TUYPH4lsKMyfsUmDP1jX1R
yMPaUFdhblJRS0UEdlcJGMOC4L+LPPySSzRdN1lzJpTN1eIsHJaj1uKnUFg6ow1TH+Id4EocH5BK
8P5w+P62Y6agowHrnlBTn775ugGgspbCz7JvkyvfDgpYJDRgOAkqVQxRUgkUjvXfGAMXfmyK104A
WWByNSp1kcn1JyBjFZfd2MNuB7Fptv7wWlGnbJjMviyG3a2GqOMCtyH/pWG8jG+Exx8jWBA1BnH0
A2BDbNf2+Bnsg7tny3Cv0VWgo7meSVgKe6Ut8D/UI0bnPT7EzQsVcC/P6u6p4FrPonEsOTl2hNr6
v75Go/gFyEIAZ7gmdACvYn4Tr+s4sSfNeSCdPQSeAnctirvM1qQTxldHCBk+tlbzjcXu4SzNX/2Q
ji5LRgFSn6yFcFo+/xyjx3KHtWRVNuhBdeYAaE8DymxNWVZtIF+QLV6p01B1RQfDOaBcFnFCkoXg
gZSVHWomzkLsFX3XZVl3XR19iC51mSx6y8ZqPTZHCph/oMb+9ZrM7JjQTd1JitIcSF8/CAn2T78v
eCQL1+tVzU4hWud5G13hSAPJujzXEJtqo2ZkLX0v8bDA0dTlzFvHTrxZBKDd1PSBgyF91GCTKEKN
973atGLBz57LBEACgIVyx570kGYh8Zftfhw1Z080LagnRDymVUIvstRyThICx9uuKKmRLNY1yJz6
G0pnJOi7CYgkvlsbnf6i18OQfLhLrr2pUoUUStw2KB3x16bbb/m1po0m6w8WpDl9l7gwiacG8/J+
gTBAL7poqSSgls07SpTNQn1sPqqJNJr2jQpjWmr54c4zho9dXj2vvbqCEkWSZ8TsIB1eaQRsk3EG
fonEiZku9Gpsy3oQvEBxZKZd+Y2O1OTSzt6C463l3naR+0VQDL/ISO1rCkQ1NaH/CShVetyYRbwr
N8q7ie/iKm4kyBfL/Ye5+Xa7jBvhYsFIcdgddApxOeW6PZRtT09njHCP/CtVKq4+VZ8upvZ1c7ZE
Xpt598rFdDwUV0vJUwKyH9VaUv0O94lQYBOJKjrNVtFEUta4EWRWRonu1mAXE0+UI+TCN6rV1fSS
iCdXHkQUQBpbDjGAFeHCyBrFMk/ghzcbHmxIcIPEcu1oykVCU4UJgXvarVHkkzmHpWqpAH1Q4UH7
P1bjKZ1ClxZzNk7DNh16PmtyiVZN594YKSI51uuCEiGmW/BHaXIPdniNNk7C4ia8AcpcXXTzFXLf
6k7ndKiJniIiMrYobURPalBckxzCyCmLHtTJDuXHhsHvhPY7CwgM1yluv+oS81NY9ID6mE7nd6YH
3MDB+llDvgVMKrgRaSE3LxKiWRBARgg5mXozMFHZzDMtwFZZQiIqVo0/G1LVDCj6s0yaJ23wEXkn
njLHf10ekk1WpqVarHM+JSHQ2GYDl8HhqL3h4QXk0TuXCxsKy5l/a2Ck3Y3zmsWHoi+2R80llbpm
p24M9VvnOECkCcrr8XTQkvmtGQshIDnjGDaQ94I6uDPpihQ5XM/d7DSvESHsWqYTmtRcBRVqe1yf
yVRMOdUrnHkjyXM32ZEIDpcpWBbREWjxAIEGiiH2r2pzK8RIaR8Ojwmlm9lr8oC9anoT
`protect end_protected
