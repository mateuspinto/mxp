XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����QR,��Vq��6���#b��m�1�,���T�S#�(�ҥ��^�N㜡�r��5G����W��2�F�dS������^.zP�s;�@n,�$Iz+���ãʜ2]Q�Us�xj��l&{j�̵���D���<wN:5��Se;4}���'�*�`@&5�({����QXH �OU^7p��G��a�C䓤�! '�cΩ���p�{��c�A%W�� $'E	@g?�>Y��U��`x�_4��N�6�yE�ǰ�mb;#AmF#g!��C�J�U��qK���
�+B�R��w���G�9�HWzCQ��7[q��ϒ����jڲ�9��/��o:7�OvߡA���B����!�g��ـ��E�N�"�I�˺|Zj@�P��]o�BP����\n�i��2����cN� �٘������Z�X��Na9`��NH ��ܠ@�P�)�s9���)Җ�֋=�hs�D�&8�w�9#M�lU��N���2oc���"2�����9��,�yv������h"-9m���(0�Y�~/������W�Eg��w��Jߋ�~��-0#�y��r.H� �@>�/�A��R�DR#O`�1
��qQE�d����>/ŝW�re��g���ҟf�T��ٓ�7�eW濥���)~G���;n�4Ս�[d�׬�Oy�6Bߩrmq6�#<Qi>'� ���������o�jJ�"��n	`�˜��#kr���7�XZ��Ԋ`�C@ �:����1�< ��`^G���8ՍjA�:3`TXlxVHYEB     400     1c0'��y�Oq�n��L�;{��VoF'���V$Zs�,�r��}��F.�O��Wݳx�q���!�q5Md�Z�a?o?Oe���s�X$�G9����j��+;�^�u�p�Mw �--�Z$���jJ`d���i�#��\��H(JY��A������GI� ���L��1ٌ���l)M,�>����LGs��P�R_�[�m�ݙw����tw~=��W�E|�)� L\R8e�L�ɻ'r�Vj"A�Zb!�DU!�zh���Kz}���J<ս[z��:�%SY����8*��VE�բf�3&�d05O{QN�*���W��4*l|�V����
ʒ�q!x$O+��m��P��+�!!�mGgЇ��)crg�}~E��s�o� 7'·"}��3)ңw8��A�U�Aq��{��^��g���^���(3��&OJWuI�b����XlxVHYEB     212      d0I/�!��x�k'���;C�q2Q��\E��^���� e�[_�m�m�YzOwJP�t�T������������s\�q�ۉA
��H��At�D�s�!�xKm�u�x{�XK�l���n=6~R�)�7c���"x�x���(��܋7�k�j��A'%w��0�;�n/�駟s��ط�29��U�[�bmO���;vf7sH`y�� ��