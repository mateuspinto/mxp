`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
tZ8rbzGu6dq5saYLHTP66sSq0FWmIFgKRskjzm5Pb4874PLeqC0kMR48RJ7ZX+8ZlQqZCeAGn3jM
QkKRc33M8Hdz7d9L5KUDH65R4Y3XuBjG2jzbDaO9OTLUwk8IcD2bcfWUzMfdMWP2E0w6LwoRb86i
xTrdMIMBl9xJ2ZZkONRilGBHyWYvhAaHfggA5hYkPzBuo30m94w84d/DssJXE4Z7SWjhpF6DD+if
mS1Z8Tyvr6nplApB9sw8dEdBOayD7VQQQN5OhUz2D6zVldn0QXJigBStypMAWGHEBf4CAu/8WrpB
240oaZEcy/i8/TNWxipJ+R2T95jQ1baNm0M9Gg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="nrVSdoB4OihRv0Y6yHVZp53UFQMKMccNoXm8PPX2yIU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18064)
`protect data_block
73m6Pp+0gtl6WPgsPQZU/tZopaSDW3hjiYYb8Bccp4rsnAcvnTDRSq/EBywL6e4gg69Eb2c742yT
EBiDNPDcm3VlHffxXjJD7ULhAnwxTOVVxQZlevF+zD5MzRhU9UDM2tsmG2Wf0iLcWpG0ZxZWsRGT
j07JDC40Qi900LxcecCKsZ3/POkAbR3/5wHLyRjpt4fdSxp+IC7xc50t9f33zXilJH52ZHtAxcHy
Dzh0wj2KlDxqUv6GnMYTwfK/55Xqq4IBCHWn5qA2o3dQsbgpmXEHlevgg1NFLmZOM6Res/3LSCk3
1pBtavqQ/QZf8S1VQgo94UR9J/trQbdqzjZO2kvppTSwCAV1GMWCK11cRRBIwpYAvR0r7D1VlsNA
DV0RiNYo0VRGw2quAdT9VDwueWTcfiTQ1UAkgRv0FpxDapiOLNnTdU2az6kFwUeXIUI12zG49xp7
kO0pt058WyG4jTHg2x5kqP0zAVs/R6dYg4YHxUnk2ctue89Q+FJJf+4d+MBMlGRDfHHA/nL3fJk6
2HCzWX7hxTNtApDijJYql08QG6nIDzqd3mz/O3IDJVOsasF1sB0DQGzkW/n/8Ilz5jPc4az2rtgF
dQgO/lawhbg5D7JHFrrUYvf4Dipq3polV82XDzqpmIHQf8sVRoSEuoL1Rg7ocehixe2Kib5mi2AE
zy9JLCOfxBO87BxPxCKG7YQ1pyT0HKe7FJI1Ih5rkOukTZK0vLHQwzh+XYklafrwCv1AN3ADcBPR
r9rqT8h+Te35EJAIxiIZD0/OMlsMwNnMNWcXB5f96IpXqxojNmLzCZ+vJe0A6UlHF5BbevFjHVOQ
edv0e4t6xojp/9Mx/iZh4FhVbVwrhwsF8rpbyop8kllaZbeOEVtMgFsezdA1NN3rTH8Lmdc2Kon4
okVOhO7RWjRGl9Wck5QK8ozt8aQ8HMG3scu9tbG3df6pDFDfg90riUndrqozlMrDybQd20PLgZ7m
k5W94k/V8FSZokHXg8eAV5XA3NLi8J0cZhTN0gWhy7e+T0tQDAIqVFPH/AlaBE8ywTGa8mXw3vXn
6SQIetcGUq6GfxzW0xCplPISFjuZtkaefGjmHJj80chBD1zgIhYMxVMNYAcZIjwozbWIwBto42BK
khclEmAVddWDGDv4Mepp/IsPPN6sgmPHBv69MYZAQxaT03O+Fu/kVynyhaK7nYqbTQ8hnKEssxe6
LTLLywlK4K1iNOzdpPxm8v2z9gqmGdueY2/vZYod6W12OTb0AnMBNFyW2Itt+2pnYwv1L1U8YGFj
WNfKXlMWLIjxYgtSdZ0w+jUTuWqmVphO5lw46jVNi3g0zRwNhPzfin7QFDlHw2Y1uvr9y1xOE3+t
cSGljuj0BsvzLEjmjIOcsRDKsilRdAMYUdnQWIsVWTIXSSO/JsGF+yzDuDL4+cHpw9u7hylBLOcJ
0bGnxecUkTp3efm25k0wLze+k9rsrcbbYdXT2dgx54qYb8LsV94CzNODBj31kgfrEDU2D/MncCsg
955hZy8CC+IB8Dkt9S4mjarBJeMsCl0KaaI4U+Ny9OzSQTQnC9LVVTa9Jw35sCPPEXZ8lcqrd0+e
rSqrmh93+PwFSE+t7+UK/C6CeT8ua+KN34tHZxX1lWy2Xb9AI4MjLHTYTkM0A3xI0dhVO/fSSljI
dq6RgoqsaDCNGiNE7Jfh7PurW5zlM//uA/GcJyKFi3qZ601qHO5JnBxQWze75mnABQOFkfhgesBc
LJtFM1aQIb+LSmRbUiO5tEd5r8VTqk6wFCMqfsB/k+dZaKlKyfNZp8L4bzrAYLG2vzpDm3p3/g2p
xoag3Ej1vQP7rCvtNf8AcJX58Pt0myxMkFfc/G2T1bzUSOfgbdwh/uwM/OF94nJMt+LanQ0aVJdb
2SUqf8SDqBLpzDnLInSaJfhvTRTheLGwNZ1NQ4V9uT+lxiTo4rVAE16gghJO5ootylviY9CytQ1u
qqB7GrO4NOH6j8Atsy9SZC5JYgfwnuSjkpfxR1lQhDsoWGsxcQytJae8k6BbNXDDWsVk/wjpAszF
HrVKhHB40Y26WIs0vUVg5+4WRgD/b1MaTwjQaIG/YeHrEqWNnNBnL/I9p953qRhBwsVn5cWB5/6f
tVhBMnMYA6bj7rm/fXo/amZYC98zQ6Uh5Fz156mlAz97UVHCKvpbriTVeoKTplxAZMFxdIE7bVQS
KrFB/CuTqngoa/a0nj+NpiSolvOE29AGcCqCgRTnlLp2S+7CS14kspvhjbzOKzO4kTQYe4IB6eeZ
TYmsF8Uqup5wteZkY8hYeHbBuKVsM6qzrffRamuP/MVqw36rnzCve5NFRq4Mjl36QeihCz0puXmV
JIGvKx5Ul+kpzS18TgJhwEsasbeuTIO3oTnATtBTjEgujauNUUtkA1zyiIJSh1pjrlfYRp/f65HY
uyjcV7p0d7Lr/MuozM4PU1vBOjMsz9Xi8beQcqHGB3k/bTTEogOaGYyQoCceE6v60ao5+e519S6I
gXhKIRvudneKjI+9O+QA/OyBLAVc6WS/zNiogdjhBfWUm2DCFiY3UZ4o152bGo8y3VsX0RDKfz4Z
Mmc/2W0mYJbnyaJFBNzENN/vb9r4msyIy3gQXqTyF+YrJ2jgy846CDKAHOSSe4F0msViKKdQF8NQ
ebIBVtLscohAhXtWzKpnuAVmYAwsQ9mZIdFxkevnpjtR8AdHJWT9viqSGNYoFBDS5h/6Epenpurs
wXZq11pJO6jgAA9wFX+sgpQkELjDxi1GyhQM7sQSxpHQXvGIFoajwaSf1IaLBONl8cKG2J+JeIgK
BjqM+Warj4YQvPdYqNJva/Wl5Wkv42YaEPRJpbqz6PRlAbru4C3YpE/wtR62JSh72GPppE8lhYto
7+YIfD8FY9CJTtYU70UHkgkFbwgxhGpJaGRXuLCH2/w++NCYNDVsJdHbWsA0eeutQ3k6PKVlUz6f
BWmAewTD2CazZ6Y/mAOvgQ1rK3Bjk1w1yXePso4NPayoU/G+U6dkBiiswHPduz87RY4OxgNUS/81
hDlCcNG565zJcG+MGRw5SK63B8Y87P1GhM1ljIM1BQgd7x5w4/3LYHWEI9D7MnArhTvZG8NKfOWT
qsMvlYzDQEBSXGUfSSX+6sJMIZimNOjxhRAdD/mtQen62z9mDu1mLKE3BXERCLxcjf97OOVd+cxa
f9FcfqAuVinXmiNkF3oqkvZ4Qej4Y47Lk++HTxVv35rgVyVK+W7QFqqxGG/Acm0y8SI2Do3F2iV9
SVRZBpy24Nvt7AsGt+VjGw8i/oOAzWuM86c6hWyLOww7oXynMSX3j6wSaNrxV7EhpaKMbWCKs0Tg
LGfc3NWQN0kI6LNLM9+Ap2Purasq2ZpqyU5YCvOAEC3cjB95lHSP5SpKBxY4GnoREc26eeVnq0Ox
SY4ve4hsvKkneJXEcnB98y52cxlMgWineR3ohSgzkxyuJMfmFtuaX/6onHOO5j5YOQG+STYWj9+i
kbH6NNd8NDKH8WLdw4pHlbtvzQpMohYT5PLHjNhKmvvekZn8luTYgF45uPTbAa7uR0UjDi+KU5FB
Usr+0rtzqRb7VOzt2vGoOaCo6jXKbyKVc3puWF8bscW+NNWUoGuUX22MAfwF3avu24lt8Pk/lddt
eH05l+rcA6NSENOOsqAOLdXdukmFucC7GTkmANzLvkw6Zn5QE42SJkxiQP9DWUpjvkIk4htaiG69
AgCSUyLVuRwSpeeI1+9ZOxI6A8aZ1vd6aV4ib8iCqyj3a4ENI3309xbuorY5WgKpDcwgCeunGK3a
2Dux7wOWJ3wJ097wK9kpm1SDoYtdgM58OImVvJFVNH+M/rimFEc6pnleXmtyQ2JChGSFqMZnPquO
AS97Wb2VMBy/jrlMqew14N0Av00gS+Gdt8mIv7GY5YcXm3iD4DpStYvDZHNbFTe+k2DjNogEbbvO
zq+6B0WcG6zeiYxG7yJJdjCFXWsritBCO8DxO8Tmq7kJIIEnR7Wx6Hjj7GLuoVBAtEJFQofCnWgt
i+NIRSPETBf3wCfOKrYkE7DNr/sis3+xC/r9q0wLEwoASSZxWVdpPX93jUHMlp6eK0es+bmIroAU
rXquMVUZm2UEoVbXWZ1Zo6xyNHEnaV9wmsm58aDByE/hhMC+4wdug/bRkAAQjpfV1IuTWRYpzuSn
LPSsLyxL6TskJyh51V/lCpbNNdAI6guMYpJSRTfs+s1OoWR82ks7DAT6Ixk6i7K7DuiVLXVfCzAV
1gHf0+x3hNNJcLctVhnxczoHkAgUSYh7pPA45vMHu4phbSFpUi83LT5/l1aIj5XzUbbhYtEuu4mV
u5LjeDbGlV7Elq6nkQ7yKcZFi2jdYHzVT+NeCMVyTJcMViMcddf5gwtVXPNK5TdIPJI8MsW5vY83
Wl/lgiBUFWJvZEOIZiJiYfIyzYBnfrHXh2IDXH1D3/cC8cx8CPXuLB50+yUXlXHaKFO7ExvsGalO
cJofZ9QlPVzVeSgFit+x4TRY80Kc55aMRvcZMxXJCV5MH1HFw0NpX2sO74sXhxcgkbceiSj/hgkr
1dlwWfp6iSBXCHJJDA5JmANTK7OmqoDP0eB7cFjYKaEHvwNxeB2BYTPe28G9KYFYD9e73NR2ZwxP
0i+WCCq9fwbj02jXhGnzOsqhjttAU8mQcktm3fHgSnE3NoOJGYIt6HCBYovLLIr36MNG1nQo/k0Q
C/FLcMnuRNTlgsjRVIDz46An5+ei8H3cP5/G4YZkpB6aFsOSE277TeFdm2V5Z5pv72ZQ9j9+5Tt0
MDqRYWaYDqkb521353c3u2j708XNrvKmQp2gnJNMY6TQplmxx5SFNvT2ELwdk+3hwGWWvdCWGo7s
wNoDMvEWIzSNzRX2nBObj5a3XWKtRdhUMTOr4PvxEL80vZ2U8GxfI3kuuDercmZYNvsBbCUTRxYu
Nmschr4+Dhmu5/RWHvCAMTIJDMrQdtqiZFt7hgmTNWXXJASOeUw7LSW9xlXCCqlWKWJxJYCWevSJ
5S3dQeewz7Ire8ehVoMhu4ajD+t4N53iYJ8Zak0PIvFf3dpJMgqguBmm4yP39pVsQFIR721kEQOZ
ECGRjIXye8Jj3rXyUP3y+orlN4KOF/y3n+HYbh4CjLK7EbKsRg7H7B5z3EvzMatwr2wTexmc0r0p
qiUQQjc08QxR1soxOEk5OUUb8qFcEmu/L2HVH20AP0zp5K4Klith4XyJP3WjX82EApuKiQerBx2Z
yKkbWheht6CgP8OzJCDXRok+JzFL9V3PoKup554WJhX3pPIwvmzuMQ+jmzyy0rJzD/cxOoa919lw
FjSeTwUcIgdAx/fYIchCG0/jVxYGuT4GAlYOa945T4hQYTv/kI4QiM6LkN3HdQd30rliFQYX56BK
va5qqpR9tZOgfCJVKWzcXAYkTFf68oEki/zbKzfRveDt4QLyrcHb60o6+2Q6JjgvmULjyqVaabIA
AQm9kg+dE/m60JSe8dkiGVNez+A8Vl6SpkwT5x8XH6Ubkw0ZqBHtvTD649tHrkYQRbe3txs7DITP
2uolVSAGSh94saFDwZ6OFZCpSDgz1ZSPHu/kbW0ZAJK18i/M4vc/eylioCrY5Yjoad64hxXo77bJ
vY6o3ihW3Y8YsYLIhh+/DwCPdLUprW7e97p4uAeMRDL0CczgD8qVprbFrlglnsoY+A2BE96/Yki6
X6fhWbtUhTipCbOCVgTtU/+ZhL6EP780MlsOP+DqF3e/E0Cl427SspxE0/AUm9ZH+SgGanhxgScH
MMv9TtCPoqiDT5Vji98aZ0d3591rcHWah5RfjG9mPbDNjgcNDTJ5um/6cT7IcG/OFB/0o3/AP2Ku
gqFR1yqB2uEUVIw5UgjTxL6eruSD3eWfz6YwQL5AEmfK0jg+lwi32hExgrv5hBWYCwLk4vbFyuKl
vXW8hU7GObAGsh4ECGb4/SZybEK3FhUuteK6z8EdDDmrq9bnyVdbwVgBLGcQGwX/9nn0jOsDH9se
bI5bjP+qihX1yvfmQKiiC7wv/quyX2FD4xOqDFXc75KuSYW/sbH2BruXL75SbSgqcFyOcRa/ELw3
2odczzONNTaKbpAOSsllbDg0ThOUN3xaad5LwnrNJYdtr8OpxRgHumEHs9V8kxTsMeNiF+32SYCW
pWmlN59D2YuLWd8Y6tSLS4DErbNjn+anojsDaKFvlf7XvUS5zfJEfL/dJF8z9J7iU/S+icF2swka
cwkw/Q3O70/srTQu5NZv2o6EHng34kGiylDN9yWSF3k6MHKSC68X847h6NW54CM/K/w3ZEwvYB70
xqrKvJ6tJ3TTncIL61Dh2oA0L7gEOmzF2zkieFNwxSQxEut/03rlXNqGDB9fhr14JYJnbdx631KK
DbZEY0XJfuojQkZXCfDZCxpPXUPIypeY4N+L5mTRQVmoGxay8xDvJDXlb9UkkieBZ8J6tEoXh6Mp
1CifofoWiUMsVv8JfY0RjvMsnsG59Ky0M+lLDww6n8eMU3p1FWjNvlCjcl9N+c1UGvQy2oFbUkOX
Esg4FtXXdM0ODAk02X59cZWDqukVIy7fXNKqMPBQ5hmv1n3DRlomNYaNl73PruYgicIEbv1N5LTk
h1ET3BhUefBUm/Iq90vS63pGto/2bf3qhIqDMyNfg11QGKGHoN/hyJWbi+Hb4ilS2h/OZa7YApPV
IfSh2t4QUgOw2rwrvYNLftPcFS7UiiOZ2lABkGhhKDda+jgNSKzZbiUdR5jJ5le/SgHA2UeUlD4Y
iGiQckF9jxw8dcMR6+ZP4dvCplgPbAAR8rhm/wAcNQ5DMPFt5Qext5Su4eUBy2nJJZeg9tq+XK5K
LPz/xYieiOX5QGPOlFCHucLzBfbA2OpUxvCbM+7A3hoS3wyqgToEv+O5y4gr/3xyRYB2AsXWByKJ
9EMl70IDTqOcQ8KCSBJczAL+0ZF68HJtmWvmledc6lNFYHjY6AW3axiqEhisbTLtUNUi2+0pVlB9
X1Gu7xvE5NoyJ27moWRSqtPfsQQv5Qrd/R1QMWLqzLwyaKh3gCNFVg8J5TfhBsfiQPsgV7lJKGIG
lv1l1Kwi5TN+MVbCspGng87E0u/RIeCItJfpgobMNEIgtrbW1j1vB5/SXQIJzPK6fG9NPhxxrqFk
STTev/OHNWrRh2Y3jH0Q7pt0zJ0yhFH7VsnILyPziWXHzTvuOB7IkuDDA5sDfqpETcyLP4NESOco
FnHJ7zY1jRcXXwhd8tKCaOz5UICTPKxflhSaijv2I+SVF2Qycm5fUSlwqp9fGf44BcIPosWRWoD9
Akq7sDjUlM119/XMBFq6m58cPjQ6saW7jf/e6J7yhxU02hAcHoaNeDJUIhH3iA5HloVYd/j0nOIJ
fgQHxMHMfX1ZgxOZHl2WZLgntobypzvqJEXPY0w4KL49KlkjUWszWIphNa8upICVApVOGgF6w58f
347tQrcJBLRlf/MmaNPg2L9TbcLKQTqmyjg+2At26Aqg7R96zclVNF5Nh/omvPuOKT0ROLYQnIgm
aV3HivsGo4SLsMnDzVg0tr2cH8GSAUZ5JZ+2dSYIsJkbLkpwtte6JgOLuoUNguzh+9yEbM8tmdBk
1YoJmkaP9qYCKNcx4YyxWKz7Uz6BB6yOvXqM3WePdKYRK1jtC3tkTdvR1SZRMq0LMByxkV7ORVBw
znXLcE9Ez8J7HopHTakxIuuW2la0Whsr4vo6ramcM5FIUY9QBraFqhKo7BLXO2hhBcCJqvJBsYd/
Q/D1buU9t6jFCXiOYw89tu1rlN5VtcTSBo285NY4ZLqiuadMTEcxdQaCS/yKwyIN6cP7JIHBAbys
ryk8nCV0qZv0w0kiF2k3HKV6dxpWzd+EP+aDJ7oUOK1mKHzJlrMB14PQfmXdRXdXF/NgMNtOSj4M
+rJTkDBW51wS37Qs8UCJciFFmbFx1MTey9n2eet9qkyPLlXT09cd5gaHoi6sSLAtAinMd7c/8wqk
1EFsMxn38iqkELjVgswH7CaGSdIbdGVqYU/NHPROp1nborefqNjwKydb2HFS59Y4S4wToQ8iW5fF
ZZlRnmw2rJcW1hSDZZM5HilDDN5r34IHBa7KAWaY4p/t0RKwZ8BXE7Bk/kwjKB9BfaSGGxVBo7QU
F5oIWWf6z2hGTCxvTS26sW2n2MuRhDDFvAH1jaHp4Uy76/lTKtKqX/a9K6uh9nCqz+GagVfp2xkA
ZTNDLPCc5yFeaGIxvYLlP6unyOqtBA8OVSrVXl56WgGQbPiEf4+kAEGOHUiwxjYU0a5JW2uSWaeD
Cpc415A3RocP/MYzFeujGeSvPOpKrwLzwO87mdloyuvCKJG1nf1PrfFe2WFOPtJX5S05A+HRsltT
9GUdQOE2QXk8bIaEAutWLJpIiRI7QNc/sCW3FZ1I58oOjYM2K/AjaWsZ2Vrx1J+pocHsxWZC2Lh+
oq+qeIOA39dYvA8c0SdDEkmXx4g5LshjwGxcI9S3xfgTiI0dAUQakPXr42g1g8f3pVPJK8Jk7pFk
MsueTThRpasims9F7ccqQ7IIB77FlIC2cXu/znOnjK07IFtXnZAF7SV9qJuGjKl/p+hG5UIkH/AT
sNKtTGZiw25FH/f81lV93jKSUZCB/pW6KY3Ya6vZQtsypqpQ0TTlTuzzYmiESPgcU/kIfeXVnre3
GWsXc6n7+3tz0uE88D+Lvdb8/IpPu4gx/bFOxZBWofX7byoi4o/I7pCHpULC9+rHTloKfqI3wNxW
5tkgeJjHwNSit++cMSgne8HDIdnTvqGSChnPl73N7XPkKC9V/pm5Nn2IB3QJM/fs5Fk6oZ2GjaU5
d8UhMgYiLTKVf3kkxJpVVA+1fvocHQPn+BQd/Sqs/BSpLuj0aIoF0HNK52fpy8nU/lP5oCcRvycm
o7VjSMS8fnS2Z0H36frdZOKZUe1r+IU0uHhWn3qrkFaAuRRb0YIlnVterA3MnzBuNEaod2RxMLwX
j6+bwWVXUPH+SiDXqzgAjllv4hOwfGfnP2y/79a//+qBWM4iulWgA/crVSTo69yNV4KxvFqQ3wHS
0ERU1VTM4ryys3USTNmT8hShIzjR6A/B6dyPU56tr8jHNqmsd7HK5X0rhv9hGEh/KtpVKKlJynB/
ahZfETirfdFTk/5FLHR31k0vb/7aqD5dsZwSHOnma8pHF6hCFsXb74MZ1GAw+GFCph6p/zqAvMk4
0hyaSXnlkwHl1KQbQfdt8HGXUI9utDtiIoDll28feMOzihi6vokZFqAEMoHeEbnA0DFx5/1MYsIQ
XD0BCnYNDy6kuYE+rYy4Lf3AFGtKXDpwDwPst12HdYP3RElOBCh4NCpDzjJSzNhHZe2l7tbnf1/A
Vzhx+dkxWjiENJtEyqD27ewiNvzFQVpZoCn6p/empH/fclkigbXDl7OfNdaIYymfkySequcYsle2
iGwJ12MFhDEQ35dpgja7fJcmCfkvtz6VNt1xQUHVtg+bTx3a7dP7+is6cHfBfDkyg2PE8ETSo2eo
spLXOnEU+iLZV4U9CjmbNLPuGA4P4P9FsvCKlHvSiSETkg/b/J2ZHnru8mbuA58TXRzB/ZlD1oSF
fhNSJ6RQxcqcIUDFFPlOKs6MGkuBrCDqw0ODo3Nd+BaWcQmKwHklRXnjbCxZYE863vNLjxkYRTan
SFbuJ2GHr6afMaQDZGeWfv7Nvev7UC2hM24BZWI+TMmtzIeFtVCDoVAdolxVNQVp6BdmjL/pujKW
g4YuxH1jDZl3U3Ec0bP7ngXfWA70x57vCpRUsti1QTSkClFDiztI7zZvuQTiHcfxO3heuX/lxt9h
zNugl0YsA/qrfpuUh78OZ1s35tSQStQ09Yu3gFeL4m/X/yqbA93AjPW9g8hS/wvwB4690vXmbpnq
K5ST1tTCF30MhO26bXAfE+Z4bM5q/f4Dzsqk4yvvtJ6jbEw0b5c/3cDQNvBPcNm5xk19NAMIj3I0
AgRlL2WwU6S6+hIYacG1cP49wHOwmxYRLL/yOQ5OlcaQs4GQ/nuSfqQIGDDTEsBjIutr6sA7gHes
jSO3tN/aDPBd+junlzhcJMp3PjZCdp8pny+dIrSTqlyFRR9U+CVJaDwbPCIRkU/qwe+61/vdXM5k
l2d9FS2FrFZ+VgXO0zQ7tjgqPB7vNv8vtcrCbd5sGJfz1ACf/mntrPa1rd9BHfCswUrh6YSn7ALc
YbAIPxkpIMCK3NXkSekFLE7Noc+I0wn1ifqOFbk+ddyud83TKWfGXTMwhAd62DgzRrTQJe8t2wTg
4uDV5Rg9KxcKKy4aD0nj0dCdP4bPJN2+/2x/4wXakYnXTYMuAtPAL1Id0VMrOHfr0Lg9PYp1fu9G
bJeS5s7SVRMgCfxVeJdiGO05KzBLmJViYLRn+1+Y94UkgehVGUbnYLqXkgLaWwemcSua4vp13Ykd
ro/J8nJJRZxysHlfuLLcAfiXhPqxKP/9cTSeIj8HwncTif5nNb5Udy/zu9YT5GZS7j4VUAKsX2o5
O8dB5XOPgygnFchi1ppCOXuAtbyiI5w1d+Ao7MYKwiTHiuUv83mNHj0MkZ8fvOowiNuB3EoOgxY6
kxYFjT3boOQ/65+C0UWIQyRzUsppd7bBBUSHRW8uJzRO51ltNphhElKqCVMXjOH9E9mu8evOvYbo
yJtP8HaaBZlJHbGjoVSZcLjf4l0vBa7rd8jOZdhfHvDj4qR1Xm+T38GyzZ0kMae3j3Ie76YkbLss
D408Vg7VL07sYZgMDNKp4kJ87uX5i+t09DJLtwWqb9u5EbdTlnJWU56MobRQsRymqu53hxdz/61I
piTl4osi1lIPqZWKyr3MSpBcXkhcCPpWbgcRUFWztblHjgsrh6GRVfCSoV/zI6/+diaF29KJbfUS
ZhYpkMHY5ygPePLaCTWYLLv26RE3+ZbLHP4BlpI0l7vQemKevVlyfNB8H/tMY70FCCyvE4PEsPR0
JbsfzDkyT7cJD04n/ay/lzfTWXYBy5BpzMZe8F5IuVohlM04mHDyItAAik56IxDg/pDE2VANclzV
aVfByNKGWghPokCot+txtc0TQcULsIDgfidxkR5+fHPXJKgtmoGwl6V3n8wK9yqWl+tGL8hM1H7g
trlBoCNAjzg3TW0/IRygpU38O5vSWAqB0QO0QItD1irBAZDlbpHchV9E2sm55PfGbn76adIAEDVa
zsGRBcDQsN1Nf9ZS0z+TH29KK3pMwf5YcQN3StrAVnVnc/FpMs/XwIoIcB7SARcEJ/PN9gmV8fsP
IvjuHHYXs1KWpC8f5+pg6T5GQbEvIqi7Zusm7bpWive/JGWQsPZTfgg2tOGx0rQMac0yetV6Q62L
Yr02qJHzOmMJJuk+5a5+5ia4GpYgKgyBZPyH7NeE69redko0wVAgzjRmyHC+Jq2mg7bYV+szw1+G
vSy9GF+QCfq8DO5FleOjmNRqgBdZ4topp0uDTW/D6nBAPSowCeuBHjocY9pIObkiWdGPE8EUOecf
nQLSTbJaQ1nVNdUm0yCs55a/IuCae8Jnjt2OyJv7bOW8Mw8E0nrG6qFfa7Uor/X2QqvH4izrzoYA
4H/sdByqIZxuXhoFgox01/G2k+XFNGQ8Uh9OtppR/FKa6Tq7MBfzL0hgqMocVaduJHROKg3O9nqb
NwhJw7saGVq6C2/jMYsb+UO4kaThP8wC55HTqgiJxDcWNdjyh1XpeUfkgjkc5DRWN9w7k6tzkbXr
+YD4MsP8Q7cvMUSngtfNDjSLHv2EIB+R3LahjjuyeYUUS0UG+3F3jHhM80TTQ9z6ar/jZbEMQP3w
VfEfFLgbQc/cmPVKoF318Y4Zbt9wNAvt1psj1fWbW4H41+5eIRqUP97AY32kRRcmGgB9BgJi7a5m
PP5nap5/9LzdldLKtXPwHm2/nyvMpSEKp1hNgpeovfVC/IuGPN+i88j71pUbaMY3stvOzi1NRckB
LeWqaBdUb9ZE+PyhvzKDbKWIioiLdfNE/V63jBtxg+FU5o2sTWahOt9Gxsj1+aUWnXbcI+LFrStU
0GzEwN0BdrNaR36l6zYLZYBaYS0IPl34rx/bNDFVNMgF6O6QmG/svLM6S1XNWtDSmMXXRjTkzQ3X
CwcxuAl1tYGdPrRpNJMR+QJz8YXgAqZ6nADMOzQN7ZM9bmyJpU7tzdrns5jktuqtcis0AXQd8QfA
afEdgclS4gioqhYn1Ax5lkZR/T1s3pQkRvFeQ7813I0yizFPMMDKTCM5C0F/KrXsmO1vgI8PBG0I
5BeCOBuxAGfnsNXne8VY0qt8KQvYtWOArIaFc/WDhnoh40cVgBEFDp53sFtq/z1r6rBKxzRR0VTV
QOQnVLW8JsLEIX80T4jVZIEZtJoEm74/ntJao7rB1LrVkpk1/tVermEE4rmPEzQcGY5+bSANXuuC
Su+9q6pbGi9uEFu8Vrgd8Rj+rXEW4P5HaDhrMDRLv/ntab5nnHannHpLZMRLRJo5tUPHww/FkkF6
fia2pn9owq8vvq85ryEffze7r5r3NEq+KJo6D0OxJdnXMlAiYTDOgR8Qk9OARUFSBnVsJ/ySGFfH
v1+sd7QylD39+q6ehu8QeBudwzfIdAX0CbYTbNKFzrmTVclDSs7TviuiVaO2atvDIraW+voVqJbr
nAix8Fnd/ouEKGW7snG/0qkZ3Ih0EaSOSpt3oyZbi5QFcyLmPfkdQsKmM3fPBz+7X91mZKuqEIeP
1NajaWiDiEBMSJoGz7uDnwB2TKQdfMlUNo6CmGeAJc8iDJpX0DVV60oJaCFXcXp4sF5LYFV08VA6
25/6Bk1j2flI2UciWLlljimc3Yc9ZyuoZLa37cGBg58HOfMgqfwvCVIQEHVUkzRyoWRFwvNLbC8T
FfWVwF6FOlfJTmobXx+NgU7hu3PDLESapUS0lLouVQ8jAS5+Ryhn0G0Y97YK7wHmPSn6c7HlITVW
8P/KKqU/vbKcWPwfO+mV7ZovcXfMj+c6GELW3XluVbSZVbXzHWmXbzO3CkckxfZJoBfURlJDMK2+
6KNCoOdmnCYHX1TnniU57dqhAs+PoFCyHvBEU6qwcNJFWHKNVwVhMJOaJBqLS4wNwd6v6xHhOxr4
EdkGDlbwDOLXhE+P5JyVuGyCXRRx0AFXILDEDLwX1+4xUvP08VzZ3POwTSIDWKp4KAOIjgXPmwjl
Ho1rEz4XeBKD8UlAar8fWSCaebWKxESoanszkdRgefexLofu3n45rgYZnnbJ7G1WgmBMZGdBW8b/
LGPvDAX9YcvtrtAFJbNdoZXn/GG0g5y5L/nyRJu3VH8buQQIBtYgmVcQ6z6WGVQX2DIlG7hGkqrL
CwWVmj8F+KEmOsH+WsJxlGmi7/IFenfM0qda5w/jXJtcxUFsGIPdwrc6L91+VMbV1dr/9hxe3+gY
eV4sDxY+XCjL0uNBokwEu9p0QMXJnoYrLZFva/blGaHfgcvW7+UErLYHR04SVprZjcwwCnRk6fI9
Cr/xi6jeJlyPi8YuvP9432PE6xForKu/uEwj95l0O/eIfwxHNRQI4EvLUSfn+BBBu5MLn7BMH4xz
XVJQLGNKPGmOObtGSP4SmC+hT9nA5Tv2MmYxwCEwrI2Z7zPNBw+qkH8zxI887N14foeLHQ5cly7j
mR1P4B09zishHyd2N6LMuTeyVFuNMcls39E9RTyL2Strf4preKU6bKqQiR3bOzU9jYUS/Ca3L3JY
9HT86QKurNRD1ZVIWiWZSE3CqsXK8BipO11qlHRxL0faq1N/D6BBoyUVDEMGAbtyyIGYo6pkqhkD
34HC7UqiB+aG41ObN17huIujhUK4rddhRmZXtFhCFMoIKGUkwO1Ka7yJ5cWzo4upkVaurGS4IJPd
2+LNaOzWJNPXIDOj01XaOxsy6ipxwmBdGzFbInSMb6VkFRqfIeEmqcgOHSEQCYEos2SxpIU0ieR6
7z1SRpMizgoJBf4B/ZYaCeoTkqvn93wQqu/qbJmVgoEVfCMKNu/zf6yWBiZOpIseszaup7QJb9ed
53FE4mpx1g39W481fr1640y5u8qrhHgDSO15rYjfRhRm0FyQ5m6mkA3Tkd5yK4O07BM/XFaPkvoU
LAbnsEu3LxA0Vl8Y0JKFI3nyy/IjewpVDJMBWXxVRuvib+j5+3GhpTsJJ+TCEY2Vgl/YH6uv/sIY
DXbQyK5VYwJ+IY/kCCIR5hQkn16FRqEZ3rLXGhbq8a622AstKWVXms7g2z/VmYQI+GSa0LusoScJ
9mw2V6L/o40Qgep9sr/hyBR+NiUYg7WWLMFYqFYNc+cbyvrfki/S+oJvk+aHyByE5xx7crlAMb7z
v2uuyRCPOznLAXQ2UNHLP8TVyg/WWuId2J0Duq6a/SyJrFrWxpdbGFTWtWXfG+lgeK+q19sG48ty
2T1Tbj3Wwb2bua1FDBmlJphCA+WHcviKVOE0HAK4lZu3Xr1bNATllt8KYkFqWl30WiHKNgZttl8B
HoXF6+7PwABX67oDi0aBglrUMKcqBxfJ2BvaFvOH2nW2tg890uVRUiU8uwYFhr6v3XA5j3PnoIPW
NY5GfF5WsMkjtSTSDXMo0kKrSGvOBX+G4wyExjh6HNtUUHxOFSIM4BCWAqkRToVXhHPeQGdufJMo
4ubglY8p4zw7AMyN0B9W3SwZp6/q4g2+Hda6ZALd6+uxXoSAoy6rnRaOz8XEDnznHlkfLGeQW4tX
XkleFU5LCYDGDm67kJmNp71++DZc6CeA0oHevIzvcGQz8gKJe/65zkuDC/KAVgViSfTeZekMRAxt
irgeWPd/NQgyFVNBMJ5zS+bw8ONmzg9hWriX9IKXRQJDefaTMeFNZwEqyC3k67VVBMcMNIgR+PgK
UvyCwOLAhJPesjsRozjMOjxoa5NYqE2lVRRGXnK5yjrC90Wb2nJSZ9Uqxn36jcHSzqRcoe1wcA/Y
iH2BDDEmWoi2SBeMOtJwC0cxByYgcpH34DIQ8SFuZIfxKplRj/gV239WJlBw67vABeSbD0RgyAOF
gchMc3Tp+S/D/hmEGLZmP5wmFycNaanQZA1Q5mUehVKc8949Ko3cOgQsEzJSvAJA9lcHZOkjkXw+
CniNCeSyN03ub9YNqVyBL96E6zqEhEwF9jNBfutY9dIBwCFnMV+w7vro9G8Alxq6/gH3ahQvHWXj
kWoShLCRuEGk/vkfvrISYe0cVl5SsodWVCUAqO1mj00rilz6gz9SoWyUesqgnC2BuvFfXipB/K2Z
qL5LyjHYKKfa8CKiEP1WetpF9Mczayh7h2TRDVvAkt0Ryl9mOjUy6sAjPyjrZD6WCtvQfk9sjlFm
1ZDqDFpDp0eHoWHIlor0DplrucZ3OQ5ZHKwBg6j93mbxgzXUiHFwleuySd4YwDayiwVR/O9Hp+Q+
mSbIsW+USn+UP5hbpsa2pVA9cdOnG7bJHXHWeDeTUSBubMjAmf6P1omvNnV0ADghg1QZJpDqz2h7
LNiVywygBARogvQPQ5RQZk+BkjEPbWNQDZeVmUa4KTJABN8J+admjly5wpteTQ1Bdj0XVpM+NoQw
U9yiDDXTjmiv262oSYTiR0Qtj+6nrXvaKXiFXvsLnRnbs01tjoZtf9A6uySnnoUq+i/jhL/i44L9
szZeXkrZ6Lt6PiQQbZcXbfzUgaZpmJ+JzwZ8KqNl1N0v5IsaUtfotNl/7kspm3OWTzwT6YMreUfM
xVYUKWOKvby+Q7vnAwXGaWtvLwwoKdeImekcMaqUJSMnMb8T2WFgBhLMzjg5QixTW7UdpLODGNfD
eqJkFmfwFHlYJdp6NmSBRBRaDldjyU8a3efdT1H+PAQEbEuZQ8DzkL2X14p9vI4gt84XdCRLaRlk
eYqrikubXRc6qeP+bIYyO8lgkiFSAcQNm5BgeTG3ggiDz7O9RNCijNxxFBCPifkxq9Tw6xgwV8lF
ioaaVt83OIUG1tqCbSrFQ4nZ1hhZSj1+hvK2YXy7Fz5F1V0K2elU8K/oJpd+hpicB/JYQCmEFN1s
uKEe6pTqFbZPi2ZNA4ZN3BSGy3IFrfbukF04GGR+IMdVr929+BIdJhJC3AlyPWz3AZguMLKsk+sq
VCuS7sYzuHy0+M+si3ii16pL8RGANMviXK7RMw0kKeDgAp21art3bw1Q6zcx2Qtq8GFGvK2xt1cG
+sBYiR5EM+KCqk2isvoX2FNGIOP0dCShe9gCNnfwkHQyvMg+KRYl643wNLRU7aYTXBWoMG5es0QP
Eu67Bgdih0lyY6cngqiHx7IR2j0i11TfyUbzPozvfu2B6ZB4Ku0UV/JSQL3OVuMfv9CuGsGvwUCH
lE2dHP7GFp8xvpgJDDuVh7GwMNq+VUXXQSjizZJ/iF13bF7Ge1CH9bjmYhYkgYXH4/ASfMIG/LnZ
Cmptj3H4eHHsqGv31lp5U9CovkFYvnIB3yUbm9SlmkbKwgs7cSfSWQvyQXznOJF03df3QQdiMW7i
wQUfwlFdMa5b36lYTQob42pT8YZm4I1/sfjLeLOlUp/dJyMPKf8132yQ9pgEFcEWKHRa4UfRVaoS
VGi4zJDZR8y2stz3u/Woc3GFDZ3Fcxf7nF1/N5wyt3kVT1+Mzcbr8k69L31Bdv1fNgXncl2NNoBq
YMoLw8VFSxtO82gtn/nyGBTClybZctOqrUJpxJlxz92BL7CWw8KKGnWtjhJScW0t1vncCv8Y6CT0
DQ1F6dBsOJG4E0hh43A5HZD8DtVCqvUEeTRuYEDJOrZgk/qxoWAnMYZu6ykuXQVp4Ti0vsd6nTIz
BpvUmGpeIGXht+L0wg+mnght/Z8yDGxVichEoV31PQEd6J1Fg6rMC7wY2Pq8QsxH/RfCte2AGuzo
C4d/49qugDZQnHTRm0kvsgxe99SpZ7lB52gnEWpMHBVEwn/CwhyHi8JfRT9/3NGM95uZrekw6JWl
Qki0sao6w5h1EbVWkOoJIWeg8QL6b7qB34w6V+mbAQXbKQney8GZfAq/hBoeKwI0z1atiPPMBLnm
TkEwpvNIwxba1G1x0wDx4n9W58jEprkMb7UNqedDW1U62BIjknXAq5aKcyKM5hYJUrOIGJoYbOdB
2hF501e+vrzzkLU15uLj/5Q7mquHrjIyTnz5zT6ZjBsntOUdy4dT3770raJBn3XRfOgnC90XNcNY
6prN9qheKg2D8AEkUNLSHl7/brAAi0VKsNcYZ6bvl1AiXJkdGyAKBn8byyiyckD9w/x17RkX0hcC
spSUcTfd0k/Wlgu6NXLgldXH77X//zgZbWqWj47sgEnEC7oGcFnGyCiiezC74NJTMCDL6Oc4FqI9
04oNr00rygcir8Ej02MANUezN/+XocCU28t8k+AVJupdmQrt93HqOi3yKqIbwGcbvchEE6aKQqKx
bCSTEQPr6Kyr64rNhbCcGbMXdCbDewjuGJjaD8lMIFAEk68j8jOocpkpwatrg98HbNwGWXG9D4U+
QxEcjM40pHXdE2jMBI7n7l1wgRnNIXFE/HNTlR+W8c/B2b9Wzusl8TKe6AHmCHOg89wInHv6Fwnv
bbwjLYzpOVmhj+yQi8bmk2n6bdWSuwg43zuF2FZs8F2q68chqU4J9LAarM2rT+3VoC4Sw+vEaRwN
k7BCAZJVqtcunn7k8BtZh3F4NpBssnO9twP94e+wRugI9lfaU5Q5PMTyELhQYhRG9iA7oWJtsxx2
PwbCFBDnJtUaEq8iZ9kbuRqiSimnaxjaCaDlmVaQPhGqs6qEBEfy/yltyJfYzfshKM1YsuHGqcBk
+iI7Vf5zvyOYrDVFlgKL4zLdcKBf2NrB7I21029RD0JTeppH2cLvWtc60LLNDqoWqlCB2aM/RRw8
0adZGmLLa19yBNux/bd1dx+5xcYuozcFQAR0YPSDeCAuDCQCLu7TTwppU2NyO2XEgEv2lK3E+tK7
J0QW2M8eFQ8VLb/OUa/4JqCPyDGRKD7jWBjkJRuYzbOv1PkOpcloaaMWS4Cd4z1lVj+BWa7dKGAX
0YtukMUtCyMz+Iif3ta9U3gv1WswfE+nY8yYZqJRNC3WX7aKyiC1+sYp9XGA1l9As3YeVicLzZgg
hnJR67JdeySi8TXva4g/hvUJ3Ct7cfGU8CT3kW1nMj1YvxwVZfVUU8QSV2xtGO655KkQPNSDMoIc
uNNeXlCsiO2xlJgUQvCdj11kbZrqpKPPY0ZrtiP6duiyz10G/oHvq26FN63E7TmK+VBL76SNmwuD
nztnLgFtDb4/oAzGtCNAxaWaFtqHB4g6lxLHPJWbOuUU+8onekjEsm5/+1uity4OcSyksjUSnAML
ZO3LQhoEWToo+bxor7VszfwJO42lXuttEHH/+jlDBjnchY1mdwNe3Sb9/m/IgtGyCjP2BvBNTAU9
HP8xRSELmI0fystMfKxppvhByEpBtcVG17xX1GMSF9muFYHfZlJr7GxFwW5+KM3+pkAtte56Q2DB
RIYROupLAr9ft/TR84vKUFg541oqK0UzKf+4DVf1cCpFuKUssgcsL+ISVBX9vvdnjV8tpkF8g/AJ
RbxxPqkAM4EkAOmCyoxv86cYYMIyoaIB3k9BwuldKksRgUitu0v+8ST29sxSap/fnMqZ6X73A85H
XW2/Mbly0YqxbTB261jVjisvR7qxqa2dF6p2iqxhLfcG0f+O7PeEUiNZCobU7DqZi/XUX9Ws7FZJ
VWvlLap49f/LFSrevbrZyKtWvVHtw3V7FiKdRRtgfEPqpN0PCv1rnSL03j2lUuhcQ+mYuZaJDE8U
+6T6rASCxug6Oyinu7AxHOfm+uxMiK3Uzpt+QSM+4hdRI1/FT/Uo/Iu5e/AG839h73g3p6+vRPZ8
ht40o23qHZKlEySf8JcF4n00bsJqtCPefHKY1tGxVHfgPyhFrV8InX55+7HOzzr+AMMHkRguMj4i
8QDDYF0hisPoWjmNXrV6t3NeZR4XFHZqj+jG2qH4O7dGlvs3KgeLOou+ZE27FVuge3hj07owdRIp
HkiexcQ6SEo4jxRO/w8mUXIpRb2zXNj9JnMbFIlmybxmZg34rdcD86VkC8MHdTAikE+uD6XtJ2uv
KJf+paQWtMIA0alhpIYMipu04IccuZXwL4BRK1HkR/S5Njsa77W1qMGe0XzCZekfCT76bpHhaf4e
BrJNgV7PSMpveb/zRghQKbK/gWaNzwv88Q5yM8VcWRX/Xj/tIabVliMypIFiicEGelJ2R3yonOeH
rNe6aIlKrS/1LSochuPzXy5PROb2AyeLoWNMGgOgGHp1oDhul1pZ5EXWlcO3Gi40DFsgG7BaEvfM
CD1oxeuhDKTeTlVn/6/cPtZ/V8CVCk8rEox5x4haePNj7vPAI1H6jhCRksrcKoSqTeuVLwzJxvZL
GpWvnl0FWRX3icjdlX6dPYwg8nefS2+y+68RZMgMgUckGoBGkA11CAGAg8TPMYvq2lOLMkxvXOyy
boXinLJ9IzQRSsejEEtSgrBK6QNFwmM/zUJObnmycZuSsYLIvQp6db5FBS3fzUP3hMwT3d2Pr2u8
6P8uKrxd8pTNfslWm/BGKhGGH7CkuP4zf7x1yqhlaito/RG9fz9e78C+yKkV+UnsoijBw0H35Rca
KEebSdMAZ3Rf/+0KzpemAlZkvmorSaqJFkKtGcHMzFF+v9H2XOMknGO4Gf58LrLQ7Vqh2aitwFH5
RFtXMf7EihBHBFHfy1RdbJ5E9duv/bF5GAvTd2Ag8rYsabnFECqEQttbUnA0u9CMo7pNwSviJh3k
DKt9vlhHL3SNuq3ZtWuRhAhHhEjkd6OnLfoU8S84FaLNIACL97xaGSSoqpeHRNIj2lJNDNhgbm/a
OTflp9ntbyYrczMyYrsPUqGonNBy7z2Furz8s0/WLXtP/hFxmx7Pd9Jet5s6MDJfoGbpu9OGIX1V
60KslGgV/jTMtzyAWowFvDSgCu+YOA5dnCbAS0LVSbjtU0IKcibZfyM+ip7pHBMOYSp97D45n4yQ
n4p3WHHi1+C/Cga4qNtCvcBr+F4hDS/X/mqqQGl8siD3dF29N7F+9shwKp3vJ7aEo9WmWKfOanLb
KRwiMSLTexZBpNBS+pT7Rsz1r2FO+rvxrXuGFoJ8qHWEeZ9slJ/7KuAB5mrILksjHHAopLgAYXvR
lWWaqEZTpHkLsIj8lWIRHEL3H8CKgu+aQH2o5Ohx9SWL95eLiTC2Se33jMIr6r83YLhZDFkJLccm
zGqmGx6XE6CydUqdt5YT2Zf1i3pTfqOZtWAJXMYJxF33aViKdyXuMKtoH1TBTJTaILXVTai0fXW5
j/9TJDhdAYgwqbqg5i7/ccmdKkwnr4pdOwUuug/9XYv0fKedGm11iPJIXP77t0KEiBe8iarvS2s7
jUOoe/9j2+LlKC55iMg8Z+EFZwjpJhD0W2Zwr+tBmuWEmcT8hN87VwB/XKgWZZJgKu79qh3Ra82r
pn1ULBJCypG+duoyzIXcfoDfMGfJ9YXQaW+wTwHoMP10XSRxCnvPayjwgNDhS3S3uv5WGa4Y1Axc
CfL+YfYC9Dx7fL8KgpG5JotJ5QWd5b03C/FMkevG58HxbABrPiv+qsdxoxhgqu1sL1EF434eBWxD
EEseWQM2ZSSvjzalA9Q/luMuZ3m2Vd4PmIfeZ1EAmLjTDm+VdWcKlUcn0A35jpq2Q1KkIrrWrM14
ez175VT5kJOqjUsiPQaEDkTbeu0bx+XamZJB/OJIOTXcOJPNtooozIKZz+crjNoI5/Wjab5k+yOl
UxsyQtB3/qDhDfi9SfXFtVq8lLCxC4P0WwmpNhfXUUWUhFBYX0cK6LbFOV4yMVB/c9SWy3yP/gng
8SiN7jZuQQ9BMXlgU2fKC6pCPkyTRZW7FTMio7g1IywqfO0MnzZ/CsDzshvk4T33Yu0qWhrwUC7z
xRox+WQj+5ZAlf7xv+oUse3IdFXtl+f0i6yTPwNCfJAqnmpgrA+MJrMn+8zGCKqYIqtIuWluPTjg
J4NZZlfUn0RU9rccY/Md4/s4bi76lqLJ14gdKIyX2OJkeobzKkPclg2yBV0M0e3lG520QTNHcxak
rxnpV+HdF2A4OaJL2TDkZoXARBrM6y/8+d+5+apBGT5BiQDvQiAoSJ9cUQUMR7hOYvwA0R55zoZj
o7YkZxlZAbytmLOpNoNPnPt3wDd/MRHFs6HJ1fgDgoCYWbsYVWkb7QhEubpgxQxWNN2JSRgB5R0y
kT88kFaBb2Xcvd9LmyWujaqer97TOx4sd9dHO2f3+QMGX0FRPS8sCtcwNNLIUpKFC+eof7W583mA
o1NHbq/IJgj1hMDg8loQoYjCiJijx1t/reUJjSiZiVw39EX7O3DxGVwGzFgWKgz4TBV0PUfSoYiA
pdjwv2WT3RzFnqh72gQssg0KGTBfk0/x2GMc7G+ZgAhxvvfz3eNGllB6XEXSMHRvF4vRqef1Y0VT
2BiiiMEaUU0MCeDq5M+saZ/58ElU99waAK3oq2RZF/hivv+ghld1Y5tT7knm4xaWZoJbcEkyKX1w
KtZ2qYCXxSyrljRbawxcdXhfECXTzdCu32sCa3clLwvwgGZfEx4AAT8MGBwXO7JNrxQP0Qkyx85p
vETo1YCZ5kR4ggnqbF7lZdqf0MYjaC9m+9fMdTHHr1EkHKzQZXSN0nd0swodL602OBeTwP1a9lrd
QyysrpB/ubLTzk4+9olHvyEotxKKMhhP11MoJD6EzyvQMWJaSs1ae9XPGTGeWzjIAJnPCoBYWpjx
xxv8bc5ORwMLHJPr3jCzWiANXAEvbegRyuY9sIUfhOR534ypFaL2w1mEHLCTDRCS7qagc2C1ryy1
07S+0+IiBZg86mwqxGdngZ2rGCxrdJzKrw8CBl5PY7ayZwpLxb50EHoTawvMDxy0AuXEfSK4vvy/
N6PP6r88VV1C4Ro2dYgYBzPqT7MBB4yXNa9XebQmRzqRjRdz1fHjVY0p9IjeecCb0OwqOZMu6t9V
wIIwZUbKJR3BaDyFAHKK/kIXX9o5en5vK2z/XhuHH2Kww0ra02c4SGLh099BZaK3B8O582YAmPqC
mJrtB+RCjjtOel2/3vZT90YBN4EaTk7wQdtAHIVH1URjmBvQSZzIeHik8LA4F0TyBZOMgbXWQJ/Y
tE2edw5v72HZ2XFJSg9ZQz08sPG9vBcVgNiL9F3RYV9lGXWIPto7/wa0Ln9feqpYum2HvhAicu2P
5V2VuJr97mdNof85Q/9F5E6h/8P5zhOyNUcxPn3Otja+B9SWvvUdqBhO6P1yIVldmMkz6oMReRAN
jp+8s0L9PdJMiMbsorHTC1OwzFhUyFCwBfp0HD9Ji9FHkQSQZFl5frOGk/xkGFV3vbC9kyXheBi5
CFRwS7DsBsQCPT3qmrN8Olr8DvEacqf6oNxhk6Ne8xJURlH9k+2oqXv5UU3TN8mxI7IhHxXWMBUY
fvRBP5lWvyLILjfABz0BM750cpukPj3CoN1tQvxVxl7moOqSkPKI7BocGIqiENPoROs9VPQuZhYt
gHo1/V7mEw5fErAbKxi4t43vhCaO6tudC5FKpMAyI3o6mVwJHWcr3xMiBQHuqiJbXEfNEhWFFIBc
2m710vvb89HFilxpqlYTCnnx0maXoMyPubI2MU+SdAjB9Q0mQ9yMJpxCPUx1UYRAuoCO+ORUs3LF
5/KzmE+OAoEav4e/vb1E932YUXrYkLnfdrUuyksrhUs/5njWl16oHg3M4VdMKdsAM2n+Ws2K+r/1
RHNX7LazI6yvIEPioDgC2Yvu721R+SwKHkRZ4NzYH+6DHUtrfKLypH1SykrEp5v4PnrMPShyPJbR
o1QgN8ghArDGpPTsRQapkIntmc9UNdRGQCw1EF8lnFjTagq8AlSVi+nD470nnXQRBsTBU6SQEkZq
Jp4LH+/4ZMfNC/7iBWiZn2dC9965EPyKGQuDy4JTokaUwaJWN3OchR3Vs6nlWPpnmBD2Tz4+ybqe
vJhZdhm2omEXEspRV8qjljuOt083+Y7JYjBRlKK8tcP2Gd0tpmecXqyZtXMIwXAwYBYqTSWjC7XC
JkfsyOvPKPnI74V9QXYNZLoDOofVidkKeKzdsr4Y2bZUFsJk5XwFNZfz2I12TxSGBs1TgvIZ3dzt
cQPBoU1FWJ1EKYpMFpIt7uNp9EGcdS9q4fGI7oXVFdw0hsg5BON9titdpXdXX9XxwhlqSCNP9jd2
FPyLBvNmz2YFsSS2y+QdSuxSDGDUMmO10+G7BE+MXchNfAXiwbY07bevfw6tb2OUnvS99ODJOfCV
QWf2k7Ws4BwRnIsGZph0t8PqsglxgpdcqJlgc4mV+iVHq/pFENx+T+HKjVGn/1Kyqc0MxSP8dYUD
8YK1yOo8PQhb77YtWMtWH9aF9eWG89pdiDPAl//33AMxiuhaBPkIPhBmMy/mXAU8g9n062UdqKLf
LmHg7xsLo/CoJHhsquTwmAYMiBLbVIBx5raV9Wcg1wUAB1Fhv8svlPWeahmlinfJGojPoU8QNFCi
FeNIoPs+GR0yenS0rwO+HQJlU7GD1JWOggOLhUKPFi5qu2sslD+Tm1Sn1+ZQmqPq9HoDbrEyZjc0
PuRH9Pz8035j+s+wsP+gcuH3GBsAdmJYuNYYQkTwM5GjiKwD3nk7/bO2mwLL+ZepMnJ5xz6d5R7w
Dp+6BXtIIpnJDbgo/CqxPU5yZ/iwSFK0bWn2oS12o3dfkVyJnK1/OjPm0iSkjYdVUyhUtR7DNdC8
0NM5kWiiJkL7QPJJfvU9HJ6PdrbY8uYf44bmH4u7ABGSkRSr08WYDkpMOioR3VkzJg0TsjRk0NoM
Ew4BYgd74VzjG1pNgZx0K09i1Plmb6uH2rx/oMpZV/jEtt/wAImaRyMo8+SFI/KDrejEQmOS54OH
XGM6D1fyT/szV0JhtrbHhgo9QP0S9+PyShiMj0dKiJ5lWAlmbS4D/IGovLY2SGFraXCct0rAakPg
UoymwJgz4JYg9XnoAvqMoxtSf1/mCvlIje7OlvbxdHhnGW3z8VPLVM4ek8wWf7lMYZ3Z07W9Wa25
oUNduwQ3U0fjdEOvTCZJZuhNExhA5XyzA/vhwlYX+zMgj7oz8yCWPfcZqGglMwsaBXodePv02s57
wvQ/sR2qx2jlNhLrY0v9lWCjGvPqfQ6gBvAdkaY4X/qnM3aFxtsehhIlMSQ1jGjrhKc3Mg==
`protect end_protected
