`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
Zhj0OOcUQnJqGkB1eu8d2neShXyqMogw3cpGmTTeD7KNiVtdL68j52OaWSSeeY6RDckJRHFqWTHw
uxS/pDs2G2nldVMgGZQz5KCvTKA6WCIUl0eY+hgPtxBmVrzrFpxoBLi1KrwdpKORbRm+6BTAPArM
ZFUl4Cf+yHVR6i/yWrUK4t9/yXr368K2h7D1zNACsVM579WuZzEG3jZ2YOIdgRnXqbtVy/S5BlR/
jfbhDdErzmHbUZQsoxD8hJij73p9zpIZeJ/0Eqpbexih/AlJpHIRmovFqI6XRq6NSIuuNx+sVHBZ
dExko1dGR7A35v4TAUQlrbCOarzyraO2cdhefA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="FkaMi5YZGgiOUk5FiX+Q/ngn9p+Y0A393rsZwCzdqWw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2448)
`protect data_block
o07ZePCNtab4AZWY/svQFNIoEP2CybfSveZaYLS7eew4lZWk2Y6NWhgacj8mtUTc+DaG0J/yh1kZ
isvGaw/WCL+pxVgi0IlCafjzvOvIrTo+CD33DLjjuxbdPR7g0DOHaepoyQuLf6GvCOhwDxgY48FO
B1gdtJD+YLuam5a68Lbqc3XZCXUxAHGvZ8Pb7FJQV01H8MV6i8PpbFOSayCJFTeelvfJj7ccXkat
4xu8u8T2xUbEpQ5jIVn/gghfPMnMabWiwUBBJE5w0anMCOjo8BSBI2zvAKuW5JNGCDt2uL8QZAlN
Epj/Xi7WGGipRd3OHxlHAB0OFFHFA/98yiwI+bqGBODmVfJX90N4F8/Bicec/1pKQ8Vwaew1G/Kr
M5PeJZKLNV6rLL3c2D/kQ92jZmw0qIxhKKtOnxNEGEN7Pzfgm254kyOsceIN5CQu4DUJzy0kxSYA
HPBaEhp9IBeJs7lhKyJ30B4uEAUsSbfUlkscOR0iGR27It0EeVPcw1pO+ZqrCoi+A2Rop5Z63WEK
FpM59/O9t00LUzbtQO/gAfEp+b9KT1MEN5quoPbvJkacWJfPEENa/K+Oo3G8lTPPDX05yOwQeFCH
2u6m4DCqHul+K2dUcKsXDqIY8uFwzuqHFD46DSzLPpVs7hVWJXETdXgap5igldERffT/tdQtl5Kf
QFjylLf24k8Eeil0FCfxIia7ddujHJxVq69V130HFiEppJ2DcoBBkdvtPmvZcml2u7vZRy3PmPzc
AYWZ16T6HOrX4RPoym3P5cT/bLNtQ5xkz7h9z4Oc5beuA2wMvAFCgI65H5BnrxbUrS5gHrrP1O/y
2k1H0B4uNVCSzq+cur+G/85qn2aldSEyKFnIJXeA0LqzcjjxR9zbSiD0XArU9/QBEHMgOyHXtZ5z
NT6+cvYA01ApsAUo/BfHsJqoWjTBpzkYLunMW2ZjU1ZAGFZtUkXzxQsRTjK9bGm7sSmxsubXLDT0
llnItQrQaf6uZC72oKUu/qFYtSoXTJF5KIdnfnyv3/Poi1w1Z12+kP2+f7eEjUMEgSpkSqCn+GMH
9ISEUoPf/JRXS2zt5DC2orQe3eSLv14jfV11HHqW1x8ENxZOyHPmSrRt48n8CrR5mn1l5gIXKMFc
aLKhD5izYO2gT+BKI14y4IUERmWOjZ/ygYp0pdni51BVaVfFBe0dYenHkW25VeIG+GKW5qR15DEk
Q939gjawiCyfM9tdpeI0aIGTJDybTnxNVk8Ayp+jxWG4uNgVYKP6WHPsmayhCXngBUyUa9G3BUOI
qOT1TyvG1NNGedQ5MzRK1TiV/jmylL0YOQzf3LrBBEauCGoz5Pc2UJ9s/Y4j4DQ24fVeDLzlOlpc
Hg38JAKoVdOD21ee+myHP4q7EYV8RxpEsJHPVR1cf1cqy8BUBSNfBnL6QRMHIsae8ImQ+JdEAJCW
3FiHCw5KhfRqkpTcZ+U+u8AAMAwpmNMa+JSOQRB8zOAUSP0a51Z3RVOSnQZ2bla2Ax1kvv4k1cmf
g3E8Lxy/wRM7yN1OEms5+7ftw2fzPZHb+nYonnbGSo5O6nXNEpj2oCEb0zXOdoYkSaXUA1tKkdUW
fCpRB1y2HlJ33vV4kM13wZW33xT4OJGWySNGgRGe55MOyQTgQsm0IqvbVTXVRi752/QfYuDxX9J9
PlZ3nMDR96Er+o6NKShncb1GED/m8OYnULq/p8lUK0WFq7mcWbwdnN+47Jv/c+t9I3sjXsMBqIcc
/Y55tB1HHR0/Lu9Xdq1EFr+Ehd4tKlwyeUKl2+hrnxILZa6NAji+DrrP+V1mxw6m7ahVthdSi/pp
BrZt51ZXlYFuYqFEGLNZAdHnEZUuAP5PjzPolCTtc8RfTw4Bx/RxwkOVY2w4BjEOxlwT41xTGU+3
7jQQUffn3vne2KU6Ys6tWGjIWaM4gUd8/TQMjW1G/TnOqPgyAJ0H5l8yTROLL7yrAB0thYwLBK5Y
nb0+bLTed4QLvKZPQPo0Hg36c1CTqX5Q4eRjgC38H0OeQB/xRpwdHRFWpZDoH6K4KvA/I2EBH9ae
dKI90Ztw24e49wui/2aIJD1WmzKzocyyeGioIj/ALz3vCtd83sHxFHw3iCdSLmnXMmoU2JVL8RR5
0McaCY+ia36WN7xwaykvssKoTC2OaOFaqrtTzAO1vGAzUXBFzWPUuRQtZtAmyH0dbLpta0GjzlRD
dReWvYWBO2BhLp7f7/YxNIRkPyBhgc+Wm7GkmuSqQMuyzTtGUOH2WUngHqWwBzRHS9cB81AXOdUG
KTY3iiDwNxVTxdsVB0kCBcn7xedzGbtBxr+uYZszCjJD1fDPj3YlAumv7AvPFCzYh8nLYc0t30zo
gvibKqtQbqb9V3dfTlqNpKb+NfotX1INDtC8RvJd2CWIJSaN3Y1wTaCeVAbhOcpXaivYArDoTAL3
q42nWpoO5WmV4XSZHu2qv2Vfp2zVep4BxnvZ4N6jqsBRScVdL3swzF2RhvutS1Yb4kJmk+ZhcX4x
Qaivn3b2EcJU1Ns2IgFMWjoOk5uFiCaMaV4gSHVOW77kdnY+v6Wc7xv5vmIBbDJ69zFeXbISfIkA
ubAdfHMrXBjW339fBaQdqbIOv/WQBxnDZnzKamT8n8Y9urw6wDchFPY3w/9I70O7+//6U9aLmuNM
ElHAXAkep5+krMhqj0aSPIBAWlvwcOMTfUEcqLC31wVvdCK6RAaSov7fA2DsbvPkVMLUAiJHH1rY
/zwDuqclp7/FfsF9Q1IcxQjnQ4cH8pUeis53kscUkNlCRFKEn2kNGPuOCvGIYM78gnNFwKZKZsO0
nZLodtTlE4bGMFXsLPVqTLrFo5ewm3JHk5zzRRar3mA7R+wAqZ/hDXPnkQGvFdAR/WGP5Jvbdo32
zb+8cIp4v2NVPwZyxkPdBVTYySSPGXjed1SrgKvdW5WE7lei8Ul+CPseKW80QshU7+afcItbnv8H
/PiRHmxXEcBNnbKg1Lg/vH5ZuuLWVjWLLB50sc4Z/McMV0afOGFY6OXUnhV2Jh/wxWq4gLr6+Xjl
9ofBQw46n/MvoOpb9vwRQuQqc2GhKhRWZ8ZtiPf46aa/pnNL8Sm0ZxiNVkkSpQa/S7IguR4NgB5+
z+GAPFUajATLM4KdRQPAFHLQYlDCeg/TOsvexJ3uq3jPODzkSyJHEBhZkP4H0dzm0CUJbbcONOc/
a2qyJ+VCIVP4PLDB7kHBWq4zUTfQvHEjFSAtLZnlSRl4IcBUbrnHiZmlTWsKC+1IIY7FdSaX
`protect end_protected
