��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���=�^���{3�%���\h�:�0x�஑�Z��:ԊZ[�J������a���!�v���0��Ȥ�O����h��B^�Zsχ�����֫d�odvw��%k��W{�{y���P�J�������ڋϼ7A��a#~*P�7���!�e��m�"�ɞ�4�d�U|�+\u�s]��},�F�M���i��P$�ˬ!�2Y��o;�\�������{%�_���u�j�~�sŰ�\�Tjl�[b�o���f D���G\5[������u�g�2u��.�h�G<�EÛ�����N3��>v�6�7�ޱ��g��f����­eb��؋�d�c���|SD����8@]�[�V�h�
����yL!5�NK"���|}v�߆/��i�br%u�1y�w����1��\@DY�X_J��-��S�?ݘ����-s���rZ�����U/j���4��W�_h�)k�,�9}��_���ؽx�n�G>����IG�q+��;7�̲�$�����bO<W�B��x7��� ��j��������3�]�flXW�VZ�w�Tn���I(�1�B�X�tb��-ri�l�نk¤�����������j W,E"�"��.e�o����3�ꈉ��`��~I�D�Ѥ���<R�K��F3Sj��<��ľ���ء[s��*�t��e&��N���i�^����e�4�j5��.B*t�Ku�c��"#'&�ӑ����W���2��d�띻B`��(�Ii�@��������w� �	��&��AR=�Bwq��/�Bgqf�6|ן�����װע؃D���碌
:��ghmײ+Ijr��U�5����&���P��T��,?���2�;2����Ŕѩ[e3]h��p��}�]��9͚*�?DiƲ����i�q4҉����W�d�K��}k��D����x�R�-�H�fh��5lH���w9Yj`Bj&S��1�ء:t-�ᖷ&�潗,��o���W���JR[�G�r��^�ӭZ)S��F����7�y���x�
�~59�Ԧ9�ɟ���]�L���M����S�{�e����7Tΐ�2����;7�C �n����Bb��vH<��V�(~�hU�F����7��ʊ��a`���b1%\��>V��p�vs��|�0��^	����pS��*�dP��t�����£W����9�PG�H�ג �$tc���=�kn	%u5 �3��Xs�a4���ߒ�1��G�!�p�w o?v�q���:��B�/I�vW�A��^j�qh��:��^x��Ҧ6<���`��J�!)$~�o���\F�C����0��7�#a�����_����3(�Z�f��^u4>!Y:e�O5�$К����HŔ�I�fbިE��#�V!�f��"�������f���&�}���ܱ#�?�z��T��,���C�!K��k���sy���"���_��|0��=0����+jj���q���X��Z�%|C��V���Sw���+�s	c�65�-�uu��t����K�C���I��jڎ�O������XM���t����>��Ok����\;ru�~&�4��|� ��Ǵ)�0ﺮ+���]v>[d�/^}���4���B��[�̟� �@F%Rd'i�[��6 H<Y���Gͣ��$%�X@I�3�g�A`7oA�e�5cY���nA��ѕ��%�Ot�'W[Q����r��V����ш��b��s' cZћܚ���us[�e:��.}�m�=�U�r��Sxv������K�
!�Q�Tн\]jg~���Ȧ�ɖ^� �:/3�=P�Dq8N������	]��?���%vz��Y��1�"�6��RI<>*��ǫ��]۵��[��HfϮx�H=���&��@��C=�"�U��r�|�,}�(�s��S�t�t�b�UK۞(qk	����?��O��;_8���Lɟ��U��2��MN���A]��O"p�{[��'"8���$��TtKSm�;�Ng�ݤ]p�q����D�V���Y������ޘy�c��5�S�SI�r�R4�tJ�߸�W�)�ZZQ��Ȁ������g�����<ȋ��g�'�s=���l��<���,�I��̫6s��d�{Yſ/.7��Yp�X�|�R���L���X{����I���u�8q~�Nt�`�b�	�	K�r��٨0QW���~G[�qqx c*�KuhL�8���-�F_�{�B7�l"����_}�} ����i����V��ksRk�Խ��BO�OB�^ڙ����6�M�������ڈ�I	�K/��l5�!�O�P�h��#���>�`.���AV�GL۹�\q|쑉l3��G<Blt<�\��>���MEP큹w/��+Oء�ڜ�����8ǔ}a��$�m�Q�}?�+��rL�ש��kY鉔�Em��7Q߇��Z�T������j:+1�<�MM����m�T�s{$���+�H�����ޘ���l	���N���K�S:9�Y�Q�Ȃ[8��������%��Ԙra��C���~�;,"|�4�b����+��~�H�n˘�F��6/G���Z��@�z����l�4�EGM���0�g>}��6kSʩ+���P����2�~>t����d5��r��?�{�>�T��G{R��Kg��(*�h$#D���E拜�E��i��dG�ѲZ�x�F�ξK9�(��'�����HZ�#���3oD��<Ys�����G�!�6��b6Qy�U���*��>��8�C�/��E�빅�Kwva�&����Uہ����hfG�
����-f���|}r���t�Wo�VqzWRD�8Z��y�>��]9��f�n�?w���~x�Hv��@��_*U�����[u�!�e�C��r�����g�^y��֯����g�;�!���]���	H3i���곊_�~"q���m�vT����fB���"9�/��s�f�c/�t;m+M/騤\�٨�rI_%Z).���8f�`�$<��R������zG�̟����3Y )�.��[�g7ɥ%��B~����~���Ƌ�AY_#�K�aj8>��,�d�A��$��D�RP���9�0)�����S*�BZ��&4��nfa���`�lƢ�0^7@]��&�mJ-�e�Gwm>�,�e��=6� ���JoJkc6����2E�c��5]��D�v_��0�yF�!�	l���a��^y� H��(�7@�!CX��6#���m	!�n�{�HD��a��Y�R+`r�e�����O�M�ѐ@�8���I��ȹ2er��vn�O;�@����zQ�%�'W�������<j��S����g�l\�EB��c��z�D@}�����>GA�6	�́�Z��
Q�@+�c̼M�H�<,MZ�+�S���W�ބ�� b>�3�9�1�:�������<��s�U�Y*��0� ������A�K���U�eku���p��أl@���Y�?�s�#o���,SVp����"��[��C#_;��&q����G�=�P ��i����/���vz��'��PRL���X1�O3�S4����~�1\�AX螄���Jȕ}_�\+u�G����A~:���A,�L�_�}�AI�0��Z��I��՝�R�Rj��݊�?�0��J��L1N&h1�ĵ�[���@9H�c��(f�Na�0іp�$G�V�g�ru��<�#���}J�5�:�T_�w��W�o֒�rw���#�'�����~ ˅�>g<���m�?b�ηϒ�g8D�t����%R"g����NYJ"r�s�kWE)Hظ����a�݁f�4J�v�[茿�z»FוЌ��mN��,A�\��I���Q3��o�����[Υ*y�T|�l'�c>��"��Ǥ�6�dz5����
/P��D�\��kH M�,P�ݸ��+I�����pz��,��H��2�[X�.Vs��e���%��+b �`�h{,��er��-,Ó��Y�n�nD|OA����/Y��5��.6�h��Ym~=u �Q�.�qV��_�3�e��~�?�pؑ2�b�O3�<�L�,��T���< JJbͷ�}ǰ�a9�o��%oP��$��3ؼ�Q������KZ�ٟh�y.<�zq��������׻1�U�����.[��˔�ߪ�{���R!;���c8�2Q����T\��;'گ�x�����+��И���>mI`qZ��mĳ���U�gB�|C����>!��k�$ר���z<	t��8�a��[��.�m�=�I��ڹ��]�n�	�]Ł'� ��Ǜ��V0��>O>u
<����d8i{���$�(�X�yO2�D�z�}��+2�|�/�*�/-XaVs�щ20�c��u�M�:�O"������N��S�X����f����`C�D�Z~ʜ��y '�]y���R��ʅ�I��r��D�@/��(I��<�c�`A$� ��g`�� :�bD���!oi� ���T�l��_�5�a�YR�w�7}�i�-���9����@-�t��H!�b�O��-�g��!RGX��{�6�gN��Bc�_��n�*Ag�k�>V�����>�w�ܩ�_����}Ra�l�"�Kf���t����O����lp�z#�L��-�D����vQ��?����Ęj��\��"PԪpT�މܡ&(D��E�K��]=�B���Ϫtnc:B����X講}3���@��L��]�)��?L�m�۴J�SJnN��$��h� x���L�7�I�^ѳ!7�:�F� i��=�<~zE[�]���Kϸ�g-�i ����³* �����Mc�_$2��6O;ɼo\��ɪ��<����(M�W*Tpd��Z$@ik�Hf$':p�cʘ;%S�k�p��H�����6�����95� V�P�19S2ۿ����wx��=,>m�<�'^y�ǧ*�(pH�qp��uI���A�.J����b�I;C~��eK[��t�X	�$[�Q��AsK��,�Hh-���,��t����ДP��M%a�?H��p}���� ��˂C�k+7x�*���!�2�-�fI��6��@ A�=�����*�4����k��k��h�iہ��XR��h���S�{���q�����ڒ"v�4P�{&ny�����!gA�����A�T��NN/�I�`�0�㑳)��' |3	�h"T�&�0Q[ɥ�ka���
6@�o#z�9�������GC}���#�<� ��\�ve��c���a����au��
!d���n�����Ѿ|ҽ�$�X�Pu�[�t=��<(+݇k��EX�B��QF۶#5�������'�2���h�*<�RWi؇_�fٸ��'XB]3�	�9� K�}�#�]�~�H~������tfmL,����y�r������T��=���+3Z�{��9���fڣ�%������KL�*!���jk�KTƋ3h�9��;R��u�|�7.�֏,v:˄��lPb���5�Y���]��ߛ�Dt&��*=~�L�i��N�_��3�OXi���0Q��+&{�b�:��hN�"^ӗC��، �'�{�#W���7T�V,eʣ��������P�"�,�ɼ�Q�.<"�[�ߛ�Q�-�v��Lk����?�2��Q#0m�M.ao��D1�9��K�)𐨥�k���D;��
a7#����cpuk+@�7�X��څ�_! a�k֦��6��N�/N3Ug}���l$�����q>�3�� �N�W����ϗ�gd�@�ã R硚,��Xl�N���M	;RZlF�{`Y����� U�mށ���n&�}�}{�.��C`�2u����ܯ2��僺��B#��P�!�%H'����	k������nx>��0S��/f��#����=�bL%@l����ER�k;��ުf�Z��-�n�}<9%|n\�sQ8G��&��^����?NA1�����:�fd��'�w��}7YR�ɢ�0?�!@]���R��w��̦�C5w	��p#�J�p�2{6_��hw�x�$��5�I�3�V'�B{�|<!��%.�q���毴S�dJvB;�n_�C-�_!98�sִ1�z��va�2W�b��؈HU��e���X�o��E*�������蚗��\�_���.������3S�Y�j�V&i�-�=�t���Cx�xDM�]I9�$�	�<���Z�q���G�f?*�o�C[��=c�ʌK;�n����lZ�a�R����d���n���x~�bkP����*o��+�}4���ٌw}�?
 ׸
�K<6�W�;n��L/03����P�=�V̞hՔdyH�@Qd'Ô;�qdlY��?�������^�H,�К���eN_�;p.�Y�9Y�z�F��P-�Ϟ-ɩ/�Ϸ?Li�ܬ$��Z�v��}M����8
i[T.��$^�5��:�[n0fR�˯C�1�0���r.Ç��4v�m�������5�9f1Ĝ���� $ں�I������_;D��+��/�e- ��[������tC��ٚ�� ��K��owk?��CU>ѵ<lw_"�Xk�1F��/l�t۹Wuꯣb�=K�?%˳Eѣ�8а ��-�e9%:v�n�����L8R!�hc�2���7�S�C�8A&�C9�V$�����l��
���B���Ѵ�e�l??�¦�G���
��_�r9;k���*�R�$_3fC�}��D����Hg������s��u(������C��s\����.H��q2 y��pu��_���Ԍ��s�[9E�]+��X�+� �ԇ��+�!��o� �P�9���aiw]G)2d�+�$i����p��>hS�AW?IwI��~����J����Jh9���F������_�¥��"��㸴��nuۀ6-[�mT����\@�]��:�Yf5'W�l��[6����m	R)�	��)ް.�����f~��8]x��9L��I�$Og�ȉK��4����u\6����4z�S(� �~��Ql�Ԅ9�����Ѝ�Rw<�ĥQ���$^�5֨~g��c91,�E�م>=N%�^8��t��f�m�A�;Sr�Tf�-ߜR0�	�U-1b⫈��,��sG	�S���h&�h㫷�r��4����Ԥ���6���n�����Ap��>4R8ai���h7����(�i?1#�X��'K}*:�`Rg�*�k�P\��<7������d_T�j�Q��H�O���H�ƫ$ڵ�M]�t7?��������enϝ�0O=�C����&|&�� �x�/<�1��y�F��;e�_�eȷJi���=e��d��䨂}4��q7M�u�#N�f�xY�y���!�C��4+��>��n|حx�� M9r)�wa�c8N����f���O�	O�M��>X�s��+;h<PO��wA4��t�m�t��q�ۢ���-����4m��:�����e�qJ�`����!�����_���k��N��E��tʝ�q7�fq�QŅ����@��I�B:���;ͺ���P�X��=!]כr�K��da�{�=�(��!�)�����@�WI~���:�!*�[F�Yv*���Y��j���.�&���fƠ�J�X�#R�"���z��]�dӧF�.o�X��;�LlZ����*-&h��E��,��9���e9ǠGDP�%K�C��5�ya���9=�zWCKp��=�7�ϱ�o�M9t{"�qX�Af�Ѩ����v%%W�eU�5�U�����o��
,�±8���7C/[��r!T��No"�Y�jD�*D�����?g�r��˺��N��}P	�Q��A�l�^�'��m�����7��z�u@�/������KB��@�,�"B觋��SqUj�BvSwH]�Q�}��p�i�.h)�=����k�d�� �p&�GB�洬V�������?�qXC��z2��s���В"$x8�x���N�x����К�T��3���HG�s�����w):��J��b�ȓl��b4h�{���m)-O�S�Em��U��F��&�$kNr��T����M�Jc � �H�3.Gi?ا��Z?C3fG�RY��\	� u9s�=�>���-�o{[�I�T+-��1�0JP`�t�.}{��vT�ޡ1{|Z=�R�[�����o��&��0~�oOǣ]ь���b�0O�fK$�O �(Y���q�JP���};w��c���B�J|����B�T�X��8��\��vU��«'T�VFA�=5?s��|Q�Û�wt �|w����\��8bV���G����9Mݾ�.�,��[7���ceSX:뭣X�wؿ��f/4�$/O��oqǗ��J=���!���I���}x����s�SpjI�Y'h�=�u��x�^Zu�|�T~�:\����T�8�>��7K݁ٽ�<�-�B1-$7A��9P9�P�$�n0g��2�:�|ʹ(6�A�[�W�<����<x�iSp�1ύ M���DL�4|�!��A��9�1oۇ��i�`s)B�����E���X��� �D��~����ƧK��V↔7$�V0̛�F��N{�Y&V���,K��$4dQ(����S*���B���hZ��֩��${���:�{��A)�n�I�)9�6�V������LFj�2�	R��evI���u��B `3#�����[�#.�Cb�G g:HqR�#�S� C3J=����2��#�肿�)��+{u�*�m'�٢o̔Dv�:�s�6)��2_�Y�������
��
1|g�>��M�k e�F�/=��x���|��!�ˆ/���ev���	�3�G�0��;�:�Ɖ���RZ�����5� ����c��v��e���7ō�g���jCw(p�;��_d�V����F-/HL:UK�4Ь���_�+{����Q!/r�c=�\&|
X�MR 0��y`�aS�$�L�n�"B���D!�em{Xg�E6�����%o��W�{�o�Y&�#����aC�׷#�e΄1���6C�6�ryޱ�٘�n�cG�c�o�5= �nԭ%ڒ�u�s� ,}^хF	����mJ	�VQ�5K��t����`d[-��\�'&��_A!ߔ�zm��Ym��+���l�{�%?T��לÓŴ����3���Q�#U&����U��/K�\�3����G.n����9��k�O$���:%�V�~$�ū��h*%�t��9�;S'���Ը�sǽo�A,���_
`���h��P�ǭ�*��2� �D}o�s	e�O���"z����y�Ɏy�����=5W�IF@��Y��b7��R�`�n���;qC�Ά���z9�YT��JDd��%S�K(��h�;�/]���Hf�0>�\�Gr�,��{as�p���¬���'Oa0O������r��?��3^Y��v���M����e�4��Z�YE7ɐ�Di[��6��r�NK؇=���'�� �	�3z���(&�j2�3߭�/Or�e��1I�`d#�ʌ6�HR����h{�,R��%�=v\�FT��ʐ!0�<}����ڡ%�+W}�^�W%�>GN.x(���%�����a�������w,5�?�W@'qT�;1���\����`�9Qh�E�x_X�m��	
�ŕ�Vm݆��㥙�_Wk�t������UZR7�x
���i�u]F�uBݯ�zm��r���C@l��Ј�"̧A�$���.���`K�-�0VT&?��x3 ��v<�L������%�.��r�!'"�$o�w�U��b<`�ytN�k98�=|�}vm�z� ��7��w��fy�]O�|�"D(�zG��LO*�	� 3����F�CiL9w��	�Ed�\�6D<��}b��T^S��?+6�1�݄z�X{GxM�)}���M/���[�uz����(/e��®�`���q���델��
��A�п< ��}��C�%[�.>���Ќf�`�K�c��rN;8����J$Dv��y��<5�2�ϲ�(y�x�D�G�M����[��gVzր�[,�Y�['��!�=�Hl�J�����h�cp�	�ӆv�i�\�0MS��~ ��0X#8�/\���97.�j�P���D�c�AzB}�/���|^/O4F��^��?���L_ J�����Kt'�a���n>��}v���2��#��l��&��S�`�Ә�mY�v	������1�V�Z
�T�&W�HX}
������D��wcn'X/�|7[�K:+��c����8n�_3�V��>=���cB��C�CD|[�5Ѹa[�s�1;�9�����1�p��:�g��bSTm��nS��2nꮱc�!�0�v�
��c	Fԃ�NҮ*��2���On�1Q�ġ��0�������F]�8yiF�=m��*<|n�F�Gu_��[C�v��h*�i����c�>�Չ�1J�抲�!m'��}"���b?<�0���i�҃!k���TS�8�����v�0}q�J�6��ߗ왵+��׍�����ð�ʏRP.���ed�c���g�3��8u,���tӲ�W��ƔY[���1=���1t�A��9��<
H����*1#�fIQ�@�i?�0�8���ș��ہݜ����M6v���C�k�`ĩ�����?�zJ*�~(r�������}7ST��� g�y�.)
����;���i�,F}���+3 ���b�d7"�WbO�c�������fqE@���ZĢ�~8  1���jV��G�1 p@|�M
��O�`Xb]]�Nx㓼hOAk��	�gn�w�������Q��Y���
�Oأ��bW��!s��Ň���_`^#�(̾��V�P�NJ����A�tyc�\ӄS˸����As"��i�TG��ge��lT�	��	���X^Z{,����v��Zk�J�����3DdO�`_�i��/E���v�G�dŖ=Q���t�k&ɿpețn�F����Kg�i�"�����t35/��QNgG�x��v����^�?��	�i�[F����Z���֤��J%���5}�N�QȆ\�2?Y	��Udn����-��U����ڻ �M�~��O);���GD>�6nJ�p���Fc,�:�2�#i�gh���zvǤy�
M���
}���K���@!;*��Zre��C�r�_w�������������4&-��ת�!k��ZE�Ks� `SV���
�V�5�����,+{j�W�a�Q�)q�cϫpW�}��˶��$ۇ& 3{��i��%���Pٽ<G�Z��qW]�����ZE �m�΢��A�LR�s���TҒ�O�����F��=_q�:��m�5@��y��+���j�o�3�m�7��{����K(�}:EFh�b9�W�(�ά�W��q	�t�����$��?�m�0��8r6��Z��U�qM2B5�U�ZG��a{83� �d��(����<2�X�q�H�+�5�o���qD^�=��c!AA"��Cj�4G�����Q���Pf4߃
Wgy �<�+Y���d�f��c�F89I� }�㦢�[�kP1��$Tx �z`��:�+,�|>o��x0��ˀt�Dc �N�y�5:�;�-~㕳�QI-F�
��83����H���+-d�P/�R$t��2[�����iŮ?	8n�.3��3	��Bjx�}��æ�u�o~h\[	�y�A(ϳ���w�^V��
�h�Ƥi�!�i�{�!����8&S���J+g�u�DC��E�eK��C}!����6�:�WB���*f�2���й��d�a��&���<B� ȦЖ惛g�]:6�'�9@N�vY�+m�v��O߾��O|��_k��Ru����vIE(�1�߿?��z$Z�PV���,��jr�r��UʿO\����l�8\��D�$��d��S�.�q���Ƈ�p 810$i�d�"�d
���}{��Z����ݎh/a��]���P��妇��@c��R��~�\��俹��!J�9��;�s�Q�����
�E�5����&�I���53{K�%��D�Gω��t��UZ�;���2��B`>�X� �I d�0]�6�$�ec\�>[�+8@����N��L\�馆�6�i�*�b�]T�9 �~�+�$yg�%�������X��i�1��;2�L=����y�S���6��]���L��╨�� � �G���1_���x�!���u��c��>UOg�'5��_�}n�0/�m��1��,録�̰�F�B:l]������"�3'����>p�ؕ��0y�^�Ձ�nx̶�OY^��N&m{��B�5�u^���3.+D"��	�[�Ca}����]$�%
Ԁ�:�K�Z5��߭w��C� .�����~��dI],"%����x�y��Do��h�!�ò�5�H~���92pv���0���0�Ûf;;$ܕ��e%���0j�.G%ȃ��]�0��]Aj��p?+ۈ������Лf!�n^@�Q+�u[��13���D�|�4yw4U:�tGR3B�od������s(U
�V_��ɱ��}�PƯd�8k-� f~HȪ�H��*� C�<�D�>yV�L��0��hS�"��cۉM�g�U_���f5�"�������@'![+�3���|hKk�&�Cˇ�O߆qx�UT|.�6�$4�	���X�',���;"F���}��E+��(@���N!b��FćZĨR1Q�v�0���,���1�"���x5��otkڲ��/��߮jط�7-�hM������#^���4��<jE�%�7I��'i�@Jmy�p�I"
h �r3�-G�.���>��O�Wx?Ӏ�M�*��g=y�o@�S+?jr���[��+����@V��º0�N��������E^m����D=3���ʟ�I����]�}�E{�l����������W��]�������|E�憴�����|4Q��,,�~Bqv�;*�9'�b���	I\����n�-~�D�>�t���/X�����xE�lyt���qF�k��ٌ6�9e^?1�}�Mj�
P�Ҡ*���`@:JP��Jӭ�lDu};����l���=�i����]8(�EC��z�	����O��9��%�>���nE��`��C��H�c�AN�f�ğ!8���M0(3�� �G�&��'B��"����c��H�g��n7������GZ�yƴ0a� Ә2g��V��X��QjV�N|2m����{�8y���9n�N�X�p��g���XӉQ
\�sW#ef���޻SX=1"`	�=.W6����s�D\1��g�s|��7[����@يT�7}�f������<Soke6��8��h%��{8 ,k*y��Po��#�s�'́�G�!�>�f��@
��&�R�F�/�?!��g�Re��
��P�0߈a��Q| 5�{���%�&���ʷ\m��.uc��%�Mu�]����̈�J�V#e����"FT���9����Lf��ax���t��~����D���0wI��Ո�Aֲ�%a�aG�cd��ӄ����f��W��=����>�Vkg�_o��y���k��);@m��{���T���Ӷ�b�# ���d�%&������+w"�94��t�Z���b���{�%������W�I����p�e	Ε��UB�g�e��J��U��.��6U��ھc�8Ǽ1R'�O��M�Dڵ���95o���sNQ��\|e���Cu��D �qyj#-v�&ئM_���!c}0C����<P��#��a!�[<�&�sȩJ��	jwC�R������	�O�D2%dJ32;I���s�5��-v��(W�9c��	/u��h�pF�����^P�y��b��&�{��,K`�#y*��h (��I)հ�D}w�|ꡯ�뒶;j�ZԓJ,\9�\�~��;��k�9�l�I�0�"#y�g�ɼkV*���}�\+��7:�)�q��񭚸�g���\�!AȔ�K�}��3��}�ycSy;�XL�0�5>�/�;�QZ�p��1a ���I��ě�+�>i&֯�� f(9�u͎��}�a[,��AX���j -��-�iR��	K+���S�-�S����/X�٬��HH���B׫�:�`�6;Z�0�t��A*0#�G-�ax�v���AF��8�0r�9��/�Գ!�k"��,���
�.���'Vm�N6d֍�
Exz0}`TZ�r�|<�����|��M���鷭��$E`S��<_�E��S^�0��'�e�\�:«��%��1-�Z[���N�$�+����.�*�b�gQ�P�~H�rgyf��&�Ձ^����v둲�ٵ�q#J��i��<�: L���r[������l���-��̊8�(��t��c&�0tk��\#oYo��UT�W�+C�d��s3�����Zr���^����J��c߮�	>�=�NX����>j���^\M��3���4�j�8瑸��
,j@�[�2�)�L����5c��� x�wKKo�ȇd��:(�3.�������uw���5?�$�>v���;<�[/�� �e!��!ו�_\-\��Rs)�����=���BJs��q��P�D2�aV���	���jna���͋���̢�3���9��K�t%$+$���i�g�y5)��b���m�6s?�v�S�_-�Ѯ�dl^\W����� E�ϳ�+�S���!��^S:����^G׉�nT�,�����b�)A8�?ˣQ���x�K��6��{x��N��������s�;�aVkz�㼋�	�7"X��U�;��	͖0��+�~H�ycΌ��P' W0��]ݳ֎RL�`ۡA��S��
f�Thu'Y-V�.J��d_(����{4�`g��DPf�ko�y��Jg���m��_6UR����b齨pbB�O����s\�p���]Dh7~��F  �,�`���"���fK�v,�
bil�Wb-�)%ӂW�w~/�s�=t���
'34����~e*g�r���>F��{���4�@��r��j-�Z|L��Op�5�S��j�я\���q��׬�|P���H-�3ڮ��<tD�$���%�()hC������ cA���g8T�`~b_�0ne�q��մ���п\ɚ�����,w;�Lv�Q	靠���x��HE�p=���l����6��V����p����@#�]�K)�+�)k��_>�� �4R\��[z�X`�g�J�ˍ����0��"<��%e���kvm��O$-���;�i��c�`F#
��_u�=���:IS�s�a�"f]�	�\5r%��bF+�Y�.�Űso)Aq2����ɽж�k�5�;Y��<�$�s��GC�K�ⅨI'�A��^��'蕁��	ݽ�,+s��13HNRӎ���ɖ��*F'����V�ӿ=Kd'�F��&�٥_�l�����?��������G�z%�X�9m(���O�&&q̖�t}�A���b�����H����� +c�B`�B,�R�OC�z&�ähtd]�进���`OC�i*E��.Z)w�s�L�S��P�3�dMIy�m�d��a�N�c�Ԓ��X�66^��M�N����#���x��_�!�wZ"�D��qzT�k����h��T�*4c��#�B�(͋�{*I|��˯�.gC���6w��.ض�����؍�׈w��b�g�Hob$�o�j��­��nd����B ��Xk��~-%�enaXKg�g��j������FR��*�6E���F�6��6��G��hFA�#���=�} �B�� l�9��!+��+w�>�e�i���xD)O݋��4�U�~_�0^�������q�Y�^S^�B����
  ��Qw����?�<��>�%�0�^�Jbj����{����B�K��ƽm}W�b�X��@É�j�Z2���[�Q]J&c�i�J��k���Lli�Z��UH�':Di�e����8��$,#�d$}��	M8q?.8�u�̜f��s��Ĉ5Ko7�iox�2�tsAٌ��ֺ��H�N�m��}L!�<F�1�ç+l�������OL3ejD�D�P�'��@�3�yr��Z!�șRx�jhL�=D
.�s6(�<���/�"��F��|�S��T� �&��Y��~��)�KU�V�%�gL=�ks������c	��^��1	�R�1�k ���)̍Y?�Ta�z�g�*���>��f-�i�R+H��(a�P�^��� �P&��#��־E0=�8q?��[z[,��ЅV�y	�D���dSl�l04c��Gk�eOp��
�6;;�\��?`�-��̂� ����] �*��=^�嫣w2���i����}c5��g���Q�/��0e>���u��9�l�6���u��.�.�\��W�v�ۖN��9�/Bj�o}mw���s�fv����	��9p>v��6�髠b�g�w�cI�`�p��M`��r����G�F2�����z�:�ْ�c�Ę ��r��t�"vZ�����`��$${1�b ؒ\�3�ʵ��]*x�w+���O�)S���r���J�t��ֽ�}έ�%���P9;d/�%��A�!�}i\��y��
!���F�#sK�tݢ�ni�j���>�E�>b���u"�g��רC�l�!{��(>ۗ�� S����"2H�����PX��`�}�v�evm �"/ �۳��28� 3~������*6C��ɶ���%�/ �wq�#���xw�\�䚥���r�P9�7Ұ� ue�y�%��������%DWLH��&��&w�;��wz|�H�>��������p#�!��G�}=����l0X�D�X�K0����;�?��LLRX&>���A�ةO��%�<��O���<�.*��PN�~n���9I>i&�C���`���~&��zy��(���B��?QG��g���Ǖ68]9ּ����u}��d_P���Ϡ���}��gt-W��W��˸.���&�j;|Zo}�P�aD�Jt���sl�2��)U��8�p\ODg7n?q�}���O�����M�4<W�HRZeCb)R�.��nԑ��>�\V�ɪ	d��h�_��� GR��	��%�����5�dh���^�0�2��E@ǽfT�p���o�K��a{`�-��{�1'.���+��ϕn}`{'��4�p�J��>/j�>J�C�ىpT7,F�5��+��k���j�+l^t��z[]'���^�U�'@{o$��[|��u�����=QF᯶hnz�o�@L��dQ)#���m� Jy��&_�>88�0�:V���8k.K�v{V�v� Y�2��M�k��P��C'�IQ�LWX��Ȩ2j>Ex����Y� �o�U?A�''�U��..�#	;���Ȇ��maP�1�0"1�E�XQ�>�����?=�oj��;����,�9��X���.���������&�*H茻�+8G�,5�}�	#��������F�D�N�]��CrT�?��à��g���fǦ����׽�w��J�4#[W�����d�6=٢x|^�gu7��:���O驥���xQ�q5��:J im'5վ�p���8�D������9�N ����b��
��k�J6�D$+{P�����p�=zK[i:K��ڝ�|q��Uuk?��[ys�B1��k^]a���/�.��c��#���S�@=��$A�l�0���\[�pØ��)G4�d�4z�ϴxI%��+�5����cOd��Y If���������u���i�Ar�׉E���Ekԩ�JہΨǲ�`�[Σ��w7��G�Vv*&D3N}V̈́��Ab+�(S_��mf�ڬq�&��&�Yn�![NK��U��V�����+�?�s먾�17װߊ�hU��o�O�ߔ����X�'5��K��ծ��g���ǠkFʄ�hg=�1j��mH���EF��52n������/_c�����3:�Ȕ��p��E\���x��5��c��T�>?��QMOq�ئ>C���Z��J����_��p������r�݇ϲ�r�"n2�]�'N%��+�����/���Z����0��ͻ��H�ɻr)�!20�?2��m��a���Ы��k��|�ѵY������NH/R�Ĺ���lk����ìD��j�uj���\5�5�k[lo�Dm�H4v�R�;�-�(�����9V����ț��\i��>ǖ�o�v&9��C����ī��3�B��9���<4��fW�J4R�U�}����|���>'��^�A�ƺ���@���O�B�Y�ῌH�O>s����V@���͕t$�i���l���+��N�fy{�-��D��@���oA���ށ�M_Sj@�J}7�Ӣu��A��îp�?��M����[K飝h�ks��'s�{�m��)7�mt���WEG�������z*�؎.b����6�����%b�ظT��?��Nc�VB!Y�tA:�M�?�Ђ'D����w��+�`T75<�P������@h�\>\���/ Aq;��a�L�@/Vh8�n�Sl�W"���bӍ(~�I+Џ7t�F7M�6�$�m�_G53v�"�z��|(���a�{��U�=`6j��;���hv�mz��
�"�Z9�D���C�Ë.=eb�tq\��=�/��(�uT�p烹f![
��O��^%YA{�8m�=>���1a��zMdt;N6�Ӽ���C�+�{������c��Z��\���>D ���>tf�[c`�~�D��m� ��C��A4��
�q8�h�M�(�M�Rb;��x��IM�ڲ�E��"E��Ve��U5}� �p�x���N��2�|��ʠ��z��'�P_Hgr���(i"���"	��f��L;?ľe�&}@��%s������6����׿C�j�R���x_����n1��d�H����s!�]����� lh?�Ԇq�Z?qVs�kDQT�q��-�K��u��3����g2$�&��D"��{�;��ɸ&�1��ɁI&�Y9�n�8���p]�w.`R:Җ]�w�@s���<���A���Li;��fY���(�x17	p�8����F��~鈍/��B�"�)�|�IwYH�W̨���(,[��^9�;�����-q4�2N�Hw�� wúoP"A�{����x�__���X�Fus�:zx�PqB�M�9�n�y��$�=n��)d��$�Ȗ?�녊��@6��ӏ��ް�5�0\��yWAx��O�\��r�葱~�s4�^������,�����Bq�D �^�9��>V�f#�V�!`J�]��tl�<rS��W���UtUW۩�n轾ǿt�ώ���H��U��M��<i���&�����O����_���q�or���~�g��z@�g
�������򙖽Y*R�}�,[�t�,�)�{�p¦牘�Ɵ|�� �+6������-:��/����HP��6��Fo��h�������@	�$���?�:�; �Z��g�o:���p���5�`��B�ǂ��m�����ǣ�p���4�����Qr!�u1m����n.�m6#aes�k�]��l�k/%H�>u�	=϶�J����φ��P�K�[�+k޵���?E÷n��/�f���w4X�=3�rf�VMO�6�FS�>�mIM���(���Cq�=1ʧ��ұMj.&szKΫ!X�H��5,���Ü�5��rq���:u��u��n���QX1 }�s��T��J�Y	 �"i]����#ED�k�9bo+W��\�΋�c����`~7s��R�$�O�����l|�(�~[;�p�5�`��Zs�a�藎`��\��֐ø!x`���Xj=Z�hk�0SW����L��B��[������D��"��⎊<�Cs<֩����&l�Ҿ�?6 !�{��:���ZT�T*���'T ��7��k2�#Y?�	�o�K^v�1g4����T���m�b�[��pS�l�0��l=_cg6D�w��3���K�r��������ZU�����jp�}��	h%���a�F�/���<�b��UN�j��z���we��W�\B&�oC�,F�4��M�l� `�N}��s&���5�`��jDr֍�D�u{=�P�;E'V�,�}ӵ��i�i�8L�,Y����
�g	��㲲��3\�+�-P����ؠI�O�-�Z�s���J���f3{p�D9�oh[àOH �I��:Lr��\�y�8� 	J�h��u�~!ƤH�
'����HK=Po��<�ن�υ�?��xU��5�E�gFj��1	qug0�U�%g��4�&h�s|��*�8��%�ǅT�	�<l��	��4��f]�:��^Y�����2P��܌A��Sis�1�7��|3_K��h�� �=�1�~x��g=L�����r�����'���2M���Xo,7	n�~�>�tV'��� �	�ȧ�2e�]�h�m/�Y'#�eC-]o�&�tL�������Sv�K\�;_���IW�:��I������^��n�$Q�K�6��Ѹn��lŌ��c/b;��V%}�az�Eq���\�j7sz�`��J��d<(���F���A�S�X͝�ǽ�H��w�X+7
ھ4g
��_=�����E���H>XV��'�h�C�$G8�?'��0-�/�qE�[��&���
g��;��^K���:cODӡ�Oݧ	Q|�*�L�����̫wE9�2<�'�3z��.>�����Uz�H�VP����m����B�:�a/�]c�՛���-"�@�+ԃБaJu,gaG���I�½WM�W�Lu��]�j��i��M�6U���T�Q�z��6�7��Ʋ�Y�y"��Q�3�v)��K�>2��~l��"R`������5�af�F@8 ���m5&�g�&gc$�(զ�"N���b�[����a�d���_��3'�8�t2a�3��r�55�̦��k?\�Ѫ��	N]��͊���(A����h�O�ƣ#}��X�y��i�F���x�	�ףQ hVזP���S
G�/�W5W���#�M �]�:]7����e�=>�%���@�ol������8ę1��`CrP�~8���������h�y��x �S=M��G�.9o��p	r��
�?���&]���P5
@�>�U�SQ�VJ4P��;5��,j���z��%��S��k���w���N!�� ����1̪{��Q�]�"�[e�������U_��,̅�޻�)��X�0b�xl�_�W��4i@Ƶ��e�т� ^~9��_h<H:�(I��>�g�/�Jē{&V�����'���'�~�7M&���M����K~�Q�5�1����׳c6���4}�0!�Iٱ���頺��(�؇a��Xu�c�̚)���k�����l�&/p��&�����S���V�+��[�%Ö��Ɓ���W�S��zo�;� �ۋ�B֩UEza��0`P8ꀲJ5٩�0b{q:�����1�=4_���'r�Vʠ��]K��S�cV�� �F�%��F����z �poݭ�
���J�����̳,��u}���bBztӴ-m��?mʎ�j�W�r��^u�"���b��qdbާP�k�(�̪�Ƚi�t�;�n/����؏�q�C�F-V$���zٰ\8����[zc~M�'�Bl�	6 ��rrZ�%�!�wk;!�Ͱ�1AVC��k���5�<;���Ra�a:w��J������\?�K��K!�����q
���֪��բ��4��d�՗(�5Bc_���P&��45�7Q�z�ؕY�dN��*��Ų,��
~h�1^ߺH�@NU���^��8��nkȗ��6����AD�JU�s���TL���(�hh0�s�u�f���S������ǉB;����χڪ�߳�pc�s�Y�-�F�2/��l��<6
h�wU1��/|���CVX��(��>���1�k��?j�W����I♏�ǽ��b"�� �	�dc`3��i���,�/�"E��v8�d��ʠ$��Vq�u�u͋�
e��Ӽ�eQ��
�iR�0@wi��,8�a:Ӊ\�f�1˘�b���C_P��V#� FB�[e����2i���-^��@�ɢT��Z��� $��"H�a���!]�� Z9���Y�b<ȶ�'���#q�O�$��u���lqr�Q��If�ΙԀ�����)�8���@8&��,�Y_7�w�9Ñg}?��\��U���Ua>+�\B�F޺�aJ]�aQ�F���Y���0EUf����xJ2��zI�]��8σY�����z{{�����-�=��Nz8�*+���5��ǟA��܆��I� �ụ_���K+�?��*f�p^&.����l��Z�Em��|�e�Wwt�_�c��JHwY2�vM�T�Y^]Fn=SA�I� �h2 U���8�C��l]m��:N���t�g����V��A�<��L6���:�<3g�4�ˑj�"�������əƠ9N<m(�J��e���ަ*/�=-��{�w)�/����6�쯵�9O����4��
�!���,��6DD7ȝ��ޮu�8kqwy� \b
��4���=ܟ��h(&?P���v%�&/�U�'��v��$홬�1�g��vt�!z�|(�t �՛5\�2F�Ɉ�a�m�qՙ&ƝcI�Nl��	w㭈A �'3z��VBQ��T�|-��5�b�;"-{/��}�㹮Ch()_l���$�o��y���q���{�o�*F\�y��g��)?RX��Z!b�zξ�"bF3X�*t�q&$��B�����<�qf=N�N�k��Tkz�)O�Gl���є����y����-d��^��Ő�(�v.$�Q
�����Y@,E�1�\��3���Y�v����Bf�)���hH෽���6;�̬<;�g�i��b������Mn4�ϥK7���+ ��:���eD�_����<�b�Ɯ�<�rbX��E��Ciz������_��-��i�J�#���xw����(�o��T�G��/aj�S`����ّ�yC�6���c)y��Jg��u�&ZS�bړ��.#4�Е٥����k�ǉz:D��I�$�C��u,���I��ř���yE@RòЋm�\/Xt�s���ɴ�9s���,�ô}0�H�Y�*�)yX9���m����6��ﻱ|�9n���'�l�Dr+�3�nI9Y�MP�Eb"�Ԅqu��W�J��dW"�7��9�ŵ���a�q�΄�!�����T+;�ٔ��B��T�6q֦���TOH��#fe�T0�z�j��k���.d���,�Y�$"��t�������;쫘��R�"��z���)�F�t���R �����|��9� ��U�B�t��I��J�K�?3��ȡ'�w��\���H ����?c�@��VZ�CQ�ڀ�Y_/�?�G����b���.�U]/�7�/���&O����tM,gu/0��f��۪�~� !+n����yV���� � :���x�9r~'O����!	�hg��y�����[8��M.譾e��MK�w�3����*	"�a��۩U���m��y4��h����Æ��6%˴#��k��_)�c$�3h�{��-C׵Yn���N[-�6��{��y:�_ϊ�y �{���/ط� �݆�ے͑�VK�i?_*)x�Zh,�c	7�0���h��,���0�6����#�p!Ϡ��v��6Y9jw}�B*�t����Đ$|B��Js3K�k�-N�U1���A^j�o��94d[عu�x0y���~W��ݭ)&ֱmk��:�q�4U�"P���y~炝w��;*�j�K���'�]5;_N�>�<ߛv13�V,�)�9��W �-l8��ś<��	!���zn�E��a�@�Q�oI(�u�(߫M��8����U�ٰ����N7���눀�����{77�[-J�W�
:���u�#w��ew����<&�*�*e��Q1�����vCr�O^��^b��V�t�����(*���N��!,��H�F�����7K���Ӧ����k� �H��x)l��� �D۱Qᐒ�_�a:�J����
�?y�L�cP7B��jA%�T#!VB���t�"�!߫��*�x�x�B�u_nD[����x��V��ms�����9DGb��5YbaFy�������/�}uO]��1��H�N	`gf^ͻ{b˼�� -L��P;��$]�<��n@>�9��S.A"�
k�>A���g�ҫ&-��_,ȴqD5S�6�i+�ZU���|w2�y"���p�mj� #ʓ��<��D�TX�~O*p#�J]E�����j'm�U Wn:�2��3
+�8��ΞpweTЄ��W̜Io_���r�D�J����=�s\�$�EE=�8�r�D���ݻYn5�a�I<���t�vU��l��,�%�c�r&����V����	]^����	a-�&~o5K,����D�#A��	9��^��r;���(����p�rc/�l�}����c�����8{Y2@zɚw�(��Z�*ȖN��uG{!�+��:c���������u*:��V=��{ڸFelo��E&���>�I�c�|�u��I�R2����=d���[�(#<��ј��&�]���H]��L[�����6��駇|{S-5�'m3�Lރ�t�� ZȐH!^A���F����,�]�%pi>��>%3�m�w�I���*V�	�O˃ǒW�R����)��o���9�U�hD\W�N*T��Y��j���8�h���~�������f���D�K]��o�;s^C���\L��,u6\�
$�Õ��V]n-���Oa�▫��ٔ	u/or�agPu�ĞY�^�ws��ew_o��;9�#��� p��-���qh�OP%���'9(��)�ͤR�����g��HD���C�6gȫo��Q�N_}��+>�ղg���FB&O��aT����!P�#i�w���
u����+�hl�V��ɏ�#�t��ʁ����ǜ�p��n5[�S��Z��g�-f��=Ⴈ�nN[ j�$�8��w�<F�s�5r1M�1�)��e��������"�-��V �1��ۧ���?����Z$�{���+Z�3��T���|��f�a1����$^d[�12��v�?�jF��ɲ����$R�4K�]{��K��b��v�1KC��V%�s�(F�rP�R|���� �X�D�_D��|Uͼ&1bVmM2C.���z���JPc�h���� =�nq�n��Ef$U&u7���$��*rM�c�Ň<d�Fw�U�e�dA�R�����Igu�ͤ*h�֘9�r��yoQ�ndl�j)�]�2�U�� ��;��Jk������b��}A��Y����UŇ��J�V�3S^I��@�0��U�?VE��� �J�X���-B^9��7�;Jf7�I��*��[��3eS5J]��#������FT���O�%�r�ts|��n������n�> qA�%�:�� �R�_�KŠO1���'Bҕ�z0��Oz�85ցj���V��FX/Hٺ�i��۶�M
�,8>�2�Lǝ��/Ud�gC��w�i�M��M1������B�{�*���\���f=�B����HV�٪��A�f?�V�R�:��R$E�7�5�����=#�U �$r�915��*�~'wC��W�o�P�i����x��+3�}A�*&"st]	�g�H��qWy��ZI(D��$�r/c�)�cS4�/:��)�4��3���2.ī��A�8uԗ���Y^�݀X�EiP��6������n�ɴ�%}��_T7# mx�1Vm�[B�-8仅+�`��u�P�pf��@'t���o�1~�؅����d���F^+�����t�cQ�f�,l�r<?��l*������:�����3݇&�um��h��*����d���^1�q8�x�iR������g���ȱN��IE���|�J��|\�ލ��r�+�wrQ0�ڷ��h�}��O�,�5ɳ0ԋ�]���dp�;��O��v���,ʮ嬗��q�WMИ�dU�R��&`����Ub���)Ě)W����S��"�����7e�mhFs��<��0�c/��!kv�jZN;���3����>�rC�1��*5}V%�K�_V���XbA�t����@�'���.�q�V��K�:1�������;u�L�Ʈ��4I��?�
��21\6?���r���Sqg[-���_�}��)��@ְ�~߀���p�,{�w<A�sSΝ$~+tA�䲂Eᬂt&��;�;33u���"�'8�k��T�Fn��w w-ĥ���,��$Q�.\00**K@�	��c:�}��;%dŬ;��U��`����	ȋ.��&���a[�pRq(��g�^1���������Z�o���˽��b~-��� )~U��n%�#�����M���f�/D8��i�42�����?8������hB�X��§9/�'h��C��5)�����u?7�>�V�����"[4i���~F�y��HOK��gH���.�1�8�$eU��T�D�C�5�:���x~�NW(�����GǏ-�.v.	c�T��F�Nx�F+��>�"��R2�G!�Sh�
b}�CU��S�xs���EF�mrq-e&�Y����dc%��8���aFt�2�Zww�혨{�Q�J����qJZ�{03՗�}B6�eaR"Y��v��1�O��V�nj*�y:�a�Lh��>M跶���N���<K+�����p�Ͽ�M����ר4�b�KxX�4B�������#.�X@�����v��=��b"�u!ИO�yC��f���<_qQ��� ����U���������/�}vg>R,L�T�ѷ�*���r%��d��M��d5H�S�گ��~���^ǡ��	����"��ڤ�p%��A�M�%w@�:�L�:�w��	yv�o�U{UY�.���l�τY���o}���Ձ�Z�i�Z�-�z�B�" ��տQf[�&�l�:�UZ�V��<�Z�a�^	(ϭ~Bk�����u��皳2�5X����9�&</W�}�0���L 8A������2!"H?a��@�쿔V�v3 rB���E��K�ef��l�j�1|���䱖*���!{`ELe+�>p �KD����ؙ/ܰI���f�ǣ
�rH����a�r߰hnZ4���I��L7��:��L.�;�M��A��IOf`k�ͳ�,�RD���}�W"mvؖ9������&2.��8���8
#�q�ks�=5�L)����h�V)
R��n3�V�i|\�#H��@��P�u$���,f͝���e1��]�	}]�zjN�"��Ea�M���>�*U]K��*�w��TM��T�on|+Q�S!���]���n��M�%��q���+ȧ&�[ȥ�;i���C�^/G���kn>\��g��?V�ؓ3ӘS9�'��P�O�yZ�Ш�����"�s�6
�>2��=3O�/@7+P"����I����1!�5	�����%ᩂ�[+[�*J(n_uvԕT�W�)=d��EB;c��a�\A`�,�ֻs�'l�xQ�
�eH1�۔٨�VfU��HU��k�9��>�]�Iܒ'l���T~��Inf�O�>���q�C��K��������tpt^��ּ&�@��P|��E��* �Gƻ�T�%��:�:��,�G|�dy?�[VƨWjd�?&elp+������1P?�w����S���@�ד�L���]!�cY��;��J�{
�M�/7��΍���K�̤"sQ�^�3�]�,��,ncg�]'*�v��N�=w�����;
5�`��/@�2�7F��>z�:���d/s�X	���[DW3�>�YD�ٱd�W�V���9��<;(��^@G��⇣��<v�`RH��c\DU����I�HR�ל!鈣�;Q~.aC},�*nF��à��(f��>=�=N��
���Ѽ�V��\�����w�>���|��8�������`U��ey�O�AN�]���'��r��3��4|���ar�v�N}X=;�lP
3����Y��
ތq��GRIi��0_�a�:�*�B2�c"@A���L:���+�f�!��ay�I�1$(�؏q��L���!��M4a{
��F��`�Ƞ�ccBy��=���R,�B��v�;ڦL�Qz�!��d�v��7/U�<��l(�~{��!q>P�J�v�h��B����2.�"���k_D-��6�B��o�u�en�&��I����/BP�}�:�&o�.�r�&*OWW�N5^N#�&j;I�8Rww AJM��
�p�^xd�y�ň�uO���~����g��=:���jiR���Z�S�r)?3%����|Y�-(�7�a�� �f��ۋ�
&o
U�G����
u2���)_�,�p� HH��	�M^����i��,�r�L����/"��_EJ��Ib�{���> 6Ĺ��u�+���� ���;Z�Q\2o�b0[�*�/ ����9��g�Y��$Vwxz�d��W0�]�d�nT���b=Z!��o0�������@E���Zٝ���s*�GG�����@*�jb��Y��?����9�r��,�BXEZMpp��N-�E�|��� �&�2&���pả�%���:�O��_��o�BTݒx�K�u��J94j�*H�R4�;S&�:Q����D>�h�lG�3bs	�*4���%����(��~�3�9>o/j�6u'��in�| R�j���)�(���	$B��}��B�.��e)��8*HL.��j�=2���P��`�!@�կ�����+��%���꨻fᭊ%-A2(�n�.�~��G,D$6�w�ֶ@nF�T5�˨	 L����FEy���{×`)eP	m���x�U�;9�}%S�dׂ����`׿�����,9h��:á4Ѷ�^�u�Sc���������Z���m�M���1J�+� w�%<�#[�g����X++֫����,�4����!�za�!�e_AXq��6{҄R)�z�/E�?4K�`�$[��ش*k��6)*�;�A��YT,�"��t�C���.�j��QzB/�!����6F����MJ�9���_��-4��0�#��!��_�wY���T�!j?�_��{^嚔��,�O�Vy^E>Mc�����y~�6�����Na�EH�=a�&H<~�*@vת?��$�E�	Bsj���O�(�wl(��[y�ۊ��R �d䊄:��(��)�\��b)�Rc}�i����clXѽkt�2Ȋ�_�ӥσ�lzr��r�EjV�Ӡ/Ҟ�k��̰WoVdXK�r��,'���Z���OÙ�D�=F����01���!�{�*Y����qM�h�0мQ\��1A6i��T5��pdS<�M��(Z����u R �[�G�+9K�bR.5��#�8��ʿ��Q�!�,��H�p����k��)�`+���Y�[듽��\�:�+y���V���j��E�B J7K�8L}�Y�%���v�	Y'�}dkߴ�0��[���@���&�@z.9�$w��镈�O���H�O�FR0@��g�UFa/U�Ng���+|WA[���v��
���� ���d(6�?x�j�"W;ΐ`|�N�>����G���]�m��R<�1�4��&��м��;���/��h"P��_h�u�KCRn||��!<�h�.3�+�˽�'��7\�tai^-�>��b�Ndp�?�71�M*f��a�~�����4����Ȍ{�;q��$ Af���"��gǺip���5�d�Q�~��{�=ޅ��F&�ƪ���\�)*Cs����r^��z�����^z����r14ن�<�bt���I�mm�!>�nW?	%�U��:
B�U����YAo� 2���7u��u�$��T�HIn,�Ew�w��	�}Ue�g�_8�-���IN%oP?�e�x;��W���3f�߶�+\���V>ժRN��;?wӄʳ�|��i�[�}T�ICߥ��q2Ԫ���y{�ߐ���
�4��\�<�r��۾p�k�Ó���q�+c�VJ�I��O �4�p����~��_.�2��q�B�x�X9XXvQ#}���UW�O�͒>w�n��mϛ�, �j��%����Ц�
�E>��}�!��`�h��������q���2.F�r�EH�$khu��s]�>��^#!�VA�á/�6���r��I����Nn�Ǚkg�%�/ҏ	ս2t��Ql��0y����N���n�{шy�`u-
��!%8�:T¡G�Pf�h�Ӓ����Н��_u��g����+'ғ��n�Duֽ�^�6����E�8��
~��*�o��%��(�OQOtb�K��+�G�7��ź��ˮN]�b!��t�����^���+��CF!�D��t��x����w�� �)��w4Uؠ�_�@\����$qe��,�kZ#Jy��t 	������(����R ffŸe�|��z�>� �4��� �b:��.{�l�����A˷��(�"�����L��飥�w��6M`_�\ͤ��Av�g�ȷ�RIi�B]��b�z$"ܥV����tLU���T^�(؂.�
n�޺�`w
�&��6$�'r-~mÕH��?휗�@�4��-!��J�vd>W�l3��^ ����P��!��qfˎ��|n!�C�6]���TC�s��`���m����M&0�fm�O1��'7�K�B[ͤ�<Ɂ�f���@���+@p%#���̂��"C�-DJb�m�+�瘝�L�k0��#8�o��O�0��ֳ����zN?w����x�y����O*f�8O Ab���o��'��o�O���u�ȬQ�3Xs�P����.�9����8Ф��� �����i���.Kk���*j}	+Lb��	/bmT*J�.$�����C�U�x
5v{*�����C��ى~R�^=[�~"�DF�>@�0�ױi�ٝW*�C�f�z��]�z��6Y51o�b�;��H�F����X]]!�S��ρH6��ݦ�~tJ$������;��c��d��� �ђ��ɓ��>i�G�F��Ѐ�.�I>ٳ~.���u��Dd�1g���5��r �����Z��0������`VFҝﭿUo���=��5/����}w�Kz�35@Y�p?3�׹�ȇ�Cg��|Z���[��'ګ��Zʒ�Ӭ�����x�n&��-����
B����\��4��w�en���/�	���yL�ÓV��[��U�������GM��oE��;s��{ſY�e��1\��x8�GgX����L��\�5�4:��N��K��{�4
�q�I���H���@�cp3-a���:��7R��C��k1�<���1��f����t>a#O�=�z^ў����C>	}̤Q.�%��Q��恤B��cj5b��A\�����c	�	|���8N[~@�r��270�ފ���z�~� �p�
�J����ǐ�U!  �&wɶJ��=�#�}Wez�%�UUh��8��)D��:���_o���X���+P��&��&�(ƀ��=�]NV78��iC�����7�MNSߘ$z��PP|��Y?�	gry�D�ز\�f��&���dt�U��䯫K@��=E:� ������y��!Y����~�ۉ��E�f�����U� Wh��*��������E���b�3n���S��V<G�I	�oC��*��'uO�� ��
�nZ_�jr5u�3Ί��;�?b���]$�@/=��C�Y'��&ܜ܏"9���������sd����*��J����,��]�f�{����;����^�2�WL��3�9��/��Ծw�-�`/D9\�l��[XGw��s�@S�1�_=�^��2`du���V	֊������𖢙��EhM̴����A���	��,'�GL�W��A�3����_�%�'d���G�obB��
޺(I3$̵�|���XV�p���i>�%�{�G4hT&z+D�Dg]�?�K!s��W�zT�����Je�:�6�z�Pp���ۇ	za����$�
�x�~߾?�2(�бt@��um_��e���j}<9C�[�7D3{Y�NI
<2:��i#�_H���#�~��a�5�3 ���	����,f��b~�E��9��g����;�߇3�2�:u������!<��P����n���͚���u��N�w�V��'5s>I/���ḟ���y-�C�<����`�EM�g>o�+f~S��c�����C����>B�ᇘ�n����kD��W�|Ϙ0�6���)����ɛ�<\kD�e'][Z�w�o�i��-��q���>�&��[)%͵�W���.�u�p"�8.��^���P�������{v����T\g�~���+1hi`Qj�5����C�Fѭ��,Z�5��=S�_Q"��Q��.UO�z�����(�85�6K���ݜ��`�G^� @�楰��3S�Y��7\�.�O��&�;�[l���^?F4s6�E/��	�SO?��V�<H�l8X��Sx(�[ش�P�]�g����2q�۱1p�8�2�y)�t2��;�/��%�G�v@$A���,no�h�"k�o�*\~��ּ�6~c����;%̆�$���ڴ��Y��Ov�ѩ�D����!��6pe�g������3��ͣ�����/�K�.=�a�K��N�':�*��������w���Ź���1��L}+��ÿNgE	X@ ���>ɡ~�je(x0��;��8�hC3�o#�!�ܠLӽ��]���å;����q�h�3)�Tϣ�{M��ms/9i,�[�)�D������6��Z�_f�"6��>#���p�뺼��n�%�6D����*~��C� �A��XS:���T�z�)ɲ�FfH���mbDy�@�~� E$�j|�! Ek2� FX�x:)n���N�#��t� <�^۳�k�3����~
vFh�s;�ٞ#EK��m`�#�T�{a��lPUN��Q��.�Uh��Ū�k���A�4����U��	�*^�x�R�\Il�J���z�L�Vf�ަ�I#��nc-�sQ��x�膥Ď(@O��o�f���1�����qƎLi?0����$��S��d�8��Q���3Ϻm3�s �T�)���O�$ސ�!_�^�v8�W/��m������B�`	�V�,�,@Y2��B�7�k�S^���� �7)W����Y��R)rсdZ�	�Ө�:>15�v��sP�;9i�Da�@�ibQ��1)����#,r U��CC|�L4�=�d�z	E�q����E'��-K�9�����}� ���r$@]j�;�}��)�&G����>\y ��i�H���.ѡ�50w�u���]���{O>�9�2�7�Sܲ�ٟ3%"O�ETm��C��*�훂\\�wFt�=�%���IU�����66���:tk�ɽ �%|Sn2�T��j6��(�����try�w8^
~"@&���!���v�
��i��9jw���	��c�M�;���"k�AC����<X�Z��X~,�Q}����UgP�mV������M/�H���y4�>�oM8A r�����b[�����M��">��g�}u;�R0���_ ������)�Y*h�Cv)<��U�u�
�'�����F}ٳvl�j� �R>� �Z#(�A�Ч+;�'��Y�K�����8D��e]�F@K/�.sV]�@q����e��Q�I3����Y5���t�R;�K]�Y��|\��;Ԥ3FQ�$븵\�C����W��c@�}�X�W�T,;��&׾��\��kE�vځ~g�h��ڮ؃V_%+1J^]��{p1-����������=ѣ3��H���3�/�6�<����ţP����j]���7a�ɨ�����.u?��d|�� ���g��}� Ͷ"��E�+���k��TŐ��o����&�z6����=�H�1�N��wY$S��xǙ����qj�;��<���7z����w<u�����SQ������c&:]��$��ߠPa-��vК๝����V*�����]V>��,ƴ���7��vds�bP9�ul]Es�]D.��ji#�Y��ޫ@!{i�~���ſzڜ߿��J�x��%��cI��ڂUK�����!^�,l�ʳ'5�.�g�w�������М{8"^� �jMI�R��y��:��T�EXL�=R�UUB7��.����2b�6�������`S�|�0G�����V���r�{ؼ����1�fQ��������<�܌��Z>��4��/��E�Iucs,q-�\Q[]??Ƒ=o�U���:,MEs�e ���9�L���s��U@)F�R"�/�7z(-��/�B['��z �WN���T2��ߕR'�����Ks�<��r�������j���g_C|��O�2k�qO��F�Q�"��u3s�v:�q�ԶU���0�c[�IQ�ر_��h(��w4vW=xg�-���Y�v6��,qR�l����!�<O�W�bI�rʥh.Ƚ�D�kCs����1Bz*K7�4A���^����(�rH̵buZ���۪�$�M�Ɠ�F�q����;��&s�Xo>�i6U<�g���R4x����YWc�n3�.yV�#=�D�9�xv9l*�:�v4�c��DR*� V{�ACR����'+����	��c����� n��^��m��-�>"+�;���v'zNp�~@��ʞ٧<=����r��I��yD�}V�Y7qy*��ͦ�p���!P@���oP1��+J_��'���N�-�D�c�+Q��!�������F�+X�G��ǵu<�l�B��"�e�Ds�A�H�~��.�-������x:�;��3Z�D^]�o~��20���uZ=բ4�v/���jy&�Iqf[;B��{��Pڇa�M~EK�<<T[�oZ��c����NM�����Y2v��#��hLSN��-\�ͦ��ˤ����s�(Dh	;�L�Pi~46<���W0�J��%�v�~��?u��!�md�z�
C�������	��l�"I��[������^ԭ�VG���\>��$>F�2�;ܞʾ{+3Aq����5;���n�k���o�]��V+e��ˑ�S�������u�i�����:�봜���<�<��&Agjpn�W��M���Ff�ܽO<7M���ߨ^YUT�4�0����s}�[�he��DpF��:����Fnz��i@@C�Sys���)\�7sq��pn=��9{�E�Z�.Jgub/ׯ�%������C/Vy4h-ߖ���Q�	xe���3�Ŀ�_z�/�9��
� ��H2|%	ؓ��8�x/is��8�*ޥ�Ǹ�`�L����6���!=
�U=ܗ`���d�1_jp|I�D�W���ma �i���E,��Sup�c;�����3��M����Y!�z�~�L�ma�d��~�>���� G��}�W�靶]/8]�|��.�<z@�R�=���'��L\گ{���7�J[R�i��G�D�l����&���z�F��ȃ���o|A ��S�\�8/H�C	��/��+TA���g��e�y�5�O��!%u� �x��;�i���2�>�A��<�Č��:m+���8xHRw���}a��	�9���tDg�G6����C��ݹ�>��D1F����xt�գF4%�髉QX/�lq��KC�w*���{�)^.]���BzE�J��G����������N��,���,L�{Y=��'�
V*:b��C�RÌ�Z+����r3��l���ϖ�਋i����]�"X5g����#)�ڃH�)�Uك�{)ܩ�,�� /�Y��(ez۶ ��#О'P!vC���u��ce�uA�g�E����"M+4�ʤn�U�]Ya/R�h\�~De-p�� $��7>�J��[�	�H>��[;R��d��$��''�@k1۩6����릱RnۧN��>�q�3 �?,���CS/͠���r�*q�b���73�f�ɵʓq��*̲֭�N9E6��jb[�h7�F����:~��5 [D3��3�o,�[����y��~&��Y����+1՟��}�T?+����Y��p����<���.�n8��]"6�H��Y�f�����V���Ͽһ�]����͸ˁ�1��f֫$m�䍯h�H2���C\���_l]�4T�p�O�}R1;�f0�)���}O�j�Ȼ�F�e�^"�c8�s�	Od��k�%bY8��#����������2ϟh�	�P��������5�Ƿu�S	2��ͱ��4,��9����z�`�mr4!��}�RAd�N]VETY�_'�E':�=�
��v̇��,f�v�Yuj�켣�p���V@_8�d�{��e�UT֍�C���_j�r��c��l�'�|Ѝ�+�ݫ��? t���@���\d��K18$I�BG9v�'�T���g�]��NO`Ob���5m�b;�6��7��Z���!���ҷ;�{���x�G��)����}�.�Um[d(�'p�Mx��]z,�����z��o5Gd�@G��?��߮]:�vxY���W��йi�΍��g>�}�T��`��f�b�@��{C�XQ��"],l{h#6��L.��k;6g���q؃md���蜌8�>R��%�d��9�2��M�����ɣ�#�nRσ�37�i*M�GGN��?��âY���t���z-| Y�In�/��\[-P'�o��N�R���`f��E��y�/+�̵٭r�&	D����u1w����\���o�j����h L^��߶R;s�0��\��Ti�>@Ӽ}��-�r׉��ζu��m�[RI�2�U��tE#�c�&�*���Q��E�SץtT�3t�?ה�&�u:躪�^c�9$Kӝ7��St`J
��0��"S�!��ƈhFS��
JMW���TS>$��e�m��qE�J�)0����a��?nŔ�Q �7��yF��J��g�dޔ������W-H��ke5���ZX�dZ��(٥V��6@�u,��	]�V�q�x�X��I'��}H�A�r��ٴ��ڎq���ƾ�����	����g�=���3��"Ǫ�@�
��8��`k�P��D53�P�
�# ���*O��G;C��S�V��WKxqo��߼HE�|����w�B�M���+�F��]"�+yQ�?9M/��_8v�����c� }��T�)�M3{�^�	�b?�L�A�`e��8x��)�8�$-�`%�b���m��d��q7�q�@g����is���S����VL��cs'��jg�B;������򬜪_��D�d�m��Hs�����n�C��*���8T�R�$UG��;/�Sy��>�W���G4O.����pUBȽ�v�3*��	���Ȫ�U� O�r�#�bwꕪt�D��
�dǣ�֥��W|��̓՗/�jD�f�ںN�9�ѥ������ 	D�'ó1Jt1�γ���fYE�N�;m�q]�;�+1д�V������!c`)���/P��^K��$�y�u'�H�~�Yk�2/x6ؓ�ź_L�\?Q?��7j�-z +��V���9�9�=�=V �Mqɩ�;t	�����p�f�,��]{ߤnX!RB���F�'�` ��xO������p{�W_��1�.�w��4�H��1K��ڙ��1�0l��]���r��ݒ'�n�+���֔�߈o��!W2�P���� Ke�us�!�u�L�;�P��j�U$�����[���f��[�k�~3ͱF-�Q� $6�p���\k2o�E��
_M��,����n�+#�����ېN6y25�k�qS���Xn�K�I,���h7P.�Ĭ��%���a2���Q�*��
G�=O�-�΋'�5��rw��9��*s!b�0=�#S5i��Ģ�B���S�Q֦X�D޼�$J��/�$�p�˨���3U����y͕���:�𵻠�l$��дᾑ p���Vm&h��}��7���һ����b}�/RxU%�osS}�b�24#��Gٓ��;�ٝ��*�0o��[���/E/�+V?6�]����:A�BC����.g콹Jba����K��i�;`��y�B��k$H�H���v\�� X��];�ӂ(5+��O�57F/�JKz�U��ژp��k�Ș�}�U��J[�A�{$T�q���W�����vd�cڤo^���x���c�%��/7J*'�������,�aϨ̓w~7���4=,FX�KLҏ��5�q��*PE�(h�З/��������H��I������&�>�� X�QB;�bR���9�t�Y�ӓ$�.��`	��e]����r�?�¬�zQx3a�qF�Jy;�kjj=Q�qqM{	#�:�S�=���f��Z49m0.]bi��� o�jH�����S�s�e�s�m{Xh#o�QZ�bR!��fe�
�SZn�>�O{���e�� &g�%�?5c,��-��B���q�A�B��s��8#��NM<��H�	�$��8�Km^�3B�D�\�6"D	�⟰��;ac�W��L�:E��~a #Ʀ5�����G�=x�@P!ju=�k��1ΏD^6n�D#�@�k��#r�Q-f�{1����YE����'KTh��3EAW,��S�l��n�⮞�����u
��nN�WZ��3͔-(M�A�Qj܈� �~T�S����/��B���g&�ɡB؉�ENUy�#e�F�RB��=@����-�⺧�%�̿U<���x�+K�{E�
t���z�(��0��n�<�^@X����?Pt��آ�����˚&)�`ƍA��l�y^uZL~Ivb�K�.�A�y�E�q7��x�n��?��V��#�Nn/�`C���F��X��> j}\�4f^ye
`.`O�HS� �!~�U#�=���O6l�Z����q:Ԧ�9|
���cTyH��?�so���$�U�厩^_�$�8:���9Ȼ�xD2E��d���%`P�@c���������Qd)Y7��-&^J�g�=س����Wf��ELآ��Z�ld��uA��^�n:�29�>e��0�E<Ak�y�CM�w~�N�ئ¯�ޮL(�}��3�'Ne �q�R����ԑʶ��x_�0��@T��#̦��s�q:H�`k�V���*��q�_)����:�<Q����/FV��#qЗ�]W��թ�� 2�,�1`Y@p�^�YWe�z&�*��5{� �{��W��gLɷ:.��~q������_� �S��,6����S�?c����q���n��z"�6�+���Л��P�=el�4�U4�;/�7�=%�����9�^�X����.W/��k��LpW�R\�ʼ�����»�L�&�g�/G��6[
Pj�K��ce�@qw|�]0.�8
�?�1���ϖ[�
qXD�Xk��*�Y���m�G��0��b`�-^s�/�|Ǌ]*�/C�Рtt�R��S�j�i��*�m�o��w�z:���un�f�%408�@�S
�d�]�W�B�@���*���7#��Q��h#�&l��E�>�UB8���e>���^H:{��*XGS0Q����r�zx�;/1o�)4p�iK������'���[���"�,����J%By��t�b��6��#����B"g�d�X��ů���V���U|��^��T��ƍ-���!�v��h��"ܷ�$��
o�k�x���k� �EP�
�O>V��ag��'DZ)�����`	�,�,���y}b���Mp�7Éswyڽ�.��O8��)�b��F�;la{y�4&�p�,��^}�Y�&˔��ȴ��%>wY�iY��/t�*7�:�OX�w���Q���H��
J����)�����=b�\=�fH��������k��n�VB�V<p}�Dp#�>4Ժ�}����k?�DŌ�X2��z�u�F��+,�\:���
{h��~�]j#�K��c� c��4mRhώ��_K{2B��R��m����DT�b+��_ �0U���n��u���+p���5�6�~�n���M�d�ʤ�mC�OO�5����kп%��ga��\���7�c�n�I��4!:�덬R���OI�1�'��o�9�%�[ظZ:�t���?�q��jK��\�u��~�s��0&�@~��7s�1��y�i���<�H���`A�W6��Ϗ�W#��)����Ա/7���2Mq/Q~�} �,�T'�a�3M��~Yp�Z��U������R2�< �jd�v�ݴ%�M�XQ?���L�,��^5���IP�l��6�%����E?��Q�ؓk<3Z����*�X"����xk�^�Yn�Y��6��g���'%h�ihKH])L�4�L�H��|�	�Y\`I��5�NY���b��p�@&����� ҳF�_sJ�0  a�5��M��,�ِ�%�ACT�2��Ƒ����[A ȸ��K�!��93��wn｡�r����8I=�4�}cO��_�@���mw1�{��BC��_��v0��.m0��7��a(7�:U��ֱ¸�ξ�8�X]\���yP�H�%�+�D��#������;	xޡ�Ipceg^�e>�*CA�����h�^#f��r���z0����s��+֕���N��Z�󨺝���q��"���+ޘϛ�\Z���i����K�Fe��FH��h>��cOJ����u2�h�!q�S�Ķ_�^��.�Y�µ0�#g#]��A�$�&qv��m������p����Dpj<&��l$fȓS�J?G2���u� ,G;/l���M��(��H�³&f0�n;����C&t=�m��3)󅕜>������v��ߚ'$�6ˏ
Gy-��@�����w����1���i����S��	��M���U�� ȝ(t�[楛�ko��	
�!��!�,6!��[ü�b��WXy��mV�m7�^5�z�*/�\�8�r���k��p5�lF�;3K6|��oJq�)^��:���h�S�"�&��:	*�6"��$�.�!����el���QI�@�X��M7�R�*`T,W%�-��5��/R���}$����u���ҩ�n���/x t������U����C�X�W�6�x���
�%K7��"ƫG��ћ	��!��7pE��a�U ��!_����U<�5��fЊj��ԫ�M�<?�t��z�bd�2[GLZ=�V݆P���R���㫥a�_�,1�P&�Ș��:d���gLɴF/��4�����t��d�6�-���4�~���B����*[�q�S�u�@4�;͐��Nt����bl.��j�����#7塳EE�B"t���Bі�Ћ�lo��{g���$�=C^��-/^. <���am��b�`U=�ۼ6wnذ@ӵ�I��\|��ԙ��\�_�����S�����|J&d ���� "i������*V��"�@��L�v�V�"ew�&����$�~��SɅΑ����	N��!� ���nI,��/=���Dm���P�}��YWĤ8g�,2e��Y	�8�r"<Byq��$�JPl%ct�/�:�ߊ�m�l$��4U���.-Ҧ��{e�MQ�ȑ������j~cˠ0O���u�$,�2�X�ԧ�$4�`a�����~>fw����h��;G�w[AY��2�ת��PM�O�ȣ����O�yѓ[��b�çd7EQB�+i0�T�?�zJ5�y����� �ɶ�HR1�n�֚����h)G��T��B�>��ܤދÁ�|�'�KG�h,���lPvl�����^���ם�0�M��q\��Ŧ�Jt`��T�'US�|5�x�;���QJ���>;�=�i�f�`�,�9ǻ��4�agLN<L�!��eI�[��Z{�^�C��t$O���dѫ����r��7$�udA�p7�+�8.��Y\2�C0���Ȁ|������4��M�-��bo�	ͅI�"\���Q���=��P%:m������XcQ'*� y����q��X	���n�k�vK�� �k �*P�]���Q�u_K{g��fo'��^%��AD.��Z0-$j5�q��Is�^a�)aN>w��Q���ip/�z����.��8��u昊a�Y�`f5�$w��LiC	�F�/� �#�u�T��4]�h�Ǖ���I_�#J��JO�1�wKcI}ܑ �ß�hV��D�i�2��&��%��8䈗;v�\�6�O������O��F�z\�\�I�v���!�r�z4�����z �e.�'!�v/h��$곲lp���i�m���t(��ߛ�٫ߛE]^�f�&<���qL(X�QK�+
1ج�(DJ2"-�3L(~�I��9.�ٶ=���S��R�M���)j5;�;�]�x����م�F.)�ר�����u�+�'w mLi��b�P��&���C��
�#t���\�}#�S�@�7V�ǨZT�X|����2��6�)$��9�A�\wtÅ���QG�@@��Ւ�_�@>f��Re�e�	�R��yWe�4����,u[�s�7շ��X-�Q�ml�p�˲����<dk����G�T�AW����J�u�VN�Ŏ�s�8��%[��K�`?!`�-�d�0bV�	��.�'�mv3�Ꞗ�LE=��)a&��M���-H����u0���t�u�� ��_}�83�F_�i�̋���v����b�?�����f�j.�  �V��O^��^*�M��F1�,T-{sN�Z��~�ο��#(�?�����a�3�oie�]�m�R�Q^��S��_�8�Z��[m�
0a��x+�0��y'�OVh޿!��Đ��W>��U�]"ת��� ��	'挿����wxϟE�8Kz���nwmЀ?�[6�W���u<?�@g�	@M_����d�1�6MD�ʁ���X�	�^�
�q���,h�8�=D:����I�uG݌���(9�<�B̔BA���"]sa&�s����C��L�:�G�!�o^\�p<i�ː7�į\"
�� �ա�r����y`�\C������%Ɗ{Y7D#'@S�{'�m�5����M��@������E�*K�歧\~��5�K��sB��f_o� �#�iobTj���# ���ar/M/J�\ӟ p�/��}v��]���iOjR�	�L�HI974:?¡�o\N2(�y��\t�t�m����d��Utt����È�������ԃ��x��=Q�w�=�R�;z�@�}�h��>�av�9�զ�F�@�	.���j���
�u�ࣨ�t��l�@�bKd�!:���r���֥:-�*}�py��r7&ғu���)�!�����u5���>�5ʏ�M��*@{�
������$�I��1��w:C�$��,W��H.���dp�Q�I[N-�߾����1�U��Y�A�mS#�*���gtp�+ˇ��3rI,�t��l7��e����n�*���Y���b0V/���.��o����4#%�\�������Ј�I����T4h[����FU���4ݱ,Zv�����.����D��z7�eO��m���q	ky�;�Տ[�Ǻ&r(�����4�������Ն������l^Ư������>�D�'^�H��ol�����=b��Ev(K�pQ������
l
�-�q�ɫ�Ef���uq���Z��KT�3mg7cǡ{�N� ��w"f���Q����QХ"�?6�k����Dl�}������a3��5:f�͞p;Ě]��p�ct��1G�����W�Im��j�O+�p`	`,P��37��S���¹]|P+i�Xv��<k�6�G#ˢ��WT��{	/��;5x�@Ͳe.^��3g�|8��G�.�lz��
@���e�Wm�yu#Յ��F��|(�@/��I��{�1�	�&�B�ӰX��&ׂ>�D�'�n@�<�O(e�%A�̈́C;�	���	p:�h����J�m"/pv���̄�n�d-*��`e+�Q��*��}g�(�oz��[�/�kVB�ַZ�
ƅ|�lb�,腉�^8t������S��yi���E�Z�!M�ᚊ*���g� _2k̵�B�6 KHzVb$ܥ\�7��T��
�x@܈%[Nu�b\PW��7< -��ԿStʍ^R4�Ts$�P~���q@Ɔ���wQ�DL0�G	�~�e���,��5эA���7�xE�:I�&hyH���|'��)r{"���i{�~0�\}���dJ�ʋ{
6��tA��_!�l�W��1*;+�v�pWހ����!H�s��E���R�9=>M���P'X��i�H�z�g���Ԥ��OD"���i�1}V���J�Q~O���y�p�;Y22����p��Yf��}�&1�6�U�^��>�ٌ��)HZ�(�h�Up�>|.��l��220K0ߖ��8�֩C�$�$+�;I�5	����X�����.�7?j��*��|�B?Vϖ�'��W{�)��\]���˾�����k�o����ҩY��W�1��q�0FT���}��~��'uQp������Kl�+��AXD{H�n�o��:��_(�h���Ӻ�-��QʣD�eB�1��h~񨚏�G7ڧ���1�@��3q���.(����@�N�9&��6pY�M� �H��Q�����rB��'���3e�
M��3��`���r3@'�B���T��N��;k7�!�Q���N�,5�~����<�\)�l��_%r\C�xz��LLo�g���^�A�=b��$t�_c7��Y��j��7�hgj-=�s�j��,}b�?(ܨ�25��
��}�X'���Io�}�h&�������bܸc���G����R"�e�X���HE��'+�g�x��k�|�<�L��I3<��̤�C�DD�a-M�ȁ7n@�N~�ޕGDH���h�{ڝ��D�)?dI-I`4�����ʲ2]ܮX❼�4n��8�u�T�Q�(�@\�I����nk0�<(Lz{�F�y*��$����~��g� C$x�$j'���Q��UN�����v$����MXì�9�˟�@�2�7�bȔ�Q��6��	�Ņ�hwwCvO�ת�g�$�=@��-p�M�u^/��5��VE"YI��M���J�p��37B7Xt��������%�9����b>�"\HN �HO�$����%��F�}����1������2;9��u9D^=p��ذ�A�8�昻��)�$�д��xO�%t�[��_���$�|hH�,w� =�#�V��s	�M�4TSrk����^.E�7��FƘ����:3�zla�|y�����g�rGOz���]�:g��#9�q|1�~k�@�������$J42������Ɨ��� Sל�FqDwZ[|��K�}?)M���D<>*D��!s^d�Ytv��o�l�x���yU&m�z�}}[j�l�e�s����?18.�2��B0�~�>{S�������L����?f>Tx�Nah.�3�9D\B\\]����������[�e�4��?���r_Hg{�O�D^!���t�܇���o1	��H��&��^G<C�m�z,tᐟ�����(m|��^Ңo��NH��X!�Ч���S�h���N4�75͜���d1`�1es×�H�!^��|�A��}d�6�q��v^cTP�܃(����;4�5D�>��Ua�÷�������m���5��Ȥ��c��md7���zR�	{M2�-jyj�� �]`$+�lJSD��h}�W���!Ͻ�a�o��溺ދ����\�����G3�j�4�� �,l�4�ҋ�*�.��owI{9_�*�n=?��Է��x��L�Ԋ�ǰg�c�\�
,�:�6'�	�_��^���ˑ�t�'�h�M?3�
0g�� ���#��V�݇��w���=@�1,���f�D�L�6Ք̽/��[4��	<��d7H�0��T��J{Y�X��%�E�m�i§��wU�axÉWh2e���1a�0���֢�D[-�O���B�a�ً��̉�.��-�FQ��'m���7�T��P�	���+ދ�)�ۇ0��|\a���Ƹ�Ķ��쑤s)p�kԔ�ɇ@�6)G�Y�}��e����~c��t]s�v�p�&$�M���D�r�(�g����>&:��d�*Ho�ʲ�b�q�B��ʆ����L��Ȃ��	��Ae��C�XHh�S��T�7�A���}U, (0�NA�^#�x[�� ��ae��Ns��5[�G!�;v�uM�@7���|p��'P�j�s�DesJ=0�E��v�Eς���!2�2%�ovo�3��+տ�Z�${���|_���y2��|gbG���L�#Ȫ��j����K#���Ӫ��	cCو.��&o���9�8��U�=�y����\ �]�L�P�=2���q'f�\��Br3Y��z�/ڮ��������q*�˰nTZ>��^ɧF/��M�ݳks	���|�6��٪�%s��-ބD$v��Fɮ*r6��1�غ���c�BwP�����	���&��ݶ��I��`�������~
j�?�����-����Wn���l��2���s�������<�6W�\�CW�����e�u�@6o�o����D���(��l������Fz�Q�$��.9�č�d��V���Tm6'��
�?ƨ�"�DF��q#r1�ٔ�;.$ee���P+[��\H�����RiZ���\�K�t�W[-
��Ȇ�o�������l���N��e�����rw�=���#�¿�ޚ6�W�#��J���&Sx!��[�-��"����6ݞ��L9�'.��q|������Q!�V:�5�b��7MfX=.�/�m[����n�0UՆ�_

� ����{���*��ﳴ��V���v,��>on5t�R��w��C�ǣb�M^]l�P�y�9��b��ZT�>�3����x��m|bI*�"�+���b�|�m�ɉ��(Tą�먙#ͳܺ�j9^��3�҂�J���np�A�����i띞�4 �]�g�%8Q�����WB�AJd�N�sz�À��
D��BX#��[!&x��@������B��X᨜g�-�T]A�4�Z���C(�ZۓH�&�����Щ��>c� }��Џ��őpjY��/8m E;t��S~��t�1�J�jl�>��z��A���C;F3���j���/�=_��PH���0ELi���t�T��g�V����ܰ]*����f�ϑj<.d�a�m,ٝ�݉)w��KC��v��_xԫv�h����z�N\��ͱ >�־W��R�I�|�de�J�{����d�e��3�.�z䭚�aʽȸ�^Gl���jjP�cK� \ՠ�̶�	�TOPcd+L�M�ښ�U�hƣ�R�O �@�1q�p��a�u��f�і�7;i��TDZ~`N���"�jM`�B|�3��˚sF�a��փ�~�t���F� �l N�3�9��>�l�͡��?�'&�y)��,I����LX��R8Σ@�L4I�C��pguU����ZB�
'�Z����|l���LE\�.�h�a��\z4�J���W.i�+�Ȟ����@�|Wì�xx�&��]"l��tq>����qx���5ӗ����Ф��J/·Ӫ=vg�ɉ���h���蠣�j�r���H �0��._D���/#����k�n'��.r�j��u� $�X�6�l���7	wbD�%�2̃ܞ�O	�'�ϟa"���/�ֱ��	$���h���� #��B�],�%�ck~��&�o0jY�ԥ�s�i\��՟E�� ���"9�r b~p�]���`R^��҃j�RW4����/��'��gT�Cp��T��Q��l���LfI�����vydw�u0b��fXP��&ƨ�7B�ɖ���}̯	xR���>��k2ϧ�"�׶UPE�k�W+�e@�08��I�,m���Vf�����s��م��H*�V���8��ZyF��$�[�h_�Z��U��W�H]��ܳ)�GM���c 2�+���� x���F�*��D,�)=����U��J�>Z�����n��ha