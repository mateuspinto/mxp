��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���x���h�v����Sh�-��E��ϕ�..͖R�젙�����S�?��o���C���'�;e����ז��=�UC�{��@�G��͖�Z�eޚ�i�֎$��$����:ɒ1#q������&�0�`H�Xb<�;���;M�t�M��#�dؓ�y���[���J��ս�R6�q5�����
P}��Wb>c�0|QS�������<w(� �@�:Ez}�L��j#х�'Vp�#h5噢{�o�HQbЧ����a��m��6|1����B��V��߭�� ؘd�Z<T4�qZN�0��
	�Dj}��l�}be�Yۙ5�q�%�Fݥ�b��</or��#���F{'�D��/��y� �,W��~��#�:r�Wׄ #��M������nH_q�<�w^Y�DZZ�l]\(�0���5�ԑ{���!y]ſW0�\ۢ��^�h=se�`M�'��wf��!yʁ��,��E��i�յs�i]�2�"ŝ�B����m�M�����O�r��P����2�u,Ft`J1e�� �zhkס�G�����Q�C�I4غW��KXN�7���> ���B_���N4)hGF��`��c�4��kc�%/����"�Шާj�E'N���v��1	�R=�f���n9����Bm�6�+��q���|v�=��[.ƾ��4��`bq��Ә�nx�!2�!|�R���0�'ūp�Ĳ��@�9�]���P7a�kJ'`���W���8��t��S}�:���'������}�N��"�w�}����}�h����Ch1,�fb�}q`�i�.vJ��x���G�K8i	����O$�Ʌ�"wɉ���X�5�z�U̔��AN�\�1F>Y� ���/|��FPl�qx����Շ+�쮌�2��k0���+�xj�� �W����B}Pʟ��z�q��@n(��)G8qk۲����B�HT'9��b/�ǖX��-IL:Z���\.�c /D\�?x7�L\j����;��G�o-��s�0	�t,5�ax��kML�*d{��x=d�����[5��]�[I�|���|�>W��Vj&b�i��}�~Ph?;?��ɼ�Ϻ1����>��U ��l���5�Rpb0A�a���m��Q'�Е;I�2�q6SʯCJ��/�n�"l�3����)�>������0���-���O�3�K A��e����mپ�(�,f�_��R\���E�^
�DM��7�' ��KC������#s�oٳ�ׂ|�l��@�K[�hH��m�)? ���{�wQ��;�ȹl*	Ҟ���_�������Q-������cx�]Iǁ����Dvd�)o&5]RF;���+���#�����M;�Q~H��>�8,�`����ϡ�I���(�?�L�p�;�߸�%��̑m�����2�E[��+�����:u�-�&�a_����P'1 �էJT���RuP��V�jAU/���{\�HC%�=��Z'ΰ A'���`�p�gغ��1����ŀ�/Q 2��ǔ.��;�&�a߼j׆�o��?��x��^��"©fhoN��MX���R�+	GI���[����ģ�qU�;踬}(�hO��F���x��n���=�����o��FYd�җi�/�G"��ʝę�km'@ R�ٮ[uNH��·�Ǡ�3�+�X�>1�-�󇹺yvH����7�q
��NM����(���u��9e��� ���M��b?Qq
&�'TW�JJ;6��^�:�^:��a,l�P{��4�1V�@���e�4oA!d/:z�
ȾB@��k�l�(�iEN}�O��k�m�NH��<��\���FI�_����g�޽�b�����<�n�&�>�����ƽV���Y�Z��l�Άp���h�2cdB�$6�&�W��j?�Tܑ�q�T�M��~{���-$e?G�P,� {�P�����m�+͌o�J��/�׳F-�<CYA���R�`s٥(�n�ק粙fwnz%���w��Bٳ����ħϖq�2DB���!,�j�][����.�4�`Sꅾ�|��C��D�(�M��$�D���%�] rm�e�+�?N�:~�	R	G�꓂���%��2o Ng��)�N�摉�- AXl?�L�z�1��%j9���О�P[�_�\)�X��1>��6���GX�n}��S.�%Ҡہ���DB��%��B�݇��]b�;��A]��vM?�WI�z�n�\Oٔ�hq*��[y	����Y8d�n�߀��\���j����@Aq�2��j$ﮂ.E��7ƉX1x	���O�0ס�;,RY\^䅽%Wb�=�y�;8i��4�<��ꤔ���pJC�X�r#���5�:}3�-��k�b�{��W.4�K9Ԛ�]�vc!����vs>(��溫:�-F���*��g�t�� ���M��A�Aٹ�U)A��o�ј8�;;�>�t�{Jx�i�k�n��~�N=-���>�S	.��zL��/ޮ�=���6�5߉�3� �u�]�T��_hD�]��#u����β��Z�/�0���A#���L,�m�	�������^@oܰ��ŧ�
� �E�☆)Q3�� ����+M-J%z�.7��4r�Y�|~�p��0����XC[���c,#Ǚ�6�Ӣy�^���w�U��6MΆ;i�&6�WYx���$��y�C�.Ɍ����,D�� �h�2)`r�x&֨eK{�kP�#B��Yd��6S���+\���B���d��sup8E��}�^�����]لG�uJ�'��#5��T�Zj��ӆm���!ВT�o	�(<\<@�FiwQ�v��u��;On��嵕�
 �
���i���/����(}���>A��i@Z��Xu��$�n�Ǡ��LNI#1�݌�ln?�	��yW��qC�y ��.^W8�G%N�|E]�{����+���A��m*����&�m���r��u#�۔j���
��$����s�x8`�!���j���Sk�&i�<م�K����#_P�T��p�[M�Ư�O�����Gs�2�������sCγK�O7�E���cN-���Ȫ���7R��G��΋��F�>�)P�2�'�C�p����_�;�E�����s7�p��#$���T�e~�!���)� �t�/S�d��b��q��>h-���Þ*r�Dq@/g�D�����.�Эů��^0�4�~\V�5�e�܊̳ж�㫙�o �ʥ�p�7�U�v���-�ix;�k�YS�]��y5�n���� �"�S�����&�=�j�`����).�~����R�Rls��6����M�eրٙ �4u=\I�a��v�]j(o_q"�̣ 9~�f/�g^ܥO~��&�6�OԚ���O��Go��ǳBi���mM��?���;xT�o8��jϨ�s�w��'���W^�����=ݲs�o���ոP�Ґ��w<.a�bC��0�o9�z��R%#��{b��*r��O.�Q�S�26ć3��^��"�NBW������hKdf���To	P�e3x8OF�L^I�!S"�R-X�Ll\���Gz�Z ����xbȯ?4++���\���|ҟ�!�d=h��j�[���G�a��-=�)���sT\y8�������0#�Lʦ��[��S��p�C:����B��J��e�M7�����M��9$8`�#tL�(�b��'��r~���ڏn����gv6;�w�ћ-��m����eMq�R H�c+~�дW8�����p��!��=+a|)�����È:�]�+`+����}�� ��9#���Q�|'���uS���9:�`lpQn�R	g�j���>����~&z0[%QyV���TO��!�f�TQ|E3S������u�;t=#y,o�	]�{��Y�f�-�Q���6c9#�Z��h�F2K�2�! ���D�`b�&�m��d��T�p�a(h��x>E]�8��J�l敬�y�R2�z;`�"g�z�MI�N������&S���v���o:)���-�ʉ��J�j)=V������]���|�r��C��]#�����K��1#%���nv{��:��4�z�?c{�>|8�^ܖL�/cI���1� �"c�~�|NQ��YMf�y�<�=!�X촿���A���kA����J��v #��o7�3�fC�Et߁������5���ݨ?�8t�K1Jk����yz%�0��VB�ղ��Qv�V
�����.(���U�T2'�����c�1�;����+L����G����T}���� �4-[;����+2Y�۾�~�k�_h�x�G�S� � �-��m�( �3�/���y0ucӂ��4��ꉶ�<hw.�f�W�3=�� ��ko!���O�l	�B��{��&�����a����lJ8�;��Iq!�B�̦��b�@���[]Nb���4��s�=��,7\6� �01�x[��j���9ËԇOhjܟ�{7Ʀ�����ڟ�_m��cg�v��\��S=��܄VjR��O	�W�����ж@�����آ�@�݁��S��Otybex��F�d���#Wo�C�WD��rC��̖��:�u���ۑ�u@��?{�B0qG 0Ħ۟��52�I������hMP�9����7�^�ӈȔP%r��B4v����>%�*��~h)�Bʥ���f� ��.Tr�;��ٷ|�}��V��]�a\K�&yΜY�h�xe�� ��6�Ｙ��7��_��yJ�d������r&�aP}&�ڠ0oBr0轈�}f�s�?���c^-"�]�IP��a\�Vά�8E�ʅ0���+h�n(�կ���]��w+�pT��O}���|�m���^5A,�М
1�}`��AHk\o�R�ޖҷ~\-�%F�<�弌���m��h�[�_��x��ϗ7���1��;)�z��3/�eQ!�Ċ���Cr�(Ws�����C�( ��3za�%.�{\iuSm(K�gCTj��Er7�7��I�7�;���+�Hq����f6'�ۻC�鮽Z�-�	w�hg* �'�&͋��{��!_DvuI9V`��7A�B�0���}��*�3?��ʎ���I�����d��@@h��&q���T;��`�P��`�1����m3 �T��%d��(�<�] ߙ ZEf�v�Qw`�^O�xq�� جpZ�I<mu
�R�8f7O,���@�sD؇��H��Y�ﾅ7�R����n��S2���F��X�j��J�|�=K|����]����A���xN���j��n��� ����a�m��^���7j.���|�U;;4��Y���������{͌lwO��WY���\<|�%�a+�\,mS�i6$�1JڂL鷶�X�ۻ�rTR>�Bw���6��U?g������O+縦�ߢa��F��#G7 ��
!���L������������T�#MAjկ�}z�0�t�ZM�1��ura�n�t�YGj�.M�t`�-�W�!�`}�@���L�2ˈV$���
�)��9tg&����2)?4�c��86d�1ʀ��s9A���pR��>����&�ğ�y�|P�U8ω຤dR���vU���1������o��ʳ�,�k��%�`9�� $ �/�t�-(�G�0�z9VԚ�-1��ɫ��3�4�3�����s���u���u-'M���8�~��/��`��8aj��=��Y
_)�W �â�%���-b��U���3��Y�)X�x��y�V�d�qS�:�җ_�ԩn�Cʏ��|L��)��o�@�+�@<��Ǫ[�'����=b&F��(z�2S}��E�4�k��<T�_�؁�<I�4��_n4��jIN�0H8Xx��K������9<Ro�CSF���"(_`�݁�]q`<���T�*Ҳ�m5�.�3LOְi�|!-�	t�d"/ޕS`ҿ���>*Yl^��+Kڮ��a�m0"����(ؒc2�S�8!w=^��C�I[�?
�Y�� �qy8^C�$��Q���
�T��ׅ/�|:'^��p���UNlr�v�[m�]��f�oF�/�_f'�h�L�V��I�mx��i���:nfu�W��ӣ�uX,�4�� ��k7p�fIԸʻ�	dl��y�Ὧ��86.���4V��