XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��۩߮[�#p���*_��y3'3���u-�݃����y�E�;�>��9��.1k��C���=�kDTo<W�qQ�BpD:���d�=��Ȅ S+N'�\M@�}�fڮw�uƌ1ocIg��[���c��g��˴�5�i���c���x�໗�E�es/zdX _�QX�������j|��J��[޻���c�ag�Mt�2�&wxc�B���cHT���e%��G��!��IV���H3,�|�/A�bh\	@<���?�)߲�cz���El�o95ӹT��o?��޹ A��5��K��ưu��V<"d�L	��IA����F���1��0K?�.�OcBI�[�M%�BJ0�L��G�o�l��}�"1?^=[���;��"���l{�Ty;p�e����[�y�'��+��Bxτc;N�����^5�MIFǆt�U0���*EVN`�Fm�B�!�)������f��L�4�i��Y�����X&��7ma���o�c�ekjY��8FW�
�sQ<�R\�֦:f�'_o���_�Q�@+�-�|�6h�<���2֞�} �M��	!�,��܁�}
3�{���Z���wz�ҵZ�ܵ"+�2]�w����nT�d�G�"����_��D����|��R����_�KГ�R���pz(Q�7")�1���P�i��@'�o�^Zl��$G���:W[R}�.h'�ٜ��y���nFۚ������8���/��d�n� S:�H�XlxVHYEB     400     1b03�+�P�T�s�6v���p|��q\'�q�$���o�U?�ka��d27x�������㑰 ����4�ݖ�.����3��'0�i�/��1窕�?��2-��q��/��č
�B���:Z�z�L�u㱙0,R�oF�.͐��6]�拾;�M����!�2�K�#n,�j��Zi��TM�]J� �<yS����� �i;$�X��3c� ��},��}��9] ��ݺZ�(��4�	�j@������5xS+�vt��5����U:{�H)��i<^ޫ�tGK�/�{bR�^UwB�_��/���i��F~��~�=^���^@xX���V,�oо����I�e�k�	�x��񲼞"�.������C����P�/^A�g�3h��?vS�MMu�d� �}J��?� �-�	����&0��6p�����,�a�XlxVHYEB     400     170�э��*U��v��H��b=Gb���q�	��"/ ���tR�O���	���c��>���{*�K>��Uc@�K̚,��F#�J�!�y4]�MSA�X5��z�j����p\��䲸�be2^�:�f5��KX��M�j�8r�썇X�񝩙�G=-��X�~:�-�z��o��7c�~8�YI��������%1M��ڙ��~�ߦ���Z�E�?'�.|���cy䆫���q>��jzq�-LB��
e� gڼ��i�]w���`���N���cM�le73���$��2�B��眔1��K�����k�����-E�q#�L}<	�Ox�'�p8�r��`�GO�Cf�s)z��@���M��
K���zH�n���IxEXlxVHYEB     17b      f049q\�3�2�� �K��_�\���J��Fkj|Y�k��鉴����/x�@�����y%U�"��:�iGw/��簮�l��CY��Y�%hBKӫ5����,��d�x�|5����F3�l��&��<��I�:pw>$X_�y�����������oQ����d|^��������|C"y���+���1�6\����j�Y%<�WY?;ԇh�_y�KI3q���*�����d�ӑn�