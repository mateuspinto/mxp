`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
BKPlJL/2w7nGNCGyFUePtgNM/Y32j6jJy7jfSzoKGCbb4JjOP+ZKupGk+lctZRCOwfr+ia/ppFAQ
foPaWR4yA2F4m/IulV8RGvYZpzL62yzXW3zHj5Lk4aWMfiQA32N6KQv/lm/EFNEa5V7NcXKSx3aj
98MWDdl4fTzvEbYoTGDWYG82JIZcpbZnZPW+PZ5AL9m8v9lZgeY6Tdi8VONk9FYv71Z/++4Syn8q
vSLIxn0qWWaZWbJDa/cMTc3VUiGYjg+s1xmM6JcOv98ILqmdyZW0iJk5hAbaxTqDeUnZWYUd0CH6
qF5KLbfB+0MMDiF0xJg3ia1ftBO1jsWLza3rjQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="Kr9fSbjuNkQiEpRd10FyUtolk+hpbQWjYjtW8aRkfx0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12208)
`protect data_block
9k5YXQ5gWJEMNqFww5wdjIkHAQrRIu3HLCwQmvDn8E+ckemC5GzRWTmQHtH/gx9azsQKPxfPlwP+
g8Ml399URC6p+qLXZC9Al1SezElu84Kz602l8wybslIXKXOwe4dYba+BL61a70GGSsaqHLTvJIC1
Pn0QbftazQSxCM/KabOQI0PkdDWnsmnq9lw9+3WjhppZwdZ6jdhO//7fgB7ut+Y+ATrlau/cSRNB
t37YxrJ5YGx/3JkVlDE1EB8z7w/4KLK6fCJw4tM2iIlAp4tEmKcPCjwOETyShq8tbyU7EEWWsXZN
aiaYQY/dxMoE3eDsYxN9nqaMkDG7cbwUf4zUKlufSUtLkDUb9SqHnaVm3PRol2p/Cd1Hs9e9I0K3
ZiGR0aVNeAl+nKHskb4Ynb4zH1G2GFJzy/NZOmctNdkuLD50lux93OZl90+m1MNhBhrKvPCM/Npj
GtqSHUR/zjWa9Z3cPMkbRUqknj7F4PXAFQmWyIQPpyMWsr5D2zHfp5HA6Wqef9RfRw1RbtW8P1Jj
oQwIcdQsZokIwKsDlnkmeTZcWFNDsTt00W01nl0wk7h4VklXfq5vAPz5jf4sFVgfiU4aGb7ce0fX
LR5oQjjLhjudkjqtl23+MFL1QbXgCRE84h7C4NdAnnHNNvqUhaYyECqbZDPL77dQnPoh2IIwhqea
4sK2SYV4++zs6OwcQghJevvV1FUBdA28EtCM7QwS2kPl3RMFaL0aJUk4LOhjB3jb9GlMTxriwZLG
i1O+cptR0TOFZusG/ACqfXSLAUJLhJjW6RmasVprR16dTzaNPQwULqPfHeCg1DGAdrzpyIRx+YPW
gkCkcCcpP33oC4T/iI2qNLnyMGXm/UDa+nl63HWWEEr8pjLV1KaAmHWF4qpPtkt53TQk+H6wadzk
IBSNp6sNNJYoLg/xnFL7b9ccuc3hsfncxRgk9svouDjiXMu2mbk3SeTSNipewbzvRdKIb3co7JIm
AZnLI3fiJSUVWt7PlZE9RO9COsiCC/YnYZ4acrdv4x3CFrq24ETSxvsypsL1SUViJVGaQrhveUlm
FqVPR5+Vx/5bYG5+ope9I2Wo00EsGD2fnKT3aA4OUwznnUyzMp9i1o/kO8PWioTQtorWoHqnyvjq
prerWtcSNu+6CA3wAFlDqeGVMzhLxpl/bG+RybnIS9WYlc8yflPCIkCqsmfPAmZZYvWVEn4E0JHx
i8z7Hz5yEDfRLTe8ivVyhuw41TY3MuNeuz7FMs5igLyJUyMURQiRC2lIgD9llTeRrj9lhFIPMhgA
5C/imtgd9xXGRA1ejCzftCXKSU5Z3UDaAE3zJZBGFKOH1Me9tJ6kjBWSHa+SQVgRYoAtfPvdo1N5
zSH3XDiTn7KojRUDLB93+sfSYLO789hkRLNGRFhQiurXojrN9XBLE/xPeY/BnTsvXTQM42Bh6KgV
ZwWQgI1hWpZy+P/jhQ3dipUInoR4izJdghR3bLIFfmxCcoh6GUFsmS9VQeJeOiZOIuNF80CK/wyC
dXbRv5IuwQIVpF1+TTu604vD44dsGGt+u2ceXFja6JVgL0W40BtXXq/R8M/XX+kdk0KU7bH/GylW
2erEjBaAuW93Zvm4a+7zv8X4Collp0ZgHTR/Atpv8SyZopP4nl2Gv1ei8j7Fyn0GwGDbok+ydxbV
RqnJgbb+QXgR27UYot8MihlxYor9lmM8hamSiv2ZbH5g0EjjWy8stvIGrpiZ0A1aTocTOfI7604x
HY2AJeD1VjR5M08WdxZN0QK7pdS+AVodKIwEl3RUpGIj0sG7yB7k+GYtb+dh0DhxTOrMxSsX+5Od
JO3rTItz8qpwdSNc6tUmdKIAEcDPKfKOKqsXZ/gRxVHN28BvM9kbvVLM1H8L3kC11l8oUmax2hKo
3mrZAwygdi4ngs8CjTxXEXgz4ZB1heVfdjTt8KpdQs1IksWn9q/X0i7OI7rMc7+/Sxpw1cmP3MgR
ED0nh8CASemZ+eVZiTmBdNNVOcp6bI5Ccat0E7AryNtsq8ZYChhQMu8kLQ7qsYiT8PnZt67fv9Sq
YYhRT3gmbx9yPSp3EN9lzeSTD+hXCPRXUEcjxQMYoGBGtPURVhosSoS4xjiAJdgjPKF+78fIy6aM
vS+VpMLdenKkoeH/tzZOnuF16DCe+/u8wLLgSPIgrwS3/soutlKBV66aXhA1HSnlnxeRNnNJlJdm
ORm2yLaymL+g7kNjhnFEIe6tQskKEz0qNtio6p3VvnAu1NF3a9idoag9prXkgILE6l3sBX0LVtoQ
2kXInbVDh/CpgARmm6VnvulUp0VP1KtmxwLJDqnV7tcC3pSfWmxL4QoHCnXoCMdkV7Cre0QQbIrC
+h3Fhdng5ZQ6M9/Qy1G/Ei/b9aXYQWbehzceDl0yXxnMQd9rhPPmFLLtp1R+XVZFn+zQS4rQBKUU
0/+SuD/2V9/Jq0yCdmk6lf4pXt+Bve44JCe0o/5PvcHlh646knKGkx/RU9jTYj5XPjUm2lYYf5wF
/29ubML8qWAuljDWThQ9CLFd4euYTmVL/2XzLU6By2+sfoTEgxmEzyWEyX4dpIswf9CxJTyECBrq
+FVfqGA/DtWx135RDtr3zTOfM8WCPYgdYq6towbkpZLyrRjPfQbKc5gHAbEp0TftBjWs3MntLeaW
OZAQIkXPW/T2ycLFHDOW4oWlnEGAxXAgc0Do3CyUCU6DPU7yDwqva/QVb8AWHbjTOnAQ2RXCvEeD
nV93Ux4pt2qs25d274ngCiPtIZpEln263W/jzB4t6BoPQFop/FDexBr09j4YsPFhDGWqaE8CnH5q
Rz1BWHpYxEL5ADdArfkFjBDKF775phgeOhEMKQI7jc4rKx7IGrXsWPBtTsoEF7clQi4D97Dz7ih4
JwDFsgK5mj8FbvUCvsVXZ+yK1PdWLLYOWYzXUPkAVZ0x2bSDQ5REdI6Rll0Hn7TF013j+tq7jIpT
9TAGF+7+LC2GFcKCMQOkgM3BfB89SkNysLhu9vC0KmUrgVtdMZSxo31eRUxFdkOY3zu5HB/ERkU4
oKh6G0xPCVg1/ZBNvvtPb4pw2viu0VISMA9WIcjehKc8NmZwytGGkP+5sgMMkjm1WBzYLWmUkJxz
jQtlWqFepy+XrgpfR5S74hmaheM+NpioVAHpmbRVjP5cRdW8Gd6R5Z6lJ3SkH7wv0M3g2eMuHLz7
476qXAIW0UM2oZxiGoMDDPcK/rV7Iz+S+Ei0RzAXzXe3qxXJ54m1ZcAZcqVbCT6vvhMZk6Zo7VSY
0fWjgoC0eVywTMIjBI1wZ/cqoKyCooXvKRVkjEpwTQYEb3cZYVXql0+Ge2UKbKGl8q68UfWPDgTZ
KbWYj/oFbiF6xra4D0yssWIL+l59isog0Pni8I9+SIwPxx35m53H4fj10ldH6EIlG8P/UFdhQAbc
1cAzAxZbikUce31S58LVE7ov0db7m03EuwHMbW69RKIv6ooXC+M6I6bhXtRQFD6HD4uyC65JmI3l
loUP3xx0tAJezOtSAJlaa+Kx6OCQOLh2Flz8L5ZuBzA7e8jDW1IyLkV2jat9apXfn6SRJJrVjRzE
JHN16sYFxsMKWDxe6KzbSbjUsAV2vKPR1NFWjLF0+B4j0C8jbbYzpXa2buCl9vR9mdDKtnoIl94o
Q9gbzTY2dN7bRu9e0131++hksC75oPW5TfdKJD2Nszx13wefYouHR1DviNtUhGvPsGMMgvwa4feu
Hneu+pggaXkxAVKEOEvtlcxx9zdJpmIrpKbP+sAWKoxcekHZUrzZ4ZwIoOvLWUApaun6l+r2DCVE
cKbNlwextjXSolfHXCaRbc8b5TNptNtO8cwo4o626KPzvFbdO6OQE/F1SKsZQL73E9ICIx/zhTkc
1UyexhH0AaSg4TIpbX0fxVXjbiTZ3lz9nxGspr9O3st13tpr/8ZENmGzHD6Om5nyA2nBib06dIUl
wfAcIHK3sLG1KYS1aM8uPx1443WnHnN+wclsWcg1ncyt5Yi9oRowiILY6qcEG8zT+Zi4RLGmWdCK
uStx1aXKjS8Un06wHEKUFf1xFtKB8U6Ho7YvOHqiS45hXmmaNhMjKPl6V9TfZFre54PbQI9jwM8O
C7jymbyYuXE9Ky0sjUDXas56apeIRJV8QxCEhobvKjbt9fJv0JHAT1k0emhLRn/8PJa9rvGVxH4P
8xJA47a1bDN+LSgZSddT9HQUVn+flgYoIaawZsxSt4L9AlXVbMoZ8umzp4mWKXInqRZDGO+a5sLA
MIH5MQ13Ot0tGpc5LplfczUaPuKUmPeHZZi0a0oGI72mMdlbReFUjxvFfkofswhQboOM5XaXK45J
jrfY++NxZcuvaIrfVG1wm/G0bwu6oeI0t5K8eoGI4o664Ogcqb1KGnwviIMq1cu/FFVuo35IFJY8
MijBUroiJ2UFXqP0B4MuyBJ0AnLOttd2R0U4bQolfXfjcQmtXi0sWvW3ZnPIbEGu18Ty9mj8h0uk
GnhsEg5tpzHbGifvZGorSlW93wyTPXrgg/0YqcuqSIXIPLaB+JUWuYz793FSeb6aY4NLubHZyaOk
bn+AzMsGxn9wnucN+syPlBnuCuyewixIqQEvcLGOqKvHo6oBCdf6ut3t7aX//R9Xai35I/AGF6nc
Qk036VhrGEet8rkHzWlVZgRXkgUDoWrWpvvxvsdryhlp3WMKmMrjFMdKG61IjOjeUBnh+yYrb84P
oXWirUsJxBYAdOOKB+RjKK9dR5BEF8ymBJarFgewicA3Qjsozehpf4mXgU7Ri1dPUhXJtIWhanGx
s4LqwHnaYSPE0GCpT5/L/crDCwGbOFgQeCPXyhUBmloRZVXBNcqHCCvgAqaFlTpuXSXBGbx6kz00
C8o/Xf8KqgQgmw1kN1F/cfwQzduW9UsQL8D2Ysu8AoNEEk3XoC3biS0Tf1yWLW5vuDcKqNafr/cb
PjQXKuWN804defDCtMi8ReD+3/25m7NXrOeF77H7NjOoGHxK33dU51Kqm0MRBiNUFYKCQ4whSXG4
QtGPyeZhSnkv135RIvL507GO3KJY2pPVnXT+8jpJRkkO06h/Q1wTRj6V9a8WK0ZEPk2/BIl/HtBh
P5aO2EgITPIznEEGssrRye+4y69urHvg01cCGfPafPSf34sEaHQAIp5PnsxUc8U5SdYD0Rs3WkZq
Rl3GZdFeAT10XzDxoceNbKvWH9Ve3kBI9Rh/+fleXMvGSwW7bHkPVgJ5sXnZp73EnJ4IrSEQqLQT
f3P7Wc9YlCLNIRCOwg6xuWcgrvenjh7WouN9bvcKTvI7QT9AtVbyydDsZ03ML0g608AGF+9gn+YG
cERKQ9wHTurQSYvqHCwbUoFqbFol+ADwIdcAFPazVrOrdM4oSql5tpyYAlhTKYW6m9906t81NPC9
k8YfNWeXSBF6lOX4rigJ2gsbh3ef8ePOQFL45oYHBQsLfV0UP4+z6YEfBW3dTv6cWcG35EAhx2uj
CT7jpf/YaZ1E9aBU9PaY1VY8MhQbRMJLEBnEma+9u38ldiDrDGOMyR5twxZOBbg5MpUnio7lTm+W
8iSvmhopSv2MknirmjECRgjWEU3+vob/1/xzBcYgtKfL5D74AmoFYnYP+QdvyAMIG0eqRt7/e45L
WwMa6+YpJ1WaYuvnXeQ/1vciQRe76jZLiijYSmGlJz968jgq8TuXH0jncJ7wi3IFiWv/yweLWvYa
BQRLF6Tk4QLyp+z9cutehI0pxWFVK5WF/C4VyEq+MFrZ3V0hXkzCHk4Z5fe/tRbiANw2pRHEu8XZ
BdmRnKUyPJUvEpNRCGpAzmly92uOEfJz0IqoqcSMl8qIoBax3Dfw3w1wleINucnBmj5sGjEOB3Ai
nWP1BZuE57PpynWqKShfMrO590teU54s/STvRGpDbEEQn7Ry09A/eWDdXq1HSsWhDac+qsYm/g8e
/VFXWXRaalkGw5mCNxD+/hNzDjgRqC2rt/vgl6I9rggWtv0oBclZBKbZwmRrVhqsGB4Ec8Lki3jW
fgwvEbH09mR5hpUaUC+yn7auXkwQ+xYAdQaQgurHEF17fJDUdd+Xzc0zl/nIuOtOX+e0rIE6UkXK
jlCCH7LWdFCa3hhSiA6dg9XEfzcMRfzDCW7a5kwErLfR4RXlSFFrA43ovQv1qoetZNIq9KFY3+yL
HDXFZmmWd3hnD90CQrSNu9ucesQh5I1GNkhn57Y3nfJ/LAC2aQENQTrUjd6mFLUgHvgm4BNepLOi
wH5oZcj9cDaxIcZDYzeGL0zeRCsR7h9jLOA5ydv6ux9wprVEo7Xkiy4IIoqTEfvF9gQbVMDu0hrI
zDjz9aPFamK+wkxvvRg9VvlKonV31vrzkAhGyoHwBYwNz1rxE1xqXE04HTO6hTtUTCKQDycRezRr
wXOgqru6hmImlG82N8A/C5bS44WDdCYWajzFtAiTVdLAx3bV61st/wdAB0h21Qgw02qNizoVJjtP
G3nNaGKA70NxddQdH9m5SNctKAhxzGUk1oj6hX89FcxxDjAInrchNTcwczWN5jnH+Vcth543NZX2
0wIYDVWwu6d6OQWp+ZZAPOuiywo1wmfFO2jfO5AXGBzGyNC0xG+rcoQHU0Zy0OTfIZCA25uvUxi5
Eix+uWI3gCRsgW7NCllnKYRcOtSUSk/t9tDI1u9MqG0h70JTf98AIDUTqIt978IKMR5dxbz5YaM/
Zz8kSazHBGbpeSm2/iA6caqF2bjoV3hAtcnWQENvuJJcRD2kH4DlApn4Mu+nj9TFWIRG75pwLh7L
5pYR5lvuns294aDJyfYlC92+iRdB67CyctGn/FSuj+Jw2zOALlSbCIaSjGlV0YVD2B4fw++YdGwp
6XHP+jsC5mxFf62E49BKeITykzN0IQ9agg/rEWmtKNzTwWvxdS8x1U9krP2pxHAmXW+7IM+itRho
VBnHduF/3uzf8GYZD0bH6gtFgGGxy7ixaeY3EqwF7PfTfDym7SkZ6PoecMBRlQR0F/QOn90o4Pnd
W7TB5I29wAEqHtm9FC5zRcx4eY7KIhjb6nWVwuKG2rt6AphEB4chiGiaTiXMLeofpKuGhN07vu+e
/FX3KSj/BIJoFzmbxzXNbl4bVTi8oiPhaumEhkSCGDMcDyJvGY7UvBskCO7de8Gksz1WEmzT2PBf
uOnMe7VNZIbqF2+3CgaOEcMZM/1a7p+FMek/di93ZDFMzlGmzOPGRNzaH2Beq5RE/W7utLaEvVML
iQnVxRT4cpRal7Z32xKQPIikTB8NCCdt7+kChvKQ8KSaicjGFaKogDGcwcfMcTk05d8DZ9q+Jp8E
3pHTF/CzBB7DyXvFYDVHwBLg11tdlGrdmMvjQM22Y4L2vnWDNmgFYVBt9aLZx24dYkntxUTF6wey
/MNcAdwK5YHlUi3hUGfIKDOemREwps1gjv9F6xPvjP6Uxh/tbAS36jkoKMuc6XBC6Afr5RAUkF1V
NdhZuOxRX5rWu51H3jDKS1TiNcouvBwiifyvIU+u7uMdWYlva6MTnHQMz+NJSb+zxcklo6j68bYl
CaD5HQLxcM6H+qD1ljchxBs3hn1/oUxQoyq5KIPHHwvdBpqJQl6XBNG9lXUwXJuJQy3be6FjGQX8
rPJrgET+wGQPv6gj84UaVzQVeiN8rikgHW14jhwQVQoz04wOFrj5ayrnYWuxxM7rDX6CwSrmZhPW
STJFDmBwu2xT08imEzos7xkU+nJx3mhul7yarN/Vi7cNpKiVD7Xsnp+GxbLpdtonF2/FDK6ZmveP
xgUvDdrAb9YeObOCt3SKyFa+4DFTVS1qLEUojYDUdFBLB3T4iqbk3lU01P4YM3HvczfPUOflu2Q8
j1C5ufK1jUd8ZdAgm4K+P0jAekMEN5+LdERYgtMwJaWnMu5JzwlBV1FBvQINLm48X2Ox00+VGLFN
KRArA0ylbw3A8YKCKw+lJi2T7j2FDfpbMFV7rmGLHh1b9/vEGlaRForxzfpGcEcjcQt98K0IcC4v
N4i7VqVLvlxcVJIrt2Dlsx0QVOW3f4pr0S3RaRjQsMXaR/f9VHaEbafRH2+PEu51TYUFvfcubOhA
EtD9wbHLUayBcLH0uojJEDePRHUjFhzxPQ0FzuteHV1vsleQ+aL0CiM4CvqKs4m8z3WGeQrHohNc
q1PaHrkKAr2Y0UI/xor9bS/BHoObdbWJzf7pegKUGV0797LEnwnMSsWUz2eykUl9WR9hWPIw1uNi
d2NKH21l3lsvxbSXQroDK2Kg1w4X0WuumEfZDyBWJfnCuU4PN2MZlLVFpsoGie7uuXuJ7Qmv4ipw
8cvotXFtiT749QMlLMjYl0YcoHdxO6CU6bKEXhp72ZNkuMmkt81wxBaAY2r2Z6iDWtyIHx5G0L1l
yb3N5mFbjvktrl7wiVOhWVV15xTphSXepd1lroIMaRsniJeDMY9xESFuEVk0D0g1WyzsIO6Dnq3f
sL2TGmtapypPcgOrIVjEocOqPFYrOvyhx98uLIP2SUMe3NCGqTZYkTAFpWMCP4EoTzt7WFYr9N9D
//qC+ooamgjrJObIEh2NEVb4jj0PWpJi7hIYul+pWeZpJfljdsQ0uyt6AhjxS/Ld3WlMa2O8BKtW
GJuTHCAnnY6rLaZugWKnrv7F4P8UtdoUW7qVbo/43vJWu9ZpTVQQM2dvmkXLH/XCsYVpgSignA+D
XtE3yjGEfrBPcJGzULTofXN3Gs2jeeQj/45CDT9ei26vb45PTM3jXJnlhbR5spos/ZN/PNQAdcqW
BWUcl/z6p3HTmDiyEVeJRcfPImOgVw43IB2gKUn68P0z2Hmk3eGOgVvSIA3qdNNb1gXsrorsJ8Re
aVMpZoGc9dxr5bug6mwBEiPuhPCWKIYPfKIx0By4zJeVXDmAh99LsVNan2uSyK6dAcMyo+rKKFFS
PmSvnv9zsW59o3bv66xd7mkKtkdb+Z1AlKNsmuENlG1dmgr5CLGwS7JHKbZctF7uxLBHJOTBVfz8
UpNKDtohR6hC4Lw9dG2RmMeUNfLq+5oa0jX9osyptgNclHAVpB5COCTLeiDJ5FaQnwcAsgnqE1Jc
PVRHQEyrwnO9V7xxMDzq0+QYXd9cAMcizjKfjQZyHi7uKu6X9vMhB1Bv0Hwrd+FFNwmRXR8r4lvf
EADnw705JDYGBZy8+11I897jgdr52V9XS0Y4DN/i4O8ilRIkRrg/RdRIYaBIzqnSvJ2OF651HMWi
SyW9C7bHZCBFhoCTiGy1yL2SPtpAC6eDFGCf5Nh3IaqFjr8607lryPEbrckkA2ZO26UAgVa47nsD
wGOwT785ca9sRn84pabLHLd+JdIei55JH3NP2LZ6fqhefuAmumXiJde4ZzlgR4KGypBVQXLr+Mkq
Rv6T4z7vXOK06/LBmJ/0u8+C2IB7TC32o/bOhKyxf+FK1w2jbHY0pSubRjoiuHr0n3m+hGWA9SEJ
4rRq+jBLAmrs6cWn6Lsj6B2cA+NiR8CPOzf93lYVTRKQl/r+iSq3/wUpeU9mc4GS5xCwnUfLUjdG
MKr/dwG6UoAx2tQh6jNk9muN3yv3MkWLNxVvTyGceTzFcwjRW7wr+h1MRukTPPyTR88f04z03Jml
EVuHcw7zhamphbLadaB8ispa/U/mprVIkm6zRWr5smN6SGX0VOwrhrJQAM1qXM1O6chnXCkWi+wJ
PWsifkzQDqa//OlqSBoim9mY/bO0yINAPU5Xe1zFpMv14SMyt3MQ7HzzKPwbiLAdXLmw8xZktSzk
LDIFqGGkDguXbjYQm9R+QtT7oFBNLDkNcGvOhOdXtRf6Qw16ZFufCLiTF92o/wvj0VycLqyUWB2I
mMNQ0ZYM/wEiY0VYNtHmmEuH+pJkrmygpkyxzN6xzFLyn7sDpp7pRtIZRE8g52FSSmL/WnCO5sIZ
/meoEhKrj92LENm5aLiaANmCoGNLUTGY8Br+QzkXlO1NIgeYfdChz2GeYKqaAnnU8H2DqdXRIgQb
KiMtg4C+GRxhrdtRuShbsCC8dKIwH0cWsKR6RXDimkHJIgPi6kkToGewzOBB+ZCu+Z4htrtMreGR
mEB/hY0+ZzZVD95NcW7YltZt27cBmw4VDLaqWs9u+PaFanqUS6iykZ4CKgf6jNrwjaBOzUS8gBcv
Xr04ZqeEYk3zC9gogtj2jmhvdgBdq1JXb2R2LzSdpQNkpLygOKQHEMBURm7Tu6mxMiuksNsV+tMD
BGfZXuT1JwZCXRJTGK5M/2oq+/Egt8rbqGV37IrSAzvFIb3nEmCLnAEAbVSgDvQR/+AoNanWb/fW
13cBkyfk1NCztU3ULOBUkpNsJRryvfZIROgigN9h33D2Qmnlcy2ikWalCi1w0Sr3mCynaBpTPZGk
ZESXmF2oSRyEh2F8mz+7q35XWw7sUGz8u7gFbam/li3r35AysRujp7teyDLOsVTfo8Nqn3DVYRIp
FhIGSZb8qK8JwRqyS2src6yWof3ZgP3SNADz0UXAasdh3L+IU9cw3PPQkc71LaRV15D22E5Yb2qO
rQBOHEdGHMp/TNoYlkNdPs8X8Cth3i4Oh07YlA4+nmPsIe1aFrGBamHE98ky9pYsfhvfSHWlxJGo
OyZFdjNxl6JMvuHMVBKjgw+Q6NgvKnuZnmKiggzWw2uiDLfoGesAMeqb0MBApeCKlxWpnLLm9iGQ
GFOJj3mdVugF9+FDpfNCwDxfGhmf2ip++NVLBtbVCSeXMzdh0ZFARTuojMv/8UjMRquVDHE7GOqF
UAzJlQ4YIN9Y/AJI3SLOcFPUGzktPrEXo8fuVsZ6owsTkfvM7pQWkJt7dL2giV96LEqlj+gAGoDE
y9Huf1XzwT/HMjzab4AcIscrMO9GSk2RYkm2KCD9D2pTj81xl+si2Behi/4+4WREMtXIAmm6KPgN
cStJqay/fIT6UWNgZu0nmeg/nXGpvcQKEcJ96GHwo2P7yt+T2jtutTfdQ8mTxXGO52/AqEtkxRxM
jAnn72J0b886Ja5LzWgewFxwR9lT05PXQbvPwQFkrRcHWt+nsUTBVEKd8kJ6m0BSrXuI25QH2OI4
uWu98mCfdxZv91qPNiTKrg7FNkHThHzSq++EFDUhrNgZGFRJ/bBFH7P1uPDCXfUumcSPDzZ7z7ZX
9T6wOimPXfp4wsbtKxLF3WZhRUoI0WTh9/zPwOG0VOTF7hy6+dmlLYVw5osF+FzFZltwbVbMDxKv
csmTbno+tAEMmC1yxlAYa+L/FxBmI/E608/3mtN2vxWZkSo4ldQTlyypRihfvgx2epWMkxGpcjBl
+WPoixqgRK/J+mrx28Bq7elYp2dVNLg/FT/acWjGHi/O2o5UK82xD0zSVeenYCcayyNG570xgYlB
/NnUWyk2ErwpT0q96ywtQa5sz9YlnjaGofJ0d7ppXztEoS/VP9JbnMs0SQ0JwGcHtTu1PnZG/VBE
UWCrna9BuVZ9a/YyPYOyBAhpjyiA1Ognz41GjSn0WlEa0ExVQcdc1aSObEuGjgfU4sIrAJmFLcER
6VqOFiOxIvVWTipeXvVaVdsTExo0wIehq71kXorn7uVje59wRolYX4a3O5zXTfZRLYyEM7AYaY50
KlzY9bC7JCEmnZ18FBwES1y71OBZkvR36mecXdQDxHTpUA+MuC6+XZtPwWc4fsX9mvn1ZCsb71iB
gCJPZDf4wAm6av/0Vr7yHv5qLGzKDKhvavw4tBb44Qr5GkodPHbQRT26wgRdJfFRzEQgEvP89BOB
sFk6+UH9u3IZLZd//BKy7Z9nYDk52oepf+WlX2DuzRPypePK7oERb1AiSje/5HfBrkGt9KxM2s5y
acaclNd2CVXi6UAi/gv7vFizMOWXrAYCdpiucZZFjZGQLFYaXc6Zs/sbQOOe19pZLSyq8JSkzCqk
j6t/uBXjfAYkDI0S6X0lZY8LyrHpOoqKZosOQ3Fxha/63JJq0CgLj7KYnLpQCxw0hoahNrcgCWL7
lqv0Hmhr2ZuBmv4vSAWtZdNNVlDyP8Emir1LRi36WAPKkdYdpSh613Xpz7p+AGhaY0w8I0Df59Lb
Azyhll+12/CaWuuU+2/ndcivJzIFtYBN+p8cz4Fv30TIqe3PXuyTLHpmEN8Lbsoqpa07HVmgSSeO
7VwA5H62BuXt9TmgX3Kyx7+E6Pohw6c+0oujbhsrT6zKYBOOxnlAxIPhXK4K20a+QvOIiXs4oy89
D+NROlmnhqmjEqW0tUwFVfsT0eu8Fbgf1ibfSOMsxVkpmBZzvQYoi+ngv0JipfkF4KZWiWGMm2Uo
oy3DMc2bYF+lwCYf9YKEho9I8AyOk0pDBXlIQ15Sj36foYH9YSovr2YYsg/FH7oTqo8/Sjli6icf
213lEWjlAzBEIROf39J0aQ5Ey1o1W2wXMYPNT+aj1ia1KE63OMiLX0vckLFE0AoR3epI1w/fxeWM
Tmn8lra7jBVmIb4hUl4xsUjoJCJvHHXOX+he4O8NSYq5s1I1G51TyBYmnfzHoN9Rx9EhBvxLX7ZU
1Jv1b6R9JZrZ4Ussfi/N3w1qiezXkaieFaiEV30FM42qv0tfy8SxuxNt4MOGzouUFw3kR2V2KQHH
ZKWsohgATR7Xuk+k3zkOoGd1ryB2JdeqwU6QkA13pIhHwSy4rVofolrjVkld/6MZq+riJhipZa6u
GxpvIE6jcMvFnZRNeN3kW0iF6A1l/1X4qfjMnJ9p5ODwoyW+elJfmizbvwANB3ytBhc4YpihUTCo
d8+qC7NskcD00RSITwssc9yyW5TWbIBjMfYAh8aV2GuXtG7EbCDY7C3+jv2VUN6W26iP7eblr2yK
C6UqZpcEc+DrXnd5rYym0L6zzgbm8Zb+G0N2Gwg5CIGBRLsDck9rsU3ASUG/ULxv1OH2CbQbmUOS
Wbeicv4kJAO7lsGAoFXZc3rCHMdzGJAxWGJ+5JHc9DfnIfp2PB/iVo0dSFHWmOgvVm8xFgBv2I/d
Z2IaOkHWQnlvu7/QMicAFulmMqb9oS8lq5Rz11C5Esu827hq9BWNSeTR6KBzbHnACu3M5ekIj3uL
CBZqa49n8+7brAQ+2nuQkYct8fv7ZA8kFRDVBI0LvWYp6a6mhXfdDVAg4yLARZMbNl5YjtA9Sbon
JZNWNIdm6jGQ/gSY1BLdUmTmCEapuvv4GPvEPlnZMmBcoUuCK8xGXA4KITty2pYvtW9D3pf42x6W
rN/OtKe/tsas35SkIBP8Zli1WYmF1L8yv9+pTd/yT+VsKMyymd+BqL7kjOuFEyQKTIyRkxvT4eQW
bpZT9CGWqIYQSbLigGOjEpzViIzHp2XjxvX2e2y58FjdyYOaZ4PSGJQoHGOHrkeV7wGkQSlCWCMs
ynAFUOnTgY/SUUIdS19ZC/H9SwL1rp8XarMjt7DNDsJZa1ZM8/Z2Jup7bEsUhcjWhxMZr5ugpcFB
s66eaiYJJ7HkxzlIdKaNs0BEbRn0jJtNtkfYQJhtcJxby4JNAIYAKk941BEpAhLIVA0dQh8RDA1Y
bSXn1fXlfkaZ/mYIfiSOvZAzKmxHL1GFbnna4oFUfN4Orhs/1GYof4qXeHL6fnbcS7qKzmba5Z9Z
tUimrMPuAYMKQxjebkf6b9EjXVP2HQtWezwVpw0EKp+UNE71d/ZypDbh1gNGm4PrHfghs3nQnjnK
Lm/LY5eyG6dALqPfDy50eJdCIqs0l9chx689pHxyKsrKuCLs0v9syGmMR+YC/ZZri4Q+251RRMS4
F92LNkvliEBvcLwI3lmPS8YAK9htpN1bb+mkmyg7QEWcFb7kcX1VuGKKezoQ6sKjjQyW4a09Vg7V
wokUNKR5SBr+taKokll6u74BEgGJdNWs0dpZZ5LS/mUBb6WagD46fVPNLKOEsvCMXZr1G9bJ5EGm
g8RYcfZOM5H9lLKWPkOUwf1UGfGEuxvaYxE95Njm95SyAA5fA827Troyji3qjGU1W0+alvmMT/vB
7dzsznZcwIPcGUQSk+qz4JpBBPZRT7ReDeIZb+Ua7NbLlVFPEhIDe2+KhvMRR4dwdBflmIwCJIcl
yQci1/m2bSRg4zq6kQLeQma7M/ZPNfYAW06eQIBX/OuqLtQZI4t0KzNgFJzLwYN29o0oD4AP5625
kXsW16QyPdpijZ0N36BDZpRVjEWGk6HDsB5eqe21LLYersUxv12f89ECTN0tZplPWtgk4WlnnQwL
EDBtMW0qy0FmkSZ9oYm8mQHgUiTlvKDqY8bWuC+lE6q9I5TE2TwYXGytHR8pDCctIxCFcimEJxET
oaT8jiaTLzo76qNBrSvT+5hKlue2xe/WtFH3ZY3pTqsIPzYQ6f64ArMyW0U1ff6MVedk+1y+0wJK
goIGBu/cUf0l2Axdk4FW9cr/COK51e8FtN6gOSWKCOmv/C0clfLdSM9ctxuI9K+0x/YZMAoUmrEh
TEgLW3RM61W85gRkWKLqJpGGkyzDnavjPBDXRfhmykwwY1q1zfmvj5LXgjGee+a9NVBuUsAjIj3H
3r6dR5WCUPGoSYuZgit7mfLvMkDJmwr26GHuSOiJKRzet1xrzkgvbA5fmz4tV9wnNR/y/tebH6XR
CsHLB43cmvrJHORsp/Uj1xn2FVUva+Dqds7zYIn9DrWWenvGUZpYgPFl13v9UHuPWCcCiaNI8+uw
BVRTGOUYL8c8ZNgXqPDjzSJb4yt63alwGpcx/O7979r0pJRabTB3YPg5NnotbBUqVisgkkeB2HW4
jCIB50kljA3KlC2dzxo0qLkFEc31T9b3s8vmWTYJIXbfzLrxVauANRotC+OuBil0bzdu+igZPpBe
CtbF1fFJrf0FcZQCwGbP9FjAHiqV+dMP2YjPNmkSl+5mkKDVeGWplHvLqiOKeZ2ShwIOLM2UlbAp
9ZjnarK+MrA7anjgiK/dbhUFgm1a1XLivhTopt5O7W/D7zMCg8+/a2ZJQSi1xnQSQyl6/yFwyFnr
IEpzdnhvjHl/XphvFWeWldiJOk1GNQXm4Lxs02vG/zaldsdAFuNDO9fQT9jcnA5Algzb4dMbzMOy
7QK0+Av/PNgIoyUvthCCfL9sDW9YaPRSERmOXK9+Mvpzn2WZP3CFFi3/4bPez1mtFkPRphR+1iz3
WXcBtL3jVDdAD2rK46lyVyWbVcAD1b4faElbGcXlIPt/JyyoNFogjzZ26lZuyC9BI2mW2+O38MNG
BHAnsg/DmPj+VMbuiuo13O81UsiUvnoMzc7oe1TxBHPMGCwvXoW1q+XhxipEe9Lv1JaBQb8NTOC7
BSJ2Fm2FICL2yE1ytdGnspnMQjfz0DELaOxSdvhGyjKuSKbzt36+bFeJmVr7Et3WnTT+m07+4vd0
z0F1/g1chUhW06DIr0h2dxsRom5KiS6xFcKhDe4P7nGzbZ0h1LoEiriUmpQDF7WRgkdSn8I8n/sI
1aqCnbKpAH7CCNM7OQAEaDbdaqIYrHRgQbA3iAh8Le6lhcUjS6VHdMC+MQ4zicsFcJaSTzg+CdHl
KkWFjX+h7V/+vJM/ilK2nU3vGA6BsYq7MVIwWID/rWGg44k5SYwxxhcV8+7Ihvv6Wzik9vwf06sc
DAHBUiSpMcPvv20M4hb8b4XNv2kRC/T8AYpmRHTPt1wjrzSa2m8x8LXam8e7Gpwhj7Nk4Ls9oubm
LDLGWYfb2VuHq+MikookDRU5y0EX0XXG3mWTEPuOwyi+5ZJUJOQkddCjo9LkR9j0A1I/St34FUYU
EiRa0QVNe+/9suMstlZSHx+wG0h96AdO9BWPH1im1Mb3/Cfvl+J0yDhC9cIxynmzbDqpKiNs26Cq
yldMoKiJEgGZP61cDTduwduly2GuwBxoJnnh8nRQLZrtwGtCiaJcGmBqoA1Wbodz96lCKTL1qi85
OztBcK5+x5WutKDe2TWyP95M6XmvwnfFbEegARukj+/EwjnOj/JDLx4IgNQ4anYDNF6Drv1SFtv+
VCXmCF0Pt2s+lAswx0UHzYSggApvU53Udp+8xD/EMM0ZbQiRzR5ETQtNM2ro/r0Lzy9w9ngSVybA
tzizVTEejPQBmWg7AagMeuY53cfvMf8+H6XR1CDjGY/zvdilIVBadnnmtgZYDoWpC5/KB5py/6Qa
SUlPXlOWB9UvuWV9LFwxR0T29AXD2ADYUIExYJ3OCx2oFQ1J40+G2IheEOh0nAAA704U+y0cZRrw
7jG7wRzpXWa0PRSeVSNgqULck5jsjBns22qU0/iTPklvA89iKNA1LL8NY9jVeiaX2KlLp82W3qdq
uytD8I8FxTcehD0d5DF3GEiCnRMDk4J0c8NKjvTAmeZPHW7HQv1gDyHSGud9am3QT1QqMF6uWlo0
LNiprSVNpdXB1Q==
`protect end_protected
