`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
TWRqA01ZNMBRZD409uaKlV+RoWhnlT/v24hxLHfzwZ4s0Jpr1DbQChHt5yJWu9D8ydSN4/Cb1fsz
E/ovO/kuJjcIWrAqMtcwtQyQiJuG8jlt8M9I80Gyn4yjplbIiejZsdbT5Pqur3a2Ao5rE4Or2axE
DgxC1c/64SsNftRBSQuNhBEVJ+7jdWsXggd1q7EoLD90WBefL87sB5sqcy+zg+dfHWPdCGPiiHIJ
eWGL6KTQqSxVfgJwx6p+5MgLwHaxb08mv7ztdEDl0H8SExvL8cLvhBgP2cJq0vatQXp/d4lSmDoI
PXgsEPqidTqA04cjuewWBxU3n0A7+sRnrpXb8g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="pMajvRV34ad9+1xGgFb9hVZU14lOshepgCNYYy88v/0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8896)
`protect data_block
TVKaswz8EhkG3AGsnjhZmidmM1cyY+wdeA5HRExcjY06MOvI3PSx7J1ylXIbN799ifVVVRCC8fnG
fVdVDODlpfxD464LFEtnKk9Tsy7ZOhChRYk8nGhwvsitykEBISbCg0BQnOHdOc2HM/ktFD/SGIUC
hwAWFiFFJqZrfJQNUV4S0VxHTW4YWs5UJW+tvMRgIvGgx/zGO9k2t7qV2gbftQrPXWMNjpw87oO+
wG9w2DqjosCoSZu3o6vAHLkxr9scSXUyGJYkXz74yzplsAlQSfE+aZTXpDWoT6e6p5LpyFXGbyOm
wGV9c2uKvqF0FHRqaCvSNORtWcjpewJWuRCxIMTOFXV+VAaWPE+rq/LvhbUPkAFKbUth1Z2XP3sz
GsWOGREOBCIzV2c70KBtxm2VW9MX47mixyrDFx7RbEpOQ1PVxoSQBog7CP4KvDBl5HdwImgL+GUb
pJXEHr71IWq2uSD+bDBAB4976hWPGTITlHbCunBJ1BrAppCWY+lK7PzJ++Ha5Zpx+1Tyt0v/tDyB
jKO+TaRtJkI4yCXld5IESN3woDawGaBL93eVF50yYoaPtyumqhxjcpv/PkoH4AVYZkFAc6/1lye/
DGHXx2VC0o57XjELBZVYEARCP5zskwaPqVkNHkOp+/+Hy+aXrTdKf92ElQZ5sxOkz5HyPpc5zPO3
33uNd6EgkfcUteKFQ38Wa0DejWY8pRi3+BgZG4bRbMefTnGhz1aIJMYzVnvIqDzq3HNPgDJqAR0x
ePHAKXW5yxv730zRaLRyeYvAUyEmAMS9nOH0CBCE2NTh3ENdw2wsdnBsq4FIu5B7DTbSJp7A6luf
Gx+IbUR8R5qok1zeWoyAh8yRnjTJU3pjESVGpRodZGILBCEWWqC/cPIl5PTuihRMkFgDVvWh8o/8
3aQnkab2Qt8kdWAt520vv3turS0F9lOg8sK0EusnN489JekJn078vFVHQdWbbhFJTFTfzJuKeWW1
dBqG+sn3JzXJD+E5agvE2M7KCwces93TNUB5yw9pH3Y96JAd8P1wwNpbX87TDSgocJNcD9EyEf1D
mR97otGHdiHmHBIDfcT4ScrE6BVj+TEItp2CcnCmraAe0beev8sjL2VQ1bKnogiyQmu4u/2wUWmL
gUxlEe7/9lti62oUKNHUfoIacqDwJIaCzii+bDwz3e/rjwt1dLDUAuQxwx0PKODjckMYYQ0BW77j
CfCkMa8TN0Ljx1tGmgBf8Iolngpok0ni89mKEE0SJQMas6Dz43WkIRfbIs4vecgIYHft8u6sLUYv
C1OpfXB8qRaCCynHpIvckX2Ze/tQmCqra8CPEf+aSQEinAFaPuZQy3QKbQLbpR3wABBwomfxdm4p
eGgLPkjLOKXB2pDzVBAo3gKYbFmcSyBoHKO3PXEXlxXU0Kg1Zf3+7X1bIv8+A9Ro5ElBLdnmDpbd
nkTAgEApfwmsjQyygxlH0L9AHO1jeocQIb2yN6OdvKm5SIBh6El0m2SxQqz3FNPY8cLOVHA3R9do
nxOp8U3GW/EYYANJFODSnsyJjuuiDSrBrb50i2NaKM64KKLzDOcAeNFDcAOZNQ9Rr09TKh4pxSi6
f3f5dXssKFl5/aWq0qhRnND6afNObmRM74wmQeydV46M+t9wOFPk5RwKJ0XEdgSSG8X3bSR4NE1f
CKLGi0Qc7bCeSKFqBYCjGUsnafBqCmlwi2Hle8zyR3G4pK7bH8KbHdapidaEonnsSAxICdmEtFjP
luz7mYDkhDDOC3xXHhZw7p6oDEI4+gs8Dux3zhIVXziDNYLSekVGDpVi2CEw9DMbS4QTKJXfjIRk
L96KHgiNzZJtVTfT+D8Kqr/tgOTKKEtUIuo1DHusBaBEI/9S0j9OtqLqbwcnJyUqZfdJbVXaLYaf
ROjgQhRMLUw0fg+xv+goKpSdjPZvp20K5RAtiKu1tYfwx/PZuBHS2HzRgSO91K1B6oOBDXzQ0sBz
n25WYkoIgs8okmPineNi2GXTmhAnh18quErEG1LP/rGlBNGDmMGQnStfbL4C/wML+RaRpJPMv7pw
MLtrdJsgHkSs2MzPoHwaWvtyDYqSKJLyCWPDJUgyl+ER/Mk6/JlI31iioNag4O+dlSSGepCKsyIM
PSWvDoE3PLgEnKG5M9SaZB6tfdWnPNpMlLMIEMEEgywFb0Lods1qdhu+VrSRLDWjnwNvhjhWlHLE
1vMIKf+my7+tohslau2l5wspx3i5JW9INhoLep28JW1EdrTleNmkuZ/ZCnkyhG3UPg4AcELlA0It
wA8kRd4IQtJrLOd6DU0jrEGitlIuqLk8o6M7Q6b5KobtujVzYro4oo9d1+CjQCaCRbXIj8u/mUcR
VaM9T+UnRDI/d2uQhXFm9KpyUcAwZSzVCdYAKorP6e0DZFXffuZtRNLCcouA8oMgS2TTtRf9Jytu
q8TLRzpAMwlk8pNA5YlAC7YDxVlz5eY3hiFFPfuddtBXDFE99oND1b8geDkx66JhkH/091eQK/Jw
ywOS26a4VXNJWOpCmVHwvFcz6H+oOe/yRge/03cMIVtdyVhGJ2xF+6IAJIEjrNDwNRTGBNXIK4c0
EFdiucNgTodZ3fkuoL3uU3aOqBAjMizPR+7RiaHlheaxEkTCLHYCWjFlpNg45Q4lNwMwcMxa7IRF
Vkj+tg2riSzp/tz1Z41znhYOoMoWjIbmti8Jbd8psJbDLnL8YT3zdIEkdYgrMDE7zrqtk4+AYcJZ
7YvmD1uV0SWI2tJV8Rs64YV+4QBcdytgIANk7/d6KH56O6GYg4h5JHJRBWsbc3romSd8hy4K7jKh
HxahM6qA98lMshsrzIaWJgbLq3JBVdMpDXPLvm5K5IA/0ymEn6J4exA6UtB3cr8voxF1P+xJKymA
9LzmT7x00DkNQb62ooVTYZAxVJHPvF3X1PPXH98mL2+2sfYbm4xuLfvMoqgVIsYbmQLFeoOr9wQY
fyxcw5/hqIsyeAAgSghXtQ/1k2Eh1iBKzkq7t33hEXvY3qzkhm4csPk2P+VHjvlZ0lWvw9BnV6Y5
ZQD6ozKO+kL6haIbqW2TnTTj4Vz1q8L9/z62TIaML6c7jaAt6ZPhRkPYwodPd7Q1pGbk5+xp/jim
z6aK8/ujJ5A+QZY+wLm2TMCdJV/uCghAUYLnbNgBAo/gGPJUX6Aik+OHQ77AtkOnTOmWqlI+FSYB
bpv8Osq6yW7xISgODOxsd8IsKPboiL1cWApOrixlUPRTF3KkTIbWlVvr/I/czwOsVT6oJXyqz9ck
UiIa4XP6KHAaa+BltR78wUTi201YX2dd7gE72MWMcGq+jNKmLxDGZIVzafekW/7aK6QcUgZNYDTB
X7NMz1Se5dzDstlbqGuxkzAOQkVcXs2thANM2wFJHkLBGAegKT2GNI5XdaoChQRnp1G146rcb5Nj
ur4V6XodeRacvZbP51WTRfx9qJh4fl+ph11tbAhZ1oM2u71v253D/mfYYlNDl+Z5Gv2ymUrnOT34
b7Tj7gcwwl1eBj/n/SM0TACuQ4i5gNT4X4khue3b7h3ydDOwPLA+3c4DKKpTHUn4Z+dNKTzXsWYs
V0bFvfv/yUmT+7TKec095FNA4bQa1mC/zOE6h6/2REamJkdmsMC/1F5mFf95rpsxV97PgZpZ2t9p
E1GVQon0M4apoAS72Oy1zM9AoGgEx5zNJdZ7299CGayBKMEF02xFZnvykJ7rn5L4ANJozrZQ54zo
vRvz7of5n8oihoTbsQC1RPLS+3tLKM6C+w6erh+SaIJs+tIOPpRqTPgQCD4cgDt3fqD/oLb0nmcl
HmPn0StCfau2Q5kMLvX4kD/v/hhtGYYkuJ4mtwBHI5ECqhRCvVjvIuEGqgRjaxa449cod6QGcmez
qXMON7HWMl358HBYybZCeXu6oJgaj48u8yGhgf0/6542LVOBDoBAkm78+qus+mkilG1eW/aE3PAS
bUey+hMJzyLo4krFu3l0XW4KmC1Mvv4zKNaTSxCCZgs0r0XprRmh4QDzHE/BQRKh9V/Gg+wsJVl/
PegmNutKsmXb0tKE8RhaTfoXx412gkUj44C/lT4ueM+mDcwpt176cYhbMfLkOhAiB5APt6c0Ss9j
bZLgBnKZcScDeGW7V4Aotfrc6bEDxaCK+jJX7gZ+d2vFMWpE3QFCDMuhxhTNBlr+jTN4/Mq1zgbU
mnFmq3SiUdyzQCRtrOKktaXEEnUZS9AMBZRBTAcdtTc24mFCNaIg3tAR/ILvgVzr7s9wCaCnN05b
WoISsmYJlBXN6j8xzMHORL92SN0kATmObSMVk831rh2e8EqiRwXRNSkEQS6A+f5gA0ASt7DSvLaK
OUK6xGmVbjUuMS/o/MG+9LVsmqLQaZMVnCK97v4GbLqMlKpRgJSkgbR3bfPt/WmJjkK6k+JK1yiA
xogbz6sJFS24GCMDPfVvXCRzeo+6lnFagaLrGDeEbCtC20UYo27LJjP0+1H/ELCi9oUdCSkBhJy0
0HZPdBA+lf3G8xFWum5tuMBI01dN8KbwmpWSnHwYkSrvuntRlmiiKTZ+nCV5Bbe/jSXvA1jfyrtz
TkcDuQQisA29qo+k4xcchi/YiIZbJ9Wv9OrVPAdE5w0jbT9yrrWYzzJ5LwswhUQ7Vma12l2ugY1N
uMXD+OHUsHSw5tTd2ZNgWapQESjQk0JdHE9XPpWvIZN+ZXIHV6yhi9xMWIaoOh49xZpvzJJboNUE
UNvxfuW31pIhOhyUinHS+W+1a05Fz5ABrfI9IiMnOptzIqz45JK1RHBNRRFHcxCBhYpBDa1sA5tm
+TSbaJMExqvEusBlRkvL5P34BIDXyl7R3yRn/QA62cOm+kcljt1Wf2OyqIQPviQBkjimj5tMCnGk
lj86rcHXLlPaxICof4Cpi3iOoE9SLoLT0Vrkndnv/wRfQjEWazTDYoVN6iKzH/QsYnTpjAEXsKiQ
3q4dy4lSxnsdeNB+pgdb4GIgO/WD8k5u80Np0fTbn6letqGKs4xJm9s89m38+kRli9MFlSz4nmeL
A2oc8rAoAf0oPtklD03v6yu2b557DzfaFJk/uQrZF10d/6RKOikEfz7pe9DGZBlPWMerugQBwSAG
vZnny6MO+uKygDAxcVILjJ4n+c5n0qUJkvJ2FaqWdghGG/RKFiAQFy1VaFOaBbsoSnsEP+arjyLc
OUA1E35GXvB0HV1AnHTQJX4H5w73u817e/SYU/dBd0sNcM5Vh0fZ7PmUMYdfzNl4wsr3a7MYQHGV
4dnxx1a6l6vDyThckKoVoEhU3dLnFvjiSFKkegcUmPEcaSMx5BZkVGtF2hrGLap1LKSPQTq7umKi
UAeuJCh0JzqyV/OZkycmE8ThYSCbzHJFo8AYyO2JpO2+yaLREcNZbNTWnKCJLUZUJ0thKIwmMwRj
taPz1dzvWJfhf/c5tUKbSeciM6Ti6Vj1wyiOwcwO82ICCtzh09DXo4Qnj1xt99CG00iu/7LRXcfy
NGWK6oPFZY8s4EVz8Gf1Vt3psO5LhQwke5+wgh6zCLn5aWcDkDzZmGWqQMNZrxIwxBHH9k4KbhCg
GOwObVSQBL8IxJZ96TFfDeQ7w9+iMXqJ/O6SoVS79sPBAtNl7CeDR8GX5kUMEIJuMLRzPNdm5+pG
aQau3kebQ3bgZ6MrGu2bfEcIvqzfH30ktwrY9lun50RkLX06Ce9K6hpjvsahpBqkn4qXXmaUZihZ
GYdPAnE7SooRYLBk7DNNC16/hz5R5QNNioMQXSmFEL7JSlX4nJMnBDf8wQJTqlT53qEVNSi6JJKG
PqV+yHBNGp4/Mf9QihDnk0797RX773T/N/04RfRg93c0eSdZ8ROKQKcNuDiR0IWFzE2BDbenopbV
GSK3g7XdNe7i5SDxqCRyL1IKa0VfZ32wU6WfOvDlhEp7btthLbXsG/QnicBK7oLjsoNW/jBgIxki
ypJmFuVCYAPSPN8npYMT3o9LQFIP8vwvgkXTmhfNSDnTxWeC0owSIzufo7E918XyDPJLGl3uCwL/
KVYLFvZOTILNW7fNl2GUb6oR+GKUiyW+hTmNiFUlLfzjSUhvC5JUDWd8TvktbawlWQSmlKe0bH0O
nENlOc9VzaxH6+35aEx3AYfWJZRCNITZflEKkNS8jKjKXn/BW2zNsEGVkl2mXN6SGmBSNY8FHJID
gEeJqmW+nwAyJRW93cJXWxcdx6U8pqTHRzGJhxlc0vnqCUOMB8JdO3C+mhdrdYYY8BQQAnd3EzkD
u7Kgoino3xxc6V0+p8D/jvAGhbtoHWXbc+hzIU/ir+14yY/yP1u97rx7i2c1gPP4AdPcgXep/XPc
Euza8hkelft4S26RgWWO89xsgPM17ya6lELp+usE4m35li2EKhHsgB9fP6BkZ0fzOIgYbDJLGsgk
qudKb+FJwjtR8s4CCh7LtrQ9HLegjPadw2mOvlkhGd1C6Pe8QJ3j9NRkmTKBgkhhRZj+4CR02C/t
hGGa/RsSdWBZwVMDBDeBVvfVnVn6dGGU5kOi5WQZx0chKwuGNSSDD7jww4T1nAuT1kWwT+wejPSF
Gi0lHYACM5CAzPhpKCHJS8LO6rTBhgAB8htCBufpNPpT3LULD3UV8X4n/pm8VLez/cbNUzNk/qs0
q9cPDlfAoWtQ+kgzo0/kXv+SsbRjyfhozwwyDQakOT7U2OdXXNmcRj1BUt89ubFKU9aMWBFDaggV
qod6JXcvE2nYisa+wejH8PXi4KbpYZe9j//qaRJHFAr8ILqjpr0FbR0yWNU3zkHIRN7JWBWftaCo
FpzQufW3mZcMiI74tesm+98kCMUWYUdTum0+t2lP6Mc4ULHIMhcULix9arQQpNqlH/pWiPxBdp22
370YU+UXbbbzcdGddivqDjh6FKaLkkWMYxHBpBEG0OW7wVOPDwVVbWGxnelTgWhUW0a7qa/SvoVn
KKxPZvZfne+trKLMfTM5l/8/yVPs7GchlnC3iEsjmlJV1sKPr03y7e6V0BiHiiOYpr8xy1yitCwE
9qtXhHi/iu5TLK3JnR84bWNQNRF9VgD1IgMnEMCSvk4jkz9usEuDmNdfbPIb2Y5COj/2e0YCa6tW
WQEWqLd3X2lHrksj+B9DFG48nXVRBC8c8yX2nT0OLm3UVahi+poFo+kkJmXXqnuky/R/BCleIYjz
EHD1pZ2KivQY91katKnxgy4vdiPD+hBX3QgsFkQol18lAv+fgKFP1SdSGDGGnQziAuGkdL1Xyjej
l705QqnqPCrk9Zhqusuk66zW9ca8YgeafZbCpDS2nGeJmHiaCMGLlqicGQsT12L+YzxiuFUcQjY7
hnCFExSGgr7MaANXfGDYnCyDCp5Emd35UnW/NfSffjXDtul4zD61jjEvfHP0BM7tnOtROl8uMvGV
ITqpLFR6qy4eXaonYWSXlmSl9HHeUlqArYhy4mzXBdBybfD6PU+FFj3ratwe4zlS3B/rwv6CNaLa
j59IMyhKCVsvZzZZWN6liZd7CBOWJWuv9uHsbY8EQvbTWDVLsLthpGf8Cwd2Q67qOVAWdRGyd6jA
qqBKK+OT7s2LubF31ku4z8cM9d7TSdA8Kfqh7zn6NnRXWokdvKLKpCLU6ByBnlm0JXMN65guEFRQ
XTguXk0lQD0RTUPiI8sBbv3Tddn/FJUZnKGwpr+QI/g4HaAy5luaTQzC1fJWH9rWjoK+efk6lCdR
+9Toi/N7Ltku1mc/alNKPfnSIWASU3U7n8FyXy/8cf9I+/VA/ePusr1mDsOn5Yl78MUGhFI8pY87
aGiNlVLuLNmigh7pjn9oEUPhtE4gxRNWEEB+B62F8R3fVAlm5xiVJIvS+D2BMw4sjvF8kW84X1L5
hIJwEDJ4Q6XxbcI6Wtw9ScQwfo0mQ9HjqQHqYK/asninz9eX1fKvrPA3IJJgfpVKTiAF+6uNt67Y
9ZChRgUhJJ0qgqq241k2PGx3i4jA5IqzYHQnxhGwpxrhrKP65Ixs6jQ4s2SWnCXz/46ai2wzQHEJ
v270YtOOBgyneaprtEknJhRKTm/cwiKyyCmCjmLmK9lgGdg+xZsHe1ejSdc7QObsOwqZ7PcU8BCj
J8YAaldjHwCFMpVQbw2hdXn4ZoAjyvXJ990Q1yCkMGPqbHiwTh6jnNIMHAIU3ooKUQB7hhy1+Ipv
k+ipc65/sEwIbPkZrQq4a0EympNX/eH/U3l0zlGGQcc9I6d3HVngAtQlyVseLgghru0iJE1lEgp8
up55EnomvB1GF8RKQvy2b85L9b09/lVtjAgGEuNnpNpfCpmLGUQY/S8zEktDZcuG1lNwNYW3Year
pfDKOdO+aIJg/6caTxwJck8UxTKrU/IfmfhBjZ5CjK8C5lrpfoqQ7VDsemIh5AM3824sNemtORk2
pKKrL16CE6Mo40XZlp0NEUC4ZLUZg+iPjUCDRIqOtUD/fko1YCXWAYUW31iVN9HxtwsiyHVz6zHD
qhQV4AUECI6Wwg5RenfV/kLn+r0ICgGHae04u/M/fVkVYqR2DcKA9klzVTt4xcTfzFfa2aOu00gl
kTEm6FPC1EcMRCVTzybqVj+OSfQPcMdosDUdQQ8pROkrTasuf1O7Gp5mE7PmMRudtRBMINtgjQqO
Gz0pI4q3BIzlof9ZiFFBNeEyiYl94AxEtHXdcZz+JtAl53n4aaMwcTzFG7mIFjQdSB0DPl2AnONJ
F8NAdNyU2i3THPVovUZ1fXZU4i7L3UJGF72DVu0++9/DKuG7x/J1EJ/jNyjPjAYo7YejFuw3UHAu
JCGo26z+zXE7gx5MHV7N2QkPsehogEewka7iU5L8CtnuoupyDz8/O1KhrRvE8WheyiYhg+jyKxAI
IIWVgiWUv3scHI8AB/ubVZM50qCGE4ymZUy+9mjmtc+1H1nbE/czYCPX4l9q6fQdH0GMHjHiabOW
mdCLviKkYJ0OSGZ0YbHJ7StG0gD/DBDeMyybOBddN98iJfi5WyHtIY6qywiSErayJTXg7Ac+Tdn1
pYv4xLs/NpIUJuywC7C641pnkn+P6HrGDb4bMcIlJ9A5BIvdvSsdJhJ9K+voN8r+AmhI7ESipjay
FzB7XIll0muOO1eT5Qt+3llFgCmHpDLbE3pQ7xQyCNyREE6Kzn9EqZDIQrcxFjhXiP/83r9I9Pqp
LsCuoiAuV4tjMJB83m7XrhhQR/ofSZQZnd960TEa2KTikSZKfxBluIw0jDYRR8ENqM4fI/gSNGf2
8aRb/a0AXbtOeutJ7ZP5Qa+x+6j7C6vtj3RmsH8mLGeHanF5WkVoZo26IWEDfAv6v8pzIjI9suQ2
xb4CtyOpVWgw5RluQbEFnbzNdv02zlnFagkIR3WGFlFVM/7NY20KsWySIEIkejO3Nke8UgxhICR+
0DGrxEoRHmm4Z+QOMDN7wevsFO2QMuyEfIw3WH6IMT3+GXesQN3wSnuoxYMZflCThtnVwSEY2ls1
n7ghgaQrwtxXEPvGUl+i2etdO3dYq4Na02lsjSmE5SymwBTc/8uLO5GSmNkgYvBm7vEp8lGBsiOn
RYFRLxUqylFF8okteGwaP6RvrSvLhETf5F9dbhSkcCIO2oYm9pOQbghZXvC3JbeEomTpqhu0dtbL
9rU47q0RdtbPwWvFTTRRKDwatc+oghYUwShxpfhI1vUTZDK4Z90uWzsX/2jeGtj3bhukUEFOGmKC
kFiVAEwzk7gkPQ5iI9GAMUpyRBOJllLXPyUebO3aqsNCAytfdefKka1XeAVD9urVDRKYzCf+K48J
IDV4N/uMDvNGpSBwDeVSbERgXIquhwoSmBK83EHa2BUgILeyehyLL7trx2kw3Xjlc+jppOLpnxxH
nl8xF9yZfGQN/TozNBmfan5P9NEOc1q8eMYMXjUZiUsonoUaHmq5Cja2axy3WJIVAvhJiIa5Noa7
LJxNef1lTQodDt2S1PKASUi6DNe+goAc/0OF3/Y1KJudKB4eAF/R9hAVwPX9AzcAw33Kh0cMsWa7
klJeWrrbV4+uffmuB6sS2ahCLEA/u6ERYibh2H4wAoUEjOWr5tSIZ37XRvbEdE7uuBj+uTO1fFCB
xTx05Al43+S0iy3yux+g2P/7Hzi5Ruy9GnIdNIC6Gyv3oIwTOMpdSGw8ShprTY+AiP7F54j96x9T
NWjj9w/lT4b0ZR5kUrWwXL8l+XqiyAHvB7RkIgllemC1uZO7DRcUt7aUMtU4IJBHgbIO0/XMudv0
4e3T/uJGUtTCJLrxIg8lu6cWbP73npdqpQkFkXERDqs/6xDoEYOppwL2u+biFDGTvhk60IFd5+UO
o/MJq3XVTIdYIxQIrIqSKtTh0CR3elmOQHpBFoD3GHvf6PkoPJribAnPJ9mQrYPfnHiOR+CapFVp
cCToukIwCouF87INdHuf2bIA4H0ZV5Gh8T3eGtyWj0DdDFfXtJVSblGh1j6loOrX4aBFEhFzQgs3
A+f0u+6YP/+gCax1yZ3tAr8jauWUvj4NSvPTBcurWDBvMfisiZxFTjcQFoRzhP2WBjRcATGmYCaP
iROHdodQpBv51qrmD6UD9elfBoaN2eoOz97HUYRKoeMWIDy1rUn7/4k4schfWvMIuyZ1HT70qOlm
Jj7gLt66Wo0AcnrwR//AfQWu8TM+u2HBbxTmvO2kD9OMIwx3LduGAEdOewCGcpmTgpq5WiW2IM4s
5DUx+pobm+vUXWMa8Bl/JuW0RbbZuvBE09t+bCz77R8KgWU1BDAkZLKNm50KhvX0ziz9PAIE4Mcm
ffBhE7MwQkx56Ge7D4bippI6kXHv2JNFlDqYFKrplihNmANG9MjqDTUmVsGEiZhsd5clD1IOxF++
708jh1k0UIIESrqImaumED1EcZdP4UdMDa5zybR+mMOu+QA4AKyNH7huBY2ueJ9K0CtoRA0cMCgG
uEwmRbEMGw1jNi/AGTuHlNSMkJfKqlSZ5Ea0yuspNUMGTuaQ1VblneZuEqkWagz35fk3FYHLJQ2I
4mBVHOAAREngolUnitMvCua0+38rkzBATbgg+2wpaBSg6RR0un1un33w8v2KlUu4hWI8Fp+RZ/Xr
Jll6mcirF/o8fQO9IJBPhzw7APIFRSbuMya/ZZmZWuOWl+HD0OYM/6HIle2FaBxp8bXH0XscRffE
hFFmGDMCuSx3i4iItk5a36g+oL4bvChkO401NU0i/uBM9keJvqjk9Pn7gFv+72VK77rcS7cO0Rse
Pjd+hcWKfGCipdn9fdnnu2E+/q0LdxBgo/jP4ST1r2tSIggvrEQhVfqF6QzJfbHLglr4mEMaaUQE
CkuxtsKU1MOmHpvrRJ04JX5bIn7QoONb9097rfAo+IKyF/EzxFgVWWyJLgNuE/VgFMoXACZwSKKV
3skVVJBuvN6XG/ki3ib0If/1pYR92WLkoFMfymh9YVPC+/GuFdsSPUR3dzYGGfHsdN1zccAGvDgG
xe6Y2uk9XaDmkQyg7HYz69OfuqKMdOfTTqLmGf2pC5aVNYVZbIsO6DVtp0GKGzWraEYX0u3oqkVX
CXbhd76sw6M4dMIwepnu21QoK+KdIkLKGKE3vZCelut1ugmLKv8foHtuono5benl2aP/21gD9hZx
dkKkaimgAbKsB13ifXr+E9TkzfhxwfMseJvtOSmN9zRupVfcDFsiNbqMYrGwOYoZB+IxQ+U0Ke7G
HqbLQzpohyizjTshDhQRAwiakEDMQQ0dfqcrOQd5Ikkj266sWP9IKX8tkCjnDePePj+6BE9KI0Ms
A7YEAfeVrBS4Mbv3Jc3EduvL57/CpzJiZ4981OiBzSxSg8bkjSjy24CXsNoPWd8KDFiBdMPVcn6C
64AwgeiaiKa66qr9/enThoZBq3cHmNcjO/UY3J8jyiKgK5MbpX/Ucd0ex2EytCKTKGkbjQ8vUNID
RPWYqw==
`protect end_protected
