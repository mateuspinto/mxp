`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
sEvdomJd+1Vk3egbHlDWf9r/TE/qi1dB6MtuTXHTtHOEl5Z/HEmn7qrirSvPsUHoxzHxlg5Gjl1f
nSd38izJT26wvsGQAGno6YsDQglwi4FTZvX/x3FwCxUlt63PR/fa9J24RCgH3G+VExyBICB89vfv
2P6Le6oKpt+eifBbaAZMc/w5/UbYCOr9yClv/DLjphKim72PjTQcsjHuffyzfCws5Xk6X1C2SPbq
40loOL8nhaqpp6rb6iefOFNVFvNjxoGWtUG68R/2bid6xh+0WewUe9nTia+sOFjL3EeHAGCLzDYk
ABIZI/kD93e0gULOK8BsDIPXONSE9KxvHhFI6w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="c5tlVD+ak93C33WO2F4gTUK+VQSH6rS+zvIM1eudhG8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4400)
`protect data_block
o2yG2QCz5iv435lbwJ1Wr/fqG1wFXtML6BwpvDTCpR48pfeFlebA9M9iZVGOfYad8Ex5pEBfO+B0
YftstQIM45gu1IW4QlqVvVqUlWY038qMFGEdpEdEkzHF7TCKRumZmAv0EImAQHh5XX+lcGRSECR+
z7HXtAy75WwVqSOJQBMfrAHwiVR/vt0TqNav99WC39r5L8ZkZGs8vC+kheSfa4o1JbQigpamgB+E
3afchxVVWIrpUSDVWUVGMrnTshJ6sZvJs4ojDxh3tPSCvkih096GlvcLWyPerWWsCTfqX/AhEGDP
mIGXWFJbTOFGoGJfFnqKGA6XRO2qQ4MKCtNgHwOCsREXpIExBLJmgffbTvXbkZI2yn74vo0EncgI
IMm1J1p5limMcFutxYDGdtlR3EeWI27cWNmc9jISjgF25+PEezO8aiadb2SRgTcAF/gE6qUjDuZd
WwxjIjuXqhbnCQ6ztP/iRSL3NswQtAXZP8lPwrIGnRqYSO2oIZ+FTfe2FHXcbre99VMxtOy1Ef/1
Rik2IW5MVLYiWq1vBwrF4SNQ18NyiIk1lV97gxNpT5xhdeW3Qub1oRxT77kSlw4s76KiX3K85mIQ
RthajaX1brqJhK9vQEO0yxcp3zPibSqxSuMWjsPgkI5yo+bH9eisY00PiZGL14DReQthzugakA+6
v+SDlZsARPCPcIK1y2mFGfShtlOXkEu0ajpNvB7dYizGG2bgzIAmlBOrUTM/uqJ+ojPBMCUR1zaA
6GUmQImIaElvAWk/zJphkrfwSxAQ/RW7/C3GqchQSdI1BJt2K/nNE7BmNaNLQWZ5cjJAuSqXBR8u
amvjFyo8qe9enytGZ2yKkkT9k95yNtzLQREqAcmBV4yjmJ6x9kKJay183jfg+QhVLvzRRxKqQmNl
o2zCWfEIPv3oAtWwpztd+TQUNxUePc+dJsRLSBcNwNpu40UZ7ngAtOumulHbvdEvFmlyT0fAHWdd
p1mplnMvkSnITmM3/FQwM2c8TG//T1Kgt61gTPg3Hs88SCazaZ9Ko6hMABU8q5x+N0jIEwYbwgES
wULEbkIPvMh8FSkZg/zDkS9MrXX6d9k8OmAnR6UU4tLgVdmRPgWF2bTLk4ywCqvbSuELz6ftv0qf
CB3Xgdd2vVcR1HKYgC6L124aj37xRvzldWOMh71qa+XeEg+8HtCu/8NJ3zpAd9v7WynfbuSIV5OT
XbSASnziJoSq7ZKEeTmGT65yZNWz4AAgPnIWBiIG8GXzFm1ih1CJ8k5tq8AU3fdMIJ9o/Ie9p5kD
4+Te0qSZ7smlNIHhkiUkXp4G1bY2WnKZHWXpyr+1dPEKma0Huor/3gg6+inat4wmt0NIaPbrJf8B
bWE7jMj+Qabi0Hg2x/ISDBxSbn6u7hR6xtZycIT9oKG9fNjgzy64Xc2VOdEUvcbu7EDI0xHo2KqA
JgUQElN7VejDD87jbjlv4wMOwlD63uQQPpIYn7hEBfqELS5+xmZjwjKorCQDw1LPGrZT3oiAb9OU
zk4/uzfaiKanwU8eWNT4j42x1hp8COlj3c/ZCCacvgLZOQKb3FgcJXZNa753rbyS4ueHmBtNtRai
vWSWy2W3jUaVjzsnxQ8ldyHQPbG+RAsVHHCh4/tdByZfD9deKPK6xHfOqakE4UE8twxEu8v0Om+Z
WnA2xF4j+RhqFPdaVCm+x7p9V3OwGHLJ39fbhoxzbm2HuYvd9qwGCvdd9RRAB0Kv9qvuuywbfo7c
M1CFDPiTS6ig7ESyD6dGm9c4ZHaexInF/qe/XZAXgaE7ZAHPh0ds5CLvSusdd+Aiu3nIRCXpAV0f
jee/CsosV0QzmQDHvCZGUZbpiyrls/GkXKlAbLAJkeht1uM/V1QFwexc9odaKBgb5CkseYZLbZa3
x+rY7IvczUpJCkl40K7XRQNQJs3WrOZftql3ZnNuMmxhaKdl5TLjRflAClus9wezuZGKf4Gmhk6f
RbMmw5IMKIqysrRmahY6irSPA1DnXcVD2dQw1HhTHu8w+FoQ1gX/DXj3YiGHE4dc43LQz9wXRxZB
+9e9NC/qaJjdWWA0pkM4iyrODo0Xfj/No5ubwpnLq7HlfVQpu6DrmpaqOYWfzJqZyZdNcazLWvFi
c2I+WwiN1l14jhaHXuQj7iGQo+X8l6N8eq6CZZvSb1cJff33Ev6lmvUt58OvT1tByo/gqGy+GNk9
if7E7JHln8Fs+wZtu5SZogkAqK1AE6UqkYihr+gJQq25yv4FJwG13jdtaBqeVnML5PnYCRLOGkEE
//5BYWnwpLfRP2dWn2NSpgMrhAlSqFpD6ueXlQw84fbLSRBkAB63omq8yJK4A6r6tQ4F07h2do+i
TAWOGLNqEcaLAZ8s5rYgfz/09GNz74YY++rvnNjwSwBQL9PlM44EBOBEsTnjD1sIxCawFKWHa6mu
U9hI3oLtRXWQGPBuXGkuXZ/xhzOnhkp3Dttf6k+jBo5VExcEFP5S9Sb4h5YnwduglVpka1bgairN
5fUlFmgJEQbP94W78QMj4cOYmbanLul+8KNH6XqONYmjwxbF7o6IVU5NM9LindGbYaFZSkZXsNog
FYDVPyFI9tpHUDBhTE229N9m5O//Fy1zUxj62EJSBJmpWh/WaG9Awbc8Su/lEDm2QWDbFcD87AO4
7VY0Kkd5HRdcBfmqsEUu9O1GoO4832Er82eAsLm0iab0FwAKDPU40x5x4QJGOFmfc7o43DijixO4
RHxXEwAl9X/PS5xN37tXJOrOTtn2eQaBpB4bwVye9A21BcMRsS6ebhFCGhi65uojlP9kLeVAL8Vi
zE+3Aacfa/HPcX8UA2q9XPx+C8tlhVIBmpe3MaToFeW1EGUzLca/OOs8yVVzl9qYDTlcx0gcdxma
w1pSHOsKl0+DvEcuk69oDfXL7Ox4kPrh+Gavh+XLeXOFUqpNYw4BtOmGJfZtonmemDu9YgHZC1Ik
8DV+dj5H128B3LVg1ikqr0tRTqQI3g168toQCcHtCbEMzU8T+QrVTLQGCvAc4StQHFFfQ/YNm5jD
IpVQo42e4qv831m3XqrohyPfvpmEiS3TBotuQLfRXkq/TSDPkIjalc45zWX8H38/2DHdPu7skbQQ
rkAVRZv5XUkfc/tTIUJkyr+EYBxrU/uWof5JnHJ0aZ3an0T94uQK+xOMWDhI1WZf2cYceJe1vZaG
rp2YcJDyBwXPLuGuhgtLPHdPzz7brM2sd6EnuBJ6TovlvUp79KRliRYruxl2ex9eNe2zoGwPucO4
OMLt/SB7Wj1+krK8a82c9KMqYCNFlWSIecXThoEJckCieNBQzLgdptR36euhC9KOs0t/yXRAR+h6
6QdxYHLkIrSzyPhCeQuxyN/qsNIYVFV9Dblmb9yHTy0t2COWdynjQmNrli5bn0A69i5L6fYaeESJ
KlSZa7M74V/jr7ertYxNbC3R5xtvSnqeLOMtMybimsIhCHsLt0KjS8cAtCtv7212abetctVK//Dy
Uhixf3JIuIIP+jHxornuAbl6OYYEs3pFxkYUz91tr0Afj3ubHTM9R5KlO8A9of7m2XjpbpL+tt76
oT6E4Dgp/43yogUdz6ENUZ1aTBxPJMHfvwgenuUu/TcMx27QCJK8kABBpGTlNN9cH4AI8sRpQTN/
G26TD6+mJypyHj4zNZ0xi/JDU82sU4xV8Vv0aB3v5K6zn7oXnApfNbykGey3kttDC2kAhQaTJg86
p78sudHCjSpcfClVr5MQPNbfkGUOy3E+XYKkOPXfxigBml6Tyf9qqawTYZesq/NAATW063n3diFL
znRSLZ7ZAcHZjS2FQgpmG0LwiJJFs2GY0oKlSA3O3cP+60CdOSE67O0/mp3RcHblfkjQZZFsBT/e
NNau+NqqwRdqLYWWuPjxpoqucfLxdWsWi4SxqF02k7NkYpPjmYX3SODHeZ+SV4Cj4dxr+suMPzR3
z6E82ZWPXbXNS1nBA/QZgJYXFDzajsqDjKzMXcKEVuLVU57mnZCI6ykEzkD6q/ONt0C+8HANmjTs
fGRI6xVrElKVI9saRZCte+L1sn0iL/eKobi3FzXLai0L1mmo6vdGhGYXS8pJJuqb5jqW+uHKBckr
2xCnErNxmyafRgbe7ByrVfbwpBiGY43ndKDI50N+uc70RVHxxQaZBOtxNW4RAFYG5gFPxXpAHVkn
HHmnKn79vY/HB5e/BwZkN14DjhAWzFHJexJiVXi9QlmjM/EHIKQpN9UnTPInTX3QgrEiZyeh5TNF
9GDGlG5XZhhIK0xvJGgcFKG/hzSSqILz1HY0mS+uz9h0HrUx/Nq6utRjySVS4XKjOf/UTi1j227b
/qlXgHnXdTQnBmS0XDSUeVc0vGvbDsuxxT3rtF7qt13GsZJNZrJnW6JIzk125oshACTS1ufJeGye
nwtNdUJlmFCMbCpqNt7uF7SUlt/zHWhVjgIT6SiE/+91uSdBcLURb2Aaazo18Bu+BNLhlM3N+2Lt
+e7LBTJ3olaGoqLVLfh/O5gdT1j0Rb1a/FJa88K1/QgoUTEIb4LLxvEWT06WTaR94nwIJEy3iZ2T
85Us2Hj3BIm1s1HoVVvREtY6c7NjrR3GmDhu1S/p676TJYTH9cPpPMHYvDruzKzl5MOfC6mVqS+R
K3mFlcvoMz3tzFfncM7qIuFAC2yWZlkeSUxnpicSjb1r6ixw28i10p2ZTIK+gJrNumPrg5vMnee+
JtIGcz9zVlvbkMvReo6arXNVROhCKDiQLPVpFOJJXGJOVSAksBq0j5U2Tn+HWMV0vl3LIbejuqrM
9CRt8Gnhj7RBWwyqa3ADBZtcqD03sivFE2O/TIAbXKgp6gJDy7qhUHJYcVlCs34SmE+Uo2BNl2Gy
J9JQIj5HD72z04OBs38hxATqvM9Ej3OSBpg8o/10OyBN9+huXwp8ePqLN2iJj1YyGzHbQxV20sHk
yfuPoao4VjIcpOI369VrnbPiyJhAyEOM/6R8ufyPX2v4R+0+LYJvqzYwXEaeVi48oIcu0ZVPVDNi
G0k4Dh65vQWsIzCuYqKfNw3OBtmI8ICecAWEbKX5OOFTz1D+xFrB/PBIjOyj15x9CRRPrJVjGKIM
yMmrgeYwqf0baCBp8sWuFwRQg2opSkX0NUJ45ed6iQvUcNnUlqIyG0FhTwfZVVVdGzfWa3W1YmIr
u1n7Cy6NTC7B3fyikHQRr7NcLZeUojdbwl6CQ9AqK8GW9CQp+toDDDIhCsphVl+wP9BigIjSEZqK
VvjPLiucVYlCKszsuqW+LSufUWeTXXE3v54iGaW/7IzWQNQUevkVV4w8mJxP768DHNjXs6L7wBj4
MqDJDq1v+IsLl4Td6QLeCrJ3/m+jr1+CAf6BnRsTjuNCfk58mRHG48XjTXaX0w9/P0jODEbKdjbd
Hjr4DV8mswGlEebl1QgIla6kQv9fBMxF8V28+ywKlmFoaH21LziB2Y/vMEUXyHZVDEdce4LpcyqV
VauULa/hcHd8ggFEQ25ldrlXFAbxFj48rWxLlubdLmVX3doXLke472ndfNpnx8ASv2Kf2pKaVell
xygcv4MbDLSQUna2esYL0UNSrVe9DiKpqeMyDBfFFGEj5iUfmoqqVTz1XxdflsM1ZkLNUwgr7KwN
qQcWVdCYzQsZ2RTWbYlmI9Lc1XafwsML4N4VpB+s6fPH7rxmh/7nKb/VZrval9Bm7MLBAoq45T9X
Ipz/kNNmy8okuMWwWTFnRLhHQ4Q0/li6aEH4QU0KLJpHIBlNSGxajC2cPKg9BfHqj+XSCy/cSW+3
cdE4T4QNHOiIn88ZjRhlsQR4jCoHiv8d1AJZ/XLg1WXY9/x0Bt10CPrdD9mcbKiZ+jdKvm/N+rF6
vJ0vyNtG3y8nByw=
`protect end_protected
