��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���-(H�襴5&�=5�)�$�a��S�3;���@�7wn5���z7/��,���z���v�0d�<m�ݠT76 R����%�i����Yv���P9}}�e�Ϋ~�ֺx,�V�K���cbQ�y��j�v��Ax��B�*���Ħr>��A'jv	��B5�?�j���zVEV6��wgxa`*���W�w�v�+����y����+�#�E�G}���X��������)�9mI��<_]v&{��׬mD��	�>��f.�/��̝2���`�4�Ӕ�%���C����3�������L(���2�0�`�������#t��'�k�Z����@{���5z4�
�4g�wp�j(�j��Χ�������%ܐ���?�A�x�����(u���n�RSd4�D�6���~�+�/�d	�2ブ�j�64!���q.�l�u_�G�����VM���_��lw���P�`|�|�?en ϞN�7tu,x�)�\Ă
Na�}���$��U��؀�>��A9�S��8O�^���m<q�!~�u�Y�"��O��c���$���k w2����bs��&I���`_�~��â�nw7�Kމ[���?d������Z�i�}��v[��}�%X��1�ݕ2�y�Ƈ����%��bv�P�}I��'�h������j�!�9�T��^��$��b4���DA_�Mmi�s�d��x�M����g���c�зUԃ�����u&���|�b�Y�	i$��+���fע�R������.�Sg? :������jJ|
����W���ؑ���'p(�|1�B]������V��J�L�:�E��A�|��P�^�أ	��g@�mJ��7��1���5RM뾸��-P�<�P�7RI��?�.N7�-���Ȣ��M��9�$Yo乼�#�� &��(S�=���Y��%-�T;���P��,(�Y�:�q�E1lr�[��	�U�`��=�j��ፎ�؃B�y�]K�ŗE��gL1�/`���9 /���0��pU/�祫Y����a)�9n@��
_Y�{ J�l��_�ܿ������F����$���e\��;W��Q�a�6N#�*\4���0�T��/�p���_��~�^)���D��U�({2�/�v�Kg8�v���N��bPMY����r\��ҢҞ�����O��Y@Z�#��H{-z�½#FI�	�����96j�G��+G�HK�T�&��p��?c�gSX��ȇS?���k���λ	�RYֲ�cla�D1���Q����K����+=e����x�E����,�^jä���wVdr�,P��D���6\�pŵ�T�r�O�Jf�D\u�`i�1L\t�B����?���^[�+�n\ez܋*�%�(������c�}��#�L���ˠ1��~��P|Yp/�V����ag�!խ�pJ8]���Q�!��妉#ݘ-�tK�r��W�Ǎ�V�=�����+'RˢFM��Q�����qY�Oҍ��C�� ��g}������N��f��{gQr���U��ƒ�J���<����A�uсR�q�udWje�~7�Ga�RC�݄�����̅�ІB��$���J�DL�O���硰5��&���؅c�f�p$a<���@-�o�58��Ʀ^�N��F e�^��ߪ	��8�e��Q(�m�C��-�VB���|t9��D!{�ʳ!�8�*X�Ra�)`,��u�+E��$��pΞ]N�i`z�^�u)��d��<1�³x<���K��8gODL���g�L'X�^��t�(�Ə��6i/im̓&Z`%/x�|��+��%t�*��QF�]��7Z���A�����wdQ��$b��4̇_���<�n�b�V��\Bp�����Ǿ^������I)��I�/�h���ܣ/�HPjh�93�0w	����*A���zv7�c�1	^��)0[3��;1��5uJ3����#������s��.gIJ'[�@��(f�%�"C�Ss�Ή�%�6�����e��MyP� �/,�!<u�֖�S��q�r�y�G�J8�Sk�Ap���A#b���Hz��{�ʇ�����\���q�\v	4;�O/����K��<5�c�	sQE�`D�=Ey��]}�X�r������=e,y\5y�����B����Zo����j��='M0��u�Ix
�9~^b��[�}�6ES�_��p��!$�3"�n�D��9��8 ��$F*�)>�qJC�]�	;�=]��r-.�Ț�'�/o�y�����Y  ��MBAO���w�~�BѴ���:�-�qŅ-$�j&���������P��tr{F�;qI�K��P�n��`A�G��e׺0�4XU������N0�/��$�2�M�|�JS�7x��B
�*��� �6@#��5��N�"�2��䣜�:r�-}�c��`Ʊo��t�x�{~���V����ʥ���Š�3���ٖ��#�E�ß89���#���O`R���}�K��+j�:�jT����#z�Ryr(��,�ؐ�r`�Z��	���O��W����A�C�z��ǥnOI����೑Fol�r��pJ=�o�n���q��~��4�{�7�Fum�'��H�1oD�����i��o�Qg���2KW�����承�R]{�ܪk)կa����7��0���ץ��Y�a�z��^d��i����q'ӳ�M�U����E�k�A}�0��
�c]ư�%��������u�n�NԲq�#jщ���FT&��T0oy_"=8�H���H��~����'ǂ�u�!ì"w-7x��J�}5��l�G���]A*�\2�C �V�L���̢C��tb5�_���P6 ���>U����6H07���bK}�k�K=�&Y��p�[�q�ST�7L�H#*|&�g^�-�� j���n� ��Xw1=��Ǣ��i�@t|�*�&���0��@J��ƚowv�)_c��Mӻ#& -,	p$n��:Q\F�A0��=�L��K�5"�>#��+�� �Ʈ:�r��
�r<��d��<�[K¦�*K�����ߣ͎�鹿ls�B�����C����L�	I=U�״G�˃ �y��f���7�;���5�~ۨ L1 -�]�,Q��I��'��2B��*�</8
n|4U^�o% ����K�C��dS��cr"މF���Ç*�0V�gC����G�ӊ�՛�}�3Ƥ� B�h�{�f�QU�M*�:��E8����%�N��+�Ғ�����;��b1�s�tϺ��E��ⷛ2���Yjr���-l;��S��_
�B�¹�����{ڥ�z9ԁ�KվTG����Z�_��H�l�G~�_7��TA�Mw�*�~;n���{`|�΂�vK�2�PdȒʔ��EF��{h�����f(&����7��
Nժk󊢤�T�4l@�c6���L�S��D��)�b�'��F��8̶�]�mj��R~��W(���*���[�������OM�����tL^���p���̛�ԃ��ϕMm�
���$W�8�����J���_u�/�V<4(=�N�%t��x� 0z[�ܭ�8��57�y�ioU�Ŕt��Q�n��k��L��Rh5ni�lE\�R���}����}�����ZK�Q�~c���$Opj��K@�"���"$�5������T�mz���252�_8{� C��@�ںk-�~u���-K=e�K���(�_�pQ����SEC�!�￸��!N���k�!��u����*�����S$j?��+�-I��� �X\}F{�-�0�<-.7��&|=�u�wjxH����5 l|Y_<qqB0؃��X�I�&f�%}�o�(u�wbFð�z�����%+�֪�25a��Sv��بF�5�s�7��P( p"{_���~�m�:fK��MY��,y�>���v����H7����dYF�q�����,�p�|�I��7�	�z��b-��2K�[jxؕ�!��,���)е���d"~��H��-�{W�:��I\�jn�=:�:a�2�&��^U�'r$_F~��mG�pSV��̚�<3�!-�5n�nq���{1�6�F���X~�b*+.�/�:���ǻ�~��M3-�Y��b]�s�/5���<�?ʽ�"o%��
)�כ3l'Y	0�j�|�S�j7g���xe�
c��.J8V�iMav��Y�q"��9Zj��w}>�!j��	1p�G)y],6|)yOPSU�/� ��ńu�Zڿ��A9#����ե2�T�f��
$��S�3�=�H1�y�~H.v[?W�#�D��P���p��kFʹ7}<rw�b3b���U���ھ�g�������(=sC{3T��gRw��Ѳ��*Ri����NX�SQ<</�)����@~=�0�����bSb�F����9�4W8KG����vm�4�BU]�%=�z���m��tgL�=YkB�YNt�1��GU�gT	�f]^pʋ�\V;�vƭ���	-缓��i^��R���}�x�x'�+K��/�j�~����S��6~�Z��o-jlx���$�J�4��ٙԛZ5�%{1�__�j��ٲ����y��53��J��+d��CtNe��:�I�|l�ֽ�_=N ?g4�^�Hӏ� �T�!�eg&9k���3�þ���NK�x�����]� �"{~���=�>u��m�d�4[RY"rỳN+d	|m\I��"�r7N����q�h�v�%��J�|�G�f�o��cF~/߉5�G򱅎{�J�o�����a��#zm�w]�N>� MVp8�i�3�0�n���q	�4�LG�H�Q��Z*DP������(� J���[l�ޡ
����\Nk5��'��w��̙
���c>������b��ՠ9�z3��v� ���E�YY2�/�O���q틁N��=�1���y���j�!G��G��h��y�#��z�*�|]w��������QT��̈́�)COi�����@b��l�����O����o@����$��k�lo�w�8���X[�*�|�,�t>i�ԀSNV�f(�3�C��)�߹��<�*B��$G]Z�\�z<V�����<o�|�Of��o���J���U��?O�T��@��kxǡV9���dZ-�A���˴��N������G�
�*��N����m "ف�ha=�Ł��¤��%Zz'P����Ң�<�/�'0�N���e��:3�'I����pD��H����wIAw��JE�P�4z�ҥC��|"?�����j{#O��p��4%��]Xu
��pÌˀ��2Qp|��,�����r� ���F��UcmU灮��_�6�&/W;4���>q�*�W푃eF�t8�W�O�����W�U��Y6����h�u9s�Byxjp�:�O2}�o�5F��ѱ֙Ι�A�u%~p���Aw�Z�۶�܇!5�nj��
s?>�-K��C�� t� ?/:UG�2�kҕ���5�/m�t�����2=��Ke�w�I�G��yl���ڕP���_������˄;��� �5
QD����0���6lg�e�Z	�S-�zO�IH����9�����&����+@y�E�*&����x~�>�m��6k3��n��rήB��ٌ��X�Ǎh��{̴YB�k�O�\]h���ޝ���j|=u�ݑ�/�	*n��N�.��v�6RKys������:5��]�,{j¥�r������{�����3J��SML�Yk�Q2�V&�-H�;�H�yu6,�(���S�0L`�����]�-)���%v!�b��8���2�����K���)_��S��nW�=f�x�EY��l��}~�3�M�kZ0�R4ا���isKq�!'� a�1z��ݧ���.���cM�gt�9��� �`��F���Et [�!��Ff@�i����$�̆�W�?x�j����<Cl�ԛ�9Hņ�~�J�M�� �?!�+.�I����������|O��/�@e�1.���xS�^�p�=�+�#[X�6�N؜��3��r��6\{$2���;��S��ɺ0�����YNr�[a(�>�c��Qj��Uپ,9Îw���@���o���a�A�i�R��H@}�Q��Ct�8#�o�(߮�%���8����xq.H%�DK������4׏�3\�[�}p�RP�V-F���E��V�oo�T_���t�}�"D�'�3�<�Ob9�+�@,�Dg���Nv�o��vS��S�a ��H�poD�/@ "xT���x3���izPY8=�+X�1��i1|Y�|G�J���.֨�����!j�h3'э΄�����&��y��b�
9	S����Ln�.��Y�vb#�yĺ�Y%��ì��I�G ���j\(��4��ݿ���M��]��ވeBW)�� �ĭ�Y�/>%�S4��^oǤ�������IlJ(C�|I�I�	�T�up2�ʨTq򥀢C�Pp�F�	����F-�U�AU�$O7�(����dM�Z3aKu5��Ya �~�e9��M���g\??3��
������kp�l���볗���!/#ɱ��<��*;F��q<��X��H�%7�����Ͷ�Ð��X�������/��k�U6�&���$^_�_[��A�LaR�
�^E�O�ͯL�Y������H){(XT�lXW���DC����ZߩZ��G[�z�铏<O}SҘ�@s�E�$,6t���G5պ��Z�m4��%u~ӳ������	g�� ؒe���D�A# �nL�]��V!���`��m,&���M�o>dYI��E�9~�d���hY�]o�ωc�#s���n(��H�M�V�(<�0�߉�Ė�\��ထ�m� 9̠Ɵ����~�~B����V$��#n��#��J��-�����U�1=�*���h	Ds��΋���[G�ٰ�8�P�?�C_M�y��ix��V��T�W`m�GWܨQP-'���&�'&�Z;eIJ;Y��Q?��|����1�v��?1��{�E������,NN�lD�*?`�&�tf��,0/D2�"19�8���'ϟ�?'c�4�L���ls�l���bW��
�Y�m�N�y��=��+.G�Qa���+�g�o]5蓱���5:t��d����[��jBAo
ɡ���5.6�����!$��D�	�-��(j�b6��NO�#��� ��(�?-�E
fB�]���؈[��dmC��ߗ����21ܿ SL���2�6���kib�q��MyhU"5�݇���Xq�m�n�����f+���Rh�ՙ�~��g�1C��n��t�7����h`  �og��eJ�h�bw�.&lķ	t���qJ�%#-̼v�&6�S��O����`��7��7��$x� ��!A���U�{�/�wD�g�S	��@���w �گnɁ��E0z~D�ȕ��<��gÃ�g+� ӱ������v-֠L���?{��<�6d��l?�@�*wH�)�\�`��}�w�?	O�zr��G��`�v�=l�����)� ���y�h6�-�OZӉ�������C��.Q|��������kFc��#�8�����z��'Z?����g���Q~�˻��O�� ��(���ڋ� ���`�#D����a���G�Z�-����@����A-�A���!jl�+���Y:qYQP��}g�<˷�`�Wu��c6+P���vwm�H��<�^�{���L
dbO��9D�E��� ىЂ�&<����W"�^��զ��6��T\G�,/�D������{�c�w�<�$<R@��x|��X^�	�&x�1��Oq�~72�y-�&2S-
����� Ǯz|���&Nn+~g�<	�=��H9u�נK�����-�����=}��_«~Rv�C�S�B0e0�����L��ڴ�\k�#ˁ`E��o���<�1�~}g������h���lj�za���`�v8��蹎ئS1U�~'v��	��8[���2����qn�K?,�9h}j�i�i��,�G�jY�f�Ty�����=u�h��k��ǧ��È��C�>e���,��+��$�J�(�ۥ��n�d����Ka�F�[����W�cØG�L=�Dϻ�mi+3zk�[��]K�m�h��+�]��)e��5��:?�l���L<��c�8�N[8�KbM@2q���z��́��x��Y7~�MOX8G-Q��}T	!�#��{�4r�#a4�xpgN�VC�=б���N��m5��z{	˩�R�t���)H!���{B��J2�;�J.�����]�ur
�P=�;ji۷J�s��yipd�|��t���8K��/�<8��A��N���a�l=Q\D�Y�E�q�3ȧ4*�zϏ.� 
��8��@�kwY���������F�m�1�}6��^�g�12 �G`���Ѿ|��F�Rh�B�Ѳ'\'�bH(����2=�]a�C�e�rgߚL�&xz��^�{���M��uP��S��u_k"�ôR��u�J���.���w\�H�����W�~�A�=�Z侟���bG)�0�"9Wm(&e^��E�>��4A17t�%(q���R"��Y�5��A��N�T$�q�LZ���'
l����l�E's��`��]�6�s�G�z�Hӫ.��j֖ԫ	q���u�}�S�Ô�������A������l�u�v�����離��?P���y���p��,���m��Vq��/�u�ry�@�=Xܿ�<�u�#�T���Z:��LdęJ0k4(�V��q���v����ߋ��)7aU:@��5`��x��y~!$�?�҄$� ����	���" �Qhs|N��g���NVD��|z��F��Kш�w��x�z'� �9c�Si<�w/���21,�4��C+ \W�!�|X <�.z]v��tń�2��Ce<���U�q	}Λ�C�ޔO���Ni'�R�������#�Z� 4wJ�)R)���JQ�X3����Q����h�����_i"8�=��f��N��u..2�n\��U:7�9,�L�����zcxfQ^�"��+iiJ��Dt�tR�r�1��0���B�e'}n\�_,��|��3]W�O�-\�{!����C��ō�+ ��{���`)Ş�w�7��x29�O���l}&�ݶ����H7��`���@g���ԉn�(�Ӷ��ް5S�'k��*xs��}�"Y��]$$	��j-���A�<�������cz���60��J�/�*�_��6��:�N���^�Fv�Z�F�����{~&Z���t�����Ur�5\oP�S���2�E��$����m�K�c�$'I� #-F�����ډ=˜G|�mf��/���{f�:S��b����!��	;m�͚]ab�8���p�7���k?�`���(��K�r��ҝ� "_2u�w
���I���@�M�qscA5�:Y�I���թ�!_/�n@H�*�y����!�,��՘�`��T#DgÌ�ql#��?�P�}Y�
��<@1a�R���<XS�S��]�s���4���������Z�B�CD�S�'������MG ���H7�Q6�`���}h<�e��c�J��Ќ��}l��l�=���E!l�B%���0�^`��)	[��h, �m��������s�P��;���a�7_�?���kR�w
���.�C�SMi��@7N�0<k�H� ������܉oP�2N({Ө��5��$��K�\V�<�/�1���P8#����'/VWP ;$Ϣ0`� Cm�Q{N]gL�ȅ,.^6��S,�o�V8b