XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��B�����2�{���F�R�/g\���H�"d��n�OJ��J>�i�IM`弆1��S�;j�)���[��gќMn��Ӳ��2(�� b�� 3�g �s��,�<�}ӂ$�_W���Ȉ��C?�X��
�>,>�+g�����,���cxK#Aѥ& l�1FI_�c��`����Y��k bV������osR�bi!}�^������� l����]��h�F��JEb�9��x��e^��/��h�B!`/_I��s�!I�NL;AV:{�R�sR��u��ɖ�@�ˠ��@|@��A�� հ[0<��R|��Х,� ��eq������	�)6?ȑ���N��pQ��*�N�\��'�n���|cq���)=�$��R��[�6|;J�u���)d!c���*J�~�H�2D���ɷ�\h<36�pլ&��uIe����vG�s#������7�J��ݱ9�X.�5���0�{5��7��>�bs�����jF&E2C�sXJ6X�A�MO��������k�������!����J嶿���AC������Z4^"0�`s�o��x��It�[�u�I!�s���,v����v�W���K~��^�������Ē���NJ7سC$�����^Z� �"��\��F��uk:N+���<"4�b��FO}�~,!�!���?o����m���0�3;��8xjH�3�/��W��b��r5�X�9�0��8��N�����Ѹu;-XlxVHYEB     400     210�|���ӳ|*�4�)Po�Q�Y�P�V��o@���,�Zd�_A}���1V'�8��1��K�z>��ސ��?��)�V�s�VU��n� � }����S\��_j�FQ�s�'��Rc��/��?1ʑZ�c<�Ӊ�;�LŴ"�jR��6!�|Q����i���-}qHU��BF/�M�K�6 �]�Hs��ߞ�G��t(��Ɉ#e
؃�f�GT�.:6��99v�\\���]J#M�%�{�2�V`lv&,�	3�w�" `Y��1wQ�u���$	f��h0�΀��(��.l��ǃ��@���R����O��o.�՗� �rlA��j��i��;�2(�j����-@��E\�Ǜ3����#��1�zk��t	�z�H��F��y�D\��J-�Y�zA��w�h��&Y@Ֆh�r�-8x��^�T�@R�n��W���Ⱦ՝D1����s���v�_䝽�9Vk�>a�bW#B��OO�nY�f�����PU	~��v�M�Z��,M9F��9��DȱXlxVHYEB     400     100<=¨1�'H<�l�$�z8�k;%̙���p����-�c���X�Ժٓ� EZFX��,���0�:�ȵ�):�-��}r�n��o��њ!uOιy�e[n92�R�IJ�{[ɠ��gm� g�-+w�ѿ��h��-=�����vM
��#p#�|=�c\u_n��S��'W�u���%r�<� �,Q ��f��#@��
,ex�����d�s�vo�����q�^�z�F��}soH���bC+B{��W�q�q�V�%�!ݘXlxVHYEB     400     1f0tC�������T�M0��-�Mxz�s��:S�i�,�+.�������7��g�;�N˭����>�_A�PpS�/����D���%�*��AX�;~�롞�n�A<�v� ���qN���.��J����*`�i(K����"L��Ҭi��
�=�
ߞ"w>��Ђ��P*����t�'DE���,�F'�3o+�j�g��}?m�����'�8rD�������8�����	sF���p���u��*����+$��a�d}���m�P� �!pر8Tk��]�ާ����:O��A�X�G*KƮtg_@��T~л���0y!9����"��rm���(���ء�J��+� �����%ۣ"�kƀ�u�p�9N���X���:������W4,Ѿ�,�xH�.�B/$=�\��ɬ��Q�us���9r���[� ��x�.�i���}��$G��+:I�����y���&�Є��8 ��h*��sa��%&��XlxVHYEB     400     230f�̷���x�e[mS\.V��M2q���G�ap[���>gi���V'"en�D7�Dk��@�
-�nT�
XD�\�3� N;@�
=�j�~��j�漬s��C�=��~����ܾ3�BW�Ω$�Y�8������4�77�nC������ٟ[�e��O��˭c#!u�]J֟Uo�g+��.��e�F�]�J�Xn�hLy�̠Sit..f� �f��㑝���%_�M	6K���ͬ��t�-��L�Ҍ�S$Yvf�h��hZ/���v]tChޠ��/iu9e���]C�d}��q�N1Ys?��s5����-W+��3���qsROL��,?|�C���ң���9�M�" V��L��M��-赸�ZW��Y	��V՜'y���Cڍ0�m90�i9��ß��$"][�A����Hg�ԯM�(u�)#�N�;8��`M"�Z-�E7H��"���o�3�(¼.���������E���������HwX���<��DC��yv{+�YcGn<u�����x3��^�v]T���\/2�Y+�8Ƃ�
�a����1�7�|�"�r��{TXlxVHYEB     400     1a0ȭ�Bi�o�N���|����3ψH�{	����=4QxT ����r���3MW�sm;����*�d��ĵ�G������|�랓��¾dN�Y7���S��C����R�I|�'!P?�
jX���ڈ`5��rW�؋�|jt�r<�m ��:��	���I���ɖ3��8�e9���Hec�r���5%��E�)��MJ��!�Y�/Q]�c�G�<	r%Ϟ+5��Q%"�L�ev>ֵ��[�_C:J~�2tw��t>�)Y实���!Fޮ��g����b�ܮ���H`(�%$3�奒w!��<-��jeU�D��b�6bP���uX\D��o��(fh1�X.n$������
��;�z�_�`�������`���w�51�ϖ�i]�xe|��x���a4�9��Gh�C�vXlxVHYEB     400     1a0�������LZ
8�P��w�ן	H���W<)jY�O�ϳ���V~��V�a<~��HYڼ�w�k>�5���� ��y0L9L�ց�$�Q�7�	3. ׬��Gλ3�&wC9)!m���}�N�b,�7$l>���ŢJ.��]6%�h���+'�B����+���@)Go+�y�M*�*�¬o�/��[,�Y�;c8��X7p���I�u5�Ű��k:�{~�а���O^�%��^ö�ʷ��e�_{�tѕ�pg�?�����J<��$������޸���H��H���=*�ȘR��O�!��%8��/1D�Q4�Y�v��6�h�G8���X�Zyk�s�QpM�����j��8y��!�@��:��m&#��f�=���XEz���x����*�J �U���HPXlxVHYEB     400     1d0�G�ua1b|F�VX$�ͼ'�Vy��x���f�>CSC��/y�ӵ��
�������%�bJ��u��}�����K+;�O�&)���h�\G�h��:u�<��o���L�5I#�ř2-���6���3�xp��UW�?݊+�-x������\�ع6j&��_�k��$�'%f�eo��	�������m�B�M^hmo)��r�"�#�{!^�8�uQ`�ǠIn���BV����2����{ǐk�2 a�k�}�`9t���۾8��	� �A��H�R>�0K�&��i���5kg�Ѹ;�Q����rOIGꍭ}���i��gb�ul���|24p�լ��r����~Z6��˨��`�?h�"�{PNf,c4�M�V�tE�/��/U��k>n0G��K�����@p��O��H���G�ܖ�Z��*L,N�������ƀ>}9*�XlxVHYEB     400     170A,�Ưsj�9�,��s>����z�xj���t|K�i�*y�CI�a��'/��F?���h��&��˄�աt�0"�������m�q�a��*�2}W�6��GS־fb��|���y�l3�f�z���ڌ� ��ՃI�cb�I%!�9�`�q��#�����$��78���<9T<��_=�ᵀ`��V%�>�"���p�: TS�p?Th�g �P����Vd_aP��9��n�~��U(8������B�CЛ:	�2�b�Љ\Nώ�����Ⱞ�=Z2��:5����+��&�B^!
0]��p�Z R P��וSB���B!���*>=���o\2%ݛ����0e�Y��@�ob]��4W��5}��a� S�}�XlxVHYEB     400     1c0�v�-p���K�)��kW�pI��8>�u�oソ��Y�i]�?����v��
���"<hl!�mD7��=E�
�hp�w�"�4�X�'���

g�
,�m���<����!�@;���P,X��f��0�O��`�*5h�tܦ�.�^،�@��9yTl�1�y.-
�|K���� =�5?2��$λ��C�3}@����+MHqw�򙭅�Z��-� ���_�� �����Ĵg���:�&q�Hv�����(�7��	0
 �"��L�k�� �Į>Y1�k�����Ĕ`7`�R�����s0��׸�Uk��Ѥ'���$�;5�x�y���f.�*h)��h�0@�w\�r�=0��	J�V2�^PB|��}^ܿ7'	[���v�N�vt�#�ߓ��{��w0��=���t.�gL�uE�@�9)2����a��]���KXlxVHYEB     400     1a0�}�y,�@ 0y�v�,�et2T$E#Z�w����Pm�_ЭHj�t	*}�g|J�V��4�����V�I��io:�b��V�	�y�3)�oqmN�A]��1~IMD�m�]3��Ǭ=D����ͅ��uLpTT�<��$�����ƴ� �uq�~V�4������v��-Y-a),de${a9���5|�[���0������ɿ�O��>K�IH	�ܰ�`���t��=M�,�3C<��ٳ�
r*V<�s�>o[��X�L�t&آs�AdX�2rq��s�J��p�Β���+役��]�k��ލ!�M�B	 @�֙X��F0UGԐ&�}�/+wd�KWZЄ3��f�Z*|���\�Ҵ٪^�5^Kk��-s�a������]��.���l�(����/'6�[��$}XlxVHYEB     400     140�/�+�����龿I7(Su�f� �^m�#�d��bD삆D\W���-	���cTK͈g ��R�t3������W�[�iT������D��Z�.�����q��}�;u������ �/#t	��l䶥D�'�
cG���L�����#�y�Yt����v}]���:
ߋP�i���{���$ɾ���T�����1��@�Sj�}� �:�F���)M�ʒ�1mJG`�iξ��:�b�*��s�/��S\��-^���OrG3<sY�ޮ��)����ߣyNiM4��>�Aj�R϶�ua��ؒlR�~DA��[����XlxVHYEB     38a     180
F������	���K���f���Z�`u��j���:����z�;����~~�cv�����S��PD�LBN�U8�C�Y�w<iu���xC�q���}��������gj���!6Ud!fN}��!ɸ����V�})�lz��Z:��C�,�mI��{��w;suQT ڣ�S�ZV����8"砧R~��<�H?�
nhCa�6<a�~�|du8��VS[��Ӥ���"�CR�N��f~X4 b���e4̨�*�Cd���~�6��|�6q� z�ͦH�{���/�VF"Ρ1詾E?�#6�)(�4bQ~�9��;d�_"��-���-k��H�܁�=|��N�V���RmI�W��D�x���@�M*��]��ް