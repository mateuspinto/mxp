`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17472)
`protect data_block
tTJfpJuhLqV634uBnMj1dxl1h873pUpU5rlLz2sAZzaUxRogokfUl4Q79nTA39JD6nCRc2cPo3Pt
IW8+fyE6YlEPVlaZDhvlOVI1O8ux3EaT7wLFGwQfOR3BthLZh0KFUBTMh6ksFbtvFb9/PCMYdX46
XCJzSmM3CHL6ib0IUY6YejqxsCDDtub1OA8yYlAkr0vB15nCVci0CFiBkai5vDtTricZL24N3d4U
XyJtMD87sZsohVFzKBcnFBlmSM4OOgLIwP7eUPdNX3jgSULlcXte6kWTdILhoSetAgnNiyRw38Jl
LRK+DCeYURKGOTWTciF4FdJGTszw3bN+N3eGxtd9xGMHtnryOiiYvGdeh9xPTlVyMfGJAO7TsvJu
3F/QDwMNqKTe/iUNlUQP7f18dec4OBTQ8Ku+/hKOoJ/+DaVEkxSoDS3BZ8cCRoZQ6EQ3/2j2hRUh
G+c/Df0BN7NfwoLJhLGf6X99GA/rdofVa9jmiS11ZOUFelxmK2t7raAAAOlE/G0GFVcvtgIY3toG
9ppmuzYAVoU6WaM/cZdd4altFoa+n5m/HEtIK3uh1Mgva2MRPTaKMhFkM6jAKyWhgVVrOyGB1Ndt
JwdgtGLYDCggUxLgHvgGo/OZGG/4X9iAqfmONi8M+SyTSC7JfATOBbEd4DVlDQEZo11qHu6Kqb4A
OHvvk5cHRzkNoJSf4rXVasfAp6yNOgdIyvn0QSiv4Dg/4rkbYiVeYRyUT3EoZ8XM+Cd69rXpeAFH
Un9g+7LL6uC5er55eFsaa7oarBiPAVq0HroXeVfpEaXsACT/Rca9gFsXTcgOhjtk0l/9+bca/4Vw
5He0GN0e7JUVQC+fuMVF7sfnbq3Gvi1dQ0nTFG9RpBvhWUvwKRjh7+/Hp14sngLeolCGOoGmI4zK
8h0AaSG/uyuMzUq+2GGAXcM4PfMAUJbVBUi9ozTOMCgp23xYD5kaad8WHZ6Sl0qiiKON/MwHGXVT
GmAlBBQItPjFf2CJzSCO55OFusidSYmknMF5EKa2rIhSjPV++Xgk0RQdoC3BR0DBOZYzlfZ9kl/v
1xLMdp6ejBKIub2IbxP5I6uePz9ZjAX6TDpAsJV1Hql1SpbtzDxYI6bJ7MZNMMPevwwVoafyKaW/
shmTi5EPqzHkGJrEcR6l/UUT486D9sXp+ihaHgov//EDAJWK86mACGvTTU7Z1vHdbmIxU+xPVqmP
lWbRpQkndW6m8XIAppGkkFcqhroy/Mz02z1oPKUeTUBqUKiJVMibH1E26DdjuJBUgqY9b/ifhLGK
TLsJhbjp/IM4ED5nb3W6hTmxKNqK8k6kTriQx8/Kk+pC368QaMrq6UzzsDImN0OiAVy24kmIBUrb
+TwjB3AkSOV7WyZts2gnTHY12PTLXE1TvUB+LYmct+NcTgpEkKULMzq5PF/6syepL5++gJnJcD7N
ursWdl/VMaut26QdMHvt/o9V8/ihAs7XCnrKeV1BcB/IrT0Ckvdjqr1mYjsBUx0TeRocRPyIOyEl
8xrqheHnUGqx2AhdkK+E8HceFF9UtO7R1VWKkfBqtzzcAJghuioHiR0yoslMUhqHZc63vuArdinc
mHQRsOv/WYrvN85QTPDAMuFQCuzJwAGkhHO48xstTqMuYQkTciXfowHUhO3a5hiw0QatpCtnCrYv
B8b9seqVEOT5hBG8NPWcr/Jme8bzGFRkSE26rDdqR1KPsDW9h/NnC6i1DwXebOM86Oy03Q3l0Y+c
hvis7YS2QgkKZLE+l7fNdyXb92IIcHR0jGx8Iqth7t8zlC5pzpQN+6X5T/aFzKevuBOR05q/w8vZ
R134T/tVtLMZvj4nQPWJ1BrOLL33d8xYqbWOorXcrApZuch6hBkIaxP3gizFqDkEczfPH8xrZiSk
WYguVlgqHemgQsNmZ5J9efRyWRY03lzzavYaJX7+tVZ+1h1E/mfJaCKerZumXF/aG0lQOOir0Av7
4WxWSsxYlLGRa6BrsjDrgei+Q9BQI0VemlwwZSUYM+ahonkSPGjizPj49sWfCGIlmcTHl7Ca+Opw
DGCE2iCoW76jNsyP79m7DcIfM/g8tWJfUPIgdfh+mFZmw8qe8zHZ3FfSV9nngQq1wMwRExxl1zoZ
QciDMUAm/akZCeTIvOiEFnoyeMns0Da5T5JUFyVgTB+xRyOUsC+xCHI/n9CfspmKzaVVOqL4P8SL
6vDFzY2y5BDuJpjxMvA760SmaZCZC3GgbxWfulVKzr4ReclP+ZKuf3nzpKgVKMOUz70ohGKCs6zu
3bOByFrGtbZuo/c183oIH5aBHOELSu3rqCm76Vu/kksied2LvjvPIkQh+iuYAQpF8CGnBLOlDkzH
Fh0xVQiDee7V/JIkJJEOmLMb2DInVQX36c6U6bpi7rxc6mw9rMsyD/U4GdHl2n0WbaTTgCpASDQn
v9BUE+x/lNAfUFY+yZAVZx+Yjzf00MRAORGjbtzmHh5GprcSF/2Lwc7ip5qa7RIdwgiJiW8LsgDN
DSMxmnSzyWSDJzwTn4sRBvuVnzOqlLqMBHGAXrpMRrGO3iN/Evf2K0022AC/LuaANf64U6mK0rBr
IE41SO0p3fxfHL8aoTdEdPqZw0LHDHB++PF/OOrKBCnfmxxhm3pmBbBn0HQ+AHz0HpB77ZlVHnPp
Ch8BCJ9/S7yFwiwO8bVuZjdR20ZNPUBwPrSqxUwOawGQM+WG5okBb6suZ/XLT88X0KD3y061p/b2
b9rke5e1JWqS8isBqdTMrBjtPjewl6D9tvaJjFsvan3U368GH38vISSO09fVqxMgOBNiTNt9ocvq
rlqEhwZdwLxQCTsLuLcUEGulxD09+NhZCVqlXoZeIzIssOBVx27uJNcjVr3AQ2R9d9GhHTd6F+I7
SwB6N121iGrT10qHk6NGeQvinptqzCF92Ob3rvNeILDbVOAzZpZVsKklqiTDG2Yy0/1CI+NW3k5Z
P+Bca87pW7lUkIFioTaaJ3c3myxTdp3Qj294XsgQMUXerdTLvt4DNWgKx/TYS8LChnwGm8eP6KSm
RlUyUZLafyHSzjrfy/KfyU6hW4L7PJgKRIqxL9kfbn1Ndqpn9PXTqiH1TbL2Db+bzU8w0sC39ZEO
pq1AaM0Viyqp7DOC19NlLEjkKND9hYB7RTrTJMNTZJsXSqxguIkuhvf4x2WT7ukY8mCKK08sbls1
WH4ohVYUnR6wsnDZvdo9qB7HWCf1+r5JCnc/WmiUzWrax5/LqqM/75twZHbARjw/FzWtnw1PXD89
MZ+EEvya/M9bVxK7ams6q0xKhs9UqKDRMmv+ZQcq5oNvVuCYx6ltCZ2xGT1xdgZ1btv3ay6b3F10
fMvqLFG2Z5bHv1NNoYygQF9KkpbRQNwaMVbfA3LVa0liTKBvtPiBPQQIfdxX81dYxfaYXEKWvFmh
iuA1RLOBSGV3+h/F13pAAoPJZEqygnLtdgZj8vr/CDiZa5UhGHtKoMnBONVT9zcsxxiVoGtQjEyV
qfAgp2vSTNLis53amv/A5/Us5QdTUMrIkY7wfXwxyElvi7LiToytJXrZfJMAFdQrLTfzOtBKOQAy
TEKnKK7QqiM4h0T7dcYbwfXzIsIaovkeDVkijgnWEJNbeNMyeQqnARQcL9e/mqj3831Gg3ZrW6jt
D2cG0XPKyQg6SfJy60dlq6RkTSwF9AcVdfpbyILuaGlREF/H26LsBsbRmEUiGDsa7noBS78FNSEL
T3/ma59iaEZdKLGVePcr96XQpJUUlsS96o5QFPh2fUdYNHq8/oY7nM+4z0pF2mMfzTDg0Ymwz+1L
fXMsWqV8Fl1Ii1BPo+bC8r6WdczPgohcBQTJkNm65dHnrwxQwRo6m1oXGaxJRKMc43j/1Z/8NpAd
amtOMkkBWBEfM4UgciniHkWp8fM+DBLXSITsSgagVYcqzheGhMGM9bDM6Z8OHComkaUGH3jlIROG
exzvp2AcSVgeIeoxUwLKXMqrWoHH9WYG6HqVFHt4yQ+EBsUr77WiJ/+qHmA0iKNGu+aR+cNsa3Z1
sJhS2dD2U+9gRVccO6Oq4J2XYcmKbnyPRTxR9CVe3JrPfkOfiujQtOmFZ2yMkKI0mSRme6LC9run
IroPNwOwb6RmHAue4ncqYP/RLmTv4CMazxhDdLEJgOdIpdV8hiI0EJB8qQndrjr+f0vX5Umds7OR
02I08nlWyylxZQOEOGANI6KgeqcLCcs4iyx4GSXiVRQcLGbK6U0/YgE18S11tDRigWEBNMhV7zNc
KPy+QiPwUD1Trl7lrE4LLsN4jcoSwFgHG2c1023UnGCAJ9wxi8l0gQkGmIhvsmBqrX8wCxsUVBQO
HulrHzOt/GgYdmSSPOSF7hKWux3X5t4PdcoLlhSCQfdE5mc+//3dp/1GE/7q6SNCCmxOr7wkF8cl
LSF6Eu52Hq4ip9FlWJmsPJDG+4hXmqhNBig18mE5cB0C9BsfMtS3OfgPdwqBBgu8PgxaKIyQTQmH
yNieoNYGPrzJ7blI9J9hpPXqFtcwe0940Zo5HeUpR6K63nm4zPv7DAzjRrj9jS2hUvbbNhivrCZU
p0+P6EU3arwlaX+cINAv0lz/BMpi9BOzzX+GVuBXkoY6DF/1elKA3qUaAjgWY+OF7YTnMFcu/Tc3
hltVvWfzExH2WcyKdPnKTH+E8nsA9fUdrp0IxjXlidSA+ih03NuC/aYDhYMbMEtpgm7j75bBh5kU
m4dL0My7OyJ8WsOHvn66pwVvcz+no+9gX6GE85VyCpn3BGdeSlXvFoirQeThuTMEcWG/Nyp3ZsvW
NsM/qp+4wRM5nEvLR4/akONooEEdJfS/+sTeo/FsO8j4SkeImKp7nYVKZ+BOessJqlahON8sGmXK
AgcsFCn7eZW3b/uR6Jj2Mb2ciLTy4uFlTnUWTB0b4l0Hi7Hbgp2sH8fSXWL66tRsF2YYUa9WJviz
V9pN+e0lOVYFTDrDDRF8rItBVKxf2S64Da8FIYFG4f5ZijW5NQbiIO31w99SglU2Jzx6oAxKKJED
HbFIyr7SXBR+WQ6mLzG6HXBexgeyN7SdJfCtV7rFqIMzGoVMqJ0nBMXEZDPkWUAUfKkgiI1J1T6E
pPVK+W43yzUhOzcrgY8NFyHhKuvBhXlNS/TFYzKCtCuQfCYwVSrYD49Rb+765PLkhUQSVNvDt6/n
DWVXQhCARP+yBd0A5I+YirZuAyAeD3eXroE8PJ2jUXhlbmElN/v6lTNLC78VCvKFtzUZoIJmSv3Q
vIQxlxyCpGh2aU4RnT8LYcXTirpJoyVy/oUoWbjlFljCh1ZiysKCfn9HG3VAaViHHejB+yJiV2uv
KP6ae1MTp+I5thFzs/jJNYceho+80JIQYResKHigV0Vk+c9Ql6J3mPWhTMN1C9mzFifw/wGJ11oK
t76ALVZ5ANtUjPN5GMbimW7TH9w5kJJxE4vwzrTkWBiN2/Xd3brNhLDCBwJab349BR6hAMAgz7LW
fvoJDX4Hjq4GW2T5bSbmPVh+BGUxPUIS/nJTwvJS4/eIY8jWyIlQnzneZj45uXHiNxG7pOfTyqsP
ShWHgcitYy8zqYcJWfCWThTZJzO9QcUEVf1xQ5UTTzY7gd3OAH+vF8QW9bMdp7lknQdKcUgFvgyH
vJoe8DBX5xZkORBScTgaQND31LioPuUmNYgJMlgvC6zFyV/u7OSXEjGFSo3wVdL8aHmjvC58n1Y/
z7XpKMLOOXLFCvKN0GnrJ6/NHzEbh+cpTWhsRHrngi9IGRR9taRE6T7KHQuBn7ECPzNGdVGb03sy
E2pRekH29xO2mNj/SljvUdM9Kq73tqtxyoZoH+Aw0gHr1DHFK8sduka/rwTBVovVkrNklMiDKXTC
f46eTJca1200EJ/1L6xcY46M3ezzZ1E4INkI+QBSu6nl7Utf2WiiiSRHkSQtGi/TH2EMExi7t2WY
Uh4EsazGVA27hE7JGV+eFlirEgwOaggNVQQXrNu8SJ3eMCXjbwmW7CBBGbPMGlPAsGdmsjIKRu8/
u31GRhqd4mP74KrGRcuHrV2asPPmfqcco9iSUhHF+6R8HozTl1bApETwm9fzV29fNbqDShSU5VnL
IpEaTxLHVa8xRVDBVn08+ZpZ/zbyhfKUQfXr+0Sqy/tG16wOm8UFnnYhhPcMkoeXXv7N0p8PH8MO
YCHb4uIo0ZfsiJh71VabPppnihEdLwPLbAS1TM00g3zJJfGxyG24m+tA2uzLExQGWPK/0I+Q4Up8
GqgmU1gS1aC7ZN4W4kekg1OSuPh/YvA6C9ajDL8jC/IH1qMZqkVPEQAA1/Q4uWV7DA/4gxv+Xq41
VM2fW0pKABaxHLd9HcdKu7rTicmoB74Qo18ymjx2i58vwZ2q+W8DSZfhOIoaGY7UdVwYvYid/SgU
Jip9vnDM1Ap5FQoTNG+Y5VCqZUvKHp3ycS7wvDTy0VT47qwZVpCXVFZDeOi6GQd32UcMlbx63Ihe
n3ctnvlcdkq9+ZhV4N+kysfi5JVmkg+nLR2TdmIGaQQDa3kcZgUCMpXRWQGStIXirKABpcwZlAZU
Ci+c9aUqHKNNDew+s5dtV/jgenf3OpDLZM2s+SMCP6z8ZK7ITJTwQzcgJO4y/kIu+xMnPZ5eM85B
zZV7DZEz+g4FUqnibTVF/Wz8/jCw1tQNMs/sPoicg7h9tJpCat07f0TRDJoa94Xs68RnQ0SWI32L
W136ndVj6Nmkyfk4PDfAbaLmlgLoeqZkkj98Sve1xGXsdQBbOGb6DtyLD9jFCQ+cAsRkL5GZQEck
7pvJNMYkbhQp67M+3Eq3oMbe5nRciwE3HwmhBWRxJd711Nf1/WcZnxuyzUR0HSQ4AdytyBrHk8lm
amDbO0h2VFHeDus+pxXO1b05kEnU4sp2UVN3fg4V2W/tyQGZdEGZVSFLoUkVWY1lgDTgxyzdmYsF
i8l2/T0M2G/ifnc1ghUyiEWdHgLHeqagsHO6TXHP//wwKWnEyrb5mjWUXAbPcmDeuZSsyvEaqSAs
mFFq5RH71T2K0Y/zpaUoo5uXcmS4DBmbcZDGOcnEM138mEHq0J6lfeQe1eUya1jcn6o7xTAAJRP1
sP8gmmWP1DLHu1/ZfP5MbhZMU4s1KGoZoIdTWSRCOf7apiNqD5NTVtNb9+KDJ10jVSYvTrlv1LOH
Wv/9eQQG5IicNeJXWS7kmZZcgQ+UEHlvOl9eNxSgEUmzKfa3x5/zoNDahTmAj8wf0yv0P+Uwulb2
7+bwiECdvbY5g5GGJJNm1dRqlNZ7drca8LqYzSu1IA4o98gyBdeSceutiPykNILNtbranrhlX6z9
85tC+9rmlQdIsOnzn0fnB08gdLxb1CzEwyyEMSo5yCYMf5RhWiyuQaAJb4fiAF26Nwp7QYmqJz51
FBF1LgvLttPZqLCBdA/aO4MaZq99Te7K5OS5eJZNAofDv698oPPGit8ZyrW+T29kDbK+/bsJQdEI
njgylFE6IgtzjDhQRjjsB7csP2m2CzE4VaTq0M74zEYWJtLz0bE3mJG2/QOeA1T6IoicL6NAW/5f
DHGRXO6LNYkVcmNmLaVqDcvAXHOcnrjsDotdNrPe3DLYthiiYlkPBw3PimKzJTHq0uYcIDnAT6Zt
+4r7vko7x+Jt9E2L2X7am+tTxNVd5qloFKIGGPdSXoY7VAKG/7OGpkIu341Jv6DbjjHblIYZFTgX
EQqaV9RrU3qboHyphxe7nMFtvxd1vURTPKf8aVerYZyLkgDW/qjLt58uk+Omye1T2SXBRP6xMa/r
+3gLA5bJDUM7DmytwtxurYoGqQs5pE3kjl3o+du/KljAXa5MeWVQz/b/MnjU8nSFiwRE9nkY/dSY
LljUHtMyeG8AfqK2FlgqNWYSqynLbS+Dzn/RrdYZCZzzhwhppeWd1Xqrdu5WkC+stUH/+1X4wL9T
b6X1OmjR5mFiz5LhM37bdwxtKWnm1AE/6hcBAoJvErMKwgfBp+0/EhQKzW5zCohP2BxEwplvUEK+
9QnB6WnduSxskGXJUIka2/5AlE8CM+zCvFE/MOfZeOC8J/Ec/qlc6CRfkiKbcmrKWk5FfrR6qCSQ
bvC46zInwkgcGqaPBuj1UZpn0xYqnLmnTP21zmNAoQB110pAEyvwkV936jacLjYQaaFf7Pukb4sQ
TqIcbb9jh5dD1ekLQCcpI4UE9BCP6hTD4Rv+3C7qIeWqEqk+xFEZMqmLyL2JCi9E9nj5x721HkGC
Cgx7V+tVp9lGoxwi1yg1Zw6ba+aSju4anRv4eXd75VQ1+xhvzRLM2rRF4rD1gX3/q1aACJ32LI9n
ZBBiKZSh2koh7nHxec0cEHGxKvq6JCxAIaasihfDchiYrM18O6ElAB6l5jkkiC3/qrslFjZPyySe
aNl/73DEPx8nTI1Qqz6qKFihHNYWgUGyJ7swaSl8CzYtw1xLsL1R85jtFRwBIWKJ66UWdY0Er5fc
qEEdVaX0oDZjBjdeonAjdr42SWLrYQVJFAnWMch7gOrubyY+v4gy0ksHL1fS/WoBhAtxOePYrXG9
QkZ1M3vWL4gec1xRHUPUqi9V5Bl69R/mZUgkADAicGkY7K/mzj3ND7Bw8J7oE6SxLpHzjD3yuVJj
gsbLJX9o9fdyvIT4xe4UQvBeHEHTImrtCWmeKRtMDWdkVXjmHNBXX1aAxF2PrI5B/3sCJ5I99oLQ
qbxxAhm+PTrI4sOauJBfBIpNujlZVFKERLZkf2erqBCuKsE5W7tE2lU8jJBHApO+9a+tReJpijZE
4PHMeNDRRYhrq54w0OeNT1FK5c4fBC9/9OPR+c7NQcCBz+aeayu1I68G8L6funQqphohrnGmmA0a
6s9mzpXxjKAehuXJ1OfSqUt4Eg5wF2J+0dCA1zcbuWvdHJcGVkfjIINUUNm62cuyqsTROm38ByiX
jPs5IpiMHWQc6OZSMOpdTd8HvaCo0/a6DKPwJcb8K1+PwwpRezSNbvaTCo49mI7unhtrT+RTimkM
lkliT/bqV3/2TDEjmnV/qROO8d5WllDUMkYvTSb7GE904iGn7iOKHZaIDHebQW9j3ypYeB1JYMsX
BSmO/JM1uEB0fin280jROfcj9EZiLDHswf5NbyLaQAFRvuVvzrZNHv9bl/XMQQM+3EPznB1ZWTeO
4pg3dlQWvrkBXlvY+34KCR0OHSrjKRxtkXHHpYy3hW+M6bYskh5cyipBNKMqr2mB05JIuE/4TrqZ
/k19/gfPEYmb/U4moq1z2AIahpe+QG7cXCk6GhkYgqg/EZRHgrJpi8PLoK+qg+MZssv205dXNpwP
xSfS88n5YLJ9fJE+SXAbveWr17PHCTVKkp4tAxNhvcQbdboHVbuLpegH2k1Xnn8KJlgUPmlf4ksT
sID1i9TJyhwH6QJSTZMjh7p9RbT43kGwQ0GRlKajz2p96YksUgl0IUYb175oLEmcFyz61Pp0QWm8
JjmbsZPfMgfRRjt8mWw30rbwW395Uw0ho9ABOuTfUD7OIxfyVRLXjP0SVEUeOCjF11uVM/YToN2I
gDJrlFuOwazg10jM7x7m+9bBocvwuEz5SdPL0GMxzmV/QHjG2MNkZRdmIYgDC5yB7Po2AvLQO7yZ
kQlZxLTIkE3q2XLCxO1pjbZBWR3EX0ptwFWcpLyicwsedHV4sc3eFMA+E1UgPb+9QFIU3XL6FN9G
flCiSmXfZYGxABWFK0e4sSB1829U5Dh+oXVrty5lfimJgaMSUUXkkaak0G/6fCHNfgg6GpZ5Z+0n
IIyVQKulOjVD33cGSVDCArAink6aUE+TWPPUZQ/ojFzVxFB5DOu+O34pqfXx2dsQoAl+OKy5d0A5
/4A22JGJwXsHp9Dt63yiUF1XqD8cPIOBYq8AxNb9/GdqwoR0p72NELxo4h6LSxUUztk5sCsjk1QK
1Wa40LIDY8WaI3OjDJf9+lE0p/Z3mxkqQwcx/ClmcUpRln32uJSzTXp93hSWwlM4weiKYtd34VWI
i4CYwVt1Z7NNYWbA5jhrfIPxGkqNs88balSI/ar8+n734AtlQbp97n+I/IRWubPPVl7FGd0IsWxA
b7Ep37HsNYpjbr/FjY8dKRzkWx91PyxI5RChn5iRdLITmKq9+L5nHyliwgY5ONiKLLBnVS9Ov8Ux
D81/X+F1aFke9AHGvkdxZazG+6PxZsF0KVpeI6Y6tMLxfyLSHHc6jxhKVanRx0UgkQnXwsoa0cMk
u0Qzgi08QNBn6NNLLM3Io6Hy+n5JVeuPBnlYn0WZ1lN8ZMwSeXx8AHYFYewlk9hqWRcYm7CI/q5+
0zUkkmePnKIORiSXp5/lYMF3WuxgmgKNUsRcFjqmas2cXnCroOPJhUixIG3JYZFkr5uO74q4/R4j
aztvirrBs6iWAXjDFUjv4hm5yoRiIuvAWOpxAPmOY9nKkVADW8JOfVE71HHqoofrzG8/6mc5UK4o
ZvWmUfO7W5FNg45ThBPGmhMkZARWk1mqhibwiiX7hYRX9Yce0PwWw3V+zvptPb89cswUPSSb6fqs
kk3vEYntLnFu9H7mdOXGcMzN3rqQ6E/YPgqo4SLfrAiX/3TYLOdIZZWshNujP0xHCUNspTIoxCVF
GSCMPfPf9d2bNUOANqkoGoHHCL5VqL3Q127zsJnLsHRfTG4Oc1elpdMR29NCtblxg7cpGIykzT9m
tc4OaygPpE+05FbZ/wYubGIQOi7OaylCim6h3/iUhdMHb6z1ZaVCigML/OnFzvsBhl8bT/QEt2Ev
aKrVQf3xH40/Sa2MD9MTIZ8stecVjOMLwtnYdBSQb0zS/O5CjwYj66XEH9X0g/xu3nI/f9FFFSLh
yyoms5bjzIDsgeYtWcM7R6G8tdxJ2Fo/bTYlsqQvT4t9TXxk7akpUG/1O6SAWg82g0DSZpbrty33
QDvpiB6bZEGaZdYO8x7l0RzjUAb/HX4PzGry1umAm/+AKRhfi3W3Ayj+WMWwMKsVlLlJSZ0plwbO
UcWkAML83S/Kd2U2AC04LbcGFOgE08E2njuO7HbQOke+YpXJ9HIWdfb9KXWXLjlVXAILwL6ZxGdf
3k2eppptzjD/idb4QxhGjkEcxJxzyAU6vrNcu+sUeZDRlBtR2ffFg2KGCg+5RRDUC729U/JVZT5/
6rOTE9bTeVf+yKYJrx5z/Hnd6EfsGj6PTMjdsOjs28j//BAE3NqGq8zem0dNJ4MN7W3N4hfzNq4I
v04jahs35plvAtmp4EZ7JkoNWuA/PsKzGXX13SmHjQni3JcQ9/dDUrdIRMMMzz1hKrTYdwG6V7gT
F6lpAsZ8f7FozeVN9kWJkb1xeThT5hK/LMG/Ie9/PsgQRzyHAlEqTRBxcFk1T/xDYcbiUH5tO2Lf
dlh6VtGIh//HG9QJHOm+QEKhv3XEYNS51Z6WUIHhpO3+h7950Khidj3ww2WxZ4AmAYgARP+B4mR2
kiQUHX2fY0QQ+HG59bUCVlEVhFdXt9HBvU7BvgXg3Jp4HfttcraktZhIVrSLRuTMQ9Sok4F56Qkk
CgWu28zHVnTTpZCxjLqUq+Xo+juoOvXzMAiWAmURKE575WjZ08YuklZR2qGSUKkj20X60Pa3LJGY
ij6+K6tZRxXQNhDnHtKzI8LShlXeqAW8deitA68QUmNRr5jW0MaHa8zi/SQo54EseAiphZI21RSo
NY4YaAuIKz56jhhcAb8F0vGmHPAdJ3IYT+psPsI/BGM5YYt1NXu7W41tG1YwuGui/vv8ZbSuCOV4
FFka/GSF7ey7nGJX9od56fef/Ahu5vK4qxTnJhuQty6MNsMK1pqS2y3zB8Dha8bekSdiGKltDO3h
ngJmc+83V/8JhzXEHNUNE0/cthSUT29PCXZ6pI1XMdDUJ3xUA549GtoeF9sulH7Ead5fuEk64oDI
gmzubsqd1m6BX+mP/iR69C/A2Tbgr7shhhkV9iyk0Z8jrbrvJnCaJt0Rq2uCO9ojnI5q+4pQ55+5
y2wzuPmcMDluFqk5TL8DOYUBde1cc5iGhWSwTQEYfIloKymfBHsQgYLf1AgDlyKG2Lic2AqXIEf6
SP5ZhtS+tXttfF9DGX+FuTviAtdejdynJkq8zKI0xdqVgzHOo9jbxg1juupWLGUbMwrhBQJX6BIe
4xYEzfj0SmmgtJFpo7SSGCnJqQ4tPzh9j34d+iuWYma27QfY0XJPnmR58ZkBlFdIxPkmRVKJl17u
O/85if8KK+WMt72OB7Br9uRt+bBJ8044DB7X7tlvYbbchLih4/Fv0YZp+KDcwmbQhz1ZH7tShuPv
QJWaQUEjNjeYVTzO+NjcZ/j7GlNvSqQ3/lntpk56q/JOGDssTYI1ZRFPc+dI2XeIxJV834nVnb/o
mretzcRgrCOT6l2sAjnX68xctetCQ+P8Dy1/tvzBIN0tPX7ThhHrPt3pb6Ho2lZUUI2WDJ+QOSIX
rZHMZGNcigT1QjmZ5mv/JvzfWwUBbP/Pamvb7PZ1mgEdwTVWIr2PcFYKbi0neG8vvhLYi8SLboyR
xJ/1Zc1oAuwQdI0MGOUprht2EDd7zk0ZDfG8P9tbwQ1yoyTRgGdIoHDbijJMc8GmVFGGyTomxPIi
+IYCy+0ZyGjF32b7blf/MjO+prti6m4WZglh3TcKzHAYHUyuq5VJdyBs1RAG0LSf9hrA4CF70BKp
rOXsPV7mp2X8evAjt3qzUFYVjE6u/ZAU4pVVIlR9Q6dDjrhPi+0fQvVokhIovHUi1FEWAtDjjn8V
6+Y2pI3DK7p7nVIdHgs782Q2vrX3DhhhRkWyPiILJBTYtUEYOE3IjQcrq6VbAs0WVuw2Tjwl+tDn
b5DstuX6neL3e2JsRNKRndvStqRTJCm42asjqiiWazb1FRVEha7F72QulNg/ubqTiOGXOYaBiXm+
A4xocwo3yWfcgTr3dwTRfEHRt/IAf6k8MlOxVNTdv9AGU868rYhPjmYokd7+/xyhiuK6yehFS8ch
QH5xlPAWXdS6wM0d0Pxfgp2C4pIOrLbSQ+w1foYeHlXaYxdknL/3FMFA2omnkTqRtNDUQOOiNYWi
tksZeMwwvDFB0DPJjWMlvqYYsSUbI504icFb1YmAeHH7p03hzeOzd0w9pIajieQIVuQJtajnXgtC
MM53YbyERSqIWWZN4dKtJ0Ydh7goWedBUXtRI6HLx3j7/eHa/OOXok1tLbc/73ehzd1S0MNOBuLz
LKrRe7iQ/o9hT80PRDKYQ6BeYV1igkcCZr+NDxIPG5XkQkpi/Hcv7PCSzO2HnohCo16WR6tgoljO
J+US9YXoLvgJw43D1QlgV2/b8kit46aEg+hkwgpsvDzngoYiZlIO26BnywUoBisDuuKJns5kii36
suWzo5cXej32AXM9UvXQL/xoOorvg7t5xeSHtpJcSqERX5CyhifqULrPUoZVnNbKCjdPk+wiixos
+0M0iqCW16W2Bf3HvYfBk1f7cicjCTFoWX+rWDMuxWcVRUciWiXfYaUsXdq5vvl0wiS0d1YN2cws
zUeSaMQin3s0kdosVIHoIkvMUR+K/pTPz61d0Kxy39SIR4J28gqDfcdJ/HYjrztgRI+pNkgHHAI8
ArcNlvPf9mZyz8eOfAz25ipgIz048ck7CtsRvm7LKL3xtqCYgJe29NNuGy4yxVDEAjgYxL95XH5O
l2wFcNKX81O28oRvDQHJXdXF/NF/a5wvp2M3bXOIPJ8qCVselPLfJJlKPdMeDv4SbiXnfIjcnSQw
G9i/yxn8VfjcReAiowS5St4XI13S4/PzuUYIMATL2qOflEo5Xrx+YGWoPEXrJfTSJVrfn235V1uR
kdgdlF3Zqj0BWny/zBCfHTxBQo4ICQXgPYuJmpC2gtPaU2+MYWOuOY/mQWKgntxDMzoqxj3N3YEJ
wu5qFYrf0XJC2Zbi08rwUp2oogOC+ZMDVjeVBUSDjnYc6WdorW+RQcjdVmTGHfQBTev4UcpxbvVS
JOTJXQv9neNc+f0scQNLKyv3Es5O0j7ap5DHTCMScrlhY9je20yhCzT8e3g/BsgJ5w2Tkt6qicAK
8ifPsJQbCoQTOFFMx+M5u6mE2jjKhgrhMnc7JT0LG84fazoPQl0/7nLIwFBXg8+K7cPU65rxCxhK
EPPt7PdN4oC7PX0My3jtGZyZY+whtSPw3pAY8HgIL3mknCrxJR0e8RCEEDNqdb2wx2bL6nJ3+blu
x4HIYFVSHlUwnS0tAQRuxYTV7TsNhwrR14dUAVN2+KZ6skYu4YmMYhruV7Ef7w/31jJvkee/aQCz
PD6rI1PumLaRFp7es388BSOjD9Wjv4kvlwau1sBwjYtFlLI6wmcbvpR+SAJExe9ORRltOOiMbBZY
7ybDr79T4kq98bkWBs298HG29QqgPPY1px67nONW7tsdsO1tZhDwVqpdgwODsGhTmev3QVI5sm+q
mQn5J+IPkrUYYuT2279FkMCqcnSiWcg6Sxs+OvWRGIslAz8mTU5BjG78hMBbtH2ce1euEbvTgv4h
sJCQgCrwY9+LkDQ3b7od6MOcaYp3V13asUkF96kzbD+SMm6gbce652AlIOxC1eFCi95Fh2G4hFWB
YzwXdwhrHfDv5QFRt048hefA42xi1GsW21LTsBJ87hgtZu1K7a/4GH5TEH8HZrB5meA2yshEtYIV
DWNYvyqgpc79/VO2+IcDhiNhCaEIZRBMeWUh+u4JphIOsuKclhV5kOIV/i+vhiITZgkm3NPqX7vu
ZEysIhucGHZ7G80ludkgjWbGvMmUmQ+Hr42EJxpqPoW0zZThhVqbiUvJ9uX28Jhh+uA8ek8LykSp
POUnSPb2Fl8u14Fufp7HKRRIGEZS2MkiRkqW61g8fpXeDbUYmYDJMNudM14T/GP1hmLksdZz1+Zt
nTHHLEOnakjEVArJdJnYjzkuNCJ7ypWuTXrczX5vVpbCFLpAcC6fdxQ7q4PaVZNpLVU2VMacTIMH
pnsGgxk9WKE8WxyA5s6rZpGYeBF+nsPYD9kQeZxENlj8+3n2dPJIiLs7vt+y3Bw/Yq/qOoxy8MOC
TdkQ/ONtio7PH5vPAjavNXlwcK0kkYMVptBscuXpzGKA2dvLa0VBPjaZMCTGT9kT0+eyk8bcA0xA
yph+xbr0Ie088/6/FAPWOLcHLhX7MgX9Q0UDXEjCL1vip+uy/E2kr6Md632fFeZB6Lh5ol2wTb7y
x6LgiXq/iFImyx/puaYAd3soyB+QeqFkDl0pnhxWfaplY9/bxnMb5LrwvQLxazYB9fjYq7DI/yt8
UZAzLXA+yRF9R3eUh6LeK4sVRyDl9auLLJqHCUSBEpIo+/7Gk+B7KuuwdOJv7+ff2WlOM7ID+y2Z
AX8JjWtHoNf/vt1Dl0xhbXDxoRZlwD1GhFiiOiotGsfar9zt38BxykGYjqWELzbZHtSNlhmE6n39
hFik5/C9+Wdya58v0do/XD0PNIbqKIS9rZS74DYLTaPlg91yjh+DLjXDZQ5lAOx+qa7dyQ3G/LBu
YialN/7BQWOSXRpLdnRksRRZaeE4zQk1fTJki5moUVypyD7k+R2pmbXR96KM2SvbzftBQ9P4f9uZ
0SvfvFBSMTlMkAqnaMKhRgrUUihNJeRYXOj9+PVbgiAPp6Gb9mFCgn7Zy06YoLY28kT3H28E0/nL
zP7ipIjLLSrKg8Hqf9CjfvlGJhqt2az/syJfvZdNRoU3GPmbLZizV9cZomj62N2Rhsi89sx7vHWo
e0qW8U6Mkfdx/7tumF1P2DJZCIDKANVrqXOtsyLFjjqrjGhhJDMjfBn79f2U7DDNlpqRw3gvJso/
Qz8kgPYOf81qDCki0S7fiQulY4I+pXqTNISm4J8hxaocYpHSTaNis+tVb7Zmak6WdferGRFETic2
wPXW21OCtJd+0tQ5AcYIx+C7v1B7cZCBLgD7gicGUOxz2Ve1LT92VhlQ/9OccwiMrGuOcQNxHS6E
evgBSpgI7eZUcExzBR9gStP8sVPQPEpqmZWFW1xG6sogLhIsaLeyjK25cEHjfALG8Axh8GLW0hCE
LtY+1pkXMQ+/Iuv3dH1U1LkL3hk8EmkoXfYhUyduH9ZpTulv+h77Df6dPRdhAIHGxAe4ZUqWkyjU
U7UDwbwVb3krlRutNpTLSR8pP8RtNpoeZ0jX5lcrhNY9qlxPQDS56R5gFfhhjqAXMbY3dKIBqCJa
fwZ5M607VGv110Eg46oF7kzt1pTnvCV60AupGGMOQ0sq1HmoEzh7ZwxQ4ImdgEh+GcmJ6P+ecFCp
qrubfAzn/HJhbGYyeHIHmY4YBzO5ntBV/5mrZI80Qe6quPCkGGbAHZQOsm/S7STDtP/4qDe1PEJL
KoP32YXsfEzJAxxZFQMh3QzMrR3VybNXR3BiMM71CLIZfKyFU+srfBMpz1VMgAWKVQp5tBgLOtem
UTA2mFhtk5gKBjoCRZHwaU4pG37E0KQZzbVZRyRUUwMfbz251kZHUfkH5PSF2sGYDajc86mu444b
7/Bg/jcSo2UpJBEuB8CBlBipsF9mm1PNgIzClXlNKQJiLfP3q7ATsA/gyQQfi+EjCy5N65ObSXN4
ptzkUmQT+dhIIzfsel0STZ8fdjT7SAgIY3wAXi2Guk164T+0r5gfLUD6rKeFSSxNTjYppWNeYZ9b
oQ92JNdn4otdGpkDAbHjS2rQOZkvYi+yV+4tLsi3LC/L88loG06ZSJgg9crqAZbOrVoKxMn3T6Ra
oT07kXLcyA/EwC/1KlxBXe6UNBEMA1o56u9uaIMUxoW4OeymH/YZOuUYZKDlpPHOSVWNyBABGuyj
E/FR7TUb41TYswQMLmSsl1/yKEC8aPx2r2RYrF+kKUw0I4PygBivhUJy0dQxWkTsyS0qBrqZbyXz
PlRbXeMO55rNDouiAN22Kam3h5OLlwlITtnweOqH3Zm6NLm+vM17Ve7LP+YVRWffyxWH037bD4tF
be9nKGm5rfj505ls5YnRlX+T0FpVTL8/t38yEA3EzHH/MIKL1/76cPC0uvctXcidJKSKlLOvIlc7
qGdZNvo6IDzjnAMJTroQHkJGwUjx+l2Sej7/Jizo+FBnjm794Q/6qX86R15Z2Pg30CdYEJRpYH4b
i+YQcWXnwMo8cpPoVpvYp6Yequ8aeQLzcIZeLAfiyt0iuPpJfbOlTOBbK4xAlTtR6hofikX7kUi9
3f1ob/RsCVISoztzy90pfRODJSFUTMrrS5GHQ5LlitD3djuZTTE5fqXj2YvXK5QfYcn07SHH5Wf7
SxF49FD45rUSShE4tIrhiQRpccBF8To3fusNQiz/NnLYyakz2bBJcUNXS5I2N+S7QLJMGiWURJAc
5vAk11MfOhBy7cqsei3+9ulrXxB1+RJkYl0ZzDqTy8FoBJ77FlpOv5OWttKNjwplICFbOaChchy9
Hs9D+cfYa1qtHbHX/CbZCtskSH02RalKJVwI7l/02P51n2DFbzXifRSU90rZlYPOHX0Guy7NftR3
vUuMR42N2FyFy/gn1+HRqUJp+OdoOsPETUaqnJRHPDmCRneX3P/MwBocd6YEcDu/XL/0koX/nRsA
gxIncbYHSSDVnt4biWrJFio7ZGlUg2SywkqpTKnCobojG65TsAY4/0zWfO6xqFHfTXBukzVBFylE
Chu9igzC5zRPL78+8bE/pSANPPV20Cr7MymmburQ5fx3S5ulXQXNp+u7T6acZFHPeFXq1dc3aIZh
GfagSyaF02TxnwmhdkrCTwGjePdEw3sQBpm3oPtUR5jhVvx0DdT/ZJwrFnsT2Vd5u8GuqqRZXnsm
fpeXPUsXH+2c8lPPzCdvNEngxDmcCQ9vR108YV09Z9L6kRcIWo1auz5EbGv3Rh4Gfqv7P0UpVlNd
/vEYJqwC2Rg7Kvgy+RhRGS+WTCtiNUTQVmpaLxNbKCwkNQtdxLDYEKM7CSsCbPEVPxAN676+ch+s
TnqfdcBdH8iaYomjSOfsKk20FLd95Kz+Zw6c1PcUNP49kENCEn2k8t99jN+A0HhLAPbdo+hD0EWM
EAw0pKLonsHUsJFqdV/UbOHqALbNfLbWcHg737j2ltbJiCO7ljdkmG55UkChgxPa60FfvtRxRSHs
u/OkYuRBHEzitjuZiSEv8gY7caqAAleTumR/FgApZSexbBNwPPYgbRook0yHCiSp3XbSVK5CJGT/
msmiqC3//9F0m9CUi6uL9sh7GZJcCRbbB6nNCnR4casDDpDKSkfDSTSYka4Q0gohtXpA57HS3Y98
v4Hr6WpnK0sdwDiwKhcnunMBTGJkX5Iuu6aGU0uLBqNobxdnVZCmlWRWR3Vqn084zbJb0lzBsNqS
Eek2u1Z4DKV0wXq5cm+cYowwCWiZbp954tEuhVSmOcXuVGVpb0S4pt2xFY2b42VzcUKL5Hl6tAS3
xMHztsNG4lH//0JWaQgsqVblgMn3QrhfS2jq4liwVMQk6CUIuX/43FktVxkMhTHAuS+pXzp11xO8
1Qh/xnQsxlkP4AykMM4UbYRPhGQY3gLpuoP7tVl3uJeHilavX9BGVxSFwdXDGO74jsRFq2iu5hqe
nxfp3ke2YscRctOhXvlnBuErE+B8jmPeb0xfVhW+CuXh14lwZVk30DA5t2BOIbFZLTsjRAZtBKD/
t9rmcWvcnnTk7dzNlFU+JD4kuLd1P0tIBFLkTCLNROodvk+Qv11risEBI49jGCEqcmRiYOxtcdXw
DoreU5+ZyISz+ckuzJKkYOEL2WLxpzm/aQyEpQmEZD/ylUx+a1puyjqSdEMqLRfUppGS0BmRZy/U
qTTvlJZO2z1mgNlsSL7TPmUjgqlsTnqGJzfWHOyPBgV/wrLKXWHu6Fk3lW2pjy/guWek43F5Y5Is
PIwQ8wD1Py7jHxGu0yYpDur6YjuCFzHYJ0nUCtbBkB+fSdcL2IqJdYLqErtpsuapsaHiEDgw8dYQ
B3mxIz9oRjbPrWlVNfwiGFA/z6fjb7qE9GmjMx1RHbk8rbJw+iaznjbCQ7ysNB7nbWVe2wbks4Od
NRdEmyuiZkN5XibamlDGEb9KzBAZGybvZhaR14nMoxmbxZmLg3ZNqXBAodltekdJhKVLS92zQJCm
w2Moi3rNBR/U1f5+Y5CDUfE8XzH0ZKRFPvc97ydqjrGAq7ZZa33nrUj3V0QDOpBR+h59fSZUatkE
OZ/eUCAfP2eWaUxY5JF6XZ9gXkgk9WjsbVJstMWEj1NKNfBcArJBdM3+92rYs5/pQC2WeVuhu4/5
pzovms/4zuoaZOCD1O9x4Dwm3zVNzNamsEhkDeG/sGgE8u+ihC8f/mcVMazCtF9lqndmQ0GWhnz8
CDJTEoG7jBh3Wey0IKRMsQN3n5UTV0lhakjNae5WZM4+HoyzjvI5FFwFQDqsk4ECnIRu+EHN2kuZ
G3I2xauh/WnX4zq8i+pTz1Nm4O3RrziDkQaSG/vRKPXW+OphwtyB73REYCfxd8rDj7PXuz7urhqd
JpsZIhrBFAF6BHSSayIlDEDE6un5TRUFsPK1+puSmUS2/zC6dIJ5R4trT8poO6Ot4sF3oZBnlbN6
C883iQTi5wP/l/BHQWyIpZyc+alad99vRIT9N/Sn2zXX/5P2Z0UYdcstH8ceVhfjixZjIAGOD96F
lRLf09EXYDqm29cA4BWda9P9/3hWgmT9HNyAZyC0lhJPlvjy5lbieWflWBupgUTzOGqEgvVU/ZoD
8HYv49yw5eJPbujembBHLBP7PdEujc48L4gFslIFkPrvRPsJBUv5y9MWGOq54dYuxfnClXztL5jx
sUCTM1K0/Q7YHsijd3u+A8dXb0fGumgzBc4BtBOTIoHzbZiqsZpfgzIrtIjCDnorcZe8G9AjJPoo
lsyOCTiMOExxZaiUlSLfsxVmRnPeWyQX3/KrcZoXVeakQMgCTHMJg/N87MKfQ2poq5w00mV4eJRN
Q1FsbNZ8DSeDQe5pW6zJuWp7KVJiJgpeGQifpAMZKu+MbNy0nw7t75RKug/n7+lBoZdWWYMzj4vz
Buo+YE6sitn9a+AOVb+BVOpFEnA9hrZ0RbCVf7qHCx5dntDJ2gbYi9cReM8IJPPZwEvCqs8Ex+U6
90ssWgDX42spdbf24BFg3GNeyAO0WIH8hI5Q77ZvWmrDadrrnTbyDx/y8YpfYrB2k/fq8tABqXVx
OsZnrurivse8d3ab0jt8IpSoOXXZgOx5N6+cY7UlVVhTtV3akLjsVSnZKXmSLvte5qCebtRjmW38
bWAA06aBre5WpD9OV19yiu9F6oYv7isboBLf7dwFmJx4N01hzUuQ4b0pjyNTcY0wZ1AZ15qckLwk
QvmoXMqvxf7TychgHwwRXwMFsGpmUrGxb/qDXJB0BDXq77U5gm0KwnZU3RN1qNc4k7XpKLHERsJ5
Cbc7l/t/P82DmpKmPdD58nFPjwSAXBnaacu1DP7Nv7j63hqQop+8XG6JyQrxZGQWnmNSt7fo2S8R
mxQ1VuH1aSxrMqyumB7Kha8uQP9ftTQ9qo+mhkbfJTOb/pJ5M0SjZtUwR+7dv7nOEjipQjOqjL3s
W35s3qMB7s+KUTMgRU2JvnJxjHAKiT+QoGN/O6DjGWyWRIduqr7/N7ku0rhyjj423gmyy5BKNL+z
9oWq7KHHe0ckm9Xcg9Phu5MWL2PaecNX/3n9I6+NeNGXuvXPs6oKx6Np+qE87+iXkXZUwmI1RbXU
ccjX/XDcMD9shaqaoewkICPqj9+u+duz20dRhHsZmz1WIvHlNFn75VAKmyIZk1IJ5E6mtxny33Ai
SdGLtDfFlhPd1F9dDL1LGXddwhwAAvdoTvuFXStLEHqGIFHh0t130DnT3iY/H6PzcrfdK6a0mygL
fz7C4DzkdeKEbk1TZnMJSUlqSfqsGejCoJ03GOEZdPkbp/deev5SVcET43Oj66QIxz2f16TzQPN1
ugGmPFMTvwpHeC0FC+E07fx6pjolXQVdZX4/hgSwzCp8juOdxotM8I+dmObE1uzPzG8d5ji5rlj5
fuBEpVgmExV3YdmzMezqvprEgtUUgA6EAlWon5FTQrx5oH+dy4I9Qchqg7+HP+bo+kb6JuStGmHj
csNakdpRo2uI1vNDlegOfs9p0FQaYgxKKk9sGwpyq3F1cT1UMeCr4wHpbv+gDNdDHg1yOX3dkcbo
vXotEl1qubxobWYUycqU4P+ExsCOzMJ05mjzQkbBi7EURh5YE4aokFgiiNXlIQ+Y0/k8emAFE2jN
1hoqG/D96FmQOSMA4PxP+AzoAP+LtWrUQ76IvSYK/a1zVntiOsz/ZnCYVJPSnBNiqArnMBRCjibL
axhadPibzlaLvgEbVvwO14OmwDrYe6T1aYiiIkg7ynr8Wh6AG6464nYO61BpMfXw6kBD5mmfjvOi
ZL7TpyactO8icmFzJcdWeghH1Q7eIGoLDQmk5dMX0nMxmWF/yGyAl2Xuc8BjKeO1g5UwLJQQSd3J
NCOTkpdZxdwr0AEjNRumC5jDLIRSvpH2i8Ea1BIIotLnSbOGvS2uTMx4hU76WuhSiETVRkqSg//X
dz2YvDs//vuiEs9Jkruc1Ev40a6CrYTXqYFO4e8xRl2xkg2BOOInJYlRKc9A8yNEer90xNYH8tb5
cN0fG/zH0s5UPGEpbjfo6UKYXWjsiKHxFCgWwk6hKUp/GG66rqgK2Ts80Kd0X+MeDzjwgXKj3P2S
ooWdZP9u8i+P1LKPihxNq1CUXhWkaGyaJww7ET+5hSSnN7HicKj5tYvWKZPi4IU8wfj6PjN0bI+z
rE7+yyJkZLgKADDyKKhprsjfUXOeIHXt+2aoKIHCKecujbzpBTNvS6jLFzIi9Pmrv7BWlOBSriHZ
GxAWB/mf1ZnlUjwsXkxy77vnTyERFNPqgpWMGwF7EZ3x1IAS8UOleX7TPlGYS2VeWXiAdzxGPvvK
RTQAJSyP5+xMU730/4kWXHfJyv4zrQl4tozyoULq9LC10rfcmYizbGnGOs/dRyAwy4VmXw58PSEd
7m2bdLE/rnWD0i8V7u+DsLQOJKkUbW+WvvccTqhZ3Vv+0fHp5tMWYpQXn8/vfUGUsrWsMgAhRTxa
JJ3YStee6+rk9bCFm7Y7pri+DmC7vSt5X71Z2EEr8T5YY3XCBrD/ulxpkfYjIJrhwF52cw9Ej9nc
Ip9cjbY9UYk8/dwpvL96RI8o5jeu+VWE1q8ekhbM0oVeoBKmXpveRM6LU+4dB38ot6yYofBEbjOo
jrHVfGbej6DUGWa5pUAD7/mZKMPwqxtLF/P+SOxfnvXzv0k6f3Nq0xS5VbxXPx1iJkb5LJdlrBMH
aHzIaDfl3LnT9Bkpg5zqdvriKNjcPYC+Qh+yQsiyTyvGdEbDRmyduciuZ3bfRVVsMLcZcbEM+i/L
T3FwI4hcBY0U7mMx5milvNc8xXEXeA1go89WLg7qwmcsU0Bp2yhstMi6VbKEHx1MiFItaEvq+rvi
pbHfQ0ZXP3kn8E++D9ps7JW8ZJJGGy9rgaDOxB6PiZ717h74o3/m4ItJInmJEf7Isq67s+tKTLUO
jkD8Jfu4NFyT+aIOh6rQNJdPcyIVOebhSkfPDu3DvjiUgBuX+8s3zvZMzbUPOT/fYX5+V2YV4ULL
NPFqwIbgUugHU8deKvLvEpvV/dh11sFRVEdSylspCGloJnyI5U8qAyv6BHNPAABLmPxPzZyLR/Y0
CzaWZv1Myk4nhSThgy2/rPJOcOlfSuvfxgUCHcWj/8HVD9eK9VwSnL44QIhgG3Oy3EfZfAQcl7M9
OYRUGHBjZUclsrx45wU9QFX+zqw8CGTDrOWwmJ2V6UemgBNT6fJ7iCbaR4T3GMDcMbCPbaFQ4/U9
uaN2DibBRU91QoNjUB0haXZZ0FXEyYV+8IqvJTttkk3TatNlwaw3bp3i5GewBLlWD3e+yxDy7we4
bvmb6uleeTyjT/SjiDurpqSfZ3JqOGS8ywqcedmCHB49oWCdL+ysRoRKvvDokZvFq2FZg6W5cXXH
E2JNWAX6IU3Ld9911b7JZ4Ra2RC1xtnT6fRMUy9fBGbXVpMulwB9TQAYnyMr0+vkQZtdrm/2H9B+
MovczBcF3XTJkMI8onWUQi5Q622IFZ/flqUxURS6ujZdIwTLBUqCVSJ5F5QO3sScrz480/7R2uEz
tORJkccUUWxg15dTs4iD7uNq9SIv+uWrqJKCnsvTnMkibIh3Rptx/dtK1Et6xzlg0hpi+qC/iQ2i
VjMuPhx+I7X6QHcMLyOit89SqJZk3OKeFhMIkK1kk5D4CtoSJfHXFjeTQg0f/Db9keH6VYsxkOnP
BHNW4cWl3p5hH3p9ArjOVzTqqLtfSf/1qCT8E4PoK3FrRdkdNyJq0UPe25X5Ah0H4vtTngg35R+/
BYdTVu1uWTJMgwgvtAmkj8FiLgQ9X7AWcR/KKGYC
`protect end_protected
