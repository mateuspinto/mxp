XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���R����~%���ޣM����+c���W�ҤRG/ʿʀ�P���cKƪ\ס���b�+��/
<�^�����u�rG�k!:OH�4x����ȳ�"�
]��imp�˽�����w�I:l�20]�ؓ(��k��Q�$	�����������^MѶ�zk��^�λ��7�F6x��ȍ���r�s���#�\y�&�td�Ʀ����U]{&��0²ԏ:��W��K��j��pVoCq�HV�����h�s�rg�g]�=|��Ҋ��f�m�ALK!r�����Hb\ϵ�$X`������2$ؾB%��P�O{����(-�Y`�'v�7�|���+�����W6�U�dB�7�"{��׼�(��u���-��&�2t��m��SH*����K��C?��%ցf�(J��5���C��2�&��
̕2O�O�>DttC+�Pzƻ���6T9�E�{���ץU�Q�zϩ���"���15%���ͨ�Cǭ�L%@�]�Od���"u~Y��!�# u,b�3�V0&X�wݳ����|</��ǚ��}�j�M���_��c�q̛�~ma�����%�3Q�~	T:*{��8Ǿkr��T��-������pE�"��*XT͖��1	��0��@��9�H6*��a<�h2U�޲�_کN���>&Q:�hW��^��:x'm]&w��EZ�g�L��1]�g ��Psޞ��sGe��1m=%>�`�٨' ��"2+���;�XlxVHYEB     400     230�����9����wj��]0UxS�cU߉D��f�D�L�����V� :xٶܪw��Zg���l:�EQ��D����/�_v��%�,Z�'����]dG��yj�t�H���'�{���2��~�#��²�Fp�`ݳ1�y�:JX�/7@c����[��t�nU�(�/&��_(mf�S+���E	�"PlPM��3���5�.J��|؅�M_U4�]����A���<��+Y�@G�V>����8�m�8������{ig�,(<�&�9�V��Z��U�x�� s3&OH�d�ڕ�/�V�T���Od	���)��[W��1���X5�'��q����ϛ��b�cK����J�W,����*I�P_��O�J���B[o� �Y���Q1|nȴ�����Lz`12'$L�&�����n��F ��՘�v��τC��a��n�
%f�{^1��u�PT?]n2��F��4�i0�gIB����+�-�Tb�J���v͈���M)՞
�3C͜oXћ;˒��Nu�����;D+���Gؓ:�i�XlxVHYEB     400     1f04Tf�7�E��HRk��'��O}���Bȴ�PX�^=l� ��� ��^�@���N\�̔[� ����%�N�J��V�$N�,��G�Q���qJ��}�^�B�U��c���py�z~�JT%�N�ר	G�������PV|%��T��X�Chr0��=9��� 3�h�!lt���U��m�삌H���(9h��9\x-[���n߮5�#������ݍb��
F�f�w �|5C�Hx�9��]�X(�V���(^Րƅy�°�`���tV¨����YEp�ہ�V�+%�V ����p�}q]��g�&� ;=Ymt��J䡷�Gt�=�Ze!9-�,Z�R��� ���A�/�i/�֪o�����ͥ�=�c����\�R�RR4�!d`�Sr��c��r��2���L�Wa|⑰]��� �Щ��e��zsJ�>��U?}O�t)V]���~�2�ĝ�\)����jT���"{��jH�o�˅�aٯT���s~-M.�_`�mXlxVHYEB     400     1b0���� o�s�<6��~�(��iA%���j�F��x�c��:+�i[}��k�IX�m/�XE�<��)z,�߂�Aң�Dj������ �.kY�mp���)�b��`B���I��s@.����5�Q����1wۃ�s�I]Qջ�����+�"�����V��a��IJf-j%˕�K�����`�l�7����i�=p�\F�>�D���/�<�L�N��}/3�~�?.r�aV`�D�l�ڲ�;�줽+f�x���� ���t
X"�����0&EW�?�t� 	��d.����d�ΞSz5�y�$Y]A`}���[�f2��>�F�~���ʋ�0�Yx�`P[�n�p] �)���'�; =� +пH8�d��B�ez�Z� ���D9ѧ�������ޠ~�)W��-.W�pV���3�XlxVHYEB     186      b0o^�U>�R�~����	y�}��:C�$�K�����x�^������R�K�
n7@��\L�x�z9�4��+�n��b�R���u��Y�[^�&�<��4D���L�x����u���&?��)�Nv��Z��Ue-x-A��cf��D_̥h�L��X��y���/Ã+}�ns�d