XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������j2�S���֩7�� ���JS���-%�t]�6��|��X��y�,�|�ȓ�wI>�-+�.U1�m��k���uYǾeO?�����ԗo�?� ���8)b������F�Gm��2��8�%���Q���|�F�
��K�XI-�� \d8̖��C�c"�Q9�Nו^q@R�`�=�v,{�XT Ğr�n�u�PR��S������(mp��si'���F�i�Rw��~1�l-�g�;��l�EJsb�(]�%���o�.і�2��K9-z�T�-Bkw@�=ط  j�<z`�R�|=��M�fe��}�kc��Ud����ȶ����Mӑ�Á�eQ�I�����T$�0 j�����O�b2���F�J$�t��+d� �u��Pʊ�Q��G��ۜ�dbQ21���é��S�<��A"�)�h�����[B#�jo���_�P�G�%�\�G�R|ő�c����mh�*G�2��ϗN<ˎX�\G&��Եl��� l���7	->�����t�4��-��H�/�|p��6�zZ�r�AK��� ���ð��@&FW^��{=9�P[Qs+R�����y��Ȇ�aU�w\BǧO�u8)�&hF�(����/r���@8i{	�1�9�Re���!
�����R�+�\�m�GZh/�-��">�4�����N��)}���bXC6S�vЋ�mkWop���D�8�=D=�R��4`K�0�o�-���J4ˁ�@�� ݘt.w:T�n"c^��c��n�XlxVHYEB     400     1e0�"#G��T ���m����єҊ�����&pޅ&�0-��	l�)&�w���ֲ��D1���f]����'t�G�Y�~�T��a����r�'~��Ϭv���f���1	<�oa�9p�H@����O��9G��3�����"_E�TMD~ӿC�Ki,t�nQ{��-cT~/J^�'�N�
����1��+4�ct-v6
��-%O)ߋR=c����x�H]��O=N=����2��sF GǍ �/-�@9:m�?��VY6}+DTWY�:����N�oJH����9%���Q-
/�U��M5�z���&t4}�dӖ�?=�Ц��6P�(;-�
�$�@sT&k�]�b�%���=ݵ ��� e�I�'A���ǽ?b"�Vo����To3�73L���ߠ�<���z�C�D���|j�˪cv�ӣ�[�C��q��aYW�Q@+�{������rǧ�" �ML:dgXlxVHYEB     400     1f0c��
�Rˊ]G��S_�S�����_5���Y��<z�3$���x]�"T�_k}p��e@hz�$�K��,vL6�K��w���/���@ ��DJ�gWh���c<4�f���H��pE		l��t�)F�kxܡ�������P�c�-�x۬&	�����B�8HPdԉ���cY"ՅA�U/�݉�RƬ�ڀ�Ȣ=`pU����qU�rJ�8�k~m��a�tZ[|H�����=����{H�:M/���<α_"'w����L4��O[��M����u��\j}* ���K���`�[ �_������r���R���IP�0��t�_�X�ԥ˯��)R����� q����)�V6�ϔ�𠞇74��gTɚ�Jn&k�5�h�KC�<Yxό0m*���e��!�䢯!��n����=u����.��y�*�J�ڮv�b���5����x��2H��'�0�7���1DD��!L�Oz_�vkM�F�� ȋ�l�LXlxVHYEB     400     1c0���j�O��X�疯ݒ�?&�7)!f�5^��iXUR'�_�!݅�a��J`�"nu~��k~���C�(��K��l�=��m����c_
���ю�(��+dV־��f��}#78��C�Q��s�?5Hm�c�������\���5�*CP��^?���,p�Y��'EWfopG^<�|�o$���f�ȞI���ϧ`\1Bbu�pu�Y�?F?)���S���J��|��boNK��
�䃓�硃�h�i����y���1�o��W~<�F���A>�o�(���u�~�@T�c&��*�_�s�"{b6��Å�c�7h���h�J�L�S�S�p`^4���i$L�w��ʁ��PH���/�6z*p�DEA�7�N��M��ڔ}*��V���O-�{��@�nv4�< ��+�[�K,j/ulȝƵ$�Lu��F��*���VU�ȸ�XlxVHYEB     400     1d0)���a�BQ|��x.���������_�`�;u-���W_R����Ix���������� 0���	�60�!�TH��Y�g�=�i��7@�6��ڔL��r�q��N8��^Rrw���&�������x���Ku�n�ha����M�`d��G�6��f�<�s�KJ^E�ٛ$z����R���7Q�eV�I��u��U�%�7�L��&�B�� !8���^��]���,_�Ɉu[�0l�?��E�S��_!zRK��W��'^�������TYg�ӝ.,=d��l�x&o��`�vއ]3���p&r%K͈�i���u�:�<d�7#��wn��~˰gre�$�Ny�@e�|����oڡ��=�A�/�
� 9�������
bCי��SL�(��������{��C������i0��,�f��4����3A��;� �z7$O;���=v^XlxVHYEB     400     200�XHWLpu��Xdj]�
5�����+5*���H~xV�A�v�%�i�vH�H'��7�}m/;��s;� U�EO���Ly̜Õ��+����g��e��߽Z!��
�3�(��F;�t�OgaҦW�i[�Kvvd�Е�����|G_C5�����, 0��r��h���,��hj<(b�V?Jѳ�0�@l�9�l1�>�;�A���H�a��=[��\�i��Bߣ�����v!��fa����u�6��ErT�[3����2
�v�<ŏ]�yH:��2��o�|L�!���f��������@��)���P�vi�;�F1�v��6����K�� Զ|��=u&�/M�Sa�wܝH��Q�}�ҧ7�|T]��^�.N����J)(4��;8kĴYARY� �g��֮%����0�F�6�d�)O(<��M_J�2��nc\�,�֊�{�iп�������2�ġ�8�6�6)�lӨ�}�Vw��}B�;o�,[A��/)h=q����|XlxVHYEB     400     150����s 5'�/f����ͪ8��Kt��*D�V`��(SV�����ť]]���>��o���>�\�FOj�Xj�����g�l��3�aN�9�k�����
�͹�$̦Y��	�;�|��8fk��������6��=�,d�V����e-�s�=�X$�dь$�n*��k��"�FW
g��g�
i$��Ј��.TZ�'g~�'��X=%���}C�o����ګ� �1F��T�Ӻ��C}ƒ��=�����:�B�i���,���Vח��?u�?r�o��0J���l�tٝ,'~�U��e���D�����_G�9�/k�ͺ�8�0@H�>XlxVHYEB     400     170������z�~�i�duQ�>���[�k#�O7lP��d�H����FUUA{X�HH���w��P�?�9	��y�>�����#�D�S�s�ӎ��<T:1��nz+r����j�S��	��R5v��Q���lF?>�������NT+\U��H��:[�M�]u��!������)d������QŊ�z�:&7믥,J(�|G��]ZW�x\��'����^aL��wEm���e�j�Q)�Gi�L�g@F8�����B�
a��<)���U���S�[���ĩ�j>��k!�@+㾱e<Ƙ�s��%cV�b(�.����[t~�[w�9G?��0H�cT-���G��H��'~�����H(5Ub���韶��SXlxVHYEB     400     1d0���'j4�� %��A)����6Q����σ��ʕ.�;q6�U(V���e���e�;	�j	�(G_�8nmȁkE���;�Qm�`9�{�hW��1~����"l��슙`�V7w�ʶO�)a�+3ڥ
�I�Tn��~����g�|�¼S��8hU۪e�;S2X����N�x��N����z~�����#^y.gZ��FhI��9��b8?�k�p��6��`�<���AU��wb;�kx9ٞ�Ÿ�	�ҧ�h������Z�/�1��'4������$��g�Ҿ �2tY_>�$��������IY%,5����c�wq�N��,��o���g1�x*��vYnl��܋j��1×ʕM⨃�>���k��Ku=i��V�{^�xvq(v�ƐYD�R������7��N����F���\kqu�K���L��E�K�}�BA���?)�E�F�XlxVHYEB     400     190H8���'o�Ç��y��%��'Er�9���U��8}C�����\��N�]���p�K���a��E��-_�G��%-�j����q-��NW�����|�j~lUv�Gk�e���d�E	�e.��i5�Ey�J�}y��A�5�$r,Ez����FC��1B�J�w3����n�"d3���� ��s���2R��:�,��Ea��s(��Qd��⾄1�Z��
����k��n>Ye�p���=l�o �����@��×�?�2$Hk���|��}�=<Әd&*�Z������l ��q~�/ J�����;&��2����䵡;�P�#!�nTb8i�����[�kH7#>�7�&��\�QC��У�m�.4�����/�䑂��!r ��H|�W{t�^�GqlXlxVHYEB     400     190���g�{�,l��5��v����Ə8\"/c���� �3𞛇��8E��^Sk�b"����SA��NUa�;U�L���ҳu	��f�HD w4v��bK��!ۧL�v��[�WEt�ߒ��l|�ELYH��-�|��=�g)��Q��3��%Avi(���	��������К���`)����{��9�Yrh~/��ӻ���7�G<Q&�$������S0
�=�%��ƞF:}Xdf�:a��\|/�H �P'�a <�r�(�L7��U�(e�X����� 1�8XDm���ԛ�@��(N�8����?�(G�d�$�\�1��Cƈ�-A�~��<����Hi�M㊑&�V�@��쬿�ޛ�D��/ 
~�\-����Eq �u������Rj"���!XlxVHYEB     400     150/Φ|���zo8��)ݖ�������s��Dr)n����3z�*�p��-�������/\r*I	�!�d����7�� 8��X8%��Y�~I9�5������źw���<VL���3�~��P����d�ֶ\%hڤл�Z�#$b��R�$gE �9������91��g�v	L�m��3V��Y�bJ	�����ܾg�\�%�n����ܱRTL���6M�y��/<��%%Q�ȱHD���j֓�K�y��O��k��&c��̒��V��9vbV��sr?�!�4���'�����IV��� !�E2�H�F�N��9��^��XlxVHYEB     400     1506lC�������밽T�i��$GL�@��`���"�_Y������S�_�W��equ~�X�a�u����'!$�S�6��|g���������S�A�����*�O:K�n �Ň� ݆���cC#k|'���"f� Q�d=/�2Mj�#�U����A�C��Ŏ���|�h�uܟ���g�7�����Q���V�$o�A�uA9�9���D�j��eۅV��減�8�{w�:�#�J��>��y$�>����6Rn�>c��L� C��!�ΡKwC�����ޕ�#�G��,=�{�5hTA�*=@śɮ�`c+'G1��8=9��u�OXlxVHYEB     400     1c0T�+&?|�����uܯֽ?����],��X��vط�h��o��Qh�M�`ɢ�ǒ�m�e�W��[�i�٥��w�\����d�f-R���t]�y��AO�����2�b��|����Yh�D��a�f�ك����=�Ysٕ��*>+SV����oҍG���m�˯s�f���Ya|B՞�1���4~���g����bi�<�"_��Cʝ�F��J�#��/��ka�9���8�&��-�Q�����2M:
%��B�P�эa�4�m�[j��$�L�5�\6�
$�>�i����N�e�g���f�m���|�O��ߙZ �̫!㓌�0��b6<��θ�r*eˋ8��)
㈋��2���j��n�ğ5��>�v�xӇ��v����2�:�sܺ���Q��īx��u�ք6"�s��*�"]���TK���	/[XlxVHYEB     400     1c0��l�w{~ Z��B���@d�e
������5���w�W�IU�����z<�X��k�7�P��$G �ʮK	p	(5��}�i8߾|�4.T��#��6\���;9P@g�T�9h,���o!zt�R�LM������Z_/k-T�&��pc�e�h:p�)��c�m�f���2��雴j�����'1d^=eo�Y�/�#�軉����~s(�c��!X81�����=��I���[�q�1%��?�x�<�GH]���&����O$��[���c�Y��S�rfQ�:�'׽X���Q�<VIŪ	i����~Q����`'X��Fj)k�ۻ�!�?���r��8�U�V��\NS���:�)�[����#�1�y�0�?�����s�fRJ�<�aַCV� ;ؽ�gP��j�s��ԕ�_c��E \��f@�SX�K���t��X�75�K���C�ZgXlxVHYEB     400     170�
�].ߊ��4�f��X�Q2>�ra�,<�qX�m '����E����8���EL����jW0��$���t�ʪs���mR5m�A�%?�D{�5�����9�)gy�zk��X�p��X����l�
�W��!B����gW-��(���Z��-ĸ0;��Y]p�Qu�-���0?�:�b�G�k���ʩ3�a<? 3&�ZҐ`�S�{ibgF�B�;�����!�v&��E5�ba��w+#R�jp�o�����w���9�0
�S��eo;P}R����]
HL-}�WW�x&�Y��V�B��$)njL�%,��q.�pQ:B@vR�llֳ*#a�v�p#�^9���N~�c?n:A����]|���	)	(XlxVHYEB     400     200_w_��.39y�)��x��ߟ�~�_����a];���́+}/i�:>��<|d��s��j�M��������V����S>"����=ؿt[GJ Ȫ�����2�|��'�`&
��yH5R=�O��pLWa�9[��	l
(2�e6����s��:�r�u{�Q��J�H�~&4��w�Z"jᒙ�C�P�[itH���ܖ�H��Am�,Ӽ���e�P0C+�j��l� ,tGGF+��ui�F�_���/�z������#RਘX�c��-�W4�&m��EvǴ�A�1�e�	q��'�v�H�{�R*t���	���7���|�u����92���U��aӈ��P��Ww�\�Z!�����s?�	�� D��j�Wďl��3���͋ $�����r���u�2 ҿoL��������R�7��jiQ���s5&�m/����������^�vw��8�B�0w�RZ�t ����%�(��-���'��-��OXqIiPַ��J4B��WXlxVHYEB     400     210�B�(��Y�)�,7�,�)	�J��5%=e��?��;��G� �:%5��Y7c��l
gAC��k�êW�v  ����D�2(�s�M~;�!�$g�yb1q(��2�uDà����#\b�"���! ��9��_��V�M�rJԣ�R����4���O���o�n��=�&�!�ճ���n�e@�\JA�8�XA���c�'\; T�f��u�R�Ub��r�Gr+���#��G2
&�r��Tj��U�TI3���C*#��Oֲ��_Q͍<]#������"������&��W��㠁�+�3�
���Rg
\z�'x�FG�/$�WiQ�Mp�S�<JG�T�Pw�0��u}������T�a�mj`���C�F4�e�k_��3v�R0�����̔.ļ��V�g�OS���M
�����M2�x�s}jT>TEZ���*6 'sܭZv�M?7�m�=3��A��O��C��V`M�3�qT�AGL9z:������]J�[��d���֩N#��n����XlxVHYEB     400     1c0�KMt�e7{F�W@M?�X ��[Nh�p�1v��_��dx��R��/����<%�iE�I� L�tf���@���\�? l?�����^	�ğC����ќ��x�e�{1#�A;��H�m\�T*�o�|J�Ozz���8p~F����Z���(P���˓�,�]�K����ߔ/��H��.��j�'(�Ѭsd���H�alZe�Q�)�J�&��ߧӓ-�V�ޞ�:6�_!�'� �g۲z>-�
�&���D�<��*�i_0x���9>rܻ݁�!�ͦ��C7��#�>���}u�Z��J��(���l���4E��Ͻ)b��~0��g��e�Dx/JG����XƷ�Z]E^rr��¼V�j����_Ķ�{7�w���3q
��j3鯴hj$���;QL�H�_.l�-���mY����.,ټ<e����5�:���e�FXlxVHYEB     400     160���ܽRZW8K�Ž��ܢ9�h��Ki�������]bt�,����v�E�%��j�CsZN��x�߼�6X�^�n�r����Ѭ�"���'5�S9�g�We�%"E� ��a�Oőr�S�2����?���GGz�\D�3���}�HK�(��4z�:0������ϸ�$�P�zݟ}���H���ѧ��&1���d�Oϙj)�y�Z�>���(�r�Sd1�JIRoPٗ�]�L�̸dD�^cK����ڋN�Q�����=u�P*"��z{��&��|<t.
|�� n��4z~mI�o,��m7��nT����B>V{!Hėd8|@iMNB⒳v�lr�	�XlxVHYEB     400     120�����f2�2���;n��Z.�cݡ"��-@�b���a�(9�-3�9Ff��V���HO+G����>��U�\NmWf]e>-�*i��BK�CoEO��&��Wv��ϬFyrg��aL�/V7��3�`={O��0@��~8��S�[C����D��kS����.���|[Y��Ӑ;U�11���y�Z��������Y���C-�_ޒj�Qn����8����<i�X�B��=8Ԩ��
��$�7Z�jZ�bŚ4�G�L-���iXlxVHYEB     400     160<�o�$���q@�����vk,�fΩ�)^�Hˏe�.��JZ%�Tg�F*��_��<��􈼉��I6&�K�۫k�<>��O�T#gZ��Pt;�[T~t�
�1�L�_�����>i�D^��Z������@��͵���"Je[������a�L�xo�op��[�T�r�Zrz���] �<��4��1�O/7Π��� �.��`xLN�pg�$�޷Z1e"�܍=����꿃*��xt��#ڗw}��]`+Z�5�o����^~뒪���(tC /��ǐ����r΀��~�]������$��d?�ogz�i|���������ҵ�[�ö(ׂV��E"
y�Rp��kXlxVHYEB     400     160�Q"��{&b��,��H�����;����6�ZW'l9~e����,�7��?�j��J��5g����d^Z
�����!& ګUvQ�� p-J��N�/ ke���9��"�i&�r�2�r��FH��1�:c�c0@̽����V�`�`bC�+��J~������_�#�e&yR��iDA� �չ��W`0mf	����7��&g�?+g��{�FQ��:��y�9nb�3c���
���i�ǥk�9ULf$�G�����=5�P�zߴ�4Vƾg]�~�gX}{���]F�6~�Nlcο���>D[e#����䷷��j�R/��^j���B|�V���XlxVHYEB     400     200�bT�G6�����0��~��
S��]����2>P����Cw�[#�.�sfq��"{?H��vi #E��%�+*PV�&9�K�I�HȮ:~�Y����0��Ħ�b�x)_Ҡ���7iD�ߦKI��nU�4&i�"x�J�x{�Nc���lF�b�?n'�1YB�F���uI��fVr��_#�7Wf�e��]�Ӎ<�o"nlaZT����j�B+���T��p�N�Xc��/O�	���v�!`�S&vU����{�$������ ��߀MƉ�\�E�A蘔�Zߥ��|���-�o ��}��p����a�ʖ����:l"g�q�@0j͐�$!���¼��UͿ��/��7,t$�@�56����]TN�0-*�IŊ�y���b��7���ϐ���R0ABr�~�l>��oW�q-�oZa�7��,�,���vyV)	M�J��ݵ���A�<��F� G�h��|L����c�OB`&�T����hM.���9�̭}���sd�扛XlxVHYEB     400     1d0-����T��.�����O06E-bt���rY���-_Ȭ�?��h珑Sw:s ΅Q�DC���=�q���kw������9�k�V�d����*v���ٻ��@�^:f�:]���w|�E�m`�'����u���Uga�Ƭ��Wx�cr��bՍT�r`�$!	󤙼Q��ӵ����jřx�V����m�܊
8F���2�����FA������^��\V\���V�R�2Y#	����hwX�c��������/2�:�8������
�����N����2�-�e62Ŀ�x�?@Yg��6%H>�7���l݃�X������F�B6�-��6����y7�$�n���JbK���e�����I�_ �dvf��x�y¹k�5��Myt���AR�;����B���pb��;^�-����(�Q6{p���,��y$�XlxVHYEB     400     1c0/+L�<�D����uE�F�����o��M�Y^k�h�Չ���%^1d��"���zv��@�=~)�7��XDc��$�zZ��z�5j9�˅�x*����@����c n�����"�d@M/l����c�����Xct��{��|s ��A-;
vÚf�1{���6=�#���}V��f�rD��C~���VK��b�e��]TȔk�z�I_ǩ篚���:��t��}��|E�O�s!kTȆj����"Q�������V�ǲ��/�@��Ɍ�ů�;M*�7����o&������g"��:��n�������&��!+���[��3���a;g�m\�;'�c�8D"��t��ِjҝfDa/ߢ@�rx��_M,�U�6�+֔�Sq��� �~9
)z���~�H1bW�p�N]�=e)�ߨ�cP��J9'=mޣ��j XlxVHYEB      42      50�	��y+}�_M[3���%��2	$y�B�~��U����/��ߠ1��G!k"'�C�Eǜ:0*Xоu�4j3��{Lw��