`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7104)
`protect data_block
dq65nxKCFOeAWg0ybCC52Z5ThLrWiLHRTyzdMZ8tqKxxtciQcg2RmaLmShY6+O115Ej7IMQxCxOt
gqyzbpuvdXwRFn0yUlKYyTbBkOSCwiFrKXPEj7cHAfTxj+Ly/k/x+2EMlb+Tsy2LlG64VjQyvp30
AvUQ/k2vlsuTnGZAwsEw+aZ0ITfsyFw9YAb8A8LXBrn5WWXh7slFb2Zs9O8mwdUPM/oyGShdW90B
O5hrxUfYu2Adxv5E2nZxym0AFlYFYJzdK/O7nwMdZppb3Ae2lqWRKBczmmmqjoz5UqjWtoKw/ROf
+PyrQN2eYI6HFfLXvjDIEsQA3m4PEzNX2xKepwku+rWnDpgE0sCDAs5vIVTuMc+ZPuj2RsivRXoR
GaR9e/CMR6fwGg6Ypu12ZPDvT3cONoBZGR0lVMudHLrpb3emj6HfRQGOnkrPMO7gXaT57mNTZCU7
bCq+p7UZKhnD5pAHibiXVJ3iAFutClQHphYSzUA0PnSxzHJQ851p+xFO8e7Rk9fD0wOtB9ZFyPXd
2545oiDHMB3ClrV5Imbk5iQc7ZghL6rXvJy2SGAAF0FArmen+REN1gyog7KjoUqIljpn0Aa6lCOu
c9SyxXkoyhfjhBD6YWYbaLzEm9eZ4XfLTqSHiDkI0djKQi0l4E+9TN8W3x8UJSPggl6YjCgitQMm
sZ1FHNIlS5XTJj6GSVY8DXP38h4yLceKq/8P3C8I7Vjx3m2w728aqa7WmN4KDedylzOnGjUzNzGy
lRH6DiTlHKc5cnuiEmee/kXjlw8zgHCd8SH+hsdPA+UlHlaeb0blrVq+hmWkdicTj0Hf7UdH1ZoA
m6e6qRXLTl+t6csM4V9DXgztOQ8d3Qiy+xEF4L1EJ+ZuSoIZPxTCThCLW+dgnrx47sJpLb7/HdZo
z5t92ulWn6gl7Xru42pnzChAjLamPDMv5XEW0KY3R5Atqz0mW+Z2RRJNwHhJFJfKGs3rydOWdT68
Rbu8oXdP9jvsNQXwlBy/jZBs6XckacEejnXnIY7XGvbwMuwm044jfUSirp3jErXW3GlB3HVJiRbI
t08tAuGDqw1DDXQLpy7zQLOxp9/bRYdvRNjQHYxB5Z8OYV0XJ6AivJKrfLGG6xTPTCau5jcfmQhU
PKbwqhMjoy9oN7weebDcY2KovaKM9hIFdj6ETZV21f9N9FUXBFRzyARoRibFczc+5raQKaNfWQ0y
aZqcqbCNxryrFkK/+5lCUnPaR4XfM8ZDizQcBqDKdYUJ857LvG+wJtfFLAfRZwWHO+UGAkFEveP9
YbKpEbyA+CJJVNsIf6D0XW/Bhmb5D0gfLZzr/Il7EPzgvPdlLE9l1S34vpp0h5nbEF7Z2UKcdBmN
GWp/4pSCfai3egEIhIAIxsEUzPpdEaBLpP6Rf9pwAzkG60GII9KDTH1Xi8eJVVXaVagwySTi/8YV
bqPbQWtf91+F+xUm+ssKuIEfEMMvFHC/w1qzK4eav1cYNmNdNK7DHrLfwSDx1oR3GqB2px52lRXA
h2HDHH8MgmrB2dGBFcnuSYXvMBB8p613V2Op7yOqYqYeOZwaY2p70q1b0whiwoeO7yc/ESI+8ecc
Ta8oi4opiZdu6POS38yXpMtnDwH9hxHTNRs0ZltHSIRXvN1Qsg8xyRUgx72+DDdyqsITM+Q70s9a
FDbuxPs3AuOLG0ZoZNCuQEv4/mbPClnMr2CBM5Z611OAfP4NgcecnRsxiEXsZi8LxRGCaT5b3d0P
aoXLrcpqOXPoecAn1tiK2eXvJh24z6wZlUDMilJJsw2ilLg29RGtWRRCi5qo/NcNZNGP04zCCEEe
Jax1NSKQWDBC4kJ699kkx+JPiNNWzJA5ae1wuUkV1VIbhlV2znzI6B4EnjIEgIoJ7C4wd9NbpJt7
pYuB5xnNsbHdKhrVdJP3aY6tfk3d+PeXq+Q95UblDUHDVVNSawp9pfEAK9HtMbhXQmWE/JsPfitB
1CB26AjLpwXf4ScXB0FpCyi2yFuTF77Ls7IQOK1gtXwgqf6+XD40eZNV0L2hYpgrsH1C4WLZU9QV
IWHmsNeiv1uuEcu/Uyb8m5Itz8SXYj9HYHFOUR7ZK3qn2GYUq7qblIpxV5ypYdCm/6f3oqLhQDB/
Dj0fW7fOsylBgLXZ88V4gRk/Xe1ZKSa3k09wuLwOmuVfbRmL+ESohfSApWSfQtMEiZ5xdLkm2Lhg
1Rgs18demhDWxS8C1/PGCUrWHUOq5/BJKAJUMucNZG0GJ2WP82zW3qDvzEsFbFQplWZZ1Wm/+tiQ
ocwapCjm7mqW13Sz9vfr9k43IkzkUZknr6supaHrKHXtZYN+3BnGOSpOKGvcZRnM7wgrYIGw6jfq
BVUjRhs/02bsForWL0y3TptKMVq+GIolzvKrwy3sdoKPvgMAUmWUTHgexzOCiYoP/LG26fxMyNAa
icZNZEdaSVa2hiWtGuRAuNnRNpkhB6ftmgcn3DfxU2/ngfxCIKYI+dhBzs9aPQTNl3Ov1RUZCNnW
PEyj4zNyq9934qdZQp4bZ/hykCb6DSfrrAD9G0j1SuinvJ7NJlu62bF00xb8t8u0GXAJsuuFMsqO
ytnuS8rpNiiPWORgRNVYP/wmu6OJjmNATlFQahHA3KMmdVeNkjYlrJyQsBaSotZxv9qQSmydj3K1
mg7oTT6yoWWODd+3Hr8v3cHluFrbCdojWzFP2L5ADQu6nIovj7XWcvIxBP8qs6J850L7gakfcP5+
NIXthyhZzG5hcTBjkdeBsnVRptoa6hCrfs0kZ14OnIOLldJ9xGePI9UHIyhySlZRqkcZUE2BQCB1
xfcUIfEL3R2driw06GP16cGoH5rt2n6U6PTwhBim2uhqLbgQctiB0vIDhKaVeVDtuaDClQdHLpCX
lQMSjOPHwVM83LERREGwiAsh8K2iTnZQ1kP9mEbwzw5pQYFxfCDWenq01k2BOo7qjnP9mCOverVR
ZKE398bdGnYa236rMV/2siTbYajgvAlFwj4wZOKJqW3GqhOEDLUJf/Cs5qMoNXkw3BSZPAA0n2Mh
apWiLW/qpXS1oJKnWPQWYQguma3s6DXfiOpZBkvQHM98GZO3MEVSe6zRMDpSp6rXkK85qquRVmDp
EKzwv1WWnbP5ArZj3klRlerP5gC4ZqmyGjbPVkN3KRLb3SF2a0IxNIewzT6RFLhITqh8VEZ8yAvF
DK9sA++Hs2Jew77B1ZAhZXpc/GDvoe/j24Q03uDJDYcybFfJSFX/PvKnM7fK8/5opNPPHBiVEHuk
/6iQxNRkbJHpuG+BPCwdYpez2vx8an8tjQzQ2rmvvtKm6ndJWCcjQP041dx09/ASoJt9XPqpTn3Z
Ee2jNvd2d4QCALoXtzcsgj0PnLwTu3bqYtBH0uGe3WdwBFp7DSkIlR6ZN2c/5JWlZiQEAb77ZRtS
AdAqWas6XJnpOr+wVOlsX4pDg6qKaJddA0f0A1loFQMx8JzbW2nK4cVhddmkUH0B6jGfCzo4d2XW
0PGc4zOr5HxV0ga5IBbCV5+gxAgF3ELf5D84Xbhu9kXkOEKcBIv5MGNxmdgcE4Dj3PqIeztCDlim
xOa9te6Srv2kyVMjTFP7w7ZxiWehB1u8OkrZvmMNZ6Itw/1D8qYR3lOeREZAoh52YcKdOPpnPj4q
VnrK32g0Xa+3ZrQneJXmbjWKR83unZClzDVaU/ZPeDagBITKQBXilvE7LvFmFgyJ8QEHfoAsXP8j
lTIKgC2sX+o0AvG63A1n0cnq/Ti+ZaoyXFE3nHOtPIeoZacCh3roOiAsZJ1FnwP3vV0xMmmy3V7U
htkMrORsPrwADaxrv6sXQKcfsOqoxCJUOeeUe/rZjqE9vbbtrwIYXN22Eb8/6tVJAiFdhlyCJ/GE
jJyfGGzqIIMHWgPaYWczJDhX+aoPoj6v14iO6IwdvcO1UfP0n2oOhhNyWBvERN3aFoB4vEmh7wX1
tfTXUzqv+Fry4MoK5XEQfQzuwmI4qlXyDHKsniChn9O7zqE+JHWgo8EWsnN1QXoygSeIMPgYTPcw
9bzSvbN5WxuMn/Jf1fS7FHt1zRrkzuoFLxNI2wvBuO0CoANeL0VibHBEBQePqGrUXX5OMrNiJvAn
CZEqYIuGbHDSWz27QFZ/K9YW8Jiowmj1bujtt/q0fw+Jm1ezDx/pX3chpP32bEfZaHuFyxnxjApB
9CCzWn80J+SHkbh8x9jAq7z5jamAjtL5+Jr8bEFKZ517+cRhYM9GJGHMoCntUkBSHMPd6Sk+SCfN
u4jbH7GKD0r1+sN7wa3DuldW5kyBByF+cqA3RATKpYbS+T2fqxB7kp69de3xI71Z64EzwiduPs20
j948nVkdJsoSyL/s6RnIyUWZ5mJPFPwH4Bd6CIWWw+cQ6T8PS6qLWNsKfeaQsYMOl8H7TYGWuT7H
1Z4hb8s4csyc6e+QR1/VYPyISZKCh4sCKRlbvmtnFMgkkAF7BdWgmrRYnFEmT4ksAyJUsMcj1vAL
vqRLtEHia1UeHep9T+6xXCOhF7EBd10CQ/WOWlTwk1UotkAXoMPuWw15Qyu3ZfYoj7CfHEwq9J2m
pFpO7XsoEZkKxbw0IGi/Fq3/ToLOlST3xCnIDSqG5NCIUxOOwftmnKshECtkHvVekECSqm65h4eJ
gCsPLloZtxiI9rQshMjLGWWOmZr+eY96tlHE+WQhyD3ssPTr4ukG2Tov+LpRYStIEFYWP1TIBOER
qEuQGGGcRQ1VX+AAF+5LWiSynNAQfp/N6bojNYdAjA/c3NyTFst2tNlZz/SoJkIc4gkJcjNFlTdf
wU11LPVxZCIX/SbfmkDmTs2wU7hr8ifmnAKt2Fy3jZ9UFZqIV8tBKbAaGe/WLX18krIdYZ13kqtU
yNbtTUp+48lFdDw9HBjd217kziO9XpSLmgHag1UDZhnzR1XdJx9jGm3emgznam5rx2SoVAWuEEhi
vg3FhVNgebGhqHV37A/m5fIjapYvXmXsCY+u0vrGJWBOFJipZzi9hAaSF6a1/cI0vvUkT8QgJhSq
6t13Ro0nRuDgdn0nTMMIIMHpzHM2tL6LlL1Dat1Sd5SNsnc03kAp58LnuB5qkfQ4mfqZekm+eaSc
jOOlx/xCRjwT9OZGwtCENGycHeURsnetmXqYh9noOUloXad7ovVI/R/7vbCZOiIEZjdTaa9TSjkT
EKhYuuK0fXle/0VjRT7DufeFKni0EXwitAvlninRUdHuCt1MiMVjH6aLsVidhPG24mCzp1M9VY/Z
X0x/HoFRGwlpVzi5lMTSFyg2yt1BIZQDGYkD7ZoE403wPf3RTKZqqX/ODUwPOYkBksW6pEQQ+AiX
o1QLT6yKivmhHDo5jO8ICsJXn25gx+fgOL0zLVAwc/fR5N3uJYrsIdegph6kxCi0V7w35VmasKrc
Fdp8a3nbE5m4llYC/SS1H8mZ2VBP9me1fPMe4H6fzvf3IKqxM0klaC9x9SU7EGD0pISkQ3V2A5ly
VYgh4Zum8m2Z9OkokSb2PitSWb2QYrAjcFPhJUAga9ykRs6tyCrYk87d8QVR1+rsTGwRf4DuGDEk
KVCDYwAkEEW08qwsMq8U6EJXMh9G5eRBLww5BC7UDmSFkpfOhzta8VRZieYB/n88xu4tYCfk7rpn
R/fgMYNo3iLOzpax/GBRk4yxW6Cm4gFWBSLS7xlTFhNhRhKsSvMBATdac/oEOuAe6GPCVhdITyqi
i2yo2xMKrohuqxBVwDgH+tbSvLaO0Pd1nWlxS7RHwKRX4gt2IonSOd5OkqRAPfOr2q6i2CnX8i+D
u7pj6iZKIFvqjvCJ8NhFZ0MAGofHXkbGUzglsMKT3RklzFZH6UaL3I9S4TbvcaVBlEyX+QPqYuZv
HmdVfbbUamZkOtAHbDSeFQUgegzLVE1Ouf7ZjOum59ubpCzCizeKah15arimCbwkYiAM1zsiK+FO
bdL3Lj49EzEWBI8W358eFX8kHBk5U6FVRI00nZmssFqgh4oCGxdIHJN6vN230nejgcef3A4z6S8C
bko0wfvRHpjBydAiFdiFmI9DI0t/IL92ERNFkVbsIEn6YKZdTwiiZM75QTUkdOm81OlaW3j5sThh
8c3+PeHXRMCeFdWOLHPo1v+I6wtyLjdHvmJV8cU2ri1fO9D0nkd+rYJ2im0E/IQVTD8W0iYO7mY2
1G4XBqsWDLUoGmdLAEvS9NAxQs7KSkpLP22ja1ojhNAzekEozjC0P/iboYpaz3qcUgiEGruFIXxd
2G4p0InW+PCz+GAKLNzpX4KSftSeXOqHj6qIvIPXioenb8AbsSuaw39eOtTEdbdtTMk+cNSb66Gb
42s+UdiLVpkDHVLO2y0RJXrtm12cMbXxV/FXvjSs2/A+cWhXZtdoMPdG04Jzer4mAVDT1zJWOYhX
1B9SRLVqAOnj/NJghIdhEhjNbFyKQBWEqliP3OaYcyeuCFf+TKe9/j0boXnkLEUNfu6w7m9u6VoX
ptwMF+ll3A9w5GZyw7PbmVzBC1/a4BQwiT//4TjeF0vt6EddwpRd2bTa971NG6OUz+2WobupT63H
DPHLWnZWSCasZF1WVIZRDjrUTpcE3d0o3UsI8tKsmw/AqvMg7rH1mHoUx5FUSOylKn46411asCGI
zqq6K7vYzv6wI96YmDuk/+YArNbFkzGOBOBkFqcAtYIV8rBSemd0Mwbspsa/vxo9pkywgce1zxXq
RqUCN2MByfjBS9pD7OAjRAf9H8DTxorvqeNVsX2RUIdkCdlB3DJBGHKCOrFtTWS3A/homp+HEdh0
8wO8EzfPwi+npB4RDlE6dxtULJoL1H3TSqrEEFS4J3CETSA9PdFKCMYcKDgjey4Q0sO2aaSWfgl3
Mhy/MmQX4z6GNCNrQZTB5a5IpDX21HMaaEh4nhxQyWqkFL29qWz5OGaLdY6f8EPsKge5+IaLk4AD
IlxKiJF2Z7xmk/nAGHl13Kz5PDiiiwSVusjos+KBSTCQmOKTVkcWDWew1hm7mqItWJwFmrK6NglJ
60h4yzNlQCUWCLXYrkY/a7GhurHpZTJZBblcbb4yn/EdsrAqiBzbHP/K9tfnaSCuL8dcwqaCE6Jy
BiTdrU4c2DAeQRmzBsjUKdvoNbLHmf/T9tXmAuTXZ5rJYo+5zrcGfSz+M0LXrV2bZ//hsi5n6hcD
8wzndH29aXRtF9jDkmxWDjSPinZ3NNJkJ1vSFHZv5/A/J5KbcbFBtsO1NI7LrdhvRuW0SiJR6+nS
aXau0zkZHjOPjhxN6AEmXCcUdbQWBhavkdofgUcHBFPkVKSaoAoItYkmY5kIXNmmc/xcKh+1XmQO
xp2mDorcCy0PN3KlcrUbRDaAMlw5bDLqK3khqnnnTeORv3IsUA0HW+4uiy5n0iYiq7PWyp4MCsZ1
Bf0GxUqipZx3J177fcJFMMmRK46ug5rYkARwaRZaHWnPtlzxYRMl2PQkFlMN1ZwzpO0Sgh8MzTqW
uWbfYxIytnhw9ElY5139qHjGoj1YeVut2vv2JbG7dGUsTDgafz+xCt4sGw14uhkmIo5uvauHHnGc
39+mahfJsIGXFzI92bgoVjA7eQjPUL9tJ2lJ8cHubtIt61Fms6hjDpSfIpDS/YmbQ+XToEQLDm4D
R05KFq9vUcTCdQJS3wzalvZAfq9KXY8YXLMxwg5pRwaXpT3bzFXzS3ITxxczRO2jWk5tE+DFrTZR
0YGP40xucGJlNgubZZg8mErvY/weps3BJdv18KkNhFK1XZrnGeM++EMOI86+HnAOkVWx4m8u4JCC
PGSBFahPnZdLk0gK40/iQ4rk4lmm2qoc2wtZi1GG9rGHXHJQa5ZxM9+s04tJLqYjCgz+tzbVsFWE
4Ei+DZXKdxWhQAegtdHtGw8d/0gkqSoePAnJW4Ro7OV25mi9XDo10/s0T9knHuVGrGabWATq9d6J
UvY3QklxUU8FV5hhfmQwAB7ekKyxewwHOdv32NiexMXeaXIVCUlCQLRPt2YPF1zfNQnI1x/GAYKz
Gh1kiZ3ivgcbZ1vD+pjgcsC1OT11pWXBM9ZYppTbNFb6N2W9Ync4IXzImv7IRUjvTzT9CRekGRxb
FgJ+lb+Pw1ERc2e2F/qMSfIMHVGlnNhXyQwH9BjlL4JJbtFjL0eiHetUp/OJ0ljV9YMeV1v1yYK/
xkE77riE8WIoVvVcsTqvYmaMepi/W0BbNtF1G62aZP0Z+g+/+SVh3RmwmVBXYlCfiU1z1WbN4nUJ
seB1gTotmd5nuj8woYOjwquGvysa9rUj436mBkdZFlUjfnCcdX2YNiAYkJPW5LW+Z3qaDDBhSdi1
Y6tIhmmYyUzFH8DZtRK0b2XnGvvH2v0sHsq3M8EDnZfgx2oTEB00DsZBgIHMMXE4g2/z3OpKv4WV
/MCgRM+V7vhWn8Lo97Qc/+A1nkoIrVyjc8GfGJVeMaPRoEfWKukEbFgjerxsnQ9n55W0vQu1PAWY
I1Lq9+Id7wRUfME3KvzcjUK42q0+HheDahlif/O0YxaBRMM8eSfNfzgErk/Mwrz2++VPZrS03i+A
2vmScQLSKNRemEczIBaP3OtOU4PaxORslALc936APQwKMeI13ApYT6mY55SrMDzxo4S7JWNzfMwg
EDdKHKsxDk9KI003Tk58eL0WR7Ka4W8gZC91/ZzHQm45SKkWiGlxLbNGqXITOTJjL+HnhJTfjDAh
WvG3n0M5a/MkIiUC7bMANTaiKRsg1puv13lfE5L6jhHPQYhvt4c/PmC+HahIIa+5WItYxZf79jBN
t05MQzdWyp7OJuUUsR2qTQRQT6OXeSjXJp4Ikq8IOt5zAFMWrC38q0mYZqrCS9gfcDr8JV9HcHK9
FC6RWMLsLzoc5+k5rMaWaduKSHvqFWiL4ICV4ojEBZZU6npw2QSdYAx8oXHQREGff4PgfMYWRoAJ
+hqXVRt62BYWSIIR3ESe53yWweLf4r+ePVyWxkiHvoAoLL92P2dK34DZvwveYrBp8i8Eawz70Czs
wLoj3HphLdHZ1DlyPAEHplqu4WWubBOciyesZZrYhIYdrek3dUswePnkyCyQb9c+fzH0izk8Hwvc
WbNWjgYpexvSY/whrFeSS+5G/NBZ7xnuI2NUFlKL2ROIviEP8MCqWg3//0FizRmfEnQbU0miI8ir
MK1oGy8cFFbfvmv/a23c/ciZwYitR+dH6ygXaLjb66KkTpx1IToGbP3yv5nNBqnbKJGfEpLO1gvj
N0CZcmpZ2SdKfLGpy+KM3qj7cmaisJuMSlSvlGsBtlRcW1NLfiTykkr55SAwhS25Oi3MD0B6981M
KypqG68Z+nLRlm0gpQnlVfzSc762efdMxJPVlXO5Km5Onazg2QYBPGkSr89bY8vEBL0MnKqVnC6X
6x5QtzZCTU5jDPvlPWzmqu3uZSW3z/hq2dfWqpQ+QVeTT3DiH4yHzTRdb171eVVyNKSUbAOxucjG
Wl4+jEHHRmHwzLH/AjYEsc3sUC+bX2UN+uTo55QOi4hMJ7il
`protect end_protected
