`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
GsYSijc6ZtaVgLgThVLvdgRgAaqvjDETY5Gc2I3qu7FweqRTyXimEbB5n+uDBYeICI3JeAoR20xT
kFfB+mRXSZTQC1oS1wK8pvMV+Ub+nfWmEP0yBkKT60Qh5Rck6RtKpwQSwk0t+sktin1VmqXsnb1z
rhNK9eCt/uvBzjWuezAzaMjmc2mOyq1BqMbgN71wB4wBUvfzrA2NQAjAqPhez2IZZlzksxy8EuTD
0xLMqyQ8es7EbPup4o4QhIWP78ED3ekCFAn9lDjaUX7lOIsRMup9ISyRHNlTojv3wmYpqoKw0iYg
25if/t1HcxXBlLLlO5o0Gy03gJvkCjweog0P1A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="GnofeeOOjWw8fScfan71INl/L0+3i+faRsj/I4B/O+Q="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26208)
`protect data_block
mE8JP4JSiyJndF1lgbe/WY2hhKBCbG77UPYm59jfm+c/8GYKMkJnse0CKSKIataEFdRD/ffjq3Qj
4t2w9unSUIsn3v+4VaGAIR7l+ET7et5KiS/NiWbm/840/Lqxecb2E/yoIDUJZFoy8SMWPPZeL0VH
i0Bl/YqD1QaWK3gC4DHl297T2Kiv9FsnflpXEcsH1dKjgKKQTFhx6HpzcBGWMRewaBC/dv6/wLOn
9wiSvSO/hcUmOA8FzEFm1HQECnHYPraJXEp3GlKwwx25bMAA39Ofw6aEeHGdCIdz0usBSz0sJx+e
o1qg4pyrvz6M10T5WvmVLAgjEfQwDD3RaNMMaJtX8zeuz8KTwR4aeikFhoUQ8oZiQbct5xdjS7Ex
oYwh908lYvoK6R+GXTXOESOA+ZEViN4O9s7tr8TJE05WyjsRyuCbtDo0dHS7BWaCaAEC2NGTRcOi
F6ZbwPo/poq11PHp+EWvCkpLsdqesq+Kp38FP52jsEQzPkR5sFMrJJLB24nE1fbYZdc8xZIYbnxY
jUQ4P9w05TwyuVeiaQzUnq8VtRstn9iLM9/ixXUQSQOUGglvC5e6mYGzBkSOC7rZhW1OI8xxKgW/
G/ICiqfKosJJF0c1xZtUspIV2FVDXu5zF68b2fMjSr6v5Lp0GgHuDpNPKqY+18k/QfgvVnykh/pe
rsi8diwKiK/541vWGKABj1qBnKc4gytsPITjK6vJwKYXO7z9kI0/aTpgle4+7JVhKnisQFE2dl9o
JX08E7X9y2QP5fsgJDLg07066OC599NFIoNJKtkyIcDCAQYI4eO8DgqGVPzpy3Ro+V57QbDyiKCM
uqkUpFMLOyfW4wQxzCZJmoBDJ75RAI9HO4vvjHyFL7ykHfSMPa1m3C0vN0SM9MQJbbbrq7c2+/6r
XEVdGky4j4axkrO7w+3aD/iI8hw58PUSTZ7x2OshPTzBS89UCdX0lSJgJVu7OY6VlqcNB51cBANZ
eClVAQU9t6guw79psP3sGxhpkLdwKIy2YlTzJYWXvdWS1pVnoqsQQGZ2OVZE3WV2zsEc8Zi0Cqdc
+cR2elNzyzcDojY2mrKbBIhCF9VSb01Q4Xuclbr7J7T53LhId9YB2a9dFLLmNWTTVC4f2HqAu6Tn
aSJai8o3sG30DSbwiSJuyR/2F537V3kzL51UGCXR0W8j3/LqZFsQuM608WM9peFEACMmOsd5g4wp
q6+8w5DWX7WlSbJoxV0r0fxw49zoTkcTeoI7pXRhP1D0gGfFi8QQG7mgRQ5g2vdh9hcvNZEPnYqh
7m3lVnVJYf/A06EvpgMAGm3thVV41Tm2O988gvSYiuyz68ykPZ5jrCsTQ9cE4dKhvMsOSCcGxk4R
XCzoOpNElsfguT+qnSrR8l4/vWtMUqvcKODDOb3vjFTLH+CqyBiey93lvVOkrYsL12Ql5y2A2B1F
Qnz6EOGVY3P194nAoW8emy/0py7/QTErYA86Gy4TMMZwXIuHi5+9Wme5K0iWEqyT8WUNJkuGlH/5
5gFnAH2uSrocJ1Opn5a52Mubn3HNrCg1e0KcIbHCWANbNTJhVtxYiGrl0GA2GSJ2FSTWRyvIvOvZ
pcEhnZzilA+WvbZmR8aBC0HJGJqNwi30yqR2AvSvSZ2oKlnD9SAqBwwYCGc43vGBD62vv7OWyjHv
Gi3iBWWfCs7A+tqBDSJ14Wbk24h+1I/j7aTcxkewu4VEEzuDfh8mzxgNsCRQvEJDyXOKchFYIVrI
b5N9ow88tnUirfzTeqOUOT/YEzwm932cacmwh8Yyo3oWDEUXNWUdOGptZDSXPM0+D0heMGuFUWpB
nmGZR/w0+evCEaA0FVpzWKBaBqH1I4XLdzyaI66kLWvvm3Mcpioria+WZCChbT/gKEvFUb5xEiKa
qpdA6be043pHrSOuxtH1MkPks6dH6JwhAeP6tTarwRV2nlYuu5FxKW/9zb1dS13MulSPcFuPlZls
9BFa28EeOssTGElniV2a1cfJbGytrxmWhV31s+Jya+MB1QFULuxuhVgqTEkklTsT8S7Tgdn7wFqV
37ZuAScCy4ppdqNVVtSW6UZHj0YGQmdGE2WEnUb9n+GELarxhveqpqpBRy2NbJZMAxO5u2Hou8+s
uTm1divoYnym6v/rljigPLarYDuDD1oVPS08Md7Itx0m5e2qrbYPmrR6JBV406AoJFAq5jjz0DuL
CpIgtoxUwmxeNPDCPidepk/70LIFpE0ZQAFbpllm8d8IAbu43WgHE2kVSzoBEKutVQvlG729cvfg
/1vcLKr8QKghh86/TlHFC2R4bX75uu/Gbl4qEpCwfjWWYg0Z1XUdeWCais79MDwg/MSAL4MSbpeU
ygHDK4TKoyZHqSu05xpJl7EeQYKdyZrBqqD9eJeoH0zfOxeIonWGzp4MlvTOWzsyjx8Hdgjnj4dO
d73Vby6iF84KRZlWyBIH2tJ4BJ0eXTtkRU3hIMEBIg7FmtPtJ7QLSVKU6I8ZMvDj4I952eBPsW57
N+AR9pp+qfnNhyKdJWnjvBWKQT01i5Vm+6RjhBSTB3wMBki3A0Ip2+/EUAdQgbC2dzdeaFqeT4Xp
dbLZIjfMVghokC/ECX96tMKG2O+NNgDDm+tmLA3xTJq0sSIdqeduOUbM4Qk3Fijrdn6/CO0UgbMY
xGTDkskEiMTVB8gldcAwAH60sseZHf3uJyPwg7SpxIABQtCOhqwk9vgMSy/K7I5wr8jWPJcV0ur0
wjaWu1dx+OcFmUODN5uxIjbZMPHLitKa3CqC5fXslp0r6NbdgwbZmrYF+/8lnuzLDmCtJpiyenhs
hrPxMEx7DXB0qAldZ7KjpqyK4O9f3xLnAm2gntjgINwdrsJ4ylqJrQ7nlnGe0jLfJ8N5sHfeVi7c
MpmaUdYtXGRmac0EsZD06uu2B8JEl2uN0uI1eUjLPS3v03iRplo+t7hAKPpRoTSXpIypJeGkI5si
HiQ7far48kjwXGJPnUjntiMPtj8fRZCZ7+ko5ol4iNzo/trplAaIxHb6nLvv0GI5MC+L4YQNslI3
XDOp4JT9yS0CaRoq22Alc2/fGnTpEXjzd+LX2oUOXzYXOWtJt3r7IzhroDCgUD4FCB54ic2WgU00
VWNxRQz8DWZbZxv2vKwlYF47SaMW0STDColxcWeJUBIVYpYUNmAvqNh3FRWgnoIhceyB2bHwSF5M
GdDhrE4BksDYIFk12leowSrLFQD9CODRvHPf1Hm40iwDsWReKBMRRXGd1TBAv1EY5bI84mWbknWY
O6esAHjsojUx4d0MSe9FUrqoxQswGns/36EJ5JBuljiiInZAhDJQvCnmiJMWH/N0V8wnqmRRdPic
nTjRajtKZmF7S3jQcKCdfW38/vsk8wHOrw+rVucMwbvQPPkGcyqg82tYh555ESL91M6439qDhOAV
cZuL+uMrJ8cubHbDZaF3HrpsnfMoOviRlwxnX1SUg7SkirQKV2JeQDAd7QCMSA5XOQOXlB/yrtzF
mnEegVzd1kvC1qgkD3MyfSL3vVQ4QMgYkP7cwJe6LSeT2CSozq/RThtUKbTvmCW1HC/sUoZKH8NH
ES+xYQA760Vcc+q9hRvlga1DZjpj9pSYt6VodILEUa2YqlIrTVFByrlDvM2Lf/yNko/1nLQu6h3W
S0ngE6aH52nttlOQTJJYyhKaxJv0069simCA4W/De9QbaiYHqzMEZhArLyWranCs551oKQqTP2/i
TX4qDnBwIVKaFJQTshYcnH6fBWqjWh1snXAxn4Sp8fbifbQVE4ZfgXR1vcxDENvtkEaQJD6zsyYf
hdq0gqgMHpvLOEHtrMki367kNvre3O5VNUZ4QgWgSUobhHehzicHjUXKIEGfRgMrCWW//ln8zT5v
VfXduUusQmYBaECMY0fPCVCbfLzSIFyQqB6ZQgkDTEnh8yJMW+fmIMSK8P3RFsCd73EkQ4xNwTLL
QUQ3Q1NChtYCJq3eIiK2ZOY4uvnAEKXHrTVa4OAvl/pzshjkd1ydu3PvZFtECDefXXbwG2Gu/3Kv
JLrZCr+ZzRGYmob3L/nXB3WLKSNm2nMZqecNdrbrUwJAmUVvPp6OK1Uzk1+35ofIFWxV2aWaPrDu
lwpITnoRL8hapZ+0XFv/bj4GyDwFin2dupz86xLEERu2a9KmCqNh6IqBuoYk1Iz8U8ggeriC1iZg
jiYrlHJf2pF1KWng4cL659p7Eg8iGOymE3XUHBaJTMURB+Lp5Ihe/IZeEbftH9f81iQG9+zx4cZm
eao67sy7NWZxHqKNWUcqxdMWMYRlGFnwRaZ83NV8KgZ9Cl4+duzRhOcTcFgg4DT00OC+JyU42g7o
ki7QYU0cm2qkXLCox5Je8s92LUrNN/aW07Csmi6Bqtj56Mf8ZYXN20LV3HrHwTXyN5xh9e+d4S4F
E0pLSx8Q1hS9amTzhaHKaHKg9o1VcOtcPUHLaxfJNihj86hXNPRfma2X71tud/9/LKGAw6rmV17T
pvS3c4FmJwppnvsbJXXTaz8y6ftWCTZKgF3tNz+2JchoobQ7NBw6W+KozwPBjelCL0pY4JQCo+5X
janPLC1GAfd09FtZr/0A5lHAyYnOLKoZvJOgPhqKI53GHQmDYN+TiWEha49ct35CrF0Q7R+mqb9e
hhNsA4Evo7GEalSnCxPzVzWtUmcoY9g6nDi9SFJMht5xgR6AgdKKCw2oVAIF/V9YdVgyhKKq37DK
LYw/5h9MrnTXBkppY5D99XRdkOn3qg+bJdYU93qKehZjhUSH5aoMzSZHMIjbYVrVpFoeevcxOXHy
mnqY0k8ayadfr4hMiM3MvKbP1edXZmjkXFCqUGxFPAc7WunFeqZRaHI6SRzir4wzCENGahckzRHW
vg9LYCVXB76/ws6Q18AicpEJ+G2vGhYf2BwtAcKhXS2BakmjygHhIceh1KDMlxAjon3CuRJoesH1
0GMfeREmANEpjmdV8UK/8SDly/rD8vNPPO7z4CEA1//nDh3TFFZX/1CDghjT2nMey08jVdWQmZKP
ybpojeBdEC5B+gdzqz9GJnq6ENj0TUA6u71/LvsZBVkbqndNXyRJkkmXxZIA/dMC8twiiIh4PGld
BO8aS7CPgt7ShVcMFMtxy0Z51ydMT0DpIxPBA/YpI8NIQ/OWAtlNHGf/GmYcDdcCgMuVSp12LG5B
JmF12Q9bcCoSltLXqCx/tPsypDBD4dg3V7l3NzNNO3P/1B1nvW3a8RTjpvkHasweEckNFjHVLa4m
FtFDkMhmbRGzIUo6b3Nd+eWqH306YsXfP05GsdEKELcK7AnSoMf3Q7AKaFIwWLzbTRJiQbM0Yoey
k8rHIlUQjUUoQFYA1shzwM0y7LGOJTi5kupRmutCuj45m0CHPXSnqZEIJhChYScnHoSAAclSmhfa
Z3Vq6s7gQjtjwdZ6xQnGEpU4tvv9rWsMqgQpGZN9ujYzV6EJf6gZ3hAIT6V0BTSXBsHxlGR3yqO1
g8dKirTuyQEIp1cJxKtkrqV3fvLLpAkCWpP6p3S7CwTWny4Dxqbo1+bIGTxyDkZEeMhwUeGouNri
UIJBYQLnUD5JKShxM8mU7JJsQtDVnrNLLN29MOcURTF2MplrQG+ONbPXUA0AxD77e9wdH686kbEy
ZjkHANGxB8aoBpiLP5RPAQWqwz4P7zMMOILiKOnDnxoxCOX8NZfxhw4PQAw850J0G7/jOTUGFVsh
in0NIVPhCF25hNB9q+uGW9c26fpcopQKTQsuYwzdeONMj8JOiYe+STEMvQsqQXl08dcBfZbrbs72
MMZB6a9N59qzaoPjoNtByFAaotUi0bLDk+R0lp17V2YTbzmcJcPd86hMirou6YUwTLqfRheKVtqE
l9E3jQ3kDcP8LAYVx7HnuZ/gMbmWUh2avI2kWKJ7tOtMBReRQdU6WwtyfjwepmTwTSHSpVpFlID3
G9zQVNS1UjgkTAbAhkmDlNXrcTOGc34GtaT4Ou5MBmHm+U6Ci2JlpR4hWHJ0Au5dwgEIFuoiIexz
CM6Qrgy8hzwqchDjErBUWLurgN3sTJ+a1rH3rZo6zVkHU+hy9lL1EwX72CYI+pwH5C0CZPcb+OTO
B2meYwY1kPR3omQQPuZGwX+lZ3ZfTUjJk6dLNDSqnEy6AKhXSsV9iQoFTTxuN25tuhxq2j7YREak
9Mf6tP5qgH74rO8EnjimVUwEvxyVI/lHmbMhDVfwHdyP4lNQay/uVOhdnV5B0RjPwF4WCmvdRqpV
B13J66MDEUg5VJ2Wbbzq7f3PgLhvaUhn8nR/NWK0rsmNADcQ1Seh/10HctWdrF1v5WDfcwWItQvy
I3kje5pl2ypkUlVfeTG6tpsMwDeg9ePuLEU1CCHnz/K+5kk0x8igpnY17cq1Th7tDbrjCv/VjT0S
j8G2wP2n5tamET1H/yMuM8mVI/CMaqQtesiLe8MzdcbP0KflzpJr7sDGKXMZckCJ3WmSzjZ/eBet
lvwqfYRJnbPt/MckcLf2ghA59vUvjimzCnVP27GmyQhvrx+tHV1NGxdrijWcJ7Vg61nm9HhaggLS
vIzeNlwM8mr0aD29EaJKqKoivMVVprEATTM3YLU3boZjSxCltzh2KMavzn0sT+Yc9AfPpK9Z7Q4m
HGej2heuDx6SFHLFwScJXDVd7Kn9rlwhivJTDXVug7kpRAlsYVRX5Bb8s0MrCDjoKtbE0Pzo4PuU
NI9WL/guEgf7dklrnesS4SOHVV+YXLsjYTQxCJtBup+09aORAnJCyuJCvFIgBm/V1PI0GwiAHV0W
kHhdfRrHERw/y/m3XG1G3tPPhNcAtMYStCikLqkWg97w3wp0pFAH/kF5nuTCcxhXMicAOsK5SlhA
u7h10OAa37jsNgUxemaeSwKCvqWzxfQUlDi08/SZVGUmqev23e8l7YDQHWrChtFVUVg3553biZNH
lYa95OIkKUXzk6/HGdpjdkIN/KW9pBBN5aItfpzV2PpVsrxynTLwx0JXsPI+kcnwwb3q6MpjdHcc
M982aN62rjLaVqZ0PhCNwQ13EavbPcgBpwY6X8j3JSzBre6fdIHj0HOMZboTtZMuwbzLDBzJPX4V
Km4nED54rDEdG5uWWrbzmky2xB3wXAj15o4jZ+tFxFkxCMZJnAjk8NDa5n+fSq51Xc/2QHh3tMb2
q3ZGM9yFDq+a90Hl3mb9bIF15M4YwY1/treB0ohcWW4KrsyQ4wVAVS+Vk/bcIIoOSqO10rLws1v0
/4Bhd3BxTgw8a8sbPIToChryMCy8IbUd4RCt9KhkItA34MJsMkvHeNXYzsDpajfTz2nJ/JxDE19s
gGxPBTIl6yfmSGuBgQGEYQqShiYBeA3pOGd3GwUWLZVpEkIsE7vu2v5gZZfOlKk79g0skZFIv9Ng
feE02tj1uSYGUL0B1YVoKjUhofyqqpIS21Vgq4TxOGtVdsK49WGeNo2KYL23UL2rbpNr8dIaT7qn
iPWyIpQLFLgTjen20BgP+v3j7WDamAhsOVRyG3nc7kB09QEy1CJvgO5B74zai+xOq9DcEhTyGZzD
kV4/OBlO0S0fe050q1fhbiI3YzXVn+dCxjriQ5cVN0KMzbw+Rs2Wfa9Pp0uFhuBBpb+oRmlOLXYI
XlDNM2lUS7ntOCmZWvr8sXvXnX9IW4FHt09v0gPKUCfpPMyiCy7uEXCuGIK2iV4u33tajBqiBt4w
XmL6QE9petqW/Jb6PQByub7SCCpcRznvBuIeITHjR8jw1ZWjFsP+4v4sYaUnlh3s4gceMOHxz9B7
AwtbIEP1Rzd6rzKEDmWXW5EHUYxVAEPuYjNw1ID05uqeJhT9GNu/RJFJ6nOnfH2NrdHFAPLXb9lJ
KUurL3+IjJYYtl/f7Z7t3mDiibAn3/K34d5qHnuQsazRjjvVV0NtdlL05BwgK4QaRGS1O5KUSbRh
opa88iaaJrDn1HfNihvI4afopFUwiPazcwijGRANyXTK0h9qssPR3IVI/q8KE9OejR5S2kJ3+yFP
0NL3ZrxGvwSHZXW+ATAa5hKfXKI0+/JLLSRDWVsgt8YUMLiBnYifPeOEy1klUlDdrbGn+oNuPBg/
Soh1mt9afrr5shZWoogZ7c9e3RrkK7s9aGFs8O6RdHlFa67awv4uYNy81FkdUje6PAqoG521EGNR
UK1oYd5VVovRviSvyHlCo29iotS+kQ9NDizsCgWNbTgVH4BfSKtsiXHjQXGOmgQAZV8Da6LkM4bx
8sWa6CEzMxaFQFH5j5dY++Ph/hGPZWekOm16RWm1NkKYTfoCCOWyzS6wonEVbuA7pGJ4R0atjtRd
OxmlfCwGmCFm41XbvEWZY9fT4Xck3r/tMBNivNcPPMv9DSjfQY4pRhVWq29QmrSAFKcWrTkGT02S
QXYw43h6RyrDKdK51NQ8zLfVpOr++zXMuVzO92W6Esx50LdiPghwn/l4koTHVg0YbePWwAJhc9it
O4x4946eEeE3cKNKU6o/CGX+sIIO/19m15ifq+F3hNSq/w4W5NS9CWAXsOURXdHQ4n/HiDi4u9Qr
A3V+en/OkNpfP9VdHxiUUGd2wigzSMVeJSoUF5QFl1L18d9cZhNjsRTnNSZZXGAojsW06QOpHQ6W
D9qqVSdbbFIbDBbepTjm/d7QJQzvoJa+CcXUSnM9UBeauehH9iyxkg0rul5t+NDivQ5lR4RMHndN
cZofYAseB9pPE3+6UbvXWXG0Dq308VNzAd3si/w9nVPfJGeUBIYrSI0qwq0+J85GiTEsFTr78CFW
ilqqh0f8ElUXgVgQ3IumRgVAFIcsvI6sf792RhuGd9B4JBWOaEbbZcm1CgtTK7af5X+U+TTooije
/95tlqQd5VjtG/LT7x6WRGcYj/akXvFFzlxFR3oK3LQCYy1Z5958v0dI0JQemxAOHYn6wHSt4HiI
HdZGaDeVHG1UsNUdCiDUaqzg0D473BHLDEusgMaMYfuyvutS/f4pmAGP7N16QrmBrsEkhwsH6cDX
HE+ah56Vg9XyaQxhneBqya5ozRni78BnZrC4tIhrxA/4AZoLUEFz3hIsXcQG6Q3KHNXXwO0gfLp8
HTzOJEvqsL3gPSl2WkuXNRHeElJ1U+kLvHRVufSSaDZnOfkTMTMKS5RyOpPBJPsHhYz0uBo2OEPF
im5oJsVvw7WFLhjEEPplMmIwMWQMZaz840apRWoPVrRjiFkIDeNqZCIidJ4Uc4k9wPvpeFhiObpQ
afN6jfq0Wfy6NgWYEDfl0aiQAXFrXjIutCYuu0V6VehB7qB3Aq7oDeH3KMxoXsaxiNE/xeYaCXwt
5IMwkc9gFf9aHNrxm4SlnWPuKhqSe/Y7KhCtO09T72oqO82iociI7p1EAQAB45+D0Z83WfQANQWx
dDcBFeArRJs/9O5Q1okPe9cQWx5aNuSPuaiZbu+2cjqYAEpjnza49IG90pr1/Ma2YWockbUxHVnc
JA/f7ZqHxJY+7oL6FisMkoTV6OFkD3YpQ1scZxx7ZnWZuvHMzzIEK5XIEG6VTkFMB1K1NdsRUNfW
BmetjtpSAyygOGQlKugbo+OoZk9Q2kvEfZL1/BDAzro3YfhMlScCa5hL8soea9af2QTCIjjKghdY
2Y9BIWf4o049hxS1ZP3yIId/HLRsbIbyAkriYO3scMKd4qrWGlFqliKIxBYZA4EVx2MigFyzvmUo
WHxI/zh2RR14u8ucYTX8Hoks89tihJT1i4tThgnpDG18YUqJCAYyt8KZ+SICxHqH/tA+4G9+B0VL
2RUYSKkxrHs6QV6tLFbV/Yq2LZ28uDoJRYZDqgEIa85orfldcSB9UNscYJQlL4PAzJ+cR0yQzHds
zcpkf2qVJdC5OBFVDhhfSKVRitkyEMZehBYSIKyBkGGoPuJWMr1IdGAEGqswOOK4VscJUr0SSap1
BTd3NfoSv+rJnEwOXuO70c60e4IOc29jarNP7YmaMKMrSj4G7bRiK5oBYltVHGYDflymsTYZLE64
CHMbU+YV3whCHjdgXM/2jqclrvai2/PaFpXOM5su+Lyb/D+2gpCvbqkBEkdbPOns6x/OKyktxiZA
IYQinpprqohWuwIhN55hP4i0XxkB0/PJ7+nfAM8frHLkuMwOmUc25t0iItgMVaEybminaxouCUxX
NqZyHta/qJX4iDFayVoT9rdOFKM0r9GRuxUzVbqv/vABBCo16dKp2QNFeoGajlOxi+t027YCKqKv
ilrLH1Fde3LRcBNNCftA9pMFhsnDJf4I35VkfRehHNTd3U+qN6/m2bd9Y4IhdkAP0m64PM1vf8ne
XxQMtFAEeY9cJn9qp5Z/DzK4YvueO3OhwVp2EdC9ELpQplrkfSTVQoCmVUJS2ggAOtfjFld3SFgk
hpheT5HPYGAeLFgkHlSKj4bL09H31rbQ7nCB42uruJoiKuW+BGSRNrtjKz/BUeE3hP0QfwwPxjoC
61oiTr3Onc1iNaKbrefCj0ktU9sEtb6zxWS5B2wzTyF3R3IZhVMDFGhn0nY3NZm1WUGzMPcxd1lE
9oaN7uE55+ADxPHk3e4pQaUcE9EJ1F0Az4/kgj1tVaRGajZPPa4b1in9FQYMpK8Lxt0X4sEJMKU9
6C1+rBVWPXhJJYIUMQCIsJQOkZuusFiOmJm97aAX1Zr95avX2phAtlvFQc7JnJrjzcEGhZZ4H1WK
uAWKuzq4loQ0SpL8WIb8bmGTPsBASEf7QVJOexQSLBTLiZPvLswH7E3Yx7mV/uZGmkJF6TqEXYLZ
EU3Fl8bNb5vLc6LNrAKPm7GN+09BGwmSUgDb1oETV6tUj+63lKbCiVQBzUwVM1N6FCah4Obr8jOm
v7Rq3T9XwJQRIN5lF70nAsxdL70xSVczvcjJBRLYDEFfx8a4NaT5kFQnT+f5+872AP8jtQZCqZyU
xB/60lRPhmSHwt1M0k7j2JQvrJR2jbw3WQ35vkTUVOVBXn2XP0elnlSTe7fiIeskO9IdTLXe66O6
FyMbtcQQUZ0BS6Fyi+UvfJO/9ZWQGMS45BvNhHqop3NFfXPPenJTRyrttDi6WGbvUQDw3h5m5EpI
jVNZ/VDoNJ2ixGnuZsa7I3u88q0MFaZa/R3h9z9wLhR8ut4RWV6DSJB4KUsBKr51jMJMTPEyXjam
foRJc7gzYMhu7EWk36Nn+0oX6Oy16o0ByRxseJ6O5XFE3QMj2EjL60TFNmO3jvTzMkXzqItL5i+q
Pq3gd+C0wwWMYWdGVWoE+gFAYr4RX5TMl6lAJL5WAY0XOnV+jpGzjevcYOx1Y0vLKUr58UI/Ru4b
rDmjI5R41cthF7N4oBLIQEGQmAzK4IVSxSqd/u7ll0pChjNzlrEPzEZYX1hLKwAxfcHJBBrHxZZy
nZuFAJ3KC1bw+tofILP8ZkgI8XTfHzECid3Akiy7AYtJUDaWrMVOy7U2ZZ7l4iHbUNSeZJbmgZhQ
yKoNiTxLFioalAGjsRUOX7O+Xgp1V4nUZarvx79nnSKmUbHRe/T5GfS9S6Qkj84uJKLWb5yMdQPt
jWf5zfQZWAObnWIhxOpo+9gUAcLmCN9N3p9DZk9yeO+cm/X/PbRNSu2QRRIaK2h+vDoidljoBh+K
5ALeC3+71doYyLB+GZmQ6urSyFYbxJmyXoNqNFaDk6Poh1NBl6vMG5tw3GrGxCRpcGII7ZEJkhpp
O1c0U1cPVdq5ZFvM+bzHZXdW0Nnr/buSia3tav7fY4drM6f2AexhWBSHOKT+AaUiFoxEEySt1wH5
sRgdVbQIkVyaYfNVXSkNtflR0dgR7r6lQefmfYQ52CfOeQ869gc9FKXfsVI2H+z6vjLqVFgjXFAD
2CyeK5pbFVIVEzjaXZ9KsYgkh484enlufjhGxsw87uYoMlcFHMWR9J8a9hOw9XhBMuhB1bCyPfhw
19fZtjEsdHQjAnZXmdwMSyajH81OT3QeESo1eC/DDGKP7hwtstNmQO6xn1O4DF56+HfUHLhgOLWk
3wUx9hqMTIxM3EDDZP7G3a7Owd6hRXovkqPS5A+1iy1kP8DceZd3aPPZzMolpxtJBl8LDiCzIbXJ
NQSpwpPJ+zWaNQKadSWANkaVBr8fIcZPFiWWBzyQNjIjPhHPH1FomKHivsCTns2T/0az1ol1CuYF
tayC1OmuG0w/ng83SU9XhqFf15oamh+htVn4QNTinhg0Wx3HiRu4GHSoyf2X2GHro3Fldbrw8pHa
054FgMBIAPU6PftIAJQsNYgjHhWCloQ/upTt5W98aPyxOvR1EldaZmhTraMNtTrtPYzqygt7sP/E
TR0pEVnvtleLzDDpkfw1F2LcsmBgeHaZD4RHl1ZgJ0s/yll6dRtxrFJ10AqprHaXDKZcVkbR4c1g
xrAKymFwXfLJXIJdHhaUtjPUtRAkO74fYACOxgQmInKDbbUb7C4HLRYKIvBr4jtOoKSQO41pVCsL
ysXiY2UkFBpB7RmyeA5I06iaX+gjxhaNpx8IMGjoMyWsse2pxDC8x/DAygVEf4ktiT+4yjQnYHfB
WJgmMuy6YwmjS7GQnaVHLXtmtM5m+VneFrIIyOIBRNhFw3b9gvmF1PRV0qfYlSaFj7RXmAlXw1t+
KQvKSl/SR/CoSRk+8aLqpUsChy59DTXJekuzEvT3IT8ib5+X4QJ5mpfh47bRZ5gunNyJ4TlLSnzn
y51IEjYjeScLdnjk1hH71qf3A1iRfOWUpVLR8g70h8O5hvNELoT0qNyGBemlB1YQBXakVsmcmdOg
Jaw/VGI0rlrT301QtQ8CaQ9Mmrr8jVfXD/Khr9FtTYL4SpRCxkYnsKmRXPXw4DN5Q3KuZX7XRryP
IH0jl7dm+ZbT6t0yYDNdpEJpLjxpu9RaR2eWOC3PNHoV2gkEf9/HjYjgd/ZicPV2C9bRDQKLae62
s0Ze5qIcKQHaOMBu869uvtORWzqhEX04aYhLuHbYc3bnq48QcViUCrv5D+i2htcSuXBshiUqkvnz
+dUfGQckjT7m/Px5sIS4bWy/OMeirW9UV+1MxY2cY9q0NkcJ5oy0HzLbNoav605uq54pJn7xJylr
Xl74khBvUpWT9I2NDDNDbDIpfEDyLhtRbBfiXOEvhLJ6zf/X983bUMhBOTlxcpLhNJ6bdpaElFQ7
+Q1Lad7wOPDmrUy3fVAlMiPpvV+UHbOBcRPl82H0ysyaA3iFL68oXE4xsdqtebhxrriJ5qj5QTEW
AwJuVBe6fWHfL6lu7VyIcW0vXVgM92jwkyWxDMjG7KHkJiCEj348An+SeTLDg+ZMFOC3G3diuGO/
IxLmMcj7P+nju9cvZCW1NI+fxSfTfa7w5dm2Se/805wMSlBm8UkDn3W4talm3uznWjRnEsJDrfH3
JdySxWozdA+NDrBJRDaZ0j7zh2wp4xHmoZxEZc7l3dh3t0rU+GfyMLlW8nVBXIq4FsOcqJFwfpK1
ngGUUpKqjfC2jYmnbv0R3AGX9nrC+fQ67/NdgOdjU25NVL1PJUmfgHrXxdHZKYz986el2D98Kx5q
G8a0rdL2y1aN+teL43+btDdlPkl1Lc+oKOmRjTiQo7lUhnZg91gKGC/f2gZk2Qcr24c4gp/Y8tld
rT7/R3lUcFCK9pkz2O8BEzQTiCuIQnh3CSaI1bdPTSkmAN0U5voFxywbaXKwF5OIwdiDk9bQUZh3
YVCqVz0SwvVEmDoTuD9aTan7107v8o3QYBvPes67P5PQxPtYUkDrKuC71hfHTh4O9D/WtCp5AYVN
0rp/oFoKCFmw61esschK6bBItayVqQgo2qvwUm6tTQLehojwUR/IJm0AHF47/1OAZ+Cj7cvLUC9b
r2+E74nLSvBHbaJDvrIWpFw+2JqlkI3tUjZTnHlYvIt8nRUrylr9fvQ3/vVBqBj4UDTvDgo7AM2a
Bxg6hzyI+bi+zhod1oL3sIfLnqYWzInwf4meClLZkz1CKs7RGTpYNB0vtyf+yC394JLgaN8XgozB
9aGiNzbfRrnaiGzqNtNSwh3hRiy+ega50Kjrze7SZ3mvVcCFEdl8mWPON+AI/HDqL2/PHftQ1gxS
q8o5bTN6LbWZ1BYt1yQoheEJpIuW8CzQ2b1QYxvSDV4qUVrUxNzvMSvwUu0u617tXkV0pKAaPpAP
gRrzA2GiBUbUsGw5AbdoTxIcati4Z+6bJD1d8PG2tu7cqbwWimGkeioC9Lf9MbeFWQeaskMfdQJn
ADeZyWE1cEb2L/HG9Qctgnm5Jp6AH2Fi5+Q5i6Z+jD1kRmq8Dt3D3Xg6KJG0rKKJyfz9sriIicaS
GrcwjjntJF6CG73RiUsvRET+idtMBkIHWj5QXOHX2CH/1aPkkro9Bp70cd/YvNUMokousN90K+hU
N8cEKnGUS+oI5J7TrZczIQBow5SN2dlMoDOyN8RX5Zduj8lD1khqHui0NB7EHg1UYIWD5o4730DO
FBWKNDtbpmeu3kZ88pdvQwZI/xm+dHWiwRzsR2ZioJAjrfOSeuGoF1DeZtxDIsZR4sYQ5czLlw7V
GlXurKICMgUcULVQBdWdd58GpdadsusBOvaKXvLr8rnt/PLUxB3YCABQyDOlW4YDpvg6ZQfOAkYT
mIgGjvcMBGAHw/GSSLmhQZ9uwFExSHX9XisectjOYNhEeCpK1tTuhei7CXcTcI8f5DJNezUM5Vf+
odvmu2jYRspG/n5FTo+ZVSiVvlgOS/DXBQNXwYgrx1xc8hrh/nP6ceT4GirkFRzwVu1EWdJkLkJh
teRXLyZ2Thj4+79MA8NFNE1KEprDE1nZH/YqNpfKhcl3F5cYrk8yXRTT9RkLH3llxIvAIt/4eE1v
JEDUIP6phpU19z5XLoF56nT4UxgCefIU2RbFnd3PTDfQkKwTslwaJdq8jvrxMprQxnXU9gvV5ohr
i2Cx3/2naQq/2MSO4XzPSlCE9BVWnbR9EG9WgQsFGVi2hHUgHwlt+S/hkNLOZ+oi6olXAPr5mAlo
nBHcLvRz4zh13zc5Clg4xHPkdogndJBb5pnLd1SDinvvMfpxnmZmzDoB0vYQUpBGu++5H+NE+uCU
bSfRD2Mq2ASijxWJ7xhqWR0sunoyGitb/7uzGFucHhkHQ34Irm6epoiYebYCUJlHKsipO6XVW718
YL/7EI05rGPPyjY6Sm5bPXkqCPcRSJmmpOiZG2xfJObb/k2GBGq63n+fEpujYt5PZL+1W8QsJUxW
vXN7drAeXLvD8QFcLRj6zseq4pb6Lf4SK7/sjy7pjWgTu1Pr/xtR0c5y2m1d5B6ocU3V/S0f4VC/
BpULuXIybA8VfyQFa5Uf7Chm5IulT8Ek5GdIM58kPFhilgOIdMyQpYFbUkfnCN+xU1wyzs228Ts7
Us8cyL1ArOmfKQvvyRlRJ4eio/WZ13MktfuiiVRIQPjt1Ff7fnnegWuGCbHtFlp0BiuhW0L7ees3
+tvBj0eAy3//mBQCkaPyy1Wcn0ghvd7c+V+bxKJ9Pi+3H916m5NIHHnv1uOFfEtjLv1aBZrma8xy
WnSkG61rrH1JR1/qqRJP578RLh5HWLqgCY3ACNTfv7bBSpUy2KwH+QW/pdJ+kc3hk3WkvYgMfAMV
ll5B5IYCWMwTBlaWzpFsGHUfzgWe1FyFn0pCBGAYCWFz0Brcdgryu+/lBTp+PvbOBQSDNY9sjV5X
NVsU6YtP4p4afYWFXaZHL+1dptKp+68Ywi8ZaROrKkcCYbrdzo41vgOvECVAk/yp0p/185zTZkwz
fnbVabT1iHr5+IZwV1es3wdgeFNRzXx/sZs3+P2v5NkBfyzKb32Wkp3XRMkJhtcpufpgz2YBCQSq
zZqlGOX6UN3sO7ZbHBFIZpK+IcpK9IbYpJNuII7umX4fyrYZCp6GA23teexismwhkYhR63AkasbJ
hDK9qaDL6Zuk465Xt4H8ekieaMm+1GxLs+3IMHc2iTa7A0Fb9BTPo9IE7lW0ay6e1rjTAoVBdqui
/jB9GgtmS9rAMz6boXQuRkLKIuhTnU3Av1KQ6PcsSahax152Xo/5kzBApWvuEd0QpllPjo9KQCU2
C+MGQWmAS6dHALojaL0YyLRy5gpXjF6wy19bdOhmkeAVR8xgLsYuqc/ktr9uxWWX9ABaC+yhePeP
1+14j2nFQC7eMKJ/OIy3qrJzY/zwWCirhmozwmJtJtGFrcWtq8TaIpUjfw3Kdm7Kn/oxjHBAALT8
VwA269Zajr7wIW0l6xrzgbiE7sniWeTq4ga11uBNs7Y5W26NU5gljoi+Sw+/kr0K3hFxDZdOWHMW
ATdgYDRws9MGH2ynl+wnCrsrD6ifM5zqT4+7JLPgZsz6iACSJmElUIdAZ6NXqHiuqiTpR5LZ2YXw
q6MGz0DIBHCluE/31f/JJpblh6mntR3eayL+9WgMvS6EETeo6su7RJ3sw3aZegznaowJseQNZ9hf
TeLTLAGt7qhxknV53sstKqhMrBWBif26y192sx5IX/jPTH4WKI92SSAov/waExdu9jZFpbf4jHGA
gLZtuZ2xi9M+b6+RUCBSki3uFaAwxk87RKjsUXpQuo8sBmasUQS1NDrlM/wMNJ+ybEpSVc2LpV0W
qYhX2Uw//FgblUTP50Q95uSSyqRz4pJVegUAXhb+vqfgaWcxtTzIUxn5VQ6c84jOG5U5F7E8ZW6Z
PhggZ5Y8wBKw2jOeIPjxpjai4+ib5ZzSw481TIMhRg+jMGhtxKpHSlNA2bkEved6b90/+W0lld8K
TM/Jk5woArWWanPUKDulFs+sm8Ukp0qVlQA1qNQ2JMo4p50HkHCacsJRmb+cdpd56UE7dQoaycmG
OjCN0U6ufccGU72AA9Uuo5+fF7St3DyvTPoxgfY4y6/h95wtjeR70dUY0SuBDEH7KZHiBTMn43eS
2aGBZhZQEPz43KhSfDN0P2fg+BUeCnUPpibUwWPx3bKI2IWeYuyvrcCmWRujjqtuvGTumpt5fTZ6
jXuRu9+mgvQYFdv7MLodFHaPfhy4OZIKnIQl6aQ+c3PL+AUmfd29w4tyj/DxySHhwntBhW4VTOfO
PDITf4Vj0E7S0n+wapEkzQlaNAKjOZzRNo6wByuTi5XixucZMZLTa9HQpPN50dTWxMcJynBJcuRu
oVKDhOYxY+yzHiKSAJYl54c6d6ki2kfPg/8xcWpKrHFIOQ78ctrsQdrtkzrnibc9LGF23P780LJu
tOoqV+0OY+KqzNqu+wFHCKj+UMZWQCoDVgCXhmyiH0NkdHIA69H8u8exNyMn9rUB2L4jsqHMVHV6
Pz0twp9+AbEcsvHrMq0l65WYIAND7QTbiTivtNY7lOzngJy4cUZOm4ydlHrJqHMSfKT0Z9Qa5XRk
G9vWNTfzHJ50rFucmHSytV5sokkAF7FaOKNL8yQQYk/c7IQXvLpEm1E52jViKSmkxKoQl6v0c+SD
Ar1rf1PffVXlXLqsng0dpCjUDb8klj7+5ErRhOmHPSrvHhiOHNbg38TSQoQiNnHqAZTOgF5YrFzY
Atr+e7bv58SXip1sHCEdDdIou5izQ5jOK4kTzg9XF2cvidECrWtX16pEARVcYR/pwRvXHekSKhE+
ukiRef7R2DNAHl37Dfx4/nMSpC7PFlMWE6vo80WSwwfzw4y4i3vsTXzFHp1oZlmC8N3GU8EKHSbV
qjyLNij2xTTfAA5aoTGWLHrmaxxbvhvFFH1xE1sV0xanI7L/uszD6larXmWmeEdxzVAaDugSiMDX
g8An8+AaqgA/Yv5JRat0ZicbmLwOttbq9/5XxunBmqdAg2ErjrKgqp8A3OyniYLL9Iw+xFyjojyj
IcWCwtWyg0kKK179bud9uxCffg/6RG+Nol5JkFbK7m16Eq0Tmb4THKs6FrkjrJi9PB+klyY7U2vJ
Qw7/kOvAiEXJuLVLOgqzFzzboTtRT4eU0W0s8Xani6MwzyNXISdEJgAFBBUceiGuPetrij63m5h/
2J1gtsvdpqs2Xl1PBkLv82/CHOmr/ezrBrlujGADOC0JiTh0LfR65knWUTeAMNll3bDF7p6YRbUV
MvcDtCkmVA3UtAacxYBkMybT+3ILYC0rrL5pyXyOAHLznTo+llcgVKR4i/iPtJ+j6rv2r4xHpBCM
hNfhXB1i0fPSrd4Qi270aD95N75nThWZLkHdy9cSWBiBvSLBJZ4J4R7hN6MSlxo79DITjhIrBErQ
wAg01GN9zRRrBgwBk5UFHqZcPgBOheBsO42VAs3owp9csEMQF0GaOxL7k3/cq68cDyBNQVX/z/jW
rAGOo99kijm0kihe6WZ4+vUMgjfRxKof/bGRIsS7CItH6br3wK4DR++tKstBD1+WGuacy25ysT6X
7Yn1OvPjtF2HSmkvWJw4yL6L/aqUHubHGAQyQxSIY5zyoNMTxyPQbFeezzr2ddnj/p6yCuqdXDY9
IlBPAmfPuKkju648EANGQ9Xf++YmClvsM+A86eJe6Vny2PQtmjnqMxzrTxYziKwHtmdzG+SToNSJ
QV9Wuc7qKjmW7r/+LJrprvXXddvY/Jnetko/X57LXVQFKevV3BbsQT/jmMZiCzGoTShp/d0FWobZ
rT5jf7ZE8iq5oSDqWo/ps3jaaIw98zSeQ1GQ2XTJeUscm3kw1VvpOJ6j+NG8zsR57V0Yi6wiC/em
mY0CdGzz1rkNUippiYjFk0vrEjAqfR1cOEwPCWjjRk+1iIP5qpUOwfQ+KDRFS0QpBqj7tnCKc9Ed
h3tTogmNMyprbtJs+d/KfZF2z0BfA8kZt8D5OOZRMglM6TaBBbEUfsnJIMKzOIH+G03SZkLfDpE+
rAFckaIUqNrpkAo7/VzdBSsTLtfk7LwxETemzGtlEmQ/E3MUXFyXjZ3KQqO6q0u2mMO2riqwEiH8
pFHH6P5erqTEohPfYmqpaQZ/shFX5Zk+LY6J08kNIua1vqPmnjZxTBf5O1fSMYDzkkzISdOEHo9O
tzjhH1niWdbC6i30oHNzzIGh7eTnxHSjbWJpnXEKyjuF+GA4LmvAIwi9ZbO6SKCpEuiB3bbfvPb1
HwdZ+96AtLctjmPpjM/m7kAK8tNsxjjoN4usJZqFLtzt6SzjCqefCYxcL7DAAQY1VK1lJvX9Saey
rXi2M5x7ko4NUHK5EMTc5HglkQcaPCI6JRMnTd1JAc4pjVIBAmhr4d2VLA9XsvI4uonG8bb71Jba
y5Akmf/FDSw9nGkRb99fgk0xWSbSK8UhD85X6zRh73oeCgqyRi/bN+nLus5wDB7Dk0fCVCGQ6k3l
/K1OIcwXPnccy4vfT8u6c0lj/pIO+TVmdDl5jNFV9qQP87v4tON/zxKhk6cPS7YZ57F/J77JZb0+
lZlcDuyeDffriHwAEPrQqj/Fw+vUaJvB98/mYqK9IOdAY8of36Y372GLRJiV9h90apKkZjO6gfeP
QsNU6icRqlUTfJWzWWyR1zUKobRqUfZpzdxsmFrrtwmVRdQ/IfpBQ+x0327272+EiD2ky+MGI275
RYD6W6Fk36L8cuwTx83NtNkrq0w13tnQ75nzHSIWhjNu9u8bIVIMCdbBrkqzlgawsejM+Imtxnoy
1rZaXPW4pPbYUCFyCEOfOGHUQkPYtPFIVGu6D+NwdW+XC8T83P8IWmGhKkygQnrvZd3ANSiODGGk
HSVKOKvx1vMkBi5FOb1CbFTVOKETbfeLTzNAVbPkZnppLFQyh+ht8Wyt7aCXOk35EARdzzbGiJbE
UyU0tUZu0jHqje5mS9XVPkqQ4T93wAp1bpKFl5LDGrZIusDYkoLe+er5bMQXVOcu/JcK8avKCTOD
LZ9/m/EINzf+njYKn28LNAt4XFqQuXufh0o6nm1k1EmlnkhXwrRs364lvwhOZDmYIpgzAaItDQeN
aQpBHpT0Gtbt23HtZGvgoEJcvDh2cBNGkkmoaXxJkPhqt65Z106SEstbZ2i+JQaInScMB1Z+zf2P
/5sTYCfXmnkb2vM9DWqxenw/PFX1QwqYuktmlbzYy3qAvjgP3P9hvX1+60xb+mjODwDf2rfVU41A
OWBFhuqu1AJ+zKaulhKwZTO3jfbItFGvXXhqHRPgRpkvK9ylKQ7H9QVj2kRsoGBd3hA5wid5jaJt
yQGoEy9Cznqk69kgueEmcc8HUaO00/X3whOxagAJE/Ngj5P4pyrlyeCaGhw8gMIpFnb8EXMTQqw7
l2BqUnNL0Uz+NVlUuXkwsCiSM8dhNDfrHGGTgzCrSgtX+ygiqsFa9qRO7LhDLLEvs0jP+6aohQ6K
I2D/RFWXOlrR7FFfqVCW3oDeagkEEEd1x6pJoG7CYDsiCX/3kiI7lEZk/WKurN8vzoCukb70wILN
/Kns9GP7B7hDQvDH4q+EQ2lt+RyjY2R2RLSEeNMZiHH2bT3mwwT1kkvGdeAkXGXsHTkSsfrDckmv
iDh1kL//MQZUmM8bSUdTuIAOeXBIrZ6LFbJ39qhSQhbVKxfmeDnxJIEaqzHcJQSQ7qrNhrW7QmU3
xTd0RoL55YKNbt2HGOzk7mGukxbjPTpJ0kOrwrDwFFOaVVKoiT543ZzPAYKvD+XKcp2WGzEh95uf
0fW79IszUnT/59NgmIFzruG+hGD1SrVi6UzxUi8TzGblVFe2RnFZeHBK4l7/xo0pmjdJtRN0oiwM
FPzkvDMME3g49l7zbuYw5DZ2zjm3IqmcVnMyR9acaOV+p2k+k3GUSzgYPWPpaA4mrcG9dMP/hcAf
0adahbMJ2+yIpw0mM7oxmJG5ikGWBliqYZ3qDdPGKJ8ua9dYd7pGL6RLkdNqY9GJ12dJsMnRE1P3
ibRJ+N/aRM/03So9+0zAO7UEW2Xch1tJRJg7aMo+JA7G4G7UKrIsJjaKj/QBNkaVz7Mj4QCGRfcR
Fj3oqFU3EPYYVzOzxOn5PmyTnLuv8r6aKfTEhZBM7URDpdN6f4z4SFioigelZ+H44DLrRUxYm1aL
XCvG2P9V2uZr6+9cJ1v75uCiWTHMYcXVGRdTwqiD5YOwm+AMYcnBieLQFBJaGGWTcwTwvDsgRTHB
wRBtSTjG+78gNgtpal536t27nnJhw27H1gqYKMxqtnuI5oZTRRPbUl0azOd5B3R3A2NuHrcR8LOg
xccESiXMNWGEixBOKP9iEfbxDQ8QenWVZiO4GuC3m5eYK2KJjhoo1hC86FUhSeKsd4S/YyB8ToAA
Uz5vA8+gjbJwbnXS/i5WzvftSDRunIJPoa+DW6YXh1l+oVufn4orF4zpzQoAl37bd+e4cljUSSD3
/eTvsLfW55YagzlWkHh30usPTLjEKMbyi1ExmFTksI8cHXONOVR6yrbmlKRzx6CZSuqPPR0Toe+j
lrurSirRBXUJ/3uUP2dfaFKnyYvxeYJ06IgPCbqLpCaLkhjIR2Kof8XHOOcH7fSwDtFJz2KYAtKN
8q4bmzBZYXG9oaP2iCj29hmV/4iPzupEPLr6KhKFh9/GV5gTmm1ECe+6lNbfHFV/MiEFuX1fuWgO
ndWg0g6HztcgcradDGyUBpoqNFG1I370RcTUjcu+rvgO9CZtv5FeYUfA52Fxi4XT/euIwp4nyCfR
TFcx0bDTgoFO5LKcJk9LUajI4RpZSVd8zrZ8roBnFPLt/g/MaDtZjUBzpqLZD/8eJ4ujfeq2HykL
NNinp+Ng0W2zKgJQMWTtwPk/DkF6HnriSeXG1ArF2CXqB4w31dmwq1peAs9Q8PXv/0pAAmTXaBTW
axQLYQMacbx02fx/srViC/KZUt7Nj172EyLjIlwg8IFxgqEIO8pUMtTLZRAqds2UT6PF0pEox3QG
6l8BAjIkZNqNx/TFRNjkRfztaFzDk/d6bzxIFc4aJe6redp5EOnmnW1f+JbEnj/U7ly6fTfyWT/l
p9/Z6WthKDrImo27atuVGr/B4B5504ULuuYRNujix5dt3AYv7B+QlR+lW6E8YltlSAJCklx1dMw9
amUzn8AzWHA6rmbo+IlJgOqiKlDr/KrfBBjZ8Ll/3JD5lPEoPBiHFt/xHgm+Bi1GMv8MLhmFR8EM
Fj1Pv8NFPlM04OHUwypOm6MmGEumBXvtt04O0S0rp1YKDX7n1gotTcE3MuqnwGsFo0aqKGKnS/mW
7JF29mCGokRe1ZTqrBguMBIauG7sqfN7a4vyw/QIYbnA/ZrlfCzANBQdMMFc5KFVxLtQH+T7EfqM
Q61ulSy2JWWdUnjnuv34w6HeMr0RLrlwDwYgwkFDx2zBP3nGrVmPkt+5JkzwdwJO9HQlausowivU
YqSTBJuvSqY5VMObFZyJ/NsIH7hEv/M+q54SatjTXCrCcwDYZS1dPNzGTYqWNrSuapsSdsas2Ufk
XgDy4MJl3PANU6ST3yFvZTf6W7fvMr61fUZhbZ+nUo2vXCn4v7BwWryzUdB46fk6qVeR7HnZGx+i
0qdN8dnWYF1ggzzw6SeBq7gm2bYL/kyY7QK6+IEq/zPgmw3BAitodSTAmK07iw1TV5mb9yBfACDW
P6XqNn+cKckfF/B7W58GyiWA7GHAttmTeE9JKLNZqsyJMu8Xs1WItWIVrmPpCdcnnjlQypyWj8LE
IHeUUnC+wC6h9Ut8pjr+8Xb/Wg7Gv8cJyAoq3doVFrMtpEDTvgg3ob2GKALXIJG9W1vCCpObPQL+
VHVmjj5E6WV31/6T69tZ05rvC1OAZFo7R9kMMpW7gdxiiTqBt2PEB8VOGQfl+lg/jAPTzvW2+QeT
FQ2a/vqxIweCKGjGQMMgcp5//B5YNMCy/tnA+JbTeNdFmHz9OmYF6FcIgbgO+EGuEVuvOA+wbDHU
SZI1kW7w+dXXoSbLBvKGnQkep2qHAqQRojs8Q2eU9fUcxK0iXlBQsriYYxyRq375rXsF7DhZPZ9c
B63b8y3AvroFC13hJGIQVpg7XRHeauNcAndxU3LBbbQvoMCREjJrEmhcsYP+zf/uxUd3VztO1+R0
WTSizuZaEtuZVzXVG4yr/YeTEQyPT4woNPCEERhdac+oz3v4bQHXscf4oNU2wjIUqYd+QRIfgdeS
uvBu2/ohORGDFzhMu3pUwIvzGeWT6vNu+dpt+0lAbW1kM9Fq/QtyE0MeOH4p+qBL+cLyKXmc/eZ6
oCpJ5GW/9VG3WQnM6Ava4GX84hG4F7HnFWyEi7coo1sX3eZ1/80y9FrPagNBeEt9ICfm9Oj9Pr7t
FV+75T7WQXUMVQXjkuBgMoeWaVb+4jmWFdZ3JTivoutQvD0uEZlmuRr+fFS6qo9ERsvRdEDdM39f
yNd6NoBqV9OZdIfZqSmlhnaLBffgeoSHLWLJQ/BWFBKqekIyHCIsVFD+Sj80v+D0XMnEDISbBOxm
CQFfK9wM/E/Ceo5jYQgMv0SLgnmrq/lEMLHmZRm3iFP1HdykrsDPWiWZ4A6TR1+kVNZGzYTstlr8
NewSVQYS8HP5j3wZBJPlzTZTjVbPKQ22MNgr9+euRa3iFKIbhoscVL/6v82G2ZG9+mhXFsIiVmVs
6AvpkM3uBNuOKRaxnaShJkurqtkOwnefl63Y/BNPbdwtTKKhL/IIESexDdg0bHeIiLJgWY4Qv0K3
/W5oe8YEMLcKZz7DgfQkeBV/mIB3/pazZLaFwaICMxInLBU+qn++b3ecoZAndQ3dTdgU4+s+i29P
H1UzsAqpNzoIu2TghyBRwoR0aSxYwYyTuRd93qKPs/sxqRJYmnTnYM037RElpGFlQppCDTCcY94c
Q/vqCrKX0zrwIn97UhwbjMBKdlHyGmWYPc+CwhrYSIASKKCv7cLQ+XxF12U3J+dINBmqRlTgkDG0
7zyMuUBJsSD60uuAdaNhc5oJOvEvWIWR0+v0JEwue9vvdbwLy/aHCCxCsp/E1xhKf6kzzelSquXc
ilAV3anGMBx3rncUhSY+oVKdhf8+zlEUXHrwXmW6YAV+C71NdpGaP3/OMSTBkB+CxiNaw+Udf5WW
PTg1rHz4hFNblF8uFCmBy7k4CnraK+XocHuZ/a3NVqkTaa5jhO30sC/zkMDg6Xxav3nz3MVwCRzw
dmkAs/vQ3zBLqpLBUSJOw7BBe1yaFSChxnb3TGhRWNpnJQ4Jp6D/+0+mZxcf4Jjw6XdyHrNyosOE
jQOtJOH/zViENa0kCRTbZ7IAmyIIzNq9D6wEF3136twY8Hi7habNhzYTAWkUe1m+MTxnHsJZGoGW
/mCa5lbK0qa7gwCw7DC2Jp90YPiEZekLIxAPL9RowkfPv7Y84YPJS8gkAs/nuXcRdIIfl12IDYV8
nHDk0lB3VQCLQ9mV3idimzjfbsGuV2+JWEZnQ7VtO1ixA5wll6p86kHxFI7y0wlPUSHFhVDgerF8
aI1meVLVrCSZy/LsN54S6I3mU7pakDMbgSopIKtLzk7+aJQyn/ZmpmcNJbwzwK+sceIeO40Ptbuj
35gIpCQjC+TAgZciJ+D0s7ZdClT5f7Q9PhgkV2JlCZDGpA0Y9DL+8dJEC+/yu5KYjxOFldb2KTO9
6eFtWWAuNQvfqZmP8KCM2c+RO5ES4A89ao4Z/caLgfAZFgUPA2+ela79QLXvjs1a3+QvvHdChOl0
VT0SP6Fs5e8UZvdHOz3cBbvWmleO0C8cVmq/i6DrLD/i2EPZ5ttVJ1b0GpKOd8Ch3OiCdOIiCsWs
oLtM2/iDWQiNsj6Z8qweOB9aBHiqLLFNOoLKMG3KC7FFuSJcjaixOhKRPExirj7xioszry81hGgU
Mmuth6Ab9FgAjGhcceKh50CI2HH2r2YwIGErr2tuiNbnna9twixMW9ZgvXlAV2t2q6OGfWGNurKw
MghQVeCJIIKh4Ay1Lnh7f2AFUREBcXFN7Ebic49EFJXlw2z74hsrBrbozuLz+cSrANF5MpA+aAdV
E228rNF8+JMS4uhrkDn56hD68ZCo4KeH3FVi5X4gbcSSYFhlp8OlRH1Ghkhit6IO/q60WI397meS
88/KUkRKiRk3x0Xyjy2hZujyFl6jHUMZNHiSK2zZE2jh9D6iBo7NV3VFW2e+7t9rNyQLhwYOZcse
bGyv4jh3OSZV+YqZXqGid6N/2QjtdX281w8CbwcNPtztSq4liZmQRrQOzvvh0YKcQBlMS+4kn8Op
/fYjIdlu6a9aZlHg8OwtHF5FSvxlyQwDNX1dCOyLFK3E+hjNb4Q34jAk5pKogXz8wXJW5o67/QYs
dujG+RETQcUwy4RE6Dh7Rt8/CU+Yc7QCvfVCgBeAOZYIG4P/J+NVq46kWADGOi4CK6XJXLWqlcBg
iOLgalreYyCxvxjb5jf+dlyCqkdDGv+q0yKQhLJJ690+9ZNiPnKhptmwshAt1qxfDhmXZeHWFhgp
IQ/FYcD+t+PWwc1fhRJxhETQCk+q2acDi2jzhCMNg5C1thsBGqyLD4fhkV1Ek7MuyiqwrXNg4k2j
WZ9/HxpF/PFyyhhmS/KS0MtVHqUsnMiGunlhsec0F4TAoWXJfRXs7alh7iloye0mh5nMyuvi1QTh
RhxtnXciVEq+VlWbH7EBmccpZqv/DJlgxec6ai33GzV8jQlhfO6m5CtNpEv0n91d/IBmeZeXJwU1
4ibqwdytUH8qHJRfFd5iqYCpdgHM7tQVai8i3GC8ygwFDCy8raDOf4774E1+fiGDVt3WrIiyodnX
lwj7RlAwCMKdvnvvoVNMr8SvqrdtNVsKXOLqJQGbSYn/osEpKgwfEeztwll3o75t65o45hF4cxii
KaUX9wOO/2EwVRzQS+RAtShkNV6WFrBIEWn++fc4UEkesaWad2CMeyKlojNs8txcIOGLJSaLetbC
HbfbfNyhH0sk95+AirlwpHHFx4UQqKNdW7FzyJn2zmpA1cbZ5qo5Du9+/+3XOKOnj6dh068irKd+
W1jamjSef4SZ0C4pLklk6pVSeDFWrI12cM6RO1dkqVcqGZhEIDXIRDjEL3z54pdfTLnLE26dtEum
aLNQnBgOWo75K/QhUZcpYqHNVIZ0CW/cfgn3/tuIygKWeq9rURLbUNqUvtdGPQRMGoYpmHCXLJgi
+Ynt1uOHIiTI06XJ9mpvuh6mWlOYa3oxc1JRMKNVnpiaC33Y5Qn4PrKnmd2jsXo457UdikPm7bGy
4b3OUrKz4Z/zHsMecg7tdcTsy9BfQKlGG9iFsJr/Jc8kdFRYx09lNCDbiUGalxXIiEeoSHusqqBo
HkB+qEhs0dp3JXVmPwvo8bTHwHZhSq9Dti6kv6GmRVqUXAsHE3GXSwtGFJMqtJDImDockVM+k5y8
E1Hkrzq04lmmwjgiSHB1098GhYy7OIxHRqI4vkn1dCJ5cpP+9J7qEOgckV93KlAlp4319DhX51Ee
VyOtr6g1bPzLM/Pq5819UyID1T2Ga2q9by1O9gjnOUb8Hv4drYfogtDcKUoSJasFPiVVI0Fk/WlT
MEsplpbTQGsHjnPm4OssTiKbOb0xnGw69qeB8TChixQP9DxbsDMT5cItvknDADXYZ1ahEW+GHdjK
uTPX+g3C3dao040dhc6qvCBdUNRmso7hozXs6eu5HPClS6D1YWIQLfQ5T0a9R75u0AfHhH3/YRIN
MxxiPWearYB+DgI9Bna+uox3/J0V7jomPni8ZfhmlQxXCEEcdotsXi1keJf0CcBKGHzJGvsagPyE
ogcbeUbUumYvc253kwt8UMsCYQWozOHuvmMPznsxM+TVSDG1d8eSqgE9c4i8VFjmigrH11hUMoqX
g/j2ZRzqJXokMlBKzoX9Jsj3hefL0z2xiyQsJIP0dGNYYBXzU0aCZqdtoXO6zba/kOW7xZBf93AT
i/Nb48ZXigreqqbN3xvbI8Tj1bU9XYpDZxxu/rliTXLNZA+loUXVvNPJRxupyaCmCAZYCvUn/4Ye
rpeBWIKVsqlyt3s/llB+oLKyMF4posAja63B5fy/RbnGDjUqRI8SJo/ixFWXglqOE3ABK058TVel
/4hHMZ1kS0F25FO/unfIxUb9y/in1QVh/+qELbrYP+O42a+7YrnF7bEpCFD5CHB+VXZmKa+ArFe3
nM5CD1Q8n3mHMQ+V1/xyh46p6RvQ91q9pC1hYsiylZcgZuBA8ucB7vsRf7laEEYb+Da4AMO1hy1O
vMdSoe+80TMbNlo3v7wYYAsUFurpKdl/HMggDvcYp7DVBxB2UHz6RSq7LGpdCn9j5YtclOD7LTHc
3H5j6Y3ziQimWzCLvkEhfmQUxrV+OKpOHYhMrPIgMnHMKuf7x5naOqnQf4Dy2uGOjgmCPw0Os5SY
z9Sa4p0wEiA9mUCmL0QBRzZyPq+kGeEaNW6w8hJKDTtgkjuugDj0zIRSmwVr0E+am3g4LSYWdjA7
YKrarl5vDKJYjWgZnZXflGkBmZRg0MQY/Fmr7YTRVb+0imOIBK92aUpoX9iwevT+vlHuATT59JWB
ypX6nLJIzl87twFi3Q1GCFORAaP+DkiSX6LOGhoVjN8py9t/Z4kh8P8y+1zIJNdRMQlXaCVAgD4h
q948ccNZSOMGJkfD9Oy9SRGBiL5qSkag1q50OT2gdN0LWbjsGAvCRY4mQSFdiKZrJdew9BoVJFBc
G5v+Wh1O/OUZQWKRuu3LVNQEYU3SlWzLtyu6NGHaRq5b6CZ38tYIl01K9xU7umJa1QEPYQAVMvqA
/DhfcanXh95JfGs+e2fqgx3crPM0DE1R8zw5qKXDSHRSwLXJy/iWi30V97XyUeGJrFRULcEpUJLS
G4/QubFs0bk7tmveVp6y8hrBtipwpvWcUDv+CD6/L0/5ci7AF2ZlmTyHVxoOOHe0TfJFKvHh02lc
JV04fRFHmCreQG0CxJjAUXRegxPq6rcmCtLaP00uzhidvn5gAgTyzWjIR243BPU2Yr4c9PsOzA9u
NwslBqDI6YFhFFEHpMsBCgfejuqrgQer5/bg38BMftoHIROvrm6sB9sBn9cWRh7Lt0fmoV8t9/Lh
3tGJ+kDVupMFXvMzLupDB4sR5ujcw4jgqtGiXQHK8nbPFsV545IJk9m9vPZlldlDVD6vRcrjTI5X
n8QjbGF8t/0wMGJaA/KksUn1OPpMGP5YNhqKFCFZhqsxC0zaBcjM+0d5siWgu7D072IfIphM4F28
DqLDq/a0xqf7jKa/N53CnHkKpk1r3X9rqM+HBgW7zu11qHGvE7a+0CmiEHvuJP+xB0Wn4hUJcIBO
9EiAprcoziFeI53yJbvM9dIaf7kpJgz2RKN1T8pFJGwsjwI88qhIkDZwTB/xKbS8sZpfWXfpDZnD
fAzsIJenbvF4+/zUdV4g6WSumx0i3SRk6ZxygY1oMpB6OaWzu0u4wAF16pVXBmUF0j9m+sjufhFy
Lh5zReXmPzpE8xl68CCzKvW4Oto/hpbS48hTkJvS02tynGLnn0LEQSiytao/vPFvaST/AZH4Oiur
02aL+D+P7/Xj7GZk3VT03RUAOsfPDX2yC4oDkDJBYJoO3MUINvwUWZnRKdoh1wtKGtnr52R0LsqR
j2M0ZrcA1ShFchullHzOPq4zPtcItLjZPCZF1vwKzL1tdK0bx3TxAWnlslzWuSJlJLSdopD3JGeH
wecrs/nYgMBlQjaolrC6FbQRXDfrZ6tbRzy01xSz31blK6u8xibpjKAD4g3SV8wg77K3w/n6IXDb
KMHqClq9A9dgjxNX2NW8YC9CrUD1+hWLm52/8D/4YAvwddzscb4+ZN/Pk6wmqTyAPbx+qqfRPiLQ
MADR4BD5nC4vnQqBzhwsNRgVMaynnxO4D7taBQHGJTpcpZ4oQrboBTtDL0rp8qIAyEGvoE70H+PH
ftdaOOSCAN5QV/l5JALwVWIPgyD+Nq0N7qc3EOTU13uAK6PrBpAoY5dXnapJ1i/wegKCE0njDkcK
MfHcEh+WH7etgQhNig1mYxZcNmp/mAf4/SoBqcXS3tDdo2w51vP11apSpe+K82EdwZzKJOxvtPua
gYUle7BZbjHdpf1sEYboOHiWKP8uerkGoTtKVlybv90rTGKYAaJrNYMIQmlIyDuq3LK6+ppL8Q/x
SsZ9dbfSpTpGhrWNbo9XZYqlw7jf0xBis3+dUA2GW7/Te4rOrxCR5Fpjqd47iRtDuHmp21DIAzOQ
LFwXiM/p9KCsXbFL07XlT9t8U7iHVXi9EP0oCKJqIIlAAA78PjOQakK3EjIesSL8TzzHR1M9asJL
RhBMC44h4sfBad7CZ/DvS2P1VaDvHXbNXIN6k8L5PVxzxXzsDxgX81G8UxPSWW27cx5+hy9uC9V/
WWCiAu3JMY6C/7vKI7B45y5knkJkdoWVseT+XeKFsA/WO9xgjMFsmIVpZKS/PhaNguKeu/3NVrGY
sDfv+20dj/OpcR+sBwfWDq7i09nJc/i2C9SISzd2CQNTmVakZzaAZ4Lf95XmarL5bktOUkcFFfQn
LDvEKB6VO5y2RTJs8ctBCn2h5bv+/Mg2VAFsOi2+lss0r9jcdAUBG7m3LCXOtMzS7NF922k/2kg2
KY6lyTioJKX+ladVrckTwPqIAMbjgTONp4PSsC7+3qwdebKtJqAgsz0wGRiYSAK2/xiMs+UN+x7N
t0ClboGUJuUxzFhP6Um/CXOtbCdkKECKmp3t+npZxGKuc8Vk62DracjIXrjH43nN6j1vwxCNP3tZ
5na2/cVO0wPGlXsb2ZBjF32R8m+tJGX0eMtzKKIn9lW2ERsOojDxAxk+JGlPUQtQ96q8KEnKA5Jz
3CE2jpA+fsHdHfY8RgcaiKxtsa35uy6s6ySWPDFceWMOAH8QG3GKTPZcorhQJCirvENevhglls1W
2qEFLOKzQ1Y6fwqV+xh4GAZIp6vu/aZJohvMli+Y070Mw+IwOeYGjSb4JFFkW9iUN6l/sHPjp29g
JkpzsjgFrZn3jnuNVeV2PGFJzSg0iIu8qE1I9xtrtZl2LXFb1Lxw1lKVeLOqBMFrKKaiDYCeM+Sw
EGa8evRr6HAwR1Lr41zb7UnbY8GY3Nm+NOpUgHXcpj8iRDC4HPItiwribQWAqPN5Wd4dIJLA0osj
f/KuG+i5EP5yIsUbq55PR/WtKSs5hC6EFuFUahQl+YWPAjCF6shmax9Oy/9f+5joqCuAO/+wYKd8
IfVyq5DyxSivrjF2y0UrwuyMy3yGND3M/QChd3rrqWfRxfIvHBKehBro3Jx7L7UuidtmJsb49d1H
8TM8tjv/yPhsgEAYdVqnDwgg3RJrfyi5zwru86ZokdgawCkGRKoBoWiILrvW/xcB6a2WxkjTEGN8
M3aPbx8KWeNqsCEwIY+8nF0NAXphwdpu7Wn6lkzWl4xiHYjnfn7nvI679wDfP/yBCuKUZSn3V+va
aQInnP8GqT8EYh0teiebI5GqlvTUkoTz1kTVoUvFDoWMT+d37yt0yF2qNgIzX98Z/hvmvAHxIgB/
gN8W1JbHUEhZfDg4osBkbi8G1mTO1PH7xcUX9DXbQcqcolI11Js9gsRHmr2kQiHcara7cCyQsdKH
P0BqgKWPJZWH85+0A05SKsUcYzopDIKbMHyAftnbvrCu3Q/vIMFS9I+SR9+RfcsRxssY4uwyA8Ug
j5QMT6eHOwF28URs++a9JCb01TEi9G16rVXwIcVZ52rBW+wfzVDHZbM5sva85nCJdrjaV5oCdpTp
ZDlNmis+/wlfPuMI1g3IRO0D3GbotarqUi17T59PY5IFpLHf5GNILAb9nhdLY6/1zqW67q6CJwzC
srIuP/naLPVSqycR3TcnDx6QSIiJlPerGuvHXaRdCjlqteaPHm1Ld01dHBuF32hUEticxXN9NKha
QGVPsWhEzVHmamowpP66UieEgLlNu60X+cWgl1xVRTKwgy1NLStflHh7ddg6fqmoCsjV10G6+A+U
YD+/Vp3DriGS17zm0XAu+4fqqEVml3HIHsI4o3eRT8PC92tw3IHvN3NGw+lQH9oSTaiKZ8mgwsZc
wiLXTypXxU/YxNKBanTdpoYKoh0cfZyiTNOEP6S3kb567ljjqKDPmKn1POsvWw+EShrNnT8FS66p
sCJ5mGGuOyfolVigWB3powwsVQVHvK7lWx3MN9cC69+6uHdOfL5yIP/OH9GlRjrekxVGm5+dtgYf
8I5GcPbKuL4pGnYXzhCQ9utydCcb1trtEAmzoSuQxVmDkbDHakYUwMHhNFOrnSqig84KjaNKu6yO
bX6DsAipBANV4artDPfHtGnMTAYGiqYtKboVbEWq4tK9VqLkuW0Tsni6WKLkZgEbD5Mj6f6pwVr3
K8jisMiB//02Rc9PRPo+g8+mB4EjHES9DPC7fTwV/3us8lFb0+N3gcE0AU+ggSNKlvLrXfA8TSKv
86w9SdHgYQQNTGLU66+4/rABNMZ/Fh/mN5dCjm+abVnqfBNdF8VYGL+as5xRP2u4TW6bIeTvs+MD
SpA5FWgBnCSens6WFX3VBuLGUZqPBHK5VKW+EB+wPozd37qZhUXyvpTdRJmap+6KWgvc1zPtTIWy
DWC2KY0VFbgsAkm3yV+HU+u6l1u8DpWwjZTv/JKdrZ4al0yzC5qccPZBufJsMMC91SLQX/kiAZk8
R2YhuIURdgaXNwJtGRDanm+kClTRTSc//1HkRVhpFVaES2M6j2oOGxGHjFaMDURJ4DM6omRkan++
/Tr22dp6OiVuSJRnWQorY1lNA5Cgwbvl0aVpcOWadnzo0/SBd/6PaixR/GHoUWXDFS4rNRVfSE+Y
/BFeRZBRJZqqTA4PNzxFpgEFEXPGItSDFHBzRrv3WMa64bmQFmGR7Ov9HdWRwDwyZPgo6vwyy5At
m+zF3buqFoC/vY17EdsFnjga2qHIuKfXmup1XPVVi5CAHy9dQbvPi47J8n1pAShNaVIKBbgAcgiY
ix7cC2ubJHMz9458pmXEfvk/fgYBNkL4NVBuhfdGw6wl426L3NQauyQ3HINiv9o9jFo/UbNZcJRQ
O0Pblr3Me5jJ8Krvf4QPtwk+CaA2qVeJhdyXm8EV6EDjHddgehW43TEJtQV7J9Ys1rKx1g6Uxjn+
pd768wZLckTDABXuokpgSdbiW+rzKCpnWrSrhuusdUd/DivLvW95RWfVi80GAArHok9O9OW5JyJx
l9tnoUNt+T4G7MFm34du9wIXAfDXD7vad1S+yPVspXwApSuckUo5D0QOBB4Yep0PvDdXmyKO0tUW
jhB0ns2dk2ZB4mlFq79SlQPuFCYFLkrx4q2SQIbp6D3eMnFIMh+L/gY9T01145wOQQB2F42jiXVC
/DJdLkfsnbiDa8drXrTdxPRpSJhmSUOIuzXPcvjBtgiEaMeTis++wl5MmAQCxzqWmdTpGDH3a2Do
L1NvvB0k/a4IUYocwFfVYpdtL2FWiFY6M/MUHRVxNFArmTGvtZqSdtszKIWbkh4yKTlFTC97M3Hu
pdmZFUc7cBUvhrIvBBwkiuBPIDTAK+7bDk9Q/h8fUPeZ3eA6ssBmVXhi+uydiKroG+EpNSdvfwW8
qzuJm0xE3B5nyaDTBM+LoVjsFr2VC0w82OmVJr5aNUCaFv/FajSC+QzVjUoCRSsSj7N9sjjFdj9M
SfrQN2nB/PHar7bbtzyz6C8ZYNjuk9aXDzeWiNmNoeg4a6vCELve25YWnEssINlKBDDUTyWGeKt6
Fs8oSwdFBralrW1D7J6z8fq+2r0bZL079v9p/wBICfBmws2rbMW1YmUjSV4MjY6ZZhmw0riplSjg
45+2ToTo2Wz7I50vqOG0smAGifHX/HnGW/iHaey1iEsI/erWT49orKODA2uD2i3IqVLqD4wbekXg
V0u5RcnnN66+D0NBLINYjkHj9HItiKS9/uQO7Ul6b96TtC+rXqK0Q+Tr/d/+1NgROSBa5KOZQQ2Q
JefaVK5LX+UqjLz+vy/4xQbRp16joP6ua8HartSUvhyTIlVDGV0CYsxD+pSei0Uoar8M1mh9M2x2
acOWTBbbH/0rQ2vezi920TeJIoo+4Y/CKnu3zt/eUI4p4N5LHIn9FR4TAKjYJgkeqPeNbZbe1ndu
x33zq4jRiS52vOEcZWk7vnQi9yAXqMLG0D3g9j3BPd/LojVHcBQWfXVpDbbri5lb0qtqziNEKVgu
e/j7Wbpb28Jy2Tnfk7+aXbxee99v+8rsU1jyJf2Mf3qfoQ9uugScMoDpDbwBIdiky+5ChsWOrt76
DfOutT99kQH8E19tLI0CNszrwDLT+7Auv07jVs4ZGRJHnQ1ijsWYeKinsPBaJF6Ql2Se4wTe7Mzp
yuYcITmUYKSEvL2jV67/nVNI3sOsDWqMjy4lLguwK+6ipFPZqhQNeqMFdn5JsZzeMwtMu0iMFttC
kAjSYvOgepIzwdHTyAyMCTnP1pRgqiBVqhLKGRdTH9YmLzX8qZP9DvfXRpIV2jk0RVcOI7ZsaNqg
qeNbwBMT+HXKvd2Usc7r1Ojp9UZ2c7TPFATD2Bnc+ARFusuBPcskFbzWM4/5vLOTy4DgvhSlbVBm
smMNkxl+sO35SVZjPzE4jhEy0t5NlLkLA/FbzonCTa67N0yGp2JUx6jjw8W1NPCru1ZSwuluSvYQ
PB3BQCn49kmlJYWarbdN6OhyA5w+LKOhoeP/UX/gG58j4RRvE6FMDmE7B+nwlcWGuAZCUp5/ibbe
P2cGCAaJz/Je3gadVWn9gG4A2cRrvP7nHzYZdGj5LvgnWdFV+X1cK1vrnkJWJKg5SFlNxTTehg4P
U/vRvRtMvWc2ZTDeIO8A0qtTlWKGEdAnIZXQdAmgv97q25XZZblQxhwcVRJRaDWFxnqNfREIrbZs
pbNgqf8y8KopppGta1JWb3DG8Kddxvl8TXMenU9X85kKCIH98U1bR6qzKCXS8fWKGz2h+9iMz9qG
dC5dGq1duW9P/dMbCaXFdsummLn02a7JeD0DMhK8+OcGPqYXI8I8m5jD6OFud5FFScErEkMcwYJF
kttnUiqcagMQMvVJZWfXgoDs+ugVaM8oGBYp332ht90IjlUZzO/WLfziIcStV+bUjunyj1Id6kgt
/SfJUHltl0qsI2MVooY0LKlsD9VO2FAcJ1JrDSiqHVlHRmYYsn9spwqhHRj7zmPxT3+dqQ8zo/28
iE3z6VB5+uC6lUmgIHy0BR37kRJO5R2h/Rbch/jRLk/i0TzgCUBQ0Pce0f/f0lwrb7Tzi9Sce0Ge
LH2kqF3B4VjlcPturMXlsCalSbom0/JJLwAB328L7x0jjP4RWMHJr4ANSVrkf0TcpWSNlGvUtQxj
YLe4wUWG89AFNW+AxgY7OdZwXOcN0MRiXCOF1mXV0kyjH/fGbCEdC0ozAOiKqMf8Fe9falBWu8FM
g0Jvp6zH+z+8njenO+8vjQ7Be0T2sJwRxZDqWSZAacfAYhKYoEgGW2IhbPoCfIJpd4O+YzXamcOC
xVR8G7HBaI7qT3FtPhDygyqlTZHl5YmcnDyzl4cZ4U1Ggk2kR2AfIGILB+EujXtfRi56gk2AR/tk
ukYqkbfB02UuBVqjwjxydtl6sNnzr9UL4RWPlEUBuZkmeBBWSMQ2t9D9a3DjVQe4OulnvcjvHyZZ
Xjs+Yfrun342i2jA3QFiNFwyZsZW/QNi5SQBR6CIJ2GXOQQviOaRMAQkf88SnhWu13L4dPbQ6Byu
kANHXdeUxkosBEJ6khF/xkDegzXDlSQ1NcuXd8uYg5P/iSDiGmuSXTbLpfS8lGN8Pjf9dqiqC4/Q
NfO2qfTOZKVWKqOXtA3rYqu4TUGDarL6MV7rfeH0VNdWAmVKBj/oLM1vNiPJNHqtbRowKaha+UA9
cB+f97bQJVMRM+YeMPw9Yg39aeVizKNR5d/NU7eROyGUJtqxZMDIWzIoYxtxWVondBpx3d8js62D
XkKuUxF/8ylek9EwSWmy73ohbAqCHAdeRTn51qdUdzhswny6iD/yTMRLqYgmUuzag6e3PjnSnSFr
J0gNElihR3T+i1G7R5XrzcNyucH2GlJC4M00roFGZ0hHP0kEAOH4einqLoTB1QHGg4U+rYhdtvFW
PlYqJBB/WD8ZowWSLYiWYEPE32f0rpnpKrG7fokG9C8hspbp/xGB8LjNquJ1y7Vvm0ICqfcNq+Ev
f/9/uBVtEMjOncOoCKAtDIgcIpkrMbApueCC8DeiuEUIW3AfSXhF+JIFxix4ikDFR7kpQux/Uayj
4af1tqAVCrvhNma5LEVb/I4wx69mXDtBiDH8nsDdONW0GfKG0Sb8U8SxJG7/
`protect end_protected
