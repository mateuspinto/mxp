XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���6��4���"��]�Y@�o�^�{BI�����8(G�ip�0߮�J��Dkz�͎�-��"�&А����7W�H�� '��x��弋Tei������q:���%5����w?�o*~��=�	L��k�����%9��lƀ{�@����
~�H�5-yV/f>/��`��01�{�����c@'65G��`��3c_Ԛ�ח�i͆>Q�E-jXL R��;NZ
iSN�)�3�H�q+���
Q%0���5�0�\��2�����	_�3�}F,���F(X�fa��AIyqZ��I�#�"q��f���Lӄ�q�Q�n��Q��sC��c�xS�IK�t���Ҋ���8���ا�5t��@2�2�:��N��I%��������F�^2�J����X�Y�\P�G�\5Ũc�t�v�O����IL@�;|	�Wd�
Ʀ�B��7qd�nFE�B�c���<�?�ٕ(�L����وB�����{�l_���%��+>Y+I�������u��ji��F���~�3͉^�[��mJL�?g�ܼ��\�YΊK���S�cb�NI�F&Ǆq¼(��[��:G`�H���H�>@C���y�ib3Z�"�F���BeT�)�xW�[/ع7|����Uq�U�"@�IѝNb�@�Q��ԔE�����������5\̥�Q�7M|_vʪ�`�
�Y��+z�\�0�!�b��s�WbPV��4ېs�iм���TC%Q��<�� �{�y�I>(���a�9J�,�t��XlxVHYEB     400     190�啙d[т����쥠�0W��f�9��7z�7�/�۔kj�M��C�B�F���*��!�֌��ę	,WհW���B	�̞�]�t���/��QD~؁e��P�a�{q��)B�G�9��,��k��U����;��*ۖ� 
����Ͻ�Y�Ύ���%ٻԘ<�6�z�X�A�z����l�)�v��r���
�+��>Vmn=�jեO��_k�w0�2����K(�@�4$�O��@C%����\��p�S�!�Ȝks��vq�a���ϗ���)i a�����=��"���Uq,4��L������� ���\&8��I�F�{�Iz�|�X���e=16%&�#6ב�0�p�[���C�K�l3�W-��x��` sޟ�jʵ	��C�Nu�#XlxVHYEB     400     150��D�;�����s�>Ty����`b&�K'�����!�`��0p�@G���'vِ	C}9�OR7
b��h#���0�~���fo�Ԧ:��CPt.��Q�F�OZ�����������r6�\��n2�]���[�z�Q��6�y���̻ws��;)�@��,�OK����6��xp5���n�H����*���B��"�Nb���P���3�gtV���� K��nj b�.�W@���4e��,�E���F�lfF��S"/����}^}Jp�U��;Ry-��x�ĠF�?�vJ�+���J�_�{+G��:�DZI9�n4�E5,Ô)�H"|�6\��sci�H+��P��XlxVHYEB     400     140��R~�P'V�W���I��x3�<���a��#���ht��d�������Tw�hzŃ�c��5��^����C�7-�}�������Ǘ9GL�n�/�o`��:m��l�(&������s�y+j��h���j�*#�"���w%����/����wE�	p�ܑYl{�@��KZ2�����M�^��P���H��^�`�i����H�<�$�����l:,�Z��TIgt��M�D��F�X�� �Q?ϋ�L~�Ⱦ�4����-��r��ss���m��Ķ��Z�����s{P��g	i�~yu����ɌXlxVHYEB     400     180[1#�������.���(u<�ߙEVfҐ>����A>�lN������[
7��;L���7��e�b��Z�AH�wV���+�K|?�̾`�)��4L� ������W��e�#�>���r������f.��g2��}��k���.JR�ءSj��k��g;p�R�i��IΣ-!���`�mF������j��l�W՘w�>6��l�L���j����)�%=�X�J���A&s�C�k%���R/�_�g�퓿{�?3M^��HZ��p�Zy������i��|p��^WCP�m+K)|���Y̨¯��Z@�z�+Y�����=�U`�v�{{drS��X�dD�nd�b�h^�c��"���[j��7���}8XlxVHYEB     400      f0�頩FM�	8�ˆ���L���Y})���#T�߫�!�w2=�_���nZ�e�"��e�Ƭ�,����"�A�:Ջ�1X"�@��M�=n	�ta�^���u�Z�J@�v(h��B"�ǥ񭪳X���zy�M�@؋c��\K�3�'�7�+Zn����{d܇k�ʫ�[چ��[��4�|�E�yNf��M���E�@�u�ݥc���B (�F�UB���#��2`x7��XlxVHYEB     400     150���IYoO)6��ٓiփ,3��7�N����|��<h郺��Tz��L��іƑE��v��ڡ
k���WwA��+��"��%ј� Q�J�gqiTP��"W!�� ޏ�bE�X��N��p�O�{�w���~��_e�Hi���U�G�Y������J)��s��L
����'��ߤI+[�xxj��k��"�����v�0Z�7#}��߫�7=z8&��>A�	���x�V�Vf�4�Yz���g��'
�Ѥ�a��F���	z���?o�T��x�� �+�݈�9$p%�3�C!R2�(�l@�T�,dv��ݗE��XlxVHYEB     400     150�� ��^���R�b]�aC��NԻ��c�`��#��Z#���<�ۘ��hW��7�$����0f�V�a�h~�L}�$��tii����G��7e�FU�:G�5[�z�J��7��3h['���j��d��`�xM��KI)L��  ��eJ�æ0�0n[����*�[ǶN�Jb��/j�!�W��V:Ag�[�	��:|����k�7�|1�v�|E�5�����tl[�e�I�J�1�?�������:���A�*ʈX�}��RZ��.����#�W�޵�4|<j=���C�}L=���Ŷ<���K�������YZSu/�ea��\|�
}S�3�RXlxVHYEB     400      e0��ё�X�y��/�>&C�U��G���v^e�A��ɣ�~�'��F�r��&�����mX`�N��wJ� �%ckg��ߥ�S�HVeR[�Ʒ:JOp��/����p�q�g��SK�RL�/C�X����G�(���q�|ӂ�+iZC	*��P|���oa�s�u����������W��uN~��b a�c�4��S1 S��U�ǡ[=!s<��X�)8��/�1n�zXlxVHYEB     400     180�A�-�`N*���B����� �������k��ɍ3Z#*�e���J�\������7� �rn�|���:3�K��.��Q޹[����3���̿k\�?�÷�ɵ�2ys�����Bnhg���-�0��h�F)����&]��������K��F��N���|���1��D��ɐ)*+��|�/'l,cS�<����� �;J�U��ʆ��45)p���/�W�o�v�ٔ�w<]�.�)��t�A�`H��Ć�A��#52ʈº��Z��A���R���Z�]X�^>�T�\�,.�b����.�
 �2y%�7�������1#{G%C�HI.���������n�O]�s�,?���?k�r[�	cVvi��.b�����XlxVHYEB     2f4     100��$�U?�~�zی���3&C�������pja��V!�9�����XǊ�7ț���pymg]<��J������'�o���nZ& ׸�T�S�@Ϸ7�NB�Ε�N���1R�B��v2}-W�<�V6�V���"�֝����9��5�{��U���]�蒺�����vյh!>W|�1L��TPv�,Aft�9�Ӄh6�h́-��W�H}��{�F$�}s�~�ߤ��
;63V �@�jo��v{�