��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���L�n�����68ۇ�fa�F. }?DЄ��ٜ{��HBer~�k<s���)zk���1�Y4)�H�qIIZC��p�����&z;%�3�~��`~�/�2�"��7�����5q����a�p�QA�-ZG�{��5:���s�~� a�<%ʡ���N� 3��ا������~ BS�JXݳ��NД^\}`��$\�&o#.�E�Wv�?�P���,����}��������<�����b�𴨅�;�vo7�*���v�S���bH2����Kc����G#��֨�m�nF�Y ����	I.��@A�M��D:��'�T/���7��r�U �d><�)�K֤U��4�3��������n��W�t<����V��;�Jό�u͎'��׫~9�H� .v���e��E�����![`�������������˲����w���<�f�^��u����.p�	��*Ƽ���9��-�;�����s� �L�W ;��r�����qC���x�n����D	�J�]��N� ��믓�즲([� ����u�Oݢ�&2g��>�7�GZu�jb���:�៫cW���u5W~3=|�#�u��I|�'ZTQ���f��A]�UX��^���ļ�Dt�+~>�Ҽ
�tB�0`�,�d���U��z,��j��C����.���_��?�%����O�wnz�ɻD��V^eթ-���?	���5�7���ӣQ�Qy��x��TJJ��[U�b�0���L˄�*H��rA�k�l����Y�"C��p�@�4�0�����J�~�x
f�=�}<ی�~$+g}'��b��K{�c���J�ፐ��6-hz�=Z����g�-7�+w��DoC`�9�S��pFz��0�[�%�ˤ��1�6�� �\�6�Jo��i�ð!�`-�t��8�Xcl%nMR�����c�	K�>(�S��������wB��$w�f��v�]D�f�`�,Y�P�|� ���Q���N��Rʺ}�, ��S�ؘ�����<J���>�ᯓv�j���$�j��������Z�bit'�ڌI�Pm?4ߘH�WلR ����ݣ��ؘ0����c	-���:t'����,á3_��Z@'5n;ի�Ї�@�[ϖ��g}��"-ڑ��xk��rSb��?x�,��mə>U=���8�-c�)G^H�^���%�ⰲ)_�����ok�t���P�q��� ~;F7��6�����G�����M���qi��`���|]~܁/���:���|��o!o~�����V(Te��BU	r�lnݽ��Ky��YTr�l��y��EC����.��ʶ ���V�PJ�7������'{&���[?A�٫~8e)x��@כ�(��""����#��o����l0|T�_H�o����=�����}aV�D�Ǳ�|c)T���tȭ��Z�����)bo�A��A9�'*� x1w+��Ud��^_Fh٥����%p����7e���R�����!��>*�ŋ���e��%�.���\��W�m�-����v��G����
ϥ��9>�x �Gg%��vj���2̦�6ޟ�F�t%�ԇ���^��G��w玵3-� %h"�_L��&Cn��E\4���Mr6�*�J)|�1:���*Bq�=�>��,-�SH�!d�y���Ch����mʻ?�b39M-�'�2]j��,ѰJ�Ź�`1)j�wnLۋe�0)���r\M�[�����UOgIb9��"vTr�=-�<#\b"�홳o���"S,����!�S�f�����ձ�2ԩC[)�q��[�ѸP{�lT߶T� w�ȁs��"��������`7szo�Y>���ޥ�K��5���^���V�]�I��W�s���Kb�|�hi/F�GóN.����M ط�=�)��z�"�/�j�)���8$;2���!�jT���4���ꝣ"4lY=�T���s;��4Y�f��;=��C��!1�F�=@�V?���F�T����y���],Տa��a��4Q�øO z�T��R2�u���~�)����Z߬���}�^�E��%�SzP���!�ǷʐtHv��"i:�u��f��'�B���|_�# M� ,HȒ�ۦI�B�k��CX���r�]�ԅ����c���}-m�G�2ʄ��� bT�X7��A�2���]㯰/�`:���t&�}����AN!�6��I��ke��K�����0�e͇o&1��e"͓�ʃ��(sUUK�Cޟ�6���A��9�F�}�ͬ�\�wC(��*�:� �Wï�cZ|�M�)�]U��w۴�&V��f�N�j�HF��#�����ҧe�vR1m2�"n�S�*�1����_�Ä8_ﻊ��)_S�v��T#�CxYa'`����;�����VBt��2`�h��D3Eu�}����R������f�yP���(�A��3G�X�G�@�jVM�Ӝ��3L���_p��nc�&sn�1�EȣP��SƇ��s2�j�D���w���i:y``����YX�!7?/a�L9G8Gi�y���7=�}��?F�����Eb��:�)�Hp��Zz���*^h)�v������1J "H�(��������6 h0�r�5�Q��1��t���r[TYvT�Z3n�ۃ Q����$Е��Z���vd�4͐qL�Z��2�;�vZi0��״�\� �f�t
C�z1�,����op�)�ȡ��m��$zzr3�iɌX�U�b��-?u,[|�U굛ڬ%n>,�� �M�ݙ�m�h�z�0�^�t=ߺ��5Qb`?�P�"�����"z�*'d�^�ҭ2k����n/v��2�(%�Y�W�4}T��ܴ޳bA�65{$�����������Q���}��J2-`K�o�p���J�;�kJ����՜�~�������r7@��R�1B#�L�xĲ���������M�1�w�W�B�!E��UL���|#��wz��S�.�����k\S�_@��L���%?���<�n���ީ�����:����3�m�0J��`��ɍ����e��;�>0���`���i���)��x�D����o�5���h%6��#��[��^|�x]��qefs6A�v��(�b_�d���"\3v�����4����I���H��x��]��9�R	z������J��"���ډ�z�.��C�<c�c�lpH�&���O�x]ܼWp
���*����G_	g���SZ�9���d��԰�[�5{�J��F�ٽ�B��YȊ��p�'B��n����m�퇦�C�h{�-9�úT������3CAFp��`�. D>T�tEu�i/�IN�"������O�,N%s>���^���Ƕ⽚�]ю:\w�'�r����='s2���6�������Ӌ�]�EzOC��H�eU�^jwtnU��[�8������a�t)X����ʊ��h�y&t$��%��}��iG�L�����DoYFGm\@ �`��e�������%�,�ݚ�N0[� &<j��6-�)��+��� ��l����py݋p=�i��!κ�����EL�� !����MV�À[�W3r|UT`�3�MПΆ@��Q!eJ��ئ�XrT�2�Cv�?RE@�v�ˎ���=Q��Y��~5���#24,i2H���s陶7J<H��7T����o�8ݥ���a����)�x]�8:��'%9#6�����Cz�}�T�3�Ե̃J�g�.u��l��YF���]�w���a��U�&����ȬQ��l���'S��ԎU�~'ٔd~�xaz\�W�_\��}�\B���RZ�t�t!h��h�J�)#x6�`D�Xk�ߪM��L��=��oA�o埉��!(�ʢN�߭Fu�08&@��ޭ\�{A�z������L�Ro*�&�[����5�z���k-�(�k�Wn�ѭOC���+	f)�((�Y_�c!*؅�Px[C)�������� ײ�K���C��%.+ޭ����I�J�Sf���h�X�9�i�ixC�Hto�&�愣��c��w�#��½0��9����UɌ{&`�q"�$����d��T��COz�#���&rf�,���n�6�X(��i�$(�&yoP�F�1�#G5��1�G�)3�&�.a%%9f�og���'�s\h	KR�G���G}6�_�k����#�_�&�����Spa+��I�ҬǦ��s����ǃ��W�>{�Zh;8@5�KN$�3A=�-�[7٢Jگّ�����4���
�J[���]��!���B����{��|�k�.���kA�<G��+����`3��a�G�W��Q>�U��h��$F?���1/_�9��+��P�ay����&�`X�bJ�r*[���؉>b���|��|13'��B�Q���5GO�S�r3ub[���A�}&��NɎޢ�=I�*��|���%��	���,O�]�އ��ʉ�>� �sp<'������k���3�ʥ�
t���<�Fش��/�d��Tq��żrLіiKYz�K�6靊�yme�._���7��$��}�D��uD�_HH�����: �DW�<)R0?��\:ሮb��${w������|�lZ폈�z�����9���Jb����.��7zn����і+�:?:��B&s0Hpg�`�I�Wqy�IY@��-���g}l�hs(r�k�M#�a�|0D�3��*�0� ����b<D���ӿ��)�`���e��f��g�5H��:a9Z�U5�m��a�O��"�>b(.�A��=�wY����W�!��]��RhЪ%
bn&��jjA�#�L#m�Zϙ	�ד�Xu��ѓ��V�a턤8�Z�����q�o����U1�	`���������FC��S�Y���_���$��pg|��H+
�),d��v[B=���e&��2ǿ"��M����qD�E?�v���OO��..�G��=��0����$~��魇n!�P��@�(G�⤨��J�%�m����h����O�0��W�,Y��K�i6s��_Ĉ	��EԆ�$ކlyg�wXa�[`�"��� Os�
�H���[7'/����pz��Dyb��%�����=8�4#��	��.S��ݺ�L��/�1e��)�}�"Gxx����x	h;���7R�+\�<?S���1#�λ6�.�٣�[��09�IF���e-.
�����d%T��׶�������f�L_�)��d
6'܁4b��{�Av��Ȑ��,T�U��j��"�7���ԃ3���Qkj���B/Dp�FN�n�{����oY��n<(���]?K�Ⱦ�O�ܣm�o'N}ݘ��í�jD־��#HN���b��b��i�~��79\�흆xc�'���s'/I]�ԫ@���oqEu��f�d'c�v'�<�n&sf1��l��Z[�&݉B.�RGi3vC�z"����� �ID�#J�t�� ��X:���&�����MMV��3.
�8���I�A��D��s�K��$|M��ե�"�E՞�HmM��Q������ҫj�"�P��V��ۈt�g��-\$� }�����~����vz�X�;�;S(��@�)[t���G8<�,�==��B��V`^k�̋�ѷ��E�&�0�ȼ}Ԟ���Q�������_�_t�5^�[�d�?�C�?���^Q��PP�1"�;G�4�ŭ�~_Lw�)�V�a��$s���A.�Ĝ�|P�W��3�)�di'L���{}3V���6p����V�y������OOe�Qb4p�y�`,��\�Q�0@+�����:���ԔD�0�O���J=aą���4)'0�y�x�a7hYř*�iK��VI�Y͛Z������aeR���ʺ4$)>�Y6�[i�z�R���i���>� ��]8'7׻�ҟqh[c�E�fO\�G��~uCtO>�@o˯�e��Wp�[IQ�h����k'��U`Q9[�k���>���7�z=Q�FO�[(�bp@v�A�%�:�B"��^q�22�'Q�_6�A�����A��heF�%7��c%9/�Y6��\q$�
H���ۤO��ʦV�oV�2�#�]X~�a�gb���Ԯ|�"�ݻ�|-L��ɛ�"
+_~�k���i��h�%��j��a)��)轒�Nq|Δx��i���8���;�����߬
n?��L�ۅ�A�ǔ�!�9�HD��>���T^�4��Nz�[k>�\�/H�(٩�7��B֙A[V�Ɇ<ǔ��%��U���$�9A'|���e�*~Ea�0��!����Ji��P����G�a�/4��ETT�9��[�?f�b"�Z���oK�5U�]�е"׉4SX�'�p��]�����k�ߙ
��BFGlR�C��p����{�d�{��0)�f��HI��(�����f�d��$���X��)�XU!E�%�xo�0����������C�JP�-�Y���y�ő��k-�)���{znX��>��@�i�"v����ulpI4�嵣����:����m�+N �i`�@�����DH��h!_���a�j�kۦ>-�}9[���i-�=,�wΐ(��k��f0�����}�PPilp���@o.��$�;	��!3#�hq�[q�d�Buo���n�.������T"��Z�X����/zОD���O��@>��=GP#�ql�`�����D���F�C �Xe�Z�m�I�_VF']{��a�
����#b$�u��
�#1�@w�M��裏U7Q�܁�v-PN%�MDN����5ʼ�/	��<o�T1c��v�-!Փ�j���mӮ��%Z�\��	�'�T :��;��n�N�kB۝86J�1�g��;v��K�2y�����Dz�fK>9�]�tO[]d�d�}�݀D�AaZP�9�*�+��%��Q*��eŅ�0�~�J'Xtן#ٖ�"Fh��eH4鿯djIǟ��$m-$�5m�U�Q3,�nRs_�1�}���.����k��\M�-�*{p�˭��� NQ �����z�c�.wb�?�����#��v��?r��3��ڛ�`���D����&����p��W���{�ҳ�Ô�w�uW�m,/���D�����Q0�#�cg����z�p�<oz�%��I��M�NDT�N�n=�����|���k�r4v��	��@��NA�iXCԟ��ݎ=32�B��^4BJ�I�,Q��~�̘�f8'Y%<Ñ�;ՅM��W��K;�t�V-]2�|c;v�x���p�*��3K>��OG�#�}�[�����^V�EQF��9��@D�!��@�㰯��:�1�<������Y7��fY��*�g�:<�D����Bj�@��])�Y�ц<*s8Q�G�l)���`���\�I���Ѡ���Ye�ʳw=�6w�:E��m�k����T�;b����a�`y�lDj�[Ngw/��Hj)Z�n�#�tk����:�9���R�'j3#Lo�hU;�3��=��'y�)��z�2��8."6rǴ�yE�E��Tg<�����Y��I6]��"��*��I!̍ʌ���-�O�"�H�)�l:��o��E$�}�a��r������|�<��u�imc ��д<�,JN�Dc���;dUU���D���[jd}��y��+.�t0tl��uF���ݢ�;8j�1�3��ˬ��V��`7,�8��_��`�#}�i��{rW�	�-]�����/�T3�T��(�]�Ɉ�+�,��Di��@�҃#���� 4�*܀X�k��N_9��U�H!9��{��d���[��7�8��ۉ���A����F])��K�!�� ��I#[�d5a�j}��3)�J������ka�@��(�]	O�x60��N������Lqo|�
N��ROhq��g���p`�3n\X2�ě�RU@�"�A��.ZM$qhUՍX�H{4�2A��zo��=5~M�8F���_,:ۥw����k���6���~=,�;���.MPɑ@b	�9�����c� FX ��g�Js���С�����ο���#����!R>)�����nu����,��9�,,!��zwQ�'՞*ܬ���R��s����A��$�ɶ�3
(G}�Ş�&l�t����k�?��ul�9�1���O=dGQ�J�Gn��Y��O�(�-p0<�;�x�j�%+<�CBَ[4#�K�9yA�d��v����`�h%R�򰷖8��fv��n<�����\�G@�9U���v�I�)�g.x�5|���ŉ/|DnGY]�Z(t��������]�h�ӶT�ѷU�|Tm�������pЍ�'a�9fU �6��D{7B���r�-/W
솊�E�Ov�Ĥ~�nYg₠@�u��<ks�ˉ�b(�^pd
en#l��j�����:��m��ZA�������K;���� ��4�{K����ݾq����ש�%&�|�P*<�H����]ƀ�XaiWg���r�E�[cJĠ���R���0ޙ)#o^���F��;���i�S���HT\���Ә�&Y���țS�7?�����ro�@@I�o�b�33y �@!
�-k>jK�}���,�)���<��C#�g�j��!�G^}{Z#�E��s.[��B%b!��CP/�	[�U��_�ի�턃�u雱�O�c��㿐{w���q��i��~l�`�`)�J��9B[X�v'��%��ՊS��p8�̀բ	*"��zdFv�Gst�i�]-!��ֺ�p�G�H�գo]f�BbO[��.}2@
ب����G���[c�rՄ`��n'���S�*a��>����8�ΣB��g�L��=fsI�U��|�~�m0)7G�B���曌�|�hŐ.v�4�{t�5�t�\�~R_�����h�lNJ�$Mv+U.u�'��;�[)��B�&�ND��SJ�ՓZ��D��4�hK*��j<
q����=o�j�q%�&`��C�j+�5U�
�U�z��1z|d���B�-��$'�$S�&�{7����_Z���_���`ķ������k?z��F�Q��lk��5��u��@*��d�<p�:���}pg߿zvDul���N1m��	����7�˹�*ac�/P�Q�k:��yj;���o�f�/1t�"��4�)	��hC�gd��\ye��(T�$�ܤ����p���)����-K��f�]M�o�KU�"��3��q)��T���@/6�0�c��AD=+�]�p'n���q?9��L���G����w(�6}3U�n�p�P�"J}� ���<����X�oIw�����"�]f��X����N�oC@�ӎ��J/;�gx�d
K5ow��S��&�S�u*�L�
�*��d9N��;�B���x	�	����Y!��Xm���,��h�0�#�K���5_o�����c=d@����aJo�?�%��=d�}�򩝼̭R�G��*)�?��-X�������Q�d8�	ta�柔7R�x�La�/����Q�>��3Fx�<����өJ�<mzXr�o������#m���[ !����:G�WJ�;��)SB3}q"��>�|����ΈA6z���(>Ɠ�,�tw!r�98�(�����ʦ���Eno��=m�B(lsPm�G�G��m3�UF���P��� E�4�ڲ���UJ4��ǁNŬ�_ۇ��j�C�P+�+c����r��o$J��O���ݤ��v��߷��[�7�^�L�����8k���I��;��J�T�n�؂�b�4�Q4��R��	\Z��7Ese
?�	?��=g�7���?�FO9��+�{�T�2Z�g�{+��K�����}R3���yl;sCu��'�DP�wV���S;A�|CN�j6��b�@�ͩ���N�N}�S.�4r�L�^�߭���k�^ҝ� �>�����gM�[�'���UF��:=Q����r���m�ԡs
I�R&3�=��T�f��Cw�D����o����Ν��z^�_�!`���W`������L��e(�)���[ ����k���@Ubt}�?Jթ���;�T�,.4�9�ρu�D�#�t[>�� >�2 7�~Q�w��I+Fx\�D���n�'�o{���9}���]�R;��#����0z���S�]m.nO�n��'��2V�	s�r�?-&�X�^X��1*-I�xD�2?'Ҋ��rB�W�=P��@hrK�4cb�9�Z����`��
G��p��bX��AR�	U��e|�њś��^~-��=��m3ok�ʆ��.E�ܢ��):X�)����<��7c����I����NTX�6wVnYgn����}�C>(nq����[w��H�%��NCĻ"R"b�LW�K���+$W2�}v|��
p���pj:�h���l��"\�D�!�hLގ����<؊27M��bsD��F0����	� ���z�IZ�Zf�}<؞0&⿿���4�YOkJ���k��Q��Í������JB�g��3�f�0`Y��m�b�H�L<A�������h��2,�-��5�p%!���B��'�GM�e{��y@_r�b� ��B]�M�r����h5��p�^�-�hȥ4�e�Oj�/���;�A��2j?ә��t5���%��&o�4�]�RU�#uQgIP?��2�;d��`�T��/�<��{FWA��ͯ�6 ��q����&�����2z:���!�W�O �}i]ɑ��Hf��f}�V�b� y����y��1�?������)�pI��I))Drp�n�.gR �Sι �Sz8�K�F��2��8ȍ>���g�'�c}��7C��X�_D�Xk�}�Ӷ[m?�s-��[�7��N�p솅}r_Z�:��J����`~����H~�[�*�9�V��F��'�q�j����#�Y�E�+����7�+͑�j6�U4V)F�
\q�'�`����1����J�!N�Y�xGP"yZ5�2+_���� 3.����0��o�-��N:���AQH��E�He��a���̋T���^�,Ȧ�*��( 7K���F���(�úUx(�4��J,��}������j���Q��,(ZrM�m{���"I��%��byp��ʏq ܎`@E�@���f۞@�~�E����;Vq(�H*̄&CQ�����m���\0���o��Ә��BH|~kҡ�Z�_��fS��'���L��W|��s��	F�A�Xp��&�P��9:{�t΢��1�l&��M�Wx4V�p�9u���2��@:��4�|a>�	-P/�0(L�>�FU.x�\��>H�:���g���k��gpZ�5�0[&�v�U���[2{���}и�j;}�%g@6#�S����G�Ļ������$�2�=�^ڌ[1D��)Nx�5PpW<��|w�+x�NU�- ԑ���wlS�����Ϡ��N����z�@����VhH2J�sm��%'-�mH��;�$O�nT�_����0Ո�d�N+:���%uxiu]�*��J���F�!*>87�gg�XP��x�G���0��Ҁ䠱��Y�B�]�hť���S�;�n����ݞ���%H��O
~�59z�p=`L�>8 ��)�6��%<�k*t�]�����8�캏�gt�\.(eG�j>S����Uݺ�:1Af������<x�Z���L>�$�(���k�7�!z�����=)7�������"+W���!#������Ym�M��΅Ľ�߶��,#I�%��s���ţF�u�IL/Q���0w�R��8&��x|�z���̣���eX�Rㅄ�~3"�6I�rqL�$ �T�T�}h}A[�~]z�؏� ��<���宊�I���H�)Wu�f���ȟ=L���T�v]j��"˛#�ˤ�����̯U��n�<���C�~k���x(�
�Hf:D`f}��@���i�	#/���9�UQ��;�wL�g���E2�\_(&p�`�L�/ urM|?�5�1��6���G�/��"AJ ��n��d�r�)���V��f<���xknW9�P�I��JS]�!�� Ze���A*����E����&��mJ�S�)�?��95�Y�<�/瞧��z4����
P�_N%|"8*7��p9��c�@5cz+3�t��p�	(�����ƹ���[�K�/�IQ��L�eh��؟���p�q=T.���r�5�����WBdp��H�q�,�P��	�J��C?9}45��M`-�
��@�C���AO.��}�IO��SN�)>�9����Y���sz�@�%������ ;�ƥ+�&�yw�i��~r��p!��	�TId&�W��>,zÈ���i����Ŏ��q�^%FH-V�G���Sׂ����]]�L������n��H���ʕ�)�w0��P��ޡ5����n�^�"�1F_�P���X�2����U?�	1��[㺶��f�=���L�$�4L;�PȐ?�����+ہ��E�D�c�%qX�I�Z.���;M�����l~慓���5R3S��
�q���8u���h4�`ѫQI���@��9����Tz�M��<BT�,��g����|������u�mk��������f��_4�D9����Pq���9q��y���G��J
�A��f:!�j���д�Hj85�6��~�6h�q�$��3Ĳv�J�Z�'+�6٦䊉I�����"��5>��z�-���/|G�:�A l��y��EKG~����`G]���X�����^�Zg�z�,']N@�^���ITכ��ڛ�	�ɷ����ٚ?�.��i�'�4����l�XĿ��g�D�J!>&�M��<�o�Y�"Q�/m��
vyڮ�|������9Y��{��V
���a����v�"
��8��d;�����!u�
Zs��2�O����"�ܔ#�NQ�b���z=ۧx�����u�����I{� �A�؟�Ԡ�:�NP�o�Q�}?l��|<H��}d:L�*E��L�>`������S�y��M����R����7��������U۠]�oT���|̯���,m�2灨���2]��¼��T�e�F�b��:Y�@j�*G �,�D:��k�Ǹ��&�0��+>-T����(�F 6D��4s��g����o�׌��Vn0�xA��P��!��m� �Ę�Oy;��vg�'�M�\e��	F�C��^��tN�9�}[�h����[1 �	�r��Ӽ��[��r�me�M��?9��� K�\^�P�@rL];'nH���f�����~;��U�q����L<�Qz���9�+9��?f�&�y�}��E��>� [�q�����ܝE-�k��,�z>�ٴ�Z?PG*��B���u\�(c�m�b��J'��l�iw!ԅC-
<>SR��D���}Q�L���a�qZ�p�����`�9Ӝ��s�NB�Ư{ɀo�/�l�S�����>(V�K�*�<kM�!$$�^�������ֳS�d;c^{|g���ў���'S��h@�1�J���"�b���)S����J���+m�0��
�W��I:p��Lk�b_�w�(b&��@�ϲ{�v
 �����` ��C�S�GN�b�~9��qz5�0�kyb��q�k�^�"�&���ߍF��k�� �o#+�l��|O�p؁n�rS0&Gp���H�q�Dٛ8FC��/����Al�J]g���5û����;m����"�I���h���@��E`�96,$��؜`Z���[�2\ukK��Y�����h7�@jNF  @Qq�U�-�㞳u�2	��4�}��җ��4K�?��#�={`<��ŁȀ|��3.C�lk��BDw����]1C@d�d�{��XC���z��XA�:�B�������B��!��{^����ھd��M����C���y~g��+
��m�S���=TE4�|�F� ����й����x��`�a#���������v����.�=�x�h��SZh�v;�˳7��5D&�X ���G(����f� �#�G.Kďa�-x�"���9��=�}J1��d~���=am��p�G��l�Y���e���O�3xĞd��%L�˲Lm��1���� !�s��w��yQU7�<�A��QL��@��mer�,�ݐ{�%���r
�ql{�v �����9�9ե~�f�!D���� �Xی~�E��	�EV$���q��
�r�g���!W/o}�as�'�Ŋv5T�� �$����Z��9b�ch�����`^s�&� W��YT�� ]vB�0ٻ�����d67����v�A?��t�(^<��9v;	�.����s�'�,42��O���Ђ��ʺ��JRQ��EW�vB�F�QihH�$7�>�{?���v`�{~���\�{��Pz��9$��Ezq�1�p�D���� [>�Q�Æ����� +��ib�EO��:<~��W�Fy��l�{)le�5���K���+�xO8૝�<���3�n�?D�m�x��m�e�.�n�̞ku��`�����#�i�~:�k���C޲�ȸ�����D�`��~�b֗0 ����� ��� M��H,1�R1B
70W�\Se�w+�G� �#�����S���K�{d�����_�D���d���P�ԉ�\> �7ܾ���\��ĉ��c8�Uv�U��h6�ÆB�<b�ϑ����!#!6H��d��������ֶ"���4��P�>�Y�����e֌ωok�pM�.jβ~��P�s"�U��	:e��5�BN�Ȉ��c�@�Ȏ* �)�V |�~k!�=�V���g�0�5@�d�����U�����d��'s���bh�u2҄�����*�!��m�3E��ʸ����Bs�1fz�2��Ι��
>�r`1gs�7vC�L4��#	r^x���1�ہ�@?;,�s�L���g4J�x2�h=� �qxk������*6M�bO��v�Y����M�KZ2QcKza�T��N����C	��Y���Q�;�a�>_�����LT\	�RZ�g��J�9/ڭ�t��qq�\���_��2���WbT�l{5oI7�E���*�����j�K/7{�\�V���s�!�������eH}w�H
�Lʣ�ɻ������DU�)A#D�V�.3�V��u�=��MG.U�h�J��5�E!�6�5�e����ޜ�畷��C�O�#�44((p�-k.;����G:�x0��K�>���_�,�j���G�2�9!��Ӡ�8��isjì�
�*���e��"d>Hh"W�!>�m�>u����j��t;;<�D�R7z��(�������7P�<��9]��̟hwX١{�c8k{0�+�_VݷH�>�ޚUԬ�Yt�ôE�s`�[�c��^pu�C�����cJ�Q���lˋ#'td��+U�9���}��4~�L�4dzuyMk��T��z!�[�v!���aJ�`��*	�"�7B+&�����H��2���F�?�Cwc��PR6Oq��0��}\�{�@q^%(������?A�Qae���u"B 6i��5s#���6N���r��T ���aR�_^��3��7j3��
w;w��?W�
�ä\�[}}�^f��9Z0��O�9�c~1�/�"���e�{�N6K�*x1��>{|]� ��SggM�i� 䘛�,x�;~�=]�~���@�Ġ\�k��1��c���`B7-Ź����\�*����Мr;-����T$H��p��<��TPe٤���D��T��F*��S���V����:��}`����v"h�����q˙���+���K�@F1���
,�f�a.�9��9XY�2��崭-n*y$�Ya܊�њy\�3��DmPh˼aKm����f �)�(y��.N��舢sN���[=2E���'�ȶӶ�j���2 Įݪ斲���&P]U� ����uY��[�f>�o���&y�ܸ��3o��� ��A����a��R��d#Z����a(2�Q��^��S4I�Ox�� ;�E�z�5�rOw�Hs֡(������I�W�.	���[~�K�]�7 =ˋ�c0@��PT�4���>��m����9��	�~eV=ȟ��=�_�3�m�0*��3�����R�d���a���џ:`�"�4�vk@���E]�m�j����f�xH�Ҟ?��
��bZ	����k#-�\��xS�B?�`�f"���T�Q���7���\@����n����o��n0�
q��U�5E��^H�n�^W���{p��5���<N�ߑS��6E@�R��|X�oa��l⿡3�t�ƙ�h�8�����ݾ���5�˥i�#����^pݫ2D�!�F1�o�`'����jac��&�%u:Ɛ��k?蚮�U2&$��ͼ�.)ύ%_�u�=W�+�\�ؿ��7]S�[���E�u��Bi�+�DȒ0CA�Au@�$c��|�`�^�)
�Y���GS�<û�7����2I�V��o�<���'�]�V����6�'2�B�?�vXe"�
�0y?�fb���)�v�����]Es���[�lnGz!�Y�Jj �-A��~k�Z<z'㨓��9_$�x�4����	�t3Q�z�q��(\�fC����u��N���˛�~1rI;�mh�#Qh���7���߾Y4�~�j����#s^VR �Y�x�5,7�P�eH��t�^c�no�Q�%��o�