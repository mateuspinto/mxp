XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���j0�ؠ��~(�����h�0���a/>aX�4�<o]-#��7:��g�>bI:8�n!*ˋQ��ѝ� �-i,����OÅ�;ZHf�l�A�|DQ��Ef�U:M�zʋ��CE�{K�Z���2B�� k+��x�h�}���jF�$o6�
�6�&sǍ��*��[w�&�TN���Q��A��  ����8�/�<���^�1�,�|r��k���%I��ꐯ
�<���=n2���q��+p��o����O���Bo)���d!X��3-1f��$́�Z�ۆx`�`nщfII����Ha����\Ch�{	w��.Q�\q4��~��ٽ��XĘ�Me'S��j�0��+�
d"qw� ��9f�{pX-L�z�Sɀ�AO��$+���'F�����
���)�ʣ�V�wBM���b�(s!?�_cq����h� ;F����c������4���G^j�Qư#ؑS�\X'��.�K�V/;^Ԋ�`Ki5�!d�ٹլ]*��qKt��ԹV?��qrP���Rd�Q-��=�ێ�U{�dNY�۪1Vw��e���AB�C��b�V�kP��'d��a���~��S�>�6����$�᪂�5��刋�}��7�8�x�\�^$�-ȵ�x�ٶC[�%\�32�䌭g0L��6(_Y�mH�T�����3	�i:�2�����Ĉ̹]ɗB�=��R&�g�����!���=c�X㏷�^��Ӂ&�]����L�7������R�-]�9ԄFG�VXlxVHYEB     400     220�-����Z
���`;�	)�.Xj�K�4c]t�B:��)��h���XjQ�qs3zlde��Z�L� �AS$����[�{ҥ�,k)h��\D�w������������J�L���|U�<]K� Ӗ���A��'�=���4W+����Cȩ�|���t�Ϯ��f���
�t|��О���4P��
�~Y,8]j�p�b1\/�P��-C8]_��P�0�L>Yz!DFW����2^���A�LH�#��[�o����0Vl&hey�Q'��c��vҽ�SX+�uFi}]X1(�#T#��A�1=A8u�˷y]3'�S)՟���m��V��yK�� ����)X!�L�cj�Up �l��(��*�<�4㣢�^�����9U_� �6"h�$����j~ҽD�Jbyʫ�B����Ɲ`[
�2�T%%�/@���{T����8L�XE��{�)[c������fC(�iH�ė��l�BL3;̶C.�JS���V9�O��KZ:�^�V�G���.��#�K.���FXlxVHYEB     400      d0���cB����j"�[�E��I�։��e�"-O�y�qc^���ϩ�p ��qacW��#_�a��Tp$d�GQ�T��`d�¦�W��,hp8(�kNt�'l.7`�e�|t�+�7P��D���?F�U��']���0)v\���Z�����K ���?�k�mL0n�e����U!n���T�&g�2a��gaI���f��˺��"XlxVHYEB     400      c0Y����s�����?���︆�U=�b�~�DGw�M�_㝖�%ͅ��q�g�E�X4pN(4�oE��Ψ�W��b+Zr?*Z��_�Y,��-�3�X�]ae�<��`��A���_ ���M�>��!��cs��t�f�NP�Ym	"g�)D�j8�#�"'Q�Il1�}��D杷gr���I�Rb����3mXlxVHYEB     400      c0��٭�%ɈbA�����2���Ɋ������O�?�y*�������NT�#I��	p ×-sA�?|fAL������A�ʥ������p��'��T��U�_�Z8�b���\��9X��l�j��,�F'����Ӵ@�_�9���z�p��-�Ee�}Rg�0�6��/�9��d��փ���.�=ߊ�#3D����XlxVHYEB     400      d0Q,�J�!{��s\Ae$� �c!H2[Ř&�˘���1�1Lp�յ�;���$A�HB@�D9{<�l���ȠLk��գ��O��� �Rk/���RP��X"W_�j��{�p�7����m����\Le�G<�-�fx�GB*i�]r\�+H<���nq@�ք�[`�M�����	T��#��G��Mg%b��@�O	�XlxVHYEB     400      d0�e��P�^+�W4�nt~����E��;�ߧ�L��<s��v�C#=���ui-���+���/(�r��.��p~��xƶ- �.�.�*�����Rb�CO4/�з��~:Ⱥgk���06s��G�O^4^��fx����
e����L�ޣ��n�����A?� �!����~�b�?T&ʃ���Yն�����0��:��]H�$���<gs�XlxVHYEB     400      d0ς��w9�(M@rX�DW�� �JV�+�}ܜ�9���`�5cKyh{+ +1;-g��R�s�Sꂭo;M�=����A,��g#�m[�z��f0��7)����[����y�F�� jECVL����Q�<Ib�<�ѐ���-*#�Ԋ��C񤒊��	
� I;�u2E{�X�[,�J�^~����� ]�jэB`�B�kXlxVHYEB     400     170�(��!�M��K(��>P���:ge��PӸ�M�1��Y���l�ٵQ��Z$�~��㿓X��ҭ�5����e�:r�Oσ}�6�P6��N1�v�\��Z���n/EZH�|� �K�����p'��'����;0�d}��v~���i95oGmgvXe�KW�
�&���a�Vl�pO��m���YF�[�Fm����O�Z���Fތ6���G6~NmLp{3�<��@�k�1�Z��)zA\:F^l��HJ�&����W�[�>�%#BCvKK�D�J�T�2nm�ւ?N����5b͕ߕ���m����d���8~��ŝ�ڝ����LE�+{.�x>5`)
�����k�
	������XlxVHYEB     400     140ZO�Ю�>��U�ŏҀ�4F{�i	�K�B=���a��+9W�m>ZBu��{��3�Io4�齉8��.)U�u��逵u��Up�a����xG9�p-R1�Cr��z���FYʚYRԵ�ORr�?:V^�פ�_K���UtN��*X�j���(h�Zs��������viEb/���FL�|˔�����J17�<�I��z���?Eee���8�b���%Sת(w�F,�d���W}vtthzO~���r�6����H�#&o/F�ט��-!���r����	�;�S���pO�I��l��Y�Ab �
%8*�oXlxVHYEB     400      f0�j�[7�U��̥W3�֥'�"H����?8��ԥ�1�{��u�����l՛��~��d���B1�zr�v	BpJ0'Z�z�]����y���b�z�^��	�b�P��P
�a��:��{zS���M��mZ�堜�2�t�!���~`K%J#���ެ7(�m�������3�A*o���YiU`#8d:�(��9��%o���Xl��i 
%����&'��!AIa&�@�I��ϼXlxVHYEB     400     100�#��m�����xB��"���J&�_���)Ώ�-(�&�Ow�`�����9nSZ�>�zg�A6�H��x�������S���=�(,�P����|��Z��~�ෞ��	���@��1�u�m����S~�Jlq��ŏj���B|���C�τ�l��4	�Z���/�52�e�'���\ǔE�����j-���v7��=y @�5<]����Ђ�]���W߽[���K-��cF,� T�]��:S1?����!�XlxVHYEB     400     110�Q�?��|��cΏ(�R�6u�K� �� �Rn��Mٯ�|3����Y��om���ؓ����±R��[��.t�H�oɤ��
��'�8c�lmjk���K�c��:�e���*D���<+)E�;dM��W�P���`�� '�!��A�������D��:���nӟ�`֠	&��RSHU�o����qR4's.�Kh�������C�����W�/���ڣS��B���/n��oE]K����g^������s�Ax>r���^b�:XlxVHYEB     400     110+���g��X���;�A_��%��Qt�-�>�M[K��¢�溞�v��WJ���eJ#�)�	�l�k��2�v�<���.o���w�۸��/�s�&�A�
���D�p�zIb���n�l��}�!�=Z�,g����������8X17Q�}O�o�Z)����&�і�!�ks��e_J�R�t3��{���g���
��)�`2Io�/�$ӠɝH%� T��]e��/h}(k4L`sEg���Q�: ��tF��箻襵9W�غMXlxVHYEB     400     130ce��\h.��N�16��/ �.=ZU���*����I@�����f� �b����M���Q��I(�֥%�����Dcn+�}VGT���Ѱ���F"�>���J��k\�k�?5T��3�ɿ���w#>H/:���Z�a�Y������Ad�W9�i���#���d~gŘm��"[B���Բx��Y.����Dq���M!3S�<��_a�NςŦW�4g¨+Nͱ���po-��~�m��Y�S�(
��D�:#m��[���hr�;�o^~q]��"Ӻ`��p`��XlxVHYEB     400     100:>���r�k�c�4���%�b�Ϸ�K�Q48�C��y��6�n.CfMx���k���j��7�,��3pY��kp.rL������뒜���h���˒P|�I�2�~v}��)���9��P�D2R�VД]�Z��87�Cq*|&�P]��IMTS��,�<HA'�+;�#W�Ma���=kd�|�E%GơLԂH�x�G�݃S��f�8�:��H;7�?Ǌ�3�U�͕� "��`�:?��a��XlxVHYEB     400     100�X3:���`6�F}�֫���|RN�P(�G3@}C6�]��^e�/�䘈�e�YD� ��귑kD ��gi��K��Ƙauym��R��/���=O6��_�[�t�L��@�L^�WV{��1@֚�Mx�BE�
ek�����$���O�έ�i��%a�9��T��v���Y���}1�eK��r��{����\1r1��`V����9N��_�nj?[�gpV4s0[���0����[��C�ʵ��XlxVHYEB     400     100�j�A4�ɬڀz����nPi��j���V�)CR��,O�l����Mj���Cu�д���T�_[��L���&�mr�CɆ#���cd��H
-���g�S0�,]).Ks�u]�K0V�^����{��1P�ʴ��+���$f�.ֶ��#?\j�Ķ���p���6���r�ll��F$��M� ��3`�v.�DQ���Ǭ�Y�N�%S'���)�� �Y��6���+L�����T�<�`�t'�/mO�F�XlxVHYEB     400     100f�L���t_k|���8�N2���l�{����R�)1}�����P5Mh��a_��j�vT���Zw6���WYP��>���0.�X��;���d�^�X���=����ߝ��%{�DF��y�n?O����+�j�W:�e�P���¼����}w��g�DP��{Ez
��LW��G��f�<��O<��15������f�~
�[~���@���uI5�u�3R�;�`�k=ɿ!|�]��e�NU̵wY���օ9XlxVHYEB     400     100M4l���H��̘��	,��C۪yC�C���k��A?����Մ����FH�P׻���Qr���Vz��k&�mYsH��I��������{�7="M~2d�~��NK��²JCH9rX%WF�,�E�nj(���H���}���j!���n���U��,6'�u/k�8�Sb��P�>��<`V��3�(@�JĦ3��=j��=�����-��ۛ������Z�
21�O|a�4tD-��}qP��2d4H|�XlxVHYEB     400     100�э��Ѝ�3��*����t['>�����Գ���dn��&�q��º��3��lG�!+W�s	�����{�8�_�wfE8��=k&�a�P�׈��rE����5�=���F~��BwئUB������X��q[������Z����:�J0MذӍҰ�K+YE,vA<���'t2��ґ�����2�A.��ku��X6��I�r�&�+|=pF��֓e��q�UM���eȡ�WE�ߖ#��-p]��:����XlxVHYEB     400     100"z�]�KR��Ti����6�i���wE�d�'�D0m�? w8�g�d��2c�/�w�N�k�����OU�'n`.�����C̘���M���+OWM�+�_�X���	�����2[*e���i���h����`�E�����ڿ6z���hi<�>�u�+�=�DP*�fv�9_a�Hw�,ma��u��Z{xkC��n3i�ߺ\NƩ�j6մ���Pe͠���`l!4Ձ;f�q���6�XlxVHYEB     400     100����=9�f=@O�]�n{�\1Ҁ=(I�����s�0w(@|p@db-���wi�H�u�k�N����V!Pԛ�.��U1F����*\��=%���HY�8��B3Vp�\����[˅1���8�;1�ϊS�vs���c��9�8ޭ��9�!���^�>��7�S�{�]D�w��J.�؁/�Y��Q�]*ru�@�j" !rrǝ���'
�ao6�\�ό�d>r�}����9��VhP��(H��PȒ��c�XlxVHYEB     400     100�gV�ȋ�x��^N���_bh�����c��1��R)��>��PJ�R}��+�?�F�k����g�w7%��w������Tqm7Y��=�g�L�T�[�07)՛���EXh��='I`)ɲ���I���\��^g����9y��[e��ld�YA%�xD��_��:j������%RDY���W�W^�ڮ�/჉�R��>+�nX|�5����&ǲ!*��-�a��@�z��䇈�!�Ac��y5p���+TXlxVHYEB     400     100��l���	M�-��/��3S�}J4��A�*9�1��`^LЉ���z�]5�# ��ka�nX9�Nw�	t���Y�?"<��2��^�E�k>��hfxo�.^A�JPr��Gq#�S1���g���`�j7?�G,c]��\:
�rݤE��t�-Ml+����4M�Y��ƒTI��:Rx?��d�Ƀn�����:v�w�)��c���
2c,#�2?־4ҹ����A�^���}�������p0[XlxVHYEB     400     100�5��,`!q��!���3�� �����a70�	��vy���(��^���,�3N�T��qf�+� a�6��Ϸ}Wv�?�_�v�"�h蒹�X��W ���,��@�$9��c��1	UØ�6�P<
/�����\�*�BDA�
��/O��hBX�� ������:��\�oq.3d����fz�.O�n�1?�M����ס��XI�l@	�t����G^YY
o.ݞ�p$#�X:Q�F�3�M�5=�v?��S/��XlxVHYEB     400     100g�ǘ��(��+��.��DR�_2�%�i�QF�]ە(F����zޛy�F~��4�BP3�GF)�an���o�K�8���=s��mӮ��qŔ� ,�^?��R����2��)q���ѵ�]��Y��?�6��7����%!�wV�����(3b
<a����(������0�|����7�԰}~���Ş�b"���1�&�<B������L�����#��9훡;��n=ԳKA�}���oji��#�e:)XlxVHYEB     400     100W��r���8�`Sf�73K��=8{� Ñ�pUڥp5�۷���eky"WNXeO�V��ˋA�b2�ߵ%d6��*9��{EbP@�%G%�a�F��m���Z|�)ĕ-橥��Ar%p��������=�`iJ9�fV!��[F�H�P?��Z���
���m�z��WB��tzLЂP���MP��'!䍼R��'����[i(.Y>��V[�?Sx.�����|˓b�_L��g3�!��%*e.RQ����ד�\��XlxVHYEB     400     100�IK���@g�!k��b�⍆R9��g�AS�&P�->�dׁ{����d��;8/����֋��P�")jk@ͻ,��(�o���j��v��,�k�lFB��,�~��mKD���E�<�I�Qt'���m�˾g�[�"0qR�|���̌g�c�<:C��.�Q*!��Js^s6�t+dE��⣭��N:1�ѻ�3{��/ };��E4aǼ��]Rʜ�`

���'�=k��6̼`����6�V# 
+�sQTmXlxVHYEB     400     1000^�����s�*%-~B��Y���z�K=�����6�,���=���p�f \-�.A`MH��be�N�����ډ���E�F�`�@�fn��x��w6G&��ՀM���X�󲉛6؝cX'pY���U�o#XSW�I�ܽ�EaړAJ��L�t�o�uU����琠��F�/�g����iN1[�D�ïeФ���:�S�'��T4`1�|Xj��;O��������E�!�5�~{ݰ,,��%f6kXlxVHYEB     400     170�!{�b
���]s��]�`SQK?ւ�*m�Қ��ZW�n�<�|h���J*\i��=�E��'����q͡��Oy�2V �Q%����I"1��t|2{�ō\���c�6H�H� ���ԓQ�㌆|I���"��7[4�?hYUɚ���u�a��	UժF	���p�9�գ���`���F��n⫬=�h����T7_�Z ���F߷���gt������������b��OK���Y{Fė��A�#����">g7l�	t��U�CK����2A��p�+��$��<AJ�Ü�����p��'i��IO�D#��R��t�%��S�!�a�G�l�}�>4>3�XlxVHYEB     400     100v*]�8�������V��;}#-w�^X�1�<��Y��UʙD��ݒAY	uw�:�1�]}˥�	�6�?Z-UC�f��tc���mƍL98x��!c��O|V�2^!L}3�o3�.E������@#��Ŕ3�z	�0���2����Ac�T�/<�D�ׅIXr�e"aw�i�A�~��$�_܁���`���J���𲮏a�:�B� �����|�:%��a�$tW0W�-}�/�MK���XlxVHYEB     400      c0r�W��|��-l�b��S�^F�:ߑ!�t�����Գ���?oB�����٥���9���>��~����+Q��+�	�;:���G�`]O�]v���<ҥ_��-S�mw��XD@�cX�/�ê{�ζ��TA׍I��Ɩr�#nA-w0b���yE"u��O͞��{� C���f~8�a"���XlxVHYEB     400      b0YqQ.)<[�z�f��,ՑVH���`��Q�7;Z�oe�L =����G=qD��s�±qxg�W�ed��<�{�vȆ\�x�Ԁ�ջ`_9�S&���(�4j1��m�7g�}&sfѾ�α��:��*`A������왡V~W���C}`#֎����;ܑe`��EpڐK���g�dk�XlxVHYEB     400      90�O��MΧr��u7�e���n�����n`�"pu��4m�b˲=�(�.>�����'������oAՒ�6�4��7���:zGI��6=<��rkf�`~������'�N!�o�Z�U)��햮 ^�d؞@$��ڽ�XlxVHYEB     400      90�M|h�p���zDY�*0�݌�>�>.韪�� �8*��5M����g�dxN�s[ k*p��V��b�]��.��/���l���+��i��������E�\�Z,��w���8U��t��iw�vWw��������jXlxVHYEB     400      90O�&W�j�Vv��b��m��X�GS:,,k� Q-��RRQ��|Q*�Yy6l9:+Ό�Y�^�f��z�n7����M��ƌ�c ���X��󅯵�;?8���D��-�v�򇻃*���pjʧ���pp�6���Cۆ=UV .�XlxVHYEB     400      90��t/~�� �� r$c�~�y1d��de�G;V#ş�ߗ�Qn�tHV ?���u��Q�d�f$��;m�>�2Gh���iʞ��E�#�A(X3�CR��F�v�g1^>�6}	e ��)�c,Ov�C��Й��s�P�W�XlxVHYEB     400      90a B���$�����-R)Ud�w�y�:�5����^#'G.9��_[�s���8�n糟�ʰ����>�/��%-�uj���LZ��o��b@��0��"6�½I�"MI�#�R"�H�8��Рa=�7n��1�a�CAF�2J���_����XlxVHYEB     400      d0�y��
�t_�"��s�GS� ڡXTѫ"��``�8D��̲�Bh`�X0�8'B�9;���@��B_ɭF*��"�O�����mU�?R��� ,S�G���A��E�\�;�R�f���CQ�BZ��z���օ�����P9]�K�C@&p�p��K�F�����std7�����[�W5(����i��\��P)߂�B? �IXlxVHYEB     400      e0�����+�	J�ʲ0D��_�$�Ɖ*ݐJ�Z۵n���li�U`o?�������'?�6����7����#�v8h7|�DoI�(<R�Eb�}�a����JF-�c����l^���(���82�����}��VAj��'SU��y%(��d-�{J��oP5+7��zO8��)|�������bƛ���߾�'k:���p�	�u����1���.�����͒0�#�XlxVHYEB     400     100=�VC�m���ڱG�M�2m�;Z�|�+��HS���BW��3l���t�V�r(�<�VTI������J��pc"�r�\��G�7�eD��ȕwI^�ߖ�'�Q�v���yQ2�oL��*l�q�Z{��vT�%��N�2�$Z���9�5I���點u�Qѹ��]�Ŧ�P"x0naS@˽RZ5��� �����GIV�u�gvy�V�8�b��[|��F��.>	�����J��Z�J"�X#{�N��T��W�XlxVHYEB     400     160QЎ3��r�:�z�V5.{��h����4x;�^.n'+*����|և����ٙ������ю���p��շ �!Q��V�]^;��e$��@I��ѬQ�a����@7?W!�����>��D�9�4њz^�r��K�#�n�V����ţ��xe�2'��f܏���0�iɿ���:߮�NJ\'E�%����t��+�?t"FV��HE���l�.0��Px'-{��J�Ql���$@��Ə6u�"/�~)��I�P��<`�	���񜎧��k]"��MA��������0�#���@+��,cY�iS�݃���K�����
��J�hDN>I>�}�%XlxVHYEB     400     160�0��d@Xw�-j����/���u<O���>�9Ů|6>�B�#�்L�v��$Qw�Y�-ms�W���8-4E�@�����ڇ�/������m��s2�%�|�Fo����9��>&|uH���8�Ql��`jM���J<�׳�,mꠄ�Agm�6��KA�
2.�P
��e��d�@O���f3~��d)Ҏ}	j/��xI)��\����{N�~�ln��`d?C�����w��h�A������3x^��]�����g(��Q�O@�1�,�'j#]OK�MH9����^�wXn���΋��W�����P�	���5r&�s����-h��7~�V�y��s�XlxVHYEB     400     140ygw
���D�$�LU0���{"t��#[���ed�GJt�"ɮ�O߇Gc./�?C����Vv��J�� &��:-�~y�����<cSI�,�6y'^��b�?}����@��S<���`H���.����k[���q��Io�\&Sf��K^�JQ�닫���.|�h+>"�[D��)H�.ߘ����e�dO��16�=h�?u�[�G�����CU�mB�h���{!��'�A��'ƀ~��z��Ֆ/[�0#��?�G���P��RsXW�d�X[OE�t�A�{���uWU@�9PQ�%|�X��E�l@XlxVHYEB     400     170I9���!�{_ni�8a�Q�/�
ƒRI-<9�O`
x�dqW��V9WBT�lD]T�(��#�m���w_Mv����⇎�8�3�[���׋z��}h�+3�-t�ܾ�ä�����'T��(��O�p9�KR��������-���v�v��8|J0@b}CB�xx�9' u߇�6M�ּ�F�����5� a�..�=[���Pu+�FN��ma=��}.YFZ���Zv��}�y�(q{�b�5ET#)��dNVJ
u�4e�`�#�tq�5���.���)</�Ue�- D.qk]"6ʉEG��S�b������HKʢ~�,aku@��ק6�I��r%��,R���I�Rd7^�{k���XlxVHYEB     400     150V�9	�w�E�iE �� *v?jSE��DLȓ{��п9��99k+I:�G��Jc��H��Z�+t�Gi��)��$����=���uJ��K|H� �;NIQ2��dy_4���%.K��"�D��&����kM��'g��f��9�pX��[������kױ��1Z�MyV�U����#�2m�������e��Ï���kg`֑��<	�3�(���>|se}n8,W��oa��j�[W7����G�laQu�I��#3������h�5��
?�͉�Ăa����9�� t�ҟ]!C��sv+�H4O���뇭P[S�C\����#�����*�b��T�XlxVHYEB     400     190L�l�sq1�
�
j�H�2���B>�RA!�,��hNC(@{ǧ,���_�^�l2��٢�J�7U����1g�W��������U��� 9.Q�S՘<m�kuB�A�yG�RW�U�I�V��ϑ��,E�����q�ڝZ��[��$Os�>���S?�M�.�?`�zI#����[Rz0�x�$"���%�9T_�e��H�5�L��"Q5I����~�4"�M�E���l+�GЏ�w���`��͗����`WR_��T�C���^�qW9Dxu��}��Lg�fX��y����{�~��;�D��P[X]栯��Շվ
9F�bײ4��@�|�7&�E��T<��bı���ZQ���*��.��jᎀ���c������>{�X�#.#~�{WXlxVHYEB     400     150��8�0�L������z���_$@>���kkUL�P�>���8�j��.1���7]P�4���]6uVr��:,�M1��?������ـ폼jwr�"����}ܘ9D�0�V��-F�I�:�9��}�M�v�����<|Y3e���@������tVn��;����*���{>7j���0�؏�r�O����V����n�V�# �~��{y�����L��
n���r����Kl�x�^j?��y6u��n'pK����f��W䩅E�(mj�JLg�Y���t��<�;���S�O�� S1Ȩ�܎o��u���4���H�-�v֓d�� #XlxVHYEB     400     100�J��A���ɖH&�%��n['޿���vp��ǒDi�\z���d��jT٥���'ۧR��¤�F��`*�#��K%Wh�WD���<:y0],�#g^��RƅR�:
]��;h��>=ϸ_��RcR��T8��՝�p��iԉ������*_�g� Ll��Ρ{����.���9��LR�=.�O�g&��ܞ��nA+��
u�UUȳv17��c���[�}���]Ԉ��Υ����������XlxVHYEB     400     1909���ˢ�*���1��g,�Y�gd��'��%��H����6cRb�%�jȝ��%R��
2���[����M���� �w�eO6�]��Ki`ݗ	���q���)	��Y�ۜ�TA�7����ƛ�)7E�����V�8E�ш3u�V��T�݆��VM�������p�zA��"nd"5��u�V6��u �-�v�a�>�����)���6�Z�N5z'�@���|����%#o���M/�^���)xаM�S,,Y� Cș�ul��x�׹����Y�`|􇚺��RLQ9L�������l�����Y���(#�ٳJ���;�N$͍���� "�� #n�On/E��)��:J�KL���Az����.-A@���ۙ<���%�a���j	C�پXlxVHYEB     400     140��
��>�)��ʏK��~�����Ow���v6W��S:��>^t�Ӷ�Ϩ��H�+h�=L�$ZK����QP�Px�.��⛜�Ked�+-��R�d N4u�'� �����%�<�j+e�qs4��<��� ͧ�˖���b�*B�=:���۰E� K)�D��ޛ�X>\A���+�_:�O�̑�J�%���Ř��~�8���g���p��[/l��p��Q�7���>���8�%��u�|e���o7�Y��ch!�6/b�,=���&.��Co�."m#?n�dV�(;<��7%�CR�3;B���;���, �H32�a�!�XlxVHYEB     400     150vVfs�P5,�j-+[B�ܐ�WB�u���L����	�ő�A�x�
�NE�������+�Z的>�V43�|�S-1��k�8�	=��g�V��;5Z>I��s�A!4��Z�<�Mg9Z��(tU�x\։��}�!  �Y~�ݬo����۲������R����c�F��ߤX�����7RZ���P� o���~-�5�P�0��9ř��e�ϖ���4��x���k��W��,���M���ݐ؉�����J*�1Y]�m�ն���&�o#c�R5��c?���^v��苧tH�zpJ�������� s�����>�J_3�^RC�� �jNk#�cjT���XlxVHYEB     400     110AԊnͰ �f��!���q�W��J���hF�#�����B�;�v�L��ple�ĩ�R9�l;Q�C�'�0�f�qG�3�EJQ��0�w��i5�񡊤q�p'����U�^4=0^	͒�W��'8
EB7�u�]2T�'�@r��,Y/���Z����gْ��e\8�A�c���=����Q�lO�hZ6fL�8�`,�{="N�{����ajP*t#<�d)���/��#G�/�B�u��"�v2�ژ����@��V��	�,=tXlxVHYEB     400     160
�;<"�ѵ�DoN�	H����G�Zl�V U��}gT[��l�<̢�8[�������nb��9�y�,���/�oճ�B���w�?~��~�,��k�qOJ;��NLe����R�0Y}�h_�mX��G3�)�A�.\u�!
�ga�;$�Bڂ�`8���F�aEhSs�T�G�8�|����mե��y�ф���Y�?�8@�Y��af{n5���ґ��9�W��ys��p%���TR��2��'�/+�J�ݑ���	HÞ��G[�wBZ�c��އ�����|/i����)4~uWd����F�|����-VU�ب��3�y���*�JK�ť�3�2-XlxVHYEB     400     160�o�'�tty�@���˼�}Ʉy��-	���B𡓋@E�{1�5��uf�����;�=�g&L���g��*2lyA����q�F�F�x�6p{.���Ek�"_�ԇ�O�3NvV��B]c�O��H��Kc�ޮ�+?�)��V��4��-�@�w���4�DS� a*J\���0�P�'��L�H���W�5�?��I6[�+�Q*�UʠW�J�"u���+ǒ�{jZ�I��L�4�w��nF(��'�2i:�}�ص䚊�ڳ�JD���3�ok�L7�vOr8?-��r��,\R�S��
�OƢ��N��֗����s� �:�K�NhĪjQ*2I�Y"`gd�{���Qo�\������XlxVHYEB     400     150�z_&��Ӟ��ʩ�,�´iZg�Bw�r��^Q�����#sy�+�i��O�jzh�M�bJ���6�����p�'��R�i燰T��4m��.��Nz)Z��p|X������?/�LR����mqT�j�^�c��=�����n��7ǿea<|�:�|
�ճ{g<db@�9�����r��y�mȲ�iÚ�UC!n��ڐ�\�+���m��2Zdg.�����l���IwRX�w��:���"���^��R�.o�<_+�U�hɝ�(����F��?IN��s)c��:���e�>*�Ea�b!�.�1��P��n��A��H	�;�`��%:�4XlxVHYEB     400     150'��x�H'�_0��%�{⫡�6p�B�G�s-9��lA'Y~��,�R���I��o��EF��pH�g���Ջ �=���S�3�gj<�2ܭ'��_��x5t$��]�b�,��΀ Ӊ,��)��b�I����A�9V�4���Oק��=;uh�Vg��W�B�{a:��i�F����,/�#�ڝ�"s%�X�9eW^N�����o�b[�q5�GR,,��+�6���N��&�M�v>C˩��!U�s=��a3`�M�ȸ}rs$a�����A��QGPv1������{y�<f2����|�TU�[\�1W�\.@��H�(C�"��iԴS\Կ$�D��XlxVHYEB     400      d0D�ީ�S�ڻt�	3�"5�����H��'��O��S>�b�Y1�pW�
lL��v���K��sH�F�\&e2� �6��;K+�W�����X��^���R9���w��=1'���ů��U�3�^��5@Ǟ.������Ԍ=��T7��H�T�hR��I��v-[�f��+��{���9|{b�G�7�ؕ�uxo���=9�XlxVHYEB     400      c0�Z����]���]��+c�=_(�1�=�!����:�)~���q��c��f�)nS4rb��֤�E�hC���[˕����:���T��y�$�Q0�
_�k�1�2�}�'q�A����*��] �X��t����e�2*�;�j{��#��C|�k��'�e�	����)�q4�ʃ�/[9D8�#��XlxVHYEB     400      c0ɷ]h?���Q.�}�TU�֚�0:�>�9*����89�־c}�A&Qv���|���v8gfz��*	����ǿ=�#�)���k��;����<΅}{t�d�W�%����b��Oy��H�X_��-_�!yL��8�,�����k�s4&�n�°&���Y�Z����;�o:��D�O=�U�e.�$��xXlxVHYEB     400      c0B��6�4�Gb�1Ih_�����a��Y��2^����,#�����
�|��ЕHW��N!z��L��1�]�)�w�qrIJo��E����UC6�>j��F��~ ��d�g��We�C8W$��,r�� ^R*.���H���6� Lƪ�`����6�aa!�Rt2�r׋~�ܜ���2��t��C��E@��XlxVHYEB     400     100����|�_���*��$x �k��G�^X�=��Q�(L��?�_�_�,��.ae�Q2�V�N2�!��̮��
d�◐��q4[��5�#h�E�$vX6#��W��A� ��.Z0�a��-��
sX�M�|@0I����o�'�CU��;Ƭˈ����:Z0� ��+P�QU7%��'kc��4οv+�4��B~��ɝ�b`����R@H��]	��(��ֺ�e�eX}S]���p�;����=��սXlxVHYEB     400      f0C�"���yMWm;K5�� i��5Ư�'sc��d�h�vo��-�+ة��~�Ǿ�'���~�m)s�F�2�@�_�S_���K�,����^�_I���_����l�֏i��a�3�
��n��Va�\^wo����<��5��\�B�
`1t#�sd:�8�"{�$'�7q�����/������Ĳ�K�?	��?��z'�O�/�d�=W4���|�8&'{���I|��rS�Air*�vXy~u�K@�'c�A,XlxVHYEB     400      f0������`�"��$	������gf�'���I��ͬ6�/��Ց�%�0���5�Q�����yݶ��@�M%<�V>x쉆[d�+P��;�K�!�����eC��|����'lD��|E
ts�t@�C������������+&aK�J+�E������-Yo�BQaX�W	~�b2{~��e�Jܳ���f��u𹦾߻�ķG�gPc�� �
a��\���l���k�<s��P�Ӿ?XlxVHYEB     400      f0&2� �P��FG�����PiA�	)UHrm�!V5�"���=~�]��x�b�'y6��G�*�?�Oz���	�@�98�8�P4�R��gg�pb�Q<��s��Ā$H�W�"�;桒J�X[��O;�(� ��3K�4�{��i.+3��N���S��`��NF�n��m�9G�[����l��y����Qj�ֵ��c��$�Kp��D�̰�w��?����l����U���X2��ck2�hX4ټ/XlxVHYEB     400      f0�F�ԀLѾ�s����󸾆[|���������u�]r9X�B~I&��c��lE���+�呪ZA�>E�8(�N�����9&��ť�OZW��G.ì�D��[�*�C�?�,�1����Ҟ�\�j+>��a��U��g����aUK�cQ~lxPL?&�w�޿�� ��K r�8���a�[��yM7E~ٶ[�[��~���T�� W�f�C�>��m�XlxVHYEB     400      f0�xW��m�8jIAZ Gk}�6�';~�X2���šFڣ���V᣽��.�0�eM�A��T�C)��9��E/����������"�#�K0v�=(�3�R�x
���t��G*�#a�A~�О]�/�֊��R
��A6� D����l�ZжR�l��bc {�d�*FG�놡��}VX�*���r�s���rm�f�5��qK����e��������ξ滝΢��,N�j�P�XlxVHYEB     400      e0,��SMx�[���C�ѿ��z,>D�l�Z�)����a7Ǥ��S��o�wT��j�U1��a����!Z�4`�%�+�����X&y=���%L���s���N&ސ�\�Ȅ�x��]"����3��㐭^!f���3x �d�x��^�<5���i�3mFo�q�3��p^�c���t�*�qC����Q>tJ�f�"s`b嵅/��7M�F'�6V.,�ƽbXlxVHYEB     400      f0_��G'���	�uhL�(сY�D��=�cK����ٗ5��	���!%�շɅ��>�Pt$[���P�l��[��򓢟�\��9
�4� :th���c��]��t&(	��j���I���_7B��	q`�K�����ޞ�;���FRE}�jL�Ks���PkP�r����Wo��(�;�lY��qX�'mI�<�?2�QKv�poӒ��q�����(�i�ch4$H�@2�e�n���XlxVHYEB     400     150�_�G�u��Q{��&���W*��TwM��lؖg\Eg#q���+����茨��8Sq�7��j���,û�rMV?U�mc� �u�y-�%���F�.-����
o��d����$����o�4��շf���xT BDDl�|�X�e2ji:�G�@�MEj���{��|w�@\�qF��2�?"�R:�15���$+]A�*Ձ^F�~4�Y�Uێ�>O۩�|��.ƻ-12��5(,��A��`[�Y��f(�TQ٬<^��M�ҵmJQ!�,}]j���[��㚼�ڎ��[ƹ`�i6z������ ���%�x��5��CB�a�[OI��XlxVHYEB     400     1a0�ԳY��4�N�
�f½A���H��l_W7�"'��SK,��3N�T4I� �NF��O}q"̓.�o[�8w��b()���g9��RC7<�1��EalC�5�1��>䨜 �_�5*_Ƙ���
g�S/3���L�_5D n�'9�Ѡ�!�;�W�Ifd�2���|'ck�Z�������lt�#�P�cw�.��S�R#9Xj�̮wtfR�&�u�Qb��(o��c�)~���n����@Ӻi�sM����)�p�YP�P<�<>S������3f\%�U��=�G�*����
#X�؅V ��W)42�C����J�zY��o��$������\r��U{.(��f�5@��x�(���ߐ4����s��#%�^*sՎYeRՖe2��J����tB
W�vִ�<߃R XlxVHYEB     400     150d[�������OG�~g�0}F�r%��O1�}Hh���@lP�!zЀ������Xf����iý�w.�q�S$*�< ��@��f	-�e �C���V�G:��yIS&�q�5�����8pm����p�{�s�Ē�|�:q�6���s|�>$��=[r�ȧ��I9yeU���i8&���� �����D�/)�_���m1S��-�����Hm-0�)ǱiB���;�)A��3�'���4YMIgK_����2b�䁝��Ҿ�P5���e������h�1�"���
�Zp*l� T�}1��ѶcE	���̋"�-9���*`����D ���E���XlxVHYEB     227      f0~�$����(�-ؠ�a9m���YIá_�~�5oc��V��F�g/Z���GuAM����&#=xv��a�RO3�]
�0��/z<
A��j�]kf�O�Ӌ�ar<%���a�4P2g�"���hJ�P_�ɓ�B �7S��h�\0��:���;XaH4o����l��t1�}���jS�������.O��*p��,�ݡm�'t�%�����,k�e���D�e��͞fכ��5+IT��é;w@��