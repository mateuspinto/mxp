XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���� ����*u������I�,�7�R2g4)���B<��5r'k�"�M��:17Ǩ���^x � ޫ�M#D��𩡸c���;
��n�n���8P|��-w:
�N v$�o?*i��M��Q-aI�����9]0��@�n�QLΊ,ަ�I�v`��>W]a���p{Cq�\�t�ե
XEJҠ���V��|�A��� ��^F6v��BR����v��3���e��lK�M�'?��]�c7���!X��0�*I}n>7�Pj�L������I�u�]�$Hr=���g{��˝`2�d��T��K����y�����J�I���^OUbK})��X�>F�/��V�A�C*e�I�M��C��}�źD��u65c�4����kU�s��Y�W��jQ�m���b������Gz~�'����k4�f]+Xd<��4�(�������c4>�/�	6� �q��1��Vid���r.!� 9c?�kKh�2xR����{��+�$Y�O~�BB�՛B�Ut<���e/;M�I�8c����mK�L֔��_� �����L���}����J�jT{���Ս+̜?��l��rd��[�΀�f��a�;��b�����n�G�W4�����W���ɻ��Hv���̒�;�����Gj�wQyiNW2���n&c�Tc�V����%FgX�enur���,A�Y�F�:=�m�m�J����T�j���so��Z��%����)#��F�����s!�Ds�cE���xmXlxVHYEB     400     190MKhf3$!<E
�ɶv�G���僋3������cN�=޴���ܳ���7���4�ϊR��@K�j�[������D;�T�(���0��E�IC���tuz
�������q�=�\4t��p��݊�8B=Z\�E���T�Y���'��l7R�e>,.�wͱ�������4ߓ��D@�IJ�sA��&-^���"u�m JR�f5��<lQG�%i"/����v��8��ߜ=�j��`��97&mb�k/��̊�"����!U4�z眗�n���ßL�^Y���`��~J�Y����	9d����(n����?jȽtQ����7���eg�:�@I�a�z�!���u�Ӡ���P�.������S� 75�l����k��YU-���;XlxVHYEB     400     1a0�c�^�͸�D ��ø��T2�~8w�H�����*{{�p�]V:�@�V	�rXU~�{�<z�JCW��#J�B�����5[���w�ǡ�����C�a�����6a6�介ex�2ݚ�� InB�Ud��Q#�t���n����N�x� ���}� p@0&6�,�i����7�%�S{`R}}k���h
Ѵy���>����7�N��[��n� Ȟu&���N,g46�PSG�ozW�H����K
���I�� 0	)�|}҇ic�T`\`�#�[�$n�E�K�/�A/+�ӆ)4)��e�X�Ȁ��[}�0��W^�Td��ix�_:ߦ,��{5��@�z������Y�CoX���B�U�9��SA��K��׫n�2P�I���k�o�nasA�NkMKp��xXlxVHYEB     400     130B/�f�eS[&Ȋe���V�lO��S*mO֝��T��I�V�i�~��2c'Ո@��x��:�-��^XE��0�6����sq��1Eh4f5��Ȍ:�@�@�f~�f��D$�#��4�w����0�S��*�����T$�����e�P����G��>�7�D�1yN���V�-*p��H�\dod���j~����y�}��^#�>"��<�ե8���C ���`/���}n��v<��!XT�O��t?0��r�Kc�-8ws+;�@��>�!$&�F��JU�á�D<��+���\%/��� [2XlxVHYEB     400     160˿.Iey&|�ؒ��1ۼ\��GS�#G��N\�����(�H[��������Q9%�����QFK�YVt)Y�b��r�<ol��#��b7H�doכ�i�*�/#8�7�*l�Z�Ҽǐ��Ys�^�P�?��r�k�ĭ�'��㷫�S�KGs|'!?�[�j�C�\�hN�}.�jfj�+��c���Ӱr!Um"�g�/'p�4��wύ�MĄZ�Cȧ�����4��_J����]ar��'�g��<�:z����^4ܙ"$�cw��lˁ�㻧�%:EWn�Ɛvԙ�w�,D�Bo��FUO_0K�����
~�gZ��+�;OЭl����g>�"�o���-mTǓ�ӉXlxVHYEB      3a      40�p!�o�*��y�f\G4rَT�/���ߩ�ɕ�j�c�i�E����_=����̷�+���Ө�