XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���W�.<����ؿV�9������Q��ʍ;F�e���ń��h�ɥ���¢�x��-=��C2i0ТR;R%R���K[jJ�D�iw�B�v�H������G�Р��AC:�+^�5sE�GaJ�A���}F�[�ELф�f=�g��&�����c�gk	����x������*.6��Ķ�(�?�����)B�r�ϕ���s�K���9�n�t���ą F�!A*�^��5��ƽ��F�m-���C��0�_0�i%�n�н{��i�ň��`�G���觺��/.�u���?��)yg����w�j�ɍ��2%x��|nB;�R]�]P�s�=��� �'��	�ϐ��ECQ�+J���Y����	��٧�#�{e��}�	_�!��a��.L�2Y$�`�,��3�mQ	�/�
_�TY:Z�Z���������`K���J����t���RMI�bRF_�P�)�#r�~=|5�(p¢X#Cj�]�k���jl_Ԇ�fZ�:��3�T,�����*?TO�d��U.pY��8��wۖ��P���p��#(v��e
Hȧ�`B����ۄ��#z38#��R,� �F	 �)!����ޣQ���"~��!��e�'q�[��2GXB��c����p�@`���(�=��CL�)�u��z1���:i�b}�s��39bx��_��î�~$f�9.���&���	�̴�GN�+��j�u�#�c(uYwg\�s�����_�^��^�I��+�{Lv)XlxVHYEB     400     220�I���8�"�����]^�ʃ�ָ����YN:�g;��G��0|�ٻ8�6g�qs �ͳ��g����3 �`MwBꍙq��g6Ф_fq[�~�;ÛooQj�SG��kM۸��,8��ۡC3�L&t���YcC��á�Uo�H�n ��b2r���]ݭ �Z$
�Ӗ�5�b�i���L7R�jEx|�+�8p��G�vA�!�I�+�e�4L����
u�_�pN�.�qw��s��Li�Q�Hz�^�A�.�lz�+�s�7'د�����k �@��l�k#��O����98}������sk����9�A��'��7IO��s\o�k�~�������m(����׳�K%����`u����>�҈�0�@��(�U�&�4�eUhs��䨣N�J����8� l�d�Nq�J�Y_Jl;Vq~ƽ:�\1&;9�c�,r�����[ڼq,/�B˅]BI~��d��x���r��\Ԭ��e�㴗�S��%7 ����42x���^2r��N�%<�X'q6��XlxVHYEB     400      f0���	K -��2�)VN'#՘������	A�C�
��ac��hP1s{Rg;赀&(
�Ize@�-Q��Z���؇I��+?�T�H�_a��nχ��6�JX��}V����n�j3L�r���=�)T0��lro>�Ʉ�N3n׿�ka�e�����f$��X�t��1���l����H�]c}��|7���L���C�J�y�_Ļ�Oa�/jsT����u;��,Cj��XlxVHYEB     400      d0��AU�q�q��[�� �2�D*$X!7�&�ϩ�O�</g7́���#��3�#�
l�������ʰ����$ү���>�6	��0���f�[��ؗ�Y�r�����/��u*��RS�0��+�4wM�E��Y�p��=$"���P�/�ύ�D�luR��z�8d֒*�F��F�OÄ�(�$��K&x��/XE�B��uf��XlxVHYEB     400      d0h����׾]5}`��Ib���7]��|+^&��6a�T�w�������	<���7/�:
�0���V��Zg��r;9��lX�S�i��Ʌ��J���.�5�9q��Dk!A�ĸ;$��N�9�s��S��ǜ£��-��ޙ<>B$V_j��Su']!�B��^۸�'+{?�mZ�;;��1+�~nf��
���~XlxVHYEB     400      d0�1�؇) ���#�!=�)0�fe�D�z�+Nb-���ܾ%�ޔ(�\���h��^���t���S@���:����%�dgZ��f�O�MQ�O!~�Cs`���6�盍���(B���n<�	�~�Ɔ���X��$�1|d7����QE��Z�{E��g��� F����B	�{<{�R� �=�}U��!��o�I<��uXlxVHYEB     400      c0}'���}�rS%�!{Qv%i��Dv0��R�+m����Zۑh����G�3L�-�ͽR-gC�H�>B?��w�~TqA���8��zC{�Dl�v�U�n�m=��g��KD�ۉ�Q��V���Ab�E��p|�mi ��׀I-��(y�h�Թ՜������]��
�o��/ЈAgcEʓ��V�������aXlxVHYEB     400      e0<��|�ھ��g �waȦ����B��Y�_��ҋmN������;��_�_2����Ҕ��]؟����ڮC�,���G��Ψn�#��{��g�[�s9��f�`й��<pj�{+�<r[b~�p����o@���IpH�.I8X�?��~=j3��]X�*w�E�P}�N��n�հ���w1x�8��^@�g��-"y��ujkG����@e'�=� 1��YXlxVHYEB     400     150g�|H	�̄�1AZj_ `�j�����Y����C�PP�p�eɔ�x!V�?S�B��MB�&F.�@��[�`�9�J#@@�Y��6�Ӹ5��&�$<�<�����u>��. ��@V�5f��u�b�n����[s���.$�* �YQ{��:���*�����@j��u���X1�Fu�-gO���8R4�8���Ʃ�FZ\K���Ӑ�Ҫ��o����R�n�Y1:�L�P��f96�Ñg��ǿ�w���hb V�����W����ZP~1���\:����h�K-�)r�)�9ںi��5�w�<��n�r�cfl��d��6'����~�j}I\2XlxVHYEB     400     160L� �U����9�o⫧pbQ�N4F�}�s��t�c��ldᗅg�2�/Zh#ZZf��H=�o��<)�9]r���#SՂ����wMW��O���=v�����s�2�6Ӡ��i��*��4'��K��f2����Vg��iw��c��ȌT�C(����1�Ӑ��6��(�q1�W���@�H���c��Ԫ��v�LH�rq��-�#�'R#z$3��b�+�����r��J�o55�\�Ƹ`�d+4�a�E�C0S�?â;]������R�֮�G�����C��R]d3P%x?/cA�9H=��I��%����R��A�5��:�``��Bl�ʰ��c�h-�ZK���XlxVHYEB     400      f0�0��Ĳq�j�J��i;G�*�X`~� ��|�h!�<;~-2��hY�U������E�ˣs+w;���_����ڝ�.�{|����-�3��� ^ �
��]&@�~�LtĎ_o��\H��ox3�'��C������J����ز�ArE,m�����@*R�5uJA���vK�m�� ݍ�,p���J���6�����i�����U������*Jgf�����I�\+� �ӌ��7O$XlxVHYEB     400     100'�����
|�짡�g����3��ƺ5��RBz��&>K%I�
7�o����Uw���mϟ�6j���=��/U~X[�n�IV�of�jpl&��3?��ә_cMc��:BT\���c7˚_��6� ����k�M��_�:?�k+�������2�VsVw��2n���3��Syvʃ�����u��π�:eg�g\A�D���K�7hb��8W�kr�ie��ۨ��@�����WDg��c<C��Ό�;�V���XlxVHYEB     400     110 ����B�z�EBՉ�I��?��elC>��]��c)�����/����E��6��&���l�b�y�ͱӎ������G�k��'��EV�b�]��f�;�C�X���*Ӧ'�99��+2=�#����*���;7�ӛ���G�j,[|&�qs?'�Ǫ�v��8Qb�~�ƍ���c�7���o;��Q�a�Jb<�d���}L�V�p��̳N���(�)�<����r��o�mk�h�`���Ʋu�[R4�C�\�:��Vm��Ge�?�XlxVHYEB     400     110x��t�?��)p�o���j�uY�S'��>���\G0\):Fs�7J��C��bf����Y�+G㡲��(�-I2�����{Bz���n���o��q�3�WJ ��2�?i��"�jV_w�3�L\`�y��]z\H�o��$�ɻ��L.<�*ڻ aR��@���Q�w�����/�ʾ�����e�K||Ƴ�;Up���'>s�7��g�� �M��a5v�l�#$��?��Wg�C6�Cd�����C�Ҳ�5��M����"#��#��U'q�mXlxVHYEB     400     130�4�-!U�*��USq�١�W��w����K�"��[��\��&Ck���[G�瓿��#�v��)�ǩ��_�q��%b�%2��5��#g�m,�����*̹�Hz8;[��N�)U������ ��&�6� r�|}36�[ktn� .�.i����v׍l�V�B��A��j���Ty��,3�)�	9�1�&W5�u�e� _&qׁ����a(�~���nT\��E��ERJ�J�}�181]��a�z���ƄI<��{�Zў���bKJ��#˘�/]{��H���W�NM�Li����=zIi�tXlxVHYEB     400     100,=E0Ӫz��6��⫋�캋n(�o��4����;���E�E�����6(bʦsb�-B��7߰Q���?,{O7�^��2-g�^�J@��uY(���wMF����E��G��Ƥ��):�3:	�n}�0����N�}�
d��]]צ�B^F��6�̑�!Q�-��׀J���8���3�RO)�{^��)�������-��tL�ԝђ�g�T�5�U����sF��bxV��S̅�]'z5�ƀ�aXlxVHYEB     400     100����(�)"qe)�CX�M�y�bP�Y� Ւ���4��W�4��*R}�Ѳ��>�+6�&���J��w77��k�^��J�:���?"��<�;8d�FAV{x���5�-_F�d��><�+���n}�!� ��B&/� �Ԡb�X4���Z�_z	�W��)p �vLF;i����/+0�8�m�K�����L���ҝ�/������
 �wP�~wX�ː9�:,p��;Rs3���zn�n)���PD�fXlxVHYEB     400     100�'<��1	F�K��vl�FO�K�� ��vҚP{a�7~'��?W�OB��T�����v^W�쟈�]ֿaS>v����;�nd�|�X&/��
��M@��G�N'��YL�΄�܄)(�J������&��R��adv:�F��S��\�d���C���K�:O�ֱC��ޤ�C$��/�2�H���y��'0�HC��
��Rh��|��%K���89"L�~�.Ԇ���CTI2��@b鲀�\�Q=Q���	� XlxVHYEB     400     100���V���̹dU��Wozo�!�|׺/��̬�S���@�y����6���g��7]�kK�|*�Y6��T�#D7^X�9�]j:�G�
�E� �6��[z�L��m&���-�Ҙ$¹#���M���:v}������7!���v��E.{�8G����&ww�~�>�e���^����b�6���������$�ͺ���;�`u��z#�'�Fv��n_�k��'������jR��"\��eXlxVHYEB     400     100�<����2�Z�.81����IPX�lɼ��٤�)���ͩ�ǈ����>�xy"��"�*�`c�K1�S�a�k�=���
�һ���H�J�H�^���,W��v"��0|[sIꟍ�F>�İ���"x���|��_�6�����=]^[ϱ�N�8v�s��Q�p��F5\��A�%�/{<����ѽ)���J�2�v�����i��ZX�^|��MHH�ӹ4*q�`�t��㐍rC~6z���+�L}$XlxVHYEB     400     100�<����2�Z�.81����?-"�}����Η�ʄ�@�X���By�F93^�#R�<pH�{�Bíac!Y�	/������;iؠ��G�bz`B��*�E6�>/��,���I���4(<�*�rY�WԊL�{
JI_�q�w������ӭ�`�8�{�Fq.PN��!��?j�d��(��8/����#�ʪ���"�ZD{����"��ƥQ-[B���&�ꧯ�L]�.(v�j�jo�h
Pt�e`
XlxVHYEB     400     100�0��s��)�T�|� Y�Ǝ�K3VcOZ��q"�y��r+�=/ ,�Uɱ��$4�U~�n��4@�`_��_�m�����W%��U�"��}�72iAwj=c9H�FrG-��p5b]�"l�]hlx��_Bd�2r"f�Q�섅��.��M��q�[�O4w1�ŗm]��}#l �'U���Ob���t��
b�����E��0U��D��|ҏu���#�/�:ʝ�xJ>�Ȧ��c�7�'�	�h���u�A��ӼXlxVHYEB     400     100+� �kd���IbCb�5��A�ռ:9�����;d�Z�2����N� AE>N��=��'#��,tDL#4wMO�KP&`.k����B3�]�Ě�t=��d�hk�ɰu{.��;��n�,�� (<m���o�g���"[���������Ӛ�<��LIZ$ǒ��*Շ�k�"�<�&e&V\-��$L�����������;DUk,�ㆺ%�&��.xve �w��̓b���[g�xP�p���X��XlxVHYEB     400     100���IG�����}^g��1��tBl�;z�1�v Ǫ"��u+�>��$=��E��9ID2~~��{�+��� p�4a}�K�9�	{o݊�����~#�%���<4~F^nU���9KGs�GM�=u ���i���b��a](��:���5�Uy���>�բ�^��\C��݀�m+kc֒:�-� 0�1���s$�[�p6��Q�;6w�%I�۲̳�A�u�#p�7�]��l~�w��V��ۘ��H��+���.��ۄXlxVHYEB     400     100��b���GR6�ݳC������R�ZI��Ē7�h>ɇ5O��"�Z7'���w;F�A�860|����x?1�P���i��^d�[���3B�\ˑJ��i!��Gf�N��2��Lp���`�_D!`��[r�Lc^5��!�O�s�G׺y�]'��i@���ƍ��G.B��IiX����7��SB�YwS$4\�u�GЎ���POs~|&�7����N �2��y���Zh	���^S!�j&ɣ��[��XlxVHYEB     400     100���Λ"���e��?�I��9�� ߆vVD7�l�e^I����-��^�2�q�t.�Xw�]�H�ϋ�D;��:�/�C�j�ر��lV���OY�ɄvV�?����׀":��m�3{��ͷuXm���U`B����2������F�oT��+k�������u���)��ɰ�C����,�A�#����R���Ud�˭�gWx%�H��7�R����UO�hTN��8Ӻ���,ɻ��M��@1�<��CnC�]�`�l�=�D�XlxVHYEB     400     100u��=�uc?�h����z`��{G�W]�nK>���Y������&����8����y��}�}�!����7w�Y�1�Τ�B����$\�����<���n���䐋��a���v*�涆c):��0�©d9�8��;�ߊ�IS����ˡ=9�$�	�A:�B�Ă�+̵��H�\7�ɤgp4�y꽏qo�#3 ���:��T�Ͽ�W:�����${�Y��THc� H�1�Gr\-_ү�2�Hu�K���XlxVHYEB     400     100�
q����Ė���w�P�_Q���k���zM_�+����U�g�6�7뻗 B5��)��o13�p�0Y����7����32D�;����@6��_�g��=�!22���̒n?�!o�u�W�X0�>PZ�:b�:f&�^�_�ij�az��R�K'�gV�hj%иE�k�g�⃰�D���{�&�hZ���kyi�0�j�����ᓼ�T����p<֤Z��H��pR�,�-|<R}��"��/�/:�̆y
؉����?XlxVHYEB     400     100�m@$������1��U��a�t��	0�u�W�iI���G�T��(Hp����RUtq-��s�̤O��H0Ǿ�9z�����q���'ge��эm�&���� fC�A-Ǌ�o�l�f�$l���=�2l�Ixr��ĕ�����z���ڷ�
��P0��dq�qݨf�|1�"lB��d��9�
�%�P/3Շu�S���z��5g�aR�\���̿������g�b��-N�N��q:G�.歸��7XlxVHYEB     400     100�#l�񋡺mv!Z^��R�Rz>���@�f:(5����9�(���F�|qMwr@u�n�B'���(��-�e2TB�!�C��:4�80R�f�1ﰅ�~8N�b���z�u�?PWt����l�)�@�V�φ����t�!�Z�Yち���=���{Xy(b;�}ûOn@܌��VZmՍ���R��[�s���S�WYС�����=���պ��6'H��0��2�'p��V���Ce�H��
n u��2kXlxVHYEB     400     160(��JM�(?��q}�0�0�����o8�R���S��mW<wZ�\���t���A0��/��o�Qj��H��ԕm���ʖ֫��]w��E���E]݄*e裼�1Wi���xૣ7#�1��}�\o���E�v�AG�@�\m*�ǃ	�H9�5H� .(�yݳ~gz��Co֭}�~��r��on<b}Q9���#p�SbG2�n��-�pl�m�����u7F�1�3t��g$z�!-�{U&�t k�'�Go�u<$�p�,���]?�H��☨4Q�>xW_|��j�  �s��o��O��ǃ��c�.��>=���|ڃ��X�Q�7�xr)�9�L(�XlxVHYEB     400     110�
z��DƂ	0��a��7ZfM<#�"�NC������񯚀�Az��c�8��u��ݭfLk%���]nk~gb$�
�`6��f̴ͯ{��:	na��Aփk��K:X�
�~WU[�i��k|EO�'���@�ܘx[f-���1�����<��-��a��'EIu�1��a��}&�Un����y�.]�����6�9�g	��hc�zơ.nɇ)�M)��O\�E�soU�s�$��v�����um���\l~�NMŞ��_i\7�m�|R�ϓ�s�EXlxVHYEB     400      c0��ư��v�2���ʎazz�M	�_	���7@�9���잛Q���$�t�m���0ϯV�����	H)��&
ե�8暸��H[��e�0�W�&�, M@Ǯ#.��:αuI���̒�ór�5@O�OYr;�շ޳����yY=]�����ž}�i����1]�E? �%�
���\�����oXlxVHYEB     400      d0T���'�~09�Y�vTl��iu@^B�uы�zT�fK��`�`(����!��0;�N�6��]Ϟ�%�]y 1��{����Ri�6���<���g}�f�.�¢��}&{�D��(#����H��W�Â�b���Q��.�K��Sn҇0ɵw�p��wӷ=�o*(���Ӧ蔟C�*:���҄
�7�\�<_��XlxVHYEB     400      90�)�U�����̰�M��&��v�Hw����<�X�ɟ8B?�;��Zr�
*|U5���`i`�!#�� GH���(�F�����'�(�s;����U[w'�@R��x3�a#���y��n�=�,��N��`�$�~]��!m�M�>JXlxVHYEB     400      905��N(��g�5S#_�`���He��&�ԑ��ƇpmP�Ĉrl�#�T�𴃈20{�tyR���j�.Kf��L5����7�k
��h�x�̶�YnA���C�d����	��P�I��$�1iR�N���K���1���-�P|[�jXlxVHYEB     400      90M(y�KgXg#
�-R�y@��ܕ�A�����d�i�}�߳���<�i}���^�����Y���e�k�f��1.ܷס�X��! r:��/�na%��c/���`���n�f����Z[{T���C�'1|E���}.���OO�c���'XlxVHYEB     400      90L� ���	�{���~�1��z۶-��NN�}B�_q�0����e+������d�r�f�d���m��%w���B��2���z�z6��]���qs�>��p8�o`���ڨ.���|��Y?���u	J�	����Z���uXlxVHYEB     400      90�z�E?W�3�W٩sK�� ��u%��M,-��ڤC�]�.��S��ƜE�LA>E %X�{�9���M#�Y�IG5�z0��mT|6�b�h�M�<3g�Tk��YT近-�{�ݡM��Id����Q��)�ԉ���X�$�eXlxVHYEB     400      d05�Q���Ή��o�7�P�����C�Z��[�T=�Pk�4������-2���A��E��[�����+��O0A��P�O��?�	�g��%�QC�ҹ��Qw"X.�ߖN��D=�H>8��u#��4`�#[z��׆�����lT��5Hhe9�NnxM#���A�Q��������e��rC=#V���&q���������6����XlxVHYEB     400      d0��v&�x{�U6�b|-�t?�8[Z�RIK]�C���r����E��f��8E�>�L#5�<��*d�6�r|FT.C�X�YQ�k��uZ^�#�ϋ����<l.���G�������k�`��F��=���8V����q:Y�<�= ����cg�ݳ�X)�n�?5tLq | �R9)h�4E�sj�����ɝ�.����SXlxVHYEB     400     110��\�}-Xs��T�ዊ]�/=���WA3��Cz_���}^Z3��F��X/{��n�ׂy�9,NN���#7;�X��l���	�;�>�ʕ:�gw�������u*"H�63�YlU��S�/nu._	����p������'�$6DX��H������N�e�g9h�Nq���q/^߳�>�	�E܁� �m�D��Q���kQ�Qx P|m����� ���
����ҕXGf���?	����\�1�71�	�`;�G�����UYXlxVHYEB     400     130��,QɅ�S��:�������r?0������,�;]��L���m<v��Dq^�:ޘ��'���-F��t?`@y ��`���`p�\ ���QqA#�ϰJ��=��!dwA�u���T�.B�M�(��Oƨ����BU�4=X�������y%����_irp!��$\�R��F���1����2�NI�̏�R��g���qv�B��V�H���-��q�ԯ��EU��yu��y��H���6�4�3?B���QO8�i����81���,��)�/�d��E�X��9zY�KXlxVHYEB     400     180��ѧ��!k�w<F�{W�k{{�n ��v�7��@��Q|7%�XW%�W.eJ6yM�z[J�㼈X�4����ҥq0�8I��{� ��&i�^*_��NVx=d:�8�B�� ���#������T$�;l�0E;�̯Ix�κ�	��"�!0g4�"e��7����jx.��sN�0h|~ѽ�<J0�����*M@������`X�Ah�l|�YXf��JE7�u�]�JG����~�A����Q�"�&ݶ�ԓ�]Qg���\��_�]���Z��}�H�Ϯ"%�3�����I��_iFFw��f��0s�o��S �aL���ɏ�1D�����=`%ڹ� �D�<���_3�ˋ�9ލ��ʥ&�%�R֬XlxVHYEB     400     160f�8�4�Y�ryp�>�����Y�0#��������?���� ���MÔ���gD��וU�koj�d��~zgI�2� �]x�>�a���[��|�攅ۋ���Ϙ�q�0ܟ��>�E|�b�O� уMZ ���,����Q��������S�C�Zt@ �f!���� '5S��H �\�.���!�®~�T�[���3;"{�W�����+an%�J&.ܘm�wq�mHĴI7��~�vS�T<��^�wr��ܢ
�	I��=���n{���/k��r'Y}ς�M�Y@W����������u����~D\�����@�t�55�$�2�Qb��+R�&#�G��IXlxVHYEB     400     160O)�Elr�)-�l]sDKW:��avxR��/yޓ�a��v*d�t�	J���R�f��)~��$��D��W'`( �,m��׃��&1�؂¶�D�$�lw�����k�HD��bq)_8��9���_M�{jCٰ|m8�
^��BS6&�E��l0� ��\��������8��#-���~vN�8��J�#�T�8�%u�Q����9j��
/����SZN�8��*1����@�Z�h�;�nT�PW�`���[N��~Y��_{���3?J�Л \Δ*����WQ�����!v�5kyG�{W�b� 
M��=ܱ�����Ya��ѭesS<�(c�I�M������Vp��1%�XlxVHYEB     400     1506��D/.�8gT���W�Hj�7��2���[n��90�ӯA$��Yo���|�&������`�.��`���\�=vуx �"!���Yw)�#�e�/1؀�+J��J=Ւ����u�����5�0\w�H��.l�)2B��������n��y{�@�vԏteT�,�7t�M�vH�^���2�۸��Q��sT*�U ��ޚ<P�&���h���%aE��Z��-~h]����LF<�ޱ�;㺉�Ě����H��`7�0v������GĄ=��ڧ^�n�rrH�&O�x`#��;9#�O�h�S_�^�G�D���QIy��c�BN)i0�Ґs�6�uXlxVHYEB     400     180�W�a�:7(�c	Fa���%6r��"/˞��u�����X�-��C�Ǩyz����H�慞�/�wOv�M�����^�i:Ot��~��T���1E1%�j���S�]c��!���<��&KO2~0���J�|�ii�,�;&�.����E���,Ll�w,ۖrh�_��[��p��q�]�B����M6DG^���Z���B�����2g�w�O|o���Q؄4Gr�F�Sx��S���Մ�&he���������Й�ϲ[��ґ����Ly���_�u��"z��8a�D|2�E�*G�[��I���t�N�.�1,���R�g��i������s�>� �|�hB���%y��S�Ϭ	��<�yG{��1T��XlxVHYEB     400     120�ť��=_$��v=�ވ��ϒAxg��T�+�2��A��sH�y���<��ɅN#p�I����i�1�ɂ8?�_q�
X��3۲t)�F
��e���d�T�;=�O�VG邏rN�cuR�JBrt6c1�C.��g���xm�k�uf��7�uƓ���RS����C�s�pI��k�!Jԕ�<J��t�;#���x�a~C�E5^�e�Eܶ%:����@�	�x&����վ�p�hqB#!Aȸ[� .-"AE�4X���7R����8��'᣶�� �3��\)�CXlxVHYEB     400     130�qb�))�{7�#��S������~gc(�iƱE�ǵ������Y��YUh?h�A���*x줶�q�_|�p\�as��0.�0,�̌K����FFu˳w�Q�q�[�!m�>��iѧ����8�v�Zpq��j#'�2q+�Dy��CA!�3]��ҽ�媖���&o��:�8q�Ip]����9�^dn%�t-���P��}G��'�36K���$�4�ABu�\Ԕ�C����?�`S�q�>'�b�ҽ�*��za��4\|�H5����Ѫ�JSM�2�-���� ïsCX����5Vd�f�i��� ���dXlxVHYEB     400     190D'�w"-�1Y@
#���}y��8��V��0�H=U�-6�ҙE����#�N���W���@�KiS�e�Sl�f�Ac2x����xZ���ޅ��P�H;� 6χuH�w�°�sUk�)C�@���j`�$�^����>�����MzC�i�"Pz�I�p�B"�"}l �����1Io����2;���� \z�=�=���H���w$�c]�O����(	|[�m��]�\N��Sb�8�]"QS�Ur�y��q�FMT�Ǯ7˿�@���{���c�����r��"V�9�vZo����Q��s�1Ckjqi	��u����ŭ�>.1RZ0���Ļ-b�s��'��4�M�����ْ{�l.۔�2U���(X�F�]ݾ���O�������#��#q)(��XlxVHYEB     400     1502��0�n+=kn�3����%�Ѥ��v�9��Pȱ��d���Q[�"t}]�4ң�_X*�bK��{M�<̈́���n�#�j�����@��]�laׂ}����J�$9ġ�x�Ľ_�+�τ$Yn���tr0�v&�f9@�?,b˗�p��]���JY�8��|��yq����xo"�D�6�⿺�Z�,��n�b�/��(�=)���l�L �)�4'���L�@T��e�u���:����+4n}|�f/��@�����2jx~��#[hl�y:r����!X��]���d��Y�;�V����`��j���J��s�HQ1����2Q�^�}�?�XlxVHYEB     400     130���=�Żo�
a�����H='�2������J*�J ���L>;����r%ʚ��)A:s���{���)���J�=�l�뤐�;���%��:|S���T��	~���'�if@��"dP�{����Z��B\�4$�O?����``�˞���ɨhd] 0�a�+[��H�'�Gs7.�Կ��U�ï�Fny�WM�������f�D�zOj������@Y�N��Z��	��KT��eT��Y���K}��DK����S`Ѣ���s"򙨭��L��l���=i3Քe�7YpXlxVHYEB     400     150ʥj?�â7��W�;7?��oD?�� <� E@��a$CP�?״sKHf�&i�D��@à* �&� ��lgQ~�XvQ�Z������a N��������O���D ���%��@�[C� m�3��
�Ѣq �I��Tr�Crqg�_R�W�LdK�/k�-��Z��S�5e���n��Z(�}[�tnےE�V�-�s��+z����y�6�Uz��e[!t%�� %���qѻ(��rR�kg���z�I����D�j3��6�����{����\8aJ��I݊).��e�� o�7<�<x�;������м͏��B�Ǯ�5��XlxVHYEB     400     160��:b��I�Xk���[��jv~ݽ/ҴNkr�'�s��gF�]X��R��� �!�*<0�՗���/����*��vW����e�5�B��*�U6uƛ�������S�%#�T},C�M����."Jˬ�/�%��mО�L� �F }�V-�f��2j���:S2�0ҿvQ�����uw薑�yTu�������-г4�C1���L�C�o��`��ĚZ̑�7��#l$ו���h�AK�*�eО�]�x��>;@:�6�Z
t?�]��/E��n9��N�o���_��
�v����ɼ����Y�8]Uy�#ĎR�,����}�ǈY<;�c�aB{�^Q��zae�XlxVHYEB     400     180��F9��L���2�l� ��d���R8�V,��Ҹ�)�
���)z0Ң�&�)%���s��(���yՌ������Ѕ�U�W���jb3�q�{��iw0k�Z�p�ķq�&����2cIK�l��%���{�6�1�(�>�-�НH���U�M����&�o�(�X�(��s���Fn�(R+l�*�!1�G�t�cK����;�Jn-�Tݥz*0I���z{��)��@	����2$�C�9|�������õ��M��R��#�z�; #5�>�����l�-�������-[de&��WA+��ߞZ���s8��	��')����V�틫�X�i�rBSQ���Ȭ���7
�Ԍ��Fp�N����XlxVHYEB     400     130 ݑ?�Z7�3F���Rm��k�G)�_Q�Tf��7AA@ho�G����.E���o�~H��Jyu2�#ᙟ*�2�gj�W���C K��3FT��zܿX�B� s��ڮ��QV\:�:o���A�C�.�ה.jM��O��c2��~��%1�Lw ��j�<�=���w	r�J^M؁�v���=1g�79
5�O����eز0��Z�����3���j�Y��Ɲ2�.>�0e �t?Z��$C��5�O�B1xw��&-�ET��a��ty��O�fY�j��p�D��GmӪ�(;G ��w�g�B�q}XlxVHYEB     400     160�Liy��w û$UB�UϷ������߹� �Yv����&M1�i�<*�GH�[@���<~����6O#���l�c1 v/���˩�0&z�hB��$�`H�[�8
�%�I��}.sR�X���H�|����y��f���<.*�6�[�=O�g?4�P5��הB&6MA�((7�TE��%�Tt�����������R��5 �(b�	Yw��; Âi<��	r4.��jW�Ca;�A6ₛ^�6�m�L%2���U����BK���j�Ύ\���<�P����<]b�ߝ6OP��ܖim\w�"V���4����|�L��g�K�������#�H�#�*�5:�jRk~�XlxVHYEB     400      d0Ҭ?61�������T���g+��;̏�'�+�*ǜ��KN�$��z%���Q6���+{��Kś�u?�E� �\ �ߢD�LJ�m���W7shhle�Imov�'ԉ<Y�5��A���:C��7`{�o4�o"L��A�H�z�h����]�E���Nj?���B�@�[$��Z��Ȓ�V�Y�o��eW�更a#�"�V˧X�6XlxVHYEB     400      c0qh'u�09?jp �󈝫J4�R瘣ͮ���q}w7n��KYz�"�p�:��?)�n�W�*ɬu����@���ŮзN��fv k�鍻q!d��n)F�����m���^���5eW�D��s8W�����^v�7�d�(�9�-Ÿk�t��I�+,X\c6�"��B�v�����s#�_��@���Up�XlxVHYEB     400      c0��p!��,����l����縺� p� ���VSa�05��:��-
��E��?]5|�sV��{�s�Ì�h���_�!�eףk��{��~ W�Hi��je�z֛�v8�:e���?0��`�q����FU_d��|��[؈���5K+,��wo��,%N�-���H���J��k�(��|�K��ŏ�6~� =XlxVHYEB     400      e0?I���K�us����-�P7ڋ0%p<��6d�TI2��U�D�}2���5놬h��'��CW�"RC�˲�4�-nǣ8v�>�f�6�b�w�#"c�F{�(t���3KR�Jۿ�ڣ'v<X)��G9�K�ϱc^V�Av�����<�������wI&Z�� ���]���"��_�4��O5�-��>��떭u�f�i�v�Ĵ���v}@9���Õ�ژxXlxVHYEB     400      e0����ם=l]��7�3 +�CX�uI�K��+�t[��è8���9I~�UD�p9o
]Q�^?zjU�%���N3.^3N
=x~o~�5�v�V�� 7Rg�!o����ߐ�ē�g\�Ѝ���Zɧ�h�*/���̶!Cr�mW����֢}9�����&t�	��H��heTG�ũ���?3}f��.=1�ˬ UK%����6y��K�f�U[������_�XlxVHYEB     400      f0�����5�Ϝ���c#�d�˖���l:J"*=eNHzw��E��x#m_�Ϡ�AY��(c��u��!f.cwں�BZ�m��j��W�����'�T���%�~y�s�d�ܤ_d��2�r_8�#f�j��V�J�A�)4��Kk����'��a۲a�n��,���15�n������/Ʃ^n� +���M�Q��y�-\��x���R"�b����GT�l����p]Yv�0�` q�� �	��R�XlxVHYEB     400      f0Æ��F����;��؀@w���:d
Ǖ�<"��R��˵Q�*eW��?Dp4��&��$D|�@��f&)�����G�ed�J{�݇�������+1�/(]C�Up{)�;�t싦��
��MWĕ����Mo3�z��.���W?W4L���Ǽ���jG���E�����Xm!���E�nF#�gd����.�ĞF�"���P��F>' ��$s�WB�t�sQ;���`��t���XlxVHYEB     400      f0nA�X�0��M���<l������ԡ���#G�T�����R�A^[�� �ϣ�{ =Z�s�\�!JRL�r>Un4:�"��1��������D��XJ�-d��MGů�Hpnl&w�\�{��R��TV2%%mNā]�Ĕ�c'���-�f�i�����-f���y�[��_u"��V(��jf����E�5���
M;ܬ|氂��J�&-�R�TH�X�W~qT��ɗ&�+RyVpXlxVHYEB     400      f0����������	�;�x���+�1j��iyi�N���������iY�gP�.�i�?��M���N��_蟌5��H�u����v���-�_��qL� �U���;�(�S:#O�B���K�l��F|���@�㫶�Z�'\��
����@?d�m�i���+"$	z��\R�+�Œ��T���'R�k��a�R_W-�\�Y?Z>;�J�j�֞�?�a��T�TSk=��XlxVHYEB     400      f06��^���cU�Y�ȗ���~��I�q�����k�A1�^-��D4�w�bcTce����I�S�u��NT�喔�'��bzUZ�Hbs�j�O�D�1��Vd����
SJ�+��q��
�A�+�*�G�H��}�;�� ��x�]��q��P���oH>�o�{Q9)-��޻莞�ϜEa��	-@��T��qD;����4Γ<0�zy��������M�bd���Nv���LH�t���XlxVHYEB     400      e0K��2���e��e�*���ǀ�jgU�,
85�	����:�e�_E�߄����;�"G̿��4D�\-�W"PB�}�������X����D���w�:�P��q���p�G6��]�I�����щ�@Z����[�d����-�\W�(�g�B����Ï�YN9Us��jh-V�ѩ�ä<w��Z�8�_w4q�CM=}�z��6��"B��%m�_iw8Yɦ�ٽ'��fXlxVHYEB     400      f0�B�3 rK���Ѷ�2	?8�>��d4��9&�-��1�w�v�wOHu��h�T�i�k�_��TxD��
��2i7)��X]��.�7X�D��R����얈���)9F��%|��������Ȯ��!�$�%ѽ�ur����`��Ζ�2��}o��:O�I�� ��`�6�j�����F�&��.��K峨�h����7o��N��ृN�20#ѾG��s��˒[2�r�XlxVHYEB     400     160�߉��Z��9��^Td�T0+_{���/��{��MB�PNVP�|B�e~�S���J���MiZj9�	e�]J�A��ek}�︋� 5hj4@<i-��⹑�[|�� ��6�i���!��UiR�qZ�|-��w$�y6�#>:&|Z�
�L|�b�r�2� Yx�f?�ȵU�m��X�UAy����,�3��w$��� � �����)�d�/-��a�Gt9ȱG-�S�!���.=�$g��̅u���Q���?�*�y9<.�P^;���D�p%�?K$�~��7B���'�#$�= �?�Z_V��������c-69���nW�Oö���_�uH�XlxVHYEB     400     1b0G4�'��#�~�XHw�uh�ƞ��oG[�{i��q]tB@Uj'!e���q�V�����b5 �yQ�j�5���]fn��1�OE�>�����D��=qc�����e�>�*��j2�ܰT]b�����u^�G�@L��2��'��A������ќ���?��2��s�E���^- P�Ym��/���Yʕp
��:��vL�|��f��yj�/@������$�*�`�	 s�ŻF�y�L.���\R��E؆I'_+��SP�r7�]ꊢ���'hM�����z��|հ�A�x�XZ�����c�j)ϧ�SU�u���7�%Yq���CD��x�e%%v�h�Vk�RW�P	dXdB��ѓh�	(C���eg,�s��H�Cۥ��җ'��;7Ǹ�}ㅘf2�P-�摱��}�XlxVHYEB     400     160�Q�$eM�^⤝�R|�0�s��5��?��P�񄣦�,g�9�v}�e�]J���ZXu��: �C]vL��a���''�%�-rkXH��R�zQ��/F��-䥒�P�g0�Hʼ]K1cB��x�2[H�7�4�r%�k�^���֩_��¾���{k��h	3qf�d�����l������:,
�� ����Uԍ�U=��*N�o�C����FQ���wa38۾b�cN�p��B����7EyH�D�U��ޏ�������¨����!!��μ�r`i��_��~0���zc�xNS�dmq#m\-k��kM\�G��2��60u���L��ue4ϕ�6�nP�s7�R�XlxVHYEB     1f4      d02X�rd�,g.��aF�!1v��t��P1�5��V�G?�\�G@��JӤ��p4"�E�]m	QWi��)8��@#	��(�f�§ȏ�Ӛ��QZ
p�]�[���Ѵ)���%�����%+'u�}��~ �G��%U�b�
_�A1X��)���&}>�0z��Fن��ؽ9�B��dAmf{����j�7?m�J-��ޯ)o��_-j�i'���