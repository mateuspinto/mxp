`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
OKUnzzO58i7JeT7VRUchTav1iSCY8nc+RoZ//G2O3vCu5Dtv8h5Eo7sIg5OBEhYj/p57hs0zhYES
rnSMkd+3sv+SZfhKkxlKWf2h+0U1wcmuP6zRnslz2ks1c82+ikb1pWadIouwNGWdnhswyjdKyM00
gGAH5Z23pMYtkgxOu+0NpeA/3pRnIHHXc0u5Gfei8WnRRDuFUzvyBanyPIUEpOj8jcQl7DwMdX5t
dekLYl+q5EcHpKP6CU5TQ1RtGYMNgu6sfJfYmupk+KAx6td7IQ2U8RkTaXL6ca7/BEKgrwtuMwmX
LlN4bKCI1tdFPpSk5fY4gQdGnAbQ8tjqpWNxeA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="n0HsDLAcw7k4Xu5KpugibqYHXqWaTmJJvNaLKsFFqN8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 94592)
`protect data_block
GpKgESN0sfZsC17TXUiTOraUueuQ6IOnWg4MyCbjmf2UQniuLiufkuivAw0hp3Qo0kVxjT0pT9HV
YVvJylfnRQrvTMkvUd+NkloZYs69nLTYIJf9lGMQ0fhb3R0cx68vViOfyZUNhnw+I5jYPxdR2/rQ
oR7tcSNVQbVzNV/rhn4pxumTj7HQgLapSwbQLyR5jjeG7haHYJ3ocEIsM6U7oRrb7jcs68jxgnsZ
bFEke/gye39hrERNF1HTaBgVZVzO4wI65pkw3zoZ9PhYDtAgBvia7cyHSD3kmwqTk1dLQXjYoOr4
cXCPowiQJlON/H4PoTHU6AG7hcZozjMmQ40RdIKnvHJxQWL0z/EaVUenUVcXSWsSO7bT80GheKjr
z4Vr0DkvQ7seFHLkSuKDuIgSPAQzmeYGncAloyTv0uf1x+YhVw57aYJGDFeU3vuzgbpFw7uYcVfM
2rp94aHXvGXrF/6w9wBzt5YQSN097XPcwcgolDGXRBH0Sjh8xXsZwVZyTB+aJqYDHNdoNlEkIZXL
eUuDLSQ5CZ2eEVtOs9KxQPYqM6KyM8ug5OiKSIYMSSWndU3bKJvXkT/WNUfpwJUwKLErhEk5Ieyl
GmyYr5X1keYLlgg6P+RLvivSWzUOHSGhr8wzHEHs97kt06J33kkHN/6uA5sJxvvohvHoPO3TM9Xm
3UGpO9kxCK56dTV4fwWyFmUt5nzjFLm4YWdLLi5Rsoe9kTUuRfli9SrYKQABrFpakFDBlVomILKv
BAvj1kAe/Uwn4an8yYMgo2zmjV3WinFb1nfZhUO+5VNfvpgVtDcU7Wc62R17c/aJyz85a1Kz2kG5
BcezxZm13JxKuAX0JR0Rd7ZtubGTIFre38T0svcrLmWEqNkHoFRIfyAe6dd0Wecb9gYtnp7CsnxO
x/qY3qGzn8TfdYN3FnQH86uz8KXPSSytERYsdw/CYg2u+USsTyjaoIsRQxDiRcTa+eM1k3hz23iD
Xa8ozLmeiW9h5238EdXTME84BIg++pqBiTYd8hHFoaP8kXCSN0zKZCYeWVaysEY4j31qjFbVlDOh
7e+DjbDJGkX4vxaSOA3LIxHL7HFiOD9rjA3qi9ELemC4PX/IOTe2WGOkpigy0Tb7Oo6LTtWvUBHm
bFAtZdk4Yzsoj/apmdbwmyL0XOvgvv59gfLeP28JnQyarx23B2kiczUAPX6VleBZGiNxUv3s9LjV
hPX94rEFBNXY7XmpS/3Zz9VCR0xD56BWy4+9nI8ABe9rMnWziLUa2YWlzhw6Syk+OR5I8kOl+aYO
xT0j8wKmsg2NQWsHeuxbJhZgZPGypbqGcRC+13I/Vhx9YBGHZozm8LIWRitcBp4dNzk986Wwz2IK
fQfybVuz9n8ZJsIYbqPN77hnD/uZ7h4L/Ijm69QFdwLTYREXuV2ayzh4tm3uTPmG3MeHfUi1MvBA
N7CZeUf3vugsgDUbY8rveUEATaf4DIPFI6djEHnGC60kjtseNegLKx5bdZ2qcUDvgEpzp7/BS+/8
SRpCAkfrUSff7tj8b9oAQJNHrbv6qPHJHyCBzWwuul8KiutcMGzoJOQl2XYmbvoK1RSTO2l9UUD+
TaaMnmRC5arnrhsPTRFIqM9dsmOZu45IQUsZXWLbrK9BCL7dmj+uGEGhZX5GyhttnKFUisrGy99c
rb3qVfaeTq8zallYEGI5AcMuSeJHEb8bZ/1UOL35Cn6ncVolAVumWQq9GAwkWoEi3GVF4S7iW8De
LjsnByxNKEjaBReR43tThDLUyVVpCdLpirS2tDpMyzxZm1FyqxkzzW5NVor7225VH3sfFB1X0mfJ
8YVvIJfbjlImxKI3wuV6EsmqeQiBY6zgAbn68go8pgFdItsp9XGhIkvf04jn5lrPMhkNaUoWMMml
gLV3eNWH3MKv1NPqRq5MR+eysZfly8wZ62iq2ltPY5/SPcwOKd3ybRoXjn+xxL29XRZRfhbDXUwZ
e71MEYo6TlHWocstrND/EsOgB0KDqI9VYQ8xVhY7W34aRH6KJDhTgAP+j2yAtExD6dxd1pC9h/pJ
JyzYx9LmGS+wHJox+vVADKvJkEMFA7s98Zz/94x7GM51HITyJIqBn86NLTPgrUBT6WmbAPSrS8kW
j9E67+9JKj2xfdJB7osLyl6rf0CkcxD3vqg91/OhLmwULvWvUsTs3ZkZrxBD2V4FWxnELCChwlZG
zrsLWxS7vtoWmpIn224L1CNu/nOclWsYInvZm2kk54YF6TerBIRTT+mp7mY2RccEZEJmP2y+upxo
ftOXyHur5hN/C90ZJdCAkdqgYy7bSJo/JvNK/I3bnHoYGbGGZ586XAqiH8BSAv6KmtSvufjEcuxv
2UfBtRXm07dxZ9DNqETXOO5hUnArDHy+DSZYVC+HVN7A+tDlxrPhrjZkzqZbeTjrnEU3rymNRUFw
bnb8IrhtDRpjcI5YqiBYad9e/NloWkAjVsklf/S9Qt9gWYoWtYNBvDL9gR2aVNzc4HWAxWTQqRgm
n7RqjGvhFLwUJ3Qof9D97uTYsPfJfyDT2q2z6E1CTiXsASMncNrbBADOIJMbP3xSlWC/7GbLYsys
Ut4uANGbD+/QPYP8I600rJh3VkG5hUMys6UCQaO4tixxZi+N288webGk7+HGHa2jRKzWd6eMR3fZ
zV6PGm7ZMwaK1xQeASOD+lpahpbqr1wjrgT2QBw9xNGfpedkEEewf8DZWs2ejsRf8LPIIfYisDzQ
gJM/U40qL3rd258Kh3BXbw4PoCms3CrAcwKAqcTvEbvU7RaJW5LrD63GZL+J0egExbz2aDYxXiXI
WS3ORHY3QoiVq8ECgEKaex0X5cZeS+O5GZYGivsn1RWQMhf0XA0OcFC9427AWngqkZcHMo9SRelA
YzTWbRno0Tci2jliyPUaeEtWSR9GQPXrOYBCQmR8P+LfmK3LRIDI7ioySbtDZ1xKZwgu8N4Tkn38
VGPi8THDHSbtxHsEICB1XeuchbXGp9Ww5DVimla8B/ZMwiBblF57B7LNaWDL1qj8e37w0vWKOKQU
DXLHSLFDgL+iiHYNMwt7LPcfDobDKuBUrysSpJeythx115/wU3zWWZe9p1CNj8i3nOT9T/Eqle3J
f2qNQ5mEC+2aSxiN9+ucODzLIjxvGUtPjl8xQzI2OsBgg2ZBxgRXK3A3VM52IkUGSEWjkUby+yO/
12e29ybqkb6VUBeSO+xhYdfzGxH3Vwc3xOu0+tNPeCUysTtRwrCt3OA30F3+/GWih5y5N5KKv8Yx
WNBpCT3ABVd3pq8IJp2oJwoOhFIBFzE013l0B1Mj4MoJa8mS+KC3md2VTC55GQoRdZg+OoKmMlc7
cx1Z1eFbbhBI59cdU7/yEj3BE2werHv2N1IFoJGCtX0ZFUFLzM6R+Z87hE7g2q2BqVE57MHkYfY6
FMLcBKYBMFzezfWWktOsJdBMkiu+IgBEetYPdPhys2PlsE15B3m0eaX2+EFUynFW5FSkF38/C6v+
p3+KP4Ki18TESBZ0Vgf/OTnCyUtBAveGgQ6oRmP4wnQzyaDH67YHxE6BrKCx/3rcS1ITjW64QxBf
TJsyqklX5yEM9E+M+FlzKdfqTwJYyniWu3CK3FQqiSERY/CSMDCJZ78DSlwIJXJkF1bhjkrgtk37
bFUNYHMLUQbNrB3M/FmBGgdUoM+DhTlqnLXoHA1WIC+J17jKB+l8GaahErpaWyOlB0ctamWLXxuK
K9DY7otWCqVa7FOwJggHFR/XRhKifiH0tn5Ge06EXATT3sA96Yznnpimscw27wHRyXbSd2EZBwLj
M34eCXXVmrFyX22rWwbGBofIAyhmjvUJdXnhj3RhAv273xk9tBzABiyqB1naGRbi3Lr0GUCuT79y
SwmVeF0KNdRaPSDLWoAQTaJWdpQmzLClPM9OsV91G0e5QeMBbqGj6OIlW3hJr8JFbkm5JHrpeoo9
/4bnoVcHi1DBnRWyoHbjmhR798jv94xucYVyOgpwDJ8Y4C4Pwsdi2NufqSEduX0C02n/fIVdQiDU
2fs3W1c0cfm64JGuJxP7luo/LDz73MHWGxZvRNffGyx+K0Und/8m7xlmmctZpW28svCUPfaIUjHD
3KscGeAMUNm75kk/DofkZFZSonfMw4G52JHMvqu+PQXnK9WAP3rDYtSU5Fsg/L5kWtjqr0o2D+7E
rhbveuxq1O03AcbeEX4KtevtzWor8LRmdCPV3dG6GpkIWRnlgrim55q12uqsPphuKu9Jj7kELWsB
7dsXaBTJCwH5+NLx3aN+m8c4NcL9bLG5+tjTHB5G8BR0/sryWBSYH+op1bbo7mMySEarg/aWv950
oxpd++UinK9Dq5mtSm64CCm4vOjZlGzqNlREofnhQYLjB+ocv6RL2hGZNGLwWEWcFpv7KOcVoxrW
Wz2g4pMrBwY/onNTfseiLyRMn8Ly3+I6a8m7njAqWtjghO0q/eh9xa1sIL6ZDsqBDDSHnO0wpQk4
U57i3OaU5ylUnpLgnx0a4+zkcYF7opdmkOXL2+/ooTZtldLnEnpe2Bp9+LDXEQnHUyfzllhgXymd
4+BWWx0OdU8S42YpjeTyrylGPx0oyvX0Q0pHKG83d+aMy9/JTyzbvsUvaEQNwunLMGiBLZqHZ8LI
k7Mrl0HlaNCIFKDfn1miXpFIMiJhvZF994jSdOblohJaiqtLGfGehue6fahap8RY2MWRrUnTHQB2
S/6csW4MY23g/2Tv6tDt47mtmbRi53VrxVA3cyjD/KPqHEDdZJ2rnSCIVCyWtVw2ai26UklZkXQ/
v937AR4kMSd4xr7xPJjmtPedfuSV0ShwXjv6TknDe0rfyLEjnS4JMJQPht+XSN3QorF/yE0+5FUM
q/0YV0fk558HuT+e68tWVfaXxACmwQx5zFIBW6B+50tT3U0aUm3GFZkfi1+Uw6NiHW9HGi5LRtL8
xShKIohw4WV/XYqIDf0o81Mw4SPfumIyl3Noa6SNVqP2bIRP+EFrnE/3OFcUS+5TOCOy4z6wmDzo
tv9Zmw0HdhW76eWkbjpDtd0E9YqIROhvTQfSno9Xdi+iX50WqO9xTine3f50WAix1bgvlfvz6jW1
1s/UPWYio9BJyLTwuZUCl0nmEUw0bioG08Y6x25/aZZO5i6/IjaO6HrWUnD0zJOBqzMHanYCQOOq
4/eqeA+bGV7HvXuaM91MvfD8kP40WSZ6hlrTtdf73lzIqbCLpjug7st8oGL25Fd0im1030KxQxdd
UD/ff7pXlbVu+Xb5WAzulYOUSN9JGIP6ayHSocfwL13msxlURQcOH3jPychtMmkZFxzS0Zw88sYm
yFs6j3GQXmidSKoxjFwy9wCT0NfM5ZjNyJQTgH4J75E+v+oH1ugO+eARFXTmRF0ux7rs50xN0XPq
FnwH1pAgYi/TCIrvP7bW4ou8pz/JL45wFcDcV9c8LB6Jlk8nBLdWuVzVXoCI2r94QAU2M0lWmHmy
WGPEbA/X1Yoi3d4f1l5KfQniD+4dpVqA6PqDWj2rYr/Xr02y6xaw3uHhH/jzr+j5A5bLWqh9pn56
DmTBqsvz/8XG3Xpb4KCtSMvMipjOo4UEqf4CUjKBw1rnvmmd5jro/EPAZXl+OZFBGe82PWtHx0Rx
t3VMJv+aZQ4GMOtm8oy/6tU3tHHobXfoWwffUXJMzGoXQX5wUDlqzKkhwmbHIXnNa0cIB18wvv43
47qVhMQ0WmHQovgH3sC/6YEth6BGAdPGDni/jl+FgvU4E0pIKwxmsNqdbBcYK2Qboqah7mJTvAfo
FHK4qBdWVkGL/KoyNLfUskKpQcHAtkIUH0x93x99Gg4JXzIfSEIKbKyjlpNvriIT4TU84vlaEhE0
Ee1An8nFCWatuhu7WhNfWf3J1kXOHTTlAw22CtoDv/y5hyOMPLJDBeTdYwZ8DCrnabG+43/Hl2Pt
l94CQlCdavcOL7OR3JAJb+WljJY65pIsMdVIwMPnk2OZMeA69cVdBFwPKOSS5ZECPBDjN59SgjYM
UouFh7BbH5yknFr7ggjJ0j23r6dX/6yoIV/9Md0k2997o8JmI4VRsOdHU7tJRsmAAaZ/3w9PpHtn
gHQt6zYd8GBL0UhhYlBfmp9R2gE3KBtb+IyC3RzQJZa4x0S/8vTeFBbh89VQ7hWzrYUwfy7gDxhc
VVTommo+YZcaBPnpcwBfjylFfSB1J4o2OKldyXvVeLxjMTnLTe+6e5nDvBOwVzJahpbyeT+a8bJ5
rkqgDoYXLGWAs/HlnbMHQDCAOYQUwbTU6QaR/HLiuajf8XOKT2GYs0V+5Dqk6k6sSNCPcEocBux8
25geA9VjJz/1NWiulBuZowfOnzsRwBebO2SYwnpt18bWj6Up+ikLfulUtwYur2TFaOyWR60vurd0
zfL2bgjzIXqQ7hg2GxSXCHjVEYdmTJdxE0fSgBFo3kH1dkZG27EUV2jIGy6RByqIZZz97TZUxGxI
a196tpFbgohVPO/TMNDuD8QA1q0aXCFhf4pVeVcfvm80AvH92pso+AXN8SumITN7WICD4FNZMu0l
dsLYvMa4kB6aZspi11RoVRIVfNX3qq+tCMfy+DPSzSFqjVSd2W9LfADN+H3akgo/vGy0JHjcPkru
fvSC5piY9vC+bntrn+oLm/jFm2s6MWn6/S6y1KvaRfobRpOtvE1SPcqThYIEpEKpMYx+YpTdU0I9
HLMOMpZu+76XHyT622qf+/Qp0uSbf9Lo3mEp0vNNsOcKc6eai8wZA6fLeAYIs7AWi5xjoE8hFVJA
aDHeGdnzEtTxLfYhv9/Iq0SE/JilKCHWu/FkPf/f5H+h4X6kNbIaC5hXZoV0smzytFG+skd4ZY/L
9rYW4C1RAeYR7IRHV47HjGAvNlTvcd5oL2aGQTU8iCzVYYXxb569QvX+3BViyn4k1psDYtgiRtUS
KoG+MIz6Q0VZH3wjtXwPHPycE8xChWlZSlGv/xJqxXDOvpcb26wnMU3ILCieex/r/jvJ/xoRp+E1
b84wlDyHKy+XIOHKKKKTBQ91+Ai33LdbFOYlLDOQT9YSuWr0U4ZcLE4i63RpzEdgeqkvD8S703at
8t6B0tQuPhBO4ruABb0YxAA/bMFosTF1nKWn+DgqA65WkmiPD6OtmCV+tbciVGrVszxHuLWPrCLW
ChfWtvmMYRtE8sg/+yptIrdrUVXvgSeY9t/Uih3QRgZLF7F1tasRgbDCQcyZBD0gDZAB9kWzm1Nc
lbnMm2fVvDquNALqzVMs04ds7BOlRKwpSwI+yxSN1MK7I11QNbFdqQHWzmTD6R3yHHf94NxsRJWE
JMa08KqMRPhG+PoT08Tycp5i75QaeI2edwtHyDtbWjklKD0VE43n7s/kE7HEVEjFndejPqAVd6vt
OKKwq36n+cN3BmHRjui/PcZKFMjhY9tkmDbC7ftE6MVf58G7Y6sUWIgAvqriHrGYO88K2R1jQwHs
ryxGfUEdajLtPcBFjsLcKg2QwZLeKTFW5SQVWgS1ZoqTx0jI3Ws7KQFkpsxr72m4qhtCz9XVzw/Q
sKjCq6k4C3g+GFQ2JOH1NNE8Vy1OjTU6sADIFlsHNRgnZqRiocgE1aSTE0MORgNkcd71K1znLPI3
KFv8OhmYyGHFOTZ6ELobPU3ueMd5LUUiJFq2INtL/M9Vln0XBK7KyUmzLBlE05h9fRj//OIn1dYD
l1lrVtWyi+Gr1IbxtbzFYGm4ESYIhKy6zm8Oa2/gPoHtgRLcMrA1+CcekHSn8UiGTkvBovOKmUgT
IidnmUUjRUgFLIr1AzGPb+xy8bdtFT9zzN93lvxp8sYsI4r+QxTv+hHaMYt01/GXp6ko8y8ifTqD
/uZVczYHgdInInTAaS9iN6raDRoRLCpaL66WRPqls+ClBDf8Ws1sv3YULvfh84scFaoOxKyzFqO0
dLOs86h1zUMfiGlZG4RxR4qBZV33g3mb5l8g5ogwD0AUBC9JWAsLXuWHyup9hkJjpkdowpIxe407
uAO8osxq9DbE7kLz7+Vl2h35DwwiOObnXWnga2seYPkRnqXrUfVwEfHA7VkPeep37bjwiB6IEjpw
Ar17cudJmg6q1Aeqmh7Em0MOY3HHyrKjxjiH4vEzIChbmGx23gTNObHPGLwLrOyJ8T1eYIvUzAPI
mHR8S7i4AjrjsWzifEZjXNdCXSEPH72hO32qgNFtoZhX6ehUPoxUcZChdGvdyNe0A6Hat2xTkQCk
CwGHAfnoJhWKWOPiW3AGzLNfTIOkRP1sOjycrBbQL7QxR+qYj1StKOYTlPB89qTBwIdNSxKP3sIj
JrjqBd2tWW3/Ed2HWzjRftG/g1JvKDIY2WR3HkuEcIV9p5kML4AZaceI/ESzgeTZ+HKto3AMjZh0
nep/faeMJUZni7FaPGBabN+KJPLpxw15vIuqbDkz2kfRzGXRLiMhPoA9Rn6NQimGp64wnMZKvdt4
T4yI9cU4cs0NKtqkQYQNXwiVAiJfAkNPg6dUMPrLcH3Hfo9qAgunxpb3yMEXOChM9HBZ148Y1D85
OTtjtDTz0aBtf9ex6dbXpipUMYQIP3tD5cbb7fWhdfpQQcgZBfpTOwIte3q+06tQG/dn1NMG7LZM
eqVyiAgpGxgCAfOhbpsOXbhF3bWYjMmlGa953qK2PO47TUt96X2q7uEnREiA+yMEfqiwzFWQm2pc
5RXssbOkFLVrGKdmvjrb2dcAwe1jr2KTSpypvSyW8piVUKH8qo9HwKI6WcAk12EGMhzAMZshYxSv
U6drKBjal+mFVa28wmMADXZ10bgiRK3bzcX+g0+gEp50fP1XqmRJ+1V539dmU2N1vC03yrY5DqjO
zAvAo8M0fWvo2qthV3/v3hmRsI8sCxBgp9ZZRjo4+567RIaxOvDG+4tpU10n7H2sL0JSKhxuLN0k
Ak0xZlrEij1QjWKXSAkCACSBYhjAoW0Snh6MwA8qfTXwU1LwyyWcaO9tD5QThjGJcnVqvW8RKCUH
eu86JCnzluZaPkQecBc4cR6xDRGldMQlmMygNr3u2fs2WzLneDVuk7HSCOuu/Bx9vgRGJ/41J2t9
DjudISlmqll0SUS+c4ucDIHOC8ML9VB1krzu2FF7PeicjQR89QGmLsQD2SXgtuzRTxA5K/st/cTe
04TXM4+m/RXAjaCO3SVadNHKY4DsNHgzuQwGp14MM9+cfht/nbmpVeyBhGtgxFhapL3vwE59o5Qb
qj7nJVZkJyOv30NSqfN8bm1OOiU1uj7JXdzh3m25REYYAZNB8K5Aq1B1l+G0RulzBII64h5LfPzb
5a5KGYcP2swS8ZnnOVwwYgTrqZIylc0z4X17yK8p3A7zea1LizOjWpGMHnBRDHjOoTEvMCvO8iU+
eno0+pz5canyUTdonc3lzi1XCh7GHj+giWkMHLXefwXQVuJlbT93d2J/l/tK/EVGPRDDY0KEz8jR
cEj8nkQwKReCsCEasloKiLpCqdzT8Js95p+5M/FhLZJPckOsHoX7YgISxMgYg8Mq0c5FpvRSYSkz
eFl49SnGgitHieMlr8foeSORf8vl+qbaQej3SlU4GL3bTHXkUYsXw8SpkepWeQ4VhdZk1y9SR+f0
Wffz7eVX2QIaOwtZDzFU0OJelZXlXm7mTH5v/fUfJ/w84f91RvlnD7lCJIaUwo6ncLamHdkztp9g
VBieKhZXHB0kqRYtaLNHeb6LBjEU1bi+H2+tmOmyg7LivIA+CwCQXS5aD5mlgdxrKyDD6bT1DVjJ
nxCgjpl9wCVBwVmHNTDz+LitbAjL90zJfjtDZYLkDdcbyzc7i1sykrdac0SEuIjuL+NKLdX7JIvO
csfyvSrbNU3zVJONKHqxqFTqUuhY/XB8EFWJ8oeZdlLMox6HfzHKnimDXI4aL3SqeoxqYbVFAe9g
fwgrMnmMbCiB4qoyzRq5SeUOmOXWxJKW4XVvKrySGS91jMKJAv99kyYfMy/cD3cc+vA5fcXUodlL
bOcAsmqqaRALTBcmEGIYBVNmaN/3YPRehn1rgohDDE5OVe2fWykq+TRmDQlq4m7rLsebVu6Uew0Z
7ijf+Qo6u8v6qfeih7uDFuOW09i+4YZARTqk960QUC2GSEmLEQ/iQ8UXupWGyQEHccxzIpkZIRmn
mSoB/mDPL6cz9huMWudlivJ1PrslHGW8NQU2BTMtf8VRbntfyWofnnAPyDMhqco+Mvp1d1cg2w3T
IxNb3laZttP7zObwLHqIeKwARr2eyRT87yYZvrqqhW5Mg1+PU8YSGg3/HRA864EO6gC2+pUTt5k0
+1WX3++/vZU4FzZ6VnLQsnlg+El019Eh9AIY8NsQkDGbTwwCDzpEuautPTsDolHbT3V1n7fAkH7b
6iwUU0wd9Zhpy02cekTVOnrB866hbgltrd3uYGgCHaZzBsP7KmZbr4FMMgxQBzWkmm/3UkVRyDGC
FhznFYfg6f1zLCND+mf5sQp9dW7CCjnVE9Uc4EVy127PwfPol9sKlofeIn8Vzeq5K+OArhhgdgaj
g1vocQuZVUukd5emNucahaZ7+cUftUzJokeIp0FGM0OEC7LsqBUoBnQuyD8PNeHJ8GP4MGxhxojR
CuTZvtddDuCTVeARsjEQYM1NlUy3BLiEeofy0HGtGlRKq+EiafwtyHnUyAdzNrDIjASF+Sa2mwXa
yT+E2oWF3VE0NsITKxrBYaPrWuRJBYGSGgltd4A1+4PYeV7njUqwCoCs1coRLLWdJcBPs3RAm52l
evtfyjKTCbgeNlS/WyO5o1RrJZraHciBA+9UdYa2bYHVFw4AL4g2aOClkEFwr3UNLjY4lV4u5o1i
UgN/FDhb1NHXQWGc86MAU4M2CZqmggC97N0eSJdDq7u0RdqF5xpLrjB867ziLJASxhePcuQrBuh4
esgKbfuJ1NhitBylHfv5g9UGffjpEEca2bfefk0geZQ+TgHlhiKJu40M2wbHLrHQ5SLq9pI1Kj40
bNJhwpUmc+7V1Q4dnMA9rHk944fR0xxUs/iJzaVCEfgMy1aRYndnSNNhuevVbPmMkExngyhukCy3
/GUh6croHN4wfs6OWiIVvKC0Rc45okweltOkkaoZsi2GSjPuHckTHmFRZ5hFLmgEwZQStk3jikyJ
FnLpAvHA3fCfutm1YeNowohjJEPGx/eqHW9Jlrw/2k5zjc1iWN5r7l0VH6SxCFWZywsvq9g4aQQ0
TL43WG3IHpK3fVLfcRiik/1/4D5V1hNJ82n33roZ86HcF/pF8SDcEWrxgFuzd94fn+LWndg0FWIc
zeUPiFUA3ycRkQ9jDEeTx9e5gUTahHCDPsB5NkSQwK5faiaP/ZWgV93NBbu3Ib3z2JvdFcQTpkUy
fhT+OKDu799bAnoXHvRKXuJai18Zy5O1WD+/Txh8bXS3liaZzqxKVs8IcNwCBg+jKLdhguLq2tVK
Gsau/6oxDALQ9a0tgrlyHh2Bn+/wgiAQsHyTeMl3+ACLJWku6EXyToVHR7kigmoKLF8Rci51CbUB
tWS1Uu1y6FE0PO4ZTAJl33bDqb7VnLKLLpKu8w1Va3XiglQnIu4mTGItMBKxMAmq7sk8UaNdiPc7
xrdWfxRoTdX+L0PBQdqKkl4LbV/ihJKnI5aAPKPy2B1i+ErvxNzx3xlseMCthO4zC5pVXWVKFHmN
8zYgpq+5NRMrOClPSmXZMSJGC6HZMkR2SDWICRf7phwYs0uxv4e6HXlQla3YMtv8kO5gQ/qqU0N3
o3C8JHJzeliRRuxDidfcILj/m1iq4qzBaHtWTGNJWg2SA4aS7d3Y/AEgzC5dCd0XuBuIXBC6zkv9
Nps4tJHtDDFv0N9YkcRDfzvByjlaB4t5vyVAeLMsUOQogeWKUWhj93zolkCJE+XrW8iwmMIgkxmw
ikAmJaFdcCycj2BCEmZylqrouCiRGlHWVM1aaDNJ2jOZm4tTSx4m93ODLm/C9duVpsL/zf+0bXDw
lmAUU5qTgOMYHHZGoHbkkRei7EmCoCxKOiU+YGshgSghBj82/4BOAmfXV1FAKlkw4v0dEEL/SRfP
s5AL7mx11o2DaEwS2SzbmKKnc5YcN0dpJpR6WtUlqhKaoiuWOsQF4UXzKo6VvZCiHPFe/DuTQwgB
vxwaNdF+KdeadAyZCjUSOgBOxLFEjWzzmz+Xe3Xyv1U6GieLwRFpuVpNg48AG0Gl2qtIXvRDw25O
CHAY1eKMCtKmdV1N9tHqvn2/MpHXAod4wSh9iY3vpCHbN0IxKQlL6ydy30JA6SOF8UpDe43UpzQ7
Vg6fQby+F28yh7gme365omJD1b+zuBv5h27V/PP6UXxNAQYbpiipa05ISmlMcr4NYEdoib1Ip4Ze
dvveZ05ZOK6SqnWUFtnn4ipYkIYm0xg1j4TEEQZKxUzgG9wTy2SE29s3zzr4EVSe+n4M6EDe0QeJ
q7FWO5u3vXCmyTTd5aWGt+RSoyntyR3gsxPTzYV5YCrciAkbjKVe6bh3bJgOfEDTfx6B6xchhLtN
m/TqlocjNzd6N/yWpAwJY9yb5auT0jNhdH1KXv5ofXih5dQZyKhf/2Abwo+mdTGVTTG4e0ShqTkM
ydbbHBe8eXXEEyQyh0Zb/2laU94oPy8W+aEyikNsbxsjKTvn6ikhPxGglUGI5W3v/uuUZLt3c1rx
BoXrfXQBumwaM9soP0aj8T5NSs5d8eX7CWSpIqRnJPkOpvlBESyI/GWPDgnwLQARxEfdyWCrEILm
emxWy7SVMHrxGZSy53XCtb4sPeI/pc5MZ8y3pc/TD/KOB29AcXx6YjB0PWaxc3QGayocb4AI1778
V8dC3Ba8vSZGSVpueD9hQgI+Eoz8vpdRyCuKRNXU3Wg64XyWnZh/+kj4a2Eb7+Xx8EzGi9eBzINV
x5153cGl1Mas8wQGRNr1lsrlRxSru4IjcIocQNB+F4e5oLtBpuAv+e1e/A2kE20IuA0utHfmAkH/
ISupTN7ecwRLKeJQNKzDoXCfhQyoPi3K7I7m/kPD69JrB31UCN0IrVOPomnabEgEVREQl10nzAUK
99OQuPdOQrHyJ6M0TNxyscCHWLiY3UXPYA8PjGb4Q+NcfyGPK9oQXn3O0dDsySq7Z8MaZYeGfxCF
NI9024fSAkpyNNPpNLyI/0gPlnDwV8P3+iQBD85Rld8/xSPqGTnnaOcQB3PZTKeuYGZ6krofVNRh
7QZih8gjdJ1MeDMGBzm2uDJopk7taeaJgjQqKYPG9YuETIKA5SLXePLj5L45pOKMfCr2zBjaPAN9
yE09yCSj+7yxHQ45AdANbsM6oZk3notJ5UxGhjRI7jgAPkJ/X0B9QOaaP15VVWdFidSuV67o28RC
LetbpmEdnf8HADmKuYTkQ5rqn4SogiKxGZ8/J+B24jim7t3lZGs0hvj0+XuTbquqy+UzHoPcfOyL
ObqtBYNqdk0CVoD7+7figYw5AIGdq+TM5lqqCvjVToq/65cvVgv2PT7Dn/VMZ/fFXsmyKWDppNBk
nfs5eIgW6fr74+hullQ41BNDSAOJfNyr6n8OJ6FK/Cg1buZHb0ewp9wRWUlDpYoOgRvmgSHpy82H
QLKwlyydL83fNbuJn5Dm/sYEKUPyCbST2uesQc4vKnCb81B2g1wMLkwrMKnGpbz8hElv8NpDdW1N
doI0ySw77TYlFvHcJKClSivcfcje9S8HX21fdVkhEqRDKxw3Fdpw6qeMFF2bKNp1IohXYLVoqUJw
c5bNzwKq2cvCJebVkUknz+4IUol4XFWJON8eK8NF+MTg2FIuPJ8S2MGM2fIOmJX98wkDeAxR7ZK/
YAhUA6KRbz7ZiJsXYVWvo877/y327RLiDvkCw40Ii8iO/3lhvIU92acIIjQIH6Klomjj4FdL4gNM
mzQbyMX95hFVOnEtvsOcCI3gRmSN1r6Z7rhe/E1poiWy45SBYzjbLk1RvNDHkhu8jFuJjOBETyx3
QomtoANuPhFvEk7reD875XT0GRi8vhj9/0IitV57dyCSem5jxKlYpiXVyY5uICdSzRt2Z8iUYeNY
1TUtmhmcZIemjC17gOCY/NyNPZrGfPdSBIZWLnGyxYVUu7oIsXaOIbz3/SbNQkoORzJ3JJhRS0cW
kKW7V2JE3lSH2awm0DtitZl/xYkbyODoLmsBIj48wpBy090UX7YT8iDN99ROIg1SPAv0fF2RJ6g3
UDphKDIMUhKAYw8l91vK6V4Prxt9wC9eS+ruwh0uI6tuX7hLDNS6YgylQuK7MiIAcz85D/A/J/pj
0idwHS2eGErkbFIkUPBgYWmg5+CpTDTTj4KVHKBW8RBycOn9IqNpucCYW/6cISwPmPyp4TLXPFRl
T1cVvEB/n2JQB4HcuhsRiMITkAcLhDabsEBJUNSbrElBI6IMuzU9YREBurXr74CB0oh7lQAvL82/
hoLlGUKVsqKjh4Mwl5EFGJIqAwUqWgESHhEkgrdvVp4kFRpoWxGY1U9brzH9rvxJX6RI+yNducsu
it1VVeUZ2EbhTX7jkkTnx441XLiClk9iK7Ki2phK+CwFZ0GQaZbzLGbmGELZcbLoxqnngASQIGjx
h1PtKZWjF4TRA7nf1t01o9QKFlT6LGPD6EsRXqAsU3BWXCPic42TOdR2WikWmMrQ1ezMdkyfZi2c
wumaxy3b25DsJCNPwzVvOHAWo9STqQvaczyLN5VqWdmi1JylqXZtxosex6925/i31vNUAaqyz5yx
zsG69soGEhp25Da9ROaS9XuhAxSxSUkwrJRg/zw1PFjZbxsPvXSVmtVim4huwAyTpNO6M5FdL+FM
s6p4x8pzolnp7T9ITP0dHCfuIcIxphdr/wQjVQFCILBeG9rttHrAYwyL6z7+2LdSshVvgrUSVNSN
TdZjIVZnXIHhV3yGIuQCnVOGOrb6JfSr1YiR99XFkIVgsfpV8KCN71XeNZfQQCczv4iQzumbAo5p
5f5viutv2nb0jFxrMy1+GcmXViI3EPECvl5c8Ce/py5fnSQcVrFRBydyZtpcnO/GFpQOQA2jqDe0
YhxitDmmONT4kOqgkpptcdMYMaRDYu7AKE+atRaU9HmfHs1shxbYH2k8aPZwvlpbRwI28QTmRvDA
8201lFq12B9E7DtLs2qNNjumgcLJLRWckPxYEvVHLMIlZFl5mPZfYqE4IPSFeZZmZ1N2DD0ZiKjT
XfIRsobxL/rYP86XAtBLRWfqpByk+eHvwSsnpEFe4ygQ5HnjgSywF8cqTIOaFnsesPeZVnzivsm6
zFIZpWZTOWGX3VTxjBNrXLL+C/J2XsVy33Vl0FLWB7PIhwOmmrlMi8PxaJl8/MQnLocRy+h8Mzci
1fxBa4ilBYWJe2ayAHzC0HI1cyulGux64G+7N7o4KaSu26ev0NMdRMpWmnp59pOAL6KqyaLeWL/E
0hmzTTFOc7HAI85ZC7PROnMAvMusEWnpYAslazZwU9kfGOzF/n8VXFK9tYZX2G/wtSn1Kh91SnNF
Et6GV08CBO+OUj/5tRNlHTC2WH2HhIF1leRhAblUH4jd28hWzZNoPR2SuquvpT//Ip0E8biSDkXE
mJciz8q4Lf/3BEVMmJeZNz9JnQS4yfzaWMPMBXjdS42f75bSiQSTJqJLOwwEW0G36JPp0ipjM+a5
kB7oo/1aXfvQoEyog/ywZTPvQUTuyDk6k8+EWP0xr7R2gfJpF64GlBaex4F+NJc32a+cccId5jab
ijY+VrClOPamYd2rMuOzdmzYZLIBOsPbc/XgSGgxPAxWA2lrQj+9I6MROHG0eRT1m2sTu8+s2cF7
9bS5ZAQqwFmzMcOPkCiCxnFmxxPA6EmTsmZrkRCy1V5UbnuW1UzC6PliGHll7RJPz7TlJOPWad7M
cHnW/O/7ZJowI3Qv+5m/uzd0siXWrt1Nk9qgX1AfA9OzIAXiBKTATdkWbBdkhagYcp09eEhjXlOJ
9gUP/8+Jv++4pUJuVTt3gd2Iaox8pTRL09x52X4fJoihQkZYDg30jF3tiU8MFF9bDQUh2otFY/Rm
W88BO0e9e84cgTZvUSo0laCeKZTUHEnHIjv9yBfLhRsONY7ImQqLqD1VR8F4dXg8Q1/aQd7Xmey6
or8MCt5sPwWL0rFoReGr7d59iqDzsOVVE45L4/UHbr4yiWTGQfLqdl2duppsPZE7OXlHFl5ywb1k
E/81PctZ/bm0TraCbzkKI3HGYllM+gSD8qB9B7lQ6eTjYTjDDPCVikX/fhHCfeUWycnPZLxgN27e
5iQW6a/Kg4xolAshdZfsYyix6i5/ObjHOpTodaymEQyq46Nb6H3SF9UguG0mTswZisaVmLrMxSZ3
kcqUQ+Sxem9+OgLKEkc7Im6Qp1X67rqGGAqFtA62WrqMvF5QHzWgxaJYI/wDgWoRnJUPOoCGDXG/
MSrfe9+Ns5aWa1V3Kuyj3UrF02kNLceIDvqCJL3mx0VN5Wq+/70vAiCwz7j+4IwYvlFrdQ5wCmTb
DT8GGzfU5B93cGGvfzuq8OsQgcNLNDqV+MlOm16swk2u1tVcYbdJrUHDA/xhuHr8NcuGZglEz2k8
A5Q0XnWTJ61XLh5FgXYD1RBigcbLKyAKoHnX3Ryf2j9eLkMHjWEQ/JNV6TRntCl7MMTTmfdBh3iJ
0pd41rXQ/EGp3qQzDjJl5P+xWqCWmO37G6a7f9dHgE7yc5x1/5DxA2Y8SomqFTsQ5/H2lwMuSSoG
aSZ6wE+yQfo93WGsMKsURgnR28UblywqWFA/lqBFsrKTo+kkmLPXIwNbzuqvvFKLb4Uh9GrnlUUr
9qwSaKt6KM1DPJ/GVVc/CXjDbtAb43tJB70WiGbMav2r5fW1KVMC72DnTgvoi1ECxaNqO23bE76k
AXF/OeujCVOEcCiUjGcMreEfcC0hHVYxHmXgE/2NBay5EZMdSgYsMKoGXlaHoYOPFFoIQevuaC9c
wt9jVbH8l/yQ0yaFd8s0b0tDD3jtL4e3RKxvodTudF6mEF74SpVIvfw+h+LnNAKyd7Edc7IDJ0O4
fBpiR4JLhFzo7cRh8xwsZguNXjBU1BtDSCnxMMVREh5sniW5JZNM4IhUFvv6IxR9tao5DEp/15V9
qytv7ApJuGrRVjFhqEoeRtQ015JyD6y8XoC3Thd3bSzvI3jftYjEW+RkY6Pe0OfjDkoktEOg5qDX
H4Uq5SDp+XqZXOdobJLtSRbC7U0l21Hb1gc2M+shovNVrp/JDo/wN25lVg8S7b3RQ1u68Mle5yDJ
CZ7kUkLsz71m2aczVaNv3nfVZVm3rfbqClbWR0OBh9/SDBzcx73BF2lvS8gLzjsGT6eueZ5PMCOl
0ZhY94YtXP6twVs9RO6W2jViIBeiW0FEr6pa5LSOvp11ZL8qmuuIsp+s/zUI6V62U/+1uX7ZJSUL
Y5QWanW9HYzdgDQ/PfjV9AVP0VgsF1hEdGW/Pjba0wz0y3FsXDt1Jwb3mTPRrc9c12XPCgEoxvfV
GEYt3xOj+DAPLwH76rTdtnxHRoHTkXGPVD41il0MpSgUCb05XEIk4xBnaxSU81nixrZPKw3Shnid
i8Vf/D4KiiMCy7D8odjLMLK4Umk8tj/8MLhCc3tCkHQnlQ/iDIpm1zGNZbWuJQ8c9wVhiELKhm5R
fKNs/d8CQpBgNJir6UHiwFFaviB5o3ogXIG2IZ9kmzr+B2OyfPv8Es40Fk/FZYV4OYoh9I2/mkTe
kWR+xIIkW0I/xGFiE+MbpfGOt6NOZbcUfpdD53ylvCD49rrTfoqw6uPl3P6tYWyCYFtP/Kc0o2WZ
5pXMmTG/sI+7clNi0uYyvlmRF0YbCxyGDBoDgpEb+d7w18u/pPGmVSq9twp6/aIGfBAuMjZqD4wz
AHNRmQjfw3CVVOvI43e6DXOnStr7bRCgWo4dBHLrdeD3Aq/DVdBs4mxbe741OoyCKoVb8z/O2ywu
OFKGvDbtU7BIq0O/c1sd/ZMrqNsYlKYRXdHluahpd7ETYaI72mF54iy1GtcmEA9U2drxFYygHntX
+EmJMN6f9pNy5wbUPkz6IZYAoLjjshbaXmcwb63L4njC45/xmpRFVy3dfQ5JRZw7aaf7BCl910kI
ojEWhwdgnUWyGCUsUPlRxNxxyRRCsnTsWD+NGYyeXUsb+mG03wiA1rmHKaktvnus43uryGxpKrOD
eQ9ehD5p+RGByL98tXruS6oFL0wz4ZpWzIeXMfj/bdOh+GflsMYD0+Uga2h8rCFwqjIS7v74cCDT
87z7EXozffxVH4UXI2y6AIJFlxmfo6U8f3eXL3duM6eA6RmPWJe35RdeuNex4qHsdnfbxuvqKkQW
nf2gHjcHQ+nYby6nHDnI7cB48QWFwTWt0ExWPQJOXSZ8eG7wYYmAUTbwnNxmFy/Vq00guk+9CS2l
ftHJbUz5m9pA6mWSCa355hv5qmhp9uDOyXqzhpdpqH5AIRGTIu76ZUZoT1wKhkLyUO6MBkUa8ikl
IuImdKKd/rcu/0ofZtvyqph8C+juPNyZKlsCRj0XiQatfp0HeH0xjYM0yehnA20p8SwCCZSwsmCu
gbmBr5rxoVqAZTQjX9qQbyhtXc6P4G4DyEKp3h80X+YorkExsfruJEihdIlQt6J6DdAu1ILRMHFu
Iz0JVratPcLIs2sDXhSe/Cc9hroo9SSvU9bhABQ2HXWsrVwata6ky0jvliJOroe/wvXKj8N59jVN
BTStjZ3EycJuBBBijq2GBC5AFZ7ZITll9wKOsctqKN17mw0a+RVmT097obU0mJbMmsjaSEtIxffD
EvKvGuE/urzN+IJIi2xohZocAb9ypPEYMQd61qnLQnu/vSwChI9M/AoXz4fJbIOouyFVhf4apwiz
pU9/bw5lvjUpvqzc7VzkbV6KCIpuyr6i4F9ajv1UhpEof1jwSj8mP6KzHqTrLn+HMcAS5lREHMlX
KOIhdlPQxA0aD8nl8mLqOnt00joXWwhtAUOlywfm9YzIKpTkjogCQyzhbdTF8tSaNgRfzeB/a+4Q
5rlybSDSMjPrGVQiaySZuzP7jaygluiEy23h/wVP+PaT9bGUM/6ezVxdogL7Z3OWmKPWRo3gkmyQ
vQpyc/vufiRPYEOWboHoWQRGLwaTKgXOW8nqygPDVKYEldMHKzY8vgqg5dOkfFepRQJ5SxJGP7NC
Mfr5PWqqc4uIdkddF9DYSGo0VUTzsadfkYzQ/WtzwjMP5VYrPNhEnjF/2r75FgWJI+ebr/kzandw
7T1b5UXcKtuvoQ9ZLWNCv5hsgd0EH8gvbtzxn9pIG+52YQ4+UoJLRyd9LOsB3GYPLTE+/LTWD/5T
SVA/MC62u9bMgKQAEFAB1GEBzvws14yaXMYlhSgAwDatwGodlN+q24EaZxClgN6/IaJXVqFM1nEH
TQWB/aGnLVebLdK1Z/kYHie8tWmieSlpvbRkl/jLlqr0NJAS2eDaTS6sQ1X0Q1zXYdiEc1Znm5rI
vKV6M4C3fLorCzDmmWMCsVIL8KOsKMt+TO1x3WP0wX2/fBz8gAh9Xwzj9AoIDYVLozYU6aJ6tA4d
u3B5TSYFKHzGYTHEecuBNHxRmxGK+J03Df91zZ6//AY1eux4mh2J+tn9YvJCovFtbm8g8x3aILU7
aL+DSgJseUmKxzOxjqLMGRhulo4/apRXl062L2VxHDcF6ox8X/JHdbYwjnAPJakU85ssPhbNr9ZD
qBn1KbQWYsmU/UJgAcVQK1EosU2NMO0SjOTpYIRwRkUI+vzbc+IBx21Xw2Ihyki+e4aoe9yWOib9
T9RDsuIOgoreqRALaL4hmLZyyzIvCFjFi5HgS3IacAVt04ywEh0ILU/6NKacC8NPj8Vib5cKsGr2
BKVuw+C4BeQSlZBH0bqw/GUbnw2RtS+QI1d8BAFXuXEg2jXGMrr5bojjkeLdep0NO3qRloH3zzNe
xtUVFg4IF9t3ZsdYMCNImhglTYVm6EOf1yoxqcr8XZjiE6FJ6xB0NEXsl598RD0cxrmuNp7+8LEV
qz66rhCklkVG/YDdSFJ/eE+tBv8mbWmONmMzI1c4K+z+iJQ6QuUFqGiz8RjW0tT4MsWO4LIfSK9A
+fA0U4nNP+/6l24FUQXETC6n6BS4CRpTpC/ip/hD3yWrvAMZh6qm3cemM0GXrxnU/AgYOH0dBBYG
5VYd/wUCSmNdLtmsLntNWgjBmX9fMaLz9kRM8vN1iTSV1xpZjr5aTDy/AjtSi7xZoaukszFdX72m
0nsdY3NXDORJjo1k2xGqI2Kg3UfrkGBmlN5sM4TJ/1YbvOLbYAbTgdnYREjCHdOj4RRxo3H5ZJ++
m9zz/UFR0dRu/0yemMKKfE/SITxoa8VgXTYyFNsUzDGcNDhAIyoLgEIhlEEQqw72HvkJVglrn9/D
tpM++76OTsgcTNal9NQfY6K0xjiWuCoCNDpK9sJ+wFj8s7JSFdDCUwW3DhjXcvSGbUi/nBRvBuFk
LenfMZTWg1Jl98W0cKkN8bUZg516tv2G0ZUpErZmeGFwHae2wdDZxCJeOANaQJwTjdsTvlMdyOix
Z3c8RVz5hN4LL5+NeWdg2bQ+/jEcL9RyEWbrKKQaKYHCwx1Y/mWHEURcsO6j2NEaIPIg7GBakjkJ
knLD6VAP257bo5Igv9oVJJFc7YFJR7cHHnItwOf3HFNZRjH0CkoZGqj9GiiOe5EbVsNHQNQivnqC
j1mCsoiFp87ENaXNA9J/CnQvinjFzYW4DKdqVpCTAx3SoCPz04IV72azsQKh4hMlWQqxR6IZ0KFV
URWQ9zJLkiAP7CtXD0hVc75Yezkjh1lnmWq9NpJBJ+X8P36WjTPjux9P7H+tqDvg/kWgrs8SgPFC
jX9P2xOFO9m4VK/BmaCdFFP7aHMmQNjDsiRFCBH4VZD5cr6A3iJ45fDXmL7uaOjsGhixu2BxpTib
N6rn0UNeq5gMHeGH0MkAF+3VLB5bLYwjKShnYXR+bVAd+3HnuUxOZCXNJStt0Nu+LvL/d8VmX/Nu
Ew1VuKclpqx7JiUHrSXmYP3U6Qs5+WqJJspLpIAurjALqNuHFUE9NOPVoY/6gAqO1ICJWi/lOPRz
80k2NytuVdIYqNImNRJ5D9VAAjGbPbcSscNMnBbYwHhECW6br3SyxDv4v4JI3Md+tWoOmX0HFnL4
jqqY/UflFh0aGK/jOwBjLsexDwlGNl9lLdYaVn4A+j+3Gv8EVqugDYh+OuIhPXTsixo/Ds2IxRnI
OfkwZdGttBxg8oPn9cb1V+cu3ikpuJNA9sqlyybV1wih5wtM2lykG9GUA1AOtKlWmvzrD8+1BeyA
LyjUncVpmQI3ELq5j5sqgcl/FIaGTHDeK3Q9MusOnjTaLvuAHVIDkfs4eoHF/FtRmZwR3D8xEvTK
rgZbQIgmPqLn2uHX9RoEseU0ho0M5b7r5620jf/fVncZyzZzneSED/MqDkJA0pyIQmH6y+mvn42e
BtXv/SzZZPMFZHEeggFedjCJOxtAVkuUQRZD4pHgDrU2S8DbqKbCMTgKmBncIh9a1+CZioPCfh3X
wP1RvwkRARfaz7Kqwdzizz0QE3R3atPTB/KN+gkqPKTgIvIA4x7Z5uUbdOTSBFd0m6aLH6r1Yoqj
ow3823kka5WPB7x5PoJQJOyKFeJo4mjnLlzMPZw/h1+2GYt/aRL2NLpsYQ7c7FEETcyPSBM1iY8Z
465c22z+Xv6gLsKBacvaysXDJ1m6REqmsUUuv3bstmCtuYL55DSw/jl8geJjn7AH8NgrYgFjKFMc
ht31lon8GlWk6aRsbJA5X4gjawzI5saT3q0IIe6hZMm8+Q/MKfNT2TpIAHhc6DxLW6acIkDPG1ty
odTNtiIuejrJ1RaNqy7vAIbxEi1cc1LrYlb/f6HXTpLHvZmiylC3HlamfmRE9Fhx8In3HCZa/A0/
q66eOSOFyZppQzhEp3praooTjxRVuufv6nke5qKdCJI6X64giSrMNMeuI0m6RP6Wht1Yz4os4qRj
E5D3dNMaQStKEsxq5Nkfr6FR6b72H/EGM84Qhc3BdRBx1Orey9+NzIyjU3x8gZ2rZyriVM4H3gdA
GHzr3dpok4QDCk+fe3HKz3Xq7S7m8s3WZFCYcEdc7WEL66gUz1O0RlMJyL0ahXm6lG4zruMgG4Np
7mcZHslBekuhR8SIEe+9pOfSSSW3eSC7zD9BCWBvtNPu14ev37DH6RpNerOJZeepAj7c2HMY/HVC
2rsU9ObrFlZVO2XJLbvrwr9dwpHZWVBcauIG9Zi44KZv6EzSoFFLTFfj/YLxbKJSRJyTBn7z1ayV
zSthSeHV6ipd7VEyAniEr1TZaAxD9sz0alWcrBFVP9hsqVNba48ysuBCWtb3rv4YEIaJHAkG0z8T
J3hnZHYhjyJFaQz9QdLavppK2Hif5CV3/QUOQ+voqvTv1647J8QKBvJHmDaLFRX7nu1fURAT4CZa
KYZgctEA6zN8nJqUpv/riHIO8H5y3W3MiEWe8c2QGYyj3bJXkBvT+qO7BQGN0F9lhhAwGPd0obbY
wK2LIHNjmwaZfjUZPqUSwoIxOUxcsIxOLhzVOC3T2BeHkPnzvEP6oOBymRedAXpbwAsJ0vs1sdAR
I92Ds3vtIFus74JIn/wcr2Yx5c7NK2iKOvj+yPSkzRW6TiivtTdvHv7MqhwgFO0A5AgEZCnLHwAD
UCmgz90VsX0d/XtKxdzLoXinb9eu+mAZ/UzXiPskHQJTE8L4WnwhNTMqj4Z5zkeWu59bW6HxCXGN
5dbMmY+yeYos7ewaUf/BVjwszj/bM5TiOS2o4e+UqLWaoNSSJKqvLCg65UIuD9BdNZ9v41GCH6bC
cSUCeFw1kV6XXcOu2WlKQK61GLyA4CTjsx7k/t8TXKcK7iM4ZDGrdtaIhHPQ9r4jNdnMB+rSAVg0
Azn4Z/KYwoTN8zNrklNUc0dBPnTPiTifxHj8U/uZyExL5odbvKqIzwJrA/3xll1U+6sZwf7a+5uX
w4h4sUcItoW9aFkOS8pNad2mpzbDEWz8FGQSM1kQJCaE08yXABaW+1fYHbmHYUYuQbBLU8DwHYiu
xd+jnBDxCjenYBH8VAPS6LsI2UB2nh4PD4kgGIvYvwOVzO4X411OisVvC1f0NsHE4oPn2dkbLTgG
ILNtvZhwjXAvd0EQW/ULwMsFip5c2PA+b05i1zpO7o1UGUKoDZgAO0FVcRVK6c/dw9ZK5gijHGWk
XQCEjWaP09VZIAuItFaK7K/uR/g0oSddjV4CMfozFJtnSIVPamWP0f6VwFq02z3LzYmjV1qgD7o2
Jx0p+TC5art2gU3zVB3/LG1KZ1soX6+e0C0AeiMcVTDWQINAGog4ldfUOJncf43cMRfjfBq/hB3E
w7bZ5XL9fY8fk0deKbmArD2L//NoZcujtC/1cBoXegKbutYRvHeFMjJBGa+AxoUWiD05oPZWyXLw
JRIAW+w7S1ChA7quUHWlCKJw++VBFFjm5VIj6yQxx9wSGoBd8b+MCz9rrdvUHGyDyzVLFJpgHIWb
hM95KYPoD4MvkBK2FgfqhjLiHWpVSe4dUytbGo4/xGomFL7n2Kdkx84JTvuV8hqH3Ji8uxxLHcA8
+LlToUttdZgXFTMd6adE+J5FDJvJTnLGZRCop223dVRtYYG8wMfgbM3PzOQQp6RfA5/7tFjw1ACR
fOCD6zZxVFKgQV5TL6NYII5mQQSC3EPOB2obxkVna0jsMy5GU7L1i72gJnT+UTOI+8QXb4CXGSSV
kghanXnFaxVa7Wd1YoAhdcsOc1WgnfDkEMEYjgpDF4pYkcV/PQE9qMEjh+Lxie0KWvX8gBNXvRDD
9aSu2W4L7ABu4o3n0WsW1Btr9nKAPL0oJRDu7z5ruV/kS63hxseiCa7moqm0g+cegalQdJB0ZRBQ
8XA2ltveXzHeDxMZiHOO97HjgQPtAHAN7WzVXwQA3iLtRM3Rq/ZiCMdA1vHJOoZeXCEhhSeYMXsV
Kf0XilVci1RQpN+1LntxQjvP8Akl3nWJWl0LZ/AWAUF0v5fhU4JbtJ7lCRWtWqukCMFwQU0D2IBa
PhHP3DDnVGNHEh/N72nQXCWavpwBJQFulG51sl1jfDi8vMm2BZPsIUVYETJAbJ/gT6D754eyykeT
RmFaKOL6nu+vxM8Nn0XBT+OExgQHYMluU6bXj1bdfFaWynRenp+xfx9YX2gHKAPJeF75cF5t0Ra2
vJbbLKiIFZg4M1qnPvtBTEhZOgB3WFlfBSpU/r1rFVY9SYCgoK/ZvnUjFnBS0o3WEBHhmVjrv/+1
aJY0z9I73JLvqEvrut1HFoE1WvUN6H0MKwrmSStTW4Ls7GDCoQC7VVp+gYw2bhs9XGb3GN0Q5g4j
4Rx0W9oQwON/YmAa8IDO/+Lqe4cSHnAKcoBR6NsFNbZG+OU23rDQ3Qvk7tiY7rXLbSObu4bKMadd
xCC7FQ35aQuplr8Y31Lo47yC3j9PzVlStjJe4rIa2KtNCosQ11EHXRuv71XRH9/yJl4LFzOxTCbR
rJ+8Fhc+R2Ix7cIvZo2gLBz5GmjnOQ7bWuwXFYhPk2y6dd7UGfN7VEUzvj8iHQvgDFSAmH8KWLfy
VJ2Q0G08O1c/2zzLfcxPISF0AflGZljrQAcGkJk7MSt1TZ9xYnYUN6bIFWQryJWqKPmV0omXcDXL
CHTbNRVhB9h4zMVRTF095b+OGFpNJyHSmuWnJjfjzYpJgEEx7Zcow5Hq90OXXjJIMzRY6e10NrrT
C6Q9fSfOKdCh0zIpLjYOOxfw5eOuzLTMvd9alLinaLsUrKt2VOVH/cJeXxT/TRNwP+3ZVQnfw3qu
r4lxn21jYrCVfcaWFQn5JGeSbFTncXXHqB1WoLR8vNnH2BIRXrl2FvEkMGRK15FzVN7mQqWwlaYp
SkQBW9IrQ/zYerstpxXixIMYp0w3C61N/voasBugBosxLGUFeE8vtf7qdaGL6YVYcOf2OZYUpyoG
LjMza7C/9lD9esgpdBQYtUqCpjvpy0b8/HTBs+VjX8zD8FZfwcECfeKet9Y61EGdWmstfNG0ECuY
rYBvRisZ/JuT+Lcd0WX2yC05zWfAQfeebs1wrl9aNR7DM2BG4MibYmxUUCQ95pBWX1eAUAvXwVsi
bytqfv+j+8NMxSWtm/3rtgqoIGoRUcVbZGvLqicVwKHfDOLKxMkEqa+VOWcT7/fV9LLVVG15eyyU
ipow7a0eeGRBPehZTurMzM8uPS+yPN5in33oA5i8Xd1xv6R4+lWNaFQto8InPiBSftxyJ9Cs7YSg
WzTQKrxIbr0Y5zD232/9L4Y78PSi+9VDew39f5b9D2o1g4EdWAFQOofigb+xfKF+1li02MgsDHdI
g+4BertsMFcoyhC1k4KuYLLPw9rQe/3q5Iv707mOAnySSnqTVEUqtzJGZabFhf6b/Z4BYiJ9MBct
srzug56zuaCDGSP6g6dTVEs2Xt28REWZhVSboJQhjNE/lYDhzVAgvH00qaHzGrc32mEdlvnQzoc3
jFJ0w8HbMOqj+NsRZ6HDCwEOXUt/mwsAIfCs6RfiV6hGunfSDUqS4Nhc9oPGt6QFNHEklVT6Jaov
cuErUSgmJ57y+UvPtjqEQsPuiwZI9t10J1qVnlXfwDSTc8e+5/flzxWHV4eZHnSIPwJmPdKV6r4F
4u8EPT1GxpxVbo6igrtzSK2DKlqPRzGGtNMml0vo1jnI91M1C+JyxDDjqw6FwjeHAfczqrY+zB0W
g7Jp3aUDbUwllnhIbt/wkzDJj6ZSEXb+l46+4NcrL9TxMPxaIc2zPrSBctAQyuXAqUCDYGnlsQr+
JS3l0UrwD1knHrGSScanqbW/2+W0sdvTT8nKlorhp2k/bH0fjX76yi2atct10zBLlAkTlRH5bFdC
Kel/MsgrfAiX2J6irKls+7odV7wQ735Q5nOe5kuBPNpbimoOuBwCKikKKGNOvd/Pn7X6l30Zpe4u
A8wCo7NaIwW81/lhxLcz45WrxPm1VNeloGelI5T5O3K/RHePlyqJ82Ge+eneso8QgL2EvOeM0wvg
06zJ0HkGD5JmpfuIrpN3Itx1wjwjNleNDSFtHarLVZqQLfCYnm9hVSbAUsp/SNZXq0RZJJDln1Ym
TL0CkYIUEC0ydL/64rmcQa/NiJWbsdyillXJqOa8h+ywWBdRfyd4ZDcKudASMFX/Kn32tcedSWjt
z1VpeBCg36HAA5SsplNPXTn6507NgeaZH1PGwurvJ1OmkFPsex50G0IPU760HmGqgpXQjpZfunlt
yUJFtKuMYZAat9O6it9+gcJ82IXjO3JL9ujOjMXHdjaK/aE7Ct5WwGB6i/Nf2ystk77kfrjIb2ij
JtflEiIOXjMS/m34hjbrfW47V559000bOnI5haXD7sRyoaIok96VqT4ddPcfXkpON6nhZ3E/o81E
45UHU0ZezksB9XcfDO5cuvk/+Z4RoBkq4NGg7SybmwoLEOtQxX8OyFPnR0Ym6Dd5iyJNVfHPgmUl
FRMnS5nwUa5Cbvx6eqUdSPGn87BR9dr2xe3PF8+RUloZp2uere77Ivx6ZqobRVmbMoc95diiktgh
5dxKxSIGLXoAWBLIagsmFxC+Tk4UdkKKaa29rM5C2lBGy33Q40PoVyfdzn33kLqaXoHF2986ldVa
zMHqTY4kqq6Voif+lTfB/bKJuUMmKdb9TkIYHmPo0TEsv4VTN1ArMKr1Q8ue1LL/GNbIS+lmr31g
M8qAGmJPTrtV40f+GyYnqViFHifbDaA561KBS8O0oNb1LmrO9d6cgnthIFREQ8rQKFRcg6dVbV0M
NyC2Fx3lcc8dxxNRa7lNgQJtiPvnlp184zBY+YSUE5ALfZdTWTVRgEKJwcJtJipfaky1Mp7OU79u
LPkWDHABn/b+/yc4n42ovv5xrVfdsmwrNJr9Siwx+jxIerqsrrfDK9GIQWeJ8RXcONln8kz24V3m
vTcNtcQs2usarvOV3FlIenucP/Jco3EJQv6htjtt7hcwLsVu2/IZCri+ZwFlvbAnrESSvpw9ua0S
44+T1VoCEJPBBtgdeU1bKqQwzOc2XPzKWEnNJHAHrwJvM2t6dGNXD43qKON7OXij1tDpb5lGbUrL
NBf1snEpBb76GY8tpx9bU7TzXMVZY/xg39M3gA+cLEh1L/Vw6BhSRHnV/8kuHD3jOAcAKU+D/5/z
3IlemCSD2QUPa1Ta8core9/QfWHNV7R9yjFrslhDxowDSLy6wYN8luja4kUhUv9qJqluWm/ybNbv
tiPF41bUoX5f7zv5spuecpp6aey/jMak0vdsOqinPVWfIBfKthy3W2+4yg9lONduWm9p3Dch5S7M
9iPMQnICdbrFei25BpMgTEwfWebSWT8ysx8f64MADqd/LAUzJAWtKm2TNEvGQlnprT+8MXWQbbKL
C1U0oZBatBVRHCOV42m78BcjbmtKlwW4lyIbOzkYFGeLoSDZ1apkYahtjSI6SyeO4bm7zjcBcY92
QddEBEmxIrCP4eBtLd/etYSjR13WdsxanF8uYJBV0rGA9+Fbu3jKbmpTN0l/ukwPPx3iIKH/rDD8
rSunbQam6jOA+ga57G4Oplz06PhdxTDKQlTXzRzzolCzxZiigmpNbWI5OoOcutIxaOn8vQRl4Si4
xTI8+WnCuT1OhNIB+RkAiW6Ayl3F4n0CJZfAJg6jh1sI62tniwq6rEhdz+90CCU50sTb7TDa70mf
We0s5GtOf3UFwSUOgnpJH/MHQ4AoQssSizudavoX78RGcdl/EnR0P4nzasYEznsNv5Ou+iZpXx4+
cp6SkBPqsuXoRZKkvXVMk09xy2nqEVe1/sxA3+Mo6TW6avBIfUl7gquwsHHpZzfyfWPpkIAduoQ6
D/7ebKsNQfaJq5HMGG+qd/BVm9LqKeRmi958wjnPWMy8NtFzZfep5tE1+xxnr/hf2AQliSOmqcn2
tz+96Oc06rFXXLRYNn0XN/2QH/Kv0d1JjKDd92QmO06OC5HLJu4IdUk12Bqpqu68nay11N0hlo2P
JV1ftgMgzPGZnJA7W4x8Yka+6vvGONf6o8Li4kAC7G3lyKs0O2KlwfswPVXD5CyZ8TpOTTAxyj/H
pnKyCt1XNL9XU0bgtcOV3ynYMbyblYUVIrEmkEuv45AINLsb+eDJu+/6lUxL6xodA1I9F1HmLQGh
xNNmmAOtp5FKqdcXaFoBJ14lLEfhbXoOTOqYGbdXxERjGG3LrmNwhYImvzls+ggZJgKyDaQ2bNzo
fGNRGsvtQymE50je2pGfh++3oIXkjq/uHm2CH5kWd/CUXyVktVHCH0XiIwp1vz8TBiWbihPB1sEX
RR2fIuR4DkpRvINCLg69zGM2k1YjtIbAVCPGWitmOkGzMGN7rL1WBZQnoab62gwPnZ6pTigG3Q4u
Hr7IQYA3kdd/dI/JFgrhbkjcX5VW0z7+9NGpxDDEW22BVz2MIvdrdwXUc0xkqq1xizS9fD75VpJS
9VhOATipTaYoXxyF+nd0qoTtfBKCD++MH/zIMLxipPhyHWJTGbztIL+DVtsrzcPC+hQKFDgNy5se
xJ5ZkdC6syVoVd6stepX9AbLTODu0OPTM4m2xL7KfbTpvkilOxCnK40LsA1U14PdbQwVsQaNXkWP
HQSU+rAVDEugrrzk+41gtYIYmfcFaa2ujmJiKI1L8gJtck4I/Zt78MSMRbfyfb7tqHw7m1dsK+HE
GyHM/+iKefPgFIqH965AYSrUhRUtCfYyoiCebAnfUD+zaFo1TuGiRLMhYbyGw/hnlEJ/pMLG3Ec9
pGuIqTogR2hF9YtNUjGba3aIpQ7nDRuYn1Nz9LhAr/Em+qu4tVOpdreyjJHLzcoew9nzeg+BPr2J
fpAdTCn6vOcfa2JNwDNj3J+Wkl3TqDq4XgFTer8Xn1f/0o119EYdE1S2FfgtnEfniFzLdiW3vRnP
lfKhAltVoIs1o00OjSQytkjyM3Pc5zJLo6YoYRg/nwB7E2eaiFRdt7q5ldHp4DXspSJOFLowzlE2
sVLGlh3zCoB5lbV1LdwwYKeuVVQFU8mcuj0WKER52TyBsV+xfVg1Z9JmOqOycFuhSc9e9JD/hOk4
3i/i7PDdQ/3Wx8U7xc8CH2hCqaTvVVOx0bw71KcJ2SK87a2smcDSFWDBd6obCfX1JmoCKkY5fV5i
vS1lYQj8sVYpIZFGbv8o7QUeeLNYIB1oBfthX5Cm5JAarneJa65qlFFPqp7OtCyYhFwdHi2c14zv
eaEBjudXwaYV43R9J1sFq6AfAnQZWJueZTw/tMwOAz3gAngr2z+0AC7uO7FoaIVwu+01xXZQfpGU
Hfnp9HmU6XfFKZTlDJS5kMCdhh+luKWPYmsm8akFuZcQFM/530U0gX8sOBJqi8/MWV77DG7cfobp
sLR8yoIoQKFHiQ/JXmrhWmPd/sSrFnFNJRdPXyH7Jp6KmlmaAtjwM+4pigIw4ycr5leh5KTmnAyU
XTYE1IvblwVhAlQRqdrlBJbU6G3+TSErlNl9k8bdAHtv9lCZaQtxSgNXm4K78iHaaBZxlMu0LiJx
IPzfT1JMXo1ANuBi0oGqnVvfSRaHLLZrB6JUkPMpmil7zxZ1pa0bDPc+dffYYbGyRpeh6XoWr9Xu
PqpWL26p+HwU4S3jJ6w2mya/bPYex3AQQWHPq2i1gWqh1zlGTx7rvlEtpLxWC7mPE03gsZjxTiWa
mQkjchZKA98ARB8fZVUEc3saU1UAuyGTdn+QxJ6igJZefKoHv591cgZLM7+v0SNaSziBCbynXPds
C7ZEgKzQnSq6+FrMevGHb0Iu95djxr7+ExiqNCT7t7tNqweli8WOsyTVWeQz5N3jXxSZHeS3z68p
3HpGYKTpYREhYtaatikolIwdNubCBno53Bq3eMbmP0LkwH2vUaKqA+2k5mGABsFeBhNGJZB3QqNk
I0kUHy9iZLvCPUCOGNNaURrphJPPaMZQ7v4DWISCsQUg5jpvk18M9fLS9M9nWjlngrJ59p4aG1Td
k5CvWoL7b2xMTMMikLhBvjlRmUvWwyCUukv9//mb5nzQO5UfsykQY+A8kBcC21hJN6Eo0Z5jcjxW
5ZZpAnC2BzhymAubjPsEeX1wGPuvcY5dkhG/WyryROnh0xIyubMpmB9mDFypitNc3qFbirtCNeB5
1GGCZy4TsKX/ug2acAJwsv+IKdTHAEi+Z7GLH43AYkhKSZ/P3jKSB6BO+t/tr2veQ7Um48u7IzYA
epdrRiSj1JhxZzbOuMxfjWAkBjIs/ywoOPsjn7BG4bHEc/KsTIeU86R0t0XmHLYu25iuj6W7ISLq
PlstqO+WImEmBaG2Mj16Hlz6CAqf4GPIYG7H12Iv8uj+UvmdoJBc3P0Nz841qPIkC1VhsRqViyVX
+ybUVmPoGXiRjA96n38slP2Wj8dhJPyMtuHK2ngfpp7AzJnoOC5GRXCt3uTrbMtBfONaIFfjiHzL
9Tzmlz/FmNLRcbdOQR8Y6rcDLnNQdbBlu/+Pzgovf9XgiQNEy+p/W37n3DHd+V/rTWFMzSkF1A6k
OOFCjJEQFYLw5x6ryeyVqXN9zSWD9IxCsDtCj7SpZKIFCP1Hymn33o3U7F05nY+h6jjeB+StaIyk
50E+NkjuZwyPkXRFCYDF2a6Ovc9Lo4BtUmgW1GG+myYylXG5MeS3OJDKeMa7zWlKGDcurtfjhRgA
6FLx7bueGrSR5KdVlKVj5v3H7RQpOF+OddmNX8u/REbO3IPKXP8A1lTWxbPX++sRdGTXv9cGIl7Z
SIs/Tst3L6/5bCc0wc7QW3VSsrXvzyPHFpbVsSWkfujA5Nw9Ioz74Qhb6SHof2Rtm8ecNIcRHTh7
MMdt/WEi2igYe5WER3Al3UMH1iDG9omor7oqTut1LFAYFbrPX7iBtKEHzrt4CjjB7kbDGYvALiqF
rJ68IeNbIdIfqpIFEOAVMGcYz2uGYDYZspbrZd/UTPDyfZTApzxeRyAmSgEui9aLX4A8/tgF6dFY
2uNwGvLzSdKnToL30a+TrdvRgd6Qr4qZ1SgdF/EhutSOvLGZcfnN0TtElpIlKucJBoef5ApEKXbU
Cd/PrMGxS4tr9PQlkZ6HfpxrojCaXtLN/ZXVzlpjRVZR/R4oEuxU2+I3adrvFV1K/JYmq3tezvBM
l9sZpe/Ovx1MbxMm6DQY8jxAJ43lZa8WiEFKhDKyOHqjIH+ULB32APSzLmYu7TBMhysno+rh0nHM
PyFxwcCplMSjq9C05qgUNig8fzK+NOFUQhc1ARD3zr4dBqW7cpBCmOFxgh9NLiODhinrAGXBGmPO
/941ySvJYU2mXbzQajwQSBqlFlL3X6G3PQ7ZaBYP3WGHh3oF6vqYXlyj55ySOuDO+rJD5U5QoDMW
UBttA4MfxH4fDNGxkjSl834mriACXafMvSAAQwLpzbyOD0mErwYk6NqR/BDWXJK8Lt/icZSvI7Ge
09wnR6VEcFIaU3JLMSoPPsRIXCfl2BD+YF9hordYpxgopfpgK9xNSC9J4Dl0Cx3gz68CdZQwb8p4
JCutgh4qQkywtpl66OLCzOzJUjtn0361mILC9xM0Yl/xczlN3WE4nC2QO/gqWGlbvwzF1hyVqWli
KDmUYvwDOophVcuQO0fEfAt/139zzqzV6spyRVRC7X5tCoHwIj33oDWmhx6VuOdB5tBB8lsijhQb
q3RBHX/yvhPgYOpzZw/cn9HQUqEwWBnDNWZafYtwzkJ7cC0Tj5554MyPG+t/Goe8TEAsgsnL9+oh
CPUbcQwKLIQKczkAHVmrDEB1FwcnK7kZRmdAcmY8cfPg45dx+CEi2FlTp3dwKw/8M4srzqMNvlmi
uPegvtVzXCbZDuZner+eWuaWgbF5UJQlGB8VXj+byhT1DEaNcgf2kS8F5dveoBONfMBD8MKtuKT4
lApGEfcZbOgBFOYWRTGIX44PntM5s/Apd+byIkPd+2Y4+feTcU96JfMA5yt+ut7dgHLDyHUs0QDI
MbN6wWzhOnLq8NEb/HDneVTQz3mrefvEuhzgs3AN/33vdkWc2oRwdEiyn3A5Wdl9InDRdR3p9Bx1
blolQ4C8lgMg9mSzPCUhBp3Nf8vDDfgTp5Uk8wp5k3sCxKuwRr1tgbrMdF59Zcx08e4wKQLXQ4KA
nBh4yMt7fh71+MaMdJb2nHgFrSA70p/EjGOu43g13vzAyP7GAcEafaJd0vemOeblBEHdvKXynWqF
B+4hxOnonEIHK0I9p6VjLYuKqWdXJIpFTpSgQW14CwGN4xSz7FyxI2SOYHJFCmr0q4xwUWqaOtqX
AN2mbkmEkv49uGbbD+B8gEZN4Q5ufGMKTGhvd/9IQmEnZBlr0f/DCuzoZhr+9TyAG8ZFmg4JQgCl
imD96FO71xZ8F0dV40XcAYcxyEKcU7tJ+uwlE2OCndxR8jhvOlqBJcT8rM/ZjJk+um7HtIZA0Fm7
Kl3fO4p9Ey91tYqk4zBc78qNmXouD1F5dIP4D0w+1p62tzleA+442gpj92cyhen58Hlm4ycZjhgP
me01/OqRxKRuaV+3RUzOLurFBiYgJ7q8oyYql278gC23CHCmkUCV9wj7Y082wmtCn1tCFJcZBqos
1GILl+UlXlqOczQAB1FLG/9L+9C+27RDU3qk76VRpcb4xnlV6clJBM4Uab5DClEJlINN0aGK8s+0
bpWy19Tm1QjELjMQ1GrKxydvqnZUzTOTMXRGD69JqFVGv1ctfsIlGh+WxNaM4Md5XUsh5dX58lVu
s6Womxs8TW8LO+Rh7KJIrG3wXbs+lPoby4hRfHWYHjQwfvTUxl8REtWHyu4dT5eLEalWBmWmkELj
vojHxCibdXGiJHEsJIvGB0AUHfufmqyMhg8qDwt854iCwfHhYHmrAjHCKBbXE3m9/s2wgW8YF1vl
FNYF80eV/ICVdtGU2ktv1sV7zO9sae0e+KsWKJeBAhzYfK0dFHDLi9nu5yE8B1h48at0AvR/gef2
TVNGSlDr/vbiA0velYD9GNw/X0NqdRsBOk+79qbDWe/jFm9NMuf5nOnQsJ9vmv6nhUtbjD25aYoj
5sV/ymlI3rhpd6QHLovg+36+kMVE/Jvo5hoiSmosuC9WnnF87ycqtkZqlq9iOCBCVKhpvhx7Kj3X
3Wkxrc1yPJtC16Vvvq+CTSEB+MHmjUaRUzcLwWhpbvRQvuHmABSrR1lENNYsIBRIaIOYPoXIUr7s
vw4CujRuW1FCb6YBWuj+8uomYhrwsSQPvSn4lQMvATZHJzlZ2tvFe6rwok0zrH/EAGgGyZ8skyQL
VxVVWteLz5OycvH6CZSqf46TNGspUf7S84/E7jaHyMfGz1fiT5p3tIyZgZmznulI4EhGmgd4iFAv
U8iLRZQPh3nzRHaO3ktrOUckJlb/7ekTtayPamx1TQaxeuXCahGq3ROX9vIfWXieTrdDcFgFIz8w
fuN186Bv5fgJ61qYji56yRiMAMNDThqlXt/qfBW3qA42qd5YwJeVekQe55/nrJ9jxS7ZG0bzjEsH
9MpSOLVc2FwyDRroRadgXXBCA2ay01HlRbG/sHBA2pHHTPoAUHpL4lxHoEpJjA05aak23nODsrQk
whj3L9c4e4MYv4dOx4AYTs8EV3xYEXB1lQmAnV4bcy8fhBr5DF2yWDAh5/HI9Sk+dwKHIhRT3hDt
aOf3203qLs0pkMihlbslA+OZtGcoomOBXzu/yiGNRT8JbBwWM1BgHiFLVDBEVDhHSMxmtDQ+qBLa
MiEuHRzEHLlwsyWrQCw5+mhdkwu2Jtn7ximqxXjCD+GqNZygx+8Tc41FqNJnLMgFz3mYKgUGwALz
IgmNvv564IQOG3C+NWRRvlgM7Ud1krvkmjmd817krs9M94w5S84VAyF9ST23hV6I65NEOCAsh5AG
E4P5VZuHmMZa/+R2I+LzuT0EDCNP4BgcxQsfZ237M3u5SXG6fMV0RGUQBdq8SpC1duae9t7Nujfp
o7Ula+G3yJZV8N+DfnKloCtkVBm2UZYfzppHTVmD0otvUgjAsny9oxixGNu489TDTKT2hP+6CfR3
LaAsO6+dho0u9zvOIYWnu/8m2Wx48tg0cY0XNH2x3/nhf90QkuhPK0LWcczpPa5AjbW3F2e7n4ld
CDc1DX/NQm3LSF3jmDirDJpUwEPvW8+kePfkUevqj7Tl+lF2xNCJxmfEEsIYE0BUTLMa8bLj9tzj
xI8Fc2MQEScNZCrR0uGZ6mMKbfPPCjNnFoibIqlSJX1O8pxuw+mSSLviuuFDvfpxFZLS8BmcXkNj
wUnKI2GujdVnGkQbsV7icTenW6VBsMId/BuTbG0D0ZwbKgrVP5xJnUZxIy4+geReteocIKIQN+71
xGTlHy73jS6QgJUHLr8uz4G+QZBWpBbeqQseCrwqr9mry2dTG1NrT3FhfSFEBzmrm/V5L4HnUqzA
eeEgX48fIPQhCP4yNEix3yUb3K/wK3E8VYllVIy8aYzO9cKjYceNAp+dmxlJ9XLa2UZwhNEXvUfA
KW/jUicXdj0jSZ6TbGq0C3tC0z0BTaDmWB99mYbDglYLH7qfDH5/4jCxcTph+MtTYCD/bVCeZv0R
HqYup4YbYlopHrU0ELhMJWqgFxisgodlHdOo/mjsWgfJGLt5mPswnhnF7n+YPB3sLA+gjWviKa5H
QZEKzkeD045xO0ngx57AbGE57R3Wmassu8aKsEQP43Nn+G2xsGDVJBWTn6sVGu4tWAAd2CrNS8zE
UkfMxLY7ilyX/0GOV+a91v1GsshvRJftF8zuQHX09weUAVmEfy986i7fqZzL96pEPr7qywZIm+eB
D4psIO0eHlj52SzJBPzGErDY//LRvjqS34VnYOgLb6zFEJ19R1JwMCdauv3gXsD/bpcjjIYc5GM5
nt61MjPVlqPyfkqNXK945kDLitYlxWl+TL0yfhovWh/8J53nrXFfponGeeTenoZ3v3CCtfQMOQT3
s7ItRdt7iO6d3alPbh7cyqANbdC7amn/cJ9JdgHJ/pPxDZl8ayhE0ECfQpFN41XYWLS8YZeJYcQa
7XzzpH2ZHJwCylcufHlPNF3UJaQi5jsncIakOK3P+wAWpdrOUYtiTHeQpVrt0IJOJ6EW4Z9UBQR7
BAZDLUHsrYhjR6zLEAGNDAhEPAwSvMpgvyhkUgAER1SMmyqKvCtUGnOQsz/ghsfHoVlyO6aHwQmk
O3vOp7SZrqxZgElfFU2iBWNE+9R+4DXDFQewDOYq24HTwyobWON8hbqkUheImfaRNjW9spiAPu6j
vsDoahnZuAeCDOyKTWWiHc/Ujfyqt42HUXtovK2y8Qmj49U8G9X+IOfz9j0HEQC4SwKq6CGyMKyE
jJg+8svdRmY889p2lQrl/ZFvd5qZaggH1q2RheecWlTcpZlYshylZ64oIOmwNeWb59TuILtBO+Ux
FpjMXHOdiOqZN0ZLNclyMu5HspixOxMwLYrcA4Rc1tBtJOzNsqY5XlLVTQCJjv2+AvbuD4DViXbU
IGh2Qmv53Juj+5KFsH76EtwfZUXepKJUuJp6wmJkPKfv1tLqr5YDB14PwGQl+JGMfRFyJVuR8Cju
0XQa7MJr7xnffv09iurjc+ksjA+AawgnoQ6ly8w2W3GmgFTYXKn7Kov5HVu8vR+fOfnZUiXSHwJO
UCKMvbGMvOIWZQzjvZnPPDIgW+FFv57gnZrwnDtI9wSYZ/TNh5enCE9TdkRPYek39rZEa3SULakj
jumSby2AoxIYW+Jp8izR707WTGSY1yYy4N2MIert95ocJa2QNRIV2ZBk5q8pMHEZ28ZMv8jezIQn
+hrQJyESVnJ3DsmcY48kxyUkSfnd3JL+0c9yDt79CWPVNHyShD93jdWZxZz+wQTAgCTyineHMZd7
x1ewaeUhLMA7gBrl4tpKW1pAzstBhaHL1/HudG7P1CqOv/14QG/BT9NN75y8kqGplfAkWsXyTAdP
Jp32pO/FFB4KWgxzWwp6viKj7Yrz8N0CTAc88VN4zevMYmRogtO7/vewWf68bwKiaQfXPoaCl9XT
N9sTVLMcXGt49ITVEpDCio9kG/fhVfNwts3oh2Znyct6BkmDqR3P2oISZqyy50MJvgSmkwqVykH4
0E8raLI6gnDhWEwWo4yNh1Oh2HqxAR89oshLTLKL6bZFM5XBCyYgZRuIeP24rKqvRLvPgeAFayvo
7FJsbcMwASpYhl/w9iSt8vECldjCYYuebu2mM8EOVCs3XqG0lcaH4L+NacV87ttsJeDh0P2B9N84
35g7/Zuk1+FcdkTkOvh12jvtfYvrywxuMHMRLEKN6P4hgYbw7/SwizJEK0o5vSoEK9CjYumGVZsX
QyxmrHmRyTy5LubMSMRWFFV4KZI3xtmLeUV1TU4Z3JWGy8O8CTWW/NgyEffi0fMEsn3dwgCxf+lX
kuZKMPz2p63AY8dJiWx3MqjGo9PeCgGkr+Bg8IYVJHpV4PCHlaPJ1NlKqPscGVIjgqLGBioL14Ze
KKnb+wtAG3jw0Ao8YIcJpNWFE6ToRrxMHryv52LxitPb6StFMnRSq2bjizR4HuQwIEb5RRscMvUG
bRf1PPqNA0dgzbG9VZ+R92qeyWJERlA76FzpHVbwTkA7rYCJk/iKrgeCzDLcqwS3Vf0bmOx52yU+
eNoQg04OfNqlnKH76Rduy5co5OcBHmnaVRrlPYUX01lmlbpvwsOgD2K3HCMLSFjhsZ0Jjxs2tlag
aNcttKnph3oDNV+Nf6WkQtYhAJrYsvGp6R1VHI4r3kjpLy1emd1/otzA5Z9TtZ8DXIS4nDS64Cr4
4RV1BNjbCwvoefXNqTJnlcRjGtuJfV0d57F9HCouVTmaJYIiGYBufG5Vh4Esl3kBQmjDL46rIcQb
d/NcO6xH711QbvG7UYBR0fxzwAsVAdEon92X125L9DVTR5MuUDwh633kFI1g8GltvXC/weuwo3R9
tYvmPBkoCoJwvG6ITtzBdScNBxhOEqFVTuGE8l+cOtGRlNdYsgGtyBT+uwVKKSD3fHBUZ9PLySA8
0bx+alyPntwXkdFv9x05CXH/8Id3b4i4c2okgQNC27zx2tbp75Z5P0yBKhMEkbUD/5jf2wVsjo+v
K84CUlA874sIfdNjbNPttVNPsrDe/V/4c72HrYGCer/iHnqmko6O3livgx3OAK8bBfCt3OYsi4ym
21RKewhCKUhhWfjWYOeiHGbmuONCEJfqyHjo/E0GB14lsBENGXpVa/u944eo/miLkw5DJZ4Vd29H
n4vPSWtaRdBUcy42PxiwIHVIGeqWQ8qKzSCnYpE6QvNKI9TvbIqQoschXpgukE1vreIzmQ+pQUvN
UZ/Pbrqjsd+ok3vPZskMZMx7C9JBkzVtE+xEa84D/RfTU3jSQ6TmQosezo4AbXPoNkR4iiui5C76
jISwdLGdVj3cHzuRFnAymnBzuFl2sBoXdLvZQGyA8iyQ6wpM0IB24avaJNOH51l1YlPDsdLfOIsb
W/DHpbTf3v1FYzgmP2iKfIzmFpDi3tltDRIZqm1wQsD33XfFcxnscwekUv/LmKu5Q9xTWK6OwlgG
WifKVrhzV+YImluuDVT3O8FvvVbmO77KFClSeDJQ3tmKYTn305I8xe4wAOGjpRUgatw9Xc1CUzSq
F+eu73lzKtt1TsAfx7vugwwHNXQ4cYPNAwgIhEu7269fAqAPix57coEIMNGVC0AuLF19a3ylLcgK
fdR+dJijsSTImupNuYYI64gJnoqRDDJRk30xRvswsOrok4ERIFe8hjB/3vAGaKhDds0alDCBd6wn
SKcsWmS30RGidUglnFp/cWdCwE31XZmXbPT7t0yh9vKtj4wmhYISRCAfBcTvL4hEceDBODPc/GYT
CmJBmbAG8C2Kax9hidV4D4+jE+Bt+mfP6Gw+LEWTdG4f+rvnbsnpZT7PqZ8lEdlWKsXLakwHtYFk
E1zlAGI2Y456zkH3vaNVTBFzUbB57Ar/+IuMawsEhoxatDPDU8YYbbBZLxnYFBDFsBGptVO3EUNL
qKWett+oxMHkVq5QHMMKWq8ADxinDDKIQr+gcDeQLDO8BfM7gmneDg/jhs9ptN/+FzsPjF+jNgnx
budzf9wY/MIhw8AI0plsTqa4QEhLUv+XGCKEnZflH52OGtbYQ+i7dS/rCs+CBlSQ/QK+qfKM8C7M
3LM8ymyNc4YndbnUtY3gQOJMiadOrPopVzgt1b+2ylVQ8EmRpHSi6cOoM6I3Zc6aio91JmF+HNji
Pk2uajjGlnTmz+4z5QBWpsO1yWL3KlEOVnP7bWJjLgk4BqdYHDYcII/101dYvL5ExRclsZRNFS9C
tyarI0nNKmFMYeJYi6TBsOv9bkxe0LWKcmq91UOBgMl41X+Nirx6sArRtd2cigfxs5SOXDfjpPVl
lMW1vfDFlw2TWmuzbDyJv3PxA2qY2vYs6DQwtFlbKB0DuIopJ1EKAfygWfnJK+M3zZopkwM0Vzev
EAmqRYoQ9UkclEjZ4xlLsiIXpt8fQlMil2jWrqL3BxyvKDVF2Ory3LO9f+qTEufBnSrEwhZa0ia2
PmIFWjjxl8wkPrhkZLTHbZQNFTrCjy7XlK9BYSmXFo8av0Db3ezpCs9akE5QgFrqOTjNSlL+rsRG
nOey/HV19Ha5b98jfFsi3PDRx23UEIexzRGwj9LRQNfvF3R1NTRzao2+zqJzlCdCoiFguNVd6Cj2
R960/IenkVU8S6LbqGfNDnP+gyKd/aSSs4kDQ7qUUjSxmLSKLMW8Xgo2TjMKUcQvb9UtIkz0qLA2
bjTGznleef58+ZGJy8C1OAorMQNBYUhXzdHbLIc6rgdpQkR6d8Rd3Tx3FcQxlGR3rgYSqmz0KhQ1
0h1xgRACnvE10A0LEnwQzJWhxYBp175AzhLJxEyy7nCydXbtkcpLPsM6j6TSFfXnnLbh/t3zn+2W
xMWi/qgWXWj7zRB0AaE3v9th2/Gc6lO4HNifjKLkDT6rkHVNDLuS6AYeRq9OLPy8wpBKyVhuzEzP
ONdizD5BQcWliWxBvlBmKeU32vFjJemJlh8lPn/NJV14AAjxx9fLshE2yp7kuKPpKTtQb0EloxX8
Sc5YENC/DraKQepZSpUQdyBF23BABzTTTHGn/iZAOqQmuJYsSAHqnwGA8tp4zSYLaICbZ8276Qgn
0f2XSpQa2+F9+ozGBd8NQQD2KActzGZSJMwr4leXK8YqDJQpfzWpDIaC6qvMMXlhLbGQOk9HezcH
nGTDqKknXldh0ZwY0qiTRSF8sFuYioDrpbdOeNHAI6Pv0hz/wlGiER0ebJSdKFbpFtCg/E/9c8JY
VdHVKk4mWb59tC7LrID8zJsT0NrHFGnzhF5yqQR9qrRxPCI8T64Ky6wNtMjr2Z9Xtkw5GYFzheLD
pxIOtaTqRh0ERr3buWx95n3qBCVyueSr4/0+oaAe8CRJyJ34Wi+xuYVFlBmrO4B1OOmn2yzJyqhb
Xpzk3lzP+uWrU/hHZHhehAexMpaQJ9AHe5+Ojo4KBnVt3fPV+kxTkU/OqCWkv65SJOTHTFwaqt+w
iAyO/60utbUUtjHuIgru8jXG7TIyWbrl0n36hdElcOhJWVx7+zFeC0kld8S3JYJpbPuL7KJx0VE1
tvrqgoir0rI5pJoMLKsyNqLibcEil+6gRxEPBcTabh08Q+uxjzQO9qNrbhoittQteSpr85EuY7cl
Y1o93PUDQZRNvnIlnafiaEuSJ4AfczQfo1cOi1KxUMWpNX70JPCwBTkzoxpy6hNab/w70nuAmID/
DPGWUAHBNJmASrfeB5UsG4quR9WAuuy39P75g4e6o7c3z/+/E9THyyPGQbRc3DDJUEggraRseUtv
9JpNF8zv5RDLt/hiRygT6Ho6EouzZXpNcWTMOfZWV6DBoNgJbnIgaSXdn6TyH64jEfoG7pz0XL2k
4ZLvzJuou0zmiMqxz+ELvultDMl9/OpvSHKoEgpKJWE4e6WF3Wkrd7d8b9jJ+V3Ee0CDQmvHnZQX
Op0xMTXcJRH47sN4lqCBQtgm0F4HMid+1/Dfd4xK/k5Eu4PAipXtUmrEstZqadPYRrFHdsRybvnc
TwqpSeAUzMZF6UYStAp5T/u0mcW6G5LJq83k9/T5By2U/5Tz/k3fRi2IlmPIM/xihNVOKhwbiaB3
9M3VkmhhzDMpWcfr9K2nYlGQ2UXdbWCC59llT39SAuvT9ThuFF5WrjbRP24xPbit5kBPQkw24Da+
thN4SN6IgH03KlB4wxSxdYlSVUgsxxdGRijUvXRe5RoqxvrewmC+ENtRRTt0RM9P0BTiztmKgZ1l
90FWe6rdGTf5XfFq1crcBufSFHuzYsW1tJUENJON2NpOuiu6wlRq8F+lnMZArSgIlj5bYpeumWk1
PejDy6s/ghtL61GbRSI3aq3eHoUCSVz/FrEkzIpVVe3TdkP10s2tlrN4GUckUim9oOuJ2T43XJE+
iU4bptk6iKhh9OVdV3nunvxlsMcMpA0yHRylR0/LxIuPhFpfyx+AbO7cS4f8TKiwFxSCdeSTRSKc
dNwMa0CxA0iD0dSYLgX//c7AANai6JnVBdf4G+e+Wv1n2ZyHF89+j15dlP9ZOpNnF3Zf30UU8XAZ
RpAaoVkUgFCZ+6fTxkejZ74mVOOilWPseEv6nlXedgmHd7/TgvBi7E/sEVU+bzQ+gK9GFmxqwIPQ
Luv08vRhX/vz19fK/AFJCShXzN3YbjYdl1YZ0Z42hKrpapzjflDyOdJdRkrJPxw2r6w/pAU0oOCu
IlTiRUx4rVCVyU85R70h5zaOSlIXgP0gXkQ848wf3H75vcKOvi9yUSzgfrL2IHssPmdCS6REhrNb
jFJLYP1jxcZabu4nG1D02BwIRFWbgb8o3ap0zZ1yo34pEKkkR4ly1rAp1mnE9bpfug9+noD36+1L
4iZN41SdtEnVEfkgbgMOM6lakQ/3gJLQt2og4f159N6VXl2WnXOIQJtx3aBo9z2RvlXWGM/TtG9c
B/OdeL56/CLIbPA/rkzpGK+X7emTZyzigK3/VJOubZ+gWyKst6kzAAZQ3HIx67HDE5KuwWb7h6O3
OY3IT1KzBG+fK4i0KRyDNCkgjMULACghKoimgwx+fLFXfU4L00/qWVZXMQJFtb4S9hoACEZW0vG7
JfnR37FtccnEQIGqKhcOy5qj+Z4+9oYuhKH0IcoDUoSLpw9HbFzRVubg/ifUzTfEzQFIAPyKiURk
NtmWXfgr7YAEjKwqsYST1hAW3/DH/QmwkmXzquL7KwCuEhhvFze4EZX7uXohniedHosVIoYWJz8J
w31Ba9aGc7jmfVkYVPn4sk18EuasUF02SThOXv45M+pU9ZqVEkk7pgbMj7mecE++fzJgyVRLv+L/
BH1/uspXzHXr5+08LmjN1OuYuqpMJBXz1u//edaFTN6OZdTAMsmTNEJ951EU+8tel7UBLfJGN5mw
JtdjI+CRmP7BFy6CWwn33Ol0Vjafa4l8QTHGVORL7UjybS/P2hmGiGcQd4Jn2o0eaC14PU3L5I2x
DMl2XokoaxbQq5FuURobdS2HVLmis52dmojSRmDetcdyIAG/2lLXuIqmjBQx5d0SSknrlW7kDgpv
/6PIOGgmUmUzxMUX59JgwQ+JnxjvSYWJxQG84D5XV6UliqP2BkBnBivwf04BevmUySrfC6jmlvbs
WFm0IZwRUhXdnYWSdDm8lH+vX+2q5kcBS281X2M0cEpWnRzTQypmIdIbqeua1XvFrTZFh8QylJEu
UYzbaWymBEEDbdYXcrI05uZPTbLugJWi0JlKcJ7gc0Wwknju/45+iRnMog7LunwhiUIf6wHhigFf
2ad7ulTUs7M9T05CrcAQ4gw8S/IduwIVjOWcBTMO5hYJdH3nr9CWrh/CTAbvyAiE8n9VPbcSIi08
v/7QgrQbut2iDZHHnVUC0KBoXfjePQghcugQBUyULXl8ZmjTX+Rc501zLSjBIapK94DMoOJmcd82
kLD9QCPyyUyYpc3cxrvVv5GhyyOrsYn9+UoiBMi0GjeV0f4aAxgAWNkgZsGwdOQtuXLe/em0Nk1V
0cXO3hR+zlsjqksJZKBLjWd7QFeA+L14zawamMkuwTObmI3mARt9RbVThZMkuuEzuYCwtPWJSbWb
DoayjjtIK377/7D6OpYHl3FLpJ7z5azqSiGataTFel+ektqXTDtNKsX4XeNpvvVPEAtVadTEPDxY
BXIEGfWhkE4VoCI7zXWA4LRxyovQPfIX8mHgivy+TNDD4gAa7MhKTobuGxfPjkMAhRGwUgG6ZtFN
u+C9ACltcJG/1o8CGm75ofX7ibAVnK9HxFM8jEGkZ1AozCMby4ZJoggzFFaO/PmXtpBIcOZnyzf6
XWcolRbP129eX3sfDSI1QVz3Gfrs5YkRYlTYMDnf+Xt4n1WDuiGyFT9eRVi0siMY7+1DkRxxHPq5
Tc0kMPk7/a4krWe/xl5bVD2hc1uAtpTSP69LtyLK6wsfPc51Rs44OJt8VT+8t1M/SSCGawnklIBr
4y7W1IIr1UHGc+Ck7dCd9xvvv3MJXdrmdzKyUCU18Rc846b7ep1s2zLEdRk7RFcPOfGRkTWdsthl
4xmChcxrAUIYWugRPZJUKWojiOW0u3Gb+MZw3EVowDKr9AIWNF16ihgAj8k8ZQ/oBmC1oG91arRu
dY2Py5tYzO+JcB8pBZ9QvtWFP+Dhd6yKuoQi5aOPZcbHGYYsGGVU5g9It2QMjk+Ilmk8SF7eaoZV
/yNGhW/frR8cIGt7eSMREmCpnghiy6jz/g4z93/ZyahihoasMVQveILutrQmJ4VwLSsq+gnplX8k
A1w2C6J/+11QT85o9ITBsjtk9GQK6fJlWAGMALi01hkOzuV1Dc9mElYfjYpwZrYXkItEihyEcd2m
1jKzE7QR2fwbR8AZqGmR50N6XTSj0JdCWtBa/A0tkcRoe/dcMR+LiVj28A7EtYNaxuzPlQMWVtuO
VPWfvjaw+siDjRDCg7K1FKl9y6EdhjLorYvmbMyCltVtHUKYtF4Ruafn9BpzqfFx7Xv0yrj3LwXY
Qlkw5xlMqS+1A7mEMIc5xQtitDNIwEDqq553g553i5ToHXQ7/1y8QlcezuRqMqAnDDoAh3/bQbln
s4V95HGmy5Qm0M5Qb8EZFqaSQrj3b9WAmKwnK8fpa/Q6hNl1b9Phj8SVsE3skMSavxuoKCay0YUx
Y6AvIIPI2Iz1XFU0Hcyzw7epjYDxpDq0rx9thv47YB9ecifmYOoNRveDAPvE8Qv6tPrNPQ545m4c
ItG+p57OuX0BfisZlzf86zS2FmY3lD5H1Sznt4yvLD/OKoTrTL82METk/j1nVI8+/aWqcfM82Dk7
f2LIkJzEpRHcC5213tCrDuwa1DECjlwdPbORxJCCCDTlV1MgLRFxGPrfohKHawfHcydXbqzjgDEu
CTapwdDDGicl02/ACwwsQBAsYeihPUxMmRbOYobmPbkfzQ5mKJ/a3+e/ELpPcbe5MuTS44cORg7E
zXwkDS/oNPONMVuqN33Iz5zmIjAsj07Byuals0eA6IiG5eqK6fE/HdjtjWTEYTr0/k4u6uK/NU61
FKYzNkEkRLS9P8V3Bugn31qBaXTzhWnzesRzOlHo3APnsGbfZv5+YDisPBk1lshfctrbVN6nxKtL
IfhFGiiz8dZdR7CdsnD07xmxf8Ivsi+ptcZZLA8jgqRv+yqR2LYWMfhNvUL6/9AHm4Z44xllOi6B
llyzWsU++cut0z3nZde7i/csFZ9HGPA8j1GIq0S4N3S8l7ZnZUpiS9BXRSMzxJ4NalDmxlqa9SnB
X7+9ZDgAN4SatA/JMErYsRzAQ+eYB4eXAE44iubQkUI6Q+apkLPxRTEzY5PSsyH61UsU/y5RsWC8
Mfzo5TTd/qraajJjozra6bq85Mmd+Q0Rxtvr3yIsiagGYYU8SSJ+clSqrXAf9NkmD1HPo8s5u+s7
/E/u7Ly6SCij3eKn63N2hixmn+NhMax1hzsmwh6CyJduZqFJT+qq4GmZoz5lvvcTKiTh8/Psdaei
gmgKbIjjJLgvVxuUkQIImvgYg1hV8BkAZIH4eYO0f75PnAqDbZxJ0BJPcBHZb31vEpopg6uZAnT9
9T+LWhErS7U0P4u41DytI/PusDDdPE4jgDaQnFcWfo1N/FiAoPLu0TnlC1GKXF1gqYXSm9MOQeyZ
0teBDLpD+rbIDIJ3BsRAzBbjgEenBjJ9S3L8XnkaGsflWfgKRcv7ZhD56AILJlzte9c475kWluUn
EGmOWUO4RABhvs01gX+bYSKnI/EIbR8lb9r2tq7LOdepPEnaOmVaYOFRyxKuJpzXPiVEZtKwTgGS
5XSTPPYdNTvMUL1j9lGg7OcJbxqViuN8IMpz4XTt5KvwEHcLEKyaP0xVnHHHPEuNEQczbFPZAhuH
Z+We8jPtpDX6qphe9u1N9eCqUVgtrwPF37DP869M28UYq6sANzVigbhlDyWmUhQzCZrRZhHmbe9U
u2OcZiH/GI0vLli8ey6q9k2qs0a94Atk/DPi4wEYm2BivC78UvOkJB1jIzR3vet0KB9Rs/pEYOvC
QJtbf+nChzdtwrtZ3NMFtbLwv8MRBQ+JPt4x/Pcyd4Krle6LwAIzvBMnDAVOtza/BIXBrt83l+H2
BPOkyj0nIsvpUP3ud3H7pM40ddqlkDfwx8nI4cR2EbF2pxuU3CTeNdAwZsUTStOVZ7o95eiKUFOV
y+ATI95cFnvfRLV1q75z9jwX044RAfMhckumW8jxy5xIoKCrLZeNXk7qdfQR+j7pLzRfetb1CRco
/YcqIsoKwEH2loMZ9ia9ALEOd4eFVYY+m583YtWdtkqZJB4+ugPtvhHr9ky1qmQRh7leeTImHgnV
EaQLoshGb4a0OPazzy1i/o+sp3Auo2zOhrjTMT7cs1PBD6h56y4vTx0FzXmc5PQl/7ahZFyj16xA
RYjAcZlbZEt3CQha5QFL+iMGdPi2OENAd56v95mNNEfvObdevS1W/sgzJDHS+B4I/WiEuEyRlRv1
guowmfE5v/KrOn0mnJB8+wp24rWdn/C6D0MXEEM0leE/Y2Z2KmwB/sVBz3F2tjNpAAToruZJ+1po
vAevUTXA7wUKGRC6nA6iwZZj2BxJgdoxbd/IXaYlJ0fkFfVB8bR05N5jKmmuZ7I8MLWEir3nZXJu
LDm4Do8WUSEs/57UqpuhZMs2R8mUOAXyfpTkLMLRKJOzS4JZShhmHLeyHlaUQUacs5D4HbvULv2+
GOOPzsSQfaCC6RK7K4FjAeubOq9/BCqRwHJTjAfOjSH+5xKuatA1acYWP0ho6LZKrMUl5AJmcbmK
jikYnJG1d7mSA9v+6R2Q6JCI8tXs8Lz4oTDPKnow8BsNgq0aeWs15+SaZe3tUvN51qn1ZlFMbjsY
YXZeyjKdcCCIWxyz4DV89SmU83+GbCXHGhNCFDp/nKXhzH25+wbazq7WetBDhwoU3GEbZOVCykzY
5fDAbyYkTHmVVHTHz62AhtbgxRi+W8KLZTUzvHCsmzVZbH2OsVT47OTRQAriJRAZzgoGPtNRhsRl
5n5rSChlduR/1oDvhkvzT5QFLdHN4VQ8tfeSJnbYQ2Sl4kzshaWOpt86FMZwCaJU0eP1zCJbKZiD
qCtOhQfsvBHkU54nOumA6diQVJKo3VmgtvZbWdW5NUyih6AHouLA+SKDFu4oslXM/En2g85O8J49
GKMYdCfQ80zzorNL91PhGWJSq3ZsCFLwvHxhAW8B9HfOqDOZ2LXZW3a5L7zAdtNfI2Ze/gWlFf+V
hOai87tfkv4GfMkGZuaCdWzP/Z/ezEXRMToJAYylRuyjwlneDKPMk2/dN/m/XVE8vQgK+OoMlmNJ
tbrlcPS5i2Bs0uQBbZevOBhSW8bJjYVg5zFzxitTU8u2IcEgQ8jc4nOrTH3VLLCjf24vZ8NB9eJn
ZyYCyLJMAYFcLiTMue6SGvck3+AQEEVpmovCTZLzFCN3ML3iBwsFi0s2eHPAoPiPx5jF/30DbS6t
9VoJ8vBMFEm7UEwVgzTOwUqfGrYCaUP0OG1S/CTztE7G1SO9I7uiwJ6fEvz/4E+aczgZakoWsMpM
haRfizN/nL8+Ns24s+eENwjTTRrBHoZW5o9gVW1JXJOaSkh7pNXSp3117GYsnUa6p/o0SzMpps1i
IQU62F+o8cpC0x+AvjS1y6SCwGkwaY6mL6iRN9jxFX9XE7Hsau0Ypit8iSNwDVeaQGcVkmQqf2ut
zBhuwy8Nt2osxXnIks+DqnX+5hEcJAwwz3CkmXwzeDW51dYuPiUlyw5OWYI4Vu74Ms8KPqFv5XJ1
zxHoKdVjqVMzQ9WVh2pqfhBMvul9Y+GbOUll8X2ou1Y8UERzf+HVdz6g1PMPoQsKhMHFC7QCwlkG
TE99cJmvLGRBk9qg1PjNoIDr5cPVdZAgTMuFEO6K3bHwZgiqMucZS1mXbDvC+52cHdrxVC5tkRv3
Y6zxMFmwZvqXB5u99+kJdKRxXag/zzVpQPfH6kYo33yjiZcDHtcgW52WVW1wjaSAzYaggJug3f/r
WLtqSe035mvxv7nMtf1zHbXMhvZ3o/vbETo0ywgwRexPPbaxRUdVIokI7edJIAjZP1cctZrA1giS
86Y9LLGESKqx5MviyVhPeqhhF7aivFZm/RM1vO2fFpoJH9ra99Hzd0S4tUgevnm/mnKeaFGCemjz
Rm/FA27PKGMDtF/nQZ81h5dCjRF30J4aEK3kA0ULzSHOLoIF9edXTnkUEE0mPBR0giyqlM3CNL0j
QG0FCW1Y97x5B0zt7LpiXPNKYkl5SPpGy3Lt+WUW2dj/T9u2T1VVWbdsAYFwX2KEZcRAwpQwy2mV
c/OiVOOWIIPthXFxdow9gZ5irRryugVt3fWMU314UjB36X4FyiY+DJWcAbKpz0VMVZ0noEs48QIy
GOCoujCSgQCrjwHSuSsXcXyRYGDHUSUYLA71i702ju5LlblALBVANYYyPd/14U5P6eb8oTJKZbpm
J7E0pghdzzL6Xjb87/FAl3fa48Q1Fop7ft4MKek96OxjzzKREC5PJ7XCh82itZgBsL0mJ4GMKfpf
MED8DYwVGpesUOwP01Wrvno2EYvn091V34SaHUsFLLNdnUGL9S5k1gqzTK96bnKeIRPogGBhrzZK
b4Ekuibo04qyZF3GJ6adab9XgX4ZTP5CBvxGPNio9BZgcFAdqZRD8bE/Q+J6thEC82mq0x/HMqT8
8idaH4wRYjlcthBgP3MdI9kQkX0BmckXHbtlGxS8Z8v+G5S3GeXmVrKhZDRxtha38UwZft9ooDdR
CSB2XmOuQm/DrMdXXqfJfXacoqp/GTyxCWq+2M6kYFHN/Zs4IZOqeb8VLz9jPgpOj8mrmgHWUrnW
QBn4oe3+n+CY5WvcM4rCU4K8eKopZ8arlOdEGpbqVx9V6xzzLnB0vz3WFfYsdrbaqS91FD5LVs3Y
Xgq5qo68rolIs+X4NgmzwphnLnEdELCDtGhcMdC0Nsui3UW6VhKTZjFFRKS//BZAM9Wrx0VrjmTK
507f4LMc88QZo3UtnZmjSxQKvYIQly38h+8pmjlDAT5weEZl7xaZRb4o4as8XSkyOEIcxAEV/i/6
sJfgY5tTxsS8gre95DEoAXsBhSlmHQvJBGoswTKR2TqMUFjY2DJ0eOTNClEu/vl8S7gb3p+Ueesk
4mNAPapvSWT/+5TGcGgFqg680oqF23vc3sGhFnWDFXra6L0/cjW/g1Ai+SPF1kCZfiLG3easSsn4
8iH7D+qZCG0F2bXHLhZ2JQcUVG4htEYHdzo6qDLk+vFU1OGS/LFphv8aPKic7lQC+dF4lmzBkgcI
UXR0S3s91UfcGcmndox10JIf8VYQkqeFAgJHCtW+YlrZ1jOQu9czhLCrVdUCeBZF2/+tXutneTqm
cCM2Uzv1jAxYdongAseDY1sttTjaBYWLWiHYUkMqYSU0Et6apNXPCNFxxsHOcheIQjKesfTBJTQv
t9LkhkiU9MajKP861NDa2oidtK69IiQV27Q0Gh6xO0sXAor7XoBGuBmYY+ftGOuLBbYPS62lEI72
qBKmCnq22aDtOo1oh3EYGnqggQoNNJloiN4uHv9NzmsG1u/QIMJI/cktAu8/64p+sd0SwFpIQd+6
rVUODQfsDDCIyoMYRE1c+LP6cex1UX1oMS+pCABwidym4qeBQu4aqd0XSRIllaFR1Fa164AWSXwH
Z7WAepYJjEfGh1ggPjFp8z2gWvxcbHj0oO8/UXymlnZooAyHPlqhLjkmqrzjT4PF0ZdoozY+TyIM
II2FTdN6F4QP29m8snC4FRIJSOQmPCtZCFRKNGWF7AnmjUeONoane3vzKSmgicgDQ+4a/khSX0Lp
vdJ15xqIyeEpRiSv1r2EYIW0lnKclj7XeTwW099M09WtTpQAW1eiEHwnzQEAkPWUIHxY67RuhW+x
YhI6ySiREHSqLfiX7kCccsicZ6v5eusPifx5Ihqdq1glBYhDkVcCy0Xj0pKc6UrGSnuLvHJije9J
NVE2FXFWy6jRLdesFqFOfv1ZxbnpZPlFbGD+De2mtdKPr1jvsmxoCtsf3qXsEfJh3MPKjP8YCknQ
RTsa82svZ1gP2Goy4w2jzotyFbdSI0E8HWKFt4jlj8BzOjZrC/em+ah8VYTA2VoTPBMX4BA9+VF5
LNPZaZNKsDA/0zRo5SKkYohnDlNM0oseLEeDzAdsYs5JYibCLsKPnjpTie2y+hyMIACZWY1PQseF
D653XpuXfYxxOnnk056iPkcnV/+Ug38FgScFcIdo3vX4VAtBZl/uVOjRAdNwp9CE/cDPw+mXrPWq
02qLD9//80YoOwglIu2Op5idvZsMn3KoIfIjuatEBBZH1fSOo43wVGT3idUSSakiBK54vZ71jqg5
M0V5VPoLqRmdIJFc8jglkcnfMggAVqq9uQTz0WrtDfBhDDYAS3GwGMfZUXwwX6B/atwBrsxGML1C
pjDv2jfCKRtkK762Yo4qMiwbqsf0O+vobiRtHIRcOrGuGJgID4vJH5qGpPlbAmI+DjBOEKikXGVO
WunuWVv7Z0yjtHzf6CdNmVUm3tikX2nWK37AQpkbVntnd7SwGh8RVBMS1uk9JnbyLD/X5jq/jMbh
Il7ZgNlib9joeh7vvFNhIcPBiJZ/vKmnp5SOI3kzdtS5zxybtD9BtZb4dZkHy45VdjdtdomE5jGv
tOsHEMSsqIVViwT84y8CW3jz7N1p0kUPMqxMSAjI4KBZ3UwXvMdlUsProQhfZmAEU+3/PePallYA
so+TZf2vSnMH3mesjvuFu8B99AZGvOPjffTLfE6ThcbTMVRJ1Dg5oZCkMFmMJQkpSrpLDofOceRp
vFPpEw3zYty8prmXsmKV3/XwBWdr/WflBBUgc1Qgp/duR5kJ2jmYz9ottWChNrpb0ILKlfqZ8nA7
7A3tNWE4s7a7aCcUBBOFnWtv4eWZ/Xyag2Nw3S1i+mIqp2zGFRQTSrXtEZy7HfFtagU+5ckDRl/T
7wA83ApjqCNkf8N42cQS1726Oxr3jkxLOaMAcUGz6vx4HjZoytqG4H73ygd+rcJNf5lhYnJrgaA/
gNYMrWilTV+vhLTVKteSaiip6quDFrLNipJ2xnggV8r/sIV7lWbE/nLOtrneUI9Lwd+tqV1QEXa/
hLZAgX2CMMZ/8AU+7Y4aOwlrmIXHQzM6mbWxeAfsR7ouqh8zspDTx+3sHktou7ZrNHBu1s755XPu
A1otuIVyhdDhkynGTviRbceov5V5FEBaKJFSX3qRNv4t0ms7oJ+fwDm4gyc+JqKxi0bmggm4812i
jcvefY0aNcLwJE9UlrvHFeCh25wAbcICcoW86JZ8mEfvUwAIHQr9d7g1orF7U4D6nhPVXszuo1QT
BXYq9Td9/lUBE1q1vcF4aQO0nEb2iz5sWFKc1hjEe8hWZkmb8t/3zaUFhQITjc+ByLVTixNlLEGl
rZ7ZpSGnx0Snas+XahOAQYwRfPYfrHY0BbKZYqhl4paPnUcddbxED74j15K5suycXV3l9jasr7p/
ZbLCg8SSmchXH4TMFefX321DR7Tu6lVATPxcjaMY+CFr+e00v7o3RCamhb/tYs4gIvqCLmo21ky4
8WoPgIu5euj/4wBQRxD0+eikQSrE9+4NFDRdDWl2e9VOFnKOZMlH4Erk8+Mgi+C0edRghYPoj8bj
JA3wJG7VgdzaHjlc6lRJbdEQZKhEp7tffhcONxJfQ+Br7Z+4Bwh1D/iWHjE17/Z8JHQq/+f0/KDz
hLmWghiolAkdmEsQr0X58HmI2Y/tKDeOsq+xzK9mFaeeZkKdPir6oCtNI78/hsSc20GdwUvuSz+A
F2j4gwWhJOdWPrISz5LG4eXQPMC21Pwy5uEqndQsh/h9O0ki7nuTRFcOZWvQdc4Hs7HUiWxjEAG+
h0EXZTOcWbuW6EcAWwkGIrNZGFDMFubnUv2NYMgtbuPclDABZ8OjwRrC9Js/FFraxH1yUU8fMw5s
3VBunO9FVKQAfvx0qWc54xWxFRk+xEp3AIsBVTDsME5v2VVb497nd6Urz1ofbiOUZGgivpx5KYuK
Oakq2MMeYx4h5nE6GVwmF9gIutijrpuAP52VYdQQLTYvL6FUHSEc7i1ze6OJvKBgeZ399byvW28D
jCMZQSPMsdBqE++HwLgGafGMlLz7nnkYWGSqHNkfLvgTYSApLf7PTWtbUrHbx6f4qt+EGE0/YbCx
00Q+yUbAlOkrooyfxsD8LDeO+EJBJdZCiOJgHa+WIqAC5ikD77IH1xZy7SASlNraWfy7iHh0mqnA
XRiSm+YIWLg5HBNFkNu4YD+7M0MhuK5KSNEuCuSGcXv4v1mJUD9sp6a+SCZAujQ+Jq8Orej1NjAi
vEC8fnnSEqE55nIzlfw7Vv4YpXNUtn92BZhCGvFZ7txMugKoSHHSudjEavTwBm1K448Ghguzsj96
Id2T+KQSJylhjCtGZ3f5jM3xHhoDrMnINwbcBiRKihMao9AyAIL0SHhenry/xagjX/ACjZ060gcA
WgvIKcNu2vnum1he2yiu7SaFC6MgC5X/W0bDSfusRB3/yLw9/K36hrJVNEMWWrU4Wz0yPoItA9pL
bluEvqxxWAjX1EEJPoUauzqOpKN+TsPK8vYvtzjThvSdNX/XgCqB2XTATn3DuRUYfgNLOzS/qfFe
2ReMGdQDVwXmnAkJ7VIorfCtu/c99ECYY6PiR8agA9PMGgh3j6sO0EEN6lBhgpokLBPRmsdof4q7
VVOcscG4Wovcfebey9ZQtCf9z4RpdV6VieCIy2EPeDX6nufAiXOFs9NFGSF71fMZ8VK7c8QuNd4f
cK7Y/qtjKz+c4Yel2tK5+/h35zMQMWrLmw8XSYd8tQBcpLsu5cGLUhEDofGLEge0MEimkCksS51o
+JJnoMmEOQ1LbEd0556ALvXDVRvCm8JS46W37dZKJI8rhKbMBVsB+tcYaNQSeuyvfhCgo+1i0OY7
SVKZEqH1KeLvnc2k8LlnQ5Ar/xXHQuHP8mOa5u/m8D/ecymYf9hLZk+5Xg/w0Mv3OY/fv6J6EEZv
l8BEEVoqpmifxjOqFOmWITFmvNX9LS0UB/O3N+GxAYxt6p2fSe5UxmHTqO2G40PGFCiaakoDScQT
Bf2gYjW76ns1rmg0sv9vg55RKCgvDUDMuUunO7osHabzhU53/rxM91ztq7y8VYx6l6KpW0Hhs0cd
zkdx2STOxznsd6kZavlBLWXDe+GI0hDrkkXNPBj8R/DeMHYJ/IcNBg7V9PYGXPf9vU8Xv6OPdOyX
we7jnZNHonC2/RTSVNVqXaIE5m3MyoHB2rsWndIyTEJ4IqiXZmhwVQanTvp7YJRvgSPfMvGrPFiy
Ac1GpQ9b0dbjnsAFEOoDoC9UO8hDRX6jdaGsLRjYjD124Ea95qGLO4MCsA+EP9bkQPCxzHJr/E0U
M7oly7QBa/wm5AfJMA2fCgQ605slREQJY52ftcQIb6CV3cAgceAFLa5foRtsA/QOWNoU1MhXoi3i
j6NGeUv4Ofps8eWOrqA1q1uRfjVGryH62b2ufo/9Gcv90J/qTwY1XOdmm/SGSONRw1oVDcn1nSod
Sh6dTAHKEu8qsaYFix0Fewc7fO2fTfP+mEMHCemQcgK8K1TIwlSDW20YsPUPqunaOqDLgu/gbNho
rH260z3q9McPc9i42RIaqahQOkKYb6Sa7MNWgYLUzIwfepvvHmB3hXxRCpEZ9otMCPYnCetNyn/D
F2IoHpXQi9mhwd3KXL5bTeMiygWjLp7n+6ZwmtLVb5bHi8AKPCboKVBsaG9bWiwixk8CsVZWOWmn
ynm2wnssKZ4S9u3oKy7QZFzH9pKV6s07JKRkQmv4cy44/AYIw+j/vOcYAzO2Lrsr6pfS0GXwQCgk
Mgn6GDCzIqbUSSafcy7m2QDR4hOjTFwTRt5qWcYoKgWSHfq4G638i51MhN++okYgs4ZQ1/9l3ad0
feMuNKZAi1yoDAqhjOueZqxl6KNXMVosTi9insIBCEIBLY/3V+8fTV/00F7vy/X43AlOx/RIor45
CDaU4eln3IMGjx3th1hM+dJhkYm1snBtZxy1DMMm9QX/RiMHUVDslnzJ9NyzRJY1xsDixxOLPElV
gmoeHUpo/ySOM+UnI2zX9VlfHISegwjK89cyAjscYkxKFkK89vmYdsJQwCnk/nJQGdDTewmit+4l
bY0oyU9rnz3t1IGI3WbuoBCM6exl0HuIBpwy4WxkZ2T8IhkMFWgzDeHegc16U4FiZaGMywOmztz8
/R5Cr6tdPOCTwapxZuhThtmR4RAb+JCzAtW7Lum31sDdP9bCVDJMzTJHuVGqO0UGc86arrcb+C2E
Z3npl3i6tHYyPJREZxIniMsrc0xpqd5afz7QjepKoYePfEJ+AOl6kB8IHFvffaEatZI5/ZFjxdlO
rIFptbhhNeA+BnptPH7YO1H9+cWkuIYBZI0SDoQP07h8AtRbwyEz5Z7XqtOoy2M67YkB1BJsozjQ
5Ru+/jP+biaIFVWBlQdHDOd7xFpJkJzYvYfOydy3VkixB5uh2VJA34oRBhoK/bbC1bfwoxnvZLzn
2lTzcdUhyRnPYEalpPH3gfclW8wgWMWe6rz1AI6pHSFUBxGra+fLQjU9xCyan8osjPmPBO0fk7+6
KhcV3l00ap9wuS1pAn2gTLDpquNyNrjwbrYpJWugPC7dd9TtCUSmigl42pEj+e5+M9n3Qislfy6K
rQnXTxUDbnA81u2XTCc4PmH+1+iIe8Y/BYcN53918ZkRO6Y+Dj5yQeyhZVxHPADnmoGqe6O/3iaM
CTzNXm0eCqocklM6XzWY+zkPecAG9FPJlNRnS6R7iKYzZQIV51u8ekpGetos7BZaF/rCTabRowd0
VgLY9CW6yNaqEUB/tQXSUjoJoSjHHZksnfDWGCP6FcTXvtoYfakA7ew3isk0UDO91LOMqCjp+wVT
/nN5Yno/kyozDYkiexdSi0TwjDzRgaoBUpDffdz0VUPLrAcsgQGnjRxWcSt08EA9OsD8WZwUVpTx
XzF/ZZdxmHXZhXwScab0rAKvDzkV8e7MB5FtDwOuUQPfzMB/36hGISOy/7Nd0QHvWRrs7nsUUhR1
Xqnm6rmIat69NsBg9kprqwp/AKxJTZsZo5tIQ3gas/B1WMai1Tu68phaVsxrBgjG+7MJIndP0k+w
vfDZW1TwZm7jRriK+dWgedFjJsMzjMXLD0n2QPyoiIAAu81o0M0SkMU5O3doL0W9DKvjLG2c6wZ7
XOKEMiMvjvg9qAvhvJGdcRuHKuOptPSc4d0H+WqiSij/NeMv3OL1mGX0B4d40TZ1qqqbfxVwqTB0
T4BzGCJw0DU9xT/PjLFxCYJkal/Ppfz/jZb3XfLcF5KIpDlsER6F0Lyqr9MgONecgNbb289IAcje
6HOR67FjcidyMNzwNz61la5U1TYeWBsqzp1zyY0+45fSm/iOCae3gq/skT4/8/kTZ7LBsKqdo8Oo
k964/Ox7KKzT7k/4Wf9eF5aTohIf77MEwyxinApZhPFG+VwQtXuuL8nwlhAtwyJaM5EUxLCt2JbK
i26R792lSCOzSlbmK4adbi+Hj2Zc7kFwC+6UAawKrFRUGQkR56V/rwCwR0CFg/cIcMtKXHbCJ52C
sVCCWiEwpDHj9P31t3zAf2L4nKaWFZoBse1ZrRLZ8CS1rBaiQT2b/ZrPVhWyhQHJRNXRYdBlS8OA
HQoFHRJrv7oFaUivhbokxg457VoaiD6lk+pfFcqEKCoo5grZbNVfVuQC4lCsQOxtc/l1Ra53BwQT
7hmMqSdytim5JSFNA6/U0xLFu1f4FZyRVbQsf4FVzA7ArBNgVX41sI91dKMOXqWz6ZvuZ+d4QAEm
R0TfVKEeuEwIpBiQYEkxFVFzkZFvZkVLU8Ld6420hxvVfMyO5Rqyr2nAgxXF5ifW4BSwI0eK4C4r
DZzYJRbIQGKYizn9U0VcqqfI+Th1NRA1U7wONcAKa4Hj+Kdvd9+5HhAAkk1l/XYc6evGsRBsZEaI
DI7mU3fJEy3fSNwKbCaFkq43dUiloDU7TPdwkTLNL0MxNeWRfRFQT2lIc0jt5Ixa/SrE7h8qr3+T
zJc439/PEQF5Jyw0L0OrOchRJIyI/5W3PvLsjYfE6B/r7Gh1MfAdMp5PgPFcix4u3KuqOdjpPHSD
d3SakMjZIBaEnHR18aW4IouTkiSMcCKjYi8u2llXyaL1BXJgvkvb/H0JeCW6hSDFhbJLy9odTmGX
+T6n7KiBxkcsPcIUPxSI7RWRcN81RJ91mT3N3/kWucRjL7kI0Y7swXnfn2xgk70HPcK9uxhhutPd
bytieT5VTyAxN+9B7OgS150WPg8s43ADHmdCQNi9XF3aWuwRMvcYfXwQmWgpb1B4oBtNdugogEDR
9V7C1SZxQ4F8jnBo9lpjQeZ/xFCcGM9yxjzYMiKl1uUbzGAzOJtPtyQ1WsBUESAWoycTHG6MBYy7
Q81ks9GGVRVlY7HCQOnOxcx3H3Bd1MzzmMz3/qDHqPE0xr9wfkClJANF/fBPFGDAyRENuyXrurRu
nygHBltydMPReCeewPspw15/AXKDFqyM7QqWmZCDguh2SQKgGooHm6fYJykiKeUXWhOSCsL2wp9C
F+DykZxBFrA/V9cALH5Y2th+USdG8PZTuUDHYTa9wIMn5etyikcKIkQV0ha/DZDPgbA3xBQWhrBZ
EayZhVOExOgqjjxxHTCG4Xa1NlwD7q9TntN3hxyDUItQqpPdsXVXEM2hM2pv61GX8V9PnHRjIzMc
nEkTzdZOSBkSLIIv7mFycXYlYZ8MWLSK3PiUQWxAs/aJ69YTWWbtrZFZEvRJZpN57/TP3uiU60Cp
Xqt2TOkuEk+Xl6o79MZBPyKkgMYl9DVR3qdFNvlrwpBKcy/b19BYSJgFpICtHfBtHb7maiHglV+g
lnc7tdXQ1K9hvv9R5Ri7LY2jt1JMNvWiK5qV+ez8ELvcrtfIgwNo/EoB/8xcnekucDib+MPoBxja
xyq/d9pyOH9/gAATkJMmNnK5MZ+5bo7gb2bqUzSWRq4cxQrvpez6yDZDlkiPYaJclSBgNDUQ0LXo
JMJnfrpD3Q30q+K/p3Y6AdMiCPGeZN63vOTj4HdigNK0sa61a1Vu/WrFWbC6aOjn8I4X6a2hbYak
cALPN+QJohvG1VCea25YK2GyBJllUZfI9u95jlW5Kdb+iP5n59UJPaIx0Pa+qjbp42hWG/dRqwNf
NZEeIXOH6Ja1yX5aMNVerPGKbWyiVudmP/8Vcsi4PA7OyH66nMS+LWm4y7WNlPPujs/Py7UpkxSs
XY+1xsRKprZTm7mSzYu15HRS5SwHX9DsAwNcvjQloeQ4xEIOYq59ASOAgVoVZHppe5sY013CmNC3
m+C5VnvciF9Hn5ImeNsy2i+yH+8vpSkpehrBmINDdAu07adhaT1flEiUs76gXn5CopJXN5mntuTG
hW3W2/su1xMfvpOhFYGaGyT2FtP3reWvDBC+c4SSOF3mVkV9Lk3Vrqz9g8S7YCghM1J11azAm9J5
D9ASHRaFVaKCe/2ZyELcPpwLIWE8uXtXaIMb4il/WXInpQEggWJEVVDmE2+JdY1D7PBakv7WZ3Yi
STu7sJJCStoH45tFiw8BrIB+ORKhQmR3yNHp/bvq+J6Cy3cf07zd7xyqXL1NsijtreSI3GphtH5D
s/ZONaAHGYInD/jgXXb9rbNN/SP32snNT7IXywKPRzUY4D4e/QUNXHVQyVXmy+rskiF5eAYpQ6nx
nyS3P41IxBycSUxo5hSVIpyg/sHtq0NEuI2Wv+zJy/hNDW/gv5MJQiDL3t/1jllmPq0IkyBCEwvl
qJZwBeuXhyYh3At96AyFX4QkGUGo2PfAe6aQzYLUs/GZjbJwqv/e+zQ0vu9zuGBtGJOppDlEptlo
iBmBvrYvEbSqXAK4bhu6NiZyFakwffrc0Lya8XbskHyHybnBiQYXToKfAQN4d5ioAT9TrLl5xTGt
sqCZU/HWVfKF28FLoMS1jXengtk0ACKrSQqfOShVIKlQNKGg49ZX269vVWIZD3PbJEiLAhhZB41K
Xu4/sfnyB5dgZhsJwE+ZDmj/KNygV8joTLhHvxEQOtL0jPMV0kjygk43xIp4U31ShzR4YuR5Rr8k
hu7YP5Rd8xV8TK+7k+FYfGGBGTK15qoqxRswZj0a1DWmO8km6tH7t4phfYSk4yg7Ui75a2FKFpx4
u49brtYn7uKImYmY02UL1ZoV9thLDPKsrDvAHA2XsugZsDPaqzLxwkNTPVOwUnEFrS4heDNApMLY
/UV4fEboV8xeN+q2Y7anhG5gMAQeM75fj5L4sh8M7UGzKedAxH9OfG5IDPq+34YFtuIzFKPt5CrC
7pqbPTn6dZKVIPj5DYWd7pVmdOS151b8oNf6gWXFSJE/BW9dpthrmC6YOdYUGlgW5xFSGyBuj844
llTwj7XZXZ1IhTK8YYzjBJQs4y2Da+F1k2nbljW+DLel6l+Kq7a8rDiWPBOo7bMkdzDdJek74lLY
BYJEQIFWVM233AOw6XVHoGfog3Z2hYrHJg7F8rvdpRyOlYqloM+uGE8yvou6myL3ZPD85+X3+Rb7
vmMOJvifs+a1WbillunEbzNT1LJpJv/MZvAtg3j38QqmQCXWWNJoc9kaZpACV9tBG4929n1pTULA
Tjbt7EOBmLkP3jfMicweXYEPjlsIVB8Q0NAxh8Awtk9SYY/Zh4+XC5UmHEF9LXliKsZ7pxhjvIPd
ojZsC6qoy34SsF/z2XaVqg6QYG1qy3M+KKMtTngki/QxiY4kBwK5KDvDsGmIusr1Onu5DxW3e873
PRzx0zWeW8pLIaAyYzxxYCYiaqmCIKHb+eDt2obKWGG3zTb20WY7hWT1lWT1T8OCWvZusu6vuJYV
6GAD2FC95THnbsTOAWAqGI7DxWtlEDaWLKYnw0DDC72R3yCQGeNiGMu6GzXvqb6dvXJ2EfqsUCWp
U2ucJUI/O4OpA4KuDjrW7gddzM5hC05+/HkBoqdaPu/iEC4ArQ2AX0w2aHyLANF5r73jZ+4iGrl6
TATEjiaiuPyCN3zIEn/EJlyHIlBkzKtsEpvNuahcCFJpvuU3pu18YfYU7ASz4MgMM8zjRKp7o/Id
1+xXlea7nxK4YqhniCBqcHe+/W6bqJR3UYZwbmj+vYuOOoIOmfbkr9Krmn2eXLellrQfRhGDlGW6
GhGVbr8c88qeZUYF0CInV1qfFVQ/HvnnXY79qrP2XYFKWi2/z6ZmYycQFFmzl32JIYVaUvFNhfBb
KKmPlS2TDLTVcff4o9EVJ8KUhjlzSIo6eDIYM1y2OtACFM8CtJSNx+qTMtMmQGnEvXPevyKx1ypf
UBgVzGbg8leiA9Uz8v1PUQi1V6b3i467yrT84FhfWkjaei1fxO3KCLxrrk90IPOePqCBI35ftN9G
eMuAAhNM7W37hjPDgR7u+TZ2l8JD0XO6Tyy6bQuaid/JV9pz63W7mdrp3h04h/XfGJ5uwRADMYbA
Dwacy5eBra1IKejSIlGKWc0Bb+MKFmTcZckkE3PjRTNdVChan+I25tOK4QmE/xfidd+f0vGNWKmK
LwneMXgcLrLRrBhx1+RRgcoYJ0rhREsdenB4Av3bscDn3FsxLd1rOjkZmEJ2hIKAs7GIC7R+V4rT
qFwuQbBZMN9GZNEDf9GkXHOIbKLAU5LaG6o04XJy2Q6ksPHiHp1ZSn1CMW+1J7AB+erIFPh5d/+j
ZQzcEr8GtiLih+hz3gDhq0tqc88q6B+DIr8c6KhNVBN5a6NtwUEACI5he+JjgrY+pMI9l/Ok2WFo
OFOmR18n9sH56CnbjmhHhzPyKRK/o3jSb8QPXDb2hj9jNbpiTrfRx7mEYSZc9nvlCbvQb/ad80gE
xwrnQb2aD/jxxpcO0Reh5UDOb0/0hWrkY50eXfZ6XKll90l4DdQvz53o2eblZac3r1j3NQAV/Vdw
MrcZuua6akFZ2PPHauSHqV00iZ4zaYnwqSLcFmy76ldh5GUoOkjZ2Jb2xFQ+bwwYMpfD/pT2+pAk
FOcaKmINxEIjv9pxnQlGTFXs/iLfQpm0VEdWxAcm0Axvp7HKWBSqkdci9DtcWMS3jQOg2TNNo7bk
/6GM/6bLuSxXcw0VV8nYI7e7GEXDeqDr/zHOryHxMAH4b/W0oVyYzFEJ4ArMT3NlXMQ1Bgo9xlKW
qFRA1Ec2/tNnseq6mVI+XJNEc4MyGutQsA+7yByFVz+Xjpj1Tfzrmz9pYxB0rsB481d8feRcWnbi
51ST1OrwjNk4HEBBC3F9lUex69KbN9p+xrQOqcX5xn6XUlQwdQZ4LhL2LziZZANUmJmtel6Hvxs/
dcyra5NqazcGq3PlSaSexD21Lb6JzYegD2sZihuhlOGdq/dpr9Ps5rh/9VWnuLwRFGFg34j7WFxG
Vom/smnS5lWKU1J1PqoDUxn/PrEMQG0x5fu0w71OzprGtH593LzYhWO2tRaSUh+Adg0Z9Q0Ejj8+
gKDrTBTmq6pIcb9uvauiXS6wnYaRO7K3K88geXYqcj9hX0fP8W0+0FcI3BwTs5j02RrSJpZpeS/o
OwFawQ6qRDxzVIqOs39i6q2JQ8zGhYz9LrypxwtlUBk2ZQT1UMJbUo+npQgbLuMeAoT8YGoOHeDo
eStXa2H2hcc/0+GJbWGTe9Wbo+jjhXg1h3rtNZExb1Dvl80/6EyFYMVqsRNOWZOUlZ726gbtoxkt
T9hg8QGG86RJBrrxxzYUffTUpgTSmWEHm3OVBaHXIDct6jeAYIIqfJruFLGVFvY7ktSMExX0Wn9+
zpxOix3RyXP/E3OTgg8mGNoyWJ6Llp2+K6bE2taDYSJ4L48IZYa1rwGnewOvryRoslOBGg5MsI2Q
XraRKFKM/Xo88fOmbbYo3uR16eKJNEvMkplQuYbp2MnGtJ85T11cMv6DqL8xpkpJx4oz/A4WBTnu
rlIePh8rb44vC7QEew6r8k37LsTWc4OtXcT6R/tsSZMQkymYBaIQCoifH7zQhkwM+lIrqdgClkZn
GfJHSF9VhY8PXEeIn8KD56dYKVRVXWoL35yOAgUXrfA39iwGnvK3VZasYsWoKE/6NdUAzNQCkO+k
wnVnoMpnHsCzLupZXpRiWJo/V6YWTZvYWFWbghRS3SpLEyiKrK5WX67NAmUi+yQ04LNyURZid+hL
nbXB39NehaLGJ6c5uQ5u1WuJPOWNFWDwLCGhFu1nKWAWMRsytCGzNaxsL/QNL38uHgIY6Ec709LO
9Md2+6nPTMccjgqdk22+QKqTFEWGP+TiWI7OJL0eBfxMAPyqOXBg4ihK49+pzytC8yNHd/c1NjYe
Vk74coQFLbBuRWeEQOzR8ZzFaUq/y1HRYrpudi9TXZWGGHsouvDxEj1iR6+sK9jmlMKMZ1G2h48s
yx7Tc4YBXBnX4eC2M6tjVNhkVhMBoQK3bWmcSWOuYdN1afXmXc35mn9ht9kwDhD/Kiaqgb9K1cmN
AYe8bQdx0fdBNUz3MQIlAJfJEmHzz+/ZAGkSfqT9h+yIAqAmmPCIdWshmtlYG0LOZ8AdrEwDpgD9
n1BPMlERr5I70OthSyxeIUhoe247OGE/sG4eUle6aYD0IxbDhQVPeKuRWAWgxaL76uojOs/pKJge
flzWcpT9fD9tXN4GpO2X7JUjYWG6gusr1wDJzAY/mcLlLlq7u4IALFChsGUxUgbRsMpLJU92O3Vs
53fIf211p/82/9KuFn6TZY/LVWsQfb8QnZ/j2K/RSUl2ElIrFHi3oXdeozgJeFQE29a6bFPLsG7v
J0j4u/KpBt4KYZnWI0OP7ruUT1GQioRz6zVQDEHfR5LeX41pS/Mj/bgnA0qnzrT6gqJbu/uPgzJu
pxpJrZ6KCn8VAcYLRarujVZBENSA7lwi6mQyNC7SGzZV6rYGFDzCGzvJSAM4N3i19uHgkliurhGj
Lp3RdUvMR9/gS7WYLtxVArLbjpvXJYkafJaJ0CvsSRw3CMy+GZsRqKVvQC0U9LQtVGw84ReL4AWk
9JKPMmLuBRumH6We1bOKq/LrQ5Ld+tnxY9vzTgcuL2LqoNqE/j0/2mB+Sj2u4qmUCqnHcBXZ9OxA
MGHx2dzOl/StekJlXqwGUF3eykxsOMkyv2XFDMFFe+xGzZM0de1Q5CCKlcB4BIRJ3uuaYQxKIJM8
HHaJIIBiBgN6FQwMg9DeWxcNKPIrRdM0D7CyXFhPPTAY8UqkrVlnJOm7vGU5xer8T+CUrLZxKKXu
swlom630Posg3JXFQXWRwm+kaM3EhMSupWncmm/HnJDbDFI9t4xYy4GoYWzoqYMh6Sipoyl47IaF
MxaNac+v61quvta56unaeRuImarEwnzKsy0n3IMnW5452OVMkzcwJfy2Fh2DkYv/s74Ge3MuNkta
Pjw1r42R7cO7lADU6ULuW1u9YDWix3H0vPIF9Ne+dmYv9J6kDRx852I+kepYiO35eaTDbu+1yxs0
ut55wNojwRHkbFBjVP1tiulcMU1D/Kyncdyg7D1GA20ThWlu81gY020Syn1r2sSZa/68al5pygMl
SzcfJ9Js8RWOmSnqHDipqsw/qa7AjhiZzOFnXiOP2yLnP8uWog/88bSXEubpOVWQaREnzyiufSmq
L/rFQt6Y5YT4VDVd2edSMtFXILtA2aXnZpRmKfQgZ9wOWdPNgELtclM665itDPNOnYvNqJ4m72OX
pv381pRSZLdo2D4rtLEikOJUBzrtjsXb5/FRZOwTqsedt9slSfVtw89J9PfVVioD1u7+NqAX/9JA
g1sCR259qT+YmobpY0iBJUuRpxxtlsQIkBkxNND3YUHjT0k9DLHnpz4EX8J7J6GzKrSx+PX89fZg
ghvAfiB3nUYUHV6qHV3Dge3talNoelTaGJ8Y1s7RT+3vkozyMQ8vmA4+xc7c4IT2NvDUWWWMz740
zr9TklCMpHK8E3CpsX2IPYh2rNMXT/vmu3NL//SUIsQdCGvOxq8bAysaHn0hh5WFX7hGMsEckTWe
df6Wqmh7qxnMaooS2MVE/tG0X1Bh+UoHDFdvdsRNDLqhY2wGvnmh7Cu8bJWo+1aoj9hi8iOdOYe0
oe9GDQ/TzU/Yy4TFFxcoEvfFY9guM2aUpIKJj9b3yN9j/gN48H9Y01VPoLrjO83RITRuhZKRK8kB
zlafLlULOK60ZoelTwWfAR6P+44gW8TyGFojllQ7xgtOwmh9LYWd7qdYlgqUgR0BRxXcyuIu9IX6
U1K+Kg5B/Ag1m494m7G9Wuk5RK1pyzepqQScq6bPiQ8/HNmdv0OHLPa0zJqYPv+523VHnZT8ZFcU
h0u+mVIorGSAejy0pxH3dUfjsNInOmYU/QpnrahW0a0f9mR6b6qQJzPulVgaqQjBCEdaQvqKfhI+
daFb1GzL7moivLLHjusMJdDb5hG8w9JN+TVX+NYJjyqJo6QSJ83uxMbVBLojznHXBeXBi3DK8zZD
7piZt8Gzw8nC7nwq8CwFhcnpy6Rw1q1ilOLsQX4kDBi1QU16dV8PdI7CxX/MO6dOOiI0j53hAzpH
T8g9SR6iq13YWE/b17YtTHMS9D2spBL8Q1IECaMJ/BgcYlPOSrGc5+mx3IKVuaSqa3uDxvzTJL6X
1ObjmpJz3iRjca0+NkLX8M/DLxr2H+zcn1MtgJSfPa1LZt5vv7xJXRRijXlD3Zx6FbXPU/sKcVRf
5voWxDnuqbaXuCpsEPRshWIN9rnuSjs3JUAo8SHrSxhGh4zaI7l/EBVtp37VLb/KDReW/7p5+W99
6ZZd6Lk9Qj1IJH+xbPHl61Vq5rJs16b6EvFO7360zKqLR7RJ+KS01vwb/ssiPl7qmXJ9VCjXC9/K
eKldGaivwRPwgM0F13RcqIUJQnJ2OAnF9gYRFGElqMgGqNZmVuF9pH+fZIVgPHxXp/buclILyBt+
8b9YrRmEf+VlZl+Oix7CP/+CjeewR5odxM9dkDUJNcmzaQneSp+JNbS7bYd+kx66rCdnDNWRIShu
2/Uo8Qj/7kIHqKLkguneG5UC9/7AzyvX68FpVK7QwR+CxfCgpL2uuwDFGVKtgsrIXQQT3HqonceN
0w6NHh6BcRLWjbxZ9Vbp+ZGz1h48aXvfP/DEqq2llVh5jYo6huLmaER1yVczL4NOhrxgaPbsZYW7
s6BNzr7HirtrG+rNBlBYI5dKfBs6O/iOPgv2/OgjttUlOa+nW1f61wwgRyorugjF91sbaX5ljavG
aTpFXEbdBlfM+SEzBkpoZrVo1YUcUyzM574hGLu1qvH/MwoxINl6PEvk3qVmEefk05bNG7Q+uH/h
gTmy234+Dwt+8gWNPvZ5D+BlhVZ+Lge/sRYi4OSf3oXmwq+GbzonRBP409bu82hlkpTeLXRKQ/Ev
d7pzYMjEdRZcA48q73o0B2PlivAGGveIs6T+cgNfuK1YF54lYzEB6rLIZq95YjEpTjN2C0aS5uNV
EjqSRwOL1hdwXVecQkRoZQ0nseJIry+aQ7vPn2h0Yd1DQGQtsqvdWG900g+XBBSzk0Bcgz55uPzu
S424PfoB11Scgm4AsveGPqfTkkvQBPYUsOEDC+cE0VzEwiDXm/6uAVDGURblEX7ppkVnwFbts9HU
pzd8xrSmpPEaAPuYsQzFtcrC6fQu1YdpatEfqudmaMa8hCT6TUE5tR5X4zCPAlP6ax45bXZZQ9B+
XXOOfmWCJ+02WLYEEP6gEnRuAU3ej5SGAOiVc4zXDY6LwPsq3ekWpgrIKFrRRpoC5FwqvWhgMozH
mxO0Vt5JrQf3SIaaSg+vDGxINaElfgh9lFBPqWeOdaMSQSfaSCqh1MF6nq+M4/cwr1M78WyoirNA
P0r/TaMRVJ4QpcwYejZ22nPEXMJi46bqLj1xsRvx8qgBUiiVO4FKjoRpfOw8/Tc1Xamr0vcDVEy/
cpnf08siyQix4d+tfnn1YBAcGf5I3dTvj0+4Z47Lrn1vkMfog7ayLTf3hAXx03OkqOd6SKfs91QO
BMn3mOm6Iyi1DZ1/qBcehrD2rcxqWI2T/hwxGYCsC+Ncb23bYtBVultUB+cYtk8XrggsOuG8KV63
r+hJypmVg52C2coxrmJeI6bAVnislzzLGo9mT2NFS5HKHDsfDNFhXZnGdfvgp3gtXNH4D0oib5A6
vaLKAQZaaqIqCrerDY6lRNM1YXpWUfB+QsocyRBL2vkPGmhEJPq1qGwagoCVeJNbK75jx5n1vgXY
Xh1AAUk7Jrjl6ak7//mK3PPSLGzRVJXe0dTeYQ4RtoM7cy72S9NIs7gl7O4Pi4MtxKgx+wcp77Se
Y5QuxDZoA7cIf+AHD0JO7ke/s7LuqosJbMW0jBuftBHv6o4mVtOhgIy7YLpMhkoANPLjKmEHZQC4
ZpRbclRkvX/skUQmoAr/Yh6u1Abv6nfmDxksvXdxPyN/P+9LPt4Xku/mayTyIZ0mzUebyLyjrGOb
gDIAPe3yHjIJagWcPwZAOnurj62TAxa7r3ub7O5QYWbRptYB6xRKNZMtesrqCOwAUCe2oTl45BCQ
ejaX2PmyoHmA0Xa3ep1jv51L9h6GA4kifpRUGQexo0FkwSpJCNRLxtwipGX/iJjw5Rh7ltss4rdZ
yfpNB3c76I5SUFN5rENhHcOXi8QhoqgrFovWmTzcQ4Pn+NHVmaN0sRrzztjDALfP9WYdLRU5TLGu
exNg6FyDc1QKhVPeJF7QOSIoneImLFI4jJnuyyaIPU3DOE1t6J3zQDHkbUWO99kn1aYH1Xdeg9tE
lCyMQTvytoN/I7LZRwMXrdSi6eHKX/CAstP0D0xncF9KEgdS9gzP+JOnZGtZb5qcQberWRFz+dsT
+XXWAroTTMkEHi3EMB/1Fv/Jj1H1p/sFrzx08IDNVEJlSB70uWH9tAL5x9M5gcsxNF4Y4QUYqdwU
fc/BRgbC6WdrJ5v0ZOY9Rtb2OXGxgf5xbNwo4Nes8cgz9ZsXhbmDnREB3ydOJAGyUJqFj21iF6Fi
HXMdNNx0V3U03m0cBUf0C3HjN0Kz4583RfkNlYN45ED82KkFn+VrAmKWMnygqZLdEA1tgkTziNuw
H8KIXB5w1Mk9X6GmOeGQAVnjUMH8t2ZOEMa+ZfXz+IYLkyWOvV2ZYwVnfaUAc9hh5d3ijYlxszfm
pfBelYypze6IXTlppa9xdYt2fG/wEW5ZufvhH0rehH3mA+w7DMumGqCP6hcOpP1TiLZmC8fv+Tck
qgSmaHg9CYx13yD7ZN/l9nAkjm9fQ5zrwdnTSjAQo0q7JTTqCGWMBzna0Kp7p41hPe/oRVMQONno
MKxJI7Mok9IN5nTbj10oBBBg1NGTBKw/kC8aDLvdj7tawSYzB/cV3xUqvjIiInokeO1CgMQw7uBD
UAXhnCipB/BIZshr3+FUPUOeiAYjNEGL045rip5XhHRoyC/btGd0hBLx9wyGSNVVqHSnik3NgCsn
ErFEjBHzL3iIG/WCM+/x3+S6M6aSwffXu5vTKnYfka8P+zqhqND2a9GW0ttoXkJ6QBBnGMRzlvgx
Y+hC4bWTtSOLf/RcjXcZf17OQa/DFRfsflF5fct+XWRwzKWEn/EYE1mDgVg6WuhXoZhs0ldWgfD4
C/6Rc9bT+BvTgXXg+QsEc+k2/ewOSlLnaZrQGgN+w5RKvfqU6vj7AixAsYyhR/tl7JGEG8mPNca3
VorvYhRG/kZbCzas0M/+kzS1aKGDlV9+54bB5IJAPygsZzUb35sKB967gOwmI39/hL+c8Qo6Zj87
hQsCJI+7j1RzCr48tn//s3AxCDlRzTq18quomZGNTl77j3xk6pFrDziRT/vBqoVEuSFU/5iy1CHw
szssgmjtKZWOFmrnAkWKLiyqAu+J24h8hmLilOvaQG0TeHaje8uI+vCfHsCZQ3wEqyYQ8kJn0zcn
FEV9AVePu9s1NExweHog2i3lt9rU7fBNvt3MiZmJXqrm4bTCzTDZfyVkv1Gvyp5SqGWeu9/CeoCk
Og9vhmDDRl5cvgB+m5dPPFFJZvo6S135UGOdZ2P3c5S/LKgX0filXF1HpwLSEEYFddT0YlPselHU
8YtEP7gDxarQuDJkFM49VPsKD2IT0R6KG/j4xr/mO5mbjwTyyADcYoT/WYelgDEuIgFt6CH61jMJ
oQGTmWy0Sw949ShN5XikmYXHPHpJZSzDfr0eGVTA27tPgo66vbCwNNre2K0F4qLbebeYCGIjOSJL
yUrgRXaj8sDCjZ7+TVgpx33ISHN9/5FyHoTgBpBiVCnopAIy5kIYtry4ZgUdX2SMlgV3KUOI+HBZ
M6RXh638r374cylcoVQgyO19FX2wbBHLU6E5YX4WXTcV2vdlhHKIMiZlP4HfR619syRNYpgC8K7x
10CYPDOMnNtjd7v9UDg/obK1jTyTE7a+W1pqw+/85Tr38+hB7bK/he5doWrDsXjyfmM3/ktq5EN5
tYcU+lO6GlhAvZWU3w8QKPowJfmEgb8FnOLzdUS/4iNfRDSHdURvToZOzZrO38BU0JaAq2WMiAMC
Y1gGrRbOB0wS5xZsMsf/zPELdZ38TTwT4fIle0R5xuWJgvFM6Od1RYAtH1ogsZTU+oZPT3BVYGpv
cRR7jkHY5gQQnylAaD5hyCk3phEnpvlLGklfYBZ1u909jL3xQGLIN2BJ6QoSZ5HLaAvoKHwgGb6X
J7p6J1sJrf6zVGQ876zMyIBncU0ga3/Z+nGYTJCD6p/4CKtrdTj8mBpBJkL/hW5eyWjssFkuB4vW
QSGybe0q8VvEQR7zHIFduKMFz0SQ+wNGBsliTygdYPRqAcaSWAZTj2quaNdIl7BoM0BgWP2aNdbN
cDAZknnQXf2+J+EVUQseSw6nxJYIuqRu/FkxMeRBc1Id7/+ct8YecGRHNWRRfBnl/Yd2aBBF3oT7
H/mOkCIfdZ18qKIsVfHXVl+G+qqu59FVJtTh2MMrwUgh2ZPkN0bdBrvdpbYBWVMpC8PH0rDkLnpC
wNa0LVJEdYb9CH2/q4wItcgVmCBspenqX9MZthN77hB+jN4Sdg+WOIzMb+QR15Dj0hC8bbHptNDK
JBecX8F0yAf2XrRd1ScIO0TnR5ZAs+90rJCfp3zdGqnNf8v/RAjMkfeUrtPDTD5W6z3o6hP3gACg
1q+kZMRFOvZ2j4Jp/34KJFMte3s1/Ev96D/2B1NVGrp07AnvRIyByXvmPCZAAGJ6gRiltyOhcEag
g/JGg0hXQyFa2J62IKaHw6z/2nghjVhDtGJG+a5A1pHCgP2y0cnF1FWrsthy6us+2Sz3tV/MMKQd
wPEVWmWaLSlsJUNIjn8wVEmPAa/xjfyvYrqtRpFXwGmzxzecgJbwFCGmRoQOMIN8A8vgd8pCTlj0
G2xd7Jh4Onnhd8bqEvSl/RdbBwKR3PK1uw0H2TfE5NeV13lP2kCPJlFyDIiMpQtDpHNpHYIWAY60
GVDe2v3vUZN895yNONmjbV1aCabLI1gWD4X7+d+97vu7PZMAcE1h8ZmTNQZH+rJnSvZl7Od8jymD
vVsY5STeI4kSTLOTjsbirfops9tvapXarlssfLKdvBKifhdm0VKDuRjc06A8DxdP/KUfWLp0uLNs
0fZT56DaRD3C94lnddGSwTKfzdMxam6bApZybpcyCVjImhl5nnGLHkP94sKtqoGFm+GxyuLJkGyr
FTb+rzwCCxgQOxNOK2A8yhwv+0xM6HwJG7axWbDDkwLFVQ+DrgHSaXPqilZVAyavr1X6MkYXYV3D
c29ejaIArunNl/7EgTJJZRbsY1bF143c8lGJHkJ+R3zpRdh/9y+wmKvWqlC/CwrFt/rwZ6FqpVpN
7F7rOaZUhu/rWYj6py2fCZUG3ukUE6PhJwZEaC5akQMlCnzA6Pn2zfU1BKTANkGSqHvtGU8ISSlt
czUtbfnUEzRdQtAvInkGiJO1wdmn0E6EZhiSvfkfZ4xJFMDdUnYZAKNRTpleK5uFEWgaOX3gfQvS
V9pHKiOepVARAp66BA9z52VrHWUyJMwGGgcQeqh00iMTx3EWw64I298XqXr8/BmZD1fxSrf4o7Cr
z9IEGeIysz61gvKNDaAZW1DeAYgSzGCvTVYxyEWaCSoDyWQAgKcjbRDuka/7bTSh4x4lICoI+AvA
ugJDdNgg0NhXbJ56xlxBo9gbOXEqwOWFWvDtBU2XXBW25JPE531xMRRhTh9f2rvBCPjPsn8vjmbM
IpQeweHRjeWfL+gRUkFRntsi+YhouwmjIWdg9krrDiGrEHNGp+3eYSDsoKExoj9e8GKjHy3+zL13
wP9r225SyCKqcYbM6zh6q/ry/XIsoTY37GKC5nSBHbGXU1xvKiYRMaKhqTKaeQNbNADwxb54uKYN
aMC1sHZLPnNP6sy239XHkFY2UGE0qqAPJ4vxBFuC/qPgEFd6RMD/MU7lvPAAXgtL4fOz2mxwkW3V
LvTRmXN2eYaI7YklrRibx7Ls4xFXz7i4nsxRoPE0MJDFGRBm6C35LwP291sZunuXx4G/i1j/5au1
8N3IAwB72ysVrj9p8Lk3rkzF2/vqBrQqva1fflnH4+KjnNcqDpRVO+PPl/rZ7oH2r+947kGgqMvV
LCsRslWJkMqjzGCMY8sp+uZDzUgsqgjQ6TYkkq9iTNFh19K0T3dTTSNSxGqwROoBZnqvJsJ3BAnG
EPakSoFjtDIt03+c108nYE3fy0XFn1Mc3Z0ftc4PNU2cBA1GFfPxs6nxavgWoRC/EeJTWhJt7YAE
HBB/Dq1I6oZzdVxbJksxLzeNjTmbz9isyFH3M08kFm+hurz6DizfRPVVN1J96Ldac5bxIAbL+tub
YQ0sm+6x/zgslfCC3LWzQb4jWOmRQPVh/YJi82cV2czcJV+dOsQnIykf3YIK9REHFypSe9THbAgE
VMNXETRQeQdx0HE3kTPapnA4Y5xEjGrudansSLPOukiqtuj6GshCsO7beozUNZgUlXteu24Te8bx
nrPXD1j6HVsp8++jQ1tDrfCtwh7hI5wc78hTWEREFnFgRGDlicEx4iOgdGzLYN3VQ4ItayJLINSY
/WVVy07fH2qGh1NmmFvEu24FZYK2+PJJMT+yYvwkO2NPmTeRnCblDRDTBpRrAwJNVc+GXjKlibWg
ODvut6zTnoFAqu7WTPGffJE8Fep709qhLC55mY6Zitya3OPIEULYRHKjUlG6W8tEgn62gV6dsWhp
9A5sifbxtM7QZxWyO4M2x36PFV+kCaDEfvNQ2/mptQiA0V6BoI+NO3L/9JoNl4+tAScO0Vjkz20q
4L6ZgyjmDUndOzmB2Yi1p+FGbRWhlSI9COuFwkFPpGxvXmCYmqlhY4kuHz8eS83wPsD5KXDNlGK4
fDXgnKtF/ruri72y2dJxTOqVNGQDdInSECW/6S7pzkl6DZQega1RfzOK+DAvG+rkAg0dFQzQngsx
FMALufkLjqHAwTlb+iVrn5xZl9t88RCUBpo1TXQ2gwckqGBQWZNXkfErW9A7uQUGsFViHoPoPQqz
Fk34RkdbhniMTucK7rbz/ErHvQAVJKq8hNida6CaBrmkTzDIzJb71U/sifXuHQObGn6f+bRh7fJy
4gtYum0BcjpLiDVJMRcVE1MwfVMZ0l3bpIbK3i3PX4DapMFmSGT+fnAosAiEWH7GSyGgygKfDwLe
SRCNFgXgZ5i5y0j/oC+voP74eqN/Qzrb4DFjAANjkbDfvi04EnY3j8NZzsas6HwQE1q+TqmAZb7u
UPW49c3LZKPbitePFmaA1rqc8y0Acg+BXGJopYtWkmPqpd7mnny5sBTfwpLJg/4cB3Y4wVjGuPpD
DozKN/EjbRmh1NnPnJkdQwyVR2bt/FanLVStToTT/YVJOoGM+gTN/hg6oU8+vhd/J/wIujypgRG+
SC2R8M4fiLUbfWjSMqnggw4QltjQzsjfiRbZkxSFMixuQklYqYZ2a2p0bcfU5qW5oQWzZ5OpTIq+
1hEm8TzwsAb1z0RtIaQ8BupHbcoWpocyYTUPySa76IIknJRAZk4CK4oPkr3szhQcy4cd7SVvOQqW
fvUq8AJsY5Qx1EoRoW3tu7Y+q54foG4QsSv5bBgBls+XU4slymiXKUV/QEnCeTNww4k6IU7MQFp9
fUCJnJs4Jf4UusJhqxuxIWbIb/c47j4cj5cjirVj2GHYn181xfeP6n08EKF7ua8+1q3czok8f7vp
DdKBWUkg3Cv0QW5UNqLCZQGK9cMFZfaw0ZMmHtXu/q/v92uMcwQxhHD09Ai/lmnIfccWCrFrXow0
m6jYPoAwpC6b05wBAb2yeFJ8A6nMenBhMQexfDssJQF7MR2Waiin4kwAKYKY+RPBGITp8A5i8K+J
KtsN2an8cFZY3yU5T15uD4kFu2Rs5xou37g4dNeG5Tr1PjMnSA5+yQCsftj/OrMsorOcdh7keYM3
r8e6KV/qHoHba/TfzWN9PmolKm9pRZa/gI8GWIIYPo+PgJ6oL8jd+Mq8ZiXHv9TnFNw/dDdtdtGB
AkMEAp0YbHdn/GRQqPzuXohPptmrRfSR+g9eX7pIaQ8EMFqRmqR7lyorgyqPy1isnjvRAZpm8k++
/2Y4RCW7aXa4xoXgGWqEmGo0EHvhioSSzut/Y2ettXwDF0Uo+KPp2PniLtGbQWKhyO9lnyfr/q5m
zfEiTTVg40YzA3yoeHss7V2TVzfqpjt9K02Rt9587mUX3sivfn4xx4UIfnx96ukt+xqV+JjYRHdE
Vv+pTrfPpL2CM+M71uqklNPf7S60xHFRa5ptOS5cuUXvfeYShsJRpzyRnqDEPbNowLGwROx9jgZK
XSFOlwZfKgUT9nkele9bwrEmQStjsgYKk/UEMHsiW7sOgioelhPLSYBlvYwoN0Avf16YElWVHhkz
8UleB7QGSzqDsCziDmFy9Kzu78uvjg+hyzy8uINJsNlCemEzpp5SpLRQjyGcrMmRmw/9K3vjN5IU
MhCTelea2XrsE8KgVoxGI8HSmJF8xQyJ8cmlYK3Ypx36h1EMQSLiH3gyEP3oPtsvTAUyhbngsJa2
w0RMlc03/e8/RXIEywx7ncXBkAjaoHBVvnFZfwRJau6TAnxrA3twPK0HzRdaqjZwemJ1nO7uoen7
w3OvTsGbX0ul5kD9yL8Qrs535J9Jpn3BsNuTgP0p7zqGS79kKWfwM0Yo/2KOlxqjLP8vrX9/mtDN
lD8lIY7nJwQ6HU+qhJA7evIidIX0VyMWu+GVdJYdtKgry97vLPVngzRJLPUu0qerF0Vmyzpy59+X
OdY6m5t2HjK9XnIFu8lKGCo8gaJLKj7TAQeUa9qh90k42vVYtL9hWKWrJeR+4ONOzwnvyCPwONy7
OzhUlusl8ePgCElzkrrWqG5SP66+24XZLnsGL5OuBpjRvRU4j2StXG5lWpHKFcA3so2E4O0t1xqI
wtBm72cQx1BRFsircVbcdgSFpFG3BRz49o6xtjgZwHMWjgjJbM3eWyYsNrbodfaS77x5gAccCPUu
cU7TcP3np2xvzpOLJu1itLa6cPyBh235pGZYEGHdXgM3SiVeaWxcEYnqytCXUAVaQXvKx/ABsMZX
1swv8EG//T7rgQn+Bq1jTZztjN9nrvFzqt3zBGDuZl4fFwzoFsZXNHOwQ8LSpVHWYCRlnV4jRcTd
Ywv02RBlGYTPc6G5MgRgueblA/ZTKZcLsBapjs5H3vgqCgAnomrUK3pbSYW0LXsu8V7CjSJAWtta
jwujB0xwU+mgzab2CNg/KpMhn/RIG0UVdNS3SYcTFj9TC3TuHzm5lDUmdkSdhPUG/z3syf1kDqy7
LqhpmQ9WqkPxUyPoOieDWRViYAho7z0QgUG9aikr1gXAUykFlzRwHaqmy1dF3YuxQ9ctXq+AFwen
07Lp1RIiqzzy3tgQRAIW0DAjXdbiyPbL25SZLa2pX8rkMcy+hl21Z86LlsS52aP06MpLnUmA9Ykz
H7E0Glzs1+mwVPglL/m2pEs+TrO4bUV5nl3FOFdnbaO2cz5My4FBmCJvwetU0duw1bt/3qLjaWsj
Md/U41VrID7Kv4Nb0zopf7ugOvPuBaNK6njGeQ4l3mgYUKybDeh1/Fj2jU3YIAkKR/yTW19Pgzf5
+qRlM+3VODM+jZPruSbuDZ59alyqZfYoAp3d7KxhNJj+Zf3Hai+2D4whQVg6IQPHnahDhtVT9K5x
7LXllxcIgweqdHlQc6Wqo5lwVV4x68yp+cSSCh1bBg4WZtSWjqTesDDW7pFSG2lXalfoV0ztlKAZ
rOvxDiDlDvQucUj7/aiW4ux/E8UOMZCav2VPFqle2PZqxMiBelNAg7O+uJ8+OjNhodPhhOGCKbYZ
Mxp4oTnheMBSRYsgUGDAGe7RsImVMgnsJdGEpVeLdOws0ZsYW0MgzfT1iJhgOnYRANUqPC+l9GY8
ajOVD7MEs+Iec/HrTeobKkBuTWEDwXnQC5AFoC9R8Wv+cqpsABBnsulJcMpouIpt0qHnHXfzziU2
BBcQrCFc72V5nERe612ohadxwSt5H61SDGuptGRm1mij7MzBpyo6spDBYxv9HJKZNwNtvkX4x/Y1
bXsZHc3i68Ihg0miv08GiO+5OfL3VZ3yy+Jcambnh8J9PWMzIL0FXSQkDX7UfcpEXsHkD2ngT20p
jy1Zegp6eJs0Ny4F4f4RiWCyODeVgVos6WbCQXuqn7F9Y1ZvgloLOlWj3JUuJ0BMVCLUlDRtZEqJ
bU07oHiCcoqMKYEe6kN+GOD4BVWJB68MhsnH+1SCuQALTUpXprwzeMi2ktQj1cSJqhpKUPg8219A
I8vvGnGTaluJ+2GzFfmL0wyRczWCUdcJD1XIO9agq+VqllWBw12koerXzGWhrn0U2V++6j1m6KT9
5tZXgdUXwraIHUcqQl+bUt4sz/lymD++gLQ29RMRlttMsF3mXqgU8fH6TRaWXbibLXnaViwp5TOD
YDjyilCF/fOOznQ0XsXrYROfIhG8oPXb/ddMknXpKyckVB6JuNSgo34no4EWJjpdHlRxVMnCPtZ1
0tL9CXqct4m0I9ur0/o647Ea5EdKIKv3YLMd20wpw5/IX5fy5ZCIGmnZkKJWXh6BWIxlSd2Rog8X
yRru1TIs7cLFCqF9BG4HbXaUZtweblxID6hhKa8Yg4AFiVKr93E8JqCXqNWTQ9yvMYi+G1w83eVI
MqAnk4gvKym7lsmAG0mCgEyWob9bvsUHZJ7uTSSTx0bDmX67BYEqLFD66FUduffJaIMKzEsvG3Yo
JQ45Nhp13xjeWzQxmY80vBHShLC2u+SA8PS7Q+SnC4OST/FFQ/pKdhMmyH03uyI/2NCuS77YMtup
Uoy6wRCK2mGfOZe4mvmZcD1nYHVRpuqVNWksSdHP2Ik020JmsXaUJ9b0mx6IMf+BG5mOzuBj+BxK
tF7unRQySawTq3UdjDzVMBIx9b0uL/43H1TLUyIog/3IY5rvavKFzEdWjjecl4UkPlwmKAjEo5vj
OR8QUmQ90iU3YWq10MWwK0FnCpvfBc3h/oRy6t6cWeS9jMRfpq+FsDxORh0eJGLRKelXjR69PB8h
xK0igvDJIMA92MfZW+rSfLCI4GvVVHHo1tbPQVd3j66dyD8FgCbgqTh5Lw5/nOFzkiHh23fqUd20
sJgM6k1S7fjg0Bb43/EDMk8r0vn1WRK3hy0rzlODCUuGDFTieHf24r9FW7TcmkckILYv4oO2z7//
IUqB/9Sk+XW7qlIZM6tHQQmKEk6fIRJsEi9D4hyFsp5gdIxvJFckfLI60n2vj5HlZ4TUL0/pkdEp
y0/P9loZES6Y/PO+LlV8CvxzaihCe3mX8/IyZsb+d51/2Z2IXDyiWmazeVR1Vp3A3ohzn5RVZYHH
P1Nn1DhxH2acr7bqY6YdoPRWaTHHqKBk7WhGrQKguEPoWcRL6FV5tBV8xtSJ/17Z2p/ZW/qRt7Tm
pKYVvlwHLvCvieWiJYw4k+HmS0UyGdc+N4pSfNtJIACbO1iadw9/OD184wU/+cG/RM9H7Jct3wZR
Jo2QslND5Z8591YF9G08rZZ4Sbt8vv2x/q7L1Kp5gniKm/YGR8L0R/C7VLzpRhLLI8Z4kF3kL3zs
/Db45nU1XnIExZ1hw9qjWV2v/rpEkxDyB/j08shnBBAFaqHRyy3RUJrF59AayU9SZqQ9AUdQu6a0
uKvXn57Hj+Ef4Ts8OtdCx9vAd6iWx0xQPmN07VCfJQOpD7mCaMPHlMVeBdhoxfRcwyORUlj3afWd
RVYDn2ARJk/lAxPSkJGD7nMzGYP7YN5Dw3jju7IJEv1XW0Zt7uyu4Yaq88YV/m59i5E3zHK96BW9
Lu2ATooyWrwu2Nzq8tR5xLHdfmlnUdX/ZH6laSf6699pqKkpUxgDTUVq7i25etMhkhLPeUGlnlKe
jaipYLSFOld+Ulpy5ItjCoO91KaSfnaVsBUH9xHOMSCZYecDXujL5REQmjlhLYBleKFadJ4TZQIG
ukt9Kf9drVDtKIX+6T492NW/cHQIjEQmI5ySUVqXqYTGDUO8BtuLZqzQpBvx01cNLMx8FU/iubPb
+c5A9w28iU4A/C6XU5lpoPY7A3p3ghaXcay+x9XZvJR+BNLBnztxE30NpmShumfzWU4LeKKQv/DE
SDJ/I2VnmjkkeRI39VNuA/j7MFAYP2OCL/IYLRvfeP2+CqplUa4L2xJje71webCVHHyJNyWoX10Z
SLaRidAGqtP6DTmAp1uuLGNtGIdvTEIWCmD5Or1fsbZNmw7Eb8FJurSrYYiX4KpcTjwE4XHoVTyy
MUs3aD/hhyfKA2424tX3ymurNjjGxv9EEjrvajSCpJ5EmTjDYzkMGUL0Uy2MQh/NA5YGCkWM6tTT
/+l0EwX72O+93oBE0rZPrQCzA+bndWvt27FXwbNmOnZs0sVryjUaBXhSam3te8Xnb4cO44zHVyQm
D4Kc6RLizClKsWRhhGnsZHrsWTFWNt8vj8w+1LqYqjGmkYBBQaMZEdcoXE5dps54QSUT4+vfveLr
NUa/qOS9gCEP5yIohOGOABNQEIXZ7graiUb/MK4zLn0TgbJsOGqnP1rOsvKlemx0jHmxlxrlRBGo
Dufz5Tp3NXVcegZamAoUXvXM9db0wJVh5GoR1Tf22ZAr8jejqn1F7Uc26TsyRn7ah9fNT6YzeRjs
QA3Zws5IikuZiIRFUygZipUEgXAomdeDBrQ6/1WHtomZijjJCTeJwy2WStrFfaY/IvwBrE6vy05T
xg7cZLtlfmDua+ngc+s2zIt/rXCyq/rSrekZjHh/UFypHWnPtG+AqjrPGhExn8GGkBNVSRRE79Y+
wheKn8bh2W2uFBCUEpxhSFegS8M0Gofg7cTgKSAHFk+KDnyTs9VVnzcFeI7X0RiwRu4yjrFHuIHR
IFTgHDhBzOp0VKPj5vEzKc+EqjHVZMhJFBmbZzfajnk1EBh1ZEDHdF5m6FFk97HemGp9vUY0kd34
DkY1DUIygNb5uRDvAYYTMTLhgr6ZyGWYvhbxCTH/M8OxaUepeZUSDWcIVXAOxCSe95tiCel0GCdR
AlzosJbhvGQNeskBW7UW+zo0DbQS4moo5yQ6A+Y9y9p6LnJQF7X6EEXrF9b4g+IHtbvCP4uzFcJt
s51qEHQH1tm2NPjakwc7S2tt9LQ0VP7iMI9l+0MEEKycDezvfcCLaaT9vGCXXDZOBABcl3ukch0l
wZk9sMS1tQY3Lxo/nbnR28ffMhRWeNI8PwC2kT1NymW95L3KdXTuR+kFXRwOLbTOKXQHi8KC0Eqr
lILeeYX6Ta+/Ve9FArQtLmqi+8NJa8Vv1/syAyspuJ4zDnx9XLg44oUKDdRwLp0WhSg3+iY03zke
X+hSbpP1+QpTlmh33fXx90ptIfTw5pfA3Ar8GsBrZh89CYmtCLnuQ3Lewoyggo8cYHt0ETGs5dfG
kf4M9wIeJJyM8OaxPl+VZQ9DHJkFLxLuLMIinceUMrtgFi0ePk2/oEiC22IPg/epS5Eg27597/ks
drPm620IVtszEbt5M6lTFHtP6smOSDIi9IHd+7ifIWyZB+eC1eupec5+eHq6RCwVXUq6sqFwOry9
kl7mowixmamEQuqbyh9DlpMGqtdA1KFCw63hJpHUfMlAIgwAHxWppiItzCv7OdymOq93B8X8kU6Y
GfV4KXOZ6X8SbNIvzGTNlmwEk+rnwNcDXcwsPm4XB7QzZMtV9KMPDbWQVncl4Aexu4xTO9Su4Ck1
pR7bIVCLyDPO80LTQ45W6lyUl6OxE89zoEprZ0ZE7JfJNyqQKS5pWN7Xec7N3FXYzrzl2z77cxFw
9rHDW/TsT8seXS/kFyFY2n1+8rg7D0ZXDajfwA/9kvs0SoiuMVWDMNw7ChvSZcnFo7zWV4DjVmDw
vtYOCZB0oUXHiZhbriFnClEL7yivmPbm1W6voM6WEY0pnQ1E/Uu5ogw22pBRVq2xTtKqDfDARegg
CF+3oITDY+MPC3CzYesPi/hwNaOmeaO4bdT+L3G36M5EzjXrgyZ+MujI8kQhvtg5Ap/8f3Z3qWt+
fJOHBqGDKrjMRofSO60gywwLGDsWFbirs/1+BasKF2sYddKOfSqcx+hX3mJP5/u+fJYotBqL6Yrl
LdOLeR7aEK0VyLS8FW3R9xgeP0WYtFI7zxFhwvlU3NtIc8gvjiHOgrCuHWFuKb1+uRRHmw2Z1z6Y
oqoSYLpv2+bgZSeJKXgVrHBpYCROfcxrQMyWJ2uxuUVWumkva7fSlJgGUswREUlkAu9Hd04ta6FL
UzPH8Uce/USCz81ASz7dGS7wfxcFpjeeOOiXYlnvgA1nAUlogTHtBVxMiOA8HGaCfj1zYN6c8+Hv
rOKAoiD3LyKcRe/z9G+MDdAbdQCsv3u6tuitaMw4j+K2abjhKbZGFep8kor6lnVBlPopihwXCKDW
2aT0AMJeS4ayfapdO3t7QkoqDkbnuern5ShdQtjX5XLtekLLMS3WMUkuFjiI+By5a3PAVwuHBAcI
o+h3IeVZjqMcMrPjbWAiRVDJitZJiRCSiwmcKEgCTZ54mE/YDlbh+r3KwuGJOiFnIi/zphUNLAIk
FoJkno7k0rx13DuLc4WXG6sbKXVXcbv0vip016pQoRUswyMlxPHTasOgKVlEWhCpZN4rtI7kJNTj
nSjiflwK12DAVXrJKwMhvp6Lx+oiEvNR+pSNJvzPeINd9GEkh8YBsCTGY5vhZiZywczefbayBvt/
FN6AI7mdxxnmLK4r29WWlrNlvr+XZsAQZwpxbDA5FZtEipbjPn3FE74P+CyZVzirgexdfcETvT4P
JSc6VXYWW8hCY6XLImoQZK2wYzg7XZzoUqxQJJwKnqsPWJKva+bDh+SYdALTpQ0OexrOM/hp4RkF
WDr0uiP5MqYBNWuuEUbN/ObxApUlKzdCXq3pB5O9Zwt8qQHcKqNaugM+0e/NCOMAkLZYjOls06u7
vHHJw/6Ki+n0wxpgnry3v7zWbFft7AGXoV1vJHpHZCFZjdQsLnDPhgv4IWgOy+0xPR/xNUVyHvvc
73eYKlEdH5eTwq+dMnUMrH4RBfSKXyrW8OGVgBGLEoiIsV9x7iogi/xrfI/ur2rSWLmSbx7u6XV1
lPEqXBEEWvBhJFW8SBsGoNA2J0NhPVTKBL+SoIfRnNlb8Sj2lNNBtE5uuHAis1qKbVFpMHSHwsFf
GKHcbn6y3Simn/eNz1LkGkGIj7Fh0qDp4sW79JWmFDccCtliTfZyztLJFUp7CWE8/5Mk8uPI/mpy
BcPEybB2/Fs3JAW3TTcqRfFVErK4SiOoYvSxZi+VpiQFnnMMQEQz8OqOxk3uEt/9HHTT99ZLI9l3
hQuyLECNFzhzdkETnYMIqEzhcnAG/FSjE8hdpp0VC0U0Wor2zDa7KO3b/TYgmvbPVfGbyZPviVpR
7z2QKTvwxz1g4iQtfDrAhxA+S/OBP8P5c1wyvnPEfS1S20QIRR4U5My6vNK/6gg4vAzwNbBCMkTp
og19N6QsD/zJuiDoStmthY6KaU8lt9eT5+CGIlyBdFXXdCpRWgpiihmqwzWBLeodbud4Qm0ohoIR
71+CLkvRuouQPxXCVsMlF6BD0LeUJHxk2Dv2FJzm2/cewyuSN9Akov+CFwY2BqW2Lwn5Z3cWsocB
vD19Jfph8axAypkn2RxQX/haI/h2hUeOJ2uMvAAvo8unf1VTSKfiBCYC7NtyAxnZK6TAptW5tgm5
3AZS783fP/tCc8YrhTn3UaOZbhoQessFwlEYnoDQf93q5IoTh5uFZTnznWtjE/8+jUVL2NUdV96Q
73dWDjT0JJuB9EizgSk/OO+P8yGXvA8sbRiGi31c+bVJR+RSMhzBXyksZ5e98LikAVSy1TOVe7+T
05DBIXKWE/q8MfxkbxpBjkAd9Jet1owLxLmqWJIggCDQ8kW9d8eOHS6GpImIiAV07NHaeYdr3o+6
nINwapewai6ZAjDZQe/TIuaIW7LRk8hdiPIOJuHwQ+gdP2cyZMLA/gta6FsXN8WKQpMkriHqiXhP
Ryj/Nx54k2L+UVkG2QXYkGeqnAUtXb4Ga3+AVHSBI21s00iIaCYmkNsylVWZCR2K5ZlY6S61jgrZ
NNcr/79CldEVWLNG6w3jXCe2dn+S+W5fiJvwc4N5TsMW0O4y5LeJjJD+vT/ayUp3HxDwKPosZxmf
unSLNd4jzwzblPStutMHy1hJsvlnh/7ftWecYMTGry6gXx3qOeju5n9P4fii0RQmBldEUWKXa5Ry
QYBMWM6BvmvRAgYs6IkvkO0DlKpdNeE6S8NdsxuTpNQxIrEGg30e1e+2VQBbq9QhLtAaOpKJVbMs
Cuj/08HChjm5DpNKYiD//IIrcs53l+5w7UAZB7aFrOGYmeC4pi6h0GFwvN4z2UWJKRX04RSqIwsK
dovC37+fx3gwjoQ6AMYx2B760pUWloWqchZarB3i068NlRcdffVCNNVBObYQIR4hOhkSmUSfVWiD
dI5NcEC/N70hj2+L+5V0aZ2L0cLwHuXKIElwqrDxmztV2Eo4I3F2qK5EpGs4dNL5DkkpqFEzK4yR
DPmkV8Ley75t4kMNj8qxD3AcVxXtmG/MG/ws9KWuYfBEWJAirMLdbA0NCzrFojZLbejmZLfPYbWn
S6EkT6zv9dleVvdWNCUkSaZKTw8R5aOCsvLTI4pEpAZDIHbfO93nUvFfX1OQVpAsVNvMmhv6N+u0
Sixe4KtOWOo44xxYV9C82+vxfSVE9ucfGefqkVp4DcBgdM78VTxFAXUsUyTbQ5Df70qJMrfwt7V1
rv6eImiRUZJHsTONq1UV1rKpURAhvUMugBhK0DfSZkBaaw+jI0a9Vori9380ExljDNDrwXklutnv
K5G7MghYpagZ8PKsV+0oRFG5lsS3hfoP824SC3MycJQYVwq8olnYuuq1N7Fq0UJxbkW/QobKOL5e
p6q4oVDWfrUjNbYRX8lhmqFmdaOiHE0k2LDkb3WLwMn+pw17ZxUpMgen+GXcJoP7nj8ELIlTUhs4
a6neo795uC/ByqbPuu/1+0+coaFhzJWyUwYtclXKfpj+IEf+BgTMcGKtk2D3RgwafanS+G+e9dTf
we4fA1wZepeXlImspq+9U2N5fqu7PtRJmYaMoNN7Mcdbdo8AwzvWj07LLS8ESG6bwxie331wb5B4
y+xOsCHYrDN2KsfFsPJGANxhqSLR9vmmy1BuHH+PhSX9bUfDOlTURr1coYsKVR8hQpBfjCaX/t3R
kXnm/K9AgaDq49JZUZQ+wAH66RZOx/pCAz6v+9+si48fr+6ebJSN9y4PL4TetqVamHMOhj9l+KZH
UWuY9qL+BgbgaBykvA9Uwp6bbb0efvzEmRDH08fjUF52VscRISWkzooydJaojpC/6BMuJ05xVUZe
96j8oq2/uiy/8+0X9DclFTv4MxC+Ne61onugC8ZIJCFquLfXhVmvxAQPYbdJSvaAh1rulyTmHG01
Up2tSzPXEfEZNCbUMUgYad4Td/2L8FgKmupgLuAeUd/G9tWt6kXSDiQfJXnIf7pjOhDqoazwrRcK
TudZF/HPxmUBRNV00mUqkWP/sLYJxndPTkBnkzM+o4HWhTEhVWGLYQbzVuZKM23sg7+kCAl6TUUl
+sbW71XyMQxrGlLsCJXjV56VqyHsQ1ilw4nJcsQTB/kvHt5VV6emsjllUIquX5gi2VQ890BXgd9D
RcIyZ8knJ9kgNYhdJb8q2ex2+c+ECJanNw0n3X8H/WInlVhWtWjStDY2rG2AbzK7+O5PCaDFIYTi
KIbqYycZO2D+UxNYRmwZp+lEg9pceLNtnWbxRHh5vqQJhNX14sZ5to4MVxs5uCApcSUvxnnKSMn8
YAngmjVBXQHdoqLCIkdUwZpsktNeQw3l+6m9Vtmy6hrk4G2v3uAPxigVC6kstfs9lhn2Zf/eads5
ppCOGiCERDp3pKVBfgnUuLzOP49I9W9oH9/rcoOzcZPilSc24TH4G0cRqg2xjkWTnhqAFgDZgWrF
RFdQlTvfMJ7geqj8NorI1aZn3SHAsTca3nrXKJNfjgP3s5bDSUm8IcmRpM2k7SGH7ELiPwnh9nY5
MkCcZ6mi5FsylAGI48V+DpJSy+ofBxZfzytTSZMizT3lshBkktFsfpgAzKYKL9KAATCHQqBiR9rD
Ibs+gZ/I8bY3g7iSwOzUBtYC9zDz8m6ObX+UVJTR/zGRC3BzdgqDfzrldrHaTjTQjlLLqK3xW8GY
XPkZV/IKxHbHNJ3Lld9BHdmr3/QXI5QEclAtvlXCynMyIM8gthf47BGqJBLsGylsp3Q3N+GVU7QJ
51lNOTlLJHffrZ5dYQgVBcd06ZL9B6aHrhrr8IafK1TYv1K8hbVAg04ensH23NTZZ3j+hFjMj1lZ
HlgSpWlwfbG8aDFgxAil70v5GuiH8nEXxKJ4MA05ebqCAYdmuecQa1grHgQLgH3NM9+O1ikOFW9w
KeFRtQa5H3CbpuyskfPeyiKVpHorJcS/Mlrd+UmSb8g41j/pNk6nfXXHrEcIwYYGFB8otAkaGnky
Wmit8pi52VNVCwaTSnrC7VB08YDRdvwTyCsDuwgPXYT7NSdM4owdAbFwfPMg0YyzoV/dhGuFlb7Z
dncdNLz3Bb2e8juJW9qNYT7TSohMfdULxAGBHM01uMfZleN0Qe0AY0WRDGwh7t/XPPnWrqA70Pos
yFOXxFgmhTkRxdWSkxZXJQx6i3lUUVz3mgiIZ0ZCy94/E1wkf8Yr/zUbBmDcdqb8xHUkfdSjcJFH
0/AavAirvJXo9u+COzyRc6nPwB3atGfFMjHakF/s0WdjiVRTdqo1mKTqHY5CFC3nihMS9MNHZhU4
KCKvdM1FavFS+4DvD6ELmp3dyUHau8HEWwSPGbBHnvaa8J1GjoWUu9vsuz30QYMmTIcT3bjSGxv3
NBG7ECjsBYHY5sRy2E3XSaBUtvwlbp5BUbsVvzM8kTS8Ipa6VsYRODDXKS5UL5amMRYSMfriyBOk
2u3A9jnhmRNIXC5BJvyfIaaaMnL8uqWr/Xao3zBkiPyJ9hGE33MNyBHp7Yrv6PdwjywTtKOj485O
8LE7Lkx+6k+BED6dsrXainuS7dXn3vyj0cAHJyO5swAmbaQZbnbbqOSr+69Pa5RSi981U5xwMIq/
y/c0p7/NfoYmwcnFKaHqnt0HnJ/IGJo/iqt/MVMHqyPH/CaYywOMxk4jT9eZWWBvM/w89MPc5soG
6JX53LMZCjDkkD93niAUZ0GHPMtpxV2Q1MgRYxquM2l1MNMl1WQMhoEBCZErZAvvp9ADLRMia/zB
auz1tK+wJbX4JGghRehhn8pFXHTvFiUix0FaVuR/HJm3jhfRsLRT5/C2HOteyRafe+/tx198da1Y
G5xJ7wk8HpS348zyOIuw1JCLEwFnOP0CFcR2eAlZrV1J5Li63yE6dq5aPbzsg+LsUr72/kkFQGJ0
ImBXS4qC9VxiEVXgkbRm7cxPYdoDs2Q6cODnkCbWphS9SM0Jtj796SNpvnjmbLawocWJyjsEA5cy
srJO6mgsX1Ky7MwF6pQoWbV1V7NXYq86v8jy7mbjiaMD+JbchGD9/C1wDWzjxEfFKHSmn4kV0Tv3
H6DnwaTh2mxnjahXud6i93Iots1yRpoHxbTEkstlb7PaJGzFOc8YJC0WbGvE388tv6Fif59MgQUO
0jUGtDYuNA64Tiu+AGp3nK+c0OcGT1N1kT9E/jrj2lRmZK2fOugzBQVY+wtuQLd/6RosY+1J8fBv
IdCmAgsOVrFGeLr+vyXZhIuv5MozQKaOMS/D5JYZwe2ZmB08bCaXrJ/mSM3hA4vtbOedXM/iYepm
qi5xl4pXd7qVr2S4JpEy6REkGwYLQ/hvr/qC+gM7LWUJ/Y44HJUF3auL+JzGOaq5oTYimfsnBOe4
UbFi9ovmmhvQ1ybdMzVzUpKIGreT2G8bnZAZOkr834Lh6g40SnAjqMhAzwKUJOwGgxf376ZiklDv
ts+cwVw0vUyt5UOl2L4GBL4uxaSNEcbPROtvZXxY/BIqzjhOEja9gT6hbXxcH1SX8Ehkk6hzk6gz
zLaRVuhLEE6gi3l5LMER8NXM1dkvmjqcVFtwNA9vXMPkuOm1iwsom8EGH2HjSrogs1HFpts1adTt
h9U6mT8bP9NmzaY1F0BJLvVrJXbXp4etdJL+eT/5asPimKr+6qv0Qu188CSWKrYlDyt05zs1bWKb
UEznNoIpNtJQi97/hmyZTq8sOJ21OeRFdcIxgmYz6vH2NDE8yxvIGPIfRl2tJl3O5y37FltKtg3K
mciJ4i7T2RSmD5zPTUyXXBqdKIr2w52Aqtqt1v/07qz3he0U+o4XT48qgCtJLIjoqOlY8SGCJ+KO
HbfUQI6SA2n2j++21iiBnJPn/z6zHLCzE5OlAR4cD1pdSTxqGQjMj/7vT8QbenjlCfoegKC+XlBq
/Y6ulLv5UJvMBVdvgaoW1Jd3toTfNhcsZtVirfzUIwKYzepZuBMMY7HZx9Ia/vRFUBDjFrHSuJ8n
ys6qaMXkK9iJSLbpEz/wJbl5jvlqlDWBwRZGAsmpzS7B5ccb3OFzBukijxWehTsZzN68vqqJ/guX
ww3jJmfNnJUJlrRZm2u914gjBvm64w/dbgsukP5YO9SysqTTrGCrgGvBjrWXzplQSbhJg2IMxbRW
954ouzIRckEQAbSVMpGJy8as9z+/CfUfC31T5XQuuqXBtAxFZjfDEJwO4+4YkZqcfGimcEJXemXE
TEKBnJ71itVgdIlDPGXXHqyJ5kIbw5AkoLjC3o3nLlxTw/+68/+xLWhD5luSijBilXq/wZZa746S
rle+0h58f1x/8gjfek6zNuTTpdWxx/GZt7MrY3pBin2n5dIp2XvlnkSdNYdt0EH9J3jzP4mgYX3l
jkX8A8AOHhRcapyOy8MUzJDNYT2+vlrz8roQ/W5rAfGA5GJ5/ZPASTcMhonfBOnFzIszjknF30DQ
dQ0MVuqmAYrYQba5i9q6djFBu6Kl8EEAWOW463hlunzqnOxL0dOEjRFUdNYmEiOEb1NdvvKJjOJJ
zcovAYllh+DTeAhk3Y89UxW0yWOsqLMYBGv/V6KwpyiADRu77BaKOP1nqo+5uONfKsR1EUhpye63
tdTR8REix+zQ+WiDD59BHedw9+SgAwCd515jy7uB1ajqCh3/9IfsCXwYfx9t7OM30ErmtpD97cLJ
MyTfkb0x3fPeSUyZ78WHHyGdgVxCbhQ2YmPctJ11/ecfiXiEbAaZkmgwx2gmr4eNp/DhpaYRijrP
U4O9jjuSXLNRj8BJVgV7JfJtPp7p4s1WeNhvZBHMlugiSa3Vhk7u46ZNyRVu2PQMswwT19LtkeFA
oNoKvFY+sVRDjbXa9NUI6phNA8UaKO5oWFV+FbCQBJcElI86VEEomHS23rAcdM7OVqw3TGwIIyWV
Oj9sGlaZolfAIk8hGVcEk1QBemM4KjeOCWfUpNm1DOQLUhKZnnHeXUK0osve6OobNtndiF3ZeBgY
l5NgPR7l71QNbwOLp2psgCgn9nuvLzqmV54swNwPH7RmqASINOEgjIx4HB1LxsOhFKpcJsmgPKb7
i84Cii9c0PYQwnU/XiJzJZ1aLjY+x12d/7PTnYdLqAN+QeNtussini5DJqhplQE9XrbOUcCciF1E
D5WxwbBt2azkwSg+EyTIgcto/7N9g8jJt9treOYKlY519YQW2x+qRxkP+mVoVtSodIYxQ21zRcIn
7yUsTAJuvQJbVqXiFulsnAKUSjq/5ett7J//fK8FgShZeZNyQcuTABD+JeO1/n5cqZnI9rTxp+kD
QpHFqhRmur5BkBau3/AXgoMBlTVwL2FjlQY7QJ0maJDhS+AqH6FRcjqJO/ctLFYukcbAWtV8+W4E
yesp5RFwoXOOzQTUQ+9dUqQJNoLv7O43/FFmSrTom+hoVk3q/B9PQX39hW3FNlt9jcaQW+TB3lRH
Oh5U4CTt3rtiLigDGuUPaVE1fr3RVu/0VO0/wjpyl8tqyU9+6m5mOiJntRBYD0Zw/DhZDaRCVIoq
swSUKaeRgllXPLcYebZp78RlJ7A7E8x+e4vy6CEfdI/kShAhk5gOVVrpvlcjgZ5gBplauYHf8roH
ouwFtJFa6sEpykGqS3fHaH1vYX2Zd72U1/uvfsexnxZya3Us6elRUyC2O/y7dkbkFIgfDcr5wKVW
Vjn1SYsuMYTVBBWt7C4GNovHMhqdtY8rYy6kBmJmL2kNenTd7uzIz8njxVJINQPbQtcQLemQg6zy
KafQnz3OJFxUu1FBvRtRpVNw1C/rXO5eaSg7oT1Ai+FZvFSIbLq7PQeiipT79rxb10WexF1rtVMz
ImBUct+WYWMDCCIWuEFcg/khK9cZdNAT7DNTrulBqaIA6kurN33tWQXdPYkvwSPnjsM9CYWFCPam
US1c7vJSapS0lK3gGzEu3PaqoqxaOwZQF6Djcd0i0T/o+D6vgfMZC123qXRwdTx7q+8B9TFEK/8Z
ptMl/29CNnzvqYGDlKcl3wtFpSQg0ZuaD381SeO2ltBbMn9ivye/XdfmmxWgHkfKFKLyOeR41YR3
r0ypzRCSDmiHV9+9vxzqawtdHR60Xh0wnxEKrjhcq9/jLUSPMKtXCgUsLOih7pamwj8A6A9qxyo1
sSih/1u20nr24qRPDc7C1ArSMpXJDb1/w7aLQGGTZ6USwEvJU3BiKzFNJGWlkLhDW4wcNNiuV2Qu
NAFyrLbk7bHaT2HDqtJY/HbUlIYbhqWvVtQSaHrnwzgmJQKIMdmr25OxPQdzVcDX5qhxV3+ThbN/
4lhdYrvuvAAkcB5h91EVj5HsCtOaSLPTgYRA+d6+T1gOIiOqNqYmil4H+Yz5Ib7s1sNJuiaDxecb
+Nk/lDAhWfuEo0//SyYOARpxYnRwLDrAIG31M1tttHtSt215MTjLtFwqtE/rLH7IxHfMr8GkO+h6
J9wytGMEpVRJucWvVqjFdR3WqPXe6IidPpYs6HYjlNGlV09tOZHg5BkaDc8P4gVynojNAxNAaAr7
wrDuNScLXwdnJWIW0PQphiqyT28OAkbF71QJ8u769U1BUi2MGZfUtt5VrbSsXz2FaCkYX1tpnzRz
yA2jskMelFaT5dXs3t2P0VOWYvagHfKLpISuWmjJSg2peSUwGmijZrGSAALFiky5BCJO+I0d1AGx
NQFbYntp8OEqptfu3QTu8cIBylZ7VcNt4OrLRKA9zNRQLdfkwVpqq4UjDsFPmh6j+WLN0PoIcmcY
vHL2qhCNvw0O2VRYt/SQ68s2a1baAuJKUILpI8VyTOjLs5XawkyPEK8i6g1JaZdnIctPgqo8RnCh
T8rxSE4rIa3+iDuXI/k9gQ5x4LUBHvz5KG6wW9RkIJJ62dR6h9sE99pazQHWmYy6HUWOj4eORNS3
CdEjWaOYqhEB0J06xOD914ETOrnBYKV8gtaOR6HVWWzHvIReums0OuNKedp6rZtF6kVwG166HJOJ
g9QH+trWSBBWOTFZ4MGIWkvZDZNO9OKCa5wuZN8qooEuY36vHQ7qrSKRIaUBxqs/kVvIPJhm1r5h
y2mKDr/Z0w8he4g4PshJL8mGSygTZ1Gbs9Au50vjsduYiYMo6iQlkiwW7/nQxBSoaDhDqrXA/S3B
/94tuPHum3VsSpprVTBwZ8a9nU8GIPsxozRcbhBx1wFLOc9KLZivtArLWfKe8y83GdlliwFeAKvQ
uaE9tbej9/7hyXIyprEwhKaZZ1+kLpI3227CvnHXqckUEcMk6oh/hhDLCtBg1uNM9T8zXXDCQdpA
3ZIZtIilpiqaxd6v7Nbo8RXyWaPMau0+RebyQ6TP8PBM+kADcis5QjeF8wfwqWTYynyawaYklIQr
CHgIO4DgrsAObRzocTwNWh4WVpNGjsUwNkwYkHKVMhQmRnTaOvw2tDiZqLgpQ9kGBf2UUsKbZAfM
Eqn9zBH28hKGyIlfVkIaj3d+O38pQE1PCf9e0sPATxz+/CXFCxZrseqssVi2Q3HDTqG1HnTrWNsk
Ufdd1e5l64JuB3DfpFtwAK9U/9sogY7luHWA2kaaw2rbCLVLIn0kpDzk/euw3N1Idc5V7RK/ABh/
Fwqx0tOVvR0WWiyUayRN9lmYX4LRtrZCbiQYbGlFcRyc6r1HtfpWp+AQPFqsHlvvOrwLLCIh+2ua
Zle6e5hnjotlKfEX9to7XRgCxvaat6RsWQVwTQKsW5sjVGysfzMG+yNCDArehWvbn/IsESCNsnvr
dNcWiA78+6TDkrpW0IPd9u7nCB+RgJm7LyuL83O0nwdxYla7BzbfY0hPp28huicc9ptut80t2DK1
1JKGpv9ziTJJP/YHT6ev8bJlsNmjzNHWX93RQP1Q+FPV18w0SoDxV3muTcu7NYdKPMd7C3hRrpxN
WPlqimNG6ygrQY9ONUfz6C2rgIo8B9etmx5MlCRA7If6gbi4LgsSU8ga1b0l1nntpqVkLzEQ8tkC
gorTXSnNQZ56uhNb5E3jddWY5Jv8xMwzpJOZvKzIDNPRM5xkAWg4XKVkaimlDBlLyusXm8wLk2v9
GG0E290u7AZG7Nf7F+Ak945mivBsEIgYt7XP6RxLKcfMmQ3pOXCtH2W8s7ryTTUFpCOCzIfTjZFS
JR2V81NXTUUWGiX3pJ4gaKlcAmkSICYAJFoHGQg0l8DEvJ9ObDL96YdiAQiFz8Vryd0XuLZ5UogK
oVrRJEFAO7YpRODnF0MLdD3aSvmxbKzuwbvK3pt6hSIBQu5uHfRjVpnCXmvyTcJsHQB4Sj0jZX0E
ebhHocMZiMoUNYOODeabDGRKISW9bvg8rY20tU1wLRruMUS1rQkW4ARorqKY7awhVrWHN3Nd/vwV
quHIHqqK0KebkFCcf1/Tr7FDaHXG9fNeFztVlbKM6yFMw+L3H640SoxApTSulsClrrxQwE1mP/3G
4oUe8Row/oww7NylFRUdC1ULKb2ePfj24b0iMki1S3+qEZsMqrP6ayY5Q/vXkWNt1VFB7Z3QOqpS
bERd43xjEhsgh6IWfKtpO/RwYbCLIcRe/L+hb8SZOBAHUPQTaJxehdNUHLYDzVcfFYKLuoWaUbtY
VxtnQgxPdelOx3JUmviDG6jQU34x86K7d1BERUSPs6wrYFqGnjnqUzwj8zPOxmoFf/D3h5WpSBeJ
bWGp9in9yXnOvVS+df5LjNgbXAsvsNZaSU4u7RosNP/E6ML2jUQsDZatx0godiuhXW8XLuNaXs3U
b8Ts28xfD02HVZehNJPVMmWAdykrUYw0ULXK022Nf8tOhEovgcBHIVdlIU6YI6EerUDcWhpHerBB
6oQwZUBZSG/1anYLvZz3SrWzWeXRiRVn6Mu31hAlRR9jcQx8TgFw+0/1Iee+54KJxdg5jvrgCwiv
y4rTHc2lBidnUKiwbPX/R1ojrUqgG1bJ6Q3pMFISFcsbnHEFLLPlJhvQkUhahcHPxEEmfkshol98
aHoSewlWhYanDWb72DSWiBaijwCaODNbtaL/KABsrrn4/+7hQizyQ2rtKhsqBI727O8Y+xI9KFG3
wytqpnYprhBAx8bJAd9HgSwTp3+kGketuTSU40T7IuO4C/gWZjgLx8Pe39I50geXnaLrErn4L+Pf
niyMBVwRg5Xs53MX8ee3y72s+/4oduzDcwTf62iezKHQ5J217LnEaxMlLnywAw63tRpTQLb0Es7w
aSy7L3GjyIizx0D8PCQ0q6Mb004YE/YgzpxCGPS2MzIrgeyRo/98LaAdMq+gUCxHMC/B24fxYHFA
wfexIfrOJrgSysGFoRGyIXrw49D5rAQ+QJoxYajN/Ly94xjVcl1yeCd0bg6if1+Kwan0zqxE3uQ3
NPe9ePrEV16x8PyA92IVqrq5fyZxv/qrke2ylzIwZU8dcPuIIbGGOxzeG/PRElfUVLMIoN018qlF
qMRHAi/RUqBKBFaJvWYILSheb/k2IehTDMDeW9Jp/BdSqAHIeySTT8jr4DvK55jlo/U79iVFjNJE
inkwmcw677IPOVHMOT5Cz2ouunyC+gWS4N643H3gYNCGUULqI3yHEAdKjoifUaDAsV0vcmbkf31r
XDKJYvICLS1GxTY8wVDIC1RzWrRFBUlkQcNiO+a4lQuYsds5FJnn7VmzSJEufp2+Ubi7Osoxc5tK
idDJa6rcA+rW6UhffnXg+LxskGppKciGRtlpI2T2VBPSKQj9O5+FWW631B8a3UvizaXFe8Xbenm9
teLyhHtorV7jvNC1aLLbm6sFyj3XOMXXcXbEXSh9i7ygDlWOPGdlYpIvsymIk1SF2bBoWucm+wNO
yCDB2NlVw7Q5JsX+oHJ+5ck3UdVxjBWr22uVPbQ7e/d6GsG+SZ/VeGIsp8a/sqsfcWjz9LWFYhCw
xYj6nOkhFgWyzoDTXbrLMlEEwEuTQ6YYUAvr/zpCPEbVKKNEHz35uPu9cT51h0LQFOw6FL2Bs1Hn
fTOt7Wxtge2YS33ChbY/rL1IeMaFtZjJSv/bwlJ6hBxqdrkMaMLvQIuHdXV5wd6CsdOiOlj31mkm
MPMl2WCpqLQcwVn5n+djzpnQhZ7oDBYgklCt2k0kHf1fAF+uyKKt0eKfcI6/8O5DT2RGilagXa8u
l4zSJCsfseDqjh0goHg6lJg/iMxsPVbuscMGkvFM+kdZO0ML7IoZ5A217ckXDxHHQTCojcx5QOl0
1jvUlyZxNa+0QUx1UoAcfLINvTl4PF0WNxYnzYD4vXqEar5YD4tiHPo3oEe+GL+lzoSJ9SbLS43G
v+CFZ8+jTGiIb/5BTpvr+mav8iUKsQOFM7OvvEkQAEIcTZtyES71ddDOkHGP8TgxpMM1k6bCmgr5
UYzb/BsC/Xf5uW/3W7/Xf/fE037atkuBLRRiwDQZtKbMR/YumDwhef2p2sHC/yejrYlVkI09HLOl
p13tAW7EqC3aUnlA+9BqiIEm/dj8hlY+IOCKpNE2LWbWM0k8eu0T63mEP2EoAeZMiHaAzsqBLzeJ
q5o9bwLY6gfJ86tTGUUcGuzfFikk2WS+4kSrSKPIUkAlxXXhTmUf70WnbJ822LopAGrdY8TcyOwo
cEGxQ3eJ1yLAhIbyLNrZoIujZko0du+VH1kK2YzNAYAM+Ksivy7takBIWBpvRe0wzHSvO1iunKrk
+VkEWcm0QVbIdktnORPyF5b4Xq9AhjuBeV2biJsK1pa2gxb/jE/g4mrfYqUJI8teDcFjWuj/QKJp
IUnFg53mPAjmdyT50o0f43wJKmNHR+kpCU73TAwDn+6XVydFyehhWL4AYsDRUSry8qq/94P+mQ+G
DDNJI0e3QaTWQxAT9nPWesY2N/cxJCzPUEHqYzClOw1b++0YB55oRQtRdLEAxbyl0A6jB3YdoBZA
fi6ISN36MDlybmIyknEzbiA9zo2udnBBNGkuiZwlF1KwpMh58N/KyzEaDrKaB/NFj1SgJT1ExH0Q
I/XDLNG6aQwFVs021FnW9Fn+XeFBpluHNFCrGekHXnL2aI8NpRJNHx//fdiB6hB+++eHqcgj4nlK
zcDJpGbMqlA3xxkAX7sCEhFMGeFDpC+nAbq5SMKlpOtJ2fsx3QlAI1VifijsktgKGW2sX6UVwT5t
dWLDtrn9VpPM5goyEkTzYt1/jGcv1UkzHczvi8934Qe/+Smhl4xod7QRev/oCPZc1dxAMbgOutTd
rlak2KI2DMFqEXyAvAUEhSjuFB2lvC/VkSKTkaC1vcTBnI68f9wlLC+DujQqJBMj9cAQKDxFnmWb
NPRhOEodx+US2M2mLRMvyQpGyTdXewlxzt+ND5TfhisWH1mDJYYi0y4XZOrdqVSc9IN4BUvgKJDt
m/EPsAchcWt9fSpxZy+pYLC+b6tYN29o/2I83X7r913RUGKn32Wq/8nql6+ddlEAlzZ1FrM/zEFI
HayNMi5Qyhl5ZAs0mLx/sZEng8SfopCrFyaIEBFIrOrNJXE4//egApX7byaFgyWvud/auqTrHp3S
6Lag27PPUnMxYDRUY5AXbL8IGOiWy1H6WUDi62FLSUq6QBKHGdYapbW3j7LOWdCkTLBGUQNee+Y4
/tNkyk+ZSWphZEZrl0iK8ixsK9bB482EIBgnSUCh/xfyiUj7gXjw4Z5MsNbjbYtm6jA6IOnV42hV
guORYGn/NoCK2LzqJ81AcXA3mpE/AllZCJ7Cdpoe6G9tEoXBgz8uOVrKdciGnCBSsvdLEoOoDLMS
YyMCF0QhcA6MGvMbQg2u5iAbrhnrLMS5aHrQKCvo8sYjwAXdgK6lury7VJJsggl0K9vZ3onibUET
dQArRRCPMitYP4OulmyM/CFmB5x57shXOFzXLNWbkiOWYiwMSlePcl78lHE6bkE5XZvAxXRuY3/X
Nt6cI/Iy4VY+iaeHVMsValJEd+wGpAzYvL/1D7TQqOW9rKYVr7ro+t9lj1LLMrKV+qhR2HRVHj2n
a1FZPmNEaT88Rh5HK1AGoChu5f6ccJPlA77wC4BGw3MqKzaZi9Nsdoz6LH+pPwMv/6LJ0Oam/9Fm
cEgmdV5hFN/g6lpmzyU5+N8zc4Eijj4lqty6dH7zkg8cF17O8z1sega5u4Hpl2MXBhxXEWHZMxdH
zB9RTNfQM6zjT4ScPGQPv4Q7jyzdHml3rkSRD18vmAiAU1cCE9OLayCFFGJkDcyGb1x2RORijLx+
y7YzEznfsdREWqw0+rjvHpixvurhuvl0piwYQaflKrpLQxhleCmjssbYO+pnqhqwzYWfN1T4DsLV
9xhbMdwTxD3vpYN3SayE3JClWZBw3J3J1DjbpSygFylDc0jab80YEId681DO+DmQ1P2lAxWgz5lz
pFa+G3kJWFA2N+AW0PzbYGbWpNFjNPluTROspY4iaFXnDJRWuKncGSiD8d7jVcktA2riZrdy9t1t
GPTer/O41J+eBhnnxm6PCq/ksyNcX3WZaGrpFIrsaKWGFmwvOY+6MmZBGqu6DQ5PtzJYoz6JiWC1
6qPTCDnYW0ElsOPC5B6m5GREwgqVGZiWpg7Vl7v3/11h5lWPtfY4Lal9tAnrL4llDBQcj5xl8dal
+tOCP9/D9jZGMIlHzk0b+y8kNF/kXoz+hb9JjXJp7urICh4/xaEh65glXjzZE2N5N/VqB4jV4FJf
vDeM3pcw60Yevj+ApcctQSmM8iQ4ID+tNpjaj7SQbOZPFIAyG4X8gmm/3Il9Td5hVGpFztRySVjg
G6T85mvqM0L8k6hNiW8A38ogbFAt62CqZGJSGag5uDR21pRITz7tB56ujfKPVzQLaOWMy/236LJ5
JiqmZtgDzxKK9euBn3hg1t3rHvAMxG0XyS7pbQ5XSsUxomNVZXeftFyxBckTmXSoO82XgiY63S2C
6Us6zUrxeE83R44HAWWO6XhFQ3K83c5A5mnyF+nc+9Xj4YP00/aUGJIrYMLBOxJ1J3bYkxvtr7Ga
ZHLHctAwrijkJ7KRvtI1Lvs1rQ0Hhkz+V5kR423SOb+lOrtRNU5UsAbOT3cFPqAV6xgdaZAciD6V
8nQWl061qAE/x6UFxAMxjgJkvF0oO7GnfD9pXXjleDkBgJIgEdhrZGU2mbJfdW0S0Vq5iray7pa3
8LSbDRrpfGoL7NAb4sFDPGFjy9x6rprxI94oBFpDISOz5ElT4NCtp9+GvW+aW7W5CgXweHJJpVGy
oQLnQFI0dWtdiUJ7wRDoKe9CK06svpvLFPh44x9GOC1nfa0swNYkT3KOaB3tj478aCZBbLlu3ViK
ymsRKoO+rTaPLMzDoQC4cx8yNSo/shhJs/ImJhpd2K6+iezFwKbY4SsVn8wFkNJfA4dCnEqhl+Ml
uQGXcMLzfMc4rJsI47pLzG21ek5A/gdLN4QogE1aflF9QdkXYTotH3MgXwp+JzcbaXyEmXaJzCkY
S7uSYmb7b/Ziux8eOq+qTKPU3JJTzvjZIoaWV6nVp64WBZK1BSvR7M79d1BYyNblHL4pZfoyMOFc
HpgGOiSmF/KsKkX2xJncdHRjYpsnCGck534gOEVOpXP6FGJY9GWaQ/nb2vNJgmMXbWb1LAei/ToK
g6HnTDGy0Fa7igGE1SMZ2cY8vYAj7eGKmMjKQmYi3uaP2PIPzi7nXTc9nGQmaaPuDtav0ZkgXCZU
c59OSyVqgiAQHc9X18s5DMl5/MqUeHQ2ytijy3ML4ItTheNACSkPmwC/8+WoHGhbNIBAIZ30nX+L
u518WFATn9EQQhMKocQiW2WylOA/UjiO9i8hQiuYdYOz7+u7dRi6dK2TJbvu9tqD5Nos4sA8YLWT
pWMu7eRzIMKeya35WSifvSgSOriXQrN1OptbxaNhHY9iL5EtZbiyUUXHb5Tf6k6K5b7PLlKFNoOB
HEu8Tgvb4gQejn2MRWipMWn1dUyTYSyemg679pFeHD8L7vw/Cm2fG43qKcHd+59viXrxCym4n+Z6
CVkRMd6jDTkmCR+DeWiuje5Z3e9iP4NZyKG/m1GGilpANTRQn2s97OBh7MGcpM9ISARo+o/WAFAE
CeW7RY4BtidLtxFKYfxvVWgSbElvNFgQghmLYMqvfxNdciAtjBSk94gS3CSXvVnZY2ACxUJFTFIG
DIT73HRpsRvb6dg8u960uXuZaTAA5DjuwMnyhDalM9wxhLQENIf2GJUAQFcG1JJhSXF2takt9Z/a
g5xgw3qHea0Xjs7uGFqZN2IfX1auSuea1W36SeGdzRR3KD1IWyScyjwltQGV2JqpNxsImvaFvrl4
dYX0aFHJNbdgxFrHezbogKQMju00J6I0tcx66VAnyteS7J1sLXFnJEBm0+dWJPIN5S+tzqEMZKBz
f43IKNBGHhUq0X8ZR7BN1RqPxkWRVzN7Ni+/k8Jny+nlqaGwyOWSQaEMoqUY9tgIQ1vVsheMdK6Q
3tb7E2bqAyX0sDzTkGekGbH3EiKeqRs8O91JuGJ/F5IHgCZsfluk5b06ZyVaBV5LRGWDqoJi4lSh
RrPzIXT0yhmhepioqzmxBS4L8w6WOkHPB0bwNWHWSa9MASxTAK/jQ1HQyI+EoUKxo84OTGWFaEAU
BZiPsUYX1QX9qVngssTCceavGJsICoPuSo1NKLSHI8g2LdWEGpsIgP+G7CVBCW/o40Bh6m8Q6CwL
e5FvXMwrc3FUqsqp6UUuoj74ha8KWDS1oft7ZLyJUp6Mal/nzE/4DTQOl28nYiDSYe1UNSEdrzlE
m2qv5HPhJ6D8eZ3se5Rr8N5/NwxWnKkw6Ebl9IR/62xwVLJQD3Plw2Em+Aob+kwb1Io4QSxTqmE/
BSfJkvPWdcfQzI/fmGgvMuLvHoxU863O0kCWK+Op/CxhJ5TF9mCFOu72fZUOQ6+ROOahv+FhPkY7
q0PEXAayFpMKUYSKk6ksY3ZShxZAqKOBBrJes8JKSwlysNBtK3ioxy2F4gKo+ITjvMNTDLPmxsak
b2ExB8+7Ad+4cBFRJP14naRXHo3+bWhP3GJ+mhGz7sAiU7ZAmFJ/ezIEj24cMjJerI+o9bW+S20u
aAdjVn7UEGrEy/0JjVzMKe3vyOrJTf2u0nCciDS1gFOIMWQEWhKXI3L/d07Ha3c19mcsAjJRvgqP
4G/uNXzHCzdpjASHAvQ7xXeCxgDKmbVyCYjHLD1iLqPhp+sbFiejvm0aB+UZnae2GhU2Jy62HMy2
p+2HnYSchgIZ+OBXpHfpZmAs+Ze349kwP2P459sEzWxPVAEl0SYf5XN4PRM8qYfpxkwsbHL+7EhV
BwCnZiQjxi88fX2LjHK/YPJPVGK3bglYwgQ4XcrlFf7yhfh5OZUy5+Ulkvc+s3me6xi2erCla2oO
NzKsnXWav+FStCvXNvT05+3oDkOwR6xFOQpFDq7kVESzrHm0swTBcZKDrvMOIXmtkbxUU5Te3Pp9
xzbDc/Y/Q5W1wJ88wHFdEdqqLMybwzI/Tp5QllBkZmVuUyjV12bE+lA5Gt97KWNlgBsu/Afn20gT
rsBFF8YI/cWH4D3gm8sSmMty2i3SHdOnBi6MNPlMxlLEdaQqzOAgoMxg8VECVFWStEtV16DgUlvH
Qjc+Rj45rEzgf7qPM0XZ9ZLatQTs0/s+kw8ROtPVd5f/pZsS/Do20cBaijzRxe+5ksdiHcJl/3V7
ymXOao+kMFOntD3JmlNheOZmPVBLnn3pkdOPdygsmvfRW+OgWCXFsTWCKATYOnIaOdduSX+h519B
Tjld2Bvb2tj9xu2OdzrcDQUY8VrIzc8gTRX7oU/WLoneWJFRI9LXXhiZAGzSAU2ryDhn2bQ05M5v
1XF6TUZ12PZ6tHISyoewJtcGRkS3ElhjmppYztjGx2HNYflkV1z7Of5crK+JLYHgqsKGuJs9cNkM
PSEBhwi2yjCtyhPucsikjDK4OuxVS3HLHDITxt03rsiQrTX8yA9ZIiSeeQTc5etRcr4mo9/QEo0F
nmha5QZwGMESDGKSy3/B9/XrZqS4SbkaTs4H4VUw6ErhurCK6RObUf1OHhafRjKDG5s5/8fNYgKF
nl4PlNGIHrb2NQ0h33b7bdP9MBB1nHhW2LdmrL2/BsCXNdLJ9ihEdZVX+PmghD31SKFWfCrIDSw+
CRWz/Ve2tC2HzLc71Ed6qgL2cRENzKr6xI5Wj2VxwHNZhe5h85IoPzWhMp9h4O9ms8EWhyX4h/qZ
rbtDS8aHY/JG/MOZdQhO+S9VMQZFUfJbAM3E/1qNoReRPvNSfa4EzvGnYPsRsioJh0L3SCRyzdB6
5hHfok3OC8zCfKgAgq9jSzffQndkN4wokov5MVqPv/+QptogGbQATE7i6sYHS6A7j+2B8CysQpXW
NsHufpZuCc/VJUZWHKUNGICV/O6UCBUJAVgm9JyaAGNseoV02gmFNC29ccuKrRsbMV2MKxOXOTUi
hocTqhFwvWqMrNM4nLHkzTEZaao2f1Sxr23Cm09j13JJNM6Bbrq8Q0ieaTnBIy53xl6q39KIIuI6
cXX6YtgK24dCOJ7k7v0AfyOCZWSbS7z33MKQz4W3tV0VqSsexub+fF4mg6iA/IgX51thfbAVgqjv
u6//NKqohIxK2itLatAqyE/PxEJcMuQUlE/KXk+HPJZ/7pw26Jc+Mw7JcfY79a5V9kN0UCWPmcBp
FooSti/si0IOnKHE6HooG7DptwxSrhGTtAwLaBtwBVTOeP8APqUl3blBineSYG4Q+tI/R/3AnT8r
cGo8VjsHWosbUkmRa7gFaCLrX16Y/7/R2Na6uwHDGlzRzx/rjDQjVLP98UMLHEe2UYBv0lUM8yYY
3UN0VhyaAf7xzeU9N+Ppju8RH6HQ6tL6fuiO9kVo0/1bARUS/gTemlCUQp5AwsZOdLXHM1iLJDJV
5/DKj4+T/Xjqq5cYy02SFmjtYDLAvPG2UYHF4BdkdR/5Uacy65nb1WxwqQEhoAgWuVBzL167dznm
qziM//FHSHWwFIlzegYcKhl4O4kvfCEbtzCUVFz+9TH6ydFLBb03N4SPG1DldMAgEj13MCqDHcVe
nYk//Z3hDUNItzSKHrSzKWpBv6rZ2KZOOnHJ1fptcgTxkvO/stVmsVUQv+AaWXc5yIwkP69XLRJx
1ubAk3xJ4V0vrdpWB11s4LvHqTwSWglPS1tawV+YYgGo34K7cb79z4MEvnUhLyLpl5d9LAQ1AJaJ
7/0df9zuytSz/m3iHtxJ6ChVIK9q9WeLki52prvwYbPeA3u6JhXtiERcZmPQt3B/2IrEXiq6Sj6u
tUmHo+6og1hWuJALvizC6ptuXSkdCm/RKv0YiDWuXgmV7eV6IVyotPXle8Rk+86HgVGnGL8UGdP8
sxRCSsm6WaImxwhgKtyztUYxa0lRW/HYVigIhQ4UGkGG3CKGzC7vLJ4/jPI0oc0P/vfjoV0imNGx
GiN2kiWCb8bpelMKFquveDMSjf9CrqCwSViuinUOnnpjuBioaN+g3PC7FrVV7OVYKDjqFY4StcYX
g70ejOC7Vd0ScVJSLaXtysVyy4WeBl7CenPo0Q/1fvT+DbJpIT2v9Saz9I9q46LOH1XDje9U5Ec0
bc+76SjGPyqu2JUF6JHkxo/sPDmE1syT1FBAveUv0rWIo0O6/pTDoRgCV3jweXqCrIeGbPBuuMq7
HjnPy/MosGynm8UvhIlqitX3EtD97dNOHHNOahAUwywtGExhOzSEdXd1vU54MzsVC5SKGsfpF55E
fuVt6REb0/E+HzmgQtR2i8DjYj/kK88zeZ4eFN5/zaPv2b6KJjXGpfI99Kx6NQzLHMQ9b9Ktkxxm
FRq+a4aW5bO6gahNtliBU8i6aFXHQ5uI9jP71krCVtZU1FrH6S6/enUaX4krsSjgjv/LgPKhjr1u
Mw4SGRHvSK19RzmfEvhySSqCFxvK1jod0wQf8zTeqnZFDtVNFGuBaBZjzRFfVih7olQqZa+K6zxG
Bk9f3E12muSYXLE6X0iXrH9/0NB++EmtoHV1Vyd0kaa19DcBhhm4olfyiw4hOP2FQerTeQkky2wZ
4o+PWN/VtIFhpVMskRqsGIdMiiaE9A5d1IZGnejNPVaGl8FzrnNbaAhZGLuMJN825wi4aLSXyE4W
V33KjegJKEFg3XSIPmxszBcr3RwKW8fxo5/X2qpO8Y5eWAVVffZPxT0F23fcIgNVEDuTFrZrl9Tn
OXhnmbQLNnlWZ0IzpkuGPyBhDZdv7M+bNCsMd/pUURfnYcTAdCdq6cBT2wsoKA5Il017iajtzWc2
TPxoYCkJVjKMySEnT81YnkJIQ/+zqD6Q7Q34HdBhipMlRqE6hg2mAGUjjjGddvEn49r0gQjcch79
bwZ1dttCi4n6TIhglG60KGBRsiYHBXfxMeeYc+pWySo74xyzFXTfeI4oUJ6ZKhgxBHTsD9GUCLwE
M0G6IONX+QBA5vPfbNPiKDhPP3I89B5tVMGO245gRzfpU3hE5rMpymMq0lqLirRTIdZe0EecXHdR
xYEMo4wUXL60YBVTdx5vZoTvdn048/WJf6ZSxm+pLBetEsbAng23At9NlgxBRJ1jDOa5ulbCklNJ
Z0X7l6nASIO3R6h4Tr2CgoOI3zOuwfikaRUpC3w7z50Ho/OaDkERNCIeiOsw24W7BBFxtMXIvRJ/
9Cyf8T+LVFCt215z3W/TgcErV1sBDCtQgHGJoSxgRx+nOKkZL5REULGb0ldGXwAIeO1bWh+T4h5Q
0XrPylZseZW7tZ8yDeMWTj1mghPghJAc7IzNf6igkLp192pDX4OHcAmV7btsnfLeL+oB5P855cPE
23fHuDcuMCfhEBDp1oifE0rxNYhwTgbX+cikhUxfj6NRAxvzhxbwC1YPtab6leLTtYpJbYdY+5Om
25hDNladSt8Qo+50l2fX5EhlomwPwtuVyoiU6W0QWWN9jZ4mK+JD3JlqKF+UQFqGQNSuwDwW1Vw0
IzCOpQn9KCeYrSUvlefG3XX92uwF0OCVHz0Jt7TUVUhzCL02XEKYWZt6G0NUKB4I32Mf48z3ej+J
yqm+KgHihF8AAdcDndhOGALeN9/8kmg/VTs5pm+yF3IYu9mHI5kIUAKmI/pGMg0EClcoseTlUjpk
erWt9RmxkKVTpljQ22LiVUIKiSqYdSVf3TZaXLldriyeaLL02l73lfjt7QkZqPzMYhHKm/uoWy8J
ItRry2QMjftcR0FRB2ZvqZUAQK1jzQlLIeD4DjE5YdJnUjhxIzyRojxRjgyoCaCD/PpBo6FLZR1F
dSLqz/q/mmGCdhdKxR2e9w+CPl6a62aO2Z5XVf6Soeh3qw9ycybPxCbA6Yb6lPgQsYqYGltIrKo/
AXPJw1mHdu7znomJeQErkjOjS3hLuwSNlemAGrRLgtiv5utBjzNtt1ruSz2TV3HXefCssHAoK8Py
4msg7YFWav9vcmF4kF2vmVqJhso0D9kzx8Dy9d88ZLC8uUZcEJ3D6dtiP64VfmKvT2R+0EeVZ5xy
VwtZJQRmB4Lhsn/GDdgxBImfUdWZf+H13rY5t1o6hRIpUlq+H7q7k5DNU7d7LkNlkYZXKepgrto1
32toemnTYRNUX+kAPvUQqGhD8pJMVINZutzmm9ICxRUx8ow7stVpVX5Xs0ICBvSH9H6Izbbs4WQu
CFKnzvyIblIQ8nVtHtdVfsPsM21s7oRSkito+JvieOpmqdLTUoYS2Wrhpo/RpEnBKLZ4HpZNmmV/
w4aYPN+YuEZUrcxLkCg2ui6LLZStLQHFeSA7EgAY1OhpLq5eISCHHM3NTAcToYP4/3akPn2Tl/2n
sG7hXU6KGz/3L7Gr5e6KMvMeIbw2/ECMNM0zuUJhn5beqlI4zn/qZkNIzX+SVvFw0wa0rlsQxjC1
FY+obgYZoLKBXv63FMoKfnOiCtlfwkk75sIF5I/oMzw/WgGOpv3v2uiyfXtoTiUbZUnVnlri0mJ0
y0nH+7jZr/SX0ajP3BWdK6owgsX0MAOC6hFjeY7O0fZ13QHbv7r9NBQ/VpHpWC/CdGGtexjwWmdS
epUWFrc6q1UtOhD48JJXS4WM1CMcDzyPpRWib5BUPAn3fn4wkZdUagNFARWjNGm6tOrUKcz5Qo9x
VpvUz+G+z/bCa5rDn8blhYOZF1NVSnjWebzuKxZdWVEhimbhGhXEfHeQCgGGV3xbuyZfxBRdRqOX
YVV6uYUhXe8Fl3ZIuEEy0XjZMHd/MtHFxMysX8ZRbXxxXNKdlWqPq7y4vDz1d3TjCO2H4EqLSuHZ
23c0C8KMQ++Y1dN8GAcb8aRWLrhqkQQ1LBDZI9vj6DiYdHb4bKHSWcdBRxAtm9YREq58VEaNUJ25
aouZ+Fai3mZEkKMLUMtToGU6vxM1iqmGCDuXskWUSZyDo7E3Fby+HGhVo3gHA8uI1y3nIxAVSYcV
cwJ9ZVxHyHYq8TCJreZVL2VUTh2B4tXedfVI366LhdQNuoLznAYR6EH98sALQYNvyTc/oZmyyATj
MRXSXOVAK619G74y6Y8TBAjaTeSnIm+VvgZpM79//5UPsiXkgEreKV5vr8JN2p4DfBXUh8e8Q++z
4cqlSiuH8Dnt6J7j3glrpKrwgpklZtQbYsNxouaqqymi9fkcYCHRt2+J1yAmwooT29hBuE9O4lwo
DdbOB8j7UYVaDdb/GWOb4cRWa2JliSfe0CajIzlyFT9pCeO1TJlzBm8vMK9SfH6Cgdf6aj6pUU4J
rs30V1T8MOdksgCIB/aT3vEG9QyCjpBe8VRnJRu4DcPpItz4DsmqBecIMMv6M4YnL2MFZhKCNK8O
yi2lgst4Y8/8GgB2FUus2Xjf/Gjw8vh8xlzdyqsx/vKlc9XiUOipmMxpp2VcyZ7iT+0tBLmra1go
UckbcLOOluXRk9KROILnCbObQnYvbyetSx9kyAjG5NS99wMUvPFe7pzRm2mN0eqMc+frxPhfWRCG
wTKi7wUxmX1aLt9nn+Iqif+03b+xvh+WRKYWLiVfLTlJCbB79X5GSAOZX3h98MHGLvp4GzWFnQTW
2YZVvV76Z998Dudxkh0EXNQ2dhSCQK45SSftmaStoJMWknVgg4M+UBjTA5CaMZYU5g1uS9Fe8m5f
HJCOutNM5NZkFAvZEAHt1rhJgDsxvGuRkTWZn3VrlC8bw+iAW/kMcHuW2ySIZG6iEZLX/Vl+XLlJ
HtES+1iruq80Fo9J2QTz/Nqnl5ii/HTAH9CbX+nWoK5qXN8b7bxrX2/L10r+qq4zh+UBTdjiuXD/
QvDsb/wnKAPIeRbaycGRlH7trFpB7/JYDBbrkETT/Q9X4rKU5+KwIP1+zwyuyrjwzKViicDICw8K
uANZ0YuSICr88bOFq94EiP1vjQbcH+Ix0KO1VkIvPo1FNd5Xon1y7uJz9pqu4JcYjqI23Vy1qAFD
UdIHIdixajTC7KKMD65Od+5DRX1a8bRV5vvmxKAKjWTdL8jgkD3XKxLjXgog0VTVqZ4nOzUE10DK
KkmrGGoyLbCplT5KUqq1oS9qAtpUzjM/g2/8Si9BwgO9nOgnsuj+9OWTQrqVSFfWIF/Sr9nFQAyC
4bevd5IONUHBq/evBhn7kJBRYvw0kMlMDB8q/AvpFRa2PJHHMo7jxRjgZ3jkL16FzXssj8rdoeOr
6OnM1zPpEtBUzBnJ9Wp2XxD/F+IqQPueAP4xRzbTRs38mZwNP8/1mcYksR0yNRU1u/AkHuriNzu/
yYP++uGR+mTSGsavS7BlXmbjaOTcOmSWdyOepPgmRDghon8PVBJJS1/OwqhPimcufDgFmZIzTnau
IZrU5kHl8gER2hpGUXGNzWwp7rTfgXHVfeizoxlVkoiT9yfIMOFIjrOwBllZ6PvigaGHsnXqOhZI
ghpaGqrS4Sr5kAceGXtB9qtXQYVJnkZK7J1BNbjsDvNugiU6MD4hjw+53g4aQlx9qyQvhw2R+ofq
rtN767/4qlNVuTwxQownM81tRMEbwr3hEIRt2ww3kVQeLmlI5+95hWViEfmbWF0DA99GTDIvFp8j
sP4Fy/WlqrscRxIcSrf0S7rRmwGDQbxJhf9i82c5CiXfomDuTxnxMEn3emT8v4tnj8CN4ivBE2gQ
brK0b6jeKHuCuRIIxKs0VpOkRPtV220f0EyVEuRIo1BBeNR2ZsHxGyNwy11AZ/nMno2WMOPO612D
iRhrF2jwFk23FgXjDRG7iPV2oD2Va+gtZmbgtOz1RLOcjSFRw37R8nBi9w0n5re5YFBixN8mQBQe
SERua6MX4GLMdRNL/ZLkM0K3XlmfvgoV45vunNvrRec53NlepruALrTzcuOBRqTguqIX1kHsMbpy
P0T2YWdkOGYnvrZxQYO8lPYFj8FDsBlHYz0flgf1k3AtCVeeISb0Xx+LcXSJuxF6c6E9dnckRb76
kNrWV+ij3PXGtXLZ8wJ1r0pFjkl4eXJ9jypv2eYERPJ9Wy5BWfdz6u83YuBqlRAyr1FBernzKQt9
gSNwlU4yQ7b5UzzvCb9BK05FyMcpRUSDzvDIkmkijDh8+c6VWK9Bqzm8wnwNbQZnrNsdv+su96yH
9ONcNunwk257efPoLb2rvd4AEDs5pB2PNhoGE8hVPAOrlhGeHNx1Qi7SbLZd/dJT0j2oF1mvxYkl
OaQaHlTaDIbmvzx1qAVVMbckAKqmR/zJD78YTQRuxDMPs6Dhogvyexd1aOAvKWtBHs8TjYs2tryu
xT6FsDbHE4WXsWylDD6dJanpZB3NLZQQW+IyBNA9uY34iFgpcYa7KlsOuLXI3fOZMKw/SEb4LHnr
Mt5a36OlJgA+iZnkXh9BFUKiUwAFt//Z6cn87covDdxp+7ydIzDbH0yKK2jms9ST/QJnGHMdVWqJ
ctc/cdISwl/Igbzjbe1gdAohYbbyVsFI/Pdl4UBGYtwKLZ4QRqNTCbrS4mgs3QGpLlnxwlzeBFNP
94IQnKeiSYYEePPsH5CIkeyFRS342yAnRNnXJgAkUzaQKVfThCtJt4eIouG0WQJk6DcHl8tCGYNP
QJ5Dia7qd8+OC6xhaiI+vSre/G6eoyF3xSpyCwcDQZoCcoBfGWXCEvTNjZ5Jup1778UuR++P8bYL
c+Tr8KNz9QswkLVS5ghlDmD/IPKVjoFtUwxqaIUmuYsFm+/vLHGt+UV4Jv+Ww6loKjouwnyv64MR
MDZqqAB7K0UycIDPTakfn1BA+Jv7z8xBcy4X+HXkFAgclXDMuvjc16B64fsxxnf78hZZgPTRqQKJ
sCCPYo/1mb6A29wvQNOQrvQQtQEF9W/ipXdMeA8iRSPaTIgM7mQELt2U17EuCalqw8MW+Wj81tt9
AWO0fYQztwIyxxQVT+1GEFm4wXx7qfiUWecIrUFufpQ6FUJciHzsdq0dOQQ1aKMBhJR8QzovPLoJ
9U3kGJcVKuWXknN4K0s3+sRBQnnZyg+z6CB2DBa0JRO0P1PxI90xQD9CEDd1da2GENUOdXGw5LLF
i2YeqQPVyBEujzrNRu3UumnBHsEzZev3x318S8kFGO/r74tUobTE573Kx8mXBW3tjiuAyOLKaPx0
7lopY9DKiJZjH4YRcaZDfNHcx4kW8KBNZUoI08lKZIKCHyIyL8Kq0/s0drVxXFiMmzuPhQoVpksP
mco7muB+F995oGm2oKtQBCrKbSH1AUblAh8ae8LHdQzRl695oDolJmqEdn6rpbVwZh0NelH0sFEc
jVdCGwWeDnyat6TevYjlArBNdTIDw4nhyr9lt+hXHKTxtJG6igChVzGvStQsH54Q3POSMI9RkUhU
8HHIvRrq8z9rvjlJp/x3G73SX9M0lNVP0+LjnDnHDtoXfgQDB8iMFg/zFRH+tpdqCN9kv3U58lsP
+aRvL2dwXlvNQPixLv86NcrQJlcfVjoPg9xSocRBhRo6AYQtjsk9rRkUUfKjBcC5ZWP2YJNOkA1q
QHCxkaBwzoZy/BCMmr4fHUSI8c5Uim1Y+Qi66Me0zcTwPlNcw5kzLKBbCFlOMkXu7lHnTZOYPgxe
Rh+ZbQBcBDBbo23BcC3VsLXADcpUitqDZyJeqLI8FwzokMn+qN1evVWuFvIYSWAwShoFP8sdM1oV
bLVNEQEPg27JdToKp4REWAIH/ZfhSnqlaeKWpBVY+PyjZfHKCvQw97oxbcliP61IC9gy6bi9IDvO
jnrBaA21C2nGL9yivS9HvAeIWPrqkou3MXKWY6Xz9HlFYdB1dlSUhEopT5MeipGlqZEHA9cdjSFF
4GBZAOREb2LVi9gZOL4V2yeN3gQeqJi2C/WbLMkICQOoISbz8dGbCAWAxbjaFXGBxpZDUELBuruZ
ch5rxsktW7gpMFr1TuP6N+d67Ghts7rPbaM6vZG342UuPQoCJY35q200gg5A6CKSxzoNpZyrePim
qi01o8SbSLLckwWRkOXNj2cDVvRIP4Gge8HkrlSSRo8cEq22idR5zqwvL3sLZXwFN4SSOrL4AqpV
qS0jApPQkyZvM6wZrGuZlXGlLp7JHUv5M1MlOAUTWI3WImjAwyTI8P8F+7c3CLMlOQJ3UG7xBTx3
XbIn+kbW4ESA1eDvTXNZptoO3l7MA9djzq2MKCPSm5KX4YlEFG8o8lELVJPGC2RmzH8qagY/kLyp
iYtVnVtzsY0K8MMl6uqFlJiTgGxA5d3UE7JKVGOY6ml3sa3WsucL1MYfZM/qzaHoqOaBVyU+IhGw
Qh4XE6g7vVlAH1HIakYmkPEoK2DgqvgxXMsVMrGB9s1ON/NqUw3d0AigmDAYMFnjiiRlZlOrVPCZ
+WpGaH4W329Kc6cBZkgidgQXxZNIyiou2Z2KQJmBDzapcn6drbQy9XKSiG9sshH1Sv7nvvZ+Ovqu
qIh4f8iZqgInny88Thq0QZUS3+nsHIGghfWSl4+XF6k/cNvmj8cH5MlCNUm4zDCNSCbMX+lgjBCb
YNiXUboWXgxnyfyHI8ai9EMJ2l5JYJva7fc6P+CUeSj4BXUI90EMF4XQ56iBdOJ2cwlT2hzU8MIK
iP2WK416i92ViJ2FGTDNxOK+d4/Z/Q9Z9DeIKnJ0yAP3+JoXqNzThdV0aLp9KoUcyVDFsZNVXbZ+
1tqmPwWnRYB3y6Ghk1YOPF3el7h/9BIU7VceidRX5w3ctIBFWlMmdAJ3tvp7KHCskTJdKIi8wt9R
tPVua427OEkS/aZFMOA+387+h4FdUZdsJdel1l3/sPsTzMzbFG5Ko/Cy+R5NeRKS9TdAVP3XQjTj
yvgyPMTZxLU6fZSjhANYrbvDm6QLp+NeE1kh07B0v3/AGzOGv/RsuLCoDNhOkU8PG7j/H/oIgWGC
s+rS6adFVNawQa6WK2GvmLvhV1/3lgLpIxTuV84ysOxJgCmgI5OijnTq4gZ/P3NjzJ7TbZO0jhxi
BanqQGbDFmcv+PKMGxYUZs2lCIzFo2aDt1wbllXxaeRHwMyntK7UxInD7oxAbAmNK0ybccjTs1ST
FFY3AIsLN6MBLEXJBN6rAIPzyfG4CZM7xZOGzfW38H9lvK2Z/laVOymZdh7gkmkmeLbZJquCoYZR
MdCebwhep/5qKEfnkgNdgikanQmFULXcGfOvnsPKDqIxJ56Cw/BW/OF+4So4+Rt1xjHyjy98M4dG
vW72Pd4FOXTP565PmJBO5AbfCvdPJZSOMH/inWH9QgnfojgkUrRR71Ql4hUyGmIba4iCSbxdcNjV
I7UlXIUMHipPPHrMXCfFle4Ym5qFUf9nCH6FLKF7RQMaDkeyp36/Ze0SMINg04/zJmr6RqkttQ/W
dU9KBdSEMcGdxN+CN+WvH/W3DqZbGd+0CH3q9mJiR3gTBPzNNwlKGtYA5W48ppSiAYLe9x4sXeW3
ARaKk35P1CouyP925afRc5sRK8nRmcgPO60E6f7yfputqimuthqARW4wbtMmXkObGnPyQen1gxBa
byov1ybSkaXe1W9YezX/tiZTN3IyXBlKp+odBjERJslg/9J5p154Jb72TZWSBmJf+Ux9Z4Dw5tQA
XBdFCg78zYHBJUafB4YNjLXVafI89Wjett3lnZ5EdJvhU6d0pFpBB9akNF4Zcy4NjelvgXp+shHc
9HiB4fvNupV731+YGinGoeVGP+REmOz8hUHPKF0r+UWY3CoqidlD8fz7ynk6cm1ljSygbGuCFs1q
qlxhZO4KhZddj0k2SmXztrD+oGcpSMkIBQHyOHRWawgldlKymRiPEg8ZFacglGG1FonFP4XwUwWG
a7/L40009SCGmNN3lNgBlGmg5VL2viYV//5PTm63XgqReWytp0BByyItpSYgAMrHjM8IO0AuNeKz
h0bwZBQ7aBl9aLJhq65z9SMGD9OKPDbu/IPSfnvg2RAW0O6XNFVFRGIrDwzhrCVeO3qJYqskwgIq
VfwYiBKOpxQWpeRWylvNG38riM5WS1u72diLl+a+5vZ6gcSjVIiH59ywdCJUO9gTeGRj27WF2Gs9
8eg+ULWcWwOWIZ5Ss/pZp4MCgpKIyhPKIDt/4Bh0aBYAHR23JAMVFDLsfYqHKxqTziJhU2Xuphno
qWgNvBxS8rLokqJ5GLs2Q3PCkmdBa/HnFKE6qX10WcojuhYElmqt/HayrnJwgSdNNcGjnWueWpxE
tqKygqlaCk1dT/nu6tJQN5sz8HFSQcmLliiOeZn8+CqJK08WL2Y33uWT8v/gsjl6Cl82XBZf0eZc
BjZAFtmv9Jbv4fwIY32jj8ZEdrDZRe1eAe4P4Q9OYFRWPlj/2l4jpzuc/ZLAfkgC4tFp+LJDRsRE
IRR1FG2LK0ZRaRauBycYSP2zD79f1b3FcNTaCbBpiAYK/+sHOVDoCO6qr9eY0WmkOP8dtEL3zkEb
qyLOaM522XInV+vAqEVfQNYVz3iv+uzAesqus0RSOr9ZvmHhe1VbvGF6673k0+8eVq5zKgMXv1Wr
oSya9FQ8mmFFULjUuNpT67fWZHSYy3SQ18OiOrm7YfljmlrB7FWK2qj7zBcTNUsxVVh6x0r3Lq4l
LcnSyL3NncVoH9gFHiBi0Kkcw7pdGDeorqljQ1LEpKcjuHhAsdoL0MqNKunjSuATJnsNiMoIDGZu
EFdofvkI9Qh1aQqrbKJd01jliyKwY3gbHoxgn9Ko2lyM/vQ9t3ZGPJANiLeNMh4mgu/3oWrNQiwU
OGv1n+Y73SqhcvV0uS/BX6WsUqcJAJMp+ynMbPpOeuYDjKczRKvYBH4TyeQiL8IVa/BeBcgdELXc
ZMxArU6Yx6sAjI2eipWZee6M9PftYcWeojAMhj5iwcrk9nCFSUiXhb+v/C3B7FNgn6F0eu40VewP
Sbs4LPPTEJk05WqsaohUw/302G0qasAQb+2/DaOAvd5youqDqMPYIvu+w1DScG6PS+m+ZpG2Fpkn
ESVkl52Fot5VS/XQxBQEJevQiATValsB873cmjryTkfXZ6lTB6av87I8bYY8s/HGDLUwFeyvVILD
BHA20/KM2uhC1DEFhH7VDIF+n/F1rWUQSeEL2S1VXdczfKKUoS2I9mXlSUz14uUE5gUPbHE/sSnK
pGjokAqoxzZyQ/TVt5vFhLd5laCGApxjhFb+iympLVSWYGKpsC0+QlnFwQGHBTZAsIrYp4L1OHqe
Hmx0CthLtEANwYEm7w7KxkzC9KmhoD2DJR0P1n8Y077MDclvMZRnLBszShOxgRqI+fDnzZmibxo6
VUeLiCaWJBgcnItMiJ9Oa3bSWYQfODkpkg0GOOOE/7h9eTicIzoFzFsyt2Qrx/4jGmUOT1SBGI65
GST7FUMhWieHs0bYb6hjx7dWy/uBIy2fUs/PTNmj22mUIGQ6tSyzKfo+Qx9rRXR29RSEwL6RL7Ah
2NzTslnIIzqYVsCyulXmhX5895wO+YRoCpypPVzK+JUb0+MySyTpjASlO+EKGGv5iG51hr0QBynh
TQWT8OxTyXzpFi77EetlPpj5cza3kFxRI1v0hFuq9IflXV5sWBgM0dkfs5vF430VNuSSz0qMdvDU
sPdOjhGN41mj7vqSnu8DxqE1ggRMaJO0ZjTdwp6Ow15ZHtKSUl4Q6t/WoWKSz/84RJsh6n2k2Y+v
d8J6hxD7F7TwWxEsD6jtJQ1rCd+XYiuEHfLTag9KgdYJJECMWsxwWU1FE6cHvpOzUs0OwpXwbsU3
fpKf0MXE4YwJUoK9RIudSII55DLFbwxbjue34LweqqVR2dyPM7a50WjO61k52n1bPVYT8b9WAME7
bG9p8uPen+gVGFQbaxsnHM7/XjCEoPEZVjrMa2MK4aSTI51YbuxOdj0i/fxutUw417zelmVOsJp2
a9PQFhwtcWCKLihXzBU5XEUh/M4TH4/0KnjnjpqSXpN3FFJUDgQlOUy1LpSRdvarY7ZdGxFwB0HS
7p8pE+ANs1A3xyqhxEvXnpipI70ChlWlYTDkOVt2rAmEKAXUrxAUl7EDh3L9Z5k+Md5I30hQvsyW
xxvK60FHB4fC53YrSrPfARNXNFq6MDxmgL0JDDNVpDD7Q/oMDezm7xpcsCrWYsBitHhmHtIvEeON
4wwFcdir5jeenJCj8WVcmzioH08A9Dh5oReEvZxSOQPKGQcFIMPOv8pFiAdmxN+TlHPtlxuhNYtG
DTYI14lEQLjqbwQgkMOX23Pho1OiIvxM6FHAiig0cNx9t6Ef1jl+0zX4uiuup12NfXWYxkuigM2R
lnPcXkZf253kAbuhirotGZpV6+RlmTGiplLnqIoNzVHik/C1gEUbdTCahfms1PoSwLIv0tEc1Mje
IR5cRoPjTpN+uP+xDl/XFGySR5iIzI4R3XO32mAJK5OEZ7y10/9bzwCGwDnIPI4hTp612e/CiEHm
IvYdkV+8AVVFmMrXFJZOucLyAIkNlI93pXoChTWuXbZOQcXrJr2yW73R9W+eLaLPbhTzAH8netxV
UlshOKB5kFgRxXFb+Ce5Azt3JkKZ9O5hFJ168gf4UpSveTE4bNCAJKbaLjxXIaDTOCaZ8CK81ekX
m6+cC623c5aBMbjttydfJ3GTPmhWwxowqAvKXfcVj24fFXTv5WMM1pLa6/bYmzneYaqClm90ajwn
EeIbfihn//NMipngkANVqPWwkI6AEm/F5+KGES4MQTDlI6zPMxlgzhJ/pmOYlIJ6ZYZ6KxwUlRSC
ByFwksDXS4aKgTbKJYrfWoWvmrZkeFJyfIbVhHjJjICtOaprQPD27Yhutx6t5n3ehOaVkxZvV50N
4ZdFirkleA2iKUqdbcBY0lywVsaxg+E22t4/ysBo3szvGx0mMGRpiNgXaGGrFYfC4wnUzAI268V2
enNiKNSmu47CQyB/0Uy7t5hdvZppyeKN4bEDdRgAkRJCAghGGT/4efTQUaWZA7W0mmnOwGWxfWIw
n2FdOggm2ttgTt2GN68GhjPiCTBD0OPYqIpB22Dhx+yPIQD5Ax4W7oBbmPorJaH7WJIJzbM23jUf
jgqxp0LhSoibf+Z7rhKM/PkXOREith4hkUoTSILIdqGAujoC6E0adUBfXrG1yptucARc/EO58otf
1ENDfXzGnXpTa8+k38Ij1gTbX4q4SDjXqNPTTtMq+5ieQ+vYhTn7NEjiT0gLdxVCvEYsDgwP7EFp
BkoylGmfOcbEDygOr5kuiNnTM6Rfha4wgrSUpGabxl8mwQVRG+a6lNwoCWAOgBAh1ki2aZqgZl0o
9SVbjmdKRia2uxM4NbVq9hRZ7E79qBC6I0COTLEcJuwNOSHn8kWCjiQcTBw03pGn2/g8F102djwF
hqi74o4dPm6VPpaPgtPx2xKgkJwIdIp9u3Jg2/2RgKKoSH6ceHosg1pTJA+7SnukzPblsFKK8mh2
PyLFQ4LIrbFQwplQkCs7MVYv6cKU24haS6FSqqWSvHKVAPuAdH9lK/eyMXoy8XoXCiBQPsDMvSld
FUUAytw8hJqwwI2bOmtRMJ63ZFs6RdKV/ZVYPMDO192Z8P86AJzG76Y/B3u9/ZHEKp8ai9pnSzqn
1do1KVUj9swUfdT1aJrBl9W9QoGRloPtel0tHxhTRASDLvdsT1QrV9KxmAPCtdrInI51tbbtDp0u
B9Y39GQvOGLJMZtbUa/v9Gcxvq4C0Be+y0rHSwHx1vF269TSh/jkk2wxHbOMK9y7avqfMWoHrRPH
fHwE80vR91SzmLnvgzNqiD+SFhvTLt+wC7yRpuMl8ctqror4LTOw/HFiTcq84wROnPOVUhv1GOO9
qjeJbb+yngA2O9LjZTnVI829/Ox5arA5oPifgeu1rugyCYZxvW1YUCvVA4l9IhFnqb2qCvXTOPP+
U9l1FzTu+HxmD0buUdALUrD6elSPjyLk/pWFCvzV7Kw8UqptdOmNKO026z8RqUuQZBNzgSOs1iHZ
OwHf8jv4CFAmueosPBmrKQg8gvflCg87hvOc0BAq8Bq/39y8hsh7ANYXklhuRskI5s05IBz4HPpo
F0PXcwETO4YTXt0Gu7AA2ITqrosfVz9qL8uk1+WayrNdUUlGRIvGUK+jlT8ZNqMfyaRDJzB3K2Jj
0+/hlCTb2KKwglhzuhDnEWRjp+s1Qn70bfsDRoPA3k+DvrAI+5WvGmJ17Z2OvDTkD1lu9SqbCBy5
CXlc5PmIsw9X9uz+Pj18wo1xeQXGRB06Dbk3YLEFSolkqfiKHJja3+w/Luh+dNJswsaZOY006cL/
Jgs2Cdv5IOkd4YeAhRr2ewb3I2Z6Rti86mAiynQ4rbORd6zv8JCy2zPXqxS3MExp4twwsVTwhgqE
Ty+xVgrmP/xTDuToxQ8RQEPtxO1THG2X8ocKa+vf4mSVpZ5pI9a7GDQUlA2WobYUABYPFRi7/NTJ
Lj+4pbq8G/PmrY9VgGeMiLx7dYjsEoMPVRYJD3/Ji+63dZyep38jy1Dqf5Or1g8Eb3b8+UY0u6I/
FxMPn0IibYYuANFKmaGrZ4RQ6AalvQG0P8efP+Kqcg7WHYB3BK6RUskO4b7HnLRlK3Siwapwi2KG
j/A/HEPyerySBFKwZlNpzpMAyKKSG76PcG2SVt8yK/tWQNN9T26/rF50JWa24Im1UID74FTQtST0
609Iz4Iz2J9blsuMy3jV3c/E60ZVpBsBWks0XD04fAjV4FJCV04taFNk+B2MsW3Yph+Dq6HcSODC
ZtcmaMPH5OcXR9qwvAdXo/xpScpecazDgJqk/h2R1mLDFQ57tRg1xnFEG2piMdRscY+UCJ+szjKQ
s67cXHdnonOD39H12hyWdz68A7HJPpEixIw+7d97DLHBUdo/xXZP/x7u1OX+zoQ2bwTRTceyVj9l
EhRUkKuPMFVMV2X5eYs0o8OwOSuxYK3Ekm/twieukxhM//r64mRSE5xnZyGh7w27lrSudKR2F77v
bYkNgw1rb50mBwGlVXmwAFmfW/vQtv3qKXPCcaylUe7dP6y+V9B5m6GymjTVz+dnnF2a+r1Ym7p2
ZRZ9p2XrsBLJCFVUiRLllvomyDStEoS0moN2BPNllMh8zjZgyM9P/56rcZYA50UyBb553B5vf9Zk
glNdz/7CW/dpQb3UJUDWa/u6KmbG0uBeozV+10PT0vm2NsORoFzmdWh7U1CH5BLdDRWeWVCKsHU0
AcJtLK71DDYHJ8FlBIYngNuripQyzpGvCrn4//cdAj6bY3CSwRP5JkzDNRFaXAtP6dK48WPD1cDZ
/rl/fHyl7YrZo8LDRh5wZHdqmYMmWzdX9slXCaq4+k4njSQuPyA8UeMPOTJ9dicD4hvUF9+mtp7W
1Lfbd6vgKTSl/2T2WXTFybpA9e6aY8NgFRvXV0G5kn2mm3A8zSY7lp/ouU+mZ+5GadkvwMMXBypv
/GC6fCi39qEPz//kmEBg4oK8A879GLBqyhMW+i7hgVcg96Uu6gvFBsZC9frjk4w0Z/i6/U20gFbC
YNoBT2j0nRJOqq0cB5PkG0y/Fo/TIdlYQQtI4V01t0Ji0d9ugdPl17gY6EGjSFDgE7pTJer68CnZ
1iFvR0bUWDSWZVvw8cD2qmiDgFPgaY2XdrXGFJ4TD/oOv5qDTffte7uaR5sj6SlhWVxNzOM0kyAf
z/CDiITtuWZGsU5Uc1xOgPImtCfsVfIA3Fcm0un02TcFPERzFVb6LjoFl4iJYkdMrnGhp615MRO8
GMhxW3cXvpzeTXr32q+gXiMzKiWUAdw2TRnBh+y3GvDbYLQh7ME4fUR/b2zBzRzAqVJtTXe6jfyc
fPEkVfwSKcZ4nhQxbY7L1dnTFRM4wAlQDxC6tiYrY62tVqwP2vIRcA/Gpxdug2ZJkBrhEW3E/Z3n
LVb84FKX0o5EzTTJ4sLefhPZVE0Jlzm6qYqr56PFXfZN7+1CbPTFV8p4Tg5MScaQQT5m5XALkDlx
gTKr6dniMknjyTU2V7PNthxkiZ585mLwoYqWs0/Eyu8V1D1wKyZmGUHtLjA/pLyQijwT8egA2/5h
qGYLyDoWd0PWuszZpBexH+cI2RKrdTD3zkf1dWAZFsJa7KKHyO0yjk3W07UVVMYr1qFpx5OcXCE/
iFRovcH501xvgtf6qaqvXOjUASjiu53tOZUwHpWapy6gSHKNYM+QFzUVRwIxcjjl+DhgoU6SH426
NUUXpCyFgsGfaJwtlcr9LbqZwEo4hlOfZcCecV9zA0V8Trbjv6ldGSyAKC9yAQNTz+KAonGPxqPq
VlKl68t1PlBBquoKWQx3qmMzT/nXv7QJo592oGfV7r0YaSvsj7lGCimXyn4i9NAZLgVPNcYCX0Yc
X8frwjMJxIktl5h+9d1HSJ+bmJnxiBg4Hfjn0MN/5XPEdTO2aBvzMiy+wYMlZGkt9FxFCAiT5lEU
H9nKeVU0gtHO6uU1SPct3T2khDghEHrNSmN/XjqVk3ESPewFNswKN03vG8eeIjPSJhUZcfv+I2D0
JpjYE6LWj40som1R+gqNbBixI3zTjhYifB8rfAkmJhZoIxFvoRFztuiF3QZEF5TLqlyzbIcE0kSd
d1z0aYT9Lr+FqSPH0noHpmeeepy4ZCIEpzxgPNL39RZKwSIlgIO3qLc4OtwQd19nKpaDvMHV3ez4
zxTUx27KD72UHj1WrSSbpm8oIYo8lacp4qVT2RbgIYX0r9SLssXFo0EWSVOuLMTztghLVi4QdsuY
n2bpJnfoBx+aObOpPmr6AvWyWArGqmpFxUvN5t91KjD5oxBEg7zaLXbJsf1GbryjoZOKndVM6E+E
Dglm2LTyUzaAO0om3ZB+l9IpTc91OBLyGip72VjhDT7b0ZE3nYQ3vH9MBh1T6AjX09k/l3oIayol
WKh2LVoUylyD6wJM7+3BOcxQ/wGDe0cU3OQ4yhKRXLNz/rpIm0UWQ4xIex32JURWhnyel6B3e55L
gEmgDQIm/D/7iPXbFNz+r55RJdSsHvfEHSaDjFIsdiq2l7OBNBhmXarIrJDRAjYOAhf6P/236WgC
W057VenvDu5R3lqa0eb0jquNl6MuzLK/Y6//dx7B7X1QaU/73Il7BZlH860+NA0Bf2UMjx1SjOI+
hhu8aXBxuu+B38USAVApdR4EuPSpCbEw38n+ckyvVFEswPJOvbkmErUDzmMw3AXAR67RUzAaXqji
+xqO5NcSqsjBVWfAf59FxjTZ4QdpLRKPRx1B48HxTYEmj8csaSyYN08oWPHmycF9BHi++kXB+ssQ
kKVJ2KwsKhY5U5jacG7+7rg9oC4K76HBZGJDqsOqXEwsTnLIH3kZrxsGRwYreMkRHvwFZDumx9X9
HM7H/ZpP/tM0t7aeX4hUuDuavMv663huqIC1wzf3+8BjJwP8+JTPTLiaupCQ5p+7XXkZ5+YtFyIk
FqhJOBJLeSa5Q1n9lciBQUFwqZcATXbcCSIMQHVDa6Hw/zGZd4Mxd1TnAiuxeVUlCMFp+UyG8f+o
6vgsGWTZ98+ZNFaOZ2hzGXDwCLgZ77LK/LtJ2+yzN7oQh67qIlllKTk4rGp/Tq8G/DV9ACntO5V1
h0Dy4aDuOQqJqJhPfpKjH1MESBGYU1tvZefiVQszCd8HZH3sZIDFpKfGIcL7BJ+UmFm5VMzPEPzq
B2wzPaMcyNzFqZC/2N7T5vODPmWRmLw/SuGZ9B30qmoqrpuZggn7G82E5OKKkxNRr1p5jl9GX3OK
lDsETmv+fEv+a5lzsYcnUUTZED3yFM8kbOQuv/HMmwXuXdANTPtZLtV4WC4YAp0teMsr78TDGHAy
xsaIAAYxh0CFP5RYWWPJVq/T40j4PXW91PvjrgU8twXBp3FdU1ojy7KymhmdEi5AIEryVO1HjJlu
MB5YpZt5Fx7N1vqWNQ77k5aMGHDOGPdX3LDeQpw1yqLs/ceEswYEvNLu5njK+J+Do21Pc3628xSK
HlPQhHA0Ypg7FkfX74ORiNHvqPssxCRdEj9v+l9bdaA3yy6/a+p6mZ46wTQjz+NwxOjDCIJMIDrE
iSYy+lqRyDxO592wR1HbRj7Gf1CaOGB3RATarmcEBcd0O3NYF2vtZoQ8cY6Cp+KUHyVPwjUERxp7
5l0Ats/VsuxPaUAqJggXNfmXJP7kt98Wq01+gllhXcWKWSQFo+eVfheHI39PQHRVmHRaGPPpBgtN
vvv4Bp1igZAApCgTGw3BLPqbx0ScRva5V0xO3ci39EYCj8ZFUB+ji3PrtPM6Xtw2/hEm7VP1yexT
nnZoka5HTdAObUzWX2ZbN5o5lKTr++xmh0DNNj9h7tYJobFL8usrMaywA49QvzXHtFjzn9WQcFhn
HW6Y3TCzl0Zq2TIruE42IR9lonv5CZ1D/RwQb7ENH/Rjhqt0jgsBGiGUFQaA4fyxCGLP0NfpWARH
XuYPp4x98F2LTIBKJoLX96fupKweodHm+0OWtnMM5G3pWZUsHoXtdeSYXzR0Z3rA96XTU8oDW7/7
5VOxhch0R9edOpiqrGVD2M3QbPG35J4U8dwt2x4NubSdK4YULpIJckZWu1Tz5TgvEta7j5ktQ+l6
UBmZgzbr2IIVARyr4WE22aBylAkDBjpHsUO3kejUqdZlY5DQ1YaAGSnO3DOn+igRtW77KWX9Dk6J
bcA5fAkf212o92npku3Dxe297k0xtntw5r/z693iD21tsbO5RMNbq7e2UvtZeTe9CyRx5euPleYh
RdBn+7osJNzDfb52g7eDu3x0O2aug1KcAdYwnq3pMDKKPubmnRGySxUCFOb2s4SmY/1X68JWxgT7
XOfbNKZNk/AUmIZErfKzYPrEUW1ofQ8grSjDK/GIRB9VBG7enlXve1ePGJJ57k0q1t3ykDOrXm6p
tuZ3AFUJmzB3CRcYTPMcbz568E1Q9uDba4lU3tvbrlqV6RRITbXEQlrPr8qJYEJlS59EBktYPjEJ
I9+CHoeDbnTjgA8llJZhNmsXR0mDfyrJscLHAPo9mvo5gYYV9U4cldxCxHjnaYslFcmZXTDDPPW5
16IZdFsZlpISzb+u6KXwrb3WXNklC7OJfsHwVZhrOuCbXQlvtcaaZL7GjQ3t4+Oio/CTo+RdQ1iP
TyQJlqgmYC3Ddi6EzLWQx1eyn+7o4Pw30NIZfSv1OWB7H/TXwIfu26RBQp2RfLA4Hw6e649PbzO5
YHFiT9pQot2CCY+kOFyZPo/Fra65k++xcyc/L/cJQbU3Q8Ck4RV+4WAJnW9o6AfvosFK2FSv8H5j
wLfuAncVqVA/ofXZZU6Kv9yPUByhrHb3KRt6A524XsSasqk+2l3DqyiDitqpdH9bzU+VHMfxGbTT
cuLakdUgYwVQXWjvl5vDS/h8VEA/B0qD5IwLsoHTxXC2hC+ooeGbkqPjwsQYY81MKTYPI/N495TP
LcHJp4Ymb5D+DpmSozF42hTo0fX40aZj/Ly98K7Nhq77fxMTGqhf6VEs2jN/k2ezM0HUEZAt3HYO
oDlKC464vSk2ojc8/uGeb8nHsUiiSFRWI4HKTiLAxxh56bm28dNcVzu107JluRSCdOh4S+geT4/U
U/aZUj+VHaRUJctGlRjUjKJ6Bey+9KWQ2oihrDelUqrLd9I2yeiiOPhy95dKRqpzVtbh1ZzIjig4
Zpb9zE5JmFaJrxq+vp2ciiXyaOlPN+RoiK4IXVr5Wiz/hiV/HjGk3LSCvGCwQ3MzWmoMLTbp/KcO
sLufU9JcFiEktIM5M7LrxevyvN3ZqmFt+34jElfaLcVesTt5WLNLCos+f+14iljUMui1MQe6Rh8C
TKhKja2tEFmGdfefucCxq7PHQ4OAc3narl9rLkrZl+5oAJziy6yGusHRfBssWKRl5qhv5yc5WS8b
/BiazDVCDn9I/a0himeh61PiBJ88cYQoY21Ah5PYqlUFBALSTFKBI4mUBTrnWkStCQmd7oaPiHX+
qsnaBoRed9Ks7w0S1EXiCkrE34PGccdEX4gNeyQjfSUuuSsLc2Npgduv5t0cZncJflbKh9ZCM0rO
CzjEDb8N57FQMPXevYohKSZHt0jZWJstn9Qj6krcC0T9pAxu42HLRfL01PuJXjWt9l2VwgfqbYqw
RZcAzJrPV8+0zbImLOTVgGbgl8o6G421LUtAETbIJjgC5e5ECQaDr6ZsJ508iKpOTCR6FO8P2tIA
KLdjhQVPP7yml5fcJjUyDuXhEp0WmeaDklY5aJoiLY1vM9dKSmV2VxqyiYuf0CyemnamhWVHIYAt
nwTYv2T9NEAqMbmlG5/oGjZtGA1t4k9DCFFzVlfZ5Ns5ZA5vLPLKqfvN6l5wyv73NOSxMPAAEvSS
Wd17w1yqFBRbXoLYaEYsRpIYW0YuIxCysPHtd/psvmTov+Kk71zeGxQy33u9CI9H3gbGycUr7suF
EqPCuNErBOzddBFkbYm1IoFixdOgQ3v5SQ7+kFYszHtyE0vZbpfz3m4zTMXsDKABg2XJljF3gsl6
6Y1YTicpRw3j5o0sfCedO9pcvVSWQh94ZQ+wyU0i6n+A9kg+2IEepXic8GkpZBL+fH422H4u8/rt
fza2cQNAgGFMl0cJCnDTOvcbcS1VRYMB7MF2YlV/7KRbf7hoBCFPGMhmWDIC1ZeJBUpMBNUYfD9n
8Bcd8WMs0vHpZKmc5g25OAwT+EoFL8FUkAAoZeTM091u8klttjRoqz2nwVhgsh2YWuKFCa4GZ7sz
5cpBFk3m6/C2mszkB9hECRDrUqQZzzB56B8bTMDnuFaE0bwNXjGl30XAVQVRAO1v34MLVLfdW2PZ
loAPtHNzrAdXze3H8Xu3FI5viDkQ4zSrbPEOKjm0OitmtLfGEwpVcP1zPvhTt+Ij4953XA0b8ICx
8Gba4LTTfrVO+ZAezrmkkOOEj4yWjsq/AtFO0gaplm8nt9AkzzsDsSsVALB6mJqehPOOeNb5WxrI
CSoANlU5G3VNdhU31Cby9XN2Y1aiIUPuppuCXSHBZUSYyi7fndiDz7lzO5cn994fRmw7XUBzS3Rj
sdMinK8PevqjOlJzcIurQpqn2l7mYWiiYqYq1yuWvsCL1ir5zWAlWBZ6Sfv+vwXfw+2i1ceQaXYI
JOJk7nBbYfX8+0xCoX1jEFc1iQB2yRljJtnj2lxuuzyWCbn+FaM2UsK2sDzRWBAi2bJ02lw3StIm
6/ijoU7CqUOOZoUGAPOior0QaO4jEfPiCNRebPlgQhzJSHtqwMRJW6fDG6OPCmVzOaObmFz7wYmV
23al1PfJIVVOiUD1n+Gw8of4rbDiYwTZHkKD5oKVhFN0KhzYTK8nqkJS/JQ2ZtvQ4KnVfcx7RZWz
tHaIS1SBtpZ9/2+TvQMG+u2/8K7aFWPAvr8JMxbvKc3vihojtXcH1XgVf8GiRDbM0TWgBtVD7KDq
wwHrPRaVKQ75yQDZ0NJRelC0kgzfO8uNlHRxmxpOwkoZxGf7FzY+Q7qEmqsXCGoSO8rfiGsdkR9x
adWvclZG2iYNKjUrKZTRfsbIRJ/W7OdLn+TH046Ho494+ZuTLYtx4xCE+7+S9BYi6GdcPpD0NKjw
TYDvvjGO6wAanQ+GL9NrzdZOQZXbwuxRpBPd34ZycHtG4M2l5dRtLFJWMw064FNHj9P/CERvhQgT
OO8kTtg9ClD5qnTF+J+GTrjJbZ1LWperPmWYV+JQiy/2d+2dr2T0z6UnuwO6p45d/VZNJ+LKxXSI
FW1g8rCAsYVDfW4g/47ByHeMG5p1pQZRjLqhnDqmTfQh2sjMjJY+HzWlnOj1apgkaH4GWNoZ01z3
qGgCBUGS/PwRHM9yBJjK5cfQjkYCeqJYWRPmJKWctWc8YJQooZB0SHljVaRwx7UgwyIhezS3fqLS
jJIWR10OGqde8q+R33Vjd/Ka4xeu0YHHocUcXcuGhIitscZY9sbDfosdW/mYIeEsQaykXKgRlYRA
UESlb6CIYcH/075ioBj7eAVGZUrLTjjRfS94xuAyJiMjyL3u7wzRz0wnUKSRgfb5ixiVQGcZMpch
A+KUZ46gD0dhs4E5zU+7A3x90jSw2nJy6X7yHfzwIyaDlzlhs/uX9+vU7El/HYRb8vkpLTYMLIHZ
No+BTAdF6EcM5Xsau2erSj8tRAufN/UQ6AOvJdSpueWka8dw1jpduLouJOXOuRiKxnWmZv9WGWPs
BcWu+30rUaPI+j+BM1Qv9gF9UtkE545lGQQKDQW+S0Xwd+94rPHU5CYcWrgidZUQJMyDdAwcBWaY
ztV5xasZj8zXoyGsQBZpBHCW+/2kAI4PxgLjN8DZQkDJqFpHm5OAsvHEjdRg5hJchAV0ZC+32bCy
YfCADOfX7Xaxp4ap7ZAOcliBaFCygvFSvrK1RweG7Ap58+YSoOMX1mSFLjc7Q8vBfBbaNmi/H1BU
1vLb3ECCzpurQK8r36ePPkgtENTguBniJlFJsLV7ki/KDF8sDZimgRLQqghjOD43DbgR+A4yfIYv
u/yp94abZ8M4s3zaASpmB3m4ISCrE2SzVeC6r26SRI83B7YDvbitOtaTnIN349bqPcCgjTm9zsTo
cV9f2CaL64vYrDc18DtDkZPbptxEaKjoPSNODa0W4svWvrCnuLoz4Lp1syO6FrztsFrR0OyozDao
AvJUHYvYiXP4gQMKA4fvkrFPX7Hb7u9agBIMRR8d40cGVFNF94AT4ho9MSb6q9clx7Y1CEb3lxqt
eAPzY3COJXJjEEKU76feLD05ac0FPb6F6z/ZS2pXAFe4efN/pKoxvN0o9MgQLMy3cGrh6X2LMRT6
+5A+iBxfwQsYylfikPm1aYzwETOJmWQkdMtyip4U5Ddsc04Z0++GT8ZpNSNYSOo26oecluAtpr7R
dqkgJPNCtdYLB2zjBuLfb4yS5O/K3PEh1SrDwbF66+/rZPuQQll14eFQmkG0+D0svwaUBs1cidKz
ummb7d6QLh6R7OwiAD22r+0bP/Xz2oBuBm2FZ2PiJppI3U7d3KuQcyPXCu5zOnM3dwzO0J1JSPQs
lXGAtodmXgXPy5AbTZXyEuEte6PGavhdcY+0I/i77nb3KDbi45eGbW9eu9XxU3UAhcIGcqbGpl1V
/XjIYbeB6l5gIdrv3thSeU6aB1evTROvU4InjZ4sW1Ek1xO4bOdRfwgnRQmjQZTrohA5vdxVW32g
1Xed0AshR8omgZEHcZeUfpdbrL+B7FAWn7v08nMLuOoxDFSDKf42+yHjfx0LvuLYAdc/MszKQpZN
IzSNRDSTy5g7E1GSsuC9cJPVK8SRQ8XBUnZ4pyz6igRxgbyp9GGp52NNOPiNdw+IQ8dvoYkemcAy
Tc4fe3RmPBSdo6OM0tBHVrGl25S8d1+d+9jdtPeddTdW9Apbt8xM4AsnkA/M2+64bHrehqKtd9JW
GUH24npHej9OkGa8QFqbIrhUTQbqLDxIKYfPAYHdlgHukyHGxAG7+F18hnbIZeOaq2reYTqmSdUk
AEWPLiq/Y+DL8czQx/bk99gXgq1OG+sONGxuIPva63CT9/1awkrIS4a1ZiJeoBJgffcjFkH60n+w
9dKjV7hgjJfq87vqIOlyUu5RPL6Mv9Bw4hm3FqEL/qT7G4njonEqpmbIEfLivqQqtO0mU0UY30EW
FPI5oAzXfJ5Fi+JObpyHiGTOI6vhMAfNS5ZjlEGRr5l4ZoUQOFyd7/hpkhIkdwKtxx90XJHo1NZi
9XrLTP+gTlAzbarTexSP3rgFzfy/L/T+J47juWN28aIQ+sKxdHDnytyng4eKmNS+6wOdK5R/UtRf
ahLtk04NHcCtAlK97pBiVxa7yLh1/bsbdWyO5OSqO2vT3jraceukRSYqWFy62vkynk3X4n5kbkjT
tEi3UgT75+J9mGvtgM7zz0q2PexYWK98xLFawhMAqZrcqiQDY0WfgA9rRsMpJgFb9zSQPBpCKpLv
iQqSpIi3VLANn3Bk1gEY/hldVng1Hy2/Qlv1+MIpZgiuW3IrGKJUMCXAW/+bAO2peLt9qKefWnCK
dz0tr8i4NEmHKvDMNv7w955xVanSpbO0bVjhw4ymnSsoAmwN1OEBAz4qugS7z1b2+h7hQxO8/J1w
BHHyCOMfhlWxt00MissyMPW6qkAoblQgEe79rQmsXCYsX2SoXLQMJqsIy4YnI66t3YCD2iKqBZuJ
sLLhJNBCSTgwji0j1PV3WDqTa2TMgmtGHIAWU4DspHldVPnRAQ48KLASd5RvyZ/9cY10Cp1wgnBS
LjVrIv91HKRBWCZnaMo7PazUW2rtqT9dFOJp8z1gBmAHdb1YQYXq2Uh3dlg+dipmnGBntr1Q7GSy
dMsDLmCRfjKmZKePKVaAHDj/y89zHABfWrNuAPnjZY5at7couvOi9DLr9m4EGvcmm4T1ufnd0/Ro
NROs+WvnfdLe/dIRyXam2lzAz8VhKFnxMmQBFYGYYY8nB96mVRBXj2a+vjq7H9QN74h6XSFlAEeg
TrDIPp6uwI6DhXdLMrSiFYduS+Bom3cHIjxbRFO0CtkuLgpIeW2iyp6KiSuezrblPoY+mCfXmRyZ
RRiN5k9FbSCneWSA6iUHD7Xfrdn1K/CB2moi+UmzJhVZ9Dumv6T9Rut2ciNmgulaicGP2TTg2l03
1PGfOHmyAMF/6f9XE+xyjFgUK9GvlKpgqtLXEZR+pXnAEdi/0EXM5iZppwzbyXeHGQD3cBSna3pR
fX9KFNZt6KfQa1IH3l9XAk8ti7lxRNy58ptVx5LGgJlMzTCYJzAPj1GsQntkIFDKRpAux/QNQQ7w
qESmQ3N2l+bbg1/WFbCffYKay7C3aswaUMR0pGtgXM4enlAAfTRWu/hnkgRj9kCqoePG4pOaVSSJ
gO3PjcgLqOfhDJyms+nBpK80i57Ty3hV4s48vqQZ8rHdO/3hniT6baVc8iEVRYPiIv9+VH5B6glt
KAnaLGAy7VEVL4dXa0Hntr7Fm+rg3B0ePuUnsHm5gF6g7G+ifNRMB54UTsHW3EaccB4RF+AZglFx
VAbZ8wgWBwpRKYy6vARAcnyd1qPuUctZL+rJ+AzqdNgMHNQ1pxpYmCI6677JtYA3/zUoYu6bJxTm
aDl72kkSaCbWcrKlh7xCjpUyOrbpYYcUhWQjQczmNWS0iKrJvX3s+0GnkKNhBUrzXOybmmcKebsu
DMFsvU4pihe6bmIZb/bDTEFnaUIns1RKobdWQBb6WGejCnnEq7FwEEaM44aX2IkPj3ziZPnrEuj5
1biJEC12oadBXJkcSA3CyjhAfhr6zCraOdw16cZXw3Ts6v5QRDv2O5A4StDS5KXrxNlQybaDetiH
uLHvaVKvnok1g036NsUeg68hQ10PxKyBVd0ccnPyjs62QlSob4M7TkGLdgKdRRIyxaChoGuwS2Bs
Sxbp+514PpryF+telOb1F1cKnJbjLWnyRFkfdgPPEOPUIig08ezzOfSHDM5Lrbker8cwzQirdbMN
oeI+Z5pWHhxQFZgFaiSxyV9hGQyoTsL/+FzI0l8t63UmDWOFohk1B1WxW3533JQuQHQ5jyKpbr4T
3QKiCcKUz2AYifRUL3gL7ToHu2puDtA2c6v5Is77rfcizc0lgG3oTKXIY8YO1Vk3ZrQ0gMRIGftb
e6IJYn38JKRImQUbS3JdA3ajydx6AhyEOo44iLLakT4dBMBDIuA5G4A+eZGpuoIMNPHXI+PFAwBe
VKguiDiaTM148OMf0XZV2jNp1q28fh9z6AhtrDVHU0N20UU+BhvKWtib2mqNelq85S5W1bAv7UjD
5mkdvcvaoNICBly7nD5YXpvFXWDcBcs4yRUlyrJolB1QxSId2rxpyhMPq6/2h71TKcj6HRIKibWj
oRd/QpiIxP67063BTsXWG7Odgc8JcKsl95aRTd5XBz27V0u93DDITyVpA/o8ql2PrSY3xgjuMEOa
faDlEeNfsoP5/SkKsZ4uUzFXs+SZ8Uhr2/yjzZyCq9edkr5Wq/dG1MIGSIFS9vZLPhZ9FW+7gHJa
kB2dnasVfQD3h9+BNFVpOHlx2GA509aEVdhaG8Tl9qVANSY+OSKSCuyrYDc97eAC+mpuxrh7gPsN
SRd+7wS9DVmVIla3P23iUsZqZWuwXAu/HvLbm8wwmmFQWOTL7EOQB3+99xEjv9JWIjTc5Wo+CP9J
DHT8M4C5e261FZe6P5XBsGIypRaH+nl6LtH3SbdbzMGW36VcnXEkJ45wLkovsRak44wwgz0YBPQk
ZkJ2WO6pfDzttMU5gddofJ6K4ZCVbLQUcS1pNb5aig0ZoMPlb9fuNBk0yxkdorVlUaGSOOyNebFM
+Mf/j8nyd3iGz+WqyTm9ryLwfR0XNYfXvXdjP3lPBqEM4eQ5aTMi4BOubSnzXdGg52bv5DThp+OE
uCC+I8DIwWVLJn62Yfr0QStbWvHtW+/VGCHG0J3c1AaZeSiUdv0TUi9Tep85XXinequ/sW2a7iJC
YJV7GYF0Va6OCdwOMI3FFZs9uCERBqQMDY98nptPemgOw89fHRZqihGSGnUdYSmGC1yRHWcOA33e
sO96EuJu42bBLA+Jbu49v1WICN6e0w5g7PEdE94qRZ/KypMkLEVS6sNqmzEep1gJ+NiXkJlidUxq
Tpcg4g2+kzcq1lgOIax4Sk0rHaPUNQh8GjPPfN9aiX764F4Yv0VcafOVoZdv3eNERpQgSZEAeIuK
L1Hw+c9HoclbC3ftXhqgkmhBWUuH7c+QSxR9MBYR4x1u82IpBlt0TVhY0bLovHuF89mK1soaZY4k
+wZ9HbN60CsjCWkklJD9vdRgAyLzWvBWZ3T3noC4wJpuIQmOLVVo788FAyjJtzaHJA6QbiFyGmcb
1uRoaEfRZhgvLsEVA2Etnj6GjavNdhfL1zlkezmdhAWdU1RAEWJ6SMIcavyySU/YusOUxMrMDBUB
6Nahzt40D43WzPh9hum1ffG6pA6ssFAMfGyRgIa28N+EPBY5WkEzCo4fSuQDT0u7o4Ckyj/+1+KO
f5+e8ddvVi2IQZjP3yOnDuJ6VOQCAP9HrmsKL6tljYRfV2xGpggO45m6xF5qNiX0I8xzPGHUZDF1
pA/7I3LZDEOfNgXY1NNV25TkaDkTeh5dCYMvkvPThQddfjCgSdQdx9qGXXDr1Fo+lWhlBdgF1F0x
nJWTUEMV2PmuU52xB/lmzbH57WZgiA0LsLkagdUlLDaHAkOgL5gXkB7OiAy5mils43P3SI+gh3AN
604zatlPEmr2R4xypH4rDszYJdNWSUdu48gdjyoeGx9zbMpANqWAgdHdmu8t+MB+Ia2kQ14TuUXs
1bLNXaaMod8K8w1n05ABxnP90Rx//eu+aBALlwkafIhMbdhFZleHL/OlyRFBQRUjMImhDXQRIXw/
l6MP6AudtOcPkUFJEncCLCDETPm2gvkWUV/fuwrGUSqlAG+7qLHqdEWM3JtECLqvID/T8NyoMW7d
Ce8KjgnLCp50XuITVu3tLmKGvFMK9QsyLxMGKZXADUwTs0fOPms1ntJC06BuyLnBTGOzAtCytsF5
B+Vc5suJ5sM9qjjpIBtfYSKXsU9FDU1k/WrYzNOOOAI4EAny/Vp3XDhYOwR0bFRRJqNJ6cMPPDZw
e2Gz7XtGZZDwIWnRzTjrdjg/9A6bneHSEpPhOEGZS//YsbEXDCraLh+3ricrwjCjS9bjVnCSABcE
PSTT9uxoTEzqTZ5AjdRGH9GzvNn6p39e8kgme6lRhQlvNsNvLR2meCLqcuWXRRUZZ9dIDLKDyrwe
1cZ9BW+HMpROgX+Sw1giLER1677jBMEpKDagWA/UAJspHWSZX6sWle5eAng26jkwl1+WR8JCbQRp
7nC/BojKw3liDEzupGO7BsRYzxxshU23hU2H7miaCrlie1tc8VJ/opWrr2OfwHikE+xx8/tj+XzN
Yplcj7MZkE2C4r42AYfeIxbWjW6JfG10E7H5boE4zGD6qlDRPogmGW8elxFKWqs6lm5226coiBip
BnAjswz6cnb/3MXoFnpFqleDnJUcQnSf6Rt0qrEiqUZS/Ph4PTB2UC6+UqWbMwtOQ0JYJEzmaELQ
pVjUz++7Gp65kq8lsAS26Fmh4wRHbadBtlc19HykoFrO/M1niz91TQy46ipvnDjedQ9mtLkOJAbX
jd8Yh+eKVv6TUacO58k9ZfHvCfJTP6QgIsLio7JQbywvjYymLwuHkoLvDH43oCK8Vj/y0eSBJRhg
5EvRZ+ycWUgtsTyCKVp3OaoQVcsnIZhgju3mVFWEOojMX9xg0EX3jGniGWfLteqL+/bYtTSXRhnt
LJf7Q849Ru5HBWfoGOyLLk+snAjbC6WLYWLSzZveWVX9kXZmWmcGEfL1NviBTy+RnXcfFCv+SCBP
ywAzM6H/CS1z3V4OzU89Zud3a1QNFq4qjZDgZAwtC7WXZeLiUGDLwCdLWc/il+NT2k/g/AoL8Mjy
gsaoLfXJeOtzkGUQddg2vvLav3WA9kt50r+aIEt9NQs3+eRFQq/maLyJg9H2lHHtf2PtRy0yASFb
E281ynPckSx1baMdvXM1WQrorfQxkR+iT7lsoePTK0dWp3emaXGeUtVhTGLee/vIBgvOqmlgiaS/
gNRjnrlezkzZUb9Zh8LVSXMim8eUPYSi9DCW/AJEui0Rayk/vv16Dcl5+cEuhvkAc9YezqCoyiL2
OvAbQe2WcKfeRdaeZdAa1JQ/jg5TYX17ZTmWCBtLvMtPsB0mmtG05RluOc7MBjlQSDbUeKc5f7iH
GwxjQHddfQS9JtPynW9lKhkmAyv7hNvV7FIPY/7/KFpFlVhc0qRDc4C7z8/Fs9CdvIOb05auCnFo
k5wYKdQJckPuycNl0ASEgx6ecRJdOCnYkFLRENd1Vi//C2DytNebKhRfvGsW/vuo/BN/ey3OxQ2n
IsL+Y/7S+z7FunAfJeDdILntS9UXC+1wl2lsme7U4a1RDbLB7HF8pJAc5wyrPjFR3eRgWr2x00wQ
tbiM+XpuCXSD6aSQn1Ubq5KarQFXOipGXvusFQAEYiSTnV/JY0Yj1eUVKYFHo4N1Mphpn8/nL8mD
BGLX14Y283OPn4a9ZtAO1UyHJSSrOxgnRDI7ly976AVg7CUk+GUw9ubNbfm6GfL2L1CaxUtFguJz
z/xM81YZU8ET7sZ0pcIlxUAg0PP7NUjlybnh+/q481YkcCtDJUBnq8yZjLAK5jw+IPCVDem1s4DN
+r3aXm5eDBuNYQ7jG/6qWc4r+cQTuMN2ayQWTgsQd8MigUQd/8EWhfj3SnZd6vNEfChGh7PPxh4y
T2x4xJDSEu7h0uPZJYWKifB8lXLZLtcGxuDgbrrGv8JcIZQ63RlIWChv3+ZkvjaJ2ji+LHaOJnkm
f3p+oppwScZmQlMicb/Y0/R6+1uKiTJhwCv3RR30QMugqKgyCFAnYCb1uERGigA3XDsTL0AM0+ss
2dYSIJfZ146YYV6Ydy6Gn8bdIVroEf6wpRa2/xyfDJ8tWMOMc1r4dAasrYr36DNGq47Nn157iTZx
csWlhtopv+RJFxZ4P8ormkoAo+6NqV/hK36yEgs9VPL28FPVJzRevxxYIGztoq8/JXc0eZF7HdMK
6nsqz7rAzzaHOSTqlODur7YpVuOhCk2Lm+0p/TPUcg5DnUmST64loHKK3GTcQLBx2jTvHyV+O/CP
9px6RNA9S8DRrHR27MLE5RzjDDcXAflVlRR/P7mVZa++jDFiOo5qVAGmIA9Z2CpP8209RyTe5f5Y
e1hZl/eJbUAwJ2ipfZ6BtYCpLcj7F8pKCE+IBBHdjJ01yqxxp/7UNwOgl+B+mVLRIbfwFCej5CTf
VYGism/8yeJ2NmGUxLdhYJiUP3vVWIcVUmz+zxD2puxwhFdtizWrQ+yE59r7Tq+Dj+xEw4p4oh9i
Hz42EG7xNzl5UyI6fMwlqGTDBGyW5GIgPpHRurB3LaE4j5+yp1ksFAPmhqJHDrAffjA0cwrd1M9F
GxgQ4MWV2PvgEJRiwlFnnOvmS+C7BkxFH+BXekydB4Cb97oGoCH8DagtnAiZkTnO6z1u9jTYD3nJ
/qSUa1YQiAaAM6/5UQ3szD5wD91ID5rSPgcqDvZATzy7o6ZinWUqhAnJtc76yExPewoZKIoRgI7A
NGGPsa9/Q7pBp85y+vDYPr9HFRwPDSinVI2qM9xaZcZ+KNMqKJiNgmJ0WIfvC/+hyd3d/doYqGIJ
YHHfZmIcgPRwWmrwe6QkEYibO+4Yyg86hmDEn6x8asZ0BQag6DFU0gfunKIGw/Rs1gtXbO3DPrMN
3pp6GA1qKpr9rn/YzVCuqOTMrTHkr/0EWa5Z8zIKNLBI9oywutrYgCSyzEKEsS/gr7gswmZu7QZW
9EUQz2pScaNsFHmG9UatF2n8pYF/JsHz8oovINjLLy7z/88zfi4NYtRlJqZXm7yo/R2rEgA+FaAo
L393y5EA0psuiEbtL/tK9bfSLMdFJMo4seTmSzeQUz1+ZiF/HJf0yj4Pog0wW4V09OlCBmjD6GLG
lQvUZwDpoFUK91YexLeAp6wgFxpUEBw4OlepwxgtdtRhedW8cPEVxS/Pt1akbBqWFxFlMYFGCzKF
Bh93eWXJMf9WyBS569/IZTLLwn+9MKlTcaudCNTPuS0vzq1wvVJsIeG2t41L9YNn0F34zCvYgNfC
prDJGYR1rP0W/RFo0ezOqtm6YwKXuYu7leRbxMQXvWlC3RY2ZxVcfwMPsLmgGrJXTtyRpCA8p630
HAmtJuCuKgDNbLS0m4eWD1YhsJU3X1FB/ikeRfYLwo8GYNXGxGpuaIG/0NP3EsfhlqMNz3GeMOxj
4aB86wTtzV0N19r0NShpCKBNSQcUwH2SzA3/LqvDMAT7+DrOGfHrEZKPCt/o2x3QTNdEXE1R3m+T
65j0XrFlpcJXzSSCZk4buNJcU1q/Dib4eEWOoMy+6jT5eX+68C0pplGeM8xcRppJKpT5OxDM413Q
69uhg2srXDBUx09NPzNI9Vwy8/QNk60og+hOiC5HnPi47tOJYpoW9b+47QhA5EoO1bMVhR+tA8EW
oCT0sTCSsu4DoUiaC8SYSCwGURBfsIK6dYaedplVLlXrQaDGQeAgW6yzGjbvELVhVdIJlgRdT+3E
pOIC7N5e99wTnXxHlvfxkglkdFEyNZHGBlwL+Fq+8PIXJYZdM9fKyKxnZBh/joX1Emwoia4GSy9A
ScboesXx97Fk7DKu+3/W+OFbVwkaOgSMWEegaAkQGMm6Fgddrn16v1zCiRtXa/QgDAp02KOQG9FD
BzIuaor4FdZknnt74V28l/a7ZzjjbvahQ/VlTx18MtlITnzMOrNLzLuJRuqIw4ztaN9y5LkCrEUE
S4d9S4HbYZWkVQk7tcv7JNCnLuqdMnphjehrb48sDmA6r4V3qHq7tQkZG/H/rRS7NWT3ywogFG4+
drBpKCZwWkthMqmWiWRCdGTlaw1sop28Ecux2bZ3c0aBuTAFtwuT3ArTHD13jD6cBFynqzD1CS2x
OnodFuUOTvLHBEuQmw5GALyxBkRYNJ/2OtywaP9wIofo2HC86VheDqyOp10XPHKrJXJdz/Sx+Mi2
cbI2Ctg7ZgVj2oVXFHO3HyoPv+I2oVSNc1A0xn5cxVtHnrwwCHN7awz7G9GbTE5GKCr6qYyS/qaq
/BqaKyCwDH8Wa+k9twQTNML3h0J12JYp4NTYPgFIajDs22aevHDN7V5Zjl/IovlnOT20f+55JW7L
94DOmGi8/JEcYVnOchqVmKoH1uWoTywELz2GFfJb68ca4Qn7aczB43gbW4j4Pl7RJBQRzqFqUPLv
CCmpTKoI6MTiwnTp5gfHNetwVDIlFQaQQ/d+ybM=
`protect end_protected
