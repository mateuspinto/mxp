XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���a?�2��-�S~
��͓�XZ�뢇FVx�/����L��c�HY��Y���.�*���MS�n᳣��[�8�R$סN��x�uD�M��aާ�<2�vS���w��q�T(��r��0�Ղ���u����
QV"�ܽ(+��C+B�m_�?��y"\��>�������?	ze�w�z,�{�dﰕi(��p�lq����W�s��Ȳ�i袈�=���H�t���
'���[O��� �6j
��mԽ�=`1�;^0D�T"��Ta�����ND�m%
,:���`O�����y>:բ0����+X�w�[�MAÞvNJ�E�U=р�C�)G$�~yew�0�����!�	��$�iC�6��4P��f�H�:�1��o� Vj��2:�%����@����R�����M�TDX�I�h1���׆w��>���v�Y�Vb�W�����]@P�p��vn�|X�>���*�}��_�.��+������ǡM4�vE��5��T��ҽ^\���=��M+H(w��
�-f6U�W�sɲ����u/xH�M&�[��ZotK,<���W,s���]h]�3���r��0�:A�u����}�% UP�؟�-�+u�F�@�m(}M�� Ab^�u���b��'�f4<�L25��6�ɇ�7�����Bݰ>�}�+�ï���3�/ƥf7���=���U:���F_OM+�Eϛ�MJ��r��M[tm�}����x%u��b҂�b �Ã<�^�X����j`#"��x�XlxVHYEB     400     220�g|fbTv�h�P��:�����.z�U����w�=c=l�:�
���{��M"��n�ۈ
;C�f�f� �5`��E��Bd���6V����b7Pb.5ڣ�K�$9��Z�n����i�r�S��^��z��8���������զ��0G��Z��m��C�w��A�_>wE����,��C�Xۂ������]�k���ǉ�Jk,Wޖ"8�X��!��78���Њ�;���oS��'~)"�S�E'��N��]������$��zw�s;7�ߤ�T�y�,�����O�t��\�0�cT��O&����`O�q+��)�CN��f��1��N��R�9����'��a�B f:"ZX�QC�w��s��+n�20��^��_�}�c��˩���R�uL�}�����z��
��6o��X�u���X�9�# !�Z}���}x���<�l;3��L�v�Fk�[�.]}h�.�L$�ӹ��t�E"9bW]*�\��ت'ΏVo���DP�ZfM��A��^{$����e�J��N8��,�	~XlxVHYEB     400     220ДCʒ����#GoF�w_���(��Ԛ���)JI`���@�E�}G磱��X�����J�jP_3N�����`��[6�G%��w&
*8}�z����)��A~���X�z�_+o���J����^���t�Q�*�~{�0؏����v@�@ª�w���.�;��Y^F�����f�<ܓa���X=��N�i��,i��L�+BM=!h����D�䲼�2\-��#�}��o�K9)�����������n�!��L��BfԟP�A��x�Z��1!��2�{wY��� 0�����Lhg��B�q�LI��U�J{�Lx�+�	j�%U���zo2ջ��/P���°S����9A易Rs��#��u��Jn]n�@Pu���?�;M�gY��2����SV�������?�mk���%�2�b���]����xy�qЧm��
7����ak�GK��Lns0)�`V�L�?���Z�����2���Q/�H��"X/�(�d�O�鶏�03�⎵3�M�'+6l�<C1��tLF�K��ur�hXlxVHYEB     400     1a0+��όq��Z��z��\�qen@��m<.�of@���?�B��k ^�oAm�sh�1(mc5�r5�5���?���J�`�5�s�8/8וU��pݗ���R5�ʈ�{´ t��tY��h|'"��څ9-n:j����(�}��#*	����s���X�dP����Ѥ�:�	zV��hK=�*�N��칬�[�>���q׊M��[ǀ����U�S�F�D���t�a�O��,�$a^u��@�8�0�D��,��1<�S]SΧn!.�P�(�Q܍�H��u�-2�֢}�������@�<��dF��=*�*;�^r#�0�S��98��|ڭ����ٕڢ��,�ߘj說�gݿS�bY����>B�?]����ww݂�SChSqB4Ja�����ָO1P?���c��[�r҅�+�j�j)RQXlxVHYEB     400     130�Şs�4�{�8��y�/�\W�&V��HcL�,�"�C1\=P��g�=6Y+7����N�O
.cC�O_�c���{V&��(��$fk��>`Y�����&�:���7~D1������[	I�:�aK� �Xl0j8�DT7�m����_�D;Dj�1w�1���t�}┨y)9a�:� ��S�� פz&8I!�m�!Jog�_/\	.��hs��Y���|��(qI�F��<�R��<^z�9� ����M����� ���^^KX��dRǡw���2�W��e����YS_]����XlxVHYEB     400     140*�����;�/�#A�iL�\ǽPLP(G>��͇r��R/%��t�Y<	���\��͛((g	^3v��U�_��d��*�y�5���x�V��j���P��촞X��5H���v�?�86D���K) &�1��� o��+�<;N�*B?\io���ӳ�9;�@�u�����F�� c	�؎���s@�abœ�!�X��Fa��q`�<�x����y���'BF�6��W$Tyw������	�����垏Z_r&������#gǐ���)Tx�;̾>3ОjH�#x�w��M;���I�%04��մ��a;�@r��XlxVHYEB     400     1c0�(�ۡC��,��
'���J��ţ>��U�������Rа�I��'����Zn��	!�dQ~���q�KO�Sr��R��I�w�<����.���&#��Ə��E}���Iq�%gY��N�܀��s�zb�S��|�>E���~��ؓ�kc`R������kOA��gG��8c.�n�t����Ϭ�6�H`����F ��
E�3�Q�>N~�]�}����J�>��C�����PX0�4�e�'�9DҲOfR�#������e�U�� ݖ����E�2.��װIn���3��5ٲ]i$vb*���҆;�����/b@��T*�40�;��^��w�t�R��b����@:��O	s�1)����`䢒Z�cz���1���Q�d��p��Cl���Bi�tZ�L�J�A":���!2� �
fUă7�$XlxVHYEB     400     200�`��n�N�K��)4��ȍ7.r�u����lB�;�|��(���?i��SP��Hn����Iϧ��s�@����}��V%j�3n��g��"�AU�����Pu�ߚ����lݞ-�@wc����x|
�`>&�������
����Bm�Ӫ-��cϫ�!f6B.0���f58Z�
�RN8L?lw�����y9�M���hE9X��eT�v;Ґ�R&s3��ە�.|	@,�|T�u�v��mpk��J���9��w�7^?�Q���0PB4}g�?��/3
���+��ĺ��k����J�?�A���EZ'0��|�с����*�UO����s���Q�����o��� ��������#�).�՝e:��'HXe�uGlQ�_!�oa�C��i�ٯ�n��guߞ���b�Z�Y� ����J-�(+L��j�1�vSf�졷���s���P�6N&+�;��X�Q�9��2e�E���g¬�8�,bt��X��'�"O�xy+=XlxVHYEB     400     1f0��4�<��D��.�&��)�O�����B��~�uKT>X�e9ƺ�X���E}�m�G�_�n�2��Ѱ}�"e�7)o���IP20��Ћ')�^�2qFܐd�g���c�f{V�ǔ������>��瀅k��;<~"��Ҁ��~OW� MN�ʱ��U��e2�Kቿ�A�[�E�ig��-�wR{�3>E�(�2��6�_�1J/fb�8��Y���45�H��i������ZBk�p %@����@�9�F� ���U_"�W����ه�F��w�	!�E*O�wc�H����vz�
�Pg;�����;bXl�S�$�N�|��T��UL��� ��ya��DZ{E�kqq.Q��*��:#$����h��٣~ď&���C�]�#KC0,��s A�0r!Ķ���!��RI�:6�ߝ^υuD)�0X�c�"~�S3���[l�HjuU���Pҧ;%��4�w8�{��ADCl�Q��C��<WI�u�eyU��XlxVHYEB     400     1e0AvXs����j��H$��yŌ��X�X̍���L�i�k��Nʃ9�2\�UM�2_�W)z/���X�lS�r����HX-'��H�y,c�t;k6�ʢ��V`��$��[���MAIN�s�Ũ�
�-�y��#��J�e��߯�VXX����j�c���Y�/��
�4d�|E�\�QZ#9��=��d��"� �Ck1�U�����3xl�*5���WOa��H(�q{ ��@#j��V��5Z�/�K�ڙN8�Z��`6�|U�|��w�G���'Æ�s^�U~`�{-�е ��_��4Q�"�����8鼃i��k`�y/��ajFMZ��[�>o��(�.r� � �
ϥ��DiO���^u�>�垮�ĆS�m ���{,��-#]�B��	L���!m�~�o��C`�,�Q�ߘ�]t�F���d����&E(��G�����Յ��|p���,J��P6��Z�J3�A?��PXlxVHYEB     400     1c0(d����E�"��m��=͂g_ꓬ�?�q�M�1��K����
 ۫i<]�?1FN�M"��	2��~�\T��$m���zQ�Gv�e?�W��H[�w��#���l�KY��y�#����z�:6x �)�gY��eՃ���c�#|�D�kOוޢ#V&�׆�9(rl�Cc�xd9h�2?� ��d�?d��?8�����2u`D����feܵ�?H̭�:�Z��s�6U4+|�g9۴P��+�n�W �VZ�tk�:*:�����v�(iCn=L��
!�ub��f�Ń��V�ȲѮ����M/a-��go{�O,�p�V�ƧҬb|�&XV�ƍTV�P�\>��@�����AoLW]�wv�Y+��2J�r���3ۭC�Pxڌ8����n/�n0t�ڗ@��45e*o��F	�Hi�?oA�R�#��5��<=�lHVB���K��F<^�e�UXlxVHYEB     400     130w���D��p�X�b���uk�]��u�$0��뼂���ΪV*̧ƈ��ݱ�؛���"���xt��=�&)�+x��n;���w~�]hÓ���V�P�QK����x��,+��G��>*f���U�Sƾ�r��{Ùt��==�A�CQ���mV��}��2�� ���<r_Vj	&DCМ�����u��ݨ�����{�0c�:ڱ�9�}_\�E�N�B76�qr|����7=^R���fH��7�jpg��؀�"��O<v9���*S�#�gF���/���8"0�!;�T��B����uٍXlxVHYEB     400     170���+�}�7i����1�&o��V�ב��n��fD!� ���#�)B��3��כhS1˃��藆<n�+�M~J�{PF��5MK�����|6�v��v�u�{�;Rp���=�~�I
�jz��f;.�n"H�xd��>���i(��[Pd���G.�w�͑�-j��e��w]�S����ю��=Tll����Ƨ������b�i�Qw�96ɩ�udG��/�P�v"���O�ԯ���#����|ݚ�#<��ِ�Bq��-J,���9�t��K���T\2�J��)�0ϔ����ͫ9������^=f�\/e� �A��R��O�����*�{����5Q|�V[�/���XlxVHYEB     400     110c��6ϪQK�M��(�lپ��zq{IVT`@����#���2T"~�<��4�¡?O�o��Q[6ޢ[�x'�{?Q7�郿jDq���GM|8��X5�0_���5�)o������Y�����s]wn�~_p�j��\�.�3%Vk��;�)6�[��Ll�n��ؕ�H;l�b�S7�N���(B���\�)j�b�$������6�݇�M�����$�c.XkE����*zt�uIڸ�U(�_�G_�󄗤��rU�.����%���i}�,�a\XlxVHYEB     400     140�/��a��$Gi�k73�8�-r���"p�r���O�9�abB;�v��%f�["�^��Z�3�͏(_��������uȽ}�4/��)is(r��g�_'�A�
���%�0�3��9�"�CX����M��ly�k·��Ye�T qօoӬX-d�R����\�{���0�bl.d�i"���(�Rh/>�!t�P.�������Uy��v���b.�M-�xx�HqQۀ���[ǛI>;�R��b8Ī3瓤sCqYq��}�*��j$�C�ѣ>��o͔7>�)ѻ�1�9��L�ѕZw1e����n�����͡g[u�XlxVHYEB     400     130%%����W(�d�~�KQly�eH3o�\G����ŧ	·�R�CYyB]��h~31�5]C=A�u��|�u��v��&��t���m�w�K,q+5�o��2�����ʾ�HAS|V�d=̰ѭ�,�q�h8U'ɑ�ӏ@c�Σ y.f��n��G���`��D	���6�)�D�v�֊^�����M��+�8*A`W�y����*mZ	�y-�d���>�����P�3x��N܉��$'ahPn���7�E#�z��7e[i��?� ��'�2̣[��3��`�u�փ�9�M�?XlxVHYEB     400     130%�ԋ�y��k�<hѴm�?��xXeti�F;=�%�Qf��[�AN1�K>�H�B<;�Y�q�Z����eGN�o�0�k��3���9uݒ]�6�a�q�)p7�E���$�L��&�5��P�XUy�&L��ގc���I� �_��Ͼ��xn���a3�h�T��-;BV��C�C����P�>��p��C7;jA��%��e6��ҳ}A���O���������T����\���Y�>X��o\��{N}�q6���q �4\BJKN)	�)hh`w�za�#�k�K8u�yr��#"��C���O���]�����XlxVHYEB     400     150$��������_��G+������y���X#`T���$��ꏴ�|ud�T>�l�v1%��e��j�\����{��3��j��]������uye?:Ҟ�R�עΪJ\�f�]����&w�>.u��� ���\o�wdl+cL���~	��-�o"��r1������>�z�5{vﾊ0#`̂�6n%1�*"�a��p�J����\T�D���<q��}�9�t�h8=���6�	��c�M��0t9�
qq��eI��^�P:4�y�fzv��(h�;��b�Q��DIn������Z�����
�:�N^"�� ��d%j<���+ �d����a6;XlxVHYEB     400     180���m�#�՝��Qf8|��(��Ck�~�����7�e)�IAN64�Ekxݹ��H
�5�d��yR��
�Y�-���o�/o�~K萝h6�'y~���ܤ�;���[v����*���جx�c�w ٤��*�	�V`��ty%��{ u�Ebe��K�s��~h�m��u1q��7Կ�8}I9�,I��|!�0�n��������w���4ڮ�:�sB��j�2�]*�c�[��`��~GC��\��AI���-[�y�}��I�^���p�W=��cޣ�؃]
f/�T���hqǜ�.c��U��i�}�^��(н�;��7��$M�9d��Y$�gh��.ވ1��
9����95c��Ju�6q���I�g��Ijm�X�G�-K}�x��
VXlxVHYEB     400     1d0�&�q?Y�Qĭ}- ��%�eu���%��X�^C�<"���X�Ʀ���!��d��� ,'��z���#�.�g��.A�ߡ�^k$ui�]�BB ��M��u���ڀ#21�%����8��+���	�S4����=��i7��Z��!�pH�|#_���:�FA�i �Z�G�����ڝ������D����]����^x�9p���mȜ���&����ώ�
�`{�^�Xړ ���Q)���w�J8�GӁ��3���0/����B���=?!&cX�6;K�������s��h+�wf��4gP�r�S+�����7�O%ld�Ck��%5m��=��}2��ܾ�H�@S@��h�-�C��Տ�.P;�H�P���l\��y�;mK�U�q��o��N$���`5�����o���|r�]�7�1�z�)�E��M֨�g���^XlxVHYEB     400     1807H�$f"@Ls�A!�{ �k���ͦn�v�6}	ǹ��kQ��Tފ�}jc-�sp�2	�p���Ot|K��a�%�u�1�'T�9�x�6��ݫX���H}̴,*D3��;��N�2�r����+�ȶ����g�D�\��h �5=dmA�@  ������߄
�Viq�^�����%O�S�o�#/Zm�k|�A����������ak��n(b*�UNpu�@�uj�F�`���C�#xAq��}Ap��O��I�������[1��M5����ĤT�B����e���5��쏵ML���7hE�?諗�)�
zT����J?m�}��A�{\bt@�����R?'�ϼ��tk�:�'�J�>]0WƦ|�NA�3W'XlxVHYEB     400     150S9�,��`�0�8r����>�)G�H��#'/�F߃Ž�����-��:Q��.P��x��t��CL�=�;y��\��jW�8l7�	H��@ɵ��3���r6�s�GM3��t�Ľ�e�EA��·�ÜTc��+#�	�C�����7�7+�~�I"�u�S3���8܂c�~����ԫ|-�����t��l�B�h�O�B;*0�V�]��j�n;��Xyo�)���5�L�f�q�,&��\ՅTu��/ܢd5Јm	�5��!P'���d�2bGM��i��̙�6�F#]"���Au�^/�ό�F!w?evQ'�SL9)S��\��*1��H��+ͪBZXlxVHYEB     400     1f0V�(7R�R%ꁹSRό0�2*���aX'�mT:ZH�<h?�v����s?�.�+�2�W�������2�u�q� �ôY~Q
�i�цqr��e���A�K��R#���0��6�N��j3�U�ޛ�BP�OQ��>}�T�|&�ҩ{�[CcUdP,Y�dw����Y�E��::T$�M�{N����H����$�хᨦ�[%�� ��4/=�i���t�����E�`>��$�Q}3�8�v�ө�6�$�;��3&�K�.���:�λ(�I���Pl�Cgi�F��"-��3V��	����9�Dq�R�5H�4�3�~Q��n���$c���L��t�^�zB�W�w��\�^�J)��b�5�_JÎUG�J��K)��{���?MJ�X��m�K��7G��2 g#�����	����ԛ�������2bP��!ŭ'�Ç�g߅S�~�)"h�NN��,���=����UN��a�4r�P��b{>lXlxVHYEB     400     190>s^x��}��e=�{*\��8�uU�Q3�j�"�k�֍x>��tzX?��͗LnP�"�3�iy���꾶?�go<d�i�ݘ�LI�i(�P[��f�.|�a���
wZ'	�nh�5"���|@8��$&�W�P��W��AK�#9�jKi{"����57�rM���mz��c$��4NS����1��L�ō�!����'����֚�+J���X'�̛Vuɿ7��
�D�Y>�m5����OC`�ٷ)!���Wֿ��v�V���$�h;�7i@^� ���v�����r�
k����q&�Bґ��QF�cr\�8h�&���9��Lߋs���o*��G�D?�x�
�8��$6/�����!T.��^�6�<ݓ�7@�OU��Un��r��גyi%��V&��iXlxVHYEB     400     170���t�{���_�RΦ���c�t�p@�� P�Ƴ�@9�=��Rf2.pށx&m�L	��@���lwZ���O����y`�X��_�[]��#챯0�4q�Q�Z.+97W$X9'J�Rr���T]��I�#8ßMz���DȏUj����w��D���qVi�B#�"w�FC�3"�o��[j̋����L�8�U�6y�[�p����zi��*�����v�}���X�Q�&�'�n)M��P�qb���is[i����g��?��p��2�)�cK��۫�kB/��6/"�0����)�\���%�r_W���cM�xoe,�R}�ٙ��أ�d3��Jm��Ĩ�u��"��(�o�ꆷL���1XlxVHYEB     400     170��?�V=(�(�2���Oj:����'�U��B�@y��$��^�]<�]?�7f�L���%���դGm��(�\ �V
�Cc6�;�
�N}�#(8ʤ V�����\ٗ,Ԝ�S�DF�{p���;�qd�����mL�%r��](�VFʰ����߸a7�J��v��6��^���_��T�q<��~��y���pS��o�´���x0Ve��@ʢ&�;O��1 a5w�r��<�(m�vk.|slJ~�u~�ǘ�}�-Z�b���U��S5A��l�7���,4l���?+���;k�����3D4S�B"�{(�L�?�=(_��<j@�A8)������$~�Ul��3����
��d n���0XlxVHYEB     400     110��i&�@�(�.��LhZh�v���}��I	y�/�bD�Ԋ��Gng*�a ��9�ge	�2�Z�ݎ3�K��c@�0��B��ŋ��+E�l� ���[0+�W:v����w�':<d�C��j6�uMgխ�Q��D!g�y��da₋�u�c�k����'�t�,�~�m�el��Nw�n�d���QkR��xDz�$�|����6CǞ蠁Qϥ��-�e��WR�T7x���篳5�	��͉o`��
K�8E��x����jA�r����$b�0)�XlxVHYEB     400     120%\o�]I� [�&5Ttն.E�56��W8�se1��2ߨ#`zfAX�Wq��XJ�ro�2���17��^�����SAǈ�Y��	`i�Ȕz��!ٕ{����� 2j���6�)����JI��	�[�*��%Њy�n=�cl��e2t�k/�G[�;L��vI ��бӚ+� �A�+���/Q���z�-��m!_i�+�O���c��y��EŜ�R%�L�U��+�Zz��x*�����6)�o.�	 �䁽�*$�`?[+��p����0*7�;oA�'���XlxVHYEB     400      d0�$�<�G�ǵ7<����a%�ַ{V�NV~��t�Y{ ���0X\�`�;rs`!3�����7$Ȭ�m����X���
i�E�JI�\��|9�G���A�j�M7��"-�Ê!���J���N@���ݡ�&�J�6�K��D���4E�f�8�&��נ��:��E�ə��7�8r�!���Y�xA�=|�'�F,@kXlxVHYEB     400     140O�x���34d�(�q�V3������E��j#�>j��b���`��19�B<��`054)(F�M^|G�~�v�4������1Ș��@���]2��(u�-�<�#�|W���B��C%�	Φ���Sm)ܺ�B#�vx� br��F��K_�ԯ���t��;�:��)>�pO�^�ڪ�g�̻ڶx�� �-�)��|�Л��iwZc���{C�v�fخ�̯��67�3��y�s+�����c�߲�PU8QvX	3m�T����?ӆrY��W�m�����s��1*�ҡ��X��	�� �l^a5����=KȀXlxVHYEB     400     140p�JD�i��PZ��3��H�����|K%wY�̂#A��ہ���dQ�����s����k�r���~pj�Сi$]Ɲ!�VF�?ݷ����#lʤSGր��<訑G����� ���,ܼ���l=�:�v>nG߂�A�*�37�
l���)�C��s���}���޳��0�\1lYe���ڡz",���Y��A�`HO #!B>z3�/�^)f�&r��j���	 ���[!(��C�*�z������� ��N�k-0x�4����.��������+u]t<���Fs𸀦��ԮY���XlxVHYEB     400     120|�h��	���	o�2��z\qlGS�#��Q�8D�@p�D��hc��P)1Ƽ��y4Ӊ�>ؒr��(�yx�Y;_y�&�8�I� Eo�ܣ�����4�t~o���=��椛���0�k�W�b�:���.s���ư4~��W@��ǧ�$���A'��Fp����M�F��'<X���;�f�XS��sN���7��mv�&�����m�|�����zҩ�;��U����P��*z�ޑ˂^����f6M�-A/HP ���e��ǉ�[��p_.�}�0J�RXlxVHYEB     400     1a0$S�zv\���w��}��Ì!л)e�+Q�hm�&*�Uu������q��q6_�D��!y��ܯ5ڛ�z�H�Ǭ�Ӹ�&�uS��ë�w�}L��\:aG����P�K�ˎ>��(;����ں��4Q+s�lj��qF�w���T����7F��z�[η��Hp����U�0D{�脇��̴4���
p�G�_�<�%��P��$NGf]f���;$�+����=x�pc@�
��/M3L��&[��B�?Mc�2ҁh���ӣc����P�7#�1�j,3��c�|���|o5#����2��y\�2�+��5�@Q4{�H/hF:�-�@u� եo��z�6Z�<.��@۵�U��@�����S�z�_VǴ�c����Yåњ/�N��3���yn�"Zn���8 �߇��x�-��XlxVHYEB     400     120�cQx[�SG�fݍ6H��׈e�H���m���!0qj�l��
�R���J4�x7&_��@�??��.�Z���@4Q�oY�%�MFG��/Ɔ�ZG���6,
(�A�����^��˟��J��W�'�$i�n��5��5�>��4��
j��&��E&x�k�>�<"C~��G���C���{^
����ٕ��l�$�>s�����+_�YO��ɇ��4���VYe��ۚ�8:[��{ qB��u�c�%���/��W�ml3�?L͂"8���� m�~�Rtvv�XlxVHYEB     400     180���u�F�ʗ}�g�%6��v�`������,�<d͟�	�cƣ&B���	���D[��r"$�h�2'����ָ�x(��Ꮶ�A �k��z�$�\�㧱������V�&SZ	�������|�_\��	)�Ⱦ�Y�E�B2���|��~�>���i�B�F��cv:)�Q(h��Z5157۟[�V��N�e?GF���F��'`��������p~��#��)L�+�/H �r�Bfଌ�9��|a�>T*\���18j3A[n�:�a�^S����],���]�e� r�c;���������Z������ od�t����X��^���u�.�d����������P�-?:5SU�A.CneD�+)h#>��XlxVHYEB     400     170RR��`a�2e�2<j��جr�MSV΄ҴV��9�;�i��įpr�O�E��`�^�����nCG���p���T��(�H#g�j��Gryt��$�Y�Q�_ٔ��6'�)���r�U�����������-���� YA�T7'�J�R����6�4{�"J:�.
ST���2�E+U�BQx�_��\[�+�'5Iq��4p���01>�JV�Z)�v��'�|�6c;[������q�����3eo�_0ӟs��L�r�}��+�eeA:M)��T�;N?�7k1]I����Abq��t�4�Ov��/�`3��@bq��A��uآ�ԏ ��~���m�h��D��G�4���{��&XlxVHYEB     400     1c0Jh�&�e�ݧH~�˕�Kt'O�bC#�A������Φ��"�2��_�؊���
��t?�pP����y�Sa��Γ��Ŝ�2}����}���^�W�&,��ffk]}�#M�gFy�eDO.�J���Iެ�����(ݨ,�O�pO�/�:��#�SUP�qgr�s�x�J#>Sy�/d���N��$:$�$�l�A�//���ȷ8_
U���y�1��^�~%�:�$�����i���)F8���1w)���X���X^#H
�h���h��=���Ww$#�O(��Af0m��v�~�������@�q�3e��:f+�����l>D�g�|��̊n4��jgI��� �3��@&��/Xr���Ξ�B.7�y�B�`;U�ߏ+J�9�˼[�[Lt*�c.�������:��h�7��b�r�|��O�������<઻N��XlxVHYEB     400     110Y{k"|R�7�N�7�F�>����ez��M�$����v��b�i��?�a����2%M�Z���A�ƹ$���u�|�,�]����얶���������b\ej�AR,U�ͻFj��?�V?.'[�L�L�W�Z��F�hV�.J���'E&4h-|b���Q�!ڨ5����3�d���\��l५������KM9�3�K���)QR�e���ԇ��_����+��?NS0�*X��u�c�QT�;�g�C�����!u����4�
XlxVHYEB     400     170����P��=��ny2^�y
o�ZA��C�����&`��z�m��b��EeWq��AN�D�/�M\��}#��؎��v���6/ǗG:*.�>B0�	�Z�!��s!�R t�CA�<�NQj�p���⽑&�<�s�\�=K�Nى$���s��h_�rU�{���,G�Q@���'�_9�tLY�g[��즙)t�|��6K���|w���q�m���Or<�l��P*�e���mW	��J��kC kK���m���+�1/&B2�# ;$�c$p#��DQܲ}�#�D����q��'�?�8�8Y���}*�|��n�i�Aj>X!�@��?�'ǈ��I���˙=��A�2�4f�J2��XlxVHYEB     400     170���VP\�$���9a@��!hg����	u��H0������0f��������c6�'D���t�l�:���B*W^ȡa%�[����w^�&�m�-M�\W<���~�}N�4[T�Pl�V�� Ү-v�a���_�jh��T�e��-Ɠ�Q	NSʁv����3�HS��-���������]�SοT`9J�����$�߽Ìm����6`)FL��]U��s`�7�ޮ��U���e\�����(�E>-C�*�rE;+�p(�ލ�AQ�1�;޽�k����@�@2�!WS%ᚪUu!3���-���w.gtJ�O�b�O�s�г�����}�ƥ���]�]C�8,�3n �ث��[�sXlxVHYEB     400     190�|?���ȸ�:*Ӌg��3�ytlO-���B��44�|�K4*�K�r�ʘtZ#�0��]Q+/���kSn^lQS����b �}�P_D���I���4#f�|�� ��0��9U��G 5%���xv���BVp *!�$B��ἌFE������kwbҚ��%����`�sŷ�:����nx��i�:�����_5��+-�6�k�,���/�2`e��/��u�ۥ{��˘>#��-0m�V��5�r�i�\V}����Cy=&o�x�:Fk�[�\BQ� �a�D���ш�Ѝ>%���Ld�L����4�aP��!����S�}%	pY�tI��[&$HmI+�*ǑRUMt���L^�O�4V�9�8�q)����)!�Mu��]V��ӓ�:XlxVHYEB     400     1b0�bFH�>G���ׁl�׉�Z��`�D�	�U�`��m��S�����<��=!��=:�y#��g{)�g�\��!�d��^!����\}A�&�l��u �{��6Z�+�G������7��b�����_��疸x�U0
]��4�qqF�F�c7��`|� �`Ԫ8�&!>u��~T���|��G�)�qL���H�%�f#�:2����6a��2Y��i٦��b~=�n�V��Uq���)I��?��U���$�s�wk�Ե�=ҺhAH�0��'��v����~�-q�����F0�-���ԛ���RU���}6�(���M�U!���)��F&�i�n6=n��^ꬵ�������/�<ڋe���_�ք�"W����}�L�����M0�1=����(�;*`�G�`�N�|>X���Q�(�g�;+�@���WtG���3XlxVHYEB     400     1b0_��ɨ���٢�"9U8S)��;�DiB��ȾZ�N���cҌ���]����O�u^p[HfP6���d�4&}��"�:6�ld;��9e�ͽ��E X/Y���̬_�����s@5^*gb���Y>eOj����i�[����S��ʻ_-���h�Əd�Fh�����'C�@EE�U��>��j+�/$��(��mJ�ϳ�~2r��A-��{�O�#�[1Ȇ����+��W��U���LA���1rf&]3�C� �|�����A����H%5�3�G8|�iAH����P�^�/M.v�����I�Y`;<��U�*�β.ݽ��B3��p9H?qx��tg��e\�P��?�=�%�T�Hv�F�v���][oP.3����E��M:m��m2�x��j`��4v��AL@��0��$F�ς�Nq.�%XlxVHYEB     400     1c0�:��!���ձܘb���~�V��kd��䲳�o���=<Z�F��/��ɵ� Xe��١Զ*Ph�P��Wˏ
%e�Ӽ��{��:���	��r��������67Z�$��7i���}Ȓ�Ｔ}�F�����Ӿ&!(�{(�.�dr|.�����۟�V1����-��U���F������h$���5�X��8�����/��k��fG�����I��W�oׇi��6ȃa7�JC�ٯ�5����G��<���)�m���Nn����0Q ��O?mS�l��iոr� ר�n��3���,ڑ3��z3�g��j�alb��Ǐ�t����Oҽ�dh�`��n�H��X�����P�p�zyK�=��X�c��0]�����ywJ����2��s5��&-����'�N���Q,K?�����:VBc'T��x������XlxVHYEB     400     140[�1�_�L"6sh,Z�P�"ƺ�įk��Z�9��Eg�y��_l��@��w�4eH�o<��p�߰�h�����\�/�N��E�Y���XAo6������3/p"�Z������FQ�G�9T�|~��w�Se�j43{�A��(�=��e*g�q!ͅ'�7� ř�\�Z}���C�u!�.�R��9te)����OG���z_����n�آ�t�� s�ц�01f1�8��/���w���L�yͻ�(�E��G���)\OdhY�w��s��q|C~��`J�%�r=��Ug�[|E��[�,�vo���E6ɥ ��PXlxVHYEB     400     190ۈpd��{�����w�C�Y��ž�ً���XQ�j��i������kD�)o�r�����՗�����N%���6"�.��V��ɿ �Es=n��O����cc	9�3+�h�ִn��9q�J;d.�{�����F��8n���M�������+dM���B1�-1����k�Һ����{��qZ{]`]NW?��?`Ճ%U�k��>Mj�a�o���I�@�i@�E�h�4��"��;������_r�,�:�M/s�3���N>ė��{�0��j|���{�����>���&�Sv�lv'8�*ݢ�8���T�pA���P|1ޥ��{�,��ogUf�ۗ�Z#�a,����$��*�;d���J#�	j��K��J��xh�J�CXlxVHYEB     400     130dnڰ.��b!��{�S���lx���\Ɔ�QZ32����@�Đ���K�b� �{��%H����x}��0�+Bl�	/��<�tbl��_	x�j�.���"�>3roZI/� �=5F�8��OЏ�Km� 6^�"2��dTu����dyUDu8= O�^f��lB��_�*���6�X7�t��e��f1�g�����Y�f���B�e��XG�93`�h��DE��ez�n�ÃQ%	�k�
��	����D��������ؙp&z9*�e�*o�?��F-�H!�e��V P��5r0�S�XlxVHYEB     400     150���G�����Q�/J�;��G�Uif?ɇ���ս�i��M%���i�V����&����Nvb˩ 'Ƒ.�Y���`��+E�uN�c�K�!o��8*�v�1g�ɶ��~V���,�K�&ފ81�S��;��q��T��M�\��+(
`�2-\x�TT-�~[|ξ�|�!#{UԞ������qz�TG���S����`�[�X�-s�;^�F�R�I	�s�\*���<��m0U�Oԝx�We��QLn��DI<�%�ݤ�)��*��Iڒ�*���,R%��}
������"�n�imZ��� vw��pl�Mp�al���>5�f%���x�a�M�{�{>�XlxVHYEB     400     190�6�4E�'QK�ې�9�.o c�|����Ҥ�%�4���S�j�����Q;���aΔ῀�/yp�E��o�B���ez�F��,� R�z�q��;�8��ƴ���\�Zi��x��-�.�c��+��J�w��dHՒ&;�BWҰ��8>]�%���àJbz?`ҡ���Y��*PJ5�J��l!�6y[%�p��Ώ��<1�ߣ\e�,���ODt�c^���C��M�=�?�4.lL�`�����ldP�8@]D����y��A�
m��nj)�qq�7w_�9��� .��Oµ:��]�qU�)\���p�?p�r'62�CRޙs��#�Ru3yF���p���3Ak�r���k�h����G/r�]�V��^k؊�Q@��,���x�גk�dXlxVHYEB     400     130?�R�Ni`GG�xG�A����/ D�z�Z�Uw%���œ9{z*l��^�fV��*ƾ�j���<���w4����F�{���Ҝ�Kо�*�.seۜ��	�.`�~���M�K˽��C�Uvѥ�rC#�&��"���/�/���?;��*���-Z�	!�F �N,ɠ�G;��Q�(\��w�7A�n*��l���F놨O���#��dbw;�_˱��Pq7T#���H���'s��ؓ�P,���

�KIsS� �3�N���(b"x����ϒ�x�_�*��7;Du2s-�Y��03�XlxVHYEB     400     150V��򖛌�0�6vJ�jM�prƈÎ��ܜs��O����*r}sN���>;�Ƴ�Ft<[(#5�h=WI���7h������mq��kW �YS�Ǖ���;��i��!�q�K5�/'��<c�����N�?_p�1�:�:�)f�#�I��������`��ܑ2�� ����Vn�����a��J�������(<������I*m��l��G�jh�'��R��ۄ_���c;�ڔK=L�8���@��ǫF:��{�tRuaŋT���'`�i�m�o����^y�?���_t}���NFps��)�1��ڀSQ�����_xf׹�Y־�XlxVHYEB     400     1b0Q���5��}�t�W�5�[b��}����ލ.�R1��K,'�_)�t>k8�*��I(�G�
�����@�O7�KGU����
��5�朏�;���}�Y���kǥ'3��q'>��)�\&�1�`C�)?�U ѱv�|����A ��
SG%U#�D���R��s��<�x�w����?I#����.�B���&��+ڊS 4	����xs�E2��9?�[��Q�{�����6a�5�k��͗mD�ߴ�¸i����.�V� Za6�X�'���(��M�N{�8��˧�i������T�v�:�}��.J�f��e�A����=:�N��h-��J��ty/=E�MEW���%�x:}�6d��9��mqI��ũ^�s-�FG����N핸xX\� 𙎓�*&yW4��4E�����V���B�_��Y�AXlxVHYEB     400     1b0h=�>�k�X�N'������N�W�[;���)���t#l�_y 7`���2ɣ��� -��a�� �I���G��P��|c��]�=��k��5Um�YT86��)�Ǌ�S�#�����Jv�ɢK�nw;�c\w>r��2�]%����{�,��F� �����[���޿S��d�������4��%oVK�00���� X��z���/t����v�s�!�V`������{>V՝�תuqOx@v�x�9|�	F�W�����1��dt��[8�v�M��Z��k�u�8\�@�o#�Ly�/
h���۴5�wk�ߠ�N˩��تE��H��owiRdu���ML�����Kx�`�M�Dd?'>�ڻl�=�q~�$Rfq����|_cq���!���+TǱ�����&�p�ծA�pI�����u�XlxVHYEB     400     170�g���q�E��t��EL%�-�g��,�NQU>I>5�$+@���S�thY)kݩ�l���^#7s�JA�~ �A���|+�%�ߜdŬ�M7���w��ĕ�Y��g4^����'�8Mz󥓎�����$6�����K�0�{'����0��DDBhĐ*������"X�����
��>����y�x;����-�:�|��0=��]��Ĝꃠs�?�<���9g�#`Z����td�`�r,}�'�N�Ʉ�Ϡ JV
�0I��p� ��G�Y	}�n)�c�:���붺�䭜��(���'v��5d9~6��b5�p�O}en��R�0. ����&*��m��Jeo�V��t�XlxVHYEB     400     1f0�
2�hĄq�}� �)�h5�FV��Bk�Q������'�8����ͨ/Jk� HyT;h��RN�$5�=�Hv"Cc�y��(�PIjN��M�s@{6N8� �����m60e0��wMu ��6|+�2��M��31�9Da��$h[��¨	3������﨡!>�Eш�����1{����yr�%�r��q����H�͝s֓�=���������,Yq����^Iǽ����Ly�`"���0��t.L�q;��F��d�����Aр@Y��?�<�g��0��L�~3bi���,��b\������?�#�M�Fq�S`�s�{���K��g��A����N�	�з�tЀ�LǹW��[�SQ�R����(�U�:�]�)]ℨ�N- X�L�2�%�1��/��lU�Pq�:�q\p���Ŕh��(󚐚��������)�j_N�oj����\�/hvU/���K���\n?�gS$����M������Ηu�XlxVHYEB     400     130,�'��N�A��������~i|�
��'�-�W�3Lw�f~i9����Xo�oDnF������;��Y��N`���EZ�褿��I�ꭦ��I0�P��ꇉ�j�u4.�E�&��e��6�x����=Pz���.?�L��_ ߕ&��U��e��J� �)w��L���m�t�cc�-\yG|�z�^�T9����eP�<���|!�!�Hi����y�ħ�78xY*���FO[ͺ|�Ef`�r㓺���x����vH	.�g�r��),��?�SRN�p�(�䑛~�F.��y�=N/�`��XlxVHYEB     400     190�kď�L�[�J|a7���_��y�{�Q�)��I��L�D*��J-ᴫ��3�&����̋�:�����v?�08
���83�	����;�L�㴅T��I�IU�eV2P�1[�p�Bu���}ʻ߭c#�͠5��X���l�o��7��v�h����d�H�ƁN��'B/G*����WD���;W��	�{������61��V���d$(�I$>s����գ�[Ϡ�`���s��q��	Ք�͌=�!WH�gY	KN���K��U{�59x��UyC�v,v�v�Y�ϊ������բp���L��y��/�o�'`�!vB�Z��(�:�5y��"3���}*+3��� �d��
�����ԍU��w�6��g��Qvq�,a�c�f�XlxVHYEB     400     190� *��a�*�k
���W��n����t��+����zLS�ϟ�=��P/F���P"�M��6�̺{<�G�Cn���	mq%m��_tʄj���-N��y�����pUBm��1<�G�f�ޑg�L=��ê�'���w����(��R�Qw��3
uє� �Q���Rb����(�s��6�V�ua9 ������QQ<�ZaTSAr(��$ ;򤀵�g	���B:�!�&;�< X��,�����7�O?���@�X͇�4�/��}�n~����諡����}R�;,�Z�fo�4�R�_K5��D"�����Yݗ E������
�߅�?y�71sL�%a�y����
A(4%>��f5�~w~<�05	��}��=[qjn�XlxVHYEB     400     120d��?�.��#���h�k۰��H�G#P@�m{X���K��W5��Cj�������#�]s?�q�CtZP�Er��u�M`^)�F�ie��x� \���e��\�@I�3��%٬@�N�"9a��=H��˚T����-�����^^��Y�����e	7�`�W!����RC[���1�wN��dŮ�)T��eH'��b��sA/ou���^��۩��֟qm�M d���6z�i$S�EA�R ������fQ� �8� �����.w�Z�ZXlxVHYEB     400     170�t߷��6y��o�I7# �U��瑹~���be�
�T Wpw�	_����X�Ɍ� ��Hs🹈E��6M�9�o�1�Hʧ���t���܌�vc�n�?����'��^�f�!?��ٱ��j�E���Q����40��8�*x��`�/Vr�c��f��y��)�j�!�ؤ�;�3W��ۙ�j�f�G����#�,�Eպ�n���{r��4��Bq�e�	؍eeo�B�T���������Tq�ͪ�V���������j�S^�.��Ǵ�&��[7
+�+1��$�i�X(�ǭz����S%�nq��FX��qґgw>s�d�yn�FLA�S��P @j{֩+[:qXlxVHYEB     400     170�}c�wS�-�����j���N4����],���-Q�?R+0b��� ��76���I�6}B��wpT�r8�yfݫu��/L��0�z�W&k(.��b%Ujo�V�G�NlF��0{y�ketW�7gJ��
��Kjt�n��>i���Sʗ����r��,1E�+��`S*'���H��[C�J���[����Ł�e��A�	��]�h~���&o]/�ښ�Yy��WVK�v�h�@�)�2���3qr:�	S��u��C���ޑ �Rń�M
ˌ�C���=S�Dd�uOK:��	{��߼����(h{�ӡ�A �e��Jn{��l|&�p�,\��@��,+��h��B_��}���XlxVHYEB     400     180.䐈
Ⱦ���w*cIB����
6\�����X^߿�'�K>���-8����#ߕL����o��Hj�ቴp/�9Ԭ���F��N��ǐ���$��+BӅѫ�0 ��F�O�09�L�Q�ja�l<@��g�4ݢv՜�E��OT�V���h� �:B��Ş��콋d�z�1t���r�~�Qǫ�����?����xG��x�˕��d�G�	���r�W[-Ҥz��۵N`o�(VH��r<�e��lQc��hR�Ҷ���u�9f�ZJ���Ck� ��PCT+8���!�B�ʭ�́�RR�Y&�s��N��.�-��~��HĶ���4�Ȣ_��w6J�\��a_ix^�O����={'��3���������y�SXlxVHYEB     400     100ޓp���"K���S���"�ω���.K�l�!�|���!=a"��wq�l�O4 ��h���ߋlS~�<ۦr2�-����`1�e�:	0c\���֪�BЏāR6W��OmӇ�w���S�Cәb���]�'����ϟ����'WR�&tdr����Y�䛂���y�����Bp\y�˛l�bd���J`H4�>o/�=,��v��%�b�<&ӫ�HK���4����N��<�sN�+>�]��,DXlxVHYEB     400     150�Eg���(g!�F�!�K���WڙCʳ࿔��#�
|!)�z��c�� u���v#@5���t��]���J埌��oz�C�Gz���Yyȋ�=�����ٛb>y�I�X�ph�v��I[��;��2�Y�P�	R�`���d���TEt:S�	�1�T��i��q�"�L0�\�=~���$w�4�t�t�ʁr��ܤ�9�l7��Cpj�H{��!�pq8��RBY���Y�;d:���,�ep�p�H��G{E��vȗ3�%�.�*Xn�Vg�Y=R���"�CXZN:�^��>q��D��`���������<̆�jY g#�`}jXlxVHYEB     400     150Q�W5���HXسu���O\��%t���L&za��8F"������������hOM��Q?#�`k	x���\̀{���g���#(��b�
'���I� ��4�HK}�ټ�E��n�Na�����,T,�J���ݜipV�~M?#�e��T���]��g�C���re$�︁3����~/��R���UP��k`ls���/+wf���*amu\/�G!1cؓU��1X��dO�F�m�t�K���)1�W V&�-v��e��a���"a�B��3��9pʍw�4I΋��ȋ�F���%���A�f�8j�㩞�|�{[��q�ј���ݙ�3d�)��XlxVHYEB     400     150�E?�p��s��2��ti��}�7�N����G��.Vz���J�\�v��lM|6X�Tཨ���K�2!%��l�
]�Dd�R�DrĨ�6���떢��Y5!�ץ��i���.;t_yWb��A���'过h�U��'Z�Q<`sV�����ץ��d����L���OJCfb4[2��
��N�أWB&� ��3�-�X!��oeA&��@���>উr>��"|��h�����t4$	��K����~LJ:z`I��2���h�xBt]�[I�єȰa3��)@X������`�o��č���3pF��T>�'�&�U�pG�J����P_��nXlxVHYEB     400     180�)���W��	�]F��E��n��T)�@����.:qx6�NG��`v���l��Էk��8�(�et��bH<ܳ$0g���[��E�: ��܍(�<ۘх� ���M��|W�l���ߎE���aW��#P�xz�LE�ɑ���i�J-٧(���,;S]��O�.ҏ��BfKؤ�@(��� X>,�PO"��������G���� Dk�hW:���N�s��|�� w 2�+�f���rd�F\o�+�W�d?<G���~�_�CI��]8 Ƕ��@���v��N����q���b��c�O��V�����˧l�E��B���H�uw�{���e_��xO�/��J��m����p¬*]�<��)��8O��K�}XlxVHYEB     400     160b��ҡ��u�����ݷڎ��F�FG8�?�6��g��"��C��Hn���	u�k���<��E�?l��KԢ��B(����Ag���LK +M��ݳ!�z��%_=�N�̫Z)1ɮ=�]����#�G-����c2(K��������g�feб"��`��U	���4(/襼?�D��b�QK�.Ŝ5^�m�GJ��w�S��"��-xr�G��eV�&y�<��o��1g��26t�>�Bh�qX���'�?m$P���V<��K6�X��>�p��v��A$ A]�kd�	����:��c����j��u�Z.�E$=�4�:,xܣ��:��7?�h}�6 ^XlxVHYEB     400     1a0}!-����rB��/�������������c%�������n���a����W�u5;��`F#O�B'�)���H,�O��L��Z��6� o��]�kG�O
D-��l�.�Qc�$>�l놷>�Qg.�X.|�A�rIb�?��o?Z��KZJh��[�������H.�]3�%f��O�3s�ҙ٪�.��� �R��!ux8��E	L��4HM�,���j�r�<�,����ɜT�[���4�Ȼ�`\p;���\	r�$���F`o 9�����ԩ��AI�ȓ$g�hǤ��+�l�")OW��,Jo����̲mA�~WI41�uzBST���&�u��}����:ڣ���y(�T�Ǩ&!��q{��5)z���E�7E��2:����Fj����,�xE�m&���XlxVHYEB     400     1f0�>��yޝ�����_���`qq�l&�Tv�\����|(��h%�d�l��W����}aN6��H�dRZw�[߃(�ǅO\X�VM>M*L����q�.�ĥЩ�7~<�%�.�����r�y
l���������:K�F|�����]\��h��X�X?M#����0���\���^Ų�����Z���t�Oﬦ|��0|=FU3��
B,�����q�p���E|BOvrLH���8��]��[ݙ�H��R}	�i+�� ��*�1�wY�h�ԯ�Q?���ߔ1�x<I}���\�nl#��>�J	X;���.��a@�>��#s��K��)�	�x�{�U���,B`$%��ټ	���M&:w鬥z�#i/�X�b!,a�?
F{j�#�������Bx�*�ŭ��5!�Α�'���oY�J\��o��F����`��<������E�#�v��j(g���٪����D+%i!���K�]K�tțXlxVHYEB     400     140�b%�)x�;۱u���Hy,Iz��]Si��q�~��
�5�F�>�\A��A�]ݶ��g�0�Qu��|;n=p���TA�h����KmZEe:�n?���wޒ�K��W-C[=�k�.b�T�0n�����	H�.��x[���}��1'�Ġ.����3GF�����>�
EG�����
�ːgt<,��;bNo>�G(��h#$uvA�����VY�%G20�0�Y�z93�Tp���j�^��(zG$����Q��5�HZ�C9u�V��Y�;�;����F���b����Ts=@��3�G��@XlxVHYEB     400     140%��VI;dkq�݆@4����B�� d��P;���k��g���Y櫅m�R�u���DyѢ��ּN��^����[R�8�p��<�1�:�2�)٩���?Lz�Z:�p2����f,�ԙ{KU�85��Ŝr�)O�B�m��X�>�����n��i9�ӠJ���A�#���ix�z���êN�N�7S�F�>�,4��[���jW���v�!���5��.�,u���,Ad|������8���Z�U@:A���H�*.K9�}�^�*�[�w��j�����-��@�V�$?vʢ�9�+~Z�@���XlxVHYEB     400     1e0����#c�7.2A��(f=Y�:�Ԙu�U�8U�pe	 #T�o=�U��<#�r�Fd���%�VP�1}��=U�����5�Z�L~w/�%�/X+�:f��[����M� �����̸�q�2�O��tR4
�ރϼan�R��K6c~�yH�0����K��o����?MLw]p���%оy��a��3����_ʇ�&0F���m>�{�xZ�j��u��	8RV`��Y��]������6����� y�gY�+J�7�Z3c���ϲ���4�KX|hQ��X�ш�V#rvy������=��Q���Y�9=��R��\v������dH�K��m2{ _i��=��	�J��f*`w���R�T��w}�DY!q.N*;f�`:A����	�J�$�Y��.1���5ܐ)�^��8^q�#��n��� ��_ K���!��5hEI�j�\D���U��I�2#{���A���~XlxVHYEB      90      90�<	�C����Z�M1���*'8+阒aI+Pk��\������R/N����=u~j��W�(�g�]��-Ύ�Ms�S�Dz��X�7XB	iQw�äk��~N�����9ƪ�2Y3� ���NU�b��~2��-_D�t��wU