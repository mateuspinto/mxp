XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��nfoUg'g'�8���ڟ�|�e�	�U��N]��z���ᩲ(2����/P�����NM#�=]7>��<�Jk����G�̋j�]�-��9Q�6�^�
X��[����k0a����ww�.����2m������i�O�NLp?t�v�J��
�2�>Ə��7�L���er�|>�F�KF���0rw�>�`��Fڹ����`+ϱ��{w�X�ֳ�s��!��L�Z��Uَ�ن��%l��W@I��3az���$*��#�; �P��'�ӥp�	��l��`U��'Q��
��-�Sd^V�t���c	Z�XS��HVw��F��;y���M��N�z����Tؚ˹��)j\׆���C����h�6�b+�^�}7�mvl��ZG	��\j6���/�杓�I����eo1-R��6 �)"�~��W'H����>5�e�2`����#( ���O �+8Vc�f
��K�Hq��k�u����-�X:��~.Ȉ���� �$E���f��0�R�y!`I��@R&՜����b.9H.Y�o<&@`�Y�>��,�]�	.L�h�ޘ?ӻ��8��(��&Hڇ�����m��.�w"�"�yse��6汊�j�8h�n��:1U, p���uע�n����,V��8a�[����vU��AM픮�@q�����O֚�FTg�}�& I+�4Dؾ������C��d�`,��{���ɾ�Hpm�����
�*���f��ηN�{��+�XlxVHYEB     400     1a0[���� �EϦ��Z_	-��I#\���ȩʽ7�R��'��{)v��?s;SV�]�#�<�d.��T�NO1�*eh�rƸ[�s��t�F����� �	BR�Y5�F Bg�~^���RH	� �y���wW/�ms���$�X4�Ў �k2o�� �:8귈s��@A ~��������@�~�/��I��=N$_2���54~Llj���S,]Q�D8i>�ȕA2G��L$'�����M�"��y��f�����~Ձ��=N��4 ���� x󠳠;���O9���P�Tt�=�.�&-v����]�g��3�~4���x�����#8�Y�g(�pN%2p�&Q=2�ZT�}�������>x���(�)S+�<0��Dy>�C��<�W��qs�gfҚ�8j���Z�$�i�2�m�jQ�XlxVHYEB     400      f0�n�E=ά�'e�q-*K��I����m�h�X}m���^C�M~����r���$�����׫��䑕���}%y$9	A"���R�5��6���0ѭ�0�Mj��ε�)���W�w�]��K`���P<_�J��u�$_��uk�í8�w��T�Vl�zNV��w�=��c�F��o.�� �߷�PQo�O<�R�w�ib�u[����w��e2(nmz��j���.��P_�3��K�BXlxVHYEB     400     180йhE2��E�	1�W�����~����d#+^+f�b���d���~���or��#V&K���t�w<���W(V:T��~ |e��酿��c���Q�a��-E���b+��,^���$YA��ݩ���fI���(,�$k���w?7����V�hQ ^��0����e��q��AJ���x��0��4�A��O�>Ӟu�v7�o&���,P'	+���ۿ�xC���_���=U�eP�q�V47�d3R�d|ɦ<fh����&����f���;�9V�z]�H�}�ʜӏ�
����8�����Pjl���8Z�` �2���/9U�ZT�F��oC�T@X���Z%-K��>F\�u+����x|����j*�)r	 ,r��XlxVHYEB     400     230���)g��H�N{E^��S���;��A��gJ���JY�c�Ws�w� ���Bd������i���b�Y6��7��th �G(`3 J
��H4����T�7�5Z����)��Aj�L����!������M��.0��S�4v�j�	��^��@hR�f�e;�/��1=�:�
P�1�/����j�l�D2e��.����񼀁�o���6�H��s�/`^`�M B":S&� �oA��ر�6��	�D��0���E��t�u]pM���0��*��r�����Ë��Y �bYb���,=�g��:��W�`,��x�� �D��ޑ���h9������]k�<!�(�P��:[��� ������d�q��i�����=R�WB��4�����`�`�r�(���h�%�%��lZ�[�������1L ��D�X���m���W(MrH�h�_��x�VDC�[U3���vH�&=�w[3�>��,��5��O�3)����ᕾ�{��L��Z�V���	���\��F!!^�KV�Jd�@>����pOÇ1p��XlxVHYEB     400     1c0�d���wG��T{��aX�2F(7N�J*]��uַ1E�e�A(������h����Y5%K�6ƞ}�R�yk󑌏��y���D$���ѭ���\��=b*K��t����m��Z��� ����>�Z�LIU�������h�f��{�e_Ri�7!#i�F6�
����7�{�셱���9%av����76�;w�Y�d,��r�[��p��<r��L	�%B�>�@�Q渪)�[��x���*����2
3S^�~��ES&w\��S���԰ �i����E ���υ�e�����b�g��.�s_�'��V̋����@q�u�q{�0BNrpha�y�͎��Y����35~q�V
�YI�ٯ&�?�c�R��[o?���Y����'�J��6s�IF��9q��A�sj�irhf�k�u�[���l0� nXlxVHYEB     400     1a0g�?�	�N\pk32�Y��Q�,�F��HѴz�Y������j� ��Z���\�x��P{^�^u�$(��K� �bA����iVqD��rAM�|� e��'S���;�x�_`x����[�W�%�e-�r<'��)B��������I
�KYN���x�7����ӧ�KR�A���bYj�5QtV}T��=-��z�%)�Oq�	<�w2��5�F���]m���!�%�R6Gom��h�M�}]�
�)Nԙ r��u��)�%G�0���u[?į?����E8���G�]��D��[�t+��lq�6�ߐ�O���b��gw>�<�Zg�u浻�𳚱�Dd�i�2=��½]��$�'a�y�ʶY�{l��r�6�0T�P�%H<=u�r$_�ۄ���M�x%�1R�D���eA��ZXlxVHYEB     400     1a0�
-��:���n�+)��y��?��Լ�>�;��"�_OB��\�P�y�+�1>�!������=3N&��n�(R��ix�*�nz�9�+�Hfy�y�ĵk�3�z���f�
���8Is��]���J	I�F��}���xR�sX1�-?�����dU�״r&/n�����!Q?w��w3���k��"�H��S�A4�<^ψ_�����T � ��<��R�"��l��)���aQ�</���s�k �.�I�Ż����t�!o�0i�cj��M��iBEa��ܝ!xGѭώ�ASF�mD����$�����ĸs��\�z����μ�B}�T����;���q�y=?���F�eo�]�w�r�H��Ncc{7���jc�5o��W��C�����,*�˽=��XlxVHYEB     400     1b0C�����a�wzX�!��$Q}��:�K�bh٦��� �2핬#�w�CK"���thgHK�rg`UB�ǵ'lim��r�x/�<(�۰c�iN�;�����=�q���o�Wu�#o�_x|?K�#ow��RM�'X��mc������FYGm��Z9v�m��2��y�@�K�G�7����i}*����uU�� ��%OȬ��E�=��!�s�s6x�n�Sҙ�BzW��.���׋ˡ"z&\�Yy��<QbE䌫�!n��%G�(�~�c�"\�_�/�`�c�*�D���h��������?�U²2��>����Ώb�Y�6sL!���N���,=,��]#1�]�0?bty<x �x�����{�_J����p��ʐb��ڨcH\���E�,3�	1�d�5j�XlxVHYEB     400     1e0)�=��3���\&�6÷�A����639k�J�����9�s#
Qp�NݏK� �OUÅ�m���8(�1�"�-IY
	GpQ4�!��Y��[6� r:K �M��W���jN���p �������7��Y���ӭ��op6z?����7�9��\�Z'ѥ��TBFή����	͙N!q:��7��s�H��etw�a�/'V���h�*���<�3��O�G��
d@xM��ᬞ_���Ŭ$�f�U�6�A{ei�[dI{؟�b ���������	��i��3�. Ւ-5�^4y��31�-���3"/��h�C�&2	oЭq�A9��(�~ipIq�A�k�CQ�:c�,S��ST��k��n[Q�#Ѩ��W��3ھJ����Q��u���sP=e��g��Li��Fr�|������[A����*�ߴ<���)`_���I���7Đ3i;אc� J����2��XlxVHYEB     400     170���!�q����G�77�I|Nރ����3f��f���#"�=9FA�*:�B�%}T�Ĵ��qd(���ۉ��	|B2��1� &�Os;�;�S{k��e����Ii��}��v��R�"�Ό���bؖ��D8��,e�`�s/�>0ަ��DԦÖ��Y"�=}�7q:}�%`�O��v[���+��[�l�׼���Z�C$v�{���lYx�l����Y���P�"���=h������;E���@ߗՓ�'�lA�RO6« �Q1�I,���p�ѡ1�5�/��m��=���>W�r���Z�Y<��M�gKM}+z\NFm�|��pw��i8������������0Ý��g�9�
,XlxVHYEB     400     140��4_Q�As� 8�\���b�ML��U��s�]������md����+ }��o��S�O(�@�ׅ2�O���:Y
����V�K���nГ��E���/��a�V�+��G	��J��^G#�gk�
�J�aF5���z{��Yyxl#��Ժ��H�m¼s�[;�5
�����#��Eƣx
le��/�F�?�c�c����o�����
��ʑ�G���L�aV��(OH�	���������쭵�^�Y
=�0a�7��fM�+7�l�M3(�ͦ�ޤ�:?,ɨD~��`�x��]�P��d�	[%XlxVHYEB     400     140�)�o؃���+>�S�Q�;s!U���Nc�x
�VZQJ��U�H��+�Όe����]k-��	�r��=1"���nzbD�
���}�'�.�
8&c[�'�|��qMCp����aB�)����	�)�Ãt�#�fp�����G�I	����XV�z��S���C�$�u��B��C��f J`U [����"�~��1q�<���kEq�����i��8^Y���4�RB�+���?]�w)�~G���/M��$���yޞ�C��[����-�A��^��Q�B�����.A������}XlxVHYEB     400     180,��G�iO���_���ı���������8��&��ϼ%��a�U>�%�$f���Z;0}ej�D�[YXc�`B�W�ݬ�먷����L~�� �	�A��><��(Q�����ή�$��S��V��uga>�?�5m��~��1���'�S�����\�����1���ƽ.����e=}�2���a�{!p��ݹ��<��Օhn����3|hnrO�M�\~���D�^^Є4r��F(&���H�a��.Κ�;�퇷×W{J�=l^��'�~{s�a��-CB���wˍ��n��/#�������<�� �iXO?���0=Kx
�	x�ىԶ#%fm0<�A=[���5�+�R|˩�Z'�GQ�X�W,	��OZ�*^�"��鐎4-�zcXlxVHYEB     400     180Ae-�� ӡ���Z��>��|��R��&��!486U�a3��)�S ����"g�$�S��Z��k�E��F�gLL����n�;���0LŽ����ogbG#��0�H�/���/�����t�=OBt&Kt+��g�޼c��v��Q�}=O�/��յ�ne��f�#|{,]qK���]��nF���jz �R,�8M���I�E�9�+.R��	���z:$��y2��{��I�C,��R�
���5r����Fl��e��)L�=�`�m�'�k!W�M5#���v��NU�2���d�uyiHQ�#}��r\����ql�	ѧ��@�E	|5�te	���DG)Տ|��k�� (o2-�v�DSV�Z&-�	�R��k^$�iXlxVHYEB     400     180���['Z�n�P����MB�&
��������oۭ����7��5o���#��f���KKGY��!��<8lb�
50&cQ����CKiG����ZAJ)!�*3���g��������J�Wż}���Ɛ���o��+;R��il
K�d����X5\�c��ڔ@�����ܡ� ���u?�+�����-��T�1������i�
�d����Y�\�F|?jA�pB��C5aQC����X��b!�8b��?�:�w�5�/s֠��ZU��GP�q��zh�</Y4�������*���M�����_\�^�Î�L���\��N�s���2p��KQ5Ҥ͒Q��/�4�6s����?�D��V-y]BŮ�|['��L�XlxVHYEB     400     1a0��X�k;bN-�	�:&� 2D�bw�ҹ��y�-�y�g�.�~�B�&�FCy�Ϙ�}9����8���k,�y�� �5s���h"@��c�K��Z��?�Y+�̮�':tФ�����}���>C�ŃHUùu�F2Wh��A�1��9 ��u	F�'�yn�}��<�	q}�Q�մ��B83W&HM�RG�}+*�~6��G(����*�r�~8��R���F]���0��B��c�Uu�8ܥ�'���H�&�(�VP�d4H�L�W��g|�N&�1���%?��Zz��Y��E-vS�'����B��	[�:ڙb}#��;���#t��I�d�= ��9@�.��u���/ ����W�؅�!�$|l�\!��5��~?�R�A�)����R�i/Mfa������$*�>%�XlxVHYEB     400     1a0��Y-O�����Ҍ4rr�RU�:��g�AW��fC�<�G{���q�2������c�1���ύjC��#�|/E�؜u�P���W�ko�η�:��h�g�Q���j��;��m�u4��c�)a+ �5��d�[ˌq��F��� ���, �b����t�����,�<m��#o����/\�~?�<��tF�+�+(�Q?���.����T ��[su0D��z�vw���9�	�i�yu嬰�ǳk��������%F9�4��ip�^wY��]��T�)n)�ҭ���/�x굜1���z�[~� ��.�x\��ْӤq���9�`0�e�B�6U�q�.��E��L�J�Q�Y��2��M�Q]����~�g�7��7�xN�\���]�:���t�q�'A������hs�+�ݗ�3��n���XlxVHYEB     22d     110T �'a�Љ�A�21V���T�^����OOO{N<>�[^5?HH�d�h����<��~�Sh Z���������*��^߸<�h�2�]dp���8���0��9��{$W��4x�pN<����^��E�7��R���dT��Qx��b�T(�S/0H����R`����]���X�Gn G,�g�v5����y�m1�DQ�mD|G2��Y�}O甚����U-"ٔ�UmE����1T6¬
��sFb\���4@BS rw[����Ǵ�2Z]���