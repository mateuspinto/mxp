`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
J1N3lvaLyLKoQkhGqh+d+NrtA4/m5Il5oMUd7RzR84WVoKo1GAQ01zXaDud4+jzmPhd6M2+yxfdd
0AojNXyr/OKydGI1OMBWCJkxvLkdPGFv/JKY3GB4J1Rtb0/dGg30Q0l9oFmmLN+MFpcdN3hS9DBs
BN7wGgtLtES0BZasJJT6xJsZl/L+zw4uSFxuh1KlufLwOib3tuXYtp3NaZAQjVJ/KaeaMLmlIBXO
Up5/psMYxxgZA5vJYHZyenBz78iOnX/U+MXqELwjueiIEuD33MbCRA3alpASX5PFBZyyyCKNlMf2
1SkSwPIjIkca3vjBP68HTqD0mAsXOS9FYyDEKw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="m0DDLhZzPkxez0Yyc0BQ59U9nC/q16Ws+qjYL1rIrPo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 54576)
`protect data_block
5SqmbJcc6ijABeSVsY6kGaVUoeXVSvC0WZeaBOXAsZUnirr4INvw+irFBif4VrfOYc9PN1mHv2jL
VLEbaXuC0M1rCUyhu/PfnIPgs9BdvSdZiJV5pBs+W5YzXNDwmIUwRbsWEaP2jQ6ga25mwGQzmrxk
D48Do5Vnjt1+aXR9jJiZR20QNRXLWgJFG/3UWacnCjIdT2b7uXcAa3lTVX4m2rioDRWiC+n71R7z
8NkI9wdgq4URDEhO6jaex1F4sKcO+xJmHXxt6vu3TQjxR1s4hUej5lyG6O4+pEozSqZVIAiGqp40
kqABwh6bYBfRhZv20iQOZBYKZsA1KIBpwbD9pvR+kktKscu2QSojjGHYYJZvXfqcz81Bf/AOQliA
ADJGDpjFqIF4upkTyZsqZgkvf3tq1ymJn9HAc1bHA9OuFesS0XqKwernkdCvoFUP17pZRrL9CaNW
qv6TJNMXsnLWn+Imfg2GsKrdA2Tun7ToFmUISf4+FSCk3/m/RRzxEZnWzaQAOnm4IPeCGRu5kTcM
39RvXj3sN60VnuRBg+cNH1FP0Py66JxahuvbzjVDuFv8nTPY54d970m/K9Dt2xO7pKTLBYOeN9u1
YAu8RpdnVwbbfrIjvWcBv23gfN+g29milgazvuP0dTOMib9zwLqyGo7Ss2hHDI4d/0T+S+s1iT30
YRMvChbYvNE2QvuRYczmRM6rztaODphtlMZzVDr9dk3M/wpNQ/vwXN7I0X2/OMuY9gB97ajeCCHH
zcf0A4eSvKQb50uFhd3KI05uKYdbuI4QL/VgHd4zZyi2uNYl2PZr+vfH7rS7nMgGfFnfMLach7t7
SQauIAwH50QxKTYY8WSPPJuQ3oPmdFa4JUtVwOB8Z86YRzM8ibOctlf/qJ5c20IAK2gGB1qLwtEO
hiRhq1R/eRZ8pUBmpwzRWI5LyNXhh9l5UhRSw5TDfuxnlIVhILNiHpGQ0HgvTr+jlIACzqS1946v
wP5vEu/va5eyeOZPJhRUyXIKGLHQQKsl/mw4oH5abSJ7jHqE9TPPYa6Oe5T8NFwLOLcdIfh65gvp
+fFfWfAoxqfpby8kvrOxG0OXVKqIgLSDOuFl3AUso9gngvKWwXmB+jrEuwUz7ypHvhe0VXsgZyL+
5pvjXGPfnRRvcOzmyoEjuXvew+CfJhgaJyMEnfo77/RmTQs7BHoYgaI7FJRO/S6C+2SKMt7Ss282
J0wyg+QmEgf0p1NhsuGfwZIawF+Mu+I/9rcJpkxp2nSKVqzhs68SNBr7ipgW/8oMkLsVBFfxxxng
tgIlQjsSye3spmFf47J6qmu3/bh59ZzNo5zuMhamMPQXP5B0NAlF1/mqbnTUXGgJRd+vqcMj4kO8
N2TYb1VxbsgGpfDDjKj0CiKW/01mGG9Be12kIETxkpJtDOgpAoBGYiQGU7NUggad5a3SzmUgO55P
O4MoXKzM3cLluQ0ZGfC6K6vfc7XyTcBYQsuuPTlvKI8QWWdq/T8u12ntQ1inCLf497GguriNalSm
nawQ/WJKuCkUYF9zLYvYhYETncElIsqyu4VPpe2gSWEQ4VKe5NP1onOY3x7fE8UbMqeTkbirzwPz
uCGxA0t2tXnydgjjnUjLcr/AsFBtUqyZnx2EW8fc/pOBcFUWvH7R2xun979gF93tLAGmDsxbE1Qr
rw9iHWME7m1kLro229Kazj8dfCTaIU671010ocffCiUjvCbUjD+4iJqjnT6xyCO9tPJxHVex1+t8
5S6UDvyZWSnkgIHZmK4Orqe3GbTextmcS7DkbTUCwxi3ovsl4oKftNgQrI+IOzkXHrO/TVzR19w0
Lxz1x07g7kf7RNi4oJvq0zCcXTMrJoMfUreTfvanbrHrn2dFMP8K3e9fgbY7Pozebf78elPqh3k1
FQI2xn1KdXj/iGKBBPPwjf0xQ5O94c4RTyihdl7cwub8i83O2jSXkFiAqeG07+E8v2J4m2H0WuPj
yKYREDr0RofKqUV/EesapOIRN6NSik0aji9HmRp/gQ2hHhGXVBxBbX7Z78jPvaN6rI83r5DYx7Y3
J0uQHVC5tU2GNRstTiQEdnx0U5lfRopLWJUGhv1Z/9xfGyR7qbAx9fF38tqoa6Vq5746uZVO/ari
sktSPpXGgg7ghJph6NbbruD8pi8oUKgstu+tRivupxivAHBxr7KP5h5Se7zOEicCGbJA4g/IyT0R
yqkQxhNC+jCA7CKLSF1Q5cDh29eeRWzKImRwt+M7/R1SmmKII/Eq4Ek+Zt/aSf4iQkCXjCL9QhzE
Z4K2fcr2TNH9CrW6z1c2fPkNv4/eKpVMbnDmrURoqIRp/cS3qhdIXTs4PKcLrUVEQlTsj8RnmZ1Z
OOzBAlAUeX7j5RY49lGZQYQqXVjYX4ps9HJBDXlv/CeJwYiUasZU6Xz0/FdpTYEDJb308k8/Hogw
aNrKzvrKFsu5x057ip0sudM4ffUlmAU7FBIp+xpelZwJFnEq6gl3ha1D/Hedwa+JkEVTRDVG6WhQ
mXYdRDyf5mpfKHDNC8xeDBQEcErwouYftMd3crFve7yCEIkAmuGxGrAn9Yo9U9sIe6v/Qux8bSaJ
quHTuggj4vExKIukVdQ7iz/4X2Rj58nWZ3zSbzMVZx/cFzeElGMeyAP8eQmUshzD9Lxs7rOj6HNr
KVstP3sBAd3A4a6SqLU8tfWoa/yPF9Cl2GMzWv+lefFDosjPLXsOOo6lI6SziOXqXaUUVQvEBwVW
ErK43jgO2zd/5bdPagyi8DEVshjWuj4CckGzawAFweTdRNkWVBDG/qiFhJsfQnSza1tsyZ7XQFBS
RgqlZ6fK7DQbmfRI94W7Tt+oDq45ij4Vi1aUS0B7QUV2EDNGnQoA48GApQJhtDlYuAxN3B+rqqjl
HNeOIdMobt6fmgauOBhw8ievaok0oz4PrfzBABCjeJtFZ4BlDTqqeeqllHPXuB/oL7a/Yx6s2kFZ
cXQHj4kTbJ58Rudowx2zBnVEda+7hnAAO1RNFfnKZwCkmEVtCLLdtWaRXz098N41cla4bTqJhUD5
LLa5bbuvINxt1NKFWbXwd5kd27wn8NBi9+4cFApSaf0rsG/1sJODMzVv/ECKvwdQD4SU5fzpeTwv
zi9iWW/2CQH5/rlWsA8OLYhGemUmPWUOkvIhM5L0TkbcVFxXIJvPedplRKeTy8nzcS9Qdg8s70e/
DbqSWUdtczlvxiHzlxR8ooJAXetan+49D341v+/JJf53AwSOtTxbppH1st2Nhgeh/ILxy7k2holi
HXBLefQkltxuMWAOsZ+pMh+EUfqV7ZlxE6aIjBXzWsS9uQuCNqrp80k1ow9YRNSsOzFBirvXTW+0
3kcLriLlt9HWDVNPdX7o19Ech4w8WQMQB/U1ZHEKANC72seQuGlPPrT9mgFLBQpoY/zqAe95+ctt
BZDBwbc4SuJhvMYWXHemTQGlRuaPy3n6LYVg6hSpBfHRA1qp068jPekYfNpyJD1Sm89kv3ZPmk/e
JekWVCK8CQrtecT7xRaGdZjPzjQNP/t3V1YdhwivYN+YMiSSUZ40S/mMDtLuovtGKadMtMygLVkt
FnExykMAYE0fRSA44FNF2V+3wgWUQdiVQbTiDD5aWxguVZZronAKj/jtZqUwIV25CG8hdi6swJjI
t5BuZiQCTM0Tq23V/ZnocdMgfiyMFVTiATrKhS88tEqKi/OOQ8hwgHxjVgiN3TMwtWSqAW+ufVe4
nW1U8RZI733kjk68vSZ/PEN5XDK7fmSMO1uq3CD6RLU2vcTvYF6aBo1T4Ni25VJt6oKFwMgT0Yut
xymtTWA/unxHQi/Rjg3dtGqa/4D6jdb1NLHPW4R27Acn8HIXvFd16Svq6y/rJabTIkzv/f42AGI6
L/nttNVYCDANTUrjja55xIaxdqYkiPMXt6+sD5yFq5MLEv8tFQ/Y9uVEoRTSCH7M0s7NkwDLp/xj
40uq3iCEhZQ5JFfwv/r+bLiPQscqXcwkFGpQ1rAt9gtxGL/Aj3jfDeVAcZRK6mCy41YVfJSk/COo
WjfjEJjqFLOmYYO0HS8SnGYtPhfiDkmJr+pSl+jEdFsFJonCtGtv87udnbI4ddtxeEaSnYynVGx0
rGA4kSDX9nXWGsW3bY1pRfSbEQNfDokm9w/Mg8pzieSry8978hJCvQkCO88bFwSGdAMA7dopZ+no
ATsWE4UnnhHlNZJdWXqrMxJBptvdbgR7BbXiB5tNvM/ygOSt1OFwFGnVVyId/t28qPYIszjeJBz+
kXXabd1SBzLSMDwrjborrr7z42Cdid20aYKt9n8s/B5qijjoGVZiYllk9lpyJBhQSoHuvGrGAIt+
Go00hL7iPA+jVS8wBtHCmdT8q64bi/ulZJGXrDDMI0+9ztCV7qe/Xov+pTHRrOrvfEwQvpfAKTyG
zXUSvXDkoLgQ5AuTaDwfff5XEZCBLu5aTouA8IbzBSxVqVbzTM/0+5k40rzUAia7x+NxKGS+gWxG
Yz0Ck72TFSxmkEgaK59NZiEqXflQc8fPSJEEGtqCOYlLST6YawGG38Ptibudd3aSA1CEA58jROd9
ZHGFK6KCPg2KCFT0pxcYLOCDzuK0H5vXhvotMCEa64lG8IA6TnPS/ADpvy4i4OOS9R6ZcngLOdpN
d2C7MSldtUjYb3m4mXtNd7gWj1HFhs80oE8XDTdKri2Ec6Qmf24BO5zXfeLXeQ0zwcGFPUEW5x4n
7UI7aIB7waYYqhh+bb5usfc3/ttf7vtOht54bz+63YLEa5+RoSAlbmoqPQtPqw8lMqzrzKKDrMU/
ek1DhR7c1Wtq8GMKb4zmIV6IzWTakc/+I1tg10jfeOtuiQCuGBATSnoDxAwnyygEQY4x0lP+hKko
KRRdw1Ea0xBwidyAh7uysV/mh+T/yRewYAqJ5gP0WCf5dTfRO7fxc9ASOnN0EA5B5pfr8b+w1ks9
YGKZ05HdoVToNplEdPFrflyomrVhdhhIjseKVz6yseR6NORVxwR4yd6pWzeLUIqgTOs3ICpG4HQ/
crWkMqV8MPAAz6CGjK5UVgjpGTlePbs2aP78i2PGh5L0Pa3FFAFLAxYU+DOwZUVO+FhpxiKVdVfh
xu4Qjluf0c293JFuQevfU4TcIBaaZ3XoR6YsXRcOSrE1uwy55pDXSshAXPuvmG/bT9njdCYWh7Z7
lW6rjIUZcTwhiQ+5jqU3rqYkilAxMoSy/8u9qZmtWtpqb4kLde4Zin83ev8fo9LfIupRu667o0py
r5C6HvZ50hrR4yIeqVd+mIhfOOyoCzGlzywG80RTCm2ybK5LJy0sxkOaoyQZsqa16ARdTDGs5Q4W
Y0qvGKjkBzWANGI/k+2kRfHFby6CSgnnZknIFuKgOAY+EGD4bdBJGv2CB2fakn7IOXirF9H6d9fP
ru+T1RRX76Q2xZAY+PhyBJ+9ioS5yX02jel1kbunAvUH76u48Y22qglMXscOSRh8JfODfSZmwoNN
um6reaLzJWnIUCTtcWb1NJJfVzZky1tbiBHmWVvr9JDef5cO0DJrtYBk0vmTRrSl1wtoyx6NrohU
Hh7Ug025gnuISFSF/V59lHqxOVPTkDTS64oCTSgtbqaK7G4p8DM7cSJ4iAw2laoNEsnAlVMmTLWa
A5xpklC4LeIwYijcCLTablD83X/2dO+0KQRUXv2LPHPNXJH/ydyUpIYHwOA8VBDKDgn9daSLTH7B
GMSyXvtztZc6SiEUaINQC6lyvd/bIWr0I5jZXija3Y3pdwvZEfeiqQBJ0Ph7tfF/uBgD0h8tNXd+
A6QKtvanOouT8wFLFK7+Us6vqhqNh+j9UdYL53sgSummT9PCqcvHGfou0yZqtj23MUCbljjUwxwY
Gc4qhojpzXUImBByzh5/dqDiFAlZ8SihbLbCZanBQ9LXOh+yOLQySLEudCwBxzTvKjqwpqMExqRE
MGJCjhANjslKAM4PY073Caj6ezaXn3rwte3NC5Bs9e58Y96IvM6fLqUcIJicXnn+zvySBQ96U06F
DPw2M1y8LQDu6787FPiTLxlmjGVNH/R0ChtDEqObrHAKHgt4ZD5Eu4pLzT6ssxkwMZfCXfkt/pu3
tij5ytLeNHxrIJhfpc/1jixO5NVSj6V9aCbXNK/HsJQ8AlM/MVajw6ZOCI8XRD/2+eWwp070AhwO
TzhX9ZF1AlOb7UvuDx+ZMXZ8rohnQC3DvlKe2rSW84rV7GAlOeIIC0rB1Sle1+lKq3umAgT5mEjE
D4Xx2xWUb8zCe4Qqyn6T89rSmTMVkCQbTBCp7oOFZVtAmC+SWjQAfVHv28AXognZnn4ekD1An4oj
rlTLx4jAbSOXOR70O5OBYthpKxNHpGEH8nZN0+pglFrc7EKzPbOrwIMZAhzIE6TnOEng+QUCPoBH
GwBRal2CAJQLxTF21BxjjKMhv8ChV5B70rTgy25C3C2KqhDWq/wLNszkVUZMLBk+ovd9Q6xVyO2l
jOORyVhjrBs8kK9o3KPZOBideoy1D3A+AnzH6tjSzxlqx2CiUh4XKkLQ0En14ivJKsx18zDp04Fz
hxm1TjtBfb6YmSQ59ReUvhu6LclPY8R2QpWp6JJO2AmsD4yVhjb0bIku/GD83S8cRgn7+DhLqNgl
Aks8OVS3QKnntOqWwtznp1gnN1uOnBBsdUttX8vbPhToUvXLfqR7x7LawSp+7VHuwSEp8CEOLeX8
veMQcPLaZkGY5KBxz9/Mkd+r9L7Ye/FsCApC5oB+7zKnRxXUJdFkJ2Ig3GxjFblbDuL/2dJVrOlQ
NwsrhOUMlixC6tDVrNLi85GZrfDY8SMk2i9P2h9J6kv2g3+Baf9G3JXhRzGLVTaYHx0I4/9YXNjn
WYcfR5guLJLHvoq1rC9mRCvZkikWcb7HUkvZN0nSozLddtXcPYAV6fWqkosyw4XH+Vt3TwsArJVn
O9ZCvD7D51oiyOL3qrKuPwlf/gAZzPkm/bRmA4YPeukCFRfxExYbkVygZRwzBCJk0/0fPvR3BCrb
29TAddlQxvwVGn/He2R/Zv9revCKxEcW5fsu9rIxaxMUVQSsAx2zaJQRa/8BSzXtbLfXkCWQjP3E
711yXIZfShO4u/HIQIN11CJ4iYtGVYnI9ErBZVuXH92keOmOqrXtDxlNcPpuCx3CinRgeLPUvPOc
Xt8Fo6u1IuKcKErfmdEHuL+9EdjhtbapiaD3nxmM3ezsdtea257Q0MtR2gbYKfhhZopkzl2wF8R7
9tHUXRwp4QpUjIt9a+Q0db6QuGUCNCibsSp/1YJohkQueuXz+fGL7/yxBm9u0QUOXxfNax/6reyd
LhpixmxJVvsSfu1+FxRbAYcGwduC4hkB5XNBPuhztVwhHK2eo1/PCrncaMxXZ9k5MDw1f8t7hcv1
BLhGz9Z6IXtQlQ5foSYNtzFlpHBYL0jDJPmrztpV81t7Typ+v3nbLSl7zWkl4KzCtznW4WRuR7PP
w3zFrswu3NYtK+qFXbkccDjp+FHUAvEBOQwrRmH/0DvsELsolKVKD1AL46u0zqAs5WN0A4NZmors
VuD52a4dOr+X9qyqMcWxhoe1zTf+iWGRCeODWOldvqRbUwB3ZXL7P7jN6iYeZ2EyiKMFcvhMx6nF
1obWYzv9zjYw4u6rAO3SRQDi5nSeDV8l9/YOfwhsaCB+nGW7almrjfpFwYjrRy7sfb6eUp/5tm6z
7jte+zjAluQ7WLBaF+jtqRbeqVm1bzjxTMT6n+GCONdiFejmvQcb8LCpIVwXOuhwi3SnoJkhwmJK
fCUKzh/a2UOnf+mzgZoOCQZZBlNHe9IM1srWeHTQNEZHW0/EjT4D/BqJAjPhnBd++tIbfb78HK5G
3MyPA2/9XazIou4n5nOD5B5Jnf0rtAzy57TFQzE6PIvLH3wiuCG0/XfzMESKhkm5WHZ4VU4JRAy/
CZcmPXlcYoh5FnJRNoQyYJtYef1j26bpGXdqK4Gpmov8ZO793Cz+YVJCFjNWI4PtgGnD4re8Nt9a
WpAQHeuem1Px4P2ymjniy5V/nzPGYbepfEtqT6Z4i/6iA6rD76EMpQp34E8M8dnc7hJVeJv/E9gh
xdCeLXHDNn5R3jWaRCe7fU5jRK4v6Pp+FkafVGeUvtGrtsumK5wNIafubNFCJSyPXNs+gd9m9KlN
4GCVEty7JRtFRmvbzi2vIZsQ3ca0un2TYuI6nmZnE+AE7LZKfPbh4BfO4AWWjzLOZHxOkai3VdJC
yGhA3G54llHSGLa4tDbJwpZILCQu/h455qlTVCIRg18KLRZMqY746H5K6E/zuws6RRAs3p9nM63h
j8UnV0PkFxhX/npxtfc2pLkYum8JKqSp5Ys94n8dX1UIpJJNfAeJYkuig1+NeQ9xlSWtkdG1wOuG
b0PEGGataVKiw1Inc6giUc9suWuGYbcBB9Zfp8ez8CF4GMc6k76ZDQvf/tHn5iKP0Okh16u02Hwg
4gG/GwFmsFMdJ00JggNzXA+jWWyPgn5Jt0RRc7oUX43lkhxwbdrN9TCwfD84BPzuJXsHI0X2sodW
ZMTsIm5Hbs2Fa2534YdGH/I8AkkfaSWrZVWLbGv0edfLZquTvc5nGdJo8XTxJ5O+zPSHWBsqBl86
D8TyPgRQ38rHLYCTL+1DgVfKGS962UizmmBTbnA0U5qmjqhmukXu16Dk+N0ecCo1/xq/bs+lgrkB
UPx2/9r2K9srLsxmc/izQZJDEiB+tI/u+vS+Dg53RQb9R6ZNoDldHNeeceYTT6/NzVGkCJmL1U4K
lxvfCodDYTFIKg3qte8XE/lxYU3unKw/O4fJnRqMjlmb7ueGLWg5PKxXIB3PO2lIwqtl40Gr4jv0
Rw4IaH7aFe6cPVS7Xls5xAJLmBm3v2geH3LIC7RrrzA8BhnhmeP8iCoxncHXubPTYLPh+t1P7kcP
eBIfngvvLloADdgdden4mvipEaSE1vTIPKxEANrT8C2KC5XQNqKxsIwj3W9TFxQut/sAJu6g9A+Y
Ua0uCC8Vfzz7eyj6SHKvDaL15mqVBrOevlkeW7BPRAN3IquhSZyNMT8Yxs4FAJ1TDcKot0bkkTh0
4K0Htnu80p4JE4pN2mRJB0QrRYI+zXTOBhi4b8qXsH9u+0wuW6Q3eOvfftRqLnNb4oZAghsHI7Q/
DB5ru6tuUkqvZRaNas6kXmOYA0iGjGVoGhN5F+jUBdps+J/0aw0u44Ga+uGy0oa4pgs3JzaSYNdj
s1KXfIy93Dp5aTwK7yNn+f9fX0PYei5BkVXnd/kFAGz+RQtjQXWYdYws9Qco5/4PVgA/32GGIjdE
mbphBKD22y5AqCzUxklW8aWJ56eqfDH0Ia+nn76gTLnXWjNsvP/67htZqHQEGLceOEyaQJ6iMZKh
i3aS9aQzdi4mBcsO3mqhMl3ML3ZM1GnlxUtaD1O6j7MMG4cnIjiRkd5pH8jDQ3w/5anJMjdzP2Hz
hk4ruuBxqhTu3xTQNuGnG20ES5U/95bSTIxNuG3a0jfzgA8dKUuuJWHNGA7zVMv/4yb0XsEtd1rp
AEYVdnYGMwcCXWa2j2pKT2MxIEF/8Qk8F03gNNABhPcj6SuvI8cJdWbshqRzs8ZJTeLSY8wcfKmV
GGJ6BSEuq8XLEFZGfEA203CJ/TiSsQdbvAgwdyL9cHo9HvOHVYRQPcYEiANGYDZdF+Kxg6TyTykz
ZZXIRwPDsTOdLQXcqQ/PL2wlOsnjX1B99G+7mDILLxcn5gUOBW8WP2P9eOe1pTqEmprZ54BgxW8w
JpQgJTzpiCNP3W2z+RNB65vciG3b9iedU6cxkW5So0RsAw79+Qu7HIAKPHRCjbkuYKQmyJ/0Qsx6
ct2o/ztEYdGIxarcBt47C4Tv73io0+wwe0MnZ8W015NuJinIeXwEWjoNnRk0BehdtSf/4RFY8zuB
okH+lb+1rSxpsdLg4N65HJffUxj4X3TVGp0vWlwBbj2s9hfcxNe6DvW/QEbRAE1U7/NvG4G8QQZ3
TMqN9zjq35zIV2x4c/FAreD25vy9+fNY5M4a8ScSriMV0TGCF19CZJKGhyytIKNSV8Cy/eYtDzC/
9FzEMr63LSena10B5ynsKwblRjM0+xfZHS61vAhhsIl+2KxxWweaAey20gI9q8LO0/FkeXY2gzzD
XOk0Oq/RgHk8OIscmzHXzxYDqifW8kVUXNGRp1tCH01Gl0AK4YupHlp2QscjRockms+FZ7o9PZzy
EDpBxwbx0Af5YdBM5Yh5DUnOh+8UNaePxEV6WE8CCFuTUnMXVJwKesfK6V9UYRtAcSVn/dibDTOI
4DUDA/VH29rN5c3bWGXlvJ022d6zjMDL9nFj1aw/wg49RtPav+stFSoC//4Jf/1hpLgp88qcqrOK
2CVb91C7yI4mNxicDJ0d9PPkA+Axk7Z4dlrlWPg5j9haUMEaK5AUhhDdVyUkEeLosmjsYh9FZD8b
LJkHifk6g5PNOVLBAHm97HWRCzWBgBEk/j5/V7WKUbzscHgjy4pCcFPEDsATNSdG3alFhbrZs2XG
6ssKYR+rp7w11DbgrQJGd4PNmvkl5tVvb68qGJ+zP3idXVUsjR92HhhEapocePEv8CG1R6fD6575
TrI8FCz3jcHgI6lmrK8xUVsUqdpw2Cdnep7bf4nLXta7+o+7iF2LYwIhwQg7MNQ7wUy3D+dp4LZJ
+Ubo9E6Dzz0VOdcY1F78zOxKU1nppmMHPkZ6dOy2qNIEAHmSwJI/Bwkk0tRd+rW9RU1wQEgSwxkL
DfrocSwKQNblgYGyR0mQTjM0jSKZ0asMIXMZy/CqvORztNt+KYIwVSN6HNLYs5dFRn6zbF8fBmFw
FCyCRuEgZU5rHQf7zUog46YUMTAAdm7r7dS34ECPAo4vwUgUUbqsMKD2ebIz/steoIEkNW207WX+
Mt3treHVkApXpQKZvyhxuq03mNHxu9kuRKFWdLcCrt1cfH0NsABB2YNq5HJ3tIwgAJzpNhD9maSR
1GOaM2z1zUO02hM968HmftmfOv188zrAesCPjSlzCBvDdoDAXMjVR90s8mip1r6tqbLXYbuPWRvj
TUY8DWJlQcyNwBrOL2xJjMLrwOj0goLNI0sop+xa/o2WuZJdpWjiclrPM0V1dhn9fMpTBkX3tTq7
EqCHdVSGRueLXcJ9bh/U0x5PElttYaNVICbqRdcgOZViDXeVLLu5Gx6VsM7shjVJ/Kfc+IHP95Mu
PcLWjR6SzLoAJCQ83yrDMqWJ93U6aSsyGtx4srD5DejBdbjG3GgYvVlrUlCJ5PnVIqn2vyBhStio
NSwjbOYwfR6QZ1KYgUxV9FtjQWxDy5qf5GNxA5Gv3Uy5Fbk934g0e0rdPwm3q2gdDicm8ClVD4ES
2y1R3ZmsmRI052PSFPPfO0EF8pVSWwxchyKwgeauktXtfFwWzntagWzXP80/M+/ve1aZuiYrexmG
vzDIP9aQlBzLp8cbIiMQmep2JZyH0elIAMYXA19IINtmvaizSScqPg86MFOQVOF2XnnE+yRoyDZn
G6VMw36YGe2kkUCnhLDJVvBEwMXL7ZeKfpBpEd7bJGfLBuMskyMFdBnklFicVkac8clK1X6UNyhO
cVWHZoJ5x9h19R3/S4jiuc0+3j9x4oL0uPpU2vhEeo4aav0eAPOX0fI/RBPfmYJmNOULidgxCokc
0ezQEGnOkCneQbZDRYujYuf+gphsVWSz0pnkMIGJ8qJGhsIs82szCkWnZiXtxgfLVi8UU4gaPdhv
r8ABup4hAmteKvGXbybldhuX9/u3GxREStGqoahHu9MhNAS2KRedQRJiDiKdt2GrQvpknNx/MTmW
xMBO0mKFHVZdPkR+/nZmINcCehcBHkb6NOJhZQJAZymyG2P9vxujthKpK5KJStlaVBhqDNVO8X/A
Zxg5OS/+TVJ9fSCleFnxDc10pcUHI9rMoHJBmfHUVd5IjThrFKhyx2ic6UocvkwuSZYRh8UlyL/b
I/Me0HuKpcvYJ/O2adTFU9OdgvQ78SBvSZSaTBS0iBqPi0CtWrSdkWgZQhaj6YtXqub+DlUShtV1
RN04a0Amair0ZWBGbb8RNHV5DRcOQ7+p/THPeUizh5hu6tn5/rNTXd+FyEpx2aJLvyf4tysc1wGP
Y87OOUku0rX8CxDtFk6X3TeFcdeic7tcEdCQTBCuFaDpneMa5hXFhN3gbk900zZPaC0O0t4Spsf7
wy1X9rJa5Ool3jiH8q611GM7JN67Vq0dboxO3ubQm0Bdo5werWeAIzWGO/Na/wlf+6H98V8WET/7
SFUTJQ+xqZoa/CnOeoD7mH02O9ggqJ4Vivmcky97XISQvl84SoVeOvfX6RyHCMz8+eyp3/aSadwk
Qy08auOEge8QDmFNQA+UWhViAj0kvyiVPYHaSiYw2e2QEdjbU8mBPojsQeS6VD9EY1CpjYsbGa91
505f7BqEJ0btd8gkPlB1vznvIlAl2ZWvgNLV8MUJxf1gwKF2dfTpiS6V8MQdeaKrkVJbrNyEqOLn
Wi6qjZCzf5AaaT5cn+L3lOHxmpuadltXzjxnVkloGWAS9M3XFfSr2El/mbAPqt+dDYaHWpCE4p/l
m0/2lk7aLMTiLt7RgFxBMMJCBADqRrrg44mCYqM5mpSlpQ6KwUy53iEfvtgXQBf114EsNCWeusbv
SWNHAh2CwpgzK9oApgSANq7TWqUzf7QfI9GTPp3y796OkFtNkR3mxUa+TguWiEQt/tQcLY2gLlI2
LTfFBt8CmofJk4aMHm4PdcZWggBVKlP/m44rmxmyLRVYWU1qRuPeeYTstpFRN7ZiEabW/RP72dnc
7RjJh8Teb6yw+Ht/4u7EywyXH34tdbmMhHTCrLVIYneizLTd4QMTqLf4UGb+oRzhMY8n5UcM5/Iw
mkOQrdZ4OEcQRLSV5JRJAWi7zS/m0jMUi4JxhwVCgNShJWE7NBA4iu8cY6Wb9ewyISomFzRx7VPt
lZS82naoXOn5It2lao8nfBClLCXTpgC7cto2R4I8S3ps6HtPkjq1QdYwtUzZ+14RY6+XOrYwY02d
Rk+nIxbBDTBdebAEn5JHcSvMaHOkFLRHPQwChwZcZywoFL/Jv/qiYSeNWT4L+umdRc1fD4iVfnzc
Z0rBfg2JgatRUbBXxn+pHIdHE0QFfqO9iWM4+lrNwbvSOET/uErq3e9DwC+X2edMC+gNAn805Z1V
dNZyKp3gD+iWHiEEp6ScmQHyNiLxiEyHS1sM+kh9j8tS//+Cibragkx72PtusVR8ZgbC/iRd3Tau
Bp+OpQelbSkyGVwndJI2PSKhLqIEn3bfS+XOM4mA9MZ3pyTmLfAqZn8Stqzgdw2Ck/5mUhqUcKFp
9HoVe//su3Oho1mwd+BoyZnAjo1z09rif5WZGlbbTNpMmZvUZMys3mgqd46G/MgnK87PeKy7Djd9
wuneELaKqf+AJIyr9496TsarA7Fn6HXvESdKXGooHBHxrJR1hKjUNEx5SY/V0U45jdpt1D+tKgpA
mWaFBJHy/6/BwA1fJKSOG3TfvYLcDIC3vHj6kKPpheLNpuPC5fRweF1e5aGAFb210MIglf3rXubd
8fr2zHUkTiNM6tewFKIR5Iqo+Ggw/JL7vkbbMme+1qIrorhRDptgD77qznq3vVULovM6jokzfqCC
IU+kL4KGK9hQgOknu3/f7Ns9kK5/3a0DPctLjvIs5OEDtJEWB8aqnGqxrPlrg/IPXoEmc+QEw0KQ
K7SNBgXpJcPmsoRxWKGGFhc+IS5Vx0ZIiSBhGAGSbYubnVGdU67Cb+fDfCr0aKyGXK2yf3FZkfgN
6ruQr7t5XlntL2YTRRyonogi4eulsyfVgxQqJM69CGSe3UI4JEwjNdm7NVklW6UMkAh2xVFgKU7f
+kieHNHBqPckU1F6lWGPR6O3ZjSYdNb2+xDy2p90qOnNfpxJzQ/WljYoHOVzZCHF8d+3Gi+oXQym
SY4xBhPH/uTnACLA3bPaLiLKmBvs3OC0Th9miZ928WrLXFD3ojAcCtHmjzxJq1xSIJg5kJ6QAx9Y
L9aLJ119TlDQO/zi+rrMZXm5ln2dPZGImdIsk/4Yv8xd9Ofd3ZtwP0+zSjgzdhOUQoOzvU22QXEt
BJU3J6DjKqzTR2m+Fv73bo290F68G9ljnyR+sj9l+Cqi7bmbbsAAwZQY0OKp504d+48QXqIJLhBU
mJfKdSU2STGgzzjIeyye2dlUb6ARkYAhSKngvLEZac2cmbIomNRIcryttkhZOmCeXrMEteblqbO/
QTem3IS/hvvszp5382mDtX/KS89bIs5zcGxbYGiFqDGeBtocip7c+2FkrZqJwI7dRCH0aQoIaDV5
BqQ2hJKBJIn5HybYqzNK1QRsGxt2dzh4M5mcppj0vn/cQ7M4TLIH0tE7mFq1SQt3gLllg8IvR+rE
W73RLCkB8C0dk0hI2uA9AbdDIc3KD9YtH/uUCJui6a7rwzJl1l9YIbg9lEcm7LDGYFk/2w5uVw+6
JLpLrC6SHZS2j1a/aBAZsU5fn0kVYQG1UXwkAEfBYkfegViLqvB7Qpsy1Wo8jnsqRmprYFgJ61FK
/4jm5uDLAhpDGyjYCBDFVozw9yMoaFI3KT0rJN0ufJ78OwLJKdPenwMPEmn+i74gXvVID9qxANV9
F2p4U/aDYrB2yRDCQU/8D6/bQNuZqD0AZWwYS0TDSSFrVwiVqaRXFRgG9VlxXG1gWdxQrthXwGyu
0pmLinsdX0WTAUiGlpMf/1Frx4SJ+4h6cA0XTqM/WxmLnFumoyxwhIccsZwKd9ciVwqHur5TgesA
juvyl5yM63S61ILDLlDxwUDZnvd2i89RRhTOzBuhFJX4e4qHL1ZFCgmidi886WFf5KG1Ci0UCfAD
bOjccya98IrH9VLgnJ702PgoW/bzCAXuQVN+toOVyA8Q6s9D0JdwdwTetvFLzrYDmM/IodYt4Zkq
GJHE/zdVkObofIRYN+3P3HO7h9mbKGsV4bWBvgdXVUuqE31rqtAs6VacPwawP+kF4pyJBrjbNlRl
j/LbQF04mOvq9emB9YBqAw35yTggEJv3tFv0Ff+ag6XT6YbHTAjzjmAaIoUXrCr8Vjg7ORx/gzSH
ibhpDaxM1ZxUioqj4oG1fh6aOgDv8la1w2tPX6UH3po96zxcTNRYmw8abgcVWhaGwEo5Tz45/gA+
sfFA+kAvpQkO9gLDELdaGWy0ARBHuvDhFX3paKcT5y/W0oBM6/1PlTf9Xg6Orp/klk42L4DmBz+W
XJhW3J343gblQvxInVnrgkKaIq1GpNX7ycQ889SxTnzYI9dyQvC7Kq+YUv9figXyrmGsWe4EyiYt
0KxEEwkJ0KkNg+tL6KFQsMtvk4R4EM7Luxeo6bEGecNXd0eedwZUAfpLU1Tln9CKUlOEyRcUgn4d
PPBQyfttI1niOrULG+g4fIbDZh5NvHe+faQvK3EJ+kI3Kv90DGEyH0/eEf4CeuMC7KcWgf8Loq34
nVmI1v+sV+OnU3RUvlIJnuE9nfC9QNsk8T983g/vxxm/Y8yayjPUeaOLrZqWwac3UxD/919n5VR7
HR//YsrpXPv7pdreXrkdBZNIlM2qydtIb3yGKl4Pj97fySQ+RSRQBUyh7sStCgCkM0leUel2ANZB
g8Tu6HWAyqYOQCmoQZB4CMriZMyLst6viliJNptJRBmT3D9uxO+dawkXUJC2hZxkqZsRelTzyMj/
xivOZuc3AFazPxTJg1Q4DYFnmxbM4jBJ/zUAG2Ya0NsT4YJT9NQ/jU55bxSx93u9cIm+43WE1eIY
MigejBIjCejnTjlyaXdZYXIzVkcBxfwRVQ5Ntbll9dGVBGgna0gEmProxh6tPWBNlTwqOcvzQQUP
SZ0tnPuHWFyKnxxaqxQfBNGn3ORYwt1WUEpK1robs4XI7E9XtKd28gteIvx58ZoayrOAOjgtLelU
xjOdrw6e7w3TL/C2bxWucInHxZbF71HCUfkNhn3pwXnz/3jaC+lYbJ0BqokJWZOrEgDvcFxSqI8w
BO2SFYlt8f2FiPNtAjUkxKzItw2jomm7LHhp00DNQfxI4//kBje0oV5wql87er+ZuDx5HRyuY2rN
rVjsk2lJBVCUEd9hWQYj9kffVh7an7TXnFyJAjkfOcjg02oz7q8/+cxrkCnK3HFNG5z20nfyUyOG
vh0yW2UCaE7uWA5xpw8btJMdrkIbw2nUVCC8WCL0hYXZsFOExXhtzA1sMkHDsoX7ce3zCRIL7O63
tAAzZzJAAlbPYQd+nj5F+xV14LYB20BZ0OvaulyIgeef0jFEN7VgRNRB2cNeL43TbJcMNMS4nIVM
+Ueryb+O8QMSKyRCFZLNUlXeZoN08MqUtvsHdH0TN3jlpRkJ3eEHWvhygn3F4l+ol8Ykz0zYtYsI
9K5JxhRHPWnZLt6qGQw/FG2OQ4ryjUm62KaIcKo1VVCgiKgreMQU1pElafwSxuidsFEv88W8n+65
7N/R3dJvj2EPTz6nOwbjVzjNnZrJl3lzXHlqrYvXe6b7s7zcabocoa3ET+AYcfs2OIel4/FuaJGl
LePrHMN/yk7p06LmGR+MURiVUSIfkIscNDLQSgmOQdgYDqQh/TerSsgaG48PxLgx3UvmqJCwv4Z9
LJggsnNtABbvU/VYcA0OTgN5tgGTsKlUHt85mKHGz8UMEyWkR8sZcizoa+49F1kMRne7YaDjA/hM
PeQFRhfc6glc87pD2j9gg7Lm60t0gOR0pl3sAqIfXIdxK0EXgJSF+xkIhH3Jc8DSGXlrFRYo0HRk
wcZTchZDdKxO+CeYls552Ghkg1L7SwXIzXQqlzcA68PYB/5+vEkkoYfyxetuwHEuC1ztpXq9XEPJ
Or1GK2VsPcnLnJcpS1D/yAabvtH533Zny6/65+bIF+h+Vn+zmU0OkIQ+emFCQEGOHBFd0V2D/KJh
ZuyBBVHi12S7WLnjU1dV2kdPQ5H2LZAuSV5/katxvpnzggzq8vOqzK/3kvYGtQszhbOZlwI4M/qO
p9RLsoi7Np9t1oUqtYcBfM2wCPf8Wf65IKrltMWMsB12rHzw52328wrUnxBPTfxsu+RaZQZAFiW3
Fx9Ry5zwridMqMpTDtEWs2sarErlj9RwZRr5efPL5KFPlVgjo+gRc2kBTWNIF8QZzVFYYSAXUIsp
li/Xj6eO/bSepPTab+QasYl+fhv8vKrdWGd5wd1YH/JeQUtDT8DLAJYCC1pEqzWlTa1eRkPqbawp
ujfD5cddTTGHGJ06VBXGNi5zsIzuzl59BBPZNPSHarg1gD+6QQMTUipqCx3aXoppjVkW7IBn4hAO
O83PuJwTtgl+V86kMhiR9Eug4kEjqHSS6aq7vzIjR+bqq6JK6urkc9Um3YkPv45Mj0MP8WUxZA2Y
brEYH0JJHLIF+oNu/eyP7/HLh30pdjnMzV6mBkvkEhrzFn1htCT4r7frQFDjhE2adxUKskjspLIV
q2L8B56I87qyCNu+H5foVkVzVVqg2bHwWuBnOxn5a0F7WLwo4Ei92jKVGXDhmkTnsD+XPDQq/XVw
Lbl652x+1ZKlOssZ3+Z3qi3UbdK8kUZpXFAROmYzbfESNZWso8m2UXdzz2jeOXAg1YtwupVFH2kd
6IW562IOfQW+zlW9a20Pw82O58HIOMI8SQ0T/xJBER/El/BOt1DFKooQYvu0c6Y+eb8yfGJlso7k
/cBksrU1Ny8VPL6z06ltJdZDR+L0Amh4JUW7d71auE8IcZc/qVm73K2wcD08DJjw+SvZcKIvSJuM
YIZkfAmgC0xzDkh8yCLWiB9tLlLAEAVvTxfdvQUVmRcjTnQYiNuyl5MOTwdXZLXW+FjzbY6Du12h
Sv2znZcvVdr5wcappitxZ9X7bDx7anFyn3DMoMce8Rq4Qp5gAH89ABPzgQBAvDJVEKVFrmKO/RQ/
wlw5+BfTMD2bvPBciywWcmgx4jtwEuSGf7JQh1CtJ+Lx1GZ+EUlLnxxH7ZTvfdmBC9Dar+mojr//
MceX4/sRQ5nWfn6Ptq2gb0Bq5QYfqqMcsDtrExLA2bs7IiCjlmzN6oTUEzF0Ncc76imWvjqH6RSg
NBnqMKSI042bHxbi53o+CWN4OqOVfWxxeaA44HBU8wHNNMBNwUqpZRjfReviB3FXd5dijUqb25mJ
nIA1YKN1e3WhqSrw4bx8CX1Fm6S25shDc66keyDyh6qZGnlSKtfZHkWvqzg2gvvULS503sLMEX7w
RtCrjVuv591PKvteTRjBCFwsJ4e59B2lIHW4QtJ1aUNpXkpyf20L93qbwktSVGz3RJ1YVeM1QNKM
tQ60H1rM6j9cdH6H0DZQ51GxlvAYXIxOFsiwLUfmUCSauYjjeKLTaeKifRvOZ2S50xY1F8vUx2h6
KOgo09UM1OFtV78EjijNjUYIdiQwQj0UxuUmCgmnCiSDBIyUkr9J7YmvHOISPZ0cubj0kcvs2HVl
f62fVob5rV1cHJuUwlV8XWfxyt8y1hYDdJ01xHmuOQT8E0HWL7GhEUN9dxwTRYjJIlTLTsRK4pqZ
80dY0abHAyTNawgVJzroJC802y2l4yf4YMZzvH4rBvwPHppBjEyuUTaL86UsdzRtiWTQOq5rTXzJ
VcptLDOvH5m9VbfR9fqaVrpJjxIft8hdaxaxVDCLExZvMqyG5DLwJkYpJhFlEFHN1RGxfcnE9iD4
CxoL+RbRmPy1uNbsztYuhk29a/lAclKlHDD3uYwTyHYh9F2xJIHkvcCryw23slz7NSx+Op5pTaZY
b/TgNhxkhQBGdd394EN2+u6/BWkmToe+gYwgox9Ox7Avb1K8ke/KlY695pH2TsF99P36DIWY0Fh9
Cmx+If4Myw39dhOv7eAnQb6wI5NfKktHekUpRjUeTyrFawZPvwgNwr0L22wIgoMWOfJOyR9D+kT1
6SX2aqLrXgxvuRQEUU5wmDyUb2afez+m4bUGlwfY6Gy2v+Z6bUt9jSj44PL3PQPN8qGGPuOLCHSF
WZ2HbG+QrlMCMcHQzUDS39OQ5d4bVtenbQJXrX6icAoiZPb+yH/bErLejxfB190lBfyYEkP22cWf
OQKzJie4hZ1BLbnT0MH2hNYerKYMT7dgXbL3FpAWArK26x63GQEvDzSdf2ATVowwNf2ZH8WUp+qd
5f38VKRFbcUCPkKYahfgfJtlwS4kxVuLEw9Ckrm1AfmOj8UKD2ZuJ4PQc82Hc+rGK1YL1KPLBzaN
fk0gz0d0V73daaKyJON2Ry3AbEnKwc82g1O7TCDvMuxxylxdQoYAsYqiW7limma8BraG6s3xL555
iWo/ehyyPvlyM/EBgKuMNtohp99YyM/3z7yvM4dyQdYMSZvJRDh8Pdh+VfJMGENqq//eSaALQj4y
H6Dx8jhfTwxBH1I3Wx41/Pmv0WEGHYf1oekH0TkJbXaPAkW9IOdF6aZcTGloVjOpWfOfp9dykTRg
wqynGGpUoaE+vYHNVIxYroA0+HqwOXpN9WJc76bVOOniUivxwHcJrdSwXZO51Ho2DPk6jiOXncuv
blhTvoYxLz1YVzeRluR5+TAkSVvVjyCBjJwgmfuvHLH58EXhgw0B/kwpCws5707ydW/4uA58oaM4
f5qZXVppjzVaLCUULA/HygDK+J+ezxNSYijPiKKuwwMAQzvc84+IDcVq96EbtwocaIWOlonwrXbu
f2lwPMOdG+f7WPz3oPXWpSSlcumETE/0Vz2qbPEmzmvcaJYEcov+l9xL10dr6Q9yQ7GhTfNchAUD
DEljRG/amUhTz4r8Yp1oOCYnHLIVtL5ep00x8/qHFL0UdaxpJdNUJ9yxVXbf3LSagnHPAwqqJKiz
cGJauMCX7O7Zm4vEi/5JYnSn62hbtDOPdD0R+j/rCnsxptWfsR29JvQvWTSao4+jQ8gy9U6MtVtu
sKOV6IXar07PO/V6QRfvmu81KEsOMW4f343qI9BhbaTwqZ9idPPXwgTS84e2L+J449iIEY+SBjUt
Ddw95SBZ/Oaq150dBXfqw4/JVN1GK9jBEDmZw6WYQ0mor0yuGalS9/JMpKLCNXp2hBfkKrwCXxam
mcpHRt16taFVLbbrHtF+H/NfrQN358S1rSv50UQ+ZR1Wr30U66ZmPrdS+8krq7qgn9/AxDTP/7ek
pxUt+e35LEriTbQnQ9VVP4cjE8husNWVbKCmdLUBimk+a+kCr3eol027+Btr678Xd8pruCjgUXIN
FgrNK7dDKNpVra3wkO2JH1uVWXG+EAPW8auTGQh1oEd/2N8J97xNMfD3yAgV/3CSWR0DFbHGtP+H
uIfNn3yCcITtxsvpWREXOHYLY7The3Kg4nd1G8wBKlmMkXe7tUM0cY2DPFI6b6/7Aazh4rNKiJX5
BE42EklwcC83ZJs1q2BbOeAigsgZtyBhtoVyTivIzQSCagXqU5MO7OLzVd1zzpOVCLFGQd9Gmcwr
QrLzVa+f5UMt/6ZBcoxgk1vuduHwpi8Imvto5FJvAYWZ4XVrbsuTb0JXW5LfG+l/rr171pGWV4IL
WPP8D0EOLmgtrOEFWHcO3MwcrdmLpW20CMhzJ+d+UyJR7mugXXK/ZNAFhrvwz+r/UFjZEFNIFZ2B
4RDhV4INBDgXT9OAVCN8ob0nh/5JCKp4eXgOgwtekTAoLOBMncpOe4fStw87o5Pr6qgWiNCJ2tMD
J0S3uCEAqjcgfEcK0QhiKs3NbGOdEkFvdV7q5wWOsDaCAQYzvguttm9+COFM5dTT9rMaBWwjJwCL
at23tNPV/HgstIg7djUmmUTLdIm0w256K0G5oPBWvMdt4Def0DUZZW4KbhTxpqt3M6dqMg5KQegZ
gWZKW8RomdD/RbXb6Qyc+ke6DgSjtD7Bx2MO6VI2CcYj5nQ1/5esUWZw1NViDvDtxPsPIvbDN6Uj
A2lrlMAv6KRDwiVKloojfD12+unhNowdMoWyn0NN7R2hV9CDxXeW9NDH6sJNY6s71FiwOLY7W69v
gEHxaSeCnvbOSV8U4/YnLw86C5ItqGoBvtCtxFX/k/4KCOAgAYwNcETGhaBAJ1PLKlLiDg+fUQrS
6A5YJIrvicmeQXqcY++/HWhTPx6mbAOgB9TdsW2D4wFvibr4Y5rrt3T4eckZrenkD2uBRuJx9Lwf
HBQwAP5jeQxjfBNPM0QMBNzPXqTX6rkIJoOM3OvYKWAPQAlAqJBm/oXL0hPRBuuRzT6TCi9Af2e6
NpWFR1fzDbozcm6fn4nBVNpc2Bqm42kpwSNENa4f3PrhEnU57Iq+NodghQZJu02lCCAoJNus26dN
UG+DLBcMroHHw57e2hNd4WjKlueELR6xGgCp/K2a3gd44FZv8ZrWB3VrXq2xu66d+4MN3gzbHfOW
RuDOTppbXH0d3+gmykkDu2HyQuBSDoUJEFwvvt0jzEqywqOXXEmc3bzinb7UBUh7l7LWcQUjZHgm
trXleDK7ZPE0CmwNh1CjlX3XW5tTPY62LcIeh7J3kBwrF/vBlCg+ILuvDb0aFb4y4Xc92G93AlvM
h0jpVpHtHqiDnlC5dbfWVsBNm4jpammgLIt94l43p/pE1e4+nmRc+LhdGd0XRM03oWkqmNtljuQ0
BX4HJgei2L6gJodGjZMgyVlZtX1TfQtKJYD1c6mzisXFpVP+tjVBIJ19iBrLMuCkkBs3Xfs1HN6c
4ccCf87umlH3wy7JnLZhgCVPWOxAHXXdo2ArVCflvZuUs+Ie5vJGHBaJgYyWmZpNdWz71EgXDss0
2+CaQbtiXyta1WOE+cLNXkfScB4/yExVOZCpjMRZ4L9A72TMjskhvryrVz8pNknzqvtAU7XmEymJ
gqNl+I6XGFe5OfsQk1si4+ZSCVkYNVodYP2iZZnMbeXeeAbdq7lOj+mBSLsElxOXf12irsTr2j20
NT9M5s5jtzdRTeFDMpakwVv3Fz+QN0LEe9tpuE2h8fXqCCVJcSSl1aFhJCUrftjcpWVePryyH5Hb
calFZkYcH4361RuMw9/2Dcl/oHWPsujooehdJNOdaU6CqkbSns+BElBEAZq7FaJh+ofs1xd4WPLZ
ZywhxH884GkucKRdVClKxECI3TC8kLIkAvYlw/UO6sB0ivMGJ0hCeq67NWOKihRc1TCYzH6co6A8
PfQh9wOFvummHvR13kfgmpaI0OPJQQta4amdu1JJrZjbbbQ03BzEL6Q9VIBeXRf7X6GyLXQF0IM7
FtITjf/yRGLedKA3DLrH78LEq5YRKWgFrgQkklf9PkGFYb4GEtX7HDPhEsEQjSMdAxtsIpuWGOeF
joPl7YIno78VKkvIXvw+oTgydtiuCMrcZRAwRtDDfU9ga6Z57AeYi6/CqTg/994nH3GnPZjUVJDr
yJlBHpEm8Vw78w4mQcAt42Zdtrfk6u0wf/gBOS0uybsmRQLiAWwIOSx1Zn1k1j7rc1ugJydwcNUV
NDJ53HjVyjkx26I49sAcivHcwNj+W8iy15jRgE0xnPXnCwzuBwndgwpDtF8atphPX2I4ZoM3pflm
O93nHdyHwJwm9WYVV6M7rPU04Xsoy9SaTNgLHFd+qRYkX/KVCM5QdfHeDb/k7kVJRQpg0gsurNxr
W+xSFtkIqI2GWsx3vdN9/3H9/IE/YVMJgFTVf/IHMGFv2PztPXMsuPhA1HNHn40gX+vEbC+QCfPA
GKPpuQLwiqMMsTV6QXLCPxb2UvdA8OHYfi+J25R7e+VraY8K9n0H2Hbqw1L3r0rfgp/RPGFAdFu2
HnF78NDs4XxgUVuT1K8ooTdTv2bBFRrw/xbi6rQK+70Qr+Xp/0J08JJE/VxRlgim36kQtMn4FhLh
ajQGKUJW1tsjnlNxCNeEITZBq/E2mfpZeb2tKy0HRusjoiBq+UkyLoB8R6S414WMZv1/wzCW22xV
51XR7TvChvIA+p/rgdYLbX+Zl6hEdbjuKCy34mPunzo/K7OVx9JYhG9NC51Se1NHMCNg9+M5ZkEO
UqpHhNzA/dmPrtnn8hzYbBTmuPEQv6rUv5rLTCHX5g5PFOawbZQBO4G6wm7j22zGICWolFFA/CHG
D8+gRMiZtwdKKlD250JW4a6mSiRpTFyijQCrZRLWiXHelRFp5UeLj2tB40EqDpj33KtB/hYAY3hE
6dLgJAQhxBA+x5Opz6hGeVbugJy2JOBxUPoXyQt/jDc1E0Yl7Vo2ycQF6klEF+jiKfh1QF84M5fb
7EqkkrwqLk+QjS5gf3MGJyrb4k3ZuygKsljjdIlOy9AQH1wdKBfql+xECCHOuocyUCaZfHNIzYw4
N2I+fXySAiTGCECivOC1Bq8+QGFdNJCrBDaCAlbDpvGgMeTlO4kUZrjwY9NmNp7AovhBgRaN3XIL
MaS6ig8YMd74ICJNyFJvYyeh9wxnBKcy5vO8AHeDvEnHXCzMX/rEsnHiFr/DVNGlXaNep3RvsLih
roRPHuOnVzuYFwnOeObQj5td+QMLX/8otbpc1qeb0cfqCDF3jh4uzVmAkRKj9zYA/xPOuB+zJUJu
n6/1+BtbzVU9vpklFiMQtpAqrMhbXBI+TrVmmEciUOv5qzGQnl+J5FIkyGfBehDT4Rg50BPNc7cw
CmEreSy5fJNceWjpa+rA+TgMB/DnQ1D+bZ93GPO0rnmM4ZiAjyMv6Dyy7uboRKyR+drhLetcOhLP
shVpFdzh6HfNKcwfAtFTPtpv7Saza0461lzM6V7DXOR9SC/wXjbjRDgEWWDo9g1Og2Uvhlm9eSgo
wSbVcvimg0wwG5jBT24C3odkhtlyvGZUHf7z8FHDVL4BbsEnSV5rUgV9os8ZZvRgc2OSqgdjxPKW
vg6SSOjucLvaEvig7szRZVLDiQo0ZEcYAmE2eJIt2+MF2Qd26xryhBLFYSzMMVRWWSD2THKZC4FA
p1ix5xYFzGQBeLS5s7QNf8iCEUFb5kMex2taNlEXaJ5uk4DEjV+pmWfnAHxI1UW+W1n43ysa+hG0
w77A548ha/9m9Un73Ukhmk75vVibkuCuMvX/llTCnkddaS7ei0h3j2Fqneu5b/lv8sCWyebzIQL0
emBkYksJsJshUkCr/UNv0ThNwmgNUIGG4PZjTjRFB2iTol0P/c+N1U0q2eO52q/yL0XSGnqSk1NX
w2Q28I6iXuUxnZjeJVXfJEeMWiZ+N1sfGyxO3lFcDT+Ha/9jcJvgXB7fcb4EAbU/kLvFioFIdnxe
e6AW5raxIshkDHqnoR2XshpGDQQlZzLGvBQEHnp9NDHBLKHod5gDsW9cPeNalmTfwSSXvytjz3MQ
+gJCT3gvzmMdKdr05BmcICfZL5NiaFhCgnSIFSwP7yOj//ehqBlH3+AkxP/MJVZWCmU8CpH5+yrc
mSyKuaBXSuFt4jZoYFjZCbgAmF84T2dtHVYI2KZsBtDMXCd0q45oVEqTNQDgkzdDCz+27XruOCHF
vktbC2FR7bh4R/Cryb/20WMTxBB6qKqpfdwnb8yqZYb/CJHmOTjC6Zm7HHw2WspxR6kQ7gusE4H9
E7oZcwQr/2QvUwjwY6dF+NjXIMHYsuwlBboB+9rETc71TlnvfjyvBooHyuSKnxdz2wuz/4FJ0Q0r
KpyABWxIY6yHact6Ven+V+9CgUUEzlNtT/gWPzVPgE0WdaSiu0NMcEG7C7MxATvUGEKOdvHkj8/9
O2Sxcj2sFnhR/RTOfKMFjeXmK6RfAbbWsN9lBCdhIQQIUKZ68RMV/mP2a71jp8JCmPe6+pXo0Vxj
mESNopA3fB5qjBt6IaSjf6mO03mD4p6LJJ8vZkEEo8k65mwsmJ8J1UHlH/68uUSfOp5kzyyWVuxJ
MEJfLcOe547GdQoBwtDFFo4zHs18apXwwrqvYiLTeKAtLhZQoSXYvVkOxNmo6se49WByzprdzliu
3r48IEN6kQJLgJ6QvhtAcpRF/23CR2um8HQcJhaAZ8+fR6CgkEliBInsc2kZho4Z9HpL+Em4hrLQ
gHV7989LsPiEQbRHXd0zJhKpOT2X0h6vVAe6W7HdMmC7tV6Xo3Fba8AgTDSQDeux6DNk7Vjjjx2h
OfwxNRm/00FOF+XeCx/pIzqEF40Y1BqrdWMffASAmtxdVRd5ocWoMGDDzKDp1K4IBGh+iv4+Z/w9
0Ni/Nfa75azBzLuPp+i7oW4VrEjWkomjmaFOfnL7V55f7bt9N7ZcFnomYaNxkPmA88szKVnxBSib
vlatscZdw6EzPqgvRrVqQDxq2FBfpDb7Sy3Csxy0aTUPVTnPanEEvBqsdYzPjMKBvZMYzEBmDl7B
HGgtrti/aDA6yGIln/sCL/58EvKhU2b3/7pdHQCiXiCX0tQb/FWQiLtQcFr/puFsWxnCbwulzsC3
3eDNYMMNggk5D7czeZqDABtJKMnoitTENlWsHGlyk+ZzuT8mPtjWOFK/1hNLewuVpzENQ5bBuDsk
DYlEKlHA7k70GgkqbztgZWxTzZMc9STBb4EdDkgEO0Zkh/ax3zIaOvtvtvy0SySOQyg0bUck8jI1
PxvQJvkhNJMb+UeSOqGCmwUjjRal6jiPFAlfHfx+NFiwdsmPfJokstWttR+zrPkNSQYafP4RgfrG
dDh7xpnt+YoIWS5fsLYJAOO6C9zAip5kJ55KK5rea6mMC3FNX59WBGrDreY6KfUHbCmERamVKzAL
j5sf+3WmX97koqCLaduAg/NDrpvbPqTWIzDQV2eX3z/YEZ1Ra1iNF538PBZtffyEyNkq3fYPqCjb
c7nlPiCWmV4+VPBSVmeZo9suJSPK9pRf6OMxNnOcN3jzd3TSIB/6C8EiENsmjXwn6kLDc+h8QI/b
GXS74CUMiyPUYPCzdmn2XuYhpHbcujT2ii63cnECgBI5ejYOjlqVqr7kAvStFmWaaoTvzOz6dhLV
def3gHtqGVMP2pbcBSRbtaXw7ss5LDPUlMg+QTQDUE14VSeMxyy3BuVvl6/bQVtRqxPlRZp7Hz/0
GsbR5bPJTxWBk61Wyyp490BAL3nzR+8QHkllTeM3Lu287SGVgT0x6F77mjhbEYP1qku2JYX9WXUL
4fYamAHnk41ErLswZw10rArxpStbxbuvlwYTXhcs8OxOGBFkvj0DUeEr9IYhXFnMXMzxpo8/hOCo
c+7Lrzonbm6AXCKKGvrS7iUIE1XAUshK0k7ztnXUUB6Logr6AdTXuTDHpscArn63KVKDk1eBhmnk
YhJYCJ0O6S+iRxGxpvUmn4EthKambhz9feRp/4UxM2q3gJkHXY3p9ttiAGGNCCKdJoHBreIkcbZl
5ZvOMlgVxQfK6k5s0e4vdK1OcfQtFqRwNOxBjpH/QI0M1FfzNtd/WMZtJxpS4pELYv+HVYqg5cW/
TnfwqEldNTYHERuMvRHNuY0hmgEawxMDyAMJLQQdVRK2RGOyqxRhJ+8PHaX0NQDJM8jHwNMWWov6
VmKHhFvJLdrG9w5Vqd+KWxKp64JE3uQ56/LaH6loxQn01M+p5wV8yMZmCJKs4pT+WDqcMu5h42KQ
VEgDvD25zKcT81uXh3yvSHNT1vL2nyBYZabZDWz2Ipo2Byh3L6MUXOE7Z7PgBMy+eZMnS8dQ1ugk
vlTHuNXt6UirrPH6C2viHN0obDgAnckbXoX7mFY+OSsQDw/d+5c8IErG4p5uLW89z1170MBEi20G
m/xqkC34VzEdk2T0ipEEqQrFOtcuMPT7+sqfEC5R1ouhp8a4LoGImx4wevFJMgDm48ppawGz0ujb
xzDHIN6KAMl+7kOFyFEUsfkxM7vvDnxsLWRzc4aT4vORbCrkCCEU2okcQjjbTXBUJTD4bAOvnMrm
KXuRayDW1ijUfVFEul/mm+TUk72fopLaaw7oeqPQODnu8GKUKC455HwDbiMnwS1b9F5jP/Pfu1K4
gNYq5/gmsdW9XiAXiQ4l8VAuBNIzYSkcyC+8DcZqmla1fWITEppjL79g8kJq4fFvrVjaOx1KS28+
Z1/gNUe3uhptdP5VnEeyLUjKLgKFXp3zjp17CrTkIRnYDC/P/TXC2h3Ql0A3o8iqDaVHgl1lhriB
bZ8W+k7gu8bG4Ssbsy1URgSGKhIYXFQZVYK4Zb4HSpvsjfgTfXJmxfX/F7chfDPYqKTJXQ+xq6zU
6UnFWSaeJr5Z73bKI8cvd8E7xLH8uBxcq3mlpRIXMeUw2aRSJ32a7tCuO2f4KskYtuLSnNreUNy/
KU5qkUYRP6TaV9A9bT5/eR1XjaZ3EVQKuz7c9a26kh88A+zKFPuaK8MAXSXiOAQlzGQQ+k3KDxrR
GVfVHiI//icDKnb53YGFHIdg89nukWtN/BhXVZ+THD2P+MCAjXxeD0nEIijXswUgtJ1QcmPISdDW
a2o7S1TdagyHd/FhAVNmsf6+yd7Crx/btorDfp70gcdsqY2vslzX5EtAC8PsVx4ERTWfl4QDdoXv
nsGBxNSusm5nG4u6yjzeoo04maofTwp5BLr4rYlx4XWb5hF3FjInkVB2Qvr5eHrQmpBKoa58ejjr
lqxiQalNuPLSbNv2fkJn6CDY/fMbHLIL/aPirePXmmDtdSfBsrqQ7wBtK0wtFeZWCCppmG61fac4
c0okc+LqdicVpFYRR25zjK8Ol2Y5oV0CnHWTGArVlPbEwcSK6tiiK04YXsXzLdxIuD/OSF5OtZKa
p3NSYz8FFcUVEQfg8Hy5tTN7L5Cgi+3dGRfZ5wM479rgoNh+N/hC53MWAgF2uWvGh5fhRyb9dkZb
1KLu0/a3wWp4ObsC6j7qIcDGeR1P6RjdeSQDMbDsqYWviXhOMKAndV1LPLrthZ23eJbuJyNx40hW
Ccc1eK3YkpF0ZvcUROA8jTtyXM3K4nYyKsHZIfsWlLapPL26D1vmtcnVal/UbcfRNWvBi/RAhsC0
70tKRwNH3+k2GbEhlf8R42/Z9oTQ4vef/UHuuKYELaXa7WbvkLSPHvXm3qk/p9Y/bGKwS/NR1Z0w
Zix0czrQXtgM3ykOmzCOkKKunpF1Q4do2pthbdsxB79UW9xpWuLUMyC67tNNtQCvdr5A4o2us8AN
y5TnlWXSqoLKwfCs1jGJThLXR+M9uTvvyBTFK2SksCCVJl3Q/f4DbCgDynr/rqT5FDiZEByJpEqR
bhHgyHYMbG9e3riGScmgy3OznG6o4fNOH+JB7zfTGJJlGVi8jVkHGgXtEX0+0r/LOKXdqn9ekSUl
cbWtGlX4JRKJrf2zqM8Fd0jRlcET2pyuoXSK20kKf1NFllFYzGgzF49VCJJ3FuT558x3jEDPJNqO
nuYWb+1QtqL1ql2b5lLgEBnadeAvDHPBv5nf8ZOuYhSjQ8odF+L+PWkgiD0rz0ilqsifwtUnLV7u
N4pd/0EorGi34Sql3hCEO6jghPXPwUefzC+eaTbf9hoIpXwVf9NDtlSwnHPs36H0isbVlhIl3Atl
lQUf6rF9p6yqsC2xlwCkvg9nhxkh/CrImDdjBgu8R62CfZqIpPUVdIMKtJ0TmQT5iK22NMRfzHzB
xkpNcXUUSdBDhz/dVlWb0PZ7fIY18VDtLcalDJEKthE/qoRCz2AirZOZ+jOFjkvsFf0gWTKw1RO9
byq8zDZx9+iUrHqxFwqYv06fRXJJoc8s/AfpcPNgsYj2GuKnbWvPB+d89t5w6wy0hGhm7SroTKr4
gODpXmPXUraiEuyRBPHgal2NtIiUg+UeFg8Xc/sKwPGU+D7/Li7w6Mg+pqvjySD1Bk9Obxsy0KHe
W7AXYzri5dPq3qMwevXI19HDgpx2BIa4ylD9qu3XF8MW99i3+oNZV+eDictLbSKWw1tmTIJNih9c
iIn+/m/8xNTNlc1mu9zw9JZ5mBhZ2iQZubiVtmLyQIElWPydqJe86va1RirlBIL7ul7d1uJR/Ev6
OO0uuD8ZJ1OWWV/Mmwnqp68BHLCUITbRp3nO+I1Kd6lk8sX/mSnNKOIDph+C6wTFjftf+KP7fJph
FLtHEVFozSHU0lp/HNBTIghQOysmQOd+5m2HgR5QCnetwjmxITJbGtW3kPYZ4TLdCHeamxd6sR/8
VpSBvEtQnhFEqUiY+jJpbhZ7JNq6vXb68Qg9351OCd2qwlH8T8pgAQwf7UdBN2ouNvVHR/wUEJGV
WF0QhznMJ9mCS+B+GJBI9zTLymrpQhdOj0xBsdRk6keml4gHUsNyEC9e4n1proXtraxewYiN+TWp
1tz0RLYiss8B6nSttMgjk2MfoLd1tIYcmab1qBdBXV1w2SYyxt4d15Z/+QyuC62KIxwUlMLC4J8t
T9TDQNFbRYjewYSUIV0YKQqgKVU9whNrQ9O5bgiuiVvu0+RfysPBdX5bvmV7QCUTcQdPZHBSvAxw
lLIoX15Htb10asUzZDe1Ifsn0kW//67g02n3r49vrx9rUUpsx9k1pGA6d3hrTs7wwo2IIF2+D8AX
2HaFPknjmceh2cEcnGWzXvuicGUudkAaz2nfbJnlMu3ioyMoxCTv+JaYFJUTa202umJEBBJIvFIV
hieMTe6rKiY3RTSu/FB0gl3fuJv4lfeK6vyxDcBj5DdO8mse0duDmBJEmRAWB9TsRnUrPttJBtIt
1+64q/OcoDIJUYSB2uk799Y45B6lH9/Vx5OliTbUfF/4u60OOOG3NWKJJZ5BMlZk29yEMU+x1z7Y
+2wsX3dG/rGMmSAQ0gX+x36bE4zxbZuUZAku+0BDM4nEGaMcTMrEIQK48HVGSmZO0uV7+qS6r8+9
Hg2Ht8vcdRPqX0IRGOkxX+ZtZqkgGK7M6mroQaLtLt7d+plB2vSUjRkBBHEM0PRIoNwbfUnUV1kE
4xS7pvFBpfgbGzEajZ7VC5NxCokPFa5HgKopTPx9QHa8/7LYVK1wfHR3zwmM1hZAY42Bhq33qWU+
92n91S2IMlvdWlIIOOmgjwoDeRukSNdlqVhMjB0JBhcLSuNS/KQ6nfes61u+WGTaKyLuopJZE6bh
FR6wH9Oydzs6LbN6G6Xx+G6/16PMBAkJ3aV8fhdGQXg38J//lHfBHXMF6u88rNjUKUoxQd5M9JWy
RzC4oJIMPZivzjhNGEgkbnKvEG92bQ3BazfJzIg4AigpC2k63K0fRPHcsUqJMK5vasy8BgBxc//t
/HJpnppsggtzjRddJ9KWsb2H/HFac6C9r7rskNDReA6WxkL4EMgP3zA5a/V4T17aexIamK8fhSU4
Hyvb8rWyUX//hLlvhh2CmVhp7l7ynyjvw2Dt3ydOyt6y79mqnRJO+Yx1xY4H5sQ1FhV8I0fhXVEU
LMxo3Sjcj6Eguq315fAtq+p2khmH2NVMT+rupN6Jr3fPy8n7pnxaqFVeuaSV3s7sIQa1SITjIyml
6mAZc7VGXi+PK7tyeiUB5Eo3HDFaFz/g+1jm5MHhyqTSnhEMKf7Xl8p8M7JMogHKW0lMCinTtGtw
INFrp+OYFL5ydNZo8q3DjoJvGFZIuoSNiXF5rFlhCKn6f3PfLbkwggZElQ2bKmo1/v0S0VjedTe/
R9y/UTogNfrxZMNUMLXCe6I5Dh4AG71m6h6YcuAMQehbf/E8rZOHwUo4P6w1G+0FsizB+8rQJiM3
YisyLcJ7+dlba2QUrE/boV5A7nSm8uPVfHzeT9tpp0hiEhABGgl0/6Yhc0fk8RpxmZ2se1zFUqZE
di7EFasLRLb1Ih0OuQevjgtXpWVL1jM6EYfmJ62tuOCioTJMj/fAU6fcxd5N//3q1Zthfhr1QarY
B+m+27F0ArNubfYj6+OoUtNUNr3wIxu/xY07siKModFSZhXshKH6fX2j00LJGf8MguRKeBPUvi3U
gZaOB2aBk/G2kMPNeCsaS7hdGdwGknpElJf9IKeZlsvZUHypUYt0zdnV552Jop0PqSf6dugNyejB
lJKaxcc5zBXE5Z8XZ4nt4RnIQ98UP/4VDcIlY8PFMO5DjYEEkEtEYChGqpeTKTQwRbZa39XCHo94
sEfBQapaPBjoL08pydIgB/BJ1BKq4ndHYNI8eRyr2Lw8CkOvf2HwGn8wQ/ixLIt8NxHRyyy/jq9L
tkn8yp3VupuOfn1+Wnbvn58RBtWzkMPB+jyBcfUB0IcY4KoxzW3oGBmjrrCy2nUtO2TOjuwAcq2H
cPUrYGNMcsf5T6PonRQ2KlidHwb8w64tK/e5TT7TaGUVcrvMoPZ/X3l4+qEHu4hD54p8a0IzQND4
pEA5i45k0TJshBityIKCN7+TTlGipAdORXnt5jxQcu6zcttNU6tHv1EQv26IFXLTq2c985eFPlW1
blbMRlD2KOLc//uybOIeI8PpVXNLLsFdk7vD6rSeNCKCLXYEjgniyP9+BquZXUBEfpJaBjUF9t7T
J515LeOPIR/c1kNMihkh2Sqc6I0PtDs9rI7Ln9jNQQL7ZS9O65y7Hm7rCOZXIkfge4hmn0z7n13W
1I/ktEQDXW9NhOT37RE3jpkS0J76VGjuBKW7qvhASy/oEZJpaP7af6VwEZ++1mzMjFYPWWQT/WaT
Qzt0TPLkMuZ9DopC4C3eOTrwl34lC44jCzF30AeEjDp2kIsppunY6Gt/Xa9H2hH2c8T0xRqzAoXz
FDkpGOGChcJYwoUQZJ1Ss9VY8v9H6vg1PVUQlPRUOAbshsNIJcWzLnXQWJVv82E4GgtXf/EIwdB1
hz7JAJAiK4ox//u2kYXrOYrIsf/F3orb1fw5S37OA2v00gvPExma1oa7JiyrWVQMivdqQg9dvmJH
C2tzmhjwYizVWy+lvrWj6laPH0S9ZJAtpzdwRM581fzSOV4jMGQhh6XgJm5kZDccSQ1pSb4FFAQb
dsUUR6tXmJuG5KRGPawljDTEVCEB4nR7CwzZ7qXhWP2puxOZRV6FRr6RhP1zckL4vJgFHqcpCQ2+
owAavFgoCbrvGrODDxYGaNb5F75saWJ5b2qKR1agA/uygcFZX3Yt+fh1tMNZ0GwJT+lNhe6UiZQJ
wG0K8JZeOyZiGzCbfs3G8lAGO/dzotGClYzMXlZTbzwUQluLz8km9JgU/u8esQVwFnKzxF3a61kT
ch3NoQ58Uqnne7zcW/2yntxox8AU3FJzu14rYBAdgScWeR+JDKVZX7Ejf9vKleciASIzv4aRRPKV
lghsYxgIBtBDDEkds9OmBPPkYtqY4BbLnrEwMgb3d5kHp0ytWKjTSCbDCSEcxj4k1kuoaw88aIdN
VCEoyN7Ou+hoAdChsr8CKWLqFX+GviIG8LgtSug2afTYtS6GP86732m1tX0t/YwmPC0SZqfTGckl
81XYbrhD5bM2Q42EKEO3BjL5saVH5yUwIzCUr04taUtAfOb1nRdZyQsr8wpGKlZbVBgfevlq7QKI
gvqlbeDva0wlelqL76aSldti6Qiam7wWFVbVGmYvGYVhqZijlGF17HOqFmiVGRKTAOBtez7aF0CG
ajf0kINY8pOKmC+aaE1pOJhSH86ltoQ8q4gz18rA2qg6LMC8anNDx/YiL3HA2R4VAH7lAjTUn0sZ
qHtNfvBNCRj0frHEimYuG1kX8jl6ZylrEjl3u5VxlfwB4RKMcpnVXslx1aRk/w0AiSRHUyS+iM9i
LvpoyzDJDwV3qnL0QlrlG01QagjWvSsu3bp0kvnbjFOUP/4UdH+PDiwVsNNmC79717DPCNXZM3xz
vInhPTphOAAJZ6VDuK9vfFp7vX5bpbyGW3uVu5Ax7vpXcfF879Q12soUuVTD/l5IhgfFOQTwGucD
YQ6zg1QQDXuD1mUHaMFoLcSsB+8xCu9Hrx1ewz1A0tJ+uUnIBCrjr9scG1Fw/p9G4VA9OJhDIxGz
PPYN0FqzwEvOimZb9UJaCHBJpLWj8zcbjtKyMr6VxQCw9puh3Oiz+JswJlVY89cmPG02135Y1UGj
8pN+k7fzhAR4fHx/W/ak3cGlGS0153zfTOfdwhFKDsNzYaP3REGtsLtpsfgEC2AtEmnP6ZabjYX1
xysZQ7+ivMzbHXK0JTyPqfNLokVj5MvgJj6fiOLPONQ02cbwXy6wdsWg59nMqeqejed+h4hCQPeM
xJkxcy93zdZSzfrvYh3Vz43oWVk89d9Vh9lU/HbgQVn14AdjYQri9Kn6HA32q40by1A7i+fyOYgv
1MOF2S08A4q8Vz+tNpifRscRYuO4lva483T7o8SMU81FJJYULmFoWEApSkzl5D1p0lhGuAt7kj+U
MwdH3nuTQdprUAOEaJT/cRAcGiugfynAGvL0nXZNtPCvJ8umKfMgli0vrhAtI5EZmRyoZHZ/BF81
OxT4GyAEFawekpDmvfRpJVUcEHaZtxKCBOVc5cMtDo7jUXwBnrMf7y2gybr4RR9tELyYJCFU8EvC
/y1OgAYeGoHtBa+7oS8YInEA+GPgAcN1wL7q9XfFDIZJ1YAzfEskfINVPh+Vj9HK0E4A4avOD5SQ
eM/y4F2rKap2LIESdw1jAKCX/Vseux+1cmbEBI+hIHYamahvFR4kbjqv2kqdTl8bYwMnqpua6fyd
5o26Afa7OzXE0hLzcZxofVqWThQ30wSaK5d8X2hgrX6bOGUOJjXBAh3nglkHdpow5HnLMcf/Z2Ll
PBN7dz/PY5rJxO0J0hElM5qZZG1jag342oqUMeWjxArv+RqYYD6Fmk/tmAW7mDIO6HpA8r4/a3df
ltNkYQ91Fv4s0pe/eZ/nfO22LyhK9r/YmvKps3KbMiMT08nPq00e+5FoGY23rIIUZ00LH5R4appZ
W/nTKEVKfcsIm1Tp+nTrTUxdCNhl2q1BK+4IgVmS89aamctXxtweRBE5Bg5o+IUovRSye1Le/Uy7
247thf9uxTkLHuCnNDlR6kmggz53zvoOCjRlHZWMSKfOjd2mXCPMF9CAiN9BBKyHugEBzmxY2zi2
PqXrp4p2yVcyIz52Rp8Fgax3Gaj1g/BFjOr92jhZQ9J5Cu1NdvRmVqSF95GrZ8vaOCCp3H4SSu6V
u0IlJSG3qknfUkevnIr32xBHG97LRGXnqSYb7qGG8s4NucBCUt2BOE+DJH24xcNUAIvc8uVooZI9
sRfY4DMB2/yem8uqrlTCUHRF1gbXJeTMb6qR/unJALlALfV8rQO9p8OmWPWBs+yIvb1k+J/9Ftrl
Sm3J7oyD/GHk5KFaTW/GVNADbP40XroJU9aiGj+KnL70taLOoU5gonyjmrEDv42t5XdpsSfEUyYa
x3TpHdpMCEfu3bs1UhT5QTOuuv0rcwe2APwZvYwbqKARJnHlJfKHO1djko49FbO0uzcA5M7FjO6b
DK+335Fe6yb5EbLmEEAgUp+nN6mSqaZOanWz/FHfhKb1XpdyuNIy68A7lAAoTkmAcnU+0STmF8Sn
BEC7wg4cHyEDqjA44AXC+GZaZXbAzR3kiyDce89lW/MUlgIernPVg1GBaIbyOrLCacFpmlKcXRXH
skd2LTu+bs/et1ougQtnkN0DDUWkygpm0qmyzHTLEkJ1dMw0zWJrCCNuNVAw93/Zra3M2t8g/8oz
BcsQ214L2/tIqlp6CcvMbzoBDEDB+VH//w5phPD+0rQVmPySAwb6lhuBZugSbTUd+4OgU6V/z7MH
MLRXyXEXRRJ22Lsv7aGOSL4HZr9LvppAvkBwFM8rwtbYSPIxVsed7PdhdTGBkOaUQ2pSL021ri4Y
DOzGwBnWb01NlVfotdtZ+Vo8qL7xjVSny9thV/QXX0kACMTaCwC3F/snkkwZM3xjWQAjpd9a+RTF
j87KiTn8Oos7/MFVxh8WOg959cVOfr9t0hf20MpBh0EzvxkUt+GuXu8z0Nz/c6fhlxsUX9IgTn4H
9YhIU5hwwXyBrQ/ofNwKTsfoyN/0XoCsIyhpNbMF4zQRuKc/RB9ntebwhoodUyxfAGeaJxlnt63v
PsIINz1eswj0MKrmpX7QuTz8nMguW0+g2Nd3GqhDM8vx/30VIVFrvRlplEk8tVs1TBIQBDOBJEUG
WabmP6lPSJD/amtuThoY4gJBNX9mPikoYVIlkphv517ayaQNo2U8Ck2FG2t/9BjhJPFXGt9vwTmW
CA1OuUS4WMp+IBZLdl2WBfby6kdIPT38cpiuklZ8ARkt6PMwKtFfPDfzJ9IJe37c/XixJFh4+08y
ILQbbatWN17aivo9O4R13x6WXGMNP9Rzq9Pm/30wUfAhu2oiHuCpI9fMKLdFijJqZoeBQE5ZeDHC
PNuDm9yemexYtlFz7+ZF8mPEmhOvZDr/5VIWJhMZ280mnVlX8c3agspdqWABVgHrsTAU85zgOL+T
oMHzvuDLkTIBrTgeY6B/WdxatYadZjflCoePrqmt7KQYu9KeBB74WNkkE6NHv5dtnJkaF+rr1q5+
jtxWW8lMZoBA2PN3XYM8XtDYDUWtog9xS5vKIqqlcQk8z5MtlhQbptsLZD3l/NvbKsNslObHJjz9
wzcvj0Qa2e3P8j27jAza5iffNU41xhNL0C7QWF7oUTDb5bsZ5XUzCvRfdB+7XW2QCpRhyxHSFGS2
VkKcs/LBYR1TnZIMEzIlVDpHlu3/fR5xhsUg2jlPO6FkJMSP2y+PpDYsfi7d+ALBN7IHKgHqB0s9
8SwKea6Q+w35IpoMryBzLuP1yaSp9yf632k+NDMG0UNkJmyGBm7R6n26Ebn+8oV3CtS/7LyTPoHA
2psHHYIfHgFZwDkLEjh7OXDuXc4EWjlkW7wsIXkXcCaZ5OCISWwrpg3+m5TFnvyMxXIMtmsFksTB
t/Vr+cuDT275XLWJgeuL8ib7owT4iDfNVbVVn8j3FWJsIjwDdkbMf1CPA9H7fslzIQ7tmsBB4w1C
/q2rsfhw21VGhxZOd4c9Z2Kc/GIJpOCJVK1WF5DmyGH0gAo+gKQvLeKB15/KyFYTwrRjMrVs3sic
UAvXCifLY8uZWRStQpYAGbc6ScZuIEiHX3HXQ+vWL/oSUHy1fpNDYw4ao/hcdaKL2SR9opj89IpO
AYDtIPxlrMPdcwPioXECSXaK51J8xVKhPy1cdAl0+tHRBs5BOYdRQpWQHV9R2R4A9VdWI/XVBlus
ijgSVIT+XlyuBiPynwQ1jw/eznaX5iRGgsahWfzdzk9lANmYlFOePs/pfXmJSrbXUedtnl2tKZA/
cIt9OhE1RgCcJA9ys6cMwrfqcxd7A2xTT4E9n9M2yg/bsF7pD5FzppLdJTJqzcQcm3z1YN7FMvxN
93Oh0cCFRtgHqOSx8vswG2wqVJhUVrzj8H32rIvrDMlv7PBn2b/eWaInDhfk3UsbBJ6X9oXKVjGj
tSaQPWxFeyceTvLQFJA/U9nXqdt/mXRviNohn+ZCtla/bhWAYRJyqUcTtv/jAWzI053Zvdc37+M+
4JoLg1VVBPL3UDAYVoh3Fdfy5fHcWSBYh55ZLRQW5NoRvs87Xptww8D21IjiSTS9ttasUOUt6n/U
cnVDWktbmv91R5j0zYy6Cp3X+erFwxd9jHC/+1LByN75psG1jY5uxewFgRzaa7MzT4kAxQjjmCCl
I0Wm/tQD2U5jZaFSs2SdVgNDvjyWGyvG5G5Lr1E343R78QDnseuXTidgQLx+bzWmqJuv7/Xyy1Jq
gi0SpLkRFH81XLS2ip74PIm8o+JbfwQUo3jRatvc5OwtY6wFMTqXDdYNhwLHmXUVyeAd3IZjh+hG
pkL1UEqvnikNW9CFmTVHO3iKk7GuHGRvY/hX57YwtT+kPO1L3Ad3KBpo1XIvjEB6B/sTMtn5rytT
oFtCnnkLaK3y1YCvRvkUnUP5Isw3dF8P24eu7vGORaTHGqPZohFoSvmhLZRqWr3ezZLUXEd/KbiW
akxHBO6dHEc9N6ISSc5ny80LnvQdPNAGs72Ls94jfa8INM3H86fd19o6jNS1wCDX2Uiju2zu7sZ5
++uasctplDDxS8X3Zy/RXUzaZ1NtLn/2yAG4yUHakIh2Lmqa2yp2Lg814TJVOHjUJ3dsqNCNWNmB
2b7kOAGJvy7e/EYq2dkY2ZGGGRa0ijYmVJVLsl+s1IWkbArj8c3qAj3hA3sdpGTFMTzFEXR7Toey
i0H1XDZ07yIiZCvVE+a/QNvrYR40KmiDGn1qWmFpFmlRLHgp+l7oPd98EIDY5ffBxroJ1in56+PA
egaHDGq/3mFsboJNWdwpOLQD0RFrqkiHw9lmx6KRvdHIbxzXB8b7azi62FJQ7YmsoK+tqj5746An
BR5rYZnNa+FDZ4dsNxXce5NU3wnzbIwGpU9SG7jyl7/d6lp0zO6MPKg4Zyu5BeWlSOLRFvaShP7n
Ow8PmLRtDY0vZE7kYHgkAZon/0v93hSJe0+1stuWYWfl572PbFIDHZ83Z+LQGMxdgeFBaSYFcaxt
By9ZW4JmFMlX547zS0uE5Cbkrnf0uc13lG4fOIuJt9GM6RDgkVrZrTf1TWR+fNqZT5OapoW0PyP0
b1mX3B8RBd6edW6kd/VJ1afGJUEShe1oD2ea0Ze4gGSBkr+vkNhhqtBUYGOgFCVK0V+f2sf/f8QM
qyXpRRfh6TacYmabNrHV8WMkvscFW5zW2zP0OrV7E92ZiE+cPUqlvK+spCEHqdkNvmYitkqZuwdh
jzkVhzqRdLBLB7JB8XRsgEZ6DLfctjAh5S8xr5sEKm7+fYCfPdZ8cP3AFM9/tjBjPsXdIEa29fZ7
A8K4S6e/IzlDIyMN2o87dsUWy3RlfX9bzeuM85CLMls/S9OlQmejg+ShYaEVAvI1sCcauY5+Pslz
7aO4E2oIPuYK1K+Qsd1s2HtT1LCuZsXQbB1RxB29Xeb4RFy/ukCFnBMdKWkffSqpsvoZ1E1XGglP
vq2OpjoX5M9mIozrpdmxHve1cn2w8LKexDeRxs7791ysaaBP1rccQBA2gz3ofQ4QtgqZc3mlfMsE
Heo5ITUvBIDT1De3vmtVWOsvXzZYRM+6dJ+CcLtjNKom2m1foaWkPf0uaP7l5Dci7dQczCelkMul
14TCfI3ZXfllQ2Y0jY2BjvU0J6IIaeee3PDM31nigN/ACC3oKYLuIZcJRO7xzi2BzA7o7DbLdKRz
m6Q+xwzJ5D9qEladjkH6TdVbslwEouMpcFZL4UAZoqvolzuOLT87SxZ6SJGC4nPxD+AC9P2YkNgU
uMOPmpnxYXupxTFZKSEZIx5Z0vIVG6bxN5u3Ao6+TmRBbkdP9i/aEZSmRQBLkFYZ0Uf7tzIFylR+
kj4Q1D7jX3ttB4r8Ur9xI46gFXAoqAbnWIePgh8ZZ1GAiCCvCELZUUDgPuFTr2JDceRPRYUuyQMz
Q0sbBvG/Cns8eXKOiPRms99v6TyTURugd3IGWF3OqpGhK3LkY/qZ0B3IJpAacL8WNgCvK48Hl3El
Mz6oN0Qtr6qZ6zFsgA8Puix6cjnToFCS1kUNZssL0v3tzsNGxJgbevi9JNaLcEqqZfkiHvOXaM+B
KBrFsrp1MbKpygwHuaUZjH/9e6CGISvKt0BQvWpoAYJgD88k4i5VPWXhX/s2xG1xJSzMAqMvtNx2
4aklVPTQnvR5wcXvbMO4YujkLCuZRoz+CD7QI9lVALBjNTzAHYPuzWkzm8vKDZSQ2LSwTblbToWz
+feYdfDNIRLcTk2HjPH46bn/jBPufkoI/VDHuBGvc92WwcRml+N57lSlhDjH+5vJRP5jiKxDhtaB
rZUvXD8K55wcTYYMrM6LJtYXw/g/q3a3HXdJg5wDGYUD4ovfZP05Yyz517qWpWAg8UYh5RBQvBaF
nLNUJs1PS/lc1Qbsse/fyvFb8DRz7vWtcuuBsyMSE7Pk4cg+JoJMbsiKyjYlrLiQrN8iE0+AM08J
6DyjrZHpjcPhAT2SAb1fsHolYX7A/wlaRooBauz1Ie4NKLPbjHy2Ck0LmUgdasNlkjgpPo6+oUkG
lRgEp/FI5xT0q1ppldFrNwFJJQGGUOuLeKTk8tHxZQz7FfM7l8Z7nimhve3h4jN9jeLRE7ftK1B9
zX+ZJamplzFhcBvRZWoapqeeXCmsd9Cs6Q/woCGBBDWzrz6I1uzUX2DnHlscoASiZQsT9UDf4XG7
XUmSCdyTuvh9zHhTbYiO9kZNPUiCHPm5UuJ/Z9nk+SRqhrAa+Kq0l7gVpu6v92UH8mdPy5CW63zH
3XhCGmrSVsK6+X4wD0jExi+uFB5Dp8CpDhRvqkC+TxFzGlBHN/KITyD0UkNNVPJlf36NLKlz78qI
A/AE84RWkuWNtwrptrV0bOuY6OakFVx7sRKTuQnpJm+eHES1P+mMLVe57j/7L+lFis/0hVeQVBBQ
keiuNdxeqJLBvoSGKPwxQt3lvSW/rGl0ClpVJNrKGtSr8+AirSTQQJnTbTwDiMRaq3+7W6k9uEa5
tm8duzt0wCxWJgqkbwYbEoBpow3XTjyWbtzM/E1LUUduyn0JNmyeYiLg0FWGT3uWEBA1hkHN8AAH
k9ePnYn6jo+H4pzFxIHna2g0gTzCrH+pirRmzJVEugk7H8bdzFdlynjBFJbfWl+42Q9dKbZjj7AF
xw2IDsc+lH1ntQvGsAGNqnwBaR5iyulaUPu3+7fexUEBz0YiqUFuOsdZZsj5IUKMKo+kr88RFYHU
fNfFpZggN0fFVLuwFAxsVcKJW6lCHJ5X+V4h2U07PSu5WqDvp5XBTEzXVIzBqL69efJ8MCjvw3bP
ZO3DyX8R7t6Xr7L20QPH56N3Ll2DvHSkYGQ5NcW/CkzTiL3CFDoyG0mhnU+OkONdTWcGNIeSPM3N
csRJcGDv6Wc0OM34c6Vlq4y3jxee0zOmDrQqfncrF/3RWuqtLqrfIgQqn4Dn/Lx42zKvB3704gbU
KGFbl/Uro5HPhp7QRI0OdYNSI5pP9OKowO65yGU/bjabzYg1yUEE7IIkticST1TpVXOYAseh1KE9
jIAyYLl3bNdC22sN1QvEeuuX0ldY7Vh2wpNnrDXC+kvJzrVKDQZVU9OXoogNoFrguxJX0+A/397D
No+ZmdboaoLOlOf70mhb1NsDQWeEi+Esyh2uZgY6rfQPqQXD7FJ8wKp/IZKNYWRFkjSQmkA1l33V
24rB2hfkFyJeLRsimjeN8hFIQXjytoBIi7BV42N5ht/8KJs0LrIjDOzXmQtBobQ8LiebqDOKqF3X
YoohzIvM8Kpq66dflCa8ra3nImSeZ1l/LH6ypBa71Wl9qmYVhhrM6bL8P3So66/UTZcjYet8GJia
VSUesiOHksuItiR60pcK5X6+YjfThPVTP/R5WE8RswY7AtOjKzrlC2FRoXCGxYizmod+apeThyXZ
Ojf96b/RxZt1cdf5kPa+pDQLmAW5xRMqq94zpemHd0uUOyLhFzJ0Al0XVP64R3pQrD9U5nL6avyb
C12Oc101KdzYX2snqmc1GTfrswm+OS785BGA6yMl8tAkSBONQkE8Cabgtk1Osv9M5cwaVtvMtQIT
QQ+H42TMlreN+a8h3YVCN6kJOQB0s5fCptkGqyuWjuJFaL0iwQ7Gw4gf4qXCAglK/kphEIGXGZUj
xbcQmhZMEBUvLDBuOo02N6w6Rm4Xkmjjh6735cIaiimAttugbsPNOoj8S8yEAGc0WIKr9amsvri2
r+h+r8wqMrNlcELi+B99rRAja9aR7Qbd/AFr4JYkLPjoCEXKjnl+YCheae9e3KJvlrdIXBOUlkt7
SL7F0M1pu0FutJiGk4rCrT7/+bWQXpHCM1DyiYCV4X30NzERUl0Vu6TO0YmvGiPqEiJGm/o6LSRq
CzzvK7ckM//f0jrrPdc7g8jNo6CGeyaPgb/SFJ77hVRyx6BBuFbIYsVqvrprvuawpYRhrKEw7zhM
lTFb6YuanXIdx6EqK7V1yJLcF0JM3HEHfuZ9URCS7PSO6bFko+O3Ds5AywMgMzzR1u4aHeybiKql
DD+iZzKh3c9AQL6StyeW6qxz4TulqisEeW+ghJQRThjl35oChXOS3ENL7h5V7QXQwQfY9QUeLp8E
KoOF7wsskw+sJsyv59cgSUTMd7SszofdduW1lQP+up4TIRwSW1LDkOLBXQsRjCxhZqMSv+dU3css
4nEh6y3XyjQolyafDpkfj1uXrHoEwPH1xTni/BXcFYqgneVRSR1/eNd4D1EprkVGhSHfzk4fiHVu
73sd2dr+9sFS2IAInSOn7SI91gfAV7J7YoGgbFI5a3AIPwKYMCnPe5FS8ua+Cm9Pcqxw8jfgWwIG
fKxF0Tg2IXxz/RURzY5PBEQoFmnJej35Ii59RiFTQazBOp0n8SWP3L1R8OUYiwd6ui6f18Fda/kM
k6kdKxnuGuZvVktnBfphDa03e5bxS1rIm9qVy8RvF+AyYGXnWhYTxTd6GwXV4ahKty4LV0hvumwK
vlyQv98wNHJjJMh42tKHEgC7CcjX173/LP+oPTKAcede/bzTMnwK0kL/KMUtDC7W/HU/aElAXVXh
5U6X+QRju6QqjGzQx2bfSwMonW6O2+AMSc0ngrBc+17R3c46SwxLFVzUHr5CixT16QKyvwRnPiYT
bQN3DH1wB837fImhDkpispvHZSBmGtnd8/oUjxy2hPxbOmz7ipsxgZzWjOeDCZ1nXEhnh6jiUjcn
HdUSdT+/vZstbgMzjYedgq4AA+8KoU+9su2BJDkNeEXPgay1lj8BIl5O0ewjpqyWTOpqe/yMWa2V
0z+m44kPZ4yxAn6zSYHYQVLwpOVA9ZJfb1nQY3hZr55Pha2vopZVJyHrI/BSh6f9PEJwhHa75Wq/
Y4TgmLfoSN3Fq1P7anc948h4ZdBQr1q9L2DiIT/GGB6C6QZY4rjkDtuJgak14EQdJSxXAG3nr4Pm
8APxLpzAwTT99Vv8CjBfvcrQheWvrViCH2b6KTeLaaCBj+ruhLpnUsDnoCge2cr+ssQMDO0JoMdX
5DPW1lUUGEuGX1hKuDcF67UByadTHtu7MEj/4oRwUAxWRZ1IVWH5J7yOJUdfSCxY4RNdagUAQYsB
9zdnKGmQg2aTtPuNZ1hqu2lVORKA9oKU9hNBzJUmljSGUJ9kYTM/AmVV7Jcvl7rJhOSmaP2kOtm3
wM35xtNFrwEqlFEQun0jckFbFTsryf1x1hqQXkUFyfjqFhmQ04pCDw9iFIBmjAQ+0ktCETq2FUVo
OswJfmCpr+0fWALB0K+GE/+i+wU5t3svxsiYZ394e7Zxy+aMfL+SXFA795FXCmAO4rf8A7ZdHodO
Le+WC7SXUx6U8VM+hCzRdn2eO63CvRZd/sNRecIlznMYVf9JjZWiIh3gPm58PbSRwuvsFoHwr3no
pqxrZa+RWW2BkMLgbtGupREk58YgPUiNSMZ/ZhWvpt7a69xMWm1Q9EC1x5y+jBjGXfdgzdeU5sdy
VeMQFhS8jGLIudp2GHQ/R/6Fjh+OZED4diOtW3aCU5V0BIHl7oPfSI3eMi0ZowZGNG3quY3kGu1a
hyPTQaY/h8ESl7nj6lfNrVOB2XgyDUl31Wy1B6jRhaAI5G6JAOfy36RYraJEMV+bwfn/iZLu7ES0
hCMB9hbksikqkJE6msrQuDZC95GfWNk02/TcW7Jvc/ZJh0CbVMjDbOm7d33f9PEj7899GdDCDc0A
u/mZE7VkU8eA/ntG30psI3PPnk0toCOZY85gEZVPbQQjCqQ4z9Malb9iWHVz7QtnuSoP/7ZPcrsH
4Xj7oNj3BsKtOFF9b3rIIaJPHDhwmZRE6E2thDfAHYYScepDOZSUjHkrn9DeGQQTGkqCDJMMfYIg
KpKNP0QZAuRi5P1U88nvy5YwuffTlBHTiVy896zLp/ydFfootUlHkFCGv+oP+pSaLrawCnN8Vv4C
lXW99bc9d9SwtEEyb9COeu26WMUVG9Itlplg0pNzhruJ2OwW0TZCfP7uhselh93kbGpxndUKInz6
qKhxL3Vc8+ombgBm/bRx/MYHsYB7Uy4Py52wmYzL4oVTBhVihV3z2E6x3EIDLtCCAa2PIK0XUfJ/
KKzWxjlKnZFwFZqDqCE1E8LKWDmvtmJ1xAgB0KnNQnzcexuLLZfgwuBwMS48py1QqxnEcwP+sU9u
d9J1KQX9WQQ1zsyRcK7L7Llmey44UdD7k66XVbcwWt8M+BbdK0IxObRiXOzUvkE0hEeb7VKfB/9q
i+8cWhbbyRuuNMS/MCPmKFiircE9iTO0VXKIyfiu/vSYotx/UYVMKNy1Oz9DibQxh2acHsByRvee
8H0RzVkbL9Y04bgY66Yp9nrsXKtz+MwNkeLdj8E+Hp5xkXGkyTo7JVvv50Sb6Z2Ucsu6idBIntZE
MnzQ4D3ugtkQLWYr/F1HXW/Ntl3Zen5uS4fS0xHEzr53/JtCZvTLYKYXMTB6sNSmzp+I965VMvWT
XIrRRBuaZh1OnDimcgrlK/NIoLTI2IPSOK3xeM25nEV/FDAtZZBY0CmNOGnpY9rpbC2jjeVzVYiv
wZ7l6G7mlbFz8n3UUkmDCMv6uB62ehf/7+v6b2PwUN82ueeg99tveVEwBlQWIkocpOBlSCvkMYfy
3eI+2nPbEIkx8v1A93nGfzokjecfwcLYzXzgWGl7m0SD1YAr6eAGVhi36P5CJSFhsfxwBcomcEPo
V+/Uks+s+QKFJsaf1ebZ4+/P25ExUFnwGWGzsMwWad7dEA/5HnbBfZ6Qa2VIA75JspyYJ4/QZM0x
+My7/NCIKlv0sWD2i5TcLphA0QFFjvkqVv7M+so66dFD/YuODBFHXzS+ohg2dydmU3eGfq5rQ77u
LoXYUKMP+DJ0YujAp5GJ/UF+x99VNBMzvsXi8lU0TGCrbyAFLHRBoS1LDZpsj/x7ehZvtcDy4rva
djIoiSsy7EBKMVxCbepxRyK/Y5PvjsEvcF3/TZjaT7iJZntY91Ib9UsWTouudiUlJ2WKAwRVsRAj
4uR2sYijr0ceqJX8VFYolHxrbr4qIbgZ83DBco2AdFu8MzV5ze+TIImhoXnDDYIrxvgHFZwLShYd
G/JEHF99RdHbuhGgMcLgkcBhQ58zAiXJkmwqcmkfRUp2uM3eYukHoqVasCSwh8iq10+HdD97xpo1
U3AwPKYd/sst/VKxZOyiOmtz/WKtKHMu7MWdpyYPutZCNzYUzcjqMhnbwn2lwEknU6TaQGcJYV31
xId8OD9Cr9xI451M74ULoGw7V+24QQk2jbh+fKDVInMyz320xIfCxf39AgRMdiBBRpcMxeNRv21X
1k477YDJBbFpYzzcE24MGfyJ9yZF2icGvsuMXA8isY6bTh4jAeWZT+o/B8Iie+K2e6yZ7SpTPvpH
vFTzwubwr47TZb2BC9ePOvNIyBx+gU8BW58B4HfLNWzq3cRRmTWbG2GIgpLkSUn9azusU01nX0Nl
tra1NNOUuv4xzyA558QecPIJErzKk4VUlLfW32HG4W2Pchjf5V43guGS74S7hXWOeak15A1o6sdP
TSsNDav7ZgbeSAOOQlYl6ol2rIjhhh0QzUF+wwfp1TMWV6IzPMOopeFJQbguhm9aS7II8brdeahZ
7yB529+ZWlpT5/ef7cRfO4eanWbtfEOkx4DSOijtiiZ2lHFYZDOI2IEHpXAYJV4G/Fh2jDoD/sQb
xjO1LFiu1wsexgnLau9xKYhEOpo2LW4g7i0ma13uYjsgjBOeCiZi7yZiH8oXclSEstwaLc00y5wR
S3TgmDy0Nq+A9YHa88h1iJC0BeDRXQ9/cD0PVIKvUEt6JdvZsAsaX4GC9Bm2uOTP55Rqf0wI4+Di
SrTR8eylluvJRCuzM0EsalBl4ZXfqyGE1vldctLeWSplefM1zhu3OPAgy6reOs3dtqiP27B3xy5E
fYX3wY8eG0cN6IZ2UM4mrYRjZsJUz9sZSTaeMzCTIAZmnC8IzzYtdKe2EXxtEftM2mRnBmcTiOfz
0+nhdzXdJpsCtkvgLxVG1TMYTFLB3H4kMg2QbaPKVUUh+hF+9gUT7uFT4uYbbFXL4aGvE6Vyvrs1
o/79bPs7PHf0NBuJWixJlOlzcpuk4+nJq0HARJfV7Fi4m3jUgSmw6Q7PRIeOccVzo8D7skuaeJw8
GyHrsQZJ53cTq9UHWvXQLADsSq+QK55p5M1o9/UHEVasPKxbRjc3FZSVKm3ljW4gXNXV07SMAgw2
hGWXv297+R3D+sUXI1I1n5YtSmPy/eBY10LgiIXtEaFF8b1PdL+Q1mgODfV1gGAww/pTappPvhD/
7wKKnsuc+9UqOWhJEbgBLVTf5YKSYPslj3x79Q0qP4Ej1DSfn1Cy0ZuAm2ga5hlgft75jw5US9Yo
6gMo5qOBwOLFhkmRiGaEdaC6DPjrbHip9bgXx+KsIJ7EEnOBcTMd+8IoBK/qq6h0Odlx28ToRB5m
duYp2fCHqmiyNvXq69hb1cdrCkHlkwWUXOiNlJuhFL9qtBXemu1Y0cCyGW3rZwTYjm/8nnr1mhdX
lmY0MGE8Ai6DK0QpEQBwCM1STovTKPmImVu0K13OG0bffNCTCBoWzUwyeH3B+6dnmzdTIJP5A6Cq
Z7KUef7kvxBTVQgX2UiUOhJLgSuTtGZ9+Z+pCtU9K8tKx+RZkcaCv0xkQTjseFt9mxi8FubBtGZY
VyyyML5sOyCQu0a+En5c9gjfPgNOqukWtfm1s3MCN1ioAbwkMMuq5xNch/R1SKmSVltlsuOf0zMg
ilOguHE6u5//UahIpCVxZWRaCQbxYNAYC2utUZvYCDjcNvOi3QwkXCyOZ4NfsMosfv4nn78tGHab
vf9hNy2Nuhph1Uus3/1aRj4EWMGKXoOkCa708ttG8PIVxlCFB4841FAdcV910zGNEaGmlzEvbcD9
sg2WoUzwT5+C36TQSPof4FJK6Yfc7kTszL9/cumswqeS2PN5kEwZ+RWcveFmCaug88KJ7putPpc4
NsQwpkPSXrQX1k332Bu3zgyy6HL1w3FYLKFjUwC2UC4N5hIf7hnWR5DF2RFHP+P7411kY7SLPVaZ
ht1b4EfqRGtAsxuppYYtdussCCiyqhMqCR7GF9Rv2hGq4wNQ5j3lT+NOLPqDCg4aPKHggkjK/Rg7
alN5HFEy/9O28nX3b33KRHrtWToSBGVlAlIglC6suTIIDDTH5PO4uTxRDWlIeMMiNBoP24udlUNS
1eT8EA9boYU2nFG6pNQfjX5CjrsBCAVX6/+oGDwdRUqV9nLmy4HwhgIueLreMI/KLtuia4PB6cNc
+NGs5puVqXZzkzCM8yWkA18rKq+66a70Hv5qeC1zGQYLhhajE2WAwhx627x3RebNgetw/n4d8kkh
ZeSEIch7YwpMLgCF7VZ/rlt1Kpnc1sP+pYRGYJ8ukZ5+MzhNFUSW21T+lhXq+zOGEnS1h6fkN+Xp
6uVCbj2R1ujzOVUKp32uPQNL8Mtq6n3B5h+hksiWJWfSh/zkQJn9MKaLveQl5DUOJhEI04SBd5mS
HtmQpjZRfvHdqdV97CBf4AEtABh6a6Bk6AsfevDjjTcn6uSh5s+WD9nXbeWz59YMfnnzOv2OP8oL
vWd44JLT+2P5z50J5T+LmXpYaC4+eHUnasBukqo2ICmkeNJFP4B0E3Xfj/Z0yu3rzw29PLvAxxcp
8tRq8FnRB7yE21wUh1g73YjQZl75BT1lMj3BZeOP5+B7CSM/Ckp/RI5HjoLGlLBpWi7epiB3vYLG
1cCBRkE1iSOkZklDPmm+63pN2SbgdEF2KVwxHz/fLR+JecAUoeCDWsHrsGwuG17ltJ8rDQNtupDj
I77elHaZXtzlrGkV8KSj5V/gqsgnppDl32EK/hD4slmLFg3D/95y6FpPmUNIYVm8SOvw9OguiVwA
FlbejXaAMm0f8u3GZtb/HJCN5cHsYwbiMr9/sE/rKm7W4fS5fPJoeTY+vNZbwMDFVbRvrabK0uXi
LFAOeii7LOAnZZfs9bFgLBh7G0v3lh8oDKcafydWL4aOluK5uTQ+qmT7MJv20NAv8iUVrOA83gvA
kw7JfIkTbHU6T2UtEG23RhYbcDRFTBE8r07L8G2FfEG0QYzHhQ2q30ey95nJ6hFNWS553vCvDQg9
WzyDqkJVWzkd1l+5bQD/xenfa9rjQoT3VZWE1eVSir+7iHne6KwfL+IBKn++XwNvjoXGrVyol+Lp
wCTLljtw5cwnv2DTDrTqBUQvvQcVPRzP202u5E4LmTZ8FDzld0fg1UyOZrc5pO5IWL9axkci+GZd
n+G9oRDrQtzn3mnV9E+k1WFCrsOulrFR1kZwYowtOf9xVYWMF/GT/imkuzdBxc+nXr/i93xnpl2s
2kEDhJSXdsBZYotjtMGNWPf+VHvE8xmuyl53t1l6qvTns+FIyqrt9nWMFiY5W6bSk110jY27xkW3
5+8DYPGNdE475WvVYEmKtqP1g/5Icm4P6tUPS9vbimsEfj5HaJUZBOdjy3GlQR2lPu66mZUYF1/W
tX7/IAbaXbSGKK9cds5dBkEF7Vs4suQ5U9VfG19bUqOIblw0UW3NquDMF+LL/XXT299xj5HVx2Hx
fzAH4NlNj0n289HH9fBLGveyTQ5hRTW1Ol4vciy8l3BIIyFkfsRf0q/gA+tIJKeGOSz4uPKQTuWX
Yd5beecKNfSiPF5JEv6DNwp8izfVLm0jhL0nwHH0VZyP3dLisMkF4YaOmyYMYLPCZhZNMrTUie9W
ObavjfGYVMcnijNijWlOrjjSzDFzWFFjsGMwwN5VOsQf/fvzKa3R2zH1JC1ZDW6PvWkna49DOds3
WsTTmwV5h+FbAOtoU7uUxEBeY3ZHYtzQU+z0NP1Egr1x+Vb2YTCxVyXpJ6AxV8ENjQEn899NjniR
Tg+ulXpZvXwjJTbo46c9/LZ7XhfGHAzujPCPUtvGxXu5svHEZTdNE2jq9yBmkiQvX7zQrrtSMyaK
mc9wkZSLIcNz9lvC074kuKD/ZtYtP4fZueXsn4aqRnYtwKfwiwJVE01q+Dj8V179SZ9JXWegnK3W
JiHr6gHFt4RWhkr2IUzDqX2gCS/EtY09lWySPEKOQu5yGFvd+B0iNMhb2l3RplAkJjdQa8w6Jhhz
6hFGqHlPCvAHD4A2R4jABLCHbB9Jp5X/LZiD3m8e7iBvzkAYniC26xye6zD12PHbGgQJqATy0+Ga
xwJbOdauUiL/De5SVJo/nhGRAyEvE/iv5ylnFYSWz/WhhvZeufdPdOQzAzDfWTUZ2A4yVT2aLOhS
Ze0RZM4CY0HljZrBMze2WnymKrf2TWTZYpQxQtJjgtlIJBOPt0nnaNvNvQyYRdjcMKDb4H4fuem1
+uNwNdKNX2coeA+UuHdNoCOVx5syWJWD62jJdAfP92l65Y2yzxDyMZLfvf7Qh9t5Kk73ld/XzBXt
HIO8JrbDJOHJQ4XaS2iSFwIowXupgvHVJPq19cESMXUYpo+bT67sk/Azau1mRck4S8pYLPLju4qs
qdG41NmcUu7/xzzzLFNXR12tQT/XrEnbM5+GuZuO8ZFigQtvFbPnyyVHy4Kd2AHty7POI//yhXcH
vharIRrsUoNfOjAJAod4hy3wUlR7Hw0up4ScCe3SM0vyVPlP1y635BF7ndfmGADrURQY6dFld17G
pTEMjsBa6/y356g2woxeDk23ZQrLGhg8yPcpuDNxT5qvWozywRXI7JqqkbNs9rz+xSytwdtxg9sR
gVDnuoJ8u4el8WkyVwK+zibdVdePX2HqXnzHvLq3ECQHHrlOFKhMvewRv0BmR4VYk8wnT4oqA8lM
J8fntQa1wBwzw5CnpV5hTlyJDbcIauAUObjkjsUhB5d9cDBHNiHPSqwNmJehrOYi3QT6h5ULuPHb
aGkMcTAxBPHDtZuBVeMeg4n/iFp2kDQ0naXeFJ5AHliedQF/9mX+2qM80HN0yOdKtkh18fFTnIAQ
pRA/1uoVbg6h/6L44+H7ChLa1switTh4DAjM1uzXDXTyPiynz5bXQh7IkoKbpragxi0gjx6lYgxU
2VSaqibrt+ij5Z2opXiCPq5XelmIcqyxRiO/vEWhgAvA6MMrYtYNMMfVFuKCtCZSBvNOVUeZ/JUy
tsqCiuHoS678mWxfsHy7RU9P/En5zZuPS+gLtm2/xKbVkMxW0OCYFeHr+IEmAqP3tbYWmM1J8MAb
FQhZ93tXOm8b17gjWU27uJP5+82NPphfA1T3QLaq/8E/pgap4bZlOXR2aIzpuoMA2ywHHA/kamUl
HVr+O0z6uBsx8ep9hG3bom8/hwzs5IpYZiyJRVdW5ug8dKp5oq+y2EN5PVzgLvxQ3cem5KbtjUQd
VtX1PQzdvOqAc3eE86jg+9DRFSZ4bF58fGq1G9eBwLLKenGc1bVnYuIbBkg6Lb90NGGIe1NpOErx
s1sF2FTip1uM0tRRtE5IXPfAjJT8H5SJFCxClbxlcts1eoPAfIz9Iboe+PvO8ug4gEW6m7BXKV7N
RTthwppdSXVNossddpKHy9zZ4hIyP4oDI1tTLUxe3UYHvEiD8biOopLK03neENp7BZSxztDJ/oV/
rF/RTwMs5jWDENVuKfcsi8tRLD2gTO6hZ1awEa3jiadX/kig27iiycSAVzIPLw1R8czJWwLeVnqI
+JjckIvBUh2ScA6KOK54W13XQ0lhs0Ru5igY2xp+uKJDymD6bNt40Yw0+9IBpTbkZ7R3PPPiAII5
hKWcONgR48cS6yeLEId6nb1a3+c4uqyEskKiKcuFXoPfgCYkSUKZjihBQvuSsFoCMMSPz6GENSrG
jYMbC7Yli7KYzIuXnn6M1S/A5sDVnSaV7EIJHoUc6zVAWj4vAxOCEKm78BmcTnuUXjlhX92zcfSd
kTjTT9y5OWm/MuOB7+yaAZQzV4QAoZS5bpHmwozBlnC8yo2lp6roxq4EpA2jXvBzxqUMBstzqGZm
PRFrDAD112vUUNoNm96Y4WUYFzXOLpc3OVJpcUJZ3+xM3i6xfsi+uZdkC+friZ2sUhGLLyFkcL2w
0mv4P4O1W9QxYfwoVj/yAaGfKJae+Fh6DP0gJw42QaJ9J5/D0EAnffrw6+Gpehb4EFnQtD+lz4Up
uVF2b12P78rOb6Vb58tpX9VY6vXWl+DHwwzfy3C8qSKsNqlQiEPqNt0Dmli32PS81eU6vFVPMIAD
AJ0XwNlkYNGAHNLrBzyte7kebEodsT/rji9pOovdwMrvMzaUFbzUyF+Nfr9MFgH/1Xi3KFpOcS82
QJKcj5py+nKY+RMUZ3kgTo5WVbJPu3/ylLSJ2UPMjJ7bCI9WhMmJmGgiFCjgHy5JEQ2PaqfBRdCA
97Cu31cLzjietVyKuxjGMtNnKOfaTIUi+IYJTFIX4DK/OLmu94hbbSFA9hX9Z8Ku+oGwglaD2Tej
Pb6B77jsOx0atGaQrCgAmr4yrFvoFWAtXmx/gMTztSThNPrSWwKnfWXzflCiwevsMcmtndm3kLJS
oc7MSpKa+td6o6SAONtDX+Dr81ISydi0RW6bmXQlNbPMfOGQIHU3rhR3PE5p76w6EfdfYmmiZwAo
A/QM+kX/AKotf1ahgLMneFK7Wc0tPa43Gy2oVo7a1r1Ej7Y5YHlfZDjRX1UDXOxXKXpTPvx3LNO3
DUTlYpcwxFRdZ5K5eR1NXvZg9P2iAVBR83UWnEHErxP91hORWbwNkYRRCRLTYJjcXCHjkTsDMNcj
G3O8nr6xkt8s4HG4VVouwGITk5iTldyMcXOS+jy9PwapV8R5NubfL653n0ZBC82WInTXFWfI37uD
QOGxfX1MLNjvQ2U6aNHXiOLJWk34O67KutxQF/6WrgMr0DJvhoKe8+BP9/AKA3E9Yf66gnnGVMHx
LKCNVMDm4F0tgW+QN2oAkRjsiGwnut0JOj2cEVcvjVSGrYJMlCjR7mmCys/3CpCZIENUOTTbJ7I0
qdDI5CmXYUbRCW8TkBrSIpull6avpDfPyglYmqNOkekfCeUtF6Qc8PSjT4Jl+vLp58ucWbOC4EFV
qZysDgBHsSAlz+IXGowgZ4nvgQYsspbRyN0kGFTv/IMGBrpARamhc5D3sNFDRVanI/BdIs6VDYHc
ZCDSAPSdTpZwmPTwGMnH6AIGD8KY8aapgShNGgSyvjZvvYHI5PVR7Urw4or8xWnqbiEuBT5ZbhfX
ZLEBUoqhX7TSizfH6o9zRrHWnr2l9vtoPr1RQKd9LJzczidUH1+kksnulWz/Wm57kK4A45hl+NLA
NDq+l7vESYSEvNAc8kfVEZZTD5RGchqVC0mi8n3namDZ6PNlZC+oz0iDzgjz8Eo9PZX2Uh019YJ8
jnInrNdi9hB3iZiyy3YNbopx2bPtVNWXj1EqAl5HuUTXrd6kucIVb9tGuHViA+deXz0HGos6qV7Y
8JBfEeNbNJ1tyxyMeEiefcmL9qEwm8Wlyd4UFgCEwSR/3tXQ1NM8PnCD4yKUutSqdznpvbqqxyVs
qUga9FYtzgn/NxZEs/kSH/Iz7JK1hrlMZgp0FD1MgAUtkCk/VEUSRaCvOAWU/kZRSt1QlX66W6rQ
K9fWSUwbSR1xSFIt+jwmW9YH5XGsOuMzhsTYWG8ipNSUJVksVpUbwEP1mPe1X9oFtabJ5a9GfUnR
61WaXJazw6HRS5fmcR+cpw3nPOjsDeqFfFgnFL4jMDDlWcdbmNEmFBjsBL6hZTYxURZrQj0wskS+
DbQERX6N3CQ6nU0CV1Xs1BXib/exxwSUCxfiTAkVaw4oKmtE/xs+5vrUDYLAGRMG821AaMaz83aP
TphSBBAxexsX5el3X6IiN6SexiLE2HLBmkS88s+kHJS6ZchLXZSTEKDhY54S4KXXrOF7mkXlTkMt
AdsGV/oKQjGOFVvo4yQlf24PJSOCfo9ZiDjppMswDQ4XEEg+YAUyLB0CyTwfLh17X6nV1sD6/cEK
zMWWVIQetkQKf3SkdJeicaJ9DlWnUTU8jBenmEJ6B6qUxiFi6cK9bShtfnmAeVAlG2lDNJfpzVsw
sp3zFmPkQfDw/JPJTyk3Fcl5ipveMZ6GDi/u3bVwgDmcAGDfck053EyGh5L5Squi1vFIwV/eNibi
2d4ns2nzwOe1Uhfwja0C0WhIoGBO2/PaXMgjLKIHGjGe3ZfVOB92y1wodtc/c4Mk2e41zJdIpYuN
e1LYTS+einHLeparfJeB65oPJ2spwIfcdagYoQCvZfpiuF/s2QqMGZCMIn235ZNxaCB4ryZ2jCXI
6y/Of+gGSKDIlvlD9vpzJZlhRqcynHZgc5M4zEKUrKk9WB2bZO4m4Dhj5r9bH09cPtQe868WPXSX
pk7piLk5x4Bz1ds6LzcejOg3KXGZiikIFWgHz1kb9ZnVVMRnbobPZ6ZZSzlyIN8bsuY8cesapgWJ
myzO7qJ5a0CE6FYqMyNMRat6xOR8J66C0UL20UM4HskRUtWwDQIM3P/iD7CJky8w8vsgXL1rJFV/
aqeDgqISVQL+3KY+0DTNUIQvwidSQKm6d1T/rsrIyC7BZHWhNxsGVMnzNl2nPnVPRcYrOU2S/JQ6
4/Fdp0n4m63bJJJWYXjpAhPiVYLa9krZPXva1PagbODSL0Ql4XixXiJPynw6/qtux6/uE4YTZKvw
0rm5dtXcRrSIQEFcaNG8kmTZf/O0THs1ljnx7qVaoG3DO/fip9aOZtOD5MTrferUZGOQOezeVBsy
1/u0OILLvFjDkW1w4jxuvSZ0pA7sBQn42uSgsMwlBqp6OyTZK73CU+yZSxJK29NgjEDH8ueJqFjP
KNAiiNHKC7V43mqOXuxFpfZI3GHXUECwqh9vOEv9wuQiuplMePeOmy2psG4bTewuHBUSNpo88b2j
N15+Fj+GNBfCi5GXqBgXwPDrXOSd5omb2IuD8+um+7CrFHrlyZS01dnaCdTVkjK3M3h1d5N2E5SO
0UcTWy7UiWDJhkfrQcs45jjXFcBAOFp63dKLszrLfsXI32Uj8eN7QX0n84758ai+ff54jwNAJja5
9BDRrwFVYJ5XF/2RsoH3tncKwLfKrRp9aoieuGgE3X9Q2LMI+SMO4yfwoSlmEusHTXXvktC1GllG
Ux0MkPanb3Si8hb/5VlAK5hS6I6yDUK5q0dizZH25yKSTfl5pFmKPeVsRdMRWThB+8mbihQ8Fo1W
kjRHfDmnQijebxdtezk7cFo00TzWuWZfjO+nsj8YJgWxL1N3H1me1bL3cFgB4PunwkJfrmBjZU7J
aN/v+cz2VMZiICxrR/GanLiHCpmd/awrS5lLumIoAR0yjzmWsWOXSFkcQ7DTFnRD4Zc+Q1Y1pUqR
uTLhkSwqyiTQh3U95zi99U7vWv9x0sbeSPG2Xu7ixJhDtdp36dEUVFr28C6ohTJxAhG+Q2iyzoAG
Bs83qdlvK6SraY+QRzO99O+dgsqRo1QkqDeXkKTupktESKUhPPl47iC3cfl4dMcs0Jv4NXPxCTTx
MI0oq5Z5VpjpInHQDMhj+JCqECyBPTGsTVru+Ry4Ytjn9Jo5nS8K+23weXYqUUnhJLt0WhmIfKNr
SxpwmFnJ3uuo7btoWIY3a/DD4X0wRmlzTvp8xpursz1pNUdoHIRoeoAtoso5ClbQJSPwq1x8QqnW
snIAbjBSsdo4SxW3vNKtNeRfef3kDjgCt04+VV0Avz8zjtdKNvD3Jarwy6JuO1wfB2rKh8Ut64re
lTigUaGsJa8F5ua5Akfv6SfatuT1YRF8hKzhhhQYKUO95bfOOXe9ihVu/LdR9PoGERDG4/klFhio
yUidyMYuxwb21g7572SXiCRufhIqTP8PHAa3hEVzc37q4XgaQ0QcTIdZTE+umxTw6yrAF7EY1jZq
c9aB/M/Py1ZNDrlUXiYg6U0uxxpyT4Uo58rFW7K0V0Y4PhjTtMRel0+LNVkkESmWD3/xreASFt5M
ZDM3HEOYywelpx2B/2qiuPKehd8vTDQTYT5JYajQWQPf2F6pTV8j5YV/fbgIOQK032aXIwMLx97L
IXiJMVYD2x0gpRMj+OCH+eUvbAjB+kx7vErvdsxx/IqnE712l2i4kJN0OYtydnrhUNiuKWqYykui
0P+yz2KT4UXUAqyI5Oy8BtRGyJenG57YeBiHQYdJ8H3gSTNPXwdEGSSRZuUEtgJYoaIb7glO0CIf
EbNKlkiE0okqajC2xKbPYOeDOKZ0UGYSqh8lpMofaaiHXrwY0LiIg3QkW1APQlfv/qJwd6eGJQ8L
XtIVP/UOOHY2N+dQB886L7LBXHwFpC2sdmSjYuWOWTwbnuQ+e8zM436tuLKvCbf8+B88zOS46QUv
OsgGmvzwzO3tYKV7q6QEVY21htZUZOFjwfQ98iBytx8QhVwisU97ZpDOQaXlx6w0bv1zMGMJfIHD
An3k3pEwwz3HNZkHvkSzQWgvRbRW0ESehZw9U0uf0iZ3HpXtWMvrZL7FCKq6c61aQiY1P13nKIhz
NyywJDncp/fSgdzpJIFwPjTP3MPtbAFg3EarN5OQpj7gNY36OD3jM9CqbD9rwa2Ddq0oqPwnJ5p1
kaxxDR6vIYC7ptV+BONfsDE6HlYNtcxNzROxFm6ubiBowQPPNOcwbIGqvAgTm3ny9OGtn8XHLH8r
0leL+VuUPtMP7OrRs1LNDLv0oIQM+s3Ufp7+1/QKglng1+TF1Xq/nOPkzXdM1vlUySApz4YLBR/A
7jXbktgSHXR7JHPWgYASiDyAhG60DFifr+o+UpSvwsVCqjSrRkXEHcdpxKvJwyZGiEfWE6EFo0lS
MvtkxhbJKbjwt0l0Noj9Gjbgi0y/CRGD1dZrFpzxXdwxvSXcyO1+1J3DmplEVtNM3d5Qbw+nPhOn
xFja/l7/AtGjfohAomcL/hdyKOY8CnygEQynM9FT08GKMhnFyt2Zq9tu1nhID1whxGGpzYynXkk2
LKGA2iVCdZdx3PohyFWa/O1my5dftM8UKZLXXo6OLaa9KKfVXP3k18IGb4TDfu/IG2lCC9ONR7Kx
TaReMJUvC81QnUzRg+h0MtdTbpaMXBP4al0LzL7C2yutn/CnfFKSV9G9KyK5OunQKL7OtDug9syz
EPQjs2NH0FcsmrRYKViM1hcJSi1/YhIwFLOej7t/yfHYgWdb1JGgedQUTjChSm6zDn2HJGqcy3Lg
pD5zOiBEYJjDUG5pLU99fbGxRbVX1y/NcjLtqvVF6aQrEbFVdFxRTXX1Mx3h+921S1AXvxwdtyj2
PFRCyS2viwtRyy0zoCMj/XBOUy4KR9tSjIcAwsPAPoTIFYYWXYCMyMEThiCxvwwLkcPv4kBeaSsi
RufCO/yrg5hvgER3KII8g7tQYs41lHjnMKmQ8daAgsSvyoEehrqzDnvD7/Joy8dh58Uq0dI8ocAm
Q7MccdgjQQeuBRBwbfU5X4fNpAi1hB7+AHlvWUF29tsM6O8JDisWHHB6oYwD3yGutU4kNtcGsL/W
Ezlz+wKUq2wy+irZ0toskj+PtQsN9HVTdLdMC2I3h1PfzutXuhHs+gI2zW2vjIkSxHD4pRMkvvWc
vAY5eROnqCzN+fmEjR0OYoXBfeRDUKizNjdhdiNNZp8xgXm6YabWuAenbu3PB/x23JngtKPYwRzn
rtgJhIZ7tN5mqUVI/8TPay6Gau2KAbCw78GMYG3qdtdid0l5h4l8sK8/GsM/e/KNokGTvGmCbAqn
6+e6my2zYv8cJPVr8YPAALhYqBvExn9ZmRpGIU5Lyye2Btp7sUNQAt17PHu8fS0Ebi1OJideTM8K
VLnfGpOf4fm8UyrCPjrisr9okFsCTnOIVtV2AQbKS6861U2+gEWnIH80itl69rWo6egGfKRF7sJI
laQXUB8mDvz2Nx6uafPOd/moNu5gue+3SdN4DNDzTqdLXcJY5hQqh5KT16wPYwk8/ocdn3m8RznU
JEGopQgnzhH+hjY4tOdNe2mNHUZIZEd63vWGNc+q5rJsmh8Jj1mxPx/XmYN3EWeMHowp3jV3Jwsi
dXwaur3RquqpqBdE80+QYnPtle328JWwYZfGz1GHf5rV+lTvoD7tJ8QDOn5+fVO8hd1ulVxzBgm6
GXmOrVM73bwSAs1mh34lGczVBXZ+GTuzjenXPkOxPvuHTfOvgG6TKdNMnq5lPF5kJVw+JSEEakId
BkXOCqTL/OONVOJ4PReuCDv+rHci1093aXHJbmi2kEJEmUx4Zvw5z3gE8Itk2oPgdAF/t3IH4W4K
4bDy7rdRLiuRdLdlB68r4gqCnmiP9d210yOdUbBQJ6FWyzLKYn9jHfFb61lq7QJZPoz3tFApbSoH
dYLQxZ+KAFV5SergqNyr1qq06FYkLoiyR9WhPcWABaNOaO5WQEguIM58hHQ8/IZb0WP8ZZ/zs+SH
5Zn3wuurLzRtacWzx9nVOmWQe71XbjyAfEbj0/1KIGjJ9WEVcE0Gk2a5vqtTPTNmbOIPNnsZ9ZKC
/kgyl3k7OWA1l5ke69X8k+PVK8UACy7VDgNJuzwsrPktpdNB3pVlBHx+uN/AnBX8bLTZAUvXRJx6
a/gPlW7apDLCh4NKqlT/Le/IuhRfkm6FDuMO6QEzZrDdJjaDCu408CbTFpqn//GuPBCW8eM1i1b+
s2htLs0RuccgJnitE9RxFhXPq5WzieoMI3XSDHwkPXabvWg55Fm/DjiBvdF5aPtM3JhiES8y1yU3
TwoUcQQgOW39L/gNzRWwnxKeX23rswjemZK6KwAgvBXoxnlZOVzM+Qcy1TH8YVapg4DVnFX04gHe
K3u2EGQgD4VR2Ck86+gNXgJPL687T2VmiJmypEATxAcqa/P8HJ/Z3+IyxN0wPuQKkTX6/tx1ZlyV
2JtKl7SawGan7jzLcpDaP7Rjs9lVjnBesduaOuVFcgAHIY16nVbWLVI/LiO8yPpmn6f/z77ZJQxG
ARhlSxLCsc9MvgkGCDuK9WG/dWl6gTWj0ZbKXjEajcYL8yxBvz3oizGskfEQs0LApeu3TfQILmjz
gCi8U7OUoYOhF85a4ZxmpSiMuiTfN2DdEpMrNX0EgeFFgiamnN9WdQ4oBvz2uP77LWU5QBtoeSgW
3c8k5arEo4FDcH8M4Qsl+xBdbY27SZ4V5NNKTra6KqF4+3PKSh8oil3NftEDkDSFcYrMf9S7AXnM
j52NANKK9r6CbcVnRVsygMuAdXnR8mhvTl7OAYGkT4jz87QqT7q2R7SHuKhFNReNvAn5Q7VennjG
/45QqYCy5khsKEsMTuZKzilcmomSRbxnfZi0eKqbnZPlnmBe/R1Bqsaor8nM1RtuPRvQ+BMDwxhp
4neG5a6+7MGfwbVrTFyhT3C5R0E7l4wo9TmXml/wVWROv2r0JAUzT4PTfRyNUBLBi6GToWrJba/f
dbo5QY2CDtq+zFItckMIDCQP1jKZvVZZf1xWDD769cxhO+lSUPj/41YBY+KSF8OmOnPFj0Y61kRP
jfHeeIJqKOkKcrLUpaa9CF6dcQaRya8225qY2s7IvEgP2W41ulwWVQbGHZOxtTS37l7uHVPQX4Fa
fAD7/vhgXFW8Op9OcecKdcsOiPsQzMMq8pohbY9X1AmtVBE6Uzs1xKKt5wrQYcDiGYuHrVV01fAJ
xx2ebxdS2iQlK0J9kpp9VmB3ly3JI627P04qosXu4pa6pvvr6yESu+w4Jp+7NorQoL1BTS92CcT3
LG7aTMkQQLlFJMsKu/KQmk3EnYSELRzeNeyuyXAVYa94Slxrl5zqdGXQ5n0uD5JidZr8DayIwWuI
0nHKggGRuQkbVPlEr948LwzT51BdZ5IDXQgzHuzMqWT3+XpiOTchmnsCAsjyGo7m1gy2Gf7sR3VY
wJjIU/iRwgGZ7PHeDRxUttCyCjkHshw/4qfBVRZFXFOb1lYe3hdDlI6FCt2vFmeegBk5N7BNg3bQ
DE5TFGQz2z1LQC3Sfx48Fr9buShNhrHgIEmtorOH4AcL/DJR3HWxeuTn1Khv4Oog8DBfDxoxkzsi
318NN0iWIFC4Ta6maubHwuLcBVnWsZ/X5LMAdDJyR2VvZVKJUv/Hl3IapZZcVX3lYqx2A4XKIfAJ
SQVMUVkm3W1SRcEkO1W0mUrl+9SUAwPwROw4Ve/SQCE/EPUBKBFhxI0qO8TIH6sXRUzQ+NVdIBz9
av6ogXAqDTZSeCNpPgBzfN42d3AQEacC5UrZgwrQ7aCc0pqDGa2GTQ6ojFzx3YOanjangIZzNHD6
bq5iQ5JRhI3a1wzj+7BRU0ntwa0NM+418hVZUoXChhX+JFfOww0CKdMkBe6BVd6CsP6MnpHI3SOr
8PBSrTDOEggbeyy4d36640VDp/NBnZpzP7jFwJp2EQUFmH76VeaHuWfAT+tq5+mLd5n6HQSomKxL
2IoFclz0403RMUnGXWG5v/x9+Nxujurr5/s4zRuYvv/X/zA8o/c6YnQNA65sTiFeRWYUjeoWYAyP
WCXh6DBPfM4NJV3Tvhq1h4c+Q9Mqaj5bkbTGuQaeF2MQyLgxxEf+ilYEZLHS8013o8pX31kp8gYY
C+Xm9pwoqKDZ0xGPEV3QDZWkXoBBKJTdPMG6jnMVegZZDg1WiOC8LYvcJfHkwaC1Sa95GGVqBY1+
iTYvCW3gcf6NPCPCDAEzQTciFe10Zn2ckNuW3BbpG+n5YE9r5oli0xHlVD65ylJBtgLiwRx/mD49
uRCQJekHssmNsbL4XfWL8EPMh6q0/kphUCNjn1EtEbNsOvqBJkFXenG+mRXbUArQuC9ap6IoQZ7c
mS6kjXBLtq0V6Wt0BTfGB7+8XE5lprZAHvM8BYCIK2g7JDp7iSJocwxVkeWq2LNWBWra2p++j5KV
tmEN8vwenes2lmjiZUUJs7BMetRk+hwnuvThX6M/c3r1tc6RM1+4hDd+Zaj3WIkh4WkhJGE4buUO
NFhYdI6OWklE2eVM8LUaLtztnRwf9jzXaPY2q6saGgtseFCQeIvoJr/67wtl+N7H9/guRll6P8sD
HIUa8YJpIvqntPJZUNNMPvcMWueZOHCsXuOuysef6hCcYpmA4R4FXJz1wKvV/lwfNl+SSUEHiIPe
Bid6E7qimgKd2GDi9S/vwVyOU2XPhtL8NkXfbfUnKgfBQ4mh/5hXtuqpEdtXcfjo5/dzQ3tjJZHa
Q6aM9bWRENlYH4inn62wrztrFLdgJr/cEZsXiCSdUajUHKktSmFs36udWnbo9YIeQ7XNvxK5cmpL
UntScEH8gvv07U6RMXT3rqx/ojdhh6iJXhWjFBCnexOW8WIB/7iMN9k8E8qQ07MBNMpMdTeog9DK
e1CY6YD1Lv07D+fITNqSK34Qen6A3asxvl/wGBJnMYCbcS+/tbzaAsu06ILrTwhBxXbq8ZdQ7kYg
iZ82aJaOC00tYqwNmwBa3Wq/cJID26u1puEvBct8lPsVgsVTAJzuFnU3tNWxihaHWNkRJBdn2Ku7
tCl+zKrZHqpsbTYyyYiwVfdnKwYbJlegG68uYS8b9fQg1anCjB2Rw9qoLRxj7aAOSHNXfZCQn1kS
PAWw07y0vfZKGWRoZ80BHutw1tzrjdKPhU4cqcjJ7DmMqzLFqT5ijV1uZdeERvytu5kObAIbcil9
cDgep1JBzIRbCi3vrB7h/01kjlFfr8FWEdrUY3nN6AK2+aFGItqLGMZRlQH41PqWMq+QPGhuIimL
zxasH5fqW3bWW9jhtSzKnU4gPM+l9xsKRV9bpwP5+5MBPvNNfgcsk41rngrEvR4K3coTqkBIBz/b
PZITz4f4fuce9Cuz8d8/zZw5Gk1JtMQr8iLc3SRPGklLwJc/QIipKuQZV0izgsO/8k4mFYqX9Hs4
DdfC0qER9FQ+I7D64ItjUQc4NLJT3fmp6suWNhEG3xsZoV2RhmNJHdZj4uFTFxjioFdm9nffgfZ4
QVksa0pOgpIkh6iBBQbYVpzGAmlFQqs7qEgnIxb7dWkQqZp3nnptiEeYGgYvJ0dXxNHk7Q3cT4GI
duq0hAyMXFsv/5Xrxa9+LxBfMRGb6W079w9mERKBmerf71QwGy3cgb/rxPHj4YNDy0s8xp90FePY
J6inMPN5Wb9ZYnoM9/opIK870DnuKI2kdTuU/Xxl3dLP/UdFyRSuQhlruZ6Uq7Z45Cflzx7YfxyX
6+Ek5rwey4eCT38BM5vlMr1Zbz6NYSSLopca+ikJrbc6dfX/vLmrDrYgHOBHHf4Ih9xAjAffW8wx
ANVw80h95kueshCfVkEH6pC0tLM9orZ6/XjRkKQglAn3/8bxnP+vSwZCYHWJB8W2l8r5rNV2wjYK
+PQr0EttjOHYHd1D+M5/Kq+7vSmUj3jBE7ADrTBoJ9CzDshUwJwzfIiEcdX6DTdRy11H4txiIloQ
eim6y+z+UhX8Z6m7LjyTeqqk0tsQDlNQrr+rRUI7Q8TFNYB7g2EPgY3P81zy3Xv9QmH+ZHGItXaO
NhJt6xx78Q3UsT7Dq43STfalGaykl9RT98SVj8norBw52zSDPh076SDHyCuiVW83ybIR0w8TjdJs
NgtmS30Drwf4dmjRI9BiB3MhbohreoWgZz38a9uHoEf0imcftJ6uG8AhfgLu6c0TIeTrslgYJuQ1
LQ8PmS4B+sLdifj/oRMHribDIWTbhIQuLpp1pv4xCyxgQ0VFfHyZbf5AiQyDNWM836XgktTxZQzE
8CBlH+bmG3hVZ9XD1Y18p5Q8VmKCL1FP5NK+ozBwMFoBkBD1/RMOgtI9TTir8xcFwGnOtmNgj2wy
7sni7xrERjLGl51A4xpgVRwKDiZ5jPUGMwwBkJcBY9HPzIrmZPP7p43ArgDWK2eOuJfACUHyS6XK
I+xbOns5+sdFluPJTa/No6zjhALngUR6n0CBpLspgCyHS7MdgsWcNpVXmngooWoXSr+acisFWVhq
PlXRx6M+ExQJTk9tgp3ELEAsl8EdVF7+3pckVX8kZD0YXt1X9c7r06CdIsXTKQSF6DJjBPI7a4AV
DRK+ubVLKUqQfCXg2yBYQ5U5a2/gH+geeLlU2ljbHgWiNGvImaGLCletzPXAzvPdjalR/0UDkVTx
Q+ILSCqRi2OaK97mJASa0S6mY4b8IWc1lp3RltLmWmPuvp7xgDZ967wpUMfLAnbHq+H4TlA7HTpL
9laCqkKU25qoF1fpmqzQ9hCFr4u76SATCTICKbQ74skOI0SZwBanrQyi57OJ41zX4yETpZq96rLA
8w/GLJHZAM//5b1N8DbOWNXWjum74lV95wp6oRtOpNh4xavIsTrXk3L57FC8Mx2sauYe5JhgN2oT
abTU0UwmsdKCsCrx371JAeOxxG0vQR5NLltYdR6pI+Z5XpcPPNmfxJZwBMzAV24oxPosnl+t6q+D
Tuyn+cqN9pbYVvbFoOUnT4hsT2/s849hxKvJ14m9J3YUWewDdg/i0vjDdXBBBpnMbWEJiI/SJUDb
ZaBmTGx9wftTHhJa5P4gLTuU11o5X95kc3n5nFpHrRd2wJc2LWAZ/Lwho1UpqlVMC5QoCGL+L6u8
QTmKW1LUqR1AVxyYkmjKclw3+uBiVxwuaTNHlwkMkSB9n1inncTvF9wo7YWNikk2PFhhRJ7bRfkY
sb0KsQB5Dc0IAASNxxTpO0sSD16Dd8bfEkfgGb5vKY1Q56k6O/ibPvtQpWGoxzhOT1lkJcZVfPzW
eSVEgNrDXdUaM6kNC4xn+Nz6eLfMHq1LtrT/yK0RAGPrfUP8dDAoB5fFsYjMbOgGm6+neMafF6Fi
qicgO6bHphkybk+CZ7ZlU6aT2z19Cart0ISD4F01KblWZQSOKcOxA3N11+aub19pew6fHrDGI/RC
JbQzzTpuY4LnLkT9bFCibwuYIiYlo7WIl3RA7DyH3rl3yYZO2yi+ahG7iLPJp2qlA1SC4FIyV6UT
XsGVWe+qB8Uk9NgKS8H6FxvscqzFE6Ia++dF6Zrhd04rzyjP7VM6GvKIJ9HHplh5w5Khw81NPdDE
SEPmNi0sCe6SwROZb+AvYp8jiZfpyAnxe0dCL4G2zvKkxI4xdDXKFpUzJMaFvYTNiBd0YDNIPvp8
0wpZK4u0gHpaVhw+3Xxp3vbttWFQF2Q0ZgAs3jqhA2KWsys9P2l2CPtnR25BykJvZa5pB9rYGJuv
tEhzlHcVvXOFNsYE5y/QnT5nESrdLoRd7wk92fZLMmxHw9qf/h1VmnP5FIMRDvaKchNu8auTYQQU
3/cjbFF1QKLnGAN9V2jq4tCIopXPyq6wjm2kN8XVCLvFGk0sMcz+hqGwm/6f75F3Sc0/QW8AuHYW
jU4V+SnYix3wF2kBCVIvX9BYHJlz5z/BRobSFsJ10+W/z6J84CDs2P8gUGKBFOkocZuYhMuAUgql
LYoPaLQS3xacijKn/DjExUUgr2v53l2elvjr2GxHGRxAZINH+iExD6mW7FuqY8BMHqvsMLqJES+V
fgK0WeiooC9orvVMBdt/HGBDtAqarwXZ3PkpleBZfNa9Jj2sgaNo8YvN/Me88vRlZkey3O3I4b3Z
7z5VkpADMRQaUoxZHmsHRgrBpPcq2KdSe2TnYARy02YX4+j+CZXiXM8GZqU5VHVhttHBU1pAKrht
2ijCc5ADq1HQif4wFJTmfy6lnkVzvMCEgsv5kVd5u9brWk+cevEEIZYcgFsUAEwW1lDV1mLJp4ID
NpAP6BMbID1tNPw+JeHswMT7ZJypAN71vM8eip/BCemp03hWMMdEwWC24ERGjI0S9Phnm9zqbQ4F
LEXKDLwnnDWHdgIKmy28xaiXpDW1iG+b92nh9Lw0g2QtuNyAENE7darf6OMnyq5EzBa32vs7h88r
wHKJQqNjwdGp+Xn1g424Jk80DknXG6gAXaQh+PGhei0a7+nqteKGohiEV8At/Op1uJrgCoMZEvZ2
evjMVIM7YkL2Sa1DEBKg+r6lcQP5YR6x5fPoN1rdI/6FBQF30h3zQzfqD27fLLNYllLnC3YEKPMZ
n7yVBPC0exw+rOW3BJhusjaKSj/Vkrn3s6/40lky5Egpm8k2628vvQaMkmvjqujZMfcmNiUuljUa
pB4g82joWDQ+3podh8JMC+3ss7dRUu5H8MJooLo1QInRjlraHqwZ04vUB9yJTkRDbUCeIxvsK3dy
F/9mtjaqWApPmGRlndzkJfEwKob2pHUT+P5rljvaV5axbY3Vut0gnzhr58vpwhVTjRRk2WJSTf2J
zRsLeDZejF2LBf0eRGNKof9puJjt5BrJ6GLoghqC5w5ENDkFN7AhEsBq0bfdWYjtKs3r6Guqktve
Y8g6fTlUPIbhJ5nyFE6HKYmJimK8j0qqLU0SnXEqW4hjGxr1rIg1XejBMa3u84eK0Aw4aAwd3WuM
o8PVHA0UNXcKNfAXczTwIh5PpQAThQ1MiuutIx4/MgvtE7NDekLs2W4YWxdpk0Ld50nILwYV4TY2
fqQVg3nyvuHoPxeyZ86hYFbom44XIKm8um9WtM5tYYywyJklFxwy/hUy7stmBhHBiURVPYRZXz8p
5nqz26mapZoIcEhcT3XEtlCG5OkoOh+0tExDdlg3sf8/wfKAVhnvCvxf/QjmYeSFovAUs0lliPbV
9cTnNXbh2l3LVEFZNrWXOtotU2EZRSQHeP2eSo74PSd5DZkws+Og47qsvIw5JHOIHOxDFKv3cO2D
x3tVeNy+98ssppls2C5nMildeTEbhtf2dPYE4cNqhl+8YLL2xufu68DNnXaLaLBkkhTvtpYcXACZ
0u/I8zTf3yEB/l5mdVZQWknsG08/ZRYcJOopZdnUjqmV4ltGbRinM5VqFGIyGYg6KJ9HNMEG47kk
EdP5f+/ALiT7IkcI6RXnWGq75gaD/qH/vKVnlMSkcZzNeDVlCI74It5mzi+6Ur16RKLiZGN4Nw5I
obMbpOqpEU1fNL0aXEPl0OGQUw1DX2/ypf6erTNx8CR800fHPnoN0BtcjZgyt/QH7W+LaYczkP5g
TtK4fXa8k+j5LbTRvPv6KP7yIiHsNPb5AMpzRO/iu/elyOoNUBkz7yksrUhblJPClzq8uFdZVoJF
VHg1KGRBN51UDrhbs93XYAs/Dfa2rqMvu+kTtDV5FObwxA5rqmD2RTyiwag8+wOfgC/PHMXrX4Cl
/8REMA6dEbhM/UtHNgM9EJvFy9DjPGHCkB5MhPuUyiuw7DUe3bP+kV55vN3vC55iUgqxYIHjUtDk
Z68cIBHTkapGCQVj1zHpgkS3NDJfJa8uVhf8iPhBKfxlm75f7qBW+FRK05b0sXW3Qe/9CJgseEMi
8oYDitGZ5qe0t1hSdLUCg5Qh/10Snk80JHPC3PrgCSIKrHnZaHJgJ4a1Gp73hkweLBSaBZHn0FyU
wu0PNrHwkh3qQma9bsYWdQkEECsAwjswzw4oeKE2QX6UAWpl5lXqbny8rRBFZ0uSB9BnsKXDJBjk
ZKue7yMgwOPjd8AEdlPOeKu+1Lmsc41vx2MD5+oCRYKlnp5p1bDX+l42ywbIMfi8OuehN8daf0WM
lfxVNOAwlAAJgzPGeRAk2HUiFKP7FIWqCth0hxWROMzKwe6GfdgE3yvUrTfdt/fXOfuAxIrGMtAy
pZ/71cFs/ZozTYH88W843ECayCq8YQhQNK8me6kBXN+yaB9zgBDH/XQRVbqI+W9luNNFSDzoXBzq
CAv7PAwxensTx89f1lxqH3XJiFYU53pj+IuQVV/2k8R13kZm21MPLF/8zUdYdQ57skYQyc7DCIcx
6av4MggZiFifgiViy5LS1kLQmLz9K65yF97sX1pNtPNgsfgWmRd9kKCmIWd1YDrmgENLqdrTyzVZ
HTrr1rDfCLxowWVpnJVZH6efNjyEZFLFuVFc25omkp8ViPR9El+SCHT+3mDJHd/S8MEbjsquVaBg
116xSOYgynPQ+pmE11r5mUK7z8vj00tir252kcv2D9O3+X3Are2IO6NcUm76rw/e1C81YtBNAns/
qSute17g2bYAclApDFjlFACMdg2jv6emSKsClfb9KBMMHVhqU/icNPF/z671EAXpZNLfs5kf8Q5E
+n2B29A8iQrR30VW3i4RKCWwQ002zi6otvNN0sJfWeg4/9UbeUZS/rjqJtSJxc6g7DpcLbA2eksu
3rI3RpmuwP0DMlyWZ2gXIlVXEeSZJ+SeNiMVbST0LIT1NeIMKg4cytnoA/qgV872oVkBwSf34/Ej
tHVXj0VI6Ii5YR8xDG2PtRXWSYsuzSOxeEtsUmDrlbGWY3DU9x3TCgv+uo66lUtOGXWsm5U/zQh2
RuQajN0130O64GCs0MgGRJTxaA2TnHstlIEZE8VCk1ZYK1soa5zHKxtScXjq8OQABfjjM2Ko05qE
54Hqugw0J4JSry0MvhD/3pqRFjZkpY+MxKWtVcMEG8FEX2fK+uEP6kX2wDRQh52dFdyZVkB62Ihp
r8TJ50RzHGhQpnL//UxFs2cUU5d0HeBHkiGLT/oIcN5Ck5NKwJTVdGAUhSljiJEHblkqi2rfz5mR
8wHYtiEWM8171CqgAPpn0TkQZlKX198jCeInU9OWX/iG8fxh91HQuEaA1GXKwLrMhOAN8kX5KC9F
9WdLD2jg2YiCikMlXiR+4ySs8QMWACZXLy4XZHCHVlayM+dhh2JMQPfzFy6Ohi7BKKDBPRP77f4F
nvdhpbmzz1CCiLykH1PDuTJWjcRSMqvwWm5tzrHvU5xT5mYYfG7MIBo2zqv7nJAk379lnNFdQnCh
wUPuzWxtQS7hYsYTHyIN/jHVQMBX+I8UqQr0q6syaT3OZHIGt3u0vNDpt9Lur+rfBhm2XNVJzOZT
QMuyninAMWQ0rOMN1oUSGtRsIICMdlf7U+13JaBiF85g0RBsZJpyzii5gvdzh6IvIYnGj4wB+nFt
GAxfwEeNGHc/6RseQwSzydY5cCEmM01UmZ4Qv1BaRBa4XoHo92367C9TywfKqVc6rLPCIwPAXwhU
GydXgOZd+vjcL4uEBSkhrty8DnZ3ubbTv+wyOFBGLSZQ29YoArXrSOIcLxNgtEJ5ftgRUw1tzVq5
p1x5z0oCWg0V/zaOrqDxpwIMod0xovTACjm+iafYC9oB8ozXG4XfjtS4FOqlgSpvI+8TMweufghU
n0batvdMsxZ/a/NGIaqCl0idVQXVvYnWGr802Mcop12mS4atgvYCzpCYi/gCBrSEzHtSdInilflI
ZzSYfk8qnE7ve1QVMojGzXNViVgCaUNROriXYFBj5L/4BMGuIyegwl4hoiHLKUpOn2pKF8pPgqyK
83wzChguTcDMO8J5tyTNLvp9zim12JpAFUMo6hg20l9AkFxm2NjM18NDWZY+m+p+fmFibqL3x146
vF32QGrszeKeVk9xq2D12lH46knKZcBR82YaL/lJ90X3u6nyoaGB43QMh1lloVHI4X2cHXD7tQJ1
gMpC2cp156ltmCVPdVvzXEOKoHFclaiZP68tgbxOt9Y5tuXjE0kZ0wP6VRCbH677u0HXiIpX79hn
G7/kvdZFEg2di+ALrkso/gNwFGyGbk099CIjw3J5dqur9nrUNJFx1G7emSON1+iAlTZ0d0OoIA/H
Uhs6JRFgfKdHQmwg+3a+8Uxoahes3eMq0NtAcC9UffFrxRVaDH2fJaX0g7jxJzrZPwelxwaTiimX
RVqn3IbbCrhX0psWEjvoR2FRc3X9CPQsOGMp7kzn1Bh8uW55X//zrChYSuw+Xxd9KYKbc4seZoWB
wsqplIGD9vNNKuceNYVmFWe3FZgoujHQ/ocBz50HRH780kQHQ6uaeOw+9dO23Tkjm1en0v3xbydj
wakVuJCER6U8RWfT7hQAwCqsaGuvZeeCBWx479/qDcYDXU7jCoonoINVcUVrNu1+4un+3RahyM0X
L3Z7iEsgjS1bl1HO5DwW1as/SseYQoQ7oQADYKK9YwcHY0Phasyk9PUNnGWLbYUnK8CfXZbxIii9
LFm3CnNYG37QK3oxUXFbqD5EEZEYSDnXhzcTAvWHgWjqx+zZqHX/KkHvCnqJbasWNMI+31JjoyW6
X2esZ2OLM3rw6KzQCRAu82jBVdUzsmY3ikj0LMkjV7xCGA20CgSGIgW5e1W4RyAWqN07gxHcWvoP
GUqhb7xBwAgb/ZVcfSpkfJKnVBi3aNY6OlQVk2iUmUOYm3K6UbKVlMW942G7FiNQk6S3uO3gqJK5
EH4SS4ezo7vPN/hgxj8menNgz9qyYxpWeqZbYk66JOlfMdsfSuLk0IBRNhtg6Ke+boJkKA3IIucE
8wNnx1NwWX/6S5d0LZNfYimfNDuMalYtuVrHCgcDmAPkqv+ZZxz18C9OXl6HL/Iytvro/suecvCf
R6GyHMtsS+oc9Y1RVxiTouSWiB1YFnHskyYsEiMicjsSiTncMvuANKJRRp1EzAeCKwVU05QKd9Fw
rVVkqhvSJoyVZmWeGNN7l4uN5RWSQNXw+VJXpp27RlKJzP9nxV/ZZ3lVTsa3oEjyxrdDrovbKx1g
sD1LBN6kMIK4hkfMmigYTLgCaZRHEPq4/WqpzZj5wiB7onV2sj4W5mDOnTSubjFN4qZxAP07yq9d
bpsCk9pF1FzEUiRFsFMomO/tlB4j8k3AA72UMUmmFczDUQes5H2AWk2Adp5APqbktusFbObyhfRB
fgh6wqRbSm1FeGNwTf01B1RveylfsQpwSdnfF3HpIsPqh3cn/lD9h/EC72JWno9xHVPgY+ri1rCo
p3k7c2Ib1NNryBSH3jxqYbAXWizctEzV+45RJUdxvZEhVULb/4UCtIOJg/T1v3lyVemwpP4jPWVN
H4DAXxxCG/xyjcXmc+mT/00fwfVEHMJGPejiJ62hVN3HI3yi6t4UooP83l5F3BIuOWulD0zUY6UT
ceMTokItFGPDHJmipeHBG5iSsMrByVBjrEjeJxD535sAskTqpJCY7WTgZO1IHL5MFdK0QHA3miKU
dzXk7hmz0Cxa4qII2cA8HQIKWXYgtN/hc9EAc7FGbVC7qZjjBj8aQc0Ehfoug2DLcJs12I+msqLt
GULE1J8wHgrsEWGpZ0gSbL7OLqISzweYkEk2iOvW76/l65GSp0NxdplxADxTH7JfsxTqFDvFSQ+a
zr9rSND+iOKLAdXC8Mew1WFoYtvS8prEZSPSdG9AUqbJxQW4OhwX/zsouUVYX5i/OpZu14JljcD/
pStYrtUPuW5hLxaSuA7KKKWLacozYEoOcFeb9iJ56+f8THh8tGTA7jjMVPJCMAtpaIjpmpFM+t/e
5ky3hufeMr1+Jog2VFMO2Pxx8nJwARwGdKsbX3NhSCkqYp3mcEK+HTOc8+Dcvps9PTV3c8F9N6xX
lJTJ/liYsOYNiNk2SsifxScKTWXSIp8Z/tdAxswWp0Em55CaIEalhF4v97BCsBVHaNeMgNFZSE/B
N3VfldqKh9eVIt3wOWjV/LKag/QGLkprKybzFB3Msxlob6fE5SQYBOslSN3VwX3Bwu5WlV1iTBjB
VWgAbZntObyFqvcpOmEtGShOpRqcGwAg0MFy2P3UmfpVbFMWQuTL0rifGhxfc3GjS0yb4ZwnGfHP
VHt8rFhSy2JDWttEcg60liQ591/Ad7PNmGbOVj/WDKYZgi/UP7pKnPAaRT3ULB7H/WLmC73ttCzQ
Ztpd8cvIUiTfzrLJ2u1iV9XCL9BmpinmMIdcMK+sx9G9gWhHqJ7HiS20JECTiy3MVR34qDbnc+4x
xV/cKfSMxFbMKzIJjxDcHUbgCy81cHideTzWPl7x0h5hSPV+bk6KAf2y4cW2AL/SpmHoeRG4pSoU
nlWLXfIj/ww+Vitxig+FJFvzmoHXCpiKcCkfSkM4PBT3YW+dSsy43PD2jSXB6/Pcpb0AYLJhwnbn
GISAsZyzKVjXPQirTNtMz1UL+L+2SlKykxAzDOkyrE0EZbsCLgfOcJXeLtUa8dXD8S/cc+bMc8yx
qi/SOqwXYSqrmCGETW7EmR0klkPn4LPRmRqKi/t9AHC+ZpNGyY7gNhksfC5yfWaPNKoFVKVbZ6Yx
z9k90HtmXk/mNoA1hKs925yXb8ebEBLrsnphzaN5TBq1ekRem+iJ+/xWEHE0th2je9AM+RkHG3Hh
UP14nYFXbyZYMoXOZQS9DOQj6mt9pkauAhoqv8GtkcLxWIij6qQBCxsQvVkv4x+pe7vpFfJsVMsJ
Eh8ToQt2ysj6c7B+owotHHzxaI4l2zZKrQpQkiP5Lyu4vLUSpwKlcds4hqamSMiGgzR2TFu3hsOM
rDS4Zxyoha2nktV9JYYHVzyg1FYfUHl1M4DU/deOF60S+5mNdV/UYn5KEPj5sbhDm+f0PODtKSFx
jHriAaq+YtKhy2BFbCugbmOsPAWcvpISjbFFBYgVJ2rygCxcJlHI7qs2EXvsvUITA9jghKTCCA6H
44LYNpzXyEvh8NUMjpXiAzxaHyFTXXi2DSnpFq+pNXb+KfD9gXxG7v4MAJV0rRx38GERVyceIUKo
JfJM7ysHj7W6NjBB6e1MfUO0E4Ks3Eon6lGItkQ0v3YrqFE8j3EgW4cXxf/ot1tZL8zTXSL3XFXA
mHKqFfjZHxd42lwrdf0kkRp8vAHHgA6q4kd7ZC/Zclfp9n6WHkWcGU8swBM/nNB/bO4ZvNxjhlfv
lmt7RXJ4ACvPqKYQndxHPbdNiGOPaiCwgtvok29Uq49OMTU32giqHuNQJqYkHM0MZoncrSUycUL1
xP6C31RYWqIyNRQu3VXs5tKw1wsqOiFAAj+vPoBCntzaXXhYY7fW/6YyqlGW5kznWQ4rOakHmU3u
DpfXAA6YjDj7dg2f1+tctowcT8RP43NcDjn3WEwToi+mFjnL16jBsh5kGWBNhZ8gd2hZ1KM6AR9A
lzzLtdWy7rhIrEPqRL5VA+C35GdtTAN928CVnGUf4lcQ+OAmQC/k5/+RgRH5s6Y8CG1MwvQ8CY38
FFIjOh1zjiKW1GES4P7fBY6ifmV1n9EnYaDgJYaByDR9iSfvmXAOgVAmZCUlPwY083Oy9/xrdVRB
W/Yl5fw8YZwTnD6ILTiPXMdfDmKoffiUhnYfWHrYPkbEApbvro8KY05MnZyf+XHSNCXbnRmnZ9Wr
y/tLEmFgiuaT+0Yybi7IjZT/w9uiZsQ3xKth3uLyXimK3x5PMtgR/+Do09jGAfKjQU3eCOWHyQ06
Nr1riqK4sZormxgCxUTCMlZ8N7UGoDP7pPhj2PE+xjOOvB/77xzKBy+6PJWbCoqfI8J/dT/fIXtu
XHzoHbYjDSevklKbZo/Szztiz5WQ0K38T0mgfDLLWJkzexRHRhyf0GDWc0EKQtdWU4EkiiQSAxsj
rQ8XydsVcOc2HHTzycIDMUbD7439hVfLAiURqFOk8qBKLA9bXCryn14cbz9bqOPGdAJcj+D0VtK9
Aozqkj4Ifcgdd/m7Uar12C5wQ1dl6mRK1dlOnCxz77lZR+H1AhD2bslWVfIr2N1jGjLtJpKPU2SO
NbacsupladBkg98j8B9EFvybL+iyLAWgaaLIm7rJmJqNgBPVEwtX52VDdxvOGznX1eTc5G+pMzGl
rkE3C1AXDP/vpEaBtXbtZF3+f+i9gk3Eh/5oPBBW+zvRKtZ4QfXTf66aP3G8+6695blr8rCvLlQB
XObvOLq2EuDxLt/pDLRBZHKqxl705Px5JSO4qPj4balFiUADwVw84ln+ItZb3OZMZy33tAUAosZ6
wcH7AamXeAcKNhduNfEK2s5G2ImN3u1mNDXN3soP+yTzos+ijJ8o1yPrJnYWK/PhSbrDAHMCzUMD
ozL0R1h1ZJ+1mm6qlfoAhZmYugUntTbJnNCTR0b8FkKD23lVe8/bBFmdF6Q8hj31itWSoHbvsDTr
LU2s0TKxS5hy+BrgBZ2GOZVstRkgB/DMkMgnmfczSSJmNhexDrbDeBC4pqijVeIxCXggtlQIOkRO
3VtIXjc7/5CV7e1lRbTPUU0cDO/wDNAtDSsIWg18cCjUoZcPTqr9dDkZGvARC6NUnl0APOTf0ieX
x2koBIrnRzjj7Iy3oMyqi9mMrPfR8MU9nLUdeaZDKz4VT9a824H192PR+N6Co7rTS7rFOP1SUTnp
kLuTOAXVVypfK/gh13dKTbGUbx5cSUjUiSBnUL5lhXwikD0kZPBlqkxGO2gdxysK3gmL8B3A9Qts
R+xgmjPmeCjvjXph+XIQc7zra2lUlbtP4jBUsNNtCZJ7RWOKCe0h7vO9Kw+gfdUIPY/buRXPG0/9
93BC54KTyYGB6TLdPGU/slU6uXJicC7vxM74blz+TWjn4kZ0DEV7X7ljk9Duac6VQWWZQ/Ca9G60
A3QVV02+YkCmnZ0h8ZdvVRn3xDtHqAceC4O53Z3Ae9CNxPNZYvpFFF+QuKeW+EFcLy86yS/XYYRS
vZezUuCI62te+TF5IURA3oQirrH8W5uzdHgdNbM9aG78A4C8WPN2tOTmujTmiHXqEBMl3w/5CsSB
+fUGLKCTMDUfDFUcjn2biNqapUcGLA6XoCa1ojFaVgrzNfBg21KwHEsR4Qpy7LB1MkRak4Cx6MmR
Y88Cz2D8p+eu4nJU6H4J9Wb2rLl8Fxr+QJI7Bo1zck/O9B828zt4LdocfTX3zz0P4dF6tMwpf2aQ
z46FC4NMHl+3Ggaj+ZrWz8NYRzlczKE19tcZDiKbkFYfzs742wfQZ2Bm/pbkKTcO/noJBF7/1bpT
yz6Vwi1O2GRrx/V0578T5rOWrrDYVgaahL30tuNWGzevfjYujx2AawBg2vwenBDBD7N/vUmjyHrM
Zus4K5jSEvbyO1hfa+XqYnU4F2TqwLYjvrEpKbW4ETdGlSqb+OR8uxw5l/Qfee9iIPK92cIxAT77
oUsjYRD9iwdp+VAaPWwWM9yDumc38++P1vt1AZ7NwatdQR1r3lwyWO0AwnUP1ciePxqUliiW+qxR
TEsdjPDwXl4lVuV7Xty6X+Te3OdWTtislleSC1gVJiVowmQ2RPiirwqH8Or66xXMoST2buoLUpPN
6G6234tA6tUAxF1x265ZnzfYFKkG5d/WgqsEGPdQ0OZZmaCOsp850JTk4iivIuL7n0VGFSlFhx1K
7gB1lYw3J7mUbbDJ9yPLppj3BTy17ZxQZx2Iodw/iHRWkV0i0T6o7ooVv5WVayYR74DNAmfgrrVG
iNA1HNmqZem2937oeTAWLO/5tyj3XjZgnfIHMKzU67ossE+m0lmFD7JnxOdl2fuTN6i/3xazAm2i
aQX5Tie5KWcfMdvko9U0i70ul2e2oTc5CV66i3NLE+RO4hyjXn/p0lKj+FnHVap04D+DtD12UDle
aa4C3JPe19qM2SpZ4yTAFSSlYjBi9OAANmoQ2PuH4AoGwjJryp2z4DUTm0ybcHgzjg38uyGngrRR
IHwVfBcd5+OYHpDnu4ckvRI39B+f+pxzm/G1Adjamx3FOdsTl9UiHqNRl9ALXiyf84n6+Kz+F5Hi
G3Bojx9aIaH8ow7gP67YvqmWaH33HYAx0t7I6TpV3WJ+ZXUs7DdPNc3+VRJBg6yE99JyQRgekKpL
5Sn9bxG5Flkl2yYE2Jp6EoEbeT8NNkz+ki8qCzNcvtLnRUEJngZIIeoSA6Zv3Yi/gQ+o9AcgLY5I
zgCY5yI++9Iv5F2De94hRlpIkBVHwayVmwsXyzzK1NKFYgPhEfIr0fLJmQt6qhxVs2iVReue82ae
qt+5rSWE9+xGJ+XG4LIMdf7uD5fFESBhpAYE3IzCb8lasniSoUUnFMYMuS326xuzA9QaWdLdKOiA
Wp3MidoMoAGR8JjQkzbulCNts/2EnbeJg9wnPhjCi866OhB1I6aE9zrwyvPIWqn/XVCwdMtAVXrz
2NNmuWycm3tYwAQKTxmUeCrUIyA/hBmvQ/OrybfgHuwdNZoaCKlvDMivouE3tVi9gourdHI5XOXg
HTn05zce8mFZG1H4S916bT0Sot1/dlwk6yGwfxoIYhV1n+YkOD10iFxIooJIDZ+I4Bt9r+UK28Y/
Am0b2V2t4RkkaXrQwty+iJc4JDCTgLnce/IFu1+TxElf+eC4RAM9fSmSBVL6b6Oj0zcPqdbJgAH8
EwZVLl66gTrHl3nB0sp2V6JnPbwYr97WWvoZNaOsqZLCgP/2Kllf0/22DZSXnRiZ5fRFZ48KHv/t
GFUiLw5EeMRR8skJQf+CRHC4smUWNV1g0KGCtNtEv4S5STp2DQ3NsxUHx0LULdFUhSqa3m6gtGgK
AsxWcxXHXM3ubLXn5wLW9MMw3P/jCPrTUdtlIMPuLI0LL2V34QY/7IH9mYeLV1CjAn6085oXIrBM
KAJWIOuwQEltV7XNoFz/v/0zbSTS/mcAMV2utg1LIfwV34OYQP1nwSw9ZBbxPega9A2Acj8h/9Sd
QK069jFe7bDMlI4rOqCA/Nv0tt3Qa6QPCbzd
`protect end_protected
