XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����EJ�f���,��пa�*���z&R0I��O�� x�kV߰��j��u7r=\
��2��"�Z���xЮ���'\30��\�)(�i���`z���hW�_/mU��3�H�_�`��UQ����B����{>acC�=$���z�"�MĐ�kl����Gk�r��[����4�+�dGxinz.u��>����=5���qh�)�9�o��A*��6+Y�w�[�X�tw��9��q����G
�tI�2��̯��M�G�g�2-003��Pg��+����W�4<�[᧱�6 JR��Q�����to�� �F2-J"�2:�˹��8�׺��C5'���3*S�������;aJ,���q��/�9
�*K�b�[�)*{�"yB�u�V�c� ��!���X���0��7���"�g5�"<�/�?���ex>4u9�t��1<����8TD�����Bѽ5��BC����\Z�<��� [s��>��D�(>�NKM�����fm�j*gx��P s�P^������:���֩�8��+ollUuv� ���<�j|%����?:J��h҈���hӧ}�����[�-����Y����;P���]���+x�#,ѭW�IK�����C��0.��-LkP�L���ZUK���#�Hݎ���H.� a�E�y���_��0r�
�n�*�6���P3�Η�~:���lPb�D>k@2�Za9��a��0��U����{ ���.W���)8����6�1�����iXlxVHYEB     400     190n���S�5�C��SC,�`�E�
�*K�I���5�tb#�V/��|�w�G��d�ꅅ�S�
�ш�]���b<j4�ٓ��pJ�ZXh_8��-#q����� �	Qм^��b���$&78�V�����Ϧ��X�&9�2�$������P��B�9�{ʓ��z����z����T��"Է�l�|C�o��5������X4���|?~��F��S�c���.���m^�-A#�BO!?+f�A��m;+F�^�H�H��%�Ȓ�tب�g��*(�B̾�丟�a��`��&���g��	�(#��73P;�X`�},���R�ͩR��4�%�����yi�F��t�u4�����:`��ؙ�W�kk�U5��TK\��=D-uɯS��y�)@���XlxVHYEB     400     1a0���I��;Y΍(���0Oyɬf�.j�]�F'e�4E1M�l�E�t\��G��>���e�ݡ#4�<3Z�����M�PQ=eh� �~�{���fV6��#��u��1�!=�V#ɞ{�����߱�I7DnF��&*�M-�L򭱖ݿ��S	�8"[�=R45D����A�3Xf��Q�`~�W�`P�XW�ٺ[��8�.US�C(��p�w"�'W����HC�I+�	�=[��<�>H5�Ѥ�@>3�'i*&p�=<�w�q"�nB�m���!�"�I�!���L�a�t�|İ�V/Ӫ�C޲o����w�i�B�U������d��Jdj�7!��8�Y�lҖ��{\Ii�2G$<��|�#Bp�2w�݇���녵���޵��ę���I���[��Ē�~+wP��D�h�H�XlxVHYEB     400     130 �ǉ�}{����Л&��o2����(#���Ewi'�L�1�[�K0*�!�B��٫��N�i��^/9�]Mxp�{B�{P�����>��do\����!n�`}/���2P� �����^�?i�f������jҽ���}���̄p�&0�����Va����n�@Z����[�[ �$d��%��[�`VB2���.�rKߣ>U*��q�XP�ڀ�o���I wF��f�V7�#�L4���]��W�8��1rI�r�w�k1��I���z�T6HNi�fZ���"_�YXlxVHYEB     400     160sc/���t��[ R�h���+��p"�g&��W�FK�=�C�eAq������p��$��`ZO��+N[�W[�\Y~���O�ƺ���2P"�e� #��9�_� �bp�Ԧ��=W<���-u������LF����~xA��w��lnvFc��tÙv	�¨�r���`�Rf@��[�|�y�~r�3�)T0.�����z!	����FE�?V]���0�j�b6���8@���;���9Ǖ²�9
!���2�;���<ά�0k!	���DNL%GԽ�e/�x;V[�y���F�l����ʟ9(���TV"]hm;��&�(�L<�J\`R���6��@��xPXlxVHYEB      3a      40��}���uR�3s�_�&�݈�m~_�u�`U��y/�y��Ɖ6������e����2 <����
