`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 53104)
`protect data_block
V+Wov60Eg2regMco3XLYqD/Ku91HFqCuMR7YXeAtkqw9/VpzN69qnYKuYnBqnGapnmCP3d8XU4em
MRx3EvsWrMqUe2z5VwltbDELVpmXtpiIy7zQlbRIaz28DuuecbK9MSsz59W0ywXdKUcHWq7dlu47
Rqe/VHr1xhnVJmaY+jZ48znPf2f6UsYKGneqChN+K6m0nO6FjSQe4RGM/XPB2l8YwUX9rr86mESm
jXvea4i38dndBGLZpPkkGYjKkEZI1doWsn+CgQ8mdZbGOtZW4RyM9pGXMoDFNz+MHOh0Kq1FWoso
vtZDnOUMZV+Ri0F+52DhCo4+zhxFfQyjDLVJxd3/MaEOaW+P5W3tCXLwNodlU+6UBXOssLhvDmp/
RPjALlgKY/XXN0sSCzQ39QYQTpCH0G4O0aPGctQFLF3i47fDF0hijoBP/u52sMGezaB5OI6y8i+5
G5eS3+gGU9uUCEBhQCXersR2MxkHyawfkmhpvfukKK8gvGSwlr5jSbXxQU2ZCpcwmdCEWIQmiW8z
roDjt/S9vjcqVs3fBaOOzCbwTqydTmroeTAe49kLBOAs0psr4zvCPjsXZ0dDLXtfWGJ7slP+RGUL
naLqLKCBkrzCtz+uCgWeLntaKQNUv08QxO33NFLAmhyJBf1SkO92QmukBEANTWd7KfXjPP28XgOb
IRbygPQq0wWcJadTdZlWxeEuVSy8YfQvFXp6gtxNvwctWLvTi9cGNylqxDJF4A/2HWThFWs3f3tB
S7d11qQ1O1PGcoM8jL+xcT4sl8bT5unRQz77OadQXyrOXJgEljm1XFgb6LTa3bB4qDE0JJuMyQ/U
1S8N2ZqqYwP4rRFDBfS3HV2+HCTGlJN30hQQ4kxUZuuubq229E1IZSAnKE9Xq55fD2F8iTrzp/S0
ZZc59e/MGHufbS6qwxARUF5+SoABHoy27G8Don+9SqWzTSicGBWIQiimlu3LltQy5g5+d8k3MlcS
yTDEEZJ7mP8HDaORDAJd6qziz+r2vBcNS8mebaJI5PJ4lgV1r8P+65CrNAvRipberpMrxbs+4wSp
vWeig924z/RVQmNfh6B0xnbIz5TAmjXQ1budxQmd5zV5AvykESXmCApytUFXL3Bi+LsYbW01nJy3
5F8wxUmU2+S6bohaT+2mHEc1Q4l5E2LaEV3eO/IY490Hkv437759/6N72ClVcgSBJ+MTtTlopG7S
41hmK+w0KImA+4ylRogqJhrizEMIIZkBP1MZQz8Hqs381TO0t2NhDjD3FVZEYq8T8B2wIDaK4cQF
EMCnOhpcjM1d3FbT3kQRTTeZDimkZO+vtEzO80ef+EieXUIt+e3XJWrRmCqW+Qa33w2Us44BrBLK
1yx8YNgvIP0pGrOaI8jl7dNFFPf7r1lKU9JrkYKdkRdpfTPqm89NAN5sJBYbreQcxdvqVQmlixmB
1F3jU9rnQErLhv2NaPMI2J0mf7WA2JkG0BWUEgexpDI/2Gaa84vdplTctrhFMH1UQ5IrLgpWp76P
XkTlcSTn19dtCGqsJSaAsd80zBnuVJhX+6Y2OOSvGmBCzB2h/HTc2gxb/wPNrVNPCB8hMHM68AiR
OowCXmJVwK6jfrp+JP7ZHSk4gJUl3Nr2LTEgNDzPyN7/YV5XYPgUJRFkTQvUMuHogX1eeiHlkCnx
egycS6Bb/gOztsC0iBrzxwZr6ljOApK0fZsJdnrND+Q2CKGcMBaVQdRHZ1WzEjrNPLdO1P98d478
bb7vWcdtsNELPmwyss6dz5kwP9s9sRzUTHTzvQPyqVuNn7BRFw8qPIzIU0ywmzwXLsLlbTa66H8V
FvLIDEpPdGRJdzrMv4mMWUUV8ImNu502HtjOSsDI1SV4d/ohmI6JqlNiqeGAPnXmO3xpl5BbiWqF
Ynpj5W8wHdWRPuALzmuC9g5dQBGPed7x4PPBXi/Qc2g30M5kRJW4hb3OpoDIp3H/IFdXUpqRP89K
Vx2enzqX9Ws6B84FyJZZ1w6UX9D9MhrBpmhhYGJ9k5v7JDH107il2NZcwFbLqrUQUVuUzcoXx9z6
R7S7qYPfbnElhXTGreF55An+dkicc/CW88Z4WXY2cXicc/FcGwPyM6WOIYX0T7iAuII2IZgrUbQv
2PQ/g0nqqhNGv+9qONYEA+T11LGJgXIynSo+90ezO3D+gi7aZjDx9Qr1jnZuNaf7S9xIWKaQNkEp
bJOBPKLLXAqkpzM6p1T+1m02JiQiiv1v+7n2MIlYw4+3Nzqar7XiuLbQnNY0L+KvGWbV33RKG5lE
6LcoZVqgizxYLLez9YwyKccxGMPVOd7aEZq0q8V9i49CziN6dab0TsdirjGBu/m4j2r++s4VoXOP
4Ba6/qkeAQanA5BpNMsGeCGKQxiw3/FEwilpmfyYAVFSf/LPnHaigq1aGBbhRR3qDF2AuWWyBxfp
4+0Q/uuhEg91oVcKGOOZgPVM6uMrAWhemsOzZQz2+kF53e5RJhO7m6UzjHFZBT7MZjmy/Oc/LREJ
rnNisWooxt4/3OILJke158ymBLPFP3dJRvmAADP+6yNJn8aN0ujLnKUNEPX1P7Odt32HcpkTkeAR
SDT0iz2IqaEVI+ZyEvzuSwzm2DLL2GJzfvkpjbg69ItetNBZU5pP8JhCpdNMtIym8MrF/eV2ATPZ
bHiY6dgFNrv1BYqY49ZzXAQOvBxbiK1sJAI101IiMrYgDYcx+gERYJ7PjtFcl8MuLCJ2hQh16mHK
908GBW5IMjSQN05J+QiMW72IcGSBWjzMzA+cxKFR1gBXJAtLSsqoSG4xTYlUmnbhppDCdLbLYCxA
aoxsih60kibmVcgLmgabQBd9TLvtoshiiZL0m0dzm9rZUhQrS9yAFF03syk8OE+ozqnMTrpSSNDv
FhBwC0DQ+CgUVCk6IGXZc9ikj0pjB2phRgmsDCUMefADQdUFL79sh9m8huRCwTQQD5PLWKhTwbWk
wXeimJY7TKKxPe6LCUpLHR6H3fnEy6yCiRRR/9L3ogaTN6l8aYhFL3Z7/FNQUvMuPUW2H9qkoFOk
gZpw3h+AotFqcsQv0HdMKatOjEYc5KQ7RTe4rglaRCk1KOnVN3pKDII6jR1k1xtsanYRicNbFUgF
U2djYBE5xib3fjLyuF36zRgBW+z9OSeNKXvlt4ugrgbpOIqiY5ZmXWG84KovS5Few6KVna6AI44l
LnUDx65LR4b5NkLoUxpzOsD30D0/epOYLIE9V6ic45UpZaL6eusk+2C8uff7GGdSO3vMBK2BcJOB
xPB6o8PROoPYgskXddXH1IjdDRHEoXMmfRBXmqEglZ2TV9epHV4n6InwU+XgiNX0p26AWvTHZgUa
3SJCDjWthK8ciKR2jfBAiW2ZJ2nsxlglHvwoC4M+FiXkGFgpXRdG0OOKfAIbBtupKx4euVINmo5m
cf+ATqNHXkXeQ+7Xm2im2Jrv9R5opTIJyqQf+1QWzr2snluBHM/Md9oQio0unK87dm8miLa4AVln
vR8dCO9E1xE8IuE3hwmkV72A9mPUL0biPHOc09pbFMhhakiut9qPb2fcOtZPe86yoFm3Wpj0J9VO
vArPCL/IdQqAGFLFg/Zm7cLyMUhI0TaIV7V2dqvApC8SNFBsTc+IPvvzCogsGEIa+0QTrbLC0P52
QeSt1dWx3jL5cURknJGlfx2NaQLbq23+DVFgiABoitKrM7pGKZDLzhrt1zDy/6A6ojFrBVwWT6oj
awbu3rY+e2t2EEDOdQqIS4fTfFQW2VOIFJeerA3r1YXwh0SkD/zt8jL4UZzEhJWxewj8P4PUK2fY
qcQZPpQ2jNKhd0FFJhF8xAoZ1jjJwddM2WhQJteU8WxcsVY8KfzknkVStV4ZwyDmTBPa1AndQrHo
ViP9Z8nfcvb9JfF4fiQTvrFuFck1tYC1rA1UxcmiDJk+HYfJavpcTWPAz5kAdaWVmHn5sKz7RqVn
bVOOGHtGCTemYbmDzrL9bLxdy1mHzhAJxYMhn+AoNk5SSFP1HPTGJYL8/fuAufFKahK0+jotRCct
o9Ptzw0JgE5PSp1OURLqXIKqthaQovBtv6UvzqKYy73JUa1ekijQO6tDpcmAT1wHzdgxbr96OO9s
83xFg1Q/7XYRatencaD8y1qewRb5eNI+8CXG9bLshx07sNIpsH/mFdNjlYdDieqH09EKEazza+oG
nLlY0tU1Ipw7UjEZpjeH1kipLwKhAMAGC/BkglZ/Wj0DW0sNNlDIM//8CoSO6pBap86w5kDdHQX1
27Z24mOreQjTafWbL2oR2Zq9jTu3PGtVt8O99nrOgQ0n1KiCPb6Re6EItS4HRVd6WQHOdckjdwUU
i0XR8TCBRWlAb1/jKD2cUoogh2E4/Ehx1KIUbx5Lkn1K8sCfMAIWXlHEhrW+hHWjdLsvJWch9Fbx
mJEQAuEorGUbS2y2YrKV0cUoN1Tk5DODrcscd3YcjyFE/QhtVscdKHyS7C9DnlTN+3RC0q0DLCXv
B/Uhv/kf1M5byiO63yhnxewTKEmUtF2KGryxElziVAiwqv15ezrWFEWzDq8Iqh5xTLnBBNelNaTY
mhh0PAo2/Wzmc6iedl71Vu9/tp9XKrZWCszLClLmJw5+ImJZ4nKmS3a51UqkhA2JJHLnhj+ASC03
X9/u96QSGS5UrNiZt8Pks0N0iQKdGwmZzMxsu7J/lu3FZkDZwE9wu2018bkH++LX3DktI3x5s+EX
ZP4eXR0rvK3oiUH48o82t254rSxeEJewR5zo01XhAt4Kk41DxYKeFsX7BnUl6WQn51/ELbGCzMun
jNdqQCrTik6mFHAqrYyrgbYKGkyvrcBU/kFy2x3P4t82dw1ebnhguCJrl3oJsHmmnKXgvaFV3hX8
ZlMLh2gwfRWHmTywlqx44BlQskq4knOiMksfUUJNiZpfsHlQpdysTWnWhL6qR7tK4B/moMtxJ0/j
kYGcgpM0WL40ldtd30QfsGghACRCcsigMt40fhUP0HXI00lfSbs3ns5YA86MsBoopQATEiHURll+
rq1pzpfiTIV8aQduHNo9dXJ6N8J/8x0P77ST7HtY5UOKQa0J64JAKEEQjlN/DO6N1SWPgce3DkQR
EthWUnTtLy3YX3BFATVfY+Q1w98X+a4pIxKL5x2u+u80btVn1NiOgvLS7zmzVziNzLwHB5/suiRD
rScBJNbEfaRQTH45hT2kD3LXl0yPI4hcKpYzBp6wruCYJ+IZfQDRAiu0SJ632ZAPDOeXRLLYevKK
PyyeQJc7c2/Ivf+0pQT/979YUryLrZW+cIbpMl+qvVjPtYpQ1qujcGzRA/6U/a/vRydhBDAkb3mx
pW3gfZMA0R8CRNOJS5FMYeIYWMpfooC5ZZj/8Ewd6AlyhQ84A/P6GBpqyDJ3REDyNvmQS1hzEnZZ
HtrvtnEIBLWeEe8zxzSjC3/1iXcWJFul2PnJnrS52Ojq2EahFthXAQ+S566+9gH09lM9VhUe+b+H
gJUJv365tHJjVuaX2CvPk2QaN/BRPIakSAoVqilDYCRjxOJd4k+GpvjljnbI39KIKP1IHuICVgPX
NmvqosyVnXEaMAoi/xNw7OntxvVS1pWVIVwceP4KzomCRODCHqBtWxxCOhvMNtlTK1aCUyGy5GBP
QdSG4ZjqB928E1t93G7CUVbnq+tR0iiK5d1uTWYDTp9eHWMe1fENs4f02lrmx55XsuaT+gxaoxnE
JH3sOEUwwQS08dfgb5hJfopSm7pWqfBCpSBeFbpGMLGGTxBPMGQ/DEJoS8pMV/peJa87v+sj+D8g
7RYnRgd2QhkQdHbSEwulaoTE5xSTOxNfkRjZQWp/e/s/fgvECqDt8+24vk5XaeLVE2lVCvOYIoWb
IJULVaBmZbAy3xYso3YiM5fNBML4nxFRV7DCc130Bxg4n0YlpD2fjVuBHA9sqy92OntOpfsny1d+
LaIc9mWqv2LXru/TLSrO2N6d88V2LEtzdKaCL2I61IJ/v0YtZ+B1bUjkON3H90pxIhhdEf+/S+Qw
GdORMWKgPcG5u9rpepEm/Z43TTHvKt8YhSxIEQT6hF/gE9lmWWXRwRG4RzaAXQmvxGtdhGOOxVkK
TenxgB1xIiknPCYidTEZxZSSQ7Lvn4bdhsKYngMAnfFz/Fu+QsXf82a5fGyLo95c9/PT3fDoTlD9
lJZYeZ1jBLWJEx1IPLZWFVzuG6vQtZnMii2W+DwK94Hd3VBVOimBu7qydu5DUuLLtyW9C39CLWWl
LN0Pt4jzKdWeePuEcg4pfFZbbJrqaSq/MWrlhZiDsUJz9g58a//Elqq1GF/XfZ/8cFLUUjaaNgP5
f41aqdP9gBcyKTRP/BJ9Mg5n/wi0aqxisgPNWITH8EtyU7rtU8bi+OxzEEYNzJsFTmcMirZCgqx5
jPcqzEwSyWI+2/836B9MUDL3x9e47w5xF30jC57H756zrqlRcD8I+KD/Ep9rmfMyvLyjgYsK/cd/
rffQ4lX1e/lwPrmfAPG0fblnJsQtv/261q3BEhJsckG+kNvgexi3JDeV804KluGoBKMjqjCJw9qW
Ow68iRNxTBjwNpfL1aSeKGlxMWumXN5tEN/jkw1cNOxeRueHGJi2H5PnvkeErvCYu19Asl7yoPUV
hwPa9UCXbjy1Wtt48/8JJvuLDlsylXUlIcFFgTtvUKQCzbXTgsXOkzzoltzjHxMV6PW0jV9UDlOA
3a9ZDDO1POnJUkiqV+/u2umP9FQ/q3y8kWSE9+SUEWQWYdEmNsSFK3w0hQUH95kyI3hqgNqsyuIf
LCN77cHzRiMxXPvj6xCiLW/7Bv7B4+RbvlEER56yBYczE13WBNgGU1TZSc1fP0g/Lp7NXNyPS83A
Le/xbRtcX8nPUbE0xX0GZQOpevq7HP2/CasTYC5jqvXV9pNwWwkJuLee0B/MCGnaeLQ+gZ/mGLOD
srxzy19La9MDMIyEa3wb7KKUhpgM5/xo+4YLrOaDj/BqVpIv8iBhZzYpxHo9PEnjWtGCdn38a47a
QZWLF6EJSeYXikVXBvdC4Z3ebGklW37Fhh43F9mNLLqF9gSb1AX/t9xvaMSIt+d8PpRFO6/XRROM
lyWOux/QDn0B98RSDDASV7471LuBu2/7FvUIyPnS25iChGp1NGV5sCW6AsQWBZ7j7iNSDbqHJsgL
aQC+AylCMXYOOTm1dGYqm3Znvyr5RWCoseefGvIM0SIp62g38pPJl+udhwpKV7smBtmdxIP2EzCn
TcFLBgywtbCIP7JjL25UzjRGIKJNj20oa3yfYjOBgCRFm+h1i5eJPiS0EV6HXaE/cH1MIyM5hJe1
rGrGLlh7RESdXvME7O1KU2E6o5ujEI+wb2SfBkvoXFv5G2dSz9x5Xbphxy/5+s0N0mcxk0Y5LdZ3
M96kqVdKXRLJ6FEIrbOXnE0reogHJ95pFxzHJ5CNPsLSk9neCXCg0F+VFNRbFLgioALYuUYD+LdF
zmZMGRk9np/P9Mw3owDHCVXuXdG359suWgX65VqAOI5ujymCHpbugNaWAns8aQwa6rHGuBW0lUvu
WyTVcAhVYnRodmhg/F16rB8aYR/WCNVUgmC+cbP81huHoIbSG6YZkbxYfsXUrmyotVNTocLLo5x3
WznohwPKE/19A8kCvps/m4G6FEaOzazWX/J8iwrsb0H9zCENRkxs/y5pEyuG/EQC4wgZzkqkchii
WaCfWCh+Hsm0uS7eHEHvKl0Ub7g0zmUgnlvXPK9HRfzpKSu+XgNaTALIXABgnrjgHsMb5N89bZR4
eiGhynAST/nAmxOrgx/xpBl6bDCbtXBvMZiQK2QChs68NrJr+XriOued42ZC3HDMF4a647qTxmnF
9pwF/QoFqmKNWXauJkx3dF/RndVWFIiwFdkphRZH5uddzsf76LW1qw9WYfPBaF8kWQiEmJcLt19c
8bibNkZfqX4I18Iga4OPGSEGoboNrZOaHSocLe44jJ0DaqfBvP4XxAOUMGK1F4Y/W5Yt1NoHlL8M
g/sKS1mtToJUyJRuPDnqBHSeq+K/BUB78j9cHlfm1r3HuH4Qcw9QoW1hhvl4nfnOq0JsENNU2a5/
xrcHaggM9TMVkaLkOzpd+tvVNKrTs26eK7rrR3aLXF+aQjbO9V0y0UtO28zfCZIObxXGUqdKwhmJ
G2IhIGR8gWg/W469+NyKHcdYGm04sELnJrpqL97NCjs2aoj8pxX/LvecMD38EYk3rHAHhIldXU7V
tXxeebWiI6r333xs91vXzs1e/DhbhEIF6Voc+IL/Yt+TuEFhRn0H0aj4+qwakSBsgMb502RmvaUq
a+e7T/4X5JRm4Eb3MLGVdD3iOy6y0EYbz78V7oWMCn+bvxVh8S3X3MNVGIveLMwycXW5pI2ZKDMr
BFgKc+GWPF0E/mlQWMEarLW0B+zjJAZrWiG6gMeD6Xq17FqkKfzsS/lpjdzjPj/5PBkSJ5XHGLQg
ancBhJzuFFF25JWVS6/SqvZZFYe4QeLdQkkQ3gsBuuA4Iu5IYg1kKZUrQn0uSEs29Zs9d96ZJbDj
Xn5auo3IwVrGpJipcGitaj0JTAK4ZMxmNhL5FU2ZvgGqQyDHtsmuJqw+2A3gJggEbm6/HUjOyRB9
4zTWhjPSPD7tbImjLC7rRaRESL/S7NpK8fBw3RXKBpaAaJmwW8SWeNyTNLPLtoe9e/o/PNIAfdmn
ww7KncR24hpUkVyM8r0bv+RN2XeynjsZ2Q6oXpcsANVkuxOTM+ei0b4rrEwdqTXUJXWp6Y7UlLhx
m3pk+OImlFIRYst3t0uhxPNyqOZR4z8TXuYrJadjFXQBFeowqCAwbAPfVXQayH+4B5f3WdcQjzdo
hFqKfvGj7kwA74jtgnc/QciBuqsjDWbRj60u9EwBBYfPEELttE3aatO/7Z2AcgL427I827ilJSdF
B8Goe0naA3PKJHvCcycfgoLPr+v6jeXXtwvsePXRWPY429+JO9QD2ERkbpvFIvYVwUTkZb5NMEpo
GkalTdUBOpzYigmXDSvHDpmfUHPddj9DWXwgaD+7pOOBiFz3r52+g3460NKhHnAOXyUYjwaKnpDo
GKXnK2TNNH9x/4V7fCazITxQkxVMpTHYP+8blG5IPGlO51KlpxzQkLGuKAIBk5D0C2bAUqVJ3H7g
anAKUAe6cGkMEArRp0G3zvMmTHuav6Io9vxJ3BOp3tEeyWlbjjWkOLaBi5eJuErcJ8TTzKYGcXVI
yxf0R3SbVBtB81jPHJI5jMGFXl+AcW8aBKlRFuN50lXaJdk4HhUYRLPnV8viSu1qe8NhdmRTG6OG
7wNTKzGnuyYWk97b2Dqi/7ZfCxEZ4tKKjazZsZNTvJ2Y6EZT/5Iu+PqUI5tQSA8dgNaZsVWuxsV0
5eyvq+/bzL5MxEBX/KDHb0MeiuzSS2RP6NDIlxT1mHMlThHjboohI2+AQcOzuHMypUrHuuCxEESU
8n81dvNQYoMusPBgs4yWbu42QHPpbiKrW7nSy7E1icn3lkp0fc3BCICece/Y3mt8o4Vw8tUo6Vq0
Y3HNIOehOTfckYTmTt1RSVB5NV8bq5GztdscYe6GN+GQ3QcRjN0TGFwCatXVOAuRGBvgkCsQ5g5S
bhKIJrWyWZNcrWjSaZRUDRom8ooK/udgvkk6hyCnG/nO9Zt4ZBUcYNDL0WHOsshu/i1wNGF6UliM
/cxtlcqeVdCFN8QidpcMzgZLiO9o+Vm63n/+7Vs5bS9b7WOqEll+YABVJD1QxQcLgTCZMs83JyNQ
4kW8TnMXLGynaF3FlxxMtaQWAGlG06yr9UpdTY+mlxLhWhT92BbWToldpzShFxeXXcFR/sO+nifS
0BUrSxLt1QBD3n7/p3QboZ+Fue4UQCBZDJhoA68NuAejNH+EJ9fRgRKr2ncJ4HunILO84iDe2LI2
rWNmbK2wtQBkTQ7XhXqe+5fbpsWAncCdwSsSTz5b7GHyHTKhF5tO1cjp1ZttNK4WFmU/FU2fkMae
eDUQyG5qsUd15l9XbRHnagz1uZ+dZAqWRIrrmcyOjDTmMKZd4EnjpUwrsLPQJg9W0RkYIZs5JmEg
omjiDZypOg8y785Kd8l7F+3ODL/BFc4svY8zeDdDSdJR19rFhlyAxgf9ci76XQIn1dYFHdBRCeRT
97yF2T2p+NaacwGW0lfzCz60pJjEBH9hDW7eUkWd7onlBWUZmcw4EBElUS/Fz24cNdaAEw4KH8ks
As4/93od6N9Ce+zR9/zUZJDReoqVRNxFrCEk5hjC1y9aOYqcf+9XLDM8WTZ3B3qiSMjw5Mnyb2fK
GpYN1P680EoW91X/leAU1g43nmaCU/HFHvIhHkD566SeiA97RIEDEIsHos7kM6qpNGXuIyeiYhlV
IbjD7a/LBHMkA2lCjFlyZE29EKNSnx6g9qtn5CYSj6qlwavlCPRDWShHvqDk68BnUCoDNmsfBpK3
XJQulGGtVc1ZH37lLQDD8TQbg8dnPJLiNLec4jYEnqAXQQNwXbs6XcR0+hdV8yZiQ+Cg455Y95Sd
NCFZcXjwmm+Fe+kWb3HvNtX45+QCgzNCpwv2HOVDMeV/INnJtkhKiB4SnOolH2KODEN1xmF7P9qK
tr3AWYhOSxAx09jOGOV6IISJqp6iufEE28IJUsThUpCOaeRNgLY68Ncvh31eAa1Su7s6qXYVjgHG
kWgaJuJ4RtzifYzv7EIaY07+t6IImUna/Rk1gsTR3gCqGFLJlkTtb5hXVC4E7DiJUGvBx5iL40YI
LOjvLo5pGkf61P65jI8EjdSq7koB1oqyYK+zeaXnFHx2uneemGOQDQmErCri31ZFRlM+6cVI9xFe
jiVSwSDkL2iLrgYwaSMT8d5V4NXVi3xHP6zgKBDQnDLufINFvpoVT+gusJ5hQ89rfp7lBM+kYaKQ
IyETxX1IixNteX34pCdl6Wcvn+6lvcgmbJmLMWGNL9WjnWYkRY/U3YGzcdnVQ4Z6ydOLv0zGSjLl
b5Xln2Hds/Rh08L/C+GTs39yKoNZdQ7bv2kNeJh/brsNSnzgehvBrxgD867ueTjfm22voMKShP31
HzXGwrLEZJpLUBfojhsKSiBzgBX+lTxFog4HQjfk9z3G98ZYUscRcrfYkCJtLUZLzHH+dq8o8GvZ
WJRFtuUA/fwh9rnm29JmZHMG0ufVexOLY+ma+rRPrcgLMgRa4T4kgw2tvoBOoqs7Ws4gzfZFlUxx
LzUju9wFA4qzCcXmK3BhuTeB2O5aGnxHztyXnbk9akreuwd6zWEzBRwKDA2jyJw9W9gRDUVtMfCw
z6T3e9wrg3y2lIrhTvRI3/+hQEB2GQJO4M5U6dpGmBvqSmqljJTpqozRGf+gAzL6LC/Lnwvi9i2k
2VMDhurY7/4UlWdpoQ/BcMOlUTxlf3OeRKEc8xla9+soifXq5M/c1AHlJKuIutjsAb404pQLqB3C
wkozHOK40dvDiUkiw00/05LLqhLxkOOOQVM2Mf5uRpf5P6XgVmnh5HhOwXBUQI+bAA0+o9yznR9b
zpJ8XUuak2yCdO7Mt0EtLaLH+DrTkn7AshODZZ2nOLzIC1i46HinYDVZjEiqGVAOOoM6w1uvo9WW
CXQ2XrNoa/BB/U0az3bUmdeorMtWH84Mm99WvRRqDOdJG536v3ZKJErL7xsfdzyq7lg9WuV+0eVT
E4LUyAagt7/JvYOnLmHKUZiABRD7tpYgvcuusI4Vz9Opbot3P+nHZbLyJZhzbFFVbv0KDKX8EiP5
z0p2jiAU4OtKp3wD5bRi1Vje6yXUIf9vE+DWgp6LWn7B592/JPmQRCNPmLRQsSmwI1wEKAoLNvg1
3R4tcM3K7t7NkYG3GkIRvCRS0FBdkHu/13Sgj5Z6pbvAeM2aevPt69W2C2KsDIZnga88vAzyPl2L
a3MbaiDa08FvqIemNFyrOmA6Jrm4frdQZcvwjLxkOrW54GXqOlQL/8LSvwUYJOQUtI/rMUrpU8pT
FbADhscWzsR5OQdo0RMub84+B283Njw/PB8U4mABj0ZXt5Z4IP/5Fp8PBCaMKmePH8cpZ2D+5ZZy
XAoM+xjBpUPjjXc2Ncb4FO/izpYoPKeoSkVcqcTf8aHTDKMVHWt2wOWAlSDerjoLpMWQ2sC3IRt2
k5CVuvMLsKZPbSzjrjROuIbPjdQ/WqAW/1ne83x9nGV1JbYhDtVHHS6CAmnT6PbDroqMe7JSdiSY
Giym1mdYP8OGc2AD30HpZvWiA1N/alPJJalHpKz5zrB+9grwa2s3yk7Vcjm0MTkM62PPk8dzyrIY
tSt6NxA+0fpyJX6KBDL7aFjzLVZprXJpWrelwIc6WDxsZtsIPXEj8q9Uf2EcIlTIukCYPTNL4kza
6KupQulR4lvcddg2RGBqiX43JBWpVs+z4b7fcq/aJquid+I1yTEVq80apJ2IqB/FUP4v/igKFdDY
mcnmpP6O/A+yuzO6cmgO+2bVyjynNM0M9vy/xKqTpFgrIMgKCJSH+sVf5LNyzzajTJBcfgzAsZew
LxszAUxhr0iBrzj+2k9OgsfQf+qZakPE1Fl6dBF4YuwBc6cZYnCqmMcT0o+mmVc+tikE89AfGZEn
pA5tRqkb37BVYY2tyoh4Xj8AJRG9hxXjm4BHREzT1RkHSUTRlKyHmw5mcrkGfyV+/EI6OB97Jqzs
fAO54eaB95qE9Yf+ct8x7UELUaiCMKV7X8TXpRCeEkGq1GIBtEL3Yi909116L01/UpxjORBllokb
BtNQHEbECBV81uFRLZ3/TSCTqvF2nVCcgbtIL2ok8Fn9ZuSBI8kjTYPd4cuOzybrbreG3F5tJNN4
8p9f5cKEnQiD3uCZCJRW9m8Ga2L1kv9EMXTCNa5k42+EFyKAMBzGKIyK1CJ7QKN4+7IhcVakuhkk
GTVGQfgiM3WLfSw7FBDi1VWT8PLsKPXAKRk2koTmDW2DrLrLrnc7fHlPVCBZLbkp8eBBqt5aSWzx
5TlatsGFhe+cwlFohwVPBeh5oxE2VRMURTI57hvp7qH2XITcG9vzenEl9IcyU8RMrqSOU44ghmHC
HQ1cLYQUc7zgk0QIgiRJd5RC72ROQFrtUb3Geix2/LsEYyA5eUb2k6b8avnd0HX3IbW0UCTxExoo
xYmWVrQs3EapGyrpZeQWDV+gTtibIfhRv7CrjrFKQjlMh0jL5pGAdvb4qqa2mBsYRqFbibC6sbbV
rD2truogLMvB9uavZA8E884eRYaTXH1hv7G7mE4PZRSCNaz6UkoALDpdklzEekmulHoYTThTdHo1
a5ZOU1NAyuc1Gxp7mO9C/9GyV0jlpGxGyysqzhucimHSoQzPjBe2ZOvAufuT1KnAszx4v/xoKvRG
cFx9DW+kDzJY9eYkVyVxuMf6+9lGRcSstppmASpbiG38MZbTwRTwI5fnF9Grug2VnXR0Q+yu3UPI
SmubxvLzdWDbG4Vlwb9YjoiETAeJ1hZT5tGh8Fkqs7sTdYmONyMygEB3JypmrLPXLuMqmgUCDv/I
H4+PLQ4w1j+MEWIdmrX93YqWMZCkBpXttS4p8cAplpDWTvPVncZS/bFt+hPeF2P0fc0XISuhfdaP
Kq5mreumE6l0ST8X6kY6zXw56dt8fUjg0TqF3hL+wJDXJCs4m8T3J+ai1fQifLTc13EFBO/9vk3e
YOlw+vKrQ2MORaiJVf8nP5atxS1CnlNR/G8OyDG6nk4SgoElQWmcr9KpqZH4+narcCgeNL9Teivs
6tr1PAuDT23Jx/fyc2Wwc2ZyRFohAhy47kjHOR5QrlWGAWa943qQnQNSHpEttkf3ApXTJWBLpnkb
V/m0nRdAakfIz6mojCdmvKd8jAJvFlDfSqTyYluVHms9DUAmKeb3WJt4Q6x7HbjZZxp08aWEi7h1
jUA0n74LxurB2XWKP/6i4ipLWz05s+pFcbJ81z+gOKjpy1lRQIP7x6MsgO9a98lg5pzWzCGm1fWO
HBblr2EwsT58ZslHc03MA9d7yfHPg3EhQVw8YL4mZmKPxry0glh2RqRdva/vopVf7OC4BRtFyZyg
leDHeDynpg1dVXbTzARkddxbUVpqrzs7fRqbmpHgv3NOb/LLO6E+MfyoBMqfUy/ND0bAA64PIUoH
61uAljeKqecxVajyzxXVlBzLlxv1jikYQilrzFkPVrQIJ2sFsMItwpBfpdosQAS+VyJZU9YjeMos
r9C9LCQ4Y51FqAo+/6qQjNJlWdRmT1lr4Sio9OKLmWybtLjioP2oAEmgYZQQOLyeks4qc9NJK/YL
mK/jwxtqOp+q+oquAjqWhbN6a4RlISNpw4pUV4nQCdU7A8KqaFN8LwjLjAFAS0MySdashRfQVFfX
0v2f0z/Vi0AJpEJcI6Lq+F4U6Mh1MtcXrh9bhZkRF+lyyRuJwY1/lcJoSjIVyt8sLfBOjptW6zZk
Tm09bUcUgaGaNoNclBNm05ZIio04bd4PxWvM9TkK4w0fNX3BDrRyjKrbdzKhxPlqxVT1pf2sw2Eu
1srCeJOsxWN+gpu8lfeaEayiMndoD7GCep9vPr6SR1/rpga//DlBHL1Rf9W8FLOB8rS8FyPFiqde
qvaKbFN7gpFHRKBpWer5eZOtGgG3kjgGdekkhCk7Nt5uj5wRlKEVVn/VoV1ixoGYz56RIGJDmSvS
eGqcd1e9igRRY2i3V9v+/fzeuSfhfO20lrMJG4iIAiwti5TVShh3kfBs4GI4s0ghV69w7w1agACo
ko7gcYJmm6vqH36lKloc/DutO98Mx64bAYZWYXhTaojadhCE5VExq3+N/gpWa3auXYxf4oCyLVXB
tYJ7q81lnIeJTglr8FZdWUVZgOKS9V9ep4ffKu39jc5PKVTdcNpyrX8atqxzujN9m8xLJbxlQVum
5tzKyfSEM5cD1T4NQVx8HsPBwpUs4GtsMxMEFG1hpyEAgeKgHPNZLFmywCnvohCzS75iWCj6FIVd
Cu08GX5Sg5miat+yJG8P8Tov/n+vcyWcXK/pLg8jP8COhBxl+Cd3k9JTj2EM5mlfkYhn61qEQBNh
MEDQIfh3HYFBunuIv7U0FBynaaaVrhjoQPsQR7ZmXllxp8zwM1dR5IZtbzq/JmiTspjfRpfk4Fnh
/UNd+06/Sj55WyRJUZYou3c6xmyLjzbGFN2RYTM4WltYstdfaybxPKGguVWocnM296HHWUGZGFvi
HfewJ/TvBnIJTi5R50x3wN+m8tCQJuFcfKJbvjyteinZT8rOhtyJoSXcHRGf+PNEg4xz2B0WmX6Z
hAos8hzbsS8sI+co7jqw90oQQxSYagse8PlTkMem5xh692x2FP7JkOxyQkwUqLOpD0HRA2b7JaYh
KzaGoFlmjPiUTJ/N6v/P51Sp7Oxc6i5feBw5cysR6Z9ff37vrtiKwOq//cUJF93h2L8SLLSHs48h
WEdry38Z9QrwDU0f+i7WExwmwB9ncF00tvhF7O7w/ofo5Xr40w0JfNTfLbls7tM7DRP0i6YbWG4Z
rfFIJ9AolMY0u5UjxTC2zgnf2c7hNBsWtX+SQzyIUcZjUU62wBxiYoFZUgHOeLobAMbmig5KfhPW
k+3W10reoK8SBpqThL3fSrOUWCzpOaydfEk4c9vg38DdX3azJEMI8HHlJMO3TLx7u7jsXVmRZN6v
1SK786ij9Rr8fN5fY0ka3y47rHLs7PQdpr9Eu4WPSN31EBA27je+0ts7hW2mFZdXulR3XVf/3nve
i4PYvS4rOtxM29DuHJt15AxyxMADLbBF/m81Ru92841a/FDzafmGA93HaA7EH2U331+Q+yCzavjc
npL17zAFcW4dqYF8X12lYJZha92UZWPi+GE18ZtM+XTNuPa+9qzu3Eh1H9JCHcO6wCSmbXqdgFCc
XNp1wu2x0cvMO6rDO4S/5Gnjcn+tjWB/s6rdrSw3NmXhR0bFFd8UCDKjb0kh0aoaWASuDCV5m2G3
ILPdbwCd6ecTQnoPACJeGOGszujuwIJJCHvpL/Wa2Nre79GIVXSTt+dYLKaq0W/XWWGWe2GEL4at
PGpuTQZAVJYPkEDhjXnJiFRefgQ+dRfH+lIJ+apStJKzACYxcLw1TjHcN1pnxqvpbn4xMGP0kBwh
12TGplb5AT/7vWpaCfCab+zx3l3SIcOcUJrJEQQoGds2freIffi7XL83KlV6nwEo45yPwB7tTL3h
PLqsiWzoL1Fd+d/yUjgz5wd1OAUBEzTnk07nVA9+1i+8pH6Id0LiAyQ91feYjY2qXQyQasFzygLi
kRSxa2bZTBn3w33UxptD7fdMxA7xqgz7fmwm9yqHhdO9rteb31mECtwYalx5xd0vmzsatdrRCy94
qqLdFOO3nC+11Mo9qCQ6ay+P7r+JUqOC+qgXqfu2t1SqifIQ1YbOpx0eZ0RtthMwcSA4N6kVJdfv
Bz4NoWCBKs58m6V8aXBdkiwqjnoXeY4mTvZGoOuKPlizfncfKfPbEvPo1gewk5041PPoRNbpg3IN
RNVesyVQndeqcF6yaljhq99fjg7SsEQxzf/+xlJQlMSLGpTHbrGynnNjHwVJvgipuFAnBnDUHj7G
Lt2W7u8f5coIBeVa9ddbbD1yrN6rdrhNMCCr+EWnlsBDZSGQo9ZwXm7ZsUWcBhQBrgv0fVrdLaCu
Zdl9PZwf/Z4FsjXpUyj/hsjkUdHKpaNFwokcu1NFDJXAAtSPyHdc/wdeeObJTn1C0QfmqpbkFP0z
VCPcFr0r4OuJLmBkBFf9lKykbr/IPoQLAaR9PpQpnfidN7g1dwy4g4XGjdE5GauXA5UQmu6biu7p
2qdkNNSG0XxKFF9wjSD6405m1ugHwzUdjFlEJXXttYSlNjbCUYFsVXVeVXyxR9Zyx/7RhEoLyjiP
mkM7VN2iDB+60oEC0Jk8aMWQ2lzHyKPbL9pVaFy+kJ+NAE0KdfbDFxtw600Ni4Mn6LaAuvXq0pRz
mVI4dfSnF/bW/Yq5OUTk42x6OSVhd06IidkrlgTMIXuf5NwWxHqyq+HfwvknIvUuKgiUsKGn4I/I
TZ9NCtzymppAObu+uaM3lArntZ1LsdvgKxEutfzhuijJIM5fRNk7cMpWHN22w1Y6oax9rNrPE8Is
61ZdG/fnVAmFdwwyOvF5inpyDupSVxNMbgo9h/j76p6kstqlxIbOMt7sdLrowpqVdG4zaM7n+kat
+Wxo2j7t0cEhWK8+DfkL5xoNU/wyZzwhA63uYpZcljh42IKI9eeztnNvUwaC6UL9hQTmQ+S7Jv0P
aldj5I3K11AA8IFpaTRDZNuuESrJI6kn421b4Z8W1Uks6DAoivmw2xmUwUrEa/G9LkURZ7iR2CrJ
CvhY99WYDRypmdGhugkwp/KzK32neR6KyS2aVlO3TfwqoE+mkt4tLPUtydWVFpAjvhOgK9A/SA99
WiMBnD8XBa8gwFINkIMcz760CPlMBl2OdEex4istw1XUORvr+v3yqIUSt4k1MrdZojv+E2+lsAm1
Ms4Vm3qgobRTKr8HOQuHc4GzqjNW1YoEMBFWM6KDBNp1Mi8VlmpjXQuw4PyHGZsfSWofhm3kNtEm
REo9q/wh4Ky/m9kfohjrcgTue0SkMlZUmCawz+hebPHvmOkGoIsIkaD+JEXoRRb511D9qeAb8pY8
jhnyNZhVRyENvNxCaVMbG29PJWyO7adhlKZjqGtX6EKe0eF4D9tkLhKuxZOVRhoa47s/46kORG0D
6EaMMp+f2nW+SKROpHQntA3xUYcFDtpWrw87G5ACb8qmW+DgKAwpbphSsgsa7L2mVyJc3/j7s2it
ZBfUgbPLMMGgfvpG0lAKZ3o/IPDQ1GELuo3tvgW/IjkTaOc6NNsLrH9hBp3S9OKVD+VHftbK3Sz9
ZuHD0l5oY5o1fwRFyrac5Mkjbwr77RuJhVmteGaAL//QB+wqnludWxyw/zECdc+32p0T3GixkSIB
SDYR3t90DaPemTOCF/aA8JqP64nVWnAlAvXyaZHVbc/VehT2n2D0kJ66LUdZEgJ3N4znN/9F/958
5kF8W2UQJwlZ0drxAa0oC1y6tfjn8q+5y6wsK2QFuQornVboOO5Ii+qVDcitxQ6UQjI8j3X5/xlK
cEyz6WHwZ64aDaQE4BxLLzf6aYrxxuwTVaJVvko4ZxCg2Y+jw017d54GFoFtjxIN1GTFKunoMsas
j+PDeLsMsvY7iMH6CMJdac9Bkr2rZ+YzZpEIy3OFUGonBvM4xzRgdRKsoSXNnhJuGEhM0U3qlrVi
9Okh6U4WuvJoQCqwrz7vRP3zlldQHe5onJRdAIa1ESCyU3O0vH7oYbTC8yLuTRjpAGL5Vkc6rf3r
u093ny0d6yxVTqjremVMnaST6WpqRqrYZsS2UmX+WvA6PZKVfgsQAtzefyRgVepFAchspT40R6X0
85G+8EQMs2AORTBbcQ7TA8sMbNj/7wg8dRRaffMxm9dmoh3UQjXnDjg/fQIwZEyKTz9wnKRBm8HJ
ROMivFoU4af0eF8xvBzTz/futuGf+VlMAXYYsHuRhq+K1LqpmZMNkvCQcuVaCn5ZQ+U0KZCbr5yy
ZE8pdgoaMNhbF+JsaHlGkGYt43BpAKBkssNj4futcVZbmt9+clo31IV9SXQyFZ27oOpsdWD+M/Bk
heFsf21vIAT2V/G/emLTfMNGJU/KwKYWRR+id8wMWqTBU6FRpTNwtBuXzlFcuaBPx9fKhVfl5DqC
kzMATIGBoLJZB2Vd18HkC1EDS6i8hu1FKISB7ynox88/jqgJY01hcs9+PbmxCQDGwMUUy8HjQJ8X
Th8RelR0i9Jm+VZfda/81GLYh0FV+5yEBwsaV5smWumbrC7gsAAGx83k5c97sROb/njPj4pxxt2w
U69AME0hKh6ZuTyOJD/DQLyDh5a0S/qd0Y2s6CeM5g+AnELqR9MTBzIde0kNMDZ+ZxmLzo/+j16H
yTLe1DlIvmbInzEZBs4OeuW+XKECvIoX13nTRs6muauPR/BJp9QOSgDAZFkHOQZWH9fmMub2ReF4
q31Icfjej2AeNxUVg1BakJuqTdqaJL9P1SKqoIjTKRkKZ96ZLDqjDs0PGjzL24Gsm+S7Xqy6G2zO
DEjbsPLzvOJlVqVtD70W7jjOMkRUSAKhP2/LbxP19nusU8tvdeBou9mOszaRrjHfd64VnOg5JoU1
gGMQd2Rx+cPxnEiHM348OdYjlfgZHl3xF1rGGU5ne/ZST5nJ5rIFkn3gOXWOxoZ7yTsZJh/uoV7O
dF/WaGIp9+HgY4VI+7csjgyZ5kBzWpenMds16TY1Ro69+m3ew5Vj1l74Qs5SIA2vu/sLuTrvjC17
552MIAFnm6LBgx8gMkDMKGX7KQwy872O6WEjpjncorlxMejsuVc6fkFZ+afOXzPGoe+dwgEf3BiZ
U2eo9nIbcvCKwbq2eOnc5bEBuVEwXJuu4dBgODzzBEFPOmd2VokPyCfDqiybsBjM16LwMbuAeIgQ
dcMUF3FSuNRikETo7ObKoIuahJb3fXVmk7JAnmxgm0q3lIesIVi0bpKFx/nwnksOdbyYjz5yv8y0
6NzMdD3wBkRX2uCJmtXhneR/BKh3uvyFxnMpmJYdzyHtDa7uSjZYba7aZYTkZ3zRxzObaOOWzkAX
0zgFHwLaT5a31kxyTT7UALynEFfCOkgEVKvdWkV3RvOueS+2K7l6dfB+lrKsNC/zC/1bObKOumAS
2x033cf6hxl0RYEabV0FUhaeA2HH3+1pQa+Km5Y5/XiRMnWqnrz5ucd0YkTIQT0EbGHNEispXDmM
by+/XRfu5iY9YdmJrfv8DciLIUEYrJ4O08BeUB5qEvQs9IdiICWYrjCPxrooBPgs8C0wbzp/a87p
dwqAG7qJciWDFpH8fpKjQgmN/X7PhX0oJPRFl0opTDmZ/+WVigtOMpNdPzmPPDHkUa+7FbPpolbm
MSiL9sv231xlS5vzkdEVqxvJneFn0mNroG6YIuDB6yo8JwDpdHeb7DMb9gQrK8r2VM9m8d4G9yBK
PlNjJgNyjd2UKJ0ErITiFrMqtppAM2QzJpe91b99ikDII9XkozUshpIlGIo4kvv4vzaGugdyXhnq
FN0PXTHGdTn8vLYqOzrs6pFf3a+SqpFbIyjHuZDHvIN6DB30jCXcxT81dlpk1hkNnEw6/oaYcQcf
XAsQchydHkO1GJ1c80WBzmDz38/JPqGo32n+hCj91USP+hbXjBPIyXyWowlPpdSlihCOzfyl0PL2
oyYnWPyAlDSaUr8UXpZl7lUiWDo8yVeqZ3ohMtN/w19NwTgObul2VNIz4IHmHIsT+hygHf433lyv
dcA51wvhElwlSWkPB+cts/fcr+VhGGGcsu5GPA+ha9w+monn8SQsKavZ1CR7EW9aUq3cI7M7iZgv
ybuvBuPuIYt5ZgZQ6uCJ+BcBU+ZcQfIlDCnW+614zBZsTSNXyKAhpkzYbGAo9DwSlIxnqw8h9JT3
GMLl3J6h6ZepjYaGxNAP+vboCJwxun0WTljkrcuEPmJGjKBP05+05jmeKXxFCL4yxWQ1owktrJ1T
D3GpMuRKGlNF5p9BABnuBk/Ddm1ZCgU/9RtDFRy8OGrKPb+ah7nKYYWqbrrinhynvSTfwQ6t1BJr
FwIz3ih89XbU0JiYw5NGTpbU55TeoThiQr+ZH3ApV0BxD/D2KbV2b9vdrR/aar0GuuzCnprrH70Y
5repkNvGX9QuKeMvLGEGQLPptoIyPFVttKpyT7dWH1rBg8qHvZkmATaNFPiBfRgI/b0LUFVft0Hp
r/TKHwv2Bgt+UqhiJYb+oYpO0eaug9r6LFGW01T1kgVV2VAHB4pG2p7gpS0UeQKW66wGIOwcity/
Nk0WVp2ycHiNQjeoB7WtYKZWtP8zqs4irakX/p9f1eiuhWmjaZq7jqne17EHTXgTCjj0dbLYPPaX
9Wo4gll084jTtUM6fWjCNGnM/crjywWf1Uy5PbHZVjbBK20fxk34tso2sRRH1qBgBN+LY84zYCDF
Mmm/K5eD2WAV7ZcwC5JdZRWTs+QtRX5xqJrTBhJ/q6fyjNvMPrpGC2ibRSAWy/JeJre73p4SONHn
9IY/qFIgRB8gmfohrRkFZsLvgMdbVm7TgSdxXL7iPqmjt9jVMKasIXhedwauq2fn4xZYbw/1V2Jz
33zK5BoRrsijqdoigSVFt/KkuObnH2xQKajQRZegzqsncWzCEmob7FN+XpX3U+33vjF6LHoboSp5
QYeJd/hGEW5oBcnhTfUkGjNnur4qtJ6LuH0/+FbgTshEco5y2IAdGI1fBsBTeynLGwo1hwyZCS1v
DQMXDz5w8rzn2rWDzO26cHGqchlM2JBE7Rx4ZwFXLNXBn6GTf3dlktSrXa4hgkNWBDlROpXbmMBa
Yd/LBo/dS1I8/diMw4VUlaOpc1pBbVEvfZAK/qZyUbvjXOzoY0E3ZAkR4PbYay9sypj2fDp9oJvH
u7eQNGM6XhUqANXVEZ/zfplhj4ZJKH+bqu+Fip6MOKCnS3LNWcXcTIEG421QHbVvbfjo9Ec8rlQ4
kF8YMMsPcjHoP3vAy/7u3XxtnlJ2/CvtZdseHysHaHfr6EPVpvGZ9LLQt1F0qynHpPd9Hebq19/r
sp5bSAVTUoZ9A4t+ufkriUkXTngVBDvlWYCjuZztpGiEDrKP5V3dIdG24AhBb7cfEiOv39VJQuRK
6x5vzu+ARq2deIx8SoJW2g0bOTQpsqe03J/O6dI/evpjJuVbLUn852Yz14yOmhReUQeiA6/uBxH/
ZfjqyyCRl6g0OhuW8JU22tMC07cyHucP92d7RnNIu6GGiMLwVzWKtnx+PG3vjKUvv+caipm1FRmC
7VQ8vLCnDaM42tOOHnshOxgOfqX/p9ZwqqKkwAlyM7YJg7o43g5cGL5EO1UdYTYkxfMnQTmTvj1H
5820K40H0cqnJ/aKC3e9wI3cglSL4fIrI9mfEJbYyv2dDcbJzpqIdvpyIZlTx10xa2ZcAWswLeSH
B76LLLMUEU47fqPDP8sHQHZvD3gZ+pKA+7VHgK28aAadbaGVSo7HTLy6h9TLZOh45HbzqI71Ichz
aoNgtQte5dWZG5G2znt/ozIIY3dBVx3KKZHZy5UMxw+YOJajThXD6g+P8yB6eJM9g0NxiK4IejcI
wrQln6uhVr8aYLrIUJuPptcnB37mnM7H9tOMte8LWqb6FPI2kAXKtM8yKH76LxL+jGtpxGKhrjKg
NMWylUvLlsC4/hQ2pSZrNaWhhD0N1ObEBujppZy/qdMdHVlBWrX39T0WpvTeL2asVHl8HMwYO+wY
iqw3rBgaog22mH33fQniq3R6QnZZGkgABvHnbsR7MRJqScuyjPSYNm+ieABEVVrhgOWdJ91l64ly
jIEh/hEdcVreNzTbPgVhFw3uSxmUc97+5oBjEaizbtKgvHXMqV6Lo6wTemNeMIIu0DZKmy5uvFt8
ABZkxCJGsXrHPYHJbZ+WToWj45/1N0zknV4+OU5zYK9Q9Pt3wzz3DA6XYwKs+crdLIAnApdptN2Q
VeyUXfuJpnQg1VFhG70Hg1JbOh9Szf+WVE3ADiuXK3HhEMbnLI4lV4keISLVDc/g4tn2rRDFUpl3
A7weABrGLOxV9W23QBtwmnx5tYC+rI/GF4+pIbMhwyyse8+I5W4aU0sfFjdiceAYsW7GI4xfI5B0
if0Uv9z6pWD8UsOVz31wkSi6XcgTrRG81gQARBbMauVPR0FVGR1D61a+c7m+NWoZhtC3J0RuB+ph
a/srXUquIDFhiza6Se2VMMOd/ObBVHKPZCFtrs6JcnTkBFoaCfe02psxymlEH1Pr4WU+WmzisD4l
Oz5Wbu7H8Q6/EHYMOPJ+Ln7gWvjyLWnagcmW5vqvIdQa9gAeXCLiSxokNiaiNjTYMNCuMU23NJbj
wjHkiB1r1GO9IuI9MQ8vSiNilFA/Z9fWXiBAhu/pVZFY07q+n5z9yeaA1L9f/gxeI2Y2g5pH4fBp
Umci3fFKbo7erV0zNHlZ4aKUjAWEGZWppo7rn2vLaw18tZUC7SodAIa1B6oJUYzRpKCK2aOJR77P
RJRCvxlHqaUecuCbm07xMsjgFPHtjwcTUwlwYZzqJkrtBAqpPfA4HKgq/5Kq4nmrDlps9Bz1EvH7
3t/X8hmL5hiIs9u2Hs2068pxsRIFCAZgrqm9bhhswrbF3RVllz0Hbw1M0cagM2sKv79zLd04iegU
KUmo4dDKlfUPo2zJHzWOc1rdgl5FSCm4EmSGm/eEQ41nN+SKOirdYioW0tML2+akGNWBE7GYumkQ
V5Mk9QQKvW3L0QbVL4d+2E2cVn2P7R6vYFnYr1g7XxNUuNR4AhPNBKdW8F8ZdsoguWlAiucTBaIP
3EC+6oBB19+5PW3XLoGXcE4a7gd1+zU0R2f406USg/XKmCVX/aVyCoHzKyjrbCfeMCPEcdZ0fu7D
ecZ2Ocd2fsZp71nx6f1iqdVz1M1dEzQ6wWJfSbj3DpdIA0qp11fGuW6Q3fbwZcl3//f+SU/6uYtl
4fmeybIMPP9QfStW9vuhOVHzUmsCUZNfXISZGOCAhe428LpjUphBP5tH8SXJf0Se3lqummg2+5AV
61txihVnmV9gEiG1hkNxhoT7OSN/atOr+zIYu1mMuMmw7UdXCCAREuWxRu0IZ7gYTma3qL7cWEBt
aAfXbyKRgtgPCF+n8IWkLoVYWarFH5oXzLW4wUlteMK22/TvAdxd7Zty9fSImPXgntafgR9qWEw+
U0FyGcMQxCS9xevgeW/PGuz1uj+AUXQHC2TA7l9Cixsa7hw9xhF7XIyjIfDuIOLoOuvQ2M3MR1so
WputEyLsA8W0GbazxsR4pQuVFOFqvAh2fRJf/2lF8g9vhTejMwHsgB3BUvC4aG9bCfY4DlyXj3GN
aJjl7vm14rD9zUHstUlqz7MltZA/6ns5wS4IaE0+AsH6k09y0El5gZE/S+LgpJRWZ3nV6KkoOVFq
MwgcBGtJIaMbJqjRu9IQrPlNvkmM4y9Op/nNtvr5dpx2QqYErGd5ZCZPcy3DdIfKjk5NoUYMzYYC
ARxZk25kRSAavqRc+KngPWoG1O/JLhfRpRpAtTxEvsjQ0FGOMgZDhpExv9gCLv0au5MEp9yUsgqm
1u5MH1zCp091O7IC9La5nSt/Tyj4MJPuaLz6DIruhS0LHyS+ZGDMw8h0U+EmYpsxaAMAjqVfUrMV
8ilBMvaov/bOklcBx61JAoZOVxwhT5qyujzHmr0XRM3aGNDeXQfMPdZMSWCF0dyNdl/lhuSoBn9Q
bxbBgT7cw5MpHoNDd/q3wo8mciakW6GUxuIvvEYOm9m+0lxSsihtg1QNqxTM/FitMtmbQE9MLiA/
yoOtqwkJugwfWiX7ReCbfAmpiBtba8+VmpPngoevCR88Cx3a2+Xf77hBdXsWXqjNnTqvYaBgnprM
s4IOEQbxSA7lNOAVpRB9Cc9NjZWK3cLHx2kF/PVO4+eLI1TgPnDZEP6MUhvlmOoyeSWUFL7xicwe
DQjmX22g0huHqTvCawtLR9IgebbzGZIsqCDBb0FMXTxMlxRXdy6ljMGkZa8mRZ6hyNES7Wf2ldGv
KvCy1Ljp7dT/POf30OHMWEkj6x9nGae3v0HYXGnPnx+UEA6twtOKVLqJQA+ikNnTbACMREMlvv8i
TJbjQnCxIb+qpRcuHtnX1KTQcGP2I2OIuf8asfEPT9PSyKj1Fb8R1tKJHvZqLsG07MbdE35Vzomp
Zt1/mJKTGp5e1+MAtMnGez3h2XKLA6Q3uIagdZ7Lql4SEaTh0zdb8QXp23vCZtLJXTeVds1DzJVE
ejDDrhTTV9ZvygQCH9OJM2FfS3Icx2WG7yA7asuG3JARD++jNkZ3mN2C+HxOP69g8UGnriy7nWXC
mjlvoGUPk+fy4TwSJPodCsHXaiFjFb4NwhpNSp81hC6GTIqBz9jsoq/bh6lPNesXu5V4O8nEQACS
Ye4Qk5HhSwlJNB+x2YsBMwxRYUnAYRd/I3KWaVBLxx3eMCyQEE7E/GTJSi3e0NttnS0FOvUM9IfF
DZ0qfq16yqUJI4zLEkADLKFSJrKz0dnIoFeQkImI50jh4WurICvVoarI2WHyFsk6y6iyG8Mz/z7/
riT7RO+eKZjt3JnTWQLLtxCa4G/IDoyAFf8U6QG61WBWGZl8C2Zm/TgnIdakVTDyx0MFS5Gjoj+/
Qu42JoUWFPHHAdSmGgE0Mth29eB5VAbfkaUzuetWnxZH6vWHAthn8MxJFFcMhFT1JaQR0uUkMGRw
k86YY14e+jQ8AGzgi6IzvsCq8IdWw2qmniAPELj/6g4/7/9U/ktCYOgzxHcTLnyqz8rZSHVXx4sB
+uzsFsGjZ3L9C84T6Hi2hm7stY2qhu09KRRX+k+7sAtrYQC2YMGsqEeSBcNgQDFFLo/6Ysw8r9+u
jraCrv/fXecDAQZ33ZbTqNLBhkq1zEwtyCBE3zhjMiKcylOJ5hmCw+/owXsJY0r7QTzTdjD38q2G
x4vuMHBBKLRLQPvFkGd0CoaB9V67rHftfvIMGLeWe2EmmJ3AKbEuU1OyJxievRagsb+bCxNyH1fS
Iyng8XfqpJER+WIGmH9Iwgv22zntAUGxTunxMxClVyf50MaO3mU4giWtnHvf3vfgQZc05NwH4bGF
atLelGFe5D6Whj5oPUNJZNsS0LwdUxP6etDUy9nowYE67YrntXH4xdUoLgSsbRAJpXaL7WbP2JLA
Gsdut+9bA1txRaymi38HOy0AmxBI8t/hgW54lZ/4VX6sdQW7TMiLzritS3LLSwjkmvHOlYoRnPW0
2//6GPoQK9ALCaiRZWGortHu4QoDVhONM91LoZMffgyfq6wEAlWWD5OL3yW0PTOuauyuo9KCYabE
FNiXd0CMN4cvoq3tdqz0a8o+AjYD9gSFCVH3+w0jvN8QfAYOEy4qSQMGGtlvK3O8GyxAD2YrVbr6
z+MXB/u6/PN/F6bwMKMNaeMjVsOqE3bL1i1yHLM2Ugr1XiKpRIH48lU80L06qWoEdHXB1Q4Tno5v
/WQo5MJ2cLYvFcP+oszC/9BpLpj6qH2z/ntpoc9tm6hAIQzLNYTVreNHcXtUlyXux/fr4LcrBBmz
1R5CGTOstCYKp7wTjiMviiTkHY5z6U8Hp7mxSYzuMuq4bAGVxAmWj/MhNkasuPEfRrXEA76KPH1c
h4/9H+snWe/6hlwmizN7474i03z9L8P5mrl5djJ22Pj/MiYlMtDFtFodC/mHqoJ+omaJphjbqgZx
Kk6+xKgCbDHUAPvRlqv+M6WlUbDWexIR9q9ArvMU6yqi2Alf2Rlf6qXECGlIB2RpySLTPinj/EE5
5FZkqg2hAhK9RpjLa6/M1496SAxgCVYkorJ7aGgCVxcu3oYpLd0alzg4++GJGcQ6zMHgTLa0HR8I
GVGIch87Ej75MIxmTtTQay46QbklskCvSlDuxV7ggAPPysxFTnqpxRgC8MRZKHO7DzQaeiVvuYrG
+xADtPHx2Vv+bkXDq/cCXoV18e4N/I0Zts2QeXyQBxUaUkYXA+M/VMxxKqT6d1CNBtjHjLuPB32N
N5/ZGQ/AmyBm5mbsM2GWu4Vj82fY8L7kF1JLXDZ0q6HiFbBdHU7jQs88XhtRqDs//t4w9gOWR5bI
GjenfiJsefPPunhdtQYjciP6pp68NjoY9cNNGvCVIOwRdGf37rS1zzesuFk1UZ4iaCYkkbH71X9T
mOY6iQzOtS+l6FdGt0kuHltaq1H5vNnrLGHdxIMcMJMGi/lyAotqOvBrqMHpGWqkNajPnYDla5C8
H64MyGLG3JfOQ7phE9Lzz++nG7eZ8y7s6aay9nUxXCYOnEi7znfxF1yU0bNeWpLZsla9eUGUsmsm
MtEclp3la1lN5uJdhHkxzBDiIqcUADTc0TRqBEflKyu4zN4gf9WbARbBbqR7Arqd3PXdS9toheJ9
AWxzZ0vwyZOsltah/XCVeHr1Y6yfZxlEjuhZiSyFpzt9MfHIz/iiNbsiEOZp/Sc0gLEveR1N1CHj
0SNDs1jEeATb0BgyBwtsSXN925nus+eOLujiTKZ3i21pW+RIgJRJBq3LZyx2a8ycVif9/bt4vYVi
R3raA0+bWZHLV32AWwvOsYVwJy8DPrwpla88vhUTq+goIuBi7TYbrMRoo2A/age+64qanzm6futx
hg9WZsiK92le2eU2F20NTq79MwTizLwmIcGsTrEziIOXpdiqYSXw/wmpqANgU4i0SfyNVKHuhj0G
txRoLwROL4TBo9elrgMEzO476IgErOwtc58WDbiZNiV8j7XR11YiueYntkGOYOHVbo78MZuLqfJ+
binSHWOspKzrIiyF9s1YeFoQHmCGe8pMWrcz7yFea7KXRx+kX8OaKm0eKIRih8u+KbNkwIe5jS4C
I3saSZC06WC9eTJEt5tYqF9GmApHiromKOJDb4wQlnvEDDUJ4vBiJt8ZS8BBu4Bt5m4w9zG0oQZ2
7io0NPY60f4m/3EB3ruaNXITZwOD2o7mLXMCuRRCndSK+eSaeWBjdtTMCHxWF6u/Yp71Hdc2Z42a
i0bjuXSTmGPm/Gk23iQE3DeoaPFQo8M6rvhhwCGz6SouiV0IecqXCPy67fbAWsWuGwxLQoXRRNUi
7mPN2I3Yb0jfBTHkvMgNJ8ZWWfVhbIqg14z6c/rS5W/PO1tCRbqvogcUUZlIjGo7RMsO7zyLLbCu
U6XUYZ7csXz1HKJRsxwWI29gIQKrVg/lXuybhQzlzqQqE9U1zLIKG+nCuUyejDCHCBNCkqGBxa8m
71WPToLYWgRGH78bWc8noGLxr5h8q6+kE2Wgouo87kaDqBpsIUFEP1ZC/e74gGQKHDoUhAo8z3QX
U+VF/AieNSud0AMkSTfB+fGdZKxflCu3zgg7eYLaU+ZNKkZwwrhEvvBfX3O+wzFZyx9z7O5BMRTf
lINaX7KNxf6p1Mfeks7PpyvKMFLMTv8GZNHW5/Cim35eOlSHIozY62JNESTy0YvJSEuZ/kxMhdZ+
xtvzDwZC/OtnOvhuNMteTFcWx3zltccrTSY3aSDWaIE2pi+SV53+bMD0PuE2jyITFdv1Y6pxCCj9
oK5xOdRJJQnEakOHfjqJZYRzGmgIHJvjze0s0cjjWg3XQ5pkFqkofLDtJydenVDb4TV764aur8g0
nAaYQiyxcgLa3C0bvkXV46SYVH6JHQG7bWl5yyDE2pKpPGPZGdSiHjJrbpcKIGDpj+pgn1rDvcFw
UWCynzVccYV5gI0sLCaKPR2m0+zMOgWS4DVOkKeaJm13tmTHT0oFJpUmjjGnRPXHUFCXgnSfB6ZH
KmsZfKZI8Ys+MPZw8p7l5DtOUJrbiasIQZJ4PQIx5fD7Bci74W8dQbSJAIfgXKa9NRk8d3IIrsKB
XYGeaEing+ZYlv9+AVfxz+QEQh0slxFtyI8P8pCOgCoe7ccrIb3UD3jaOPoMVgLv+JX4IHm83ofL
9fQ+LpdtT3fGSMc7AWHVfgUvnZKMjOjPCaBnbhzaT47cpwBACbvQbpe3Kv6osR35keYJoqvPnGri
7vxoazSCF/IR7IMUQgh9+P2UltYGn0CCPn30kQHBTyfyvayAY7wB/zObh7h4usYu7h+W3fAqmHbO
f8NJ+WmMQvqcgYlsoMgwZvd0Ao8x6P8hoYtj5hA9PhNu2/Mme2wsyNXV4j3TWnxTK605EIwGsVma
uCUKMDH6zqQhfjz6u2u8ZI+kWptKs4ncJGxqKb0vA9YZkj02d071s2RSHnsqW/wVavGGRgAwg/f9
CS/BlPBg/auhj2NlA7zdlL8aeBXWPzKay1EI6xej+iLCybmTmodTNUQ/kuyxAcU0sWEdUgFg0woD
jjC720qYemFtxaw7pDo3bvnBCxAjgm51yO9UYpEAKbOC4DtHYdO06IAF7+1EZvSIJwX+zJ13fNml
Fz4SN+IpL//BYgDo1ElyRoHyOm6pPaiRQJ+zDRs1nRS2pQgmh/q2JNTPYcCyiQEdYyN8cKlvOuqZ
I+sBoZmrCiz8RNf4QJFrWFetmEO+JuOOSnR45ZxtvSOyYl59tvT/ybM+ghcTazF4VKjAdex4rDgM
JyKiacE7oFQfBySJKeWqpmne43SNHrT2mpPB5raDAfJAblRHm1QD+pajpsOllYg7qD/jDrMQ+WQm
pODU/jlblUCiGe9otYEdFKieIknlQjlQ7yXlt5ZOBQowDevtDFceVLVAUO9SNRl3+Y5e6tmI4HuS
cVWhDHwPuM4CgZegeOJY56hDHTCcUXLafbMma3KiCjMG4wxuZFIykG/UiRpuwaiwsHldaRQnuDrz
rpseD856Q1SmU789f1jbNgSncpd551lCkiEwC7xFlpzwhWcJnHxHQZByELHO48LqtVfrr/aj6x71
PnmAGoV4c/QWESO13xKir6ilWfJN0mBxdD+rfrnZqNWk+ZpVrNKiad4hIMkbwhqMko3bEfe2IC+C
ek9IVewrgRTcBKbEgwy9NOMyBq5g3fJREx+CqeviAw9pFk0X3VFd9kqLsEjP7Qgi2O2IpCy2CjZt
0s6ytZroYJpcxZqRsgFSY5e49aGub1pbapyErMDYGqGJA6GpNk4yJ7re4tbIapABoejGuLj//DxJ
fpsWAvhvREt6OlgwSTzFGfAoo0cncvs5WYmqj/PgMrzVT6vHLw6RDnCmIcGI1hrHn/dxqEG8cb7o
kKeLEa4YihWb6qh3WQPB9OhT4iovTsPqJWUokGNRFVW1iQmQ8rk5VLpBQdrBWp4z5+HVMTnbHyYz
l2pCiji1c95//EwroHXTN7yxukb4YG9yVqPbU5agGA+5p/YzT6piBC3It4Kev/YU8wkYXZa7BC6q
C4oZ5VBGvNjkpR0fKT3Nv0uk40ypFTOsDcXmRnq6+L1pCxZxJE0aKlIGVFoyztMZRj74oumsJXOx
wYiXLVGUQGGblfr3FiIyjwmEfKFXDndNpP8SXtdeRkIIclQMEN6JWGZ0J2uJsmyua2w4VKlO3I+C
1AUJBVvt9E1Q5v2KM/odIrx3VU23tAZX+BeSl7eLyHACeK0cuJ26PhG1u8joYJG0BZnS6g9hACoh
2hVlkTkhDPSp7GoGdypWlQU2+qhvJyGK88aK7PjwsAhLQnp2eLg/m+e0mvGZOXaxfw+6WR2lfOzn
G1UC7i3Svy41AUT/LNUGf5TwZ7i5cK4ANEdO1B1KIRdRkiRgycU6mXFdZa8p30iEGZIpEHI8aGdl
3T8zh40fxx4oAaDp3CmESH9eFcN4DPiPNJdCfPemfbvXPc5lJnHmxO2BQy9mnM0ja+UCVnX173Av
XjLcUmNTO/qwbbRKOH4NfJloWD5v16DgvnJAjrbjYGHWXeW6L0KUiLsF4CiZH2VMKK6vuWw+gGxP
pQfHfnN7BEcOQhuhvxaeRSAgb8nfUTtH/aCf9SP7gIsJhwXKqkSJXbBLbdI4QmL0tZX+kUER8lRt
s55nx1SnhYWiX2r7a8nMd4ZAcp0b35t0+oXQCtqXfNNgQCDEuNNfieXfJRbbevgj1FLa1h5PrIvA
J9XhCrMJGBjrOCaG8TiZmuv8+FIsVr31XU6Rfd3jIlE0APz1/nEFE6qgHtXzxavyELfm7DN/3ADl
iUPc/B/AFy55K6lqXzIOIXFAHL06DXSoIuWDLZpNCIQ8JD7x/Z3pAinfWWhTandhAe19qtV8plG+
9+YKuVNo3IF1RpNZyY3a/Cf5psCj/HtRIm0gquR/oE1HFhXuy9j8mAKa2HW9yL3HTrYw/64fubgy
0r+QXJwjn3Agllxt5Z2b96+0a55lo4QpKww+xlPEMoiIRE5ZVtHksxcdrdLkr7Pp/gx/8lbMBGbd
zCm+zIvpDmRqELcDdZtiGQxNHaX7JnQ0Ab8c55t6bbbGqRGzIF+49BD1OAyXrzQqnevgkjkGwRzq
y+syIp0Z16z6uf0x4b6JHnvIe41M91wneITRg7EVCAByz9/ptDE4KYNmpzkYKvoLbe/Eoy+rkfL4
EvgNPG2OioJZu0aCJB5p+pMOKQG5XrWWD9HD/fmCNCXYwJJ0RHMMtrfstGkm5UDm+kARqXl6kGM4
T0frpPspF7fS3eCPdsRy3AJWu1SMmaJPn81BcUMSWPDYDMcgF4bNlvDblHF1Oa+FQgjSDGDAV21G
O1adA9e+qAIt0rggZCbGkF+xGFtHlZ6cvuJrb1ZqAMRsYymLEexVwmUiwyzHjqwRpuaaVhcjC0bW
uUflT8F/mzwrY9RMcyrG+BjUGGv1/iq9CZ1KwBfJsMn+qho84/saARSlsAUrO4WrglgfV+yDIQKv
A1mwiEviKwaV7W3NOhHJ+A8Zv2oSjqphIDFFsC90Ta52It3AcszL5nfQdltCJ3P5PHxaC3oLPEpe
RLtHEuzG7gptTCISU82+7+ccLcVBjDFFnMSvUANDkAmzo58iNNojOKfuVMmDNKzsdQ877A0olAlN
NUIox78PRdDouBo0dE9QFBmeasdKsNTnerHBcwDEv11/YIAc8eKLcPwEzZP8YMEtZ7XEMjQFQjqn
wKkNw3wTef171MeFLViC/JJfkr8M4ekLDJY4wW4nRd9FzQ/K0CrZyewYCMeh1OwJhmAX4Hw4vinm
kr4jmu0LzdPlel3oF20GQJpRcwpqCNgStbkxw9/F0S4TSEmIxpExwAnUhVD+3iTwbifvxZrk1azu
cTLFy7dcA/tmDl3oyGMbocf6QABYpcdHm/aKYBLmQlYGyPJ2iLlx0fSOGIfuyzrNscxc4F+6axFT
ex1/7kV3RsYqE6GLX1ZucMOysDOszPVb9Solh6L4wKP7gPmkNnhsCkk/5He4Uv+8vlFMaYP5whTP
GM1Y/NtOrliSNxh/BaqbcBeVe/Xh6I7lwGSJnkUSstJU/djtnDClHtIUlFdyD7mHH6PPt6KUmp7W
z9h9YpGufmMF7LqlzSZcSim/FiqnOOTcpl4s3k4D6TauhJeBw5NdzkW19HXx/TYmasYR8i4U7+1m
uhdpdwutcFsb7urKpEg438gDe5FRQRzqoPswRMNPZc5Fs5li0LY4VP1JiWkMwRk3iVpIvAKa7jXY
syIqofrOk+iLWCa7gLDTS/MIPFiuxsGOgNQVwjD2UiOIoy7bUotupf1Q39qq1xfcbXze1MNCo74w
dCNA9FxNfqnlcoZHcCHvN15HPD1TA/Fqw6EPbwKLBf4tiSIsjY/wle+7WfHGXWJG8b4Zz9gAMBdg
F5qsTnIZIacPXYi02OcnJvq5s8tGsyESFGsXR85UHZQSPK8IgK2FW7EeJ6ykNM6slb2hvNbtAj5p
R19tdOSxlgDQTvcy08iayFDLav+RqrTGADS8HX9W2EqkbPz2CVNtQE7RlUQxqv8840aXMIkpXT7t
QBslNrjt3vyqL8+GXreZc16wagbwyniNSJIfluP/RBPEQp5fbuPC43ZHZmRv08wnMb+u3iaR2mdH
KmLE/znadBlufTSFkWqItzNN9EUss+SftQ3I9BqSHumgb5jcKrujC3iSSWwWrK5+mGBUNOU1b2Ur
Ugyod2p78tB5kYOTQaZSe5F6+eYRGndgoYMsUB86n4yRoCjgi1KN5yIiiri37p334S78lOadxDeX
LZaU+TK6JDt8tec8IM5YkyNEvoRy8koN59mTpk7UQRnidzfs1q+tM+re3aLbTpIxtcql/mh8TAVn
pCb6R7hnc7F00GUrx0eVgoddK+nn5mN1Bw4dCrvuAfN4xNdmVXbd2zCgt6URQM3r7PwpQ87Adg+w
A8o7Ib4f0SUuINCKo7KkksWnaIT4GIhRCMukTNn4SQFiH/9pyNmr/TQCgV1dbzFpSVw7Ap2sIuoS
q0VfLgVlQr4xYUCTkJJ3UuSbxfEqRLPBWMgNzoyDY4onn5kDaLeysz/j6gtKpN+see74sS8CRy7Z
PJQ1O43ujJ3wrzLCtCs0PdMGw+aWYo1nA7c7SaMnS8/1eY/AAkQ3kMWWTO2KnRN0oZesTNhboi3f
MKkMeXp+YM1T3UmL6iPjnGlQ1fKodywR5F52GTlI1iqIM485D7c+QVb7t9gBSmZK4lBWH1Y9Ow0c
+vqDcJkC2IVwMxUndxSUvsKNS7MYOVZmyd3ve95AFYaSKyCibaj/ceIUWx0S5Vu0eCOlxKSW9Q5r
PamBzHf6pTJ/b7s60himxUlt7/BnxCy/dq6d3TS9sDrgVONiF0wH0MOIS/485VurrDH9YV4nnSXh
Chz0uKTgcl0RiUKbyo/0qVsU9TgwfQoWElk9QTbeKCwGGtD3TcmOgFEgwz+9oeXtJuXv4+PdQxP9
ixiMcn1ss+r84VSFCX97s79MzD4LYdfzNi+6IucSYj+H7aWcJ8FBlN1qRmVMY4U2dB6aDAUVMxr+
iO3EGp6REuMNnA8tjlxGvwt6P0N8sk2x+rLzeNtWMUYrnokZw68Ow0kfeJoYXhR+AfS6iZhnV7j5
f7JlkSx0Hdg5V0HxS5evjI+YxpDARYcLgmaurqkCIMICYbYxJmAbmmFeIS5EyBzvojQKu0L4619z
P2FLaAbxTurCyqyY6D/qkj/gJSy1xmAcVwVJv1p3aPMwuSZ/8kLLE1yy/eDjD4qCLEWa1nmEZzEo
DNq2LjdFBMPJAXPlGY33JwO3ID7rzu5Agr2iymZ6oYsZfKujKYZ46nvFeu86WCb2629GCREyRM0m
zY5ZMRNTvqNV3CKambUhU5BI5AgmMzQajsZxi6M/xpTPg/RoWot5AlJPqoC2BZsrw1PmLLYoCo0O
6/4NM/pT3Qpke3HHhT1DOjZvT8UKsHVb2mHIl5KdJ5OH8XaDx8DuncKsYFmx9s3Cp57Zm4cXnx17
IK5hQNwRvTmpVIe1TV5pIZ0onr96b0QH48ODUEm+HE6REpeFimzy0rAwqCCBr8YKgJE1FivDduWo
45986/YfKqx+z1xsK3wcG80xukYxqm3igUKkpZhw1XfKZ9QXRTo0gMG1DF6J2M6FWOCOL0pHM/Du
KqRrBTCPjlmxTJg1GDNCZsFs+Gp3noCvFkJRpVhTh+tDG9sLgUkRdAKzBNHGcW15qSy3frqmzx64
0bR+/EMqrJvINnGKtMQ/15PGL3uBrjoNeiB8zlddQVXrir3z4p9goulpwUE3ob/31LStcK16pMEu
+p7jJmvFCVPopyjh/8IUW2WjtZikLeY4UYAcqMNCWD92/p1Kr4qMwTYtMolzP9KyK9hZt/0XfW2W
Q2/1qJdG54bBgHeZkRmqBijp86AwQYDQl2kHe2w8ULgD50CyIAtEDo89Qo94kbNJRpskGO7OWah8
3Rll7J7J1CJNaWp23qSYh/KfQg5jrbUab2hXW23VGcpxKhQ9S84urke1vdXWzBpcxxJgEpJYY95j
msUplfVKuFxH1SZtAou5qLcwiJnGxxCxnk1auQBtPxY90kNWkFwJlNTOgtQP830TlrnPr2jjUYxS
AaDeWM95bF3FN2EleckX1ibVLu5bw2CJ+s3xhF2PIfbTcXoWGeWskMWo14zoT5qq/Ncq3sOHVTS9
OecG4qg2U7xY+wswnXzVOmBrsyrLKAUgoQEsb1bDfDzdpv3kEgOvrn3Rr7WFw8wIreVIdam2J7e0
wlZCBioUbt04udPotJSFs2imiTHaYZV1ZwKU0e3BwVtndiqjJXKsB1vzmFJDJa0N5i/pGKdSabPC
ElbSMY29wYwb8syUqzuEAEMZXsE+J1DV6zVBOp2L9nkvc5h/2OnkjFa5T4KW4E5dx9nUu7cn6xEv
o2aTjbQn9VVgTxKUhsgXItdD4ac2azuzSF54Tar0SQg0HT2F3btkvc3U6gpoYuNInu+AWVfzE9UW
Rq6unr+pTcnnIn7gs8fK2PwiKdKPH0DSiGnMJGUpzeHdMp8WYIL41ZKsSjqyGygUI9wLFnVOsz5L
xm5ovkx8psPpP00Miph6WAM8Pjhn6EfTGnqpCKW5c4AWtlkd9FkV7Ws/QL5oKcnR6fOiMocw2YkN
ljMZMzjEdHMrVaL10mBlXWuF1Ifr1lrWDKqciQyaJdp/Wd4UZYfDyjQ0EUZhKzPHErPkXgTU1si/
lWoMor0HbE/2nhjVzhlW89EuGOV2W1xEu1eu2Id9cNxOgP1px4L4ahLSVdvUVyxPbLTd0hts0clF
PVDTyuAxYvCLxL3zMi10AEBMMrhGrEDcyK3HR18NSFBpR09lWPXP4DHf1poYFyQzNYa9oMLmlta/
vIDOHYr7zGFbG8kc503QzNqDxMC2FJbuS5rYKipxipcR6LsrT0DQvVwCGcqvKEqpt++CkscTrSuv
Oq1A2ZmVD+v8s7uWh4zkbsLdP8FUNaS/B6KAJ0h/nTNnM+qfszr2pf4m7pO9AYREhHQqklCTYc/P
H0ME+7w5h/5JZmVsJ11jI0Ft4qM61AnL7MxiXQF1Vgoi4y0HGPrt7FoLjf6Cm5b6qIYzp5qxGKR1
6Ozn9CzTYjBfRxXu7K/Q888IYw9BVTGORijSFq6ZGF5Ck03ugNc/V6uQATAYGfJJZbCnYUE1L7CU
4hGTfU4QBPkJ0Pq6g4bGHS0kqsgp0oyKfLzhACVrr8gDV6lbx1oZtmSQZi8brYs3bsfbje1sCha7
L2+C2iTkey7Uo7ryTPN5CG07rSjQvmqkQOd8bfzng0qYXOmKiW9FWlY526pvKi0ggUDVbgeOrD3z
2v6m6wQWOdubp/tD4ApyvHQs5G5oAwBVkyNmteYV8FRzisfj1HOoTilTPgsG18h51/lNZ4vNZEr/
YEYLbtScERyPoRhTnn9Bqo36BS485FIzw9i2ZKwUy+HA4Objf0T0PWVSrA2LTT16puarsFn8N++O
5MwC9zfqqE5gBOdB4MU4flzx/lZS7t0+V9WqBGkT4MXUgVoqunxzjqYO64bMdpT9ry7DVRwa0VvR
ysBlvbIELszPVX1/RIkDzWRkSjPMQO8TYg54GBs89/yPtVKkWWvO4Eh0fdFp07KkQgL6pzXIf2uQ
Mtf4jLqdmtCv4k+BxYxHszg+cQGVlZpRwq4pI9MKg2tWVAhHoO2FlUNVXm3bKAUs86gLb6pjKwij
HL6n69Z9NEw5/rAGdPDwMCu0DN0xUFWQj8mDHC0qkHlCvMh9Hbfxjx1BmhECBRwsK+ltD6DchcvR
6f7WNVSVD9Y0JZSyQfC+yEdZDnK/Z8mQv0sQPYnjHOClBkt4tAk+3mAAbn+6ggzPRNbWjobbjfS+
OkdokN+flN9X9r0AwsUTFoqE4R2G4XvW+cZUw07X+PDNecgkjSEVho1X9O0EzzmelMiN4qoFI34W
CPbrou7NVBgMrW6NpYqML6kERjQA5pbFlzmlDH1JD9OUrs2dFgZOtRJaJyfnEzDoLph+9sBr2A99
pi/VDUs4B7/2r2iOczPZBErBaePxRzmPBxHAuWjjxivGzygUCfgOhEJjq+n/C/fBoVtThBKQq9KE
S+E9ZK65/Ygz4LEtteeKg+7i/EkWJsV/f70j7h9YPp0x8MyZkVKu/GfjF3zYu/LzotXACdDfwnaA
BjCZucF78Z2sRpfBsdkUkkatu3WY5bftdKy/hdQZ7qqzyfamkzyRXoLOKWyTwXlraMFoMWySCV3I
UPhC7/BNrbeavHp7OZx2wk0epnr5ThY4FscLHW+8C6XOpWuoVyF7OQ0b5y77+HM5WfJBckaHZGX1
8jlATVO0ekhXmvhlCeybRKXG42l+dIT1mOMhsvYObtJ01IlALmUSf1JJq0zHzig2iLyHn019ewd4
xqIB6U9H8wd6cTLxwLdtlbOM0ToW2f1o0csgOZMb7ptvKWWGwnYhQEVX17vt9WpzTbgdqYmw2cNU
X3XP+gRSZy65IxR5sG7fpWLQUppQGX/TwVRXpL4CeAntPUOaOGjqVH3Qh7UkjaA3yE1KWmnLPX13
AxW4cA8Lpl4aSU+8gckiyHXOB4xNM0Dte5/iDNu4PrdS+qD0lUEdxq7lRhv2YF69WwJOxb+wu21N
OWrQVE9fuwMcLrc6QLmXfBkqjxqwPLt+p4EOayu2akPXWNfQL0kuhoMB8crav4NlX/FfTGMuDTCe
Nw63gVuXP4lwWzJkhlgTElLp3hxk25cLFA0IRLX+EBrQov+UrF60DzLCciTudojLQPeqBNwf/QmX
nMG8UXIjlH/0+X5jhbNtJDzX4cwxeNqxGk2/OuedHTwMdeAYgD+skZ0VVY86BK5g7QPXncD5S5Wa
cjGwV9n62JVq+T0dpUxeLPrU7cbQ6dHyn4xwhedWvgGTyh3mbuQZRJNX1K/wO3KVvypDi+iGdG6o
TG2/UbDwb4eWaO0NoGgwydU0PQBZl11Z9FI8Qw3V1hmuugR7KdC1cAUgHyxJmq1sL6zZ4hmD/l+f
oP34IjqLHiPdVhNEM/73Efd32u0T2kC2hDeyo9ruZ5b3UgVRTMOQen/fK1X7oZA4Si8WqawdlP34
bSCTqGgp11394kag7kNbrow1Rf59XscGrA5yrPyZumnmOMNq422xfKSuWmn33FFNT84oJ08oi8VA
2ipYADONafIyHfyNM0xBiCGdOhu3b4QDEBbhmwxkfTiCiCUe/10sDalP+ZMHQu3nuZKBWdQQp+/i
RFdVstf7Ti6mss1fcaUDN+etoFnKPbkRRpHyfahVzovGmTj0bKee+7oHGh9j47Hd64RNBDkwBy+K
R1Yg6iX6zTC/1ZQg3Sae3/ulgt3cL4Ob+AUuzZY86GuQl32Y0fCAlGb9R9R1EZNMaR7Y7ZQnsP2g
2GKKUSo6jgmmvChcO1hCeBQFGws8H0ANdunzZeq0JbSQe9bpFFdRBWNWW8H+gD+uqNKcAPxTd9OV
Io10sSxgsiVkeO9OYnDQgn8fzbIJWzmiq1a2POhQPB/GdrDH86rNn87Mxl//b4mr10AO4r3Tuz3H
2Ie38lQZuklElyp6O95uGYPvWX08jgZcSr5uSRM1qtc8r9Q+9+mYO6fzW0o/ZeqB3HeThC++50aZ
Xe0W5N26g8RV7bS1brbobjXzwdIhGwIcSfZxymbuKQiFHsNoxDjPXwoHf7L3mPSBH2hXxiixOZVo
Sz1wmGccOMF50QX3AnnFIw6EBEU17MOY5mQO05ZZk6mlMYNZuJ9NGY5G7nj4XZHbxq4BDeeQpJJw
2D+t8njj4ggNTHBdUrx5Yzeeb2X/c0Chn4v6kOgYb8wpo+GxpfVJz7ExI/N0vea0YJjKeLaT45AC
C3Un6NNrjc5PyURzHh74jc1KOrZ9H27z+tP8vv6qxuSIuKNEZRVXrm6nEu3m9Awce/WFZx9i+/Lq
WfobMMZuqWAIVu2MaOQouPsFzUVNKVNiItt010w/hxsWpmjKtPs2ACmMRpNXWGDdtHYpjNJfuRpz
bis+dbAkgcIkVOp04H7hz8/1ahdwOFA/GezylKt7qfzyYgGZolDBzL6uxDb7oH6n4zHnfKj26g1C
AMDGNhFoOt3wAkKkZlkrUDYh7hzmG1R1VbJ7ePzlX77UIfF1l6DvM6M4pjz0SyUlBauXJxrMdbGu
LYZtqttGe62HMJMLeiIP7BXqmPyVpGmQfvfep7wD+ndLFKetB8Z5pX6ipz1xGnG8VuDmfUCGBaqU
2QBEgAnvXZAdYV4GIxRYkb/svnmugl/arXVUXrm7s4MrHim5zP/AcB5JXyrKAQRHa/ncMcjqMsu4
DAQMPK5IrRA55y2N6IDrA+fC9ig8n99TIn+fMPTGVG2IvWtwagXZOODzRkjoNUmKUYFy8YBOHJjh
BuJrR9fFcE7LKzno1Rqwnsi2xkaOa9Ic49Cb4hZz5Zr2X+1qs5Mqx3lOzx4BURQixKV3btQj8qis
qR1/M3jfiYovHd9GV2g3X3nBFdWakahZ9u/cltZivrQaYeuKjkhFH/yuCFUS+B8GqyjMr3xBSceJ
j6CHB7AwEHF5cPwrpbHc3+5PfubagypQgb5Edel2znoRHxnBG0XDIePMzWgGZ65plJrijs0u+rjc
9g63FxhfTuswjPX6KnJ8VueX54Ti5Yiwx5gH/+ncDrZR9E++2qI/iT4RacMwI9p3np0ILaWJ3Egc
/TBoWdHbmtnsimH98345WB96ZsmtVc//ldwF66yvY8tUkxqL3FLfLl2KrL0QTVf4QFzPlKhQWZek
kZrQUmZtXKZyrr4WP0zzR9nWp65g61YAAYfUK0h6sE4jFbQIlpk9MuJZhafDeQJepVSfRKrsa2wi
Cub0qpdpbkzjFgtjkStWTQa8LU2fX1gcUFsDVh9NvdLNnFkRAG+OqB0ouNZLfevEbQFekcHZQvep
jP6tKEZId+fgrRfeStVLHu900nI9o8G3rOJBSWefUO4+z31JWJfengBbfXwiAO4phWNIKoVFtasx
FsA4905JCAD0aRinBWSA8w7uwoDXhhypw2DpsSVYWXwzac0QqkGrvLgBw6pzM8zeWo/KHwHznGD+
agY8riyPThiFDPEuDXrzR/b90pzqzLSkl6kmbTX/xde2rHAxm28gh1FE496F1Mxz6P1yGyiUjcrr
/Pd8hI/TylFrhTpr+oHJPiDPQ/IETsCNzg0HrqidpP86f5ma+zzUquyGe6pAVcibE0W1w5X4Kx94
Wy/E9xIYMX25GKMCabTTkeguaLJT7c4VV+VqokaCTyrMt3xzN8MyAIZOawXCC/dTtlC+BGKNO+Fw
+jn+iBfgs578Flw555WgIRtHWUB3so3UDXxF5LXE94wAs78Kel2M15BVnoUlITwsljDg+3GMmOwQ
GvIgSk4V81b961A1ddRdSdVOJ64j04e6X+vjqpsihoz0Tm5DqQBMQBmqDBo3id7/vwU80xg+p4YA
SD+a3U2lH0VALnpUCrflZeD7rZlfzH2JlBtP/6x1MLSHXGLfUFWwiZdbSy/6veEIY28tG6KqGOiJ
uc6PLv/K6Z6nggNZ82oVdLKCa9HMAXNJ5Li89uQu/3J7q8zw7vNBt0sHdMVPFzXWEuf5wvEnFQcC
PDpp0FmoBRt7GmVmLu0GHphgFfqjopRVBQoG6wAfgOt7GT2lJKGbNbR53UZ5kgdhZ9FXRFHktZiT
CslJNNrAM6aJ2QqXB1WqVbDph/fdRgV5kWriPhWD6FUZjQrDUCJFK0Wbju3j/MJ+BqW0iKeysTSs
nE1JoHqP5NwyPuiBCXEAfV/lBT1rZmy3JW73TUM3tL4LUznFAGah0pA1nQed6cI/+Nx894lrOoq6
KnKynm8vWomAnIuF419zRNqQO1BqtzsmYXa+wZ9bA8QRbsUQuTS9KQE+pBRCGq+IEqfZqDvFPZ/D
f7zfkH+IUuGIrVdxV/H0szk3ycyXhLWXw2bvWRrHTAmdzKz6RHk6zOHbI994JtqeSpVoA6nPMF2y
xNOn6bDHiFO40o2kNzv9DbAXeBRRl+1BhxocgaiZEolX+yZG9QJnN76VbR7RN9xTEI0MTTJPfawF
93tLl+JYmufJBoq66WNUQCW2dzT92yqugPtn1KLvHPSmlnbFnLzGjuAei8Yb95AEBkooxCHuepvu
fU2RWCowuFUL6c6qoFe/+xzZhZsXZN/wywGfHL8qdUGEjKznaoFlZlVgK89UMrgP2mPwYwCjd6O+
tXo6hGCOuJIqKrhfIrEq6lHCrJux2QEdgof4ckEXnqR54MjX2EYgsH92XfQN/rPZKPbmAz3I2TQr
shlkLnENc73WJwyHGfvUPoQr92KX9h8EXrHIuGiOdqbS4HWo++tAGbMEEpHLFosyiq2UVDooVE4r
wsu8SGEgM0YdgPbIX0P5hPXCp2FSkbU9fk3Yr2/fNgS0k5iG9EeDDyq+OR0roIrEDuCyYKG1trJW
fnDqOCBE/rMlfjFSnzJ8eT0eZwogziVwtvhsL+B46yq6g+3XULJ/7rQUw7FILX9SFzVbCuLCy3yG
WDuVchg3+wmwLEPJecgD7NN3oq+kByYY1+HJDaWifgUqqDW5KZTDXVmOpiYIOYgcd0gclemhfsZQ
7BB4XIMBSbppA/8tk1d9wLhlc5+50LF9xqg4slGqiRZFyHP/riAxOg2YzQv7MsKcsA1gB3FnLSOK
Rb+ZMVC8NNSR9Awi8sD+3q5L8nS5t1f7TR9HraR3UqXmL1UMtjTFZuA/a/6yUxclvaKrlxp1q5cI
qRW5tQdciY+2VG/d4guueJv5KPcSCkCe+fhAjrn69ryFonSgBx/aKk3XvtSWbA9a8OKkUlvEfHRB
Ppuh+Bhi3neh61xhZlKfOUV/R/Wt6rNZ6qIihzAEkEre73iJPX9QYYyy9c14kNyyhGjnbOnyu0G1
w4NlEYwIq8guNg+StlRkia4jLiFioc98w5M0tg/8P4UYQ0VSp67rL2/dbrIsmr1aEh3xCVyos+ow
rgPxCWc5xhYuLnhOL8E7nOail/RuvMJcsX+fMDlTZpyxGX/WIquPA1BjFKoiOe4uhE+6nMaQqXIc
sRq8gksHTBfvbbFb8S4KAc8qNWZk7JY13sSkuzU1lKOE+tKtz1zpg6M3pAg8kQiTzq38OfaFQ22Y
54XWz79FCAY9wIUcU9lN8tffOh0Ir2gQQqaEP9pDrQqYaajF0QWO0WLINtmb0VlqBOxx90oHmJcs
tHHf2VihdOBTcqyd4lvuedXZP0V2l3+U4fFjZntORZctrv6khdVJ5adZMk6uzNSf/gji+MSSHlZ8
pA5ue7acToQNnFRWzJN5KTym0PVGhXFOYx2ljUi+qJx7PeEyTnytsxXLsLnJFEkjGvA/+9eeaAr5
7Ee3g/qU5uuigSJJ/SbZzShexn0HejVBf1peorEPbd8svYKa5jGWYA2tXg7SmrNoinIS0JRZBqa6
x/Itjv25+6eQ8fyaqEAikYfpVcQa+N+Wt4oZjs80R/LqSxfpCU847OViSWWMfoalrFn4Wn766Hsu
GbA6iJpSVudWQBx+FCY9e/Azoo1t9JM//hqazHKZFdIOcuXH2t9HIO+IzQI2a9KgfC16gm9hQKaK
Zu83Poi+YKCB89LgPJHSzJmIGRT8Pl2Udy3/QVaT8hnnT4Hhup5SNmAEK7kdDycQ7BSex2dTBbCp
5v0TiE2Ot5y4wEStBw1qS80yIlgD0Dl1krgNMIkWmrA+eYHr2sgB1gtFZrGWlL91G1yDg/GY2rgi
E1YOX8DY4LUQCdwqmSGnMfix5rv4vvJdwRGa6VJg7EyPniMCNftLn5LupmlU6Ow3I4HNU0i+lwMw
k366CheEwR4kl17UzUxBiro7P3POjvm5U1ZIjlgfJlaFzKq8CPLpZmo4I2JzTtQHxCRWtCikGZ1l
e8ER5uPDqi0trOXROov5LkThvenTj416QAHPyrR7uq2mYDh58V2Ry6xDPHEUbY6xPS+8KGL676bu
p50IXgNk472XcGVfVPkDwSUuZ9RpagVP9bl9bO2swZUaSaDlWjYfd45MLgr1eut+gwjeSnduSM0Z
6qESvo9RasGtfm45KznrZtcu68Cb37Ogna1oNrNGIKPq5AkIVRPAvIlF1UKGyGTHkfTy9rHO1R5W
abaVm5G9YLyJclDzI2wDdIsjGfL+4FbFt1GnYhMLAG7zQMzxsFVYfEQzSkRlldLf6BlB6cjzJVYD
zJzWXfPta15PlAcMlzyLpLJ/DWnlKttWX823BSishUuR4D0pXVjedOeflZ0cP6ZpTYnm1R2nxwXn
+W/FeTmydftsKSlJ+6fG0M46jlXq/JV+yRfKPnWxIACfvGUDQgcqfQTsH9Crl8a0DwjKPMilZ9Rp
ySCs47IHeBgC1hdHdr6jTusTP3FldjMePe6/0yQye3AiK+cOcBfMxDMm2u5YGbMO3RrLQl5hKUOA
7gOmdXfLdIDlWkacJvgoJ18OiBDT4iRg8I9S13b3/1DCn7L8bJkW9f1lnMIpoOUDGLU5uvqm/tPd
D7N8GElsXjyeqdTeBbTkOqMq3ccy76HzYVbuwl2yLC9j/MUW0qeq4lphGnA8IErYOr+bALavODrC
IidyNLgpBIeJsOB0Ytb4CEpfkVIiy1J2nT12eVzyCUU6F0dekfpSERCcgjJPx/vt1fXnlwyh7rvL
lVninUpBQSzRqlKq7bTxS0Aj906Ydzm5NSRC7BDsjnNDlrns+EEoqJgb1Uq5Kk6J/ennXn6jMmu3
NbAyPwrfKGIfdjdqGwt/acPadLaYKkNrwGBSJhJRu1MqqBVqGwpEwIqwIv10dHv/2rboVC3HJSC4
1xyZ+ZzJTCN8ViLGoAaY5POxVun8bDMZEXGcBClCB9m6M+ARVDlpEJ6sI3mAZ28sJILdiPO7WTYv
LPqerH7ZZHwyFH9/Ip9yXPJQQBKu5ezgcaFrhE5XrTmgtJZI1B2LKCkOQtdBCyf+ayLrpIz1ATjw
0a3+oVs6F6BymI/rAhtUFnY2wYSDgbOv8sFB82ruMjSY11ZGHUrNAqM67DZxZ/u+/sq2/G5OnNVx
aQ4iJolO4DzRkS+pGQKc4dUvGy18a6v8pYu38aXl11gcTzy3YUqaQGtSOFBqGPyL3iFreG0hOti6
dzXbhIHHjxBKLtKiukaAHTC3b4GuW7QHmyCQsQ+syIqIjBS+a9m6mWsj93+6sR85uYp1jrccBVJE
zqvVwi230CLLrFc8vq5Rn8Ud3Mv3h7cxk9djTrbC8a1EQTGXECq0Wl4qhgysPs3EsG/u2LQZ5O4f
2lu1bvLy2HrH5Ytazk+VI0rs1ZO6h/W8sBRlOc0PpfUUMkGezn5IhqxxLgKBWIbQAdYCyx7xaF97
6QhJ9tXV9TZmTUeA54YlcI7399bty06pINDp9SfQiONJbIZuNU5R/nFvKRA4InAWYaI/PYcp6VRv
2Ur6/W7M8KyhkBRkZ0e1i8V/OlxXH/5lyca04BOrj7nt+O9zBSoCdFPL/UHugr5tS1yxNvIT49i7
m10HJCDvWaGxbIUmq8BG3gmbWSEr7raZeoCyoSIaKiovWqbZsRspYCC3xBNSpeRyHEwXl07LeuFn
AmHGEQSI5JcuJuK0yXTqNPkAjGjfqTFcmvF1IhmlMkqbH6JkA7ReDZbD3q5iM+ndPsiCTahM/V9W
c5JWprEet+0lcLutBQkk7CnoRL1SmwwCECJyTTqhUcGWH2rgw4CxAwQvPyQngtlQv9xdoqDfNX/9
fIKr+XKTN3PDU+JHfCgaF+ECUzXh0zlvayEnwFu5hhlDc8j4dTV+V5WawjsblYq3TmnejF2Fl14E
H3vIG4pd408enbw8mE8eRBtTG9gr7PpJ22+3HdCRW88/AYXW9H/5+cpCu3DFQ/59yzix5oiofyej
7o7c5Z2we/NbCJbbMUbFzxb9HZxMCUpzezkt3tzS/IY7Cobgjs4wWIc1LQ9qXcSVfREdadc4AaXU
tXrzOrDXEgnP9PXbv26uqtLl4TuXzIfH/Zc9sNZ5FaQ/+xqlzqo/si0uO30ZdLIdHm4YbmCmBjHh
9+fa1QCoEVbBrs6p3QudSIhVH7ElTScP0TmTTO1Eu0LlhyDhgYl8RkJZBu+cX5ghfx/XFvYTr+5u
RI6E7JSdpJQCmDA6DMUgz8e4CgJu0I5QYmCCKL0ceOaIV7TrxAfQAHkXXR4AGmQHRAdNzwKoNRhC
ZnQT2MRdvLiC8Xl48KHAjAV3xb7el/TRSF5yKNs6MlUjdq2fFBkFd7gdaqFTQgC6kn+TwGzxPuQV
G2aiTIbFtYzhX4Op7ZeNlCbVI8dvUwfHDzXTl5Ff+qRcfOZMJ/KraE2VxXUQ6rr36+hakebz6/ZE
44ZypkxInt8GmsuAALIvAROr4h7MPE8m9+BU5KVhEotkA9ey++n2ExqEB+zcat83Vg8U09/Y9T+W
dXAeK7geCsKTboF3ROlq+cGAmq4JgWlBUq2boBZwS5EakiyJNYd+dB3V8JRh48V6nlIxjUX/wMUR
bpxQ8JRm6Hs1aK3pD7SfaijLuMvWqdneFUvSnSUltUKizH+efugkqIqWbTVC2I9y9+HE+SxoUecK
gkE8iiLidRpo0Q6ii9sV4d528LB5IjZS3THlDV6rsjkvani8WBeREaFTYVeFOujIKw1AOvb7iLGZ
lCNEHZbd60+3HMnLVBg67RPMOHCAKuzC5QuR44p41FnCKdjIWdXBLQvVer5dc1DV1LYpKxnhTkBx
4joq2ibcOxhNC5Pp+GQ2wgcg/Pd0meRJsB8Wp3eV1ilQ7yE6lAFcjLK95gM1/6RMp0SGrXeUG4mL
hRtg2Z4aAA4yZrE7bWS4nFbBwilZHDZponREKWSxVnghKhVo65zu3NZmwMLtDeiFlFPHcsnftlmz
Idjq101C32YPNkaP7vaOBDsqHolvAJWW9b7ySzdSUv3hqeZ3oYVGUi/hbOMf5ZMfdv2cHAJuZCyV
9Hsnp49c+XrK/aT3p0UBYZrrRWsu6kEjJDhgPfY5Q+VA2ySvv3W+DvTNKWFtWbCZd8lh7o4AdaiV
fIbFOHb6hi9T9RnsLda3S0BJYtpS3z9q8hkwLjcVeJc0SfYEqHdn6RG4VPnER6IhTE6MvzNvRalC
qdOrKNQuIMCL08md/g0RGYBJfgbN3D7vo6kRrftkavyGbRI280jRpXpWbpTWnGtgIdkxzatTAYrG
iUg/cEnDC9A9eEaAy9qKr5bYwb8a2TFWnke6n0DY+sKchj1S7f12JsOiyyDUERU4ARnupW2Qkxsm
hB+921fVt+iynrVwSfCwevUmIpExVmvAYF0uTyYqTNf1J4BnMtpQ4nI3h0sKpoV99OaGFKvcCBsO
+KFt0n+IKsWVbws0pIX0suaYSqWmypju9MF8vqlZWuoUHqU3BQW9IkzTtrv7MLgye+rtJPkgkJnu
cEQtX5GczSzOg7DyuxvQ19j+zLGNPlaUPcPMn1xrL5YqWdeE0/KL21wBrtHZrkoYR+Qt82uHSX0O
/gPIAFQQq6brhvJo2GL4OL7JlFm/FIZNFj91C7hNq78OEpNd4HP45TlvfFZSJIDCNJmi6A71WN6U
u7iLtpxOTdvcHud+g6PpMLzg+bqud6kL+6vpY0+DKy27l3PQJryZs6JCDAir62/29cfydpDLjCJE
rHvmRbOnwTPfoxHjtoEMb5AbugPVv3NKHRupTE+BrAGou5zOxiFuo4DEqPBwP3omj1/ZLh/GQoYA
Po5SfLhBSlVmTEuv7/qmL5mVEL8SJn/9bgNf7VHf/df08mVtRJEZaekXF7M42e/uHKIr4ONhiEhc
PpNEwscL9JKYNxssY8NwXhhEpqvLqnumeW6hLFpBSWKRFvYhchISLswSitjeOFiLAqpHh0rM178k
JhHZ9ZJEhZPLekf2yk92pi3q880VmKw4z7Ayh9LfJPrIfimgLVrvft9XeMPRK2o+2vTIXb5Yds+5
9P8olNJmU3Kbz8HfnEEr6gQX4dvhdA7ZKBopNSRzXTPWiYejJ8gn3MPbxEQSSFPbSa77dvLNCofZ
3lIPKmvJdSnCjoV8oxWP3XeHxNe+EfqIK2uk1X5YKb4aqL4ZvFBL5rbLGatzhfkLqnDiOzonnmXD
ZW4wm7+aOWZi0AzTfqd7TcUcFQ08JCShrMHgieJzrtB0b4dVHqSilec2VKR65Z2OcTg8YYfe0+5w
eSZji455U7PhAxdrOS4r9wgLkDGCLKTd0uK4z7NwJmNroz25m4XCARqQzOm4lVsF5O8T9yeffASH
XMcOO+ThKf1i5FSs56TsP6sJiI+f973SxeA4wzIqiapRyCe6hFwbHkEKPsBlYxqekiLCrVemmzuD
LbPFR2hMk1VmP8EmT38ZZ9VbSHwzQp3+B3pvhssTHDOSLsP56pcgWzeQq9NWJOobE/TFLTO3ebnX
BsLhnzGZXcgK8bF4RRhnCbxk2s2pcAr1HW/5Ezg+E7ntncDmyVgPA+0+8RgQNtNPwZcgBHB5iXQJ
syQlq4ZZJa1iQ+0FW2x54tNH8GvIZMxi7jFqopiYwXDkQT2kez/fFHvTBM44jrOCZpFuTX7hV1zI
L/aPmRgFnJd1CZYHv3C4FhG+C0+t6wf/RwIjh/UHZH5v6sKp7FgvF8lo56h1IHR+wVVbZA15d8Ff
FHtFGN6WznCnRvANTdTspzkPtqweK22aQ5RfRVZ2pF3sqImEQwnsWL56wNl1oMmHAkqcgl531OaS
eZ+xG2wD/8w0imVQE8DyPhJHjdr5OSi8brtvpOWjp8BgEEE0P+BtChs8JfRHspuoDQHY/cgNbaFB
LYxPCykXDUCHswnnKThnL8XkPhvVoVXHveg3RWL+av7mHVdeeLgQZFs73T8t4HJTOz73qqNmxhV0
OVeNttQL07vhl4AIBJNKjp17XG+Slpngi/qVUWC+P7zRn6kL5eWxMhAop3hmyWwbloQmyBEu521e
BbVKYJexh5/Sz+ZOnuQd5thA5QnjNo1EI7dSf+bLEm1KovSCNLzIP/rhDi4bDV6WeLJOXig4Dg+9
5hlCyq8Fip236b49kaT4xljdnpxqOwnK8KBHK9fS1N1BSx68yMhaAww6uZ+RVa6J56orYfpk4sMA
0FCPHHHPM4hLtKKIxAHFco8JBVnwuqYyH9RKgiN/5X2PtHep5zKQUMIyeukyT+x1ILPSFYkUoGa9
3MAkq9+PoYIJuQHWnka74dS0TxT58MTYHprbwS15O9RvFOfqR4AD7iae0DiLmZtCl9KZTI2kgpzm
7O7zuCI+QuLat7c3vl4KHHOanYu3/t17QuwCgyjqqujrm8+6yyljG/L+MuiWXWSsn6DM387meD85
VQu4YOGwbpJEMqb33TtFn4nbxYi2ZQxQDVD1BWi4g4VY0pV8G/zIOZOl2I1m1ztTDe4zOnr2eJHX
FsCJW+8L48yhh+H81o8czFw77vfUFImtmCWEEPfmVCorOCT6KUuou2T8jL9gTGpf8B35DdE2HvbX
gCXmM+tEVVDSZv1c99+oEjS5hKQQ18XB40HcM/a7CDwkkceKEczaJTWGe0/FwjRWW0DfPRqLpkkJ
6HD9bKAuqAtLvhUc5H5/PULDYMgeDkiuMYyqg9JWqRPdIv1LHg25JKvRCEby29EXxLgf7z527JDr
AGvmSpBh2ySkOUvATMXpc+DlHkF4JljfxqZWmNskYrO5OlXdXc/d20MOp1yWbzn+sqtiLy1UErEU
N7tdTfrG8PJFgbL/yJLMaM2pgdep23N+jDhtXSvb95sjnmFkMTJIiGRiI6DH/FKe/MX942ONM27r
JAbjB5T9lmy6AF8F1CYyklKPiUuVlJ4mc7mElmWoL/DXGDgbUaBzy7KVkq8NQYV1rbCjN1z5o+M6
2CBctCoJq5C9dBmZ9Hzscl6j2toz5hXUprz89Hz44lsnBKtrRvV1pjFgdjpfBSnJTHzsEqgXqeLr
SCPTgGEgVo0Fbsg6Y9eIuRdhI7N0h02acFMytUezwqV4ghRnxPs/KAmUAkOt5LGpuKw57hkV3JQu
QFRS5FZyNXTjH/tDbDf7h4xQURB3BlmwFDqlyGK9y4jdOIRoQExd722jfYr1ZrVrqxlQjGGG7w2R
6BgNf693iGI5lGyMt6ST1BBIauebF0mcKpeUdGerOTLdNBwOgqS6eUCp0sWHYC7jkQUeyXT2xvxQ
8iIVLGl5pbW3ceah487pMfx3R6ILuNZFP2U7bIwKnlsL+Mz3wOB3Wpvs4A/kNOslN3oIR41rNl5O
v3CaRhWrh5ICgzoTDpSxQOlfn8qm4TIRY3BbWcxjTySuMbGEhAkhw4hFVjqCTnS94H8bmHJ0bn/O
7Ve21HXs0PGm7BLk6LCM73IhqtgacvG6ZY7Lz+uGX5z2z2Nzr0KnbXjMp+CoQBNr3n/YeEWXqsEA
a9sjBnWodhlHleWjr2bfOgkDb4nt8Yd4LAaLOwEEpzIlLAwqDvg4xTPnoI9bByafoaK0xxqe1FHu
09RWbyE4FdHJpmRKMHjpDNlMtQZORoNfU1uuXCrpOm8MuqhqcLNKMJQ7boQ/yu2LG5ahEh67Fl4w
dCaCpDn6SSG4pGn5B2wLk2zdqF0bnn7iOtObXxAQ7PEz6sqsW5aCz5F8QMEuB63a1m7XxADZCHCe
FdksHK2LyFh0I4auDC0357Qd8llc+b+DM0ggeoHhnSPhpGD/T7Z4s76HezUBwalKSYaVVv9V7JSU
iuwG6lAiLQoX6dmXHhbaaf2QDtJ2AtZ+yFUTHzpKPIQI2KAEyaIS1luU0DY9GIdpsLH15H4v/NOZ
uPGwbf9CH9u2GM+1FplgDfLxUxwAdUyOe5IGyRQ0Ra6talY5fzo3L2/4uS8nqvpTMKVWHZ/8XFUf
p2ZNHNuxfq17Pf747i3HiJNnYeDCDTqTL+4jD3uQXKEM8pS9M6FF0xx7hcHkWZjxs3Qv6kmlxAr+
prTR2OZzI9hSrbQsWd6+a31+/iqzgys4dTlvW0HhQ81M5u9Hen67BYKOpt8jKEocV8vfNaOlq/S+
FEHC9ZIztrsgisUaieNfSkU5mXZ30La+9KJ/2r1RWfv7LCKP3z5cOXOZsGQqggOOOCZh3/1UsvCs
Dx0bcahBZmjqtaRUpzbpYWL2vqEXEEjgCPT+QTX52rZ3f0FkXmPpwOIfKQxsGEg1RSp6v4wdj04n
XHoDPlezz4JM41KoZHCegwn3wFMYDqDS6JuzNenIW6rQgcGtrvlOzL6+2nOi5Idx4zMbOM+2El57
nIjCMeInJTJrZZRusjT/d9My/l1rK92cArKHHpD+/bQOJLVUEBqSeJa/4hvL7Ft5RVy+fp78U0eH
38omoBkcAa8QNCvVcPViIbm1wHafP5d+7qdD3dkhUnJrDXfbRmlviFM5AueeNa0UF1c4Y/LlcwFV
La/4/2h1w7OR9w7Gz6HpY2DFGTXuhEvbzsJZzd89DFrGaZPL+I9tA/avb4PUiVigpgqgKFyH1/Im
mAOsnGcneKsAIqTpeR0es7NtUbE/yX/pevXSY+krkbkeAgUyUKfjne/0Cjs4GAieo2vRnba79TzZ
K2eHKhtt70lRT+2n4Me12tdNQTM1184OGWEYChNV3XT6hIAQV8RXbOidixF8NNjp58jbcnUJyR6/
j4NKLldQFTL1v7hCz06OmG5ZAVtlajIEnmjtM3T2TLTWn65cIJNGP4avCslRzvIameKKpSADykdn
0B74N9pY0Mxqn4FVzhHzEdTAdcfsq5AuDzG3n/92p5DdpSQIY2FP/pUjWJqRC8T0bDqRHNl550zS
80BMbO7UoaaEI9k0BglvZME9i8WIUuRCVSKOfue+QOmNrkt+O6vYwR1ys8PT8wznjhyDaPyxhdZw
I9R8XbEc330LrVHA3gRfjavKI9ASrxKl77GTy68mnHt6wZu3+NTQ7Nyib5ge/mmZ9hrnCd1mDoQo
fpyqiIgeAlH+gOqb1qS0hz0W5g1So6NNp23wce5DeAVAbUoFTdnfgtPSRMe0GT/qn5GYR0peRjqk
Cea5ffHNJfur4xv/aNDYPPCWE3SCphq+wipeW2crmlJCPvEDyymm8YweGiCkkuVnOt/f2E3yzxyb
Ae7BP/CHLG5uqM30bC/urf/cBuOKLAqwRm546ByQ/jClvBq7QEAryfJLnueb+u9fe25ljHKWBMV0
0Co3iK9JtpMdSplvHeEa+ey+S0NYF7IHPObb8es8NLDev7C3DJEiwkX2YJyNOG808M6jveRzH99t
YdO/GneDg39cH35CnsuoJGUM4c6tkeB/oHkgJqcqYIDZfe2og2LKFFyxhto+Ky9dolEDjexYaC+Q
zBuK4kFIy6j+N2Z0fVD1l/NWLipmHlXL0CZg0x02f+ssXg2oSCDZL659e8IvBnFobgGHp11AmljF
00cr3KqIhcKc4KBSs+K+/D6YBr5ErKbypDFuEiEQbfh7BAtjgD0IwTSFZEMiAVp4XpPvNRQyf1ac
NIOKaKcnpTshGNXyPb4fW7ksQLcNao1v+DkGrb77k9CXliBbCI4PmIMjNVEhELmu+qwP2y0Zz2Sy
oIDNEaZ/Pd5wHPfVmq/sjvPNyCnpUgggO+kp6oAPdLD/iQm09grmwvutfES7rOwRIDrMWPM1OAr8
D9kFxNzaxQinwZOfjeOLLx/ml0raya3tFeuHJjbVNLwaTBONO1IMclOQ6uLtCsb1sIGSHU/dxoW/
Vne1meyMkb8oRBkXRO4k80IHqOVMvGG70pwR4naEpQ4u8VN4daYz31uQ6JdJXSxGXwno32LMPSsj
7XhPriv3xez+5qqE4z43n/GLKbR68uFHz067ZJpqJPs5TlGw3ISBlGN/aX36ZlJTeOfWDfbXlLBe
7/6FE5+KPfEaln906Et89AHO9xV5RzLH9XixF4UIOBCt6RcSBSGmpa7JsuxEWu8qf43qQjgSEBFM
2NadmYo0WSkaBcOdzVuU3u42r6yGs2EA32NlF8vUFB7p74gWoR5KiyoTJEoKa7A5FAf35NOY5HmX
izQEOgPPwBVaxUm+2MsmSbBEV8huIclFUvA48vZ5JWRmSU9qxMQL7CccY9vzDzE8fBHJwAkr+co1
ULspN3XUp9eAyK6goOP2T5KIy5WSHZSY5GG+RfDKGfrEnAilnpF42P+K1/9GoJABHiBbkdQ6aYpW
6Iqmya5UNsHGUeBB8267rTu5Og30/6JDCsFEFVfgmRySbAz2vLCvaOynG+IJFSAy4UKbfMLHfhax
aLLAKAHN7K5cs8v8UmwypJtFaGemCeOgK1ViVaJhC3BGndOOPJjYXlLOaoiQMNKrRR506nr+GHJk
PjSR29yXIdnhPs0SORGw2UoFP5P9HHRFtEJoqTY7zi53y+smiFWULuAYloUXOs5UKfuHwtPjRSJQ
620c16nPIEK1QfBMriDZjDQD/ChIXxcd/pLtJzjN1ArhZxmHMFGDNhlY1Xi/vpnS6moDWjc74iZQ
nOdZJNn2dHMrnUpp60DotUAwdA4hCa5n/anmAgFj2wYeJQy1mTdPHrz7zZfRgNlZGpKdIuQ3eLJ6
qfh1K/UPG5FdnYIusOgLjolx2ldPgNWeSU5ay4hMQ96BwPROOq3t3N1RqSSpVxG8BkB+fnJRoWCS
KLqCGIUiaMoQsfQ2a/VSxl1vg0glS0rhwN3nlXOjycjRPJXZz9YQMxqcw+nWVpPjGbUf0b+sxCWn
MBszh4xkZlGz6ufDCzXQvfhdZlwHffdBAqAW1SCD16VwvFVi5VGFgUz1L1KKQfeiwaM0z//RiJ3t
Pms8heZgCsZQ7zJTpJVG6nbPiSlWwsWbeNgLQADOA3SYaFIW2pRd+38hJddmF484SeT4pgfnRtxp
5chorecXDsLJRkUg3OVKQM4tQr2dyJpP4QqfyOhm6KOW81dZXsGXsZ7frNFVwT8cwSLDVrv++F43
HcMzkPImFmuTPL8naiafONim13tjqk5JqP3S5K1Yg5P032zEwDRKKL55J1q1KQpRwKWvAOMn7NAI
TjOPtzf9fO3B2YvXxoOnIcPQO0HVvyeq1DIaiaPFmV2vR5lIhE7s+ZiDzPwjyq5jm6malJCsQWKu
GmCpK8ZAbOLiSiZRjIdxnOjPbVhNPhwmLMlU2zXv0/2d0UZFGvTv4DGBXfH/sbLbCXY7aj6BtxN4
aEn0GucvlMcBKRehmyi1pzhAeuBVtnMnoBX/yUKWrOcadBb1VYiavobVQ9+r1lAvqY+Qz3QMIXS0
VXTwPN1cN6E6JQID1VgPUEkImgFy4fvPNn97PAit8D/50KaXTRtUMq18DYbQW4jInV8hdA9ODXoD
GKnc36/GoUwBImHI3ytZQBO9jf9+QAxEd7ZLP7G6Knel6sxA4NPfJS7Z6nO8I8O03AyZRNrnV7bv
/pXCkS5trua8qbjxCjzzgrt7wA0po7CY9IPS+Mc2xnlpivFLZzkkXpOK85tRWFvwawB/th8gYNbo
bQfvJ3wIxtR+0IGGcZi6PRc1ldrIv92CUpbl2LFXN9hf99HkSkHnYH6VVQA2zo5pIgraUdsiT9MH
N7cNh11y49PYkrmRDv07AusxqLBZXShyRE6wD9IAC1Go2Q9zT0s618JM4yrjbFd9gkCAWVwTbeLL
AelVlmnZ6VczVvy4HtK8lH8EHQxr535fXJQwWKvAXSSIfJOIoiJMEUXg60WfL8ETqL2KJtaGjv9F
VQ+hbkZg2SeZv/EqXd7RNjbGlRRWudCfDakxiugwQZfjLY9ibmyxPgK4hfViaetT9dJJbnpiQg3C
wxLjapJnzeD8O0rgHF8xurI2ugHQ57opD8ymjArSB9jgT/9X4WTj1AT0LmGzwg+gs/ZhurCDDgZp
fDj+8vjpVtLADb8iu2F40XuaMzNlxaI60IM6Q2HOue5ZH6RxnychEbOmt2A00xY/Dre32DO9xWtI
w63ql8W/bETibB56uFiLQqMG8+d54epRB4bZv6YmXpaemm/XXbyxb2qgkB6WwP/u6uMapsJ3bwLA
tydeM3ujlYnnU0ZJOi8eWNoyu7ZZ60X7B5Mf3kSINYemQB7nIZr3VwQ50XhTJMVQzmNBO+T51hto
2yi5LJPIo7OS0gm2jLtanXRnF/fFAn+W5rHrKxytSU5tbqgq3GkrHofbOEuXbosSilnOJc0JNQGh
qPA+Ajse3KAqwy60EVG9wmqAaDyfOJanNEEgeW54AzfZdN8q9hH/eQfzPb11HDUMhcMhsRgKwJd1
ceHJVKPE+GzobRwG0imJZGYchfuVoaCJbF50JZACoUQZIhE8qPkGg8tqM0lIgmFvsyXoAxT+GvGI
4+6hSS7Kv/Gxc/mu8MoBmsl5wqBqFRNvo3LO1LYFXS0iMbGF/G8Zlad6F/B2jgl/e8vBPboZgAbg
evdLVAALMP8AdhbaFp+7Cw9fS882vpR59xPHxCImJxa9fMiGdCcx9/y6JfuuUzau1uHouEFA2Q4w
EEbXeYOBCuYJGX1NF/tu4nQVJ43mLKSTNa4Xk7IfchV11K2GLQN5jwtTPvuPP6qwrpaJcqVyav8l
5fmyuJX2hddX3hgcsv7LX8LGfAgAXUJxgumG0Ga9641WHFZilF8s/naiugn2Ku5W3hC/e0A4OLbz
jf2ODNBxBdGDNTXEnO7OX0PXlKaTImFsRKP9elavTf+By6/DVgxI7yHQJsoj1RKskz76RsyKKnwc
6eyTLUfnQ8f7dbptsGNIsfgq/YlPAWCZwC1gk6ph1QUMDqEqukSkh+5jZz3PDA3OTppXZwdXxErV
PO7wvRL5nvSYI2+VhIqNf4lwnycsPWJecrBE6sUzsZJUN9S6XWTJiDQZzHy12drEPC5e9wEBIDh4
aJqsB9a1a1UPESO+Wxd5pFRKgkpVdfwlP6KGAMoC672W4mzLWv0lkjVnIDG7/Pay3lbvqTlqzal9
Zx5dvCYL7z7p2UuT7/6qmcyn8y0NhexkC86SuA8O/9wZAH4OJUzYUWc0RlOdZfGeLPYCh+0p4BA4
ebp0GI0CND2gO5YEesJ0tx6g7W3tnJZcOdlYODWTpngnRSgNaE2iBkcMxzOA0DTUKcFyatm8E1Vb
5J3Ju5FggFSOrO00S8gmGYXXkPEK4IZGQf+B0et+9KAcaMsi3/JF6olGHjjwRVgzBFJPCceiQbdm
1jEyTgxNotTLHGHNfFfs77Q1HpM8VBJm+hl5HF+8ZeBAD/kBv82nx99FT85KEHvAsechrDEDh8Qw
nnxo5i+Ir2b8hvu6i8ugWJk3HaOTAW6BUYg1v4s+fRS4Wmt4C+J10XuypROaz3urPvCROSph/Df7
EKQtYTFQIdf1YIHOWmDWWaScQ2jXJWxgLtgngjonjZDn2fJQ4nqGqsksVMZSsPlYaGCVzx+6Jxd/
KcQFFq45eL/39Y10lq73A9HCsGOXpwa5oRujtMgnzWMlzqSnqz6iobx4B5oikvv4hZkO/+XHW6/x
1yXbd/Pa9WzDVX0MlN5tg8i5wcXgq0a9RFtxOWs8L+b6fW/B56XNlzvU1+2scNupTCdScDnuLA28
kGkoyPyo8nGFgbzfzcLBVEvT736ekaBwk+DyQvApK9PzFBuwTmOJtg7dQkuVFXYywaNDk1ibZ6Jx
f0+WOIkQClVNYByWD7o2fUDv90+/moZnpuZheI8PyDzNOfZG3xfm/wog1HUxTs2xdwyicYgedUHA
qfHD/kguH8TkMYFKti1FzC8oYxRVxBr+hIpTCmocJpoV8uk0xK+4DyO6zMw+oMrMlwnskivFSThQ
E8HKCtowbjOhZwkdfld4TzMTWVBzamsACb27zIg89ckJrjj2R7KelSRrAY70RRUFwoqJ2D6FiO4R
WlxZhcOi64RlbBLk8myRxPl7hUaCLaxYxhlfx6vp4hqEhbOvGkqftJH+hy1zSZxzEM4dRFdCtKYO
NUD7XwaCfhAXwVK/BgjusNKCQOYqCidvTfKQbLgbeOP2QE870Xxh/2lSa79djnhB47kExUZCSkfF
2DRQfjxwpLBUEnNFd/0I4pyHPo5dFO2x3CehNhx/kVp+B/HU53nUh9uV1IYtFCw0Ua9YzZpjQyX0
dD2pZSVkezyy2JTWM5ZCnJdPEFN8lHXpxhPNgn5eSWGnrf+ppIgpJMK6WKkaw9gSnP3ErV9anYqc
oOVLNTzJebjEDFcMNoJD/Qd4opsE6qdzeEHHFZQO42zW6nixJ6qOJvMqPSIdZcznK+yyM1msdeE7
OoxgkNTOMdudQY8M+2RgzWdxM+DZX6WHr/FJDSmEwU2Ufkjx4r2tp8gkkehJ3MhpFWenhl5lWyFS
2zA0XP7RuHvXNDP+6QBGzBEMjQC0uiVcGGmGVp2dsgZkKUwnzOE7eg0gXa7BXyrTwiqVWD8afTFC
i9yTXTnch6VkRcqUE2xkXlK7rI8zutIFbzGA3xn7JVd9QqYzWzbxcgbvmMZHCt1XmJv3GtHTH0Xi
ucfD8d0Sy4FSxA3WFH6YUzW2rt3S65XjoqYb4MkzyUmFUkGD1aTSi7z5XbVO1cIsu2PNsZjA23kn
aV2cun39PRgYTxIR3vVV3RmWT2rk3nvHISQ3p0BcxzNvBYYTHuJj2EOXag1Pq1APGuvm4lmk4CM3
tHKkGz2i7syBoVl1UGuvxAYPn7Vxff0/lZ7zjU0lZoiWRX9k/f/kay80K/Pp75gttcEUXBMjmF+J
d+etWX8/XCo1NDPGM1xVBq8k21fWx4aJvmQndcRA2tWigjIsRA6iS++jAuTtvdDQxmYBQGfuRiJs
M6m3HNTtaj3J6tzMMc6pAQJLIwPrS29ouYrNe62ZZYKVxaZwY1t0JTh6m4o7n9QuUoBaTOCtLp8p
KMub/vPAkRGF0Gqd2LYW6MJ8HixFi9a20anpTPItoVmObsyYHyaBoF3I8JLdwHK5MSKzr0XKoTMG
Tw31ASk6QwUHHgGN5JiySaHmZkvxUDuIARpxxgrTXt+f8EIrkf222zXsfhKZMj8CFdfeJNsuFvtM
V0Kv0cyWHjT9x1jENKkOITIBQR4IRPAst1HAZ1YJ5J+rtkWQo7wn+oISqTqccacOiWvWg1t8mmek
8qzyZyhW7moTDocbii51cRZMhIopAHwkzO6j7JnqiJsQrSw7SA/o6LCKjt+nhYQ7rkngKFtrp3Du
Jx95yOr5XbGSUCWGRbr9Tg0wwMUBOeIBb3NLYLxdI/I6S8c2BgRb2q2v6Prd3fQW8y9xHlSRR0zp
F4GJgLYX8e0CbjUe0qjwBxboKa+TurOsinsWlxaHKD9StMR8oWmVotKuVETmi2vmj5r/kwPzL2fO
ixGNYaSjEJN+OFGAqtxFuAiuNLNBvOZI5aZ/hyT51z4jArqhOBilHfFTJtpcHYeuA5nd2l5dB0AS
x/Pd6zejkzDs+qb+/RkQudZwwW8NiJ9w46UdguvIqpGylQkdAQjID5acvyaPkDv3C5mItEB6jCQh
C6u0gxMPFgzLl44DDyKR6WY+AwChJlkrJ0Rog03fwtYcafCVtexaWSl5PV8C33ToKE0cEsuPeBLZ
pSe/BBnU/lqkjnB5VfMyRJ3sN8gJXZDaeZdSq+DbSVMO8NWmHBaGF9lX3qVyim4uMLBxll3J/R4g
urRp1D2z/dGE1sKsP4l/w57VflD9wMvJ8iFqOPGWi76HaYz40fIKQGRhIGg59bboMlw8X5BphLaa
egLq5ycahY5JX3EBybdzGBUMPsjn99aPLYSN26k2HndA8MEk7fNgoIa4xBQ/BG0kog/IuM8QDIZE
zWRkgGlAHU6voYyhjP9SxmH4cWHRLysLwqZbOGS5e2PDMhskjH/xoX07K/H35tjF1PQ/Yre6oCBo
gCNn+T2FaQcjIUh/ohMcsxwnNjuPcHnyLOLxv/6JDPAYS9bTfDyIFMBjnUY1ievvyNbGibHdmy+8
Mxa3DIKVSIb4oU3JZrvUl3Csmj3hCGkvCuCTzOXxBZ4qxErELIQGFhinJVKP+C+QSW5deuQNf7a0
Vu+TsBkul30v07qozwMW6tgY1yJ5r6M4134hpdJuAY1i4CEDC1XWXbYTpnwVGjqcWWeMkEM5YNrc
TcP6kr00UEz+ji701I22wEYQJHSpdB5+iOc3pIKWlvClk+Zz05LiiDs6eudomYTDW0ZBeVtkq7ne
O437sKs3UOgo3NHut51ciFWNR9GigVSRIK7rxVXYNNwFef9uOvJNSLQRfIK0slYeVG8ZFURz2DIX
IRO5+WD0LSMRS3f8O2m8rYEsDW+eM8vfb9hwTAWWZ9GE8Wgu32kbLyLoMfmQbfiIzaMVSdUNxunl
jSizpbP3kF+JyYZCUA8WfRfkuZuCT/aPnDDJQTDKknwKrIs3zQlDBseVjUxNVqkMM/hmHkNkIPgw
9aombU1RxcQ0Tf9RZ1XZkvIILqTypeLNSn+cFLVZ8SiGTIqULSd/YIqZms9DNYruPOw8KMc9AHdn
l3RIWrZkTWMv/nH4O1ptB+KGPZ6dB7KXt0riTD581iyZ7RKoidxETkQTpXlpohl0DQyCPOPUqR8u
ZyPz+hOpMrA4yfm+j20ZaI1TD4w0EDInP+PV/XPJsqNxZ5bX5Tk9NqUJlJPYEosrzopuPZ1CZ8cE
6gjRomdVtHCFIusy5Ot8hT2gO4dQw2DfccIGslFzm/IA/HK/LRZz84rGkavw0BTD2ajQicNxa0uO
EdCyusbcn1zl0Iw4IoZ9E/2h1LYcqLfV5mNEsjbGauxpL3s11EVfkz9G/EuIld4QN24cIYf2K3U4
fnbP+g5hbBzwGg3Tt9PTPigregmADpqOmfLMZSI87z6472pLl+axLOnIWYK1TkaqjVKUuGVa5/yL
/V3LJRemGwR9YfHCHxGDHvn9/Rf88sohBNCABt3mc4Di4G+BQsPuOE9UqujYpev6QdN+aolGLxD4
1yREhdlPS0SE6mAYbQHQCmdlUjMxfRXXC4Ena+FWwsiXn8oE0xws/8OSPbxqr21ONdIOkENF0e5v
r6QpeUVW2bgIBoNAYLpfZPSg2erg1huiVp5szpinrknS8fykp+Bgp98sWjOnPNvgDN3Rs8tZDOY2
X7ESZYb/Viuo6+u38lmXAgB87+S6XShBkbMxKoH9qHRYXfOjLhlatbtXacnFEnsWvpF68JkcDkY9
NrmPAV9Xy5SbeMLi8MeLwW7N6EnBHL3bl9jHhTtdYCyxsCW1wBevyQpK4+XPFkJWmRuRbKcxxRHY
BrMulh3Ki7CGA00xI/LT897ZCCnxDjOSfv4lKC1BpR/USugXQ/TGSomeUQ5EeEff1RECGr1uiiwO
WvZ0Rwa79dr/VHdwU/Uiqw95KQzWSIkD79ZuuYwJUeLEFeYKRCVPLz9cGWUoyFvKU6n8KUBzACdm
zqS0JM/T3DBI9Ty9zQJ+0TZFYfH7mDk1oFPU0fz2xTdswLVwtzmGIWQHOvKerW0vwXJuZ5C8Y3qD
q1oEIkxpjUxAsOgjDQ4aUQVA4q75/OntzD8KRmOFN+J1je1EqLO/mHrp8aWxIcDbEPUlfwGPkOti
6eLzLdJGEOgLuTEk+WBhU4U/O4yVNQ0j7xoOSaByX4cxdSHn/hgTxblO03+lcIpDvm44cWrGyKAx
It25awPQ17dVKlNhhUcpfoDf6JkICXi059VMJDsEar4iz/JW1itXaPfAs7BYvxRL9+ed5eyz8xPv
8d80JNPGlfCNzC/n7KsYBI8DP8c8+rKfGxiVNMbX/qMBQfWOFzrfBZ6hil5so49V0fsTsFg5CQx8
nCsei01rjaQCUGU1B/Yf9ytYqKWdy2BIQBJERzJ4IaXOcg+v7bi8M8Fev2xQEWY/ed2NJvM6HlzN
31PpHx6YyY57AAfe4xrGKmTGvkUTsOq0gszYrTZchitPz3Ddrdv8WrgmXaY0wA5sv9WpFSIQCDYD
0wdjn476hz3ffB0QGwWi77mThVEqtt/4ru2jVDImDaVO5ZCXkRvVlx1ELj/DP44Parx510QQz5mE
ZQfrybn76U5nBevG6FVwhSc06Cmgga6FB4ISBF25Sxh3aioQO4pJRl+f4DOx35dC8G89dAbbyXgO
oTADlF7DMya6dpKQk59rpFa1I1eEHiA5VVGxz0hr0++ynWBsW/0lHRq4ZX1yWL8PyYmz22Yw9wa+
1AuXo5L+lVsCS3kbiVvbWKjNAN2XhQiYuva7nTCON9OrEvZNjdZSVyaXwbT6O5eg2oWTrci1suKU
La34CDeAo6PhNRnGYyeLwZsRqs2mi8+EXwBtOU+4BX3yXHSz0O+07tuBZWmHgMKtzWoEx9P/+wAK
ziC5pYGkZ0pcvXh6TinhwEnR9TIMEpljPwlen6EwTxh+l5CEkp8MXY/FovsGsStKCGCoG8GLorn3
9uolMX5qx79D+jenSv5Dv4TxcHdxGO6P/0v6EH8rovBEcUATZNkWErLACv+C6kVCPTfSDSncooYH
249SQvsMQYyeDcUUtlQtDvJ9sDG82Ev6MNv2o3HvR7UuaIvC53p24OrcOGef09V1ufmT/Gx5PRII
5emt7BV+G/wHk7Iz6K3PM8dyWKBXdFSfSMX6q1zATHi5bFGhqSQGPEUQYP3vjA709E8Onw6iJYgt
0FmyngwWglpWPJeFJvZwsCmVgVwPeqaOMWfPDGHmCS7o66hilWMifFXDutB4IAKUh5LpmeLYe1+P
ZJsYyqA1QBhw+CXe7fhIFPMNgqtrgvKdYpHRnZbOBqrNQ75w916ZBAnt6FyvOIEZ+3G4hO5fqcaE
U9I3ebFCvpem9rPYfZxf0d0BSKno7Uv8H/0A1SyOGZCKKt9NeLPrGmJpNlHoHHw69yOPjsahiT2w
tsIyf3j1lxDQFgOwXEpcIpcmxxwdjdEStkypXYZlQjdvcyVwT/KxcelBErj5WVy5KQ3LGvmZiHUO
8kPxmdBGyMFIRHgoMAVZOvCjwguESSaZUjznrNemQnZncPSJhMg38re9gt8K+FxJicQJUfBKvaPc
LOB9ppKkWNVjTlC3L/jkD8scPSKeZIIwNwd/JFfSS5SdBtrE2ipYE7sGqIFx8tFu8cn10Cus30w4
vQ6qu6bKKarPIWSe0ay4eUyYDQ0Lu31esQ4n6O0YXITZhbyYYGsPCWB2e3cJxZCZ9pTmnhDQFdu8
X1C3fz4+pFHVud9UFcVxg00pPvP0W07pw4g794L/S0uqfbXtkNLi9Cz5qlcJYzqW1sX9/I8HSMnM
IZAsbzTHlYtmg7Dp6YdSK3vkmwPbKDZS1lljkppaiGiQqzMmL2fVUL3jQKNqdV01Bz1Sl1bxZmN6
kKr2dZXys56EnhHAnHH+Aw62H7jL3d5+Bf0rmyjsSj9fKwx4IdqWOLf36Cr6qgxg6jYNIUxRfMDO
+jDmrGrTnzzIjQJFG2ZzaYaVh1M6OK5Xb/6f1HIzyT0YcJMA0BsYhr+9J4k0z+B4tIAbsbLjgEIU
hR0Cry1p0oj+/abLotAo+l45JP7d3f+9FLb5gZq63SH9H4gtJm3U69Fy776urjIMnUBVvWQEdFGk
rDcVx0vNu7lTkB+vBecNCTUPhtRc6kNwoVQ8qV4ikVYaiF6xclPQdDHK/wWG+j7diNMqcSDJc1kf
n2YoF2mfHw6HowyQTRaE27+6q1EOqX1gKONNCYqO1xf9cgT6M9Xs1gxNW4S6kdG4vBeJz/UDSWZE
vB8qUqogPREo4+QUxPGk4bADegcx7eXD1YLqwNhLiO+nSdVI19fx4ugKOKvde6gPJGkanlurOUnI
JKuig0FWUJZjavZ0R5cgARtAGrL+zRa0LW3yIOQPMKaGRMnMT9JpOQN/MbpNzCK5WjLp116wiGFO
fXXdrSnUoVu2X87qpCSK7SBYPAQlbX8dpefHLH8+aGKG6O5uYPVzGb06OtSknue/KTjAEtoBpRkG
JHkCHj/45jmAf1ICTI5qYtBVzt7SAgtsDOFUiZBME5jysGqGquJOypTnFM+/yHaOzTcNP+fzGywt
WOr1zqbDDSyz74uIDqTg2u1l5t8lQpIeV58ycc9XiYBfhKS1lYx3QNOn018+oR/Oyl97avKAZVDy
e3t9/7vcG0mo4jR9gZIQQxXcLCJMs3thci//IJOid5TPJq9GRTP9nIbYY71nXkNKMefRLrEG1M9k
rKJpMMXBWrXbCr/OjKPrkDkDFooqi2nctSXu+hiB2PDcFYlp/ssMYhQ8A6yXHZiCQGlX2ZPpw7nH
Qtu7ffThyrubmGA6/dDTuwzAGnkCMjoI+bVGfGmqiZzC4Ogs0wv50x4ttaPVtc8KTxb+nUqcWKdm
jPVXRZe7w9Dp4Sf9RlCD9a9rxofSyUjEriBZDSBGTd7B4IZ04pT7JPXBWavHV2C5SVvSehV8GIVj
Z3QWL7BagdG8zldESMx5PcSrEpFAWRy9p1n8MoQyjMVn9onUpiVHDFIkug0IoqPGD9huIOp6FLA0
q8gNhBUzV1toMhkaYxdkkMR/hlKcOmT0jJpeNCqZ7KUh3PpYvbMAYvqe92VsC1VhRhDS3w8vrdPR
b80m4HhL8w+yiL2hh60XXcpc+SOnpJbiIYxBbz6rsaBV+mlN0Edd6GLGNx3MWytCBXnyuKqZpHT9
lRj7lMeUtEBP232DpLG39OPCv30Zuf3CM5RT7q5x9/qp5C8HVYKVYeIWh7BJ6dGIvwyFLT3E5HrN
kdJbfbRHDLBwToYAABJdK5QBmRUrxyspo8BboxmzIebIdhI4LJiyKIVaWxzLEUs7+orrwn1BFG7U
+yCUOXdLV/+WAVxU6JHXWZGDSqZljqIq+iCSt0GkxwW4bF4qLHftbSuR2PWOGCv2JtltVdxbOHOK
VNAdFvnxD53uL2q+2kdTLjg4m41y688Uw3gJMToCs5hIHQ8c5hKQcQCQfa7hyCLGF2aAumuKy0oh
efzPwUi1Oo10lp/pVSyiF1ghj9fqeYG43suCymtO/Pa74D6kttUkq6WzmyZsUk5l0TexNSxmln07
PFlZ5Xc9Djhwbg/qrKLrpVes+Z/ulJ+5l+nNtzHTCPA+Ksxav6GYLndV1I11AQ9NJQGzdYOwt/Wl
bSSYU0n8vZ8FCe2AR07kqFJMAXbivvV5hqbQ3KUZWRsCJ8RbTBQ8+R9YqPT9Kn9tyf3ma9g5dmiY
HV0whuee+Pc74gU3tnHPVHwQT80CgUluw1sfMp60liBiFz6zUDQ6HEkOjOSSrrfN6HJ2Eh9btoOo
08XwwBTwvtqT8cCNL0+V6x7bGBxnUH/nNsw1QHznLDsAzG+Pz8jLkenrr4To67zudVEWWDVfOqsS
sffqaE1jN5++vmzSHV+XI/jpiMTttYeX4/3QeSnlCSY8G3ShMcoxYBAXQ5JrgviQKNWdDZhopAIh
GFaMXppufFPirHPlDUNQQPBUJ/8oUD5lXDAvxge2F8yWbnHdXnN2ukt+DG+C+GSViBLhOOMW1Yqt
sG4yNEpskYtebKTXNBSBs2li0+9D3OTADDYEXuG0R85cK7YTBbhS6Ha/Za9V5mT40Z+rZ3gAofwS
rwjYObnTQPX0GN+2yOH0DipMBoNZ09taIXqUXneyKUqyK3VBlifQTGM9+houxG8DIP+/b1vaIbrj
uZ7cisZEpTwUX2Bw26eed5c+qLzy7BpbNBOjeZ/h7JVYsdSqzs1txZvGnE9NUiJzgmTt507hsoT+
5hBkeHwE8MmEL5WjqFYFZoFYChbb1xqeQ5IO7SzhDWE3pYDpUo6UpFrOSJvYKdrnj3am6OxwIQA2
OTcpoL0JVxOYv/butAr2gwguF1rdVYzNitpEQQgSyN7OLnQJyRXqpHlNtRDHPF0s7j7vy518ZPrd
4J1MbooFQrWVaq63yUaZM4n1tXzC30eSR51+iALaumRkYcBRuzGkvn73HAiTUdmLYrlFDT8aFotY
OdZih0dV2rXpeYvFrtqMgvL6wj8a3zkX41nzSUuKxzPDQMSdfe3QymY2r9y4oeHQi8mMCX6y66qJ
Z8YWm1VRAWejHK5/QF/NX/jfWR6kQ+6cKjHRbJXjSUIVPYCSdBrerfVUk9VYO+L+HlBFyQqjozIL
0b+cW0nKP16UDJlS1AuUSX4ltcmbeS+pXuzwtbaDPK3vuTtm/fZ5yfzU/LPBCvB1UG8V4iJvUPdh
UtbbuWv/HGSP9qznZnSDgZe/qT3bhhnDvpL2TOKw3t5FCTjxIRyJmSQaTXmocvMQT3sPJnTGTAVj
nc03TDhanHNkgdjDrydbb+XhrXyuCF2OxyFLjNbvTYusQWxXxJH7ekKaqEsNeD4L5gnG+o1cLq8+
RN8aEjRO4Baqs/sMOH0UaUp4/dSwiuNhVrsrgrTOxILpq2tKsr8gAEH1UvBByGDEyOKonch/Dz24
irf1WnckxkTBXXnIzAlT+0GkaIZA9tWDpEX4Qymb7Gj+qP8NKmFCn9TfKRloNYYJjoZzLUHFf+Nt
ciYZ9MAb7xGLG3Tu/G4y7iXUMuDrRGP1rhOBDD4X65RY9b84sI5Cc+SFt7iQel5pgOP6qFKKB0ZI
UfOKTOa9QJYp6A5X32Za2xRagO+L8MSX1XBR8R8Lw4UTo57TdpVgbzDQsGe5Ty6nGEo1h1MfDXvt
HmRHF8MbMLXhl0001BFvRcZeTKZiIjVjodwMz3lfk//7RRA2v7jfKGYCde/NnBSrsnMVIX3jHlt/
mvs3yXlE4txUlawh4252zchz/oqpaqUY16JXapvm8OQS25ULRNqivlS/FHXDlajQQnz/iRm9eqgp
4UjQb9oZeKjIq9JTBYQdzweAmgudzaonlTfUP9FthinorEM3tbkTygjaCr6dJnLJ8pjOTi6H0wNG
+fSjWTvkh8jh78QGt/fQWdzdmvpFSZQo61/FKcehrxefDh69fm7gtlV07ya4acCyV/eIDBZsqIAv
HvWibCOUZj+kEjCuaqOyt48XsjEhmt4IgpsvwkyIyvcnTQSMCN+0E1kcB+sSZGRpxYOSa8WHSbNx
pdlDKJjQEFO6eYKJQ0guIdvi+nn1M5j8RmSrwJV/+vFnwzwfqA5GsvBQPQtUX7NEE+vmpCe2myLB
KijR0yJgSdnMY/12r6s8DbCGtbMGPr8fppvrhJdXz/Dz7IRTvmeQep42vcNgnYNaIWu03bJ9B/GQ
5xW+L1uwp4JRZBrEj51kKOAmnQ9mzH4Jj3CLwzM9zZ94zTRVA6039mNAVX9MLFVfus4mvmmAsEFF
3gga304YVuITOjom52Kf1+1vVS1Cuc4CAf5dFK6Ua5jtKv4Io7Z8wITAui3zL65e80BVbPxcSChh
L0t9GKXmwmWLv9b49WIAX6U+jb4ca7f6kn0jfVb8GXBsqtV6BKU/gf6QHSpBKmKxR1/+kES84ync
cjMtyOZBye5gdyWkbmL9Iu9R33ntoxLBY3wRVJMsEqVd9YSfi6KhHrF1CPGXjZUQ0Tn7YX1BvYBx
aWxqR9RbtEs8ywZagYq0QeD8ZTxt3FQR7vr9Ig2EtLLVhnDEsBCPuPWtGT1OQnV+hU3kQZK5z0KB
TDN9pSqRDx/LY86dd0j/XyV3FSH2OnrcBlYm/mH7zuvXaIkejQTBKY2a2oPqsP3BgohWPdhRSOfy
JQAryM40RH3jUykTkmyQml5c0JnqSMDbF2I+bxPuPH6NivhgtwAJVs09A/KO2CQpEvkRmgqafrBD
zalIJMnrVSComS04ZmGrPX0KsBsgXazktjVa3PL0Zh1EoaqfLMAvg/N+WCmjdhllbCFWf3W4Ruhn
MYNekg73/mL2d4gH7JdYwVbn/v+KCB3KHjkNrAUHWjlBK/j2svtX2IPcAdDvKBLUvjA23PLsxIGA
eIZE3d5QMkxaXHK8msnAnwAnEM6Cq+snhd5366TEInqm+w0iz7FQtj3kzAVKvwgdkMPepAe4EpFQ
Gw0rRUI/XjFX9uJm0bKtIIZdwlEbQ4NIlIWPFqiURFiAW5sQwqGRq+CMVZU1eGVQ5GUxtZun8+HW
GUoB7SVonbLD552g5JtZNNOaHM/2b9iT3BEq6ldjWRZmyEv6fm/erRDNlRQX9h+/IuRM33bjqdaH
AtS+4LjOWK9Vum8QKem1zrQsYRP2z2c8AwXzDzPcAwhzMturrkXhROqSYJo2fLL8mkT1ghELuAaP
f9cOwbr8+SZwFLE2NjiGNDxPkB8yIrRnOJRJT4JKWl7b+NfKOK8+pRz76liB+3NXuo/bO6E9G1YT
oL35qiSk4tfwblvYrdQF3DbHVg+cq7JaC3v54l+K0xlyAGgZeYLsy/cJSr2CYiN3GFkmYVqCZ2kR
NPMGJY/l6CfQK8XksqFQGOdRYHKji/Ud3tIWecfAf5r9x7ti3B4rNGxXbZszB8vShG79wR34Y3gi
Dbqm0pL16ynvJiwJ0Mtpq85Nm7eDTXRGyKJSiYg02HrNj4fat/iCQGvhIwWq5ndIXPFft1JrrePu
RlauIUZ7U1UqM8AWkbEf8XK4Z1anpuPvFhUFcBxaRglX/fI0EGNOIMnrgLvQThvzTU/sgoaK1c6q
UtJBT/FuPcB465DzmL2CSRKV4B+litCKmAXSnMWry3K/G8j5hRNvkw7RA5JiCO4QtaIVrRnR6Z1l
DdbLJ8lxxQNeqRnmCqIvPzNbqXswtncHr8OKK6Pi7Toua6OOJ4JMxdoWe2Wa3VARSDYM5MFA1Wt3
Q5ERLoOPAgIWs81mkR6i+r/Bjhglxp7ozu691yYZs9SV89bPX9LlJzCo8FeNVBbv+jY8oaR610gd
auqKTSgcV4+Lz9a+TeVGsuFmJAHlnJDLhldXf9HtjuJNArrdY9+BafBViV28ON/7cE15ebB5+Q9m
MzAhjZMCjQr8LIasyCIdjFIaCYXKD5PNyQv6fBh/SvlIdHgAWo6W/fGg56JMULX7VA8mcoVjYV5R
HA2TQgixVBSJYHxs8glq1q1JQCVCB6hgAbO0TcMzHsF63nbhhP24hl2oKcVf99c1ShJa0CEj10EM
AiyF3/ztsMdKgcK6gIV++YneYoX1+WyHK6Dn7hnqitlxt57g8wgV76VV/f+A020GX58VMDttjdpM
dx2NQig0npvIf5tz11iII8NHNWpEsxxb6hE+LGR4sNGedh+ULNkYUIzZVBBheZa0T393TeC6uyyb
U1NpiC6+dgWRo1+t07TlKDqRqSWwptohHJqo8fJFFP9sd7aavvxal8wz4dn3wVBcof+bU+lH/l8E
zdVgdKbymGRaoNko7QDWuXKLN+YlnKVAKh6EMHntHQadh2ewklgKQLJtfYvAT3srwHv9phBeQcwi
ikuNwiEtWZUFOuT70TmbxzWsKR2Dd5tInx9am2ufXNlvkbBBcJK96XR0iqUzvccwNf4h1tNqaYt6
zdqTKwlNg4BR96rUjTAKy1WysLlXr8/8msjSYGnqdV1I33jWfx6gwcl5Bhz51LL0wg38YaPxFuS5
pWuZ++liEw8l59+KRsMX/n6BefuROernRCB6vb/2LEmaxq1j1v8eR0nSPc4maxbRmugzUp0FXOw2
HyPWRH+wAAmFcPpwTFNqgqOw0doSz15G4C6ocrLFZ/230LPmZ+oDG9DY2ZTMnh1egw9ZPbSrhPxE
lnhwj1rXwdYq6X2jJC6fIAqB+gxRzzL82wwzzOZa0hH+t1IOFRQmGnJA/35ADgrpUQMV199HAb9P
UxMwrGjuUJpFv0EJmElYcnLTP5XJvDGoHCcfv2U70V7EpqcEN7XZy+kzkP34pJAeI0yZ2tpSevgo
fw65E67emz9x/IBs0saeuwejIOnafPqGEuuFlevjzbylBlyc212UTuYMkrDD9OqR67/tj9L4xTwx
c9wwho+Zuza/LOmNrLViDRWqUEF6EvjBqPg/e+dm1g0nYG/ZomWU7yBiMatUJ28Lbr2oXmUhy8sq
3C6qzGLvWbDMwVYtRpYIVIdNNsvz33HPd8Np5Ucum6UvOWZBqdN8EsjP/1z9Rdjga2PAbA9cv2Zf
7zsoFMGfW8mizhK4BG3IHSAei9omVQ1WS0Vwh92C0iOH65Z7MjlDvRRVjh01e+S/AX086KOe+jwo
UPaffIH5PCEoZaPLtnpS7SKam1u/3PnM5UdJp7CW5BoZv/FxAVojZgsMln7kdAcvTzt63/hVtutE
VausvWJESW4K0Ud/2nenK336XwRP9ep85lOw4YuTZc1vy7wOfzJF29s7IyiWCSz8SZg6IFIdESGK
9Omfuv0dLkvCqIsQAp4rutYEZqlF+hicUlVyNiYByF0Q268o44g+dCFW09mfKrfQelfyvR6KJdqn
H1drVj0yMCj9ZMMsZIoG8NToqrAJuc/7DhK9eWCVbRKNuFfX5WA+vw0LPc0rsTW1XaMkcaxUGG+M
GfbrJdssQ6UuzJKERlMf/mnHcv6ehedhfwxs1Xa80420idtm02dX9xEcsHvC9GAlDe5D+hdRxGI8
0/3zUNNqT88ItLcLGRWM3DY2IPEZ/vhWvZMjU3sEZeY8WU2lGKoBaFWVqOmRZ3enVdAUWbHZRCWV
K9pAFOQWp/Nd3OEEUXZvixjhpRHHmUaYfwzIcqVpatGehrCR2GV/AEGYnYHWqUWRIHIGasuqlDFU
yLsGYB306x7dpiVUVIoHaNFo/h/9e+TOOfqzPKIiwjNPQrb+p2XhqJ8eg7QyfMnVPVUnrhqabY7Y
OpEQPsffqpHnErsfrLRIaGK0eo3I85Nblpn61+ACUaWxu1UxPTlbFC4g8RDu9QFtW66e7QT+RLw3
sBBa2dA27Ufb9kH9Tjbn/CX4Hpd76hEAviqymYhhnEe7NX4pjSNITZ9rRnmWRlDwz/9vJuSqbWFu
q6TAXws229hhmlbItyrcuBUW3p1KTUXxM6pO06Wbc7JrXIM8qyKifUAaLBxp71ta1sCmRTSSNGCo
UWuJcuwP2raIA1BdNiK71+SfjAD8Im1VYHS/t+R0ZgBYZozrAziQPDMqEXVxYkWUX1nUqFWzkK9P
Ep2FoWM/B3ntKyKCUYX9WbPLYy5w6lgk/0XGBfVuskecSzEYiN8nZpn3po+F+kMIHm9jb3Ov/hCn
wJjnFsKi8OdiJGWeZteVujS19GuMIP/X47fteLkwPxVcHUp9LZN15HhlZ+mkFreYkRYhniQK1Kax
yctRUiM1e4TqyrTGn97eZRcnL//6vc/+WodwTiAIzmXqGQLbRLq6HF9Sc/hgaYRXwK6yc/1wu3Ze
6SLRyjZAvh/9bTd2KjuQnrMct4BDSX5y87Cuw1pe2xCTW/6k2Tv14ezLgjn+rnzH8RWadywm7G9L
pUpdsEpbVAxYb65+7vIAb6iROSivj+NUkh/97voQWIWVvDmlLqkb8RE9VztaLIUdDfO5YsuoBaUa
AMtgxMzQkZn6yenlSXt5HawuQmh4gfYxNkgi3zLvaxaxMsMo4VUJF4jGuLYOagsKzDfHfltZwDZv
dNNGmxIjwHYqrMtjnEDuJ/+lEhYJ9ixk99moqjZ2cd3SjIsED4HAwx8xoOnZvwrXFUhM68b5Sk6v
u4GdKoAC2C9bzlucza+7+1CFsIRUfMoHnZOjTF6mBhYFgRfUXpht8xb+lChcQ8+qUI31z5NZXWYX
6EnviLSt2F4iNx/3s2mwoed6MvQftxIv0BLNJLgNfQJ4a5fcrfM69ZzgDUu9xg4dp2KIQgh9K6GW
lFR0oiwg2QAr5LPTV1P3IxuQfpCbLRcyICSiJYoJ4UZYVLZ7MBWLFXGc99x57yN7H0VAhWa7Nl/9
SSVE5FJLtyPlehyj31uNSbwtDs1feGSKcrcZo3BPosTda/+xK9L/Y5SO9w+nA5LijtfrBdU+S0JG
o0QmA+E9neW1S5lVAQiwsXLeh2P8/bPDSK1iiXMWZMqIO83KY1zLkHSxwSZp2b7h8Ah/Iv617Cbk
bmg3AMzI1muSVt2CDU2XJqGYF7twi0oMQzt3lQSUPhTC+RVvvOwWgIZJSujVvyRLaKPpYfVWEpR6
wn/mL2DmecjRpOHqDgPLB3r+rMOnRCIYm2NIfei+3buLscE6RSPr2Q3uK/Xceur94U9QHk3FLg4+
0UgHyfr4+ZakqoEXv8wCjzU64WMc0F1bZ2kE/FXkkAhyBWmOeGt1rSZQLHHCxOolpQonVBqeFVdX
LZ+BsAtsNfz6FqBMvTUcf4Go14C4prrSTppkcSjg4UNmFYk3XSyBK+7HXWGPQ2jf1wqUvZgiGqHH
xpQ1DiOPMuuT1800PBQ1soLT6qup5AvGwb+dDJZc8iE8LOWMS8dMrZCHXJGOUPFSG5u/wz4Mwavo
kT5OQ1tKogPOzj7mPBq2TpEb8qVAox7VA4TDJ3Fasd14Z1VCEf9XYVCFEEUbRQXgBD1YGNWx5uGs
v5QWY+ElTKNgwMLge+g6d9EF+7y8DxRXkcyzAwBKel6zIazc0HQvIwRdGUF0DKeDgi+WaiY3dm3Q
tTzfX1jGwdzvweEjbA7E2N6Q62BufGUva9+rlQxH7hPI47TurEQute94gA6f7KuIUIQXJb2Jvh/j
+9t5weDqnfO/nt55D5aYLEmmsTz2+fNzamzEo1Ljj2v3bNkjLRlT4VvjMTzpeCw6Y5XgW7Cbo9+i
44aXNAWZvfhYzaZsafl0VsPSbAzztFBcOF3CeVxwVQCw9D/aJGO6JSdOoRaRSNWBO7pi5JufHMWo
HoInL2RAtBmM1GE/rMRnGabsuNWpn2yjQnq4oapoMdEdVRLTQHYQhqRjlqZMSbzVNknZ3F6kINrv
YhmNP7QFKHgYag+TqWdzlujQ1ekSY0tOhZxtEI2O028YTRY+o8s01wqVxRWCEpX39xANCnlSGcto
TG/A9CsgmJl1A/2/TR+V8e5XvFC82PyJqm8iDf7KUM+BWkZH7fSmTlQSlvpDfDTK0le/Bpl/b1Cm
lioUxxBOLaVEGNEZ6aLNdjt1a4Vdcal7H0WmwuGB5+ENDtlTGWdYvXDKjZsvUImPtKH6ccuBwemh
1KB7Ziq/zkMP7qSkPRvr22noluv2/f7myyWDqRMBc44hTfy/eadU6hlwjkilwgluxoIlIUcqjD6h
2YQLnDFpfi8YF5Sf73jb/d7TpRYEnI3SOuqmH3rPgLhyZKPxveP8B+YiLQVVfPi7KAMFC1QjQbL6
VWN9m4G63rM59hZwmRwwZTbi5Dr/rwNoXs4HbuR+hv8ineD9eVULkTl7qRGRecb2wdcLSqazWCnC
41EEpFWRwyTSZ1OstP4GKY6/TNIpnl2gLvP3B6VMXWJY7MAWfuiQ0VQESIWqCU4xG6inL5sBUs0j
morWg4q+RUi1cYxzLnI8sdxkM/agX7nqaRg0rHDEiAKQE9y1XH4ev3XdHpuPZUUqvE3u+dbQS3Xe
ywzwYCvCge3UYK6Clqd8+ByuZr6T0U1h+G6kzBL1+1QLUm4vQIDIwMpEYYFUwXUTcg9yxdnqkLwX
CHBVIKXEi522XBCf7F07zgACMPk3fIQNqxF5+77Ilezq8TUK5Twcnd5iBR504doKgZHCQev8ys9B
snJPWZxzehNXCJLH+8s5wWDQGfWM6DnCps32x8EWGx9aDeDjv/hfyMEPgc9C5RqqT/BEfodT/Cu8
N6Ajjxhh3YRA+cr3n1DmbKokYp0BJKpVHPiQnU/NTGruaAiDg5TtJs8lO4h28WIEZtNTmoHJT7wX
aqJtB2VYR1o4ZAz1YG83gJOTfHx1hCd3wOiLLnh8/PmGjSmk/up+6uYDJBK1uQ5HUi+NFVgDnOmS
TqhTRLH7p4ApiYatdZOgrfxKMg+2cEQeTbTEMNXbaNm9XgWRoXD7ii++boKcrl52HORjrAxB+tvf
6zWYU6E8Zqr27guhvvw+V+MVKzTMufgNeCia65+ds10zORLvRpH77lI1P9AvLe9/z043yKLK11fp
3f5kHv6kl+D9Ut2sc2fOvIyPn9jlX0Z8ATqY53PvuxPleNnIew==
`protect end_protected
