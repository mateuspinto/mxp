��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���^���IѼ�E{g{�^�����w*��0�%<�(���Sh=�)�5��	v���㧿c.����7Bo�^j8�P �cȣD�}!�,��-�\��"�g�:}Fӵx�-�[z�����w�8�v�����'9�j���9�����\������ ;)<�A�	�n���ZPd��Ԥ�V��V}C��&�������\@0P]��M����=��	��n�5P�J-����z���ˊ��%�&g�R���vV�"�i]��jɯ�,n�2��k�8�ǆr	� �f��椯. {Zf?�1��w�,���4\��'�1�����&�ɩw���1RW�D�0�hJ{�� iBG��b����7>P�����H�� ����M�����C1:*+�Z�A��3)f��'������.��<(Bp�k|,o��[x^E���cO�jK��W����K6�;aڪ1�B�!�&��oɯq��� �/��D4����6��Qli:ۺ	Nڀ"��UHN��zᥨ�Pء3�]��,PoPV�76vLC~m��s>��s��g�?#���:���;��?�!�O��J�����ߖ�e$���i-\���m�����J7��S����?3��o���;��/�bݶ4@+�L��d5ἄ�U��K4��<�-�ً�m���Q�01�i�Ҳ�P��z*]v[��O~����M�"E�C�P�T��Qӯ�z�6�:��:���@hT�H�.�I%CB_}+�-�l`]��������9n��P�)�#ѣ������b��,l��}�ڠ��
�[�W1�}h��7��D�L���-��IE�����H��0�O�JS�:ƎDM"7���E���EB����,P���P��W�]Ö������2	� �q&FO�=�5����Q��oØ�����gz�-2q��g��n�~�9Q�)��{��'����ɅT�k��4L�.����£u
d/���\�@yᣕ�����,Hմt+4���a@�\��uک�3|�F����7 �W���K<�\j
�dӥ���YV�&إ&�QHZ�u�~�y3|P�O�]��%YLc[K�K��X-@V��K�fB���!q#��T�9�l�,�w�e�UE�Ր�~����P�Cޚ+����
c]���|#��_'��w����yr�}�j� �)ӑY�<{��d}�/=�e�B���伒�[�I5,F��P��yP�� �#�E~�Gܲ�t��lvYx.Έ ��J�
�4�oZP�}����b#S��K��b7��D^��rK�r��b��m���4�kns��2�~��q�}���?�&d�_/ �j����%y!��B�	62�F����DQ�t�j���&��7F1�u��u6ny��1�R1�V�O���k�����P� ְ$q��Aa9��Z_9�E+z�TQ��um���afM���2/o(�R��ws��ϸ�8tk�o�`�Y�F��}m 5���VdԐ�"��*�싅}��;"b�3x�Y���j��vs��Ў�~$P+Ăj�|���ndp9%�q�ON9ל�9��q㹉����N3*�B�S���D�k���&��f]�i|f�ۧgLT%�l0��t C���A�cC�;%}��y�	C���8��I��9,�i[#���!��&)(i4	���m�`艒\*�Ϟ�}���\�$ K��vi�RPuyǳy��K�A>��Iq����!�R�|u�]?���st��K-�?95��\=��� s��lXZ��ZOB>-�s����<S�(�̎��{ٛ��E�F���\��9�h$ȟ��	Bb,I�������XDf�����5Y^��-Γ�qm�vIb����h o�,pJ�b�+�y7BxbH8�_�M�yL.�8��g�ؔzcy�Ź��f�n�L'WjFd��J�T�2�_!T�L�#Ψ�J�Xp���v��O:�5�~ ��kր��s�hM�>�[���RU�� �7�)�&r֛��e
�c�����@��L�˻��Z�=�0J����9�1�+`���T4�!��]��{.�T��=]�,�U@7�A�#�uw�i�V��Ɗ9�f��'>}�4�����;�_��I�v�&��7���z�~C\�u�����;���O����I=��t�-��g
�#����7%aJ3�[���+��d���[X�+�"�X�
��S/E��F�u�n/���V�?Ouz�-�I]"��}�D��0���V˗��9���%|S�{!a��F/j�K�=������^U�K|+r��5F��8Mbo�Zk<�kq3ߗ.���`fp�w�2��_�<Z�ݮaqS�J��z�Ez>l�xV)m�φ���&�ĕ��Rp�*W�����|S��u��̛��~��j�|X��~. +�,,�x�ih�r,���[��^��{�)/`X��ټ �Tv��KR�X:"�'Mf0��\�-1�4]�0�/k��>�S�S��Z�]�hT<#�Sܼ�� ����c�O}��]��]�	�$G%#b!����zn�6��ǬvYn�X,�_9�m5���v�4X�:�)�#6����
�il��P��=��Y:M�����t%�LnB*�	�
�������� �ox��l�&����_��V�iؚ���k~BIf�a��IS��?������R�Kt��9⾡�PBu�H�x�����"�a��C��M�L:�C��0c9�'m�ū.�<��	���k���E���/������mu�.@ڱ'v����R��L�F�N
�8.�<�x���,VC~ �C��g�n����N[d�KY����N�"�o���� ̈v=�uIՌݩ�l�⣙_�B'��ڒ
tZG9�Z/r\�c��s:C��+��3���_+x�1)i����)���ޱQ>�g5c]��1[CEN���y�m � j:��|p�@����6L�gm@�ڮ��rɨ
t��[���A���@�an���q�`c�|���j�'�U�B�:�-�=���_�	�_��A�@�o灹�����ls���|�܊�ny���۞��h�1�����_�W�	@;(+�������p��~�w��@�$~��,��|��6дG��E�c\;����
�T�%A��'����� �����Ʊ���&�|ƻn#9�Q�_�?��h�%~�NgѨW�kŻ�'�%#������ۜ~���	
j��8Vb�oe�MY�%o�l�j�T	~���UQ�g���!���������X����^�9��>!9�ڇR�Z���d_�ʴX֋�I�<� �ݎ�w�i�V��7H^��Y�k�֌e���؉��@J�ʷ6�w���퉡�(��p�#lmK֔38��;A$����2�$W&�FI���k���b����d������L� uO&�5�|%�<�;�DO���� 局������p��c+�Ƅۓ���9��K �-�ߦ;>�#�O#,u�,�E69�'����cH��B�S����lvV{��d���i�iաaۧ� ȸ4zwΩ
��������!�ÿwEIu,P�YؤM��Dt9���o_ۮH%Ùu���C�	IБ����2ެ��?Mm��OQ�q�v60_3h��O�z���Vǲ��g-����L��|���k��w��a/R��݃^�����>�DѮ���� ��9nR�f�&;hR���WQcm_"�s��7o0�Z?�C�Q|QaK#�wҿ��ܾy\TV�.��#����3*����ۺ��?��iI�s3�
�"�����vX��ɪb�%L�8��U6-HW�j�,�t�ȏ��!,X�A�$R��t��ؘf]h9j_� �{S`��f��2�(�^)$����7r�tD�2��fG���d�KL�G	����`
�O�c ©��~4���Bŵ��e��������5I9��Y|���TF-,(=7�;��d�t����U��$*,���a�e'���}[�I_�$�)i85k�[����y�o(I��7�1i�qr��-�Xx�t�fȪ�^I�5QG=uVF����A<aE�^�j͊��DY��bc�x��Fe��$��|���E��wUs�$���S���ղ�[���p��Lg�<de��@��G�����Eb�Q<C�EVB�>��x������t���X��*�-���;����U���F�ڣ
�|c�� ��y�gN�v������ӗ�Ͳ#�Һ9�~+TTt����F�Z��W�c��v,w�'u���y�@f{zR���H$���W���b����6{5�"*�4�	zS�7|M)m���z����g���Jm��@Ĺ�ϣ���a"�Y.Ӷx�4���#G��g���k��V���������\S@�۝�{�j.{� �p�?���*�^��6�A��mV�c<`�����0=�_�sYȡ�/�jAm��a�M�X�Ѱ��Z6��ҳQc(�#�N��Bʾ"i⪌)�5�PeU�b�����}?� :��N��OXw��F���w�u���F�ؑӍ���5}����h`�����#Z:��W$5�T�Vq(A��&w��ks��w޽ظ˛���)IRxO��w����W<A���f�t�p��xȋW��ƋB���06�p� ��c!��+��>�l��q�p����X�p�E�P���@.��\6��L�}��ҪI`��&���)�9�H��N�qc����ռ����z����9� `��X�]��og�_��{�9�m�m�����>n��YRH�ԛUE:�-{�0�C���7aJ�h�9�c	��o��4��$,��8D�1�+k!V;A�����V��0<'��<���Ӟc�C�9�6&��1�͛�3�Oy~�����Y4�ԸDsD/:��pXRR�Kh��I���ԔQ�	=xA���(ɻ2���Y-�_'��2{��	Lz� �sxĖ5�o^Ek�q�-J���H菨��,�Z��'�?��#8T����#4��JG���b�rG���p�����W2q�9^9!�nC�N*���U�d���`nUP'z�ƶ���,�F��Ⱦ�a�Z�$��;8�0ld�g����`�c��4T 2�%�+G�ƛU�՟�˭\H�R9�]�\_.�K�ڞ��հưص��%\HZ1����h�;V�K;܍��J��A�b���3���ړdk-&y��A���>����w�o�Z.�D��6;ug��;Ԟ��Ų��p舘�ъlE����
�ĥ2�k8��(����p� ���ݲ�1��x�<�U��GU-vX{�EU�,8��/t�G�<�� �����0��\�q4�=�K�7&��wh�LX�C n��9��ɬrw��)@|I<�4	��RZC�vf��${7����1�����E9�$3]��i��I�7��bC�Z�k�B�I;��v}�˥�/�'�|�L�����/T�|����i0Jo��qW�l����.��}T8�i<�S�����=ut"�J
Wv�����b�v灢�DO��f��A=|�2��+	5,��=@d��-���*���G-h���Q�Q��2%�s��%�=|�T���������Xؓ�6�
Y%�o�d�KS�`��� ~e�t�ܖ��}ɡ���ܭ��������g�Ξy�yx��&�P�$�j ��zg���ߚ�E�t0'�A�*�H�.m�t~��C��7H�V��l^��K�iЯ8����~��"�\�z�$�Q�0�����*�Y_;�G5�ڽ/�^;%����w������օ;��}��y�Ͳc5�<�������c���deՙ��8\V��W�ls��u�İ�d��{~D$e2eg���'�м�SR���w���c����,o
�y�_�8v�ͱ��*�rN��T�qLP��/��4H�8�K+��2'���c��V���_TI#0-V��?���O��|���8�鳹���=�3_1�R��*��ADG�|��0ykؓ/�U�Y|"� �7�[���Ā*#����>�)��So��]q��?�QUq�cMՇe�.��� ��uwQ���}/��*�F�$�T3h�Xy��NU�]9��NLVl�B�q�1~K�5�������{��\�:���<~usޝ��W3����L2�����f��T�ףf��S���/	���`�$�I��ߗto�{㠛Q�ɬ�1�`�%�b����0��&k��ɘu���DJ@C�xӲ�ϒ=�ɋ����ۜC���w��,i��U��mݳ)K�&L�'ya?���tD��xm��W�?蔖��AyE�{�T��.n�~�x�Y�32?���n0;�ծ���{BB��*e4`b��C�mA�,{R��ۓ�46�l�-v�'��}�^�,� hI��۳ ��Վ�@x���]�%5l<�"��!0~A�MpO��\�����d���/ɣ�jPϫ��{�h@�}ھ%�_p�ю�U�_�B���nת�����Fx��}��߂�݅��z~1��:�9:$��ag��==~!�	���{^���%yk�Z��#�Y#?�(b���+_%�X�&TM�G��y�I�'�w��I=��:�pFfx	�)8E�.qi�Հ��@�Z��+N���8%��8��w&ŹX��&�@TN;�U��}��sX��+Cbi��#p����L�N��|Tf��mF���;�����\���dK2�cw��_؞,�R�c����i��@@��t=����ب%
��.���3�M���%[���#�3F2��,����Ǳ�nN܁�6�eݕ�s���K��U��)/G��-��i�\�1��x�tْ�g9�X�x�dl��,C������ޛH����<|�
�Ь�U��B~�Oy�	�H˳�������0�ۢ��ٶ-#��q��ԯ�����@�ZE�����8
0D���<��(I�h��L<��|�sص��u�C�[���ԋ�^�e���y`PC���Іx�|�9�<z�������@�=���w+�5[ؔ�\�`V�8����	P!���Je��Ar�"ȫ���'S���{qb]aX�_�!����`ی�	q˾5Pwf���O�n�n�/�J>Y˚��Tc6H�qh��u:�* m��V�>��6�b��N,�ź�L�!楰��/`.]�}A1�롯�O��|�tLsP
f�z����G��׀��8���-�ui��W}]g��	6� >iX7)�Ӈ�9���A6A�1f�����d�2�B��O�T���[��HO��c"��~�7|��Wψ���|�Ơ�S.l?f�}5#Ӹ�eF�aK���������th/��q�����9W��7
���#�Ζ��[��M�!�ۑNa좺 �Tk�2���ݏ��N�ܘ)������hN*x�&���Y�}��@N6�<�ޒT�z0ݙ�A��LJ{��?(��z��D�� ���~���g��E"[�5�
rP<����
�4�uH��DK��WC7��U�)x�[WS<��}�ҋř�%��y�(��W�0d�qj�b���ĸ�c��.��l�9�����i���~��-/���G��b�T1���B��i��d9&�{4 �V������[�[Ly���?��z5���$S��5,7���IԆ|ӌ?��"���"K:������$�)�����x�e�MlC22�W	{n��M%��4���^k=����z+X�W��]Q�X�f��k��z<Gg���;���we��P�(�їC;O�ŀ��G v/z�3? ��x���,&g���C�'���ŕ�	��D��[��+����Ӝd�(�c�4�p��צk�k�>	� �hD�n~� ���ZN��
��!�����݅P�s�`�=�:��D34o���7�%9�����	ܞ{����l�h�+����*g,�?�q�1G���}�5�5Wb����,�d���g��%�rP�3"'���C
Mp��	�ND �@�8)!
��uj���B �� ��vf�-�2�)���VM�rV�ȃӆ~�lx������hSe���D��_| _γ5i9��s7�|�}p�R|�9ip©�ݬ��P�����k�d��݋�$~����'�^QS��,IW�i�anA�A�"B�N�Q��Y�/�ӳ���f�!����%z�G���L�����h�=hի'���&Ǣ���3�ZS���c��8w��ڶD�9m�frT��9�ۧ]�߀�چ~~�NY_��Q
�oO��B�hי�cijL* 4����:���6A�A8��f�_HmU>��T�b��)�J�?��/�ɣ>6d�������Z�ÏD�f+ȶ���m���{'��p5��^����^[O9\	�)t��ѝ&*hΛh�z�q�&:�l��-�=�H]řI�6A�'ς�W�'(`eQ�1���1�BttԆ���(�M[�������Jҽ ��$ rK lD����SbI����Q��5P �.n��i����e���Wq�?�X�y%+p}SKU�j�-	Pk�1���R��J�Y.�4���VC��c7V��Q꿪�t}</b��g���Q��vR#�E����;�64�u_xl���K������{{S��x��>�pؐR���i#����>V(�օ� B�R��l�(=��9��÷��FM�L�ygj��,�L|�>�����cF��c.lA���|A-�m����"��u۱���J��m��'�:�mK�L禳���\��A���V���e�$L�P�m`�'uE�y� �
�V?`�'Ҫbrަ���+iL�"9�l/�e[��3)ss��1���.���t�O��"��?���9Z�I
���K���#j��I� :J?�e��%���<Y�曄�&x0������6��cU0?xA�zP��ݺ���V�|4)֬=�~p�3�ڍ��W���~B���ZM��nu��e~e��Il� C(���g�T6����2,Κ�H=-�>Aq�.����
��p�3�#768<�f
����%����tA�76�hB8�g7pCTq^�0K3�.�����cdn�5�M�Mo�4��\$�,�e�WE@�(gv��ՐZW��R���p�V�~�I9u�E�B��S���/��98��/���X(���L�{A*��$��%��MqY� �%�w��I��g�x#�<M��Q/�� ӓ��|���Ew<;�Er����(�6���:�HA-�k@�0�_PjG}���b�.�^�MY�'����-8"�_J�4���	3W�_��&h���o���ԏ�S��R�Ю�О��7M1�A�ZT��G��k5{ɦ�1k�p����j�M�P1�(�PFY���ǆOۘ˦�7,:#˷.2�`H���ъ���'�XP	[����p�־�9}�8H�W�L���D����1'��a#���!dYj<�S���'a(��Eq�),��Of�7�Ќ����u!���dT�UT��֜�E�@��.�Y���{��r�k�x��t2�`^r�1��e#��I)\�o�;��3��q���]��X�{R%�,�)�8��G,��Nm�s)�X] �~�e/��
6�Yo�|O6i�%�i���a4�'x�F��lHTKn��iZ�}���34]���Ȑ&{������v85��Ӱ<-4�?'R��)Yo}2|�dⵂɃ���1?du�?�vR�����g��)��Ɠ3)q�{���BҲ4<��SM����O:�,b=��;᝚������i7��)X1豳!�C��	IL_Pdɳ6�%����X��:�{�Pu����ʇ���m�:���������C�$�7A���X�t�kj6\��Is������W�I���ITI���M�
[��h�l�*��XZ�s��;-�&��C-���cvٴ�q�c��J�N��#�Pe�|�b[=̼$���]�Np6�+s��ʻW��XT��i�p��m��Ux��s�5B��N"��홳u��p�آ�Z��e�I��P��'���.NY�ݲ��+y}���"��Q��"��[-���I����Kġ���6�+Skf�<����{B��MR ��52Qw{��ѹ��~��֜V��G�[��)�8�fph:��c��-)0��I�ۼ��;�����-�e����sY���� Nբ�dr	98�~|��ޡ%�K�`O���B::�e�h-��� H���Q�������q7���S-x�j�pVO���$A���	|��f�i���25�Ɲ�#ŏ��}s��(��~�Π���nU54"!\f�%}�v������9���L��$#�#��{:�<ә��p�2��\��O��ł�����"�r��0��,OO]F6�|T�x}�g�Lݎ �:�<N�����`P�7y3�< ���5�^Aۑx�H��jZ�؅��ra�'���������C� ��oZT�H����B����To]S��Ɉ�{e�,�62�)G���g�9*E��h��`�5���[����RO�YQ.�X���YEb�x@P?�0V�Q>��.
g�-�G��ի"����D[}�#��\]���@�(���U���58�s@��<R�2���ߥ��sCWe#��2��|���wݩA��ݞ�-^�r[�"Ph$7�Y��/������{�p#�q_EF:8�(yjMn9@��WX-���*�r)-|�.���n�P�*v��XbR�mw��c�`�SrK�?���.|]D����!�����Y-��k6��u!���>�<p����3-�HH'�+f��P��O��s�M�d��y�c.�8�F�ȜOe�v�"6a�����T�'B�8
�/�Hو�R��P�ۜR�Z���wػ��ǧ��0VO ��롽?�J ���H��=H� �ا}'C��uaĽ����	G��~^_=�v��]׹�X�m�ӧ!Hƕ_��O�pӞjNiĔ�j�V�*A� (���_�b�?>�&Mo����?����'L?1����sT��qD�Ȯ���x;����ϐP����Yl������]>���\�T1@�m�ȍ	�-"B�AaN�ĄCb�=���ctg�D��hX��X,K���6�b]Y��'��r$tW>�����`��(���rut������K4J���t6��?�[�gI�.�Q�LQ�Jp/�,rJ)�|"Z�k�"
ڬ���Z)�C/㛗�~8�<p�B]T}dtJR��p���q�k0mڛ�S�%e�ǋ�������&���c<3�0��)����c'��s�=X9g��܏Zq��-4�[�1ڑ��ge����ږ]N�#S�������F�
i�8*�����������=�������G���'V�tm-���d(�+!L�� �否�s
m�����'�	C�n�������p��
��cw��T�[��K�-�a���r�(�Q�Fa������X�Xxx&�S;�	�`9K�Ө�3�l���Ź`�	yǐ�P75��p���C����U�SLu)��U>�{�����UT/"�SpY1�$M��v�)����#�V(�� V�;\�M窶�+�Z�A�@�ڦj}ʣ�N�3bHn{�n�/R1Yӭ+�dq�e�H�ŕ��0udŭ�� ����'����l=oWT?�[����3�'2	+��V�A<�#�/�i$���ںD��{�E�h�$�d1�N#�7�iu��f9��d�����*S;k���Ŀ��V��Xĥ��I�2����O����i>8;.�z��	᲌e#3�d`��sč2�؋���]	�����ԽK�u����Z��x�`F�=fT�޾��RD�P��J&<��xzW98}[��}*kyp�_��;�~��7�D;X�g��Qex��[ǫ�a��-� 1_kS�]���q������yP2e]%Ֆ[�ͺ�<���=����(�����|}D޺�^��W"e�)l��cP��vQ���!uu&�Ιk@�Q�4����JyKL����ԣm-9��~u�n�T�ү�	�E�׉ �Ɋ��bi�|m�"�{EИ����x���Y=0�V�н�;��<����Vz���@Qb-/��UUŌ`؏%��l*77Sٓe��`�ߗ$�`>[��[��&Z��ʔ�Uyd�L��Y�0���?v�:p�SO�mQ�Ӂ�Ԍ���.d(�%1dſHvgQl��R�}j��m�{�|��	a���־�A�;����H
&����{�2>o��>q �읞 HB~+�ѳ�VX�Ll��a��k���x�P$Ys
��Өڳ�������H���Tgod�$	��IX���t�[�h��+��E=>��/��Я���f���؀���xlB�?b�$�u���f�ہ�?r�ʾ��wn�Og���ף'��4��/��b�5܌��g[G�
��|�f�d~z?^��p�ow�E��������w](Z�5C�������L�P?x��8��c�}n�,�Ȓ�����5�cSM��B���އǸ�B�4���D���!b���a$x���[֫�%H_��yP���h�'�����v�B Nf�H��v�i��=T���&������qn3RR�����S�o�X[����V:1ƅo�E�Z����B���z�ڗ�'�ۅ�5��?xUM�П:G���yPr�O�/Z"bPi��,lH�ҵ���er�-Z�K�[���g�^-�+��47��t�6��0�����T�~�&`ʑ�(��-:��O#ɔU�5��Lym�8Y*щ�ą��N�"���S:djBV�l�'m��f~膕�w��|i%��-=,��Q�XH�p9=��Y~�,�����߼�KF����PYūI���E5&ڭ6��lÅy�6%��������͆=�޷l�:Ԕ����k8ȴc��]��_���r�м+;xRn\����������r��5�J$�"lȆe��j�1`j��"��<�iB~�_�A3�'|�,p+��������<_&���������3-�痖�aN��ށ�#�DRZwumX��� ��>i�Q�c�WQ~��̟���Aj�nC�lh#�����Lc��OU�� R2'?á��|�����m�-�Z�k��e�#�\�����؛F�t�T���o��<**�P8��(��A�WP �4_�$�ۑ##÷���4j:&i"��Oi��S~��>�X��r���s�hyF�(�TCSdl�Ou*�R�}I �?�L�3�9�ȃ87���PBB�r2�F��ܫ��u�8��� \͹��u�>�|�	g%�9�K	qi�;�B���`���64�#!�lt�8�R�p�Jb�/�p�������&�Ύ|υ�n���4�
���턽�x�O\���Z4gf;��9����䰋5�7Y���c��mi5����P�