`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
M/cEFqflqvWxG7AUDs2reTnAKS4ZhNiPtArBFnGUdbAwuDd4TtumLjbii42SuU4+/l9yD6JMECCv
8JNQg989CGxkW9lB1sQN1KvzHHjJKcrdzZyZK43L2buvn7Bc5bNhMraAguS31gp7Z9SKuBvyVEIR
s5BBjnL9mDIONfL8XIpUWk95zuPXg+TR6U3nuokwBJK25FrW4McM6CBuWNGqE5vKwD84GPbBLOcm
yOOcHGLzqNv/uRijo/iZJx0tkaYAJbb+JfLAxxJTkxfdbCYoVsuY6L5illTHI947fnM9zyKjvT2E
Fi6v8kbKbUZNlgu5Tbrh2nui0Ku9E3fFFhhorA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="ktvtArXWo75MuH79s20H1dBASmepFXm20g4ef85k70o="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 928)
`protect data_block
KJw8ttXPMnpUUXBTzLMLcC6MPWx2nCP/VstkGVAGmuTotZdVTZs0FSR3M9KjYFc+TVPs3zhUWIxG
IJ9YAFTxmFVTJE92vop52I+ZL0PbNnk95LejOMADD7TiyIrXZ8owgW/fCq9CDmsoiZ4tpvK3s2il
wmc9n5PGg1F4PLV8IXudyAaVyz2X3E/YqHXQI2fTrsHmd83Q6rKygVOcvEzzeem7tRwe5UcD+qlm
W7cBVmjhgyvaBB8gnkWeLrIBXYBvWNXZlGbWi4n7Yf0ngX21F6B4I6o2h0X0LJyicj9wgt/gk5lz
gNZphD3TWUNjVpD9TKXL3+4QQPYQWD5aQeC/ECzbS6MomZ/osS70v4T2DOGUY7gt2jKvCUHNhgs1
9stKs6my7ryaCbv+j/C2cLniXNmWJG5xqWl81GWI9f9CdXuU6+YueCYOZInIMrnrWWzLhCmaYT2e
IN4+Pesac1NrWSlZNeDSW48J5feRbpcCDhGXriwXI60Zji8AkcWrU57eJr9S0er2EKE1axVkFZf3
rFpkW6BldJi7NHybipHv0yjORLMEHuiCKMAmm9NUhVXmdEiAyh5C9HsH3q9STgHthEEYvnHT1yTV
iM1Wk0ToXnLN+P+Yi6Wxs5E0EfJjOyqKi9FCs01d6UevxZlcUHLTLxsPaCN3sacHCFo6KB66EPjV
H+iw+KHweo6+eQxP9foC73HO6UOKJs7lS0wLn5c4mUcyCOoOfkHqotDmR+Zxq1nHRrcU/c0Bo/R4
XLsbjcu8Foiu9rhikkmE6cZiYaXm32ej2hAWgZxkOrNXSnG7yWTKkpVR54sDladP2IFatoZOmXRQ
wDzfwtu8lhiMOlYh3R4HdiHtDwZwxBM2Aj4UwDscu0g69iU6kLj0/GWq2KQEAunvYciwWUpjqc9W
8zb4j51bRt5sVaaISpbSZR5gIiL8SYDXQMnd3DwTbkSJ/8lGRDKCpPcL5iiJyyfv+LSxDiphFXh8
lD84vmd9w/0MrenLo7Wv11deg6iSVa1Udp9k/K3Sf6z6PuYM9P5nzw6QWgGA8qVfJ1rojozUPN9H
i+znW5s54cEREjNO93tAIbP20jEdFQ/1jvOlQ42keNu5G3SLHGWzl+J6DmivEjqnsEI/XgvCVnjG
is5vYH2ZZTZ3yZ1RC8qhd56W0RUy5JIOLlSHGLtXbZqH+5xxn7WJ9Y67A0MWLD/DzgTVgDUpAQy4
yYpht/5/LPg4N0JjOAM5MQ==
`protect end_protected
