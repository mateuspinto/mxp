`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2448)
`protect data_block
Q8KNXBxooZVwut/AOT/hxv+w3PJsf/ZbVIXqcxRugTGAufah6IlYYOT6Uh+g31i6I0AOuWE/gSvB
0LKib89AljO/PHq8hD9H9B1jNN1ZypudnUH6MpEaDniylDOxkQqoGSl0kSjNIg4DxKqu7pvpUb+j
ygSzh0VT6T2o3mgl0cmo0tFtPJrxwEO0l9e2VLxV33SW6/UMaMGKqNImKvzabhdBNKTE3ehklZ2Y
bDCQNGTn3K0C2A3vzD20dlWcNoElXtK1RaUrDrYrKkqJx96g55sP7z7xP452KweXYK4V6K4jubZw
soHClYQNVx0eFwArommwAOowA5MauiZY/b3glkBnkenYoDLDCk1AUQXLJDe9j/4bDMHsHp+lsXdL
ijXhhZM5+jbuGWm4S+EZvy1PFb3Gb0zWY6+bi0nzNWeZBLbU6meBjyR4D1eeumBZlozhjEhXU1SU
H6gOTOjDk3rv5gpdBksEKVdMI3rp2yFFtU4Uk8Re9qqQpXCGptihDV9r9cMq1hyh/r7oZxAQQHrA
t2kNF6QlnBNzIMEdunueBq6EfgCrfFiwrvBtuFD1rM0Wks9OAsYW8AmbEt/IhMcgFquxtD5kaW4a
WZIdNiuJhnB1JLIjjWD9qjE5ehk396hLPU30/ISSN9AbelEvklxrnfPwcGMLnry5GhazKAJM5+C2
VYwvwGlLu93JPkOMj9olz6cg6TFfg89NFyXGkaAGkI2593cRB8WvQsiXQgucYfVCL8gwyi6vgtoT
0C1EjKYCBrkRsnZJN4YL4DWHUX/Mdosj2OtUYPkXoXgKokeZNcgzkoTQVy8BldoDRUQzb2gb9bBb
sGddLS4wy2Cy3q4B/fuRWiIhYIIzY7XdP9gCnV82xFAurPjYCVg4upGAHaNs5JEWdxhZeSiTiL/Z
uCYXIyyIDc2dprYDTY6nobNbiJTJS/yQF5NAZhgOsmYEPSIwwM8dbiO8/V9rwBzXpO1I7IAtZSAk
q9AHMmug+MP4kEBncorH26t0S8QPzbCR+2+HYFcbaW7LC2hr3r7N+b3H+EzwVTAA/XeyR4Z8g7md
Wguk5H/HvL+kwF9n31ipjA8twEXvpjk53jdv/6IbMEiPXaFQnqjATQ3YbH3ONWYx9NSIcnBH+9BS
0TOY/7b0RlGhEVnmU9ZI7YO/s8rbp0W/gfHJy3TGUOzBflzwiUAacudvC5lqt7gKE6oMBufpdE53
T1lvYGMgLqLEi9Z7nXVies5uTsgWL2em9Ke6KVTmbk6VEj1Mm5BDUCGZnWgIcvYCrG5emH1B4Nqk
ZDSRduXXBZLLMzJnXmeISOisCAuSy+C6u1if4MGjRj0MifZRtZC/4hOUWq4Dzb8MJ+AE15Vo73qb
TORaCqfp6VK1G/lK4ifTLQhUkC4rR+C6EM4wIsD4RjzN7o42Q2hndd8ELM5clpJLoVo99n7XKJKE
n7y3Xfy9k/kMSruJRpw3TVaIXxlWDzyXhKQWLe+n3rM89xxaroYoS70IhAKI5hoksxl4hPkinj5z
ZF8tjG9zMdtU9F5H3qadNMSw16DUVARjqQzJvlfDrPS217K9eJkmGCBVk/jSvo2t0LfSORQcEASi
ZzmVr2vEi/vE1GPm8z3WYqY5S9Q9T5sX+bKR/mb58oZceoMCioJMLKATalM6qFjAiopKcCZIcL9l
HUn7WItxR4xuw6CJBCl9OavC7DO3J++AP4N1J8XLWB/Bl4rNaE8Rni+Znj5utsdz8BImW6onWpt5
UZOeYtG9CqyHJDykpVv9gxXkZ5cKvU3pRvrKLV79kNiCNALqQdUpigA9cO7RMlEF0iCy+w0p6D0z
coAB27IODRFYCfQnk1xL4iZw1vDbsKcNViWGBZnY53+HhgbaeTKtRknX7mZXeGnOkdzB1Wq0mMXe
3Gn2CdENMGpeJfX8C0IF8ASARdLObNzqzh+HXSWlL26Fj14P3EnTyoDsyvYbp2iS4LucJbw/2qiM
6+p5GpU6KvBwuTSuJ7gunEV1Ji1hLP+bJlrDOfhAdyLNLxh+VKS7msCTZWyh34JQqMkcvVNQ5uVt
emXEfV2LgGeFMR3z5dpj9fmUYUldHdXqQU/XHLtcdiI9FztYB0SH97QCTRbhTtBmCH14NhBo/r/v
UocE8PfHnw/iBuFFmjidKA1gH4rzA1g6rbg2pH9akGMAJMr5+fAUYWh8RRSHUdboDu3ZzyrlzbYA
76WSPap6fcynCIAJioHlFknVL05pZNoFvRHmYuNaeuMJAhL7fKtJUuQg9z3TEgparJQEykHRUS4s
GIIOp96Ayz1DKR6stP8N/8hPcK9IE9DtCTbsmHDWdTkumy1CaIVh8FJrzIQh8gOe50Dt5JAy8sGS
CEHc69Q4DMlUB47J+zBxhbCfUNa+ly/h1nnqueX3f2RMXS5b19vSa3q7nvkbzbKLj4X/Nkli/NI0
BP3NiGPMjTQomiwcOGO/PnrelRJWvWigN9EnUAlnHeZGMgwQUeHjqfvoQdabenuCS74fmi3JnKOT
A4QQndZsbmGGcJMLrAGOrJ4i4V0QdDxpI4AmlNCA1JOp3hTVSVivzoQ7n/yO++H2ZJIHsswWTGSE
mU7Zmrz0jtstJ9hyWAHxcGMcOELUItbWh9EJC83zSePk2QyyoK4bR8o+wMh0NyJ5N2UQRXddwW8h
NBxrYlbVMj+El+UY3vg8oGiWAw5eX7/c7+gNn1fN2gdtFxk0MVNNqKki6lt2LgJDxb2kIXQORgGm
MeugvErsE9n8i26RCrtpx41uH6G7N06ZSyUqOszeqevTLzEDAglxwWj/dJ3plb2GYCHK24VZ7G5f
yBUsVC3d4KDerlMu56DbsNg+FQprLIKclXtY6SRfSrd13mvfirWEA5cZcRT+ahE8Q78JHuOAFPPh
3oKQl5UVnaNiTNDBdngW6VG2KKbStXj/9+K909gwAyaJKjteF1I4ztp1DOni+wd+rlO9z0e9uvFT
tmqgKXM6sPnDUoIhshv4WJC69Ylv5Ip8JEMd8ioijh4rP4YMaFI8z4hfwD1C1BAn7ngFHnklNNno
X7zo/dw8TVuwjVH704AZlQYCRCDCi4ylUz+CGsu7B1jJ40YUwJl24HffEqPuhj3H27HfjUWhklVK
dITpa9jaoz83ECbPafJDZWpIIF4GBwHmstBb/R1GSpKoveGrg0Kde1wdxfcSZsnlNmGPozr8cJHq
XxvceWPCNWh1Wf2E8uAZag7+7VIVrdWipbvPcAVi9Msk24H+7/97HjdURT1s+CPw37UR0afE
`protect end_protected
