��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���đƼ?F?7�
�=�Q)�Zi�#��R`P���qwc~._|�ѝ��{3P��,$}�,N���ہ��dtq77cE�gt ]��~
8oP@�^p˲/T��[��vq�3��	���\$9�7�
b����׉_2UID7F,;U��|�e�#�R9��TaD�.�Yv3� `��BG;����RL�FH������_t�'5u���؉{��;�L�H�-�trW�n�V�8��"X	�Kk&i����b�*H��''uY)� �wK2�X�*[�yA)BZ:��2� G8V��䤕�j�Q��%3�H_�^lpb�ڬ/�~J����
�ߩ�8��~&V#���V�F�������N��3��pLB���gU�%������K��A�I�H����R+�^�T��]o��Z�!���*�َqc�G�'���:n�s>K2$��g!U�N|%��Ξ��*�B����q��&�WN���oPØzj.��Vr���6s��_m���ΤEE����)�@=kI�c�z�#� ���/U��aA�@��OۡXh\P��4*�c&�>Z�@K9~`֬��A��+�1Hd�>K�6���5�.n��G���"���o�a�f����d���5f��R����x:����Lu��A}�$������N��BO�G����蚕���- ����	{��k���
=͕Ŷs��*��8V�L����]��Y�U��i؂?DX�e���D�]{��I6wıG]43��`X����M�9��h�z�V���:=-̟g����S�����*��7�C?be Z�seG�1!���Hk6��jy���-�{���}��i�_����y�G��\M�� �"����ׄ�^�,�*�b�෉��۪����3�X�q:!I�=���ԉ&��B.s��T��DA�?�x �sH"��P�ݼ��v�F��
����w`9:�b�*��]����b�6Y6W�v�t�'$���W=�����y5�f=���T����Y�[��uB��	}�KL*G��q�q�t%f�����:%O��	tk���2y(k�ث2��8�iq�;[BpM:f����!�c�^s��B��o��,d�>)�H��	�%�8x�vB���Z{���f-RFr ��i�<=V�߳��?6�u��d�_���It������׃>q8�U�s �k$e�a��ah����=�-~T`���_B"��c�H�����0xq�7��}��d��Ǫ-j�욬�$_��:��k=4��n�<(sN�xْ�Օ(�ڈ�[�?@h�]��8��ZiJɩPb�������VAk�.�]4C��h�'=��#b��P{��X�ҽ)�Z������6��.�e��'@O���?^�[m�<�#����սU~�5:\y֙���Y~i7��0���5zo����� <�z�ŉ_&��y��$ơ�nRq;{l����� ��n����U��F]����b(�kK�/8G�q��͔�ҹ�6�;-rgau��߿:����n6TGR�����clH�~��kVl �f�D�NE�ڲ3��4{�x/�N�r��vw{}�%yνo3ɪ�JcQ�B���_��;[A�C�s�?����{d����T~ 7Q��7uƒ�/Z���q����1��J=5N{Vs����g#)��52}�l�?�R��ôoH�e��O8�kA�,�X�{P⎃Y�l��#2Qjm��=VLΫ��a��QǎH�Vˍ܄v+��R�f�9����s6�zUd�;�L�..ٞLY�2ۜ� &�r�1�fT�M�ɻ}P/!w �K�l�$vE�pQ_N ����$/�Q�2Rm�,���7��$�ݝ_�[1QH�|>�M)/a�M�2�%h`M�q0�����2䵮�@M ]��bч���њ��E +2J5|��d��S��wS�eG�����7�K��yJ���-�;4���{c�y�G�7D�H�I��iY?�O"bw���P�'�<�B��W1C����!oa��P�?a�wO�SbP6$��M�ӵ����F���H�n�.ol�L�I���V:n�6WÙMV?�Efbr���}��dr��=Sg2��O�5[:�����0-���N�6f` �;���O�Y�����={<�+f��3:���ʺo�jj��27�M��??��OiÔ����$�SS֐.�i�����^#���K�ǟ5,�8�����3y".�#~.׻{J�n���>�me%c�31�>߅��#�/ӊ`�F�)/ihar�	 H��g�ƪWp�q��w�?Q����n?�Rczr��ר`��O� 0�g�t�Z%i�%�����-?��ӎ������2Z������OfAc>��_F����vw�D�f=%mQ^���P)��{�;��G���A0*E1�]����[g^� �ܸDd�N]���O_f�U���T��1I(�x��f��)���	����dn���Y���lf.������)���*ݗ��e����W��'�
�i^w�W�|���8MR�s~d�|��l)	
Ե��#�6uk���B���\�dL�10?K�"���W
�36�Q��J�~�F�$�z[&%��'H����`PhU~a��B��	zJĺ^E�QSơ8��鎌����|�"n��M��2p���M���3Ҭ�������|������JG9ဉ����=Ȩc�e6������9�^ �����
�%�mB���Fa���ݪ z䔁x�1�"EI5��][��J��i��,笡M��M*�$٠��5H򷸫v^�.U�{�蕵3t�QR"V�(,�e08)�A)
�>������=�6�+���a�]���{��{|���q�Y���+�}���q�- rnB�l�u�\Q���fVz�&`�_��AG-'%�SG]�����wy"-��$
�2�����1f��Lr�D���{ߵ?��ia�i�N�'ؑ��U�B}��O��`��b�h^m��T��;��S��~�;j�'8FR�́=��mH7���}ʿS�%埅v���FcEt���.Ф��U��5�����[�xy=i�ek4}�p�k;��h��Eu�`�l��\h,�5���Y����K�z�3�
�Hb ���8�r���}�s����a�w,�{�ċ�:BZ |����ټWՆ̝c#��m��=��3f|}ئ�g���J�Q��:�\�ب�;�M�H|� �.*0��g����+W�Ym�^uB��
�<ej�q= ̔A!�kV���e��v��t�?��P���"��^�ܝXj HCE�aXMjw�4 �ʗ�0a��O?vsJ�Т ��7�bLj�~vBB����пi���'k?y�4��a����G��\/	O	p���js��z?��y�)�x��8�ߞtq��^���0hDs!���� _�m���P�v��H:�ey-����N_�sA��zc*����+#H(u��,�N&)�����r���D����n5?����� L�8�>M����=�mK��h�u$�0\� !=@��0��׸vRFCێSsK����_��˖u��Kf,������u�����3h@q���X�?^(.	/�����L�+u]yt:�R{3���^Ӳ+���m�6.��wΘ<�+�2[W]P��)���ݖ,�9J��2��-|�!�g9ĐR�]6`̰Cʁ��qh=����V�6W�:baB��� ��V���	��-E�X#n�{�g��5��q��?�Ҙ{_%.�8b�_�݊�/��Q�Tŉ�u�Xa[�i�_����$�!���d~�t�`�F�C���7�z_�˺Qթ�&m�ǵ��������L�C��lJH���<M 
���?���B���h����P�����ITa/VA���m�t^ɞ(D���w�0C�;3%~��jڅb\��d�:���FI����C�w���������n�8��g��`N_! ���״I�q�C�)�u��a+k�/��ǲ���>��sqA1�U��~�FA�l�#��
%o�Y�'���n�:�k����4���F!w��>[9&�䱇�ř΋TVT��@a`q����mA�kugľ&��0�X)D�Z��	�k+��1���<�wp�Y8��$L�B�D��[�I�v�i����Q�LB���&&Oޟ������<��~�E~�Zb��3d�V��=bi��/i\v�ʛ�m�#����^��z�Z	M�S1� ^���5b�����08������ԫ���X�*�4LwFVX���ҧU(!r�H)�����0��8Щ���p՝<Z͐�B��d�&'(�ؕ��6��|���B��m=���9.Q�z�"wv�W@i��ˀ7��	�-��_f톸.Y�6
&rsz/U`��W���'=�ۍ�������)yf�(�<�=ɧ�o�	f��MIp�#���!�Ȣ��E��QyX�4�nK�j���({3*\����_d�@f�ҙt<��ǰR[���B��zd��4�P�b����i���τ��]{7-��9w
o)�)���`�R����=&x~I����ؾ|��l���n�a@Q���@�P#u�k�h��2P֫��^b,)tb��d8�3���؏�����+'wO�E���HK��ʼ
���V���wu�����q?����x��Q���6��*֨��m��k�����U����(g�h��k�(��A�#�A�"0�:�S�/��L}Н�~"���n��e�l��i_����''��3�DUё�����^	�1��2SV��@9Z��EK�-���YQ�+?r��*I��Dc�Pz�e��?Jܰ{����T���8�Q����K"�H���?�sڝMJ:�Gq��V��T��y/K�a��7�k%㮠!�ޕM5�4s=���PWd��E���Y���'P���A�����#�: ���# T��b�X� ��QK�wǉ��X�XU#��Y̳��R]ˋ�E��݅z�
#�B^6�+���!�ru7c�o��]v'{ �HG$��I��]0kWe�-Dǁ�c@�?`K��� �riH��&�[�=���xŘ�so��1@�F ܤ'm�.$�i�O6$љc5�lwZ�Mm��'��5a�75��/�3BtX��u�D���>#�R�I��1L �"_-��V�礢;�[>ɹ�7j�]�cOW*��>�@�-<b�t�F���Y�VS�`��d��P�L���xH0�LCg��$hD<��w�P���%ВHV����!�2ޛ�r�JI{*�B�4r??N��Ag1D�g��:�u/jTJW�W��6�*��ל��B���Z�r��C��}��s�0��G���ד�M�$^���"r�<��P����IV��q2A/�[ܩw2��%���zBHu��	L�D3}����2��}��=7���y��x.LlO�V�׬j����͆���S�7C�m`�CDmUo������cn?e���=��gVɢ=g�οV�(<@1=��gSB�Cl��W,k�*c⎌��l�#_-�N<	t�眲*�j�ֶY ���1�U�{�^��"|�D�&��\�~�䷃�Z�
|ԩVkB��68�K
$��.���f�'V�Ѐ@n���ͥ}�7�����[��D���Q����o
�mT�����f�e<0?��n�d��O�|6R���B��wxC����UNߵ"��E5'4N���>��J�Mt��5q6����q"�#�S�x��dge��n/���7��� ��˵?xJ��
�O��c��S (+*�i{]�9ǅ|�Z�-�Y��"A�:�װm��_�NGC��X�n=2����;Aw�ߐ�s֍]h��賂l�h́R����Q/�1�s\[�B��M�DK|�D� oG�#�O���P�7谉ۓg�~�*�B�~gZUn1텼 h)0;2	i�־���^'�2vD�K���b����Ў�,�SnD��y�xZ��%�6e��,(\\�5~u�((�C��$�	���c��%�pGw�c��WY�I��~	ϓ�@�l�
"}w�1S�rs�w�M��s��0��to��P87�Q�}!7L���S�#.@ra��1gfT�w�������x������Ӽ����4��]e��֎���	��"��,O���j 'K|����+5b�玱��C6Q������Е*6�}`>�\���B��U=ED*4���[Qd����Д!�n�)\�g�fM�Iv{���bᬋ�p	��d�������j��G�Z=�����.%��}��)$�=X�=�ݻ��������	�\a��&���XF��e>�0SP��i/�ã�����w��CI�_u�K�*J"�\3>�h��H�%q��nPYFS�I���KTiݿ��(� ���jX"8��'}`�I֎� N�|\�C�hfMR��OB���eH�����\�C��� ���w�vȰ�'����e%ɞG�9���(`	���*k�`����=�6A�)*~qS0�L���=�A�҅>�5ɝ<Iw9B���_�A����J��p�.��3�)��y��:��BΖ��`aK=�����=��A�Q����ag�}��6���3���
#�ci9j�W�{�ʵ�=�Tw`�ۗT�+a���L/� ���nt�r�Dw˼�r[���Y��ph�-6S���h�_pJ� ��e�Ó���^:���o^�8���Up������`��4�]�͸����(-ut�y|˯-���J�di�˓$�8?b�Jq.�2���5d���]�l�W9���̶��+r�)p��=�)�,���t�Eap� �u����G'e���W
�Y�_s���agݫe2��+��c�D��}������-�f+$.�:W�4~�6E�U�VME��!�7Td�c��L��F�6`�t���?{<����b�~k~�|��:�\)��_ �&���v68�L{�������ł}/��j�|��Y"��n�
2.;Yd8�"�Ga;n۷w��z�Ӿ%�E�s���%?�μ	�OZ�E�{���,��E�f�����Im~Y��R��˝w�.�-RP�	0�<�����3�_ޔ?�	-	D���!�!�>�WV�3��K4��RN���4����]،��%=yc�Y���W�3���� @w�2N��U0_0)lDշ�����rl� G�$#̵�HD j�8��F��c�9#���`�{z�ij�3���}�E�FS>~y�jRP//�u�=�<�ɳ槫��[�w�t�XZ�1�1�۴�n�.�C"�4��e�#l_�
�"3�ch�s��U{�!�+���>.�йf(w���1��݂��cC����69���,YnQr��B]X���f��>HU�"���h�Gᨰ4�=\����mU�Eڠ�!��ɿ��`l萔��{0��6{��_Xt%��܃1�4;&�|�[�k��J�:�Xx��C6��&]�d����M{?8���qW��G	�J��>r�n�`G=���-0�s1��^�0�G "޴��7�xl���5Xd+���S����Q�[��2p03�F��!�C0�& qo;y�TO/d��%��G2�(G�E��(715V�����U�P�`�`[�|¬��f��C
ۑ����?�mdy��AҰ������(�-^�3.��a��C��N}�BTM�00�Ʊvn��<qJM�2��۰(0��#���8��N(2W�1]� 0�ɶi��n�qS{���7�x���^�(/��㹃n�C�,m�/��-X��t�@�������[^	"����S�<m�����eUc�9-��j
Cc��6�=6\�\`:u`]�Z��Z:�A�2(W�����6G��Û;w��1���X��91�����_@��i�����돒Dӯ5�z��H��e�6��k��o����@av�`cX4p��g Nz幁�Koz�nBg�'���$nBuڥc`������.���eGŰѝ��`�[�2�/����~a�ҫ�� �]�=�zn��֢W�Ƹ<qŤ�q`��oʀ��2��ըg�+L@���r���2�	��Z��ӢDy��'w��c��<��ߖ**YSMPRݴ�n��?�y.c���5�?Ǖ�.S?E�;��AF0U�Ar�Q�]|��x�<ٱ�oX쳬��L2?5���v|��)�sJ�$n�Bν�JuKj����ij+�v�����+����p/�O�,FY�YA[?h;�����Ŕ~B/�2�IX�;����Pa68�֪Ֆ>.�-c���4P?1e��2��{���Ɍ�$��P��,(�2
*j4D�]�F��ލ���҆R�k�r��(%�H&c!��aV�l��6��G�Ng����cڼdyź`1�_���YF��� k�E;��Z�փM9��i`:]��D�4�bT�=��!j�|U�\JUUm�P�%��M��΃���^O?g�Л�	�;��s��ɸ̡�� �k�zC������� ��(�)	���\60G2[L��R3� #B�l@���7;\���nhm�s�6C�C����u��f��C<ԛJf���Yz�j��� "�ٗv#��<;mN��`[z�,�,n:�<јV�B�d���'���*�o����n� '1��x�jw����|V�]����ʝ��*�
Y��hQb�!�Q�.9;CL�8���A�����q�\9�[a�����������x�����m�6�%�"�����Î�E��+��C=j��<��&Z���1M���cq��f7=�FZ���g�(��$�� !�*�n�:�e`�g�5aᏀs���.F�P+4q6���*��Ⱋ�:�Q�B�!�V���>�W/��ת ��(dό�%�Av��EA?ފ�L�-�.��@��G5��2'��o
f!`��yu���8T$bApBI����:	�-=x���u��u�I�%j�3B��E�f��k{P�>���˙u.J0F�ןqx��Rm���c
Z�c7޽x���Q�Yja�����A~���@�
��p;Q_ʲiIS/�'
�8����\C�j�I��uAN�E��Xe@�JlRR;}߇���D�^���ՙ���@Tk��3z�τ��XQx��T��z?&1��K�-�̼�{<�����.Vu.�� p�ޢ�B+���~�|�u�X�ȫ���Bc��"F�4y�r���W�� q�KE�W(�_?�\_.0bk�Rc�֜�-ͺ��j�6^G*l�l�>�X`sk�@Xo҆R*I�2�S��(+CX��W��1SEY<, w���Ff����E�rt6s��u��@�p���@��^z��F�ϱ��f(�!�w|b�aE��M��L�p�b.��\=��Hb�7g���	-��R�D ���*L �M��'�S[Qy?�$�_��ɝ��޿���%�&�;a���Mu���Q�}A�e=��	.� ���L)N�ˇ��2q��������lV���;�(���^}�����~^�,��tHc>���ס6!9X�Ĉ�ŝLs
�<\�(9�6�,Z�k��eԆ0���xc�
a���� ��5�tv��C�� ]f?܋���Wb�	JYe0��Q[p>���Ib�9HBߔ &+"j��_Z��-��M˙V$4�N�����,eg_V(�U�gK𸺂���밫Cϩ/*8j�4�巩9ᦃ�/�d�I�����5��S�w�.���_�$]b�l���rJ��ԥ��q�dLĦ�ū}�(H3\r#V���S�}*����{�Քuhz��6?��z%�I$W)�z�M����� %R�/�c���� ��.~��עAb�B��
vT52��&��@��A�<O՟،O)-}*����ų�Ŕ�@�	�Cu��K:Y��l�#}�Qͥ�v�l�2|�iϛ��E)�"��|KeFn��l4���������T~�"��
���I�$O	�qm�C��>�rL�+{�_�[k�xf)5�'Ob��2�t1e�b�7�C���oyI�{y��N��ŧ+��DM4I'���Q�Zp�M�4~p�"7���M���lC�%)c����#g#*g��r�A���t`�h���&���u0����݅�{($��?Qaȓ&ˈs�*��o>I���81�W�����j���әɚ<�nJ��.�x`�Â�|ل^�����ku�D� ��d��S8��S�5t�Z��?L4��Obg?>XJ�C���l�j�s��>���X��ȷ��F�-�w�C����]Fdɨ��(�~�TM,Ĭ�B%b�H\k���R+�>q#��?���V`ڇ`&���2���'�p��oa�T�(MVo���E /��P��g�\܁ 8T-����jnݮQ��n��|QN���}��!kD��������&[������d8�i��Eĕ��a��#>�W\��(�l���T����]_`!g6����KO`h��
|r�d2+�z4b C-�뤏T���HUugL�"�^IK�߆�r��;��@�������"l�s�i���pH��ci������������"�C�At�7�Ӗ�}��0|�[Qu�W��|��<�u�M� 3�܁���	OA3��1��Vɉ�@ϻ{�v��U ���3o���(I"��pj\1��W!1P񐞸}gQT�$�0
<A�i�#�.`��h��\�h\��wR8eF�O�`��2ԮAT�b�ӷ?�o��x��=���-r�rНuqq���x�D�꺣��E�V��n0�O,��|���^�EＥ�e��@�
���OV���\?��?#��/ͯ��ϊ���E����o�l�˾L����+DGi��斻=QM�>|z_p���|�غ�Q<[>ejh�|o��%�H�e�CY�f>�6�Dn��S�T���6�|^=��yԋ�?c�떿����$���!���k$]�1���mlo��QL3��������pa�SPn*��V�h) �ѸZb�e�����I;R��G�p����@�;��s0�4�.E$#�1������(C+�qۙ��%!mG������#Ez=��d�7��/�k	�Ӷ����FMEѮ�sZ@���{݉�@܌Ɠ�%
y�s��r���~�·_�Kz��%Z��!&-1O�0�ҭ�M�(	����E�N�Ӹ����� i-��t=|_�N]�\�n�_x�Y#UF���V?���\󶥆�� J�lzO��a�s�z��=Z�'��q�8��e���>�C󘚁�1����-�、9;�3Ê���Ձn�]h���08l���5�5,���t�h����^m��^P�9Q�� �����vU�"Ka�P,I�a��H�ZQ�������E�:�qp||�	U�A5�kMf����Q�u��O�o!�)H?�r�A|�m�n��剦�����(�_J0x!�E���tŤ�`�dW���[,��v^5䲫�-�_9ۖ���+��@J�����6eeaŶ�U��$�[���l�����a��Ж���!� Fŗ�3n�╇	�
*=��0�ٷ��8�M7R����C���oD�����b�\��_��)��3��vǀ Ta��Rմ�A_�9�B}\��d/�\��(Yf�p��p��x�JeVp�[�7M���~?kP�(Qft��uӕ��{p( Z�e���!��R)믉>��UK|��n�CeS�F�3S���o�I�q��L���O ϯN�f�T�:V�R,J�0�t҇�O�9[��ۦ�����`�EQ�����\&�a"��-S�Tٟ�nA���[����H�l��2@��;y��p�o?��+in��=��0���y��ntp�8��|�&U���<?�w5���y(l
z�\8F+ĠrI��U�*V���7Ct�&Is-,:�"妠�զ70ku�\��=4��5E�IT����P�U{/�sH�rH��xP���%�d"T@�'���q�� Aܫ0s��X�$FH��V��6/n�'��ꒂN���]��G�9 ������/u�e6[0�	���D�N ��yP_C��������I !�ff��I�'�D+p64�<+�������G�_��٠y�"���/E&��a�C�Q�w�M�Β�ނ�$������h�(#'`Z
�V������ R&����j�n{f�64��&��]'i��]gH~�0sk��:޺H���.�ނi��z�]¸�C�i��j�F��|6�?�'������w`���l�WC��s�
��O�?��!y�1��\<�4�H�:���X����.�U݁������m�M�����P�������VTЩ�6M���E�z�pH�֕��$K)�ԋ�U67�L!2=>��H�θ<����{VȤ0/N�����C�cK'e�?7H�VƊ;&}���'(�|�bN1Qh��U�~�R<��ˉj�k�7��\��^���+�^�u��p�)���Z��ߎ��i��E
�������K�R��ro��,Q��! $:��F��X�-1q3���#T�	}�Fr�a��mMR0����Mh�N���Vy.D���>j��e��u���u2p�jm6