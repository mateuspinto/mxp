`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2448)
`protect data_block
+/RNe0JkEI/StdaMlxKma1XmAz2OeIH0eYa0hT5/OzILzUKePJlXEMwxairKjUUaFzMah7s4PgP2
CmAgDxabAO1O5ptphQjq5QPcvllWT+kWwLe6kwDGqCMQErCZvh5wUsZOqGCK06/UABwMKqiicrtI
GfSeJfB+TsYrY02X+UdX07ED345LP6qmR23MVaUmqITzjGTBFQyJYAF6i10VNpVZk2ac1SGR/jJG
klIq1PO8UD4Ba57nT1wfjlXLxI9+MWmKoujhaqFrXJfkNGyfl0TxOpcnmy0jLuUs6rz+W1HMYivn
zET/xxyNZMNMzTn+Zx7JIwovR/X3BcgenRFUi+9oBo1ZKvmbpOOclnLn6P/72CYb1qacUSMRogaj
SkyLx/mK1W++lzbtqprkg4vgX0s/i1/0XACKLdyVRhugjbFjHNP8AYnFa5/MVjOI8fUD4tqQh9Y4
UT9c/VTX576DC8UCa7LBkEryHHxwJkEbrMid/cvJjdkcooEpVx+tZxMMQVRRUZwVa90hq8AC4Wd4
xUugU0p0N+XqE2jJNOr0Kz5306KI8vQAEhgKpalygdUGDNTlaZTZczURQXrc7Eh2pXSi1XqFBgyy
gXc3Ic2TI0fx75sGlUIWIXa/jiHOlYJCg/wBsFM8ekadsZAA4n9gJhd24kYTjK/2fajiaGCVikBh
qYRUEF3Kyk1R0vB/rCMrwidmXQZKVo0JYghT5d1bxgb4z3hjEMDB7qCfuSZemw9I2XnBTBQTNXgg
TRhYyznzVUbKDZYMd2jAHxVvd5BM+DnQavRCAeQoBUg4yIA4+clb1y/37hQFykOG1IcnCVQ5t51Y
EADBEUtYNxVkT8vW5/Clb56/xE5idh9VxQ7Ntmq3qKn5bQjVSec+8Lo0DiXf+9QZehFSOGmgh9s5
6fEU/nwWfLsmdm95ey/fqBU7AOIhBX5decgZ00sFM7FRIQGpy011m9qyq0UTAt0TuoH9OrVR/tqY
I76Sk71T/ydPWe4evJdQB2diVVsvrI8jTZ93vIfOZM1DWrSUp5uOyflBLwMIBsil2fUOUDVYzJNt
wUjN06AUormb8Q71jT1K0Pj0cg3QuhXyGl6Rz4H48BSrr2wOwjjo8efgdBiZkTMk9PQLatDvAkvh
16jABMd+mhNIBtUN0Lj2Knmka/kSAtS3T4OyQVKKWFN2wz76xAxprkf2ylwH6JFaHjHyBoskyese
pN7DugqI89sY4eTJg5K9F/5DthBTSqWBDLXT0qzxdL9dkK4Geg/58JHiyJVV4pHlmocyIZykbc+h
JaQfgYF7crl5zBw2KZ5t+fvTMHK2HVMNlNfy1jdomqOyLD/ZCackHfAZMVRWRo6Lvu78zELz31mo
USOGTZYiwcEK+XgeDwpEnNX7JM/+AVK0u51U/AvOuEtQvukTDn0t2paxaF63t4X4Wk7m67Zat4M8
XMoXaKRaq1FQkE+J3vOZrBRVNv1VHFW6tehnjg/bV1FnEqIOVA7USFXoIOHSi9udvYOgFvnHG49P
PxpLl1Lmx5HAQuQ5w14VGImyUsGOUdylCt+y5vtxA6Y0kU1d+u1bfqXB+PO+yaw1ZDV/iwMVSFdC
GmFXXWNzRxArXKYAhfuyFmlmr21FoJxDyVUlJ1JAqipXvIng15AATd9JTbwnANlcxtDNSf2MjA8Z
GmLMVVfVMk8KiJaGEdByEidWX8bDzVm0ZDvZwjPEx0S4xCtJ0+KsoZpx/Krph9R0pL4ls1cc7KS8
xFq1WZGH8ROUfj0zdXVuOKinjY3NPLI+ifkAjX39CembWwzXp+RjAFxHTNVEIcyMat+pwQjkMygZ
SY4evrODWT1Fz43RtiIEWvMc47z2NBFwUVE06DeCDcwGBTWSV05+RKl0ogWktY6sGmCyncLUhDg/
EPulKFBRHcGtND4UWx58MuS+sqEx5YsLQ+2QPOeZRX+MiOdhuN18dkVyVlKFTTHSb0ThuvI2xc8N
KfnHCLoh4XzrfDVydYoGCy7zT2rlxowGq27bdYUrapfnqQCi9OZiPPgZ+NSSm4prjmgmxx6xV0YS
fb0ct9le80Z8oSnBGMO/X28dLS/B8tgC+7brkA0hl9R6T/fNIYU49AfZvMxXwJmgGgAQ4AXXy0Ex
8vcKi5E84vOPgKB4RyT8gRyt2YSVWHq7zRRHnfSU8XsXswQH6j+HgEtns+qfpR1EjnwzruIL72hG
flqUKCXGuZX7SMyaYWPQJkTlH5fvgp/6VtrApf4EfPTY/AYjKdlTJ+y1VgrbsdF7fMRSvNamIgJ2
JQuTV9Hc4pdzS3Lwm+c/iPwyIrLEcPbAwtQWCDhwxrle5Gg9Jztb6Meqd3FLHje8B/f1A5dTrL3b
N0TksC1Wup0136MLLqnVtWClneLWXk3FAnt5PAjFG4/alhwBETKlA511mWPSdUnCkVLFKgW+cYQC
AirjOqQ5COvgMBdb49jukViU3Z8ua7MhPmxNymq8H1UkXECICyBQ3e1BSmGahzFxgw0S3WDgVXyE
YLlQKvDVWg/ktuOtoKbjgFLUyDst9Yip8mo6N92J3Gx03MnptisnLftZgyPtTjO4L6dWZ2tD0UI9
tHkeZjAAx927CMnmmk03Fz1LdIJpKUrtpuLuFvya1SGoxdptjq06grh9tT1kv7V05J1r36+s3UyV
4VqJSp6sS2x+3ywAnxVSI+SSzDYG/BIZFofDVM/lnTdVOgXR/A5gKsYqf7MWAnkmPAqkve/Pga1M
NTsBW1pvn+bEnnR7V5MKK0ETR4wm2HMukE34MgHiFwVJdzRx4+OmaiYWvoDCjqXN4OT8WIOFpmZU
SBEIIARutLjg+UgHgpm/E7zNoNyIVUn4ZTV8rovGkUN1bjf5SHj6VDM3ovLiAFMlMHv3RQGtZ3TK
kPijidyYJ4M96EoTU+/XVxwk2HQTsuUpZu9lqaEHaPAMdMOzNuTaqiiKCI0nE8056DttGpDAHH6v
332JZgFllJfgHqPXr29Dhg28IU63BHOO6wQ207Mi10t9dfqw1KiN6dOaZustQ/ftsWh/Kmszjt7m
9aDHPcKQZgZg8z1Ps3JdGrMV5BjK6kvFCH0k4/oS+s9dB789ppA6uuO641oGr8MNMVBBB8fltU2l
NNsfGNFtKF9KMRNsHObV8+DUnQxxC5hB4+Sw7I8hxq9q/UjNll2mcUdPgan9GgmWvxuAqX2gwFnc
32NQC3xrdNZ+ugonla4WZNEm+5apTv9FAUnChxOjU08obrQaFGuzttBXWzNOuBtyhZcNVFSv
`protect end_protected
