XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���\IF�~���ڢ<��v��>rt���욈�.3z��3H�!��M�c{���dB���q���s��ܪ���0�!d���ħÏ�$����Ֆ�ѽx��o�0���?6�<lJ����f-�R����/�f�Ɨ�D�3�Q�aZ|��3��������������4"e��/2R�Vc{_�r���0aܾh������=YE��� ��F<L$�M���'�ܵ�'�(AG�J���K���I���7�Tt�g���%�f�?Pº{|_g:kqِw~X�gR�-��?��M�J	ꄯ
|�'��?���uBW'S��]���F�$�o�֮��
����.O� 9�q���TO����{���'X�?ha���@p#7YRLk�D�̞�j*��N���#�\+�`�jt&������*w6���}�3�c=,j��Q��~�X2<���B��"P��Z�{���k�Pz|���9n*��5��锯��sn@����^�V��g���m�OOl���L}9���]�c���4$e�L�XQ���D-� 1�t���	��$ �
N.mq��x����X����3���r�DJ��%se*��BP`"��5�hh_"�J�\SeG�*�	KV���'r�~�	���-��O=sM2ʳ�/^�aOe��wƱҶm��;��c~�������u �� �-�`�ރ#^`}�~�&wj�OW1�*V�c�$"LN��/B#Qo�T��_"jO�b�����(嘢�XlxVHYEB     400     240�&�(��3Ϸ�N�m%z���^�N����� �`�/c$�N6����k� >���yVisu���.;��W��T7��eO��ހ
�B�w!�ڴG��G�]}y��܎��ӫ��}Nz:^Cӂ%�H�f� D�
ـɆ۰,���	D�y�5��:3�5�+����o�t&����
�z�����_Z<�΍j�[���\�d�%���Vyp�Fx�Ж�Ii��1�r�o��0�k�̐<ۤ���_ÿ؎`����}j�3�UL+���m�4�F�S=�h�x̕J�4�k��P���nd��l�W��%l"����=e+�J�:
a�Dsn/�6�`�ڼ������ϟ�Gy�<���}t� �O��ǣ���o��H����j�ǸR�e��t�Xx5���� ��Vb��e�g�CF)����ʻR�x ��V���I���*Pi���]ن����$pO�qM�E��K`]�N�v�|%X,Y|��H���I+F�H��9�^��)�`��p����C��#���CX����뤭d�c&��K�0$Z�*���x�a��K�����XlxVHYEB     400     210��	Χ�ety5Y��rMc��f�awx.����<Qv����$
W��)N�Փ���e�N�$n
�q.d��)�E ��&�Yn6��|�z������Z<� a�j2����m^9C���e���_
zc���5f�6:1W�䲘{�U�f[f|�&_�0��P�v���;���v]PJ���	ě�P@ֿ���v�;��;��>���5l�m[m�<��7���V;�5��sU��>x�����
U�����,����.e{��M��2�(SU�!�#~,h��ӫ��{���P�uK��̕�X������?�ΉW�(������X�5�w�aZ<fs�h���R�z��A��T_5I�=�ܕ%<0�q��pٟ��]طz��}v]�sq�nk�i=��K��;GJ��fj��4�����qfc+:*+���r�Q>s�Y�E����{c�j/�����B�d�,Pb8�_MySHF�'��F����^Ҋ��L���oS~`�g%E6�|����O椫~ќS�qw+dXlxVHYEB     400     1f0�]�T Wr}Mc�F#'��8�Y=*�(�����Q'Qދ1R��%��5.1��b�+�y��U��-E�(��*�����:�ʍ_|>�!A7Щ+@\�:���ңq[���Ⱦp�,�G �΁��Cq=��z�������/;j�ʹ��-\X7zK��

���Žb�C�ד�ꡪ��Q�Kxt�.�3����%�&7��>+y0`s����Y���5��;��YƳG����y/����T�>Jk��u]D�K��`��8�N{�f�2R�;l\L��� /'��j����O�� �s�iXK�i����~r�#t�U@�@C��x|��6��r�;��C!�I���
�:���֐���=F��u�����a��8�<�jy~�uF|����43�Y0QE��]��w���'j�V����u�}+�h@���s����:�%\
;���]���:��Ʈ��L�:yv��Es�" K�ޮ���[h���o]XlxVHYEB     400     1c0���"�@y��T���Ym�b�^�zD�t��rc�H�e��Ӹ�GDr�&����= �l�%׀�����1^n�i4�ʲ���#����'~�]��>�UY�\���8��X}@�6��V��v�6������2 �=g�O<�u5F�x4yŕ�P��fZ��,a9��^ ��%�17�5�)�]�g��;��#w�f�.�q�y[ȱY��,� ^�rC�S�9�.S��6YL�\~��VB.�r��*��o�O�xש�!�3�����i1�&0ǡ�����%�$?�?�3�-&�I��9��� �ze�nDt�K�g{��:-5񧩉�y�����.ZC<%.?��F)��%LW�n�����}|�e��M�`��˚�,C�m!�<���~Dg RF_�D5˜Vʳڏ�:_<�5�X�-��������,��"�JZ��XlxVHYEB     400     200*���d2�~�eL\;3���0�#I:UiQ��q�����؅u��a��k���@{4�sWHM��s(�w�;�j:�p�v6���(��>x�R�Dv҅���W��>:��uj�`�J�6ψ�B��@�����Q�KI\R_�b���u�v/p���Q��ԃ��U�z���4\p**���{U��u��|j��-���`J3(��QxF��LZ��H�E#�ώ��O��x�<�G��4,T:w�~K��?�/�i�	ł�h���>�&D/!�Ƀ�����
`ʈ�(#�Q�5�8�
N��w��W?P+�p��yZ�Z[�8��!!���T��<�L
�ft��X���R�E���vY��ٜS�(�<A4��o�i��D��L�2l���l���������5$�@���Qt-�c���Ȫo�6�	,�9dNF'��X���?o�qդ����F�^b%����Χ���'�/e����(�)��fcT�Y������
�1��XlxVHYEB     400     120d��q"֤X��/TQ��p�9��͙_���n5��׮`�YgXV�͵�1RC���v���h����.�p	�7!�3�X�}8�l��D,��6�SrxU�g62�{V�G��̠������PD3*�7ٮ�[��͏��{��]3?�r�[M~�0����!�2�9��F��KT��x�:3POʰ�7f��[O�,�?�-]�U�\������[�g��p:�@5:��,y��Ng^�[Y���u�4�����rSS&��}7[b���<�x(�XlxVHYEB     400     1a0YB�1�ɍ:FUĐu:�j��\�����?CÚ��(�=j�Eqo��3a���Q�-�e�l�j���� ��M&�#O�h��X��V�{/�|4��q�9N8�A��i��"�x���Wa��Ӈ@^����3ӱ Չs9��� T����0<J��F�����J�=��H���甇����>���lH(�$>�����^�pm�SK�����v�35��^���		��_=�-�8��Z��b�}5����h�����.�v6��v8��:ڽ 1�3U���'�%2!7�� p<w��k�7��%>}L�D�F�'�NՍ6`*��g��c3�	�yr�f-X|�vĆe�K�jL�x}J̢0���h�� toA��YC�s0��$�o�w^e5�h��;+JXlxVHYEB     400     110�.��-�8xb�6.٪~wbHO�Ҋ�s�y�Q�r\K���:&�&�Iz�G�!|�ʫ�d���"1�f�}���7u�ܷ�TU�~�����D��x�F�[	h��n��_D�7E~�-�K6��g�
�Dv���]���:����� �x�^	�]-Eo��x�w���Z�V8X�I����>�g�Ҥ�NOR�W��d�''9�ft��Q��,$�ue#`h�9 ��1�i��.����:�I�T��Vq.~������H�R�K���2��[�'��vXlxVHYEB     400      f0����<�k$�z���3�NH��a�W*ܔX�v?�Kf%�(.�k�eG�I=Bg_j�#fzX��a28/h
Y^O^�
}��īb7 ��vzכx�FC���-�����w;�m�.{��W�)Fo���E,��9��9u��:c#�C8��U�6�~Hk�1�3(*mVi�t��о+A���͘(<�F/�6�F���L6}�-Q}c��o��ԋ� ��8��VK�FfX�̂yf=XlxVHYEB     400     130#t����;��&���q$R%M�C�i���6�	��Y�h���/HZĊ��뉇v�B����f�����o� �[Gʴ�$�v`�$-|�z���+a�;�S<gpd��88��L}4#~l���Q��ī%�I�����DIRjĲ�Tǆ�_#����,����4�#�1ܼ���~�YrB���_����OL�q[g#U�
aZ�n��J�ֺ	��qGK(&���u�$R�~�۰<D�9�$<ޠ�ڶ؉�E�����kP�
x#��YC�a:���'�`�"���Hk��XlxVHYEB     400     130V@���A,c�����1r4��0{_�K锍� �c�zr�����ޫlix>gMbrBׯ�5��籷U�E�a\��|��^�&�'+��&k�p2]�����3�rUn��Ξ�C\��?�~�����m(0�<��C|�ǬSA[S]��������/&L�@j�^ 0�$-t6,?�'�����5�w7>oF��_��p� ����Y��(G/�w��=�����������3"!�`��m/0�*x�1���� 	&��%Td��-^\�y=����a�-ZG�HyCx�����u@�˟XlxVHYEB     400     130�w��(x�4��V���(��Uh�K�k��[�y.sױ>�߉
Z:,~��{�3�>ػ��.*�Y�+:]�l����>�}�t���r��%����ȴYZ'6���壿	��-�� �F�WZ�B�T@��/�&�;��Ɵc�X�E+O���*�������ûm"SLg�#���6X���1y�.N��B�����E�3]�X;ZG��F8~���2��n���;p}��F���Ȼ')0�0�m������Qs��%F�x,a�M$)��v�πa��W�D���a=�@,Nr���e�)�?�XlxVHYEB     400     190@��LW��Gߋ�[� D��h>��n���T�>��+N�&��+���u��? �<��Td�ۘ��y%�� |��N1�s<����W�F�/�U�2ՒwASQ9(���5lY��Z5a��$�Y��ύ���{{}|��X�V!�-(��M(��W��)�n���uڗ�{� 3^$��5?�ɶ_���r�;�q�U'#%�����J��l��+�na�9J{	���%����E�vqn��8R��Og8PW3����X���G�VH|4N6cl�Dh�7����] %	���n�� v�1�<A��g���#y�x��wۋ�wV<#=M]M�e-�z]>�W;z5yj��H�r)#q�"�����㏟	]d9�÷�߉@����}f�q,
t�K�V5�h��.J�+�vA�XlxVHYEB     400     110bv��
������O����DWbX��ж�s0�����)�0]\����tT���H�f���%��U~�HK�9��V�}�Q,&b��)ן�������vj�0�_��h�n�@�����[>�t/��ƙ��?q2�j`�&' �U]���_�,h��Y�~*#���0��:���3�X~�<A��G�+��wj����;q�Z�|ee��0C8��u1������I�ٞt ͅ[D�µ$��)�hC�X�� �f�-�����=��(iD��� �XlxVHYEB     400     1b0L�Mq�=@�\�YNB1��ۛ����"���wʡ/������]���V��5�,�������e�j�'B��� �U�K8[��%�JwqE���ے.�U����� )�m�-��nOC.�%\�c�|�-B�)ؠv8�>�C�;�|Qòƫ��{�x`��$I%����@pI�|�v7Ѭ�݃�)!���X!�5�o��n�@�M�w������?���Z��?	��O���4�٦$ձ�^��yyN�8��`~�2��J�����p%(3��ί�����'%�s	l�l[����A��~��_�9��(��@��"Eu��ǈ��qс5Ы�u�hy^�AT^�a��b�� ��J��R��,�3
�{�uAן8nWm�(�\�h�w�f��i��`$��'.>o���Xk� ��0dZ��XlxVHYEB     400     190yz��o,C������L���Vh�YN0���R�Vu�&�$k������d�˴��X0�����y�mZ�t�I	����vzv�l�#��|��IY�U�c��'�Q�t&��J'�g/V���S~��cA��uN�g��m>�a 4	x�_K�!Ǘ���5%���I�.��v}%q�ű�@��<�|ű����
��Cf�&(���2��l�p�����dF|~���k4~���aʨ�˹1�r��y��^�w���'��k���J�kԶT�rY�nQhn����ᩞdB��G9�A�
�\(�������*�r�2��FIE��������5�L�`Դ�*�F�F����=�8��~���RJ�n��/��*9<�� c����� ��`�hܿ�XXlxVHYEB     400     120$9�}��lx �d[_�婆��EH������o�A�=���iW��[0��B���BD�9�N�����m�)a��Y�B$ި�t�&KA��s,#�*[��t�y�;�zF�	���
^?�޷�j���z}{��B0�<�Γ!��������緾g<���@/dL�k�k�莼��.u�Rz��J-^�x:nQ�k#����1;%X33c�rֈ�N]p>��m'3:���6�L����R+�r&Vp)�ah(1�|�����m����"�[�\1vQ�^
װ���XlxVHYEB     400     120�
�X�j�,�Ƙ4_^�'T�����&�p�dۃ��"Dx��]+0���Nڞf<L��Zc�J�Pq�r�&lU�0?ni�r�f�ڪK�j�,�b�<S�4�F��i?�]b��s��",�$�-����u�H��Ŷ���+p/[�{�=˜2�O0�P���� Z[|�e΂\��bm�z�1m
�I��Lo�)�,��M5P.�[y���ڏ��P
Ƃne�����Ơ���
��xU@ԬO@�5�guA�2�#)Ѧ�����q�C�����]��4�&�g-
�9���iifw^XlxVHYEB     400     160e��}��m����UN++�J��b|���h_��p�T�8��\ӸhY=��@�Q������yEHN�bl#��)�ɐ�_��z��*f��7��Z��9���&ۃ^�>���.�yS̆!�8HG�[á�e=��!"*�C;���f�A���
�y����7�뫔V�z-H��7(��3Y[l��)����w���l��d���X<0��bZ$���AE������;q[��e�f�=�0+JEr(�;q	��~�U
��fVT����7������N�CٶD#���"�1�P)ޛ���Hץ{�#��r9���ޥ���_)U���b�\���l�z,�fM�d]`XlxVHYEB     400     150+���ssl4�k���@jy�㫡�s�<��*�&<�e�o�~��.�i�*����/x�^���{��ܑ�Ղ��;<���~�ǘk}[u�|�c��8��g�Dn(ط����W���Q��Y�g�>u�)� �CwѬ9�$����<On����1#S�T�N����Y�.�R�N10Q����I����緗[A���"�������색�#�\"�X%�!���U?�ij��M�����W,�&d���P��$`U+�=�Lolo]��}�~#I�R�5Y,��Ӭ{���"�Ke)�~N��/=���J�lUܧ���S����dM�	��A�XlxVHYEB     400      e0�}�i���������	�A�s�}M��2�,�Ͱ�m�K�]r�D����r����,�y�X��Y6�����gT���h��D���f-^*2����0״��,'�wo���S�+Z�"�8�xe�b�ʝ��cq���S�̮s��b�9�M��Gm��q���&��EV\:�?�R�y��������R� ���*��ݺ�U�<�S��(�-���]o���8e]��XlxVHYEB     400     130X���Cj��˙�%C>Oi�2n&Z��p��ճ�f*��U�)x�+�X�[��9�D>�p.B����]�b�C!��쉿~��~0��p�Q8�ɩ(���;a����2ۖ%�G�v0��-Ȇ��
�ج��`�uS�+���>�#`ɠ�n��a�k0
r�T��9�>�2��,@�Hvb�U��Q������?��!��oEo�D[�x�*�Jw��o�b^c66we���\1>x���u."�Z_�ӭ$�.ע�s� �a�)��e�fd߈q\SW+�tO4��R���&����5�w}XlxVHYEB     400     140t� �(W��H���n�GR��AP��9��� ���p �G��Ca���!�ÂC��f���ү��8s���{�W�'&�������>�ך)Bw���YnE�e�����
Ǥ��(�
+�~����߉q53L��_qi��.3i��qɓ=���4��&Pb�}{���%uZ�Woh/uL�	顿a���?0K�_���t�a���\KI���?Fb���O7+��8J�?���i��A'�»��j�b��-����IkK-Ǣ�;��׀q����G���.�I�y+��D �9,.Bz��.�;�Ԯ*���=-�XlxVHYEB     400     150�0�[�*ׇ�Ʊ��q��:�p`���!��޻�+(�J�s������ǈmC'�RV�@�
�.�uA��e��{���i���^��v�g�� �,���ߏy�f��,�t�W=��*�ؕ��2o�]U\��E�h���j`�oo4���\ƹ�;`�u-�\g�!`[���}��$�ߴ�N5ZKJ�Hz�6�K*�����e��pȺ�Tc�k�Dd�3�/���ʈ�՞j�����/ ���u,��;`�T.��}�^�n��V�\�$��&ԑ���V<*D��g��]=�<��U��Z�x�0��۩�ֶ#�@��y�ݳe�u
KV�4�djk��XlxVHYEB     400     150J~Z���A���>�F�k����sq�7���휝$U0���_��g�t��B�OY���DSD�U���8pL�	g��ة2ߣx���l�ø����Y��ʆ�rD��?��By�`Gݠ]X_��1G��R�Z ٤����y���{�q�yC�ͫ�.�&ǯ�(�5�z:���f���7;���]9��X�x�������ׅ��t�ś�)�N/Y%F�D�%�^~�����>'
���b��U��&Mmt	>���k��s�k��Q�Ա��V�[�Υ�Q[����6�^��L�F��`�?��A��錍y�����oB��ř�A�\LS�<,�;
�C�XlxVHYEB     400     120�O�L��'��}=��eŌ��1�F��L��˛q9�~��c�Bk��'nw���B\�h���Տ��h*Y�q��tD�P�q��a9���c�w��	��>�/�b y���r�?߉�� �>1H�e�Q�|$0G׫_��R��'��:�H<;�~g2ʴE���}=�&&�0{ws��n��2����Ն�6R^0��^@�-$"뵔�춮���ٶ�Ii�8�
���N�E�&���B|�%�?��Ԯ}7c<�YP�����b�0R)o��t�>Է;�hD�XlxVHYEB     400     130.��y����aV寯�U֌�-�4�Hf���}O�����2�	�;����>*�t��2�7�1����x.>� �W�M�{X$�7$�:d���f�h��?�T��e����io\����;5�-�:�����z*�Mʻ-L�ٲA:��|]I�����]��y�9��Q&5��ᷔ忥�0���y[2r�r�O��N�n3�Wo��&�"G�6ʸ���'�
'䓺dm�]�=Y���d@�ڻ�}o�e�P:	�l��+��"1�X��p����������0��?[J�(O�`�Z�OćXlxVHYEB     400     140�{�rݲG��P�����3��(�wmCN�r�ت�hJi �8$t�B��v�u� �����^4/f獫��ݦ}-J������)B&�Ǌ�9�Td�,���8�I<����Dn�����L��_>��~N��,x۲":G�[��)`r��-�2���ۑh֥�"ɢ�L��\|�jMРd��0��4y���뷼��_'1�h�k_h���,�H�[�62CJ�}���>��E=.D|�ԝ�O�ca`B2�2�ˑ�MEf�R˴���M��,6�b�2���jI�v~
o�PW~����f�?X����d�m^��js���[�hv'XlxVHYEB     400     120�/����m��ӈ�����P���}�+���,��ϖq��� �z��Ҭ�'�;�[��ܧ����*G.�S����pA�)��.�GO[/���,���}��~�	�6(�?�=��i���B�c#�=�����5mԒF�z����}���V��i�gV�k>q*x�i��\���|
)=��jAX@j���q�lJ���+bx�_�Yt�yH�_A�q�f��0ɣ�^�#����i,�2�?k#�7�t?�����A�r1$��P�FO�U0MN"�������A��+��zp�XlxVHYEB     400     150ʣ,哒�?z���+��r��j���ʱ(oؤ��<f�#?�	�	2�u&c�LD#�2�$�ҭ�$���ߠ2����a�7��m��Vdb�H퍦Ͷ��s(�%�ǻ(�Q�Ք��o�<��E�庤�r���㲥e����fݑ`T��~t�xB��"���M�>�n�nn��9�z�DGJ��S������U�c �]��0�?u��^�S�е�-y�-[y���.�v/^��篰�&�u�=���a�e0��=��
��v��8LV����麕�>����_ٱ� ��(�*=��n�U2b���*�u H���q�g�3T�����2flXlxVHYEB     400     150k໪�/��S�� ԋ��aĦ49�S�ld���*a��._%�c5V?�R b[���8��[i�e|��@;}��HO !C����j ��՝�")F�3��V���0%c�z,��n�\Q�t�v�%}�������d��WgO:��6�Z\|#ٮS�Jl!�IrV��Y�%���)ӤyL{�38n��alT�؎�pDB���� E�ˣ���5j�G�H�	l*��	@pYu�Q��%fvICX�Γ3v��؝ӎj�F�ۤw~�5&�
-x��w���߄� u[U��VL�D��4���7'Q�(G(uYh�Вc���XlxVHYEB     400      c0�]�e�M
߃h�Usf��d�5rd������Yط�D:~�hļt�Y���"P��i�n�2`��̰�dG�Ed��Ǜ�K٥�\t5r�ɬ�o/(��s��5���?#�ܘE�^��<G�$��z������9����rg������Ҡq �K� }\��v4�3E9�*�y�$��U�o�;�M�g��n�t��kXlxVHYEB     400      c0/S��o�A�����'���ݺk;���׀`�����D[u�6zμpo�pNx(+��N�ǰ��_���m��tS��w��U�����{�>"��;׮K>Ѣ�@��u��} �S��C!�GxL5���f2:H�f�/�,�R%��s0,�&O�Y�@�-p?^Y6���=nh�<��5}�KVP:��aXlxVHYEB     400     130k�7Ȇ�WN����(���~WM�H�rU�f�ܰ���:wX8��.�P/:Dc}�iK*������tׄ)��R�%I<rV�	����H���y�t�����6D]&?!����ٍ9G2V�J�ǚ�L���#�O~�!Z	9v�zUd�%��W��̗+�]�dE�f�Ft��D���#r�M����w�"F������ʶhoUbl�}�x�8��+YϻA��E�'��� M�'�]r�&�3�EUQ�����OCC�����Mlv�fL��&l����曺4Қg|��9[
1��,toW�8�~XlxVHYEB     400     1200��K�w4FJ��	��{�����5���oE�p}�F�H�c%��ԑ�d�Х���|��"�*PC3f��>����{����#pb8����� i���z�?��CT.=�ہ���ӄa*6ct:�5!!��W{^�!i��m����r�����ۃ��D�RC=|�����l�vA�~"��?o$�u��q���e\y�vsD�������DK�;j��,�}t�h�K:DY�f��$�2dۗ_R���+�8mN�-��}�E9IԮ���-����N��e&?k�$x9�*XlxVHYEB     400     100)����>4*���~�$�,����;�LP����L�t��cߜ��]�3#��hy�������O��0�L8�٧c�7�Ě�Ĺ�Y��ޠ�*��.�j�s~����<����.��ŉ !ͲP�`HC$Kd�=k�__��h?�`TM��Ù,#��.��֒����p���7��3�l�l�|h�:$1%��\2�u���;\���T!��0�/,����S��pP�2b��te���튾5?��= 	��m��XlxVHYEB     400     160��^�q���yL�쑯]h7F�Fb(�#ZPA�*�c;�_��wFz0�F�/ \���*n=(�KE�����d�h�}a
���uԈ�R
�����XB�ut�@�
�T��;D��Oۥ�뚀>�[�q�f���[g-���N��r=c���jh�IQ�y��4F��'�(�+��?��e<V�V�/y����j�?��kh���Ht<�,����zh.û}D$��̌l;~�[�(��(��(�X���h�ž0�1�4���Yt�yߣcQ6)ܖh6��J�OH'l��*>�"х����V�-��5�Ѯ�ܞ�m�\�N�4�{�0xW���xe<<����QK�p�7Ԙ���Q�XlxVHYEB     400     1c0P"�7�U5 #H�U�r��ɀ��bw��%n}8�-�9<�$�&��lU7Ԉ�|N�h�>��V�M�_�K�Ï+�a9�E����Ͱ�+����9�C-T|�ȞŘ�`��;�FbI��?����bȣ��u�z��괘,�8��/�3��r�1K������S�6�F��	�Og��?9�����g>0~��*��}3Q��]��w
�!zo��h�'�<����\5[�8�GL�3�b��e�ͬ�Љ7�pC�wԢZ��Wb]k�drp�_�zx��� �M����Y�o��Y3���b¢�Fd\���"�Tf9��R`2����a���$ �S�ϰ�La2���y�([>����+��o��@o�F��b�� �
�Ͽ)s|t�Ή۞̎�����a$�B_N��h��Q�����l�O�{�F�ꗿk�)��i����ߟ�l7jXlxVHYEB     400     1d0r����.'�v!j�aX�	��z@��L��`���~�B���@��w��x�O+e�[�
��8���� X;���)��2g�����s#r�?���;������e�O@�znG��NH�|�O�r/�*9&"�©Kps�m<w�7l���W��8<�s�|�`��^�)ŗMS��	c*�)rF���\�4����e� �vqQ=_.sڧ籨��FZ$\��K�|.2����؀'�꫗������ 2�-,ڬ����A�ߠ��Y��{.=1�]�?%��PnJ?@���:y�� �����9_2_�oܼܬp"@�R��t=$��i{��Eq���se(N\�B=<lgL����6V	�o���cx��'t����yzelϼ/i%�I+��q��Pf��#h8��H;�~tBZ�LȒ�6ܸ�{W[.j��D�C&)�9ٓ�^XmXlxVHYEB     400     1b06��K��r�u�čK��n���(��P�k��=4f�T�,Y����r��f��T�޳��@�d��=��g�t$1ZX��I��#1� �����Ry�|@�N$�h�讦�/�6P>[ ��e����q�!�&��=�:�LgJvcba��$|���|]�B� s�l�}�(I�po��,r�˸�K��|]�2�s��j��*��mJ�4�i��a�'�Eﺓ?0�Y:��+�Z��V��s�s�d>��fJ�������"�h��Y��H���?��N���v]4V�&�F����Y^NRȶ�U\���-�������s�h6ap�Js�MR����sm(`#���P���{[��m7vqaV��
) �d�_��P�_�%���g}�@�$��5,RmX���(�EB1�f,�夢k�GY	3�ΏE}�ā�S��F���XlxVHYEB     400     1a0�1f�RҔ�흍$��ɭ�.D�,�j���^㷼gR���D�	��]nl�oDR�d��'������ݶ�z�A6���<O�B���[�d-]���1y��c�fIВ�+�bB���	�\���$񠈮>�5ԍ��r������C>_��2�^t�®��0��q�.�Pи%��:Y��P�"������Q�]j'*4'��0�P����1��ނe]����U���er�y@Ey#���u=E�g/q����n���O&%��� ��W�h�����[�K��
�QŐ�/��{K�����
�'����8 ���ʮ����A;{��8ے_��w6UB���\J�tQE���C�BZѸ�����5�Ҍ�e��G����%�@/��xt�i����u2�I����O0|��l��Sd,q�`XlxVHYEB     400     160��+w�����6ZzLf��BtW�|'j�	^��r�-v��l40�*j�������q�&�?bk�drQ�c�����\�y˝�$�M�2�;x��'��	J�U�����2!{��j��Vx���ٿL�b���`y�-s,�Sne�{܀�䃆OHt0�-��\�G%j�P����C��k���E�G�4��ol�=ho�XE-w���0O��&;3_�Ç��9a�=���9�<0_I,߀w�
]�9��*�	L3�Y�ǵ[��KN�?n�ۣq�>�Ǚ�y� �l1B�I8�aO�&�Y� V:2�Fq����	�F`~S�)��¸���:tex��XiPXlxVHYEB     400     160��j+���p��M���)\��f�(�l�0�'�*�e�9-��z~BT�qx���`̙�Fw
cY��g��S6�1��4�k����,����~��D�"�s�`��d��m?jK?�����1>�!��RB�
�)f-ţK�^#�h�@}=�w_�N��Ҋ�ď���m��C�_��"o�����aQQ=��:Į��&tK���R�d���*��N�d��Dτ��nU�ǧ�{���_�|�m��$5��ʾ����� K@O�q�hAR���������)`��m�����ۍtl�eU\B�lg�/x�ԟ���%�
M	�c�*$�]3/&@� ��G�.ٍ\��ȹ+�͝�p)�XlxVHYEB     400     180"��ܭ���=(�;?K-���w�A�.�/�,�0'wc�PSU���s�v�q���8��Pv�z_L���D�FA��P�0�z��0j}?肶&S����!�S��PT<-j�x`r���=�ע@U�՝����e�������%���%�nb���`Ȏ����?�W�׬lG��q5��Ɉ#YI��8����A��� ���v���wy!����r3�׈P�
��H�6�΍�-r$�E�����5���5�$:^�o�p37����OB&Up� �kU]�㭿����Vj��e�&Xzآq��Sv�b�9A��듿'>�KY�e�GI��ɰ�ފB�H����1{AUj�)���,z��bĎ�n��a ���M�����#Bg�XlxVHYEB     2ed     130 �G���Ho�r���P�2���Cf��6����ǡ�*�t��,Flz k#`3Y�=�=h�]Nԯ%e�2=��l�{G"���i�O���O����e�c�%;|�,�
Ь6~�9}��ROO�m;�c��ຩtg��@�ι--"豫uز��[��	��1�^
��bnil�>Π@�b���A�pce4{2E���"f�z'��5�U�0£�����Ϊ624�W��?�|d
H'� �����ys�u�ǀ�Ia7b@9�F�w�ύxWә�v̤�[v`�?�q��=�?�'Q��lv�Z�tU���wF��