XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Sr}�)����2�՗���#� ,?��
���e��$�2��0�^(�\�|���ODɥI2�g0�[��^8VY�ԧa0��b8�d~EH'\ �q0+��yیɁ���bv��6A����Po���~�&�Qd�iM��HP����h���Őb�����%g�=��`�0� ;�4�,�����Y�IS��	2p!�j���PO������Ni�����&��R��ቼog5\�:���N�}��",�{P{��/�-Qq�~]��B��xvk��O��XfC+
���_M�~ *ry������0�ߎ="��*��ݏ�+Z���~��JF`��=%s�i��F1�\I��+��{��W�q&��e��U�� �<����6��H�Հ�PF �p�8X�UL?���UЙ+&jS�ח�hm	t�eQ��La��͘�D���m�$��
��&(����I�F�RƁ]@�v�$�"|��J��A�d~�� ޱ$��F�윃�E�/Ru��tj����vڄ �?e��ʷ����`��Tx)tK?Ws,��$|m��KO	�\��⹨�j���ώ~Zh��m�f��/uYB��4��)m��(�5��/Ed��x���F7��|=�ux<�<g���(������D�pRRa�\�#�&|���`7���4�&����܂�e��Y�q��Xh�Q~�p|�2y� ����9'�,��M9������`�[;��(G��b��X�D�~=��g�T����#\-�QZXlxVHYEB     400     1e0ͦԓe����&��6�L+�.��y���fd���(s���?�C3����+�4NRg��rL��1t�/=�P����U�������c}zAN�؊<����b�s�*O�t�3T=;h�kP}f:E���jh�t�7�>M�3ۯZuy,0���F8w({Щ�`"Kd�Nf��~�
:d�PC�3���QN ~��Qz��_b`c�~1	O�I��"�]}�<��mhJ3�䨫;o*;�Rq.@�#��xfB�xxfE#�p�^>"N��(�`��3X��C�5*�������כH���\���J�fƙ�3߷��P��s�_�N��7�%O�����b�	�*��7��P65��(f��27��L���)o2~&�cep��M�V��i5c�I�j��+���2J^;�-��8Q��ǭ�h0���
|�(�:1A"R�!�w�����-�]e��Ǫ��,�։{�Ȏ�z�˸�E��FK4VXlxVHYEB     400     1306R����������m��D���*b��t"H�����'/>��>BAl�Q> ���)�x��ת�]���M)�;l`���<�+]S:��:_
 ���o��*��o>���P9��1eGKi�È�L<R["?����	ku*�P��Y�2Vָ̂A�)�,zØ��X~��	Yp(���ZI�JFK�3dNRq�!��ɭ'��Ƃrw,�z��[W���b���so�le���I�'��bn�̋Vד��"�cІ�R_�$'+e���r)+:�����	 OxE#L�F��L�FXlxVHYEB     400      e0�˱n���4ܫZ��s�(�
��l���Gޫ&�'�`\"K/�+C�F���Oxc��Ըk��;��~0w���T�|.Ǔ�r��t�v�5a�����oC�E��0ʴ{����"�R�"|$�6�*���ΐ4��x����/�,FSlW����%��A%�?�T8*�lP��<&��u\��%#L4T�v�q k6��UxE��C����Zz��R���?[�XlxVHYEB     400      e0t�U;�`d0p9'�qR�}���/��O�D�^JT�B���$�
��H�L�h�65O>&f��ˬ��E����q�=X��MXtg� sw-=x�w���B�3Y�E;D�uTW�1�����T��j����m��ƿ��U'�)�w�9�6��ִ��`��o?l�~ᲷL<Q��ۗ�t�S|��P��ѧ�xu�ӪS��#E`}��!��t�D3MG������)�Y0��"��sXlxVHYEB     400      e0^���eQ��g`�)˼�y�gh�l���hv�|l4�'������D~�`?*�����������ᗃ�n~���d�ǟ�~�ݺcỰ�B�4r"L�ѺCщϽ��C�B��>��k)�Y��|�����jAJ�;a�o�1������ *@|�0���U+�D���)� �?O�I:V��!�
���O�R���/�!�)CPj�\��|����нz�Mʼ�9XlxVHYEB     400      e0+@��	��6�L�	hM(}Oo`oZ����$3� Ղ
�����7j�Re�6�§�%�N �D)8F��ft��[�����Ou�]�*uvq_�x�oW±{`q�|��Y�(e����p����˛x����fM"㧪��Q��ƥ)jMB�ې�����7��yAY�����)���m�L��I��(��c�㽔
z}��<��B�Szvb��d���/���X�<P�XlxVHYEB     400      e0�#aޙ��<�)�I�_I�`j�>C������l}ܻҟ���6sO�o\��2�Z2���B�(xN�#����F��$ȶك��x��0����EN�!n�K,x5K��8.1!�<X���C��7�X���m�4�n���a`�i0���2����/����{�=<�?���q���8���N~����#{�:�`'��4��WK������	eGmC�<�f
�`���MXlxVHYEB     400      e0;	�Y!RY靵�j_���K�I����	�r�s�� p��,���Gpd��Ւ�AU���N�x%Z�1p		*)Q���mRS\I�D�L�����KPg�C_S�N=�(+� pH�b��ş��d�oa���moY�yɗ-ݤS�K��g��̛�w$�4|/��J�^�� p�p,S����s�Q�������pѫ�aV?*�f�l�p*�ֹL�GƤg��zh@���XlxVHYEB     400     1a0oД4����ؾ�?[��@]u��/���q%��vL��TP�̝8����
�YS���約�=��"�!G8ߎ ���36E�i2�*�+"A^�g_�5�za�"U/�Q��d�@���U� P���E��(�������˥X ���V(��ؒ��
�Y�̄N[E�]�):���j�N�[��}v� ��	E�`�gw��bUwz�<&�4�k�[SQ<K_e7�6�]�s1+x>,77'��L���.��T�f��W��_��&����s���K���,����Wi�z�Vy<�p�l��j��b-�B* ��H��u�Rڔ>���\�2��jB�qaF:��vG4��n3D�o@ԘHp�ء�
ud�,����oc���I�U!�W>���AooDM�n	B�:�4�j,g%��JXlxVHYEB     400     110P�t���D"R�dp��F�%5GXmߩ8u`	��$���B�D+��.>�H�r�p�q#�,V��] `�rװ��U}m���|�D���E"X��N�c)+l���qh6���3�p>T�/<6�3���`���h�ZkJ�!�4�yP_2��dx�/SF��~,ʳW-���Ezx�JC��m�հ���4�T�(����v��vM�&��s}�w��"-��Y�=7w*f�8�a��Lt���;�]r�Ѥ(��6 ޹�a��!�w![�]�)6�XlxVHYEB     400     180k'�Bw���D�p�ou��C��y �����7�i�Mi,9�_��
,C��x:I�,�EW6��K����M�S���2J�vQm�
~*�yj{�܀��;w}o�����+�*I>��@|��c���3e�*�|�WR�R��2��C�V�}�6<\n���ڈ#-X�Js�D�	�~)�;�Z�6�l/^��g�R�����nͿ��f�z��0����(�DF�v�Sx���F_td�.D���ѯ`r���F \�����i�!�bal9��N����lѱ]EK:�#���w�d/�i83o7}�t)�����9�r#31>���sV�Q�L�X�@8����N�=�c��G�����:��I5?�EM�D)���	%�S&XlxVHYEB     400     120.}�-z��0�2�2�'�y@n���,��3%֤.�" ^�0��P��!!�z��7���ƅ�A��Ô����\����)��R��ܲ��* ��P0����6!�h�M�jŪ'���Q�*�I���C�t��z��,���:�I0K�X2M�ғ���}[/�ɼ4|M�����a�c8B W9��\�L�IJ�����`��jY�(0^��}������]�?��ɠ��:M@�]{��V!����{lÎ~ODb�[�������ݖ�K����X�ld`����3"7�VXlxVHYEB     400     130�S>�K����_m�3'�ď�P�M���Ւ� �X*!�g���ӰI�f;}�v���)�4�4�`�&���i�A����!/_���!�;8(LՑ����SBIF�K$os e|�v�(�Kb�o����
���b�a7R
�]s��Lك.��P����ﾜ�l�)^8VU�Y�{d�w�~�!���᭒$���N�N���H�#�v0O�Ar��'�z]�&�ĐG�e������a��Ժ{�h�eE`GR��	���B[���_�h��D^��嵧|�E!�����e�Tx�ݕ�\X�a�XlxVHYEB     400     120�k�_�^�W��ao��x�U���rG�����$Y���v���:0�wE�3r����YG�\1�[�ܸ+������\�e,�6�Γ�78b��v�\4�h�^��1���l���
�\�L�
C.�U�ϫ3���ɰ��@띻�1|jg�M�7����V
��-_�o>�V �A�t�T��X24�-��k-�vz�/'Sk��uP��7���:p�ܣ
2��a�!�d(pm�6l��;o,<��f�Z;bg\F�Y�n��W�X�q��a�v�a���M\�XlxVHYEB     400     140��o�3iD&el�'����z󮰱�Z|�=�Y%��Ot�~7 	��H~�;$v=��4�i��ChXT��x�/7$3h���>mrl������Ȣ�$H^A�34%�.`��<��Q�������T�0�>x�M������k<̲�*w�`B7{A��¼`m�x٩�y�_-n��&!���6�AϹ�#��E=ڃ����/a����is����+)��7&���(��;g Q�5tg��hS7B��Vb��:x+Q��s!��c�EJ]�xAsQ^w#���^>�I$*�=�x2KB.���7���q�j[<T�(��t�B�eXlxVHYEB     400     140����W��H
lI ���ԥ�#�}��!Y}@C���;��>����������β��DB�yw]z�E�[�s����~�j�������F�>z�4�؏�� oL�5��qZ0�B��ѧAy
�����W욂���fdg�Q�d\
��f}5	�f���v��1��z-C"����`�k;�d�����އ ����j��R޺.���NU����MD0��18=����DD�h�l�ȃ��xyK��3J��W��`��'��[����L�H	P�-�e�B�9#�Lq���V;t����ye�r4�wMa��JM��x̬k�>�x�gXlxVHYEB     400     120&y=�d��Q1�	�0;�2��Ȭ��D�2��(-5���l)$���g���1�M�S-�(-�;ԣ��n�	)	�u^�w��[Ev�q�.7��������"�St��%~'��l�ac�T�#�k7��{����3�A��h�*ѩ����EV���Z2J�9�K�5�K��������j1.��e�2��h��������(�o�7����)��b����Ui �w,�D���^��o�ŧ��⩢1�8�!˥�nn����`�<�{��~���G}���Y�dkk�B�mXlxVHYEB     400     140�y��a3Ū��<t�^�hd���Q��X��D?Ψ3��	�<���ٝ?���,:Ф;�`��x��^�4sF��:z8�Q"����Ša�G��b���e)���E��=�LJ���)�u*Tћ��I�{U����H>���9�-a7w1Ƌl��V�E��{�ӄ �1
��H��uL�'O�p9�5Q��]sJ����ag�����)<��_��)��]�RoZ����Rw���s�j=I)�<C�EL�p��2m�6#�Q������R�Z���(#��c֡u��p/��3�(�1���PL�uz�Vf��j�c)��)u��I��XlxVHYEB     400     120���e�.��
����2�T�+�R�]� �G�D�0b��11L�+��
Nf�4�˟�����*�a �o��7#�	|l�o����Pb`'h�ߒ��1	y������F����	���� N�AG�Օ�w��� *�Q��)l�;����H��ol�`?�c��Dw{[�}jT���Ӥ����g�������N]Y0�����Z��?۲��dw˪��7��nr���~S63R��v�������n���:�豧z=%%]���hT �q�8d�&*b	�N�6_�D�O�%e#��XlxVHYEB     400     130_�����a>�Z���>W0��7J$��bz�1��W�-hS�����l����1L����p�=k\��aj��s��9y�����bshǘ����*:Eگ�)`]tWp7�Y�!�D�]�ԭV)A�iμc�������]?�U�Ѷ@�p��"�d�'�G����4�3����Gg��o�(��qt��S�Rit���D˧�v��C���%�0�F�M�8��b�����~��T�	�v�GG���w��/g	"����%�$��BK���d]w����7�)��+�5t���+@+�̕����XlxVHYEB     400     120f�ml�8��_Q��/w��9�O b�Xtw�[�isA�UV�طc���E�R�ɰ�ɚB,л�U	�~��]Œ
 �MQ�I�^fs(N5��m%��bb�-�~���G�~]tl�;����c�
R3u��~*s8��>��Tp;?F(ؿU��@u˦��I	��ۓ��mQ=bY����W9[Y���7����"��{�l�u�oQ� S����>�K?��Um-�boΏ�瀘�����=0��L���p^۽�s%��L1���5����jLOoYXlxVHYEB     400     140���d4�e�s%�hv=d��RД"|D���$����/��`�*�P9E��Ozzf�M�W�*G���!\�$%�ı��V`��ˍ�o��"����s.M%�O<�X%<����NQ!�SS�hz����$��Ă*���n(���0R"��OZ� ?cL��VS�}>X��X�X
$����a��m��-I�����|�P�"��} [��|S+��&���%@�0���Dr���0�,*�93�����(:�N�̒�������t��q?lyi���]�[3��o��ф���"H�����{a�K`c�u�8ἲ��vL=XlxVHYEB     400     140����W��H
lI ���wYL)��C�jp�߆�LBVQ�Lp���,Zw,�m��Q���Қo�����+N.�mx���	��6Z�P+XՠJG��q]h��> %��-��.�2�&�����|��o�kG�����f��L�w�-�'5=��&�ٙ(#� ��_Ť�za8
ƺ�L�ZL4��P1�[�Ÿ���x�	PCIf+��M�-�q#h���7l�<�;
� �z���o�ݡ��_S@��tv��������Ҍ�������}���z�6��Ͻ�[S��\�$T�×�������ƴ#�d�<(�'XlxVHYEB     400     120۱�4�j������X[�a�RJ�����b���Fx^yU\|�)}1z��E��/mbu����#�j,��W��Z��B��q	�]Q/��w�^��F�H���~�
~��a*��?���Y07�� ���db�&5�̾~����{�>H�X�M��(C�A�RD0�!��,Ojx�&Y`L�@�Q�tTky]�\w�B�t�[.�QtV7��L>��=�a�B3a�T�K{g�)ujh�������F�g2��:��^j*��*�~�PL��m�����-�`6ժ�XlxVHYEB     400     140�c�F;2zV�S�~�i�!��
��Ay�?�|�݀y0�7�����Bf����)ۜ��k�I����0�,�1;-reI�v\��O�X�;�.��M����f�C�^"武�m���!ύ��K��r����2%<k��&m2�"���R�R�ɩ��N� �J��(-�(���m��D�}�֎\1a,����]'�c�n6���U2����������9-
	��VE�ӎ��*��U�J@3"eXy8`�_)J�=O^��v��Oɚ��K���kЀ$F��d38��@�_�8���u�� qR����j��"X�XlxVHYEB     400     120���e�.��
����2�T6�=�����q|,)tv�̤��Oi$Ѝ���VWi�܊�Yzե�n�U�i��E�Nti�2��`�.5��J���ف�S:� ���h�����UpGk����3�����P���T��X�P]�!������R.	ŨN�p��By&b�E�X{vЕc�]#��
)�6�8����5���h�ʛ���p^#@�m��N�Rܿ!�-��)��s�8V_i>�0� V[���Dī�C3�TIWbz6 P0��u։cF��M=���ɏ��XlxVHYEB     400     130���l�dӏ����>���|��'V��?䃊����{�ՠ��	�����YB�j���S?O��$0�ʀXet�F��S���g��^D���+f�[�<��2h�`��ε���`�	4F��	y����/�� �h��kh�ѳ�-o�\@�8Q_����FL_���L����0%rM�x������Itzeû$j&G��c�օl��S�I����g!Z����^�g�큹+;J�4����A����^��o"ږ~t�q��L�~L�
p��_%\�=��X�����?�i���J�����-��������q-GXlxVHYEB     400     130怰�A2�H`܆,��$�)��"o�Ӻ��}Ls��ǰ:����Q�Xh��r�wd��'���R\I�����`��~����40�>�13�K������P�Eά����"��>�:#Z���Ϛ�3,�.�qn������w�#���hJeS��z*����ʻ#���0*�q:t8����n.��.�e�ڵ����E����F����J�Ie�<P+�ܣñ0���ٵ,��8O�_I\�g&Κ�7�-a�3[��U����C���:1-����o��!�iG`�5���v�m%�Qx��ڦ�XlxVHYEB     400     140��U�`y���{"�����5'r� q�,f�s����}S�A�����Q�'�׾�����B>$���Nl�);�xv��=򃋄3`�t��(J�]CoŢ�w!�~{�G�a�#�m_bX+v�ڈ��(��=��L� 6[h�i?s���\�K����x���⺺�)��^�ׂpײ�8����V$�PӖ��)2�Яl,��P�;N�~�?|�&/�A�;mر�*6�?���Y��,�Ή�vW�
ᨸ��X��62�����퇸��}Y���4(��75�i�S�V�k&W� u��c��	O� ߕ��O")O���~\XlxVHYEB     400     150����W��H
lI ���o"V�g�C���uS�GR�F��92]a�m�	ԞD�W�_�ލ������C<�;�}.̲.��r�T^x���xֻ����nV,Iq9Y�N�[8��!#H��h�lnD�ú��-�Tn�~����-����+�B^�<u���O����<[� u�Aq`����>��=E�8ЌT] 9�N6�OII)k躟���aF���C 
Q.���o0��ђ�;����a��������8k�Q`sB.,�b�y4S}Gú#agGV���K�5��	̢A�LNM� ׏�0�+�4DV@F��9�LB�P�AP��fG�W.")q�kT���XlxVHYEB     400     120�w8��dvJJ<Z�D�(�ɲ�!H�{r춥T�0�g�s5k��D�mbW�H�J�Y����-����e��oZ*���Yݨ��r��:
H�2N�E}����tK��U�ϛ��b�at���~9�@�J�?YM�Q�*QE]߈�� a�M�;aθiG��F�|��dK0�N"��|~�c�c_Z�C9�,@�
�Fg��9������Q6 �t#=ߠHX )�ƌʒ�m�Y7�"
�J�8��=?K�U����� )e�>M��6�N�'�q��J9D��F%�+��4��P��g/XlxVHYEB     400     140�!�$;�Bi���A>_hn���	ܛ�}�^i�.��Sިz�Mf�h�EB,
���?//��n�y���˺�uOK�!���x^�eM(WWP�@k��C�`g����X��Z��bS.�_�R��{�"V��K��g�lw�"T�3���h��^(�����j��f4z
��s��e�eȭ��M����B��&yE��K?���i�n�D��W�ȉĲ80g�����{�Nn��޹Q12{	BX]˯G�梡�t9���ϔٟKE�0-�����1O=-tYb�PљU���kNS}��o�o߲�e5��fl` �9�~_ro?�XlxVHYEB     400     120%�ȗU�s5��P���*�X��H{��"�	3��IP������Aw��^T�.�Yo(��W���A��t)�-�&,���$�JBcMߏ���`Hy_�q��X ���)��%��̄(O[oRn��i�KVjȀ#ͲW�16�F�����Wv�Y���9c�?Y������ۨ�	,:�W���J}&�V�ȏX;�l�����;3.<��4�{��K�j���N�!ȓF�ɖ6o}4a�T��gV�?,ݝx�K�n��W0l�UcJ�#���p�)�o�lXlxVHYEB     400     130_�����a>�Z�����΢�柂�e[�\M]lu� $��!�2��}�1i|�OF�Lx4]����Q(�/�7m���7e����PշQ�Úzݛն���;��� ��Q�cmG���7q�*��.���(��d�H��'�n��a8�`���RԖ̶�`Z��wK�p�qnv��O8�G�����O8_��Z�LI�+��Eb�:��n�� <r��`�*�����X��Z�0S����`s�ʈX����[����\�R#{ck�͗3�}�'#��Dާs����@�:��XlxVHYEB     400     130怰�A2�H`܆,��$����b���S����n�2��9��N ��������	�W*�L��c����`�4d=��@�Ǔ1/�(i��ܒ� �Td���*)E�Z$A�Ֆ|!ޯ����e�g���`'܊�m�2˃GvzC��+/���۹Ք	څ�Qh�Lj��~�A�J�q��L1�U�Y������
U��s:��FV����-�O��Md�E��>��0P'j����8���P}>H8�PFT�
~�h���7��M���F�%A��W��i�.����HrZ�!�3�r��S�|�r�)�FC�XlxVHYEB     400     140��E�6ܪf�Թ6Dc~��1:,ᝏ=D�ɔ(��Tzx06�ơ%K
��l���n�Y��*��)��j��F���x�G�7����u�0�Ӱ�7���Ė#�>��wV�ɡ3Il���0�ca���ɢJ��D�H�cYD��r�ѕ��3#��]?Z�N�X�U��4��^���\�P�oD�F����,�V��^}iV��n�KZY=,��Y�����L5M�~D��xG�q�H�da�{_+B�I"�Vk�K9`c[T��jy�)��%��p��3�
�����j�֣GA�S/��( �S�=�Fr�"d"jی�XlxVHYEB     400     150����W��H
lI ���Z-��Z��tm�(݅3��Ѷ��	���o8���+�=�����'rz<I8⪖#t�|�l��z�&�����FF��Iꏰ4"�<��0W�b]�خ")u���{�`z|��?`l�C:y�\���2�?|xǍ���b���w�¯�#м�I�泃������6p$��*xܟ| ?̷Xz��X)��/05Qfp"P�Q�� ^���� t��1�\9H��g��M~�����G.o����@�K��0OUd���σ?��
�YWd�;�����^�0T��ˊ�k{h%��wv�bx���;�hR�XlxVHYEB     400     110�OTC�L�~mֹ��ԴO�5#0U%�l��SI��N�� ��`�D��1:BHxz�x�n���ܻ)�_�	��M���+R�7���������Dd����Ecz�<��#p��"�,����2y�$x�F��0������"�U��%�iUN�ed3�M�'-��%~ѳ:.?+�N�������H���������fF�Bd��O?%��V���6����I'�n��}	,4�Ԥ,���PZ�Q��0V��̃ǒ��:�M���q�XlxVHYEB     400     140eEY�d����dH
�����p&f�l�9�p�Ɇ%xƁ�Y̎|��ڰ�&��pt�aQۺי-��
�0��vW�D�_�[|���5C���69�[�3t_r�?���0��wh���X�Xzf_$ԵD;Te��]�ɢUTc�_��+�h�-�4�ܹW (���0�O)4����k"�E�	�:+��UQ�\U+*�wD�z$����_���d-�6WI[��M��4��@��ι����"z6'��>�5�j����N�Ɂ��,뿇{��[�)S���Y�3uȜQ+�ࡷ�;F���WsXlxVHYEB     400     120���e�.��
����2�TO�Ve�L#��.�޶�f������6Y�)�9\_�D;��7ׁ&���㧌,+�}��$V��y��Ӥ�3�5?��?���!�I ��	�D_�;u�$wKj�f���i�T8��|G'vU6q�1F0!��y56�΢/6�V��?b���̢Ю���I,�]1��`kbH�'�t��<���"�����v(T�3g$��b2S}�?tGp��͆���6��-_)�(ޠiT�ԍ��iE+���Z���Dgj%Q!�`(iux1��bk�Л���XlxVHYEB     400     130�o�Ǜ�P�'��E;��D.!�F���ߌl^w#z��*A�_�j�7a���XG�c�҈/���Nܲ���5��
o�d��?>��A$2z2�\���Wq�#�#U��/!�\�������Y.I�����>����A��T�������)
pK��(�P�m(i�{�W���n�	DЫ�b`���:���q�hT�����������b�Ĉi4aw�7��E��5������B=���2��c��?Q	)����k��6u��W�<Q��di��"�������l�w�"��-�Y��O�d1"�oXlxVHYEB     400     130����@���n�T��^�i1h-ﲜ�����`�n7ݼ��p��z��r�����ǲ�,8f	ܦ��k;��qԡ��귘�-g���������s"�u�LM�"�U"@>�V��=�~�$(��2?,�����;�pf���#��?�_Ϩ��� )�g�JvG�'�sތ��&�<zs �_�m8W}{}4��@
%�����5`Pڼ1�fB�B^���Q9���s5}e�����i��nn�����t��w�
��&IXx�T^�ZaV��u��_�{����\�L�7N,L`XlxVHYEB     400     140��,�UK3�������Ϥ��.�I&*J��9�y��c�#)�W���C�߹��M_J��#�3��u�8ݫd��ERb�gb���V8?�2?�>�6N����6q��V3ʿ.7��
-A#��cdH�� :�F$J�B�<5�M׶��`�d�dK����(�4�CN��ƈ�k�}1�2X[�����p���_��P@I�,�8�P�ߢ�X���Z��T�#���T�Bڨ?����ذ�rO-�&���O����l�:���6�Ӯu�"_
�tXb]�u?�Q���+�3���?�f̗�{�����Ufg�;�����&�k	��XlxVHYEB     400     160W�P_��������{ǁ�@a��3*�����G�%:p�`�����a2X����(k	����v��`ݰE�>1�Gɕ]������'U	�(��b�mT���,.�����$�M��j}�g�0,�Wr����v�ӚX&��D���9A��/����c��$�� ���xʕv�o�,�p�c�Q8ݐ=�)�
*n�?�CkY~a��$_����p�c��J����l���K9G��a��"nel�ʔ�oeh��T�_ �n�p�p�0$����LaE����<�B7�mj�3#���&!��-�;�3�bX��g�7]�dkN9Nr�S�3��3ʽ&Ww�8,���6�C�vXlxVHYEB     400     100E{ɎlSǜV����`=�o��������lbF�t0;����R�܃���3@���o�D���CT����vD	`���p:bM��t��������d�tZ�#1��=m>�4�bI�-��9.�`�X�]0	�0������>��n�����_c���(q;w'��|,��(p�M��
=2Ł���[5l������[��(/)ܚ��2�B�j[ ��t�u�mr1N�l�9g�H�u�	ŘM�'���ސ�XlxVHYEB     400     150XL̼G�*{ah���{�]�|�.bqP܂�M颍�ں��P�#Z̲�f�^Ԡ?�����/�b��a���z
�Ax��E�t.�'�g>�o}�<����s��۞/;F��D���#�iކ&P�`�U�`n�c��^��~ ���g������ذ�;����O'ߒ�Q�hm��.-+WTsMM�����·� 嗚a��>/;%m��P�� v�(�.�Wx��\[� ���NA7y��B(U��64�����5�e�eոm *e�'��;0�0��h�t��	e:D��ܞ��Y�I�*{G.�{a���F��Mj�nˣ��.���T{���!vXlxVHYEB     400     120�Q߅m&�%��7�.τ��_��1�1�ti����h��`��K�?᎐�\�#l U`3%�6!(��%�3Ǟ�j�������CJ��/�u��9R��WWǊ�z[=�rӟ`-��ҁ�힅l��eaI�q�k�D��m�v�g�Τ@wH/>���:�>��N��8B�C�P��\V�5�.�_�zڪ�O��;;�&��d�?�j�"kԹ|i������C�81��'�ߧf��J�A}�{9�,`?��,ܧ{Z6�o5l�W�1�WT&�j���C��c���&DhR�h����$�Y��XlxVHYEB     400     130���yK�۳%~��y!�1�ۄ�X����G�6o�ӡi��o�qvX&x���Nʚ�jhB1F���|
���y���ݤ�~B�(՛�|-��Q\�q���ֺ�,o;:I�~}�ע����~
~����fQJ��{/�.ڏk��.}�n�O3v%l%��͋�p_0����eRE�����w^��e�3�gHx]��l�שڮ�Rb2o� 4��q?�1Gjb�_�T�z�I����T���� Z�=�q6<��$���@�&�Y���j&�W��B��% G��F�z��XlxVHYEB     400     120�ܥ/� ��ɡL������6ʀ����#lv��'NZ2zn�'toΒ�ל����J�����-����ͻJF�v��@Y�\����9o�p�)S�6wq۟�J�Q.-Я|@�p��s�P�Ui`�N�N2�,kHR*�@�� j՝.\d��.!�o��ހ�_y?4���	F�2��ӵ��t���d��!Y���v���zq1�dR�5Z�V���.�)S���RH}�pp	���S�4c�0iDU��g��7�d�F���h�ѲJ�!�u��aӏA�XlxVHYEB     400     140���a�N�i/��Ǣ�o+i�z.�L@���x��?@A���v�ʏ|����Mȟ����:�B�%��'�����=8�����V�2�m�G��r֨�%>?sB�~�8��@�� �G�P�侌@�@`,��;�̇�����`zƁI����C	��Fd����B��e)b~��F�f�9VE�kH	�uB<A-+�=`�x@{�]�R�d��n�Q&{�Gt�B�y��w���BƁ)ĬCL<(��_q�<�	D}�`�M;�W�X&8�d�ع�8�y����������e���������~�A#�w��ar��3O!XlxVHYEB     400     140PW������?_vG�ꯔ����_-��|� 6��Aվ/6�]	P�v��MJYv�a���GTJ,��f�~$�����^u	!]�}iSp�p�\b�8���r��$�NCEX�d ߁�VJ�>���U�*v���ֹ,����h�=`�&�@�P�������@����0O������0I[(���艍���w.��H�ɛ7�m�z)B<]<�	Nv���n���[�|�<��g�> ^�q�R�j?7��ҍ�0E:������X7͵�=܂$e���!��in�Æ���ӣ�ҡ}�>$"�9ϼ�5�k�|HXlxVHYEB     400     1203���-)ͨS�;	Q�N��J�P=����D'�\��� Y]f����x�4SI�D��eGh�6���qc�v��ΰ����z����~���T���_ �f�Wg90x�Ľ�Ҥ�6̧_�`<��UnR5B�R� ȝ'���_h;E���c@��n��oؒc�vs��p2O���.z�8����g�	=�d����Zu0�n����U���,�#�٠���#�z/ۡ��L���/���z��� P\3�PΈ��6��'�Ŝ����>{�X�uy�CsXlxVHYEB     400     140� ���N�2z��8w��
���C�Z�+gtS�~�/�||�Iu,/0��P.����	N�X"}���=;-�2Z��� �O4�J��A�9���SHC:x�=*���=��i�{���~kMuO�2sP�<~sEa`Z����S����'���V?ͤ�7�b��u���	Yy���+�[��<��!���*�,@7��eG���&�O=��3�R�پCN]u㤶{�������S�&���N�vK�����v&�_`�S4j��K髶|Ɯ,�Tű�tR2��e��1<:d��_h�Z
�hd���P�QUoh���XlxVHYEB     400     130�*�/C*�73$���B�>�9=�iP�H�G��psh�d޴�J��>�ϗ��i�T�c��K�k�t�,q�Loz���KÀ����6�dw�mE���2����_v��}��Q��7�C���G2Z�:XO�J�a�<-vۏ�sry-�v�ԲVb�[hU*<f`�-�*�� ׄ8�k�#٫���u����]�#�pD�1�+�.�{��{�}ёZr������ip���5G��P$��K����2탇H����>���ȵ�3ûO'Q�� ���������\s�Vs��i�p{��K��y���ٹ�Q��XlxVHYEB     400     160��w��\@,%�뢕b���ǅ�)�2=��Ą�����HO��@��ԣ��MC!W�Q�;s��m�!;���JXA�M�Ya�����;S��촎E�GI��\OV�Y1�5"�P�f3%;�[�.�
�:�o�ZˤI��t]��a*3�=���^�X��>?��P�N���=��Z� ��!ߑ@��������nPON"�B�*��OG���c�C�w�?[Sb�R�<m~1��ȂP�ևɠ8{-�+�Z��f��#�^��V��_Fk�ţ��b������<�2��=��h&��g��_��>��o�oA�s��)�r1	��0~�B��00Mg���S`{5XlxVHYEB     400      e0�H���6�������vО���M�2!���X��~�N�*<�VU[\#����i��KɓXX�$�jVI�J���$g,(ٛ�2����v����C���7��ܦyOT�K�1'��X<��q~缷ow��@��X{�@��.�����:���T�x�K+|��p��B���C���H�����l��#��|i-}��|6?�
�t/G�0�*� �2ͱ�~��3JUXlxVHYEB     400     150M��Z�sne�mM�h�d�j���&UvdzV����d������"}����":5��7���$��h�3�2�#爀�$�1�ܻ��pff���R����_��\F�_�.E�"���a�_fLʶ�עLBo�	e b�������B0�p�Cߴ��4�[Z�ɕ�+ۏ��L$�� g���)_�����O��+
��(��L�):X�#����z�֑�>�,.��r�!��R��=an�ɫRc~���F�n�C��g��ְɘv��'zpr��@��� 	g߭WQ�/D��߷.�E�t�?OfR[�.� K�֝�-��ŷ�� U�9XlxVHYEB     400     160l�?'EY����2�(#�H���)�ST����;�k�.YL����D^)�B=�#r�������Sw��s���qV��ޗd�
�
[k#�C��::?m��=����G�t-+�F����8�M�n�uS�ƚ{���MTمޯ}�"wN�)�(���0��ݴ'2�)Y�GO=�g�ȝ|?f�� �X�F5�}�w
4�I����Ao��i��gf����)iK�cW.���[��X���=�W~ZƄ}|����mBMĄz(z��m�0��&��cj$J2�r,��=o�F<dR>)XC<B��x*"*<�D�L�dX��ւp�O��W�ؑ�/��'��p���XlxVHYEB     400     1203���-)ͨS�;	Q� 8.������> �����h����' 
v������g&8s�� 
��C��S�f�K��_P�xs F�,�w�x�
�Nס����g+��@F��:��Y�3�m	��?/�@�N"V�z4�$��a�n �N�!���#�j�8����"����N���g����t�14�ĝt�L����ơ�;h�O���\R̹��͜
����x�>�K��%D��c� 2돝�1!��}V=���ցRY�39���W����Us-I`%A�
XlxVHYEB     400     130�//�n�#�kl� 8���1҈g�9p�cM�LZ�;���\.k29����#pV֬�n;�f{��$BF^���j�Ls/��W��VV��ڳ!��B���� �/"Q��r�.Oʑ��H��!�P(4��"`�%�"�{���9�ѤK������"��g���4~;��?��AǰV	��#þt�sW�	j:�muh��قU�f�3����~�/E�Pm����1EwNѲ Tcйqƫs�U�Xj(A�S{cq��'�ub�X&4~� �w�p�w���J���e�ٿ��XlxVHYEB     400     140��2+T��OD�q\��Mov��\�r��=H�8
Y�x�љ_!
�^�%���b@�kJ�e*���3�B�ܫx*(��>Ӧ����?s�Q	�Od�4)ܗ!�"l�o����+:�6�=Ԑ�k+3C?]]CP<.!���}y��(��ݱ�|��UYF��h:F}ބ�k���GJ�� ��i��S��]J�дF:�S�3�Q���ꂙ�S�8GPj̝����NK��PGkv������Y�V��gcX�f~�?�P��l`�tx_!�p4A��sx�Lp�Y�5�KxY���ɟ�arڑ��a���t��E�CXlxVHYEB     400     160�4Ba�'�Z��P��B^�|�z�6yp��t����oZ��\�t��[��&K���Q݋���
�|bl>|���-�+ߧ����檺���f�Z����$���v������`�\I?,�S�&�1���	E K�E7��]#�M�-�۝��
�rؾv�n&��C6%����Y�-F Lo�4?����ӻ�x@D��J�!�݂[���� T}|��#���k�[�v�v:��;� ��~;����Q�����됈$�w�J&�XB���v��XTM�/��1":0�8;�'�U%y��B�,s��/<�>��B�U�B�kd*ff�ek�&��0��ʘVVXlxVHYEB     400      e0�]�߻��	?	3�G4�r�{�����~��w�9p�v
�O�� ��N��0�t�)T��CY��,d
����F/vh�s �V�o+����Q��d����{�)���h�$�Q�0ў�-��z'�u�etk܏c{n�bXy?B�љ t�d�]'��9�7��P`(j܋p�����n��U2L��R�����k��]F��$��п�nm tI��o���k�XlxVHYEB     400     170�O�F
��|��	���v�F��j�v�t�k�8��
�*uP	ݖ=Y�ۃD�g�O�OH�����ݱb�p�kA��^?k��މ�Cs�s�#ko�&[ 4"�T����8i�}�T�Nkqh�S� g=��sW���H}(�ޞ��[�q��b���g��aH�
�I?Q��S��
�sCC� ?5���}���T�RXW�]��pX���@�6��&����aֶhZl�؉�?��:ɴ�>O_�������^ϥ�=j;n���z�Ws� �ׅ�b�$ث�O����c��0����PEȖ�k �9u.�m�Øϻ��K5����2������²�i����}���9T���Y��1H�XlxVHYEB     400     150&���� ���d�X7�B7h%7���H��[e��~��a�r2�b�,y�p�9 �@+�$��溕z9q�&���Y��J����v#](���X܌���Br踃7up���i;� oK�v�f��f�#����c!��ǈ��;o(SA�)�5,��y/u���\���?'Ys��k��eGe�"��<�o�\1��tBM��䯞�7i����Y��^��Ͼ��D �Z�L�=�J#8��x��ow��0�Enl��5(�*�l�������*%����M\�ڣ7�� 9s��S��O�w&t��[�A�\ p��Bl�\�XlxVHYEB     400     130��l�ZIO�H�Fv�0V�tk�:�Z���,a��ל��~�ِ��`�ԝ�^���~K�r�Fd���I�l�W�7v�ɻ�=��H��R-�k&j�2�N)E ^&4j �N��&�5�AO������(ZA2&�*-C>�%��_��P���G��ёbF��1�^��Q�fm��s�����F�Ү���3�����u<Sz{.'�eZqY1\n \�u��x�i���MC�p�%d~
#�frQ��$�w�C�wv[TCKsh	�1�y!>X�{�1G(t���������t�>qo&�*w���XlxVHYEB     400     130��Q~��셤�xTm[�g+������%`d&�'[�	S��>��N�ق�D��/}��l�;�ǣ��ؕ3�n+$=ߕ��>.嶌�aO�[��H�H$�=$�Z0ա� �Ճ�p�1�G0�T��*Ʃ�����knj��ѝ�U��>+������f�t@Y�NY��;��2��QgU9�.�����c����)X*�N�G�7�"V��"��A����UK�D�1d"���<3b?2=V�٬��X6/5`��dwH1���/ឡMR���	���¸��ߗx2G��QK)��+�5��|��XlxVHYEB     1b3      e0���}�j���!ӳ��zϿ���ºq��g�T�pw��4Te�e�����x�)���Y�Γ�����|@��b����G������a�-��{T@��$��|~C�O��m<9�֩ޠ�{U�*E}坍�n�0��Г7CT�`}��邏q*Az�T�8��Σs��z=���7���;�|Y�S� 	l9�Ԣ�Z�C�F���)��^��$5{