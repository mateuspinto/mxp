`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25184)
`protect data_block
Ei9E+igXxaSvURK7Wuu6QlFX5GgAR3nXKTl91b5b0APh3vHfv9me6tGZ6BDREoxn+BFB4ohERSca
1VE9yWA2S692guP5MwJTCSgHHHG08YovKWV8dzPXH86LtqG7MH598PbgBFjjusX30qEz6JoDsKKq
EuwW5+3vp4KjRkDzzEQQiw26DRdcF4pm2Jip893DZ1Wcyt9RNNVaikDRzRlnSYWujrEP4j4rUaOi
H4ZOMx3ipjl56QIyVG/hIv1DZJ08M2FdQ16X0muoBfzdaPiRs0y7PXQtMn7XzWDIMPduBFOonrB4
shfpLb1BwwLq9fY+AvnX2vhGPCDiVm3apz9uriRrMSbNLOPJxJcyIFkwHsxNcSSQekulHllvKBeB
9Q31BbuNnbei+4oiCTmWOVxlG4qGeGDrt4NREvIxNDK4dmGS6ZWndNcia8x7gBBAAIIG2RdBGtpK
PLP1J2tQRINXAieISkLDo+ZQZa7RoPMw1xwzWM+/RVgOLV1FD61QiU9YGMZfHcgX3gykS4Aa/L9l
Cjx+T2fExiCrTiS7hVBxKROeV/I79ZdJlnYKXPVxY1Ry3NLd83Av3pG9eV6iIISSgswZ78p69aYd
R9YDFhzSaZLU2rqRESkM6h1KV3kUwcK/6XKBtucgV1t7iftZaWLzK2lBn2cUJ+jSVqOzR63zrC1o
WleOn/MIkXsEcIUzxhQis/m7M64x8NpSw8QTyvwYODrmJSf1AqxnE+g17E4DOF8+kk4S4ltDsqpk
Erh/WZCISKZnAZNO+VmcEpJWWYuG5m9AUbRoHu3kcVdOQE14OYrYtLrfY09UG+R5xBNioEJiBKKG
JUVfz9a90yKWhxJuIdrO97ezYQeJKThEglq1m0KedS4N/aB9rPO8CTXC9xQjkA5mXTJjvX5ceSoa
TsmuGuKRKs6L0jCbjEkO977MTH5DKdgGdXlO+W/7ou4SbmBMIKuVid6ybEYgSddmxWcaChUkVgXo
OnrBbiFTf5x+nRgMdshnTJiYBoY5JAKEleaGVdhYy6ujd29fwmnO5Ekvb/7Sj6mBJi9AgmJKSY4W
r1OVmIMk/6z/dTJoRoKIfcjhl2df0J2t6dHe5IaMHzVGuexhDkGxHZCQIftHB0q0NjCRLYB8aSkt
DL3xbw0Gjo6n3+cb3iVuIc4To4Zq/PO1XSg358GP0Egp9wHvpalvGgUhvdIoFDA67mqamDEdH5hc
k1PGeGJuLCJ8oQs0PIwKxgxZBsO5DHrQAf1xdx26RQ9Jy98qYhLbQ6jSsxVJjB2lj3MFbj7XtIk/
K0T4/ipG+kcZjD4k3lb12NRbxlYjQHUxnpW7dmajPhNHmqCNf5JQK25cUi59qOph6wuwW4gjwYxP
LYZlwFGru9RDXwqqCuSuRU2nMVT4nCV0nXnidZO/sTcPFUpwloHnid7K6Bv/MRhvLUfCNFFrv/Rm
TeHJfPx0Ccd6skYrnxRtJ06krp+VdWpiikghWwT4I2CThIGJbAwDhcW1cbEeEuWHE0++v7XDSYwv
++oDvwRLCo8Ef1YZ7miy8J2BwiiJ9hAJ4jx4owcJd/HsH2zX8bhsOobU20TM/CpdecAwG6NVv8Qr
55ba8FJ/y2dhQ7C78pHmpVpxKmt6eO2GK1m/u+qkkUi63VrK+W4hFHR++AHz5PLgqLjKiMjhn+NG
CKpOR8zSawmlM1trMptvehfm5iBFtWsLpm2TYLV2FfFBD2M4vrtwspJAwqcQCf7e9lmtcchcUtZQ
UtlQGFxI1C6G6pyILpytE0aWS2pKHIA0DBb83IF62F3EJN9SfxDgBBMfn4SoFMUgZe652zoFdAja
S4uy6fO4BTVHiQWqfp1n6MoI9efJoP7jHDUzwNLfQUtZ4L7Dp0OomdZ8tiCPQ7EOfhMku3radyzs
OsXhK69+zIl4px/APsaGFBfHy7mpqCm4eUGliw9iyHFE3wP6P88eiA07s6YqQVG1mWKyQZqABjUD
4S+ls/4d1XhxlBGY6s8egCnMpeh9wH4Rli0Bocqwaz+9CTRrgdG2yuLqnFtMdIzIhQM2gcYr3PWy
gc2Vu9DZSnFBdUkjhTDusqbRMN6XCGSMyqyEAeCtHSWCU3fpatuA5cyyeWwZWmdvv2VFg7/guHwF
lUvcE98DxWWDP6ipQJQU/9+HS1Y8bEY0MGLI2xJ3N5KHs1kRRiB9IjyS8369ISo+/nG3ZdLgOHbb
5+7Clx8O63eLZywg5QoUtbuV7PB48Zdz54m1wgArq+GWbqBjtnzEJ8OzGpXkf+MJU/HeHGQXKc0h
fZ+L3mLOJgiLqRGfF9YB1ymxwYrhDQdMuSIu+jVCu0QxqFc/ZIl0zq7+NNLU39qk2CGJHV8qjagV
1SIaSL2i+CwW2ksDjCLsE6wYTLX+Z+3PKG5SCpm8z9Q4H3QVneTNmmVaZw3GD+rCB+c9oXvgZNEO
0qQqdC3chtBZ59KU5vBIQdFfKw7Y9AgUdbLxS302LEZTS6w4BTZzOj/AmvCmMeCXgoGG8+Xt1M6Q
DXcjfTLlaWkzDrcYVVzBKw1L9XaTIcyrXMgDu8zBcRaW/sO98vnLIRFo6FpFn0Y470pPDZxlGd+f
oEu6Aoc+YUCusypSZr2XQ+kyeNrUKYDubxwd2W1G3WVjoG5aUPv6gwlkfVk00aGMrqSlGTkWLo2D
JZbfH812XHmO9fLda8CZhUhscI7LB96weAxR3CXTAaJoGPOib6u3enR9vzEjqa0HJMl3wiFDtw34
xd/fxMoClmDER2AWE0+egoQiUfuirPIDSjU4x7pzLz58qL/rYM2yVr5a2Wi6PzcvNDUiYbTTxShf
dsX+9biIWHqaYOSgSWOwNNhZH6jc6BF9QVzgx64948c4EQL/d3hCSx7b/7MhUb9biD6nhpIPcywo
FoB/3vvtuBvyPTm1SbSF6SeOlIFTg9yU5wxv5GIZ8j1KhBbXirPXZtHFBh5ju2gF3Mi5wq5sz4EM
9CIMP0y/xTJmKDkxyqyaHXVZ1RmkVJ/0oBb6fVFq4g41PqLxEpLs3Kg1yD5TcJEFvJz0VCZ3xemN
iHaWdCWuawvKV0Qc8MYnhENgg/zg/rvvWGRalZhSL8G/npRE+r4LOXU1C4qR0dzL0i23whyHk1US
0mOnD8VSK0oBALEZGJjOZyRTxpL6sgtOcTAtgYWtPbuXmadNJU7R/K1PR0Gj/fuzT0xzBOJIiXUa
cc2U0I50L5UtsT1sfc5nzmL1ErIuzra63IbL+aO6M4plmWT4LoiK3KFKb6rM9R0z5EdVFDmts/we
KpCkpoqVzxPcIo02sIf+nf0mlvFeYw/eou1ghS3X0/JltXMZOPZTZzqR7P7NK7YYi7t3c+Y+NEk/
iml4B8rzKFZ4+ODdjdJd32/O/zvdpJBrN74dhRo3I7eXacmTHZInPjVRJDnDm02vvbgsj27vO6hW
zqiBwrjfhNVOJ6in4P0xFvtODLMdSmDfzc82r1/R9mMd6JTTvhFB46tKO+e+neSpqNUShjrUjZbL
RP39+ZZnisuLLMGfY+aVlfDFplIhsvWlvpVQARLi/K6Cmtd87xpbaz4GkBhSzPUKIHpwrVOykhw2
WIRikhsldX2ILN9yx4Bg4ZNLqBtP3ze+sQMZzdqmRCroUAq+Ca4BOoJRfkv7wvRVHdEqKcpD60Sd
ZJIOVu9aB0XrKgQoe2aymNuc1WS8GZcbNAqzYA9LNgSxaPl6uD02zkKcBPVxYofZ8d9kHBthuNz4
4myYH+/DIzPRlkq7ELvOsZSyHtL3VPP88ye5A7B8JWP/oPuz/xdw7nfKZlTWcgMaUy2Q17/8BypO
LPaEnyrC2lNmuBhd3pNGSmStjqRpE0WG9jWPy2bioOvaklgOKjAZ+QA6xWcDV3g4aZWcmC40RbfZ
QcSNfKNnLZfZ/VKtUp95yffSH3w1Jl+Ujj1J6tgi2jZve4wBM56SdSNBdlZd5tnKwixXWwaKm6f8
NsvyvKzYBA4NlVBhyiqWqAN9qfjE2Qa85XcDbr3HkBjEf514Q61tWZhglH+JKUvdgpte0BMQuFTb
wwDwxfPAz6LheMn7fzDAa9zVhfQ0pDnXjVz2FfeH2c/Z1a4Y33HB6EPJLDJBzmBb22A64YFhXcmu
z6xzGqUlZlOfRFrOeatDomDu5KtNbk4qwTE6NY0A/LCewr0USXnvaMDMfkGOJTsdSa3EmrYpUmGl
MPYY8ziiKjdGklSOhHOEDCNa+gCayPLZbCMJA5mJOxNOh8rTu1nS617+aI8XEBGzcDo1XjYvkkOB
jPejvD+/1IM+Cv4FfGFnypoBxKLnowCmmoLNpFiz0QdTQgJ2aCEt+N59hXFlS6WDyHkZt1NaWiU9
XwLkg2uC7/CEEGyeLXDh5dYMsuOtXG9zttKv8iLJPMudF6K0u6Z7FMyZGVFWZz84qYJKT5WjQl7/
BGVo3Vq1LfkFNQoFcc+GRVKHlMX0k4LZ/lXIAWxS/ZLJyOkypsDFoPSnyGiFvNu8jFQX7e7YBS25
ZcyJqvuFTSgvakYSOrrp0zVM8TinEf9+SS2PwyZvodlZyjbxWUM1HLDJt7kpz3t5LNhIuC0ubptV
Sr7NH3KrbHP194sDlJDTqWZOREB+WQqRL7bGCbdICOocxPLmskaUNntgJndDUYwRpqyhgXS2JNMq
NuJ042FINNgzbwnf0g0ErtZH1ZlRsUnnEKvq+54ypDjeMwGOKB3u9A5QK6sD6c/RP129Kd1hn590
rl09lmHGiPWgYExVZ7yw2540TRCxsofeNvo01AEHNCwaRiJnEvadbViN+m9oB5SpkYB2tDyMn6xA
rfy7eQc3p56vUhT81Y7mlw9RgxzoAzJmmXczZIRkJZmDjtarKL8qePL8LBJUIVliExZJXhnm1AdJ
Xo+AJd1AkJ9epn48P1wwj0Ctfzoxefqji0CD9RewM27RiO9sV0/7TDJ5n9w5PC5xQdkY9+H59dD4
hVZWnwdpNNGtIbnghVjYsnwlufC50TnvjKjlecT1zADK2dNlHukiBDYd98BP+DCPMyVP38lWd4Nd
iQgsq4vh3TVBw/99QvKgMNxK5utSZ01xlLkmcZShPz7qPyCGd3CzBuKlwontIkjSmilpvw61D7mA
dfFEYyIMmqEpxQPOR5WJpiN7+vLuz/6ziFu57CLouDVGKtzMufhxMbDdY57RCfS8cqZerh3k58T3
ra0i7zSuu/MkFwT9tH3O5MoPblr3mUP/IXtyX5ce7/XhFYP8sSGN/wQDMUSTPukhbB2s4N9MS7JW
T7cghioYnuyhiAUVFDh9jGzaMiqRmpsYZFb3wwrephW5jLn9MLbQQ/ovH6J8C7Uj3VxCOyJfyDT7
e0j8/kxPxXfEySMaw6TIchVsGeKlh6H+yetMWNOaFUDiG5++l7AUnNtOGoQweUO7Z4CjgnqG7w5r
81bDhTfDS0NzJol96auXbah2bKRZ+L4GkIWVtxUeNz2Teg1fuUtBBEPxuCw6ytqnGKqhBYxhCXSk
3jxewr1mlYSvr0eBJ9EvnnrKOwFlnaL+zzOLS5P6sn6DP4qD7SqLtu6vNs2K0sx1obO0D2sR9+Zr
2Hmkkmk/KUx6WBXfPXeRVmsuX4jAEXO5l8Kg/SfsjinQuMonTGbXiDG0Imt4IHXyziLXv0VSU7wC
raIhySpMgP5e6a5ZLgp5DT2WhRIynpoJQ8Q7irc8XPsuPpzbutc8dAvEv7/e8S3KuVxExg/LAqjd
sSDkRymcBl8J6pCtoa0z34HXvDNnWiknW5JWFVEIyYjSugp9RwSpfN2wE22OMq747XgEtWmECL+F
g2hyBjcDHKpi3qd+cKW6InyRthZQXyB9TswzPw64U9gTvvgUdNAN1DJdXbeR2CnYvt3pOabWTSfX
1nkjSP9r5X4wW31jMj8rUvIdPBGNzkmdbYfiv4x8OqIUcOM7cNPzU95jhRDJCzX0THsQlwWZG4+j
hR2AV3Oo+MKlcPUOjrjKj6nzVi5o8Vu4cNumhvbco1mXSOKMQJQLzdlcsxyOW3Xir+nOIxRoOYhe
GsZihbHh/98Bn/UK+xEu3hoQwfSyiBNSZhyP5KN+lWgFwnbXejrlT70khb7XOekYTWoTJqd+wEB5
BccB1XzyYvBIHRUND9M9IdtO8vS0MVuBhNbL+Dz3/8A5tdDiyqCYEixVDRTnZvFmlsNXpK4b0p/s
FSHvm82WEB5SGPBurxdpdOsW85dlYRChZRmZ4WxI8zAKYSX8Ze1rTOb/Sl0G9bDjVwG/aZRYF2g2
acXK05d67nudZf9h/94IVdRi1V2xOf1QPNwm83/QdsHKwoT2P/GymNawfpYqYSOkqyJbCxz54/xA
z6+zRGmmz4UEc0vGgbtQcXaJCb+/nFlLOW7ZfwPUG+nd5edCpgduESoCUvJfNGGaufCcsYDGQAbx
dE6/X0O6DCzi8gsEG+G/9kvKauP6I8c5SGKArxO3BUqSlgPXmx6B0BACa7oClbgnpjhTIS32NXPM
VUAXgxgDndGY+eJaRcsx3Pf0zT4Y+mRAe79OnEK0uMBUp0eYsjMR9BqOvL6eoovGSAwJBb8l19fw
bfJn1q6fpUDtin7YuFNJgWHnvmW9TNkbfz/JpfBw6TiyQNbx26UC8VP/RDDq34e2tnpbGJkPR5i7
feFhhfE3rxvFpoJsLeKUOFVAVAgq228pMYpKT5uiV5sbRW3idXz6Ztuw2RHa1S2uEgtDJXzaIonZ
RJtc6nizpFwD/M7Z/+nTJNqmC5pXrk0gePBbeuhKh81d6CWIky7QwlMMGdD/kRsIb5l4wuZG2dQb
v0yUvK1TNi3h9dyqKGFw4ltxtZ1MmrK6PBZkEutxyR/YfCgKnQQiCTyQeCWPMHQi74zZ81xm2U+r
iJ8A+IZLWGJd0mdJcBMl2E4okw9/+y0Qo/DRxcTO9W38Ok3nkavLP5cieZlnMOCabLcNEhn5sA33
e9ZOvUfoF+bZWYjek4d+Ckvmehye993d6X/a3wBre5dN+K/CmZuw4NOjHDYiTLbwyw5wDFUsp+C5
P119zUtOjvdg5IwD0ZB3Opxwv+IOCwK5Yew/eg/AGqV6CE8UxK6I1IYvgUpTUvnfAx+QkJqou/B9
j+nBioynzprEqd7XtTe+B7CicRCLs+kCG6uGb4GEnIjpjA20cr/CSZ3jI0qFi4s3KgTp026ItFQR
7kIYrCAXQduy1YcBAJsXJIRpxPZdB3vGTfRB5YMeCBoJQT1iRHCAurFnYixuwZ4IM3HmKlMz+DN/
5DGKJHKrxvXzwoTrhKXbZX0wYuO8UaAGg6sFGc+fIf/cHib3eaN8Ij7gXxvXikY+UdxGdPW4YiXY
+X/In8FK4vTfEjBtJOS50D2MZHnyeySNqmAXZtTzNKkGzysMYg2bNRvXf6DrPNZyQ8lbN0/zWtiZ
EwhsS0qDUZKmqpdjIWZOrU77p/S6J5OycHjt/bWP6fqOSRPm2SH+arFV2gFgoCTs7Nb6aNTrwrbj
vK/mzoJmh0421rftxJ4C4Dln7Wp7nqvrQGGaFBa6H1Wklo1lzGSaG7Ji+RnofKPMgTEMGVA71xhM
1LcOpmPMavLf38amyFBCJtTWTka4i8neraF0mR4x3p8+S4LbXCgP7PJSW3f55QNJETHnC7Fi2Wt5
z3I6AzrdtbU8PqFi77orq2k49YPPf5kuk0xBkvCrpjofLAtqM2UXD4MqcA0vnlWF4fnUrL2DUCcZ
gX/8ZJiYtWYBuWHxaIfpziTzL1FBv3S3jEZMAMvTeZ5vESFdrTEyrdg1cN5rGRJcjtcfrX6ee0C4
P7pFGzQ7Jfv53TnAnSUtkjXfbi5hfhLKgNiFluh/SAnLpDYDaHAfY7FPWjQXcyvYMhg3wr3sExTL
CAmBs6+LjP1c/X6VrEVIJ+F4htAwmeqPPgmy/HVnGnmd09vevCF+qxLLVzXziVhQwoFSqhXrudXZ
xWU7/VWzqkR2sAEhGxwfnGnXZhnSJyezjTzByq4PfX7poJEezoikHMSd8Gl6vv0JK7Qel9a4BI6W
OBp9N9W6YSResON3943HhqjVCL7VP1V44ksHtCJK5LTxUZC6voWi50IElPJuVJz/88Myre4ZVgMw
oCY50UTT4OnLmW0qTfWeQbwZzPN1sG5ARwkvrl5Xua8oupfwH6F8zABaXrs2wXdxzbn5oi5i7UMD
dBTHGm4CJufkdNo28nkmZglbEM2l+BPS+JV0BFmJ6wNeP/kaIh/CW4QT13mphvz4Rm7oB0d0tLn8
nnpViYCNcX+UwQU9S2LU9ULGoVHuH5R6FfzgkTxrYg/JP20xqk9u2eDL39lWyuyAS7jvAJbugolM
+tNtpz4ozEovNEyDZRdtDtp7fCjDj2oP+/BK2ydt553Wr8ypKh8y0vOyI6CRZIQN0nl4Jdoz33BA
7apO6R7BjR2Mi9uCoTUlTWVDkH3KGX0Jng5zbA92GXe/L1kQdvQVjnyi7IqQv+fvkOthGj8wYAXV
Hdip1AsEPUs8LMfl8lUCORHK3Zd2bc3ZxUZ+1nO/ly/yVlAhqqHw2H25DCT2chE46JRveFaYgNxD
uxycXFWLWfFHloJYmqLeepO48joW4evwrKJVPalMK+ygYKVg3V21GhsT3DqBUovjJe6b7vNaFagz
TrEFoRrW0w84YIGCZ7lGQvxkXFte3gk0iiodsBatuF1VfEhiaayzSWTIlE0U0le3Ir32tlRl1pyL
J/xB6KkUCBquypO07kKiPwjfvl+dr6DMKcambbtCxUzxDuZgBsXRU9N9DVdjFww30MGqRQFp7hhp
3Waa+WxAhtGYwdTT0uqbx1t2HHs1yYeo6N8wBJsqrno0DGPONVdz8CSKXQcL/nj0EEdNunMIt+Uv
9csSufdIbn7edpMaLOP519U48P5KdVb+4ZRajkIwy4Fp+FwfOBs7yFYh4FrDoyx/bIdwdtPbBIVD
r1eyBnrl3Cpczk3zUzPZHzvl02VZA+ELk0ejkxqQEG2AXUZ9riXOzVXbGtuOEuduAgTcjKI0BKXE
k9GNirj8X6gA5PUOtbKR+2Y6Ih6yAl0tJ5HQopUiusmWYjo2fHDyaPtEx9qjdjk05PJ1hXIG4LCN
fW+5KrlUozYGt1H74O4FFrGk6hk4lfVDUSXItS7fiEvnA8Zk9eNCZI+bXdxc/OW5a16z/OMKJwMo
xRJ1xneKjICZeyVz8DDYxmy524D3g4L478j6+oST4Ccw9zH6IoEmdAxQdEJcoAeaU0M+DWN7cVti
rm2wXjtRkhWwu4zaGqkAafyjps7G1/94IqpxzS5hhpmISrEsESWTSucp42lvDTdV9aCbf52K2e8T
EVLwq4ffAQs0QZjE1JWKuYjAgVsE4GwEVzIIltHrYl5MKG8D0CIdXo4HBgCpyjjegb9I9lwr1iwD
kXx/Q6uqfHKgasJ9JxwN12xoNmX+rJ6MUzU+TWmHTJeIbpfJsuucjqpN0NIeOFMSKTDvF4S5caeA
KIijPBJrJUxmPGOHNkRamezVh9tXEICCtb5M5KJWmSm5pnMaM/qS+yVcrYlTZ0mF8exvd9co22Tj
BHxRZTBgRu4B3/HWCPW8dGDwd9AYzf+F5rSrCvdAI8UcCbu2LFa2BKZdjdSV8OXNAyWtFrbhsZfx
tEkUvZg6W3+NTuHH1I6Ko2+m6jzOQYosQLBlEFYgfBOw1qX8SGRxG9G5cPioUFFd1FECQ2sqcS1O
2RYULSa1sgfWaq3IbGyQhJVMMxTaedqTOXxXDSUOQk6qdiiDLpwBnFPOzbDgPeRFzBAQN6gC5L1u
jzk1+g+/MsAfU5VCrEmQzaTot/hqw5KOWLobnhQ7H1BTF/WuHZL1Oj3Z6oJukE/dVioqLrEAZhw8
Z8l3/j5ZIqjvp+3qSd6W96cY9BG9NiXH1E43md8vNij40OgYZqLCN0xaN4RSmfjHom83KV/tdkNX
4ruHK/XU3pi2q7fw/sW+RjQh9KCT7648q14tdYEiBbLPShlCfpx0vUzlE4cqD22njp5y4Vk3yqgt
J8UezeK03YnOOP8YNlEDAY2gzmAzLlcyk7O7xpiloUutF5qLWomxCeNke770k9BXq0TgEoS2XEPp
ETDbqq0SPNGyA/vTBmyDpTLLx3+yaCzdSyWdEeELySOCMuNmEiVBAJvwdMw8IRdnbK1AHdXLNMbZ
Vheze2p00plKFG77kayB6PvvRgDArllsjblrDzkPwWPZVRsyYjHxRHZItbWpliQCf8QRoDIODL9U
BzDJvSMllwVYWJ6eEscSVW+xRfjloG8nZgHsf8gVPnseqxIGftCRllSPNgjsj78R6vHcTr9S7XNI
rzO//DSA7LXPIHcv/HYUO7O3BcHB3+kpgm5vmc9sZqA2oYHbPCv1GIZX/I1YwejqgSE1/5w0OuwM
TMqWUhVRK1E63Y8llUOdqvVTlZXd4cn/uPCcPdYqXj7NpqcbFK6P7yT9BIwk8be8ebxjEyPdoxkC
YZscKxMHCW0P/Ym2WmE6yTT7Ri9tWDl5PTRqXcsOizRpbpxyjZixI36gRdO/4wf6hE2OuYwykhXg
RPh+OMO7rmcXU9y8TnA0dtzV/MN7INpc2pNyDEQef41jrAOy7MKjN6e37IaMao4XePbCG9qc21o1
QDyiPbYOau0Pc8cn6Qai5Aln+q+Pc9WPTRdu9/iuQlhQvrCSSoplzP9lyq8sCC8SvQ2rpClKzi8h
msXD/jx1VwRNUJIIaJ1oWRNd2QpoRSM19ondTC1RxYdc2lkF+dhunuJMROtTisAqwR68l/NZG5+Y
eB3XDirhGl9q4Jq3Oj4PmFg9wmkXiKeUD87triDsESnXDX8TUGMeBu/+Sf/FwVu60PdML9Xfc//W
whipGqf97avZw4zp4xWVklVaMAiljDs3VCyq0YpR4n0v53dLd/B8aQcagdsEMDrvICcYIWtV6hy+
9fFOALcYSMzTqczCxYoQsmDJGPBF4f1iXVNl4zieI+x7QJwaEetaXua9qJFmzi4Y5bWZHLzffHSO
JKXAwb3vwQf8jdiMab8WN9oULdR5sHqPCZsC4q7UoWMrCqaeRk7H5FOnCLXasjvEZHngiEkcOxEH
lsYQw/btVvkAekLOKQ4xTlZvBT5ogntcJdsfGmX4yBwzVSE5x+FnYSKiuOGX3jZbNeV+WcD8XyLg
mHyLqL3gESMbd4ynKYdGRhV5wI5YEOguPeWmzp0y7cPLVywKBptsjFK2lESMJz2fLY0zVzL+Kc6f
x2aPfb1XTlh8NdFlpZTgraMd0P/CorOEA5zvd/bGt12x61bwspMC2sw/GwQ4w9JkgqChX9nqeVb7
s6KRX6jDUbLPTz/HihZSEDnLrjZnKCRmguPfE+eCAqEEIisLXCB9hkQKd/xBNqFVTBTNhe+PkEo8
5P2z4lNGXMiC9cClKEqng+tCrE2k/O0w7Wjsw6YrZRKNjEhrywc5ilieDFJcGs8Qv7BZhMhJ7bW0
LXwpAS99ublinN2VKSlEDUKDNc04Y+z44/5z8fy+yn5Iwj14olNhzXmjVwCk5qJId2WcAzrjl1+W
m8cu2o0zB1G6RCqyN0+SbARC0KTFHl++J1TTxf2p7Mn6K5rFNEr9V/gGri7zJtycPfMiZclqW7gI
90xxHTytVX+QjTgaw1DIHzgMvWS//MQvnfsU15msT6R8nGcQsEw3//FwrGk30Ej8aSgAKyWWHFB4
+0rU8WH1KBPPFOuz01gkEKQX755RjSnlMth9bIjCwEoX8cMxeDaFcek73iRaUYPiyqBvqTtDlh3k
tRguvRyoX/HxDrJ3CboiLFvXXeB+9k+wl77Sz61IR4/bhzmzkoX0fS0Ou6i/9EN2cziAXRyJXIYL
thTG+XLt6BLSXbTTkOcSuxPLQLktTfAWmsEU1+T7aXoGTvj8N7CgaUhlsB4EI+SQOuARqBsu9RGX
dyABoHcVHMYAsMCWJEmeDP7cjq0Y36J1ucdUiNc+Y5mYHU2bJrVmCBJqXxs1jbXrQNptKMtjLWhi
gVBqo7TZWUKsgCD88z6HFQHg0bJYdPJqUYcO4GDTk6NkySLZK5fqE5IPwI+tGIHfBHbYLRSNyDqZ
Jhj9ycDsO8Ewq3srEY/iheK0XRs/GA6fG+0vhl0ag07SN14Y0lgAtIjMNJaoJILEYaBl5nLfP1+0
ks3u8Th0bGZ5NTxtWGWl9wz12PEHfGdLMwSr1PV9qRPc5XOvxIwKPy5+BRwZGbicW1nA3dWZqsrx
2pcn3qTYkTrjCHhHxRT/cJ3vs0/d7QWbIFt3D2gUVvjG7mzfLe+7ZbEfD0eoIjpNP2ZMZcgD+/L5
Yc1PwaNrUVjtkaY3XghPjtqUKL0++JdJrtJ5aHhQ5hmIUlgSEjEBr3yJkB7mRCwUP/XaEnOcwuAP
hv7Gjtzs/hUEwIs1xmQV1TO0zEkGdlCAfIb/R7l1sDIQiFfnDvw1+Wk35jWc9pCNbsuOYR37SMny
INs0YG/+4+cRDunirC6msULDgyP1BPfri37DQq+HuUrzUku5sJQg/BTrW5uBcTsCpEOVoZap7HEs
bRXWdmYC/T7Rk9IekRHgZ2KRvWSeSCYEeQROUZpIvK5jUueRE5lkptu2PvEprAZ9IqyYefRzAol1
K1uBMtAvlSxsnSgbQNXaIpKRDTsRwHAFNxQFD7OdYbqjfxL+tudXGPBTmBeng+78n9F1yXdW0+lH
aF81t/00qfYyzivHRSB0kjygFpoTyAPGMFYpDaaWbXqDEIEqXML7+gAeIQSDTIC+tu8PZubDKnU5
KzYaU4iSxMgOIRcTfyhljcnFWkgIaF/XbMt+HFulU0TNlgBheERmqVYElOyBkhffobtcNgVVp9Tg
qXwBQMMNxOoQN1p8KvYFwFXuGTtaL4mJHzUwggphJTJP511omvXCOXKUCwooE63tKOVCmf7effFe
+r8fpNo78CDx6Zua3ZZt8IW5jZWq06mb7mJOoZwCRspJhxGcGAUCqbRa7A9vXxTmLzuMgLntPOLK
nLFBEqPHDFdQSa/1U3B2yV1ROyQoKT454jCOUz2fI6ng40w8MyiBQ9rjYViwNRhNOX37PLT/jjfp
zMQwLHRhz4XqD/K8fLwg1yWlXfzk4BExabDmSBphQHzQPTXddMqJL70faPEbRzzsG/qCnadJ+TFE
F71FX022Rop2VmLHba8E4z9v093FYKBFk+ZTJ7SlCNaD6Bb/u1FYdd462+Ju+uQAC4dwlU3aJ1MT
nsPDhdfHOZumlqCC/LlO1mSL4s3Fmb/V3HYt0d/6flAnwbrun+UQ3jhD9fPvsxVEanlW/D1Jfu5K
TRjs1YHrjOQDvNVVB7PzR1pGYV5yYZibNi6KdPk/dkchplVg6j8qr7l/nnfRXwxPlV99fZV7Dd64
n74wPxz0swxmb9lJ3H5cnUCMQFYHyNc7snaHguoVlEmCAxYM28TCImkbbXEs4v7w3tmZV9DVa8Ta
gP4/vr+biyUlFZK9xK1mO9G9VI8oYXkbqi7CRZFwiKKSQ1nfBJXy0pOA6XIy23QAYHMqgN6jy3Jv
ZaDBUFgtJVZj4LtNetqCKbgFc4C+zBZAQ4STsdEsSWCbJLSMjxb+HTKl6s3i79o1xpidzEtvW9Ph
XqUOTxYMr6HlnhQhfWYpjbhB/pXWtBMN+y0HlTTPHI6lexK8KdCJPa/oGnqeVGC2Y1fv9gIY9jZQ
KB/51ACK9SJA4eL4ixSwpXaKnaDVkiGVdt7Mj4ot1VpTLeXBNWadpYNbd/iVoeHIQI5crgphY+Fz
E06N7iXuRvTOlx5U3Fd4Pqw7P8Z1QB3hhq+zc0e2amf4xWZI5cLE/PFY8WIcmGWx+QaBIqlhiVKh
EHvp3/vubnEtaTPQqeSMDzeK2giJQ0/4XOrapncU8psSRc0qQW9VeK7vPkbb2h4+fHIIHNMlZaOs
HyhAx3vZbGnVbIRBhLp74oVWIysGyNeKDocKbI8IzEl+0X3Mgocwn0z7HXCvIysMtGxdNTYdSafg
0DJWA2qhowHaPs1vmZ9dFaGgp8S1GqS6yIZlwPmsytnvhoJvq7cBNHuBhgH0C5nNGPjmxyKnFY7N
G2wpNud0gWjWpF7yVruj9afreWbXFeSQjuIgYlqRsYGLn4lVy2Z4oXAgWEVFxfIH6mEwA3MpIBmX
bkqxv/nIivwV6hpVFMerIPjq3uGVn+JqpL7JqPJxV0eLFNKaE8jRjSd4Fal0L66U/pTOgqXus1ZX
KmgDQzlJ0Up7tlM/mjvOotWmjQXAW7A6zsrm4VMzffFnAWGkCIMyf2Zf/WvS9RymJPtAeqf5vMFX
eMKVg47q95eURsIM0o5zHbKWwMGqwuFCSmZkqpVT58zHSPxXixfjJjLCGbTakLp3od8p+8dejYP6
Gd+8Z22aHQrueDNIyPQ5vn8WbPkQivw5qm+TSqyzt95/UAPW7HxvBdd4D2TV6cjT/z4AX2cRUa5x
g+7W0VhfGDekqroKMTI9+t01nunuy/OQ18szyLervvGCsmrCiGnhw/CKGoqGiYnIekFVQ+R7fQmE
1UVg0VOzrXXLWhGEHHRQnJLnfs8GNP66tRJ2aeiHr9jwdnU1DJ6/+PsQJbteUQRcr4nD7diCPj+/
hs7jzTU47JmzCr0tyLHCPRhUu1MEr/AZE+Lv/Nnm0vps/U4S1e7yrQ/E6bA/n/gKZtb6pCPgGO4t
4NvknDAVv+k0W34OdiXT2BbTUb4CyEpkLMEcIyq6nCexhKvWgSMpXlwnxwuAMuzuK3WN/TBQX7V/
jHcwjgBoUn0zMwTqhNwfblOD56ca1N3amw2aMqLIF/XEhH9rU6MQGAbcjzH6i1iIT0vD0BgjxdIh
P1XyXUmXNRaDSlilVtHcH1fjfeWH4hHJBr89gx28HhQJDyr4pDYEON4hTP0vZe+ip4ZzP9ATjAEE
pib556bHNV62ryjDZpgT1UD5J9awcpRH1ohJulmP1HAuk4n2kkhVVkziWTrOG7/+AtpEcfPvT2qB
VlHzNosro4Oq5sGOmdAInMQgwoWZamlPeNYml7O4Lb/NiYTCaD8IBoLknK3ENIpT6use0rSfPFp1
7+oOvZ7DxxZLbeWE4Isn+MGCNI8xg27uW3Jfh7v41RSC46t72RKrD9g9TNPL4prf2vJjNH7AZwXJ
5cvDpz7jm7VbbWdC2Jwlty2nIkzikrwiHPqlhUQFGfXzce/cTY2+UlMbRcpfza/+zHsrx6mfNwB1
/OEGQPbY++BTeSCFfxoLoD6Tx2Xa45iSNNVJF7CAT2RhP/TdgnCQK20fLM8AZ1cKTUy3+fhig6Bh
Il3V3psXaM7mB0bqW6BN5//jQxriTD/7/wG3eehS6+d72qyk/WCrqXrktIOBmzjSM79aibU2aSVH
KFadJ6QZPPU+1AdqvBTGeoY/LXdayFLLF2pFcPtBGHobLRId4NL/kUSKXukGsCvLVqyeFZAPGJGv
5dc5GdAxl+l81rxkdU3eJ+5AkF2/lN0V+x5bpn+JZRFq6zTHKcv2KmaCTIFHn0bj9cPqv0rzi29S
4ccvxWQcC5tZ0wVbNLK1+PNRPlhK9X5JAAkGsT0/IFq5iR2+5P2CC6LUCTBwVygV5H/P52lDwTd6
Kiv2NBMP4xb1G+h/xDjuw6UHFvjpFn2rTxG64VWQbdFWBTNo5AjKmZKoMN0yPycTGh51WR0nKUrk
QX4q65ydSxs/ZDPNSdRg46RTw1a3CL63DeVCuaVgfOnl2JVFyfvwX2fSjE1qve8MkHna2EaT8kGk
yGSqHTeDqN+r1/kKf90f3Q8qSrjrTNKcFIq9Eo+ZnsW6XgQX7pq8ntedPBQi59R9NFhtxtmF6mwD
Za4GEmN9jiPi/lsvpTMQ7BwgMichMd6D5T3YpJkJ3BzE9uLv6qeQEHbP3GKRP+V+xx2lafgRx/RQ
OCBkYJLx+mpuHYDw5V/t0luWDhrWJewFIxEGnq8SMU3hWueVePV0E0nKm+AL5TUP3KDwAJjc8WaV
rVA8LVzodw04YbQwAj92xurhf0KxNz4y6O+epEUYUedoQ1xMmde9qIIT716wNzSc8Ip7ZkiJv5Fs
g/+F2DshIRY7bLBYxTZLd39FVAoRC/rWjK2+sr4GPX6WHTtfefcQZs2UNsYLtTRaFloDwxtAmSRi
Helj3pJZAqXS1T4FLd0Q2pjwTewSnYn2lqzvciX8CH1QJXYFDnnJFCZ96sBcstwqkGZn2VFH2L+J
1D/qbibt35vgQVVAdo0sbr75QTjU/00ymkrxBSxwixrtlOKYCSH4PPF1eoQGrzhFr2kBMofN0HYz
rzvslZqal5yOi3d9d+kdGX1taDb0Cj9xgpYTBDLuoxj5Xqi+463izBUGE7hNJTliU/DRJPzA3PvK
xKIF+F4CMKEbY0QmfzmHmdFGyYXyiQPIKE+IYo+NS0ZAhpBbyuxRtSvqcRtlF+ch3r8r0/AgSI8I
YIpEfYvFiQZ8mrUbovvJrqy4ICHXqpRA9NsbsfZ60TvLLU2LMEo7UNOJY7h9+b7c3a8LaSgNr2G7
QbZE0wfz6QHWEi9HC0dF7cgHJlTztkwqGC2/F2sODA7O8VRq0LGR7TkwMyRiWeUT2amxxRlC9Y5W
lIopd8Kw5caSIn2muUQpZp62f3x+s8J/HLbcvuU+kj6xrPKf7zBvLFUJDuOa3CsmDOsY3KMoW67o
AJEcY9NMTVznjtpnbSBuyQLzhcLvB8IFS7irRiNivM7tccFYCDsaySx+zMKPawA+lJ5hz9hUn2WN
NCJPt6r0uQaUutoDFfi3KQYRqp+hFv2yHt9UwTUqp49gDz9+PwstXIQ9EZPbaCCVI0ApixrFnnTJ
/qa9bRyc1ksrFBn2A8YN1TCNM5xmaIy0zKJhw4Mw7H2DiiU5VLSzE4DGURtvV59QyCpjDKIWqBDQ
e9DaLjGtWwEVIpB1LWF4zIUX1dIgkQ+DEXWeFsDh4cjAYe7ND+Ebr6XYknXOoeuX2L9L1cT7vH31
nZYKC9vL5kuUlr0fevwQAZomIVBMMtiRHeZoI+gkSTK/fNcoFGtb4LVaGlUg0nrKdFcC62wfsnz6
zDaGvyopoHp7gzGTqFkUG2wVyUU8tjXWywbcGcKUGZ32THLMOYoQbVy6UVMSCRMrUSvNC66Ao8wQ
Aneu5sWCfOwsI86X+u/p9t8yaee/Nf1ACgg6fA6tGIRrdF89/v7GHUPjcUPit9scJc3LjlJhAg1R
Rx6KsmGZDhZMTw8TTLPuP3fqUvqucAKjpRFZZ1y/ES6QPvE2HBTmKh1I8FAf/hZ8TkQ4txdaGwWp
t5vpAD8/7TLV8mLHXOceLVxqQzX+tzuDwPbeocp6WMYsE+ZpYJK7zp7mJdjnbWNiwaKVG6DO6Yi4
c4EkQqq9LXuzYRS5fxCO49Uoif3PgOL7vqWOG5fGKiEzqgck2NWBtE8OMkWuWQXFm5MDBI6APgvi
25PhiL9oQKaZGsEgHj1hWXIBBmF38fytwtHoli9bhF13grI/wKNXzQGtXSV0bOGxpiZKaWhEnsX3
GPd8QkoepnV8LprqGOx0HouU0aug2oLkKPmFnirgyc7TxeIBNLr3OjeRo0mK4cqwR81/SFHV9PFa
KcmVU8JXDzSRivJoIlEA6PbF2ZW+Egfr1AXH4OyMNkajkoKZ7VEKOgRl+Eqc8mWG7S+7oS+q2DP3
RChDtQSWNdLtUz5jn06U/i1MeUgMdX1BO44U+rWO3yYuvhd+rTtt48XDLnmkb25Yk2i1Qn/JHwms
DqSCXgV6UHcnRr6wLo7I4C8elVF2HDGMylkfFzdU0F+LxwzLHU8TmCUzQctKgRD7g6QOHjFQOGHg
Y0FuMZ29uZdQTJwne1CupNgE4PIW1nluZu/stW5J+ItNZTezgaQJjDohVkxF+Ndu2dICTsfVVOLr
votcSB8GaGalbMrCv+dL1wgJCs8hivkfDlrkpRmmr5LbL+4449j5iVCVisbEkkSMSTJgjEtJwv9m
dxo8HNo0ShJO7+BFtzlST9I7TZx1lqBgJlFMYwIgY1HiPok4ocR13OBQvzmocDVwuI1hJwRWhy91
3ev4K9fk2UDHyIY4dLDMQTlLzz6NMar0SdqujCGx5Cuo13YWLOM27dL3nFCCAhxa6iIG7Ufmjryi
9vtiM8KXcyg8uz2XdNewMIlyrk+Q8xNptxUfm7ZgLchRjzSxRrdu+q04ejRxYMJbHHerf/zKCVWk
PQ8QcmYcs+PLjKR6zxD/9nqxJvuLJhllfFPHbodlvK/72Da3MQ6v7Owtj4BVW10q0BeCFexfA1py
cnHcICdvvMs1rxYtz7KLDGJAejm873J/QKcc35ceojU2TCsbLBcP3eI8RE6HXIJAEV2bWOeCKGHJ
uncdrP1UoleHQ8brrWHTmrl5p1IbxgJBKliAq2t6IeWnUBgRmaGsTllb95X5wrgPZ0sLUjM2cBhC
4XTQkcxjmvWgdYZBEFhA9/fo6s6pmfAtQJ1F/V3MvvRmyG2uCq6x4A5/VkIAXaEjIm5r265eBSg/
i/Jz9yASjnitTOX6dUlR5bFHuUzs3HV7XDoXN2LTtomtRsPSt32DdqYL8rEnEyN3TVSFWDqTQU7a
h0A2z92d2c5Jnz1TEKBsTWx8+ILFvNTCoffxV/jOiVjQUEqt4YGjXomLgfAUDjGN9mqdoJTRehBU
TN8SNHqaERuv1D/WfKkbykCl7QvbxVE6z7G3Su1iHlIMmwdH+DuGNaTwUAfeLULsETjv9yWV2khw
4kaEw6a6bVlHCFAhieTLVGnU3QROPfJjh2QMvPGYJlJyFA29NwH0X8E64sF0iNRLDcyTl0t1g3XQ
T7gWFETUKLdmrqN2h2m6E7LarTnj6aunIMxYzm4rITNkZTfxzkbjY1jIddF0dxOK4iFxs5qdobMT
rBXjmv3pGc/WSkklHqyc6WLV3Kb5XhLTersy0kK+K6cs5/8DkcybyknTIYi6bSnvPcohL9XV4aN7
g+XZGvejzDNfon6zwdbpCj3CUKZ45t+tTEWTOcw9+BSP8pyZUqNp+EOyN+SUmVcFLo/tBnDHMt8N
LlaJ2E3o6IAXKBx38sGLwUM9pxbyLQVi/i51Xj2GZp51SyuF6bbtwwCk/XRvqQ3jV9kHThpPWb4T
7Gq4ySnYIbK2ZO96FEfr8cp+q5aQWSNO3yq9Q2X7WFiPubqae330Cmj+8c2mV1O3QP+Td5X+d/H1
59km/J43Jwz5rq6wjxrGHCrDF7v7BPJOsY71o46n4NtKv+7X3WWfzDlCtXfOK2s5fpqlC6heoGc3
UFhzw5KpgL+eA4pcsAhfa6/3bZQL8CoMi3oFxxQTquLW3yfDG5Lqm1P9MU49BSiHPwNQlXyoYDY8
ny8EL9zIPp287X1z1gM2MkTAgHW9K84bZLxdkNeLSobnfr/8OW8CyzogBlUsrCuceakVgGQ2X6JF
5zN+zjniPXNNA4IcW7JOVrMbyCyEcdD7nCpnqrdoEogBAMjb5SN9VSfKUiYTt6O2QXyDVNiaS8mQ
eT3n2DC+b7p+ZS5ztjoQCU53kYPz9yOF9x6v8K+lTs9eLV9GBSIsxiou7qM2lU3seNffCPEqSmQW
PCk9LdbJc57nHZzdtnYpc3487+QYXIwHE8b3SS8Nv7Y07Z8u+5A0h46R3X+lMc+QxfspDGaGTDOJ
QF8D9b9CUY/MYBhSNNfOXW5iyy8C1zZARJamDvPpq4L5EpnY3/qvulw+M3cV25m+e51ZCtNCvTXL
8MEeApKtkf/8UqUouz3MnsrWT8fZ5OacgCiL9figCAg1DAPBDk1jw71IgYebkvuBJOV0nBqKITOt
5DvJbUejSHnysXcJzmDNq58enSWHpceuXuRO3jrTJfoAmK0aeMy0Aky4RvJyMN6yt06M8l0EztNk
vZkLymcnqScHjr1s5SsY31mZDw4BdPJNRk5qyEh77hggYY7vvxsEvLEAR1qXPrWTsuJYF1C0DubV
RN00BlFluQJLOyWLpnBcHCGB/VD1H80J1Yq5qZpIWpEuSFm8k9EIC1YyCxUBIN4XtY0yfkWB0Ehs
WE9LcJM9t98uzyNOklha5zntsCausaY89m8Yi/pcGXD4uYaVKGbuXvho1jf4U52RUXYl8ZaDiJ8F
7BHUjuqZ4Xq71L81tyaBTDL8ntMr7WPInHPHZBDzHAU0muS9fqSFQpCbti3ESAzhgfSHgeHhylqk
mHo4PS4GuEf8Hbm1nvDwwjO7tbKauL3ilCD7npQYbotGPNAhNmQkLlT2EZVjN50R3x9BhZSkYyCU
kYyBuxQsW9B7oYfP+hEXq/f4GeeOmFPFOEbXb0J2uZpVnV2TddVfC6LxZeXCWNDcwCQ4OUgU2byV
XtNsCIK1+8+HYi+sVQtp8CNl7xB3R5/8kxhe2dkDtxScn3XJLMd7bPfYrhfUPoGmWFS02hwW8L7T
ZMgGkkpVI1dx6++DRMyJkCol90ijeboZ2i3LXQDMpOm7sLxISC0KaA2IvCLtdUSCiFKRPSw/UQ7U
SYOLp9C3lNR12wKiepmljY6T218jD+aPA+MuWeYrgTWbkgNrfSEI466HFQ74Z0bdDnANNiVByeQ4
Qg1sBzQpB9IhjP5dSOWB88caAMO8nNYpINaQaz14FpMJGTabWyMm96JSKzm7i019jIu8gZm9SjmM
2UvjmBLCmfUNEXv5bF7JIuqA8ssTXwQAosk0abXbz3c7gGOg+Ft+DRd426Cg8qXcVn4TvP+/bVP8
F9lcIqDiERCPjBsQyAyTm0MQH1f0ciDwhbnPbBPbOAbRQ2PZz8KQOsFqemwHUr3UnwNyYY67vBkj
YnZwE+wABoD/vNA+ldDpCwLKQnjnduRA/CSdwCj4CZu646RvkRuM2CYYSZfMcmsIfvIE0riiGXUA
Ei3fWKRaohEeGgWReH5E68llIKb+lCeQVAdtPwPU/zC3wbAc/+MR+/OL43/2nY/xDPe19z62d6G6
HrsMQRdtsGZQ/XaTjY3oi000vhZ70iknlDqm260ulvW7MYRQodmYsYbkdjRRz0CPR+NYCp7U9FSt
ydBd4zpAHlu9/r2Fy6KvVrDt0RjFSPjNIytbLRCz/GYeAxWdtopa0WnqEfade6qB6ypPhQsLLcL0
W2hqroY+3Nf5BFaBdLXH180YZhp2dg+JI24QmETjpcjNX+ifF47lSUirIwrmSFF3DJ3LgDwJJ84Z
BeR+772tdgMKlEVjAXGa+HmOvk2AewRHZyLm+5Ix7Zeo9IUIx7vRs7UzjE0GN3Y1NCuxQrn/usEO
fkIWDYLHsb+QVRpgtjYkkhZ/YeNA0sa5wFtGe/xKfIcxzTNxQt2a1mynhusYXHrJgvGC/sL3F/Cr
7OM34NI6raNb9PtkisKtlfuEoV2xO/B8/dMWrLor4nq1J+3fAIRjTjnmuTjcHwq/T518OYOOgB8v
W51WomA1f5SQRcZJsT6vxSZ6gLZfdypu+yuKv5MXLullCiSdhypf+752yN4AaEXTqpHfQ8baSIUg
HxrX2vnxjEMbvy2mwzgsNLHl5am+WIl6c8yVmg9CwtVmy1QiIXP9DQnCZHcN3pcM9CuZpJkknXKJ
fM/hbZ22ARKokokEVbiIYhEumEmLiZ0g8pCsr45fw7GG9nsP7Utmdcy0bbp/0PN0VPZP2Vj2iyuX
5zSr6InCOenzgKXGVdJsjnbltSkB3QVMcmBiS4oKAUBXGLjWnw0mWKLw1q1UQ4LyHI8rdklKZdS9
gYm6Obw1cS1Zf+FEgDx3ugdDc7JK+LysMd5OS7wmQh+1t8+KHqez4I63we0uD5GRG642SoXxmA9B
7RMtk4PC24XGO3HKlE4rQ4pihwt01LYWE8POu2u4ucUCBzzckR6NSRUGXFdb+sMAz8NHgC2DdHie
oBirQjSnL6ngPPz3Ah90hK/ax/K3Gf1ltYC+LGT251BETTbpBLI6jf9BzpxZ860ZnwEZvMgwSjhH
CPE+ngRUmLQvL1vbnn/CPkkRUnikFBvhmdsNuPW57yeO9vLndCeZ45WfuWjclVKPvvGzg92qs/yk
KrBrqiUMzevlqQgcxzlf4Ot/mxANMZbtClFKLhwtKvQeRj1WNL5pFMuxyB0HAq5ljDV4Qy26iRZJ
3FSj9EhgpLPm0FWfxoHJmrEQMY3baQTUtqOf5Q3O41imPsnQOXsFFgC4xqqqDybHId+uqo4ODrhp
dIbcY43lSP28xdjPIY4Aw9V4sZI1g6vJSEeIFRk4hP9ULI9lbjEkPlyADPlEmsSh8AIUrb8GwBhj
E/X9x9hcv4OeGXzfNCbgntU48pq8BXULU0idDia071bIQdTMnD6ktv7P00MIR1ER6D/Vbew7aYiQ
YXU3p12MoY8/3KgPdXZgnKFHmmtFKt3qXxcy3CtTwiEfEAKJUvIomH44Ir8mAxhTocLUGp4ueSL0
3qLwTUW74/kh8I+f1aXKwjGHJ91QV1fXoG1OBFUZlUJJS5X25u2VFUSGRinKGTM4aZvdzNRJfEs0
odxVqNjOFcs7MGf9IUdVWe1RpriiBC3kOTmp5mFekPNJrzVTSHeSydnD60mmW7b2VFJVz1WGbHvV
frwWM/Aoijmaa6yF4941vEALJCPlu9syqgif4C17vut/WIVlXYnhIcem8/1BXcMD6dZiZe3ZVCfo
zgJotk9QvJs2Uq9ORpJv5KPoSV53q9BSgMpP30dhmFZjEJW8ILrc6S8Mw3KEHLGppdLqn+D3xmT7
N4oe6b+jUbCHrTpC7LxY0FZr/x+jI9w+aJD1LDjW3NraeYh1SWHks2eO+5IP/vJUJrfk03Oh/Atl
JG6RSJmzf3/KJ9tb0EYZS+wgmWjXuZtxV1WC4QPyA7196LU95VwTrfBtoaRb5ES8Mk4Pz+wGOFv0
Yq4/ns2Ul6r1J6xmVYgO49g00wucBXPNeTGMiej4UHiALtihEf66wBuPKwJ+M+nfCso+Kqm5e8Sh
zlrDRcQq086g58laCnbPqMJpi+B34gxmZir3yYW0PFbxg24OaYCLfIW1oD3HVGukoF1hmSHvXz3R
NFgVDpSE3svGR3h/S78c6XTWNfZYNsMMkwCHpMu0NnNOVKsnRmQzrGdK9DBjyfihhzKptTc4kcdV
nk5ZgTG7rxvu+hx2i14es88TDJkbWTbFEwDShfJ4VQ8Ixwx+OQ4P83ahnfpzSnLfBsM5rG9GA0C9
+GXPSaf1fVyABAXz2vowOS08xdSMDzjMx0DauNeXWoLJ5rl4CMUz90D8XrUjFjQX2+XmIrEmOu1y
7xO+0pqfQrIZRKoD29sYUlpXtLn4Hhv8FIDi76AdHH1I60erg/DfhL6JfdI7BwUmxkCiZKo5WmL0
Wpp/X45LZr2htAXpg2XUbpTKxjJKsAYjeUGHD/goldBcjTpEkV0TrfF0Hu1bcEeokUpW+6BZIDld
jf4sXhIV/6ddNEO5VX97lyoiKrZjkKhdJ4FlSKom+m219gc9vuZXHGr91TjgUu30H/LlYFz9pSwJ
Ml3M6JUpVyCFkUkRXNe4PZfRdO4u/C7uLbrOUfqbHSkOI1YNJLZDi1sUddfmaERCDxiVBRRayqxQ
iCAHfaSTCeGPOrlpDNyMNzC0Kpc42T2UsPfbSqzXPXxIyTllU2M0H27y8nLgOvYGeygMVljT1cUt
E14tTk0/5//Hj8/3kJUoIu8T1fWcRC2Zbplb258la4Ux4pSyGOR6ADgRMs1cq2gUzmfiA2d3LJca
7ZZYzrsYT/i684X7k+N/e+OdRGAQ+uJdD6lUNFPuMUiggwUbPyIStt8werBT2LF4mdy7zvKXA9G1
jBLKjK8uAzcteMcOq0r9Tus7ZT+k2GxOlzeu7t7pbjLZPDxeKCVIWj8PuSItB2diIVnUd1yvxCj9
u/M9mD/O90g9f0RpskG6y2/QmOi7RPugJdT/DFeiXwRRYe/6t4NB+sjTgVKv33m6q17eLn2d4vZF
34ZgwfqwxsEHDecQqiRzL/rb0P8S6KGbMCcptNondmUPFJtuQ/LJtVnIfPmkyl9Vu3MbRExMMREt
DpFqEO+7zG9DCuyvWb7Ny7CWzezlMOeH5j1BsnZISUB1yacb+8UXXA8H5KRF0a9Z9nHIU5BnhNIE
uxc/JBkDgFEsfZEKTkFbGpgDRgE9AV1FPhfBSkKvWknsTeKG+evjtOguHFsZtoAndE5GGldbClMS
k+wx6Y936LerQ2t4sHLckaFuxoPbWUQ+8YS7EBNaWaRcp9O889iIXkxNt5Eqc86lu81LhzyJE4GW
mZig50sVj4ZVQVNHduFF5QdLb3WgZwT9LVrRAlpvVzxMwFQy78Isq64cLWGTbgX3sXPywm7D3/vB
sUuBgq7XdujN/aXYGZHL4eqdcqvS8HnlXYdNaL0UoWzsAcwkuUJxeq/6NGwvf17h6WxQpQ6FL91b
AUfwsz7B+ni4NLDvUEpC6YBqAs73572ok53bZhIUk4RDTKP7gme/lnI9EB/k+eofDdPw+zHbXRlN
uUNEqplFStTW3WSFNKhNmZTrkWadAGYZrZyhiUOrDsdXnJGDCxWwqSqmNVcq/4Sm3Rq59vW9FTxj
JJbGNnSUnin10O+EO1bPmXtyIDjVKIIGEulUqZHhZakRIvJ+YRAbrygkANOM7HMHkXF5zoyeYR/A
lbrUt+f9uNTiS/F6aK7uBFdcxKUg5X9MMMFIA0d8n07ZcPV52nhhm2dvG860vNYDa9d4YCQa+wPN
BbNOsMqe2Ny5GeFvNc3v+ZX5sbR5DHUnR0a524fP1yj5VE9/3thzVn04/mz+SHawitimw5uds/zU
+ruVJZTDLeNSlzXAD3HTMBC1Ny233HAH5vbK0SQFaDkbVrv/90TWbNL/LJ4/0cm4ne3ACkTx5zrJ
WtOL+KworcxhzvuhVaOfPB2avTVAr3+AaddAO4TT57aIMd2TQXF3CdxsD75PVI4dHLQ84rjMQkK9
x3WqgLUelxhJJpt/LXtzu1A2qd6MtHdWNb7v2ce6BnoKOfFpNG1xZmVCocb0rMGB2ydG1CdSYePL
T/GFebV5PvHMx9aBvHYUvZTi26x1mbvQwrB2AS0nlz6ZbXz/m9vS6mv5CHBrqG1aSdGH/QTKbIAs
6aamFmHJY/b+VqSgyXfQDGVhmGQeAysIbNKrwASOzhW80gtPdYf6ILNevX8m+ZQeVQZ4h2cMkdUY
Je2k57TqzSzoxzFUjXaF2qj5YJmT3FZtt3Mc+ohv2QywIZ7D/xJ+nEN3Umob4kl8SMbNCLQ8JSRy
3UPkEvJP/uJGXCmPDNnOZKtx4lSU40FSFhF2Zvp4n70O/Sd2c+kHLrYXlHYGzNrx7hIIjlP+QATb
7vQ9R3+ck2FQFAtplD3+9LPsTsDCmi3b1lUI+X9/AEW+M1i+BcABhKoYmNz2/yM94AZABBxELVt8
/xxmVMdYSCdzB6krJQ/zP0Ldc9wjif5RYop3ypfxQ8u5gAEkYXsgTeQlcKiJWaxtwM2KtL/aI/Lm
1llyFXLhnZ43pBqXzM2zaC+kinCv17x2eCcu8woe3XVX/1I1wVbT0A3yHvDV/I6n1ZCfCjNd0YXR
WWGuonTXh0rVhY8t1N2AE5FuJe1wXSPEC+YOwJbq731EF1AtJW4E5wC+h0mHADb9X/IBxI6C+TDi
9Qtb0MaB4riY3JTTCvyIBYtzQxPE6cs4grwJxgkZ13Q2nmjvwBRGlXFDE7PyMK+5HGpfXghHmroo
GSW6IkWKz524PJ2TIoXnB69o54EQqMJ3jblCr6/w8NjDAI38fiH+Zf6oKKzXrMJGNsbROUMKqDWJ
YwOI0N0QqgbJVCWjEJgN3e3yASdcKbOW/p5NcVRkR0vEGLoC/pO4laLuhXssWmXoWN/ypSAYhZCv
YIzq2gKDLRh4uA3XIkTBTN6u92L80VsQPNLQ3D7S5LbDNL3o194XiTayxoFfhybnz7Z5gDHgnYbH
xra7sSMT3yANcoENqhMThd0AMKYHgO3r7ljvBDt3usCVOi5RVNUxIGpzCS7kMU0NnlLt9YFf9UTg
Zahkj4wXUyu9hRATaOYFGCti4QoY94NEUwFPHLVYOUvLOk0aS4KlBKA58njkEzsox/HgpPTaFU9q
gpIyn8X9/ZjBpW007yxg8HDNsZs+F26pOHaK63xF9S1XQqCyPnVBLs6kveA3wDPtxFk1Ceuvn9ce
txBOGADHColwtHF3P4XqdIx/l5JuhAYkSgDdw22+qUKO1hQIhwCRdqVW2cMJEY6JUzoJiio1IOxN
FazRDansZcy7oKqxnEas/7kVSWIV/bx0t6GGtrO3VQ1jcprpxb6K3xGrMipb+JMzL5ZI5hAp09CN
D1V3pZ8Crku9Qu+fquQaYgCfJXdbkA30ynhL48reZbBzuT6naDGWKpYwY1FmPgjAwS/8sR7wijm2
2hHYZTWSl2nZh5XCMc0zeK78X88y+krdVTLCbD9LmG56qmYj6JIASeOHlB/nTJhjuuUng3s4+Ejd
4a4K1qtgrS7cgJ2bRL6doz2xMBZhS5bu/p1mU4gMBIPlzXlC4f90NIqZQRdo6xA4nMa1adBGhVMj
PQhU9j6MkYPObY0BrDJmg4OxG9OiUOKzHGJNBpCQUTYXXRuUN92Xazq/a1yP8wLSqPN7Ino41tnu
Yf1ouEfoex4Po54EYxhTDphOQE5ys7zBBJtFDiRi6SHCgoOgOkII93ckJH5wo0yeLEI2C+WwC3sX
snJpxw8dGRtHkSoBLX0KUSXMGhGMro5rJ3RQ4AMVZuGsxoQ339Ht2/pp1gqXFdBaDLoCH6Qd0cKi
XaA8SDDJqgDhU2aQ/rNrmUyv9euLsHl3q2w5JVbLRMi6DC8zNUIAPQx1VTzq8VMA7xeLbzAkwygN
Zqj3CZA/f8uK/rm7jg0jgzW5W68B8v1BuyF1B73r7MevPtR0eH9exV4ws0I+2vnTAF7c8c1lKikr
biK9CkiZu5p/t3YAnODpZalcY0yOGf2shS18OIpqBAihgGEndWoQ5UkzhpYAHv/Ut0OdiUvPVUqX
3ECtPCvkK/cSpmVVD3f8ogULRR+uy2RIQ7ToWgVE1ducw0LDeqGqc0Oa48DAfXbJs1Fs0MJZcP2Q
VZgvBo0IeZErdmwtjiBz9kyNK7I5bsdCeMOpPfxyHWYR/jccVrXk8nxBbLqxcNS1xSuc/rAEbTf0
asYWrmEq8ieZecTyKXFp0NO4cZtcjzPXf+LO9xz7wizz0/AFefly3q20AmU95l3Zjwd1SjV6u9Pk
m0YvPEcnyxYKDf8fMMvszkSMLFp4AJocEdbzhLPxs0XaLMGS7rvHbDx4bnNWLYfiS7Mogc/J6Bo2
iRSOZ8cHSFY1cnZTCWQp3aanYS8mnoIcOaxJkfaHe4aEZlQzzR+llRdKHdKQ1jUCEXLI+O16joM9
6d61Zeg7/oua24KxsCO2bCKCUySb3/TS4+vF4tBd4wI26zAwUBEN5ptCVZ5p070zYM71bsHO3JnN
jGVZxyHMoayW5Xu26F0TTEHGcatu5CrVtUsqLxEGcv3AGwYHq/62tAOQvqZJ9eiJes/0dsJhO5Kl
dx0UZaOyzCEWBrkR+vrvhJsT5FhhJEasRjnPkxOBx8dEqHq+wkO8mS5zOc7LJX4FoN1ntmqkkXxD
LqDXZ3upgyTONUxCIF70Zkhn+qmNs6X2QdgTVxpOQLTndM43U3pipj2GJ1RRuAdjzFFv9jeHJI8n
qpHMa2pzrS7EO3a8ATdIhLj5ahBCzoc6qI/tREr6pASjiiLL2Q1J7kInZw+4jlha46vEsoC5+IRN
33aTf9c3O5zIFpwfF5GESdgOemi7NReHLy0CxL3reqquWyEVs2F0eub4pZtgspVGlqWOJ6yvkAi7
vbjVp7blFTbxFPFjP3YJnWdfKfPGTGP6ISmBI61PIx/wSftLjWMHUyZxPMnzMVZqvax8ai7a2kEL
95BtNsSY891+uYm8aIETqlbzY5kNmdyDYozYCaNoCfyVUiO0BGqloILDl+wLjfOwNsAXQ7shkTnk
qizznVJE+Ar8NG5cRDKWzN0Rb5oibf1dLg1uT0tVtaivsC4nmheoePDB9RToe0GsCPGQJHFmXm9E
Vq7bkbPYmJtlDal/uX3SD6sZifwWm8NUAny56Vx8yn+KlkHrm+iBSmK234S6jdxf9Su5NcLFAAIW
/dHjOQwIlI4lQcawcnlWk5PUnOByJQoItaPp4Ch1/IywQQRDjBGKYCH9JuYCeBeW+dBfTvPg3e8M
8SA/edILKHJtLu6GwXm40mnMNnHFGKMLzR/HRt4c+eRIk/RD74CtnjCcZv1FuoiCmR3ziFKYRNW6
SbnDSyhWphIA1mPtK7g6pXZfHmu7/VHmfj41XVKhJrsfzJlklL7e7lfRrbry0dxqaLR7BdLWw8Qj
Og9+6rsCVEQ8bJ4YqJrzcRia2zw9kv8mF1evuEbbn71SL4HUmQ4AcOOvJ4nviWbahY4XPqeAPGoF
9avTu+FOlfXtSgdCqwMK81RHrKnQY8iOXNQ9/WoBOskuV62DWlYod81c253LGuID2dAY8s0SLmtS
FLKvF4NTHX/HrAEHPEUIQi703eXtxmktzJH4DKubICyaMkjCOA1pN/Z+DfjeiXQA3ZmHSb+JIfLh
HIYb6VxUVLoU2Qo44kIudNKHOI/JOIOan8XKLfFxXoSG4at3YKeKE9nXwp+Gptsl+9LGT+Dxk+x1
7X0PDXMI+Z2I4Mce8Ad/JmA+g7Je21dFwM/AarvjaCCteWfkh48bL2DfJH/TdWCoC7+FjC2yh+DE
8qCV/fTepNt5pHcogCQU/aCv9cN98ErctrQR019XwQkbgrqJabfdETdwsy2Ddk+8C4T8x66rPjQC
yj/yjLu7jkGmbag1xVWIwCAFAei1guIm1LwKW+ThzrR90qaJh74BsHZILdpFcQLfBvMeGXlbjoLV
sli3CqY4h3Db4KOo1d6wZhA/9B0jatXp/d6JPZ9uSlj30nNmso3ADrf7xlJte8Y3f7vQ6ePywHbZ
wHBO7ERracV7KepL2+eSavfGC5cXntilbCbbAkRJq/FGas61r4NWB07xeuGaU3GSjUMBMr0QPJCq
lKZ8Ow2N+qt5lqgmwF6AGSFinbf7cXmWp5qb0g4GB+r/T9tcpeXN1+2a6fX8NJ7QjTZVomnPvRxT
Eu2wQ6GvMSQM2nbqPQ+rMqTjAYnzg3UtorgDaCI08i1+btgbv7ktH68SjETUiJBrPyWQQRqMR0EG
v+5qp3USidz5b2ZjPXG/VckO4DGG4rmjau8XOTlSc+EMzsbA867CzSpZH1BrZ2+d2gZin6ibRD9E
QEpv134huaiMqMNtjy438X8SCLNxr4ps7wXQ1fa6O+W1/WRTba8h5FDR0ty/G4Aq3I9HDWOXk79g
FGw2OzDM5+4VqxFu/SLe2pFeEOoGQNriD0HhQtMk1CIUKJefWQJniKblvyct7q68vYRqXt623DXi
oV+ebKoGGnJA8C/r50iTpRhtKyIivUtrndhCDYi6AF8xRais9AXoBhvqxiX7Z/oT80mNHPx8nU3i
twybFtFyUIEg7XheOtPZsnK/H9KOEMMfyQRE4KigGhKwnaO9H+xRcUlzgQr1HTK9+w4sV6psBSDm
oUg3ln1hKUMufrF5dPXBPL3b50+jUqW5KhtZgF3tN2ayj1/ueJIX1ACweDk5B6FEYwQVgeQxNYP1
H5847EurJDv9RqxKcy22PR+KMSbQWm1sQhNQXCCR/dWVbb94LY4q0YFcnPp4b268ybt5/IFEO8pr
SmEwujzOo68bMplX2pHPEYFvMofyP72vNjBfQKWrRCffE8b5F8EVDqsaw4o3de2Joz9XhYQVGFP3
hRg0uaD6CMkOTkyv/Hcnsyo3aNH7KEqLOc5qwc8D+Xm136eOROfHyn7Hd0kaEPclSM7XzPKDwNUv
8owOsUEP4JBFd3a0QMKvc5HrKYMqSbiAv7O/cl76x5ClTECqXNBgn+crH5y2cTlcZEP3btIBADu1
4tJQAwClnkzAWDMcTPnnuerxvsAbAsoquWd8FQj9ePt2EUUhl1Ux1gT2BhuchIBCmZouQ3Uc/fpL
Evn/p6tyQg+cWGOi7j4FlNatX3491zZnunktXCw7Fi1HgI+5d+YtNUcA3FioOEqYJYaVovyGHPBF
50fdyQYSNsHqX1S+qZiHdtJmMYa88xvQfrkAWEW8p9cFDyczEbb3GdtgV/8c7wbuZNsnS1IB47qb
fkoUIeM8BFBE6ksiHmnV1fRKZz0xZd4sYNNzx/mfNmX5JX4J9y5S7VwOt0eeSnXWEVzsHdb2GRRn
FzgBWZt2mIDq5CLwVqjSZTOUrUDfBZ16UcEuaOJRqVdIz8j6OHa8lZtecdmF8+HSdzpyAN+EiBaD
p0UH0rFaUkPFzGano/LdvzWpHKVDNG4rwme22WbORg4oSyUBzKfnSaa8fbJqPaOoa490czyf3Xdy
Jk7HXiadGRkU+qBpLmC9jaKs7ZMvu4oOJ1gl3pfmcJmEO35+1pVmsFgQTWNqnPFYieSb3h0qNBKT
c/0NXglwWHxStVF7QTBoD37YKc7JFGKu3GJvqYWSvIJ2Tc/MWyxo2p+6eWAWCGplgirujxN40zQF
M0GKHmXdvS8vpUiW4f/3SnfVZLN3Eut5jaEyYuxBbSjYt1nL7wJbKo8NFvNLxGtEWyI51jNXD3+w
/DEuK3OZP4ya28mh7B9aYIx3cbp/DTiqfr+OExJQ9a+FyF1zixB77xugq2XLfRDhHlDBq28bbCiP
gYt9FlvFX/TsAmXHQlEOPryhcpgKGANB+VBkqoVjKOVzFc5I+CIN/CSdUcoRbggYk0n+L1Qpo58o
GZO9HOKhfiwoBvn8Pd1D9XHdgC3K/iFBOkWMjvjLGR2aGAXhGnDqtmakcZTEJEI4JPhpccjIMFGT
33SsIIXnJ1A1A9y5TP7E96dJVA+N7pH43vp3hOIo/0CSadJPE2JoZKXLIHRH8DBhUYm0H6JM3oC2
4Qt8n+0ZMa4ADy4HtalL288I4cX+Gei5xAqNCTO4NY0ioTVexn43bCLMhVyw/pn+A4Eqxi0NOPm1
Ra4qi9l4hfRatB24KKExaIyqXcUEsvftZZuSjAd7IALsqv0PkLlbuc21H7hvHUKv5LjnWTNnTXw3
134s291W0ZF1fCPeBjVkVB8fSS+Evh1iA3B7Vu+AsXoeHWI96CdTgg/0LBmrwBARI9eKwG/zC2Kj
jPsGULTsfnJgZiJtcaGT7Y+Jxe8EKns7wMnC0K3hwGnIbC4afzwY117Kvn0OsNI6cvwJtT5l32dc
+tPVaK/kn57OMBp7pY4tG7TPnkxtlffGX64NDhnSLBnvW+DNxm/KHma/mewxlN4GY7gP9Hoy6LqF
j9+l12+JWoXjLO6NW0w8WBRylJiG8IX12hEPdrhaJ/H4cQtSsu/h9bPYYYBSYQXpQ4j9ISSu83oy
IgkTzCL0ccGMAN+3zK0TxvtlG9/WAo3D3j/ac1DTPlJiShiNcFFDEkoUqBzMJEEpXUrCS5lncHJN
hsR87RoqAr2FiRUDoJEeIgn3AbqLGlwm0jONInAs4SptfKqt8zHFYCE61J6Vyz4RDUwhLNDl0XSE
I5XgbRpQW0kZTjEPM/6pEseUxDj2emwme6Va0kRD+OcfqJMrYRBIsXqZXqs+0VpYcydTFDTmy75u
ROsXf+TzRAiu30gIVaXR4j7j7akankZKN0MmX9M7RDd9soNer+Ekb+WOjzZfm35xFkoFaU8N/GPO
FjxCJEvnb84pojI2wct4G468OznxnRUKPYrlz6aXftCcdREnI4bX+MXIVRRhBAUH1ens1Pp/ejDs
DOoeYvZFDZNVI2pbPbOZZtnVcASFh8jP9r5jA1hiO4cfeubfnaWFVjRjxDMazCpLAR/O902lkT3V
UZXXmEP2amNu/yWmruORbtKbqekL4G/WWsaWR6uGfrY6VqZ/5dKe/S3szEXjLsRDeVpq1/w+rFbv
kpHjnZm8okSDDSpV7A8YQLfDuMVxommitdvKOz2KWRKo1yuT9G7BFx8BXjDj3UA4B/7MQ8wQBxO4
pUlhIOzVCS6kOSivNKWJGV7DsqNJ0bvDentgZjt3KTUMWTyR6CsPiul4ppF5eC/kQv/lu7/gnv0M
l8aFa8pwiMq8c+vWfpEx1ZZP0Y2KU7E9FZE0y6J2j8FGJNO6R0PbvDbXyNHdcKlhX2tuFAvBXSDG
ir5ExUrH9qHuVaMkOZoREndRVwYVQUQjovD74J3kvaicgBY0f4qWd5Qi2Ra4OCbhtmmCPuZldykk
ca+gMQxsS3w1eORHhTvVhG7qH5cb2Ryhwry57GKz0HFdoCeheq4w9ShJ7HkcSDKqXRwbsQ/D8wyC
FWmh6ExcElKKjXGrlqRuvNv48vpKj7ncWKQpiZ6bBijif1/Tk64N36bYjHebUE2Qnu33VnnGfAG3
zQ4v6LLf+SPyaO1cmUI7JF4pYJIlm0+A3AKYW4WhXU6GKqjvX9I6UIVQA2XQUvtwG4gDudRteWif
JbaKpSxfEo4BkK92aBL7W8PwziF5+HXsOc73SYvmLIoeZLHHfvyj1u10Ex/gOguu0lTw61bRYU9Z
oMVQ1osRG2Lwn9GQ1SbuuQesS6AL3WzzlHm3gg5pk7yGirAqHzkG7sJCmEIaDVxRdfmoncKQj4sT
afCCtf5pECoyUkaWxmsUY+7DuwcFTVDiJr/mUTX3afp3VosAMH0JNJcKrRqrt4E3CGpuFHxM0Pns
fxgdPMFJOEoQtqaArxr8EnK4kjDAP+2Gtrk5Plf6poJJF+0/l32R21erBdcidhlM+X/cFRqr3anS
XmyLrCqf7ESbCwnm92UCBrrCFggn6nT+Grle5eNxC1DwV9Wlh0u0FYZVtfDIUMED0UuAzYJ3LfAG
haYdmS4fZQ1rXN7w6Q9Ip1j+/rkfwGSulAXxg/U7wyEfmozzVF7Ee1lnkQn5xIGyDCMzZ+BZGz/P
j5k7qCa2rTv/e4N5fx2+gbuamoNc0PI7HurSA5Y4GFeO1A78wGM/g1F2Zm0x5DU1H7T79PNGceg7
jMgsh2H9Dft0dRQ8iSNDBAeoJy2JfosxRyD9QLy6/MVSFf40y4Iwy/zXHmF8NEfzn02gb9vyq59r
hfI1LJqQ1AHfIQ+/J+bem4nXQKsOR3mdesq1EA30wgoxAIndF8DNLuuoFyV2t8SksGzIkJgeflhE
JXB4MxCp/46aH+DifLbdF3LRmClsz4JvRK91SyJcbq7fVtDnTMtKzCbH3ZKCQ6tQBBGsjIhRXogx
GFZn8JfyI0FTC2RspUC3/NxDtRMTuQeU853qgQGFFYdqaSPG/0huP2Ytfg008ZefyR6dYW9wZhRd
mz9icvN07J+7VVaSSGKOAwlKzufKo84lQbhiKsbm0WcwUz6TN5s5QN9v6VEzN8t+2Jw0KX6uv5K7
cPMobM8+eKPp47lr8SQ2xYRRrYJmO/tAN7buUMfG3Yq18PXpIbzsGga49dHiBne5TDgl2nYXA4b5
ktSiKJ4xGChufe0i24RlkscFV8HlEoFIPzfZx6EgTRXVAbQ0q3kzgtWJR0DCbmxIgaGX3S6+uozu
jYS0uKJKcNPTUxhpDAoeE3wJW6XLnsK/rzC8UYte6aSERn7ZBNJBKPWCl5fzGiHTWUZLw1eWVYZr
qf1nZx7rfz8ol+hRfuP4bbeAWoGhYmlBM9g1h38xfyWSu4yJvkWzJj8PinhWyAiJtwP5fl5kteyC
FGDn79Fx4JWpMcusrpbQ3CycPdAl8xQDrD8y0z6QhVYD/xrM8hAwgakbGEsdWaw=
`protect end_protected
