XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����*BcW��M" ��e�~���op1	���.��'��`�<�4ጆڲ�-���uJ�X��uX��`3�C�3ݠh����^�������*�9� ���\�Zo��ݕ���*\��r6��
o0+3.$��/� S��*��a�5Y��~i����n���Z������f�a�1$�^��'0,�CB���)|���	/Qb�ς3U�)�$� t7�ޞ���s����X i~߃	��ECNh�_�{Փ�p��v�n���Ư����w�=�;��
�b7#8�����z�n#��4V=ztj	A�q�	����`P�XG�H�hރ���i��0���� � �ﱕ���9�$g�����3.B���m� u ��s���p�L��Q�ۯc�)�)�6ۨ'8d�6�/6ǣ~���ܨ�.����L���:�¨�Y��4G����e�o�ρ8�p� �ij��)d�_OI�unWEdN1�O.P�;V��z0+����#��]�����7"�'�*���.�I	�2r�G���ȿ�9+�m�e� � �ݙT�* ���g�@��tC.{/�4�Bx����Cv�l�J�o�-��OX)�ݏBJ���:�d���7zW�
�7���@RbJFC2̥5��xoF�{C5�[�^+3�l'\��'i!�H3����̘H���]���W^�.t�����Ez�2(�yl�94�U��@hbC��7ڢ�n�s�1���XlxVHYEB     400     240B[]ه:��҃ޫT��mm�4K�{�~AN 6�n[X�ʎ�fN��F�����a�{�1�7oi�#YXU�AI���G�h��ڝ�Ε����v�c}#tYS�>�*��H��J4a�����t�[0��)���$@ij�}�p�����K�EJQ��_D@�
��$<->�f�F'���+w�7���Rhjz�Al�\h:@4����*g
�s������r�$�> j��qg@x��%��Bu|�{*�?d���{�6���/e|^�M�����Z�j�:��Y)���*5=Tر��ÌAzt-��물���d���mC�96��`�O�i��ί�*���y�����!vm<>c�N��1 �8(�j��3�o�<��G�m����+�������)�[g�լS�����| ��l����R&⬐��;h(i_���6�s��擘�������~%�(qQd�����I�C��.�?h}��\ݪڧ&S��au5S�K(Q�=ʚ�����w`��p��Q��-�ST�m� Q�t��o�4�`>g�(�F~�I���U�ȷ�XlxVHYEB     400     210Xp."lӞ��s?TG�0H��()"�����3>
���^��QC=4b؞�-7孞;o�_����2L��V�G�޾�m�y��Z�X~�Ȝ����X��kS�rB���\���K�8�yv����A���ܲg	�X0��Q�f�tn�0�;�j3�v���f���uFt�<�l������d���g�?�o����(�r9Z���yS)Mi� ���'g%ԍo�&�Sy���	"�p�\?,g�na�*��`0�<�|��;R�^0!�zHQ�Ǉ�]"��x^cۓ���]�v�{��AAE��2l)�K���]W���j9�%���$�^L���H��2(�$슎4�f��<%$�JEL���tj���B�N��@����X�qS��fd�\���L咮�*r�hW�~�\V�9bd�oY��r�k��(��J�,k$��`�}�����HX:���W,+�*�������)~/�H��c��ǄI�:m�����G2��4�ݜ -[�ภ�8�+��b<��:XlxVHYEB     400     1f0�pԂ&;h�N!���'�j?,�@��;w���1����y�3�g+�LWD�;�B� X�,��M�}h�\�	J��8��3JF~d!/�ϰ����k8��D������M�m���,Gc-�;�8��>B�X����놽KW.4�HX+3?U
y��u*<��2��FI�k_,��[����z���p�[ۗ%w0����+\���e�ԗ�akZ�
�c��h��M���œvǿ� ��ͬ�72Y<����W�^0��F�S׀\l��	jD�m��ׅDgĢp��/�#�Ɩ��8�΢�S1G��F��ϳ��T{�Zu�A�Q�̛^#���q}��|����#��Pl?�0�c͐"�Zn�~�|	"8�M�j=��$}M��G�8|���A+^����D8+�{���-�,vߓ0�فu�eaܿ}��/=Uzۭ���Zs]�
��67��"�i:+���������ՈoH���_���	��B]��r�����XlxVHYEB     400     1c0Wm��2N�?\�ӹw^�d�a�1��1A*��h���}|����=�9���W��S���E�N/���$�<c�;HW�d�H�4؉�'��u'����s*�O�\0X�c+����p��JI�?�`	�y�g�p����h颵,�\K`�{D�:K\��tT��>ܸ��-��I�Ý3�!N���x�l5���=C��n�Z[��n�е�d�}bVh׸]5�p�K���!��#����jY���k��y���5y���Z��˸(	5��jH���u����$S}b��U�ve�������?s����m8L�L*o�2�+aO�,���ʏ<��R���������qFE��Π=Y��r ]���g�u�+ ,0�a2
.��~>�##hӠ?�.�Xn�{#|p�1wW���IT�FJ&�����K�x���ɱ����j�}����uXlxVHYEB     400     200�Z��\�%�6�an�T����YX��N�h��� �J
�f |{9��}�u�\*E��t�ȉ�p|�/���mw�͹6�EpH�kÙ��4���F����}uZ���[ۇB:�������U��|�u�����(�ꊻ@�[�Nג�`�o��҆wBl�k�@�^�S�]�����c��05��n��аv�*���P� ��h��1aב�+a$�	�L�Y�(���US���5U���]Y��x_G�[��+j���9c��|�i㗶�]1ִ��y�}!�}������<V+Lt6���C1w9�@����_��Q4��~d�Ym�H���?�B�!O�"56,@�#�I�aц11��D,.�S�x�p�ܴ���#����e�'��P���l���h���iK`#3��c5c#���ӳ�'E��5� R��i��_|`��4�$(|!�ʯ��Q����Du�<o�5)����s���`^�`�b5Ʈ`��0�sXlxVHYEB     400     120E��_-�:<ws�	�%�E:�j�Db�Ѥ1��}"�-������*rEp�gr�d9Xnf�<�;�I�闌��r�	D؎�j9"�ŋ(�	~����[�QM��Ά���J���t\w����4��y��w����p늏�oީz=�AH=��f�3v,�7�"k�dH�y�>����v�p�a��H�T
w�3�}A.�<�U��C� U�:�DB���\q��I1o�+�8���X_��1\n�Z��i�<ř8X�O��W-$49��%wjJ�w��XlxVHYEB     400     1a0h&�H��l�������h����O^���@L�`���Ț��g�"F������_�O�Y�ΓO�kY�wX\���9E�y�,4���vSqBqo��,`�9-�?���*mf��2k����sG,��)���9�u^��I��C�wr\D�.C�R��{�ކ��WC���ǌ0j��`蠒9Hs�ȥ�YZ��B��0�u���K��D��zvƙ�~ڏ.u�^���B:�Ւ�8�°��B�yͣ������t ��輣��w��?`���ܧ�'�;�>�R̴tD�p�MP�.IW����	�� 4���t�75|��-�)@}�[�
+��4����#(�4��@K�h�)�;��T�7a)�XST�-�2,?mF%�3��:�����K;��ƣ��k��׽��S�����ٻT���a�U�.�XlxVHYEB     400     110�%�t���L��^��>���A���z����5 8.^Vm��֗l��U���ab���cų�[q�	�0�$	�"��z�tu�X�BP�[��ӵN#�!F9`h3�S*l����XJ'��S�wLK�l�'
hY�b���#I��d>[eծ?��M��!��ietx��)3)
�d�<�X=?�~�t�	�z%�� �����(����{���G뱬����A��9��C��̃,��)u�wG6i�^}:��'�N�>��_���Ot��zKFLXlxVHYEB     400      f0Cu���1W�"	 �
ƛ�p(n�����d}��z��Y�z�.-��GЇ����(P�z����9uU�{��7���M�V�W��,�ք���Am �Fw���w9"�d%�ΡF�\k��ky�ꚫyq2���Y�rN�.)6�3�/���?�W�H�a�u�+1��3�6@�1A�GG3�HZ;.ŧ���	��e�ʹ��J��@Իv3���s�%e9�^�:@��a���E��%�Q��\XlxVHYEB     400     130%?{OP�19'�'��A�qR��d�����+[����A�sEd�ݏ�f7���_5H���?X	�5��(�1"�>o�\�Ŗ{����!�ԫb&R$�\�¨�ReC$���#����V{�k3E�/l�:�G��sE;h+� 1!ت�U�y���d��/�����U�TXۓ����P�ꤍ���Tͪ���Py>6
(7Di�i8�������� �π�@h��N�(�oy��9���⳽ӑ��M��-����[
�+�jv����x�Hi�u�*i�	+��m_�)������*�A_1��969XlxVHYEB     400     130K���ӓ�����l�a�9���,)�E�08�`���tz�-�]Nty����g�c��B�o���{n.���<A�D�@Bfe�r�v&�J@�F`�ObŐɕ/���x��؝{ﵢ6n��V�9d}��c< �n�.�E��~NF�\N��*�<�ip�VAg+�T�j��Nj��V"b{���a4��Vk[����!B(������J�)��X�)��u��w��'))�%��Z.��1'W�C�TnQ�#���f��y'],���:�IP;�.P���H�������[�w�l�6�XlxVHYEB     400     130�k��s�ŉ�T�Q>Q�b��IO��i4;{Cy��T��s��;�r/L�-������ӡ���J��y���L��_fO�>n2/ʄ"�p�Gv��gҫ��r'n�m��9|Aubi�kP.��MM����;pA�K�s�$���B�Y"� �w#�2;ϐ�[QM����I��Z�OJ�u�a��i[t��de0���C��w��'��6�]��*_|�����Fq�#A�8�-�D��t��HW�*>��>2���Ť�5B.�Q*A����䬋Tw9�N�k`�����}���XlxVHYEB     400     190�m!1d��+�A=m3:@a�ap�Gx��f ���ςG�㐟S����p�m�T�:~��b�J,�=p��7����?�<���H����0��՛��!��"��@�R��\��_����T��@�2άϭ�`��薫p�~�z��i��ke�d��9� ��n+�~��l�d�����!�j�D�&z����v��iAM	߃{n%��"Y���-�4I��P%Pn3)���a\��0�H�EU�{E�,�@�#�T(�"�!�.��&SQ"�}8�`���n� SOd�M��1-��)��Z�H��(a2�Շٴ����B��.2>�)��/x�	1�3����:r���Ɉ"P�[ZC�X�I}�6M�/��^U �d��ҙ��U�q��0�AXlxVHYEB     400     110��۽+_	��gA�7{�mdY�M���&� g������Ӥ�@���apqg�;�m�5Xl֡XM�؁��G��5:#xT��z�y�"1+f���TD�0-���d\��fa}�Yf�n�I
����m�sH�^�Ϯ8LX�������P�X����ԱB����-Z����j a�=�5Ԩ���k���;�d����<<1�ߛ�c�10��Ǎ�)���yU>ϗ�����V��Pp/g���h|P�A2��&@<����oi��'���~ؼXlxVHYEB     400     1b0�?i��[�9G[����ʹ���OI��ܐ�j�˄\L%�S0�A|�<���J
q�4��\d4��^8��]}A�OÌ]Jb�w+�k6��:5u'lm,~�k�g�Ru�:�,HRp�R��ڬ��]����zh)�s񢤓�h�����߬p�P�n�0�d��4��/�o��uQJ�����B�M��tA�%�PRm�1Z`���&(�}��m��8�S���=�f-@L��P�s�zD�9�7�L��W�c93��Sn_"�#�Q���Q0i]�8�>��g����46�4���*$L���D��]"W���L��Dp����AUk��GMJ~��#�"�FtV��o?�g���?|X�[kZh�+�a��b1�Z%�<�1 ��+�@l�Fy����k�	�i@�1mz�Hcm��戆Y�XlxVHYEB     400     190yB$�`��˪z(ۣ�%݀���s�=����~ �%�l��1�!����=�I�����ֻLѻ�������?��p,F��y=�u�B�c;�f~j��y�ds��@T$�9�ã�^�U�����SG��GmTL�W�m��pY�[.����^�7���ŴB�"�����2K X��D���j���g+�-ap�b>��<��ͭ�FO,��r�>BA���G�Vq��X2H�g�-#3���e���w�b�t�.�c���������?�� ��M�-%�@��ܾ���`�u�����2)C.4g�@��(jgfA��WSB�N�"�Є��;��/���Z�f��Ԥ�p֥��*D�r\���p�2JȺ���:�jŏ<I0�${�y�XlxVHYEB     400     120�������p�ZĆ���r�w�v�"AC �������3��b��=��p�6ꡣ�w�������MC��� ��O87�px65��'�j�ѿGb� �OH��BY�Ə	D��yr��H��K�'�����xv:��i6��2�6&e����+�Z��g�R����``����EM[�K��K����C�|(rȭG����p��q<Pt��r��[��Sh�ޘ��%�\{
	`�gz�E"|,Nٞ\铭��(W�I���@����]	ZJ��|�������R�I��k)s�%��o��>XlxVHYEB     400     120⸺�T��"Ϩ1)���h��Y8��n�_�q�1X���rj�
R��\�#��!7z�i2�&�c�KO@
� E��f)z�V0���u��������M��׾��W���nY���7x
|`��*]�FuY䑒�9��)�&>��
����a��Yc�6vQ����Ь\��+�2$��b0�73�ա�S��G+�iub�� J3n��s<F�@��WO�������E��Ԃ4��̪��uܣ�Ub3Q'�%� P�~���}!T���W�3�gt��Mi�XlxVHYEB     400     160������3�1��k��"��7x���P�ۋ`��\3\�3}?ǭ���~u�Z�ɶ�����W�}��&�}�1�y^[�dOI�7���&x�[�TP�Z;DA��8-@��&9� M��Z%��fiw�_��&��{�1U�S4�Յ��p��2^��wK�-�e�l<�]��9��I��.��ʺB�����Y�ѹ�'���&*دn�޻���ɐFR������u:�E]�fw#��ª�=�H �Y�_�@w 7
Y;+k�h�`�F��9-�>޲�ֿ��������z���U�S4/�SM��P�M�G�9�c\�Ͼ֒�<p,�����8�-���XlxVHYEB     400     150��SbD�\�dp<�u禫��bV�$��Ϫ3�vT�X6w�!-=Ό`�����d�\V�a��H:g]<Cm��)�"�yI5�8Q��r6H�:(L��0�o͏5���]��AR;~;�!���lߜ֪�G����t����ɣ��P.G��	4�IGQ�Q�G�J��[)~�;@�7B�&7șA!s�����;�lTZԅ�N�[���>�G�����e��]�F��M�2�L&�nT8�A�Z�C��;�%Ͳְ����2���0��]�d���[�d]��g÷���Y�����z�����j'eC�R׸�#��Y�|���5G�>�3�eʔXlxVHYEB     400      e0�D>�آ"���L8F�u�w�_�No�Lz<]fS��A�m\w��3��ӝC#c���7Y�)��T�@E�`^����><V'�d�)UKYk�d��_Ů"Ⱦe+}����r��Z���M�4�=�!w���;���蚉�vb�iPv��q.{:ΐ�]q@�a���3x�YUH�@P���7�y��ʤ�����p�}��wh|N�2<\p����C�XlxVHYEB     400     130�`��	�t�"yĐ[,��K!��PW��~T��-h*���sI��v{�r�y�����5Q� �(����⌺Bm��t�r�;!�<����Z�> �}��-�e�m+�W�,<�����+���֤@�o���v��Ѕ�LX&Tb�R���0
:wI�O��Fi�l���;?��W�A���R��aJyb�)����VgcF�y�Q��5,�n_�&6wc471�[���6����7��Ai��K�??֚q���LһS�i�}Ŧ	����b{~E�3�������=cT��D'T�XlxVHYEB     400     140�ך���c
���=����|�V��-�t��� y�P~���߃�]=��'5yH�d�$���[0+��W�������(h��4�Fq�0�>�Ý��8�� lFV .��b�m���}�����Ҫk��4T��Q,/G�3�;��㭤M!牅�ՁV���,Ӏ�p�ޚ	v��"���m�����0� ��;����>P!����ѐ�}q����J�,�[C�8Ô��u�:8C�3~6O/ü/_����E���6�K�nM���l���3߁D��EJ�a�M&V��ح3��-C.��J��q���OXlxVHYEB     400     150�V��X"� >]6��~�rIĸf�Y>�g|K�Z໮�}�t!d�'9L~+�OfGީ���[z�˹`=�h�k����f]q�琠w��R��;q̰�h��&6g��X��O=lY��X6{u�B0>��<���żƼ�%���|�_Ĕ��l5�`�P�:�N'@�R����[���f�X�����ܣ��{+zax2�,��(d���:L�O�츘�jiq[i��ʝK�{;�n��X5R�M77�:̹����t.Yk���4�Cs?��D{p �\;�.ѱvBzw1�G}it�v������x�wA�g
���/h/A�8�Ã���c �P��XlxVHYEB     400     150��x����Iu
�|e/�4�\��nZ��t�7����Ufv0k9<�$����>%h���Ȇ�++(S��ە:�G�����=)��o�uė�py���Mb��颚����Sz�%��9��u�_L��+���F��q����.'�/B!ԘI?�~֌ZB>=��w1�JRg>6YJQ%
��Jn���aP���^�����<��Ǻԭ���+��	��Q#]Z�]A�s�w�<��W�����AB7� �7�\Fb!��r&h���:t ��^�\<V��v?�;���YU���G��O� ����o�W�yB(��hfr}��� ��*i�_���8uXlxVHYEB     400     120�|^,j�t�����`̪�kyv��AS�`\^@�aE���u׭iy���=']��hUb,:p�H���׶W�������̂�7�,���u��k�51�t-=S�C�$Qxҍ)�p��W¥�iu�p��yp��=?W��]�F��+K14��ud�;q��đc�*O�ޝ��� �A������3U�z�L� ��M�OL&{&��Ei��b�a�x�_s'A�0��b�LZl�$���������I���L�m�
yn�Q��~�۴^�#XlxVHYEB     400     130XB7�Fk��^P���r�����9'���ᙬ#�)��x���G������0Of$3�<uŲf�����@i`�!Ͷ���T�N(��8��	��}�\h.a
��!�,M���P�F��������*(G\2�\�=TG�P�L�Y�cc;�@(��V�Fo;�Z�9)Ó��0�ޚ���ֲ�xUq#������VܾB��!�@R5�_�+��;X�AA��Oo[y����*-�A�A����-A��7���h�u�:���	�=Zۺ�ۖ����A�.�a~�HjX�&��fZ����>"Oƀ��iXlxVHYEB     400     140��s��	8/}�ǆ)h<l�^a�	�̰��(�A5P�t�Dc٦o'�V���F�n�.�O�ų�����:�Y���,�t�J?q�yB��1�zo�ʔIw<	�m�歫�gs��Q�^q�����KhG
@"a�������԰��F�Κ@���@��U���I�x"V!?�h>���*x�ƪ#Z%:X���{���ʩ@���ڂ�W0b�2oB�X2qO
�"7��%qĒ��_@ö{�W�rz?��"�n��v�e)�___����p�<���q���K��E^�A�eR$K�"��d<}nš��D�� (XlxVHYEB     400     120��Χ���sy���9��&q"�'p��W-���hv^��ڃ��4n*��o���y���������:v]ێ<�?�����9{� Y_��iI��MX�㬤���2�S�o��I�b��ol�nf�^.���c��9���^I�Q`A\lx��M�<�-9 @�(�h�-�����\P����xDp�h���S���Fg��%����,C薋�^�� ~����#��C��������9���i_�M&
�]*?���� xZ9jhz�~1�{h���v(�&��k�XlxVHYEB     400     150��żo��YV�iV���8��Q����@]��bb$�%��O��/̲/YQE~�c�H�]�ǿ�:"�}�%�ψ�
�Q��*���}��y���\�wQXiRG���f��xIVt��ɂ�}��G�c8<��B~��e��Ja��X/8��\�2{�;��iSB\I�@�E����P���.�u���s�Hܢ�+�[���*
VZ�a\q=0��Xñ�~E���/)��Sob�����r�\l�$���{����]���o�;?e�;�b�-�/���0�<���wa����!1t�1�ހ�]֖4o6*�\S��=���X۪e�6���B�O�ܐ�o�5���XlxVHYEB     400     150#`�뀣���x�ô�㏵(�:�Y���<J�5�7�����は>@&�N ����?�ͭ�?j �O<]��C�@����K��T��*+�]U2�f0�4��¿')�^�����m�����3�h2�� f�����$����L���L/��8c���trS߶�ف�����v��zW��~�u�}��摚��ڹ.�pw:^�]��iG
nҧ���#%���B8��%�Z
@�ջ�<$�&��ɼ��۵���-�`Xc�U��w��(��i�B��c��ρ:���IU�>'޳&�Ώ'�������@�\?�"�6�4�B������+t	7XX�Ja�|{XlxVHYEB     400      c0�-���ԼMot�!t@��Eׄ�\��9�j[$EH
E�&?n|�5?�rĠ\�:�(`�dN�L4j�J���cu��EIGßqe�S��(�>o��hp��6�2��y�`��'w(h�7�b�cm0`��
�3W��*�^~�v��H=�S�dy�:�����H���uN�:��$�0����4�m�W���n��BXlxVHYEB     400      c0}�q�_���^��(XC�;��,ޙL�y��C.�so��N$�
yځPTs'���2W"��%n\rv����p�7��@�G�����i��_Sa0WZV��Doc���O�`|���m�{��͂�A�NѾ �:�����%�'\9��6(��l�`փakefIQ�~<��т��1��f{��@h��?�XlxVHYEB     400     130/����o�j���b쭍��
����%$����>?��߯�g�LI[U
|+�:��7�FjV ��~L��w)8]�<,�I(9N�b�9lӕ�W�EZ���
�+���YŠ���,�:��Z=QWz����M�هu�pR�)նa�4��6��BE���wH���777i��V�e�����I��a�)��}�kWo���àJJ�\��� �XǬ?Ը}������d���{*u@}Yظ�EBMߊ��1�m�xU��Vsd\�T!�uǒ�n�3����aKl��}��lu�ݲXlxVHYEB     400     120�m���!��acډ�O������rᵶ�Z.Đ�|���	d�sm�ܷ^�n.�aW���������z�@�}��ov��#6��Ԍ�F�,�K*����K�.��8��.��R;|*6��0P��%�W;�1�bp�̩)AF�in9��o����N��*�HMM��d��6?mT9Ջg\��h�j�/=T��O��WKJ���ʹ�-����P���j|�$�!%c����ͤ����/ŖQ�U+{��m�]��g����	N;N��D�= �I' [��-4��zcXlxVHYEB     400     100◆�|�9�uS��LK`�d%�/'>��3��u�"^J���
���h��]�5<s:�U����5R ��lG��5#$��޳䢗a�j�Gq�I1��Ai��V���9|i�^�g�u�3E�~ӞZ�[A�O��#?a*�t|�/���Qe�Q7#����i��_���I׹���2�oJ�i�1�'�i�)1 ��!����(	�.8@���-�X>�QYb���7�/�D�J<�<^��k"\�#d�V*�4�3�XlxVHYEB     400     160�%5�Ɉ��� PU�ߢj�bcV����6Yl�]�.���5X�\(_j��}�z!΍d�n���8��V��ms���yä"P�����E�He���*�~� i��9KR9�$EY`��$��9�ť�%9���r5+���#��?��vw����/[���+�y���p�Mz3j���y	(!	'�8qVٌ4�;]n��%D6�3�E����pF�PJn�](�VodN����z�@4�M�NK�[�N��F������r��,h��<븲�,i��=��]p#F�*m�/�]d�;&ʩu�����Oz!�/,�;��*:pM^�I�m�������l%�� v�ǫO���Ҩ/YXlxVHYEB     400     1c0ҐĐ�k�+���IQ_���q��O�pY�g����@c� �)�^�:�~��R@"��:t�����_v��ߢqA��Tl�Ի���o K���'&gdĿTg�59ut�~^PO�*r$?-���=%��k];�`���'K�����(o͆.��v_�$g���|��O�	�R�Q<�J�׸Y�(є<-$���DH�̰�Oe�9x�n�����/4����\&�끘�����)�xH���a��	�/�?+���O�U��$�q�&��b~⑯�ƅwl炴��T�g �1�U�h:��vfٱ���3~so>��<����Z�����*K��y�(��Pc�c_d����<�m`��1�W��q��M(��0տ=�E~Wa挊�h�NU.>a]�A��e#�b���KT�t�փU�S%�L5;���Y�jM�\�ho�=XlxVHYEB     400     1d0B��9��\��f^�fǒT�S�?��.S8���Y���6(SwY��Z�W�{�c�t]�h�5R})��#NW��A/~H�:쿻	b����?�0`>�P�gv}
��>���^`m2BGx�ٗ�PW����uq��\L-�£�wU	�l=��.�5$'הS��U���:�gD)�MIϗ�W�R[t�7��:a�h�� G�L�r<�ݺ����$�ԉӓȣObs6o(�����3#��$	l7�Z��h�i�������f��k���D�s�`D�#���1T9�Z�xvs�+���b����k@��ZEw�;]@S1a7�_�
CǑ�t�o/u�d�8�n��n����D�͹����l׼�t�]-����GK�ŗ�vw��qkq5&ҍH/��ݼFu�f�AϷ�^� ]
���*h���X4�ڍ���!_���c���ѡ5�0���{!q+�l��,v�5j_��<��iXlxVHYEB     400     1b0��u�C,����q8�A�m�._�F��( H2������<�n��$�L�E��pN�p���g�r��Y�s��j\�d��<� N8�^@\�j�����.���R�����w$Z�� �����ZV �_]]���O�߾g�;ݱt���!��Bہ��w��m���:4���F�%�� m�L���mƜku��\(�k�n��|U�'H[W���+�`˒#�Bu��� �S	�-�?�|�AP	z*%�Օ�n�)B%�s���N�q^t�uy/0�V���gA��(���kA3�x�����O�|�q����_]�1��I4����8s�7�'�����A�b�T�Nbǖ�Ąs�3��jk�o�(��V5O��d��}j���B� U�`i��#l`0�?p��:%b�y􉧶�ї~	)n���q'��t�q����XlxVHYEB     400     1a0�/a�fdj��`nJ��}��u���`MӋ^>g���;���g�=�"����ĵ�J�Mz��)�S	oW�ŭ5���s��WF2�d��������D K��� Rk�߬Љ]�������� .�
ӵ�6L�Z��.�����tƽ@���j���뺓z�ip-@��<�H$h�̉�6{.�v�����͍�V��ϴ���b�A4Y�7�S��_��XP�y~�dtI@�c顭�܆�Q���˜=獹l��O<(���Q�=�i:K��^�j�n,[ϲH��l�iSq�p^�c�F��9o�2�I����Fƿ�G��c{��jCkhAbш ��p娇���z��ųO����ъ�5R��$S��!xH�[>L�*��i��6
v��5�U�(�L*�yg�l��exd�6�yM=�϶XlxVHYEB     400     160忴�&K��5�����(zs��+Sɖߒg�;�۾�jg�J�R�ۯq/�s>}�-�+[GaMY�D�6�9w��)��?��-Y�i@>p��ʖ��:F�Ӝ�^��X�S�"��g4-�b�1y{�t�
�1��Lʍ���2��=q9T(�R���7�|v��@��9H$��C*�Q;�n��;�%h�$���!ϊ�<das�5(�6�
Y��ul�Zn�m��J'�EJ�����\4O�6����s�.�Ρ5��*�L#��']����������������I:��Ǭ��rY�6�ȗ��j@q��q��o��d�h	%?�eIDd����LWƐ�u�5�r�Xūg��CXlxVHYEB     400     160��4�`�P"���V�U5��!��Q`�ޘ�T�c+�A�v��αw�����p��{o��jZ��hY2Ka���5̾E�V&��è\C�һW�
K��{K�c��)�nz[a_+I�k+ȕ�$�3H���t?����_o���#�T_>c�.�l�	��0�\���N���]7َX:�ys����UN�mU��_Q��b �IZ��N`E�����}�ۅ����(��B��7�)D��{��|���$9�C�΋Ih�$:7�%�<���@�|
ha�tƊ L):�M7=$Zu�W_��O�7�'�s��!J�<Vj�.�Ͽ��
�&��$��f��yǾ�&D*3qm�WXlxVHYEB     400     180��E0�r��&C����F����N�B�]4�v�i�Z��tM?�1������2w�i���+S���N���9�����Sx��g��F��p���x,﫥��7H��y� �]����"�{*���e����=�{�s[�u�*�!Nm7MK"s��¥�}��%Z�!}IH4�ƀ!��W*@�]����tT&M��V�/=`��}�v�ȼ���z_Dk��=rD��d0K��*r����8����%GV*�-�Hm��(�H���1J���D"�p��T�����Lup/� �R7�KJŬ���7�XtY�4�3�L�{��:k�o��y��5�L�FMM�V��������I�%q�'Q�c$�'ȥxXlxVHYEB     2ed     130�g�Y��#a�)�9��QX�H�V
��"m��.�[�ʮI����q��FM2�Z�QV�c���C��ے������wTS=��D��6��;�ɱ�F!ec�vGy���!1�W3�^�'�
̮Z�?k�S3�:�@�SσAn(��{3N�n�>���i�� ��l�&��C����=ɿe�������[k��R�S͕{�l@?�B�buG3�N{߅2���NJ&�3}m�g0�W��.��K��:�rg��]�]�i=z8�ޕ��a�.��I���O#�E�$3��