��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��а�z��+�_� ��#,n�x삢~��3�[��'�[\�g���:p�C[f'�LK��Zٮ��PIy�w�БP/�Y�����ݛ���N�Uq݊��m"Y�>#��n�t
����WW�Ib��lH9�A�k8� o1���'��д�K�J��&�%9Y)�;�`�����pr6$U^�h�N�����P����J����!?p��q�:�f��C�D��)��UPD^t�MA���Iޥ�M� ��4�� ��n�A����qI�#�riwA)Sm��T�)�|�Mf���X��J?~��}���999�����H[�2��:���<v"��(�a��ߘE�5��)���?�%*�u]9%��d�*d�S	�;�%�v߸��/���Ř+�V������N��f#�+Y������ϽĆ�M�<5'b�D��������6��-U��@Gz��%���:*7T�z8�7T.��'��n�h7댎�F�'�+@�+�<��Wa0���7?J�{q���8ӵ`��FL5�.���(�RO��v^%�<C��b�����t֗0hY�D��Q�s�����m�X1?�lx�~��[����$6Y��0�?��,T}A�J���k��(d�A5�l�n/���mZ�ȸ���a��=��;_,3�v����sT������(�,
��$H��~"_ZH�0��n�}��AZ��4q�e�պ��AOk��*ٰ�xf��! �z�LKD�)P�$�7�T����\0nb�G��i8Br_L�9�`�eK.h��Sk�d�&'����Ơ�j>�y�(w��� �ˣ R|�ΊK�y��i���L��_���zE�X;�)z�R�s���e06���<^�f�%�gN,�O}J����9�����_��Ul��[�e���`���SA�ɪp��5	B�x3��-���dL,�! #����'�Hm�[���)��CM��݋5;?�@��l�[�ka���폱e�5�է���9���{���/��_��	ǻ�Hu�������C��L[��j�'�	@K��2՘m^�QX�[˯�~WZe�mYj�h��_V/J~�3�sBAG(WB��������~���Pv�C�������-����l�8t.�!�������f&��~��+d=l�ۑ%��)����$�=CT`�,'͹q o��Ox�i؂崷0��D� ��t��,99ϯ�w�k�e;�M��_�.&K�3�;�!��!���s�$I\�0��C� M�m��9(R`T-��,t�б?�m>��b����d<<)��#��0��|;k4@g���@�F��e[S 0��s�K���O���k(��9��!��5�pZ�9�&�4�Yd���ύJ��k|)#1��z�u��ņ�6˟&̬5U�6z�7��;�夠g�{�^t�ۙR��3t��~��/q�}ҧVx�x�=ڇ�R�f�G�K�t�e.��mڟ�`�!5¡,TV�\�[&zu�l�&�x1VoUr���Xhغ�dܮ����,&��d�z:׉h�-���P����~�����^=�}Al �6�/���)��K��ln�>�F�`���ς�Ha--OX~����V=h
��{�"ػ$o�z}�|:��>5��<����"�JZH�y������,�i�dm��3m��s�
m �$m������qY�M��g��&58�^[�6-%g�ux0���3�I���<�y%���h$�W���f�*�� $�V�Н��mV����5�Y��X�	��)S�җ>Y��b�9�nb	�#f�3h\Ȧ)�S��V��� sL;���*%�=�VN��\�@+� Q�,�؄�V؇�VG��'�1�E�4����0�:ū}�J�Q���{�(��߯���3��e�͝�
�D�,�;����郼Y�C7~�޴�w�@� [�l��o�Gl= /ue(2\��!�%)6�2�m[�G� ��v�u�5�r�ǒ�h�(Y����r.j�eA�Pi$F(�"g ��` ;X���{纰$��$8��C ��4#뙆H+g�����NB3�GwG,�쿡���0c�C"G���yR��Jt��-�ח;�/%��M��!5�-(kUr��-w,��t���O�|��wQhI�v���F{v�n�L�B��}��3]��PO��׺|�C��?d��� P�h����6��	�C���T`�K{����37R�փ�N�1��Rt�L�a�k/��?UR24T�|n��j�-eL����)i��
?ۆ�,�߰J���{l�t�T�� R������r�ZE�sP�P�
H�<�qca�.%f>�Z�H�9�.S�{�#�?�`��^@��]�E���fzԊB�*	"%��#���#��ލ���#�4�� 		��gY���YM�?�:Z~U5i���� !i~}���E=*S�+lO��KQ^�ʋ��p�L��<ǚ� ��:eq��z�03��Q��o���kB�W�55U񲔛�HqZ��l:�~�&zk�x�1	'{�X���/�*� ���L1�I>�:���H)�"��5B:&I�ݑi`�{^#�����]Z��7Ơb zQ>�I�*'�+ۯi>k�2�1j�0	?IZ�b����]���#F|ڣX�g�$i^
�+Ch�$�3���@O��?���t��J�K���r��>yQ^/��y�v�>|>����q�
�G�M�'�B�:`�ٯu�{&&��o��:B�f<��+d��c��C�>���!�+�w�W��I�5� ���!��M�y���U*��:�)�4�p��aaZ;"ǅ6������+l�� 7��"�UЅ����̼bS�.�ү���������괚��zt��p+p�Nͫ�%֣0<����������8H�η�U�T��dsE���:7�jc���Q�Qw���j#�pH���RG���M���Uq[4��JRŷ�aʸnu���`ϭ7��q{�)s7	W����e퀸|��Գ�a�ϓ��%|��X�֝9��q]���o#��`RH&I2Wcq0I�EaH  i�lT 	��\��ﭞ}�'7��1⸌�����e�c�i��,P�X���r5B�i�-H��/m���ld���-�k`�O#��*�If��a<��s���H2�Ҷ�㨕9��,��I.���.ZH��G\����]���Uc9b�n�E�.E3�m5��n�WvCO��]��0g��%�}��Y���U�x^ZBv#�ah7Hn`-T���$�]��]骎�4��������:��څ�r���Z�xQwa�P��b������T3·!D��.�����n7
���R��q3n��H*�y%�b}�R����B����
e����L�%Y|���|�(�F7��F��v�k�옴�6��i�W�����$"���U���L��<��Di���Z��3 _/�#זׅ?���,��&�Td��/�[����܁B�����B��t<�wv��j���.�aU��Z|-=RWS������{;�j57�P+`6��S1|Ρԣ���}A��1�y�ڥƽ-A�Zؓa;���b�We�"��f�7��h�4��Y�+��f�@E�J���}�٦�Y;�f�);m�&�nLj�	H@�r�a�\��|W	�x��ê0i��0�ŧh-�$�@���-k�1��Ir�,sF�����P���jT�<�%~���Z7�1�/_l���u +-����$U`�}�t�o�e#�g�Lv��JX{~q��ėe���0�wPpи�&�;��?�6�M�z��q�"�|�Q�YYSqW�0[F����G�D?	N7�3�#����	�z������jJ=����X��2Ӣ���F��VQZ�c��wb5�R�h�~ɢ�sR�?���0��fEj��8�=��7�ɑ�E���mn00��˙yQ��Z�l����X��[�7c[o�Пa����ҺԞ��u�L���޺2w�W ������\�N a}��6,�c����b���S���вSz�#�4Z���?/Jd(��0Tc��/L��o{����ܘ_x;�������ae⌟��z��s��}��Up�����x{�Ј����
�_@�/i>�M>�-�����P�EV��롭�����dR��Ik�����Z/_�:65���\5����rb�bE�~���d1yeMu�8��;m޴��HLآ��3jB�Xf�脇����ⲏ,+#fV?ʼ}�Hr�}�-��䮵�W��$�����V3�(�c��5��kn�PHg��qYn,����x�\C$�;`,�օԬ�?�ᚳ���Ue��fۘz���{�0��!`�Ј2�[���L�(�쾆Q�7^QO-����K�.v���לR��]��ә>T)�8U�戱��9�@j4*r��yK��u��:��ʍ�4�6l�:�����-��=h���l1/B9�P'��WȘ+���Ǟ!d��)zꗨ/�D���l5����L��V�DCI�:���Q�����[{>�"��K��q��C)��ν>�
q{�FΜQ��.O�� ?�2�2GYx�$�F?��/I������/��j�<����{j?�����}�;p+�Dnd�@+u�t�օ������+Zg�X� e�`�9�A��x��K��+�8W"-�=~���+��P+�yαL�7ױ�33*��!<Z�2՜WpJ���i]��^�Ao�H"�`�zf�g^V���eo��� .��xX�̇<��h'�S��ů����$5Øms�+%!���5�?�%�z"��Á�9`}�=|�ks,N���l��gc
p����.��٪q���d�
?��|~;R��+�OР�R=�ʖ����
�� �d̯���G��`�f�m��ᥧ��<���.�}o���'&m4l�,L�,��Hͽ��d�0���4��2,�V��a4o'�u�缙k�v1�������B>(����`S�D��1yY)G��$'�ڌ�y���69����� 7��X���3�Fy�@�2��`w�r��xƂ�qT� ?�V�A�J���^�q�*�HwQv	s@�����N ɤ��A�e�B<Ҁ �.���o܃�ٕl���*��I3nw�∺&DMXB��dc�䅂x�'\q�S�(l��b��q'��5�f�T�K- H��x�z��t�^Gq�c?�A����Ie���d?�FQ�>c�W0'T�]��6���/m�27�����.�x�ꎝ7��n�Ԃ�*x���	,C�u��I<`�7���`���!�4:���:��cD���� �7��V�J���d�bq���#/��H	
�{��\���S�'�H�w"*)b�~��pݞ����@� �ʘ�d�k��&h��s��[h����w_ݮ"�-A �N��d��MC�!��(}t�����2"OgN�G��-A�&-�X�m�����\U�������b� �D�d��3�Ù��TcZm%�iL��oZ�m�~�.�\s�����O��E���)�O<�������
/�S�[$2%7���o	���7E��ᄉF��1]Ƌ�+r� W�4��b����#�;n���ɢ�<�1����nw
������1E<�վ����q�DZ�{3J�&���~ }�6���'V��o��Y8�& -�����q�F���:�'	GR��̤��[��	�y�����;����,���j���Ǫ$��C�4��\�d�[:ݪ�߆��
�����e;(���b����q�	_B6F� ��֭Bר���T��ĕq���çB�JV�ª�^�'Le�Abn��{)̵d̷��k��B�?'e��Kq��wC���X��
q ɽ.S�9m��ڭ�ݖu0n���XP��Ƴ�W5����=	������E��m*����qZ(ݣ�z�7����-���v�E�n�b$Z#�J�w�_\E��31G6f�9pܑxs|�H؊��� �*m#�[�&2qv�1��S����"�$�>s�ԙd廵����+���S��1:Ob��A9Xxa��e��??��.�~�(�e G��5�Yt���(�Ά�ˢDxx��-boci���l=�zЩ�:�r����T�v�r�}!��r+�C�$����0҂
�/l"q���aR�e*~����	��6�2����V�����l}7l.����d��~�#�J�r��������SY� /��q�Ě~q�7�+	,3�>�������q�k�8�\��^"7Y��+��i����ާ�;a�4G����֋���G��gq��r��:�,^�5�������C��f�:���;�}�k��5�8Dq��sC��E��7e������kN�ן�F�pu�`*�5X~��u�����/	|O�J��8�Su;�8� I�~C��*�I2=^�k_Gj\��َ1N�����Y�X���0���R4�F�܌	q��"��aH4I2��L�W�rЅ����1�EVC RNc.+�܈�R�p�[v��EM=6ˇ9�2{!f�s*�g��}�z�vI��S�g�$<ļ��S�܏�-B�<�8WQ{{�!K�ܡ�!�Uo�	H:�J>x����|t��2k�#��7�����ȁ2�j����W��>;��5���p�P��1�jw�O�-��At[��5l�~N��
 �H]�2�ql��K��0��L���E�\f��?������TtB]�{_)K�
<=�W~��7*�pVb�"b��	xF���Ϲ�Jv,h�j:1c�p
�%
�$)��ME:����t��
a�9|���)��wI�g>ZaM�?�ZB�ly)楑|�N��v����cp6u�+-�"�-��{ ��׭eL�3:��<Ap�i����G_�J�b�߰�ЋX/v�����5"�N�&o����1�*NI�|�ظ���wnB�e�\����mJ%�雖@:�n�_�8X��|�p�ς�i�,���a9�=ձR R.����h��|�
�� ��?9�才�P;��f7��gI�I|f�TYj��� �e��j�S܍�j�y�!h4g�Fn���u&��T��B�+��@��/�ucu���vz��=���n|���)z�G���9_���*���GjＴ(
��V�e��3�ۊq��R���R�gT{�*�� �,��X�Z0j��3�"mG5������o�E��n��U�,�B��Vgy�����~��X۷�F+�\I�i�Y%����s�oi�`�ih��a�Y�7@%'�8]f/|F6��;��n�Wм�~J��(���"�����8M�Tp�ll��Gg� ��3��W!27�K�7�	�����׵�:�:_��0������:=F;�TwAz��_!8V�kE0���7��pU�׬�¤�v�<�h���"�[���g�R){9���&�Y�Go��X{��6�Q~�q>��%�j��T$�oA+�A��YX�7���NE����P���w��n��B���9�HD	�X�o}o�vP�k'"=qv��zo�b��y�q�c�C�۰py6W?y��]�,�5����*_������';���B��&r/�tB���K�Bb�Β����D�(���u$$����������@����sPL�145�L5]�LH�H�t�{F�}�����>�RԦ_�P5r�3�@��+ѯƣ�_��$�u��A��4+��_��Q�ղ

��	��ءNXq�\K�T_Pn������HS�$�E��]n��7Ռu��[�̂��7N-`����՚���腲�e�7@/c���is��C���p.;~���Ʋau`,	~͸�[�J8w:��_�����@����%�*ђ5�����9�"ɻ��{���o���-�Dۑ���$Դ�1��d���6K@,��:�&P�������t	��e%��KpRG�,���pt����
L���X�pL��D��Q#L%��C���2�~����:	�V�8,4hi
�2d�ܰ)�Pz���"��� u/b�E�P*_Rk�E�lA��j��`������g?2����s⡜�����ɺ���?e<�Zf4�j��E�*��Р��Mf
��ǋ��]���u�+�	z�> ._�Xٖ�w D  ���w�/�������;��Jo��s)"OVnC�C�3!��|ۺs�b}�BF4�zҐLzVw��~�w�ԠLC�%w��O`�W��ty��+�W���F�c{��1\~a0V�*O���\LK��� ���ϴ%���?-��Y3{���1N�}���=�"�j�o�E��;���C��_���&p�,�%G��DK�@�Cj�̗��/⸣j�5��G3��cp����O�'�ϲ������u�|i�L%�-P��e�u�u��m�;�0ux��$�f8�Gê�u�.1�"3"4����YR�=qTm�|�V=Ó�U,�K�GHͧ`�R��\��pU��������yq��ת�Mb�ϕ/�2`T���[նA���~�ͧջHM�	��D%��U~�Vm��{��6 ���&��7�D������O6����j�B�#�(v��$�P�G�4�t�iS2'6��=�L�C�L�����}���S�ݲAGk?�9���	���cǛ�P�tѱ�E[5� �Uf�_{Uz���"��^���]�ϙ@M�c	hPie[}���6����2E� z���r�2�-x:X�����51�Ѳ,YWa�/7�.r�!��]�V	:�%(�Pf��+���;��x��θ�wu�4"����]Zօ">ӌ*2���J���A#�Y����n4�n%��9����(G�ZZ��L��z� ͓�!���dw[�{J:m��m��ܽ3M���豄��{���Oȗ�zVMM]`hH�T�y^�@��I6��"�pÑx6�!�)�B[!�$���]eo�n9����[g1�h��=��N��,�=�:hxr�)�2<E�����_�'�(�"�Y�φ���0���ڛ�y�s,�tf�|��ETu>���_9.#;8�ϔ�@
��_�l ˠ���I3�:#zW�|�R�`�� @5ȟ�s�R��GX~�A�3|�$п�1Ky⑋��m�6u�~Bϯ5j+��,�w��x�)W�����R2+�ߡ�W��"� �O�b�5� ј�\̺�!*<^��J8�E�k|c�%����RM����C�w_��פ���Y�Yy�9��AJ�����+q���(TY
���Ԁaό��d��/!X�N�&�hVCpP0W�$�>ـYg����b�2D�X��i�w�p��p�wڐ:��ns�)��-`���������7~o�841��-g ^��	�2Y�:�R�J$�ƺE����'�K(��b���.��_��M/��<B��$����U��2S�H�־̔��l:�\�{>�G4ݗu G#�#�4Sʑz�C1?�S(H�Ó�S#:���Qѕ�Ē\j�fZ�/�T1�"}�P,n1B�ߚ�h7���Rv_c��^��vw��L�������k/�r�u�h��y�LW�������]k�F�v���dFK�ԅ[�o%EJmA4�Z��=�Cv�P�yO�Y`�9�� ����Q������J�ʏ�*���l|>p��C+*�nʨ��k��>teʞ�� �z�^��{�t�ך�9�=J��BKN�����C~�h��X��t,�1�m��"�>�"g�[2Z?�����^�����q�h�I�M�I�]�����Գ�W��ox�u�����তN��8��Y�_��\�gz�;[p�Qj��!J�ٷ��p͎�Ɛ#�
�[���`1�a�M��2���LEM��`���B�86}P��*�vT���'�#6�d���(m����sZY4pG\�
�mã�wy|�1�/��Ka�C˷�T%N�P� ͔\�������L툍�[��	�p~��_�fB7Y���rR���0."��.���.���p�r�B���;�炠��O�/�)��4� .a�t&��ե�����j���ň����:���G���<X�N���3d@)}-����f���1"�h�JRv�`GA7�ig'T��L�Ĺ��7pH�>�@������ܗ���4EX�� �P�X�VRpb%�o���0R��F�:�+���i�?U�`�(���Y��{�0�.�r��4x8���ر�-��#�گr�t��ZM/ԥD�\G����>���A�R��W�����0e��f��cM0���:���X����"�
ڮ1�{|^��:�����#�^�%b�f ���^��}�Tf�SoZ��m�ѵ�Z�đ��/�R�:��Ae�z���ey3c*}���g�����ҧة���]�?�@�K�f[�=0X�)a*�V+cR� ���I�s������66Ր�h,��U���¿�����{<!�#��e?j�,�ʳ�Kyy�NËB�@��
tpLk%�C�`	=�NfO�L���,�����E�
ĉ@+��xlAF���*M�D���@��[��k�����A��S�`8��������X�I��A/��èN1XN�ҫ�fh���J�L�֢�bh͟�}�6Ncl�a"|8�01�ep��@��֯<f��-%�}l(!�.O��zvh�ت�:lq�uڜ����	�w�$��t�����ஜ;j��i�SP���,�y�=gLVi�ݸ�qC��d��*+>aʐY����B��n�A@u���e�E���
C��B�!~(G_�:�f}�?@��쵂�w�!_Seq�������n�*��7�t�Xӽ���� �`�ѳ��\�$�L����7w�º%
#�1�l�we��+nF��D��Ɉ誄��m|�ڒŔ�
��KR"#�4���Z�Ϯ�g*U�M_�KS�v�(d���wmS�-,���kl���k��߸	ڰuk&g�OH����ַ}�B>��Z6߷$�y����
W�m�m��2K�UB���c��ûۜ��߂�*��%��	�P�}�����W��㿡8w�-��=�����8?�y���;#�웠 ��Q�]d��0B�6�ߴ���ILV5�7�!&�~Ў֭=a�~[]`x�k�%��c�ED��	k'4+����X�}3:�L~�Rս^+ꓭ��p��wߣoV1Ǯu�"�1b	�P�����w��T��Iq�I����2�[�C+3E��m��D�����3(h��w��e�>L^r�v6�R�5�U[�o�|��+��|�`0��d{q�>�_*A&̂i��8�.�NJ�J-��%�Β
�F��Č�8]���u�.�7_����"���.���jJ�
�D���}��w ��1S#�Z��1�Jl����j)�M���%��P��+o�N?fR)�uj(������
VK���1�rn���4��������ri_���O��x���J�'�^����h�B<LG�ԣݞ��`�"��9��I�S_t.�&q�S���T�GU�7���o
��s�D[�ś(�9�&�镗TS�Y����F���R=���P�i�J:v��������=���#_M�����I�l.���c_������=�=5��[�4�?�o)Ɵ�9�_�~Nf�"�G�ٍ��e7��ˬjN�n�;�b(�J>�����a��MiWlp&^o_�9d�9�J�'[�-3�bm��\{V���=�|���,��S_�?#�P��U��@�4O�ԧ#�_� `,'F����Rsv�|E94j����pj�L��K�n+>ޕP]�ŏ��I�������Nk7��d}z=&�rBW�2o_4���<$/ O��l���H��O�?�,�^�Yfs�"����w�fX*�$���a�E_��$Y�8`���&��\��@K��%�F1�׺	�퓰T��҃$=�-4�&��b �����p�d����[R�w[|hL��[rJK`?���N���hD�cL#�J���O�U�1�:��zMǣ�?[ 蔼�jRdc'�@7��삧��� �y�{&�NHu7���������Ar��Ub�n}��^lu�)�3PV>�v�N7�[�A8"�fW:��������w��/�!mBsU!�#��"�9�K�5�M�����D�H�
��0��n��U���	6�����m�q��O$-���b����jMTT%Ɇ	Ը�{W^ܴsξрZ�2�0���|�yg攱*㍔P�
�r��/�r}R��]/�z�%=���Ǧ*]�p�0�x4��Xr�EČ�HƯ�B}ŷ�`���>�*��þ�­�|���.y~-��:ʒ�mkB��w;�<��2���ef{;����C��F�v��ԩ��h1cPG�Y�
��o�1��6��!#�j[�&����P*��q�	���7�#\��K�S�xjx����M����7�
�[/o �i�n��+�W����H��a�ʱA[������
�9�=*�It=�$=�lf��r3�n�.M 1Y}��4��@���l8��,�91d7Ce-�>*��j5-������}#I�A��oQ��o�|(�e|E�-�@u��$\�z:M�s]���4�i/-�6�nxcD[�)*�K����Nuxǹ�=$����Rƌ���#�*���:_�{D����R���,M�|KE�($k�1�QT�qg� �zvVP��h3?b���͵�z��͔�v���|�<����LכZX����}�\���ʊ����Ѓέ�Xh�ϑ�9)�H&�ȡ��a"��/��/bSv!V��%��O>�IZ�8 �~�� ��q�b���`g����"T�	a��!R	M ��ç�������'��{:�颉��]������o")r�=kp��tDV�9|>������bjZ��N� WZ�B��|��y<B��\�n��xM|O?|��h��P�� ��\q���A]4�`lV�\�r�����(��V^³s��F��*P��^�uk�w�������^yRJ�wb2g�o�����{�
p�J��h��ð?�5��Sj(m`y�F��
o��^��汩�Y����ğ5����Y�X��<��.ަدG��Fυ�����Q���/T����b�4�N^,�d~��f��/�ь�u7��Cɟ�O�j.n-�b���n�wgg/��s�roִ�{n�D���7� p`{-Iyh]'�*��G~x�~l���@H�ċWQ�@@�w��Ez�"�!2�$e�Z�]�la"�Wo�j��
���&��zE��@����s�K���w�3��/�FU���hKLH��Z�fdP#��
=J����?$��Ł6��V�����y�B���ӝ}
bA����0[!������PT�n*��M�n7O�a��dF�N&�իP|Q}�3+�����?��:����������vҼLAJ�	s1������v���>������d�'"��X����V�����Ru�Β;N�{4���.DN��;+��9�h��3�p�?ϥ&k��.#ق8�K�������<�Ą�����|qC�-q�զ@TXm�s��z":�}kl�1�b@�˰��:��+�!X�����=E��Ԝ�� �pY�&�ڙ
o!Z�PXr��fC�J�/�b��z��$No�|r���3!�s�ߐ�