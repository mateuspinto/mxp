XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��A-Țn_����$9In4A.�J�]z�9SL�X��"H˝�5����2+�h�pwEa}r?K$r���8���Z��aV�xr�|�!	5��D��K�_;\�	��@ӓ���:�q��j��s(Z�]`ғ1��*�5R�F��ģ�)X�\l$����0��&].h��&��1wP
�v��z+,�CQ�:�?7�n�j
� �����3.9��<�Y�o��w#3�#ocF��4�: 8�gs�k/����(>	<�z��ٟ�EK�h@k_�玪7��Im�A���Q�۩�c�z�(�"F�d����Vw�6i��m?����ߗۆ� ��fu�[��2m>�J��r���$7`j� ['	�fk�jϫAW�+���?I��+�����;�����p���ީt̍����I.e�8���C�"���Y�-���,6їnC��~s��������:�P��ۜP��Nᘡ��s�^Q��Ο.�U��i3W�	�`	��k�dp������b�#]�0u n�`G!��������6ue�(���5���.k�̤%���D��\T��ӍFW5��1�(�ToV�KP0d
�Y���2�[��L�DJ`q��y��P_Q?ET2�S�蹷�����V��4d�d%�y��F�%QK��U��8
K��P0x^�&D1��i'¸w�wW,JO�'^n#�,נLQB�(G�K��Q��X�~^[=�$�IB�-�3�ήh�	�#�N.�Jx�H��,���Z�]�	ͼ]F�XlxVHYEB     400     1e0�8][�mq�M�д��@FeY�}L��K�@KT�G���M�i9}�աw�[�����+��O�s!mf�aں2�%���j�!ANJa�S5��Fv����o9[����� �uX�uaM#�k��XV�&T(�cS�z�iQ���ͭ7%HW�]d�=�4�S?��;�	f��m��� �nR�Ɋ[$d#S�� \&-�H؛�l�Y��0�)��f6���4�����׺b��hB#��/�����gAQ�J����9vD��ML�c����vK7L�ЯɞW��P�/a��(7(�,ר�D �(��v$�ƉX�m���$xϦ�2W7,׋?�lη��c)	��+.�I8� g.W��H[F�s�v���������^Zc$��GXI��h���c3��ƵDd�0��䐺�d!+Z��R��H��*j�#s���*P����y�o_<�0�>�ă�1���ԕ�����e��0y�Q���
"k_�XlxVHYEB     213      b0\���(�V��46֑�b?�L�;��]�<pީ�FaB�A��(5L�T�nl]���Z843�P�\&x��!%�0��oE�[��C����?+���a`�/0����[0�
�t܈c�+����O�k�ٙk<��K"�F�0A<�kQ8C���þs��
��	�(1MF]�bW(]I