XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��i�<�R��%3�_�"�Dt�1���ہu��������$k�~!p^�����[�P�L:��g��è��ùe	bcѨ�پG2C�[�����g����ϜͪQ�2��P,��2OA:X��������G�9�x�7W�
�5~E�L9�Q��^�^<��ڈ`W�ԇj��	T{���]���{W&���)%�?�|�{�uc8v/�f�FH�-7E�W�]�{�*q���J��I�Z9eY�м+��I�T	~��������V�0>�X�@�[�k�*�� �ym�=z���g��B��:��5�,�y�ﯼ�k/��N��l�I��Yv4|I�q�}�6/#����¿���YCs:{|�ɏs9 �Ν�d*A�,���бl�5:哼��nxJÊ�Y)R���<<�D�!�3UD8G��p���QUͺwy��X�ѕ#�Bz��n`����3(���R.�0q�?!$�ˉŎ��nWKBG]�����/N����^�U^&��v�ut!��9�-JvĖ�PKR�0A�)I:��u}<������T��:]�(Wh�[`���l�����/ZB�Z[�����Wt�=�lFt��E�F�����{z}	q?5�|�e����gʬ�=D@�H�&~A�J��XuJ��>��_R4&U�ܽ�������؇���Ps�?I�R�	��L�M�F����쥎 !�<�v�ߢ�!Ǧ[ԥ%:�)�81�Y)�dX�|3��Wve?7k��X�" '�/��.�J��)�m;�cs��XlxVHYEB     400     1e0��ɋT*&5��n�*�e�T���.,��X`���u�Dg���T�c��vTS@��f�ܹ\Q�R[_��"�P?y؏h�_"�U�|)�Q<qБ�����ğ&t,Ct�������
�Q_�j	�����UW����'�
�I�[�C� ��^M�5��|m�6�A^	(k�G�|�{w�Ձr�	]�gn�;V���%Crۢ������n�	�x�Ei-4�G��^ť<��rEA�F�`PN�mm]��rr�n�gfaʍ촟����Oދ�����m� ݩ?X�ȳ���;�_pvC�F<����`V��֯d W#����CrH�B�}5�'������h� �gZ�r&�Um�3�pd���"�v���}��Y��9�n�/%�#mP�vN�J�LZEZa�����av}�����z]��ٿ�@𳲸�>51�D�߇�sUͼ�a��I�k�zԝ�XlxVHYEB     400     1a0em��M�gw
"h��OX�O2.qVA9O�E����5�f2��s��s�jŏՃ�7Ѥ��ޡ��S���m�� #�K\�g���	E�����D�"��l%�}5K�o��,X�D3
_E��{�̄�I�s���Y�K��i�z�M���StR��!~NO�4!�)�?�F���gq�=l�!�g�=B���}A�9����t��YTY{NL��u�y�qkB�?�2a�@�8��@Eg"< ���kl�r\�8��"��W�֔d[)�w�*(��&��{1�A%�gY�Q�2�WGֺv�t^�mIs�Ӂw�p%��$��0�61�����T?z3�]e �#j�f�Wu�l3l�ʄ�bҩI��:=R�1��nv��&1v׸5�p��5ݔP+$�i�]�+��e�V�IȌc����gXlxVHYEB     400     130�F��9k�U,��/�[E
�DioI� x�).#	Vf-#�i��|�֨bs��X�Z��!ь�%��CK]2�q?F=�^S�"����|Ĵ&�U&t�9�)XKE����>[e�@���C"���:HωT���T,&�pď�`,k\ra�O�@��bY,� ����nZ}R���o�dɿ�R��m��$y��9{`��z��$�fʮǣ**��a�2b/�,A!G�6�n��ޟ ��2�:�sts6bfi�K��!��=!�}���Ґ��1�ג�bZ�a%s�{U�"��~�3�W!���O���Re,�o�XlxVHYEB     400     150X튯-Z����(���)�42\��{�b����j�r�q�r#�������;�cъ'0v�0���;5��SsC�e��AӤ-��ߨ�ƙ�-��xy@����M��� ��
Pʘ���H|��)~� ���9��+f�׏(�Tc�����%���臝
��<��ܡ1ǵ��O�2Ѿ}%8+כ�iH �iՌ�kHN��;���{�� �[	ݯ����o�`o~lU�>E=;O��ªZ�u^�����+��_<���i�`x�b\s�3T�����lPl�L��]K�t*����'�H��#�$J�o��I���6S����Gm�XlxVHYEB     400     1a0�y�#������Ws�H�X�A�±08�!Թ�����+ם5�v���J�sǮ��T=��'YQ��XnRQH�(K���!"�X�W��c;��v����zL�!�,�eD��|�#q!8��|�ьr�<��������8�4.�����1��Q��?��`��e�c�O{P،����R{�%��+Y>�Jj�n:��hDúݟ��3�/�>�&n�%��#����0(Ho9 �9��MQ���(��n�
�}]�����
�3�\�k�	&�E��=���K������z> �.�Lۇ����'�i��8c	���y�Mʐ� ���u`9Cp��Ϡ�,��:�;w�������Ѫ�K����MU[�h���E���6:���ٟ��(I��W�Z\`p�QXlxVHYEB     400     180(���S��t�pQ��h�ա�����_�&���s�Ty���e�/	���}�}���N�`Q��]dK�¦��H5҂��s?sl�I؀,����h�N�6�q��f�����o�b�=��P��נ�s���Zr6�����O�H����ե?��l.����f�?���:��7���.�EҌ��m4������Vܒ�%O1��Ӑw-���?n0��|o�']�:�����Z� �(���Ӣy��Y��Ʀ滝���
�/�g���w�3g��g�-}�v��\���ϳ�ږ�A��>�)�S�̖@|����
��	79�	���	�,��]�D֤۠9�v����s �$ڀ�����弪W��q�2��1�g	�tu
�XlxVHYEB     3a0     170������IAh����6�q��h��|�F��1��O�&�����	��+����OŦ؛���,��H�^�+���Z\)�N���/��v�Z)4M��/�ǚ���7�f���k1f���q"���rV�du��39��jQ��P��-�C�Ԏ�;�r%�BN��k ����6f_�̨�y�n�ȧ�W�1P���C���/ 9免��FeL�Tk!�D�}�� �I����Ű���i��КIP�����+��2E5RRv� �΅��\cj�ʓah\7z�pI��
��HLf���P6�vj�2c���&_�j��kl��4���������ڛ�z�%?B.�i������{T��
emt�u�g