`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12176)
`protect data_block
BrB3B2Zm1bhZneIdKU7cUTmS82YlKCAKd193jZtt+C4RK49I1d2wZPpGEVpsSAWjSN4108JHmZDB
TFjlZQrdpfpd+OipqZL533iiZSFeOh2NAJ+TDS9jnxw3JXNlDxgStqPCFCrIjvzBRgZbd4ZRJKsl
y7JLOea120j4P7O1FEoqEMP1Q0nzdwTygl7s0vmc7jl5fCZ3ubvyN4k2MuLUBxjnHtSWsAU7L+PQ
U4xrmk7HDKTfKyrGocfLSUZjUYBP3Zztj4USXnStZ4uK+8ga9eQ1w9PudDSSEaofBLPAiMrr00sF
WhO71Tz/dZAwmrm+xTmbiI4SdVjYw5jQl3A9OQvgM4JvmUOsW6OhudetmLfqhqMWObzUXrEdaZat
ZlUN9t3QWoZ5mS33uasCwIQO47VJw5EyRoHsTjwSUWLehGELNOwxLoYp+YCv9EC8OWsugw68+dWF
43nknSSbZU2i3awTySJip6V4F1J/Al2lBRwK/+INdxJFdCpeZv4FedDq1zaGJBj6I3IgVRllsM43
QgsXTW8RnNEeQC2XOMGUDh0Sb6ld4i1pbbXxLbcjk6LIx2e5DoC/QjGgwqBzGG4noEuhT5oFbUrl
YqPSE+ROUHzRNb2sdvcFYHpQoEEk90OVc8IjfS9GlGCQZsjM/xMPCxcZm5ic8hQyGcx8YnlDopYq
GKFTvVph5xBtTxRco/pW45HAdhHqIFMItCoZcD1x41qR/b4hZ9LDMIMP5SJyjHEv8mQRProcU+hv
qzkgoFL6gf9EEIbOXmONxxGkyuWDgTC7iEWjDfQepWPULr04I0nRpDEU3OclY9FcTfbNY8QFjDEn
ro6W2yZxdny5IhJUpdWU0AYECvUJgNUz7VzOp5PQTevxlr9tmM0rlLojBu4ugSFnbbH8CpnFWQ2U
zv4bMF74KAgoFsphB52AflKePC53wk1Vj0PiiHXbjJHSpJ/r76meTu724E+lS+75dQKtco3fyr/k
EYu0eMJhC7/a9maztBSxK08ot4d+k6bzihl0hnsXvcmVEtF9VUKYZBBbRfLGMz+07QhcRq1lgUsN
PQOPPvktlHKxu3C+JC6bkuzmQivQnpoHv+HmO/R606rn7Brhc8zFM1P033eoodOS5V/WYXwm31OS
+QudaOxgkY7tH0/jrIxFar4ITgb/Rv9LZFXyVWU7aWZ1IJgcPTtsw98fQktDfk2CCFyxJ19PBWQ6
KjNPfn38QTPGOEZ53s5HqOH6R9Fz0Wadk5PEXw8RIL+hHF9ztrI4cfM2+Qr6d1dcJIQk7XL30wIv
Dz1XLJMpySZQKgisHFUEP6T5XSkH3HsAMrt85pzBdoWWn1SN7qm3uYdXqRzfJwSz5YhAAeDSDN4L
zy39qAGfn+n9VAtdp3lYsNIUvwLY7pGehNLOfZyu66zRVqb1Gm8+0i1+bP3+ZXzFF35s6VayR36F
2l8tn2oWpIk9X0ytShojUPJFoaVuVgYI/3hjuDr7s9hcKNSUiCCSjpCHCA+a4Kwb5f6HcyiwtMUA
nUgQ9DDcQ3TtASPNgLEpj1rQqjbyqrxDQ7Nm/nRoMKx2R0w6Jbz9qsyqgkm7SnYIp0rPmxBQg8fb
BFEm6CRJV8ORRiRKnE6UrxdQsvZIcduOwWmWiW6PtcTi3H9UIxwNibPHZ+QM+lbMeagsXsPpOJQW
aj1IHZ+XSJhWzaigeHvy6yrCvPbffih66MRpbmoytokq8yVIH3JFp36bOlFLZZsUoTLGV9xrQx1H
VSDphAg3sOAnk+NZ1C8CDr1NUiXAstTB3AsoswONaIfsnqQPivmCuy825mgztvSgfvQliU1veSb/
JFE30gzeiLE2HwZZ5ejoq4f6qiYMiik/vyyoHpv5onhpv8FDmxAqJgrq9mmeibQoxmZ+x0Cx0lM6
A1jQ8QVz4GzpE465gmh0eSFpYw2Jq5wpn192/2Mb2RbIWuxlRNKu6iEUT5TZ6NREbRKhklbIO+nr
sUFNA7AAMk4295OoyBo8fn0qk3KZknoY/jTQ4kiB8726M8XbqrYRnZP/kpvthp6X+vO0XwiPut7u
lUkTqLM1FDZw74OR/ch6e7q6LFzlvjPAVyw9RpLjky8ysmTIRma9AMgKk3rzDHcPc2vsSDWfjpLd
Qbrl6r/q/rExEg4W5eXFY5s7rICb/80XF5S9/GCt2zJhhLvN3FUqD0WYP49nsaTXkZ1wwzuqAMRu
GKUeM7ibrj0AWYOzoojnEXKVqSpsHCTFN3GmxpUQSROPvb/DxcXyJpvwCW1n9V0p0Xt+AakrWrNb
bZO71OICVEXN6AVNVlMjCBw2KvdJXBeiR8r2Qd4TaUoS4O+CuokDVCMPgIHyuf94KMttHSjHTe+O
rsLTLiZPTX7YB6HrGx/c5t4yE/OEBT7y9cG4P+fiVCuDJQiL/BmfE7dOm+E+GxdBsy0oaDs5JJli
JztNokyTWGajK2iZMixrTTk9XzHMbI6XHZ1yOLfHpM11MyhCtVh3N3oFpNlpc5sxS+ECgZyfWxCt
oyvzhJc+pXbM2wF0saI0s85OBYZQ9o+w3qlN9MXRE13lZFOMBlafZtAxrgSmzFYh+0eq0RyoO0Si
dkU7d0E0FIaCdL8pmflBIG2joB33DMGycazGWYmpKl9yDaJ6q6gA5bqaG/+gBFJLJlCOus5zazWE
paDd3B63bxxwbViTCXNzOz5d+CuCbLzbq3jyWuUkrc0vDqYZy+Fo0Q1hrAQly0QOWXAtoEp+K7ay
ij+UlfSOVn4HfbGrgBWPCxv4qknIbe8jA0V5YYS59r9+O3prjYXGvO7RUiyihRgGJPikuJYa6lL8
9GewnDDPHv8Oow3WiPiwHrzmPQ6bEQGLwDQ3TCv6b9K2VHj8NQTkHBhq4XuYPPv4NDYE8cK3458w
f4Ol2YnIzJ5Bk49DyMSCk3s0KgAHGfCDsLgMQAVA3zTADi2ftP3zM56OiEUIX5cuGW8paUE2zjlA
Hal/pReRuyMQaC1eI8VWaB3CCy0BMxTnOesvRCm9fGyQx5gcce9kTQkEefwxmdjUAPRAH16xcSsb
Uxcq6T/FFUCetsnCkResQqNFC/WfNB2LitU0AG0cCUYDspIpxv0ITuLsH/sgThqMOU95x1S5I23c
6E4sZ9AlUGXGcT8vHNPdXiNavvx56VHaG8R4GcKDUgozqx58NU8JlTxBA8jnmK4ZjVkyZy4bl09T
CpWsexRv4pOkZH4nB23KS9ZfRU51tid+XeU8znclu2e3E6Q5Wi2YG3TEwUWuWjOnNeY/cdfHH+Bs
xQODSTOa5+Xxuc1eWsOf/zXwrSOSupYyJrr13UeEJkbMbQuyyluHx16akCY9fJ4lylhZZ/7p9DnX
feelMZxKkl9BiyCfMOJWuH3NDbm2hqnALgfdrt59jwFYYfKpnAYIDSSc5w1sAVAF6OogMXEY3wjH
LhwvtbaaL78XXUsPgGLnl58gseZsWdEuhO7c1Y03mLQygiMfOxn0JQMxLtnMSVv0RKv/MG/yFBdp
8aFEJmNIAf2vxL6+q15eEiWmZjb6uDrUBXpUcKMsRPIDiycbfSOu6byjEYCNJw+IfJrbiYiCwVUY
FbZOvad+aASST30NRs2LsLErvs/yEONqK1jN//okyrSxUb2yyMo9ePVZrN+tj2flW0qgJljRn/19
1OZigpb6Z9JSdooKWPUFMleL4mPhsVuSoZF+YpeG231CvomswCLVACdl0coVK+oZVs/LCoUrZawM
InOk/4G1qcoreCg+NqqDGqTWP6Wc3ZDoLSyIj5MboIljhRcc42u9pBLl/Ha4LQ0h0aquSk1SkeLp
h7sG16WXcxTIqlXzCSoB/snM4pqpmy5X39YqVpT+eUGImbaU8cSOlfHsX0Ap2WCzvVGofqc3tWHP
GwAJSEq8WQlwcjbb7vAjXjjoLCK9Xz84wuUCT4w8h1lz3ZO7WTqPE4Dy3E6tntT8XDYT2vwJ/ghg
+AHVovZmgkmSDTA8yn5U4vUQu8U4vundpGX/b65AcG64FSnW+IE+zQOajV9RefhK0ZBEyXF6Ljzm
G5jf863DNuFb4KGzRq8P6Ksss5VthT7BXWaqKIXU/eumSPYokbpGlB9frz8KbQr8tu4ViYyuIHrP
pw0ZU/vFqB9Ek/TEs1Fhadld+t+Osd0ToqgrxKMezAWx7yfFt7S1x3xXbrXVV5BUqodyrtIN3YB3
x9uPlPH+hsmhZWgzCL8nYYCM4hW1C0w93HQQ/eBvUq5virE3s9rdOukvCISnTRzzVD14DhS3gJ4P
qZsVudR0wMpQtlGeiHBb+5f9pSbkhzcBLk9xKmFEkWBviXQ+avNRn1coXEAq91E0gSHUQISLP+NO
/53LatPQ9//o4eNDCPg5wev9sFY2N/AIs5dRSml+slBTo9hJvVHjikFYA790IM6+/CDlDsJCRIMr
WMM5hhRV8B+nMSe0g7hIdh/BhwU2eJqvCb050AfRWE2nd0rJf3SE0vkxhpehSeessI0fDZiTTkY8
X5xedtLUjAScRGMst0QCIEsiuo0pzjeFiCIb0QcxdNqHfBuCUj94ulV3se+8Q3psDukw8GB0+uMY
Tn5C84izCv5m4jU/rA3Gltt+pdcsSUPKaTEV6Pkno/mrDNo9TEks/G4WS8/0r3vaeSbxCCy2Luo4
Wbfe+fh2DjPuwdkgd3w7QNcgv4VQ4dQKxEfqIEgIv5XSS4CBRhQ3B5jVbv8I5tKO4r3Fqzj73aGv
yJZpSGj59yizUtutrSzeHJQwwuqRgtlEMWFKtOyJtaWPvjw9DFgC7eSALqVUX8MuvVh3UvaWi4Dk
HDFJxWOBzda9hP7FL27FrJMNA2RWdNYA/M7eldcN52ygXQnwYVuyyAmkeudtlLDHbjDMLQgzkUPU
oT6ErUitClfmh7Rt6KlqdXYaYwZZL2WZDyanit/qH0PeF02jYM8z/YQUK3ITTJKWTlv5k3Jzi+4f
qcfpO7DBa4W4DQpWRCN8Td2VwrdvdSvv6F1RQPhHrJ6nFhM6koAnzD0Kj4hH6zINe0j4RBdJ/3NE
RJue29u3TWtFbJf6toRtfa5x7fhMqcsLkcHzyoS91b79qa3+3t0+TGNBJvPia61oxdtetWGp9dUb
Bp2s3Ef/uvLqscI3aWa8v5jGSEfCX36hh95jU2/0hcJmnLTh3mW9UJ9cKQAWJJ8uzecXrBgNYnA9
KWoU/Tx7Xk8+zhDRz7xLI1kCCtQtq9b0ivOoPlMoyOEtEc2p69tE+UJxgr0B2Er91ysoBmQsRWwX
fyLdsK6cDVXTbWqvaM082g3693xSFKIJdn7+McIRBkFxdCwuWL0GXnYjx1fprAiJ9P33nf1nSl8L
yfDmjws5ZV6okR7Df+MR7lZK6cu4/yeXxJC5vfOVWDYWObkftBVOjPcLJLNr4G6OqzRt5jshAQ+B
QaHEt8mOoH5DTjz0x6NUlu5w1gvvV+65PASkgOeu7q4fHt+XVv64++3OcM2ttpf8+Kdmt4HQ4eoU
nG72Zc0J7KQXddqEJTMojLzsAxAXcu8Fdh7HtnfcdICk2EW9lcUOgEQliMjs44BCnbVZ8YkN7GE0
zkYAMSw+PWrjT6OzLE45B9gvQTIQlvzd5uuM/Kt3GFTQlYjN22QurnNJHGsGL4bIPFxw9K9VSxSv
a2cpDYzyjKQau4L4zzIHBfGdbnZjU/U4Gurvj17+DbB1SHQvjj3cuqhrBOiIBtDH4IbWkjFwO+ap
A9Fg5CAPptUEMz/TmQzdo+5fFtFYIMrTYG38Yc46yDo/6YnXPvSlUxHAN+P1f2yZuE0Eonm2oOZG
IEjt91M9D2o9hhYy4BS+3Bn0r3BLoGSLtrFdZl48PNJ8riBA9GGg9fDdG9tq9XNTQ8N6ubUFrqe4
jdzIcea0nW4dYQcVM7OD+gug7nqxpTi5PfZycTS9zvUaLhkaiCP0tHwtw3NKhDdxMJ+OAYlV/N7I
T3dmw1FTvB2fMInkDuc0bP/nqNbryGWMuDHUW8aM27a4aFc4iZUFpATzAAcmwaz+LsmgBaknMjQu
eQb07QGw0g8fMhV08jtmA9oV37DU/D+84acr1R/hLraoPePh48jfBZ6wiAtBsPZojviVI7oZw48C
ujBnnsb098ZzAftTBMfry6XIapMPzTF8DWMqcn37shbd9ullUNB74WAfVJ1PTgt35k4L3kMrmuoM
+Baf4D7cYOjbOk7m9VWjasy6ha9Ud+YLo67cJM50n411Q4C1mN7lIc3rZAvK2+lULKjeaqCIyCpB
mOWHT8Fs6SOMj4I65KKf4prHxgkJTWTTmgihCHGeS3QqCO/O8u+gN26r6ATtpBMdQ+NcjwyAzSfc
Drq8+ARjsn76J49YxOt0LYZMh0MW4ZJ/TwHwDj05oeHsrd7PLe0NbW6sdvl2boj8tDv3eEaD0BVA
8OKq1jXLVbVF6YCh5dhopHjXp/u7wKiZzdGld9dhG5CmXuxkPLihZxAs5AUi+C1viOWKOe5oyjma
UFK3BQsA0ucLcNyiANYw0gxUFzwMCG33lv0bK0hi2hB9vS0S1FNEp6OXT66GbUKj4cT1fOb6slHC
Uf2LIQEV9HXkyDvlCFQfWnp889rYtJal+ECHroeiezCp5idQ2NPOPZ9D8N9uxI734q3dBLM2+0yo
38snDcNb/oAaP1fNcwCVm5qEC1M4lcG8eN+vIvHhAvVMtNFpyXfh9vF4a5rJFdo/jzjSh4I3jU/A
yZbhMQ4km1w3GClc83bF7sMly9vdslcTzcR1ybrvLVTHhIf9z92HM3yupbVd90BM/mqnqK40GVxN
dDI1LuxpxMZVhmCUw/oo+YWonEAtABc6aV5TVsciRu8WlMWEfOO01V7hpYfBqXWijlzOM92/7yqM
n+pBHr75leTZ0UtSqUrlSw8kRwFIrOrBnQZuBlrHiX9vszHdTnNkM02SvLWAeISLjUzaZayF8caH
11IzkhHke0rHjY9NygZTlBJL1sUWbe4i4DNtC/vFzg9theoyHZOz6aOdGVflCSruKCYxFcfrTZZn
78lf2kyEmzLxAK4zeJjRDBy31XvC0hCxkpf5NRk6RhGwhkhxVNWD2JFd+7PmxOzDjJbv+Gwqfujn
3LxVuanjsRyVZjxDiU3VyGKB9fGf2wZXNw1REcrfNyEgJyFX4z69juD8eG2YMWpUaWEGlHJDN+6p
Y5Uy/s4P2kxgvSmqjq57EqqP89sWrTD+Oovmc/kvLWaxzBWt/94OdUMp3fcc4z/ec5Rw6JrFCGYX
0IY9ItwXpQo6Ee1/1wY5vcilPnQ15TXhj3RSHtYVBHykeaO4pnysbXKXJPQZr8/0sN88eSnXSpuI
UpVa6FG0PgWz62KR6LY+fzB+X4xnFWxUb+ZxtYfLkc84t0wDTc1/ssJvjA/yu2c4TltsDkD8odIJ
buTE2eXVNqwGqFPZorSxZiTVw6gzGpi8hCnXJ2KDhbzGEQgkFz+Xf72C+I0b3v+ETPXsYB/yNWlR
SCX9YkyRYzXKwuMTpbY59uHcwRHBeChpULLgyauSR4RpkhZxiK2Nf0pSjyssN3ESpgge/Gh41TAG
iQQOZer7/sFwLs0XLZpZsHy1ndIG9fnpCWLcQXpttG80t6l61OG3HbJ/d6iGMtHPP+AF2uPhqEKt
Zod62gadKdKiJiltySqduxjurXtYZTnWUKfvAenudo9D09+2otqKUNjb0jOpdkIiw341LscpOZLq
OylofE1W1XmceFfA0qZRIQbh80pTHvrPitB5YujSvcy9XJRPN6CyeLeqSMBM4y+q4l2mVKqdf/K/
x5UREvuX52MS/yQI2xk3vI+EWZ6MjLppTE0tjAa4LBsqgmM6MJtnTpUFvQ0hofZdXb96DdyEgKjH
OMgpr6H+FFyY5AkuRLScyFeDkC7kUcJLzlWeeYTBcXSBjXoLJE8jPpUxgmSCBO/gHTkdgS7D6TLB
7U3rib9yB4a2S9lbYbESswrpg9Y1pZgV8Z8zfYETYb4Zi80eZQCCzJ8UCEpOKsXB0Yi+PJzeKHnQ
SC4SgEC01zfryYhDnqwFBXyVb339H4db3OZ3ZsEhxqLt+qjS42uL3igBFlDMzTTNmQtLN15fHE+8
06WFsDtFWmdBxHRXRFe8fhxqB9LcLlJvo0FLiakL098EEph7TUW1umdbRh178IymhyOBl2bjz0JX
e1A+dSwDgN6DO7Dn7C0kJYF3m+gxF/+KJjbdngZY23+ITJe6YG7nK0ti6Q3dipzLSVhekGc/2rY1
f10SPJ5EW6pcvyDCi8jyA4+NDQPKjGCwcgbtoDa0K7KV8Td93hdB6TC2GAPvXY9A/O7c2hEYVbsW
20wMMyxLue20+fBccro1Aq0C7FhvQnxax6oLX+Hg8ygU2mQxO0grF1d03xttum5knHwdC5Z1SZX3
+XmbOIfLBYKLPMY62FxkWnas+lPqOENRmBmSSkNq3UuTpWgCeiXsB01wSoECWeejuaZ+13aBXtxk
Y4xRBdeliVRLdxG9oRRjuiK3NFdzl/wRmS9Azu+RBeHSaDE0BEC8EyQW+2ZM8PvFTK8arr4x0UiG
2Fo8BjykC6mcSVUMs+m8zBbIULTaDBcQzFtBdZaHLgpJrGAF++eqip3ASt4WbWQBwt+237dhECZS
MwGt9+jPKjpzGrhrey7QZbaQq8g6+LiHSur3YYKkteQH6ufdoF/KgQcDFnHkXCR2n9aZ+iAuvUNK
4hlaih/CC/44W4GNPXPlfxpxqLFSo6Rv0tf9CsGn/0HVEFOM/1NU7/rJpG/ah9o5Bc8T5yfKDJ6+
wwjmi71k5fXWmYx8IEhWp4dB44zi46Nqyxgnpn7lfBLG28reQ9Bgm9M4llFIQ0GaVTNrf5AgWfGM
umjMvhCv8+FQ1nSIXsoxBmHSPdcP+XUN4DkCMTjTW8nmngK6sd+hIgf35QBaMipV22HR9KA4Bl81
kMBSN6vqYUnaHD9Rh/PyVLp3dZnQLL5YL9Sh+km6/PpjTG3mYcU6vO0oN63ITap6bGkUkpj5oh2+
TFLGHkxEFfK4s730ZTN3ALaVMycCBU8toZ6Pm3oe/IrsYcTobFjEtt33fE6/RQSGrBsE24nSMyiD
ogoecJ3QnQJDnUkcQxfT6DUx00eERdN64jQLpStZYV46JVI3UP8R5OWUJDUbOkkAUiMd+NyaS6b4
xioDCXEmRmQmvwOHMEpDGwuf8BU3kVdGCLwvYEQv4P7oyhcOrV/rrMCOrt9sVXatXOC3LILD+V+l
QX7a16vBF2sqdIoJvuEXSrQWEFWE+NrxWTCq8QC3fwkg9kgCM593a8bXo6l/nhuVOCvsU1hLaQJh
wWsE4EdVWltdLAru81FojhBfSmjEMVoLr/oA4tq3j1HJwH8A69IfOXXq9iDRsb1IqyTJpGbxTWhy
Mn2wf6LeYF3SsxxyjE35RGiz+Avep3r/JxPutb5QU9UCdbYV64FR+VyRkkl+Xgnhgxr4QeDWdWaR
OuWpFRcdBSKTBYWr5Ov03DqtvKXxU3H2UleyECngnfgjG64h8kJVqFpZIvpNS3e1RLUnKivFXBTC
CpG0QG9XruPNd5unOvw6HjrZty0/AwGiT3gMmPcivtBqIznHnTxJGugl9gnnNiOS0gcSVDw127WR
TdvXQoyfVeqs2wwjg0bWE6gNogMuN33sID2L18seauKgwFif72JqA+1nywvXMUZ/6lgBNrH5e+jU
neZZ8Kvlc+O3zP3ZCrXlTwpysxaA9DgKwi7A0nH7dukYU3OoLmoH3hY1Smw4qimWNxQEd3bDXkZu
VBc2F1W+dx2LqJz82Sg7HtwgfJsbNk9SV2tTD0VkRfBJcFaytjhxORnErZg7YuXHbKMhrU1QGUMl
vfympInXB2fvkh8QcgRQqSWZnAdKKgyDwwPa98nrIg0GA/iMDg2/lVuaTNhVy+ajGmtXeqErAgqt
sxHSG0omK4Z6hpthyzocZJB7VLVWToyerwzdmsTkJ9hGrmt1/CifW+uUiBYWzCvYwFnpJlVxU7Hp
kFB3IWLWmQg2MZKUI4B3ABwjLnmaNZrUHmmw3erJsDPnPmg6prtcjIb43gx2chaA4Y/qTsADgh7p
JaZF6RIQKsb3VUjgs3UghOzsaxddyEfsup/wWHo7mr0Ynzc81mvI0HHnmt1dfBAGsAQcmUDg6Y3t
1FeOSY3XXz8wIk+yhEIAACCP+gEE5dNSjWoFfT7R4WwrlLeNXuIFxvFtFAElf2+ZnovQ95XPanoT
z8p/HjeoE7SahIW2QBjN150kM6ggXL/ENgwQM3Fe7GD2grdmNJCmYhSUNPcc3A8ExmknXxr7CQZP
9ELTG+bysVp49UWWTQcLNMf86htK1HDkOT7rJjWMI0WbSRb+qCDQg3RtWVJS9BLeeyJmILtMW/57
CbEXNzqQ4EWJIqqTK7UK7w8lcN0UVIxkM/tMHTw5LE9FT1kZKQhURsha2KCkwOS0MZuaeZ0xK1x8
4FuiCZNYEqAZvg/SJ45oEHkjB4x0X4WtYW1hOzb1Rz0f5/vxEG93WgcPznGiWAxw43QKYO/mRAkc
yGolfzre1VUSb3M2afPeZTcycE5g2MWUZULZIu+NNvV6uw8yZSEyjr5eBxOdu9hOFHiuT32QrM13
ZOAwY9puBe0pkEIPhtwZ11bN0oQG99GXTguqwvLDmD/B7njbp+38liDQhdGG15+iWyfck8S8M1Rw
6T3z7V4VBvNc5L7DttbXDM+iGXBGSq2mFh1ECBKYiSs/6d//v+7jEAEWtdIBcyLTA+HfCqN0vci2
EUtHchjvRCMvhuZnNXMFTVq4iu+H5g4bicSFKloqbM31vJ+fnv2wXRlk0bGW01r8piByl9brti0u
N1xZx1kccrvkRtUg2QV2ho3PccUFdQvS2saTKhE69EEcM3lzdVZXInFoTZAsW7PuHTZZ57pQ4seX
kODCQo+aLaj9ATBoa63ecgmqFHx8ocHHUi5F19yhbrIMLKY020Mn/4mo9bhTsi746vMeuLqbUa3B
pkNBrbnDl3Iwar5/m+MpE+GkJ0nV0ow6nLCzNe1P1jcJ5u7AffuLeLgdxbPGcBG6H8FY//g5OTpd
PWCr90RyezMGQtanrr3cfyRdmdZvaoe29sAKzdwfgzgAjHmeWlVM3nQ5/zx0KictTdUKzxTy824B
EW3dsrFyDniUr6Llz20fnzg3Q1YpJPsRLAW8lymJ0c2aR5EDiDH+IOfXIGH3PIudG2cG/rG8qH8P
UeYXBHS4EJaL5Sd44xDAAyC6YDJ3EReXCQMTM5W1MkQ0gifN4AAU0UtRWjlzASnGKJ8VPaHtkPy2
qAjLL6xdPCQxKQJOLWHbRK8a8JIBPEocEAWNg7XnQ4AfUwOLKezMXcleSma9D7XWjdkouenb4A0J
g8k88YtWbULKReWyIZJ85ja0EsYk617TZVGHP+rw+hZEpNmfKVaBeL3OB+CKphErH1wkICfUlWZH
tl7utKYMJBQqB/Vza2Iz9Ea2y6xi5WQb/ha4dQ2UbsmaKRmdbR7OaQLzzaDhNUUId9JMFfHyWq7y
EAQJpIw0soGkze+KllJ8cVmmrhWZ7xzuevVllHyoS00fIpLEHIfbNKtJuiMyJMQVObCNL4ZbNB5F
ZASy60FhN5RK9cFPYLWbVMk5Pm8595DduyQbrrA3ZzrUlCfARm/T1iFVfPFkZ/NGoA1f0aPNE2V/
kjr8Q1K+ThTabHbA1ga8sQSvfQZB60nNRK/0FRWdQkzZw6DMjI1s7Vpka9M8hxohDXFSjnbje+XD
FRx+ypQ57CDepbCyRmKc7BId69e8PVJKu3ZdLI11Q1RLDwhIS8n5v0y0n0g3Fvp8oXvuTAmmzUI6
GtWnOb4deI5H7eAQByQFSuHwVP+o7w7M44YoYORRJV5LBWvUUo75n+oMAw/G0XD8UnqDZMAUZvPY
OnGhmI7tsY/k3QCX+rtr0K8AG+qKmGwWgfCrBd6CP9K7+df1dWDbKIzFYi7FSUi3OHAB8ZJ4Tr0k
PSz23z2I/J9ppkgrYUoxQs3azUN+uwjMENAWvwOpqO5B27y2Kmgc++Ue7CaSjIOz5POReLD71FtR
eRYBoXGnbGGw9lso/9AxecgnIMqBgv0yof2wzYe9tf2G77bI5rFcJPrdJEUNK3NhHC9/rJ4Tv9l1
wBBQIPxvOGf+94HKiRNvym8KFAFkZgRDTH//KhVlmtL5zyc/GoRGVV/uR4IsGOznG44lQMRBpQBm
2ngJ2VdtaKk+NyjsKAIeIHYLaIR1+BMvSKcrSkGEDvA5CPN0BhqLXVu8pswQuZHqKXX1e8CFNt7W
pUCIF31eEhhFtBp2//nIzHgjiW2630qhEcUAwSWv+oAm/HQzYmB2/Fjq5H1Nt5kEpcY783WxGl9M
mPmeIQxCMdkKYRG1Z4LM8DaTUnJgoPAFWeBzpbeeKxppr6eUGHRxOzWxJvbNmoHFa40QSvt57zIO
LMWK1Cyxg6xe8QhKIeyHl7TLWfDunk6m+4lxt83NUDx0AVl+ui1Naz/BCLoG7cTd4LRNL5unfCYP
HXA2ZqF8o9NYmRbmP375Jpp6cD28Yy3PmRMSvzW20JAzzwFXq02pW821jeT9rgkklwlpvsfpBLTj
w5fqADDLkkeL7jHzpoA7l5o0fv2bfJeLWuI9fyXDxlXXuECVjg1yYkvqi4/n/3mPacFXAptSvGJh
mSdpzTTpvM8Fc0p6ebY1aipPLG95cF120ehQmgIyZ82X+VEldS05Csyh7+X3aa01y5zcFq0hyrBc
sFHKl9O7yPiNS10zPCjGhYVgJvs00btqclBtKeInKZk6SKpjoFQg/I9m/F8zEQin5TEkbbiosBVm
H4cjmY01AnM2QNI8zhEk+oInA8IEhwe51E/omWtG4n5298cDfm5+zsWV3YiPmcA1RyR0Vpxzg1Ya
OwoK5hpFPG5WjnWhtG5ozYEufMjKvD4rjHFl9Pal15wi1B1oYLrxlGSVXGLdHWXWbP4+Gi+2SscB
APnlOBg9Dq8cpvawLgJ4ZUvlImHMBqQdaA0Hwo3gjeoaA3ogr4VyaePP0avyN+bCO9qDbXmQlCAl
lmBpVGvqB599ymkZ/myp2gSNYopPOfekxgixHh7Qp3biZWVyQQSXgqxAkyQxA+QkklBlWJ1yPYDH
uNBB+ElHWsEH8Ws4vbKnPcjGxIKXay+d8Dd5CLBIZUQrrxgYZM62AKpwB12UAggnxEb7WD08jE5A
tW1GdcXBxY99H02jOzMzvLmrS1b6WUgthqLg57H8QYtx/20s2nJzy1qggdrVmV6JPQNrg3EKAtbE
4Tegl4m7X76Jwip0XBsyVNf3OTYxtNWThK10WlVyc2iYCMB4lDzCGsdotC9entTqJ4xCaTIJvxNX
WnsCuHg+F2HeE5/X+fRuxqmDKh1tdq4kHUkk1BAIU5+AeCvv1kl29NX+ZS7LGqRVHTYDAaJws1Kq
9iwQ436TND2JS1ED+M+AmX92w+bRPF2jFaC6JPZmNrC9IBlglNX2m4b8bfkd3TGF5iO9EWesfk1Z
3K/dtapYsVvme0E2p8wmQZ7lmIXO4B2TQb/Zv/Hq/ox8evbNogi2/qsH/2zFt31Q7bjfw9LLfa8I
1fJ/Z9OvKxGYetm6TRHAWhMqBVanz7zRn4JYCCiLERJv3g6FIcujmOD4K5kIi4rPaBTHLewJ2Waa
XMtn7cBNNUWnIXnsmoZ4e0IWbQ5eOzeyQuxUolD3fluFFGriacmovbBMF18nmNY+x2berUmXydOO
fsCAFvnunKRmxflC7UVr21zuMYr6EhAj0jR36HAyPlG7QkwVG2j4myzc0UZ4KxjuNqmaRFABjplx
MOiiPW4+L11tHya6U5/5dH69ugs3wkbw/GuDPeU29Md6Hc8Pnw7k7rathd8/fET6UG7tN98IG765
GxwLpD+kUS8siPieqj9AlLXNwVPb949E+nN/K9j5VtKzgzX2oS4/bjmXo5H735mO4hCTmCAxWpD0
8PWYGXThIZbfWKaC0tfS8cq7urgz87qCKTl5QMzRcT6QPCdtulMwdn0GMSPdyiE2JOm8LZoUmw38
iXrm2bl4ty6wdKE2tqnM0OsgvfwEkFRYytjfqRuSfhaoIVb7jCfkiIKh6lYtCSQ5fYvS88Ag4ifF
2NxeAOySnRPuMdpMb4ufPLgnekkcaMsAoTLNtABy0VGjiL9eU+roQXaAu/WgRJl5IPEBoVQgVoTo
kVfYJuCtTSlNGqhPhX1MCIiGouPDjSkXIbeRIDEpcIr7/hN9r5Was7o/akrZJ+XE+asILKUP6I+S
UbsW07FjPsbCqav8wqiWs4zVmjTFYsA0i08Fla50GdGKYQKVZf/qMebzLuyOZadERXeA0o8zMDuh
xMtQxXla5TfngDl4wSG9V254pEmsyM61Jbdo+FxcHLEXCqlopAVDAtM6uM2h2rKVqS5gicjnzdmI
VVJl0Vbz+xBGQilva2WYiVcTa0gF2KK3iXk7nRSFQnob+o26OXg+H0tCyDktHUkrtlzT6W8OtEUA
SNhOGFJkX49Lh+v/Ila6oLMTZpC0069KuaT4Vp8OIH91304d/eLVNnTQZO2tMd908W5Pjmz8fxuq
zy4wRHrHceOTxRq4dRhDZQeZzG1CJvwtDxe+kmPZwuotwFyCbpmC4XvWFM8rWYf9dovIMpkKihzN
usQXE+aJ178N4+Rrd1qKAJAmYwmJ6epelRyhTmA0BoCzihF0La1J18z085nKk+OSGISLhuRSUCwH
gs9goFrFeHrx79tJn+tQrUpoQb23HS7a8o2PP0Le2sgwwMR7P/cvCMZQkL2exAxDPcXVS53HtcuX
tI9ossSL1+PUUbHLnNjRX3bD2hT6qorBrQcBgmNTSwTTHxyxJWTfBnOs5RM1q1OLxzFYKszobAGP
jS02fexq6lkHT+1i+nY3FLR9O2swrfQR3nXUfABWAM7bES+VIwa8bSjam+4J/npqmdhE2EDTnCJ0
isGaKe+Da178xduTJ4KX/190ymrbShoTklPELbcnH1GDvmw9pXTyX6/U1r9zWkmINH0CPamnaZ8P
Jtp/sqT8rjnoCBamG0tVVWBOa3W4Tz6Z1xBHqCIVs5YRtYhPZLe0u94AUL9VtyBL6jkILzGkSiCc
ld+g7POjQx3YTa31aIp4qHE1z0VIIZ13BbiAFHkb3EXordYvEf1QWkN34hiWVFdNOm2ec4EuuueL
MGCnL7+oo3Bya91SvVYKMDnabcJGe7llKE/WStaNk7z9D5+MKIF+6DVeNZQe2GSUynbfKqLjOFRM
/u/cJfbpp0ezVKyPAXoDKbDGCt6aDPCmcPe7TJ55IwxG6UP+3T9okHYrQyjkZIL9q0W9x3fPiA/+
U/+urYjbQYGRahYJEctyN2oNeTUvH3Yjxbn6ZDl/R3fN5spcKS1MlwSiGpSldkcMWNIsxKbpNwl9
Z06T2KC9D6J7eUSUk6IuTLyHgGijH7fY6S2kbIdnAg5sul1ue1drdlXSRAwDu02QazgRPQLh51R9
zfxUZHHIeUIl8T+6PwixgS7FF9aOUPBUeVwRwHvDipNJOGQVxTDpdGfNu2sQOdBKkg1yRU/FpSc6
7FIfYHWIuNoMMAkmxQFcWMQc5tZ0n0gpK0sCm25DbUN6HQSphrRTszBnM0y7eb707TQxu16lQhQX
vEFS8qYReSrvXCZz2xbensFofVVHucik6dPls94KzR8zU0V5waqVkkKj8g8niZmaIOIGEH9K1EtD
MhrXRw6OxHX5qG6C90TkH+CrA16LBOawL9uWlVaR+7aRZSOSleojfM+01beGgCKjUAEjC8dFdcZS
91wHHKaRtOLQodKelp10GAU57knqLVDIYerOopBGHkhiZ2DVuSdHsVqoW62z6Z6R0Ev5dXxjxfwj
OUHcN1TZqcqY0VUSuscjr7+8q4O6AlbXfJdUVAMC/twfo9mJlmISSME7mAACVYRfo0QswuFidhXf
wsTNWyROLNvyiFfA0qswF9H8bsNiYKZodsMq/icxZYyh6Yoq/ePXw5l5h/zuAkBss5lGjNisiSmS
4ODin4Ab/CUAJSHbe5nb/Tlc+RAmXgDMZA3o21P2NTFpwjP3vFQdwpp2Rx57YHWOm/LaJZu+bFfr
tYagqmlDfTbbr8uembbuesm5QeeFIPkhp68grDYi1FnsOjjHDaaVJHLoxflM90qlSqu9zDhMut6w
e8ugw5OsDBpktH5HsB2cJsmcEhXRwPGkcGtuVgdeXxi8cfo9hufADBppXVsJBOIP+LvLvWGIz4ps
eUuTEDSq+vnmysdgq8y9ERIkeXqxB6JZ7fyKvGlyzfR1luk=
`protect end_protected
