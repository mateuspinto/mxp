`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17472)
`protect data_block
Q9RS7jcaEbFaqt+CL0LPJISDid+XyFF/DLEQ6hCC/MYEOkK9FNbQ0gBYBwrZIeVXzNg8JknnyzhY
jPzvJotZJDQi4XH/Xx9342H04I6JFfdeY9D+Xq9K27M6MRcauAPcYFUMPHa6F9hSuZz++Y22+IDA
5Krj9gQlvHe0zQV7LcX2eKsp6UTwJJRjuV1KB+zNXsFn/luu15ApyIY0X3xx89SbWA9F6YAkZ7jP
3HJyW1s5OHEcU+6xK8MbJrbTRAdTgYY2Zc+wyFTmKFad5xKAwI/QGETLyzIvCPfl+gZnSB2iKnvs
r+RcCX/PISUEnptcb5m4F+qgFhhfWtuADd+bXuj0IXM21vtCqmSrFz7Ql1O2ODUxlysVy1JKFJAa
r2uHjWrBPrs9MxWq81bMaDaJAdxvwl/zLII8C9q2nreddgQQRsJx7SCZjKxy/byz77yjAJnJNGKe
CgjjPE/DvRfIL1V47lzi44uvmI7+x53uvUBoAwOrrBsaaW+YO0vl2gLbhPOrFNPfJrrsIiG/XFGQ
vvPfoPEQyplX9CWt8O+nSWRV9Nj2WeUgQcADleOCbMVxW3nB1CUDCAzTGEZoZkgo6WUazDRhVRaE
2bfZgP0fFy+zsmh0SqvU19AejPYn/d9wy53PBf16pgY37msbCCJoF7OqkVaNv4RHgYPTgd1VwCA/
7ZM66LTsbHkTAD4D2BvN/cAqDKFO1TW1qGp3b17EUHdF+WKCZpKGa4izgOtFVPVQ9TdxjKzgjwdq
BPxhcAm+M0y2InaomkF9dySIVE0qYmwu944fIfkNEsX5Oriy3oWyKBlvz7DtFlhJgvjDEODHSjs0
eMTVtwlM2HTe7dKxAaYIHJyv9LEbCwrI0QU4QGP7j1N5Ktzm/GBSQPCWq+O0EgbjGm0Cq/aSrHD+
6ofyetnTSZEJ4jQ4PAJbqPhiC/2iQZ7pQaw6ZIXfclqlaLVlj8F1NqKfoJdSw/rlp26JIOJKYzvs
sbZJHOL/nLgUcEaQ5vip2q70xkSuSXma7P0Nc4yEp0kb4zAj3lLdliFLkVWpsvvD9esT1kZqmvrs
Y3NZsgQLkBszuYhuN+4T7Rpeq+D5VZh6yVjXQx7ZTvodaBHUrZLzyvDfsjBl9MIh3MYLOwF+ModD
vtQnojuUARgD1/o4KVDxuzI/7fDmLRKgxCmlQAHs5qjXEUZTvM3uOFDc+UpLLgLfgG/xsBQbo6pE
MkIPA5YLJS2p3oTbc7vlgJtKgf38PA1L7mdy5jjuxtzlPX+1sToinrtRJ4XZuRsFi9L4ndzJDzr+
j6iv8KlL+mcTcuGjHTcPdFOI80azwIPmvDPBfklXBN8ph02/ECtG6+8Zu/yQGXZNwJn8/eMph5uB
8EnI6MGZAZrFGnk/Tc6PUqRSADBmgr1KfVBcPvbeK+RbVwm0H9UZXSzS2WvsHG1yzZbDNnfa1fok
BYj7WJx/vOeqKUqSqBEyJnHvRAbgvLUXC95rr1o75KuJbdIIMexa5iApDJC0vqmtmWu6Eto91oEt
o9ndW/Yu5Ei28i0qP2QgPe0EpHehUljfECt/AmEnXVH8M008YQCV+zqFZUxGeFrscx2s+nhIUf5W
+gkUAcSf9djuSrqdJiWTp1YUj7gNs0J9GBiY7E+uiWb3WLcnH6aciACNdTh/rj6fC93FAFln7KxR
66WOWVf8SGggLPDN5VtI4BWsQ/us4SBQtnhDIaLSb+zun2tG36rgskvCZ2BX+BkxbupetTgQl3vQ
i27foF9BlrV+EbVZLXTl/YZhc8AXxaYzMrpDWjZUGvAkNZXC6a7VMLhcG4s+COv2EynpA3OlKGzz
5B2NrYGqwXM8MTe6MI8xYZohA4KFej9eJMziQzxe7nnDPJE4+7JyD4nN46Bjq9129HXELiLqBgO8
30BFkGyNSFdkPhH1EmnN3hwf1sXGwUyk+O7IYYfebX90AL/ZF+67uYcrmT6WRmHQZxxoBUWGvxE4
O3w1UtPRcbXcMkNsTaFGud4v9MApbf8fjP7lyYK0sUyzhuCxPG244U+ARpvtfElT8a1D4ast1RGT
WgFfD8aS7W+A9YHsSbZrEeF+Ps4xeiV6olFUIN3qML83U0EdJLoG3lqGCnaFCYhRAnpAakzlsWCI
AhV95nOgCbI0Usyn+QcPa9MacSMBRtB1gVi0NPCOABCw8sOhlXH/BNfbmPbe7gEBHzEBInVhhk6H
fIwtTiMtCnSz/4Fb2el7y9AdvegKireqdNvDm2FMxiBkewqhGSfNPwrLs/t7Ka7GFbWpbNjbR2Ih
7BD6iJT2UEst0eAQLF8kidHQYyKMPpSQiEdz+KQKyuVBinYMX2pULXjMdwQdoKbheA6W56s8JTbC
plawo8VEobBYE9TWNFpbBp2dUjCGsN6P3UFq8pl7ABOtDR+v0I2UMCNsImOW1NWHXOjg6pBcr9BP
F70DGK+YlRk5DLMlRBMJ+qhlDR3UGjRoiRTMlyVJApdexX1nUY/kXcF5QqXKq42iS2J6P7odOlLq
qQSBc3edlxMlL96BsSwg8Sr4dYQGM6WapOLlCx/lGapVbQdHOcwQlCZ9bTFEfDMOf2y/hhvfovh0
eRkEFz3Vt6S/yqwtAesvb4MqApaWOAtz+IYRMlsy20jfUj3ylrjrDjMfVe8PfYQAKqZgQo4BLJZL
I4xn4zbiw86cK/i8LMa56bmLEzgGsTNLJshnsY4TNFC4vlAuLOrL/F+THDDXpuozWhRtua15NpzL
25M5ZbawGHQqwh12xTCHqQ2KaFToTWoqH1J3n1LFnnFNQYb6Zfz2ls6odLyc7f3QguyyvqPv6H5m
dcEL+haWWnJfYK3AvNiRhWFprZF7U0ODvIEWkhSJG1yYu/G5hBLB70b/tbnPWMxodQ1hZMALniEG
e8e8pNEbDrf61GhKxFMhA7jMPUrJgzZQsu8Iq8rRLTWTwoCnR2bQF+5d6egbPHMD3u32JvIIxIOQ
zyXfN9dQLebOqFjjRwxm1bPOco9aE3bDQD061WQsb7HYUBr2IXibPLTNNZS8dzKAf4Q6Ko/BP/xm
1NaBjrSMmrZxo1/PH1RuccRnmPKVvYXu0bv7Cd8noffQvbiFx9vofix2KHuXB3UXNkEKgiNAiQc7
e+n9Rv9ByHMXvrBR19hsV/cFMGpSF6FGRrveoCLBj1Dw0cieHe/Q443nSmWgmiZMyIwlP57vayVb
zF6jZgxBjOPIC5CjQQBLdKPu5qbR0puYcVjLdU21/nJuhfiMTDZlFnK24LDnVY+wHjMb/Q/2CQfw
o5qDNX3Dv5veeYgl5FKdkF98vYxRYyTL2VLW0PC2rDvwzNI0i8p6PZn+5oeO00sEziHrH+QxSxn7
5T9oRzpEhaXoV2cB3+FhJFvVifP0l9w0cXbeNCrw1rv8S7sC8Tiuc4YLYrGiLzz6TLNB22lj8jie
HL3JGkIjic6pRlAwy+2VFkLOkacbYWI+gAsD8RqOGHfEMeg9DcEAtD7kLKF3dj3vPQWfqQZgtDcV
QuqhlF0v0TD++HHcn7btxo7O79NYGzELdeKfzF23HTGZTgY5d8cZzyCWhvc5KGWZjTABkp2Qf4ln
ZmKWk6+Vyz6OmGrbKwcdCv2MQ1ehDir8jcl5FuRRHv2RMQPr6SDA6azzRF0MVgP8epoOdpH/l9Jb
X/sXAaxHK5DqW6QX1kJaFFgGLmzJJzENu7tysukUJmESlo966dBS9pSg0WlD/WL3VR3dSX4/EtLX
rc8JbNp1O1ted23JugSumb8MXFL+qAGnwJuRwg2dgxRaDXtdfAuptGuh/Octi7nQnPmyGvZazPHd
8HCepdpndnMlu4TzDggxDhYj3+noXDLro8HBsk77jed7y2jyFa/ikYlE3B+B9KKpfLkVl5+Cd6xf
ihAqY52/4SCHoT4d3wB49iP4oDdvbnliYxzHMhLBwTRmu38jxEuPzjFvBbx0lWEWfxPJwn/5AjVX
c333h0wLsOrdKwdS9r4thU/CvW+zqwG+rj5hEQBYvPshNqv6cpvgYL/7vkNLSCv1oPonPuhr/3Wm
QwLFm7UIif/nnwu2oXlIAMRoFWEM8bF+vujtTOVA8m+/SdJqeA+tLCVs5Q48cnhfCSx5C7RH0RQ6
tmZWtfEkZ7fF/4l9sKz4U6CJOs7jhOPKI8vf3zmswJReJqPTqKBEcmIAbay9UeblpV1n91t6jJsA
P0uyKdz3BHd+zclfoOni/pwdihJmbKKsANck2Q78qEEL4D9HbYOx+MD+hOkg+TrM5N3AE8u40HMK
sNxPvsIts5iTUVgtabm5RY8/FKlvhVAgQ0yYLrTRQvlMffGZSscRxqOvlf/yYYB7GOidLS4V27s+
pDFAx+pYalRu3c4271bW1tP6Dw/oV3ArsfhvAxxal2jMVTZl7eulclwtFBaAn3wBeeSi1uoN5LNq
YYZWqYcM47+J0lNUVc0Jc5e0kC8p3dsDIIO5btGoOfQp8Ny7FJIsLlT+nXSLfnY0CHVgbANExn8F
PupAudSPnb3iSYsDX06aSPOAQcb1IbyuHI8AvXZgzvE5/4t03Sv3LvjRuQuuHdwB/hxCx0gqoJZO
eMLMEGlIYuFCMgtv50sbKerZpJqY+28sZvgWbBt5j0OnhB0BJ44R5KALLWNmW4LRWPEquJE/aUQW
94sn6Y8ip1bJ3xYtkKGIul2bMQhb2LYeInxuhZ8sdcfKdS/HkxK9aVRzHXybynX0fMm+MF/i7V3S
0yHZ3PwFgZuhFwiPJLOYqgJUHX1KKQwlkFJP2ptNnKijwOy1RDJwm7R/h7wHat4S291jqcxp7ikc
VDLbeOK5c+1w34P/sK2DU4sINsC1kD3rRxU5iKZf0+268gGJCWbio8rv8KCRHsVumEoF3Fml8v6R
8YgA/79gmelFYYToYjE46DPvXINmdLsOdFvv+jrzecaHoZw9GNK1QETN2ABiPXn5jMNl+/FkokUl
C2QzFh0nsonWRsiU9PZp3Ps2Wjo6zKBYECxLvIW7jYCCVunJ6y9gv/EVTM7lOWMKGByrpNZxunqE
hIoTXSO0BssTIMEk8XGut9Mlw0DQ9Dp6mhJ2+WfYL3vbHCF11AQOoUHdsXrM7L4qj5SPyTZnVZ6O
KHCQuFUIuWyJ2/Es8zSzpFxYpnLcRcGknTyVYkF8LRy08pb3Gc4WAERRRi/6rMyXQ+cpSvVSB6BP
4qEH1VUrFvr7hOPdV+cJTy155TtkHsWDmS+ooO90rkA7sc2RGal82ZwUAalXk90rZTFmIEfjy2wc
zlYVI0M0HHzjqHOSbm8Hk4p50cHl32kghtgf6+abHlDylGwGYoBBDa+c1IBF6cWKu6Vu4Fzra4pW
9AZ9GNx8JuQo6G13tTur5TqzzNWG063PZI7vSOwBSsArb5ACHlm6AMy9osstR/NP6VWFq0vDU8wP
GgPo7+9O7+yI26GHZ2YdshlmKPyIouUnngPSh4OTw2tcMC7GOryXhRdlr34vlzxli1Yk0sI79mp4
aij5ko4/2UKdFEBERYMmDhDIqRFnVo60EqpElh9FxvkqP0E37xonam/cEXV4BNR7oOMU9n7KcTPH
LOye10AfiXDdbyX0ldlOb/gPRyHr15aAihcVDXbOtfMLGKnGk+Qi8Ua5P11BgNNZEGdlge963vay
qjsBHN9QDJ19A+vch9sWdpMkrtnhMkg2ZL+0CFCMJ5U8/xEeno4QlsYmzFWWfJIIAH+4lwXQnQfa
DgE5b93ubhUXV41AkZ4kGnSbio5bE5nbDPIypXNYPcajfq6T0YkC1eK+6HhjHLSUQezBz2+AiQO3
BttVuwXXZJXoHSVRKJSPt9/Y7AG9viLNrJfLFBK3JGM9J1XtLN9ymO991aJB8eyGpMTWg4yM9aTJ
d46DCYJfaduXYsZXD44827Cx+PAIjILbfcXA/1ofiy0R9HI9Eejhg1b+GeoYOTbrcAkhh+yY5klt
x8AyR/nieG6igt6zBrUwQTsRc4MHATeGt+VE0a+zSaAe6JCYL03nytuph6URmGmTdZ5aV2hvsicG
EHlCXdmKzGpDWsIZjRHv6wVtyKa6w00H74jnK3UqYSbHvMWQ9IUehWu7lmUCl5X8FV2Lyhpqx9+I
FIlonhtchngHPIdle8ekgbFdrbAtBAINDdmNkeQH0JY7CAxVJlB0Lkemor74bvT+3N07/VKdjj5S
BwBMK1vO1YlEf6YZvaAWIA46wY7x9wYZxmPMApkgcsfRaa1sm/L4QK2JuZVP/kjR2YyNTquVFTF/
GD9pHK8l0UkRa97vP+egGC/Dpuy01wX86YwDwrEfA2LSqTxLoK5hpg0GCrXuEpPqNlLdKQ/wnvHY
QBporgVfoGSFPRPoLUc2wrC1sJmUPStzN0QK3vhZ1NI2aPyg/9GAJ8NnNw+zW9M7SPUjf96lsGU0
aJD/nIt4ZvYQrzB+Hd1CzVXMGAIrJQCTRWzXlKiLFxTZ8c0K22r6PIeZVJPV2oKsrTR4V1zsCsOe
dMz7eWiM1c436fO5jnJoXu9HMeUySWoTmtF3dPq+Xxcg4AHfYKvW6nlkJ9LspRvizosRPM++gkHe
otpFoZGPaAoFCaIvThxr+amaPWPFQq9jpIIU1iDse/pnfEjBdWTo/oxypSz7p0Iw3mhnDZf2WLrQ
I1DmEzdgM0v9ex302LDzoajyqUBXGtjt0tsSwvxD1rM9iaf9MEP0r9Zm4UJzQx1vS+C97yxXl3pX
k8UEz1k6EY9CTsHXz3Dhp3DnJcAtJk+ujyKqn+zj+rmPtoDaz1TzBrjCcrbnrHqDa/gtxowFhBif
9s4uJvAooyMdsx4CdyZxZWEkT9hVWgIbUbSIgkT/0hQ8ZDgTBldy6jTw2MC+44D8oxWop2Nh8rLc
sDf3XVg84c2xSBjfkYpgXJZ0J6e6yMgOzUuTsQ2vSuMSvawaPUg8++7RJACV6GWZ0MjXzSVu+5AP
tYN/w40850m6/5kJqKJkMcOvh+xthCvgqQp9GPBseyhj1X0UyF40A9PrCroAkb4pxuZcT7RAP4GT
5VtDEw8Ec/MeyWvlbK8Wsl23jtZEFOFOrfJY90ij0gUiUVHNK2JZGFoZWSc0EwTzEz9Y7tbm5Wic
6hNnfu5TCRS9GLXMANGIHcktCPZrbK6njB+Ah4h+SV30YelipbQPg8OZEaloeU3gC9JDx41T/2Hp
o1nRHbZ3vCSOb9w4ZQv1n1h3X5iLsxnbd3Q4DvqcSpdNm6lbv38C44Y271OqAUKmfKGuVJLuEuF1
CFdinyLL/p0+u79lyHGKJ7UTw4+SthF8PRSMjUe1UzrKuPkTsRbvgu/s0QWPki/igMK69l0NdvNj
+ycmrFV2rMbH2i1c10UxUkWBThOGn6W4EYIYnaxpmuB6xDK7Ul2hKyOVcleRVnc3pZOo3jx5CknF
5UxKOD4Ec8k68tZJy9oMJy1jGrfGMkeHeU3OmSnC/5iRhWWC8CI8NqHpz2KXOyj4dWxYrOjHJrhx
pwlmiEu8mLB1C0k/tvH+cZUkN2TVox1ihFP8n/bBgrAmaSjseLdALnBl2P9zLaKonldMzlsisZvd
LhxthDuUTzixKSEOIIJ9Od8ZQ9oWC53mt5fOOteJeSh3Rk504xY2yL20yP0rsL+IeIiIv1YsXPqo
a2J7iwYuVO6v8Np5sj9IgEjbLFAkOJL7J+9nsm8oVx6XHVOjxxu6R/nj8Fa41TLU/Q+1GihyfeMz
QBgGzNa5QUq6Z7DPcwFXAnYHKACdqyQrfyveKfGosBRPatGwOdybjknA/DFHV6ORYDWl/b609anv
kvYuUznlXeUYf8ayZyGEG1g5KUKGuRBmKrsy/4TzLnzUzachKKfgCiloDydCiVdk0O/H4gFUVYwP
xNdhsA/k1bp1XXEXbemJUMT3XlMLoVHZXx4Plambp/xEZ58eJv3gld4olwX+sNkdEPZVeatsIJ6O
4tCbumjGiVkJ95VsqkWJH9oqNTPDgLKR0oRzPz1uHrJucOYNb0y5PzC5kfpgUyOCSCPVHN/+vpdS
jA6P5cxwytI2teJRhYsDtBdh5QAhWBChlsq2ltiBzyxW49DPjDY1Sj7FdW5aqmcbAskFqD4YLi1p
EMGrGpE/CpYCJaUBcg1Pg94EnMfKm6RTLNqILloykHGqJOSJjc/qS/ptuqHeQ6u/Z7iz70pd0Ikn
IIBRNK3cFqPzWkTIhqr5WwvDymDvCdQD1AGGoxTDWOWvb77u4zyv3K6Uq5Ti+qPkjc7Jh8gdrHYI
8D+TZeAFET1jQMMQ8R62dGgz7jUW3UEVZKaIQ5jn7hHC8Xdr6QWOvWQee01gmM49qnhX40XCMfkb
guTUZtccnxElneJYZuQd7Z6fpicMnGyQGGWn4hRM9YQHmDEdImWCnIuIpV0QWzqw0yd7N1hd+BAP
mNfaVRqqD1YZs3FJ8VulFd36qAdA5cZ6GwoDdc3Jsg66oK8Iij4iE9wGw4Uj9+p6uqL/UtfoORNk
+uokaAaP4tYFpYVunb07zkoHD7WkOsIrtNKvWtCrx2w8TZRw7q5NBbMr8g3uRDhvElMWYcvDKZhx
IdqxK58K+8VdYE6x1tLKiSxEP5JwCd+ArN8olIj0/PMVwk0X27MRXhI/icqdibS/UOsSmyF5D7sj
2jwreVuSL2Oj9vrGaDOIe4weZtkKeeEc72RDqAG/AG3AsDpyNlDZrqRuTrwhiLMEbvuTZJ8wFXfn
9yEbVVrv8tH5KZOxwN8uyxJSwyc/+YgCqAnWUfn4CiLyeH3h3RJzdFnfCkTnPAmImbfHUvuyeRvA
r0GXFLprmTOUPfd+h/GFCc322UDVywmSki+A1g5Sx0sZmbNGr4LjphEhiFqPxsc9jxU+giK+xCjM
fdO6ryRJAGunmW4QNH7rqFiyCGWJpUd+mnbJ4zAwKfJV4eTOpdARhXcDE5eyfIplsJVcHl8qoUZB
KFIY5a4xkxn3NjqMHBE+Z9uiSzQ3Bc3paaKFkifS+Ls230fnZxFxIswVfS4vd8oh37WoERZAwRfA
Vk9ARaax8QkHtTCQmsmYQSIj/Pzn4KYeW99aGbdY0ExmUkZb97avjvYw3Px42DgtBYcxMCWnqQm5
epVmUgDocowftxPncUMR3j3GElihAzX+1vLxpw8qWmID29GmtFoTcJew/5kc3Jv9SHldtruByDqe
pFKVCLvQIPjofItM64KJFiIJgy9xJVfsj9ZkAkpJ/h47f4Cbq+J76fjHIk6u2uVjkHfpglULD50w
N9XtIA/6Om9JsaaZpqivPvM1zuoUSplBkmj8wDNTlkliT2MYHAF5vRxgT9RkGdxRfZCeRopN1R4M
O4OVge8R447tWWIE2kFgE/+FG5YMeX6NwbXSYW+vlMvQKz1tzFIGwS3980vlmd9KB5rPgKhR0pyQ
Kyhe0bVxrjPD2GtaTFc3fFWVrqSjarXCLGYfaX/qqMWxnOeKyTnv0Xk7QTlQECOBuWDRcQdGpTKB
Wz5UNJDJsey2uYOTV4rROB4IzE2ObECIbxJl0WKoll33Yp1XX2eLpNsugRPZj4dc5mYqI+96uaLR
UCzDtn1HDLWtJogNkGRfoXlCCHYMaKu/Y3+VXqrM7t41p7zucylIhyonMrJ8xs9g/R3lJ5/qRfbF
LvDjTOdcvmK/QaNqyCJ5x8c5i1yQTXrvc0gfeC796CIDXPbYcM5hvW4fHjXbbLAkii2PlfPcH7M1
nJfJp6PXyoPuSPge8JP1GeKiVoXh9807ZqYLS1O3G66LY5J6TJD+3D1FowSNvmRdqDLFOAPUbc1d
grqTCn832fzE8ALyQEglwwvQUjOsdQ0t6C+TiXJ/pOtso5RVjbgPa00PGaxXdgdJvPcMW3NTO2pN
p/kRTt539dYhTlR7OK78DFtuMuEazSAe1pJEUk6a1lMYdqi1+S9D1WUR44pzahP6u4aXfzODggYE
Q2PkMPNdwmW0sh2hBYeiIWXzcdf+0tqw5dNbSdIfyfRzVQVO7FcFi625Q7yEZvK8mzBM8zsetKSt
n6cdvkpgBJEwj7Lesbe63KqRbPiHATO8VrSiJln9Vma/1qR+zA4CAsT6k4zD2K2Ee95+RQF/e5lD
qcsCbK7qYZcDdPWbmbPQ7FYzEm7UdrGnSJFHtmPBWtvVxgcOt3DLFp2I1Ih0SkIdlDqaL3iNSTul
s98HHq2GdsyiTuXRI/+1mRXLUkq5Xba4KF05aO9hqVa6t1fJ2mf+dsbNYGOegq1XjkYeYX5R85Ce
yKz81NSnxnXu6aqCkNjGNg8bQ1/ge5TLQK4egjrt0I4KijQH81orBeYnEfeBDuOe9VCCAmCnM2n4
OvTk6ulJW9MgXwu3f7qzfP7OdgrwEPTv24xEDqmisonLz+d+OBQGUQUijcTBI1EK7Amw5XmYqaBI
PJTPrsVm2TFg4YaJHmlykLZYs8kd72+YD7ijm3f8gj01VbHWto9k0IxCRzRopI4H5/F3plL2dsFA
JN3jNXHvZM73C/iOghJIkcIHGeb+wzYRn/nN91vQc+fcB7UBu1FWaj89b2aeLFuoexYmr4EGCK3K
1+OjofHeE3YDM9HGx98ZakAX1/TdBjTZc65HBHC+JzxH8bBtIf29N/HLt3+5FTpJl4PKhJJVWMT5
XabX+wSS53JQUKDiU8ZXo9FD4G8bPAbz+xyScYDnDcwpVnwP2KOpy2LlbyjrEB+aoN7GCseUc7Q0
bSwE/En8EROji3g7x7K6Y0scmRuuc9K/3biXKWSkqZUbWCKfHuiD3lORypRBkv+yTGv0PkXwfYqw
3d5McHz6zWCrc/EC2n1Y3HJjCJ4wgH4bHguG6RZGoBwz7aUsXGImwMx8ohSDTWa2Ajp2EoHSehgt
ymx1eyIQ5f/LO8Yxxn6qazQ3EeV/ymsIoecVdnZtAh8ej3f5l56SETjV6x5ykBpd+8hnSiUVxJr8
7qk26LILn/4CbOPa6adRgUTpdMntxD5vbwAuIfMgeVSASSGginlMvTrXSCMprMpCEDsg0+3cYzqv
3ic1YS99BsXZsE4JYHc/RD5Mvulw+lx3vthuTNe1uyQVMIgLeBaSOPX4wM6uOsqPNXm4xI+BC1Tl
I3lhH56O2UJSe/vsHr2WMuEphhuuOMS4mioC+q5rA0gPV7OXJ84PiwvVnpqfstyVW4rjv2jOuMsO
H8yhMNRdHJTo0PtihyiUGHB2EYuq9B/tWllkdXvKoqkjVsPot+MhSc4Rqe1xBM3wFNY5IHz0usVW
p0Kc8vdRsmiu7vtyZkFfgnx0VDaH59HENw0lR2nkFJ4r6NoPFad3lrhrqh+5CFq1eVqwU2n6VMf5
c/+gSz8+3byS6DHyamLaU6O2i9NmHr9a/buCd2vBYjY7UZM+sSCLJ8N426mnmSttYao6QW5smF2h
zx5taWSwzz7E41B7jkn2TdlhSLRWeG5qbwCOIrrxrAIptfzWAqk1ZrvXmTId5SmVjrJqrUJszH4W
ZaU1vqk8D37LxL2I/cCicLk+vqTe4f7raunu9ecAWt7+ytIRXxESkx4pkSlVN6TvIC3F6ENMqqZ9
MqrawqXs2xGX8XtUjm8TKt+Snzx4abINFz05+EpiIAM0ZwxV3h66b3Lsvmkw/JRq/Jx1JnCXCzK3
N8OZzLKDAHnbbtixhdVNpiTNL72P41zWLPZOvcJn8rtRFnO6sdACygWT5U3Vv8e23XNN34qwknZJ
DTuSVhGuSpfkEZXDHLwngPJq+/P7RwaxgLfpliIsotxdxxHHckhdgku2aqYWlfzw3k3wqUAp1qnE
UtYJhAXnDnqv1v5lc39whTZAywy5xUoajiUpCfsDJhVhYFSuYEdhRnQ0t8jfllLEGxm/Z1cwPYd3
TqcSliSICH2pZ8GdCXgpXvJlNtllatGxoFN0gjriCrFrAAKFgUcZpn+OpDdEJa37t9UyWBqAJwVU
Wh4xXk1HpiPwPpQmWtsLbM6BpiK5Bw8+pERBj/lv+UmlMWrMomP3H87VlAzCwCngsD8n+P0Fznkk
ULXl41tyv7MA21Bw/Q7lDxgWDHEjeel9TEhg62z9o9hTYaKHEyhmj9y4ziT1zLvEdpFxghY/coIF
rsIwTOVfTK6GmD52BCsPAXwcd00+uYARl3KmoEtU9Atnse+YZYyvNcRt9b8k78DnbGu5eOfgHsFm
IBgPHeiKleweELDFX2AtuQ6/aQO9aOyqsA8R4h4EgFTecP+JRq4uYbq8X9LI2fwm9sLjnARJax/4
Bc7zHuntGNrFknFg1leFuVzO96HtdJciA/gSjiPenxCLZyCt3U5pdBaETJBFRjzJjPu8OtvTBnF4
ElMDXYQnf77ApYl8mfqP5gZdHpgP0cRC5VWpgBDz1v66fvIyr6K9LCvKRHxWNyHu/q4YETQXhAih
vl38dGm/aNqFmFb4qSMBr3SV2+qr5k2xI2+WCwxRg09n5hc+3ebKYUDVYI1W2QU9V8BqL1rpKapS
ik2CtgBfaQIQkOEKkYebUAdimYVGcZ/6+1G4IJfto0JP8Ty3qLh2kyaHXuOcUUxv4GCUwr4bj2O2
rlOehs2//Zm10kHcv8mRPp6m2fTLatAbdTDpRHTL6ldw+qdOjzIUhDtFgx8vD2RYrqKTfJbB4YYk
qgTcrImMcAd3z3gONdvcsxePXc4wEizlbfADhPH6zU4BFhQII0NEwRygZofMyYp02/IvqNDQS6eK
bZoa06pkIP+DGL3OK17mz3fH4SCd62fkLypz1Uycyng2WaL3HXTXYbW+W+K0o1LBwglFQoujtPKL
JSmMvIwcKr7S/jb5TPeA+aNsyvrjdsgjZGXwWz2sCh2acv7c1r8O6w1LUmqvgphIvzUtCcniL/Ai
7uA3ikZybBqSvXlXvrVBhK8yBm+iwfFEVsNHS+nnLfG1W14PoIQCYFNVL8cnADB8DcA2VRqVgvGN
aWSMGhuLvsX7BmU4O+wZ7Zx3zqWl7GXsTzR7nirUW9GQzp09tQNmAsE7siEhPTi41r44gTwgAgbU
jhgfUEMPsV/ahg2BIqqS5HYpHNxDr5GT35zYPs5hfyVMc77+Vvmw5nY/0RePHejce2ne6ReFq+hT
uvSBnoAeIrBEFKQ0bwkqmjkJqorv/jaokJaS5GdBtrz0U0UJjDJ5OLkEY12kfsHNbXqx1ckfM2q2
1vAo53ioTlHijoxKt5Pg+57H0hnU2CxFLe5iTeQCQhQBvxivixZ9e4HuGQ4fUXsNDBdbuh6PM9Nn
phNY5mCCv+kdRGV6/OkHCOXkpmkYI39jB/qN0oYrZRLYeRw6A2MK4MBPP8zz/5sKNimCD2+CT8Ts
zG5QfAoAjQG+A5qbWYG3wxygtVzja22UkRJ2DCgT4McqYvrRKeNaX+/LF6zYA7T5qnqDiOP4a7OL
CjhTPADmJF4krWdTq1+tkm6mKn5xzYd6GUJ5xlYLeq/adLPF93+M8CaJblRmVwDppHitS4OmzCNm
f6WaEyIF4iErVyxtp1aY7vA8IuY5IZb4JJkVUX9fRM+LAprruuG11Z2rjqoOEIv85nNFbc9IVf+I
dHFWyQ+dki0/PF+egpG9KIi9Z/oIrQ54eA5z7RNmNssJply5OdHR5VI/uh/YPP4kxhOd/Weh/sZC
a76QmUgLSkxyD7yLABDBZHvtM9mviH4Bn5Keuv34b3yisXskqBmWi3jcPhKffGHGoCR0W4upKysY
99qB1lMM6FIpAPek0QQ4LFB1OEeSLynekOoI/1jA7QS8PNuCJt/zYCwl7i9ppyLhfz5XGZ9gYPUI
RT+tnFfpbHF337k0tvc/FXQ5l6ekDwfB2LMGLhKfRuQd+8XYNjZV9PHVQ5gz7M3EdfekoY+HOKqI
lW4gAcfradhbqkXTAMQnzQnaN63/3UiZlhz1if7M34CVDHgXUY3rRH7Ecu/ccHdzWraIsp3xaE9k
r6fdU3oO7UVoE+xkGYhhGL52u1rFU328Sn9+NBkQ0WsKL4LUlz12+kNwBp5vjqiDdrYFMnkG7EJ0
LPNxAlJlj96yKFpPCL/bcI2Hxtj1brTKcmnE0ruDC9LbNpN74sbvIE+aT8cKn2BXk06IdH6IMZFH
PtuGQo6CqWux7NpbS9FTsvlRMYG6flNDB7Vdg/pmoblDeee/MyCnk0K2sQuV9XCJIFyIOGmU6YoF
2fjgaVheXj1kWg7NHDbCnvhJ5SnDxbDVzEpqo471SvwcJum73BDfcxojlt4bYlRJhGJZQWasZzsw
CbN/wqh0rRXdFOFznXShg2Luugnsy68jAbCHT9bfldEzJTLzIH+ApUXchQjCwRjJ2PLOqanMrQon
vgRDR0sNAe5d7vEfEmxmfSabdNg58OOPfwewUA1eNh6BSIr0ezvfHy/GRMtiee6zgKqLww8Ojo7W
8fsvM38cqmjHGF381ojJ3xY0Fsh6UUeI4MKmZKrU+ZbwUKI5MaNVxZhhvnnS1Fc9ialu+wtd24Hk
CmvwvYOhc9iytqLhT6k08yq2CrljCi0qM11I39BfiqJA87KdhWkkHwqFAbYdtOjD8yKMjAfCQ8c4
nqVO8+YcfinvwKWsaSSa/OPfclfOm5VpJokBVNrwNL4aPzOm+ON7r5iF3qLULp6+JF+t+GkVYMkX
QFHQ3JYR2aN/pNaykz6aHuG5bZ89Z2pYDlDEcht4wty2rtiJhGeM+vTRMyVoEL4+CJF+RUe4Gv+K
xJj+8TvYZVCXR2bY7wbAuVYwQnR1EsmGCC1d3FRSlt8eEEcHShxlFz0cUgbQLVl2+TzATUUx08KV
hUGSf8x5gjrfmoat/cRxz0YT/iToCMs9lY7LRbVE0J0PvI0NTvW4sn5OwZ5Rpe2MsHaRLDwwYD/0
Ga1j9d0FA8F2dt2+4DTbkyFLsbjXjwdTNdLNM+B90oTHE1YbL1JBL5XeRytR8L1XmiKRjslwtG/e
GO/RyVSRh+z16WFYpKDizt+J/d3cH4EM8iotgZw6EAwuik8wziyw8ty66kZ9vTdAEVyjoDTwPXfi
L8bvsdvPkd3rmTGI2EPhjqAmwYKGvfYl3qXgE24nGNThK7EWDaYqxiep6iEIdHXMzMQUQAOtvS9h
2jd8VKJmqLvXoIf/JRkiO8PGrqEhNR/Dh2MNMlNev+1p/irRQm7fgpfFlNlVHKylJPtMj3WP7dzJ
OhBg/JMnwlZPntbBJfN479n5AwAfrfdm/WHNDcB7ttv1qzidPg9k28vPGQsBttyAWfUrH6NdkNf2
KFKNYSclJIKCnBClW8GTlcrL+TVDxAHW6NYuBm7ogkPpBqPDIrkaaKbGpciQKXxzX9ejwjXqZFty
VKXHsFmwM4ZfYP/1Wcl1+Hwan4OLuvsspjF7mVkepG7nt+qbwjad4Sw2tgnGPWTatfXSwQs8FSTn
iF3EvHWOt0hBSrgyDN8Y8auIgIFzXQgOQ3n1pSEpCLO/Cfa2pSkaVmBYm3ks7GTBnwIYIr7BcYyV
JOEQqDSoxAth+3TH6ToINZ8xOSXa5goYOrpfV0hObs20rqlD69FX72YQLvQL1ytuUMrI/UX2n16h
pWi1byqPpkjPgTDlD51AsnaACigutx2YVi3N4KG+zvjBVy1NDgFk9PT49vrtP5h2k2v2aEFdTK38
CRL6lpwVlMOxQFY29joA0EFlghWrx1WasO7/OSY2tSB8ji5engXh5fmU0hmsOHo1u+tfNw5VUsbu
nJ2i+KRkuqqvGnyM0jGZJ0gVzOLS+SCqWYC1dg5OEwJq8ZGW+/RSjWlp2LJmzAJM2Yj/66RwE7/q
n3xfAIMeb05mp8FfEDtbaIPsa4nd2sG6VPgG/kkjM4d37l1sg6xhk/hUY5ClGSp4nhGV0LxZJzDC
v8yUWiET7gq6H3y5iNTpqnExblEqm/cB3LB03eGaIx0kJBFS20GQNp8cxosfRqArE7hgrwPUp70s
PZpAEcEf+ghUXrmfi5aubf2N4LgHz9i/gVaEdJMZksQvK8mpi0xTCSQUX6Ey5oHMU0r9MGzij8LQ
KgDSeB8pEN9ZqkVn913TJxP0YtQyKNcbtql4FvJw+134ypgeapJIVa/8emhRAwFcUEahdRzPIgBG
aEt7TnfC48IsAes0MKRg7kLqlv9m57t18KZEV8jJER82/8DjSAshUxQW4v18ihmHvjJaWe/tFDkE
7vRsCE9IV7TohUGL58Q5YCtaaOLeZ3Q7wslvCBTULZlP8uQopn0OYIfuQ8TevtHKgmnmMi+VYWzv
q4oLm0T82m4xFMd/66n53xRBZinPbYJ7TVxfw5+eOk31Mtf04lTYhA/hfLunba4nPdS4EOwcRi1r
Kq0JYrzorZkTn478EcHadc5v/dacMog+BejIGLSxTc7An9i21oYx2zxX9v26w9duZm87YxFDrJVb
FKzLz2JhOBrmgIIFws+K9qIoHSVSbXn+Uz1OawI0TKFfk+dTLS2TpjcR04wNlh9uy6SewoydU4Fr
9PTPIKaHO1U7URicfZXohr4r+tmAkcMra7x0Cv4rQSVUuDzQyVOqtYJrUL8eVDwv6zU126xJMabD
gR9Xtrk6bp9CN9yJ/auL7QYjxShdmLGMqnuFJL6BICsTml1gjDW9ex2HfVU9Gm/iHIRmUEbblScv
Y/3a7ZgvnZw/sZ24GxWBiHP6+TBnmwhD02zHcBuBsaq07LJZC3pdktpkm1eZMzxkSm5gJjILQYBQ
L9f/jzCvoe2gJJgzGudU2en855fRkU2zcr1ax8AkDKDu0uooHIXEumcogmstKvA6jOUxmTdevjVz
+rwB7ETqkmwTyfDTsrPW2yxDWZmWpv4Phwq72FWC8aLdxJQV3PBxVPOhsDcGd9DJX2ulb4aKV38Y
65p+TGTupxr54zkrwUnLrnYWvGjucVRRD2nsajccobSaCdEzHJS994xzeacEEhEBWu/sAYHNDjyJ
CKLmLPgN5ociqlBhe1NUeepXSi27t4jew2gIGbqojTTJwBSxzfzyHYNk2nFy4zUCi9J0Q5ypSZtG
QEFaEHl3chkdrG4vOBc6uU/DbflkcvAiascpNvrgyIfBiF4G3NaZKs1LRyb5ZD0rLMtuxi5xni/b
0FPBHLZO727l7quIWbQwiSk00Yj8we+2I0JSOeJvChykeO2wjK0VKrM0au7tMNn1Kd33UvN6YbfQ
Ci0wiTwu8D8zbbEhZ9On2Agy8kb9xjJzywrDisbRr3Ca6JhDqbdoOA4MAjrKdkEFqUgT+BPRaqr4
Yuj1pmLM2lyTs9MhVVLCvyze0kqrwnwcWVj80obE5KDSQtybmfaRScGccY/7HTRsClcp5z2C75MU
SkY+x90lO13QMs+iBJd9GNc4Pnl1oMhF8agCYCpiZ2372kFad9/9PKoaLhHUD+o3cLffbdSFNcZ/
wxqp4InbCQPXzcxY3sEBaQfn2ArH01dgs1iclIJ0nLMjBiEgG2FwawKwfx791ecykGbjjDKOEO8g
lkzvB7WOvDrLRbClP+IpjhL+ryuC2myvOXeQWRG7giRxJgUmqKb4KqsCoLXtRU3CZ7oPINc2RZbF
XTAgO+CszFNIn/AdnfalJ9sr1wNOgqGZLRQP05QQ4Ng9at6ftoX9if5Ot+rzgxb8XEpnpTkyQeoG
MKPEagL8YAPWtznmkS6ybq3pHMw5YpauD1s8GiFo1tcWc4TP/40/FwiAmqQCDPxafPrpqdLZlQKe
Pf2yDAw2iG6bDevTz9oU2DomoCkM2igjS8DZ7GGSG0gn5RTFtkyAeNkSjHdB3dHwkdfzyvVcn0hy
mjjzF+FxOE+Lw7gGO/ZwbcB4z+PrAe2YY+qmRoLxowANam7iUKite8Taknz6UDsFnbtQrRnjV6kl
3kcYHxILOdaqpA6BMOJeG2oBdMPbSEO+C5AYajAfsMv2ralaYX/BLkGKXS48VXeECu2SdrQyULOQ
oG2mhbfauMFQzuFaQenjxgyCSdWP/TDAWutoK3ifkj/89krMhDC+ju14rs3x2K/ierW2d1MP07ST
MUFf0B8/wjJMFlbyUm49162MBifrRATbIiYxC4Ho7auT+OKNOXvAtVCRnS4s/nl92vIAFyV7x6vy
fGtdZ2xZvRcPt2aWFRhxXDuUlh3fab5eZKEdxdh/2aZJnM/rFv2fGpb2f5LbCXd1nle3XeEpZKgn
r+c8V5LekPNH4M/uw8/qRkEh88Mi70cPFRdVmtLhW4R7NJod1P4CND8rQG0qqFOMCO0jvdmJMUoD
R1HKbBQWPAyfM4fbMR3FXY6+y7dEUpMXClfNnNnLJkFujCxk2SkiG4uh5GwvneHlfCQp15vPye9p
eValQOLr3BAVurLzKbxoZmhW+olzb5FvSF9ba5VpxhDTaHbmdhvBd/9viJpwJrOtns+qm087iF7g
Pdfn4ehp5itpSETscdjSlO7onL8+xnzY9KLKd4Y34r9rSlRsYl9TWoAEVfDTt2RLWIRl3H8nX4Cm
2e4iwEOTf9lSy+NXmjVBTt1E63zqerTtsD5GmaULfATqkwIRIPgHBzk7NKx+mOiQXasyLbOnJonO
Eb9vCobz8jkpWWiDoVypmRfyJZHZezusZU/r4i31SamERax6LEkStay+35LJrwR3YkMOhDIc0z4s
vCHOEqPPrrjhZHV0mHynDXN40aZn7atg7UFC3ZxCHOn0DoXIvTcvdHKk0LykcZUBWvVLYIYo87m6
od2xJsuUr8N3dnRWeMa1cJ+rUYlty7rkph6zXZxBQhZH5ztFgbtnxJSejRZnSLA2KEJbcbabPS2M
XXFlnfR31qoz7IDvOeopPUW7sbNlgLGww7kdEXyP8a5acn5ySCnbByrbuLOCawyGaFmMW/Zxd3Ph
PUasnd8WhZf1QRJBsniopiDo74aP9J8CbGiRADCIE7yjI7KYcBLMr9Wf+Ml06OYnd6XkEeM016K9
6FVdo/fL6eJJAbsU33soFL2P6DsJxpEE68tqlFwZJmPz8GGMO6w4h3AtAPU3aa9bDWOP+S+xLGTw
jVc831Ufj2PJsoorOZ7UH9MtwBpq5Xw6iOf13l+GD8FyERm2MfEdD7MNnIjIAyqRAAhBCy3vcB+h
I1gU47ULNqqcjKkndqHPi1ZG52WJOjRpoWQl7TTLeAQtnqDNaCRvJmItxn3BFowIm/jZ+4POEBZZ
+yBy2RACV0yT3B5QWHWH48FbAo8Pp+RaVKuClM9AHyXJE7iXZ0sILokrzHh7A/BESPt9XSDceGOM
QMmOclB8u/WcEuy3M3j4U01LuPKqWWBLJjK9y2Y/GF0i8u8pRGxWgIAZq3e0yweByu3aw4p21/pW
7aoIF0o/5tB522LrXMhmSQ6JEcC7qBMmd1fO9Rjkx+E8xq677dAp31lDDCH492IoQPWEjAHTWH9B
WMK3WygbIh3B2TMOflcnnTFmfIqvIN8PN47nDgLpDiGJG3DWbMKxgdqyd0dbn7EIvA1ZHl3Zi/FO
Z93lykVakXndqpLiUjKn+8uTbaXDl0Mu2rIhc1IXZ/TqmWMrGwx28kdkGGAgFI19OfodYZ/dfxDk
Hp8+20FwzdTtM3WQi/5w//cQTPimcGX4rO5koha1bXzP2ozQH/YWZMMprsAyNjsljdhTYcONQWLu
G/JyxVUwH60lDtJEJJhkstliI6R4HuDVDFBNUbd5QzhcppFx4vLd8Bt+hODidcDK8j2gaoThLZDj
Br7zYzvFU+ZdM271djlZ8fskAaiurziJI4tnu1uht9//uSQ6moFLKFKZprFq4Cu3zFdtEQAWY7Z1
o/iPtFrW8IgGodUeWKJ5cPZzwFtFo++cRzuONUL8eKJ6yPc5MrZto0H1dksLUrOf6+14KgkHe8VQ
H47stZVJ2Rzpu06IV2msWA9HxBYfMiaIl81HcFQpH9HmEZRZguP5su37dObcI1W8SmwR8mrbpoKU
m3OqqziUnmjudmYRxhGacPPl2cxAmSBBelUbDvFaO90j5vGkdmbA9a66SPEvvNAupCjH0tylz//k
ukYk8rHcDGM9YIfhccG1IYF98pxWMAbpH4lPNBGfN4qRP85PP55j9Ehsm2Qs3nN538+K9xFBQrFa
fjhstSBfPIeNtYMt/GSGjLFJAfVbuk5KScDFc7c0Ug2B16xoXOhg/2gopqDc+P5uIal0ziVLa+Cp
qjrwOgqdTqKgg40BHdNTMVXAqkJk+AOKptUevI5kC9qZzuNWiU/HUbZd9KPnAds1jKFFEFQkbpxS
Za5wcs90a2jKJKnA2BMltraYrst6CEiRf8nkMWMUaatXlbUu43BUwhWQ5KWCMlxBlYF1AQ4mE0wQ
llT+CMnLgwuPPkAiMXoRlNE1mkv+M+EtCBQqKXTt31paiKsfWLBpX+p/zuCpoJeeCHYQeomEHJjZ
arTe8m27tLe4aNuIp4jGNaOfIiyBQJKU50p08ftJGf3E1JQqxXhYAxFZMDkBYGu9xh8mMmrqKhvi
O3FxliozYrDWVzZAEPbFKAxQXY2Mu7tfA74wUwX6UUseDjCIQMnkFVeJgumKIpCaBrgEDyKEHTEY
CO28N6bmV0a0uPbmllzzWObZGisuq6H5VAqrD04widLpm4VJ883NWcjsJBbLhkScj4R8yUMtBqdf
eUc+dEIJe1w/f60rGjORjoanJW39PhUYva2LKjHJ/dDr76UV/NepKuFDjDV9+rDiUJTovjTE+t4e
Y6RBbNxteefQfbc4//L+jqAhFMP52xX6TMynE3HZxhzZg59Zyg0DLI2zu+w24EMF2hvacYLchJcz
a7BQmgTO5GO/dAS05WIstzwsMlVokVqgG2rENiAbCmfZ6OU6Ax/eaL5iVl6RdgRlLRd+ooKJEldw
S+Kmon+Rvz5+xtLVj2wrrXHtFReD5V6Zh5bt3K+oXGJh5qHd0kYYwUlc739YAzGDdmMTowHidz7E
JReE2VdRJq77bUQoAwc7cJggFzz0TCpvfZ29M30ETILDudnBES0rjFSUT92ChlbyiqbTCt3K7lLF
XMKDmSmMMOn+D04P3AycxzLCv8cmzcYfDpt8rqV9Xurv29+ISdcl8uNpt55P1FAlg+8Fek00V+ma
0Rn54s5iPyBo87dghoCFDB2JrYIAsh/7JXeg2MCfJaMKqh2AhoZjWksuzBnhU8drdddfdpX12Pco
L90Kpc0sctdHAS2mL7QJj6Hs3lrQYc6MUK0qwj9yXXrn8XMoMatZUY9KYRYiNoyJDbOGySGslzMz
h9J2tRMZna9UqnCycH3kMzNWZphz9c9/391LR8tTIhrs1xUCplb09ObIeVv6hO8dE08Uked4KIiB
QhVH7gJODSTrd55hA4IyxLpfkvPNtOefhc/mfhCXkpeafmxmLbBinNaqd8a84voV4MbIBHpdN+UE
BwV9c6ijGHXXRE1JtT1Vt2DN4ZTvAiICTgTOnm2Ky/cyK2cZ+w6wNAW6Z4khDMmU07NqZenimYnr
FPDaJHS4s5Upqdh6dN3Otw6kouM/0iAT+tMb4Fz89d9+T8Z0sg5DUQg/XJUxz3V/qP9ZzWYzPx2w
IYKCCAbW+QNjZvEDAZvuSDxmCAE/B9omQ9edldGFLdDHt8nP4NyIKnmebNQUnQ8xkjoxbNNjNXYX
TMDTmmd1CIa2dXKjEjKF9zV95XHAao/A7Vyhr6YQ88vgaiqgq2lEb0QTAl22jeA2Eurw1Sc9K7X4
eNN4sQphTf/0NTiTTHh3NLW906WEs5aTI21GLY+uHzv9OSe3RNyJ1Ajbj7XsfKywayrnsCzZ4UCb
guYcy22u3DW/Eh5RNIoRsdF/RInUnf7tBnAXGMmkstwyAso1WjSqiQ2hhVk5qLauF7LTUWocW0cP
dgexW+BfGRDi0zr6UQZ6ShQ2fkJWzaOX1cbeTB0RnaedQQf2Oc4ex4TuZjLvxNv4Q+7MrDJkFB1/
5jZfzYB+Kdhs0vi1obSCsaVtNtoJCgmZGngfMAf4eFxGC1JpVDMh5vsH0KoZ9qGMLwcZ5K5YseOT
eZomyZwbvGO4D2Y7g/fWoLxprvXExAh7kbLDxUMpuX4/jiMXH8K4gI3SoRG2FKTIzQgBV+P9Rzs8
k3jmpQGNv2GwnNIT4meoxPJI8Wo16aJsommv7p9pmiyGWL6wHlntAG87JDw509WtRLsTE4iMqcp+
z85S97UiJ/VMTRWoPGZmgSvuR+Zb6TQWGvj0aYmTsc1z+WrVX7ID5cv3/uJPBaFHNgiIJo5a9F/C
1LMI0uFRPpfx+MDp22IoROJeqSA2gGeJPnhfnmuR9ep/ecAYny9XEFN/hiv8KsUAJR0D0DleGBN0
kpgdbqaLJJGkEB2loDPAVv8NpmIScscgzBKxnjQ0+tCMsvwTqF+n/dVbRec+CM382ws4clFVNWFg
m1R1hnE6ACvi4gHI273liWfOwOIB/xxQnA4rf7iOLjtYIgFF/O9MhIYhaTioVtQ0Z0Q2MrTk7582
YjJTSOr1CkE0ch3VvSEqMvAqn0NkQKENwwAY5X/N7hrip+/IdmngvIS2C1JE6Hc+nUbE/o2KQ24q
dkaMfVHqO8cUOPgJrJg/Vk8t5YuUMv87XggndTiF3tAFHpQLUMdd1U1UixqFDTL1lOJUxNYcWcwj
+VbvmWZvq5akFcBne1no4lFws3Ogt1jdgnZ9khspK60avjYpZ8j4GXE/Urbb4Lvn6+YeU8F7GM9f
y18e9t+gwevyqHuhRrtrHNBq65qVLnXo4YG+eY3kvUEbu9lhQvKRscHeXjAoz4O/dBD5O1LC2bPl
rIEIIif5jUrnDgDd73Pck7ej3/BctjdKPLXhGa+FZjCxpYZjJ+WFN8ylht9ZCJls3/KZNNKtsS/h
7ngI7mxrxMMtzZdEb2+/7Ib8plUlprVguDFREauxaGcCw1o/LIPRGSq1FHj1iu69Nu1d7RMpRAgI
fmUznIvfIqSnYIUazrVlQuWIfhRmn73STQ92t3qwVkIsMr2Jb2+xF+mXGE1Rj4Ow68HQ/nFivklX
ZI+70Cgk/ovCnI2TjyhU7ww3kF09V1CoQ5H4EH3niEdPeNHG6tHIGC6dWPquHt7ZMeMff+BntItG
ZqDaT964+Zcv/iRaSt7TZ9g1KF0QCE+EEbzK4VXFb8tEmKH/xMSfYbSeVYczFNk0iG7ynlxEdGsk
B7Fxxxsmh0bUJ7rIySrpoNkaDW4F/dKwFk/p6Zhz42MCMThlLaAiSe+iu0brCGyxXqhuDBZRlwEu
gYaqg71Ixoywvz9bHF8pdCH9TkM5e9W68eVW7cp+9iNAkmivKF2vmoZMnEs4J3Mrs/wzzFShOcMI
j1/zlpJcOl2c25TSUZLGJMU7/K1VJPRB59bqiBC8VVSRfb4ZTd0X+UYggPd1lq0cvJHpOvOebuwx
LRYG4tZeTvFsrQ+zcROLRwYKkV0Z8wTenkU+cgT2LZTkClN0RORUZETxyfJ82+TUQ7AsJdEDw3sb
G9AL1AxCiUidJG8iku9hfh2AAJKYGbqYcTkSwlMC
`protect end_protected
