`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2448)
`protect data_block
0USWSUGxovGsyBJteYpEobCIoMYi+tILFGIzaJMw/o3UMenGdX/yveblBx0vXISifigS8ltL8OFg
RPa/D2WWrEp2BggyecqMLxalc4Yn4CEaUi8rPncnXGf8dcv8kdl9IS2etxlzR9gv7EyMeQnRMp2a
lmuzDQb4ErO9YfoA0kpUnN2PqZmyG/pMtd6ABvZz0Xa2B8rJnaiTqb9ZDLCe3/oIZfuADZsdVbss
x2PkGYz0G4ECXcVX3ZIV2uli42jbExjv3y42s7NU+1/GjAc7OJZUQmLHRKuYttoXdttp8bye4c6I
o7Rb+XOx7fWT4a7DYl0Tl5vk48rlHgyNxx4p5YKej3Ktp+pa4ap44KGzU8GWqKkq3OiqTnUU3sJz
V2fRnUonpC7vZp1ZETrFGNMLFLUUEDqMyPF3ptaq84WDhF7PDQFLuYbDU5z2jv45238O5dPXHzie
gdi8vB6PqX/5RBgotd9vlwzwk5cFntYjFwKBTJtuvqm/Kr2BWV9PkF4fo48lxZpaePWgplBA/qN7
CbGj1lFZezzh0pUsqtnZuSDs27607LagcHctb7fHJpKAfxNap2aBWF2AjvbhFiMMm4URD1JC5Kfm
YMKclRNlqjj97wvJqzJhxIAqjetIaciuzP8nm/8GSlSVnjV5Jsh65pxtbpzvCDT9UYNFZdao/rmr
RtXgzCR1JmdaDZBUPaZtLtgKlX8TIkqAaaJib8qOYLSbdkhGZnJa/kICUECDT9PrUxcJhacL9sul
+UeMhG4PiLLaZfhOKIS+7helLZQBpZsWQElrhIJAdDZ+WQLoKzsWVnhA+RdItIHWC5l1YKs596NX
kXAjTux+pe86KRfb0m+mp6QIQZqv9UVN+JnyFGA+lieSxcqwGmIeLbMC2aJ0KVv9ZD2ov5UZ2i+a
q4lJbpsj5Di8INU8eylrSpmw/LWjBTCtZHq2EvlFZtWDnyST78qwe31Z9Ak02zzJAyqESDz5bnF5
ZoyoNxo7DxtkhyR4XEjKN94a4o2e1GbrJJon8FonEtEeFm17OxnqbPjcFB+X0Okt+vT5heIyVIB0
j8QZft2XsIZwzFNxFlnlqR0Pon01pGPkSt1cpNh3ApV0ZE9sPqYNol+eHNW7rbKn3uqiwd3T1jwF
tw5UUeQMa7ZTah8v7Rz/83UO4OsmhX9JEp/SGGFwWuCNj8XN5bOMYTS5yh6SPvZgnj5mjjx6nFsU
kFfC8RLq9nU5PRE/GWaGv1wKaGHZqt0pVFzTquN5d8yp58pB3zn7o0F+8/oUu7j+cdB++H9ij344
OW6mU69uZ5gErmU5QhOMdTHpC4lhiRxxvYtKZqb7x5B9Cn5djsWItm8HrjJXhScMxrCrJ06kFHum
WnG0NUVfFcjdxjnK9qh4IUfz5Z2DYWhYtQiHLo6afW9OJU8qTaZ4eUHeLolx54XRx2+W/D/7DlJ0
bu66nUrFjAiRPm+6qZ/nUv5ORtjbF2A5+TBOaPrTbdvGM6NIW2MpO5D/LSdYTkyU/WP1Uo+ez5N7
+GUi/LDdMCP3SB0vhqVz/+aMT/ao/DpUU8Hn+/LM9Ro60dEJi8Izecp4Mh22cUQf9+D1kOGWUws5
o2HBC22EyK+cECWJ0kctlaV5hrvregUvavxz7lGj8Gve/2CDGPs6hvIe030IYcd5T8wayJm27hVL
2lEXNHORvuqjNC8TQ6485JrGkRvLiF8vfCghEqUUm/vWN1pOM0CtWRZ8uR0sd9nfTziOLXatsjUC
UHkATAMYi+G8thuHScgrvJzvT/1qlAcfX1CNTOFhnLxpPS18SlZZ+bS6jxAlGh1n3zlpvOxIf7eX
453YQi6i9PunzdFuoQo7XDzxntCexa1tAD0p+ogpP7syEMh3Y1/CIMnSiW38b63WTSuId++YOTda
IX0CWlAb9dQ+ipasU3V23E8BIuGIA4A2T92x06gygB9AmTV0rtz3kcfcE+VuULR7Oidqn1j1w8W5
pdmSWahwGNXIr12B0PGByDVbkIXCg8U9yK7FNf+1sC1iWbcwvxCVHipHyZCExz90fY3A+cZcPbem
tWJ7lEd9p1kqTyUiavfzcXxgiTfISEqLOvOpNnt6m3VhmFXTbCxMk63WGIMZw05tI7/9vqX1CCvo
vK26kmSnjyci8AmNXiZ8jXrjH26NAYq/J8d843+gPiQtdM6iTzdjV2p8swVab4Kf80zSUEBI4uqw
RaTmvQicyIfPVceiUtQuEMZPHqa9SmMepRr6kWeIOzK/q23IcZxn7JGPPZ+UdzXBoqUZ9zC/unS0
jVWlr9JdbgIYyh0Ej/LtDO39+vJ6dgYg5+qBXMPCiOymTE2FuLRhE+FxOEs86L94h5dxTzBnrekG
AgM7i6Zx8tauoP0bpfQEgbNRK2O/S/F+QeUgdZoHos1k4OA3l2OOa1sEIdPkYNhBWsaHNJKKQ6Oy
OMc4RYg8cXO3oE0vbXcdIn/V0jtXw9Q3098U3JYg2tGqYb8maMscST0I54TzQ8MNSL+rcNznIX3B
3hWXUx58GtyOeC4bpkKQ4I1RLxE/fYY4nS+wul3j0NHMoxZVgZOjLTB+yOHQQNW3XGsc7cGePLPr
BVACctP/BcHbKk2njfydTZ54vH4YZR4Bfmx7VumuiB5IZi91TKzB3qbOAUuGs8pCTnMjkPNCLAZF
cBVbFjIzpQczyAgqiyhurTjei1asAQf0R7GFbX3rM1SitaWLjjB8odMCzXZMgSxIfjAV3Fcf3up4
skPlSgGIBLZRQk6UguCmkdDLd1MqPGer8MNrLZWCQlbg5cEcGkD+sKfPH1/WPzUM7jfs6Igvkub1
oCNk6MMlvbJCzVGrGyExG4B3iWcV2dINSk0KZwE1JtVwsN8jJ5+aYFJurcOQ8my1ohNXFVSaZAqi
x4WDhGzi07gC6awylk0Pmmrbdd4gfYi20kqJAuG757nJcAHfrRVIx4K1kz0MzX1V+M58NBqvQS1N
8a3f1E3RdZliVWcIsorxup+Xry2aslx/tVZWo7vBZgfB9ZpWYsHcoFvW8j5+hWety3zHlCYXdWet
1vCRYhZfrMidsQmeXQIc6px9QUi6zq8+iLuLSo9RcT9WYRLEEIgSu/J37oWtzqx/mfHoWP5VtYgV
iCqGXUBPAyNWYFhgJZgBJN8X2ahul7LyzD0f/YXtFnE0TLcYL7gRshrgW+PRStBz1Hu8XDzcmlra
R9HSkVHMq4/E1izbaqsWpyAteHjkuj7uofh3vreAtxrOZ6mtAybkaJESgDa7jZmInv9kyh5m
`protect end_protected
