XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��.��p�J�Q�^�~oI�y�����xYM�&F7[��\~ �T����VȢ"�@�-��4E��Nm��o��3u�������3�t*(����r�!���n��$�xL^�f�}��d��_(�XǤ�ب��rm�t�^�҃,��!#�������7z��O���u`r�?P�}��1�֘+�eZt��RV�W���E�nA�g5:�ˤAGL��<(�B�W�lҊ�AB{�勃Kr~EGŘ� �h�Gq�U��,Ey�!��paC|�8�MQ�#���Q`$�M�`m��+ޘ���1!,gD��p3�`���1��="�#κʴM���~T���[u�Əy�|�Aj�v��^��՞�o��`n-�o�S�	��:�&�YS4�cEE���AӪ=�(j��(�P����^iC1[�"q�;_����S;�>�,��-��,3k���`�{U�����.�p�q�����v��<B|���4�I�����С)�����-�%����"����n�M�����k���KEʋ����f��=�__H����9㰵��t�p��s���U��#M��9>ŨE�io���]�Iȴ�#���o����Z0��%���O>�o��ڜ��)��^�C�!�?G`���-���L�������:�`̔�W���ӗ���~��I����t�����
Sy�N80�4�S�־�Ҿ Q�����f��U^�Gc)�a�A' 4���t��T0����"���o�TM)X>�;�x�R��R���XlxVHYEB     400     1d0�P5#�LU:��r�ُ��J|u���M]�A2�2�`�r7��uJH���T���}�R�ƺ�a����S4����L�L�˹���P����)H���쁐^�q��|����W�1P&ϒg,6@��Ki�;���b�L�Hͻ����ʰ7��@���A`{�N�ر~SRZ��Kb{���%\~��Y��J�K��Qj��o%�;���ˑ�s�O+$bh!�45ف���ڠ}�s���/�ϦWW�M2��=)U��z��/T&�Ͼ���u�t��apyd"�8�[����=�����{��gI�s��n6h��Q���6	���t�'Aߚ������̍�S�M��ɖ�*�S�X�د���+3�`$+���XV&��<Ϳ�c�����̆M'�k$�J�)�6p`A�)T'	�6���j����z#���v$��yGb�ua�Z ?�`K�0-��XlxVHYEB     400     110�t	Ae(d�Xҽf�ZB��e���Ej�����Ȳk��j��9�����Q�S���ҹ�/6�����m��}���I?j�B��������/h�/&�r�,X� �xoob��rQ�2eqx�v
�|7\Waö�#���5i$]U�0m�\�3��V�hh~"K�&AN�~�����?���5�(�2Y��������X�J���"RWܒ}�Y�)I�K��s��*�u����`袳��,zޗ)�5��i<���/�K�~�,�Sj�XlxVHYEB     400      f0�ap��e�2�ȣ��������)��,dtoEq���p�a��깣I���X���~e<�Jm$����\����A4���28C4��s�P�����J�1���-��,�':Z���~gܨ��P~r
��Tn�ה_�^������]\q�EMM��R&����T��u;��U���4��'Tv��<�Щ���URp�Q�e�����/7Vw��笴��u�kF/��Y���(Bk�;�XlxVHYEB     400      b0��L�/�(U�2}�:;�\����J�q"/���3c��=�Q'�ы��������&p���c���q4/	��Ȩ�7����lpvJ�]��\=n���'��5������^�u8)��(.�ǱE�q�u��Z��jhhֲ��a����<p�r���$17��S?�Ʋ3w����|s��|XlxVHYEB     400      d0Dq�tA\��r:�����ɽ*�����H�fbv�
��������%��pSFm�����7��EA��>��\70e
?ؿ�g������zz%vTd�hE�I|xS�f����޾hl��N���+�脘�v�s�R���M�;�2�W�g_����˿R�%�����n�]�Kg9�K !#p`�E����&��T��aN�XlxVHYEB     400      d0N����/��v��O�����/s@�.Z�$��X������@3��뻤黕�7��+@�#xe_��g�^oq�Ԉ��ˁ���{TE�J�^�y柔�g{s�u�� k��.�~��ϑ�GQ��3{}�)~�qT�I^�ɇ�Bc�9�Vq_Aè�z�k���z2�H5���YE�\y"�@��#������?Y�-�]�5�XlxVHYEB     400     120gI.�y�!2�75L^ʾ~�d�`�ʦ���^#����.������t=��O�j����E��8GDT�tY����qjpа;�xa�!���dr��4��Z�$�sz�WUMv�o�y�;?��ծ�pQ�z�K`]�3]|1j��_��1�R��ڰ����ޔ��_H�3����l��g찗�a A�De���lk���Ax�J(�V|T�Բ(�4���wd��4u���v�PyS	�>��w�����wq��\YQ��4�,���W�d�c=IPan��J/t���:�dp�^�0XlxVHYEB     400      b0*>{L�!I���j���9pM��j����q���Sc��t�`z�����2C�g6.[ai��ǐv���t2��c:+��M�J���j�.v0:��m����3��J�-�-�S�/M�V��t���;#��!���dbx��-��h@GP-6��+��Fv[�X6����ˠ�~Nz%=XlxVHYEB     400      a0�Yu�,\q��OzP}H	�l�,����ui�{���\�>l[������U>��$����ܡi��W�c_ÿ��y���XN�- �`�s(�x����@Y�gy�fX�,UUDz�\��x[Zi�z���)�#��>E�ʚ���ְ%�ۈB�&��E���B&;XlxVHYEB     400      d0.�y���m&CmnX�ʄ�V*һ �mD�S����J?��� N���P*چ��* I�=���p�r4N���SB���P�߶�)��R�»-�q���"L2��dէ�6y�ƈP*����5۱��]U:�5��:�Lc���B���"�bL����qϠ�.�����qu�J��`t_���^���>:�:�$�)���ݙ�J����XlxVHYEB     400     180^(TA �4_W,�z�,��:�L�6�����C�56�.��š��ƽv�\l���P	��@��LḎ������\N����e�OUxͰU���BnL�ɤ�b��ׅ�_%�VUz���c8��9�c��t�txI�
�f�}����*��Vd&I���kU�{F�T��d���`�	�j"�!�>�,�	���D��ц�9�ʕ��m�^����C�BMD����P���8��]|����j�LIc�
�m�����(I|�58��W'���h\�C:4���Q�J�uT2٢���6�VA�&E_l_���8$K�72!���+��GAo�Ӕ���Ɇ�s!zH,vvż��Qq��Oج�������Qg��.z;XlxVHYEB     400     130�p�
�X,�A@r�	�E�V/y�����p�퉄X�5K��ձ@���D�Ȍl*a�N7E$��Z�Y��Ton=���f�5l�t	�� ����~�v[6�3A��T/�	`)~&�[��5���;il�2 M�EF��e��g��Ѕܹ��@FT���I�]03�ENxy*�In%hWw�.���)M��г֝lUue`�[�dY��(z3�M<ר�F?BY�d$W��=�EWa�-�e�O���ݡ�B�@r�YT�ꅯ���A��:�@� '�V�}s2��=J+i|�~N�A���K��>�oXlxVHYEB     400     110]�FCo�cq�|�E��H�=����pn��\:�V�-g���E�Ca�gEe���n�e��I���!iC%�HX�ݭf? �j���˗�%࿒a���¯���x����6�*��L�!��T��,��b?���t��ɳG�	B����o��Gq9�fŗ�*�1^��BD�`���OW\k�a��uW��T�Ҳ]7p�j]k09}� �{gׯ�B=⸠�E�7���:��2��)����T��C���Q�H*9�����J��M~��:XlxVHYEB     400     190T��.��	fo��:L��,{	��);�e$���!)��<(�39_w@�AҭXx^&{�8ʎ�����V|�N��hOw	�G�����b��p���6�~0�	[�I��=��Y���۫^��yd�CL�*O�}��a��vqUPZ ���
a�'��9��ńf��%��'��6�����]�C��A<�Ɩ��"��	��J;2Gs�h�ɬ�ՙ���qlX�	e����9f�%jr�,���
̕�����x���-�؎fr=X�,px��]�4��Л� ���V���8'�݈={|�{�!��p�xmMz����*ս�MFYP�
�HǈS�=H���C?�	V�!�}���V���x���_�"�W���͠�U�,�.F�S}�Cx �;XlxVHYEB     400     110����E�pg�d	?*��,�R�'� �����`���`8I����-\��^G�2�f����'մ��_���^�+wa,�8>�Ah)ʡ�Lڷq\����;�\Q�	��*�������&u�[��-��	f�^�n�_b<�E�n��<���K���&�k�����R��p�Q5�Rr�Ψ{iMV�>�|�Rs��Z��[l����T�}�Eƒ:ݜ�ĝ�F��*�(�9���T��6;�� �;��5Nօ�:?J���e���ع�NF��������XlxVHYEB     400     110ɠɎyr=1�;�?؝E���S���&�J"1����ǽ�sRJ,$x Tl(�`��9ֹ�zaONA��0��uo�(���^�K�T�:�y�Λ;���3�h\��x<Vn:�o'�$�0��[�b�5���cul���F>5��/��ü.+Vt�-֎�/�?c)��}�t-�ר���D�'�� �Br����9YH�K�+&����).Hw��y/���OH���)�Y%����B!V���� ��9o��;��Ô�` Z����pXlxVHYEB     400     110�X����h���-؄I�*	��_!LP��<�w���YG�@ژ�P��wv��)q��������9�=�v�.���ݕx�K?D�ۃk��ǔ�#�b�$Wt!pS'�_O1�Y�����ᯨf[��{+��"m�I���=?#ȸ���,�e���qt���u�͘�ں�Ru�-XΫW�c*�zv�R�%�&r�{��f��R>+ +�gHn���'g)��}��$���s@LȨ����X�W	8�����`*z�TW��:�P� Ka���ev� �_�XlxVHYEB     400     100M���0�4_���TW�����i��r�H�;�c�uI��?Q���E���o�;����#�Y/���	�VD��R�wP�Y�9>����(��3KYRs���Gie{�<�� �����;�X~ T��bI �m#SP�i��z�ag�^e:lj8;��;��a2)�鯇KG޲ma���}C��L��P�3�����Xx��B��PQ�y�q�X��R���7'�{�c'Id�u��}�M{��bp�m 0���F�XlxVHYEB     400      d0L��0���&�5nnX$(�+r����ʽ��u)�v�> ���ض,��2�@�M[/�2 �$Ӳvq	�GgA3�;M3}�|#O"���`���@��p�o۳�B��1_�	��*�ne��j��~�c̓��K��:���$qdh��\��3��B�E)���ӳV��
��yԺ_�g�Gd7�' iN2<���@`�֕$~"YdXlxVHYEB     400      d0���]�J���l{��Z�/6c`$J��m��p��D��<k-�a�e�H1u�+K2�gw���b�s�M�ߐ�$�޽SҶyՉ��\�O��~
1�e�� %$H�r�C�1~�P�7��k��������Ԟm�e%%`zx
��F7�n�hUr�K�5�q�2��V�[�s����ݮQ�p1H���#��J��I*��� �֧�D�}\��XlxVHYEB     400      f0�j��ĻK)MqG]���Wm˓>˷���/�y@,��ե5s ���u�3r1�F�Ǻ�?�}r0�Y=:J��SN��x��)(�����^�b�i�D(�\�N�ȩ�yK��XW��|{F/v��k/I~U�2s�vb�^*����{H�萝X8@d�K�,ؠ���X�XߊBW�aU��L�e�bQӢ#QCFjqqU!C*]�lq�E�S�k[ל�^*4�eSґ�;h�(����� -�XlxVHYEB     400     160U�T���c��J�*� $��L���-�����^m���j+k2�r>���(�4�}��F^6M��,�}V��ms2�l�����!�9a�eF\�T͉��-ž ��7;̎-�S6?;Ȥ���6\�dlvi��up�r�n�W�7zn�fE7@�Q�����H���h��Et�41�GT�l��d�����B�-ZJ.,}�L����}�.����[m��C�:'�����VH"��u�z�S��c�o�X�ML�kyp���']��s����wd�nV���˕|�4������js,�DgY�OJ%GT����5����o������� �P�����
�XlxVHYEB     400     150�P��E�jb7�?�-6(y�:��}�K�h�c���ӊ��P4Oc��=w�*�P7egb�u�/���&H�����W6SjMr&�?��/���ZR�BQ�'�?����/"�֩Q��0ٿ1r e�a�`SI(7v��2�6��8bB��>S2ˍ�]	t��坥�^���V��3;T���)�������:A��sbT^ }2�eg�H��w�����,�Xt��:@��p��r��ʣ�0YI�����I[�����O�NL��W1�vht
u	�а��{ܼ[�Pe��R�~��4�a��\YoMfgBt}p>q9D埜�j��bt9�ޭ1*.g�%XlxVHYEB     400     100˕���Y��x��,U��f��#��f�Ad#����H��� �*-@mN��c�1���O �W�4>ؾ4c���*��fw���|��y8����Ql[��1Yo�GDM�H\�\�b@������&�_X�5�L(by�|���S~w��a� �Ȇ/�!���60B��S���%ą�����U�kY��TQ9fj-�	�ƎJvu�T8�@�o�?a�^��=ޡy�ĕ�3�[����R�c�J��
P�xS��YXlxVHYEB     400     140%Xw�����|v�u�u������=�Uf�H�ai�
YG][�0��4ye�P/s<͹&�;L��K��l���fI�P��@���A��?��O���-�w;w/�@]8��BU�F�x`Q��~�߸��~�J��A��>��4Z�1k���m�NA��":2��Y3���/����0 ׯ�ӡ0���/,�"6ڌTATd�&/>�J<'�*��!}���&�0�>��`1��w}l�X3�d,��
E4��Z�d4�nkɯ-�S'����DA�II^˞�q��:R@�37���Jľ��7;���6�}~|K��s��</NXlxVHYEB     400     140��uݔ&#3 �Y�����Zvx�R�B1�w¦�]�+b�-i6�<N`��i�̟���n3f��CQ�NeN8�3��*�E������a�*�������i�ܢI����+D�K����݈l�K��%HT��qh��ą���}�c��8~ɻ0�_�_<h�6W孮&�|��H�0�ɖ�Kn҈�:a���l�JM�i�Z�Z5��������E'ij�t���U�n�n)u���ٝ��f�3{Ft�2�Zj�}���BCϱ=َ���o������%W{�:�N����֪Ȣ@�|X�1E�?�c �E�*��P��V+XlxVHYEB     400     130�ܷ�K_���� ��bI��Ws�M�g5l���\zڋ�6FK�&��(��cGB_��$��ӡ�jc��p�z����]W�U�'�؏�wn	<L��D�ʬ���>|������G��W}�(����Jj��>����/��NT5U���_A�׮�
PR	��?������:<~��`��@���cn�7��71Ra�4?�|J�כ[��u@�؀���c�
+]�PV�$���+U��T�2Um���0�5����gڥ�|�ǡw�	확8��Y\'���b��i�<���%�a(����.�XlxVHYEB     400     120 M��D�8�7��?���x {,���w��\��.���6� Q�h��{
T,"�!"�'�;�Ç�I��a�@�AW8I�5�Ӏ�Ҕ��'$/����<1�^n���ZrO����r��MU@�m�|�B�b�Y�c���
��9j�7�ϻ�� �'�Q�OY��\i�~���v�����{�7<��R @]W�~p�G�j�pm4	�o�F�n�]�����`rgu�`ͽ2���a�9�h�|�� >o�:�bŚU��w5Il�xM�Ҟ��G�8풃�XlxVHYEB     400      c0�Nܖ"�o)���|����w!�2�/�;�)	�O\u��h;S%�\�����2[���5)8E6��7���E`'�Х�K�����܌���;�)�@A�h�����;�`��4i��7xs��խ4��{_y4�e��p�A��C�ien#�~D?�D́dE�]�?ǅ��?�=��;��"~ID�o$���:U���=XlxVHYEB     400     120��s���d�L�٤�i����-VX��+���]{�R5d$}e��4X�
�¯�1?~�x������݅�#�WV/��Ԛ�d��j�@d㿞j���w9�B��A��0���gW]+kv��Ρ��ў�_��+E�
�Ϙ�F�q���TMB�j�5jlr~^U�ΏD��8m�V�80�۱��n�f0Q���uǩ�|��ћ2�4�I�H3���"����''U=���;[Y�͘���iWRN��D�d�cb�v��4.+�L8�Q|���|�b�b�2W��6"5k�/wXlxVHYEB     400     120~N,�Y)5E�u ta.�Lf� S��ZE,�.�m*QK�o��[]�`��L�a,�Z���O͡;����ˍ[���
߾�A����dɽ�P�� ~�4q�l)|6�xE)c�V�K�ԅ�HaT�
�ov��Ŕ7��[2t/ݩ�o�aH���z�@���0n�U�O��4�%��ko��hXI��{�ѩLQ���YW\��]���^,jd�5���\ܸ>�۔j�fQ����@���0�R�N�愬��.��ɉ�����c��R�&b��<� �Eh�s
W�[ӖXlxVHYEB     400      c0d�3��qR�l t,��{ ������o��l��=U��ȕ6�����i�`u���l�w�h�L�+��4ʫ�(ު�}s+[�u��SD*�.fK�-A VR+�G�n�����9D}�c��}U�]o^���Յ⤸��<|�*���������N�3!1z����4��>`��՛�{]��2H��AD@�����G�XlxVHYEB     400     120�C� ˥��ٻ-�p���f��#�f��ň	6:���S�ME�����eN����b���-ס��YłH>�.����l.g�eQ�aԃ��
=���H9n�l��v�A9�H���k`��6�Q\\?ZG����������ܴ�E!tck谋9��
xn�x��l#�j��̆x�e����%�(j���Ӫ���rf�
M]?�A��3�;P�F̫��M{�"��S9��@_(�fS��u*�O��e��Eڽ,�~e��|OS'�B�{�b�h�`M�_���H�XlxVHYEB     400      f0k幐E���2s�sgBW,9c����R����ݺ�ʪ��:bX�O�f2�!�|�8��qܼ j��$WJ�7ķ{Z�5OҲ�2�FJ�����
\Z��Ϭ��^*�=q�L�2z"<�y:[
��O�Sx/�{},}��\�R�C
�I��MO؆�z�QC<��$��lV��~�=�\���&9��A ������	6ͽӒduE�р�73��_{_q-?�x'��x��i4XlxVHYEB     400     110@��a+��c�3���Y����6q&�on�mȓ�Oi�� �)]�U��� ̸��^��e�K��g�KD1�.u{b�@� �7��BŇnL�������0?8q�3P��-��	�t'�q+��r�#i������b0a\Ȗ��a8'�
�³sb�kt�����|�����ɳ1�Q̾�U@\���I�T��A���h�� ���B�F�S&�!�viyZpv��&{�$�p�Q��H55�T�C�c�س��E��?��h������u�^r����XlxVHYEB     400     120��@q5%20�n�q(��7�mn�٤�E�/�.<����d��[>Z��K΢>��?�P���~O�v��W��Jd.T/Q���u��6)!ڬ�z�
�TQM�{*^��)ە,�FKD���!Nt��fX��Ho	 ���ޛ�x�7���)I�ȿ�Q��Ԡ��q��qBQxѩ��'�3Y+'k����������F��b&���(M���]󡫜H��Q8M�����3�n��5t-�wX��jw.�|��S\`�$�8=�z���c��}آOq����ڕ�XlxVHYEB     400     120l�ɭ�1��m6G"?g�+%�V`�Y�h/s��	��q�sS�+��Kù�zUZ�������*�B�Hχe�;�:l뱪^�%B���m��4�)�UI��OU;���@B�n�'�#;?c�l$d�D�
Z`��C�{�PE�`�9������o��=_�G�"�h�i��ʓ�g�_<np�Q�G#�n��{���Fѧ��� �3���X�d�r_J���%�\�'qּBS�u��%��Rnd;���Xє)}�����ӞO��r�J�l.��t
��DZ�� �����WXlxVHYEB     400      f0�7h>�x������B��vX��1�@.#p��M^�	�3�T��,[.�V�3_@"���m=i���o��|"+W�ߺ.����������|!U�T�/Ѱ�YD���0��#B�f��]	M��R�(x����aB`�;^�xa"�WQ��IViNd4x�y+��Am���Dt!��:�nW�W:��);�c��c�2�t`�ڛH��ۗ׶8�g~�k?�t��k���!��K�P��D�XXlxVHYEB     400     130C'x�Y#��$??��|a� *`q/�=Q��b%j^��nFW������+�JqNc��7�)�5���h��<]�Uڵ��a���MQ)N���L4xcr
O�$2�qu�;�����X�w����^x@��B?U�OE��X�*yA��9p��aFw��y�-RX­�<�}���՝�-(��LLC!z#oN����x�&~Z���hp(k|G9� ��4Tr=�
L�6�u;T�ϗ����&;�P��G3���"����ۄ|=6鯀�Uj@S�?/`]���~��NɊ����~-��LXlxVHYEB     400      f0~��a�	J�y�}iԠ���D�x���+�-��1�9Dy)��� �^r��>rJ� .[N�E�4��w�o�J����6}�Ҋ����'��&��!E�֎G����ߤ��N<'I�$\'m,�;�x��^��5����a�Y~���z���o��I�_	�s'[��J�hMn �υM�::��lv�m�כW�'t_�ns�����I1�y��$��n�eа �Zƫ�AOa���48I���XlxVHYEB     400     150چ-U�ٗ` ��Y�u��ЎOh�}(/?��o%�ۉ�Yƛ[����$C�����x�h���}aӸv�K@�&�|��?��؊
�B�&7(����!�bn�\���8���B>7afgr��R5c�_O:���{�>%��^3�>H�YT-�Yս�g�g8y,�?��1�ݞp0'����{�^�]�֢<�륬mMFr�6����,�����+�W����V�#� ����H�9	��w�$9�Yq�$�/��!�Oר0%o
�T��b���(H�3Z��{X-g��>A��y�'͒�� .z˝h�;����ͯ`��yr����V)��j׿_(@XlxVHYEB     400      c0`�yi
o8��E'iA�
�Ze4/��]kw=�D��� ���6r��;�/�M�L9u����D(�-2��w���n��^�GK�n�l�Ι���6���)z�����UiKoج��z:��W��g5j�Q�zh�^�1J�ڥrV�;6W�Rm�&�p��5e����H&ɺ�?NP*�PȾ����\����.XlxVHYEB     400     150�e	�&Zχx� r���������;~�r��~�D[0{�����i�m�g@�/��ڏm��+�KPu�AӉ&��!�foqQ�z�O���u��I^�8�M�>H��Y�4\�� �Ѳ��e�%֦'���%�6T��i������oP��e���1{��ߟ�tE���Uc&���� *X2�
��n�~V,�x/���1�PJ��4�a{�E����Ʌ9��V"h�c��/F��$Z �G�+fw�YR��$e�wg�(��*����HCod��O�/�M�?��)�/),Z��k]�y����V׭�]q�s*�g��2(�v:�A����Bk��XlxVHYEB     400     140,փE��� N�d����Ϭ0<���������)��`\^^�F?�9��&�ﱼ1l=�h����c�W�f��f�/����u�:>Ȑ���%��ۋ[��t�=����Fԍ���\�%`��h�L�I�oЖ��wŻ`:�Ί"�f�xX��3��c10��	��:d8�o{8X	�A/c{��D�Bq�#�2�k���jV���)��֦�z��5y^��6����Z_�>��4�|��s���'�K�?�7�K6��Z�c��.��L���P���� EI�m��0c�Zo��B���4b�c<r�t�����?G���XlxVHYEB     400     100 �q�z��Ę篯=���l���Yĵ�A+@���A�͹�E)�`�Րm��f�"�����G��`���O���#�Vg�K����� �8�]UOH
r��z3v`J�(���eh2.�Π�>Ԭ<���*��$�O�&vC�g�_�����M������n��Ի�נuw���ѐ7��ƶ鰳=y�.�����6+�b�V |to=��ξ�=�͆���GUg/d6�F�Ro	|N8!Fs����šd�XlxVHYEB     400      c0zm ��ӎ2 .h�$��kY2�KT(�M>SN�����8��H3�ɰY�f�����	-o�cV�pm�7��Ȑ�nKj��u�j� Y#�Jr7��}�b�[� ���ψ�?��IY�������P��T�X�-O�%+~N̒*4MW��[Hϡ��5�)C�y��Z	��ìg����)�}�(D��*�XlxVHYEB     400     100Uy+��3Xژ���(A�ʊ�1�6�K�؍���x�'\4��``�()�|�ߜ��%�4Ҙ ��8X���M�IG�'̫J��ŭپ76��fil��m�NM�X<�2�����h�;}Ҁ��*�z�0��^���eLԑ�d
ӱ���������Z��F� %-;c���c��$D��V��Z��T�����w�p�F����!���V돊7a�Z�H�:Km��S���.�e�RXlxVHYEB     400     110�\������K�U̓?�m�Eo�2g慬��^󀟧�SKy�yk���L���>v�{ ���@9]�YI��)� �i�p{�o�F�bb]�'|)[����W�G��iö_
,h�Q�G�i�c;1�k��t � ��sjoTZ�t��gl\���-jh��ZΦ�a6G�E(�1�P��P��lZO�FKj�X��I
%���w6, P1��Y%6I]��A�����/_�%Ihw�wv-j��J����
Jj��S��)�s��7}���XlxVHYEB     400      a09�7�,��6���ާg�;�¢6�)��tR\Fɯ��و�ښ��w�����������0
�K�s�+���D��<��̶�X��X��'*-���^yX���P>!B�L�d`�p-�1� �H�g�~�Lb�ɕ)s-/+SA�������;�I�n��s�u8asXlxVHYEB     400      e0��X	��)� F\4Ǎ���E���!�I!��+H�מ�)y*�T�H=P��h�z(g;XX�݀�=��<*�jCKZ�1�KZ�J��[�E=n=%�N��W e�֖���\�(_(r/b˙�+�~� ��E��(��"	x���g�ِ�D�ݚv���ƥ�y���6(H�f�R��N?���Io�6��[�J��@�j�\�z�u�����[�$Ê~������/�mXlxVHYEB     400     1a00I*��L3������y�#�I��pٜyjep>��x~zYk!�U{�`OT-n�K(c�y�ʓ�0iC��U��hcm1��
Ԁ������׶Κ��3�b
��"�h{�vG�j�D����	r�5�,���w�Tr�4b�hŏ�[gJ�A�l$����b���9-yʹ�G'8�Tm�������%u���Mh8� j���V����몡 ;��ˍћR�T{sgJ)��vnR�`���خM�Ʀ�Bv�~Ij�T0���M����'��
WȉZk�z���i~Mi:�{��1��>��]�d-��:�h��	�=m ���Bղ��s]���� �._����!����r�z�u�����(�V�֍�z�v�}�����7���
'�p_4���aVw�=`�
�;;��ӷf#��C���XlxVHYEB     400     150��Ql�":-�R<��z(F�n�t�?܂%����t��sn����q��b1,���Ԣ��= �� Z�`�7rFZ7̅mA�8����dG��@��3Ğ~�.��Ml3�qn�0��\I��LzǦ\	�J�ږ3����
xl����
vE���pg��D��-೑tT�zV��&�~�m=?����яR�����S<�!�[���DP2r���hJ�!�ia�Y!i�(L^��ڐK>U��\�d�P.+���3�u���a���:o�ds|�>�2Q_���X�?�k/��"ǽ� ���?�}�*r��!�؈�[�S�y�H��ӈ|�=XlxVHYEB     400     120�6��>m}ӣE׫�����-b���6}E���0|R� �E��H	�D�,�v���|	�d�$!�2+�����Վ�?͑�[d�H!��ظe3%?�P�"=,ȣY���/�T-�?� A�7�߂U�9Ŋ@�K�2Ŭ��"5��B�LF�&:)�S���q�r-?��u�+8�>8�7J�a�U�vk�:��㒌��\ϸq]�o$��ە��9����ꯢ�I"_�����x|yB���C�`Y���J�&���Q��*i4k���V#V���'���Kpr�N�<�pXlxVHYEB     400     1d0�k!��΁�ޛ�I���ջ��0��y�!� Q�NUW�)�&#5+?U�I�J]%����Д4Ǣ��n��2�,�2�oC��S�|�~כL�)�l�����~��"����4����n�$�&D��?����q5WG���۱@�0ʄQr���N�W���n��t`�V��[�R��aB�)�n�AX�fJ��B�o�̯��'�:�}�A�F���$v�c�1�9���%�$�^�)���C�誂λi�+����= ؀{��=B莤B:���؜���'�8E!��+#���t���tE��s��Xf�7������;ọ�*�<��gSC �PС�ăT\��0�\X�z�k��"fd��u��n��EF�C�=�Tw�����qc�>C��Pp�	!U%�!����B��E4؏{��7J�y��L&��t�Bɧ�rg�u��<чiP�c:�0@�Ԡ�XlxVHYEB     400     120�cq��C��a0����yWY�B���ͭ�}MV��@0���3eieU��2ڎ�玥�`�Ʒ��h�N.� R�}I<��n��VӺ�z<�{�[�2��:�KFg�D��Qq�R�n5ӱ���}�J����r�1�[��B+�	t���̣�BN�v�*70z��o��x�y>W�|]{��|7�g���v�t�+J���ᄒ���Da��H��1p	$��$����36y1�����RbĜ�QT��)�s�J_�_���Ftb^�]n�+>�]� >T�XlxVHYEB     400     100й^TxD�8)� 2����mE�V) B��9O�ju�l�P;�B]*���;DB���5Bj�J��:��wE6Dp{��L�{�(s�`��xLl��@�Ƕ���u���^5��m:R����O��~}܏�CU;��-!��[���ᦔ�W鹖Aµ���[`b�F}9��
�RAʱu�\������;웫S �(J��x]��+�Bi�� k�7�&����/��΂ɬ4kj��.��6������K���E��)XlxVHYEB     400     110)1^?0�{ֶG,r����6�~�_Z@������?�R���~�?b�8W%F�ı�HE�Ŕv;-@��hL�s���y0�K��f ݾ��#�-�gIS���`)o멙[������0\ͳҾ�U���s��lz��$5`zr�i�k6�=�A���M���ȝq���N�DcN�4e�����4��U׆�zuo���GG2�/F:9�	vl�v���$�P�G�̻�<Kt���Jt�
�%8݃�{b�&~�����bXlxVHYEB     400      d0��!��C��+�0�%z��{H��(�w�'V��Ib�_o��qN�`�M¾2�Vj�kU$`t��H�V�t��9�{�_|oi��d���m"P��'����J�T�ƚ���l�Y['�û1������5s �X�<��ٻZ��a����j�#�Es���B)��*)�Z�ķ����t�t�I�'�F�Х5�,��x�+�7]�����XlxVHYEB     400     1002��76"��Y���*)J��I�B��$�5���u�^g{�(��T-��o�1��I�[��z.��ϋx��_��=2�N���I�5E����G"=���:!��T�D3�"�i�U�L�Xy�X����hT�ǃ�y�J������?����~A�5���Tw×��@���w��\��O�����m�a�mM��u�L�����l��@����aq_Lg|*y�в��
M�"7%�/�jp`XЊĽ�˹x�XlxVHYEB     400     130R����������1̗,zy�^�H��ǟEQ+�������HdV	<��/�! f�̚���pkk%����Vu�� v��7�=I�K��WǷW��I���Ӎ�@� ��;ň?�.?���U�a�yj�&ܽhg��o�}��f��FLJS��ٶ]I2��R�V $��c�|R�f����Ř �ӯ�.��=�Wj|������-Z�1K�˨7��2�ea�m^�uwU1�����2�k���Y)���2�Ψ)��!�L������$�%��2�b��0�%��!A�K�AY �$XlxVHYEB     400     120Q'�uBN�j�)�1˲��Ӥ4K��@ʅ���k�d���ګ�ʝ��b!FIsC��5D0�c��`�zv�0|�G�e�A�f:��}�z^��Q2
�X1�X��5����=�Y�^�W�oBw������N��D�
�Æ�I���Y=]����B]Ɏs��6�>�������ْ�	�}�Ō�g� v-�8x�bdȐl�0�ٽRE���a�P�(������`�a�>6��D������νI5�+�]j&�;�I����J�DqY�D�vEb��9�\~]ٞeXlxVHYEB     400     150^*��!{��.�U���JqX�!�v��nuy�\�$�tA 5դ堐�}�Oo(.'�c��Q�тhu�Y��?��a�Rx�� �h��K�y��p�����l�G�i�ԗw@Vg��F>4����c�ό_J6@Y�	|�wm�����q[z\�y���q{����,�IwK�>[3�P�$dViJ%�}�OU�9���c�$m������'�Z�[Js(v��]��fx���7�m�.��pd��k�pkuu��7S�T�����u�� '�b.�iGc�ą�iR���X���d�a묒��f]Z����O�7��XlxVHYEB     400     110���n{Np57M��$�oY=�V]�U���V���jh�g�+C�����<on�o�$�+��?uw���
�BF5��i�@��M�w��g�!C��y�D6��[ O�-�+��N�i�Xx���5C��}Y����h,(�&�ð�ֿqo~��9�V���N:���
����mzd���A~�YI´˨���*j�R�3�=��;v�
%��P^�мfI��^��ײʴ��2�y_�G���E��L=��F��U�+����
!��1��w�(����k3XlxVHYEB     400     110��D�Ek��w߸��d�X�n�!mV�fhy��
_cGY�u��p��ѩ����7+f�?s��m��%a���@��4�u�-��.�W�h��F����u���b;��O=V2��l��N�l]��;v�*���N)���ב���`���3��Pl'���:^w��*��uP�yf�� ���t��g��UJ���w�B%j/l���X��j�4rT�6��q-����<2'��$�S�%�&��h�=�Л��b�Q!���J}����VʀXlxVHYEB     400     120���Y���ջo��jq���%-����8�T��� �r���A*���'�ag,��:$�E���|�]��ɮ�A�R��!�9���N�<��#�u*t��|c�����KU/ƙz?�Ϩ�"��7%�y
,KWK֟h�wDM5SI%ޒ_�taJ2��(lo���kf'¢$Q���5
�����v����AO]#��>�k��Z�ұ���^\�݇	�K���U���R���FV�-y����wc�u��I�Z��$[�*�B���/����O�u+�׿~�����n]�i<XlxVHYEB     400     100A9F���Ce}���rUc�Ң�^O8��KO}�)3Z�S���M��Q:V�k5�oF(R�Ai���Z32�Nz���$l�.�����!� �qq��:U�?���!�9V�hSR�����J�V��$hz���6�7�s�=q�GJ5�9��Z#�>���Ś�E�
8�/����&O�=Vgz
���@f(��4^���sҩ�	T���%ȲcK�d�6��u�8�U(O��<�O���'	&Fڛ��7�Hu�XlxVHYEB     400      f0�E�E�|��r�>��Ðc"ҁ����*P󧏖I�A�/If��3��9�o����㱴{,��¹	�Bl��]|�=�\�+�r��*sH[D�=P��Gc�lڑe5��Հ�#>�Te���	"Kcc`�`����@����s��Ka��� '�
X��꼇�^����}hZaMXr�_���Chp�Ē޿F�o�5i$� 1aɵ~Y��*y3i⽬Y���ع�\�6��=�G
%x9:�MR��wXlxVHYEB     400     120&,�2
��,��?oR~u�/-
�������9K5"]<���_sJk_gO:Ğ�y#�� @��OOқ��W�$�u:XV����O�L�'��%�q=�&���>e�V�8m�*Λ��u �D�i�g@��b�T	�+���^Xi׮�52�n�`��2HBl�5@�U��
 �#��B>���%��ߙ�l��8��S�����9���e�4���$)�P�f�E����_����U��g�R��`�߀.�t
���ʳ�GLe�Dm-�iM��	q��¹��n`r��,� �g%�vtXlxVHYEB     400     110I�1�٣J3�� ��= ��ނ�b9�;��1��.�����':����1b�׮De^�R�r��C��*�*�C�ȁ6�k�nۃ%g� Ks�rC�� �6�S��ѷ�!:�J"zg�dt���`���%��-!QJgm����c���<�F!LS����F�����h�;��*I��K� MReW({�ݴn��?諭�������ѥ�� ȱ���͟��I�d叜��i�ui��!Oն=S�-�W�XlxVHYEB     400     120�hJɞ��J�Ӄ	��|�c$��橦~�+���Ea\T�@I@i���-U���3FB���!v������h`wk�����=�5���z"�ݒ����c9�)�#C�.��{����%��m���{7R-3(Ш�}�bW�J��^�8~��M�#�(c:������U���B�������*�y���cK6��#���_��r�@<�/����n��.�r~�%�&U�A )�ef��a�}�g=��k7 �kMe�쮱�"{�d)b�[��l��$�g�@������XlxVHYEB     400     140=��uEW��KN�`���K��U
���s��F�UΪx��q��P�Ai,��^�r�mK�s��Q�^���Kݬ�,P��'�}�'{�?��M�P�"0e�Z��ȉy�>�m��4\r��v9k_Ő���Cܦూ<����JQ�|�gz�s��@�	���"dQT�ӫ�$�*���ܽ]�#=Vd�E��V�ke~�$�[�ֆ�`��jN"�ax��TCA�`X�l�D���1�%�Psg��N��ͳ�}��*��/9�`�V�\�!�*��t�ӝ���=T��6^o:����w�=��eD�XlxVHYEB     400     140}��
�������1?V[�Ȗ���G�bu�1�ZjTK�Eŭ��E"�s)F�𷨸N����]K�i$��I�J :R&���\Z�S����(yI,a͸(�ɾ�i����֟p>~����W�[{V����kd��VS�
R��cQv������N��i���Q{�e��B�L�5k)���)������i�98_䰟�Y�ܹ�D8�Mt2w�9�XD�RT<�;�*I��q��z�	��kk�J�Yn|��w����v��q��SMr؎�����K���z��R�v<�`�����S ���(���qJ�$��,���7�XlxVHYEB     400      e0�5#�Ǎ�ڹzC�4'\���N���IjT( 2@r���Y+qMqː���]���d@�����X�L���а�|#G����A���,{�׈Է ��Lh|�T%����k�p����\K������
+�#����G:.\���k�b��<��Z�5��DaI��B~5�k���Ӄg�?���yL���,k��*.t�_T=����5�~�<�A"�
W&UXlxVHYEB     400     140n�yZ���d=��P�Lj&��?gf��آq�����4y 0��tQB[W��r$/�E�e;B�o��Ɣ���XX��/�A�C1A�ő�v_�Ʋi�IH&������&}��X����o��<ǹ�H��N_��o$�8lɢ~c�U��<��U�`����?�cȖr��M�:74�GW�Y��Ll�f�o�ⷜ�"� h����5'�W�>�[;kj��Gb�o=�J)E�3-�*|LR�ec���^S�r���\�_`Gɔ��2��7�5<L�+b|�P	�Ѓ0�MKذ1���G루m�g_�٪i�g�$��^G�XlxVHYEB     400      e0�DW�wJZr ����x��И o6N2[��(��r��&�]��*S��˼��훰�ÿh^χ�+�E�͠���$���cU��`��9�k��%Ϝ��@�(m�j,R��c�!��XlS���.�*Jt$�+�Wl�(՗3���뾋�`����Fԏ��H��;�%�fr��������σOTӃY��ĕӁ�p3��B���y�÷�&���&�ؽ��`;=��XlxVHYEB     400     190/�S��a�>g�=��*�-�~�H_j�ע�y����	j��=��.c�z�ﲝ:���|�[F?@_��Nuk�)Ȉ�j��H���"���gx�,v�Z�`m�V?��Kf}C�Ҿ1'AO¨�6���(p�^��-���Gj��0�?D��8��$$�d�8�Ay�γ�����>?�<2��k����R5�U�!T�[[�MP$h�bPƿ��aR�)�4w1UnY���k�������_V�O?���3Ѩ]�~���磶���'i���	��c��ذ�?�?�������yX���`�}�c�~A+�N��Jo$����;���L)�ʈ�vʒ�S�b��[«jߵr��?n9��BAx)X��L����W���m rl&�}~i�_b4�ɤXlxVHYEB     400      f0�A�Ǣ ���:L]x>��x~W-)@҇G�<tq0�5�R8M��\�����8��\��^:�2:p�ܾd��9J*Y�r ��\Y�$��#ѱ����Ю��ٓVU�V����弟.�x���Op�Zn�Gw�N
+�^��\�*�S=��7K�h�®�����X���{0�t@�z�/�X��4-�g���Pg���Pp̔Y.��VV��k-y�؉ �0��XlxVHYEB     400     120@�B�iE�7�t��$��f����:�g �Ap�̽ZU��Ps1y�Ńp�6�Q��Y��-0��w��ll�Z��(웬W%剐H]�&T��Oz��"���^�[�k*�o�;,):T.�fǑ����ӛ�y�Ɨ���oj�h�х���/�P�T�?[ҳ3�%?I�שEzt��C�V����a�"�F�HxUڞQCB�ʸ�b�L�24���S)M�5D�������\CWgca��d<S�ٍ5]�����0�!�@w���kY�4S�.�@�O��XlxVHYEB     400      d0��3i\��'�p���yY
�%Mܕ�7��_Ў���?���.R�l�^R��lE뽌��U��Mn��O1��)�KTC���z�L���x�kg-W/�B.���Z� �K�p��M���W�!�+�~z(�W7ڦ�
��juN�\�~�S� U�	�I��#k���ja��B�8r[^e@�Xa���y�WA)�3#����|7!%��4�z�ŋ�XlxVHYEB     400     150ڿ�[]Y8x��=R�+eZ��O�\�!5M*�<�:��]�줷��97汷�U$%r��ӕ��*+dҐ2m��^��5-�Z��zѣ�������uB	�ς�gZo��}�YT&��SbR���@�벱j�4���7�`�������ӫ,�!0�vs��gF����zx�~��e����PW�7��)a��,z��l9��Y;��P�� �'*���8f���Lp�G8V]�TȘY��eT%��mA��/�Ygr��C�m�Dʓ��w,�1%"5��3���K�X_E��8˂ٶ��c�Sk�N<� ��Wu�����{����^8/ ���z���wHM��XlxVHYEB     400     180;�!#33<=��2 l��D,����g��K˒������~���4v,����5�šh��é�{PU���0��	�{�RLup�����e���v���Z��z�P�ԂI�Ȟ��w�������iA6��l��Z�)c(l� ���g&W)�����!��5l�V7(�2G�[�K������2�S��ΡRX���$�$0���1��kӮ������/iw���������u�� D��2/��5�����o��܉��r�m~���!�=�7
�:E����7�<�B�,L���l��A�S�5 ���1�]�����LU"7��H�Y�^��|��̗�ޅx��SLR_-5�񏥭x�eN��XlxVHYEB     400     120���P����\9�e�Bک�����}�����[��?�Pcҧ=�Λ��v]��Y��d��{#���!1.�خk���7$���F��I��]����h��H��F��Z����%��<x.�r�v^
���4�`9L9�����,�|i��=�2l�f6Fn�nxL&�g�$��pv#��GZ������<�.D,P���x;݈�h��t���9jQ�e�����` b��_[S��I��닩7�.��!�Γ��o�2Ei^�{-���j�t�s�kK]a��XlxVHYEB     400     180v��7q���tF�쐠��S��쾵�A��F���Vtq���W{��"E��M� ���	���OZ)q��|���Y��#������g��c&<��/�<r��/�J���(p\-���a|~I�`��R�L����:4O���L�	-�Uˁs3d��0"h#�k�܉I�2���.S2�煽0�v�?��}��Moq��0Ԃ�%)[vN��ě��a�A��W��^N�S!�җ/1��+t-�JD�?F�|*/�Yɮ�[�Ҷ�Ķ���iG_�d���s��?4a�=��+z���@tzΫ�_!�	�V+	�+��.,�,�$(�L��9�vT!�ę!)2ï&q��o5��p?p�E\�h�a�0D����_y�ôT�7��XlxVHYEB     400     120����P��HE��K� ����v�J.�Î�97U��
F�a�π�~:D�TR�Vd+;W)X\�rJ�U��R��o���۫�
x��%ьK$���a�(G������dMը�/���'	�G��co
x�)�ß}0U;7��{���	�V�^V���pc{@��U�#�*riT�ϯ�Ţ�m��JǱ�ݐd	&M�m2�w��
S�1tv^�G�:�}����%��w�2�i�&(G׆)s����*�~e2h�jD��v�{V�'q�c!~J�4���n��@XlxVHYEB     400      f0~�`hp��.E�Ц/e�N_�I^�o�f�ӷ	�t��Ol"�`���s��1�t�����O �҃f`��r�̱="A�^��ȳ��e_`<l
��0��(�ϩ��"__���sL�� �+D��2��?Wc!����I)m6½��ey�1\�XMۿL�rסA0Nj}�Yd)dm�9��r�%�̍l)쇚<�*�f��[0߃*�R�;��bo���mCÙq#*W'�$��(XXlxVHYEB     400     130b~�Wom�a0��!�	���L��e�_��,iH7��_�X�\�d�E��3��o�WT��M��
��~�PY����8Y�o����o�	�c"��N���40K�d]��D}��E�NF�07�k��$�Sl!j�:�Ĭc_t���������Ѝ�͵�����{�P�Z�-T�E�X/+l�F���dVϔ�u�{�����h�;	7����s:����bH�E�����㌿��ՠ�<�[��+8�suX�N����kG���k_O�d�C�fƸ-��bG������@�͙�ʹ��ˉuJ�@2� �2,(XlxVHYEB     400     140f�����lL�x���Ն 1�T��6_�)G{��n�w�$�+�����N��U����m����˾����[ݶ`�|��&��w<�A2[��Y N_��+Upn��lյ�?�=��nf��F@k��"���s.'���|�+�E��Ҟ��`Xğ?[��M�+{h%����acôRR]�&2@�-jTs��y��j6��g�&�� �z��2+h��2�3xF?�O��3��[҇[O�:i�c�Sav����y�����Dx�b̝; Q�$�ǒ���D�T���h=��(Ypp���r�$z�k��m�=*�S�nm���XlxVHYEB     400     140�<h<��D����@�F��F(�@v�7�MۃM�����t(1��}������b��
ڗ�I\�G׹xB4;"D�,���� �)��h���6x�ܳ[����ŗR��,l�����ؾG0�d#�"��$�5{�������+����U[�EP�y������$�����CO���z�Ҳ��Ǯ��� t�=Neܠ�x���T2	����uM�,�9)Ib�ő"q:�Z���+.O��C�}ቮ����qE�֩Cw9�ɞK"���t4c�[wߔ�B�w�8��G���[�(�nB2ɳ�h ~ܶ�L|�YF�XlxVHYEB     400      f0Q^\���BBD�5m��;i��Z��}�ք��Lm[���N�E� �sJ�ʲ�Ӱ3��1�<i)9�kɀHc��x����/ �Ǹ�]bй'仈Bu�4@������D�����jm�kz�w�$Τ{(b� n ��9j >����*��S�m{�l ;ऎ�kr��\�������ۿ78'� ��!�-����N=������?|g�4~ φ�����!
��<g��/��S��_DLXlxVHYEB     400     140)�o�z�+bI�u����{[~=�]Ue�W ���o�d?�e� 2bi�>���j0��̀�k)�d:��)�2��в�x�Ʋ���PM���������o���8��>�>�Ÿ��I/�tL
(�kB�Y�f����@��_8#�H-+����ꎠ�W'��I���.N���W%uc���[�#p��|��L�Pςb��׭tF8�'�پ��o�3/��H
�AzS¢��|%��v���	PH$������VP�����t����U��΁�c�$3����o���K�<n����젼���"���@�'�B)�XlxVHYEB     400     120qM}b��"��6b?:$c�&�|�]�j�
´�9�v�o|�$yc�/҇ Z�BcL\��b2[�ݔkT- 2z'"��I�XP�4e��k�M̓ؑ�zw��,���;!Cp�yLZ���X�A}e�?0êu��1��l1��W^����Q�N[s^1 YMi�����|n�$�g5�[��h������,������ae_��,4w���g���z�w��:����Tk��~�����Z�̼�G��'�\� �>H8d�2��7l�r�ޟw��\�yaXlxVHYEB     400     120*����q�\�1��q_�9�������?�2j���}��Gh���#�hV~;A����E;�]2�����n��"�}}�
V�k�T�i/_���� r���LE�i��j�A�����Y��<�l�@Ǿ�A\�����:&�/U�sl���j�e1��'uGX.cIDE��q�s�Z���T�y**�R��iWWp��M��9������<g��HR)DU�0*���,ʹQZ���fqٯ���`*@�}�q)�h����\ɴz�ϳ��n��
H�n�pܖ`���c�<XlxVHYEB     400     110&��q�����LfӭR���W��U�wG3���Q�{#�y���m�mM���6��`�Z*�����&:a�;������P��3��'y�4![F���DM�	�]>M�Luo���&!+^{�)�?m9�+�iE���q�������Y��CZq�/3���Q1)��d>'�a���ò���okg`[\5*�I�dk
��`V�gu��o�W���h�5�s3�kږ�X<�IE�a�+Ѹ���#V4^�GIZ5�����=��_���\<UxXlxVHYEB     400     160����yX��_	ґ�^�t?kn�����|�PJ�sۄ?������:�G�&:�}]۪���{���t��T����哪�.ƒ	)�@fl@@�ٍ+ӹ>��s�L�+�U�'�%�vFSȕ��7�m��E��5,��Ī1�P~��G���u�sֲ;����b3�T<�⪼�Ё��ĥ}�G�V��2���|귃�U�s�k�v�г�I��@�.��4p�H� �R|��Qj���A��N�;�!Y�A�^LU�9��P"�7�@D^.�ʮ
�Zg��v�����
�>O�kI�?�M���w�t�O4�˔���U^_D� #��_�>�H �gUf�:>XlxVHYEB     400     130�~g���0VV�b0�]�.ܘ�DE�<�+��2�g�"��as�[�+���ϐ'V��w��GW��;�^S�v�$#��>	�M�Ǜte;�N?t��dƄ�z�[�АV�qK�>^�ͮl��N�0��}M��H��?�D�CѴ	б��r����S������3!���Z� +��"�@�)F���Wu�p�g������j��Jx)%T�(�L@�}���/*S0O63���m�g&���2_���Jn�35	J�qP���Mۋrr��j��.xfD��Z?>{6�������V�����#Q��,�BXlxVHYEB     400      c0#�b�PA��.v*�|γO8���w�>�S��a�u�l�q�N�ڬ͡j/�ꆣȃ�˃�	n ��4ovB��?�cB�d:��+��U����܀�2��R�b��F(�F^����O�e�$j�''�h@�P�r����34>w+4Y�!�|�O����c"��Uӳߎf��L��� ���3��oQ��ctXlxVHYEB     400     140;��!��3#X+嫦���DX>N0�\�y�j~(���a�	�D�jon���MK|��^1x{ �&�
�X���
κ �`�m����B�F0�2^��,������Pz���֖��ej{��g���_YƷ*%�����>��>5�{E�&�!!�a� ����O攺�C�W�/][r���SEB� ^C�@*I�jbV�.���_����b`��<�� ��Z��W�����ː,�IqtĹ�cEnW�"\��@�5L_� 8�ֈf��ܩ�b����|L�gf�����(c�
q*}9V=?T��"��� !��}�7���XlxVHYEB     338     100�>9����}t^��X}�T���; ��]p��t7:u�h��[yK^����B��Ҿ[Z��I{1!%�s�V����X)����C*|ײ���^s�L�_�E����;���Ǉ��b:<�r%;�a�4YxO�g���������"�#��E������%-`w�U��}ŐC�J�%����{��HAJ����aJp���o��\��*c��-3�e��9��+�~��q�)66p���:�v�X���(W��k�