��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���{C�%�P��%֚��	��3;�Fr_i�<a��R�����j�*T[��*�/�yr������9�8}���l��f<�EB�j���\h�Rw�F��׀V�~ْJ)��q6� O�)1��?���0�l�[�!���4�bȥ/�$���i3d8"Z�@�/�dh���6`�t�gÓ�of\�S^	�zI�����Z��$[�s
�jur���ȵ=�/�Y+�F~�$�БQ��K�1���zS�а����K�=	;)x��I~��ƺ�[w$a]V�X�o�)�%Уf�.��������\gH�u����r�u������ʝa���Ƹ�� ~1���_�A�MG���%��V��l�����9�e:ǿ��xS�dt�oh\T���|��
���}�.��$% ��%e>�ܥ���R�x�cZ�
Ye�w��K(.�X	����B�%�	�����̙��~�׀�2-s��GC
H�V��BwI:���C�AA_9K4��Y�I��˯�54Ǣ�����$.����7RYBrX�Z��\*?�������V]@ǧ|�X�V�
�s�k����0�ݎ�.�]<ʡ!�����v��xMj-�5!z5��Q�J��NO�>Xwy�%�+ �62G�P*�w#
L0mPv�5>�۬oG�F�1̸S�r�,�[*-J��m�|��h�}�ù{Zy�{�q�t���f��m`����a��%��J���N�ll=����#P�{Ԉ�U`#Cξy<?ݦ�J���	J?�n-�t�dȑ�����?6�����6�/��z6�ϡF?�;�	�j�S�X�H@�F�'�BuAP����>�����Ƿ���`}a#f�HC�5R��īc�M7�����l��|ׅn�P�k".�U�S���6A��s��9�J�'��PR+`f�ܸ�-��[�>Q��Ɉ�5��L���e�^�=K=�ɖ�e	��lZݒl�Uy�iW u�Ȣ�2Q;r�n6,<�� �Y7�@~�,��.�,4Y�Z��J�g��f���Kh��(27�����g�0�=E�_��� 
�[\b�rǧ�3O���1\gEĞ
';�,�m)��b}��O`Γ"<1(��0�!�M-�m(�����������(��y�0q$���CM_�]e����s��&�~�M���a��(�;��oWo����������%0��ɐ%�"M�o�Ys&8��O�h*�;'�@d9IK@�5��)֬|���Ћ�7+����UC�t;�3���ǽ2�d?I�)�ù�h�?+�^��O���?����e��o��i���Z�C�?p��0%k`��Ћ�^#|=z3�zֱ~ݘ�(o%'��\�VnO.԰a"�-�'̓/��B����?�U�ډ��&�d��O�������{I2���3��⣿��6��,/-��a��R��?�C� +-X�#:��G+���,T3�Xj	�_AT����:��3�}�bi��B���c\�hy�(��O̹��~}h�\*,R��m��|SG#U�f��:�23�R���N������۪�6k�*sAC4���������M�pi�7eT�O _u�\7[�Fm^=��F�9�\ֈ�s�4zl�c�O7N��i� ���	�YS]j���M�
�q��&-1��2�T�cq��4+��]�e#�P�?�@��{�I��$�B�m̫�q+:KIy��K|t� � J�Г���X<��Z�]�tn��TX����p��NU�kMt��S~g�緓�"�G	Ugϸ�`��e�ĥx��y/y�k`��vD���ܜ�3�@�������`�(������˂X$s_��"���L�����ցW�I��>w�GcoI4	�hn오hcSuu�T��'1bh\��ҷ��EQx.N,ک��{��Md���/�.�������"�y���Ex�FK� /W�m�1��t��	�kl7�Y�-�K䭍���hی;��{ q�j�~9)7�N�K`����a�'���B�L�f����@-�w�J��$�I������D�2�%����~Dv�����x�lQ�2.Ft��m'_�kZ��dD�ahBJн25hܮrj�(�31��_�o���L����S��U���6ۨsQ�t�]5d�r8��x�bJN��H:���.^-&�{*}��Q \j& <7ގ\Ǿ������a�� ��*��z!���<M�[�w��.ۣK#��S����X� �d�dJ-���/,�  m�}�WC��w�śu�SG~��C�^	���z�|_ܔ�&/N����IY���G�xn~�6Lf�������XP�+ǣ ����X�Ӝ�;Ɲ\�N��]�1����e��?�J	�9!�&��l���;�2�g
=l������'�����//�S�����!�"��:'�v�Zn'���nBv�Dg�lS �9#��H&D�w�VKb�A'� �?@�����I��1l)$⚾�b! z�2�*��^�j<'�߉��:�iar�o��iM��p��k�ł�������a�׽����ޅZ��eBJ]a�tC.��M<Uw�M�FG��)1�a�,-�*e��>�rU5u��7Zk��+�3�Qj�P$Is�j�.�����|���R�g�U .����@��lV�F���Su�y�-�8<gwc5���~iL��o�����|�3��c3��.��F�8u����b�[��w["�5�.��Y�&���=�נ-oxNL"��m�tP�G���{��#;76Jo��z�7(�pE��l�娛��c��/���+@���3�.S��f`Zǒ �