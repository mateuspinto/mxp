`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
akkyovSPXBM72Kh7p++rmP3ruHDrcgkoLLWC0wTKaTXB5M5QlCcbvw4O4IjJS+hiC6IyCFdg43Jr
5zfIih2wMNW58Gv4Lklc9suaEx3XAkKFlQA6GaR/d40QPHw5w+ap5CBEW8y5JRVZiVR6BqPqQ559
rZY/nc6KLpRp6wp8qXzeQMt43hysmMDcTIzIf7lk8HGGBE5rP/ZliubfHNn061cpUoLMd3eSK1QP
QwLRU8YK4k0XfVqfAmRWbrkaCGp7ZR6XWi8keWRfvr1/eWnohOjBwuoIUkRjjzCU5Yi9UGvONgYb
GaNq6JP7XHLgM2CI3RAmg4SVjk+EjqBGPXhvEA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="EYK8yB9gLGz4JzVI3h0cs+gBq8/4r2zdK+TzCb+iVOQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 54304)
`protect data_block
ZQLdwlpu/9OD6NSokm8uRG4uh6oPSs0DExCin3ILIw2JsTt8EI0lQQmVTZjQUJaj6xI/N4828e5F
/Le0LlK4LYh143+XfMF0l1RUz4GuPCIdU/XCzzf0ym2CFUo2RZ1cJ31fgu6izYjcA6Z35j/kV5uP
yTICUU7tKnudYzrSScP7Q84vD0c+TCgNwnmh7Vs1an9QivkXBuzHwp4uC4sZmqr2Vij29Ps8ypSc
7xGucR7a2rkJVhYbo57Hs6t6V2MEcVn5sY7/DokWZIVXip+Q0AgxmfjyZX8lle6CSHT1PQ8mKoOs
rGa5YlWWXBEon/VflLx3ALBracjCaXYudR1DfdMqhOdl0ZH1f1c2mjVLfpa2UViIMlEXu2CE1oYP
E6FTfxk/MNatqvcMirHP2axQGanfxIYG9k4JczQayYxNrZ4r2G5FyNefQL5JzzKokzjDijGpezn+
gcolOdk6b5hAT+1puhf1qS/sN9ccNnKGZ0HSbG3tTadgA90QZ43ZnNszT7ZAyu8uPDmbF30BiFFh
I7vuke5GjVBci/Yz/6vZZNKiSSYJX0whNTCqBXrinUpOvsAg7LuJOStjxMgl7Jycn0Toj7QYkcDq
HM5gZPg7aZEFOXBfxGJXYcw7kGWNfe6vmn67wJS7xdHaMKeiRP8vsL43afVLKy7DpzTbg8oBwhTh
kSdtUT6MzFin54jQYtTKHmzGNi+E/Sj3GuY029VdF/D5dFFjcgZ+qgBzwTK0os/jkSmjrmCQIaW1
vgIlCXAqAC9u7slZ4IoaY4n8vxcTBzQetY2mwkVav9LvBe2fHKv8WWFQz0oP/+0xJ/bh60lk9YhX
zGHQlW5kyxXVh2HGMEbtKXFQ8/wcy5mfG6dV1XlItXLqkva2mkhJFQPbjrC61QYJp7NSLYSI+Gvq
iWj189NRi5M222CvUWSjVq/APpH4uR94PKa77yhjJxa1kmHzBxNrjSsyi917rZ+mTrfW8bWQQ5FH
VhNYCLJiVm83bpeAm3DzI+WuyNZKB4/iJ8Dn2Dw7/4NP+8HcUyLh2FIJpjGY+15eV5sWuyH0iu4X
p1Cwt7oOAqcXbWCLjIRGV2Kbey8qyoRj8Q7i2z9ejufPVzpdoOQn3AxOTZmy6J0auyCL03nWIEUN
xiWJsT9MBJGLvSZor2Hc7iHUNu/xNOehc+xTVFWzCvroz/Z6wUTJSG0xUbrRdSzcU+iG7RYVXhOO
qVgOmaCAC+edj0sKYG+5hfAoyI+Oc3S292Cuc8ym4JdHJbmtWNqPJxRS56/TZb+ISG7i55/JQYvx
iXKoW6bEB3u6BdQA2EFcMO0hil9gpLzlwZ5kRqhRlSpSUfBlsTtos460C0InIdLuc4CvKaPt2hVl
ZwiLbtucOe8tf11gs6zxg3M4Het+Yexc0EDcPtXA6s+uXYdRJkfVuAFaDmLMnolSXTsMdLDiugdx
3zp3/P555bZ38uyEl5Ofmkjv42WBApdl/LQ/yCgDzEh4WSKLkCD42eheTRivPmY1YYtBVVjv5/QB
B8uUdLLqgnt0QsWZrztdyqvk5HI6keea5YviKQkit3Pybjrj48Z1WSrMr36yjc9TY3jqIoH3Qah0
qGO2IpSyDS1SyjoXItDffggHZP4slgJCTs5fngiTrCrQUNx1J6g3RQc90GuBZTOtUa89a3AnhPH2
rZ/u+aSAGm47ue8NRaVv3Xl+vVpYmP36+GJPVf0ZaMpXR1mK306w9oJmVwp2xn7XBWevYK2ud6U5
cRma97PVAOzXaOO0ynSO1KlAuMQe9deEacLKoWX4t3I4CWK3RXTRtpduThzPtGjsnAH2gWSba79b
yJoX668DRcNiril7S+WEHU+/rs7Htn1/nHgdRGiano4bZnHkrF5KyxJpjUhjaTXJBeIpCHj8Affl
7jQNbaOR1vDLS5iVZN0nPhMn1mukB95UN7gZnnvTYf7XO4Jmejko2yhaGn9Uixl+9H3jjw2ZAMed
ge8n6cyLmSDW/qiCOllrfDiGPwif48tAJA0BciwtPqWbsKqkupoRLM7nTtRVCnqiXulsVMqRELsq
cRvPNSv64OQt1lyclAzDN+iw5fBAAf3Zycw8cV3Atc9tEhWpW6RtrT/kznfLhHIzeDif/Teio+PL
k3bp18s6gTQa/zRjH2QYyYlkTuKmbA5ICLm1hkhyzpbHDpBLPQ0rPSJXmrFDZP6Ll4yovDT6IUfP
aNs6ZeDiLBqMQLNAu9ImYq+Fg5jEcEzBuFjpIL1p3YMXx1UWGkTcoYBBjqs5dIGsVfnUV/ObWVlQ
K23r064F/v2ej2IQDCX1mqmOApeqoufltHEB6TxYbz6TiyvXSxhMyKgMGAK1UjFsV9bw9kQUTQdc
jvMQ8y1WsvE5IV3gXXKqPuHCCsI/cDbK4/nQnVnQ4gPQjvYvW096CbZaTDE1ugNMH6YfVbDA9GaZ
NA+YAyvH+zx/2BhVW8KFYpQeRv1DQ4Dss5cxmQ3Up52EYb/kFaNCWpnacjmOXpDAtUbz7NC4uEaM
EZwoZLJvWJFGhC9qORqSqmD55nfaAoFmDwPfZvWiw9GGltdB/wf+gKM9dNhFsZARFPrZuywcKPm4
spowqcNTrZOOGvCnD2ff6fzAJOs7dZ3kGZF8RaDVEPg8a9ydodQSHGg0YhKlT9ujv9gABqMdbOc0
5gA5BV46WAZqWR4mpfzpVm6TxWuDT5gkbHuIs01T9kRye5Chgd7n0kJu84xu1KP1GGVZxhmjE9qE
MrzkbtXA6vEZW0xXl29jGbQFB5O0U+wDnQsVPZZiEnwpyvKwyn+CWdQXLoIzatjmgVZh55hE+PEb
uWO1FSkqHfd8ywBmcKjunOqd2xqYgsAlkUfL0FIv0Kz+cD+Duq2F4EG+sf++RpDJTcnC5Qr+3y0w
7+f/rxjzs0n1NP1FGzEOh/970zR1FHICf1caKXvgV1bkOxC4KVRNscqXVfBrWtoXfvvdign797TM
p2nW9kxiKbTi4y6bGo3dNtbeJgs5A/fnZee8Eo4qViws5MIUz68ktvrS74wnse1/dAG+/z1FO+2M
rXrQ4XjUT7FkMoAgmmfIxNsD+yNOyteOIEQ1JjVDme6uisjvPKmYYFeL/HZJM4yTTUT3E76m5Z4g
08z8tGgwhIHM6hJbYqpD0Yec9iJ3SnqDJrTaA2We2WUKUAkdoMrHxJ0rUHl+YUCji7g8ZgHqS2b1
J+s01Umw+6CxspCYPc91LOn7wZGyflXjCE48+/IqgT/p2gelO0K9xwUJms23UNtQi80Z6cSpWS42
rYGsg9qKH5IvQbkHM0OAYEEkPInrBVteMTkQj7ig9lGV0qQcV13kUrVQRlWs38XCm2SnSpFywpjK
DSvjiogR31kAu2r9bA2OQnBoTJn6k+uqGxzqqkDLVNz5le5840lSu3eOxiMn/1Xqn6bDkikZBTrn
0F2CaGRVjBVvfGTVbpyqnps/Pp82DEWBJx0lD5Uc8WpRZKUVmTgwjCBzOGHfqv2ViD0RPKazBf1d
gxkJ30jTSkHVTaeLgJQ1ChMzU93S3mQFKOakdt23hS7reDtwe8KG/Encwp1sKVd7bFS512K0L6cF
UoTfFclgKnpODQD6JR+Y15IS4nGQSF+NmxLXNmqtMKsrYEZC8oGhTiW/mE9hkeuEoTzMnZqUE4+F
96e3qYsvYpIV/xN6u0quvcl1m3b5ClYrMiz8VERXPB4iPIxSALGs273OUltef1OXouzGp9P941D2
veWhkgNC6qFKGcJ6hDAVsfkt5GsKOsGrQP72L1PWQu/H6QZRg/5Nsom61I8LQbfEv17b/oC+dj0A
vXWVC7JMGbUw7OSfC1V0ulQ4d56k3odzquuKpPn5OQ7spGbS/ILpkMqhj/gHMv9X5Mz7S3K7psbd
+g8Q+A0L7n30mOwElgKSfp8VxZDx++rjAx9iKoe9VmVAL00hZwy6vQwO/JELbA99s8V6fgQ/i97U
jk8MBMkcvsreGrl1AufLnYftVpJ4te2M/NbO+q0b16hvjdUMkB2jjuH9JVQn2b9yLtGUl/By39Rv
7oklRWkXTCfdji/npsSYAWV7pNWXHTSX0bH5Urz2V6QI4gUJD6eTn3uNPGanvTJzVYne7/HIdpi8
PIJwBFp2D7kjtG7cazR8ao53BfXX4pgWivOgArdo+ksSGf/kqS9l6kV4kDQvr2E61e0StsOqdTnu
XQF54EKWOmy/SjqNAA4tMJ/nB2bhN0wccY52r50P6GK2KNkaGJh86+PF16fNC+kO49ET5fNts/56
Y7fZWU81+SO1JQHGuYqgODQLf63DEI0V11mQDLFgl6L17Z+YkP1uMAVpsc1SmLHY7I3SibCdMv/N
6Z+BVHVyum5V+L6GpJAtAFHlVL/DzFRBRQp1HKzdeIE4CSeeKV7SWoJo99fVFa6SDpOaT4ihku/e
GJXVrZgHPJle+yhxiwSKYjUlS8G7kKvEvDj5m07ia9qqgWfLPdS8nk7yCqsEUO+ZBYhIOGyrmfOw
/wAOvbBk3Xh/K8cpmLzqbrqrOw8AUefrlGS9BBU4+8Ix4wX0C0yo061oN2leIZc/SFSg6iEWvWq7
xZnPBuq9c2uvgRW7rkAp3zDHrpbZGCRU2F9lFbVDWbUTI+qetYaieSVlk+xm2b8ngv1hsbvc6l5Y
0V9XQHkGBwSY4aPwA5jARF/XuXSpwTk+UNHh4ElpDt8gjwjnJRpQZsz2x5FyqNCLAOLz4KynPiW5
tNl28yGM6OzNEbZmdOYH/nNWkqnJz40KRq7w96vXhk8NgSdkweTu+/8mZFZAwDuXqD54bOU878nQ
scv8MHE1pFvcf7gGZAL+k6kFURLBPg3Z45iKB02p7pLnNx51mHKDcMu3YKJusElVSgUKE7nOsL5n
sAV//gGwTGU2FcWT01QHnuWjIPhifWZ7fHa98xwY88JhvB01FWBd8h4MEHHHB5CDcAJGWnVhMCrL
CM2C2F0ApnXOINqDTJUraC/9dL+FA9Qy03jHtge/iAB/OglV2gaHO7vn+1v6DVfsDgwk/9bcA5ZS
yxafX0vDrC07SGgLcLOrRenY8lbeYS6jxflhitj8OcdKNFNUin5g2mn3oYqNeZDfpusu8SAUtqr6
yEIDTsuvbcX8g34bdxp5jLNn3ObdcCh8vClxstK+Y15ptPbOo3R2YiuYIgOHbmwCHrGrzetfPofy
lWt2w0PlQYS2ubz8kcQ5VG9VPg03UfWi3PSoWCf660lznR8lLLLR3BqYITd3/jmEj6bN8HXkSUpH
08MONQDcD07EHb55tg+p60wlCE3iNGAB+q9K3URKNPNtI8jbjGiC9BpQuGHIHjxFyruJ0ieTLQAi
kDc9dVkmE/aDyn3JuXz4YQD3qgYtkY1SV2oPovDHf5EuiY+XTJPm+h7SIGlD/0a8wKSpzCG0QIkG
gUfizdOjbHqVoxte8qxXA+eZGuSvY7wOm/uHb9cCgU2dnH2U9M4LOnc/LC4uPL9WLXF8Nq+qPG2c
foo27lS4oLYGPOj4QrVk6VbXU2/Kwtvp00tLEOAj99Oiod6YL6mGseFTT/knRuhupaQmhwk4HoQM
w9n34MmfnWZyMnpejSecS5eIIh+DF7m+iIjFsp/W6bEINy8c5Rpkii/uUU08kPForb/74J27yZ4f
p5ua75rjHhmRXe0KHYeJAn54rll4bV2dDMKoIoHb8MBAOTuAjfeZYpYBqWYOsdwcbHX+oP0RCnMn
E5U4RYEJTMfxQLJpsTn3MMzTaxeWntbzSi1PEx07k0+8fwlfQPXTdfrcisUVtF3IgeXcfa9Ds4GH
J/MuGrbAW3t7+s5jXsv5hUMn6Y5obYwjtgnq/OrUclUJgap7lDJSsxkRnMvMd1bozA80UywHMo9O
DQk9qDLRfBfYQYeF4Li8tgroAQqvuO30nWmhpLFnM7fcUnp+g+3WBjBZD+t2/4fzLQNREKaSbdns
Ya9hqw/7OCGm6spPicgvQdpsEiyk7Vlg1EpVDjaWEnmPWMUZBm14wwGg/JTqoC4Xk5rRsi3abljy
QhNzvBAXDSRbURNJluuxfoNd7F4yws1yDjbX5MlhlaUukZD+haIzBZYkdDeitOiiYJMtj5sKsRiw
ZobKX3qblqmNHkex+gzJ5NQ/F5D+QaTkVfgdIhZTyJj5peorYNnGPK0jXElaNOBKS9IYeDCSag7X
N7gHXLL7z8lig3UJz9z+U4BwjaRZrmILL3pDj1Ts/Yps3EFOpReWagJCFyaOA1BnCXMOfFnZ07YD
IamBHORlqn2Pi6VwBsEU2QZfCoJIZJPa4qg3KuCxva+fD2CudwL3pYQMYjGZYN9oWKTaaKBjnpYa
dPkSZ2gd7SiH5m7ttooGR6HBe4zoooGLxOvZx4ip39N4AGFwjSsH57neDKRyozrnEiqP2kU74QaF
OwNrvpa8XqwdbxAQS/hFuD8fCwNqMt9QBXvddcqb7ZflFYaAyXH1k8JW9VRI6ojmAa1eAzOwTpHN
w97tNnwfq182Tp/LqSQ6IqxkwleL2lX/oV1HdPZ9STm5TSOV8jwyQqbc5inOV65qm0LI4VbGr1Ef
j40dAk6iYUASvgbqH+0ggNv8+aXh/nv5SL2J5BY9NjTV0b9CQZW4mFWHyNL6CguWCDwOLSu0RQJG
6k8RWOQRU9fBG51v15dUJiyQOEBQyJ4LdupUUOdnm+7UvrKe2YgxiMWLtOMEBgOI9n8LGH21/dM4
0tOszJ1H6CdzVmOxenp21zoujSnW2A4nw2G8JvnyOJ5SZKeOrSqk+MjdYcB6G3ojl1BphYSNUS2q
4PgU75f+wqJu9/QpCb9YD/X/Mb11BevqrM3zoT/6M1V+tP/6Z9NDxIaWcU68XvMhdE28KIOvUi9A
/Ic729xAE3c2A6Fk/HUUEnY349xqWkBF5GB/Li3WM0YIx6F/GIf8MA2MV4Rqk79p9Dkhmk/Gw5zF
OjRIjkCNr8uv7rejfG00zQlTjBop8BIMfsnEbuCOW+FHe2GdH76A3Y/lIeOANDAgcvcSNm88yAzB
hZRGj3M14hNNWCegQzEx8EBNOSJEiy9fnNVQfjVfP7OCTRBhmC/96/T52qDdeiaj/7gv8j0npPKp
gCvbiNOKpDdB3a0ZBvRIri4YOMakNyx0n+cgDs1Tz1tHMOjBelqGRScwX0AqjETSpy61WYpDkvB9
C2EexVXhd0qrGYUDJZLuxZhCBNI6IcpS1cuHetTMUL6ABNcgmE/5tgLUtkD5+7zO5mg6S5hWAqVO
Y8YvepF1aSJuJU5zA5IMRiFRxTS6KUpScrCCScN2fSFBJglxb8WZV03sMl5PZ0EI18HO7VYTJEwI
GNc3zcfgK9y5pfweVnzaLb7MtiL7WCo9Nalbt/TxJpS+2Y0qQSsy5HjGWqNWGjXwbdLuCCy5hGoZ
4TPckTo3+G9W8wxeX1D8o/+UcRhydyKgy8N/mwyLCwbsWOiyqmKqdEBZNlIsqFZzCIlSutqHHgtI
ZV3ou+wefWQ1mQ8j/DK9nk/tz57HNZcUBLV6iS2TdgglfRGR8JSC6hJzEowoLztvp072UYQk0OE0
qVpiCZN2j06cUbiOC7zBK7+Dfvlvyt9/agTkRMyNjF8PikNzK3T+A+NDfe0jaN+8zvsA1w8FMB1g
pO+JveGwJbSSyJkM3NFZFd6nm0J0pPkzoiE1frVD3//HuU95izUdGVRhfLmWzSLKsSc75RLyjI/h
QsxkXhoLgiVBwwLU3ecHgXxVI+fgIqhjo1pRnrsfH68eHBPg2X3mJ5ud3lQBGbptm1T+3hpyJLnu
6BjC7+nzowXFiS8tHZ6gsZsm0CxDo4zCda7b4BUzlkQxax+rYQMJytn1Z6oqyHUwAsdvAbTVJB2C
T3OWMYUKuZQbhsvz84j3mX7uddKYpk19g4qLb0aP23tMh2QRuQJAeksIRIGPesiluCjTaD2B+mlt
Ft79eml0S52r5w9a6WUotC0Le/Hh0k7OrjapMXV0yNW1/tgHyPhiMbEG448txWLQW0dlDqdgap2r
qxK6quTqY8xVS1WCl3xqR1kXUNw94BY+vEHAFF1vIpV7bwykTCoZw8xe4vukGFmnVGQ9P9oVU2L2
C6WuRTUbwUGtv6L9pJc4fzJD3adaxohBvJSXFgwekZgZW90QxuH++9gk1I1rZMZyfQQPe+vm4V1S
N/OIQsPuPURYPKmXuP08KSFZhtalomBp12YRPOzPTTcrVukTvlJEQJtV9SwSq8xe8sqkFldtzm95
7KFuRCrM7H0phPivvMSxCV9/RFGekCTobBE8tArvwxnZQ2Bt8NG1VxFD8VNmMdIjm1akX1dW/k/5
CwLYby3LNul3xLkRCHRje8DJl7AL/LhNKQf/LvPfP05KRW8s0UF4V86pOtl3E1EA7zGCoTEAfV85
uKibgicvtnMdkNXQMQZLa91fXKkzeS18vgBxMCqii0EMwHl/AwVk8+fgNDrnmO5EpWx9HwL1wiyn
uZKpdZOBTC47pKKBdB4TsuEXyp8S+LwPgD/2+SjQ3DSj3j+tDIT85OKCB1YxyAXUdCQE65uNH8Fx
pUQBj2rRQVpsyji86C/6szV2hV7Ux7DCrMXPYLZQOUElCUfp6mfcOGhfnedyph3vG7NFDSp4rnRs
aGcfUjG6zeKDpAszXfznuF30LidDV/dvbFMKC94gdyNaDMDbBgLmsaI69Zr4KzbZqjVDPZvsnSk0
uN278i9jNUSa/TxzVyps+foKSvQOfqjUHCqtf0F76J3U8THMEd/slrmIhfgwycgxKwbPD6cVjI/i
kOQl9b0CxFBgNyeJB8dEGF7CSgW68OQJVuuL5X8JgOH7DiFxyqCnT8bY/SnJaYpTNqPJs3jHrD6f
gntx2BUlutczQfmVcBAOGsE7rADsDKNVODav0YNA/IL7gwPImUt3H0MdfKVnqCYvxmmcsjI6s0BI
SwtTSaWditgT3mrCWPjzdoN8HKPHRRNhNstdUXSZA80nmYIjhkaFQsgmMxkJUCTN5R3by6isQf1l
ULlQ4M6vzdBGiUm/0JtbWMChGTRJDzMTEB6zggrYWYthVaZVFd/euHpn0CQY17XWFPGa+NEK+jDA
7gaYifTkfkZYKoMB9HAaQlyeypmHosn/NSwqSFFkw61ni8LyFmEIz/IySyNMM5p4m8RES6pj4TLU
YlRzr20+wzxuFT8uIgzuw3qnxtTvfMQrktSQHOZgfvLCwV763Fib2E/FOa5VjDsNDUt5zKznm/qH
3TibnhEamWJHLj5WMRa7sJfVQPDXRENntUWxj+JqDGdqLmvSOfjsvWaqWD2shgD6gzINyETUnKtq
XjUfVPMviyNF33K4g2WPqz0fx+v4rV8dNEwHAon4gHWvAD+/CueT6BNtUhReprtaBBTuQOeK7zV6
vMREUJ07rxNtvRBAiEv72j29u/Mpc/IGYdR31yYnMxe6XQMvfB2NDWloBSyUMgMDmkuXy2vyEBu1
FezLb9euGru8iyr47gHBZbl3kOtXBfIZY20Ao1iBbtHeRetql4Uk/72OEnqLy8vlfnjYyyE4e1Wl
4RBYPgsQiFaLM5g82OWPakOOBcipNlV9hoxVP9rKM6PXducC7vfJUrB2H9uLve7eEDiBAiAEX3Yy
r0yJi8k5gvvoQoxq096nboc6QhbKBlVAR41b0Quz9SzxBteJLwV2Q8kuEoflmWFqrGby1/YJKEnW
jcV2OnmWQxdfAiJjYV14Cm4KRzr8QOOUrJPG47bO5F9ZQTpA6bnforku9as80L3lBNYwH/hqaDPH
H2g4bz6rdC0aVkplKdcJZSKbUrZ+S9vJoLXAArquQ9zwC0EFsoaiA1IetL7/s6cm5L7T0N0exEF3
C5zJZc5jZAvx4buzfgaEY5HO6nUB2Mv4SFebp5EHT1zjnm5GI7PB8Wv3tPckBRDHcqsj07X4jPVA
s18ifzKmFzQQ6hUTBvtt/oM1lWFkTrXkO7P1cnx55UXFscQCFzD9JLiXYZSyUznbJpoQYqG4HMtr
6KIed+zd88wAm4bZp7AU5/BH9XQO7lYLhf0s81gjpp0vdYXVhWLksaGGEE7oEc1SlhFPw9TXmH9S
QrwFMpRCnP0bLi0MuPGIiDvXjd92UlAQZV8EWMGoLLSUR8KiFApLu770apKpGwQmht768z3TTcmG
GlcvhEAnQquKPpwNOhhsmtEpFe4zzSHgXmxhq1l9eGLhTIoGqVbhVXrcSMWe/w5zCZJ56Zfz8CJ2
ZMu0JwHqtLnKCoh+bb4qX4uNvXMg2leJwZ4gCWW5quJ5KA2HDlKgd19XPEjC99+nlbd6yd4TD/tq
/nmsaiNwCfhZ0oC7OIPJvlBfWflVIHvPGutttZSd6czR3oUyhVA6wtIko4FELs/852c6yyz3XYDY
QSKN0h1SeW6Y9e2DuWtN1Dbbbo4ceXBDwQm9fRvSgdJRUkWFK2v5KzjNK2PaL0eB0hbKl/OZLifF
i2VcsAQ7BmkVsJrRChjOb9039no1P4i3WYC5h4f0t2iAPMumn11SCDMkCcsZNhzcF7jXaPoup2aY
W7lYhgc5tfk4dOcZ42g6nSRRmua5TEEF+BhSSZSt2eH9lsTrmggCypLOObUFT5x5fmsXI1CWfiQT
qUF5CgYaUtyUm343krSB5Y7vbtHG3RP4c6k5KWq3m2b4HhebM8JwbuDHCLPAv952Kv+W2Yq8aP7k
P7ILo25pXnSrpvcCfoQIC5RQDJXdl+VsPDro9eKT5itFmwXhrdTuNlEM16yOM2a3gp5405XbPl4f
mRSY6lAZHxALEoexzbEy8fffVQoprwPYpsyutaViLGFzMsC96iAJyc0WotP08iagiS/+cxwNRGfG
rS0UB3V/5ifImosk+IRUDbm4ASNVGm7sc2HtS+MWlb0eG0DJd6sQSbJgUuTVAUUwbaMWXzhObmOx
EEJ0mb38b7Vs566EQjKq4/JvrW0FTY6HcxusqwDw4Yep7AsXzbkxAINSeBfwwqrJrkkv/0EYOEc5
CxjWtCgNeEXBz9r9SyXmyxxOYlVLJiy0qKhYf8Ug2TVNtrqo1hKHqWcTcp2g/wBTHEEZfUwaAxes
hIv8MlSJR+TpB9921QLhiMS30rgD7xQZfT9e/XEY2yCZk7QsMZQrQ27ffnvAyoYzg1jg7NF/P15S
2qAwZkITF2SDcisIAFNfMTojn4ZMIGWNEfA4HQZnLq1orMJUUTNUw0jBOiai8BWcGxFMyPRJ5zQx
IYqICiWwVDHJDIspx0c9ePYhYXrRwzT0GRWGhY0K0Q5vSjKdUtLjiLgkWuG7Zk9vq6rWBsnjICg4
ed/pzsZq00/2tmke3Fv7r79FOE2WcVGcjrkz119hVkm0C9dFZyXB5X3s6vfIwEzk4ZA3obH8dIO6
/TJ+zj391hwLffxQT+hD74pcK03Dn1NzNaXtSbJqc8D1se6/Z41q7VtqQvydcqwowz2Ccyj2OwdR
Ipdv49rDhUAF1230P+5flcdgSduH5d1aCnw9g/i0K0DPtmG4W4lpnV1E8EQ6edw9xsWsGOga/pPf
yboE54phwoU5KnvBtRmOZdkAgvfYS+ku+vL7+TbedGsZUcqluhT3CLx9lbMVyIVt0R7HyX1Wkwix
B/EnOP/hzUsFWeC+EqeNprpFmc0OfMX4JLqKy39w1WG7xlvtaLxHoipahOTHSwmgyYwDf38xooMj
rVnKXuUAtzqb+89EbqliA1YwsdREOqjKuAZkGSZjOginkUjNw5ygdLZUR4uvMccgskGcd5sAwwKK
1LqgfFq9Hx2AFBTZsuOCg5xrz/lKrYqAUJrQEbcBxWIDMH17T6sbXXiw6W8h2RTSeQeNie+f3AgF
eVpSaLdzumemgI4eeyt6n+K91QRa51Y6qlxWvbRhr9fmTKOIDyfD5S5LPUxPM+H55fNjpGsRoToG
wflnmaiWZMaeHydX0wfpIHyHgAKMY2wZJ64dbkzMuVBeJhMdA+HMLQtplA6Ovaannga9ixiXibAq
glp39gd6ajj2pMkqFBo4JXlKB7M57IJKs7MO/WiFm2bKLTjZd4qbnHRMgtEfUP8plM8vmrL75ML9
DCtH3iUGQV/h5+8ZWYqWY9K7Ez7d4/KknUe5hAKbFeuRIdkH8lpnn+B17jCNN0uq89ShOyzAsQ6k
PXDerzeiF0pN0/qyX13tR/fjumwaUbJkIcqfwjVkfadOx1iCFY0O83DgalKacLFI8uRQ99Oc3PPd
TaMH+s1WjmiItzuxOwJscBLvvBscw4vqhhsa8l3KZyx+2C0Pvd02ctj7D+KZiAKd7XzSFKl9VJ79
o0zJ3wFzyw1zT3cvimtQRl8bdSVZQB7ussF4ZhsKOsst2T77DUNFs9Mhs36CAD0tLumbKwPPoNle
AD/3gluL9gmQX9xnrd1oNA70cT3lZzCwejKmKghXHlSeG55BGtK6yta5xcNTWOrjv/viO4LGyhQG
FzF10DWvtXbJN8i+/yt9s5kNbq84lJf++ni9HcjKXy58lm2oyK8hMV9gqf5OyFqmp9v5E3jcGpe9
muN9i2zKy9euGyxedfrpA/qelrgBGQIAbmqknGPBzr2ntSfmSQeEHEitmFTroIUpg9F64V1BJjhL
Cfx+wZHJ9GUCdQMpaAMU5XVZFV+5RynrZkuJHCRf+AenLcrgiZ9wUEwv8jNRSE9UrAfNwnc+Rzwn
DnihAbrcVQSKxtyH0Ym3u/2Wd/52/oJU++HW32o/f6R7Sr3pZbuyqvZlt+9nFh9QwzxQVWhLcLsN
/8tvNtPw8yhc9Ol/UqZ8AlPs/5AQjJTNqWaYyvYFJF4/o9vxMaztCjzyhxlBCd1bOT7fj1PscAjB
Xm45tEoY+pAKi7ouFgTk+Hv9bLZDeewDyrw494/4uykHMOPHcLeCbXd4gRWYwfI7nNlQ7tvazwfB
2kBTT6v8PRJUgmtZ5SGCHAnNtZbjU3/x3TwLBXNH968tS2LjG2gfskiOff0iPiD9rR0wOMzpwDvq
Q4SGFT9nHyw6ZNuHue70tbaRKEkgwQUnsNPcPtRPVyjQ8BTFlC6V8vH3aMjof6d4+v+wTmGIhFAp
ExUZ13wqnkmHhbbToHZ1TGoG1OgFaob93lbHA82Qq27NqWlKoobOoPR8uAP5wvMr/07H8LDbBGvu
ob1lpDakD7v9D/gBB9NEZUkED8sUjV2zZFr85b3tRtF22H1+WUF8Co/spQX7SIavYYcHV2dnXhPj
akfUE8GajUkOAx9tn51ZHq08dV8qpbXCVvosiWtNItmCkO2BMGeRlo+KQLpBTlSeSaaPp6Em5+oc
337j533gllTdiYTf4AIepyzibJqDjBUrSBepGOzwFWoC1GIpMJ019fB9hQCdd9759edqycyd8mgv
vQ/PUDRPsda4jVSRZrDKNd7vY9Fs72oO97hwqPM1JBXJJnHx7egzYayhRfC4yizvIoTpT6zZeRgC
SE77LtWvlNjpWdBL+dU6MQytLA0rzeHeJhB5rKLkm0karjH21OoomQ3q1HzzO+URnAd4Si40JFLH
GyGKXia2KvSs++Zl0qDg3gp+UZWzo9qXH9SPeZlFO8MVxgC/8Anj7X5jtWI6muhVapNkvv1/dEcG
MKkefDecwIQLbRt1ZkXyNb1SQ6/eVHj6BhBLjVQqh7YhaWec5FU66HBPaitxLicly+yC1BpIkS/+
DVfmw4pYAwv+727QhPx0rSDFgKnxxhuRi+w6+ZTLC77OI6Fi4S6pETfJX8o4StzE1pyGb7ia+5rd
xOwa9aE6pnWmDK/jW3apjkCYXZ1fq+tRIuj17LbNrG0B7tNllirBXJ0iDsCUCwpVbZEcFLoK4DKS
wwgDhKHsPllqO943lBhqfZ1VmGVsKE6EnUwLMjC+0srXYy5YlOpjsXlMmAQbN7O7Lgp+t5/cCuNq
u4HN5z73WMHyDnwKUPQKFGTSqtKMbKby2GnSrczHKRxkvcnHb6ixhOOdD32av+seCoo3RBbHQave
r3bvJF4UShG6Cp/DeLTDSGvJI8AkP5CljDJc1sjhYON9G1OS6AWlvMNf/a2mUXj06sSfQ5owgAyR
GbTzwboNaEZw4K+QeQ0TDj/8rAuJcvUS5kNzGcJV4MNGOHZ1FX3ldY+kEQQVtHwV9QYpoEkiexzw
8FmhTEN3oxR1ei9gUUlEpR06KcN+JZ7S6zEgqY7Se4c9adUF970/PUh+vfQHeKiT6nv8pDuhN+ai
hqirIQrTxwAeI2QmHFdBIykPWxwuZeahtRbMsj/i6pLkzlZQzw+bH38KYCf4YuKs/mGBNLYWvvLE
TkKJPC2kuNHLPkmGIBsrPKqgHublZ92Su1HQizGr1i5omoJTyDORE5KoYcpZ6ICY8/PPS9CEE/sy
PuAUkPHT/TnJvxORBrcOBKB8G02dQ+s772TFR+BsV+zWlZZ/kOo2KOt+llHMGF4Xq/yshsQpHoJE
naF2EzXi1TChJUTSw7GMFoy0J+Otabp5RaIO6MvHR9Ji2HmYOK07Uu1bjj0cPXvBVZqm/4Bd069T
JCRKhox+j2rU8ZwLTTqs31353+jvphQDB3VR711ui4RJRCeyQAOgEtd7uRwzDC0GqzM+hTvZS8AG
DrAR4+2nwppz7kPgGgx5mDU538Fqn4DipP4VwljRe5WePZR/WXrElUzJ55TldJn1OBk4AWUWFOIb
V2dtfoX4DnMwDoaiYeiDYDGt9B4gGwNh3yYOzRPRdgs/+EvW4qnxYsHkZXeRD7EljSPwj+BhWmID
qbxwL08QwG7loTAXfn5RTa76CShyICklLhunb+E6GBvvrT3wBlwLXSJH7wX4dCzs5gKLgGJ6UyVJ
LTtNotxz8SEZEDc2bppQhrx8SH3q9dfLEdJ8p2QK+W7SAL6wspcTc/3BQMeh7gYpvbOM0mvChAWG
yYuTizgr+Uy5GsOHQTstJICuaa2jUAjhx3bvBPLFTvowiFU5j0NcXGISeZI2bAmMZVKalXKqIlz+
dGTrVF5NK6s0vKmjSUweeQBDtWnrXhFOUTJ9VbPg7ZF9V7qboCwqxyfsy8CpNRBaV7dIKCCBKEnV
mAi0TkmtcoH6FrZpG4lKGIGca4nT9vGEjLx/uFYleqzarAhxooVGCgfWtR6ZnexbT/vje56szdl0
zum7zip8/x/NIaJ+c99S9KVhCq8PzMHLrKmJU1XCGVa4TMBq6wiPpBCUSLtid/yv+qa0+4HYW4Ml
lqFcs3MroYtMPsbSadZKzXrDaOt/CCKAJ8pu4LmgBPiGKFICVlsOmhL+iTHQG4NDtIygwYhEHUMF
mvalEOz7XJWUU8dNWJu6BuywRfOWfLTQUTPABEUsFhoQTsa2Rp6KO1pnFBzmqfXW4pNUPq/OVkUp
SgJ99oWAU13pWiKznq0uogeM4MGkJ+H8I8ZhXgCpuN9mMvcdt79dES3hoUeP1bQJIU8xqZUnrUCM
ZsPFkydhx0dNbf0yy5fbgCM3tiPVOGNCOYtxh3rwxSQlaQ5ESlvGO8yY/FdvwNv+CaQTeDIK4rJk
ZJbseRQJRFNzgu8gWVwhcTg4sTD1Qh9uYQL27PQ7stwAFXBE6M2jmQ80oWzStu/cFoJJ95U/QW26
DWmaMZBqJs5G24bub5LmJLvdgeCen4+R+2/1qMfWXox6Sfw2csa+3MgKOm55iWYksQMZgPcUY0FI
5eo62bWHd5z6h7zap8iQYLxG9XgMIj94KyZYzaI45TSy9pVlFIw4VU4tH4Nn7icBMVo+4chAPRbu
FfXNsEFChupNoy2li1ystmFKehzrO10PNwnNfJeGlHB5T62rgqQS6A5CuzuLwCdxBrx5b3BP4bY8
trSlewqYNuhao7v4qcvZBtWKEVRHfMY9ZeUwDUWs3VQz/Z4aYHhjXj7NLlRka1knIQeB8sRvHb19
8joEYyxBs2GWVa3+uJfR+DY+tBie0NLddUZKbNVv4LnqhZHTC6bMfbKD3z5NlC/9/tnpq1GkOt6v
ugHr1uaqRo9C8hJONOdIxAgM/u5KMZ7ZBJbL4/bgRoXlFr0R31ih9TJU2hG2pol4OntdBFM0K7cf
zuCPIBaybfM82TCSi2VpjE1T3d+GLrKJsjz1LYFi1psKzPOSKZjBvXrHD6oze468Om3SX6+5Gs+M
Nc8p3JvrL0I6gfElfLd2Ftkgt3VqxDjWkeg8hVN5OCw5PNZ1SEU9ZcA/gTe8tljk4CNTQ3zhQS2o
Ox116St36U8fIt41AJBnsSrY3/ICZsKK0UTGx/JD7NMVZRLkxRx94v+H6s30FIOtlP2hbeJMP8PX
TlvWP4IyKTXLaocYr1/tbD3+/2BabjTswlkk6N5ZunIgEf/M9c48JFcl9RrJdOo3XtzRDjcNV5ZI
N+3gkwehcsapqmJmI8OujR/FiaMRO/SHHHlsQJ8bv5V++SCIhmiodL+y0c6mnZauU9pCUFGQhYLi
jm/ZqFTcdy+PAL7XDzKXwjiKE0ahqTosus7FXD8gpg1LOc/jZKbY8udgjCs3i0j8BQ+L5+cTatgP
NA2Be2m2Z78AAdnYmwb6l6ZTBfiS/hlL+z/PKnwxJgbVzNExatYzbS0gpFKAD4mbzaZVKsjCmI3j
zemnqoTQ6H+UoiOn5G3djWMt6m1U4O1HrbrinLQnMgpGewtfvAZUqkqMMB5EshAIAFqnNb+nRsiE
fSCRTcb61WHdp9ShH/65ggQly2jsqyY/DCn58QieHbiJZWM+kcy002ad2yDTRRfALsvn69R/+6Aa
NboWYvSm9RwKVpuzXYb+3PKGaT0q68Vj0+s/F1cM3gJWTFEFpbkfaJJv2eHqoKuT6COu8Nhs+Ykg
IYYalmoZGYIQa0G5cd0oCERRJhQ4AVy8dBKYEsNh6/rPTDvYhFqD/stXgzCWvIBSRZZZHIHFDHnQ
NcKt57S/waU0wMpOBgvaFS550gBZP2WNm5Tt9QHy34ArjEt6MZPeKcqk67j7H+JmZeC9KhUvzekr
AVSNfClFVnFvoJYmhtzQcB64ho1P4+67SoANodqECkQeZvfxwIJ41VLP8BzTnVHZOVeFa5IE+6CK
oUzSqzcYkG8Wqp7rINguHtFaeQgaAMq+DGdJdS2Y1s1lolr1afPXozt9iPmk36PSVi00d+1zs15B
tND11VXKqFPBFKRF74Io3oqM4jSMEYF5rqye2MfgJppmq9hrZITr5Tr/f5dvfbPBIda1li63YeqU
e7/NFaHcYqrWFtawB+Bm4YRrNpbAP5rNv1Ecft9OX0pfwCHn3v6w1nAqrLLMdznV90KDgjYDIh1c
GKE/+ToLwbZ3iOB+GKKoBPsPjP5y32XqS2j4P7zKZqM9BHaTxY78Q+27NJG/KaFSCf5G5Z0mnWrB
YC/uZtn9cLCSuzMTV1u5NdmPuLFp/HG5RskM2y0ug9HnrtrbzmYmrnPU3rCKF3tqdmkUcG9KA6RU
zHT7/O6kt+UuVjnfSBXkxgscpczFiNJ/uVWN9AIgZ5pM2ez1FB6qpOEI+luMQHvVIWXm45JQFwt8
02o0LLy7FetkE5n1pewn2GSqcdbq4XZL+vgD7WU37t7LHkWycr40S675f2Q74EKD8fDDFRTytRWC
rQXRxEfjcpE1Qw9WdN/Jv7DMGPY7AC2zFurA7WHln0h2GN1UDil/uy6jhciBoPFwNAs2Olcophy9
B6wPRlWuPwYbujm/FwCErCUcvB4y51iToLWZGRKXpSQn6kGaeSPY8jJy2p+0OgZU+Y+djRdHKAPH
KP18XxsqTDqksdL7QtyG8jAIRehRNrqHeMAFC/UlYfvtezFnRof3kNGtEBYWSIUjIvcvu3CxRPZ/
Zc9HCI6hQLZEMYQKJk0U4unuBmqqDRE5sYUU7Tx0qn+ajT3b03oLm4q3N5+eOAfWJQiYQ/BlMdEc
l2o5Uc/lOVKuMLw3T2PmEJFa2EhAdhOIgqCZjwYrQbQtx7z/UJ2kvJA1HUlQhrdDXfrIsO/j0nsa
Xz3Eje8cFjrhpnba7fQZbAh3sUPzhNRvQsfjhPLH8lTe3UpIgrzigwGcxfXjeVNfB4k+Jwk2adOP
IpOF41+LunvrGPdGay1qgTtlJ3FiH1zYHniUgb0hCcXyTw14HZbZhxIlwjMxQObXsNnvZPuKrVe8
YKVVcjckj5xjxl3fhg2mmNoS3kkwIvra7nB8hyfhk0mMQfVn8ohiRUR6zBEPxPXflDRJM0ZpnSRt
EZbuvDIRE5iBoNclmt95kONFfhjBkT58Ji/8L9ittEWROl58cerPKcV8RNk5AICKdzxnskfeg5vA
JQX2jKKbl0ItP+bxOvyXXHGmBc71Gt4jsaFYwJVHAL95b/Nckq+xkjh2lHDSMbcVzULSAWanjgTt
CHuHKEbNKJ8fc9x2/Cpep6l9GXEFdTBCA559fhLNRa2EzI/DeDg/bpAaKjXzJPHdVdh+TkANGtGT
c+VDD/upa2Cja6cTtoV7YlVhcGeVI8BkC31bD0p90Hk1p+CCo362S8QnmKj2prnMPnivOM4U//ga
GK8D40GvJNYEFdt6BPX4fR7qCBlPYVJ8C4YnleV3T3fq4c+StMnohaKwbcvPdS82Zs6pOn1ez1KQ
3pnEGUuJNnkOQK4ZLv8Cv1RGmqmt9yH19//ODWkpxm8nZOaEnQ9GQd9nKrLIiPZAnezbBaNpK6Ug
8DC5S0MfeJk/zVzQ10uNaZ3MCGIEqxVKa5hQm7kS6ZfBq7HGKN2gQcU9e32DCsYP11CgQl8WPXFV
RIr8h8wEFilZ+24sVK0//mH2l2h+OrtfnP0F56pDRd62czPjuNv15MALAhCzfubxTetadLs1qAmC
xTVFGLmCBUHUJmfRHEDH+YmDdBU6zAZKObaLKHIZ+LCVHF0yIpNuBg6IDOoXOsElBq1j84S/UgQm
B+37zAE1RVOCavxN4X65vU/QINMrSk730ZlBwD2/10w4am7urZ/lj7aRqpVqHVuABSUgLXRQkFnH
VbJoXxPBJfs5r8Nn//eIavNas9/lbOFi/K3IMLsctGrlu5xlUHVfDudLE7QKAb90hJ6sNfmCBAZ1
HIhD9qh6haaVJ492c1xoNJ832Np0BKg7e1gNBsR/czhVRGlFLN6lsvBEiVYVF5xdSKBg13S5TF4c
GEqPN0730YM3tcWR3jr6i7Agf7ZSH/nukWVPbmkxAldAuSoHHRElDAlZGz14DTU87WRGs+rFejXT
HtVIt7dLNJPtK1NOaXmta/e2YVAwfJSm6slxlxDfXEBEgPTtt8LAXjStlCjWdaG3A3gIbl01FZhI
oxpqBh9kLyj8Q6FfXjTx4iVmNiHu7e7iYE/jMcXeeBEaGPj5yGx8/eThAfjoUg737caa5FYy9FrI
MPrOw5fa21vHLlM3UZU4h/7g1a68O43Zw5VMjaOLA9FX2oPv54A9pqc/jd4DxuMJqpj7+lKoZeVZ
fRT9rMNxRU2iVEs8Q2nZkBeNiSZ4bsoJjeizbXuz5HH0LjZmDVqHyckI00O7m7DxQ8HCUf0d9eq5
7cMzLH2DcWyfg52rfsvFwW3SJX0iiyhkCmjU4ttSIETAhHtmkW3wlLNGD++zck/CXORUGrBoYF0K
ONbMx+raAE1YFewy7yn6SjngpMjMwOT0wRjAPFoRfDdBnjPiRpwZ/AqMgKMLrOK4qlrhLUc9rE2U
887wT+6d0RcksXqAcPSdJnDeothGy099T0JrIBJTc+sa7bsoqOuCGkiPEJM/RZyNsaEommZ1ZXY3
P8S/RCWetLpj7W8MZkhtFb1id1z78nWy+nR+uflIWlEBLttRlOsBqntj3cvpbRTKSO1F8IdKIqH8
JWuiXjDZO6GJe+qB+QVI01xSj+7EIRIoeTmCkaGJS6UkoPXPDMU4+Ti/GTbfcRWI/3/ltx9wFEi7
O0+FIxqACyKIpynqHgUCYb4wVlBFFyKylFcrzAIz27ejiXaUm6NlkA2wDR2XbDDdK+2vYJ5U7AwP
1ksNGmus1bgw7tJ3RJJqWwd2kjI44Lwncf1LZt9qfBAjoOegJZa6vP/hGefWA4I1we+SkhVDjauv
z+8qEoqHRtB9pHnIpjY5ZHNMsNbtnIbqBVgk3pJ5YQ9nVnk3jCfYHSsdEQIvw1cyjrPNFDgUScHt
Mz1hr+yBkPqqSNdUUSGiNdip8okPw2+iojp20l/4Qw/9OvreFhkKqoOHPkbFB7qIgsLu0MRQ8k7V
BuZtoBm8rL5Ej8Cq68HWdv3KiBw+SluWQh9TTVyFEUe0Coa/odX2QRmecBe9z79DK+b9GY9llche
DVUPbGHeJMRqbQopKY+NJRjIUqTAPkNfu9A2Te5wU378NgxekTkEC/jtNO9ulsfzS/YmZc0nci3A
uI4fm11wUrwriCasEprSYyJUS7lXrvNltN36EHuXmi8sAUdjb/swU3a5RI8w7XhCZz50DhjzH2eA
wEopS7zeLmGzisBoOnNw6kX/gq04E4h9dpWj/P/s8l1w13Upb/zHR+4XP01iKkZGjAjcfDLbq5LV
nKZFnES1RVQTl2He07GPIdNootF5BvArw/VpPAVnnnV45ja5p3qZafhvOUCMCOTDlLpIEFrlPaUn
tH2gIF9gkZ/HX0gqszojSAc+pxO2+Bth0M7GgXq3RfRL2Z0itcFJF7iBjBeuBREu4f7PzrSkagLV
xnvAXmUZSAi2Ree1StOQVv0X7U19rJT/QQ1zxdIi8lSdHJonNVM7M2Zwlrj7Tu95u9pxrgJeTKOf
iEJNtVzaS2frkfm1Lrnb9+OgS2cgUpynxRadGm5Da5PdK5TXYZCokV5tFSuaMbE1uQIF5bbvjy1M
1wwt0la/xcu7THxa8T8CD/fl0Tod8E0W3kce+jQ/UJfrTEZKSXTbjXE3e60/P+sFSQGE8wlDBF1e
bchA+WN3ljpq2TBou59M+dzsTedud1SEd2cHbkZntq02KWj+UD/NwIJms7O01HpNUkUt4tYWjLdy
CVSeSm43XZWm3o3hXDZopvst9Zy0rcEA0IgulZIlISoods0LDcsZpTBdLt+Lb0WKIqsz2bcEQPRM
3I4/3uASZ4vcBogrj92iCTpXpTthBdLSjtt6+ch+dhpScx81XMy0NcafZL9UanqkvgSJQ0Y+VYm4
1Mu7QbSzSqsb+76DrYadPT0Emv0eEU8T1gU5C/w+KFj5eZWNJgOWt2YIk/TZCGAl3nKlJsyHg5aZ
7k+8F5C9/kKi/8e4bwfWi6nJSAZJs+QzYsAYC2fA3Pahleuoxc7OsxrTMUMssUYqvWffCPzFuHAF
ET6Evn3ZZhAuRqs2Ne44HKE+NtQluSRZ11EUMUV7cTQwQqqOFALCYGBznmFf8xnvJTdJexn/uIMm
70oqSwxR0AKvyUVUvhSoeERaVJ6S8OUbqlz4DkyAe7hEvfM8dEp1/qO0RDCyH/rs/LgvRSiCC1La
1wweeF5ZSIfmO3ICFAVtLrwjYfjOGDuYNLC9pXnQGYduzZIScpPlzx7Bgsug+KX+/z87Ft/4zkI4
jdQc2I4mifUSCQqMJT/fFd2t0IyuGJg/bcAnotIC1ZDV4XiKwInfo+BHFsNowgqJ+cus3pQo+NCX
/YhRgmVulqsvg8bEr1E/CzW6O6/4/6ud9FUFuqC6uLLEG6whet3wAgPhXyg6xn0kt28wKRupj7xC
LqsJI0zljTbrqmh7IRQfYSBKwG9TeZm59xN6sEpvoBnfGK0m9+LZABAO2sZOkIJZiZEsurzLGNqx
b9dsuLFjzAuoEe7bw1Kq47qS58vxbsipFeUltHtLtz5IQskgN8YJ05PBwcOJ+2fmod8FFq/3oZfA
QyDFuGqQZZwBnMUThN26SwO10aPfHe3cA51aGz6PLkx/m8OXD20pPS5ujpNYrtwD3cgNbBLOMOFu
NhfF9z8+1W/AfSmcapwEl+dorQBDZzeFpMaY7RlHXmT2Qn7dhvelYOv1fWoHUvHA4lL+EA3JESiv
grQwR4bGMi18W4tIpUvW+PTzBP5ItdwPUr+RvZpm4EjFlGq/iwfwMMJCGslY3NKMtVyo7VQKOQkn
pIgHm4RcOfLWPJzZvrmMreCVClZjwexteGkeAh5Z3okvASvu8iVJF0075UcRFn6wgYFrjZ4Bgham
6cFwdNX34AK/dc8gAjPMHpifHAUmG12gsUbhWHWKHGxmjzv9SeUh4s8CfuTEBZyIMUpQWvHF8F2i
96TFR3gbHIW8zwBGdfY8b/ddyFRvF3wmImMQLqS0IudpgBsyna5lA7g7qFAif/VDsXtzM2AOlynI
IItwqoee3bSueL+8as1MyZRPaVqkUrBo7F+BQUAVXJen3tDP/8ECfoJR2XKSWeWn/soRoX0go83f
uBpguC2EU7QMpJ9BNyfyqOSrq4W0DDVDv2sKMQgFjGRhtdn2iGRavGVjjfKKddnroklca0mycHgY
oYSLZrW93yZW4dXsv6R4I/MMrcUy/KYcGUzbV9ZmjJZOFFNoz/o81epnnHfDc4ZVEQ7W7nIcYQv3
2RzWBRqkqa+zIwWgwnewNcMt+vYSHbnUDvYWboVHZ7dUrQa5eATfvbCtMpBctdgbAh7H1Ugw9S8U
ysxir0IiS/v2PgOUc4lv4aFInBT0QzipJW9xxBWBQBF3Ecwi1+1GwweT8EHARbEDPPl/WdQaJjxa
4HAUz3CXCBAaKldahQNK8tQCNHtX7kShd7+Uf/iGP5GRJo34p9RK1AuChz7ydvTa2xuiTHvhBoW3
PnUMePHHAXxFxTWWZdMo0YXnlp3qLBjjVk0Aa7ZQX6PPUDJe+ouyJnI9157hTzCT44Hb7O8sF0Ml
d0myokPzKsbxthU0iAmfEJ17IgRXBUv07y4JZXDxcSOS1syoJkBHT0H6NsHNiujYV3RDWHY7gEL7
lQDtP5zTBcN0deMNK+4R2Tq83RXiU0DHhq+nwD5a/L9ticotGVOiGPIZ/P/oAkRgJmbafgkqSUxI
4MtZYfn3MROHL/VZ0a0YCNdZBVeXg/48qIgAuC+VX3k6zKbfXH+qAul5sRkE7OZTDSzbVLzjIjuY
w+E0YFvnsDzF8H/+8gmyATldA7tnBub4QbPx72Iio76k38aAwW2NQtbligRxh03CVIbsibJp+308
me/K4uX66bNXA1kf2/PsxuqV0x394lhRZbTe21vjg6b/I+V1yc9dvnFf1VsKpGiFuDhyuZHEyoTi
ogSV6sYfGpm1/Coe/6w3mYPiaS2ZydXmWl9BIfHBeX+HE1toVoy9jzBnOwNyJyla7Whfvqu4tix1
QmoXAQJSxlacVOefkiwv0v7mm5OT1Y4/ERf254GCYedARcaFCxqfyURzObkqK3MZP+qzYMqh4SeJ
NEtrlsuMMNpwZGXcH7YoEqPNwrEy/HCfTi0WjssWJfYJyT8kC0HmQCMm2SDN7/FXDz5p1I74OkAd
CIcv0BNQQcXo6dYeTVkPpS4vVnw3Iw/DZsjphBzWdLkQz20LgpMUHwFsZx4pm34WSWclRU4K8QIR
xyX6T1zMKCJZBU0NeclcsFHfu/qINxsITmcEa8ba34nx+Drg8VmY2LpttCjqu+9zp5k4F5weTWpl
Y6ao6NhWQDFEMZCJf2j4fH1tDLU+SADr4Xs9xNo8ohCMJQMofksOXpLZJ2vVvYQiUDklEhhW0tqL
mES9uZZrKBots2DEac71x9btRp+S5HFLqlxMD2Rtgrhw3Pv4FndINrsymsxsXUZt1kVB4iDjRwLE
GzMuckIKITMS55vkol6oPYB5qPdjLlawj/IZy6rWtMOYQYlwQGdZSSVxcziYXdhkXZTMy8R4Gw0T
Hw1VubN4JpNIVlpHpJL5gbAwu1eSa7g4HRk4LcOFt0mim3oIyAx2jTvNJp3PfI8/kHM57A7O5o4w
LpA2/sDmIPr98crmq1/aAkY2NHXTcL1PiQTQQogUKOt65yFA5HjDjypRJkkkwWIjPN8S84eW7Nxg
IO7isxYOtN4g7a7jIRNX6ylK+SIbAal6wwdLCQHEK4qvgYKpVSXNoBYBAXgTO7wf3T55kJfz32rc
R7Q57PWzIau/YKaYvmNTgAeBi5LnnojIAz1HDhykYCisYB1lHPDswnVyTMQAMa29wOCISAREDtRT
edm3Q8kJS0frnTbSAQXhHFmbLXEvihna1sOqrIeqGO3wVPT6mrOymrtVTTjzBrxHrFBlXmuo+xb8
5vzjMf1aqZQ9Dz2W803X/ESNjGZqxyqnJVJRroe4FEmV57xMGwneSoDTFKwOP3tqinOQDYEKU7ut
hKo3/spEBD9HsMnbGJOiKdZ6+SQuV6KIW8TeqwN/Yce2zzpEd1BBUC0bw3fiFOyvfURjsIiwzpuH
sS72xcmiSWMqMMgABrE3+U8LjKANe5BzK7EKINVL5rinzSLAl3qtA7MYg2y94wkmawEFIGPxSeWM
oDQl9bFrMOjDs9LRE/A+qp4omOeXSc8VAriQaTKnSsrfECk2NyemLgb8NLEkldaZogVe5ngQ8P8c
vx0hts5Hhzsfjpwvj8duRFFgpQQMqh5pcfQO/S4OGqOEalmNWlGGiszegC78qF1qsyFscjtnQiXK
J1DOCz2ebHJhEzJpiAiCSe1xzmgNfHu7IFHxZiJ3OeKuuomqa7CyjT/TZBgNyMw8V4LShpwBrMgV
Cf+xLidm1puQuOGtv9vWEJHfBgSP43wWeiSKQq8yBCS7r5HDUMeWc5wMH1FsBBWGeWKV8yNVKo18
FLpjP97uU3j1+Lg9Vv5yJlPNXrEDQW4PHIqXv87T415MMTVSibg2tKTublTobOUIN5ZFS7zk7Zgu
TqItYrWkAsn09De9mZ5tIoCXl2QD1FVIWaHVFcJP1gskt6cWPDeUyYcyTxrJHlZdAbhu9Fs4cm7Y
R30IoveOb3NRxSt4F/c5g5MxBqcymhbCNne6obOedeqj+Ea/WDhaI6sT4d4T/AC1UFYSXN14BCka
8qA9gay47kW9/rD5za8nxi6YOPw3pYcx7JvbPlZiON+VMh+MalPzA5Yi+ypWhcrYagT3SKuHzY30
MD2gStGjjy0KOBVdDTi5WnOuABWoqi3cHmYS0cgG5ER1oFq993Vl4B4t0S0xiMJopLxHTPQNFMcw
5RHAhTcEqyCS/THagkXuK3ojRoNB+Jdsn7Ec4z/7scna8qKiWjd+MkX2B7/TyZytYbAv9Y4d0yip
SEIBjfu3R4afFeXbyrFp9QJzEfkY0avxO8UMERBGW5PDNa1gqgYuWr4WXy2HcTS3uXSfsahBrI7d
62k/Oribzc4zyk2vldjrc5o4eX/18YhRDyaFGBpbqDmGFQtkvg0BDRJilcU45CsQWMX49GIdOdF4
7jsH1GuZjmga2GUok7l7HBcEnXOatnAAMiZJjN4K4PEmaK4m2YUP3afp0VlwBE0nMy43Ae03YbKd
1tdUzxT7Md8kROPaP0tJzsl7X8M0+CYHv97L6ZVB9ujAAGNBQeMIjpNIDRQMXe8e5/2MP4JwwC9T
PopmFvhLXHbQ5esqzsCi9ovrNCqQ3+OPWtNp7Gow5LOXtn+bfr2duQPthbvYgLvs54mLxovXLZmx
RqvbLsd39Youn1hQSoFA9qJ7b5B09LvmlSF5+bmi0J/wT+CBp+xCLd9XofCWzJrblQLYPliQR8gB
R+FoZcF5iLOEa51GCadgc5nveeM9jAC86nJ1GBO6LlHlzwmIA+WlsQPXfrQsMWtPQft8gASXk0C4
Lb3xfTHjO6yJNM2vaQUY2PejaPMFBJ5CUiBYmJ1Dm7+AnmThhax7erlDwoqsYk/YPdlbUdTLAwri
I8SQf1OE+856P/St/78gG0Zw83BHw+Ut9o+Ew1Qr8nooqiYFk2cbDdARUGhuSKcdynI12TG4CQHm
YWW28KyxcG+q7cHOLlIYEwcvftX5q8Uh2LDhVy2TNwapZ3JEuuMiWKClv4GqUwD8EJlqqG4mhJSV
XFblNPiv8bw7oGdmdOsfdUoMYndCBkz6Z9plNnxXQL51ZwbFdWlsnTVRFqlInIDZGCyqAp2HoYQ4
OTt/NSI6dx9kHmTUrvmhI1Bmaj8jnsqZiZ5s76+Uvz7wouJ49k+gkXRNiSi2LLoVn83YhPRzk/Dx
Ch9xb4fpGZqBZNUxLt3GA2IM3sGY6gH0Mot2tIj6fgBPyJo9vWHI2bfK6liPGZivYL5TYbLZxYx3
buNt21WqEmGqy+1aSYI2iYLRdDp8RAZTIrJq7mgIRkXNUbt2VizElk4NA1Eh3zuBbs3RZC6+bvtw
YJlydf5J1up8r5PkxYdb0J9C652YI3+88MXteViQIbyEuIWpRbAwtDXsHVdP9cDDiBo1lNcIe8EO
p15GIj+DzIVJG3Un1W+KjpplTqnoowb6oP3iGlcQmbS0ylqc6rLlWbc3b8JLG3QDlNrQ3pHcwvUS
19vmAvwnW5hMT5UbiNFJ2tjleEYFOw4UaSUKLT0sGk5aQMlbjeJ8abt5cbjl0ySlbB/5fEuVP2/g
naNBmxAP+gKtewHDzHFCGNWVEp9lIfJqplFPRReFUIbJrLf3j2mhJ/J4RCz++xHdnGIXDmkiHgNu
pBJAiS46vmqAP7Ob7guHVg5bwhAykRWAWPKKz26jGcivpy+RIH0lFJBnjK+s5MfaVF3IcpJ1s/n/
bQEOw7F7T0rd7ipux2ENHzreYBaknAwrtQjHoEVS/vHRoGSomjegAQdr3EN2HnPfYBQbEpwGKzoy
PuSrrHpG4oqKOwOoxENGsVyYZ667tOGQRXCd4H3+0nH6Xr2fhql/86+ob29WDxemyU6FyK4+OeRX
egs5rhQ6wkCnE+77KEWNSi6oAavyRvoW/PVd1+XQ4Ft6gtYi7Odz9hAICKMNPtdP37qVeX1B2UeB
20J7vlA33tdermj15Bhyd2JPApaXcm70OkCuZJhG0tX+atzC4JGuGMr14o3c8WsFuuVw/gvk+eM2
0mRBN128Dvi77D8x2HnEisnIWQRUBotiz+KNAdSYmstBmPDvu0o9ruYcdxR1/3l1Wv6s+t4H4x/v
OxOxkT9hJGWjxgE+ge0i/9FuLveoL/nkU++ZA2sbsLTduW3wrMpe6KSWGDVSVInRbiP8qVz7/7dF
PkOYbzJ7ag9w0LpewZj63JsR0DMYUObDLXhzHXl6slz3w7TboKiFwslXIbl37X+4NTZcni8xBAfX
3ZyZ40PBDJUW8ALoz9O7uC7mjSCoerdmLNRdxMGyDbXuU5A/C2foakfsi1m182G0gZCc4QXtNkgk
O5JeedBRnU6Pr00MifuhDWsl6tieAR7xARBuBXtTkFTOfhbp4+WN/bOjtqCMngxBSFiD9fzZNFbO
slEpi4iOTYPcsojVGXJoXdczZG57dR9UgEgmVMkrY31Sn00ULwGyJnzpaKy6xT6YwqldK2FwlEpn
ALhlTCA2/HiXJCp9X7IzjlDffQwhkQxgsheZEmC+1XsnButhq6l1AQ9naCtZLr1pKQVwBsWTRO1n
kvbig1d3fOs3hIYdjyX8ItMP7qd0x3sqGGyjC7DK37kiGYJ9aMg9Gy4RoWc61PacyPd2O8Zlu2Lm
N6lG5iys9yHdm1xXLHHzfogw9DVM8lWAPrjJ0uFMOi7zBujc18mANegQS9fsr98HCFRpX00LzQKS
BrHQXwP+9vaNMVgWPAkukEDMwUSPcUAPH2ImQre6HD6gpBcJqW/3emKEQCTTBzp20ocCUpTR//+y
EXabHO47Q1cs7mOMLjjijOdifsbBOZ4X6KynDG8aEtkSPADDLC+mn6Duq+jVM5hgm/CxFcpnB/Y0
uS8DLQuJyxYsLHiXqMGWi1ZEAIzWKuk/4UvBVTjMnB9PR8EaPyc5emfbMyOuVKD97LHjOoSlQ1/a
8UcFYqrGEDv4xNLd5U9kfWpmhg6jJLpgSDqPr6dekqjyhSrOK1FwfE0dh/NHxjltblhMYDg8Iv2H
pagTlWZa7CxTiRjk9MGcnuCn4CzxFza66wyc92H1w0SM0KlXJTrsaEifm7tw/7At3PWhSo2QprAW
2rKfbd9HGxGWNeSXjF09W0tfn7jq0fNMsR/u/FkMQH5n/o967yZh9SZLzpfnsvZ3tUBizkf8uH2X
i714oF9ecpl7LLfZaREOzkTrUqKLKFmdXClHzWa3PxTHNYUA7vi6GxRVNhxzzWON9Pmh80cnwskO
BB0iMqpvRObynThscaRUJyC2YcYdk7qdmaHQXsVLI1Ii9n/p2krFj96mlujvauj1aTx7H5hfxwjJ
9pEIE+s6aZawCaI8wKDxSWKu+reMIRzBLhpKaBnqA4a1HSlUEJ6+DDw9PDZFqPI4wOSlj3/9L80e
Jm9+DZHlPz/NXgNyvy/5WbVub1e6aGgg451OdWA9o4UABljR94zI6SMmjL6zaSX0gYmdFEjgfcyI
D+M0u+35wuXd4ZGjTGRiS4btRRR9Z5wl4kcvPBabJTj9gVRW1MPzUkAJ5DnexejniCmjsZiEea+7
6YAoMCwRtWDznwKruIytFycq0YQV+kr2hXBwLnYzlhJ/iz9Pe73SyuXkCoHtA+moPi0U0y53vTeO
zz8xkD0tpN2T8j8KyAbURsE+rTDfmwau0fmFMycbHpIpHLFjD/pXDMTx+meDMc9SrjGWAG/5aL+2
WRwqtYPAhE/OiDKozd0uVLIu/RsQiCr7KsCXtDgxKERA/kNdscfvNazDEHzAv8GBugghMfTYhtVt
jSKQXHOGMUGcYVf2OlH9B5UscE5yL+DXLmAvAwsfvuZmlBCcihV/iyeej92fGrRBLPNEmxuIKqqa
rld+1tcCmuMFCppaHXV0LlzWUI0wavkfkpftc04btTlPhQT897lMj33qGkRUy6fad/9i0jKp2gpw
l7hygz76EaEIC/kUmDGqs2Md71eXPmDTLrPAdM90k3yF5fq/Ca8S0kQrOm9T2N5v0J/4UmKPzCRZ
2bFvO09If4EszBQHwll6VncSdquSpydncUgqu4WBDs5K8Cafzngae5+/wINg/zywd5mn5cpiPRvn
QI3rFrykzMfbQNIB8Pxt3k2fq+0DWVBwE30OIlPP5/vcXx/7kc9cKJClDkNnEh9DiyJUBRJDR3hS
gU0k/v5V6gth80tSp2HBbeEO2LouU3JKXm9aObcArawfAaY9Y7NhVs0iq5FXoUgIF5ZLMiCBH6fC
xnq1ABXa6b6nbotXe7h4QKXP4Yfhl63PS5foxiODtf8Q2qRiMV+0um7zgRHWXEq8pxJjdryCIeKh
80V8hS2+5eRB1FRNKnmklwhWqd7AjwTnQ4CuYpyuQTiha7kBMReAvHSKAIgvPHWAboePsTzEk9OB
nITaZJvMfQh8l/jaUAlxc2qL4Gg3yNffTqtwwEXgDWDaec/iB3WLy4ssSYuxMdzWLJiL2MHosFCR
iKSo/s2fHnfW9Lo1EOhXOuNuuyK9sbmenCuQPGS+XyC9iYXr4iyH1qvusw276kRWU9XUK8XSvJ+z
DptqTukIO0L5SaIglr0uYvoZNwwHPh8VZq2l0Bb9ePKjpHTNHhQDtLtaDcggxdpoOcxIjPpmiiiQ
PHaOUTE2fM9pXVitmdQd09AR1fW2veUwNVpOWNo2AbIWsfadxe2Ud+SzQ8BgdJiUmYCUk8X2fE14
zfwl+BBzPEYumynYQvTwjI05ZAPAAj4zJHSoOm6t2T9+daP8i83Ugt9FL+U6zTcr2EXZvbEtU+WW
FnfMUjLee2/m+X3S+GE4tLA/69+SEsGComAZdyHRLRXMm98/XO4Mlx9sI09i8DvlPJNZKONBsgmj
EV4f7ZkQ/KPN41M4PyxqrYEZJMoNJmB6jLqxTSS/YbdHZaB7PLlXbp/Aa9uXTnn1OJl68wn7gGA9
YF//Aekh9Wfeqe3frtB0Jl9TaLzlMSi4bZgIQkSoVfGKz999obv/qMP9OAybTrnx36zgSVNW16QE
4TXSKLZdXLd5HELnB4mrLF1zuJPbJczFPXD6dbgphwjFpjo5YbrarzkRhgBAgkl6rtFZvlF4hQtW
EWNBsDsN07V+T9EnbvUQ0V7o97VBf8NZnAcwzAvd3ubjNS7ZhOv7SJZpRT5G69XKDB6Whk/KD6KT
k1Cu9Vg9p41q6ERBLAIWK3cN7BNWl5JCOHYR3sUPVCdQvnJGDYaXqfqFBCkY6uqTpsPh3VO39X30
9eQZ4UChQzWRwzp1qTUBER6XWJZniJpxeBcFKTAzZg/kGhuVr9DWG1lY5iBeWMkJvDRBh8gtTZjm
za0DuAsv6WLZJiFZh0KhdODniWHh7+cqU1iGDqiMgEmAhj8wXqRNNqcAwqGq1SYD99hMjgLdOprQ
vtfprjBzpLN7MrRS/K3bwMSepTouGr2Wtb6LqtTY3JWUKbv8Mw0WAmCCkSunWNLZyO76wburHnhX
QCXMle9DZSCjYkWQGIgA+t1uMDwDH1phUxZCn3qCyQp0JF/GyEylQy8OW2rXmml3y0ZWFz0YAtZL
O9vOSt3tGoILGEB0iX9EhexB2jVlXAu9BjAvvJuRJhC6+d0jobf6aGJcEbOw1098ZcvtE5Mh+ln8
93tYIx63D79m82/hqaOSETkyDqE+YVXWYVK4wz4G5HVFYkbeV/OZozsGtYeP7RZEyIJFPNEJ1v6f
LjdHJK0jJqJZSD3/PP4rJLA1GaZR9qDqmgBehy4a+kX1gZISjg4hTCB+TwFsVIHIsV2riZvs2eK7
fkLBg4y0wYXDCvgSLWMIqqmpO1iCe7YMKOV2z05A1tAGf3QICTijDOCWePmB7gXpo6e3PZ7T4Rdq
NIRTWYfHR4Jcvhy0DjQpIZ8R+r1HbynelkvRA8DQIrXoHZMRVVTJlqvzJfxrqL5RMgXGulmcmSC2
xR+qk9x20avVRvjgaVmv1S2LDN46LfVu1LNFCPH0Zt3SV7gABpfAQB6ChDg75Vl5HOi//5rA5tWM
TIWu69idTgfWlQIvd5jOYAuw6y/3ucDSJ1CjVVcLi+bme0I6bKT72f0R2rl2jCrwR+lIW9ACA+QD
xedQEajjKB8TU2J0+O66gHbQOJnZPn3l5uSI2xVlJDHj7AHaGhDwmKPL1J7su+IFrTVpP823h2jj
ShcrXz4nw6ZC+WL6upKaYt5uDvA65hGKiPFXU8+0V5bbQWrvEAYQ9/EAgQp1Li9JNrhjIlkpYqOj
7neeS4ThIk12iwmuET/tEqgNvsY9E9MBKru2PtJ/ENmdt2kCz/yzo7TktqqOrYNswjrMo8eTSmCA
ZnJsqfU8qbw+3PMeYtqDPmS2P/3BZOWanslvMIoTeKCts6ar+KZrLScH/fOCO1oUjUsiqY4f8i43
lXaqhrZO5GlwcPxWNJlw2HJeOh0R02sTpK9xvK45YFlSXBCoCseS4L14zN/fB8H2tflroTThfw97
AN6EpVhkh+lIWyDCItXzCPPzNXeE7ZHvr0JJsQzD8i2001aR8zIRisA69fSXukP9g7wcW9h+3o4x
Vh/DxiW7fbn677xdZ40kgDdWb7DcHbU3ED+6vQezcBgSE/vggNH9aT9oetKS7ZbdnbRfCzlv1lov
ewR2sy0qhAzgB2ZNgOe96c/kbEJ1lD9eEXylmRnMy/V5yH26hLv0vD6wJsewd7LDGNxIoic/2THS
W1EH+GTn4uCN2KIhcb8hiDTjuNo+AfrgQn7OmcAu0AjuSJV0MRXgUBU5/yViCkrgywGQay0SYh5V
wB1a+08E5We1p8DwGzAc0pZ92Opa8/NHoyubFDC26MfES8kYckaJSyoxaFynCNw9wSeyb/6VmWx6
louwe2VHleJ4f4jhT00Efo20254jUNBhtIWfrMsd2XyxOBiPIvIjAskvlrUwVWbIU2NhlsCKYKvR
Ao6nwIhCxFQo3tGRIf9BwTNfD165SBb8/ttkPJmGl89EKlcFI0FwxbkASfmniCMuSg12VLtI/FpF
diwZX5uSI1ysVhrNPm4Kdc+L1WWLq75WM+fyeCV3Z9qlXn77syW47OfnYc72lq8akJzqJlxe/k8V
0n2j3yp+s0StMsdnPTHh1p8x+M0qK8iFLbsme1XfI7DNBW5YZDJWlamSvUSmv40QmFadN7CqVfnv
gkNE6lIclnmzbXn4gpPhaRUEhG+Lg2fcOlQv4GbCMstJ7UsP9hkJQm1edaO2eOphWBRvtqjAxyZC
GgJ/Z+r5stFezKUsPafM156DT98cXQfdBOoBEWFMCyifL7krfvdVZoGUJFcEib11BXDjus8RNxjB
OuJcXZiMnjW3IzVVuLPqdgJ4lKWH2Ei6RCEIjExohNjq9qh6dqUiDvmZyotW5Ksb6BYWY/L/BLT2
stPUCYJlvhqMHfNewnOLqc6XRG7bdSkPC68mx06ILTw1fknQ0SrZYEJMZvV7eAzvSF6+ef617mnD
ET94Naw7M+C+gjPTHcqHkTnRtjdr7I1KOO3+FWrxPUnujpokBE8jrAQUs4zuJXzmgPXlobH4eFif
dZrJ6M7UrlDNHzxyJ9tvwwbYlt8YB/JM8bYMHNGUIHU8NMwEOaxs1sYj8YBMDM4rMk0Sz0wGz5Cl
DcIXqwmb1i69/tjEYumu1ixMiCzmdaStG7WPwyeqQ0QCLVONhsNjH9WAMUjt55W+3kquaK8Z2kqN
/gQX/HxUVgQt0Yn8Kkuz1QFhtSrpsK2OgAnl3x9LVZVZi2FJNnkZRmTqba/3SxsQx+wpZ+H8RVkN
e87vhBYrEo5rXXXKzO2Lb0jHTijZ15Pn1Q1uW55ggvPb/A5eRb/OiwCrW70B0FAAz4HIVEY3XmJJ
iltMiWStcZtzDYE1BldSumMaWSSAbO6BUFby/knHpm28nnILhH3IJCw0thkK1IdEWVCQbYUAMS+T
9Cm0tycBDKJRBSx0LU79hOnUXXPIwIuTG+eR5Ka1JFnnMWVXfBP33PHY6BzvkkQVXHKBudjxBp84
FOW1d15TnfJi0jbs6rv5Nh7+XCOsN5avemxQwLYOD9dcbhi4XCajip8uCTXMERDBT8YUPtQzRkOD
sMiwUbSsrf5ezy0VzdTCm/VVcrs8Zf7TRTRcvoc+4nBpTLo7vzwdkW4vHq94Sh5apTIzwoniSdNy
cw09cBA9wdU0ytqdxixJLNZ45Kh+WCw/1XHrfoQhpT17Kshu8/pO6nXeYA4knmzh+qs0P4bTItHH
XG27Eytai7A6mmfizDJPxCVDjUoU8C/Qo9fmKH4xLAbVn6fIhJJ2rRF9oDsA4aPQJrKhMbcgX5ep
hhFLv1im+3RrrErBzWTKzyzpYoJI5RSOzgmrMBO7MxKAzCbmm2/h2pHBi8Pj2LeYdAQhZj1Dg8bN
O+yXDPinPlr9j0ZmtmQDVXbeztLrl3gtz3cWoOSSjTFrOa7EmlM/KY3oWSW/ag8EY3Yud+Sftoue
KhRXKaNE2MX69p2U0vJtskVEA6AdBmcvJiFQxxaWz+sRzYffE6WX6mWMJhmVXKv2bbM54+1n7prD
PT6GuRcYp2jDRTIIJQE/nUM1kIDjFHJUCdUlQT5Ff2BeimER0t8dLI0aPpCXd04xt1QOYNe+ti2F
6mtKijfDMNI4hxQ6RiNAmkV4VwUSnAE3XFGJDlbUBddBmw4VFyIxXhWruAqMLKGJhmBRbm8iiC7G
vhRNVsd3VAPkEXLqdmnFM53qQoWP0zj9cm/mPy++AIFvwWF1b39um0oATQy8wmJF7bs/1dDZygpg
BZP+FtOa7k9Itlb91HcNACUVJWgxcQ0FMtg6EOrdq+ticWBAzkOSWra4+RhIjY++QDv+5iMlHLLh
px6zS+qB7YFEYOB0Fd0ppfGx8nSromF9ci6tejUPYBq5HX+bD3+m5mGbiCEdieMz0HBUVLNYgy4G
JkvWGp5EWvjgHa3Qh0VGLbpX8ttNkKRXHV8ybukPMXJb9kpdvq9xtqtBTFp+JJFN9PMp0s7EzapH
pEX2wIb7+tKDiJnns3bnwYqBUdTbBVD1wunf1lrQMD0yvM8LtYeg1iTKI6vRbytFPL96SlqwY/YY
LSchbGE0r6zvsqjww9VMbGh8t7kJjNCzwPhmo5h+e84rfWVyJaS0jEMT1ROERAe36zMX8f93jGWr
8OwfRJXPBnC8YAP55n7rOwZMhjoNikYOGrXY8eXh1RWHk1hwDF50l+yVj0kwBpYTdM2gUdrj4/Iz
D2S/jUmUFE7DK7cBGzMRNOSlH5jGRUTheUoKyauIeVN3iS4+tYLQ6mQdZgN8+3+O0Y0YRMySRwb4
3cRctWYwSUDbniMimnZuUlKz3tKLHp7dWiEdD5e/ODil41AwWPsvciIX1g8taUALnpGtiT8VTc8g
lg47YWFnpnkQxnLKrd4vUFbywJNFYk+iRS2hEfEbMlHYHp7/tLq/kBveItBfmWednGj/lbcyDLU2
27uEav2waM+M82R0Y7mMWH9Tp34aej9QMbsUBE/MOC/Im18KfvplX//f4PGaZyTy/v5daMbC/OWW
JaNZEKEDHRIl1DMUBIGsxUrHM35Fybc5g03/DvD6x0MUHv7t7U873ui9EsfWUHOcl9Pp3dJd1UrL
UA9tncajm90/CNB4PEnZWyatTUD9bW29tiwnZ2Afr2K0KbHblUjNetrjIWKpZ0ZSf+UVLxStDuAP
dAmYjPwbELJIuasGXXftOdaHi67/xcEXs6RWejRF5rjn6QbvmGwHli3eW4cSWVf1FN7VhpTuf08S
vwJIMFCyGDEP3s9mL21BLDRZJRDoz3IH2LgaX1dSxngFSzWm4hoMpoU0jyXr2rM0PLR07lVxwlqg
sAa5hqsR0le2FDsyZhSj2yBGwKqiUH+4zNETY/+rr9tUZH/SpdTeengiqPCXJ0aqOc4bYVEX2EyB
dbA3ZDn1rxE5ki5mtwCqhdiz7hFVmN4ATUpPACNibftv37qpyen87t1pqt06JzZn/q5gP8LkkF9V
fUC1XVgTXrkLXCfQQOGn6wgN5tZa4Ezqp2NjecwJDYNCIAVG1RMAkyTjxwelVOppbLLVADuC+cXK
bopIWUjUNxGRSdHKOVe7VYm2U1kMog5UN9QsuucIEO1KWM89i6WoQdwOQ0bTWbqPMMyWdHEsYujQ
qyBAAvBdlCozWW7lF4A+4DiXjI9O0DnEdv2FXlKaNqfKs9qeQOWrH4ppAODU8XbxJpJ0RXp8yw7O
fjdKDKHhzV2PcLpos5dWdwz1dY9rrnzGvP/thwywB3b3F6BJXautrO6g1MUt46nfrDPE5cWCMCYO
wkJjJzXaczHQhtrx9p47RQ1DLKrla2aFXVV7F8QpV2YKYQ0I3QNRcg6FLFWJBpQUelhCjsnITt50
MDdaV89XdXpctA0XnlhKSn1eR4G2i0miOqqHA7mX5KULt1fRVzYECsmqPjL/wAFxkTgPaO5jxpVw
mfjCO2thPBdDxeWSeMCAa9pHEPUzKwh/UsbuqJVhcVI+gIFv4WSPOXfSux7IzMIgeMoJtWbfXnl6
ljnImnrLYayQxufesJVV4LLW5OT6292LIKhrYoLvJ65Rg0BQiej55Q/dtMi1P7D3zbDoJWLjrzp2
HEJrTf/9uMSNhUfZ2d5U5LnSwtbKMH4Q9VfS9sXpmWHB9bylumWbBTbpzfsBHRuiZQOYEEoaZzBL
WJHJ9BQ8DfYvkCjQ84xnI1eEx2cLPBGGRNS+wERXpnvR9Oa2gRe2iMiiOVPs0cCOzx2vVGXGxj9v
ugDo2r88RD23EfNEYOZ5qBspe+keKYdCjlSbo9vmFqI/gI4qVjkG0cekTrlqeD1CrRf/Jsa8lhKs
oxQcLmoV4xPFTQLrb4FSZO9X9al7LmEn7d2BY2hdExHamTOL4MS0V+u5IE9efD2fgrNWBN5qYeI+
InPwJSxOevoErUo+RvhEwsw2OwKbA/f5YgDGFyTJikmJASHdKSypVhkJ+L80y240BJOd75JjeWqH
1goNkBWVCqmSoM3ygRAPGlUtZwDCCeczvt4GSJQ7bn73O5j+M6bRjou8zE0BWVUO8W4B11nhtJT/
wvSfDKlX1Lfj4JXnuakPaGXpvd1wRWkCyUK5JzgHyLF28M9OQVY1/otL3xEpjOA8HecrU+gy5IMp
3qwG2v1Q9yJBpKRdh+C+oXr/36KGY/IcT4OQOMfmo7sCLGv/pcZr/6rnxgU/+S9S9/e9lN/sdhg2
HhEWMfLzkNVDHSxchJqLNyBy8fQfFO29I6SO2UgaSXoSN0MovFwNRHbuXukqC1uRj/Qm1w40wEOo
n18y4jxa4Z+MV7xePgvGrBQA4/OE2A+oyrLjDU/bSyzBNWQ6NvXnELTa14cvgZFayeQQbrhkp4D8
U5dU4ydDPpwPtvs8oXRL6919W8MtsFhLbJrQV7jS8IDWVMQcnhXJoGPNdZFr0/q71BiWpLc4xHmQ
vEvvaNJbcT07gw5bJNBTgOzLN4ENpJCa8cY/tHXmtR+/t/mmQCid/sHmiLZ3GkWSEfeXMhbY9vOV
3X1FjvBBZfghcw6Hog6ZYKY2MiIIhDPtmK442+iN6JNCE5pIgpxnMDld6TYKdb34mrNpSidwlkfv
dzzr+ZXNT+jLuEncatrJdNxUW9TOOmriHQFM8dE4V1F00fDO+vvc7mTFpIgPOkPjhY0REzHaYpg/
VgJnINa+ocFLErr48ZeNMHzFHNGqDNu6/6iUyxrrKYNJIuT9kSo3lCQBx9y2dT4XSk+VrV9oEhHP
2TjpxfPQSpDB3AsQa+5IpPcYenSSfFn2ONTLV8UEfLuUZd+ws01JTPugJMJX1egpW18bdhrXGfAt
7E40lQihh5tSBb56zGzS8hwe/lPZGSLqdCd7/dyvy6G5xaFcdEU89pLVge78iw8Vr0HbZLBTGQJb
yp3shHr20SIBGvuluSHc0vbtwOOGC7rqjFaUUWgpJba6hi0Rh3nujBqpjphSlyuH2+/vTKLLBIZf
ec0nQ/bZRXfyS3s2hnBb+ciYB9Mrk8aU4LD3zoFr3+g3LaNnfVbPejtcmPhqRCytGPmfBC8ZCokA
lPI7Brp0AZIIV9AuhXEfEhMxPHxewHN+RpQZy4/CaJcN2MtRw+4Xb/xEd9jlmvGt39iKFgjQItA2
iRs9WlcwZvAZXPxD8SvsxchdMEcT//CybgR6rK+yJrewaTHnVYcuwtDV6F7u/JyMsgdT9PtwczAA
1Pz4puivogSTaXTSMCFOd7xyAUfkg6U7ndKHgKNbPthX1kT/ac0lqmQPXCzuoA8m9cA+khYJYwMw
IWM32qUQNGri8gVPiZSVkGYSP3FtmUbRM+8VmrASCW60inqDOdTCk9i+WF8QdTvWX7+NLGKGHtUn
bWtBgjUpz2BHWWX1swi0biApyIVnNa6hsKePT7o0V8+ZqcOOJrc1JP3k9z7ZlwGhmGxYmuahOmYn
91i46akZo+sdXVirycCp4Zlr8X/VMrp6AnROc7mmn4BTYrr7BYRKa0M3M22dmJTrfEA74FRo4GLZ
c8/ipLgFFups2r2DklfKfecsc4ZKKUzI0b5d03g96Oqu8dp/rQ0zINbuzz44rfcsXOEFTD1PIppg
cH3gxjbgAUbGvV0vyPISix8hWKoD6AtlEm2AR3b5m/c/scAyGAfNpQDjxZx98Pjs15SxtKU8TNBp
x8sLNCgKw945x3dtRjpukf6lHdfUsdYHMTD68r3R0xIe/y724Jn6Y2lnsXSvn538xCpuwhmjVCZe
P9O9S3UTvWnHPpbuWDDe59FCu2y/S9CnVGtvSiYXOxJuMxwQNHUxE/e3MNsw96M/o6cVixrh5IYA
hk8oMXjOppDmpvtkXwiB13DUeT6wsqXchdHMX1gCZyMGWi6gbFkbg1LWvkirlZMtGvJb9denlcPp
OxRBGCZV/4dtL+SX3kc37xeKq8aSSCPaDWCo38qD2q4HjEEsvI2NuzgxJUJieIJiA4Oui3do4ner
0wUQg0OSPcjsWAqZPMo3Yac+KdqIhNlrE9fMkLxVsLXca51iVGDcHfTnJY8Tl/HIUO/pGVhXwabq
IU3A1ceuwiQNBPmVBeJNXbUkNdo5JkIEkr2cglMvGK37rrVoQUyj2KxtzfPCPezN7RhjHpn5jR3Q
n7dexgLOX0Y7tMzqd+/BS/EM1Zkoei+F27MbKFgeJ9tqJ4eY3KoU1oKe1u7ishQRiIr4M5aa1WiR
bX0zGqJsxqx7CWtptFc74mVFg6wAsJnoqS497GIXVHqlNmumviFeY4JwqTZJhJJ7Noc/oqmXQ4fK
UdhiI4Vyj7CYrhcfH75Jb/QMv8evOsJDBav/dbBRDrTUbTj/NbWFdcV6TxDnLw7GXJKuEmwNi4Sq
iUktO53ggOWelhwPTiEZqnMky9FbNCdNXo/4MZmp6mauiieQmazeo9Xn/YrgNR9apu8use1rHIm8
+EDp82yFKoKLvB2pJj2CVJBUJXEcUutVrrZTWrO6Vw8eebPDOplfHP6WBePGkGYxg36+CyUMgWaY
e1iJQUOqkkt0VqdQKBfQ4wg2nPH2CrwAEDMdT8TjtB0i7F43z4dpX1BShqbRfqITrFWpvvDFls9o
gBZXnwSs1Y052CRX5YhwwIiVtXtHhZ3Dd0EGApgjuGUgFjebcmqzYOZRGS7DhGzHmEgS2XCZMzoK
rC/Bg7wAHUokkxsTTZsmQHQr8yDtVq/cRLG2uYa7l1krdIOgjrA1FE5B9FkbA2dtGGEDW+pRgx+I
iN2rOIhFWFdcOaAoez5GglkQLNt63FlnKiU13r/QDR6/5wa1XFSSPOZfv80J0pRxDtAtik5GEB8l
8FE0zEKCLjGOrGXNU32BooJ2N53amkk7VUraJi1ZHEHDEzzEum3rpWyX+nOhs7HLz4DNT83cw8Lp
jmjHpim378DSwyzrhEQ+FA/OtgsXolJ3x+AxLRiT5+pS2b4vd5VNrRMqs4w4pjK35+7ng4u5QeaE
AVKOBEzdiNTnI0H2yNe/GfQLRWN+6gu2vTOcIy7E2JpPPSgcCgkzJjCPLAHV5WeA8pdonTP9bBKU
HdmsL9/kBV3soLX2+9eSg1qIOgQ6gtyIruZ2m9gRYFQvXymV3U4BCLTF6RjXtbMxdXaZ/gDhAcVG
+mhMdcoFbEh61ti/FOJh+ofYy2AZjsGg+XgBy2gANRJymZplzZ/BmZCvp+tP7Po5d1nyCDDOiMLv
51l6Sn6+c48ETYxjbu6Pil2bUqxmWWp8586/dXGtJcITeEg4sYYpeyiuvmnwEbF4YsfaWn1jAtul
/M+GwDcsKgW5AQez7ADW5a6H7y2LGdjXP9Ydoz9VmwOUgkmifkEVdbKoy/DaAAthQ+qpz/uaz9s/
VBsSl32iZVyf4Ax9V+xd5QJA126wHg7CRXDvGTcOZr3LfFpXtOuyiy8YCRgoE7PTVnjL8mDhvs+F
/q4lGGVZN8FvPmJHUXVcLeTa0AZiWKKk6o0ids+Zrj6aO0HysuRlbIM9ixcL0XoIgjOKTHV2jiN4
SoKCUBm9xKyO8BBi4J5CFEbNXJsrUKadJYdHeb/zH8uT8nji/2QYgz2YvEaQLzaWwkkGwbQ5krG1
EXSkvE6REztdPk/XcwGKgzmJlio8Xw4oHrqgFXhC7NzVOmzkkXmMRMlPMuDZCsC6VTT04d5x56H8
ca8o61mXe/sZK12uwKYx5qBB54EMNizWy/uquOXOq75/CsWqJuN8Z3IlwLO1QoPtk0g7bqldUUaA
VCLq6pMcOjJPcZSo79kRwAVmF+huQspl5aUXXcKWg7ngGbq/xufOxu9exq+qQJKZ6DBt511nfQ8o
WiqkBYHKh0ctowv4IV0+CojliX/GxB3Gj22FKN17x/TQhvetGUjB/jU/gmOLEOwKPOty+KPwcV+M
UlnOT3q0wNgKu7RjqDePqzy9/WHoeIWMisee5HxhsMecQOaQLbk4VB3MGc4M008GTSJ1P5u7sUL2
QtrPNtUwfIhwiw2/XiEVxp1iFLwPn4IhOwut5oGzQ33K16Gy3ahxHHrwZa0z9ZtodkS531jYHH30
mrGHu4tArKthsC0BTpvtcmhPQEG8QZ8YLSJWt0LoXdvo1ZS1Vylej+wmq8RKpNu+mkCBDN1HvP49
pJ6daswWxBVoOUUSif77pZXW4mi2jYD/k8XmTSwNoogABw9DipVUdeFz3oedSaC+zlk83IZys5u1
CIPX35u/on0m2+XhE81qs40JH7KW7KzaUVmVYIVDaFzVmLeeY71GaP0h8bCs+nVvNvn2U4OB/Sth
32Bgos8o4ErmtEa14t1iujdEGHlNB7gAoFrLhnxAQVd6MxCWqhjLUE13XZNkGBMncv19/pDzvEOD
wjO0DVKwhPvv3Ky+ZyRwIVRH78uyrvOD6Bc0X6fdjvu14L2aEQOpT864f1jXfZR9gh1xK0MYLbyo
YtM9sYGeCjIZGl0jj110tLqTFJee06sAKVgqibbrwtc4iVg1KaDBWQDllTDE5w+QtGk/5Y7ia5bD
Y5nrQIVv53paeSdidocPu7szd2GS9cbSOThJMpo2ZWNH7OP1H9pzoMKx1N1sc/xiNzfU/ogvO5oA
jN/6dHoT6J3emAcTMLoHC84kS4A78nAMEMgrhMTmSU7t9teJ6Mj1OyeOlXbN1hFWL5yn0lWpS1KK
p0SxzHEvl4z+VCZ9pzx6gwhW9X7vAk2h+gm7EnruKSYe0a+TVw8FeBKZS8AqUDzwbWnjYtCpC/5v
lMZ46hzZFWyFlVjB9+kavzaVPkphaLgaSHSkJ1tiyNHZhKz/t9MbSalKuMPlubN5tIne1JqjBTxs
8AbnVmPQNf5UDSyLFGeUlSEWzSj6LHDi3ukn0xtLw+VEA2S2b0aCi5Sh2Ow3lliHmea8umhf91cM
IhkI1Al54mXWJOrDVaXEBmhUMMJ/+wFqoxkaLGcKQrNmv6dREwyRpmDQKEHA1cO/TUlXoPqxHa97
y6r0zohglZVfT1gj28lHuI6YBD9yiFCyzhUUsFO93Tb+wVbi2xfzl8vBa9Hq1y/jqxdjd6zTyanf
IEOXYPrN2aV/zOCPRCVOYkNTY2++O5X/ngGpOD9DYQTumhW4xV3P93wkEqd9tBZo4Zy+Ly5oAMA+
DiuRPB1rQZuN74sbpnC4Y/PvVA4yf3biAW3n/P5a57gSCjzsAYeBNvNHALZNfHTn/N9TKSOGwXY5
P2d8hAlVM+jJMGP6rwTx65em4uTrK0aZuELAU9QBHkJGYYdysGrKsAHvsKnlPZm7Db6wbVWM17Zy
VjfKTmlO8zFZjwx/6MrzkmWx4ljja1sm4VTNP1dru42H4WlqwtP21W3+zy0tZ8yEj4nMpmkZ8XN6
+EVUXqQ5R5hsNF+D+R1ZXUxT2xaSwk60HVQerZPtpJ9D6KmhxPEw8Y5H4kkGxA9XSF+sVVEwzHL0
raaHL/2Y7HnGfawLpEfQi9pGFpMhRDbujrbCmMRYmqB44eBg5NL86NO2xT6yAuBOLwruvv5qPnbT
q0XBFk1NfxkQ6kTlR1YIj8jDGaPTY1U8u5JXeocfGmAwVLsiIVFMtn2+DLcMF89+fzW0fVvn39uA
NlLfWzIw5cZMC/B2JEOsWzOHsHysRVq+/Yhr8gcDmnEbL4Oo5h6LqQd/+qXwT/B6Mfng71Y6zLwg
Wp/kvzO9k2xR/vcad2itkmqg2WKNR+x/L7z9rvyXfipgJ8bBflKVy5ppPyz2yssJqu4P2sheAu4L
O/brtJSbJ0ICzuxQca+6rO6F1NfsOBS7blpMEtY2OlMKG7Xte5aT1ZEWq4IvJOBLFAt3Jf4RzyXD
CzP79lmxpfFtPnsj5Mi8IO5ql/LhBxk+X2Z192lg8cNuBx1jV22N/+4n+PLTTHAtU7rkiAfZuE2t
/c+5JJBKZfBuReHwWGmPcvZi+/aRqYQ85Ekoz9qJ80TELw8QaULZ2XygunF3h9JKqou2bZ+PHKMo
22ybFkvhODPAa78wrYNEfdsZoO471I6/sIWfI3NX3n3Ckfl0AI33kRMn7DucxaZfo6qKvUK9QoVE
jFNpSO0jKK4JMZKnEt5yqiGF9WA/Mw3fUugcnoPym5qCB31oG2pUy2yzlKKYL/WcVctuNgXe88Td
qocTMmlvK62sXseUhz6l2z90TbVScPw2/hgynJ1dTBmuyhQtMuzX2beKj7H6wPmULSUXM7M2QApH
C22w3bMCMIrsfaFtaJtc+roXwb2J38T+vU5SayJn5EMSi9ovuVVDPztSTz08koZYNxJGYFpWCfER
j2BG+3RrFogDuEhQXso061hK701kjJQXZOkfhhUq9YgcvcL03lCzqYUwyzlXVFTbRQZ16ihd5hqK
Sbz0c9NjnrpkczJmt6OiS2prUqGbCmy8wll1GOvaZykiYzQerjbhFevsjiXYLC+4jaxGSnhFgHkw
gyJ2ynVg6Hb0bWhL5r64ruKu3yUyUkFlvW0Tic5ld2IkBOkUFuH4KUFV6jOCvttSmb0jmoj8u2CS
ueRdibT6t3Yr8pBL/GbKfHV3nc3GCz1VQjc2lzxQnUzhImwygNcM5z7K0UvBHetONGQzxYoUeNCn
t0ozFFSfBSHF7SyJARy9BV1cp7AB8HUwENN8mrQ9z52kSBG1O0cWwlP85rP+wqccJsK+nm79ddzV
JUJYWp1wzrPD7nh9GUZ5I4kcl9dyowwOVkap7q68OHAekNkFokkmwonkViEGdCrMT/bM/ENoWJOm
QeJ7bn8KZrK3eirWU2l43BFpUoBxQ/cva1C7ufM45y1VbdJ/UeiZkRJjGlrC1tNbGsXa3JduEpmQ
yx2U/0NUXBwKnBVbNmkVGf3P+mLsgCr5YVa0PYm7ApKrIK0+cCDwnyl74b8h/3iYJxe5zU9iXvH1
aQgCmEKuQPvKxUnLhHJoDFsRFy4UtUX81B1hWAIEDh8xE4XHxDqqLcJLe4Cea6ldgpCEl4gNhtdJ
iKOhUeRogXj9BdLGT5dT6Fn7OSgBiD3tmpSd8M6C5o6RRoMH+vtDTS3HD8X3neuI0jyWu5Vv78M/
AFgDkbCPA6tKR4MVGpoky7KOTNotetcTlxRtjfSVGAmEjVvJAIOs6cR/bz1wIJ+m9VBp92pETojN
5qYmmL7ldtH3MwSpXrCDKai7x5C/QRf6r7CkdnQxDCtFVTgs6abWFUspVryl6PzJXShOW++gHHvP
IDBrmPzmip1u9NmkqpWLA/GTmJwklcZ6WaCoH6b8vPoNK+X1ZTjpfh4bfMiUvuUljuclxSxpIwWa
2wbw2k8LBzLVUr7arht1qtguJsvxSy6HehzKaE+Brny22ijRP1haTkSJPlsJEDLIc7vd8oL/Gu8Y
e3AGPhH1BNHdMqe1Fe7N5bx4n3JaW9o2DeLznbmE1YrGut9b0VFEIGFwlfkTbyrSoYs+g7HI6I5U
LlNeGUPA4LWXuuzlmhxJlzjbkBSeTxMhhvGvJygfpdtcLJUmRGztRYDMHhDuYMFdR9j48d6mX2mZ
tr9D4FYXhQhbWp97LMpRbut8MEGIRgn6IbO/MJpO9ENpc53miepno5OiLiL0Kf6yRI3E4zcZTf+e
TJZaYSjhMv6ypr09c3O9lZdEndPpYpHU1nYJ89N5HkXsTtER7D8ojhl3rDAYxj48kJzmj7tNpbeN
JWdTA7y+8bmjgMa3sUuOuuMxzb9fx0Fpp2KTSjug2RB7x4NCMErKQBpA6eulzCQAyOzfR25EWibu
RR9cxjV3dlCpcWkE0BauxHcU5CyH81sLFqTkC0OYbC5uGboLbFDjbErr8j615iuPr/l5dAkHp7op
cSQMTE1mrXWZaUpbTYO8J1e+nGJUVs7Bqe8ZlfQ69Dxm/RLxidtO5ddyJ7fNWmbJAxT1Mveg6tD5
gbSIkq+qav+5p+VVUwJhkODbb1zalTVRVf+JfvVEVqDkahnyaMlPJ3gUBhRPGsHfNOApbgs0ZVlD
A5ruRcEH7VIjd9q1gvgRL0HrwFMP7Y9ilT1xomAS3BPn0fsM5AFYn0lM2+vxgbzcNKdUCu1MURFq
W2pH2yIo6Ft+ErCRWoN0P/XYUKNRbizGqDFY+eNQoxxOxFbhr+MhJ6v3nDx9U42zi4SVFXkUhd/Z
TsQfQfF6prqMLGhF8IF+vAgWzsaOtl961NtDsezpKsNxnLKLrM+XzTmqfGTuBBwFA1MPRBRA/Aqg
UYWkiG3+BfmaKZSk7LZ9hPgb9eDZhPO11+s99NrQx5XCs797XxuYw70sAHachNP2tqNJyeNV7Vo0
Jwldb/1MjnklYejozRRxtfE6Q0RUa3oC9P6Q3z32Ok20w+x/l/56DPnuOKYnUtxtclnqUumNKPTU
SAyFeBYwbBku2hUkaxOV7cc55/wDEVuvqo5U35V4iOfJgZm1uw3Me3M/7CLGIzJQC4bZqMtndakF
rB/cZZru2Wh+n/Q1GwtV560D8+Q1DBl+txVlL1K/cqhiF1+B5n+G1E1uxy3FAZYSSm2TTNzv+ROG
SwpmFhwPHwpSwrjMs0kjEpOCIpVNu554jkMPwKwrr0YQ/yK1j0oeLL27Nb7teL/fz4cMLnsvCnzX
4eM7Br8lUeBU4g46ScBnfYGW87VV5oPR84j6KMg4b9Aw2YaG24IxUqSLu11YjdotWn+eQNrUaeZU
XdZEOi5sNd68MvvfliowY8oKuNYQrqVWXuQjDXQirYvFcoh6XgrUCR+e20t6bbMiCE4kRIVAtyxp
sB+tCzRmF4ljTx/0LdfIi/5G+5ZemOlGNfo5eHuyVxlK+WhXLFZ8X4lnksuMa4aSauKBCbBPRsfH
6YFjogd4WXMDvPHSd4c+zdXL/6x/pYaf1vJsWBjRkGBg3EcwhC5c0gBuINJ+HpzydaI5WHPVuKbK
EJdgNPrmd7Q9NuFVhghR/V8SweQSBvzUKxUI83/pKu/qYlhLcQi4CTVX/w1zINhdrfUEZ4B7vRzL
j1TmOViXdlIrAF0XSM5eibrDZUjWLZEfKzVULBNm0T3dqtKGydqn3Ay+B5fIorF+S3Heip41a50M
6ZdcVODW65ixKRnsaHrs33KhGgHq7un0QjDTQX35wSskwSLfTeHvWhr700ZXbMclrJcRQvOD6Yf6
tfTMcHvedBRipwalQtjJWgJuyaTYlWDv6PQiqSXZI1f7WRdUn7IrcKc/uxQRWB8iyItVPzCnV3aH
gxloHx+kHpDrArYcAJSlbetvVOzXqs8ZI36WudfKbqvia/QCcrye5/uC6BGaEUUGQ7K9/vzoupO6
MVmm6Fe0pM7N3sDwsGn2HfXt0GhPqvgoevs8fnCtUG1ZPHGDM2/agjPRzkRnsWQTNGZzI7lPj+do
qvnQtBmMgm9MCht4Z+YoysgZnTV+qBZ5l+ceWcOzR+7pTE/ibmnDnetwmHqPFizzzquKkwwtHCI9
qFhIcKoot46pHLIaB2S2WxXr6hZGJ+jEQGZXrs2Yjwjy3QDJAX7hLoWmpoWhPAuNNn/RCYwmXgDy
rwMmQJrsI86QIIPWH6GwQ/jNLPcyvBgNoHBBnA5BfwDsrZ/7n1hAX/BVxC/JcxCkuGRPm9AZrolW
ES/6fhfMWAg9gK5Wg7fnVxIVIvtSQ9x4pLBMOIfSw2E9Z3uGTZwkcrDA/huv+dM2eXNklDeX4jwV
SIcOvKGS3iT8Xri38cZHAtcllb9Ish/utJDeMIJ9ewN6S3KDLn8fXBGQgSUQzZlXkY24HVkcaTuK
Kd+8vsthQOMxJPu+0ADwwJTWJTRkemhIswyKHxpICiE+IWG79vLZEShVuHdP8abJbQCtlEvabWUt
uGmkmmCCJMF7pVCYuE4F2HPmPUCVacF6C2pYFhEN7RsmO6hkbgEBmPZATl+P/I1e/FT6NcOe0/gT
AnJNZ+jgO/qhi57m5SyXosfi0vYVUnZvV+1FmPg5I4F+SUTWd17RfGpVHc6VZqmwcax4/Pr5BoNT
Zwn3T8wWFKs6xWFRXoLsKxLPpvbXHSP0/nfsyRE1vKGzoja8Tz+pQheghXGksuEBAhZIkj7w5JQN
wZtmCHTcjar2Fg3iW2rqqdBHG1Y9ZdFyA+4WDRD5jQhiDm7yK0+5WmuV+XiAjvZNUgRxRNQY5L49
U3zag+vV4vTceq+Qt0mxvSuog1JfvNd/T3V6MTux6pbnlAS6M/sCEFuuD3qMBnJ01qICyQGbpGpo
SdErYElTzeZvXIAtQQ2MinnBXy1j2kHUfDwhWS08D+KxWsLoyhpsMHJmSuEu7Cj1p3dbP2MkKBZb
CBnAUc9/qBKFKZesgbbJ3SEq3dDK/H51X3eytAVDGoRHnPFVvfpLVJNBu7h+tVQCSxN0JCu0g4EE
9rvzUlA015Oh50EodFS4qMaioiJb9Wz4Am5HfGWWaWdcqjnduizJC/MFZ/kfKppy/MNCguf5fA7q
gukboBrm/+nITKo6+06sDhVy0Bc0ZQoTR1bzVhnojqBJArlrdC5s3LItfnm3piwxChrjSEbDq/S7
0UcDV7WVXdlFh3cbQCUA0lg9lg4Eok1qN6LusPAMt+VmiNtLVAf1yocSygK8toDbKAiiuOTnnVta
SXAZFd9M4GtMtULI5PITDaDp3JhxfPgNwfJ6iAcoW0XweehtAO51XsJe1ErLQA/KDe7RkUeFSbzq
1KdPhOFom9235Y9B2sz+HA7x4Wx4wurcpHn0ElrqJPAk4qENI5OZnuVdtMxSsJmEs7munBaZtrbn
TAd3rlNDT9pOpL1517Wz54FVBWSbYzEvD5qtNFoWtdqs/P36BdvZ+ECjekwmX8A7/XEVPFlGVM0K
CPKcFgnxNVOFpxJ8CySvi1MCuws4TBsCEZQiAW5DGzVpEJ42UHvGBaEkIHi01mfDZmPVJNKBKCUy
gdRw5u15g1RU+akIktkqkjS1s1TnJVk2W/DbvRlB2dBkzmnY/CK2eZdTamQJjziVIZMOFlNmsQRb
iWTqr6fD9s3e0oe+dL9NSZftKo1VnXQu5o/s7041ddOSTZRI7HJzkea3J18pmgU9cHQc4b+bci/7
4vW6Ozz2rtmX9JAE57s0J6gfX1cvBPv78K7ufPvAaj5b3ey/hP2SZEgt4VmnTgLL8PxU6KXdb7C4
gpUgFaC2XercYmD7C676+paqaBJFDeShlbEhXeTUMxX4d9bmAPcXVezFVxR1weEQsUQ2o19MmnNq
WjnjiNpnviyhEd2Vs4v08a63Ukt6iIC8VhtMsFTUMd1z1vWUVFwh0u/uPQzyo9xEMdbMtXMn+hcu
EJJwm2Uqsgo1E67LrrA+w9HOPZdaxDhdoCctBpDMXITGhAThMXu3KgzUTwXVp++wSxE3LYyFhDt7
EsmhjCMFPQQ53eO2ZgMj2TVdyRLQXlJKAlCQV4ZZnmXuwfNs+YkCI5Wr+wBaZTZgGhgj1s0SN9jM
8WYQN2swcrynp0LKO76IZaUW+HqrrzMh7q7lZ66HzxqNnLFMTTolzE8Ri/6rHhhVmtvnzyb1Q/iN
NIgYntJRgUWH4tbtCJftAmHE2Fo6sYI06SD4eLQKcZD7lTLwzSPUVoxVRpDBqd4bmDZq8kyrcZ9x
ktvJvuyJDXTo6VXx68hURBp8vDP4+7svfxpk94lJLLu+0xm87PJbvuXuT5CtG7SNvtpPw/LZG9CO
ODUBtrs3fGpOED2YJarpaqUd623wQsC3LBP6VUa4vVAWj1qUH5oFJ08qTWw7sn/td/Bi7q/wtYLL
wMrmAGa4gdwyM8uZ8YLhO6HPUwURFWwt3KWYcwRcLLscVEjk75s1DlyNR3UFVjI4ybIN9c4y3fXA
TriTzVXduOniPjgc4ufUFswfH1uaG+ZDAGPC6dWdCqIBpgrmZeFw7SjEPZ/0vvby28JyDXv9N51Y
MaDl/ceCwHHmAG/2nSUJZFh4U+TfUf082MB4Q8jophNcAqPIty7u/HijVO49GsIXgRamY79qJz0t
bo0kXPe4/vIPAxbIWdACSaK06pkeVbiPDeaWdxXYV9fBLC511EJZ1ZOFB281HuEODWhxBjxbc6p9
1Xt39Zrm6EkNcPHZvmpQxrWnQiT3Nvdz76MgseHkcIBAf//d5nnyC+f/u+LOcEjfmNGC04apljM0
v9poJ4jqvL4x9AO9/Ev1RdkY65LwnfSeZykcee0bRymB37zHY74IE3fa8plbrFi+lJOTklKYARxe
5NxnEi64OcnuylGq68Mwuqe2+l0HlU/lRcXtqJSxj3xAqPSsFKcQ3c27G5BwtXTzFCfk7ZVb6Nup
KXIdX7dsYyx/MDfDFzI7ZIA4BPsKpxa4ukSMbD4C3+w0lAIvTUEXQtSI28Pyi4QLkVBWI+QulRMU
vaTX4LkmxnUjVBUNTvyhikedkF7FBZ7fyx0m2oy3wNumXGTdRvO1gLRFSHprF/1LVy6AkAROtykN
ZOjCYWnYx5ltXYcSOA6cF4aoo3PCfn+Wrom3Gks35k50RA5tfeTXFD9WpRVXknU+uU43qLDGNZxI
kGeuCn4XsaLtS+k+8e/KbJGlEPyDOVxtr0qC7Hk8PwRCuRFtqeS9BvPeBw/Gc8Lw60qBA50eZpID
b8MwF9oQLEHfwHf5sl9U8WVT92PG+v+6TE/5/QnFCBZB4hUM3wgcKWXJA0hpgtCpfpN4GHyRBfRf
i90XBOyLdb6FC5TYJHnQpMSj06BogK7jpX1uG6GyVYmrBt4h+0B59Fj1oVs02XXTV4Ni/1kSZ4Ag
gPnrls0xledg3eWQ6ncAn7jOFLpmPP04jFgnB2jmaFQ45PJpcFinbHM9unWF3olFgAM1TzWh/vrp
UphMCl4HoTg57WIrQpAWm24FR1LaX3f2EjuY+wUJPiTU0d052PM9I/DdlGVB7lJfkM8IMthG6gvp
3tKkas7+899IlsuepWevfw33RZ3wkFRnJHulc6+/xSPaa7y57JmtbkeULhgUiu6VSXT0FFtQClMA
9Chxicm/+cHZ0p71nU99rX2K5uBrrNHIacwEckkgG2xk2GXTep/qZxsNG2Mvf9xbr9uTmJwdCdl9
h0GensJVRCsc3TdVykP7fesqKWu5zOblcwh34A5m3uXyH7ikEZ/09Zf+RyD8RPAYOMXGX2CKqplW
Wp6zt4KQVvDMSQ5aemVLtvAMHDuMBOaFB+oGwB88FU7qHq/QaeG8ybsPt1q2n39lt8yfnOMgj4Or
moeGCaLMl4+a3KiseJrmKYurF2w6kSN5nbjSSi6Y/auDyqhuGUzpBDmZs01+MsxmfgMeeD2ngVuZ
qdBsaeuRCYCv4+KYJJv7sSOATQPv7wGcCVlGxu6gRS1142TYZGSCt7UCJkG+iPFWGWFPn8+4AnX/
DixZGRiJ5aPIxBMJvmH/4zXjNHjSEpbyBlQf0nEDbXzAAhjT8OlJwUR6R8D0D3Vp0JU3iA0sbVU9
HVF0jH48v3S6/5oFWe9fP3q4dvODxeJLG5tLWvpuBkHDU7koOuWlSxINghKAUqLSb2E3Mfynzhfn
uDuoB9zqree5GMelNiiDGgPzvRIRnAGHDsTah3UVRvUKkL7uRBk35NYwgnUqHhuVod1xb/vYN+5U
njTZCiW4rbq0vhLu8hydY2WscKjlxGROKuZCbrlSdNxrJNmL4VJn6dASgJySfy+Jub+Rdf0JJcH/
Lwp5xO3VjQSCYBK703VX78MO+fWjY2CjNbmUXAKGCli5kTbPIEG8HE72cwNn9LTaM6qw/NyAle6V
ukpRCRQS3/CVvKom5o2fBf7mcDrqWCjrF3dJacZaQuQlIp8Phh/y+r3a2vrL1V0Y1xdc4CyDZEAj
AndQ2hBK+AD1HSdT41Qv6CciRAbE4Et830i2lXQcHumqMmiYkZsE2X0AtDAOrU7Y8Tu0DFESX5YD
E4Dqo/s16++iZ9oT4vqS0uBQqJCgm23RLHxOTJYtJPNTNqleVp5KuviEifulzIwL9fK5tYGBpjGA
cAVMkxEHlVF8ziiuoSSQZbG/omvVg3TVnKAdWnHx4DLaE3OubUZ13EpCQUHSJXC9LYPjBuYuNsCK
FOZLsVfS80lvGEbFXPLfgLPopT/yNsx6P1RQMX+fYsLfpAxkJcdMAR9sg2pOwesOg6LHNqg4Kas8
dKENOblN87FBaQ7UvIlZv6/awue9R/m4cTG44d+3vW0W96lI1guBYz8p14C94txjtmqq8lYBeULp
ecS41pW1bKmhVlK/Jr7egZFPo4mHBDGbYerQNIAJ+qwTPgpxdq6OUkMxwTknkC0v6FPiPJf1va+T
gnySv4zuiPzRNwxppiRa2js0eg8mYs5YJBs3HzWfdL7b4RDILr8NCGxtDN8nZ1o1GEfiuSHQbmwc
lPakWuaBP6OsN0bVMNg1sELKBDZ0kqilN71Fd1n/0X9Yd9JhGUtLTz63sHVmYwdXgAvcWxwN9HkP
OQjZYX2pjLhdpY2WwfhknSXLYzK91XdPBQHQ2H1NNDZ1LIvWQhv4zfbDmj/PrW2s6Shhc2ulqitS
gUKzbuYbVoyUU3ojSq4UFZgZ1AWz8ItG1wpOEIHOtNc4rVaV0ByT2k8c3P25TYXDYy+Q8cZnJ+cK
1dxWD21D/2lBvsDKIciQ9K31DtH3UvWa6jFVIZPsOsuNrM3J2YtLYpe8wPwmo+XVgvNBTP03oBTe
ykMAWh00fC5ahYmVzquuQpwAAFUvhfL1WYQtN4/hZSuN3REF8/kk9SIku4Der0e/dp5uRgbtc3jm
h53SShX9d9dSCpCAr5J/vJ+a9cFXblH51W0aeTetZurehDcd9nAPNUe4NXJzVSupt7lf+ZU9bswg
5nV5iaHANPgbLf8mbB4+ZFuMmvZKzR5Qv2I4NTu3EXTBz6h2lFijZFMVDK2lDpifQND1xnZVqU/I
r7CIAZkODJlsFmEMreUHGzbKz3Fm2SHoID7iXUnJXE2RyIh/DNHFurqWCHdl4aYSpKVol7V4nTSw
R9FuRG0by2BdCJ1Kwbd5Phj+tnAH4J5tv/m8FjEU/GeCrEJNPFMkYK5DP4Ak6L5kWf2ePGQp/Gl/
fx6N9zh6KH9CAUT5pdO5ZeFthx9+lm+jvMTERLKSsoy5dlPHdmd2O4Bx5idUQSI2x+GR8ZQJ8kzd
Nj/2yhN4CP7S/lZhLd2Nko2kcy3cl16IZ6AywzsIp/gxVMuYFEjU6OVzwsW8r9t9r4OFqBbV2/Ly
uVsH5NOAgALGaPvBcoYDqZaCNno6Ze+jpb3KCJxqvWv26TROBXmu5JSYwvnJMnWCZ0kRK5n8Rg3L
D7Xl+8UWwMLvca2czjGUfuhb9dS+Gx4dK5tDvOcD0SXsiPZqV9+owXX0vF6IOP6yffqcaiqyuglJ
UdaoCoyPtCG7aOdz+XmaG4feCAlkpWw6kEUKqaI2ue9POm2P2e7U/oP0Z9B/MmAq5NGHpUz8o8Q/
J3swZKxwTQY8ap5OhN/RTUdnn0kl6MTg1zfGyPg1H7n6edGRo+VKl5rtw26FfebqHl7ErwlPxlXN
bHh3obwRYcuxPVvFBqv4fh4d8azStrvGmttsZdciRsEqWWrzHhRYEGPyHgloXinXG0invtnL0Zfz
SL+JYOefDE14fLIUAVr5bI/fUoeCTn37SeI3pdcwcqzQq77zAcInhw+n1F81gdk9wJuvcsFZON/p
6BIUNRJOXPt+0paudaPbcnaFDPnNIALPoUqMHmY7S5aszlJuN7L6t9xC2Zl8umv9V4lU4leBzXXr
/q83tKwNa4Sp6RvebJGB/cI2RYOdFcUPn5co3v/crb40sIzbeCVFPKzM9pO503K1DP3C5gr5D2IM
nTyomuIwLx0RkO7L1mH3U568Xoda9ujs2uaDKiQ0i3WVrEMB96n8a8WfODADJYLquOTrkNL/zEii
2WGYDc2IQKcbukFZtMGjoPQJDrLWNz7FVr3nFk8EqNg9weoeGVvIXmzETdJaJxVwqwCVmDqMNPmQ
dgDS8WpUISubfXUBgfeP8nr8P+hEsYGTaGhwz6fBN6DFXkcKsNL85JVXdpAz5qeKvlWN/ovmXJsi
LYUDvVaqnr41uyKcTW5XNOtBuPe5d+FLDwCs2V5uUyjxQWF4LNH9FM2ZKhQQU9Di5GkdotDZebf7
kFY2SBgLr/X3TZc99Uv15qyqfzuXytbGLmcp1g4pbIZgd4jpDxjizIGRH0WLiWM/49bgozkz1Ns7
DQ+OTVWVvifJoiJwH7on5Q0FqxgxafG5Hn9zOgmloQlmPtfQv0IzBZb3+AOOQchS0Vnk9V5Rknsr
0vOxTfTpHGXWfvkxL3A/gOsrP/skUxwm2J1NZWjzto/hCwUNTXU2JBGtMhsQGlQtUntQmsdMZUHd
k1/hhuAJC+m3HOwsSIw2u4gsNX1wUDrEv4UDMZB16Q0Vfos4qAGQct3rC5jNKZZuqhWUu/1JKN62
UVHk41OSugaxtkzYtQm6hgWD3Oa+YIwlFS/5Ry8fsBj6dFhWdlzwOpyHsGl/tRsIK4SfNLZQQKHf
XrhhJ6yx99V2HFu2Iafk81WkB9QmSLQQib30i636lGTqMThleCsbQqeKX0+5Ej+dkU65EkiKfg/2
TjMaeZxmMa6kneLb6YmMun4NXELDbl2jsn/327CBDkAz2fJEpNFNTX7351t5InECg9xJ/xXEnUUY
Ssu3Ow7cnvoBUgMlCtzESdbFK2espgsiOaJSwEP3oNYHnOCfySC4ULb2eHMnX4aplvEmnXk+iSFS
udT+uV4smm6rbGVu29voE91w/h7q2dxCHIm5rLrgr4x6nyPDyWWSLQwtQBiTBquuAxGArZ4OH1vs
cI0pMJsARGqbjZQO0hZt3iHbQtjjlRKETaBEYnpefD4rOalfv11asVS49aUsayvOvI4qIixDTer1
L38Yu5rKPorbTloLm8j8QMCApm9LHTU3MklNOxS3VRj5KsS2hWpEfQ5SrEVFOkQQT44KVraKMTWP
cmOCzk7bnbTrSccP+8qEcthlHoEZJXBeF8RUROLeJ2d9kllBGgOHh1EbVKxMQkxDlwhvmYu1f0gu
nm/AysjcdMC+ObgfAeeZx1L4HgdyGs954v0tNSqmqCW+fDqtgYqaqnUM8HNUSUZSqV6WdWHYpfvU
QnCKAFoFIvk1baGjMiVMTv6oIQmdYyyhKLsioPsj8LathlVl83/FeOWZox28xGHWATqovaKUDeXp
AtMSvwJP444B8075NOy2ZF/CD0xiKJz++INn6ICSPdQKAbLYLc653NoVSN3rq4VVXbh7DG89CuIk
M0cMVA9/u+hNImd7ypldoOAUm4OplG5tdhlD0+ThK3srw6ieLj8q0/HSMCXphXyIQ3nr/dWq/Bpi
JJNxEv4K4sxth21vmZmZ2ArnwuTDEdPI7RhQgCBDsbAJE+wuK2Q9zO0N1zXcqzQBLchU3dgr4irb
1h1Y84gfTVD0H6HQFej2Ykb71U4NoRCwEJR3cvqutPFOnoNPOiaOwkcYQop5NMrK95iUNnSZBu4J
sG3DCotS+jn6Q4CLgG0hjv/Oy1ZHGaPCpQSmx50/qn4QAF+PQ3qPTA2C4u+ExLB4vYd0m03VoJ47
JHoUmVXyTLJ98WAIBP0PyleB94KEthnHpLVfliWuolIYQiTiSHVmZEd+4UtT0FGX2uFrLBg5te2q
cl/SUzg3Oq6jsuQY2Z2xDvS6o2dTc5XsW2ZJo1URFrNJwtak2jhva6ZaJuTZmbVIxIez7xCXrQpO
2Jj0AubJzZrpvhX9jj1hAkKCdwLcWhQjG0E4OCC7KN79TTcGePVVKLuqfLe+RZVGekw0GQyotfzl
+NgyKVQw9SjMNg5FS2KGBOvJeCEbkA1Cuvg5dZOB96QfHJXkLh74Xglw83Al+losrDU7BZ7dwAvi
CL7n9DDxPYddv6jy9Wku5sEpPH/ljGVimPq0jyuyoGQkhvFiQEJilkLSXQR9ZLqINtg3Oery0Z3v
yA/EA2PAZXMQJe62m9WA8CEQMCBckxQKNztj8shHk4R1IW1MphEDtERnnigqB63S+5TgpIKyf1Es
H/kPjEdeJuAuI5H5BWb2VloYwWHVmw/2yn0EifH/KVZpMGUbdldF3bbqqXNJN0Df/mAfS2SUNhjR
eFPkaf2FgHwRJvt6aArr17ShEgn1Ozh8eYNg030qOf8N50/T4PddZsBSa66KrILtXoNdOJuoBgEq
8x4NL9SXgbXq/njekM6hM0JtlbRTqz2d8hTUAdamhk9hSfLQMTOi0DFZOp6EPrv1/Rlf2A2wZYYP
uYHESM+IzTslZzPDcJ4Wh+ElA/DwON2UTkoXTl594tU9bK/n7MDTtEj/1boMARJEwHlQ5Zn20CsM
VO6nrV9+zlnBf4k0uQtq2pO4xH5neflHlGn1l9ebC+dtNlNYFUnZsRyPi9FNR4xTg4PEhJh6tEDj
I1dH5ENMrFPOg/NJ7c2X3CLbxkELNdOV2ryKby+ooe03JVE7X60Qm0Ra9OhDBQggXjqWpcjR3sSm
789XwhIz1JW+DtLBNKyICgPYMR84DKSMmQfhsBB0/nO9Hgw3ljJHsMlYVqBy6AC1Jd22rYFR6kTi
Q6Hh+heCybmQrCNJdcLVbCfd9RlFgF4E5eblf2+f2+oovGlqxzVh99REnE6bjcklsB98S6vFsNhz
bkaGzL1F04HJpqRp/e+n+p46DpX0QYbAStrww3shosQb1d6igTFSwgiOAX6DO+TNvwi9lIeb3qIT
0RZl44DHgnSrt/ogUow5l0SotV3JiI68xpYwIz4by34gS4XW/DxgaqAybk8lYNsv431E8sN8DZeD
J0GpIoQHAYkEcEg5Pr14xXMTjRaWwOzlYBUCJ+pMUrnbilIpoSWFWu9xkMXWJ6VIK2tzwcs/OvWq
k1ZEE6nL5CSDgIvta6vSKPkuNIp7BMBaK74jSI1rCJeOekBPuqdaj8mTRudEiybX0q7h86piQ+Ow
Sch5vy2QbanqhI0eijJo0LOvMUOnK91LhYgBCde8bxEvV8ar9w9LM43SXuW1ofAQUgGZJdjbmCj0
zsUTDLhadWuXPwpKoCdzNjXiKifA4NYi/DCupYB+vAezUKQTqkc85kWMt1K/gMDLRvd7263w1J0V
/RwxDmWnOcZdMwEyUOWUd8BzUWOzkcpx7drmCYW9xIzo0XUAloYArh8kmPU+fqUdePuqG8BCOrWz
tMQ32ZA60GVnK3akxnhH34k/nC+umlaqQEexAxk9IYBvHYzvdr6od1WL8oaqfVahQBvLXqv51y72
pyrFMVaFj9JT4lFCWBGOnDjfI6hKkW70qpHrpjk+oo6bf6eHsZ5DTmkCDZnCLsPiEKqSEaB1Q/iU
nRAhNgQ+IDEee6WuAzW/teaW4dCnt97DeniHWsYOiBfVkyER3MJ+SdQOPRf4wDhBsm09l5u33D5X
Tu/eKdCB23RrBSGGdeLv4O+uJmoK8tdRosKYsQQWRxBe6Eniy7eHQrqoEVUkrPqUC71bUNQ8eLZ/
lV7bZBoklhqWR0Ye6Waf6Vk5vpj8IEyyea/4/6hqH/WRx5gbTA4xKFvVizS14Rod3QwdyPqRvaK0
dvk19mB7V8g+lc3DGyQg00wtQVTMF3A9Tg4elbs5pyaUq6L7l/jYZdl2imcIuzgra8eFbEyZzwEt
DBr44Kr8X++ZHzLj+0TWj/suRSrAqEuT63sH2WpmOGxk8kJ0KpXjTfaSAxL/pr0wH/0voxEinC1q
kSzCEN0/5+moWXnROOYkpxKnr1iREqmlPHzrTMrGDlIWIs94S6pvi18B85QUyEqSycI/KysSTE/b
c+8oB2jOOdhy8dplGRVt5GiNHZiL8U3bx4Mreip3K9D/3OZYiZn7yclPqH65WTGxcZ1zoHIBwi+U
8DgoPZyHb2vsek2EcRfkq4uLPx+O2+B6tOg6uwirybZv761S8//26bsXrmcudDF3fnAXvF2qbSVN
O0+dnsHbJLmEuJjWvIEykm391IC/dXeLluc5Upfc67hM9BvG/XAhi70sAYzlpMZZ3BuwEFC8LmB+
8iGwRnVbjpGy4tGtrNf/KDo3B4WIBuS9s0NU4x7nAArbVREGm87+JOJU9uVd9XJGryXMWzyEJhRR
z/IiCIW6ScY2zdueitHWFyX19XyKEMoZITqWvJAEiGpMDludJKzEySqcl89DEQTKVztshaelfvkD
fkptr85uS+WDGxKkZsjOwENiEq2hsudrT+hVF+GRWX6BWGeAhcglNc0l6GpMrzusYXmGGcINpzFw
F/DhL2/tKYqSeX7UPh1dYs3vYMcAwxQcOTJBqher3y2FoHxZVbbLM2p6oS0zkgBepqfu/6BYZyyf
4GbJnTH47hit1Up02Gk37XOLYtbfVdHi4JiF03/5DlVxJEqalfSf4MGINv9pVA4DqWfFXPBbnR3W
I3GT1CorSx5+zbhje19UnF+A4ek1IsQbEjOgzJkWY/oQlWahSza2JgaBCO7xyup0/HwQZvUBdSPA
KfuEq9+0mFQxdHPhn56AUA1HoViPAruQJ7rx5Bo6GCMOhjzFquIw9xev112Ka2/Os9VanT8OIX/f
SdTg3DjmgB6wed5dN9uCOhRoHHraO64Tuin2Mcl9QwAJgk7E8MyLKb5Dvy0V4icUxUrTHXJ+TtXO
vd7ZXdrKKEUrFoEkmI1QtE0TGkMIu7mzKplEkix+s/xel5XNMetnb87IJhw09labEoWblGRu6kdO
NIUgtwLJChZAWyA7J3X7iBZh+Azf3aJrIANoBNWldZQZvs2h3lBGikgYeSWo+vt0FU8H/Uky+D0B
N3+38s2CR62AKMegkbE5wFtoFb/eUu0t8fkM+IZZZnjrgZCgYwrtCPqOsqilA/jgLPeiZrvyUo2z
1XJZuM1Cj4DnTKNhuX6qZH7kUpN1/M8J5d2Mw1UBQBckgT94eQs/TxR9w8P6sECAH3XPqaH2pDih
+f7Ohyi3Bl4mykMp2OM9c3EpPNYB8MyA01bJ0sWRVgsljmmmjSDzlWKzOYw0bPYzKsN7x1uyQbnm
0xZSrsQWxfxwrA2D0JXoCc0SYXCJmYx37oavGkIdGhrjH4s/OXumUY5+33HpO/07DcSCADDQ3yvY
G4crmzVigfxIK48G+QZd+0Z4U60KJWdHTCKygrDvzbN7KP0MsiaEVEvQRBscvJ/t+taEbLtOerph
vql4a46jnVpnwJD6ErEzBOYbzHIcJ8UPXqmcA+86y1FCp1IK+Q+AnERg9qG0SFX89SiDBEmkxFML
zCmZE9EZlfAtiXfimUawT4VOnbwTqQn34Yzytbt11FHoXKxRya0Vw+9RI3XuDCp44XbXLIT6MDYT
WpXxNjaZJEvc9XLHDTB1y9pmt+gKtsc+fBzZ7uWwYmR264p8IQar8n5blljESn7nXopcczkqsjI1
73X73P7QhTh0WIbpJxVqG7z3q/XDp3vZCxw1bQSCJuYmFsl9z5l3YLpWnrSO0Xdgn4yZqowLOIJy
m+W8bV/YUeJbh/e4bkA7gdjiqXI4N8TuRsxOGtFnsj+15CKNUNvMnIRb6fjoEJHe4tR6PothcOXp
YRuZV1uJRlaaLe9ZYfMafUo7N9ttvxpoVQa4beYZKia0raxqVVaIKCsBhAY/dhMyodkIB2SidT2y
Poo5yFcnzxumYq6yclZ63+vPN152d3yb87yYQ793UUSZM0IDuL9FV2VyNyBWntvHyzhCNc7hCRPq
81/fTp432CC1GpKBPk2KD97nUpse9z5do3T4lr6A1v0E+maLrwZYnuFRbCd0MTlbiwh4d0UxMAVv
ipiYWvYkdlWNTRRz7AaVKUp+AUINFkcrsIRQUDeE6e76ONTk4sZAeUF2vIKjVmwJ0+rJV61KnDeD
cDyTx8GvRv8lIaxy3aoj974Hw0RgCVXTJCq2gHQulX0ASvPGtND4GMAwR14Kmk3kXKZYvOzw3O9X
EubDM6szjii0dk47R4sawbdxtrvVBnOwmzL1cO4kSKqet4g8jHxku9daIazIStfTu9vTQKyySzxS
sJ8raoTJ7VXmn7DzNcRgB/eH2uvXWmKtKGsK/Q1dRbvnN9Gf9lrYCx3n8xjkYgsTByOQtVrpmuU0
PHFYe0ZMG4wHTnzT/YAn09L3/Vukz92Xn3zaQHpHbzIo9ivWUUXG245awpwtkzRw7BFz1aIL4eYw
pB9SHwoLknymW5sbZsznmgIjuSqJ68XDkjasPI2+cVUFCuxb3LhVp/qvPrPA5e6qaAkFpR4JcK/B
zC6TBskfub02BZYB7ZOjIm2PhJ05D5ql9zalHpFkodMy8PRKUwZbXsctJm29VotIlklu2jATrXBj
lbTIsZhhnRF+I8uO3vEjC5a3w3X5+DzknqliNnqkys4ePta/N6c5XaoHS/KH0caT90pP3Jmnjq6K
R4F7a3oSj+4nlBduiSRcZBWYLR2YUXpk6ttexlC/gxm78WOzmck51EW2cP/cGlKZYqXtg2fAzPua
AK8smUF8s31/JuPUzKOa4i+8aRKbLbpvPLlblRPOxjaWu2Sxbh0VIpC4OLZhSZl6Dae1h0Jqt7dZ
zP/CdLNUQP16GFbNioAKSraG7OE+3FFs+uwFVwrzTJWpGZ2nVx8QbtRTS5F/MqLdt5a68Ip0lqdm
pEj7Sqr/s0e0BlAXc+n9E0NQSMeQmUKQLjpvTNQrc9tKUHutg+Bkyj4TkgMuOgnKCWfNVH3pxC3a
hujQTg2rPR23OjeC1WXAjR8i6YQlNiMywLa17HUcEnEkljKE8gy1l57+pPrFo2OZ7EuLGp9YhCdo
Nh0x+4mbSIqbaMa27TR9cqTGZfj8ydAFeFSJD83yzCgdcGXi+D3azoufEt+cQDBy858yx6lagozB
wYAGoX5qwg7zGf0hYi3o6tbjGtNCcR+ZKYJxKK5J0CGN2Cmbc3jOVLe/3fakA/znZmuTJfDWxxKL
hH+o4s5YEdRu1bj+O4LPrQb586WqPU4YHksYuFcjoh/ZkvAEfsUVJxygk09zDz0CBItWwTUsuIIL
PpYkXwD7Zre9cs3YEc+9z41YgQZ4LGj3jZPaGQoEseMKDQG2BpMMWwBU4eeC22OkSK2tGM8MKbqx
XJc0WdazVZMbwmvs1Z//dqO+88EYxm4y2gd5QU06WxA3jt7ryuyrNO1jVeBQKx6juR2uLXnNzouz
dhAXtGCt/dlnNHOOc0OJqAK8zHo/XsulGeCEckGdqiMrFTnmdVcB4DXwyWwNY4sNf38GCDnyhSuA
s1NGGT1MINLySSsPFDBIlRAtUpB+dB9dEkiq8axCFSBMe0ZCj77bOC9BErfvQGTVXavvJasCooqu
TmD8zENid0v3/AfYoC9EvIELbTQi2uAB1jLreKkK+MEqcVXlb4XxhAWiGoyP49Rx/t0LvGHcAfiP
y9Ma/GS7duTC+mf8lJx63jjcnelrI0znLR1oqxsHGd/bvrz0bidYHhTfEJxgpfBE41WhdjhbSzUd
HmQadZKWeAVLLnLQMYmi5jNRdPAaL+6K2Kc/rqBT8XiRuNr+wWzEXLzoWFQW1UEpYQMw2UHUwIro
2SSpWrd7BIZ+l/APTy/t1M+HJ+VddamO+o9ok3iy0emqmELYIYe7JV5XhRc3lQWYPpcgvA6kFq/j
pack+qQw2jb3yrVhrVPU3/9I1eOTFetTFZwrtGnfHK6EdgwU+JDKBYuaZhmr3syPTHuFfHJSVlQ/
YEF3ISD04rgPAG/tsazdGaiAKBVwRrBG/d+3lep5YkF9o0tRWL5v1pgle4a4Q1Oo8mqGw40Jf3D8
TSlZhg20GAKDGu9peXoeUBsvnwd9UDP3wx/F86eCF2Gv42u+Le9qaNI7Ajd48XjvR1WOESsvCOys
odOGsUaO/UMbaRJJGnqhW7Qx15ZsTbEQ6gwsUum7jvp5IunnWHkVXeFnJL5xKs3VmQR+dwshkEKT
I3JI1m016nVTjYDAs9fTRcgthS41Jj3x9wMge51wJ2lYfZtO+ufvJSDHDQPeBXAtUSa4FkyseEKe
ZOAsXyCQ0ZNnzl79sWLQDKyrg6OqnmFCsIDrEKNfT2uJps6ZjJ7aDbYKOQ7gbeWuCRh1nDI+h6Xu
Elx4Lf6lDzy5bJFqRv/KYmItfaNgS4eEa3SA8thxHAFrZyr9BS+E5/jCGtnCGP0ERaEmMKXoXPSo
XU4HoYQpApHErFmzQloB+cz0uySuxUzweohjxyu0FCUQE2EUDX3GPL9GVuGxhxzpm5IsWf7ooGhn
jARchHv/NB8fuoXBDHK34XBYOcUYUL+jkLXdbJ6QHDqzVj/jFkQAiiadnNEwlpsLu3S8Zd064j5r
njcXNdwynRA+eBg+1G8aqmX1lnwS8xjFBvffZqGIcE8d/0scUe3hqLRki5AQ29Dhrc7ikNrMZ8iy
eM34TamX4YORMPhCh6ztqv5TsFcQXcrspPSTMV6c8lEcM4fBYYrsJvY2UJM3KLfWKs2aiY2Zm/iB
HgD+0CmxuqSHSePKyzKJ0B7+aloZgwrxKVbnHvtSfvPHKhNKti8+WA2PXRIBGWNZhIvhvedjVW2s
ZpGjak6tPzLCHSOFJ/HXUEtQeylSRaSc/bZDemBEbZ3OGd6zRCEj1jL7tF8dr2asYz/DH0Dt+Z12
b53aMJopLqCPzO7N6bgSwW058Vos+MRUVw7pwKyTwMyMJ/ykp2cEogQgiz0kVdme8t4IXWfwojtY
8Z7CgnxFb9/aKkCt4mi7xmOZHSK0jOgmPrN6Uo3h5AQoV8CzcoZjrGtmH7EwcAxuaMwFdoiJ4Fn4
SvGqfPeLUJmodry6Z2ElH8NtIHzZGg4hNvGrubd7g1PCLrCHgaqLgjpvinB6W/xUKa91fG9vDYDm
yEEbkOuGwzKHarg0SFwJSrf4a+vftNmSrK+w0//ITlxU718I0mS4xaDBoPeB1ehl099CfSdFWhbB
XnBtB0yIiUyuaBHdggBfiU9DV2UA1Gyah8DNZp1w+h4FyaDIWZug1m4HW/icDigRsQg/64NcLfZY
cDEDQSe/wTktCpzTC83pzBeYUVC7uc60M/LP6tLje9tnciQUyH+BlKps4/2dbaqzXeOG7Df3ZyL8
szwTVf1SJLZAJqOEoLs4Tiy/wIZcv5i20IiuBiHMpstr5LVd37Hx7aZTulyABCQqvgfGmzQtFAyD
0v+LbOYlA+JUZIrir7LwlMMePCNbWBCVAR7yhGLf3vxjWF7FGYb5ZNkdpYXfZc0I1k6eyMXuUJI1
pzaK0SoBLEmRWw4AHIsff1qcya9cphXvDXQjMDJIiDkIPeU+Ob5bVWxsDPhRfwhXMuWUE7CnK65G
GrDu2TwyQtpUzu1YUXv+mleiO5GCDFuPiWlFejBFgExqv/HsmquezBTLV+KIgtrlMX8xAa11COBB
k/zI0NwKw3KsOwfIVaEOKr3U8X493u+Pxzu9bLUIZ+KiwGTWuks/V6fX+mLhmkRTa+hUdtBxLKir
OYXx+O14cJkTgUYfDprT/B4azWYESBAjvBYw8O+V2+/a4nwhCJTPM3Fq4QZdmquNAi+gwToQPMYc
ssPjPinYbuOq9uI3YkwIc7Ky/vnnctpkI6JcqdD1cWOXmgLMFxAWRj+gbcOlDhPTh3oQf7m2SU//
kjERFN6iB6c8bGxX5whc3QrKWfH+FBTemsbtXiAcpz7JCLrl7idOpuUPo+KBBIzFNRr7OzLIRjpD
LWJVC40BDHkVEzESebvR8i02vFGyoDk9V0evM3rc7QAtLllsC6ddaf99EDhcevDQI4Fp/+pegM1p
42AsgAqShz/PlKuwrpWlpneqtLR1zrD5jgxUlqfgpD40p76wHED1vAWQmZ1gJgEV9Smhqad0rq1d
HmTTI3Xejmnozup4E8kJz2fiD7TeOVEQG/f4TB+TOa4ud+4Psh/6glLm1RLJI01ScT3EejQJpAY+
swdVCdsNxwcqFN8xfh8AizWgTge/j/oacSRNLl1+LF4ZClKaNbDm3wJf8sn08wzchzX/ArDi5ps+
V98lUzfofgiy+FP8eYqKaq6Xv7ob7DoXXuCKN5hHpMeB7LjSxufU6dR0Fa/Vs1Pf21SUGvLRBuft
DFAKJ3+f5r9qo9I6Df3aPyqeBCpxS6OD4Ar41DKtFqyuiHVgM02/HQnHFMv+mJUfORhtGbiVqUEg
e0lfCADvKSpYTKGcd4slFBgbSy3/4xFfSZrbTGQQQyyV/GUFVXZwYM3LvC3i3wHvUaogrMeHdDeb
hyNsifxDQhxuoW1tU44alPDV5GO52HupKf0aBjUseMUGfKVNUmEQJQF3D+E8gyfl7WjW0408foZi
4It/jleRIoKcmT20jP69cqDmAAXx8+mNLdYPLo7eFJbNi2xFQI0/6510fYOkLtr/1HkoG4z/3wcg
mtbOWiIXkgV4rhMSW5lfV+FKl5Me7atev9I1wEMJ1ClYU0g1iwlUjcLbudeFyqaI3nxlzxmbcGSx
vRs88Es8tizXP1j2qxwFsFxv02qh/u+6TkL7xfnJxWjykqFzsGwpAEIK1gflvxMroYoGSPt9xcDT
5L006NgudgIU7MpW53sB8SbCsZnBTSeTzslubziyZR/a5LLjXk0sotT5QllJ+Lw/BFi7dXl9fzPv
aFUPn9zKoEpf0gMZtKmf8evFRLlsUfpMfHhqIwlb69p5NVJsxyV4D7C3j3kFHVElGlJu30JG3kc5
UeOZeToQOAwEQBagoPPbcFFw8y9hFcvC+cD+hs2kl1i3WQFleL4K4auUWTUvn+lSYnOUTAzx+bus
02ODMyPOjHUbDUX1GOFBYeoDEmYLy7y1R3PvnJedG+RL/UwE6GfNMAjEIJYoTvlOrPwtCEphs9DL
Wi82Ncy9CXvSQFsZNLRl0BckDVPVPilIknuP5YdtnL+J1wy5odyKPSTOxFRI1LL2P7LQh0tuXuNe
J1geIoc3IVzQQGqowxJa7k4HYonbJqumHFKdOw8zj3Ef+BkL0AwmOI8ysAGgOy+Uc0Yzj73XjLX/
U3ErExaszzcHFFM0gpmy2jGTIEsK3VdaPq2NN8r3Y+xu/8annDERx9hg7JYveujmbgTnDQw4ncbX
KryBJ3t/pmJwBq3b9LXodjyyjQdrDZZsJe5JgRvbkjwliYdlHlnCtqVGNuAR+JcWK3a6Bq4Ff6Nn
MCvGrB/QtqGjBiXzdgEucFIV2n4ofbjPzgvlSmCT77jC0chpXbyZDneQ6WOz6cQDOkW0NYOcFzHT
x4cR9ZqtLzyqXoOgsAhBeUjU6hxOsmkDrG73Mkz3xB2AHm3A3u8bZSzATZnUAWEyqTATZJ5q66pI
90gIFJsd9c1+BvjHqRy9rbiiNJ0/pRXFXCbxdCV9WMoeFySvRy7qWkR4KX/QnkBgdVHOmwZO0TfG
lWyV58PCn3OaCaxY35M4aRzxpb8P9IMsMW70oAefwjOuHPhI44wcuBBnuNh0mOG0PD8WHKNawja4
zChOwBfhwxtO2I3nrk5NiJjEVmqB1xUq7sQ6zvnuofZ6ochNNpyPRYT4WkFYRxMTKpNAIpfvtK4C
/nk1hOe1rpt7Unxi/bn8YoJKNKVbmL9WJ0BbwgEbcmR+75dwfgUFly2N+Zc7heXftIOaP59PEQOr
4wIs5/wuNpPTwkEDNTl+qf7WmPuypivBaFfw7kpzbXinps105xBBj1ZE+LJIpsBLjr/0Z8S9hD2d
yf9xCc9gAH9xUgX6g9fkW7NwHWyLFILojFXlhbUyjaym3vWp/GCuFe/Wrtw2EcpHNraQ0EDviS7w
5AQowpCJFqWPbXPiajW1D1GQpVL2F/SSNbu08QCRS2Ip4TokXihsPYqTXnMzYTrrTZ4v7HCtPjFP
hRdm5uRN+Pc135OB30WCW6DtoSPmWarzjAphTrSwjEfc9OtHdnbfdKymKPBby2gxWdc37dPnLBff
x7PvHw+HDUht5zupsa1IgI7PXzjHL1EgTO2ArlUIdq6sA1R/XGnTxtwIB4Tvz/amr+kBlDoZ6GKB
XILom62Q7kyrQWmLhneIvp0WZqxK2J1U2MVSi8CJ1Sc5LkrbPWzRgYlzVzinAMqlcgRtjyaUmyN2
rocxNAYmiAEfRXMWjnuGhbA6iJNSVb0AYn+/I3Q0juNz+YwWPM2MyzXUAAnLUEB/o2emzyvLVrcf
Dba9Zng7i/skfiautmDuIbzy1NIiAMKSShgIu1gsmk3I6LUa9TkkZzb6tKANALfoboQ2mqsoad83
p3nUwCliA2aW8bD7/iKZ3BdjWLnRS1Wevubr6WpVXLIlmIqOWCOoni10/mwQD5eN12FO5dc7UQ6R
Z/JQgxB54agS2Olbg/vsr6xmrQ5cuWLE5MLPUk6PF6/H2oOe9NKzVITrFWvHdgrhWrmpJaQariHG
PrUhH3innwSKgR+1c7F+svZK+dKantebkTpFoG9tsy2bDC94bLBUiWjxMY9RoXYmBjoVqix5u8T0
WzOFLDOpBB6qaRuYnkNvw96UQ+m3WikqDPZPCBatmvxhA3km54pLojv3AcvO9qACrSno+o747Zb+
l50tjIfr/PSyz5v41ZtVE+WE8l9rWHG0Dna161HiR4CITQLSMveJ0d3IQlqEywpsjQQzTTuzpdpO
X8TwCZNSGvlVaeMV8yoD3MFG0vABw/CxpNppmMfTV+8fWHbIEfEZL6tV+QlN+ykuQt+cbCRGdabX
O8j30wdV6aXcQoysrrfL938VyEPN1Ob2FcaLZqZe9Muq3N7kZ1ZF5n89WoSS25jdqxLbSB8AICtY
tuXtanASwZ3sELhUTjBAHd3SeuIas+YWDH3ItcYVtUIQsjO+XwBy1/YJ9Rcluzgy+/DwtCJ+WEk/
I7IYKQxYxHQto/0PXrc7qGN7zB4y24yUvPWqzV0hFG7tASeFVj03Xm6GT3nj4RDtyVGoZj5JXN7K
XIw8GCyEk8DHIXfgUI4EGg27GwksVkcuUm6C41DfQceZrfdFPUv2jfpIyF7yaWLnfYrUy84RzXu7
ynMgVEnKdPwyq+7Ab32kgpAss+uDT9DR7Tr7LdzJpXtx1g4bWbZ56k7dopOeA6BB+ujx2YKx9oBc
hkQrQScUVtAbPMDjUC8bvKZOIO3qBzpCI4LHR/uJJDZtkBh0DcL+bewx7CGmgbWEXU7dkc2gLLjk
dVVkRvZNqUSPxgWL3OFKVjAbJCxn7jMIvTJi8VB3GG2hBXSSTAO3KxFIJEpCmjBAxLsXvQpev5VH
9v/jb5wcAyzySv/cn+6dUs/KAUtovTQtVJU4Wf+yGgZbkS4KNV1f3nxuLQffYHBtRRF9jdZOY9uB
gKbG/80RF5ShmUgTVupyy+Mehq65SsHNbrlBIRZLRZr+g8jKKb7q0GtDP3gf9RynAvPQFsiwnui5
97iH0Q15EL4J7v4QxQEvtiE7ObNkL2rPnTzgIRwWmEtgTnMSSRDHPSQgTtAsIb86FIpZ41QU/7dR
kXTlmEl8glTPyBmDhcr+AlNqxyU0XNfRphavl6o4Lnmh+Ku/rkMFEd94Bvy8kpJNx7/bFFHUy3t1
C/eDw0Gpcb4GgrIL3k83paWB8tHOyFQp/b0bIr043CLlteIyoTX38O82YhRJpPWzE+HNs1P1SHk6
24n5gmm8oDnWo5etMA+O4LAezGHrSLlDQ8pEWo6GHMZYqoEe+SMb61gpYzdfhmckNkF1XzIhWg1M
oedxBR0L43yuA0/rVL+KSISIFokyPkg/OWoUzvXmkc+sNxw4iuhI5neZ4Z2C8tZ2KCTvwD6p/FOv
y299Q/yZj6fiN82QsiHe+X2uQ14HniTaePCgGytuBSBFz+MU8TvpaQ7Z0ebltJHmo2DEKkeWCk9M
xZ7gxrVWtzD7dIfNT+rWDDhxyRkcwMJi6vIthEaMWCTVtGgo+C0nAwpSwcmnw/slcrb/wb/j7e5Y
Z5HOeUXDiLfnYBrWkFHDXMaxIyODE/UEG9ttFDAs2O9foWsc6CwJsXI9iktcY8zgcSbBaEiW5pCC
dq7PnerikD2BDkeZ0hLySkbrpW8Hh4KUHfARRC3s9TZX2KPHTpWVNqh69Wgrskg9QKYdo7NJeMAx
2n8zpbyRqd4IKECTrg3LGljKgF5wswGULThSPmrhGFSXdXDG68353MIZFJpNvntqEvaky4LgDzpg
3XZ3l+FMfG3N5yVpq5iezYvoiIArjqkJsr6jNwMu3afX+dWuohepepXlPn5g6vFiqcrzdLmrGNJk
RzPTLA0+93z9TgTTEgxBjUiVkPfkd2lG3M06MIH7i8G2huhWLP1Io4UFQYJBNpxW6J7HdH08u9Ae
RT6vDBUmGGiH5LsqcCtwgeVj8O7u+QqoSmyPrTDh7Fpzn9FSi4DeWDygWCr1nnNIDgILCv7nXH+q
tllmaHmrIREQOvPalLQKhHVYLjVhGtvDtUSLQQxH4pA2VEEewLZPdeoqXSxOoXmFXxWNpJ9S0tqC
BHiE3UXE8wk3pM3AJWa2OXh02rR3MHBV8iSOIKiVkXMNBMC1X/D62B+VA+/ywqPVKmYSUuUf4Uex
8N2ikdCzc2auRHLtFCdQ3Tab2w4IFlb4YNuuEJvLLTM4zUzZE/CMLuemkmsaANcVes+IS5lCN6ux
sGr1UT8UQYQyfLh6a9oTNreMWYlPlh5HED8SKBp2vUB9YITL256r3TS1+L5aoeIksd2uLuQWgOgQ
2myVLGGkX7j6Aa3i7735XFdM3gzzWbSxKueowbqn1oIJ1rlYB90DhARf5W+/oJ32DE0pc74j16av
YXA9VjSOUeamDCk/f+uT2ATFRGgDDOqRtpw/a+lTNLF/lW8WsOa6TpuDXAF1qA2uhx/Y/fIofDhV
/Sq+zw+ObjgH/1RsfSbfrNeQRnvLIclgTUnhLdIN1D5KhFtjjY6aoUnxC66N0z8M0p6AUONpXbhA
gbhfvwPivntyszDgNL18scpJVEmEucL+ofsv41eugIJ7q+LF6cgtLGjfmjTqa6SjwrP2FYfPQKR7
PTYTTab0lnlxYAL8aeUfY2X8AhAplhniemXdJAL+RpeVMq5/EeIPYpEzJOI/e1lLkK4W4CG/HvZs
Ss/nPGR3/yB1OopDz7t8+XM+4HqgyeC/H37KmBMI6PSEsuXla1JIYNdxFawUzLT/LioWhYCN6a2P
aVdom+gc7vyRSpWdqVB4luddj4XuhDZAcXJ3qcJTvGDXuaIx6Oz6FjSDtbUEOBpLkC7OLFYCG7eh
R76IfFJ3np4wG/OSSZxk660RxxF9JFXENiDu42e03K+N0EOm8PeeJSksZd/lfV2ukEdNm3LjrItt
VAO1yzRs2xcWUYEAn4pW4yHsLj/yOpqwJbD9EEtxPd2mkRDoQH0lioPdPriuga5VAwr+9W+XSqM/
zczltsCL7vea3/l4tu/qL6VvLfs1z334k/Yff3HdLHLE5EWsR4urMhkYvQhCLo86dOSFjvkOm9nr
lfj0FGrbtwDMZ9DCEf2tnhJ1HEPEXfZYKIzAxi9leOsLVTeLGLf0iR73fQtzMHZhbGleGpie03O7
iwOJ11GcbZl5O+AcaEXJM/M+WwjKBZmoTE/mrxt5PEXEubKOBeJSm2sV9VysZZINTyNgNhpte4TJ
alJm0UfMu7I9e0jDscUygbnytGiU+/qUAAILYY3KcSVoo9EeXGhdYVIqPpA5zH7DfD5AEJjYQpYP
1Iu+PVdKEoK6V7AUXOw+OUGM0wuGCI+DtTKV8YnnlXyB6ivA486BKkPKMInmzG7rhkUuO4MNdsz2
8odUjloKJnLyhJzTX0zl/S59zbZSn6AW/a0+bV0el/BXfOGnhqArgfuv26b9QpeSoF0VL7KfOjBN
a2eul5XlxJOZuMFstw5EDeEB/fppZi5sEqmdq66x1FcgytZoUMRM95K5CdGGPmpRsOnXnX1vcnV3
DIiFXXjRbY8fHKG0pDW9ZPCCJ/k5qhrPNew8cQm+YfZyKUknVqA/ON8iPPcpxU6qH971FxW4jCNE
mmZ4LX6M3ea6QRKtZncZlgwehkQjvFn2neaSohnZNR7kfGVGv8nUmAQx1ljL2eVsYpjsA/P0mCkf
r7U7R799w5byqvctMcXdNHObHn0RPiyLQe2CtF2osjMP29V3Mt2OQuRmR7ixUYdmsia/pEa0P4Yg
CeoaE5h/DY4qm9wCGPudn8YNyYHR2RxfnsyONCq9OBuI0BPQbWYvwCKo5kF2Nm81hvNadNsTvusW
JwoXgV8axxAq/RRzprXyQnJtRnAFOhdH8Nq4CW0zH5G6fkC1UMaXRXoAw9H24Qi1NCzPv6AOCcRY
fcylrcSC5mFhQzsLZtSijUaEpgH75Gzq2Wv6x+v1+LTpoZTT+OaY6SzqSYneCHli8P2WsuUTtjQp
00hflSSHFxcFDKgEY3R1g9q4gesgxGwSQIIimLW/oPlu3BvGbF8jh10e/1piuvpLlKLobbxm8Rxr
pTAU1wkraHH79SVfBaYlUQOgzQW0crtQXTHbpP5b0xypaccjPcML6ua+o9HLZnulvF2pCndrEyIE
em2SpFCP5bck/i2T1A9TcVVbIMcq4yb/W3c+mC9GZlChZ5oY3jDLPsYOVCtwcx7PHtNJp+fBEpQb
FILMuCWNJv2LLOXde6BYyy2nGSaQIe8IvgQDVBQCBEuI12rXirWsqYFAmtBjLqCtL4BOxs9/iOuj
rXxsuQhzuh6r3W/nH2tGRaP0DT2lmXKWo9GqvehuDvks/VLEyT9+1CZXHgzqhjJZ+/XYAGgdhiDC
5AZfp+lpG7Lry3tC522NcWZFd2DQDjkpUJNpQHfub4fWXyI0XDuQVf6loBeeM+EmhfiZOK539Iyc
FtX5q/9F8R7QPTfqIwb2ghdM1TkKYfTUsoJ3Zxenu1PhP/Hs14gt9AukfUN/PJsBEkLIBqizt4zm
lBx7hevX+kOTmlGbiNNZmVCp9dAfKBKzzM1S45sSe+Ht7fx1i2UKuKmGFqlN0sezBUVF5hmfRwgM
agraPjQbjuDJEv00PrLd/2EN0NFAoYHlBSI6h0L2A/43YAQpZj6U97uz9SvORZNSoe1DzK453AQt
Vvh10Eeb0s7310OGFucAvf4To0N3fVfuvMrOGKX7T0CmsHyB+nO9TFTsMCMhLhEoBYyeSY1HWLGW
90A+807XeoZTF0dqoJBjjyY1gDQwIh1sw2RrpZ3PqUPH62O40/hNGRrMFL6OkMtibeCeiTyhVI8O
aWN26mUPXQ8widS2yFK+Zn63jGXxazncS7wDM51KC/G9poEQBEg8WzAaUl7lsghU4RaaEf6AV4RA
8pmHZMw07PpgJlH0ZXIoPIf5FRuUsMI7vF52M20DVt2R0Z3op+riIx5pUfP5ZvqkO8xiLWpErZBK
cUXf+PQQJXOD8yXUOLc3cRikm4DdRSRnfEVY8yAa5sBnj49oO5kdn0Htj/dJ5c5Cfu+U+ezK6304
gbnQoa/K5FTSwHn6YJk7cMM/4xQ15tCbDb3gL3OYzFO/Q15aJa1NGucZlh/KhrvTOwKrQp7jqofT
pQ6q/cPBFQgF9drHrpxGQaVRCEVazZj5siRY0Cw/GtYz8L4qwDm6YbjG7fd3yX9tJ8PRPtrLD4LU
xy2xsFiTPbNf0FlauKBFz2vFeZfObrADu7/UDr3cbAjl4ewWxN6LhMGq42A62nM6ZG4G6ARcTVoK
JNGRiZOFKgbo56xGFeJ4ZLMCDiigNkHE5el82z3MzyqBj14Gzk0DhrUSPSGH2D7PzPb866arCFA1
N1u43KzaVtFOvFeSvcDYyfzY35Vkn58/CzjHRD+z2babZ2GRXLFoh8lk3kC/Xw9uWz3VykWxk4mq
XAbT/dr8rTDdBIXsYBlSb67AXNi9jOyD75smiyneY4s40sclWCNi7LANgu/17sQ3D3atQd7qeVcq
HpNWtenuBqpZRKrNLNGA2Em1M4FzxFbMVkRgPV+iNz+HqGbCh+YGW6GzmtSV+mC3oWYFnPF/zuw8
JACt18pIlLxoS9fEYd+V9wjPE24X/YPZ9fOPWp+MUDlyP/ICfNOIeLbUoFsCKuQYjh7loYlyBmdB
fxn1vp4vTrz4iQVYpnbZwi4aKkyd4K12+lTfw/o52NC7Suz1ywzQr3EZGqfKhLJ6x64chJ5PYsWa
rII33LwES7yYDpzK5VlgNptEZ9NdrTq1/Jcs++r3DPcUgFDGQjT6JN5u+yB6Csk5t+VrVwF/ZY/P
MSdZ2e+aEaLcT93dYGp29I6/a5K9Yn0bK4mopd5AE/WAZgqbJaDAzxQoicaaPPJJeAEZ/kurHOLZ
py4PwSEFd6hB8vDWIOkmatTqaPt9qL014RFJpMZpDkJM1E7Vvlx9HELvpsVSBJHHOWugtpJ66wpw
jGrxUtcPBXhxLHn1Fx/37IJbX87oQp04sMYHdjabibslaS1+iYH4LLFZo+DNVaovabBxqYM5v2Vx
h7weri6405DS9Yu7ZEsaXKZfQxL4KT5moB8U+ShX39ceGQHvE9qX9k/gxPSNqDj5QhyvWxcCGZ4e
UjoXkoaglfT5DRlDr4um06fYsJcyl/BTDhfl860WIxxVIZuOz4FuhQ1FBMErR8oLHmk2+0cUXk+1
9Ko2N4gGJVNMxP9hR7ix2cQQF0TMtePKbM5OltaKX8u2jNkV5ZdTS+ttBUegt0JUAhbZjGlHp+KL
0Kw5CnXH/G8d56kBCDPId2nRaw73nI1WtuwiZJ6bSUv1+3BtZLjTlOFq7IppSFyB6td8QVSSbEls
de0q8gMudAsARg4A22GCFLjdUY8kIRZphzUdSdWMLYp6F7jcpJVK446Jt902wYSSStIZqOxpH4Sq
iCHxALb9+hYRZtvJiKC15kHPBsRSqM7PsYGqufDNLF1S4wPildKuZn2hQQl5Y3TsLJ9FYUqNjuoK
pWoaOrZ7jHIp5tAIF+wEKogzs936qUBZXI1vaxwwSpL73HArSUxaDyCRDqZgDjb6pB3ZFuMRbRBO
BxChCBKqCHcJFyu452yQT0fuZS1oaPq+92Bf7XhuFUp4RJFLMNmJMdEewDMtIB9s9e317qG2qcLu
NqLPh2b5ddyVbBY+ALHPDEX7Q2ruYAsjrrLWNdEf7WFwF5onX9/sGJ/nM4uSHvGfChNuAqnTg7vm
o5delnzYzetKxvjpRlDXsKabhr0pZkUjMZzWAoTUWHPil2IVgnVRHEOaFQbIJ3vPTLI8UGZPY0lD
drMw8Xpb7HpAQBqqcNy5BvMVDaRMY1+WusaIUBZ0aVkQb0ZNq+IcBksH6TBKTCBMZksczpY7gUXo
EeaI6N9gXoiLWlp8Gax1Ua73di1OWp41L76xQm26AwpAN/waudpw+sBHwBkb3sEh5F0Grc9CMpOi
PquGM9kDLp853N/DebyCcN5O5Fj6AFOszhDI4ApHViYdUy4PVoPix1xBc1TJkz894DJm80AuiGEf
5AfSru+wxQKTNpMAAZbuM/yupX8+70wb+WpzHbtnFMRjkab6YZ/OOuVRzBp5qd7+t0ayCOU0EXvO
tIeKcJejB9RHPp2VffRL4mxtBPtcWukhw56KhQ/Y36t95C+whfZDI2ywVfw/bUU21WbhPh+Lihml
3wgY/zUMGKF9SNwZahHzu8OBrJl3Lq6O2CTmmZGyywMvG1euM3ppEXwt6pY5+xOh7Y3bhZTv2b6x
Id4t3LWcJ/E7HCVUT8rpr8uZXH1DFcLQQDywHIbadsySLkKPrKmIxHvwEsROraXA5fJocveV1Qxm
A2/TJmg7T5DTkJtn1TMkDybPQ8FZfy9wPDvy6JSPOQKIEoBjvnInj8bAZb0oRATnKJbjODVMEuHx
p16//RAK8lHGCddWZQ7F609iYSN9socXb6ILYItDaB6GDPZCsfvIfs2fyoB2F62XG3Fp4UKACYg/
qzUuDjAwtF++I/dDWBHjQMUHc6UQISMiHwcm57gSDdDCI6wE/sl9B/tiLkacgwjWkUqHMtT7XkW+
kmk3kLIEpeiqAvO2DfwdN908l8aIATwAOroeKnLq+oCZGRk8+Uk3tAju/uWiDLisbbmYd00S/QDz
bNt84mJ5suJyQaQCBhK1JDynregG8/uI66SX2UwQ7QKaEzRyJ7DoDJ7u3LwWOS7B2nE3uhjxV6iU
PlIW2ujkLCPCTj1GMh1s2oLwhZHVGcVOzKy/rlA+jCfm0/O2bSxhPeUi/t00y51DrBX8R0HO3YC2
OPI1fZRCW/G3QvLj7jrfAyw7Vp+Q2ix0B+zdCNh6jXp3BF4XHDlGS916yeDybr8GaSciuNtX5ccB
2IHNAbwGKGcG7GvsRuxNzoFaeAdDF0NuEYUV+xNcSBu9BsxEXkyRLIqfuAmMziRsfPF65ELn4ACV
F+wRg8Q1jYPEMBcTzmdetyhyXpV16PHuDSsYUSc8LXJgNvmde5b7ljrK4vTPz3YrohlJtO/WkaVj
9typuDQnismq7QjtaQVtP1LwedKrfTTHWwJhZ3HywQJc3j7Z1C4So4UnVqrLpXB9jqul4eAgNja9
doei/1GCWnhrVwQpM9PyYyycaL1RPAdvH5k4MVvANlzsoJIvPXK9t2trgrs34N1g5rk5cmSw2KXq
3uAaZlGAqcs9F/x2YMzPQUZSzR+7bUB1Rd1Ky2rF6fKMPsejFOmm8mPWdGepPC0YXhC/OuSmOPlB
vSG7sNYzJLItQhcf7jeA3TozAQIVuEBAnIuPhRPxExmrfflHlAt6R6gv95w6Df54yCnWrquSLq7p
3Da/zToN3nhfJ3oNFwS7h5TTO6EhsREgiSl3xCEjqIJgDXwo55EqbIhQXmLYmyEC7XamIBAmiCWz
f3+zMAD4KHV2BFmqw6GwMkxmhX6oePb/UCKUUolbhcbbLU+sUlA9yYDdwZ/X7hNK0NDGlcOX8ulf
fvrpgntW/L5wcEBVyff6Begv43Q8rNMdxaF8VbSwZNdKXPFXdRGL4KZ0fxZeMwvlObwREWv0Y+M7
1ioK+NdTH4QR5tRxe9zgxQzsY5UGdLs39jtreHrwJeymwR1RxWXwMmbjWJkW9ZdmnRkDzWCrV21k
eQGrnLcKzJvcrWosIURUQFZJdkShnLBjN5tSvYIaL6vQFMye1Owjtw==
`protect end_protected
