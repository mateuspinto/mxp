`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
Tf5aEBc3RILFaaTcafMFPU3LEL2iSUnqhKtcf8yUHcEJbUqvyLNZr9tEqVF41eZB6ykrpYUjjJ4D
Iv3U50o7C2x0/S2IFkAVJR0Xv24oCr3Vk9NzXkRdd9xBuVssQ30vjUjJ6xfTrEIxJLiL0wvHBEsf
wQfTiFdqdqhOsYEn0ye5rLopChGWMpSJ+XgZIFYckMUrRSDwBtW7Z0wGLPlM+F/9FzjhkwJJmH6M
X69uEtJ53L/IdAzVrhcNsrFHwLSEExB2MwmNjLWsCa5s8mVKcqPDVSqFzYcK59cAB3BO+dL5fl3I
nD2QCcsH6hL4sffWBkTPWtPj/tPLNZJSqzxrDg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="Ud/3CGQXzX5XReZ4vXAbbJBfZnY7CDqLhpAuBPHsVQg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17584)
`protect data_block
s0tkrMbjW7uQZniZ4yDQWy9E0VzbLSqN0z55eEY8iYq5LrO834qib1HVOGTb3xIRxhX1mqykVT/q
Ztun08dkFOP3OSRNdHEiKqX/dfZ6JpktbdxdBk0UasDxgCBCoE6QKLup/dJ+S6nOUpj6RgbaGHlz
rBzO6ukTPuFtD7vuJ3MKuLNjZZyGdx9XlCt+4N0UK0LTK4zD7/fwV3Q2cvmEFfFed7uyAg6pZnW4
4m2vVs49nM8OE9WJwl6JQikSyDw7pKEv6YpQTCJzLAoIT5xw/4hWI9wffwI2/k5ETkcQcDW3vX2s
8cCJzEwRCIwk1iZjS2gkP2mUlYhGBhbaJiFH5h2CP+VmN38JazT85skurNbP7E6QypuDnzkCo5XY
q9V7M5k30W8RG4R8g9oJm1vVseFulrWz/SCvpmAUEU5PnqR3h0q1ZI5ZpDhPVejzZ17PKk6Xx/wz
X6wzVkWtDUcQ6mvvRFUPC3FAejjWssDQs1Zn/vsmgINrrdp4vmluIOzj7h9WcVogqMc7ZF2zgS2S
QJ8rDgIvyRhEDeOLSvqk184tAdndFygPuu43s4Jnu7+ehLu+TCCVjPm2k9UIm7ANRy3WJOcr5IfN
KHQKnB0LZ9rzbfPXkmLdg5+X1Pljrm3eKWCPcibHC/7FXR/n8xjaS/KFBodpTTQn5yc2wS/8HSwE
E8S13vuAeljnuYC5WKE6kfjKz2A3hW4hk+HlCbcxQEPYARxNEPeG5JDhBMNhJ/RdObofntQIX+37
6CE17NRQUMB/SEdN7pkyd3HAzH5BOSHRZXXyFilqYlAmVXoxzu0emtxacfdwPqtQGE2Vg7VQeGkZ
Hyw/2oaJzhvVhseiH7NakV8fYZ3ZPaHIyu6b74GQw0iwjTpRbOnMhJzO0Fpd1E2gIs4zFRv7Ypyk
ZqYzQrqeXRGYn4G7D6PiaCINYeqvZ0xaLWpdG3ZsT2z0ftTZA5GAeZzcK2b4mYcEVk9KA+WghZYf
40ce03r/trobPLxhvbJkY2JkBjIs2wavNZPwrcsFLPEHNiHsgRlEbQB7PGYMsAdJoxxrolPezLJ7
JYR/qkzOsfbg3R4RgA65ViEFb/XYN1DWfc116eQ9yjYBd7IemG7Sd5+qlHs3HzoAOlt38f0oE8Ub
JtDTnTn8KSzQgs+cxYg3oL8YLuxEjbBi9fsoWSzZW7nlgqiBArIWXieLW0E9/9uxydwdjfX9eDPF
O8ngXTQZQYkT1Daqv3ZLbLYPth9jv8Mt15/EsK69CX1cakNMgyXR2IIEr0bg0xWO+jL4O4REoPhs
9MNo18LuUhllLkGI1EWSDnThYshrn4CMTXKBZHo+GznDC8QTit3VKwxNhuBwrLM3XZngkKvrBgB6
RIVg0z2kbaht1XeWnGfEoNHXBA1NwS8mUe98LGdT+z7eIszvp2MwHcazYoN0F4qr4NCovmCGuiVu
18kQ3mnGYVlOkPaK0ppqcqTkGf93r5qJazDorz9UYqknlv1eBpu2o9Cc/EfHMkSacHa6pOv+jw13
KUMZuw2voILV43hSLVpIuUqxmtnzm33ZZiqFEDKEgb6BlLwRM9r+GY2U8LkFy0ck2IVJq5U13uq9
fuEQQ+6vKmE4fsBGyFWczfZHWCqHJ/Pn60GIrgDfwh2lzVJJPsNXImn0nJtk/yamsJTkVAVGP+5D
umx5Hjv/sYslOPYlE50MqAPwc7KrHZp1jONobYL9/yJpLppo/TspP8vjq0lU0puFNbXKD9prVXpc
GBg1U2xmxWXMg1jHNwuop+LsjmMgnjRikHuoARTDPoiiXJdSsPz7saM0zOy0AR4bpbX2HAZL45vn
Tt2JGV5dpzJwiPHAdf7v5Nzb43zksZGFPnUAJovDFL94lwoRJrZ+1WDTwsyiFWY/IVRo/v6Ygv9s
E9Rrwypqqeg3gewxMWYtisbPY8asw4AVXQlv6K4EzMdamB80v47e90IdNfiiJGRK/SEM6YewTtAY
lYEnRKItI6RLccudkxL5kU80uLu6SQmq50sNnEcpF3BV0ylwPPbviONUBfWcecq6bbLF2iKHSuOR
9njhS5PmgM/qQ6GCUOcr4Prm7tZHgdKvJ5m9Jm/uM0/uAldwcBKmHppwUW4O0/bzHfVzPPJPKM/a
FewrHinH5JA/k/o6qt1PwwG5v8jRs/chv26yk2jEI8YbYI1jmZ1FP80hzPMUGhsLz9GC30ASUwxh
o5GeHEOhnKiA0cjZrldPSdaowwSFCgG1vQYnhmnz7FV/hyAUx8btEJIdUFBhO1Wc9YJEM50jdy+t
vpnvl5QjdRpWa8ZWP4HpBdp7YAHkwS0BGPs8zv2ntik8RkRXMlgYho3/8hmIuYnqLnsQseWJISKO
uKWxVDaCvYxUobDyk4/NOLoBN7b9/dDo64lY8i64ql0DKqgrwv9Y0/1gbY9rxo3d8k2o+FKY848l
GdMjPoLZ6fUWTDy3rfq0khSYFwWdxojtk97f7SXSqBs2y6omm/x0H/hPZUDx2d+x3OBlxji8NVcQ
gNSqX3zi+YobogRyX4qjlNkn33vHge289UUteFV16Kqd/+a52JknBhkCy8nvMJHG4N/Sd+jljoOt
0RvHzYu5loIjmFXT2XPzkk5zPCM1u1WXL5wMoTYvzqbOtRadPdP+1Rg8Sbo4USRZ79KlfcqFSYC5
vmMBHCS30pV+ywy8OwM0mML1Ma7RMcnhps+mPWnoYmIcWSiqr4yiibvfKYYuQXA987M2Uu3jPh/L
8jdoxn7Fi3G8SEvgwRR0nQqtkNYZRLcqmcoB+Yk9AtBxY6XzWLvKVETVerA9uBXKmquKsg7zhEYS
2hz3968K//fc+ypGTgRBsog8doVy6kdZE+ge58zee0GiY8dvE3GWtruoLXYkMdC/kmqLPxIAg1mn
YkIOts7iWkBRioMsdVnA6wonv8PpuqNrGSZKHlkHQcEAyc0q1Fokguk9SnCC5nUAfLGbR4PLwHE6
0Wh8mHaIOop+tbWMCMrO579jhD9oJjxSIP2bP6xMvbq1yXpXm/KnEJIPCuLPLrSCQ5JqEEUk31tg
TkpSfwcik/cUEQ9pwpFlwYuCBA5XOo5l6bA2uJzS5w/qiGnEzgpIqZU2SAlh6L583DgtNCzMB+lt
ARa5394kl6w49sIKlZO4lktOOGOu9w8ICTSiKSKS1sRooNQsb9v5gRxzcc/GNlNRP7PiNUAn6IcG
OaoBQ2h6inGQqECU3llKV5uNBJXYRUeQVo7Ymy0QEpSpWwD2x+uufmI+pyf8ivp1YWUjDUUaXBLA
LHBj/NR3cd1uwIlhoTN2ACz8SW+FcMHn6Z1MocQ3eJRS08ryT8yWGoNgPL4frCPr8LTd5fTV/OrC
epqlwdXF8F1YF0xOU08YAaaHijdC5GgojBVjQZtfNERe0MLqx4lNLA2jzgSPH7kvUoLH9bhsgEAy
/G4gnVzZPu8ZbxtTyH6eAPM18LZp//MfUZHrG78VQmeb1A2pV8EWYZO8d0bUfMMQiqbO9WcAcajH
Voe1POQxPKSFgrW7Gx5cwkKd8gikJzjaHvtBeJcVfblyiyG8KJ0duz6RaxR6kqESik4nAsrVv78U
1AD+BQ7xWCZTCfCavqM3N0YJXc45DHY0LC/i7/79NhxdO8Qg5eN/3bxjhwo/xlG47qqtsPHM06AA
ErH26B59N6rhnrxXSQY4SqTfe6k+TiMOuGj/5o9ceLw8+GdtCkBXaXm+jbWZV0rrmdRGm0lDAhr+
F01uru5pcbGIODnk4f0/8cTh5o2iK43O3tnZlI7JddJzhr8w+K1Z4jBuFEgR3gPlntNpc1itX6gI
TATyaLkc444CUvtaeaAfjemK1PsRdMLBAYpRnevSe62KF/eQWszntoZe9LdY9w7i+A6T7ZnvudQu
JevxidzIkhG87g11Ss6FkKtmwBJxs4QT7YA55mejrJ+6tonSr0slJ3PKpH55UyBEW41mm+gpH1/Q
kQbX+qeOi0NXW2YG10wtAS/icr9i260FMEHuJLPL6yAOeEhFycHfHjII7vrcOVPu1EBdgRmf4e6v
169hHHGAjsNTaGIkFh/JWXRsn8GaToGRxzTx1Gs8A88VIIoUevRZv4V6OWbALAL23X4V1cpL6MGn
pBUI/47rlRiviHWsyviVtjFSpKvmUjMvcCftZmnPDjlpPDPKKSUeN39e7iljzRpao/IB8iL1oC4l
87DH3DGxCE5gT5N9qUpHVVskGUnU6TU2IfMNovK3x/yDyAWVVZka4IfrsJizbt90yo+AqEW3pfr9
J6M4ciN+mixeZzEztz4tPK3hxhoXlBwjPSuwATqx54mV+Q4/1IqgUhMP+7/zvbtIlC2ZrH5IVDuh
JmkkeDJ5txWjVtCVQo5VoXPG7pad3JC1AIs8f12sYpH4uinWNJjXeLQ4aWzYUapIXFJwVk2Hs593
AZ9KdXaLE1KLPMWS7m2zoF4Qs+xBRnfqDebwI3u19T0/TS9q+sOBj5DJlIO7bKWD5LMtu5i01Ry0
ThKlQzkPMABYbyOBTdXaDXUILzYNG96wpIfs/b18JwwQ5fdbeV1FeCmCxxaWfEJipm47ompfbSvK
ay8IqVp1YTU7tzZ+/etKaZAnz0vxIvvMh3dbc6N7+FMK5Cw1N70EwcPBcCd+f7Ralg07hn8dnERG
9ygYcc6VlEv3UOZD1RRRr/1O7hChywT0mCdA0zY1FUX1GLYk4xa/81vNZJb4AKgcTLZ1a1F4E2gi
VCkvn9LOqXcBIEgcgSvJ2dJA6nfIu2LX4ay+5KPqO+EiLGh5XfeOCYLEjRMDXQYY6vXzKaxY/woe
gHTXbqO0tttLDuHJJqvMPWh8xCXFzb6TJxKf99lWMrJ3ukUufcQWO3h0SdyemAoSTpVMETaRFyQt
N16C6hL33832YOuzav1MqlEazGzmDKOfJ2Jj5nSVCHqWVjhHlw2e2FAFpZRjv14xRwcfnqUwUt7L
H7GdXGtR5Tqk186LYk3wG6FmEJb8/DBTe1aX6kF64K7u5pvS4ywusJWh7u7xnSy46jpYjiekQiso
o+pHxUJdirGmrWWm4/Eocw2zthWBwOHTapeX5Ot9EMCh8w/W7KCfDK8eoYH12VA8A3hPWRyCmqRH
K9bBnPuIwIiIBeUbAxjKzXcPDX8NALBLtEatssbwAcYT8rort+UI2GNbv34m7zRDxAYOJIomZyZK
ijyNqoU1X8pxJWZIPOinxuLOiXKdmwFQIZ4E0XoEteVS7NM1Omcfp7W73pQtIrBfhrMw4D2KDvC/
hFpsDpijfsLJd4GVIB5fGP43dmoQIYzRbBQaza3YEpcj74DGhrg9YGrluMhF41QjeqW2/8tMFEVW
I8cV4l7U9By2UsfvVpO1OTVcaJzGuPPrPME7gIcbpWS09biZ1VwFsizQAczHKApJGQgnYJ/ShnGo
B7xTHFDJBD07sUkrYuI1H79amUsZikr1GLP/4KuoafwD4MhdDudiJob2LVRdy6xskEpcSs9+JlSZ
z67jfwjXRk9oFTYUAdxvkO7XuyhcDUSuuBPa/Lq0xZ2QsHeleX4jURVP2RgVJin1+zbwvi+pmMWJ
MoaS5gclV4OEhpZZ/qTmMV/M19pHOLibN+QsS0a24gkojQfFRV4q7yA1N63D3pKkaT4RqOrcBhRT
46V5O9haZQgau0woc8PCVSYvtYCNZBk1waegkK64njr4AtMApLMygi/psurzgveFF4ErDZvR10Hp
mbt1iqe1NpFQM5hY8/DTq2ieNC2Io39Eq8Ywn0doGySCriyiOhB3XBV8I+Qi9lry+O7CRdaaeMkH
A4b7jg6F7ge2rVdSZDPQWjY1UlTXf+cZpWAT1tiN7hQ/jrFzuQN6BX+XFMtZNlHDg0x6RlNK0RNM
zpN0zhdiyNTo/W9DjkHsiL5bT1+ALKo0YaWnp462jarkubTIJrA2/Va9hFgqwFCR5JVUwqVYMjKH
jbrIIZOFxwbxTdRA0Vjn/In27GF6xZWcwhz2YvGZBmSc32FzYeAwThRCE7bPxZ2d5keSExdhx4tj
0Bj5yF6ZeDLYIqkINe+LSBCg7FHiRVBycMjVq/+stKT6qPX46ViTz0MP/rKcrYy3mV3B81OIGfcL
iy3nQjcYxe6TZLqDci0D9QHEmufvs/DOkdN+chCWEUgAti0GhljeFTDRPe5la8EwCupdMPCMYwa7
+sFwc3UU52/w6Z3bmwHLmmZq3hjBugn2jf0X0lYaZrtUmtqYtH/vF/xkdvQ63Q/bnzLb1ky2WxE7
+xWQGK/8bju/YLiXN3snl8d6fGRMtT+9EuuNM6vl1Y+mCM7GFhj51k76fH/BfhEZfG0Wy/LpTOFz
D7HWWzURY3NHsKlZPqK8ggJhuhQIqszBM0twzLEVJkPX0dqS24XNgUvDapMaTURxUPkXSrYxMfCG
BxLmHgFSFeQPtSBsX/xlK4FYeftCuQMDBPRWGw37UZHid2TvvKUPTwTGHy1q6OPZg40xuySkNSzX
bN38u44joLBy/g+ktNFkk4Mpf4ygVGIYmZZGtXkQNqdV1z3WNGzFfwlQ9wcU19OfsZL4nLsVH6Bn
5YMR6NFb5deBRv2MW0VItgW1xuY7+9eD7OhGwzsqp4dfFeUgYzHYmYSi6sxXRL/BYXppYg3yKgR3
VH42L0Bk7IRGjH5mca+tuwrmmIUh3+i7aGgej523XztAooEi4os1tPWD/UGiqHOpQCsWQlPzOiXJ
oqGouE6/5xqHzxj/3svbpV7d1/43+BVlrJdhVwZZTO5EBzGaXbFHipBwcNe/QK16dvEC5hQXOdTG
QMZ6d5fC5jO+CJy1hUnsTqcDil1a4BxOlAfUDJJ47pomyFuLTB1p0pFZGR2COpSSBdm/JG/7IMtn
/0AkbO3zBDXIjzflYKIi5f6rb2eiudSUk61rz9KGPzvP+3J08DhVB5kMxUxlcEOpxCxp5vu5bQua
6YYeTpHV4uoPzPr7p+N56Ju7rAPS+RFOlgFwhClH8IwgP6BsSYEwGncKk2ER/r6GgMtPQ/kleAwY
c/lfwz73IhDzyVK8PEvR2AX4eJSBKKhHhB/aaHjKU69ZYDV/oT2CHWC2m2fVt/dTkY3nkABKEVnB
MCmRBrX22ODtT4e936GOBsNdy2tBGCD4oXgu0LeqNiseZTetDZAUxED5h6YDCM/GX+xl5s2ADDHr
EjdKoCGAGFQAqtjlkVfn7+RLfnh5HTLjv7YtAR1fZMvYLrr5DpB6miLHgDHMZl76ykUA2erY/F/Q
6E7xRZem/6AGifB2qAvsHSwPNsrB5N0UGS4/yvJVjRnHW62afiAjM2CYQELKEsxI4SHkj64rV1qY
zylBUUZviO15WHTjMDjxZ6fY7PJ+oo/YgHVabHCdHo53gOyk7XPjh975Yli46CuF/NC58pQWr7vs
pwPcgVwBFN+rGFiFshIBS57b4aFxLQn7sU4NA3Jd9KZ24PHePBblpOd2SjReUSRtqcLB7vEDATU/
IAn4K82b3JejISlvRPchjR+eA1i0l6D1BePmFhKtP3tpOxC5EFy2N/Pdmo9FqYr7Ajt7vMyTvubb
bhon0Y+aiHgpHW6lNdTjNOxWu/sCTOqP4Wi1noVi6+0l6SeHPnWsUDWr32l44/ZRw/PjhJ6/DIaP
RMz0C4WyZbCSAv0E3cIGTK+4AUQyXRDGQpaXQYcKE3jjzTr6fjZ+dNT1Un3gEsgrHbaz8ITsYpTg
c8OTNZyW4LHeVx0RaL4DDbKq+ki8gwymHGKSEaAC2je9+zNip0ki/hdK4yiTd4LTzr8txCArrt18
PziO6zE+UFsMJ6QeDM6fxB8MSLJdo2zIlSl6Z/2Ju9Rs58u7FOA0IagDX2GxSLL22m7bEKJwk0zM
A+GzJzNNgEsyVjt+125CIAHlXlNpfZM9BM5qYVe7LEYZs93WGac2OPf/M3rpi3e11/x01h5LEXsK
rUKOjWXi7LDICxHUWbzc8vQeOtN9DYQ0KO6aW64ZWK6euuydDNL0EFW7iBCruWWAxtUF8pFEpnCU
b5vSlfi6z/PZS/eZ9H8lLbNVF8tvWIVxemPr9P3Rw2jZI8nFJQf6hFlOz4OymQw/wYy5qGLrlpIp
xEAWbwvHC9LVVctzHEW/zA/sHiVaECkd8pwiI8RF1RokMdZzj5pUWJF3N8YIOsMHnrv6lgppYkyz
2n1ZtqssSNlEW6LeJ9z1/ddnqc9SMqbe2QZi/XFlUcUa8uialS5SqLoZtNsfzsY56CGwYOFFUBwQ
35ACAYssRcQtoY+sRinWox1s2x053roMdB6iDhPydPD4jXTC16ygUWn7K0ci67YyA05hXDRqdMKO
DR/zNyUpirNhY37++bI3luYMJAHCoE7mey5huXd9rmKB73Y2mfvzB+z9cy67O/i7DPDDQZoBp2Wb
S5OqOl3B9GekisujZENVHTJSbEH9GcDbcDg2ejz+wf8Qso1Eef/6szxzN1srWeNIKrj4fcs7EHKw
30hyUM3BhmbJL2FWOLM0yx2joV8qtgtKzb1EPOnGvI79JG7KyVpZUySV+svIeFl3kt3UfhhRZWpx
eoOH2L82e1hkyr+pi2KQLayuBQaUf6Hops2j0h/V3kSrfdlsL9C4y7x5kW+J3nYwf+WfYNBy355I
h+Ol/GG1r0gRfXNhxxp/l4N2BUx9565wKSbkPBHhXIAKI5kR0QN8Aoq8EY0nIccZGezbgvlWH2A0
bA5gyvfUq3dO8S4WkimOiVlZCEWOoMfDaidevKXFpCxZ0py9d4Tbx9CjoNKTntN3iuxWtwXMW4eW
0UJLQ6Q5bJHv30m/u6yNwEkCQ5S6dCXqhElzhtmysvcJjUip3MIEXk330AVpNb+CidB6xCDw2hPB
WehZC74Zx0qmTftEKB4Ishr2fq2PLT7v/Cncggv0W0oQV480IBQQfyfyabVNR9NurEQguaAuja6r
2IwpIr8Lf/zliLj1P6RLXQR4W/QTSO+5XR5d2EnkFmVAZzsqu5uqAFYag6vzhERXm9H6/Ka20xwH
eJwxlvAKufi9GOh+R5wnijafO1y4IrEnia/fxJeOQm7YEsitQpYl3ErX2TqZ/Xda/SJvyvjWGz+S
MejY62becGg4NRIX+gJrzphhCLaTuB8lfN9XpPvWhEsyZnbel0CiYm169/IniRM0M7Q81xJJJp8J
esXOihOSQupjJxPgnP37oQ8owT2Q+DuEmtd59B9PQSr/5ktmbuFbKuxUEv5hYIZDTiVLset7SiiX
CCgDzd3chAyzZ2Z1xfH2TED7gQQAISKANrJsUqOMkUiAgqJJ/P6AIhx4dEVkdGhx/NNNQX1B8EMZ
FI9XVOnM29Fyg8H3gQbjIJvl3BxrQNPJ2/zDed/diw36s70sXVwnVDM9zyh4U9u8iDnItTocrtdD
maS8uMqbglmZfkQ4ilHLfGqRSelG19ri4RPwMUq9fqR4uFyeN3nQGLX1R/Vq6YO9lmXKh/f69yH2
zPWy2CPMyaVIzBvISAwcyoJRx7L7vw3vINMklcki5EN7tgyIJXxlXYGZcZkiOcHY1GafaYAzyBFn
Po/F4Nkh7W3oBraYf7od6iu7f5cHV5+pwBRom+kf4mwybmJSWFN9LeJI/ASHf9qqZ+LSCsvSUfH/
vFjXM5JgOi6GxUC2EkqclUwZjr7fPxu0JdonpwcRnXape/be6M0EGWplSCdS/Xf57lZJk5OqZiMP
82u7ZN2y1H1MEz5vQNtkaHBKqcQBL9lmaCXm3IDU3hC7YpW/aPcovfhcwu1FxYgV+fchckcKLY3t
iMzIin/7DIKmh9Vha8bgO5HhScIhKjH9PVklP6/cgM4bF/nllTZabJzN6epzxcIuYJfxbMjPcthy
ri+aVem1IRFUlrWUfE5jjl4qtnC7BCBPiEpV+JqERZkzH7TDXYzJyyVhqRHkSegHjDxAgB4IHcY9
Am5HOet/83BoFzumu0MiRNK7szj5V7J7mdtfn0/bXzdt5y+gFeaibJq9OE703CQQmatRkB3wudlP
PLOpLB9ifs5zB55EYItz9Jhi1tn5JCNkygD9BVTp8M9kyf6IB368sZjE1gMNDYj5VRGXaC0voxNq
w6vxe6S6NXblNww90RWabJiHRI312FgjHFMMqyUd6YXDmDtsjj3k0MBrBqNy98CjJeZNN6hmyCV2
+W4BWSvHw6nbxB7gZpIQIBmt0tzV1FIabW5AugeN3Cx6SSyPh/tVvuMG71IKGcoUTDr4NptKjjzQ
C3a7rl7a+NAlrfOpCTL/xuD748kQTN5IAAYvXmy+0uU7VJXk86PkxqB4diuEPoRENWQtJTd1g23K
0mOGRkPHXeBBvYLAYAjwxksEsUIucznlK4hQZoEDLCvHOE4KMWfaCNVv/pcQp5EH9ISfJtMjWmNt
VKrO73PITXsrZCM2X4THmiSd0RirUoLF4tgCnY0Je1+u/i9XG/jRCijtmQfSah8MSLOKHetz8gEw
chYwx4dCXX13JHp86VjQRZs+zWjo070+Q5q31tlwkk7IMFzss6+EWEm7qvmTZk7f+2UN6zUpj3l+
yohvM8EqjrHbqYymvAUutnNiRxr6bNG/aEtX52wQLUNr0d1iOv+OhuA9rvqJXRildp1g6JG2yWKv
GwO7M5AKaslShO78IKDxKC8EYiu8okFLivoI5rITzPhzzGonxwWF9E5iy7RyNL01AGHb9JpY7/Za
vpE63DYG3PfSX0V8Ht9nEH2xFyByI+I5bqt5DAKyFON8MlYb1adxzjD8DtDIUucNZhbjp1A+qTlw
DlDSXXuVhu4/dZ6DNBHOFrfm+9VrBqXme/eYop2z6CMte3JMrXu2ydT4wsI2UF3SfTs/PNfO7JYH
iTycatub6MsVIOud4uBrrsc826UfO4rkc0vABxxZD3lbbPpcskEw2Nn/y9hfZU2ppIr1LvZsEfzi
hV6vDeV+xAFlhOXyOxDCnIppXpeh1dlRdGs8JGj4xsc2ByQDJJ4l1txV1er6v52G2y4fIVc9hMTR
3z3EF0+zVROb+CBtKHgp1uK5kIFNwvy5XYcCsWS+IitKqcYLH3GajSJ7MQiofMt5IVjr91S3CvY9
5Er4e/GOJPv4vfCRnpvneyC61EHK5lg7oNA95t07t46tI9M8yCeWYbbls5uMS8djRzbwegUs5o8D
qo9aAKEYBZ4tGTe0QRbUSsjOXZ+wxuZkZvlBq5GKX9cMahKCsV6j73bLx+xcRgHJQQrlPjY1RA+l
syv6iNaTXSB2e77KbxBY7U9bGFEiQ19VZfqyvGsYEy1xznDBfAFe+sgrzCVz+/l2toimnPkGpDf/
FyPPGllg/CRbrCgDnzwol6Y3FXLYmVu1CMJ2JuwXXgsJSTJrv3lHJYqk5N3oEMs5VNCQhoSHFFL5
JJzT+JjEbhrKZE2b0ICt0Ka7yIUhdz6pbLkxiv9UudXRll3A9vClDl9Pp0llRKApkohIEZtvzD4I
aYzc+cFtybbZNtVqzIJDDo4BscC1pLcldEiWGzWVlkkldQYXPX5V9y/1nB0Iki9KeIRLtQ7bR+Ad
D+nKgOOqiyIFrSbajc0woDn5zSQrvXjXNyTXEfGhLStEgdaSZPBNPVFt33MwQOajfzSW9uuQTbBq
dGFsxBcX+8Tmjmwue/NMPX++T+CigCzUUnVqkY88x+LSZAgwNUtuSpmEJQDODoDApq8xIjltz7+v
YmdD2BbEJDZdwOU0Wf0eupyxxSffx10BF+uPyBYvhD+Fp6zTsividnF5jjxll7f55Cyrv3QsU1Qg
iVAVUYQyRy2SSiZhO/IfsaS08ERkM9KODamVoUHqh8umuZdfyFuWvdEF1NPAQk6ALv+0M/2pNEA/
ispjCvUCrQ6NtjJlUWXbkHzt3pxWQZ6wn8+jvA6/BnYwdFF+ivRFw+o4a8BVnJpV9gHjViK/dPDs
mIGeQsZG4zrg83pLbT150U2Q4rHsLnsw7pna4U/9sYqVzT4BwNRUyTfuwAvRKSzKKiZIEaKcexPo
47w1mtwJtn+x2y42q16N2OJSqn9PXtM24xzbynw9IKnhKsjShP6Tzw5s2N2KCFpIeB0Q8pyXy6n7
FLSgHKZ/mujr+7KHrffMfaiRt802LbNUh3ZnDyG0n4o/hgL47baMZ0AnPPKf9fv18b7hU5AGHoZu
ElOctngVCB2XFUjly19VevLi+U085OuYLvwBn/BCiQD5+q+8Kqo2bbNfhrPkEAr+KFZDKoS2KFdK
3dftF9rSkqEH4XS43prldkQA0X3gydURCoDkIp86mA5s8rwpxMxEe5rg6nr15ZikqbT9rc+Yeh/N
tNhJAn0rZTVNh4XSPxtGakP0PRm8p7AyePjUs336DCyC2+fSo9Ww8rEaihy9rUKV2nSa5CncZrcv
fQnuIiI2GwXQedy1SI2/BvlC+Lxnx08L7emAs75cFP4tI+S8kwT0A7P1ml37pooBdO+C/LJ0crHw
OYKPemYWQeEoiihrC65CbVMG8JtLZiUpUkcmEQzngt/5dzA+yCfwWRxpJHrxgz+PwlkEVHOZMnvR
btdrGQxG0laZnDxJRr3wl+a0VclpXY3B8dtWWpVInJUKTpZ+PcRDKuKETZtDHdOSHZsSUaW4fs1n
h10w4kHaoXY6pCrKYMtsGp8tsOCByP3jLt5r6em29i3DwS9OeiWMk6zvfLRUQRyBvF/rvq5ZHfwn
383Hh6KpMtfsv/KQKv5DSwIMuS1ewDVXSZuQHiuRH8RYaIr3J6mY7lNQUSDw1vyfQhvxnHMlnWyB
kNSjRSTN35bHho8mTECSucjtXVkgcCzbkcEKhmactibiQtCPX4g1HWbBzjKqNkLsox9JK4XDgEmE
hpq7iqtAX6qkfKGTCUu7S96jBCazk8F/0EPrG9rzgh0f+ZHYMGxFtHG0VQNDJ7i/AGp3gILelb2Q
dTjsv7ov40klAABc83ymQo3zyBXL68ZWLUPVnmZxGHrGsXF0voW0jZdtzavOmYWUs2TttfPKk9Bp
45UKRXs/akQH1QM1nPtrfwrcspWzOHXmKwtfe5zONWFSu1RsGW82EQVxC9bKOqk3rvpFwXbDb0o3
0DIVVYsI9sRMxhpok4u2+Y1vk34VrgxLozsLUwYcCrfxZOU29Mm39PiDwcyfHLRs+PSbcD5pG8Zd
5/jHJt1p4qUG1rptnqso0w1pbhRP4I7NsTScc+X2lvfZYEbhcptmA93qcaRb3RZP3oTgTQeIQkDw
86N4v+ZK+MbkKvY+QEBffBJK6MEdXdLBIx698+fLYQG6x7nH9tL7zYUHQZbOyN0RAjANHRdZPakT
k+EFERqbNOe06yWCjTIVVyzG0kBgsgXdxzpAYwVS+sW0XrSo55eEevR3jy703b8RNmiwmK91WD96
86VsrjSf3SOxumqlaPRi2Wnj9kcAxJHAI2rsH/BE5B55pXjs36KeM+2CNZPTKlYvP0hXv0A7YvDz
9iJxDJpP1UeAlsRPdQrmypWNQ4yk4YWLsYvOw+RcZNaDkUZmI4ti7OzY6VSzR2Z2HaRxllBUw5fw
O/xFELMbTKs0C47zkdJhj+kTOYIGyvmNuf3zmxoxbQK8mpQrs8YUhFzD3aZF9K67pUncn1FMyJDh
L13BfFCzGmcsAGC4KbAYJBKLhgpi6QZsKkVFBNH7DvjQOQvAWvonzK3H+GksLKi2PsxfPuqHMcn9
2Eyo11DhXb4f0CJyrAVse6DDAQO8stPlGDPwd57dPROL3Ds2vUBXSW2WQFq6Q7F5l4qXveIMR57m
vmKIamKGBb3C0kveU2xGsgFzfcmEEpyJxp66qOPPrb1tt6+clOgPdNIuGLIZCfXKR8ka7/TF+muA
nhqyqpFprOOfHuf5yIErfv8o15IM3EnkAc7gDWBBmiDPIu/DfSuvoDTjhx4AziAwovrHFhYJAAiU
lG3iatW8wcEsHXtDkEEWQ7DQlgUIQWFlWiRuJp2BF5WNFpGZNPYLhN9cK563LGMIbQQw6I0L+TRB
lCdIFANy3CvJIu0Ybw0CdCBJiEVcszaYk+iCwah8OkODr8jLiZZoux8eGFSs12gEaUbVrK8tay/z
UnFESYzAb9c3PNXvA5lTIi1DZWv7WTyqN4VyP7jpD0IwTpgV/ebQSCqx8NWEz5cgQ+++J6eM3pVL
LaQsU6EJC/kcbO8w9hlBoNkMdW9m/Z4cm0SU4/lnOjR4BvAGPqBiaNfXjOpOecDscKWL7tZFXTic
8cUYOmM4OEw8yM+PJO12wJz3VsXrYtx2hNlU4hfcvsBoibuX+q0rTNFlCJIhx8et++8ezpcpolOS
bGMLJJHbbYoZkqy37GXV97wRP5shWrJVxFg7AhAhxL/2FSUO0jzCwT+tWMjasoVRjxObDukhKXvo
isqfOdaZP2xs8y73YF3CQV3RSxbZjxvZCN58cc7OKkyDkgCqb7uXRlphbjc/DMGzxLzqcj/scKiS
uvaVUxSbPvl4yaIjHbJmOL7i/kgwRTpanwnwGDcz3UhI/9awdtlB3Fh/jsybI9GAxeUoHYLrMiWj
rV5UFRhl3ZU+rLSSvyi2vtV5NZnleVVxw/Ho6+tDdIDL7YPzgMsVabHdtFHm501FgDTpIZJOdwAp
wm0f9QeM/SPIayCD+HgT678wtxmDIsAznHVjRMj3CR7KD9CX3ras5vKCS5Ruay/xUfvTDEo1XKzr
lZ0s9PRNRPHNdDJx14fXXZGxFHZYZt4IKFgvUkQOgKZfJ+0sXskHMm27gR1IK3wWsksbHF6SOIdx
FuTW93Ynva1AIWI6s94LeaAA8yq6xcr+pdTqXt8DKWqJQitbMYkzoE5k356k5L0051dNNei3MlVU
kvhAQR8uOk2bqIpacEo47yg5bPxjvirfYmXFyZpcBKqR8pF9GcgJlioVVWiNZHD+AfFXhBC4p9I7
UKO2XUYzGTtckqi6/des/eiEbbNAGWbUuaXTkYS0ieLiyWXswtBCn3iUEnD+1Q8QMlyLIqcOJ2+B
qt8mc5jD8fG/4cuUEp1sRJKm4IGXNz/PEVKWBMBvsi/SpKS+Nw66y5lFuneHRn4tBlyIY8wklbff
CJMchFvFPww03Ghac/esYzMNSzfmMbkcKf099K9m2RdyDtc/69FKYbahAG32/SYHDSQLvC4ffFt/
RfzbyZFGK9aR+rWVpgZrQu0QPWB0oWAXa9wl6nmIxEGojE9yAylN65aDHiZ7iZlF5d+VZAvCKRAE
1ptQDBrnuSbgppksaQTOisIc26U73Y5+DIRxQwf5XhpXp4UPIJ0EJjYyncu73dF/dbgYMmPCznDT
os2+S64gy6YC3Q5/71Ny7IIoNTmQicLo7ryO5p6dV8XIPs2fJucZBLqaIREOgxpuP1irZlUz6PB0
BC6EKQ4ufP3K1SLuVsxdX9P3f95hUurLWvYgn+CeFjGhsgfsVhEVVamVZqOPJ7g/ALZgj2oD6mC5
JEaVO5aMg5bPdmU+ttdM4odKLXIKJbwH4Q99/+COy7q1J1/Jm6hIiSlRVA2rfBVFCcxIXF2jIMJ6
AejVyMN25pxB41bPuTyDYUksoTEUuy8FyhkCBU2wUOKC81kEwlqZ08I8veE4hQlQ7qfmizTms201
g54Gp1wbJ6MPDQcktdiO2jqWqfkXNp/l2mZFBv9YINgeWbZyQvAneODQzUi3tF5fIUg7+td+EYk4
XJ2vWI+vDzS4a0j90w5GQKmUf3qcjnnB3J5vQvYEBarz/sKBr6b8JYjAsfEAaKDLDvH+3+Ie0xef
JeRhjNzew0SJRyAt27DHECNZx5lC6fTLcOqQQZRgWQwdsZpFlNL8NOdwXyGoz3vLt1CHeRZMZR9a
VndBhjGeFWH3xmlZ2aOVqdDbo9MQIIqmoJqN9Td0GGFylkULvP51dcBkY2C1LYRm0svJzBQ1NX5J
oBgQ+l23FjLWYdnbQ1w8lbqCDvik69XiwWzroexG0Wd7fnbBWY2Hf9RwQi391Du9rPG0HFY8inFa
eOX3sx95+z02DAhHdGYHCbu9bjSu7PFHzZLisRlBBjUpVP7PUpL4ewjR6lgX+i8JPK+EoxOsVQuE
eg4zi+uRxsHxCwz3e6K9SG5LkGQdjPTL557G0iyscTbr0kl6xSrfl5YgIqYIcc/rvRgaUTGoGtJZ
wJDISvvA8+BGRfcA/DcpoBgM4d9d6LDYlHeZhliAVWtVLR+lb0xK/+CrU3tx/l+uoyKE6bMKI20k
yUywJbmEgGwG8l21fvWsnAoWpfIDc9CgMVBNGOh06zrpcU9U+eBCLItZT0RviGqpUB4ZT/xB5oX4
ELzZM8i9mlxecdh0trGLR7OEXovJJzbZxdPMUQOrP0eOM3fQHtR7z6bFOhtf9Y1XwEtS43i4aAIz
Ola5stnbocTobRuf+GUCT5oGuw2dL6/A8yRUAlFcYgh1tF/mtCMuJKRgM8AEyfYcJedHfwu64d1K
NcBSMNQpiDCKZgaXdlJCk0c3ve5JF3PA5SZoLrsL8BVpA2jbL7jpGt54yPnZJvMnUemO0yedQlhb
sHgL8OVDr7hSYJaNQ7X+rGu9ibGu1+Gi3DRIFAkPnyo0YVK9dmrbNA/fowY8IqiZuk22x3Do0syU
d6oeMXPX+xHRZW4iZiaFRW8F1xbODYlP6klK1oL//FyQnfrE1YzaB57EAE41f2E/MR3vynTteml4
l/3kYOnQQ2k+BHgmEIgGqe+reE49XOZWO9LHqfzTQgpUeYLYgS9ByK5frAkWF4HyZg0Cvylp0xxF
IpYSUjai/Icyt659H4eTWiWu47GopY9thss/0yBH7pUmCBrfThnnGLXs8Ibr1JoK6J5S4ZtwjgSg
/850fd1MPATqlbahYcLoSgrXc3yMb0q54XNVGgbk/3OoYCuZ/88Vrj8um89uiLxGwaczr8kr82u4
dpvKHKpESLGE4CXfahUocEgWlgwdqdR00ryPG0h3SAkH9gZ2I8TdsyIcuv+nZ5vCPU6ZVZYiXPeq
yyBBtEDMcQlO5T38VtFYKwJGzoH/FasgKgMYlpadqpDTKVo/bPXT+zHySmSY1tmtbVNN01LDCprW
CYMDQkbO9YMP/aI1/ddhbXztWVQ0DyQ7IAY3vDuhV0Gi6XK8sDmh1LXisojziP0kYsnWXsE3HPwj
cdET5Ay+CYmFtYVGAc+2jYpHCVmBWzbmOY0gEbuPny9pHaRTd7CSZXJPZkk/c3Ed09BjkOi4Fqho
+TYtonRmBS0gUOtsxdKELeYav/JAAoqrlihFJtbQwdKJJ4qNqCFFvfZvI9+WeX7ADTJzKXk/IsPl
/3K+Tozx6KCw+1vgppcGXZLUFHQ0PLGV1IdnSN6JBI09BjakyyN4lRt9hvYnc9/gXG/jfduOhJJs
HdNLuG5k/YlfG++y7OV/yRmGPmoek2bAkewYBShxticMxcLh4iww9cBPp3SAlxJe83Kv8cNo/Ymn
3/0PCUes/lQhyFWrUCI2Damgn7qCYOBw5Xmh0TsnklOxAZ1lHQY9lcixAmCaubCUl/TfIlBx9WnV
ipcofgpjUsQIAGChWXlF/olIoGQwBZRW+T1yaW+vy+1IWiNcS4lzYrRq95gDbzdh1BZQ+6B2qYUO
r7PnRUDbj+jmb6eMqWl1d9dSAUNvBcT6wrdd8jDtW3troizP+xn787E4/WXcwb6ZdVCAaDOHN3Ht
Hbu+859iPY8JtuDs2V0w4LDSVMLt0s9yQ6EA4Oz0Tqv1fBtTEbLdTrU+Zi9MCUFvbFyhdHFu5dHY
RjN4E9Olt15WF0zdNc7EVWJ4KD2COsll8eDu74a5aMua8MBshbCuqBmaCTX3hq48shcDYXAqMJIC
zakBYGiwvS1lnTM0m0cO85ns5Vgz8lQf5kLkgLV9DMKXeREI0x5ZvdjDH4Cwam3ZFvWJhSs0Tw3d
uKVv+H9/MlawP72EM5pJy49iyISC+sEQF+mjPTtuSdhsn1g6eysUjnO67cY20LQmyhbhmbSKeILz
wIYU3hFpIczseP1wv3lmFMjvGfFOeTYPPnxJvJRXsDTWRCzKMJLgPWWEdDB0W9BwfY9ni+ubD4dl
Pjp4/CZ2NPLf2ahR9FIP9rT+8aP1mVuEAzz4jkvnLJWmBa12Hz0NYseLRUEXIVDM8igA2UFN/pJU
iEVEsOQnRVtr93Y2lIqOx9N8kDKrdD8YDJiwUig/2CUtUKgWUJw0InmDt+90CLdO+AI/N2L8mEay
tjor6Ql8x1Ow6LxOiEwV4htepSM5al5KlZd8WTMFmrGv3KONVZfcr1+ewhTBw53FTgaWKLWSRmv2
SmCYKzNihzo/RM/4YCN81lxB3uhAXmvqyziUSgos7Z2vjCjOu5J7buxDEkCuSSnb9ar7fq9bpssF
Gxbb7TV3CcB/CuqCCRnxXk8BWs1CpfdJWqCq7c2r9mnWiJbmPKwpuPlsaP8DSLr2NpEJcKpHh/Yi
HUT9beGbcYitmEsWyBAmTzVnpJt6/39qbbCWrX/A2MdKlLBGDPo6GfPxlrzgr2FfBl42VLOd6DnJ
jscLQhcvYYbt0Qx5b9GipZ1cPjZm9fmMLDTfv6LBhwxoY4ESBDJWVf0BljzxzXj8vslBPzTmC7W3
cf27/0Mc+OdrDn9qcPyFub6VfYctsFt/SXNuDnZgRms0r4v4JWxHcHcn2QIPoAHLAyK2/YKKBhfz
IM1nE/Fu3tjmGh+3t5M9uyvpJmyeTesHomq1cHrn0JQHqVlSLe5BqcVD981KK5DHnLXklgCMSS9K
NjAqyJAaTpeI1TsX5JGQ4Ohsecagiwx4EhrtGtL0Ho0DZxJpl8EbA0Iq6r6a9hwwkGFb+PXFGDUx
M9WPmbzjRIL0LAw6Nqzdx5RI4uPp4UuQqbReEK3hZERouQvrhHmZR80jkGpyMmbtg4rhCQtsV9ca
+s0mH/6/ApS7H5whN7SBHP1USW5rgIV2GzfQNB5rYxU2lF4Pdm7RHCvzafUmahq1bxyFJggsek+f
+yfn8qIxXgLHyOK1jcAX/R14kXwo3c789cQf2xo1OZ1oZ2l/2aprq8vhevECvtKt9elCzTd8ru6f
omfDLY5IJCO1oUD3cQo9ujkUwsqDfiFss0Jjb3ZOsvO0W94LNz8v2nBZX5lPBNf/i1PPFTiWhtxY
T9cAPYy+oKAqxee2uq6i+pu6BEtI+7JL9GzzHwsHqzr0jB9yJiZnG/bmZMiK48xeKlMywCbRfdzF
9rhzxwUNd7b2gW3krCX4zfnKlcwCrN6Gaj/M+T+Enzjj9awCP0gy7GhQpNIJ3veh7ugW4mZM27BZ
0HosSo+V9gsCTguNWE0wwdnwPHexE3bgnhtBcD9vhePS8+lEzkUozIsw9+cfmjvWBRNSeETZG5E3
0iIHy7YNmhJP/RJRMiBmF9EYt/YuozXssAbeUtgmuhH+y5LY4gLq2FBnb5GeVx9Yd97cLNpR6QpL
vM/ZbCGDIjp2/LQL1Oj57Tqs6VDxvRj2otbVkf2V1IJ1WKfD+gngBpU1shHy4O7kQRjqNXjVwF8r
qWLO95KBJqAtsKvMQuglvr8sSDzt2f9fRYCC2MfoGyNXx96BGXoLOiZJoNczD5De4cBp81cGL6og
mhNU/pdlBL7GnysbN1aJnfVNEdbLyNZAMw3w44nEzYDg2aMEWKL6IpqU4u8wVnxoI6pOqOSeYJbo
PQn7Jh2WXcCI34fMNTo2785rSKARRSCYf7y+tNFvsDJU2Czst9Lp+W6+EcBYbbsmllPGeESqM74J
lip/pJjsiIgePGPfOC0Jcq7XEa/CQwxGHXiyjDLFZeT1U5dSDuXsgjNypqrox+3blKbgJg+1JKoW
BMByppDudGF+WkTow0LSchRG81EGzdPsZB6kx18E6BNHKHQFChSfZbq1b/u/E6vserxydaerpzUO
EDVQ2Mh/+wTfwQWlCzDCO4Ca+v5d6rmQopawx3povqWgovV7JhBj5N5+EK5SqVMuCJxikTl4rjp+
rvyOdShcQoaOG1dSrXsbKVxGaGLUysNtmLl9Uo4THc0gqdKWomJ20C0AXCsZ120O/4fPymXjptbw
qBvRNfUoRB/Cv6ZeWDV7JttJ2e1PB0mYgIveDVOmEWMXUdh482wGfT+mPPRy/lRfivAD7XsPqBJN
V8x9YHf+MbOdC9ZGfkgJOuz+x3NcSMH0VEOZXyzS/inqj9npjCMfP7xO/zlVLwQVDSZNreiOdo6B
8KgzHhDf3yveS11IuxeqOLjcKWIyU6y2/9TS18sZSS0z+huGG8mOVYFBOnZ1anpil4/qW4jqaKqw
yS0FXEsVruu0jUHELmWEPsM/QU50t1VdPeFBgWZSpAMlDUAD/33w+zsdspd6TP71QxkA0RtZs66X
sBFYxReyvO4Jlsdf4CNkzICJjafBdX2rvXkQsiRA1bAfyg6TWFwnmMpZCL/ZqiJs+hTQl8AAzMl4
tHN/lR7mQQyd+6Dliq7OnwRkpnuhK5RJ+fZO4ZJNfdJr4gx3V3zl+gixV54k0YW/d0Qavs4u3xfJ
oZJl+oxadXTpXlj4LLG4qGm4uFVAQXVr0a4NJjK+IjY04PB1qvCMsfZbJ8xyyRl0PIk8Gj7d+iff
rnnp3byOUtaTmK3s1WrEGC8KcBsyjpN5oHJ6GokGxLwrpz1pXZzixSpXo+Y1MtXpCpv7mz1DSwLH
2q6ZMBcBGMPcVfO6qa9JiUc+A4zWVULp8XpM5gHUYo3Lj53cWHnEDg6oBlHvAkIwVok7KPxAqg8Z
lrZ/rQM9K/ndGrUBHhrNLlka+HmAZ+oKyha9EpDzv7PK9kkPHd8pegw4VCokquTI4DIfWT4YLz0s
MLhwm0Z2zjphyJ06lXyYjepZgrN85tszkTtXMIOl4VjcczYXybWOdkMNhuukMyEBAHlWkimacGzD
6Qie3IyXJQfIjNFXI+Qbb5wkTXQ3FN7MN7SsaRI2XUs7TJCGsENXl8+qZT5Hgr4zEd+HEQnuXlwl
rlnDj1nEQSsTJxB9zrGva4m6rZFx0QSH+xHhmTIOfdSj8sBdNKz4o7tJ5XNXakxAW5ogHIqCl7IW
+YA9sXi50TVye0wNgMQr/qTlCnzonqCnZGNcx9zt8KQnQIlOykicSrX8t1YL34wZgtaGkqpfS5yL
A0YkMGRGQubxQWAYey12QXWBus3WcPVvL4p8VwcHsbLuvc5RHL/v00knKmNgDG/E6hYJ4eMRKPRQ
AOpvAz4Sf9t87ldCPrB7IRAEJX+6gBbtG+TS6HOnt28LhCf5bHEXDXr5+PHy+7QWaCKoC4Oh7Qsr
MGPoPcaX/1GIiig0gH6c5uhlqT9O5kFL4pZ6W4Az/wHNlJN1a6bFye43oUuGUHMx7WMhTUAakZy2
7vv+FJACZ0JUUp1m2Mppr2EplA6IxAivqx0H1TmHTnVvyfTZQCQ/exr1rXm04+4t7zXmJa6QniCq
n584a3ylSGuEVn4WlKKzJ454HozK/F/giGDIvWx8+i7GzD102Ja5PMyCbo2mcprEcLFshnRvJk+s
k28QRDg6mqGDEmhRVzYiEKY3HWa5ZqnWGfZOxRBmP8ckq4ycEcu4lMAYeWwREeoi2zMX1evb0vnW
lFd7J17YePGMstpAmsxCo3LpZhnp/SHGg22At73SH7lmHnZQsgG1jF0qPSFheurYZup7/vqTF08D
62u7BUCItc5tcOe2uzSzBlvBbZzKTHpLNlFtZaRkdeWVNnqg7vA9lx4/reblj4PgdHLkkUSuj6U0
U1JykOyQqB8i36G/PUNal+/WuQKmrW3BcZ3SoQzdSXkFC0balFx+ImfuGvqtYkWGATW+aGEm0g0p
rUp/BSoMhZt7grEmFzqH6D8l0eGRFIXGmtp9t6/ZS1Ajsy3AejDMrJMbvHTk/iVbR9VCdQCrAw+d
1fX9C6QbVi9Gh0zjwP4UHCL+V7+zbv2LL20Xs6dX19JZFiMJY2jdpZLo3xwLxykAFPFFH9StQOAE
DZS2paQU7C0qkH2R4OktrnmyJJYmwWJsQ6JvyjnV0WUkqaH116rRQmdMLB+QTlKrZ8FgMKiSWEfo
WcI2aNU781qoCRLzHhqgakvGcwFH3L0yE0MZbLdl2V94Qw3xK399zHaGmsJ/0ZilVP4QCdnx9Yax
KiAEx1zSUrPtMoVMZd0niaaGWo7ZL7hJZOhYyKBvpDGgFc7as6Vf8D+ELgICtHn0AUj7Royc1dLI
V3IPBlV+D/4oTO/zWpIYpO+KE7bzELqlwtkfF+nOoc2L3Pl8XAJjKs3/FQheXooQKSB0unqOBcpn
m/pAHxD22Ypy4xR9wyo7IEYV3sp3EGWZG3E7mtGTOr2m6o8nbuurqxWJXjVkMJPrqzrtltp/ju6T
P9YtnaR89JzoemU6qVgLCG6xUgG/X/QCtSd/C9Qu7SNV7tYg+vT7hm9spDFX+W0C2ztCxd3aztxn
op8XEEeFny9O6uPiwA3EU+WGodF4VbZH0WyuIi+bsYO/X28dbtiGQUlJ4G+Kt6VnKBWcYeU+z1w5
Ur++N+34pV7a2KWeBUW/h8Fvp+kLWsjw3/soyCIPZHH3jfkPEK1tBon7Hbwioaf42d1sYDCgUlHt
ZEKIgSpKmIgex5qyM5/o4ev0j+xnr3l+DOVo/j4VZz9Ao/Wc91+67LFx0dliP6fIXCRk9LktbuVw
hgDqcAco5IJSVL1If5P9exAoESF3Z1Vb7+KOq73xv/vCmlo/dUrKC5Aap2Os3oOHfOP7YwAbWpaN
Od6PWGb3k+AX6eEo4hIFFy/43NQtGkk0rdbKxE71qT6ai3VETLfK3cRgu9MZNK+A0oBgJJlftskD
12oa1S722kKlkUi3f4d5pjcON3Xfk28zw21AwmMOvOWAB70QQgFR1FLbfnmsql1K4105gR7FYZS9
O/wlqeAlHYT2L+VPYBWb2Pej6XAWKbzT4XkDQbjTiB54EsiRWfdlUvo4UwJ35M+d5Vb/2vB+lNKa
BX2DV8NB65XSqq4fEM9I1G4/BQjW1FeF8k9F2bMCesirnbhq70o+bDlVYNgSvwAlpHq775LNXLXa
C8C1cv+BR64U6nYFoToEjZtoqm6zbzkqBZtR77i+cox+qEs4cSwkLlAd02XtSggxYwlmLmXL25Z2
+0ZXXJ0oJ1O0sI+dkGljAAKTkFrAX2ll76NMWeIIcfXcorPj8dg5j/IJoUVDeyOwswtfbf9aRxLl
MhODoT/DH7WCJChZTrZisHWaE4Wu4CdPJQKcpxw5fYTQx2lQNl6K+hujPclPFBkIOBu3XerKW7sb
Pm0+TSmNEgm4vhI8yP+tf6CEyZQrGXJlDY7x+9VE8GdKiOhPuU5i1O3AteWara6J0ZkLscpHaAGw
wg+R6zQ6EJcNZXr1hjYez9VFTzzc6tPsTonK0YVx7cJd4TPTxJETYPY7kFR36O6v+tCQBH4FiFuR
RMnNgq3f2MbhYX5g22KoXf6B9cSL1jrIuuAebPts+DQnCj4twOPNIaCvG2TIvlXV+rwfNrjEuBbS
Ze6dwCwhnQ7zQOMf7nx9C1CTM0fNEH4B876Ne5P6HsjkEoq3uw5l5ANRDYY+NQnu0hNCS6CR4JVh
Tw4Um83gqmH/4W+GPAgjl8blSipbRJN1WYjYjQ==
`protect end_protected
