`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
2qROw9/+OJdOEjGBwyDAcxC5FV84khzlKEohm6z2fzwvXaVAt8A+T700aM6+oyhlSMGP9OBrqjSB
n+6g948muK7fwN26H+rLwJH8sni0/5Y2PRI6TgZMg2lE//B+DDonJRokeMKWcTI1ESVozKwN/5Vs
tsiqHknlzh26yNYLFyMr9FgZgj82YZytZWlfYbpPoj74681jolJNdS20vJGo9TFnpMWW+PdDhKDr
kdEDVvkX7Zb3uysttsCjBrr7omw/vCb0j/Z/yYNkOtRRpSu4ix3aRtplJvN7ky4Cdk99QdiPxdi8
z7gHZpz3vfakkZKSjOwHtdoBVLezwKxoXMAFJN4Mx1FOCwYOXOF2KgnMCCHSOBpGjynqfDFKWEz6
gKTZC9+VqkdYRiNLzWXqPDdqDipFCUuhmlP4j/B84uSRnmESCqbM6bIOmgKCgeUJFh6nMYFjJXss
Eu56kMObf5OJNl/Hyb2Z7SHyWDWqArW9zE6xz1bT9TIsejfcMk0RG3C1gt8OMgz8X5tb2H/5dtuS
wo31qqCK/y5F6GOJWl6HxiKLGuriPHm6FuH+T2So3vd+HjUG7fgu9XRqmiTyw/m2TVvNK9KOz1qZ
oNwvXnsYNXC1eYrdgBt5ni1k6JnKKihQY2xvyvo2V6Rmp8G9YbgBJF5zHCUgwXkuolbIaOByo4T+
x1XnSOmXurt07nnE24MHEzLzAJgSGQFOHTnHGXtEDR8VpIJEXCmKi5tiskp4dKVI2BeEsqnb0tTo
dx97HseZ8vWLqwci0Kn9nX0xwDFCN+CRp7UTJlWUd1G7+0TkPdAfAbqfB6SLWN9AfWC/YI+wcx10
zYzcH0rnn1AdGOKif0tn1d+gsZs7f/RDXPSdsY5xFVaOANZNdpEtdvpeCmKVNWZoEkil8+EZDOVj
FaBUCZe3rhZ/n1RsI4gs2vbzXA76ldVvNDcrb/ONhe3v1bnAp95NMotlULhFvsDuDlEYYsRtBudW
+y5it/dYI44feFlck/aRr55/EiLBkYwqYHL9yuGlFyFDayss3tIF64WauQNav3+PekIXIe2VkKMn
VGRvWgY0W7JI9jd4+qRiOfhURVmo4AFjKYgHhjT5DjrJjqFF8xIUt9B9bHlX5UjKV73U4tczVp5f
zPv32upyoLNNmASNWtUe0v41QW60awJpB4LCsTCHFPemKLN2TiGrT6YxPSUs9844WlFWIWLVHXGU
tOKXMBnePdqy4JqSScNfUbyzTXMnAjuP5V+TJXBBvj0JL1lXMfyIKZh1HUugv8urPQHlkfZrMthE
UQsfVKaqLOuSbRjGfu78ueImtOrDJO2W2Alw6JujfYEV0QdNUQNigrTQnprF2+GiO9Jwa6PaFvl/
39oxFTEZChx/A1WWa0KR5nFeRdkGFGbQj3mwRrlOIf5d3BjiFqVjpJZB4OZcCMHajgDqo+BDgZ6L
1wKBx2L9cooD8hZLMzEsVAB+xT2SZ6fCFjY1S/6+XplzVIae9J3g9Vuqz3vm0q5s7doY4YKTRrnt
hQ7dsKGzfZtK0XjTWqDGUnEErFmpFPp9OubTnxeWFh7U8kw+RQqsgSCB+XoeVypvUbLTalr+kVPU
Q8lAYiP0sjE1VDo0PIlq6J0wjN1fKavVfogpzZ2+c7a7F0mcAczf2sN1fXyta5smH8WTxjrJRSgF
TmywnowP0LDQUbv1NnckHuoQjsBy1SHQC8A5zbmc3sxzSe2CehDWmRyITE/HDWBumzxZ9Bc+Gmzp
UM4nvGQtHzXuU2Mp8iuMynXFDi/CNjpMGvixpIHzAqMS+C8SPQfc0YFmWiC5du8TJ7KiA2FKrXAD
LwCRAC36VkWlDfuZHjG2ZjJc2eUX5zOUyoTClvwU2Y34EfG4zS7RrZ8uScV9Qoz3SGWZ0LVQh91j
76cQciypjErtyTmO6+Lt/DxVjR8dx++iZ+f5BGDPORyl4NIuz+vZ5u82d1IxzlsKLjdyWqErZnbq
e3QAkIG7A5XIPNXlVQ9UGVj8L10hCYhRb8j5wJiQmfkO6ZxaUpOjr4Olfh8tCtG9/5ihLsuHLY69
DbqUWXg/GgfnKEgc7YoNJLPudOyD1bRW95AG7i23AV6AWX4TJPGc3vMnr77b
`protect end_protected
