XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���	&��S�~�R��� �� �	�]i�x�&!�fX�r|�6�ox,���	�z�X)��lnvۀ�*L%/E�9�u,�������Y�ābȣ	��yY`o��j[[��s�M�gxe-��l!JI�K;�U�c�e B4��ː���r�a�<X��O�[�G��nUK��,:�YO��s�����l�� �,�t�{5�(�:�:�{���˴�w�v�<SMX2D䘯�h��\$�V���ֺ�\�������!�V��>�֫�;+%�ms�}G 2\�8�K�6�ںv�JS9�oD�)�RK�-�/�]����MY��x��]l�1�X�bK�w��T[�ɚ�Չ���z��̿���JO:���kQ
��`�)Ȭ��_���m]23�a����y ��7�G7�z������?���X]�e~Δ�8X=���k�`E����̷��D��9��Ӫ�F����������L-�A��^D f��f��U��`��B�B��DϠ���'k9��E}U�ZH��*�$�ܹʅl�U�V�]IZ!�}4�1Vҝ��cw�6��C�Oz��J8�w��']�ܹa��4�~����O?�/��f6�?��v&<cB�	S�9�Hbn�c�Ǳ;C��|��1�|�r\GK�yQ 0��.2���G��ւ����P��܎�V>����ٷմ�:��48~�=�n�f!ݡx�@�����E��~��!:������؝>&ܳ�^ $�}7eD�l����|�����NXlxVHYEB     400     1c0�Z�Oe�%qc@�1���&00L���Zr=�Z�6�d-?���D�������턗�tXy�-T�ޓ<���08ʲ<ԫ��K���f�O�*5����&�X������H!�^xK�U��h���q(s=�Ti�"e��{Mu-xY���A�2,+` @=����)x�L��
(G���12[q�iPUP��>��&kU2M��
�A�R���Px~GSu��Z�)�!������	��'d��I���������sПSL^��Gh��4��p�b�Z�y��(��T��^�&@,�FæIO�7`�Q�g�חK,�!�le�حbh��}H�u��T�_�O����Rp	P�,o���Y2j�B���$	��[���Q�_%RU8a��u�s;i��DJ�K�&^0�F�M�R���/I��b`��PW�$b\��H+����[�f	=XlxVHYEB     400     180٩2��ғ���&��5�RU��p�1P�7��s	5�T'��j�;�H�;>nǙkcQUcT���1f��^v�g�p�&�_�����P�ح�8<��3=�r�9�ݳ+|@�D�X-��Խs�@��*b&�9����(N�:H/��A��k4�����j������7Kh5{��J�8*W�����/@�$�Y�-��q�S��)�,�R�3��F�4��e�~�r�I~d'���Ipr$p��L�cԞ�9����i9��#�.a��7Q�F�N\��s�ZZ�C��m��mߡ�������"/�.�O�'�!�]t�U�u��:�	�gF=ө;4�	�;K5�<�"^v�/l^.��G��{����mS�%T��Z7�
",5XlxVHYEB     400     150��z�di9IĻL��]>�3������������^z��i�NBy\�1.c�U$�\���=�Q@E�4��K�y�M%�l�!4�|�
hU1�@�ɥF���d��.��t$�fC�Kg�Rb�8�~`�K,Z��1̓i'�#��(~�NF�d�3#K�����3���.Iy���\1y�3��l�Q;�N��o�$���u�=OЬ�2f*�nY	(z�I��a�N���ﻙ���3���Z��^um�:S��O����(h��9ro�w�˚�_��ۑ����K�&�`�[�e=������������w��M+�=�i!F�ѡ��2��Z���XlxVHYEB     400     1b0^��/\��f<	��P�K����Ya�@���\|�� �'W
'�@Z�n���A��wa%��=�<�RP�<�*N9�G�SdLVo����0l����fwP�q�kH�p|´��#JDZ��"ƶt~��z.׍>D��~|���e8�7��)�ԀXQP%��Y#��O.��$5�tD�{�ꄝ�5�RP"C�Gv�J�
`�V� ����Qn�zY�r����L�I��+��x:�i��PRj��a�(ד�ʹg�<)�g�0�%������P� � �wf��/�w�V\���YZ��i`���kW}@��z�[�HVu��VǟR�P�&�Ω�@�魹��ׂ"|��;�O#�O�{T��1�k�'U�"r=^
"��l�5h.S?PW�Uns��/���S|B�Z��M��
���Z�s���_�֕6Ҳ#��M�{
9B��XlxVHYEB     400     110�~����j��N�d�6v��S���C�48�@*����&��J�%����@(T�PT=���	\*:�WF��˛**^��o�7ֱAH�7ޠ6H'�i�V��jBY}W���A��� |`����wO�=2�?�`eXN#����]Ĝ��<]0}:�O���.�D� }��!	l�9^��a���&����9��ʬ��c.eH�E=����uǼ��n�5vQ���蓽�N�� �ƨ(���]��������N�s^��	l�XlxVHYEB     400     120γw��޷*�!\�o"�j8�����l�$���/���t�W��1�q�Tt2���
X�ʯV10I���%gM����]�����3,/G�B:��s���"�Sj��9�kd>�qu�ne��g�6G����ik�F�
��pP)?�	ݶ,�Wo��L��� ��ԏG}��n�j�R�Qo�2%�a���&��b�nf�7��^��m�K��D�C}�2!$��s��J�!/�c�s��B��f��>#΀󼗺Je�6��������+�,S�=XlxVHYEB     400     170�e̲M���xS�ru	�j�'(f;��Y�Ε]{��IUR��9Ģx�a��좟�c�+�<z���H[�uק����D�ͬ��W_'������Q>� �ſ�m��w�͛����P���?�����K/��7�b��{G[(�o�č�t;)�N��]�2ٞ��vM �.N�~�t��xr���]�[�>�E
3D��y��Xy(�
��2&s��IR��Z�'Z�O�M�nI3�f�ߊ���o���c�4gK�:�vqcjĴ�BҲ
=mj~b�lK<�3�Ώ`O��o�OMܓ2K>��Z \��9���Y�1�!�X�Err�.��o"�Т�h�W���W]����}�7n\dhM�"�XlxVHYEB     400     100�u� �[�@�1!�p¯�� �z�}��L��m��n�$뭣��f@B��,6
��()T�1�?w8
ONq�Gl�~Q2���2���^Qfrs�u�_�D�T�9=Arb�
��Nu �@�4B��Q�E���=���n�c"=���L9�:���`5q��ܛO���yX\�s�Z��e��n|{��")�3�Q��'vO��<f�>(�J���ݏ4�Uo���T�;b���2f7A1o@A�/SO,C;�ݺ�&2꭛E�q�u<RXlxVHYEB     400      d0 ep��(V1��橇��������H�Wf@Lճ?M��н,��uŴ�k�$���W2����fɆ2��&��5��ǀ�����z ��k��0;�H1rCWzsi@'���� \�|ַ�K�Y�j~���m�q�!��`#��9s�r
{&�#���bj_L��� ���)@i�d*��$<)��K���0�L<O��+���f�C�XlxVHYEB     400      d0�[�\]6���e�-�'Y�\7�u]�_��P;�=�����(��?������ț�7u�-r����ļ"�]Z�wq��M%/8XsY7��=�#\ī�HĴ*c#1��ш���!�$<2Q��d.1�+�-����2wU�t������� ڒ�bkJ%7('�bXE�Y.�����p��������^�L�1��J�+ XlxVHYEB     400     120EP䵟]& 2;�&b�4�F"G���~���ì���)oZ���La������++<+a΁T7���~�3.���	��Q����uj �Q��c��+�K�*ZH�p}��������!�B0ۧ%Y���|��\�q�����?���v�3!�<�T疳+�����7�:|���3S^���h3RP,��dP��w��`�����)�/���[,�W���:77,��_�y��>HԑKej,x6���T&Ks�՛�b�u�Z�_�/6�ׄT�$��i�F{^^{XlxVHYEB     400      c0���d���@�#���1s�]D�F�N6����OO�zOS!�=X�Ps7��v�Ջ!�]W3�*���H�eE�v�.v�>��+�b<
}:xC�A�S�I�ޜ���qM��0<Ύ�J�h�Pt�{^&��I��.�v�Y�Z��@/jZq��yAx�A��9����e�|�V;[:v��U�qG��c�XlxVHYEB     400     1b0T wp�s� �Ml�5��Q&�m�:���r��
��C��f���b���@���Cv6{vE����H:������.�1�P�:s���h$1�	��h�r���Kh�c����0I�:�qv�����@����p��R=[���+�n���.!�����Z���+?(�y�.a@F̬�4*O-�{�3��vH!�5���/2�̑���	�o!H���:ک�柪�
��ڳ�jp/l8�,�G3)�P�|n����4_�����n� AQ޽?�g���w3��@�뤼�x�b���O��Z^���a��o/���ŀm�m��nn�4!�����K.rf�O"f��GI���պ�*l��^H�6Q����o���p2:��kR�ѿ@�z�	��q�����Ms�7�j61��=�&cf�Jw�� ���	V�P�0>�XlxVHYEB     400     1b0w��3�|�{����N'Ds4��LdF��{so؄šC��OZ�$筂�8 J��*���c�~W�Krի�%ו�@��A�����×�F�?e�A"��g�y��An����1��`ʉ>I����3�'4�RE�i���.�r�)�&�����K�W�,����b�3�aӊw�jpoK�5�k���۹���R�K�֖��*�狱��?�u~^8�$8�gi�XX�H�@�s�\�Y�`C$���)�"=<��ӭ����"���vb#���/'�%QW��#N%�M2H��UQ���GF:�5<�Q�� z�X��E!���������ᨒ�8 � �,�V������U7»}�� I�얧��f�.�M:�~���0��a��(������R���f��9�u�И�V�X�a��~U�r��G�$6���%~ک�`�XlxVHYEB     400     1a0�4�9�`��pz0�ꓘu!Yg���@q���x�o�L��KcS�����~�X��)�D%��Z#�l�w�r��	A)�l�½��x"�M#�ˑ��'�Fhw��N5��zc�1}� ���y�p��"��ډ�R��虹Y��
f����<�C�Z� ��5R��Ղn�闭�n*�CO<A�D ��y�l�n6��z�`��
�����͡�1U�
��2(�'��2��47����$_lI��kN)���M.�uA��d1K��a1Ŵ1J`;�.}��;��N���*&��moy�7���E�_%6������ဤ�E�s�/�>Wµ$b��@�ӈg��"��Ty�W�V�ˁƲٝ�g�j��W(2/.��;0/�b����OG�{#���G�z{�XlxVHYEB     400     140�h�5��Ё��?�B����`�ˑ3WWtTi'��2����D�VS	A-�܊���w���"�	`�RSA֐0<Ά���|�*���o��b[v�C�&Z���N�@���c�'�B�f�/WvmҌn�ҙ��G5c�1ɦD�	�-�w�}��J����y%]#��(oКV�;�<��j�U�6�Z3��}��]uT's���$O�D2/X��h��(���7�g<S.WɈ��B�C�T�W(��_)0Ke:��߼-��p�=��
H��6=6J� -�/q��ק{ٽ�;mjT�tţ.�o�'��v��AXlxVHYEB     400     140��+]b(;M��WMEB.%�7W��U�<?e�3F�-r2ud��~���D��Ҷ��G�㢅�T`�"������P,���vI�7�~Y���\�&��������+�<;p�Y|&#���t�xohЬ�m�����z��X��ԥ��H��	~|�U�둪oϊ�ט}8E�y�b�,�����ۗ��2�CAccC�`��^!lђ�%P�_����֩z��?EVV�o�	�oN?�ZiJ��j X��$g�>4lɩ��.2��f��W���[�N=���<qn5M&�����F�M5�酺�����ǶsւexGL�XlxVHYEB     400     140Zvr�=aX��"]!�Yƽ�s�+��)�^��v���yє��~�(�@ ��a�lfH��зU��"�a������gE��'T��ω��ͭj�=U��0mp��hް)�|���M�z��Y��+x<���*-�A ��aR{@�,u��'�8u�7���L��ԢaM��@�%�e*�qD&ܑ��������r�ŃJ�\�=�E�/����	7rHU���U�j���}Z�$L������H�;R��f�X��G>� ,]�*���d��"\�J�#b)K*��w���(�g��?��T��1����~�G1#����MZC�O�/�:���XlxVHYEB     400     150JF����Z�f��eՑz1�F���p.
��)&�~b@�����4���.THKګ/���{�:5���(5�
48I���%t��.���󫥯�k���{�@m�Y��;	����	������X��ŘD�X��}d3Z.���`	�9!E�Q��EM���G�K�v@������N�IQ���Lh�n�E�=�T��c���H����p^�~��_g=z!��	�W<S�Ai�'�e���VJ�G�����R�?�lwaCA���j��E� ��������WԱ�0���!�c;�;;��xB]��,�Vfx��"�N�	�Xo(��ܓ������?����=;�'o(��XlxVHYEB     400     140nAaZиY�,��ڇ�&�&j�Ow��0��%�
3x9c=3"$e5������A�t�ͩ/!���U���p�^@_U�Z��Оf=GÙ	0�9����U�8�@g�1�0��O��C�!eX*��4i S,J�·Y�#h�넕�9]B�3����D�(7�E%���^Uħ|� _�(N�uvX'4��fIC�#���bț'�g&�9$�=q�D�ub�[dg�3 ���6���?:���>�q����58fc�q 7m���+%����w��Mޏ��m�ץ	IV~�i8y��=�l.��7���n�+�c3��z�E��hXlxVHYEB     400     130�T��x�������)ƗB�۔��4`��7���\�̠н�X_ èB� ���U�!P���+߂N�8��w�U0�i�=i�Z}&�DO!�,��zi��ɲ���B:X�������zMj��~�<���
�vX��ChXX�$�N=���K�۱vp~LE�^L�u�Ġ8���n�Y���⎊J�(���m��>��{b�)��/F�|:b�b�Cb�|�:�*?�ET�?�����^
S��`<�I�9��~��G.�r� �ۃc\:�9Q�C��n�������g�$%[�����q�_׶�XlxVHYEB     400     140@�{�D�Ϭ�ؘ�*a��	A�'�i���!%�����!Ŵ���a�C-�L���7�x�)����Y3�-ɚ	4!/zX�U��(F���`+�f��1������MC����V1(��`� �c�KS��9I��`﫼:7y_��o�`��y_o����S_��k*�[��/��=��ي݈��O`=��x&��ݲN�e��[��Y C�'ѫH��e���a�q����T��&4v�^羔�7���^s�_�Z狔%�o�EqR+�H)��w��{�æS��W�Td�[��;տ/��tb���!?N����SXlxVHYEB     400     180�NW������/o�[/oD&�/#�Ezu�O����э4y+�vų|�,��>���}��}Eh��2Uw"T���Im.kW�"��_p�q���6/���J���8�׾��Z�A��pulj6T1^���G�9�e�.<��d|i7����J�v�X��n�r��z˟�����[f�-�g$���zB0�� �~�R��7q����,�oB��-aD�NK�����D�\�"�ʐ�{o�坽w��_Y�,��EX/g�D���M{��~%t��GU�Kqt�)��*���o�L�OJJgf38g��Q����~ڲ��Dc�������ϳ������m��J�Et 08���(7]D%?��
�E����>�rXlxVHYEB     400     170W2K4��[�N��c����ν�0Ƭ�O
Q�l
���E�h]JH����{ �y�o�����US�ܔ���M��FK�lE��F��{� ��ֈ�{H�g6[L��]���:�`��X���>f��͌˔�<��VYS��zG��'M���!��k��N�/�I�z�~�V��e+�kA�>`	,����x�2��g_��f���>�|�w��q��'2�]
�P�W����Ǟ�B��A��1�4_��V�L]���Y��H84u�K6���?�}�<zet�L��5P�������n�c�N� ŝ����j`�����M3y�E(����B��DYx�*��FS���	r�A�����4������6�f�bXlxVHYEB     400     160w�P�vn�v��v!���;W;v�_&�gݵ*���Χ?s�.��}�ykE��3���^�Y�vEӭ��G�Y��5@�����I�֭���$��K��\K�<�x�R�H���̶��!p��)a��v�Ẕ�,�TM_ſ�11�5�ֺ�o��������Z���q�P�Iv�%4|�]Y�AF2��)	��+��-�0�M�L
Y�?T��d툖iR�s/�P��Y�ë�����%`��	�a�d��j�g�� 嶦��ʪ��7E|�~��ޜ��`[dE#���V���Ȫ�k�E+1;�5y�
���C����<a)���k��L�n�i,)�\����Θ-Z��?��XlxVHYEB     400     1c0O�.��v�����?�!c�lB��z̓����$��
aJ�8rvu,3Qԁ�t�t��/�a�M������v�v�o�[�`�^V�E�x:𲴦�k�,�7��F7�g
�a�/��\��}H[՛oD2��6���]Q$���s �&����-��{ <n�����S#B����Cd�0�������*�[
H�������w�T�z74���jМ�8c&�<s�� ��S��K������+�$ٲ�X�J}������k޿
����`�����Iz<�?��Ni�Zh	�H]Ӻ/�E�n���[���k���,�0���(28z�NG�c	:�_��:f9��q:&�SKy q��BF�k�Қ\�`��߰��3C^,�����6x���Ä=Sp��SbYg��������J��s8Ռ�9�:F���a���9%�� (RUD��Eӓ�B��BcXlxVHYEB     400     180�br���9�w�"ʩ|�r��iW(pv�n�����oH٭�Ѕ�'�^���B�z�N�����~�K�O5��<��O��JY�c�P�B=��#�A[J���W��d�`J����}�BI.ܰ�(-)�TD9��u��ɘY�I�����"�i8�^��®�3�y�ȸ}eQv����y����L�6���	��V
LT���r��s�V�]�,��2�q5�4�^��żb��R�\7��k�"��/W��Ȳ�i�:����5��m׶�r�תđߞG��1�QY�ǳ���e/����/�(o:��dW
�=
z���"�0;��}"v�3���[ʛ��x���X�v�o!��*����5+���E�@#
{���XlxVHYEB     400     190�=�gT�n0*�_�l%T=3��ct�}��'�?
�W�#c��!��rX�\g�+x��k�(��.���_�GD>�T�����*l<���zaZz!�min�"�or���s��O�WQ����T,��%=?�z�i�ê���{�3��"eC��d̡Fʷ�Ѽ"xr���(���ϽQ�ѝʘZz%����h�{��
I������I%Ye/�%#������D�G�<���?-���M���ò���/����B��"t���_B:En]5=cS?�Z���;��O���Oi~N���[��z���˺&]�����D	�}�G�Zd��+Ş��Vo��f�EW{��Ԑ���k��X�D���,�5��+��dj��"�y�tn��JN�����a��XlxVHYEB     400     120���qKw��bF���Q��!��cX��L_4y	��b�Dlg��V�1�殤��kpdQ���L�w�)�B����/������!o�hv�XA�~�Ɲ}h��ׯc/�%��y��@�.C(C�����/Bj�_P9�B+���~�/ЪW���nn �₷{N�_TEﴽa�r��:'�s"z�<[��6�亡jX=~�
�0��;�a7��7pM�T��Y��e+��՗IQp�����s���:�ݗ�����w�b@�	1C��xn����E��q*�b�5�C�
�)�kXlxVHYEB     400     1d0eS�q�Ty�#<?hg`��+?t�3�4k��P�('R#�P;	��x��Ay�o5�֩�^�5z�=ƚY�)�}�Qc���b�|vf lF�@x4�mN
�zC0�r�qV�e���da.��`b�����a���sFU�a
��)��nO1��P��)nv�Ŵ'#�G����x�=%jH�Z !���J���ܽ1�a?�\Zq�l���K� �xq!��IL")&$8���?;t�����Yw\��:_�2m�7���t��(Ʀ� �#:�{4�k�t'�~4ޕ�UOH������,X����h���@��7�ދ��c����Ʋ�[Ԏ�]!����m7���JJ���������M[�f&x<W�q �GWm�J��zB�U�l�vO}5A�ކ����5xj����4��I���	��6s2���T�����4���<u��`[���0�fzXlxVHYEB     400     1308O���{l&iU*�^��¸,�i��Dzj����hk�$=��(	�������u֩��M�>�5��o���F���ӓ��F�Y�o�-N${N��V5�)��L�{�������Y���p[r�Ti����&�<�����U\� �砫��g��ʂ�ע�h���
��k�[�P�:C'������V�ξ���@����|�{dg�L11H��~
yB��R�9%�Ur<_�,|���m�1^�������΄�9�ٚ;߸R&�l�a��C6"*��J��,!"��U-�o�Ԅ�q(iXlxVHYEB     400     110fq�����^/8�Q"��'O��#._�N=!N��{���b�uDM BcA�&G�����a}�Y��
	�R�yj��s"��0W�[�I���<�E�~��'��<�6�5�}�ëӁ�z�p����&�Ԓ'2�La8�]�j鮣wK��ج�!�dĪ�����Oy"��f(���V�U�f�lY-���L��c��M�V_������l&Ra؉+lO[��Ƿ�l�#����2�w�:��� C�
������*�7�����K7ω`EAXlxVHYEB     400     100�}�|D�>3�{q�{tȟ� >/���ۇM߾��Y��^��;��<TL"��z�7H$�|>�b۱cm��j�
᪱�?�嫪��D��x(���
�K*
���}���M��M��9O��vrr������?Bo� ���➃lh�_@���p�T�#�Ɣ: ��"��Ь>�3���ݷ9*p������Vt�4ɓ�̶ݮN�eJ?C���wO3��NC0`w=2�v^�����ӽ��XlxVHYEB     400     120�����.�IF���Кk�P��MF�ȅ��8)�(�]Ē}-z�T�h�-=m;�Ա�n����%����������w+G�^�{�m&+H�o�yk`�X&���ޯ7W��,�	y�_�rH��""�:\	�Sڇ�ʚ�����hf��r��!��Q�t��'���!���0�Ƶobǉ����7�d�G�y�w�;�}+��B�(Q�����'���tWX�b�\�~������M+����s	;�č���#lq~7:F�0����ɯv�g�5�$XlxVHYEB     400     140��}�� ���D/�������+�%c�ϴ��1�{��e 2}D7��jD�04�OS�ݗ�v��T#��V��j�,/?�H���B$#�qw�����*XN����[���VN�3Im`����b3��9
ys׿	�<�:���8�b���4���4ZT�/^2�����"c�_ⶁ)����m%��˷|����TtS�9��{d�<�|{p����|���# �a���\ip��Ϡ,RٸY2�����-p��)]�·���� �'���"�_�Э�π��tyw�8���ZZH	%%�\p/*5vu�%��?�a�S�XlxVHYEB     400     1b0JT�6;tA���2�nQZP�;��t�\VD}'�S��f�Л$ueQ�h�Vkܤ�ȕ���`���{	p�BL�?xL��3�ҽ����7x�AwW�������5Q�2��^|�aV���.zwk�R.]�8�ݚ����եѮO�>��1�:�WʘЦK��^}J��n�约'0��}{����t��i�m1n| �z{-[ν��^�)�Ù@rMt�"���l�}߰�BF�wF^ܐiN��>�7�2�%ֲ������켪!nb�Ύ���M]�_p�`;�-H21�m�H�Ǜ��ԷF�eU�I6� ��'�#�����'gO$uﺪfQ���Z1K���²�����4�P�UH5�. ޴�y����0� ��ெ�p`u`�AM0N���D�h�ڞ ��V6�9@���?3 %7z�hfT!�XlxVHYEB     400     130���D��~-��ĕ��"]�A�5�l�"7��l�r'��]�������l�I�In��N�mF��~��C����;�X�v�"��ؗ@`�Ío/��o\q�-�j{^d��Pd�b����4J|�|����'+�|Q��F"�|sRaOү�Ss{~!������OH���tϜv�"���^�7�# 4�עQvm��E	��V>��D	�o��˺�����>oMi¼��x4Q>�Uj�4���}�{�+�r7�*���E��e)���~B���#3f�>�(���r�^À�iYXlxVHYEB     400     170e3�w�Q�
�$�+��X!w(Z��
�o����c���VH�,PAP�s�:�����l�7`u�,�)A����Dp�w�xnG����齜,�%Cm�v��&��-�k�&���G�iI��х�r���)a x�F8S�R��(?��%�17��c_)���+M)l�r�+A�GU1�ՓH�=�o��J�(��Jey#1�!4��ؒ���U��^|7h�l:�3�b�.��p��XQBp�`�ځ'�W�I\��=>PK�..LU���p�3mIn��~D�l�`�1���,_��,w�p��4����ݮ�y� �O/�Y�a�)��8�dqC\�g�qS�r���* ۺe���fEҡZ��� ��"(�XlxVHYEB     400     120����v��d@�Lו�Q8�(�격�w�"�D�^*�c�oaS��E"`x��u0��)��O9}K;zVw"� '|[��haҿ�:��e��N߃Q!�ugdٲ"�4+��ô�� �X,��v:�ػ����zj�^6H�>��E iY�`��-;�d�)i/�-)��ϔ�d�D�~�D�k�-$nB%�&��^䅏%LåH�#�gy`�'l�Llf'��:M
������|�1��V�����.+�j���c0��Î��\���|4_Ҋw����CTQ�ϙp��f8\.�(�XlxVHYEB     400     170>-9+@Ѡ|��+�jl�t�^�8�m��@� ��i�C����p�E���9���p�����/El��� 	}����O�Yp�_ ��u���!!�0h/��25�� ��೻�2-�<����]c�b2�� {�{��-�*� o�@�"�8���߭��h�墶/Q욲Q�yr�gG��#�� @��o��G���ϚKH2Vw��E�T�Em�x�S�d�Ợ��XG��j���^x��I���K��R�e5iR�^D��4o)��}��p�d)��AQ���%Yv�<�-GY^Hh����֦��l�����$#)	�s	�YJ7j�0֍�bJMڪ�c�?�Ҍ��`������"XlxVHYEB     400     180�s�[E*���U@�hj��������⚖(�nXtnɖ�)��ds��x\ہ�d�fhף 
ژ�Ju��a�册��hWF6���z&[bS4M5|�$�r~��r⊣4�[�4ԙ��6���g0���Ib&c���)yS���C�r�	�y>*��́���@Ҏ���KE빊3m�ѮFc*tu�)���dӇ�dQ;���<21ԲG�D�#���Ypl���,������N��<���?�7��|��c��P���	<��޹�[��#��y��A�d��]{��p��
=R˘ۍC����Ur��h��rj�]�=Ut��k���w����@@��w�n�n�l�~�&(;�EY!��Ѥt�c<٧Rn'!�*@"\K������yXlxVHYEB     400     1804QPs�(Cg�!?{��b�0���/���K/t��� c>|����ߧvfp���>�ih����]�*��Ԩ�����4朇H\&������͙�:6��$�"�jQ	��j�?N�Q
�=�����i;hT���r����pu�Vi��~Y��2��@�`���i�\�
�K:�+sH�^��q�.�Έ�*}�qi�����C���:��a����ֳ�������t�΁|3�{;b�"�t�Ǫ�nm�6|F}�̡�"�¿�y~���趬(1熛�d��c����Iq��йl��%Y��yQ�mƳ�i��KU�i�s�l��o L����glE�6��n�L����8�T�!�NM<O�Y���k0!(��=o.1~yӷfXlxVHYEB     400     140�d`����������h�'�h{�ց�<�2�>y�2�>��P���ܰ\����2�]��lS���5�j�Ǥ0ziH�W��$Q%ejA
\�qQ�D���Bh�2�EVVEA&���I����LU�a��`l��:��3O�,���%Y��y�O�jj��/r�ͪ�0'��0o9�~�<b������ݨ�Dq	8�Ҷ�����yn�d�J(��p�Ӌ\ i�� -	����� (�����ԛP9��#�(8�L��H��Z���>?<lQK�Z��1�P鄤f���h��M�r��ӱa��Y�PG�%����\�XlxVHYEB     400      e0feٲ���-Lv��o��aCO�;��V�
C��-��.�n1��Tlu�}��x�VG�"ŀ���M�if���/EUw�H����~S��-��Z��'�ҡ��ql�(�B��BWd��ڳBL^<��>Y�O��ͣ�o����]&%ڨ��X��� xʯ9� Ӧf��bԌ#[�$`�ftxJ����	�_c^x�e�_V�T�5�G�S��rs�B:cӀ�?�XlxVHYEB     400     100sb�Fy�pM$T�=9�7�oaD����	��d#@���\~q�|<
��ӈ���a&������Y�u����1�� �����q�P$�z5�_�b_�V�B�@�J�3b�I�L.H��x
y�/.��Ug2Uv��q���2�VRM�.�E�btt��9=�o}L�a�L�;'s��m�g<}�o���`e�$Q���6�F�q��=�z���?cH�%.K��zmA8������u$�@ ���
Λ�}�/�p:XlxVHYEB     400     120~�u�	tAP�wi�fk��z�Z��z�����q��;3ש�!�2��"\d<��{�� 8*�Z�&ՑDc�p�r�yGf��6�T�L{:H,�_�?t�a�Q�"ʽh �q��D���O��
�zнFTIΦ)����wc�߃��w3��͟�jxi�����8}Q���[�0$~��o������5%�F�}�~e�}�%�-,Xwd̀�RO�����ir��n�����e8y�� "BIN��D%���-9X9�Ņ�8,DLy�����'����?'��XlxVHYEB     400     120��s�Q=���<�'G��Ue?�Ḷ���nK�j)��q�������P��~�]��l9�L�����NM��,���O6ݫ6D~r0x{�K
%��C��\Ո�.@��>!�C�:�
Pa��<�1WiM� p�:~M*����&��0g:P~�=/�ț ��t=��aiJ7I����D��kq�G�Z4u���ݤ6��W�9��z�{�D;�J�9�:��
�~�s:h�V��WB���C^=s�&���̗~Mnw���T�k[��(F��D���gU�x��w���]M$�1�lXlxVHYEB     400     170��ɻ��ɓ�4���H�Sf��WLOW������.����`���A@9��$��Dp�YW�;��gN/	�8ʯ1�ʥ��2��x��Nd�U(�FE��KKz��vq�t7y)@�?Q����Y���-8+�Q���4����#�Ź���O�%sp=�R�4�G�/�'��1=���vW(����畕-��� U��f������Cɜ?GA�F��{,�����z��-�H�Ϣ��u�$ܺ�_�-�Nx�2�?^sΙ����-�a��8{����G�F���!fC�"L�d
˔����e��yEe�c��$ĭ��""\|.��t��ǑE�*���`m���s�`��g�J PS0��]j#���ӳ�C�Vc�XlxVHYEB      87      80tM�	
�@XcvC���W�SB8���X:y��\�.�겡����^R�]�E#��7xh�V�"Ȟ�J�7x�ۄ]���X`.��)�{[L��N��S{�@���x,':?ûv�G�(1ܿK�����