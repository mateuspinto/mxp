��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���>`��tvM21\3�f5���d��(���ו4�q8".��<�/\K��z�EZ�M*���*u��mm�	��Ew��!����r,/*`���a��ϵ�Ǒ�lAqt.l��^ܩ�M(=m/
��H@OG=�.�Ǜ�Y�C#�����W:���Z��ˬ�r�8�<��F���}G����\%%�r��Ůe}�2T���I�/|Td�Z�{$UMW�E�[�U>�$��׻��kc<�L-��#e�z��U!�Qw�~�Y���>3At�<1|�#Y;���Vje�1�n���*�ڣif�~��~8�?���N�(�4���&�A鍵���7���A��/aq,�#u\-�|��
�rՂO�Dj_��e�D���*5�aw旧@������ fs�<�j[Wc���\ߐ5UBڌ|��qm���Dsxm2����"�/�`�.��ͱ�ew�bFְ�\5���&�id���c� x/���س 	E��U,ד :��2=̠|٣�и�zw�F0;ǎ2qW~ ?h,�Q�#-V���r��� �׺��g�yPǯuE�3[��c&
� ���vA�g��ֿ���H	�����Z��trRÇ�uu.�eYNe�6��>X�K49>�j�IbiȽ�SH��H�yc����hI����+�ǼۂpXo��l/mGF�^�bE�	�).�N3&����ߪE2kCZ:{��Lޖo7^U��N;�c�qm�r���<�d������9X�5����B�Ќ����<@�� � ��wH�/b���]�"3�'+(0����Dd�`-y�!�=t\\?��>_��.d�H o*�e�r	�Ok�� �ʢ�>�G�6��(H8\큔�m0m���g}2}J�P>��}�<��=<��3<�k���ު�|���K�F��%�逰��s;g��k:��IKi���G\��-dM�������[����?!�����|��sS�F���51
z_B���:�	�yϖ�E-;B����}�����K7�鿒� bD��z�Q����r.�P�o�x.H��_����wA���%5w����u�Ґ����1h�B�eL��[��0p02�/%ʰ�n����5	%��ک$�*�m�A��6ޢ�)�nxT�nJ8�ǫ܄`L��~�]Y��Y�hq�U|��� y�S����т�Om�琺��G�T%x����"�$�tg�9���b�5,$�S�$s@<�"<'����3�{��֩�R����fF'��u��=b��b�N��4@��ժ������z����5��%Z�e�T�A �.��dհ�re-xr�ӈZ۲Qh���63�\w�*�O؜����Ѷ#i.�����v�=��}7W�
 �+Ī�=��+x�
V(�Mm��Q2Mب��)�����Ψ>��܄ew�