XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��@R���"��3�X���\b���
��m_VL�4��$`ٮ���;�4�1%˧��Y0�1��ju�V��T5sԟ���8�x݆��T�d5])5�(P�������>��z�U9<q���AY;�h�������C�d{��&��z��=X�O���AGw�A_����q�����{�ۿ�ƅ���Q�=ץ�$M��H0�Nu�V㏝�3�)�dҞ9/�D%��@�xT;	,�-9��y�D-(�7�U/g\ �T%�Y8�r�{�z����+�,�Aܾ-L����~���8���@�[�i$,�>G��0�ʴ#�g�T��^@s��3��Ɵ�ϽG�?������zQ��V��vqZW��y�"��C�à�m�\�����I/$���_�|>M�HF�tͩ՛��ڑ�0�v�����#���]rS��"e���.ST����k��;�>��e�n�R/#��n��2W�s��:!'�FNw��@{��.�8$�Wrؓ�'ǰVQ�bO݋I|��q�oԩX3w��e����J�S
6*sFF�7��,�>�5���J��mo4�#���$C�Ոi����5���yT�O�jfև�/1��o5`9��/9�r��x�,m��#�b����a�G��O�����;_ jݎّü�NU<�l�e0;l��.�|��H34�sA���D6ã��z��0+~î�*�;��!ً�]����G�p�&K��y08�"���4�5��V Ղ��r@1�߿��'���(!���-��p�6�XlxVHYEB     400     180gm�'��[�i��2g��'-L����F����ϣ�k'��r����b|��1d{��� �^�1Ô����h��[���
$ !B�'���<G[G^�KH�vD9i*0d���N��-�pS�D�j�^(#��_.�V��	k@Z�3�NF)|�Ն�#��	�E�ƕ-�Զ�
LX6���N��U$�9�ᆴnm��z����J�� Z�r�P����'sÁSm}���F]�?�ܷ�^�s��P�@`��B �� ���	�e�-�Iapߪ$+8JD��U�bg����%v�ZӔ�fX��B*ڤ�0Ç�B&7���>�t��Y2�qmWK��\�㑈����{.���������<T.�����aMӌ,�XlxVHYEB     400     180N\W�p���5�~O�ʱ�U�&��E"#��շQ^xb�Ǵ�
��(Yvv�e��f]|^>�BR�����o����7��7��t9c��鑾��;���� �3����������"u��?�o��k����]D/���e� �v�i$/DIL���q��\d��ӄ�z��0*��X$��i�
�
��)W���h>`��p��A��v,f7���y?y�n��\N�}�!�B��Բ��cdrG�ß�WL�1�eEh)�e�B���|�۠�x��BN�2�m��^��?S�=0-���O�3SO=$7��>��;��bh^�� Q7f�WP����}Me4�O���?��0J��Ke�t��*���p2���a���%�A����L��H�K������{OAXlxVHYEB     400     170����	�@�9z�x�|�'{�P <���3����z,-X��HƔqEᾑ�H�"n��>�>c�������p:�fj �J�	�z���:�1��!��W�k��!5<���&���!�Ɵ�-g�����cs¤�8����?�`��vs��5ڌ�$��7^��� ���<���`����y��Hdʒ¶�;�ퟥ���i��_Z3ں��)F��k�T��m8�i�Ia~�/|n�,'!1��������d��4 ?)V�+hq{�caM� n�L�+!��^��d�%���]��[T,?�Ƴ��-�C�\c�kh�)���!���ī�ˁ���\��5�h%Mc-�	�Y�=ҹ^�n��XXlxVHYEB     2e8     120�PI���p��Tr����&���Z07x��:��, L-�b����;B�b)��~�����ZJf�W:����AD<m�c��Z�#�ӿ�#������.&�Lчȍ1�Rzu�j�)"�A�%��1�g�����D"���F�PU׽,*�!���R��[4����3;��2�nU��㸊jl�a3����b#�5?7�|�^���b�tY�������_��J�z_f9��=���\��eY��%t(}��3,)�.zC�H졧R�f�K8�(�Z-g�%