`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
0USWSUGxovGsyBJteYpEobOPsPHALRTkIVYh4iRGuWWUv0drAXttl0httZ+qJlyqfroXecGJBKtK
oQP3oLkM8WFamCyNIpxsDOUsdgk63BrjjsiBoUxv5ofg+wNO4siS/2CYwoKmFC3V8ENpFYq3odla
O06hU9ae6oZ/7DC50kcmnoot7FiRCm/A4GOCGrXw9jEktsOFIVwbGjB/FB8/XZ8zv5RymVVNPt5Q
M0dI7untjHAM58PnhvEGbEmFyobYVhg8aZhPeIwNWLj9YLWN1YErJE3vXweOVHHuHolr3xz7G0M+
4vuMTaD97GX1A7OsD5Z1c69lg8VIui8yvBT+ZMAyOcgkoBCGT38TdoHtNc/M475iRiJ6I0R2ONl5
3JtTt52exV5BbXC1PS/SUmRFZLpMUG9gRBAwBUnPa7UbArYxgayklAVz3/soEfOSHGcwSJsPJTS6
srpKo1bhBLnJiHa5z90cCO5/4KsIq8e15ZdbDWilE3ZPANWs7+0Sv7hOhXQM8frDhviSAiTKLVjo
HNpXDG0ilRXPtxgEcBMy88pr6GDxcFca+FIOSRgTDMOFDqXfhIp8xsY43hlix0o01GrMeQY1jvQ3
hWzxtfkegZv0BV7q5to0vUZ1O8C+IfcXzaEIaZfKu+rN6lEmLyTVeQslYSPvXCimFLP/Lc5HDJUL
FXKMWSc+ePHSF2KUur+9zZFNNfmF8ylhp38ut0VgZPrcHyVweUvY/K7e35sQGEcghaX3o/K/LxJN
XwikT8I09hvZkWPUAYcEorEiOSJW8T1k6bhdJb8d50GKHO8aRSgTPwZEdi4V+XRUjcLsbIXMb+uU
TY1ru4JYrpnlHlgFtW/zkIh0vdlDI+hhAoFU/v81kQmxcj5YIatli4UlrrmStCa97Pz1cnjZy4w1
fIHNXikVFAcdkux698aMHyi6/AwhwM7IloispL3FvyS1or+hbH52b5OFVMcYlC0gjw+uPRq3GGkd
Q8fxyw0ypDJ/venwdxulQyd/f6RC/nkSUUza4V/M3eyV6rd9aotQ8n4mmvFVxN79pWFB2RJHYHyM
VMVy3cvAN/kcyMoreYP8OlTa0pxJxgpSC91O7WgW1upJ09wDLu/soPwvc/94o9QiWWGVuL+YdJxU
BYrb9H9M+8nG2ukjRRcZM3j54Aa9oHc24Jkzu11r0GyRzAm7Djk2hYg2OyEH5CDqT7BgOhJujnET
b7XJAN+tMPAk+tH1xYveAzkAoGT5YnoffVqMZcolq4DXLiaLdbTbT/bppHdmTbZaDPvr2RPpCBmZ
Vi4B4GR5bqiQaDYmsi1LLZGdFcN9a3A/jRRt82GYZYZ5VynHt8VjJajOKoOtBEITW5Ps00r4TAsR
R0towmkYsfADntwbuLKaod2IBAPeDnecfp78aK+gehofOjMrLF8/FCqEXNuICYyuownOliarjY3z
3w03RV1NhKKi4aTu8OqVcPQMZYqXfRT3JUKI4dXtAtlW9D2xyCuar+lVwN+cIGtqKrEfNl9fVAPj
UdDO0PsklNGq9qeU+en8SU7XkM43dN0l9IB0GscVM7VPOuUXvbul5cH+VTvwZBU6+Mw8Oa6Lb/iI
TsOrHlEPx2TKlGpJ2oD/EkwYAg8XMg1cKmrrpt8HHIBMQItXKjVrrHEyNTIbyzEu9BCxS1zuKiOf
RLTESUwQ8XO7UAa0QH2eVfowYfpNBDgF0oUtkCoB+Qmytaw/JH//X8V+BZirVX3BSY8l86UZj8sY
uhDdWnMSOsHqxl/aIy3vxle09EPw99R9411+4HE6MrqMtE/htstukVlHcnEh3bD7nveMzChqCNaQ
BJ86Tkm8I8nLBZYMWzDheHmJEnDoS2W8E9ocBdqqdVt7+pF85Rqgr5JQV20OWz6Xtpf62+Evo8Tg
2scF6H6pzUF+5/jSE/SdjDc6dfrZ9W/VCsCfk9/lqyjET2nu8XPm6d9yRtMXKOLZ4QxVBzO6OuCh
JOB+UfK9w0YpFeO/KDyvZH0i5b34aUhqJgCESxnH+pY8ECjbtTueRnzcpGt9O2YHzGYwfKB+IARV
zGH0QahmW4hBnlH402vWLfD4hclBI8yGNVUxskGglhdIb6FjsSfeXK/5mXWF
`protect end_protected
