`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
k7iOFCkgUuIFK5j0J9CQKNbl4M8aHANORXclFkscrhctS4RxxpYcHP7UWi4cFGVXucvIobvz+C0w
DC6mYGQUNzw+jDg82/Wk4NVJgtrQTPoA7bFfs1OiWSQ3+NxBK16FCTKvjF9fsQNRPVrR6FkHU7Ji
oWktuMNWnivR+A4231NetxB3brxtiIcDJ2jlMwghvrVAi/RFibV2Bu8gYwNoYnNlzc6NpCBsYs6N
RUMrwiuqc3UwfjtYwOpXXun3Kjq8eQewWSjSkCOyTuBv1jQMnPRkwBfq47qPcehHf5zVXpylLqWm
p+iGOaFn+XdVVS057kDhuQ0pBPb27louV3K7kw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="OAFZZ+AIDb1/EZ8q4Y5SHhQJCEE2iJKRUnFxL4M+c/c="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 49152)
`protect data_block
elWJOujVcZGBsJdkq+J+NzeSUgPI/1DC4s3Xc3Nx4ZiuQm7rGadRvJR8q1qnxaj6sCkXREGYNVIY
t4vgsCDD6VgtwL4e3YOSItYqY5n/2BnenzP5//Wd2ublr0nCtsXykI7UYRi8ftS9AGFw1SBB/qzz
RlWUbXiO9psGDvjenmr0v4KZ0aBxmMD1SqAQgfK9sElpVR6g6JHHOcIDah2lT8DTfVy0BxjYBJZI
msQ0frU63fkx1btKbqZ+PUpstQrRLeEObtnxjQ10ugrqzWT9iOQ/oz7rwyhmkVQze1vjI9xDR788
OKAotnz9tm5E1HJGWI+2MQfFbPXRo2TvAWl4z0IbnhXGf1s8TKX2V7+lKbS4esqLGSq1nIlSDLdC
q94IXXldzzRnGYcZFGZ9FrxE9B6tgNPyWmRn4GWTB9JCABtjReZTeoFK1v5k6hIUAkwv8xFFiVoX
0rM7yUc9BoHfqcbnx9zizJ6ToqLnTrdXENliC1SRKiL58m0N+6D5SD8HVT5WghUILzVbFQPOVN7o
mCPeSdDy9lk3UlZNOzjtnfkwj7CV1zzBz0Yt0TM7t83LSLJ3x9vhkhVV820qeXlEZRLiCBx/Lc+/
6lpnvrPBVW7WxH25WtGHw4BbQGvQxFTFy3IG5qAL5UroZK3vQT5HC+uITheoVbqX/HYWc6jggm3n
7X/+11xiJB8cBjCMI2UJFGzp7bzl9bk9kgguyMnBYF4ksc1S4ol4q+A8qpDATh/eznD6Cb3UbEXp
NBQS64s/uUJlASBDtQeI6jDQdA8Mj5h/gz1X+Ly6n1EcLO61Lu6E+rZEfm9rij2Q+512vSZKJCs5
4BxJQMNpKvlWhdm6VSggHiMkLHgdOyOVuZY4h3nI+qQGPzP6RMROwCB8Pb17sCmyKZQVodVjEksu
KQ/JWgwq+TzimMREfgv4iPff0GNIYu6hhASPE6ZDIEfCCqbDtte2Z/a5HEaAKV2soIFE64r30rBF
AnfOVrXX7OtiBfYFACSEK6oODV1AmaGTAzVtB2WMZTwh/Fl0TM3EM4FqpzF0ZcJaUlX6p2gPQ/Hp
fjCQUQfNqvMyU9wqtJdLUL+q4ekEHgPwwlfEQEVkdyibB0VmeIMnm4eIMBM5TfCAVnkVQkQQghBm
WiDpPLEqy5XxRyA2hP4+hduMFlstS0Vd4/KDuZGGAjp5eSaZblIi10msAwLY1QMan/3GQ/C+M+i3
qz7EL0wndqHePLAmPrJ+npJDhrG4wHB2o9M1zIam2p8fwZkoAuQFGRx4SnCszyIzqpfptBsAi/Oo
468IMdwJ3HFe/0Dn3Ll3dHAs1U1TfRb7tpNXvNgHWK3vrIQYeJkJVknKTZvubfUhbUvZR5nm6V6i
wLzOcgQ9j9/XxfkJqiuQujzWuDMxckOo6al7o7ZJwhR794/RHN7wp4PeajXx5kEXJywWkDiBuI42
bZxXV2djgwq/757ezNQ22opitlsSd5Ecu3RQAMbTgG35hTFIb+hu/+pw/da0BXVkhU9h7IF4KL0C
Z2AfOP2krvPLrhR7QPAfuCFv8vaYHSFjJ1e75xPItu8hM1FZOEJ6wDAWKGlG5Aj9L969hMU0IBnz
v2SDRckSfSJsmEmqy7LfYQYcnawwls4w7hVzt7kT/TRQe6J0FEPqLI0rpDjC8u0qhpl3dlLFUGDJ
nYv9Vipqdk/w45AXFQoXMhhKlwxAiZo8Kw7E9P0XQGoPDF3RDOxIQlB+LTWTebhqgBvY9lW8QUKM
A5Zk4UQU+aNqfmJUu1DEBQ+S2b9kw7jYLaPmC1bToGseSvD0qA8BAqCke+PRhrTuUbJ5/8KqRPX6
x7dJObx1fVUHSPcWYZBXrbDiJLHDWbUvwYImIY7lBqRbYjRhJY8D45Xv6z4FAt0XPTQ0bY008rNA
t2JuSKxTFedmqmctOD76uIrwLmn34KS1l0Qll4a97YsJeujUjHelO7poJ3TBK83c9GCf46Qw/ezp
o3gkFyGRuitZ/dp6oBa/UqbVtn+i3yOdTkbcRGBC0hfNPokNamft31QpM24jShw7ALMeHbFAojWq
u2dTQq1EiP8RogpsoERsl0nNRVThbayCKNCM1iXRYr5SBcqdoPC2XxqciK9Il5Zl+KyKSqsmjMxz
lFKtD5ueInEQUA29T9MZCrgSU1Ptf37BN4raMUrEVNlocJuvYl45Up7d4S6B3VyUKqAGsSbSb0sj
6tZTz8hp/9O8tLhiZBcAnHWrMchunPRNbGInbTBG/5AqX9+mZqQvfol1RrzpFYXscXorL3lbBACF
RGBbcjBqpu6pFAITZFwqUl8vyuB3l1GGhRTZ5pQcuIdMznnwsGhKQHG1KrUrCcPpgF1mElGZI7UM
xikIwG1BJd0/MUmUIZyOemuL7uiXrnfw6Y7pSrY5Bs+E6c/dsPuMYAjtJ7FCAKUS3CEbZV2zFhNt
KUvzNvmKLu2SEZW2rIYtRNLzyU8ekU7CsAVdBfV/zXMM3NozI5kxP5qp+Yu0bUKeYh/IlpQ7o969
Fi9lyVzus7m5QKPq0P2IdxyDRT1Uu6s0/zahD3SPUucLNUWD3FQtw/QlfjykHzaQVUZ50akxEckG
da9V7ndA9hgPHYKZFOh7sLUJDR3AtHpUE8uzfeaTmz/qwxD4oUmor2wq0prVPjjGwdI2vpD/yj7L
PL+xyhZNWtFGv3WNuETx+AfRJBdjbMXVvlrvjak8+bRTOtkXDabq6Ilmu9P5JD/f5W6z6X8Lpfqw
gVFZow9taAioznCNcYJWmwRkqLxOG3yDr6POuvLIHyu9yHZtVfZbJXFsLXfrwnfsLmWcql6XkiMR
mUNNo7x895pthy2AKD19QaLan2raHmNCd1mxfxq7NMhx1gaDEZAgeSPp5A5nRMr98PuaH/FCmVQa
8UDOAnElJ1sTmxbMg5STyvZhL6YC2RaV1t+9CdlU0GbK7LUiZiBb32XmRid/+nH1I4kVA9h55lRS
QoXKwIkz7o9evkaAC1gxHBjyv9bWLeY1kd/uxoPR4zEMsneCGL+f2pd2B0QU64HlhIXUWjfLjixg
xLHaLbvtUoy5jGYLbsBdXcQce90TxswSpUlAYXGCIVDwzAuMarKCc2h8uHsmUnBgZNvmUokCZ5WV
OjGhw8S+3CHGQVM4z9o4MDLhRvAf0Q9IQxbp7ZxCf7lpy8zkO1JYWc6wLOWRnSs3tov8V1BBZ+Nv
ycdsjPgaiYTILfYsmke728HxgII700K4X9elcBLov4wTt4f/nkBR/Y8XVW/7Gx6hAxwVjiYfsEfi
ap/TKKsoaULEO1DnRRSLImLN1qgInuNza+8x0eO+SJT28MJcpsHyZ1JNB1SdHjqp3+l7Bw+3tuyL
ttYIiXvbayHGYnyzriZtLcoB0JLgo/GkvbBEbgDMqLHcRIAMFG/jazQQjyCco/I1F1sDragUwnaU
JtYwpdwJzaMRE1U3w3apKd8aTenIyOp9986MeG3FWymOmCXIO0Pd/IyVRvqo8jJ6lhjSR9fA3h3x
FDUlKcDhFGhmDo/V1I3+XDewG/0kJdxL57sDmLXjHskor+nCGtIKj1jHXjBTWMCdcgfBtMQhmNxl
rYqPovMdkLPxo+GV+qBjvLTP1drkoia89gT7D2uPJ4+0uAdhwzWAZiL5W/CfgUJrgalMvoER/zY+
XDC3JGXBg7dyYlho0gE0jtUEhuoXnTv1EfbEN12jXXSR4TUt0JoiXTojYxAYtDJxZoExsOGDUhGX
J+2oX4YItrpy0eiwxHxEVR4JmOkZU31UrKqLuxpJL4TjaTdgPFIs1xWb6DH3h9bt9EcxqPR4j+Kg
rIW3VnsLaBZz/lr5UdYuJw6ZBXOA4vlz7BpNrJbSOw9THA4uI0u2TTBIFz+bGv+coOJeqVq4ZL0G
5VEfascr0rcCJf706EfcL0KoIWCl8lJ0cc2G1SFIlfhOstK/fpKejdx9hs2FQO6Dum6vpl1YKxeB
YLjfIxpSf/vFUysZW3yCj5KavUH/Dm6y3VUxCnmLQyNHATTYcZ8II3OogyXe+qHtCEPuqSW6sS2g
5TRMdfptjUKo/MyZOwg8GzP6IsrFKchAvjNtdwvj9JPODk01ofJL3eHVQkJHgzHqu0C/DpK2FRcg
F2r4zbA55nxfgzgf1vfV+P2RablcOH4J+CwLQLHpikf5TnF4/iQDLF+owcO6DTEj1KIjch2FbSAM
kVg76/meGxYfjPMjesQhPgO+mBTMi1MLDyXCirF7NOXTL4erEkMZOGI6Dxwi0mp2QtLF775Q0sKl
9Oqa15TAhWgz8REF9Q7i5DxiP5QoPHGZz1cdRsloEpHoMHhH1403wi9GwC6MEIIVaEYcFpKL44Hi
32I5HelQXpkRpwJ/pZIQVW96nv9n/aYsdITYvgB5lz3oPHZnrynMQrEegt1KFjvlLzcoVp1fpj62
AbXS2d0TZ/nC0dBDDnL8FQYxqFiOJVKB331c/rWRsLh9L6Dyn8xscW7QxsC0+uRZNROwadXKvmP4
c93icBTwXwR6CGz/Q9V0+OuquaSS2IP9YWD+HI/vvvq0Ma5DUTWN8F27vu9xWnRaWFCSSv265uKz
dYQNcyqKFeeF53PSDnrm+bgTlAWrL24+K2HbYJAsPgo+3tyV2HSRORMaBJoJg2Dvd/zCuifI4QWh
qYmogkYVR6AY07Vyo6bE+bcCuRlXO1U2JEWts5QtXYnj6c1zeN/ne68kNFm3HYjYCbRgfsTKAiBw
STKqwXOvGhftIgKuzJn8LXiVjpefao7sJuxl340/d4y+5JTmdwwzr16D12C3Iy83Ru1djAT0GXzC
9s0cBwOmZwidH2aIl3DBwcfXsC8E2sqJHUK8MSHl3P0PxRA85KSBzVFt/wNHyCp//EFb2ixvA4F5
tq2fH9fH4d7n2dEOd5T52m3cLI+ckSUV0zPukEKyfFtzS0wKWI+M5FvfMQjo7oc09kWTRuJm7gxs
HS/8ghj5bHD7sKUTG+oaz0wcRIetnZq5SAGnZmB09moxokAoyoPjAlDLg90c4kvRlfI9miOmYuDs
p8rLfAdGhGsUW3bgEo+ckZXssLHmzFGoMv8/99HcQF3Dd5uD6FAzZ2d6pk+bzZIAT5iv9O9uJ5Fj
r4MDHTTIjdavbjAEx/kRxpO/0nCK98po7FC5ZepdzI47iE6/kdTj5n95mkkHL0SnRHN7ieknSJni
ofEcJ4W/F1fRJA8nFAEbX46Bo90Y6n1Gkee/yeAWbrmt6KN7C462L3ryVqt6PwzX1eHsXoBNwoIJ
Qh6oG13PRfRc+m4ciCsSyuxhlBQrcJlLtfUgVth2YRnteNjX9kKe9GodiXQIUKnsjMtY4MHTGU1k
VJ6IHPcLe/vp8oExFpGhNURUZJz0NkkG8QRINYHS/WUzIVujPtMELAGVDTvpBXLBmoyWNPuEXjNA
Xj9213gUO1U0G/m9bZDWphHK7BLHu7c08Kn7BFg6Zfo2JppOHMVkbg54aacW17b7WPW1+Wy9bWWJ
CQI/N6nM5ecJne3gHmqSE6eZiKCdimYLcs2LN8VYiZ6Wyro8sXbabHvG17VWzI1N4Zzmu4xsPmDb
BpcuSsJE9ADsBFp8zR79SfTLbUPd5RV1bKrmwZdD8vWYyyvhNE6o36gs6PcPzKOJYPcr+/HliBNS
PknsDpOU3lD0f8AVLOrMegfHEGDX9Kn+E94eIkCAF9Klk4kBsS1upV8PtQVwxwFHtaE3Rnq5wiH+
iErAC3Kt1UP01vo/6p3GM9QVpeYpEZHtuhXVH1vX4hIQcrOehXoubY0E6bPl8ExabvXdzlWYj2aK
SzPqZpQJgwiqhVlJ9eHG+Aq8HwXTYjMrYyfX6wMj0JNVuJ5I34i9VQrcpYpZcaHkfTYMKk5tCBDH
D1NYoDNtHt3OKwmseQ1Wuuo6Vq9jfjN9pi+A+7w4U09fBrnvplJ6WMKX3yCXPpmhOr4S6kKQTfB6
HX3poMLSQOYt6cFUGDoNnzJsRE7Q9v/Bzn27dR4nPQ1aHrGLXvhaL1GQAVrLD2pprTLZDC9jH2BR
b5Oo1a/JefHISJoK0KBbydEQQ0CtcDEa1wM4wSLCpEUqxV/MIoNAXrV8ihGyqPqCIGJAs0evtd7k
/rffJxTZwhGhIBod/26nBWxN4EcIg0R/Qlg7i1rpj9G0NCJavmjDAahWtmk3+ymx+ODAR3vPj7Jt
AH1fX+BeFbKRTUWZG6cxD9MGVV0v2SFc7QUYDZLyAaP1hyy/S/oPhPAAPmuq+45IEewbV+KvdkWe
v43pYTpY4PAX6CKLZaLB/sz5L97NErxXtN+8NFi7QapCGRhZTs8oTHQRx6VLs1NvStBz/uxSkDg5
mEqMFiz8OPo0QhxguZSxnj0npI08zLwmCegKDi3wCWShvqGr2EGMrFgty64jHXOb+RHg7jGfKaoH
X0M8xdSmmdtclETXE4kAZUQRkyV+GeRMDiNl0eT7xYn7CrZqpp1tVByrKQ2iqGtyRh0iTw5rZV53
6YpeBWq1QDGPFAHM/mYoLa8iACQOqNuOqoXsyXJiqKQWo1cr8j7KEMqNOjU+K5PRV7UbLPBlBSwS
0Ie1v5uvaoftPF+4ozHzM94W+UBhk2m1gZ3h9RCkRn55xmTw9Qjcuj3CNRqEwYunsmBia//fM6nQ
3egy3iq78kjpVI5jcMssvTVjwdKELilWp02m6ndOstZYwqrDyaqDQTftpTQTgKdSpec8ofIrPkmd
lJ9wLEZxNe7OqvWuJS0e5sm5watiym9GBJPvrmeELhs/0Kbt+G7CNTCzY550jmIiWpRKIjqmxwBM
ZJXGMJgRmw+//SihcCILB/7vWC2friB9fTSqw5QhkybQVxgCV45jtvZBd1aR1uXFiHgcke11SLgL
O5t77Yq0JCXQgeh84LBVCBLDuyZFsw+DWe/OZISM7NBr8zTSCaBhuLtxulV5m0nkIPyNRGYCJtiH
W/LJL8eMtLSHEeWNDJQneot+KtnU55ebyuzEL8R51ZddyV8l3kt0CFUQIthxglhEIT+OeR0+2U0g
89Pg86s+1YVleBOHgjo7NpwaqlUR8wa0+t9shSwNDBPOanaqvXpuT9CsvvbfZLav1gI7uJaM5kad
xUQr8VM42Rv10xOeoSf9X+43cHNGAhQv0Hvy2M4j+u6T3XgC/OXdtjIrhFxYlVuVBYeu9i/ZeVfW
oiHIQ06DUNer3pX2z5yUz4B59ebz3oQHjw3Q5vJZYKYUZMgm+tjCDKyES+rhQPbZM+uH5D37DGkU
OnR2Xf56yfxv9/lpMR4hzBZdcBJLf+LkyVmjKWfKTI0J/jzlvdJiSfH3po6rChawbQkZq4mtjfdN
vrZELDZ33sn1m2cvUL+ZtRTc4mM7VBdCynH0zXqWBgkH/XKcu+OQRYmXx4W9k3vCQbg85J9aJY+B
oZm9TlTKinlkBFz2JWYPbO/51BEptPPblfvIJ1tzLG5vSOU5i3DJiXgUZ5ZVHudBkXJHeBO+v0R0
BrnQmnxTLWJUyrCrqEyWXlqYs6v21b3WJX8p9mN9kw1/QfOS2DbZqCxqZE+TDUybbpq5FVaOwVr3
bqFFljsGH1V39VRVlFjL0p+muGV3IcphM+3AYoCQeMy9CnN7lSqyNfbNY+nd0AmGVH0fIsPRba7t
xyzal3sfUnWm2M+iuaDTXgYefS1kLFsP7sX82rLU7TY3Ok9+l3juaN0cjTTKkyJ7g9kQYZ5bFi84
ojW0tHeqWA7m9d++COWvouTe8mYwGFmZPdJCtk+Gek+wr6L4nLfkYyyw1ShCN1B+whBI0wcFW4Qd
XK4ehdvuFZTn5BGjs2mEUyQtMiFNd5AyQmS2RfvyKZLA+eY4akDPmFoo2hnHOXUVGl58+RmZrXPl
KM+HMVasEqInzzLcg5R61mQUnmeY338A5DhmGw3F2xNLCLlEXR4+xlN7cYT9RHVX97/uR3vwdCTL
XPWt1VpvU/T6OuYp8jV4yDB0Vei4aUavr9X30c7alMbb5DwMpUtqR4/10r5+5Hyz+8pxL3taQJqR
MCtDtTT8kH1OLNhjki82VVphL5kz5qHzkM5JxHxBvO0oClcQXSD8D21TXTYFU4PgfoWSbiWVEDKd
C2xroKocuyuyaQmyhbq1rJsCRVl3gS3Qv6FUhTUOVjlSTwbfBn0DXUPXhn95FJi3U+r02aekmaK2
cNUZeC+XvJWyQcDNoK6KxMFPvY1t2cYPGuL6rTpApH0l4hb4mgoHy54VGYTdz0ozv4d3hmvBBQIO
iO+sjfztUXqze33nqW4umOsDAk55BTfhQ3vIKGBLm1SL9Fv/Q6RgJQIdPtqdMWDVQnlimaJyJfWn
+Q99SlGp4SR8/xjDmuTnGUJifoCytTdsNb8ittzAValqmKEfqcdfmiLHmmvKEpPPZnJ0TBRcB/rZ
Ear37tlGRNJ85EHh+h2UVcyeqIN88Mb6u12Z+seoLX71SPAPUzobtnTbKHQYlti7nn55L+LFfaLP
k7QTmG4Wk53QKia/xiszGJZsvypvsxzjWAtaJm8zc5+tzGn3N8ncVLXUlgryhBOMYWhIB0QOeGrl
rsqNJcAj7T8PuAqBidHcX8ch0Y4ZoTPhXx8xQBV2J9j/7xbF9zZKqmlEoGAijPkkkX7SVxzao2Ps
47zTO4cUDx3GJTk/35yhAgzJWbYsBcXQdvMZmiPWtqc22ib+8D6AyB1Q7XhOsLnW3Afw/HJsx70s
9P2bGpatpZqXqx7Wi1nbv/VQfZ5q2sPmEbXbiMvzuoLNgTYXKhAOT+l9MZhYus2LvhvUui1vBcSW
zJNvmRTBCXPMehlXiv23F1Z+BfJJuCY40ItEvQZz3Ma5SYIjnPzcbIgydJP4tKF6390Y3+kvph7N
bZbHKnKAqZFHbB7eQ2BegraRJlHdFi9Di0Yw37DbZX4CqIQXLkaDaVCrmuUrBGN0SS27iDWaBdpY
mVhN53PBgXKiCjS2bD3CUx0qjv8LnvP10+WOOD0UMqfZhp4sjFk8dGKLPjq/6r8+KHZy40LktNWq
N22Yif6tet8wF8U15Wnpd4NgxhDXCu8Twfa5U42k+4hAyCaXnhH8X0azGJgNkaZew+m3BnwZ5vfC
avd/xUnfqqUxGWSAp2WCqY7KaKW7sEtpSmY+gtckeT7xAqswAHyskPH6LRcf/k65TOTqAvFWUS+R
8eGANd9TqNOjFvnji8c2dEVSWR/3OmcUsqLXh0EAlxqKq+9S7rx28L43LUWZ+sEidbXVrCmx3qGo
rrs0DdV2Zye00zs/fYsRRz5VE4uqfhFyX0cdDcMFiqUjwoqqh6tCQGBxAi1oycc7YSJxil1FTAY4
v10jbdN3nr+/8dNmqIjy2bqA2wATr9EIhESGaBp8SXatITupz4U8oqWMEZMcB0QcqjZJ27dzB/CL
FHU+TN8gaCSQM7dpJfcJ2hUB+trgA6EJCvqJJgGezuvoxpoDICPvyp0ky3DrNtoMJxZORwKWo8KZ
yV9RUVXIROBqolH+0q17YLoR6Gu+rZBhnfdJ8oyHZpKJb6O8yjsLCbf3I7Q9uaP7pdOyzAzeZlnX
OnhtErriaUcztYOQilAAZ1XEuDTrjV51batiiQFLZ3jP1BslOyodoSQlGHc9vcW80arWW1XT45uw
aEyTyCmkP/2EGAZswQBcXOHLBhBZlEEF0iyz5LqvUFWmqRJcZXAEofG49FD6C2wrBQIRyejXqUJl
vuGROCX+9HpqtLhok3X1WPlGPF16bxU9FnN2FEjoEMIr82iWLACvV2rNAgXe8TrSQrrJXXsZRk41
GHLLdwMcNn58ymnqOCvt0oOKWbtpfaHgO1Cfxo/zBDM1FHi3U4maYreybKAxs9LZdUiwk2KvwGbI
DwL46726VOnLb7xDrraf8Zss0hWzN5SnOcXoWix6WvdvUQg1uFa18HCX5qQC+gFdOvOz0R4nMTs5
TBEirjelN65cbiYOLEgzre3UzmVQ4wf5YQJcFxiW9O8KwMUXmoSp+p1tf4QhXNzI/ZA7hnXPMO+3
+gAR6FKPFPS/dHxW0/Atppx8lJLe2RAj9WpRMMC7/zMksJNza1bVT6sVPXW7ya+4qPDKBRA/gsiA
abARlugoSugLAywJUd5lq4mbbkOQ2yPom4HZoss8c1rRTIHUHL0sIfkjEE0pbW8+TvyKuIUZZd/k
mkkecmIkfdOM5lUP/MjDW7JV+7aJOAP5Gb5FwB2DWwxaSrunfYDJpiMURXrY5RC2X62LK5P58bOF
VlATy7bkPy8ZWNuKIrOega6IyyU96/RRszeOsDmKbUz/kcnteE74msMZrvc+EBZSPgauwp6Vi7dr
J1/W+FNetRsV7thVeO8uZZy9Sx3dY6l9JB59su0rrw+9v595s6UpWOTn6hEMS1KWEe+EoiBeWdhM
KBfvIDxuhQ/Oywe7Xd1fdDZniJn1CEboxCQ1eaQc0aulqxMaX+rJwHysLtRQ0P+Mu8l/Uq/jor9V
5+ipmbp1gbGihjB6V+zo8KwK7JOQYht31mGQfcc1lvtuqhAfUbG3TDjWnudXnfr2leEbR0EvP5HM
v/wg8Iezk4/DOioeCybUiD3EdzhPho6FvfL1xXuBCCJtwovJc7Ogqcn+wm0ddXYjD3QmPUPnydkV
dm0SkWFqbLlSux9QltbYLL2viNno+6iYVD0gAxTuhwgOCODVM4i4apSjlCXJvZtfHstZjP/sRiKP
bmqAZNiE/mE5WgCXNkFJyr5CezNMTj/BcyxYA6lcYPoLta3m0vBRLJHOxKAE1l4FLEkHb9Zx6rrs
4tl7MJv6JUU5HAyilva2IUSVbr5GdZGrKm//g7K8LHtrpUHTVusV3tV181JfNtWh0FMXup53upjc
/x5z51fLnJpyrLlxNmzIf4F82mSZ2i36I8igO3x38gCyuATg0IKxzlko6rkAu8M8Xl/IddwxbJ0M
GCV0jfr6OK6rxiz40vcBROPBLp91O78TnrL3WcaJr3gfzwdd64tyOa2qQvReOEjBgMhbdwUOvCrl
PPnlfy3o+uPcdTH5LGeT5Fz8WeH64SWwfF/5I+ZlElx8d3qQdyz7+Fqg3Mhk2eSLlDbN9jq/lRas
Bm9xFpqNFUfE7vxCnkBZISQ2R3fNatVsvq0mghk2Wm3KjgdZ8n3lu44f7ZMtEgJpoIpkU8llsgfk
P8uJsfZjW90SOZitXVeUnSh1yUflC5qDRuGtoaagWkl10nVh5n92h4+dS4doGMVjOQvsGZx7ClvQ
JKz2C85vBnypwbJMfir6OMOjD4VRtQ/vNJ/nLlFu9l4QC7Dr4mLBjNynLUGFGfyWxgKisIgrigvR
XqqGQvFXgdvJH8gpHMMZRqCc4RaWjeVyZcBu9SBhYg6IdIiTdSGb4qyQjufaPxrVeeu5iNF4Sbp8
2Bku093wvuWo2JINaPRSQN+IiLYRR8WSTg4xcD5tRKM3Ooo9upBWuKEpvXyaXRw6uIu0/8QP/5Y3
aq/voonxZcLi8uZRRaGsLc2GzVCn9XgJ40dddmmBWptV+qVW07ZLbS5nv6XgqWZJvTZVwMqMBLz/
CjAtEn+e9qHbCCTUXp47mQtdE+2xcJhowpuSQl/ktL0y/civfsVMJvk1LK2j6NbTIYUi/G9Ge8Fo
Whfn4qScK39Shyk7sjR3hnScAaPJLwfr5DBtLl/I7K8Wnp6tx75r7AyImxgNjdB9dx4BQtHxcBlw
CBdfc5Uyn0AXIqrOWpfgEjCXon8l9ah96DRpUHH0c81vUglJrQjHPAWW1XFZEh0J7u/bwyNk34iE
vNYBxSjOnuuPeFW0k5j5coAj8zHeuiAKGI0dS/r0i0dtoh8EdYGABuuBHGrLrManYR4CwOB02Ha+
cbgNzKagGblB25UBV4diI9wf0MR0lRV5GUZ9bpZFH27t4M2pVuVg0iQf+HpSpqDV2YYMviH3irIF
vUzs2XGpSYbl1RLLYUuj41qpSILQQoVzdzoWfyirkL9BbTwB1UXMIbqg4aHcvos9zKvtBrgTTyGX
3Gt/0vSHaTLVZC9le02FMGNa+7JE45+ConXkAAoHCREfgH9T/bAgz9Ec8orxdCxZf07mTJ1hRHCq
W4AsRk1lf2ckmgRTdcxZTQ7+J+q+27ivI59eh1tz5HyXUL1ZqtEBaTkSn0VPCO3bLEWiapSVNcBJ
Y8QuY7wU4srV5vFa7Ap3PhM5E0e32b4ZLsXwO0EBclGB0p3Nn8sgMMnuwTKqge3PHtJsCk2ZCh9J
xVpjrfV4qwXNDtapcXeN2x3BI5LqDzVk+7bwo8OyxAhNflRMm7oYYsVfaPYqH4bBmbqDj4jCOT4k
1fBFgWsNIh5OmY9Cvt/bMYiO2bHKhNOrj3Be6QZ0F+OR0jOJgTfCk/BjtN0xq85JT0kfymuLqXX7
9aw1tK5g3jHWfrz2o4ROQw5NURCWxoa/uqXcElM91PwW3bhwfzSwQPbIRuhBfXa7ZfBlIuH+p0ds
Oi9VjKEU/JWPa+Bd+wZ8FHnMGv8xQ6elEFuD3ys5X602nDysHK+7DPaxiqj4Udjjc6XcqWRwxT71
5mF5qu6enpiinOnGs30QtOwCkMWiBqmEI/wHL+Rk/QdxrGuzJaXBoaD1u7T151vCUnnkJBoes4/0
k2GbNVu/LCM0TWLWlW7STKw9P4Gzm1GVuhPga6jP8LZwfUTmThRDdJxw1lhh8YRJ2i7gFXmk2ksW
nIbJGvEWWc+/6aLe9Lqe2zCxMThqPqTmtTnCTRkoHGJlAsdync44UERVxoVZsQPSMpeMls1FTHTa
nArTpKSAWJ+CnGEi7k67s/mZvsp+JIEOrQBHTwlYqYbq8D7bElqqd7v29MHoc59lZwOsjUP43dyK
2TuZW4dTzDVhsjV3ZSjy4Dy4fLy5FuJTSclStt+eZKhljpPh+cWWn7zTFt7nTuZkFpQevXqlPyOi
LNdkIWpKVBU8fFMpYmI+vYuuOg7GNKgxjJvHq9zxAalmtDXWta1DIBHB3veM5IeYIFpItX5lIaCE
8YsEUli6pL8DHGI6mVE2kqpJLvJHGauZFjjRyz5dq4mgaiaHE2MygPr0kx/YsHtMIRtSlKrxNLtp
+lMFV6RvKomU5b3de+2LtZnr9M/QsCvtUUX/7JEZyPNLpvHUT0fI+YnYBHq0NEqN3+8o3GGdS6H2
BXulVBIwdS24gs3XwyRsWX0OBhvu3mpJpkpOzu6CVnKjRU9VKjjrc9Y1mz/qYP3Q+7OedQtqmFn7
YnvreyHoRhEjTZNy/yZGnzQ1NZ4eKkweAtrWNlArSdk/1Y4dkpguK/8xCiuzxhVYCGi1ardx2Nrx
M39o6pZqeT3hd+pTXbrizFmllhG6bOVaFl0gJ/tunKD8GmoVPlqCYSmWdcb2P5rSZYwlJyuuColu
kYPGQLbmLRquX5YjhVNkop//UUp/81R2ASLUqyTUDWrYtHqrUnMdgM3T1ZqV9oMNveIUQzzXaTGx
7447Xfy1zBgj8+nqcrTMa9qF+27i0eLQv4wID6YA6U/ofXoxyfc5XsvQMWDv3ACqCpv4vv4fSeCX
4cqwuqV3Hsz6Ka2+Zl6k7T60M5FmyhMzJXzP3KF//Q1NrjvmjNkVHJInQH3Qlf0EHnUGLFgBQrp8
RLW4MCTq/EL1f8csAvjS5BitSk91HCLH6UANeYdGOUp9FWU69Zpr2+IRPF8a4P8zTG6SIBEQAMP/
Q+OpIscsNIIbJ7iSN6EJ62PYEEIYLCrXOCL1LgaYDLNKPgqEUhCKUrTpkXyqZeknEfY7bTI4a41s
B5lTlFgBrlNLCb9h7oCn+O1ZTXLpdkxKy0YaW0JZNKNpNKQqMnTWhxKPrwIO4L21v7dD5Z6VA/eG
T9qFLH7DkVZC2MbdQZh6/U4Fhi1H3cSPe5gWOy5XwpiEZNTbcSbFkjzIwGePXqW4QwAN03kFQSoW
v7Usf52GQm7VdJMqOf2nVD0Y7HADzwgIVTlfhyuhzu+I0b6LAzwY+W5qgbkXzGd3NKn228SriobC
PHHvhR949/YAdmncPVIBp9ioD9TP/nLT7Z8KvuKuVcLHZfIYDmpPu74hQJ6cb3jF/TAKaWmKs49r
iJgrc6wy2wPLmlYE/KyndtfqOG1tZyrKVDF2M9ryC8UFNvkGMsFC61e8IdRRNqVbpiZFoCRQHmtu
/c0OMdGFLNxqw78sJdU/W/65teVjraTFWZ53xjny/+/mxQ+iJ3s3rs+EcpHlFD8yhf7uCCe5BNPg
2UU/Si3WNrF7EaZmHL/CNIGclZUDfbAW5IBiJaDOs0C4v6F6I/dJJ9JeSI4+FyoMMC9uEjrKuXfy
QjdHmpy1leq5hg2xDhRLktYT8rxTxKZmcMwrSHB5wkbQB1+4IKsK021/FPjZteQzobsYfco/Y1DT
maEAKz3B3VuftAZrXwKCToscpEjrPu3ilAH5hZ24yUJUb63p0Tw4zfDUp4P7zEjQhaZ3GUDwd1M4
1XyiwI6MBwPhSIiptvx3f6+TPeF9UVw7j5y9FFYU8AtcqRFI4iet0j0BsSLdQ+sZeizv22dSadMx
v17dg5TQKStxd24JGY5xvFm/712h/ydNyojs70HWBpACLpMuzJ/E/LznDuCPidQ3iWodSWTVNvks
+sQIuW+mJQw7YYFX89z3lEyKrBunnxWLMrhJhITA5jqOsCzW0W4/dltnbKodWJH7lX0HvqAwh9b1
uRc/x9+KIBkwk5KuGzg9Qzem6DUakMDyBC+dMtePvdg0o2ASbgcZOshP/AyurqC5evjKDHihZRzT
1oduVG/2TAqZLOBbjNThsebWgXTKs9umaEanO+qY+nlek/v68RWoKty40C7pnATcvmfpPLjox1TY
gAab9KRFOa5Omat65S6iKRPygQ71I5YVqXcm/8roNTAnIp2lelY1J6cbnBb2pb+zYttEkbYtcVD0
462GzUzh6KsKZso8yHBBoxm7QH/W3YCKl01xFxipVISskVLr9LlF0OsJey8kyQkYIws/Iwu84/iD
ewtff/9QUJaqk0L2odkqnwl3L33DvwjBNVxfE/ia9ZfESv3nQ4dQPKsV0Xby8THTKIE5fv8VVxxv
4iLBZkInn/eCi1TZOlNpdV43C6HtOi3ZH4c//PqXUG+SwtY2ZbTazpb+QmQETFiLg7KWAp3yVSfU
iW39/cTFyLlBI8f60JpF929FpV76YGw4LxpIG2UaT9ai8ByTsNvgJ4gi987h2IMNAjpSQFlAY3bu
UaV8gIp9wAo6aUedE7kCe1S0Gpa0Z0tkFMivObcSBsa/x4/f/VEJGQfqCviXNRTHL6hJjKRrgacA
yQTKqv4Mzf7rGUKnaldbtsMdY1qlPiYIuHqI2Ccr/PPzF8lznquvyphzLUXjoY73Mm4vdw9OFQNd
4V/gR+xncEM3gnc/+twOrESp4qaVRg8oggQ1vBW6AYsyFtS4QMK9NPP3UIlf30/dc0VRXsKAN76y
wOCOwQVZAv/n0OiEZwpzpYrbmIBDv2iu3s6Yw2QGLDk7cDePHVGLxArGrs/7zRKEZy3/3SZM9yuJ
wejSLBpCs9c+85KDvcpv8IFhSCGXo+IkS3lupTAXu5AnUKlRU6sw65elCAT3htYvJDGrzYyW5vuy
m4ru6oTNLzIGnkIoTPJKcZ4HA2n6rANlyXThU37QJ3geL/1qER+synpYgCek3TAxBdq5aG2uwq++
1gsLlOPTuOAnJwQdCfQfcBJ04Y+nGezHAMzhQet6Dti/+zLqZytrBLZY9gjsNAjOgwXt7iavJHf9
L8n1qdbMX9C0UWWyuMxFWzrVj6RYSchDofaRok/l3ewX3rS/cLF8hGlrz/YdVIMvz8vN22crUTJy
yBocCzq4Cbxdv9sd01gCtKfEknAT6saxiRibqmN6r5uf9zX8FRZyhpq/FTtTqmyJgxH83InZ3Kzk
odEXamMQHjQfCPYc8uy+UDt0RueI5shou3NtDn4PHZIbTF1ekReksmqtSy7quYmwqx1pgzuohK2j
UB3e99NLOZJjZeJgqWgz9smlh8eo0BfpphoGv/ijEOxNjJ65UdmrCXdOdHcARip33vbpQjCMMLqW
RRhij51THIoxyVUkICX43PiheLRCT8F76oRWvyCmzmQeNUmphqcl44d0Jbu0YQqAjKT5PRsHixax
GTBlv3dxfrbJ3W+H87UrIWdzn+EKBmbOFimAVUWpGw7Lw7TjtVm9S5dnR9N5Vhwg7R3TEkSC5cjr
evADiJl34pi2kXWW72YSTPB94cc0ks6R3jZlFxUw5oXLnMeJCXzsiiujZLQF8hNJirwbhf2XgFUa
IAWqyZIaGv0spWPgdMhUH3rMdBdlYMqkmpcnBVng1/KrTay6owKYLpXw+nrdTWE8tpY0DFVPPK+j
658yotZKmnOdiuL+jidH9SW2EpZf4nLtzo01+fBOcvr+u73kL4ereuygM87rG1FbdSQ9NE21LSug
Y0iuUJW0yFsxoYcgl52YKrc18W8yOLdlWy2OzoLEosczJJORBTGGIUguJdgV/aHK7wgU0pqIEEyS
xTUxjl09lhwSGyg+5KCUUAZVQjAX8l0ZILCDWpZ3e23GBVRm5vgtfOVJ4G+gDGN8D3VZhtkvcQUs
XTsDX21ku08ph8/OlSifk3a9cfmzKgjjD1U9ZxunpP0PDBSndEOFlSrCcrIENyuT9WQYZyabEHAe
B7WLMtRGwNpfwz6+7AHdMq7itTm0qqN9cw5ijyzljYsR/tX3Ck9YURMThIPaIoul2Xs97b41/j7W
HmmX9uZeGIjNWazSglAhmeVjYoj4MjaTouy35QFxkzOSJwjeJt5+eRuCnF8v3Ilh5i7YA12+MKm9
Mfip8l212gvWcbTIRly50jcEBZZt8wQjgCAdRV4OgBQSCCoqbScR8epaJKvfMRDFu3Dg28Ny8s3z
M8Cpg0p2ssIliAPLf2R51GnYv2vnazQ3RGX75qTuL95qPtX48JjYsuJL833OPcWXzCuCgZvkeJTJ
0wrGcbXd4eAfzBHTGmUrPhvAfzbwy9X+5TqYneZGnkrH9gTXeKc7wX/1jRi56oQvzCdX1pYK3M5r
TdqQhn8AKAp5iCEXERMWA8sS0MaYDEQ0/vMD0G9a2JCHZk1QmHvXTOiVPfmaCTN/BAcQHH8vx3Oj
Fznn2VI72f5575yIaWnI0orJzRLqrMAA+WAj78c+oA2lwPXPdVQ8bzaFgjbW/Kb56DLAcTmdWZR4
1i2P1xOL75gRPA+TSQRmyF76BQusTK8/JJcixpfC2OrZvCoNhyubikR4BunhCpOitLyTYj31X8ep
UlHx3aUWRcXQNBTe4h5CEA4Q1R/wpCr91gfhbRfm6zNAIPBELuk79R6ZPqhhCe3w9vzdMjWaRNZ9
efXAx4LGW2LUw6aomYRlDKmANpeixgP/LvVzy/L2GCA2jFt+B19V6z8i9+Y4nnxdnb3MSp1oWXNK
mG3g9JapOIGBA/0SRhYyRB3fS60ThAD+8kyYAGQ7wDB5u7VRDBm4ToNdpG8MCT2DbDITh7Gy9HZy
hIUlIlcCI3vq2B41P/o8Ib1jTd7k8Wn3n67YUAN/FkDYTPhiKTyzKgFBEcVJeTMw/+BOD1z+E6bG
zAFvYWIsH74/QPl8kbwUDNEgFHMJkAgGWzv1ycuQK5xrLlOvSkNLsHSyz8aLef3Hi4fOYtbCoXVI
dPuRnpp93rcsReEwH73AYOFLod1AFtxj41xMpD6764OKcTIjodXU4YgotjINQ1m2VVBwqmsz+f0x
U+F2wqt9MLJ0BdpMhdOaPNK/Z45s33L2eoeGYZJ066kuI1XZa5YoGMmecsWdi49Zm/dsd8gCog3b
8jMvsRngGnCe2RypG3qMnjCd9P54LFHW/bsp1jgEMFXq4pvb13oDS6eWluAgAbTFFL3alf8TWVuP
BVSatfB55b3lIR9EPJrT+CAzHRp0H5jzN9RzcnNYWQK16WLnxb5JVaQe3nEBep0pmjgo1+nZG0HM
C3KcOlr3BLkM0dHPvSHXn/RQepB7z5/fqfd4J+aSzH+AjEqp+KaW6rHGbknxc7Y9irtac9LEDLez
Uv0piMY6NIBl4Vg2shz3X/yU4sg1aeaz0KKGYC8+hRo89qF0wsF3NsAKCWsqp262C9MmttLKxUSO
TRWfvzks4jSbzrjQjcEsCLl+A1Qmg/1l+fOf8D5tibRFanOJlbb7UdlE29XCWsLQCGPgCwI9+qN/
DIpDUF2UmNdPi0jYgGxMWyoSS393XeYR4RVzC/wrAsn7ac8pEZhzXxjOHe4P07XaBPqOTgcfQ7JL
eiqTIJoVDypyDqXZbuwHEAZ2jKkYC9LNAm+h6x++zzLIzAT8tMQ/tYr8564xcZyqxy+H7QJDoPpD
VUPg9/tlwwX1uyjpt73kHt8puqWUdR+CizEOIwWCQsFfQS/bojWBszMYtYA3n9krwUXlpwNXTm/h
VgKGr42o8KpKw4QCOuuQtb6o5AbNH+SffsCNiOjZ/gB9f+tsvXbSMgodY0hdDCJqNt8ihRkyNTMk
tX2j3um7jQxByh71S3QQPEEo4NGFF+f6NpqiyO4kkEgRAzK4eI/a6qgnVbJz/44AhJUjCnG1FC/u
M9Rn07ZnPrDnZuWpLzIGUrE8/0WKPaW9ktgxcmWgt7Ef6nZoKQpEhBQ2oj+mbJSqNWV3K65jTywY
gfIQQVsGEERYjK6indclwjk82Pp2DOy3/cOC+Uz7BJaPiRkxPliSXTKKEeARBsKrDb0h4TrKoq68
jMlPzB8aheneF0DC57p3zwOECYF9BN+yQdFD67iOPOK4t2Prk/Ckq0uk6xnjJNwHvoYnPoUKDEqk
EMzcRlqeYsSp7dXb1hbsxpggKc8ZDEvQfVtXVqKDSFW3xCzzt7FHL4u4e7fv+cE7srzXLEprKZul
euvT6bFfszGTQTKvJbkWl7fQ+WwVMH2/euZkhQIdZVgQ46ZCu8yielAtthz39WscAdc9/6MYAjjc
/4V/WAmDu7D6R5pTnwRdKMUwWOyjS4T87WATBnPXl7uGlQCuYcc4nD8+/Nod3mwxQzRt+UXKr8Z0
cjphS0t7mH9ukiT0wHV44MBZPay0xR0PXk7uKcQSFmJsKiiwnR+ofL9oY7TQrJJDStfPLi6kAv3c
iYb1pH7o7fLx+7oNLPZrfVRSdZvTXeXXdOPwpfWAELgCR5hBOao/4Wtq0eprdYYg02WX38/tA4XK
E6nmTReHYF4mQfgM8PF0wnPb4L7/W1MROYqS/VY/SNfzeg3iDI9NiOayDD7swJuodaLN663dSOJq
fTtus0eY2UanccU+T09jEU8hUrbxIcBZpCfY0vSWOFQe3eiaWn0il/4OFB3Z8n6Vn1XMctgrOi9C
ZMTL0aBbLzVdDaRUWURragnTKUh6USHPpMoy0KElcsvK8MDnjUXUhNdWqjyBw76HTQHDSl5DOQ9f
K4xjTLh8q9c+jLeeb/rI3Ii+65iDcF9wkoHG8jz32IbD9NMf48aaiNexRujYmjKDYTpKDo3BYdPZ
GdKWsnHRMbU2z+zMMdF+SkFJRVyGm+WL7kIU47RHbn7csqS5d4OE8TGEPl+nSHi0Ha6czS5GmhUu
LJ1rHpvyEMCtsV/to1uGONf/cs17RF54eeOtVW1nyP1EC46Z86ZTidR3FdKJ6j9mI2Vt2Zi87mTS
vhJ5K49AcBvEirzEjwb3fLj2c7SOSPEpmcqW+/q1sRZRtBmzr2lsocqGNlN6dLSvIIFZRaluaSgj
M76f2H80Oi1FO5rCgUL7Jq6KOubVXwIoQUNTQGuHOVnLpE4wbgqbB/WM7if5R9JclDtbYJh4C50d
UGod0vcokc1kl0Tiy865txL5q+em5z1xoMxcsxg1pA6bXMFLULpDxvuancxBtH+GOfVba7dsD36P
f+et4lM+ihMgqCPbm0P69ZUAa2nYXme0gNPVCCag78awL8pSS2VNKyHxH0sozbMvHq7Cdv1w0Ypa
qmYdDshkYqhmHHht43clODNMsn3HKnV3vxcjAy5nUHW+wRyNt+bgL8Gk7KlJr30HxyQ5w0MkH4lL
Z+3WJqyWtBVsT7ID3oCKN0fFPTtTc9+0qAAx/OS4CTxHv0sKRKfaEQgZ9CQsHetxRxMp8TFsjbEC
w8YLhDYXH7vBJMGRUwiO06BnhZCVQr9iW/zUXHbQ0/gMgYiEFZ73FXPNtz0DapwGD2M0pupuxf/h
d2ZKqstq+NWQcQJt9bwLVhYj5S5OQuQYTHmcyrf9+YGXTPo6vokyYCgs76MdQgLz1N2vDAdjRUBc
AvJzor/IN4Hnc8aVQzlpbe8VT9/FizZQI+dAn7f1VdO0fzTzVI5i33C97bKK32LEhFuI7kXKHaIr
3yjqKr5+CRdtEPZ+4AhZICSwNsHhj2CuXLPAVA2x9CtwTCx33eVd1In8oQK8/V2m08Yui/wtNPDB
VTpdxY+dMhHv2ky8XRQEy+newFNRoWtbeAaSK7c2i9I83AZOTJz7MAFF/+YldvDa8ayIQwT/UFaX
HcGTWeMaUzDCddnYUKFiDj16oE41H4ldCWiJqdgGz3AHiRj1D26m/YM1LaE01Vf2nrd7afNjIBg2
ffseMtIxD2mZNoWCwTZHYCNsGJsuDDVI5GXesSdQi/qQlX3VlIiA49j+rXIWvCIx/lRRw+Dgxp3G
J+Ncw8FvXuJ+jwziH3PJrhvbJnWBgIQrJhEOd/upr9YazZJoFqxE4lbIUdJxatK4qVoa7kVnrRrr
WLpHmndxu0RrpPGET7cnw8WWHOGE2K5hHkVgoqvqAv+nPbOg/j9rC8tvhPkiR/6QQ7ZLggaqgaxR
MScKmFouiJel1VuvhUcq3ZqibvPTJnQTDMmSB6y31lmExH7Jfcqw7fon3H2IxgSw5SoU1LLSBwE6
sPUgpBFGf8vJIovPZtM/R5dbNgDgqLT38KuXkyzWr0MKv6YKHtG49kSDHtWtXrEaQFbjSPQe7ohR
1TeJTo9MTJFbiIvQKhdoRZRnoJvB8QE67HRwZMOuyqNWDMqodCtWS3czhpGtWw7asaoTCzI8/4/0
LHipCNM3dGNxXQGxFmTHNz4v/z6pwixgWaMcTzRU39KgfVdDKrBuxWXpyBgrxGogHKtfV3JEuW1B
mPtYZ/ZqufcLT2r8nVO0wy8lvBNH3XAB4UMLTyZaFa18b59b/YK+CQCZ1K4DhyU1YG+c+psLRWOI
45Llkos4r48BEiJriWU0HBS9acLf+vqr+JPw2lZdH/gnMmDK+wuM+J9b+M3RH6jUTKojvUxDvi05
81i4PeF5elAPuJRa+VYWNDJp3cSigfJ3QTnIbjeeRrDa45jyataAyjm9SaI04Cx+pXa9/ww5ENtP
9KLbi5lNh4+0GXSZ9k8TBuQ87v7LY7rwp7+TPxdnbIzg+/dRe4LEsIip9U3FO8XjWCWkPDqeDlVw
KQxZxLjY5YHw4E/0Sw/h6+73Y+AlmHmlNE76JZYa5wGoToM20LVsqZapoHOYtOzmTGEz6FDWZaG+
uxnExPfK+sltlgtB7hD4aNnMY4BAb2POfnnVZBC1H220Zi9zcMMIWkgTZMwROKfwzHAvu66fw2Yt
92tGB1yuHs106tfMewd/EE2b142IeUVn0o4VEWNqGlVT21UY7QBUj8o59Pg7Y0BReip9+0sp4wVO
DqECpprbuZHinEzgSrZeGk6WvgCAYUmZ3X1CkSp4pMG0uZyeCoQxoxQ1rrHYJ2gAvvBXFwTrMNON
+dlTt7zR7tz7XONDPrz3VqircicDnY0/hFrzzD3J+t56D3yhwG9BmIitLedrFpta4aFMyYc2pxag
pdgUaNx7zE6ikyVc7MYbuuPUNRcfzEAGYqDrvlgi+5u24uuhF2i4cd9hzJmFWsHA3l8TyONcoPZg
7Z3Oy/eT2a3PQ35qAOvcrxfkrE59qhQRZADE2WxmDI0EmpHrGfIH+mUZM9xNsU4ZJpb4lgw/LaD3
yqqP1/2EDb26jIEnQLTj0r3Rtxp3ifFDxrLLVn3SPcxtFwoupWnCbodhEjzXM0VwPPoUpwkeSq8J
nkMa9/GMV8chX+lFEpZUVd1RSdRsOI1t39+sgOD7rwtSMjNd9j+T7NSO/kDEnHjFZ/lv8srB3BLl
geCoChngvju3v3BkEb1oQsvJqOIbL18EZucZU7vVnGnVbjXO6LVfPfHALh+UcQ2X5Me2oa9bCvhH
RWAfb7moUaAObLw3Ltwtb2hU0i4Ay9wY6bx0GKpC1zF85OmBbikZokPF/U/zLf1Ls3wNb3atMeoK
1Krs3wLta1duT4OslMgiLQPYpmwh/sQ4YZ+ac5ny+oqszUv8VNMwMDZNhgxR46FQ96I+BOZAz5L0
0VrL4/GUyMUi5efOMNEFpE0CYSX7MO7tJyoab3+0YYcc48ocIDTJcnAkFgaoZhltjEz409dFH+2i
6/020UfBSeOK/Y/Tj5OtBoFhfuVst8JVrFn9Qic1cqZZRb1shJBbUKWY71b9Oul7WG6iZ1Ww0yXD
QQjlQEGcnbWo74Tdz+0H8PwErdzg8zj6xqbOiB/7MnapwImIi/Ku9r+RKNAkWviue9Up+KLb9aKW
Xx8o5Iv9u55i4EtJAkxl/1qDjgX4SOE2m+/N5wUcs/T6v6R1pUZAzosPg+j+zzLrwK+YvU/QCYp7
MlUBQd1jfiPFEGdVIzFT7JremzcB5WObAdra5AIDx6m6fjjPvVajBgNb5f2EZXxWNoo9VC5iK508
zNw1C5cc/ml2G9XPNCPbqxS8E5cllDGKlq+XTXj0drIK17Dji3AnKp3HRz4myjms79A9lCGvW1KK
UDx+sPDPFuCa/Egj42P+ImX9jIPdtBLUZvwz5xslrYVVPAKM9+d+2Pc5Wdift7zYw36diu1DuZ18
wtZMV01Sozr0a8hl5tV8/m+bv8B9FcBYc03Qjn5ENfyiBL8dpa5p9mfpdefBJ5ssSjVyQmS2PJ/Z
DAWU6KWa16Cxnq7/Eeur0zKCwaHkewXU8W0FvI4l7DcYeATTgpxuObVYCYtIYyam+6tOYUQ7Mydg
x7U231JlP0krVfAcZoQJtRhTbdNEVm9Kbkh0ThuuYCF1X2sVFa4AP461qsAu6epnSNp1GROyF/CG
lAgpSFgqvvrBOdTTIqpSMGJSxl/l6CPgK1Znfwk7BhNUxOslQAxvnTnJwDXitTlaQ98B+zvIClEa
/Vea6HIbaXoAZrPQIWfkOB1hbWfODJNV4PxQ14kqb6C4qNmKF3JRGN9qTJmwyM2FVLHCXhoAf+Ky
FMeC2n21ABhvoac6gxerRl3UkaKecikhDQnoPO9dDrp4Q93w3C9o+uGG92xfUqYODLWKoDTzgVxu
L4SZmEdiIyCPVbDzYagP+0VPL4jvQb+0GFGup1gkyw17aEUihK6a5SBGCtwEBghGZY43kTKqS8iN
mDtxMFHfE3whVHxorj+kVCDbcK9nBbfcqHbK21Peft76WsNV9To2dIWkpoAtzlPBoEozPrlz93wM
RI2zxLIKT3IHkK3tm5rew8LoZhR2VJDf8cAXb++YKHkxTnKoGAF6cOUbWMav/p0UaIcW5+wR2O/f
viquBcN9HYBUYoJj9/JRA5FvD6ADWsca5oULAS+zA69ZL97V1jfYZ7Li37zO1OU4BZjDA7vl8y8v
8MLqpveJioPfi8UwnZQWBjt+MMarewCmne2g1sQQozUQHRmraWx02jl79n6lq/zCAociYblGlCP7
V6j2dFX31eDXqFDDK8TzMTeY5VT0hCBUDdnVAjQDeKxxAYBpuEP7Oz2VGscf5xrIbxG2bH0aLm5z
9yHmFeEF3XGoFBcO+q9zBkvACiI8tLsiZomF0o4D4qalxtLRrR7wPLVlVg3Ke5A5b1+Yp9QlaaO5
el2E6xI34nH7oMcyGY43ZSwGt5O25dExsI9inFzsa5KeYZjDfUZpCp5pie6Cai5OirOy57W6GZaA
xmA7ESTpXj5rspCEQgh/02IF0Y9ZQ2qSVzkMwZcIyYaJiJl3m2bOk/T6OoEvniLs/x9OttSPaoLb
F9JugUc+8/sJU3ReIAqa4XBlDsGWtNQwA0REpvKKl0M/JGnQZHu4mmhJ2fJgFf1AVhrOrOXR9ur1
DjEU/mqbqNxxeJ8M/apUXUlfoMyp8IvePMyzlTidcoR9qxX6XQieOeh/X/alFoGpJQ9AGvUgbkYB
FmWuCINPj2KPcAazl1j7bvq6rWM72n+qf8L1kJcj5SojXo1wPlvaLosuusBGufAN4BuJ4qKtdIe+
5ewCCSGyVFNTKHxpTkDJU8X9VYODovMAGlYqCDQIkkKz1QfXUVMLIGSu/DIweDIA5kFnbmQ8VJWH
qnR3GV6QcUipxDyrILmyKP7OYSG7dJudbjNUaRsvwxwvvrAd0MSo4rXWfSXeZSTPxVWd8gfhxNMX
yGrqWxN1JZeLCB0f19h3R70Qhczeo6KAzH9uwh+h8qo+Ryk4w86a19uTMH86SvKHOY6BH7Lhz+lG
SsAY0la0icj0PfDHZmh2sr6F6Up6H/OQZNtCm7k9QfSaMHLgVmNTLtULp8CTtwdYcx7MCF1ZREaG
iGHVDYU1ikNi0FS81iaDGwyAP/l7eBwqbhN5pMj7GoYMJwJnIuwvFZrxJZ5mAQWz9j/YVnjHwVQs
iGAIzfllAnuBXGn9X3J5nF4OkW3IMRrA6vFla2vdue6Mr5r0TAD91sRR9Xd3slhuwe6nEdB5KpoC
t6R83EINM5fSr+SnFv1guXLrZX3d4orJ3M4UscMFatxwEdlgh0uRKcNYcIPnZiqMpOSmG3JAVdsd
c+23A8MdRwpS9Wd27ZqiituV6fHo/TQCBl0xESh6ROkERM51AKVPqv9uyuii5fpzxKP0Yv5fKI1a
ua1zgwG2QPGiAf4PY309qTTjgjgjQirRFM5tDNx6XvLougMRhipsJ+qgtL/faB05lJ9okiUL2/+I
csQKPveywV8PXQT+SlK3UPO2LxY7OVYbG2Ql9ruS29R/ipF132VdPK5rNfHkjhPemdCgCi7QZ4Qa
iTxM0wN/D8+AXww6x24ynS98loLKw0jY3goKZFbEOctVXpoxu6T2hDQnUP07YVMdn7eyFWLIvvfp
dBKT7ZVpbmc38BQShS5pY0JYZvzRwaOuvxj21Ta7xvC4zPZ7NsLNspfhE49ahuYc2df18X9SUl9b
ai/HtXSUxGcQXE3XyKUvevqHljt4KryAhoCac3zQjui+ooQSPJzGdxGNvVSCYppS2bpzDNEChXGU
ZgHmZSgXz6sMs2+gEkuqAXqumffSGmY6P+SMvK2lHWdw7Hdg1cnp4brBLZhF5YvZXiJpzcnA3pm7
/Ka8MZdClLfrQ8nqDHl80YvJ7In8uAxb0AV8+KGstGwcuIeBrll2aUObJtNAcdCP5406bY/xmcle
M9okFGQqwe5dRqJZN3nSm6WLttPm0ARdEn2U9AT9IR4Vw40cFm4a3r2v0n/2zok8aswsBZuAMjjI
bYfCDNDq1ZCF+lonGcudfPGkw/OCgogxszVweihc21DDNwVfvWJOS250kEPN0xGV5/lqO68w1W7r
uGMl2Oa14e/UaUbmzJRA4fKVGwG2y5lr5lof+osW9tpua08OvquO0lHGTydifeYQzHS0pS++Ck4y
1B6RjM0fvPU/EieTJGZKqnhqgFqy/t1XZ6AO7KY42Ib8lrN78hbqecQfYxIrwcr/4k1+CIU8SDCa
BbECpZfPbEf44UyGRvRsBC63PwG1L01bJ+84m82M5JvXPW9Cpu/qxhLmN3GEudAYZi+pQ3YfMhn7
1oIXHu/TrR1rLd3uCQ5uxxjP4FcZV6YNSduQwubXd7V9IX6fKy2s4GeyAv0amTJL1qftvnxf6Q8C
dk0QKDlNwr7RjnU4CeKPL7xLwZH52ElDkSKNFIfdzjxyfvynt6xfP0As2CLb5YpBGzh2Kg5uSkYt
C/AQToLwsOb8mV5TX1zko+xsyk40RlA65MViMX3DYwbhuV5AiLk0+kldtA4dhyLdiplhqwmO3Ikg
GfjnqUNUOJYzjhnlzN6si48CH7Q3VoQJCWl4fndW7HbFFi3cf4W8I9mAURfZmUN9QBvGpDLhSgRf
Nxh1+bioR8T1bxA3T78MHWIWZ4iuwjcMFTJljzzwCgxR3w1rcBxMFUqHtoKkzSQ0mkCoxJxtoHDa
ELvFNtq7Wn173sTpv0dG3aPl1mpyGP5QghCQSn8OsCDQXnJw7hz/JxdQ9bNMLoD5duS4OiGfnSz9
g8fG8JsoqrbxHrJRFYhAI10fK1waflQtFgLFfKVN0o96+UMwVsf/MLQNoXA0JiCv2dxvDJHtldPU
rosdY0oryTH+9hdiUGx+S81ETx7gLYhzCzOaKei5t4sWXELIvVLIWLOXTJ7ft6K32iheRkNGZm/l
L7SkUnOnSA3S+2MCdtMSy+QCNhDwX0z86kEChuQvfLnJMhbXBmd8IMn3+FvHCxpc4byYEDdU/NEw
LYXK7eoei0k/acrWsh4Vv0jzFEuVw4HlDwFwHNxdE3m+U2g79B4D7iXeWoRXzBdRemoYBsWzMJqk
zorWE9ewE1IcOf3kOR1oN9LIxet5GyKnVrD3pd5QIBnXhJeSrNcqJAIXRIH6Q43I7GnEGP4M7RVb
lagIzqul3yDzLMlNVX0C4hi94BzGh2MB8+wrC+n/n/h0zYqgNRilIJUthhw2+eZrPBX46aD1Kwv0
Gbuh9xn1nyMMB6BZ3cQYv+Qx/UT7laQep0s9lw0Y8g+7s7r3oYYJjAasceXWpZ7hTg+mJVyC/ksR
evbD9OD8tqC6vqoS2/mVU2SKxysFxhZijY6h9S9T7cXtVRVMz6676WEb7cmD/5ibmWSwsI0tvw9O
NmrF8gISdstS+7bpaf7Ff+NSFqWVTuaAlOLgJhHKO669ZEbBuCj/UNxpGJMGpWXnS/Imtf6XMxm/
yVyvUI0JZQ4N+0eYVzPvw2gRDOXDYh/TGMsnVUFPAJqUPOeDSTlRUuNQf6uEtwcpbt/yEMrZtVPY
ysMHeTss9zvuExStysigQrkqZCsYk/VAgAyM0Lv2ZykE//bR7bf5/RmT8UaOB+d/mOO/nSN9U5vk
kJctEGmJ6PQEsuUuncCPiYSW9Yva49UduCeczX1W9II6g63XccRjTYWyLir2tM4IqFSYsO8ooWIA
6ZhsQo6HixBR2aM29y58xY2YahJx5/az1KbxF/re/jSm7ha2DzjMPC8/aIM2Pi/8DqaZi4fujnZx
5//HwtYyic9B0qXEOhndHqp9ExnGaYSRNKvfZcv0o+z/3nPw5fZMjVVHIqkNA9M+/d1IbQVuK5i+
crwvG+r8BrU07buqIZVNposib8O/fvRwRmEmhWKkb3QFTv1LyMOfEzkwttZF/P3b7FHO2eKak935
3CKZ8reX9z9cDTH7ZyQFJ1ai6LG4jLQ06oUVB3QIaecJErdbKHl0SgWsTadHuDZrXcEhkfziPNBj
kDsmzzrPabvcswqORMjEIPsaYEsp321OZIU8A94tjRvrd+WF2vHvxUdKVLWDg22G7Pg0qshYyMpI
BT8WkojbsI3C+VArZeUGdCIij68u5vvvgaaNCNUPovpyfmdjQN7R5+aH6VA8lNTqojHJqvTebJeP
e7vd0tbmLpui82wgVhR5RwdY08iDpYVIxU3gdBkWpGQJKnAEwqg1sI+wtUEfWWfBsFPKxTUiyxSo
qEoagDVCva2/Wk4aeivVNyZ9C166XkglLz+/iI3+vBhmDN7zL0/kw+y7WMLr1YjLBQpitRn8Erx/
xiDUid0DkvA0Qi+Hip3SWKj5kuLtvn5fjkGrFv2l/hdGQOgniP5/bRrVHgcSLyaEyMFvLei3BMyC
LZVy5f2ZLNGdlbBpiAVZEtkzWeSTBA4Tf8mxTGRt/c1G11lWYV8j7G4qm41NJPNJDpmi1coafU2F
XecTmaKQdnJRhvIhxkYv7Gh/FYN31IE/JpmlQOC2Bc0oo7wfi2Zn6vjj7ty7W9anUre8p41zed4N
bGlWtu0Rua3Z6mAPTgRAlcBmTi3PVVdgdBWIkjAww27OYZXIPf343KPlL9g+WI0H2LsGnV8y71qD
7E0o//Ze60BnLtnG4XUVjRjVVsr1Ake9Aw8deLDp4gtTCWD3ZsO2RAGfGUBsHyocBLOEm8Q+Ynx5
xSEUub4YLbwE1BLUln0mXLgSqpX0eH/227MWfXco49YjOZLqQc6I2O/8mU93qaO/Y4JnxF+41QGx
y5/SF+wucVjGrpAml9utn4pQz0o1urTzTRvS9z9QLbXl9JWPhHx7a7QLxs9jgGPDA+G0zmqk97Cf
0nxxyyyxk912g7j6VY8sler/SwpDw2yc2+Y/G+Q0Um8Bp85/8z3hBa0kwWJUBPAYjxTcMZzjl2dG
sMOrGHiepF/Ir/2RDSImsR97BBzvJuZNDu13QkpgKYmkSjQ4hvjMV48ZE9KpkEEW71Htr2AeZ3RD
w7Nnf+7jiDbzFjmJdwKMLraSusXGx82J2/kFi54IV8N1jVf4q1o2IYJFfYifIbPS9fQjaKxlWBAq
jCm8EKEMFSmKpcQdYfnFW2tjwKx6s2sc4TFF0pjkHWSWNNvcdqkBpwUIjzLUldlY92g8KkMLGu5y
Z+xk/giC9ldbU11nGKdDg9NSbutTDoX7F5nw7lID2VYJ8MChpGJWve7C3+q0Q7gw7ByxPLwDBwfR
Sjnc0FCdD9lDQ/shZKM2Jz0IQ+4eBdC+v+xY/HOehVGYxwcurejdCz3Jno6JsKx0dXd5+WOhUUwL
20MJ1V+f58AX/Pu2aixP9A3fDVtYs54Iz7g4On88xM03OWAfFoYTSwfm/IZBXs59Ps9RHXGhEVEj
Egdm44LvpW9ECCg5UT+1jsA8MNrawK5WdyJ3eDY9olOyGz0BZS97H/VCmDueJLGrag4TP0DSvJ6T
3lUYkwpY4OW0A+knehe8kA1s+gyKsWj/XWqj6Y7YRxvh2+9LrVLbmjMTAMbHF4sf5R7ElFIatSN1
7TM/j/3JD9rHed7ozGQu7hH/JV3xFXVtc6huNOx5hpoHIdtFcctmGZoBodavSSNNTcsH8m3OUZCC
UDk6LtEW7KkmQVCQooQoeSNpDsCMm6KB2FCd+uocbFUG3EfEarpceXqpVPlIqgSyrjvmwt26D0/O
oNL7qh4NdEUGBPT4w76QQovX2+COj2eZll9EWFJgygTh0+uGetGW+hSs1lewEZMZD8RBOCiy26+F
UUo/ZYYiVY316S/coPHCDgLeZ9CzH8y7/cHDtYUDjYb0sk+XnTAnHIU1nxPh8XJ6epwqQv1GFn1r
liX5BqRM2xM5X2XXtc3XitPsas+HfOisRGtdC/e9nmopqVEDwWzl0uZ4oeWOXEs4ycA6Hh2BGEht
L8vYPmMY25rdml3pyIr/pUj/CFhsBBbtcNU4cqd02zpXekGQubPZoYL5nCCPfaAv1doJfEClhEyD
WjjPoQUsF55lqbBY/8+xyIlaFGcBZSfifeusMj8bM4RX7Q4untPmq1Ktc6nK8MnStMLHpkVY/XDS
QlMTVErn/1x9n48ZFmF+6P2vaAzxB96MoAufFiQG54RPro63Nvd7LJY/Hsw2O2yyyz2SyOQX8Uic
4mew+lQd6YZM6a0OMGAX+NqJBZDLDu/IDAGBKJ3zHkB99MqQfe/QWPFZaOFEhkRKxCRTh3rz9p9K
Qr9rS8+uGa2hz/nUuVCIAEepRVW8VBCO8rvOQbPjpY9wx/xi3capMynPjemAlxmI0WVZpwKZ/bD+
iiiuLl/++KiQx5uZ5bJ4nstXAW9mdeJqqZqCXCw5FrAaymxahahRsQi78pFjOVny1ujQ6KnqRIOS
czZSuMkMiubG9QHthD1/CGYXdxcrAL21UJjUhfkMmAangAApD+97trhWFqswMVFgEV20CrRkZZJ6
ZrVsm0anPfMyL4Hq2kUJ8oNJ7i924b7h7RtSVMRrWMTI8oNO+u6mBETBIkC6uO3SlWXiCygzsTB2
hOuyDxuej87nzBrjw1UdYO4O/ujAlx3q8E5cUoOocEk+NXZcM8knM0eRkpEX1Zts3o5Htgyawyci
kGV5oDGur6AlOckZvUWiwGh5iye4Ylcx81IeKfBCgiLuL79rq1ZgT4l8seRF03Ab4cPKMK2EuTSU
c2JROwNNwL81vJZ/qKHY7KxcEbNCY4AEQAnC0VzpfUYHHuav3rK5h3Me/AIeblJcGaybwMf89Jke
HUV+O89rAkZp0rOhipRSv3KnKCL8l72uVDo7azm0MWCBqwTmHHJ0ndEqTuHqcexCcJ9pkmfp4sqy
drabLL7ZrtvqNQL3mopeFamHZp22P7d1qbIByu2039WADsNRLp4rKKzJtwsKl5QwZCdJL4e1kmkn
bd5px6N+qbh+SwFPAalFZS84dv/2YIK1oNM4m+3fPpKi89OJJ3OCdMtQacxC5MNR95IEly8xzlV6
cn5zBRYhOTvqtDfqXDpiOxHPmReRvVecwO61o+DvgJQDoo1GKT/HOOKFZmBwHhDvMYaPzE0GGqmf
u4jS1b6AbXmgfr7HJrBQve9zxmfXjMhtmqaYr60Bk66NNiIlU7Srs5RqA5x2cy5e55s41g0vuMk1
ntY246LZoKIj5ZyQQjiXFl7+7UozHml6SdF9RDSLRGjAQaNi/CbtNEM9Q/E43G7HeYfX3dZJeJRl
Bsr1G3upSqRihLrN4OonBL7VlC6RbWEDtbXAX9UbmitwNBiGBdmv6VwKSakzePg8Z7mAiRKsU8F7
bHc29788QvZXNAug4eOob3Xa98E/9d9Kftx2Mt4tfNG5vZ1yp0I/9STv9292pSc2yzXK1dGgqlI5
ULe+46N0WJn95DwAzA6dJIfe2aEfjYPqkGYNByLd5+O/9DeCnl3TN389Q3wOFRX+uChSEOPx34uh
7xBlMg67Ld6k47+IJ264dnphMIoT/CRIpiYiyotxqAWadcD5Lf7EB+/Bf7coI8AeAIuPAJAEsx2S
rVNtZEf2TAjYzDvGxy8USAN9unx4GEhk95EMvbppLwORfj0nCYulu9JzAR/ZNC7WAj89jZqT/tk0
H6cM1TUwJtiiEAKblXRMXflguzlA1BJymIyDMa1+AXK929JHD0Vcft+V2EtktTmfcD/Kvj1gH+Cf
7IkRha/J+977VG9aJu4LOtG5zYz+Ka8GrpvebyJLX6moA8pLFvX3IMvWVNwNlxwVdtWOwU25NM9d
tsIhfHJm7lAb/NqgDzuTszcKEotvWpfNry8j7OdTBHce36guntNOSscaFQFWo53NsyJCU9wZwyr0
J8pCSLvlCVvpj8i2tQ55DU2e9iAcW13AwJc5gwSDIznB4HSoWDZHPopsyigVHTzLc22mDsED9bCJ
R0B4rjYTJr1qfaYRi8Uyz2HqIaifls2tFEZbMkeR8NBcGZawcotkI8ePIABTPmUAEif/2zWZqbgB
axjCu/jtUAki02JDhoBWDrrWDl/jl/O52ivPJol6EWYRdRvSXlUg09xPV/Hu9N8eDAiKD/yMrmoP
1Bb0jzI7W7C3B4GJ4NkIoCq6161VrCaiOFd4cwFLvTNl7ychb0EbQoTysQqn/YXF5TyB1JzCyYzm
fEK/cHYi/r5+Mmik4040NDCCJIpyV+cBdl0IygPuf+jMMAgJNMI5PSUv7K1J1FT7N+/bo0I1Jnue
94V4G8Zxs83PFMJFNLv+VFHfQ84nJOWsawFGAwLBpZ4vRT6c/HBWdbw9x/CD4RRlXhAmuRH1BH+b
y7MCcTZeeiWueMPy1r1nf3jZ6V38rg+32CkVumTwhhkOiOb755YhUJIPqY7mzCyR4j6I6hui0/nb
qlCjS9u6veUoGPbiEW8gXzReLhQaCRmTCWXHvlM/xpA+R8TrlqNiSwKHJanaO8SFtt9rWLjd0mYe
cRkdI38Ml1/G/qe7ce8v5AvUCsYCdlYEaGaBe1x5rgMPRyadJ3ldMlNpcVPhsk7U4VC3MbuF1Znc
m6lcHolIdoquhJELJJkiSglowKeJpcPP1HE+K04NNuLIdP4eRVXt3pyBu2lCa+elZPzJkwCD+9wt
yylcx+X3gdF1zMJHlpcV+G8ArLCew0XlSyI3ix1W2kaVk6yUt90FNtbP8i8W0d/v67fgZ74P2w0l
N8I6WTNBCcz1EkEIWUI9Lv2npBvqDN+odKvgT2laB6udvhwzljHYX3BrKtXvpmoBvXlTkZydZ9lf
IKu04XPhMrEqRYZ9ndJq35FZj5ygb475RxGx8am8UCiw5eNPShJgxzuv+BRlmQ7OtrSs67iL1QGQ
q4m5dz78bw1vAvHfx/8sGzi9oAJ8Q7EINZeLB3cPrRyBHcqoLEL3kg4frN/fHaPtULs2oKRvB1xk
44T9v2f9yQquXdywB+RS1LnyijFkpr24pMyefNdi1kgqEyvPGLER+E12Xvgo0WaEOMMX3U9w2wpX
JC0ZegEOO0k2XTnMkPLLLYw8OIeVX2/RCV2/Uk+yYnHXdXSCXRwlLhz6nruyPiBdFa8JQQ8h7vMd
heYkUMsAA99usVy164p2ONCQ796WBGjuLnnPtsAGokNNBYRTqwr/1Z5M4/0ZHQATa4C98l2bIPVD
M8gGobZGPAz34I74J9Ibs6ts26x0eXUgMgXyUIvXQdu2nOx9hdP6ramwUs/0R1te24C3zU9AfcWN
yhXRhKGTyUsMOqjJGHsUNg3pRpTztOShUp8IMvDuSBi/qwArQZrL+UzzvPPn+7TyE5eGNlZTy9BF
l3bZc0JMIntWYPOT86AIZr5d6l8wPdkfdQ5gtGp7WGuf+ySxlsy/I/jKKip26BBiJuZaro0qmLin
/RDbQ0HueTHiM0L1tdyoyQV3GZukS1MrPqPgWpxChbNE94UJ6Twox55WynPmi3y3ru5PDgixqszC
N2sGS0Fm9FPlI5ER2F3Rrz3UZtSHy6YWnLGsnD8BK5NqZultbjKqlBCQ8dx809dRXId3gxJkxk6m
2IJRKW0Vbdvi4E/40i1BsRjLfrTELXuVeIiAde8ZTg2TVGQU9LNJ+x+2YwN5cQXOwR7u8K8YbWR4
q8nmFqw4Xmov7zrdYF9VleYVh9Exs45D2+wEQKqop2GNcdJHUbPSa2qov9c0EoEFM9k2OQIqLGFV
WZNkWFnNamlMciE/144xrz1FCbQ+jGqNr4uSClJ6mwL4d9ID7eFEmHzMyVpi9vzBDCWAeuBmb8Gu
xQxYF4kfvPqV0IKDb11hcKA3e5MKdervgnlJNkaSz0KDWJWZHhgYzfKIbQ6x0B3TUpRCNmC1RDzR
oEm301NN5tltgtbQTIRicSB0Q7BN1uXWHQgNQOgtg0LXEd4XrDzdo2vEbZgxB2M3v66+tHGBRITA
ClouVHet7/rQ5ptZ1fR22y7Rua/F8P8VkkZsKYN6jBsTlPO5uadIYm5NjlDu0ew6fl+CbAq2Qghb
MWPGNZBlXbpkfg9Y9kFofblRK56X0ooPtt9hV3BeiTFtUIO3SGAYzdnXAxme1EMYviVgNIAavBYR
2SRi6Fu/PlN/xadUALY8zI30b6iCb87mwDDhr4z5yIrG5Lm+cgnCY8r2malZQagYqTp2TJzNuv49
zpiOEiMzgCWAHnq1TwCqiViLf1xcoIfAUZRv8hQ5mbt5ERXdCUk/l0+VZPh1d4tAjlyrG9RBb73Y
R/VEGVCJ5uuGjC4Ld0okKGUO7XNa/4pZxONr77jJut5+/CqQmOkSDTgMcnB1xKowkpzpBfWeg3OK
6z/QG3Pa4bUZb1peQvr32yUaTT6qDi8jxU+JWqdcl0B4aarwaKJrvZSjMRBZkaGJtEC1Ky8gSZh2
5Fq5GMAH+Rgr3h7ssJ6h9lq2rs5zAmzlLt/3tl8V6hs+rce1/eSINX7vJ43lLwoabxSXHayJ1bAC
0N9tn3l4v5FX+SJQQL1jpX6+dtioOPeX/duwkH7dlVwAEqH3Gc/T7QTGFx+B5TV+86JITlVdnfO5
I8+W+1TnGthM59dhUgRiX8C3PV9/YgbKIa/Dk2jViqTsET9ZRhArTCYArkCe4t5Faa4Jb3DZRfjE
qE05SktJryNfSvUqzR3a20iQES36MoXxr2LXAYFowZAHW1qKhA4CpsesY+9lDGynzKuWLgekuObp
Kh1bcQiTJWuPamvouVvuXPhNoseXnmL/fXrEDuy7weL1oraSc+0F/hwrB9nSNrEtix+GHh4Vo3Jj
DEuNOkUAQB2/YLzGeFD5zoLOawpi2prdhpr/XU1uRWSpfcc2Wdyq491BwMdmxGLqMuzF9aC3XUC/
mY1XX32KDnReVLvnvWnHH+glZ7+AnaNRuaPSha5KjLAZYbSTqz8uhj7IrF/cbul+q960EeGM0gFK
TouD+AlgbjoddMJ32CGiibE08QDFFPvQMIy9H8bsRbXXPUqSBMe4FawfvI+0luwddGdSH03GLDM1
53M7Hih/fPElzghYw5NlSKTmTeP98h6mZfGnEfCE5Mos+GblMakdTBvNbY+dBZ51wPtz6EPMcowu
x/poJI9j4NJlNVjAbPfwJuMjm3sLIZGtYR8RlOmoMWWiLR2+leyfjEfNI7eltX/7KDr9SNQFQHTE
MU3Tuelb9Y55lP6RdqXo3e+79x4irBZLV+IAZhlb8Gced7mY5GxwZvw7PWXwe1K5tUXRjHfUA8p5
LD+nU9OK3YQAjBZDcWfn1ZiucoC6mnELFcz1x/zdFXcfyWAZ5K1vq14z44it3/hvNwxmTd0MOkom
QZEBkJEDDqErFCvtKtSN6jAul2WCy1QJprM51MryuEo0lXNH0NYTw79s7Fczf0zwFVdGCN/0zPQV
lmTPj44vAWdSFUJWOed7MJLhtWAI7dIgMBg0LZiprBClpAAJxJqN9ycG+glpgNA4KJ0Y8geE5DMa
jJTdi2wS0nGOExvi9TWuJ2SkgpPXBfls2ynGX42uT/rYsVkLMj5Ru0iZa+osgmuEZvidGrpyET4E
4PZodLafj0c+mP1QbshhOUCzct/PFxVU8XwIP6WsOLgDZO5u9HkASsbgIkK99n9ZseybeiIczndx
GtetJpXTFj2zlNWYcyWzZJ0q7Be0L5OcmcxVvYYi2fr/4qHNUQtXANKCO7RvuLw6hb4HY8zIT84y
u68dpBjUJoSvkTATTi+tnKd72dKHnhjWrvs77Qs82w7gQ5nqwZbiTlNWJD4Enjr7vYDqXpP5LyGc
LdZczfJkBrt5aSJ1ucSO8VcDnpEvP6p0pNhbkujZA0dcWiSsuFbZFlmeBusEcqjbd+pdmQljAFf8
I73KhxdjZmd2TE79AM0mNqAQGzavAQEohA5xSl8RbhuNyFDqROkMniG+i7LsjmiBkpm1iDTtq6E7
Ll8Imy5kabUv2FMLS4mKdn/n84rF4Gv4sLNuy3JQ7T/Xf3852sStmGh0Xh2j3CqY/dQF7Lawu/Wm
VS58K4skoXXrEq1bxvzjKD8prkK+96bamjfmAbkWaCz3RCFzpnPczgkDpdHtchU0xFQGcDAp1OPU
HHNklla3zZALt1HX32tCOgqOAb7l+13NSEC1qbQ6gYkuLsTThUxPrjc8hEYM+/Qk1sxvjthIEXns
froRnkyNbPH06FIBB3wnR9VkmJpzaPU7q/O2MRL9Hv+4P2ksFO7i/YXpVk/vpOwPhW/C2DCGO47B
3izYE1QvWQrrmrS0vpKA8Z5vdVtbPPygzvMnjzGKDSbxmeNfoHYiyX0e46qEhJOjKWkZCpE2YjBg
kLvd8uakqkeDUcARmbGE+xhcEOi+p9nx0Gsqub+UYrFnnL8RXN2xNDppbq2xnm//iVvIqvZ9yFtw
FBOxt+5Lzkn58PB2tz34oMtGJA/CtTTG8Ly1oAHiFx+O1WX6ZuBCuVOi6SfJx89p+DiE1Us7gv2t
ITr0AIdu4d2HBRwSmCyJ2Ms+PEmI1NHguXvsX/vfZL/4P/etownRSgSG4zrwJljy46LYjieW/ku0
+C1+XEgQn3GvcGRUQVAgno+ryhnvjCA+ACMXv5MkUoCgWMhmLo4iVH5Wv9noYlcs4LoRI+5VXkwn
LsIfR5FVE51a1Ojw6ctI8VfW2q0dunsw0qtwMek+7+IPyUaE93aixZlkBZ7T8hcGupsNxjcY8+g+
X9adik5NySbXPSccPTznvYBSidoIOkFlA0tUC7BNYi1RmRTulwDnJROqHaZAvCqT10YW0oq1wogp
iyFSnQZTBIpZZWyBDQ3jvswUwKtGTzl+RUB9+WIZAa1I8ESuybH18PzHrcAHOkf8dD/+xirs7cKU
xpeeNlbMNVBzFCAlZCGdJJoD8Ea0ShoTIx3/46er/Ub2NwN1Kl/BaaAqShnCesXxg/YdMiIjQhg8
miCJAwQ9UgMUU+QML2TEsfZhrBLbB9FCbc6bbjnl+6Rb6D6PeJp4lYSuQzhdqiLJ2WyoD5nuDBXY
v4lsFM0PNuTFp8Zvouo91Tnub96pIos7ZS3/WCFxrdAyY6KcU9JxXE4kCxiVztOhnPJyhHHI7AKh
lillRAXoDJVrhtrwcSp6JJPowoe8zPeT2j3HPSxfSljMfFvZFSqfNdVbi+AgBSdBOqpGMcfWd8bj
yh4BXgYofxvz7cidu+x5I5xuThJLSF9T7VpABYMFYOBMpy9are+XX9Lca8VkK2yyLn/wp5i8i4yu
NJGQrDw556F7eOM6EKrrSyRjYTYTK3zESGEi8OFfW4se+yH7NAoNGW8QqEmum5jHskFWfDb1tfrN
jUTmf0BLBXi0VNENoI/gIs9szs27trXagoEICS4CATg/YzHZu2rT58O2buPFlzSp1yLHFJ9882q0
7Pmq5XtB6p1g9b57mZOokRKEi6hFrLGuhA6Jkwk1wRyNrGQ4nkFRUYGaeCIUbasbD4AC6Cn34uA1
I9PQwHuQsxOJ7kXSzU7a4lCrWaTCVsUGM2o30GylZIGvXWFJftm3nfz7jgcc4W/Jkl6N1EmVwg7I
XZhiwNoHCvQ189KBY5b4YH50Q32bX1neE765g59WFFs6vl0Q4W34KR/a/ZdPtyykaR2R3TfJUjEm
UV8G9fgT/OPrt/Gq0b4z+e4Q0jiFgYQdqyl9kH+a0qBh4ImTjsLDnP2Du580tNHt5JqH5/DkIBuu
xbFAWGPWJasaoCdTdnxwSgMzrBZisUhOZN1AsB6HiXB+fVh0hHW+OjWh9uQd23A8b+JwFeHYB4v2
lS9bmNLBBEje8DkGuVpNZZxN/y9lRCTx7PHrReYJbkVEdvJdXQq8DJ4Xg7UYjnx2qGtkCLYAmYHC
fjCm6YgmQFScMBxHq4iR2iHO2sM4Rz61oEmh33uZ5ES+FaT21/Ud6V0OepIbugjnXxt3aMyby+vE
1LZrL2P587bOtj7Zlu4UIgNr851ID/jBKxcjwQXXeZ3oepiMm5npUHBBZPZZySqGIAahw+Akhg4a
uTvlCDNuRaIWnOy1/CIWYDg6NhcgTSp/SQeDlr8rqBT/oKP2T/QbyF7TXAtldQhST299koCObj+W
3y8DVH4fl4LtdtccHBHPccVyUKYOjBO/TouB2od7iXinLuC1e6ho7tLEeUBtv3u5uwVIFXie7V4P
9GnCkvXnJxEhDV0e+pbZh4whoTsjI7PESZsbTgBDb+fRpMgJ89xrAvfkmxq4aeodcwvN92XWK4FQ
Z/eXyYwNB36InnlH/P4gobz0aRUwPGPkShkNq389BLUaPA82MKT2d7FA6G10NcB1JqlsolvEIfmd
jgucwPdgxg6lCcTq9m+o1Tsanc8wA7Ai7/3G6etQw2/thdfu+phjGlAkna0lVZpYsrhoRcpZLUnU
e8jrOpHydKYffO+NIINg4bAa5wABQWErxU7Q3+QSFjasUo+I9fUFQ66FBeGj/lSZKclLBOcG0dAQ
haH0madpXCadNGJA9V63PHRM4oR8IDUHEGuLXxdemWPuUzpg+bwoLKYQzgMV7Ju1zF/UseGii7hg
ixNaxbPYNQPhGaZBBTnqhpm3FpkjMbd9dRolqf60YC1b09IzFHqFcrs5HgHFUUkW5WQFm9jEU+c/
Krnz826JeylXLSXCBoDvv8gVwJIP4heORa6jCQeTx8KXmlFzibYVX5VuaB/0LwqSpVDH9TOiUBgi
lZtuzW9Kg/XgHBg60tCD46Im4i1MtOkvNEA303gc4/gKAX7jPKcNFggBC/Zcgjdb6R5cW12ggGCk
8vqOoXqi8824FZUQx/ODscmIQwf96k7pp9D+lNpVEG3sJGK/ozfc7sITPZ2idgzk3nhslRxZcqEY
Fu660TIZxmfI4vL4C9c2ax0YmC6CKzJDKzJIWWMaTDaGuJQBkfPG0v5Y/YB+NrXkj2FVmU4h256b
YIUZZ98SbVUs6Wv0Y2k3Us2UHZishGmpMIQqxKf8JzN24tTW4BCfFNrbb+Y7pFv4FQTp7igYx8hP
YeQ0LFTjJLEfTRX2MpffWfsLF1iBvVl1FQDL3SUmIHXo5mA+bYp16ilF/63/Ln3mvPaCuwbfv4Y1
ytVQxRKljNpHh+B+MnC09KghEMOxAOIcjvi//JPHNRHm818whgjE1nks9+yQH8XXpuH8edmfjJMt
e+nBk+yuH2puJ+ULIFMcsOMBH19mlBkWZotwm9vEhnRY2mZ/LoV/pBavAv/bUWuXP2yqXoUWrv4J
YFs6ItWhGNe8AKvZndGKVf930Env7H30KPjW3L1J++VFM8mpN/1NfksP9FDiV6HcbZkq4hJDSXLx
zoUKDfPZAqdX/W/0v07LAxO63MCvuR+kcB5GKCOEQ+V8kVDLaY9+BW/3ncdta0eUQinRWNM9y3Xo
xd4wx1TjEpNSbslt6FwIVGmuy7UCksSF++RV8yqCwMnMX9eCMFOU+j48jQiGJbWOYg3CQEyHgARo
slqW9FRwmqMhN4so3nEmPqGCpe1fTHNHWqgAzbhU4vG+Jz3ST6Z+cH6VTb0Im6lOvhdVG6/ZEqeo
pBkZ7BoILQdLJCghMexI9/sIPU3KO0BCOTgh67/338xTr28RubRq3rnx1hreSDssmlfkhb9WXG2n
vgPacRhnpz8OiAl/nXn/1V85E7MYvbIHDD22msfnnjt5fLc59syDF7HC4FEcjuZQg/Ve77wme1Rf
oYEGi/ooF6XP2XAdbGu3rU+bIkTMux9qZZ5lFqRcxJWIHa1fz41JSE8TdvTnmesj+7qIpPpEU8A0
bVmzBeEG8rJ0O6jGAQ4QFJei1YEzc1YZN56B4iJSeqMy1zVQXp9sIV96Q1ggQLI/bkaMclr69qxd
ia8uMXVuLpX/YlV2AeFujjsQdD3A1zIScAC5wcRH80HpNcok7HBDx/4+MYp0imqCVQ2N6r3QL6u0
DrcKLueXPXsDW+u+upVEtTMgYmR9YJ9fe8MxRwPqUw3H7UW5n0SSvfol1QB+RjABXk97moEvwoRC
zaGw85CjBh37uh4Wy91kM09qUh4XgBhwI28ZTrz/j5TiL5XgbSClxfsppiuyulCD4RF2C1iD6FaT
C4VyrKdDZ8tV1lw8IuEGeVJmZWWVHCy1ZzhjrjOKYKsqO5CSO4aua0rBbXgXA2/F0eQl9qIGR0R2
g+H84Ek6GJYswGI9flInN6lW9T+jg2pThccupnqHAVpdyxI05Sk1YQvZ7kmf89OsaPR/S0E0wMwd
9crj2KxiQ4BCorjxUqhLFxlc5d9l0w4Wjocba28TCY8KlyuOrVlrG7BRU9hpGBYvrpEy3a8nYKBq
UVin0pxp5icYiyMFpOd2Gi9hw0dknl0XmktEqPPD/EzDI98W/XMsejqlNRdYUhvtmXua7Zmh41Vd
epdLgUhHSP39+mZ0ed4y4TU9ksWnI7i1BFdN401adbcVa2EfvW8etNojkXMyFLeCvJS7llWZksiC
JLPHc97zkeK4xCkbmq2SpUcYZQiV+D4mcg0EhjjWEJdNRtJD1HguQdfex2qKCM2wm9+p8O3W5r2N
C+WlRRh+7B2UOZ6hm38f/WnDxBaMVnN5Ke1wwtOn7KOhrzrVp2Ox8Zz3eHetrsPIKFDmLQo3wLh1
wRf2redEYX4cTt3jqELFnaOWl7JdOE3IRnx4qu/spZ0V2maMd2jevyOD5+9VKMdoTrT7c4dzixu3
DBc0pKXjKxgLbL3bxnLczVf7HUgaSOqNmzeGJgPAMK0O5OM8wdIUYJukfHacW/j5VYBrm28J9Mjv
Eln8baSvGuwicBaSppSsZ+PiEtuKINNk4I+rizgbK6o8ehJj+ZgbzwC+rGANd3+SD8z4B/2l1dsS
OF+PirgavFkaeQv7NVcNCYWSS2mm0ndY93vZZRtWh4cISzwo5/zZ/FbNTSGW3MuaJYgFZ92PpQWB
aTawgt/zXNKj4zuUU99T/UuuT4JpdZKmqna1Gu+td+Q4JnVLSuhVhLTexoMfBjjDDHevqKoNYJBD
I8JKBX/jxANoUCUM4mJqmX115NPDsy8J/qUlTJD0YG9QVGGNiOLqbrbdQuUA9yPNYBHQZoX3Gsko
pMBDyGYzBhgZJmtg07vA/MpGPOMLfZ1jSoCBRoT+7JlvEwoIz3XIlNUDwrfi8pUF9Oykrt2muGHX
1dosjhqDMTvtWeH8YfPbnf2KYymSbHkly7NQpm5pKUBtgRhNKxx7ZYhsn7fLh3tbnleViE4GUNK8
icaTLFYt84vq3EyJCR0noQGZjkdcyojjZmnMSSWMmeA78xNuGRLiTTwZMlFQmuL9/ICkGZnvygKh
V6VGCz0HBIKPAsPxU9DQLpx2iiV3bIW0sVHpWWT16uCLGTfp+ynC1U82CPUW+iGtvzVEfwkngpIj
IkqphHG9TSj2hQis3kYNzQLT+OfGSB4arzaT54SIMuonlU/vTnBPCYT3/n98XNIJnk35NOkRdZuK
VdCMF8nuvbhkEAlajxb5sEOL8FrIqTFx3sqzTb4qGVyPmTgK4egnRXs6B3Ik1aZvYoEWgTYN+JRm
Moa0c84GjR/ypA1YZXbUzElL24qrW/1XAjiCruiMYxNGFJfgAtoj35u7/sKVh8Y0Ha6PN0TBPY0M
HinzvqJPmaAG04vQQkUiSrXQRlkFnZtXM6Q91oyEPW2alEnfsMmlwUGMGml/brZwNxSq8QvFcX/4
i3tBQ5YxSGdAs3EwBlSiwa5tMQBFULmZU1RSIbprtRA8TUg+lAGWrf57p0F4ozIqUbXiEZJDsH81
TlN2R/mCd9B4VrjE5VH62adeATM1bstGgDPlqJAc/cBugpGKgyA7wqbeRXMe0Cn1MW2dRIF277lE
3n1OBin+U4STS2e0zjYJBRgZSL4pRxVjdJZhyA5flGzZZbVwiGLa8c0y0uxhBbrHYPS+poqlUumz
ocLUski0Vxgn/EA0NtcG4T0lzogk6DApNycyTtmrcL0zzC9P8BBWFamk20y95+Me0grTeF9zzgbI
lZYS3yOoW2mis16F6HmtuL6s9VKLYgLay85OP7FjoDNLvHvVqcajG0uJhDHQCszsiKGQC+fc8FB+
hz8sYWvZoAli+ccKHMnI/MTbJ84eDh4sFyIHf1fUKMDnnMw9hKDeRy69V1/f+zgagVnbohTwmh1q
OcRxiBLSxjv7a8jQk8zb3Kt8JjXR3MrfaV1wLnyRrUIvSGj5tahTlUtMEeVGrLt9RzIvI5vnPdKz
ly0s6FmL5T6sxCJ7ZfcS4otPN2pGQ65tRc8Ud1uO0uCmAbbrC9DxsDO+JR0ixh0zeHtfL8PTP9j7
Uux3ERiU6u/2ul69o91WgNnK72zK5qHGiV10sC6sPwTAGyTGW4NvGKJDp1IPFjekPyo6djyI2p0b
TJEMgKDsetp+6RAHg8PGYdxTc6XZpoa16sl+gD8cjDjWY7iSy+jXGNDYRM13MDCSa7ZYV/Cb8Ork
eM/9MPauV70FUGNYhvFVm9a+rtlA+1N2ABvzCnAICAfn9HKi5AyTzgs8y30a/uqGoqt81+NQCpGO
a49XzEDJD4zDpgprq0hq4iZT/58NWUxa5IxQFnsmHHHcjWCHqED+FIjdXPsiJglarjJi8GxgVW7o
aX/KWWBqydNM2Zz6SkE0sPGG2XOmYwoTcHd+blDiQeSNsT4BLVymjpQLpqqwGh7Ke6iJX8PDA8py
CrimTrO3yGgQVL8WyeNG8+wa0JaaTcmjEpj5bnN+/pqvgKS5kRHZgrPD+KjDH+wrY/fEzhw4s1fV
hgWbCWe2dQ/rxaquZ83VvVZ4JxTGuidvMKBJhldxryy8dgXxjVoLWdNCjjMiSK38Y1vNEZzfbjbu
GeQLfkodRRVremnP7TZIlKO0jEjL8HaIa5MFL7R/c6ZYzT7ggO73+hNPo5IQeCcnrzjHo3aLMPJS
3t0GkwHisEsgMHqLtXPshaPHNvNRYUEVjEnnRRLGcr4kg4dFAAcLI3/dFndmv8cah+g47hvDG7qu
76jKdQ1+LFeyvihmn8YWZfDGUMolVYG38HXgTHgIwZAskY8SLHwr52xjSvFuc3s8rYJcpzuTZywf
4h1s2fC4oK4sQ1tRfpNgiuWTosx3DhdPNdO35Hy6GU0/68BSzqizDubuOC0XE2MilggDbp9DLrQb
FMLwqe+9bOJGavXR0sb/14VX3Tz2Vza0Cx6bx9XmBInbQXAzOo/5QXpuxXwA3+xFEnODqajwT8az
vjeDEhccAqH3CuwXXskvjofkB2d5qt9cq4HiP1PF0zq0PSZTKeLtufWLQ/FSY1dAMkiuHif0O9Mh
7jW/Tg3gMRZiP2+h2KJT0uCLk+PfgHBAeFWK75dvNV00D61wlAbgo+c7mYTLBT0nfwxICZ6CP4vg
fyadMbUH0ZuJ4tnGYjplR3HFKJZI5S4OnEkYpVk3lgCc3J8GYqoay1MVQr1GdeyDFpsyj/c4Ppm3
UfnQsj5Ytkupp65d7XVQIIgz7yU+nk2UTAgrlkjxmryuGa0TnuDtDpbldDIPZqVwbqQanLThGtlG
uZn+fdDCv8R2QAjiguLYw/KXIgxZqBs0Zoa/ALNLCUqn/n39WkiZJJg68DupTxmTm4HrGgadMfv6
8zG9x+YNZor6Ozlcjja5yhNZ87y9UrVRrBFT13inrFhXdbgegRNyAqAkNeySKPxpTOQ5OHdNBK/7
4kubVrCuRqxpDrgG5sQiPtHlBWC2VAW6rz+gT0LjYyrXSZ45PfF4q0lrIzdbtJLFSR4au/FHJoI4
DgftoOAG7O5d1LqYsZfC5j3lh1p6wzo7y9nFxaGerWly/67tpi1a62t5qzucc1mHNk/fQmV/AEhS
wPuBcc3yHonjXkekR+9lToN9K9QYMkTkoku0fxwMgcqgQPIX4HCeYjnFYO+PnJ4c/HsvGyBKEugJ
CPHeQyAxzZSzS70EGCXUZylZ11MjMKlrBd9ngBsBoiyCjXuLNtvQUfW0SDRtgFZroPAxKeKtmhIX
jrjpiiqLW3s9P6VQCapRrnXOxFyFaBTTp0pYTqsyNm/cAtmmhMqzbxPJvoTrwfCBk2gJSfrLKAVj
tChaL8C7M4/1Ya6d2+t9ZNP4YRUGE0x42KOK3caxJTUsNF5McXaUnj8KufZRn7CMvmRPYt1OadyN
MCJPXEIsMwa7NKd1NyidvGezvd1j4uITS8pvworyI2a4R43FDJEmmCNDlg7CbU482iRiM9vB4ZjA
ly/ej3tRQotFDbDYjYiZ8wmQMznRN8tJK46cw3wa2hmSA7CPKXn+rlHIa2s0LSAcVYtd+wO3k10Z
Riqa0N3X6JOCvOufGqG6ZDpMW1nbA7DRSBhI1qxzIXuOnig3Px8f7Sgv3KI3sXAGXa7vcrLuZeRo
Dvs+cmNWgUwbffH/KunwIC/4JAdYH8H/RNaqJUS6kuwNmw6B+w4NOmY+F6slMDuzY1hhQx5IQGP9
6xEIGoaYZRZnuDZOYyC1UPNi0vFRafrBRzFXLAQMpc6txpMg+DAjx8m2of035rWuQ3tO9gyBAv3W
kPL6YIYBhU8/M1Hx0FdlP5hMw5lZmXyiwxiQhyHeM1BwxAYpfRp1GiDI6Gn9qLW2+s4m6yJ0xqrT
anEJKykJB/IcuBUNkZD8coy9pNtE4VJi1wxfMg58PMyL8uYCaK/Gwf4Cj0vgMYjwdcAyxOnYj2M1
sdKfzzw4x3VL1/xnqU71l4E9EZx09pgEruXZ5skHPM0dZbS9M6Qh2feAB2vtPxT76pfZi7eV5C++
bQyQY+q/NZ9wfkj1PpLrpCCjHhVBkotRyxrkH5fDYTc4RTxuQDBktf9bZlkRJ5hlJTMjm8qaaF3c
vbGh44l2oK8BEomSUwa/n5kntUATyZGzj/KR9Wmq64mWxUFTrCfbWbwbYUZ2HjHIeX6HnT4Qawka
9E8Zjm789igGZEFDX4Sunc3Rrx/rRCgYvxSGsvNC9NDmxBvWzSvVLDRgKZSSfZpQlJ3RFyxuepcM
/Gl+lGfQ1fEB9B/EKWqT862jAI5egjWFrSimB5fUnEZ1h+IhaTsAVmjbCLZ7on5Nca5G2GOEFMrW
ckiUDL8VW1OKe7I2ZLGH3Np716R5FY7nfuw9c7+zwHyVvjJD0/asHXuznHEjPEeFr/JL6+iQ8IIC
Gxw1DMzY3V6EsK6qfJ1DaigemLNYxU18iOzVGkmhN7eA2nEGAJcm4ZotHEtmNbL6vnfYS6BARYrf
1f+z0D86R+FmcFlslGv8qnrhr6Otgy6ZjMPmWBgEKpncMX896KMIIBgTRo3o70+OP6oRRm0QCXny
kVIc6dOoH/PUsGLGgERzInQ8xRK+nIyWKvJFiTNUet24eOcFrC5u8fh20nQMipeeIFDo0FQdlV2y
xPDcQohELPQnr29UxxARWlRzYcxPDmXaOOJajexFek8ZetMmOl9s7yu828RpBoUTWrW6EBjahAul
iVARxAbOZXkXwd/qi5JvxVnYrQNxLxlXWxzPKNX/8PV/NK0YqDD9OXO6bLLURTkixam3DyJ9IgzV
/WeNmETIxU66Vk8csIv/oga62yEYOWdaxaWLzV7KClePV7Zi5EFYAZg+X6lcqGRwfPvGBzO30xrT
Pj8x82daFlBP9ctE4ad8Spsq+vN+TCxGcY0D021Ik2X4kSLHnRMrIGBEer+a1KptenatV5L47Vi9
X90uhFBGNIcNYw1AkQrwwSRHCDSekUD2OZa1OFQ514bvLPmgnQtXO2W+7DBIC7CoS3dDey4MZxC+
4omISLuVWbmpRvjVkcIBZi2ytB7R3fnAv9chQ3KgQbvZWUBa3mWeho5fuceI2s0g0GtvI56jfMeP
RDUaJCZ6uwcKK8utklaFamT1MIgBEp73JyZmmRTOSjQ7UyDjyNY26IC7WI52ZrsFF2aSFok2UKIC
F04g4Sk+c09vS6PBLENWQkB9H4DynlGbprZcaZfTGvkaaltIkKkvyItQ/4f3bKKzC3TE2czlrQ4r
jxt14sQTkC9ff5cSS8rEfXkumwUIYyGGtgsXO/1P/x5fVfrCCscYYUCb4xBNx/2ISaM2sCNvV5Gn
JUyZMyd8uB1CboFzlHieedylwE075rnfSTBNn8Wyly3KbSXve9Ke+/QM3omrb9xAshSDJaaD5p02
JUZ3DbIX0xYDqWnqF42mMI5M5syB5MA37AGA7ZKxub9bEpsOghbINVCwf6b5ty4oZMnbtq+uVPc3
AufCO4LWEGRS3Nsf8mQ+tGszjWnU+X+1TB279U372ScTy8XB/fiv0CJsmk7jwp1v58tfUpLJ5GuS
opTFwZqNh0vcEqgH9Gvg6X2TQGpCc12w802d/Piy/ighbXSuivvOjgYDFuIunGnowbSplKlU965c
cLBrAzCsZiVAlsCE2xvw2DrG/7e5Ai7XxjbINWCqlVgDJgZdC4y4vrS2dDCXd0kTIh8C5LSKtHCN
jj7G+yxYgCR8d3vhrIxmDcHuQJTXoWJSP7O9pnuexhQZgMNox4qjv/77rdXDIRLdVG/s8tuaaaAi
m4RJiYoDmjZwbihlxR2Nw689hIN7bMMqZ3+zfJo04JR1i2BlUYG/s6jvqM56K4vQ3HZw2vhNWAOU
SJcriBYvxtghHvcwaRSlC0IEMRXvp6TARswwoVAyjfsjz1ftQDCb3XmWKHBUPOHL2RKboKMoemnG
YLoNuyDKLAbJpU5YVrDU8aMJ6DpFh2u4ESlIW30O2nVR74yveXJWdUTWokBkAkwMxOxgeXLA+7ci
MLmjSJxxf4xfSErK5i2jGnFK3vWVK3RMOdsl0JAnVgxmbIqxtSAKigVGtoMZARv37pu7NAhwu5Dg
N41eT6oTjwUQTNX+sKBys9BrKmWA0DPuKibUSgb7c5SvOf1oMBPEmIFa9/RdtV9TPv+OntFf2x8t
Og/InKHdzYEiSWGhoGgd0FXevpjdFjy0uQFSq7tcwJwMbsWGTF983vRkV772FNfM1DT24p1Az2tt
6bVPk1Y8MXAWCRcs1RcP1KCpr5JkV+7DNuLTsaq4sfxb8StNnJmRvlDBhGxmGGvWHBexWpHEAkMM
idWwbwSAWvtnsrq0K41UvnUndc04eBnU9RPZhF4eRtmYdD8m5xRswtm0LHFXBF3dGptjHkfGJPVg
toZHr8z1BNr9jXDMKMUFbIjTl7yjZpXxP99+zZaImOZa2aNyoc6XGwnXn//Ny/RO6uDl+YdSX3rY
ILh9QO+3wkcbm9H502Z9vUXXLX3gETXwaUm0UKMxdQU58VyslR46Gb0wKSCOd84V0annQqVkPS/c
jlTM7lKdeLy5Jq0GrNAYOAqLmWNL2v7cAaC2KkdlSeAIdLB0JVHCmHo1oMV0myRR4gvaAe2uSOZ8
UbDQJnd7jlcb6C3ZuiVeyJKnTgwo8Xt6bbG6HBJgG0awHfXpwxRjnEJ8DlbUPb3pVqIL3KSTGPG8
n3Hg4pKqTp0qgOg9BjX8U0/vOz+3qzZ45TwLrQclDj7tcOXfzzTu+Mt/h5UoaAMlM1KsITpITh6i
AEbPMa3v8M7a9JrBA1VmhS8CQU6UwGPb04n5+LRW4W6bmWZ2hVuqAyozkSbKtLCmCIgQjvEKZmMO
CjryVaiiRrC4yxatKypYLPsvfir0j3xCA53o43bMUGvabuPrekdJFltq92rxNRkyC74Xjzpgt/X2
OvKN0SxT5fPqxDRU6cNeCqN38mP+QzvbfMJXO/x4g268eXwcu+JsOCZwDsAiZx4Jwllo9x8zt5us
VKAa+cayOwD2EcklxoCvWc0HLjK61e1+zQBm6sWKo/YMUSSTR7M0eeWfAcyKPgh3oe0gd81YCMsz
mdL2rydT+qcnPF0uKlOBfJdm83hFKBcviEvMK3/ALl6fkDoXJV+IvQHjciWJscozb+c60w3PXb2g
a8LDiQbXCdtIoLj++NJfL+SnwcHrCUxGQgrz5pGkYKrSaS/+jqzcWA4x33CVQU/xgaROPNgaHnbv
EON0nAs/qp1LSHg4LXtEWS+Y4dTQMt6apKRhvKBNozMlnWziN+fatyRwt/AMMe3uWMpZ5FeaD9J/
vDlqg51x4ZE0TQn0oc6c9pD/DEriPj+J4seSXCJZbctT153QNm3yO9Xq/LbS+zwB93ABLF4FIxH7
q64V2+8ljX6c3YL+y5zOhViCx4GKxr3E4v4HY/n0QxQ3zAzAhNSMPcMyAWkJ0WbNCoLDAHTuYR26
oVMww2Z1rHfCFuH7Z8YFega+HDCkP4pl7LExwVe7JjkQwlNAactJt7aTvLHPO9XSHerwFgFb4f4V
PWjDbr4JF9CuuAVW/5i1yUWq6+UepJbX4DlVbBh1GLVAYnOFofS6BOhyy8AXwz3HBQTpPGtTYl8o
7rxEsOaGMNEllOL6Qk7IMAkHULy/w8maLsNiq4BLvv3NJNG8b7zipTdfDfuXyCiqH75u3XgB09JQ
V2utgBoK2K6uk/ViGxhMDmnFYqgGVIqRm2VJpGcDBfTnpn7zhsPIAud3RIuv7tviYEOiXpr29VG9
rzgZkT5/JisblgNz9LoK+7AQzgiPkzR7tyvjW2miYgdu9XCCmMRGH5UCx4FAAVzESTgt4BxXK28z
X8zuclQaF5/1OxT5Vrih7UBo5571Vu9Ve5J+PQi7uXhEhZ3TnFoTksxxf859IN7VCIqPZpNDjTX4
5uQoTKxA8LWtZSKDqtxs5TMXdg1mM3aVVYT9iVgUOyt67RTmZ4a1xONMM/+l9E5YzkLR0WzglX43
UICaUaDjtuPYOyYs4Bx5N91WuDL5rxaRGGFOL4m9xWYhdaB3RFnOfst2yn9cyXKi+xWeDd+2lmkl
1kknCga3G23++rouKyGew+HEt+oIXK6KC7LYT+ASOw7MiU3KPOYrTAa1Gf8mFCalAot1MFVTTqfK
nnJH3q7H2FRI/jOxqZU6upCu6rpAyyOWJ1KuVHa049AJj+qDQ+xArqLRhQvcDzEm18kqpTJ++1xm
t9/h+q2HASj6FA+xCdo+mlTuGXH//NSEkFvwGUeBQgXriW6lpHKdoJDYhp86VZY+EHPc7X1o20jP
UvGc7YIWaz5wsg8p7sQ7PO6I6+01KZCE/sJu1yUTA7cbQR+I9YzVXc2ZN/K+m6i4BIUBK2Lg3+Bo
zh2hk5BWFCr/WReyxMwxSgs4Vpn2hZ0HV7pz9AFfXF6OdeNsdw/6ODMzpZn2vb113azPSRkHK1bL
EIxKPCnJLcZXKVFuh4E6IeY6feuCXV4HA4c0Vd7XkPKltkcyoP1c0NGgnxNsihvdyvjoGieDxBKz
KHSi/hNi6wkG7ArJUtPD1xAguxRfChD+M+O1SdxxffP83jeHrtxymP3V+AfKVrxtavwcaAUEmH3l
ZO7xsl/sXWHXgFkVGN7P+xcswN+QmqCK0rOHd4Ty8RuTSTagllJ6K7puMJB/o5ji11Ad/XzsSrGX
Q42ROgiq7RpEYjVvI6Nkapj3Xo7Wd1SCHPbYuwwD/7gtAaUROPY1QvSSt2muQcxmEwX3L3YvsKlL
SQWjzEmdeBi0MxGF2MFXX9G3msmqLzjml4qKnPzVn7yymWBgwHLPLofwNwguTbs9OLOi8CCEQPRx
nRIL1Pco0V+PmpXgOsnhcnFh9BFNK6E92KBbP7nILzNejSCJxGjorhKzB9mO+JxcgPS4k6hsxLjU
yme4JnwxPVKun+bZl6JvfJHLuzlJcIMqRo40JOKiSQ7Q3S6K/GLL5Zd5jBcjE1aBKAh5lfFRQSYc
79QxCFLKL0Ahz3gm56SiAJDJIm3KACiRW+AvzRr510BtGEYAzMlLTq3KmpUbffvlLoSakugyiFCz
E2MP+G2jNCV2mMjPipUkGKQ/uT1U2qCZW2bhf2poZVqBZPk4e4u2jrjLg1nIsgYROGvSD/3Xq7/W
NT+I2LTNX8gfdMSThvxl+VM9KPeRBLhKrCks1T9S4YFOfEho6RFSXAkXAhfNybtjuT29MSq9xfWw
SbQdX8ShHX0zXmXMp94vH9FMbsRZPtN+3VIZm6HIV8RbyxzuA+dWBHyvyg8Rn/A1xXvtye0p22vq
ffnLHNjMlBoIntctLYVxSMBY6dI4HgMTZAsfS5gfkWqTTbfvDBoQQ7L4XdyfcUr2HTbA0/nXOREY
lXDvNZmKFKfXE0jJIom7BYQfg2delja8v4o1afxnULXPleHE8m1AkxEARxriI8S76uGSGAUqaeSx
enoAMBebZBp/W+m/hfjWDHY5ScaCPI/OtdnJMw6O6C8eFr0gbrmyjBV+MHHXhi7pEjjK0zU7FzOi
hPBLc57HmF9P57JqDuCF0aTnmT6iI5W2AbQPVD9XMnwCVB/v/ZFFyjXby/b2qs4DhaUcX1sEQQao
CIZcyUGA+KW/txatg8NuFSUbo44TNGQdvBpD93dx/kZlQ4+Hl5zNWhzQbRfZD/aEFzDB9Lfyispe
L7v0jP0m8Hkbb5P7BA7Gy73Hp8dKrYJc95guqMfkUP0k9HOvnJsDqn7vZDdBN45vfDRkcZD8K0Z0
rd1H7pqPzL1hMYWnoBybhMSDH9jC/+FNV631JKR9W9b3Lout1rWDMCS488iKU+DzTBGppFBGpnBs
WAD+AhdlHxKx2KH7IDosJ96MHvcP/0kGa1hGVeXGr4FAkPBGs2Glrd0OJS0ALBvuamNJ/ksEl7YP
BKGwv88txzL6ifIBBhMKfRpd9I73QcOGE8ap+gmZeYK5ydAFhMwQAUOY3Xa78wo/bZvLrU+yQKYK
tJGGNpasxrv3meQlPXccM5C3ZiP+Iy/ax8JkaFPW0cUiy40teLuu/bfmpNfNlsORwcgXSZvkWWy4
uph1c26sLqyOpitJyqgjpENymY0Ef+q9YfO85iMz5usJuv7632BDE1qkKq5+Qf4SBtr5et2YCtNf
AmYq2bDcKXvSzquKJTMix+vzDffrmPRnS5c+CqgjOyc4WXMIeqdj4Cv2zOxoUQGqQPfMF+VI5Aeo
vucQZyrWFSeHGk7xwxI/MaF1GxjaPMN5bskCBmJ4Z3wJ2Rvjm17Qc7C1LkJFYBkSePKPFBaPvT0H
Jc4NuYdaT4gQnjV65/w4nS8eli4yeObSDJEgILiBh2ArHAIHz9c9JxP8EMhcYeih1fPGRWVEkYV2
pYIcV3gbwz9rvDw6xm8meekoZ8d9z3JkgbshG/JG3YtPHkRRYrd4RVyJHoD93FAJdeQVVFNdPz9x
gNJix8IW5t9WkTYZX5a+yUXFw0UESfie6L2lZdNfziYn2jy8kiofiIwEZ2Xu4RN29F1Nk3mGSi8/
XtXI0TXO8HUMT+EELcPHbKk5ksbaXkAhUGlDfjjE9a4WfPblKYuNSxjkJZD2UC7sH6o1WRN7NQPw
WnqnzuibA+gnq9V8g/JTEOP6GUHVArMKR3mesvWcZ1aaVmZhe4ziTXVehqvEMuQqF6V1YoL8n+tG
XUZq5NgD6eoS+fCg23GbOLahupb1CphuaVYiyscgDr8rjAK80vDCTO6qHX/evNoaDz083Nbg5tbe
ycumVP27Gf0CZHWMUIUO9DIMVgvOFWHrM3Lq7AARfuG0kFPd+7K7ddlOto6Yu7eSj2RkDxkIp2fd
lQcMJDca/dBNh121YcEhoQgornKwwDnztC35vkHCAf0eWqNJx/OxonA1S/TkhXWoPP19/DBcVYTg
ZY9b7b/PKa3+V+7Rf4VXQkmoA6cOAu2E0WJcqXo86v55xscPVmjiizuIKZkiLZO0DBJSvYzJ1TQf
RMunYQMa49HsoMBa4w88iC0Tv6XaMDLVoW97KjuUv7b1sKB0GyeOsMmBqI4sUh+n/b7toomwNHYe
8kRALs2LdNmyyYguiiGd1CkTV08G/T8u2Y4EW0qvZvlgljpSLflf+sF/KmBFK+8KNgaZT0RLiheF
v+F07X6bGLQCLVAyTs2XiErc4rP/2OS6fV13DsP/YHmAfnBGkpXRSYRZLkPJyv5Pj9Fbv78ui4/5
SFPGdfu34FOnpzmK/hx18mArsS81g+SsijBrY8f1cWnzgNLFyN7MD7zUZaF+hDPxysa4TlIGCzL8
mlPSFsmh3FkAOXM7pHLGVRACBUUF2AS2MtC+nGB1r/kmzLyuBnJXm2c3ibPvBJX6mKttgKgcDkA9
xSf3QlvPgViNcLMbsiWHa9+s9c7tHMK+Mtk5qXtOlsKLwlyGDcJMqAm7crcu7mYX5wDH5X9nyo6R
KDG6f983ftMcQ+V8Z/yFYxMtQeWoMbQWl63hAwohesNkEBxxqBaW8DbCdOu7SfIMW2HCadFRK63u
7tDTSDz1snEdfRFaNykVZK7a2KzxH/DAOLm6MKQ5lsIHphyTipONmuxFKXSqjs9YcIE0CgXaqvoY
H64ioIis7oAr+4XH5yRTKlV2UV3vn2lA7DCX1tdQHNoVsUBkrILiv1JgF+inb3XPLXwwKyYeq98j
MQTeK+fF9804mr7zHU6wXERxO1okalfvmbUwnyiD50imwYW4yxTeSnSIFet+TPfCHoENnEgm5OpK
FxbHZwJoqb+wY8jHaHQKFs87Z8dZjzxRhQc1nJtSPb0ScY6DXq3F3xdo+5P+T96M3sn7fjFkcsvU
SQQ2JiKZmrvpBMsClVGiOXyM73mClZ9Qcagse+GQKf7V8cu7DlBrYJRzlB3AE3+y3OGcuqv1h6P9
WQJlqjHKjb8F2DA1zpoNBWtHacAmDpQjsndrZ/dMORoI7O59Ql29jUo/3ujm7L56vFL5Dt7S8ACQ
+BrxhylZLY1wlxlhJqZHm4YwChNjCSfs/flUWDgAhe9Ld6XZ+g7J3ce6ju5uvnMyUXGdI65JMyB0
Je6xcZZsr6xDscnuWWbQQZbUZ+kYxS3SeM6mbQfNxu4AEJ19xYxwaYG8g3X63a4eMBUES1DHVwVm
DCth+n8YptIAhVmMVFmzOFP8zPrP9TfqmdeYJIsFlEERxD4q5XomG7rB3FKp1dIeCUPRm9yp73/U
vmgysTPlfad7CdfcIt+XU1nOmC4U6vtbKZy/dCSnDrc8CP6IijxZfsK6Nt29PwDWxcTaf4h9e5gw
Wh/qmWkrekruU/YBi+LWu9d6TszdU2A/yUBD2DrPHqZEokWulW5GJKPPcb/MPqoUz/rf60TjWlXd
eU6/VEJEhcutd1q/PPmA5imne3efTFtjx4AXAimLLwtvEiCDxZj6g2jri5bf0STzAzV0OappbeCc
/YmSzN96ILdIbvBUV+2EFq7eMgjAvvLgxrIEC0ZqcYSvC9meiKsQoyvuApAcJoyONnbEr0iPm+Np
txZA5rJZ0CyfajnQVzOxdq72pmCRHKS572EuIxu6k0DtMrDDtNiEeCVQwlYXsSMR/GAGqGlvPiw8
kMsNFLtUWzk3ffh68GOZDFkWD4CITkaD7gGAsxxFhBgcwnEBfvGjrp00qR8cEOISdJAjDVMs06JO
8M7K+PbT2KkOJyjRPL1NNpOizMyuJRn1+bvUjRkHq9T9yHkM/h5u/FdJf12FmWXQdzYvNdQU4h7S
i65s/QKnvHvVVMTfuLs78BR68uRW7N/C+jcXH5qK19e1tLhVsjAnk9vej6Org60h91JyywFB/Bzk
umEo4ugqVRVCIv5r+d6H2D3rqMZ9hPldKLdLF2WT0LAoPrwJE7L4YvaFlnNqCG/d4gkvrd6xoGWK
JPCL8Vj3tHjAqW80fcLW3U8lMNZI0tD9Bz6cp5IpMDwxakiQpGlE79/9IMQmUnUUVJR3nLKebsEE
bPUqGaMYj/w8rINzRokBPPPT+k8Fjp2b4mvpCr88mjgqIRr3UKjJ0QLGcsMGPQy1bZEW2HvwlXrK
RsjHrW+syouRd3kzIhQeapsIi4xGk2ckZMJUT2iCHGfYOSAeZAQOpVaH4fIGEF2wub/qA4imm3x6
UsuVRaSqD9APbbOcp9Ir8Hebto1HXaF1lzUX/Swwl95GHmCJKCqhvz5ICLzq+3TP1tbIg06teZTR
XSEwcI9E2IhEjgXitLz0cae7jWvuhuwBxniNDnMyerA9jtq2GtCQP3h+GJG+o2QK3qBpBIiMyBV1
qhif/YpXKymBxbJqgqTsE2Kj7nURCoV0GhS2uvPp+SzWEepQQr8yS1RZVIjaWtHT8E3/r62Y9j4g
/DhQJRIY/zGqRYGetOd58sdniQevLCr0LIGtF1MB4pcbb4qAuQxq+XaOyt/ThzdtE+wTUivDwQt6
6QhggOJ96cacEjbwIcDSlPR2gBy7IFS/jI0JRqD0Bu5kC6hf1w2H8hGO/1MbD78mdu8KO5fdP9oz
unaDsFJqm8lLJ3KgSsMAqvzW9SovW2gwTmi572svUjThdYJyRIPqIldar3EkG3JTwuLIDije6BW0
TfJ3efC3uEgIOTZsVN6Eo2k9i8hsrCnBplx98mryvjch+02tO3mu7xCO8eHkf7hwgiBFBItf6PXr
w/hipqnSA+knWCKkK7xWpyBF0Pq+ue++CyiWaDo9Qx8jwhnhbxLO40ZOOqX6wdVYNgbeuYUubddT
+lja0laauBcssRK/zEfUNyO2j7TUjd3bYXhae/CB3Y/NfNQV1zrDb3cGPgJU4F9VgRPsxHsEJ3FP
Qk6xw8nvC+wMbSwU1O4/tveVk/aOgeSxCxbI+vPlgsek1PixjZphiZLtFR9fKZTT+52oUWcSIzuq
6VmxLhtxmIouMuPDG7zSWjURQ1nUGsOzR1u4DIhCo3Yj9Q3dwML00uBz0m6+Ion4KLhPhSinnirc
92doFl4jtfeP9I5ZN6rKAFOlk8XU9H8UmobpJF3jAoziFL6b7LcOCsB29+plIpNiNzguYJNMPeLN
stjXSPq44TXnm0ExsltnMq1BDzW8MhCzy0RCdC7xXQXISf4Uai83GSVUoSefN7sumO8WwP36TfqD
SyfIuojgXuJYb1DV+9IjuEhoLxJB/HsQZp49QESyPoYMNtbMwS6Vpp6wRBmdKpBmYjBWac6o2GL2
G9CoSip2TOKSrBRgwIvtxprXuWc53AtqnY9gfGNQNJY+5Oe8UFw8ei2a2xByyCTEnTxgcMNfYwSD
er/pVmpWCQCcD2/2f9FZB9k2lm4GSVtHztyWIEjsuLnpwkP0wdQQh/oUYxMGsKiomVgx9qXCguQ4
b87qfXAwRNl1RoP19MF+kH7hRhVByVh3xIyABoofnjqJO5qSX+LvCtZ2Y5fVV3h8GAknEkBOjrd0
n8pQ7A1/0Jpa7BEi96izdVnfgDvXvbNH2JRFi69HLzPK32LOeHyFD/1PqXAJXayIQxIcWH+coibJ
241g4x59GJEhDalPxi+bCqf0Rye7EYvOVCQ+5B99/0Zx320Gsg2esHf0P8mwv63oj1WpDIEAHj0g
egaYGD9CpmiPtOMtpQU/bRVl8fc1NNN3y55KhEMOAgN7DgaI37D+jb37gtIW/F5lK+71GZK+0mSN
mYkCEYj8ps0/rus6gu40CQCd3DY+4Hvrtx3MboeZg3BrVne1J3JxYomXbL4vjRJaTNEh1YYyKf+V
r3kuhXdhNSBH247lBpZo+6DBqw7wKHgkwVzr9+2jE5ax4BmnC7WZK89NesY9FVXpNsSEGCHcQJr8
AybO6jcL8dOrwIM+FtZIFW/jt7xzd8Mh5NmcgqpojNv7xSJGduyD8Jgh9NQVfDZo8hQLQd0OPKmc
//b097bMJMIfNUjvapuvoESKrJCMEXKx7NlrvgxKh8uAYlsbQOkaPjD0nuf6QdEayAEcz6G/RjzE
JBbUIwzUtIE3ciRf2z9eGNOYqSUxqqiGPIZWj/+v4NF32J6JAeepXKgQfv5Wj/UTPN0/+/JhQI5V
+Gch+MQfCgAPMT1ztT1Noh742lW3E9DMcJxyf2IhSMubgi8XYVlAXi9zFO0Jrph4W/itwUoa83mD
FkGGNO9aDAIhGMuRiLPvlR/1+4Q5EvlAfPBRjY0qMu1Vu7acXr2kYexDSsI0jEylB4LvrS8gEu3B
j1E0Xc4yxpMvf4X1iMfxBi1gma6VCZe0oJ0/ChBQEmqceg20ermSsW7F8wC8PF/tW4uFmEuIEFbc
y1nx2a6MBET/0Pr9ke+OEzgYqxGL2XW+QMpWuHBWeQMHGCEwl2adbLJanpjbKGAlaOZuyO/ybFjN
DrqXe+qfWmIjBqMnBocfZA5kwtA68FLjaCfJ6bsQuRtABNM6MRgdB3iWUzQbQGmoJJhdmF+nW7Rx
jJKFDr8Xn4dIcoZJqleXDMkCb0l4YQWFW5ZjqwVW9S+8JmlsBdTp0pvbFS8avv3OD07lQSdqZuXe
IGzHEzr6l2rlCewsMgYY0wfzoCdYbU6+imFYBdbb6RR+8CcMZMAy7lt6QG36/bCiYmM0Xhn528tU
iTshvMN5IDImftaaWbsUKoMpW9ztQl5TbHL3oY7Mxppv4lC9raZPXl0dGsnaxZA7BAyby3J3RG2U
pbwN3C4e8MBlmURUZGl5xD7SvR7RvfY6+ZrHHTi0E0H60RUNDq0QNkh06sj8VZMrx9xW+vFUpDlw
I/ThnVyzPSpH18+45J465kjyNCVCgVzxb+AqOA2ebAVAAImAI2gx1es96wymPszTAJcdZT+tql82
2aJKRKFQ295qBMloQw2/ptxjL1F07a44wW+boDiPBHNPZH0gadVxgEtwi0qf56V+47USAqE3obQm
FQWO/TJSYb7xU92c664EPDU00Vxs18nszmJsrm0BUfr+KHBi63JdyQNKpJ53CxFWg984wUvMd66N
x2PlchtTCUTsadDTwcsL6Z0/ImLlIS3wO5Ji9qGk8XEzScFOYz6rvbaDtVnmZJutxntFsyw8KmSf
pCApU+rwO4XjUu4TzbDRLFV9uEBngF2T1AMtT/Nv/4So4xwytyqHfbbHio+uNnkCZLl5nwvOiCU+
LeTyZ1v45S1fc4tukOXqPXilkp5EnEyaw3AlmKlPf45EfywcCWSJ4tic2fWEwXQTorPfAvcD1YWS
4uW3+xh/opbBQz4jHZSSDhGWveWc5I4ksXUK+NgTLn/sPnMVXg5S6k1/vgGX5MzpiQG9FdBiHGO+
xMYZ7iQwlyxR/3XzGySMLuefhaZIJhZf5W5D8GxGBDa0C703DO0poWbC6tlBW+QviGv2cY6macMl
NegnLgSnNECS9l7q7jTvb3QzpvkPM9Qs/dP9vIj8XNiz47c5DmKVN6dukP0ZlpxVkD6aDUGCUMPD
7cvpYM2dMVxXGxTzNUUL1SPCsmJHOJEmGY2PQKWMnfocRGH9i+AulXOtW9Olvafe67ihu4tCeq2x
3lkjeG5gkrnucE3vW9NctkXxp7iwEkq978PAHvPEuSFps0JZyun3u2pV0wDhIpN66IogXH8gvE/P
dIWkxQZySRJsDd8HcII8YtlBfmMBr7LIY01YplqRvzGslljWrHgx6GyUKuV1eqPfBd8F8QfBSwh3
cj/yIHjXUzmnVN31DHKLQK4IoJCTieiJ+22UxZy9dxlbnufIqCovgekJNisxMVNNVgHRZYLhGjSP
VGYHVJLiTj/t3j3N6MER/av3k7m0Z5JTMC41kyEICL7M3amXJ1F9OTm+onKxarqG9h4pC3f8ugCJ
vMa53ChWEdKUOFYnE/5A8FBV/rv0rdwU+w6IbQC7rIA26KpJgnGw1k69kA+zQzIgIG9A0HTgIqhX
MNbqgfWBdjzFUnUKxaVgLp90I0ruXsaz5XBcps1K6K0YGkgzJmPkuBFJJx7n16pdqgvor7Btw2W4
5b95F4+N1W+Dp+ROyAwU+NK/Xn97W5oBRoO5h/owIFgK975qL5oLnxyELTArxl6f4H2ZAcsnuFMu
s3uR8efxmnPZ5JUOdT6CcRu7qyzaM3Sc0+h6VKoBm72uJgTb10EyT2jJ8PmPtTLREvR0da4FAlO7
3GTM4ZlPRC/z6sj08ZNO9cR+HoV1zPJakylIvXTTo8pLnVXI1PZM7dXN0wOGycrf4wCNvHLqoJt1
Q0O9ncxGvPat7jtBYxCPJR7c8M3FI6WZdh34OFxbtF79U1YRjdz1GmoRx85K+hGDBdJ/vgoLuYR9
zu/5L7geBTRHBpPRRql7Fq0DoFgtknCYX99Y+ejeCpndH1U4MefUD8K3blWQiOKll1G1jGmyzAz8
z+edEe6VMStTvSZ2HIagFuVs+SWftYDRaFevH3lZdwS7Pg4uK1p15ghfRY5RE6rvAjk+9zughlXC
Kn9wrJ31vT9n/BGElPCNDkwdjWpj/AU/yHtpmy1K5y2S1sng0+ZCcOSKzx1i++ZSLzDLceuFWZVj
Zfs4sGsM6IAt0trv+xgCy5q8QVDEf1L1vYYNhEDHep2uxbMV7fFXm60M7Gfs2RwvdLaM/Q17h+2J
cSzc8bIl5056SUkEMFsnm5JemjVxkJS/RJb5Jv/w9e8B04ik1mf0xxrjwwJ+XiVldN9IAGIKQBkt
aQiCC9ApXlgzEdeTDXZO1mvr6z5sNE2vEig8HGMsvEnhmOdiU3PC+iJfirSDo5cIUVUANU/xO4Md
D58eBM6Y19u3wZs5+lncNKn0EBzwLW3djV8HuWx5VgTbfPvka9OZtalEuIlw6G2qU5QmU+E5wSWN
0RgDC3E5gfxdqXS15QGInM5Ghk2dZ+zU7P1nERQHLBErTSdbNOQ2ILZ/7Gi9aqC0+I+GwcoWV0Ny
MUJe7AjFTzw7IC1DGoqh0ow6y35bGvKBnMBYZJohmLr4L5E7YDLbT90aP3E88zatCzuQlJNf5JnT
eA0/B75Qsz9chDcq3VDQtfv1tCeQ6f4RaO40JLF5rMF3Zp+pNOsdQgf5+ahrEBnieIGK41Qk5KMQ
T80aZGc3l1rXx9/2EiVMMr3OSvPS0i+oYGB7sEFR8Kh/mn3nThPxEVI1xa3E7RwJIACBOVCF/TC0
FnrOi7ysSeDNGcvwLnyuKzWg+md4jrMBE9Pl8hLkKUPQ37IEfFYL0SKk7AyNvP+kXY+hT1NGwCGl
7SLg9z3PWDMgSR3/JLl8sY8ueiz7Ny06D9hGXHAjhpNHvp+gZ9BHjASexhozUpaxBrzQHZHtLeNE
vpnTQFVKxY9STIzhKzd8j52LF0rzknUQsQnBnAs1vz9AGlU0MULChSm/EsbVcIeSSbvPN3xxrSaK
AOWsA9enu4SaPlNQabYwYySsa1kiiPJrQ/2gfSnUWfyctYgC8TSXHxKAaIjbUNYVSpJabhMWDNvF
23Z8p8hzNgpoxJ8np6bbRQ9Hd9qrP4RIYzHstlqd5DLyzpyjSTPCMEG62i14jWMHh5wE2w0XvWm9
mlZyzYmjIrjn/B3Eh5e+/wmbtltxhFxal7+F+OS13MeN8+py45C27ZHDGhEGDuakB3ltPcSvMwwg
KNEiKyftx6LM+omzpojsnbYxIth0mKXqJfIYsVQi7btU0wmXEQUuR2zvWN6HD4BNOg+dJYmMx3sY
rhJHvsN2JfejiJYS7jTe8+DofO7GzEuzLPId/oYEUcpX+jLGe4KltGzhhdY1R8N9tdqp/QuJ7mE2
CHddv1W1vCXXAd+/HWlNyHxJq91S0TkOCj77HJ5SUEmmnjDrdv8/+HKqUolbXBF/AvUHQN6mJshW
u7nyQaiA2zBNjUx5YuKcxL+letNIGbtGe+PGoxQaA0Qe2jgfSvil9QsNnvblPxthEXrMFbQqiFhO
SwaiVxINyQv1vVWQM/kK5zo1AjFdFkIM5ABAGSryfsQ2ucjcHinXdBSdeA0VU/PxpZPrvWA3JXjc
9L9em6zdDLS2rrJDX9eSdOZGkUTkVK5vk+4ii7yaoawzdPkmHRmMset2F14lCoYzB7AzFINEW6e/
qK49eYTlpf488onROBtWTmuG6SdYaYRKqcjZm2c+lo7JDpbqg6GKWMd5iqKxUk5WoJvQ7CJ13AF7
T/dJkKxqPtx0S69ciZ7E4cziXHRfed+L1SQ31NaaVZnNZuUFMzB56APBQDZ0Myezm8441l9nlrvt
YHD/3agpvv2cBNazsQgzy0BTeC5BxIRVbmpiDVEHvSjqzFn/eAZBP/5DIDQDaaDVJhBdVBpbAt2i
prjsBFaAK93QAJEPKZuYdD/Fpg2RiXH0XO/y7RtGTFdGEofgF6MbBgl+e0FzMKYBC/DmzZ1VFqFr
NLyuMcsidoDv++awK94vE6c0x7VxwPg1lxyjU0zuxYH94cGWvLDwIvKxWw9LFsKyEVZeUuNrKEYz
dUAs3zd0EjHoPCIRM1frewwl6D9ghQ/3kF0vMyCD0XWnJSSDt8LfFCUruNTSpWS0kuxtf8xkw7HM
2DurXUaO4vhNDyRYyHEG7vxZ1Yjw5tzOwAhacIwt1ZWGUsqJkQ/KzXvrrUdcERw0CkG+ua3PT2r2
/hzYRLBhVs7tq6NieLRWsdyLZ6TnUrvdUxjgUMfCtWfMixeP1kI2XEkAqWzIk8lMJlItdCtRPZbX
FtqSKgjzjyf8RtepiAcSawco2FO5aYxpxkaoR+DRW6KhGkYSklIIzp1TxBqw1w0fiirrKq09dx/2
5MGVrUOb5FVr8aY0tl3RER66uz8MmnSb7v8FrxVO8Yu+wfR5hQ22eLJCg1O0cUxEgawdJrkEqaOX
kaSyKPi04VATH8NRMXjAZNRoI3QpV80+eWBNsRHBaXcK7r47+g1eWA5HyWSH9IQ9F7sDrus0unjU
XfRdCyxoB+lOqwvhpyyKMn3+/vw8DaoOB4RwNqYGqyqWogYCkDwFFo7KTfgjUrLjhMjN3ZOt9asn
ejMgzvesGukqb00tBJRjrGcMLetTinjB4VPwFpe0RLby0SdbEDwm/uPfw2zN1ktrN9UfOFAzWhUG
ZyE4BduPxNg2KyPIf8RV073tbZkpcTMHyIzgmTr3Kp5FZBKT3iceuGUJe0JFTGQeAKZUvah87Zz3
fdjCc7Dj+/xtwtY+15CWiOu55T/xJtnexJLMsrdS/RSIPrr9zS6dyywB5SmFpcJKDnN5m4IJatCA
Y4ACRDQoXZQoPbdTCTSBG2fjzeNcx0wwoE32GP74oC37EwzfSroD1B7vVYFB4zY597+kt6PZVwmd
lswd7MAEBze6mqioqE7QXBfhfeB9bfiZq2I5oEmwTkBd7vYN79zywyO8EtfgxamA2C+uuVitNU7r
7wpo9LIxNgNEyd9ffMpZEE/X8KFVumniWJSMsMMDLKVO3eSnZxwEE61xyh5VjVOjPhqXOA7QWdN3
piOipHdsgxEeXip0b6qWYlDz8x0Ynsl+nNYhjm4IFIcuCsotN1ZwVgrJIDHDl9m6RT3IWtG2l+I3
zipfsHMNgcwGReJoJWdXuqwWpkplImCqdP8TsMQqvP/ja04Su0Gj484qM9YPaK3vLUluxXIhuvgy
TDymkUFXKRvM920wIS+JIPp1NuAZ3tWJhgKToG0rtIrIlosUr7Lpfi2U4A6J/h+6KYzM59PqcqUx
dRyKyVzNBEAbUD3aRyx1YsLUX9P/NZWrF8UIrxxl3JzJEGITj5MItogVzxXjsP+O4GcprLVlPXRA
kcx4trupsXUBbEwaM/ZF/pUriJRfsu7sDOtgfZcKQanVbQU0M+0Abrrnmh9VB3JhStCWj9ZxJRRq
lOLM4D1PgEIv3USi5OHAvyrNyJS3o41Ma3Z6G/cs6ZXeAMXI0edvAaBp+YN4XSr8DmUGsIA8gX8M
w0/2WtKYftRhzPv+RSClmOm1XbBi5koV/TfDHzyuFxxkzOAZjtYz0C3qwkchQLlIvksEjoBOOWH1
7DJTIGut3uXyRMqBcOBk6HmITQI2eRXFNP9+iwRjm57nSwd7DPAmFhx7IBARR8qghRG9Y0bSvmnd
G5SJnzA554YmZHwXgCzwJ44jMwkvEVs3J2qveSw/QfZ9dhLlhDY3hvTg5lmRRTPd0K/gQ/wZE8l4
WoVOFvxq4I7g0M3LZicXD1PcADjb6NGXQCCrBk2L9Lo2sbNfcZFMVGkqh7d28nCyUMnOhfNq2tAI
L8O62s/6+/0oDGJiKk85O1E8jUKPZvWYDtZSwt6imrFfza7d55dRDOaDiFVfETGA9y0XAkN7ciU3
nvlHqPMsOy/0PuM8SWATKPlKizRQjwvFH5LGsGYwQWxXMNxx/LhpgErSL3FzxK1thVmHC4lm4rX7
uaVih2V1HGK9BBi4Bos1b1b8SOn7CRBbV9+mMx8iz+CooI6U+S/DIcDc5iJG8UMJeNbPdlnAxqsL
P7wDjJbzaiX94Ms5WbqsLGMtVWuSJ2T89fbfArc+CgFDx6pwgpJFkxhrVXHWRphv6nrxXWPb8ov4
+sLf3tzwUyug7UxT9CvCVO8h/eCANCIwlI3VFpA84dRrmOYkrfkNOchmXsKKSHntEXHN4Xfz7Ee0
5+yZuONwKaocCXZys+r161Z6ZbV960q2Yacdnaz8mcW02iLUWVh9+gNXvL9HykpICeFqr0GinlMc
HC9tHy/eklBh2QtBTeT35aezGvJnSXpxfOeZSeuIQa24V9oHnoObjlq4fqg+cShn33KWuQuQDZnC
TP7nvImTZBifaAPc0ZFZzjwNH3KC/6XgOL1CQfIu65x6MpJNSoXzU+3LHpfMiYPm9WmrPeh3rBOM
AGtmK2QD2Ca+DIXfntWCiVH6hK+rgXZs/DbEyznfHiEHCrFHdHA+i+KGWGunpU5dNEbxIWYjllWF
m5+C6NsQqVLc+sJCvXkpLYE/9aHAwYzjLFoql2cHGIRIIxBL5v/ZDGlHTxzmz4KoCV82N9PkjL/i
QhLBpdIuZ7larHYElvFeh2puOh0La4QtrgQv8LfmWIwYza/MosUddK9TWlzJpahFYakTK56OgkGL
ugzIUlpkiLqw+srHs1dmEiB6xCvYMiWA0NuzjyBvuBV+oj4GngnP59hKWRwgbskbwoJrUNEqnNEP
XjwjP6hWtGZUDoRWC/ktlWCcojAdv2E9Uj6KEZjqqKlDvpHc9YO0A2AaVZ+ppp6Y6LvX9DJfhgam
n5Ev5nGUQqYjbjv53TOyghpPg+SXFqZj9AkeTqqVm3ZV3YQ8unQzjUFLBWBe+lQSgN4Js/p/CEU7
q0XaOdeRHIwSS9ZFrCyIgl+DTlZKuFZSE2PpFYni7IV/DVe151I+bI/8VMR+MFdaCPWFCTMKYKoP
/4stfz7UQ4F9lFvszlWEorzRtJCNal4rXuCobDPgVQlz0AG6dwRX/u43YF7NXLx8tqMA7SUWzDpI
axIaF9hgwVSUpnk3Qa6f96jHc7kuCwlKDQ2YMgRihcTrRyRGKWN2jAs8tTnd6TB+soiker4+e7W0
LHxu1FldpD8Zn1jtqeo3yRSJJB91EAQiK2/jVMvENLjJtC1QxyyCOWCGq5TZP4OAF2gDO1D5ba/P
cRnlAZOybz6RE0HxqrdcLI8Pb7xmPu6g1Ljg398BXi2mPSHqsk9Y6NbaW6eKHXpxlNS6cFpqICRO
NYV3E5JJ+ynMshje8F+JhwOpVIZD7wySWQ9VKK3qPWPH+3mGr7L5rP3qLjx5mDwd9Cgsm9ednozT
yG0m4nJ6KeKjRqP3UKDrbTIba/UmFFqAHbcS7mZtAcaSrF0WAPRPN/cFgB1Soq5QujX1zQwVVzYi
ZuyJQVlsAf+lyAmsTIhc3/Gzhs3rTqYOZ5wUw3pgunSxDKQRwQYYz6wv0fj/3VXHBNLdTnmuD9EI
IflQJGlge9wA24b1ZSI8veaqhGf3pg5PxaiW5Xqcbt23mACfwfupuHG3EVOWFjII8nDd994yQ8Yu
J/ruzk7riPDfFT422yApVnsN6bbg39rNEkFthSIOfgq5RxpX/ePRYgk+Qi8MJ45xgjESeZ2BM8ZD
MlCT6c14w4XKl0cg7+05IDlmn02a9lDW7h7yZ8XxVJfwuTvxZHNjpR/yjOq74NnjNsIrqfCwKh8Q
byseBILzbLfOmROHsJC4tJoQJl5bVFXc+3ea/nQ2TEod7lNnnTFY0SNtk/d2u612iwolzLjwM69X
uLbXtqHEMf3M4YixDdkwWYw4rebgsno6q9oZAbo8VZ/9KivaumR+JGcX/hK7NhAHKcrnaU5mgd21
lryB6yipvPDoVY0BFFA7b5lOJ6zyFkxu7geS4oxlD2m3vxzahK/3hnTj16JywCs1s7jBhKRXYpKl
So+iV0VRCR9GVQN6Reqm3Wfj5OA2DJesH5eKBA4cGNgpiD4+Q/TYUjKKP60AL7wCGGupnLb68Ozn
OMe5BBo437sQ13DFcE51HgU6tsAnlLqAHgYfixJIkDYCHZRp9cV4cETA3ee9YnGFiYY+X3qt5lQy
76dTjIRmSytYU2d0H/NmiM8JtztgEZ7hyeN4dSER6ZqdILZ49QzAvGwMeg3mbqx9wlHYUphNQmTl
j1NAIKzGpvKwYL6P9qLJHhwMHo4G06D/7+Eux35kIIlaPfCT6yxgthG1uoyFd/KHWFMUTOJgtVZI
KsgLi16r7Ze88NsEOxpmR3mtDjyQFQl9AQwZYEMmJMVPsK92B6WaFy8CCmFooBGE9lDlala9fRO9
9Oy5YfiJ+YTnV2rOLAIpdi5+oJ64aEZqP0f0+z8FaQW1e3+k0tqhjCAmL2vM5AIvFhjBI0SO0X1G
/IrhdtXrJkO7KaPiHkDtM7Hjw9KKezaOs5nmDgYVLXYc2cc47A5mak+fj+ZufG8iWCmioa3SVkZi
QW1mrQ0Br5cPxQYQ1K8VSnfbs0/1X8hcRI3ozqd6rtn5PQdeUv6TD5cVPbWgtjWphZBl5PG5MWGN
Neze6HvgyWceMrMVZTtH9Dbv/ygbZ8QWy2TlJD+hFLkF4XORobWZ0Rb8HP9t7PprwHmUidCi/bFm
9+ss5y3DzB7PxRZtO2hkWYvW/4DsgzJyOs+ZweYSbsojMG0/IvgDQq3HEdjrgNSv42aMWCkI+UL+
JoffesS73ygG0bmrFsGryB69ReLzPTqPxt7YT68L6WhXjB2P8+rBJGa7ogosCFuXOowgCfTiOSni
Bs/8NQZgp/EGcncI4rw6gDdM7YS/gD34XZ97NJQU7lrUsYJZUSQrgQ8/eklebLJHvfAHsiXpM0aq
6PBmYOhEPOovLil5qGKeAndBAC8/MdzgstN1WH4GmfqnIeVlXV1RPqcRdUZ9CqTasg13sE4WAL7v
QksckmRfKswM55w8UA3Yo08DMQcHXNIk/Z21+ySNnwa3xy0wjRNdColb3oHVfNIeAt0KhDZZY+OC
9zr/HUFjitr2aXgNnsBU0BZUJU/fAxW/k+2zE9HoNZWwzWTG96l1wRAig7rURk3o3R2rcgZmd+ku
3MTPV5jYhZxAdLY54IgcmjCvqaKwG1IHR30DWIvu0ytKvaXDViZoEe6ewXiTCC4TuxZehHEOX4mZ
TM4bzZDCHh7lY+pqm5cSnWSyVAoaq3BVskbBbDD1rRG8uXtY82kF7lMpzwN0bRSugLe+Vad3kKeR
74LK1ilgiIq0QXBIX4RhEZqkqL5Bow5Nc7HrGK7TtIUrs9WV4DC6qRJAcHDokzVLjb+7tGdp6tnU
rj0FyLeRfauj5X7jZMOVI57UzoE3QkAJq9Y0VoBkRYvrMnkXxQZOc98GGHufu25PZr9xo4vZSQfj
1d1NACNlx1F94uwAN1fmSWbkQ+fwppZO52aWvMgZ42ZbZeWWs92Lnm3ovmV6giA4KzrVtW5IGU9a
QNRHFm4P84M954UBvUd16LI9T8bz3LWqTdCoUTrApZxb7khjZ8GAi4jxknhIVyYHta+8tGKASudQ
Siw4E8ASEfpSl4QVMF7xg2XTQR7GOO7LnxcPKe+SL4NMQEKjKuyOHn9JO7NQBbwrPwPXRyi/iF1m
FZhhNXAP7cdVJwxvLa1VHKyk09J7cBLqia9BSfNamEcLihJruECu3EC7ukGzBvgm1hepDXWFNy6/
1OlWYDsSIwzuFK+xe0UGU9VUz3tcV8cpAbc4JDBaGE02Ef3zezqYeVsZyx7jvj9dQU08/oprjQKo
rxOTeRkxvTQwpMJkWty1Y7wsMWA30Rrn7Yyls8Y/JQm3G/9HIFr/53rwROzr24wTvBuHG85L1Qzn
pYhC21xTZoEXQRr8fRmkasJV5yVjRR2I5VEZyCpDweC3ZRcHQbo6MHLPtIjSTFKCV+kb/Wq+KrMv
dXbvRMDsltUoU+9jJf9FQPNw3FIxEiMXG2gK3BhxH2QwnPbK23Jxd9eisLveLsmGruEC3r4kk1ZH
AAcfZ8YUU7oy+wylyqTZoMfzseUFo7E/GDZo6Q1XhxPmJcSXTLLLWle5Kwibrvk0rXdaetgV1zt/
3KH3nsWZCZFFj8g78SjyA1RsIeLBHNi9/DzzgGFDj1NX4MLRVyGV7mNE6StbBtqepOY43oZnLxW/
52ug7idmcLt0x0OwFYsgqpRFEUCbi1AUTRwOm0n2+mUJCLN2zbEG0N1ZKa65begFWgKwPFHUStgY
dOfVGyOCo/qaMZuWmgQs7Gy99+hOEKt5ODNYd4iUmQTuQSXxmlh8EBvdZhK3geojva+7TbSBOWo1
++3YO7FMs3CMLZLX7B1CHTobPG0oKmkNpMxp+RFnbnfdgq2ZTBgUtyXih2HpMT/SZDoH84Yp6i50
DnMxUZbHsfmTHJMY0d8cucSE/xREeX4CVtYMwycmaCAcrrjX7dl8vJ4FB6ScnPttP8YPgxIqSn30
e49ycbM6N6jQmMniVJqYlwCv
`protect end_protected
