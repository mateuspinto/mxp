��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���莑3ːz~�H�{j8���_L���-Z�|S)�\Ίy�:�W�!s��z�>��1��G?��Iղ�\M}���䫮x�S��`E�̨(�k����K�B�E�s{S6�b�0�*^.�IP{�be7v�����잡x����d A�07�:��U�"m��mN�Ӄ3�����~����-hs،G�0���sk}�l1�B%\+���L��l�~��u+���m��jBX�V�K�)���7�S3����̭��mٯ�e;[GPO�ՠ�y�g�U�͂�6�tA�ۜ1�0Y�����2"}Η��2Kig��W��ќ�[�ŏ��;ܤ�;�	�uJ6�̈y������q��_��:ř�C����s~����"�`Pѿ{���8 �jQ&p�0?q_��6I�l�`�P�Ɯ\�8o���֙j������ն�����WB�?,��O��U�aP�x/�pvw.j\?2-���ݳP�ۘ"X��w�=�{5������i�2�����l�;�Y���oPRL\e��;�G���	X����l6�	[Xm�8�h	|��XA�X'�:�WJ��i���27SQ%C'\2��n6n������p�g���.�_Kϐ�l�:c¨6|��a�$�HM��Z݁X���x�o�F��c��5�k?ձ5��{߄�cp�����a�o���2��w���"��� ,�4��/�qD�b3�h�W��/�]QVӫ5�p��a�A��[��h"l�
�
=�G�KVVe|;���#��^�|>ԇ����R��c3�_�i�����	|(�O�?r��3�3��e�B�5Қ)���d:���ڌD����(J�7`F���@v��x�:?Yh�J��(��A{S�V�~u�)�Ea����闝I�u�����P6���ҋ��O�~Y%d�i�4ZS�I#&ݪ{��߆�ֳpGn�!�Ҟ\�L"�c��Yu;�8�6s�9I8���aL��*2a%�A�&w�T�h�gN&�/NwtzQVjTp�'��2�"g���h�*��7;0�Z������ ��X�M�/-»����G����o��#b���
%�.�B�^\�@js�$��k�J� ���<�PHE��ڥ'7���ذ����`~��!Q��Ć�:M ���_*�Є��Y�
<!t|�>%�Z��J�*������>�<���]���l����x������K*m4�s���-�I9�m�o˭~�11��U@O<���e��}׭q1�����ۙ�z��e��^2���N�z!�Y��&}Ds�i`7�V�j��P3�|$dM+�(�k��e7��Ӗ�	����~A�A�1�(��0,c��d�]�ۜ����:'��
5rߎ?h��~�ʽ��`*��d��sTz��`��'y�|���w�O���k77G��ﻭ�5���4Gb���}n�΃���f"�D�>�}L���ô㟅?��sjݘ��oz��qb�z��&@s�c��J��	`�z$��)\��ըVaa��J�A�p�_+�)�8�S�)ߘ.g�|A~T��j n�M�u�@f/":s��&�6 (����C�U۲d�z[�%L�=
ݯ���e� ���h^��ׯJ�:M����&B�//u���F)��4�,�3z��$q	w"�Yd�l7u�N�J�Okvk�	~�¼�MY�o��w��]W_r���7(7Ax4P�BC�ΊIP$0��p��;��S�g	Vc���&ْ��6e�.4�^���&Gy�?�w�*�)�6��yl#��J��HS�{d����*s80z�1NC~^�G:��i�a9K4s�P>��,Z|��Pz���X�OrQ?�w\��Cz��{�H�q8���z�����/i�z�����������fٳ�;�[e��)��'�� �U�P=��gu	5):�?S���{ ���@,�J�u���A�m�k%�Q�+�=w#���iM���%�KҖ�ؿ�7v�rKf�N9}([Ӽ�*E嫙+����l�������eL��'�*���l���!�28���f��D$[]
J"�V>�
T��>�:��U��F�
V���J33.���(T��]�+�����]���xX���}Ôp�+j�)���N�������\y�� �Qhh�%����Ʋ^Z:��U�Of�9���oY��%|`���3u+���H�s�m�	}�~��$�EK�ٕ�4��oU;�ǣ��Q�,��'A���M$H�'i���*kB�B5��}��j�3X�9�}Y:��D���FJa��_�!GT+`^RJ�a\bb�>o�εR�K�L�hf��D�H4���� %l��-V���+!����19���n�#!��%�.Z�Wnޙ����_v�6j�e9�*�G��n���`!��o:��y�t�?����ˮ���(ju�>�qM�jR�rˑ���5�_W�t&"����ϏZ�1�����J�� ��'iM��Y���ǵ���K��A�%V�R*||��cp5����IkK&��.�V�/K��t~P ��p�<b34!��+"o^�WD[@��6�Jџ���k� o�q;������B��/���P��8��fN�����'���x�a�pF�݁#�Z@��uԋ�*9�@�t.8�nuoz���,!��I��p�O[���S�̀�0{�˔(O�#V���K�4Rx�-�vҗCM���Xr4PGE�\��.��L�'m�Z\�c{���<۰�Z����~�IU0l�%����1��*��P^;+�c:�ya%թr����`���Ǆ���,E���w�cLZ��7-���� ��>O~5����-z`qH��Q�+��C�t#�~pl-$0�[��	�2�e�#��n��r�q	���ٷ�85A o��)$ > �7�yݖ�ײ���/$�z�R�vɇ��F���- y*I�yea�C9zwu����/���܃v�;��S��k�d���pz��9�M��&pP���@��M� /�t��%�b %{^�O��_�l�'vv���ӣ�t��BT_����o� o��y5[z�����ӥ����
��N���\!'�h�\I�ϧ8yu�C{:h,0��X 2U�ZQT�kBq��< "���%R����IybN���Z���C$�(���D����#�L��U5��)D�3M�����х�~0?�c���c/�L��|ش8s!�m{�*���"�{���N!�'��@=�[�gU�����ͿQ�h�	�#�	�ea�^a�tLeY�h�A�SJM�z�4M��>��'<ّ��WZ�5��_^�)w6����������TLB��GU�ъ}����1���)�} 9�jy�
�GҊ2�Vf32��Mɿ4�����e������u{�J۰iu�ޏµ`�`�'d��������:�	9癆�5��_H�J0��Pg_�����F]�� wjʙp�t��-�Nɳ�L$�����
�vw.\�;�nAϝ&�Ww�f 	��\(* P'���	ă����5��o����8t�p,9��������vr3�BE��8���H�XҊ+_����Ļ��ws�9��s�oqd��m��i�M�)��
��w���泩|�Z%�F	/؈�+��|]����g��3��D���,'.����>M&@7
|�'<�1��	K�4�gI�D����bʣ%�2���k�y~���Y���́�Ң�q�RHwó�eo���L�o�.�۴����y���S��7�15_�`U�)
|c)�P>�K���.�w��`hD�^���Z�Q�M����"Wӌ�� -���Rz�����G�R~(=�˽���Po��Ճv��i���9M�� o��Pc��A���9�lq���U�e����ޜ��_��r��F0L���dl
�͢��dJ�8�4�}��|�ɣř��iN�ĥe�xy�R����ЩC�E,?h��yB�w��}/�����I������U/���9U�.(�m���G�/Ჴ5��/�q��H=42%��/��\�g�F֛͑�ֶ�.�#�O��ltW�_9���0{"Κ"s�pS��w&�����7�n�v7%�WGA|o����K����PY�/?���`���!��h'y?��5�N��^%JJ�����J�gA������#����q�Gĺ)��u��	�T��ۉ��}����GWs�I�Z=_�FZ=Z`ӲC�׵����~�TJ�R��^3grݹ������,>	�n%[W�KhM9��C /�c�������r���`�(��&�^Qs���(���J�ւu��f�I�H�`fⳒ�<*�=V5~ĻV��.�]9s�c3tN�&�z~.d�#�1�r�B��5�2�+a��D��U1D)�5���N��T*~	0����٨�wyzqV��m��z�RF8|���i��ۋ��h[���S����� �r�ѥ��U��0M��U�r�� �2�z5���8#R�cB����f�6V~RL���7��y��&
�[3�9��@U9��9���R��ʡm��YG�2�ڃM��-�&g�TG��wo�۩�v/ϯ��9�FQ�leaV�ߘz���x�T����S*4���F�TM�����4�y^n�J�{.|N
�zùU�VS�>�P��W��t6>QJ����^B�vu1�7�O��Б-ٱ�ۈ>��O#0��� �j�D�ci����3��>�[����OAڛ�xmA)''��/�}��FG��DFFe{��[4$�*�_8?�K���Z��֮| ��ta��i'�$4�`F�5�o���T�cN/�o��4��
��p����;/�����V?|,�.?�y5���@5�����A-�1��o=���WW��f��e��K��*�ՓJӶS��ȺH����嬕jz�$��}�x�V��"0���71�ێd�s�=Mm����Ε�������M8��١�0衈���A8��A�5�y��j@&�m��L�WR��U4<��EWG���=G�xP��-/��8�N��Ky�����k����ە�F"�v/f��E4�0�Ġ��N׀cM�� �X�Do�8�{9�ޥj��b.�.��� ���i���m�g�������OԼj��:(�ı{&�#�c��K��{a�e��{8�x�oXv<�[M�閒��~�  WW;�ڎ4Ƙ�$^��Ԑ�e߻��%��Ż'%O��9�0��<q����\:�)�D�~��H���	M�����!��{C�awO�tD���1f��ݟ��}(AV"��e�5��7r�[0PG�u~pQr��?�cB�S$�&8.�:/X�ʥ�,���f�ך 	�5�V>Mحw}ގ����֘�A�pU ���ʰM��/�Zr+�o�;f5�m`Qߡo���z�AG�BȰ�],��±��e����e�F�ͻn�]�T�)��%	�v*;��t�0���J'F@_g���
O;�Sz��o��5�����/���>�a��ᢜ�Op"�6cU�O����<E�xk#���Jg���$�QW���L��*�����U����DA��G�<m��� �~��7�e�Y�H>�0;h�7`t>2�R�儖��mGB�x��7� ʖ�+t�$���h:���h����'�YOp�\���R�~�c�*p�2]���`��Q��S��`MC�7j���N��.QPφ���H�|�������������E����{I��l���ŵ}N%����t �*�*:KB�[	rx�v�2M�b#�m$u��Q�k�,3�������9�>�OT 1�?f�!b��Ҧ�� ��+�\���rx�.��� �m�!���s�{�(�`�-�����e����]���X��$b�
�2 .^`K}�qЧ0/pF&��)j�>YL�Cgv�-�A����}h����!�62n��?�`E��v��P@�1�添�ȀA��0�ҎG�A`���xA҇���� �������㦿����)��g�!�1�X7Y�~�4��j�Vxô��f�ym�EE+��@�a�b��5�P�3�%N�[�3V4[x�=��H�"����o����k\H�b ����G}E��=��ږ�x���*�Ϫ��bˁ�d��R�|�S��dg�V�Z*�}m������2��r:��j�\�\���?2E�Z�Ӂ)vķA����9>���t�֎�7�՘3���Q��˗�@8��}[�[wo����|�Z�R��Y{n�æ�Ճ�̆�n��	�ʎ��f���Gr4C�o
�w
`�}��n��gQ��d�l���l�i;��.��8��S�1"�ݑ���'畋��;.>�E���"�6(��woe�^F�	���gx!:�s.fht���v���[D����	:
�]a�Je��i9Q������z+NM�sP��;��+"rg�� ��뛿� �^�`ަ�	����]�[��3�Q����ț�s��)�1���"Ԣ�GKX�LȺ:�6��Xu\\�+�=C��j6�B�Ԭ���xﲠ◩G ';*J�`����T�4���r�>5��̈́g��/�N'�{�'�e�1GQ;+�	}��^,����!Q�V6��sy��Ύ
@��&��;���t���&s��$�#�va������i���d�,C���TE�WO%�A��/���"ފ�:%�^������;Ō7d��N�������qՓ�D�sФ ����]�W7�j�eM�h�?K��%~yN�����VCsP�(_���]����gO�5	��p����c0�s ̺�������N?d�`��|�`5�Ѝ�o�~����h�/��v��<{��R��Ȕ`dR�ǫ�7���<4bv� Kh��m��?��:�ezt�2�w���ȆTZB�	w0\=Da�P#.z|wp|�����8���f���s2S�ŀPB#n���b�ud�kR������0�\{�,E�,����;k0�Z�-N�V� �J����
�S���:�>��~���g��J���=:	#R��:�H�F|���nٔK~eJ4�Կ��۴F:��M�0���c�e6�5�]����'�Y��e�����>7\��"�v809��¨5
����zR�\,	�x��xci�T�'
w��.*8#�,��Yg|��\Jom��l�sW�Jo�{m3MP�m�,R*=�0�����J
��W���"�:�|;u�K�]��j�FW^~��p�����w̼�_��j�Bc0U��g%����=Qo�3lMB
��O���$���0�
s��7%	�zQb_�Z�Y��r!*^���W�wn@�nT��#�拉^pЯ./�2bM��%���m��6H(��a��UK�ʣ�z��t��wZ��Zw8�	a
c;o�"�z���v0��&�G+�8�V�|�wR Ա(ؐƩ}�τ�k�l?p,�x�y\K�xtz#;X.x�;�3��s������_t�0mM��?��b��{����^%�}u�I�w*�u��ԷW�b�Af��5E�&��g�}��T��R���=I7i�ї��9�h�9���;�D���(���v���i�ǉ��g����a�6��q�����IMil����t|���ˆ:�z�����l�I�)��ZU�@^;Q�}�'�iL�]���������^MϷV� �����Y軫@ћ7������ z�� fV�f:0���k�e%'����_Y��M~w�=��C�JE����?t��`�(D����%͜�pIԉN�$��
q��n�� o��&m0I|��,)i`�l6��&q�;=�F�1�GL�ۙ{/�1c냯�
X
uNð�~����^>n��LC-e�S�$�ck)D;�#8�l�!�ړGK�=n���*yq���lW�� ��:���oX��b|�>�W(|�&��S̭��a}��&������b%�Ƃ1Ag�A�0��g�7�_ԣ�AM���J�H��G�b�rI ���;�~������M钤 �B 4���z�4YY7u8a��ʖ��YF2νE%��G��'��<9a�\�4��|��~���bM�U�����ZczL��]�r�m�� &��Ô\C�f,ǖ1��;\�Jt[E���)瑊���^5�f�񈏷6{4��ב�:��jd�he�]X����役�eĜH�fr�ѫ��v5����ȑ'$#��mu7�����#�ҫF!7�x�ȾU�B�[�$�w`:1,��W�׻�E I[��ɟ�F�����)V�
����X#H�Hk�Ɯyy��x����"b]�/Q���tŬ�cn�oD����I��§�m���Y�S�����j��:e˥�3{��]@�q�n6�]�AE��t���� �2��^��"�Ǜ��酿��p��G��hl8k�� IOD%#	H"��jX���	F����x[f1�v����\
V���ʷ�]�8N,^<��Pf{H��/����Q��Q�PoR:3�s����9^�I�d���F(rq�u]b�����jc�R��T[�2L�8?z1aNUI.����չ���,)ǲ�숪?�?��?�_�M�"S`���J�Q>�.#�T���i|�/�Uw~�|����D���iwق���Q�'��y� ��H�^ϓ��XYP9'9*�8�_p�W3R�}9��A��:���o��vK� ��oaa�l�,Dv�M�c��Z��E��y������^�ݠ$��|96(S_l�ΖM��4��5ߠ[N��ڥB6�]�~	T���Φ+�z�m��j���8�U��FV7r�����Qh	�_�[�UT�+�s)���*��U�M0s�����#��vt���v��3��]�O�c�wz>2i�䯪R9 ���r50��
�'q�:�]�^�_��Ѽ;)Ѽ�z��c:�T[R�L�2�F�����-��������Q���2���`��ŧ����7�����{M�8�h��(���
;�������n��$p�3Ńb!͟�(�d�^/�M�{��ܥ�D������H�2��')q �zr!`j�!�8n��d��9�3)��BF�J��&��-�SEpG�&�B�)�\�4�8�l_�.wLbv�9^q�<���;,2�V�`f�-���2��}!�1�6<$!�C%�è9Z&>ϛ�̗�U�{ڥz�~��Y6eH�eZ�{0[_�;�{�)S|^�S�R\�����p���=+\��ѷz ԟ~m�\���,w�TD	>��5��%}��]5j+a���Hj�k�_�E���~���axb^;��ra°��O��ͪ%.
����$ �>����\�K<��ϋ�V�4<VoQC.�W'8�%�H�5}����~�	m�F�h��"ж�OSS7s]i	��H`:nf|��w�W�G�Z���R�pj�}X�����77EsWs�+!�[��%A=��c#�|u�T�v5&@|$���x�"�3��o)���� �"���տ翝�����i�q��N���C_E�sJ4v���u��}
b�1uY��̬G ���D�uW�$��mЖˬ���输�lL�ݫJ:��'0=E�r�������A��C�O	lY��:�{���h�4���V��]sf��{���(h=r��
��4�a 8�����|�A������؈ ��K)z��C �_��\/���n�%|���<)�:̕�uZ��B2~�x]F�%9�v���G���;Z��h()��a��B�(�)@�Jl3D�p4����䤦Z~6��I"��R�-���j{�	���g>n�vO�c	&B$;��˥�)�I�8:�({|�����`qG|�S8+l:p���zb��c�������Z����,��#D�֑˦��4��u␮�퇺t��{�/��� W�A���R��3�����aVl�{�	� �8�����xc��~�=m]�"f[�{ujjf+��@����F��7&��
5�����gG�4��-����nG��zT�!��Z��J��|��˫Q�~
P�M�%",QteLŁ�`w{Y�t��c��WUoR9�3���<䓱�Y8*Kz����&PT������>����4=:j�꧋�ȩUbJ�0�fx�j0LbJ���nE�bES��34ٌ�B$�K�Ϧ�2I���2�C9�m��5-Y-?e�n��H����hww��uQ�ؙ�O���Ĝ��ؑo��][����l��_�o�@��REhx��pL������jF�KIN�\��Z��Θ�o�f���Y&L��-3E�����ts���p� ��n� ��Sl��������ԏ�L��[�ʔ"�\���ʘ�׺;��Oj�W2% �V��	� �Ԉ?���g����E����!�z)���@_�l��M���C��$]�n�Pni_sq���a��l$�����% �����=�Ϥ�|}��{H*����̖��
������i\���%��Po1OҜ;�6��Y����c���C_b�P�u�ę�v�o���]��x8�$Yx�'l��U2�ԔR�^���9�I�R��-/�a��i��xJet�0^�P_�B��iO�65oI�Z�vu�D��j3���[��0E�\�\� -�Ї�D�.Ł�}��к�� �Vb��>�C{𬅧^��<����<�mBin�+��&�DsB���'{�@.f,O�Jx0�t\�j��:=i	�
�G���k�F�oX��y�-�gx4��;����J *Tg�Z��c�Vu��N	�����m3��OBK���#�^�Cu�;+��
P����Ed�"Z�(�`&�G.>�G��;@��~��3a���dHR���}wY�&����զ*���Ƚ�� S�UYko�=��v�}`��ڐ��]�oJ����?��O��0i�&������1���(&����)ߜJ<�GkN6�U7!D;��26��;��=2�{�GR.���!��_a�6�C�+ ��o*.@���z^
TH�Gx�>�oP*�f�.��^3n����ES�̰MY�P��89�1���>ڦ�l�}�����k�i�o/;R��j��>,�"��[�?X��[xH@(n�ڛK��g����+�_����YXI�&��u��o����N��}4�d+�}�Vp�~�\�+�z-�#�.g���L������nmE4k�l����Ke=_��eջŒ�1���]ȶ�Ч��~� z}�6U@�R1�����F�jD����uDM�Ԧ.��%_�E�c��+I�t�o�`on�C�>��FKGC����x�2F�>N:��yk��Ak�VO�D{ X����v����Gd��6��~�wޱk��::��i~{��}v��)F�;$0�ݾ�w��G�Qb)e<����NƖ��_3���&펏'<6��u��]��ٜ*�9�>̽7h�|����Y~Kt<D��Q7�R�f�bN�3�nDCef���29*֧�	�K�����u��n$.�4kRc#$��~p*��2_�n��PG�)���p!֞�5|�C�Gכ{f4�'�H��g����:����AW��:��k{��U6�Rng�������Co���}e�Nr�n! .��3� ���e������Y6�aB�=� ��+�s���Lw�T3�'�X6�֤$��YI�#*6���dL/�(���v�M��%�����L}S>���uΕ��G<�_�;���"3����e��|C����^0�)�����nS10�܅Ԋ�	L	w ���\��$�����O��S���]R�|9 �s��$�����MƎ�
M6��
�j����ۯ�Lo�{F����	P�'�zz�S\]����s׍����w�(��|y����u���El��,�ȏ���\Ĥh[��LalFē5�5*�:U��! �0�bk��=��K2�L�5$c������I��M��l
��pi�H���qA�?
�*��������I5��Z��,�{�����_����<�3v���k�=R�Z�7Mk|� B��X�����e��p�,f�����v���K�$	*��x�\��х��4&�"�Hр���jBN��~L_��z�&>��tzAQ0���v#�#p�!9Q&*�0eš�ྙD����&%"l�i��gQ�̫�t.�M��!����U*`��F����Ut��N�{�)w�����V3����qv�Q�}=���w(>�`� ��!l Shm�Qүf����@�� �WEDk-��~��8 gu2e���*����x�k��RE������MX�c{~Pũ�$	�V�Q<�hЊ�� +V^Y$�����Q%���}��kє���˨�AwC1JF����O�%O����5}|��=���85�dƘ��� ˲�1[ΥVo�\)Z&�H�C��3�`�K^�
�����w�y�d�ם�9�?%I�,C]���< � *E׆��AD#��[�w��.d�n��BT]�j3���"嘦?<�8��y��bP�p�'̢�W���}���t�q���_����dДH�h�m��3@9�ޱu#��l����N.����P�����!�r_?0��" �k!
�$3��
U\�]��ӫVmv��׻�|�Vo�`2�
Ý`�G���F_��37�����Q�<����ĩ)�K§	�F�枀R,�%�5�PĖ�jh��w����Jng[TW��.���+�N����k0}`RU���2�P�Ev}Ʀq�ј���W_)�m8Q�g�2�ߘq�s�-࿹<2�������+���	��|�^j����G�t����Z���i������~��<�y�����V�c߮�h���l�cku��J25m�q��}޾�o��M�F�Z����������1q��tj���$Y@�n���^�������@Q��>���|�&�4l���s�㕖js���oS��|m(˂G�}�����>ݬ�W�uFɴ�\�:�ߜ�_��~΄J'�Qa1{x�ތ8������ҕ���G�-<"��w�]��[��,<*����۹�6�_j��^���Nf0�m���������)�>1"�_�ז�� t������"�T���A��d7Opr�.���O����J��r�D	k�]���Vm5P�P�W��8��j��f�p�ה��d�^�"��܍Y>]u�t'�"�7�g���o�=�@���{:�kӣe��e�@C���c�R0�c���vw���p$}��f�L��|X�/�cK��Ʋ|���٦���I|I���*n���1���6���kr}Dх��f�Np�Z�E�%y�w�a�m��q�x�Ҏ[ɛ���'��1|hT�L 'W��j�M*�K�
"�@�'bઉ�u�MWHpN(��Qj;�C��D�)D8�5@�a$���ԇ���\��ʸ9$��-^ţ��ړ$A=�ִ�O�>�k����h��w��،�R����b���\����� ��JtigH3�X0��d�]Y$"�[�Y��<�z��?�??jORQ>?�fS�F�2>C��<�]���u���C]nT�¹J���Ru����Rꯃ�0��&�w�:b���]BRz���C�1a�GsS*[7~�%w1��1B͠Z.!�$>?���Xp�@Xy�����I�W�p�y.��2=�ng�DZ�E�-�n;b��t���ck�� ��e�m<	s2I�_ÅHv�[!�-��3��l�ݽ�K3x�z��ۀևyxY�Z��:�#H��Es4v���c�6�<NWyD�o@�w�`�9����q��A���@�H�I���]�Io�Ȍi�WfY�F�E�n� #��\�@�}�z<ңM�!&��<�����A$kjv�O,�F�0�iڒ�Ck����/�@s����Օߧ�J�[�%�����y�����|,B�תM���X�c��B��B�l�),�}���?��^+� ���Q�Љ(vԷz�C����+�tG���?_aq�x)x�`��\	������~�p���xB���sYG\G(?�����)2C�$u�x�2���n ~�">n����`����58]� J�8X!o�즏�.��֭)�Ϭ�rJ9-���[�;c �_����P���������	�<�wY?���v	n��K4)&�z��	0ooN	�kz����f1UxK��Ѭ�)}"&�Ĥ�����vx�Z� �5@!�H�����~�t�	c\E�N������A�'knܔ��EA��2K�m��)2���:�~;ԇY�o�iD'�Kr������M���O��B�������������Ho;���C�4��?Q!?
��f>m��������j�(�Hy�A�e~�ِK�]�
*hC���E�7�9��:<:��I�։�� �Ϊ���v��b̋X�I��<�/�YT���-{�.*���#؋�V�Ѥ;5�ߔ	I�T-�f>��B?r��׋�� uw�/L㺝!	D�LY�\����~T��r����0A����o�X�l��"5����J5��s�&�M��e�ճdV
Ta�{Q��ES���"��I��mL�j�6�IG��-68VdNq��}^�+R 삑s���F������ch5:E�<ס��E�a��'�����5���А�K��W�xc�js��ݍ_t5�4�W�п�^�(�>6S4j`�O�C�XXY|!����N��:�7髗'�F&1!X`L$b��Fxm��E���2�hg��n�a����j*� ��ƴy*m�3��!sY�[�Wn�TX��������╡�X�k����vo��ؓ����c�ζ����nD+�ŉ�@�R�Y����o�u��0��D��jr�V�ss�h���[�7�[���(.<r�k/~�!�$�$V����LEk��Ke\%=.�U�s�x��~ᇲ_R����T ���XS*��Q��K�Wo�^!�jk��R^5(�	�j�Ќ�sv�ؿ���&A����8ȷ�M�Ow�c����
��i)�q�kK.ɠ�`_7Ӹ�l���������e�'�)m<��I�Ė|t�üFۥ?(V-��lhF�����:������$�M�;�e^�e�������-p2�L�]��]f<�o��_<x�M��+9��3MܕM�7&!m�)-��߈��د��Y��
�p�L�~�O%�iqeJ��������xV�;V���-Z�E+{�7�U�����%3z��Z$�)��W��BFe�2�x\�@y6PHz~<���73N�c�^[�.B$�9�/M��şN�26)sLZ�q�9[��	�F� tN�:��7͋)���ᶰ�dwO�?��d MӁ�ҋ&Py)��L��k�� �J��6ytd��Dbr�Nq�͎i�sJ]�����p�:� �����~���U����B@�UK�����b�]�p�(4���	U=��O3d0Ȫj��0�i��  ��_e�����;��?<�s
��q^|Y����/�w3��<��P������lO�.���zF�S_�ן@ \<�^����)^U�9�h��k�C��j�f�H��@U:���m�*A�:n.L++^Կf͹�*�H�7H�m8��並�ߖ�6��-�LLTcZq�A/!�m�^�^�ѩ������=��6�8e����Xx�<*��lJ�!�J�;D.�4���K�%�=l�&c��0��xU�������!�\��j�i x���v�w��{��=�9���[#X�\�{/+}��X����&�Ïܜ���+�����`���[K����*���d��N��D���̩�S%n;40�sg��<x?*�m� w���":�����!�{Y���8&�F>Hb�;�ͱ	�B�dL	����eG�	p��F�Pv�'LUཱིc�>����R���1�ɞ���NJ����o8��o^��G���c'���������o�y��"5�p)V��Ġ��p=�L���au�E�-�=S��Ī��b���-�2h'q�� ��z��I8�Tu�)�B�g��K����4{z�?��]�N~���D�`b�&X+^��K&lA���r� t���F�Z,2d�=�!-o=�ø�Y�syMx��z�cB,֋�.(�������cu)�Q�Y`�xȺ��aђ=��j�g��b���M�m�����Ɲ���xbJ����a]m�&�ǯۘ���ތhԊ������#����������e�D����`�͉�b,)�ó�-i$H��6Ҵ����(�۩t$T+J�ʰ<�OK��/vVY���PxJ�w�e���Q��C�~;�F
$��m�
��D�G
5�����v�1BY����bӦ�t��YAf�oXV�2���s����`v��TiiT��g��Ě:�������la�+MJ�f�P��VKj���]�W&iF�d,�s�i䅵�ڋM緫����r(K'�<�V�	R&X�qΰU�+]}'�7��K֩aN�Q�~.j��O!���ܝ+)�m +����l��{=��.��9��(�eZ�ZJQ�WoI;���x:�~q%���˲v1B]�5(n<��a�1��3�HL�_/�,�	�w�+������*�8k��DK#]Sw�Wd����d
��@��5̧l�t��6\9�i�lgXX��p�����ÛG�ښ�|?�v�H��"S5%�~Zh���]��A(`������Z=��I�c�D�-iӐH�Ӈ���lO-VW6i�>��#�;��~�K�8I�a�7�l�6C��e���4����<��[</v�>4�5V���&�h:�1���R��p^����8��	j0o^ �V�Q&��I��k>��R(4�z���ã���.�_6� Bj�2�]O3�(q�@z9簐������OZ.��ԚG�|}�Q�UΣ@�Ib���-�B��N��(�HA��BV}}33-�I��ut� �=�9�+:�u��gh�$@���m�J�+)��R�
�&�
U%�˾jRYB7H\��bc���O���{�?%<���Tl�t��os�Q5\��m��~q/i�|oMfNS7�*X��v�ǜ�)�v�S�ʿgt�z3�
�6
}Uw��J�?�wg?�>�kP-��lnK�� B���H{����OQv��tx��W� �p�<�LDS��0#��Θ�ӹ�ܡC��N��˥9k���qG�s��>7���g�=!?P�T<żBR�[ǹ���LW��v�l�Ֆ��~e�W��,���є�or��v���i1��f%.��3y:I�.Z9���y��.�TG�P&ޢ�G���,�5i����>B;����ļ��'3e;��u�fh���Dxtl�Y������=|��:��5�;�j�^������Q�h{�xxI1z㚠��|GB�����GPa�� 2��9�6�!A�7�[�/r�@^�H��9�/7�"-l��m��;��	k��|E�E�,�<��������*7*`n��^f���>@9�����?�?=uW	J�Ђ�������&�y~⾵l74�Z,,n�nm�s�|l�n)�2o��a�b��y��쪶7o:���[���V�˹i]~#Iaĕ�����(hQJ�9��O�/+Va�{�Jc^����c���MN`d��>#�� N���ڽ�/��|��5�'���g��kpy2CG���Y�lI�J�XW��O�s�q��sK�Q�tL�-g���E\�i-�#Ů$NGʰ%�'a���,:c"+��ұ�N��~�q�)�j�~ ���������055���oQ�C�>*Y�"�s�Uv��n�����HVUۭ��2~�co�j�Y��9�dk�*;�`d�J�fP�G�R��g+�i��Wl�+�����W`
Ęy�+�pUQ9�Px�‵�^��b:W7��^�H�i�2d<������+�$Ɣis����K���F��[����A��S���?j�E��U��ʩ�w���&�2�r���w�vXN�N�I�%�Mn�`����D�dj?�פ,���T+�=mN������1�_(��W*�#�0�:��<u��~�;�烼HS-Є	a���|��S��G
o�'�,[(�Jbݵ���c���o]l���#���e�����J<.��!�{���C�#���;t�����ߋH����E5����~�GI�aoz�O�/tŸ�C�Ʈ!��SO쓤Jq�����v��d����!+!-���U��(n�9ɬ�X��Bib
�2�(G�|��2{���XZ^t�k�0������&��A���:qx���:w*��<�[�⃁:]��9n*s���	��_��~�yӧ,$'c�� >b�bq|G1������U'^z���YdJ"h��A����L��M����
�l��>l#��(���Ü,s�o��H��d��/�'�M�GAO�jb�� ��wcgA�3����o;_�w8�Rf�Mk҆_g��ܣ7@�)+�dŦ�X3�����n�hc����L�+:����Մ�Q�۷�{|iɉ�d{6��iW	,J��1��'QU�
�c��
G��Ϩ��/l���g���Y���sdj�P\i���jjV�9�G���@鮕�������N��/*��6CE_T54��.1�o/ ��T��U�.aeB�\��kbK�{Az���w?/�_U�(k����&����x��6���s��!p����|a�չ�Y)��V֔ `g>;u�	<���b7�t��v�-KƑlG�%�Lɬ~`�'��T 6�q��iLse?�4+���{�Gǅkb.t�k�Fo���&�x���4Tx����Ypp(b^4�_F�k�5ʷm�sw��^��ѵ�1;�Z��IMދ��di���Ō�3�x�D��U\��ݘ��;�s@4�����5�	����5r�oS̢��s�¦L�kx����t؏O1���|P�U�M�MV�Ao��ݏI�8�R`�?��U���D�`u�s(e+x�ށ�q�(,�<Hc�X��R��w���j��;�}g	�wI��@pYG�����E��\*)5)��$i���M�����Xm$h�\�g��Me|�!k�t=:IP���y/h��G�#po<tTY6JHS�N�J���n�N6����4X�t���O�Mٺ�J!�	\U�(Z�㙨Ϫ�P��V�UP�<���,*>� [�7\u
O�<xx������]�.��۫����nD�*�[�"S��ZɎ����]aWl�3!�P>i��L4
m{�����W�#�f�thn�r`�-�Z����N��|{�O{l����fr3w���
t���s��K3��f�|-��̜#ٷeT6}ւG�&����6�=O��$4���|5�����瑻� ��hHR�4/g�g�f[��,�V�fؼtS��&���XݲnW��Vh�Y�M���
#����D(�����!� �����;��]��da��9i�lMCa�4��l�u/'��7H�d6��]V jX Z_�+���>�Ml�F0�GE� pf�;;�|4)G}r	Q-�~ ��@={F�V��3����!��g�C�u�6F����I�bl�λ~b-Uz�k/�[!���w�޸�SV��rԺq����DEU��`ػm�6��G]2(e�↊"���`I|�3(b`�)
�ض��r��|/s7T��|(�)�����a4iԝ:?ZI9�h���.�܃��.�B��u��7��#���L7�f!=C��v�Ϡ,�5ZAg�f�(fR����A����x��q�b�S��
�(�����ᖗ�ڐ�/��I�$��k��ޔ�D�ɕ��Dk^��Tݫ�Mь���.<����;aR�i�~�m��$B�S#_����E"��6������B��H]�	��	
�t�4;\�T(�=y�|���>�Xbf��	�pN;�|MxJ[��M�6MAZskF�ZX��{MH��7qt��Ś'���E��};�|�/��L�ڂ�D	<��J ��mt�m �ۧ=����V�Or0!N��+�L5]w��� �3Xr���8�)��>F��J��i�-�_��$����j��}��d����U�p�X�%��X��u+��GE�I&%>���� ����8q�{��%5w���aԽҍU�����M��w96b��
�&���N'���%��<t͊��Aa�p�RG�q�`e6<Q�L��ng+y��9�C�#�b?b�Cq��ʎ�{��L�?+�����=�j�m@��;�ݝ�t>+p�$	T��K�!Q"�s,E�'qD������u��5=`�{�h)�
��N���(-�V����0�l9��]�=��HTW��LD��	nGiGa�� {T��J��n���J:����A���@�5e1d�Ј�$9�ʇ{�Ǧ�ժS"�J�� �
J�����[�2��)���<{
�$����$t�lb"U;��Q��	:�sb6%���y�?��P�MvG/'b�/�J��Z�����1�'���
B˕�l�u��a�M
[*jJ��8S4z�&�f΅�"��LV�葑
d������4�#��Re�g;�fg���v_ݯ��$��x���QeUj��/yT�/��+�=-�0�1GN2��bN#� J�ݳ���s���׾�#�Xy�-*�C��z��(t�����痼|����It�hx*D{!K�v��!~{��=��w��=5�f��� �9툒�8P7�3[�'����\-d���4d��H�ټ?@��A
��C��5��õ�\՘��y"4	�w<��V����F"~b��EB���̄����N�r�u��R���b��dׄ�xj��ӭ�-&�/����3���U�^ Y=�tHg�����-SZ �IPDf��3ޗ�s25�&���9��Ֆ�HB}����V�f�.��[q_��"3�z��V@r孑r�$�Z2��H���K�+쮳n���y+R'��H�M�]�x-���ƽ�k����Rߞ@���!�Dį�ϒ����?�e@����:1\z�-z�b3�c���C����P�׳뛆s�;�{��,"�ù��>+��P������\���*I�%s�U��H�?q��=�}�f�G/�}�jc*��}NFs<XR>Z�&�?j/>3BE^�*Ir&%k���P������2`���k�2
T�re*�X��Y,���D]o�9g������O�`Tgҗ�A�J~9�J�_����������B��.3-�����g�t����<<�B��h��|����B^�Lyă���6��������/����XÛ��E#�Jiʳ�=��<DB�]��P2C�ܬ�kT��bNU�.1��v���fȚL3��0���$�������3����S�2T�Z)V|�6�w�0�᫽�n%�	%����g�X�F<ꊕ�V#
�`�q+��b���]�A�b�qp�j�����	�wt�n˖/����[�I�+{�t_�H�_�s��:P(���)m�U�]�v����nw�=��m�����m�fa������y3>7)��u�"��-��.j�,��f�^@�n�\ha�������>WFR:Z_!�]�S!գb)v��Rg�HLh����<Fg���܀}��d�"t�lZh���9V���C
?-9B�����?y� �ʴ�:[��~�����+����CW4&�4�!gJBܞ���a�RKe�\�\*�M�`j͞��d�',.+�>��@�a�,������	?�㈀`�!KZ_Uc�	D��5+��(,Kd�2����!�m������;��s�9��ݘ9��/.I���f���/�4����4�;�J�Ҁ52�z�	��Ǧ��m��ߵ'a��)1�!�)��t=�C�y��c�"�at����ű8����D`����[�F,�NZ����w�d��R~���t8���r�G�x�ex�����, @%}T-�12���U�y�Z^�>=aU�'%�}���躢����V����@	��6����B�#�9բ`ǔa�ʋ	Z#OJS��z5Ϩő�X��u�/�{,դ�8�琬b�'W���c-��Bj�Ll�Ŷ��]��-�.Sr��-,9)Հ�$�"�Y�=��E���������P)jS�9�{+��z�}
��7\ �����G�[Z���]���*�8���>� ��'a7�Z�n������'v��X�{��'�O4���Zd�����=�\F�A0��hN�p&��;��
�8��{H]s4���_����6��G� �����H6u����'L�]�U���v��Wm�:E������$�w0�k�p�m������u?���s��/P�m�E5�VCt�Y�2e1��z<��0.�t�ل�}�~*�>xisX��������0�i��ɂ�S.�{ɟ#�6�oi�8	�}Ȕv�5����O� '�ܤ�����j@�����:�
N}����:��7xw�Y����}X����'��R0��m[M5Y��L9�#�,��՚��:�H�|����;��N*?x���5�-���ӣ��Q6Y�.9�W&�ϧ|TĈ&u��,Ϟ3]���T�c|���՚$���ח����w��?�+L�+���5J�9�Gj�G����EQ}�K�"��H�u
�4d D�!��qFX�B�����
(�����ہ�g�Nn�k6\x{Cf6Ә��C�^hC�;���G/�̃ T~8����8m=ɕ�N����$��nF����9'?�>C+�ok ���N9�!�;�v:�K��D���ԨK�)8���F���B�s�5�=fY"�'�y��^G��a�w�;���Y���[�<�fC�z���I7��6J�U%�[���<Z�-�n��ŉm���m�h�[�d�Z�S�	)���p�*cR	E+v�^7��r��_1c4�{�u"�lk�N*[��d��dV�4�$쎳$={9��Gޓs�^ĩdV�"Y���~���k�,%�M�$!;�v�ѵ�VU� �*���襾��֓�m�M�K�4�4�����}_��+��g1me����T՗�G!��rK/0����͒ؿ��9�`�#]�ZY�y6�zMxsg����
���^�I��|�{�U���^��*ni�~w��3Yҽzb�9ǐ�����d�4m
�GI����������W,���n��cX+�O*Fz�u�/�A�S��d�(0�9���YyTN�δ�����s�[,�[�zv$3ܤ�%b�1��i; u�	��0���SK��G�2L���>8=L��/�]]d�;`�';<��s���tY��p1�6��ݕ�����,C�Z��E��,(T�[���g�ACt��>��0}(�Ƈ��8Oo.�g�C�ɢ���6I��$,*���exySm�&��)t0cֿk��ب�(��5>�%�6��>~]�r1k��e@�"<��@3��v	�g�BA���$G'��"]��jp�AY���~�[Bf�E ���)]v���}��}-�-M�ϲ+���UJ�@��:��Bz`��C�ϸ�9q�;\�K^ {���1�ʸ�_��i�{�{׸2��}��٤N�yG�2.q�Y�`��q�~���e����4��35Ӳ�8�K�f���C�R�Nƫ ��I=�ѫ��M���#�%{m��__�v�:�hN�>K���ʇ���d]�J���]�V���>_�
}���!�*�tBz�8nY59�<VCkx�*��{�]��N���V��lu%��������$y^���WP�-٭��Zk���A$%�總���a3�����%��rB���e=�AMs��A}T��
���"N��c���$.��@IvH��W������n�a _�����$�*(��(��H6��X��$e��N���H�SZ� ��s�Y;�������2Ɯx�/V6�����e�/�K7e�4ĔW���K���O��y�y�D�W!��MX:�k�!,g�k�jv�	�^���܉Z:<�Нv��+���\�82��y��Q��B�uV\�Yet��RA6聘w� �'>�������w�����X����ڟ�#����'a&4�+
XĲ{0ʊ+%7 5ć<��d�&.��`���`���>��0��Kz�$6���8X�Ϥ�&U2�h��Բ! Ϫ�\Dl&���3��+x�� �"�O�)H�>��':bN�n�;�?��<���'���P_A�1�~s��+���z�+�����W�����]X �FYa�hV_�*�/���� s��h�|8�J���,:8]8��0��4,�m�[��Ag8�q���I��@���|,�,s�� ���S7�D��曘���}@��q?c�uiN��5���-qK�FU8�ŝ���Љ�zr%�X:��)�Z$n��O�a~v6�h��C��QW��̿H'�oqOt�7�\�
���|��^�N�/�����dџ��F�ba͡���έP+�0-H�AB�2 6��*���(7rSM2��6i;A_�P!���t�@k�#��H�e�����`99w�������� Q�?
N{i��*��""i�=}t�g$��x����4�dT�EF�)�xiGR�-a��
�B��I�-%�������6��;�����EP�'O�h[����d��)����<�!vz]�:"��&��S� u�Ջ	��h!�_��PB�Ҝ��X�.���~� (�3?[�I
]������ͻd/~Hc�1��Ɛ�w���@<˃��^���k�d��V6�o%Ec\6H2����T��d_�k��)i5vM����
��18B�J�t̊��s�J�{�O�s��&^R�0�����)���q����Z?��"��l<c�im��WA���2�'V{|��r@0V5,�';� ���Rӗ'5d�O
�	�9��������=P�F�T=a��M����w��Զ8�s�a�Ƀ�h���Ol�W5(�h�={�fξb�������9�J,qGJ��ō�g�M�������������p�����)�PN����{D�a,`,�ڹU�
Uӹ<՝���"3]���v��$��������K�S ���X��\��R��'s�39*e�$�ʂ�#�P2ˡ��c��#����o��}�w�Hn?���X�1�������HXIP#}(�%c[�81=J_u�q�vV�x�g�0F�����/�5��g�_�e,
���9W�D	����(�j�Xo#B��NiN!̰�n�Sm{�q�G���1K7?;h���@��;`I<Zen�'���r��N͞�#u9|:\��|���-�a|��8i~2���z�L.Q)G^�訤v�tc�LpRo�]�hR#���U��Z9�˱}���e�i̹񽃔�uA&��Ӛ9�3(��vuk��TE �|"mk�gY��%bϩ8�Z"��<�]�M`�Z��ʞ�����cVA+�brC�<~ϕ.��ͅ6�Ǻ L�D������hX2Ҡ�/<�tr���d�l�I�qٵ��R�xe���ݣ����;F�LK(�>mRXY�U'�,�������[�����{�W�(T�ѫ��Ĵ�	�f|��n�SɊ�j^ż�~s�1e��zz"�ؤpZ9&`.��ca��m7�5�n�	46�w/
�|ڋeG-pݱ0��G��g�LE��U
xGO�?H�z٢�ʐ��pVo�mД�������k@8.R��޵���-k���`زV��h�s��mv����$��J�k�&0�G�G/���U�R��z���_P�%'����T���E��e���C<���<��V��7�Z��x��\Wگ��h"L9�{ҳ  �	X�n�#Cq�YB��v`�������4���<�ȁ���R���1[�u�r_h����s=,]�V8o5�m}|Z��k�\֛�}����>�mj��}���
3�<c@?S��D�\�ɂ��*�0^ޒ{�Cǧ���Y�Q�����KLD�uj��6�G�5�E��̉޺���{eO��qB6��o���!�EnLZԊx�J�v�L�Ξ���oQ��,0n}�(�Y�ţ�9_�J�\�!V��͵p���ٲ���ۖ��r"E�$�А�p�˥z ei6o�!H������	*WY�])�g��"H4h�G���a#��,�hm@dS���Ot��9��G�Y��`��4E�/`	��hh�f\���g�QY�l��/�6Cu��G�c�ƷZG���U�KPŨ]�	P��)���0����F�{��X���#�	5 ݄�k�^^�[�=�4�~,��g�牒�@y!���$��3�G���g���D�������P��E��L�l}h���o��"rbt�4&/r_���b��m��V��i�4��<�};8�%�晻�ȳ�F���B���/�d{",�߈`[QCThY�����8`���졛�I���N��?/��AԽ������f~�~�n�j��lpQ.[O����=f��V�K_%�n�X2�����I�K�m�W����.�pmj�˞�#����-��=0�_r��B&�+Z����T��E�B���"v��ԲX	�Q�@��02��������-�a�NY#��T�q�W�MK�Jw��:
E���w�ۇ��K�gA�Q|�jSA��{|lU�f{����i��C�z�K���j3�p��S,�i�F�9��1��a����I'J�p��)�	�wtZ���2�?�i�w��o>T(<`��� ���5^�z�|l�!_�=&��
� �QKR��~�e�`MMh���o��hYM��w�><�j���Qi��cwx�	<�&<V�:)�ɲ:�8f&��d�쇵��{�ߤ.=����A��L[�=�<Qܾ9߶�EH�����?Tt�e�v�Z;�>�.[��1\��_�n8���:���cf���E�����-P8M�аS�%--1�h�bx|�'�<��6�~��Fp
,Z%
BA�T�)��A:���i���68����"� G��m�>yN��-����c�k�CXE�_�Vhm��#:L�i����S դ�$N�4�nF���/8򨦧�������}�64[�=������$��2��|����Po>SQ&��s��ӹ�*NQ�ħ, ������&����\ފ�?i�ܒlW�DԮ]ʫ��$�{;�������Rn�	�����&�C�$�H������@s/�:.ԊT� y�I䄾��}�[�=��m��.ҥ4�?Q7Mw����Ml�F2��j[�%q���T3ಮ��r*�c�&����>�0��7ܲ[L�R��ZcY%�+��\N���X� �h�P�5xb�՟hu��ji<0���?l�x�I��\oR��n��i(y�N�6��Y5���Zl#㠒�},S8dÌI����y?{Cz��m��j�`���k�
!�L����Ԗ�$yu�4P��
�>�������h_/"VB�ԁ��Nm��ulbVrE���N�10���]{��4;�����J��D�B/����CaP߄y�K�ʣ�>R�vO=�{���^�4?V�?r�˞��%=2�-�fP��8h\׾q�8�l~�`�L6���/����<����(�1E�O�Q'�I�a� eU�St�Xy��.�PF\F�96��7���J�3�b?�Ŧ)&��p2p_�k>,q�6�o�h����ᛝ�_U�;�����R��!\�����$�%֣~P�ϙ����z�?�5���U���f�B%���>*�v���D����LYd�k-A�R���{kZ%Ğ��LDxO6OH�mXħ�U=QtGw�$%��5+A"=88Dq8Ol�d@�>c'9�=������ã#�f��T�_H
��y+dʈ�?�1��d�t��u%S�ʺ�O�1�#��k}P��)��L�Zc ��߇�Å��޼~F_t�\eB"*�[ˏ�_�I����ɝb�0������I��cȬ*E<`DT*�r|#���;]�JK6��b*��ZP&Z?�Uy�?}�t�:���r�1��3�5r$7�B'�cR�!�%���X&��<4�*��\�YZb��Q!�t��X��Jõ�?c&�Ϥ���g,┪�S�?��W�oV�ޱ� 0�e�3�]� ��E��v����a�0��k.ڿu��V���t3yq�%]Ĵ��彔�-�U��kI{n�8E\\�|�k�q�!�U�j&�3�y�ț,;Dm�/Њ�Ϭ�>O �,���B6��܂]=
������[�8�I�\"s�����;�Q�"�ZC*��1�*Ic4�:Mƥs~`aK��_9�߹E,�i՜o�\t=�1 ��l;�47�X�F�p�CfZ�:q
٘1lq�R�\�����Qϗ�'ൗRn"��Gg%��s�ՔYD�� �$`�ea���J)��y��K���>l�k��6���d{���V�7�*��kl~� v]�%A�L�l�ĳ]p�!��������./���y�J�Kǜ���	Z�+��O�~�B��A����.�;p�t1� n�`��y���t� �܎�G3��k�/,���ƌ?�.{1�^�τ��t6m`,u<�j\���1��R>�l�X�2����p��'��;� 8J	7�;
�q�s�5
�B@�`�n;"	YVm`,���l ��b�?�l��y����r�|�9��{�B+|�h*5�|�ϳ�`ώ�/An��#�#?$�m@7�����/q#�N����b�7
p��y�O�~�H�9�!�Q_g>LO������o���>�=Gz�/��Z.l��vO[�fl{G��=�b4v��>;�v��3�ţ�H�w#�G,mn��0�W�̺JL�0�m����朡h1�ߗ4n�Ҋċ�E�0*�n��`[��a�B߃�ܩ-x�6�zyr�~UB0M����r	YUH��u272�:��g�������� ��p?�aM1�1�\K���L�.��}�}r����X�Z���6�
Fab�Pd�v&?8�Wl�{袒�����X��c�9�	?O�^t_Z�Q�b�xj�d~��&[Z�$?�c�et�QpDr����2MR5�<��䓚5.�9X1d���3-�#Y:RLk�I����g�� �㌜����h�`I�!y�:��ǟ�|wQ�^m���+��>J��1�S{41�9@+��tR�q̲���nU!��vUU�q�g������&��gH� H�Q���c*��5t��k|B�&+��i����槙�mx� "��ywJ�.��q;�ji˨�ۡ��z�<������Z�#s	t�����x�FH�Zi��KRն�7r�c1R�� P�"|�VT�W�t�O:�})�lG(����莋�$=�?Ue��<��d�ը:hŒk阗�X�h��?�K�1��`��|���B�#��f�	Ɵ����T��){�\vbW uy�����'��Jo�V��V�ݜ|g^�u ���})�Dg��M��p�͘ἡ�]��n�ƗSW�<�yǖP�\������5���R[�o���;�l/�ܶ�ɿc�յ퐛�g���$��}C�}��¸ҵK��4C9#�ds�xf�)5w��~��2*tm2�R˒��*�����z-49!�Be�'��}(qi!��;Jߑ�Y��vB\G��g��jZ(⬸�=��T�?k��"��I�gm6=�w�����?u5�]��k3�N賬v�=�
,�����~�0��=P^�y�7�q�(�ްơǖ/=�ec%�I�S᳀n�J��ہn���-Z��D�X~֍2E8%��n��g���+���g-�9�`��r��	3{�ܢ� u�!�����y���u�_Ua�4���`I�-Lb��p]�;��ԝJ(\0Lu�~:~zV9����V��6AL�I���t��)����zq�]�
N��-q��X�*�b��q��/��o����*!���}aR��+3�Q?��yU1�^,*�Tjtne�i+��94���H���P�. �8+j���`�6w�j	�Bo��w��`��mC��F�0�*Ī��0&�%�偽|x*�/���D֫����o�1$���2���(�N�=������I�#��+�P������y< J�����x¼�*�Oո8�WH�](l9T���IA�0=��I+��̄�A�eq��/5,���z㙌��7OT�0|��#3�+Q����<��$�p(U8���x�K��럸\��p���J�� b������؝�� H�����`U��7�����cDu[ki��Jx��	 ��U'��JQUȞɌY�o�*>nĹ8��ڮ�qD��9�I<j;��!�=oǈO�6C�nG<a`u�+�˳e%�&jR=(�Ͷ�W�����^G.������7��ڂ%<��i�J�Q��Slh?CWS����K}<v7�o�)'Qo�S��+g�-��ѯ�dK�% 49]�������a\��Ǉ0hS�<�� g/72����^��G����B�{���N�/`;�$�d�q��EN�,���.k2;�ym����C�����&j� e���)��Zy�gYa$�5�{�s�w�.�����'�+L�i���0�@L��G�Z`�?�e~\3"������ڏŃS�җK*���Q��Z��k���gAy���p̬��Ҋ=輯��A�t��	x�!��N�*����,�W�lO�f�����򭉻�s> ��z�T�x�fR����pB�)P����^*�]AǨ�9�Mg[��Cud����6����R�2r����"ͱ�(�QX����*드�ٔ9�}��~Z`�C���	k���ncF�n�*��ɛ�=҇}|G�����^�G���*����ߔT���:�6�V����g/X��9�&M!����r`;�Y�b^U�yP�a/0��@���?�p�V}v�3���y?��{Q�	�(�3<|�;2,8q�{��YbTw�B�R���݌�!P������^ͷ<q�:��`#�����0��C,�w�N���$�bC�\,Asdp.䔋�%���^�RD�^ܱg���	PC�\�K��͉�N��ߘ� պ�N��j���c��N��]�G�t������x`��V������Ә�@%y���xU<�Y��6Ez�+�)Hd�1���Eǣ��+@��i�Գ\;���/��7H'�!�I���Z�É�P���WV ��-JB"�^�5��U?(.�ɾV
Ħ�+HDg�Zֹ�p>�n���j8�Oؗ� ��Si�,�dXP� -��c�AtDI�؄�_��UCz$�!cN��隦]d�Z�;ͭ�¥Vo�eh�"�VZ12����}�A��c�KTa��6}�T���3~ׯ�]�����'�3)#a�+����!�PO^]X�J���~{�5L@��8�E��N��ͻ��;Q
�E;,Y��S�,SS�JZH-h�!�F�y��_���7�GP�B$�Ƴ��6���e_�*�r�FZ�e�l	�C�w�~O���cѐQ3=�fe�O/���O�Z�6�$���S�G(G��n"ǒW �m�=|��%t�[�\���"$j_�'�l�7�*�$�R�t��;���,.��s����I���1neC��n�|�{(�@�=8���jy��X�ozD�B��Dx�g�i#S�@���K��CF��E�H�B���ڴ�����'vDG�>�3\I^}Z�w8V^�A�wm�o�f) v��8�Pv���[���k�]���+�+$�?{'���xx���m�����u���rv�)�˦m`7����֬� �eM�|, ��k>Ҍ�Q�f
��>)jX׸,-��"�����xI���3&?�����4|����h�L�Q��In�[5AB(r�@W�Uȷe��>y�֝:ϞN��4����4	 _�MN�)�D*��U�v������6�b
He��V|��c��*������ߏ��ĩO���L�__�\'�8�����3٭�18�������K�y*ѡ��p��\i�2g�\�j��E�ӡ��\�W�(�DRs;��w2=+LI�^�OM˄�5���6���.�%�_V����Ė� ��f4z�y�ό�)���jfgY��US�<���Ǡ8���r �?���	F����wTs��j���7Ԃ��i��%]�9��t�ֿP~�vɺW��ժ�+�@;��ߚ[�1�|qzd���aY��Q#�2/Z9�co���PJ����YoU����D_�Q[:k��o	�
"m?�\P�d�G��Y�k�?v�2������$���\������rv��E2��x,]�6ۤ�X���.Mjv��	G\Y�J��ͰK&��c\�0��2�0`�/����C��c7͇���֦��E��Z���	���K��E��� �])�_���E�c���*�&4��=������z<p,��M0�έ�Ց:��=��,�o�?qg𞛛��Zr�#,��������**�3Jʅ�+R�}�:� �N}3�[����G�3��z��#�΍��{��w��7��ͦ6�{m���LݺGz1%2��ܶ^4�8#w[J�a9�0L��1�P'�w%cX鷭��`�l �h��S���G[s�u�y��X<a�DVlr��Fu��p�z';�i\#o����k=cp���+EZ�ڙ�oM��3��pB��Z� ��R�qXڣ�0�t]�<"�caʽ�6K|����mw��덼z��,��S.@g�fj	�iɔ5�B}�5��G,c����ˑ�0;��	�M��|����8ڭ㾨�$W�	*�u�����f����X��e� a�����ʒ"�M�i/A�1����W�E�/O�>�*�ja Ӻ&��t�ʢ����e��y��N�g��]&�L��6=�Q�v�P�6�A�R�$�i&�̙K�\p��>0x.����`rg�p�/�����Nn��3|Ay@�l�D�K]\���%��kӉks��:�6y��XٻX��p,�^��ݵț[�{��趧_g�K�(h3�e�X����3NO�1k����5�{QX��ސ�<��J�@�_mζT��S#Uf�y;F>7���8r�ŷ�&;����A���I�T%��T���oC7�]����+ӵ�b�D�	�L�'\W#	�^WJTk1~:grM�.���jc��g!��D{�0�sS0(<�����O��:��3�0S��tF?��J[�FϿ�_�v�Ck�Eb��w\��5��y<�Z�w3�I� t �շ��i�Me���2����Dgf���\���� ;J��&�O�g.�P��^xk;�;��c,`���}�,�Q�P��[%q�>\�:eg�����d�adfc�Xi-M�8Ž������C��Z��fW�
˜C�J����
���g�b�;b���va_)_�Ȏ	H����:7�l�j�������Q��G]�+�E�y~Ji��wN8l�͈����1�)B�֩a�M?�i���¢�!�D�w��HR*�Z����ia�\�f8%�nz:��
�W�5�V0� ��v�Tl ��;鸰�hM2����[���mUZ+d�[�W�縠���l���Q��H ��^YJ���;���
9��!l-���y�Y�.���]�P/f��r�M���)�Y�*�v(P|����stn������#�L{w}z�Q?
F��1Ѓ׫Do&�-_�+k.�((�h������,o��l��.3f��!���آ�u^�\ٛ��>�X$�8�/J��U݁�g�'�Ra��RHſ�S��:�S�6��lm]zw[�8Hx�&��DV�iƖ�����]ͭh�����y���T�9*�9k��+��Cs�lp�@3rS��*�i�/�L0�N�*L�9r�jy;�O5Bw���ߕ85��Kط$���0�=u}���"	���Wd������+r���p��l��{7C���}PK�>B�\x��To���i��������G�1�Pyʴ�2��M78�Ǿ.)c�L�j�9�XA�6�x�q&�/�!��t������H�)����'�������%vx�ۓk_�����/����년Fr�Y���ӆ*�h�w���q�������*]�鍟���U��+�Pzp��3�)��_kj��^���8 3��28�9��T���|"��L�i^�MR�|�/_�������+.�׭�(���@�t�.�v0��&}��Ul��J�8�h�7�DQK��7+a>��A0��'��r�5t��+h�j�x�t՜e��(8&�N]*�����ܟ1��W�������>@��Ԉ��׳WWk�$��2����P&*-?���\փMa��74�ц�̕�����SI�&q_l��Y���Q�
5.�H.�W�˭�~R"��g��_�>���(��^�)��@��KD`��O�>!�o]c��V�f�	+2TZ�?�3S�׿��JxO�Bl>0l�+����	�sf�ͺ�	"����7��uI���N�L���'u&#Jr���n�%�h5kK�m,��/����6�V��e�3
e�������C|$(���ͧa'E\S�ف�%REhH�}N�d��o��@�h���%n���B�F���!��QQ�*��ðܰ��\�p��\����u�6���F�<)'J�D�=��7���ʢ�L�'V{|�"��Y��Uk�)ha���8�\kѯ���M�X�����a��rΐ,?��1�L���j5{m����Zo`�qY�D6���Q}�=��u�M"�%�7MO�����31�!L�ܗ����r���'�ϟ�n)��>�"U)�l�wI�$4������ ��cWDɱ�m�,��%�x�/��B��N��о�b�wI���A/��fm���+2H�B��j���}�*k<pq�^�V���O �{?
��/$%�r�7ex<���\q��;B�U;p�Wһ�#찵Y4y�K>m��.̳r�	}1]\�Oq/Ӓ�p�z���3�#'�y=�C�p-opGK��6��BZ�U7 "�t��;F�9)��t�f�|6@|1��k��:4����Yh���i�����L-�J2��`����+2���K����+�q���	���:��<�B�`�P�<dJ8�POq�Y�����z{���\�QB�-��	�LQ��&�ۘ��{�_M;�7�N��z$UFX�w�K>�2�G��!ώ�a�	E9.&F��-ָ�)-��<IW��i'�D����/5�q+C*8աAWU;��� ��Iؽg$�c0�/b������F�ɑR	�bu8�u�����g������FCCf^���ie*�*��j�Zv�v����H+�31߅��f]�{DViO���q�c��u� ����'�N�< T6>��`հ�].�@��8/DR��;'�|P��~���b' ��^>�U��p1j���k)�)˲|
w�_�3-�+E&ɠ�i�Ej�\jL��iYn����-M\�fo�z�đv�ٜKM���?�{om�8�C�ȼ�TA��en؟�&�=�|�F�q�bdyV�� ��O[AB�G��P�Z��#�O�+����JA-~f/�v�Z*�N������f �_�#)M<5O%�ƏM��ia_mT�0�Î?]����)�2�_�~�M�h=ڽ��-M���^����Ʋ�!���,>�<v�?�ۗ[1��9��_z�g���(W����:�'����'?+�^�0Mıg_��x��H�G����x�=�S�OL�9
q� ×!ڽ�YP�0+8���vY�iE�r��(\��i�n��ɸmhRC)��J}!Ɏ��ب���#4[���o�G��OXl��~ �Hn^q����%U�:��N���:w;��V����7'� %�4��ߦ��`��K
�s������d�Gl"��	��0j��]�)��WD��!j3=�
�d� A7�n����ǋU��T��E-�R���<�#���ʣ0�t -�@��/k�|�-v�	�M��9����L�k�c;��c��R��Sy=�;���T���~z�P8��7����[���?���9�Y��3�C�l�5���T��G/��g4_@�-�1�^��=~�˂���g��ZC�7�ȝ�2v�@�ex1��/m�xҭ\M��@Q�A�4�`<v3�i.�,�޾��qG�ËK)�����Ԙ�����D -=���-���y�G7�����P�y�W�|]�g^#��4kb�6�]�仱owY���'ntW�����������s5Z�X
��9�B�]}�2�+��_�O\�X�G1j�T��i��
��O=� N�˗)����ҤC�xE�=�l���n�Z�rnG��*}�r�m�tDَ�(M3ov[8�$��6�C)M�P����Q� 0�\�TVi����آ��ѰS��4�$��x������ë2'�>~.���&3�"��{�fZ�|9Āެs�W�KZ&�Z�����y����	쮱�jG�Y[<���n�'����I��ӵu�Ѥ���4Cv�'��;�'��f'�g���3�	xE��}\�ZJ�>&ɪ�x��V��d�q^$ʘ�21�b�~�I<�>�8�n��h�;Q�q��+��Uk��j��[�L��2�,�Z����,�����hF�a�MP�J+�o��V]��F����X˧�}
ʓ�T�����S��@�}AZߐ/����ЄvQX�5��h�f\0dإ�R��W��V�F��h�iN9�/�bI��z������*�Ԏ"�~�h=և��lPdL�.V�ۢj�������ը�Cn����b�]M4��Q�^��67SK���[��KJ�zKк�1�)����82�Uf��G=��_9@X�ҿ��^,r��~	t�:��{SK�ǅj��K�LE��&���6C�,�@% U0�A���Os�nH�?.�`�z���fe�X%���{�M����!��M ���|��5ا<tcS\o�����+Ay��o���֔�#%�'7�{�:qW�9�t�@RU�n��|-C0�A{�����Wëad;�؎�E�3����l�-F��SY�5I���@��1._(��z��)4ut��������Jwt���u��=�E7��ґ��n���2���C�>��`��r����4�Ҫ�-��7EC�2����w1Xl�*5��׏n���(�N��5d�+EA��Y=�o�ߴ�Z�S=�4�R�Db�q�Ҵ/1���Ż叠��y�
,i`���-�����f��m	]QpT�NM��vL�u���]P���ͽ�ö�*��ؕl��X
�|B�>_�T`Nϕ���O;��������1UJ#3�7j�6���߱-�11�]�y_��iY6������1��s��l�na��x�W�N��Vy�o]��cy�QӶK�D���F,7��捈�c�\��I���617���.�i)f�/��w��zLc:�NAn�
��έP͸��@ oV�ư��[�y)1��|�!AH���n;��g���Ҭa� ���s� ��4)A���n�9���G{���:R�a�m֦�W���$�+���QLf%_��ZgX&ucN��d ��Rē� �ဆhwԽ�+&Ι�����p���Y�ls��/��c��R�	�Y���`�-��b1Ξ��o���?��	$���VK%�Nt�E�з�%�ʑ�蹦���P��N�4�ݦZOڶ��S�X�+��4���ទ&�MB����� �T�Gıp����g���Y��;G��	�.�V��K�]�K|�TR*lo��oEo��dLW���~�
�ae�=v�$p� dq�D��a���rS��H����!:�9�����.B�o]У��n]�����|)��!����VeMkō͐�����(gF���r����Jt���J?-2����>u�v�/lA���$ :����I�]s�/) C9ͫ?v!�~4� �x�Q�E�B-,�W��髕�� �.4�W0�������S�Ti
o�2r
�0w=S�ߪo�������g�O�"�`�����$�<cG�pw��ڝ��;�� ^`�	�=�t}H}ZZA������g��F,��D�d�9A����
eЗ�0$�kI�*I���"Up��u�a��S@R��(E ���pڛ��ELS�P�|z��a��A'>7��#���|��3zhC��jv�%�=&��#�����VQ�'�����>��ך�aW\�	����4��C��ts��B�
��k��6� �)Y�gLs-\�Q��c}��+�UNsq����)a�u���5Mfб��0'>���)^��Xh�(՜�Ⱦ$�4�x��꓅�����6C��F�H'Κ�q��LX��~� ,��� � �����ě�X����M�P󶸶���q�ƛ/��^w�c��bz��!��$��׽�T�*lt�S;��>�u�C�H��!Y{�l�DāL��1�Ӗ� ��Da<	gD��{����c���ڋ!�6Hև�
� T��Q�N�P�i<�E\��#�٤��-�K����<ξ��@��͢1&���VX���OOy�C)�J^VE7̑�֦<����i��Vy��PC<�s�
B��R�Ì�����H��~?�����FZ���,_���\�=+�|FT�s�l�=�̀5��?۷�yd0z�"C3��g�����gS?gP���4��~&��t��I�;,2+	y@����f�҅�A�ë�(q<�,A���s4��\)rcMzO-D>v�|#c�G�U�2��P�y�c��O�C��2WuY��j)���������j|���o'��>u�r͙r���e���'���h�)JNB�Y�{�Y���nɥ�$��8!Vĸ��|X6lgA�_�n��K��3o����3�)%����|%�#ظ�>FN�j�xT�I�Ltms�+͘\������	��I��^{�O6!9�������ޗˤ�[��m�tx�|�Sd����@gW!%��8����,i7留N����"} ���sI�u��(����yGϣ�[�	(@��rQ͍�Q�:B�|7x��{𱶺5g��s��(����ե�}�$ǌ��Q¥}�e�j����`���;5L={�4�9ڄ���do���n��>@�}3̶a�CE8r l�P9N�b(�,nŗs��}���̞AW)�[������t�$x�y+qM�9�����'�Y��n��i6X�f�+���>�w�*~�㖕E)�e���r������q�.?��)F	�!tv�l�Z�- Їc����j�"��"U�k��(׀�Ou��	$nP1��n��k�4pX6M��L�-wԠ�`cW#��ˌ��������I3�W�����m����#�X*���E�~T-JZ)�RV�D�C"\�S�q1����'b��׉�]�Ւc�vkޔ���D� y�D�����do���oޒ���j���oC� ���y7�=�b�V�̕�A����%���[�Z��h��N�u��\r��:3�J� "	��!ty)�yrO�8]-�'�,8����n�,��5ҝ�Q(���gJi�F����V��*�l'��v�����9�io�z�_V��!��5����n�4�;�����&�@��t�������0��5�_'�[����إ�=/׌�N@�*���Jw���L��[�HN"�:�Q�J]k摔g��j�=����u�����.�����U��la��?�W>z]�Ց�0��]����>~p`[�x.�xK|B�r����MkI3��H�(�Gt4����0��DQ%�R�_�`j�J�Š�����X�YK�T�τ����R�§�ML	�e��	ӂ��������c���� 
X|Ѷ�r���Hi�����/���2�'�;+��s�#@�pw���DЀi�#��Mv3�D�n������n|��RS�� �v���[�Ô�Fo$&�X�s �N�g|��\���CS~���HQ��<�1��:�,���}�.��҂�mb\�9J��Έ�{X3M�@p�4)Z���˖�[h�]1f��w�F���P�V30��������+�P,����xiV�h�қC.���(����OZ&ó�5ӸV�@�$$HW����O�]d�:� V�Spq�IqM�qx�ҭ��ݎ��O�o���9Dx�QSK�M��l!�Z��~v�Ծc=U��I7�u�$��6�o�Ϊ0V�u��`��D�s+�Cg��Ǥ��Y����ـ�=W��Ք^��p�z�۰��y��1ƕ���F/��V$��֕��@(k�������=��Ī��$s{�m�z�f�V �Y�.���&�&?���`��"]�d���y�j���}}�~���=��,|�@��A�R������tnyYe� >�`�2�	�|�q����#�_��ưXɦF�1��'�����.t��N2�p-�{p��?��s����'�z����kAI�p�5�B)��3�gV�:�W$i� �T��%v%��iO^XR|�׃ڂ��� ��������)0�k_	�v���n7{:O$f�a�|"�����˶��!<ӹ�U�4-H�Ӎ�e����J-����O�eܾ �ب���9Y��$-��C�������Pq�w���C�n�1��%g�)���LB.͊�z/�C з�$��"ͼ��b�{�L�7�'��8-}!O���(���~6q~�Jr� Q��5���ߊ�Ǆ�A����r�p������2�OF�:JH��]�a$o��{c�U:��������j�z�C�a�R�tu��7����1w1ʝ� z�f��5(�(ص^��[0�e(�W�����?e���O��J��Q����bt&�8���������i�H2��W�*"i&"̯V�gI{&*�Q�Y�Q������k�N���� ;l���ʰ1͂�G��� �`Ѩ�ޒF�iak*ЍD�����Gen*�wW$�k�&4�����2�J�!�tl!vF�F
��L0�n�4��#�٫�ͰшH�}�X��:Dp	�ϡ�K��Գn5��A���o�o��!�X*��M4��*����A���3��`&˶�>2p",)��ۭ��dt����K��UmrW#��5��Ġ�Al������t!w]�$�|؁�$U��N�mn�㙍��ռ=XR�8��m�ǟ5�@��%�Ϊ|�l������Pv�0%L(*JJr�� ��=F��ܙ�[?����ե����X_���^_M�	��[zH�����,i��GH�ΧE���̓�m$n� 1i�#ה�=�Zh$l�b��ƣ���NE!�������@��U��Z�^����	���-b߿��{EЃ0�c=�Ig��? 7��	�� �J	�=Ŭ�^��+�V�siAI�EY�r���H��f#����$�c]@cy�k�Wbz}�Mi$�7�E�F2*ȁ�N����4sg=!!��s�.̢Nj���o�)Y�t.������D»��}���^�n&�K�5}|#�~A���y�Y��|�j���Q5-ڎۿk7�B}�}7�x���4�Dc<�_}Gp��+���H#��y2d�׽M.2����2A�����.j+�3�o-����W�ć�_�[m�ɻ�>����2����m`�Q��%iY�;�b�4���� ��C#4a�}��j1��@���!�u���6��"�ۂ� ����rh5Lq�hFn|�F��a�"ۨQyO =��,o�ݐK�U<ɨ^���>CI/�Oְ����[������ D�A>ߗX|�ڋ�l�*��KqRIwkJjO]�3���`�s��� �te�����x��0�X�0V�
�JUm���N�<��v������;	��>8M{紋���.�{����.�3��0���{J����V�j��<���W�2އ�9�"��ڂ�;ދ}z~�j��RĚ==��=
��%�eU�\�bT�qQ�E��PD�2�8�>A�������Q���v��6 �{c�ͳ[�p���+J�o���/�JF�w�$����]��`X��S�[s�n�O����� �u
�=�Td���� �15�H�@Z��-�	]�2��?f����"K�[l\�,����N![�:�vQӟP�����2:f��l�L�M� %Q+֍*�jW#7o��}�3f��>L/�4z/\O�����ƞR��͖3���?��8�	�{7���W���c�4��Y��ͳ,-YC�qO�]¬zL-�oy�4���=�U++������_nh���!���� ���Щ��	�H��֑kPzr8���*�ᯫ�iX��	�Ù*~���!�R��U�+�t_p[�����	2"[�Ə���̨�������b��eT��X�<3��8�������XO|��a+-���ҫg�U,�AO�n�·�6�Bj���f�*�is��m2���=����hͪՆ&qH&Y�A1��5�Z> rQ�"���pq���x)m;�?yؼ�*`�OI[��|1�3���[�,�	=��{�*֐�K�L���]�5�����I��}�����J5��
�?#ρ��r�h�8[�m:w
H'���������	�̀�pc� P�8����G�O<��G��&�x��[��!�$�P$�⎥)9b֕E��3KP�>�5H����p�~_��b�7��;]X�W(W��-ä��wb�ƅ�ͤ|����t��&�9Y�).MY���d�T�| z�����ѡ�h>Vȡ9`��yY �;��!�54�E�ґ*��q���m�g�̝�.$]�U$�� (���~{��,,�|�^͍�B��|R���֔~G�7f�̅>��@��rG��Ō��Z�!�kt�p�a�$A�@':@m󑔶�]#���	ǵ��Z���������vm�-��O	L{�qD�߆&�f�:��Йe9:�ד��K������>�@�v掁<i�鹭���],�ǁ�~���.T�KMӾ�S"�3�aw.Z�x)�w���}��Vu���8�F�&Z@��<�3�wg�N�����:"v�T�M�HZ�Y�발'���S��������+��Ft˵H��CRp�\7�yF	a@?�*� ,BE��t��9�Z��n �3=��VK��D���\�%f�,E�]���n~lq�����"w�l�i�x:vr9�}��+�j����ŧM- }_�f�����V�*���#�I��P ��@D�D���N#�EKj���
��y�-���2�/��c�uP�KN2�'����Rv9�0?��S�}�ym��AS~N!b�{��w�K�����dY5ե�
��X#��7��1��)#y�]��Ta盝�/�����)�A{��F(#h�c[����r&9[�N��oE��Tɻ�K�!�J�6��9���?���kU�4��Ų�����ƺ��^׉`'�/.D�s���!Y��� jX/$d�B��6f4Q$��LD�[�wa³�绲a�=��NQ�Ss�@�(�iC�]��Xʲ/M��ӣ��ۄ�M��6 �]��`簂�~?@cW
�k2!�@���_�!!��~/,L|d/
��	פ+XpI�uh8���T��
)����/���"���u�N/"�����P�#�z)^��]	U�������Vņ��J!�P%m�r2���$Q}Œ5��9{�YzB0�X�JS6=��/Ƥ11�؅�w�9)��Y�Q�p�Dt!~���6׈6��G�3����f�0	������N�$�C3�XW�]D����<hZ��I����ۑ��?���#� im��u�RJCx�v�]>�Ym�^�n\w�WX}�J�� ��Å�P= P9}�fH��|E���	賣]"��
��+�)9�I��TW�$6��Â��s���3��7�7��Nl=��vZ~Y�w�b��P0�O��
g�t|B�ގA�WkZ�\��!���ӝ��MP2�g)��Q2���z)�Wi?�x��� ����zO�H|�����^����Y�X%��'ϩP�l����3�?"�f�{B\��'��I�a���D�2+(��u�)�,q�ʺ��:z�`�<��I5Ĭ�5�oߨ���V��[�}Ot�4î���:3���#�i�����k�$*U\���b�a�^���h�RD�|j���Tbs�=.�ᜈlJU��B�`ՑF�i���l��A�����Q#U�(��G�,L|{{��bp�ƙ�	����Sv�,�#o(�$UE@�wPG)a��*\<O��P�x������WI���D���E̓1�'q�8�Q72�(��ya��S(��ˈp�Sk�7
_z! �,��#bki����}�Cװ��vgd������q��&)�@m!=��+��*J-$�#��(H���k�J綵�(�Tl��|�����GhTs뗨i�����EE���kb��)%�p�9zȩ*�'�z��`M���=���A�X?DK龋���<��>�h*1c����"謷�UAB�� ������)��a��t��z]����w�M([���0�U���/�����gy���Ϛ�_0�	��T��r���w���Ǒ�ل���N�K���٨���m���=��{�{�H�*v��Õ)m�4x��)�3�̈@y�s�pŇ;�^r���f�>ڭ��ex����<�gڕ�֍R�>g�g�� �1�A�H-nx2�P����]���ޞF'iծ���)�����@�!0�������2H�p�O���yFl)�5�������CX9L|-��p���~-��0e��U��5�6�9�c�6���@W��Ǿ����29�AUf��޺x$8��Y�+m�abrz#�K��lS�#��q��f�L��?�B;p	#ʏ�C���>�r��b���%�ha�
�� խm% �01����ʫ�Tn%U�4%�ؠ�9�8��������fڭ'/K�Q��)���H�+1d��e9�)�kdXP>F��o~�̟d/�LZ{]����xmx��>x���wI~j�yE+R��A0O�n�$u� f�|Sh}���U͎�SS���2m�ɱ'?���E��c�
/JȃfU��K�L`�A��7��߆,n��a�%D��f)1))�o2i��S;*��I��e���ķCC'k�i=n��~���J`�ͺe�%c�/k��~�a0D��S*��Eu�7/�"�y�������2P�n��@r4��E�,�}��$MM4^����(V!E�JOO��.�A��ܢ���Neos��r�׾w_���Z��
���@��E%��Qul�� ��%h�OP�un����Wg1�Я	�������R�ўMG��m�E��cT+�O��3@T0���ifm�3���f�ť�(����8�|YKb_3C���b��~�l�J���c�&P�X1	�9���\H�&A.U�EA'����q0����
d�(�h�E[�4��j+-q`�[�!�?X��� ��m�a�!q�wV�%�TE�5ϫ���-�"]��u:�6�n��J���
�I�NX�4R���V<�1���5��'a�������"��l�Oaϼ��x��[d�/03W���L���\�:Im�Z��_|��4��)]_EJ�th��@�R�M��yX��zC����r���-���ron�LadԷ�V�r��H��S��&��ʎ׌
�� B���xЫ�,�u�-f(�e�����^&Ƨ���X�3e?�Q��i/�+a~cfY���
��>���V��n���Y�Al{>>Q�vW�Q�V�S6��E^n�:רA���s#A<��nw"&[ ��pȦ�>5 �{�Y��a7[�*�c�r
d��c/����6u �|�z�BG�fqe�3h��:#.��:�G�8^�D��5��S���n#PŚ��g%%�=��M1ٯ��8�M���0�$~3g��G�2D\A��©	/X����4�{���?[�`��[�8p̟^?�����]ߝ.~3a�ѵ[�� ch2n�Ĝ�sQO)���Y�˕� �A�p�đ	�i��8���+x�o�����'~=sv�j�D����]Da���-C�iT��+.J�r��ف���&�9y=�ܠ��i0�13���[3���M����.V�խT��ޖ��|c�gI=Vմ�j�1��h�]n��`ѳ[��7�o+ު��@��:�p�~��8��@���N_�Hu=��[� ������ԏڣ���*HN��B/ƒc�ܳ�gۭ� ��0�?��H���{�
*8�:-tC��X!���[�\C|P:F�$�#��T����	e��A��nxC|�ĳT�I�7U2�I���rv���)`z�?gYHG����Q�G�_뾛u��:wqX	�϶69Y�0��x��Ss^�o����it��"�1�o֊���^�_��< %D��f��Nl���DF�9v���E,����RS��?	�W�
��h�ZB�>��s�N�e`��#�u�A8g�˶�;�@R"bl%ƃ ��'�EՈ�*��P4_W(K�%l�a�p���Esm�~����Ky�
�	�]�Q�Ih\h)xk��*+�F��Y�AqPn���/a�������Gf���F���ˆM�u3��C���{�i�Q�1Fݨ�ӵ�J/�4T��e�U�����%f�&�As�,���k��;�ll�=���=f>e�V)���t�9����g0PO�1ǋ�
 ���v�lyF����5��G�'R��; �u��1�#���%��q'^�߯��s+E�[�7d\5�=qs��	�[���[&-�
7�5��xg�����C�U����7|
�۰x���0V��$o <�t�Vb��� fp񙲘8��{/�����N[��n*���st�怾D�-0U/���~�ī�~%�2�\�ʘK��+��39�ᄲ~�9��"(Q4}�ԙ����ʚ�J�U,���J�m5X�g�R܋o�VE'���D��-��N��;�ںCU��0kוڑn�Ӽz�@̿���pW�����B�7�e�"��
f�Ϧ�=�al�o��sx�6��P�,�<{�uz8S!�_ۈ�y��#�d��� J�Kr�R�N��f/[@���g�V�GS�0?�� ���q��m<r	*�T�jŏJ�X�3vw^��u�F��o@N{�u���j���E�#�;��b�3�t!Bi���Q�ڡK��Z�
k�ͻW�D�����Èƾ5���$���A��Ȳ�������E��r�@����y���;O�7Y���لR�d�AL>�;A}~EYW����(P�}��
�NOqT|�d�ln_� �ŉ ������|�YVy�V���0X�Deޭ& �#xț���k	^��FY��q5�+P��\��Y��
��(�#V�8�C�#\�@05!�g����;��U9D�1y+!K�7ഃI[�&���<\0=o��ֵ��W��.�*u�w� ?�ﳮ�=nK?ʴd
��`��?���̰�m�c�!�,g�i��q���z�P�TX����2��#�8��v��5�~�n�@��6r�i��i�����Y��9�$M�9�qiQp�%���Q��.�� ��Y\4��˴x��P#�����UZ�/ih�����{Ӕ�)�u��~�ſv��̠K��E{f����&���ԭ+��e���H���AN.��q��>[SO�+����Ľ"�%��i��aE�,�U���%�°�s���F-ڤ5p%�uS�::���;:Q}�P�K7��pW��