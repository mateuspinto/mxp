XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��]�: �L�����|b;��.0͡B_'{-{<�^4����A�V�9�m�1,G���،Q�#�1��rY����y������I���ҌW/��(X��
����Z�����v+�g'GɆuK����8i�q�E�LZ�^�{�����C���w`���TE�	e��@wY��Q9z�ދ1�͇������z	.f,ώ/sls���4
X���� ����6R�T�~'�F?V���'�wxY1�I�F����)�#U��JK궉�^-a6nq�\1ug	�s�RŊ�Ք}W.�n�Gwj���V�ǂ��b���)?9^��X�Q>ႝ���s �ʨ���WyY'uQHU������C�3���	k��֕wV/�����E�O=�ϩc���4��L0��ĮƗ���eg���X���;t���hnұ%-2�>�ؤ���8���j;#��g�_��c~�ڮ�K��b���$5�I��p+.�W~th[حe��e-�3���:R�������:i���`c��,��c�퀵��!8Є�{��?%�ҧ��(��~�y-�ә����1m���Pc�����v�Ɨh��U�e���j��"���̚%�kD�gwv�@J�_��F����I����K���^�U�=)�l�gm/�i���ۍ+߇b�u_�^~��B�m�-�xͫ��S�Sj�s����zCo-$А��1�:s���|�ߧݎL��ꩤ� �r�~�	��8�EhXlxVHYEB     400     1d0� G����@�{	�|�i�Odk��Z&H��[��!�7x�� &<�*��,���+�ұ� �l�^�	O��X{l�"B�q�iO��~�%�a'y�p|#5��Oqߌ��+���}����ҝ4Z2 A$V���������n���pȺ�D�TU�,c�,�_��m�����O��;�b^boO���@�Gѻ$׊2��TY)\��B5�iaL�ς����F�f��|��yJ;��e8���0*��~G�5.Qč��.�O'���9��.�2�n�l�l�fvΗ�O)�	�J���<'"��`�T��OH��P�'d�.Ą�VQ�4�j��.ҲZm�qBMS�z4�K<R4¸fI\f0U���=W%�U��J�g�/P�n���Qs+�~����O��okey�����C����#�X�i�Ȋ�^7�)hg�5;�z�S[�)ĀJ�W�!.%��.*��.ր�S�t�XlxVHYEB     400     180*,����n�U0W��Y��p�y7�'��c�-����I�U�?���--���m�C|eP����.,�a�V�=��e^~��H��4�"��� ܲ{>�"0�����C$���&��93���>dPU^�KY��W���G?��U*������I�-ֻ �_"*�J��N���d@K-�����%<	�︉���?�o�0v�������v+* �\�	6�K[q�})�
�LV�~=��9~P=�ǯ��p�F�l�E��
h�����.�XXo˴��K_,-��<�!A�H�J�xi�N)��+�e���1k������z��n�$�5�p�
��ggb\9���E�Bm��3P�ꘚq��?9h�������q�j+l� Z�&����XlxVHYEB     400     140�ު��f|��Q��li��y{���s<+]�!<���I5&��-�/�#�p��$���2tXޢ^4Љ�	�.�nJ�"uAs�~��q,M=���X��f��f ��Ҭ�4�c��Gb�@�zC�8�aar��my_i��u�A����,������!.^����'�5�-�tD�y;u�5�n%jq(�P
h��o�8���j�8�V�}S�xgkI��\���N{�+6�#3��D��(o�)��䩔��cc,�_]�=��n	AuBG�%��`�Yf?�xz�%V�s�gz�G=:*=���aXlxVHYEB     400     110������`���d_��}��_�9x�]�uCh��W�P�$*�Ȉ�OQ���U�v5���H62����J#^�3����?��"������
������-I	?��P�騌�+�����������3
)l�~����L�GM��A����7����eS�5�i刽-K11D+���*�|l�uM�j?���do*��m�xUӋ�}^��,-Z�E|�%*�5�+�	����
����C�,KW�6ۡ����ֈY4p�d��O�¶p�o�XlxVHYEB     400     130BM0hM�Қ�ύ��n�.���|�B��	/�q�b��d�C�ŃO.�x�o�?�k�zHB�9Pٟ����Q9���w2
�7 :��8�^ P	�hm
u2ܯ?���y�
�p�8�o�D�0���H`��3��s���=�5V��6�K�+��_�����W�/�&9��-7t��$�b�5�~wh�� %�!���ΉON�Xʩ�1���LnJpi�'�1�@���r)�k�d.�q��Yt��%4L웷s��D��ƭ^AC�=@hzN��JYs�
.�@aT< ��F�ӧ�8�7�XlxVHYEB     400     150w�Ȼ|��Æ5�W�R3�܏r��F&r(��8&d��x��#��K}+$�3��u�Y�^JF����.�9�=P�hO}!ܥ�l�<j�	/�FM�>�S�_��l,ENaFFh��a:K���@�&��Χ����6<U��+M���*W<*u��K�������VZ ����+`����y��-���żi�칇]����)?fԒ7�����+B�^����ח���X}��n'P� �R�6�:
� �7�G?�5��B��M	3�������`��O$�ʲ}�X��B�6�z�V�(�pe3�v�=��)��`�����hJ�l�	�礉�&����G�XlxVHYEB     400     110��0T�2i�$!�U
oz���Az���G@>e�7{^D�{Z���Uy�f�}m���4��8�:�a`WD�Sz���9��p��*���9�;^��4
 ���&�/��i��K���nl����:�ܹ|>λć���������_���x�c�j���\���ߢ��A�O�K����H��+��^�B,���&�߳�p/|գ��q�Dj��M��a�T��xB�[��U�y�$�)'�y�I�:�,̫r&��6j��/�j�=��5�$]XlxVHYEB     400     1c0�e��TE�hԝƐ�E9X9H����9"�E�=;NM8��f�E����a�*�xM0�L���㑩Bgo��z��]�M��NQ��x$��uʽK�0�'��2hUx���<��-=6�|��ˈG����'��.xoA��v���iHS��G�r�5�m�Ùy�x���sf�,�ל��U|�´6M�������	����f��0E #��Q��)L�w{$��v�[ª���Ǻ��Vbu���}�U���͛o,0)Z��mk{	�2�w��J�ָ�y� `��cڡ[{���P�\�f�73���B#3�R�����6�u�!��XC��Tr:g+��s��4�4.��g�r�s�T1�d�I�%>_�l�F  ����ݤ��_�N������&�v-�Оf��B&�g�C����w|U���RP���XlxVHYEB     400     150$��s������;s	_�/a�+�w�������P�L��
9k�,�m6�fiʗ�zeQW{/��� �٩�DM�6?F��|ݣ�:�H�[��UD4'"�zX���lO��<fΌ��^Y�f&���i� Na�\�^�>�S@o.�U@*��@K���8�o���[�N�N���<Ig�c�����Jv�;v7���n=�E��?͟,Is��=<G�#$k�gh�CW�K���/�axE*���إx5�#Tdl:��������	�������nT��5J�v��D�Z�vf��:l/)jO�'�)�������7���#��C\tՁ�*�G�ҟ$R	�DXlxVHYEB     400     170Z��2B!\�`�dm��6'ل��Q�\X�9ۯѝ-
{ug@go1�\wH���H��Vyx������	*A3�.Q%3�����0�'} ׄn��z��"F���U<�v3s��'�b�į���}H��QE�c��?Z�rϤ��=����o��W���P�e=l�5v�w:��NFq�㽷0r)��J�M��c��gQ���r}0���h�fO	?��}s_r9Y�;@�����Ȼ>�k�疟A>Ԋk��N�'�t4�q�` ����\ sG7������G@;?������B8�:���o��d�97B
+]uu'Cg{�w�9:u�f9ƚ/<h���s�0A��]u�:yދ��9��XlxVHYEB     400     170��f��C���zSs�޽
#,"9���ם�{ߛA��ä�7�G����;����I%��V�F��₎�r0�,:��a�����z�.-<;�
!��߲��s�k/�s�Ho�&4�� �f��-����Bg��������i�h,�şO�L�&�"���P��>[8�@%V�-�����p�p;�G�	�ջ�5����nmT�3P�(�?��or-�8'@W��Ǔ�����?�&ã̷L�h�M�$�
4��~,x1�+���ّ�������l�Hw�M�\���sGv�Yڲ���2k�;���qr�� �[�Q*}���s��P{F�
ux��*���(�����^14�`�Iei��(��ׂ�4#XlxVHYEB     400     1f0�
��	$<��f���7:HQ�.�G8N�0��i���/�9fCz�f_�P���O�������&�J�`���w�$��v����S���.(˧ fV,� D�8�S}��<+z�ѵ�QJD�2&x��m���|Io��i���T�W��
�[�_��^eH�q����t�z�G>��-��a^�EU���|rY��f`��4��+!��/j|Ҽ��0�
{5/,Ǫc��R�d���������g.6�����>5�I*&� �H�P�E��TW����F��t���{�F���hd��y�O������pM}���XPJ�ӌ'8PB�'�/m=����	ѲC4Y�e�$\�8du����|tV׫�{�$�P�h��}m��,P'�&>��w��k��kʒ,)cy�yW�},���_MMf��)�:��LL2v/K�M2���rapr��S>��F,�:��1H��{�p�	X�bb�c�5�TޜJ�4V�Cսj���1]"�B���d+��XlxVHYEB     400     170�;G�I��0O�yl
���K��f�_�3�X/DЦ�v"∟HT֏�
�f鬏
.J<S���"#Xp�n�h�r��	Z^��{�r�)�2��.W�Y�I�����μ�������+(��T�?N�A*Ҥ��W�����n��F�V����W����W��d����QT�~y;�?ེ�����)݊��$��{���GH]�>�&L�
ʸ�ֱ;D�gk��Am1�<�h����CB9-kq�Ͼr
�X�{���T>~�:��zA~���ۤ;����H���P��Xg@\W`��؟g_�5�Y�K�y,`ར2+30��R�EΊ�J�6Qk@�/LR��t2��u�)�h'|zj�ݒ$*���yI�P��XlxVHYEB     400     190�8(QS�����q��-��)�H�[E� ��'ϋ�%�PTNU��|UfK��e1��O��F)g��!��P�����i�f��)��M՝�C�GO���e>� p��M�F����ݿZ��| �����)*��bs���
A����\U��&;ŏfL�찣*�R�<N�c2���nI�0����u�x�� ��,K3A��[�!0RA�����_��*5��<��UP�h���ﰻBC�0��1����}[;L�����H���db �3ێ�V����0�'��ݘ~�{�*����kB��q7.�xh�R=�
�P$1x̊���7<���м� ��9�N6��;*��j�#�����Ƀ�l��Ţ���+��01�~m@���&�m��:\�GXlxVHYEB     21f      e0�i�Ɍ�&�(dz��J�b�-��0?����vm��ѥ#��ďC�~��oQ���w��=�8��z9�j�ql�З��AGwҷ{/&�o���(I��eK�]��A�g,3��q�muu�SC��"H�u�Xo���d9����C��B77I��D�����51"�@���D��D�F���=5�)���軚$UF�P5Q�6|������RZ�/Bf����'��20]�~�+��V1�