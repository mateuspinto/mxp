`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1120)
`protect data_block
1OnTS2BvYi1UPB7DFloPJXQGFxBOZicaeFkTFcmacXTj1cKWhaC5F+Olv2BgPcUYy8LG+GqR1nlL
fbCTIjC92GrN93N6+2AdUHJ6YRwHO1XMZkiiqETgjJRKN1ppycv7dr1efna3t7nFI5d+EqWVEkJb
HmxHQPSSzKpJ0ul9HYa55HrOfR4uhys7XNeKYjleqJwuJLbYKewVpSG8/N3Q40REuaev1AMMgIy5
2b+agvSVvkoz+hG5Ae+Ex2yXiCsIlw5qEslZaLyTwnUMfLjO1d4LD+UjklwULAHFQo6b9Vkhr3qI
PUhk6IVcQP595rrnyv7wGt7WwRgtSydNwbmv4GyIrsnM9MYBEF9tiLV3jD4kNdVPHP15av43iZQj
tjVZXgfH/KlWUwPXowO4JHe/tBBa4UVgb/6P7m8NLh2U7k14p+QEKzOHbYjJpCpnStfdzQj3orvj
FdjNC9jI7zTEtlDuqxb5qVNyfT12LOLwlvFzxzZ8atjo9LdWtAEEf4mh4wzqjQFDCD8VCylyMcpw
Bl8XCMLEoAeIoO4Uy6IT7bRq+z9aJEVFYPfCXdqKt96J8Fal2C+wd1EhKcDatxdOrhbNKDKroQ0J
uMOM+HjB9WPBEjFR19Qts3RhFiV71V+Fl4kWM6qsCQi9FUJ53oqLAczE1bCGZ5CVNDW9zHWJAp+6
+eSTZGS061VJs+Jl1389g7H52WTvRRCbvlRV6WzNtY7zmO2MR5ko7/EjCRvcF1FZ0hp6BytpUuLV
eOReqZflwdkP5BiaGXjN7Ypt0tx6fnKruR6Zzo8Eo+vJpvYPHvrV2QZo0fI0YuUC911E/mXfUm9D
BDV76RIsEJsD0NJV/B4rXOL6FVuVUj7Od6vxopM2sFyKUnDDVVqZ02k+Bhe7Ec5hb0d+nRi2+U+O
+JTregghJI4UDvuBU+97hNyn28kEEyeJvaIGbulVpsbmEDlj+EuYwdqqB4Zq/N6K9dllX12Zz/I+
6GCed/iNtbB6GOZlM5pyuykBRMO+2un+1mlaudNCfGT5HeTQ/vaj6rV7ilUpwQo37KkAoS3jvvN0
WBU3DSE04p8yC6THGXqVFl2zW9UT5SzSGBHY+kwx0NT2T92hHyvTal9mva0rrkFQkZZi2mfBkYtP
MjbvdIzuA2Di9VeFQgiQl69a2FxZmBSVWmP4Onl9WatpIO0uir1kL7qRaSXTSFQWQaVU6mTgMqyp
P6YYfOQy20HVSlvOFyVNxqIWOQA3NT3X7rDIj59korNpQGWw6PamUihQW9o+pJDqERZXMBZ9b1Ar
fbs53pfZhYdKKiX8d2X2r1WfokZXZqNO3JjW+n6xUb5wrkOpBUVmHUs+jUmSreTNf3PwdZOd0D70
b0Oyh1JeRacUfxifEBEyOEnlh8OHlml4jat0Ia3Vxrzxrwe5cPN+oNIK6p3eDh70uaTSwQUw4ghn
0jmYY+G2btGxB7348ZFok+q+6GqJOYjZttbnliU30GkxC5Ds7A==
`protect end_protected
