`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12176)
`protect data_block
7vj/dezox/xw6tak7hL1nOJxnDHk1yqv0sVi6jEcPLIWbpdFS0qsreW2xc7vOluAZ8LvVciThxtP
kg3B3XmbJ11rRmXPM9no4BwPjhLk5yMmv8ygyK36NzDEFCQ70+WlaZSBNIKyJsvwK1USeilwyWHy
k5B/r8km7JGRold60NQtWe9fughNiTripXsZqsR+FB4LlRZw+Wiez018gHw8/P2pJIuAW23k17BC
WMSN7+IW5oIx7yUghVwDK4Ozi9YCnj19eS7AQQjRBqbdANY2yFxEWdSaCMIx6ybhJcdfdlxCHQwB
FikwoyPPoi/qEe3zg6OiJvXv2LA9Xl2JmblIZeYI3xVwIq+eDdGln7k5BfXYMMF+htpy0+UwJhwO
IOxyks/MMeagamSPYUxXN+fqgdtB0CV5YXqMid9yexXL3kNNYwggqjt9UwX+IkmxnKcb8UWDdRWi
ETaYo9iLmM0AL1oqqeJPmgbj6mnjLimIzJkVlgv59ble7cs/xmOHJ5UGqu1zMis11+HqdzSkadR+
ohVDwOMrxmwr82nQnWssVaTAZuaw17nCDql4aWay374W3oLG8ej5yTo1Z3bBwtVBUpksTgcjdY8b
zSqmch/TR9bypXmRKsLP+XYYUDwqdcZxyw1LZdaYt6hI5iVo07ocbbWJZ0D43SLjrhcKlMjvB6uo
/HUCHyAZnVX7y66nZVPkiMKmKNjZGMbPVGvGvPH79LHehTQGh9hvtvsJIE1fnBTNz2xqQyWcrYGy
abJ1r4xRWDbPkuxSopkv/MQXkjFTyussZmtzbS+sZywURviYw+MAp9qZM+o0u+hXyW9X/88FKI8U
TZYP++u63sxfxGxiiwE1uEe9AUG1Yzov6+cyWte+f2DPIZsT6/dVT4L9ws7DCKHJr6aGR+tCLDOW
fQgSWwzcqXPs1tu1M05lzTtQOKLGRspPIgGJnCUdPN9REgUc6Jf1A7k3W5mtnqLYa5KiVKpfmco/
XgiTvUFvdl3qY+n3xtoYxj3V+ePCo0qFOeSVqRnbfv6Xk0tnwN3JEhiMjrQYaTuf76AmrKaTA1nl
kwd2GlPlMHLC4ZKbfAxHYq/tYmhxJLxmzFPawvouR4NqZLTR7zN9xHKu+F1rJZQQJv9ZGbuhVCXO
jwH1grnhhTYNF7y+VcAGQOPB/o5Phx0qn3f6F6QNTmOPK01/7qL+6DzTmeXXw9GmjaVd4lqFuzg1
4ZCefxRIlqir9CnM2jasVz6R+qkRoU95dvCCMVFLqKnLOCdHxg/QRm/IUUTw8501icf0mtxOMj/E
yEuPt30V5QRFx4HUAil5+e09LC/WgmXvdIhgJVua42C1u+eDuBYSuAbrhPU4BW3aBo4kyQIl6vhs
806rAAXIRU19KAvgD3moTbyymh0Hg1ZIjljIchHpQSjRuiFwjWp1haSIL8bkHiFVg6kNWmQwiBq6
g2U/V/7udmrcpO6/teBUmoFpX7DKY/tM1srWOQ5743z8WEGM0OKUTZVitEbU/vxxZsxFFUvExg5f
6phWfj3a6rKQ68CuQoHVousWc7omZvmHVvHvHP/NUuP4522HVjkaMi78FKi9fUlPbXog+Awq46Q0
piHAxlFz59q3ZxUDejIBnnuwlcY8IHpB9DWrIwUNseND39ebfFim1uHdHlJlIyftxTxANRABPckN
2knpCCjPXwPwJx5FGJ99eJTYXFw9v6mjlcepXBJvimzU/OLkuTtLIOMfwMsVCYh3eb/EJgkkv43b
cImZKd0Rtnb9GwhuHySfFG+cyJiZXQz7dca7tcdKcp0yP5f4P4wWUwtvs6sIhqFtvLa74klF3leJ
r2tR0GE6B+J6POGx81r1RHKfktDDorWYq9xrfjqc3sJgvJTZ1TVB57jSsF69u/CTNMnVcSDYWDPa
VWzdUQpowxcKOowQSEeIzBaiV3AJp5ykDSCR1OgZFIVHJZFkhrk6PrlPR5l8buzgQYR+i97CPYKc
IlQsAvCFq2PFCacTTDAsbxYqTe7RKVWBULUa8RCzaF7GQU/tW50RO0uxSR73iM6h20UxriIzSBt3
jbZkrWy9daoD6rQeJAuBj2L7Wimd8bpKkaWVAa2Y049n7djLfIPvHF6tD7N3NPg73S8/5f/ZS8G/
3mZueRX61GQRhIzG89CwqPb252+74HBx65EbOuomtIBqJJJaqRB7XU3FJI943E/ga2PsyHXz92nw
/rJOigNC+VMV1nRUi91dFYVDG1CUOQbo7SnVFZ3WUz50nZxPEBo4wJgSDUyB1viUP2TH4qsKtclu
xZv0LR7qr6fMT+0pPsJEMXNeLUyaOibXXcAFYi1QQgZhp/cxiiVEvWh1vXekHFYdf4SZ1yGRY5sX
BhgoJT0yVkLRWV91BawIj9M4cfmT5ljBByayednB+H0KIKuSuufq9/THZ0DTrubA+1wQrpqayHkG
ztGpnM/k71+JSgNc83yswgFM1GRCwM6LE0FEn0SVmWLsHrH+EKzlRC85bdIbN1Ham82d75v/PK+4
lbFPw7t+qt342QbgBDhmcHUKHMlkuK6NdA5yj5dMZmVmKrTtvA2Ymr/3F9TTUqQLyCqdSTHgG1IP
9ORHTLXellRzMm5BGkyU7y+pZVRC/f8TAwx8/yPsGNGFqOw211DKhQt4l+Vz0A2P8JVgYltXQAVb
tnhxBD0UIWZjkKBjJnVPg8BSqsLHv9uwfkDCnNoM4icG3iCBr/z2D9yM8kqh3KTD0aE15SL4mKAH
X+lDUeV0P0fz5VCnCzUS8+3iYuuZ8dZWSmQjzfSsheF7md3EulablrcEBH/lZVMQpcLuNMqVGyP1
6/OEGWMZeVf14qarlw8y4TAeFzfod4pYG82+8c1XQK0ClaTNPpxcTCycCnM1PVDNEVD9S9Ws6jYh
hUHQuZHrA862fl5EWebcw+GypvICeE2m1KQtSUBzcLIYWrjLnRveehxS3eehFxOzPDzbPK7cI39E
4WzlU2JiKFhdiTQpxnH/Xx9cJHwLGLDwNsNol2xw7WgC9rjkIPTYNIm5QJcW8WKEN8g0LooUx7Dz
dHQHEBoxUeShxXUMjvKMmaBnnmlUT6D+907qIp7phLwJjX0UIhketLLZlc5rvtNZlyVhrTfXLrrp
PJ5oVI4GNCZlqYrQ0gc/1EVdkVlN+oq2AygsQZDzV+M+79QuKams5AqVYXOuSlc0vApzgvGEWlTV
iKhBdblKunIG3GffYLeBvAyCXXviY+hULGa3b4A2KgcipOGBOqBwbVP5bSFsEv7wXo1ODc6CjuQ+
Kx5+pdVxhln0QLkTkopV5Y3KGnKghvrdeIyPIFDbipaODpBTwnnPgXeTLkofQ9OU3R9dFrQB0EM3
WOssIXwBT3SGHXyDDCbMtzIzwSDHnJ/RQTb7OTExnpJgImnQCrAn+PDeLEUxnfFAhdYvwu/q6dO2
c//nJqtkr+RwKZ3qdtLuEghE+WDulhl3fYwqEUOP7p6kmQ3zHwn24AR2faIB3nXwtv5ahTdUGMNn
PrvGQZFWuBbo7RKf1IPC9BljuDcR9ao4/2hv0N+QlBgrO+R+c1ON8n+Gw0m1pOh2Q70VtbXw9p0O
KhB7DPX+sE+BhtK5irEi+YGgFnRWOCFFkgh3KrayytmI17SXcPiXJUr+G47NSQxjEDLD1gU/f1US
cMf0nlQ6yUrP0PXLis9ZLKMklMnWGDX/ov89edVOnUNFE2GTj9pgzsBpOQM5TAERp6apoJ6QupMY
+I7q8nzaooFBDyQwr/eSiozNIFBKHIZDZSi/FR607nHZY73pZSSLa2cbGuw7glYLgGblXfS//SGA
4FNvK488Vb6yDE/1QSAXMQ4XdSQ/KEUpWbNgyakJ5x4FEh9jjpw0QYL4urS3YwYRe1v7flkbT3Ph
ZEWGSxpmtKmHlfxeeBSHxbkD5j9ZS6KX+mq4Ms96pgwfYuqre6DjLv7DN1qgaEY9F1oR3OQPjuGe
tQerjxLutvhuWlCpbEkkdgs5MbX/mGOwSHTCA+q3AIo0VdOjK3jthxespVhDoG7leztpwvjVkT3V
pII1syigV3iikW27ee5udNAqqLaJOB9Ib1HMDdqxLfsD2+mXNeW14MGRAb0HSZUbjFmdkubaxuA5
piUJ5Y1VYE1e//dHICpPeaZmEl8HwTdtQtFxp7MMHibfM7RetvAnBbNdA0ng7uU0yLPJtxXGato7
LVkqGfUpkM8t5wTa1AWDvFSlT/WRwYi0KL0qFIpvZp/YpanxMj+2wOKHjn6DW+aD6GodMRoGrGKS
BFTwgdd+vP+vMGVnEllKqHjqVZG7eM2wEzZUHUGlF96++eAy1TXN+6Pc25nCmp38Ck5vC4U5SaSP
b1YrtHnU4RZGeu+LxivttzGI6wOClFoC0lJ8Elw79J5CpwNwwhSRlA8lqRTCPbjNNi75SV5Z7UoD
sn4hem+Q0SQb89lcFkkHYW16suDdY2mrqjsFzX51fnPVh8oMMZl0ZC5z8nuYuohh6qV6GJEyai+V
ditEdWRsE0BkR/gC6oxbCffNu96ZlSkOrrls0H4KGXAsHV+Ex6pOHNGs1IlZr+BNx8sGoC34wNaS
v4ovqEHPrif5i5fgcJdogA2hBgOojsNQBcXTkVwR5BLQn872urZtI30nBk/t438RhFXEIeLACP01
dNsay4mxEYpPtQhz5jP7KmPX3l3hoVYa24G8auJVTK0SOep2LmAuuUA6OXpDkfInubJKgq6Ou2V8
svqAQ7cddn9UZbOfzsZuSEm9lCqWwk6ij5ge/aUw/OuiLGgD00L+6UVIxzQvAbOG8vK5OW8fvUtv
tr484cRdqVAh2I4TBNX0/0RbU7QGzd2vSAR1X+WZMlX4gOVHgcnLzNR+syv0nIAAblpzR9XIWYfq
OGxshdaMMHdO1O//7bHtareAcTtsHXvdyTfm96e9lUB5d5HIfqd9RUG2/0wcoosfs/x+gyhn8Htb
Q8KF29jKarSU5OuwDMjGd30d4i6S3/pjM5gOWxv57mpI0JMJJT7F50KzFR9wqXAxdolVKS9jWZBA
HMSdNX/pbPXn+LRUkryCEXj7Ri0p32CzlY3oJkaBnahciwUnbBVrkb+az4iH8v1JLx9HsXliwxwq
jKlnHt5Gbr5Km47i7jQEADSr0GQaW5pAArpYl8cbly4Tfecr+Ew6HtbUNxjfEP+fVy2uXij881An
qlIeQUpvsE2xnnsmQchXfCX4xQ91e1SxIK+yMG3480k443/Fll+WK3AXcfIUSttpGTJLyBz4ds8G
QF40oGJlEnA/WthylHIFK+6mesfkuWbGOzk1gLzE2X2nXtkNv2DzUL7AVnHkAGZ7vLUrccni88Hz
nucjRUi4VDjANhFspjmtyoGTQHYyPY4ATy8vsrvQ10fkFBkVmO+A0Hkwf3eYCfzUnnTTd7IcrFxt
nlAGy7sR9oI1pqWDxaBOMrmKKY6khtaA47sHwqpSimWWGVUWogGEvvS48kR241UNNw2EI9NtQynL
eQkA1nBK+NMH/ADj3UjBGeLirktc2TwLe9ZrdAVwLNkbU97iGE2x6paeN2VvqOjyX5AgYVIj+4Ud
EzIuIrIpwbc3fuvLy4Jt8j/5MwTqYyjM8lm4vSjGm+0rWcxUq5SHST1Vxvague2j+Zh2YVpF4F8N
D9YHjIzeQ7w3bJalEwsJAAs1N6O+AippNkn5CaR0U4HCOoCWFWK60WXi6NL428sqCbiHrKKFq7T4
XRFVQ85FwKDicGcS5IJq8gTv5kzTsZmM/fOGrxEwWBmHgb/IZ/bXsgkm23TB7WrzAa1wjJ7FgwZC
dMTainDyQ13A6jGQ1OKWCO2A9XaxBO+0Xi6zY9xF2pv92B+V9c1SZbwQ3TWqHmhpDfMl6Y7b9om0
8wTtIoUtatCNYqubOzCmZdtWrh5W7OQpSM0CJcwebPtoTeY28hUK5wXuf8sLXwka6sPRuNrGDNqm
tqkEkXvD//LVRAxEvc/PpcYy+s8kv6SJSMAw4BgdxurArEp/15Lc/lAc5hji3iqaWBvVkE2qsfxn
6uq72p/ah1ocvjM7wb2wspZpwjegk2FycT/JaVNZqEvXZJwCqCAxqjA78x/s+AFBFQPzCNGv1mLO
FLp0HVwDeI2gvyiTu5nbDMld52NpTRcxSuNj38tQNXQW386ZNKaXRe1C2XsRojcgZfPYSlNOz2wz
k1Umi81SohnM9Qmc24ysbDqvmjazPX7ejqrze87LQF0e3SDqJWGudrOz5k/Pi+xbCyzZVcrs25nK
yEbn+oaiYRHuL7dfUBpPHMZIdMUkjl4nhfc9hKxRc+ZUyLDeW86MBIRwdOLKUCNak73XA1BcuONT
F/bmOA5xoZW+T1Qp3B99KqWC6QLSAos9CYgVk/BANzFoCMcE0cmlQP1oePkVd0xV7ojlXM7R7qjO
Cn9/MoIqw6ZxLt8fJoxKOtJSM0tllW4WSVvU0vgvwa5GfEC6bfs+ZfV6FAD5NV1NZHStV577fpI1
7ZIAVjPScONSyCaFjoVHpVXjXrvFGVvX0WgZkPyjfLp4vTPDR4IJ1jT8T1jXh0RG6t211hPNCC7i
ZqxSTY1Uj4eS53xHdw0y1R+YpRCMkNgcPRkw7geu4ArImgtStfAh2MsfKZ0w6Hb3M/TZG0q7kvrQ
Apd93C/yEB7t5qJmv88jUM3fifUieA/bgAW2Da4lWAq5Ux7qPQMwwsSyCidXF8cb7s1pR8LIicVK
xkEK7v9VCjYQf6xhQGK4eUDyb9QU0ooRWQqNi2hwNH2kAiv6L6WueUtYlWUpGF079tz9BTrSKHrD
bKz7D73PiIML8MoOPM2n8JTFSwoQ65kgM8GU2vY0pumta+XTcDylDWotrH6VSeiguKTdhrySZ07q
AYkDicBO6NDFQr55H+lTDm/8bN5BpMqZ4f4n/2eqk/zOCHfT6ej/wG5prW8OxnM9yxmkqdfu93vX
fp9/Wq0OFBfPlCQ0xCRvIvtqOaqUerNU8F1QzB/kqE8xbEv4BBfJVetjRCBEtCJDU4A3p6Y0BbZF
dT/vlV2myVhzCL98wMx7FrRlV8kEmpFt6QN8ACB1MytJQrc6R7qewKtWvbyFitVeHGmIgUxRGocv
E5h5b8b0YYDa7CR9ax/zbBS3LzVM1YoTACSBpAxB8c0nDXUou4gGS0KVYyCdlVPAYWJSS1a+y/bd
TGO1U2R0y+IZagqtWHUdpy0wYyUHveINJpLdI9qEkg0/tG52ZB/PZDNHOj14XVe88Nc1ORqnZb+E
m5Irw5MXVeRxiMPqXbmsGyfmsDbgTg2feqYLxBGYxsQTV2YLFg2EBaArz/zYdFG/mLORP2Bis9PS
k4D6wqSdsMXw1Dl4/pinFQMUhnHHNxQtsfpIAcHO79XAQhODUBu9jl/1K+/trCt2rJ25HilBZiAf
pbBfzOLfddx8ma39ql+Em7KmT/OZdF0SCUrwOgJ8DTavviOQgvVZQAhasR40jcZS+Wh1FBA/ldYH
Vb9cx9AbkXknnel/rgIBQQYXdhAsTRTqqr1FDsob6gTVhzMrRXbRZi5i4fvdidKDbNIF5+ANGXZ5
aiILRTDR+KPdWb3j+qB+vCtp3C99r6kycobN0r03ixnhn4WWzqbTqkRny9zCzLsHStyyYsSMifaM
rbYwkU6HoQEbRMOkBr3cb8Or3i6c7TdkxkrB1tVQyuIqRG64UpsxD67WF4KMk5hInwwKNUkMNi/h
4GZS0ioLXFFdJSE4VFN8t18saxA5IGq9gKRfehcq5t7UbMo3hx2FU1+TBD+vleDTloZhZ92XQ4Dl
Vx/miu3P6svw8s4UfXLOyn95LFFKpW0/V1cu0dPX1zd8jx1nRr68N6rbW8kgIg4gW1kdcWwOA8a5
YJxu65vrUNiIyi9Txf8YZPMe8meze+HZpczMD/M0MqdSKSsOXCAAeXUoqj7tdMiApqboN34MkxEx
SL7L0GnatMnpYyuvU44jn5+GKgpZrSwgx+ZjSeNXAJznKZUZi4WCrYj0vLZOrLW9cF0uZnzklhIe
8QCSnC1D+fC3aVzRpOG/BDj5fq2CfbFCzKZiYoU+mELFjfCaASGuKijBWGLFqm4cQvSRCykKnDSm
L62X79EABpLemIIuy1+NgvwIY6GsdE1wu0w4KgvXGo2LQ4qho/ExcsXPCbquDdR0lIef2Qj4EZJ3
CNj9gnbqsELFSx+6paJuxAk6T+7feJ6IOFfgw5EH4QzT6WAm38BtXzfU3IY0ICZnCsGK/15Fr3s8
PvwXNUtp8V31y2g7IFp0Z+0rfMrDSQ48qwrz/vTZpfrNgJCQSWvUSPOtEOBzDVw/j5nA3HGUPXL5
3jin23mm9MZqdmDxjOTEKfPMFpi2K2HBelGG6pXydkskItnr18d0aCNpQJXJMLNLnbGN6hD8MzeK
6hnaPxY5M97hKEgomNjDK4gqDoR61n0s86DCdqOfky97HLHSqfDrUVlTab0lDkqq73RwS66uVm39
khiTZoUVNygUkEqFz/XBQLmdXJo7Jate1uL2C89fjU0DMsN5tgz3S9/o1iNBL47SJeGIvIXdRtcm
TSo083i/Jl8C8lcoRIyNN15IyOXAvauRyLDvdCC1y6dAF/K69wx/Eho87jVCtlOPWoZAILqIIdvG
uMfoM3tZYs8O9IkgeWwX3M/BnBzRMZ7bsLllcbLzQC8o5bv+OHg2QC9/hFxG5s+TsLqRrI8pwF//
QFNVMvV+2iNgNRiGKSUhJx1GqQA4w/3wCjah8CkYXMddIIIH77Hcu8abT9dnlgqtse2FgYrJyEii
x1Xzh2d9LhXjsFKa1iIY8fBK26W44g1b350qH/gK9Rf4DF+ROGu8gAsr6mBY3rW2agdxIlOTujMB
Vs8/iHLCD2++j3DffGhkOzcJ3Lt0mdvLu9zpgq9Mmli6vYJ76Wgi2EAc5MvzmjBtOVJAgczq7ovC
Iz6KyyZimt1ME1BcpSURBtqi85akdYGl61v7ATSAv8EWRALVrLz1bJKN5Fz/4S+UxS3Lk73GIBxf
XtIHHgLA6fMfUMq3bnzbHoP3HYUrAr6h37R7O0TXSzMfJxrYG24d5N8g5R7QF9d4kjvRovXEQ4Jb
YqHd6Wi7u4vLjKEDel8J9bgM2pUhEWqYGiRIXVPhiIxUdqKNus/kCeXCBvIBKyGfs/betlRwAn25
2t40ZzSPmhNVbrciku7jBUa1qta5oU/1I0Ww+Q1iR3iXtz8km1HFCgWpRAPXxM5s5/nSweFHs66C
ER+ZJO9LyyxHmSoV3W1MKYQJsh/jvK5FtB+/0vZW4/5+w/H4grePJAVS9NvuRcoBlt9tIR7uBWn+
SLEBtRczCETV6q/xbghfsNIAFlf5QmWFdUnFPW8J+pmHPx1EfgvX9vrakKJh2A9xkv+wWq7Yxisb
bCMTiqZMjKt1cYVUxnmeT2LGUMeRHHFscJGxyj+MJQQ1idhU3Jksj6RGrIax099bWZ+YGe3Ke7mM
oBxWjx0dOEW+Wy4GQ0fCWF9VbSMnJrcX2vhF48IClPKB1u/o57ijfoemr7Q5xPbTaZfG2dmsuWwN
YcFuvtjQKJvo1EiVZA45KzDVqHxNAk7/4EAllU8Dj6zcksSJChkLNE7didQgww9mku8uI0LxqOU7
+4XLMzBAs9amnTNp8NO/o5pkEHf36w0YVEnTLXjvgIrnLVrcI45lP7LzkyLB+v3uadV7/PiwLjrd
dwmfbDQdzB3tstU2QNIe+Zqu+8/qeHnzOBBpI+H03DXTkCqjbfcqxm8xQlxGteMACTwFSc8OsYAG
Fbk1dNG2lpPSAefXYOZUcUaAHNBeXMDIOfFQ7Ol8Nv2W1/YFGirz4zGoProQ05dhX1xGpE1VO7kW
2rHtEmYoYP1x7ePd+XtSSicIpea88Ks5pb8xDaZ0tEuhVgy3QSeBrErsSj0+ydX08vLP/gdnQlN7
l2P1aCFX77T/4lrEipNI8AGCp3lnfvup7y8w3U3d4L0c4Nn0oRaU/VQSmCrf2nTtccqNcBiYUOXV
8SbO7Y/B3XFHVZGGIbIS/nMCrDLRuhfxvOkrnt1H9smYusGVP9xBgkeGJVih6PGxYbQhCqWCFXiC
ngD14y5DgY36B3kVd+TiU3icFl5NGhS2GzaqqyiqfJVbrz3jUU/VYD6IvAgmTW7mDjYheE8ICPxZ
TLEukQDhm6/kfuKopE2Fr7brjdksWNEdtiasPl6dy35XBH3SiEyslLqVWCayWi66y4jT1bWBPVnz
Y6D0kattBAtJeO7UF7l/y8s/YVjaSfWBKSNT/4Lh+Lv7eBUj/08tWnzIasLn+4cy2GaO7yfJaUBj
DyDljI35STDStPf2HxLjLN/vZ9jmPc5oYhpKbfwNaSPCJkc6P/q5kjYvaR1j+1YbbvIFDknwdqOk
srHTxIUv7HLNwQTJ6S2VsABPAImSfxpJu5QfRjQKlBeBlcjwu+DSwJN9vN9S//gAw0xn62SOjoXr
1tg7wxxY0J0AcaWnwcsq3e2MB6VDqN3umMmMN3O5O9sbhMj00YrEnOUK/JZQRDpb3eunIKw1hp1a
MKLdKPnMQAw5UZLEfQ0569CcKhbvEIKzrijLVBQFH5DxuhWXBhFdVcZZ3zYb0IllWGx6LxqG4/rd
JYa7VYRtPVkkyR5CjikcEshyMrlL8BowKlTXFysb9o3SmXbZ3XXmY1A6+yHQORa0bXkQncJ+IS+x
pRTJg3dW7fNr4J1zixIXmjln6USMQBhDm1PJRT5rskDHfSpkc27NMv5tf/IbEf8d6eWHsJ+fdfbj
lcI6voP1yOULSbDRLTGhtPLEGu8K5KS0V70AXNBHVn4p/e1rRQH6rP+FY76wx/nk50mpTWW31iNG
74ZWSCS9hXyElnPEzCDZ1CnhjD+0PGPTlDnsnwvLBAPifDBKOsfU+rysnGw+gHY26XJkFpTPhNfJ
E/baOjUkCEVerH9IFTI4gyHXNQkbvY89j2PqqbAdK/qEWn7xzqOucKbx3C+yICUXdIvnKgFT5TE2
cF2B90Dw4stUREPc/DAn+h5UGA/+ACb3GpMH2LznxS/thdXQRuKTJ7xnfGGlgjFdCRX257rhROb8
2RnBfK+a2FRHOVTVC6ZapQs7Z4H5mBb6lCy0hUMcWwqzsM/gj8brnDiq9NeqZSzmVpDhG78IuGij
rJMGLrkysiPzTbvAJZDEIyO72uxDCt1ONumzDpK0v2QYIQzIWxJY0R3ks4eyJuQjh6Ywv5J/2GRT
JGa05cYDAWVnSrZRY1fiHrkVKw5VDKPWeJ21Rpb6BdklNqwYWvuSu54zYCp1ImmuIwpHT86w0mQs
/0RaPZoZe124yiGQG/dULZqGlFiL8JODaTmfoWaDrNd9PILwFPvRsGxGydugH9N77Cca7mR+yorX
vEZe6DbwIlWfUV/m/p/bKZlJ0JXRdp0LxTQf9+jYlqzJ+cugVzLgDuwwmZhJC06RB82I78mwKXfj
eodlOFh4z/YPhIDZDvDTaOP3zKcNj5fvaVwlMn5ECECrlPUoWn/1rX6SKxbBTs3tXAD14iwQp3No
J2prH020gp82QUkn5C4wW2Cgkdwuf7hFWkybo/OfsmN5CcFQRth8UWjiQY0wyjJgbLQT57yAY1p/
WgsUW0YMzbCLGYwrhiFxybtkCaW3bZYWGgylWtdN45YGLMt1CiMWhuiDZOw6giLek0ikpj/4YBz1
0sJd4XdvZOxmUIrZTvQIUgnctRFi9XO8xzhzKnULKgh6+1mqOIcWWpxeKxjd2X4/ab/+LDhBzI+i
6itS6Gsn7L4xrYeEwPPX/OROb+nyIeNRYBVbTXSiXlEeqz72I3djVo39fePxJ+9i16hEEjgS+7mT
obMSb1BXH/ynnj58ilEzI/UKDgOiowYtzoSSKpB0Te0Z5KyqzdPBfyoeEy2MBwQAgJksndjn/QKX
Kd5sWob4ZshZDUezSA/A8JKCcNTbkmKwSJj4Th351KO7W84KOJjsna41TIizjB3OOD7BmIjQwTQw
Wz2I5oFZFk0/mZ/v5ltXa1VOk4G4MjM2UJAbpBentoZ1mn7ELN4Kao/troRl50sWqgx8nPyMzdKY
onHUv+rF/9zIweklsCI9wDmuns1Wgrd0SSKulh35bz09281rmvGwEvz2NrkzNvmuvNrGGAMZQFrG
rpfWzw+S/WysC61zoKbt/Nb8LwSThSiAXkCTHjukC9keXJNICANExSiHHZzKzZ50t+FlS43KT/Fe
wHAbhzJc6eXex8mzZ4VTOy/7yrW9pX4N4sFGAbKwq4BJVr7Kl3tnJx/9GCj+NpZ6fSWhuvqlffKb
CIml1Acv/tTHroCPnpHMG5KwO5LETYg576qDoF0iiEmo8++LpI1r2NxN03sfshpj9D7fbwaRhrpP
bvaAz4bTHOon0lo8kGTrVtVPHB4d7nAJEpqlH8JJk/3YcrSRH7TPrHUFkUQhZ/aMLTp5ro9i1SvC
iNkDwoRNey4iTmIfjH5Eaw6ctPkwtH1rCSIrt8QRxF0PpAZvrslVeabK5NLQ8LE3yu+04Bv/V+BA
/SwJ+Lh257Ok5dnslRUfM32+EyCLgCyWU0vGyzcA1lwb2MafE18epECR3rlgqScCQueFHM5PmrEE
yvoIJI4L30kDy4TOcmKmitpteHnIKP27PWEPRM4lOhDhhK4mRQZU6eavrqKB63bY4DHz8GDoQQam
YabMpYLu8mvfj8mxTeKamtGorLjLio810e2uWZ2Momj5d3CkuO5YwsZsaz8dMuqK9Ank8r5QMTyf
jqhPZtnM40F87PCtd44xtEHpuPoC9FkEakEqO0C0bdjaJ8/fpauqDJopftGFGrbyt1KI5JkLdMKS
+SXsIR6nQZZylQOWwQWw5YLEpgZFzmHAxxwlpYGpOxypqshcqCUdMMDk0sAMlrAEQMmGWAYOOnth
nrHun5PwdIkk5DqbCntoDMfP2DppRUj/+kkJjm+5eRKqmldR9aNr+FqzZlRl9RljLuDySTor90Vw
RAVboB0wz63ipLFcdmHtR1ywk/bVkFtSCghpqRc/IH774zrncTqXpQhBVx2dAVv1yUSO/9MD+T/F
tTUIIWhFqBYLbgPN3z6FFLKsRVmF3wy0eqZW1DI3MaSHAKyZW9XNSaNRMWLAn/Et2qhJ5mvUnQoR
EhwFqG08gQu4q9sZZ+GC8Swk8VJwG5fmDsdyKlftScA+DXaI+r09H+cIc+g0A+ZOYwXHnUhurgIS
Ivb+7gq7zi0a1hT87EmiGsy6uo6Kxt65VMtMeO0FE3TNYQ1Mp/cLiDjb342RlwxAkNlBXwqJHw/j
AUERasqC6d1lEVc1wbaBn02epmPHcJIRL10DedRgwJ3XI0Amum294yzyT+h+SbiU3kSMyTXyLMuK
hhPkUfsOHKnKh26+n4KrrNbfEcQRggAbsb58joqIJoksKp8TXoPXl/RrbY7CLCI3hp0voJCMDxAj
pMcK3Z3+ABauX7ZPLjIxzvF6ebxjTqZOVg1RVkCnbGPDjdGbQsnYncUUoyPSHPANnzgvPaPJo8Zl
Sb2nz6FfFnOy4BOu7BJY2Ix+Cwo1UdwrwABxa4iFuFHUWXiznUkzHGDU4pcgEi7uWnX2zwhL1GUl
dvREcXjaSeNllg5TjIR6z6jpOSeZRUK/QR+x8Mx9f21rXLYByQQWJKFzMQDwImxFKCGzsTLSkRFE
9FDGoKxFKOI75cqnhe9fQMftS8ng4tBcmcsPwdB7wQ/7u+1sv+5c+DjziuMm3VEQym+sVJE4aNAy
k3zbSisDlazqZhk+0Ie8+mAmPTN4DK/CEjpQKD97PvlqSOYNFHRpvrsl9bQFdzng0mvG/mZCde/n
vYjrDALgKBQeu7Lj9CD6vCasce9/TILm9ltitu+x1O/EdftRHr/090PYjR4ZN1fo8zdJQuXqoII8
8i0Vlki6nwKoB+4H8OJnYQn+dtBOfLREgpmefHmR/El4ELTfRCVUgdw84XKzmjxTqsVDqRgOZ3Ck
aFW+8cAzT3Je5TbCZ7ZI0wPWWDntYcyFASUZYaPhZ0zX6Yy5z3/DUsAkOSWhec7G9lYZ+XMOjJgw
UCydNdAtc8JEQyiXXTsA5t2gi7u2LPuV6eQaU1KXfNA0X4qojWyzqTMmUebNdmGqi5VDdwJXaaYj
hJvkKapgaHZmTw5KYqbEHPfMC5dWWu8YZVgHG62cKTbQw8SqxATW2A7VE8E2rdc81cn+tcRivf2O
PFViCCllSm+jAWkqdWnX+B1AovC2RgMu8M9mVwxi095hdLvI4/t13AixefTtCcTZOisQBnhzTu+C
yapNA2P4pBblUUMkTdqNE84rSogMpY4vTDqLcVYUsxQoWvgebVJ3Xno2UorTUbZtUdqmm1wS2VtF
BzNczyPrMEAeqUwgHW71qPP2+51RST6ElCfQ2ifTg43aDmVXHIHysgBYqtnzHXgALVPqbWdbtD5M
Xmvd+c/tiDm66r4un+QmudQ2wXr8EREt/ZNuOX3+aJnLcyOK7KKcbbbpVkRkUGOWW3LcpBsGmq7D
sSBY2mdHiCnangEZssaMvdpYkYybK+t7Kfx2JAPGxuSOGtX+nLE7S78r9447eCPliE2mwAgQLknW
5kiIZVpUrMkEwTNuPO8Bt0OQ7EVMaIDipVgx7mHD+xC0PyqjSufNy1/xiTlKQcVRAHeYXC0JoMho
9MXdxT4m12Iowca0JbrCuunLLHFpUGRdKc4sMWlDXFq1JX9LxfDzn93ANahAtTG+pSqobbtCCqcx
Af1dU5rWiyEjyU7pNirSbS4ULH34wkWr3OHXQzJ+rf/ZHN8aVvPXqdE17ZvJVYtUtBV8Z+Nhr7o1
QAJB0ie8IZyGQFYjVNZMDkq2zBYf+d/jILdnBUeR2nm8onWCsIj6IKO1MBANOH1pnLWGxq9oA5Fx
dIdtNYSyZFxxTqltj6bSoBy83mVHjRyBzveazdDToe+3ZLhe9DZwlwEmIbTFxUgKP8+o8w5EBCFT
QxnnPvSSpxPeuQZ9Gz7ttMEJjasMD0W194TnQGBL0eZ7Kz4WVYs6QciMUpAf0sdDkFKXvfbFgn4U
L7A2skqYG6B2oe83tI2EBGVFfSAeGrb1IYo6zQPMSgZoYi7Ak2BmSRoh55Hp6VB6cbnOa8Uw2frw
XwDraPeY618LDgNiB0ncVn8mYMY4+PBxFOChDwuo/lqY+hjNqSiLjWWMzgd4V9lsukvAX/qNP/ND
FlgUz1ZmfD6PXF5WEl9NRGpRDA47BRXVST6EkM2wQUMxaF9R4VcSNRZwW/VRsAR8EQVhs2LwO7Cw
3ipedwdbPB90hh49cAn6ZKBdIHYKhycmGhKP/WULQwPhjvTxgvru1C7IjkqtlRfbMZl7fWmrnCYx
2fozYvRnUmNbs/5CVD2SNLkLrMbwPsIZjk8oIOCCHIMneAZDkb9lZh/nHGC21JYh2mYEuB5Rm7gN
DF4ZLMGG3sx7KLbXfE4270VqcJHNMC2rHEvXvMnAQWw08LEZOZ/xoc+6MS4Ku4oaS48Z2EJ8JzDz
WpyYCHKMgNxHhB2HfP3n75FX5VtDySJsKb8AeNdeJwlCA1hTA70qcjr9XwBAEdsZx3lsL4jgVanX
dEo9MutcUxmdem0gD4fIqMtnLRqPKsdLL3pMhhTZPitX54Ei+b/LtBZgYsDmEJLEGXLoncV3E/2D
hPjwC8l8md0Xk9BsBAOOEJw+JsObQf0MWPm2+ICgkSuyXAu6Qrh2dF9oazDFQhClMSuyPqC9YQsT
9DIaOw7sn5LPiTaaw4skLe8raLmbMiiyQcTgP7L/XrLczhvOG8xADRIivWtoWN0AGnWSzsACOXCG
ZsUo4VIo0p6H/D9dcpnECS+ctwwD4X09C2VwDLEoX9fLnAHHFOcKP/bl0z6SXd5f5xiOIwpxja5C
pqDCV3Y6sH2v2suD8egkddjCe+7QqOBaigEInJZeb8Dz8ravAPmBqpBfi1UTcLTnhkGf46zlnqfg
aHXEbisME1yDwIxm/x0+fGC1vrDMvescRbzkWQIuQyW9A5+Ug2ifekmZC8A6RM/agxKmhkCVHvPX
DWnW7stB7bR2b0IviAnOWJUsHGRVWbqevmaVLJhGiS/FxCsRcModEyrQ6nWn0SEeeSi2dUuBf4Wu
xRjA3p/tSPGyazYXM5w9sUP6FYiuRR/zoCd0hN58znnS8xHCJzZjHXFguRMgnI+Wbt5yh0XH12uF
qzm8Z5IQUhuZk9HhrQDb8oCqtyO3009rcDjPX2J9V71Ki1EMnOOPoEgx904aixA/JhqVAUsu8PNj
Qed1NHAsCIvS7IcUXFPfy3uGnISa97ch0j923pnuJcU3vBc=
`protect end_protected
