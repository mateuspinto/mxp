XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Vv�5�V8�=��0��#�f�fu�:�+x dO����Q����(��(�N�ꗥF�DOG���9�J
�����ᾡM�0E�>�#J��'}w�oJ�� �����/E���gN���jPnP��I�3>��W��jIɗ^@�0�")$�Z��C�8�R���E���D��6+�1�X�-�w��L�ޫ,CX��y����L�ݠ�_D�Qe��G�c�����i�<�>W����3/<?+u��/�a_;��3G�l��p�@���	��\9wt}�d�f[��oH"~�F�*���r�=H(e2KgR�+��N�"���~x��@�z3�9����a@�L�P֖�fd,�S�W�0�Wk��7���yC7��eds�b��l�X�`�4���9b�D�dg�}@��#�}WH�EV ,�k��+�VM����a�X��;2�b�exX٣K�CP�a���}U-TK��L [<�)v�t�(F�����VQނ4D�-�V��]�;����;��Ûq�ܝ����p`��	�[P=~c�%m� �ԃ�
�ԯ�-����v]$���j���L�=D̶ed�H��8'9�8Oyn�x����.�B�UW�	3�w�����P`m�	3��h��"�#���S��y�R��C�?����ˣ�&�ש��ozOͼ�Օ��!�6��M{s�o*��,���L�ڡ1�w)k6���f3�ZJ�����Ԁ�u߶�Kt���t�!2Pu�'�m�N�j�>��+�$#?XlxVHYEB     400     180��~9�2�
>pv7=G?���!6��<��<y��چ�
�e��7��q���`x^�*��IHx���;Y6�YE��a#��E0%}��rq� JQ�&EH�C�]kv�P�ԉL � �t=��% �
�
�[���e�y˃�n�;�\e�:P���u~�iJV���e?��7�JV����x����q�̀բ<E���-wH���[�eX��8��9�̧�y��3��D@ e�±s�B�z��܊�s ��k�1ݙ+�0���{U��a��&�g¯�<_��k��j`�@3��|�:�rRivd��y_Mv�o�u��kC��P�91�K�#{�b���S_���K���x7����8z��6SH���kңvح[x�2j_X����XlxVHYEB     400     160e��9ɪ}��$^�B���r��/����δ��^�Vcr���I�#E�-�Э)�������B9`��;��/.j�_#�ʣ�CH��wLll��B�|�c)���t)x.�Ӳ��G��#9,�x�����&�J�9RL�I�$�d�V�u���S�f/�
Wu�ss�REnƠPQkN�w� ��J��4�C[T]��;&��R'�Sh��1��zo�+�r^am�%�H;����*6ԁ�9��u����܈P��qX� [�	
Fu^v$�Ll\ۉ62��2��# g}�ނ�}!¥R>o��XX_�)�b�ZKHָ�{��a�b��igT�/�7q	�ۿW�����Ԑ.bXlxVHYEB     400      a0o�ͷ���N�Pw�o	V��p���Z@�o���!��2�޼�.~��l��� ��*��9Tհ�L��ӧ�6JTh㧷����Q��g3@���t�1��;����e��"��]~���8&~Qc:lkw��7�=�2����J�I���FXlxVHYEB     400     1209'��N>Y�>U�{��w�oG.�oK
�6�l��ؼ���S����vK�5���_��? ����+��_�:d�����H�>�H�0ˣA������x#�:�6��ա�\���%`�:��-���ZL��M��-�c���!JF���	t��ք{n�pS��5&d5:���e�ޢQ���c���[i��_�1V�M���{�;1�ͿI�\���t��t��^$���1/E�K�06�Ζ�4~���eBz�Ya��8���W�K�>l�B�(@]��7K�`XlxVHYEB     400     110�&{H�6�Iؓ7��ǚ�v�T97l A������*M&��6����4KY�v�c8�Vov$͑X�ϴf�,ME-AC������m���X�
�.�K�����H!|�p����C�|$z2��Q���>3��]��>�f�%�!���1B�W�\�^3D��P�y7)��ne+�	 ��[ƒe���_���[i�/ I?ߌ!֊��=��@��#;�@���dC��0���K��2�_��]��O��d�I\�Ņ���[���9
�� ?�L�EXlxVHYEB     400     130��M���T�l]�H��m�����nD�����"d+=�1�|����V�FqJ�_L���ga�
����^sф����}%I~����+��<Lg��x���:��I4}K�g�=�(
����ղ�Yw9rc�-?�R۫�2���?H
�(
��:�g�k�K�3���0P�z�9 V��R+�Mw�#��iZ�c�j`Ӏ(׿.wԌ�C��&��B�CW��X����^"���ah���IR�m��I�_���g���2���6iy��M���4�#�`��q8�
�M?���l)�.��V2XlxVHYEB     400     130뿊��*\x��7�+�X�bZ�7R!��1�ꢴ�����ӫ20�3�T�)�67���42�-Kh.�N������ϤM��bj 3�	p���pڜS?[+��r��+Hh��|]U��zs^��c�P^xa��N��_d����8Ă�ȁ��1�Q	���H�O,A��$ȗ=@���/}�JE���#ʴ-�����d�qY�p7�U#�s����|�?��Q���"��'���H^I��.�D��7e�[�r��(����2��O�0�E<���8{5#������� �팻���w�
�TLXlxVHYEB     400     120��'�a����ߵ���3��u��vd
]~���ǶTϢ��X��,簃�˚M�3H����o��8n����그su%��f�����
����=��˭)�H4��J-�$"<)����JH���e<\��9�b_���:,��ԯ�c5�[���Vf|�Ǔ(ѳ	�+�>Ky0cP�p`��ڔ,�j�5uY�� ��lA��_���R�>�&]���J���K7�Q�\���mh�٫U�T)��_5lw�{N7�'ZN���>��JUW]ir�}����XlxVHYEB     3a6     180���2d����V��YF�"kl���������4��ϛ+;�b��K��}�a�6��P�C$2��8U2R^'9`{(ՙՄi��l��7%0=�W�\W����s��#���T�����x�v��[ �߇6ֽ��_PR��g����DI�Pf@��}(�ħqEj�/������nb�ah�r�s�`d�[�[�Yp�N3.EIKrB��B��j��DdF�����u���hH�nd����ٶ���C���Mi���a��<��%�0f�+��"��_������/ �`U�R���Oe������a�6��^p��(W��z�?��x�&Q�Z> ��\,�Ş;�Ó�!b��2:��2�
�}��ز&9]��e����E��G8'_S��