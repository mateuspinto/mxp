`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
HwNHDl6naOxlRGdZtZlV3nlrRk49w21MqAGFR696TtmAUaAtjm+QvKMpYQg36V8/s7yVsqDzJRzy
wkO63PH3V58UrgsL+PjTBCxBV1CXbTJHJRgksLAxyw1xnz2ySZyl8N6PvSKmoxvBzs6Yhq21GsNs
EYFOGxiluSQ2vm4K8bu76E2K2mrIRwFTmaUa30qEQZ2dRF4scHBXZS5v2pTOJH0z1zNS3ZAj4gVb
CffHP4lobX0OxNPgSGQSnUbv/LinnT6taXKt9Guh6+Yc1P3luwnmHD1rM95RlDsuwZjZrTAnM0j0
HPzYfEYyVDBwM+hbPhL3VMAJApuQ07iqtCce3w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="kK82Ibcnv5xV58idC6y6xj3MU70nGrVkafMLoW+tyTU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6528)
`protect data_block
Xo8FRvaK7HdZJntGQT+Ne7ewYTp7tcrjujGuAYEI0j90J4k7HUj0X6eEu/2J2IYi3Pkw02xjaTez
2GuzfuHFZnlZkM3jU2Rto5FqpGuVNqkCqPCDEFuc3Vy775Vop2K/2YEVsf+GVKtxq81YbVRG4/vx
QjxmxRx9ROd2ZjT4Fn+60sGvX4RJBS8YocVLyL6hcg2CLVzFBo9zO138b0lADnNWIHBkTIK43gy9
rN8KBEgqKq4ixLDStLA0kB/5j5KGXT+NVvEGS75HrVn2ux1/Vt9V3PKcqztUJx5FFquaDb8p9BBs
LX8Srrb5FgD3XdUNTJILEl5LRywauTqETQw3EQ9D2qLKnCAwWsg+jTFv7Il8z2AH5Yps9febEaun
ER8/ef3WfT/HtadNTKi/tB9LA4wLosUhA57Hb8zb2hAlfODsP02J6T1cpZChG/okxhLKcEFn4kkZ
uvUNCDUKs6R1lVlhUXxqY/G+IDDHNnbDTpCGw6YaAonbWzJ63Kcy5ZVxcq8B8szjcOQ30pmTqN6W
MMQt1sRnq75OUcABIM0aOAaSbezJE2yqKrkBMdtVgATyZRwtFYk86yEef6KYK2lPfSUijTX9zdr4
Y4Gi7MTAoYGNed3CHjVhDrhkpBvCbrw/ILHe5ePLjEM+mGgAOiMsohcQdB/Sj64A394rgNkVP2Gb
Y3LeKULvJtITFnpack7YzMV5EEXb+X9XqpJ2xFdheMHR0yEC0N2mjMRkX8a6dB/G8ew7FOz2drNk
PISdyxP9gdIxwpFzKzPHPFeoc57ZjA2MPNOXBoqVw5fk+vAQJvmBaxg8mlY+WLjSPFQVTXXt0HfN
4+FmGN/Xd+vjsr5E2KLzVCEt7CLzZoL9JU+cAk5DX/bTgop0F/0GuEYZu3aspXTtkFH1JKEcyvW6
Y9jscKKUl/fduW+dyN7L0yvC+8sIurDP9CB8FDhuaKneKrFY8eiVd3BFtRyzeWiLL2lpFpaHKTpK
/nmA00JFoIRR0nWXYyw9XaqaKxaod9RL3i3DFTFiqu7uetzqh98W/DrZxyAHrYJopsfo5W8zomM5
KLiYl7DUW9sTnuxMMxylQ6cYNo/9PpKkgMyP6Vx35arZ4evOeRdr+w9lXoDMaAye55NDp7TDwvqk
cUqJz8xfS6HOXpCDmcZibeufsif64OJfWB2/cSJfQzmJOtXR2nAXB01YSgNPvxiYNhVIdqXUNgRr
NWISDbX2da7huEEJeXVf07a8ojs1gg/Y/ChaU/lhbofLVJtgyZZpB7NkNNG2vrRArDR1ZgGX74Th
cf3p5NvuLkTT3Ioqmgo0wvsw8yuk8L35LWn8EtDDck6vEg4iFdIfX8ql4P7gRZGhRQKzY3jp2gE8
7F/4Xpu0WEOXpgEh11/TYH77icQEInIVbQ6j7BlaNYQC8+ba3L7FAq2Iq2634idU5WGChGvadb63
wT+IqwKmQ4S+eiiHxBQzuuy/2D3AFiReKqOeRrLXr11JJanQqwLos49Cmr9S3Qwstt7QA68BfGRt
kUbySVd504m+kL0nO0EIcvW8OzNrfbbDOf/pUr9JPTauOdoOI4sQjUHHFbS4gkv0wWvlfc24SC2O
34oQoRIpAiMaMAxmrFuaV1lCautCCf+PxMPf5eZe1oCN+TMb3EIegcJP4zYdxtS7N8K3uR3ysl0/
mU9QH7ENcQof51/IC1cQ4PDHWBE90XGWB8uuGcpyhzPNM++mayF4gh4mFY5+l5lK99PkW1A3b4cU
fyTdlzPSGqmxe220raSkwVvZ7oiHNk1i40wfyhsYJogpa7TDj+XQQQ/2ZKq/SafG3GYyjEzrrxuY
gizaTW8uezmCorE9+3uBvS1dU+gLTWa40Fh02iRcXeitAP907TXDMY3mWWn0nRw+iSvvR9hg5+wz
I3gqUjVP5CavqJiY6mGeQhSs9BvEsFIxx1JARqI/OS3qZKjWGBHaFOr7xWwqyGkowpG+g5afZ+kb
NQKIx1zFRDcCzg6lyj0Ab7y7UXQ+rLAvKC+aCsWk2j5aVIOY9FE5OxPw93gRGY6LTQATLYm6tdT3
W/HKLQC9zGj1S3UdvsjAsJ875r7lfP2fp/YE/PNZOd+Dk0CFSXBALsCKW8JcWOTZ9t+3pWHljtM1
dmUsJQ/7WQ7uNMdAzROutRHmrh3uEM5dch57yg49khp8N6LgdZNN7Arylr2ymC7zWdLpWMmfbeNM
0+WRCpDTXeHuYZ9llOMMuwtZ2/TljikJeXDplcQ9TGgGWteCZPnuQ9Y0TuTgS2lCIq42BHIryr4m
XtCtvx5/y0Qx00LAnpQZE+7aBlaHW0vok2f6ykf/em2wmsYBMVWkaoWYxmZ+ormUfHos+A3n/MNK
TjK7sk36QgqMIAUUGl5GdslnoqFg94x+u5O0F22pLBDtFV2TO4mxEia8zd9aOwDZXxXe9KcXhXZ2
GEkyp1qTjrs7WTidMaYA/GKkIdN4GqgzaVGlJfOx3vPGPgJiUDI3IN/OscQnMD/LeSNqe7Ut9EOT
TSvkEzY1Tv799NrEVf2MhymdjOMYIO+ZBl1sfNKnV+63CvK8eqQ98qDmEEyHvGqLfQTpVCd9/FE3
P5k776oYxAERjHvLbr3Q5+iXunj4ZA4Q9fgt9yNUM4GKQKV0ooJz5rtt6eh0fI7MJO0xEpWTNCEH
7aAXrcROAY/AEp4xGElpTHEmAbhzuFaQ/peVyiEkjpBFa6kbB3zC3jk3yBbd/fwaHl7Hcs43o+uM
YZwSiXvY9kNnZFrNkdrQvGmXElIsE0ngK6/5zm3Tp3MUXLvYE83lyhudLL3R/Q8Qq7cEleqpHy1+
BcPmqj9Oy9MGUEjiwkCXkzy+BbPt4df1IAkZgzFYS7MgHHYQV7y/QMEWlJuZbwNfmnoCa+dbRbuK
eBmIk8FD9urpc87zXeniVh7cR/vm4hO7GsqguOSFC8WrKz2tjc5NwIFv676qqRlfx2xnHLlKwSBu
IJmh0FLg+wLZVfCS7Oeu7E201qxq+olICgOSkSEFd8bwzyDronL3b5ekN8y+2bG8/GVswQfGt31w
K0CESM7u2shbBKGMWhegzJaA1j8hy7JrZ9KV7L+TjO79Ci1Uxm7Cpt12ZThPQ7DjLCUr0vsQSrb8
70qcBXpZKl4Y5FAmOwGFuS16bnRrxeKemtV1YVvnw8cQm+nq71HlnR5eXSd+ZnR6is+mtFto1rst
x1IDkATgVGGtha2EXVK9OgdDWzEM5bxA84Zw2qTxwjqZAT4pcqTjLOi/HEM01Z6ysSBf+ghUVtio
BvOq/sFJHcaO9ELdWFw1ZuunyQV/9C0tN586TnPL6HM+fOQxMX9W+Tid4o4NWnTmsCw6FO3pXWyP
KRncDaPvE6w8aFUZJuP+jTFOcf0qg/n10Sj72ZcRCyvY4p1/BDYmNc4teWhp8ARoZ5Vbf7EYQzEm
IbS9NPTZdrZ8HUjFJbXi77c+rhNG8a4tr2UWV5/hlPCTyFESD3psvXTz0gYVOx1w6YlAmV6syTjF
n+tpmrRhzoWYtKzNMWkOAlxnLg+vxNhDcXyar+Y3yd2ouMs9Y0iL1gIY3Nn8H++Li3uITlRbRvS7
siv9SdKGdodqQVsz+neHafzeKMqvMAA/2A7AIq7kxgRHLz+PG4TPQgGBM0FQU0Fon/jOqPwShCx0
K9xBKd4ym9BPQ8ftiCcCs4U0cC6WyZGmrZpnkO+cMDGrtfoNvjD58f0PBmyVvo3wc3PsPtHvkGhe
Jztc02pvDbqIUDhyLfjF/Z3lsHd9HU+LUmQmtPN+QQpgHQYA0iST2SN1YchJRVxsZTJKXcWZoDjN
DOJrJcjYrPRE1V1CQDPA0RTNu0NbqPuEZgj6C7PaiWMtiXYYWS0E9arylSAG/rkjbGBHbqQG1w76
MB7MBvUo1W9S1U+0LJFD4U8nBsjrlOBlBa428R+Srz+FElLfUGRp8MOD4YYye5dBSJ08pEDiXVnm
ZIuGUidujl8KTnPWFEHUgjof5TW2aFRywGipaxFNe/dq6hg03lfoaX2jpHVqXnJ5TN981ejJnv9o
dxMbSgW2HnbZ+dl7EeCrE7DU4n6+pO87yqUafWWKjJx5pVPW66LxRMmAnejlYAnOqzBB3lG2vGlj
+wsk0z9fH7QTakrseKDqvnAX3ZemGfLGtkhE8xRHejj5CiAP6cRXmJb+xXMav0l5U4n710IkuPoG
vf638oTJpdEjUNaDy206LBTIOs13UgDFz+LM+6nPD1E/upMsSzhjhAD3A9uprH/xzGM4aG9Uj7iv
ZG5A44kfXhRdR16GDj41GL3nijJEr8NCmnzDWhELV11uWDR2HmquGW16hUbS6EZWkTATSyBb+Yed
8Wg/zob3LkM21hQyiCxNKGTiyngSuobyz4rAYA0WmU/PR6/u7HPccbfTrT7SkJeeI1+dJLCwszBX
9XDiwRVwuAsmtecsdbaBcYPiOUbKAdskNSAFmcBd3ZSpwsTiVRwgw9gzcXX92IFXtbIKbfmWnjG4
ev0qstvozRTffmpo1irL2EIw97PO5ayQISlJ+P+T3iRQQFHZs29Oro7DJE05FP6AkOPEzw8HvU36
DOf3yA8d0pM8xDHCRRat1hToWAoEAcX1vQEUkcHvUxXXuDfRfOsKXRstG0RtnC4i7rCOiC6FET7c
A3rdYJUtSuyxiao7fFq5e0YoOdK2FFlkpfAeJOohWMXdFdnIhz627pUe2s8OPY5NV/1KMm9AYcUt
5dhJitOKVLm39yiswV/AEahYPEkW9QLBGuU78uEek2lnnuR8uTXz2cH3Go0DFLIDuU0Sq5p1amP5
VgQ10g/mhTIxPPZqzsFyihnWT8lfOhA3XkO2wH0UwaCTZcB1oq8XQPb21mefxxY1u29lANwEbax1
7xpPVY9dPjAA87uKskjX8u9a16qAxh6omLJL78apq8HogyZm5oHwYmG9JnOpuzI9kxxN5Om2qxuA
SNuBnjXXXuzAlPzzhW8Sjmx7tv3CbiqtglAcUVIbRGVVWpppWOesnLxHxX/oj/qUHzBPLWsG6N/Z
uKML/AhGPRECRrhdmOVpD6kdQgHAR6ptqOKz+mV6Pff6EwLZWYO3l4UbO9u+s3R3/8ZtpEwa+GH7
dy2NKXGYAGF3NbOfZT290vEYtno4jGH5m1LvigHpNeTh4b2Qovsv2ELmV6FWtAvX8KDvGFViMZpy
ukm9zsWllZrdj0zryEJgvLDIkTbuNV2Sb7tkTHNVDNAaPM7GgCcT74TtoQqIvGXEBn6yaNdqL9KT
DoZZomvMwyzABEEU9Rh1vJ/7cGWEIjA9ockJpjubG9FL0yLhMd0ns9aTlQYEPr3+MOuPgmrfXEsi
80XXTs6AnFbpwWjPtJ08AGbedMNSMsigH91uXIy4qzDsCHJgDjWLKtzZX8uTMKY1KoVWTujTkkif
Z4oEJweHWTLu6CEvBsbwgBq2G7Wt/g3OPJa1mRCf+kTmPrnfTtmXzRS01tV1tOghAy0R9eJYwCJB
D2WFXk5JQ7R3JFSnX+jFclTESJPaEqFJclo9xojCMX2IRuDh7Q095/bPxcjQBs3qhzRD68AmA4x2
QD9EIrl2OTS15dum/MejcxTsOXGBuvb4whrdIFtJ+d6/dc4eJiq4bmZnJexWuQeUDSVlCQeGGwEk
yBli29/dV4s7pXKWAWhk/Nf2zI+x3tY/GiuG6KgrhR9hw0d1iaJdtf8tPsAbC0xn45aTXM1IScgN
KHIK8rvAa4SESdv25e+iFyMY1O0IGxhdCfKXYgNnRUjC8RFZrml6/ukFyRpSgiozOPOPrtFJNqsx
1RsJ0P/goq5uhQkh8klzhhN5OkBcRKJLaFQhld5dhEyZ37rxWmzJ5qeYxsAPo4DxwhItdXTyczqw
MFlsFktji+rEQeS29VKz7qFdp86hsIQ5LTpbrpfCNa+eA1D+kvURd3DJXDkIXe65gLrM1dAkYj7O
x46fNA3xrY75cjW3VSpIpsnP07ilGvNt1hI1OrB8osyJDuhK+WC7+4NREDVmbCmlFJjnVqD8312c
F6QcLlBxkSALTwGLOhp3pRjh6Knyjyu4COuoYcehGmmovlz+385HgpF8YuEdl4FECZQeCB+I2h64
NgCui9GqJbV8pv3buyBdtr9HjbyKGxAAO/IOJe+EsYYvlySPr0CFQ67jF9vmhaj5TCXZP6d/+ywG
IPzum/E+hyJGpt3JfWwVvW+7POkb1V56LnGr5SlyPf/eeprT70A90/nYCGkQaetqHbcDQBiN0vOU
BIOhNn3Qgguh3NgaMZNLnguh8ZMdDnVsHtXL5Ou4ipspH6aLG/fegMHkMqvLcotrz4dmmxrHkYyq
Q8wjS+aL1UPPbBpJ9VEjEVTC+FLnCcQ+GEPm/ZzNF/LckEWYJ448eAW6d2gumklqNoPykSBnV2ua
LkeJgikcyg6DDDmjlJLdxTrPBYOvvuTYkxKKskmslBXIGdx5tcpVV4KfgVFMK8fIXp5gwP6dA9C3
kiOlfzzQv3nVRH3o1s74rQbKnaZ/1ygY+6OxrbtH7a+MciBE2GYCfjdQV/lci4/wTZuujrtskVQs
G+lzP/q6BcZFflLLI3s6nSApCADGjYpG8y9zSaGqnBYpgRwFMMIHBlhx7WpsLR03sa6F0huULq1a
CiJy82uVUEdTA1hZA9aGod4fF7ql9kEzcqrSuv6daxvZJLh6c3wuz0/OTFB/I7r2zqr4SgENqMZf
wrjLw/o17WbMA+jeiHC6i6jZ9MBuw35MWRferVRByjpHmpvmjxiwD1+726E2Q6fMkfWoRtyE8L8S
5bLhmRFV/T3N3BEeIovwBLjCQQionEQHS8gArcf/DDayOjJfZdajnI4o+Jmgmuu52mnZgSwwNzQL
Y8AA660fmnZCu6DnbtTN+BTk+UcqyDAoSixdd7u1o7/7lhgwjLYx2VzCqBsptjjOe5z3P3iQXKhh
kJxe358mw19Js73XNkH6yxFlg6K8qV7I0aXcG0aZ/4w6TlB4PuqPFotgicHycACZNdn6cmL5G5AI
DKguRiMls2aIFXzXz1YEjLmYDq7rtvFc7/BA7E+S5w56eqpRpcMqGv7YVPbwrNoIv/F09bkOrYm1
1kerAQFlz4/Tsitsv8XbNH2XiPD7vqrY9WN9K/Qgd5qHFY5TQc8xNl04hwD2du996rmdk5uxcbbH
+9b4fVWDnIO6n8heJ7ENJFRJC1RVk07mqeqz7H4/rk4rAhHeByAotTWIdiWBtesIx2tKi4lvjzQx
vTfKEW3RKTTTTz9ojSpV/IDX9hMWSU41Bzsq04dZJMyFsyjkZG3demLwKj5txG80Fwk5iozDN0lU
QhE031QUQIghe4byNGsVmdpmDlQh2B4wNymrEVBMzgBHuoUnuCphwuOIHLjXQfZjP7un1PfpAr7P
sDNfj3NdeFhbaGbSsSyw7ZR7uyXhJX5lzTPvGQ+0ChpLd8iHFeTN2t0uxSpUv1XBRmwhgncj9shr
lTaZJfEJvm0+3k+60kPNmSG6we5kUZaKvTAZsJM6nl4rlJcJdHHAJvt+dAfdw7eDWdaa52iIWu/R
v7diZp+szUkpFwwpQraF9x/omc5bU7vIyoeavgOzglzWsNSFZlQ31zCvxaGEUQ5aIl/A2IrmTv/d
fnDdqyiCL5Iyho6wpzAKOZPTakZyfG63P4MvC7olZikSiBZQvz+21/r+GVSgAaEn9BnpJubyhT3A
L607DixGyeRL5V3VNx3ldr06dGhVit1Ol9XJx/8m+cxxT45h0aLrbRY+RMkDeNX+TIOvlflJIetG
i9oTPEDlr5ZJ4MAU3JSka6CQXFmkhW7vZC0PqERxYJrwqrgv1NoodNMXBbhq9WwvwOwsVJDoxwAE
8NfylZ3jK4ep3m9hvsOThQsYI7l9b+WWjd+rBcdvodsLejbDBjT3iTInLIWSr9Hxg3xwztRXAruI
dz3LTuNykes5HfmVS2QxuwKL6srJsuC9AQbbi19lAv9Li2G2Z8GM/TBDH3V0JHLHbfE4Y2dplW5G
+m1x5kaYuSgQtNJWVf5TUn8wjhuGAphlTrhdVBjkRCxK8uipbxyUtadmX+vdV5F21RYO40UyLcHK
EfhuzPE0OZzSwP+4AisVTlwgyUYc8w6YKVRILds55/9ot+8o0oEAOEOFbosNQgJWZKSRQkWVGe/v
FQwvZWNkQ6bflQ88FnYKZB1mftcbligki7gONa2fB7C8ki3lggT4rvNwuuiWVr7YCs8qcLuOF2q9
nd7sHfLo8xxF+L6VJuqdosY4kZ5y/zeLYBThZn+QL8gEY2H2oGWoFCP2RhiaTOBWhO/b+VXCJe+X
7FwaH0aEQxCYylGMFItW5j/jsGEzjGvVoDoxJ9Q8o1MfMK9tZV0fKfgKZmg0Kp/J3hpGkXRurdNi
UTRLaE2XE0SPF6+Sa7tgwpEk2pWWeVhCxRW34ebDFyy9Z1TfDjGA2AMWWeQbI3aJy9zrCSD24U52
agH78QNUknqL/wnV02ZvWUOYu6WnTWQXBr6Pd83nQPyfnqDtp3OVWxMqv+XNimEoi3Xv4NlNMlF/
XN/wcUoTO+p36VFhjpS+7UY6BWZJbkr+N6efpZ/huKunRKqc6qF1Za3GtAEBS1S9E1/ECEbk9RNR
zwRx4Nvq3US8ZDbOIEmgrB214KGdMjU6YS8w0P/LhtU4vmYU22YUdotKJicZf9T22W3tGsVpL/Tk
Ur54ly2k5kxeWFxRsWR66TrLXfesunulUnlnzhcD
`protect end_protected
