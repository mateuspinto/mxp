XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��:D�rJ*�U"5eZ+K'`:;�I�R�f�,;�s�μ�"�7��f�ƛ��s[�!��e�TK��w�-۱�\��C�Q,�׫.�v2/��.����݄ރ�v���׷�ZdC�(�I�0#�kȇ��jN����Q�Nz��)�w�WX���mR<�:3��
zu����Ư)�~�̞*�J%I)�T���d�i6&C�t�8!��Q�3�`��ÏQԧ9����A������Q���?a2�@��n^��Z�n�@[m������qU�s���9�+��9��
��ǎ)=��w��G+R�d yE9߮IRbUJ��:�=QS�\�%"RC�tװ�!� �@e�� �36�f0���96|g V�p'���a�x��a�x[�He���0��TC�E�*��ƻ��&ǬUcT�F\Q��G;�:=�&�~q/d?_�/�vټ�BE�ʏ���*/=Zg���b؁�����*p��!���7E�M�S�D���/otr�B?*�蟺BcE:B\s��2�=l�c��?ϋZ���U)���9ӫ�X?��<g
��ˢ#8a��'�[<{�a�o�ȕK�hhx2p��\��bI�-lap��w�gIܴ��a��0�Atf4�����m阫�3�UGj�n	������|��ޖ���0}ŭ�[d�#��7�F�缨"��*���'���?49&K�(����)>.�Ы� ���o����+��pk��f�]=��[A����v��>�&a����T��-�'(:Ɣ���9O��"ɿ`�$�!6��Z��\��)��]
zף���1(XlxVHYEB     400     190I�{�·�KT|	
����r����vAu�ؽ���!z�-Xm�LH���>��2�S�^ p���f��&�9W�+<��ǚa���9s�&��4;� �r�{��ک*P8 ~�!�d�$�B�����]�LK��}E҃�=>�.S��G��X�%KRi^�5֑ZU�ήWX��"JKJM���?5�T��K���l�k�qL_zS��K���z�#�#|z��mpxw��=�Km���˙A
�Obj�y�}ِ��(�ޮ���RL��A�e&⧠��9�0s�qj�Տ�ڦ"06�BS���:��B]��G`�Mj��[��h��@]6]�b�9�ۆ[A&t����D#�Qhcr��R��{�r��.F����%bCe;�3�HG�W���ٖ�p���E{XlxVHYEB     400     170�V�ێ��8=��O���Л�7;���{?�?]�����wS��^v��hO�6K�/�x��.����5���q@�E������a��n�+�t����̽�������'e밒C���
�n�z9u�7����}s�mXԇ���djpY,�u�r��{Ց�"��J��vv��o�=���Gs���_� o5�*�ܻ����u��5gBv|��#�ʀ�g�j'��F�:=���:@~�Z�b+^'�cx�Ye��øꎹH��	�_�d�T�,,1?^�?�+x��='L9�B�<=���;�t�k�E/�_�.�'%;���y�Ղu~��n1ޮ��b%�.�W����o���%"���w;��r���9 �^��`XlxVHYEB     400     180�oC}Kp
�\*��gM��z4��h�F�jZ��F���I�U�9�>#��tI����LЄ{�}��q�n��	0�;���c� � �qn%������,Z��c�Pbx/��q�<jnGO���g�¶I_K5e����-d
_��N������Px�`��9K�g�a�'����B~�l�cM��a[�-񤅤3OW  ��v���֚x�ѫ@C�,�a���/��@}��˿����ʔBK�\��PY���8��	�`c<�&�bu�m�&N[r��a�ϴ�"�<�3�3
{h!�w���a�|�W�$Y��1�,�q�5a�I�4��FI]¦G͎I�m_��i�H�H���,��t<6�c�ES (�J�XlxVHYEB     400     150!D``�� �!���Ӏ������^�Ɏ���a�9����?Rhe��5:2ׯ�I`�B�1�^��m���S��e��tf����؊E��#8�q��{\�<� �!)�d`�� ��j�����>�`%��-������nc����b�����X����;Tw
z޴�k���3����9Z�:�& �8��!
[��	�`�_�@�6�HV��hb(�f�FF����I|F9E�
Q���\��]�IQʢ~G�{����O�r��	ڹlT+�@�nf5n�\�w���kq����|�"n����}`�;��A)�w2+ǉ��K��h�6��ߊvU�P�Y��K�B�XlxVHYEB     400     170����vȎߡd�Rc�� Y���j<�dc<��zp���p���j�E0��%���������n���%�7�֐�f��5�n���H��T_q�]j�x�u�Q�`b�}#6�2Lݙ�iFbMD��Y�i��Źݟ6��_�A���|Uh�<`6�x�2�]]Tg���}���x����Ζ�,~Z�5AL+���~�߈kM�ac�V���yC=Ȩ����:J.���;�������X��Ld��ڃ��Get��F��	�&C ,���tV����h�8i&a�,��4b�#��YظT�z��lUr��Ə���5i<p���`*j�>~H�R�C�wg�I+�Q�h=����Φ�dK�z�����2Y��XlxVHYEB     400     1b0e<��n�2�dvbL/w�ԎQ�[����Q����hS�l]��,Hi݋�U�J�gu��(�27���=�ˑ�"_*懋B ��ط�W�܂l��θʚ��/�e�}�K!Ґ��~5�x���[>����f��:�R����Ƒ$�ߢ9H��>D�%��
�mU��t�"�y�6��;g��C�<1S)�"-��I�ʗ�rq4��P����|��<;���ex��P� ��t�3�<\yb���k8؅"��3X�g0�Q���R`ʎkL����icԌ��m���瘹�mu1����k��h�����4�쪄��DB�����f��6?������Z���7�O�9�["ټw$'R;��>P$��#n��z 	���q��3�?% ���r>�C��A�X��4�
�A��xڰ�ż��#�XlxVHYEB      e0      a0짭cc���u͢ZU�-1�C{�w�Sm�I�S��>��!��z�92#=���V�WI��h��,����؄�$F���H~�q^�-D�h͎3�.��(��0��h4#���q�����.|���ܖ�.�K�j���}i{�ѝ���PP�,�|���Z��