`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
op76uB8dP/Oo6RwDFw96U0l9mHqwp6JqFXbYzeBkK7chNTfsZX/nCotsLpPdzsS0TecMVvXIbECe
VS+fy2EUZ3e2RQKvpkho5ubAfZTXYCIPqwn9u9oxRVLBUvx88yFEsbsXFZQcPSiR9oT94gYvDiJi
/ehExfpOG7/HHoqNUkA/1qa6jPmYFCcu93y/ClY7V9QcuyuQ9bqexTLH6j5DI51LXkgKQlkMHgse
e9SY+jylKqWVJs31mMQwoD1ciENdYpEA7tnwVvtwVanyuYw6mbduBsUFzH0prP3p4Zj3kHvYGryT
+ANfAVGi8ciyOyK+sIKD4SOyQTOuPg9CWREolA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="UyeOUSl7p94f4QcP/jgmSniktWTDYhhUIWqm8oshj+8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2464)
`protect data_block
YL2e618SgZ/NAcByvTtF54hNGjcGAbNRelItFWyzED3/bQVWk2093P8Ljk6flBanZGxDjuI+0z8l
r7YoK3I3l4VK7e/Ge4/iTSSQQuqqmymXK1h6sTASeDWUpV52AvE3/zxysN/NgDmDsxLvTp2nfpok
3HBpR8HWl8R5Zl5D1UvvBDsPwWn9x5t9Ce/1ixJvreH+y2I/Y9eMZLtrGY0gZQsc7MjKIsguh5pT
VrqpJkFIcS737PSKtlIAMsDYA+xIZ269YnSzjUtz1id76PXpMD7LAFQ0AGFwo70UC0treVhXbT+f
w11JUXfs+d74UxXejLl/xanwshdjUbaFsS6AX2YKUEcZUKl/G/vxBUHLGge+jtytH0WO1y5Ho2SX
JTvNKT8I8FlVNcd/RcneZxFO08RGSbdnQIjgkqfYUQ1ERfqHpqP2xMZQjWbIe2+Z0dxVuPxQhPrG
eZyWb33dUd9Dl/3gbwb7iu6BffGsRwNc9w6blVUS926Jg11huDGGKGpXugktwgmVajtQYbV8QwRT
LgTaJTVDrB7tXtbq32WA2I4hacvOlgOhsUhL5XZ3EMEviZ47z3pa/fiOwcGjqk5zcJCr9dC0oSHC
0si28uA3r4HoTNp+eC76FywMMHUXNo14+iLs0Nu0AhZMQO17hunsQWoEG9O3RCg+NO+A44D29+Fg
pWWLsDHzUKGBo83y7Vkx6nFNtwvGHP88K3wyLv5yy5es62VQ6dSya8A4K6kvd7311hhqvfX2TeSA
2FlyzcKkjEnSkkfou+6uYbMUUq342y1/TFZ8nyni19mkTKQM/J/ljThRB/H7SgroGZxmkFfbxMf1
HTNOrMyayZ0m1kcLPbbW7YPhe0EhD/Z/LhRVtrALi4JnYQPZGlVDGIgCjBFYnwtxfBLWvQ73YaWA
3/CqSqRW0JAFUlBNy1pF+ie9fLoOoa36GouBV8/gnIdJ+5XDmWfj1DWymPqdlRD3ZDkYzUR0xB1w
G58BdLr0GdPJ2D0z05pmBYdE3+xY/+ppxZCAYAldU1c15m+QiOPABjq9Zs5STBP1QxuroqJCRhzI
Bh39Jx3ZJ4VC9dzATq42t5WZlN6CIVpg2Kf12KAO22ch6usfq+V6P2+ccFDpEvrRhXTWI2VAkUjp
1e7yqyZNgRGMy0iO/pGbGGoH0um65mpcVPVHfVE0m6Qbo9z1vV4YT53xnxNcwD424bGvUZl9T9aA
B3NTHx/drZaB3R07fdR2ywlPDSaBZ0P7C4yqgk9sz3XIoRMCdxTonK6qQFc6zbCVYc74/lD0m1a9
kMT5TSnQAyD1MSp754Uj1X7zxq+DKAZ4WBYhogdiSy5VyrbBhsJUH8xHASP1G9uD3YsktVyKU9pn
Kr9QsEnQcoswYfd233fsCYE+jG27orq5clPz6hEmU8DRR28/VwuY+wNmvv96DPv3ORGl+2Aal6/O
tYozfAa4VJ6X+4FJwcsVBr2HQfbaO2kB9qltZk57Q5Pr0a6vC46VDF50ni2jGsTfaaJRD2K3WpNV
lQNJz00Ic47R1gAtJVsGazimodS1K0yDxfCAA1nbOeglKo+zlI/JYrJYXnJPZzKwLt35672UJqYZ
nszeYysSredm1Whyj/jAEsAjpFti5l4N0LeM0yxkmpLkyQCVkcz2wQJ7fLkEojlODVevDPpM/Chs
gNanByR5A/4tg3/s8cNtL+kvQW2s/hi9dEIcxJICmVTGhdPq849sd0oinOfLkF8j0FOW7k4NMl5T
WSVCYBlpeelv7D2z+ITeNKKUxQKYViRFu1kv2FDmZzpAV26thDT+97knkaQE8UeeSTP3yrhtHcKi
B1sPykGjCAdQBBcngBtNQM8d9u/b9CjE43ira4IfL7/OpxzskHAimKlhZc48IvlkpgC7DQytIc3+
jKKzMGQPWRfNvzeImEFxvak4XiSJXisKHnZL9uaYPmp9ZCiD/3TxNewVIdy7115EXLqg9d09SMEy
K+Ql0z33LtLOlCo7M53FNezHVTEsmCPc0aC+gYaeLeNp2sWf7rgUEuILfrhXE87YIZeo1ciOT0t2
sZPEgu4Z71mz2kBxEEFPA9G0OoKAa36TRQ4230ylZ8P9QuBCcED9WiGvcGd58j2D8xSkmyE3XssE
j38oKXZsnBb3kHu5i6WgdpLKTeA7/w2kzdnRck4y/VVob7GiVmSooODX6W+GMn61GegLGcyYOp60
XDYMoOqweM0k4wDWOs1s0cH5N4tBvCnDzdR3JEdpyPOFmbf2sH9J/utUErno53Nt5GSQHaeoW5Py
XIIRo+fdHDDp0ySNbSQosXUm4KUERpkE5w75TQQAW0HViRpYjN4ytWn/4QJXz+mZXSNZcXg1asvP
9W8/59aX87NlDP1q/gSlJ01lP3/vTXUjaoVawDNKprtM9wOFsSpDuIyvKnJ16f4a/7xKFmcgLiYc
/qmxhECKLo6i9zEB7EARgyF6PQHs3MZeOA7oKzCCbeXkqgVHrcDZOm+WDFa/FkeKqujTqkAgRNFw
TqGOjdbaYm+QXp9nj+3A/wuwuQy5DP3d8rKFe5g9dZ6BTBBHsWJnVi6jYomkb0KWjWA+5HdTzEkT
yUAhABsKFL0NFQzNRBQGOcXRfrmB45PyF4pfZfclzatH9WkpIASKj9v0L/mEuQY/JB14Ht2euPiY
s6CzEn6DhFFPE7EiIrjeMuDzvKhw9pp7rj+XnlzAfW4EnD5O8nhjk272VnOIQfcUrgq/s5WnnZHb
sU4wmy6Zfih01sIVQBUL+SvRgy3XSPMkx4urR/RNQeFUXxGcDjwSNF5Thw0FvEJlP0+f864iucFI
OFbOKBR2Co5rJlYm2L+dd+AIl8IzUl+uyWzD8VDiGuGlv3TPplYp7gCWMXUAkI6/+gU/Wal1iwRt
7bJpMFih5fjT3T7YK1I+OZ3kUAVlAa0xJa1Z/oXmjzjYt720UbXe2Q/Q8r7x6qFopT7mYK5dp9yJ
+y55hKZv1IifoQRh7869Wos1ukuYUjWbQWoASDIQP1K4ypVNvdq8PEzAN/OsC9E9a9MFvtFUZE7f
v3x5ePznhoKBwWN6MqmuOKRIq1W33nBaOuTPv7ZO4qfePAniwGPWwiPMR+QSjODkCT+XPIpKGXVT
dZX13YFqNN/moUyGcrrnlulNPFU+Zuq/zaRysWOOXPYtoGaCkMbrOmmRb7WQkGmePBI+iPpi3fyX
i2HBEp5l0eASu6j9iVXmGLtir2GIo1NlhM27uE+aHlvGCAXPl67wK8UVCoVuQ+6arMDpHL0SWjCW
PngplIked+EA5UfbEA==
`protect end_protected
