XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Ѧv���<�J;p�{H<^?�|���ѹ��2L���*�� x�dH@�@gw�>�D��|C<�Su����'5ʋ{���,\�����$CT�9Z�&�e�cC��Ě$ܝ�A����ђv�7���L�\��Y֧]E��w����B�o>D�U��|!�����.~'�������o:%���'Ӵ�%� �V�HÛm�I��s�ӕ��7�k6��@k_��&O��7�_�>
�k=ǆNM��M�i�ھ]�|%u���� *Ʊ����W#a��a�������K¶�p�*�u%�ڑa���m��"����W�8Y�;@J�$(�o���]���3�f����n͇��B��z��k������z�3a���;���H�ͩ�K;�#l�� �`�`�K,%��T-�C� �>�f�@4��cI4��2�n�3B䉻E���)	#��: KlŊ��!T���<���i���ļ�?U'���*�]N����-s6\{:TGC����[[k.%�Q�,�?N�0~�� ������H�{�v��@�L:YՑ��y��x[."�F,������{8
��㘩���o��Ӳ9����f!kU���(r695�HsI��|%�GTbٶ��q�,�Ϳd��z���~����n����X��z;}{|�E���>>�3C�}Njo/2�ap�2�ѱe�ڝ���D:���U�~р�K$��K*��O�q
�et����¶ua���v�R_&�Q���|�XlxVHYEB     400     190ր���[���3�%����@�:��6�y����Ϗ��Ih�L�A@�����Z�/_2�n����Hq"���Q��D��^��J9yNmG�2|��XhXG���QŰO/��l�i�n&���u��1PU�����/��L8ֺ8vE�_�_)��c�ŀ2�.q�����4lrB8"�f��
g�Џ&����ް��s��(�V��* ��Vk/�\e.���kRk�^�JH����u������-�o�N�iQv���g)�W�N�g����?N]���Wi�����rںq��w�ɣ�4�zX�W��L���������T4	��n�ɵ�	��E|���51��L�s��M�����-��Xo��2r�9@M�KN��_'?�|[+�	/��<��w*��T���XlxVHYEB     400      b0�H�wSl<3Rrp���&!)zclD��e:W��u�D`��Gt� �����%V��)�����GUn�)��@a
��/B����|ŵ�� �H�$G �'ɚ��M�i@Dr{�S�Y�A-�b��sL
Zb���I2�����Bf ǧ��Y��m������\�JR�%�XlxVHYEB     400      f0<�yb"?�z�#:To�G�6S��q<a	�ڗ����Գ?�ু���S;�K���,Qu�$��* ���)���*��r8H�O��#�/�U�uy�z�aA�f����Ĕh6㢴h��N��wOyiB��i����=�f}�h~���iR.4o�Ř��x�+P��P2��퍛�^�`���T���&��q*��lA0,W�:薏�P�-���n"E�⑎?ثmױ��Xb���h�G�XlxVHYEB     400     150&�~(?�\b'���j��<#*���gS��)Z�����:�b�UB1T���=���I�B���-���(�꟩��;��E�[�U�߿�8� �
�A�*��N�[x�A�����F|s\%�"�=����U���vNz-�|��L����`ݳI�&������HV�
���s�� �����9�v*"���N{4���ީ�nJz����GB���l��D�a<�R]�V%:��r����YF���',pm�f5��M{����jO��+<:�k�"?U/".����&����1F�Γ@A}�-��^Ύ�|IMQe�R�1����3|jj1zXlxVHYEB     400     160Q��g�ݽլ�}^+�WL��R3�D+�|������X���/(`��_/��pv��m�?�t������9]�B�K�1YV�T�o�p��T�@n�}�%4W�n���ǵ8�$�׶X,�m|FZB������&��2�Q����ӵMĿ@���#4 <�b���x2i�&�9F�G��j̠V�c�ڙ㽈`�-l�.g[N��.�U\�ǯ�JT3p��ȿ��F����ge�hq��Zd�l���ϗ�:p�,#�x�mt=M^xGH\5rq ��YՍ�ʌ��q��3%�y;��^���<�5�O�\Ԗm8����	Ss���FV�y��n�h�C&Q�\-Y{kX�XlxVHYEB     400     120D�Z�0�ϖ��ZGr��3�8��tE�NOC�� h�xK<4�W�˧\�+"�7�C+��MC���EL4�9�a����/����-�x�+ݨ���y� �t_C�EF�Ÿ\ugB�qK{�l�����>�[�{���gIb�[��M�����ψ����H�bꡓ�b&Ȕ-g��� 2�zE�J?N���ň�Ɏ�ǝ�֥���yy]�>�D�g]��K#"��gX¿c	�	/Mo� ,a��]y��D���8?��-8A�sz�����UP<)�nuB��XlxVHYEB     400     110���T���K�!�,2"��!�7�/�v����Q����FS������;���T�+�ڼ<�-�xE�i�����g���"SjI��7�%jT�0 �]��Q-�If�F�� ��e�(gb|"
����s��q:D�눨�7���c{t�P\+:�
?a��&1�t,iE�����i�{�<�φ��e.�)�.�O�:�a�uԱ����M��e������z 
n=�Sh
�_H�gz�9��xق�
ν�N�I�j��pQR���j��P�}n�JSXlxVHYEB     400     110K�Q�W�6���$�K���$�*	���	�D �"i��F���Bo��7-�����q�ؗ3����Ҽ�Ϥ����h�����'%N���"����7��۟u��@�m�]��dL���M��G7v^�rԬ�ǎ������ $��x˔�b�+~���䣚>���_��
[%*���i��R��O�s.��{���&�15���S?�9���6ٙ�OX�� �<˨�-Q�O@"��#���{`X�RM����0�#%�b56��a;�<i��EаXlxVHYEB     400     130���_HG�}d%���P�]�����oߜ0��M"~6����>���]j�k��n\�]2{2��π��O�3��u�����1hʎ���>2"F�^���S)8z�x��9�؛�a��	�D�쁏��Z��>���#%����(	MT\l���Ϙ�M�_s��u�c|;NrM�iZz��`#�z�\U�^Xu�%�q$�i�����Ӄ^���rϺu]��� ��$8Ȁb]���F0@~��2.�
Ҏ}"�Z[d^��P;<���X�OH]bc",p#]^[-�Y.D�m����Dqŏ�qXlxVHYEB     400     140騴_��b��8���%����VK�k�"���<�z>q��MzXw:6�����p��!I{C�L�/��	���ь�ݲp>r𛂩���/���q�5��[+��9R�"�1���k=�R�hb�����gQ���	�6���I"���S�yI��w��>��x^� H�x&���.�LG)U�DL��FI����3�X�h"���}�]��D	X}�1(�`$%�x�  ���	u��v�<���q�7��1�t����t"�}E*���"3|�A]O�v�b�ra��`�	���s��������!��0��$XlxVHYEB     400     100��03p@��r��DF�T$�@~&8}��AK�3�5��N!«W�.~�����S<���d������X��`L"�Tb��������9gy#'֟��jKyO wPHw+�k�M�亐;������J�Ǡ\� +�N��U�\W)��+�8%�XI��GB�������hvBm��<���<�����~�C��3^�fJ�
3_:���h���-b&�B��4��(�����zY2hl)XlxVHYEB     37b     140��w����eڗ��P�O�B��"+q)nwRҒ9HG�0~=Q��.)�$CIS>��=�1�A��_6��z����Da��q; ��9��U�Z.�ۥY�^Ͻ8
WUh҉>NQDt��o"QE׹�b�]42����`#�D�a���o��0�R��^�ӛ�m0�`�L� � �Ft9�� kb5"$�L�
�.?a��������o$6�&�d��?�{�Q^4	`䉻�"z�yٽC���~�~AN �����fC���4��j6䇙>��6͈��>�9LI�cF�2�?D!�ɯ�����aշa���qq�����