`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2448)
`protect data_block
IqDPSwFvKNyNQCfSB0aS/31ZWGRByitrrhX6fgaK4PsUiUrBUPJXtSYi5A0Gm20oEP0v4DwzCRny
+ZeuPQrDU+vsU2T3sad36egRPmx9ITO4xFmnFCoC4/rRsItxzO8EtB1Jy0K4tNHYyl53RHYkJPd0
8ucGck44OKkphMv0TVRM1oNSZJfBpb3HEcQff0Bd6WZpwpzqpZwCJ4md5nYxL/bNjRpZpoohZHX3
bWaUcb5i2empG5IweVCWEK+HFgJNriQdJrM3AeypKf+HmOvQ/9dSpIUhAwhObU96XiTnZRO13on5
JyijRd33caVk6oZ70yK/kDBoCurnee9+F96278KBQeBvxR8LYNx/zT+ta/7xeool8BE/5du7XdVY
Cju4uQnVlfOi6xgo4tzKwmlHt6f0RzdM1N2LBczf8uCR/T9m1tR7ipXTMWB22gdMPfO3JmMKWvP+
udB7HisnPGTmDG6GP1EHIXpFZuEnGSExO/gfdMiWMt+jhDktUCL7LTc6/Cug+x7ZLd+iJyxoK8Uz
L9G3YUmHtD085nKFelWhRfKxGIznM3Zy90zBKgLfcRN6zVkpKh0Wsx9Lo0TlC4tdd+c69MTFOX3r
0uX7Z4Ebd4LUoE1yDSx0qKDkySF59TKDfq9pF2jpIuWuX3TBcPeJRkqJpmDgiQBjJEH42cIbmCkA
Z4/S0/RKyjUQDciTL7nfy+mNZX/ccJ2d3EsFXrAI5co4iAZAYxWaKs9C0O1EKPS+X62VES0a+1jT
a+q41VZJdC0Pa25yuKrfxZaSaMCPkWBxbRZi4ljNu0/MmmZgpAK22obYl5gDzSYhxEFIjsf3GEqg
BYbMQ1juPzot3ivT7YBEzdZmkvd6bl59KvwXeosCBGAuac8/vb61A1P+q1JPQyN3uKdOa4qm86z9
JgFz0/j9fjIdmiuvDRv20MPd/iEP6KYIlslrJYRJeH5ON3rxbAgeSskS5AWD0105TYSJHiTsLi24
NTdYv9uZsQwUb3bGdwLixAAOexI6cA3hzhUjMnI92aOYcCWsyxtIPI0qMhdunBa/PVNLPlV9ZAIj
eBH7yF8MRMU0bmFrBXdOKepEc2Tu/a96QYqBlzlvJaYrCPPXyhChGPXly68zinJ9sQMxjwOYu595
gpuL2GsyaiCliOeCKID9VhXEdqEdHUcs4yY+dXwewEmp+8pOzvKgBwluDp6jlqZ6omB9JnffIaxA
7zjv8QbJxYluw1ZiYLo3i+7TP7VHKfU3NGnVFtdahT0KhgxIJmRRUEndw5nGvcKAnmIKKplTXvfW
v7eVwydpIA65G0rqertR/DwwcNprpgRxHvIjt0wmQglCSDZ2EctfyBhG8QGL9vNMjh1KDjWcwzqH
o+ZTlrHTo38i79/LfhuC0ZDdoYe7gdec9tjX6vxIsPnJAdZzrShuT8F8XvGlQoqsk5iYNy7SMmd8
yTSGMgESzeswbr4/k9W2W4A1ECtNZ3GDVA7n+rFH9xnQuLvkegUagWkgyouWq+vRGqoUykfNBeKs
21cYtCl6yeOx9QK0nSmZdtmn6++Q0wMw8uVlgPjvl3OITFUOJHBVymagw+LY67H7JPV1P9ngBC25
fBXLXaJbAxSDdTfZX1QGFrfWmG0DePv0lZRnt+1FonjR2Rn6ISJzs7wwzGU24nSa01yFXg17OzlY
NY/RtWRCUkoJs0U1MuHguVklFjvZBGtBAlX6AMgrQzeqLZTPTAzV/r/kVxZ/pgJBwdA6b8Fr33Xv
gviCILEmYt5dXFaui5wne5q9eLbmFteJ9dxk0XT6E90xv7dzOzNxopYtlJuluDMtUbKX4XepLe6o
NKfO0siKKpM6wC1fYAa0oWe8uBkDtFlNTU5uFSSH2D+GDdqpoTthJd4RTgqCyYiSLNESW2AS+ORe
5voiO6dasm7B3VOwjraGHHS7c/1fCAI1z4OzsErPI1UkpHvVzcvoRhxrWbqGfmhFMQBuvAY8DYMA
bK7U/xKteH7WsN1RM7RAISH630TCd0heJWPFRf+AIfc/+C7CRxyG5AZdF2SfALkF/4YZuML6ORHz
UIrix8PgDmEda9YoSHA4/pVc26L6LoRjdJrh2RKmnVgqwHzFgahMlbezYEtqsC7RaKjwIdiwzhm8
Am0QSlY5V+S1Ikv7585ElEKBl1WSdXi+22+o4/+BFZAAGES10vQG2SiOzy3PkfkLdGL6fpT7HtZy
KLJf/w6AzvoB7b4L78rV7pvFI9alIOwQJnQyTgNXSJ6CWbZ6jSgZ99asJAzQ2TU1QIOT6TCjT5yY
qF4nFmTaiiTe0qX5c/X2LAAkdtyrUsUvI0sNSS+Drvzq9bdfw23grgWCkFEba4tRk6bfjE14cSCP
ur94yO8mgA41RaeBuzMnkVQZrrg95far2ZcirMzuPyufOaEIaq3ACK+c+XCZgtVbF/hbixm2c0+4
NmAxJfdLzUIKDqIySkhwmWKTd12dxbRs+n/HFWX1gPCgXEAogwdSbqu9RKq3mwijWbbzuSzMwG5w
DKTuq/zFJKMLxLtLRntqVLdRbZOTn/za98WEY3wDi4cWzu1fVzYjiW5QcNdBGnd8LoupnwRMDUW5
3YTX8FfkTgnf3hxQ1PXRnE19fQXMqbLMcL4CpgZQ1bUzTgeLN1Wmokw2cNciOnvHWySBk/epcCQY
cISiB4gMYLfVW+7mwP1P1hnHGS51Dxy3ZTaPb0hZZgJPVfT00KBk+S29GeJMrbOG+PunOgnwzFy8
P0p+iI8os3vVU6TSUCqTucb23Hqo6+FlRveM/3yZcGQKu6VyDzL7TcXRE5DHD8ZRjl9/4n5XnjI6
byyYIXWqXgtc3TMlwZr2iDjEVZXbuERXwG7jLdrJWmWTvMVXcFNal17vL9dksYhrvdev/G+os5+m
lXV3mPuAqcw9KoVNDvuJI3n0BIJpFCCh2Q/EIUp0W2dDk+IwMlAyQi4MwtUMnDqnlnhscXu/9wLj
P8mVIMo0xrVuzmIlPsPgLMDh6YvzBpv6+QYx1nytFsJEdvJE29+kFKUQ2+qhP3XKb7tmXtAQuJsi
Q0Dujtya+OCU6gd/TrWiekPvFt04isPDoBK8WD0cD8IP8KY9cHhTmdZsQANu3XFMBkWB0ta7HoqP
ngF2IHm9wL8Ak6nrNJXpm83roBOb62OYYBqBDo7hE7mP29rAuOqhO8ow62ITvuJGV+UPww3SGLzJ
zCIj6d36XUkR0ABjManre25mgdAPmHR1BtzEDoAUtSf+LZvcnwmryqyyyJjTzNH5ry1E2EUg
`protect end_protected
