XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��9��A��
���)�{m^�w���Kﰻ�Y!��lv��zGB��m�k��̵�X�О�F�����28.I�����]xo�E{��
B����f1��׳w����@tl.]��M\P�����#<��'��閒?��L���~�����*���j��0w��������͚IB:M�lq���8=rٺPoҹ
������-kꋫ��~����/ŐZ�DTi�ؽ+~�
b�����
�fF]-�"���_�;R>"�a��}ɼ7U��k�djB��*������Y�#����Gǫ��bY7����6xFJ5�8��5B�,�`'��Qw�R4��g=�rt�:����+~�q���v�ա��
�7
�������O�Ck��t��o݀�d$\��%>� �e&V���KR����W�A��e�P�x{�e���Йt!�ۻ
�H��7�+���m��m�u����U�t�T��![�"��.�y�H���d� ����2u����<�!g�Ψ}fސ{;��h�;�A/dѵd����Y���(�&2�z����Yc�)Y�v��u굍��^��%'Zkй�u/��}���g4�s��1�
o���)���N�"��
ȷ]>29?�t.D��}l��JA�#EB��TZ����LL�Z\#k� d�u��@Xnt/Ja&��z�Ԁ��ڝ���~Q��%%0�J��;�07�:�ˊ�́/0�Fq)96^�Q\�T����zJzn>�w������!�������!kXlxVHYEB     400     150r�G�I������/��d���n��0�b޹��؋k�X�Źd��l�i�]"�'f��:g���}yO���>�P}�\�2�?Ǧ}�{�Y�2��o�F���c�W�	�$ä�ƙ���ӳ(E>K@�5LI+p��>Ͼu�����G��2�&3�8��4i3���m�f{{f�o?����l`�޿�<��®atG8�����,�=��������\��"<�޲�
��u�J���lPb�nE�6ǼZ=F���RђW �k�7�%�p1;��`����Ή���1�zn�5%h�chO�y|O���4!�w�d�+\}t�dS��
�^F���CXlxVHYEB     400     170i��	��̳5�p�tLq1��T�>����i�"�JP�K��l(D��B.�h��.z�mku��\��(H/�i��8�+bC��B�V�z��|��Tjd�h��̌�Ε=�l�njV�,��Q�S��I��D��q�t�O� ���T��ԃRn:��c�/F!}2�kЅ�G͇.�A����$iR+/��NJB�	f�5$�Nm���`��*=����;6��9J��È1����O_���=K�T(�I�g����(% 	�N w_n�
9���H�4F_��d;�'�OC){���Ex�IK2%bv	��2rS������gۈ������m�S^�5i��5;�Q�{U�U:H
;�sg|XlxVHYEB     400     130��	>T�
�����kyC �AiP�5���0N�u�x��lF����[��Dh�Jgc�.,|W�I�uqWt��`��P\���g���|�*�R"�F%'�(�IͩW��xnGު�|�K�Զj��u�c�C�U\�@�)���LV�ۄ�Q��[���nEb�Q���&�xn#PMU��g�8������h��G'�tA�ɳp?���1�����	�5��H	U,3*�wA�<@kg=&eu�g�����l�:'���$��v݅�v�@}*ۖE�E%�S�'Jg?C�i�|5=�<0=�XlxVHYEB     400     100�S ؗ�(ҏܻ[�t|mAT���)E��:�[������AՊ���	j�,���D�Pڗk�����Sژ@H�	�>CŅ��7uQ���_��p�72دc��A�<
�"	�)<�-M�s9r@_�wk���<�D��$,1��В5Ea"V7�lA��$�<�ڠ����1P��Z���1��3�B$E��k��pN1Ɲ���5�\3)���P�Z�;Ш%>
~�v:������K7��Z��gQuOXlxVHYEB     400      e0�ö�Xx�m1���b�Z��,�~!�T��� �uxBfD�3�=��g���S�	=A��TN����.�,��Z:��2��읡C��K<��JNB�bKn��kgNRM0�ۍg�{paHyX\&xIUz��wtDRj����2-��IYUcSaJ32@#۴�ſ[K��E3����IT<�Ěke!�mѧT�%q�V+�d�!N��I�ـZw�v/��4V��!��:s����XlxVHYEB     400      d0�q/�����H1-b���ѮeW�S�S:q�I��V�{������F�������i�W�)D9I�X7޿Ivr!���:o��-s�{{K�B�/B��?�}'iş�^+.��+x��5"f��%ͭ%�6�?�ZV�x2n�n��ތ���Y��OiL`F����ZX��>����_^����A\9�u��gf�9JL˷�]PXlxVHYEB     400     120�V��tt�A�^�:RO5c�CB��/u���W����1X=���9��I/7��F��HQ@�`-ߌ{�~#��0��H[ ����dTf�I�Gb{K~R��7��kp̉N/D�b�Y��*��?`�Y�����L�h$��<�<��E=ap>@Mp�����c~L�aF��CZ~\�<N�a�R����BAv��ܴ��)������r4�څ���|�&J���w�V���a�j��iZ�c`9��y~�?�X�h��RK3��rf E;�IS4z�'Œi��|ߚ��[�Js�J�m���dXlxVHYEB     400     180fT��Ώ��H�wa���a��jm6�����x��Lii�$P�G*F���+��N,%��)bR�P�0�q/����<Q0�u�5��ѷ���z����r�����P�z��uϱC/2�O��΄��y�w�[y���gM�W���I���������S���$�¤��,o���يC
�&��)���C��O>G�a%-LZQ�ɡ��O�O�Ju�10�,��I��UJ@&��s�g�G��C�2�1�/���0��S�]�F:jꁟ�(	���k�M��X8��0�N���z�`����~nf$���p6������
��in}82�e�OS�Rf���dgc�`B�(���9"=uޅ6��[厡Y_%/�9Q~r�c��	iZt��k��XlxVHYEB     400     140�[���^�<�VSr��I\5T�-�0-�pg�>-0����f}�4j�[��~/� �l�G������4^z����#㍂�0��ks2��*�D-=���Rr)Q�+��!��L��~qۦ}L�����[��G��֯�6��G�`�ʎ��Yӆ&��|����{�:��x�>�Rp��j�kT��y}�8Â�I}��&�z���A�*��ҳ=����DB�=Y4i�?!A����Y�b�D@�|E��g��+IM:��G���#b%`Qf�:� !�M��xD���r�?�FRb<=&|amW0�4�����aXlxVHYEB     400     170l;�H1�S�I��L�,�3����f��f�$wVx���Jb�|�դ�ld�D ϯ�ޗ�1�9�>��!hd���FdI�ə�hX��@��DV�+5��:����L��XV���kN^��{�������� �B!� ������eelY�d��	�+	<p$��V���$���)"��p{��t��_�B����7�A���N�f_�lJ���U��˄K����W�	)�x+:<;�vϚΏ�q
��Q龷/��|�q#�`�}��b�5Z�ꤷ�|ґR{Ed�.�V~���f���C�����0������7cQ�)ά�sܽmn#�t'�a%F�l��ɘ����t��IS��G��td\�~����^�#��ص�XlxVHYEB     170      d0�S���w�^/I�O�� a��z�g�r;�7AC%z�<x��R�<7���^ʸ����.Ԕo��Eۮ'�r��F�\_�3�v�Q�,-r��J��9�}�	ʽ4�Y����Rk���3H]�B&��6�Hx��q��Zhc=� 8,���/65c)RP�5;q<���yP��޾�z./J�˔0+�~�D�1�mP����3���T��O���G