`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
LvIP2AR4GQN4haxnGVoEzkX2hmbnzfqWW6gzNKxEaaowykee3XP1fL+zyH4SP7mIRP5Z1pXDD2vD
5ZQL8DWu5w74GjoyKEz5wbprGifKrj3TFExmbOpT2zmb3kJgVhh/AFDO9oG2vw2TYuio9+ZwMwyj
4bPZrAKOmKW+LcCeQCg/AlGG0AAWBmdY9mBPoykm0iN/VIg978iHmpYEM2iqRG/VGuo0+4loaRqh
rJ+Lg3xAqBOTOCHcBbccHdjYs3MafzDq5O6tB+VM5ar1DqWsZzcOtJoQ3/BEWSsl65hNYeYHLp3T
jd+dg/xx/cLSG8f/8LuC+ezxArmJ48zexTvOxw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="uQdyMOlkeL7U0xEcFKWgHvXg5KcTyMhgMXXIvifMM4U="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7488)
`protect data_block
U/R4upwzNn8aI08nPmQfexnstPw2dDZU6ul9tDAZkH03dNHLRj9SkTqzH+49Q2idBPkLNzaGM7wP
UBFps4UwSTDM+Qjf9/3xlVjyVaH/UKTaWjkf4RIFiJdHgwcz7rppsgy78STLQ9s8wTVyYyP0Lo5Y
vinDhGXI1/JpLISOCYYt0S/kziABKJaCF/NKinTr5RB6BuPf1Xuyx6yc6T029s7EqlO26i/bLwO7
/8FdHsKZgQpkGsxpQ5qoCfdA9w41fNThlOwaYR4H+5aJz/Gk9u3sNTSYNbMhM3D1rDS1pNx1WIA7
Y9WXBHOO4RY+m04tuAzPnY3HDJdnrzIe8iiD3GZAr+ZWGfmhaL325m2IW2A2/vNYpaptgPSweZuw
uV5BDydOqnblF4A5OQlekph7y7zNZQpBMu4vDwwmOy4h6Xo+h1/7N7I8Q/Q6RTJ3oDUxpCNGF5jD
cHNbTAEh19DdrvdTLqj7PCrhv3BjSgy/i4fxREE0KX3h1e2Pf+Q7gZj72ZGE8DYANDFWZMvIPWRW
k63kaTgz0m8TGTW1DKfGpTyntqvjCrSKPFqPJCM+caDqixMXu2ynG39hQeQeT5L+MQXkd2SxLceC
8Wl/dcTmDnIUb7yCnIAyd1c5Q67upQssaH0qQhAUnvmZCjUp/vKx14j3QhgkTwcjVTHuRELPenTi
wsyWOpWm1LEdVTyIyi4MZ6D1LIbjvum520BEaBMaMSOo+7iG8TkeqOqBFHq1yUNXO6XHxO18UCuZ
BXDsn05g1tt/NFv/G+Zrok+5IJRnMnRzVqh/ZK0S7RfoyqgkDo8MVyfhtOvh+5dGj2gEhGCdyaCg
C31ITUThJGxYgPYN+ZBtXKNtd5kpyEn/Xm1/62JeW5tFyy2AOLCdFfXdl6nTTCWDm2xOHPWIoXJ9
tyhvcM0UGpDw8pp5Goz+kM4Qz8LLDqBP6AX54UyR/iouwdfy4ErKOuJebatpRgedWtDOenwmvXuL
3xp6WrE1+nniOeM+bur+AaQtPn9YK0DzKFwbQe80UiMYVg6aNlin9akGoo9fShH11reht8dU1AGZ
e6Xo97TrggS/rW3Gx6fuet7m+BqBV7bIHNkeNpvddvffO48wHFKIFRor3SK7oVW2lSsW5x+3HFKD
bnKT0NRQrBkHenkWmSg2mIpPJLUMospxVM3ZG9xSvtxL7NhXvyfsvSduTYuJqi58rKqZ/jaPbawn
Or/ERxGJbY8f1+rgcbz6FsvkJhdZ1bBw1DNCFrLOzi6QT6AKIruU9xZmIU/O50MuHKOxKy77x4UU
wqcvEclW+Jx8DUtoF9v/1tmjuVoXTpyMGDzBevNlEIX0krJRt576++3Pz7RJ6zc0MzqzP4InJqaL
tgdfFZa31mVgapasM3PNRuXigvMyMnEOg4M+E9dzuYqfW7e4L7u8CM3zser7RJHj3+ai2MHBHaot
u8eAPr1+TeqbSYkBuW+AdXzE9uJUBCKZbQSD1GwKxXC04xf86Gw8YSL8tsGXk9BATjiZw3Qgi6HG
EojpnY8n6X36g03YcFyi1Mijx0W8p3nY2CZJ5ZtNeRYumusNFmD7w8z1hbRlUVfH4KLJ8edBxMZ/
hXkvs0IAX3fqS1WY/auZF2OhwM0u/a7j+bIzwXu2MAcYHgJDMZqFVc4lHAjkeufLmHqOST2ySGcz
44JceDcq31vMDJ8JGc71xJkBGbn08KvRabNZif9sd0w79Fs7mTRojwZXR+XrvZKRnlv0PozuZ7ky
pbc6KUJhdUNcU+M+CCcL1gt8e2R5AC26ySv+5lTO2M/kZaWNrAWO3yYtfDtbjwRxQcPU77fJ86+E
RHZYE2/azAXnrTfSLUSnwV6jSg/VjhqImjBeYmcOhuO3I5Imdws6T+NzvPASVz5xc5CV6pip+HRR
d72M5CaMeHL4CTXcKgWJj5ykVLZV9LXoQxiSKWKXju0tUZf0j8mHga5AqbxHTgSDmfm8Y6GJFt8/
SlyN7/AZbjMKVGz60bR7VqopL/B4QFfAWiV66jr2MBIYiLuHP2tbPhy23Ua+iLMhSegNybbkRpFK
ZNVwa/8osb0amsAKhBJoi/ro1xA1K6XazyL9o7hkL4i/zQIJ8io6zYXzFGY7VsMbPVJ4xxaHMIoy
4wgJPCzFmEmiVm1a1rWsC/pticGJaLObXrnz1e++9YRLkLkfWCPB+QbRjNgPAyQR0kkBwecZj/hI
HO8YOcYHfHpb2TvwWqnPqXoGZY3e/ayj+77zVY86qfiyDmotnRWtt6jeknjq7smjuQ15FJwjx4HI
1OBijAyIer5ZlQV+GpixMaSuEqJJgXg6Hlb9C2b2nure6Ls/wt8uH8DYf+DLmI0r0rg2RH2UBUfm
hzEtXLhfFXWmEFurm1zf8FcRIxaZIHlyCj5NccK5f1OOTXZ6fMAtrojYl+t6U/C7LKCzEhntslMS
Fmhg/Ehdf2R5vZTLT83SfaU0/w2rzbb9WPPqkTQOH9vXPJQ2uY6rfqxHKQuFLhlnHOZmkEXNhNAH
wMr5CTZ7hIVAXvAr2dhKh0Ru2/1mT+6rqLyT4ud3nleuBjhEXbP9vgGjDDABOYALDoWoU05qYWJK
FJMEU1+rfQ7SmvnuSWEcTp/9nwhVTruSzzRpZQgVWgrSPPbLFGSUYzZwjhsdDL3CI59UMXoyXKgZ
X5XX+CdG2Rib0J4qQuyCemaMr4O5N8in3eJ3dxGZJ8ptK8gih1dOH9x3OADi5NuP+BIhaApJOD9g
c5cRhOX59AkZXE+/IO+IFzvPxyvuWhdQWo8xFHjX3DerrShQVJUibH529q+Zveco61oTCbIp9r1L
dKBY4xiWTd/TbiWO5BOiw/lSvDBkWNpTe4HQxKF8T8pdtaafL9ECa6BjGDYQRb4v3dNPUiiuIt4e
vdQKnDv9uXBWhrd2vd0TpCcnxXQlbgm5w35I7jGte/2lv/f1h4K3feekgjQGj/TbhM8fE4zFGvyV
cPja3o3GhivqiuVwXdm9BkqwxdE8oZJZjGowPIm36O08uMQE3hk5k9GmNtNnbhDRdj0Fz492H8ff
1KYzc7MH/JmjIddgw50lls4ExPwuf5FJzFHxZG1w4/+DB81giIQV6fDb4xXOHGsT24gVIZ2LgLJr
j0R57tp6xrK4EUIf0Zir3pXiRbESk6727wI6H5O1Ye5q3UDAc/25sma+vzO8Wr39eO0T2uif9Qj4
ZFUQzbPJEI1LYH2WwBvKgNdc9vgKfyGU+EsZmFNmCMOlPVRDWVenXJejhS2mhTjmew506mlF80zq
1NtaYR2TkyDxPDTy2tm9d6Im9WmZQFvb77u0pcZ9I33reKBCsMkStqoCZzR5Tu30bA6CwTWMbAea
Iwbc8vGkRHsEeQaDbbzUXonq7G7GtUt6/qaIKENVKlxwYWlHa7p63GoQ6Yqr5+G09Cy9oGeqUUEv
qgbKOC4RHB8q/kaacSadxdDSASnI2ydgr4t6dhYW/LcxqjPajnytCkN6/hW2aF7XXNkT9QmRG5QL
q80JklXnr/aWNZciq3ZRLX+qTJ9MptllOtaAT0rkW4pV/MqRXiwaiHrflC+ozGxGdFbz6WOGZ0OG
kTb/KwjYooSe78zK+dnQiMSOPuZgEap4Uw8fSjI+sDurFUE/5s0NXaOCwT61VSApY+pn5fXy2FAJ
FuLbr5tQ5BLCgvNc12OP32eQhJJgwfdxYObLm3Nmf8ktR7fcBXIFdmOGunq48SoBefhHuJzw2dQe
PAs68OBOI9St+9zEF6ElJUyDUitlg1H5rzqOHG6MEx0KLBO/4CS/WVnGQlUW7sR7mn5RH7gt+WPh
ycALEZ/hkC2BOK6jbXNV5H4LhnoBnNUigSQeJCYU7ceyoBLE0SkSzZ+LvAJwO7lw/Nxr40K0ih0O
ZYPET6u/UrnAKAEXZvJWAmzFFk6VDwrdRegMYYRAw+qED5uwpmSRs3L0DcN6TOIwfQ8r3hv/le8O
i0yJI0dQDi29T3q+v1sE/jRASDMRviMgDblx8yy6ZQvye7yN3ZIE1R07MquN3FdUUQbBB2vIU8xi
kmMoT4OLIK1p6YA20Cwe31KK7tOVQ5I5gKAfGJa8tbgaPTnfgT+ExuGLL/ZIwOqleylR/iMjt7Dq
J/zes4W4H/fXjCKKZ7opsrKB6nIWL342Tmtnk4bkrOzy2487oXqhLKAOp5CUG36altC/t+KF6WG5
XNoIfh0z+CUn79tPLQBapWD00PV/5ZJEboQHvTzVWXb5wfq6IEs9tT7b0whEVhUgIkKd6jTAD4Bb
lky23bNaY/nklckCf6TkFShYYR6uAxH+L7XgwYB4hpHYpgeJGnsygnEIlzbdZd90h1bQHJ8ayQee
W0dIUrhT3WCwj69d2bmf2ZDkrhK9teAx1qy8wdATDHU1IRwujYeHG57Ndt8Cj64yprayDqgn7iWK
A5SW3b8XtyJ9BrarC1wtvUGMFoLhoBXPaFFkb4Nr9DQrpx1/n5yaRVhXbWpdeR1T6NvE2xS5tmE1
Qm1C729hMm+/PvEwzvYfOUdE9Oo4AYx0tXiqKLc/7L6sf0kPjWR3PYvW3PhfCIAInb8WXlmx8ouR
GbCfrNEb8IJi0CWHuM83mvqa4U4QiJ0MVmog0MEATS3fGMbDZuTr8XV4iwcMnS0VDPleaKVfVnv/
iuFgLekbvkHsVyXDs3PE6WoneTrExE2YaaHNJpZjdHyKGFh8S7tsfJXJHM0aamZiPhb5xEe2Lr/B
uP8k+OxKTtnWgT0Z9qFePwtM/eR8/NWH/5ZI5PqZQPeQgqKj2B7YkPYSqPb8xKn2tbNy/jKU5ptE
g9nocD5ywTHy70cf0VzqjUKp/RP7NnmDfMoo/Kmu2nErcRSXGBoaEU1kFrtgy4WJ4pr/6z/x9KOi
CUeFQj0uX7nmGoEYWavEnzVsEN+/ltr7T2oNBEhZzfeg8IjBnbr4hrX3CeIP+UVtt/azbc1/3qt/
fTcFmYTuTL8IYQAJd9xwfyZIviK3LZlXh8nhOCCyJEbBYr3sNDLtgIhgJtMkHIVvaCe9NaNqP5Yi
QHze/vj6KSZgDMYfqhght9VGRJNSoJB0D9EuGYGG47ycbaQj+ACRX5RtqC02EMSf21dYx1zVYwJX
4BsepDhYWMx14tJdIlnddUxFAZxnMLXWOJYj1NWYmhxjFtCNb0pFnyuYKwjpmY6RWVGSW5ghe7yv
yk74BjdAHXXb2jt5jRhNyTNy0985mJLRttac0WKBHBfnRKcnl5i8eJoh+u+VVIueQ7GqlMVpVpx7
atOIQp4xYOVSUEX4iZ8InZCc6ZbKHT4mxsZ58DpTKgaTHLTAQrly8dSC7AkSX5n9ccyso7q+JEhZ
OtTRI4USpiRifaWeFL9JjOCDWg4SxbZT46PZH5OIuSpOiJfaciBlJ8m6OBLZTfX7yh9+D5R7v10w
KqT/6Xih7NaQL+CAdSqnRoq9G4Xlc+hyKJIojjQs/sOAAVRIj8WCLMNonh670I44hLkFu5POab0i
UgFuSzvC6cBtB/eUt9Gbm3uF2r/gYgzqC+f3QmxVJOBXYUDbYVYUW4eF+VdwKSHtHlFmphQ5JXjZ
2C5UAGTOlMATXWD8v0Ct9nNEvLsWWFhrRpFAeVoPuWSDqEbBho2bbIOjt3WpHN4ix3rz4D94MGbM
jZZc7Qu2b5dHKlLEwqiTmuhGxUZh6HC69T9sw6nIJvNaPsvzFmK1U7Ip6C7KyjtAbyhbkeElplIk
m0EUNn/WxqrWk47skTnuS9K3eCO0t8nkmlK1S76AqU2HWXfAN3OOjSUaYn1vsJNATVnXEPISIN81
YwiAHZysD+bK5yZKMeCoeJGuEtF5+WDzpULDnltagDwTUB43W0MP/3d3tUkN6/fGexX+sfRusHvC
cjNVtdMM5wcAmkyi/Ju0AsPPqbk9wZ81kFX9cIdN7mKJRbm/LCVOJAwf5Iu7wnScWA8ko4JuYpvV
T7j68BbAa3Bw9s9pUUh4ZVq7cGmDB61iZ3UEnShim7JN68eQ16V0eAglySZysMFWmtNaZc+KO4AX
DXctYgfa/ChAi9q1rf/db9XSyBb0UNGZo5G5kNTD7Bf3uYu4+WfA+LZLU92nGM7wOWQPT2lpPKoe
X3dm8YGEuPsXwqgxU7W3O5L/basf+LQlzJXB2MfN7XKWAiGpQFN/30pvismIKDfgCzyyaIIWK+m0
F+C40OrMznaYcPQd+YnijaH06/s7qRd2RXwP/A8PVqXylKR2yv2SCOFMjyO4jNHp8sHILbqkD8rL
b8LGKHolPh3t3XUi77cfdUxls/VH7Vky2UHbygM5FbbkJ4tp6sHoEX3AhWxaif/rRveTwza1zlOf
hA3o/oFywPrp25quvvE6A+BYd6pYxBQp/4VZWno5OXRW/rvpn9O5NagwGpwuxijNhXEwb0yb5JhJ
VHylP6GdZI4grI5eElm/G3GgNH4MnWGWjtnsAKN5fOjE2Pp3jAsduz6fr3xKddndyg1EuMn9Zsg4
9H8avfd1syiQpe/LCAjGOL9RVIh/EGQjQdQF414HyJw9BxOQqhNRq/rcLZyk1PMqPmRuJNpSFgJ8
Cq1bgFsVUj/3kuqmxH7731EiL6Vrwvss3nh92nRCTxnap59Wi1YQ+fKU4nd4xetSDWYqq/50fz2n
pzS22iYYzrNrx0D64Fh/tlPeV9YIUrP/MC8xJNk5JXYWlEVlOlVJHnRgSTkiGealFC2GAcMBvDyQ
Sc3kIkoeaWjTisAy0SAri0pUxOOoomz3+tm/VO00cSOHGuqvu3/XdvNLLEeHbJNzxjwQndW+d0Zd
YoKOOlKzsnaJOpUh99TMdryZm7d7PP78uWrFPpokaMIHIPxPReucoQuxW8NwsJxK6FwL6cuMGG6/
eNDOsbIhWacH47pgAgBa1edGBK8Aag8LWM/bnTz10fczFLfmtYRckXUtSM2E4NP2wVwcaJw2/R9a
+AITh1xNyXAWEYINlmnqAeWTKlR/JulgGy3WhkJ53iqxokZAnpfN5Rs5CPwL3LMi2v+KoRliVG1T
M9P+J/PBVykkTIm4TlLWR0e6NTbeqVkUwcXHvDC1XZdgh0B9GaFCShAwQFLogucFwBbiNAzjicjF
2S83AuFjjPNyGajwqmHDTNXvtPTYpsuk+ZYoqHe2dE8nCxT+REwf8UTJuSvex664kNopVtNpMi9w
t+dwY2MP1p4DMv7bgOj6Ywx4kUQPzpJa8HMgaKEKlTehvFIhOrezr6j/kFO7YWQAMFLbJhzbs6Aw
XRMfY8GPWBDtXinzEMaXWtbY2/SLB+/ymgmFi8O5fTVo+BZTe/M7cgvIH917fAXIxRjbcVT6c7yZ
txsNXcM5GfEXxQTP+BMO3HVVqnwsdyEeqwqRghIWXVs/Bj06K7K12CfIimVPKi/3/8ZOga3ZleNk
EYRKgnZH4+IIwF1ODoXcoE91XrVdJtZiuRpoSHSK7FHB62HP0ZYcL2b74odhjpyn3nEAvJrSLtdW
OrL8/fu794vwNfajnA0VkhNpEqJ/E6apIiKoSD8//+lsudbvSiUdTnZU2gtQm+zHEeuFGu3Td2pH
pAyvEibdC8xgc6RFOg0rc58LX84iLepr9o3AvELe4aROHaM/i03YSmHsb6P9k2Hg24L8vIaeY24j
MlJln1/a3rjN9UXCjoVpFaWHX700m/hs/16Zh0HR2KxyxThJ73Ar73xsROd/qX0uSEnKSE7KHLKL
BtBV4hJgZUFdmd+JkSTsIlojgs+3uTVn4grExeAALXh27Ef2oxHYcNbAUyT8fKePTzhClltq4KRU
zNosmLNyEXRaSSieYRa3WFI0acbeTg/AIY6K4aPno+czb9T8GuA/6PsgZhQWCRdUTZ4+1NM+X2Ay
VKDUdsA5ds5jGtcdYOEIL8JcIRk3n563WzbR6wRIYgN8H/H3qH+Task7OY1fHkcGWN1In79EtLU4
gPLQiiYE69su85lZbYdeTT4Dv9FUnulOU7G6eM2Hdk+fdNmSTsHnSyQu3gN8GpVOsGcQCDmpF/nl
3M+acNJHNzd5Z3GmXPytL8K4+00oE3AZkfz8h5vTkgxLtONOErD4uX608yUqBNIoH1RpZxZW4N/E
T2x/0MWWCSv1GnSPti8E2tGV8T48/FCvpGrjW4EEuKZ0jIvBwzONLsn+qmWxAgg7A1gOniBQHdqd
X6tNolWZhdTV4P+f3Veak9IASHM11n1qSwziaKl22V2nGpEnA5ENIh7Xno+GjojMBGCeMalkG2l9
QQkemKyTPhvuPN7P7IPlmY4X2ik10GMndyNEJI+mS7F3ehYskTYULeRnuRMLuGUM4VwmEo9dC0At
loB9A5+RrAusS/oZvwChx2l7QSUhE162wSBo/nd1cDXVoY4vRWwW2nTD5aO2xoFC574PL4tl4aEi
YDhphWbhLauG7Fkf2OAgcEW2ZH0doGl4GYd7hohZSo1dzW00ZTxsJ2dg4aiY2o+rh3Z3ISRQYEeY
+BjbMTMl427oi3VtnW/Zrb0jvLLzFhxNspvOSh8UyhxfmIBuLoELPSCVV61GxE7WqhtXnX8wBmi+
0dIrysMUBGnPKvLz69YmzzLWr9O+ZJ/dqoCUZBBNXE2K7RUeCjEiB5XYknFL40GBQQgxxJzp1tev
DLz1N2gxMyePtNneZPneWX0AxfuDB5Ykr6sfl5T8ngsradeBsjqjpCHjNMAysVunq1S2kRujhk4b
6x+CIJdq8ugInfhJ3JbDIr4VawnF50g5r7slaNmt7FgZwRttsg/hgUVX4EoikMG826O/LeQmI3xj
5sKDGhmZ2y0FHh8whFNIcUAcb3EqUQZKd8XwT53+jbcQXkRLBqQqAMtC46MUcBeTyCQGTBHfo2uM
63V6TvIcYQqidE7nbveOj+t9N2Yd1NqGwMwAO4UGOff7j8bJ7zw0LWNNTpxH6Bm4KkK6vob0kAl0
aaOpK8uXyWd9Y+uJFE6uzIiWl4AA50xYX/KUZAULKLGr0XJ85XkcsaO0rNfrbiwTcgy+SPZ+pNN9
KYCdzUW4ZwYH09B8oWJnqalmmY9JlII2HTMt/ef6H5j7Czmd56GQ7hdykHea7soUHWPjIzxHQJ2z
u+RZkGCuLYFEwvj91DKL+sLtFwsla6rw55QiLHg7RDJ1c2ED0WW5Rewe6N963XdlyFOWl3xxZ/B+
Dxg/fBvF6otbjHOIBbjei5nr3K56CyyVgaKyhg9pbBSahFeQIWGnAOTR6oLjrm9/Xb2rH/sNs6dK
8Jjs1vFhsDSUmwpG6LGVOJnA/Lmyo7d6WG6wsfN7ANpVoHttHxhV0nOWuoQ3gq4iovLyC4HLvOkc
uzXPM1HgwXLT5NTS1xXm3VY/rvCOSvq1bLyLAjOU+MrAixPyb2Gou952vi/vys/xPSg0D2yI/i2+
w0fLkyqH0+Zq+WosLDe9Rs+nALa0c74YxOOMS2Hl6aH0+m7rnlG6Gk9zJ0oKtS71p6BiGxvVeZfZ
mnv3ugi53z5bi97lyuGRW05Dlld36lB/zXGFC0ZNt6LMEArUxax86WkXr4Ex2Jh7RLVVMzIn2ftM
eGe6J6e9hzy4gMNofHQ5IYVTBXrjK2w/iGeCSzSYS6L59PwfU+/rs5D7USoyTVanbd0E1+6jaI3j
K2SBqj7jFHK5TtWJ8mCYeoeRYaYheoqzV04Uy/GbygGewD9AyYXUi8d1hGtlcYUatihO7gyPe97O
ivxX7gxOsMkHsvAFuWnue7UwzwWByWV/dB9IOoBnlgbkwwOut/L8GGMtObMIQM/30gCm8Q6IdKQY
AfaC6D9ucZFX8My/TmEK+bqb7Js99STNIS5nl9LdeoVDozo5qOV/8DdpQgG69V8G5J0LFy0VXnhJ
7jYTdMXErCWr0i3wOyE7aBb3mYwyrLsiV17pumzW8E6h9S5MrVN6rRQ6DUIAXCGYUQY+4gYlkDWL
aEFKgIt1MEMHVUapMQHSZqlTDD8XSCGRD/WfiE7O+mCk/vrsSKfCM6UVhhNlUXQlasQ/nkyTdmVL
xx3TP266xols/6oJ6e6J+BLCZw60
`protect end_protected
