XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���6k��8�*�\�M^�O�AWԶ��w�~���������)�,8�]��:۽�[~�%]�C�_�PXP�h�UDG>����q�E��\a�A�K�H�Vʯ4�y��S��[0�5+`��k��X��@J����@���}�y+�v���іk�օ4�]W��J�2r�G���e���GJ�r���+ʼ$�jN�T�l�-nl��e���K��>ac��5�D�eC/�{���7@��h�]=�Ϗ�� )9J5̍3�I��G��ȫ$����835����W���=t��\�ay_�]����������Vxp�����G#rP�#���T㒓�dvn�����PZ�9�lս"
M��cs�c����ppS7�D<��r���݀�6xI�	}���x��c�zƛjPB҄f
	�(X2�/���^׮ٌ`���$�!0�������l+� @��{A���y�_Iʙ�+a�BV:�B,����+����Wt��������m�9��p�J�ZP#_����^�4n��x��HS��` �m@E ������"�~=xWw�\Bw���EnN75@d8f��,z�v�1���)��-�r��ƢX
4�n���9m��UjWC��x�o� ͂i�eO��}�Q?/�S@n��i��T��Y��?"L�-�.�)�03�:Jm���裖S���~^2�G������7Ro�]�_�,�d�jD�YIf&���w�W�r� #䧣p8�j/O���Ӊ=�>Q�dg���|XlxVHYEB     400     230�Xt�њM�o�6b��J�Eu��>I:��Ц�-h��@V�(�iRr&�
�0e����l��0�]�����W-��k��ʰ3
���^gR�\$0��� ��#^c�����|<�]�3!�a�g��m	T���`����w ��ߐ"�y�U$�re��)!�ol���*?z�k��ʂ;5p�{��������:0�L�0"��3�܍�{X�N*�B��wA=�p����+:�ז,���r�Z�?�{�n»'&V��żG^��3���瘿�����ם�hK�y�|�i=w gG�n���"�w����l?-����H��ޥluZ��FrgcQԀ�U@��M(�l3�j��R^�,�Ʀ���.W-C޲�&q5���LcOe]-ƅ�l�t�=����=W��	�Ec%iw$�9�O��
2i=����[�w|�ʸ�{XGN}�h2�;>H? �h	TWq��(�<(��v4�nۙ�_вܰ�o
cئJ�Ԯ&�G��D�Z�N�ˏ|�i/�?�)����#D���O�E.�i��L�۳����ZS>��C���#�>��()�qXڍXlxVHYEB     400     1f0��@:+M�iBIQv׉
�YIw̜�(�@�>?sI����=N*fa�!�ٻb� M����w�[�2��.�H���۹�}7����62�0SX��ɟ �Eysl��Z;�p:o�Ӑ���Y�ґ���
�+��{)�Jϋ��Ɖ�RR�,	�b���7C�jF?��*� Kt��v��G���L q�2�l:�<��;S�`c�+�����HN�ON��a��j�����m��A�|��&BT�#l!=�ܪ�)���]�&s C0b )#�����oU������qL�C��e�����������Q��)ϖ����<�8�7+ߙ��R��:#�}����P�����˖�����,�(���!��&0���йI�L5%�0��·���?�ji׋k�IA��gɛ�P$�"��k�v��J�u?��y�����oΜ��{]�������Nw�\0ڪ�o�E�߉F\7h��s��;��6;Qgq\j��PXlxVHYEB     400     1b0�Ԇk��L��!��A�O�����F/��'L����Yd{t�+�Z���Υ�m	��ގ�oJK�_�1v]���(ۢ	Q��<<�e����u
�'�����,���F��\�,C�?n��^�x�Px��ɛ-�zI��R7����5� mʪ*w?u]��G� ��%�}9���.oD�Q�Lp�!@3��&0vIAl���T�EMc��qW��B\�2n˰�PV͋q �����ɵ���xj_)��ǭ:ຯm�Q���X� @�")�-S%y#�dkU=��EO��#�-�H�)��j������H�Dc9!B��#�����kL����ZFHU��"�ƻ��y:.z-���qf�Ҍ7���l�|�V�Ӹ�n
!�>�2Y�jG�}��,Te0f%t�"āD��BA�*��*�Y>4.�XlxVHYEB     186      b0��	&��};{9������R�sP��x�o��R�"0mq.�u�/�=�!2k7Ғ%��a�4,�|A�of]y�)��|7�)%�ʬ5�x���`�����]W�Y�m��g(7 �F�h!/}a��lZ��Y_���s^�6K��E��5�꼧t�	������v�O���Z ��f֞�"�R