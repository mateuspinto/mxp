`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
Vwg+qnodk4fUtB+VGnvOJo5uIGitKMzpr5Xkxxw2K1nUnSIjaHpIxuDtsJC22LuLEttuakgXlKOe
NF72iC13VRJtzger1MaKNuBwAwvm94/xRV91PsoB8mwnkMOcM/LPeM6S01knpJP3phY7cMs/13e+
EBXIC2MPe6yRCUdIMdTqnE1/ZioTG5YJNeCP8Zkf25vKZdvaAT4vs582oYO5WRS5Akrw4mQQZMW6
F2BBwluCUyWydSg57hW8Uqnr5bQDnZxbZrfajw7i5Y0SCPbHCwWRj7m2O5VR1F4iDim+rx5gWF3t
+dx+2G0eQF1swVE0FQJf4MxFvUBXd26YPOKwjg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="1GwMFSGudkHOlkfFCVYNL0H4/aKn5j/0mRm1hHjR8nw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11984)
`protect data_block
tGaPM1EA67dm0y3IyRjpo6Q33C/TYlJMfmVSoC18aybxb7Qcuv6iCnMGCK42NegV9IHPjrA8qpKc
diGbQGTeKiAVbsg0vvrC/cnaCboKLdJLyNkBl3W8MLrMKf3ptbmyoomGwmaekrcVRzRfh/tkkYg1
lh6BTCTRdY8AXtCYW2wGB01c3VNLm7NleC8vxH5qBf4wTFg1oWj6v9n/4y0cTJd71vnCIQTvndPZ
+6lpS7w4Ne/ILJY18GoxjpU6tKkrBrAzx8uLz1asdL8pNeVKrai8/MpvcI0WLCboi/D7o0dfLT5J
Ep157sLydGLeqwtCAuQa8fqL7dvz/h7ddQSe2w5uMEr9i5FsuhW5yEVR1HtTqsjin7JMP+QLyx5A
8V8MUNsvek9TCxDpflvz9sH0BRR7HNp+3bAgAbs5JD7zkGvGN673oJtqwGMqSq7BEPFwGrVxxJM7
aYK8Ve/sJpkaXxfHPAeZZ6jtm8FuJKfl3D5AsCxIOkbCzJ6Fv/alAnk1FZZ3BlHyT9pdAm4erxNa
26fz5z95zoXND6kcatiZpn25E1mHQdW7rE4cW6bCMsQmpoSf9RkzU101UEYbLiEwIvdNMzY17D9I
NhaX02v16+xK4ou6JEVFkZzrr2Vn07FAPNvXIm8m8ZEeCdY6jLLBTTXNCk3VvQ6HhLXUcrETB90r
0HTXdWYj8aQpvMiP8pJ3fe51N0zW/kV0ShNv47vbtf8O/OAkWrxE/behzLWxn+1x8wzbCh6Ovbcv
ZFKI3Ft8hODtUN9mDVZuKQiJOuKjAkTrV/zWoNIiKWUTMGIetLIr8i2t2EpomTn7IX4TwnVPKVtH
vE+P1UPEOvmWM+OcaooZ7a5Xkism0lLPOOmccIrpO/zoQS8GKp1tE8loKljOwmfhlTUwBgGm+Ybc
giglElLWro+mYjq5TSX3JDP4oaeNnsPqyW8NS8bzy5w7qTRrMuuqICXJW1x81fSef0KGopvC54cz
j1jLKEtoxhPzjJWHmWtxZyJXoSw/S5vP+tOQhkhGYUQCfnhsIXCIexT6U7r43w5aAk0jsHZC5Ic0
tRo/93wefI03gz2JyCcCMx5oCf09JFwjIIhJ0k8msO0Y0ePtC5jrUndSQ1LnTZxFWGPYW05vH8Gn
bj9x6m68u1mrY0evm9HtzvJxwwhiz4cQvmDuyFlWpd/9/qwVfkjzURsiFTx/ab4dhlTs7/bpMefT
c4UlvXjF8pdJynF03z107xyYoMQxBa4ZQNtZoTal5jVxfL+xLV4GsZ9y6jsDnCSVElE0rudNgt4j
ElS2p+dZDcgFpYOUy3P+IRD6O4jEBfb75KkcgK9nRT8YaGXyKggl1kWSsykSgi254/tZUiBJ8Q1S
Kz/CsMPJ6azbo3zYwFYRhP7dOu2la/eAWMT5BwY/LgrqgNkwGKMJqE5f1jxK4j8Bct5RvFg7LMTE
RsTigN1ObYvgG8iPUrZuqiYLCZ8jFy2CXJcvaCmEBmz/a3kALzooxWR0bUVIu/WiCoWKQ/a3KfEv
hWrbFNI3s5ZVWVUeGUvimmLT9D02vwLO+sDeYxOwHTxOQK/hs9/URudNjCt8ftJEYVwZO4G1a/ZW
mSVJywEum2EqY5Ad5jkY3Xf7FYrtakjlAgP0a6y5fr2PQuFUBCT//iVc4Xm9DncDUDEqEXedCxbV
8bLSVWlOzeZAMz5OuhcFEfMRgTEjm4RI0RGVKbyZiBuWnO6KLbLk2DELdLPwyngrM1S4568Y7uHD
mAKz3fyEyRwT46JP3f5LG889dajJLQI25J+/dozn7WwaTP+gjJzuk94o4Sfh3b1V7gWmifovqYEg
DQlbpcX+G4QyZ8Yf8oz8pXMCC35dQHKP+UmE/E1F8x+HOZi8j3kCvt4quT5iwbUDTx+HhqoqiU6+
kQBsdc7O8AOYe3hqW22bDzF29h59KDvS7DLRUmE0w9rLWopKRmPzghcy6WywEVFAV/Nmq8Q9rVmd
yMuaVYncJHr+SzN3tFAUSvvRn5N/i0ZvnO2s5KUTKhu0BwU5XUxrS0hrd93JXMolY579MgFQHrA0
I/FRbVReC0Zi2vCvTcOu1Ri3caf3bbphB+Oa7mKcnaOXApTHve+VLqwc7LhlguG7LG7mhWEU4O9D
3oLi9d34THZFnztAo7fTWiQ/GJBcuy52eJvCfozZjwM/8/EGvvZE440RokUYVOGVWwCi8yOyONH0
cOs1QchYbMmSE1Ko7ZfaPQ4+VRFtDG/thud1vtph80ECxBQ8Cn8KFfqfi4o+p3RBY+5NT0EWsl+k
fWklwOqJY3/DOnGPRIsEOFkOf88REz6Ben8pSjWWxkEZL1JXS1azvn9+IBgonPAmNsRosrxFU1Sm
6anzrDBHzop1YVbeNb/CM4/8z4iMhG0AmbkXD4oRWJZ7DeQjFqYwx2EJCDCH8AFvQ9iYv5BZk1Yk
p6hGKCL5rLZ4nofZacKBJldavciW+NpDUHy/UX+ZFX3gEkn7/HhYmg7T2Y1r4bJ/GEJnufmzS+Er
wXysjoFTswpk5VKBbe4vtkTJ+VFvfwoCBfbUfzRTGihaJ9TICaBMpJQhqQDqkNOPQsZ6t1GAUne8
vfHjcdTnjaOy90i41c4X9YWx5h+jWsXvso0dFomHbTECUH4MOOQK2NjKlcuUWv0BdJJW2ewlAZc5
6p9FNb2hwNRzKBaXoaS81gB9qXZnXlPH5s4FY8455sMZ6Qn9xPDbRfxR3so0ZU5Iu9l81DzzbYpV
b2S4lnbMchlfB8V1Q4KhoPpp6AlvMKFP67MIGvKzTGb0/+FEkV38ZyBE7fXAjqRb0OIQYKaEnlxU
ObJ10PRQxlsk8HeEEKrL0M8UV7ucnysKyGkJqkhWcFOQnIiiMJlEAdESxk6mwh8F5eMzx03OYORL
ZCpLw+KgNeQLkR2hiI1B+u9wF9JMCo6ZAuUePDE5oHZOU/GMwXlRLQAcYxLkA0dzsRI4h5yasBtJ
OJGFISHmHMLsTWiUFrEOQB3nCt1+8oPw03Uhnz9GDm8eSt+DBxPWd1Da5REuxJZsDEfUUgoH6ba7
GQSYrc7MjFuOdTBnUejAWeipjkj49bRsI/ajqJs1qs7xLLn3RklgUzcBASgyndYhOov8N7+uEg+3
9/TojJ7GientRvDWPQy4yj4NoJqn1X5tZZcfOa7tExgntU1sHWQnB3RG2N7u97WuXzv9axXAmfvG
6yL+34mfbtGDaKFTlFpa+wNY9TEuWPx54MOJMRNgvV40rcadPQRGDEnHoUQfU1a521booDV1iyhd
Kdk9qOXW+L4yoXcR2dg7f0k7YePMUZJmKeeOv+h9U+ZgkKNyb3j2F88ksq5wOZNvV84zAxO5+4er
VdvGnXFoaKszttSpi+ldQnLdIEaiWfxhfBzZn2Z9wNIOb4UG/IYEb2on8cHPr43pVO00YkP32Yb4
int9nevclW061A3Cs9oixljWXzYT/xHS+Ix9b8XUonFgkdklsTX6AcahpLthGPJFSWg8OpgltND3
G/C5aHY8HllkSYSBdFlqh0zJE5cPhYgf+ChDi+DqtK/D2m7FUJmZsQvD3sFiAJ4UAVQkPXYNrE2N
QrQ1kRrpIQA9egxstNDLoviy/74YxiGEl00htnbWpiA/N+lMqpMFMJW8OzvLOdzM/wzCsATu+7vL
h2FMGONAFxw8IPDVcCg00QXIzmTSSkEX0dVUbL0+ubbBnZyovoIlcGddet0UebF3bcSWFnYl0esa
osA+i9t2CN4OqLzJfC9uPxbPGs80Gzf62ZbIIIsdzlznpgWg+8/omh9a+Mjex4legBVY/ab1xiXp
Nj1MmeMbdDlJQ4CJ7eDi+wUawL6hj0ulRAFkTuNrq1pyNb7pOk4k+7T0ARHsEUuKsvGvYKEyFDkU
/zFfgaK21ScNPpGhnaVpQ6dqCssl3poOAf4UpiQoIPTzaUexQRPWua43JPjEuATH0H41bCdIOPm1
d7AVDdXbgE/cQ7x5MAjIWoARJHEXvUHgZM6mwT8GNb6/jBWrR8Qis0ZawhiIs8SLbcX42y0LVIGK
mvjmK1ZB7c3G+HsXlWZLzHYR0+TuVllYyKIu3OxvUlUJHd1rBsvIIO/8InT57y/UmQG29w8xHVyw
6rjh57x0rDNlnv9/4C+SXdDRYW/RXb6e9K8xSctRgTAwnGI7qeJaoVkqWV1eJzT3qkMbBZj58sQX
VZnp20nsJYyvtjAmrUAY2KnlmU6BcK1xDF5f5aKYG92v8ZhEOH2OdUuRH5MqQGOuMrMgT2FZ7yXq
nru+Sz6N18BRLN9KI5NMpV/LwImq18sVEIOEunpnnXpex1TZPg1ZHuWr2u8IWvAhimx90BAittFR
j11DvfCDJcdvdfcxaGcLOpuf8xRH+SKzJNYAtLcSxf2de+uRA7Ay+c11lES89Hx1uyI4Q69iSQN3
zufUghTLiCQfcjFgVupGhvEdNcw9KAxf0Oey7U5X7AZ8aUuorwr8ctNnl/S+If6xSMrImyOjwdS3
7QwxR5bZs69XmdXXXwzhyme7k+mXYJUF4MZhqpxN6H9VVRlKgJ/dNE1+fG0/vrJB3uq0F9lr5F4+
4Ok87iPjKdt5ggpRbQLlrsoXqNe4KiQg2Pkf0IP9h8HXNvoEMVu9ieXybn1/Xro0ddajOypm/2pI
+WzQwcCaxtCKvQHwVMbjSeDftKrkuLOOjvid5d76BLw5PaoY+pYhWrWAnEbsPQNGMi+B1UhXsqRX
RJtdnTj+Ed9agObrs6OD8mrllFK2LZxPhkQ3tVJ3tjtXXBMn46NOg+q7DzxaEwSSjM2zc4lUw+J2
9bL11EFi9t1My7/eyORJYVFuK5mok6LmepMpltdzTUrXMcjzZRjjvwPH2AtCTzn1SCizb7GqIKqd
MyB3/15gfLNheireIJ+Snu+6myS+V0HAXdsEu5CVCGraJL7MeqnY9mGqGwPEP8OXwkqN/ISzDKp0
ymzGMfr2RHv+OdewQHU1QSJo5A0mFYIm1aONtOl8PZeVub7TG9BuNCDTAVYsum0s0xx1vrPuFp4O
5bJjo/wzd2LRTuZkUtXqBr7osmBc+532quZF93duJW54PPDFBzul3hxd4QON0Fexg685A1cz4Jl7
n3tIoWWdMwD9KYVd2AetKeWh0CO1j3MbQOBL5xoPtAVTooJn8GdbkRvgmtk0WkMRH0vCw3ko4x/d
BbKY2JBnWAAIZwFfdCMpMNf+mlG8Lkl4uwgzeWQN3LNKEesK5esH/KBlrvia5cZsfztFIBlZPxJA
Y54QHqH8T5Y2J5KfV4STxPQ1vvaDXbnZGMQts8PdIwfDn7368bkKpb8Lq2LY8WpsXKIYjKl/xTHE
R0TRh45+C4Y+YuTGnUCUnZOwVgpzDlPxF4rxfqqhTe7DLHv1yob4DLjILgyGDOMa/yH+5DlQ4Nxd
hWeQgObRMh3fpU0NHKEz1BIY2mHeb5PSBiVT9Q1VWMgTvXAjZylbilaS1i/rbWpqGwkU+2wWp79V
SeAgPN3j3wmKHygm+FZhft6mzQ55rIW+ymEtG+m2k3tDcvqMCEWuK8URl80eRqTTr9TpJqZkqr+A
Uf0hSwTQEd3/3+lays7luVteKwiDhuKL2YXBLem7mKPNeXvegeA13R4PjGr6NH9rkRwoSivIHemA
5+y4ykUXp6hY9WTNaXK7qO4h6GdrUQvcoztzZmTQKMr7+SYv8s0Dae+j/AultvrenPpxBzKjTChL
M5Kg1k7eF34O57w535Dzl25h4BCJYEPKaZ/RvBdNnRqpHe0yOEr99chhp4cbgj81H/Ybc1BOTDg7
Hdg1fY/p5LumkQMQm2sKOvvCrD63fZS1oOA8NJqIbRYVvAJ5lndpC6m+l/Z70trNITnFysUcgIdL
I2MdUSYkH0H8WntCCl1EF78DYvd+7KClVrHW9HiMuLO0YMNJI59BcmcGat2d0lRoalE+PrfM/tej
Hj2671mevQfgdGlv71l4UE9aJurdvvAUqb/LEC4YCNY2GANKjXaaembaIdr4dzkbL4xxQV46EThc
0kMR9EdV3lBbwel4Rqv9RbilGGsCEhhDji7xVsO4hE2sNUzKkoMc2brR6wH/Ee89rJ2ShIU9fkhF
QfhQGh5QregWC05wkpI3yEOyHJtUCYX+vqe2hAKkHSOz9m/HDHFmvj5m3e8Q/25fk6x1p92z1vEn
HiWtof79S7Ih5Ilp56OC7BpgDm0AR9iS4VR6UUsYoU1l3SzpjAVlBzke0mfLWUEE8xLQ8rzWQSDX
FiKnVDyNJrger53xPlhEpsTgRX7n9UGq7B6rUrt7ZPdjH3MeuLJg0Og0PmWRb+zBXpeCtyRLgjT+
wCNV0n7YMGRVk7gJPf+bEHPxcDao7LYbZ859mz8d3d5GI5Kt/jGgwtt40U1RWYe3iMfkOOBanDND
ixmrbffA6JorxfDKPG9SY436ksp4BxGe8/nB6HitngoAhbb1DybId7ul4bDf6d5+9wAWwwVNVP2l
v8YpazV4FL2ZxgkLre+bVSpAqp9T0Is5vDys2U0d6XNpC8XX212UuYfuSaPBhAnQJRrzqKbaIkJb
8MrbsJpIkwV++RGW4pIJNPB6/YNZSdP4wEWfXv7AWxOPrgZUSGJetNF6vVZtYwJaLfOVMlsKZ9dj
IM4MUwF7uiTfJLW5eanR00AuZcywCL42xXfXQ2W12K0EpKEBSjOUnqS1dm4OW8c1lxAEaZ17xqJk
c3zmvHbV4I6krr9xY1rZGnK9CgLQVeTBMDz1PYqfhqhVk5bSsPgt8Sk7IJJycL3vX+iCDeJaA0ps
Ob6JBzZuuAUcNtIuRmaMrjnE5dQKGGeno9VRaJwZCpSScZDvZ54kzAnJPCQm4sxE2P9J6XJTF47L
pY5y/26fUoaBCUnGJ84m6DFTAcAtysnQhtvU/WjPiL65QMjIwKOGzPuiY0U7BSoUkaEqWTETRmrX
qbn7LJ8QT1IbmJYWuRb94+oaH2mMPrVGB5SR8vM/MSWoJML50LZ68C7WQPbMtMzCpsf+/CXKOJAG
2ZKf8x1cgSO/Aziov8LSVswXZQ/25cIbPKmb7n9Vuisqb7dpxlgmQJUKeab7oU9GgSiFhXOY+YlC
EsuoEbLHoyd9mEb5yKvYjrk4gVo6m6w9IC/16hnC0QtdGzcv207O+VksdVfRDekiqzRFFVmJh7Y6
4UvZ3BCtUKuP5bOdaqH+vk2SpSK+r+1apbWnPQ4RUaAfqtXq6d+qFv8R1hDCmbfDv6AxLtPVSMeh
ExPP2zeGaMhKTa+lEwflV6DLCkEvQeCY/a4bmudpS28D/wfyYZMAugRbxKBsyTO6zoAdLUTwyPnl
NOH+fagHwtN1x1jfZoLnmCsRmnH4r8YR6513hanpM/cG2yWz71lzpfpBM0ydL39xkOcPuOWgWk2Y
c5+pIrqhke2kCopzkFCTFP14mSj6vBQPvXijw5V7Z8Osjupl16cTNAyJLgVfKkie+TkcHGzYIEXV
mNWO/NtQgZ9DS8dR/vrMEVO7Ea8DHNB9qhF0i408bGoTEdYQAdsqAwHcNyD44k/Mc5pZ2a8PRUgx
xd9DuXDzlF31EQXJxrtWIpzGGOMfzkvMXowMyx7LSNiazgMpjnZeZTM5Nhu4P9E2Rn0JoawCC4fz
53MXLAo8+WRsnOd38qtYSIaJ1yAxE2NL+h2RjV9RBy85Krh5iUo/3dbDn/KlqPQibC5Jc7nve3U5
rL2cm+hfkOTIWrldQtQtQhZdTXfyx2zDbNovAZUJGe+YxPQeXYcKnsxn33tfWimAVdWYK5WvJizW
7WwQL/JgVN/SyRu4aqoIA9iVCEzaTBBkm4Kb3ovxdMCSxhO/H7rgVRqxc4JfpzAny/2U77exMpCA
9TiJXmWnFoqoF+92gewcDEQX7hYXb2GQLpCPkzsRXFxdSAZLMnCTKepfdbUbozODkOefJurTR9wD
AfxA4UVyM3bOh/Sx3ODhFyfYHy8hmNFkqWIUNzaoKAg0aqSUuOBx7f/exsj+pCnTzrFQjlzAXTCl
/3xQdOcEH6e1xZvoV07q199QqyExfiqVN0QBgqCylzx6LOQOcSaWAQcqoU/xfoBq67sGzmvPpVWT
QhnIrPTMTsF6Dk23K0bIa0HNaElFfspwg5MADYZ5rqZY2VhxUAilDvzDOaHV/vsdLXiI+XWbfzhU
P/9buQOhJJBOwdFYc+TEMJ4RI8+jZZqGURRxzYanahI82DEE5AeKd+FoaBxrgEC0d2nHUtI9jZt9
tbZDgFwsxi9MRiznDR7BORgPr9zyiWgzWUbA3VQeyZz/FXj//FCt8zPdatfpT/qr9Bj4fmPQqCVr
Y+3e3oCzuvCbF7lsljSwAkHX8pIg+UH2yomD0qoQChLSx3rUwneMMEhiMD9QRBNu4HSDAt1+UmxO
OybN8w6PlgAv0yGEHhFmZyq5iR6JABMQgukhC/ttitXj7Weg3h08pMjD3g4JvcRL3WnLRbArLtM7
T9KXfNMqARRehb6jLEZ4yshSEiyk2xa2tKvHf/cIO6ddAUpXcQ+UUvETt6cmJu0DuLYoo9h8jXbT
igcxyl73zbNbP4ZWmUzBZVshFfiEcIFCLsRM9QurVXMGKdtLSrakPh5jL2z33mHcRYmvsh5j/YTC
tRAbjDQGvfuWBGS6SCQ2P/TWZs5elNWrOWbYahBDWBfsU32luSNL3KEGte+qcNE88RcX/rbWj2mZ
VCx1BSJ05rIyYHG7uK4ml8W417jReK2z4sV7TLRCIvHZIYxLSOSPEwFateaCzi1T8i/nmziZBFyB
4QvzKXDBhRpknzHJQdiune/YsF8Rv1IjuwCnVfh0eKyIzYpW+gTlAVnqACj8Wn3s3hFo/h7AZ6Xm
vhVncc0/KJGLyT9yM7Ssbx9+AIiAtMIX3lXv8GWUAMbZMHNPlyX9fOTdpXb/L1J9iaaIC44xOGkp
PZ01wNXc8f6AJomji//6A6GF415TuyPLXcFIW+BR6dLYP8IBqmIxeRIp/HrxdfrteaysuuPrgTWJ
Gw4iXgLQr6TS54RwiVE6EMVyOWLhSTOCkuSHTATlGt1Qnzi3eF9lW2FP4eqhtcQrh49yiTxIKMr9
RHiZNnOC01F7EAIZXdRjiHZNaPq0DoSBeFwbGEM3hSySHsvft/no3Qi2/LCHKGqe7gVKeovjdmwQ
DCt5VH6ubmb7NWLGZ6ZYuyFDwejqb/snxxZRCT2ZaopmgmvTSboChzBlO4jztkjsT6xVNbOEV28P
CwIuwBihQz+FtGSoo9kmdshgVmyu2rZZUSBy4YrLxH4MyLGqePr0cLH8FZFEPZ/eVTNMpKM5MAFH
S+euDpmm0ycM3NkQxZuqc+RnlE2n7wBaP8wlPU/kvb/a66IezC31KBrmbQGKmtkrgp3dBMVAD11Q
AmTY8bRIIz2aZ5ywquG66fTbpdvSbzIxD6Yx0Hz00cQJUIl7hthIAw6R9ggb/cH3rqpprhktGAFG
d/tYKqiLxOGmwUs//HCf0jOffHdXmhek12flT1kvssWyTLBD9kkcmxcXanv56+rFzmvEuEbtzO1h
+PGCyYV0XDcas0a0E8C19rFpOH5h1hon9WORoqxWSUt3CT4j2Qbrmb2HMafCbynxUFWcqqlMOe6M
niC/ahKhUP46d+Gzx1VD5mJbXEQucEYl3ZuFK7OYGqqoYe0z1cd6p/UOoTE/dYDiPbV7HOy+nW/P
a4M0T4m4YPWDf2U++eoEMngmXbEni5vbjA/jhInezFE2LIXvuiJMnkElBBlCVCUfBTnXsd3CW5d8
GghpzanEWWl3RsipBqguATZhJJikPmHhH9t5o5Tu2TisiRYjVtocsPV3gGH7vWpN2I8Ii6HAOg0e
SPE3NazFpi7PsJPETpdwAttTtBLSBX2NFNIL12IDmXRaSqiPAZYynvflijs6CwjVfQD326esfmgA
8HO/XBQ3x+JzHjtm//WYHKT8bZF8AHmJvmJkHGcrr0DXSGdMFhZOZRzO3x+tNMqLpHhxqbz/s9jw
rVw1p1N+GnO+5WfekXVi+L4+SqiGY3Xil1H/JKWBWjAY2Vp29+juJLWCJkw89wYAGGEinaR5TVaU
7r1Y85hyiWnPGrLrzMZH6ihwBq/YcXknlbu41pTuh7Tbou0JPFqiPQmUKygzVVGUJuiweHKAsOWt
dZPFWkyJ0DiAtfDryEDUoCUJRkMa7KDvu7WpsfbolYp28BxJj6Gw+9B+DsX0ZMpoxNuawcBkFBol
bu/TiNZ7ykCwrxZtIPwBMDbZuldXoco1lE6BvfUuscKTDNsRr16La6tDzpayfx5XKowJwasliv/d
eqvsWz1U2G+Qp7b/329gp+MBJasXNSX3YVb7rLnBRzlQSgaccED7p1lDt5ImVyRWr706QOdDtAvW
GKSIKzus7xGI/SKlEDzifFh7o3bsA15TPaiayGTblys97Rd8/MKZh6/AI0b59S9wAK/ptmuSagx/
Ek6KiZB7iW0zmSYaIJ5QIlyd+a0/QDBu8DXqH+loH1PYAkyF7y9DMs6SbTSPpT7UYKQyxu6UN0mg
IGhbzTu9aEsctZyXynHTd0CfvrG5sYTQoQvUYc+s4rPrsgUqzgMG99gqFZlJ/PXeWAIqcM5RxL/q
OWuEAMSMtwY//PVbZK64L5KWVVTh1Wvtk/mEyZ+ADJesq54QW/1NRF3hj1hDeN4gdWhu0LgKITje
SOn9n5PbvkWGSQnt8qmnXCB+//rSVqo3QkZ9ZIpkc8V3BeZ4FR1CNKM4TN6d8IoLBKSK53r1MBr6
zRmlYyLZYCw55OYfsbl7+Ks1FH7eK/sfCYjzulM4nwqsbkvJloYoNVu11HE/9odrThMjZZqFheAV
5pZBlUalSZE+pg8kvSEK9F5p3axsE4Xg+crBHiRCTnFpdAqTXHVq14wyGE1UNtgAhXatsk+eF7u/
LAhMX6yocHDp4rua1akyn7HfqKpFwIHmeRw1oLlFbnLnbzLyU3S9SCx3lVaQjhcWjzim38rDZ+FD
/gKdk6FSr4aDe4UDyay0o0x05T8GHY0Kbs6aVNlRpBUvL82yHf9Q5krlAYIMcNLOfSHhe+xBcghY
q9hIWPAXnpz3+QyzjrhUukOU8BPiQfS8Ws/X9G50aWXq4205qXyub/Ahe4nMpZnuUy2TVRP669mD
A+PTWeg7/Eyce7AQxSOM50dbl6LsvXurB9+Uj70v1IdnEUXvn7igC4yQRidNf/Ar0XEOrzg1oCqr
SrB/KIYQ5r5i+XhjCtR8gY3+eZeU6ffmCFXTjAQoNMnuagG3G8E+B7wG17rib5WoSW8FoG3Jq/JH
Wz+t9z/1Tl7zBSd7DnQr+7Qe1+h0suddJR/2pZBX/Gm58bxOkApTxdPjRjkjA3xADh1kQXLMGvTW
c0g8NZDcOUmHsOJGDwyFoIa1sOALJI4yr8CvWLgt9Iwu+xYBqUUzbhV2Sh4bpdjERiDpy7HFBXdH
3nCEOBVqeW+9RhWWmxaPzewHqpP+N/l2Z/yOPMmVERGk2ok2k+utVbTltUr2ZXEY0gQBARYEl9AL
oiVAKIJ2k1jDnPuwT4IwRYBIT20XmPnFmp1pwq274RdD9kUnmdwSbA/hrBVqfap9iTKkcW6C1huB
tVAhKFbb+AvPz/wpjECTTns9EgsUSH+7f1CftBH7SHifj6FNNPxntcghKv+jHxvN2rORZPoKCHKc
zGrd4gzIkorvRuizMHt9mlfTrC1zT2b7mRj5YA4CSERXcbmdkQX/WrpPAvDPXrpf4njxYrPmwjqX
35zy6vDQzhhpnKziyn5hnIatHaPycm7AChY+c9Jb9QVc6qeOFOreae5HfzIZdCvfu6xIrI6BaFeW
cDI/8Hsj46RC340EbVHhaM9Di9tUOHmofipBVS4YJ0MP5nPK2uTyqeqWoQMOJ8JOU9DJTRvtUND+
yQZkjIVaQ4Jxaf3sClXNrNYs0ZfyKO0HeHIp0yEY0AeerDzHVz6bNYJcB3YYrqVn6qEbVsZy0r+J
xdafL09iSs9fKoXZtPbIUEHWfmH4ayShQWZJSH1cXJsaFz1r96iQTUUpqBqwfXGRD519j5LstQVx
UtecGH3QNFpw0CORrywPtIqjFMQXgtd0AFVFXqjZLdHSVZ6fNntlScV6gw+hOaBm03nxkZZhcsrh
jPmlENGiHACs8eneDFiUaSnaiDE9Wa2ey83FSSyqHrB0lYafl6UKqrVT08uzHu2RO4LqG2hJDWB/
NDzNrwVgaoipwTELhT+l/Agu+JUXOsmm8MAZ25hAvHrLVwgn9ONPBx7N+MjnQh47l3FUczZH751M
gs2VI0Fen2N7N2bR6wl1fwbxjk1U9B2Vjs9mkzDwzXQ50etvIPon6Hgh97Tp9ShZ5Kk3suEtEVtz
6kfLIGhH0R2NIa6S4vBY9lUEXtSstPDm5uVwBcUa+O0dZWf5EXpuBXT5ao5DplSLKkCypOZ6MIYj
/hnriBwpdoh1rZvZTL15IERCxXmrjTewYLdyujGDR9NlFxVBPhw2qIfiqjDAc3eZgzOD06tJ2pNC
mYszRQBslycCV7Wjh2C6G9T3aBmpxMM/MXYdCqcWGKanNsa2fXQ/WGtVnImtUN512AAVOKaIUelV
xqXdnrYow87WvFtH8UyFDRArheXAYn2njzTTe+H0JWd87Zu8FQRfIVZq8xAdET0KjzLAmqLIMDb+
954RyrMhA8ai6avlmWj41Be/rgh+P4/FpUogaQCVBpO5DL2Vz/eIMEA4UaDWgMwE+FhNBLfy1RU6
syfzdb+mFEMPxvl9+5yJn5DdTISvxdmoeZl7HeIwTN1g70kDholKT8qaq0Nw9W/KnjynfBckDbnO
lESlqik0yiTv/xeyItzTUbT6n9SGwG5yJ/s/k4LcvxRrq0pehyiYB0jeIjR2fSAhY8P1n6aJ75NG
pW2NQeBKX8rtyt1iOPG8mpP4orhFvTzUXahehOCOmzCSEM9VAI0j3Lo34yjvqYQetsDv03fsY139
4i8QLXy0fY8Hpm6b3UHmtLJtGDpRzsi3A0uFjaC5k3FXbLRhexn4Fh1hggeDTDK3lEaPETdvKh3o
hkSnhuzm1IAD31gxXfVagkYawfMh/mLQGX/OG1BFqkaW+1p5dyzz47YQFRrJ/t6I9NtIzxnKVK8U
2snCcrkTl5jBfYRZm26WciFLTEcASAZzPkF144yj9pnp0jOzOHpCs2cNFWK9CNuAvkIyz/KlgWC4
GOXypkX2mSbDlmz6AxmX/VrIoE9EGZiQs+6G0Iu1isz46dJ5gocVCCEI9SiTZ1TUGjK5LilsdDab
BMXu6mf7aI1bIzfvPiQf0luh0ZQaTla9RqpeuowuRsmecxZZrh7Fa0f3k8kZnODo6npvpD5BIfvP
HJk3j8MXvuAqZwgCOQ50FwxX7UtS7OqYmJf9BAhF3Gzqxrev+5D4zWoYvi2MyT64y4u0s/iJc04i
8xHR4weJPBK1YWsiPz3W+DJnfc1XkXaPORmvNyETZBAc/8EYzVPMgrCDZkt2TnvILBXK4gz0b7KI
JapxRPINNjv1begrGq5zGQnDFmac/hoBxi1klcckOezCaUAdrkzo1VHbg7kMbtbn1T+xjQM2Au1/
hg0AWvi52yRw6Zio6xXvoHw5lQ8O8j+l11PHQpcfP4LNGxwTSqqdCGyilIeLCf7aPxutrxW7kPRy
EWW2hOxVwFEo/LD2C+p+TQtiP0jtsiWd+nRYZ7+3DB3tjqYvrNjqle8Igc8zHEYfkdIzmTOHL7PB
nrW+N3g3ttvLcmEEXIKI9aFvyI3tXeFfq1WAwv2KSKXVMV1DakHub5xtBlbQ6YGFl7bGnX00s/VB
dz0MVQ4OyRdJhe+UsXIeUYynDRSrYtopE+UukRFC3M8Hq9KXgJjHqNUpydn0TSFdV1cSxjmLXEBn
e+2EeiYKQgFgVywsj0pOD68xEbz/SM3D/3imf/Cm7rmBBCFKcZ+CyPuTpV3C/2aws/IbsZ+tidoa
Uz+orCsMmxydT0oKdFl/TEkowFI8Ir6vbQeKBnXEO+MSIcq0XRpVq4tZVZSGrzS8eKNSUnEGLCKo
fRYOPj0bzB8wZ+Wp9ZUyP9er8GIu5T7HF7SKKP8Cc9o5+LZoAEc7pCgCvLM2IrlK4fxV55r6EpNr
yUtIy/e29zbnmUjelmv2nwszBaglYJc4f7/7XTYihthwpLsDLAYV1qNswGkkTDz7xIG7Yk+JsO/r
0sLOpyNsiSxdC0ULBfunz589lZoPgd/qmFiEDhQ5/Re66ac0elOcGKyMJXcMsNW2FEaIRSNk27I0
xKegeM3LPoUATQodamKjGKguDuOKyFFuNiQb3a3cHVQT4im9w+TxQJGrTi4grAZCkwsx1hZBPgNo
LG64N4CF3iXr8b+LfWO/eJHndxiCS2LRsDQca9KAoWTdH0+xE1Gl1HV8rCmHs+5PKabQEXRjj0u3
7+s3TyG8QXhb5b5YlIx+RB8cwNHfn4Ktx/KHXkqf9xpIvYKyENvxI+SdgjRv1TptHp4Q6ic3aa2W
U5XobnuthvPDDBJa5lBJLqM5T8xggpaO63SpQjHIP8U5UzCSBThidcqBIdQgE34KVKc29wcl9Y3l
B6w/KUOWhoVggOabDEJPbwBx2lAnDK51YxfA3xuLEObPgXUN48XESdDpUqt3QNrBr6CnY3HGtBS8
iwel4LhWeolqHpxs83DLGgTK0x5t50xSt0C5yVkM0dSbN2Nhm7mhXGN0Wmc+gM3SUNfpCJtQsfqU
RzbiJovvqt0aSPcEYWyutAGT6N41Wic3+Q+7PXkOTab3f4DyiTZgwNXbb7Cax+z0lw+cCJDQ4pkE
1Ta7I7EWwf8g1MLj7RILefrZ6tYzfXLdpuD4FEHH9KMEHxxC2qzcDyKRByYqi03uffpdn9Gvl4G4
Y9cei7E+XsUT96ap6rz8oyB5xBrNK54ZSq78Q4eq14zp76N4QgaEw4hfGfdeewu1HW7bqUSAI/wj
ao86zTUqU8ShLGwXafcVo0NOy0wmGnQH6pitUBvfZOY612ZHIJQ9KKBg6CaOLn7MeQ9hedmkuDSH
dFOrQLNd1qYHBAhJsOcqBvc619pHrUF1q85QkhbECmGC6euX+fhafkek3f0qXi1icDCrnR9X/h6q
P3f91d/JBhdv9cVYQ7b87DpD0xkukwg/ep3+PSSDPTt+pg2/sHQSv2FryGOGb9J0syRLeWIj03Cc
8Nd8W2xVY4jNHxVifuKDRRIi0v4eKNo6aVca4FpOpxGHcn94rAT5TJR+nlLHjxrA9m+kqyGycXjS
yjbLo72nKOCV2PnFtF36Ce0mFP1xCUPK7xzT3m/FJEJS0yYWjpdwafhTXjFOTZnvmmqw5zI8LSE8
dR8e1y0qQ7jXXb6WTCVS2NukwHBbSSNx4W1WFFL5tXMrFv8+NAOTikfzNnDpLec5k74axnkaY6Be
xNMlaf2Pq+qtyRcyHjeCSVJVAY9dlcLFAtxS6M6Kd+P5yvEyUkO2iDk6EkVCcUtM/BimzrA3IA1a
qahBnRrYjdmDeJLmKF5akxDRYao3Lvua4IoW/SS2LC9U5h4MBXBzOOlEfMBlOv9dpo0x1pn6QLGJ
iZ9Dnfh0G6IYmurypWfFPOL6FIN1JvelYrYgWnMmqzaNfC/XMR1XN0AyhedAOoUG4WyMtIo6ZNe/
x02nKl9zm2QlLKuGMi9fKqrkH3bOXONw/tGGygux0FenMu9CWIMKDPBVXn4D2cH2aMXjSkCr6/OY
VaqFlXrZNrFpdZ/oZHgU4CLxGYp8rlR53kPMXoAkjIS4tNNu55LouGseSd49T8Cvtm7/nreVZtyn
Ky1gDDZLUba/AeOpmogVbmHPKQ0+XRZWumkJIR1VMNtKMTGZ8BaJPBvrJoaIHW8vGvzqjxV99Dsr
xAwmM777v6N2glS5i7UsNacE8TPXf/cG0t8s4nUwOJj2vGQRl7RV6gY0QcWUuOj2WlMNqR47hL1Y
RlpcwiP//iCp2FbGaRZEQarCyRqfOM3JQAMnCECpDCXo+1j5zWOAPcfmfqwobUGMxEUU6PGEnPy3
g+b+OLFNysneKJgiU/s=
`protect end_protected
