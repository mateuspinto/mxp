XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����1r�IpTit���|b?�;�������k%�.*��鈧q�V�e���� ��c f�����)eҦ�t��#�]ս�7riOW��.�|�����K�ԥx��/�R�(���l�zk�����7+�P�_[]���"k|�����J��*$��kK��7����!^H�uՖ��1M�22~�H,�W)������1����}U&|g��DP��k�9o%��5Dd��D�so,x�x,��a�������u\[������Wv�O2JRC���?��Ю��9\��Lŷń�^�T�O޲�4zO��6��8��&��82�b�w��}��u��f�{���r�A�F`f���$o��s�\p������K�fgڀ"�4�e�]
�Y��\����%���loiH-�7��\��nC�<�|˖6��=��>���Ee��`��"�L�2,w����`!r�6]�Ve�6 ����[�@���p-��BR��f9^_΄=����F���V�F29꽄�La�^*s��L�y�R�(h�t?�h�S��S>����v�F�ou+�3��>����Z��֊z�k�����dm�&�~�=;ao.�5 ��v?;�hN�ϤW�~�?7�J�JG��Nb�u��X���OR&y���s���J�N
��&l���Z,sp~[�H��l��>[�>؞�Tő���V�fO_U�����ʝz1��e�Ӛ��H��EC(� S}<��Kz6IU��kK�{XlxVHYEB     400     190}x�)�v<��p�I��{e�C����.T�/s�l�6쨰���� A.�<:h�U�7t{X�L~�/˻���\
�na��S�򋞔�Y���TG�'�J�f��"����c�l�~S�8S��-� L�J�g~���U������Th��M�U�|��_�r�b�A�XAʯ��i'��N��ϗ4x'�Y�[�`�D�aL%��lv�~3�(Q��kG"�E ��t8�h#�9=c�!p$�C�8���Q��w-5r
��WR.����sZ4KLDnN"���š�.8�9�
�5b-`��eޠ�`�pg.�gQ�˳���h�7iS
��"�BC��f`�3�r���Y�����s޹ 
�����Q5߮o�RKI���(Byʷ9���};t/��OPLF&h	*�B��#�SD0��FXlxVHYEB      3f      50��=�.�]����c�u",���L'I9CWk��k��Q���T��$p�J�qC��uڠ�>�OfX�a���&-.EHe[7