`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
aM1oM7DftyqlUAvzNs4bh+3zw0Tq/Esl2TUJCssp6IWK2WrYZqTFd/WOKHOO3ah+LiQYuVBmSiOI
bbtZ5xuiJAl7gN8C7nFHoujZkU7YERkocvlIJTtyMG6hBbnzdoz1goXA6CKTBXv/L2nsQX0g2/E0
L1b3X2KXRLvWKQe1ZOsr7cBwqmtwxX3KZxkpNkwVFGDbm5iKMWp1aPzmBCt2FkZcp31ano0fx0vT
sA0HIHs9qfP3nDx33nebD8b64v3NJxsHdOsZiXAzDGqqd3+Kvld3ZEhDMu+vG3U9KnD0qGBDdCm4
GxADoPYwKnntCgChB1+yaisHIQKqEckPf0DqVw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="0Uk8kE94DgkxHov/IUJluH6+qFT6QDX4QstY0nNFyEI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12736)
`protect data_block
8AxLewV1zK7O2znDLRU8G1dBoZebSwC7vmma7fkMD44RJLDh8WKa8CD5IUwvLGUIcRtVkGx9Zz0O
5uIgANoa2FfTzkEaG27cFze4KASswTLFhLVmxEMjJSYoaO/0x8JNFPOv9vdeUl0s0EPek4J3TMXy
O53w4D9hgEU2au2WvKo/NiVYNCO/CsSzNWF5Gn4VgAlqG5fqIyiAP6MJxvWooIMiZ+HK8Isvq6jm
JswNZP3jghL8E/H/RELZ35n2gZ0CPsBn59calzf1X10T4KTtMhx5VzfoDRmGxMJ4MJjR0UPJ+t3y
dW5XgHWDEZncrsHaCAQ4e5q6dM1MgoAuV2jiWBcCUc+ySXjZZhGrLIJkrnLTIqKWCSpycn05DYfl
mEbJyJuX7VWzO8eJAGbbmEeK1cJlDomlxTcAp7UyOZ9nA4LwzxyKBjxqgCb9rSFv2I79JAsLYcj8
vQUHakGqWzk+2Eacxs9cgPqMUgIgBHZLWIkxhpOiZ1qiDYCliPevKtA1/0YPgi6egwgSN/euXTns
4j+ynmw2ySr80Uhsb5KIm/sQ7EZLx53p+GGZg9OFcukFNe0jQD3ilzsAf4aGXfRSPViio8tdJlR1
Pbkb91hPfcvG0RL4Cn/2KeC4cAfRFW6rM46/XSw4QWlt01kjcxUPnMDbUCPndr06XzCGGoskVscm
R0TwjiB1Tnln5hok1CQ7M/9QKm6m3fQfwccf0bQkwvTpH3dP0uGYi7HN8sDpbRfUY2KztRGm6oiT
DOyn8wiEPF4RzNkhIDgp0kPhTeSfSyVq09Ap8mENcIqjvJCcNL3BWNXxkHOvDl+MykbiYWit+LuI
3pQYMLd6n2AjHVy1L7NSiJlfKaap+C4V6JgdI58MdcW/ObRN440t/ZJZxX4RTNxOOp1ssC7/pBbR
8mz441pzJmtzt1J2Bb1QQmZ3+b8gNw4PwSvAsiF662/LkT5M+oKN+QwOva0A78Urh3ffkcQcXSOs
SAV8R9gKh8CBcLInZMha+Caoirs6dnJ1s/YTYUoS/3aaQKZ3VKFiFCRIyEikdgqMuwjob0PdfWi7
jJ6LZHd9VLCoVBfJBum9ax65SX1iA1j6zUtZVu/d2Sf1qSfoO9K1PTxUN1v2c+B2EtaOB4IRYoI/
tU1UgCMDBbVGGKaQDh/Pu/94b37CdQUjfRuS/7OLI8zzCJysLn3RhvLAy4KJAVvdC3wx/fnjWltD
doEpjxe2gb/31b8Nlq0fbS25ubt1v08M6QfKYAiCCfnTbXfIGY2e1yFZfv1vmBQsMUF4kYJ/1B2q
FlpfZl7AsJW4kNSP10RSmM/K+sciQwvBkZwb0W2ar6O1Y+htK3IPhKBJjcsxSI/MFrf4kEQxu5R1
UjzPJEeQWaAbzI8i+LqXve8nfGd3hwmdKUAmYev4zLPY9YKeUfnJE7/buG5CYFG7YZS3G/M/7ZJA
/vvUYgjB4IyVBBppbQU12U3gdMnM0dQ9oqGDUjp2gDxeTEa0jxq+7jVVgvBoJ/SbLxHjahgHwNYB
zIQiHVCiX6kTMUdTb4XKNrBVs0qiwFFPPPK0lolR9cp2A+4LZt08o0/4Tt/4O32qLOFlxFbkYp1B
ispyltCGdYsOoNAX2XdTZoH72KtTWjHC389z56TKVMQvZ+AUj7dChqZe3L6wZpEfsWDrKmpnHJm0
kdsm0cCdLsYwY8w+wOKgnbxayGi7jeqTGndyKtBNukHjQvzuGazC9QkSRLCQwWvZh9W3AuUZPb5U
eMsLX+2JQcasdlHdxxGEvgiYpW802CZ4j7OK7EXmZZ/jI7dtXIT6lLjQjUW9Dv+PhLUH7zjaKAho
3oOaFOpTB853Ma2oTmK8xnQwHANJcOSm6PB7ML5FKjusfZ/xVrNQXjOQEJ/M1L7A3XSgjQVYy43Q
+gcgqGNEWkjCGF+wmtxkJr/HCmMqn5ytxijXnoQuNr8VPEn6M9k3UGt00yoE9JpGJhfDyWoGIAdS
gl000q5M6p5Nloq6AXyT/oD8iSIxGC4jkcnb3jMMdcNfN0SCSOp5tCoL1I7kTjExV3XxnDD2RIUY
qnILiNUOAOgrFbUssjJtrmHtUz3x9Zd5rWUv7TdMm8QrvbG1sQoJdPYyfBjh1YCTF8QAZ7Ef/2x3
w+wmBCDX8qPFmlj06wcfdF4DFiHprKHCNIt3nlU5xIdyXtiCtUD1AO6A/0XVER+AGutNr+XOKlZJ
bwQTjtJ67Mn0Lu9aVpg7cDfX77eSXF154xvuAcuSWokmjE6BqwL1NJVXjcPk/l8bb3F4JbJ17MIA
WudEld7F3hVQFugCItcFlqtYuIzXM5HlV0ZVUDyUIXG+8j/CW+2MFmPqdf32H7P/wiZiSbH6R1mH
lhcApHYcSEJGpjEfRbIEqmnJnVATv/33lphGLjCnYJAC5sePh5Cig7mAgzyr9ieJKKCSRx2YZxJL
JW2OOeUITT1T3NePqTzlpdfSfUgQ+DZNaakVZn23diZZY/odZLCuzwqwuUCVxMV+1TX0R/nUeo1w
NFoW0yV06opnbChhL9xRZy12nf0GqLq7p25q6bLBe0STfpcwJkCTNx0n63M1QDcpFf2bvtETNM20
IILetVAnZvhf/KHb3im5pNEXxVrBZZRhYn2nelTnAKFiwG2188YudPM1LFqBCRURNBn7mR1e9ty8
GingT9gPiNRAx2enPKghAynZ+O0TU+4iikL9QFEpTpAJm3U5kkvceFEP0twO/St2CB6k8B9KdKqj
D47TCnRJjSa7//2Lmi4n50Z8n/QdOU1tc7C9B4TcxyY239ZNaFJjgwwwyCVjbXz6nMvU5qeU7Ng4
kyMcZueDPEhhDazH732fkH0fvqRBcPmcz7oVgiHK2XPCMPuntmDtzWP8i/e5QQ0rkSMU888NtuPF
RtlUWTxVudXnTkdtCe64GGX06olm7+GQN6xzviRi2BwiV8ea1qskNoFmrWcuBqouqHJhlQ/Gjy28
dZZVWXvLhJctHraEfnV+lI1/t3Fi9gGk4mfH90o1QG+a0zI/vF3AZ99k576hU3XZOjV2OBIBN6bi
FQNGrbXORy37dcMsIuGFgEPwVm24gfglbTQkuhB+guS+7AGbdPF8k236mw2QrJUgvjM2yy5nU8YP
SnWzgLrV0NwFHeHFgj7RJo++mAnjx3D7g8jWU0HoQxPwwe8eF6CQJiQOyUHFK2dzl+HoCJv2LC+w
OVenv9KuKN3iCiNSUkXV6Hwm8UG+wHco9GFHgG/1VK3RU951T58o1qC3Tiib9xnmiXESEDXq44ng
/+jYDVyEsbpW1pkpy8cLaXYOw9V9D4DQ4Y8bb2GckvW2ebNWJIWp2HaPc1BTkr3LH8Q9F6CNk51Y
eq0/Xl3XsVnfEqtvGmBFPBH1LhtNkMS/n6OA2/RzQcvBO2naLwPoLNhNthQeNIAnPfCfwDfyGu8P
f6sjBWNs9A8Or/4MMLHlCsh+QC/xdXY/koYKy0KLtyZdNCEQy/m4eP7qYogbw1RH3QvJBwO6drK7
x/18Gk2MH+gxfCVJ5LQfvoh8pI3fgVsRqWWw19vAs2Fa4A0Ok36NqjRAhN6l/uiq7MV+iXSIKVEz
lzlgroeINFH6CqFkSBjrOaa26qJSk8ZU4l3ulWDWC5+pDI1QT4XpRO6Q4xt8E5o/6xv7mhTBGNBY
+x16Vy85IDyCQ99bKrF4+dC9PVPGLgleE/MzIk5xtRu6JhxI3ZRBJ927ZQdmNdejdzEmCZb/hRao
9eKfcw3f/GpQG/6/uloCZrN2GcD/r3LitlgdXHqTZzKBwMJ5ogZ6JmZWf0pdzzfXRhn+CwRdRBbw
ZECoOeC0Z2ipQaLRnAADL1vyflI8SKX1KtAtRtJ/9jltFH1ZMIVoSbOewsIhpiK9s2zXexyRhr8f
hBDJa/i0gWwqZTk1QM1XOiHfZc5FCOW3WpeExvfRcmEfyvm7SU7nEMEjE5snCwOMSVpQrLknPPRw
+z6frLObtDyRlxYKFGm7f5VhvtmrHs1KKvaMLK8lZqJvGpRNRsOMdjd3RWAdFyLsMNLnpzy0bfGE
miHwptVIVT7/CpRM2yVSGQsLoz5/eSusYXjb2wC8+wHSMGmQkKKf72vrO54HD9Klkd3pQETo21UA
RNW1yvTmR+a+HryqAI42PlwBCYuLBwmDpZSUBJoo4m43qaqTPU1xZTt7g3qokfUniqPCVOZXx2rO
IHCej4X+aLrMYzT2qIgc9se5xPwxTwLtxAx5MoADKdDgVVA+RFely3MuFZInF5CmHbgprpb9Kjeo
2XeXZyxQN1yztY/6ERG1Nt4CuOZvoUWZ06YixTvjky43vF8pmoysP8tc7G0uHasjUFtU9eryVUbq
S/tbLYUG/V1R8r9e7Y+32j3lNn2G9YsgjRnbyDNoNAhg0RPJl8HWFqhoA0TjqxjmPekDYTrg6go2
23TF3arPaIc9atvxC3yaN4nP8ijaskCGTMYyzhkgjAawAJ2NlA5soXHyTagC/5hrb7AiyRItc2PU
ctxuilG8fPqEAG89LMExik2qO41hAD+Al8oTiJXpTtxaGQNig/RW9lzjo4YRUEuTnsqddXVlIN2P
AksossWpSJLCNbNihKBECOirIjuJLkoL1rX6LrNqyCXZUILT5o7Xu3FlgLIOLBVkOzvhAvepYBc8
XHqd8i1puvKAWI64hcATy6peRxBx6ZMUf0BMu7rZOAo2bxNXBNnmP+3ckvG/+x6cg8BfrAbvCxvz
RDmN/Klx/gt7p8xeIZBNYNqU/QSRHF5d4kvSWjYW7xV3wsUoyM2qn9U+i9xWYpOknFNtiymxPKsy
b9U7gpLec7cEB1n7BaXHIDcZMhbZbTmZ9djH+rRLI8qEYidns80OWAouphtjOz8RKOinFu/eUMAf
NAbhjk0Oie6mkfyNf1GJmbIpmuNrK22iZcF0wU52lSndq3b9YE7bnIDFe4dB2UEmbR6ySr9RofX0
MN0UNlclYHR8m2DKBJWcC9tKOJw7r6rWNgHy0SJZ5JbKdLBOQHnLu+4DhGR0uranOv7xyxqb1FRy
0TiwNpxV7eGvJbIDzn/NwtYN3WBuyX1UzkAlO2eu92VKphAamy8ubmajpBrv9HEB+1BuCEYF0wRw
xIFqXuT7mNguIc45v1ah8NeEdLys/0UI6pq3k0qDjSC6IpfbN9IK6a27eO3hRARq9ZBggPCc14YC
8xL7b1I1zKHz4vp5kMxAuGXu9Z7Der9O5ehDo8IqehdZQ7b3ip8PwMeER9HJJTrubMVnlEsK3jDR
YVhq0R1mkb0EFwo8ZO7cv0vA7nokhkmrmYsfYevWBBi2Gyob6pVB7rNSj/D3lm+iAhf/56Cidg+c
9HD0nyglyfLvVyF2uzEe+Kfb26K0SdrPA+25vUqJr7A34yxaYQ+dv5USL4KXd+Py2jYVGcfcE0zN
MMC/6feniHAzbV3GYS0TTKt/07E5au9/lSyYxHRjeQA1NO4MC0UrwKd7BsNkz0icXDVrnMo31flA
gCBokyBAmOAi0P4UTI/ZyS8qGii8X3kW8Rdso7TGR08G0rJL1xrhSsfDgFEXh1/s/9WYW5tFRL8h
JCBBwZJQhpoorIDMidBYFEgpW6LEoPRFksZh1/ZFsoywIXBVSQDLMYS8Ma1wwdArghKey0QMp+PC
CjUQ5nRhUsHEuS8a+9S7LNfW+tj0fLesJRXKWSEa3wT0NY2lof7TDhw1l93fD475t/asYJkXNgQT
wYx5qlpVjbCcH+DqdVJRf+7b6F9dI9nB5BSi053xTlS37zpOc9W1w5tQBbmb6Q7G+Zkzmr3+K9GP
7uQACeetsivGqGac6168/t/YlLgrya/6SYJTQdo5RtE7/fAAFOmghDTFwDIQeRi8vtkZnklQB8Cn
s6JB1bh6LCrz4LuKvkMAcW+h1l20nsmVPrvPux3X98xCp7a7Q5YX+mtyNKFXbslVHZHMk/6K32II
zx9IMXKumpCiQA1xvNquSotnN7eTFX8v1ny72zdK/eNmJ8zNMyRCIlieXauHLbExtufCqBcQ2wzz
ZRA9n+BWN0i9tP/cM1cy49qH2e3vczsuWc0Q/R+N0v8+N/8gnswLlPx+P/Tib4/GqOdb4MvOR+YT
y333EuDe1Q9rSXQmZ4u8ok/2Bt+cHqyNLS1c4o6HffU5xl/1kOpYhaSc3zfxI9pxoFHVnxZ4U78T
pALq5LRBKUWtH7ie0ip2GsV1qF9XrXZwrDosDaGYogS+CijT0qWn5R/EDFMlzfH19bTW9GYEem3Z
IlzJphFn7QUVn4j0UXYnqIMr6yzsoh4On4tvyhd+C1p0pDo2EzdLA0Zj8xBDzxMsAB6j6ik4GXBd
02pz1isP3yOuVDu3Rt8/RAnm8pRn9nJ29KOmsXNRIynkbfmYzz783vULimETGEKzX37/fV6I91oJ
U6w7QwW1e1C37Xl4g3y1O/MWnZERG+3T1017++lpmoSPrLbC6Luv+tcN4uimL1KLZ7gDoDhpasdc
g0SIexSgnl+lnZSYTaO3idjUGDXqkzExGJ+50oGVoFA/ZovKGrHaawScp4LbL7BeQe8wMczRZs0n
4BLE2nHlz2bffS42rKKfn0dkeLLtv+Aw+tREXEl4eHh+yrJnzPD+f1doqKKq3HkY/Rf/O0rpVbeY
VaY6PVl1aVU6HDF94uq1tE7TyAFrUd1M82WNRr7UQb78P//EHyZVjp3WlIxK1n5hLt4w09fUwt2S
2fAq20e5cPOBlco3GXXaT7FuGcGto2O7IN3i6orNujyNTE+/mMyW7GTFRUiIuH3gXxz0MGyDL4I+
aexIp9bl3owneTR6XdDzHqxxIQX+MbBEBI7FF82p3XFygXxoom85ltyDaLTPfuRTCjCfHEnIIa3u
BjhcfpV4DzcPgtBnHNcc3oZZRXlNFLpwDT3n114NDLxcrq02A7kUJP49rTlGSBvoAEkEcD4ESTK/
/9cKl0qwUDj0aSBfVH55taJIxZPDVElAMKsWA831Hcfr7Zo8SubpziwBmuLbm2dCoEcPwnJjjNSh
rtR5M+kKvXGi1NpxJMlpR56F9cN2e/OcUzVGWjICLdMX35mIyL+2dv57FOzEQR5eaKOlPOn88hfV
vtU9w9D1wa44DzWiVy3mYfkgWzA9a6iQ6lY9u1vfqgKj3CbloP+IwOIPGalb+8CK0rwlEzLjDpDd
+DIL5afRLrPwpgQYto4N1gFRlRtwER+sTZLq/fpUW/L14Dq8Y60nGSyNPBvzE3DIYD51ut3C5ziT
KVNuTv0o3bz8I47jzUrWsOJhtqDCSEd8JZHhyg2eqjnEBYaPQ2OB6yqLLMm/XwULH0+ZqiCONNud
j6VQTTsncRr16Q+NJP+dalS7NgxlajOAWcWz7PqtUdHO88Y9ieS6SFOXK/o9icZ7tBiKFwaDq+XM
qbQQgdbdhoIDGFsjMmPtbBPnCxPcESuoRLWRFmYrONpVY2twSFhHKYpL9tWM4VyFujt55JIAyFAn
kXyyrsFn1P4WHls8rX6ZHClzaSIfwgakXoPh8MmDIexxtrCYU3PHI26awUC4fqGC6JVE5ADZSAe/
hGCeNYzhhck1yThwDRMQeWGfqPKTlzDIZF0EXsvHVowK2ZQ6/kA2ANrmo0r3b0xx7pn0+tNw37TW
b0jf9qsTn8zkDICMXlEZNcX+VGQLMgOUm+b/dsXkrrXnqw53uI5uiNPAb6YZr72v+J74mw6ScB4g
DWecFVg1CPU8rw4vI3oWWJv6XRUDlpU6ayXMGnwQ7gaZ8pv+0N7GKXQEh+BRfw7sNL1r+iF6CZSR
RflNPqaMYfxx5Ym7tGuu9wzKAAqwtobYi3KvIzeD3HGHkJ9WN7rcHxwIew5j7iWrXQBP5x2s/vJJ
3ufllaZgOFC/BEGtD1IXAExg80OoECPA5MJuv8hGsvQnlz7wO4B3E5m9gd8gfjQ1nZL9z0ecMolf
LEsJB5Lh2kEQKYtbXyBVRTmZ/0k6XxmrEdiBotnjf2WM71woRJ+KVh/CJ6UZSBb+1N+xzj2d/+vf
L7ORWUA8kJ8XlnRIkt2JXlToXk/jz7/r5N9bacw6OTCA9R5X96aE5zs0j15EYtZKYqxk/iZDM4px
n8Po8f9q3oxHtNXpadgnmGBkYHdwYk6U9KJsFOSyojtZ3LmcAqqrymbhE5aZsLfiw7YPou8GLPSu
MFN9G7PhO5K87Ua9BbIRfrrjoiPXrX1eIdHfaoEvUACnCi/AA1VfETdPp+oiE15Lwi2LJKt8cFds
b1OMasxwdyjpt15vbvVcQ+6Mq0vOs8/gvN3ptLwGe0mbGHrkGdX/ssaRwCER3t0tTD3HaCfK8cKU
eU5eoypULA27Vjk63icDAh4mhztT4U8VRbi1L6E35um5FC8U7lPkMuuw/cr85NKl1tP4KckcAlXD
nSYPxata9LKHn5tQfNPHjzmvsgI2Ej76NzZ3gzHXxVru3xtrxliPwhs3ip/Ljvtlwcsy/MZDZYfe
UsimI2zECPhECRUfGG+/shVwEgl0Ozj0ziM0STXpN+ngDIvewAKSKCVPwYrYL0FsvJGOK4i0rGcT
uA4a1MywVIOXSS6/FgJ03yILS2ATK0m677Uo/2/MLmzNnx4Y2tS1KNIaoFnY3fKlLELHQt7BFgJ+
i9VJ5czGST7+/GGyFarJ/tf/SWey3zpt/Z7ClAZTTPOKNB0jK5joMHMLzsXd6KrMGLq1TaFYWil9
26V06G0jtDz9gNhGAYYqTk64FQH1vO0by8I9X3Y4C+/0Sb0r9/W6qxPx8BWporCfOSY5jq7u6A7p
/9p3KYKgEbkRcWPFIX8/XSmepHsBWUY9xG+gTXkpWixVkOEmDtV8OIEllP5tS+GWktHZLaCnj8/L
7hoasucJrXBcYpqS9jxuLizRN/r/KFMFcSd4aVFgvOAXmncdzQxT0m1Yc6toV+PFqV1UH0v9zK5U
Q20bq428dwsEs2erCqo6fWOI+IdFE0kH6DwQSeLOIrViR7Pxzdh2LN0QGdrl6Nn69KElFGh3aDol
UMlaooYGp3nPy5BDqKH7QLkzF5lpwsZAf5iVVZYiqNEo33nxf+/zbNkgifYx2MC02nD0AJ+v5z8A
XsPo892P+G9i+AiDSosSfcd/hI5XNGZTBh9ez4G8UhAMEstsf+2qCeNiUOu0+ZEXjl9cnYFmKfI7
HNxI/EwDhlPOZWDPEc3WUp3HoguzeYgSFtzyMKibY0Go91QR0gxZaHeIsVrnoDKcur88hqPsJPo4
KlVSrrAQ/PLbTOIMozlanz2jF+OBR/wBVeuaKocA/4ClAjpDTvaK7bmjWhR4arKT67ebNYKspHzY
yqU14vWtKJmSJj/2rnIa1+z0pDrDcSDQDeNwmH2iBPx1Zhk2c0cxlBFFqsDXm2MRHNe7V8UHzcMV
V2VoeBiwL/Ntq78z72CQbVE/jvCCld6ultNk7e4AYrj0CPu4aRmRHZBwgc71iom5UYuYhCjaX8Jg
5+hZ2Z7cPeBrfBD8PU2z/xRVJoJEAAXfvoABrP3ForH7KEPZcZmdmeiOynNspFqCDo/cAuTRcTaQ
1CTnJ4O3mBAngT6g0nm0nN5Dci8pZpBDa7PEe2p4bUKdSHgY6jxIe3NE7WCtJHqhbdJwfl/1iCpT
qTX29My7O+wJ8hAC7ObG3krWDrkY3C2lvtaa/g80oeGMaUymB6eHgfjOtV0zAANH+XXifs9Agmqz
RJeXWP9IdTR0aDAZLk0u0ojLw1SaJgKT3Ih0P6KeYLs33FDD4JXgDrmJ3yAIVbFA1O7rS1MxToBg
9J3KHGYJ62X/Jd9KXbo5YHBOL/lE8jET+LJthwoqhWUWAkxEFcc/on8uNrG66pnGVganAaNxqH08
CxynsBsCzqHYnfT8yRp6or3aobzzHlq5uvQvGegMIk7qvOqclY88pTdi4JbDqdkCacADv5syaqYq
Egj9xvn9NLIt9ievk4UQ5/PIRUuX1BXZ+fmqrac1tVvPJDnO1yRVi6fAIHWhFMcV0OoE7Uin931y
sVnVfzJUwrHTgOE8hmjuSM0cJo91+38Rw1qyZwNChyRo5YDKaofYoeBVbFqQCC49S+k0fLiaSxFl
LTDghrQ5C0dIYboC/hcHm/ympUITBmT8a7xsY1zsyNxjdFNV0FpeV4egPO0YSYLVPMaf+L9wfI2t
6nYIq08sC0z7fbwLFJNyuFeWX6E2lwgWb/6UOa0ZfkUS3baE00TT2wW164F8+UuXvwINKckGLPt6
9gKwT3C39qmSjmYwo1PKV+EnkUygd1PKfEbsH2IRpa0sZgILnC/2BrFBZlAJcYErdODtDgW3eqSw
dEk8t11P5ZPktqub3Djg6g6U9Pqr293L4PkR+FXnsaMRxtsKtvZ8xwJipTTCZmGDNTpYRrwDlrs5
+NHROYnF7Nq3xDlk/1DyPAtdn9k4EzdtU+j50qGy5ewDjYXJV2GeNuIHiR+GqKDzD/aBKWcOOEk9
0WTz3aYEPY85s3gmKOdfGuqevOchkpuKX8jbURVt4VXYyll3CyAfDHIknU/5dXWMsfWdD0rukCWL
n4V8kPNtHlnCT55GuYFJI/KvowPQ8cgLv1JXXsa5lnGBLNMZHPJ3WvD+ovao6rRrfi1antE32uhy
//LuzzM/VXWT31XWkl60UaTrjVCUT0O6BELlMu48tjQw/rrHqveGDLlDl5wm3anxMBwRIuw3457m
GlGZmtQF4r4wNzfHeSW0xMzoNeimfeORr9Q+tzZLE92S+r5mmCLJ9HlseHSIaX0Q10MRKHnk9Puu
o0eOMzpseuF2fwqufyQRBAsU3EwVg1NOCOu8r4D+pmJMDyA9zDOVbAKbixm0NM5lQmAVPdpBYcOJ
+2G+tVIwjIvvj0cyouLUuuIOpAEnyAQQPsxNh/hEyasEl6EFPhJ8nRwkS8Yn/R0HTxKSpZ1OUxtP
kPko/5QNrOKAZCCO+h5XI8dVfPq9feII5LMTYv+DCUXd3gks4tnXDlUNK0Rq3PIcGJFC4E+dHEOw
5EBcq+axlGyh2oNCEYD/rPmbLxlgDujKGSud6AcrgiJ94WeqWWIh91MNyVg7YaKukAffMIxi9KaY
QNA7iwt4lO+SZ1wMMuB9EuU40DXejlKapjISMCmxrYYWuCOefJm8TcuoF2SqZVxC8PxvBE+SMFjw
VjPVAfIOaHxzfByTjGTLrUFkDJEfvAsg2XyThoMzoNpxmg3rt47Un9/KKm6ECAywmff9SONN0jJT
kqWaTME55uOz0eaZo+JuI+JtVXHhYv/FlE65iu9OhGptPpaYtMtnrn/AHHj8IOF5lx5DjvAIxdz9
yNbaNOOpj/nvsVRFYtST6/Sy1vaNBtSi5mCcdQZyZp4rKuS8jfShCpnl5UFK5q0R0sN9+2TObjhf
boCtjOTaBq2YyPUhpevd/hVH9WYrwpLwvzF80PQMDtRyU1TZuB+FFBss2a9gRO4elzY7TjfHFRHC
ihlOf9M8qj2kvo9VaG2Ta2tCmh7wh8tT2KNLb+B058KUAiOqlAzjbnWxAolUvxl4VwfRnhe0cfcB
OJNpRqfSPZ+R4LVPE3IFBaElIzRs4RrxcqC1JfHgIEKnzmhJlGZfe9xXZ83gptJGXr8LYL9m1vy0
603t2Ynj4Sg4eA6olyrCdlaynAQ+f3PBWlveCT1KJtTr6/8S1DdJV/9cqMWgIl9JTWLiii2RGSCt
uVlbVkbqn15rjYZNK2pFHEwfAF/AAoWAhM+KQUuLakJn8BMamN08qvHXmR0qj0B1Ywkrix5qul7W
IXJe3PSrmMk4g3HepNcpIz3m2mrqnBexjqsAvVh7RimGSnZ+qh+3XqRkyfYcujRzYrtaljN8/4pU
+vd7770A8oQKtpt3dITMjWghayKqYNLgZ23CXHvjxXrYM8J3gc72n8+X+WwNU1vSg17gmXlP0nwb
sCsY2T2ovKyZxati3vPULnrB4mW6Z2dAgv7upjLI7jU25i2jxYRlJth73mYpHyNaikfEaITF9/3D
gExzGGeMagzCMlMSqbJaWCccJIce61xPtHDD7JaiI1Cb34IQonks8RTzxQufe4Mv6wLEKVaQ4VM9
XY3PhmJQ8VRLZxV/wIy8sn1OV8dKVzDTvXFzJSXbJHuB3lEAHsWEhr5vdMjCO/QBzz30bEYQA4HK
wsDKPTx487aVIKFPlxCZ8LYteZ/6yAqc8RPNrzlLQsZRrLZGA9Kj+E+kjh/Sg7dIeD7XmUEc7Vln
8bNs7tY0EuQi+GF+T0B3951Db+IpKRfZE9x/Xzu+kARItqGs5Tg2kaNKpbsHjdRSPTZgtZI8wk4e
2NMPbxv4xHBWKHEffwdj/UpIkpWhMJz41s3fbymQEFOtdT0L2MxRKqjyTtp9Dl6WnobyzV9FCpxu
M7LJbaL/Os/gVNNLA77Pl1K6PNJDWJwg15gHwuz3W1k9A+ZdL9/g8wFwjmXUAfEufWczJ3dNH96+
hUbKGypqKw7JC3YfGFxxLepmKR+ZKNhz+Azk1EmzDmx/hUsf37P/K2fpOxOFq2Hkp4xYvsNezewL
FOfD4BkxxkZsbmRGPb4KyqZdPc4EByqJw2FLFO9t89GtrT5OFW75O56nS5TbQQKgyZ/gETGO0yw1
/pe562JraRV3bMr8dtqZW1X7QO5M9UFlcgyFyGi0HD9X4RRYHiJa54qMAZrjFDo2dONouTKrPTn6
0pebe4NZi/dxfA7B8H9j48NXe6fv6o+jM7os6DyTh5PZqTg9fFlaT8TW94CetKfbaBQcQTGlO9mT
/f9dvbgQg/2eWY5cnRjaUhdZDnKNKj5KUnv5XXDZixCJ1Sv1JyjlIA11eikwbRj5PIMfoNMFx9rf
kq87VFDDDrxPXvd77zJ4AGjc/kgOWYB1BYF+W+e9RbzRE8j+qzrmzEaZds9bddG1bPmrQpYB4uSu
ZjmkfMEBg116gxlMOC4ZW2MXa6NR+MAXJrGk8bkQyzu+3ey9fFET8ucvXyOQ1fODZ6GV3YhMoygo
tJ+d4a7Y9EW2Orkx43zwCrlVs+OlTzg2Oxd4rtcNM/iaQmB3WinMEQqbiOYJuBmhaCpnQEBSXiUL
AKFhtAo47fOvJjDrgEpTKwQbaku4YA6HJXpYgQIUSaDZ+o5ZFwTAVRGgKU8ndLHAYR26Urwntu3W
ZkeV+Dpidn8huNwerzxWgOELw6RSIPK/BWB0BKRVzgD222lfIiMnH6M95JVEfoX5LXgkVMT0qZam
J2VIEeBRJpqzxGU0/Gz/nFKYmjZ5t4z0hB66tEDgmYdvshkLfzzXZ328WYh+NGo0/vvKhkUef2rp
7Ux6WpTU3gFvSIylt5SRBQ6QxjLvKKYGA/Lrm1qMhYclBPy+mPjswelzlFIuC7aiOB4cwNnwL6gz
fDPCucNi2qTsev+LhSc9FoHcGxQyvFe+SmVWheBR6yUMKuAI0zsE9M6+27jM6KM1bT76Zb6Tq2QH
4tl7eiCGidW1YVP04pOo9AZxbdR+F1kzh1ER+MDRJFrz053g9Xxgnml4nxK2Qb7nZgog90HhhieM
GyM98ZZlPKAR13S2dc7BIZNILIOR8vx7yfc9oMaWJ60/uhwzSexysfrl8x0Ydd+a/kjhuqUI508p
DeknDTjEAmuTAXdfYvVBjNzJStzUYNRW6NSULIMpyy0qfRJFM4s+iaAT/rBL/V3J6mDAGp3GoCvS
EDbm2MypGuCrmCJc3UChqAc8Y6rXaibIOULW9kwM4DCiNsBH5eUyYi7/Yj8j1YkgyEpknDqO5Xiz
9j+JXKmWCbRfaBJa8wh5W/PYdT8sS75GpOmlQM4oZGiT3xA8fTX4+h4fNqRhW/DqabgzSielCd42
D736QVvsadOnTvZcn1E0QOfIuPCZyG/syepRrMUYqaNNRwmjIOCjUD2ZA54uK/m1l7gm84o5nlWV
Cl5IfNo4leNZKFYdvawjbjwPFpFxwiBPCi3WyProHnW7hyunl8vPnTgluHsxpyIPuWGVy5go6HBC
7Jq/tnM2ZWoKv+jasJy0bK13QHtdthdC8V5GqtNHcZOYP24a/KjIcDfZlVKy73g0iBh7bnepivmD
XDv3CZaMVAVizUil5nu+TflXF5/F96Z1T4BLq2NERTlNKFIE3grW/+DriLefa+EoeINwJ2iJHxdo
Df8tk7GCvDu0o6iSJeDdSVhUqGuATUtie95J/xvjkJ9V4K0QxOuD1sk9pVcT9gemxmnBOj35AaJa
MwwSs1G8g81QHsUdk4UhEgXtLqOykqneN71rsVtJl6/Wt/c94A9AcrYMQJku1nq4VEOtp37tRcTp
vHDSuZeAzVzxcS7WUxiisBk/wuze0MRm1Rs6xkEWmoOx43bmQJrtVghXIzSHyDlgJripYHI22GnX
AFWBycRURAnczUqASzSC0uKCytmD/8GoipwiLdu44ZWUerxjyrQMpa7ZXv78jSDEdwnYDwU3GbYO
WjCGO8AvyKnERDwvMoK2gXqmhq4PFR/fhDMs59lXAxh8Apv2WhRQDeWuSwpYQf1387TtEW09Odgl
I3I6+Jz34NXf9l3DkPK8CqpKEktaghXOzTS9AATiGptj762mxcuINKdlPnXqHcfTxJLuFJlJeK+Y
3vDWgFzQROwoCFzZXCQ2RDLKNwCVeEgOwaRcDorKrs2FxzxydLVfsOXxl8pngjksSPK+MPbjnkWx
uYsaZ37RE+qvtd+4OAC90yqaQ4/Dt34m3ozxCSI+47X8mVfHJ+xlm3p1DEH/AWn5qCAGhyti7HlY
YVD0fuh/lPjuhsI63dyBUU/Ikopu86CQotm+rgUnRT1jvJ5LWBFhHZID4jmBme4+0AjslRjGjM4H
DHzGZluNr8xZ4UMf2m97CHZt0Gv8lvrJFhGGZ2Uj2+o0xmwBWSHwWgedM/V7nC3mktE0bAaU3Ix4
11ap2iEbBAF6yJwVzUveTedo1ezqc/3uxZAgEBY5dY5g0VQFblQu+AdjrXWtmLfOZ5rTulWO1UPs
KeNtEnOghVMibyNSPEZNPHPZPsPwAq9pPT+BU9CbgKs/vonBJa334UHLHgkv/jzVieZmpIH2s/KS
aDHgCJ3OujPXZxSTKeasbSkMadh+t6WpE4Z+ER9TZIFG8iJ2sBbKFZde7/sgCMGcfGRHxScYjSoS
JzgeyLKqOIVR/VRJrsREX8GixgvcT9KC2W75um2GuBT2e1aKnYMysYnKyeFcQN9Yc3k/3k+jM7H6
LkRdcJKl67EIWtWlwfRbdlxOILgCEA/IdizEpKDK2OdQkCuFcyiwESvIcRC0SSlgMA5PHfbOlm0c
/ldeunpuSN2fW/DPLvmaPaQevKWzv7s0fpXtQb85qGeQWdeFROoBO42mje1lrDQalXhPqG6i772d
MEVv1ZDLIuzRL6yqm9znllHfA+Rlxvpede9dtnQbtpRqOkTjEx8HUPNiAlZ3U+e3sAla33hUW5W9
fTt2aJchYP0UHVtGKMUZyVWMXQmQaGFcqdO5+1r8MTE+uA9OYAFEoQp9lByEQZapVyQUf63Te5Bj
fUUeOemsff0/ip2tVaaFstpLDAu9ybrKwMVJthXzk/7NGoz0LZ/f+oOTZExvDj7zFkrdiQ0UiULv
hAasR0kwmvbpUe2gd8crz4XiMxxaY6G/ydlcf/j51NX6ZQXDwu4hFeNYk3bv3FfEuO1F0AdP0Q+o
U4pCSdRLK1r6ugINTRUnuPO9pHruU6X1wqzwr7ZgbQ4ggoGsquUlWfQST/VtOY7jm7DUKLLF0xeE
6LsbY65dJWQ0Z4qUrhH4ZQ4j9SNkCcd4Peot/kNT/1n9dNDAINDRXV4jBNLORk8X4t8dVgB4vL71
myilQMmpo56tyOrCh28ySXftv76jTV2Bey4IHdM9/SsFdFg/rZLETcQL8HGuAUk9REBEubC9am1q
bG73zSe2T0WAkotPzAMzAHNueH2S4dUc2j7HUs6ViSDB936EgVbkW29MWHWF2GS88HVE/t3WoocM
4/8v8PvmmOyxx5dkTTMFvb5K83enMd+yb9/KsjSTqDTZ9jEogi/08eIpQiHdp7DnrCry0Vi8lg0E
785LL9FKsQ3JhmQkU6UwQMxp5cejwlDVul6FP2TA22bNCDdEnxeFYuaER1HqOeMHkgcaUeTOjy1z
jzfjDL2oVEIL3DDGZ5547I7sDw6tUoJhJyue0v5FkT8OCRgKl+5C22bqlmIbcGJ9W/bLWFh56l35
9/YosRmZziw6Xt+yVYTi0d38Ye3USa3pnIndeXICPA1uJqWSHvSoVfDdMbhqSxvzdlxgMslkMi+z
Ll8fWlPbDVH1NJ4dqx19Kw6zmOwHms7tkRTeCaOaR79impD1aOWIIwAdD1UAcEhNJ1qcqGe0DsU7
FUDDbuZyVCcRs0y2XszF806Hs0/mzvZVS0qEMRYvYEdtyD+Ab0a72rb37gwptgZpX0ut6mIDYx9j
qs1G5rAzUXKZzlxwMmxPpkZOv5VaJQLjyWU5ve7yqcWSXpIomwcsvUT9QWFq9PMzj/p7YM7TR0aa
4b74cG9l8jiqxlmNdPEs4fy60TO7P1bhLTHgec3EKruayGjrx/AKvBb4sdP5Np62alDoqeiNOQ7J
E5CfG7g35Hmkrp6Pcqm/df3g8xohrz8qpH16XO/NWVVwATxa6q4DuhjEsa7OA//EJypRzJ7llJjF
rPC8drO1U1DtOCNWAFZ4rO+vFPS6OxxTqxaA4rn3Nn6ujWq/dGIf4ETGN1TUcNDP03+9CqgS1ETj
YGvmpd3Xcf34+MWyXKgFl5ptJS1BnxrS2bsVrNPnJ8wkPTsgPF1tL4uy5C56yf6wrLQOi3F5G+PW
DDNY9dRcjThs8Jjxt6oyo+qcblQ54sS93rJyNr/O0owe+HcmCc+7AW9zSXomdw1poS9VKUrJ5CTd
R93z4eM8hOQ70ZOefx3ay1qxMpIZULC2fpfHtteeTd6wtxxNePKwkRNzJOgHWgUxSRH75rBuqxFD
gzo5XqK7VLs+Zmcy7Xyy6JzgrXvx8ShPqFUAOGQY2jOIgHb3Ezk7zCDPBvBYkR2LmxSDW7xClz3Q
2szt83YhQLW7j0lkOLNp3gBdxRbZuYpePQ==
`protect end_protected
