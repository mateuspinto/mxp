XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���2�O]S�.�ļ�)&j�ݕ��£���u)[���p�u�q�x�92�	r��o�U�s����P���o�ua�hdA�X��Ӊ}�	�B�t­ 8�h�u�'1��	L����ûF���4��*��0��{:���	z��5D�.�i�=�l�%J;��"h�z�2O<`�� �\g^݁�)yr�;���*@{�vC���S��[�%����-�r�D�| ��2H=-o�ad%r�K�A�9I7���.�j����i�E6l�P�|Lx�8m��xn)�&���*(�n(`�?i�Zߏy1���(�#%cd�4�Ju��*�8��1�D�(|9\Ë��/ѹ��D� �H�6\�pI�	��XFk~��}���}_5Q&� �!�t+�*�|��@)��ű��_�83�!�t#o;FԺ�=T���$����$����*�y �Ѽ�d���
�T�&�f�(A �n�Xc��ܳ3B�HQ �qɒ���<g�w��x|(q��>ů�K����(`%T�wDG�e5?����cΦ��1%L����� ���_l�e4�����ZRY�	$������ v�f�ȝ�d@�ď�+h�z_2����̨���=��	�{�8���+����eW�E�k	���-.,�4#��a��g�+#o}�W3)Ѻ�Jj.�Т����#��K`��y��.?o~U��
��C�grjܽ&x�}�R/f��J�F��^/�P�]K���P?}�E"3ڸ����k�o��h���Z�7��W���<СXlxVHYEB     400     1e0Q+eb�{��V�Nq#b��%eR�"��^J�"��tz����#+�2�[���S��@.�7���M���I?�/jԍr�jRV�s����&L{*�9]�#j�S21\'��^8k�
SD�@@;g��S57�>4�� @��po�)3�*�?Sf�[Ǩ�PI|��z��� D�_���\;��lD�ݴ�\ �%�����Ѐ�6�A�G�%L�FlJ�üt 9�H���K�R�K !!��f[��D�j3��ICNЛQ�,����g�����`m�&")�o�`{c)��V�y���1�h�Pz���Z��e�}|m�Ok�!	`��ƷBu��/1�|�jf�JC��v�^ۍ�Pa��^�+�M�[v\����
:z��Ѓ�fr3CK'Y�K���,�J���m`�?�c/�g�P�s:�@Ƅz�� `�v၃�������=��=%�!ոL,t.i���軴ٗ>����~܄�?�BXlxVHYEB     400     130@Y7eK�sU��,�%c��D!��I�*y^F� UW��*w7�5F"�B1k=D'�r��TH'=�r�h.��6�gW`��oYDS_O�$O_�_ʥ�SJl���j��1���dY�G��c��@#)�@{ֺ@� ���xS�f�����dF���[��75
�9^�Y���ŭ��27;oXǞ��'���n�)=���ۙ����@f�7�d�Zl��Ŏˡ�i�ӏ/\H9u�� q��Rm#j,x�?�*U�$7}�b�e�9�� �Q't"=�&�GI���W`�ڠJ�q��J�� ����7JXlxVHYEB     400      e0;���0�3};�@t�d+U���	����̏x�����e��GM<u邯�r���B�]���hQ����3��df(�r�񦜡������B?@WI{��.�`��`����d�6�2nS��! �w�)6���`� �V�*L�:�������j�=��\�t���Jq8'r��t��&�Ұ��H���CYa��Ɗ�����Ⴝɨ�+ۈ� ��eȋH�2*XlxVHYEB     400      e0���hJ�ϯWtf�N\��j=�w���&��e=���*�!g���b��N�¬���=a»�G쏽o�/5�r�Ŵ6�g��_���W��op�jV��\"��Ū��E)p��J5�oO�����XI��D���)���d�8���4��A���ټ+g'Q����� ތoj�/t;R�v�G<�0���C� �lP$$��s����J��r�����ъ���c�p0��IXlxVHYEB     400      e0;2<��"
��p��X�3O̓C��5 R˚�~\r٩ܠt{w�2S_�������+R��,U=����۴��Hd�$n�P)�)<��>�1��@�uc�g�oA��c�o�4����	������?���y���#��p�W}Z�[$k��M�6�d���ެ�Z�!N"h��0��e�?r�瓂h��N�q���*�Ϸ0!�_y�C8ǅ������9fIQ,\'/XlxVHYEB     400      e0LzZ}���ls�S�����@ry��4:�h�b;����l[z2k�Q��L5v����s��"*O(�ПJ9�	�x����ig��o�*T�日2������7.9uQw�?�����n���'�eKb�K.ɢ�@������(�/�0���z��oq����a��R	�;'G�ހ�\ A�c?�.tnY�(|S��L�)v�ҳǏh���
>��=����n�B�=XlxVHYEB     400      e0�na@k!Zy8^��e��)ɘʜ�'Bn��W���$���^�<5i�/��~N*�qd&yy0�Q��>�RL	x�ce�B8ګJ��p���7�ͻVJ1d�_�����&�Ll�lp~���&A$1x<n��J��Fp�B�΂�.��% ��1���ɦ�U�28�R-�q�{�~虍��<�My!w��}c�勠u�ar�#Oϰ�wx��:���W�P�;XlxVHYEB     400      e0(y�m���nTg!@=��M���������XzxH�5��QE��\ �R��_q O��z���j-:p%�.����]�����3��P��p�39D�|�=-Z�-����:=��K�B��/����=���@%+�Ĵ�=KT�vej//������U��8�[$�`�=�M�a��v�.g1$o��-�+����ƸR#�$Xഭ�Po�"E��"XlxVHYEB     400     1a0�����=d$0
�Mo�G�I�R��otY�ЅU$�M�2i8���/�����(
N[[��b���p|%(��uj�_�E�~�ȑ�y��`[x9�6����T�W���sSX<�]>��P9B��_�S÷:tK�	-P�ѭ��r�*��h`��w��&U��m��ɭM���>[1F�T�WB���`�=����)��MGdZ?&[m�(r������-��L�"���K�����}P���&@�]8%.���Pw�<��6~��_�ތ'~��A�ZJc~=%�O��V�'�����|��i?ET��a���.ڼ��a�r�Ý%:�\��4w����ǆNi9>��]ߡ:ϼ���U'Q���*Es`�-�b%l�Z?���S ��K��ݤgc��[֦B.*7� �XlxVHYEB     400     110��V}����P�+�z��u�	M`��H)�#���5� �9QD�5����Q`���!ʰ�c}�()/ �̷S���y�G�{�S�*��_�}�[����IÊݣ �'��r�1^���*V�+p�Y^�q
�+��1X�a8^�����4�����\;�$Z�B�.S`��Z�
@�����HS��V"K�Q���dU�����R�';����ibtr����"N���;���B�(g$��8��W���>�+՗�l����cmK�:Y�S�XlxVHYEB     400     180r�.��m���]
�z^X׮7o�um	U4�YR2k���Ձ�mFJ����4�29b�i#媱?w���=D��S��!YJ �b���b#���(>H����f=�n%��E�շ�S�7��5���EKN�M�Z��e'~b�]�ES��7E�
�FJ��z˃9/���B�,k/d|a�ș,�|@Y��{8���''�M��O�wĈH7`2Z5��r�]<���},��ѯ-��	����)v�1� �թ4��	h�C�k(H�HL] �<_�ye64Y 8X�@\T]�7ਛ�^�&*������֩%��q�&`{�Z��
w3��� �����޺C{s0:��݀���,v���K��R�y��}Ьy�}�5G���s,��=���XlxVHYEB     400     120��P��} &3��$��@D��K��wM��yr0��cHFkP��:�5���dm�9�{[�,�,���QTӽq�&�����wDcL�m�Se�0��������o`ԪG%T]zk��,����oT-�J�ؐ� |�tm��-%���Я��:h�<�QHF����y�
���}ų1��}��� �y
��.���w�H9��"�����8r��I�{�Ý��� ^Ͼ�5^���Ы_"�cB)�u����"B�yD;��z+�b�Z.�-0�)�3�a2>G`(˘���R�A����H�XlxVHYEB     400     130����_1&|G��W�?'�2��߰�LX�'c�5`�&�eı�&3�U�88�F2�$��Hk~n�5>#�>2��k�V��V�.����\}��s��4��{/twV�O�B{^��o��Kkg�����0�)�^���VF<�%$l_�0a�ǕM�R�Q��Q��kX�\�'���R�2����`e3��%���n�[#�U%��蛆�M�C-4=v����`-�R�d 'By��溸�L�
�4T�6񄼄ww��:�}��S�3�% !��Pt��~�]�-8�S���㴱��v�M�9�0J���-��]XlxVHYEB     400     120?��<o,�􎝯3ʕ`�i�Ƚ�l_�v�5�L+8����e�����ʋ4-�lW�� {��A������CX�3�h����6Ӎ�M@np�Cꖂ�r!��:�-#�	�o� ��o��O�:��q���r��uF+�U�ªS�vB��Yp�9K`�B-���;�,��(�퍛�䛗���]
էa!WOݻ�,an�ZwǮ-� ie�3��������&U]vIɫ*��3��r�MKv�\0���*�|F�iY#�;�>�y+I��2yu�?��s����#��8n��PEؠ�5�XlxVHYEB     400     1404�A�Ă:��&���D\IA��҈�����>�Y^G���3q�[>[`#�:W��y��H��?�7�3��ra�䙼�U�2>�펬ܹ�5רK��C�0�;ۦ�����\���w%uy����x�d2*�i��ۏ!��M{��.�ƿU�ECQ�Ms_�)���C�X��-����s�&�{h���{��Yt��F��`y�ٶP�N!�L��������"�w�9��7:�@Lq#7\B"����D@�o_��/�*�����0�-"��%�_��"Rp�����O���k���\#��ځ�XlxVHYEB     400     140������]�7�~�F0￦D0�'�q�=7L�DhRɞ�	����@�^�n�o�˝�C�o�Qۥ*��Fb�c�<�wC�b��`̜����kx�C�ڹ��Lw'۽�)��q��#�z2�0�e:7SO0&�*�x
������#���l�$76�Ƹ�y	^jb�e��h�z�7��|@H����	x�%b�vk�D�Q4����������βtz��BN��6Ku�̚^E}G��;i�S@��V����х�������.�U���u2ku��u��qLы�X���Ñ��MTbH��(�s��/���#�n��n!�XlxVHYEB     400     120��nhgp�E�m1��c�#����c9�8����A���w��'�[�@	K&Ps����{�dW�2?���l,�jWw(�����4�9�U������Ӧ�O�Uf���$u�d��}�˵H�N{�革��?�����Vj��%��%#ba�7��;�%�;T�.[f�aUIH���a�3�u�-�u���:>k]V����i�1uY���7\�mH'[����x��WCɞ��j��C�����a��l����XQF�C�.��nJ� �4�ڡ6�Z��`�E���b]��&�{�XlxVHYEB     400     140�����\i��|\̓��g~��ap%Dŷđ��m��,`~�D����
�9C��T�_���.f�\{0Iَ�TU����F�є<�HC��z7�w�L�2��Hxo��,�8`�0m��~D�����M�y����r��]ڦY�ʆ"��7֑��n)xv��c�t6+Ӊ��0�h9����H��8J��+�|�ߐl�-c
���ѯ��IC�N��O�D���Bu4��[�z�>�\�&5{Y_�EJC��������h�?+�4�����v[ŋ2�2i���:ګ��m�V8	M���~�5�E������h�
�:�XlxVHYEB     400     120�{�z�:f��ɫ�~q��b
����`��ٿ&�܅m��Ő/�j��C�.�f�z&� �?�Z�@G�~��*z֑Ev�R���UY�ho�C����q*U�2��hE�������or1,%O�O[��O��lįʺ�50ۗ�I�k���j��K�>{������mGP�r�=p��\�J�c�ލ�ȃ������ס,���.�3J�.I��C�,f��QW�ussp`���[U�k�o��'IJ!`G+f�g��ں�D�t���'��ѩ$X Kޚ�ۗ mAyn8�PXlxVHYEB     400     130�늣��}���LԶ;!'J�iu��q;�ڿ��p쫻���}q�JL����C�h.D�#&'l��?N��#�ɭ��߳ء�O� �Y������k�Jq�Y;$S�`�E� ���g�8�Q8<�Y߳5���B����9�=�({a�yC��� ��e�,h�����Υk󪂨`/�$[
&ua�����D�i ���5Y�m�K®�?�~.)4�	k�A[�Nq�i�Rqx�"�-2q�BT�3�Yx�!�Ѳ9-��*��[�}�r�/���W�~	�P�/tdp�)��	xlZF�;�XlxVHYEB     400     120�Z��	�3&���oV��MZV����q�[f"�a�,'��|G���*��v�֩��s!1�+QVra��ϗ��8
��>ɸ�aN��2!� ZPF�U�D��/ݕ��C�3�;G<M>�$C؋{S	}RWC�7!�!��'�6S��Ԯ'��d*�&I��PC��nӸ��r�Kp�Jr�M�/�2Di\dT�At�/��r��Luk� `�z��#֖�'0��q ��i��}�(�q��!{#�b]x2_b�ʓ.�U�i���L��/�ٹ0���Ƙ��h��F����XlxVHYEB     400     140��96��q���fh��R!���E��B����h�ax�߅a�!�
+tP8d�9��M8�<�V�dTT�;�w�F��/�<A��g;�D��:��C�]��p�ևr�e_\����Hs���\a��t�|R(2�f~�ڣ-v�u�:�ʑ���d���<����j�ji]�p���1�I>��FX�PL٢���-^�OD����s��Kg��R]���LVRu������[A�J3ǹ�b�H��O���ƣ���~S����洷)4�ޕ�f����me	vɨ>w��E����)�M�p��H�r� 7����Q//��JyXlxVHYEB     400     140������]�7�~ф��̷�Z�(-8't�H���|1뗆����5����Әb;g9�4��c�:��|-yi��\a���Ġ��
��H(uƣꏕ{��1#��JYCS������b��#�Xǐ=v-�j��[�Y���ǣSr/
N�@*��7�h�$���;�����ۤ�����S�|����'O?2���z6Y'�!|AXiO�����f������|౏�Ӽ�EC��~�)U����#4��`��$�������uL�CT��y�P�e�6SN�f�����sH_���{�֏���7&CV�PXlxVHYEB     400     120�EN7���`gϊ�M��E�w�6����s8k�O�T����DW�HnuA�^�}������l">��l*���4�+��=�Ll Z�,��2w���^Ṃ���F�JHw���������^߬���,ue��.��#�v!����:�˒�%^ID�E���q[��}���+|�#`�m�׋�Jt�:c�Kk�G��cǚ��|�� �p8pB:�=���M�A�IK,��+m,r!Ltm;�d�
�����Dy��������/E|0�"ӂD�6� ��XlxVHYEB     400     140lK^Zܛ~�W����1T�r���EEPS]��ѬO�J���2i�5G��U���K��aߢ Ş;st?����ٽ	{yɟO�����P����:�d�^��g�υ���(��~��&��:�.�O�!���iG��'�T2�U�jȄ4��t����9�v�hX��R���Z����u����h�^���#�Z&� ڀR�ݨP��f�����~z	́}ʫ��-�C���pM�zǏ����^7�O��aS���r8Zm�?##.V��u�f�$�v}��i�g���+�2�9h�9�y]Aۏ��E�"Z� �K���XlxVHYEB     400     120�{�z�:f��ɫ�~q"��Z���H`�sh�b�_�{k͝%'�={�Xa�3�8VY=��L�{�	���Muwm��ޞ�l��d�(C%��#qǄ��Gӥf�,�� ��5��D���H��Q�oE�`n
;j��_%�r�]i�V?ͣ���z��S~�J����T򘴱��P�I
c���4}A�s���a�c�&Q� �:V��#���@Klrz��#&3c��ّ����B(�Ʃ��B<C+��aD��(�_Y1��p�L٣/pT��6O��m�i���cXlxVHYEB     400     130/�W�R��K�DB����Cy��;�G7��j}������@��=�]KB~Ǘ<�OL
��YOWa���|	���,�#i�+J�PRެ�8�����KdK�[~���ܤ�u��lIR��%����lA>]�C4��x���ޙ�:D�x��$��BJHABP�!�O9����o��[�9���\�>�Y����sNb?�n��q,�'lB���LN@%���+�����jU��Mm)(C��k�1�'|x��h,�\�|#�?M�͏��k������|)�c/Jˌ�J�Hw��|Ƭơ�0��Ta��XlxVHYEB     400     130=�e!=�r#M�"�.ɕ�KVZ�FC��Ӣ���J��a�{w;2��kP�2��8���}+.TOĹޜˌ��yF�1�R��&2��Ok>.91�lC�T�j;�A����Z�9��X��gt���?#ϕ���g�6��|���u-�p�La�%��,L}��}2��58�+u�Ó4���Ȥ۬���5�^Y��lp`a]N�a�V��<�x;���̤�A�5g��d�a� 4�滉n�|�'5�=Frz5���怷f8�>݋l�B���kC
��R������WR��K}OP!kfrN��A�	XlxVHYEB     400     1408��m_VdD�م�� z(�7�xLg��%D�P��I4���V~;�ޠCK�l���L���B�6[�E3�]L!u#K����~��7�:j7�pCuTA'�\A���	�y��$h�{� ൳��r����1%�M�w�˭�[�<U��o��k��IY��!Cz'wG��'h_���(�8j��{�CoV����#	=�q��*�����^�v,�f�O�2���4�%�� ͌�4��}(]��-n1���/���~6���m�W��2��oM�.���;?�������:��6���\ֹp����O� ��DV�rz'G�rQXlxVHYEB     400     150������]�7�~����t%$c����+�]�rt rQ���4���Ix��"��:��,]�دnqX%d�|!y�5��c�T���Ce��,�b�?���JjP���=
A9pa�G�xiSݧ>:ґ�C9����Ӆ��0�IKZ�N���`jE��6���kU9��-��&��j\W9F�F;��33�{�h*��_���lND��3�sz���ڇEA����O=<I�
1�b����M5Y��7��Y.񆰿��Zԣ��ZK���?��>Y�q�)�{Iϼ	�r3���7�4����������k4@��lp�M��J��?XlxVHYEB     400     120���}����<����r�C�Y�>�D�����
�Z�e�)�57�d����S�<�*�<�<7�v�dw[L��;�iq�Ú������Zx�]5/m�Q�Hc�M�����YM���z������H�j2h��ޑ)�����_?uV%8�]/l�IBn3�?��dT�Q<⚿��AA{S���+����$��cH<6�pO��~&'�)��?�����l�p��<����Eї8E�������Qoh��elʱ♺��caG����B �Ӕ?������#�wY��XlxVHYEB     400     140�5�����6�D�6f�Mb����W7��\cF�+B t>�8c)�K9���+jx��͘p��(����s!1P¡�t���uSG���pˈ(���6���a1tȾ[-u_<���j�z�g/^דv���§���7��֚jE�f��5o9T�[X��Ϡ3�ABԵ��5����_�V[!g�2�?�e����v����o�ഴ{��܈���yVEs�Q����`4�"�nդ>�;�~@u�^�#�"�͹����,D
���Ġ��n��l��y�.j5���/n|8JQ�Q�i�w��Ү}����: ���XlxVHYEB     400     120�[��e5-�>���
�(+S���,�x��}D|�@�c���H�4=,�81�#�܋�K�p�C��S�fxp𙲾_~ы�w�*d��2�ݲ�&̂b�1����H�e%���|M' �ũf!ǩ&�K.P���G�Eu�z7FL��"�kf��E���������ƿ����A}�0�[����&�r�_��I#1z�X};{|p��%|-��C���'2���`�և@���Wa�gס��.Q��)��πω%� '��@`��%Ω+��a��k��'ä�*XlxVHYEB     400     130�늣��}���LԶ;���G�|�Pm��
SY��S��ߦ ���m�"}�������=A�u��77��`���L粨3���(�� R�VK+�*��j�];��7�ɵ�4h�W�l�rk���)pAC�����"�Ij�u���f�%mD�-'�Q��~&s�`ؗ��ޗ�]#Y���L�K+Jɨ����[�*|�Q�o���Ҁ�Rn{�������"9̮�H"W�C�(߱�����?��P@U�bg��
�G�|W.Y�G��?A�,���W.��� �[.����):5�ioXlxVHYEB     400     130=�e!=�r#M�"�.�8���_{�}�7 ��{NH��������T-�;n�1���i�b�ę֏�df_P��
؞�Z����*V*@�Ev�
UC�D��z8X���7	����:A��I�s�c�J���D������	Ƕ�ڽ��1�z9�U�w�B,�:�N[��*6I�>R1��5��5x��X�{z"������o����:�{��f���<����~ֻ�rO8L����?��(��=3+��?��B�Bd�mi�h�o~g�=�&�2Bz'Srq�q�h�9ۼn��(��
�KP�4�/��XjXlxVHYEB     400     140_2#��[��pu�mY�b��o��ٖ�Mco1�W0s��蔌�o1"OT�m�a�'j7�`1@y5<�9b7H�gO�q��G��6����	���v;9�@�x�B��5����r�/h6 O{K��bR2����i��f�`o��0���.�8$�Y~�*6- ߧ&&;��'�<�b�Q`�#�)m��Ɛ���#��$7����}��e���]�d|��Z�Qo�WB�빁��x���~�֍�if5�tn���F��P���/��m�U�wm4B5L�}�Hol_�v�	��wa���xڪ��%z�CXlxVHYEB     400     150������]�7�~����<ZP��8���@�#���-+�L����8C�a ��tk>��(�-�
X����T�<��������j�F�����Ls�]z������2��+�\�5f�F�L,8-_�د�YQ����^lxO�|E��0��X~ߍ���.�@'V�_~��B��Y'r	��A�<2�o�!�o����2��������Zd|���%���S�LP�C$����Ƿڑa�H�Uκ��H3��5�v�{�]���%�[oB�dQ��RX����)j��=!]E}���~�����6�M*g��9��>ć�����H�T�m�����a�XlxVHYEB     400     110��z�r������ܯ
@:�8=75���k�J曫�Z	�頤X�ڙ7Cv�ۿm���cO*vf$����0��{�~��	�S�}ֳs��ߤ�
	Q�!$fE��K�������H�J�e�5z��=���$�Y�����k-7�~��q \64f���kdT�Kk/�"J��
�r�k� Y�\��R����`XK;�/��3�L����S�.�iRj�î?m�+*���sQ�5%�pƌ*�!��+j��Ϸ���U�m �Q۫����2���f�XlxVHYEB     400     140��gޅI��X��sh�[�QcX�\��T]FM�r9�.՜�a��T�9^%��~�����v�
�Fx�c� ��{kœM3{>��ظ���m_k'�����_��E���g��+M�>�E�t��O�t����;��G����Pq-�·�e֫[����Cl�EZ�b	�b̔�]h�*�R�"���W7s4k�,��p��EHם
�i��Z�� >����)b��a�r�yJ �
A��T��H�FZx@�X�(a���F���c_�Y�1T���5U�����sVF��'��%��'���-z$#x!J_��18����J��E�XlxVHYEB     400     120�{�z�:f��ɫ�~q+����*14�'~a�xԦ*R����%���݅�$K�{��s��}���
H�Ia�!{B4a�T��z\�`|�bO6����M������˧��bt�&_��O'�W�/q�X>�"�d�N2�H�m8��|q��A�W&��ӱ���#D�N�R�,xe?8�{8Cv�a2�7փ55�TJ�s���?�-�}�Lc@\1o��,%��<����@�:���� 6���mη#tO`+8����,��C-A�F��LlВ6w�9���1XlxVHYEB     400     130x�aE�P!���tz&��[���l4V�RT>!�_䗴�:�@�.��͝;�{�d�9��;�;]Q`3�Ih��,~�N�����!�J;ʉ�l�A�{�,ʊ��ɊB� 7��/D�� \�����m.<x��:&�(D	;�����]��Ћ�B��|N�9�.���D[4��B�Ӊ�+G����و`����~�����+��6j����Fy	"2"��P�\��x��B5i����?:��p��P0}��h��6S^��tQ��pV�
��~����`0F��I���pd-�*N�;x�XlxVHYEB     400     1307���X�\��jێ��o.y��j��-��Р^8�U����� ���RԘ�H��;\Z��8��֨�'Bk�-XA�>����I�;Y����IN�K�,���b�o��l=8�K�����r*Q�^`�eXu51���x�q�`N�̰�`{�Z��G*
X�y
�A�C̭Λ�kFi]tڔ�|�]�b���D��Z�=Jl?A2��KK�?1�T
��գ�u��
�o�]�=�#�T���r0�7��=��)>Z��(
�y�(�V���>���\Z��d���F��xZt���!��`¡	�*�X�2�XlxVHYEB     400     1402	��+��o<
3�D���D��k�t�(� ���$��УȲ'�)�/\�$UD	��ގ|��Tf�ҟ�;���`��,>pz��s5b}�"	6�	8���\p�<*��K'E���X���_(h,���)Al�I/'��ضjg�|ὲ�9/R$�@5�+o餵�%�Q�DZ�.���mB��L���J�2V���������/�����pn�K4!�������B	����Q+�9Hx�W����1hԔ�9���7���<�a�&��/v��G�p^���t������Ԃ�� ��{�c����z�	���@�}N-ϧ@�ś��XlxVHYEB     400     160U:]�Ȓv�#���
�%]����Y�	����R�$;��Y/�ܧG$��+��@��	�實��Vg�'D�6X'^�+���o�M�q���C���{�e����P)�^�'��~B��uE�[w��vv�7�}M�����ܢoe�3�����@[Y�s�7v����~�/��P��2W��3�aV�]�_	�tvv�Q����Cղ���a�EG�����Vܣr����I�<��xSK��M��q�.R�Z��K�NV��� Q�+d���.�_��U ��Z-P7Y�<AQ����n:צ/����j�сe&���h�$�}4b���ځ�������<q��1Jg(�"+��DYR}�XlxVHYEB     400     100.���7�#�"V
|DVj���8,�u"�:
��|�d�*�cM�^�;|K��.�ޮZ�/s`E�ߒ��c��|���R u,�
KI�X7�����i�2�k^���(���R�L!��(К����E%�[:�I�:�#;�h2�����φ��v/�r;HT�r�cUP���F��e�"��Y��or��v���>��\�3!c�yo��=��[�<��|띹Xᴍ�|���u
D����ϭ\�I�c]��.e�����XlxVHYEB     400     150?Y	 g1��G�5�~a�xv�c ���:��l\*풦Z׳�n�n���@2��芺C�h=r(7W
x�#G�f4%��67�l��Y3"tg
MU�~�1w�\��?:��8��"f��iTG����J�i��<��(�'���`B�@��7��;;@�S�O
R��9��AG#�^�:�L�C����t�t��kj��6�xHB���#�J���S98dP��{�H�AJ;�&�!�������ɴ��5l�m��8]��xC�����&���m�� ���z����6�'��nX��/<|k�8j!�������"g]p���L�uҜ%�XlxVHYEB     400     120$(p�!y`�1����ݘSЅ�[W�.�-}�%'=�gZ��MW?��S.��-��fsJ����`pD6Lg�u���T���(�r����)��	�n�)�Wx>���SA�F�Q�Bb��@�&c����e�ud����j��==:oN�o��¸��ӕ�L�7K�	�}���w�ڂQ�!e^�.��-/c��j��t	��̆^���� ��Q�ϭ�Q�Q���(� �G�������/�z�k�������j@�|�?����8[�����'*�N)��}�+xXlxVHYEB     400     130ym��ϛ9�*h���V��Y8`X���r��+%��)���ī��p�Y%�ݭR�<�օ��Z�n}
J�=SNJ�5��"[��T�g��#>��ߵZ���6�MNa9�1�s���E9ny�A&���=��@t�^K�̴tA�!?4�Q{�Cdw�\�����J8#}�9�}<]����t���s�{���f<E��䜍�E2&�~;�	w;�iϸ+�k����!�{Qq����YcE�*�{�2�4��V�DO��
$� 	I�!�ur�x���ރ�}A��,�8����J���Иse�I�[^�`hƒȈz�8��f5XlxVHYEB     400     120���V�7_`���Cf3{�����ȇr&��"��[��y2j�[���%YoT1~ͧ[;���p������x�H�7�y5�jD�hE��t篜�^)�(g�Y�����F>8�AQ��+)r�r���h̥ݳv�Y��MW����!�pS�K�Ņ��*��t墆&؏S����C�UuT�y�,V�W�r�W��e%}��#�v�7$�ެ<r�B`Q���uBR�z,oBT؍�|�x�6��0�&�W�3ŗ�7	z�ԉ�7�ԝ�I�2�EZb�H�]1�~�K�QEM3XlxVHYEB     400     140�ݡ�5hM�����*��m�ӭC��(�k�d��r�f4Q�,�TQi�op�	j�rC�Kt��ɾ@��z.n���?���
װ�~�6��`�d��DW�c�?��+Vg. {*�q�}�qb������8�:��Y�p�}���/�9IV�o1�\���+q5�k&~!�i�1.��Ν|�U��Z�oe/�H��������(�5�F_/b�⧽s�1��+	�
>����\�3���eІ���&JX�N�
\�@�,l������J�O���tTTBȋ�=~�9�����I.�f�r����HHT�;XlxVHYEB     400     140�|)oLh�'���v���U���eg[�[�Tv���HOͰ��`ۉfd�)�8�
v�@�)�	hh�b�&��l���?Tuwm�Κx6�~A'��<$�Rco�Yf���\��?R�k`���R6�Ob� ����p�j3�� ��m>�ܔ�R��Z<�2	�g��C^��$�C!�����]�D��x�D��G!32o����EA���H��!�>��'.z�r��י�&_�[u�PtV�U���;�F]q_+���'�c�Y\�%����4�����/(���Dg�7��B
2���i_�����{�u�gL���2��XlxVHYEB     400     120P�*m�� $�>M������k��!r5(���d�3�d��v��O�� N�DtrZ�U���K�(0&����9����8����1ϣ*S ����,tL��.ǣ�F�"	�`�T�u|.8���ӟ$� =h��Y���l�g8n�"%��41qQ�}XKL�����ףZ9׻��f=~�bar�Ѳ'��:�n���Qϯ&�`���-CU�&�"��e�*� /�?�FGT�϶��A�`y:�����X¸�<�A�4 CQ�4s4?� ��I�����AHO� �U�XlxVHYEB     400     140.��N!u�G]�%+�w�Zj �i��ϱ
���P� >�:�1���~�J֎�L��po&�e�T�5��EV�[C�ԉ�u��k�]N޵:�ꚙ���O#RB�`5�R�~���� �A�/�9ǜ�D��%���j?ڹ�\��V�^�"�؄����u�m��2,�n�>갅v�0�YXQ�|&�ȕ��Ú����
ݜYI4A�	]e	mT��U���rҗ���;QY�'Wm灿u�=�a�� c$��� ��r4Űw�>��~�L��e8�L���a��Y���_�Ae!�<I˦��E�YW�\�%ʼiK�XlxVHYEB     400     130A^�4��11 ©��h�����c��1�hp
m � <x��u5����)�"BZ;�{��t��>D�<u�by|�k,�&Y`w�����!���'�K	���S- �MZoB���S@����u��ᶶ��}9����B�r�� �e�}U���?��'����d��n�2��lwl�z�<��X�YU��xb(:�k�i�$d����� AJ���}��V�l�ɭ%W
�|�L�V�j'?����:�|#
��1<��V��룼�Kl
�G�;�hi�܌k٧�D��+#SaJ�H��CXlxVHYEB     400     160�7��m�ȤW!eC� �M��dS�"j��HFfo[/��CO��E�#��ň������rR84�K�5ד�pTi*I�c�%�����y �/���*�V��Z8II,��O�1��"����AaB�����8�k<�UAOKG�P'u���~��|Y�S2} <1�"VxCT�%�H��	���+4�Q0Y��q��STM[��ZěD|ٞj�L��K-�aX^�
�YnS����80��ڕ
*���5���ۊ�P�{�h��`��
M����c��-�4�t��w��By>
d�2������<`>�����}yh�>'mv��4f"��.s&��BM4���[D��L�߻�����YԎ�MXlxVHYEB     400      e0u�r�t���;�C�9�8i�=��cO�щ�i����V�a��&���~U=���&%ĭk��14+U�����<+.�S���$a�A�b�w�hֱَ�s�H�p]i ����?���/�{��R��$��Ey�͐���x����B�|v����M-)��m ~S& ��r� ��N
��*�K�z~ �g�T͉]~t�E5�Q�
=���:���[XlxVHYEB     400     150TAE��G�k\�Ƕ�*�u��1�h����)�^��	��|�w��C��Xh�
J.�*��	@�iv��Y��gS�Nl5�Z�-Z)�(^ Y� _ө����0/�jP8�����"�
i��\���ެ)�=���J8���ć��r�K�>8��X�����X*�Ҫ�"z6��҄�\Vn�vA���p>9��p:�P3Q�l�U������DI���&�ex�A��-��b�����p��ͯw���l]�	k���3[�(���H��\}ST�z)rOA�*�m�� �r��6�c�<C2څZ©�C�I�pUyu��?Xѯ`#XlxVHYEB     400     160�@-�<�c.n�3�{?)l�FLH��'��&����f�����ٷ�����M=��H��Z5�Z�ؾ��;w8���N���"�_���S�4��s��7&;�n��H5T�`5lWP`�e�Z��t�J�+`W�:�� C�I^T�9&�v]����a29q�D@�wE����4��SWo�bǢ�,��7�~w�f����R1���%�}�$z�{�F	B�p�݀���i�h1q@��<�q�����)�Li~�K��\��q���n�{�Ʊ$~��LK�iT�	2wk��,��@��ʠ�`-�~�v�H_�{|g'^��<���ݾ��?5�Ql��_"a��"0l�XlxVHYEB     400     120P�*m�� $�>M����׷�x��r�N<��T����az�*6�aNΜ� ?X�&Hl�K@T�P֦�ϱP>ř5���&���Z��m��
M�Dcl��R%���2�=6��8����sX)t,��	�>M��*.���ܖ�{_���v>X�)������x��6��H�
n�X׊�[�J��g=-���/-ޤ�o��8s<�S�V��OO����>MpLH��=������('�n|޿���>2Bp�h���oe`���
���O�/SI���4#����~����=�~��XlxVHYEB     400     130E��q���I3ߋ�ef�Z��3�$�	�T#�q�]
O�H��ӷ�#����p��Cq�?3�l:�dQ�A��׵�U,� ��;t���ч
z�����N��D���~L�:@gv6 rxF*�w��&��(�|d�݊�oY�K����~�FY��p���IQ���8���bt�&�dtչ�d��~sn�i񰅷7e!4'VP�2� �.S�Kl�>�z��"Q�\��d �8y�b�T�M��d��L��d��J��;�����x��:�2����ᨠ��YA͗DH�|�:��Shz�4Jփ�XlxVHYEB     400     140+;�P����q~���1�J"�xT��)g�/K #"�'����.��v�ΫPV:��Zs����fEtGتD�ٻ�@��;0�)����.M�ߝ7�C��
�bQ��d>����h��F��8z2[�>�Z�?N�Ɛ�QjmȖ�H~�.f �̃{�Y��{K܉1X2��N�=keJK�i�[,V����b@4 ɬ�z��גG�nk�#?\�	t�Z�9[�>��QJlq��]g�ѯl�}rh��сq��
��|FsW|x~��JF)���C�5;�����0�0�4����g�'�,�������?�t�|�7� �aG�ߗ�Ż``	XlxVHYEB     400     160C(��Rj���-=r�ώ��a;�U��c���Ӵk�1�, Y+f���X�xwZ��+��ꡞ�.����bƜ�K+ho�|^L~<�I�)^;A�$�x�� �ϲ�#�Qt|mA�oE��gUc8>�GUw6��J����2����cbQ�FL8
i�<f��э�2u�XN3{2Ai}YyN17�;B����ԝ��"�,m#ӆ	�c�1o�����������sn]䔝��aJa$[��j~��?�3E�jȢ�e����Ot��g ��JP��c\EI�1Dtˉ8�b���smJF��� �7E�n�h��Q�Yƺ��\~^�f�����Q�jh_�3"��ZB��q��$3Y�XlxVHYEB     400      e0�U�W���MZ�Px�Ѫ�tu�%�;��t!M]�̏ o���a���xN\!�s	�-�H�r��+�\�$�W�C�$�
�^�7QXL��c{����w|��b�Q�kV�"42��x�cW.S!��|f\�5�� ʒ��=G^jct�~� e'��*�7"���v+�5�'c=?���k�0�ў����N'��6��ڌ,�hu���?��}ܐzE6���XlxVHYEB     400     170�L��k�Z���]@���y����y����.
q�:YL��`aɏX��c��~�*w�6NB.����q���^Eb26�U�2W�����-a� ���j�ܭ\�`��x���[￮�H�,�]S�y�O�P=ɢ��+6U�:i�͗���)i[aM��D|N��oɢ��(���}U�̴���@��U�b�OݬL�
4�';v�nn+���$���)�ug_L���S؉k&!]�����%�ykO�����+l�/�ݬ�����%�������9*�Ǽ�"��=�'�z5��'�x��I��ܥ;�t{��8?(�Q;Ą��R\�-�7�
N���L�1CB"���eԉ�%S�u*e��?P4�XlxVHYEB     400     150l��1q=�3���fo_��U#��
JȠ��mKSBN�O�S����86
�C&�!�i�1�i҂���7I�0G���X^\�=_K��һ?�K��͈)j;��Q��RnPiW�Ŷ�������{s��6�6f?h5K�x�����ڲ�_�FǄλ����i��1t4��!gΡ��8�}����^��[
Hi(F��TQ�g�ȃL���｝ӰS�4��.���HFY@ީj�ֳ���r��:�)᎒�G���xAal��sv�.�� 5(~�.��Y� fd��
YE=�t������BR�H�irgE�����ə�_%hU#��փXlxVHYEB     400     130����l�卝ǅ�
����
H��;tC{,�K�#b���8����*�Z�S]����]#&׬k��g����o�7��]�8־�T�rÉƄ&0�r���/�k�e�C�`K�"��K>��K�/MU���f���7��'׾۝vv$m/)0��t%���~1��� �i���7bY�6Dy�����9t��ٚV,\��v�&�8��ɝJ��%
I@1D්���fPxJP���������:U/=?�f|g{G�k���҉R�[{��?Z(�/8�q��F$b��b�b8���?a�UB'�XlxVHYEB     400     130��_�=��:w��nd�D�-u�.�v#����K��t�CT&__.ҏ52*G�q����!O��%a.џ9��Vn��C���~��YR�	�i���xUh����#>��l*�H\���s<���?���!��<�l�o��M��	U	5��!_�^ծ��M���1-��Pm�����wC�1h�����ů�|�A~��vXJ�#�ՙX@Qi��½�uoʪ�v���o�oނZ޺���Ԣ�< :'��\�l�g'�5�>���r�gF��t��<�NU*
��Q��}�L�V���)�XlxVHYEB     1b3      e0b�����x�x��c�� ���()59�qڽ
&۳�_���ǁ�J&�qc˶�S��1Q.����0���xID��M�E`jKޟX�6�K���^���� �`�)[��s�1a[�m`�saࣽ5\e��W���W�비X~��$��jy��8�ET�l�|���|�ދ��T���*�O�5{�+`\��x���4k�W+���j@T���kkki�Ş���?�Df@�