`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6416)
`protect data_block
0USWSUGxovGsyBJteYpEoQaa2n1c/ocEqDLqgCm0eLOiCHivf0SVmqYH3O0tgCHdrY04Lpz/KbFV
bHu1+CiJGpSGPyB0hGwN5Y9FxvaVZEoK7xBUNuAEEvZrF2i4ZKUCqv9te2tLGzbdkCyeAjrljKga
209+CIlEzOUYMdK58P10v7DxJDEXtEku38AR3gqivT3ue/GbSTr9mlKOfGahXmKyI7bK9DcZLhYv
aWKokdqYObFFTHxzk90UhdWnJ3p4WbGeskP8CyXfjdhahRZjeMuyopvIXaV2XEr+D89KAVoqP2wg
GqFy4P1i2AwbQnV9WEu2fQBcA3QUCV2YsbebzgeoXxNvXdg/rl399CGbPW6A0BglMfTtgfKidLG+
xwxCa2wNHUWhh4xcpMAKyMb4yHsxUX1kKXco96kbJMCSb7m6uxKyHgRKJG1SOAyu8qAjkX0GuW0g
YS5r/nD22zKovLAKrPwnEG6qCUNbm7uZDq6Pd/dv9KDFZ/Y+F24s4kZEXtwI/FzOOjuUOonjeNsI
W/W4U4artFpZqrTEdE2ALjSLaBTfCjQbJAz1shiO7x0ZP666EUlF9lj0Ue3fLI3qs4sS6B/cjvw/
JWwdpAKFGGllo64NMYTxRd8he9QGf9P2D9qZG6Adyb1mdZqSFgdpZXFVOjnCDJcu+RdOCQtfe3xZ
GKhCp6aE3ajMz7amQhhlTvpVMR5VLUe4R1+IydCeUHh6n5SXUPTn0J2+8rAzcaguQAFyhjslCrZ6
o3ldAyp1vAt2JNUqA+3Nf0TFfgvQa1NgyI5KNSdUG80m4CJLl9TiDA/FPb7BFsgAQyb88HVMPTSH
8UBtQoR+Dz1HNxvXjop2aOl4bpW7wcbMCp7fDmlSnGvhV3QIvIIOUJr81NkBiOAmcThq8n46eWgB
a6oReY2svthBfAW+GfNii6AHyrQ7hmw1sWn8DoRIqfPrysdcAzIvFBVAZ2qwvUFk1rlD8xLhkzf6
lnVsZl+NqT3IB+YOjuhx4z3uQDox+22JyUaH6Ad317n5UAN+3cCuGjmuIm6o52y/c6Jou1kJv8Sb
z070ca/0ZifQ9MB9Bpm2l5h6i31ESoTUh4ABnW5TGKlMaRpHKAoEdlqgPIPnjj215esfLHyrxT//
JmnR6a692FTaA9OXvJSN+JQwO4lxySYDmDFFjhv/ie3S38sVBh7iF3aco4KsDtg/UZCDVqTzDW/D
PAIBSdyBRZ5R7fa42bOXfQaasWUjfomZcKMwGGFVLzMHyf7KSt7jLYXYIyWbnoBSkcwL32ljj+8G
QBVqrJpXrr6s4QRtAM4Ixv08HUNhCMbI3MAZjOH9EgHuSsRU24qtIow5CsNrJiKiFEDoPuC/K6UI
nM0einzAILTA8dtUh9fcZV6ORwyJQBKDush4btoIpph4dh0BOiPVJVdhiEpXYkvKjGJ7SRzChpN5
6HDnWOhv9zMNvH36Ab4FCQUBoLht+LQxCSkoANzNRtYZM+X/L820miIdrQH/SlbAjBS6LiJrBNPJ
Id7OHg6J2stjI55yoef73XW8JbTJtc7hwpHDfWaS6VGZglRttTWCozWT1hxw2kK3p6LwN/u0J2RC
iy7XBiXqA+hOK2+9kL0z1ZrZEpWKaN0Obo7QfDEuPI6X0+6tEMYZ0c10EM5D4BfBMAPMfjf4QYnr
qd7aCJVHw7KdKH/P7nHXrPW3vK3lB6xL6x1RYazVdr53tUCpabkBkm6uuFkoaEHjJANRMejsRBtW
C4ol4jAxUuj2huKxoPuJvI/XT3GRwcjxXta93KEBAYWAsRteHE7eqe/qAyegX5W45NqQo6iGNn8M
UvRnQUbNpb7BwaWoMC8wUMyVGylVqtdelizTmg9sXYwpEe4VW+c8k+xFhacWJFEXH9DtHzR3eUFE
3JnWzwBCQCCfuzflGBojdM1U9BeV+9R3WPv+2btjrAOmtXU/h7IPLmCsqKJ4jimAnw6W+eovh2Fy
VjX+2KHoBxIDBv+OI67eirrcV1z8V4GmnYfFTqUoKV+ksQ0DTTlgXIZHSnkCjRfaojDBGwWdvfqj
wrfhPbiULl0ID8H5yvUFaJcpN9GQP8LWoVtTLcIPUE/ChPAZ53USlFmNt5an590FnAjjK7UOSdwa
ZutNW2ZUeHqPH2hSP6/V8DvjoKWKpQOnPboXG024bI9jkBZJ6IApIoqQfLXxjjLZ8hHDvpHglCcM
EohG3PYluxEWuIHRGhFvTNsDQkHo67R7MkRw8E/DF+ta3AEmfcSorGiAoa/PFusSZeZjZaGn8PRE
+C2nXutDK02RwrARlCwy4lAIE8U4tcPQ0leqYv6cr1jAHSmKpNRy4UwrUDzeG44bYu+pKcMfmZH1
tOXMqcZcJL2X0EO0RdtVbKx86CRe/SIIO+G+sT+3ycdLy1oZvtOG/m4VZC67kCLl9umupKAUmoI1
ogzWuLUUUi/Loux6m5w5YYe0K6T4r5M2Y1Wl1+357TdtRZyiiTLF5yDAu9otN1D8a/sK41Nkr90A
/v6ZdvWh9BD0KRzAQPiI7k1ppbYy3OSld+TCd+VUl3FudbkTRkXoEcS0W+9zd8QsJl6poDDw7WpH
wEWFDZ3D5sM/3ifgxSOQsOoooG5BRWiDflHJRCntlCElseLgC3gw7/J9tT74DQgwEPDrcbfYqVDE
ST7o880aAybiyRTEBkuAD9m82p7vi8mUJZJ7IkvkRnPm75DQmMDkJIYvEM1Y3willtFZdYiAgfvq
70HJ7OWY/Dxpn/3WC0drVmtRUN9ejVmOS+HgZ/qJnYns233TsQGZtd8k+y+cOkdg7ToXSNpqKKNl
T6aAiJPCA571wzXZxWLZa5kgUu63Xp5gsnZOQ0omkZtag9wJMTQEAY57fuuUC34fdTapMS5mqUx6
iLiKnvge1lu7S1IZGWDG+bhnzxaduD3CvXd0glnX7KfPHOFNQ+GhgYffRXt9FQqC4BwtkEM+4uDZ
QDj7McCjbTVKIdDgDRKA68pnQEHZ03TtzuSpUHnk3ujoQM14sRxAXBiSglqKYoaWZeXdILYHaZGV
SZFT/iFH7RW8NjbszAszOzYOp3kzpdZcPyvVSjPCLSr5UwkzS06l5/LNCLok4XJjPLjt4GUZUgWt
sQWSsQx6rXWICKB+S90o+hqz1vLcGs7dRZPC3pIZh6AnuN1R7+JgERY64YSi9x7AELkjFLNtUMvC
zDjAN7ypdpH8bWyDPP9ytMjrJDdQbHBMYGkVG+IKpIbruYeW53rdhTajZaapg5/xvMgBaa7cC6ue
UoVLz9Gwg/Y8z68bqmtxtIHncjqAXSYJlCpCvV8jSkc08MGJBkh50UJ6Poanr0wjcGNju4/eQ1Ga
bs8KaKITuFle6IGHUmEESSi+4bRPVN2GMZerpol4LriPDaudE5LBm7uq9DfEWli8BSrgty5ay/Ov
WzBbTBuvd7ERSgjKXCEe1aiPHXjvL2FnW7zBQTbedDO7W4QfiPBedMK7fwVCNAW/A8LGq6SMcxL9
ZFzoyu7dAIDFWMjBaURk26dhaXsW8UcI2Ufrots4mKBVeu9MCcQd2nNj/09tdfW680U2ejDF1teP
JwaE8WblQoXX2qd5bXqo7qakYy4bezzrCKMQAG6nsRGxWqw7JWhMc57iyPzkFLjjS8DEe27DJqRP
uQuoX73cd3UoBv3bLxpNofCIJVWFuUkDQvh95/mT1AGL+M6e5eZrbor2NnR6dO/deiTrIz3p8SLF
QKQOZpLarcNL7QSBbnG+zuQcCsVvn2icO77jhve+ynIsUdQko8EdtIGYn7S7KvVphxJHH3kC9OYZ
l5sXhbphR2pszzZPmCDJHquAWF5KMTY5jnHisi1Rb7k0ca2MYrVgW8/SxsgPeJMdUfEy0+ig01QS
FN1Awieboox0l+Q5oyUQEiDvEOp/fbVxJnuTPOz5DabLmwUSA+nJvECGt+vxqYrDshEBiopEEGTY
Q2cPbPU7snCWaRax1g/6iG5FyUmco4eH4p7nZX5fw/2YSIWpRpenN0MfaWGBsjGnBOOWBuGu6jin
0tdxoWs4iRTdpZawMY/Gfu0jeUJmYP7J1oTQY1mDvJGZjrF/AbDla4gCtCj19G3doyIujZcMd1IZ
bCvcsh/iqNpXODBcUR4ssC9wL2qq3quWbj1UbAOfHEWHbs5kuPXwzRm7yAduLOGyEwpyb3NpDe2I
D/ZeepXv2Ctw6qeS1TiHnzIsuXNpqpQ0KrwcdyMWMQ8u+vSqCeIU6prjI/84o20+SFQ1fObbxKjj
yHjh0ZdZBFCAVuC2xLYdjzhVGHvTAYYaoKSTen0ltihkncjjB3XnCeVHCV9i7mqL90crpFoo6Qiq
4ybuma+B0kHvNezqklAi0pSTWHRSAIOuJLiJ2EUEI9Vd41XjyQKk6WB+Yw7xqxVufhcY7YTagnjw
VxbfadjLykOjEq+gYTanj+v7EbSIuouzF3GOItkG2+Ghazi5/3VGpq1g8p52gYBGUDXhDh0RPdHc
NtGPyJ3ueNzKCUHz/s6k/X9h/zKw0dcTLpArU978cgAVSgfq35uGLftJ7dWH7ERGv6yCZ84poCDU
CQ1zBUe/lwg//yuUD7cGZqWWgfC2B+AxQregwt/N5Z+OOw2QbgPNgVyXTR+6VARVv+Egct8SerJr
zlyDScAby+8lQNyTb79XwRCmzuGoQy0yhfCVsf+zrbEiuRwGeQ31mLtVReYJpwflbY/6YxhBSnIC
FtmTIgLzH903P+pw0UCMQiX+OiwfZhgmVbY9Ww8Cu/R35Wa6PSwpVtkh3Avn11CAaIjpTo4brPXx
mQttLjvZiv+6jGBjsTzW1kAR8WqTT0xC49+Q6nkKkNFznundPx27Rkg3oSpRFR3NwDQB8hXpdVZB
VKUFAVXGnT2Hk/JHNoCkEo7ibkLWAkACOKy3LD52tOp3V3l7O4e4v+atzKm7JxHfbie3kJkaW+b9
9E97CvGP5vL9P/RpKTb/DO86VeO3BQfEhetncDrmfROCoV+jzW3ubHnaKXQLrtoYYCw+tubusdV+
XSzGlxqsygrjJJPAtPiWpuzKGMZyZgyfqpB3lAXgN917mSJEK/+c1ATNr2WHq/VSVFTpdax56peE
3gdkb8l6yELZu42JfZ41SC38DSQrlCz+S6vBX94O/xnlWOhAJnZhwl6fQJ9N3NkCRbiObXZOklse
MzRHYXIDAUGaciZX/KicHJ6UtAZ2GrfqZEk/RRVWmEKPRhVp90PlQA/9fS1Pp2SrMf6iQfNBe9yY
OLdcjNZmcoB/wO9Vfq+2+0VoWm82WPfOBXgpksrN7opUo4TpHpGNmXoiJ54TzMiAu4R7lp98nEtQ
egefrXLW0WQIAn3EBNDCXFOpDRF9Nq7f8jWOmlguuJe3jAmSXLUEl2qq7B28xnrEGbU2kae5avIA
DzcKtq8sl1Bx8DxJnhdGsfeFnGBWGQ+5lDv72zqgANYhjFctFFk8rrOcmGg07J533K5PfqfwdioD
K1h992qUQAMmu8rj3Uf3cuUeDNFN2nigA3XdWyMyic0PkqWctIM16ZF7o/NqZYUrHLeu6zY/OGM8
yaB4lYA2x659fpLVM+yBhJIWguYvHpRmPtf9YoImcGcozmnvqbiJFS9ZFEA65lmp5+gHLFxFEJ3x
MW/v2fvbgtIkepGc1m5V2+wwLg8SFw7HgSAZ2mepPIXNna9u71Dg2dhfX/3ok6AVt9vinFDFJJST
kBYKdKU6bHLcDMuYdjx/U/s1LvoE8iE0JzsL3D0sdZ9S9pZYmh/OpBzebIrUmHEv//9VBs7agfub
Pdz3D4Gd+qOfyRzms/BZyE3jTJ3FdkW2xHkgNtCMFRiji/1WGGRrlqwydTlg5a83tAzA9HqteffX
dnmIPRzDRpTME5AZxxik8n+5PkUf1hW4y9cLgaRro4GPkLEWDZV6uRCU2x/ZEcUT0Q0bzt+59zUE
YlqJ//axTHor3Zdq6CwOJXr7j71BxlBC/3XUb8joP+hIiQIaCUNrs8igL2FutMQmi/9nHt6TkYQc
ZCCqjnld3sJLOwCAe72mnushjt4nXgIQjF96eHpL9ScIaxRYieLCyF8r/NNOGd2OGWaSQuM0++ra
kkqXITZqSo2rVuBqnrqNsTG9nG8/jmJfbjL2Y6r31icABHDTXmQvWoetGD1xyQ2XjldlM7KDmUnN
QFore2qigUf6lQwaNEbbyuJlEAaUSI8Dfl0LeFfsq3yYkJ/FHCRREGE7pGS98Wc2xkZVpMGE2bfX
viYKFsJaFcuX8fXlWSCkQrAhU1ahiRaI+6b9YhtN/zEdWNJuIChZjgcPcPp0Bamwir+1dovgsb7n
4fM4kiHNfEAGrDzzOl/Vn27xClRY1ReYLrXJBl87McwF9WXn4J06W7rCnxFlPDvDFPUUfQbudaG9
WDGkUqAnhAJ2qJJDAWo1yDcr4r50rHydXYp3WPu0xoaNG7GeH6zfj+L3l63UAjsSvaiHAqSCA/NE
SUR4vOF+A6pFwTr25f4lD6E5VhTmxMpJB27dvwcj3Y079uUPp0wIM0Qh69dXicsZ/CUBJgrnXyh1
QFXXwvZPfTy/9Lca5G+iZBUhtO/aAIlCTOOaZmhVmSYsam1HNLbDhm4eIhQyZoPxPzO88Qu9Qa1Q
CuDBIGpHqG8oPXtC3n8lT1Y//rLFeeuResUu9k6q0RLdKXTYQdc4DyYRYP1+gZphBA7MgQM9peMF
gMjZUPGuWvlfbagknZmbQEvCUH6VaFWTCtL7heLlj7rkx98aNMPLQYgtvmxNTkWZdcIcwPX4Gh4b
GaGu+nG5kUZrMOS6uvYUcPrlfs/QjnC4ef+3yLcgZX77rjGsJAoYDtJm6DE91JiOho1EE7END8nd
PoYCZxDdm9nE3xOQ82ykuyIQbk28k52ZWwJ6MQhjDzwh8/MRCgTvJset14H4estA+xTeImH5xyhD
y+MIg5a4zXl2kije6gIucFSbXoQ12XkGfDWqpMelbKuz+yNRegs2WoqLgcg9lCpD1fe3vBz18YC9
QdTvJJVcqLdBqlQqXmm635C8PGW6/BYOkN1+daZ/N8JjqwA5OKxZ43Caq8mvquBlxgB6fTczWrhV
//kK6UvMgJxGKXGfYz/w6cN/W+pjrgTwinB/utLmv56g1S1dMXzI72ttYuMv3PjIcB7F2jF+ToE2
hIrzKp/e74+IXZhiLsA5yp31tqx2mzUiUEbgQwCKR8dSApIFqI4MoeJ/y0VUOZ8CX4MMwZzRD8NV
A4nZcgNf8aO0eSTR3CCKaowdlhvKEiBkiWuzbPsTqEyQmS6VA2TK0xiuoPEsNnoCg1z9ajYYB1tU
VhCf5WMGjpNq5/wYcDBOUq42SWJ/90sX/j0Qe/R42NXL1vjTqhM+Pj3EBZkmMa3AsNIIcwS6imG9
G27Soj4Ka0W/mp+GpMPs4YB5o3W3Sajvpow+WvotNPPyz1N4RbhrMUYteUfBVI0AKfYIbtLSYyzv
892iA/PcES0moHby6xWbq9t+aSQ7Dr7aZYSqtfn3bhS0/bieiyfeJn3u17fUDcsJ/lv5ivzOXh8b
Jm2+9XJVvCOd4bYSFUaKzDhoo/0YqdayMs9YWkQTHrsg0Oje2FnC1BH2ibc2yiJCyOC34jBJyGws
X0XyK7O7bJFZ2ElqcDkqzJcHa2+4+esMtdO+NSLN4tSqzW9ZMgFw4cit0/mRo9hMYQWRDsb4Yb0k
ydNRuNInyhbjqut0xiB1sS/qQMQGKx6wDOgfS+6bQ3KNTTUSrzp2nxVdZoPf99ikS+/6qW0SiM/Q
VLPGuGsGNGaBhjy469U9O4C5S/eK+rMrb9a+aemrqfwg8Qhqd5Ct1EGluBKEfFxGkk2UZk8qOpJI
6ZxJ9KDJnEXwAsiA8w8Pm5waNCm+LJsxN0DIbQ9a6kGC5ufaSjYScUPDyf7QDE7TqC1F4y6MARQx
bwceNH+8T+EMw7ZdkiuPfT22EB9KhrqJxvCHgrEcSexU8c+GYZ2zxxcXtNvwUKafumYX+oRF7HL2
B64oUmJiuRuLuMKMtJLzMyyayR7LvKP2y6CVYiYCwZFo/mtTS3vq+Ic8t8BjC9nTXsWD6hMumPpK
ZFDxTrPx6iYH9izCht9bzqgcJZ4aY/WndY3IvJUp7V1cT70ISyNGQ7z9mlm9QjthpWMtlx6gVfXd
i1uEsO7bjHuBmKruGNLCZRthNrnD2L/Uxj4am4qwC71sFO58YurDQujoNGVNO1ojr+wfgw/8io1z
chgMx9qvPB/fnRDD2yKAFJuZcZY/1YrUm12lU6gyvHUGitiaru/VXMgsrUiBjHx7FrBn+jJKqMue
A/biQt4lDgqP/z/BjE0Eulmn48q5b2YbFpbOuVKNJPpOxMMmqirUT1+0jjYsunNjv07JA4rBp29x
p5ok5UTCNRbboOpUXTs7fOG18fMO/+iEhnDqnMvYClOmWlp1YwLcE6FopmrNDAFsu9wmwNYroGhn
gSTzQhQEOZGg8LT/vly5ZXHWfoum8Fcd01BtFtbdf8DaJQrpqjgmJ0RVF1rg9r+kYNYgOIV/nnTj
y0JZCwURDhu81OOVTUt1B9NMqAZmzeA0FWuiGytacMI=
`protect end_protected
