XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��;�M)+o����m��9�a���.&U��d���K�
�e��$���7=+>����'�����R$w+��c��t�F�����ZC��q��R��M� ���5���*L�ü��G�^��1{u�Ƈ.k�g��W�G6�O\��i��0`�=��]�#��쮺�kf�k%�Ѝ�,�ߪ��'M�'�f]Ƣ/z�D�C�<O���r i����9����>~�����T������QR�5D͜4
Pv�j`�?:��8�nI��+3͍�#�i��	L~
�O���x[�XҔ���cZ� 4��)�/�!�GH�
��z��7�i8�VnFOI���O.������%{��AX҉-�}�W���!����"߷��tZ�j!g��J/]uN�9�9�_�n����w���>��	c/���w���Qr�Z~�(m��<(��Y#��{���q�c��	}6�b�,�_��M:n���j�얦{���{h ���4��WQ��g�%o�\�}��(N�`+�v�x����^�FO�%#k��U#��xp�m�v��N�F/E��J�`x#/t�mmt��4π�vaD�l��*��}Y҄ӛ�`���W/�;B{x��c�h���Fͽ��'i���M;�KA�}�=�je�Ń~Y�&t�e}=���@Q쵥����+��������1лU���$>u:����}W~��?������2ޑ������-�^�z����޲ڠ7)�\� ���XlxVHYEB     400     1e0U��U�-/(:�Bïd9FH~c9��uV�)�#�#1/���[�p�m~L���Yo�4��!'��˚��/RW`~<9g32Ox�aӛ˅��[Z�a�Ǯ���*l�X2�֯ZBs�ɜ�l��TNe�L/���8�f���/�**r��y�"�.�ݚ��2K�]o��#:G(�%.����^R�����I��&��EwMI^�oY�剘"�H�\�g�b�s�]6%��S@��.x�2�(�ZCd�3��3��F��W�h��y�!�6w>Jز��<^����QE�=�����y�+���~�UNs�M-�<����"��mc�l�|��٪��Z�A��9��0��U��^���H۱ >�RA�:ns�����1�i���!�������c[S~�iӲ<�]�g�mA��n&<O@[J5��	�1�Qݡ}!����[ ��(��� ��"�G��@�@���gd{�,�<���XlxVHYEB     213      b0ju����#\?��ӔX�!c�;�vb��d��,�t�!�� m7�?4��g�7��I`��~=X$	.|�i���{O�9y�f;�z��w�F2��_��-��cI.�A{":ݳδ1ۑӓ�X1:w�8�����(��խo� �9[��C�8!�ޤ��#Q[�P5�|d��/���Ò