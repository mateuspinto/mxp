`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3488)
`protect data_block
/4n95xVsF8z75Xbww/9bs1gotv7UnH8/PbTasiI/KXejOSgtoM8B7bzbRx0bjbjKb7cMobk5frQQ
RyUn7TBbXDGxk4kdTYXXnlqvWXFfGa3LCJAlQGaM5VrFIawnkLj80ogAJP8s9EVWLHxkZpq1F2S3
EHFU36Zfe+Subc9SYV2kTsUwyCA4TdwEulQtCPZnJh7qsH8mIm7XXrytCsuNjN3RfJZkqzpwrQB2
UFBVsToyUWb2U8QnfvcNSUX6JTdpJrQgRHWeEhcQCJJNT7H2ouQOHjqneZ3CGuOe4wjOfQzeUfoy
2yMI6ZriCOa7IFwjkzhajuB8Mw9a1miDGyJti385afPGvtxtJZE9QdhlXOSjAgseegFVgpYzSbwp
F1iWlH/XBuwhguPlyOrp233vGbvVbEScRTNASyPTC21UzRwbLPDWWXqOWANuxBiSGeaOM7wAN5ii
D+8XR1Nktz3lYZOk8GK+tK+kAqNPeu5Vw36lyNkdgEo1IJHcS2ufEfMzymP6FZ77dj/Oorx4Eo6E
UOra4LZVFPiu69crqaUTjAzhV4dtk922FwugLz1MNnv+Ykazy3t1eqI/DtPwABHYpFUPy5jn1GA9
U//kcixK1fq41H1JR08EsMztlYWPGIo+MFtUuZEO3mtBwUbJr258WBA8PMcI3Wl3vur6bt/OAVCL
9WbfJIwgPVXr9waYEqPrlI5WqrlAYX6yy4xgiqTpdxrEr4HCnLc/wrfxE4V1zx2fOE/i+ctAQV/l
vydQLvf6PBJxoeatbXOcuWmETTp1a2NY69llfthUYhQEzHVpUTds8Nvx0KHXBebFDAiTzjjenqfC
M0/AwjC7Tdn7UbSdO8xtP4njEq+0s7442ytfXp0DqMOXbPex6qRUfTyZnsFdr1QIeqoGqsIVAGMf
ExRGmmAxyftcdNeBCXOIBnJsWsEGeRs8COhcNMAr6Pw+oIcZX9UFn9y3sAaponHf9+0XqkLeehnA
Km2cpHIRBHzm4emQFoTmyJ6KlXirj7HB/xZe6Ldxt2Jsvle5SKKUbJG+/pV5Losy2LxuGWSXhwoS
sEpKe/GHAfg+gwgxdry6f5YQc9KeTitTu2G96IA7HczSABDGQvbUCrdRur/V+2HmFBrapV9sTSj/
cd65xfqwKP7soCBjko1I1/CGiOtECi+cn1PhYnkn/UxLCD2tVEuwZ7/ZobRVuv4hGmvjn+7Qxuuy
vJOVFPkxbea4PS8SiCJfZZE0m7wa1kmjKkYnAjTjWmNRROKZUSK8n3AyFYYnBYqoTbrRswhnyHMI
c1Q9nOAJBBcXrcEpsHQ2pyzrXt1xAURBIEBIikUAgLW7GS2lb6MwyHe1FZpfdzsM6/cCdnnIpHis
1dKNE6QV2/ML5FVINNf820QoRvIrucnpVFTHptVNnfv1O9OoOrHjnAEb9Dx3zrfa1j3iH6PpV04W
maGw9GSzWsSHif2gA/BsKenfKUhfZfwHfmaHXoZwVlIkGSJLYGSXfYMcAP3PLT4uXjd3bMdu+Xqu
a/ReWT5DX37+BDfO1ZSsbMc4IlJaLD30+w9Gmemln/9Hvzv6fKdO7kwXv76cDxGduZJxP8nomz5r
RndpdcivUlBy8L7uaSRfBeZa4upmp2Cl2MRZhMjda1yNSNssetocL+G/kw6EIDC1D7U+uezSrT6+
eLw+WwA//Je5qAIYwtvTRh+BYk5oAY36OyfnmMxRS1EJA+YBJvEAAxRfj+Q5F+8NJfJjFBqSChSr
NMkN5mBHCVjFfoOQpjaGLukk3LEAKStGGTh1n2bOTYnzXfy5V56AMynO3AstztC1GcIhPrBEoJnu
0J6x8Mq7d8KxRIhKca6eEc8HhfbIIsKlOG1Kv6ggiZiLc/UNJhWFVF77s9/mPpMdPIRJZZCuR/10
Hg2vDHkPQEwnmayo1fon3Um/rDRvkO9ZDCAlz1geh/WaffyYNoOIZMMpft6fWM+ni+xvvndUwU+c
o5Mx7ajGkYT7FrlSryQo/Rqylf3lBEXA9fj8kOjCRvLgzuAQQF2IMN1IKIBQEz1DYdvQIcfk93tl
iy1MNo8Hc2qEnWo7AKPq3QR5wNte9wv1GwmsPcUtY3yQVnAJcebfSiEsQ91dzV2HytSUIFAFfxtv
+n/vF6M4UkcEP8d/Gl59VI6sSQTGw5g9+yat6x6qe1Qk1PI+fiheYWXS/qYSIzUR36B5VdV3F+PW
4BOSiRPTz53v4atGtr1q/XGSzJ4qq56O/XnWOl4Vj44AjL4nYaLCCuu+K1Gi+a/NG657r6gbEq/b
CqfVxpcnvow30nhThciBYsXnkH3CUZ32PJehn9dOnGEEpejSOon3/Flp6jnpU4o8mlHLw0coaQh+
GezHr9XjK0RMKOMCONwNLtW3Dxb21GqyNfmP2J/wZQZzBAKMN/+6Zvhw8RhbAp534HqVCn0f4HOh
t3XIUOdmpITLzWDGaDRtP7jLNkc0iCmmTttyi1CO53FJXKK4DJd6vBQ3smwiAUxg8VtKOf8NCWZM
XEu7q2LaD3KtNQ2QxsmNUs47JpMBHHg3W8x289STVbQ8aDpw/IMXCvDhqNlT6nyKyKfPW3YMUOtN
e9UH7QCL89cY05u2lxwSMWUoyDxMkagsbZ5x7wnPnI3qvlc8pg/NmE6TVx6ZC/nTVp7K80xSHl3F
xVoxG2YnZTeX5DXka8hxh846AcC6RQjcY1s/hOgB9cZbogAqjgikdnGL2WKlKKS23yflMr4aIVM/
1ep9oEYtCwsuvV10CwGgrVprUcOCo2jMPvezjy1uX2JMmfIfbUCwqCo7jnryJdROzWI0G027Y3zW
IqYptFVryBVBIQl2NMS1nTK+jvAi/F2sDGscvSZGwUccvDIbHGZUjgvutnugUcCzYwWVt9wJaXNR
gye8GKrpYIcPB59gGbJKfKyZqPCqQ2L9sKPbmDm87EB9qNLF2dK+du1mGEeacQbVEqHyd02RqpBd
Rkb4iMAeIDQXNdGrMc8g2/XIrGfvIjy6ko0Y9AwFJMccPGS+FQswet7T019RoTqJrFsVP0c04Kwm
Hnv7VeUEHn0ULXcv0RGCbmPOIxk3DZlwCa46YcqN2GhUm2qvcxzhLXcrbFCQ1seZcRRwUUlEzy1V
X/CXHXNpi3cktZkGVXEbjNAptmu7im6eI2MJul+6wMXTDMtX9aha3UYMPjPYIbCwmWRofiCof1wp
Heq/FvYZjLgzlsnzl5As6QSa1W/XLf/IXsGhrtq8sFaXgCFeUE7ewk/F1kM+0M2NtFHRXN2MZo5Z
K5Mdbnd7nC8O3oinAp9YW7aCcUsmfnhFWborndYcG0az1PdAEggoYzSPKwWqUvY7VVnJbDukOmqf
zJgASZo1oMcqlcQYNqo7FQpY1AA/1ib437WIcG6H5+8eUYkr/ek8R6yvKzXtQfrhMFYBTX4vb/sk
7AmE1KeKFZNh+Qg91Ha0MnjwLGWiwy06yjbXD/bQ00XmP3wPnnremk82A/IHsqV68uS7E0fgHYGO
AHWc8+XWTXhAfYMMyguzKlrNT6uCnbkzIS3se2ijbcVTpR+B6SRX/fwTTWF/yQCz7w19llqcwTRk
nowffiBPCSd9gKBNIvtbVFWtIo7c15C3nlXcVvdYo2aqx59o6YRB2Sa6EPLR6leZZ/WXU029YTBF
flT8wx59zQ/CVGtYyddkChlpKdvwwf1BqdPsNsCg33lZHSjK1biKxMLvaD5rJrcziZSVHNm3Ptyj
9sq5vHCNG0Qvh0YYkVAbqd6OldXyv/LtH9Tw1sV9FduEyKFCGwm3IFSGKE/lHLq673eeoCbVz2Cc
pj4O22wN6T1ug8lQSSmxOZUbn6zUUaeeOGIbkdiQHdWzTpmjdrbcb99FDZh06lWbCbwJpFwcuCkM
eP7iHHu9AcupXES7S4A+DAVv6AFzL3hkurpsQnCnVGcvF6p1O6Px+AdV1rtAAfh2ByL+f3lH9Uv8
JGUIzT5EwJDNDin9ZGydKBP84qHR+p3dKEFxtXVn8dbdNhhVUmXakqbViTD1pKqOgQYVYm8kL/54
85r/4jgkm0JW6zDvewqd3ergedE+pXsDCMXLYnrhZuzyy7AbdgQtPxYUD6zes+RizIPO+ddNV4Vr
f24NMj8fiC1aOuuHR7zglQtA7N5MOBkU5wgYpuOnx9Mt8FT1hP6JhLGlfGn+Lro/Fk7qwXxtFhDH
/XfrwBcdUtz1SzCWKZm7lIjPYm5BikP6lE8EcKLMSz3lVzaUDAY+5dkVDfJOZu6kkqYC2CtXNX4k
/VHkVZxjdP7Yfnt8p0eyVRg8zL0LVoMcauQ21p5vUvtoBaEcp20YZg4YBGYpnbjGbXbSn63TVT9R
yVfcXu4Oki6GkfeEmpf+c/Vjd+ajDX8YrTeaNoo/oqzLcy4aiBdsHc45yelX82T6l6V/Tx+EV9rb
X1WABnPBQnaCu5ctPlG1CUuQkW/GQQ50Oq1skd+d35NObICyASYUzCTj2Z+QqTq5kO/oL5UIcf3/
H7Fmy+fVUBRtmraG/WSgw5FrLDdq/z2Kb4+in2JW08WxkEZDLeRE6D1QM9gKW07n+tilZxZ49JF5
ya2DM+DxQBZOfO8X+lYq/T9JjkGriSL/jJY7qb2ua7v3N5Rycj8ZXZ+UjJZH+ZW4L4Hmeu5ytnFu
F9FPjoCjCtbWHnQ=
`protect end_protected
