XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����=7���������c�����y%8����m�*�yb��׽4�CF�S"Ṳ�T�Cd�:b֞�������(�k Y3s���6Ze��xR������pG�� �C +:���,c��c�v��0��zذ��Q�zA��R�S|����81uz  �[9p���Gl�q���ګ�c�$O���o�#�.$݆k/l��#�,
p�ujq��{�t�f7��k:~bsqfk��bA�����WysY 3[R(����N�B
_f�T�id���=�q���g�����f|��ԟ��Uo���X�49�+H�vO䰆h��V~��[d��1.�h�8j��J���	�&�)�[�_6��'�f���j�|��w�%���MĻ��$�q�8�iY�{,�*�>-kn�qm(I#Hz�0�E;l=�{���0Hz�M�,�$)�'�h�刡>�lU�����Z��m�������ͱ�!�(��R-<F)�&&$�&�1���%�+���!��ـ���y?
�o3X�*���*/m))�9 \c:�H�7�:G�����p�j5b��"��T�����r����m!a�CC9��f3���M���&���++F��+���}�;�J����Ȑ�����T*!́��L����vd\#<"4��L� ? �����{��DO��[`x>���v�H��G
~���)Ϗ��^��Jz*��!��J��-n�QK�ʎ�O�ǝʐ1yxrq� &k��T��ܧ����X�����XlxVHYEB     400     190���Zk�fh��|���R
L-�P�.b��
:��.ui��r�S�Z����_�8|��.i��Tt�]%��B��ǀ�nz�u��*����Fc�i�#=�HwKM���C�R�p]D��*v�<��@�Y�����e�{��)�������*�'$�K0�S[Lz9�-�3�`O8q��K�� �X<�������MnN�bTvM�tH�F���w�:fG���!���c���ŚM�ݚ�����YF�8�cC��)��l�ҧ̲D���/������QCm�۽�u�E�1���̘�WN�oG��:�Y
W�\�}��@sc��TP%#�Rx�ǔ��,�3j�3UeZU9�E2� �*-���-휪ՙ���.\����Tk]JPk�M$�XlxVHYEB      3f      50�ޣ��/>�}�L�9�g��E.�)*n\x�J*o$�%��{m�t��P aJ���\W ���לZo��+%rx$��E�