��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���ɋ�q����DI�"܃ �&�"�r��qO���e�%P�j<��g]6k*�x�H�.��`jd�ƆP�6}��*���]�"�Tq�L�A�5�G�"��R�5��`��p]�/���}!:����ȥ`�"9%&�����1]��RZ�ɔ7T~>�;(�M[ �	��f�.BB�$�cz������@OP�^?�.~�ЧAF4W�"�q��Fy%���[.��C¹�)���F�wC��,�Z\�0�a5�]8��Μ�V:/a<l����	��`�i�,�h�6�nJ�Zv�:Ӵ����ꂜ��oe�����s�}>��3Fn�ސ��YO���>�W�L�8��!�/��jX�"��4�S`R�dËML�!�w����NK%��Gn3���-�Ah�%��o��b���m�3�Z�H����U�]�Fi��}�'��f�/��\6���z.�d��o�Ս d��������$��@�9
K4 ��&x	�&
E#�s�#v�	鷌8��u��`����Őަh���c�]��,I1�륨���b㹒$J��F䴲�{��e?�F�����Y;ک	pԈP���q�h�[Ȁ��#�=(#��Es�qQtԸ����T�a�����vJg�/]I����c����>�ny �����h`k	r삻�aZ�j�S�d�;��cJ�N]ņ�$!Պ8���M!5�6
�3JA{:��b�`}��j�&q���hA6�<�:����)'́T�i���W��ǫ�����
�@�&��zz��VĜ��g�ў�H��f��%C�T�T�ĺN1��iy@��B�i���O�6Qƅ��G:��@�}C��H�lG�`�b�2�=AT��!���uJ΀�\]�G��*��(\�
V�7�o�J�f���?s�u4���Z�5(��������"��#�@d���8b��nO)~Њ����I@l�`hW4
a�Z_D�c���_O*����F����E`�!��m���U����M�5�3�����$j[
�`�Br�]Tl�A����Q�Y>��\RݙNi�8��@�u����r-9L���y!/���a�k��(�f�4˖�[��uz���!�Uy��'��n�:�V�B���^E�;Fl��=|�tF��&-S�V��0�V2MGb`�W���0󐒐vxzW��Nj��@�"���)1���#f&E��n��Z��e���o_������F�tn�S���j�Y]��YmC,��ے�Tw1²za�Ӕ$϶̆� %9���ևh��i|��
V�͜e��Q�MB8�U� ��+O�C� m�yx_�יBL��P��A�d^��܃Bd����}t�V�`����4���س"<� ��
�c�:nk��l�.�D+hz��w�ʦ�&I<��uz�K��:���G�p�QN�iا$[7KԵҌ"��H�ѷ�"��ͭ�%�`�oZ�"/H#s�}��;O�W�773���4��ŕ���mek��9�L���hD�v�h��0z��˷���W��34~3<�jz�>��G�����#�0�z��w ��}Ʊ�t�I���m���
�-kk*��������=6)�J�j %G�	R1C��\Ӛf���*�T�l<�u1j��ڱ�}M����T�u��Tb�V�ry����,�a��U��@���u��a�h�u�Q�8��mש+�7m�:0�d!�Q�2�>�	��gsK�Ͳ�Ub<,-)�2�ڰѷ��uy�}����X`[/��8�\�6C�4� ��N[��ճ�'��y\��������FO������x"��|.Qᾣi�	5NEr�4%7Y�����_>�v])���wO�?Yg�f�z%O���|Y4�It�G"]t�l}l?��K�4��~�T����kTl����k��	��k�f�キ�1����Ə7�ֻ��t�@��]6����+��G4�8�����|+�L~���Q'��{��{FT<��w�4�:����k��j�F��Yb�E�ɟG:���䯻#����M>�3 q?三�N��S)B�>�i⍠���\�D3g�|��x+�4bN��R1��{�G"�56L��Yn)c(�ֽ~hy�C�>����nי�A38�Rͪ�i/2F�~ �=q��� �.L<�&�[�O�� X�ũ���L�3���,��O zo
^	o�����E*h"�?b�Ȑ.��z��6)��k7Tcђ��$��=�[�p�1ӱ.���Ϗ[�,&+�|�xؘ��E�\:�*i}Ag��joVey��̜(Ȁv���&n��B���a��9��w��j�9Ե����l��oˮ����%}�X%?�+��>��$n=v��%2�h�aEE�t��`)�H��NK;�����D,�=����S1�TE@�Yh��m>���_������B�e�aƱ�mۻ��g��}�3DL�y8P%}��x{)Od>�&*g��ǈ�±�ަ�LY�����[v��J�b���嘪�z����v�w��k��N���v� (k�'�%F.f��d�UE���ؓɬ�#K��e/�OGͰ�Y��H�gg��ܴ�Q�Ǵj���F�M�����hc^�)V�m�U�Ȱ���8`�XddQ�q��9)\e�J��T4��@���H'�o����ހ<�7�=u�5��4��ڬ����z��v�Ֆ�`:�#�r�J^��KM5���:&���]$\$��~�71T����vڛN��8�F�%c�f��=�[:���bqǒ[}��<o.�7;~9�{�WZ+�9��ҩ�X��SoK�.s{�7.sc����/ἕ����!��H;&��*�zt���a���'vo��WZ{�Z[�!7����� �\¥�J�H֊Y}�{�Z���ъ(����>�.��j$��"9f{�*Q�g��_M����I�v����J֪��}дzjG���0T?�TD���Sub��� ��L��	���{�B\�~�ЧL؉�5��V�:�f�Ӟ�hE>����|^1����,�����VX�E+dZ���T����ſ�p2	��~Щ1O�d�V�f盞�>��>���O�+��H�J�Lo�Fm�%����eE� :�(�5!<�����ٕ�U�
�@b��h����q�A&/�pH؅�K�/l�����jWc6��+�G��!�A�չ����+���߸�?�#VLE{g��*_�XoC�تl�c�K1��n�&ԟ !)ĝԺ�1{�5�Lvkt磻I^�� G�+?o`�BN���E�Y�`��� ��3�;�̾�d�F^����C�v���x"��=G��p2�����g�8�4��U�g5�����`�$l�S�F��3j��α^Fv$�H��W��5�ػ:�a�_�=�:G��&�a��SJ��f��j��<ʾ�7���6��K����cr���œum���\X� qJ �Y��qC����G��a��ބ�k�Iz�q��~��6�wY� �qf�$,�$�a��"�*)s��s?OU�t�Mm� �����Q�5�%�6�`���'<й;J�^�A!��Thrd���qu	��Y̝�6�����Pk�a�`p��g0�x�N�K|��@iZ�����՞؀m����[lѹٌm���_�`��:9� �e�H�+�I��|K��QX}*Et�)ߦ��GXW0dҫ-���oL��|�'%X����{R0G���85-�FG�q(��P���HG��BJ*��0�q����is���+h4%�i"I�PB!_a;��)$zXIM��������ͺ��F(C��A�XϘ�g�A]�ʺ��÷���ʐ�����х��4����d��s��^��Ԟh� ��tuEe�G8�b�*J�1��[3��e�1��P�!�&8$�8L��\oh��~5�E�=K0s����x?�0�	�>B9� �]o�E~���+}&�\d�˅�a���x����+]��I�����`���S�@�N�Q��q��|h0���1ob����
r��^5��i��:Q��=ؠ�3 ܮ[�7�]�o��	xMТzf��m4�K�4�9�;�M�1Z4�=+Yw��]=�Yp�·p^y�Bߜ�OޅC��\r���A��Z
�@k��i-���o[����)�E�
����,��gR�~��(a
�}&�0�p�D��f� ��i�|i#j=.E�ki����q��˨�x�`v�I6�O��ʛ ��'���7<�J薶4'��5G[�2J]��E�l_铖(�R�1��R��E�������]`;c�!��1v8��Z�ʨ�~AcZ_%����#������Y�-w�����צ"�^�6w����:�.C�M��<�VS�u(8eǹ�F[0��p�|#�u$�v����*��g����K�k�����Ras6pH�d�-`�k� ��elwr�"�밚���Uo��cr�U���,�	$9��#|�B����0r�$�rɸ&KQ� ���=b:H�S�{�o��Io������ǘ�tPj%M�kO����
Xh�[X����Ι��/��`6)�����d��C�!�d}A�QK�<�j��<>.�65۵�0�V��U�s)S@�E�i�8^%e��6����x��� /TAO���/oj�8�O;w� /��ا�Qw�z��ly��_�T5(n�!C8�ͨa�=a���y�0t 9�	�{�\%�Z��7y��ȝR���ucz:�F�|0|�j&i���q�2�94j^���e����>=xQ����F�LWn�{�Ms�PZ-�8�`ߦ'�FA�g�e`-�6M�{	b�O���Z>o*o���K��Fo@7���T�G�ʌ&<��TS����C��xKt��2uT����ߛa�=�s՜��X�a��[�͜C�"��o��z���1u�s��߿̴�z��'�L9@���!M�<�,J͙֝�/ �=�>���4M&C*��#!��2��#@�"2��!�1�iH*m*�5��7Õs� �8���5ɡ�)�X@� �l��?yTt��,A����,��������l�֞)��R�{*9�_����1A��s�[VɈ���	��0GL��FUm�%r����"Eާʅ �_T����UBvr)�z��6��n�\��E<$S�[c4�p7�J={쇼Km�,������(�ۛZ��M�E>�v}f4ͅ';K���G�G����>ŧ=
2�:~܊��U���Ǽ"�ˤ������EX�h�Ǥ �\^�"�z++�E�"jΗ�A�\�o���.����
���2����h<��\,E(f�Uv��`ـi�2!0�7*�q�
?KeW1��tByjP*biR�|��+��4z�$������I�J�b�/�0�#[��|�p�N��3b_Mk���4yD���)f��M���e��\�Q�,j��F�A�)s��������F�ܧO��K�p7�f�����y�/h LF!�M�S.�1F1ģ�MpT`�8sW��P���r�Ճ_�+��x�=�y7O�d����X���r˪�
ڤF�~����0g����i�t`V���B@��cz���Vr���ՉN�Y�B���ЫR[Fd9���#���Ij��ѹ����-&q�d��P�).c]$AHs����k���m̭�0�Rypv���U��W��h��0�.�WC��_hH�p�k�A�j*R6~��.vNP�&4�a���W�u����
�&n7$(YI�?�ۆ�Cv��Y�g�Ju����qk	`���bwRr%_0�k�_j��;�5�X|���U��9���G��I@�LnZ7h��ӆ���B�����\��yN�Q����=�u�EЀ�x������Mhg�?�������^UJ�l�IB�ANv�����b�4���V����W�L�TZ4ТY�=8����~�Z�QD�<`�������]�������k��΢��Ti����a�7z`IM���Ƹ�뎰tJ�
�T."7V�G��x��/ /��F�X�~�)�=� J��w���2���c����i?��]��i�R(��8�c>�-���n�A�1�� �' ~�w����Rg�UCv���n�U��>���﫮^�[�S�Ț���f}ɵ���>���H��k~�|J����ڢ��� 0ՎL]#ضf*J́ͱ��)_O��Q��-*J��6�?L�d0c2�qH��H�JT�,�uo����.m���t�(����]�=�P	i�kmq�'�2�
��'Q�8����F���3%��] ��H^_"cݑna�EEYE�	<�@��o������4����*[,��v��U�V���>[[qT[�����ۑVW����	x��� ����qdޫTRc1��%|^Z����v�h���d���� �S����K�4�K��,��-�]�?b8�LW?(U�g���}FqM,��t�PzuC�珖-�jS0]��o�T�r�9ϴ�m�B���Vħs��7Jm/�w�I���h� ��s��陎��Na{�k�u�(4�ƪ>`�2��Ǿ�X�to�l�)��ü$o��=�_�Sxko��3�B��C��m���_��U-UJ�$>H�O��C��"da����Эѣ�+��ڝ8.Նt�M�@��[�+Cѫn��2N�%��ҮJ��Q�R2��պc�ƾX�*p����΂V��!a��ʡ�KZe���
�{�_B2ˇb�I�VS��y��I�7�k����\�N��w��ʑ��D6�؛�W�y44���\(���q�5y]/wT���/:��=vw4$�I;���5��������]/A���%��ޥ�rJq���y�K{ ��T�"�s!��xF��6�O1�k����N�����#N��rh%��S?̘��53�w��@�~~�#�	I�~o����]��(|�Oo���
�M�v��$�(�K����Uf�K�/=+��$տ5f���U�rx�zt��ߩ��;�������_�E��}��ʵ��juzR�Ȱ���B��7�-�G���d�(�^`;=�򕏖�!̑{Bkv�o�۱�ƻ"�w$��$~���J`J�*��+��X(��/��>5+����w��4�W�6׏#��T(��MѶx�a�%����.ji}����$�4;@�r/FC��	龇��@E�}�1^D�ja�o�`�2��{5i,��@tL6)����Tb-�XIo�r�Ut�,|mn�o81�\�9���0l0ҏU�!�U��ؘ_2U�2�E��'�U��(���J���*���-C$I�%����xi舲�/Ĵo�LV М�e$Ǜ��!�͗�an��坾�ۚ!nB8P[��$o�
r覣�R�h��c�v$J:9�Y��a�$r�S,��/���?}��� ���Ҽ��@��!藘D��^٫KbH���O�e�g����E',���uM��ޢ ��k�	��Dv6���$��KJB�����L�����r(����1����pm#�J=���#��"Z�w����v'�]z�4�E� !7$[v�� �'�}�V��X��U�l�o�/�ydm�&o96��I�j(+�-�Dq�xW�tbe�y}�V�ߦG�;X�)�E��X��>A�)<l�<T2��C�����pǩߺ\�²��pW�`�I�H|��+���ɐ��;P-�!`ٽ�k��4���?΅����P�]�X�&� ���A�.�-f
��w%{�<R�,TFR@>����~�v���)�ro�k�����o���cd�Pku��*��(��?<��w��+�
�X.6K�e��!���^=�ќ��F��-�ߊ�+2�T�>�����q�{����Ɉq�+�Fp1�Q�1���qh�N,����r�<74\�>+R���f97��� �Q��e��[g��Zz����Jۗq{�}r[ W�Kw�6I�o���7YL�m���Й�2�y˖!$�؈���H�w���!�I��u�$�p�"���|��>�������YRH����G\������"��kyY� �K���2E��/���޳9M�Z�˜��G������,@L����	�M��:Y�Q]��o��՛8���4:����6*"����ZT�*�5����a�?��;
j?:fu�`�$�9�v�.��5�n%��7_�!�ZB�0q����N�!A��Qv���&��V�Vn@���sهۀ���O��v	��H�E��muʏ*g��&�L�>5�7�[B:�S_F`��O���Ej�&gS�L"�.BVY�k#uc�̮��	���'�eqNR`�%3�"�M]A�@�(J��LR��A�?���Gۃ���>'����a�u�G^� ���.���|��A�\Vױ�VKIrD��zߛ!.��>G��X{���;�Vk%�G�}N�D��е6���C�9�&�o�G||l�r_}���H0,_�� Q:+ �����`;\��d�[d�1�M��+�p��c'��Q�y��
�&#F���×/x��
��ߠ�'<pyZo�~�5;��܀���Wy1�:��x1y-�^�u�m�o�b&��q~����$"��M�2������A�x�����`�(揊j�_ w����3w_�XpH$k��nX��{�����\M�'���Rer�3M'�L��eY�rɖ�T�2�����5��>��g�_7�O���\D{n��r4�<^��ى��DxQ��+�w/��wJ�+�X�`2�@1JN)Z�%(�V���1��j]��~�n�S����SB�Fs�V/�4jFu�]t�,��si�-<�mN���uL2�U`V�[KT��K�����?2Do�j��$�l��O�-n�+{ɻ5ᨪ����+�0N(�7���er�E�ƴ*L{�v�5΄x�co���8~��f�*j�Җ�+�x󅓶��j����#@�g:Ե[d�ů������t����̟/�@��/�0��z`��)k?�J!a_ҲU���{�3$\��WUyT�i���<s$�e�������*����ja��7U(�-��6p�Aȉ�"V��!��\�A���x��(a�_��n\>��r4>\D&���ݷ�҈L���)�tJ�nPAGp�Ѹ��z+#�g����9�{�V2�9��=r����!9���s�?����{�F��r��_s�5d4�KT�|s>wq��Y����Kw���<TI~�LYJ9���Pa+4��T3mqj�n�����N��P� ���Z��͑7NN�W�\���>Ŕ��|��L?]Cz���
H\;� ]�w0��6.�I^)���E�̡�̧$���U/�)hn'ٻ��x�R(��)�KY
�U�S�L?�#���P�wGO����}�m���Wd!�r^�8ե�$�e��!ɍ�I��xnj_��ϫ!f_�豪�';����&wup�7X	�w)Gj�;DRaб���,� p��E�����t����T�k�<:ޡ��h~GV�F�R��a���䜉��ԫ��'Y
Ga�v�0�ba���_��W�n����i���I���r�W.��Hh����8<�f�	�i\���25D���:ql�=��^���Q܏��~�?�Ms�u���Ϊ"?��$�BAP��jV����c��K>�(���+���X�h�� EdZ�J�o��_�ǮY����}^r��;c��Q ���s	1E�Zf�5�4P�uȑ�(�~�Ǥ�k.K_ˀ��߶��4�]� F�{��]�9�uvOy]|R���,G�!u��"$"1�>�����t��^E�i*";Wx�!��Z"�2`�#�0j0���G���N �Аd����}U�?������o>����^��5x�@`�����'�����7�����l
g��mٵn
u�O,�:|?MZ��0ʍ(8{�y�v�a���ނ2�:���Io����8���.�{ ��Y�rD{� �ͷ�]<����[�\�[�U���>��	w|�h���Т��zC�����m�y%#,91�f�=���6e��y�c�bɆ,�7�E��Z�m�����qʘ��:��Mr��`_��+�"�k/hb����_�����-�G����4���×nD���AP����ߢV�ہ�9x��ŀ��S�\�h
��K��K�`##u�r�Ly)��$���* 1��Z,����c��x�Vr�W�n*EBkI��F� p�����z��k&���L+����әz��6<ps��o���R���ղM���{����J�"�=g�Cц��O[mx�T]��'��3��[��P,�<�`�q�+b�^\�<�Y4��Uh ���=;7�����%���.F�I��,�n����r2��i�ʚ���7��g&v����˫�r��u��/�屢�����E��t� �什Ŋ'��/i�o�}��w������_��EA��柽(Hij��<W\��m���C0�X�k'=�۵a��Ў����R�0���,*h��2�Βi@�	h)b���|�I ;וC�ٹ���C�Y��5l�p��n�W�2Ό�4EVXH���,A|��R��֋�����T�X��2l������[l�#w���"��k��׿r?8L�֋����b�)'ْ�1�;��Mw�o�~2�
@�H��[�ZM�{{�[E�y`"�$�A-hx�	X�d�Z+��(��f��E��/"5�	K�k~�O��?-Bkg:�T���ҟ1���q(2�p{��r-�l���r��u���#�$���ڬ��r�)��\�/�ݿk�9U������,��G�6t=
[I�[��%r�I�C�K��$G��%�3�-�!z~�2��I���7����$� 0����
)��]���;/��/_���O��%B^�V��:����`w�$S�o���I��h9�S��$l��HgV�	�/��u�w��׵�*K�-�~k`��S��^w����L��j@�ᾜӄ�)���7D1����/��4'��\mx���c�i|x��-��o}����$��`�Ѵ��o��'�Fr�NXȜб�*GL{�m��*��F����B{Wt�n$�HN1&�*̽)	�2�k��d�j� �/���K�kS�r�2#��䎃?��b�4Ӯ���1�����t�e�5e�T'������!�ԎĦi-�գޖHP3��x��%.]�	� ��ؕI��l�C眑��n�/�縞{�*?�^�E-wf���S�͈*2����k�%�Z�2�9��'��ۚ�H���E��hs�Æ>.�J��cL�D�4�2W��I���������%��H]�맜�����oQ��9��T4������H�_=Wfr�K���2��\�n|��	�Pb��]q�;�yu8��)��I\�^F��}%�ѭ�+��/�lWh��!��������}"<��܈�6<�`$!���=�*�ͬ_w���&H���*�l�����V��"�X�V�G³��ش��C�>��s����`���PAzg�����@t3G��q� #UΧ�,��y&����0]9eqQM�O���~�fQ�9��DTv������E�4��[� 32�(WU`ܙ>���VQ�џPdSb/=z>�J���6��#)�sRL��
 {tCE<���T@���q�`38*?%��B9�%����`&��=�ེ��� ݐk2�|\���<���h�(��H�Vg5.A �{��Ս%|��(jT�bF�,�rdB���1%��;7�;%�en�����x��o���@��4�*��~Ѩ�]e�\#�q�k���۴H���C���:}W���ԉS�kx^�
�'������ꁠV�zd[N,��?�^�  @����!��F��/�Edk ��aˏ~�_M�_W�#	��)6W�"s`u(8��#�@���f�)���^��0Z�g�W��*���"ds۷K��&v��� �B��TOLH�)����ύr�P1�B�I�Ͽ���4)�s��B-{#���T�6H�qm.��}�6��+����ݜK�&y+����~���C ϱ�M#�WՆ9���7!-�ut;�y��2M�Ŷ������qn�e�{Dv]���r ��d��)�z�`/C�*Yd�~ɧ�o��2���~
�t!�/Y��ˋ���=c~��Q��Φջl
P��q��^G�eA�(��%�*���(�Ϡa։�xt�+x�i���*�,+���>y(؎n�ۘ�L!��p�xA�*i��[�7x�rt�1(Ay�1���];�L7��rk%�x6�Te��L9!�+�P�/ܝ]��'�
z~>�|���%���&��ʟ\��i�ꆅK͟Oŕױ���Ch�򹎡�|��cQՃ��q�wA[������CԇI�ˑ��6��2������f��o����2�cL�Zo�0�ϒ���Q%�;���"���|�*����5�D�@�(� ���������z'4�R�|�%/U ���9��s�������}V�r�AɁ�)j���]GKdv�Z!+��u%K1A��Φ�6x��){��+������Jc����3���un���^Y�I������P���F�2��,9و���b��{u���
 �\�ڣfgt���ؼ��<�k��iWg�������-�o�/�a�;�'I˲���zec������tmP�/yUD�`�1�SQ,��B>!oy�.��jq�����N�Y��;7=���2Ǥl��M��˰�xL@�˶��6�ݶe8.���,�H}�95o~%�9[t�K�\�����Rl0�No�D��{2����(��Y��f�?�ߞ��Ə������^��^Xm�3���D͒��7Y�k�H!����(q�(Ή$���Nx�	z�� ��q������~Pl/c��K��'Yi��f��K�vxW�����z5P�}5�������5b/t�=L��zK�٭ñ��(�z���j+!Y�i�?��wT +h2� G�#�A��u4,��cc�M �~|��u�Y����zch3v��	���4[�ubc��
QftX��0PZ�}��b^�I}�G��x�:S�Y������=7���d��d�?݈��Yw�}�����Q�>��k3?�<�h�1�w�k��������$�\��}#j ��C��\��EU]eY�����og.5���&%E���ɘ�-�O��
���<a��R4DU85Hr�װ̫�E3�k6Oׯ�n���"<����P���c����DOg�00�{6�ѐ���T%��;)�@�����@8���c��� �Vf�Ss�d�y���]�!)d,>��K����#؜-���~2:qe;����B���,���2�ހ�q~'�AݪT�_sO/���^x�%\�=����lɿ�g�b��[Г�vʥ�����n��	=9�C�ӹ]��H�K1C/���g�̐|��)���Ƹ���5*F{K>ֻ��2L[-�v��z:��^%�1� yu�\�o[�'/��[���I?�������-����"��8)K�]��6��)����.�c���'�:*O�09Qߙkv��������aV1���F
w��O�)T�69��_�r��I�E�?9Q.q��B ��R{��*��*U�`��W�)*���
�.��Ԯ��)���q�f
��8I1��q�M�K�ü߹����C���|^GG�5t�Q�M ��+-A`na��!lZ���A�����|u��:��'i8���u��L���ݏ����w��p�V�#�
A�%ߍ�U�����b����9�����ؘ3�V�