`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
alTvOzx30BTCY8bmSS+i91lKQ396VnyYxNWvYiHrXw8UEG2XzpIgvADxr6fmq6EfxnhbpMGipBNG
teR7zSpCT8FI/5jojiRhzI0HK3+1RVB0Z/qls/67a+SDdTgdKQhtkkEP+d7jE+j/kx90Y05kQ1Pf
eashQgT38/PHeyoQUR97H0rSsaSJ57ezT5mekNqMxzmvO9gWwvX6fdycimg0SXnLrFV9HPyr5AIR
W74PPFBQmNYy0ISKsDbX+eFKjNU7QSoYxF5YC65ND7fBzmXzVSDUNFsE7npsjO2JhK9iUudaRM+1
IMUyXGt5pYmnEGMrziZmTdNATk+ANsLzIdbMTA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="VztnpiXpfqStbuW/d1MFHLyUD1Q4YW60ix6xHgky1sY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8992)
`protect data_block
IE2K2r/ykW/YgguOH99EYax9Bt7+389l7mFoam8fRsRREgzcAeGd4Minni2WiMYPOP0tinGZApL4
UZ/iSz8doY1VnSuC0NWEEPchp7mlOzUwf8oq2NEopQTv1hfdQIA0y1sUrl0CGamAG6ET0E4M7VYd
Ta08UHMx0HGLNePwlbrzaJ4lnOnmDDhEPNTsYMC/Ir+XIeZaDp4ajZVgdV26lGQraeUeEmwwcRtZ
iT88Ujghgoj/XHClAtYuIrUvwqmXRNVqTD4Dxc87KlLUKb17MabPpLRu/FbHF8KGT0EHDyQabxNj
keqogWEZIC/b2ynBDmrK96qDvp5M3YURvdJ8drIcCDwOw1szSaqwEEcyTbWKO7wCz2wDldkrmJYe
eMYQJibt3H299cQVDFShK7nUHxt8GoAmoQEcTeSXkBABO1BL7OIrLxCpF4Rcy8zh67izCCcjT4xQ
dh3A3PthaL/gdZMjrRtRFYTB5gy0Qw0jJ4Vwd7FfjdzPqAMofbRQGdquRZO17H+ovWBXdYz0o2ru
8Ja3WD05BbpPpNcpIKmWHbeP/Ix08dYb8MFx5VxrhZCT1qm55PWQHv0mZmgEGJflRoLzA/PrPQH7
xijNWrNkFEAgPvpT9quIdB5hZsayJFhveGTm52AdgwawMHs25rzKu5Hc3XWIz0sHgNFQ3d+uPmV8
frP3NAe9c1BIHtFxbegnQSRUwKMnRDHnUU9vnNgWC18Up4/3t91b8B1Gp6KQZC3VCmr9XNzCsTaS
2DlAvmg3vk0qoHfz011gfVkgk/Vrts+m1dX8oe/K4Vx0bALwKjvgdvrVLbanZvpAcxb1+RA8M8fT
vT9sl2aUOdQMLCcKgh1aT79fmQqPqLfDWX1ig1O10E3aL9g9Rg/E7VJWhqwK1YO8WfupDKWz+BxO
U7NyReFNN7l1ulCwcnM7ngm09JQNAtFOseXZ/9+RBD/AUiC7mMg664aKQfhuYefE4La2h4v07uhr
Kkjg3dpN7T4C5dC8Cocqm0jy1MojAM4E/fk57G5b8zBW6GMYls3QGYLlzHNSdrR6WWQUSxTQGBmm
kdJZWmU6MQym8LttGs9zK0/UjPcsBCEPD5H7smuh+HjCxD5ReTmJu6s2DCRdm38GHSTelOrovpsU
QA/lZOVG0tmrPKF0vtzIKBM8JXiaXQuf9TlqafAajSiG8/yuENCiQYRe3OpRS2vHqjwW6b8DP+9p
nZztqz8LFl8X6aaPmNOR+l/KobCcXvdE+Gi/XrvmHq77NsNcrXQXCKDQJYF5OIa3IZToWyGTlOSw
SVkkC+NAtbkhKZUn/vYv+avoipB+QnVUPW/zeHT/+LOfAqYQNpkbd1C5TDqckz3UmHJWhVnB/Hf9
POTYvNgl4WHT6ASBB9sK2IQAtkODnLmXM6C41rJFctKBVcUP7X/c+tPmkBD33S6TDmbgKV++Daa/
s4k4RDNWYuDW7KWmipiMq6mKLBJhXn7dXUVAA5yEVg9Xs6loPZ2oIqQ2ynuzJoB5sGfwxQuE10Iy
Ur3+QoVu3wiSefj5Q0+b/RjYG6GBDFWWmiJCP5jgmYlF2Y+NtItq/2+Bk4DOgsMUPIEZ7dDEcu//
EgMqcs2H+2r0QCt3y+agge5+BAOEYWLKJutWibNTP1QyED2dpch4SLUPbbKRphnuIZXsFfhmN/hQ
aaXCQCzgZg7Jn3YneIOSfVo9Rzkad+J0YGE+5z3OYy386zRVIz1m8GbJBAHvBoEE8YjFpJZLWdTa
Q9n8dD2wxLehkKft4yTJMsTl/OIxRlfsKGbsoca70PZUUX7OlUyUEUtKWUqxydry6PPD+KJzvGmT
vQZPmAdTq8AE5y750PPPdfE74r3/pKAUBI8jJxtp750H+9ZjU0Y24F1/AgOGyTyjpMfm7KgtMtQp
g9wNLvKGu3OCMWSV3Y0O1dwPraaqeETM2IFEjdjjqF9g9GzolnAZSh5L1THevKGgmpxPk2nqVJv8
CxMNqxFxJBmxhQvPl/nnCy3+XQZ/jTSjKzrct1x/gbSYNMvBMi7V4pc+4zCzWIaVBvNza5VdKAHU
hBoqAaBNgEGRLuH0c0PvsyG/Lc07XS+t0ntNRpiCcuYVbBZjH2T3k6GIaXYi06wkCpkyJf55ezz7
v1e+HuAh7Nni+1CR8aGU0Z55/SsKeGyN+I5LeGVQcEFvZ/EQiR7RpDifbWtPixe/qxqT5Vgh/Q1O
eyrB0CxS4K2A9fg+pvLVTdQsvQlZROW7LtuzM+zbScpJ7q0gb1nAhWrGKZ3Oeb5344vpIzs/hbDY
tNgcsP2toE2ddQ4F9+Uu1EA2T6ipPwZtEXc+fnLZ4VIu0omOq67qnLVqIaXYwUgBs0BWsAWXZm/7
BAM7yxze2Op0fWST6uXqSfs+xTnkkU00JlZo9oCvyzpTXJSU+UHrGRceORt/uZDyBvJcyEEecTJf
mjKh2wZiGwKJ8gX/ju9moQXm+o6bq2qkyjRnx/ldlgycXThYY8JWZCOILUxS9lYgqTij65yMrDrp
8O32dTLIrQXWr9W4Mk9kF435ru8/fm5MMiP+kKxekx6PnQ2CMw7lsIPqpVIpeyD/5anxogMy8ZfK
3Y3DYveXWTrAZWsw8hOWj80QynuCsgLocaowhax04ZRXzzXLYxnyiipYa8ZsMntysLlmVrAgfXCt
WZiDlV8zvOZeKa7qQTeuaeCIgirRmmf/2RfbfNtBQiUcXd9JhQUQLrZyMqyyTVndXHxjecmwQ8Z7
Vo6yzAKqp4Hy+V7NkaX3Q+ebGfr2KgW/JXb4H9ui3ikbUhCLekshEe0ApuA7M4j+vagUvEC8WMoc
Jc2DbXJyvbhcvaB/49ijejiBdNZKaIjVHuZP9tyDGB1iAGkdqLxNEjUV1o43s8ebrP6mwN24mv+0
RUqtW5Kp6OQZAFrxejtEt+cjJ1PGDQHF8sA/VdpKFDNQTR97uZqGkqkmznU+FFwPBOPLFmBWh9KP
y7NHtQNuH2Ma6CiVgnoZgX5tOtw2h8g49g1O5Vc1h90Lkzuf4PoxWh4UAthtP38+A40m/Lz1g+F/
YDIhEhy7guRJVz2+dKvKGvlXMQmgF32lVbBhd+ftM8bEF5TrlAK4P+V95t+unsUhsDv2WOjTX1tK
ryz/nCTO8WmKFiHPtifoERhX2oenTCM6ItvwdYP0SKYQVp9Mi+skBK4OTxa1NfPirwbEG79xHwPB
FJZft5rNqzK8198pEt4UhVXtcS05q9XDl8EvDwAJujiCOMFhY1RLu82CJqsl85DT7SogaPdeEIGz
ab3mnsAkWSiTnbL6cbcMnlV/8dLe4jJLkBMrqnYO5M/NbhBzpRbpBkVBvePzjcKBGYlqmV6Xmpbr
NHx7s+KKaak8bUZkYc9ladI2zHz5wF+2bWou6ghb6ayEL7QJ/9dyVmhDGD11hjthNp+hoC4PG3vb
b0H6wht2SVpSzIfe2xLnZZjF28TgPvuWBZGgPj5X/9uEL1e5uju73F1h7XPJhqO6A/Ei1/6F+DVu
WuT+0et7HPJ2EzLgaLZc+ixaBZyB52yScgx4J2i46zS9L+r2SWI/gzSIzH4t1hC7S9daV5NLvlFf
FoMbZtkjuYIxgHuTlBUJei8KY4gDPMScRXtv8hUpzVfVHWXRbWuylgtqG8rvZyc7RqExducu1Bn3
lwtPWbydFdhokwgye8DXpM06W6UcFnDFHIIDw+hbL6upEPinuZ22dTEJjB1yRexxHhQWpIJexSye
ugQVXmMPCj4XY0porYXSy0e9TVz42tSPQIHJ8ysLDwFHGqyed7SZg5A42w5Z0CVtMKAcJT9r6KSm
CE5McGjxlNrbs8JYpRv7AHbwVjWLAcz7Pv7xx8QX5tCGXSEh/rpVZQ2Ok2Uj91iWc56wMfrosL1Z
ySQz04OJI7JRv1FJ5yaAZNM6M6u0VJuMQeUXlz/t8g+A6Ip2sXPZ1OKhrR6eEN20/tJka9HFmtV3
zYKiuo6RjXoEu7+rPJtGWUUWqdhmcfV5A6Bwg0lY7ar9/3eCcB6lBX7pBSzRGPUuljgC4WsYLm5s
NMlPRieGSABtTVGs7gRvfJ/qy5iUHmNIN4iuIGdBKqPNvjnC/zm1hZvQQa+RRRTJ8cmHxMfJcv2m
feUMmkJhAUJrBfdP0xMYeimxz8AFoorE5DVI4muC8K/JMlb1n0RihVdNNRzV8SKaR4yd7I/yND5E
YyiiJMAGcoMt5CjAbGZcDF/hCZcLsmHcpiwOxeV8dSeQCsu62aQVUmh9BUdI/5hivk7kYfWD6LjI
OJfqAO4bFMvrmDATWKmJiLZejeHIjSKuc6aRPNQqcu96qEeOAGc4yoAMHBvFTV9B6r9cFp8X3IuT
i04LM0/5qxPsjlYVaYFsBNS8G1aqCKcULUtyQMIIUDbEa+VHro3Fm9UKdRKfncK+zWCVxuoor0ou
1LdiwCpO7w34O4DWKkYe0YTBZmUyg3vqOYwgZ1Rc1LQhNAgaIvSuyAunJ0Y0msGNS1jLYpUgJYPZ
YLk/poA6IJURrS51440Vmu0Ly7/fQSyI/y1NDtDXqpQN9V/jJENaPCBrtR4Yfi6jSwZv4NufXF4o
qYjJL8MtU9OSQfU4qOb00CZS8eX5ml0b0YiE1AQe3xfWWn5Lfn7P4JXVdDGBn8cv70fLXqT7OXdi
jy/LQo2fvq4zPAOrBeo9/hGyO9rgqHQmzeOdDl2gCl7IKhpYTxFUwNV5leP8djlgolD4ITKjdZt4
T+fAMr7Hux06oLl4PmSJZNOOeaf6X+6IbAtf2rcUCWv2mxOJnF/kBzqW0Q7EYaQhc9zSVdW/dsIq
I2m1POc2qgvilhsfw3os1A2Kw19iRu11GpMo8G6WLjzVY0dEPPia0Ji0+TiLKl7/AIo1aYaZb5I1
PsWbFYGeNncyWCq+m0N13RCLqrlrGGi2VZRYVYmi+goGZWuJPQ8SNV0+lYdSiVFnLb9g/fxv8dcy
KMrz0EGniV0JnBZsscNR3UyhYSNcKI8OgR4co972wtIoBAD+aNUYEFLRxhQly7fuNIJwbFbR+rMh
ZzQnhBFE4PabzBchN9xRn+4uXC6iQfEL6UE1bEujCjZSKuftgvlS+KXlBhNNsc58cEBm1l2oNUC4
sifz20h1EBZdOfE5HkeJMvtFpTOSDlekKocYikkQ1hDC5xI+843Qf9eK9CznRlBX3mw8wVOvTkZv
0cheHRosP5QkTOOZziLYv6D6JrMgcPSbm54VZh000e49xRwwt8STaG9CY+sE52iQpRNMD0RsEz/N
x49YfCavxHamV67uZKlx+ZztYyGSBsiFKb7Nw4wM68Af3nrjxUFadYXsrmL+aGfJkptN5j+UZWP5
Uh4ievX2x5iHVUyJH8GAHIWyKyim55U/cRjPCiWwBEXLIpyruCCUCNWb7WXdd4gEKX5gXl2PdYQC
18NDrpfcm83W7+FaP6JLtat60DpgBblnxWAJXJEj9vSOTXkXRVe4e6B2sudmfkV3vgU4VNMLzUt5
aGb726LRMyr/ITcdz61YFmFz18oPN2fmz0xgNZxyu/77BUumFldLkjMlqbEmd0ZuI8SJ0xCAZfzG
UejYbqCIkF8r5nE6bSPV75S4GWhX+XJmT9J5R7jusKXQIfPeVQtsvWgfyZzYFh3ZBkILbK1XSIl6
JTiQo3we2KTNVsCk4TsROFV/RYIUJM3hXKWIZlAMkdoYLWYwFApCOs9aNd8qzMhJfS7QccZut9Nd
vfu+st6QuPIzzAOKuu3ro6WMTWc6/cB08lUQvl0LUh5UwX967n0xGssyjRFcXywKmUIpQkIqR3Yi
8XXR8I1FSRByo/Q36jcbSae0X/gjO7I6vCwGBZBEVgQHaHIjAMhzrvJekAiF0g2Yo8ZDEMo7noeq
cDgLV8nJVdH74grrEVSh0C05BZUkMs5V4fqD9b+GYmtX0WILKb6sG4FADeuFplNujn9rL3vxUVfG
G5SLZlmLKYFBOfEL/kknMBoSfJXTjISXYd2diI0DoIVvCqPI0a0N30Cdzoafca1ZD+3FJBdTEgrx
F90eBr8Flu9IvcO/BWuTWAH1RFQULWZ9x0/3HYiEukQEOPTBEjwIiYk3ZOQhzVr2lr4gIg8KpBf3
W4mIx1YZrevDe3xuB058tYOaZ3pRIKRJ7IJht5rF3TO3fZDD2iqNdnhyni0G2BQfCHCnFW5mW2qr
Cl4XqCiJhdSSZjRPsNyVXxgf8Ej0Ibzqjess+VlSmjBHnUPTQKd3QI3hiGVUs9PUTIBIwXyp07EE
IE7iuz7SgzBCjjyov0vNIfQKchvj494aA+I+FrGv9oJL0clHwqXReYyCCifShE6jV7v2qf2e6GKt
rZ/NRJWUrASeTAZ/DVEJ9Fy6rFZgREaAqpH2vSD16EAPidDvEriIxy/GT92UHV9Xi7VO87qI9DM2
gVIWTFi6OvYgGxwloktgU4Sti7UuM6nbZv+cK3SveArWU2Lr7z84qWANkEEEEHUPwKigx1CF5VO2
RdKBJSYZ/QIPdIMT5gpqq3lwdP8spmpM/cY+g+BVvIi3WIByPnilFtUq8e+ARcsWtswfwTr2wdRl
EEZj/ehYpumU/kRTn+Ax3gzcRFWJ/rJOefsQsUU1qmeTckrQSws7iA97faTTg3FBGf1QyY/LhVlC
Mq5WiXUvR/i94aO6wTBPeml2pwvV9GeArxZYwOtu+6xzf/wACZ6pubyyfBy67J8+FWChlQJe+g70
we4z4m1qkMdPe4cbdwIyzAFS6VFnNO1aKqppDCTphyXtWP4/BYW2hAj5HdiWHMCazbe7+QFM3l2I
rjeT22E3W0A7UIPU2JzrWxo1cIxVaVGjUccjFyypnsaNHVriadz4ybuuAIGXMie5pviLgWi3ewoS
QkVwVAdODqPc3+XjFJfl4H8zQZ+eXN+MRS0KFbMIew/AcdrGMBxZwnsruL7r3IRrE5A2ctnUlw82
5tp4BbSEGETgOKS/cO6LenW1WwjW53ulyPD4fhjLrogYXnvg2ZILG2WmnShfH53V9kCP6v0x4FiI
AszcfiNeTrz3+Uh8jqJazdyfdJcWwwENe1EcxcIjaa/QSauMlMgJPt9fPP8Frzj2pBQmyL1qH0JY
bpfERBBM1+WwQV9Gps18TvzHcoZVeeVL9Eo0PiGFm0yOt2hjun0zYjkMv+L3hHS2LSWD/F6BS7j4
tKxJQ6dsF/1vKCSh4DhOHVsWAVeSDdMAOGwvLiftAibVPatsvyI7GlYsXIKbrPIgiX0Xpr/hCXVt
OfL8778LbNlasP2XMHvUDzF9zObiEPNYvxOtZI+UE05jjRcyKNleuVTtdpVH0vILx3Ln3qSHula6
+eQWpMtIs6TOvf2d4vyaeqTugf5Uftl0v202IPlj2CO+OOYGuaeVH6eXkXRcvVjhYy0kC5HKfOAY
w27WiOUrE5zMSPjRjCporgnybTvkt99f/4YEzYa1LX31FkgdIHp/1bTr/m5Tooj+0OOYL3ieqP8a
LeJeIRkvbxM0nKEm2rpfJh5yy9UwZYGv16xdeGUce21b18pBKYJVNfKbuFWbVoRkW2xgvdAKXEe5
u2zjMQXNnqoWLOGNge4wfN09AXuoV4RjGuLJcDvWqhVJpUaEc6GONKe/7v/LbUuHYcgOqUqIqMrB
G6mHLzblq64HNtV/OWTJPWWuziGs3rqYvFNFg55t/dEsUtZ0Ianvi0jmkSXVrclJ+b7JAHJBnM3G
S4h3wU+2NqMxdIORAVuVuiUa7Ss+MFpmzIx1ye1SCIrUe5zwYfXIRp5q9XN7hldlqBhJ5oSv1Y65
oREVO7A+ZUFhfzjZg0EZxvb5c34Aqxwb1lMq0JilsIo8Yrf7CBauabPNYW7IzHoBfaRkkN+eDqJp
8iFJGCtwnd45J5cy1/61rsjkqVbVC8N1OHtGMT91KX5KAGZrLK9oRSca7OgffrVS1F92JpNtA9jC
tZnYRBTucet/Pm8XINTVrwz+JHZGUJhgfA+J9Gjv2SbFWaYIOCviRH/qFOEfWzDpU7Zx6OoVs5cR
VQYglPf8GcrsqD2H2DFp0dsGKfZWoINP6DVgEmgMoa2h5uyCCu/Q+Mm1rTZ19o1WEKm+3vxPE+Wo
RRWaHdWA1X4MFz+82DljexkryGAKYJPJoxUUyWPSdh1s4kzpkEIEuUUBBp76IWFqRs2JuxD5RfKZ
NK1akNoJlzD7TguOFblQVk1vUoyrBkT0pAPM6ZNQu1Wl/TN9istaCD15zUHVRdf8lZeCRAHKb5SF
hhDPy/CLIPf2RJ9KtuXRTOme5hd2oDjN8lduoZO9u1X4CrOD78dXeYcSuPoO10DJgOqKRX2SPoyU
BeURl+cfYoqGxg37FBp/gszUD4LFAKxlCN9frDlBb12QdbIFHhvshmaoAnG1k6bgbo8FqUvyVFw3
dra1dH6HCre/1/GpfZm5c+r7rSxzFB26LajxQ2PTBxz6jD/6Q3qbktYimvBAaKzskYYXjyuxsX2M
RcBo1AzApFb2eekpm5f8Uk7Yp403N4wOQzy8VYPaMcRdisNEvQG4IUS/170wqepGJfu1nwyK3sG6
RYXigdOGbv/MIUMZ1m1UT0UVUKFoM7rwo7r0MpNa7HCj5UIgYfK16l29JBPzjswfpCGM++wGRLRy
laBxqvnF55exTe4sLkYOKaG5npLJovzJ/XoithFLQtBNFe6JdtQHTSh73YS29TZ+P+r9iGxJRG4E
w+jiamuwFJh5Q6LHzyqPdh3gZjLLrSha+pk1OEFDr1w/TtKBjkQJRqruGTKCN0yAIEaBSSoA3qBq
OU0dPcXwebLey11+B92JF1aee9i/904oFVZyG9TnhqIHJyW7PDOQBOpDR+ullwjGhX9FDgnMt42b
7fQDbO3p4Ce2S66M6WKCEfeND08fUQd9Npxi8dm1mpJPgSOCnS+DfmX9YxhfvHTALMgKERLV8sWG
vKj3aLFhsCuUrHRZxLEALKmF0pnajhZxSGT81gxrCoHv+mnYUdqgcQfT5sZoGI0Ch/En4NfXpJZL
VQrdOOMIZjXgNOGpcgzz3IJTJTrBZa5X1oO/V6QTxf9orAt8f0VScYvpkAWTwR8yOkkNqnTJI/XS
iCUIyk59kYYHDO75t2pEtc8rwZOcz8MtZpW3R5QNc9XAXGw3+XH8FW0BH3F1OhIM3EYgTixybUBN
0ojy5gZP38sCypzghWF/qEugCpuFLJrfCXY502gmUqGHrZccvGDC20gmg9cfFcVH6X+00D+vVLuN
6o/VTy74IQPObkeKnFPcsKeYzxCycHgUYwVojq1/XT5Ywg6Iu3U7YvcBBWGDi1wWR43JO7zx+tGR
xX1swlvjt8tMIm+zmVzpx5m8Q8K4kX3PVV3alrMlidBFSkQ/yPGI3cjy0uFgDzUDR3C8gU3M9k5p
Hz7/K3cPmsOzryk98GTBefKUmSO3QaLLhkWs+RRgxO3BaQKz+38B9gKaxu+lJh/mRCymdhlMCRMd
vZdR5VsHvC0gMAYLx0LmPpFsa7/F0uV0jcjqzDWE8OA43Msogcp5QADQ4l1vreBMje1ifpwojAnz
TZHRN10hd6H4y6XvH7MDeJwfAAmorgfR5K+6hVmX/pOLRadfLScH57HXMpdxHvTXu8bhs782shXO
MIo1X+Ge72okpY51JNIBogGdli3yhy0wf8UjJLzs6MaSTcf4K4bP/r95uEveQJa8je0d5vXOLD1S
jXLLyvLDoawtDOIUJVPWoSTM1N3HRHE+LNnPXX+vyYUkP82v/36n3X3QGM2Z2x2YXpiDxeBZoDat
J/Er9CFYSY+d1vgEEiESM0Pb1jgNRyXAVNWXLYHXWtTzsv12W6ltHLyWuoP5ZVypYiF1UcmRosVi
ZeB6aMyI0kllkifHp5qgabN6R6DlhFxJFVYRANNxATHoQ68yBRu/6YrBfiJ+qv42og5D2FE/tTZW
SYpiPrKlLh+75lhSBetAKt7p3y9EQ3Lou1LIkfpo9Z+2MS/ohjI5Y89EWy3myNHO60BIL0AHsYLg
NiFV1mbBpKee1yYCxd3yfmOiFg+WjTuMoRYDtXJdKWvOfrYJTGKmjHLGSzpXEiVuPB5wFhDfbEpu
CVtVi1qcKDt277yvqNG+lZUP6OEeOUfVghIO5k/NgUf0KBH3ui+JOtxbg5g6kmY5m9/rwzdoIMcR
5M27mmx24hFoH1/l97puxGDzDTsKGJiRtpphF3XKjLQ/0kzbHD5fDLP8xy6uoxnJ0nEvIBLO84M8
WIYu7QsFj+cYtsX4tWlbVMB0ylDEQmlPjDjW92Z/+jrFJJIzg0N9ujQIjmypb6kyaX9Mv8Hpnsuz
YaB1sZhLjqD62B/ZFTZIrbmpbOpuFM6LxxGlkW/MjzCOW7sVeDuU+FEeVQb6gXon9VQHgBQ0wJgl
4Igu5Brlj5KT1Sm8CAIYzsI0wb23MXLzCSyMNNFI0fEaLo3UNMgDGF7oDTA0QKEjoggLZNtzxhcG
rUgvzybHZ6jDS/zR96V0fwf5+B9nxjQXx8l9fBk4WRuE6Q83Uwkr7DUAoPl77EHwhBsgko59YlY7
Ex31Mj3nrIxFlR/dmK9nOatkOdvKQ3w/JWAh5GLpeKrc+ZrHt4VaQQNMzOXORIiRA2HyONeLD7BF
bsh5kZgy6IQ1Jew7z/2FAxgbzM0sL2mLopwLqpXGizb4+ip+c6TkAh+p0KaDb9jxfBOxb3IeXF3I
l4Qm5g+RCCzgV3sUbt4tpn9aV0PvAKvuI0bQm3l06W2s2C1mw62g5YfyvWAu/M3phK+BdV/oyrq+
E4P8zcg+jYlnjcF8CxeexqKUVYTA7vrmzK4t0L/inOAEyOSfe1Vu0a0ABhU5Nnf1d7vxzbNKRiIH
oS22pNTqgSY/M2ogpS0UP3gzgMGOf/+G1A21k2D0zGJwoqrstewLOJ3WdZdfNNinJeglo/SYnwph
ZbiNmHLqT7wCxfjvN/fpdcpuheZixoowHm4g2Mgc7N5+9Cx44QjdKDiKxomKkBb+haWbBV5YbZgN
KiMPmjveFW/SNJCvt9yknP+a07PyX1cq79l7Q1UvIR+hPz+6Q/KrdiXs6V2oDgvyMScfuZReuQzO
wVqYYDGBs+2hZofaEBEoFbqAATe63LWUaed0v65RTFeqbO/T9AEznn3Jl6j6FZeYfIwKJH2ELFzn
6lxRq1SOzH5xBwQWBRa3QQplgbCsNuFYTib+avQa6xekjGnGhzUUebvR0mOagPBXedUMl58Jko0/
95jBpnokJHsG7pev5SOlkvFYJkBDRkHSZkZWDRzpEdAONq6urtd5uHAo84CgBjHRNaff8axdHJlQ
fKVctKMlgIEgF4I88jzZcHJOPErOCswvOlgCvS2rtFOokcOvG9K9l/upXn94GQp3bppK0vatDr+8
iuefNdbBYSj5Uqkvxe9KT3fN23t2VbvWzB32/C/Hyb8j6TvdohNPgYw+mDgY17zCEGScdRzfoWH3
eKNIFqOhU6X+X5hsaEX4T1gq/qODsGx3dOxRPvYO8jXS6ZWpu1FAdbIH/NyTM4cIeSU7f+LoARNp
NDcKm7hIHTdXUEKlINFhzX/BCXzHJ56NiTLVzeszlwPXLpK6uwbRqs7+WkXqSkxTyVGMYCD7OKT7
n7OvtX1c+3nMm43XI2zJ+c26PgwFPW45zoDkCmY6Ab+dzDJti2nqR9f+5m6qwDCb5Mbn9A2y4tbX
8QDR1165aAtY4Qey0D8beBhWYHE7T/G88dGD02VW+CprrST3QY+TRgLLCrKyiU0Q9lphhW2R/Ay3
aftOEL2sqyxlYvuKcUPXqmkMq1KS2WB8Uhs1+fzml/vsHS+ij9BjXeBxp+zADuwtWpj8BYXC+NWH
RgBfUWxm4syxInONiMf6RgTATvkfbAZ0GCWooGNdFBNVPub9mlBorAIdXeVDgAGJsLimPB6ZNY4M
XBBZ3a7mKQGw4vYtPuv5DqrsfILd4x4qO+qJ/VY7XqR7Tw/gPkGLeLPg7V4W2eKt7aiZLlqwZEK0
qhuXmylIn2eXqtaM1AmgC/ckUdRofbiyGElWei76zd+UEQBHzUMBT7UCQw==
`protect end_protected
