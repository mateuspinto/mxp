`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10000)
`protect data_block
5sBAeA/0lZY4q8EbknHcyk3nHHY1kjpeA7xctpG7k/5pXge83IXk7AR6gaEGZnJw5BXnV0Zil3bj
B0N+moxjcLiw56x2ORnf4V2b8SR7DsXyRdFFIYP4kBC0yyG94I2M1n3VPShC4sfYaVBZeKI4INi0
SiS4UJgkOf4cAB1jiTpWkEHxPQTGK7TbQb4S1iOEiD3zKPN45Q3BYbq0fx1ssJiNfyP7JSRypsDV
GhYUDEpQHBy4ukLqdlpMsn2ZTa/a3c+1GPvHiw43armhrNuUcTqEoMQfqccFh0kGFOehcQv8MDrW
q6m5eCyxNK0rbIlqECoAgDneQdJXlRRJ3GLI9du5334ESKvdLamV7UFhRIMSecezAzR5QIVNzR7N
6cNgw5VTZJUxEBXom4rsYl+ii4w0XPLctgXDJBTY1ycHzuvItjYJ4y62b/2J/zkda072foUZcOTC
SYP7aIXmL7fi+4URoPeI0CEk3Me9egk1eABR7OKA+bPcLOZE9OQ+JepHtntvWyOPd/rqmew17LHP
IbSgSlFi880Fip9TVqHEe5QRV8VTu6bJeQW5eU8JwjqMe1q8Cg59weuPzRe/zzobDLqpSmA4iCg+
Z8rOMBltYoI5XjQGSVT3B4qujhbWykh49mXnFnlJqcv33+DYcccv0ACzr1etBE44ExRwaQG9UE4f
nhC0vxA6BEgIdgCjOhjY0VI5CJ2fvxK/fT6nw3dP09gEtbxSe4ARd7xfe62pKxV3BKp5x/K+U0kH
7VBQd6RW2yFeXc1UsyjqW/552UrBykBaCEvlktrDhcfeetkrXGvInKVpFRqGfWdjScnRlg9IO0lE
guw+RS9cA+52q5CCGXccN59YDZwX2zChwDnIJU0ekHZj24ALgpsZIicazszwOozyR8ZGE2bZaA9E
X2ZBiEzakwoMIzIwKbJkNwMGX0bGTogl/TQk69Go6T19E4MRT3NHJ+StAFRNSJnPNZkUbZ7LK2S7
pbHrHbEHmr1UE9yDzzreRX3lmpxGEusKIyjthBXIS40tAp7LROloucyLLZ2kgBkhXt1k/GRU+hFk
a/TG1Es2o4WqmxU8aw39/GDKAcnNqkTd5GO0dtfrNw5vDfO0GgpePdSfHOcAJjyzMfs+6XCGjnN8
s5xOtKqZtvypVCKCJlJPRSnSWaEOm8jQW1T7yCc5lY9S7Nx9kZlFc0P1eFKYFk5A24qmF9RVu4gd
Tyl074hRZdK6eOGc4FKlxi/c2X6hwEaaucxUkXmcxhRKyFeCHmRt1E2vpgXlIV7xBsg4eFa3xZyc
yc75Y5uWxepNEDUlSlzhH00jJ5Eu2+knGLwSjsbqRwQCQrszXMqGL/cL3fzBH51BKzWWauHffwPm
ZbKBhPkDXtBuYHMq7BWuSxx0YxwkSE9pJjQHGBefIPocK9tbcl4waqLUZtS4GT3DuHymXz3rE4TC
LHCMJmKF5WTaYgDwFwShzD/HydM+afQTq1AURKJ1PzzTWXaiODo9OSk8iBEu2O5S4IbTj0i755oY
IgbD3pPDO7BZiGr6q8EdgOQ+IOk4qVk5989d2zKwAqwe6h8D4BIkoZAjHEsW5kIfcppbMso/42Z0
BCVUkLdwb8R/KGlfsdp5Idw3MJ9kP7W3KyafI8dcp+WM34oZX9OmAVgFjwJs6FlIz/YXxuaxjV04
ckmm1KT1Q8TcLmHuy9ws2IRONE1GQ/WbgP3w73Xxpo19hGMFafwackJ/gktsCfcVXDJxBtqUjcL5
UM1d52+swKioWDK0Ok++iUDHdlNc/JsB5EYvmpv/4Oh8nYQZeMUF5v/qZhoaM9EpN0+jmxDeTTL9
vbGh/Gvpe+vWZ+xotQ2rSRMffJUbw05iMSWxtr9md3PTDk/quacZVQXJqoNqttSVHHCXMRKCTewE
2UTl9B73Yw34vi6+GTkKaA7AVJkshGJvjH+0mP6NiJ6BsvCs1cqFtc2jhH+I3VKX7nSKhlgsQIP5
qujG5Be+KrOJIkP2SDdcBqcn3gFC1zvsGWKFiQO1h7OvS6d8Qj+mJoiK+BsoZFKGlCQXX6p+DPAp
eQJzoGa5j/pUfurgrU0956hyMgRY1t1DIi5dDSHDNCCFHFcUivEG4CuvrSS01RncoUfyeH5JldxN
HUOnra8z/663Gz/yJ+TOL/KbhVaHtp3Y824WH1yMX4JdBqhHn4CvV2inAHBnenzhu1I3LEpUcOnJ
Bs62Dc57WMTUn9DnE6YoN4ep2FO7f8Qu9hVUz5wsEu/IKkEESaMgQgyY2tI2o+CekXo6z5UaGbV3
K/UrHlYqoRKDDgqiXZJ0yXPV5j6YjBjAVhwkqyPOhiFTPlm7gVbBRKfnG8jxBRI92R7jO9hufdU4
4ppqWsPpFesgT5FxHj/8Wq83G7p0rxLQIWBR8JJO4VwiTWAGzTs/2Rga0QIe+FvrRwe8cJA1bo9g
JE3B+CgmZSVzcqe34MS75hgS+u0HBHwcry7HWidNEMfqM7G6HAnq42jqOOtf/qpwuOsPr/7RKaEi
juOfZiOoP6G8y0VvvzCHRXDYHYmsmw2vBBySP51B811+kdwWUuIHkMnM5cq+QrWlQsa/eZB9lNzO
5DZYXqnrEB+7Al1kKmK+LcQv7Jo0q4ra4Y0u1X3QxQi1GUSrrvH4Dz8GtnKArZs/bCZ1OnojI1mv
Vm5OG5U7Y+0CwM320oxMl+7Jh/rWatqs7b7sf72/MKTinqRxGHeEZttc22Be8GX/x4CzsLOZe3jW
a2XFKUxKZZDc+xq0NaIY+91IpZ0+9tQzXLXY325LG0bl1ubagE4VeCTNIee+ZLRHP3JwmYnuJxzK
KcZtWvcG2yrpfzjip2tY7mHFxoJvxTWTVXyyJVrDPamMTjVTibwjMcqCu6fl+6B7KURDClC5gPy8
ltgzfAjXv6h8w8WaAZcCzTJ7oiynrfpWfF6EJUVbNri3gDeBJhWN4sYUzPPvqrspHc2Hp5NscKTH
1wErFUAwPuab6HTrR+LqUG9E3U6dKWp+roJbl+nt2KfJFTNiC3VMBP7gZVcJtqGwd7f6JwA5t/qp
9Moisix29umqU4/YK2HDmolxKI2KuwKizPDVw7GSvR/nijIMWE4lfsBSOmTNqMfV9AEK5fbUl0P/
zjPUSc5iu54BBZ42c8alRF3jGzKOaO60EQLkRua+a4C2Xc4/8Fr6QXKxgrS3obe4YHAh3X8YrGZU
zIE+bwTaHuuZ6/f/bTIzKrEnw7IZF5LOALgQ8dk40CTj4UYz87TAWPEqUEzODvhWoBkCHnwPtK7O
vKzc5BUfPUyA7SQVwE+NjxQWvBaJoJO1VVyhlnjefqOU2p2Gz39U8I627iJNuzWVtx2f8THxaowM
41DIOeoSG/R6RxrGMcYYwmx1XX++yHShkohIgirz3ns4KwjdlBt29E0f7l8XNcGdOcCQGu31Wdmm
b7qVnncwzCi+7MT4NC43nobeCl/JiRqCofCpDiULYgNyQmK4A3dIS7WNPkTFaeVEKkRN2KMlQvDv
o9H5bM+/7EKV/rj9dWd+a8Bzkpx7oNajDT8UM2/w0xrAC0zaq6LS1y5L6MCElr59XVHqYT0mwVYU
pMHJ6v7z/0vu1SfRP9mn1VuAftIz1Zrxxw1wFxI2IXDp+QY29vHpBBLr1QMhC2UWuuKKzBbgHIDf
ThfgRwodE6qL7qcsIWDsXwO8mvEtuINAhmz0HXhw+D45LuUCVSxD7/5KfWgxGJg+RLbwarZmBxFZ
0emM03/RUVtnhjBRoTr7adiRjYC/Saqx1Jl3OqnekMea6Z4bdbruXebOKMlNeOdJzMMV3cYo0lBy
AkIqrfxQxoAPxdmDfaHrZEFbJeCdXAT+1n8DcWFSKK08/YKF0xfQ46pmpJFu9Pt6bh/B3bIzag8X
fzrk/lWQQygUfyBPMk9ogP+/LP6PcBhlOU+qRnLSmfLl9iyhD4mMi/MerHXLkiTSktYoi0QPHmKr
bv4hVHgnsanhGeIAym35CjLy6aQclDtj5pgxWfZvH+j6nCGKgqgh4SdqzlCosML7w+YFEhaKhWjM
rUN9CrGGt135jkuk+fAhrZ+K3Wl9BICqp9yxt6RoS+dkq8Xh65Fg/nI1PdCP/EMcV8JHnDhZi9/C
W/83MUTZ8I4M0eZAykphYzjSRpzDi4VLYXgGy5ivZ8AVx9HDKk/H0Vno5Ts2Ktl13fd/Sovmomva
tq0IGlBnh3cpm93BI6rWSmiuw5SKMzaxvYRmy4jPNqDwESabQN3fWCHmI0vjZggfRcNroTCiE62t
KyNVBGNb7TYN7XY3ZhzjZOHkCNiMjPnejD8zD5fBmO8M9EpJoMwZ84acIBDBR0GSAGg/HqBVUO/9
pEi9fhCeZezP0EVRP/oqH5kwjAtXW4IAcqPl1NnklTt1eJqDTE68rkoOiEmH7nJcceqR70PXsWuO
bYDoLxGX/hymtzkTIguyF3ExyXpRUp9e/mRCu5Te1L8cgiZTEwxOTnyanHG6rte0fDVFL9Szfe/o
3peu35hZF3udicA6T/rULRmcfQQ3r7o3imJxmiYmb6mFI9eos9i1cfldjZm61iC39O2yPmtpemKS
K6CSMbrFz0HPEeRWVWlN/wLlUC3e+4PlHWnZ9z0KCNgdWfYC1CRAEWg3Xi+NZOCkU/Bpi8x7HoJF
cmJyqWmnzpMWUPAlCdDJukpq9a1WEiClA9JJQvbqCjMHxhojf1ZFVs8PRR4C8nJ409P+VFiqlUs/
MlSL3wjjDxpcY0zXMuRrGJxGXOXENVrY/RVRZ+J23pzsbNy6mgMmNE03IQary/dKfS3rXOimVf8s
bAceobeMiYZW6qZ8vosgzuPA8vPbWlNree3Nlr7bsIFQWmEUYafQPu8qjs9knJAcFsAbYs9K3BnG
j0TkyCzSdsXcb+Cs4OKBbSddaYXndov9zr5G7YdC0cfPkmMr1KpJiRufK0LgIWAVfdM+8U4ahE2Y
9qyPtlPoenxwSBQs5AVsHZewA9zR/IVw2LhD+dfXXwnxLblkVwUbQq8JsSFYw0/TwkJHlmNbjdKS
MbSX+8W2/NvqRzqjy1qwpzrMb3I8MS7dTh/0FyGKrMMCYFZUIgcNZKFz4A6WO+Y98gS7oEIxELSR
PVPMdLDY90bxhaXxKI1XZmZRWSknntPE7CeGiC7rLlQ6OviG3lm0C3wFYcQkGEGBXYglH9GZnrNp
RHACIcS4LRA2RKFqtNg/F5N/fto574eH/sIx7nPT4/nhE8wJDpLJzbJlqiIAzfWjQbgYg4UkVELF
+nsffKyiyFfw2Gr9aRP99uOIjpGekKmNj3BPv5OBC+8bmv0OW8kvMVR9Q3lELx3iI96wuiKG4mcA
6CvPBusXhftXLLAZvDDKVFQUIqX1hpSXojD2+UFTT+k563rISI7ueedeLds2WhO4utO9p+eAoOF8
lWesD4hCQfz4aG4b+W5wGXHylIQHMT8icglsqGb66+ZiYy9bHbuo47c15bgRzyYx36Xcd2JKJh9g
u5cGeelghXJ3jhUQnslgVHDXur7NIpbrbtXse+tDYshN+/FlfeZh/Q3tiR9cqVTNCxuirFD1bprw
ClWCXyBEIMy2LNs2HO9q4y4wnm87YqDtC/BlpAMW/YK0yCAW33EQpkoaTpwXy4U//9Nj72hHN1VR
AZBvEwb9erSrbJ5VYeCpoorzoXX/EByEAs5ccT+MY5GPS/lfWvxigcfVYjLIWJLiHw6Mhg5JOLjT
8OLpZIfgf64ayYOmF2qoffCDuYBCAgqcpYnLnmTiFj6Kio2TPOKP8lqGKyz3r0azoB4rYzWGPHSe
5piV5rY81E7UTPHKVazECEtSH3XyMYDqKVnqJMNS61Avtpf70acmYN6c6epOKVdT/GXihzHTQlzP
HAkaXEttEI8iF8bia8EcfCVv8JuZkqOOXGuDNQolniGpRAdNR7wjht7mkGFA5MfDkHIZNsw3yvl9
lcQLrae6Zsq3lPW5IWUJv5XeCbrqjNSHpzzjB+Mh82OnsYpHBBvShKdx/t+2MLQ7H26siG4T4Ugc
O2EGExTr4CRy8DLjwE6sgMIf1OF67HCWTSD2n+tCTnnFbQytNfaS73tfSuH0D551rAymylMFJ9Kq
43yQIjZFVfpL3BgCx23OpDTHEBy17oL+sTmwMd9edPAOomCxFzKXdC8TmDXV9yepWE3pWATzIsJD
c19zR7BwShA+Pp19LJQOp5fKTC6OnwC5wUwPtua0NIcpW/VLXj05nB2EPHH8sEZQuWi0iZBViQj8
6n7bxk+exC9hhBaBRpD5nHGZhdpxpuhLKtQUNyAa6MTRObRz8WUdcyrOLZ6hvSec6B48DbqRWXT9
DBs5dLQzinimKa6sjt7cKpm54cSOZG+HTkxXYnu4Oug0rBgE7TyAOQzvzWLrPJ/UWjwAaX4072wB
cjKjyKC7xeijmOP7nMmQHXHX5n5IT8uZ4RtKVU8D88kUI4upTnxFsYIW0HIPbuNl/UI3J8HXr+dG
wkJcKzyqOHbdg4pd7Eku1lHzzomTNwPiw2zwsUw3kyDdQqPrG2AO3qTLGmL211a1kkX/l6e930kV
vZhCOMDUwoRR6zmAwfv5zJj1FyKmcA7RclU0lagO7qH8mtm5olBmCAqpaq4556Q1gPfG40gLEXvo
JL3W9mmdhCXdNyhXROsyj/4fXSg4XabAO2jQ+nMgS4M9RrfH3vUQgq/JfqcTQe3xWwO/aP4mPaa9
6sb0Xo9frh0/5VkyHGxXRefrqatj0dYy68kYLoXShQH62RfA+q8CeZKQvCa7qfVquwvS4U4gIg02
uljlPOjy7uiEha5iT4b0KAHWEEpU7YyiyH5Hrse/Cj/52/Gt99rRoGD4CCVkXgZb6DR8zASMM2uq
DZK4gaodBdIInV7Y4zs853kNKHPfVgBpMfSYVvczWwiDkdPs3dnNP/d4WPOwbXoH1B+zmKyV9oBl
GY2gTE4FCSGVLTHo94io44UX6Bm73PyDHulIQZlJchdPvaBGsXPEjs2MlpI1oCBIILNQJ7lijfV7
j3FRYMq2SMTUuyM6XALJKyzfpTGI1sl6gBIKxq0iCQ3SGv1DRZXtdbP+q9W/dyIhF/mmXGeyHFUs
jhL1j+sdHbnlhymvaujHpYRxbK5BVMDwTf87d1SZVbLAlDAJma5YqUyNFa4xWJY+DoAi65v4y8SG
kRIqoNdisZKp7jSWAFU4nAG3ynG8J0qpik4Qz5FndS1YsUJYp21WLPbvXvh6CQ9H/SVoE0Z64ejO
XEMdMQcVi86q1Pybpo7qkdSBCqZI3YNb7pWquXhsRflW5dUgtRMpQdAftuazzfS+DjS4AlLRGwxX
tDmXZi3rl4Kr1XowZOKd1IyS0aT1dSKBsGdLdZ6f18gmXIyhgctmAWaLq+NlAAni1wow8naPrArP
KA0inyNLWXpFrXmgzysv69uKW5Ru7lHpuN0E4OtoO0P9wJyLojSzqqie1NGxxBy+CcpC+sbNmR97
DSEwTo6rzpwhsDd6zo119Sn/ejgFPUeJ7Lx0SGXYDnr2aser7d9v/x1j8UGxhILzQC0vPhxUDFL6
PRRJV9M2S3BtjPgddmmFJIpFHOy+lXZd+7bAMxiakujWclyv0xKkqJSw8yW1K0BlRd3yC770Ttvt
Mm/vHi8ocCR7s5cvAAm6WDiRw6vIfKHZIns+bbgvBUDYHfnkU8sQZIDBqmfj3+MSEhKvAdJb6UnJ
tJMtxNQOr4tPO13LQ84x7Infoly9ft0FFA+5QQDuJZdlYZIIHfPzayT4HeSM3+XisAZGxroD0OjS
J0QJolK0NOZsbETNvvb3bLH3Uo6WNWoQNNbK7DYkkD2T9ofVW7ogTlmPEXtK53VuCy0No4oPBXSb
3qbbxbZ52HnU1iVDSSNpTCz7zsER2JpdDNVIg8EqYzSlOJcrleFdtZvZv6hhwLuJihJTTK7C1rKw
sb5swiGEF6pKsn/EbEqDAjU1mnVMMJVjggEPhSgvSN6ICVmvHV90FGu+rOcXDoQWPw6wq8YCK1cJ
2liYMCGs9pXi8RA1CJiD1SEhm7uOxxDQZUxU1xtY/VL+nS0VmgBNgqiKfuEJ9k2Q1izdHjnD2HD6
FeOb185JQJxMX9TPk7nfsLYhCwv+GDwDKHcJjtJed06qo5NpSbaq787RorVxOC9y+NOgGCtIrTI+
Zi3AmdJpLRjOsFSLr6cTXRYjLIY7S7JMEWmJgUbWcr3vZ0z1GlOluOvqmW479StBuXXR5tuGLU94
xXr6jz1vJLLeZKO6xEVmpIHL6k8+avJSD6wSO+abET4cbT0hxHh2aeTAUZdPJBZN4xInmeWx69FI
38PyOtRetXsYcR+ZBiUAPJFryNlJuwbC2f4R2gpl9aITbsfgOVpefke10SH8rcGh07hdKTWSYcZx
gSNfA+J14yPnuaXKwoHlq2yrsiHQAZ270QWk0Gc2/MuVPv/IXM+egPzFA74z5yjQoQCW9xZIb/ig
SWczNZFl1ZjRMESjJX9T10WDzVkrPgD/dMvAYiCL1EOy81I7/kS8QnjeO8Hp4aNBtE1F95pTNFdj
nCjm8N5pSeMd7fzwnGM6899qiJpwWNa1LQ3mqoC/2Qq/ltdf/z4oC+Atccyi+opA7ILiluWPSDJX
eyUm99xGEvEqBcEQDrNJUKxHoIAECasl+r8YGIInLBL1hLhs+SsQfFeNNEXtJ8E+S6V8UJ5ev95F
dEUigLQB9cZ2Kmm4S/Kwxo8GwB6myh21eXHJBHQeEJ2zFS6Bxyb8Kl4y2XGiCKhY3w2FBU30g53C
6miuOyJLGNRGI/h6Ih3QRlpiB0swfb86u+v/PUrmqCmVSDRVURtpCmy7lH5s2nE0fsFa41pRvvpF
q7rh5kG5HIO5gLTYc+carQT1C2nG0H/fGOX9K3achKMcm9f/ZZjTJVwS4NXX/aIG4WVYoGacRRqk
CIpxyS52LK/ClTYmr4QTcw575IfFk4Vc+0sd6PyqHfCxizM1tAbKYl7qAABueQzF62+MY2GkQHdw
0knx6nMpalL8ZqQm//twCOIwGWs7CrHOI88XCX5MSyQUNi2NfsngbpaxHpgKCLGlrW1v6sAxpa4I
lrhryiggwjhVxNr2xQvwQnB/EwmL3VyDMbs8kmO5GLWNuq09giS4JHs1hoalxERWHiSu8Bwu0Nrq
76ZZdgLV5lq7NH/FDUDrLeNqqkiLlDok6QTgd3xsgghYQGaytm0wORhsZOfLlVpfPU1vsowuk2f7
NWW1ypCOoL+jYMSToN/H2MZUHI/wD8AzeSsyVBIMBIHnQnGudplIWn6J1bH3xQkQQ9r995s9tty6
VN6c94MAER/tcb1U+YPcPMZAbyPVNVN4amFlSPjc36u0YtmQknEVt9NCW0e0uwKLCZfsMz2aycXE
9dPjH+K3pLgwMpV9wAzaT/CmFH+hI9DjHww7RrttdD9UiidRgI8NxqxtD+S1wMZMa0ouRj81x0ZN
cPDzcWLugSJFvf6lci1TzvB4GhBqS5+V83RHlCJJ+wMJ5qRMo9lbxyjFu4sGm9teGklCoXWfGwDT
7PHhoZTLFoJERsrZhJ9cYGohnw1pFQu/lQleGcyhE5SQpHsK6UA2RLa/Kfje3wa/NLTbIRtgxKGQ
XhL65is1AiSCm3FqUb22qGKARnMbfwLXFzdZ029SgR1mRjZB+esbTN9fG8V3VyY8205KuvWQ8/5e
x8OTy2sTG7OTpW4+48a5QMQSjmx565G95iSqmP6YsLrbkRrVRAKiVZUdcfPd9Z9Za6hhMrJcI+wR
4/C2LhYLni/NaKhmaa8V71qvc1LbkD5ZWlCj+GIndYMjB2tX7DqhU4XIzjqfwhFyuDPxTJzEIEJ8
uM+Dgt3Y83mkXExi+Ui9G9oB0HTkJ7RT6TF4pNd31kVH4k/TMLoM9oXxQSZrFM6DFpEnzW+/0/15
fw03/D9CXaCaYB25gaX0b6x+1Fjyz+84eXJ8Kw2tVuDv81nHc6OIGnr1jcQmF9q3F2EsGC3YA72w
SLtY1bgG7/eoT+FVr5EzNr+/89FIE+ikyytLfnlDTxpG+bjHPT7PzDf9N0rA2IDGQf46cSFua+q0
+K0qiX2sNjWP0i+5lSdO04NuusPjSPuo52ildlsLZ9goJNWi64O8C2Nxs1aK+1LtLvVMb1MsXEQ1
ldPAxjBIpHvhGQVr5D+9f2CWvTovO8S0eMpKdIj69AAS2y7rLrTw5xndJn4zS3Ou+Ry9rVqeR4Qo
vXU5VEFnRKGqIrmlxzuTmtuHuy6qugKLmv9mFBPUN9D8uR2bsjNu8hNshY0qNDfOKAuQZCjWybJU
hb3tj7Z1eSCEMsN5SLzHFm4hu5ynlvvle55Er7X0SvlNWjabO1KtpGjxkt5n+a4/wq2GE/SKP45n
FIUkSuz96dOYpmRzsDiQNdmGKfqyEMalq7Ljg5/Rh1avFlAuOQW96qroJTl5mUGg5pBs0H9xBzI8
8hzN4ulI32Bm+T6H+PMrHJyvAMEYDu8quS1+Jl/TtsPS40hGcpH5KKylqOiIMVZ3fo3cIiwCDT37
4GmaTxtTJ6KALfN1ACxhgrsYcwtmxeVmnBJgWzd9NOX+CjhIIUiKGvR3Z5e9TsD7BMSJLNZ8eMgu
l+yr24XDEL4w3carDYTlFzoBBKLqKH6B7YrGbjTuEjpzzFN56dZYF4yHOua6+5GTaCgOIjTLEbdd
R73CQ9z8vpF91cMUor6p/d8+yiCt4u7VcO/PkmOtYmYLYqRpT452ATAo4s2oEmuV3i2KDiVpmt3c
rarGFxxZo/i1NZoaAAlLftQUY/1Id3UYtfd93U+wOtac/I6+pVPDNrRw+S1rvTyFTAIQk9mCHmjB
LlGeovoeXfm8dYtkb/iVx1cm7kiksK60psHvhCyTf22ojtAikSRX3GDzYVa4nhTkXdZjT8itkLa1
fKOnZ+mxOlcMYpnEw9kzalws/Sp4hygiG0e6Gq5buU9iFGvQIschLkaYklI/fpBgKczkETjTQFEu
2lcZlnSOi3L/y4zxC87R04K1pboESnlZKoacGrZ6gUKMh1qVv9IcD97OMl0KeJHH+7YTuZn38gCR
xoCrCEBTnZQlAE9F1Q/aA4DYoli9NoE0Xf+L40bNifka64rRkL3sltkoxlT33ddlYHnV+2P69Dgu
nKW7+7L4qnqbyCdRM7eZ+FXZYLXiEWqEWSF7gofBzndVRDyrbzXmKxVmZozbzrArgwodJ8xa1o8Z
9z65MwACNQIbdOgqyxZgKYXcbuIRAqVPk4IqzLdyGamD31f30R+ezujGFYaJjz6VgP2/VCRv9Vfx
fEZk/SI3NrCekCIIhZ2h0Sver+bNgjB+VIbhzUdGTFr9ZeihIhIGkosFxghJgRZCrPE468G+rm6n
MpQXrvaGCl9A9cpcaqopglBh8+/WtfKRyoxAjBlOPSn17SE8N8zW8NAoN2Ny0lZpFwwuFzaqhAwq
2pfzSvvdT0nMTk5VSWAFBkznAoOwkCawVFviZyH54NDpElez97aY9B/pEYZPJkelKZQLY0J3hamb
7WObcMKDji8MKezVn7YBO7RXQ2HtMa2twWP8To+LwclO2xXkPNnGd4z/xFXfTXgjvNQAQuRXPcWz
n/ud4AiuTIvMpfWfOkTBsQ49Jyx9J9R0q5Hhel2R+eJY/zPav7xgaBZGC15+eShtS6Ml6gM7AQsL
3f0u7Mroau40SkuTU6PD5wtpNSguutH6kc99QGSsWsGE7kDsE2yKXr5OWDYTyrXv1Mfe5f5QMTEZ
oF8T26r1mEr9yjz6N445RL81Q0a4Im4pG1EE9YpuYT9bKi7T4CWUpDrHo0mcTKbOh5YkBaG7jiDw
CasJBxa/R7s/h/Vv2Pn4bsOO+c2cn1sX/eenfW/8Vvni7xpQ1OEd/PciUKJf1ZmjlHq8YseSZpQP
XQknf0CMAnmCH9h7+wKhCmO4BoV/5yEqoDGgTBQaFO9iQBT5srrnYhPXkFTRsqmnJIb6ffmE1EV9
3fCEXL9BzGGbpOD9ztJXSc1hSyvOrZYT80PxMYxuzATjFLnQWCx4zQULCySTwR3lEW9iIdG6dkGd
UR+lg86R0hN8+gYHltbP0pZjw/SIueOWWkpxkOgzzjcclrzlyPNc+p6X66DPXC2lLo8+1nKoJQtc
v9hN6uZod1boQZnBYqNFSsUwQiPx6vzCXYWsDOBgZv2HjeUuMybsH66gtfT4lIq5puPyJgI8qPdP
XuyEW/vrPjeMfcudOVvk4My0jFU34f9SfKk5ICYHqyN8u7fmbPBmjesvNHDJN85bWZtSBvGb7yAS
ef8DBUwz6+C53BxLRk8RDxEHiFL0LGBN/TKfk2k0F/kRFsuwbSnwBFLfYOcMlrXRYak4lyrkXHv4
sVwDx3JBSn9uMTJFS+G5p2Ov3ONkZnxcFLRyKLmrxkw4ETL9Zs/k7uZIAN05wUlOeMKng7uZqR5V
gAbG/QK9nvqubnnDuy5tRvJxhyZWdTo0c6weDVfCk1PdNvM7nUYnKYQR2mUUtH6Fo6CmDp8CxhK1
3YkJ1AP+EmNmSH8Nz1PRsd2KnqXx9tIaeoCJc+DJsIM23mea6JXmLUPVlDOI+tBskVo/+8gKHbi/
oGRlNJTym1I2h+I6cAW/Aai1TmGkn5kvxT4AoUU8deoDm9pJ5uQSnVhrI6HSUGymHTcCx14a0AMK
2WGIzmcxoCPzDZd3jcJuMbg7kogolE/1fC+1brQaKQ1l/Tvxq44bwk7OQtYgf4ctIPkP5wSbGGyg
znciFctJTWFIcH2IBmzLxkLkLWhe43oZOyNxC3cKyHj1VuyaluzudHbEbJXKAVx6yagnVi91idH9
UsR0vZ1sxs59lOGtEBQAepxoeIR3hMbT/CxEYWLMlcHIdsL4PCQi7yNAKi/a3OoHnCZ0QrnwgJGS
Ndsc6Eiv04xp1bj8phBGzw1n3YvQM2ujbyutCPsFuuyRs/9OtrBOGY+fJGywOK4qvjZiCIESGP8o
WMJPY6UqynJAXuHyuNdGvPNC3nhKWctdejcB1HJiyZO9TIIlp/vsLmm+TCZSx6Mse/VbMycu9gI0
TEKg474d/VErD/OP5YAY57Gri8DPPCePUCersk/5YMk7hoMw5KFrzCOZpFFtN1cmBRWlbrzZ1sLM
+hyl4+bnS+evm9qkQF11waLQaWDnLj/CwIhFnaelAiedJ5cWGM6oW7YDWZXwyYHV5VgNL32bBzeU
K1y4iCmbTQhBQvZQQVbLFC5V/bXFV/ISMFteMsu4+oL98ShjfSi6/mlxkXUNadqh5VQ7qY49MkQR
BclnrBQ9PCcpv3JtnLefUjZXAd9itboIuo0/Su3KCxs9ttC87B7vw+t26ECsRGbf2tl3g9UCtZNV
w1P68+Bewuu87RpFeTJ2LVMOl6Rfl9rwUQ==
`protect end_protected
