`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12192)
`protect data_block
+cVTiW6rcBWDU17t2tXSSqrrsezP95uB4Q2ncCetHzMbsTm8S0MJY98zrPm0gU+L5VZFkxzkcNst
IkGac5fW3iUWbWZ+yd8KLbRXHaHCf/QKK9oolX1PunS2mrfcEndQOJjWX2xL3II/M59/AFNkk7Fj
Oim5xb78oB2eAGBNwwuhmbHpes/0G21cvnu3n9uV4Lwa37pbteDaJ5vGc+whAI0Lhz41evebuhEV
Wtnqeb6c3vvEpu0g2qfiVy9vTKIaVF9Q8RYZS1hUbIO3YAmYu2WZJcoYpAaCoIiHavImaxSEuA/H
RYgh+ezeI+/WGIBCDx8nxq+bosjjFC9mXuPvSZB3d2p+nPspTLD83VKZsc6JvlXn6WAhVgmfzbZT
7sCDGQsGz/uDOJR39Fh5VU2PP8+PCVLKbXSvKM6hP12IjlsfJ5y5PArTfsfepqZF7vKRG0FQDGWd
eR1c0kWdBU1aEH8H73Qd4fbgmZISo66S6dN2urU6i5sUsmPiD0aOb6i4HvfBNujkuMZrE9WpUARG
16S8yrVz42CwXXdKMCWT/e2zTwQAcKf82Z8AIzHl0JuAqnXJfbiklDm8UlFyJb8PtEi2WK0eqxuj
daqFgLkQ9aky2tXPV1Dl0dyaRQdpSZT05iJLbPWdz7nZn4YkjRMOqpfEMeujy0HeM/ooHsoNL/Bv
EpquH1brbRt6mYTCGF5rl9OeFgzlkALdEDMhouFN62hC3Nt3ERufejNwKh31r15gp+AlBFkOYdMN
poWE8jHmHi3L7FeZlUm1xgmxRACMGAqS5tSgnebWZv+c1JmGa40ZWL1rJ/zDpIIuIXcBEEVjzUQM
CElzdFrtZHni/v2fFHBuFOPvMeEtvEw8rsWJeyMJcAE4Fp/kAhWVeM/fd06l5mUQCssVQmYC8b+7
YfTQ8k6+OG/PLLD2KhSIMI/lLqhsSmQd7JEqktsfqNdYiH5dlgeIlH2qrZQDEN/CEY16gyeGOiys
XPCWtjW0O9SJY7JvrrA3b2YjRaiMDlQ0FTzrSk8H1/jeh1xXB9cZbQTH0z0KNdRd+KMELyPI8Tlp
tt8/KXFVBmE1kGzEKa3zq1B6PCHp3xIyBr1ktQGVml3qcJ9llzQRIptTuRv8YmS4xUKjBV1H9JRD
2NTBPnZZZ+9w2gyWE9IB+kJY25i3emxYJW4e9AEPx2He9Xondl9Y7e5Ta5qUgVWXUvq5guHnFKRl
/vLQhM2Ox0MwCqG513IjFrWkzYGO6SRZXIidvM/fS4SiZjoh2q+lcl9ZVkD6KpOcW236PRPMobuC
ykpeJUtIKpl+xIrCjzboXyp68mXUhgIN8NLzqCKpP7dEG7xJi4PuS4UbwwD8sLwb4yCQpq/p7pgI
7CzAItCqkz7zpCfuuSrLw0sFj1L+ZPUpDtiGGQoEAOxHPtqKIEU/oWaQs+x47fjyBDWomJumOL5x
mCOYpiFADZXSTPn/s8OWghSW8X3SLSatgmewu1JEq5eMsBKfxyqaJOGHlw0zgE+GQ+DVYe1Dzuof
c/kgBigfiJbaZ/IMBRrBYfNlNUMAAzaosjSRtjB1OXkB2RTzI3sFagSm4i75xet+wdCVsV1g931I
YVbPhFYW/isbHHNlVFvbNyiV+h7UNVqYOiDSY4jwX62uU2EriAqbAA4GZs3vAhRmBuAtGHrXPcQs
2ImyD3K7hOw4DAXG6Ne3L8lMp/J+AvFX5PrALTOlQO5nX/YoJt7+LfgqXa9q1vHwM21FF/Q1pkfA
7h74lad4jGD1VtJHIzstoTw6WUCjnu2WQWfWeVKjkX6CO5j34hL4jlxyrkUq9GzGnMlYuGOPbmaj
lTdY7kGtgHE6l1cBIf19mVhmbhmcu8OzOquICvgzb3raL/xfhdFLfgmlrpAwUxF87502iJ2xxzMe
HhGdlYGhmyjqC7oXf697Qops6vRBvMRwlVA7kZCrXjISDHLZJ1qXHNTc6kpy932A6CSYYvYJR20j
JSyGQKQVnYY3FhZP3VJmGgVpkohsYSjqAW4Q8N/YTfDRWJpQfl3RQ//PNHys+dvBKFu0yJ/IpsX1
saY6gZbq+wTpO8KfxTbLMHjMr2A11WxVdlejemSDAUlbWKWwfX+Czz3XXLgOrppH6WYGXQQKZ6Wk
leymgzPhQFWrdT8TkRmI3oBUykDMrNK6CaWRm5nOaNkc2H8mMU3KWeltLyXyZxJZXEyilcCpsH7q
3mmQBwzwH/XhUQMwZnWgBGppNyOKqqPMfTMsmYZ8RkHCtEnzb9NOFR1LJFIlI+Wm/62132ioRtXc
8l2Swnwou5MwxoGpXrLSdieh0mlsh6b08MajZXLsIklaX3LYseZmo9KVP0TJ0GBBhsTt0uGkUi8p
YfOCXRRmTjRGAxdi+jaxwqMND1JalB5eRV3bYohJct8P3W+NrdODM5O8DY7c5uI0Ab0HB648DAKm
TqF9OVdLdSzzzGSKFPIY0xUKeWxGWlNV4zcK3EZr0/Di2JWKRgigXHZNZNabdLT+W7phKi9osXFU
xjjlKEaP74DtXcP1mNxboLZU4ADHmhyugmrLvRXusGUxz2p3xwTGZukATxfxdHPPTKsrVXDEks3q
G0+jSYe8p/8ry5YJ2YGgpBRqTyq/kl7JLYopNFsJCoD3lVE5cSx7fBccXGZtGZHYWNuHIJRnO7U7
Drd8douHd5kkM/R/8CuJdmWC1/69zeLbZcOpc1vcUbAL16ecbqgxReowWZvTBn7HimQpTwf9Xiew
cKWaI+A5MQ0f8PIngxh8p4aYQDF08FfeItlh9G9ZjhjntqSs3TtPj2i21X004asNfGibk8ajfWJ8
kn9Qjxylwj5OQs7F++deUhjIG/tF6t4qTzNaiCPDBhERXmswOlq0PnmDz2bBweumVYZW9QnFOSuo
J8gaDcbZ2fPVOH1IhSY8iC7Oy5F2EliPB7CoENsB2XGgsVIPULWcZfMRQzUBN30U5jFFHEcqHWoR
8N0Erw0w8m2CXcbIl+zr/uqIa0XIqOFjXyOOYvjtRQw9vxtxkfirzU8JzwQS/ECoJqiWJLdD8jW9
CHC5BNhkELwFRyyn56BRSjLaoTxv5vnS6eZBFOc6rWsaCnPk4p+nu9jDVMM/19Q5Y+CmI+7K6E7A
RM7vjEnIDLl5hV6DF5qTE054ln9e7TpjnQ9rklpk9s2jBwIcOmSAPF7ez7kEaS94aueDzeLnrsVe
zsx1woaH1v3terJZgy7R8ggFgpbjZluoqgVN4sEOjRMVe/cewQ0tw/huHBrUCkVS2umztAx4Axim
1Trc9AeqZR28oiBZNrRoUBW5eaU35NODDnWQt1AKYhRdt28QHEZh8vjXwu8i3teCbHNn3FK0mMRf
AnQ2EFGk0h+qEAnL5Ygkvcp/KhJQ5yi/pKF62FGDvSd2/YZILn0wIxdlMl0UMb99HI26Z9UrvGZC
PL5AliOQ3DoXkPHY8JpOu3twvBc1XIw4dNG8X4H9o0yagTXOaGOviLoIbhgUwHj609vF3w9VhBz1
5JbR0qVVInCiVJxwFe/9WRaLWr7P3I89ZlYUx5QV2DdLEAv8lWjFbyj4RMlbrJFUjYJAVUpZGx+A
NoxcYbikoTuxvX+hCoANnSIBB/6d549F5eyKfakmphPoUm7a4JhL+ngrm0OLoCKHn1/FslYys8yl
XvvUUPLJ8tkS9tzE48ePzAKdz0DKCWXD+AvW6JRmynnWTTlBFOkkxkLKx4bFCCdFtcvQCnsebJnK
VqXdsKSCswgkKw3Z36a9D+8pLu0aiipMIhMLNLAB/zvY90PqzU3KOwKNlLC08fz6Mm1Rv5oWwlkZ
ACAjtSjq0xYuhScdupIE9yo3DYAJmP7SA/4a9/eLUX/2usSe2M9sQHCgC+oZKUG9Dk6CPPXuoL7L
ToIA6xzC1PNLNRarATlV4KTaoL1+qgBFov4ULCHpc+OjAHUyuFeXt28AHOh5FAWYkgfQ2hfW+26G
NQJ4+iZLWD3oWCS1g9lrwQQhOcs1YPlQOILspkzADlS4ReWPHiCvZk47iot41LLZdAugyldT6MYH
bJNRYkUKnUvy1tqpC1a5zaByHP087pdgS5Mq2ADko6V/5ECCC33y5yZENEw5dMUmuDrjaJ9nihmH
GVPQV+GYNQwL5la3RkvCHsiCKjeg8yiPU0X9a9s+/WrjEq0Oud20EGfLrloSRrxEQ/rMdfi2RfMB
muPbBbOXB6U2LmK+cG4hLdqNnvfqQkZ2/D/CBFa7pSvDS4CHgbMD0ctcgnKSD3k5KNwAQlQUMJ+7
qlv+xfnVhW8nQlMHZRNFlwkrZ2o/FLMUlGph3GvQgVHMfi3akKlGw+s2kQgptkRu40Kl7MrIlBNh
Tz1Riz84rKgKH3ABIxkNq5/5Dx3lJgkxclyB0NlAH3ifQThRCycKm/N/fiB8XroOyEBCkN/DaPmc
O+5Eg76g3cbGoSruuO2gG8QdM1eeM3nh2V04Y6QATGYovI6t38bIyk01PSgSW1p6ZXZYDn0GUZsm
nBFnujRdNpCEy8ROtk8YynS5hPJpnWpPvmSRfRGEH0M0dwPc3HjZV0aTMSw8csF23jaaSfCPr0Jw
4EaznaZm5b6BfmW0wYCchZi5ZKhnDZ7X77M8+aQZoGiNOe9p1mTRvvS4V7PiclmW3xPc6rmbN/0N
mv22ZGmZ3nGAvS9GTgLlQzaX95ss3WyZe4p4SkjwabxtcUFZcln+K9mPMAkgXu0x85eNWNWujAvc
t99YU4Btnxg5xHuiNoBXiKjFOIbzvA4topFpLIOjPWx8BAEYLSV5o+jPcPG6NZCW/jQ5R31w6P0Z
f+S/amkPFSHZWG3TGeFVLCqflCFYZHi6IVC1Lssyb9vuvPsIUeT8F3dL/qNfbLuvyfJVzP/78Bc3
lT8YpzwmcewZN0urzof6EGT5NC+fJA/kn09lU6NIS5RP2/SqYkCtny1jRA2kau+TLcmoniR/tw2d
8YQAoLCqjUcQPRmFqN56k0qrxqo00zBqTsPP+MBmn6CkJizcUB48xakhIGOXQQ/QJ4BWmcGJptYe
K+24fmb1SzSWOX9f/OJNK5fp5IVRt6qKDEjudLoM4eLXU+mpKfolDcGY5pgDIJS9IWNqqt8oMS6T
zndebZVUHH9mJJ3dY5LIk9yUw41ghSfJCmpUfnP9OtjrkBJtxbo+agQqmy3zNxO+L7tnh0rIGCcC
vf3/FOoOsR2MHdR6rZi5UGgvylvAvST9QtND5SksXCnrA6o90HWBij7WaT2IcLwV0fN434nrs2tH
jwfEFogQN14TaLAEJL86iph0t7kKny70pRT/IMDT2JYxBq/HcnZhoHY0Njm3Ldw/Z/5+l54qNOzd
MGTilAJuDq17dnpCSVY2QVAyiEqAwVpOCKjh5XDt0/WjIPRrpI+zdCzVPhcDFBKQ8XNuP25k0Cvb
JjzDG3tNkQDE01ueoFg53PIcG0cgjDeQL6+a0TnOFaeBAQEuFj0DuIo1QdEl48RaMDbCLuiPQXcv
oo5SNXjzffZCiC50E/xf9GQO/gVcu2d5QudfWWYUi3D4yG56I+lu781AR87ZnuhPoy18SIH14JCX
OoLoyX1zmtV7H+DtyJFzqLuRLGts8pMY+WGhS5QeQWTuHLaruXH6C30+xCnzIg5GCdl+IrYvsCvu
fdD4AZ3ncR9pndYCJMuimX2l+8MUMqjD8Aoy8G0WpL7vCVYha6mPO2VXvr/7NZWSeMzJBylJZQSY
cTo5vRrjHWEE2ItheJEIKlAf3RLoQDh25+k9xk0N4l2BKFK/3pOspls8k1Tfr7oL7k28zQTbtbNP
UDdLRwJkhY5e6+I16YZ0S7wD9FYLqIcCyjSe7pMeGTT3RpViDGujwq+603cbQ14W1+nj3laIfLk1
RfAu9inmF/zjVMiM2d7O+2SN6yJwwxGu2uthRv2Zq7iinOWrVH5E3NowhtjOXj7s78ii/SIT5qg1
KwcktyVg9pHRshRRgKOoOEaJurXe/3efLa6vqW+tQdYLbsm5W5QiOkLfycMA8xv/fhz07U6blaUB
3lo4vLiXHoUyf+xITOd+gm7YCMQmqqIRpZpnqgNqsaDr22bT/wMMDmWHTD3WqAki1BtRdwWv8OuH
wxKBNgw1An5LVi89/dJ3DtmhcZWUhpqBh948J0GH0Qzn1snwWyWiLrlv3EUnRVH5iGt8135fdGgy
Ah2UP/Qa6B89KopEMjtGlb7ejIiEyi8ecwlf2TGIUw9WSNwI1RzcSP1zDhgDvdszvg5wuJ5hYwy2
LJ7hU+MlL8TZndFpGCZDck9CzeKK8ziNbLkATor0jKsU9ASuxUFI/Wtsmdm1/1wZalUJTHgJmEHd
kSw/julabcKjXzEHQhftHfnkI2sJjIqd2sVRJ+fYvHBJxhheGkYxNIHsz7JMp1x0DdlspRTlTzA3
zNEBZIOVWpOeaL/qCFhccisKMPo1OY5LbIH/mL3nRev3hW+w2iYeHNMcXxyRt3nahT9Q+Q+ZH0eu
YQBBdsG5Wvf10H9AF4+fEMj77caW5hg6Hb/429KOeP7xx+TIbwVUTCsKjqF0JIwsay1J0A+nvtjF
UjqBQ/ytXSV03r/au2reGRyFlSYClf1ml4jvUTsstwOHRxeerFd6jPgXA6dYe78BPS3pd+nfqUBb
Pul4QLh+bsi/Q/250XvRpjWa6yLURSsmlS8ZvTjZEDlNebcEusAn5sqqZUNzhzrjJk/3WHd0DYw1
lQVz9AQKbaBxYEy8K8kj3qbA+9nPKE84u8DShzkel/PsdNQjPYu1NuTXdJTTpU7Sr6skCmwkRhDX
HNXZ/K6GfGwtWzPVFyNLojkQXfmP/K+a1yOn+jlKP+bhnCn2IMsogxe+WSnXhUb2BnRwFcYlh40h
O0wOlHkUsda4fZJ9Lx7CpHuGmFWw3vm9I+fnjwXoYMIjoC9nOAJ8VZzlZ4uG+RBUGHpFdkYNWtm4
anIWwH2wOKANjRrovzHBtXqoIUWKtziTuvkyguGqaSeCc9IoGXoI1STJeXpPHIK31mXpebwJve/j
LsvVw3NztHR09vNJBLkyrkl90HZrQEjju6OjY8nv5dpBkBaS/ggBgEjlI32kx7PPBrwGEmWcZ4wn
FfGULoBsMSdgGNdfKNgRlGY/s2FyDPmNDBhlzzYPmXxQoPShCKIIpzUHnIdJ8ENGioKO9Q+ADW/k
pgrQLcn6trVx3zsaf/EURlFnENGSdTvxyqaAJFDA58uKGMuKR8JSIglQYfS2hWcD1VFT/tWdfeNt
mgtMPQ0wr5nb+MNxbGc46YwAkJ0UrBx26WnytFYZ8/mrxPpTLo2ol4NvDA1xIh4tR3OGJRBicgfC
wYGVRAehXQ/9abJbiTkR8lncyHclelu/yN+Mxl6eGLPQasybvqAbg6W9DfwulGP6BS7MJT2QRQZ+
SdYB0hcrAba+AlWtpTDU65TNG+yTwHyLQqozJH7Op8fyp5BYV2W8jEY/SPKNc7MMdQ/BUU0K34BQ
i59yN2HpPdUOc88Cpey5VD3wokWRCZycFY7SsCQJvHs7YTvsYFVP4lOuTVxqbJ1l+XtXX4jFRr/9
QHFgFs0S+Gze/Gwpx/SEmjpepaljUD6vLIvxpfJnq5X3K8uNdV7I3UzZxRQ4qK9POdGBdxpLsf5f
rAVykSLzvKz0Kbv5TOC1IL2fPO3g6JHEL9L7hwZWNaHRjEJzT/prYcmtJUpJ6q8ztRtovDFun37+
mO6i2z/FWLfVK8d6gqY+//UBH/+alq8UtYtq9drgaExvoD6osd8Y9fN7Fo5vf4piaAYG+4ZAg7FU
qafK7Et7nNmLn+EoaSCiKarrEz8yF9B/6ls6md8mRs8VoSbHTZ8g7Wx/xsyvT1Zmvyw2tU8AETj+
VlICfg+Pqi83drCTKps3Q3fc0VeH4Yx8abRPriWmfZtUeFcEGY5dlp9XWXHRGACtuvpkEf717yiq
ulSesY5hyUivX4RWjMT/KYazyB/UV+9OhY3Km66LPEbVBRdbef7RLBGGOZ5q80lIXFM2DHBUjdDI
0n60LZmUgRrJaRLmGrlTKYGnKRrD1VE9L621K8HU7ooRKL2UDAC0Uc5vjUYRFU//SVJQOUWE5SDa
T/uAO5kvpvWeLm1sjAJXSB9XQtLt3QAtvANxnE7fhhC7xcLS0qJKXbY4WCrDUdbyMzUWkAIkafsj
XcDgx5OoBA3SPyno/dwrbg0zYWjWYpxpLS2gIMGtTxbUlywnD2gU54sHDGygOTmxy5MXLpWUBBRP
ffBM8Pg1b7xSBE0RYdTvENGr/yTwHrIcQUGt5mxX6lP3IP+WwIY2NXtFS15ry7aP8UfrA6RSBsC4
kINeFxoCMnMZRldVvLUZ+N0yb2cM7BibnTe4dByW9cGMUJJafp60wtlfrzM7BL1V1WUMy0wMSR8P
fzck2G5vlMP+OD1+Jq49NTh2IkwmghXuCrI7pfNGHelXD1kcLzfoc1UeLmK5Sj9czFTZvakceoDg
K/iAqrG76A14FChDaVwP/Mr812x/hZlSNv+8ay5kFBN4j71g8tU8ROEnMHIVLPckEjLqNaW1ZXUv
1zG1yIaEMHXS8JA1SBw73dq0YwUEtZzFmAuPAfzumZf6aV6KWRbNIat3CeGwP6c9WF5bqhfqGcxh
YE38Yqg+vACpmgjpAkHN2BgyAbuPSCk+w5Rdpr3RJd71s5eXHe661Nmy8CQ8gZOOfMFxAwcT4gLR
AG15nFTAGT83/LE0TZAZmePXiEoXIS5j2z66hUyj3KP73ToF7Bkqx6QFw1ut6ZtTQRVtT8uW0+nH
PHFqnKbBmomh+uyHSo1lVtp1wOwDstdxLb1xwp6+ihCljVHi020tWIym7s2UZWz8Z9TrmSyKO9xg
jZOYc827k555vVpwrlaWsAzxJq6EFmAVWpgibO7LBWoVqMezqDOxa0vEVWPtVanZ4Uc4ne2N6IfI
Rv5wfETbZmIk0AyjQs0UO9qoqfW6f+F81FtskCf//ojRXLGGLEeIvgHUqJR7wvuOokbslE5HId9b
B1ZLRw7OKrEZBHNEUvxYdz74zBmzJ4Xe4cPZz0JHDBiuShPoFJScrJH/Gc7qGt4c+EfIpDbnpSSw
AeDdF+yHTEZE1zwFkPh0UpIS//CsMu/bK7zG4e/CiewNp/7/8W2SxfdV9X0W7apg5lloaTBIR0XK
UMb0dxtLDguWuXNm/P2057ECr0UlwMmCKMqrqP7ycA1BjTIaBBxbNsfM3LwhS8OJetY12BWDvXro
YHPCP6AUBIfo60ufquA8JJrMrhkjUlxem+eGP8LtzwBjl5mc02BiqMBhNhyO2it38y74gG15Uojm
kRv2yTmzpWJ6968VR3zyXp3tqbMS80cP6eT2g+AjR2xZ3TvQnSL9oXtO3ubCRX8ZZtqxqQ2Z9IGp
xG6KQdzavCpUcZq7lzT1qU4Rxo2jHsnsjuh9rRktjVJdB8ui3mmkfIFLHu7sXkA36I7QvZqsDC8s
I+laPj7P/mwIIok5TpZBS3z8QkOOD3lwYPNn3BlspD1QD3TfiUx6Y/+qpNJoMdWknL8ZRwbk0lW+
DUzvY4d18nMmF4AuprCW2Fs/SIIaqSwu4Fr9HrEWFyAJtvOmO312aN3hZon9Xotqg9OhoSwWplRG
cKo4/hD3GEg65f+xIwE+AGqAaHzI5yaOXRKSkseuaoP8QuCWXrGfA+yXUoecA6glxf0KwJfbKpEb
cn49kz0Ow/KebDUFETOtXk0LPSB/L5VYYfZuTeOHNe8xoBVWH+xihbYePb/M3y42ijD1+t2Kr6hf
YZDqJC3i/LXoof9uVVna5C02HVHPHg7sED2s+0YD4bC3vu6Sp5NcpcBKeWYXuBonn3X7/WJRR78T
WGH3D4ijWsrqo/onfhC9WKPnFnZ1KDy137tCJIgpSqM491Ppyz2qBk9fv8dFd9BIsdAn5abLhJn3
CYDTe1QCEF3fuXJFriOuZ1z2KuYdJA6VXpWTXG5CQoHOWk2t2XynRReEsmdIc4UNuTWAevwbdrPW
9T/FP2toAJflncAqd8oez61DZ7ZKHJqTjCrmHohii9z2v4BJvahYDr3S4wrLSwaddyUfRuFpTWxg
tFePtgNJnhffI8hjJwggS0vyOWVH62j/jsk9B/s7OwWqWpI+pOOyvpZLbXDz7tfFkFu1EBCjVRIO
b+i/fDgR/Sm07WqwDbGXMQuuQkUuH6C9so/avx9EdxnaEjzpoP/eWWehYICRo5BuC6d/zcIN8I+A
wyLLtoZfWP89UwrYL9dikwKJNheYqSFeNCXnr7p7QDCkK6CpzFC9FpRc1oJRGuGkD5Fm99nxB0sR
G6lmMENssLMl4yOqJ1Ca9B4/MbyCIaOkyOHB3+tCYmK4kLQKST6mtuooLyGMMWKLdreptsKpeVdq
iByMeecgEYRhWK2qpN5inYzcGBq4WvBRaLEyTBepyuTBuYeSME4fvIBS4T9g/jksSWPwNQZoTRRI
WB4QJnB2H6Mns2bU9qFL00ECLHoUMdJXTqIs3HJPYQy9oj1HpyGSmskf5vmR9JkiInVjqnD7+N6w
UE3lERbC30k2HBQmlFq9PxklQc9lFKXwMqyhl27XsSdT+2ZF+W5wL48q6nIMJ5QlngLZXne/EgvO
HzwqnWcOVMWzcLWXGFP0tj08qXnIMJqgCDeVxXpF9yKhUYWqlSMxTQaHsgtuuSZcmlc1UBCqqqS3
vyy7ETVs7aIXhDy20w8Q/MumeOOletyJAXUlzIihFjLkVdFHGxf1kU2dbr6LHZXFoxfmquJ/BNnd
KBMSHGKG6GdWbAQ2aVNofXn+UGGRWNZX9WEbwXlhDJjWsKnKSjQgJX2QV6UwD5eHwRyGlElAL/do
FCJBsRyd5fbSrQdPfdJyfNSyTtKQ14TJlrUcpGqF+xYskeDCflsYEbdFjljBaLHXRejL2ZjMcCTj
i3cSwaJ5C9xgTgO52brnxrtE6fbC8Lk/HwzbQCgxQ2GEBQvHY/94Y6+SHn3keo5vjZ+DiGgww88U
F/CuEY0rCE+KILiodKn0gifUfUs41OVS1qhpyqenDsewlHHR3UCQMMVhPrLv8aSCLYcR5+8bPpZC
x1BDGqGhK8+sSMylDfgWjz3AQxbQh7O/8/dH+juDzRMqoK/7GwoL7b2ZY49KnKkzSjdegwfPG0I2
KMSHxX/bJi3uVIJWB6LYQzTS1VQS0h5y1qvBmLyZwNdXQx5xZxcwB9xG/JlB3YhFAidT3LZuABly
R9LAQNnL+rDpeRCqpeou+GHAlyByI1ES8mhp1JQZ+RjZ96SHel8lXr0UkFtY6ozuYGoCjBNt8lPX
T+/3OLo6vaj7Uo3R1M7Mun54etsWBZCsxK2nYOgqJx+RFUcYzJaSMAvdo3NK1bOKl90UeHtjWqla
bA4T7o4ZCUgcsX+kuEp9hEZnBsGJvr2ogVFxBrKl7am0yH6ZeYqEzv1KeUiXDFWeZMxNROknZeGy
Ihee8gAYraRYHI8IdiInRssJ7JhcrMyds+Th8oGEakZCjkC48+t6QEFif9XpXDPcaf/f8Wn2Z1pl
XZ1+kUvAR/KLFwu02Ptw56tOs5W3s6DzGr426EL+UqBe3r/uYJGiWXLWBQ9jgrvwWW/Op+Cg6ThG
QHMm1u/3dVOSrgsAdY/XWn8O0FSo7WU54fef/sf6SjzUaA7WT5jvYHrAtSFXpPI0WFc//yrU4+s9
70x+gd8dn9r+jOy+8XeepC7zvFowmU4w5cBtdfjINAmvbdVl7jWeG3xDOvzHaXLCWXieoYRGjuLm
KJUa63K6pQFZmfIx4uo1vzwxSY1BQG4mUUvmYPpZktLFvqNuPHirZPHyo7/nHHTq8X1EASP6FXQl
yI7jlnJCbK3SVbKB6Mb+4uHW8wDi0RpzwLP1cQAynoAzjPcRTqOhRfCRFAeu9KP75MsffYMl6bsE
w1V55GrAglLUbwRcoq45D/M2FFDDqE0vxtPEuuxH0ZR6BBlpWmRxSWim18rJE97t08UZ+KuiD34H
TYX5EyoNX6g9YcTgkAeNZnIuNmBAmvR0BNTMq4qIrx0bhCGpF15j4DTkXmxlDL9/zmPAZ5Hn7fs2
eXERpx8agSFgQrKw0faSygUeUoVQH5hvhiU7X5Fles6x6WqUkRSxpUtPbyZV6atG4ZwruAuHlO2I
WURA1456SR0bnN3EAozAqIIeLrzoxFuEtZagDNnQb7b6xqQZN4qiHZB5GM6VYtac0CyDCb1o30if
S1N+SDPob8XkOSoSLgMuS106Wg/+XrvZgkjJWC91MTc3ydCziDwhtKi/B8s4FWRtYY4gkMVjsaIv
W/5K05vPVz4wU+tGjp0S+8ESSrk4EIgXk/qLu+pjpX4XjE+KZklrsb81f+aIKbSZnM2O7tVTf8eU
5fx/bVROGK1YQaXkBY1fbkvPvobsYSjAseZzip2cR/fSHzY5LeuGwW2JzxWj5onUpo+EohHEwfzU
v9Goxa4Gl4QumzyvTPQRllamCw1i2xDTpY2XyhW9Gzt6XsY8i0wgOtxKM2kJY1Ssiy5O2XqVtzil
+oAu5rdAVI8S+BEoGzn68R8gnzHEDJkchbILIRXagfZg5pEzYlovBZmUwKUNEteK48IBr1WchE0A
zdrXmmg/hzXz1vqk4jPfZP51q2qIOzSh/CQs6J/vYUh+0brJCt45ixu0pCIcwdLHpznyvk3lBJTC
wjHXgU0MjuuJoLNLy6Dng8cp6ueK8Ppccsa0plTqXASJscQAJeX9CEu9KyVz//s9VLdlHLE8n+pE
mDQAU7zDYlaLe1YQHR2YZSJhex9MplTTt6s54748VisMqZDkb479bRdU431eByolgucy9jxP7qd9
Zmznhfq0ZX744UFJjYH+6olOT3jqIhkaWdjTZjy+DZER2qDWIUSg9zTZUHKLXXSTIgbIvagddB41
6xSEQi8X5+gC1KTXuMkLAFOF53jcvv7Th8wmk712apekJD1H7EoK64LwoFfZ/473W1M4U0TlgiO5
Mery0JwK7rh5Yb9n5r4MVpF8kTigpNImyYjBCUMnxppKZIMHAI9T/ZtXkDsT4R5YGYwH8E8y0Ojh
DZ+1ss++A9xByScZCoA6IU0xPbVt1UC7Cc/QKGMMlYps+knhYrgEo2R/qAV1VGeCvlN53sRUVRDF
0R+3iH4rEXbJOAHXurLDANJOv7CKQR8w+Sh4Ff8ojrTiklNpzLwFh4mXTzIXb7xU85zWIF3nwcoi
Zw6wOF5iEWmDMXNhm+27sVn8mt14f5nWG6k0WirGCYlDkTqtfXX367sTknrJkZecRTiZZXdfXf3/
5XHoyx8ATMid+d/D5COnuKQtE6GQMtmJHLrShzIqLGa1iEp17yTpF2wY2C4wwtaabUP9NiimeZLe
qoqBT779lT0lnr1fazWvf6TFCe/EyNlY5ffNZYOh4nfoWRTugwVtYGDwPXfBBb1P42kb4bf1h7+4
Sd42HV5RVTCBhS+fR2t0SfzVAgoXl1gJ7z+2oP3eYEIcg239Uw7Glbae6TC08k7fIW34kuzW3Q7+
X+3ar+giXHxglyiythkpU2MohKEbQwQhqpamJAbLz6NYmbjOvDzfLcGGSq03w4YS7aRV2/P61yKQ
5geTsnvFv3RqT4DMhDUx2JcjN12KLwDFU6U2yeRn+C0QiJwQOZfaOofL9dVNr0agu6z1sQLXFq4X
z6OAyLO3ZoTzHbZ4PIZu/FU+Bqltqz9aaxc6ulN3wwvBQOczJ2AkbWc8Hfuo/oqH/1RhzA3MO4IN
GmtHG9gwe1Cdf/DvvpxXnPx1KKoHnYJv7IbneKi5UkYn7FTVxwkxR8MTjkaYpEI5V3sTxkdCAxzr
k9GwnZ4n1h6NKod6Hsgccnak/GEQ53VUbJToIGR2aEj6TfVu22hfjttPNtD0NAlLvz5PFL0+shEl
duTKnb3rXnR+ukXW8SYrf3U1pEzqjUGx5oSiQ90sXyCMhcT/CSy1TfHoTO+kSjpfjEVRCrKs8TgQ
yTi6klHEsyXKRSW/FPwRXh3mqXU1yixOiX9obmwfp+zmIYJEhnD3yuq6HXCiX5XvuWn5dcKNkHQT
Bh4/m/p6SOVIi+Y/UM52V/+09USB/tXTJAmFk6WQtkLZzgwreRgPnRaSDAfvXttfBDJnSP+ba1wU
WwTkXWpm6IHoxq0UHpYcLoQH4UEht4OKilbTjqp3+oxa3yDQH9PSI+WYnNTaxMkB7Hk1cefO+1qc
twyM15cSq/YrjrLXVVGbAJs6thM/RFfg7qMFFbeICKg13p/kPgTCwt0cfzI7CyGOQRW1f5P6LU55
XmQ9GNDG3qrMx7s7SyOOD/enebHKwwNHkFu8vIxRqUmWmoOK9rPD3oYuklAI/YKfY9TYijxY+bJC
/+SCJYvIWiK1fSYKFW0YloGGzi0n1OkWJmyn6iGNVEMVzXGif1uakcgvybGIUuiYMrec23dUGGz/
Crx+SNET1XAtoDKPWQGq6vt/gNQObNdD+H1UZDHIWkE03BrYolAHypE5wKk7Yf0q348n6mHL3rnF
pj13SSChSA8s/FMqCrLoKaaVUPkesL/FQf3bBZzgQ4wqJ6uM6ytFmwFg3jeLMhqspS1KziLZXqhn
388e4DlKmhBmJ2LXaf5lbUx9iMo1qVUZrlxRgvzq0Yu8Z2sedNexCd5pYuqb6TXTmTBfy/eHpRbd
0vYNeBRLfNspnplRXwAPoA3ZSTJWc/tSOKe7H2GkO3AVA8cV5c2ALdgl3P7iR6YfsS93Hvh9hlbI
Xy2lcplHCJbRfQ7isZd243PsGtwLcCosMQSwBSjFgp9rvScloX9B4cN4AvYO4LdPfRlG3OBlDdup
yy1U06iIJV2LoDrU1VSHNDyOg9RWHqWum6ZTN1tl5yn4rDxMGOI70TVTa8SSGzDhBTzynTnQy6Ns
Ih/RcAhh9jlsJ0ym+nEf9DztfqjEMVNelCLuJNE63+jRoL3v/Ww0hOptbHPxE83GoZc5X1AGDkaH
zku2xzpjNcLFrB+zlGnj6wLDLbhG5RRfaFgPGsDq++0q7EFMK8dclm2q2RPV6J5OWx5bA0tRCNLL
DxfW48aeeFr3bSsgcKeThkYfb+aoaCZqGpITX0uMy7HzWye1zf+/1pFcP8W4MsLSh4oGa3EG+w52
24wYL4ecQ6pvzYoY6IGMp5YIugCBeExmiRzNhDPABLrt32w3KYgAz9N5XVmBksG8O5TU+iyf9TIZ
vSfaTRP4h478ZH17cHcI4wDXRfVhCXb6boXCy7R3snh7jo2zSMJxoRvGcpTUKx/M9L1VCIIrHdrY
/ZRYGoTYkQSHWNW5gFM3v9LnGb1LuRoCWT8FJhtTRCjr8PkSfZppsQIYNiYzCYZwsQXCcHLdHS+y
ine3SkWr8rFkUAStPsQ6Okx32F8GA9dbrJeriC/0bFFRWF0HNyAYRQq43b96qVx7DSd2KglzuKBE
8+aED6h8+Y4Bkex5ro/WCBTphVCKjA/Qj5W5K/sxxxIyaDMr65PB3o7PfIh3iZqikyLiNeE2ecVi
17YKyjayk+eEfHPkrKyBILhRzFGDl+ec9L7q3Xvvzy1McEBahLf8qCoRV4os/qHpUhZBldrhwSnM
KczEtQwTHKv4fdIdcrxtYxvyAu5eOyecg8KpwPi8W1Yp9IuSYl1+67ZN/hUCGeu/kATdndOkUPsv
4XlSdUnk0VCYZgEVvjsdiRlE5J2hBO35DFKJCT30ryiY2c6VmDyNXSPoNrH+V4k3rZpsKd8pMsWo
rTABfdaOV16jYC0qhGV8apxJFJ66J5EUFdTz6DLAtKOJhN8plol1jpTQpiklybNXz+y9Zzg2mGaC
8krHzMcViCydplpoypvlvWCvvT+EWrfmcFX/1i/SVTTWd1+I53tXrGGChz5rg1QQ9brXDrUe9jbL
C2gSdH/2UMuUikzuMaEmGnVd8lV4BWtcWJsLISGarIKU7OcpDmzaOlhCPwgpz8eBoWnXMXjufQHb
nlWA7i+GcXoJezK9+JlcFD8LUBjo5rzwhwDOQFqVcxi6kH8pxGf+RkPQyQErhCF+POlvu7NlOYiO
oF27mWjUqnnJtahOqqh57XhCQ4gEmullPiZdnKQAXr8S+btp7h1o0TnwfcfeDUZtaeVxCQi6WyqD
p+QYsp7wFjNWv+3uJskJ0h+zzvS24Yo8KF/CMnZql3s1x3Zzz3FxxKY4G/Gr2+oUqgYhhQWTJGSi
qFPmBvwaOIqQ5UHAPvv0YJMiY+76K8lk7YcRjSacWsXlgA41rbYOKAxB0p2F6F7lvMeAnqcX5Tue
d/spOQKghk7tM2RKjKAui4B9WGWBijPqA12hrwpf1pBy4MvMy3+TAKbslC+NXCpyOyQ+
`protect end_protected
