��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l����$�8��� �-,���#�bW�\�Zr����]�xi=�i��[<T����Q}�(��cr��5y:�ʧ_o��G��v:����`��a5^J�)BR�7O����#�S�w		��v�-�H,*T�(�k���m�|��R}�*�DR�Z�}'��Q 5�O+F���qp�9�Ԫ�j��|�Dv�#��Pc�,�2{~ym�,ic~=Z9��-*i��ɘ���1{en	��Na�wd��!O93��[X��}�Or��,&�h�)�>N0�Rw��NL��bT:��Ȓ}��&���	�ÆI��S����X;��`��yIZp���s�R��Lg�e�ߟ5�$�	��:�I�=Z�F��'z4��5o艞��R�F{�xk���>�Ϣfj�w��o�np�H�P��q��m��I�ۭ�͝�O�c�d�&�}y��T��Nh8�0�R�{�|�S���*PF�	߃�&��D符BAr�J,Fh|��%|��Y�l!��<h��bt����o�&�fئmY���{���p�i{��s|-�@�$/9S���1��T	��dS�O���3w�q9�id�bBVȏ�؄�?`$��!��iɰR�f:7�F�G��P(���b�稚�t��#fi���y?�]vpyE�E�#?g�>���V�u8>�B�	�U�u���f�a���^p�$��6�f�sC�PeRK�U,&<���۳U9��@���;Ln୘�����(�\9�ݽ^�h�r6'���/��A����v�h�iص@i�@+[�5��KӁZ�Q�߅�8�	�N���k3{yk�{K0p��?!�=��.r��
���?�t	��w�����2�5��q���88(���4HÏ��i�'�u��#{~gE��c������&UV����.����v�u&'="O�����3���4��&����`E~%�?b��������ys�e(���1��|W!*�W*�6E|RŠ3T�0�F[�EL�aTDc���B����&����R��kGK�����k;S;�l��A�������ݠ�������v�d�6^���� $��7���ǯ�����z�� Y�ҙ��Z!�q��f	O��(0������#���\�aan�v=��M����SLV����p����D'�q�/]��V�$)}Щ2Uح���p���*�^�V;)��;o!sb�(��(�\  ��䎚�s4��=C�v�yx�H��6]��p˳�����F��n:~� D�9#߲�
o�h�q�/0��0��p�1���z�O�0�}���R�?�V�ҕ�cؖO �Բ]�	bK�r��ؤq++�q�%��9� ހ2�J�*S��CJ��ц0c�FJ�� w�I4�&N�8@����m���{QDkxB�.ژ ����k��QDE��3��1hw�����!ĉ)4��e���%���� m�t=�B�6�|��I�˼Ջ��Ы��R���-;�C���" wp��/���Tg�X����'(b?.ə�Wl������8���~�x�=�!��v���d�+��4Z�J�a=@j���v���e�P�E� 0d���q��u�k�Cr�;2	����D<k/��݌J7)��%ņ�ې��g]9k�������7���� 3���G� ���킆Z�G.Srn#Bb��
_3���������O�)W�[��v���Ṇ�yP�#l��u��ZUJ̔�.6����)�u[E߲�]p�H7��}����=X/���zҢ���֓hF��������KI�R�+�ʹYN�&����R4��̃5L����2l@�g��8��/
O0�M\���/iX�T���-;1~L�1��Ql���w���^p����j����?uB���rr	�y�����\Mz&�xQJ8��I��b�#�G1MZ��Y�OQִ���8ˑ7�}��@K�3
�N.5� ��9'��JJZ�Ч�Q	�����-[��_NcX���դ�B8#��i�S�[x��K[/Y�JfS�_�G�ĹU���Wę̼�k+�/ɍ!}���
"�O�a������.�%qK��q9P��M60�3Z�\^�L� �$���Rm׀�[`��c!�^1��m=�_��3oQ���$l�-� W t��7�:Ǹ�?H��d��ٺ�kҙfs����P�ﶗ�a`H�XVk��,��J�!K�n]��w6��m��:�����h�уg���1�3���C��&���eZs��9wk��u��,������d0)ŕ��2e��.��>��TƒsE�:;�ق���|�Cz��ɛ=���7;���*f�.�����E=-r���-��6�rG��|�?�X����8�!���+զ�K	8N�`�E���G�;�K�j�����kGu�	3�j�d�a-��֎��b�@�!=�ڳ�pd]��<��B�,"�7[�
��~Կ�ů)�@��lh�RdD��	aE�m.MOr�*�<�J�d�U	j/kW��>Pe���Z��L�ǆ|�#$G&y�G�܍t�&��$�-����^��S5�Np$��r�D�^�%&A�r���;a�6(��� �kk��@�4qS�hOL�3�_���ɷ�AM�Gľ9<�#�L��2tV4/`������ɔ��o'R�=
�c�]A�4 ���WKSt�x_�0���Y�|�N�̅�= �*�˟�Ǥu��%pN¿����L,����>�NY3�m���^@�rbܙ)�[ʵ�Ѹ��7���l7�ȿq�aNV)�%��ދ�����M������;�������3B��-��4C�ߖΓT�lu&"&L3������G:9�Ye�
��<��4>�б	x�V�[�7D�!)��g�]����7'qxB���R#��wc�p$9>��v�s����7��_���>���]얓����yr��;پ!݃n�l͜��$��|����4/UpTG��*S���\	M�I�j���+��Fv��W������`)SP�=t�e�YG�(3�D7�4<�<a(6|�>-��-�_�jT0$��%I������ٲ����;zD�} ������5g�f�ԟ�im����5"PC9������Gɑ� ��S.�y��@��eb�,�;�\	��BG�])�Q5��Be���� ������-���#ؽ����/����4ng���f9k����';h̦�-g��=����R\m�t�#9'$>(�}�um0z��c��P�eh�_�B���/�Zɯ�\��*�����[Z�1�K^��
&�d!�(ڬձ#�@Kĩ�VC�n]���y����:(>N����ʞ5�l�n��(_�ou�d�TrH�Ȍfl�*�U�;�l�8�C⦌����rb3Cve�{g���F�\S,�U��M��腟|��:�YIޖ錪7�ba��[��r���$��nd_���{��5t����PH�g
��CaAG7�LM/��UpS�~�S�$vK
��0Ef�F� ��5k��F�sf����N; ��v������fDc�G�#L0�'R�w"�#��LII�����x�rT�@Ӷ�O��y $���a$@t�G��/h&,]��M�7k�^�E�z;y��6��y��0�0��_�D���H��~�ulq�v+c�l�]�7���mj��j
�.O5��,�䰺]؎�C'I�9-�kk\�����+V��
ч��+���e���,l�~,�
H�b2m6�6L|!԰�M�;ن�J�P���ˇ�M��F~��.�>fj�5C��^qk��C���͛���U�������Φ\6\!�ϾJ��D��7֨�K�e�aH̿h}�e0Ń��<~��ꄸ�g���E��O	<b~�h���I��XO��0$X�S'�q
�+H���m�_p���$�ִ��w���/�r�&��))`b*Z,D	"���vB�j`�8q�G�j���s	�oe�w��|��#$z��0�Nw_QUaL��մ趫��I��k���$�C��s��>��)�}��Qs��Z���T��U��A`�GP����uAs��� �p�X�j�Z)"��5D-����ɳ��\��W�m���hd���)�2M����V����;Ƈ�s����QF��7�B�)���[f�
�IuT���-�j�S��0@���8G�TL���y;��w��t~/��]0iA���?��ˌ/}v7l���Z��{9b��V��c̇CF���ድB �$�}w�>H�2gNI�0��<���5��n#o�:��L���<m�Ƒq�u�-�H:�����d���{��b����- c �
"Q�"��]̧���<��c^��3x�٫+e����������"\[��͏�D�a�O9�N:�W�M&�U�}��n�^{�O����.wO�Խq����\D�KL����A:��Q���i ��`��jvy�V-��30�e ���m��h`
����1�:�y�I�����A�گT=HS���\]��V��'��O/[ЊS��89��J�I�jp�!�ۋ1k�]6E��Vn�(�� lo��8[�С�X �� }����Ha��ВD�S��f�䙋Xo�����E����D�r0�e��Q��Y��YWX�	]e�<l�/.^�Py�K��檅4��%�*IDB#�4_V�|%��4 ��"<!�y`�3�'�\,��2����_���R:.n�k�Y�YVڛ�x$��?gD�Yi��du)�h��ę�2�vI�╊J�\�"�`r�ž�),� 
/���űqΟ.�����������y��;�6Zў�u��6��~�š����E�8xGG�����"�
��|��Λ�J#���-�m�÷'uw}��U�x����V!���V߈x�S�K����]���Y�E���_�����y�	W���(�y�B�T�6���3�	E���w�9{a��U �w>ſU�s;>����.�D�4kEP�i��J�8l&��5MD�"�-�V��ͤ*(	�S�,�yv7|�պ>淿�s�����������<��]�Ca��T$�*q�}�{fd�u������62�>fX��t_�;5gb�P�:�<�2�v�(B'�=��3�����b@�<��G�y�r�~��/J.2�j<}}ŝ-d�'�fW��п�b7[�+L�e�*:v|�B��Y���F&���F��%��^�0[*O/w��^7;��@Y��z׉��i0shx���:+���^��k�+|�I�aFX�*����z��_��Q����,,����t__u��,�L}�-��t�����X�F��tlK$)4r��U��K	{0�H��A͋ߞ�*�-�.�5�-��pQ�
?��x��,(�Ҥ�yq�Y��|�&æ��'�tiz��@�9>S-���Blz�D��X��_��-Ƨ��_�]�*���S�؃%�:h�5�����St\�bs�����U?�@3�՘�+�{,\
x�� ��jY��"U�6�'�d}�����[W�i=-�[ܛ��6��v7����7�Q�O���������;H��������/��o�M��ٷ��K*Ne��\�T���?�J����6k�Gw��˅���.��D03M�yzl� "W�F���i[�!7���br]%�Đ��.@����9�.(0�|�L�
y���:�+bs/)c�aZ9���7$�m�g��3�yA܆�7�A�<O�Z-�Z�!l}f�|dRݶ<Q��G���-�H]��pq������� ���S��p�ݺ5Xj<�����T_jtDZы5��NՅ7�/��2�޹���Z��4��1$-�$���?p����J���*XL��k�L���Ìd�I�X���mR��#���;i�`G1�eEg�5g�m.��sp���c	��nپ2����Xܒj
9�bW��`:�΋+*�v¤H�����GMc�A�#�q���S�k���R
��mr�?��ǥ��+6�"l��U�x���^�6�7�[�A����P����-8(+����7��dCB�0n$:���1C��?��@\����'gQ�z����Xُ|�]��2�|����H���;y��&�a��[~�V)�7�D�<�bC:�Į�,��s�9g��;�ΟlD�U� ����G�@���)o��c�G<�E�'g[�2|m����Dw�F>�8+;����f�i%���7 9�4T�b��I͐�oΫ�l�4������*��"޳�~��KR���l(���t'�=#NM�v�Q���q"�0N�[=���q] j"��3Bu�I�-�vup���������|��l��v@#!m���.�dq*�� fC�� 8��Ŷ��Vk#שYk�t�1H:Gқ�-Q�&��_[-��/�n�y�� ��pV&�����D���z�{�+�0�U�0���=��Z�Dx퐏���^ �3H �:�HD�"�J�h�5cHj3m�:��Z��C�+�P�k�d'�t%JU%!��)U{V��5��J��M�<��#���
��=ōg�ߺ�5�J�*��-�@���2���[�훂�����m���ѧ��S���P]��g{J�ˢ�g���O'���z���'��d8��s�j�Ɠ �K��uEm{�K��ꜫ�pEi�{���!��L$l��&��'�9�k4�#��r�{!�����`a��V@n�.�� �Be�������פ��ɵ�3��k�~�H���8FI���� Y��[�	�P���Y̓w���O�	�)(�1� w�]����@;߃qB���(�$w���S�v:���Y�^D5���2�P��\�}��w�py�RF.�#�P��QE^����A2>�ڤ�gPs8���z�;ya7r�G<�h���j�H�k��¦Y�n�8k���P�tt��H�*�y�r�dV�	@��e_�W����&��Ҙ��ZO�r����:[|#�Ź̿5�A�:ã��{���Y��^'���mQD��5��1�f���߳�}��+�p��C�{����;����~�H�G[�N6BC>x�a7�LJoP�1|룆���+:�ι#)��B�5���$́�g���`��"p��2-�J����z�1�A7�j꓋Ī)�,3���]�g�8:�p7}	��y��g��IͿ�`��H��ihp9�q"��n�,��s'�7��K�'���8�1����܍�P,�2S�~�����[��K��5��y�۳���b~�3廊-�����4+�N���I�%����ގ�̩�&S�����Tb�BR)-�5wNT�@�ƪ\�Ҩ��f�ҋ�,Jr.��3ln��m�@dU #��"�P�;V`p������#^�C��sn����� T���'��#�jr���5�W�
�~��V7g�8kh.?]���V��ެ�kz�u�jgjǈ3|��J%�J��_3	2ϞQ?۫��;���]�wG��eC`�ּOq�.�=�h[L��a���'h\d�|7�Bu�߄�t.�#}�r'�C�� �?���cH���"	X���Hl61��҇Z��~����i�o=�k-+_�%���w��%�*�糤]Mr"?c��j���۶���B�i�O�N�/Q|o�%�o}IRց���;:�Xe�_گ�`D�����W��b�5$kP¸��K���da�;�K��<�w��Ť��M�n��Źn��� �� <�<�
���J���n4�g({�veu��k��v�@�H/�ZƔ�ٽsr@�����:wL�rS���@�KW��^�)jv�
���wc�6�D�����o��N��oq�O��*_M=Ԭ
b����V�Nf�37���j^U��΃4mm?�	,GKۂ֝������H)7���az�$��N�~�#gyf�tV�H�~[�#��=�D7�G�dA�+0�� �F��o�`�I\�h��&T�6׺�i5���"r��U�ͦǮ�zc�[?μM�]�(�xO���w���wJ�;�N ��>\��=Q��͂ʐQ�v#�J���삡�Xݺa���׻z��YNS�ʍi�P%4�Cĭ����f6�/�G�Mף��k��MF��;�f� ����e����`#� D�eŴ �BHuZ�IyR��O@V��2�CjE�XqV��B��
ptW�݂)��d��`J"q����=Byz��o���_��!�hi1��
������>��A����w�5�d����4Rn<��+����A�dd�n�8O�����ب��l��ǯr� H%��5,���3m�1[[��&$Т2�V�-L`B(m���� |ߞ5#�u^��n�.~���y��@b�=+@|Y���p��9�Te�����3l��ڍ�}���(H����K�T[��p!���Q�晷:�� �`#l�����Yr�>���͑i���%��@��̛�G'��|wd,IŨ��
�ג|O8/A"���(<b:���'�����8]�'#��?5�h�R���B�`���SD��o�xk��_�6c�e
��4m����wm�Q����Lu���)]�0�Y���\�r���D�Y75��B�p�MMX ��4�U��#�WF�/o�eﹺ�~�o�~����^�]8P�LM�S��jI=�%�*��e���^����|����x���K
��x��eaY���X��~���x�S�s���h��|�߬笊Xtk���D�h\];Ŷ��k��bN�V�?���o:m�n�LS�����We¹�B�~^��c�x֏-����:�d��$3Gm�iR\��z��x��gk�`a�&&�X��7��^5d(I�,bw����
�4��N��]|�0���h�ı<md	�B�K��t����e���_k����܍�k��]�i�Hꩍ�-�fC�Y�3�-s��p�Q�b���w-;2D�f1��pw���3�;���̔����T�q�v=��q_����r�)_����Q��4L�A���E��=�e.,�e0��*
�&�c�ᢳ��k�'�/6W��]8M��V5�-�a�`�M���d�%Ε��P��~+��R� ���WeX�u��V\��+�F��gElaP�O��X��Y��>��!uxo�;1�"l�%��'p�(�z�_�`3�A�㵀�8�a��*� ��HS/:�%�y��ZopX�X�N���ũr��x��{m��Jh�x��"{ٲ�x��-�(�h�bu	y�}7-Ol�k�	�	�����cñ�]U�+Dd��n��m��D{�:��:闤��~W�`Sz����2晴*��^�X�7�>̉rӀ�����G�yջ3�Ư�JP_�ŝ�T�q�$�~��-'EA�j�y^�r���]`�J��ݷ��y!�"4Г���Լ�~ש1���ݦ��哯����v)(�29"��J=���1Ҏ��-��E%9��=�X��V91��%]2�$�=$.~����7�ZH>pݡ�xG�n��:}X�7A�b��fX��$�P�&��\�9j:��jK��k-l_	,/� �{	-��<bqf��(��ǭq���t�>��_�:��VOh�L�噚�1��5�:������'��lq������۰���W^�G����+in����|�\ǌ���1����F,�mن)���rX
;��!o��dX�"�@Z�������r�>���~g_�0r��z3��5���i����}rEU��z�����<%�2��\P_�#��B���5��B�-ݩŃ2����3�r	u�;�d�Y�ѵ�`��:[9>���:O�!U>�3���jDk!���ڵY���^G�o�OL�����EUG����BP"L��?x�'t�3;����
t����H�so����D�NP5m��sjq6t�:�L��E�\�s,���iO�C��;� �5w�_�v����r����N�����"S���wͼ��1ǰ�63��
@�d7WӾ�u����I'�!������1��~p�+��Y��'��i�u2H0ސNH�#t���wO���^�EUD�^�!�>6@�X.������S��U�o�J(��½g8zg�ǚ3��3�B�W��9!��7_�(��C;�lLq�Kv���;���*Z`��6�� �,mZ[�У����{>���H��ɚ�;����x��w	��h.Hݶ��H*��z�.���{�[([��>����D��G��e`8d��0l����7��>�w6��_w�̅��~h���)r4��jH_�yBΨ�b���WZ���q�n��xx�w��Q�#����Z�����=�cK��m�@�S0ў���Rp�4�e�j-<��A(i�x9�b��SS�3z�c�pcж�ɽwԵ�+�BS(�ej��'AG>�|s�.�ɤ�B����m;Xh�KMm��!O����T��k,݋�q\p;q�/q�}�̻�mV������^�sg)N]�0��r�d��!�0��M����"�ۊ��hIjm�$����u����M�pAm���ܹ|��$u��c�_����m\,�`���4H�n ���bJ��]B1nɦ�ɒù*��L�s�*+�������>(���	`�>`�[�72F����De��r�ã�7/� sf�Y>G,tB�f�N�V�
L��
�B�o�_�*���o;�������s�Jʤ�٥��� ���UnjC��@8$57�,�=�aa`cD4�b �Z����Ѻ>�O���pD0�z:r���F٧��sOĻ�ȋeI�qzQH7r��驜��|h@��� ����������_���F�k;��݋��۟P�6$Bk���L�p_��hL���P���'�&L®�n�¥�-梸)��/�=0��0��B9����4����
��$O[��IdC���	C�V΢�w�����9���A�(��#�2T�[��\99��7}H]2.	v0��Lc<�/Ii;>��]\7�
�3�TY� ���+U%fm��#3��2�R�K��6�K�Z��1Z6M{6�óÓ�3!�m&� s=�� �^u8|@���LΕ�[U�� ��������E�l��<T+�
;���\�4�p�!���^���'	l��b�~��)�)�������ͣ�*]����\�w���=���_|�#4����<J��Ml;iF�Y�+8SlD�,�zY}��c���/>z]��X���TZ˳�}��yu[��^U�wO�'�-�km춢������\�CBQs���ÆU�@o��	�"��^�C;@5��lڏ�Q�O���԰2&�3�׾EPIg�}��5W[��(%+A+zo�x�����F?�8���}s$�|Pf��G� �Ux���U��5����K]C:?���hA�q��g�AG�������-��K-k��
f_��m�!�i*X�1Ę���{�%mvr��TC������k�4�wZ��ٟڊ<�ZH-3��(��o��-^�G�LP@3��;Pl�$���b۫�c�"���]�S���3g�Ұ@�W���}KC��"L�W'h��Lڧf?a(Eh���4�+�kU��&���\�~��ʓ�ēh}|�:�V��\W���!"�?�TxRF7Bvcy�X�Ϙ)� *{�QK���M�xZ��w�N�#<��-.N����u��T�$hfz���NO���I�����}2^�U�Ϝ�k~��y���(�0�cg	��'i�G��BT#�(0�!��cd$B��U{�I�p��HU�CH�nR�Ũ`�d��J�ظY�����ף{Ս��W�}�Ѕrڟ|����%�ޟT�0Tm����D{,