XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� �ř/����� ���|&�luiC�'*�r�D��E�f�Z�>{3U4-|�y�Jk��pr^Gonu�[#�����^�_
�u))������ �B�k�����`}�y�:�ܒ���mv��� ��xn��
+�F�C���6!:��-�&��0�|P�A��p"�U.^�w��-ơz���'ognڞP�o���F�6�PY�4U��rRD~y�.����3���bi�l\�t�p㡧����N�����L^)	`&{��`J�/��$l�|����f+5��`R���$����.�p��\����{9I��ey� ���8)W�vw<w�',�\=��^��YL�#����)b�v���BUy\�I~�8�Z<��y�B�f���A��\(pls{���u���lG)O����{�/33�v��`?~	��G�����<=)��Ҙ�b���u�j��%&g�e/�7^9�= ��y�ȧ���n�$1ӳz�2Nq�p 5B )�ޏ4�����E�O���Mo=q/K&Ѿ����e(�_UO�3z��ՋX>�ap
�K��g��˼��`�s5ٕ��&����7�Hh��4����W��~��r��ߐ�P<�%L=�l�k��Z;�骗^97ׯ�
�:ގkx���<�0Q��z%�>��m5o,w���T�*<���-Io��]���ݩx�i,R¯g
�z�X�k6�|��2�֕�l]�d8L��l�$HD?3s��;���K2�y��Ѯ����1��<sN3N��Ò��"j�\XlxVHYEB     400     1a0�� śPμ����������cQ4�����T��l�S�เ*�����I�шg*���@BK,�#����_9K��'����3��cUrF��یiи����}o;��wH����H�YSwP�K=jz<h��o'��j�(<�IU�V� ��C� a�E���;�6��׵��ZB��C=�����u���Ǟ�0pE���<�\ȭ�gd�������OZ"�F���*�����iK���� �܈[n.+��`�s�tjK�(O9��+�&���S�H|���Q��J&G�ȯq��ď7gTv��͑����C|�
���r�������g%��䬕ƕ:!�ԣvW�%��4B�6����d�9�U��Je]� �9�:)�ޞ���Y�ҐՄ����������e���XlxVHYEB     400      f0��i��3����_4��Ԛ2��6�W���2�F���i��6�W����ԭ�h,�ohuȭ,����,� �'�p[?s{�u}xq7��(5%��2SF��ЪUk�h��{n��>�����p���n���7�K��)�1�0�'f�l�[��֚擑+�K�X��	31� <��b�Mg\���>���.̋/���Km�t���u�JJ�$�ulz�(�gxRm����B�DI�d%XlxVHYEB     400     180�^w
px�!;�>�����D��"���(�I�6�j�l{f>K�+ �P `nX{����4;� �(�n�ȅ������U�M�`��NfUg��.]�<�o��@�������q�`/���J���%��=�"� ���̫-����$k;�������k��M@nϞi�dOO�L�̲<�\�t(RR�
�`>��������sM��*����(����T�g���Q�MY����aȽ�D5�lM��)�x��]�`�u<V�t���w�4���Y|nܗr��Bȫ�W���m�U� ̞$V�b>��B�Q��Z#x�7Je��f�^&bޑ�8w�|���e�dk�δZC9�nl��)�"��<⅕րY��S�ަ��[����Q<�Y�C��XlxVHYEB     400     230:��O�P�-ۦi��,�}�Afnm���ΣV��e8�J���\�(�g�)8Qn��]�ũߥQR~�?���׬=�R;��.F�}�\O	���Y��p�A�B�F���f�/Rh*Y�~�Q�_��Xۿ���)ax�/}�\vA��1ѡ)[�����'a`՝\����j�<[K�$�{o�+�s�Y��0��ج4���H�kĩ��N�ɿ4��L�O��ŅI�aL@�@�b�$h J+�WD�e����Ӹ�.ֆ�0ct��(�@%fƶb��Ub쒗 ���T�W���3-$Pz��Y����L����i<g�YX�;%Il��4)�r�~�\[���Db�Z�f%jN�t��k�U�"a��9��0�iW[����m%��=��'޸�]N����kR=S��&�X|��@� |{�vG�b�i}n��V�t"��)���"�V<�v*���k��-ٰ��^�h��EVm� ��\K��2fdw�m�T��+w��t]��x�7>lA�d��o���D�n���)�ޗ r�����^��lDXlxVHYEB     400     1c0�7?�3g� D<٩뀡Cq���Ql���_���2RD=�>k�X�(q�>�q&���S�S�H]��R7=��U�0  �itY��X���E���u4�`4��eGue���/ө�s����^�Z�"�{�| ��~�O����nG�~O}=��r�X�շN�g����X@g�*r��H��r�.�ui�̰ ���i�:	�ji��W=�f;�[c�/v"�G�I���&��g��	�r�˳�R��jFn�ڸ�B�G[�=�Qd��L��u�!CL���#vTM,y�.�G����z��w9��xn�ipi��pGMoh�M�?���ï�nA�҈�A������6gIf��m��ZF���8��
�Km�����ܽ�xg�`�t��g_��8�5��,k��$}d���ww���Y)�O�����,��-�������P�z��b��+�ȓ�XlxVHYEB     400     1a0D[o|?{vZԳo����؂��<4̇ܲѕ�;.��;�I��m��z�f��dh���)�Tq�|48Ӈ�
���H?�,FՊ�k���r"�,����IA�ON8%B�(�Z�{���X�3e�oyS6M�Fc�ܖMB@F�EY
�T�$�#���X�)�Ɩ�0.��q�Ѕ��p�7���7A/�͵fj�G���&v�����(�r@G�@2��c�+7��A@�nA��+9_�W��yeA��u����)k:�:�u��X�#6�0����K�.RN@�\�_�� ����	 �xo䊜�4
,wo�a ,%	�]��	.���Ƿp;Z ������ڔh}��u���n4�\�*X����|(Us�]*z2"a��6���#��RҖeܞ:����(�nXlxVHYEB     400     1a03��R�2?��6*����P`�`��N��)�;g��@���`̜{��B���� �{��o�i��P82���5����/�|<���J��Qm���~��~Qo��òRD����`LΕ�o��������8[�֔�c�۷���J.���}�[����T�oM�2�lq�}mc�����v&�''��8�(~mZ˗���$��������,�CX�(�8)�����Q���x�6��(c���2��*���>o(y�}�n��,���x�p�~�É�yh�T5��R��]`��d���qws�H���:�+!�:�����3�4���<�
�e�Q[����E���'fK��s�E�z\k���`�
3����T�	˒���J��#&���9�@�e���u/���}��NR6-��'�nXlxVHYEB     400     1b0)0�r����Y���-7��0"�.��<	��/==:<�	} o�X���f*f�������n5	�礷ڢ�V���g�gbA�q���0o8V����S۫�Ȣ�©M�9茭�A�R�AemN�:� ��@���i�Ό��ҵ���z��M8ů�T�Xm�=`vH�:�E���X�Oo{R�z%3�|�%&73����tp��N��x��*�O�gjoYӵK<�����"/%W=1�����V���Z;��2\��usxЧ�\��/�g��R�c��H����W�&��{� f_�>�{�ϸ����;���z��j]\8���8�B1�D����㐙��FݸnC0c.�=�u�T0��6LR j*�eD���RM�C��f�b��ل���G�۫���N�(J���צ<����w0sH�0���/<K�|>�XlxVHYEB     400     1e0����w-���xk�8�8���*�
·eJ1���7]�-�:@�Ǉ����(\���3G�i�����@`����2��k�6�!�}�����[��q�891��U����[��x%��	W���<��Q�TOI}��dW�g������βd�d�{F��f���.���o׺,��<��,�1+�4�}��T���׋:O������ƪ2�޻��fq_<s��Q,Uw��\��v�{���[���IB[9�	�$Q&c]�/37as̐C���n������Y�]0�	�׆��n��8�����R�H,&���Ʊ��/P���z��Ė�O�%��[[�MR�0�!�����F#���{��ހ�,����<VZ����s����\@{��2]f���: ��ȅj���%��@��*�B߃��Y�{s?��A%�C��	�P��܌���㯡�^�m9����`�ۖ�XlxVHYEB     400     170��V�8	���X��0ZNR���;/;+{���O0$}�{�����c��u�zu�ɻ�K����ˏ��-�*T��}�\O��jR��K��+� ,���M�A�
��I>��!=�Dy,�I;D5Ƒ����5�$�*� D�#�H�{s�y0�邟�O.�LÆ)ɔ,������z� ;�.k6W�- .{�du�c�ڰg5�jM��#�a��]�����'."���4!�"�u�yٛ\��е�E�J��ٷ�
k���_	R)`�������ȧ�[�^[9Na���4�����҉������aG��1|E�}ĕ0�|p�f�����Ĭb)��K���(P�5���ќ� B ؖ��aXlxVHYEB     400     1401��3ea~ae"��?f�/��`�s�"���+ ]��?�SF 8Ɵw 6�m�����(��2F�!n48k=���<_6]��	�X	����=3�d�a�R9F�V�k[�g�u#0�X>O6Hzٕ�9W0K��u���V��7��\�:LckMyk�z��o���#	v�f�t��E��BZ�dc`b���9ă����X���kX�g����u�@�S.&_�%�:���s�r�u:9��^H̦�=���wŘbc/77�9 ԋ~PU��Bc�̮�9-p1��M��y�/��"��j�zr�+<}O�XlxVHYEB     400     140P
��ZS���j�o<�阒䦩����Z�8_�N@[�A�3������0H+3H<�������tP ��S}�ԓ�pm1I`#��U�a�	�$<�w�zj
z���᭠X��s@Cxi�KA}¹EC�=�#��5�ż�-�X���c(ȝ�+'�Ҩ��40� �g������"F��<��G��R<���z�W${��*�}���{�0|�������OfɀT]��˧�0�n��kQ {�GmBt���!���i��P6(0���o�

�fN{a{9�pT���2f��ㅀ�����c"S4�]FXlxVHYEB     400     180�X�)`��ko��h�|�*���4;�ԢA7z�F�0�.�.�����Y�$���濃�t7SO����cɩ�@'c�7_�^i� ���63>�SŬ�C���Cw0FQj�܏����u�)��3�j$�(zd�M���v�^~^V`JCB�n��/�^hW�����z��H��cV����P:���lԴ����0G5]Q������l�:��8)�tuO'��U�X����*�5H�������唺N^θZ/&i� �G�e7-��Rby��3����e䴺�������^ �&:�'ʖ*Ԉkq��v���}f��D&��u�-�Y�ʑ�!6!c����g�Ts�R��x�>&��n�,Z��\�����x&��]��XlxVHYEB     400     180R1݂S�2�!�n@�=�St�z���;M��%�����mq�g���-����/��Ŭ����P��]���i�	������hȣ�@!���e;�>Ӑ���8L��oJ�R��c�el_����S1y����A�.T��j�ei��`H��q�Wƴ��,G��2��cR��')�>�78G�XECL�7����M[ö?qbt�"nd:��)ӗ� H��d�}Ǜ?�5��X�ݞEg_e�3����oR���91:O#B�����Lhř���|GHBk�Q)[#q_������E��p�r�Z��-���)X�阊{t"IT9��L�T��y�2�A%�<ϙ��-�>�kt��	E��bLe4��k�7�3�J[=��EK����F�JTL���QXlxVHYEB     400     180#/�tK���UQ���h ��n��>���B6�D�F�Y�o��ˇ��Xe�f5]�߫/��K#kb{e�GS�l�U
>Y���Q�PVr+_�")0n}K��A�:�W$`� �f4��m4�-D[�6I7����U�m����D�5&�A��T�AM]�'sR:���!С�4֡a�����C�Ź�y:5}:��j��։�F�Ƈ0ewf3���"d���`�"Љ6@�,9��7!���<��_!�h!�t����q�:E��}�n.�����'[p��VS�G����tx��t�`�7��,M�ݝ�h�͛�W�}��юR�2X�8����"�\�|��SW�xcX��-��֫H��4�v�9q"[R��S��{��
XlxVHYEB     400     1a0jd�O�Y]��."V�c���� +ȕ{X����=������r�-��o��ztyyx��LL/�ߑ�[�BZ�>��J��={\�O����D�-$���`a�ʡ��UE����~����z��vVk}��_�'�5�#{�e�ܩm��p������K?Yi��X�i�29�_��b4&�X�}�CB8�YQ�+��F?�TR�8�UI�.�(�3������Hz��T�6���4��<���	s�u���0�w@&��3�߄o	PfVP$z��ձ�
�i��� <vm�֤�����V{�\�ӗ��1��_��n�4���/v4<�-:?��7?K�*�i�W%#�Vm���t�JS���s�~�b����kt����������I�S[j�7U�(,�XlxVHYEB     400     1a0��<�,2h��)��'X�˕����)c�Dp���P2ۃ����& ��*��]�H�k�}��|�4V�w���n5�G�T��AM����b�Cb�N����+!!�>��"w�:½1����i�������n�on��&W��<�n�k��`Z��"���jn��W�iw%6��
����Uq:������ƸN:D���-���?�(��G1��Bů���3�B�s�g��G;]:�u#C�c�E���K/�N�s��������r_�^�@oGXЉ!Y�}ܻl#<��dќ��FϱF��%bp2ʝy�嬦!�F��l$Κ$-�W�cw|3��F�Q��Lz
+�����w�:b߭��FUr����.�\��H>�o�0f�k�=�e4"��~FY K��:�*�XlxVHYEB     22d     110�;�1��������}[`��f��}S����uָ5�����`�{�A�p�OZZ��~�9kWN {���O5ߪ�sC��3��^Q��!Z̿3����D�F�t����s⯧͎�TD����Ԗu�`���;&�-rm�`���2!mJ����C���TB���(����GwaCX��l��� �����0�b���%�׆c��kTk:Y�*�ώ��+�i�Ȧ��dP���h����m@Oғ�G'0׷<\w����?j8���׿|ЈK�