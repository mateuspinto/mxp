��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���챲-Ȱ?Z�_���N�^�J��6�Wgǅu�9�Ճ.y���Y�]ʟ^p�bc�̎)!�y���N]RM@��P���0�����w��Ђ��َQt�NU���Ӫ�K��vQOY�
�рR�̛4tӄv╽o���U`��o�mz�H��6��iOl�G8�y���U,G�f��𜦳�i|��S��}��D�aX�]e�ך��g�d��v�q��x�����1�i�� t^M%�]�ہ �j#��c�.�x1�2rt%�#]O񶢦�����=*t�05�G��d�����׉��%[�AZ�g�u
q�ge�b:�B@n"�,3��U�y#��͘bր��CQ���A1��ƘS�~�Ç����PC܄�4���&�vN�dWNy��UTMS�f�����Ȃ�����i�s�Ƒ��<K�L�̖���Lf>u��$�����p|S��·<N*QE��kT����h��7	��f@rJ`�6��G�]�<g+Q*f���6g7A����:��۫���+�n0B�}z�=�0��aą�� =0�o�	�VH�B�#��u�?��]��9�����9���4��M����%���2��:�~�A�X���nT�Lt��͍�dF�`�T��$��N��PoG%O�;��O
��qd|��}�Q
D񤌄3��Wf�ߊl���ɯ��C�K��\"�V�t7�:>��=��������!�	������꼏�;yw�"?��I@�kN��"UD3IN69�����*ع��vbr�8e��\���P�eIh��Y���}z��Ҿ�`��E�Pi��d�@b���8z�yFK7}Y ]=����-�W��.�Ry�p���|G��@��d�_쌎�C%'fTN�|ɢ���&
���6ۮ�iw��(�������N�'�%�;+w:�m��Pb�8�����đ�}����\ ���.��/��F�K����#�/v"���t��}3M�.U�OBk�2�����g���|�w\�޹]�V^�]��I3�Vg���|�E�@��s��JYG�vJB��IݺK��ܝJ�`�P�e>ܤ�?�
O��Q͝o����Ch(H�6��n��G$�J;)�98�r�fڊ��/#rR �M�8���Xp�5B5,(1�����UI����h!5�|񨩱!��NtfE�	a���%�?�VS�W�Iѷh>?v*�&o�lW����Rp.�=�������m��Xm���� �(�_����ΨD&Ҩ��r��i���6 L&��\��՚���e6���'�L�t�(�l��?����4$�#z��ݪ��E�B鰗��X��`�p��	Hq��7W�)���������k�6���v}:��^���>�?�|�:��z�*g��(Ji�+r��¦�~o�Dfa��k4�ʇ�ݭ�F��@xUV;�CT�l�1������ �Z�ڴ�4׻��c��OJu��
�G"IA�SB����WH�J�G�=/{�x�:
�f���>���BYh�u��jW檊�:k|cʥ���+R��Ҷ��ˏJ�˰�;lZAV�cK�����E=��w�l`X�����,�,�L���=|��kx���a�gTβ0m'o��'LF*�#cy�����i�B;
E*��Zx\
q�\�I�6p�r�`��ș�V��� Ռ딍f��+B͟��������e�-�~A��EGL5KF���Q|�Cd�{*-J��-�SaԺ���${��P�Ǖ[����p���a0�����҃;����;"���9ݣ+�����tZ�ox2v������&)�j���N鎸�[S��0ϼts_�_�L?�7�;�t��~A\Ip�{?����h���8,8������+��[��m�r�WË�؄�rR�9��S�C�x;��@7�h>����xU	�Eh�ˬ���t��|�����d!ظ+�PEJ%+�I��Y³�*�Q�]�h��<���� �AUE6qkp.2B�[���v�F��p8��&���t,k�j�\��̊��{Q������Q=h�E͔���d�A�j�Ζ?�"n�r1��9$� !a3a�E�z��`�F�8F��	G���|0gi�`ִW�:7�! ��/���TA�4+?������4q��$,�NkVn^�9�,�p?-�#�b�n�#� (��O�"2e$����&^ࠓ���0�y���cI�Dq�����ׄ�m�Yĕ����a�ᛙ�`T�wh��~��|�?&�^����=zp;��R�n$���Rs٘kOD	�l��p[�s^pP���8���j�P@f^`��_r�27b�@�Vn�p��Db�.�9�E+MM�v�N��/0&(�r��D�H����M�8�<��}eB�p�'O[���ua��cm�����dl�G.�Vd�9��(��J��O��n��ei���W`����c"�v�%\���]��IW�E� ��E�T����&@R#�u�w��IX��$g8U����0ǰ��#
I��v�Uu�4Ǟ.v��nF|��HG�����t�3S�|�b�1|5�c�U�w{9�V(�į�m���A��N�F��y���Pu�%S"��g�h �1��9�b�8"{�y��q�kȧ���zXA��.X�t��S`y�~睍���]G����,;�o� yw�q-|��4e����	�s�����d!	{�����趸P�����e�ؑ@}s��tZ	�Y�}�8z��(���` �$��R��b^F��p%3P������zc�)S	��sd�q��p�����ǵ:�GX�[m�X\������_)J��a�1UΛ�8��K\$ۻ��;-^������w�7Ԯr�N���7 �N�T�n�wv��$#��/���pO���a���������{H���ۦӎ��"/�	��Dm.;��5�GSSMQ�~���K3&<������[1�����˲�@T�%t�fS	ˮ�,"d�;�.����E3@1H��E����$f���WݔЊ��v¶da/vc�زP� ��/+��8�-?��r�k���:TX�$�J������b	p���]�}�^/u���H��s�6&Bs�A3c�c�l��в�E{"U��Cs�4�\�56wF�a m��Z^���p�v�P�����y���D���=�f�Xv��Q��&�����"�c��F������(Ve�. wL7������G����y_yؤ���B�R�gZ51��HD+�Z�]䠦���aL��m=��0uS%g�*�s�-'XȔ��cL�OR�o�K��E���g�mB0�7X��^C�\�J�?�L����cŎY	�㓇�c�a�{*��e�V���Ƴf��${ĝx�Wm�x���c���n<�Wןv,?���-ҩ�G���:�%�nH|.ف�7���W>D1RVL�,<���
W�ӵ����]&�8;�ΐ����0S)�Ԫ��>�Ȃ����1�8u=6��u�DO��t�_�"Epj;�� z@_̘��<r�^��[��uY���kE��nW��q�͹,j��.����3�|(��d"~;?VĔ���X�<K�!�=�hc�i	 ͽ_�_��&A�2��zH�J崱�?Ŵ����t;�w�l�2Fs�Q� C���L[U0&ሾ0��gl
.�f��}�n.��V'[]9ևz��OBw�|f�z?���ɊS@���cDԪ���>����u-k�HP+9~aE����c���¶Z =���/b؀�[����-d�1���l9l�$<��_�eJ1f�j�$O�&�-����a�4695T�������4R ��0�C����=��PZ��5�O��J��'�EkM/Q$c�\'����� J\��7��'��Gݼ�,�X�iB��1[����Sb	��љ܇��ޟ@y�	^�!N�qu�xߊB刾��%/�]?�� �D!QG7
��9�
??��i/��O[n=v�;k�B��I�����W>�M������ӑ�12x���;]O5��q�??��bk@H|X��q�r����`��K62��g����H��Nx�|h�BO�E��E���.��9�]f1�b3�hܴ�%�Z�*,�ʍ��"���@Yp&v��m�$u��u#`�l@n2%Mi2*����c|&����_4$�V�t��E�P�R�p���Wv����up;}�ͮ��<�=�
r:�ppbAR�ε}B�F���,['W~���ڙ�%Hͷ'99�_S?E�+Z�~��L�-��/�h�n+�1G��C��4��$�]�?�:`|j�<�VHV�m��J�"�v�.��>m"�b4��$%V��/>Q1�#&�\�@"G�%A�'?��j����0�'}�V�&Qn+*��ړ�%z�1��f�ݯ�jU**������W��C��l��S[�b����F�'G�;HϚ&v�^��vҢ���Ji"̲�����~xT�x/�"�t�[8���	�����x�e�y�K���xG�R=ԅ�[2t
�GѯETB|�����U��n/�]�
Mt�̇��I��h(��ie�G�NI��������zcy�
�ښ�^l�=F����K;���]L��Ю$��0��0£�T^�2f)��^�*��f�G����p�3h�9wN/x����ai����x�1j���|����'��|��Z�r��-�$P������X�s�'�\N�?�Q�T�����i��;�3�_?jK+x�o ��9��i�۴���@V8���ưA�Tu���Qj|a|�V���P�N-+�ڗI�f���R��X��d,����5^���h�V*�-�L�W�a	��z� �` ��O1p�E�l�5�W+��(U+v��U��* ��qr�,}Ң0[)�^":���C�oŲo�~_��$1֍- �WM��&?��)M�w�J���po�)���] ƴ��q��$��B�8&�Z$I/|�����2��'���]��A)9�m"=vDtژ��Me�����D�Ӊ�M50	96Vj��ZYl��R�,nAЇ�^����]j��?�� h�;�d��Ê-Ķ�ĪMwQq`f�T�`_�M��C�n�x��mU��� p�?/��%	9jO��Y�!�ز���؆�@|H?	>��1@.تf�#���<���M�a<0Y�	���
���qb���><e�]0��GJ<.�����>�2�g�ż<9��N�	Y��I`�`MC~�u��B9�2�s�'d��W/T���l��������R�M�*���C�n��yz�Er��>��,taR���GxWdZr!G��H���H\��+�VI�hX�:�|@�U��{?M�`��_�7	���)p���B��=����X����|�k1�X�#T�U����X0�Q5��H�'�$f�n�X�<�!�)T�9F�n�k�r�_��!�(%3���"ܚ?���'3HISD,"�u����vY<5ˏ^�3�Q^X-����h(�׃�j4�zq�=�����"_S��Y�eZ�;��6�6����n�_
���ԐSS蔆?>!ݱ�Ѫ�3�r�|�EV(-��̳U����pЬ�np}���c	��"y�c½�~���%hD�0���Dn�(�,�32b�I�ȶ ��&�D�x�א�����-�
/�?Nv8`@�ll�����,}���,� ���u�I�_G�ql(UW���u`��u>\�s��g���EՄ���(�
�9�E:XJiw���in�2LCo��N�q�h�.`%:["k��>Don�?��7�H|ۨz+������S����h���2�r���NJ��-���e
3��q�ʒ�\�|z���Ԭ?���=9�;`��C(T]A��㙠�Uw�������r��rpcߘ}�8I"f��y��4��ň>aP=�q�n�`h��dՀD��߂����w�O��y\��MD�a�X�Z�R�%=�T����]��߰\��9��6r[�m�-���CF������?��|c�q�χ6 �W���v�w�r˾�Mư��́�9"����cH%�f<%�2� �IM��p��t�ڝ�*����|�z37D �&_ժ�f�ZaB�3hg)�ΝA��;�>�E�=+e�8���Y��6�踯�Z8�z�B��r�!K�*p^���Q2�4���hD#o��\��oNXy�Y7٪������P4���:K���]y��%[��Z��Mq9�RZ�n����?^,��3	7��@<&��X�& ;Į�aaUw��j ��CPc3�|w~>J���oP�â����K�'q �nN�)�*ҋ���t�,��z�8$�Y�NV�]l�-�/p$�ܡK�NWl�c��;��7챂��.�}ċ�Z��D�b�i�5S��7��S
��Lyb����%x�]�tAW"@��*T&b�go>�qBi�����w���c[m��(�zw)��xޖ3b||{���Ì�:��*���w�����?�2݇����~����9�p�j���'$�7�
� �L���SG�^8��Iݒ �w˹
�P���0k�-DV�|]��͙.Q����:�Khc"�y@%��
i��	��Qs�"�:
���0B��|�2���uv*�xYۚ9��������N�M��2�Aa�/nS���x��@%6��N� �K?s���v����ŉ<Ɯ�NM팻��e�k�Ǔ(/H����	w��I��8!2�GE����$����*�V>�}(���:��9��4H�\%.)�S�׉u��rz�P�f�c������d�~�㮟<+b˜�By��������
�'��=���W*�C|�s��6�&�[�w�?r��&���*��5*��,ֽ,z�D�;}h����kǾgWZ��tV���M��m�q��|���1m�B��n�Soՙ�B��{es�����	g�d��E 0���7h�]�y�5�(0� �J��M��y\#t�i�Q�����uً���<��zH���&�����*?A��v�q�Z�)I���P�"���:(�t�=-8�K��Y��L ��0F&5������4"8�XU��՝��
�R��ט.	�ޤ�D�Ӷd�5�Y̕n/��X=Ӄ�h$(w��s�W�@�tpy J���ޮʰ��ҹ�g[c�oUT����_�:�������y���:�E���0h\�mXmo�x�����L�.�y�j��F�@ �WԠ�%�Jw���-Ψ�1�ܿ��F匚�϶�;��q-�ЗJ�*�}�⽜^���8���w�3[(h�\������ϊ��>%��!�5w%1>A�������U|�6��"9��ӻ�Ѱֶ�VA�m������)SD'�����C;����Y0<����QW��#*x�P���9KI�jhH@��ѦQ���O��u��[��H�s>#1n�0�������M�`G\��iՀ(��Z����Q�+���V�6��Vԗ�t['拾��Se�:��8���&Q�8�����W?���0ʿlv>p|Ɵm>���H9B]E��mH��ڂ�O8�ʶ>I�Z��ڿj��w�	\`���#q���q��\��w�&���^�n�g�����Cj$��Kx�:-��D���|�	�������s#��گ�p_�b��Ζ���_��N��b� 0����)+�Blg�q�S�k=��'��#	֥������	��_�I�P�4�׹��xtX�~͑�X�`�9Yj�����1 cx��YT�Z�`k�,4 r9��b՚����r�SPW\����?�9ų��K��C-��M�NG�R��YW{��jQ�P�=q�8����k��^J�xk�R1�w,��2�W���Bz�Ü8��w�h�6Sk�ސ!f��f��Zp�܎�c�g��i���uJ7�oY	:AW��Mo61�q?��b3��N�\n��bˇYu⾠�_j��b0a��w���w�ut��Uz'`���}�f\�g)�%�m>�wz��,L������{s�����y�U$�?� X�F��'�G\��FZa�/���f;rf�z��iJNX4<ζ �^|��İ��#�G0�ܟu��UJ��
�6iR3���bӉF��M{�����u`m�N��5��I.!)�w�;�}�]���<-I�iS�	@��4hh�e�iԾL�W��l^|���h��5���h4��b� ���O�gc(w�u4�ï�u����B���AJ(vH�;������"��5o!��V�݌��ń�6!1���?!�琣�� �X�}C�wKCʉ�/ݾM�;Aq9�6TD���h!20�]��x�7��-�K��5
�=Bo��D�s��3e�� b���X=���R;�P2Po+0%;!�� H#j���sI�腕Yf��90!����O�,��z���d�s������t�,�8�|aD�0�U��r���	՟�=�X$P���"z���V'D[���[߆���I�{�&K�}~2��}w�>��ӽ�S����
�h�bO��p�]�xB��E���� �V%:��pJ�o� !��*mv�8�{�"a����FpZ�g�E�;-�`��ZLV�eq���o	��k�pl��P���q�%����o�8hD=$!�!��KTfj�����<u�;-�x>�_���
R:�E	Y�҅R�/T��d=�6�:Z��?�᧰ uޣ="A��i�9b,���ZI�sM�����=�*ev@�m\�� k����"�N��7� j��qs�ppzl>�'-Ja�ZZ�H��=������2�=*�Q&>�Kz�+����cHd%���>����4�t�X�A�M���kuw�y��u���~͍�v����V͘���.��nÌ�,��4��Z�{�h�9>fZ���a�=OrW��ᤲ䚃�A�3��St�-p���z�)<b�fX���6�_��)fd3W�O���c���%�k<?��X���t�A>K� N�Em8B�g}Q֏T��5"�c �2\~����!NjF�g�L�ߏՀ�J�Dو '�e]G^��J��;�8X��ߍ���U6�1�
6u��g+���h}��Qԙ!Cp�W���������%R��yP#弎��T��ys�q+�V�z�8hd�^zS���=I��wJ�O*R�L�/���G+�y����I|�M�<7}��t;���# X�?6��.���a��o�U3mL�TR'�:m+���
���^�NE���}O+���C�f��l���HPK�y�P�uS��-)�>"ֻ>��b:��?�C����H���p������ԅ,?#�q�~��c�A�O��^ao^n�}%����!g���K��=/#�Ƕ�2_7E�;7Qxt���@+O�	�#��	��Ԗ,��=�