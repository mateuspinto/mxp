`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3168)
`protect data_block
X6Sm4cPUSBAnElBLtlFVHFuUd8gxcTqJn3/lMQY9Xk00WZUPraeGXgtKFfyIQOcxoeYR4Ngr2g4Q
3YxNEMryJdVAim5OkcI9XE9pv9z6ZdToDqQke0EAKhsPVlmfR4unvWzzL6I9erUpvEP9/qExL5Mz
iFyrZBhj9AyZ86x6t9dje2LzqkwrKAqrOwihcOHoZETTYufFga7axY1ym/qKdNMFeYwsLWeOSN4f
WANr65SxKXVkx5Sfe4dJM+hVQDvlekeYP2BHCMJvS2jaZLhqhox+YOMZtYoc/aW3eC3OgAYcfvrM
+7EaTtk2o6AMpyWTFEA7t1RNmblQtHBNKV85hluy5/sv1qpjS9y1HlhN8eIH4WYhV5DjpLr6X42A
CGbFS2NrkRLftyZeO05UTOJNuJFimPSweL2y8g/SvSMW1dExFNSaiErNoqv6JltdBDR9479weqq2
YogFEOe32O5iZ3ADDNNsmrodOCw3wo8FjwbkGSaA2IOhzWudZBu2+b72TGU0ydGHXZqU0TyG6jg4
b2Ycwc5DNQreSa+XlrGcafW6L6/BKoFZVEjSXJR1PqMBysDR1+XpCD64sM6k+2evBWD5jgXNQIoq
ZcASBkPP09GZ5Oe6DUKm3HFugL7gwPDJEnzn5bLECDiplgCDtPV+7hfcOtNocFELaAAhBjza5kpo
77iZTqSBbFDpN++Hx/jOb6ws15FWI+tbbQqFyDTul0mCjziVql7D2RSHN5J7jeyz7Flm4EV3meNn
dJbGcmJE47dAaExUYp39f3XH+4n2E8yzlY9JbKqXRX5rsc3f2UYeaJVyboOQ1UJn5q8tfUEkqt3d
9UccmDHoow0ozEgJHAliDSbpGGNZMTmsrgBeOpk8WqyAqFkTBmBUln0ubq8LxUSHbOucuybKyy9Q
L2JTYBUSqxzJSYhoqaHjrpdzSz17Q1jF/s3xKNi2XxaDHTfcZzPY8VrKbdRilZBT9gFTEeyXiyhh
qoYS/PArsbqiJBbHtYB/DfUEN3G4UOv1VhWgrXg3lvG51JOU9M07ncViUo/OCq/A86OWGT1kp5Ja
74I8J/FZ8QwKUIVU53C397eHW74ZZhWMsIFmOAttM+XL+s39/7JP/VGjQxZOUnABBgIQnRNmVaUL
mubrdfWWGhztTQ7rA+HoGQTBIshf8Nr7rbPk5LN7DMkLIOAjF8VgGjy9iGkjr2UWSjqvsr7wgRXm
Wvt92y6grjPNTaZUBVHoxXRt/oacu4E1hD2fhnAZU4uyZdOAk8N25us8HM6ardIx6iKIe+HmRYu5
4JF+FZF9yVG33WPzH+z/b8zHJlSIpLmNK1rQ3WpUaQW2ZagcCxM6qdrCWOvQAUf6um+2mPKleBb3
+QGpEWhbP1lDiS+IHpDbZIVr0NpPcCSNlN2kgEXJkjZ5Y26ZwDig+eMZtVIMgupnHIyYNc6LNrnX
O+aty56+D8EyMkVBmfqce7rV8U1MjefGYE+dpV13ObFQGv7AWBVtUQEoxCM68GyLZow6h+XbtmJD
8oIkV6XQ4MRyS2zzD/mxqiLvZ+lmS4ErcSO5atCg1eIVjjH8a9UH/VZkocuTMAPzj4fObY6oOMND
NhCe5hTT93kixre0f/0fhBSBZYVeEU1tcMb3A1RVnFz0eJqIZwhNhplt2No4yrHrdRqVSBTzSRMc
ogg1CTp+F02ojLcPWqjZhWZ8EHRBo9792REb3vdtYBRfE9w8DdBfuv2yHFwZ/9A2fFCO5XPAWMiE
0KGJvYC02azWDJBwb6dkmxKYJr/AG+DyY0cieaRGReSZ/eXWhdgRo/Fni1FebaDaTREEZC1FLfYQ
y5H4W3uqOpmF5+1psEzl6POkKtqMfpbJf7zXaXrL2P38oFUgP9e5t2XmmjUm9x0It8pMQb6wOb5l
1iIQKg4I6PxBCbg4EljMEk3NUHg6L+O6Yy3LYsVpJRqpDryBCTIdbw6R0KMkrn3K/2bWvKDYCIHX
19i61rQJLP6FxZAJObKMlgjyhzlGLO7uJMmFUfEBkTFDPTpnPurgpukpliHB1D1SpZX1gP8JWIGj
86oofozSjTIN7es7CF1v6KhuF6dDN35i0GTfwS4e5ZMGBNGI4yH8VngNJdLJFugQAAsjoLEqQdkw
jHD042iHmBFJxc+KBL3YFMpVUDnsFvt/1VrZlqxxYNWgdszjiLAeRo74GeQSOVgyYL6yszN3Z3wc
9oUUZXUAg2YIu73YQvMdIra3RML851AvnLqo3n7Ty/NBhKAtEoPe97ZS1CW/6G6zaUHx23e0dJop
Xbhf6G34pU58rupik3UUMA1LBIQ1j82l+8RFwzm6bhLyH27UufuIIuFSn20bbPad54Sjr5A22UUg
6msrcaXwFhLw9DytNKkfjUvCevsyIlkm65vVj2EDYU68xttTfGc+vI4F3ZFKCQqjPaIZczVN6y4+
t1TKueYh4zh+px3Tz0ACEo9KV3SHU1NSWPXL6F6/5O294PKNXENGon0B7UEoKNPr8A8SSGCOdeDU
N9IQg/dVVuvT5Psw4d3mXf7ek0LGvDW4YpWpBBy63Z6uxKGqjGp0tgVM3lWjVW3PeWUEbUzKyfO3
D5DhUW7amTt6B2Uo6veQvrGS2v3Yu99n+FUH4cwV9aQzYgJ0e7TzOnMVdJdK9+Vkg/BenYsMIxmC
DNsCV3j4zie1dJnkm/yFjp6rP5zGKLsqJ+QGKZND63QS/GBMtrFKy1AOaO2oiM2RhAzfc/o8mEdX
e7R6O+ULFANF+22UiQiQrE56/Lu7k7SQtNNB9Ev6sifRQFNBSE4uI5WXPlMhVHGyJzkym2IUzyCu
qov6sm00khgJ5yazlbwwyN9BbVI3oKMjz/Tv28v/uXFSszQxMrS+69Ect1ruzQOT6QXf+LbPCbis
CIejjeig9Nse/HPliYqPRtUo4udh8ybc3egVaVytEugeqr5Tx46zsKLEgTG+moK+aiJD6jn6l3TF
eqOZ4uzvyR+EbpHqFeA7FGrTPkTGJmwH3xjwYFmN+TuqauyyX5r6SfxleqQu1YqR7BwJpn6Fb/jC
FeUpizliV48+cAEYUuFNAgSk9cwlLMZ5AMP5UqN5A7IpnH95F+q2SfRK2OZRhp7p1wQrEem9opYB
b4np/IVR5yWHP2PmI/Iwv4GPPvwOgr3/zAaqJIkKQBl6Jyx+34Ez9z7hePHXlwkwjdDGNG5/TCF1
UnZyerkuKLs6zlYvmAVROE9JOhWvzfa+coQPTtKG4DINTcKeouk7aM9J6vQ72k3aPFUHTKsmlMDC
uRyC5s5T4EA9uxyYfL0G+rPMxwUlS3oE7ijl5sd3lJVKdeEZE/ZjcvM/RyTo93zw9U2aUVTACDPv
EOZe5bZLHlRCGcNNJ57Mn72/WbuAoCMZuo/bA/G7UrDI3GI4r1HXe4jgDzFPkbvLoZQFDv0IX0GA
Fv8o90YYb7nhdpOtDAJ1lxjBAhK81qgdaRJHbUAGnK2B+5GvFtcEfq+w3dagF3N8MDJ0GGEiYPj0
Azb0xGj044NVQLiOd7q0O40AJr+R5QplkqCiJFkMVo03GgMouganOKN+v0Jr7Fpe8sr2B585IjJ4
ybWZki+QtkYnlz+1Hi/ARSSOs+eHa/W8CvBymSxBRpmVf9GbMJl/jBxNl2hPlgD5KycBYPOApa9C
wT7nK0yypp6Bu7+rHA6oUECNa9ueJT/fHU3QHiLKALQRoiljFNRUL7b+lmGvXLWqLEis7vWAl41z
i+0l3rBm915Nm35xXVXWG0d/vaOwFTqWq1wjIrPfulKRevf2qsg5YUlQ84zwzcgDFg429YXRQBCg
/qQlfwzak8j0Jf6TTbv3CqHAciivNKaqcNnWrlc7ZOHEqvCpTaKANmH/IGT2UKYa+z46nt2dJ5a3
XDzqC6QpUmshKvmTsREL9AP+Z9NMjldqyjVu333B8dEFFpcI8CFF05edjbPKWAqkbbvq8DLoxtnu
q59BNHEB6/UkdnGdNNWEgIzqzRXgTOOGU8uZEJZumI6S2XQw2pMURAdgn7cGgv/YGxcKeGsbwHoh
nvNG1dhmtfCqLMQUmeFMa9HE+vWIPF5mATun/JywtR1e7TOm0nUEVeTerrBjtlW0f2cT1URNh9Me
N/Dd6UORUkCJCioMbhxG1Ng1jkCRvDlO8QLXhbJpj/lDkE9xFxB4zbNM8IwEwKGPMGMzM0hHChvI
haeiLKhvZCqdf17tXfBJ1BIjalGVB0c0DUCh43fPwdUi
`protect end_protected
