`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
GCaujQbBatqMLuyMBNAyT+DGwRF3XTeuvZVuJsaxb2ZISLu2+joreHr7W3EpFiCyiSfotVbaXa51
9bRPwxhvJEN+lQWxB3xJpfNzJMBdtdS/iodptO4mO71xHp5t/zXNeM6jKCrG1ypEE5rHqMl4PttD
8TMDDPZh/h0G27TibGjrMIcs912lbjaRuk3vHF2iyJtUxCgabR5KQZ3TW7lLTr4UO3Pl5xyANhY/
BcKc7N1pfW5A6KlD9ctVs2UpAFMAL3ExepVWH0T2xHjWgGUX2cxrK08fH2lV+6mwb266hgF5wMW9
tCc9N7/MczoA+F9HEiVosYNsYUBzAmdmGEpQmw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="jl0nqmOByzNveOgNcgy4+0/kMo6rOtauCvzoeaM1M8Y="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10000)
`protect data_block
F/OtDlWtN3RbSL3m6oqOvgAR4mU0xufeM1PO1ZUIPUOUg/5cXLvmT0FTegFxh/1E40UwamkfpWz8
yVSV9dJOiWS1j+Q64Q6EsEGjFxA6Xxg7FDCM2iWNy3R2kh+Pfnp2Dj1ejLyEQLVUYQLs+HtpYa7s
AqbD3OyFPnViNyskjE81Ksh3+c5N9kuT2S7+dXtEOzfkpCBSTpXk4ty3e+fVt9Rn8+yHO3nTLFJ5
rlireAGUqcyG6JVX9HL/ZZknMDeiiXSXHkKaZAaHjFAeoMQ7U3AgXDCJ46znpsXf36tPdyeesOjA
9AArFihmcXrEi5SXZz2dcCHeVX1djIuiLZTV/D5b0DpWUCnq/kfQeqW5QnVdJ162KjvfDMJ4Xvhr
5V7AmoblUt9GMf1uuYOTbaiu3GwDPKPB4L+4Sw+QgrZLkfKHolvefnjd0qM3MoSAeBle8aA3uQOt
5ePhyn+kHDe/pKVWDg1A7nDLiru2PH9JkjsTrsCoYn3+qGwbm2yGD1sZVRc7akvXKcC+YiF4M2+W
0CE2idz79btOiGxKn/IU9ZknGqwTqEgpA7fTq+Is1DXaONnREuITfs847ed0i/6XGWmrfQNwR+xN
8A4jt+a4alAj4tBUiVVMo5qjcmWh6iiJjvYkvfBz13Dcl9uZQe59OPHVgKbiSpkHXOvpr+8Xc/pj
Ld4OOAIkWOlE4UaHGO4a+7Xm/AptKmYZm1GNit40Q7H3aCD5NkwpmDnwqF1YVmF+rm4kwhciUGPs
6OTePdytKHhcJffv4hcw9XHdVKA2JTWgPZm74K9hi8z0Wn6yOH9rFu66mISCHdGpbBalUEAKkXXz
lwPPhi+HgQDC0UBkR2Da4jH1lopwRp9fmWFo29OsNAxwEsjTjyh9S4U7LMbAdtuoyxz6d4ww7SCI
ab8LO9zTCokSgV8N/kEdofuy4fafqOMC40xDP2KTot82jmrpm5TjUDzkNu5PWxfhaY59aWw/jS9g
N2y4x/LRO2UQsrYkbr2sNx2GOnyycAyMgotrZixeyTqCRPfTHtnioKwlGAJ2P5Yf8kCELtv+LH99
FW7NF2HPQPDDLr6gr59qe1faYl08skuknApPbPIrt/H04XMJka/+7dcw9E4Q1zf49cGBIsUTpRdV
Tc2gm3MhKTyelopP35c7qH6AM8/EnB2Bhht9rgJBFnwq/QUjQUlM6PGA0XToSVIpM7zx1TGJ8+Mu
tDjG9c3lj4DIOiLYHriCS0xPdvkEoqLJO/WHkSMGhP5E1BFuZJEWAus2Qb+guHasOZ8su0P0adU1
55ku1Udh0+rnL1QgXLiOGMmFp53puT3vWZ3TbHpxlk0+8jW4lyPJYF5/GbyXzvi45nuYA/q5Gf+d
6PBRfymP2ipkd/UaMrkLm01ioQ80ZJ75q0mpUZ+vkoH6gEyDOas8vY4jRyapf3Ekbm1t8xZfu8HE
amtMsOGUnJJ5GBdMPQ1FOfo6OsoFouZr6C1xw9JRr10Vh1Pc9uYXsjXm6Mgk6+hK+2zb89R49Rc/
XeaWOuby+QeNVvrJwiOF222pffwgrpvvwWX6U16UuW1vkpZFdJOCK2KqqdTRrgADc2WNCd6n803m
XRgmtbti1dmjb8UfsqRU7m6VJ2yMhzd65uqzVnfQuy7c6qhcNg9ZLoX8HX+WMU3s0Xl6rzdrKfhH
rz+McYGUXpYME8ukQHzKqEPfThEHNsoyUx/zvVddqmoXXoDFhyemxzYjnq162iNeJjxx2yR+gflT
j0bCME984CldfBSyADR/eaWqXy2HG0hrB6dumvma2G4esaUi67f9crWjQq9ZF/S3O/wEZ53k4X/+
/D6RxbgCYWmaGtCJyY7QbZx7ZI429ipFLx7peKQn6OwsDpWLTFGWKowYJxsUUgvyOE+k27phaxbu
66Waqy6swiEZZrFWJg14MrVgFzbGJEuN9wvySwY0pAUK+9h7fCeVoIGoeGqnztVAHj+Wfi0TwDSM
n6B14nwQa6chgXGsdIViEtJc+S/G57CcGkiTdL+Xu2WLwiI7GEq+cgIcsDlYzloFQed9FPNcuIP5
A4rP3v8qYL01H21fJSpwLOgQjwKlcQkpJgTJD9RQTcYdx3iIpU2K3LDsFbp72GMhTGjXovwLvd9D
VYzwSxBOag6pJznfGEx11WSjfr9QN2kdgVRuCiLl2GHn6ZdaO8oOPYXdR3Z+JDDRYzYE3pFgWVsN
XroPab24OGUT++TokQLO3cfl+au6Mizq9BlFneGN6Gd09PpHfEl/Ng/iwsQe6FSS/MbEAlkr7zDp
J561Z4aV+kWhZrsJODU1dgEhUygQLs77JzyUZtHfbo9L8fVd9ysYh5kBn65hf6ohqyolubnPL9+i
Sm+pCozmuD0T6QXh+MZqXwjksDAAF4G/2rhag9gTEWIyVlerxlx0uqp8a4nKK4bwf3iaUt8rD+i0
BrMwaG8IBCElsiSx36kSC/mFpjO5ShvYtqYr0O4VW0RFTxeJ62F90xwgRrwTxp4ZzjLQVGn8uXRV
P/01SA72xK6l8CdxHNi7/hfHlfKRw6FH/2ev/4+qV7G6BSvJHHJKnAvifmYMAPnRFnw6ShWrI2Nm
AlbdMuePqT03gXao11hW54k01uneHu/A1WYe5o0ExnHhad9gutYwALQYTKTr9C6qeCwnHrmXVaWf
PrNz4ZiTL7iwYIoZkqGut98Vj/w0ePDWf36SvlTraiF18ZT5ZdpaRtDUOeiAy8J7WajseA6ZZBGg
qnlazMbHE/NRBVPo/ZmGj8aAuA2WcVPcz4xXs1f+jrLHkpsFmE2JnwHED1k0YVJl1uPfs1QYcrTX
al6x1tqJxeVojtnC/Y2XEjOYJxg6/CFBjAgLDk4FIS/LeVOqQdxDSX/B1S4ChQA/tCSHIFUtuVQf
I97+OVc/ltYZlbuckoZa2qwe/0ngkQAGhmMMWjjoiv1lCuxxFEUsaOVRalIUiO3qurugJ3wrGnFz
ah41vuOp1qOJa+/4XpuNx96PoUqLDeQdA1UHk8Pg8XTZmfPem+5kujk6AS6eambGnoqz5MTYDcFg
bwQFfwonb3iIMc/iOz/JKmjEMaNEaRY6Qr6V0IKCZ6FWnG5yysZuaD8rNc/Lmo1peRxvA9m3qgf6
yvp+afeNHA8OMj4P6XkK9PtDJ+w1eWXTjS4kvTOwUmBnQ6yHDtY8/G+1rhVcXpE/tBoZlGNvfHuw
yNe6RQjRRfPh2KxKklrjnKOkVkKSze0zbesqpzpWAEivMJJxPiprnlW/1PpHBqgqYEms/3i+vIEq
gpPHEqxgX0/c+BKEA0afb4qMOTgqfWDTGxjmpdm1ShoA0CAbT7FfOc4xLTOI9qlxUJqFUaolOabn
c/23wNZREC3a1kARg6lfl3RvktoJKNp3nCPBNVgjxNTzf/NgUSsWcTGVb3hnrV2S6VBoXgtsDKLO
kaqgrt+Sp650KUfEDpwO2iIwVEQTHRoKjw4QsOm4ePDbURP/pa3ReoK2iBuMUxW/PG7jJPFWVQvm
FH2YnUa4lVb7eM00dGntLkrrhOnyi08IC2D1IYvA/deBeNs/LW6syf+wc1+YmkL9e2OqSLXW/Lo6
Ev7uxaXDVavbGDm3Je+4GzjyQFhtaUkbSGw5hMC2FkneymB6PnX/+3cHQeWxvdxk9AY3atO7jiKb
Dl37OWgWHXKR84NcVHF0YQbDR/OkiV6KsSI7Z5eEaLC2F9LSY61Yjsn0UPpWxmAjIfSbpok81vna
lYJlZj2v5asCGGxWcwvCZ4TA8mgYXsikri+5A+KAwwHRjNk7aUYhrPQ32pgboW4dHcAHCPoRygcE
JnaOkoQchRbqY4/9MGyWkvUqSQ/ufjNdbCtkg59h6+ZkoX4y7KkLQsLLHcs/vCAVPFr82kTcuDOf
MG9XD/dSSyXsYfAS/LSjpvZnxUyrSo7PBo+XdLFIhwfKWLngryO06Yw28j6AjEVhVqrdhxrj7s6p
aokOjDeX6kEIHcbuMn8J1veQ8IZh+4aEWEnoA9W6c3zGQvOa3acQc/tGFmrYpRKGwQGm+w1aZQks
i8lEHlKrx80mmZW6PC6rI/H2w7UKFqqVcTDN2xW2j3EdbN8bpaHf2BLmw7ikxjSaZB8GtOv1hOAn
QUC4ZE+gnp5rwfNDZyyqJPZN1rbwbhWV5cwfqzXikv84QPnEM6onp7WJElfdhwxTJ5n2a8Vt4OzI
7syZwYP9UTUdTm2bA/qtpBWZ+23M2PIPn0oV/ydZc00qTImKHMoc4EhVouhzJOaktjkvLVL/4ey7
a7KpuEgScQDNT4jsPw6nE7bReMyLH//mvZptpzSS4cQEUSe3uDdTQGi2k0ZbNe8Yz1+BSHL2JNzu
A2Oxl4menaaSQJwzLdSh6ifHJqI1XZZsiAlgSK6aLE9HANRQ1nkDoDF+4wWMUIi+d/Cgx+QSrxuI
dP1T/spOV3SHCLhbTbLl8VekDX1P1GLvsNm98UfauQiZ6U+11LLFo0ecB5/U38EQeNQwV80Cc/D5
67cYknpHNt12ndNNWzIC9XYBtmdBHnMydH8uTmZzflw4dljRj02thqIa0IBHQLCe2vi8F/v0PPt4
ahfOmao9ckzz5qJoWn9qol+jgMPGyxIjABLY6BbkBck0YMYbYB4WFcevLfikFR3QN0vtFG8UG+UM
Q4SeKJTbLBDrfEVuLdWTii68qwS/8hKIIFX4W7on65Pdh+RYmFeJYRsr4nTiJ8GzHppN8/b/Ysgy
I4rKpptzqO7iTQqNfuE1I/8CzG4p7RP3iXCieOCL/daml4T7A1rMgZfkbfL4GCs0QMIrfwoSoDqR
HLjd+jGWUxj2lIG2T613rol5xN2bZXtwN/z8GwhaGFSxTNhiGJBbmlMbIm8DX4iIuXLaQ/mjckRh
PrYbYTvttBCd/05l1cRzILWKXxfoVYiIxGVLb4nLf4+jkZvcKEGetzde80kQ7MDmutyTnsvP2m8W
zTRpee4eIJuhyTrsDKdebMa/eVbn7j3DzQqu+IefAiemIFFkjSnZjq1JB14/y6E5ns7MPiDrE07E
W0Kq6s02+62eo/gn8jBzs0i1tQfaBYUYGbA2oT0sBns3msbL/Rc8YJ23e5XRYvL1tJOghgYyw2fc
J0o777j9fQaVnrUflF7Orsn1WqLkBXfqx84dPfPGUdL8Gpdiuo2oaljDXfEHbw2LXRj7emqXNnIu
j/i9SFNDMef3Oab+WZwkyqMw4ZxnfKIi3YEOo0fK5DMCVn2A/cCD9/ARZ0LJfo9Dg+HmwV0/T1tK
CYJjlQCFR5LOKrYr6/uFiq5EoLmhzMcP5hgBqjs7dTOG28M6lznFSsdhFaJ1t/wSf3HBKFaXyjJO
dy1wKzwHp7PDu0OX1FDmBs0xLYKxp3zcQ9aivButJWu4WomBv8l1kfFSu4dk5BkReFO9GVjFNvUA
u3/vNYNKGy7GXtnA42j1UNE8koy7XiGv5JUgQV2Exq4obA6QgmkmnwUZqBoxm/h4U+C8jNMgaIWN
rgnHygNZPqA1nbfV97toIDok5uo0fBikXnYnKJpG/Fa/h8shS7TWBarcN1GIaMkQx1hqHgK+LLNd
nGHK58QQb8yZggKdiFUVi9QG6qtBjEjajuBDEg1pa+g/Aapb3SdvoEi3ltqUs6+XFOJ8iB/8H6AU
gsvtYrdgiDdYc/U2DeRK7jdirTvGi+xgCs5MTk7WRo89abs24fGGFaS+EtTN+ANuVAwE7CCKQWwp
4y84bk+4ZkFHBLA2LwqU9/Kh4ibklXcMI0bfi6GtmqzmFtU+XUdjXUQPS4tEMvTC+WgSOLxfkDBt
iZ9PhGhWG59Ly7t2WYUC2/aJw8qH+KDXePaH1V8gJ9qtUV3pFgjtDWmmbNHlF6WuzhZ3OFB9/eOj
hsZ+Au/vTmwz5ziV8KZci9nfLDkOAfJMXwM+iYw8ooYnzkPRD9RryCgVU8akTqPUpUqhPzG/2LUl
SbLCBnE+QS7NB1ubMBuZXaTjG/9h0DUH68IMXGOyoOohy5vIJwm20qZ3qipMxUO7Io0QERLDGi9H
/xA+LaqnERjxCkc5qbGNtMgeAQpNdARAKI8z+G4ko1J1bKlzghzo6qYXsdnqajuKVWMi2Xf7hZFe
3EPPtlSKlb+cmoLPswooVuOb7ziilQJxaZkZTD+OALGa8gqXf2h1IwE/t+kkn2hZeCNNXmClUkTy
oBoyBiM4zkAwLeqOWTB3O8SUgs5UlqniPx60nIQZ3BtM2vle9Z2hF9UJoUHx4DJSvtnpNynlIeCz
wDhSAQPuRYvqicst6oN80gf0fc6AiWf441Lkjfz21jtUNFG4v0+OpwFD5FvejyLRrze/3uXYviRI
nze/KdjM4S0AigTOLScnMGQWvXwCbIfd4ZcsSxsRMZQ0pnIPZKbo7tA/kmXSk0PNvkssXWvvqHZn
WTqppr5jh5yLqK+c7LXlI5GcuNlz+a2SmwBVGpWKCp0LOJsHShkt3xeDJ9cWLQNqu16yKu68GWdI
Z7qHzkiSqqzDFTkPQ/vqXyPLgFGH+ZvW8c6dyIDI8VtR3zzKHCC+ouVFrB73pmKv2IkQhtzzDt7b
PWjAVp1DoreiO8IkO7bWAOM5ymeblajZe+ZsH++9V7kRa+d482ThgcBDCB4SCTCaAgMgcWlY8dI4
XItdT+ZqqTGS6/+eDgVpoxVLmYU+/9Za1+FfCFHz3kz/FeTQVWKc+aosQs4jOohxv4H31qzGflIH
aIbIRPHwHHPQ+B987b6PbtUmRpVsRa2oZw+s3Yv9VEpCiffa5CZ5GivpJRyY2PtVyUqas5zAM6cR
7LuxT18cvV3hPQvKLvAk/S9D9uyyiRaVi1VXc7THUNefPzWwMUBTvj7FWG+Fj6h3aS4F2s5/kMqE
JNSMsVOAzhSoPwCnBVUj6t/CcJZ62GXVhZ3MuhXfL6l6oTmrmGHiEXcqEkfbx0nlMlIM2WvQZOiA
Ms05oqat3mmbTwE/kpkuLeGNTWfSs99YDbzpKNeGHjMAJQ8EKCFmeT5N0nrzd+wRM9UgtjeN/CZZ
VFfLGFYK75ZfJEu25K2djPmj/d+21sO9wwfT9RGN25qK/M8KE9j8yI5CP3UMl8bjDjaKyTo+9Rg5
SDwlkv339qkJ4GxWF1ChGJjzV9XTfVNYM4u1cRM0gPNxrxa2rV3TPYD9Pq9VBGx5nk1r/+Qtd4Vp
lHMj3uc0h3YWgSOU7lWzaskeUoXCiNNSTGCWMfPoDDMJWxIovsmLqXmRmeSCvkavowf6C/Ix2f1q
uleOKfAXBkOTib+AVsadx8s4OYwjKs41835+OGuVsFQs+h4Jy4dkbwkuQcWatvCYNpUH5Bz3lYcR
x5HyztLS354s1U7S4KmMdBhWWGPlmqCydMkheG0WWhIf2EGgmgAKkDmR4rOTpT1dP2u12uC9Rpky
s5qU5TVw8aAOGiX9qlGgl6OKlAgSyZNMbMPdtjZOZ84lhF1YfVw/3ioyq1P8dZ8tsptBBO7jh8co
qHbRt5gWudDab0uSqHxj35I9c+cFY00Y9rXtv6xN1O9GgLi4zEaUFW9p0N3wZvrCtRkJ8Md+rSaW
dl9LgflvRbCgAyGhL38WAkAnugaefcVNAUQ8LwfCGv8EraqlrkWXJyktSdQiajHkpoHeeAso8z6A
v/2QT+tHEJ6SQYwe5lt7XNidSfL9+QxYQPXKEctaAitCX/G89/eMvidg0etMd7967vvAtuuCRC3F
XxAicfjKZU9maUz2MLqqLzEfH19XsjaosL9Mk6hmWDLl8n/U3/fL4i2OayO7Z7KQHmOpCCKM6PO/
OqowX5ASaK1gKv8sZgH6MEhB4eG7H/Ex7srQq0VyFAHvTIkBgOCRuWZB4+37QA8M5v5KQgw9t05O
a8AcCjJJbwcZOUIIWUrR4S/5ASRZUhKXHlMlvZX1scEN/wL+pxMRxIOfDofD5vUmqay+VK2Oc2dn
XQX0LoBRWGflgPPuXQwwPhRw4vKzwM1TNoal5ibasrCMQQhDFy9v2mk3hDt+0/TthQHESr+AXgjT
UZ/mrc0E8pSLYNvOYxr9WHNzCmhfTQzyTTQexn/vA+Sdy44zgL+reGK0/GurwXuoVqDzwhVAUlS1
GN4TDbqhPFCLF9d41lCm3kObKkAAj2qWd45x+jtvl1otdPMeFPY8uJnaSO3TrYIXh4mzu+DgrXSc
ptSiM4M3QilgeXH98iwsSXB9dzEtbSex5kTlA55ndanSXRJqlmKoEaJYYhwcGVTjjl5skYISTg9F
1xlqXbF0WmAvDPOOsEQ/NECSe03U48IdtHhzTczvWB7VErFhJME7Z9Uv9LPzG9G8exxdtTueE3LH
Xg5RX3OnjnaySyuMPpCR0k2BvaEsKiaTCn2RUwkptMGZ1EiWERaJzZ7qbIzfMmdHt6o+tJd/iD3B
Zs9LlJyteooFZ2aMmMEwDRWvKKWRAoxt3MeEe2b+rwBRTJFMxzju6BAqnXuKmLZWS/7s4koJMori
E71TytMUSw2S8/iu4spMh+8hk57fCKvsbewJU1VXBq3gzR79Fq91PaC9DDTvjTLJUhhhFi75QEDo
bN7ryeQvMrZqKM+ocDaR+/WxiUgGmPW7URKj6OkqzPJdK0dL+G5VGMumSF3EtJc0HTHYdoJHiQb4
85S5icW8x3ySrj4MXMHx4Y5QcPLTwcsleCCbQJuSm9JtSxf6hp4rqA17jxP/Pw2J5w/qs0r9ZDsE
qjqOx+8wyAY4VCHzRgV6LU0BlnxPrHy+qRZbrih8Ded97bCvpDRF2MnewLbsqDBPrmIMHaqAHENl
PX49hHuMBg6JLR4CZ5Vt05AXyIyTwS84CyyjGkDNPBRDmM+MpiLCXfXfh6cXvZmt7br8LvXWIvpH
FVjf6n5PTMR9eTMHXQgx9leUIuR/rPJTewCvJfjcrJ9j4IZA4vZGj1Tnwk1leWW81mSqYb/i2vwN
EC+sZpgC3xJG9DcMoiG2b9469TD6V3/qdEA+eno4wJDfh8pFl8p9SzxyRnXE3IIf2WD3KT4yU2ff
iyaUREcwjykUe+wUwZh/jlGWJo19p9vSNBARxocXkYErw4k5yMBFuHe3arKxE6FbffOkJ46PGDqy
LrUSqBZzWvLMJ/5jeeVYILJi5NBW4kF5uLjsHdtRrzrFuwjwVTUXdejnU+EZTa6Jdciz4UTyApwz
FVIi690JHMyi8ifXM7t1Mu/lmbebxtxI3M3sTKuGtobYA6jMM2MyMKBTxxHz5SlBWh8+1W84MKCc
L7WGYPnfco7rNSlyewpNcYgy2YC4II488PdEXBeXHzfcA0Lp/Rkm+97S6ql6SWUaT8EmWVBBHthq
Lq+zHFcYrjq6RZqvQ0xSv6PUoOk164Zc71QJ4Hx7XrijFRuygkIm9SIB0Z0/+xlHFIE1etCg+8HJ
SS7Ra7cncSxdTBQql2b3Cup+OycvGxQP61+Gp4swIQtrN889MOKplMgRTQKAmNW7Np/bdpmVwO6K
gPvhqEEAUmnp75ZSlaRyVtDhRmRsX+0VPzTLtinxWM5vM9LDSJGzc/fDpavrehh2RwRxhZ26TAqA
HmFx6uYFfvXGvuNtFGO5Fx0QXZoRO5L78DAtOmhgkgC+5STKvE7ZSxdEiyTmD6MMeNXXrrFABoZe
5BuBeaZkkwNKs1UYtGiK8g+6pl1Eo+f2bHmoqu+l+sQJugvanCfBOyhUwC85ZXCg6hxndU8vYCMM
SQ4KLji/hopUxiilIpInxrzgEQdEBt//NbLFfK11moJr1ELiCjhBAdUd7yTWY67J1fgbCsPQIGD8
QOMCrrANRH7HP7RllGO5WsnY72i0mf06XFcFQMsQRtzKomc+cl+qTnYVixHNprU9IH6j3go13bCx
3Qlfps0ycec/WqptslOZQYmR2gWCr62FIJs4X9RZKEQApXCIhePYkNDXojJxeAdcxUUzSB4Hvjpw
SdRnpWGP0Cc8O7yAeeQDNp+1Whq3lajXMmFMjUmiZzXzmGXm7AGPH06Xl6n6T2TnHVEOn8OaR7BU
ENrWME2xoUVHPsEUI7a+WgC9rFuAeKYqun5klu1WujiX7wZd6norx6V8cLN/bQ+4V3582Oot02j4
Rh9VI/1aZC20pMbegYmnX3bOWzowxIPLd4ytm82YohXokUzOOMDBkEwZARlmY90oHaqNZcY4vQOx
UoGfkyJTsN+tReWCq9ls3Uo8imbzblJPBGH8ud2y2cWstrHvkEAhZjsmSSPXsuAwtdwD1KocyWYE
ySh8HwdRicu/2HzQkhqxKv5zTsyPlhFqNXBH9M/WxL9aVyrwX4Dqg1+NI+eoy5Bd357pqAxw2FDc
kFOcJxsauGBJzx+gIaHEtqh8I2H8dOrbaeK2IWX9oAGFrkWpKzhjvDVwn+sMinSHetQmnnTlTkRX
3eKLBvJ1e2+Vk141OUm01qhH2NDUSg+rD+RGVmwHBt162TT2WVED0rU7MzJvs2TdVOm26IvdUM5V
S06LZrBcEkinayhZX+MLYNHoQqoSyZv3YUDL0715G2nq/57wR50Ilak5EMOiewbEIm4pveRuc+fl
JmvX0FlpXVRQ1ZynwQjJojWUKPBn4l1hvJy4c+10UKBoAfFm8EbZNZKHUcKOyp9VEWnWfa9sMGib
CKoGdNgRw5yOyi9W3tCzWqZzfOiUT3nQXxauJxCTMYN4jAsPdbgUgCHVwvXWvfzKPQU7hI2T2bJP
6BUOYBpuArWTuIa7gQHXjSM7riv00jJZ14KJTfpMdNmiy0ujBUn2RxN+3q8IzNyxvUcLt/Qx/ePw
wKCNoF6skTxtcb3dEdgygVbVl6D5DYPvqkmmHOgaA4F0LAhZ/AIjllTgVJT0moN1p7g/6wqTFIPv
M2yzD98GBVtYUNgd8G2oRQLvGafZxTMMO9L1mnUTzkhmEXgVG+KuhbNzQOAemr/AqVe419JDvcN/
tiyn5tEtI4/WodVYeMzWZnvRrIKlGb3hMxB3DXhVLzxt5o+2M30+bmxgT1ZPZ50dtLpzcyDsinsG
uV0fkw1bSRE5VNMR7R74YdZHCOfPETN3CZcsk1vyyBRXLmrah30Yg0uz50euWclld/8Y/FJmO/re
wBYIBxmOJxvmrSTFn/AuZGevVXLVNSx5JLWNRbgdjbta2pMvaHUl9tILeQmgUAJ7Tr+w/7BOuihn
MM1Oxt4EVuQkCQuu+ZJJALtnhG/I4cLgVe5bNmXr86pHA8gfZPJf53whtOIQdqjAVV2D7EcurpLZ
IEM9XLqCa7CRI0Vsl+2JAt0KdZx/A6Gf/Ps05bZ6HofeBAs7UFwOE+Kmm3xuPTDF0qH8PZp5HEp4
riqxCt8P4mcrTsiB+0KDzD4jrBFEZW7fAbGv/uHGyspr7f+aRwfj5rQN41KXhzi7i1P+f+5AQhmh
cfKqgNdEhpBls1P+8kcWXvnLsJ/ovHZAzOEme3d1dkUT1YBWElkZwPfLXg22CTaiLu71YZo5LDNd
NgrrgPswa+2RQbWJSVcPVp9zlM8hsNJVovWbI1twBeqKl4PNubWHNE51mhBp4J/FDFDkjZ312ctQ
EShK5NSM3TTDbpWWaK4sAlP9tGiMAB9YQwj1BRiYqgYzW7EnL62ZVkPfc7mTIireYeD6CZqXcKvV
Lo2JpgOvT/ILOmnxBycywoUS3KIVm25c5oy7vZXDZdimGjQgRlySe+QUobMBbfoRGBQ8NAZwzDTu
qLFJbstwTmDvPtaVdssnwBU1awGyv6ZwpA6jzjsJiZuPez2z4qDQmeE55/iTy1cWXsCxaGKGH/ba
QcAof6h0jVSR2NO94tezyAdnp5ankKvP0AJKM1Se0Dk6rBOjW3a6jyHMpDbh1nFxK1j+uSi2ud5f
w/HXvYXbscFwtKh1277C/cUdJLtcZWrBblJp+34CbokUcWGdt9WQzqTWfIeV0Zy1gvfDUQqdxOxb
cstnYIiB+Cn2OjZNgQ0qIWioVbUseOM7nCRBowu7Ad0pQZP81iMuj7E8QOoifmiFsOJOFjgZ4t/7
nANcsQV3+OqkDoWOQoudIAmXFkZkl2k0kEbZ1wTRIixlCQjp8TTy4rXLqutH3pdgz3Esmcxvihgd
cWOhH4um2jRpVU/rt8fwtSn4RqmEd2iFgTTTxYztR6hmvGcI0iuuWmSfWY9fA5AoXv7VS0QC+kpO
W0EGVtCe3uKcshWGcq09/4W2OnHpXJkx+0uGXny+tG2nB6covM35uz+95WzG83+RoXoDeg32+xR2
j5zHbV3ngjbUc+FIDKIZas2aPfaMo0ovbmJYQxDQ1A0AojYK7ZprZKPcOi1Qwp7/dro2rElDrU9P
lmebhtfDYnI7mpTUW38iY6juZhXmjGh14ztsbQ/v7rP4sylD3XO16qi/2f3rDfCLnQBthvpFlKmV
cYDHy4ZycrUcrbq1nfYtdjO9K2uHbY5yL1jD02ebNsaMn0be4nj8OtS+8UTnxi31+Ib1CvcnUylb
3W5GwJMStHg8YEQxKwFR7WmBfHPeY7wPazjejlDbXngcut6DsrzzxyskUW3jhPjBjNhS3ud4H7mW
Xnh9A4/v0060U+bwQzs/pheyhHGPasFqDMhi8P9GIoOSb3rdedrvjRedMwXb3Yjy5dCgiUkQLVh5
L6WoPH2KW5kbbzApFvxLaQ7zk7UduRsQk8Dcgev/URU+577iUJN5SHqPI5xqhjZGccGcM8WpBTnJ
4htWSlyfCMcyld9Zh8tZaYLZYxxD1DkYcsWfZZZF/rSZ/FkVDt/BnRver3lkg4qqCc9n+tmEuF6o
HsomTsixkugyp5IVtzlVlzPnbyXpyUqPv19pnOObB2I5Xu9bXsqVa2jpSvQNLqJBXcCLvtHX7nqp
WnP2R7aolxLUbK4XuoLv3snBhQEphLcXbnRILSVMASoe3IC4GREsCs1CG/4IYQkU2cu53qDs2zRC
mLB4248y0Jv18puvccBq+yrsWJEGRsVwSILwDVUI1RGAWgQsRDvNMsb0Wf1b3jsx+9bZSy3Jqi8S
HLjkzOcMD29w8ty5kmOCIdPt6ytvhiufBKovxL8rYHS9bDUBgmnzTUBQLKj4mbyuVSV2QBMu123C
nT15QZ9kVVWCvAzqwupUztPQgO8t2SkV4w7zt2qFTD9O9dQxXoEpeN3nBS8+ArlD0X93Nis2OF8K
GAGgacVijxwn0YV9GjyvF6YPogBoYx5P8L2qIwrnaMjQj0l/e+8e+Np6EVK+jPEqk3O9GCQYjG9U
jQtUDwcZHxq7cKD/l45FukxjO/pk9C/EkVOAgI14fV3+HIHus4enY1A9pUzd2vzUrTsLLN55ZCFb
7GauHkoPjXu3TlDueRJ0nea6GfREEo9oWwBGM7MVuT1/s++DiN3PpBzX43L0LfOUymtWnr/TASq9
94chTpyZ0eHTH2VizT1uPAyaVeamPP6tdg==
`protect end_protected
