XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������j���ol�;��]�v����i�B����\8Og��@����@��S@4c��|�j��啉4��ϣ��UmpQ�wP|�$XK��=;�V�j��o��W��ɛ��d���|���._�K3J�c�x!:V����o=ʚo���Y�;����{1�)�L�7�=��C8������&�
�?�l�Zu[�)��ʹ��~���F�0�����ʽ��)P+#�������.7a�Q�����ڜs�h_�k$�kuA��O�G�!70�'r��l ���AN&� ����yOe�����T�����mߨ����˙�8F)�M�,��t��������T�����/�����;^�f�%�q���~�^L��͏�&U��<\�k��[��ᥦɽ�w����V19�'��ۍ�TZ�}*�ߥ����c��qtx	�Ȉ8���XE���M�v��-H3*]X;���&��S�E-��Qh-�öuN�#DiC6w��к�{�H&r8-8,���������d����v��I�eG�X���Ϟ��F�20�9�Y�����t��Afa�\�tB�r��F��J*������1��:�?��������r�"����Yp���
��T�$Z�S���~��!ϘGN�>�몭�X�h�V����U�^�gY�ݧ��v���� ^�xf�!�Q?�3)���ԡ��'K��d�L#e��q����)R2���WƢ ��ǂ<iҫ����	�����]��N^2�Q�o�AXlxVHYEB     400     1b0�B��6�6�'�&cy��P�r�s#�C������u��v�z#��|��T �����9�R*��8CPƇpA��>9=%Mt�*(J'K	m�௾�]9�7:m�糑�Z;���D���v�羆ko����2�r[�{D�J���qK.Δ�fZ3����Vn�	�U6)�am�q�1P�����z�{��.�ޗ{�B�_�"��0� j-{��������\�#1n���|Y�*�
/ӍC�1y�p8r�KB�+���W�az��a-u�$R�A���(��v�7�Y {�&���3I.��dnd�0�p��G2�%�-+;r�+�;��ѐl���r��(��.��Q}���U����P�~f��J��
��r�ɨfg�31���y�ac�������@B�Ld����?w0�]���)���iS��*XlxVHYEB     400     170ȇ�����D~�V]k����%{�LOK]A�:e����I
.�BA�iTo����+��_i.!�/����+��l�1&�dOc-���;V�Q�A_n�	�g���)�ԬF�^�_���/Ƹ�Q�"�jİOU�i��Y󾾃��gx:��^w����
	��-��u�`�7��%oV���l�G�8��L�]�W��C���%��V\Bn�,�x�}@ٞ�{�6�z��z,?7�1��RI�q�f3S.�n� ����� ��1��t����2*��c��:rm����&����!]/�U��ֹm���a1�*�U�����&$�4���O��O躮�NSJ����h�^N�9�FЪ�r�XlxVHYEB     17b      f0���]�g_O�U�Vn�'�4�:�e<��B)=}��6j,stPW!3�E�؝��'2uϓ�VY{���#d!I��˯q4QQ�C>�R����X7^,Ԇ)K$� �տ�~P�V�?`��j��{E#��'
�/vI>�{Ib�m�2�4�( ���U)������e];��
h�1jJ�.a���i���?N�(ަ����VsY�'�l�*��CP\
"Hr݃|������<ԝ�