XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��S�C�mO��#�O��׍l�0�V�t}@�o>�@�i`�laL�b���-�.O:W��A�Jɝ�O���Dm��GY���X���_�0B��-ףZr1��S%����ڧy�S��0�&?��6Ǭ-Vè[!��]1�[x\P�l�>j^������K��6xV�>ǟ��w�$�]���ו���:xihL�~�]��m�m�eO�m��'�6䪗Թ��ON|�����?�-��?d[�f�kjrg��P���)V�.��.�5L����o�CV ��(U�|��pz���F��=L���S�����4�Y:�68��DaN�����4]�r���h��悚�$2:�Q��G��z�h�gy@�p����Y��f,�U���V��Q��Y*)������k��t��T�
����^���U�����'9N@rԖ�
�YxF2id!u��o,FD4}F;���PNW����4���=���;Q�>l|��D�W�?),�<툼��	�� ��mn�\bf����8$�` �]��!Z�C�/b��2�_��%�<i1�Z㐧��c>	�J�Z� G���#�R�� �c���o�e��bd��~���X����W��D�?f�#�^?�Pa|fC����{,�z����n�W�������� ����ä�c����UHW��oٶ���&-�Z�dN.�R�{���m*�+?��8����j��N��3���͓O�ި��
H�Dq�Zc�>&p�T�)����%��`clL)��Z�XlxVHYEB     400     190/6��n�I@ؼ<Kcġ�/bj*	*���$��_�����żS��9G����K��}�{Xy��NZ�������E�~,���xR������?U�Rj��,o�1|Or�1�՛ߝ([���v�ǥԢV�&�6�Y1��~U6%7f#�fziJ�|Es������?�cw�1�o��TN�����c46�\RKQ{g$S�Ǔ,ݟ��[�J|�"iP��J��J�Yn�̩+�e��O��FgS�\�|=󢕤�a�W��3ˆ�����G������`��#���:'6^^~iag�$q� ��.�n,Q@Ɲ���}Z�0Dܗ�@fQh��n��P���0��1P0���E>�`��,��	��e�}xUɎI�39^׸Ӵ�־�^EA"�F?��p*�zd��}1|�gpXlxVHYEB     400     1f0ZPnI=��i
c��?�[���T"��C@QqD�c�& u(��Wl@�[��Q�+7�(,�?ރ��r^�q�]n2^k64�0	*��B�Ͷ������1.��`K:��<@������|=n���qD����W)�� �0��Gw�mݒ��ol��`�92��=�A�oV�?���1r6;a: �v�D���'5���SO��y1X�/�w�V�!m6Dz�.z���Y�.��J��AQ��D� �P���χ@Ĝ"X�����,W����/�l���NH�\7��)E\6�|� )�`�$H��,+���}'|�"t������az�"�6��?��*��.��^���Q�^7�@��b�sĔ���E�	�rŨ�����(kd�X���Gq��r�Y���\<+u�[>��s�c���	��X��u'oZ��첍]���6�����	��n� �6߇b��p7�er,sI�&J����ʿ�m��jL7!b�'~�0��p>�YXlxVHYEB     400     200���Yl��ѬZm�4PF΀^غ���O+����˪JVr�\�a��Lj{y�kͩj�H�7L���	1��(by�e�=dm/'[g�vJ	�k�j_z���c��	ԪMߡ���!.���=6��<;�w��aǖ�ɧf�����֏ꐳ�t�E�WE��VV�Fd��>:T�-�J
��Y���-������Lv���=���/�*� ^W��@�'�J�k��ǥ�Ig���뫌������M��M���A��cߵq��uc����Ib���U�Mgz}'E�"�k�t�����nWn+�$�KX������^`�.G�r���";�aE��aBo�.z���f٠�:Ј�p:��j�e	[Tn�0`�ܕ� �iYe��Kh��-��<u�f̀H|>����J��g�逎��P�e8|�t��nu�O���$����� N����68X���߫^9�-۝�$�j�9�T\�$��}�k��@#X`���#��_{�i�����IXlxVHYEB     197      f0_}k�����I�5����H �l�<҅���{q�3D��oAZR�)l�|�_�	i������C|c!�#�����V��g;���E%����gd���3&	�������t��h����� Ne.����������:��а�c�H�)ן���7��Y��!f�����\�U�p����Ұ���2�%P6���o�O�������m5J��j�;&6����`C�m�;k!���#�GQ����