`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
TNF07jgQap/nFAhsW0wnl1m4/mfLXMUJ0ZAvqbUSO3ivxki39FBQgrOpUQQRgtlCgIDdryoljNRS
VWpM9nJzHmcTyDQymxhhnbdLPXf8aYk+a3gmp1qcRELIRsr2TollGgzfz7yxnhfJ+vUoVg9GtI7y
N6FyHj31L13XwuSWokPrpiJyXxzQOVqvD3p5NAaFqXvdU0R8aQpIhhLkX762q0IL1iHQrG/binVD
fj89ZKVFodjbH0pUOIxlEZHKLVGcu+1lUL+w6ALS+jI/6AOvUO/z8p2bwEyFCU8SlXRKC1eGWpPO
/yKVk/hKAZ4gmslDNcW31KToSssXYMuvYjCyWw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="RPi4zpf0SpUgobMtGnHnU+WgIl78vE4To+NYUwMGZR0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16464)
`protect data_block
e4y8JFJkHruCRzFnLwsuNdXqCCagD4bvl6jRsxxAMS6ExuXCyCNZc9+wVUrMQKLY0sLwMsl26Fn8
wzOq6qHNojgwYwkRh72wuPPfXbSoM0B1oN0tMajJYMKjm9/pKXCbKseQfsPb2JS45rx/yzgIJ0AD
C2QtjimjyX9FTOGSNOp0eer5sdyBfqiZD5e6GoQ3e/MjMcdvzYqqHgAo+T8iKCw3UtYNLKmZp8BR
EpPyrYzjL51wu1wJWoRVAaVw1xw64Q3FMuON7SI2wLC45RFWJ+GriWKIRUqFhjadps7XBKZoQUKJ
wIU5WmRXEdwst06Hmjf5D/4eySIfT8A88F6F0MIUYukCZ/6jQdOf2sHpuRk+95HFTTO6Usmd4IcR
IZrPulCaxDozJJlUma9b3MkrZO9e+tEzS/L3UDmSePUOfoh3Y2nIydRoS8iXZs9q2LEve6mYN/t5
wHJ3V2mlLIlSM+ePFM+1AHJud6jFzYduvvSlNiOS7DzUwJH5RpnSmdmmZ8X2muQmhOprx4u21agF
XWm8qFjYLRCeL/i7hnvIOBmvlvsNDqhNUxB1/NZ35UX+H9mxe0arBfqvrggLBYoM1Vo8iCxtKe5n
bdrtTPdZhDs8rV4UJKRk95KU9SMrgEQCM4ZHJpFjTD4S8UDs39DDkb3+BXgFT61A/LvVa0HVCrvG
hAsbiz/vBuEIV5VTmJyPkM5VRcy8AZKJMmOd3dS3Sj0mVUH0i4u0naIutRxRUXPCsg5duiluKwKt
Hmd7Qy6p/e63t9YogMhVjKojTU1z0OYfGYoN2JWJY/heJJgz3Vf4/NhVMI4L2/Gq8VhwiRX2WpaB
YlNQVtYX0jlUUj1oW3/51vi4Kys647hAJiqrQ9BJg65AE+RQIV24uzR1JQII8WGo5cCSIVVuYyWs
kkHTpS4XWudNc2Xq4b7Y7PVLKUArZbiC2PFvSRk7PQL7Nc07XnU0vMhNOSX9qj3r1qk2mH6NT+Ph
SIyZoyjETtyFR+l9Zm/geCzekSL9vkVhteRyIj2aL7qT9I1ugcfetvkzVFSnW6YEBTT2F9DsUOy8
iQG5PrN3w1f347S8AKhtaNhk9W0xLW34q5xGpb0EmsYn5BbQmfqnUT9N8SidoFCEl/Ily0qherl6
1y7nT78mPanPQpArJ5lBf/Cteg3QOltQVeSFsCZSGsFH3iBipbEdtEEoe81bXmYtBsYh98MGLM4P
uYs0ADmynGikWu5is3LlrDWhClupPQd1rLYArlxHoVgT/afXJ5Dzc2nKwthSLQ4ZFI47UYiU3OVK
Z86n8yHgqGI6pUqLQNwbTYnN5IhblnfRPOgahJGnQMrmFoBGBBe0XrgUqvKc3JkdvIZdCH+vS0D6
fOD0y8dHHLPaxoY1aOiTW3ylInxsbCS0x/jhXYLqNjis9KUmGePuXiHtdxHOW+fdIxvt+uq7B0B9
CWbIB7abe3bwqXY19/UFKZ8gJyl3balhJLgvqNQXtB58o2au1gxh3K8pgT4O0f67bBGfcqrbHrEE
z28bNQyYINyVPNpyn+7JH5VjKrBsc7UDcM8Z8DPaeaTfVndVFhESeMRe6o7WHoeRt+mbCgq+5dxH
s/V9Hf6JbGhw28TP+yuE/A24fE/bv7ssgmS9r/djJVIvAdP0LGNSt0pEYA1vYxQW+G4E4VzcxkTn
73CbA+RMxLBzrDJmSWHhSsyGZhfd3Gw0Lm8u6D0o6aLjRlp3NbjxK/rFu3EJG4rxmcYrwNu4vEv7
zEzNwS+LWt1FCNWEFe236Zlv5kR2AwAj3u/nZpy7jk7kqFWo0f+cExwu42b/jmAPYtGSycz3Ms2L
en847WltolkQovaithZ6oA2N1iNXKDmqB3nSvqY9s3GwWpyPi3JZTAA+8YHgwRcpkrbZoCTo8fgk
M3FxMdWQJfCYtUnxml9831av7iqtTosqKS8BZ6lnjO9dNO6bRHsJdVbN9029RqI9eSTaqmvh5Cfx
ypc+ZdrYdy7evE7V4IZnpa1FkHymQPM0Cqf8w6ZRuVpDmvgWpFYmNb6MEVcdy0htCGAxWMeXmYdh
QIkTjSyjXhsl5DGPlxI/R4DqwafyLo9TJlgHtGSKf0DgK0jeKqhExmiiRRph1/hwr7hNl3xuZBun
eRscRoxgZEYdwKA/8bHxJZNfDDPeCQtO37uARyla7d5wgEko19cGj0wBntYPEoT8Ob+AJzP5q+Xl
ikZaIIw40f/ZR+7bjup7zP47cnBda3oqzaiC8BSnjzkMDczzSnNf5en69hOW4/Gqrt6LveAoUkCJ
HI+7ajj6/1PwmqN/L8wakXMdbFtBcDpAUlH7Jd4E392t8KnQ5CZ9nJC4ncgo1t90xzAGHLLZe0AO
Y9htY9Y7yo71llafwllmYPUeSZrjXGxmYI9c03gP0eaqdAnM7t3BH9HsrxFS+qHDktDQ5ODJrGzw
/AUZmhonXtdhfglW54WL5AC/WBskPX9hx7q3AICO43N6qGf2XVxsSz4gB4zM33Uyd+JVV4XRABWj
Gt9ENm/7fWovEHhL4XbuHozhAqhAI6L0csFI+UZh6d9OEtKMVeVhTY93CEt2CkVYVCzWOhE5JHJr
2GMw/o8cq07Gwn+qlk6zVC4ZRfZzrEaw6oY6A7UwlNUXLaq1AJ6Hr+CPJAadMwLE/usHe3ZUu/2U
J9sOYNm1GRcLRdpcPvcuL3vnC4+GFQDAU+3I8BYyRpXFk6hlgCV8PCTCCPqALrho0jpIO8DSSNIM
0yj0kNsyWqb9ZwoJ24iasfaw2yhj3kA8usxcL/1Hsn+MW6QNZxrEBu6SoFBnxIwQu3W/x4GXp9hU
1FrJO8MN07Y/X0EGXxeWvSnRTz6JHbIYFF1f1zVgCsMzKxRI6hchNOGa3DZz2i4Hhqg6BExUPrR2
gVqkj3h8du78sDtqMOlwOlQqCRcd373k5G/sNB+o37gQ7jjLkXIWP1+/A/DgSBNAJADHCjeagzYu
FtyhRoMr4NW9dJ2TmQZCnWcIq6kGlSiQyQKmtFpjQV6hyX7tTHeZu7yLjIGfVODPC6qLE6jA3P9T
gvK5ouBhlAwFUQqWsnhkw+u8O9w47xk+54uC9PB4SOkowlSibi4PD+u38VjDfCzySdUz75oOYmOK
3QPbwcfB2zBPpRnx5tjpVV7B5WiAvr76ZOEBCbhO6Iv2/qRAvRdvcEn9t0BGyh+lRumlrjc6ryRZ
h+mSIQ5sNYPwZ7I1t9oheYofwgqWK2/aqjWljQEMNNXTdEADYo0qXgdBCuk1AgDFB0j3DDij1qWz
4jhcypC5PGZEw8JdjLuTsLip5fMTQd6ejnpAfZu0TrkEThkJ1TO3Lo8qFcrIE8LzzMsHUUmVfrcZ
/7bYHuxFx+l2Sgyqjx++xv8xQ2l3J0VikTuS9hFNv9wJh7YLL+lnNeHgBcD/ILsKI35NMmTFU9lY
/QfzPFChJBjHiAV0CHnYmSDAPCh7nxeBQwYqMpEihejXAZjUOVKiYyhmddYb5x3WaMLo8V8IfR4d
bAr/myWRwCjZtU2oUOKq/G3n9Wh2bQLIWQgeZ4az8/lg8DVa5Ms83Ykrzd7cnISMLqG51wueZ/GS
v/80fL5J9TV3CpnJBnhfhWXJGvkT9Soh8ygkJD5qBjuG8AqVo/VE0LVTtQR9mxbYChNx/gUbPw9K
Bk/o4UgdSsuqwvabRWPEXGBTTTGtQp10DForv+cSYnV5K7ksldGCZfEn1f9ulitL+g6l2ysEj/V2
dK3Lec/h9dIshAQZGERLfXPNG/gu68q8Dp1aXlWgS0ttyfdjyX559GBBSMCVfcs/Syd5TGpw3paV
Fa/ROfPLFBnUKPTyOOLlhrYXooGva+T25jacr8qY5jkHpTocjMemNVE+YoDEyexqnjUJByvGAwel
n0pc5lY9Fi4gTCdETpkPXZFrSWI6GyR3BaGImnWncr45d+daMEVtRa59aYtQOhuVEixd6cuBfI5D
Kx6TmHLKUaBJ6cIbBYuSijaleTXeBbfN2Bl6djFnbGPGkKVgcBk0wqxhilHGxnjTaoVicpobdqry
ovk+BUaMSuXmbBIN1B6XXeCMCCHlCen9ca6lBe+zbcNDgv1B9+3pbVQYJ74+tGt9pmVwXkb7Ccpl
7mw5mgjRw5mnDMx/j8BKUt+apxScmZDVvkXufKhdI9rZ1u3WuUMJTQj8111plHp0AISENIkR8Mmq
S5SqoIatuzjy2ivkSBTJyp9niwEWwlGkj1Gs1kBpzR+WteaCWOSaBuQaFtJ+XjyLBvJSD5YY5E8L
dWrjL2ZuMuzx1eRHSFCGUglMYCmZbFb+8H05bzp8SNp0xI03376QfADbQUpOA6vEv3PTtBkm/iYH
9EOv42KtMsCI2/55qC/iRELl+hMwi7pBziYJPAYyx5rupYtj/08s3BjrK45f3Kbmq/fPx5DRlFBB
/vMKtdn43+292iGQAsmCEAVEQbCjDAd7grehCF+tUec1/ytlNMPafi4N1TCQJ6vV2LSgxkeP3jHG
1NlobPSA3nbSnX5eGsmGvaRmAe6pf1QBbBnO4re+z/uEJ4z2lvUpRk1iJUV1g7y4joa/qcJCgOBG
a0fMfmLYAU+eQHF3A4PlvW+Av88r+SehnMud3X+/7MsP1z7wAY88Xc4QvVXD9R82LlsqA4rHHyce
CJsqiA5EoTqU012fVrSy44PVIxOBUOS3NAG86U935tUKvZWbtv9NVWpHOC70nMURcSS6pYB6o+PV
WOe2L3XpbIBbyn3dgno+4LOC/4F+yoLXIAumbZA4uci17s3FdoO2eyJYBLOGIungKKl41Jv9xRl7
vWQpeXJAzQXDVJAeD/S27WktEHYcYFprzhgcLbrpo2zgw9KuTSPcTXP1E997kX2sq91KIn6k4gBQ
ZdWd3N85ZDOuTRYJGLi0GTB/pQ9CXquIStWoQNtgypymItKGNbU3CL2uxYgMs1TRloz5RJFoK+g/
r0AEooIda/tslwh3OfmqzJVjDquE910/oJpvAYMqbz5sbC4eIG3rvTJo/Q8PHYW7+MfBjGSnSNlJ
HPQw+Ex+9d+9+lMb6cbMi03Bo3I9FY+1jfzIchMyYNQpH1E29ly9thUMk+H81ZZFi050m/dnHWDe
iO89gDtUWbp5fjLpMzzZbO7TnuEQL6z47e7Mw3UNFNNk9icPlSC+3Bc4gX9FOPbglcA3V/1hr5Wy
/dgeve1El3/bytzAhouDCFfgXKsjM8cciePud46DoakaY5bqpQEpWfRlJCATAdjuE5XfTP7zCPH8
JSvbx/4TO/NEy+cRyBPBV1yJaXoYR4leYdHlR0bAt1nh0HzE8VrCAtl/Aon2DHR47ttIva/6b3Kb
QE+P0MEGnvFKib/r1V0GjGFxRw6OxACCls4+sGZlUWUR60f6AWfoiqv1eej5ytPDQZ0rRYTwf1Cd
ctj6lOWrqBfyUwwKu9BJ4VeS4Dn//d4FXmpgzdgD7kNdUlCRXVwJ/jFwWOkuD+MKSuDkYowZr9aE
cO/anIchT6eQ0P+a6PGVaFl7zWpL8/cYIEgg7RVQGG0ounQoR0aBKnITe6vdbzEtE4mBOR7TIyc8
IxRYSkk0e3Ib52B56VOozNVb/F8paXMSyFOiis3DAYTfXx3141EvTVeeT52skW+n5qOzPd1gSVg2
mOGlDbZ8fsNQbftQplAUz3K5W+8MKlIPA/uxTDnfqNHIbU4K9XqKXkzIBuaeuTNoQXwv1uUeYlPT
uOs+Lj7IBewM9yq7mm87XxYvWiDPKt25cyeQM1v1DPzkgdBHjT1Nqjp7N6qb7FEOKtdlygCtJn9/
OWq7T9GHUzXrMgW5w3DekNbEBNn92SG1PmO5r2tgfKe9Tn9uYXe335jzWgFFACb/lEcTbjoo+Xjj
HBnU3HZuPnIDH2AMigUTQg3W57/FwltBGmsNhK1UjnAavMBNdNp1zTzACNhoi8opDW2ApNvI45oN
3GXcRcihKr2SovXRbOvft+Y59q07w1QUuREBbNDT+abvakZ3CT06gZ7CXSFV7USlBAF0IHfHMZAD
SGNwjmjnM9CFhB3ALN453fG+vzBGZ1sa4o6s4//l5pt/W+LU+fNVPC65SdgwEIY0n8M4alsaOVNe
w62176Zdg43P9QB95qdsj9lTRweqpUnOQ8z3Lul35L87jG0CykX3ND6DcOskIRZgBDTyN0AIKw+D
/rGkkglC7tOJwSMPb8vWblakE1ybhkOFvsJ6cPvDxskWU5vmd7379Tk8+H9D3v09wtLcoAY0oimt
78HnqBm755C63sdwZW5XuQiBgeMCG32WrDRnK8ndKzKAovgtGQpBGub1IT8vqiSsWS7d8wabfXYS
mO8/PwagrMrLw/DqIumpejT1IttAaXgrcCKtP2rqm84M40/D5+MyaJ2z0ePBq7cOcIdVGPxlqOl1
+osABX40hxusxqotczr5vERsTQ+BWUVfCvGLx9SuB+pqKIik0PI+IzXCdRm3JFfPNZiKOhI3kahm
JlDWccMD/xt58+HNb1W7aRyz94SxOWTyg0eKxg87LtYLyqRvSPeTy1d/s60oVGaLt7XXNsiMBDb0
a7sZYAR7izSJhGHKMF0vEVCJx5RO8nopZSF3Ts0c/3c42BD7Bq2vaqMHN8cHP5quiGygIqy0Yc/h
MvsMfRTn3CcuPHT+YGIh4JKavvuRqPNaPtvi/X1O3VBIBSYYRFUPrCLsqZijNkdhbET104dmiCuY
vDGqFPR8j2V3cWzMcsFpizXTAELnSz96cSFh1GFAQXDpJiUoJtCjprmDNFtyAQuS3cJdmpz+vo76
3GSciYBG32ZPPUMFQ0GRg5sV0fqrWImIMdpWTCQYgN7fvOa3J8I1RgqiZeiPP84Q3hgjU+OwuqMI
S6iFV5F9j9X1j+OX+6hMhLdNO6U2RFVmjHSKupgUm96cIZjIuy/6BiL+2nbMNqtEoLCfuP+1h6xw
8bqfUYFPemUtOY/dv761CvSek+oNHw8zIl0bEHfeAl5dkVi0Q3+2AuLq3dC/2jfzyQRx7j979p4A
nQLK3Q/vtifeXArpxcoeFPyP7CtfSrRu/AqTWw2TJp7UsIjiu5mhGx0SWK1+Xpa8jZZHIrTQNeId
8fYlKm9iIvZPphu515mNtlimk5Vn234yQq8tyEJ4m4UO/Mxt2Bv7IbPHMFDAaE2f3l/xvD+rFOsc
vjePEx+KqhImq7ujvGE4F6kiFRSbWrksNs67k4PSTfqFNkhTNZjJeB2nYdptyGGY7uhS4ALRJWXO
pl+s9BgpwZc9tdc1B7nRvE6At6p6+m/V/IMDNXlsXsYWJgujq0s5NWZItYxJywWE/ogqMtEwZn3o
3eSaVkMkd9sQH0qCYFr08GQoL2YUObzw+DMig1Uctn31FGrrLtbz61U0fukThuxX+lghfAjV1/WR
3XY2KbBeznVOnz8Jmmo77v6bnb8ZfGtUWFkH6VVuYv5wZacMI45GNgBkAZOyGHh4PlBT0zOhml+/
aHEXE/1OpMG3bFH+L+BI6YudT9mZnPYJtdT0C2OitAOxg8LkG8ZdGwJjVUaax/t6sQCAwdeRNqE2
HARnqRXS+Cufh9jL/ly09zLNLMIJxJByqSxMspAuthjCQzRu6UA1SYY1mnugVRsphcq8yG1F0XY7
JHi4zy/XPZ81S5AjS7B72q+XGOzxS8ZGsJBAxNoI9UFpkaTOYvNIeLM3qdCJ88l50AhtowyNcXl1
h+atz3Qu3Ns4OAgeQ80aCquWwBK+hpbYaCUwTszdLHb2lv3xfKUK/8LBZM4WhHrBgFZJqqhylBh/
NafnJv2IJHhSBfNgGCgQcThaiTer0dnCigs2UOotY6x3YeETfPcyHtUEP9gqFLY8UuaG2NB6CwTz
lL6ibMxlheb4dpP2HqtWbnMaDUOioLEWLldYua2Do6ukkEw0Nyjua+zcAg9F4AuPIJVKGXE35PE2
80oWU8gdPYAdJxUmbYJABt7SB5g2YE1M1QJ0Nsi9PTE0Q9Zs/8PFT+I2KbwEgcmXXPI9/kjbN5Qp
WCEcuQr7vPJ3UZZNCl3OlKv9ZLBeITeG/IJGW6BDGaEyVqrtMbCD9Ak9GNolmu1lBz4LgKQv48Rz
36EIaTsmz1VlLhauUhPGUj9EuuBOktub881UNxDUMHh6dhiCF7lgn+Vasg7NZQkQI253vX/OwR71
bj3ixzmryplF26U09Ep8T6pa9L6WCnDbSvmYTtFIakZ8m0xnuAXXQrybUV57C5E2IjAeGiY50Z0A
R70jM7xXhP9ochIgZYRWRxysb8B2PN53KrwmlTHIyjKQ6xApxfddh+BepWs5Ts+dT1q9KjX/JOh1
JZcLHQzLj6ytYdMPsVKZUS2DKpxjb0pqs57oRIabVfTdUvdo1qmNFp42yXib8/V8gHL781SuDty1
ERg/UA0HhCKJqCcRve+CdHyAkiOKIz/w2QlX7N5FpLL4P0wO9RXOTsongELLwCibYA+RRSYaXPjT
xwER4xsXtqFBdIoByQBnGJKBL0QiXasxwfLElNlfkG/XjHETaTLGYr4yzZgtD5K1Si9P6Kixbmrc
CL8DZqDw1F68RoY2d9jx6NEZTnYZy78E9YGRrcH1N1aePVqfG6TL3k+3OvfSU7tUndqN+9f9saeY
2TxgiThOmQgK9QZf1mStWIcdLqU/nypjo/pt35b+mWCVgaOCseG2M92KN8T7Dt2q9gTYKb6rj8c+
vHkqi2P8ixrSMC5H2tgPtxcA0QMXDsyawoqw6ogJklGu1ZLD7deQGeWbY61cEHJAbVHAd1daZI2T
iR8yfoxUGJi+mOpkQbJyQKvhqlhv7b7wVNAyOwUsvY5T3pfZGjl/qkI8QZxl5lCQ5nkTuivsnj8K
DOhY3fs+gNZFTAxrudL0Lt70FZfzfawcV8HsJIFNVNdAO9B/vkkZcO5Tf17qpwn3YaNvGC+0kACP
dY2qC66tbRfCvYUH91jqTcdHgYonFmgmzGMm7gtsTAPa9PYrb7uqyQherRxQ7+T+ac3cd1+OzhAw
akP/lEHxjt8ng7SzW7BhKEHgVwzl0pZncgpq4E3bNybSDg1vpQ+Gf5eq6n7q/zCfDRaulBxNjLL9
kPGfx7lrfLhxrXBeJNpl4wTDqRaj3lZntk1eZpdvifzGM4klCV1zfzt9+D9FJBn3j1PrapIvXglt
+Z6PFO2grfVYyuhxHJrUUqUEvl4pv6hPvc6/kiJKZ6RY7dlkwOyWmQTATBFIaPB9FudSuyQf0nbJ
CGJaJKNDi5vCflQTeOwkdyieXoSYh6p+4OeAXRfR7XGCTWJptlsrvdyALlheGtfehosr28Ow3Dk+
qqd5It5a+6F6oWxXyyEZNT6UaGfPkhuGkQXCnOwVjASTTlmGZhRHarRL458Wyx6xGPTpnaIprDDc
5rHn7j8fyPTaKbh/DPLEU2DwCasMkJ417YcIL15ssvq5GypJsiOnLNUMJLWLbTqhdkY42qL57jKS
+0vI9TKO9xAsHjDYC93l4QwD1PcSeMggv+VP8h2l0iPTdPzPQU+0rub177VBHSvrrhbv++3fII4E
k1U1XzxWOQBpjQqxKNn4qpPGbaJ/JM1J8fgOyoTWLhMrBIAGnXzwTXT5Bfqx3GDTTfrmKdTzYuUK
qqAt3awIdFc4aNc1E0fYpl8YdPSbwT0MoFi0r40W68GDMgVl4qRcONN72+/I2q44bp2Un+ElVH8M
yc3y32okS/ufUNnuENp1jI1g9/O1JaLZNwgss64VR272MGuLX/9BqQ+V8Ls3aLI4gXm51sQy3dtR
t4pDEelxLlmJ4S2NSb+7rD+wQ7I17t4wBnazi/kfAfzZG4lj4vseYaqPc1WC5D44WLyxoaUlZS9z
GzBmqktOLJ3FI0msOD/wPxJdrmwwbzLuXuVEOKPutsumF1OMq+VPPsVFroVRpuSw9ffO07v7rtcK
DFAklcnd7Y/2XdjbI2qIO+i8+Z20L3rzsImSw9UMzWbJhE5d8BUGXtdDZWU9MdVPWsAOWRvuyHnB
+SRnRZ3VCGPCku2cDm3qIjcONnjc4L6KwG+14dTkHwWHfsx+MQm/hnDrJa4zvtFHAvUz2Q2QqSI/
OevYxlv9L1elzYUuiFGF8qS0UULbT7SKxh+cC7vv+KGYzhDOWvJwqd518ATJ2yBCjobjFTobuGx4
LSPrbXtkjxrQsmqKUaK5/bH3QPt8mQhaO2/+fxUPQM0VAON9Ra/XhN00Ayk18rx2j3WGCb/VHL3W
0dC5UjtIc9GPQZnZZ1N3lmaoXEkNVOTlrHab485AvXKn+j6t9MqN3NohKVnYts7+b3lN4TeCF/zR
hZr9UcPY6hLcPg+IBIlqQz6VJ3qGT2vT487iYR5DUh4jJqgoAI9SorR1k3gILTvbxsGxZlsZaOHe
xMuVwBaWfhA7zUnsZuclT8EqdCWAxka9ofYDYSFlew1k8UFU4Gjqxw6OhLbYSIeY9bdGKDWw10AX
bjic8O02zAgFP5o3zQ7oOPRp6NDpt769oJClw6+H2ylC8TdMdpdRvF0ccc7y0feEfAaULH+/ywT6
biGRBq69DBRzEs3BeFIvnNggFKsh7GRUPN3pJXE6SeOuqzbcNDagdv27e3iMk+NM2ftpx/6jM/xl
n4aUq+nSoiGXoJT7yX8V/7mDY7GkosSq/tXIEfI/Nmne5K2IboF0f7WfeY/PJ0D/uz335kNFocby
nncdWJUNKlyUnjpQjyjmYz2YZhiQinQOqnM/Gg3v/gmpdpOllSaP7W6cavd1jEgl8hHlJFKz+2SD
t4RAhxSTe1XpIgxPYCYlvfBM/5+2pVxZxykGdqpUel8rDtHh86ZZFAxQbwpGphH2JWRIfVHeqCOQ
9jjdwKqOe0ob45NC4EpOmz3qfucMo/Nx1y7bqvxqNDOKq7JW4FuY5CqRozz3LMLiss+QKlJ3fnhf
ZLicLxSwadYHPENfMGGthZK6HAc3d/ZBSxBOplPs3DCyzIsGZe7Uv1W8dUcMQgGmInKFA5jlVAFR
JdtSZh9MC/+ajDy3kXgLHoa6an7vPU2gZSv2yztDE45jWlEZvoDBjG+Dt3cJ9kJW/9azhpZ/M5xW
g1fOywQHGRvA3ZzSwHrsZZ08lyXMyzVbmijje6yX6ZHPS6tCOJRHqkB1RZEPBHls4HlsEXTLhuAz
nkyDYlOc52TrE2Bs1kXcUxYih6J6xERcf/50sGEUEY60vymKmCXhQWePvVZjgJDdq17vb5pZRYxz
9Hly/qHPA3fzrOpvdyidUUx4inntRQOgXOhbJ+v8HcwD8LnnHJhbn8wDh8fEqwzHyOhLnZ46xX9K
xueLnqcZTsojlsqYUEUGJJyNpf5jtc52QzZKP/akVhJO+zai6JmpPyU0mjU72UCxvYfUyYvJxRht
C1qGpg4EnwgWbAUlftLRf+k9o9H+vWkYaMVndLsYLx/epQSEhjh8OZgHWaqXuRneqHLZCIV6uv2/
lNpvg/JKiPcNE6OUXEh/ns44jpwt0BD+e+qkTFRmho2ZybFa6CBsltvcPZigcIf9X1BUrzfkpCSm
3FFqgfJpLI5VlE5oeGWHfO0QuCkXcCB97JqkM3/Kp6Fh7sLW4IEee5kfqWyNSUBaCP3yB1WbUkWc
Rzev9odKmXZYiNW74qII6Jhi13g1pC4omr4zBtMh87uPzYpCATLOZCRHgIDu+cUs7T6tt7Oty76R
WsD/dkTQ8jgOoSW5xIU82eRmWn+JBSEXxORyvVjx2JBVProd8m8iiaz9hjbrDj8DLULrtA5Z/6Mo
W2aRdnyliXSGv0QjvEfTXHf+CNK3KDxFI2xhlczJlxD0whmyQzEeqMgo9Fksg6jaT5MNL5KdILJH
OtRjyjhSU+SIfRrSD2tFO9t5JbcxJzuNNZDMPJhFcFq7VFi5bHDQGyw/QrBsGp5mL+kTcXRithkE
9ZtQwy66L9MATuDiqEquhz9G0HFqBGhR7AVprQHXpMb6fp+3AUpNBB76n+KR5r15baHYLQmKP9ao
9JyHY0Bk4WptB1n0/knjlXbvcaFb6ydUxtr+ZsucgGf0Y51Bb+HtnFs4HBlsXa1ZpucNg6PnLIWU
KsVge/dGdh29cDkFcOrVF0BhVvUT0agUGvHorox4dwElfNgKTuCTn0SXtzZ6KcdcOFTP34yUfv/t
Ps1X/p4h5qzCGwlXs8LrRRja0xIwM1qSUvD43tKAcUkHQR7gQ0DfiYyrSOFmk8HVZd4mxpMxWfKc
Khi3cAVL7aqW/r2rUz/UZdWy4ZCxfPgmyLiQ+dnCzx/8FfKMi5lbZ+8uBUsIKcRiSWaSVsA2AoMS
D2u79kGUBYWvvAjjvEA/tUNvevEQzfvHckzN40FRt7+gNtpQPG4aVU1uEViQmuB26yDo+ViuUrxv
SEXkyGj8hENjGy1qAuXG0nEIVDOMx05pQurLsiEmxm9tJ3YUBRzxVj5qxXra2J+uWZg1nkmoae8T
4wmkfVdr2fp7cuQm/Ul5OlRj0y7zD5aCU19etlYU6+BXWzjxvvx9/DbvkCDo88IzSU+ILMjDrlyd
Bx7Lh7xa0q7cMz6p42EY1tOuRak0zohiKVSJY66EFEKF//DAc6KpRx5xGIWIxqgkr6QmJ5dn7wTM
SrUupCgMsorNKCkDGojbyV3m/8UiJ41AFYV1X2udMFiAmKftQReTmxrlXXnEy8e8g8frQGQnswre
9mjhlGMwySNo89nPMkwTUPVPzGGCavc8reg1oq4JqDPWYR6hOQIGcO92/oUiyQFIhMtdq52TSis8
p8IKWf6NMKG1df5nXiXj7bL0ryjZ4dVnt359VsmWMs5RQYfXIofH/Q4tZVyuGWoAtAtlyX8ru0ED
07GAC7+eaxV634AH52XLz0u7j6ECj+iuOLazhfF2L5Qqy4gH3P5yqFighGQB1SFHlYippcbvSM/x
V3/7pUFahaNj6wBGnCns+8jJXQarEok6bkyx16o1CZh2PREo74DbTsZHyWPErbYtSWdjn6eiAnAK
G/Ik7OWyRbme7j14q9uNs5Dzkcen18P+yu6qI23OE40nJdvEUzaZPwKJdKS+Uy5+iTFKA2Tt8EFl
MZsqlF8sPIYgwTDafTQn8GWS7E4KtdEidgAiCx2i+JJTfDQz9m+zKRxOlzBQKcSWHxqVm7B1z+0V
jG6BOlvIGlSf8hjLdedFgGUnujBRNl4ThAIYrct/NKR2Ea7yePtYba39YeGFlog+Rg375bVthUth
FAOj2/qfTyOgBSGGZkcyaytJfMpqVcZGVTxHTCfXLXISvb6AoHYhnjw9CI8pjhOYCaTD03eSAuPu
O2qckNn+EU4ULX3AilM7gbtzlwCz93WqMQwsuO43wJWcUZJdOaNuzJN2rS34zYuZ7TLfk0CUM2bo
RT+yGPNDLEx3H55ZywgRpKa+IgFTiNTlri9yhfMfiXOMWJh6yitQgmmcED+cGzolbDaOzb0hsF0u
irX/f1GEcfe6FnBsCCe8vegxs0vn1syCBa4+1qqCgYC0yXgBYkKIhDXdiDDp5ChEgCQ3r8me69BK
ZL1l0gEWBunLs8klSnhWiqm9aPct52PnzU0Q76f9+gryrzXK+Q28HS6WUzSpH7JT5cF/v2uSmRyT
4hLliRC0bm61DN8tFdLC35BHVACqsoXcMqzzM+argPnBMwC0RUW+yfe51TU7kpzpOSyOMujfDA1E
mttiU4aYp4P532cxBdx5tGTPPuvAaX9UqGoBJXE2nZl5nqdM/dSOYoCu+jZ38QJJxlNN9CGgm7yD
kWCQTb1+gf1hFO6+xC/EH7OmycZzSB9ThzNDTdN0TexaikhJl4y/u9G+BL9OFQi9yYOD53IUdfhU
3iud5lRpYpheVgdXYmEnNSHrsFvRLohzcHIiFmGO9bjE2Ys+u/ZBYkgeFVvLX0AWu2v4MbqYst0D
/KwXRs0At43HL3Hbb6d8wZMcsA4tJjgtrfnyDfeEAvS3j/vYgoX7ssLYwFQF46+Of+77Aj4yuNpi
Svl7CKfUATZAZzRJRbOIzPGK3ZTQcigbKJBBYBvqaENVMOEvmWi4moGkZ53AA6xn0AmauadGyn4E
WP65cq6LkVfI+uO/VYASMmzDph5N4VKWwUW+iXj1DaogwA9ZAeDd+VtbfPHB7th9woHUfCIs3z4c
seXSaMn49A3oPM+QTrI2BCj409KLmZ+uR6Rl321kAmYw5zN3l1lbWLAst0QoQ4rJQKvoz6A3NBqh
HtjyynxxebTJL8ppwumBOSvgMMc7nRU8hc1U8pJRTbT5qE1y+RKzWfMqxefg1fRr4enqsLpB+K3k
WFjxLVMGaBQnIIHDW5QC2JvD7x0G5AeW3WDWEl5wKEw1+gSjHFzkdRodOXGgjUVez7pdkTUnjjiI
cQGoXl0Y75BS0hMBrJrXOHvTQgiFFyUvfURozIRmPhkFA5tEpX1SUbmCHlZ2VfZSGQi3fYs7WJFb
Mm76CVeJEsCV9a/BBWXE/+6w54HSlI9qMWP5nygj8+ChAQM70Z3IJ8Zh/ROTlqKUwv9uS87pBVyz
f8gDEEeHDAd2uxVBGhhIpQ0+tNhcEojkUFzc2rcF6brujL8vfdZnoiXJcXwPSae660FRrsy4tViG
2tLo3h/bZrKRMKQu/wKHJxz+HfNFvAec7Yb0BYHfC8c+TRzu5kUalRDGf4UQyuG75mv4Iczto89w
0X4Ex/ArFAa01ufw8H0Qp82/6TlNApaqmzpT4AE/9fL1fywxxo76xyoKrHxNhe0Evlq48upaFSeC
Cg7LiwfEG58FC4pizABU0YOBvgOdmxjW6Pvd3wuwEDMAJEmULlwbRbK4nIG8kdjX4Nc3JST2BjQQ
1ewym/IF8zGbEwq0Qaqedyg5bns0bgtpmh9NoszIC8Kk0REMPhVtJbjNhcQ2PfZLqn4KbhmzKYG3
1lVCpeEkB879XpzJMN0cHMp94PB0Ms8BEcavt0bdNCdvLr6VQja8gpWmcS+Ues3xKFtnjXDomkpy
DbEHz8NNsQ/UkoRvcygFR3nV0DQtHPIyPCbEE4l3sbCyPy6JYtgSghSS1CZEPC3tmDHlYtHOVEWu
gSEek3jqdaOx8oOBe4Co1PtEw16K9uR9ckja/uX8QjkLDNI8+jztnDBIkCXQ6MTo52EMpS5YY0+c
qlS0CSnqhiWbUmeut61H4mzK9AQwSuz4vz1tuxZdk2D5E17falg3AzyWFQPp01KlwvMgR5mZ7Cdr
ut5/e3Z9Hfv6Tk3YlBNUti6cwhwYrgle1pYWWV/vMWlUYvdMX8TAPTVIlMYqU5nanShrAu4kUwRV
wMCfauxH2HCE2YVDXycnoDmnfLkRsYD9NQ1bD2Nxo3Z3dm31x1aj3zftzRd+d/Qr5iEmKsSaIfRK
4wzrkNPzPvYnlq3JmoQGHXbbuTjGFTQEcRqbQDCskeMF/qNdIchlphb4U5V99qoniu+fAWEWFvPm
LsY7gyC7H0hWzl92c3TT8mnfcG/8Pvs68LC8MubmQ8sK7n6EnxK95UdC2YWjkjLMrQJQckFyd+kG
qfqhCKxn9VQ5jniqWXZci86yx53is6RmjxzZ2W6NobFFKznCixY80V2SDkhErFsmzggBMoSeLpWF
9dqJzDxcJW+h6KZg8I1oFDnIhH3zxDLu5UrJm/MKzivtOHDvYHHzPrERaejoB26yCiWvijU5sOb6
l2nvdm/O4yWftngHiSxdBxOMWTryv38VAdvRCtCZt9+yZIKS9Ex9WyKW3jHKx6o5Ck+IHVdxYmkJ
mpksaV90b14Ik2JXsrWfAemVukRKsHkg5TaT3nAeMy2uzmWm/EQtWr/OM1yBQ8WvZ9hqrslQ0p9m
BOwpNK+I6l5j6nnSV7iW5gmNNsl21l8Kno6fxULa2CHNZHrhQlqa4t8I8WWSvglR+otM2OSwa5xw
BWWCm7rpdEdFHSshHzvaC414jfqiaOP6sAGfiOq8d92gSVqRsjtGB2l4isdJ3adqDUHIEob9Cp77
PEbXBV6wdRZ5kNIpjmzAkUyhlD5NrclDUiMALccB5NdBK9qq8dvBq/IAawQ69bd4ASgMojs+sXpp
LlK3Vef0+cjjfOMDL9dhjnNj/9UgtMIJe34VVRM4UDh8A6mRNDIjktk1ihfAWDRHkbsCoTi5PxSa
KZl5FlMXYB41/XqGLinqv9K8VDMGZVEmb5uheTwdqgn+e1gTXDmvUb3rV3Z4LsgMv8LX40X5yklg
EaBGeSv5FaITtWn0TkpAItwFSK1h/BvvDZcP/xDClLJHUx7Wmzn59fDjtJTvlB760jO1iCGp1VOm
31vio+kcEekrwFtSodkdLKlYWHGwT2lV3Rp2hwprR3lEpyct0b4YDdqNiS9de7FapnRKMxuT/kR4
XDeHLSEpvrR+7nWFpj3KL6lzIGEsaoA9dzt87OWzC5wpxhoQqO6t/E99OTNdw+r3rJq0b9zm4WXP
qvUBxqRDARQTexKdvTeDrA5x+DSg7/G839MoA7rDTN0GG2tj8+uflvCsZ2hUYNF1vgS61eaLBmyR
P8zi0YzJeBzd9Cu0cJJoPNBdiauRmimMAqOFEIwJXLi8Gog05+qAUAcwydg8MJOFfeaIVqQYde/i
5gLsEz+3Pd8htLfPrBgQ47FV/c+/cxpiy+/SemwSLOo8TaUjILsKCqWJ9BpLz7Mf63c71+XXMf5z
0jNjP1ISMu4Ja7aKCduFbJatQ/rmgQCDPG33D4bsN4c/ADDcsEs8Zmo0mWpgyWTbJlfCWMZrGyWa
bzlB1wy1KzdKEcCzc4it9SeZyZoFQPXV+Ff6R1Ew7mc8mjCyfbDgQBKwCHEpPeLLLy8zqr5HKTR2
IfA4XcqhlJzUCVhwBlJYGfo+URVW8y3XHqU0DnaBKy+h417hZ8sffAbzi+Vggm093YiaE+O8ipWW
Pse/G8IW/u1XivajtmGV3oOgKVsCGMi0dQSz1qnrkiikrjncIxL62szIlz/8rbRzhe79q2eQL9vv
gFI0MavJ5S8hT2GXfii44vM6cRswkJXtVUg8o86ssCgZrP351be0EZ9iumdRAIn00x9dMXWAuYbB
Hl5Dxbc4n4mfxXyxSJBX0BP+R/y0yhlUoOTDLvwRkW0Kq0snxcOlJyV4mpDlBRFNze2B1ssT6QLV
1UEcghtQPajp/HfUQDypOyaZiZWd1cdl7n0oXdKywtXkicigHESSq5sRQooWc9/Ds3gLHTzZogQU
+RpoPyoHSovnNzngOsNlVUMSXNQVRPT86tOXEkgmJR2lhqkyARiA1NnNroK/jPUPZUkBfZyT+HRc
JBn2im7mO+Y6JvqLP8F9WjDAsizUAKEDr2SAqeSMtfjzxqcFFbhIIqusEcZK6RFvHyou6qiYonmc
9GHVfK2IOXIXWnpa9NsVm+QhHHLWq1kj/3RXA4LA4i2zJ88YkmqqtyLMvQpVkkd2F1BNePAH9AQ9
+Ah+9KKrXlVOB10OvqNmFFhHVYwB8l3CVZBLxKy8OeANYheTc3MEBUI37oD5OIKXAa6kEspKn7ow
BSh3lRCUCHt26aHcJF97pNQKsUYVDA4Smg6ySQ+kQiB/3n/FwgYqaZlwGgdIDRds9F9Q59hEK/KL
KRp/2QN+9xi9uSqggWbCZhTYg6u3F75Wm/5b2gRBC2t2anX1vAGvXzKKK5SNP5iAY8PXZfMkZKGS
VjsvSAUHsBB1gpB6h3Ui63TR7El2Wl3RkfnJCVwenbd58pBx8RtEi/wpOxsbjn3ZwE49FoW1gu+t
PGBCSG0lPlXVRLAYRWmTuRuef/iBovtczCksF1BxEj+M0YIerm+KS2jioT/aCqH1claSBbqr39Mw
rqMt4CtB9OCGZ5TV5UUN+z71O985ggIvTKWTBpv7M0vgN3Inov3EXU3uf4YMdPiNnU+5ee2o71cG
KghYQPpk3Z4T0sc2nF8KUg97HOsuHLZI2VSUs6l7p+FR0taQL18g2NLF9FYeMHjXCz6aDU+6pLan
uS+izfAyEhw/ZI5J5kG2dk+7VL/ICYxSmPW09HNN3Bzmm0COYot6EApHY52PUNeAnzvBDOtzJabj
+boZU+NGC6Ph+oyXOJSIJOcclxTKw3mgyu35E9umxufsafXuNOOZ3iC6mIgo+83PS3qMD0oACZyf
R1ddDOZjb99D+N1cPWOCHdX13YmhKtrVy4bvmIZmUQL2s9k075pQ+jNuggK++xdCH4sjZURA0dBJ
WYhpdd1dydHfA8BqOdK2/kdl66abT/4XlkzmG7aHW73PHgHds3tkBSv1RLCjaY4inc1FhZSSTmbm
/j1HBtLLErNd4+OD7VO8C63VmnYlx/1/Yn2V0CmpcmThVti1XUx9/5Yvrrpth+e2r6UoT9CojS2+
hbJWMd6splHvRipDSe2bhFn7HR1hiQaTOC/UMImvf1T4w98x04qZk5x2ExLYzvs9VZVARliTSdtU
MjbsTiPC0R80tDqXQJCyQGY+MO4cxYAUxE4DUXETsmdL9ND1lpaHenHxra05OD2VzIr7tgFkX+Eh
hfWntXokCMKheI4qKpwi99zTpqp96L5PVREVb/FrX7nS3RLJ8y3qFJqenoV9kjlpsIXx9mJwQXiq
8D42bh2eYokNJHL1D+uxhiW9sz4Futy7QIcqldjhox9KqCCKs9pJg0f+AV598OH58v2fxoQ4YZBS
/E5s9RuJ90qHDru/DmQjzpHnQCgv7IvjbVFpxWfOxRv+la63N1dOoZ/bya5rslX2hvF0BdUbHp9W
YEsrGnJRg0eiNV21VBHaEplEhoDJEisZdvq5cql0i4VgchdqZ9CYrFTt9WGEGoWTejcavojwtX+X
TC51JP3/Pfyiq/JZXRM1p3f8PI0QacfX3jPgbX8oXM3S60WxLKeAz5Skuz25+hUkM/lFpFivE9Tc
AUFfaWYd2loGlPGMrm8MZJ7l3ebdg1sGwrkjR786ffI4bku40fW/UnC61aopiDXWGVPTXROvzQZS
HQMdSnJgvjTY25riteBnzy5ygfZBDJsJagoU+zmhicjdfpgxrtJO7XH45z/UJkuRxbQLP4qmKKau
IqMxdOxbH+xQPcgsRgAYm6Bh7oJUgZcWgeLAQSncJHusFCaG4AZtX/+lb4F8oqPeLEro6U7ht90J
Z3oXLD/njkJhbX8rWJuLCF17t2sqdUax7m2sP1QarstkmFnuCE9Mq8l0+eKePdJdQk7bhIz6PZIf
QHLZi+uDO/2KLe0kudaXgOwz4oH2nKhJYXbjdAgbM5JILETjIGJU4kSw26wBoVFYXhKlsBKN5j5c
v5kEqlSecc3Am39QOdVoqQDYXO4CQr6R8sypyenslPK6p3xjMKIwZxllKLFJv6Y55YFdX3bUvP4p
bxR8qjKhov90TndmKIrOtfCaNgKcuNOWBrs/ut35kpYwJvZI7ko+odWhdBWmgMqYn/jnfvYMt1Mw
1tB6SdWkPwgpWfd5I1af11PTpArX17vKYf954B5BfYnVLQwgFfUy/LflPoPAcbahL3PI0KqpPEc4
hsAzWPdf+qzIKYEwHbNQv6KFW7wdvMWOCRuxJBrRl2PVmFujgqY8xurciCIbhALT9Rw2DIj0X4ZM
wg68irsGaKdhqAnLUY/cX6AcC0ipxyBJsAFpGM2/h7k9kXDKYbYX8xbXoq2aqnb4RBvzuWV9s6wc
GH7RQbBL5iy+VG6ljqETQ8XD45t0oTlwpPrqZsq4s/qj/EZadO7wgdUiSaYUbGcCyWeTDcbyj5nP
vVX9Z0RBME5S6LpdHulhFIs/tqEEh6DQsSxJDsrq/P3jVXRd/VatxDuQEUTRCA9gy6vunEEvSkOO
Mq1AH36PD/N1yYfi+95OHClDBZ/GBpIZ+FNM2d84uwCx7tAZA/2UiGnM0EKNi/Gc/JOwSFcd24TI
ijyqXT+nuviR9Uylm9+9okC4UwEOLRlzp/SR55s2Om72k35ocgwXWyRVuHLS/FOv5s6k7tYuUTZU
YU9sRHLU5GhLqtknjN61hUuUEhFVf3Yk09yPW2lvW34ZAE3VD6Z55A/GTRQjOPN1Cb9HS2C5TkMz
6pgpL0rcgnI40KzPXMda64lswHShScj3C2JsebJd4hfMLtucJAOvuSrWM8uNtYNYnQDspLWlwL29
/cqBp/bkc5X3185JAenwtC2wOWMKna5rpMJF9P1Z/NcZKUsRFA6eq2xP9RZ0wsy9UWoHqnymAnue
vK81gah9HONZrfRxY+9VbUxPLwRKJcaoM8l2RtsCGeRbKSoYq4EFetaqeneuiWrsrKHlR3IjLqMk
b2MIZ26RP6dpfdyZizdUJrUH/B/lvfNoNYS4V4k/xp/fz8pDmyam30eFCPyog6tRB61yaGz74BzC
xwkajYmdY8bXDS9ls8gsWHcQB4AejDvK4072eAPgwCCP9qUTZ1CH64q0NWWHeqqqHiTpha1OS1uP
Ro3FLMh4uYM1dsESlM22c4KzTrEN6bZC7y+w62/1JPg1PQxan/sIrmfjF7MUKn1Qfkbjz8ZbnKbY
uII4XWDbw08t4Vlyi1aDcWEP93CTMThn2uShZgulikDLYG3AXbo4m0sT9Hq5zxRZqAmji1H9+2V0
WVnXX4mFasikF+u1GVJhF1PJL4+1O8a0+YTCIJyDA7pIirnCQpN8UK3NopPbkk8/b9zTxpI8KaSc
eRRv9bpQ6iPIPi6FO4wjP9NzcB+ZhLDQ3E0D+THtLjFC94b4VR+hpYez8Q+seJ6+92zzBPS7O+aV
hClaX32Qwrosc9vTKgDG7uHcl8iIThYk6GWFKmZSh+iIVdj9NgVI7aG1XM++zlC4lMWuCRaVUGyd
Ye2zToCbytYnu6txA1mHriJKRtFR3IHsOaUFZCtMTIwA9VP8UnF5edYgpFsrGw19KmgJ7uwsO49I
0ycz8tPYM9ILqYm956JXnsMizEeUrhtmeITNIBe9Q6e3oyfKRUywCrXMAhjkOScox/redr4eb2st
nO2TsaNeSVeNma0myiv9lbxPhMDJ9XttFQryWDqUrTLo7c0QH6Gj3poSymP6E2zMs2DGwQgDIMWw
2in5ylDmqVoaT1AAH7mUNT62n1ppTgclOFFrHWu+TghbuOvBH0KCAWKvPHC5Y2f1MI2ko8vUh9z5
fAOcTQvPwtFI9zfEU/q+3hJts2WILw+EdihHTZESDLIX/gzw/gKkyPD5keFiZMWZnOmK+Zz+riWv
DLShDpp7zLnnnpAMKgcCFABjYpgU16vxjvcwKtl+Sa2QDy4teurIUv0gOMgpGmjUofSbHUFNg9Gw
E4WiRmqNGwfVBxZHR3vKjOK0r+4IN/wFT7LdpJdD8cM4HSbLBBrb3PP68ITRgKzR64Rr4ZlwNgi2
CAzP2LjM/b6nD/OOsMNRmlexRn5mz72W5NcIxXKpKUA7lt9Xsz8fz69r4A0bL6oT2lUABOqV8+KJ
DdOvPFhXHshgKDzBiGXeBGZLbhk8bn7d9v7uXqZb+x9CI/WkTDmuGWkrPn7ltq0FbQU+jf999/qn
HDwvtj8uZQ0i314KAuA20tTu3qmg8eLnJEXtpGY6Ihf+w+fEajZwc0/DS0/aIDCkjhPUI4WT07rj
nplVAm4yjc/aweUmqQW+mPyhr/XnETLC0ycFPXyki3bWzJA7sNh+ASthBorA0FBmrLs6FO1W8RnN
ekjLWXTW/goNG8g7emObbFDVh6fjdqxG7JnwTknQdiqsVYTp5mGHvjVin8WOUP1/XhXDYuylRJSe
dN6rw9cyKpm3eztMQxQKFUhw4w0GmhIyjOB9o+HJmruF75yoGDIcCtpGEZ9ivqvkp13shTnvJCw4
LwC02OBaz667iPsaCxGxGTwFhg2bEU9lPD1WMkH08QK795GOsnqmooe7fkhQ2pLlSGTniRzFalnV
DzbYoR93lOayS8ns3tpoej/Q8BV8fio2qwPAlDN2H4g62FoEdZw828rJXtN/DikcuEttug1iCwNx
KMsacyF+LWvB6tQ8dTKuqjQECU7IgkttdO7nILAZSjCldvhXyJrjB6sJwjijtDshW5Mo5xJoihc6
xDdDrkgrnsvV0SuEu617gyDfuf7jkum/zoCUkEOgRQiKnw9FRbrn8DGG/YGbZPKA
`protect end_protected
