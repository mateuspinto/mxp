`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12176)
`protect data_block
OIcJePc2zH/3Ot1ehQMs7qZ4myxK6+5BYlimtyNgF1+lRFcOL+a+lxaf49AD4AN+PIb6sF8dgPkm
sfRS2aYoJeJGX1M8hghMJHGOpahtOvDWTO+gpf5kpstxsO/sJEPZlppKWKz/BPG2idTqWGIx+ste
j4cFhBWD1io2I/ZK5hgBnNnA4gI5PCG21ipLGLLkxK/PkbM9JjZxXojhYraGjUURR3Pt0uDPT15K
USnxUoCItMWvjrj0TK+fAPYKcus0gGTXBAXAhj5ceQeroGM7qDCtDf1XIW2L+6t6tnt6pUXl30Wu
vr5fFosWIKSPmCJtFXYaicn9+qFNzB8d9d2TMC5Vi+XQpHUDQkBNmnL6YNnr7qyf4JjBpm15CXUS
KpSgxgddqjpm8huOINUYEnoHieTlYdkghGaAXFwsK86qjhe5WsIANAoqHqWQujrYN0mm0k4tT07P
fhp/gzKbCgQb6alMzDjHq0Ii7MivAcO05ScKFY1iX9gpNjKsgTriJhpZlNVVpFODxjvNWt9Q2UQ6
g1UYABx0V7ngqQLEijRWXZrfo2WpCKosagFZfrdm0oPYBqlCjsS0y2dapCD7HJAkfS+GRtq159Dx
/ebhIX+nlIs3+CdJ2czRhiC/UAjjOYQibtKP77cNwvLNIdCWfHG9Mou5SeYZwjWIUdweHqesL/5i
YioMFXkg6gHHghgKKpXKPYpRnPPbY1RHTQeu+rcRx8okn7nnCEmbqxDaoG3gY94de6Zv5VcBTTCF
MYE2m+joNlw+MLpptzhdk7CyYtxS6tKyfxsJMG4C7lteac6zI15bfh5urboxcNkHQGs0wZEcm3Ha
lZB2JN5pum0NQPQafPNXGHgY0Ofc7WKVSfvaIUuGahRxs5p2+WZ6LZdvDQdOC0cWTkF1FbgNQUWC
CWlXD5IHSE8vgu2zfMUXrS6shXtv0CeKdBbWy+rtIf8NzNdt/rUX2/zItkXKmo408VOir9DNhWJh
PHAgbeJFXVnwg6f+eoUms4bi4cGE+cV20rQW3luMlMWpkg+6b7XXw1faaQdPT/wWOJ2D6J4iRuq3
SSaMTIUUPSYV9xGsXwF9dvyaSz7JnE92ag4jhP2MVVofT3c71RLmhOk0e25XW46ouv9FJT4jb4sq
J6M0oWT9pojaxogCx9Y8bVo8nLV2SK5xF7l7sYX9ytVhnbw1w0kpws8soUvQUlxlvJ+QPgdc5sHJ
heN3p1gm6/C3DOlR5sy25ulrW0IvDy89aVa6+N4w+IcHZDjwWu2lcn2NotCK8eCLofD4o2hHIQOg
5KDJYSaRkPTyfmoc/RFK58ca5hki438SV7s1FsjeyWZsElDrqMo26aO1b8kMTWgJgQA3GU+LZYT1
XLTzYAyV3d/8RRP64IY9EcVxJp1AOnL0hjFMxCdEx2H4ny8TEU8Tbj9EOIVOxazg4PwpLY70zuJ4
MXqA8Yq9XeZed6LcoHB6ArpXRg3w4SmoHs0JLRZvgeuyNOHM2L8W/Xcv/UnOw6B280gxckt+Yjlu
hpmTbxtH21WEriaLhddXg7kFf5TWZbe1eZ+soFGdpCBBxbPsj2imBTkz2fYB/KXgG2eub84Wvoge
4R1kUL95oj/5GZ2ib7u5Ja29uG+VSLAnODsUYZk2m5otYwtADZFaWR4THFGFOMibzJjsISw8AgGI
r5C89Yno/ndkbNzFA7jhZ7cV4P0Y4sixqF0v66Jm1ypL+oSnZsyjX0IgG3G01UfInFETelZK8+Qd
pE3AsDHSA8YM1dL34Q86LMSYiZvmxRnoHIvIcCQc2nksB4uE+dG3MLZVGz09CFBt1bCKAcd0OOpC
gqzIhhh5VCvFhaCxF2aN44YarYTFTlIqZOTJt0rtlZmpUtAjgEsy2EGTxGRvfpi0wFgEzsw07sWl
qCRl0zx03wCPxtD7oBl5XPyUvrxa6ceUS5QvFnR+854xd/Lj8+ZhpXQfCSyiEnOcdGTXhoU18nMA
WZUnk04L87D/wpnP23ramxaZgkIVQS+tUuvr8VvQO/Sr6/ll8SqMc3vDpYnyEmoREUYcEBavIKF2
FPn8s8jtuzQrJkBgcehfRkBi0/tgGG8UAnnZJCr5i0WRKyBHzjDI0dYtqcMToeyFJjH7CaLVJBXd
4vJKQkvDqT1j+xbLGO4fpmYCOjH6rV5ryRAxcAVBV+ZPJawdDmGQqQBK8YEyuVRzUh7whW2TRScO
sIfWg09blVL5xoWr2XFLt0kGVyxO/BJ5nXYqpQlGZfNddwjEs1xuKBMCPLZSZIfEzuPopegEzM99
mgmLUzywjxNCV/SgXZWNEoEYx2+vO6gwpC+JGuBTbm0U89kLZ6eCOzJFy2hLOsok0gZVn60kCyoU
IGdtJHHdUerlGtO89t6zYJK4ChcIX/5RRK9XM9H3CkCw+kHOFyif14bynDwSFA17Jl0cEfu42IR4
EQD801XE6r42fi+IFE5f850hPAAB6aE9+/iwK+IorwFM/ttRRkRIEsQYQv6NSFdS46BKE5SNYa6U
qdfe/he9tCgm9A5nDqpaGAafWcvS3Y/aS6OvHoNN/bfymT7SJ6HNLQ73z8Ix/vSQFEKrKnBn7VnH
RkzMf5mvZaDit8H3KGDoF5OQyw1YLqxJg8LNFWe+j9vQeduk+3nPtc/OJOtFXqDqSzkBqc4+9tlQ
LIk39rJQc1tjvvfiA0Y6D1UPagnqR23ccxW1b/4Dy8Wm/3gXu66TC6NBCWX7GV+b+iKHXqDh8RsI
sJkZClugQPWrMM2I8eAWllMxiFGTaNBE6y8scDBfqc7Dk9RgmyAUaDHQi8zm9qJ+cVPFDqQFEi9O
JIB7M+EfgWNeQM6hsrr2emRvGEvyqPr9/1gye21EBnTAd4mYQXZbDGQEfqOb/t7uTwbmU/SvFr1B
7Vs38QNk+CtVQQhFloRNsV35ZwCCfmD8/PE6IWbvI5fvg3WD8FlTfDGjzj7OxUv+ZPPFUTIJJIah
bFPoNuIHn/nxqeZe3GclxG15ZqX8jmZvyRyDeWmlPg5ZnJhMFEkd2B+Q+elcUlgBTQTShQs6ZAYW
K3s70aas8wbzXugrqM0vbTSlqtyDfcj6WILDuMU8nzwrxAuA/TdQpK8y2DIUPq8hKJH+w+cSB0KO
siOrKVmW8G9pTZg0ullcD9/1TzPitxJyP7GJewLXXATSEMhDhTYrs20cBm/H2hfsjt/HhirWUTPR
uQ9EH7IWC3l5Urr0GUUBiGu6BLiMcXAGwq25Q3sfTf8e02dGPw/nFGjXiDP0oNdv0MldLjnZVajx
wfTwdQhvLRcFYezGLg5MmQo2oQhyOLjk9ysLXzJMvT7laSM1O6HzJxHEx0xG2qd6QtMVA7QJ5NGc
xswpTqgRH12+itGV/spoEuodhyNocNwM4YIxK/ktt0BrHGsOwzkg38Onm9hd9AvUAqYKe6LUPg8+
OTs7aFgVU7ikNNqADuSgUTmiIjmnyEAFNt15barCvda1fikfWR/ceoQ8SFuIOXAqDRuL6ULPV6kV
IT4Ai2GoYXRPGoALX2AT1+83DK4X1QmwkCwOrlATdWMlMhclFZ92M0AGI9sKuxBXMaxH+Cdb4WHs
0KzaUetBTN3Ahh37wlhN/ebuse/+z2SOM3ZpetJoGOEGnWvgwtEzQw2YSBDzoa76kM3R8vmCGB8o
2EUBCxE1KmcYUsD95Lt8ZwSIBrDgJt/NwKBBYBIYw7F08tnfGSZ74IsaE6YJbWi5UCIBuoGvp0lS
kVmAjd92Nmxg/rx93Z1pK8LMKoooI13+zw6mU0cIv6q7Qt9Hz0Kec2MNyc8YUAED/K0cD9GEydQm
/ML/PpMZBVG8kH9zVyEXsLZyqdBm5iGh0wxT5A04wiDhcWKwkr0pgZjAbj8FP3PwwqIoR6xq99g2
gaIJtL2G0fgPhOs+sSZIdfGJzlQxH0wcoHdggbpExU7IJifIehG6cEJ+siF/+dTMKMaoFapynZVG
r+50Z6g2jYQG2wwxGkYDvYMjKKxImPaz1FdlBh8pPiR9ClZACCXmmIgrVBHeSqlwV0Dqx4xVAl1u
qSgpQG/NjRiIMOQJf8plGDiv+TkBK3YUUiy0my05NQaTYbDNTNwGOBe5dryooWmePB4EwhSHZqyT
49ooAq2RSI3c606JqrD4N28xr9++GSyxX+56+ojHudbDVBniYZf05OM5dACArTnpa9EeJLW54Oi9
BrkCKLRq1gpBCiX9qtvu2Pi9qyFo96z/ZO7+kl0NsKibCGNlFPRkxGxpt1ktkK3mtSm6h3PBW26h
9RtF6GjgZc1prINUckmyx6/ASY15hwbO9Wybrk53LDC+w0oFK9ScyMvq/YUn7dfrjqH4BmkvmWbq
56kpz/N1Qso5Ng1s120otTknrG29k+dJXdW65Qfccv/lG2Y6fx4Itw+P9cgwoCVFsVFDfmdEVWfC
GHv59+x1a+EM515YlPcbX3bcx6ubEBn1H2AOyaemWUPDRfXMQSpQA9KT8dqYx0H+cFz7czeSvF26
pQHvjU3Zr0iRUFupALYx9+GVrvPPyYOJVfGt2Qx6t3aFLwNhbr1NiyonNyzpR1eFGYvQW+0z2dz3
0eoRTfCZviCHe6F6KdtnwYXgClF0IsZfaIZ7IRbFRAAjLKnEHnxW03IJD4M14k0cft709muP31S9
W0ItKCvurFoc5IoO+vWnuBFGztw46jyT42O1Lf22DDyW69yw/44lgj4s07/vUfZl1k8sTxSIJaHl
BpVaTNu9BiwxB8OnszJINh88hkR5TiNqoNw/vdlOPFNGnZy2Q269GzhsV8XBrU+wXYcCj3sYLvxf
7Oehp/sdMCRWInbxQJeCweketGuD2rzdR9UDW8YfOKCggPPTl8O8VRBkOkwLCfTRbrRP1F3msfyW
S/3jizYfyegNXY1OfuYlm9tGwTu7EKXtN0rCCkeKL3XfF809OSXYD0X9xzc48QEsWCjN90lPmfz9
n88upd0g5N/K9SlXrb8RLCNMsIWjQOUNKyYz5MofBGNwO0XFNfZkBjQwDePudtOBqPWpOUM81Md+
pvztkQQNl2T+zcLnsiEOtbeRJB/LI8eZFlvc/2AmuWPrrcINVZoJb1+0USlaA2OxeKbQkyvZQDUb
dXr5qT24QJZ0A8hwgvdWS6297Isfo6QKZQ2WmGhYba0FHijL2kg94gyMyO75NvSVdBzFyQsp+BvY
eccrPn5KHQAQE4M11VxHlCxUM+MK0einhT99sz5TZe6PSp6alP9KTd9GVK82/FkljHAYYml2WRER
rHfZBXZFI+4EKaLIFrKkZ8w956Er4UR/JrBC8Wev6CDgC6rsMOAhiT9K92bReXZrhdiN80QpbuTt
Xeye3dhTs8dJqDTGHRumXCLLdIy+4Ra6ID+ynrMWu778AW2aduop/Po34WjtjNAsIrJ7aP7T8R+i
UEW3f/So9pLSM1lvRXQ0PB5FvadRgAGwc3PJqbh7YBA3pAFcehvsZsPCu7SCjBQCJchlVghDXcmo
qveQtnE3GwvuGrdWTokchoRXCB5hKEOK2kSg+fgduD/ep+wofVoAym4plR3UOQaNFyOkGbbpfQwe
n+LUfGZNHXnTb+9+kpajePextgxQHEIzp6CTDYpxXnptnZrI1x+Csah0A5FHdyGnDiYZhcjeaCQB
jC76UyvdJwoW5FXwH/+/P4cMda11dD2oM/Kea6Sv2ZGUf+b3zA/oB28WXwZbxgpStRb6/q3gUN8f
M18sZ56FTuCk0E2bxGLyiWmaReIJQIQK8iyFmKDvh7kGsIOkBn9L3hfONbmBevRJMvx9wGOIGztN
4EtemO8pJUg6RGNL14aQzpzaAgADv/aq1hhcOQIlyLOfA7GhwtETqUVA+U260THnu308Wum00Fd9
hzLDP5f+KwlDZ9cFLv2AsFASCh9oZghXoBs7CzMIstZuZ2wVopzrjQr9zt8VPrHuy+/rFv2TFj7U
Oc7SPeYKi5ags+SKUPgvCnJgk8kkap1HYwq6GHTo6PorlV97octr8Z96l0E4VIxazF2vjXcHd1QJ
ST2k1aP4KDaa0pjbKtjTU2ShuSV7CHKOsx9EXqaL+YHHeP/8Jw66LeRYnxF0H0eDGCv/S4A+1x+4
eha+Om8IFxfxLWAhPWoHuBvJGrB1YEuAMyevdn02dRBvmShldMsX3MQY2DndVuDpfQo7X38H+gyf
SogiDsu1k8IC98gyS2WR2KLbNgVwCMbSLCtRyk7PmaXzRSZtGMGsulswRSkCvOPsZNslZj2WTHAs
kPQPpBWpXIVmVibp9y8LhLPs/+irAxYJazZwyt8Ml4eU6V6wPrG4rIN4DtN5I8J7n5ikfPk8bENP
LcWEw7Bzyz/JJwSgvPRXh/Fj/ES2/7CChtrjlPKWF4brlHdL7S8wraulwwyuxZPKa1v3gDkTsQsY
pw5ycqVCikkuzlzRvSiKxe1/1qHRhsfgGPL7i0M5swqmjIrW8rMmpe6CvnKgM7zWGfEnnhAR/Q5c
KJAC1468YXrjcqVk5KiCOV3nKPPHW1jhFi/fC0MDPeCb3LLU9L2t4pPWFw7SFZkjTn2DJchhKrdX
qihOTyCOEpf/b2F6sO/Xj1/H5adLCqSRQA+gsvG1gHMmsyEuMjzZPFAJSuASFRmFSg7Vzg0W47gx
sk9pce1yw54XOx1skhXiDMV78f3n+pX34XIcyVUDU97GW8A+sHk5TixuYa0usmbuVqMrMUT4BuFz
xhR77+gkwTGqLHF/9zK9DWCjKhCqPnvOrt2LH8CwFQKGV5EnhLieB1O7ycOqzBQ0MMlHqy6ajQk2
gBFSLRcW5UuRaDe7acuKsZMg/Rnnmw85hfAUxcCx+4mOW04ptHUhkoJen/WC8RSqkvu8SQ37uDhC
Oa7G4TZbyJiFplGK5v0XzgzL5/0IzGV0RzQwPmxfYcmc9Mmzud4x62/6mnvX4FEhqpZEiGrq9f6g
pCW8zrHTIV0C7FSmPZlkbo9ZMz1gwKaGIbEiw8IRYbDOO1sATfkhXjNkWPYi9RTQTo0u4CCIRNZe
WB0/eGrJ69GexpdM0tgx1BFi3puE/wGsuRApy2IOpEkcOBmW0dR5EdvsCqDpBX2i2J9W/xH3K4ys
nLKugrzsAXJnSZdn/UdCANpQ/3rALmDcx1uIHBf+4fGP/1ksA3LnJ7k714dY9jfGlruuclcUme5Q
KENVKkZzdtkmWOpVauYVtxnrbSDSCoLMm1us37ZNJuVImEzq+R4nPPi4Ff5FPuoDoqLyG4XyIFHJ
xEDVut91GfUghgWon9EGJGA59/Ugt/Bqazio+lC+taf3ocipO9lPcf8rtyJkLMRGo5x+X4WNmP53
/uJ8IWcQ5IDy6FM0weB5zrSBzbm+GHE8fS8HwAmTtVDFO+iuehz5HA6y6pSUQZca4C/xwbpLg5QV
gPPLv7KKWgZsZedT7kpE3G0Ifaum+dSTAocbxGziYXjEcaNezALt5QrYkDHTewWhdouEy3rji4fU
7HFIVLcibd9uVlUHeAmQdqyGemyfBBciI0hfPCzDdSQsuRsrjMHE1rSwrlJii/Ed86k+uaOZc3SC
wGALyflQm+GbvPLiHit+BqBnr3xENYjgmwPpiWHrHwJcNyDHuE2PjY4TvNLBBXbrmnn+rAyu+S9Q
2a1irlSsYRXXBiSiO4uQ+QackiILGKV6PRXUQax4FHebE2UEeAGBreXFqNubxKPKt0iYCTj2Wpuf
vEImB9sVXVRgGf3Xsx4YcjiJa9nVd753WZEa5OcCjdyFwYWj84U1XOltWh9ie9neVGlMbaCtsAGP
sgsekjpkLG2i7Z6e5FZxTVSeBNv/CeG0CN5lqnscjMoWopuR3Ml8f0SPDs1d7ktSRFSDBYYvFBb5
oYWfYz+6ZlMcQLYtobZ8hRWc5iWmbL1/rlLt6JwKSlbPOGbgXL6BolLPjP7dTVZh9j6Axvk1u4U6
jU3PaBCGE54uEi1muEn77pp2aC00ShTK42zw6d+PZiX2zz4sxDKWZnkzjqb28AweWkJ2SPpo0NG/
+HlsF3IiHYrx71q6Rfv3O5MBOzPBep0qcryec5DqXk8XMX8B4MOeEAC7N38+4GqSx8J5ASTiHgI1
fQNB7s5pT9vyoJ9T6l4EuHycjDesXmpstULzXF0AHA5k4Hamk/aeZME1kJEKGHM9ErKgOvWzR9Rq
QUYp8DKI6bKiQXVA/8BdAJAYPQ/ZxRiORKjSoYk16o9pR3u9FXrKXklza4ZXCoxPIoqcDtpkYzs9
URpaP42mGG5yN0182M8NfAnbEa2C0abGZiUvrEs73oEuluDZUBkDJkQcxANDyvkevssA7d4ntxXU
9P3Pjb2Clg6iZMPxM9JpGtWTx9FqNSr8beth0umNkNkZEj8GeNoLGtTkjb0IwOyRL4mj3V0KKAIh
pHiDwS1BjxBypouCYg8oko+Hy1ZxuAOn89bygpu2RfO6DJ1LkLfb4dNOr2V/4oJ1NMhSpF0jIWHe
fNNsOs+s2c9E3tiRPNnUIlrMIxrGgd4MHXtzuap5ZBG28DeeOAZXXPO3etG4ZpXLwajA63cyQNxA
zDbJAYzkxCJy1ARane9a/pzZtUMhLCqcw03ZytDoKUGpqjljCr9cwsEbxRd4KxPl+P6bJ8yMcJcc
Nuhls19lHZy3xqCVgdHEnTq3luTtQH+xdWGvP+NbJnoAJgI5/G4OiwxsUnwU3mqc8DpCWjcxZM+a
JWarQ+/4tNFAwicaZvrHqMWuL5TU36yUC9A3lv1ptpEhT4FI86KwGzyp3Q1iE79vFIGbkUJbd++G
6LCQteNPqyrH/8/Fo2aCRhqJYqHw68/PgDnKEOWv1ob5zpd1mGoCGDvs/JlLHnvkVMpFE2MdD3KG
jaqcf/uiEpncCxRL25hnQdpfPu7BbIMS4RhD6fz3CwXCX86TTjxOfEicZd5OWkEvDK/pr8xq4slj
8BsKIS6MCVdM62szqyeNwuGkHGI5ZPCRD0D3zxVIJ41bG8sAog1Xnv/RlpHbfUhhCA5qJdqrDAVU
lTH4rfWdNUOr25MjDYRDQMMNYkoJss5kZfw1EfWBEl/0Gv80v1zh96D7P/H2T3XChRP/bebdtgVZ
MLJSYuC9kvsSkQQ45IVLB4hNCfu+3xLz8lakn2Eg6cS6R7crX+ENxZg9T9tUDXn44qtgrx8rxSkK
0bwTimzppAK1ifQjA7N3+5MqCtmhJHZH1ZkQ3+uCWqGs0PD1tojHm4YbViTNXDwsOerEMhB03uBK
A49GzFpx/qgGVKJXfaINfKwPCPgQQrdxJX17mCAZP8FSX+C1j3Gw7qMB+HvSrodl2Bw0rhqnyNhM
TAY2mQ+dq+p+idW2A1ArQGQkymyVP6VdHXdmVkoTqIQLrjaKiGqkwfF2KVWnDzq2/64giGpPkgde
4nF/gMaaGEpKekxxwO4ZeCrAI6hYBNvrWgEUuH2GzYIm1bv/F0mOVg9Lyy5JMJtqXkFyjlH+4gvf
ftg2g2BWpP9TZBLfG/6I52AUrZ4sM+yiFQbTiUVJ2qabrYdOIB8I3mZFWpmWV2sAe0sTJ0onVBhv
9cJSOUq6YHfYmcwMgQgl/sSVpjeMPQDmeQBwJN3oP1cySHvx2GfD8RoZa4fOBvmiST+37vYO39QW
73OFtQKyuBYeEXkPNyz0O0yUvwKTh7011ulRpvz7v8/yEu52mG0s8V+41d5TgEgzBbWwlZywiwfc
qsK9I9cWfK9159ZZRSYIQZnaa6tsaN3O686UbCdTr6RV2hDtPQD3uIR3+2i+MT6SmYxZLYxMHmqu
TvbM76vLDnm7XdBd+g2TJ2mecPX1RTQstrxIPUkYCrS4ZoUb51I+NkW6haImaVDsAuq7Y4CfbOXC
bivbqnzWApBoGeOZReS4o6z0/RqfhWhwj0x9Jc0u5jePVvtGZpd/B0a17/O0v1WnxkvgEu3oRFvM
IOX94xG9DMg8FMh59lqfAWTY1GOogLz6d3EwyThnsORX3by/xFB+0pUMy00amAGq6nx031hcxtMe
XtxgE3mIgPPd0W75cY5kQ07PZWjJ1zgRExqJEkiafhg27fK9dSR3BmtINixFLjU+RXla+E2IlGoJ
91m8hNCsG3jIhBMNHHZtlPAE+SjF1Dq0zioMBIZi8U2sDW5k465qmQfBsHpm32PcgfEJ7BJrjSBz
5WjRfLJeIAwwtr5tcV68XtscZNy6DgbfZBlo7hXfmKWw3Eqv8jaMIuarXVqOyHG8/qLLI6iwrQxm
eqGq/Tjss3N/bKiMoNTdofmR2B93DW0AXVS14iuk4FFQ7Vh+gm7LB6t3wN1swfdQNT+TF8EyyXf6
MdFWkdx8mApk4r/8289hyJnZ4YkIk7ioWHjy+rSpuNlHpFuSfKRu/V58e2RhkExHTR2jx5ZXi52/
MOwmZHOZq2lU92GhUs4IGiDV65IbVVQ56sy7IbVIBHkFS0Od/kSR2I7+UKS/5V+1ekmtoQlOjEfx
dRD0JjABEgtm980gaEuBaz74La8OoTNdfvVieKI/w2Ybt+zgJg7DzjtvTu+6GNkA4UOwnYCqVvVn
6ox63bLePwIjKCXpq4IiSPIEuUeaUw5Bhr2iC/K4mwdqL1HFcyaqZwVFttDOxzgVvcFuoAPjg6l4
2/6sdQilDNRtsaYzWVNu4g8xvW/K7rloEUyADF04wy1+DPJamHbmwuKrtk6UB4o4O07KwLR5I7u5
yIJGCUtY/6TPkfUiXzz0Z5SJ7MaX7sERpU+ivzvQRZSoVKD6vwAmT9c0SbMVHc4kjWz9i90hNR4x
aLJpXHBrLfYXUnpGnsv51mmSvahffj5/NyrH4GB+RXAfzqQ7kXsn157ijgMksj8YAqsy+NfLxNW8
Aqpqqa2HSSS8BhcbxHAbc3Py6eUknynybEmSOajv3kQsr2Nqw+YFAjuLYupE5h15VD+E/NKxFWtu
O8OgPTYzFSGvkIYZS5vB8mbgmM4qKAlJpZFxEhukbUpEgzu62L7UrJKvjaCB8f6Xw0ljLurVcsMy
E4z6ZBtexMDHgw65hiOF1hZj+/TcvPG5wn4TMOda25jPmir5WbolQAlFHxOAQYa7gX5aSd64yQsg
hH5JsVK9sVEigHucnMVSvRJHksRrNFdoM3h/uetYnYjUS9TSwegHg6yIQBQIdCtmQ6U/+Pd4UFyy
beiqZ1sO2bu9lYPJH+UPlTTJEzpbflb3XmDNIqus5EnECp+szx65/SlKtHIwaaddjRzWBb+7tH5o
zsdVKm7meqEsMQnQb9qoCuLIlp/MR+qOpBxwGuxlc4B0VHfiRezdb27wkE13Ahry8U491lv+tFTx
3BIT6P9gep3T2cRy+dUTd8NeNdb0YxSqxYHkVRy7V5jbW5QcT6P5aMU7nlDQjBMCcqIF/YgvDW4w
2/B5eysCMC5B5YpSTuYSF8KEg9bD6wo8tU7E0iTmgcAZUWsnU2sh7BYdBGvOVOougxlNYu5XasNz
HP4Xfm2yZFqWwbtAB0EV1Kw6Fgvvv7flPF5U+1p1DEhFhHUFH1qkoH7r+UWLACuUqfpohwn5IwRN
7q2Cnh/g3TheFW7ZIFiuMdxNYYqGGGCipJrPNKcrT43RnYUB7BlRDwJrNJUM1Dfg3p7SP//DsTX9
+082opvsyncniHc5+EgAP5SYia37zxG+XXIdgBG/So40OJPDjgGzYZPoiumSI8eUjvreb47hgzIa
kANwxexarcZemyjoTGnhmV0AOpgwqRMj+DIqgONk3MnlHwRHVsH1VWJbTfNTV8V4bdrWuSeanb25
E60m11F85ax1k9S8Go/U4UK3EpyvJLaWrIG0OBxsjYcgecPrCUtVqYzLqHmEj9M6d1fUpQLqkPyB
ySnJvEsIUjB1uRKvEzxG13EFhTcX5Pqah00prvhHK3FpvWrzwU/XX2HEYnpR0fX3tXSj5dTWPvww
zjeQmJ5junirynDqpHbliNfMZ3JR5UGeyrUfs/McWWQInNd8ASKPycDGuVwJoMVC9uab+c+SbMeJ
j/Y1kFV5b/KUX2FdPpd/qBMMmAX+K/iQnC6i4jHM9Tz6Dtft4jnjzF8HbJUnLxvmWSUXb28plhGX
II9htPb6olA3ZIiBW7deSLE6TFWBaxJQuWr3Yy9JshKUA4Io5dtcBBaYWqlqe1Tnc95Y5lplCVFk
79wntqgTKzdzd5AXP+Rw0UDqlru95+dr1kv+RvB1FNLUfHfyYHK03qRRYxn+qqpAZKvhbemRHitQ
AoFSein8dnfwD1bSATK6MMpdqA6ZtA+xGDlI3l7tDIQm6vRZL8IzOLElbFgkG5rJrBLkKy5L1KC/
Tenq+TMDdD6uC4lsqTPOKAi1u0Xy9hfavCUO5lqs7s0G8ROu7WWPVUPiHtC2pSJk097BPYVF8NDT
h7Rho0q6Fz8nLwswzCPlD8Z6CFHM1YQm5tsDsg9XFSac8vWxaoqYg8IhJ0D6hdKBqjvAuqcPoS5q
TMNZUu8d5MQdmFF6iWirqVcOAJTvXdGuwawQonwsh5IK7GaYwYuhYSdwX8mrNg3rSGkdtjFPvBrb
Nz7/2SjsbE/QrHr805zLzrxoe1eo2V+ImPg3zKrsMRNhP0bOgjsqD0wQJMsYmYs95PMVw5j1TpiF
V/1pH1mqxiLgSecCLp4yLfdBdgQqC3t2JXfHSSZRU92UsNf2N0N/wrD1DnuUBLk/Zg5jAXRI0MAw
n5C4hOofJ7TxPWg+u5rzfN+RfaRo1zl8WcHLDYBQyqTJ8AyprzBY3BArYFbHP3oo0Y8qGC6AMUeU
B9zqpAKGD1eznUWkL16qt/n3EKzTJe8MbRlPY7I8NfRzYVGwy8dS4yZW65CclTWkK9FyGarEZeZl
cS8GHWJoSVtfTI8bP2VK0udoQQgvhFhHidqRECvKFe9p5V7tjxVddKzqOmiZK4jCmBRY1Amp9Tog
JUCmgSKE+M8lcfaHl78YypNXVuBX49u182yuBLLGu/Jc3ExmWRr8AIiwL65rjA6cuzxWHtUYB6Qp
2/Ndftd7OAj8IlalDLy8p8iAHGshbS9KMjKj1t6/qHyqT0yus0enU35bdoCsfM15yy2w13iTKjry
4ArWTwkff3v/bGlgT0NZQXZHr3cSvHSv1tJ3zAbKvbG9bDoqauTJgIW32pJikiNvuMz9RV07xogJ
5m9kWE9GU8bP131RZesFaQK5N6rMu2TX/vZ2hBYApsRIcnPn9cRiIT2zlhyS9FhI8duNuBPXEGCM
dddLO3RAHjDRsEJTLfVIFQCSk6xIxdnINHl3Bnneyp6gifGSZRWbJkvF4GKfNN7W4FJ/v6MQKLe7
vp7Y1yMpbGdbfCeLoa7m631tUmojhh9dtaMj3pznwZHMfyZYC4HwyTnNkSiUjKJe4iWsP42Cfvxz
NpmAJ6GOV3/13QFYdAHJQOITV8TSEvXpybCHxFsbF4UG6ft0Ot8a8YkIeCA8TCUvkIb56/OC33qX
ZnH3Qf2DPh2+Ry+U4G6bWke/MF9TTs3FYzmQ5lvHjsISngPbBtyWmv1nVd6n2wPUCF4/e4x0s0jY
+KJRLobs8GItQOoE3cXbyjFD5BFBQ0kg8m5syIuiaH8RnkMOviPS6HqY/tTVa/AoZmdhpsbFbJte
95iYG2G4GqvDcHQKMJUYHRHH49p36Mo0kLJJaYxQZUoUz/KuB1DnXa9Gr5CSxPEWlimb+o78yctf
HlU/FTZtzk3UySvwVqnwdPa23//0KqAKPbjPQhSVcFU51sFGmYPAeTvIHcpcM3UKF7By9hZGGfTa
6PukAbeWCwczDU7/ZW1AVaIa2B4YF57gl5gzBXN1jvz3ule0X3L9OOQ7MRMyKKt2itaYUh/jg1Fm
AigqzEHydH5uOYnPMS/dOEza6se1VYEm1AH+YVVJAhy0AWnix1/RGMjsF1t4k//JNCxul8kHVAKk
17gR6p/XFD38Wln374vYnrA2isnJbwCyWRjvkbWaQ+y3VzLqIgKC5yU+9ok2SDEO9NYOd1U7jA0R
Gfuh8NeUJqqPugv/zM+iZuYOr2/3pUepf/GTMGQ5a6z3+KI0/PEBZI9EAetengI6T1vKUi3jPGmY
iVv4/zmBt71mCZD1+hT3cLInPZZ+3T9nO8zM9ISWE9P8bsw4gGg+qGd1F4aIN8j2JbfQS3afWQw4
4Bf6oXj/1hepqqFwnPEUTw/4OZ7EUcrN2SQsBi2d4e8r4j4kdsw7X3qohm1rc1ADEa5p/vHL3aWq
K1QxdsJy/WULK4azhPmxX2sOJb4ErKcyrIygTceNplgJ3UvBCyrk4MbAgVcotA5DlapJ/yn+9id1
M7UDEaF38ruvc0a3Pr+Kl0j8vMXvrThnOGCCCtOahT99GGL3OLl6YhIOp0QVH4DKkM+1+0H6oQqH
vVychLaad7sylqzyL3tK67c6W2TqvwBX6JGFNzmVmnVacY2wa5UDzuf1roSXUDF0G2F9v8PpkXgi
GXG3SX6eAFQ/UOny1W9QinN1hWRFgHCieCspA5pi6hpcv9UKeMt2/PtsZtNJ0DSegG33l1BDZM2Q
lx6YMRsldWa2ZLLeGuYhr3mop+XoR2FjpL7zC9JouB6gw1tauNyVi5YF1fHK50vK2JN4Vdpwb90K
uE5m/eaUYYFQ0Tb2WUSODq+0sCpodWL1XJMjhLYkiIZbBxByS+lLNyoWTEFAKqMQ07aAgDKtV5kG
DFGd3NtPz//sp/G2Zv3W/hyv8tdrlyjl8hqvi3x2ziJARLkdRLoj/kTW9UxXMs8Sm7Y1ew3o9xC2
6lR4sj3QWl1fFEzEw+Eush9tpUhs6/bq+Psvr1IJfOKP+wPMH9jNHDtdOFtZ6efFu/jVRpCmYHhc
Ur9p325BiQJiCYGBQOSYNvTwFLJB6etyUPpOhfNQrgnwrIdrN0aFX3vhtBZ8zo8/3AsU1abF+Ak6
WehrQ3Pk74vOLIlGUbCgnY7K8h6yZVoFPXTEKbYUQZlBjjcD1lR3cyGRqJ6xv3l9HsOXM+A/gCz7
7Az4Ia/SgsfYUt+Ekz5J0oQNUrGyptG11Mj5sQSCtR9pr4LOttxYJ3zhEG5qwekB7gPrKKvy9YKo
fyQSy2MX1dOmINYUpuGlkcmbWXga+yabQYQPHnkg8ylB03/n2uJc8IXKLRIGpCis14nqAdShWCQP
cIX892twpgEHvtBXvCKBBVYyAt3QyTFjarYusoUBcouNA5HS7BAjOWaPgz9+c3HfdjpgPnoQ0b2Z
TJDNmxCoT78LwQDG1d6hYXWwTHmbbpXiRUVJSnILycpkxo80YZph10EHPk/8XjCQeiUVunBqV89O
txFpuqK4nqRgskKzXW4Sl3GHV81SnbyxDiVvMxfjGO9Um9bFO+uNqpMSwF5tqkh0TtNN96UmI7vo
uQLMywqrY6jRE1yQ6Ei/eiyb0nvjndy1FbTmlawXTeFM4tbMqfE3qbMpbMyvbHo8Vo1d/exDSVBh
zJ4W3BVcTj1PCa0DNfewg356VJQ/h4R3fC6FNWBw4IuQz/stawZtR1QCOs7R52+AhDc1ibb9p+9w
+fsCO+f6dT03zQA3bc89rw1WYZ+XLDFNUC6q1ysFEVtxmP0QGh93WdXZ6HMx3d2V/wEwG5aGAoKz
X3oxNbg9gwPTCbwA7oPrCm3JF5OFu635dhTUUTq5d1hNshNgLI3rh071H5gc5FSH5nAG1yUUHXy6
IeA7xY3vhDIS43gNMRMvAswAzwyd8HS4Gi8CWIzHeMpgFgiHjEnBxsp/7jWOfA32ZklH964cLKLw
cGZK8XP4HmxCtquXjHilaEkABbIIPlWlK1FTDdXbuH/51iaEGO/gtzTHIeY/z1pPOSSZADb0HaR5
IKo17fhRvMBxRWB8rAzRXLVXDi2Mj2S6pMs1Kn+vItUaS9Fyj2cvj92KofMjfBRaG5eJdAAR4aH/
/wo1kBmsuEbt5rAw6SaHcr47qYAlOxrabM9C6DN7dLOfHukHwg0NMvlFecelnHsvew+kmanw103I
GUcfyoOY9J7Mzt/IUbbd2hE2+MDiFuyTmQs9tHXot72tFKVAgI1zZEor1iehp46jxxVG9fkZmWVd
p5SSlXF7gmouOg8GXbmzZUPdgy+ZJeghMlbD+Ay4xLhyc0+g0WCd7AyUWEeCDkWG/BwEijsZptlg
1XBKf3Vug7s34vfUz4Odz1O2orOPaLvYtsb5c3X6zS9aeS174JkyEdapXe8Yu2ERqk0/FwjyTlOH
aARyHwuIVTsgJW98SNmWqFI4DSB75bqntbT8w/g4wZw9utTJePpdM3+mGd8R6Pz9JYunCmv7ukcT
qH31ajAuzjl7VVhAV8m+AAvNXOOH4feuwOKUbKRQBsKwbZ4=
`protect end_protected
