`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9152)
`protect data_block
IeD7QnSaLHKmI4OX8+ZQTCgcpEglMphdBajNSuJkK5zmBWSz3sCq8hoQYNTl+Ngx9qZal/5iVuhM
GpIV9rP+AHuuvo8mUd5mQ4FzlkHRnyl6OCkHOyKyp6hgNgwjmbguWiJfErtbnbjg2yHTUwfn7m+e
B14FzZmQqj7pgxJWbg0sFYQicWv5EXBxSAioApP8qXOJeKvJiTNUOxptP78NkpM6LV7uF1gLXfdD
hPAxM4Dj0Lg+Z/+9eKSTWjXdzCnGePp02iwArgx7rTbrH71D+5yZI0/R9TZdi0JKMKtyy74Rqh9S
a8GWBIwH/pcoHnAChbbVzpMH2wEmGrubimL5qiZ3cLTO5ssA049WbEocOsFE74GOu3p49B7fH0ao
PWJDar1AlpbICE+aDkoFw7ZAyvh+WCyHSdXMwfixOlnnatvolPkvOv8cFfmjqPFtgLXj2HNa+H8b
HdmadWsaAcqqnR0Ds3xAoeSU+PQHfFctn7jyzqi5t+/UeQ7drs/oJIMRKQdst6YWx55BBUp+OOX5
CfhKdD3pQXpdZsgK304I+owwq+OXhj0oMcexcY39IiweL6uIpeu4Pl38xqLfOyePK8UFD+NzfniO
7KP8uocGDPjwlkiWNKFMUFm9ycTNqh9JL8+8ZgNx4mE6sSVzAVdlk2sXba0iGU9BEB4ZisEESA9E
K+DCiSjp3pfWO1u10ijAdhxgKs4KdcMz5zZZD6ip6BnlAkSie2YYXM2sd0R2Ag9dPzh4pDdm2Bc6
SXmBcF8F+0l1UASiVRWhihbp/Og82t4FwuM5vbvawVMo4fSm1jIT6KqnlmYpykWcYxm76aSBinUZ
x2m5Q18DZHlk+eWlqxH8+i35p5FbW7V58/V5NrFwgsiqRJcbcSpstOqYzi64OsgDp/WlVA4jCQbZ
nbGA313hNVmVQIMIjuKqch7HPY8LICzFzI/G36aLzpZK+sAQ9Bd63tXAg46u+YxowmBYN/OCO89w
uxUoGVftVRgMBpch1DfjEEFgBGe57ybA5mCI2gpyexsPZ+U7LJ40Tn4SegW1e/fl8T8JZBQPD+ua
4eqL5ZKLApFE46v84lktk3+EuUL0F9dUeaDx3tLI7MBa7SeLGzZ7HcKiWQLzeED1RHcmHfaFCtZa
a4zZtpIi6wfcEuRzvixy4p6+E8rpdiLGuqVMAyemDdn8rF6g7T1eykFhHsjwxA6Xys0GhuMZIjdM
hG8k9dgjktvD3OG30pXCBihuMDa00Rpd4RlBq5jPXlGGAaC/T44gjSduAXNiJtIGMr3WMuIxsXMQ
tZoLFS0N1f+kQFhz8k6sOKVFHUf90tpezEdKAy5Sdk1LyLlG1f2zVaVLcfvthCQkA0wTpRNPveM1
XJtmW3tL2uzVGTfGC4qGPCbRB+mmyZmPRuFX84t1WULJivNnIdH8kB+u5DIrjWjXViOOk0Ffx9+S
kGEesKKsA/8Yr/UqS0vdJS+D3Y6yaCShSZcPq45W517XnzLnYFGXEhRzr7X+RwlaZGIenSV7lD/D
5DbTJyNDNsWQsv4lvIvmHqUD9ptwb8qU5Pji7FRVLk0pVGZOic85KeVc3qBWkvov69MzJ946/R7X
/KdeT6Oe/6GJrxmROR8uKwwk2H5ZygPYO/zxuAjjzhwwG2BWkOFehViqPgDwdBlg/mgCqrfw4Rt2
NCcL8s/LYjYEDVzkohmUCdxL1NHwvxe06C93nJC40RcxRkURTi9uMt4572mSpmqrGfjKUznOIrsd
U3kjzwqWwIQm25vUu8IPcV20Sy++pYutuzQbASU9nyB/B0vXcZ7VCdfdvB7mfYGtMfIKDCYNGWMT
YNiC3oKgCjUcd9QTyz+zyKavnyiRZTUqggPqoVwEYjkaxrKajTQcDnuMy/fs6c8idzYKQsfRsRnj
gVCz80wAkowzrSM14KXJHAbmB+pim/DtjnIcTsnTURN8WSE2NjqYgXJUIYVDuWP57IZ0dmlIO1YM
ODhNCl5E6WS24LY8Bbi2cMoiV6EHb9t7awjPb3lCc3iJz23gR1pgNyqs+0gbDRJ7a2lZe4/hzdCu
5tGRmrXo/ro2Z2aba59/yzUv3dQGDFruUkQXRAnwlDDV7gvKuZYR87x4rFbUXAnMlB6iTIaNEauW
f69+aLjhC5jA56EkgP8UNLOLSHGmIdGbZD5Nr5oO0SVnzCY/1NajN4JJNQNzSgNZva+xDKEIIzUK
9gevpWRmjwvl9/SbLPI3hf3JynrXBQPGuGBEwm1BuL166VxyrDDC4WLR7bBh0vdRiD5oEze0PUIs
Ye1fubWr4psw3/uJh/MtY6B2KyCtlS/KeIrWpc2KSQ4ReUwackOS4fKXfFVrN7VlaXUmjtdVqV2i
UcvJsfAGsWLgT21YNU4xcKlGyW7c3pJoYzvEsO77hK125lyq9QDWIw0BqR+VbiVTysxPNNlPO7zp
g0oyZhzM3cOypxU0qbNxn4F5r/qplRFjBZqhrn3iFTwjrpdZVXRc0+TYDeJ3IE84S6hzKxyddv/W
TUCYu4tiBEDJvFGKHQV6QZiqHsXfDCNuwWgtUxh2xG1paIjzSGxswlXjPy+aJS8NHLIlvUubj1ET
0Fc/XTuhr9CPrWX0A7IVOGGQqlx2g9DYy8Z7ZXjI1/jhgkdzsQ4d0+O6UIkjwPdaTx28CbDndbSV
wckPV2UkT8zgjlN+5KQ5HeAAg6TfL4zQJZiQakfVbSaHCRZiTsdRWPAbrqNydwcNvEvSK/9yEfXJ
cv137dNlCq4kXgB2esGPhyclWCTyVxDLsN5e846/sf49IUbROr5PzxSCndNDMCiK3j01GEpM/+sB
1YT/Yz8mcTSvKMCLMKBBIO5tHMXhKHWsbDbo6y6YAaoaooIAxFUA/oG1s4qf1VQhnX/kiKg4rK/8
tnDrARYcGGew1jfWw8QbydO42E/JbwrE8QaGD0gruZi5MFUPUuF11EbOi9TbJ9IUar/bqSATa4X0
7Hk85GJdDZNBbfv61TDXu6BEMvIZ9qe5RAnsreZl38UxYU2myjSvctNVjBUASAbMUGc1jr4LkmYa
ZZdyRE6JGQIK693fcjdUiv10+z7l9c2lnOjvN1pLHlHCNK8kz9NyLiJlLMxe6FpXP/e7CSD07bop
DqxraA16+8XhGoPWsRWpmXy4+tpa0a/BmvKLLyro0kRLJ+W/2cOy3PaV2qu08yx8KeuC75T03LBy
g5RkxBucWNRzBDBo8pIcSylvjDgwFLkUl96gsr0xsryUweTAKRQwqzmSUK56flxJ3EMivtJUfeXp
GJJx2vpwxMsZ3jIuP32q6mJDWDSBkHUf4d0h16tD9KQ7+JvlkA2Ypdq7oRCOlcJKVJxRlNj15GUg
Lt7PEXEwsMRXy+CylKH3sAaX0CdDFnBQ7eH1lWcBQ8PiDzYs6zCfvofqJwxymU7GZ9hk6A1vsSxl
PkFTLv3EtlKcUmnaZh3lVDrt7nfVri44yZjDLaihzXq4GtiViRCPWx4Uh4F02oXGrfKkCnQIuL59
gby4TEIOmV71Nx8Xr33fLv6ANd5KB2yLF2opTF3bT2tHOV6OEEv7NrOeiljv3R3vYGND2ftc1fn5
JSZn5qYmD53RiqzJMg88AC2jpZ+rpjuYhK17NtC3Cs5T5aICFNj8HEJtlHcYly7R3hwEbzJsgIvM
NkJ4P3H2iIJu/XgyzzT3S+YN0aOoMFZO7B9lnKGHeiOWcS2/g3N8tXM1ON/vIHd3Vw1zv477bZQz
pu91hH0i0dpJzzwXTFyECXEU+H4L+EeWPunB/1q8TeCFRgyFu+2Fr2i8EAc4UzrWaD1omzmlyZQ8
knhkfQlzElqNeiS932o4PSnEFHscjmEndFmWeqnek89u2EwayW1bjWpMjWknxF6rVwmgtvUb+BRk
Xf1MWW/ZiWDgyQiji755Y2rf+zncPICABWodPypG6QFwV2a03LK0QF3/0IMCHnM+hgmabEIkA3WP
yyIQaNI462OOdDu96SwY3Cabz3lPrKRR42YLj8iR5/d+c1D7wsiivTgOJNVjU83/XSXgTHIVJkqh
zMrM8Y1zfZhuKnu1o8E22azfhGg2LFKhZhu/WVXuaxU5iSxX8IoXBM3q0Dhu5jXdSp6LMneeh+Lb
0HL+n6hpyb0IEEt4L1GAw589EiVAWwv1V/wjNr/KZC4HDn2hoxgBTnSsLRy5JA3YM6IqGTo4lESZ
waBxXTmkfNkJy/meIk+7ak5hwC+5VBclSlnzpNGf3cv9RnUM/uXiyX+Hc2W6tMl7SiAJ38z4Ccbz
HGGGfd+zeYTtN+7fPMxvwQmYybC8gqVQIVbzbctQ6PvxtqY9jCagK6Jd5KHWySXkG3OJRUiH8zO9
riW/78LXrmKbRfNOiP6De3CJdXOI6uET/VjmvI3YtU5wTWI5SSNQteDLwJ+Si2GJBvbVrEDeNcIz
49f5kphKBPPX9JPSKPKCQ5Ak89aDJ2/EyHBzHxDl5rboawmfUiOdZsOy02Y0seqjM/aTE2CGDh3Y
dmbBA9DSIac8a84q7VBM6EUoV6d3LHXQODKLA8na/GWFRMFrX5ZDOmY1KCuW1R7tFF+0cKgpP1zu
HecgS08UFEgn83QVWuHgD2sgeSgZNYrEHK5ch6lCl19PjddVHLxtJbX8+qTk5hh4zqbivudy+MY6
LWl/OHy1U/f0UZl8djV8Pw9VAT0MnYLx8S22yMh++95vihmG3WauQ+56WExXuSHflF78QfF4vudd
vkJjUE2Q6TTPTW9zWbC4rSuGoDkhFbHsMLiIKz5HeVJ8N+uugsKTrg55TTQdD6GkozlBm/TYUSyG
7mzSjjdtoJUs+DEiTk/21VHwykd8vDBYzU/xxs1yzA4rB5+Y9jrc2e4dyymM7s9pJ+kvIbk4lxhX
teHgtqvLdtsETyrE1aWXrkBL2aYje/UoqRYKBl1/JIkuVavRDO6Vs0UXjNOeu80Gibv2IAPVOUPq
He5wjHFLtcQE9QArRYph2HrjajfFMSiqWvzpwYrHS3qzZQ+HlVV3qg9/BOX864MmTiLFZzI3rvOd
BhZqJTVZBD85qugGM4f1q9iXxJ992swpViSAj6Y/OIopprTAd0K+Ihf0vdEhB6b/QZztNpm0dqaV
tQPni6GdzVDAEtjtJcpdFV7nwQTT0tVyjJBg3nqvby2KsvCBnRSzE/Qru1joyCXdAmtr/w4AkwMX
mZCfGpCxYj4YPEaU4APnqrCMrHLUD816OCz4q5Yf8MKVzlatx6pdrszBcKhRZ1hVbO0z7lW1BAB8
ujGjn4/SsIS5REpUJFSboQ9iq2J/nFNsu/9UyyeiQB5IJDMjT/ZIR+yhu36B+GG4I/XjlbICvfOT
N0NgXDSIp9fYA9b1XevJMAd7i49vxJS0Q+KcF0ZvCQpduXH4STthlgmCH6lRVSXFn5gerLcmHwFm
pA+1hXZmvYMwYouVbzjh6TFjVwQY7pVmOlkM6+hwXGCDjk6XVBsu6U59roFmhdodWtDdsl4xwQsy
kJ9SH0xPBbOTeLxP//Ks3PKvCAaKz2S0n2SatyYIFlKLnKMBtaUcCGE+SMwMh36k8hWiCDPyBnaf
GfcmzTHKvVkuY4GNJgXrEe3JKF49a0xP3iBgLebZ6632HBYwmhY8zmVkKpgqDlDs9jrc3ECA/dNo
LACmg5BVPGeWHNbQ+B8eCdSWvwDxRdjx31zMWxtUs1BsJ6La2f6jHrcMHR7IK8Ol2JfhoJOeyNL7
lGMwXGt2roGVN41DJem5ejB2zRD/JnG8ohJj+AEaLkVH3nwfqT7MSONUjhryTFBE20pe+TLP9LX8
ihC8UbHcCdI42DZ4sqtx38tvBjmvz+84abTVI6YtY1gSSgLy5WYLb8+ndC8DW4rdvB13y5V1DaE0
1rz/C9mNVbVUh9JdIiHC9ylBObbPdGHjeDOZCimgbw/ey89+SeT+qGv9eKA6XS1JH5d7fVnqKaZJ
4M1/M/OD8+qW2RCbwgd+yqaO2EuVOGrfvM83HF/sXYrRywL7WjURdZ/iYN/XEX9bBto/1Mn+3DgI
Hu1RfYxzcSRL5/EO8cE3JK00zDItOqP3GJFLdAzdfu8vMLCr8LM9vthcswWO/7vkVeD7t4SoIaV0
y5OJxZN3Xfom2XEpvvoOX4w4Om2n+fENAKkJjLim3JoPiYyLaR1A/t8EK1ogwPlJBP+rmNcuxdv+
7QIKDUdzHUGuWswWGQQt19+nvl+wqCXCj3t6DAb8qeqcrXlEZquKc9tO04hB5vLdqkuHHr8UykBB
rSncAgNbcxFjZ2pqFeKbzkBg4a9kDqQ0fz52b9vMVmV9hBnyLbvjFi00QURa9Y/4MLu1+NPuD1Je
h+nw6eAn6Lr8pF0lDBZQ9QHFtjb4ETckovN4zVzL5wRZapNl1/gsSYAeV4whMDfGQsAwLFvT53eO
I3/vYN+JkWAcWgO2zem/Rg3tB7p31NYEwnJIcI+PIlfB+XOfqc26PXrKi9fYeQ5rzpFKtAq9akJb
i9nqyJMROgLfWQrEI4r52UkYb3b9PiFOcNcGGHtlIAB+02YE/gGHeml50T+54QVEQdg/JNh8nAYb
r/Fls3ir5+RKaajKaK4Mnl0HMyGEvcMOxMO+PmDs5qrDUFHNteIvvduhdu0MYcDqHH612zNeP4FI
+GGBA+n47oU8Mm2RMbAHITglXk7XuuNLx8oyAvw0XJKXxwtNUwSVMeETu6C4vf6JzFWZKJVu+eNG
l7YCyHt3W7BwmpOX4AHoZZTlH9YkfEABQFgisWtSjYIaBehZsC6Z/l2x5WB3DbaBbh9ft82/JWCb
n7LX3+7KzH0pQ+dRz5Hu9QsNTUmoMkMpBWpsllQjrWIGPGZZX58GA4QOF5wue7ROkQlpvBjeQuTs
0swdUNlbKQCbkOgQCbdorSfQPxlIfAiWfcDQ0I2plSCwHqQN6sm4tC0HsxCUZx3jwPd3AxZdXDDa
XMEsrTSBHiZaAxTqwHAhXdU2RvJBWoQ44krQ0t2XKphjWEadz515/VlrH6qCniAHF7l4g7r84/jM
lro/qggmiZYEwMEJGcfqj8rq6VyW2ABvGvbOttfs914DTY9fEictFQGPyuulo6/RZxBicr3UDO+j
Y0jHyl+qUSeyLKeOJvguv7ZQ3NIXCmT81hFP0HwXvPdEZgOqTR+bHQQYQ8Z+KZa+h9mdIAif9mKo
alBFaDnK4UDoce7k3acFcT/ehpJADLdFi9VPKQh/S1qOq7MbwsMLqJ/2fiGNRd1641RYssB1QdN+
BbngEHG/iNLxOTFV2p2RMaVuEJYEDODTUKqbWyNEpFAKE/YcyF+Fj5Z0Vo66rJt0SsdS5VLaFR6G
KfQPnaXcnLo1YTPRxrjrvTnwuOzfetFkG5bmCnbwzcCQ0TlzGA99yjbsI+KKkq1/Qb5SMPEqwa7F
4CVK5Vc001HBnw7a1tZTZnSYsk7ge9RlF8mwzkPWPov+n4M29tfQnhLIsZQuraGlSAZTxulgPvp6
RNiD7gCAWKNLOF+If4H/R+xB1hL+4BetF9PKaTMN/jLMg3rTFb+rnBhHhzif/vIIcqK9yKCwgzv4
c3i9ETIpYmq8oJllz7PGwzONhuULjw3iWJosDfJWXDYOHL2tBKMEtnuhWP66fKhhhoAoMD9qahl7
tJa+/IQXvFCNS5EVWLrkNo08nPo/keByREwHYfigqnLnDd6Z2C0HU50ad/X5aHOdk9rlLrDAPgoi
yBpWtqX9IZcnL9CddhjE0+uFvooOK6vrnDaiq07LCfV3kRJGZ5JFbxGFzbj6irUd+XkpvXTV/K1T
AJ+OhNOCFVpEeba7ZkxKLEvH0YAAiFbPaYjCIo0sny2og9OJx8MSwNRK6/XcBjU54zVg2MmhLGuR
xLJBi5LWzGD3aVHVazk4PkdT4GH8+F6SlHnltRdevsb+7Cz03ZuUrwqcJcKT1QhbFQGhSFIxWjZv
fKr+zy7NtBrjJBP1fG3/LFtoyqS/JZB1CihVq0f9cXqqrzv7pRmm0qtyToveS3ocSg2liLC1XDfi
es22zfjlERBCsNJRVZZzwG5cGeb2ysagHdFhj4GqgTdf2a86yiLpVN5LUp0z5qH4wesfhJsEN9Bv
qfT3cuJloQmv1wqvVRAr+Con9yRzaEadrnUOLr+4UugDLBZuKgP9A6FxombHWfWkPgthvikP+nsf
XCVUoMXg0vaJ88ZN1EbJXG79K4afbgdJen+XH/R2Y+kQJUdnc94tNp7s/2FkywBG10/mQEnAZuON
JmVzmfPudGOel7kbmvvEkF9tO8ni7h8AmcIZsMmOUmKYoPSOJpGeaiDO994LmI0gvA3qlOSo5Xos
MAlMOYa5MwPDkp/sunz7iYWQbg0GXQ2N0+6LVUijsJuE1IXMOG+KHlSTtvs4PjSlV96KUYfxpKuz
cRuBu+96sGkS4msjCZ9Tqc3Qp22ihxLhlzWfJe2sKDlc/ZKzxCgseF4TKxW3x1n5Vl1p089LD0yJ
JkMl3v06sR1kpav11UzJcDzY9VwFotmKJr+2Ek54aA0oyCTwK3kqwpAqE+kD65iBAIIYP1D/8dd9
YCwx69X6Vdj/ieO5YqJ86v9gAb1XP5pIvbbXzqTbkw5PA81QpTLO+xIHNKwS2avSDZiEy6PIRP+v
dI3Bp98bifdhH9M8jMqkJAxNMuNUX9VIy0Qvx4oiCjaLYBUwWfIj1zyZ/vIhZ8yKDVLfToy8tciy
GlECG2cS1/AkufTyxGWEZukNZWGLNEvPmkTXId0vPImXrmuRc0qNhyKfspTIn53x3xWOKnNH5vHu
d1Z098Abzz5MbUROjHQbLsRJiy9L51umjkHiCu5ud9e1O8OwnHs8uuWCkzivK+KhG2BHzI7DJAj4
m6ongEDxRW9WUSS/e/Xmgj6GfPtFiBiRI8nxyaW0tZnGpfs3SJqG86lf/EDoG2rkDMGvuyfiq4LD
LTX/ct0ss9BXOcRydNbGOCVeg2b1oqkN9uELbYIYCidNorWIvBttDuxCOc6A00GA5n8k8DoLw59x
6eLnn+mDjW1JpI2PlG7zZ4u4esNdLrO5fhpMNMzvV3KX4ka3DHfPM7RIeVF30hOezsrg1kjz1pL8
ZTtawg/rKWA0utZJvyf1vL0fFMD0ABYxKilRMzLz95dH8jVtrms7PHngBFdzGB67t0gtDBRYrN1X
qVcsGHsI9pu9/Pkng1gUGJzQWIyK9wIaetOGnL35/Zl4+mBzehLTvtG3U5SBnYF4VQBRO5fdurBc
LUR8LXCcCbxq6wZpzji/nzenMN7vh2+HsTWVir6uesCBLQWF1W8Dpn+MpieP7NA65/O43cXA1M+o
p4+kAWHiIQajo7kWuzQK7M3jBlS5sexuBg1X6V3olOCKe+dgaUCzzHgVRlJK9iptG/6fyaFNS2m5
NrKpLeWKs0WvpznBQLZ0DJXfaXYA6T56Ro0ecpPIj/VFyGZpL1eHkGiGFlQnsXjt109kXAI2tfzJ
Kqe9+xkamKUQU9YBnWRNOM0TcOsM0nQuZJqzLlTOPc6xOBnjyjr3ybjkOo28NKU3cenK2mi4mWgL
cphPnxLU6zviULC/p6qo8/iUKwGdO3k3VRiGS4AJ1dePIzDfLYSNn4/kMMPFdzpGDTXP34Ut8sIw
ZMYCo4T+vk4Aj8Sl7IbH2r0ouy3ItP0PQKJyaPYWopiPjisuUKvQbDTvxW6u0Oei32vgdIvM7f1V
OD0RUZ/w63Kk52inL7WWBXLM4DHBm/P3jvz2cG+1IlE/tRoaHT40KSPEiuiyjD/gizcOtTzTf58K
BUC8aDAfnXvNXUU0Vdj5LONLVpKte0fbkJwOwMhk6oDVvo5NycpZyCzlj6rciA/EfmHh9CMBLpJf
ThRfN77pGQgWow56GGcd0PaNdyEIBTT3JczlEfdqRKstOh9OLJ42MgaDvPNLrFUuk7aBntCY04Uf
IMS3/LamCdLc3ArfKK/az5fM/KHqOrPELVCnldSE25KW2J6QSVK6rfc/1coYx8TmGxeyrwN3fba4
qlGBAGU65zFIaBJ9bKTuTQZWquZFaJ+YIDM6eR7oUdWxFZSh3NhFPTcmdQOETs3PUHxKObshnNxU
vtnR2kguYrYUCNaJoOjdxaeKQa6M6UYoc/PdOCYd4fEqqOP18TtOUojhDn/dYjC1gkMCdNVMmAQ+
YdPdzRj1hWJMEen7ynD4XHuaTYcDDI9f4gSvWirYBZ4D2a1MTGO6baaeywPyWb6ihMS2k/iqQPiT
AYKSFTeHgpW+BG9bVLwZFggCPTJYACBV7rFCJMlMc53W62TTY5RkUj8do2EyvP8im6jkaWDttsG3
ooVUP6JfjIkEIHYu7s37sk+IdDhxigzSqHPE1b6ynksVEr2kvdrmhcwAD0YHBnao5L16bq7BKgHd
szSS2V/sI4ll/jXYz24txbdxsZngDAiCo8767xm5extiqoHr7biNUQbmGH2vVOHYmELbvl9Wd26X
g5p//9BgCTMyWkZTujOUlqx1YJEGpOeHv8VZkRCD2KT7EoCdxv2Z2tLJWCQYmyGZdMLmCdejc0PZ
+dU/ebjp2iQkofrQdAv85v9Rkzp4BIoalTTr3aymWCpp8w6qLXepspxZFQhDDLxwbjkcEwHgoSk2
63OTVQCNKvKmDdMKzvzcn6uHsH70/Yf4X4QTKiF7497JBZflAg/KfkThQhVHz76z9OIghkg8Szi1
oafcHEUC+NJ1kcdQ6nw+iX4L2ke7jt2+YxRGfSL1l7kpaE/IChT4zxKBPE5BwsurSi8DzaXoW7gg
996NXzNvnDPLBdkh9hGDV3VW0Wp1ctEUhe4ErQY96YJ9vbUBa11C3SOuHpa7fw6mMb7TyjAXpll0
ApQlARfNU7Nd6e4f6xkqp7aCQPds0DUt821Ki9kVAKTu3uW04LZl0HKOHKeZ5iOLnYD+wImf5lTF
oVQM31MGZ3+xRvOm7VJpePoXvctlXzhnmhI9SSmcI29ku7k9EEGnsE6tFdTPzmQyLSJSyWxk2cMj
gYMWAyTsm3vm44csCjfXrWX9HcHBQASKFy70oxoewuuLyMaTEGE45et+JttTM/r/IcpfvzZB+c87
rWFuOA1jrkOfeAN+XiUNrLLBSxYK2mtbbah2D9hNLExBM+J67+gJpt+mb2jAm6SSrE6FCWeOpmtH
TQmsHrRqM0C1Iv+cAdKU9tqde37QhjGAwaHuMjYoYtSGRNdOqpFdmgm1Zp+A+sYlIhPvN0GdG0UW
5ZVB8cul7WAFawexQjwQtUvXrWDiX1rDTowsWm8Axj7TmapKRk+5G6/KrgwBj1rTMl03qsfq5jae
fzlyi6vsfVGvtwWqytR6AmOUqcBnSWd8dzMuCtVl/KbSLGf3W75651acGYscMHWRq6n1yrjziKum
qU87BGhfwN6PQOgmM2rPf0h1c6x4272rpPKcBZ1GW5D4aTmJxqXn7ndeFITfMHpXEG0kkkm3sxSj
mNCaJoSYOGTtJnud5cDWKOiMHfyBW6clhUo9mSDpyLrCulxvICa0y1sFX3xT04PNE0Hfl0ZGrib2
YbDxTuNIZ79WjuTeX+fEGegkFaLTsYe2zW1U3UgCHXCjUuAtjmmqtKozTGnS9MEuRwhcfwdiQyib
WMxkpK4k4vaRa0rHTM0fFj45nDCSXne7qXD7fCT8c+KKXkkGGqDf4y1o2zqMZGw+oHkyx6oCnC1U
HMzJwKhqqWjoJWPnbnhnXg3UgLS42sh+P3xBCXVaLSsiL8iyJJ7qRJwq53sOlydBt2dcRByo3BBG
BnZ5PHb+/ywySlx0ZkDiFaLB9dx9O6pCIywQmJT03wAdPE5QvLZmOquzA7vRWEWDwrSB4a548R8r
9h31eAtnlJ0jnKjCM8jvOgHi91/Yz9vljn0fLvYX4Ila369bbxbnwS6gTzUJ0FXU82ziLDt7fNrJ
XuvERDx4PKZ9XokRouJV0pAbI9Tkes/BrRsWTue83fgI8YI1ncWkA+xm+6R7PrZd7rmqCuXoeL/e
VnhWzBrhFkMDzTsS0gjmkQb4wliGlY31miBXp2et4f0onGKTzmBNB63NXurUDMt79BJgLrPsdrFB
Pt2Bv4SYyPR626/5fVxImYNyXbLnbCIU4mrW7UoyMpoh62AFy5FD644dNSzNUEldmJpYQwFtm6pP
qLZXNOrD/NpZ/n+L0QdO9eFMp9171EMQtWFDYFJW2U2XUq5KQlVitwuEO9PUj5BHf+/OBa8iPltY
m5wUP4pII0fYENqGD/qfcA3io+SimvaxTcL9uvdKo38=
`protect end_protected
