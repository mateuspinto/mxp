`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 100176)
`protect data_block
5t9A2Qxqsz803eXYe7/PSwvAQRPquncIAe6SM4+be4NhkvJ/cAhUOC7UrMqE/UQdb4wLjrPQ0cM9
d1biaJuKfAYksEPfVF9jI9Ym6SdpPtBGG2PZjDaQ0GjrWnivHEgE1lTjldyQaBdQDbiWrbmhQY2D
MYXUF2lLtn8ABEmU7u7/EIfLNbxLzthlUghkXasfU0fa4IUETZ/ZI4fAqkgJ6to0ylfXE2RfPopG
bXZ3SdgrvwBZDVGnumj+WzI1z0808/KrCZEKC1jBRD08L8/rU4yi1FjoBRCaM0uK2/hO8/8vzqFt
d1teTmqWMg94C/uYGbPddzO818AC87jL+S0/Mt0+NgjlnomaKsS1bY17QPmxCT7B0iL9qj+z7smT
cGhX3P0LqovuUyiOTSTq4gHLbEFQiX3AB9Gb6D+LeM8zU79JjZl6GIN1ds20yxnFfmHfRNgffHdh
kD7THtIaeQ6b07drTOYYTt4da4xgjrIJpHGCAUISt9zrqveC0govXODH6uWcjxOnMrKbynnSpFL/
MEE7oc1Q6925ShGLmhWaFswRv+FAxEuRprm4qNpknHs0HrloXCBnqdnjcJJpj2/W+CHzSOHk/CKC
5nLrYtTiV1uWWGZVodZyb8X9yNiE9mGOcL95hGamRNdIwuD5dwTTlzlGzzdF9AlwMeIkFJtHPY1I
Jm8DJDD+PwdXcBbOGSiM+xUtD2e/saha/Bj8NMdPVJvOFDTa0Yd2um8dhXGzGGNcJAlNnS13i9V6
Jj6WkjjNR1xMKOKgThSbNY6Gs5hOm3iwC0LRUTio++ziG5LBTL232LwsXc6FaHEuB6UKx7mnvhEC
T1+orRxAPYoTiQ8HHdmykZJsPUSOfNd5Rk1obO0LcXU1vQsuMNE5SeXd1Dkir6md7DgajCE+ZSvK
2ZrSBHEzZ6VOhbehgNAlfFTyZMc901+948i1lpW3L77NZbz7JATQCWVrwadJS4G9kqL0Fswg9CVq
5TNh0fm0EkHDm3NEZQoI3FJGP6IUBj/YO7XLAAnfecsLKBMW6uR2CXuLKhj1DezRXhP/IsYv20v9
zoni8INAhKFfzsjxFrgnnHLVdNOByM/vROXFsX2LRU4O3WX1fsIXFGHuqb7NMvQ8KIuGaDUxuF8l
tRGAdKEA9SR5Mkh5dDuCwlpjsjTiuyLIMKhdQMBBZJdSSB0RbfScRyoxz+OGlYm2EREQcNBS6H9l
lVEpsDkjS+GfVocjlhMKab916tj+AKfK2wuQN0AJPxEYRGLhGrA7fwam7G9npkEoj/Bnwd/Ixncp
oMtD4ed8uyUGeIbQg0R1wiN9vwmmw0XQdlIjIHb9B1AMT5UWA+eUwQnkaDwt3Yg2kVSBgUQtDCqd
+qYja3YFu1vo2VALCRte0ydjRyKhnRIGt8nJikSkb83h3WFrh6k/SyV0q2zaAf+e54hYY/L6rraH
Fa8ZuXGbxt34KqZbbHjfS2b9H1y+gR+vTlpVqWqEd3fALMHXBNm3Wjcr9pVpe6Ip56uGallrOy0F
TsBTHthdfdxUyCiakcVHyEMt8wMLoeNFWO2HY4E6JPGZ9LwBqhhsDVP+7Et6lmSjTImiwK5vgG4Y
PzkyEgAgZC0UEIrrEn4QAUP2w2SQ9YYtxOa8pm2cMEdrV+YJMVkkgveFi0B0YlUx7weW6IHu4aU2
AUuOhayMQYCFfwralMeHcaLfpWqVTvVKsYyK8Xwwfxn/QfexdVAp9aCHma3GqW66C08LGjsQ4aeC
icO4cg0eIXwi/tEh9TOhFruiFR/xJIOsb2SX8DBGYXWY/+yZGluKf6OTuvXvqjNOYW+hNXahdX2o
D43fN++o7YmewAM/1tKD38CT9XZmrbhy32DdYwXvzWrDA7pVGFu4m5YnCY0gdDRCKMbaOzcqH2IP
/9yrgg2plmWQ6mzuoXYhGWS97MDjyk4fdZ7bWzI/TgBQg0gEs79aynYd+xLihsM/bTcYX0b40JgA
4ZZWw7S9tHlfhhhNFX2PgX3BihNTwIH3pPE4b6ci6fRpCDS2ZFETh0yJMH+ClRlezchJTSLuHbNF
AWD7XfbzSPW3HfMabyybOZscTvgXKkkQgDiHmIQpmhKVsXGSXw3R8D3YKGJOUtzE3QttolpGmpaX
LupREA6jG8jmWd+aKV7YdkOtu9Z11iK1K6YZfQwGyyBs+yFCyTEc8cS7cs1yV+Xf9WD/D4QKNZgG
2yhPAW7Ao3kxC+O8mhEtvgEk1LlLf7e52sd6mXNWKZZDAW2FR5evCEmZf007sqHoTaFAtOw6LTB+
cJzzBsIop6tBqTIUvlDMLCm+VF6aioGjs39QPg1GIOXf65o+Pqe9OzusA9QTC/pkWQE4+x8LZzLd
SBdRMq4M3+SY4k9/dmmIsSrst8d7mHP98aUEeiefHn404fWq5CnN3HzKPRMOd/Obnl/LbOooCKow
NDQXjLbFN/4fX/PgdGdM8JLq+KyMw720RmzNgXkpXPTpbR9qLNQ/aN2IxGYHqdKRT8UxjDQuHCzF
yxdyv6HNnafW9FpJ3ssAckrMjll2Ypea2xbS4/a067m6+uVSG897gh0yj/lwizcGZlKosKFPdgat
3VaUAcL/fmoLbo3rKfhQ02Ylbr7eLqK1PT3kHfk174EJ3yrnU5dhpuFmxB2NsCwI3EqavrRRliqE
UQapc0kqBOZLIRBdzUA76BU/Mb3pWma8HjvsZJeEcHpWeAdijQtCSqBLKk0XgzdR7+ccxP3g6E6x
t2XEfNcFYOoykd3rsG4/lCqNvt4WRjZ9JrgK4NYSXHhrHQ+ZxXjZ0TEdJEWHsDiINNxjdcci2PgQ
UQa9SgIiJM6/+YQJn9norHy7b43MZHPb6vRf6jrtV9mHQz7lqoxzSIxOeluQEnrb6c6zG9002pqb
I8sUQBnb0oJ45oxWCNRF8uJzpI6ZJcF6bF4CLGF+HciCAUhtQN6oS7oollMNljFPuYCLt4lBloXf
GMGPJKqkwSY4u4S9fC8uIUdY9nmnlQPYiSZZGhhJr2bLHr2T9O5WV1PGxkSSYnHjCsbEVwdHWHys
IXWhcSJEVqd6vpem/+JyU5WnczUd1YFDvEhwGW/HhBTgExQpkBtHWLGu3v1l6l4wBal+y9Jo48Ot
PZxd9CDxEWRNmCUAMhjCSn7CArgI1C4mwGPINSFDsOAWFXeivmwBWZRXKdL3jWT2x/km/r6X8uVF
JK3EnYtXPaEgme78wswzUh+aKup3mbCJ2KLATzz63/eBFEWsPjvrVpd3hoOJ0EGKC3skS7KGvp1N
DoQCAn2SCqhwsHSCG4Z0V0xyQDcn6Ey0icIeeKWLOeQZkOk1nYXOirUJK4yQH1buG7RZluKriUCO
wjXwlCQ+RSD3yj2Qi60eja4wbTDb25NTf9m+Pt/B57MHDFqs7GUy5D9wOg9nfBZAVkcx4+6ijTG3
dHUvPPSJynOsNvTezEZtFKWUN1K5A5IBTJekoXC2KBVGEnP2jGuFMQWdwnSD0d1EGVXN3KUYZsw5
LCzYQBH8W6lCYppuIJRj066FlhVX8XVCyjftpudmUdp4zGWVXsEX9evAW6DWapw2+hK9fuarGHf2
TYZnkFTFLT4+hNJ2pPmxuiBXAGuX9p6TtBNVQncwIcl85wEiirvAdguQ9Flw1idfH4ybMBEpSTX0
YAEsABWymJJzmojupnVGzOmnZB6RrewRu8bi3RbrVc44xYWd0GRYa0uA9l4tZosLH1UIBgfTlHTR
ll/7bZCb3FrinwIMtjzddBi0rOjAna2Ksc7uFPRb96q5zatJbRuasq43GKUnaFMipey24HlfPJP8
IBRBg34kQRb6btdImJE3q1e3Pl8Z0nTQHoiJKvE2UzNHL4gG0YfrHhywzHc3lAMWG11adUxY8iwA
CP3D8orwZWjKDA2RMytkMCquYaiEOmL6QH3efVD+SZCJt9FwPJ9bXvbrVEyCxqydtmjmnW4JiuX6
PKuechYsd+G9BJY8IYBWWkc69pufOGQVSShlsWwTzw0Rjf0ufsVB2Ya/P6OZ1g5mWKMUR5jRfLbm
I4LRO+NzcbFoUI4gbyl7/r+hFcEki5NpNx3wV0XV8U7L/wKvfnpabkLrdL7oFwMQcUhcZcKWT/JZ
w1gWVEPwC6/0AsCQf0gAGMs5hd1d8laWQOC9kEDf2adF/ist6gzzytjAEzS3+Of+43LuVI+mj0l4
gM05KbFf41AJBQ+5QAFCuICOmr/Am8khh9421ryJ6rBpJPdPYrnN5i2FMk7aE/NpiAyhkh6n4F9I
obmvgZn1pxzA4L7dnij7bH40zVA9yd8+gAdRxXGuu0rwx27h69jaYCx/qLluW5ukbjmfY+l1BQJa
XOnXUluTNQGGUSUVjmJ/UK/GaNAIUpoM5cFEZ4S7Cew6vwKjMmUk9f/wPWk/KifJZ2pXOq37Sr5F
fL+M3wQG9f86j6oQEWBbf5Qw6pIJUTQGIeJuX2ckg976+pzpChBoqywQoiqRStLGZxhljzZG+DsD
+MPBwo6EaL0xZYhk1t0apvxBySh7XDQPObgXHTUs4DJiuMt2wBZHFbkHYuwIPf9Jsl2OuEZ5RPtL
1ZIEJA9crkyIaOkJBs97PJFhN2bS4LPZ2YqaQ3zLzl5O4xNvXU1wfTyoqe5G7tczXYzCL2J84BZe
sJQgTkxwaF3YeXxd/oqa7mMFI8SS14+YbkD/R+0SZfwfhSLIH3lknuA8DUdgMGHrX8D2OhQ/5NyS
cNaKdTExyCnNz9zf8Fu/BAB6HyVZefRLCJzuRSQZcU5/21k6Q8qN58WPki7gFyYwsJcVKGWOC4FC
hwtzpzXsqpKhneIPkAJIXf8kC3bC4uB5pP95sQfr+2BKHj7re/vFHySfzYRb3860gfTh/pbDvyRo
+EYExhT+6w/k5qps4qz/3vWpBFSkOXJ7Yo6cOC+v4dup0LT2yrh5AJH39vywAsS7kX1aSqP7tFVF
oA91l2QpLfUqE/RfihmM8GRcPP6fIMAm8JW7iG6o497z7Nhn5AJSQr+Pq7fya5Wllu+TwTLEdKXu
BQmAJzivj47qlBnRH0/oBlM1sCuEOLsXofKm+VZj7iezSRePkTw9KNlQ2OoMggXmT5CSDRRBSPeZ
0rXDSo2YS4MvBVN29sma/RVNWvj5rhgJ5icAvK8PNdciBXEiwo5LrijRR8JPqLzyjyskBnyK8uQB
5SHY5z9BDese4mPr4RwJq9Tjs9SX7uZzearu9KiwQaAHTp4o1WogP3i9Klj+7iMUXeQDxxGWiB2m
GQ1NWZ/4tdZxNQYPZTGi8EHFiI8wshTdd9uw+EQLeW9cf03XvetoOVfT47bmm3yMrPizvHgxzFgg
19/69/q6KnvrwO7bOWxG66UMNbiQxh5HxPkj4VRyqUf8nsyKIuNwGptn0bCJRyw5GNpKEjRRQqcb
0wHpgkduf+/ykSg2wAGefNTIg1gYYDw9ifsV2U/6r9Ss58NaJf7XQzljaPUNKOu6YYgYi57fFb24
ant5zeczDBQkHQG4wmLAMc/oRoqbMyyruwPJhWiA8m5oO1mlL2SiC4j2IZnf2KCHuJCEiJY3ahUD
mKi3mt8Vq8mwNvMCs1eCLrSiqGzMBVNY7JJbFuU/tNl8Oj+SdDLldAYqqv7GwtJd0kcJ/M0ScZYE
3P0Zpri2ULR5KWqlFq4HH/s7Sk6LIAvhZnMYlU+b+e8IwqsMXz7mgqm8jNsYAQWrsxQTCqtYfaPv
2ntIJcK5aqKcQUQK5wRbff572GKjay8YSnfRmTFURWi4KFAFYKT6SvC0zDhP9pPW8WHdk/hpP+H7
nOQOAA2n54mYzqb+b7LdXaqcJ1vov2ZJH9n8b486jAFx7cRaEixyq9robxQPiqWIwsBnmiWp//PE
odtkkRYgVKf2/qJXc7J/F4mb1tv7tTTNTY5X5iShPs6DBr04SGNM2yJYDMcrNctGqLemD22A8yzt
WbwfFDwPs8RnL5pCqxCikgIEoLgBco7OUXW4zMd5G7WMJS23u3Z9Dewz9Mb9aJwjz+rKeDNO5P4v
A/aqo1CoeDxcTas0zhpgQw1mW7cc0yI2mwyMrGF985I8ieRg2eWDW83O1qv4WINbUbH81oWwIHns
/E6SdPs7Ya/l2OrO2OiwxR1J7LH4/66/ZY89Z3Nb8BCw4UHoKbjjnAuNobuf56o9aITuP947CsI1
t7cxfDeIT+Vqogo65/kEgLVUhsT5DuvRousV2coPWWHSMFS607Ex3MR32pY5DGEHEAdzJKeFzROf
uXjnK+tmgNHM1DzxjGfxL/7AMc3gZGXRbhZ6DYRJy3cMnggH+4w9Msv7hEW2yqZW0Um++POgczsP
YYQVWPUrqzAWF7m6So1zOGEPnjZXzm56pQP/a7+JmOcpFkWeh/AophvsFOJGYUxWvS+4SRzoYgde
oey49Yw/jjPda+kOhGQl8SzRszp6W/DRzkP+gHtGKBQxOA70edJzvfM8ThGSFzarUMshNIFqgQvK
vz/Y6qB0M4Hhe6NJZRoS5dp5kZFS4upfDJkARDK3NDY63Fpd+4HzBqBB/6cz3CV5lP0CE0HMJ/ug
C97oXND6aIM86htH+6f7gkPpP9+KfFsA7ODvkG3GE6KkNvskgfkJBDCMuwG6RMVHf7TzUmGDjtQk
kybdclkSoKrjpvlsgCyiDOQ1vsPcdhm9mQkjCsg9QD/HxlGAC3olcP+pVTUDBf6Xicqp86JUnss2
RE+rm0CFWx8DsKkYzFxvy1OdFT5CP+IT9rZ/EktQYLDH1FHh9fD4/iIjmt7orpGjfxizMMp68oNH
qFyaVLlWKo1eG3IMV3CMKUNBlTxyJXRPOjhKAW2ibkY1CB9jQWe8avPEzaKiQM1LyVaqTblmdAO5
AzmC1MRvK8MvrLaoopbSsHIjEFEpKUd6eILIHtWah6CxZowJajp1q7LhZwN7RPNhwXzwyaG+JKxZ
/VwSsqSG8ZtdmMMc4iHZDUTRvN4kVAPPVd7N9FOEPE4rfq766XZOegJe6SIJloi5RIDu+rHc4/7N
+/+i26hN9l5KrpR5O98QKxdPBsYuy+qZ8xJdON8lhEmcMhsyhFKOFcoZFb3FI+4NkPdWf+Mc63Ek
e/DubDDySkMg2x7HXXkJMH+6ahPcgoH/HOP0JH5QxHPKdmmcS2T2mfvVb4sGQllbwdnXOEPT+ruk
qHZH3rV3Vx0Hzgh047l+8ftzmHTuBXsf9hWDtusTDZfTSePw/jJARLj4Iv284pZcCVe63PInQEyg
NNWUbg7MWDkokjzl5Hs1ros1K0vroQUXwq+GwdaG9Y1Ywgaooq2aCB2Fn0A1+qy4w67PTvYQ+mib
ToOnRfzkCY8uUApQpnkRGn0UxoRDxDltqBbP8NPNcBMohIHcTF1hOXYdN8o1scwsJCZ3tFt+iYC5
rMy+DYp6WB4OlE33gpI25jP/Ut2x6TSniATZQxXSEDt0r5/fzRCsvuGGnlhuGsf0PfyIbxwEAzsA
ANovbzau9534xX9EnmVsxBhBoGVmAxIn4favVuCfuvRsF3qt5i2foT4k38q4Tntpv+eV1N7RISJ8
mXAI0qWcR2bmnIjvFQLtAkyCmWBp3QbNw2w4Qtsx+ROf6gixveuCOPDeADIq6cS9+8Lkz4gXuSYc
tylcZFzVkP5krTZieJdE5bG55C/VUCGg0jDivWi7gpxUK0PXEw8Genfb1Xqw9F8BxnSnC7t/I0x1
u+Lk8hn49/FemDctHN7hTPolP8Ybem6z9UvzcfnOwE6B67WduRJoqZdxI+dO/XLJM6CmDzrgsFDC
nTvPFlhPXa0eSE6sKq0tPJsrZjzhBJEk0ZV07iub/PG4u6/9zsyrmAtfm8kmMN0mJHKUCleWVtHH
odpeIUkAt1S17Tlpipq2qs8IUjAyQHF6EKU0q1yZUoTFJNd/8fCPkMp4X1vY3HPy/HBbVj9Uv7SR
f37TZaF6bY1b4Qmy7qnj6480TtDCwOW8jDSO4qjYK9uv6Ni384Oy+mLlwKcvDOV/Xs/rsAnMFZR4
HnhMCQdrBkdAMHQpeF3h/Ibp0BGVkXUcmN5Sg5ccLhRdRL+dGOZFFcKBUucRwzGpSXLiY8fBHBCN
ByHR8xkgpK0hvaRYhYtsxqdepOxGuMKLMf6mV816Dhri9rKkxCJfU4w81z2GLJo90NWHkx9ExRmS
yTOBudb/Ggz5IRbokpk4gs771yba0R5nJU47J+zF9n7SxoqbkLdObfcaLPINlUYrcr5ciYVJaDBJ
U+yJabkNhTla+xPW8Cpd/r3eHiP1tQzRNtPWtKb38+hvGAYZATK4e//bfk0kAyLU8WHbQTn15TbC
01hE48IcRRVgvj0fsTvHI0owNFwlVggiu9TpVsHuG8e6q/8CuSW9Hs+nzWzQXjWVQxElDpqtRMB4
wOX8NrudtF9a14acrfw+1hwJLXz0J54KB9B7TUrPr4gKnTj5oofmQI3JishwOi7xpERo06UQmtxx
xCPo33poYPEBPUM5dqT+gVouo6SeQ0nymfQPCp5m/ixV0zUjDXkYohNFoiRM6kLihjuPKZmbS5id
eLSAZ1iw0TzMuURnCXEVKoduKiMirCgNtSE/PotBAmhM2CLmgoPdNc5USXDz/NCLfsPZABof6CNl
0I0jJXOwHMH7YaPpgH9DgS5fTrCsSYaVzJw8rxOTckNiW6PpFSeXFvE8Jgifhvz1AL63FcYLroKR
YdRFtFuMxQkrACUuz1+l0B9AZL0aOhmSTFGHucIU4D0WbxhLp1Hkl1hk3UJkzlji6uteXrAguii3
q2FUAPj4Q9HOg5TzrvH5VASlXqMRCud+wDEyvICNdlhMBnaLHYf4A3/7ndBuUoIFIKNszkOHUI1z
WTRPwMpkSc6rs3lpPDQeoGrc1Nv7TXthBvxFASzbfrQdVwx9cNXo6Tb550/Ca7KLMEiIXaY3RUyM
x5nK+Mch69ehsYnwPc+wsQHWvxG5zsb0SUeihVoxvTyZrwWGec+Qy/nV5D5IJHfFOraogrrZeKKr
trDEwO1E4t78lfnAL6X+xFsVUGfG69sVjdUJQJ++pt4Gy7lmhXmgRzcjrR8mcYrvD9PBzcNm5Gb3
fMHJN0vAEEy0REESqbKyKgdM4D1ahvjVKV5t2/CjzrQl/YMFm41bgrPTxX77PxbyywYNEyZswRHW
wc16zY021DSx5fV2L0c4FeTeclXUaQPHIbChl5WwV4Ygc0gAv8gEfgvxzd3NHxSmM//uZeAVxkup
7GoqoRSRDv+M/9dWF94Fsz7u2G81akFUJBMpLbKyiVyJDTEW2Bal1u3tclBPgq8isBXu1YRyNsYe
kzy2DlDg3LKP7bWL/jt3FT6Vpgzvk0Jpn6EElX4hFbQOGaYI5NHZZLeDnQh4VMCtV07lqEAP7Ii8
EzE4WR+uOhyvQUZtTtovq23FVzqL6LeADCbAMi2jb6SFGvvSlDm9ZqoBwCnQgeSOsvjzwVnAXLO7
N/CbQRj/egTz3k2iM1VxJ8k2stt7t30ABuZcy3EXhAy1I5uHdLdvYx/mTH1O1oST9oeoicE+4t1m
jiTo/tQugh33Z19Jl+PTJqcDaVvYsZTehcIpQk6RiGuD1f1VOxcIYkaRuIAwwa6IqTFO1lXptiuz
lFqFipRvvLbpYBM+1GxL9zxhddKoFyGTMoVKQJ+GcCy7gLX1ZYbYO77utBdJVXJqd/J7BPqrcqs4
Vbr+GFFK6flbQah+RAD79K0dhZ7lLRXCQ4VkS5ywmyFGVSUUrYJkpLXmJyCvFLS7eqi0jkTuKKIS
SVz0baqdfhCU7lxuqS5J2agJYQq4eKM36t29XKyeaDpV2eUZPpV14pin4V7l0bv3N5bNPITo0YtE
t9IDkOhEorfn0o8z7Jfzd/UwgWaZw1ZPfYLwcPHPWvjjkgvKUWMRAfRKFM+J67B+Pwg0De7C7FdX
3p5vDgIn61QkH6zp1KdVjJ9IeiZVGS7dZz/LY5BfqsKic0OQfi4ZviZBHdfAvM19Xe9uIMV9GCd3
0DvqfbBsEt1bMcm9NVBvnJIOzBr0EJbejcQaYNyGwfe2wXDi6H46H2miOa9u6Wby6L2nZOvhTBKg
GfRrRbAk0YY53hC3l02WRaooO5AKTF+wxCaZP8tmbmLKfIC1vMQWS+FnGwucsowr2y/epQCnY9ua
7WVnd4Bl7a5qWfsNzTYLBPdNoWVN79OddkepZn4C3yOs+8ELp8nArwL+BToGlX1sKMYztHvlWmFY
cg5qquNgLTNL0UMC1DOhG5L89/14XfcgVprT3GMgrLapZh+V+Ksup3z5dXNjUpMgbmQEMcP0OLAo
4DP2W8qZbaQmo0DHRnWRsRea/HbYjPzIpRfSlly5ZOoGzh3AN9Dn3jls3eyQenSoXYy0Jm1q5NUe
kY2wqDBuDOUIfu6zY2heNlZcXb/vbVDHtZeiiZnTM+rkb/M9XTkkOdGD7NAOsKU7IS24mwFsQ3Hm
D984Uu9bKvgczfxZZ+RODuX23k3Bqwk9of3qUYseW/qSMkrpqfzf2up+0yFqhCTHvlfbeSSwSHty
l/e+n01TrKs8Wm30AeN32p0E/cHf1EQNnlncIRaHoxk8TvMr7jl459pYW0TRXP8i6MYLv1mcXE1o
4zUOqI9YjqkkO3WfB2YyYfqwJry7A7B50YyEvXwm2osiupxZYjBmBSt3zFnBvWJhsfiYH/BDrn/N
Y7Z6NIYv2hEG/p5tr96L6/kTwthrpEsz/Z9klYr1hGn3qP7ay/jCCiAMyPy72lywCO9irn4agW/M
6dY42pXUlKXzwYcKpgnfPdkmL9uX0yOYlfSrapOLQ4oI+SrgGokguZFFoGU0IGnh3IUaXuKELnuu
bB/JbwwRtxXzo5LtTXqxwEFFm1T0+JsXOg/3lbMhJ6qdvHX14ago7kxsbKXjjH5vkO2SNq1RpxXP
X9IlCWqRWuXYcZvKnYB5zn6s6ao0RZwYFz7kxqOjZGlB3MmDCVXl5wCHs7Y4nHLAczSNdL7MZif6
xgpj33ZorzSHnDU0I11pzFPyVlD0OjDhotWwP79kAkHLHlusy3M5FjI7Y7cDd45JmIwxKyrFy7ad
qIWpg7JZ5wvdfGgV0kc3FYbuvccAs14Gik31MEipu55f28+vGMg/5tfSh2CENZ0sYOlueWTTKt15
GKV6PTiEOJYDVgJ1KAhlIJ3e0+TQf0PhY8Nz06cnks7+FbOlh4ucXgNWwUrtahstesu3Qt1JzQTZ
DGaOGVJW/ihHP8JTC1oV/wPNTRy6KXDZzeR2n3TArUN/M4KNTmTYanpEolLNDgMDRSuvySbwWLJw
Q7Dr/fcbyOn4KKKK6JWjAv6VshroauiCl9yvBbzFRSYrI7HD31sYfITS+VJYbzvuLVmawJxjif1h
8ejQB9fR3iRDiHPhtj6kHIPv5dM6BrpLIMmZfyZuo0nHGwgwcreypUQaNBWXsD1jzCMWaeSWLWL+
A7TMncCPV4A0/dbtMZT3+r9NltZhJSl0lwyWZ/G4wEv2mSmlKsaJM5R7oCPvq1THVzkPBGuv9U/U
MY2w51Rlc37+jTsHQoWhzaZwVz/VKqiM34zHyR+dPHLzYI+wYPF3DaPit6zi6sB8Hh0D+9DRkmTp
CyRTa6xHdlAnENQWlg4hb/lY7/lJI/4QCP40jmiMiK7CFlTDR+OkAdljPD2VUMwvsrxcBcyC9OVS
dgogfFLjLrTNewBIp9/MfIk+VlGz3+pyo6t/A7UYV1AvvxZrwzH+TKN1Udrk/ytrkzOTkPWEVy0o
rhKIxqDW1TDaR5QJM73JS+o/6gtamtacVw8VQTWd4YvfLjeYQWInnNZyrNqaKLUbOUsowKuK811S
eYQtaUpO1Yum/BQqMe3IN2B/3sRsvPTXdbnVX/HmyNk6aRBZiQGrzQLhqBZ+9UwsHS7eEbRHEI0g
GalSSm1gHYABfwUjTX5csKXyx4TPA3coiSrw+e8jFH3Sl+UycKKCB/cjBGH6PayyTVzXkFmK+PKN
9FY3CTDi0x2NKM+LwX5bUGM+QJzDU52HU/fa+JNhpi90CPlD/5/igRiizsRMMJ2PFIaeLmNzEVhe
YDnTgCwuRm6Q9ErRFQmfmoJiM62kbBzsjR00LNwvnqAQP/8WzMw42uWMuCcWLmyka1HxQx4nz5AV
b1rw980jCfR4LUplV3vFpamsLVfY0lfwN9S2Y6v1vRe/zBg3Il/ZV9fLZDKzXAtLT1dcP+57ymi9
k91hnO4+ph4i3hUiOegX8zSoXtmDDEPSQNpxbI/EISCZkQSQM36EFMjLnYQzbGaGytYibN7wmUDf
uD4+D82iMW8aoY0Mhlxzbvf7F5C9uHEp58FX/Ti80VSOy2o5MdcDwy44mcvG1K/C/R/WgVe+pG5h
/9N4EQBv4eloZLqyiEGiSVC/YOGVXrEqym3xiGx3P5YFQ6K3xdX8lvuyDb3r5w65hIlAzyL7iEyM
YdW132r4GowOwUiTp//SzwVtq77OZkm99jFyr/cu05UTfxnVmMchI1xJkMjD1+Al2jhB5gx3GBPD
kOHpJKMt3fX7Sxo/gRxT0GTzIgca7CI7HNIxiPUfSYN/vWRek9B3eIA9kbBaFrhKTROMMA+QDBCo
5ui/d4ok2s3ukkTP2kLREnwBYNJ8YOp2FWiY+qbBYwdRG69CLzpDRBGZxi6Bh+tOHOMnI9yBcJ6q
lPMi3r2yVXg40d9ai9kKtmyItPvZ65Gd7YjTld37uZuEmQY8Yl59S7G3YVuE9kfFgOLw/w+QpZyK
WYrtLVMfjBK+Q/jbtYnDh9rrCplYWpPNGZDzRW+vAfLB6UFOmqujlOpW0LC4D4DTa+J9Ux6ErGP5
YzfQonBBgaZrdANppdao/QN78GxQ81aXoAYWMtWgZVu6oTdg6TO9Ql3t0nmEpCLMPGYEaYeUbbtr
LKrGgb4quj158fG8OiGovYPotNP+S9JvuAcWXcdfACAH09eiSnHIOeXjaB2ERA+uTXsyLWbbfbHT
CG+lCClB4ypgIq99WAy4odS4PyZxtMRtUlyJ7q79Bh/TSRSCGIK2QrmXMCTeO1yAhhAWco6VNLfw
AStxhGlmRyvIgSHYHo5HpRAD152f6Ud28aIo7pH6M1higVgzoywhs8nnUsJJ201rvAbuR7ZCmqoz
6RpK/VbpTwOFkU6r5Pe9Td9NsU7iixFLqXxVB7sqq8dZ8PnfyiToakhaZfr8WwURp5OGecTMEarT
NdvaVkx3O42JNdTSPmKlzHSgFyHBPBvXtNnCsftmjdp7nuvfwgxI3/QVKfyhPWx7uI365OCjav8G
bJ1RzYnoymiAKOnBmWU1XJOcn+CkB/snQg71a0gZKz/lETCQqJliavAtaw8eCU7HohzFp6FgmZ/d
ItW4Bo7iDs77OBA+FnlBTIFRoZTD1LBjRt7R4lPLQoP1gIopu0qTrheQp4Wrq33xks4IWtU5qf98
ovZVWn1ihss6Q8y9Dp3ScKO2/dY8oYu5CFHa5CsGfN5mPDTwMDe/gJooMHmBZgWHsU/xqfB1a+Hi
IMpo+KzhaDYekF4OKDUJuuyHONf08WUSqEd469ibjHo5kI2YEPK/IY9e3jXM/3Gr9+TtA+FJuFNa
bFoQCzh/KwN4S4CcoMjP7Ntn57YuIbJhF+UcTPozvYgEG0FyAEERoymXcJ6Qz0fkxZcFCLmN+704
e8rJ4sARn4f5VzdNXrcW83vTPjgj8YN5OevBrBf9hLZ94lZiuN8eSxp6CLaMJ0Cmyd+SbTYedc37
Dg/wlSxaBgjOlDyz5hMyOCQg4Zr6/Z/m+YroQeUCnFsrX9Zqvo7BvjuOFx9NtvilquiI0GFbranm
3mWZeBjmKrkW/2zbeSeQt2AbUybmfmELyafc/jXSwtsDrMQdcEDpVIdZ4DLDPWOD80YzHVlwGz8m
67kVdzve3GxXq3Ku2XP22T1UFSd7IFIt+tNNHvguMfRcLae2nCS3W3fac7xs4cLGJAEr9Ee1r4b3
IBKE9zKWN0lOVWFiSW9pi0wuO7ATO5Kw2Q6PcO+a88U+QfoAZD1EvmOCj4b38ZecEinjOZP77aWb
erTXl//P5O2cIl9F+bzsaR8to7aNaHz2WkYFE6L62DFX+GMi59sM68sbii1Csc4RDQmo+gc8svqu
OmUcoblJRkZDCvZRJD0WDer3w6Eh9190aAvzNcj2jmLzHQ8X1LNae2dr2i9bl14pmQrDB/UdR/d5
BQxCIUY5lIdo9ACt12DyN72CL/ZkQ7y15A3ptslyJdTomQ9q/yD3QjVy3UCaZGlt3s5A6keDwEJg
B9DLNOQ/761g8qa4q9TRgOoMXBg3uURbAn/kPjgUMKTQ4J1DxgEfq0lqUhCbFR63cs6x3tSThXkG
c8TSYCnqtqD2zFtLxir5dDaYXycRA8s6NDXsWK1AKvtcTPZDWEcTpTBzZJdZrr1IaI4qOar6jyM5
Eg9P8fWpdDxZgSoMD9SnPtRvLc3pABzO+sQyQtOF2V2hg3euNh8xD7wkDfVBJEakJnZ6HZlGDxr1
F6FGTqCrD9wYYTrFvy8nvud70xIh3dIctiLeW6EotZRLSHZlF8i4weAlWnMYZsDcwYalKc8hyXee
S7gbtnKNtLRK9ueKuOw+rdHr52gVMb+PXLWh6fVwuApz1EKcFwKcyTNkY986KL89WkuF1BRx7Xei
X0qyCeLjokDkrbJ558iKdiKkrXZLMZ9oZIUgyjnwsBWIlhM1DjXJ/yEADnMXmngNLxDp6kRXRUl9
j8O7ljyX/QFt+ZwadUd1DK8ruHCPv9i5zV+5GZJZ1xTMVHFlQm6PfC7Q+cSQ9p+NAoA1I9vHFI9W
23j3+4TmU+1ZmWaHT5PP7Lj5xuSFtRRf8sSuNekGXPp2tHLZm7bd+UOA0lFFYTJlJTbDwkkt3vKY
TzbSmrddO8y64j7r7lEifYBXHexxBA82aDz2/InvxTIJ520eJNPVE6q/RHuKJb7KHHsHHwD3WIJR
74b0nQ9OoiDsxmhcvBTuFRSdvjJxyEzqx9tAkXFVmtBSjM7wd5hkcK5cmlh+gt6UQ3sHVsDfRNFm
uslIfbvJXg8JylQc/ecBtzRLLEqrEKX2TMLygY7lTHCSZHfLepfJG4riR1D94WL/Z2Yq3lMF2MOR
J8EtV4YRzdomsRcKmKv0TDfnDO9+En8qGk/2Uh2VF1ZyUfC6U6OOM9WdjohIvQqvawA3I4dRG0r3
2veVerD+M6bOYs7wr12V08k7u1OyxgYXXOP9MUH+oRAacbpEahYIkBWoTDJ/DNlmx8GgrcfZjwZ1
7p6EkGsAWQfArzC7CH/E67YGcEsISQzuTLLNWeS6YfN0XIbB/OXEMvJ3nafRfgok4Ke8aBtXD+dG
uhTa6d6FC70VJumYk1bwOlwQNER7ibmqqj02UkoIkH0q354pbZ3GWQRMhurfwVvmL8b+zTHFADqW
5ur5vhpUZLCZp28OZHQxIqmpRpM/AcjqOAHD6rbpUquZgSG5POXGhOx0Zev6tA1Jxsqoydl5muSC
/2SE6rbxza+zE3enn1U4LwPXPKMGUQM65JlznaM0Fx7okphWcHYzfh42sL8jfr3kCRpyTXkuv+e8
WS0prtHnIyW0ix1qquq3qHbRG0cV/fKjLrtkUWyJVZLKOT6Ly5qfxyy2WscKkVMaQcbsyDlzM8dK
3lW6sTk6G1+TbaU29VLUWsgn9qH7NsJ4jW4iPrmx24gwXaKM4uNeHkLfubfYDSkyrP4+LmPgeEfF
cgGjbxrkrBA1GKnrHzisshQwUdtIH5H++U6ZieLxAzZE4rGDlV5tg/7m6D9ChfrwUPMb/bBPdx2h
oPte60JAX3e0NVXiouWeVq+fNde2MT7Co0Q9L6W776iSgXjz7EJ8E6EsaHYXRQ2xjEukYLZdRiNk
eIdHVgeyfC3YKhXmUwUckFCxL04nEjO0PfxqAWdT0y0ugAAM/D+huIYQ1AF5kZUpxaVr+kLiVmbE
xFncbTs6y72iER3I1gvUtK6eUF5I9fFtrOcEmPOcDkJ6SrqAQw/1geE8sp2+eJNcGovZzt+Gqq+B
yZwegRv1Jswb7EOUS77N7T4FejTG1fiNqdHXYKjF50b4aHP9LHMWbStXJFWyjiy+5b62Rx+zDBOP
Zucm1SYbX7Z8ujuuTKQlaSJ+yYabbpRfDxjOcZGaDO0/ary0zSyXBntBK+cBZ7Vn0DaChqJRdvrG
tnQWSTjQpEFasQEk7NmJ1r4R1Opbz5cIoIltKkVcYK4FwwDGE3CktGBI5tGG5TX2vvPkezIEKomI
kDRX6ZSj7ubL1wJ7MNHNffJdRrOFIRR4HqYJW+DoCQsTGrSs9Zg6XaC8DVAgtaoPgC9F7OLAdEUD
6gGG6fDolXAWTfCDu5X7xzHWCpmgIKfMCy92zpOu98YuWlJbml3b4FEZqsZ3AwyXCjVYHtHASC9l
aMeRTvHODGLBUR0LPJx4Nx03wo8f83jxx4CT7AYvuYSs8TRFhJYt2ikVgGhJqwg3NlPNHjcI8Nd2
xi/LAQsYqIhr327BVzihsAO8a7cNWgj8rhjhnnUfdjh09omRrF+sUVx4ZR2hfffQRVkpf95W00bT
XXal83OBdL1my7VAsMSWULaxBtrYVTqO6G4tb4YRvs8boj//BY5XiPAcQ5Yvmn+0kXEOWdFsZqxz
OncMVfUgXitsrafWbUTMt1Ke8BK7tRsiEB2TAIBWOUXXquevDmTuHwq8a34YjvKqX7fcVxc075Lk
SkCcChNVtg8SSru8bkVi/ABsbAdFB9YhpIVFdXNxkEpP3hbuzMi60PABvv7+4RrHhGXLoyndBgqJ
C0tvSJkFtSDRkVzF4sf3xw17zy8mR9cEnFu35nv9xS9BCyYJ6AZSRvwUa5vGH/+N9KuRm+yPDMG1
/MGYDmi94HlpjFrPvqmNBaO+KlIQ7UNdeVAd0dRzPbvP572mVUlwI7o674STjR8Qe/wspH+KoFyb
nzVwyYPYfX7P2Nz7LMu4K6Awx/LogBqw9zyG4z5vk9DXUdNmQt9MzTBMC1CzkPsT1pUq8+7GYEPS
DQspThWNtAS/EdY4aaKsboyKrpp2OWS9CO7vKx8pc6Gwi6WXLboUOM5w0RwTezbrMqG0K+S072LH
Gaw7hZ0LApcJs8LiyWD12WSM89FYGkVcGYpHMRvdIF+UgXNxAGfmqRIjVSYLUvleHoQSzGt3+UQB
BfBanQcdNSopsjQSFtUTpdHVgZ6gvPVyJjc/Zqeu/efeoD8Zx6mOXp4+1Rr0bmxMrmsTdvCiY8bu
sZ2WyrQrqRVwod6aw1lCtzWhNSceg1pyepZJP889LaRYBy83iho755ox20vVbtbtVZ/etCen56i0
OT4k8omgeEywsT5Yv1MRFU5xa0KVFPXqb5+vTx5HIVZdMANix/PnapschCeUGFtWbZYxh5/QKOwq
1KA6XR79biegbKFl1vhkdBEeBR5REGRK4ilnwMEqRSihBPmMbcrIomsanhx1S8SwbQ4uS58R/jdG
rzt8dEIdNtTSwzX2ZDtIoo3X03EXtGlKNHTyw5eM/U/9aujxBrrjYUO+K8CVcvmX3uB01Gc/QTrH
JWB7IccBhvjXYIJFuVNm9R88qaGz3uCij85+aEFp1WPJdOK6+80OZi8ou/g6KyiuwEAwB0RILYwF
ge/Vopjk0Mxkwmhi1oXFooSmSCsWoKnZjXp8++w9fRvtr2jK5ZxdfMT2qyOOfMWEZRXQYDIDvr78
oqzSXOvE214Vk47CBe9bPxTRaYFpF8K8XtYCRME4iMyQ4kCzZSCIETN7lKUQZ606SEweAlYlbvxr
8lULOjegQifKE/+RmPicCrnZJMVBsJeatTJV29+VGMTzhpIEumBs/FNFUlHd0/mvSg4Rxid9bHSl
7Bn5yd5AzcKIarOW35/l21kXl6Bb+Tc9o4G0VBW1SR2yfRyIm9bryECYbVKiv5vKtFG75J2neU+w
acLB8DGyh0MXZK7k4fZqgsK3N2NTtqjOJuyfKJ2SeKLpur96lMz27RmKyYIdMhRIpVSp+c36NGP/
kl3duN72qfka61W/iUEd9BbYCtYCOkvxmb1OrG+seb45yz0ziA+DEexLDlWCg+D4VNY4Z813GKZv
CSoG2mUr3Pzz5RHWGm1X0R2silN4twLH7/njV47zmjzbv6Ba/xL6Oqw79SILVM24CTecrY8dpigX
jFHpYsCsMhY9yioT9A55jy5m/fkoYxUCC/aTN+UrnkfCuJNrLZ/hoLSTzl2xdPal8kyDVeWmwLha
RvSStlnbg+4/wh//Pzgyp2T1NRN2P6dVZjj2BJbiDWbaB8MQve7UN4qpA0gr1+2+FMICqdTHiGO0
MXM+nUZc2eynPQxUJjVa+COptCoxmuWV9W7oCkgELGf/IZ8nOYh4H+t2egvNoJs4Y9ha4nBNes3J
Qw2tumBUqoxLg+8ITZ//UaH3861SGBYCFkMmg5hNkV/JKjyHYY3Ak2M28qNH6o6MRsdMsTOsIxlG
iMp3VUm7DCSv6CM1/UUDdx6RQT0WrKeJuzUW9mmOwZiEV/NxTDKcmVqPfHApKnd32Vy9mcftTZ3k
826lodZdYLDcsmbKDvsrcF0AazhafpdEklcAaEBji92/eFOtygeFKDAhCutF7Q8DqlXWeDgwuK9d
CtMnU3lhkdeoWYaWknnnjmtPLkbsknvYMyjN5UUgdY185ciBTuzk4ynS3AstrgJsO2/GisHo+oIP
Hflc21tfJqTHzFwpMh0BBmqU1Iez50K40xKRgWX+jWHMktX32exOWcjZ3DtGgkaLZw1ehN1ss5Jz
hJAQTY2Yt0otCqLr0LGurzml9e5Y9nTfTV7Jh6oN7K1ekW+qzEYZQMWCDjLigJpb4kymscAwF+Fa
XM4WNm2SZoumUqG5sm3rhZOCl0EUh7f2egeZ4c+qida79YRHygxVI2yYrZaDkACeJ2dX5FSpTpJd
BEBTCoiNlDia1X8vEocKXCEznxWcg5f+opHTApYoAOfazDlkOH30ZyEnmYhrfNta7oc7so1dHlUU
3p6x/ar70pOTBljDc1PVD5ALwb6gM6h/U/DLMC9BvO39ETaCvdkLTR8O8KGrsMYULYIeGyXXPrvs
tZtzJlk4PCnvj633d4sRSTL2ljHJ/maEg5xTEM78mHXuCqeuZpSh8RpmQ9svBlBRvGEwYnehuvAX
R91XuvoOhC92Sr6H5lOIPul/OT3ktmkzafMhKVUOsisFjLGt1m9Q23odArOhp1oSxf3AM4FKrv/G
31o40dvRO4L+EybKrCqJbK73K7VlUwOypVLSUnE8r+Oeaf4mF/tyTcSxh0Kyuqmyk7iCAkxmCaeB
rxA7MnpHxJFArhbflVqiDX13FiijgTg3H0x9uR2VMjmDO0GAl4aAh8kDTRpOKPEDVTZ6qLk8LQkf
75ovCa5CaFCeeNvrUEblGhtCeBs16KeFnSPMTdAMCTQ6VjaNjoZggc66D/g0A2urE9jS/6iadKkc
Hj1AWK0qRP+iPpBEEBmajUfpvPcw2G96GH0EsCDw/+nUzl2MCxGZSD85o+BD7OwY6Qr9xo9v4hZT
UPjj3BMqgv55ix3MeshFtxAKd1v3VdzE4PcNAKbS4GdPAoqq993GfhlH7el7lHWV7cUUPAMG7ZRk
xYTqE9E7ajKe7zBewpmwwHsPSaRqRhy5Yu+rXVPNXVd/+7w/9QbwWeUE+Jyzkm9u2fYJta26eXp9
AweSPTdT9iwNeigl0f8iDx6XIQNZeTCEnPWVRB8jPJrzSNg/QGYPnGc2SU2hEnhJCHHlLRA8W53J
yAFIPYCESn919GNVHUlvqY7y6PSt8RBDv07wzJx9fGR8xJ0HWCsG+42zoE3KK3c75G8e80JK+QVu
nitPnaTzMNk22A/6zzgSiNu2a9RP9yjhrtV+iw1faT/G2chIBZPHS3ZWnxoKDuNTduP5v/r/EFMV
2nGho8DmntvTJCyfxKwG2dY3+Hd9U8ef2SAPPD5GAyfph2wm+/VwUCD01tONBRdH2CYXw0PbewEv
uuvjSpGUzoGpU9TDboFapEYj/cShBN5qLuDMalqc6qmXmncYD7noB02v6L1ofu2I65UwsSZZ65MS
MriUIfgIZLyWpmBJKTPjk/qDt91NJ+kOB8759TppLF47LnfPxo6CIcg0g7uDevyrYUH+sz8M+jw5
VFQRQxh5GMuAWMM/9XogDf3ULvY7JqWr3FKE1ObVzkrRD8oK6va43WDKuJT4ZwGGnpvecfYxYfXr
BJLuFMiAFHMvPPrKufAXMvSPdaoY3b9SdF9F4Kl6UAJKIrQkViCYhtl57dbZIAPnSjC9E1yEEhWi
/W5TjXcSI2jNVo944Q9xNO9yoQo7hkrCvE86GCxeX2X43T2pxitk9BONEn4X5q4jSwsyyc7nt4nw
WDklN72WJYMphNZ5eKNwAwTyRT5cth00LRAmMZU+qb6B9FXRBaGhauoYbR+vjsCJvM+xgsgjAZ/e
2bVK89VBS4TdjqCseR2OurgJ3mJdKBRs6taleS4fHQgPcHfScBsEe8ZI0LLdg2vGEDvBZc2gDU1y
0sk6uU2KXssS1l3UVfRBU79AqdIZuF1HPuIYMNeYTmjXyzefBCJYEBVjM5RdG1SO+WZRtIBMD4SW
znjQ2oZ2bRRl2+82HlpReR+XWhpLTkf85wGLf9xneUkJB6ThKzSy9HRpjZ+n86dX3XRAxw8DH5r+
EE9PItYeaTWvnNwpIby5HbzBIuuXM5lXsxtgOC+hR3oOGBMoIu6Thij6T2X+pZd/qrawAV3FmSA3
fBn594MjvqAdSZbDATnBMxCqg2iZJg4gOWs28avHJCRUtw3XYvmes+KmgIMREf14llvMmkzuoUkn
etUOREg8ZihM7H+hwMaxd8dVpVqxLWJIWiJ7nzQkCh9mfqEaQT6hauJFwmDT7EmROWWG41P1q6m+
ZPNjWeHb6HxDRtCU+uLj19BusPaVEviipQmkQR8zDDIjbm8cZ1TTRfoRL1JekOZTP4INPmXJHwbb
a3JGtSgO17/LJF7fbRQMyuo9NSmmKm41Nl+N1YS2rJ5nuYulFZx4e6Ff7fn0UPCZNPNFaYLf9+l7
C83sVdOc9Molc9o7/JSQJCT6LXlXy6d7XLN5WErRZ047LP+Y4Ei6Z9Xvq38a1Wg/pi5D8oqHh1oW
89/0Y7ztEEEeh0qSXQWguNfbWfCva0kLUx8Vh1I4LAfXqWqP/LddjqpEHZwh6ell8YJ3IxP36rK0
UYdudfoeMGqZpCLHmqQZnF3rV4jjlYUjNfdYLyiY1ufTqqg7ae6go4ZuENqDdbnYvFc7bBTiLF0R
ECpIlg/kmteq3zEc3LwqxHZ2nU8pyzTdIWC4jlFSQM4FCJnl1RR33cVpjw4huSs9xsLrVwTRqmW+
ADMkjJfVEheMNSV1Sj1DUN3pGVJAYT1aKulXAtaYkOu68iGWH95emosVuw0LNQ+DtsATzVBOOIpA
ACpbYh9neDfwb37M5evzip+MhrxWFHUBnt0LAajZcPtipQais5pvugx8+kw9tctWEGOPtfqc3AwR
KjRV1Mv88QDpQoBuCIWRnYJ0+lFAMqZkCvEU8zSrW3qS10GIDK7FW9A+k+Hd2OD2zPX2NhKEBIxO
aOaJ2Q5sVSQ8f4PyCqZbdZJl/Xj/19nmBLs0S0ZX/X4Tvn5LSWSQkeX9oIWRt7OqngqpypyY8ibk
n0TQ4fO/WgQtIjDH/NSQF2yvVGyvLq2OWs55NWZneeCaXuK9AqN2cMunCFzK6PW2DDLrY3TNFesR
hg4GWvyU2BVWEwia6P1vlbm4Sj1U+hcFq90sLqVUIi/wSjJCpmiffUr46V7CcwOpvb138OWYU+67
1wx666ykx8CQ1EniY5lA9S0R1JNJenNBzTMipiL/FVDXvrSOwEoduU1qKlbaJrSoTpReHj/cGfEn
l1Q7sMb9RPtXusoEYzWZErAEOi31M8zstIQw9XWs2+fFUAUYHRXTSsD32PZc8S4uzkuJyg7Ohprw
YJXjzRDnWCcO/HTSnnM/qNPWnY1PrKYrmqiug02d2WTUK+qzONSzdmGnbxtUVM5/y1n2JP56OjgH
EC+7hR4dwEjMflr93JpgyYjtknEpSS/Sp//V4DQM4OP0tKjrgj4hOBRyOkDzrGnfVpfJMnT6fc1N
CHlmvb1S2qQ0QoOjZhxINELxy0WAUz07ediyIToqY5VK9b9UQraihdv5SjXVc1gZlWzMlmMN2Eiu
543CWDXdk1Q4fR5J1RTSff/+mtlis2lc+ZHVo5J6eCntDvPXJ7Go6cu5nqq0u4Mn/a7ipOlkeqQM
8GR5Cjgdi0sAQeI9o+n0E8UpIUxR2W0NJNU9zKKAOPQl/uoaIFoKqNsyEqq8OVrEPVpzXtHNAXgu
/ByeJvVl1g4Gczx6z1j2QiHajgVfhtOU0M3cR5/RwETvOzICIrh/zCTHsRTdOvpgsyulouM479qj
7cM8a3c/p/j651atdXJSUygT2osR5TsISFyjM8LcF5axGE6MKJJajbxSY6gc6uKWfFpg1xLB6H+J
yE6ifFCnww7lJsuoYPtMxCFFty8VT6LomPauh7+OhaFa5WHXQYExLkBWbboueycGt+3nvMshrCFf
5q3q+rBCu3GHHPtKmkph/zXSF1Mn/hVNW4QCBJl1NpKvTZ0Xor9tvMEZbGt0qbpg0nKJRVxT1XnK
9UYuNTXtexnwyfzwiRiSEjBsjMK5bxLW2pl0HPPxRf3yYSHeb59QLx+VOpARpP+OPrfA/KbYWr6r
Q4jLTLwg+k4IvaMhoo9ZvA3SPp0gVR++8d/LIUUTiViEEToy3NIGUns1gFQI0r7dwEBsiO1s7+BF
wkF+swtmLiZl+pU8BnYKBo7iJ6x5etGSQsm24EvLPX+L7wr15CQUIPzaIsTeRpERS+uvL17GfKDZ
0MUoicwIPT/ZNiWqTSDWeCtcUfbm9gEXiPZrBVMJ0ifK02QD5EOteh3W55fkcXWCsdUtQyDBB9og
iIVszjpL4q3GY28cPRptbhK7yXNBgqwa8XXwnqXxFPd7j7i8D2bFmlBGIrai7AVx3OynkK/XsmVV
VrV9SILYpG42HNa0vbplHf7bGomDvRSC0a3D7744Xo22qepmAkeLZfG9TLZoDcdEuWES8PwyS26q
axbgwmTGrTyw6GReGUpi2q9GWgKcaARfoDSK3r2afJEhiR68L29zUsFyWA/ctCg0OSMzbRur0xjz
YpQf1xC6NHnHlHLts6lPZFzSRxzc3AOlEQGGW2hq/zMxRsOE5hbjWKFGTrM6fA04H3YdVA8kQ9Pg
+Cby9nBlrqNTVV8kgkhJwm/tUgrtzUDXJj/3USM8PyKhg2jzbHGktSYwXuy8NAl4ICTpX6J6lz9u
I3eQ7DMnkzhY91b9ReM3hWAz0ShItdf09QRP0JWUrnfupq7+0L74zXiaYySf9FzMMV9JueLREIp2
eOd3kxfIJXyvH2sa7iutOuQHTX5MlVhqaQuGo044vUmZ8oDXpH1La2tZY/8UhntwJmgkfFn2biRQ
5IaH092kS0v+ENNeZU74QZUZhrrxNRTUjaCQjHXJmHEBWAx1CmLu5GlD8whmxVR43fIKO4zmb8qR
aw1pwybCHfECBdiOMX9JBNxW/uyMrSOMo5ZPuflhZpQicmckt2+V3gwp3lAbUHBaF+DLG+swvLz7
GcsLNfe1cWj/BAYiOxXvmrCmAOxihl4Sm8HLJ8BZmeGJovKVfv6ELj75O5HT+gy20fcG+J4L9c4S
PbI9n8W+w6GUPvhLXYU0jv7nVgo/Kcva7nJFbsjuRRC7oqBeomDhW42/71mzPlo7zWM4IHUiMU3u
5eneZhU9fV5D5+636RShyVyvsgIoGeQ3B5bip/tuqE77a7BQaSGDc1RwLPiLnENMNUIGYPpHuI96
QmU+nMH6RoyJkUg9nBq/MRqO10ERz7Xj0x3r6wdk4cuGnqhrQ5FS3txsniNYPBOBywGA4DxilGSL
GrrAtJH5jG64bDPYuOirY2apl3wkqH6SkLzgT5776ski7iZV0K2USgafuyQtAuHAtdbLp1rPCE0Y
R+H7h38EgIjqpxf2Yff59HIh5Pe/EFiyPK11dhwwPW6fz06ujdAu+AFCXDAbxDyGe0xCtxVd5Rj1
/GTURRlCaCzPfCt3Oe0ViJr55kHJpOTuri7jFKtLEnlxa6dfhWxfKN1Pd6OKImevEh0vd/6ravXL
CeNA2J2Gjy32/drbq+/yf+ex7KXkniA19CPBECVDHE1GshwCFB5E37R3YSsF7Gm+WBb8PsvTbWFc
5Y3jIkDLu2ZR6r4zJcRVI2cJAC7IH1/KS9pAlIsH9vSgmeYrOIjABWNrPIX+N+ttof0RRd9r+8zT
CV7hbgFh8cVBcTD69fBtRwOLgVf58F0emXp2vBuXnvNAVHRSHK5wapGmEWLpF3sbq/8cAnFjfiMn
YyY6pOWZoWfvzZnB3Ga5xNkuB0GoLkKiNlwbWv1ftpCSPjfuc3121pwB3J34kGoW/BrdaJ+4dYhe
ONRcwFinygsPhXXZlIjDo6kZaxME2qRFR1yO82XtO9MNHxSeLnRrMvczQT9sMHwI7bhc/t4nrXIK
N0aRpEmjnbvSp8duZedLLeFrOZa8IR4BXZHrDIb8O/pFVV1MCkGlGFmEJwkdkgtyi5LplQrl3YcC
TlPDRcQdzHuBLQD/zwnFpg6NsM56EQwpVOYu64PB4tTYT2++eZBXRGPrlvAmN8y3Ub67evTpBrkY
aw2NJO/amCD7GTyhD3zgwG5rh7mdogQyNm6KEfiFQn8rb9EV90BFvt+0Rkrc1X/flIjdoWzWzCGP
XNhTPLdqTX5NfheXKtREn59H62Ra5glc61TFAQfN324Ydj6UO9HvIC1XAiX6P7ZYbmk78JVbYkw5
dkvbW/9LW1VN1zWXFj/zWqxV4Rk/E0uacDCX0BXCBS6mRDc0RL3jO5s9JdX+zsdBTkGiMu1yx+mU
0fWilI7BGtZOkS8zI03QUZ7t+nSXB58SOd56SdTaWErCb3xHJlMeJjv8mUl2mGqfw7OAuY1bx0g7
WMGqoX42qlE7ZA6gXjJWsNcfU8HlXm/mHLR9O1Y0vN0/nv6SE24XmMMtZ1hzeqAUX9Pd/gw0sGCE
0zoQ0AtEkl31EstvQ5ltESJAH0U7SVH1N3cLwMzI5OoyOEkcoGYlao48KpzhZEtxeIBjSS59lVgV
0iRTyxGgI/HxcNtNX2itchVHPBaO0WMlU5+T2/x58xn49XGRp78p1cXQWt2oUnzc6gG1ZBd0NQji
4pgG8ui13lJO9f6KSvzC2HKkBLl0q/fly84Rr7SKbhiW0H5C/ad2lWuzu1UEkGSMBKXuiFienfc8
6SEHUtimtfMkIgAwXXzzfUKmrM20d0Vxqdhg+0zL0PmoOkRZEyE4UMq0uU8UPcv2Rt71rYN/ltBw
bhMFuRPt7eprtxUVK1GI+KkhWIxiJBzVJeYJJpluDy5LxPrP7xd9nK0g9WURo6ycKY0zJq7AuLnJ
sM6+nmU+FGcGK1aXon1JBWprwsagrXekVmyB23wn3rNG27Xixb3+cQPzkClg4NOGvcwennJcHgr7
0tyHlm0yp8nZvGRl50SsJaUDa5yHSajySHNy6rBl6/SLV7w2Q+n36mXux6JcScfbRkE2NkzHjRh/
bvgwLe/lRJDfOnOAsSC37fF/CV0O2mfsJyoChuqurbQ0WpUqAQTortG29wT5u1RQAqych93sZ25R
9T2JwWMRyIRe5z8wZfjIiZhy+JSE4DDbi1nPRGg9Tc8Rk7F8hVFfZSnCSnPmnfffdCeOd04kByFy
HPZu8mCIgCpU/Un4pyjnzNw+DcwpQJfPtEHalpxCxJcyE2tD39bUMpJkG2T+kpJ/oqw4ogUsvkdL
FpieqYNyAU7It5pH4NzG77xMEXdhnnnFIwkP8wzJKX6P2zs60pzRvrQ21lF82BP+Nksc+zPP6YZP
zlaicyU3Al4pc4IaWjYyqEOR6CC9ODth80l+kPHtylgl6cB0Jh9Bg7ImJd4MDe2yLvuspHCp7Dbc
dGmbMPCxnMGU3MqSrIPnj543dozEfwxVShxIceOfMooZeoXwYyVa+1f8f6OAz4B/mtPN5l5yrdEg
WjRiN0ASYuDnAEt0XtgqraMkpWqPVHeH0KIOTC3FTwRR+UrxQ73/q7HBDdQle+3n+sWeaEVvNsLG
0ywLAgZAzxo+4gYLcUrxK2vDif6CAXu8LTqzqWgy+4NIayf5WfhxFq0BMNkefeybrd9n5wn/hH2f
B6b/S3R1SBGlqxybtcxBmBmaOotEzGlbmoOp+d+GJnl36dVK+aSc0vLa8R5HbMNi1g1l6lRzo20Z
EJ7PbgcIFsNR1SGHXmCmIW9HhWy7XR0vv137tDtVNyMkSmTdVuHoysEOD2UI2K1Cd/cjTDereH3W
tkbJF//y5DXp5ZlQ2KyrTFFm4jJBz0zAXOdgw+SMHZCKgHRfL3KbbNdOd79Sz+DuCD4KyoAhGDWr
cZRYCu9JqLTtZCCqzw5z4+3RXbxFSySJGzALgNkSI9o9G7X730uDnxcA5S7MEqZDyGkff9Qll5jD
epWTl1W9mSdBi4aYH+Gr1Iu39r6dKRiVApyj4lgiB8AoBRwxywLTDGuTRJ2cwy5XmO0QcU/g7djN
b4qpG2U0sgmv6QObMcMzvAVOTtn4pXXiOXCKQe3CksKIztYIgCougMutv7i2s5RPmA02OFr2qnNm
MQq/UYNuEt9AgorQY82HBqHKzHc+A7PSFTJsANMBmVRvfiTankpgJkm999UoqrbFaKrb8vc+EFik
XzLmRqM7B7UIfCo/jIYzznjHh1z+8M0uzP2lWpgz9W9QA7kmHAJZG/pkimv+nY39qFLVGY21llDi
EnOJzjtYtQ9WoMvDoSne/Zh3LFZZitQIrMCLf1E533ACnmuZ4BzdawfuSHzxpVfkyHfASbHkKGfz
3J2sxyd2cOmjTqFANaMwjhmaOhDmugVKk9Olh5Jta0mUCz4Fxk7Gaw9Bd9ei/FdqRoaKelk6YEY7
4lFVkC4l/C3+70x1KwBjqaFMF7HTuoluv9Vmox878jNE6MovalPRfCqDJ4IZ0JSZJj+BBzjhd1zG
Q1UYRE0+a297VBGwsdZSYG9fhWWlc6r0Be/qwos+gRlp7ID4+aDWVsdgJ2KZpW23dO7qLPQJYl0A
W6wGrCMhfK72lluarKzLiuKZeDzMzeFFn3rxI0IkfxvAD1SFag/3EtFMusCVcrcbNEbuTM5Uno16
Vh2eDqJV3CswVfzr8LaHgIEBK+2p0GO6/IKnXleMzJzf55WLrn55cJSwYPYWfA5dGA9/LQDj7qDG
kShkk9vxq3w+/aUiV2bEgazLCgav9zh7GG/ILK5faq94RLXRgyC6Bzgax217rCVJ8sFvuJWsFrC0
QJmzLx2g0Wissmga7/PinI+Ep3W1e5rMg91cKTZzU+6mwm/P2tF0Ju1vnW4FJQJp8Lc07hdLa7JI
33G+aU3SEF8c8a+xnTKjBtxT+zQ+iyrkTUgzjKYPl1+bh920jOTaiQNTR8TXO3NaZIKOn/CCIdB9
iQCQh7UAQzigjLr4MDihQERYyy6A9RoIrh2ExYtAVBzkU2f4TBfQlYCgENB441zKUaLDFNOjG1fF
ZRBQjAz51HEwc86VwD5A7ypqwHjx1U/ytXEaWh2wERCi3kuM+yj8YuPZ9nqRAq4brVYHFwF3piWB
NYrCI9QRwfx+8hwjo+MALnOi+rOQBlVDGYrjgXnCllA0wUwoBHiOBQoL852uojpOz0iOkPBYrqIm
GZeWMl/lvb0LR4ydJNGwDJHPwK6i4qxrgLAaVXQVb6gzSHt98JS6R+V72oAlth1YLnsqYvhG/MZg
AZ8Dh6xlRBUarbCAa8szOXvbxDtzvXHHY7MWDwx0xQY+jkR/CxymrW/faOz83yNeohE8claI7a5a
LZGUGOKNGGc8A4gVLGkMC8aMSS1zXChUHfdmK2+k2vTLXXBXJs+DV8YFCjcbizKbMf6emOm8kPte
exBKXTaV9cJF5pDHauHlAF2fg2SY/tPk7sbIcSSi31PdBCIWM/aKujSIan8tjPRtXUcGmQ8hCJrx
p4kDPQM9PThR3HsiSoDztoAAusFDEE1owQhgA84Df6DgYr/y6HV3pa1w9kDfRjnxbaoFbgn0DGUR
xZ1+ySx7g6QSs6K8MtS08bArVZuK+4kgvvum+Y3cbFzjvO5y/3IE2BQ3RBci0U60vEqD1V17+auP
SCAFQGhx6xz3p4IoRisq2QYsUBPDSMFP5hRKoD3By4xq5GJMbhOjc164eI+uKVZzwRcUD1/5QEZW
3Fbwdw4MpzJfdV420OMOiYjF+q3E2//zuR/OfiIcM0yowvH0nAq60XzV4OjOTTCXMUH7n5/mekyy
HlV1XaqEJhPmDMvVS4OEIKZw8q5r+S6RVasOzAQd4sv3xx9Q71k2fXJA+TwAUy8mlKMBKjL3epB1
8XJoH+z/f7z/eCrRlqxuYs7GUUj0fq7HSuYLq/nhjQATxvXMkBcVVfLyJK1YuuYZFKjahTjGSJJ4
u5IL9KG5UtbI5ru0WU+UE8LGslqpgP8j9Zn/rwKyMSX+Q4h51zq5fiRVCE+LCGS+eaN4cigxpz6E
wl+iOvFp4fiYkd7kfTY72S3ke5on6BhW5S9obFTGPIO5ebB0JXDZ9p4GyJZRin7jHzGPrPX4DWaQ
yC5UEpJOisQN1JKZsDNZkN1aKlj6lxsTinTRxOQEhJTrTKtMDvuXK1fsK8+Ft7TmS3yMGI+eFP01
ipgeQSztYy+SevX0z9uXkzl1dNjS/eG80d/uBEtjNeaA/5/nmX1beCYoch8DYCcmt04NQXxI4yZ/
vqr7H81477kmaLAmtEp2gzFtzo7zle94M0ObvbAV4sOoViQr24yLXXHJahHwBRTcRTf26SKAP3Y/
SzrRJ0y7pj/OudPMe4XjgkDRBJ6RJzMWYcoabR+vIKvmO+90UuYSWKnz9uhOVrR8tqn2O2JbOTTS
IU1UEFj+uGYRRUyksf5jY6mrfq6S36Weg1SZnGwEk7nndPIRn47QjR+xswetYdX3U6UKCCv77QLt
ziyXirtsgDe2bTv8eZU2zEBf0WuUpC+N1h2fq/yWM65fqLdxNkx2mrJwGeXzgfISkVGzwWpnm77y
OHXtpIHi57iGyKlSD4TisVP7YBFtxXwylOhx4yyjAAGpkxOfQT8+P62fXZ6IR4WCu/iZ92SNpQWQ
AIJcG3ce0eullxpV7BQORbrd6WaRIOu8rmaIJ/STFE6RlBz/eJIUfhGxcWuHvsRFzl2nWueAtjiT
xRNWrDKKpd+tfQ7sj1c95cnTq+q8k4glBC/6eHSs8CfH/GtjUS0PGv80Q6PaTwsWxyNNOXzQxinA
GZP9ca20e029rCz1pFhnXH+1tCTA4LfHS21b7wh64ziQtJaPwhvqLyxjwT1DqrvKWgcZeEH1uaJL
qtdO5VZ44tW+zVrw0OZG9idRcwzIMDHszMtzQyXmdgT+Qk+hVzJKFY9Ra4oy8hpQFDMe3IRUFdFW
Ma/ntVHPcsL/4BAMJmXArjDytM00rQ9EbdCBqtOgNflpt1ziu/26g5shwqkGfcUo7AbTqidag1PZ
Lp9tZY/pf6H9eOCbEN31owZGVvEP6GJgwgakHy8bPZEBPv+n6udGWtSoIy+EqNKvuSiNX1xb6lJo
rMpiXpc72cHsd6WPFUWW1bt8z+WU4eNUr3C+ia55zS+vQIuTZKO9iuS8AuBwl0kf75YH8Y5o4YeQ
ApbL50C/7QE4u5yTOVzEcbmScOQrVM72jZrsx60qE7cb8rtbcj9uQtoUxSk0axEgFgznW667lxZS
45F9xe6yGbdIwVgTivl93lpj8PObn8W/IXNBSoAf5LbRMLUI2reWtEsGBJ1gUD8oZCdsmmhSeqos
+YnnAi5HpePbP6qmcqQUZprUZ9CFnNBQEILeG4y83HbhmgEWoIkPN6c6o4/m3nz53OUeGNVqXcpy
SrOaji9h2OoDDuQjflmIpccAtuV/81kEGEtZbCXhApzqsbJyqdpVD3n5gua0tlUK3SObM5ziERr5
jgCGb1LDmstBHnKBnXIJnDwWXlhoJkfzFRzbhM/smit58IekqW4o6ZTJDMYBPhlNMOjA1VuV+oek
R17Mbjo77KAYVUwhPuPBm+rs5xwBJjbF3u8p+tSCELmwGC4Ku9yncKAt4LvmUnhJljsDSrrUrsWd
8Qg+s4nzQ3eoJqBJapsSvOfu/MfjlFoiwRFeW2ABfAIzhWDaUbreiSTo7agq4LwZxXda+cwSWD3F
rnelnUhJkJ9Zq4D3T09Dkrr1Tlq37zlOFpHE3yG9w5XwPaqNEtRF5iM0EVoUCpyWUCWK9zNj624S
/0450xINnZIkoqY3zFX5hAat7vcC63FHUdtDNRVFCEyd+uJx6fAbAYSZWsya4zzA62B7zjpSoj8M
n9/6Erijk22xfMFIVpSNaWz4TgvxnN1uZIrkemdMSydg+arfnkjXd3zpU4Qe/x2s4pexUGoNIxY7
jPBMoDNFlzVdJtgLQCqVlbV2fXFf4ZOEJMIma6ggOwnirQXGHzffgTVRc2jaK0V5/hd0DuKelwOh
9B/6fJHLpdThGeg3bhGWir6lWhVsgBXh7BNGzbKH1/EPbZT9pEHvruaWnbqMlwxhmuUIj4+/ITca
K9ZY9ut6AFJiOfyLNqZalqrhDG6z2cX6OdbrJNvoSzPnuSt/+bvfii+yCIv5IIajeyxZopwaXKUF
lYVsXCVbWHoIZ88/keBRtWDZYdLvvbh2KFTETgOxSUhiVblNKaRHpWumkG8cyBHysTg6ScbmJalm
wIz3Ctrpz1zHksnqlR6isGo+G92KK3F5T+UqgEDOzfGw1VYI/p7Wpz6MhmIG63JoXJhoUpScKfGi
+IaefPHNFqbZYMpNx7DD5SmUviVx2LILjae5vN+LyclHkyoHBTPeN3G4iz0vIKCvt+L6ekK0SO1m
mMKZFwwqsm2WuCYMqbw2ypHDB4whVZOPNYRDRxPQ1DzBUcSgAJzvCnPzCrG0Ggi0b5k8lrMkghDT
VvzvwRKhcM7+embX4eST0llKovOUUvRS/mkZB5qdQEjZOEUTy4V+LiRy2fKtfHerYn/xC8eOKfpm
BWwq7wWvy7XJe4OlUUWh9zA/LDrfQCqYkbjkdPZdxRqdBnE1wYOGcCUEzWshSs8MRH8uPkpCh2MF
f3pBix7sPLdM1CYuzL7k8b1SFy2RXRQYva/+vk1+chreswVEZlNPArSll/HKrwzTogPj9Mzbb2hE
iGoe/PgUeusRVxYS5PaIkCTzLP+lZGmXJK2cJEs8Uff2lNAxUJxia9z8/LC+tSZ8V8dy3hRYmLuX
2bymROg7s+O8iw/fTiuc8TghnqF975CTJKVjEHf2zwe76Aojm2XXXmORm0rWizL0VwoRwgbum1ut
mxEWVrzovehpxd6AxqR8lIpmRoPFTA/QFspImfLhBeiX5GjaLkzDR3nXrGwa7LBd7j7gCkAmTPqw
pBFgXqTLL+Bo9RXRnbeVvP1IOifz/HmQMNCMhb+M8BGh9ar72XfZSNVxk5ZLIaAf2kf7cgn3juWj
AYHvqjmu//AExhjUxjU/0DrImRbUl+Tuq/oDrG/0drZqkZWjHVuGZIYYhRDEg1E98/lqH+Poi3UV
tDNvKXMJsiKogkmMl39YDcWlms5q28xWrjSJobXZcMajS9K0jHv2keoPbJ7kSMgXgrT1Vg8x7HpG
3hxUOcng5ORCY8uOcCMJ6GNUE28wbaRKTnrNtJqCP1Dpj+rCsJvtU7MfjHM3wsILHMrAadCQ3z2v
uCfwpW9jBkdHsld5xj7apJ3Xv+syllIvTaUjS9eyy4V7Yi+VRJFabaPgZTfLGeXZdQfgnwl5ADnm
uLz8yQyu007QxeaVKHkFG0fm9QSpgpwzMUxXlOXVaycE1wkzPftp1+8+yl6qni2sJFY8pzaGLS64
cizfKES0V2tw2calckENh7LYUs1DZQ2hLiizYybxlHExqiuxcARdcxmxlrYKDjjqdKERv/NweCZi
87qFVvRv3dcO8WPBaluMoWZUbhTJ9/+jq4QiZ9UhO00Fj6HsrGbdqzEdXZn29zNc+6w1OQG0PPWw
9SifMkoQDFwOv7WzwTlZdl2jysFyYd1qbIRhOgzXIaAkaFimeOSWxY9rpaKbg1ORuOvFCSNLD2B4
ke7tm/JD7o733OmFsb/KZfqX/liJCtWQzr3QFEq/JJ5pdhId9gWA98+/rSFWyhI/u+X/Sls2rU90
/OnZZDpTpIqj8HX1C+KPFUshCFnxLcjZd0NqTLXU9iAMJupbwlJ5sZ/OmU//J3nXEOE2cJd5sIRR
C+SEFoPI0tMH9bDhJS6hZ7OTmnLDmGP6rQ4SqLYtu8dYAWSG1vB8hSVmDymtLIpoL76QFgkvkWWi
caQ0Do2Qps0fOX9mYaCG/UJmA+HNBmPnC07E3zpWGPLuyK6zA/brg94xL4ejvdIgm7WwSvekNsEt
p5voK9tVPu4WqHquhysir4XFizknQg7pX417X4DkZmnSNSOWlOrCvVXfStsPlWLWboMWUHdhjuXQ
F6z09M+mIVPrrlMzfhamG8k0mH+52gz2oBRitSw7YUXQ4qfM8NmUhYQyTyuLbTCbgNBkmsF1RmCZ
/4YkamZoVSglvb4YfUc5SQO20kA9PJJpp+ZRq4NL83h13rhudaE8sRMn3rA5wI06bLuENwYcZ4ws
KX0aCSvRro1cAmqJP3uJwemUE8b7+RMz8bFj+U5FWjs9SDxvILgCDXtS5hp3L8ZuA81Bv5xtK5hj
wYkgIRfkXg2KVEkYbvqT8FvyGWcPB12OaGly09tk/w9xwz0aDMniS+cMhP6WvG0l5ynaCVuwSMi8
jbLKdH45Mrm4lAaWZCJL9n5Gq5dYHRpS56i/NdnKuIeDuTn3VBBnop4As/NA/y+dmRP4fefPAj9h
5eKEe/zJPsQ5LtZ42XdnUutWrH6DXSghQpjLcL4Z8VgQyabyFeINAaJjXGZ5GjGoYDxMrpht8CDj
cKQDm5/81UwAyCTewAPelk1WjEzjP9rTdI4eOust+2qbBdA+ztMU6OOeFl4ykXsWnycUqVAEQjJt
CoqwclmD1DoxudnTiaHaGEmegnQQ65WrcNsVfmlpQsm9MJwMs1afodH65Ao26K8Ct1PlsPjxgBmZ
kSJGBXePDiwM0SKSuc3/O2QZBGoWSWLaiVrU6qkZGtaTdKT4sCRooS977LWm9x/u3SO/ElwbyU4S
wK0ti/kI5wizw8PQHTOV3zPS3kYpEDefv9S72+v1diPMqjcHs19zbSE3nipNFsm6KwGtzpj4y/SV
GfuA1JLkzm14Hc4e6054vydl0LzIUnDLGCxZkRYY31IJ7/AAgDFsNdWt3KJlsZxFVns+HDehD+0T
WL0L5+6zm7jsQDYQ6tfaR/5/b0OEq55SqlmJ1emOQKo9N3DCUwfqRsJtB1XcIfOfN1+c9giehzvM
eXIG9M9basoisEr1Rl9ViMwe7E2EbUXDkfS1Dl1RIJ+2RAxR/PjbAazJf7ZtcWhSa7PfUD9wAex5
wj24E+rZT/5Ap2cep6LDj4vGdp9NOA1TsSPR+DjDiM6cW9vASBJs5ZKjBpg9YB7EdXhhJiWMBIA7
MCIe8ggCYa2y9p8/ZN7eLjxjTts5d99Nf39fyfR+KWBUULaylMENm5FM1khTioIjzm7elB+xDGpS
5Kmb6zEzpANElrAtg9P1/f+pqvfnphHXpq71blmCZ5ItI5zfJPj17QOoVDW0ZvlId5kzyEAbUiZ3
Oe9aH/cW6kqOs2ax7PMS6s4WkAch4QpD6DWnBpooXUYWU4qdQJFh8JME9riNFLGzxq61VJxLUCHu
N8vzW7iigxdjuyLlVwEsrg3TP2ejnqg5XwG1foBCvEGXxuF0mbvD3cf4cutor9PJhzbMolXgAxAP
Vlna++VBfhrmjjMfcBqzjuVJIpHntzA40+1aceEyCazhTHtqFgmI998lQaSlumhGks4+COiaC4LV
DX3nDtmIrGJigH3HynHLHLpHsBOqaalir0g01m/wKdeTAe0fTgI7CtS7ZXGkFXqSltFPhR78kZyU
rzVWs2gMSd9kHeLBukDuYzUV2rPtp2RC0Y5AMUNT+nw4PtvmzKQbA6RKn8wAP4H3ulzF2j/Tr3uU
CLpTkRAPznXeQC6D3+TkoR3yCbEC35c7tcMEXv+U7Dv7wn3RXKz9D6ub+vrTHEtWLaFIYepecHPk
80Y4W0kbwSm1yUHbEZPyxifFLvt54i/V05/eBYBLYsXlIELMvh0xXWrHhGpcJDEThqVLqtFDBNui
AZHKZ2FU9fD6LQ+TRFV0VkHsbsTUjVXRzQC5IXPCmgNuSyAisXGvKLBadrrqvIUOiPoDx7kPz50D
ZfEYZpONUOYQSEKqv8XCs6t5b0+PxIy+MYlSmfH3pX5KejAtgaH8XwR5ruYL7QfFjujOy02P/91e
jqEPvXRVGEk+AZbNDYaV86sJ/2JTLi/0QVIsIU9eE6fc2Rs2dtKMWM31abPBAq0W7+xSVxqbHuzf
RwYz5n92EYRx8YF7AnYZ7CBJS4zp/iIVY98kNIDh0RvA8ae+zAfpy4wb5sX0mfLCoExnZyMWor0y
AMIQeY7ubNNOowWDI8pWz5bqBqN6olk9puXmRxWw9iESJRi/0F2ADHfzJf4IMhJDLHBpO4Q7Rezs
oE4odEIP1rVoWaZ+OaWz7cDLUtSmDXMuZbY5paUFbCgpnyYwbArLElOoULENss7VDHFZY25KzlTS
uGHSN2cnGf4kiKDJiYNeYzFIHO5MmfqyJKkUqpjZrM+j+nic4zvOXElvUEdLaiCXb834aZ985Rjz
wJNJjljo5X5DZJS0x6uUk9KKNMRueyfrfCeTMpJXF/UVv/iCcTW265rLpKO50JLZQHWYzrW7kodJ
dkYYAIOvqcCK8B/qkBPA974DVUqXcbrh2plEpXqH+Gvfkm6wMjYad3GS4UMQnscdPLhRohjdY82u
2BeJ6pW590S6FC00724PhzjKMBqLKyzOOtyaN00rZNtiR0B5jE4NFEFOAeKH8od0Q/jl29Nv7ojn
wKw7PoGhhx29z45zdsu2oTPPxQlUKMwSbBIWRw/pqd1SuhqyggBeHXgxR9nluq7eRvhMTlW1NpZz
CAbyi7YUqysdp6/wklM06szhTWwpHNjZLYMNLAH7Z2/VLD+OXpyKc8ffhD8ZuKxCnZDJby+7b0Rv
xGADxDC369gmxc+uWtvTmLcXX0KHL81iUy1908d/QFWBXk02j7b9KLX8/WPNjDxTVo89SHTZEujR
14ir9E9lr9OFGvMcuokkHR8BAR6mlQ8fvhehf6fATIaP39KE31D1U8sw08hIDM0OonIv6pDNVDzT
0MkGqoIZfa6vgm60D1jhI887+BQ2/7+yOzgVi9H+jgJqv0klIsykJJprmFsM83py7DpnV3appDW/
DAOvMh5DVydFFyD+dFH8SiF5BGjUtHkFYlabDg73iHguFV5LaCQ5oyUTfeOxKGv3KYUZ8Xb1mMzn
q9ksyZ6gqaqn2rEg8WM1Cv781DJywWtxJm2trdghFWiKlHEffhUY/zw97t4tOvZsmjsC3f3Lr2gi
ttpj/wATCxA2cDQCZKYMVW7EksFEFQozWtYheS3xvGRR9Lgl2xY17b/HdK1Kn8wrBLGGzRc5U8w7
xCDkt0MRJViAJPxUBXZvvhyNPcuV1diyiEdC1HsHAClMA3zarljsdYTsUB9H1dcC3CmLWPGXjFho
av8KusutjLldJIFOwoS6o1Vjfyl6eXBHexM07yADd2N9TeMF1Y75HuQfqXTB5nLgai6npUbs8B/m
4ep8Y9iRH04mH+oBqa14XMVqDICWB5hLx4pu9V0kVqpLAIcv7dlKAXu1ISygru0pAkO18i+oioFb
2mrTtWXKJIOAqn2+t58o8Zbp03QO+bpQI9nlWYv5FCPRRK/1DudtBpwQCHln6NX3qbaR1xOBe4np
Jq4n4QpJXHwGgA8Bz1JkknQeqcD2+StEM/eHaSRlG1baPXZyLENRNPcJ2X9Ipb75jabmDDji9QQg
8bP+BNFybGe0DGbVUgVox5IeM6CkVdffPtI6V2NmW8uQbt9P0hKkWRoeSvG9Pld4FScrSdb/wQWN
pE/eDqvDaLzeHQ9oQnRQexwK8lLxVzy8qFw2tW7mApPpM+0d/LL6e1ZwHeFcUwL4FVzb9bDiCcrN
Aw7BsV8eY83TcJJmh5YuQCWz90Ifu9eXoGPQfJN66INF/fnsqz4cbbqm6tST3q0AQztirDpJfH1V
f7vOzdqtMsytwNPqAurhZx3cY7ay8ylAUTvnmnQHcAu0Ufgo31eckJiptPdpuQ0dTyE0CDJTOO+/
mgefITegeCUzZG2UjGufydZKPDDFWbikgN4v1/a8iV0p/wkafrhR2LcJIdKSc/CVWKu7ZOGDMlCs
/K7kEIHvwffbc5tFCZYb0RdLbb5Jbi0vSsvblLGAwkxcXcsDAvQ5GTwRPA7zDtoCvRyoxG8uXHrT
CqCepgeOcekEX20/2t3y564neuC/lzbksNUH58n63s5aKGaW5QqIJiKw63tKrkDFFSY5rYnIs8pu
AmYX29OlN5+VsX3/T0OOKC+XE0x+rI+BJPVVMj7Xo5gAyWpKX62/pUxlD5bpW7aIy7a/o4zGKWiG
shWCifGSFP09KjXIuUcUf9QBE60mMMyKJcnEIc7ZZAFcNGwhYlK/GEilCm7XAEJdv3Imh20THOBe
O5xOVFzvGiV12whOfaWgIv7S0d9gZ33k1N89Y0Pvrik27WBuEUzM2qttcPX2Nihw8f6nZ3zuH8Ht
9sGSX+UzhAUnV8IbM7FJb+ObPyRPXaMH+3PZFGt5dL2VmjqWaMKrlU6Q3RXTD+XuQbPhRSvBJIlF
MNVOIMzdL6giKrDsjYuIUule8DujfDR+UlO0xWkqNuk0idJLF19WPmpGIcjltXbiMcZ2CX7Wuxu1
V1NEaXtvvMcXzBqm5qHZ6CKNw/LjODAN5u/jxvPBBfP+ds7xSzh1Gd3ctBYav5MptwV6DO7S9EY0
p4sWBlatNEoXyLgdlYYHbRhavLT1UaAPZr75/xoIfecD/xxFCvcgW2++46vbIBfT2Ih4zdulEh+h
/qQYfXTSGOElGdCkFBMaMm3F9pUBoXk170S1wdT46tFinWcvC2PYG0h5Y48R2HvpJsGTDXKOpvwM
szyjLvg262kf8rLrBCKy+xir7dD/uPRT6Epw+RTXSrAbr7QbbPKp2khizK91t2NxBn0D8zUmx5xQ
RNx5KVoryXbHwSxTZsPJRn+pIQ08HmOC81t9Ug7ZWi+nAbBG3UVc5yWMqnntb76MH0DUQK/tgdkN
awyHAoQ75hLFRaQsP7RMjAPvcCvu3hPqWRmB8Rsuld3twViqp3avdN5377iopfnHErl+sYcKwgTM
XRsVBAfzVeRyqYDnaAzXirDFaBKyeZMjoeolFwE21Qco8WZAuY/7CshAXqfyq1FSRy3LTkZXllO6
wAEUH1PSN5FDhcIK9ezizqMgvXPuDZGpHRvSjQSuTzmwaJO+cqNg7NS9YxD47RBm0eXZe7bgp3E1
1J7VOemEePrgmRSpB2aMz1QTXNxKPj500qUbanvi4/RcbpJQ1GvJDu3IK5ajZM+F4aLmwRtq0gFZ
wRgPNJ2FfOGWzuUOrJjC4qiCeli2m5HqF0psTq2YmOXEWQkCEVsku9odbpsZLJPn+rpr43Sby1/G
5GjTZgwyJLlNHlUeAxFUlIodjHskHCyQJfGzBkXC5DYBW3zFqS1wvrN8cPaC1WNuHLkCjpIU/n4X
fbN6ZnDaDrjfeFUH+gteowakbFQ+41JedcG7v3n/4XgpNmi1+IJyiooUYLPLG7PIEghl5/4R/kwl
FvnAaTFtywxWTsrOKoBmgbYf26/LNeB0qGQoOMcyr2VLoEhv8XQCjtEVvlRCASr+3gqPxtjpiOU+
b6QhoXjfqJ1o43S+BLDLIYleaEjvTlQ/i2F1VRtx1yTN8LKrZTu0gsZP6XaeWGCRRWzXqJwHU0Y6
XgI+WggIVMdwNMcjwJwS3b95Ic/f2J7zjcCpQNPrYgi/U7fHhv6cksdx0k0Pga/71I4R1kj2jlI1
wRFR7WgyXJbCxm8LqW4rYINGPRLaJD9xaqPfoaD7cWASMmXiV065HLEdBfHZneVuvaLA8+sVxS9v
P9emO0sEkqheEnidNmjf3SKKiDJk/xlYs5jTIOH1aOt9bvnsKGoJY26MD9KgEDIyKxFdMC7slMao
YWAMavH+W8eZOMRIlGXnwy/TwYLk/4Op65zqWRfY7/xphOi5EQYlAz9jPP2pKKjZBqZkoVmDs7rO
xP0qGlwC2krn9wRkrysXyOerUFCS45ZdWjWCWPDRWzGvoBTKFloB/thU01XNgdkXi17EZ8h9vHc4
Zmuq8V97iCQpc414kgG+3D2vkENlZ1rYX+hS6HWeqOlQ1XsqLEMcUIrQ4uDU/gat6V231JWRjvfJ
OZmrAmdczlf03wx4Aq3vjTMr5lMsl0mi+RvI+TQzS6eSicfAr5tpN2YAHL1L3hGUGlzkg98X7hY8
ZJ2gVE9vvco6lrpX/EEgyIh1Ko/zppjVYzXKY5SlybNl5MjY7JQdL6kb7jJ9U0Xm6MPsHpgNnoFo
zKoVKSL/Yq79CuU9xMROSIWTBm5Uz2kO1CaTZqygfIFnZjqBEsR5ewwxrEYqWDBOCsIwKq8B98LX
t0+ZwG2QLygd8Rst52WG905NiT+/mtgywSa9dCwemh127qRyyuNzEMuW34NhEQ3iHLdYMXY/l81o
wLUoKKSrYLHx6CCtSYJ7Y5N5bVBvbpYZGzYOuMssw4oS/Ql1DgI7uaBpI234Fux7fqb5sSuU72Wx
3T3O5AWQ8if47t3yOvaAPVLnF57n4/16iEmtbJI/b0i/f7V0RHjr2QsNWJZV8a4BYWms+cv8pxt7
mG4Dv5lQSq5Z7wz7uIFAWm4jwG0VD3gjUTcX956BtafLcJsTUP9xTAtkv97fQ5ARPZ35O5Ojaw6A
7bl2qX1muX4EMjCEqHmKOvRJukfdcAgdRiTfqhCls4ziIy0D2E8PhnXF4LAv+1g9dVT2agkh73ub
x0WjsjEx/oQuiIaqCaLLkKH+dNZwyttLcRpPmENHFt/8qBArSF/DwY4Uz57ufWjrNh7CwokEgoz+
1qE8vEg/eidbP2veoyei+QFemnnZCuOz+oD/eXJt4OGBph7Oy5BHjX7e77+TDTjNLVpKFqQ0r/BT
MhLa8DSmX1m3q6pX4bkNQKMZonkn21qRUjOobUyAqjlmRST7+JX95F+HeHWBW52xVtUtKBzpvqVu
ZIFR2PxxOe9V/h5A0TftP5NZbwMdfxAVelpW7K27OkFvjzr48+bdTLZRJGsYholrtiOapCobkXRU
fNEPuWFtH8ssNKwdSYx9d/HwEMY8x71dW1qUiJNhwHOBD3axSDnIWjHIFehfWkzL2Ld3G2uXqhyj
pvGuH3VKKdsk8BjxzqLDJinPZwk3TAvsf8RyDWmtZoOOdXgNcdLRNoI1HaTGH1k2+odnVKSwOKrQ
OhFV5N+YjSAzys0dQf/7CLiDThWHuCUm0f539H5Csxgyfw8Ly/qk9HIhvQEdllW+weQmxMr8vFbc
OwpNxygp9pl0RBI0pfOo7Ud3v0xy0XdJoaLDXcm5TurK08utiBUDUSGJtsr4mzm3dY3mtBsJ7or9
TuqZ9ymZm7x+rkBAhg4lzsPpI8/bjdfwuFqkpoaOh6KqZ8My0FKttqFXsfVahsueHXL380GP/bGE
gTZX/M2MOLEjW5/5f7cjzT3AjXIw1rNMjq25nGvs3wSKDxzKjs+/aB5XVOCtZ1uE89p0JfR8gDTZ
flORK4gl2GK1HTSlcy979DJnVmEyGMfQkZfz2lzon5LqjJUxVbrqrC+UaLND4aHvZ8F+UwyTgJNw
h8lVut+dnfI5DoiXFGvZAD+0aqRiA1JatknMad/xkQ/rg/9NcKLjBvRdqdS9vm3cRv2BnBaGi36t
ajReYmjeMXpZhqRB/SxVjFQypwCAuoSFZCULgBB9f0YzKBAfexNIJgX7bJR6kK3Tyf+FFnDFCQkb
z48C4lSzelSMhbUfP9Z4qD53PFRD76XTR80F5mlcAHiW6KnChFRfQmnlgcJwb3Pnd9YpJW+MezYj
+lqADY7sKg9YwghrwoaHEv+jCluHMypq49lSc1t/6fwhyjf+kPF847BivIHX9FySDACve2etgioP
S7BWYFdZn0+2mxNR/6+5Pu+vTeRPG/xPMDvA7chChk4phcUY186muYfkgU15L9lcWkjALebqwZPy
pBlTFV24JnZ1yxk2o5hHGYiSb4WjaBE2+jsZTUNvcPneVJ8E0fGh7PVe0VaTN875bP0HX1TEfTN7
ISQhfXpsKat7pSCacdUSKlFasKnGbahnyKIi6QZanVRGqk3eHqJruhSoubF1HHt9QuKKEw+R+gkV
QW+BgQO3wHsbea5nXpqihe4nWxXZMjYwYYTfuggxBfRg4OX0oFKaW0q+BMg9H2zWV9u80B8kwocX
FU6H6ScrkLG/N+TnyZt9os5bSR/jF0xQOOhOuMhn/9n8hfvM15e8GNIg9Ai5rg/qfI0hEFzFZePn
7ZFenxu/+zOVoFGA/0ZS4YdkyWsLABgynSAogePH5KSJFV5x0Xr64Ph3w4CHrtux4FTUaaQqmXo1
1/RIOdaCzy/6+ZVYn++CsrxozyobshQFttCyFpFJRs7xosLkcEI+ny1I5+AjhIxsxR9B6djEyS0u
KNU5BwUn+xMnqp49fUS9ZbF8SxDAAyCHdYS3ZB5V6R+BAcD4XtQFIHQ7Pbq5jVpjpxoG2CNosoio
pTplLsyf215z29I+lueIA3naduqkQ2DbOTiiJqF+aYu4Zd7mmh9sQU52jdhXdNgx4L3IZsF1Yu1q
nSR6hQzsHTvcqjSeR0OF8iMKvmMcl57e7T5ti9i1h8peSjNe99oPZpHrLbwmFCRNDFPsjzi0UIi3
eQVb2vMtQ1ifpWXEzgd1jby0ta85BJNE4R9Kruj6ILz2HzgPT3C3aHcI1qRGVDJTAVahxOjaW/Ca
srfSVXEHswgXbbvkM8pKwbFyrCxmisjGMjZZTTurquDC5J9K5SK6cVW7RyABAL8+IIwzRFvw7/Wx
jJZbW/4ApdBo7xyeMyJ5BCqXPWWbiJyZwC0blxQ+GRYfZauP1yOxa1dUXWCyKfRd8uIQKKNvrMt0
CzZkEdb9ACTw/2e8ACmxe7ERizNXaywG10VMEuJi8ttlVUv70fe6GpyBdZKY9OmosZ9RQ1Qrd+xe
F4S+vdOYEwkgxPKbjvXlXJxiChg9Jutw8FYTf1964xzGUbZ76/BMgeE93kjmRli79LJnlHJ6d+no
fhuCSX7WOKeqONwfd7yyyoO2D7mkWaAnan1GRo+tWtyLhfryWjZ3lMR/BoK9ZR4A96od0udMZ7gz
Npw6CDy7BetltSBYdcZrTHrLFQjJU6Q0gEKMt+MD63PjVJNxrXQXPeZBfQBZ3oIWts34eGKlSBwy
oaz3kpaEWoDXUAhVvWE9Zs6Gc4dz8/7xgX1OfQbI6CzqCS9zqp5Fb67EIHMy5Ai6g6LwAANknn0l
k/OX8h3LyPQ0/XCISvOmD3sDO0ZN+haSE/eAqgVP3YXERIwKSJTw3Tt8kyNtsptNYnTQ0w8RDAWJ
4zcuRNrhuGP2vons3xE9zmLiV+6DPfGUuQOwB5UN+2IuhF8u5awhpOy3U44PRPbY18bct24FEIuC
Vy4yycj5TfGyeALDBpc27sKR8iEyB0sVLFCX7WuGRn2R8KkQP6PMNanU7F8q/sNuo1O+BJpT1x7A
MwAKcq0vXgXr34JJ3VSrGcso2H07pV9bGZvdnDWxuKovepboVbP/gDX95Z1OiQRfC2BSyhdJ2YFc
DVJFFudb4VWg21izqzN4mJ2yIPWj1yijw/Gq+fUzDF3I9t5EqdN4mvRe7UMQVxC8I1KrT2QHuwY8
C0xqFW2g+IIPygQPcLgIG3esd9nAURTlJKrQFxzOBmz1HVCdQHuWShFfIfyjrq+SIcMb1zYaMKpp
rfHUKBVU1T6nUOZ/zKOXfZ0KwB28Mqr+hY/9vCofP5iSglB9toIMFDy0G+Ft2mLWoIszaS7c+nWu
TK+OgikxoaGqcZ6TTw1BZT2SblX1rPScwpNL34AFRwGMjNoq+p6J95npeZOtwAoJp4xwI1ekFoBH
2BxpissWi4FpUeCofFAq+UWs4EkLHJP0qWr98SdcEMHQTkZ0Fgu/TzZbLXxWBn5UafLGms+FkkJp
DU8pMx3gaL/H0zDkWuH6/OMMfOYhzXGWoJW2NkkTTJHWKJPKCe06zMVZhu7/DfRxn0pKAjjz9sUI
VaRMtDmmmEVOD1xNxe7leztQjeZlu7tZ8ML3euyRZpfFLfM0MDmxVsnq573bOF4Ifs3UzItUJguz
v0BtxHojjoqHGyptFVXZChz/cLbk4HaUHH2EYN79iV+NR2Nra2krawB6oAOzVtFqDMR43/pjlUiN
OZebEIeuETXqrX5r0YFVijuejnm4qiziKntSqG77dFgxSVqPODRPqgc7gkfGGNPfFU/7AH4GCHLL
I9/IVjuA99nW3dlLRNlyVWN7881GZTsD87AtFzPDEpIlvZm8FNDujUCOzRJEwdEfNBLB02zsmqS0
jQKUg1Iz59j04OFs/pZ+u/eiB198RIi44rWWWFSMCMeaMjrY3HnuBUHMkS/njPRhsIJduxhOYAmP
Jtu52Pnetkw04GS1Bh0GWym+AmYrQRoErseHVD2hbhB/owhHYoPc7UyYp3SH+z+SOki3BXuE/1GY
YfSWwyy0k1G2PBdfPVKfa5UbM876zrwAWRub+32/WZJH2EAbpe/kSQ1IYVekDDEwCQR0mGQPCv5f
LVc3u6qjPV8F2y6WUC4IfXweHEMwKsvV9zZfZgQkyTOYYu6dqwhOO2/wxux+qGR8ZBGQvl8uMlhY
d/jd3ek5SH/Zv71qWTdcBskSKZVbKkXFVHd1qye1iuEP59G5+OpXZh70Tnhm9W9au7RqO+Ht7wJX
p0KL4ym/WhcTX1abYIN+rDh5HKVM8t6MOoOCQkcfOBTrcFGI7j5pXr5NrSUcRlHc1RNfNzx2tnWe
gju8nC8tjMQu2fCwCB3B/z4O4bmyjHMAK96ahc4FTYdaYbX2ycxV3dhmfyPfw3NNjq9AbqBq0buN
/Sc2pb9aehs67CuX0ZTmCLYiwGdgkIKM3jxna50VTm9lrsf4AWSXNOHM9QaqBQVVp4ay0XGmbEI3
uyIxa80tDScqt+qRAxkGg/cj+N34/zxXMFiMmUFYwJ4KX8asNMfgqkBdn0BTuU4OQ9zYLQO0wYuv
OtWTJvT8Wknm3J2cbh86k8utPe5jYz46vgRvdENqqhALhy6xZUJijyyAthAxE5zlKMK3KDJO3XGg
QM+6fw4+asXlsOLZC4xUzk+su5OM6G0URzAErncXRseoZbrcLnpNFVEn6Bdia7BNft31h+9o9Sfd
9Si+qEwLyQ1KxQlCK35TfbQzQqIqb620G03obQLBZs7Udi8DjpHIWbTpLfGbQhWRR0550gVGDEW/
INTZLWq5Mu13LHJIQ+scNeO+Lsr+7+rb071LPPGYK57ZqVL7pxTDu8ETVuzLnSf9i3OAkyAu/oDU
z0ZDnwiaa5y37o/yIo/+LiY+icRd+VkRmXTSlQJBmkRHla8uocKJdI4y9UyoUljusdWqURfxChP2
p4FU/XwO12kJUj5j43eUz9L+stcQdcYDYBwcr0BnyjSdp6WNVvRZwiDPWSzChzL/GOSTm5ttJ+Ln
xpMTNCYQUF2KSTlz/+8BYZuV1KkxVqkiFLG1gEbTGmGnlBrW/3rVsi8ZH77ypRAMBaaEgDgYQvkY
abU4qzElepT50ZTEh41i1xGvauy5gkJbe63wS6ULf2YnY3uRx1C+GhnxItMw88qSuSrSffSQNed4
XY+EAmaQd68HW38PbsDd7fhrOoYyHseZQFQE4MUwWMzePaDxrOxwdX5rz6EgYE5LhFzedtIR3JLa
kFdjaRSEh35dMwjse1Enq9oh23/kEsW3rePVTViHJt/3+CLGTarkWu+CKC5xDMOBc8YbZ76Cc9YK
/0cDsWkqJAxN3z9WdO/s1RkuVHMOoOTfwOiyekRPvulHBKV8LccdUZP27KtmQK36hjDg+nLZdz9A
sFdP2FLm/1AKzvr0sfaIfu+J/3wyaMpqCXZNbcWOgttMWnrJ470zRh2c6NOeyzm2c8K03ilDFYrZ
cz8T0bWVj3d6xp7R/JTjmyJfVISJKQsBLAXmB7hWCs2IcV6XscUmecIpPucVyjozOwMeF0PXd7XR
cYtBXrl68HyS/tFVcjnKgYIRcW5eRm4jdFyiMn5mQ5HXekr3K7SJiA/X5OlWg5isifEpFqcWNz7k
KJ/yGX+ctFS0r8UVSeOO2zQZn8o9vHw7lCPSFMtkDKYQPoI8IWmiinpxLNgyRxS10tkXajlHcO3d
DNJBxuzChGeteypT6tWjCUMEWybd2Vij2RC0vy18/ZXgWy+Gdj3CrQzOjU4uE9+UQeRDXJuddGRS
PEEeiH/nBUSa9O6Yonq/KmflEqlSyH+icf6dHi28Xb4dx85GYQocX5SEInAEbF71LGP7btksbO8t
UR3VAuRLXIXGH4kCNvCblWdMwZCY4iR2CWFyNlJnnYd0/06hZv0Gi9Pl2p+lyzfuj7PmqD/LsIZT
Det0/GjRgy8zqeYjwQ2ZSjZr+pNfcpGgI8BRk8Rlx371v8ak4n8A5A6UYlP7G/FH3N3SKxpOycOw
Rmr1V6b5/TmacDbSdPLIAtTftvVYZZ5f4B6ZkVisB4N4Iz440OQ2ctZpdzElAxYJ+uJ0qLJwa0Q8
Qa+f/w8uvAodBbSaiZ7rV29MB4aHcJKMUJBpkgE9oBjOOlA6me6FFg51uWGenpfiCCKrJWV3upb1
GQOhS6EI1xpv+SSuFyU5iLmHJF/zXbtsICewHQwUyFWgunPpT8L+DZgo/BQZi/8EAlV/a7+K0aJn
5Qh5zzuZdplIE0XVvGPR+tQzQ3rHdtfF19nqiQLslSiO60o/MsUVX+LEGJL1ghLolAY1VLcrlzcs
hXzAerGerR3fqNvu4PIlCqZX8xv/jZCUjV5l6oJI9rfDKHbEAX3N/AdRFXfzmlQ2I5MtlO0If3TE
kJzINsLsoU1thnLOTASDdJ9deriqm0fTbaPR5sziI3gxmMjVsAf2A7WDf7aO6Z+uM4SGTU9539ar
TFceCQj9uw8dDY8JkOu1kGQJcSVQOhBc90FsHzU6RGHa0YjHkyemI2jZnGs73KcdkAL16HtgMrB6
UHFy1O75slaJYDHt0OwRqXH7hEAhyNIr3JJjhvtzQOipYfnCMo8L10aN6lTpKY1pFwp6sVk2I8MR
y2n67aIKOudWiDP3MU0OHW29WwjIMPigEwwStw7K4OltTzQYhCjtlkPaLBJTNOrfXgFwyp6QHrDQ
QYZTTAkQuQAHbwdWtK8s6Ti3towLM3Lkh7im6hMwHgBz9sBihsrZ84K0kxQG5BHgWQ/HLeOmNucR
US9qQWCcNwIxYoVuEZPCfSGMq/3+ggPUGwlN7mRIshXd25ZFHRlpD6zoolu7klPpwColmY2XC/Lq
bFL8fR9QIKmDTEs+/oV0rHimlD/KL/g6mterAR3miwCKSDWCcjO6KLh9DX+Oo3CpbPMIvfs6qqCL
YTe5zedghzXY1/EEMuMloUFBVzaFkKnTGieAS6dlnOeCZ4AD69evH/l+B6+8t/3qhrT1hpd6qZlg
2AiFJMBQFK/GWkfvlcKIh8b0OOJuYTKUFJ9hfmF3CRCBwBE2sKG5aqOwO5EUacI50h/5NtrV5Vop
UVJhjjC0RzniKfCMkeSufJvvQRoCKJiYA/2Xg9IKTqz2cdVU5yFz1VyiEclihD4QufiDlpFR8FKl
z2Az5w3NuCVLqtui8RbHPYysNK+bFbi+lNNjZhtxypw3Tavi7QXpnWDFMlXV6LOnEpodl0nHGjQZ
NTNb43HboV0svcl+4SJZPCYmf7boltfO5BpnD2pGMHUGCRFomQPUXuZeQExgiGr4+PSdyWwlKP+0
2FbvYCHmmvw3KW/8FGEMVR2paMyzKdjYziUaSMBzQj4e4V99ZgLpobhbCkGyGPWz9HxfKFqwe7Dv
RE91yTxEiKcx+mpEu89dJchKfip7RauJiZ7Dd5V1DPkpv6dgAGe4Fe5KLhg51VxLdESKWA2UO0uF
2CGaoYYNSkR2x9QPdAOOVRvcYUkKBrdjCoOcwNUXRz4bCR0QBAZPYPmlJOHaWcxIskpqQdoHbsLM
PwTTGpbOyU5QZ1sBZh5l0ztLSbJY2xu6zcmyd2sT9nGvW4popom1l7l5oq9xG6wop4FT4AwES2ek
5QR6whcfqcPPwwQksLgcOOzmorUqCNalfikDSSF8ea0MeOtExCgouYb17GrREF/JgjeVLSCG+Irb
sU0ph97UFRLDGLBYSu4vRV+0YX85aTtcgmcLnG4kRmSyFEIBPs35+PWoooVI1nVSOieLbhZCg/7Y
F1NWk8gTMk/0XY3/4vzLFyU6qOpWEy4c2Qa3ogUPbBBkVHqgHzwLHvRK8ww2OJO7UFqX1hqIevO5
xY/Pjq+65F4+D3l99zWxA0ZX5l3cZFEO6c3bsXr7IpEN68bcMbx3hO2nLjlouKDWfd5v4PF1uhaw
MMVgO8rETzIWVG2r1MVu8pgSkSsmR6Jxe1S8VC9yahE7bcpclTSQm7u30Vg5Yo65mlR2MeC22DFt
7Bg8sL/SXbh9jj+3sjCc3WH6G7l0asfS5DqJcTQlcjeS/9nVcpyFFioJpAKKInjULStTqmqIJLJG
ZWTuCoKDeddJym9CQQAgcdcvG2Q/TJqS3s0Jnz1AlIszpVS6+nRvB+xj6xu+WMsigEy/t6fIzwlO
qeVz8KUg/08kOoBNZE1gJPl9lLxZoapSNMwFp0ri/0KGoviMlj/EI1EX5AHNaYmJZivH6vB5r1uB
55zWXWPBUBLjZxomaDwDPwiFHM5rSAdCdqSQTlAWJZI79yL7ONLKghcm+/3iu7q/PULFcXMLk3D4
UfeqoU9nzVMboeaVLzDAPOy2Lb7JxDUgezP/7KTHgIR/0wwZ/6mGZ1dNRAOruNHklZZhFocICNBA
rKZc9kNsYkj1Q07F7ylhPGf9U4/61671yfT6h9+I3CE4ZkRtWLCTa0PJVuG+ucrkrlMStIcT/Vw8
9zcqeFFnKwTiR3mVjX+CoKoWO3u36O2C0kv86WZe/E8pkdXcu8ejVr8sDzjnsoeE0PRcpM5h5zXz
N8ZQbvQpYgLQzn7+NqVeetBe3rvsZ4NV4oGXcNAjg80/eZE0HF6eowR20pnKLMBshttq5dbsX+qR
6LHDulwv9QMFbKAeRyRpqbyeMLU09dYmlu9AK7n9lOkumaMvoQlydhd71enMDS0vlICtpqjWTzBg
kpRv3HeU5vR64Sdl4SFq3+bRNYFr0xipc+Bl1HKeOUn5vCx5cHE3g0CZ817MaBqgO4CcRce3AxVE
+Y81+vvN24/L93ElKNUmiXHdPBNxcciMDy8QitUJUDCb9cyoCofS23jVZR+oxfDhBIRE0A1hNUls
RwJ4dBYCZ21O9z+AMXZByLHGpNvD3EEKWfwyCJpSgZ95oGW+SZOFdQTF4vY8lw9UFEds4TVDyyj8
2cGtsxZtQ6MKXHPTtXHfv3TnwtTE3FKlbYU2Rx0aPuamhjti5eiD0aqQrIkpK9drezy2jW663ih+
kyIzRMAUscEjtWPQ2fHuPBDrdxHmT5Wl1wSUctSTjHIZ5VmC4FnU/Hv2Vcwm61bOl5btOvthypja
Y3o9yKrInxZx/LkQi+gpQnist7xcMrV/Q3jIb6ExLRvIK1B8kZ2hXkp4oDKda3QdI7mdGwTNYPK8
6fEHDVXJ1BE+s4OdNZK/H/JSNsaAa/EkTGtRo8Rn8OGbvozoDw7RssHmJpsal2Uy1NM53Aw+0xS+
xnXkLTiIxr6lWMPFQtotZEM6PWLLkYjukS0spnHnYfufO1aAvR7JSKPbhmZdW6BqhwezUTD8xpbx
yRweJZejdBusXD733ecb2ZqDXfxJvblo6eGeCL77mSq/uBC0+Usq7tP8U3zZLocXgE1wctVg+NZJ
UpXavLhQM+4KHq/PtS3zqNxnAz0ySXGe8JfGQRBYKs9+KZOJpjVL3s8Zm4K+WmKb8coV7rY3ZBS4
daPCgp0z0U/bfebmSP+Y6y1tCSxgvuhT7sr25jryFXLmumYKua/yDvkAET9IH+Vm5+38dsg/Lb5/
DdlDTSYn0Be63OJUrNcFnTjLdqnKVl/weS39nFQihaI9SHJJFzyOI92+5sCSGL9N9HJ1hKrKcL9N
8StUZATymSBg34zGKAB7a7/yl9nbJ0dHlRdHQiopRXmxzfOvPVr6v8xTJW+nBElACY4b2HW/FMYJ
kO/6gGnZt+H7rgkr5ef1WOqgqC40pQFQhnlMjx3sgkLWN6ygDmrvipdoUeYiJmufi+S07WAmo+AB
IzmKF3A6LGLyzKe6kxJFC/VNcYGXRHK8u2i1jwqB6xGtCIySXWEc423tmmMFRXi7fznnWqb6bcb7
tf2RP4pSkJjerHVhb18R4cFRSV6FwtBxqCl7GqJzEyx1BI8Lmu0nWqyRzOapRfSl7VFTpGuXNlQc
dgPVK/KtlOY+IdIM9gNy+URkkkyv5se9i1iVXnWl4/iEeNDY8EIy6Xp9UXya34zCqF5Z23atkIhL
MgWsmTs7QWr1Yg+2c8w2alO4C8V5qxqUvaiglNGmqoCtOrWW3JOhUVmCMVX1ToSULybN3C5HfMyb
T7qoimpvBp3pP7DkutAXbN7SSv8r3PVD3/MqzrmbLfGvXX3nP1+Cv9vVg2CbER00f5+JhzTqHi0Z
lhl/TU+N9RnIgQ9WPCAqS4hyzrU99Y99dcDihWvfO1Rlua7YNM6hHO8dhrWpSBhHzOv2I4rwfuCN
Rs1rI+DuNYUwLpHiYEZZN/kGQYhYGOsYB0ev7HsZO95WmkWTFwts2ZkqljZX5rStwApHlk2OTdU1
SAnFNIin5kcXxfrd30OG0lq05WldlnSlFOqhU2KgR4Gy7ZfZwla6aI/QqY0V49jdFlRryh0m8L2f
4C1+aBArlBQKNDsZqI7SOQ/rrNy8KyzSsMq9C2R5YbfZJ7uCYER7GShLfC/pnYwdxxBx4o3N6vIz
slGPe+3/SgUJ8TMUmdA/j7Ctle/5Ah4Dqb1y2Nd01o68GJ9BporNoMWQbSt+udUIx5Fbu3Lx7AIU
R+DrwuqJOtsqfKmw0TJl2Jmmw1mooVHt9Z0C8OFSMEpvbf00t0t2h4L+JUZxwgQf09y00iovdz29
Tw+llnoriHMiXBd43x5ANJCtHQP8aezC9lQY/l7vmCudbL28XBzvV74+Z3iBYkI7U2hQMDfNmkVN
lu6tdh2177kpZBHrEKWpSY7TasYnEcBbHpJwTrgdT8tD38t97RTYFyOk4EFNkk2IPxX4INky7t7V
wJsIDQp1RmBrEZ3MPNcfOK4fyrIdCPm8AOuvEp5Wtm3WDZSE2FR6bvM2FiaPLUFQHFS0j1M1a+wO
3/PQkGo6ppDjJlsY0i//sAGOYyVM4a7G3Qw02l6YLv2cRpg6wNHDXDzlJ0wgd3fgAe0Mq0HzHlB+
DUIXbCv77HIJSGTCAi+oBADvSe0NapMri8SZTY0dUHXc74jzVh+RfpxGhaLyTkchftnopjvUZ3xC
gNmpE4N2k72uWQMrYEOBbFfttxS6432+LtEqbhpu0ZAlFmVTvfHtMzTZa2x3pRxBzrSUNM1+9rJi
O5AAkA20Jfs0lE8Ge+sPxpNJorz2f+nRdjDjOTupRf/9iHVM3XHo9M0NlZbkNrL7lhiXAuDEXaHk
/kXZbpEbdhfSxsH3F2NCFO8DEKK9LX5MMi1xEDtAw1ukIkqisOIPPBpIIanR01+mYrppuoRopFD5
y8Rn2wZWTDs0FrTcq7IEePxR5J3OLd3P2ya796+FjoOvwf2+0shKeQdujdBSGZyyJu7fQLXcKU9Y
8zeVQ3RLcRbYs94q3xjykDyolC35sSEnqdrCq1LOm87UVXvFij3RbHpTgO40N3d7H2YUAs0fkk36
N6zhdcLI60T87hX654hrPLevq07AZE1IPpRVQl2GBryjR8k+83NSZNy8JGLApLCdUaadK2v1Ft3P
GS5P+oq6tWrZ+x8CexOdFlblvvLVX8AW3Wc+8sabBr1VudGC3Thfut7tmPsD8z69YcTuHeMTXSUQ
dsIL1xg+cGWQJpklzVYLEBDZNr/ttA+x4U6UmSxMGaKoj5rIvpRGdaDINsY32O8DRKgTbYwzLLxt
46u44Z8DrDZrVsWHf4aS7/i7HVb3+Rxkkw3NPlKIevzAoPrKoG9IXd09uZ3ALxTl280btpcm3vUZ
6p4R91kRfP19NgIUNbHg4ClEtfa2xkF8XqAwJmzWTHr+ypW2UHDLNAJ/fnfqILHr3dlczmMZVaxF
el7BnIO0Coamonfy4Zx31UpWthXGIp1ZkqWJs/E09wMav5FtHbTjUyQpeF5B6ohrhWdhwrzQvxlc
zKD4AMwo9SD5nIqNHpCTJSpxIGLCEvTQaZCIy4en9d/VnNb4+gAHtqH7ze/meE8dKmO0sn/p1XjZ
pkt3hF5ty8eYfdX251dGIeW8P1GTdsGYjvTWto7u4lbr5KclxRjGyK4w2N7mM1mTo8qt/pgZyVEX
vfM6ONqY7xL2GORNSF1mEaEd+zvjVacKmTrS9NAGZWC431YF2UuESNt1xhSDDOj8XpzXbS3HIivI
ybzMw6JyjOFxvHUOXNUw/bedB9zgR/YKVvi66jJi0gzFagZQ1UOKuK6oTmUAsqCUnq5AycIM1h2m
iVKsOWe0mFdxq3IT1cYyTa3RSS/H5JGYP5oAtaUOtAfpHbXJXTmD2uxIHHcwjgEfQFjoIk+BTj0s
DFYB6Z254bEJe/BJoNQuY/EAOjgGOfPnw7f0dFuQ9mJjwKagvJQjQWCtnwge1IYYUOi5fAOT/bLv
NXytDdqZUCLHIkac8b8EzjsmJJnBSh7V/yRWeOxHQJtEd3q11skPt/xGJjMlu1G4bBDN76vqfoYB
7tOPpiys1qr/0lmUB5jWq0BdcXAUGKL/Y4o2N0BECYQPQ0rU3fJEcGQxTM8esEDdXkD7jaAkL4w3
vXm/CMDu+qXLBMgf5F+slRCb5JfpAOU7p1arsCgOiyu0UCikE39dYTDVDoM/0bndaEu7z7z2aEHe
FT892T+U9gZxZSYTYJ5yX5TGCGRMP2ZIEGLGOqoOuHjcjkMnDoh/72GSlxUTnqYcrqo050tiZxLo
bVQwOP2wqrqyvSlz5YabXuGqBysk57/i8AoJKHGopEykoJTb5JS165ZEBw13YtTxEG7UewkP20Ml
zN6b6eAfed9ioVIwiIcG55KW1VeAketZcI0iXd5Mv+7sj/0WJeNgKTYcxsXAzgRZRYsbcjkXDqLr
oeNbK2Pik4HYD/SvZRkLSbySHauFPa3DPNgxk4oxSmb8qwt6Hjb8G8xBRmJXQcdTSaWZMD1AIgKm
YGLSa6NbRbu3W++fysVF/KIuzb+uO2kiXMLZ+lnMx5V94lLBJkVdUANccVYTyJmd5yPLdDGAtdLU
GAQeHmZtpWP3pXjL0uWsySBjgJqE+Kc83FrqIxaMHEfd8Wc/kg5bNBIBftonqqOXT7REIU43ZB5d
QzhHC+6zEZKV+uJ4uI5XD7/UzyO4a0UUZCCnVoLzI/A2PRN7ahYEzLjU4C+EG42fL/n2G3V0ybMZ
Tsq1AyB9qTpq0kYv8wnoVSsTeXIVXsmhSceYjMarfhErjKOiOhLohsWt72ToxWPFLFBErTOcuVHJ
8ck7hHjjNgZ3+BXTfk0pRGDDGAexUWgvjLZacgNzsX2pD2jlCwhmbvLIlchPZySnrwdvNSZgs0hS
Uk7qG9GNX8ttuABN4jW3ewVqq2RkD6HVfyQpp8B/IZ2mNHIw9hxXQ3O+M4EKnJmFF+DcWVyjXaa0
Iwl47p5g9u+uKUCBI+11zWcJNfjxhOhRV7h+BuDuT77nE9c52vMUgxO+W34IfD+Mfyd+ByjXRC3i
2nuoebPV+4FN6uwRJcxy7G1+1gTWrvvq7UFZiVHALplQH8tfSKMnSoV6dUOufoR8EH71OAwUyGNT
ZeWR61HZHiMhl/aykeHumST7kjM3onjVfcmBdqej7IHgExU0KCYx9pF0wwct19M1LyzNlEvXRlJ7
To6Q26lSqH1n6xUBqGrVWCZ+Jha9yGW1CH6+VxSfeNhwoi2EHNIq3HyvCX4vLeh1eri3rnqOPKAo
lkv3p5ozEX4NZqVxeVIm9NZdKXCP3tOWLRpwuwTjb+kGiRWP1WTa6ucsTGhi3c0628R8X2/wuPl/
AvHQEj5YKPRk5uff0wLyl8hytsPQldVVxfpdwH1lJ779SZvXacQm3/PwFfF3XxBrKOxqJyk0TPpw
/lCmobNeFhSsgMKowFrwxBpOvWZgWajc3xv31+7kL6s6LSN8RXxLpEGliDadjLgv4+zWxiNd2Rxw
vrNkLwfVWfIH0h2L3zcDlQNRx9eHYjxQgUod0tlUn77nJ7iBPLGx/zRf0CM25ZQfWnzg+bJVdEiU
IalG/FK7Q1BYcY9niAzGu3yCTYuGo9/fQuY4eVv5e1f9aT49NOPVy4KTxq2Xr+Vxb5MHFEoLfI6H
39Nh0AbWGZ5iSntOZW2D7YzRyPShQsrq1xslv2mpCWEWW0qWXPiVEir19T9bBhaUQbpCQzD6sg+O
MLXbUooasf2fb4zEehJSQRP4ZH5tivdPxduQzECWZ/+vOrcEpqNPO9hC8bRZbnS8w+a0wc0o5fvk
bL1Dy8W7jzlTDl6wKtp2Fw6zxsooqszsOOWEkzpBGNDC7O/OLDo3reRsybp6zJR0tEl7etJ8sueD
zo2lqXuBqCmqtv0sMmWMoKU1xGSTxExLcCi4maAEvU2EBGTAPaAlgRwWsJlQEoRyQPOIavyAbAHK
wdsPzjiFDxvTcsGc8mhJi1GTbBcYKQE/1CYv0M3c38n1d87XhX1KHEx0SsuIg6EjcAD92tjlqTCZ
1yJePCh6JMlzVcFi6drOBgnWdCu/0N86/ZwIT7KVcTlrG1JpSdJQSUh9GIIZbDZxESU5MG4OCPg0
vkvgj1KhHSJfrUblanVA2E4ZsFsVDrOpkEeYJ1SH1/UywVEJkzCthJTUtxfkD/LZz5ppY9x37ZMG
VX03QJuiRS19D17uBb5hpORuPK16rQFnu37bXmkK8fDhuJJNkmcCThqSmspR7WZSoP6YN8gFHKdK
v1NXZ0BIWyxE21XQuxjNGFPhEeWV9zJshjRaAWEL4LFSmo6AMM0PT7rlP9IIawMeopKjSOtzGxfr
XAEpqg6P7eXgEUx4vYSxBlD9PYBWk5w2E6+1CtXT5KLYzqxFgs9ckLUTGJhjrIiOJmPBadNv45pv
rYzbcsnqLnh/jylSysSPAFaxomssU8Qax8pOmpREGytjz4bYCGfMzuHhY48f0SzhYzoywFadTJBe
EeP0m3H+sPNY82Mywz39n4QDR5rilj50eV8pKkij0CYCZp+bB5pMkgCCuQR6Tv/ADqhCFUk55wUc
CJtumeWwtuVT7vKWH7f2a87CXdRiLLX7yjVs7vFdTYlhI1vTh3pYYOwZuCEAX7Q/K2tWS6MVEXag
O/0eJgAMqkdmWCky0UbjMOOJAq0G/p2987nCCWapKnYqZqXHxY8AH5gx860ZQJGe8ngWvJbr+hQT
sT6nuf6jpP5mxPxv2TwsgXWyNQUXcdj3VnA0BxywoWLbTP9vCL5FgKSEWlclFNCy7+na6ZPLgvm4
BX1KvlIjnFIJPzTt4ShtbRIr1AFbrCZ5uVsoZEqgDKGJ3ZoRKePtkwDvrSrCYQYTsSBlpmuM5Ply
+xp01nMXrZFY7mbRWVO1aMoX1ycwNukqJck5NWhsbXzCU3w8dT5mjXu6P9xJv+GRC7plXVmLNMZv
hotIGhYMEUTGHlDtg7zf82KxUeAPWC3SbjgqMcKGSlFShoOzF9gY3pdet6j725G4Ql17jibYKb5b
S7BYjKHpWdNs0EgNzyJr63hKCI1Fzx/WjJSTVe2AmfLoYo9vj8epl7hhJP2kyfh0Y+AKS9dJ6p00
YBAEFOJWPTVRccvohmqXXiTcSJfm3W2H491SnSmxTkeZCNLDKdM76kh6UpM8kyZ/v6C+lE8CV4qw
OPinyoCUUK5E5D41TUOI1pfnFOYe3Wz/9/82eVd20XGFavKIW9VWZs/LZfrFYQ7RKXKJfbffimPe
3a8dXepj9Ao6PdwP5wymqgcfZGHYYu1HZWcbuwEpknIBELKVFqBovN4KhAXpfk7Bt+Sg8AVQwOT3
yvnkJ0jEQ7bdm+JkV8uBePpWnr0Nle6yckeemZo9omTJYu0i4ftLDnIloxbcUKn+f8u8SXFxWJzX
GlPLYCguNfY/UEor7FcpafnUj0g2bu1/iQbiiYCAZBGDJxo+Wt2kQlNKb6Q8KABqUE7rnHtKjlL2
uiumZzo0tYmzPlI3CCdIR0TVQo/vj5NOzOIEAjS3ZvVLnTqnIVEiZdms6wdCc91x8cU15V/SS4Bi
tyBS2FHnPCwEfFt9xtiMDpcB5C6xYcrPuHKKFl/cv9gCQAtjMFU9uCjPajME1H4+WA6VuMgGA5oT
mSlJU86m4vqfOMPilVQZz4AVM/4G3wt8eGRrVDRTVF1JdznqYd8mukoerW7nthvHl/fNeryEORtA
yqZ3aDYaN5ktIMjn0MfBsw3rgslJnrk7H3iU/UgOF1zs60I707EtYZJIDJhZ3JlT3u1KzFLZUMoB
3Td9yJTwiI3HPhzdbbF4LU/wpXRlKzw7yyf72Z+f+oe8G73RVCkxBswekwwuGftO+aFViB+k/KAY
c5NWbN/+UzqC3RH8wULP/d+2BGr0r6rVLQ/1ZAu6eIC15LENoH2RyEk1ribUmjSIoulWcPKltjqm
4ZDwjPxSHyqNTl30lcoKspPjiLTo/nKUpWsqh5SwQPr5+EVwQN0gmQlGqs2Z7KUTnpz44Y7infur
Tc9y0ECNT3bp0DDy5yRuINZIeX/H9j7f9yLPbqAj2WYKhIwmmwBROmru1QMbVNcWPkh1628Ni/dN
3ap1ZNv1q8CUdYRAaRfogxkBDIx0afeheSv18jxKVqJErK1EQg4UExcui8CDtIR943Ss69b1brCc
k2+mgRZB7LqMRJZq24wIqXdAcp10CYJK7UiMQRUQm+sPHNFmvChRxZ/AULa5vSKi82jZDSfUFcR/
lqOOWiE9xoVQ+eS9f4y1U7a+LE+BXONxUwNH3Fjg5Li0Lp9tF3IpT6JZ2T3uZceuPV3LL8cEDhiR
kcSOE26HuGXwIdaBZuI6KfS5ZOqBwiHtc+FjKErwfGiVCInh9xg0Zk7ckQmrkJ3a/b2A9lSG7NAt
Dq7eLOeKkvyPaFjzVN38Hs6C82Unt+Mztz20DqEU8B9rU6VGUCVRSji0ZLL1mqfhNmpyj/NphJCK
FpDtwZsd7NSUKfmyS0PXVVudyO/PqKZqV2WUYLan8i8+X14CEwz8DXz2rSpFFt6vPooKub6FAFzt
L9y4ktnafEeEt9hN8gospfT+96aI4wpuvLa0L308lIH86buld+8R3VPEd0DUxWx6ROYTEgFwkF1L
oAA3YL4kavqsecFnY6tTGwWw/nCdxhIpCwj3B/4uXhkV6Ir6auze4Xj8jj7kyKUBBoyDOAnISu4J
pfbzYBpxmcYeGcRgHuD8yTJf34bs3eyM/hLnuZBnf0GaJlpKXK0tVmJYvsWiMT2ahw0sXkBmnd1K
Bl8DGnL8dXu6VdXVpq1T5LOMM3VwqDbESv7MY0MaOo71hnEgFHkeXKRY7tWkeDiRwbizOnQ61lN3
//cC1nw2zxxU35bNAIaqk4jzgMVMXD+CcgqFREETI1zY6ByrqjGyFIdP+xer6R8maMjhcfmeESeF
WDyGZtdtKXnTA8uPGDSsRBIQWISB2w0E0OWuoM6t+PMJUPI3WtJ4g/nCMnyf6vZgW+1/hKQY3fAf
NShl65carNhKovOL9rf3gdL2Nwxeb+6t2CzSouPdF7upJaH5D7QxtJPTIC61CEvLDWYJkOUW568q
LLCEGtDeNYx/NsVFmpsySIry65qgnDp1Ylz/PKhj832rz5b73FGp3MWXSj6G6MnwcuF1WQD6EXW7
MsPVGMBKkYhvRyETfv80FkLkzQk8qTeI6ZQiRzIoOFBJ5A2cM/Ev4WmWZwtQL/8qbkeTPufsbZDZ
78GMAVA3aQ+VvECN+uDgO+i+ZWQm83p5uLoVkBIP+EYT4FNeds6W0RvYYUPZiqDSucG3UgTwR3na
8cZHZ+0udEqGNXpDZ5gA/YDiB276VToF74pNmC0liM0aIXiD/VdxhvVXm/26YOdmker+a5eKVxjN
f+D9ClA87AS5TNvRqggy3s8XSCMkrpkCxJ8M/ndQEHT1xm8POpZSz+9TMFUhDkszf5ucMfiwEjM2
lTIfhkNH5rW6Axef8zQigNnTujukoWACI4fklz9BdYZ0H/4IiuCZ5pUOE8U/8LrutI6pV3+M2ETn
ASfdAN7j3ZZthUQsSwU3ImJ+jg3bGya6ddeXrDI6BSfA/V4SdxxoKZoMVG95XYgoX+4IAOxhybFf
1i2qOGHvnbaHeGTxLd0gWlhh074syvUcM5V99PwkOtUexWOYS9H/A4rMTgSjZL5PtS22QjpNLrVb
6M9czwg49uFbzuE488eivbwoEWjLs0IA1OixmBId7Ajwqv3vU2WXy0+AJ1iDXF3xeNObKd+fg0fs
TtiZ61B48twXc2kfC9al+IE0tRDgjantMj8NSww/c0bUr2RyVVDZPKkcqhUHaQEvlPMTXAYDwNOQ
nRgZhSX4gaaHhxa0Nf9O22ObNAWMtgVNFYQjxaVP8gGmc3/7Ww0kCMV65smJ1MPBKmjDFlCVsudP
1GIbBuZ+T6Dr0eg95Uo1FrRLngNivlz3yIYmhyJlsO7fH3WpZuB/KBaD+zd7twrsZqxtE5qyLC7U
UdBkPp3mt469CPNTMBGVWijmhNgyPEFoKoig/uvD636XGLiZ3Igfs89OL8gJwhKuH9SGpbHXX0R7
oFTN0Ro/QSH5UYuVIU0TLUVP2/lTR86h6GodTrW2XyPzbWi5THdYsvmRGZ33ZcrpbE4rRP/Iuq5/
5FU4QEQA//cnNV2YyqhlAFAM+uunYKOi2EM65V9Q3eKrY7WcGZyyznd4c6D0KSDLPUFPkUB7pYeH
8dLv8FFw+NV9a+grkPYkiTt28Iek3ovWwI013DA3+7WsnBEPZQJc4/UUdGIkFa1bONfkt611znfe
5RFtFXWWg6X8trkszfekLGRexJDeCzzXjQWVmwt3zpgPf5fdDfuazxo2HtrSuzl41N9dPK431AXK
LENq0amPfN4dcXh0jU/I1bEexhLmySsJ+FIsPIMGx3iIFsREPuYFK2+ahG345l/9zhsL7zhrxHvN
aaOPFv1cmnX7ElwyApRKwjjrxC++UBO97ibk0dY37dxakF+eSQ7OseDs+0PXoJdIWT98TX0GapCG
6Kr1TV4FYc7oWdMAcu4vVpCKqc9Pg0gTX/mw5IML4OwK8dvHAGuBSA92TMA6dWZXN+Und+blXe22
9TNcuF4arfMTnfOS1+1qUs9oa/Zu8cxtF9ETz8hBtjRCRFdvfshCwlCrLIVsx/N+WG2QP2wYpdAp
vdqtzLkBv2w6sdvwHHSfPL1qUgYLazcKNJZD4Ce8HX+GhmzBPciURqaNU1+zIhvbKfVol09xu8rK
JhIDq1sImqeaj6Rht3rbmiS0gmCLXLoaR5mTrzNJcMDAYic4sbkQYcriadYK9XVdbFHgsJvk7OpS
PN4NdAFqWKDrDXuDzS/kGE+UGukmk24puedyLCH24/mua61xnPCxyOM0zUq5syVA22GrWxCBmDHT
WNISVYcxhpfDe9+XJBY/6fDXgwEsChigZ+VxFgLSfIG3GGFa0Y+4l6/Jn1tnFwRO6O9nkUDdqsRK
jy7RXhjByGDdDatQ1BHbEFw4EQb19lAYJk17UWSP+4jAVp3pr87QWtsSGLknzHZ6GzYsrGTqlQBm
qq0sENfJ3kiFq++9kqpgBWfGg4rJcFov7QVn/qv15SdJR74eQedMzMfWbqC1rsqysd1ABRajP6VC
WVV01B8+KJGGa+cZlGqlgZ0u8GyeFsmPSIAWiRCsW5cFH7vjj7Jv/tSfXoxrXP0H/aGBAweOHsiW
j0tlvsZj4KPKeMZ+W9KDTQhS8RZCt8H9yBTmV5x8kcCU2UkNJ+jSDKS4QD5trdiDNsqtO6rrFfNH
WhN7mts2qieNGcYH/DjJDFKgqEiGCORbrP5dYcxmFsY2Ji0KWrYcpRNdRBeertwrUo42oY5nFeyG
ZiNt/lTozJXzBFliQXI48B8Bl46bBK+M3Hyc8Dz71TxDW5o4L16LKvIftz8tpWyxxfHJd+zmHO0D
MLfruToPNBssOGfvv5bBRHKUt57zWm/UqSUWblUkSlAJDkRJ1FZ7Urgy6TpSSfWzzhASaBOqvPvt
kErDb7G3U5no+Ag1hFBCYskCJh3qfLbaVpQ3oIrsjiWJG4+ibvr3XdtL0kDYx4+i+BeNe8CkWP6b
KNHGh7uAj2EM2MMKG20ecVpj/3ZzKSbTWhRBoO+qI74uWgW2yBoL0pAPqfmS8+7YrBEyqhEK5XJd
Q8m4/+BR+aFvSbQz3poixAtFGFwGdX9I20ONfFtuGNIbBQQoXYN47tMtR6ls/JHpVDtyTLhmGDpJ
jE1uZS92PXfsKJajw/jRPsMByJU3hwO2bIpSwuTJbnIgIeoyjvssycvdpLJbFEORK09WZPkaIj1y
PSUWWc8HpwYNMGT+8kbVpvNDALlw7AfYnUKkSQU7r31wMqlaBs/kMpu1vHfaCGRVlAurzeid0aBs
AmpDAZMoTyg5Ixjyz2i7+qHk+tpp0TZ0gnlpIpnkyh//bZZ6NkYRHDB2Q/adiW4pJdWyIhwFA3tG
GySc116CqFsdRBJXRuC0TLpFJQjOvCmLP4PHzUzMrRseRjUpAkvQB9xhzDeMk2VSX4XSyk9F6cuN
DwAkjLS6zvh4MG2lm7AtPY2uvcV1p7dlEbKz2J7t60CI3PyLwizTWhfmspcsUIuqtK/fPTTqBUWZ
iZK5+7bQTp9MUtN2G1L7O6EAT6VPin26OUD5FIfhgdRHe63KQbz0+t8Ed6pxqIKb6mcUePrFQqDj
uNzgEHWJVZ04G8AnRK+VTQkPNAFXTj+iHacuz1j3nmxKCeJstMbAeO64iWNxJZLt0g5ftOz3ykAn
ycFXD1/Afzr4nXn+dYgVVEQYTFaP9sWFLfQ+HBa03EBKlB2ZvPNJQwTSkpJ1z49fPw1t5yvVvln2
p6JtLsyjjyvZvZjKE0JdOXBQu5aZ1iEc7blFkGqXV1D/7JUIxeM5mS87fr5pZn30Q9Cv/fS1brNL
hK9K/CVsdHxxuQwHKKcX7LS0Y8gGvKJAkOCRrCNpq2W0KOW8kWeyNdWlmeMESClANfijfVlPbmRA
zwUBiF1k589YksaVtT3XxMzMSxhqLbzDamVWxbvM51S6y5KT9LtcrIm8OAyEoiYnDwSv1TVjpk/Q
31CmOyxCQ+gT5S3seiZ/aaA98siR34JjMdoYEXAUJfwqvZO1C7fPGPXC90e7/TIZA5y6i0osN4Ok
R8AU0L8a5OaXqCsweZ5VegBFInLCzw9LyRIzqlAqz0hmRSfOlBLJ7tTERYIVzXblaxJVd4XX7E33
kFC4fmEf6I1BChyBOPf9zvUsmT2YCoe0M4kFXioPxr2nN5C1ewosPa3mIXMZDqhUVhf7UAHot6P4
dtO8KCpz3mA/KI46XvrqqmLfmQ4yhwq+fGmFEjm380Cm7FydN/EbVRYDOICRvJWyI+YBJ274lGyp
ZGz3z3iJ3SnOIGoqHfHywHly0fuCg6aCMTf7tbNguPIlDrK2Qm/nOewxRC8tQHXryOGWxp1OYNJa
RUNWAlatAvJKW/GLVhW7RxU6Epi3Bl5nlhi7On7w4UWmwQKmi0JtcluD/o0Jz7iokatyOHuYh06i
9J7VIE6MuxcT59COL7DNE/a1JRkgt1jNstWv4a1Z8lWiWreVf8yJ55EJMCWMpmCY07YKCp2PM3ai
LueDy0UjxsbxjyZOo22KpNZ94f2iZyydguG8xCCdU1NWIkFtPE+83hN6pF9URmTnYeKu+VfMd9V3
FF6JGuE6use3zo88wsDjk/i+0NvprE9QtV93AUh93I2sf8fR3iDd9gBk5zDTpV8yzCSqh/P9uQvh
eG4pOwc+orBeno7L26ANbKv7XMMU/Zjm2k2+TKd5AQfRA8jllZtDzaY9Ksad8SCWpjfSNHFCQFYq
F6nVu1zYMIgT7XRg9pnkBNkaCvpO3n9H5B+xQew+GrErUgy1IbqOCxKK1sATJ2o4+qUe2p3qMZjg
ro8lsgbbrBCDvhWATbIFOVsjTG4WZkdYqstOzrnq3OPFegCVo0w5vl2lgsXydNuR1PEJR32Biz9a
jwxoRvdW2GmNt7RIXRDkYTJNcRSRylaLO1tB/N69nX8cVSiRq4JUFpo4zZf4q2F/uZY1lHOGmyQI
Ts3QHkhKOzLzXZatD0lWABeCu31kDHw23Uk0gXbJMeqHIAIUVrV923XCwtF9PorOi9le6gj1Yq+2
wXjJ4u3b+qZrBiFgeE8vxViQFJWpWrysVi0PrD8hW2wwo0JJa101tpTsKHJ5BcQd7mNEXRo9Ibd2
AU15AHdBGC2SkhKn8sbaLbvs9AUeWzsYpXtZivq2BR8wi8e8kAX6mzliaZUM3ZIAOarLoNE9eUFg
AkSX/HB5P8Whw3c7pXfRTr28krePJX4OPxxqFoyAN3YtzY2Xq7dOAz9otDtTFnd01S56ujed3nsG
tSd6UJeyj/tQYgN96fiU27GweyWcyn/Vc9Zf+aO+tAMEv9tbhd0MsCF6lgXx4eMNrG+BKB9geocn
jOMmXtP+g8I5oubvWOwaxjvimbQnQ368FDwYWRwm9TVnj4hrjNQDLCej1j9k4Y9VfCCO9bUu64Rh
hoELm1nzYsJIk5g/w6B7GxH5vW1k1VlG9JB/QbuiSeZhgS8f998IeI+erwHVuO9cywOt8DO2qSch
qEqAsYWEBwLMDTdXmQR99h+QgupNlCCfw0wF0gwX8WBeEoD9xd6HHTmgQDPtvXKET7IiTgf1NfBF
V4IvN8Ts/SkZg1DorS/dPY3wtWzjkJNHOpTwK6NUpBZRFQudVO4HGl6TO91a8IgnbjQ+xcqcp7+P
RbLDJzwmUX9SjY7SM06NagOuiPbSGccaKqj6/Wmn/+qSz4l+zObQrmik+nzt4bUfFvcn753rw0B6
BWZ3f12sK8vRsKizDRWtIT+3YpdWyhGwrriIxxsIEk57WhqSCkDMgKleuD1XHSzD8o6xZY7tDa+F
hsFBh6mrLoNauo3J5IKmLTPTU2dNgAfhbBVa18zdyZjiualUc6G60L1vllgeP/I1JjJCYTUswjYs
zwwxmsnUWZu4SjeUU61P09FM69NMLoSK9Dic3u1u1Qga57NnLABbd4ph3yGLsd7tUCdx0YclZMUZ
6mNabGON6IGXpejRRWVe7MOX9TnUN31eQJLWxWKkr5jCFFhb6xSdkKjuVlkxN9muLRy5YH2rEpWT
Jyt+uGnaDfi+6/0rs73y3e4bcICd2ShlNXQVFpBX8fZlHac+BPiSlJ8/ecAwpKQSuOX8Yfn0mmss
ndQTXJXnjgC+D27LrxjIjBkhuJF0OZxuareYKlLMn1UGgEFmsRn3cMKM9shIsQ25Jr6blyRipHLO
6iE8PQYKC6gdiKj/o+5+bPNvOjm/gZRqwLN9/H2selAfWUAEJrbdYtq68Omrg0360sg/Rd/PQu8W
+zlT3SBOoVe23Qoe286mrF0NyixcxsIw1x00UU8AQb53iLzOf42xxffY54V/TTt1vMLBkdmQjvTh
hh+IVNNhWDoKPKoDzNQlKYg1BTrTHYuZ3CAnGnDOKuWpI6et/EwDdZ4pIaMEWE02Ntsrq7u4eskJ
GWqKmhEG87Rz2lQvsRInTdClXD736c4UfAyZZ9XWDmsvtPu1uVExTxlZI1Af0YuJTHN4GvSkTW7/
gFR/yEJs+wd+PyYIJJZJRCsgLyiddfDJDZcFWrhuCZCye5wtMLe3Dl4ZUf2WHmfExYayGTozH+Zq
k2I1adm3JgFPUiit19sx5CyD8lvZxMZRbER7Zf7DnMcM1uLCwp/XBSIwCJKAA98GthA1MWALugnJ
bHm9eIdDtBAEci2Gi8+FKL6EKt3aXU5/Q7n+0ljjC4m+yffstuBC7SSakGShGGIuJpdnc1zcJwe9
alsIDeqoM5UyQW2+i1nCZIWw/syFPlwVzJpMdHpoYqlqKGe7b0Vakelzrb1zUBA/d6/BLg3xhq4D
lDlfk21cOy+0HsZ3U+A+kuF9KU0whbdDEKjA0ModGQt0dqt8ZYp8G3LUCcxF1mFuz0iwOb7B0nVe
R7tb4RTJgVI3p3vsOkvWvZMOzW/xklBSWzcJihWNzjECqJvIlw3RBEgcEAv1Wn7r7RzhvWGgQKow
AACEWPfvrlcBQZQfL6BdGtIYayIVhWkfb68monBQVTI4NohVZrO00wtWqMfJhp9mbrmurRaa0a3j
JA5c6TMWGjlnAhCIl74rZJLE3R5JlzBTmAMVgjC7p3clUnV+JOrO0hr9aa1VGdMIW5CWyhTzuZQs
Z/KPNHIG+TBwtYKsEhB9XZGWBwjxHKd19fL3mg1E2aYeetso8Pev1nmc5JUF3t8SD+kMgBqhr0nl
qG0db6P7x5xQu/QZ19rCIVWboGCWJ7/dfarj27K+Xy0sLtyLXYMpoGLZUbEoF3WhIdD4/LszarL5
2alE4Rydna8TPD1xrNrBdZJNnj9oJ4T6PH4nidKWQ7Hk/2uB6gMGkIrCpDG+EkKcuPS53AJ8MD8y
PLSzTKRhdjdUSKN6vPYTZn5FHyUlS++J9QxM//CaNKyPRvNuSMncRM2sr1t39osuEOZaHPD8cPm0
R5BFUE0V0CUbywPkFRCeOiXi0M0mMepHJ3Wa09xohalxdRFsiVjj+dQiYaS1LgSwNMTAq1gCLRYN
pPAQqNBk9FUyeJb1xUEHA+fQchb7x/oJkh4gDYvN/3VCpCieMm6yCZOzjz5CDLu6DpHrwQrxdr3l
kTJ8p2SlUocBRy0FLgxmhFSRVcEfStaHncpjHwMSb8fUNhlq6w4ybfqqJF2GXfKSF630lMORufpP
8dlXUx5SEPSN/ZSuoUQPe7xVjp7ZLIe/nG9sS0GjobKlKuMNEB5BOYaVTf0KU3tTq26LxFN9BdDX
GtPvkyg0ztVkJiBel4mb+DepiAc7Gd/mGy6aQV7MWKtrZV6YIV5bvO63U7VJZBKEwZ16gWkcf7EM
upTzyg32sYPikja/xdrxhK1Rg0MMhDgIptuxjHmHo4H2mKWdHKljfTPjDtIG0SNXBy8bJaRCKO5I
q7pHuyTalYIRz5sRr4AvWtzFjC6vMK8JBcTXWu6qpfZwnE40ZUkkZVjEYKRf9y76lLgx/UfPVMsX
BeR85g8SvLuSZG8oroIJEkEyzOgMayfpw1ey4Hxpnugrx1U8R8+2VLAjta/G2ODiJ9HuiutbgrvR
3i0//G5pbLEZ4o6U7vEQHqWfteia5oErcv/h4uRr3FKKcCRWqV9BGOW4VCZGay4LLYYm34XY9cNx
ZLk6Jg2oGGuuMPxssplsmonAldisiyiWn3UQJRwHByHnEdFgctTj8EmM2l6vcYkuV+CHqAzaUqkb
WEXQ3lfb+vSWvgOGcZYXcnlaqMwc33neSLlpdRTrvgpesadZK6xax8npW3yirVeqh9scCxHRfIGe
+a+G8VVGxW382ed0r97osZfviXXbXa/qs+lbZY3AQqyWLqrL936NNO98lSH+7JW2QIf4jhm2xEOS
kYwERwZHu+SlXM6fePSGc2gGbtQkS8C3n1cgFLHgQctnhPp2P0Kxg+SgUuoHki9xNy34dSchcASX
mV47mzjvbu1Ct0J2klv9QJiTOYoyLyrMChsLehjiswrgSbOOdx+6rjOCaDxYw78pOs2a0PJ41Prh
YLyjqvO0nb7g5g5zG06JE5P9QDxrRTGLQNYngGQfFsabz/jw4z0MC9NDKrFSo04z2mBXHxBn8owy
Snkr7KU3z0x3vMahma51GOf93pOkPO8YYJbkXbRTeYTVzNfl6enYG86gFi08/ygGO7tNMBj4dq8I
iTL0k59qIu2i5nB/3tjY/tk6rHk75z22T3Mb2AaPXfhVWzXFFWq+JdL36RyOpQX/Hb2huF3AZQLj
I8LhyddE+IsuSu4Zp51oDamAFAhlmR7cVEpRsEzAqPAglNIUMhtDiGnu+lJt/4hs/O6EkK/LTaQJ
olS32UsFAJyFudYVuBbm4L7AlfzeJu4++LTozf9bw5IoJfEGO3mssDfUXLlLqfs4sd2tjKY110ya
OaY9I/go5z5acWYZe9l427eZO+W9XaPMxh6rTvAdcSLtAV6HcTEYOvm9F77vHvBj6kosbeNPmxvf
XIwsnGzSltjdk3YmuHqs1OQOf0M2gVIqAWGeGZ+X2U5espgTJj9sgb6kS3iBZVE3FcPlhwYMdf+q
aTourw3R1Wzrv0GY2o+MOZqA6X8ceFpIMjsWlMi2C3ly+tHaoC0ABXln6vrV4p+HC6MMxQWAic3f
vs7t7902SytcEro+2OWgGh18tz4P/jolQkWma4KwMLkV/64Sgt/xrS78udle+zbUu9JiMNPB0UJS
lGl2lm3hmbIGWKkjgN3yLPO6r1iuPnQ+N18rvRzkZTHU1JXLtgj2XxyWWvRXub3L4ZPYxIkVt6pa
K0d2rJ9uc23BznHi/Fl2RxA5aEgzWVZxtLu+05c2XUUiVN6e+FUIIDCfnMEAgOE6r/L9h0f3uHtJ
kjQxrP8KVbkhuIfZPGi1NpaEeFSFjKrvR/f6AcSlTkwfK3kKvNHSCe3E1KEezNEf7d/94KS5slGy
mg9M0rNJMg0n2GL0h/+wqdFe+StyZhCGaX1Wz0QNoeppJY7ABh1UwPpNdlloIJVFVV6qCz1Rz7ku
eXp2ubHz7OmI/WpW0cMdqPnwLbUgh+iWKge/7WTMKIpOkwrafCpDni0bn3Fv22gEEAESRa4WYQB9
UgPBOmLsdzA+cebccoV/PtE2UmiVWY7ODgqqwDSuLd7LoHN21LLtx0ebRFMKs/84rbmZ3r6tXD+l
k4TmA2GaNvBRS+dovvt2wURaOd1G0b9/XI48AECJ7wcMTEt65rlEZXog00G7onC/dwz83asPmYut
QrRIy6Htv5FNOqUzzipSxenM1a3L49s3l61WWBlL10zMXpLydBbdF6LFJTL0htZb+yM+Siif7dmS
lcQE5qXCx6qvrJCpX10CR2mDM+2GRDoTe143/NkAJEHXKVk9FLyNmtLKa5z7F3K8JBZC21jQ8vV0
v0B46tU0ckRemi5aGwNB1FpeaLE+HodHFXXjPxVuSrZScW+hyHPVfq2fnxr07bJKajyPaUzZlsyO
xHnH8vjwQqfH/6apTqP3enzIlGjBNlR0ZQ71kRmEFidf6AB4+WaB98QLmmLIFR7iNHDqHJCodwva
fQdoTi/jmRuKprFmoonK+RXvB60El2TbWH9/TZm2MbN8fxgpiK0JXB/TYe0ziCgKHhbVOw3Cvpc1
A2iWUecUdwGaxvzkgsgchpBjudnmpyJxN6xl9UupNOvwKFoQa9TQUbn2vcavAQIjYdTllKYMhTgR
J+wfDE5n0TnpHVngQ82uCZ017Q/5UV/uj+Sd7Du17rQidcLWAXRqlCgwRF3tCCYGSStfXHVsbb0u
N5y6EOaNGLa6mYsUang3lVleZ5JjMA6ajGmZh6iG+vKlqBMfmOb8IkmUbsn65bQT4r6tIBRdlfk1
vihOWcqEVxATl4otSoJSjvxLdxOr3xWOBkli6JuZqzci+DeqaFlmuyTQVHzw7u0cZQcsppDRdPXC
VOnEiiznZvyQTF18SPAsI6veyLqMighjZlal1ynSzIkJwIdKvk4O+QOtj/GvR/zLRi2NLlfmZWwp
5PVE8csNuvwamlmttAirmaagb17PGQDoHideYo1hqJNduUAHn5btXE7ZvbDlcvRwp9UPp+wZd5Xb
p55X1vcG1vmzwBCPhEWi6KUEo4MOAaXtkDI1zR5yuB7ahysjp0iGz4BIgffSSJ9KqNPje0nji0jc
xlU16jD6hiJgdgcO2MwTv7CTt/n88HnKrRBNsoQ4qN3UXpHW7KfNqSnwg1SdWMDxMptZY4ya6Fw3
PdQHVU+872LGGM0uswieOhYWKzt6RUZZuk/JwuQiFdmNh854Mwt35NCXRFk40XXK32Qwqp4W6pOz
+z9Dr3SnSXqptQJvXfb+LQotwl+X1uhWja27nDsErG7EJ8Vr7XOeMgMF/WVnQedVEt7r+0rvwckb
ZmymGVRJ8NvRevuqvCiE1p448UzX2CPkfJYkLF1AtjdhvLlfi3jrSJah8jc4gicKLjLL8lh8JFMn
IL36AZOoEdKA5ww8ststPryWy29IW1W3cOsibZz+2J6kxt7sephE1zuaYT2Rzt84itGV3qm9fPx6
y+6A5mzFMuK2Vkrn8LHDgZz40hDSo94uFpfTiVW+7E+4OzslOYqOIXVy1Bw20bVU82CmFAWEI//v
hPazN/QXNOLb7fRSYGUBeC1RBRca+TJMLGOYDOWdeQ/GHnsfh0PWc7iBtmnWiVksA+vCfYBM5ytK
uz6j50C+JhHeiJleSsjSr8P2aRS1Ezc9bVq5Y6EKoUiTFBJd0iyW2NPPu1y+cGmdu5Lc0Uwankma
rgaTfsfvhNgMBz7KjcLRQtUjeXcM/6LI/SvOXWQyY5379DsAh2fX7ihP0hhyiOMl0np15M166x39
3nJPo+2XNJErb500ILJHgftuzJDjtpYhFAq9yesvnHsxEAdBU/iiPVrhmKgXqbOsgdvU0RHX+/+u
w1kaz6SKCTnFQO5pjU7MV+toGyvCf3PjIw4t6r1DFayaHcmGDE0RlEAQTRf3Mt8G2FlLWsSb9TMi
dVM+8H/gMM6XEKIr4aG3u9Ptb1JkVszzh2nAD0yOeyHwgEGM8magvA1UgOoRxPHIaaLCeV6rqYop
7RVYnfq4kgFKrlnGXMEiVJF48FOSoBqtzkhnq9n6oDxV0tDU0cvxm/S+r0Z6AnIK3ya9jxg5Ht92
rsOzBtDPrcDurR2cduty/DIT0bDfXY9yFOuo8qSo+n6sawFMt7OZ/j3MFKaj5/D5EQDupC6A2WcP
SP2+Z63+4XNQ+kH3zxGqqrVyo6NrnFCerOd5mXBL7zKPtiZhx18l6Jyl8kxTLnagg8dSgIEqxTMp
FksfaakdqhaJ9Wy0j6/DbAJBSza4TfV+g3D/V2EpRVDeiDsrE0cse3Dhnd6FLFCmSSufiRhpqXAa
VHL1FBHrfXPy7MivvY2hFnVihQyfhTY1R+YFNkzIC7YzgxNAchJ8dotkH5y9fvtWBEdN/9EupZ/L
p8N70G4lR58tiFCAotk96g15ZTXHe1cEo3jVs22yUTJVVoCCTKeM6SYf9rjRBpuZY3H1o8Ku4A4x
h0xZYbijZmyQmRatZX+yiHGztZrA5zY8TKwwpJc1WC6hOULNx3g03N1X1dudQBgWq5hkq4uiuq/z
p4laAW/uRAHPjwaoOesT07eiAuPJrFob6b6ynZtoUzz+JNXfl8R29wyg1orVfAEv82oPxWv0igrN
qJRhcshzgZOjsr1n3gZ42NJNQi86GZsVVyObbTf8ZeNrHPg3X9ECwmW/+fe9GriLzdL1ajUtUlje
8I2bpW83DDRS1wDv5z/ImAhteDIzrmhn8yw8EvfA6dVY5G0vLWUGljcR1ygCxUO6D3JV0KuIPqDl
dVprqM2m/LomKLtx2cb/DNAKtLpLoZY+DgtiWf6ncTXkDzQebBi8ijfaqdxIIPYuC+pAZVR78Uch
dlNUiOnFaWHI3EMvseglZ13C4Ux2xo6kF6Mwcx8l0akF8b7TpMONlLLcsyXoBMDiJAyqUmU0gWTx
E8btFnNfZC5n+nAMzbdegDu4xe+zVP/IpeINNFm8sZOUvW+roE/Jb19pXNkIwchK9LlV0kdeEWiJ
OAbJnbY/EUKvWFG/2Z7c5kRtt8YJmcb8S+C7ta9Q6ahz3Mr15Kr05vhOg4U44YR0FKgHZe6/Vjyp
miRwqUbDhlpJFjh+LiInIhreGauYXL/pIfbEXWJ4GYVitiOBO60NT6JgYfGztllpfEo6Bf1J5H2Z
Pz2ltAByyqu/gXGqInC2J0OmeVXv2q0wGN64WPoIXQgEVW5BKn6HqYJJ8wWZgIYjajPu4Tc4TKsW
U+1g3RiA2swSyAWS6EGpOsLHEn0gBGVWjInoo1grjKY/EGR3xGO6o7fgd4pCFRArKOITb6Nfuac0
2uOKnoXr6iRaTfbBIa8ZIneVhgjMByIMAAaHq/fmm5TZ125Xzdsvq7x84xGGwHQ1u4ChxEtUcUJ7
y0vrCTivqG9HuKvh/+fhecgtsar9tEQeVnVo6p1wp9ha3CvOz5WHkJ1wSCBgZEMjRDn9slFFCXUT
lAHE+YZd30QWUx6kiZiv0CHnOUI6e0yXRxBNxUg9ehcedRAPOxuuULlHofZLL7yIvPCqeQ15ykXm
koTnk43XsKMCWL4dkpE52j7LYDoPgIRcjL/ZhdMgdg3x9IQuwctUmQSTNmjetzzUCiwa+Fv1tS7N
KwyYPS5NSPfbSsb/YZUWO+mN9oPR3cW8lnp0Mh5NiOGhF3l6oeLq+L24g2vvcqYIvP8J4BVaS8IL
/bF/qaa80+CrLj8A48n9Pgo+YHc2qcNg6ackYpCEYI7W0xYy/kpzOsU3QcnEjvlZuE91vdVCnswR
HR2LHyGN7EgdIZ9UhfqmB4R/IdGGI9YtARoBAvsnnDBUlj6SICfdo/KIdOQTaQBd8fHpAfgqNIFV
ii/FH+qg3CJ68CNjSFvidgwE5acqLydk/pNb1lPYB3HbT4AtGxUByNzwlIVqAvgc8JefxKQBoj1+
0SnNLxaP+WdxNkTYnE9KPvTYAXwHfAwCnSBOBnvrZj92VWb3BDWnQtFuTWS7iSNwLyjyF+1n23wF
+dQ/CvP4kruWHH15oxdhFJg6cZwCRW/3SPjewb4nDiZzJDcBUxtmTV7Yw0EkpgeuqvHZbZFGpl2w
GYnDsW8EGh0RGW/iCNMJWStOJMCUZSiW5xSx3MWqLfBjMlM/EJmI9LbzBhe7/CCJVNKJjjkoJKWS
GQSpjzwSKmscqYLtS/mwImc+9nMc2rglH/O2AC8JIN5IrdjTMj/tUYyAPoa4qqLNAr9NKEooAvR9
2dZcse/TuSDGgACFW5Z/1nj9kD5W1JRXdEi2/8qtRfTcYX5QjVb3e9jAIVusXkMmdkmkgbYduHem
sHTqIDPudm7uHxVWNJb3N6KmAxTABx7NpHa44iHuK9wTQ4QXo5UgY8yiPMz+gKI/U7rzDTse/1cd
nIoN+a00v7AgeuyFjNG/fRHa57UcGZMRnNIxpY2yr8ncM8RO4lQCNAGrDgSxJ7ns+r61tvqVjZLm
IgShXX/fTWgytgkOaTAzr5JHeeT88ig9YBE+spAnmlSxiwihKc9xniM0qZjBcxIBNYuS1Cx6DACw
XdxJcWyfY6Cglo0CUE0NlWEjg0qJ8dj7p1Gly2F1lSOkzN1xBDW++bePFxb6xHMJOo++elV31j4q
BZbBnk8v1Dpus4xZp2d6XfqYBxODRoTo1xwsgz1JXrAiSWx9f1uN65TlcAE2dLHm4SgsVC7qFepl
ma8itEEYx/GpA5TwYDYIYr7D+/zd4xt2XZdjPM9FWt0qIKXTxR0MKOtmPIMVxQ2bpuaXzCIO/eKt
sivmKJIvbhZdXgzT4wHTQ5+XeCOAZKuYTsHRgVUBhdYRremKoL0sY2u4Z5wPC45QE6BP7tPch0SE
ur3vIf0PEGDMDGYLxqbkydUeIaiN9XxmPS0D6NPsk3DaReInums0x72zB4pMqkBM1zpBcUbOtcHO
xkMPEZbwKk5JS9R91JbfaYXDYCYJgjG971hfVP9CuYorb7Xe/6pyHk/Vyrcjem7yfZ7krA1UzN0J
yHlYj5QRufvgtg1kKs/POczcH4KefxzIzK1kaPI+iCIBJIQLH31BzzBDf9KoswsISZdwmZFc34e1
eRI0JJ/alznhEBVUu5FbafS8OCOta7rA3JS8Bntl+kbStXai2yMfOFbvlI1DYdsCKnZDj6XSZfTQ
YZ8UbzdYGWyAvqwxYJiw07ykaaH9Q2sfKvGZPthJ6304h/CogQxZT1WJLWPz71A4YQJkVbs9tqbf
Olumk7gyV+e8ZH0OHFob2WtRJcKR+w/Wfl0QSTHtbC1VQ63G6Kq5mDAGYheIJSDePlY6hkHgQh27
q2mIgFNJJxn/fGXJ9sHYYxNhqYKdApucUUekxTP/g/wZ8y5PlaQjrK6hssUIzsOzRkmtA4tHfaIq
B8PxvYc7ndmtSUvMgGinkCWaynkXnBxZfnRCRYEUzCpw2+c7xqznrcdcgbYIPb0ijd6Isi+vjBrJ
ki5N/aTagWPAF4cpSF3gKxyFaN5XXYCAXoofAmbHHqcSeWlUOqO7MDNJwtu4ZGUoHe7q+ATBAZoL
dDCi32F7AU7QvcgP/Bi+bJmQmV040xe5gGtT6R6X2DOczO6K6vNv73sXqgnBPCKiPt4fqviU21Hl
nzQLFtIq/QutEe31eTTJ/9xrzMnWYs8Z01tEvQb/26Bm7D71JFfctT1x2MtGxx1Ilg5MkRiCbbvU
Z7TOIyC/aUjsgGpG8ygfg5NKDjDzx+I/BXJONh9Mx+iT8j36VjsiiQyAR9njDwe0QnCE2J382Id+
Q+XIFRU6riu3NUqZyY8KhBUnPMgwEExoh6eF2rWLclF+eZOafL8EGh4gHdAE26bQmVvjuf3qTPj8
IY0O3u99RRSKpTgJjTiqdRRgziFywi9C/M80T9dqaMNr9uZDqV1UAzK0nq19Vd8vQCYhjezbYOLT
/ow7fQvAsqtJ0ohbrFbDtkbaB0WysK1lX64aA7ModzVhZKnBeYJbFLR6oxwoKUQoQAQAPQjNfAim
xet9yZRXvvz0BgwXyzu2Hm1R4tTjwFqhiypwfNyCw3MCNABtup42f14UcvE7nAf1phcyCNOYYJxP
sorSLM1VcfWPnokQRuNkm8GsBPRAlyJdg7cas7T1ydX5zNtVu/WhB6IincfqHM+InD0jyEgbx3Iv
Xk73UuPFlNgzXM+Pin23Z9WKzPh5x/0IWLESRsA6uzf+CzOSQYWSPmG2OVbvyM8hU74mKxQjnWgX
OsR+jDZmCWY82sADx/KGcMvC4mF1yBRME8cNB7ik22t7A3I9VtrGQix+o+wTNuh/9HVMI5wXnb6e
cgbrFyg1PVIaH0G4qIxhg88B2R6SB1n/s+p8yyYR3JETupBy0PonzS92XlUKG7OBPWqm8bDNDDFi
qpEsF71GCTU9eQ9duClx5yh0xiD3lrYHEHVOIvwAzTJ4xu198NIE2QBdKLZZyzx0dovGIqx4qjNq
DwnaJ/oYrbRnwotWdecOW7pSkouLh3gn2NcTAPvY3GOZ+TEc970e9PizMOgHgaSBcG9EvIMTsf1l
gTMIy63PKz4Tj7B3i0TSVkrHvUnfpQ9zA3OMTXUkHsffbLLrENXehxUV2WkSuOF9RLm4fW10kGdi
yCikyKqPyEk6fSzx/+rIItNLkcSmayJmNp1B2rEwWnx0aM3AxVPk+dSarSs02mvEROHTosFx1OVq
eVlIqwQLHOVkjbsbb5ez4zCRwCk7Fw0z/vUnr1N4oXoZVw//Ps5xPp6ikdtD8/YqMgs6mWsrTlYD
Y7j1IcJR0AsvZyih+XEwYN34jAsKPQWkp/1eMD31H5lhduUZBSqW/ObYBYwElyLQFTQGKFkKtFOO
Pkjt7rYIe9B/aZ9gtSNRaFHR1ogcIUJHizMPJ3XgKPuCiZssg0DU7dQTZBGEDr/cl9K6wg8ixPjE
Z3+2S6tyM6Wdex+PeE5kqecRi1vbT5QdftpUTITzFoQrE0oNO46q04vmf9WRD0/h8TtMYKiKHNuh
dXi9uR6FHvNVO45oKX2RAaYZ5m/zRELn7xTC1oqUmLTUt6LhXNOzUN65+9ium+u6Qn3VOAFbOk2I
k0jimoARxjipHj/Z6crjme0FLSTgJIvN+3N8L+3k9n2eY2He/9aw5bXJ9iY5Dq3OonYYkiogV6mx
oyky7pnDjkbO7PqoLUnSJmNs3yAKmcccZHAaMMCDCoSlaRHWJnSxvJhpaYCPVODp3h4RfYrNCBio
L+SMSR7qoYxtbb5tn6N6Ln6n+dSbWzZs3A4RVOfxklsuO31eI9sWk+YQCR836mStNW5+ibXRPL8Q
LBZMCaVCDZKIgmBKw4xzxODfIdJbDdZLKH882PSUS+6nfZIi+ymk89r538UqvdhiFUAC/R43aX+K
GaIcKI3Zdybd4VKpcmPR0UMB8VUswe8u3nNIHN40uoATwAGss3kF5zdH2lZnt6o+HvBv2IpJgvhS
RQ3LYox/y7gE00+7McfkCqCKcarW8ExN1Mp2RBLZFLh80FwdNX7ZzSZ2OOKtExasvra4Mi4tjYRT
UD9wT5D5IuA/M3Jet4q9lB++cCpjizd/8oa/vQW2EaOLQ6k+RFhr7+I5+uKk2spgAwPzwb7ObYP4
hD8g22XiAbcUyrBQKfYq1yvPDrz0ZfiVa+pDhSIjOs5U6WupWc16Ma6dAZclUSNEBI8Lsy7iltCx
j0VIIXteG9MJLKLeT1XlPFNvc6I+nZF+in82duIYw5waoV79WunrQnkVgK1Ibd69XnIUIQmTyCLa
6sMdOov7Wp87ljqkbbYqzcfQTzJpyuyFNgI8WN8Fj4czHjlCxXA7pCasSVFVJ4OevCs5n4VRjX9Q
YKO1hoz9+9uq25UlHbun+RAc9fD5oEZL7nFaq/+azXfcgqm2Min20xRPZ+/oj4QfUqoUCrNftlTC
CyWf5E/blS6RfNFo9hf2dFrnDZRwg+/tH8juHo2ggW5z95F6Nj0OD5H3vpebi53IxeuMxb3IM3Aw
Rt081nPV30ZxmwFDvKKKc75bl6RIf2S6QBTRyCrghRYFg0Q8NDMHqeZG+i144Jc59xX0Hk8ZjXVZ
YGq0vdzcqJ760/zqzOrGAN9w0KihNJqlKaPBJsk/F70ib0CEo8jlUDvzqKokxulTl9KmN1LDvMCL
88txZcTV6Gcb0OEQlnsvT9Qe8+SopPcFGW5uB3CSDpi3O427B5xDsO7QfakYUbHMQYP5A9mcSwBy
fQmw4K43QhifSx8RZaakyN4PxMVZQJlO5AJakFgDbWDrwP+62ir2qg9x9qoXqbej523b9nXeHHA0
/NsLDx4qH5c8HEnA3bmcGvo49P/mbzwT1pqMfVqiC2GLk490wcr09Kn2a/SWxq5Jkj0qHwREdbd+
MPox3j2lL6JmNSA0a4KVFqv3ymPEc6pNrD0bHkT9btUDaiZd65QNaCI8zle3mO8RvNWVjwB7/98w
yvvzTJrWDT646fiyDXthZrO4w8KPJ6YHoRL2c5J7vsLhDXe5vQFzcXA96LOF4nPLiFCpuaPE74xb
72kpkaO0rMyWnBARvha78tQt3vpynhO7PzPzWtbdCscRXu73lSKBznXmqC1Fp4TIJVUcjmlXgrO8
MSAG7VkfPUaju7IPXCv4bjZbk7nzDIbdIu9hx13VADJu8pR6WT/F5fc2UkJqxNMJOFVhjJKep2qR
NuHBAfOdwUpIIR4SJaiHpt/qBtONy5YW/sKLfqUuqMwwG5CnexA9opzR5EBXNOX4tjr4qLuOPkUF
ntHHVlqMwoFjy/3BOxNjqcVX16RqDkXaKSHUHRKZXQu9K5cqVSeBXHtGYcZhECShhiF+OIqW+xHx
cpErkv9ROBwoUkCem8ilfjwvqZKDrMhR75/Ommz20kLLNlBX7Z3aC5/5i+AeGgEuUmG0/BDVTJsu
smH5R9ppiViZnD8hqbw1SvUaHg9HFnhxMVVL10U5x3LZYcvpePJ5+UW4ZplL/1GDp1F6UgJYUo46
SYo0E5q4kZlPPwOgYAjLNJovGYvKbufNgHq6e6i3sbUK7IxIhMT6LvUI82tG1BNmq2P8Kpl2OMhn
Hp1ZSEgX8ri3r9C0fKJ6K9eAkU/eHNT+vGjcI7jNouKaZrKIK5tOBbw8qup9DlzESKhhvByckqUF
6oaVapLfSV/Hh4qkmoPIeWoJBOf8DUG66ydN2RKnVcg7piKNDIFedn1gk7do8YKi+jWDvlCwnM1I
7x1Z56ZE3WoyqtEDhqEbitOA4PcvmfIgdFiMlXvMN12K70/eLHqA5JsF+AA4c+DbhZYLJLaQL49b
x1iAlgoM7yWS9XRODRWKofi4q5oS2OEpY7MK6ij6MoYpdtfaQqGjBxzc+Ye0ksXLZVEKb/hsQckD
8S82IUaWqI4gBpCBwmkjMFiWGzPaU6DAa5NyNkgyDpVJUFDihC/h8SzD3V6K3MXwM6yoWj1LMWku
cemlyu7uKS9Mw2Pwd9VvBov8Ae03nsGoO2lTIdcGrh15eZCfpIMQ3WvTYJ0Jgda/UDLsnjPhWzEn
XTR5simgW4jf//7219KUGeOOp2ihn88VSEo1bKfzzG0SMkCf0+1eLspNgHJPpge6mdazrH0TM/kq
fwKW1krA3lGL1ZJJn1tbsmgb48phuxyhCsU8CQ5CYmgGN9C8P0rv0ThUs0Ns06UZW7oKqXQ5bYwL
NFMteYi1Qw19/AF6AN0TZ0o53R/+zueejd18MnAwXWffCLctzNven7XzEJzw8hjhK10LxgT2cQq0
ZpqPFg5KAwVWJzJH34BGHXXMyK9bD4mrnE/fB2RNulJDGuuxcMojDmnAs5kBc5Z+UXIzeS94PHaH
gNaeui9ZD2YeRkDO6lUHVsXojacFlt0OcMZ6m+cYk2tWZ5+w+F0DqHNbAa3e0rDPrwqVaB3/h0cS
g6VfQKfZ4S9qQbQARFQ/xcSVKR/1Q5nl/soY/b/tT87OteKGgA5VKkinjb8HInXPYzihCfc34mpF
jICb8JtWT++xUWmAZn3lKcWY3WEq+12NVju/o7RdtTFpXDFv/6YRcfJdEzasyFPXvHfAdQWyYXJV
eeIawS63xJrqbYuyjZ/v/pMW3jSHNGDr4rOCij8+fhwC9zMr3MfK8GiCEW/As/GOp00BjwR6OkFL
E8DwhYH2F1TTCa7xiM9c/i7HrLanLwJm/qSYUFpQwU/fK+Ei0v+6Tm/ssJ2bzhRGYFfsyoGSVoaf
qe+nhRh+kBYuAdc/loARB8XQ5DYYZIh0D4Wk2MiUOi5b68KGHOR9krJveVuPajbUC+98PcYihO31
Du8qYvuUKbz/ncPxgm79h/kjnfN99WdI8fHlEtpPCCUJmlH2xiN+mJ0WSk/8TyXFutNV94zWu1hA
6MugrA7ucpZmuFdrDrUD6IRbcIUsb6EPdV5hwOK8ChfzKazdiN7nvuEzzN1XR/Ly16SblPaQK2n+
u0BGkPUIzsWSqzJFvwbzUFDMSGf5yH0NLGeQKZBRM8QBIJT1qpHTOhqMdDjsAFGhqXmm1Uv8K8c+
0FAqbWV5Yf8WjMmLGzNavlKMTXaBb8ciLqLYwHF8YOgPuoeUsipIfkZB1srLTRhiq01HEk1Lf0IH
L0l1FuAx63efSU6gwZ4mYU0LeembG7DbFH1QIJ1yptYqALXSgvGLgOcI3BwsEDRtJ6Djn5ft4Rif
CY6cAnnXpVm1/CVuywVaxjtMn4JMrJhT4gg/jQAmcejcRdUIXzUE+hgrZ2EvDzq/hup1sYfGf5MS
dRSL/fFbOXkUdIUUzU+MuKRN7zK0c+lX/fjVX88ZYplpckP8RItSm+0Y8JAuBpLXTNQ3r053I24n
UN8l2NB2pVmt5s7gMri9mCNOGzzS6yD3RvmFd8YC/KoJ+s2AsYzZRRsZIx0bUHH4ekmlCWlW0/8B
zCqkFBsH7dkS6JxAYXEz3UWol0ZwfCdnmiu9crLpDJ6YP45FvGQRg3Q4m7lXHSe3iVrfEpwm6RTt
offIQcHh4papxaLR47+CbWh5JphTI2NHkBBS1BTt/8ATeSc3QM4JsN5K4Xy73YLxb0KZXvuhDmcr
t3m5AGtMqTiOHgfwXs2Kg1024nZvuFfxH7boMLJHAe7f4M1AG6+lMNWU0GeROp3uBy433wrlAw7C
zS+73xLi/t9Rafg/78am1T+pzBbqVGUSqzvUbW/4g+DQC09Z8E9Kbm+tbt1X3qPqZdfGKaLYtI4U
jadagX1UpbdglFByajsPnFqTqMUpflQ+P3DcS9eF39hzi9LAN4YrNc71fNRA9ysNfHm1JNvW6Tyb
RbjeULK9DwXOan3wuC+24LEUlUM6sSQL8CItCbIN0uVkRv0L3TbyUKXtQD0Kqi2PEktSfXmeRuD+
m2j4I389kPrLy7Kjb1mr7TmAFww7iwDzdEW6FDHk2DzR0adiMm4h7QHi0f0h35YXIlbmmfoLzsEs
I9ipy/vX/OK8PC4kTWFplmfhNHDkjmkx7li4uz34XKIcOSRrD3UMXv8jmkseH/HljgQy3XGKv+Iu
5X0ZXPygGYBxv48xqC73gk0aSDmkZDb5GsflG7g+eO3AzctkJVrTTUlkvqP9jg1KJ8HtcOX+qEdp
n+aLbnT/hG1Onj+e7ikXzbv08If9yHKzuRejpoqhcBifldLzob2ROkLPgIBJx9M/0efysAG/bZ3m
IgX2LSDltDgpEO+7wl1DFqZBe+sdfd0LshbBhhpsuwsMtiCjroYkJ30d4DoFaLy9M4rdGyWSF6Eb
H08gm1iU4qdw8h6ndXIEOpf/D+cZIhL08HU0axIiRLyuk4Rb5DyEN5fxs3vaS1oGo4ceRzBzfx7S
A8Z1qZ6kXl9iY0w8fUmU4HsAQK4sZb4dWguLM62aQlzipVa/EpTTyLsKPmaST5nEhqZIhsD8TGIO
+wgCfHt81LeIMy+H9LBt/zNGnBDSrdKxRj/Ue8tguGkis6pVPFpWnKlW5Im66pYyneAuvt5SzvR+
3Wsm7rC4jfOr4aseGCtpRhPiXPNX2YD3XSRD7RzOVaIwQOWB8VgrWdcHtYFMfbhR42PXwlI38cmw
/B2KDxtrdU5fViSFwvI2fTc5YKUtgM0Py+jijibx5et07LaOKUOhEAiuqYGfTIMLTKS5UywOXF8P
obIt1OjdNDVwym+RuSI2Em6F04vZXgQaPYeWUALycCQKupFVLa5YQpO7+MRL5YpafoYJfaI1VDgR
jXSfF1vPnLYHDOGsm/w6PseUxshwOVMu/tmsy6l4a0JyFPW1lbB8EOATrS5/NpS96jmdqtxZy9lF
jjDYvGJe+/Ml8x+JLvrNZKM6daeMwPvuZxyqtrrXGHgl3ypn6HQhsIO/hwshYgAaDuNuI5rwJEIT
7VRnqy3E8yPuhX17WsZEVkYVP+ZTXYQ2qV57T3fCKW3cN8MHmXTNFw2Th8/OYXkL8l8UsLxFttTK
I0EhEuGjRR74dETpTGPd6rpwXZrby9kar9UJHmLxp/TCwCgr4x+WDYdPKO8ZRPEk8bD6c34nXLME
AzMLPrU8MASbX+Drhb75nizxvyKVwhB44f/sLCcqX0tgxsG73APtFJe4Jwrg0faDVdLfDQVLAYlb
cqOp8YMUQ/9psIpRaqn8sM9H45cLD36BfNUYdGISe4HBhE7fmbwX04XW3VaA92urOGNJntmjf7d0
ddPftGS2x4Dym64L+X7rX3PgcVILcrkffECYrQ63o6A2gO2gyyjqnf/xlWEEQobpiGTqBNJ46XJW
qD+WXUxk7E/jfrzchyhYi5V50oVROBplAWTnMxdRl1070O9tPz5of0ZbVM0sG2xELmM74O/Glsgh
f/LEkp8lidKwSxjSJekQvkCs9oAFBxGFNEnYUE4W+Fohf7dSpc4S+EHetmG9f3+fp2vbyCSsg+ji
WDyuPikhyTC48rd9RFqSsYYCWOuk61XxWjmNEpOD/FmU7tVrAgjNbPg6UbbdRDADWLjbcR4f9+oU
s24Pr/2uxEj6VakbScqos7Ppcz9ULZE9McIMrWkGh4V1r4ax55X3iFDp0Tnyhk3VuFce4JKgqOR7
m3vvtJ7IaqckV83Iq0+RZWlE4ffTXQ8Uk/1tHoRgt7XINVgrCZKpfb4t26ZHeECBrYhSgw//wUab
dW7Z6FIz056wLjXnPnNR2ZPdw/f4+AF61kdTM7EGyR2gvmoW/r1otvNQaq1nxkw9Jzx22KM/bCqn
bBNFwwZ2aX4hRxZvTGOm+CPYaltb2BDtlVkeDKU/2JHjGdiucB3kzjVOApTeliWp1jzeBkqhNkDG
pvXyxt/no801hyvqbgELx0n4vNfzk2KtkYweu2zITYXss3ItWYGRCk9A+wzzmFc+elRuGUPA3ONw
St1TUyXJsh+2GtbhNOSCpEGXf0GDJTZRp1GJTor+st15wGxvp516WnLM3zab82yl1JlGOxTVxDqQ
ghdn9qKyOvEU5DOWVa7FXgRQtwTYzcvFoH5CpMm8VFXgrEME6z/j9qI6218Bs4A2TciOytKfBzdL
X50Xhb0DRJsaqc5MorFO7VV6v+9Xod2Z6utGmYC5M1gjOnmAau/74KYNj/qT3ZcZDcvsS97NcJOc
Oh/rdBTKl+n/pq/qEiHotWNoJwgDVeSufLFXIQRv6giM9f9e7APv6ve/CfL6OyOvCY8IGShFuv9M
RCHanexYXNOt6IJifzYgMoB+L6ZTeF3v/HHKxKgMz6XViQPu+uX1GuuAXkkEe0p5aXBKc0WOadqK
LiHI/6vZipvLVmlqRC72IVFMui9myDE12zf2yWTLsQtEKSYo4BYx74aoJ3012P+FI17KhyPGypqA
JyKeEpaYS+qczfcwx/YlgzkE5GLQfZI4b85VNvfA2IxV22i8K0Onwoft6tkppOquDpmS89H7PYHk
UbhRFEfWXnUb6mObApjqxzcEF/MUCL79XaxEDL4bodPHYRMI9+sx5G0DJtFLsJ2RXLy1jfuQijCY
PmYIIzn1I+zJfz38xNgQqsj/3oGGcuP8DQJ3DVAUDEFboHIrtmv8JMGsDa/Q5Mp8yAK6pvzYvo0l
STKDbGqbYrm1PZJn7NdM5+KSh5uSZd2qebT+7XA1DbgjATOsxZmjAwZ5kDDvvdP7gOLG6sO1zq1F
7CtTNAvzMAgrvuD7aZyEX92LhlvLNSec102SoIKnUK+bDlABWIc5JDS/gk02Taw6aZq6NjDfgpwr
vNGk3xks8t4Wu/AoLujYY0RhpBez52Hpi2LDGGK8Pnius8+cqL1PkQJi3adNLfmUW/KDLnpM9dhq
2wHvJ3h+8ySallzmOKApsEl8jRq5u7lOfaDISpbX5nU3J/M3Rl0uX9TVz7sSN63lh5Zc6V4rve+c
vKGoz8mi0Qe5yr6Gn93T7WqdT1kZyIfK5i9YL04vDLqMOSFL1hLDtZrA6E7Bah6JnwnBhBFkD3sy
G8ZusEkwNK8g0EUG7JOlX0Pvve7WnNFmN6eVGjPzcxIgBzyo17q4lZyOvqF2nxLg/evZjYUEJE1X
5xeeUnEbXbb2cPmwT4Fg7gL7BoY9LaIW0iuOTp8UQbh39RkRPbJennDRYKr6kZ2qU5PW5nlpWnl2
M4S13aWm6ZWE2Dk4iqoAvvHp/09+Ne1bj2NCdjkCbXfpqWFR0MLobVUsysNe2tkBi0hoeE85WxjL
wjcDbYOZWxeAKHR19HmdJe53LNSVh4Da14yTA+/Zbt5DPdSojDmYHso9koyy7GRHTAQhwCkTKY1W
129ubnwU5DsKrtVq3+ABkj0K2A02rAnA+g7K89Q56xkTaDuhAwu66PBd6EZTSrwKeCI7ctPGprRK
tZlAkuP9Aa0xjzz3VbgUKQFpn9H65eBp0QoNsvI5Exl1W8U8LtbaghMz7DVShyDVg721RRwugrO/
sl2Q44SvSV5ouNLGppgUS4DmLHeFdM9E6xi1rEMEDw4pnYOBztiM8BfIjs2OkhYOH9a/WzN6FqPJ
SL1IqlpOvPYpYVFSnw2slUInXp+cHe+s1NQD0ST1fQDd8SfVZrGcFHGXPmzhz21Riqbp23C+15JP
zmJJiA5tSX8tqIwnEXVe52svZqMTOpQM3Mo+w8yv77SxV12hRPh/Syd6pM64PLSsCf+vFugIh6NY
S3G/hnG+Z4tuJoQjvQMCzm8ArCMB/zmvBZPybybey06l81o1XQXmZAtCkteFXktNrNfxAJzr/gm2
U1ejn1kL5OlUi+ZDat2UlKwmVAgEcGLjPM0x3MwzlEgP1rL64WBsP0rO1pHUSqd4Tk9qrV558Eki
SNe2qDF+Rknr3aVNefGMFRyXkszfFWZeURwfGuPiDuPbD6UCGeLaAO2f94WNESBLDKJ4GPaM5pHU
fcVQtjivdpeKp/LitWRIlZL7bkr8huF5xKK+v8NwipwWpHkanyXDYKPSZVUv8fjB2coIQgTftcLf
xtq8g0K/uaE7JzRI/gVY8tOxW8BRJ/6TsjM83SolIf80j7FMeBbRVIGhjBmm+4GNISynE8ln1OtR
wCf2pR4ExA47AHCayHRBhe2fZHbcUhsUEVe/WPlLro9d0BkCTVxFmgD0Nw72c5L3cWZEysCNF8vu
bnluUA6xpwVyzfUb/a/MsvoimMQtvIawpsckUk6xkjs4jU4dIk5tt8GEa2fmYOYzlmMK5WUfGdfu
Ae8Ru3L3XUGKGg1VrMghZrkAGxEDqNv59/mgNy74P6zQdXEj3GnTbVIyc7TrIgHRXWcqkQsvZfza
Har2gSDwr/AVr9le2kr7ZBGtxZ2pEZW5yVIxgmnlweR1KAOCkpjP/O9J66ZwPwdoRdwqEGHNOe77
JUMR0XBZ33xht9YAbD763d9cxK4S6jpYCsf9NNiUKhKiLxqqR/1gcf5YNzBpCPBmXgq61fHyBJmh
9eZHPLjMWxGB1nRfPr63tOEZVN7/9sJxZmr/iddu4djAB5E8zaGAXAgM2Zx0d5urXmXoM0sN4R2z
ezvfr3EhhLOf6T3nhqru1o01TFDChwaMxNQIsgHAfXd9UfEOQe6b7TyAsKh7tdWefh2U4VAA9M3W
VcVjyofBPSvIqj40PihMPRz/SrT3u8WMYwt5iFUkVFF5q24k4CtJM5XLZcZofSEoEoQlAzZ7oS6Q
oPi4YdthXdTTuwo9JadLgZxaxDdR39KDqhIwf8yMavVk21/Ol6X3ehHuzDYkXSPng/DM+ZisMeSw
gxzFgnUsLGkf/el5QcvKzeGVhFypzsYLbkURmp8jgRgNoGT60R2LNyC2MyoU08+alxLGOi2N22mI
DWMtQl26872MbeBhLG0F0ZsaLUO7MCk556QTvN2rH1yAmtSwheh9gWJbj98LYarsFnxX9s8yenzg
ne8KqiPOQViThZ1HRqmpkd3YfoViTPqwvCBJhuqnMi2EE8b+PY7nd9Akt89GDv0XUfXp2O5JI2KI
9SbhfsJ5+Pmk+bTUiieStlmCQXE00NteygVTo06VPdOWyAX6B7XhaEiMxcxxaR0Xu3LuoNw4jzRb
Xd/4ihLE5JmZZj77DEm/9oW95ycyeHDKTV850bmEF7TCOKQvgZ9eHb9H/hwmV+5lXN2Nlf12rwo/
QDY/q3e98Iv0kqQe8tYWEFenptmC+UJvMyJVfPrCkjesIp4FUcH3BcOpmkshkJQeQu+LYZLFHUjK
w5ODv5ZDXhx8Pqabc0cRz7vAxTME81oX8G6dcbRka65/sxbJvxJCsuzSnaGY3KSYh33HaUKjiMVp
TcKwClNDr+D2wIT4zfaGNPL9doPBdKU8qfiEtmU+OrjOd1EVZijmlIn6LaGzBbeU23OchZFFlE9X
sIjNIzfWG8tsyVsg/7boLTUza2mTnn9GWNVQ7dppfpZ6Koh/xQXr1s2KHazfmiG397e9b0dLGk4Y
XKh7+khse92iKfbQZImxndDj8pB8fS9/1kt83PVZYNnqYkoC9YdE0/l2LXhWdHuax3GVUlPlYxk5
xqpWIgmAd9mhiIge+KCoBz8FuZTTxC1uRt79lt8ux0FJdHm6C7fXPklQ7VJEbgcoMZxxgNSj0JdK
6/IOJX/r5Y+E/8kl1JY1SsZDBCG0ZzLg+qLaRu3n+QIQ4LEPiOAwZ1BsqCB/lV2KxFTyQO2+DtnW
lsuhCwWycwwIsfnRfM+w640O85TsYywWHqTib9tt00nDrER5GKO3ZYJVL5WxDwbFhg934Hyo1UWe
KE2Rs5OSAdUWfCraI+EMRuKF2K7kENtzYCc8zuClKimkM2Aym9rdHnrQfhPhFkxV2Hk3rkANMyGu
qGckmvZKo1jsaa0W/QjwEtvWp4MAVe4vQSugyOZHQ/M7VoCD7UnaiLaNMHMIDKVjhgVuNoxwBt0L
rQWONO2aUDxD6SSlXzmIf/36WhnVV0G/T4cTLQiQ8loKkRbO12NTzMiUBqd7DNdWNg7s0f3IMIOd
ix78H4rPSogG9HlTd5OeWfTkq8DQ63ddmWIztDvwqlr2PlXpJGmE3+Squs0rkl5IQcY2uuV5hGx3
KfT7GbI2gwh8umsmHxh5+WFjGXo1oYJOcrvtLviCh7q0b1J+Z5H/TEO6P8Yd5+XckRBlmwwWPzqd
x8uGRnyzCIT69GsV0U1zEpfayWqWBMsilNPY/i7SHTovuuhu6AwJZ4jmwsVSmcjYzZOZn1rTkrUw
uheEWYYm3GidR8jhVTx2i4+vdo2mQH1SPu35qij88DW9RUujqBK2lio5qgIdoGh32ntMUu4K3mSl
CYDBKPGI8Bjk0B6QzQYM8dDTw3heM9zL3lLZykq2Ofj0WG/mFwUzenaaMfS6PWZVHSjDFzsQngyY
EKOFpyWIbeJHUocYr7kQbDtr0Os0U+xvK6EOeaPX/4jlJRIfcVteSdXbYu23S/kislh+4p/pCShv
7SQgxPM+vPUSQ8WvSyaR4b9ZHS3hbBIzNkq0hOh3+KXaJhoX2+6pRyxQSxqfpGWE4UTxZGCtyJoW
uWTOLeclK8sNxgvwgLzruOBCHuVfkp7PRyLX30/WI9X0mGKnjsddNfshRoUhNB3VWCxigbmRknMW
Crd3Kj6JP4gbIzOKlALryMd6h/vXa6Pd0k1aNePreUOAsFqBDhMOYYk2ynIEx/eKcDBEsU5NBFOM
pw5iFB2mdHC2iREDDU7Reu5AQCXSALHdw6fGkhg/VSUJTcX0UHN3wJsTIRPmDB6hhP2DKxIuVYMA
bYfQZ87Jt1KIoTOwYSPf+/dzBwbpZ7V1HCXvlHYefhma8yS1jZcw/gqtHbmA8tHsxRfgFlai4Mih
2GgnRfL22Q7jETHp+UFIll7sP59ytr3mwGvtl/SN+hDH1raCoipKCQ06TcvUJiN7jj4pZ1ZUREBH
wWl/aL2aRbNPK5zWx/uQetHU/8el68Z7I/iUKki1wFPrxOWLO23Q4fIEisRJJgxPVml7eQNmPsO+
VbBvJ8ilQvhrGHE7ScGr9FKN2F1AkBqXV1LA89gJgn7h4D5oMI6IxWxC0kCymcI5TyJNETqCrWSA
TYQFS6fKtfU1zzMbl8iqMuDuajr1cw2Qz8PcfD3Z4WY8bRgVVOJAc5Hg3KATLKepyC0UfhCw2epe
iR3TjA0p5TEWASNYg8SlW/MjmhtEylPFF349CGj5UhMCZgt1/KS2qIWZjQrhTrVq27m7shEN2wi/
EttkEixZjeybaekZ8ocfkPsxTDPEuCcV2tQoPjsz04XWmmyhHR7uHuomV3DFqXoFOi59j0RGheDn
6V4MgWakMA4TKopQm9U0nz8um3azbFcgwQBi1+cHE9ryjuPxl+vPywRqVwpDvBfK+02TG+Tm41fD
MgH6+ZznCA7ip92/NpquLxjRyl9HsP5Kpj8HIYu/pkcT6vQt4GghzeI0veijk5rSiNBy3LVkJewn
MhhsG7maLJptKiJgPthYxUbloONXy+YKHVUzGQWbf8eovN33ioVveWNjaz1+VzCWEQlwJVhwOiB0
PuXaN9nfdRGgpTAaBZhmM4Rvqg8+TttD96+/2Ht/98yrlO+6u1uKiEGkdxIvqHUMqXIOdSkJbDmX
2vxmmKDgETnixASbMhTR2vGd1CuSKRmJ7pNLrQ1FwsC5dO2FP7mwcrrJbiArPH/X7D9R0Z04SXLs
4fN5wqbXBWyB6yQEA6kOKhbBRwCXz23eLY5xecP6xyd+phj75llJ4oUhrEotDsdpKqODzu7o5HjU
dQQgGzIlPYGcpg0csI8MEG5CEWPmHtmlVMGkVGx9+Ihrev98/PW25GbwBcCsZSRCg7DQhFmkDulK
lltdgwuw1uJWwmbbBK2VIIHMBFIgc3zKL0isLNQ61h4rWZIxokT0v3qVrAoNcKCa22Isod0HXWGL
/od0/4nQCVgWA7GnTBTID6JA9XlXwX279mreFIsASRQL1fcLuNY9aF3sQgn8RgOI/bDXRJWRALFW
rGKr9+F0ymVmPs7vXXGj3+Cr+hdgoM/fNErprqNqTLL1yu/Wg+QzS1szQOdrXaPcg4W1lTnYHJyC
OLoQJ+GoTL6M8KcrxJ3wbwyuafwv+qbnOaBKS+M/ZUeD4rqJW4dRzSFGGeEydVnh1uDzcWXZMNxz
G81lqAKKBQsHsksa6rRiMsC7+RCK1OB00wSoh4yrj+KYmc6ocC8oIhE3ROU1CQkALm0h/bQwm41s
5+Rqiafiwo2VBXNa4gBg0YbUuSygfqp9K4kesDdYMmlDUOby5Q7LaLgTD1OwnOq5bqLHSQkcUQb5
QSCWw4srbeH+JzRTkUHXp3bJjdB/qmiB8/YFc3TdzSn3WD842tN5jQonRTka9cZzqqbdg0gaGiC/
kqGqMdxYRLEQnVxbdosJ6Ty7lKzkpcZ5vn+tKXZgJFPaWDQLQ1tVY4wOeVjtBsPz5ld1DEI3CYxd
mQ9e7tX+U10tEcuX6CisSL7EKNNI8BXYfzwIug2Pg9Ll6DCSY//3LyM5za/RWZQYhXUxk36D9BX5
LBl4eux41zsYJeUg+5RpmpQmanfrgaG5lRKIcmAg+1QGp6D8odskP4Gdodd55G9ycG9CqQcjnXL/
NnqihJx/TCnP+pP2mXyqtjTrg1UPGEkckhvtT9cTuYsJDzhp0W9UbG/seuKwM1W1/GQKqCA/Cxkb
FYX5dGsxNsrPxRQ3NLfMRZGQcQEpm1AN08JuSrHLCFfPNZ+JwWxu/33CHBIf9kCEkS+dvaYTgSRw
5s8dTtDZyN+r3kuRGnTdmp1GcKaEcsziQcY6TYmfecEjYrKFP4PhPwEeU2cX+/sfGYWxwkBTZvVy
+Qat3fsZpRx5jKRXFTCXd1Xh0iiuD06b9WtFoShbkWDgwOZ/duXCfz9jVxGZtLOg+kAEyZp9rlL9
sATcCqN9/lg/VUdx7FHeNKudcmYte5V/Diqzxs3GkACqlssBTJmrwu8fm1OiJoYvGrAFSNCEbdUD
IiqfExaC1OZDyjIQa+4gJ3et5LHJufFCnVhp4KG2Yj69b6bR4XhuUsXQdr3gzaiRFzhC5lt19ZMR
VvGs8KQ5MOMLcGSVmBEqxSthVUzfkPLcaxESmlRd7XzeaTdxsLpsiA/Uq0qDB8j5WO+eu5SMGfBF
QKEdbcnSWSS+pv8ncvr7E+kfHo66EkDu6qLDZTSORXFt+3KSQhWsKrt2jzzetSj6Iv7qHjtANhMr
PGP/qNlpuirbckfSIPWL18y+5dxON7hsxDqSybgU1AXz6iYQSTxkL8NG0YFNOZOtjMhea2JUmB/a
yKSWKFViZAKciimepZZnVM19wxfz7JMphmK9NZTudAskoKTfwUZ1vqLK5gXKn1zwoib/uzrVjIxe
KlJSD8Lcw5s6GPDVZC2OHKOKmlMZJ9WROpk+31IZh49jplCkKntJQE22kV/ASb+yNdpxUk9JMn/E
GxncYHAXLgZaW0YKnulEJrrqzevyBTcfUEgq0jeDe9ndRTpQ9lYIEhda5c05hYJX8Vq8eoUKXgXx
QaKG22DpIRbfk/cUzyxKD3OFVn2Oh0lUkDHV8m6DjoVDEb9Y72D/fStG7tuS8zIhMKop+f5jvVwe
N4BlEkdi2K7l/mnk7Dwlw+HnfpJIgn5zONaDlrzQqvl6opWHDh9W6dqXKP+3Ro2ndQmfK+sryyBO
QEifp77i86mWvg200drn7oJyF6Q6SOFs4ed3EPKHJl3xc83MbQqKtiJa3Hv8zi3UncjankdJjg5e
9LMueEZ3LuY6TpKYZupeYkYDO8oVyNOjQB5oSgoBzaoPoP0VjoGJ39zdiLYHNeusMHZEDOBTamn+
dLDb17GsFkjPawor6xnU5QY4bHekmbyMZBGKIlgWdIMBCXkpvG7SZabiX8mhxKwki4U8TXoTNIhu
EYy/7m739RiiYU+h/4taWiTsQsMtXOodgEaB7g01y6oyvcY+BgB3xgWiYwEqHOeQxYCYsWTAwDMf
Hn/f7beWaicfQSjYPg1XkkdnnI5IwvBFl/paLuHRt0QGLRg/rpN1yjGh+DQN+GF1zYbMF/9hcSwA
sPi/oI6GWmPdVI3rxT2e1ONun0VJDw/1KeyenfJh1XRxFRa/EuE5bn4ncAO7Tve8X1dqn6p+vgjD
KPDGgaSQi8EPBXoaKlUsGMKJAI6ubKGOkM3HWbJz0JhFr1I2w/8jNeuNKHWiX8BplKJOsHyjoyEp
Q3KX4qEMBxbJUDfQ0Ung/6+hPrQLKaPMMWGe/RHAVYqm9gwlkSTLo2AddxfpMxTZrKpk6C7GKgjv
ez3k++Zx4qMyssVWo6Sv/jJZvTTx/X3EHCIDV6/e4pUpfo+tg220h4oxgZYCUUwp+oDkvnIAeSf2
bbfCdOOMHiRd07TmQLOQkCqZjD2xk8EhHTWUQuUlVi6pdHsrZiJ6cCtgqFMyOXu7rqYBF2j07PEe
TZskeFRpNKBYWmQfpWQI/AhdbtvI4fANwWnMj0/+4x6DGEuhmc98ziWH46dADgl35FmF4cFAa7F1
1jWah3RRIQz2fsZ/VF5R3JimaSkftxGokvkdo9TZd27J23kz15JPfVwucajvjjrzjXgpFzwT8aL8
XecvJiCLpjF0Dslrt8s4xUbOh7PId6ob3kxU0rY+eGIoMZ/aC4Gl+0LdM0R4srNKOlG+PNhy1YjX
b6Zhm7KCQWkFj9NFC1OhC2QiHHur0nHOWbJ0Tu6svagCT0aICM1EHYTIZlYyoPAmace5wpHAmCuM
d/HoYxSQGI+L2O683o72y+2Ecs/VpTeqTQsQmFdMVmdMgTt/7hmmaovJdgDqDfMdvLF8pwkd6bsn
Sp5abdpirQO5FpbcITlJHZJyYy/R1HZfMNVNwspsGprK8JVc7WcUoalooPwORJPAfS7zpyv0d34b
nX2nla3Emw+sADE52qQA46fy6Y5/b3etyppWpPEC83s/yWBhBAJQsiZXGrzegXb87aitmWSOZYy/
UbZQUfzIwSr/an/D69EUWazGeN/8ooaFDquCZKkTi7AotCgNhlISwYk/Xor0TZB2/lm8pKd7tqJu
jUy3Vqd0vGMRP2JzNzkk+bqYam4fodQRmASxl8dPekfBYUc5/w76cAPF0IMg02CgDDgjKo/rEvIt
9zPIeI+Z5mD64seUunxn/V2QUAm6tI8KLknSH898mEgce/1xDAHAwsCzl26zJIhugYOPwDf1yQDi
tS8Ph/m5K0AQi0ygYbmZKVZPpTcfOxegmaDnm2rFhgbR9Iwby7i4okRhJBxXU3tFeCuzEC5BCaBK
ClzDZuIHJSXa0rd+ZZcWGffLOcxAQoDK29GVSEeCpVo9kaGiS+SgnF2dKRhXa9P46ADXxKmavnee
esVy+8iThMl5C3mbQRtW6vvpJY6tyMd+82dmHEw9Q1/iJwD8ath5OktY5JXN/rsf6WQkXfcgai41
Txtp28vGWlFCA1Aa5IQqtR5Z9tdnssIw7kbau7aOxQhdpVfdTXikOXuOohSoqVNhCyS/TVdAt2Tg
+p7zfpcQ9vskLzMrc70918TCyyHArnf1hS9yguPnDT8MsW/zPT150Z4MY/AZET00qh5M0dRWqZ88
/4zGZiX1nkfLXDmBRXn54pKJfDuRyw9X51zo8/wwcrFB3UFP1/Tx7CBRknd9x4HyXFDR7WHRsKdH
aEu0ql8rJVosBmrthEdlsN8zzDXu+iDQg4JNiZVYyiT0STXsKbU4cpk79uzjfx+SN7pfMpu/Q1kv
mA6mDMbF1uaXCZ+B6VGFzhhxUiGGxZi44TNly2vfPNhHlA093IghmDeTir/+NTQ46ClJgm5OgDZ+
U6uBERYr/v1Gm2+HMLrMs9oGgWUy9aP9z6z3Kf0WOXWhY5Sqd/IGmVte4HV7Yn2RgCd3ZxEamHOG
tXcWmc4EV+D7lvYAwEiajat1m/GheeC01hpTQqMEAvyys8sbh89MV3GRG0jUu52RRQW4HML2vNFm
LNjL1ZGhyK3oEzXXXGv97QuoYMWy7jXBLYF+QEYBy3ETkACPZ0rnCk6MJqxSWvi0BpXG/M8Hc3qg
mlX2LRVZ50p+DwdNDJAGqMUfdBQrXJSxshIWZwBl+3r3takvx8OkswRgbTM7VQRBfLWuvt/hyKPB
niIQOgTvBd9H8cA65wE4DA6U7w57/zYK7GCcUpms47mwICglKsPsPdqF88Z1MunBb9z8IwE+XC2M
XE98kIKIP61FSPyH20QOw9YFrB6vaL1zOIZWmss83SsHhRTBkmNE2R0J7YigyXOgq0PsiNbbj0Jq
DJDTL9q+O8l49mIQeolLANVNjDhPv5m/RpHSpESE8OozbuNrpnyUlfh0VihFivNqeMu5TnlxgWdU
7Vo7pL5xcrX4FcKvv55nbJqDbjUv8nRsRkYS5wzjr2OlbkRTL20Nl/NkLPDuM0DEG5rRCkqXF6m1
jcE7OVGn/oijIiEaP1HfEGP39isOfLCblBCbtFJom55j/Kmj2LrVKvQZ5b9wkMBi5QNEHx9iZs0B
UDx+zrm9lmSmTJe3gHbDnhxJ7qgaVbzPng7X+RjOt7Y4laLHlJga0tVQXTmqL1xF1eeRKbAIhGjK
YmLtFaZlfYIU8cNBECDIci5kZ6owU2typm2YNm+x2XCWK+rRd+OgksLi60mo0bQ6QbOrWeYK3mt8
5BAs20pSj+K0APo8h3oKXufHPryXaclmqR/cffBcFwTvUG77vPZX9XdanrIHkrh6Yiuybb6seZv2
AOyv1fxrVsVStsfTEMjzUK6R3WqWEl6c0QEDYtnMrOW1D5un8oK5ke3pqurfZtZHFMuG5oB2iOUr
PvbwYsGRL87qyEaETGrlR6+OVq3sshuah47ZzwYn6nCs5wtdc906GyXvFsXnEO2AfrYrBHyuVYYV
NoIlntWKXxvIj5TU7ktOMaGVVp6cyL9cwU2m/LP+ZnKWSWHt6OFLGSCcxGE+AhIuWxsrTm030bfy
cIVvu4WYqPmLjG5azBO4UXoAAIZpI5O82jdWQ7O7ZStD5J0kzyGTFi8DewfgMuKT8Nl0vos9ZmkX
+/TprLwuaXmoatqQMDt+pXXsUqE6cf+dYHC5IC4xRZTzgQeMXeuACYoVTPMmfyswNhbwoYy4N7NC
apiEIggg1K/0+LaojQp9ho3HHuCBTlyGo3n8D77/5uLo65jQvZCjzZnSGUavWu4eHWhFU3z2HkBH
CCA/RWKfKJeQsQcS5GvqcnGJOWyhToLmIjxn8Mq0DjBBubARKR9qlASHlxGh5ShTq3WMo6s6SIDg
rIxhtGHvZshbZ9LXec3KBrHlNDdHd4Y6tsC1ZnwfohXydQuttbWNWYlsQXVwGEhMwN/fnyCBOSlg
mJyt9SnbKu0nVk6DWXG+JnKgWMCU5S8cSEKPqXr0UEAc3UMRbgE9UI2Cd63NZGZAUxLw/uDaC7ol
ah/0NL3W++W5kRsKZQmuZ7IAsIkIIVqkq2LesmvFbV0gQ3j+8Xh8M0OexlFyB77p5sXgYJXJM5Yv
wxODohn8dM5D1cFIFxK7zr2nKC4n7EUf0H97p8A9sOnYB2F5A9RCCl6yyw5nvDLR9Uy5RvOmOPz1
pK/f4D8QQHDbVlJTeX7Qr/L4J+GwTNTVffHguVsebYuGcWa2CXM8lD4qXW3zxnx8W3bnyEaWC0c7
YWDWHfDSakZ2lUfULOR4DTGPJ+lCmwmDbt6dBQa2gKbn1nihz4QcFOzm9vPkce4qvuvcBa2Dd++E
ar9WbSTTcWnsFb+Ygbg/jEMNjQ5N7KqYAhHbSFRcVLu0ScMgUviP4aCZwdT3QgUg7Lx3YGoOPLP5
TGUSzG0gbqDxAa1locDKZ4WBfq8zSoS4rwYdIUC4bGR6+w604md4NbmL6nPopbTZbsdLgbb/lxgG
a/huBSaDNZ00VDst4HHqVMoN6KDQzzLbIo7u/Y9dhpBPcxuDhjh6a59zUSKaGjATwVxik0ZCqTqM
5fLjKHkuzmEh5GYEMbPoOEzTj07/lOSGUWuTYAuyG7lRZwEOaZw9rnTamaUamoIuDS6YVxAL28ng
d884AZ1KOX2VBTLxy6qg7+JpCXkuEIk7hISZXatlZuBb3FvbZIuicS6QvgY+U3c+J5C6Y4j66/sY
D5H3eoOTVDLOp+hB/tHygZNM6mAKzs9KYWlCOBKnvQ0JihJ8uTfMBp6+CyVWLkOqr370wKsh7bse
T3psqnZWF8tfLdUhGhAsOdwKq3m++bSw2wCGaZvKWtrTIdvqKgpDkr1CUNORNcAHgtE3d2TVJ+eQ
sA+MOOh+oN40xrfj7FUkQAtqtAD8K+jvZSiwS77IJqX1aeEA/fl2VwY0OSPbvnZrklZkMtB36C/y
H4zG3G7qP5W+3IINj6o8m7ftD0DWFoYEdccQLMeqpOkZwDDFN1VOfbXegKr7ChxkiunN6T1uW5+c
AWN8KY2SeXv2MFJzL85I7m5b4UxwjqwH0269sbBRIgmSMsCkMgI/wagF4Fc3fn6rVoHOwDW3lMBO
KkFGzh2hihC9ZtUPxOn6z4xM+xjwsbvkQJu+kkfVjYRmT0/couzjXrboGtAb+P83KNxGwzZLOU0/
xfqjXUchoBq7HoLvRM+Rh/6Dm+k07IZiX/ezccda6MwLAVi4m6JwTGrS0ekTBXau3KTxD3tHIlUn
zL8Zcz+RP+ugcn4wXWCe3nZ+Z5jLeJoMVDZPZJVyNFoDwTWffQ5rXXfJeRyeBfixVSGnbSnJqtHC
iS5qq3Dffs26RPxK0Hk9iBcsuA+pXidPRFuLoVPn/DZee20LMJ1qCSL9iRJAvvwaM2+54yHwyCnh
ytp5Ikbz184RRCXZ+7o/wahj6sAlyespwac+qLIwyx3AK0K8BQjpSuhhvV82bqXW31EfOCQWrKQ5
rrAdWLYrGDcTDgHsxmekYHVPlZs664DqXF/RaR4pEIJq8MthLa5x7EufHH2CyneitpnphbuPx3VM
lXMQCiqqAooqXszQwPCaUnyCK17j9I4MVNH/JmHPzsSgRRXwTvi+tw3QwuhWkg0iz3BPL65g+hOE
XwIzxwCIsEpDi+9D2hPGfLAKTMXMtNF9+hpwZgcgYIdAl7hR/qa0olkyAO81RnGxsAcnsgtnHIYi
7+EiEr9mZJxfeoL/yClXvhs+ntQ0ssVRtB0oN4+z6L/H93tSyjOfzRXmV6Z5lV48E7Gp0r1FOOo9
WYgWCTZtyvTXzzFL8lMMAZkU0KRRikDyX+qbKll6mO+3PwPbltfRqgurydwuSmVBbzR1Y2VYkyx2
HwnKxIEKQiFWQEjNaDtMwhnNEE6uZHUogYuibIU3h1WnfX23/iLgDOvD9wjIrZS5aajuqT1awNGV
KKHnbukSU738dtffTwFr5NwezNjOov84x3ambBumBedGo9nBO7mvlVwjAbkT3v1Ytzl7lQM3FCCf
P9Y95kL29nXWpt4Ity3xTQa0DawNLG7yFBEMY3u0WPEu24t3Jz9AxIn0Kiq3m6xBUo/7WrsT1Ll5
Bpuyx6qDkiYYHoi1V0KMEYKi9QJNLWdhLXSKCpFutIzJvRv626rPSOFSjxn7K+olMpmYW5w/Kx8v
X//N57OU4XjHy/dDBd26jFWrsBt1SRcaeW2LaAjYRAiqiwqWlfLlbmr/Jd8GIwyh4VkZF005rjvN
dQ5aLcRCbs2mpvezpLwnVs3KgtPT8q84+zbTyxnRUew1/zfDQ6oRAMSYjF0sRACHbNH/L7ZQD/ji
O+6keAtZaE+gxGHU//fNlgdofuCWGtV66SObM4JvLlY2pJIEaYrTGlnZ8tF8d0nyr1d03SAU2vGc
42uiXNiFlr9q2aYmTT5OmE4S6d5J1/fYvVmC6PI4DTdbDSlg60BgZ+x5Zm+TcmJ9h/sXWVyT+CXX
UPBo+3mWckPgskYEhmkklJaoEs3aoytlzZ1Hzxc3fYM7iKcGFOSPC8m2wdWvymjWloT7OOfowZDJ
eLctEFiPlTMjEIWF/cYb0ng/35hY2tjDbepchFftuRzZqxYp3zv9AvF0GdJ9WjLOW4KAFPOjPVeo
TzYSJB8ClrPMAmBZqqRRYDS/aKLKIMaxW5Q16bpxrrTGUPmsra5k3EQWa+9VCuHav7gyGCZqdWzJ
Q8Hk3glwwR0EQfQjxP7bdHR+V8TjqCjn1K1RInsUr6lEAxhmhXdpWs3i566rPH/95HbgugQiy213
PZ5r9zvI8XHbDPZPNbNyrTa0QiY5GhgmRcjH91fobBXXo5L3p6qmw0KPhSz5A/06YFsOI+y6gKLJ
ML3O1WcimycmwMtNO6BXY9UAnxvxRFIrELyjQmiHnp323SUnQNwHdLZhe59mmbWWk7a/RS037PKR
jI0LMG2irxUaecoeVafS/Sn2a5es8XIrblt4ooIBdxecK/igDrzO22LVmqmLjnNCiw5JX3zEjYZO
XisLJ1K+B7vSVVa50klUL7PR63RnuqC8FXiwZlXveSzurIJHWYlvSoYLPo1z9MbD+sOSIczy4i0w
tZB8BJiQQSJ8VaHWeKZiM5CddT7ZClpbnkMoxngitaQYNSmGs4pJy4ItmRfu6bAYanBEHn4UDboI
0Mx0eM3LEr+gq6205zOSMXJQEU02UsKGf2pADKNEXNl1g++B6AixhK7Jlqguuqh75D4CZQcFVoTW
qlOrSfKwh7eFbsu5mCT2BqbbNLxUUuHIVQuIPVrBRhoRQSBLhJmQQf7WBzt+Gv4TUPVe2B+dpXP4
eFYWqobjESb4ugMd7jNeElrNazWnlTSDJhSUtcDPAzs7WgEAt/G6KWlqYu7/AhPqN+kzRBp6s2pz
2MFiT9V+ocnqOPkWI0gcpCUHRbVYyEFPpBnpxqivt8raK+A8u/A+nVI5ZWfiTiD66OIVx1qk42u+
43yp+DhI724g5bY7Hp4FHQuk4tLAW5t5JoIV699kw8CtqOas8zwwHFrcdZnEzP7GQl4/0PF/HVVJ
IrRF+nEvSXfuuxuKa5gPcw5Fn4O8LlNgJGA8XnvUd9ce36AWP7f62buCqAgCx80QEPjShl01s4uR
TMaR3kEo4atUQM6WXNyin5k6M6EZEA0ViUBKlLi2AdXQRwWAlglPo5mPf0LoL65k1jTkAfa99hWg
2sGrVp/Xa3+z2cBoWndlEBlaFZUL+oNqKovvFJvQat9R/NUjAxVPKB96vj324SwsN1+6YclBOFs5
l1f10FpvTqGNZI0V2c+RwtxReugBgolHgHVSoaCOW+YBmwndFCWXpwEvNlPQvHICYRufQQPcNxQ2
pYMKhzqO4BrqTJCnmIfM33UVoao4NM2na4a8QGUXAvKIawFEa6semG0ogqo4gpEeeczLLLjfbMa5
qAg5Mf7vzz3hZKMWbkdobrT9UesP5E2x8ncMYOQX7rtahfg/y1Nq/tZTY9JswdbkZP3+u0xQZxGY
ACLViFjDaQ6tWKNkBV99iYJtkJTCE213UT34Nd+RJPKu/FtrcFz11o7SIH5oL9DSXjOxr9cfPKwY
/8181PMcPcl9Q+Aw04Sy+NHvkDc58QtPqbnMUa/eEqXs+gQj58OZrLPKsclzBXQBNLnpbe1sldR7
+ge8v+huCEPIzv9V9sSySt2mGU0eth7krIcqBsIduFKP8I/yj+OJ/3x1gvSsPJ2rTnblOE0XF/C6
WV3dJXV+UM2B1NtR9CO9jPJSYBp4LpjTcrwynNZbn3NlItePYQacR6U2H5fnLL4lyQI3OzImwC5L
ZHCk2Ca7u+IXMU8vrxkn6MTrzQ7uaKGfndfYF+1kusswF8DMi4prpuyFuYROJjgrGlxOeKVYrXUT
hVcK8agVNpiP4RVHqy+xcpOuIvy9yZcRwc8wQzxOqxatUOyle77FeHYk6RRhShdyzF96+eu4hB4G
vjeK5FIErdJxYbspDktLF4hSW+PPDgOdq2KhgJ9lvhtxXPK8IS06QRTpRN85XdPm/1goeL+7h40H
vC7ZxYcdx86PMqPsTVgJALoV5+GDaoqvaknfHtG6vJkBSLzunQ1sy42eNyqiNzFsLcDSuI/jbXe2
E4e6oeNa8aXAGa2HBzFET/I2UIVqywoY5IYaOuexzdI6wgn1F0b7TEwmnvCycuNrL4kUTbIZsvHk
ueV3x4x/sKnzvX7NaEHdUJM1N7MBeLYwUl8trFieRu+vKswDvT4JZgfMFKO8CftgYVvoYYUCllsg
PZPaZrYLB9+WdSY3Pm8wgX1OG1Mcu/58FTvV67AX8Mse/B55VtOXDBuUXl2k9j6+o3SWm1kLVtGr
2UTw0N+mYbYWHxCqBNBzSh9pXuVof88niaKP3lRNyiqkQh2J0ChDkhUCEgGXLvJn6TzzpJdqQTi3
OWjcv900UaQ6SewUaNh2S/PoP2lyzrhVPam51tXqbOe5WrFjxH6Gx32vvZf5JCCaSv5kMcEi9RAJ
C2vRaRrBGq/UV7deAZp6uZEPGkK5Tl93p3Qb23twXf6XmzRbNc3wzx69Bi8ZdjDrSIRhuVNHqCg1
UPuHDrOXqa8hqvci43jv/SKM0veGjLcGsTXaQlEiaAbUheRBDzfcQMxB4al1jMJphAycZ+/bfCqA
WaBMQ17rKuJ3aBh5xzZ/+LvXxsw97LzlGPSsIlHg6Z7fZahcncu8Rbsq4HWv0gnSTmS/d3Xw9waJ
0YXcMQKEJK1K0H5haCJE0gCttRrU8VHEqotn03ia6ud9v1lRIAVn6O6PxepgU2tTL0N9jQ4G0aI6
y3e+P1hbjaao5xaBw1f1GFn8xQDIRh8WjLnefMfD42j9FL4MjI6d9sndjtxlQQV6kApHPiEAU7NN
2R7TLcyRAHOvJGoA8dZ59omh5sGv7hgqa6AFvHuHCk8hprpBKvTjEriwykYo/ZW6yVSAByo0M+jZ
yKsdc5jEGAr+4vmJBnNnjY8bpTyoZBa3P1bChxrwgvgshLIIUJSe8/0Q51qTgBDKB4j+fptG+vyI
M8wqoS2xk4mJ/ZrgGpK1vp6VVmGyYEmmD7O+g6fDh5RRgqRjtSS4UFooPLscr6VRhKkLMemSJ54N
nnG9klNJGQ+ytr4R4HVeo/dctA4OsYI+7GVZ5VQXW2JWcDVMEx/S+nAnBnmjW6Zx9gUR6yjTBnGv
6aNSgl+u+4D6HEmkYbLr8UsOvqq2ub5rcBFS0esrazAUZRarxnyjMo5WvVEOfKo67oC6h6MSjCEF
SSgoSbs8KiC8xzrdL4p7YfIJhlO9sKRFLLnVxH0gGERB8I/uxJrg4qG9/bGz5G2wM5PFnbSIeOA0
AyoEtl/0nBaxHmjHNYCGGYh8yMkSXSg0D8lKX4dVf8du/pLg+d7QLAwjYLZdFTp6LFCvApIzdxaA
7pos9P0Hio8vdpFdhcn2vMLy+ALrCR99CiEl0c5MiyRWlpOiGxlGc8SiUkNiRyjxxsb+Bg1cazbi
jbHIMPKpD7dTRj2yK4ee+O2dHZ79H4uiHzNYbq0Iz6popijYU1W6kEycOCJ4Kz3n0mvHLD7PY3kS
Oi3QfBM8yjbMaq9QIeQqqSARBt4DX1i3tWmboB72ObXPPR/BxxSktH0Y+53S8ajZjyowFVMEOYqp
2ObKRSUZMpsFscnbbkJ7Y+VLcaPMMOa3wKtzQjc4QVvKpalT9nnkW/pTlBVc2SQMlZ4FiiUetIsg
X/Kb/AzonISKkUutF6HJzD3FK9ph2pNT0umJ37N3f+gJqPNss5b80K1TNlftHyGFWfCxwZ3nuxin
1hMcQIU1poyROjUz1obn1tJBjpmXkvEMEAYsjVf/7tCQvoXhf4NPzIEprNE6xcEgCHN7w7P6qOO2
OLtsw52TT59XSS+aJWdAue00oYlm6wsrURBBmWeSSbc7Dw8bajo2tfaGTsT23y3/ZR2ZxcZd/yOL
45LtBA33PG22HD5AnYlfUaukTi5KbHv0D6T53teISvbd8ZQl+lgkYyb+YK+ZClOPsoVSTmbdHxaW
9yR5gFLrepZpsmOVySo42y3i8Z6ThtvlDWAdVyLvqmYQWcSchX6Na49D7M5Hb70PlIKtBOl+BEqD
kT/KZ/xlrFlW0VeHJL0HuPWUeTaUM3tjmSzrMz5RvACEZ5TEckDN5iA3FKf0N40Oj7yLd6hSVGOU
lihEd8sDTbgT6qoB6+zGnxqBc/SzSEvWi5HV9M1kOPHU1iKahcXhA80PdATU77vqy2FcZBpXJuUF
Hw/aBgNXLGFPWdqtJWgtXNeVBd4Adt+YY1kxgtpHMHu0oMnO51tkbacUnQ7n+hg2/x2ZqJ9Q7s+/
xCLezew4Zn4ZmUCj9Ho1ztarrsMOUWLYjnna+XSlW5IJx5gfv+i4d/S6ab5NZF0vzbSPkagkYc9a
R82ORvOpzHmEn/aFTV3TMT5DrYrSglnGsL6Mojk9yKMgYxtpfc/PfSmY+3BEY6O/2I3F0L36tk3I
Ns8ThTn/VCDqZJLbN8nW56i7l/VpuIVhdBgZV9K3o0vN4GGIBdYes6fu7RjojKUi3yHWhOIKkw3c
Hfbb6o1iMHOtqvuNgqPpEH+Hu4lUU0ng8jJd2BUDoW+rpxvuxjIHqsgQdJdkXTNtYx7/zZjl1tdI
c6QUm/w6OpDyjQpqskOoZsBg1t36BJQxABdVp1I3xUSIEFqBsaeFUoVf+ExxcQO3u6HvNjdR0587
sf0G5uc9/g5UIu3HS7YcT2jODDvNwjxwt5a/P9oosubeDnKPrsLG4qANWf2c+cj2xW9qQQP95j+E
H1jQLVnlu10GoqK/RrIEgGfuowwS4UxTE+LU2CcozMieLKZ4k5zoHX6r5cHXnWX+0zkh8L+4XcLx
sXypKdyel5GiFMfnTPCIN12VOb62Vc4ahHTWURnQmiLkVC5v5s8CBH3febvczxOP9zUwzA7tQNrs
fNk++PwGvDVsaNk9ldDXd/puV+7ycQlMa0fPBYf8TeshLA2X2rD77k484v3oy7fcrmSfi8T++7rP
c6ihyFC6vC6oaFVKbUkUwUOPjL+8jIPp+DXQ3plKu9s6+Kk/qI30xVe8zRmNamIEfKXCiR8Vm0vO
bnK5D72k7wzA9VVP6W2Kr+RFe3TpRsmg6LPqpKhO7fLl/52eviivpJd5yKQMYlmF09P5mRkd4a2Q
ygmnCY3Pq/APWjdW6oLLNejeRPVNKOL66TazmfH7SrIQeHkveJftOVXFrNA5VQXxaq+VNcXlnCWi
gRxjj23+3pHF7pmgjTz66E1UaQEDzoyjvAXeJ4MmC2pxmlLuvJ+eMyNEOhQVWthdd/V6GU/bbZY9
pWQJ+KC3CV6B1de6Uh/eGD2TsPBCUh1fTqDSfymbZcU31QXR8HCCbtFh5IF0jGYuTpdZiyrXX+9E
rgOIz2ynCpaYuP1xGolU9HzJpYRgD28mApv2wJYhEp2AuzjjNFLp8MVcGGT1Lqg/n/1b43RORJ21
eeKNR4YbkRccEQm+8NANFaTtKz3pQ4U/+v2oTSl8k0z0RwRsYl4tKkdmFfk1bZmh2B7rdo7orWMq
aEkYmvMr9KTLkXY6KH6/1hcKb2Y/y8vwreYpJjm76qPXT0TCfLsHPERopPRKaB12ZEEBnADhSmrt
hqLbHjjYASteC4Wa7kosP+3/La98fvarMg5812RIEhf1+J9pjfj0tA5fCQWyFLe3rVqbd2WuFV4B
SXDz+UkIjT/OQWXeH6V2i6tESUwJYZCxV+/k+0flmAbr4nn+ilI7W8cfi7h4oZSnbBHaxPVVOvgg
9pYFQb1OsjTiWs5mPKzFo1FK5cQhLpgeP4Im9Q8XnH2Pf3cNqb9xMDZCO2e28qh//df++MGZgs3T
GVoU4ll/+2qjkVrABMSKei3satcHMJvawA62wWHvmnsuezlJ/pWyi7qCi4YRgEvz40eoDy9ZEVqy
pdkIYuCk7zM5f3NPMhAvBCZsVejI7O2flW8ER4GbsydIZ3KFx5gbrjjBMHWtpkbIgFOvpz2NLS1B
oluyN5i+pVFafcBxogrqnaTAWJ2jzcTsE9NX6rhD/fQ9L7m9lmqfUYzwiSAJ4mTZwiyaUjAR8kfQ
JsPE6KDVWijAvcOQR9XE+/dQcffhFQIzdtbwee5WCoOc5KPhtLtizcc5teB2NO4MejShcfxbt31A
w6N4SyfBprBQi2P13gSHuzjVbC2NSJh3S9nOVRnygja9uLhZcrs3fQ1V2Mpp8deCyxhyCNLfv3Wx
+QeYJJSoazLw7qQu0LjJbxWJsINwh+KdiV4ZwvjialjnpWBh8CXrkNTF2dfLxyR4/eLFUkSlNts2
wB4SPSrqNaC7xN0GzOe/wWh7LgGGYsWV/yiyKXQncnnm4jtjn2AUVt/Ty2uN0CP+r2J613pU/gZj
eT9zgnoHufbRrMZ737MDsBBQ8OBPXjNrLCBj7Ie9XdWRpyk2VHLVXiPD5aP2QEZTYODjwFanuBUl
RpevfjLWWneV8a0c/+BElc2EkDgRW0tjyOxxEB1FWvRiOC2QWXRIR3u+7EgXCmiVs3xcRBXa9gQH
C1m53NYd5J4IPlzEhhs62Z1mLbpem6vNl/+fIfD0vsiVPrmMKwtIZhZi7PFEM1Em8jUD+yGOsXRL
Nk77eFxUnEdjrAL+o8aVlj2pH/AhSvZdfKrMIV4ThWp1RoGsUMxvKTmZxAb9rN3uDglUJU50s8pS
6Blhdon9bukdCWdD5yFJHywux12CDclulY1t8VC7LN259TIPgbWbgRKnAQ1lilII/tg1NQOeKLqA
HFi9eOp356gZ6WyNhZU0n75dJz4/qTSvfNgtx+y5SWxRX2adEPn/GZlZq3ooXCgfi6YVo8ZkuNTw
ACHD7sNRSDJvizV90qZqLu/+6n+5pS2r6L91REGFNjagPnV7Kpb5lxUHDtrgrOF9XHNCOQcKlh4z
I5sInyuX2JBrJhHnbYZUD7lPr29K5MDQceji33cPSsH2zAuzTnSDuHulu0OgTiDSCoAetnNYdaBI
MvR5Z/zn8p8JpYDChT8iC1uZu+yJdRMqmC/lT5lr7+HHZraFzA9Qcu//Ry9X+DnsbTJnfCe3GnHj
2vLUmBb83+DzmyWji2zm2hAlYoSYQ07OQ0K7iCpMjkhP961sbg/6EcZq0/GtWyyd+xfL3q9ZRJuW
pKyhO2dPatL027TL7YUa0/n9N5EuIRULInZJpVi18FMMwfSOnfKTfKpHUjTv/biC17bZD1adUGD7
xNVdOKJ9wbNni2ZZorkpqkQxLWZ+6iLNsELN/b1O8v/FhqrKhKX/v52uqX4+qati2SW/OarxNMAP
n5SNfIP8cmC1nafiVR8epsJZOtrq/GoF4PY5sg6MOotTcbYTvh69QrNm6/DX9iRFMOBLY8JEzit5
VbTquFBLNjytH2QcrmvVv5O4bXXD9TW0Im9qKZ3VEPMUBuPJaOytg7Jk5xkJLPraagrpSoyOQCwM
ayLkwayMZ4A1uTOid20oObglx73FRVm8j6UZaBALzSXsAlonndMst6JIRK6TynEMgFbYw0nMgPQA
IzemjMhDmTQ3X6LtGJag1/dorioezNj7HEC125H2Ztx/6ytpGHqMnS6xnEMiTQHXLfgvJs5LPQwq
GyEWnA4taxGZWaUjdLFHKpydE531fcpHj3J0+4qDTQbZJfizFtid2Bc/EFXBLzaw06DlFwWCVPnA
qu8LzjYqSdIA7rK0UbDR+Fg0qkkN+oaaiWoqM78gszD0yt4x3gDjjV9U2WMo2A/snCJvOCEn34Qx
iFlxuS7YPFXUWBo2Mg4N6Iup0tRAnBo9ePutKB2WmWAud5U58Lx4tdZlC2B3GO2EqupSFHeyzHhk
0SVpKqXv0yfcCXtQFstHFiBKQDcYpGOHk9wFpsC59uMmszM8EtIKRo3jJ0gaG3MapslZMQjfXDIZ
6eVQbHhozABNsCnicGnZzKnG/A2THRw6YWAPQ1DvZDfvaLZZDL9lEW3IWinwGpWNyjMhQZmWZPuy
DWS/VZPrLAeABnePEDctnMggqk3GiLXsdxOZ8GL0p/GNLEmuFgUVABY5ZZwEMm1w0wI9BPq0besf
9j4z0KsPjxugCSngff2RQyEZEl+6ebYdvfkmMDHCRbM4l9sRtVE1F+Sbox5x7AbrVyNdCnOEoe8H
gA/AAhum/C7tGCoJLsnd3eoMYMS2PdRAsE0vbnjA22iD6KHDmuyIilwCvkoHK98+a3iRObw9Uee7
XLPgMXE0S1/2amHOX0tRFR74EZSSPtCZkGRUO0iEoKtn10jlXCiyuEXWSLTsDt+SxHL9dEXpoMGc
KDOLyRIDMzmto7CnSbAY0NLbnN7LkJwGMwF40d4SVVHrEG6QksN8LkweGDmN7sbuwp+rdlrQpsAe
cOzbvPeNmMGeaECab48op66J3nRdrZsjDtz06VTYMNXxTW7jo0OkbcYQE/P+ki49eap2Rt43bUyu
gq0FcohEKy//D7SYDNPEqKUWjoZmnsJdhkm9i7ZRJTIc90Q4O2nFT9wzkuqcF2cuNMiNnu9bSmqd
tXQeSSpYjrsGmRaMe+0RLyQfR0rqbC+AOU5D3N2YxG+U1ewQzJpjIL3SC2IYGXXqci0Gesy/6D/n
yphgG5AjizFiZ3ElOg+NTmvBQHOWCO2D+1RJTT4Wxf5ZNNcTDkpkbp/o6F/4meDxUFZPt1TzM8++
bt/ACjkc15E+yk5KxGsIcCWfdiMwYphU9yx/VJ2REuWNw3VwNl7xSKxHw7lLv7L1iVdIrhvRG7Vd
mfHByhZHa8X4JvOjAv4NJ1okeeuahJZ0WJynOKVFcJ2jNZ8MXsjSXvCFgd1k3CIYeOkxQ6bbZR2T
Iyn//TqyonXkJrE0qQPw4jDgAS7wd27kq9IhsS+OicQBD2VeLpeVnVzNjLHDtigmYaXoRyHSONi6
Loz7we37ZV/h/V4X/YjTvH6arDofvIwE2R/xwYgby9OX7S7hBeZ7tExCT9v/v/b4DLXAfmuxCyvq
w80NhINrfm4Z4jMlJGWJI/nXcT2F2bz9SHDwjQTWTrVso1TuktG4gim2qL2h102IGb8MpUThMvyh
Ngb6TpDyNqDkCtcAlzYhE1Ano6Wq9OFBtIRIF9yAU4jWrIQjG1iAgS91GUWdSru09+OAAVU9tKU9
+TEHthq56XMK/V82XEQukBD5KQ6Swgtbss29KmjOvodlW+fL1Rn/Wvf95XtrxwLU4/PMj7Jhbcpg
isvS9yheYLfAT9StmCV30govpb2oNVUOW0VNa643X9NrfsnHJiZy735yt+OnM/zTfuuPLrroi9uK
poNH7zC84FqewvEx9xeWYFIetD/83x/Oz7Ac5PFE/Af+gCZH7iQs0sM1oRes417s+keBQTAZ5B1w
rbEIWzFw3stme14rwZHY+MKH8BAIePN+0PPzZuNoozlYtCAxgBE3PYYo+aUkT3dOIjlqK94DwdUC
1D/hEzzICduaslxjlMres4hJS5DO6AVYoNVfxknq+DNCnKB3lS0Ds+oNIKA1lHHlGeY2LQh/3AQX
7CFmtTnEy+vLtBxs1E6z2exKjNFu9S/yBPZSvBZXX3XZajiOI0/neJhQxPdqU7WvC6xwb42drfI3
u/XzFDBqFxgKZb+cNXD+HGBKjzra62VobL62XkVEZt4nAGLWuVT7zcEl57R/jB8VTmkU5yWyuGWI
8aHzfXF6auroL2snKdVBCqssUb1iuDDFfJ74IVJbFGD8C/Mnfn0nUvuclxE1rkoPbIe0iF+5jR4A
80mX7Vsh9x7QG79PoWF+0vYhwJXHqYdzvBMHWgaUoURJDX1mpOvy2ivXWjaVcF5VvxJ6QNJTFxmB
VtZukVqVTCgROt6okFYh3QjPQHBOzww9/fWjQw3Yy2pcwrFSGtH0UIUjNXdzPucfN+30qJWc5xNF
ZLWecaFFrkAkJ6WEJwY6YhXOcrVCGJ8IDDd/Yd8n9k00YMOpZUlOvV32gn0l1zdG+BUvnPWt9rb5
qZcZofpOeroJN85xwN2RzT4CgsMn8spkyqnLiPiOIqMzSnDTViT6/S3c/auLiR6v315pN13Nc3L9
z8XPyL79m790HMbrZaNhG19LrlSt3zViUARkw3SXP5fuKs6ok2j4t2Y89A4AtZersp1bVhL5skHj
7/RXZVnffuAerwnyOnIgMP71neIyBuQUK7dlra82FVhLsdNeUqOyCZ94ChtKh7OqAq/y11U/dGJs
XamBSbbyDpf297k0mWj0IUeatq7rXYwhcRG7JSvdNB516SQUw7U6CCw8DnBkh1hUEClDUqgaTHYL
W9jh8Gzg5PO2MV7ko2R9XylW4QGvJcusUdBwrVqTQZEmRkQ+R7WUshw1hxuPKVVVpuI5GT0tIe82
d3k2Gvnt6G6NBPTnYKBgfuScuJWCZ+XdWaTrOMjJFpTc7xmxZr6eqPCnFyXw1doi8xVs0TbS1+iA
OjzZA2Ar9XKuRtUKmZDGW2PZJGoKGNPWNs9/Gzx32bv0VGMMy2UQ2z6GTuCK6JIuvSt8f+yPkuqL
cjZc7qOKgVvsiQAkYImUVjhANTaVYiwZ2AvgTBdH7YLGcHeCJoe57K2mplexupoe8o2uu49nXEhz
H6ygqD1DXGThXl/OReWIjX3hb54o8zaVgxAedUUSazY6TjbfjyFcotTnQBUq6KGpLe2MEgpDFkSg
P4nASBcmfHNC1ljzktIYgm+pk/rqzRoA2PdC/jeMqLFSwMdTYGBfr2cZeGTK9g/zCgXkgeK+ho7w
RpdRxGiM44MgyO7yK4xamP9ejha/PEQknW5QQPdVygcsy8LVXkFc2Cz5lmzL0kOKUUPIvEuK2pE2
8RyE0dFGEziMqoZqxFpHMzkrsVcM/BXogOCZS+El9PHf9M+DC+/F+aHBPaHGlW2J4q+bpleeYKX2
tZVInSDPju6HdqmW8iFbrw5h63rPqUz3zKt3Lf2hmhzUwYuBQJeul3iIwnGlQxo3yDMWhaPIMekN
aN45Zefp5wz2iYvy47u/yvr2kuPUCIUfUpnuldorp2aI3jIm1wcCVutlFZ8ZA7KP8ayGagefU7+n
MjJGE2LFdHwKl2wimh3wkPl72V68D/iH7rmKMRxBz7U4b2i6vRbw4NFvTzSxh0MWPZv2XacpcarF
U50YPKOFnj5dwrKoP/SWV80zQwaGvsGAs5+XOyHKIhm+QSULz6g0g6Ncy1fQdudq/MuWLXrxp62G
ZQHweDpDLTkaSZg+fZ4uQTCdJ+0OM+y+afZTA1OwWN/IhL1GmZMmN+uaT8WuA7JdZ4SWoIutcihx
mhbr0aTZRmjobL/fuIxT52ID7SoV9XSvt5LUHhiDMRJybdu0roRS/u9GSb+J1Lxe06f264IJJ0C3
QcwRKAS0sy7qWquY48Gz2j4vnUJ/0cz5Pnzo/8akc9HVhNAzt4EuST2AKGqbCbpKnWI+w06dg280
Y0mV1hTsWeLR7ws6bWcbSN+qRzLpKh+vlfhmduRmn43+vVt91HtiUsFKBhMTTuI6v5OGCZ7nIOcs
byCSSEAxJqBn007LIyDf09GlES6w5FF+TO6q/Re7XngOqLF12kVfH0dRxO5dplw1vLmNdH7BQzOw
juzlPjc5kskW4Lnjb3NE7uPk+eZtGs3sdgzZzxEN4Y1KZTpV7TWIIZkCTUX79wPwSui6SSssT39Z
FXgHd4VhmjY4hb1TyJBsboLiPyLc7iX203eErEYV96V8bxKo1QN5dcVquqD8pHytsB2+2dTcABMS
gMEWqebd6pv1KZ+Xhn/Z3APPIcrPlIGeGaz42aE+2Abc7kRM9AeIUOtwDJ75EstklOGwx+ocGSgx
kcMhklxdLKpgR0RAtOYG0V4NWSbzICrbkxELcK6KC+cWICj1f67tLMPl2COhMT1nKMt5PJOvwkK7
FM7hMtCPvc5XYDva17EWFijC4s9jbFDyGpN48J/GnC64rEpTjjoch5dti2r7s96z1lY2kKJFdoOY
J4mXVutjNEVgems5f8b/9lqx9+j0o6SvzMJQFL0JHRYoLoQcZIJAmwvLA2E4YNjjcTot/qWkyoEQ
46nYdS5J9bj+RLZbidnRsC9ox8iKeoKDdudRjCmuM81M7Btef3Enr8LL5zF/H/ceyf5dI/vrg84u
DTcDWQ9FO12dcsVP7j8M6lnylDmwQnpNSda/05L/SUV05vmBH5tCje9ZBMMbbK9i/CGbfTv1MkgJ
KJO1MBr+MJaH+1VdM9o1dTRf9XJbk20qQ780vxePQguvi95lBtlhH0IILPz+nFa/eXWR5Uer2xhl
xg89kvkpZMOhdxg8tpL8LNvFua8RCyzoTRiK+WPoemukX7flS+KUQ/9/fgpFm0qoV1OCn/y+pQBn
gan374W/tj3mXsi9+OoqPTsvwADqt3JBu5L1W3bK4ZAwIyP70WAIiyBa1y8jw/1u6kq0TbtfC9fc
B+sWGjI0oeJq8+4CNo1KM2CBZqfmiwlneksEMPlFPhgl7CG+59pnwEJN7TAUTVDODoZZbxY9/EQw
rKewuk5XmXj/JIY2PdKqqEBWshUNSVZmHacGavqrHckyrm/wgbi3H2DtFdh7aQTAKSnzjGLZBwcl
KNAKLVlCSSlOnSWLBY1FJfJtLjIdPWjCqh8Yj7lGdwU1rSP8NHUwJjhLHN3xj10jzLwrpvJ4rjXa
W6achNX6uXe0md57LVEksUpRd9VzVnLDHLhCQZMjNf7iPoiJoUU46KBEOI0/JMV5ru1XfzC5FWQi
kXJPuhKqPa4KyNtVFMh7gqZdl0JKGxpyTAWjNnVf8/Ve0I7qew/h6LqDP6xKfCSz2rwcPOoqO2gt
uIYT2ftnjJ63qQFOVenl4+13ar3Uc007QuPv1QEwFzjIezE+yYkSFg27VyBcpO0IkJ6g0e/+3hb0
XcwZMrOiNJG97NMjE0eKmjfW483Jxu8nmdnao6iVdtMv6XSDDbDu46VlF9e/Yv/UaZmA1PAtKTWf
dTI88auiH+lwvMezKT6QFTGKgiCy9yyLnJL24CfIV3hvP4IyEZNhkiWD9QEtJV9ENGrBZzi3hswP
0c0QgPxjEPe3rmrdkrR3lmVxtpsZSW7f10JtRAIAeoncpJ4Uzn4qiOd+ZJeX5w3mHC/QzGnx8qNK
PTyv9CgwT64/1NFNPaWmQBizLhyoarmYjuriRT6cIPGWMdv22SNUv8KYMNWPZmJo8SoIaB6K1roE
OrzYVVs/vXq7jZ0fZodRoAvAVz2Db0mfrYTkSxxz/X1WKtjEgQL+3vJuqNFvt1fGve4i1x+48ODO
fmC85WDdvCxnWZ+biAtdMY1o/haO5pIbindUeS6xEW7TTyKzyebjP2qi/N39RADJA3FeT2784lvo
jTzG87p+Tph5HtC/Edp9bjMedZq2KEOvde5nCminW8U11gwvrUu0vEBRkgWsMuq6DsP9rjef37E+
9CLUBGkhWqCqDBtc/mK+V0ephvWuOUtYxvH/xvLR3TPapfbnEGKVoH9ztu/ptN/I2E/VYHWR/hy1
4H1gOOrPLnTK/EYBPqha08wVEgSqnQPhptVDdDlW8TarWyK0A9UttO3rnEQ28zglm7CmR44A/5W8
FmHxr9HDGBttWrL+vt/3DjxTBQlm0q2FBExIfEs7KfHj/6ILx5lPwScToPd8eOC9yKbVZkwpAsY0
5RW2eJsqaPQe3+rKp2zeKkFa+MkByCmJT0z/T01Tp9ug3QbPCM2kZMNfXz2A6zZNn2lqKPHzklVx
NvChIpkAOLgiKxiVd64Ud2qe+Qr8aa/oQ/VFqEp5+ZaDqxr5VYCgh7iL8H/oBqbs1cGNg66yUDSM
EFGC7DZCIR11mrxeE1hl2kDJ9W3O1MktEEUkdCnIjjEYsV3BpgjOV8WJo6AHF1GEIke47EeBwt/M
eLHynXJO0UQEn6/W5lHbEsQuIbl797uNDuRKiVfIIsnBEzDgOFNGz1IIr5PVv5KT4XcIGJ2UVQ6m
UnOT7TqifO3B2PkVVZ5VxBv75x1UKIvWVwyCeneZ91iy5fzX4j3+33vxkqCbGS9Ppu/imjXv3m+1
GtgH0JG0p9XR2SXTSEKUg34S4Uv22yg5THcOYNFPG0Y8njrFEdMf2JW8YdPuiUhho0K2/W4Hz7Tr
kxxXXXC3i3d4rDkwUv4ZO3qykD3+soBKOOOi8uQJRsLM9x4yXy8o+gLOma4GJRnvpWwEKDaroLJ1
CGJ9fOrdxOmvaPtpDmuZMQx7yegergr8hKfvnivdXIEWLsgonwQ8YV4WMbf/X6lrui2ip/zJuczD
IpEH8PTudXgawFCtRTfpRp2UrvBjqcRP0FjhzbJZ9fR+uZ/XkgCN37aMMrUwMHSnDaZivjaes1Xw
qZgoZgQ0wjY1qdv8YrsyprFs0l+JC1wRMEyn3PpeTWrMj/mKrIL5jACehImV/XMvyw8CDbWMXXzZ
3GhyeNlPAwdbYjtzO9WnvlTMpZ+mqTw1zzSZyLFbb7TeWJGOSSX3pW9N1wqX6m3RUnDnWCj2MAL4
IL3qbOkbYeeq31qAVhtzGLMKU0O+8BKEcGYU8pwiWAY3c4C0+W2R/xDKSDvkpC+ZinZ48o9a+Kz3
hfjV1HDfmslk5N/TBLBfILIWfNHWbekcnGmPkLvEr1eARZwKxBAXIZqjUTugSCCYlOfQCVWV7aBP
85puvtBv+YHQPBn+ElbjV4GfMlQ/Gz10qk8EPIma7O5U7cvldvaj7+8+L5/OOefICYtLR+ual5bR
87DOL5fhYIXQejBQomcExg2aZnf+I52OTBuvYLULD1ToQXF6i7fNS0Xw7Mc1ctmuZaSBSDGUJXBw
dL9VlZO3/L7EykCeDlWuWvv8ls7zcMzfXG5ZM0zvYy0KGIDkAPpB7Ta8nGOWT/9VHASaBFgSO4rt
jZGX4BFMER6aBZWntL5Eoq1/Usj+1iE9M7QMlvMvvGHtp+WPbYrLNrj00LJRLcsVr5q4TMxO/57j
6xIgQjspbUpw+UoMgKJcJfWSejWI9dJhQ6oIlI5mCnevWFgXqEGZNtVvJVFGRmCHRTYrceiev1m5
qm26his6P/Zk3MN53QxzxwlK3+JMVWNRgHUmNrdwC1XNGzMEHEJOnCyX+2h+rHpJeQzWaLvnx7rp
UMofIH30quH+QFTbCKySpfNzGX9Jb10d8ELVSfpG1nGZW5FlxeVdEPgis4I8wf+bDiAT87kjWEZb
T+qnnvbtTbQ7pqgwCQpCXnFxJocHWZTZNh/vEL6zPOjY4/vjsUoVXic5GOrOMM2tREy0c3g1fkA2
f2dr2/W1JAz3sqEtXRleYAwhpyvbeLMLiIg5+lRzaqVSD4jTxfAs4bY9G5KMOaXvPHtUmceCEXKL
hPxmSJgAc2QBCRXw70WdrKddAUA55AkOoBjAdjzXH14YAQiU39FjrvbohjZU8PSox+gtKEHcAw7Q
YidntIEYaVOkcFiHUDQfWcNJp+o+8+7JVIB9YHqk1yWOYm7b/3naDId1AVBiN4X6b9wVqayB/Lmu
ZamQB1H4jVWiiKCwIQ9yihz/NQ+4qTDK5YjIQJjktGyD0LPjbb6Ue0UDGNNuAoMZGJcXl9KbweFj
CPSVzOSPeFuH3NVrSYvEfWJD9G88L2JIKzHxigq8R+x2rE3nruRx1ZZVr9CVi1iQfBmjLjUyg3/6
oK/TgqIZVwnuimkkaDe7PdYAZRdlQF6PUiisZsJyRCf3y/ZNEsc5kZn85VWAlgPKHpHMTDGkSUuz
mSTLrU/NrvSwfzlTvce+Ui2CzBZ4A4lIyr1IbAHjgagRIqdsMndt8Tmq0ZCAGcjgJqkgLv0sbYjj
FqksEM/KMgcM1O9QIMWU3oeaR+Foj3MiKXnoOskvLahtDqB0zmt9ULVrJpFMj5c6VwFeLAcb/C8v
sOxAW5xNtn0jimy07HTKU1nul/pvcc0cvKvmL7GXrRAW0kGM+Zy4dDv/1EugzcJlzZTLO+yhtKDB
kLmCO1FUAGHQF47MtfZYEqhvGZaWPA4w+dExU5WFS5BskmWy6oTC7Vh6idQgYUDNcAjTxIpUmJpL
lbPLpkqI7WREnrbANlMHWBaOt/Suq7Sdl0RQ4l1p40pCG4buwfbtsowQsykpVBzKvRESUUMtA/2y
oO6Zq6q3kKhRuZUwzs8Pj/7MwqbyiltiTI+IAgKnNmdBG3MCh7e2Nzazo9594CLKwZMZs3IhTAbD
h1Mo4mtQY+otBZgHlgPTEGq91cl38QxCXZdOHNBnP4jLx2FRakMpUrkxVLBt2ZzL4Wnp2jcrLesm
KJnyJavLXfW+hM2TbtIlivPdxy8KzaQFB5s+89gN4fh1LjORyPpm2QgI+U02v08PbacH5teRPHWJ
qWobEjedfPhFxQoiuuWt7TzMeGWNDB52x6zfk/qyoUy1hjyrPtnEb/24PhuT4iU9WgnR9RmTu7MO
Y80vTTst9p0lmeRbcm9v4ZNsaeNuROOJbOvajjmMg9GAdm9pD35wh4pfOd973wQCKwNQ3tcNRlKX
5Ra0ogxltWyB/oUlhVQlAi1sBDsh646U2znM69/UOu8VGn/KiXjNWVqe9Z6M9L+sNifeZH6OSQxg
Ty8iGYn3jgfjRvu2P7Pa+nsm0l7NNKVz3zFY5p3isqoiwxx+2wl8lwBGER0fxTuldWIyXcQu3xzF
ZgJmcUO1qDKoq04SrbOZniPT7Bm5WvYETXXAB5AyzGTG/JQrAdKNLAVL1PGlUtolcJwUxH2dkYPV
bdx+ZeJBQZRZgDhfv/9Pfe7UJklsOMB+YB2ayOyAfOZKklZ4EnAkd0aupWLyX259zfVcBLCsY/Sj
CyIJ1h/YTNI4viD0/4tLTuh54V/wMCoNXNa8Kl0yrcjOl2dJdmEakWuDvA0hMHIb+itbqwNzeVls
TnaRzp8fPaPqhwzescNv9vr1i9z1ht3Gx3vwqS+9FYpIzUckVXn/IPBHXBFxop9p3hAU0Gz9xTcF
jvm1/s+0Zvc+oOUgGJBwBLnXEHBZFKCJ+i+ECg1KN2iM+z6Y0bT4HYjyBsSkhuwTmrMNPP/Nu6k+
XcOulkCmMh85icc2Xs7MAMnXfxlIM8Tb8eSTBp0c4AUvn83sSLnugpMkkp/Qsjd0oqUXTMX1uPPB
UQxrQAGFmH532LMEBpCX7Tnjaf3kdmGPuvEW2GneqVEFCdOnv50YBXpZvqkb4I2DlMxdc70dbHjV
xkB7+V26u4pewWs+W+qURGJuvSxZfji5SMP0Qc828/ISvDdb4M/yHPiWYmShqT3Ds4pdU4Xs3nub
fEhh/T7ayo7aJF4w4Qyc6r4g0+lMZ6FrwCKLxXkdM9YVlJKZGRYvIdq+f+HvO/79yQtURiPGggNl
ZIVU5EcnQoucseM2qPaxNEV/1C/EUo+9oLO7iZqizoziEkxQ99qenueBBLyqtIBlzu06PBWLCeyD
EjA7huXyEUZoxrtsU5ndi9UaMT5u5EKrKZun2YkXERE4s+nUMENCsUhqeLaTJvBUHQn5aCXtkHZW
MNEUZXbs4HYJEFrpXd8uCdC9e/r8yLP+K9atWYk3r25ZSz5NMrPj7ZoQAPbfKA5Iy3p7jDJs1uXJ
cu8spBwfVzUAirHxxb6XzIy4e1tJ8u1vuB/53cC2L7knYvYKgcz9Tv9uJLrOSnUsMJxklgl7V/AI
lxqQQALBY4ypwuuzbJVLuwTk5+5XgS5ErdUdiqZxvdkhYlZ+irBWpah9Icl1iahk+LMK5UqDBL2X
hVLAqVc6Jmxg2ATuLQWmW9JyWjTZh8pbzgdzA8Wi05KRtvXP/wjXqGByQARI4RUx04Rkpf8CUz8C
gr5w1mthPdoTcAQK08eWrAqsW8YPyEX3optNIQLGo9beqPKlXti1GC+fH1rRGydbKYlyBR5p1sqr
Sn+l61Edvbbr3wQ2nkPEhexToXy107pKDARiNk5O5mZnmEDQmDZUnXx7frQNjaLlDf+ccoOgwEvC
brzfMvSrYuTQLH0BHlX/dj//0CJdyABiRBeZhOI+5t1wlVzep0r7Bnr6D/WsgGkigNXVvYE6N8lG
aSlqN/1xtkCCmIPTEwgB2DuLTCw0LrvYp50wOl3K84LZZIe2fE5jKY6+++ujpoaii2ddgYNsvjPR
8zqFABksJLWt1KeDPnjfXo2JFJqnbS+W562+5tRsxsmfpxHyV0xydAgBfOUeY45ykI7N1e8K6heG
BmT4eTOLro4RIr20PUAITvdnalnE1/jVCELzIBM6v5w+DRvt3r/rCWzqtBouO8mfIe9D8xHyBkkL
kNh1dayLtVDnhBMMrLkzOaiK0WfHyaG4uPLbWsHCeVvcDFUpFEXVtgzzSBx77hVCaIhi2QnixFed
1dsuXgS9qqRHlB/dS62n/BoGDLfW6lVxhKjjQNKqpFzUMJZci6l9IDXJEm8mfnEciHdiNDxlIT1W
MS9sD4VqpDm6hsk71OKlc+UeoxOig+EDSf0adCrhdTIsfI7icplW5wBCKUaOh9NqkH20QuJvwu6j
d9yxolb42RRMfPpHK7sNfPzVxUkX3MWUYjU6EUSaCx6m8w2Z6dHTqU6kxmxhg4Y7blvXA2L5ULPp
W86s6yKGorofiqD594ffl2+Rs5lc1Zw9b3TPVHZAaE0ALR2oOLI8ZFPDBtTDrODJrg0BX7zoYQ6p
JiVN9PXqy0ZKCEaAOLwJO4zuCr9givETH64iz3hGCnu27l2qrzjXwmboxL6lUNuovp/m/mLnO287
Ghd3uaQ53a6o1i6doKDX34tM9I60Hh3o9lG/ldk+8dHkrXpHm8Hs9y1VkZYKVOuzFsCUSRx0xvgp
8H6+S60UCO9y1H8uUq3vylPV8Cqk8wMtfPFrG4rHmSP67muVcuPCqYxKQsWtceY8c0x682wKt5DZ
QFErEGCLj5UdS/P5eOGGxoJ+InXnb6WFi3JvpcjpsPInObIisIp71mlwlUXOQoNl9siSb0mZqWaM
hyfn5Esq+UOuPnnqF/CML1E/TzsBsX33NwRHHxlph4ICzlVMvTOAlZ4TJMCJB+l4n6FtKTTnXHXf
lVZ7kjvA+1Fb+BPgcf6I3giuTPjfMzkIilw9s3f3hMebupB625Lo9y4eHLVK6ngB9g1Jm6jREljC
sQJPB0Z2/P8iSfk5xALFnyJjl9VOYhZGwWkkL6cftmJWDv5zefG2jXsoEYzPrffq/wEElDypIWGQ
FC8Scph5/MxOAxgMYEXZB8mat1rdmYcJSQF5Nlxr1aguYEDIatU2u3P247P1qk6cdlO8abXI6T3R
Cq+PRHkxH1PUDU7Qxt8ap2YMEeamottowoIx3xGF2XsyjsGI0E5cSqh0DIxB1utudIMK7xSe9sRi
EW69kAJgj75AYao4w+K6KoSlwVstdSi5qUIgVHrYzFxz63SO6FxlkiaXvpYzUdBCejDskczWBDb5
HwsIzQwWcPRYO4TTxnEf18uXXLYF+R4ZnaEspHA95X1IP/sYL0fYLa7o1RSck/6UdXDHViSqD9/H
IaH5xqYCxXUoXgYYGknEiPpfdg3l6midbpXXpICNdWOFAGtCaWSRf1+tX6WNvKRqzcQzaJd2/mZh
muVQ8WMdy32Xvfci9kRBHqZ2g5iqipMIyWx3BsXPK5Ox50c90Nwc+H8ikw9K+XNaHjDBRso4ja6r
f0Xs2R6bzNSUobgVA1Px4cO56GnxSmcVYLl8pj1c1TPi7TPu6HGxN1E+qMW2VACxfXoMtdDL5JSW
rEIEmJX2yHn+G1+stWA53s0IMvr66HH/FZwVN1ECQo75PKjNFFzF28f04aDNBGx1cDpysKB9c28B
J6dUwGmrJLb/kWt6p1XI13M7eA9oHsmcmUWWvosuSKGDgTmDAQ1e2/NaWpHFJOpFzZLPpRsicB0S
jQOsaUFQ+igTg5M46dVx4EW01WuXVORwLMhXdEG/ghT1xRD7nQYzMzVyaLBR3dPGHDPdMYja+aqc
+EfgsqADtdyQKhOZ0ZPafGAFrEZxiwQvy2jus0PztBsn0/XQrHk9xvFxNvq31REV6qOTs6aj9aLs
8I0D9fNm1GsZejOtZrhmT2sToxYcz4VyXAr+uIr2LiRtUN1IdcW1sAbjyjaPkmx84zUo92S0OEs0
yp9Vj9IOPJwGDpbtQrJJa7bdjorgdz7TuMnh4xyHgS6U4v1+Y9b6zIg3cBjM3JvcK0ES4sdC+8I8
Vb5Y7OdJKNVkrBN4PPLS6vExnI7AdGpFvRG2QCq1XOpyhSKvKSjRH5M7i2wmwrAr3B+kbMFlHJ5A
rATw3FR2JJECXXT3VBC6slUWWioNSoRPVUkvpQb0kSZM3iyNjwkPYPwocAD79D3Q4fnS/pjivS+N
bwgFc+2GwsZ1OcsLKCJOfNdrMAUPxUhayZLChuptG5WysMG6vgvUcxXcOrdzqOIr/BOKxtX/FsB7
MwzUK5ZK6YfrhE63WqWkCFkjS3ybsJit+uAGTGJDATzOVjGFPjvIdAIpZC9ZSpgH0HSCQDo70M8i
4pBsxAvqOi1kSOI49lE9hTYC8huI1I7tUPK8sLALPm39VW+q9c5+p1QZQNl2CPuDgumCMTZsrrqk
9uQGbhQfpCKg7z5yHQkduDTwmCMl7qj/3tPsRDW/ilxNo3LAT1KHLy0Kz6aKSIhvprM68FNSHAC2
8NHsq2ZhYVbgG0ugSo7T/RWPD01xiqFchHyT3Vs+TkO/GhWLTO6ig43xhlYXshrJk1C0RBWSvkTu
hLXJX0WgnO3f/H4O8C6ANUfoDg2N/445CqJIZvGNQ/kMYbLCVg0pMFdEU7XHfuxXHkvFhkpErSlX
h+B9fwGc2JZANcWyNWNzPYalDhnCrv/ZJA8i02cR+UBcjA5r+R0Wk+M9TkShYnxuwJ2qW5eKeqfS
IiiR+q1qLH07k7i49lu+0MJ8Qj5giZ31lSuoWxHpANWWO7loY/OY4M4bDKGhDr7qkYSobKxXff+r
c/IyrZivXT12okjoE6wRq6AEyawVt5xWOu6nkr/vWVIqP2xUGufo85ndDXdoN3q3QKeN6QMxKaFL
WyF+LJF6l4HUhsa+aHIBpDOQMNKPk+0lCwbneU0nxcQC6WEU3g7/6/A1mCKm4QdWIT1al2/OZqRa
sbzdrArGiGv+iQsxf14McIde/6sJGwiPlZJ7NR4EoKHSYeY4KusngYscalvMYSkY/gMb1j18MDOJ
Gf3bdENScc0wdSBBa1EyUxpIS3ojxWPzXYX6x1oXnQnKC8O3ML6ZaTAqMZSYATKKiu2ATI5yjxnW
Bid1nfOMelRzfMWnuikQUBTmUrAgxgg9buC77u4sYaBuSLFn4oxyjaH2SWDytHiPME6HRnEjT6pz
Z6wzHo6UQV3fptPVCfUNqQFQAEh6gBrNQ79ALlq5MH9Skheb+MJ1rWMfHduTGXd7pMmbwqXHtuxQ
k9ckIOn9yzqn4Yk56akUGLyl/OGlwLNHvWLWPtk7BMOkwMSbpDcjACOZfTKD6n/4R7azWxmdyKlT
Ve8hb4Fsqh+TebSxls+R154AHJ+a0UvO3CorCcdyxQpjzLvQ4ki+lkqntjKnhN+uYBawPXEj8wUO
a2qkplMU3vT1zpu6NaBYq64WHKFdTLuOrbUBourBv1IwQ7T34H3x2jIY604GxkhrJ7y4ogQlnfmI
tjv0piWyFkRejvLci1xPTerOL0YMyJIfHWf4GHsDcq3k7R/m8BXAKVPh2j4r4JSwQNLyxa3nQ00s
AR57hX4z1jCmHH6nQw2X5L4XFEATKZbfVuKo8K8kqQTKwyj1cGNHDa8KpkekpGbjxdrp/1tyHeRW
/SFSYtkNB4yzJMhkk46/uzVwhM+87R8Tgz6bQG1+RquWZBxeu8fhd8rCaoovxWxTlZ/burl9SP5J
pzSgkho/lZwcv7wBlW6VRMnXETKb61VFdoLXi2IGBl9+H2pViFUcNaVY2xPQKZ3AgnlbZBDzNc6Z
tbx3kjm55sPBt5domAdySzjVgvB4BNhmgcSg106nYfizgRrrX9xg5lkcWp8rKo/xcaoIDCh/6NVX
nxx8g1DG7vBGFCMcj336LeU/ZjHQTB8hryvdeJj9jQCB5JKwfb4tJi5vhDhlF/VLF81h97Hro83q
G+kt0nmTvfWBqjJRKcmUsBzbBaZmDhLxU/qKjAVrsS0Iktcxb/6w57Akk4cwOnSVEIQcWrzh5ln3
L8pqF/XYX+fZ9c6JaZqftthDdz1GFuM1tRs+bHBtDtu2AEeKid23bxBUWSHYCvkGsvrb/GvEqsJ9
udr1xLSz38vhYS/H4WkoSpLOWN5YmpBYTqOHy24e/LOAqgdgstLz4W53qgb9vSCv3hxwQ1kU59tc
wW1cyaxZbItuEC9E6a2C0bCXxhS3e2NGefcOHNB/0p4zAQAkC3Ogiy88VvZi3SG4jIvEC/K0mv9x
ro6qTziOosIB5CONvsCrONVW24zPSmK7bMyxBegfkg4xVi/SIgOLxDHCmVIxRdFk/hlDFqmaM57n
AxNCkU2q+5C5XtKobGQ3WZhtXVJw2IgqwTXoUMeAuzCSnLhdHBwMQS0ffJ53hAVf/L4E1/sYalJy
NPbUXU48eBaHqXX0nkvkMIYkjduabHfhzvGpWAQtAWcjS0nfLpPIdXFtAmod974eIEqEngGeqAEy
nPzZhTzX1k4oNqvYBCEBX0KLp8AvDddjksfJrM7XqOeqGIsdkquNCmMR9ByWtgjuJSDyh7BDO65a
3dX87AwOqJsCi/mDIRGZ0pZ1pFs9U+4TuDGz8p8847n3rQMrvcJ7pFFpcZiVgwfOnE8daitN/jih
noa/kr1cK21K9tc9B23FQ8c9N/lSo/9Rls20IIYISjmNKa+juxVBYA9vUhDY9eyjMZgr1CuB9XdQ
7twtNbz3TFM26KZM/96SWZFzg4DyLArxKGChzAQLit6ucwGiD+MUL/hEf9llcrESuK8vnKWuGHOs
jwkUQWYXcCWqNzfAmuwMiyz4bFajmshKFPwFpl1UuY8sGS2NDZ/f5exk0GMs+h061Xe1R3SxGCaX
RTktCBjoXoT5BZ/CDr21/Fo0TtM/3hxkmw9/X0TUBmxZnCOx8D4xW+r7Mk2CmOOXU9WjYZOjrvYf
4UefYCjg7G3w6szT1TtFvkhZW8ghlENwJMxugZ4pXwMRIkge1KQSkkJ63fRjXlRiiGLowk5xAMDi
HdR0ejG5Ll+8K8yemO7RhhMCP2YRDzeEzKPFX1FMtdTmrxuVb7AOsbcfe3BYwDsUf5rhAbhUUHNd
fSpjqNuJfNFZengCFHRD825aixs2Vd0Jp1G/0S79DWrgvq/1treHioj/RsOrgX1GfXeFTch9MqUO
bOsWdxlqAXgy8E+f9GmGOFK07+iPdU300gGJTBdBwlPl6aTo1EP6MfAsKKScO9b3AuISInYmVB6f
oow6PyFVKDeXPOx3BAhgcgfNHpUJ+f7X5nxAUXiobTgXyYvQum27dD0qtT/8bUP+VABiFel4S+qS
pHkVsmAjy2kic6cPqIhJo20CwmZdTChtYDODbbaYLospJtkLrR+ba6kxgwsdFJgeVM+zRbbROxmb
oFVtkGW2KltvaalQxVxxhGhCkRvjY4Z2sT/fTFh8tWGWT43DzbOjDaSKKFyeT0s8qIscx1ffgGBY
TDQbtuD1Vvxub7SCWYCzAH65i7ArUzhzs7fZ8HusaKqZd+LKvHpyNRB6Ikokv6BuTmj5FXWTb6JC
JVuyNT5B0buWh89TBPLL1/wO3/9UeJ5ZWPLZfS7eGZPOgE5ehLNNZaynSw9hinTa+RBYqQCSNW1c
pwEeKEeVRXEMfRdde5cku6Vr/ZvkRM65oryGbFGWWw1upgCGk6becN6QcG6rZ40jz4aGmSipgauV
2H5+xb7lgTZnv7tS1MrKZ/CgQQktyWQOwKYqVSvLcAsiUAFYy2LyP85HfPpuz5/hiy6ujxoFYXVG
2GknCf9koRPH3Wuj2uv5wqQ4Q+0XWuOktrqkuM5p9Wr+A1S5vIxCH7/ZtiFVeeEgv+lAdfRKKuJc
SaWdQnE39nSQ02XbfYmMjTEB0yV/bdzpdc0R+KOaqTnUACElj39Q5+Bk47kVfARLwd78qefEINUt
EGcnbhrBqXnIRLlyFVEofJRzToHkKAgu5UQ48lXT7MoxlJ2sGDhVBR2cCmsoTgSvhnoQ77DXdUzf
mesSIq+X/6OMaMqjZzus0ffJYY1Icj5AVXsdRCjzHgEJ/KmLmi4qHeSQP6sqlDHBUvDwfl7WE8pX
ATe8BuZpbQD6ZjqwSkFcsOEjS5YmdjHmlaUBFuFHZdB6QmVlpIyRObs1jtCgcO2SPC+asGS3KlrV
wX/IMm7wwrHUc7T0jXC+YNGs/RCiV8HCDudayE9wLC93TJRE9i7YcmVjZ5gVE7FoX2QvMIHM/ORm
/tFfjqxvZwuQimusfdTITFxt8bwu3F4VK0gQr3NOK8EpifYkl1W48AxzpBhFgHqtKZGbCOlNMrHe
RDawacSd7C4Og44SyUXIOSQ33cbtPtxQpK0wTZd1mOP0q1iZzxL0R1U4Fuo8H5LPGdDoxIX/ka7x
UfOcPslN4FSFLZI6UXDflJwD1NjRNBlg0jVIlAKqLQAeqPBdF2WeBSSLFFqmpJ5FKylqNZ/rwHDk
f54XA8hTf3oHaY+IH/2LI/LTu4lWNfoCXOXNazw2Eds30trE9rf+NrW4K4Cnodit/JXMNrXKtG+M
uc+EziAiqhjVhY97JboR7Qm/y9YicrJ/XbGBNfrSDmv0noDflQTt8+DwnAxN7CPNW8IYVAnip9Tf
msC9UfXLx1VEMKOjwU7aiHC3VmCIHvoRCg/aG5Lo6S/WNbvVd5q+dJpDeoi0JUJEUz8UJuBTPl9x
t+WjCRUwkiS8PK9e/1vczeGq/gKOSsVqUiRi/NPYukXrEq29XjquoC3ZhK+77kyHWEo4kpqYLdHZ
9gH/1cNHoshn4Wn07NlywDXW0biKaooNq00P+kscci6EwuH1oKTnIjLkQ3B1y7lqyIB2o7AT49L4
jdZ5E7i3TEap1kOPVHg96tAp2HeZMs5H97PeXMAsbWwegZEIrRQFB4hKb56wUVJ+CvwAnRjlmmnj
v7qWw/r1+2B3NOwaoAm4ibt+y/JsNaoly41WOwY4JYs2HWLxcVRrQ2eHg4lYj9jWVPKkkXIkA8UW
DOHZ7QLWFx41VOx0PIieoV8VRVOb5rjhVYj/vfy5llpQpbOvMpkXcrgQ5G0lnsY6ib+mKZJxWj0N
1+NgfAbGGvBhJmTnDIT2Nhbpt+0GrTpC2t35hzgNMAtVhQ/HDNzI2+swokRb+nmOK+3s2pNpPgPW
3RgQL4UbMbmFmGzMWk/eKO4dTejhoP7bCyXnK7tqBzNQR4A85qcyEiLo8vYPj3/NOTrHxZz1yOSG
0sjvaAkIdMTtouKuJSZGeDN8IAOlHuS5naPVXZHStSpWXjm8jg/AAUGD3Jbt+EadC523b+R1nbzr
vwzUNFDM4Qp6trv1hpbfWP0qC1WCWM1lwnxOzbvjUGPbkCM/IRBW5rkR5XoalBr34dZ3Mfh+lKIw
0R4oVERFkIU2dDAnQy6ZadiuxzpluxjiRYiXcdv7ThHZALs5iDqBXj6UUIXV/sb5sbL+9rpGhfgM
44KnyE2ZlEzd/lneHiO7sAU3ahEDiI3Ek7uGiPx2dtSo8RcZIJBAr/aMd7t3FwOtj7VuD89RDIPm
GY7HwHj4jzvLGfIC75vOAZ92FC8M9xcBxvUbQhilp7NPgft58UrABgV9AZfGWV6HiZCsevbZTz3u
l7hYWqw7ISRVptSNAuFqFXWFXe7oaEu76b//3Ql0eYQFvnDtkz5Dmeu5vQ8Sbz4FHvF++Xymp9y4
ANlpuBAsRm6ccGt7idUitgyEw45dO2pX2sLvvr+S/S6azRuOX35vpD09VBHauO4dlLQNC8tl2D5k
WXSzQO49jjAhuXNRPeB/+eJq4OaQamoZAZkJDADzOfZEhbosud42eZdPRpRs8KAgIGa5bP2wWeAA
+t2akAG8aKwShVhGEbzUtLeFE+9BtYkC1c70bJQkNVmZIRKLnuQ2xOmS7OJge0j80sfKigBiVf2L
lzeq3gEMV6cWyeXZkNh/H6FoudCPFNT8nYnnGmn7bAY3QSZHTJsaHHbmXWjlUsjgi+GMnkh4YCYD
Thzf0Y4wOhpHI/0CCJdATOaLAkk1lEYqFYefOJ1pBF+5frjJ42z1xfUkLKnbmVmhEIiaLnrSo7zK
d5BrhhVJ8UqY1+UDXBF1lxMapIlgbjFqm+O6JU4P9fasi5ECo7yXIin4g4mgvihWYRFJvgypLvyA
B3JH7LlnG3UpabU/M6yb6EGI+a0syT7oNK23BsWyzAYARVu1spiwyDQ+g/zLMBzwduzm9aTlIkqa
qlBWa1Tbbnjup9oORBd/XOUt3SKHhpxLKhqtzq1Jb2BpTUjBEotiVh4xHFmb1jTVJUbOk5/fmG4s
rT3tObAPp6BX0E1CPkx+/ykulE7V1qk8fwT60sw+DT3+rR7PK/V3yPEiiGoY+ifDKTiDafQDhhVu
Sso74d9+ftZueQCsLgHzDdGI/pT0LjpMnyvWzPxTszGHuUNqU7swx2Ac6R5OT255Ei322YFM/8mK
Jc8Q3jg6sYUFyvD2k+C4Xt9GwCpLK/3vHuvVICWHWFNSOgyfLm6TqSwFcUobDHqqGImsLeaRiTi7
D6L8RzaFGlQgM2NCRldPQHDld01GCku9dTjSnMrq1m9nDPkVqMuXVZJVnJ4DmFLqfSe51QVixCPP
5jZ1qeushgQMlWzYuOKiwe2dMsOCrfvLbK7Ef2PNFlhw8dpH2i491RrWj5Of1ZwSOYqn9hapRhOF
ptVc7LKG1q2ekuHSMjwWxSGCoBdXitTV/t2gT5Q92ErcG+ox0lUERYjBfNgfINxQdkB6E2GbHI8u
QIYDhgL8Roy4a0FLFJJiPbWtt0js8I7xyKm9ntYkrJyA0wEPKvHrpnm80z8W0o028/MtQchjhRdu
0Qo7wBIqXU8GbUmhXs68tyVrssHe6eyGW1YcE+hzps7jClI1OtRQHg31Nicoq+IEj9lDlT8X+pcF
69xXBDpgAWb8Q6Bn97V98/EY7V9ePv9uoxnRIvdKBys72Rvpx+0/K8AdmBcplQH3uokclAAdJXyG
OhG135zslvkAk9vxo868+x8HSQVrHFRMdbiLB8jUwGde+uGSWgKEFWfKuF00yTVIBfpU2RDgUNho
0m8n1iczT7jKtbs3JAtv+sgXGNkZvBb1IPuZXjVqrLI013GbPfF6Qespemw1RNshagJ5MlLhOgdu
57fbz03M+BOtY4qAFkftmSvVgD/zVzejz1xpeAGVp8jiz0RDbemIB5O8FsZF3sVQmiKcErePsQU7
n9GeaZ9C+2QD+sPK93EqA6Ugw0wjYIu0Xgw8mZg8Msxi1D2UUmwpa2o83pyOYpB/FFQsxXGvYBqa
vQPX9uQ/JI63dFCcXRyEMjafC+5F9BbXiFjO3jkBLFDfKb2CjSV5R/UjPHdbW273mfvbTaS7y3mm
k+rwd0kdKyQ8x5bbTaIxQBb6QuNJvxdRIj25woMX6ojc5QOUKqgrsIQNJxzkk9iVP75NnlUSfZi2
3oWrPks5MmYVuzrwciKiKcoFDZVJWeVyrMpuVWvFnbQ+pTvmZVA9VoFhXzd9UU7FydcRRMdkvwVR
h7ccV6PvYUIpRZOtapOFTqjQLbNui2HD3sfuB8YhPoBMe3s+K4ybvTAUtDpWEgRGqqjjQi4GCbht
BjAtOgv5Ao2pMVeaG0EKoD4KToxtry4ZA5EeU2DttWRK+JBhcJn115xdXQZTlXXWX83FM+4kGQ55
3RvyyZFgA00qOAPgXcVPxguOdxo0awJmw4tGOuR/XvajwAK3oDjZyBIiYJCbvJjaOeWJ9ZJsLCAH
RX34VHQJcNhLAmJmomMAdxjRfYu4PS4ojghk+gmkVu6IgvvqYcHbqvdq9jYqKG7O4i5CWrOv2GPq
Ze5rrtHGxQCKYWt926JsnyYKAcbcCSXlIhnlI0uZ5ibolnhrd5KeNRIpKHjhkKGhcSO1ieTwICVA
eQ82YKTx8j18QVgB6CYVk3Et9gA6xg51dt0OH6cO08iwVjCIrfojSgCHhNKMqbS4tNpXvk3JmBA1
jUDfOw3kiqN7GzdKaoB4RA6Z8KbmrwynYy14L8AUf8ikH2U+0VaUk/lk6tIafvTPhJrjUqTmJH4x
z8cRfs/7pc+5KY5qzOC8rJRbS7dZFscp6lO3CBGtKjmsKI2nLFe2n1abn90rfDTZBqTFlnTgd7DZ
M17RexM0Rqyib+ighRd/l4yNcJbHibUVPDl0kNZLrGs06qT0mPEqKauBHcKhQwHWfYvupV22d08X
D+8OMVCSfLd3PdFC3QzpQUjcZqfiWfgAShuMjRPl+l8/QRuqc53tbRG7VaI97lG5v48rekpyFWPR
vmX/qeCX+BvHm5oiQj3WO9q775BAq79shz3/nBcecfSNQ0VHA0uDPu5fhUzZoQjPhnl/lY50KxGF
/79xldoucT9NiReaEDlET8AMe/8TWPk8/Om84O5gnUPK9BKtLuUoIDecqFYTT0bHhoe7+OMR+qBI
WEyKTcghBlFJ2H1G5ZYzv3oowb00zhsnEdrmGRtyvAw7f1oeT7ucIENNhlbsUjmVuX1wjNa3CkOf
KUWHF1PM9rEJfBqMmQco5jVwJ7Ucy1I0HgejJOiPaD/5R9y4rUieEy1whAYb7SYxzv/luLpLi2KQ
vU5vzw3A6CyqdFEajK2fokCjUhPZF5DB3ssAjxQtzD/WumNLNyTZAN8Q1XwhH5+CUmEF3n+OiM5a
X69EZ3w8wKSacBsWMxEJ1kqHH5MWn50UAE90bGufffxzBGoIyJUgqA7/8o3SklAEdoz8vXa+cBv4
RIoISMlR0tDYrJaHfhRLx8rze0fc+7zJZyvZ2Hfy625TJZ8rHSGmSDIJkNU7/4UZ7FqX4vZB0chF
bnsDdUAXQC7+2xnH5TMUm9MX3YXAj6nb1nqWiy9STZx6sfcdnLGMyMY/+ZJEj8Up/t1bVxm3BNYY
tmqmYUl5mY6wbtXRir0nKBnwur94aFW27I+v0eeK88E7GVyEhB7VuLWrtQcIY2yKp1ywK+LZ/rrt
sjbwDQpp4eZiBvawMWU82nDsJgJALclQd6aYvKR8etPdvkWv8/GSjjKxLScNliTg06qiCKBunBOp
iKED0yt0uZ4qwtiS5dASNYuvTzNT1u1dk5G+S8pWr/lUiqRU4eXEmK+g+4sKRYySUX1EkKM8TT9L
dkgX4TGmCosNRu0rrJ4eL0NDG4vVpRSvZhAXj25YGUaE2o4q/NOdt5VTkLvThkpBFmFJqI6eklW2
WROJYDtRL4cNR0ejf5Wr3fa0kAVMDFdTt/Wl0h7S1vEppmWQVy6C4+icr8Tmtakdu4zzHvByNUZH
OWwMz9kCz3UXMcqbIz1w0cHEZyrHHqbOQHym81TdIqn6F6D3u2BYMKMg3XuvIZNNNelupvAt3mHM
ew9qgAGv5mdYSpXQLtb6S1dbi07Ta6Hn1TXqXj3jJUEHDQNCt4HMqM4AY9Qzqca+bWqrsud+cKee
k668w1xbbgX1Zq5N96ABKWcCmS6UPqmgd12035xhpHD6UKRCRsEf3V1EKCxagrHh2j4JI7c6SGUh
2or+EEPY0H33WXitfJ7njGID2y6qo07OvUDh3vsaOKg/wCx5R30YtpoVBo00uwC17wK7Mg2rFvuu
bnDiHFefFn5SVfNvZhA7ILIfldFAI7g+38g7IGWBUpX7xDlcnibxOfJgrdGJsB01LVTPuTRr1ry9
aduFnYj/ZXGKCZ26n5O4+vMRN1+Er2iDJBrQtSWxid05TAoGFfgawE/6lkznIko9zDwZRoXil0rm
b6/HIV1UvrOtvZIWGD2LKARIlKFmJuM82ECA6h4gv1jSbZJHzaFlce6sqf8fh7dMk/W752h+fGFP
0KEvBkSiKvhrC/491gwA6rbJUSKeHfHKMVEtEXsyqEXncIgB55h1HkKfRCkVWbRDkHyqG3uTSqG9
ssF8FaNz0wcl5f78BYmGPIh3UrNg6v4MaFwkS9gPzAh/UtdmcEH3fPM5a0W3uKVopLaA/mf0WLzD
oz60P6wmRh6X0/jJEihrKBvQWMRNruRaLvbxTCA8xQ3s5G4yBy4t1FCTKBgkiz/xEV+uJeEckDZW
ZTqssvdDZyp6he3YZsm9rXeGTxY5Ai0JxCIcg0Zyekf0yLmg+5j4JoNHAeZmwlkUIUu5XPfCrajS
FeLubgBgHdRcJTgCXnzESkoeNZDNkFE+LR3mNQdMlc4inJTDJjuqFwVkhH8G34GdB0yLuWQDHGhr
NO7Mnbph3jvS0YIhCFStGmXF29NiTZKZECAk27XUgWUDAERX8GgnrgLgRcLPak1qeO7YcXMRXGsJ
NSb/Ss1CcUACP6ZLrHlyPU6wb2JCtjFgswWy8JIWf9KKHPNLqb662QPVBh7oA0SB+GznTtC84Qoj
zpzqdh6QmGvA23rojMi4JRBo+eApKTSuLXIBTmyLj9mjM5d0tuOr+7kJiO6ZHZkfv/PwVjN1Ao5n
PYD++CvHdZOmFtsL3RuC8+WN3VDtpSDr+IVfx7EXAYt8/B0YlC7BI7VdUN0lNdr4WZX7Q7addcrc
zgsgCYGPpUPjcQ8vhY0OrLF4nVGL9GRKzFG4kPZk/y1gaRixax2N00mVw32bufRUgKpTIfzcC6hU
MZbsj1v+1Xfo6JZ1++SgIe0oGrLN5j8YEq7zGIAl/sVCnRhG937uun2KodTmcwtBylkZQCo9sGsL
g1/jum5cnBpAKMP7JePa1H588vGzQvaWnoVjag4oH/yzWG1e5BjsPitjJrUqwXkrp+fyHWtx3sHc
zUUoePkxbdYUxhsWujW1f06ppkVk7b/BSLmiYTrWu6RgVq+SfodlIw2VSlS9uYMZyFgthfzEybRk
k6tsfzS6wZd6oahxw9uH5EplBoYxT5dNW/N75LEbW/8kowlQEMrIX73/tMYLm9PqXfByhQ48uboS
13kE/MYUzooGquZbFauLxpFQDtx4YbvBDs8ZKusOVc1zL/9m5H3rnyWhw13g89BoR5InJj0EoYki
yeG6/3+tyfx9n5JKfTPZ4Iw1vNg5xH7Y2FlaLAYbuqY8ygy1CNoHPOhkCxCROzy2MmpDyNkaykb+
Ci06PBGFh7/EQ56Ru/tCgnfR/oEZgZP6RjmJYTWpKti2Nqj+gqNr68rl08WlJr5sVKUUkiCrpInY
wsSO3f0NPYYleDIGeE9ABMsg2yBSCFryv5k/ruPUwKDUhZHgmjSq6KFCDav44lrYeqSJlQYVXYw/
3RFyrePtu7ut2IOqAM9IaOHPDdHCR0KQOZdSM/PBgc2Wd7S5BNRI+THOq+aKLQfqUyfToTbZS/tW
pHGWlyx8qA1HSekRwBNaOoSjRzz19Mf9H6RocpU7IarozocvOcnbqv1gNcwI8MVkUIMf0bt1DbUn
X0t4pb1qFeL2IZKwpURiAS1qh42e7uphUkkUiva5/KVd5MaX/N2a8+DDzgfS+JDZwuem97hOiVhM
xsZ7rvsrAuG0G4G7qfkFXktwZbZgVMq8u2ktTUx0Sg+Ie7ewIpsxsq+1btAHReMdpppT7o4b4ssC
OLy02Bg0h44yb/WOaaHRtKBsgPAk+i/u2wx6rZMmENMZ+PDkH1RnSU2pJFKl9itUyxPJ6/J1o1zA
jnSvA7t2qoQ7/IE13F6T7dQwYKfw95OBf4dmN1KqObgeGmUZ6kqGXxmqgTADz2JuUJyvJJ2gA70Y
wI7GesGZIYyp9R0WY2Zs9fb/qSA8l74p1+PA23Ozv4IbYDpl9Nf85KYoEuuVPFnQVq25A3+oEfS6
KxE4MkOetXQ79+OlU+2UuCZkzPbGeNr4eEgjolx67qQdCmKTRaSSg1P9VNPgnE9vp/23D+GoebLo
F6k8en7aCm3SUg6qi1ozSFAkYU4dweVh9I6lO66lXFbHbOr+nEXso4rjUJXR88OGp84BEvw5OULd
txNS9u/F1V4snoo+IyuzehTTjRvLJ86x3FrHY4Ahcx8NkTKptciuut7HcBr6rROriTKETFMTczMR
1bLuzVsgm6ZI/XmhS1NiKXHQ2DJLGGAlSFfrYpVwlJ82pKN7DjiPtGHKmmel/XOioF3F33v8gQsS
B0LWI9nCZfNRoqGQmiIT26/FHxvOI7YXW/BjJ5NmHwOkylooeU8gm8ERvnRJfW6AhnFEfLi1WmL0
S/zycqWg+qGQ4G9mLH2AB4/Diwhh8V+TpggfnxFJj/xD/Nwv4OeRC2Dup6N6xKD7RCcRv6iYF+BK
mZwRObEAv3iQhcZWcic1ORq1+HFu6eiR3QhHC466tTftjryvGwiezUmNMsFz57Pd0V5LZQEGaXdB
Vxlga+Bza97SoxvEIX/rTUJyfQsGSqZEXahV7XXOYSUSdp3a549gjY2fKzu++jmzqIGeXWNjxqmb
NRyzO6O/Xm75TYeBG1o8VtPnNyjp6avlMdDsJtoLDl1afdbb6sh7kdM1IhwocgT521fR7nPBz8Ct
TYTWhSKz2DTymDAEMmGRDQ79iDRec5KfCzWD/74vnf/y9DiN/NfOGp5WeTWD46inzZT4594SUlV1
xdtydG7rYL8qNuLyEiHMLUhXEO9vgwaQxCzA7VYylEWY1Z3ea8sC4JOgWIY6WhS5RlAC2uZAEvMd
jSjWYyDZi73UfN+Zk7VnR4j/qI+f+3c5pAa5nERHy8IflstY8iLzRaXcTGOzaypQr7HPRFrhl0Mn
IzxYJ/vRJAiQCBQs9D9ThcaMJW2SV/hL6GoyKFijjS4DIHzn9A4t4PiAt0BqfcRBWUGZhOVjBQrf
lvfKa8CqZ3WSp6Hu1SjE9nzstLgAFXD493s5Zm3a/glLq0dpIa3+bwAdjy9FTk86xQREzrONNHGm
MZdHQN0AeFIpdMQMahn4wluqPVrRu4nndESdilO1ARDEbx37WVIrSmxno5TayLkGooV93MHYzN/f
xXGSzt6zASXul+e2NP+ASPOIWMyuqDDFmHeUVTu6QmQOIpUYp0ewmkP2PeGffJGpijd+QfSSPKtC
1oYl90YBp/N0UHuV4NpY1Utg+okgNcoyz5DfpFcvtya3wzUFQgaOSoVEgmKie1QZzZdmbvgOLH0h
WoZBLRdmQ1y8WWGd8UYeP5bLDepLtSqiSUBGDJycs+Mw9XdVxQjLFqZ59IGguNqRn1vyHMoXuqzV
pfwBAuAuXRAc0wP0VJCBkWcrq3kfU06Bp5xfWtf4sW5DMW74get0Kme0+ziptxZzroDNZeO5ruIu
gfNvuHBk2uM/3ct23QhC/Y6Qg1+Wpzby/tUmYDxsCkq3++kSyPL8YAQCej0iwxdqc6hM/C7lvviG
B1Y4d8nI/R0o+p9Nu020JEK/pgqZ5O480OCFU9qBlTmQsW0HZt6zI5WsMqMLG0/2TW7Btp6h+AXm
Z0E/wChtPbe2bxB8qkFsvna0XXImqdk4y0NELwaj0r+hSsuJoqHHcq65PVXOx8uAZy1ZP5UY5l0C
mvFXsUcXOwOZomCqj8mZJphtJnBZOHjT4kcZhZmfSF6pqSJLSwEWosksRcEwPwUCstGOqy9XZjBR
HJSRr7jWXtP9WYMnxUMf/PPXHePXdG3jbXk/JoWL5zTkSAe5AXJobdDNnDoRHrCgZMalrblZwQ5s
hefln34YcL8q7t5iWgfk7iK1rJ6CtpYzdFAN97wDS0UjanLBX08B9FCiQgfgq9PkpnDxeYTmRK10
vneUIa41blTHIrGYZVxFbmmu3odvTDZFtdZMlfxCMnuYGP3m7uZJyUqmp/AK5x7Qq8fxXJJoK1ww
zAw2hBzDre3oev7ckEKFMqXCAorAmKPU/aey6Pgq14MUew3U9yDFFbVQcKHiLRkT4mx7CEQL/ePC
gcBVlJcvo85l7K/kjzsv7hVaWkNXoBhPClsnmVnIiXTKHshaIimZzAWx/oqTx56mt/xG7X7HRTih
Vbsi4/9eMrZbh19b4iORsRnue5XTCdjwMejCKayc8Q2DaCzBUrvIWUuXeR+2YdQ4gPHabbkobycz
zCXme45f3nvxaWaAXRDiAsK+DyQ+pG7joPnqNmLxeQk6Tk+JWgyrt3ybKL5QqWH0QMJbD5DCOq4P
EH/GaishgJvNIkOiEBd6yDqDUxcClt8njitKHjoSWHKit1VknkpY56y9rFQywGJkhypcIEm5gzH9
FnZMKo+gF0tUzx0hLGgySlOijNwQ/yV2RVaUYKjsx8R2VGocWem6RE1KEttxuoF9duwUQ6xdWE5H
6WJIHxgig+L0wd59bYMz6rspiSvHFQtuEvKkY3HQPzfphVuvQBoeiTLfWL5kVEnpNH3MRf2V4EfJ
LXdoRCDCgXQWDuk5gMw+hPR47MAvWoMSMIwbXPlmUZJE/2D2vMou1Jr2cBSd0e8+l0A/st7MQg6K
e+zD+hyX4jmbCpe5ISQ3G/FCFEBzR2AdDDdHweU5RlN3zWBF0jMY/V/Z2v2gK4yFvZ+eOIq8R6tL
Kk7hBAxrs5/NRVVLUc0T/7ob7+Y5O/C+b4HShasQoCozc20MyB3TvqNIwrVwDZFAu8Od5ZfvVEAe
6bON6yJ5oCiU21Tu0VVGjWasofaW4a7ogs0o79Z4RsPlqK0LAC8CBeoS+m3cSMxZcODN7p0D/6G5
Gn4Pxnjlr98zBHRdhjfEt/peHAFtthZS78Efi0cerkLmRfpkhRI8S7jGEO+u+eGwhtuKv8WlgGfA
cW4TBGuvV8X0iH/xOpWUSarO/zld8ZNtBbJAugh5BxRqlg11BOb8HBsM/DEEHTGF/YRzamnBnvU9
UxWyWV9EEOUoj0dM0fjia50lqflbqZP+/wWto0pVqtayzjOUukfN4eXoWQw20TK/KTB1tE+3v7sW
zm+9S2/DlLJAMCVG3DjIHHMNYNE5BScQ+/gWhlFVRuQVX6o2H+nZJlGCLJPFhU1+0ap2zijCX7Pp
PlpPF9rMUj3YAvuzWDrPseinZVGQeYitGOBS5u2Dzxvk1UY27aZA7os2EzLCJEi/pri9OezJBJsu
nuD8o2ojslIRYMmC6OAvXrTjbs+1/qAJaAzQbh9tExen3/1hdSNtEEvqHlFb+GsK33cFx21fJUbb
YNzpgxRG5xfSgjbC4Az+sZi9gFgGme166W48dDU1QxejzFL6fH5wQCHjTwjsEJzcMrXdIAM7PIQT
X3YJYeFiKazLfrUGaLuuniQ2TfFsLaSibs2U80O5NtVRzHO1D7JSIG+ip11doFtk7BjvUHEx2LLe
nSEcKxmllzM6mDMq5GrZyXfOb0Rec9j/3QRKLWey9Jugdbj4t6DKVAxaQttImkw3swUTo0TdfQhm
gJE7g8R+WGOU8/IqPaJcZB15CUmrgkzfJlT8Yd7eOOWYqzMUOPsJFahc6txrPYi4CHuJbmQ6ec9J
8unvONRAFnpV9hJhsOfyA1TIx4hwI5pdjrOEf+9ejCuTt0nOjJp1ZUKO96lXnsdqSgzX/f4U0dHM
AlrtBlhcd74OD5WDbwSZY/ddwq9ToJM5TwCfs/RGeOaBZxptuGrZrRfLwiu66VU7CTLAaGDxe7w6
6meSADoMqoDyvsk5fpfeqG4OGcabErwsoWDW6tdZD9mgL58LO0DDHZ5xdL+IwqOlB8BPVldG/DdI
8dFnWmB5/T9rf6aVOMnzQj7MIig40JI6AnNe9+sNM0UxxRVokWQbVp77SmbQkgBRM545rig49X9C
yKoUPMxHhdKxMXFilWd/SgyXOL8D+Mp+huQgPuI5pl4IxzVNm41WZl1MLyej10a7PK2/Q2Y0SHOB
P6OavxMvpueDGRdFI/yDMkf7qzz8aHQNGkaFBEBrcv4i/0xkHelW78P7R/iXo/kSUOITSQtKb7YT
fxGnuOoR/UKj7ALM1gAJBeadxe7hxNK8cMSZ7DIfaRUKKuc3TEuTfo4v1VRmuJi0XBJEnZrQucJo
xME7SGToV11jyx0lvFae+5KPSmQbLu8Z1aA93tw2w1zakO/FGiC55ryYVCKlwiUStCMYlAQe12J2
SwYcYBBTgoKSFSQH440iAVMd1PLnC2yVfASa5q7rTKSTC66C0jDhv4YkUtXkvlWBUnqv6PP6xkbW
BtTnTd7Juc5KStCyXeUQNBIs2jneIu5z0SlzpEsjT5jLmnF6DbKW2/VmrswB/wok6+IwZ9omblwX
mzifXJi9+EiJegmUrjg+evO9dC9jKXcR58Vd8XHvl+ukPYw6AGXc/BOsMYV2UxekTz9JkkRZSGmt
mFw66mVbXgAAqIfjb1fsuQRbCHk8rtrL2tBC2/cIuVxLARDBKqRc39wUtv/E6Kfd9aLjyCVJFei8
Q/bxEPGQrvmlrcY1YxFlDURZgzDSoNnSR5v5Ek4xXapTgcyj6uBr2/iSWP0+7C1G0X6jW8RsDmiQ
+gWr5+JVQxz8ZWlcopvVc4CV5dfxWiqzxSQfxFQwP4LPwUsb1fBc0Pv52ATQ/ufevxQC6uHv0zcI
ep4KtqhRC+NSNuznwdAV7GF+yP6cgL1fTl7u0vtsbw1x4fR781UZGD8hwrPEFStG9wCgUn+kQtuA
+j4wmRi9jg01RWl5ZZpJx99Stynq4u7agj0ymlVw7t3UZCXfrhEANO2BLisINMaojQQg5AbFvmUf
UwLfjniAPwXZGYK16KKkMzn25FfapUqbPZ3GOaJ5coGSi6tC6bsmuhAvCl4+vPol1IkbNCKvNEES
nXI0V+9EqdJ2W28okQit8mqrnOXDFGcOXYfEsZKJ94D8KHXsOY+0pun2kSVQ6npDuLyru6tNWBo2
2AqSZyQ9gWpIRwCgP0z0xSO+Mez2o1U42GwGc2WoLvMOlmfcTazOJOdxes5K56OTRV2MUY0Hdv2q
zlNp2E3Or3axhSjA8iOZ0uu6KO38RGOqVqiJbtK/tCKFGv3OUL2tvaYjRq3oa6TNi9DE+JqbaFOh
4dusmfeTPNmI3P7WfezZqp+NMQi/NtXEXn/VHhk06yyyqVRttLzl5ix1lMDFtqjZks2sl5TCtFu9
v91s2g7pvTA+DfTSI8UY/DubaynoI5njKBGMhvG72vxkbDYj4lkzftgVAtu0gnfrLirz0277SQmW
nv1+4mojSq/rwQBV8fyy+WWaVgbIJP6vln6vS80JB/g5kz4neVOaIpihD7SDcgurvAi4qV7Ts1g1
ZGNA+YU2E0yrtND4iRkfAXqySeet1xabkiH+8U8KaIKS3w+MlPt0WEkeGMYBPB/DsHRE74tt7jxf
kbfL6IuE1sFTqG1vkuu3Hbb8M5emHjS0OMhKXTjo80EHqdYBAcz/GJswtgRVccsEOXDXyCFzw0RY
uLVur+RsnG3ptsD19AdOyDZOvPFGiA6/Pf5PzxHn/Ordynro8LfWjlfl6sipPZesiXKmA/2oD/8P
jgVQKPoyLqojai7zpFn13CJARH9seye8TMgJbBHrqFx7xYgLeepuMf3TE6SnM5h0v5xo2LX9jOE0
3ii/XZ6qT2OQb/GH3pYJ+1izROExlrQcHX7FWxc3T6QhqHVeb+0iUcBtFO2WHa22GCkYE5rCKq3B
F9ct+UbI9StVVNTPNS/+KGVA2AuedG73XG3U79mrZ7/wcYIDnJpH9bNVnfJ5vq3twttKt1fucozh
hLrDvz5NvSzqXneC3sUQ8tSlexqR1JVzs0zqP3oUeFDD7wOgLkPnFz0Wq38PmRZQA2+R0gtZxfsU
0MvhtDN/lBcXF46JLc6UTYcVbzLkt0+m1b9qM4UuWTBL9Wr9jxCgqDQ7cfOKc2kRVj+LFNv9UU+D
5rxioN7fVCgNweR7itUqo/nZr5TqcPbom6wVYFRS9y41yerA6m1N6VjwLgdozn6qTipB9Pns/veI
za20IQSa+DJytclOgMkKIMgWmfTTd/UFJa3sX8KTPI6WUVuxuFMI9nchADWR+JMGPohamXNe3t2f
AYTk0WYOJLuEtBCRXLcLlau2wqTuvxoeuE7CME8jHMRBEFTNb6hWvhm99Wci5YpJ8s5Ksg8ZiXvf
n/RV3wEs2VWn34VUZ9sswzI+pUmaVPUpjQWy++MsbklC/FMNDZLcZZarN0N5KoXcrzGeWiJw5f6h
RS/hxB1Bds98+9h35QEvd70O7zAhHM0EvK0wTrh+5v7dzElG50Ed7mN3FfBrBxLAqd7fEKUigtk+
sWSp7vemBlkT4qTiIEDzEvcN02FbP2fB82TlWvn6bj2el2jZfDb/huSdGj0a6MAzbIpZbG/9Ka2g
VdAMRY5oL62jrWakvz63RLijRhs12DLglsYJpctQYjRYSA9wmntYh3pjjU4OzWw0W5gY/fBoRaQx
o0cgWPbWQMAYWr8dW82n7bU1bHnyYVOBe04+jb5s57cYnGnX8aVDkTCr5Z41bDDhTqjITOjkxHsu
WsbpZCAzeXG4wK3rXAY6Aun85rK3/cYILyYFXxhv/zq//6KfuCMwked2m4a/GzqWknVi2xFs0a2/
PyZ4YctRVjqdG9TFWAD/S1EqfkkU1dDRXw886f3ykHv7wag0liyX/1lnIM4sMmJrVS7RNIJpZmHn
ji6PM1QwC7TLnNXOr1LA2vS36ODEP9kmqlrI2ccBgnAEs6CKfyRnfxX0SASUuxFPp6Z0yqqjShc7
nNF68q1c2ZcL8JLRzewc3PO7Sh97ACYDU9VyDqw8DqYL8fXfLAftdOXxZcZdok20xZr6snW/iJOB
zy0JH6ryRzXcIZk+LDoJvYLmogX9yLIkIuKkN7/wK43Nj1mcsHRNgkxD0oAooyUQRiJfPuzGvb+b
mwK1i2yJAx9n8291EKYycM9Gg3CmjcBuKsmg3xkj6tzpEylvGFog6CSaEOLh/4NT25eE59CvfdT/
rgv2TjyQ/eLw2geKsnwvXjUEqs4zE5G2wTqx08w0sKdAzRF7gZO++nljybk2xFwqUppz2hK1ZP69
Q8WlB21KdNYdDJaGV/WYQVhsTv5el5ozeJov8rIXAAa6gdziftgT0HWHQymlZi64raOHNBSQD4OQ
aN28b970Zui+7sb2qQ8p2zZDOL94AjAYExWkfxhowmIxQtWLFZM/K1FJqXAcOrAZHREUu+HTbLu8
mSDjhmwLIDhUls50zp5uQvgYWw0TiS34/1xpsQCphJEr405xQAtx0RQQkaBS/DCEIxuVl5ur2/7c
UZG+shSfTMPFplOdYGA7FP4VhrIFKPX0x2CcdnbBkYAPMIF8GzbWQVLivCIYIkxUjj+hzjp/pFUD
31Y90bVyUIQM51fLmKWfsEBNkBMiXAQBaKksEHNG6cNcZ9FQtg7YrqG9sGk5j5LZidiwj+pWYAKz
svrLixiGTuinB4rD2iWN5PhNoKWn3nEQfpRBhTP6YFXxZlyOIzTsE3fDvn3XqhfGMJkxhZAdKc7H
uT5vvT0+OWVsXOnhiNQxeUyEZ/rIqhJLhN7sX5TgtYDEsvLg5WPYWMZZYhV8LYpV9iNUO2gOyKyJ
5vCwJh9iua1Tipb5Ltpk3wPgUr4HvHETSDl1/zz5xir7+cagFhJHdcZKht9RIvhxzQFb/e1gkvJk
wSPzJDE+xNXs5KfMFAiMbQqpJFa3XK2btyidl+bQA9srVarNmNtyqI5z6n88MSDiHDGuc2MqTjh1
pe0hIxKucwVpFrPs01I9kqSfIs7UxRm/ePGPlrz6tZWaNaUGSyNGVW4PkRzY3Prs0Oo9j6/0a6ij
l25wyRCq1yMz47T4+Dloo2VTJaHbVWBxvkS+nWCUakpmJIZWBlPcF0IUfix2q8CyN9OIl+tVNqzZ
MXv94Bl+mNG8INxe+wmEnE3t1MNqoY28ICVdDBjNYZrqDIr7sKnuojHyb8mPDoFCEZM49pSdmdKs
yoJqLkBNW01yRNURsCHkdwyzlAcjtGiK19nL3e69thZCC9qoPIzQYUeOvofgED9p7SdoG8bN+8YK
5nCMAzIixSLB75qy8ONsVp2QlnMqwYn/h5qhn5/FfsJM63HRYjHik1rVkQbSXgXdrl/SoJ5BipVh
rU4ZaUEmQgujmJfdYOZYwXqPbcNz9s4TXYdhiGsB5Dl/1be6H5rt0fWeQES3AHo0dseWZEzP2RQw
okQEZeBL8LoffvH+eKVzmktqXvfuJ0NipO4d+N+5mp9GkUF4UJt3E+7x0+p/P6CXFkBFt5xdfh7d
YeWZfClMpuX/99EMkLeK0ysdU0qgEsZQSVKtXNsuwlzfytslbslPm0ejGw2m7fDmmFsui07xs/N7
yTFCwAQHqjTwUw1x2TtlcxPVEg0tAFQed7fvow28KptflI9RwcwOQDsVPLy7JVhhZN/4casDpNJu
BDAa6qBRd9Q52bINK1Vx5gQJTTny/DCsNz1hpmicY28x8coHZtY5sN86ljmsh7pnnuesYtBoXjIi
21Q80uWA3Kp8eMVr+RP3TYFJ5B7unW5EZpS7ZqkDAj0HnBF0wL04oWkEUxsxPn1IdQW1+nKm7E9i
jsANS71Y05Hs4ktGA8I2p8EAhd/L2/gj9ZBzQHOZ6PtQmUhz2F3VIB7bE1WQevvfRxCC/zlE4Aqo
ucQDAiPTD4sTrwoOUhUORNr7VgXCN9fWLpWJGCXQtYNpmeo5ha9nKzj7zQPnJpKZI1OfM5XYl+Xj
g8X5DdwA+eHSQuv5c+lC1WLu0rMP+31oiyBdyZkIfgxM6NllPfUOObP1lQEr0unPDASbnB189Eo4
NEH6WMGPY+APTAuAHkLgiN/y8+eVm990nUbaKOgzO/0zPZfoIsVdEUq+Epo5drM04vcwBl2TaJRk
6SVvA4byqUsB+bQeEGU5XywqWCypnUlazhfrOocwlx9P5zkmhBrM0L3/3c4a3+9fR7mYCA+DyToZ
Nnp9rVPchO3AEyz5WY/JK2t3ZuKCh8AzHTDlwXnCBe4ajEBv7JSwpJfz2Rtp2tk2uCyzw0cQryDb
xS/PfQBCepsaYs3j0lEZpRvpPe3tWDubnkHhsCVJt6wa/ywWxAm5nMQomuXZ3sip8yFM+jRGoMNY
eyKTkA9wNGK204srTg01inHYMIIUJ9PkhrLB4hcR+JKRbqwOC89mPhOwdRlrv0Nvp1zPFvdNxyXX
OtI5SXl9cN0wK/HAc3MDLQWM37huuAIT6zwI2Bu+aWsRicRHzmDWjew4YOTNI0et0BSCI0BfkGPJ
oQpUshEuZHrAXwI7UBQGiAuKX9mRHdRkYyMTzFLgSPxUixoQspLeurl3BOh8WXdlnnjy6IrtjtJE
38BusOnDAPpbWV8PdBLhQOw8ZpdaV1+pDdLf3iNoeyh3XDzWEMUe3QtOjKgytYv+I8LWhJOONVJa
zYCDVHPlcnClTaabEg5QmkDYTTQszd+DhB/K0T81gAauQwt1skmQX8g+lXCMuGYlg4fYjLdkWqwg
UaeSkKPvFU5VRYIOSWPofB5pb26TwVyedZbYHQcgo3hHuc5Wmf08XUHISPIPceMB7pR3x6y08r1m
cyGJXnn7C1xsiLpdTHjJdNzkjE9KpekBVU1pxWeBwDZvLsilM0oCtlKZ9nCJ0CYwNZdu88tbCAbo
ujtFD/N5t9Clx0crsqJDW5P5GuwYe0HmpxGmMod4YPlAN+22W8r24/8yGQQGbwyoelbu0FmCFTDN
trd44cL1LQoG/t4DJeN5pOU2NQNw0qE+Ip0Q
`protect end_protected
