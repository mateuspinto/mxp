��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���Y�oV`jd�#%��B��"zK%�L_t��~ڮ��O�o�4�9J�R����:�H����w�V�� f0M�|�(B�1��lt�A�B*c�@�΋7�}��b�r��Z�J��y��?���s�0z�~ �'i���1(êƥA���V0C�p+��0²��H��8��A�y\4�p��<��2�r��T ���K\n�a�J[Z��������1ڪ)O��be�v7���������=�b{'�r�1'�ר|f�H�m����x�9P�2����wLO�� G�%���UV6�z�`�pL����i�PQ2SJL�F��S�8��P��Ry�2�?=�kz�g8p.�Wo7�JMǂ���?u8y�g���\
B��^0h��C#�yN3�u!�� "�#�:�)�_�ti�W@6R`��=Ǌ���iI�&��ٶ��Om��J_X�8����*�]O��$#.������o8>��C��3!r���i�Yޥ\��S/��{�}z0��H����\+�dQy����Џ �`�*.Ed�̥�������Q�RǤ���g��� �j�3� >σx�͠��1�2Ղ���l��a��d��o�?
R�c�L���?_[̦Z��;�/>�;�����DSd�����d���P�2��]�M}ı����S��qSO/���*}��]�e��X"b�Iע����f�(��=�jx�YY���o�	3L��cZ�T���#�;>��]mV`�?gc,����`��l�(�Z�``�`��$[�n��#�PAH�K��X�+�A}:�yL����A���!�ʍO���p�]���c��&�o1���L���Q��4f<O��%
k�G��@�B��R���bm�f�h������-�3GG�b��hOl����	#1�#U��)�d<�3m��p�Ó�}�3*�jc.���5�E"8W!6=
G�E�������[�F�>��4݉P�� )^�"ox���'�MV���"��w�?��(L�W��U�)��K�Z*��\��mx[W���p�>�}�6���3�VF3�@�l!��IVMFIL%�:�z[p
+�q#sE�!<��,��u+�u��tF���M�AS~��_������	�-�;�ʕ���T�Q���X���yB��{R���ԧ9�o�ޡ�ax3��` IV�V�^`��;��V@� '��-A{�D_�ܝ��9bI���@�u�����gCb���[���Rz�}e�n!ql�9byA@�W	�i�A`'��<��� ��Dw،�POM%�&������I�k�)�ɦ���՛�`s"�}f����$T��b��B���� �Vِ��w��o�.�u����]��F�hXf=I� �BM|��fH?�����i=�I�S��c��D�"5�\�
�LHl� [*��Q��]��=�@���ސˍ�4�s�#-�,-��|�-���lJ��iJ��Bz�����ɓ$����g��)���ޯm�A8��y��ң��8b���4�B��تs#�u�������h�=)MۤxI�6F�i8<"�T����פ6�㈹��(���2������.���]C/͋^$�@��gL��4�����������/Ïa�+�[6�T#cF�ힹpb3�و�������λ>�K�p�cI��u@SV�a֏BuZ4ݎԘ��EZ�Db�4� ܁�Ww�*�ֶ׺�� �o�����)4}�ب����� ]ı6����+��K>�<B~��<'~�!P��ۋ�ka��\����2�Tv�E�� M���1(g��#����&��c>�q��g�ѪP<�Թr#�ӱ/A�+�z�m�w�L7w/�p?�S|Qzjex	�}��i�Oz�¯����8ed��[�v�j��0�HS�j��i�Ԫ�IIP���[J98���!�F!�
 �S^�Db%��8 ¬��g����������S�M�N��䗂2	��-�n��M�Q�Q5[�J�a�m��`]��~1�pA�!,��F6��Gm>)NEk�Χ6��A{��Ԁ'�C'__"#}^�n�b�೿������_��&.��R�����y��M#�x���:],,��W���}�M�D�!#�"C�8�F��9B�'^.���`R����+���
H��;��KW��BFG���o�τ2��g����c���rQ�t��=T˒�kI>�X�'&pT�`����X�}>��Ys�`4$x߸c�&G��>������u[/јKF�oY_�_�/J��6����m���Bc��߱Wk�vJW�Sqܴ*k"���-=��~�+�(�v��k�:HX��n��+�i-8��K�#�L=7>3�48o�]'찵�����wS�C��;�D�t�ùc(��)pA��q�1T��U����k�K�i�0�=b�|/r71���e)(~��Sѣ����'�=,f��{���~̯�8�z����b���(������ҔE7�C��0��䖱����Y�IgzI�!�y����b�>�F�~�D�W1߈���$��&^y�^R�Ԛfx�ùD���
]_�.����=Z�>5�@�!�$�j�������f��{ t��ɓ�<��,q1��zQ� �Q)-K������OE��k��/9l?9�.!IiKY[xZ6@�0��mp8 �7�kA���>�/N��D�tߘ2�So
<r`6�ɻ#Գ2�g*U��������~�����rBC��Z�wŁ� Px����ؠl�-OQ����%�N����ɰVg��V�0���I���+_$�������;ӱP �eJ�Z��x�N�z�zܧ��l�{p!i�y�]w����R���Қ���/P��봡j�{��W��V�� ��x�������%�&�8(���`$�	����t5� ��Xo���z}CG p��e�6o%�'�U��Q�:,_P�����z�z�0恩�������/=9AB�*gF�>�_>�u7�@2��GiU�rp&[�zH�c�!�s�` :�U܇s:7q�F�� �Z�ϝ
/4�Jcۤ�
��2��@_F[��כ�ʯn�b<|q���}�:u�XZ�9�F��Uiz�����o'�D;���;.m)�[�������!����3n��H,�!Z.%N%ܣX����D�q�$��Y�W��:m«X�g���EVSѠ��ct��>�_���\�,yd냵�-���t�l���
Χ�r�xV>Uc���Cp�k�w	k%���!��F��hi�ē�Ǵ�:�qU�����rh��(�阎�M�~��;+����A\S^���k*|49�Zj�T7���/���5�_pڞiͣmp�� �#�����0�����A����2=�A��u����b����\�Z�����Qo�?�q柘�@杔x%�)�uFZ���FG�p�?A�Ҙ��lv?�6�WvC�D����:�S��6!x'�#]�OG!�~x����_�y�:S� ��$�(�:���t{��g�#&�����g.��s8�G���s���抵���� 6�-�7�#��-{ހH	C�	\k;�S=t��5o M���%d��i������l7���FgI��<tOBNl�Ƴ��]�sD�>�CΗ_~�+>�7�C��Q�k	 >h7e~d�|�$"�4u��5N �/X(�fk�-�;3�(����]��D�Z�5��ͣ@�}�r��]���
[���N��l��fk`����_�K��Nl���ES	=�nd�Rj~&��5A�+��\Q��;�G�c��a&YMʰ��p �/N��	u<&3�AHE(�^�X���,l$D��"�
����Ɛ�k��?��TA�XJ��y�L}JhŦ���PKYc(p�	U�n�S�;/��H��؀32l �E|��C I���d�����+^m9`��J7SD �0��,l7��b�`E�X^�2�0��r�e�m�+dإE�r
�κ�ތ��8	�z��}�\���O�kX�wA���՞�_&G�Tvِ3O��2u4ҪpqK	�צڭ7m���q���Q1�	��F�٭�s��|]^�Y]3���}Ó��.D=}��ϖg����,׌�t��@�M�'Vg>�S�Ļ(��t|B�H< k�~��%Pb������ߓp)E�-��7�<bW�T=0����j@�Bo���k`���jd�Z\��ѓy�AxB��
�n%���̲��4�Eu�g{[�?��DCC�T��I��-��f	�.����?�I�c��`�PwKKyT�MC:��f�"����/	�H��N��7��g�uZ�B1�e��{��ݭ�q�,P�j���cD�n�m�h���)���%xY��`h�C��_`ꘗ�p;�p�V(ϡ�ӿHȯ�+�	7)o"��R���s('`oz�� �_�������������D��r*���y"�~�*�=?}:��$0 �I�{n��$3_�% �c�G;@S#�b��������)���p���5:�v��x�/���}5rz��&��d��6��6gi���*��g�iȹ�jB]���B������CA�M��GRM�é;{Fd�����,?��8"S;��|�Q4kȓf��d7ñj���PQ�������  tS�t��V2ܿ��j�ay�J��x� �p:�f����^c-ڒ=�BA�ڮ����R9�^H�>7��)A���_�����륚���IjǤC����A�S3�B��>�ʝ��x�~�	o3�� mP�W�"b�����jS|[�幁�dpj�ä?硎��H�������{��5�?��2��d���qc<���K�-A�*�8u�dx�YI;az6��Π__N�B�$��d��'|�S���1�]0ѠXS����	�rVe��5���]>Sn�.�����Ŏ��?k"�i4D�Pާ��2*�"��`��h����M��hy�t�S��<lo�H5��R����v����J�"1�#w�(��X[H���N��e~,�q$5�ic�o�bI�##��h�����T�X��\��D��Q��5^��j��š�C��n/k=�RS��L]&���,|����7,\^%.��Y�d�ܙ��d+}2}�93���z��vܝ�e��s�v��'D�d���P�9\��M/Afj�a8+n�f$1IZ�d%����)T9���i,,��y66@߀�ּw\���?��!*ivĳ�E��LbB� �'�ؙ���� J�UݔgN��"�s�@�B�+��f��4�%000�^{IxB���L{_Q��d*��E�e��i����`�є��1�D�؁�"�F|}4:�<�͓5Q�F0�E�{pq���ٸ�|�L%�~�a.Eҝ�ŃoOf�@�K��*�![H1�\n�(���({ס��n4�m�|ʠ�l��Q8Ѽ3�K�1��|]=CFӭY.�(@�ߕڴ��$JOW;�>Խ_u~�V]�R�z���|VMp�f�ڠoQ�
`0dQ�*
0�/�梬�I���9b�������T��ؼZ:�,�*bJ6�&N���A�Y�rL���a��4r����^7G�P��2�e�9s	�z��:6�J�uu��\@��� �Lw�	���f� ���W;�7�#�5G�����	�9z�H�e��[i6����޲��q�d�K�,�pXsq�O���6'�t;s�q]UÍ��?2��C�됗�@ѣ��s�����gˀ́��y��W�@r�̿+�/�B����Wݐ�|�1j���Z���C&��Kx��7���V��D�*�m��&�u���b���Q@P��m|�����w�5�[N�,���׋�V{���Z�&�{���1#f�^�DF�g�%��	Jn�I���V=�F=n�#�C���w0��>�U^0�_����4���]�b�ȣMΎ#{5�2�	<1$�9cF*Vb�Bޫ&��X��|	ͶI)���"@�M�(�.A6��;ᫎl����>��Bߜ;t�k.g����<7�&l�u��]�̺&ӜI�'��yϺ�9�6A$����J��,�1'�D�		Cm��D�(=�;�t%	�׍@��M[��"���f�0?��(�k�QTd���G[�<_J�����&t�l=�iٲ�t��h*���D�67�^���o��K� r9[�F�������h�ͭ��ۚ��<�H���7�C��cD��r0g�ov	��f��{ҋ��[�42q{�O�0����m*�s%�4��§|�����/֫���F	t��JH>p}��r�����΂� �C�p��E�I'�F�Y�쟪S�~\7H�~���F�O{1��qCc�� p&U��N^"��i~g0fN6��D��@���������em�H(f��X;���£����+t�Y���Wy��B�v�B]����.9<���b����<m�$������. ����w����(�ي���q2XK�)�����%F|(��B-D�v�CT�L斑b����P����v(l���c[�&鸑���6 {��!�
'C��6�h�Ƶ+���j�F�u�vn�p)eb��-��W�(Q:8�Wʺ������x��vL��z�e*��]|]3�3�&xʆ_��u��\�I���@tT4q��H�K.�KY�j��c���\��JP�hS�s�B��@��ׇ�����j°���\wu?�|�`� L��|�GMg�;oMd�9�y����=��V��3�<������3p���#��>I��;u1}�΃�S������*��G��u��يӳe3���3 6���E-:��8��e{��o��@���`��f�RY���-�V5#ՄM��O�i0'�0[	���G�{���,]O�  �z+�n�P5�UV.�Vȁ����N�� 3�v�.D+�E�Z��5e%�Ԑ.��|`����3Y��Ǣl?�E3y�qDQW�[Y��os��g qsP[��ND������3��[�݃$"=�w�
�u���A]o-�gK�h>�܂��f��,)	W�h���֊N��\�=��%w�"�X)]o�h�q�5Y�����@�՘��N���y���XI�b����Ҍ9��e���`���%���؋�~��Г!��ҧ�%���`)��X�b��kH��;3��Pͼ_x!���S����O��S&C�C*�&Xo�k�5��?�k�S�4�"5���-�sh���$� ���_7O��������~�?��{}҅ �(c�M���P�==`Wc2�{7���s��l��!�6�
sD����xH��̶�IW�1ZE4���Q�n�/`ŀ��E��wB
�j$S@5��y�=hV,��k?�8���J���Ԅ�`�3����m[������A�ӓ�|P7w-��"��-赹��آ��v"d�JJ��=�%jX3%5�
8��m&�Y�����O��!f�K�M���;*�r���a]���{�X�� ���2f_.8f���{$I�4"3Lx�ʆ��� +B=Mn/ą���SY��� Lg��b-��;�Y98J��Lr�H7��~���5�X���k�LT��)�^@^I���_��!�z;�&���ׄd4_H}|�/y�������ߋ�a�a�t�H۝�2�q�Z��g���YYv � �a��'Z��ܑ�!��ڔL#7�R�����@%Y	B.&Ci�{�	�>�)����G�x��>Y�jj��~tOM����\��-�������w��A�#�����_�T׃����D��?���� Mm��=�14�^���9Q���c��&k�r��%�7:������47�e��n�4E����/+t#�zW=�&�o��0�tf$�*nnw�=kl`w7?(x	��v�3���M��k�-��ɇ��^�i�T�����7�0"���0f����� ��uP�	��kܸ��H�
���;7F�%�ЪJ�e�{������K��K��?E�xy���V�k@hd�D3�ʏ�6P!��5��Sr���?/�����`�xmy�׼���鵗�v����YE�.��9���2�O5��=��,M�>IJ�JJ����Q�ˢ�\��1��$K��_�f�`�%���؜#Y��6܁ۘj9�MM�����:@��W9̸t���`ߒM]#կ:�*AcBQ��ta��װ��aƆ?r=$��@�~�g��I� �qL�d����"8�r��0Yl����>�(mH�2L��˴g�(6��c�{�'�t������;�ۜ�S=��&8�]fe"I���M��W��g>��� B��t{�0��SJ����a1�Л��S)�G�CP,��ߛ|X�k�8/�E-M���!��`j���NX���AF��Q'��oaW.V�<��A�GH�bV�`�kA�W(h�W�*6d�Q:�����jY4��PA��誄i,���S����Ǚ�� 0�t���:����(]˺D�TV��͵���4�U�-�6(I�c�+�D��kq�#���b#�%����؟hY��vG�_���}˄�+WU��ؔ�_�Ŧ�A����]*B�#��@Q���U�ӧ�-����b�@��cMY�Z�ғ�M��_�8o X��i�xZ�����F���[���	Vv��
��s��	{�j*��+I?I�5j�a)��F���Nb.��IP08\���O�ѕrF��΁�e]6ҕ��GΜ�٪�f��O���O�(��b�v9�m�W�9���<���aj�u���s����;��1e��%]�A�"D=��%����Q���N�&� x����J��l���? 2��I�����@Ԃ8D}8�M�)q�>$3�I����e`R�jd�k����q'D�!���0jK`���i��o�F�Ϫ
y1�l���9snx����d���dP��9.�e4|N4ZA��HƯ�����9�HM�	<,ƒ�=1cY��Т's繪TIT_Qs�xi�B�8�Zl�\�CrK��l������,C�`�i[K��
0V�T��ۑ-���KC��Ҥ"}"9����Z�e~�D��0
��=�C���{6����0�8��s��_�l� �x��GD(���=��c�_���sZ�>$cv6��Gi��e��2�N@��\4>�RW��n�f5�<ҩ�m�ٗXK&I���ٌ�B�Qr��R^ �Z~]�EV��V��pWi}�7����3����*�)�7�oe������f��wHJ��c�����{���Jh���ce |ofw�LGe��)p��-{yn\���㞥��3-I}�RW��<�n�����p�8�3եU�^XcH��H�ub�W{���;��yaxIܧd9�>mw�]�	Y&sC��k�Ф�]���L���=����������f?�/�g%��`&?��:+3(~�����)Sz$p�����aP���>�!�.fN�+W@jޗA̲���o2�������?���Ｚ�(�#B�E��B�i�_�A%�f�	�r|��)Qz���n�C��*}o���>���Q2��f v���}����'��'�%P�T�^���ˏ����W����MV	;���u�7��pm	�p��ذ,��jM5��0�-Dĥ�����&�I�������T����o��$�{�+wv�dWBa|t`p��Q�#�������-����e1<$�1�ٯf1��PN�̜�kcܾ�{���쳣'����R6�\�PW���S~�
[l.C�}� ��?�g�D~�D�ҝ�����p�V�t�����,��S��V[��/�:�0���qY�IL�e��|@��i������ĝ�Ր�|���x�� �o���=AI0-/��V]
�r=����;qn�
�z揎jj#>�w��4�O�d�0YL_5��0�����_�\�wA��n��`{(�@�H�.���D�|� *�~���?�Ϡ���jj��2�4c�{ �����_����V����a�V��� �A��^��-����J�7��̍�n����X�7栃Y����	sY���p�bb���f� 5k�K�"�|ti���#��)�\b�E��$RԐ�ɖ���F��f��2�l<�W2Ͷs�V�^��u>���g��qӇ�۴���bi�R�t� 'Si�#�H�ם/[η���*�r{T��N�5W����t��ށ������o�+�]�KOךb;��?&�%��.�7�Q�99Ia���-��S��=��g�'kb��<<��b;�f��-���Dp�/T�,�Ư�}���ZSlu�*)g��Qh���{mz}1��)�z�\,���
v�s�r��%�?g�Ӈ�8wasc�s&��qΒ��s��v�l�Xژ,|�",R�|vd$�oX@���|JH�� ���g��	u>c#���Ha� �����0~5�a(��S-��hi�S�Bf���R�.A�S������j�r���C��zuӵF�ڌ*(��z��+-+w�(�K;<sw"2.���狦���lY{f�`�	�6�	��>�%�{�����C�3a¿��f�g�$����#��T��Mj�f�b���2�ʩZq�q%�T��~�n�Q��TbkVnFr��<���|V�-\{"a��zN�h��� ���Ƽ5�]\���1(��jq�8��.�o����˂�<90��n�O��]�a�j`����Bc��O%c�3 N���a_����6�M�P=�K�n��~��7��zU���|*�c�y$	�vi��[ш7�/!	�P�BӫPEf*�#(�>Y`MO>v5�B�[qF�ߨ磞'��v�'��۶'.�f���{��AV��c�	b��g�9+g��%ξ��#+�Ɂ���2�$\��}�;z�O=QE��F��`����{��J�4�K��rxf�׷�ߟP��9����j)\@Uέ˫�+{J��rƀ*�nԲ<5��
�n5���T0�0aKHh�� ���2�:��w�&Jwt��
q(eߔ$�%��cXiqػ�*��W�A�j-�e�̛��&V\�J%���0�)p��Qo��>Ob��ƞ%{��,��Z�=n�e�h���D9�9�]����8��r&��ǈ*(� Q�s� nmXP8�_k0a|���,�Ā��*q�u4�%�R������b#c+���m�j�^v?�8]��\�j?�&�ԛ�V�6�`�~�XP��n�DNt?�*�	�a��f�虖�;����ٗ�;��~�ʣ^��+v�P�#����dtD�B&���h��|�O]�t���u�=��:��>&��ώW����5`��)Y�t7��X���c�w\>�o�E�*�"Fel272Fi��~��J�Yz�e�W��#�:�+[=7x��}��'_,=d͡b,�<y1B]���0����6�o�U3\�j��#��+q�h���
���h�����>�O�g�u���Aצ��r��w<��DV�Э�?
c�~H3�J�z����_��b��{�՜��`9>#F��G�Ie���w�]J�-�h_�Lr�l.C(�5�<��ps�r�Eȍ�����CS�FeK١樃�D+�B��)�[�WN���e�T*�x�� N%8B ?��K��[F��z3W3].���f����Sbo�g�n�/�IAv&;DB�e2!�<�����R��W��!!�G��4�`��B�X�3�|��-V�p}.q�JT
=Sh�����N���2��l�	���>��[�J�q�fJ?Y+.�̃ �{+�:?��x'����6V;�\i�5�����ڥ�;�Yp2$ʤ��b�ˋ�;{��-6]�o�Wa�јKf.��ll��7y2�m��(��|�_tߵ��
��a��/��e)g90��3�u5�\�l��K�p�+�B��ESiڲ.f��*�`���.g4��w�F�����`�ϵpv5.��w;���Xv�}_��i϶*:�V��5U���� /���ֻ?
����.e�d������M>�[���ךh�GG1�I�L@�a�Z0Ͽ�FJ"O���׿>�Vj��ސꙋR�I�G��aB����x�ޫt��-�D�܍i��/A2�[4���Q��">c^o5L�,F�(*u��PK��At �kK�'tI���T� lՁ�	����H�K�4�q���@�j�$0�r�ȶ^�XR�L��푨Q��=���Obw�-�f��1C�-�YMR
}'�zr���W�YC�����u��>ȡt���^C�4_Ң\�	�.��6�}#
%x����Ҷ1�aS��������&�Z�{��q0����;��ɚ�x�3ӗ5O�T]K�� ��'�hTJ�M��f��e�3*vs��4+L���� u,����-ӈ����ڼ�{|����5�y�z<��Fnԡm"��~�];���P��8D�D=�$��q��6
���q�]g��Ƭj�w}i'�BT��Op�ᵀ8s�T<��l�zv����ha}��
܁}�c�S�u^�_HT}N�����9j��j�D4�G�_�~�Ѷ3���d �������0�k�A�N]/�?ԩnNّ��<��	[���D�y���{����>�!�3��~uk��+8�Z�Ț��Kz����܄O��۽�*y���ME,� ����3۟'�>�E=��5h{����N�~^�*�(�ӵ�,H��+筀0�*�|ӽ4�KcjH���@���7��1Dj�[rK4��A�i��J�I����ͨ���A���7���A5	��Z�]	��d�|�v�,��rS=����-I���B�_8���)փ���-S���I�7;:^����ܴ$wc5h�l�PSH���a�%ם���ג��iK��m���S*"�.�sm�Q���~�"�(��hQU������.c7�Κ�@؏@�����L��R���ݓ�%���-�K�y$�D�8��S�-��ъ�8�;�֗g���1��x\���u�?`��$�v�"�xi餒h���q�����;'b�o��M��x?R�ws��'$�϶"jI����="�DG�Ճ[;�T�� ��%I���K@��P�'�(w[��a-SF�Հ����g�d�hLB\��W��Q���H1���Ȳ�v�RпxV����E$��eb��B��&H(��SP�G��R��9w1�Bܵh0������mx�"�OR�o�rf�O�mc���� P&��8���xC��)x���`xw(��d�w�Ƶ��@[���N��߼Mf��
�!�;/�չ�E���R�){�s��yS��)�>���������,+�J�6�Fb�'01�T�u0��4zn�L�|w��z� G��ܵxy5�݈��#�S?9�K�"~�d��ӁҪ�wU�B�d��Ł]��?�O*�������>?���+� �O��I$$�E��YNv�iԞ�S������$Xn\�iD���_I8�$2�����$L���p�6�C����/n:����g���S�M4�2��[5�)��=�ing]�,ˋ�wY��q|0�|�q�ٔUb��YU�\`���������俘��^�M�F��
ی�`X %��j'bW;zPK��9W ����kȍ�5*2<d��J.g�����-�����,��������_��fD���1�Y�z�D@p�=�yY�ZN�F�����ʫ���,_֣���D\ �f��a���T�C�d��w��&��TK]�_�*w]�ԫ�;|JX�����9I-`�a��~�P�yR�!��aDS��t],O�6*֣[���/�����S���{MH�ur�=�B<���H�-ʐ�^��ۈ,�W��o����N?TD�6)A/:������,f�@@r"l�Φ���	�,j�Q��Bʪ��n|�r�)��c��g���Hx(>]	�	�*,������i�=*
|6�������vA/O6�����ı M��r{ =��ڭs���Df����	�����|�hP�ȵ��w�~0杍SI�+4�S�ٟ�r�FhH/���*A�$�b(p��򓮴G�o��}�@p�Z�P��{1�Z�U4�����lp���0}�u���^_�)<ӑ2�r��٨/��X*'�R�Ё����+�  �ks$㭛^<!����h��L[+8Z��/0�ҥ�ݱ>H�a>|d��t��k��,���<i�KS@�
)���'���RL *�������K?�C�Ga��� &� K5��g~wzP��,.ܔ د?�v �z�K �X�Y{��Iܮ�9g���=�:j��ظ�t|އIgS�"H��}��N�jO$���H���&|�H�h�p��O��|�J���z�([V[��U/^�b�{r�]!jw�[C}pѠ"�h	ZQxƶ֣�9]R���3�,]��%�`���	.��8"Z��(pd|!��k�?�zu��Jl��{���B?�x{=��V���$�S��̶7�?R���n~*��L����~\�g]m�L�57C'�˃\��Ss��f�(��v�=Zr�4��'����,"��<�%�;�UI��3A��o�d@R�5N��<��L�Қ��Kf��'+LLux�k�=��zʿ/�V��wC�0�N��G�q0��:�Wo�`�K*��d������=��nL����d�#�������[����� ���n�n��q�J�R���0��j]�&��Z��%�$W_�hSs�%�<��SJ	a�q�����:��r�B$>�j�RX���`�Ne�>���U�XJm���ױm� �Di������ғ�~L���oc�)?��!�}����J��)����N���5�� )O\��O��@�š�+>_�Ra`ݓ�2�����$G�9(�\d���/a�p����vQ^�.y{$@�7�c#��O�#��n�jO&�����烝���ZՙP#(�g)B�����׻~�	�oX���FD���H��+�â4z#Dxqn�:��}����4J.���N� �W��&ۼ�3<F�hE��0��H؆!uȐ_��G`�D� �B�T���Z�����V���V`7Tt,�nJ�8R�|3Ay�v�ǜ�֬r�vKgEp���Q[HBl���V}#�|dh���S���rߌҮ�u`G�a\�,@g���Ge�W�Nxw~�~0EЇ�*�cf�@��fS���+�1m�.�U F�����ނO,�}���5��&3ؤ�Rs��u�C����X�G�bv�
��9������,k�һ0�6*�k܀��Pg:D��׬�cDC>B��X�2�O�+�Ӿ̀���t����b�V�?�<\���K���*���Q�����-��E?�_I�Ӂ�2bn��5��֤��,��,��
�1���On����*/�f�Y��4�Ē��OX�M�@��IQR��i_�,�ѝLE��|���1����e���B��eT����*s�,�T�G��O���~y�[Svn�&��E��`��@���|{:}~g5U8�&@�ח,��cM�ʋ����wOWP I�Y3U7
���l���U�-��#����W��,+��%{M��%0-�w�`�����I
�ńڎ�v�
�?
G���}\�F��c��ߐ����7J�*�X�vj��e�-�ң񘓔��#�v��	�6k�3�p؄�|N�%�|ez�$�@������`J�:���bUǒ/�N�j*�D1�;��@S��r�'�7<���P,Œ؈w�e��Ƨ'�%�oPa����OD�Ove�,Y��l�b�O�	Ɠ��>�����p��ME<�h��m�ED���M�~Ǘ�Sr`P0ŒU��`.�݇=��6��m�C��@�e
�')\ލ4��Ĭ�e�7�H3�2ыy�5�G[� w��V����?G�ʄ��e�������E�����r�d���h�PY���a�VD�{�.�{tt�˹��D�EϱA����y��T $������M0�2 3G��p��hvJ��ݢ*�H��3�L��ۖ�Sѽ���m���u��~�%l`��C�Eв�idW�XpA�ZOl�0X�w��磋�����D�@�~�2����슝�-�L�_�[���$Ok�@����.��Ob����K�9���խ,��r269�4mM�99��4�Ɔ�"��<O���cf�rMQ����f�9h˄�Aʁ��M/���&-]��^���cK����~T�� e�@7R$��0rS&gý6Y(*?�:���#s��T���M/��H\�kR�_�X>��#�^�L��w�θ A�KT���(2��V�d��j!a�캳ϫ�P�beu�CS�l%�EI����ZC\b�q�K%��)&>��-��m��ܬAN7x��j�"�N��G���9��J���f��)�]��)��=Q�Oj����5�Ӛ�~�5�ͅ�?�W�h�:}��Xh\{�68ǙG�x2��+���-��ª���i?5OԮ�A�f��P⾭0�p$�=v��t7�8;!A�^������a,�/p�Ϡ�%ɂ�Z�b�;�:��*���W�NN;��4dM+�Gyr�}��]�P����pߕ3���tM�ܱln�ց6M\�)�|�Bl�H7JCoT��C�z/��и{}|٩����1,�hθ������"IC����j��wp�7Y�yM�e��f�v�<��z�*{59�;�Ҍ��$�I ��Q檘tR�9��s���a��8��P:���|i�y/m�"ލ]Q΅.�� �O�S;Q ��RҸ��c�c���Bt�֐���㰵z[�5��٪�7Y#�m���� _�b�Z�#�!`7�r�7!��������i~,��y���n��DRD�V��o���OPI=�S���`np]�����@�]����f�(C��$=C��L[_���ԩ�VQ�;�1aS��Խnb/�,�/3o��D�N�v�&��kc@X���NFU�E����1(N~VN��L��<�搳��g�UZ�qyP}��@�m7 �Z��ڭ�ۂǑ�@�p�_y_�_'Z�����GB<�����S�~[#�%Xg�ձ�Rq&?Y0�u(MCc��6 F�{���26ݿA���G8������GF0T�g�Z!<c�`N�{����Z�"�DE��;k�F:ao��]Q�<��_�6�x�U��\�����Y��6�|	"�"jӯ췝!����W����\��A��su\�}���1S���Th�^l���TS��~�/����K\	1�j���.8]k���X���u�u}�͈�ߙMS��B�ۨtG��E�#�X�c�O�����K�m���ހ5)�l�T7� ̺m�m!{,}��U�çSe٤�@�~)���Gލ�:��,�XWd�]��m� &�E"aҬ�����K<"�>����L\OJaT�V6fk�������]Y�"�v�� R�"����.R���D�b=��)К�[�g��.g9���'��fz�T�; ͫ�V6M��!&����F��י��{��h�<�Q�#�M`�MMY$2�N�7�Ĳʪq@�ӯ�?n�?�Vj��~w�D�Yl�:�'����2��x�dZ7i�n�6#�4Bq��7	r�k�f�EOf]��y@S���96~�}����(>eΚT!"&N���{�M�������������]O_� �i��rۚٱ�K����еvC!zQ�'�%�ڢ����!Z4�e�Ss�ѯ^h�/`�G��cؤ��B�l���3�5�����2�QE�u�����T��a�WU������#V�
�'m�hc�8R��.��|V�R0�DҾ�WоoO�I��}�����]Ы#���+�?qC �ߑ�h�=�f�Nl���������\j�gZ�RimA��{ ^�~30�����0f'Z�Q��3��ʹ}3r r�g!��dm"�����u���5&��\�A�av�ޕ�]�~	א���\���G�^�4�a�F��2�� �W��` ��ud��ŷ�qFΨY3�$���[@n�)v��Vi�Ce��e��%$����p�e�dvR!�0}�+�|Gm,A$}4]��c] �[^zRv��Yme���8�+��^W�O:�I&�M]�!���kX���MMs��b�����s�kَ�/=��(��M�*[��7I!M��j�u3�q�U65(ق�G��7	��!�[��8k��>q^Bv����=�6���e�'�HG16�aVX�ӳ�yq}^����p��q��N&Y�qh���d�(�ՁT��-��]1u�����Y��4�PqK�����smm o}L����֎i��DN�n8��:� ρ1���a�lԿN�f�홷���c��T)r���(�^b����Cv2ᬞ�^ԙ5�w,����Z��ʞ�# K^;qG�uJ�ջ��دq�/��ܮy?ɱI.�U:)P�ȹ��3lC�߉�J�񮱄!���ӻn�
���}`iĠ��(I}o��!�kA��e�9$����|�̓l�V"1�QCOW �n�E���䚄$Ț��d#���jCU�ix%�nO����#�գ��"�gI��SYB|�4B��CɽLiթ7�'���D�E�[��(Ve��^J���A8�,=��)���"~��[�c||I�y��hzkF�S%���#^`
\�]��0�4W*@�z�f�Pij:b%�#V5K~o�⿝z�m�7�~d���Gc]�CBl��-���0�fv+���F���aU`���e@k.}�*ƙ���+e����_�#�ˈ3X��ă�j�u������X��H���<d"�:t_���j��#e�8��C��i���,��_�mtט��5c��QPm��?����[�0�(�t�(-Eu�F!����S��ow�C�*!��[=���4�ܣg'��S�̭�'l����,kW?���p�����$.zv'����u�7'�fGB��ӕ���ez� ��K
�r�Q>b.%�B�����S
���?� �f�˩U�PM 	o��+�N�����"�6�W@�fkBCM�iӛ������4��}-7�Npu4 𢍮���{�U%}��i���-�6N�����vo�s5��䌺0%�X�cMө6fh:�_���-A芰�ȀV=���}�LI+Bi��w��T&�˶�FJ�؄)o�!�������V#���KP�>_��%F��.R.��a@J�Mȶ��ѼG��wG��i����?�ϋ���(�@��I,׎l]����������c��P%��v]��Y���]��(����U0�z��]�����4ƻ7U������a�^��R����Otk�t�)�a�V�L�Q*��M:s̭�~�wO�{�s�սeJΫ��W:&l���_-�:�V��Ꜥ�:�Pf��}�T��֑LlyȈk��6ug!}	ԥ�8+��Q-��������
-���۸V .)�h���aV�W��qU���ZgӜ�/�������s��;�5� ���z(i���H~;T��]B&��#�©��ϱ�&~�,��� #���2��
�˖h�!�f���}�z��@����"Q�s��/\y]� X�^��w)�f
��s�V@�i�6u�i�7Fmq5<v<W��|��$q�rz���q~�����S4�A6c���1E��~�՞��Ј�ؘ[���RQ��Y����}hMK�� ����P ŶWl�J;B%P�ߦ*.Z$::U�pl�R��)�%�Cȁk��gR�ʄjBfiP.ϑI{��90z����Ā��#�_�#aX7��:q��i�
��j��bD5.$�`CʪӾXe'<_�EAu)���g�l?%bTD�U�K��*)�;;�έ5�Tg�q֪pGB g��dq�њQD��@'%�C��ۓJY�/D��,����u%s��$]\m���R��9F��u-R�͔Z�#}��(LYJ��9�i,C�$L�CP�P&[����ع������I0���D:Wdi�d<6�Pj���?DBɗaE�@��������0r}L����7Ũ
)�f`W-2 K�H��Z��AJ�-���l�񊺘ze��J��'��U��M�ǟ��B���8ώ�?[*r�3��fs�Vwg-��"T��M�8�����;���+�ٗ�}|��${-d�9N_Y�K�0��x�.���5�W>,/>�|��|_-2�G\��xߣ_�{�e/^���;�M��N��Iծ=n�J� �YZha��vR��2�ȅ4������\���"P�q���Ng����]��Iv�98�����u��T�^�4ﮘDbuRJ5X�@v�aq$��Vq$�?�ޙn��4�*��OB8�ô�ԛK`\x"����!���� �š��X�Ɏ*9�VN\@��9o8�����)�� �q��V���� ��p�C3a�j��#[/�K&��ݢQѰ���Xu�"
~B�E�p���h�s܃�ׂT�_��(��C�M�� 3Yj�pD���ǁ�+M6O���ߐ���%��J��~�����	�2��� (׊�*�]=mY@j;A�:��$�%�D���^V2�3;j�l�7d�O�a,��3�8䅱E���������w��ٶ��i��}&������/��Q]@��
�_����R�F�$O�Iw�pu���S���ya�a�a>\�ts�B"������`Cܹ����׫�m
�V#�H����WW�B��[�u����!I����4�S&�#���+�7mwy ����AX��E%f7Ɯ�ABU��2kl�}�f+�wZ�����`��'��z|@��)d�㋔M >o�C�-�	�ؕ���	��0�����������_"AI�A�z�Òc�0�����5�7���-�9�y�˱��.� ^�����֔�2DBZ�e�SZ����>�N�h��3Hl+~����=oo#x�0�QV�xA�jFJ�TtY��W���n���o�yFH]�������{__T��
89��}t��/5H=шD��$�T��cW�T�٢�n6�'�t�g�VaQRh��6s���8�Wf�4��@@߿v�M�3v-ʳC�	Ǟ���8���d��:�㔁g��b�}*}�Ɇk���Zq1�]��P	�H_�E|T�+X��׫9�� �X�c��ة��s����R[̂ܝdH
~�P�h����E,A�����l�tV��A�!oS�k+-��v�����Р69��}��ZՔ&"�/���?��(0@���\��N��:�)���C��B�(Ec�qgz��Ѕ*3d����@3���3���'�<�1+F�W��MX"��	~R������?ɗ�M�b�^�!65�A+;��?N����bx�fQM�7�w��*����o�U�f^.'>�}e�Z~�nk��[�mFpF�<�eex��ބ�k���E鼕E?�5KP�!Bx*"c���6�nn�������L�J�I
iM�/g�j3S��j�"�����a~q��P��IbшV2�3SӃ����s�$�j2�tcj�������^��2U���JO]�t��Nݯ��6�mN��:e����
��
I�W���5�����.� ӁŻZߊ�+&�Tf	��������~�)GΖҲU+�>�������(�h���O��N�8]S���l��zZ.�8s|n��⸣��fT�r:�2C��J��cH�/w���w(�� G�1�cZ�;h��w����g7M�$�������j�x�H 'h'�T�3g�9��z5�����P���v��D��%|'���K��-�Q���Qræ-�g(}i�����E̤�[ ��w6�ΦºL$��KWƵM��VQ�ce7܎�����q<��L}���o1$#��������Ky�bZI-���H�d�	�89B�n�¨�Q�>x�^���֢*�����I:��hz�͉w�Q�_Ah��e��qG�7�f�;M#�v��� �>Ȕ�T��A7e��`I���τn�j�Pe ��>��/Ǉ!+O.�\О� ǻ̴ok��'��ˉ�P5���-�p�@lk�����vV�1�b�&f5&��l�yI�)g_�6vʗ�@6t���%�mS�9��G�K3J
~2������^�.v�R@+��se�O�a>�U�U�>�t��Rs����!�!q��F�LRf��EԭX@Hv:SBX؟��������9���+N1u�!��X�_�\
�?A~�a��
4�D �=�ᤋ'�)�������<��rNIzp����EgB̮�GQ2�0 pɩ�.�߃�*�@�I��|�@V���=���
��t�}Ӱ�M���I��YFЏ������,0���ܲi���_�T���fA���@	���Yh:_c�YD4��z݉rJ�Ζg[����*=��g��F3Pِ�-�R���� ,O�,|>,|��5�I�儢�P���>	�'�Ќ�Ng6�K֡�'���3`�Y暁��*Uc��E�PՔ�~������R�֌��o(�3޺�Jo�������@윤�K�H?���XW_��&\�`��+:��.����8���Q��/��ѢG�eb��ꬭ�ؼ:Y���B+~O�.�ì3�$��y���j�Q�{�6�4�c�V�bS0FB^�3�AR�x�A-�Z�|A��w��^k����Y;u:�N;�?�k�7O]�C:�b"謦\��`��
�{鎊B�{�0�-DJTK�}����>�~�Q}g�df9�fzG�:��(�Q�۹H굺������qR��nR[��Dٸ��ʝ�j3��[��=�hvh���3mT��Qj82�O�A�J�3rf���=e��l��N��'��Y$�>�����Hl��ݾr�s�'ά�V6��r����;��u��Q�I>rY�B��Y-�IT�{v2*P�j!׷wMP�|I�<���霂�aQ�q��ΕH�P���A�.��h���r�Gn�5q>�:mY�b2����N�{�{5�R��G�N���7ۗ��hQ|������x�5L��?�ex�R����E"/����ܸw��ge:�zHI�!:` FH��}��f�c���V�f��Lȓ�����Z_F�|�'`ا��L����s�F�����lݢ�X�0�uP��)e���Hr��4��鵬�����qֲh �%o��ģӊ�K��g*V7����ȵiTL;�G�G���Q/׫Ֆ��j��\�;z�-�G�'u�X��b�wϫN�ƥ�R����8�K#x��P��6g��w�+	��'��B��� �5�T%�spܡCM�������YF�j���ϙ.<�U+H��<��p�è���� ��9>�0�31X�-W�@��	�ú@�j�L�9�j�S`DtU���,F�}u�}�,�{|N"Ŕ�4(�=i]�/ף/y�z���z�>[�}�*Z�
 ��Es����0��hA�DW2�j�ml��9�F�$��[j�f�aq#b�*�b^eD'6�/w���s���*�� � g�����#s����;��~G��Q׸��-��	��c��'�>$k�ђ3�I�S��9��x��t�)R�[��'�G�z�>�P�S�g�U���O�Pl>���2��+��Hv��;�S��N/�JI�Vw]{��q���A2�u�C��;#@V�n��Y8��t�D���-ۗ%�P�J�|�5=ζ�@°Y�S3$o�	�f���T+�j:��l�^#��1H4��>�=�D��0Ryi ��c8��ӿ<���0������� �|\��І�x�cP�̷T�!�
x�t�)0�h��q2=��K�F{t;�̦���d��%��\�����ܹj�|äZ��jM���X�W\iu�^��"�	��2e~C8>.�)4�\.�{���TQ%9���J
4�r��/5'������V�7���(^��D�X~>���B�n�^LT�8H��Q�y�$����A���Ж��^c~+�DM�e�;�?6H��Y��;ʖ�ȓb�������4�bM�L�֏w@U}���J��pߠsm����r�c���wf.��D�����T6F5�u`��k؟�T�H����/����M5��s�,�G$��@Ί�}d��Pd�L��i$��{Y��1��P�����u8브��F�W�t�@{!B#͹�F��X��~�U<g�PS�&RR��o���/��'vI|<x���w���Ԇ6�C�{��2�#T���]���D����x��Y�R���YFwE<��]��X�@�pt��:���DG����s5���m�"�������_�^�I���R�.��������p�:��=.t�iU3;I��iV�<��t�K(G%�x�{�k51҉7�"���/�i�4�J����a`�i�#lT����;dEnY1���N)�<©J$\֧,�Z�vo��	`�7w���^�e *ĝ���G!�a� <=�M�ש'�G� �ǎr��r�9J�Nχ&���Qk�:�69��?}�� /先D������W���|?�;z�b˚�3z_�O�m&ׇ��4w$E=�La ��Dd��2ov���%�������Tw�Α�e-��Z3�r��=
6iW�3;���kƟNBH�L��v�)�Ep�}��R4����m8&�v��L���&e������ib��f6>���8[��.��p��g�n���A~�0�6�lQ{^t:��b淵��-$n�I��)[:8��mg"��9�Ie�����a*0#o��9b�2�����ٝ��i:�-�Z�q��<n�i��FX����T�����2���"�Lz!z;p��8��u��4ёZ)!�W�ι8����때��S�zU��Z�x3/6��*��B�u:�3��P�_�v7:s����7E�#TXD1[��I�lL�2U���糯0~޲�$�P���69������.W9ݙg�	�0~� 3�������a�f�魶أW�{E�l�x�k��ڡ�e�f��Ø��})��Z�J��N��{��S՜�z�A9C�wRY����RR[t���J�x;o��i��5�)4�M�KF�i	�d�Q��Wq��k�(jī��u[����}��|7ݣv�P3�:Y���pq�?���F ��"���&2�C��x%��uG��oS�2���к�?��'�-[����j��%]z� ������k��YΜR�dL]Ҙ��48�� ��8Xc�t���z'V͵6�衜
��@�8@���{i(5XCdp�Y;��D�
���x����3
��I���ޝ���)�
GBs�L�����H/|�V���+�pu�.�5���\��݂� �~s?��L�n�Is]Te<`�^�'%Ze��$�?eE�3��>&mm0i2j-�4JTt�M���6���RK1�K8��|�׎HR�T� ��&*��EدW����'�^h�#�x�<��,�����*Izz֎T�&;(���&r��z&��7�W=`�|��59b�O�������Q�~�n����ާS����6.�]��+*@�cċ�>�~ٶg�n����YS�ݒb|��Tu��o�R�� �D�ؠ�����z�ͺ���K;4^���W�E;�=�i.E>�H�'���M�\��j}��a�{-)�j��/V6juʒ �I�oa��R�pIHB�$S$�v��Bwq�X��,�"M�qJ\O��_�Ցc,8���R�"a��b��T��^?[�4��kF�`���u�?���s4��N"�ۀH��?p�G�/�0)�ypzY�`@���\�@�Y�?�p�*|8������������b8(��C��d8���t��Ṓ20c� aG�{1u|��X�ugQC�^���?n��� �i�2i�\]����ܰ�U���Bp���$0ȾkE�?��'��J��C���Nu�E-Y��c�u��\�b������iraY�ZI�����U�3����j�q�
�����!�6���D)����~SgR�&����4��Z�)�h�	�l4!��ȭ���^��ب%�z�ה�¶uŮN{,F���֖�$��!���
'�JMƻy�/���׎)v���}p��Ɗp��l��zG?^�G�K��+9�7�DkΈ;�������C���5F�����w��[T�X�����$�G��S��|�	sF�^�{Te��+�u"j�o�_\�4ǔ3&�ej���Y<�I��#��XN'��;ɍ�ĕ��IR����Xk�O]"�ٔVһM/�p����T�ˎ�kb��9�R\6�w�X��J�݇�eY_*���?�$�;�k�����a�<iբu&j��{)�w�z�os�h=��4��mK�AI)�>�2ءPЎ7qbKe6?����23z^��C�:N�z�f�]��P�(v�w0��:J�YJ����ɿ�PP�^J=�ߴ���z�^+1S��
���z1-�d03uT����M�@L=�[��{��}����7�0[�ĩ�F�I�� ��.��/�;j����kT���&�T�ه+�Ѥ._�����HM��O�[���p �	�}6�#2�&kD�e����������&(lK���[�,
8=��swr�oٙ0V��)��4�r(Zk�ßc��a���.G�r8������(�,fG�Z"�K��131b��7��ohk���' �B�g͉�`��� �6�\gx�/�(ݣȝ��(��vS/R�?W��qz(,O	�
H�|�¬^3i ���N(�,��P.I�0�4ÆR5�>��N9���1��ŃPh�ev���-��d�b|�?B��	�y6�DsŐ�{w�2�c��У��xCi���}F�[3�Ϻ��������?%��������9�N�D6"�<[]��+6�Q�Qh���'����A�	�)�%Y�y$Xg�z��]���i	o�O�����Ap5�r��]ތ4~O�xF9$  #} ��L�9�w���ZV�6X^��9T)ӱ��MJ��a��]DO&�%�|䍨��dnn�vs�XP�.w�"� ۊ��fj�*#2O����6+F$�����H<c��"0�����D�зhp\�v�`��c2��@|h�>~r$��~
\������gS�&ԃ{�b����p@ԉ |oMc۵�pOaiW3�!G�C�N_�c̴�S?=�$�\�aMP�ID��
��E:8Oi�o,��a�pi��7�k���$hi%+���V���[oP�f}���:z��f)z�,IEs�U�����q~�=�n&4�L���Ҽ*�'4$S��Q�v�)n=�H�;��6�|?�?��&�4^6�=����^�l�4��������{���-�E1��ӿPB������'�����y���UT�`���$Sd�.q��G�4�d�m<K�g��Z��9^p'�A-:�A��M�� ��Lgh+�-q�Q��N,q�s9�NP����7�,6,������L�nغ�붔Y7�6w�2�Q���%�Ȧ��O��8DD֊���ͮ�D�}�"�"�
wF�4|[��+)���xBt��;�9aoE�Fk>�d�Q�uO�X���T��S���b�+R�-U��*�iO�`�5��-�lQ`Ñ: &�u LG'��;�w��f�V�l%���j
l%��� �Xo��͒i�D�ܒ&�Ҷ�rW��a�O�]c���W���J���/Թ]n
��9��dcx��;�(�q�������"J�K����πEο"��{JG[�����T�}Srd�uM �1�o���g#J7���~=�Uo��`��Ixۂ����%]I�D�IQ8�u��;8���;���"$�ʹ�ǳ�z�����'/�
B��,�F�)kW]`�����'��]t�?.0���%+5���&��"�@���ؾ�@aT�K���n����_�у؛&y:��[~��/�%��Vغ9�~�B n�~F��D |���D��&����Knt��#��I���ڬݟA��O�O�⃤۴��U�X~�h��۷���݂�^%w��FBK�)TO�퐔'��l?�PX-�]�/{r�%��_r�N��>}�Ԟ�<��q�6�k����	&��`͈���0��$�Z[��+������È�뾓^X;��J=���7�q��ҍx��O�FڷH�Pq��!�:B����1^!AQe��ɎG�Y$�F|K;��U�A�9B>�@��v
����s�s�E�g�εw���or�N�or�0q�=[4r!p��0����\�U ���$�f8����ے��2|S*p�����U���N��ߨ�R�C$����,T
�a�W.8,����]//�t��eM��*Θ7u��-v���ނ��Q>���>����)�9�OG���ғ��|y ��K�(�Hmp� ��[�M���%FM�MC��[�[�"=�yq~W#���d��cCA/-��o��W���]���n�9_c=�{�I�ѷ<�{V��x����� ]��3�J�S&w�옝���wV����V�c[Q4�~��$� �i	KʺN���({�?X��������|�3,ֹx_Q�v���y���r�&F�kù���d�kΕtx��$�֒B ��K���3U��>�B�"��(���� i��U��-A3끞���PB����ù�UӔ��զ�U���s���Wa��Kx�3�T(��C{�)�ݿ�>e�������K�Hs~,� �7U����MU�RԨ:{�Jv�=�r��X�5
�f؄x�����(��z���q�{cu��᝼z�+��}{l��qS��_�:'�l�E�j�8<�X�S���H�Ou�MK�Q�6w�;��G�����a}U��֙��K���t��)O�y�ɱq���zć�6r�\��/�%��cE���o;�<�醹Sx=
��� �j"���y;^%�=].�v&���ԾP�_�A��^�(ܡ���DzX
����2����*�T]$���C�����
�
���"��Ƃ��e����N_44ѕ���\����Nq��-�%9n����,4>�W=���
�TE&4�}��M�9K��1�*�XI��v#��-N#�T0��ؚ,j.sFdh?7*�B�0�W��O��I�$Q��Y��4kpV��'��|��'���m������7�Q!�p����1;�,PL�M|��h��]���K�O���@BHS�vk9��f�A[;��Pq��&�
ީ_�G󲨸X
v���ט\������`_R�Ir`�O��#FtEñ���)�?���E^����K���)I.�+�\���oq�w)en���&z�n{��b�DǓz8�B㳰: '�:ʷ��K�O9�&�&8Y�g�"d��u��^FFe�Ѹ�iP#n��e�!�A̬n�>D����I)KN��R�V�8Ǥ��8��f���������p^�qE����b�L���I	Kb�*���6N��T��inI$�t9�b"_/]�\vRߌ�)��-�+0� \����z�8���4�c��f5�Y�̪��M�S�/,9�w/oWO��aC�,nǃP�C�q���dG�3Z0�މc|�k�eB�_��>U;XIH������6�Rv$����C�nO.$�iAœ�٢�y�Hå�'X|�i���1�B��h ��)Z� '3�%�(+#<h�����f�+U�i�����^�'�٦\g����r��d��d�nr��9e��'f�;c��yh��T?4q�i�O��C{��
(�����D�4��U)4�Z6��`I;G����'pRuVz�k ���v˸�{0�[�6����}��S�$�z�z����<gAC)��|fv�w�2�4�pV�j��c����s]����$�e	�X��1�׼;]4D�U�wg�m9�P�Q�o}^#@]��@�h��N�����
���ڸ�BbV̂|
����P],�
R2��Լ�*���T v�����ōP��G�����Z���stI���:��-�j���
4N�$Q%P��>�ÿ5�s%a�Մ��)L�:��.N�-Y��͐�3�A5����I��f
0�o���%e��_֤�ݟtJ=ږ	1]r#
��g�0M<�R����U�O��K�5A���6O� ..�L�0kL���@�NB�ᑨӫ��fiL�e�� ؉v�E.;p6/-��Nt67\��$�s�K%J�Q�%�+%+������*��t�^�+���zt3'i��z�U��k6h%�"�G�$��v���E���D֗ƨe7��_p6�B�ȵwk�PX����$]��";�!�#�k/J��~:��p)�r���x�ݧ,}��9&�nH��ۡ�* '��u
,JX�7X�z��S���#�d�a �/@�rU�N�����%8�c�m�Uu�Y0 /_�����䰸%^G�J�����$Bi�������OC�����|�:�b�L�N0����8(�	�C����#i��c阗0s�=y2�@��L��U����Je��1v?_�I4i�t#���c_EBp�C��V�i����"�;�@��?��o:�̸u���Yd�Eo��D� +R��b6�.�#0.�iS�/D�V	�u�@G���ؿ����U����>�s������4N$���ɣ=��!���K�R���٦lV���?�w[����8J���i�3�x�"�!�GH~�umSS榢�Rʩ{a�촗;��� ����B1J�V�����b�������@{��^�bE|Tz�U<�\��uU�0r�3���1�wVN����oKgzD�����'�g۱׍""�r�	����~M.��Ax��ɥ �ݧ�E�ٽ7��U�)�h��cw~�����gv�&AϪ�{�`ӶS�����w1���K��k�;� ��ֳ`���F>ޤC��ӓ -�J��э����E��N�B(g	�Fa+l'䯤�h�c��=~7��\7X��ñ����(l���$
+����6������P;�
[�C�i���Cy�/hǔt�c�=LU\��vBfe��C�}!��
X]���ǈ����������^WR����f���=+�8���g�`��%/��fB?���R�_b�ޞ՞x~ML��g�㭇��K�)I��vq]y�G�E7<q�7�����{�����ǅ�4�����~Lw^V�/z�f��5���*{����;�E���|b���㣱X*}#Q��%����ɴ{-�o��X�VZ��(�V\{z�A�#ff$;��X��c�Q���� _�jn#��e�q�Qm�#(����<�
�3��ɀ�K-A.K�{vY��`�5��=c�y"e�{/*|J�Ԇt��e�Wwr�v3���I��D�!���E���Ӝ�D��wV�t�0��Ʋ������؏����P��xf�|^�s���H׋'�ժ��[��i;T>�.�.T8���p�*[IA��q!��������j>���4#�^���T?_J���Ķ;Kr�����N{����ן+�f��mr�}��hF��q@�) ?��y�����80�I9V�.�(��HD4��Ow�p��b1)�W�c7�
���@�:�7�m�o��G��u�މDl����/ڰY����֧�� ��:���J��#����0�0���h�|.��`�%Y���j��¾A{�K=���FD��h�#ͫfvT��|my`%C,�<�U���r�d+�yi��Qx�M� P�F=`w��$���-��#g�
2 7��\��Q��[��.�}�C:S@�0e�Yy��V�&Ol�o}��:4 �[j�%�]��s�gz[���z���~u�g���h9��{5��5`R��QS�
d��|u�N�88�!�R#�#b�cd2$�gZ��x��v��b��Ocs�xY4����Ӹww�8���Y�o}�I� ��������U�MQ��.DؒK�_�����J��l B_}'�z�z�IxF-�q�(�ǜڅ+���\ѕSް;�C����!����"�"���_dp��K��;�W7�L�W�?�eD�����t�)^�o�<�(�w���@�\�sR
�D�y��O�
{.j궣�/Q~(+<�V����A�_|����&�;S�{�7~��Yx�I��C}=EݟЪ�H �<uEf��F�]`=�mM��0�G���ާ2*Vm�P�Ϻ@f� eT>u�����H�����C���	*�[�<���/�Yl#��"Q!ML1������X�1�
�n'�pq�\ǹ~�V�=�����VO~;��3�J�&�h�NEg׳SR�Ц�x���c��z�
"�k�xi|օk��Tu<4��i�(YxY�t�9���qgv8��u�@�.H��`��_��k|D"9�J{�7C5���1�w�3-�B@�Jۄ���h9�ŮI�H౼�59�1�U�!�t�����O˸ɍh��5�&���<�h�!�{)��`~�s�y�q⃼B[��!ɡjDJg�aeEI ���
�H���'`��b�ߥ�,M�`!��`��X�q;�l*�����.��*��7�ȣ�-q*���i}�P�/�U��I���S�)h	���ڬ�a���9Fb��&§�fe&��^V�L!�tf�}�⻳Ja4�NI�?/�,�k���1x��^ �&M��	k����R�d�u����`���-�����(l��;�U�s�h#�g5=��On���\2J�oO@߰'a���Eٲoȣ�z�$�A���N�bD^h���8?y�ʎ�՜�2/̴�����Z�Y-��v�ɍ����pR�#&�ґ�HH���D���z�����:���$�^+�2W�ԑ�fS�X���n�=����7�ªOٜ�g��D;*�*|r s�h�0��v:���!�a���8kz�����CH�OD_�l��m��G�aHx�&v`�Ġǃ|b�Y�M︖��q���fQ�]���d�EP}�۔�t��Ċ��ﴷ��qu�"���e�y1ԅ�G��6`O�����1��D�o��|B�'�#��l�.�a�^�"�O&×q��T
8cg�)m�_۱h�L#K�[����B5�S\h
�SlU�!6ve���~M7����f���]�F9'NY�Fu] 
�<�5���esXu�\�RXF���K�>�hN�M_W�*$$gI��P]>J�ݑi���7E��Ӄ���-�2�����G�u�-Wz

�<9� n����i�"E�V��L$�#.�@�p�-� D���:�{n-;�ĪCѸXԙ��c_4�V
 x�e��LhdEM7��
��I�7���0�ќ[8�Bt[@����%�U�8� �1���V#v�z���9������~�<p��7
迋ql��hn	#r͵>f����*u6q�G���T��W�Ԕ�97������h5�=�ud|k^ƞ��e���W�{tm钵*��UP�/B�{"�;��vP�,�e$H-��|�ow�a6�F���j����x�<r���#l���,~�L��fPg�s޼G\hHl���\'|T��z���%�t`Y9�"f����2���V�����fHV7�c��@u����Q2�J�R�ʍOR�x�z��s�p�ie=(W�H�<���k�����CΪ{1W��o�ͺq����"F$��.O��`��'����~lQ3x��!4�������z���w�'7�&�؂��J��ٵ�X�hǖ�Թ��O�6���
[]��J�z�lA��6��|sX�,*���.������?<8w�0\��G��������Ͼ�V2�� 㓚Ϳ�AOI�����yG��ˉ���jh��-a�J���*$X��6�X��C��"گٓn�f2T���岊c6��T�4>��H!�@��I u�/�����R�V)]��s���/��ST�L��I#"BF�G�0⫝̸�Ĩ�v�Z�|�qMH=�x��P��ު�L�g�&�����m��9&�S�0��|���~�0�	����Ԯ�ؕ��˃<�g��� >�����W��x��nsa�t�H����Ô�<��.L�X�`���C(�;Bw&�����J|���� e{&�N>���%2/��Ф��K�� ��P�}/d��M6 �˽B�Ԑ:AJ�	g^�g?��4�'�}`�~)��0_U��6tߤ�KkF]����0Y"ü�ӆ�={ax�!-:3���"�Q'V ��0��x�ߩ�7���=��؍uc�K���y��_���0�8r�\"m@�1�H��C��"�*"_g���UK�q�!��캦�),���5�7q^������e�Wf냰��p����NOoP�O ��ղW�{rM���Va�n�M��f	�;a� ᦰ�z���TǕ!���B�:=;�Q�G	����� �|$�����Z�9zǎ��b`�[�,�÷�
V���)�����H�1��NHl��"P�-~��5n����`��e��ͼ��%�U|Pӹ�L^��E�Nn��k	9��>���혲6�*P ӡ<%I�jȱ��N�����<�n�q��K�]�> ��c޽*/8h��`�*c��/�~ԟ0#ƈ���`A��4���4�R]jS����P�y���G+�Gm��G�:��L�6z6��	�1��9�*̤9�	^������s�m�+�&�Ae���?|I��!�δ�Z3�{��)hd��D�n;r�R�bH�S"s+�U��� O�����O��
F�|uo��-�$��_���e�o
�RF�tG�ڗ^�[�]_���O�B��y�����-���Ԧ�#�/m��j]��kDO
O3D9��,��zG�3�R�h������[y��~{1o��w�ѴQ��@�S��틗��4GCT�n$&E����(���g�L�a} 9�s�X��[
+��H��*f�r�4����\T)�����g�oZG�{r��]\N�Q�$N�6b	ٚz@H��蕿\Z!]^���|�Ϻ�}���E{8�/�2	uK��(�G}وh7_oeP`<� p!"�dg�Zg�t��HW�� % N�J�3���UU}8~F�W�*��iʋ�����&:��0g�j�s�<+w����t��S;o���@W��������^c�}3O�䵬�P8|�Ȉ�y{D�-NQ�� �;U�|��K�����`�/P٢���?��f����nW����]��և��_u�o�����V@C;��-��"]��\��;&��V�E������ϛrm�T�?JsK<���c(��s>Z�T�����_�yc�3���E�J�Sh6�:��0P�?�	˼Q����f�?�a���Y8_��^�
�����[�]���P�L�m۶�|�^��߅N��S2N;�Η��^��I!�I�� 6��5��Pp���C��y���j����! ]3]��W����?�iw
�Ni1f+BG��|=�z�X������:-���'kC�k�5�[):3�M�lRi�����5=�Vۢ�w���Z�����
��Ox݊1�{}��oM����K�k�\*9u?r�-�q���u�S���	r�יϝ��^��$'�5z_������O󔁐�*T�ؿ����:�K|�����>w]��;5����_����`�S<�S!��!�;��O�|s�U�w��v
�g�r6U��K'�m� ��mAX1ԁ%������	9�b�����#���G�DFÛo�t�'����/���[�w0������(���b��a�3�~��D`���E���S�=�)��B��z�o��ۈ�"[�yu��������?JPN�y�	���� �`W��[��?/�c�������i���DOE�b�G��w!��3�^P�No���T�2BY���~e�S����6�H�V��-߱�0yėBK�Ҩ�,�cڵ_*���|���u�^&/7l]�)=Y�MtR*��q��	�`�X�^�g8�^�'��ֱ�B�Є���ϼ��Wk����޶3�Z�����K}_�k��XfWq�]�)9)�%ܧB>;y�)X��T��f�1�&��4�)��@-�{�-�"Xxfb.�fMl�E�]�x]�E��H"`@�����M�&�ïC�1�}�ZGY��+�d�E~`�6^�g�b��ݨlCu�眽h�9Q�m�NV%�����;�li�)mFW �GF��e�kI�v��u/�i��	�q����[�\��)		�]`/.0�{�e`�Ƨ�W�t�������*y�f�"���J\b���q�d��^�����bh�;M����0n�E�X�|�o��q���T��[�\�����Ʌ.��v/���{t,��X��� ʢs��t�w,۸�V<f�+/�Z#�R��ڜN���Ț��;(VtQ]9�p��yӒiPF���-��oP�hԯ�vUeV^vS�UFy#���c�*2ǵ.B�sfQ�����?��]�\�����ŞBj}�S�3_Ўk��۶������_��Ʒ�,�@!���Z�W]������}�u;�B(�[C�e	��
�:�K$�w��\ݴ%�)?���OCA,-�/f�7=Z�4�`��0</�x�o�%DJۄQ��wų|/%#�'�2��7��s�.E�X��-�^��x���M`Ho8K��R*(-�����qz�Y�bM\08L���{�%:T��Xg�����p��L��^~�;6��^��Z�����U�2H��=�;���3�&�yV�C��=W�U����tF��/�z+3(ކ��Tԟ_�D\d�2��?xM���)�Ԭ�u�\~0LQ��ٰ���>�t���HoB�-)�eu���%�u,h�����Xq �#ޞ���T'#�� )��/�#���<�ꇊ�]�4�5�"�0���R?V7��Ո[�:�R�aJ� �����
�g��Ty[��	�hG$3�*�*|E��+�nUG ���۬�~���ۚ��;ҽ>��e.Șz�xiY�q�a���͉����E��s 6��c�0�*�?��s�DU���� ����s"�ېʹ%rm{?��p��#�쭹�� �,E+�\bT���Mgk/|\���uY~��aUY��*�[7h�� �cq��/��ܮ�ωv��!Tz��"��_��6������y�� ��E�����)" x�꼍~n~,s��X,DB�m���Wf9���ucSYz���:[���Y@"�!'�=#	�u>~��)�<~)�E����Y)����X&�(�fm�u�
�Պd=�d{G��L��sG�ܮ��`���i}����P#R�4''�V���DN2|>e+B� �#y�K�5!R�tl�'9���>Zb������w!ߙ_t�
�V�8�d+��8�%����l���Gutej�Z�Y�w��a2���q�D��KG[s~��{�dL����| fs��W�iG��;jyX��DO��E�_+l��u�@`��H����+#�JS1M?Y"��J[��.�ͬT�ed��'X���,�S�\>2߻��"��J�X�)������̭��.,�a�peW�r�,3d�r/XD�2�}����3���C��{��Ґ��a���HĠ[L�K_�yVc��c�
��1��E�'*BY�I帢�+�|�m��3z�x�������(�(��<����^����_�6�����{�΢i�ڿ�JBf�����H
LҲ-�y(܂�M}������'���ϙ��.� !6��کx�y ~U}��%�;��L:�ʕ�mR^�%i�v���g�\�c�.]������b�uL�RC��3B�
1݉��.O�b��Gu��7�E����@ ��bM]2�>kUW&�x'�ܛ�'iLy�$�-�׏�e업�q�V�i�\��GRS54��.1���˙� �8�7�͑y"�=��m��)փy!|=�>�2X��|(
Qd��d��y��XiۚH.����׈/�o�T0���弘�<f��)..5$+7�V�v�7)��8^g?ȵgXb~��7a�F�Y�y&	�E��`y3��&XHwd%����GY��V'�����=�.��,�^��HZM.�+Cw7R7�!�	�,� �}08l�(6c�mhqvı�c6� ��$ja�uzg~���h!,��h�hd�r�=�>S�p7�Ev�W	`(-T��z|�_�����jM�BP)ZMeb0��9�9�l�q�5fp`@��%��a_wh?b�C�*L���}1݈������6�7w�n̰���]��Ҥ�ר8�Bf��Ѱ0���E��']埃��\S�?��D�$�ɢQN�#�����p�Z�0U��SPɨN{����_�Y��t��Y��ǲ�)�hN���H�Jg���J��B�� �#����丞++�"�� :9v�XƩL�[d�7��=��|�����,5�<lG��̇��m�g�>�TvK� �{7�w��d�����*X;���.�o �8+��u���9��w�̟?wNR5�:�E�鴾.�;�`�ot��A�2��S��k��Pc:�5���JQX�3�P�~��+�y��y��V���yke�'!U��w������˹~F��H��M�7o1�ub��uW_�/�� ҽl��mb�*��$�'��S1_k�X\/�/9����>]''�ƗnR)FM���IK���UrtKns���w�7�3pH>�O�"��
��	�h�;Q��^�T�3�P"�L'�> �l���3����H��8���S{;P��	]#�=MT�q>zd��K,$�k��5P�ؠ���1��Hkj\�f���j�ǽ>$IU���e_���h�S��Rc慰C'K`H'�����o�A_X
���lM���F\�v��䐧C
ޱpt~Z����F[#�?sҚJm�I�k��\/sΟ�b3j'0��_ ��˜|�r<�ेD��{:7����N6�6}3rR8�Ѧ��qP���H[(.���cJ�|�G�F�d5$`xfG��H�"Q�z����ɀ��\i�Pnw^~���6��	8谸-�X�&Q�qAd]c�
�@c��C����	P���Q��q}U���	!�5�M�#�S`4�9r��~��>K��*tO��q�HF�mfKX�X��,\0уb��~���'�ػ/�D�ٳtD�1�wIhhf����݄�x�w���z�����
S�U3�D'�
���u���3��Jˡ#��@iMPj4��!���F��Ấ�Ud�� x��i@d0���TT���e���Y�ǧm�Ќ���Q��ۨ��k���,]&v*@Vꭴz9���e2	�{h�zA�)j��`?$�P,��� ����*ĳ������������Z,.i�M�eO�&������,Z�4)v��}�
�� ��̢��jM� ,xg�� a8R�"���,�|}�>]��э)K�̨9K�)V�R�4[W7?Rӂ�AaO����7<�1�-r���[Lǌ�Z��2�����R���3��S7z�=f�����g�(�0������<H'JU��\Dܺ��0�EA��;H�����u#L-8ȇ�<�]�t�3!���GM�K��s��{nյ��t�"I{U� �	D��X��<���{�`��CAL�i�ew�$,8O)�=�`�T(�E�_GW�p�a���o��ص�מ�����c���<69�ߩ��j�M�Ғٽ�G���;��������lǡV��[��K�H)��>�g9�/���}ups�F��m~�rn�י��Ԙ��p�d���H���R��$�Pd��,|%��i�����<�i�f/~���	�fs&]�v���?K�w�Nq�u �vk�5���l�M���Ѡ$k���\�kĀU�|R�����=�u��m���,�y$Zoh��AK����O3��w�|��^�,a����|̫���#tA:x����T�$��T��4�Z		lc[#7E�e�\B���aPqmp�u�H�)��OY�^):�6���>U}M����D����E��wp�r��7}��4⭵�bR��u!ʦ�����0�Zm3b5v��1���[Cd����خO���01Ek24�����_
��gx���U�٥�<a��<p
�=x%�o(��v)u{Oy�w�Ⱦ6����j�O���M��f���&V�`������0��e�jE݂ؗ��`�O��ݙ�'y�uu�WqC[W}��t}H���rY���3��P7�>���0x��hra��x;���3�1N����R>-�1Ķ�\�K���W��/����IN�q$*�V�%-U;������a��0\��uo�e�2 P�&�,` d����<kG�����rZZ�c��4���y4,�H��ڋM�,!}�k�&�w�^��H�m뷳�rմ$���]�Uz�|�mW����s�#��F�=�,�3|!t��F����H��b3���,�`?EG��Q^><ګ���C�a�%��7���ל���è�M~������c^:,l��P�d� �YeDH�'=��1��OI���·ꙇ<�y��-�J��Ɖ1�L���Z�K�(*�Y�N�y����M`��XI$?*X9���}뎭�&���t<8�,)"˷4�CcR[WQ����)ש^�I[~����2��d3i�C�<��U���*��To���lIVj�A[2�~ w)���p����fN�㎹G���l'�o�����2�3�@f-@\�����,H��%���?$���T�YG�G	�����e���)�����w�K/SXY��`��a��>ݳ�]�њ���ڽFts��87Tk��_�y���M'�?:qV#�k��;��bD��rF���w7ˀƝƅ��T���a����R$�I�gc׮+�YeE����(m��N�Bo[�;4�sJ�f�,�dk�����P��D-(�SF��\]3ce�����Vt�1����o�����n7�����Oz[�xR���K��eII_��*͉�];j�#�z��<��cc�8;|���	+�G�|���������4�����,��x+��0�p��?@�Ow-Ъ���לMK^*9`VT� �}U�w|�8����bz��Ԩ�^d���K�y�Y�3���\4���$Z�,:}�5���-�.O�+1x���B�����.����z��o�h��e�M����Q��H���K�c�Z�`��,��{��F;�<����t����4��L�nu��Վ�����Ύ' ���ҙn02�_����"
G�A�z,���n+��c�:"�8�s�*��e�Hn�<X�u���*��@3� I?�Ҝ���Ï�cἫ7/j+��q0<κ PXʮH�l$įt^��	r�d�bsPU�Զ��󩐒�8RY��a4�5������R"�n�P��F� �rٌ���ܗp4�A�����k������Z�a���*9�-Kˊ'}�*+�_��C���)Š\� ��E����*W|,O�ҫ*+"�,Yc:�)��S��%U%�*������' ��4��J�f�!��m������=0Պ_U�Ş���;��/�O�ض���y��;i�ޜ����Z8d�j��Mt3	��(�߸-�9�	�PPc2b�i)u&¿��;���?:��_UЙ��K���(���hɐ��(�P�P����:4���v��X�N��I(����e܆�����C%#��4�}�R�����Cb;Q�9��F���l��/�~���]c8�-�9)�h�)S�nBE9�S����S<�*C�����p����}��ȇ6�Vy1�v%���~PL��?��@���O���1R��������Ԁ��"@��ؑ���1`> ���1!�R�F�r/��]�T���noA��-T�
=�yV���~MG{���kF��g� ^�����b�jH�𹷱�2��EIQ��6�h�c��(jEnc$�]P">5OS�moq�^lG�/Ɇ�����j#K��MX^6{�6���t˸������,Wi�r��V�����g]��6S�����ޝ�@i$3��CNĴ��퇂�oR�.�pk�(\Rݒ?WDehƳ//���n����δ^�~����{b!A�����x�Yײh|��7��#�[��_D.�x���`O�wN��q��d�SeM��l��7��2��V�,��7KY�/�N���qtzy����ZD�?D�3&6��[����*D��;g؄ #?c��i|�)<�VTnAC'SN�Z�hT�Cن��m�9�XN"GSAć���#��f���J�]�z������Ӗ3���n�����0��I�Q�<>l�V
�<!3nu;�����cKm�^\#�.�������F��ڽ��V}8{���Uf�#�_oѷ�Ԝ�w0�~�Q:X��x.�������A��G� ��l�G�K�z�I��`�w���0�?(#�H)u�Z�Nd�[`DJ�~ӥ�|��.�ȚX�¦��*�UMy^�zG%L] W���!v�SoS�y�^^ئ�9w���FD?jO�nd��,��$Njf�m��v?�W>4�;E���	�^<)��n����
�+և�G���nr�D����cN�O������
�q!�㼡�ۈׯ}�]t]�����wE'�y���/@�c�jz4�\dBW#�O������\oё`��Bsl	��T�Mw5�`���`<����.��6D��6���~��	a�G�
��������b��@L^l�;��ӻ�?�_j��,�j�7��
�%G��wVO�,h�W�@o��塡��=�����o0�Ӌ�3�<��6æU�]�5}c�I�}ɀgx.������"���,��PH$�D �}l��l&��V;�L���*�O�}+�M��.���M��A���Z�	�a�x�x'&�.���Ma:h �mE�1ic����ʿ�\XR��a����(3�k�Y:�����}�I?Gw�Q&�@+:�o��w%ak�N��A���+��,���`>$�KCY��n����5��OR��.���%2"sBP"�������
L��h��m���p��7��W8y6O�U��%���U�WȻv��9�&���
D��n?C`"�dy��}���}���a�"��R�ޱ0�h<aL~����Y�Fi?Į����2b�H����e7*�ߐ�2� �RHJ5�����w,�:�U�	�:+��Qe�|P��Ƿ�v��a,�E�Ǽ���g.�y>9��V�5t�%��Ӌ;}�v��dsj�&cݺ���g$�/&�	��HpΨ�N]�� ���L�����)�8��Ty3{�[��Tދ��
��>��_N�'=Ze.}���?���+D纯��jd��#1�"�I����6�Dl���o�'x+���HH�c�zp��M_M�1��V��M-��AϵG�D\�4�d�QJ:��A�� _%O�L��Վ��d]�q���7��E	Au����:u ;��7���2��]����'$����b�tL3n :\Dnp���A�%�1Ek�2�J}�" �C�0��,�܍�'�wB�W���Op\o�oN_X�c޾�������������j��"`yB��`�_�]8�L(bl��w Z1#�s���N�������TLL�1�Y�型�%��]������B�x	�ET'��I�M�C�N{���r��Y[0<]�k�\�M���u�4:u0~FD��'�������K#��~#z]ڱq�ooq��\�'��	������L�?t�@�o t#c�D�3~�w�W�c��h������_kz>rb���ؾ��E����S�i"����8�)�B|���R)?n=Ⴔ��9��h= 
���;��Oф�52�e~�ߧ^M�x諾U9{�'у�B��7���$��<��Q���԰��Y�v`����p�ω��w���na� ��
-h�};(lT�����3�'ʑ�h �=фm���N,+�6�:�r�S[�S �߬xݞ_�YZ|�,�.��*�f�M��bs�(J-w唹�R!�����	�^i�dв��qy8Cf���"���
p,V�Q�[��ZH������@(
��E@�[y�V[S{����e�A/a��qZ�d3R}p��T��In�jc��8���}7�%T*�@%.nuV�/��b��	=�`�h=�o�M=�t�c�Mww�����L-�� �(��\-�����Ba�P��� -0�)+��"=P��d'�ҿ���d����pLgq�q����Ot=�����i���y;bs��v���<h��7��3������5Xx���<�����J�@�cPM~��k2� ns�P3��ϵ�I��2	2~�VajC�9���h���D'Mgx�%ȝk��I&������n��G��H6��/en��	�6�w��@�8-�'���b�D�T�v�M���7L��e�䂉h(�/�p�
�����i�r��2�R~��\��sN;vݸ"oZ^�=��_}���e��h��X~u�����t_�t��!˵m����Q�G׆���������YE�G=`�R���� ��|u+o��n��"�$�Ъ�#�>��wBs3�.s�\�F^�Q���cw���lҴ�s2ߴZe�e.�)̸=�-�+q�L�+�T�+H��P��U��@��emv�6�A���x�?��L/�7�H�0��#�ړ�mv?ѳ��Ͼ}�rR̷�Ř�h�Ҷ̣�s+�\����\p���E��1J�g?�8W$����=�X�u�mb��z>�?&���jN�4����Xm�8<�H��@+_K���\�&����!u�z����ft!�/H1�w>~̂���w���.�{�ret8)dǱ9o�˹��D���T&�I?�j!+����r��`�Z�&�>���U����Ą��H�x���xi}�E�=<�N���u���yA���Ay�\�W�p��{�3f������(�ů]\p�)��&ߛu��j\�}���Z�I_N��T��X�,C�7��A�-��ic�}$���_鬕���PL�]g��&$������ z��C�!�e���С�V ��`_\(��;�(�L�cos�g�-a=z�1T-a���e%����c�*��S�(]�Q.�h����Ǧ��ޣ���h��Y柪��[ɿ���nLm(g�����ޅs�T������<g�qu�:��d5� V��|R��5��~�>N^�˨R1#��Y>�a��P*�ŷ��%t��rU���zt�\V�-̵K~�O|V/UI�J�h�� �v>n����vЅ��01i]�X��H�8��s�W�9��<>��t���/���(��q<(��a��%��Kw����$~	kȨ4|#*����9N)-��j��¡D�A9z1%s(�Z|KûR��&�#|Yx�c$b`_�/�ny�
l�,�����l�i[v�7�s�<$�����z�y)��d��%pCx	� ���Œ_I�-��|4"��(t�'Q^�ظ�%E������X�0t�Ӓ����~'�����zud�MK�� �w��J�6=���j�_�	�6W�<�$�jJ������yW(m!
`�FR��nU�럒�#� ��Ѷ��JܑAr��.�n�=��_y�����v�{�e�]����g�Ү]�s5h���Ta���������ae�A>�%!����8�d�E�d�B��w�;�㰫� =6����0��d}��q� ��yK�\ K���}�"ŀ��d�>�G��)��pT����V5�Y��o����Ta�`��`��F	��HQ����3;���&��۽.������۬���٣�uG��I�$�"�ZN��80$�y"�b�L���>20@P���O��%�����H��$�J�zX�v�Tpw�@$<엕@Ĝ?��������w��� ?��r����d�+L֥�4;ދ�	LGF�!f��Ֆ`ཆ|\�+9����2�Q�
C�d	/�-Ն'4ލ�8�����`r��❡�1f�V�]�K�;Z��X�UX��T�t��z�Kω�d��3x�sI�-V����pM��Ϯ��]W�������b\���3pR�BI���Sܕ�]S/�/�0����n����T	?���l�ǚ��w:�N���~���L���� �����D����T�!��15����yM��c���F!v�E
�q@��:O��qgȎ!6�@�����%�)����Z���?sn`1�=�uvU_D�-1�X�a)0h詢U�>q�8�upj�ƣ�MY~�-\�9p0�Q�_�-���)������/g,1sNIX%&�͏� 	}8g��՜�k�W�<��/	�1Ƞ��R6����9��������U �=�d� J���&a�ܙo��9��y#Aɩx����b~�	�*���B�*Z�Lbއ�59��Ѭy�Xy�w��1��T�}����M��N��5��p蹩@�F�O��#�N�O��i�wlG��P֒�1gm�-�Y^���a��\��Y�b���^F�el�]��#Щ����}��Y��{#k#��*������b&��d�+�H�qn��k�csJǺ�;|��Hu7�P�e�7�BF�š|����V�0j.L�+|R��[�V��,�'>�:گ�MZ.��$��ܵ�Z~
J��5���D�A�X�"W�L�Y[z�p���(#��/��X�w��aѬ��|���E%]"���
[9�����ăm��7\o=�����б����Y�E*W�&<�x�Ǿ�~�(����2�T�h�	͉Q���.f_o�!m����c^:ĕ'��V.T�j�f
�w��%���zez�[{:�\IO2Tue����D��#��4�*�qE��F�����4ԙ$8��6���QП����)�1�RdP�օ�IxP�0�HZC��r޺��ި�Ac�E �C��,� ����'��2EE,T��{�DC1w���v�������b�aZug ue鎼QC&v&��6�0��}Z�����Pm��0s��w��Qx�Fh=�|�śx�F�_�����	���2����ܷ�s�����b�@�>�����q3 ����&�/s�=:�"�/x�3&�ˬ�J���n����N�3L��bJc*g���2�7�W>o;���Uh�r,'�` �荛\��NH�3P+
�L��jT
��u�/��Z�/=��4���x,y��������c��W�W��>��ƏwE ҭ	x�s"����tp1!�P2mJCl4Y��;=T�2�P�f��2�,`V>�BB���vV�%#��2[�P]W<N��w��	"���\aţ'x�|'�Sd�`]S�<l=�zk;�����r ���
�1K�c+�S�|����H��pᒩ����d�y�Y��iE*�#ԙ�q�����QR�<~���v��I���S�UE��kX�h����	-�3�T�_����r:���rt�rn�ˀD%}k��C��@���pK4U �y�j��l��k)2_B\M=���.x�1�rQx*aLM�$\�N>�WX�X���H�1�d�g� C���O��g��	�H�FG6X�|�z�p�\�w!�B���]J�z���O�H�'>�c�G[���j;�u���\��Z������D�����{�p�:�&Tm3�P$Oz�q����ۣ��~����Q�~�j�U?�Q%`�l�`���p�ۜ`FUr���J� 
��7_�j&Fʊ��z�('<��8U��|c�,c�i��%���a��0��:����'��È{�>�,�
��S��O�q�Rn��G��b9����q���cZ���*u���I��������L�OW�� �;p(9XsH��1�2_�Ե���ܠ?d�N��!���I|��)�m�Zԙx]�H�4��z-:ٙu�\����A��O*���Yp�0n:j�bg�O]ys�{�̂��"a{\�0�t�t	�д$��DK��І�D=�s���Pã��@�܀F����u_�TB�����(Z+D:�V�E�T��ʍ�+�HI�^��8�䭣�إ��`3�����G	�y��5�;��QZ�%3��_ŷ���h:�^�֝CLޢ��S8  �)xD��F�U�b/�(��'�E����A^>���=!��������5"��(E���h#�ܖnq��x�>O|���@��r�p~���K큜v��5wD��2I�9���v�oK�6w�[�68uF�$���٢Oֈu,��bC�ڼ��|8�>Xq�"�t�-�?1�����T[N�ǆe8������;��e���B
36�@�s�/$<�;��ڙ��p�6���
�ޯn.Ҷq��r�\4�����x�M���a&Ȟ����$��Y�s�F��GٞP�#�H�dދ�Cb�
gs��ɮëϩ�iɆ�f<R@�	� z����R.���s��ൽ�-\nF��X��̴��)���j�kZ`?���t�_/��e9()�,�����;��%U7.���}�;��N�N�Y%����ʍj4������Fk"�P��oNAos�G�XI��0O�~�k]��~��
̛'6k��SqWJ�:Y�7�����'in�u�Q�Y�	Ŀ9����cZ(�~>��<�+f�XQA��!����j�\/��D����"��}���(ŧ��pҼ�qN��:u���}t
��Z
�;�Jz�N�.����q�}�-���N>��� J d���xZ���������x�(��z�Q�O�ҷ4��vAo7h5�Y��Hi������/���Q-�Fo��Q&)����| ��S+�K���8RP:��7�ĕ��_/�G��,r s1�J�v�����g�����F��gl� *l��R��Ӧl��ʫc���AiXm!�%\o�Rs��Yj�G�8o	�g�:!�A��Mg�-�w��Z�_�޵ߖ㑯��[;�k����0�VMi:0�#v5AU�w��0 =���,4�����-�*Kf���'#N���1�قUo��Le�m���y\�P{���k`O�
N���ƙc���M��C�n؝A'�e�V�ҵ"����D��}�P��;W�.F[n��Km��;��&x�T�Q��$������W����f�ϗ�7�Ab���1m���	���%h92���6F[U4��LC�br�O.�z}M7��1�и���'�b�P��̰/�V-��<繙��l@�S�´X����m)\�w'ң����ם/m�HR�nx��T�'9Wғ��q�_��>3�E�C#�z�b�L��Z���p�~�"�%^�εX�!��[ˉH�Z�E�evNF�9�+�o;R<��7�q��DU�">A9��R�c���F+�W)L���6�Z�.TwL`������k?��P-��J�#@H��IL����7!�j��=�k�D�E&���/]d�ڰ/�G+9���=�A���Ae�T?.I<�\�t4M��S����Ż=�s�+��0��s��gY�T\����*ܿ�/hdA%��3�g����	ct�L(�X��X��qO���yP� ���$d�r���F��-5ܸ
e�T�¥y���WT��1`<��/�A�{���9��s� z`���J�D�©�ݥL�ݹ��~���5�!k��;+�DU�X6��[E��Sm�M|B;�H��Ƌ)�(O���P��MZ\CIF�q7�.�3�/bB��.�"�]�mK �=�ӚM��  vl��jd�KP��n���d`2��hO�)F<m&}5E���J��hGT�i��0=G�.3G�;���[fD׼�x���V+P��HQ�l����(5�p��4z�ѧ|i��X5�K��=�x{�.?���?�N��U�î�H������-���e9�#��Ώy/|�W������)���˳Æ�Z(q�xtp�BoN�"�/�p����Kx �Id-L��5�
XUO�!f��'���Ѧ��շz~�Z+���qC��h�?���Đcg��X��?�h��/�"�9�%�T�y���Bg���y��\�8�^8�'}l�p2g��>�b�;FP�������� 7���}⪧�����r�kR�^��L�4��X����W`k�ϩ���� ���ϒ��r\y�e����&ݞ^%
�ȸ7��M7@m��W���_��Y �Y�dK��4\j�!�&��&�m�a�,z!v���DY��k(�"�bZ�h�l�	�o�M 4�ANج��?<��Lm�V`��K=pf�dGx��!u�|��ś7�A���utwC���5���|�y��a��[�?ϭ.�ce���#)ϙah?w{��FI��H���qg���o'����G~�U�S2��8���z��4+�ŵ�� IU�A�ҋ�} `� ��"N�E��(��v��8��b\8���fn�C����(�'��y�{�e�"ND�ߏ�v�����S-� @���τ�f�����r���HR�2���z�T{� ��K��]á����!i��(H��:y�W�ȵ��I�1���+��N�A%�>���M��SlBlCXяO��cϔ�S�d	���!�&�*�'��2�-��+�B�E ���0�	���qz�2{|g�;L��>պ�m2ǕY�&E I�1I�֩�LA.� #;�=+9�,yX�����O�(f;Z�*�f��1�&#�R*�O�IB�-@Yn ��@C�#kua�a�IEk5�XLՍ�LFsnA��g��<HfOlQ����{(�ө[�i���i�uYB4�ku�H��.zsQ�m��-=D�g�xx{vo����
w�ø�}�u�����#&����vPG���u���G�U�Z����I�ߖȸ���ws�]	�3A��ROU�Uao��.�5ż��Ux�"Ĩ�	��Cx�s���ex5����Ig��!OP�����|`���qˉxC�/�ZWlTj��l��V�a�43I ��_Y�9,|�Vՠ�<���ˣ�.B�{lճ>G��f�?b^U鐝j�tVY�	��.��O���E] �N`���N@�7.ݯ�
��\,d�{�60=<���s�@p�o�:��x�pR���b�B�p�r!�I����)��~GU.������{��2�S���M���9Y��ŀޠ�qG�<�? p�<���`�º���2#�cҞFF��lHP�M��߰��Uwހ������r�&*茧E�%Gar*��yó;	U9I��+�kD�罪R�$���ع��m5�[�K���]��!,��=`���W�����E�����S��i&�"OJу�Jܨ��������v�Q�"���va���z*�fq�u5YK�|@3�\�O�8f�:H.P
E�Vnp��q����,A���C��wr��0�2����C����	�Ӯ��r�.����:7�b� �ϟ�����su{��8S�s��ȡ��J�P��L��i���{?kg��.�s����u��[ɏ۫��:��8�[�rp����yR�� ���m�2���=����û2)�~�����f�aV�He6KWIM�n
�<;�1LnT���
�'�e���4F6}�����>BCJ�c�H�D�/~'T��M�b��˥�c'���"�6�chy[��M+R��å�W:�u�zsf�h��|+�A�6��M��qI� -��Vn^
�ƇNь���_|�pn�6.
�o>V���+�WCrIƕ�Yf�E���LmJC#��x0��e�?��i�ޒc����D�y�0S㐀$�W�s�Q�)��Whׯ��Xn������2���=j5��z�#�;ӫ|E�Z8��yM�,���}� U�?R��k�l�O-�q�"$Y�MN)29q*�2}82�([�H��KMmF������=��݂��i-і�u��ӊ�^�䷈���7(�r��Ā2H��W�Ƿ��\�__���~x�gQc4+k�Aʿ����1��q���d�v���v`K�M����L.����2�f#o�Ǔg<��=;Z4���R4U�}u�]r�Hwz��#�ݓ�����YqKOy��}C/FA���9��|W�%r��g��I�F�I@/p�5�5�q!�ª��l<"V�_-�G�jR���.0al��q#�� HJ��p��t?(A5�d����c���={�Rl-��h*0��A�<��^<��s<����5k�= 8<�)�SS�-s"�d�⯟_�#�v�������|پ�����t~������{��Q;�}
�=?�MU�T#�I.�JdP%>ce����e�p%�"�����6��2�7�SH|�]}xb�zV.��ʻ�L<4O���XV �mT��iU6��]CJU���k2�Ax9��"-7[���]>�䎢���ׇ�˴��>���T\7�u�k+�$���	(F���4Pͽ=e�V�J��EB��`�"s����r,����<脧�[�@�rޟ�W��.KfG����,Q�����}��d��=�|�O�Isv퀆�K�߸8|�jF���ճ��z�Q��'W��wRe�5���n}�Y�4	���7�8c:W�x�a>��(�B���R�8r��P`��#��@ɠ_�t�*�����64!�C`�	�Y1�����sL�o�VW}����c�Ԍ!�f=�j3�va"ڼ֛�������m����l?��2U�:z��y�
��6t���m�I�IV6z���PI�[F�"�n[��GNA��T%�1����ǰ?��r�����	�eTm+��?@;Ӌ�e��ti��5
c=�.Y��uM~%}-<��C̹�;0iD����n�T>[�ј"����p�Z�ýb���)�n����g�+������*���gMD(��jDFƿ!�"ۈ���I����٦��}����3%�!cC=��D�`u
��mj�@�{��DH���F��}�nds>�}=g�l����Z_m�^�P+��a��*Z�"$��<�zz���n
�y0�҆�u��F���dw2ob���l��YI���G��8�y:����E�0�@�^���qҭ��(`2)��
�@г�����2jɐ�N�?u����v�'�Ch�w���i'���eI��w�o�x��Ziî�l�/���9���M[��Abz�0�f�P��}>-sC�z�6 �RI���d5V���K#C��.�ߠ�m�5�++�n�ꃉ��g�'1�P�Ţ���c[Pa���UtJ�\?���[��T���O���қK3)���p�,xt*�UD��pQ�����1�=�gY�V��`ZR�Hr)�����#�a������؄�;t�)�C��DC?q��s�H�GE	��J�>��3fד�/I$��(��S�vsu�A���A����(M���z�~?�@VC,I�n����[n�ߨ�"�j�O2R����FJ�k�W����Hf}�'�T��v���t2��Ȃ��N�����T�:��F��1p�� �9Mc*7�+ �S�0A'����aǿ���%��r*�4�u�Q���FW&u�4��/�b
T�;�W�� ��\E����^�-|��y��R��	1;T�7(/�!4��5W�J��V�tu��8Fp�$����k���ҟ�u�Lh���S��%�M�\n�ĝ��C��G��{���ʫ�K���6�X�3�d�Ӱ�I�,Bށ��e�v�(#���			�¦Կ]H��4m�s����������������oj?,�.#6��;���2~��]��q����q���,>oE�N=dm��	��A۽d(�P�T[��-�/Q~wzNE�h���8=[�zI�0�ق��]��X�z��Bl��J�i��[��%/|�@�(w��Y�Ԯ��ď��A�Er|��/}��Ld�������Q���q�}I�G',��q�1>j�U_wo�V�����dB���Ǘ��%T��i��3G���:xlSԯ�N���s�_X+P��f]a����Z��3�2]�-�8g;���S=��H�&��Q;ބx�3��W<�ȑ�(��+6�a��6M���]aF�D�%�v���}�	w�-�xg�V{edrs����h��[2bb-��A7��u��9��Cၘ6"�J#��cr���0Ÿ��n+8`���Nҿ�A�!�Qئ[aN'�z,pV�Z�*�
����оЎ��+}Pz��S��Gd>��f�F�6CYP̽3����ߕ�?o��c�Vuѹ�� F���>H�~�JK�^A2u�7��>�2kMɛ�؏��ҫ ��^J�	�L��Q���8��xOhK���/m h4���.���c�"NgNVmx�WQI}��>�p9۾s����N=h�fO�Ȟ8u������D���\�]'�%@�.�$��N:x�bc�G�@���SY����`�A�_����K�0λD�\�|�x���)&9����v`ܘ�¼Qeӛ��CTJ�&}��M���w31)0FYd��ȧ[�t����''j���)�_��	f�� bR
!{�͠�q�M����14��~��b�:ېŹ!���\�R@���yhk�?}��2z�#hjU��y`����ש֎v��-��p
g��gp=�}���4x�՞���]��Q�����6�b�5��{p_�������2
Cv�Sq�Yo,3�Ҋi{(�K�wn2����X}A:���f*֯h������'gT�B9tuNJɑO�"B�����������=0~D��~�����T��l��B.h��z�+�P@���9�-�����^/phX���}�ۺ
 qˡ�}\ �5�����½l�77�4jveS\s����̞�4X�_�\Vf�[ʦt�ֱZ�ذ5�gS2/���]�R<�`R��<E���9Xv[�/L\�Pp=�ʋ_��*kU�H�	�.�G��M���k&��԰c�u=u�lwTn.��������F��K�˿[��}ط�^��G� DW{�/��|��ƭ��{��?��h!cI@�r�:�K_Iv}�$���rP�D�I�f�!OC����I�R��#�;H�D���@��x`l@R\������3)���!��A����49�T�|ED��f��ڨ�.�:�p��)��s�����A��f��ᔬ��P�et�%�Z1��ǻ��5�U�]�8�D��d��m+0JJ��Oy�h�Jq����􈐖`��3j��W����3Ǘ��^ސ�����"vƒ
"Mƾ���Y҂X����Fş+����D��s?0`�y�&�dG73=Y�5O@�ś�n�'&ݿ5V� �%ɐv;�?t�`����� sR3m[�D�W�)j�q���_�$��h
)':u���#,�����Y��9먮�LpڠQГ�7�`"����ƚ�0�Ŗ�p�`N���.�r�
��rv(��L!bo`�4Ŗ% ��ˮ@�-d��?����K���x�d�U�a]#���m,e�Ӄ�����ǵ�XK�<��h`@u�ېP{�˪�E����[{/*g������6�l,����M������������^���Z�S4��9nq�a���[u�ڞJ(��G�y]|_��ͪ�.4��8���}�����غ�X�˓�[Zۯ7;��܈�J�	9�:�'���~��HHļ�0êO�b0|�slC�^!��\�K���hé�<�$�&#h����{���#��#E|�W7�q�������Z4����g^h!��<���S��|>惸�#�{X���+f���
�Z$�~z���E�Xi\���W�DeW�e%�Na3�!�u٘���D�y ��S��������3�,�~��9J��=f�Y �1�T���J��9WVr�ٓ����WU�@�̥u��q����E�A/�c8���oVL�<��͢N-�>����z!��a��@P u����6��7��5I�ג;�]�+J�� �*���.����_l�p(1>W2��Mf��&oh%��J���j�Y�kv�+�B+�V����z�p$w������^�۩�1Z�aف�c[�qQ:��f^(r�Sd���͍n�\���m0��Ժ?��+�̮"�'Leٕ���:7��oO���O�0��%'�)�h��F9Y�K����&�S�'���<;�uL��yM���H3 ��@���T=�����E�l:�]�I�j���[�p5�Ӂ,�h�0LԨe�KK���� �L�(����zd6�ц��q,f���/�]5`�t�(��τ8�7:���۩N��p�{�1P��:�Ft����g����]��x�>M��:/�ǆV3�Nv���JC��X�u1��
����)�����θqÙ
v�i���0.�l����l�[���2�}���X�-0bhI؁6��Y����8X��:ʮ�p���&Ro%IG�4��
vV]@O�Cu�_���c��PO���O��O���s�^��g h��z˛���뼐@�Dx��\14����T*��B[μH �yl���c�������Q�?ڸKi���r�=r:٭_E��X��ˑ�R.�|���Z �
�����.�w-9?Dc
s`���m+����S3W�y���ب�J����n���Ԋ0�/�<�]ے�ݖ�X��[XP��ou�fn�|�=m� &��ڇGb�l&��s�R��'���X��5k���#��>h}o��amGI�bo��$��D��	�_#�eG��pL�G2����ڵ�PJ.��))��a�(Ȩ��	;aמ�i7k�f�yj�7h�Ⱦ���eu{�e�V��^l(����x@F]��zGWj"����~��	�T ���A��� ���\Ϝ,���9�����~T�{E'��������� 	���Rd�L(���$�@�V�m/|τ��H�����;�nC����]���x��gX�2�zi��mӔ�n��2�%�,�Z��*�V�݀MW�Mez(�Q]u��W������ź*AjJꓢN��s��,#�&����'	��Q�S)��<Q�~��S��k
;V8�l�a`cm��O+���(��et�B�^wig�e4gσ�����)}��Z5�̝g8�����Gu̩5�٩UԾAUe:�!R-9�����+y��R�b���}-h~x�X���-��U^A�>�WI�1�ct/����M�D��w��k@�T����� pZ���G;��ݳ���;@:vӱ�O��9Z�(�@�ٞ�����9���G�%ыi�΢���aV���]��k����eI)���C
9Yn���5�6~ŅU�n!-���nE����a9Q�� AX�#9��3O�����`�M��x�!�(ܻ�l���`��ۤ��M��#���;��,�}H����:!�����L>��ҊJp��t%�ӑ�a��$�RA��v�[���	�t�ő�W�~�S��¥�`ds����\z��ړ�4�����xv��Sm��w���4`����`��[�D{�У
���y��4�}����E\Z�I_�)ó����]���:((���_�m����~��;�'x�Rs,�	S]�G�B��y2?'�D�<���`}��V�C0�5��n��fa�Ϝ�:�Q�E6�J��pb � ��(���p�Y�;�J�X��������++��2	��j���J��T���!�)@L��V��y
��*^�w�R�yȪ8(���ޤuK�X��&��������mO�&�OE��h�S�4�V;�24�Cج�6�U/E73򱚏����A�<�)�F#��#0�A1�j���8�XM����y�g�� �u�M�$_B�vO�'3�B����2spY�sk*�1�r����b��!�w<��Fz����]���x|'\M�zA���8���cY��`��l>��7��.>}}O�X�����/�q��g��3x5r�I��](	b��rĐ��שy��,D�<�����D9�#f�&��k$�⧢��]%-J@π������YIv戮�j���{�������#8���%r� a�OU4}�G�I�i��[��6��r���x�v?\�e�V�?�?F$�0��,_�LX�)�\���[.e�'l�Hݾ{�ͦ��+q����RY��] �\,�%��}�&e`P��F=�B!K<&nb�h�H��@(-'c�_���>��Z$�v����~��wWe�}V\���gC`va��R^B�`�9qV<��q(	3c�+u�g�v�ǋ����-�T���r�2�sN/-�̕Qڨ�Ɉ�?�ʎ��`"'3���zG><�M�'�j8��V�����.K�I�������&�X?4�����6����z�Q�O����c���m8��0af����i^�Ә�4��K�%���1ndt@3����m#�z8����r� ��1��4�������h�`O��;��	���q~�N1K�)޹e��b��k���C=2��"M�H�_*#�m��'ͥ��4�ǘ͘��Ig��_�m}t��8��5�ˍ��S^�И�;o$�|�FmVA&������K���T�j\P�j�=4�&ng�F���qtR5bC5�(w�.X[t?�$|Ȃ�TP}�%���{���g�����Ҝ��,���K:��[��rnr��f��H���#��0�SVs�L����*셻����}[��ݐ��)V�D�h�8T�-�u�̋�b�0Ʊ�k���i�s�C���
�dN��^^=����P01F��C�"߲qP��jx�F�T����hT�mٮ�؛@��OZ��wI��0��*n ���r|s�~�=#鄆
^�jaM�1䍷��g:0m�\۾����Q�<i^F\��B�~z		c>��AZ���L܆^
R�
��VW�'��q(�jY��"[�����ȌD�lb�|��)vM���i�Q?>Œ�
BV�3��rv�Ĭ�kk8Cd����ڶ�ᘔ��<���(y�Σ��&2EC�$�!^�&�u+b�(���G�-3����T@�1V�%t�|�u4
1��W�s��N�����-��ς�8�hm��J�:9�BE�΄�����K��Z@�t`1����}���a;D;��M�0���Vwz�e�<�3+킿�]��jV�th�X��6���)�_���kֽ��
i�A�W�].}d_��_pT�7-�	R�i�8���[�¥$3���ZA)��`�Q�F�춳h`�XQ��U��ۭ��p��;��p"ƈ�.dR9Y^��hIWD�Z�D�lB��4�0Z����+�����M��'%B6v��y�H�|���'�(�mD��C�";V>�C��!����^ƿJ�"�@���,^��,G�R�Y��~���;�չ����5m[��-�7�H8I�*�b''LNn��,K�}�����1�b
iZ�.oɒs�23�(��<Z�����h�C�*�
�\�"cc��`N����L�,�vk�O�,��8��:m͡���v]rh������ubF-�~���_Ɠ.�.j=Qgb�c-��5�G���5'��9>�t2;X�x��&�[�4�RW���C0�>'�2QYT�Q!��G/*��}�3_����'Gd����`�
a,`,����pw	�8-*)�"K��G-��[��9g4`_W6j-Y�~�F��_�������:oo�U�O�S<!�#�6
zWu�e��K�ϱ#ٳ��)q�}ࣳivC��n5��K��������ɖ@���|�n����D��q�_�3[}9�#�5�� (�b�|�5�6�@*%�П����A�!w*�@����,����yW|�H���|�3�u(��q� ����
�OK'�{Ol;��)��9۷I�mL!e�
���R��I}U�a-�1gx�@���N���Cr_�P�m���<��&�*��a�t{F=xHoʇ��P���I�r����x����+��Rz�dQ��_r��Ҏ��sf_&�n�U�9���R)��[U!�:��|�9�T"�t����}��mO`�q
�����ܵv������Z�6K�D���ݚN�}����3���!������(��d"�@��t�\v��i(��᠐hƝ�܋������QYw��؋4�y`��5�_tض�]ɖ��u��)��Sz �ʏ`"?���\㿔I�	�F�~�f[sO�QE	�p)���k�^w`"��=�a�" ѼM>]��D#s 0��� �;G�-edqܒ\�ĺ'!����������/�M�d� ����\w��b%��vh�]X.���4�ф�v���*�rN���i�AqוCs�U���H��7�B�ή�"�K|v����
r��67"���F�x��l��C4�CZn֊�`�]ԛA>=ڰA�
|��>|�bL�!��!��A_����I�1.�}��q(>R�)!��L�E5�A�׮E���k���!\��ו�5�T�I�O,���RǞ�I�R����ߦ�5<N���bx�	��;ZD�p���V��P�ʡ%?�ܰ��жK���ӓhY��u*m;����Y���0���
�Ŕ%)�8�^����U�TC���T�78��z<�$�L"�v����﮳��l���((�`C0�t�NZm�U2��8���w�ꇞ�wh д��XP����w��|����b�l� ����D�yT�����.��g�|���	�Y���ע.y�I�����B㶹�	P:4�P�%�"���IqUچ��(������ǰSD�Ŀ�f����l�u�}��t=�?P�ez���
���1�c���X;��zj%�����=y(곍1����#�4�(zs��g��0���V���*���l�42߹~��\�����p	0���ܵ���_js�g�s�f�}�8E��?���ۏ,V�#�x�k��4�@�~��@�G\
%�ٸ��3BU�f�v͌?�[*\�\\ws��CvER�S�E�,�� �v�Pk��ە�����c�����N��e�n촤&��9EO�% ���c�"��	���������VH��G|�$-��oXyKK��͊�B�;c��(4Kg�ӊ�ȕK%>+t��\���(L��w�� BK �6wba�-[�!�� 󧡣�3%��	��v��z ���M��v_f� r�0]��I�tSgƛ#��h���<���/�ܭ��=<~TL�
�K��������M�?@�I��a��'I����Bwn�5�7{�4�3�IG�|��9a$F������o�X �(}�e��k�}�YAE�u� ��!��P�E{Ȃ�MĒܚ�d�	J��[F�w��!lBIڻ�b��5؀e�I�9V�U�5@CߢY�l;�P�ˮ@DgIU��#|S�(Q�j,Ue�69*q4���щ�(U���B�d�-�M�'��x�)���3n/����!5Y�c,m�����H<�+,�i�����r�����\�L��O��=!�.�6���T�I荔��!Ԫd��'�~�y�؋�M2[�&*T�"q�@���|o��Ȍ��#>YsC��vi�d�%�g��z�-��B%���13�����3����(ڙ��G�m�(Yg�Ol�3BM�%J7�4(h�Z�"i0n�¬�B��3�u@4,<Ϫ��H8�[%�af0�e���_9��L��r����f|ŭ�8j��h��6�>,f��_lŮ����b��!>Ԯ)#��W�A�r)Z͖���P���@�����'��7���F�E��4Ϳj��/��N;�MI)��'��6��˦�(��������k��`�8��I������a;w�v
�����*�@�����]#�c�K����_P�����)���5�u��<���g-!�Q� �����e���Bx�	<��D�u-ُ�����_$,Ӏ�����X�g�&)��K���Eh!Yw̄�6��,+"*�ȑ��E5�2�P�T?�&+ �����Y[f�tA71�B33�"$q�ec���� �����r����X	$�	փ���N?��F����y�;�+�[�e�?}"ƚ�}��Y2a��W�L����U{Ԍ,h���0�^ѿJ��s�{�)�YA�s�g�w� oC|E �SI)��U�鱊32Ƴq���SH���{��lq�-h�)��й�k����;���j�T��b�7�
eY	�j�A����˔Ck�[2Ii���.�A��4�!M#q#�pz�hzL)'�(�R��������ǙC��z1U)������Q�����Sq �k�X
��L�q��\E�K����;'���c����%bI.G����$�**Q7h�ќ�O��t��5���X����>Gf��u�7$̇9j������?`��1`%��JW��O�=έ(<��g�A׃��Ӓ/�s��%������x�ox4�%� ,��F��������.S:�_��=�l[g���[�e@�(�����RPϾ$adӫn���TY.��p=���s&��P��˴liQ'�k?�R�z�*��O��}V�m�7��,�b �����Z���˃�3��P�`Qu����վR�s/_?��j���q�c�%/Y��;�<�q�m�i��1FYy�ղہ
"�޻�i�����6����΋��	F�K��ߞ��1އ�s��Z���yj�]\���Xq˚R���R������pF�����v?����Ҥwfp�Þ~��C�^go*!^{�N��;�{Ն���h�e��k��$ ˒�g��18��q̳����A6��b���������:�V;��<0��jJ��5ϰ]��Ƥ���:���ky�Y)4�|��a�q�<�n3 Ʃ���ߤ1 �,3�6�����{26���%����[�xl~��7+cS������8N�k~ x�5^��!��}E�=���F����j����"5�Μ����:T�56��Dl�0�q&�z"�.�2d���w�N"L��z����R����b����]�ʑd�s{;�J=��;�y��/�W0s��\��{P���K�Γ��$dE6�<��p�MQwA� ������Jl��Tک�XD�G���1?��`Q���Sg�C������/�N�Dd%��c711�ݯ&J�<yζ���5S9V]ɖ׾g�Ό���Pƌ��	PF��y/.b���N�}*�[D�"��+�n/w��(�"���!�W\sQ��3W�?0ܷ���l�-�~�w�6�[�;D���,���z*G��ݷ�\зa�&'�>̆��H�Dú���:!�IC�=iɜu.�����%�,w�f��ד�`z��4h~ Yu�޸��c�E�$���# ŜL��#��a=��T��µ��	�ސe�u���HV�������nN�P�|M�sΧ����3^s��X���g���l�=��(�\U*�t�ӗ'�ގ^/6ޯE�taa&G�0d�Y���62:����η�y�W��	A���^|7�S���Ôj�+�h��g ٞ.Lk��/Mq�`�L-N88�~o�����{ �!O�T�3�� P*�1ZD{��"w�V�{}[؋��,�ǿ���:�2&�2��Ǟ�4b5�"���fLD1��X���B�����H��A8�sTr��dF���"Vqhl+? ��2l��1�@&���?c^{Q�
 t��9�2�v�x�ˌkhR,��ú�HQ�^��Y�],�X�@�'g}>$����x8=����鶷6��`��S%��M���xI:ܻ�����=4i�J�%�[eQ]�6I�à,A��(,wy fc�0�v�T-]�@2_�4���
G�����>�-��E�MH�m�	�Q>�P4�_�������!lGm�'V�[���h�y>��L�&�xo��IJ�k�{�`��2����Rd�޹v*��ʭP5=�>�� �U�5��Y@?�?Ku�B�+wҳv4�ͳU{��	�}"���������C���I��*�:.���W�ԝ�Z�J2��(@M9=U�zꋱ&�����̑���2	�� �����y�������)I�k$�͡Y z���[�X�z�a+�HK�"D�Ԛ�����9��0z6X�K)��&W�̹�(�Z�s��l��C1����`����, �%+k�,9e�����0��uʐ7��цV_�-^�%§���Ib�@3�R�����J����	�����L�J��O��%�+�hϩ}ȅ������<��GL���*�'���(��8�@���BH���}H���T8�aa�){���9C9L���3�o[��G���Z��&��������|(���Ep��5x��e����Lu'��9a%)���EPv�����,��9Rzd���րL���W������=%�e��3�S�;E��`d����F�k�h˄�g7�T*�I�"+���a��nT�W'SNT;��c�M��O;��1�J��1�����oí4�3\����� ,$����\�3:��7�9-�3t��K4ϯIC�6I�� >�����V�KX��&z�9�Mi+8��+x�/��DvG�6Nh%Ǩ[MGV���`3RҚ���lS��U�v5~@�?+�,e�CBZMd\k��}�s<����7ST�k5��(�o�P�T�I��|��sf�&2��7k����E���O�З�g���/)Ȓ�I����-�݃l�) \�aKK	�6@��Z[���ߋ�C_(��0�,�ˤyl�ـ%�m?�)��Y�c�_��=x���>7��r\��có�斱����bCz�;�p�7d�Sy��Ǽ��f늤��7�ւ,j�QG�+������`�]^�Ɍ�g!���(���$e��+厼�BA6]A(��z���_u�l�v��Z��.�=/ӯ��#������Lr����.k@��*z�A8�e4�����U��_C�~��7�.ȝ�3ä/�AP �����(��c{�����I���b7�dVaִPQ�
s� �V��E�g>��v���
��4�]
;���������X���v�����'�7��˨�_����F<���K@E�y��,�q��r��%���m/��!�s�:3NҮ2K�[�lG�N�b|2��L��-D���]��M �_\�}��0F��|Q豇HT�M쮶���7^2�����V�͊H��)Z����Q�$�9��%�����Y��«D$S�Qg�̡A�l��>��ּþ�<�1l�%h5,�G+:���b�雑}�[������&���j�����3��*��i�c����9�Q'6[o��:=���^�c[P�$��N,��s�ڄh���T�ꣲ���e���gO�)��e<VI����JC�:g�M���Eem��0��b�������|�4�e���E��W�
,s���d��	�	��Oj ���i��to����dۭ �U+�e��$Y���C���M�N�����l�+f���C?-]����_�ϩ��4��m :B9Nb�DG�5M�!�I�r��l���R{j��AQo��ձ�s@�ӿ!���{�eSr��ۀ���S-+x!����T�r�e�X���4���S��
dh0���7|�P����ߧu��H����Q3������ ��
tAwj	�|٠"'+��P |Eh7�&�lL[w�O@�N�n� _m!#C)�:D �	` ̴�F�e*�ʕ$eq�D�_�B����f殞|tھ�@Ta��0�i��p^����Px�d��Ͻ�ӵ����<�zu�&#ܓ��M]�,}h�6D�����Ƨ?)A�З��y�,��D�?p��	�ԙL*:��;CH�7~��Э��|(�!gsc��8	Y�'�]G�B���)�2<���(��'�bj���.���5��Fk�|66$��د�SZ�!��`q�����~�ݫ=�k�}��&kb�Qj��>}}|�����<=�:T��3�%�ݵW���21��+
���/�}%�v#�P����s�-Gv!�N�� Y�Y���@@qN�pP_��W��K�:IfF h���~�g^u ���]���i�z|��:y�Y)Y�z״�!Y�C�eo��RG�n���l;���0�d������̋o�u.�2�p��ki ��*l�N�����L0��IZ;��ׇ+�:7�մ4����5�@�V�e#5��:x��^2*����In�;�v�V/��ֺٳ�.�&U�=4�n�`F���p��FP�AR ��~6�p����{ʀY@�o�RF�\��G��]��Fs�̚���Q�6]L}`�K��Y��O��2�Т�\�j���z���t�}}���
)��.o\(�.֍����;q��t�-���1��G�}H�\ڕ�kI<�Spqm�N`5��_Ь�a�'�A��N��Pl�Wv\V�qєl-�YT��u�/�v��	���g# R���/