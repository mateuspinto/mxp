XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����`p�g*g�ۏ�0�[��2A��b/D����강՞J�o��h����ɋ��۪���<s�a�;���.�b�zP�Q5�n����%���t�^���q�+�d������)�NY"�gk��>0U4i�J�em�����l>;���B���ZD2:��i�Q�[�`Y���/�<���R��FT��Ọ��.���!_f�}�r��\z?%��'��ǟ��]��k�n+/��'l���;�U%L%�?	�c57!��5�S'�i9V	��Z{��68K� ���_�'�s6ja�f[�h,�t'L92=���ns�h��a�"�"����G��B�c�H������z�7;�v��v\u���*:$ �μ���Aʬ֜�����-�+��3@�b	c�3�ǅ>�L{�l�A��2������^�##Ǥd��Z����̽'���ձ�Ce��4�����Bx"H�r���A�������g�8�
���K�����1޶c�N��5y����ੑp���׮��fauCE^�L�_��	���/��������Ng�)(����h�3>�ikcD�U�B2������X�7aZ�4)���AO�L��J���M��N�,�u���y��-�w�zꇪDp�x]GuC�~��=\!"�^r�<��2'+,�B}y��e�ѓ�l`�E��E��bQ��H@F��LT-�=��C��@m�Wڪ���v>��~찟�0ޱ�Q����.�,�K��v'��XlxVHYEB     400     1c0��)mtv�:��<:0�Hz��d�qK%���C{G���@��riNW��8~|/G�^>���v��]G�;�7B?XM]�`9P�ݺ{w�E�uIX�~��33/�,Ego�0-�7��y��SM���WA}F�����fSJDς/R����v��@�lVT�� �褤[�����_�������Րc���9
E�V;⣎���d����{�Zk����j4ЙF2����0[�����[�Xt@�4���E+��2:�[� JG<�\ׅ�
���;��
K5 `�hg�7iM���GG8%=ސ�Blٴ4�\�~t}�(5B�:��I�&4� �u�z����^�
#���(n����ڜ�����%T+x���O�44(�g�Q�����D�V����͈�YU���,��c��$��YC������D-����3#s��JIW���3��_W���#�XlxVHYEB     212      d0��9ukì޸��g��(�~�s��J��.���T����D"�) E�H������:��X���Y��[��^&Y�^���B.�^C��G��l�̅�z�3������4���A�\��#p�����p�I�W��T�Oq$TWv��켠h$SS��UIUtc��0qf�	��.�O��Ej_}f텘o��a= G>�0����&�2�B}�=�+