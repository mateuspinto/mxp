`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
ObhEvU7CzT70wgq66FUj98qfmmUPZ+3H58ynl7eg3jTWgTRK0YGmDHANVKMvFiP9JuTcbsAQH2Qv
9H6VO9M89F4lL3wTA0WRTFXUszN/zhcCEkSo8VXG770fc4fDpIpRhXauiyvFL3qTMWZEU2p5vodZ
fv18tv2Q2mf9zKBnI/pNuaNPqOwK5c5Nqiu4uhLNsMQzEHrs+I5L/Cldf4pdU2lHUPhxyulsTnyu
Yc79oib50t5EcqdIwRtSyq/qOJrTNVwOohrhawU5dobgsmjneD98geEp4VzCcsIVR/ITi0N0hW5a
sSEkzjb0lTlciEeRA33ntauVqq+MWmyxRjJUkg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="XC1qnibC5Ob91AkJjV+/U9Y+zUF+Ls1ny2ogj7+quQE="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
yHj2fn5xEAsv+Jz0neEdCvzMT6sGxxIrCwFJneFuVWSScbGUxri5Ot4HYUhjN7J68mewTiGjdval
FTTrNl/VevTgSgCqu/9qb7n547X3pqNf55tIwD3LfxdH3FXZdcZp0wnbv2e+7x2uZDZ6WHhz6XfD
SYn2ANrNErmxfxffCWZ09LGrA0k6Q8YizAH3yP2/z+mPvWgSxt6ct3ZBYznQQAaMUS6rtYFtJXXF
EnqpZaFksnstoLrnuxBsB3/YTbSqNe4wZD0rsQzT0J3cgAgAA9Cq+LdD/+LuIEWunZFg7B5Mqcst
syoOIPrVUSkx9t4yX7z7RL0jIptuOlo0/kYcHb+rsfYGJzXGaRF1cT+zaRgVDGv0PkNDSIcsIuF+
V0mN2KI47HyDxcpQ/BCpRDICB0gLGcppQqgHRAtlPO9weZB/3gjJ9K5hb8V3uAIAhdZx37ky6+fg
hANN3FLfMUwdEnSJNyxmlUwzh7oDkRaTO/J8mxOTii1JjWZ6nTQKWc314w4b+DTYjufQhuA2VEs4
fhXOjO3+sSj7XHc1zFvWb4CXfMs7hNxYKWhxVUUwePt115/S04J6Pi3uItTHZaL2KWv2hnZY/Wcw
kNoMghZOduocAsFY0H08bWIgHZfH8m29pAhqw55uMhh1bEbRnJh9RW9FrxGUCAyAXaCThAwiMMrY
xipWsb/yHLnUVoxOlB41YA/X/vUaUdTOHgvWu5lJo7dWzMbhowHBIy199mlzhsmpgzRLrYCQCD0w
v8k8D8yvLQqDJP/F7q2zKZbTe2NU0FNWNol1jukyZvWjr4pWCVgYwTh14D5mpQ19trp2Mr3tUGN7
YTNyHjrUy8C968+chkKQMnVs7aE5o1JASB0fzDjfMvZn/v7u5aXNpbkMgiNMezUue2yj1qMqnQ+3
cRLimB8LFeUDim0a2rDd4rOCcWriUZdI6Dg4vJEgCqhGZaJcHOM/7YoFc34nZSH8CIHru5S4xk4G
RnhgCcidXOEUXdsE62Oa5LUmTrlA3w8m9/HBfejvYHK4R4yiRy5Mq/HLS3Z9IWKFJN8073vg9YdI
lEqFOzqJnGtR16i+eFydTT91urCihyhcAivNgwfaSP4tNz046FoP0nABoTdK+BHdpdK6r+L+ATfv
JHM0SBRyTyoERaVnCoh4e73PjKkdPFqv+h3IqoKgFRcD9XBVgJV5VZTlfrK6sOMfDzO3ZekbQJ8T
E+Khf9kVFEtCxQqS5qWoCZQv2gtTeDFMTyae7XRKZMuxyRa5p++6zqYkPx+LFbTKiGIBrXzAYLWU
5Hbx3GTmP97Tdzkhj0otjFM5Lq6C5/j+Hbhb9iPl1dLN63Z1sPn38iZB42qgcdmo3g9cMGR5+8Da
bNBUfoJQ2+o+iM9RZzMMgMtQMc4mP/+9R3Vh3CGPHn7E9fum01vAgGk8v83D6cr3Fgg4iUJBzr6c
AMiYUDr8Ta66XbSQMSHIuChTm/mW3R83tMvKRnKXpjenhnD2R0kkBk1+5NNvzykDBy5DuQoxqbqr
/HuJQBsaM2SqBjb+kxhrH40bT+zafovoBaFj/y80t6YQzfjSWoUyvSBFManK48d1DN9t7OVZxHzw
BE6CyT0uxWldXR5NWHJ6w2QWc/hZ+tRoOCpwBh7BuB2EJjnnLzs0YoiEbgvEuojqfbSR+HuejJKT
NOBBjD8ccAzoyb6pTZRsA87ciPzlHPwy2uFiELlGlAAZUlM21EcpdxUs94FUs0cx/DBxogCYuwYB
L7ACjjCZtkYPy0qgWlfyz2tS2DRup3mzKukuY0V/wmSygONNYuxBUB1cLO+qtmtcnoyLWWiO/Cs6
naiYKUEPUXhvHa+a/evsteR5nv33Vslf9BjJPS4lpfGKAZ88n5PaEgxMtVoiw8DhlSa5e9bkVRs7
DhaS7qDEQlKFiPp6eVsMw74HY8uz/2U2OmDno9ATwIs37znJuPYdBrPKBdSx1xlDtSvTbj8GUtnR
MfKSRwzcLrwaCZxmv5tME4LhYjVyBzZ8T5vk1sYSLAmJdPd0Dkezdrbdm5mfvJQILSKmV4otsA5P
5QjKjuerP22cUtirnu5jbfEFgsgLA1IMqRlHvM7Yh/tILTFtg1YweUQ5qFSdqCkAAnMbEhvkWhAs
MyioPynCu5ejU6+BNYj3nui86bim8vVn8N7Cgj8QE9zIezCBvcp6SAc/MKHfvCI3Wgk4/VCl6B/C
OY0aotU+h4sQ5T8hRfP8SdOIX3ZniWDhNPXfZZYoXS20+RkeHGM7Ts5Tf6ZXfzGS5Sf10SxDV6rd
lINc8nR4TZLNASeOSdaZJ0JH/OjfjrgN1NAqu5YHVIcu52WRToNYF0Gy6HdH+rSyec1jAAXDCRhW
jnZpZxzo/7dOlTEFNobgORdY5jC9mUxj29Am3BoEuRupBouKuCzRUrdp8XXk3/sECG6C8UXeKUz9
B0swJHAYlWuSXPi0Tm5X7gMWzEAK1oWr12LFRE1IfHz3glf8032gOwewg4BgWys8JvG5v2oEGHqq
Wh9qZWHvRLPPWP2M6JPZrht6VIiV+vvHtPwKYPCOcuKID1xZr9JrK5ATDTAT7jF+plzUrD8gkpzH
ddgddEwiYhA8XK141x03YB2+1QqMmV7sTXiS6G9kdcXNxSkuhR+1CWwPZx02pYhk6GkBA91StKM6
+Mlv5Mi6j4d05cZHK5tBVDYApRKIxi478QOLJAgRSSPlTwWPRDsSbg+FFLf+UBzUAa6mVvhA03nI
/Ish5VwbhEUtmSv8WEcj49RPR38VN42M65D92ksBujbt+9sgHSTpLdt+y41NEFyeCUfMeQcBHlS5
WHNf1F5rcWihoRn5gnyoBZ8n8jfjP0M5+grQ0D+dRKr91ofKWiAg3ooyIcbuyVFJJNaLTg+e5XXd
My2VgphAy7mg2C561uDguoCuCgw3Rnhe4hsRI/tAPzdfxPRP8SW+Rr3+aYb3D/qkJNJmNmUAs+1t
UFYAO5WNjydHAMTu2bVi8lMnGCQ8fVM4qM1AdoYq6/da4ZeojALYCsjWn7maiIFV1XqESblIYSg9
W4uNLxRmnQZM0sQ1NgJXcSRQQTvUAH3N8KGSbWVRhM0ZT8pK5qhwv3u/L26ppzqKKsQDRSLZkSea
8xFDMM7F2tIu3v4MPhPT34u08thTDkbt1C+/3hKXvV4QlSa5LUwxWkYZOukL/f/lCeIAub0Grfs/
p9LbDtoYC1y+758raGNNpJNBNwNhZL2zV4VR5aT4mtkaJ9vxSWL7e2I8l6p9U/a3xs+VfDp27tbb
OQYYwnuC2Ld9JsCleM7t7FaISV5F1q6u8ilkRoz+Z2AOevVfv66py6zvU7pIiarEg73mxzT6YA2o
qvgiL4KvK9TUMAHwQPO/a/QlkfwUI4Hh4jk4fzgKIjWQCz4aIEHJqE9c2u5I44atlXhICRWUetle
Zk63lJ+eqep2/hqc0McEea2IRnzGxS5fhy9c+57G9MH3j3YQs7GIHW7PBXUoj9in8gPtHWyqTNOa
6rpyT/V1DbdFTrPM2vnv0kYeiyUm2oWOyeMMUTKtYQD1heNf5jVy0isfUYOhLexeSm/LnfkluNRf
8blFXhjrfVzQVLCMrXxTVdzvtpbwC3pHL6dBvFOGyvBxBDlC4FutMrCdymtztPHy584x1R/owqE6
gyVxnR1wa3gQd0qjLK/eytDFNqTeQpmBwSERqropx/vJ2CZr4pRb+jKmYoQHKHN3B7zt3U3L0dQB
dfKK/VEUIDDFm2+Q0hVLDk+LOICSR1BIkEScbKvZzXZVXJwfE+lTtRoLTSg39ejMPTJ/aeHiDL25
G2n9IoqDQ27NAh5Fvwgs8tYsNvW235ym612cz79pR+DvsdeIC6rZ83NNhvJdSSFMpaOSAK9lLd4d
NqvbH0SoL8XPXEO686/KdGIAxYv2SDWU7RA4GI2kiInCvIifaWPZNhhWNL4XjaSSrVEDVDhWQ9r9
xZq4S/AG2HdVPjMXnoQ+i6IyE+DK2BRrNpOWtRhZ62kon+Dpnx1gmBPxfPEuCq4411XDUpAged7I
rHTLk5E83xizwqo+RgvVskOcOSUwDiCUMZFZRzmFP2/K+6HdKvSf3Enrmc+4mDZHo6eiMG57eW0t
WnhG/ehfdPmiX8z1mwZX+w95nu+o4K2WFT489gG34H0iTmWkMfUto7FCaU5xaCEHvI95iPaVVFkM
A3e+GfxGPQ8DTLzos8UHqzJCckoGxMrWKQZwArP1k6JxzJIqMjqCeMwOU0oxYwTaHjIwC3kT6W6j
voykNYzqhp7DfqNcQ5fN9KQ6raaFPoWkF/SmYaZOii1sonZsRliEYcf1j54nHTQgR8fH0fMgQ2Js
LpCOQe78DRDQ+iRBKrAMucizYdL/couIEuGkkpzggjuobs90mtB2YFreZ8kdc85wRTFe4Ep+yJB3
+jhezDJnUFmhPq6fQaWATubIsbd98iw0HoWIrfioYVI1dTWInyK7zxVYzuqijxFxGQ4nJ6OwAjp+
gyx/9gQailkpObhFR/xGE4pBdTlcto+dd1MXHCF+ynSvCfhM+KOb6qZMbd62WpM4jbgLqufZ6UxP
xfkF7yQkXiXQb7m407Bku4z4QroD4oGlfdzyMsnuJQk9cFzsl2x0VF/VM8E1UVFChx5i1OreXIyb
HrDPO5VT7bwy/WMDiLkJjkEtgo6tL3veKS7VJdfUHAln9aHnInm26KtWP/3kwt9VGYocsIUkeTnd
YBVPo671x3BPCW1R7/v3vXF/tpVH4um5LA8GQX9LTHP+tQ5AKsxM7USB+5/jyz24QJDs4DjVMkrt
Y0+P77gqFMfNxJsROwNHJUQgstadbwKv92qu2MKDrqFl8L2FOEzVYtJScl38d04sS9zwNZXe0IXo
pXxAYMPMCu3GOvRhgYHE2NZMSzi/XnQ7wX8dCLJzuK5xSd/WZ40iD8wY/GTYQyoS4PL8vboj68LE
a+cD4B/bG3/kzrfXav5tFafORMvp/1KXmrafcvbACaYVEDc+/yF5UPDxpB5gKUeWVMSR/KXld4pd
p8b+2xp2LGSi8+MrVEF7kF0/FFf2jAHT5OUXcZfwCcrNAbxzSVMTyd3lxDqo2l15u8M9r6yJD05L
bxZqYdxja0wtXAJ5gZWLzIsx1MaAr5SVQJPp3tbYW1kc0qOj1hI1vCSbaSaN0ctOI4GufDQUbBPm
E++yvjWDJpdVzIdWD0p6vLeVlU/p3ba5Mv0DdIYrWaMccBOtZiFp/DNJe80tuLCz4FePwBlxew5z
0vuDs3L7ysXYGFdljNLYOYVs5MU9jKxKNRi74szfC2IwxtvWXYOYmANbP2Eangmn0T15PzkiP83q
8ZVyk8Go4P89pW28d8BtZLpS/lvYwZYaudx2xPvlaWPKxm4xFjhs0ujdBPh6WSyCPtXdPZeCvvMf
LOOfQcdEGXtnV+CWg2AgfcK30tYsMmMsyXEkkgWSNo2/49mxoCZnKRVPMT648MhLHvtwvFsgv69m
nhi7pKCpvjhh9xdH1aLpgctr8p/fhUlM5EQFbnSXyMFUlGgx6KolvVe/EYAop2pgocc6VaHmpq2d
w/OzXav65oworvvQ6i9XaVilUpwIcMwD7PP39NewXRIsrlKKaIoyfBf302+GsWKOfxb9YoVxnO9q
WK+5O0kwzMzagKP1g4JyWbGAEQD4VthKNmFix0T7dflJZSXdWN1pAZbRPVEcuetfk8M9RqtpzTit
wyTqigtRc13AGoG4x5s/T9NWQG1sUu8kvwMTGo3e8KEgaYaXHsWb2pQYe4v+3yrq4wmtOVrOSWbd
s98h9Hhv9/6FREKNJTuntXNzavHW7fYeUKYUaN6UNDJ8cBzEjaWwevjew9cL9PIeo09V/WXZiuc6
g+ItTiRFv+KBkumVx0ze80a04nUWbDtOfiOizI3yPhDLA2KWK2JY79B0wcXVRhQZYNhoKZP1iPVD
HBUv4G1lE/HdQYLVFEeuZKXqO9+oXYjtPcf7pB43YYKjAv3rR/xomEcHXET6UPrBUraQA2T6GsZV
Mj0Bc5wezxb0FkL2vPzqGNThskKxvt2UBNZwZxAIx2nzgF4xe8wY6IwwCT01RNGLbFofDVJyKQ6A
oryFGAUQafoJCjmfT8vYNHFVOzjlrQQCxFoAIzLLzqJSANPMDr113x+t9QuMq4FZtotWCABSYXA1
4RLEybWHlHHiH+PtdnTZGSuFGlhC5ZKl4z3lJADiHqM7t56WXxS+6l3Y39pmv9NqNmScI+/AxDR7
infh4FVNIMv/nrplx4BxSeg1cCDz4dXrJQ3hoT7mQTnBTEj8kyFV9jfhsaspGiYATl82fzgs69T/
z67bsopv7Jl9S/7x36jECpTDMK1Hp1TuvxSnmcHL0ugxOVOtC684ETGCLsGZcf0wQBpwKZZoaiVw
FYbrR/8LiY3J/SkwAmZHFIoAttKoK/HlenO/FhNFmk0oUJwWNlIzrvlaqO7BmcVqXhLQMTAG58xr
FMtwpsJVoihe9eQRDRGx/MvrIoTFUVcofArv0S+9diM+JbP4S1i2pEbt4GAn9mVkZABA85jCIvQa
rMxZsb5WEPDYjYubAOJpLTsdTKRJLQJ3B1W9OH8AJZR/Btk/V1+fEwQwcBs9/siP5WU4a+7201k9
ZIxAY9rwrT+0lhviscb7x20smVT7Q6rNyth+lQVn5bqqux9FxKL/hx6aP3xqD+jJpntBRyGDNULo
dn6TX1eNjANvZl54u6tF47uQ+cj22j8L8PUAYzkKYf4H1HvkY42wjjLXuxT9pcD2/Z3wzRaA76Md
OWu4tj4nIsB8Ilaw7K17I/kSNxcELR9Equgi+LTUtSKTdQTYrsUx0R4r22SF+ZQbL+kXlOSogtZl
/Khm362Q5uZtVyG+BbYMMX6/HC5WvFj7AAasCW8WxPUD20oBja/6tF3P6GNTEP32Qqp0i1Ap4zKX
upwDsGAr4OAw6xPNKADTQZDIumfxenc8lv8pMJQ/Kora5Ht5y1KmRk1v8cgrxKHFars7l67zj8fm
KIy9eTC1XO0dBgSD4qBdUty16fk9xt8VO55FS6BT4OXnhvQFaYjQNSPh38GkV0rjLGGtWfTy3XVI
9GVKT54wU3kbKA6ZJjP3eKpGD9Hj2e3avk/IGO48qJwGkhP5gGh0as0WLIOSMi5eR6CeoM9rb157
ad65G5Bw+q0/K8bVykIV4HTviLWIWuWx/ZFmWfY4PQwhGzvx3k+4VmwZva8dJ85i4qhGBHE299X/
xf4oxo68a8mUJrzD/mYEx+61T98X3DbE5+f5vKXEkUsDol12c56A62D7aPI39wmwWqHSxFgT2u30
6WqfCGbC5jAX5BQ+WvhiwQZWdH8w0MDygsU0UsCzis7rOjOZqY/+ZYAOp+0utU12TZ9piVZOP9CC
ZHCS4wNwrZh5ePh3Yrs/XdKKiAx/bWlycBykOjLgxWHOFEJ66qzpV9/RMm/fmzKK2lJrBsBJPaT+
y64z2X6/aqcNYFeVUkfDv7idfewdtsHYbJbVFdYo9QDwkmcb7DzTy5ueeb9BtH8GND7Lvq5z4twe
HKLgErn5Uwp+Mylo1oAyl4C1+/qUgTIJ7nBpc5GOU972UuQ7Qqd9b/eTBbQXidIKR8fRt9DoGpCL
xp6j5UIAos/2nM0CIeXwLr1JDGShxJfXIPKHRdlLbqzBG7pccam9vfkX8ee3hQIkDtN332XD3VwZ
bV+IGP0h1VJ/Xv8JGJjNADGJW8tE6VdZQ3EbCas9S8YXxkSO5Y6DEwraP9sIl30yD188lE3oJpq7
MMSfnXCO4eKFlgO41XnqLH1K7T4ighhE8uoSA+m5qVOjwbGMgosrsx5ac4jR7Ara00rR4fnEAacW
d9G7r7u0tTU3UcinEgC+DdGH8isBnBzhIfhu+d+gTp9omNDdZ+cRv4LjSHKXDMehaOagMBuA3ena
MuA3LXBhyh7r0taT76FiGSxUxBc4tuXP+dVu25CJ4qK0uefVWevgWgJo1mVDptvRFXfKmfNPKAd2
66mXo7Bxq8biMKiENkAB8h8Wqa18gwSKA7iSHIGyLilnuteyD7OJ9nFZdszlSkBa5WtJhayLfEqv
F38w2qbH0omd04CtT/FXg+WxOANSctHiTK69RjuD2hqWOEcMdAuy57VZ3qCo4zxI/7pb9U1ScOac
xayKyn+4D8b+I/KfWfV/2VoDBGn8yiwsbkKdxIFlJU4hD42oljAiDNyMTlZK2hBwnyOHuh6V99aR
jFNdRERKTonU8RPayyi5XBb6sGEDPRuQ4xbsO+OHSez8B2b0udmPvyHnqRh8WaBU3JCpMxFl79bA
fYe0biyZhEVCcwf73sKxQfDqeiGp23Bm35m+hRAr7lYzhDmwJYLv9dX2D3UV6y1Wmn5HEhb8sg6z
zoQyue3p2jhJSZ6Jx8Qc9dVepFAcoi6I4fg8Ew+CrJDUw5jNyCqHtVHkrQTvD6SlroT281pqdP8D
+LFNId14WnTbS/p0qC/G8hpbu89pviYOOb0P/2/Ifin6jWRuvDgaRlEesJcNnHezG9P9N2ulMajo
SnY/Jla41EZhWwEhgyu5TA==
`protect end_protected
