`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 73904)
`protect data_block
31N1MMnqwvl4w8xq8xm0iP0THu9L8iat0MZsTd0UPziAnVCNVbNxFl6ZELeeB559On2GQLs27inh
fCJZHozVLNHgvxDJQ4pqd6BQcBGPPXKb5GqODIePLZhsA7zcfjbecGUzo+9TstbXbbMXo6SIi+SX
xjXNGb+KNeTFqfnOP9IOnInm5YfJkW3XuHlLlakfonEGO+NQuMH+wVBO3uXx8rNG47aGNG4y4Ghi
bqfAw6D6Qct+NszzXW4xDdHvI3rmF7h5dTpssWzDSeAO4j13lDo6GxbCXw75YGb/ROxuzzjPmHV1
DCrOvooxSCc60Zpadn1VIEqMvZHxX6m6GVXkin9JL4yEj0OuonRDlQznZG6S7ZY8DpzMw+Xt0BSa
DS7dIkubk1rZ+BAByJX5m3FK0mbaM30+H+o5GRLX719cR3wurKhvcZEAD/hq4UtoXlXkz2pMUx1S
TLCYdPDe7UaR3k8uRTWi+uxwO/TmnHmlnU2/+jnj6gAe9el2vJvhGHvxIae2avuyX2DHoFx8+H4M
ypkOYwzkksh1YS0av/4XMGf/Jtar2Fbs13z6MRTdQFa1ChztffUMcWbOJWK3eyqJqHKW5Bcuxj7F
kAuga6Q3OhC37fxfCQCyW2cBki6OHju4B+T6SjgLxALzhwGMYdhO1Xavh0qmiBPdsnfSeZP+020j
pyvQB5AJVgAKMRhDooRQgr/892ScPNXRp3A3rbSNc4npHarKz7NJMOc2aFiPNJXV/DbOekBP5QdY
GX1RtZmYrSDXsPXnSVCAESbvOl7w2jDPY9yLeoOsjTSgkJHVyWZ1onUoWAoL7jnR9p4y+FcaaRTW
ZCe0cYQXPqTBvDr+SsjCnA+aENQvw34sVBFIPqwAM9TFD7yF1Pzjts8TzpJmjzmBc6V/+znY4LwJ
VRQqTxrQu3TDK+eYuDqEyNCYlzQX73XscW4f7YHzmLFJrEMMzCHWOBF1WRFjwFcQLvscCI/gX7fy
AVuBl6u5f/ZzyU9OfgRxqSaK5qVcVkHH39B7bUBEB1wAyGjDfn43rsK+KlNO2I7zB2HK/K3UfuIw
fZOtUk+uE370tbihgYEGfNX5iJsp0k4HrouMlPNGL7YrTWuEC9RrB3C5jjkyDZCEUDSjoFYDiMsb
xlXb3yQxpfjTAD8/bOPmuRb1h4fMQczI1W4pknmR4KvgNMKcDBHEMyCA0s4VqlK4ylhc5SiQM5BP
QBRvM7M75S6aHyquLkKDj3ySMjefRNtKpSiue703W1yiC+MEq/qxzB5PbRwlS0inuQrSiyV3GjmH
cSE5IAQA32Y+CMonRpF9+sYdlR5I7FT/uF4AXrGDMn06dXJdg7CXZyDErv3yr3FXMFhWhVeSq2Hm
kOOqtGb5dOhgtJegSWWnfbeG/jK6JoBcYwzbVL9WHEc0jrCXU0o2kWMsSRar2heLeyJplLB3gWFA
Z3mAgQS7hA3wRaC6iHfS7DPpLz8SKO3jrDR65eTLNqoeQFiTAhI+0eTubIjtkoGO5uI0vmTxHlRE
F/6UAqrU5LrbO9+nBf8t/LIstUGu3SKBGJD8jcsgVPLF2n+DoWP6t3waoKkDY7G+M0pPk2zS9Ozj
u2Px6NkKHUrzYY0MkwRXwmQVTDR0nyYqbfY7MvrSa4VfCXVUzXSujCXBQqWhZplX7zfHCIKyYcz9
KfSjiUSBRjmKlIROIHUw7y+4tSI7ABwKTAgHverxqU/TZXMxf4CMFkUb/FpYM8Wtj74Yj3KAHjrs
TZTdsqo7SUEhoH84TQ/YGe6VWg9l1v/aVssxe4IV0LJRbdgFp5TNVgtKXxiSP8ml4FyOi7Cfo4gB
b3Acwwn2hED4Q7E4hDpSnDUsOlDgBjMlC/fCHB/kmU3dkmaqEDOO5DCqJQ4B728BsXGY5Q90v2HA
OL4Gt0pSyNy5pZ/7SmzPdyYEubslWtcwfWEz8Gm/QjuzP9b5Wlw0l6AhJyvQ3XnyT/s+v4kDQFkX
oEWCPa6TXpLzGiaURsdOxTkrUMJv1yq3sAg6XakCukSoaANac/IkVBZ+s43jVcZmlvJO11YZu8jw
PzaAgNg3AEixrqhzgRLq9Z6+SQbQ/JztQDYCD+NNDTwqwnlYpT9X9/fHguzq8SaivQqmT2zN1TtR
E6N6+PgcDx6LmgcDGu0XRRN+vSAux8DTCprrkpmK3uU+wq0jUjbKHY0ACiwCcGP5IuQZ2cUOT2sx
is6p6l0U9xyyKK2IBYDHOx5QXJ6E31DCIesUQpcrhsLd7y/nVFh85dxr0KUCUpKCv99RnTPf6G90
OWa9fyRd+a6ja0sElgC/HGYvP7vmDg/bcX3e4la7GUMOmilMIddhXpKG5g+mY50UwJngF5ExhnnG
fJwMrjpbLMejVfasAmmVSTh9skjeb9WCEnOBpdyi7fpvhvR/VtJEZhmXxeC0gZ35YmauC/tQdvnz
oI3nHX5H5lL6HCSazmlWxybJ01H1+4G84WaxW9E9EvJoBzdd/dWAPYKaOeqWzyMqfn+noDWbYtH4
2FQFQrNo81Fyvz27rTZeTW+JIM8f2v7Dd8jvNjqJAasef16CbiyCWRR9JzUX/5uPjVjJ2VKPKgId
VrZ9cB7SJRm0O8nLRGj72dSDdpyGsfpzpjcIVC8AKb7MaHxNo4PxujBBcCXF/we3nIs0nGQ6p6aR
LEJ0N+ZRBTs1Kmq1Uz4NDQe5Pd1WhGOXo5KMdg+TrSt5pEwWYjk1OAtR/uj7ZdtYcP5N3/CIooye
pzjGUQ+ph/utFaZUnA+OIgiW7vCYcU6eMJDOfNQ2yVuFV1qoiJX0hUGOfS3wPAx9mCSAjyUjS59J
+TjuA9mEExyyirbYfBrMee1CS2OINx0Q7zJ1RtARCuZpOV84OLCRD6uOPmEnRFJL/AHcoIMWdwVR
teqDPjuORcaSSWX5++cB7hELAbUCO+vIAKrY2J3ERplZ4tjMbI0MyqCox/+Fuc7Ff4OB1XsUz0Mq
Bl01ZR5jF0khmhS1mBIsM11nFEEicJnj6wsNw9GhQcBwEUpU3U/zve3EDezAx4aQKXgkM6O4mJ43
fMQNBbRhkrPWxiZkeqr/woMCj7wlctJEcHsbxmzYh0Lnb7K1yiywJqP/Vu/xcZ2IBBSKk0HiPMLI
NHHZ1qUuvb8Sduxxhu4Mu/WvWhmDK3VRyJKh3yLtq8q4o0zZMN5BZC8J6YdubsPmnVqgCzRCW/cG
fg6MuIX33W/Yxdpq8NTzvPRoZZ55dKFRqeOVl4PbAOGFExidK+uT7Fmw88CVOLiRPUhRrDTYFpbB
cu9yl5IoW9/OGWhGMW8VHhLbhuVxlTby9cPSFAiEnfo3nL4v2yd7V8dHvPG5VZq7deVDRzF9VDik
zeX2hlMbTnXm9nJQrlXx9Dpi7kPeiYfIOMW+uMZjxz53y+KlPbWWtog1VNGp87JiD/VfBEXl+qMH
LlxoPEWCRvIbOKgvafCBFQRmL7KtGtB+611BP2wEf3eCH5CqOiqwjtMjTe5NZY565pi5L19Awvct
MjWnWBpEnFUWldf+7CD1ozz0ukXszlruuzyDtRVzAPVFpi99NFvukjUrt4G+P7MJCFKfd1Wj2IPL
fgfjaIFvyGF9b/wo/2eJbx57JWR4nmXKOYPjxQFDzoClIDQWAcf34Mzn6f94kvVflDYg/C1BAdT8
jzBfYTTupb8wIJeJw+TnDE8kXrHfw9wd+BW9vdpyLevI45hcH0odnuHSXnbAMN3pjB2DcBQjF1Ga
FmLQlBdCpS7UoZL08qFEayql8zKtSJBMQHZ62PCsxO10Gu0W5fT90SSl6usa4NHL9s+87n/4IThi
Y/J+QEF/hq09aHjLgYZnHaIE0jvubqk/2AfJj7k6KihEBZUH3D0Ve9lpR9ctdZT8cHeiJ2j3I7ys
iIGP2lAzfc+gYYsey1sB48wC/Sk75zCztS8xkiK1wqtma1kX5chcmkeoX+ucajCKdxvl0By8AN1Y
s7ss/+mMYSjdp+Kk6iHOKmvHosnHEcm33zUJJEj/19N7ex3KR7XbGR3BAnqU7PTy9wxbYF2k7xLc
rZuzPnxFsCu+Bhu3cNv19sqpW9CbJqVcIqEh5ZaeCIcz0YUio/GxGMmKVwT5eDduapJT2YGX71zT
f2zTu2V8h2ERFUOfSGEFejEvPbyxJRCu6ps0qOJH8L5zhvdHbAqj3mdJquqG9tLbjWrU4m/j1i5g
ngMND+qzffLcP1FRtxjmlBNT/U5583chYuI6wB7aMYkELjhKFIeHG3RKuE8nG2YqXSxmLCh/40JV
C+MDnmwOyT6waeb/pkbm3F85a9PmXTog9aEw8qE4b9E9Hh17kcTwO0K19yN49Zkd/HrLlx8S1dKF
qBoh+WN6agDiS29c1Lnr9mVfKc6Eyvonqg1Qxfr3kFKesATUI0D0QkHjQ0jnlkC8yZQ/X2U54niv
ihblvde3RiWbBwvWG8NrkFtn+NXDyguNrTjP74XiKuBuwR9kAh2I1G+CVYZFXG3TEH/DufCbP9Ay
Uvb2++EaOW+XCB38r/DMq7ZbgexV+yUkaIubgDPMq9A0kk1FMdjxW6SLXXGf9OzaJ/rXl2DgnERw
mrmwi05WykjoWQ9zA/kq1KLLTB19v09sxManHPYgsBSL3bzI2cF1ItDjTwSx3qGvwEWGruw2OQAl
7WB5rj3abG4SINbhT8CGTP4TePUldJsitodV/sSdXbAw7OCskQH4cA4BqoTRJV+GiCiBip8CGotx
GVU4mReKUbmmM/m6PoY2QfhD/h1iRYCFrgpFJDeYrO3mNRJZPivFYhH4hplLWTk6ydvGwAkd6maw
hPIH7P+1hJIG6Ekk8LQbNRWWIJa8cTTk9eP5b6wkxvn7hra/ePV+LKfByVMdnf5cJaTDRZ3VMTxl
0MHvTtcOtgVWren8+8pgQTOJ4K+cJxHRf9VhZ8LPRYSR05OVEUX8vHbQLWbc4evzuek4yQUH+J2R
KOV7CY3lnZ84LCaNpTYr1m5qbFYJ7TJaRoZA3CElXGRsWhrWSgNjgXyNo0JHhlzaw/IJ1sC+d6/o
kQQrg7Xysgrl7BZxoCbzX1bce1G/X4pstfcsJFTaxEl812Ani3nuYvmV1MScjnoPKFnpOLslFHdO
uweRLJDu9dVv+ILKtz+3J3uB/GhQLpg8h8prUQCh+X7l3sH74uEhq5pD+4Wrbl1Zwg+muivE255g
hfSywX8rgiCh6llOXMUAuEkIj35kmfs21xVj9Any4grt3eoApG2xXOmjmjxr55NR2xlGo33hVvh4
7WOTzpP6HnSLQite2W4gQtCi0jP+AXjJIJNtJVu7or1BJ0cFkS/cwKlQSFsV9vHg2UnAoQAry1+C
VJXEzuCuHdmXKQcIbhw56Fe4KWSSVIpXrGR4CXvke3kbsa8RZxi1Tirr/WuW+RwdkZvPk//C3U9m
e4kWbnkcqZjbTbIWs39IsjxHO6j4jMasP8YbU84+HGtb7uHRc+zF4eQp/6VqXAuOU3kxiZDqat6p
FBPAXzXIN/oxvmwkv6sIBkQmjcQUsAqhRwBB4fKPlQl9u8RK9o1XNS7+boQWAnLjVxhkbZHsacLe
9Ls2d1mPoBmUQYAb0KiFkevhePw6nIvHEzgVVsIxPIRDA1e8nNrMBLafhHBWuOEQLIAaN/+8mho7
BCSn8qlsVpyqLnc0JBQ0FYNiBz2BhohU5tk96eMbHC1qYP6w3xmtFoup1UlnLxwxdCjlH/v3Olix
eWgI2fGCffTwMADF+kwGOFERZLz+GpkY7hAadXOOxNEDWeXo79am5q5fU/SxEZ7L5/1t5EKK31MZ
MdZR53Jy3uBZvDkBWI2N63wUT2aOApcFNVcSYLsjFU5pieypN82ZkWKJifXr4PBMOkqZzDGlisB/
dVtrp4BM8tAyS8jiB2if1QYHmDmiXHUBSqRIwyk4TG6dXVvgDFE8Fou24DpwlOg/gwD2YwxbzyoB
30/K8sjs70sFJdZMv4vFZBs8obwe5iolYpbkl7vmd/d8Y1Io2ZszWTo5LWfhT2993MtFVrdNkwfy
lX1yvNK9kOH7YWqNdDXy4bB9lqSEKVknHBvY4NrZyo0aCNbOJUwGnAN1rq6q0IBMkkchGKXoAmpw
ddslou5eBlHcjqovWXPagv9oaGiMviNbshV1BeMP07Ir/EdrQu2f5dk7A50Yp2XgVUfYhondCzd/
2wnUAIA82J3dKqQnfWQphTuyYnA2WUSDEqWhaBt6rEseDcj1Dr2bLDkXdxOoGkb8v9SqJxeEmrSF
zLNBUuySk37BZOGKvQ+FpkvIIKWkGumwTF0N9/NnXULXPN/kl7zLSxhUPAdULTtYJj9FJp2SXf3u
umTa9SlF9RBBV11qEbNipyFKRVCmQND9A7sfHI7IKL11gUm1bXvFcnMW11yHwvLql7IFGUaWElmF
/O3HTupiv9f/VunDOfgUJnkZYqQj/b14RJiPX8muFcKmJLuzZbmpBlTmINYE2lgWIrB4+iUkWa/N
rUgrJgYvRTOwCv/HRO2NOUBItRdmGlM8r/UTka5GFvbipWl6JOHnz0kNA+3Gprnpb+/3scm+xdNc
ZLb0iDCPzCiWbt+frRGKtTy7NPZyEMY7DjwFT/7DThz8lFRs+zHkmceCWjBO0uQEmsw383cAljvz
gZ368C5otuNQutpyGragj48+Db8NC+uNWfU3g35dY16zWL6irBVcKtuLmJiAdTYVwlRwhYSPE+D2
CURluvpGAXiXlK059y5LCRU2nZES7+rT0dJt9QkZE4S9+FcaY5VvofSxEioYWgOzafTOokV5pz40
/ZQaIFMCRua/+CKo7dnnoozd8UYcVvi3U9Tu/+YM6+uLip2Y4URWETOthd+Z4UbtO2yMxbOYxQAy
3Q01Y3qVQ3rfaptepreGAwBdohvkVMa/cBa830S2wvVcsfeLsqnUMofMUk4a3y4a6bhX6j0ML8xj
YYKKMU6gOfuHofbQEpAWlBE2an1TE512A8q6nvO0JpHT7MZV/u+PlPH/bVXeY7ao/D8OL8gOCbVY
xM08aboAnBV4CfiAD0O8TlbQdorRI02FTXGISAhzVBQrC8+oPv5vxegfyRPNPK8sGmeMO0EZclDP
G425D9+kwaBugi6sTn+TWIZiJfVnHAkpViwEszN8Mc1S0DyrpSTS5RzBAwX+RTTgc/su3K4dyrqs
JgXVtjz3/nwhQ3hbUFzvKL5hUyYPXmm03650ocBsTlMwk+QD3gvftuVZqrlphQQA7l/VbR7Wvblo
ZKhjjsVTL4s0o2EGTCrqGphR+NVm8zq5dn2eYo4EBcDr9X2dRzZMBwGDmO+anZQ9cTNzC9yE8OMP
HW8By0zFKPyKcZaheQ7HW3LRLKYpN0+FkvbPFovb26DTMs1/v0Z0FlBYq4Oy8UqYXrqNUafHb7Pk
5GQn+QElQiK1mBEUWrJsoSBnOOLx5VhHBx/TwDeR1ykbydgP8Bc92EOgAhmAaQfRddeq1nICjZQg
HScW0QfCiRbazVrfdicIRGS/y6lL6m0j6VLWfEGixXsUIDoDwV2nFKR8Qe2doe4XCgaMIPqZ5QlS
qM/NlN8v8JzlYmiSVI11OkxUSrjm+Pfn9+20TUZIJPfc5ymooqwonMSvLfJel1VACWtkOumlXQ9J
tmpm0nTxc0Ng/PYDEdhU7bcPR94K+gmsiRXtseUTziScYW+/teO++x4D50PT3WGhdNXJ9biksTh4
j/gapMnVc+v8HS52e846R8C28d0PFfLD/uZj7DtXa1xh3iG1bah6i8xpp8W7VyyETA63FFwa73+q
6uy2tAZGeWMhdeYZiQK1vsv5sIurwuWlS/IVvWDWxbn0IU53Rwf8jHemKvBaohif3PHkkCC0tJfF
RH291kAQZDA9iEthKTMZYPlcwDE3CRFRrB4wDdaCzdL8KiVlqmLK+ApiCjKPnxhqvfhiS+KvFQ6J
QBWFxjEyARhlC2d96778l7iX5DpLTSGu1KZf8YKsfGIlSdu75MkbZ66d2LWvbLqD5Cvy7+58nVot
PnvMb/zuuu80nqZeq8AG1T8EthEC/vweGH6Lv0sa6G5wkDoDC1g43SQxa9F1K09o8jEN5VLKVjiQ
rL23SS7DI2cCaz4Yl/J8Ll8d2hLNhYPdOf7ZiYyZzCYi6JD0gsa0R6yTG4TBqtDm5cDw+xSbqyn+
V5NAeRaK9yRGD3W+AbDg3/EJIytdsOCjB9xA1GDWBZ+6YYMYcLeqAHUEZjtlFoiV+9d8jc4p2PkX
y7mhjXDvGQl+4GLolpvjIGQbpGJEuacJU8ooTYgHlfXukCEW7CnrSBJlSxZAicnD6l0GPDQ1kk1F
2y8CPttEPcCfvl5l/AQ+rcS0x6fa0STHIeuQW0ImnC1fC1E0Bp03T3QNPMuGAdI82PLEn5BqhSb5
mo5++C4KyK1HjKHM2zprWhQJv7lQZEaEcoDKkqY2mc5nPiyxbRp0YtqQAaxBbIXQhmudDZtNYrgw
h0GWviIorX7Q/01ut6R+YDeqUmWX55Tyf3uVsw0moT3J2YsOUgNC/ijo7O4dO7b1nW8YqZSncAlk
2LPihwQ0RKs3ZhsEOtos5TLwNjOasYPeBHXVExszndzllBDMwVXX3Fy+UMoQkrDdhM2ZFSe8JRDd
ixCvrhrP+XHMkPZTQ9Qc+EIl2bVzeClp34Qm2Y8k/4Sy58MTFYI89LC9WXhpIElf9GAjpAzYC0Kn
/dNK2FEb+mF57svFIPrQ6REof/CbbfMcZyizZf6Np1f9jNQZXx2aUv24rM0+3Af6VgpbrKWH7wvt
CwNj1/AylW+WNfEdPcZw48hG/pFrAIutIlhJGGsUeKa+XFyk6cIzhPxWTstZYgdGtCCqARLoAiqH
zW7d/X8qUtaYwLE0biPttmjXvL7X1p1NhdquXQsyrYU/BwDAXl7QZQZP5ZWoFpscS49SOnhIYCmi
VuSNyTzMDqZBH8TFcfAYjpoQfmPoNlSArm3U11tFabpfkPdk1gr0BzxmBRGMoCQsNE0eLNhVYeNA
KOw31o0HTaHhRcjltUEdI0pPsi8D2HyQZ7s1NPBjxQ9NYn6SyzQZ9b7sS5No/LEMcJtbj/LYyd4G
snIpzyBqr2047mUEWSvkEVSTgTX8Do8nZMJp4TdOJS4byHHErpYPkXi8fkIcB1ckwnWEVpWStq4y
u2stEgqXUm0W7ePOcrYIWUt9yqXrYeEXf+DJISOjUxi3BceIWxGWWm94dFRVm7XrwI6Ce8i1BW87
d77VBeoLYC0Rob1RwebtWgx8SwbVdzTMoRIfnnHHN3OufGVg0NOXfof+1Vtt+WBCtY0WP0rnQrJS
l0lBRuAEGUsHXzmMOUxm9d2Nh9Baz+upkHE4JCwgbjHb6v9107aRXOxvac7EbA9To3oo7tX6UDoR
X76dnpVc6C1XQlnT+ca1NJrpLlTMk9ylE+K5wTrlkgdo8mv4v0RPvQ/AgIXqgpjUQr5Tql83zNlB
9AObB3GiQcSbfMjZQGZs61ru78HLWt4xLiCrN7uciRIaC2S9Z2vq5DAo3dugGtG9MKXd4v4Kjw+8
0j2icVVv7BJiESfWqyI6EabVqtYfkUnl2sEZVOPzgAWQPr+kk7nWiQEel/cSVmoGsxcYtSRAfm0W
YMlXUtgoFlx4GuT21E1KPOU6WbRQVZKI1lr1mQ5YiEHN/WdfGSNmqR6QbGZfwia+fdOmxscHBahf
vK0aF+uk96GJ3KS7LLI+hB/ZbqQBdQtlbaEkM6wmOCIROXTXtP2L6G8QLANLIJzey7DEXLDGs9W/
3uM12gT9aEY1Hzfj9M6d3bddKV7e7ZwIHLMGfLVBwplXVZGYCIwvJMjwQqdDVB65iZXMKya5jic9
8T8iQceW0XX48LH1k6gvdSxyFW2h1G6XsQ5iDMc6/1OJTUNZa3fzqUomRc65R9sARNHq1Ih7JHQ3
jcotZp+NV7GjgVP7qCSdVfbpkqHvFkMZ2Gf4Hoz8WVIbNhPrBqkQS0lsrSyFtzAJSdUE+nFNQq1w
s+1ANXYBsslRf+IBJ1t9aSpQqPhdUiZzIFKBrWRr6uOw7euMNsIR/745W+XUX1A3Wwjdz3BBCcwX
9lFh5SFanF05t4ySjAI2zREqFTrGIJbappGoHVIpSp5RqlS3HvSo5u/OIutdC100IcTBsI2BwpAY
Xr1lKrPzDRq7vnM15kBUlfycN6I2O2qKpgUUQgObINcwlrebheezwSn/MJy6ndk9HkoXw8iPMFFJ
tQrIy0tFHq2DNmw+4kb5G1ZWLCy+9bZZySkcCUZzIk5MbmX13RblAyfcCgttPsJgoDVGjuZpmt2b
N/rEvxisuxSbiGoqWRwErisCgOVsunTWE6xNw/btgN4FgJ1+/Gv7kiWQ9rU5YHO5GtaixGR3VHy9
Qj5xUTgGcHBMm2sgC5kREkzI/EIymzfzFa5jVYxYltn2tU+xNAvt1YNAAKU/oIt5uXjXgPXbvVE+
xQtymu+ydTYabiDE9TTFyN8bv5ANOhv5fksudkq2h7D/mKRuVWASFTGeoCO/qm8SsjDtbCAdrXGT
ojU/d2bYABEAzho84jMdIWxm2kuVW8BuzbV6I6SEEtM1IYhWlZ6gLOMlzhTAh89dX2RSwgS4zmt+
jkFVbpF2h2/yTWZ2PrNHoZCXmhWKOqrJ3QFC4FWC3T5Fj6cYTLCTG+I9B8xaALx8KtblFKCJ/7/c
EUxuQ/ozU5NbVTnIxq25JVaAnmUAX8QTN/+85a3HFBjHxFIqKj/QcNJM344vKpMKZ/LxSX2IpUY5
S1a/93j1IQDXzweU6ABbz8G3ziWGSqk3WtH5B1uLA8iUVNdgTCqvJrI3ARO4Y2X8vOdThlQQ+JNu
o+5zVPUccBf3kU+M9X2mEX/dBpaOLnFcc6OPi2Klamlsbb4HYbCWZloAdolC6frkyLsigBFeFyYa
Yo9CB/RgofoRpORoohCqAJFJ7ys3IB0ZkeQs3tat66Vavxv1F7L9w4jeBHalVymdMQ3/HboP8NxF
D+cDjBY/Pmk/stuKnAjd9t1gaVpW6+7ir1vyXpJQhJ9vBWHUYd5BTIGufwi8UpXr36UehIPbKS4m
0+AV9Zw2kwf8QU9e1LLb+MMu+GK7UTgVs7rYKTEz/eOnoFH5Ree0f1aGaT5v609GEtWAro5fBEAT
f+FjNdIGYQO5URf87uDSIM5+gBTrNbXiA1RdhxYhN879g0ERiXyiJ55wzYsaL3Ozcktggrd6cEEF
OuQ1b4qeFemkzAomUEj9KDKqN/r1ZMUtTnE55ktmrMO6GWSyuuk4gpeP9IiWJ9WUZW3+w0eNLBnD
WZiC1plfJ++fqPPyYKk75Ed3x27NLUgbi0N1i+J/Uiw5fp9s6sXyohlaE6P5K69SlQXlSsfq2h8n
gGpPYSLpiPHnMGoUCDooYq5k7Z9vbIBREPENwokfpQTgcqYB+YpRQjhcx6fjWgN4/EHXMvLSRU9B
dRqUvngdkN1ZEgTCRqWKJf7yZMfaNwms+xQZWRyiSHh7XNoKr6jKqg6Krw0toQtxQhzyJTV4oS4R
jjpvohueF9ANOUqxEY3CIl6atUCZEcjAun7BO/6+8FmW1auwwCNyldM9PNLCILi6HYy+qASTwOFj
AuQJV0mfUwV1cOrAcyZq1YnlikKK/carmxyjS+pS/Y46fl8gfQ8XTvlPGXU9NGmjxPMJGVXr7oHb
/gmI6fpRhsubBkydiuAD8nfOgDhxEZ2krflxJz1nwxf+0otgEAzJlq2cehgLnxKZJhcKa8nyRXzk
fzMSFioY9wegxUJ5htYCbN5tGwHDJtJ0j7PfLcKy0M7D14RfdWyq7KA+kaxEa6GuLFESQ85jDNhN
WOSUMUf3HFAzr9NXIYqwywsoAkqE0CVidTHzzy8ZXs6Q6JmY0PKQbsZVm6kBWrefwzmDnNVjnLY6
o47NtsFn08AepJ5qioqfk1inXPVpdrbiYSdDijPdh+OyLF0HFLnuCUyfrRzSuJCoPBEwEF3EOUTP
Ef1e2ChaCI16CCfJSXyGIq5aSh6d9WM05pUft6vPz1oZgCNsVJ+CkXmKC/K/BQYoLlMsUIbxuwVg
/NWKWetzTpz7SpBPAMXLw1UORQRlO5RiIHDRQUX5QCkXNLmIGKs6FFVxkGHZAE5h6j4+TrLtR7Iz
xgmtbaUIw9Ub7Xk9BPNZ5qp9wbKguSu3gt+ni5SvwcF+YE7suVa0aCpHlqi7/cyKJBHnILXM5a1I
6zLBKtfa9wpgrKiMMCt0vVBuanR+zQG/Zz4/7+YAolMw9H2ZZaniiAvwM75dR4oz620BLXKgyMnd
nBTSRJjDIt8n30P+wCW7a81x9TfjGALaSAI2LhI35j/ad3kEZdLR39ih7GItDgvEyGRr/tpQ9UEh
8nKMyl8pcAPVYDTYXen5AFsSalSqYP9ljoVJ/t8AbdAWv6GhN0NCKBnsBu8tKvXkj0SBDQpkc1WO
s7xNf/XMe2+m3z0WNjToy9tk6BWGV1m7kw4b53bWOKFyAXpj/EnF075edGpd+AjOqLQmkIz+LVtj
9XkakEXLmqtfmgZAFHhcDqEwMg3V+rzoj5WxZRjMWmVFZB7tYsverWSMRWRc0+opOOHeqE+Ehe2n
0yWmkyFQOmP0SSAtWQDgn7laoBaTTueMrquJ54MC7eLDNdReBMd+AJXmEzLZvnzimP6wYP13dwcO
8xgjofpG0feznaYXXF7GGhFYzISZTi+mC6BIIM+mO96OwKJVyzeBkJ/bLwu3SLFaSfTBMEs9jgKf
H1kFXz+alUfVIR9YMDV3ICjlczXm45ZCMT6Pfn0wHugpJRu77Dtgz6xebwrfMg6ooVHf7yPolIvZ
3VqZXFVSo5XiiEf/3GHstHf1Y9e8A9NsNkL3f++rNEDgVS0cCXcAWlmx5p1AvLl64XxPk5ywzWvz
R/H+EVCFvH6OstQMSYfxpJElVp+4icx+zfb7B7xO8uy+NplXGUkQV4PMI48Xh2eaymby4abCHipS
km3vZFM7JLUwUDvWTw/iig6OFIfBQSY/GBl10US3pk6/HUTjrRMWhOhhGmap+1ZB8/zTyyqJuKxx
7xEJbXmOVPAU4+SDSUrfmyCZTUWpQBwwp66UgkiQONDmqC+J3K9N4qoqhoDivMJVZlAeprj1+hxn
GLWNuuk+IrONpXs4BmkXq5Xkbb2LVxUrPQ85usWTApNkd3Uil52PxFHi3TQGNNH8mYKGxbZzFk7b
m59iKB1wWMYaFIPU2H7+wz2jxwcClcI6ix9qXGgJ1jiTrr6awP3+KNPxOKYJfdXUvqqt55nRh6rO
VGHU+ARUsxThWf09fLpUbRLUgJOKcI3K43hunH2frbacL7YOYrrzLl4U/bgXQDOjM2/fO2FalsP5
F0BwDM/xgjFe2pjJurHI1gtYGgAxelhkqbgDKIGZ3SX7QLdBnmMNsGaBLF+xIdMEgBovk/mozcy/
t2cfVkj/mKe2ORq1+oXbF2qy/DgbRiAquZkwYSULCAZvX/eWTDLDb/l7gLatZNIqDqZmcAqCFqCR
bZLrR6zGSPCoYuQYhS1COoJazEY9AdBzkMWDrxzhQYgMhUtcSiWscqWir+1Aqc2QU0v7ASbLtl5e
hvY3CtZ/9uXy1lVltSC+pm4YmlEw9XpARqW6XJeGIyPbzfTQv/JZ1fe+aPhYB1+7zUscCYKeRsog
84ABNJymT3mbavhYsOYBBsWN0VDNCvdGnD5dnxR73aRnl5u771KWj2Nez9Iujn3Mp0gzaDOwXzqt
VBTNZn5keEDCnFuBQaYM98FJCOzeNYUKPd+uet3YD+MVw8yyg4xMG4SZKJtTflWOXcyDKjAdoH+X
7Qz4s92U95mMtVqplto16DFNGZuG9DKXq9JiBuMi+NsMn6EwWRgxjZ9BVSY1IPy1N72LQkvWGYLn
nFGonZzSy4xOVXRuo4m35S/ibvUXul+Y8KLtqXjIwNvZ0qzrf9h51sI0jUK8th9mev/0qieJQUQg
hG8EcBWY/V1gGeB3cpcY6VF+7gkLNOQRK++UxDM6w3OrMqO/0z0S4wSGn3X9eBWw15WIQY29hy4g
6gEI35j+4QpoAuG+/4rYISXBdrc+Ibou6SZ4YqloLKTFgIXfaE5JOvst2aoY5JDt21IhW/O/Aa22
vz7aERD9UFHBLQoww7GEN4YJHsYuYnnFd5PwdRPvoB+mpZdDpPQjTztYu4bgqGoNHAIKKWf041PT
XG+yLFy7O4BxUe3GEUSLuWlxXEvlYZd9UWMP3vHBKanbbPN8RjY+eQSmh+iY+uUi6Hw52fgIOYCN
j59OatWQ41fyad8yuCkMPj2RmtridFHt6ig5wVqzJlIbcvLijw08/S2nKbGJGDyRLf0DQrTStyWN
msEAtcWUR8NS3HEa8182Awjc7kjUqdBMEItOvCW1Bgsl+s3IRDLFQdwl/JzJgMV9t+DzuHe0L6T1
sWZgubgd4XFKLxgPo+eb/Sj3nVWj5JKCJ6toUgIaBqfnbcXQ5OOLDuhnpQq4ii1hNLL37XGUQHnG
9u/aMACrWpNe0qTeW6FDGfgNv1S9TeIifTFz3crChXsVlM5FBCts3MmOh6wuvIEFx7aZ2R0pU+Vy
PIwchBMjmvgIXDsQ9UvB2Za+brmX3jkx32m7Jsn+eq3UC07bmimVWzYNjJUWv2AVwP50L+p0jGxj
5YBOBFofY0bQ6Eeq3WKYMWmX/W8ZG9Ku5JcMrb2SkkjvJI4gAZhI6hVtIv+OZZG6AMwyPgQcwo2a
mlDpB3KjlZkYMJVIrYNHDAqFjYBqSWWFg/92txHM8tNh5OVKfMGk34SUJcEVtKbuNbz6BA/ums+W
mMJGI5hBxM4dhx0ah+XXYSAySYBwgMK6dJw4fll68d6XGW2o/S69sLjQzQLHvgsXncQ332j3EggF
o0cQTOBgDlyqE7ZF2xTAp1SUJQTkdqnzzElFxo4DT/XsZML3EYeHRgSJ3qKqcfO84D6yat3jbF1a
FLqdK4zn4Uz1/LFjCZ6hSWr5nyPKPHM7TnAJeFGpNURAbt6z0QyOmQpMQWNxpfMB0dSbRp/K+BST
uIE5r3kXKg+QFAoACav2y0Fm17E2mZ5mqC7c77eh6Iw4o++gD/JIdRGr/3JocO8h40QTDKf1Mg/I
FEPrlMYFsJnbCuxZszJ8RBm3YLMW3RSf41vZ+GDt6gNVcjY4zJ6q+r0IgpM3GUfk1GuKxvNznXpC
R8Yvedh97OFLS7KzEvNSnCNXW7d4j2hVDfKR/LoSMHapJ4U9wK/UYFNAzatT2l8Ayjw3x3YOocm/
plWEN91akCNkBoEHej6dfi+h2qa0P3CRd1/Ds/e8QdT5SRM9+CQLQX2ajWvTRM+P0aTU2ewmcdcA
WM9snVzsLOyu4lMJS/9YZpu4gu+3t8HAXJj/uImdNy/Cf8V/IlqtkOQDbsMVtVrAVjX3kMFZpMtw
A2Kx4oAdxWm7dfyOkzjWCTxBaxVyCHBuw6cUfiwnEBdevEWMMnCpsqFZG+vXkKzX5TL2XJ2vKQNs
ONtTWszqOCTKCc2IBba3y4eOBHKyWNs5lwJKgsuvHMgL0cIF4wu/++3k8tYUqwWc9huN4lZkf/vv
gdjNiDfvbvdRSppXltGc4ViBZy2/cJ5Att5fZHMVX/q+FCOLI0bkLcvINdIREnGGZ4YzqDGZO10U
NKOr3QB11O/PcJeT7KgFzMtXm0KP8ynPLlZD5FCGLVnUwbapq1gDqe5A8VrkJkC7uHp2qtm3HYY0
tSoDc+kwP9eyTD5MVRdEKvSJmdU0iaInvZJ45yUHsX/zlFVGesC+Qhaw7fBx2mJhdyneD3l3COB3
NLIaxRkNMFe2yW179Sqlbk2Gb+WN/leXcCy7v2XjvWbgSBoOz3jDHk/3aLU0UJ4pXtlu0XtZH54+
j1WlKWYPbP0IegAnS7ggg1V2Yn5aENRBPrI5YIbzMXTfCL1KHL1Qq4vx/TotcXw46ypJ1yY1Ucm3
NPrgNRKjeV3Qh2odnHlz9gCSkuuMtQbVe44g0gxaTzegTuHMTlT1aDngcEpFNrLf6k8uxYHtTxsn
Tntemuz7IgqRxrHGchncoHyTFzGtgLmf9FQgziwZqo4jYoQpnNSLYfu38cYZIJlzXNmTzbL4tVLR
4kHQpUGezJkMzjd0vCIx/2NK0cbbaFi1hmAk9MKCLliA7ujSFn0hl4HXvNmFfgmBCgljEWFS0CjZ
xRQNiQm3lzxgRvaiyfCNvLFALvH9SHqi7TF0VW89q69xSPTfkZsa2agr1r2jVldEXpCM3Oz4pG9n
46quubHkzrqZUXG8kHbEp8V0PV/2c1tirnSP/8ctdHfaMjcg9P/J4caapeMTmzZJZgfahFi5czJ6
Z/ZBfOOQecY/LddEQrwTGXiWZhuNUhkDm1q4omBbOsfV4b/QYAPeWF8wXSxIYJaaM/VNOEsDcsOW
wvpwIQP2CdOcD8vuLUC+EegJ0AsSRKZ44Bmioc9pkF6OHrk40OxjfA/35KFjTrRUnLNQIotbI84P
tEvZpcWQC+Wbrjt5mpM9O/dObCBgRPcBzQIAgBIl7uVAHp/5BaVHiuUW85jUPJK3bLzTFo3roDIx
7lIpICGjiTPKS1qQbeLHwfMUEb/7DBEQvt+C7j6i2pOBPlgOvyhNm0BEz0GboOoR0wAARGAL1LjE
TprVPm7NV7pQuAoQINym4yPLWW6TBrJzkU7oZXAlmyMoH+swOLOgXbKuogOapYhE+e+UZWaNUP+G
6bd5w7jhQpE9K/hPqN484VX3feBdnbLu5dl7vxMTaNvVdwNlRAY/8+EPD4NZLi63GKMYoE/PnhUv
r8nWsw6say+xxbpbZDpgakEU/HWmd/S/cnNGhzW+27LzsHNlRSKz0xE15a45i+jbupkRUKKI9DWq
wvMtvmHHnFWh7DjeE4jnHKEfXD4Hzf0f83eNm0wrCfa8ngbndxcBkJlx9TZ2NeFvwdUUgvmKn6yh
mTur+qtBfGK7KFLSb3vI1QGwOTBMM1blUD5pnuUCxMUCS1LTjS6NGo2J7kC6HZF3MXUdpE9pTs9y
YJ8G7Gr55DirtIpamEjAKPWjBJXBgVrUNKHAG19Z3hR4K6MXDrAhTJ8phbvmVBNrmYZ2MRnUjSRH
+fWftpV0oTJZBf75nZ2R3ykHfrDXQL9PZMYGzzCrTFRmahaYpY7nNWo22QLNMGFFT4zgY5wn8+sW
ECeq5wEPZHyc6/Z2hUSsKswO87Qb9njcF/d2mNJDnkbz32NBQix19mfSsvoVimx3Z+ERwX+XqsBG
xB3eNriQaxcebOHJOLg/EzC5O0NhsAe0QKr1PWjlhYjeVBo4w5l6QBKttPaU5Rx3MVtAAwC4f9Pt
x1cgiAQjTs3unVqi78cb4Lr4b49NHrcwarJd5O8fPi7n2DfHzxjZvAYjAFoq/iR/J4VkvBK0i4rq
hEoswULXkaEMb6k/cwUbNExKW/00hH6TH0ySpNfmdT33Tp7ve0UVAAB0XQRLE7EUiu1YKQwD8oPd
UuiYbi/5hDoK13UfH0srn4hbo2kqgJt1uTBnj32J0ilPugBFTS87fpskhYYJBb4/DxYjcEcYcGzi
VSfrQceEowWOMobCapo+AnRjy7I+hvi/aozUHx1YS6i+pC+Cu9ohwuNqrIP5yiUTh1Ku2U57WkM/
ROL65GPly+ioZFV4koy8lZU0XbV8zzbiJCBqooETT7vDi8uP35RZSNiOD8ySPrfAltr6m9B9AOlV
C0r3KzLB7G199LdDc5rAp0U3O7aMOZGbwY8vtb2fNvSbbdVeZqL9Z27T/NG5IgHJkii/AdQJB9fO
wHNj2Cl7lLKDqc2PcpkKTf+rxeerScYScO/oP4lM7zYHDrzdykNZY6paL4TyiAVFK7LJ7diRqHNr
bHtlVHc23KhmWIULsDxqu4dZosLo9PUhm+WQ8ovEkche/w6bH0OrGNu1nE+XlkyZAxHOEOZ7Li7z
rwSkapbO5vy2Sc04sD9uEojh11xoH1u6UK1hZzXifBmKHBQ2No8y0uxnhPnQ7QiDmUCz/TUwWcNq
U/Bml0VIAunBK+6e3o4xsUucp5pJ3gGcNH2jmXcmfw79xb3uYfIjiA74gg9KCPF/1l9XIjnTNV/u
O5yg/2miEvWapazHq2WacvadYFXcSo098U3WZX8F/q8l1ncLbs074tyGquAu7BfJ7RuETQR0kqh9
wYio0fN9BVch2lbrFJ9BFk3gpB/tFfzV2XMxCoZYKTnJMIl2yvS0WOCqwmVp3NNqdAPnk/zsjBEp
+T578fnJNwUUOwmoVttli2ATWSaSE0EJbXIsw3rbnII9+ferpidlNID5zOypASAxMhzvM20lVAFi
UPZ7VabJTaFrgMzLHoaq593zNM+rPGW1c3Az1yBqfxhrq6cvrFD0huc/scHwpBX5WCdgASEvqZ5p
hIuJz8SMJFJSeYvYbrWWF9EEYxxUiYjO0qpoZ0qqxrzz4kZbMa5sZUpRapR3HNbj3oeRCgfeSE1P
SpjNal/4kibilPV7fp/MDNBDQVk7/MfiQUSx+8J067qsMUj+QkqEdQnXIsic/LiSbC8acmKwgRxJ
QGoWXSOqUXaCUKZ1oGCpaeJEt4g3A0H52A6xgt7FlcF2CnQkECV4N3gos7r8Hd7lWiVibFvv3W7S
jC8sSbtPAtA36rIJg1mRIg21zNhI048xOwQz04NBWhJnm1A3mKACfQlokk/GSXNO5DYkJUtdB9Kv
UDTq5/wHLM2FsP62YUsdbjl4j4jrQNQT7qxnY2OZkc4SrjWyPypgc/JnGwO49ni3ULmINp79KdRV
YncwfzEGCgq9igs2oKRM5ivWeNDf2cEXxEhCeH6za2wwVLwwngnHIGYWU/oGmSIRBMroZx8B5yRE
51HHRZ4iUIADUNbDp/ZrRIY/aRmplOFNg5cynpNCANT2WLTN7DPa/AmEtzyk/ApR1zamP2+dAV/Y
ccn2bVqSJRp3FUHULvRmncD429iUtgEJyQ9TWTcFNFzKyFks6iE5SALYMUKW539Zkf9ucMW9BFEI
Hw8aUlUJViZJLWj6vPjItlUNIbgvl6tOEiwO03hFGYjh07xPG+0VXTiszUSSZjLYbE0c62+opjNL
eFtAtltvZTNJb1bR2XBr1+pSH/SM9TNmvS0ruNihzD27QfkORubZLkdzlrnhOFEW61vddXiNIBP1
EBb13SmNBkL4S791qYWxouXZN4byyfSXa74t5mHEshm/4KeiNa83SOqRYsAqaORdeeii0ph8XUIL
3mN51w45WsDrYQXp/eD89zrm91b/YOv9pi7+RZHSGR3Oz4nT0Q0PbfPRSsq+8FyTk6bPtQmgSyKO
zW1PWao+iREWkQMXKOjZmwcO7y2EoVgxuyX3beVaHGjiv/V9STgwbn6KBQIa0asNjliAbAMyrQrQ
lwbUbgIj4XsJUAMxW3AFZ8aAOGYACR23Utr/nbxUgo5odDXyaWXStCRbJWBU75UqwSFuyWSWxtOx
yu6gjEU3Rc3uAdTd4ZI79kstLn3HSmrwBq2ttN/eBgsD3kVgWvNW+zS0VnIdv65ak8rnsjvlrajG
Q199umbjYXIFTV4TV/W0h02U6gRWVmhbTUFPmjRu5n3V770+fg++MQFmlZVzMLVhcFPdja4S8RHc
7Gzc4jHP75i77xwTjUrTI9p9TI67JKERY4TMqwTzE7NeLiBwJnjeKXrR6wrm7wDZVh9xUqI6kgeo
4qeKaZf9DhUz53/gVH+waFb4frTUrshGACWK02OHAoXSzgLB979JJNbrWKUm8x0EQ63o1OO6FE/A
674c0/BGWol0b/cfKAV14O3k6UMC8tsx6aieRKcWv3i0Q7p3umROD67JU1ft2rN6qzqF5qsItlhS
V4xZqjS8bsMhUCUXlIbZ9mQlCl/MDob4grn4js2dW3bRt7ItNheMBoIK2gxxoAtws+Af7Eqd1ezC
KZz87FZtwLtai1bqCsYGPBi9kOMF0O81HayL/ZgBG/6EJSdxqO3UEMqF8B6dWLXk0TdmX1T8QJKs
GFW6SDKUodKns/7AqP8WOOemi6YZy/5Wyn1LTa+qNr7Tm4bMsAMtHPaN1KURnWws0SHvUu4JipyH
9QjAkKGaAQN7e/mPY11EjaIASKdHJZ8KZHxdaeZlWuudOM7WMkCpmVpaS3cskCgYFPVeam2IZxNU
ga+RZiDB0q5S4e9FzSh5KK5xwHiSw/50kZRbzWw8oS143ve+tPQfrAYVsw3rALboSPxrFdhDfWtM
NJyefiYpgQQ8cgMqE7oBD+wnFFyYhwOwz97a1Nqn1jOemY6Ew6jPJKKoTRjiCgrbMaa3QZQE+1tq
5mjPymjF/M/+iTjSotiCBGxd8ziKoXOEFm1PbNn89oTudYCT9K2dQfw/oAPkZGw3XJuGcbCt0oN7
t+zET0f0kWiLWFCTMX+5BE4rTFq1WnoQEucrFDlIAuJHh8ygv/Wwm1t3DDd3MyLXUEt4GpxIqC8s
GKkd6KDPhnh182mfhsuc7oxkMJNjnAhYKPPy0LxyBt3EJHowH+LeCLyUpY55EgfchRVWgDtW11m1
uyz5h5MuPG5AS/hhn/p/wGj5yfDI7KH7ifCJ7zb9+RXKvLZ+tl075ynrJxEAVpMGCD+1O10ROxCV
1nNXspk+9FYOnMIATxDx580yNsFwboNTEP5KlOG7cYlKlA2zUyBWXEEg3V7kmJ1iVC31WpTearsj
oOy6jd831jUHvvYJlXz65JWTa3OWThSX/RRHS1J6n5Ql7V57b1/AdR731Q4PW8w9AUUsODSQCaXA
JUx+QZab1UWOEeRZjD2I4uzh+BV2n7NSEtQiD7U2wiV2jZQbZ4b6gSUMGFi5Sey1GftUCrjoe3Xb
RWEtqXXqk5Ug/nfLN3tRYyUszdDs18NVlFKSP4co8KUzqm4rGidrW0IDu+/SjDtKpzTX8W/U+cVw
NkXIzdMzt27tV7OcpVNA6BxpXBoSD63uTjaANoOFNerJB2Eh8JkzJicXdf2hTQF40ubxICx63GOv
eQ1dl6VZzpR7JMLWvobrCwITLzJ1vABrMkilgJOZlDf9c9cAPIWSLWyNGj/Xp1vXBM8utcFuFt15
4qYdYbFAyM93Mc5VO4aNgjKg0viZLO2KXT9sIZ6REDAmbpCUTUuLGyBbggKkNix4eQTSealECSQE
qMgl+X9Zj8XkLwKyPx3SH+3lQvwwghAIwzXeEadYXJL37iKCardi+tMa85ED52m7O7zVSU82BSN1
wj9s4/Zh5d4PMPyrcrWGm3CnpQVtRcc5xKQWBCKZvDdx2GWPsjFgxICO59dSeOo0pFX75CNgov6I
Lziev5B5FxuyChXHcrD+WqTlzBkYnkBCaMpXUOUyoRFRCW4O4zQAUGcwIiAnrN8mUnMyGLsJqzBo
kvAuk/TKy0WVs0+7ILjdHkJaocjPXszWIuCSzHUiXOiL5OW6/Ry1sHP5e5DUXZ2AgMQ9ZsKd8+ji
42YCD9sGnxCV66TmXvuVdJRHLhhunkdchSv/yeGHvvMEVsDw9k0Mzzmc0BOC+PsgSonCoqr+8rJ0
jFoCucIFGVICtrSS57JCMzqdFkJNcq8KC6qp+n492rbKaasRsaqsRVRc4l+rIgIdMIYjTZ8XXPJj
pNrvOPbZDALvQhxvSh/XWHbwRsuMfW9zi+6h9XRkS9dYPq6D54QyMv3RlaiaIAVLRrysdKnV4c7t
U8gOF98xOL8bNz+beY48lbEr7iRCaHl4zMn0985UyUQgt+AGX39pWoXRdwtucPbXOBi8MnQnHSZY
nXIOHh22iioA+olQDI6z4Tqpiu0mSwPZtlR4cXdE1izj4LQ3NbypQgvWXvKHhrXjA9+StNujn7Iv
kLgbH34wpwqiK2xdRw+bIdFW+q6wPU/UOMUdvGm9YMJYwsmxXFAvvQHtzaBGUA+brQxq+1jhIK4a
5uoD5tWKbJuwgVKOkMdYoe0DDPdXVb2VaUZDe9ABKSMITtYk/mWcUYHDi3wLzIMjxdZ9gni71Eap
g5PT+HrNsJCP8ElitjqUcDnK/vCPrYW/VJdm3wIrDS/N+h7bhoI8Tnniiyx0idcwYRT6VK35bdGE
y6SCHKTCRR9z11gM6GkGgU953/UlZL0oX1DX0PfjEuNv9CIFDT6CfQuoY4VOJdDMs756AKwuPaRS
/oyML7Qv36UHPiX81Z6VY75oxAJtqG1mSZhT3VrYtYW8RJO1a1GnCk32kvrDIwBS0OUVQf9f4pEG
0fOkUyf3eUIMv60xXL5epwL3uC6EvS1D4eBr0qE9Lm7hZxWn+gkorbkXX/5RBQVplvSDc1xqGEIl
9LiBaienBzVTIuDGCCs9uGgy4Mg4cf5xWnMUsLt36WJ5EooXoy5VOFeK5uKabh1iptxrsnd3qALL
H4aY5wdCCWrhlYYGMyG+Suh5h6jILGDvRhrRK1Fcb1spf72qqwEkRaveAkjM00imYjX0g9rYLIiP
0Fj1WeBKkXOtM6ohvem4xfEYQXR1x7PTCsi3N6BCbDna6O4D1fXQ1JamctzCYSY5QZUdOP7Zio01
qurVEnHbPo7ZZZ0RsMHa9KhDjC4EGAgUZO9qVKlfPTbnXlvp51l2hJqAdzAfWIhWgbxyDdZ12J/C
ipLEwlblaJkGKy+raNUZq5XAHqid1libiZeY4xP0VFFOUX/j6hRtaN28ke/ugaf5831dxmUmVVqa
y3KkikTBgirkKuQmn13S6xHhkMe4lmgKJUCTxwiYeDgb7iajbh0KyxMoL1bB3did8tLtYSv/qfSj
RZciGbIiPZ6Y7IA2C2KEnlkNxD0yzShezVC0t8t3bNle2203t6Tm7pOHhyVSFDel52LWKsMYothF
0nD5JYroGeS3E531m6K5+kdV8h0ow0i0V08R1JLtq8F+6JOkh66MNMYcyf2vC+s3Sv2tiS5yGaWw
Hkncte7TDVGm+BQMc6AVhdtK7bee2nxj3coqmQJZJXEjM4dXpiR6i3/xd8TkOIieK5bgSP0oU7iA
4v0Ka91XJ5BkNBEPcInncYvd5So5i5SaA2FH5nS7LnaOemBWTZMNSCiEFCJX6ARvLH0CHJfhJN5g
PDuY9UQuiAw0rEp6wRIIJ7zRw0alItxQ7o7F2IufXxKHv12JYimLFV9c+k1rdjNyHW92gm5E3vSX
8Dnz8bNZoadxEf9NSQkHR9vEGjmcN7pD4D6ufwB3CC6Fg7Qv4Kd7MQdx3mwMtd39YhDDp/UWOPYo
8nF5cbH0i25gmC6HzwOUiAA3mrKno/k71Ec63qG4k0gWqP3fuy3DUyByc/rByx+kSyRtOqJT7Pwc
WcrDhE1CSfHYiu9e2tp+LFdi3NT20eSkw3/0HAwou9W3fLksxdYf4N7KcZIBFwpWsyyFukTvw+hL
Nc7oljcgSuDm04y0IUpT+PLRoQq1WjkQFxbq+0s78w4hwrHiDfXlqRpZhGWt4sefpUrseB+yBHx+
SQiN5XCLrWS30B3v6Arwc9egT9N7wZyWhp/n07r4cGdSOdaWkIeQaehen6lFhcgK5swJDza6iEFO
uZnRd+mS/jkx4EsMXkZ5rZGa3e6fqNhvSytQMaPKUDXE/gwbhB0Dx8mHhJPIEzdkCehZ0iaax+wA
kH6g+FLYCBZSBoAGauuDO645Nkz+3DbMrixhGd420ch2tCSCcLapJ4DPYkY5zukT9P8rqfvC92Iq
g4MDC34aBiduFGEmw5NHyAMku59kyjoP82lUgsFW7yfD5+8mXcH77uv8K7HPMrUPQc/hxEfa2RlJ
JvVVD3yVwFJ7NGcuNkTJZs2d9PojKY8s27luJJYbidl4zxzD70K1CJmet4nWzFoIe2d8F662XJtu
3Q3eRwDApP3RTo6Yx2GmVec5xWTBSoMekehd4D4cdzWGaoyhXkrc6GbCZnRQxJi7v3M4EsbtsG+O
45oOvh25D0qpfETBjBlM0ge9C9JtEWR2auFwKvDsk7FwpKsxeTTwyiDNPoZoxX42zaZiazyGKUf/
nM791gaJgDCz1Uv3h1hhuqCZE4unnhY5j4CSLPnaGBVYHAH753RL8XXkNdHTgdaBANz/9LYuV8V9
NrSdwTxhwZjwNV2NBOa1n4clLhgIlCRVtVORicHPoD2tRV08BV/b5I00KxPqaA5idcY2kwXQVmdP
+lq2LXNHI9wFTQhG/j4gs5NEYuSut7jOA25/JBuVsJ1+8PWMK3mUWUlMDvrdXYcyPOeTCkdSS2iS
/SfGBYJdPq5If75c0vvzVpop2DITXjGxFUgd3HLMTw/WrVWvezcb/inWTKLxAqQmrhQnrCwXLWpi
68tnHforOkuLbg8ny8cZxU7mLVeuxIZbS7iVrWvLbfg3yO5+vBn+hvXUR5zNH4J0DTrJOaD9Aakf
2nS6Nj4dD0O+PumiyFcIxtbFrG6YQQFhygOIBPk/FsXTaOu2Lr4ADzdsyKWTXVA/40diwp5nSy9E
yNzZ+lwotk4f75N6Sl6nOk2rQJkdXlliwXDUPC+9cnLi+W6dLIM15z/1Tbai6bIQ8xhn4Ef1gc1x
LL7LIyN7ajWJGW90KfGXxjO1pPgGThz8DWHQ4LiAfWxudsdwSs/GoC+Uf3yrPs1R92JrsGvqoDAO
MWmkIlb000XMUEO0cCBj8cnsnqB/eHbu90zne2q3nrDkMEhZRkehxjgJpexW2gPCXmarotP6cR0m
a5SrOjndNlwfg71QAvoXUYZ16FHrFT6tf4uGf0fyA9uCcFZ3onV90eW8vLmxZaSJ2FXtxUyu+I4a
ALasRLL+gOZfuSzs7yRTXS/Dgtdci3gFvkaCKF+hzl5KUtaszS5mFrdCrywdIg2TBGT4YVjpp5Py
pOt1Wnac12yR89jxFTJxj7IjiUZd5IRlyyMs3+XEPIhWrqHz+K5sRQZKkG0+MaBKPdU9E5U4nc+t
IqPNhuCJwhI+9SviIEkMYQyC00k6yzVZtQhepremJetyL8hB6QiklMBANf7lntkA8l4ryV0rzRGb
0rgi3+V5r4tScbPNF/L0XJAMYbEkkXPDH12xAMCKrSZmkTC7IdwfS/ex5edPR4oOIkQyAKNpo6Pk
5vaCQgMly/x8wPwg1dWPmglpZIXSnqbXnZnadff5wXSo9IK2bS83J1HcSCJEpBqgDWd3dSqh0ccS
iuNF74TtYz+y2DIX5wkjD73ZCBQowI4NX7AK2t6JAlzVlI6sOi+24BHpOBIOaY1PV6Oa0nJ1bSUC
c0cHGyF/EQ9ZaXA0Efp9xwZVnEHHnQjLRYbEiDwbT9vLvj34QdrcPOIfJpoi2zwRaSE90SDovvAF
Z3L7rqMU9w7tdVwdmePFEMOo39U8lOiCl38w7IYoqPjr12fXYi3c9IsfoOSQa1u+v7aChpFETylV
rgfv7pZZq26xrNyP2LSWR+LVrmv4ENK+bbebUxaRiRBdqum0ptuyox+HCj59HSindtCI9IgZ/VFv
N2NoxwO831BHRhRTVyYSTi9o3LByeFnlQ/lZKf+uDsWHgvAL+TWGuSctLkIS4O8VGCPov57vVTfK
rmfWWBOSDr2xlMlBsSWCZHMd8LcveWhUWKe7neI72ua8DyOwXfgIYT2qAB/fmnsd7u7ptOoYZNxj
BNx+UwF2SIOCqWQurR7DGvYUI5ldf71DS5YJYg6zkyLm3QCVFEtKseudNn8yYD+dawUK3mOIGPOW
xhvh/ne/94tSdok29qywKRGdlLSwBQ4oAUNRtUBSF9WuxakeL6b7aVCgCLraywm3bZgKuj95qNZf
xHfKTyRbZGeKWqUP2e7SL9daiztGksgpHF3y5kAdlOAku9jlTpqe2BcYajteZQo5VQCK6WeMpsu4
x9UhR+rhuQZpgcuxtZrKV6hZ2x3i0TIGHDxCYpHmQjcbvN7xG9C06SV6LgOM8i/zver6xRGZJ6xc
tW7hY+TH4syh4ENoAk8oU++NS6Fxyr78CDoi04d1KlUMCzBsZ62ovyYFWTLO2j/5lyMd9TTu7U0u
/pSvEuBhTecvynGvdnvbjMBi7pt9ZQHZJC0zEQGjUaI8N3aAFYR/Ki/gMRDCYG+sbfkWeys7iOVZ
3iOFX3cr4jfAIEHlS8jy6VCj1NOPCQTNfkuhfiA6UByVEnKGUis4e0hAheLth+u+WV+GlFL8hu27
OUMy1/cSjm8dO0zeB+nrTm1MLmUNWhAec3M8H8VUr4+bUxlb/cwYm/NFJDeiOa6bLqgR9mp6u6ME
0gefu9SqUeLXeKNdev8aNcSU2CtzQcL/ulV8TJPcEKtMjJThWZ1HgJ0VAj8+sdSk+ew40Rb+rv23
dqoAhc8zoYnGn/p8HJXEHJORZp1dpmi20XYDQSIfiixrBbelTwvNWVh+zMtT9xHDtfeJ6BwcuDlz
L9hv6USiB91tOKKp2uxYMWtjMw2+lLbiOB6jc8v/M4mjbsWB1700SaGHf/zjDB+rPOklVMgopQnz
EMv3/9hPD5LLlgvlnx+DbIt9AGKttSKIRTjMXS9lH7sGg/uIsnrgL3VwFwJeSE307TEP/H+I8nel
ro7bbuqxCVsxo0+Noi7dWs40de7x/jUpNtA6tT7tRMlNeMrTiZDjzmOxkMFHDqDOjtZMkaDrgbaz
iTT66tlvM7qU6ndaRmvj1A0vY3xY5z8CyweOO0MrddPzCSR/0wAi5WZGRBaTFehM/iesfSRCTqCH
AWJ3aFtnXGuXGz38/A0r7RLD3mKZaDU5fB3/8eppABM5i38LcvBiUlZgREsHsXGatzw1LfTNz12A
PVITxecZDJsp2f62pveidGo+LGGdQO7WRpgVR5Xv97kHcR59zel6/Fh/qeRMk0Jf6GkzI07h2fWe
yuDS5TwN//bwhzfCYlWQznuPa20Pb0GCcdcbEAP4EoGB0XzkuAlCQD/I42XuC9JNtDfWoTT6ik43
FtHgtabbvqnAeMlnNFUgoAYYvU1uF8IOTYeTbSVY8p1GZLCde9hdiUHpAnVBPCrPS6cNUUyqTP3a
SxC8bRHXPRevnq5uzc2x6dQQHwR+Cto/VrTdJpTglIs9omXLPm9ceB9NZBTV0KWBQCUI4REWUHnH
FNfHIDjHfgrpfJkjlN9A9tHYxkKi5A2r9fyhkBWbxfaHPo9W2YzBFfnA2IBIhN3/B4ojcEAvizRt
0JRSBG9t9c8flXVEbeAWJjIC5CpCcliufvZbTNbd9eprr1x5imoh/HENeZJ3iMp2iDrKe+ethQr5
g5DzBlylTaNgCeIr722MIDb0g9fyTR7+Eidb/fqxDMYkGmlEzoHisgShWTJVXMxoLuZ35+bW8PeS
upeD5oyuK2Vsnh/6fXaoOabCWBOPnFH7aBs83deM0lkPsun5JLGRZU/EkRGpiESeMgCgjFLw+hz5
i8BFX7FX/EH26WQK2K27TYmag8cCSrWg46dgM7W4FYwN0mYS09WpkmWMRraAusFUWyJCci+5YRA7
Sv6TaOeQBDdF9Yes4aLmlTtTq4mN+LretJSqQPV9dXs6cOviK2KppedujeFwGezVVS1GzqsFmbzn
oLEUBOF44aguJjoGDCFq6vKICUE7XjZ7ulhLE4TWEy5/OMdLB12K5uWcJkSxVT7EHV1l7abvUvMw
fwuRQjDzcqtpvtIGv0nIORHdEL+h9rAnXXqzAEs2Wen4oPoKL9spjyFVECGwKRyVkO4mXi28Tb4z
W3y0UTyS5bPq8FID3svFyvSNtDIIiKXd4Za9dfkjGFxX0r4XWjhCrRfYJajG1QfWCxNBD3azBZGy
lVnOj7KPQvt3xYdQ1eJuhfH01Q5pju71Nn+SQSayuAge81WEboRyb06FP4RVnyriIftecFxhZgoF
mfldLWct0OU4XpmthRsVpCeYYacN/1h8JpWV6D6lkfES9evfNyhEBqXSZ3PhMK55omJXw56oRzrM
mv2rrooOQAfMefMyDlg/Schj3rISZTh7xx8R/w1vmX21av7THLl+hjDCEFYxeeJRRRbqSKeZJ/j6
npt+ldr8d6vrGxHCjpIeF1cx773FlmPv59JbhQ0x4S+pRD4cMkQaVqCOpmGRJzpyEuD1NbdTykA8
v9DXJnwfkjcqC+0sszhkfpkuhGV/+H0QeX1GpuUkIDB0R4h9Qp1Wwmm8glJE5mudJqccXPXrMkzH
q1RPd9xihdAKvON45E4oQ29Rtl49RSc0qkQmNkyI2Fn1Ta4fQHpSk/dLiJ+LkXi1XIMUGAfNCzPc
EDZLsfoX3OxZQJ2uRwIOhLp3Xd/8XwX2qPDGwCx99HsQPQMmwkrLVDBCZ3B7G0InLfcYKmXx4/Pb
5BmAUQgLNWP0imlKO/aAC+LMO452f5tu3ljPb7IZAKEqfHPUcrsO2KTphiWe5sLflARf60Oh5rer
yIbGreE8kowQn0rUdy35o+O3znMVRkefwardOQaJ5eLoz3gTN0vUDzCn72f1QZoVcig0TKv552M2
efHunTw0dz797ibv8K0+nfjXjGuZdHTpkUGlkGfs2PYoI1ByVw7+IvBPTfxjKcjqOqd4fARzmYEA
hPaxhekSVWW3Yfac84VfXjxkkAKTSTlaEjGRsZsmTRBVB6qrBuF0ptNx1n/8jPJFrgQIt43dqpU7
8CbxakHLYcd6z/BOdnTN4/jvglBtQi3xBCzECQoJAKNFDRUqRQyqEgRAaWmFinwvkTNuACwrlH1o
aF2yOWco6QC/2dvWw7I//K5ZmTmeqGQxRLrmeIFHTgGREWmP/R5h1q99tPKJ7gdo7Hj5L2uvSNb4
DcIK2iZ3OgyAa7OG5unebh0N0WESdM9Z2OmQlLNCd6rk1d7gJQH5JHdDUv125EsKdD+Mp/e/RN/S
jw2GGRNda7WmVfn9piPjmgewt6dQhYdOQUlj7s93qosSulCpGPJrSsKA3goVW0E50ZnEkhX8jyA0
c6GpNaDIUJm2ilKIuqwQNbPTK/uObkq0oxsOaFAn/ItHI3a9hdgfWO9FPdD4Sy/GFP6LnFQrVtF9
mGUkJ5KfcV+cQuzkRFrwBHooP7U3EOn1il0bja3vzJXFPDR/+FGaNijvejQy7qSR6tpDeHAZc9y6
wONcbruK8rJUq3iX9/J7OGC+Du32HWHhtsPsPE8mezTfkmokFxFbudLwlRNAasZmZ3C5S3BGfLlS
dBY/3YWzZ965TJD5DQvZVDmzjnkWEMaj3DHhDhA7ulBdoxzvhLt1Tzun4ia3KlOLGPLQPUGyHMKz
pJLENdMA962hQBd6sAGk8VUbZrzp0WNh5LAgKVjGp4r2s6iaGGlTuxDh/1jZ2c4J4kNe7aYF8Nvg
DEtEbWIGVrXsnv1Bowp9rZe8B9R1yQEmD+44pWBdXLlSD5P1KCOdma9FTb7OWgMHlZCPD8Y7i2F+
ESQ8h6a89t6W845dtfIiWmjTUFMV1CDb6HgcoX0SYpy1Iwi/Ghf2fK2jmfYj0r/YiUKuCawK5n6g
rlOKcea3NoDIEjvn8grKvLOUUbcdGfKRz2zGxFzgj6+NAvI/DFgKD+k9MornzquROo2efLarpVCw
4sq1NSHLgIturQ9DpqQMaNivQ1vptRSSYaYNi7LMz0AOW9dzKFkY0Ay720KN/CSk5DLH71LxQ0Of
34wv4gd6fmdADrxEsT+DrpDtqY1zgA5cQCO8trqCFxBa7k93FaD5EdJs0FJvBJfmJvoM7cA5LAGV
PS1fzv6/uQkT4Il914TjZzEjpMf/npza4rxgO2UPidHoL3hQP52pr8YsY5pGcxbL6uB7EW3D/Jrw
LU7fNwEAC/S3kkcfYFoY3kthN/g80D7JeH3+alY8KHP0RupIGFlL6kx0y8mcnQe+8n+KFqtvH/2Y
fjMehxXkEqOfqnuvwT0OXyI/w9MqCg3v1BS4ewTei4tGgsteipeNCeMzTdJgV8jHcoNAbB+h4QjB
ERTM6/4cpUoLm4frLPQeDhbtZGn7FOCU43m0hg25GCLvEmXTl03gM4139pd27FLqudvy5rjxfyaz
XOsCX0qvaWYxHgB1AyLYQnxXwMuAHzpY3qxtQux2DK7R6HA8gwfY8xAnYdPrwLz/orB0yc0LpMdY
8OFORIJ/NYXNHfmCbTmXiLs/np1LuyjZawa0fqyLFUeeJzVIX0bc808siEpz53NdaSFJt4zkxXjE
Nz2ofhJSdCIKWg1zICq+hTpZNp0cm5uBtqwrUxc1Fm7oXIJFR9xzNxmrOmd4Z1i9zHXuT1PoKRAl
q+iIp0/drP7/0KuKURcijG2OXHn6+2nTft6npSW4OiRLA8QLo4M1Fsxck0rlhc7xQj5/CRJWVjc4
p/FMR68Fg6Mq7FBAT1ON9nYULgIKYDZwdxtz1iCtdipnwgfiKIblXEbPfnmYPWby9RS9IR/tn/e+
h2zaF1HjK+ewCULcnlMVKvcJ/SVinRKvpKT9lbeiYhCF+ZeghcnYvMI22uNjvkAsyXJ6zzGISyLw
nHD+kOLadt53xnLoXe1XF7qLDstuUba1fSuEn8MgVFtI48rBh0/zcTrMLa9Fa77sOzSbpZJgbKpS
95OPOM1YXRiUq/595g/y+HabyG4RcZFelL9Dle/QdBpvxPEGtWkz/ic7PatTyx4VA8+RjsxBkWDC
hTYWoiSFFSMWIsYTfnNykgcswn64S2J7dtCQ1qf1SNfVfdLLXznlxs8vN9CCN3p27kHoA8phHn3i
qAyQyaZH/psrDd0OfQ3K6QdNb8BB07i3OuChw7kHhh81OdLlLbALdrUeETicz+YEX7HnJDgKGpQn
4U1Zy0L7N4SaHJwnVfF3TTYoU51xxzyoJx8JBE4i8o7KTk/YyrrPnLDSg46BswxwXJUtHRt+cErp
PdbU+mXIOhOkfgIxxyd54ugoGLXs79tMHZrSAVVGwTKwc9a54XBzTPha5eG2C8fnF1SuMeOM2tsp
G5hSr5eTt91MdYJzGV6PZ0K+k6Lhv/mvx9TGYu5eONn89PcCPWyhyVblcxlDuUww9DvgdO1G2hjB
fUWMoIjgwYEnX8I5tpQOSUc0XML/NURTOsjDxzXbNP6b1Qbi1mewTHUnwCS/hvhYetEpEORRQB9u
qZYdhK9T20KNtTtq3mKRY3yYD3BU2zLP/zsCg80ZVC2rQM4q+7GVCxJUL9q/KR3g0q4q4jOHM7/T
x1BD1PBM5/crA7FZMCMuOlnwa4o2Y7QVE2cmxiboy2tg8fvdbVEzYVsD4q4+Fm1f3myrpy62Wq4D
hLPYeQraCQ+J3voLulOc1xWGlxdFuQLUf3JPFv0d//sXa7G+2flCLWWEsT508b1Oe6T927KPMG2Z
Ut2RcI0nHWE9yjCAe4aou32fDS1vo4fPZ3I2WyTTatLnUkvadn2J158rdqsd5Zc8yeKjURpmEC8N
sv4zfCCEsUlYZiMyhYjBdZ7Nt9EGScHgY817gi5iMO1EuZE5JHIZIbJmSDPad+qOoU9RCwrhcZKu
5MQekmBqooIHOXvS59ZwerWGOi023yZBQ3yYKRbMW6GpXoOGcD8S3KMcp1e2b9IRo6rNpIST66EB
sRPr+D/9qw+/lZz3FzKt3BklboQjwz89FiyMxAPHcjuVWjtro/8LYxolWyFpibXL+4BbVlUEMMvL
rNCfGoF59XSKuFwxmJrX+/QGbjhFhkC3srGH12TBESWqIl2pIcT22D4e5BYlDwd5QwAscNCdPist
f7nhwSk9azbFMgU78cT2EhF7SRAbuUimDR2ZCuZAPQao825PUKHq//2EH/K4nYalTk9jbtaRS5l0
hs6FkIcwpMH2LGXvvLCf6ciGJCxLUtJ0LgnBogOE4Nh9Q7VTIPN1yHJbYJDcsWDno6HRAY65imOE
R6JzHoYmnsGxQbENuC3R4Ao83ou2EJLR+Wzqdn0XT6DaUcATnEux6kT1Bd7q+IGL6YsxIvASTCry
tk1A3yaswc9b/LMqWWs+tGkgnZ++LGA0oIFVwGvqcV2VLvsPKgQGrC2wYJBaXADEV7MTXTXGHxgn
tLBeThY30W4rxiO2ZjhhjISpZPsEKZyy/GFCXTTxkc5agdVWL9BRTILdg0XIv5KMB/BRNwrzMDIn
ZbwMlEdsbkPSIzwmXZZm1F2PyKI9tBNDVIec5HhH99G716IzqBOOotEedP/5fGqfzS5RJ4pF7KdT
arR+yQgjqbx4poP4ntepPortVuj4ONqSgDQiPHctshnmW8q82jFp2O4Hb0WRFWosO0/H1IMzqCPI
njICFZXs/sOoRcJCTo8ePvG2PiIega8sheL9SDSr87Gr1W3tmNnQjXhABawRCqf/XdgR1ZxLTxQN
R1HCXfE/Yhm92P6HIhzmDTpO1gTP7O2VKNP2zCuX0Q4HTbqJ5uJkzwmaeoE/uGL4q+t+r4tT80Im
+nmjnXCH2Vn0tka0YY6JBCIsyOHYQyvejvyat7cuaHCFNkGEYPYwRG51oRe7Bz2Hg/wpSe5ZZz/8
6OVQE2vUxEdiEkyEI53SZhRYXRmOmhtP3Ue0x0o+nTmTBqJVvAZXH5WteJ6dEQZFwM86lMOuvLPn
8vYh1Xiy9gqMEq21bsQ44AirInSFLvSkbb/C8H1XorQ9tl1BriDPyXN7GTSLjVYmwynNBlr9YWZC
qHwD7+xte8ve3G7HHm2DClEuVYantEvHqHMD65PWhrd9Vs3n4mleDuCfs66lV1JuYrH53N9dgJpP
j+FIz2rE065qPc9wLh1kTgRQWOuQ3ZAoo1TrNpq2qwbjcat+BTtbIsx8uPxLAWneDjbUXmp+owmN
bwLcSf3zHYztH5Q/z4Gi064yJQUARmddqyAZ+/YqJeN38/evF/COa6TpV/UWmWfsCdWzkW0KI7O4
/YRxIS0R1zEuYIv0RWzUPkffJfVVfq4g0vpizTObGaeRFWFFAiy9zKl7mudf1tWX4plKBrhYxMS1
NXdL6JwIQ6sjNMj0eSwZq+uyDP0S1KSw0tctzCQg5avcpLeZR7PpjR6XgSe5JPrdkAjAQx/IkP1O
b9K22OyIaldzQjmWzVGvkE3KHT/30BleltVEcUcaJ8NmBaCOuFwbZZMvKF1om0CvxGcCZuTMns5c
XQr3CHdDBGUYwX0mGtC1VVZoMOl3O8Y7PbxMSoQ6vMMS+zUkFjeW5W7YfDP3J8yLDFsyQWzLdIOV
8iCG5BC2cW2DvURjuNPcVaeoE3IVUHNpaDFIpkCl1THlwII69hrvrR4quvJ6fLyQhhcyk2BICwk6
kB0/dys86frc/3SN6z/RKJp2kogZJgd+cQvka7t+5fh/CrewHMER8a7jwMeYTarrXlIvuurI/sox
hLuZt55HBaIReSmqKF8j+oKBQbv/BADX660pNWmXel9Wt7Ny1D1nXkEFMsqGON+vOFU4eXk7t0aw
JQFSESRTixq0alcy3cV2bqvhwPXBQ5FqsBG3Ytzk+YUApC5lYn/KAiqe6ftlcRI6TG9ZELNQ2aIi
CiCjiCnMyY34dc2TXo5Ispu0tJXLFdvWbGneHo2KsVgnrCdDOF3BS1UkL/akXMLHrYNpuH85dVi0
Uz3aHTK4TsIRmSy5B4PGIu9FjldPqlf40GcRSc2XstljjjKj8kgUg0uerEP5QkHdNr/oyk2vIu2I
RfOZZ0Xo5NLGOD0NIjaJJR7BSQ/kLUAoWseRVHIVH4u8teN338bMllqC8vVh++u+cwpXmGXk1VnQ
5/+pKQoBQ88VMzN86JOIeYmrXtSDG8IIvBYc879JUCM5GQOkXlWIzouaXJh/y8lGsp/dSnrk5GRH
Xce69z/AkhBNPLjIg87vrK9sRr2sWyBqdqkKgICI+fwU6ruK9qsDiT45qf14AcKmm//BXS4wY3d2
cDlvQVHpnm38LtxxXW+cRwRdvFmsyDbALSt5L3kbHLvS57ETiztTEYhJi9tjvIjMtd+wMk6pmHE5
u38aJUXVU0Uq/17TjRxhe2zhGs/Op9PFsmuT1Ffhq24EyRxC/8sd9++wIjAQZuNigIwxfpjmJU8E
G/S2W2y3kqhWmr4qKeMMyDHcZIdyPFHbEezFudnWxipNOnB4Ej4JxHi8y+8CzyQ1VAOlWd2JINzB
ZKoNQcSH9pmhoYhygSEZ8Pr94I0iNJzqoJ5e6GUDjIcbUoh8cqNlvnNaCoC49VtDaxOALkij5dpN
cxtqi/nWc9REuI6uBewtkuTbV555zOvWySxquFQEf/wYFXaoeICh4KzDI7vGf8EbMhfYZUxFCY5I
saJt2j1EdnRMQT/fyG5AAd2JcgEwE36P1YqzFUL1lAmuScMJGGmkwsidy77f+08NqP6ykjdu5jBC
L+XD+pFMzHxpwO5QaLaTuJy26Ps/qldP6ilPVYSy17kGrnPq9Spmc23CGuxm3Q0k4xTdvXZc59lJ
MjnlstPw3pw5ECsIqvesZGPjvBB/vs0grgY1c7GXygekIj9K0+rKCeaT7DTDAGaXzVQOTZsYhOME
/Rvz4b/9bZjMesgmanz4VpUiTB1uF+IZcELtJotip+rhFJbgYAsI5nCujm5QfASwXVcsxDYx1zYG
ElDHA7Y28CqRYYh9s6Ka2GPimTS+X9Yi8Bc+1JrH4bsPZeZaBTmjovzpj9zOaCjbYBoexMHES3FQ
aiw8b3PDqOuIvTZS7nG9phslqEww1fnKi68TzYmCQuX/X4lp11lbGc6nf1VT3XGmyI8X+p8xOdXb
JyeeWtazc2gldlXUuSO3N6bkeg2+WRRA2hD6EUaMV4UPWNTC6dmAL1W332FGoUPgfqh9nSc+Nn/3
5F9d8bp2fEkITtc/pE7oZEeLoiRk/YZAA9Rxg3jPrRaeIDawcFsgMvdi1xPdrFm8Xh3wz5EuUraa
U7B9xgjaI/vDUMl/aw79iJUXD3V5hHHM7v9lXYjLk6DZv2AiGlWVkpeujXs4GSdk1Cvs4cMIf+vM
EeXI6LvRwn/WeVa/Fi81emykoOufbzrRnKy7FapwiA5kpdLM1UgkMygZQwAqz23N7Aj7h66x5Jju
kRWMd21H7WRsIdkehutRLEZtuwqR2AtnzYilFsBps6cm/gpHHMMuRz88WBAm+HOi/lLF8rRLQZDT
6NmljkRV1N1PltyURW7NnnbB1Ct2NtmkrGsLgm0vhmddY2xWCHCw3gEkeYmHxzUyH3gRA1sky7gF
VR/U7dqKoLAJPdLv4d2sIXn4zLI8kg6R+RkdNmBvVv8Cfbwe/7MsMR9sgWOXsX1n/dbrYP1fZ1JK
mZWKTd71PmMNV8dd3NgPZTJ3iRgmBU3iIS1EmCTroeOaWMNi+8oDP3qCs+BAVHNnam7kxsgJ4xkE
qcMnzwXIWZLNh3TVhMasfP5tCSywBNVehFQlts9OZ63mwZ2ygc9YDN98MTUElYqAL+27xBZa1VP6
vi3VKVcgp6LO9UNDucQ3TECgxR5eJZT9avCaSckVZV+LCRgbEiHTxh8XDz+BoJKjq+mdPQzNLnmL
fW2sYeNrU5YNfe+itSKW85RmcR2kKdMsgl1W5DOHMBbsF+1RAi14l88Ap+5YmdPYSxvc59hU4Uhj
dlqXXuOmirnsYLJaIILIc3+K/OLh8bDip+sYW3+bDbVOzS2zimRP5nAzLGQLbA/MlZosKl3LdzEr
mQWiQNTOTTliKB1jxhCxJKHKeWksOzVNj6nwqexCtUn/G7NqO3RjtYRjW7N4Sb2B6+nv2Tb7bBhR
Ep5VPkfLu3XvxWIjKLSSTSOaLHEQEXNjBMmUNH14xYpTDoq5vmroK190Jrl0pmJz6KxXjXWmeshn
18+Tz4RJtlOxLD9jhtH8rSwzWhp2nRZB76FBgm1Moc4C0WErGkH+id0KPhiV42gbdpx6RaCWrvyC
TXv0Ti9wBEvfRPQFV6lCWBOHWXIVa6aGM9hOP1lzAGynlkggBt5vYYCenjPXXAb8tf04ponpoyKm
soT7iv+crRpYG8fbHuroKAC1jo6RFV/IGLNu2GJ1C0/eyc1sPVhiec2u02bH0Z91lWoIl4eQrAhT
SplvSJieVH5RDc66GQ6LRaoHRu5HeHuaUvtGaMN0D4YIWumjEraYcPPKXGeh1+vlqqI8ER/E+CNs
v0tc4ohHNjjI6E5QSp6XzVqLlpn+LVMsY4iPLony2WNAPbLCUtyWWBSYM6F0WJvVD80pXcjKsrgT
AJVqbiCuAgydsBmgi397Cw1m/r+kMicSav2qZZZlqVhsdWMOwpyvn7lNqqy7gmG7QKrzlOwv1FCP
dOGMOO/QxXWOxdsezxLTcmyWzC8G7EimH+Pi+UmqypU5vfpVIgisS5vp8TFSOXG8vF11+6Y0Gyqj
LwDxrQkIDs+3DG6o95pBXZo7pTN9ZYs6pLzQBwkxH2mH41Em8bfNSeemlhdJZ+70KLL+peVfzenp
exB1C9CsNnNgMSQb8aa5/c9K2txnvWG/RkURKqkxW+kywJRQdCe/mSplLFv1R+bfqOmv6AiXDrMT
Nv8D/cKHq7kXjSaW+INiNIeqQ0zojrbxOb6n3n0n5GjnGJeYOoIEhODSC69Rx+8/xTJvpRNu742I
/wC3ZUp+5U37FhCvXh3wPeHeTWEgQcm4YOLwbwuHzYa9VvuuOiQXVPGdTGnV2W/J/9XE78oU3gIe
iOd6oZpVskbfqSZk+kTau3q7d219ZfPt0vjhTKFm+URfL7NG+Hug7aovqL/1KQOx7BdCv1Rtl/j4
cF+a6Z4Lx/bN1Ohv+Cr8JdbE5ebNSbryGPlJ5Ibj07anz7qRLhsKipWb1WWEWNmpJwNxhP6jIgJ7
AsZAnj+OFyANMYyB74bnqOaQ7iceYP9l/6YjuFmkOkeprkjR8ccfhDEjQmxgfkmIS2gE/3MfJAyU
mhwENIGbmo/Kk0/VyL0G5XcORBUkFdC8xJb96bp29aACh9+EmKnCxCo0dXXcRb8Vzp64v8N5bB+b
pxwt2vUsdLuWRrVCiwl6Sgd+RBOpXB9rLwT9hrW6tWv2hh+/OOwfoVkF+SFLnjzD2RTqg8OXsC7A
0MknIzp4l3bvhneKM+2Xm/QrnbPzi3hkVHu2ZDR6j8a0ywZe2Ss6qdgArJYl73Er/wMknJoRoxCs
vL2XxhdC1UJifwl3Fcp5owqCpgUdCd0Cw/+QBqwyBWH4PZdyrpcmqR7v0BM1JIwFFqjxklIkm3UX
ajx3FFoxOSYZs+zbo6YxFQJAGA8pQY+UQRiGreaODRxxocKDgAloQgBFoyxgIbbI6S/6+XVLWHmL
0Az5iAF41OZg5aDr6DI/8SJKHKRQ1uNMvWDv/fg8l+VTTSGqHwkL6rMQQT8g5KEAgXAl8hbSXR3J
pt/3zi/6bYju7VXyZ/am4o8C4Mk/ZMqMeMAJTA0gpmMTtiqQVrTvoJUAZelPAFE6Ymdysu8dvDFe
BAS9v8dQEZhmOy9AD1kEiWdoQNBLZOhkVJ8I06k8ly4++XpsxtikolM61NmXbIM3v/f7piHb0cAl
Fc8rgJlbD6gqcSWs72tib4pJhQnGA5MXVVt7Bqjt+n0+MJuUhn8c0qxMkGtMAYjHjcGK4prmroLl
g+zCTELQets/yw6OgxV0FBQQQQ91BRZHcHUGqY28Ql4o2pBd4bjj/PbDM85xu7Qixhu2QK7XruLc
Nm/WKHTLjRix8VJP7HKzKhYeF2j4TN4VgmFK/uXGoDPf8bmBzlYSv9UiuhI7RGGV3EmRddxhMJLL
rBKSWW9Ojyt6hWPaUUXiQeDMxVTMoVVi/HEw7gAfFtjSAtZbzmmiEZ/w5Tt9iSEATqZK0fMXkbii
uz0duKPSn+a5py1Ade2g8vXiaFiCFuz83HlNeNH4WRfuikSWkkEuOQlUqtJaqRqaTp2O3cTfd9r/
Y1VxliBpMVglC54CcQwg41cPk1tsFA2tqDNqs3ExNfEVrdVNDIM/MqLKFiFAsaw5xs2MydS/Bg2B
NHt7zJlOqixBX0AQO7KZ3gURgZMoJX0XCvj7rI7qwRoOsXh9pkLwzIYxnx7H4WFZViavNeFTBkMP
tXm1ohC5oOYqSzhwYjkwKFwuPCrlJgh54rLd33eCVqCAupHXrtwXMVBvZR4Nw2ZopJQ3rreNFZVI
eb28h3QWZQOZz04HJ5JqQTOZu5+h/2be0BZNrtaI+9nLvGn4q+Lgq9x+kqe0Lj/Dw3qVZu2Liidw
lPT5kZVt5LK9aVx9Ga4Y8+wyz7cvSsXiX/FPY7GUoHI9Zkd/r9Nhjue0DD30sQrP48KJrdxVK5vR
nvsjGR1nf87qlAuASOEFxSqgjtvtYUSx3bU9zeBfl93vWFn7WrVReGsCHMbY6ajsJAUCjbjO+iKk
YenB/eMei3bwtWKngqug72QUIgnCvZtztdVHv+Pb4vGl9V8keygh5M7mKIjmFfkBYQ63UqnmQ+A2
nX626KrRZ24IY3HDyEE/LNSxYCYSrACSDmmSQYUA9izfhG7THNc5cyexn04dYlT5Bk/QA8zQMUf0
9s3I6tnagkGPH/rdY0Sm2cPqRzFzpX/wFqb0SRUvYVwl31m8CcJOV27RYUagtDlUQZ/DsUkQkiNp
OTxJaRFP2G3rFO7LpcmcGD8kN8gfx7qSubc/ahzu484cihob/1ETTq/xJUISm7CvZzu95IGxslkH
lp1k2UdgQIIxfvsHPH9140HB22KtXrnLxcEcqCbF+v9yNgv8Ka1S/ijlLLHkIcdPtLug2suKi+Vj
0nxjay7wmwsjc7sXssFh5WAwqpPfxNUjT8oOhRv6PhhakTa31bPahuuQtx0hUaJOF3HO/mDK9yWK
xWZCVT+tq1ohVEpBnOYWj37HspZ7vsiwtVnPQv4XtFS7HzF4yVO9YQALLSNzGhrlAkdCVfftqcUc
gmGb0jNhDPfIqfprl4N4Fk7ph1tnR7Z/3Ij9xi76KIDQRbeXLnwN40QAxSA0zw77CQnhn/+u5bfh
MPDfVSy+wFW9WxNOIKj8pCAchHrb7jfz2xEHpUIUXT0IwP0FoP+gkrpe1HC4y87BsuKqD6BhJuvv
Kz8WS1u7+WYMh4zroDn1S5B2An52oIQM6zSI/Gpp9TY5trW8jIIVPyswQjUAaMmLgkb8uaH9b5vs
PwKdOYOB2Lc6mTuUDp/HdrIEfb9bLXlP76O+B5yoZC4Ew5dxJ6Bk4CEBEVGlrK4CU2f7kwWGNcbH
c64LHs4eC0outO9LdMs62WaNfdaFWQpzErWfTYaFvQkzkDbTKvDJBJynbo/oD68BvjBt79tnV5/4
ePWIVFKhxdHR06sOKIMn4Mq7+4mnlz2ZDb8xS3dZPnEt2IQEEdqAc9TjL1BWZowzbi1ROdABNy2l
kEcpBgpuoMNyiPJc5P7HD3u3ZluJvWuLj/m39v2VVDYW1GajbEEf4FeX1MbQk7wmcJxVXutocPrR
eM3lqQYz35ieQKtBmYJmztyxUMrkjR4krOKAfgnruBwYJeg7gwoAj1EYXdK9swTqLUFtdAtqBj1J
iZnhvW+11m98wHSiNzonYb/vP6PX0HO1T7oDE7hmGCAVR4q9FPF21XFyiFzhu/9dRqQwAl44jKXs
WJxQ3HB9qBAKcBhsr4g7+kz7SyvegZgf4kW7hYn+5R3CuaLp5vHLEMYy3rEKCVWpzETGT87VAn3O
+4GnSIaR+SlxOE6lZ7QN+PoPCgBWKiG8vU+H9PJaLz3o4HuV0mMv4vwYoy2iz7bktheykh7KyurH
FHvy1mMdWzQnNgvtz/5rDrBsXh1UGZCfvatB1oxPy7bNckEalxUBR7cnzCJDKGIbBLaGHvfYwsSv
NZ5Ux/pGDqF4OmPezdFD6XpLxvQ96AyGZ02xIpHzMg5USzqI2bZf9PUBIO12nlT0DKI1S6kK0kCJ
kCzHxX5/mWYyL4xUUxunwe19qUnYRQnhHh/f2B4R7epjB3/FYqXKiuP1NF/a+0of/NCSN13/Z2e3
PVyKhAiaNrSL3/BOQHPk1d4ROCXruQiClAVSvEeGyn7dZ/Ur9pPw7Bgfn8QvPL7ljl2GAX5w+s1m
b6/0MGNSmeJJUs5ppbrqTPKa2NqlVdkKHoDJDNBX8QdWVtT+HiL17luX4A0KkCUSCJQ/o1J6sh/i
T6wab2Jb8qTPHlO7Pgu26YwdeoPQwreYHHxTtZwLmc6a/hM6/HfUUV5mC7JiWSSlkUHZ28ezikkE
7oCpeQjxr4ZzEVVXvfHultpcFUREAEo1Juf5y7B8likgf6a0vGrEw7T0weLFHInTO69qcdW3nqsd
0x5lNInoijeMobDl+aB1VNJ0n88pOyVwppDaShPD11Pj2xjDlE2rfReAEpBH1p6am0/xGv64LKcS
YM8yaKRvqR+zglLUKjE31KrZtzAYVCSzNpeznLlaDkZ06QiOOyXX7UNyP0HKHzKS5aWxHn+mp2On
w4M8s1cldIZxwYWrCRDV7BMxgBpTA8N5fTQbp6OA0xOxk00Woxp8hmE2sojc86PVcj91lxVVl4/v
Lu775+QFUSMBrmjbNW37KMIJhNnhWHj0U2MjzHAOsey4tbeZcxlJQkVI3o7SLba+INBa45zq2PC/
WIwsy/AonHTgV42KX0rO1q37iYIGHLgEgy9CHj1pWc3ygv5iQCD4EzDGyHZACuvMq2iY+O7k9J1A
b1lZovEEs/1LLaJMeNc3xxS1s9uFiuo1B6mMY5fgRMKglSlQrPs1BU1uZi4VAwJGnzV2KBHStRVD
3dhnae9mEELL/Csd2u/vivcE3MLBxNAqNVrxEJiZ7q7fzX3zhPle//emXbE+DyvCxtxF44mOhVK8
rwNJnhwVJxzJ8lxNIQU2/jVZmWWEtOrydNPhTDGmTx7AS0fQie/FA6Uj4dMDTqYr3OJY3SfWTSRS
qkDCcxWwo00biP1GQhbHcMiS37IvVmfhwHbxpj+nzOz7+1a9Il4beOXF8HslyrFKhrzWNY3p7GBo
7942uE0SebstAn8Uu5G5hLPv3aE3XLTFMxeqKKwse5QROs8yyXMUPIxhEMFUur0MkPBg66eIUcZd
8fwS1qAEenOAm/GA2Vf7GQ+O3fSdKFMgMVtGpIKDxZWnat2uZpgoxNH8JPAc1Bk+r47ngQ+RHSU7
ENBAaxMQwlcasrxRkpvwP9sCCpJ321f1JnrGf8VbtutDFNh2BvIHU/ZcEQKRTUkzb6YHQgtXLzAT
lNvfLgLZNLaJdEdkcL9/MMwehEAT5TFJIIw2EtuW5940xCw0qaefghiw6dKclMHJlzdr8QMO7QYs
SJLRE0ldtQEJbjUrsyRR9Nv8X1epTJ3kevvDFaKZ1ZcKrTkl5pkoYz/W5Ls6gZElZNS8hjADjTFW
KeRx1myqhWw59iGgF501Ummuc1yBcB0D/jxzzhoyL1UXatSReY7Iff1Qrzo0jAW3drZNp8oQ7EtD
KwB+xWbH2ognvRzEVMpmbVk3tUlC0KnCQlGtid9qBVEi0RXxqsYl/+DmzgYUebwIbEULUjUPRi/w
LWAxXS64SU1wv7u/gIr18DGKuNnlzfbLYp82h0NZ7lNQNrqKVLbFEJ3DgdR3vZ3IHfZi26Y55NjM
hIA7+zMXIoRkjEGNSL6pi5E/5eAC/GORGxSU+6HiGNINn8iWpJdQi/G3/ncFsQDowXxt6rX7dEfh
Ifrzca+SX0NUpDjShNzl4Dtxzau9wNCtDOkOU9EJLmE5Lj5dtp++k5vNQOGifWJBku6jLyHluAFu
Y8gD+7r2rxeZIjEZjTs8rVPuAKoK1X5Vgqfduj/o/UF1C5TbjBSz4fUkl79XZJP0nMvD82iG5YFM
zzVY35PXfqRqiUCDis5OjMAKl0UFvlcV2kRq4fjTzP9Mt9xCtZr9VSupLWec/q+1I6xoZb1W27EA
r41hjNz+sfx8uOblDUcaQoNMerfEah7fyXw0LIXGnXiT75NGtUz4WZewvB49D7a1VXTwiF3zA1lh
sNrnIfrmFWg+1MvHwpZr17HJzSfcjt6TTtDHl6xSDGBJlXJsxKCNGSIimkDTWOmANTg7S8VJ4Saz
OFmpKUxeNiXE6xi3zIJdG115OchiKs5jyat1c26PyoXfmulWRmVuHmbYq0H5MwM4DJknB0W3j2se
1nL+iLtsux5CmyDCCyWiEatDG4pCHRY0IoBVSz2mSmCcdgClQCBClHJesJFZmiSV47PHLYGXbzx+
dHvopVzG9ZwbpFRRphyJmUZNDpgBY62ggTO9joNwrpLkYHIK4lMtqVUhIWdjeTl+QosiHodoliTk
LHdGTXyOnBeB5SBPscGo47K/28uJjuVDFxcjYyCCrJ5m/MJekJjJ23d307UsrxFJTmRjOsptn/u5
WkS4aaPAn6fJaP72MlQp4D/o03Ux0Wv7knU4ftsE07ioBAzMzuKDc7ufPAMO0bCK3ujHqviTWBfp
Mxn96tPTZPvhhV9j2n5nm7TzdAbjQ3MFoJl5fxj6CwwqHYCDNm/JQ+PSXLptMnNpnyteV5WV2u8w
uZWPaCG9aLWxiv0cwqQ7fyb7nUIuHWYCrg/mHrlSslm8f0IjUBWR2LS6K5AD5z/wK40HvZL3+4wf
c8h7CX87+UVlccjFjjLzb4rDQ7p/Loe9yX3hdssxI88Y12U+m0wZW6tPYj1XK92C2/lNYilWbGVQ
UFPMTlZg56eoN7mmadQD5xIIgUEfghgW3ZK0gdrtqhJs7Br8yTAfv4Q2Ie11RbO1EwZKovM+IVCa
jFszFf4C8F9nGJu4Vi8gCEiMjM1a+4cirYTrvzVhgrH8G4IWXjGyXbrTrjPxWW5lJDT82O/xZ1xY
z4sW8agq9MsNZCNraqeOE7KS2Q39LxA+0xJvL0alZOLJDZTI45se6ohugKt43R9rKlOR0vxFVF5G
fwaEocAk3RR/qwYClm+oWs7PCG8fVFI+thkya+Czs/DLITCIR0QmHwS+m5G1VBdNETzFIojKIpAu
XoYATgfxeTVjoSPEwVOjFR6P0j8TXMxvIB0V0Gm0RZZbzFJRyLZWKfofG4i0f86ybH7R72gnzZc0
fQnKTHTOY+IHYVQ69FgoK2Bke5XXQUCTgL9GDEXHfDeU22jO7ircxw3zmTC74ixo+98sUJVsXOUo
Wfs4SrPVBU/HUYdUereMdIVZ7EZvntwm7uF0QNq0CUl1hqh164qAYWAjZBWmsIEJXEF3/oDfASAZ
d/smyzpC2s3/OJn3yDrzT6HSXgESN0N0qH2k2z9++YX05SQ69fPDd2fX2Xjey8iyC3n/iKMHhJIT
yFw/Ncbx87DEn8izke2BVhDWtOLN6Deiz9GBT8OybmZHs3Q5iMVP8vz3+Chy0fJR33udqpU/TRRl
SZ2RL+4GcFljZX8MSwsdsTL2oH/JGoN+wWxtoylCXAA+69Je0cC+waHOiHGzs+b+W37niaoE0d9D
7G2vIurxM+IEz0ZsNAd2eNUDyyFaJh7F9neCCWLDlEaXQhjQ1RQZ71oXRmbGJDiylopSdIcbbBWB
CeqYfpoHau1SqoyQPaGLxc+M9hsyQNCeXGuc2f2TF1XJOW9bLOz5yata21xWiFjnMXnKh3L5hxX4
JvuUpxHblwXsSnfWWgoP5oZc1rXBjKL2ps5QmZV0w2PvJg4RSrflYke0+XXSfAYKk7EIu1qbX7yR
4CPQL/iFBZKgl3N9FB/mpjbkh45vddry91sdtR1XJuIzAgyxLeA5LdZ6+mw7A9BnAROzzcIZaLqd
iSr3rac9o5EBdJyB2oHYTFCJZ5vNNSjJF8Zl2qtDavo6NyR3WWERJ+8kNV2RSCHCIrod8VD3e2p6
m42SS0/JIXV5HvS+YH/TcrghpxXp7TV5FDH/rRRqOZPXVskoz4gjrsIxpX9D10GkSsr/zRH4bxqQ
dzN85JLr6nMYzhNwMiPX9BuhwMxzhrTAF6gUAipAasosoQ1DZET0W0Uf2puHf36NswwMYzwZnEZ3
iHRUVNBH2UKHP8rWSuhHzkJDwamCkE/B2jlhmI2QINPQRtAxlai+z4uWuFpgDqmCVzDm6rpZy+XG
ZmkEW/AQ8e4KVXJFO+7ZQXSC/ffUIwKwW2B0Tm69q8qc4ZsXAVI0Yk87D9wx66hRxb1BbwS+5cH0
5rcZRtWDiqch2VGqRmBmQG75mCi8KX9Ms0B+9Ap/r4jLI94II3TYYGWGHBq8l062SRIZ9HPWV6Pe
iSmqoKTBYNHK5OBI3wKwFDe9vwpaz0bq81WONgy5S0bKtSoaDI8NEstFIJS1u/YAm+g91CoElaUj
TMJypKUh83Su3ajmXXv/kS41vL0mnpdANIZRZyDm6b5ezHxl0MT6TN+2DifAJErAsRLN2ujx0PIY
meY6W2pnUl4mnNwcuOu6KJp1g60OT53mk0ngIl93ZwIoXsBHRgrq5z3ftBAf0YKl1LrrR4KlDvkx
YfNoZeHRkDk1oy6hQ0Uk4hCq8XCXgmk6z0MbvAiPvaary4DH4PEYAX6n9+zebTDvYQEq+TAvlt+T
VXu8E8B0pOUSa1WOc4oBAUAcBv9CnQmPoH2kFcS2u5I2abZIJL+nv25RBmAIvkpQbmntQPS9LFt/
3SX92lZ7CTKUabb8O7qtso7Z4gS3Y67PY/lVP6w0LZe2UindDd4uO6j9cG6R5D1r+mc/iGk+y7pK
cGn78BaQ9C7Dsmq8wwCSG9VyopluES0bVk2RoWlYp6jLQ9BbsdMymweibQSuTF05USsNlPjtPiUA
rxhpVaz4o8dmuJr67GuxI8ajE7XyWtZJ27m9tJpiDu22pRz7stO1hHDZYcr2HmoOFj8fT6/2j6SS
f73qJ8iBdQTlEpaoBtcRUQMc7XdgJaAeyCjHimMEfZF3aqZMN2fZuCSftsy3vako+7h65LbQl0sN
ylhsZ4sxuFFZ2Zmua6yMpZbA1XsSwrR8GHK09BYkEsi6w8onwlTNSexqIsPXKuahkXt3jA/V0VUV
fpPzB+EaWElkeW0udJFQONGp+t6tqncKHkLyDlToRw+XHzUn85trk9EHcL5CggcjuNXmq2z3RPlk
2JZdBsbCKQtNVHHXFZ32JhtaZPByXQhSV7IpXbsryDsAorI5pcnSL9UJj5xBicL+lNVOW54EPxnt
8YQOzdFFbpMW4FuCED2rraa6irzn8SdjveuV40HK+GbY4X3AcUEmNWCr0YNGhgCJD41WxskCfeTd
h+Qov2zNzFq7pAVhSH+7Wjsj//TpX2dM2H5E3tKpLzsXqRsX6cHx+cKvV6Tram2E8pKAJHBdMjkY
LPwC6rfwW96jDEe1likZLe3Hs7OZruO5NwwL9jfm8fFdkoLkzJf8CmV+RxoBaybBLguGH7x/7o+v
7KHj6o3lKXOStVM5LYSeLzi/VSFF+TWsZ2NQmN8YAiQlrZzTtb5FTPybgqSOske+o69EJG6pJhwh
mW8UbF+TVQQx4gCPmXxqCTqsDKplD4/mzQEcTI4/apHz6UTJPlii73aCrx/Y3hWzmmcxlwVRwzdI
hwTfcpNo1ycU90qwHeQ3q+7Qv7ZevhQoPDkaC1XCiKws7O9n1LmuvYbkZHmZYQBby0zZfy0cafaW
5z0UcpvyEgWMULknUmjgiQ+eGdTYC0+cG9/YShOlVsmTK8fDmHSWtBBWCEq2QPZAoMGF0tVRzjGH
qeuetR0VU0TxST1g3BwkBxPD4GgykYMQW3HVWuwQv+8qx6qIJviinhfmQd9JhPhkXHCrZq3dlRms
8px1rNx5z7u86RMsFeuyvJGugcApZdrRzLtQUvgUEtkK/kI8KjFiess4RgB7H7YldlCrzy9mh5tr
EoeeEA9uuJ7njJjnXKatqPVHQj+WWSR8vVVAQVTa/AwQR+k4VsfP/hqyiuLmFqVsIUmdRZI8mxMi
dsgTym/RR0TMgQRTtTbhyP1F3H9/qU8+HFpp9PGPsFsoH8+Y2hffkwehKaWRsy+aVLljuUBKsV0l
0UIpCuA2ePQhVpBwr9du5RukJyFGzpzDxLN0cf8+/6+UWVdEdI78VfZsIynikmFWxHKnFQWe+hPm
3da567bOsdzNEgTAeYNz5l3PppUHo6kbE/ko5a5yz2o9mNbOidy2ycJqbG8NjlVGbZLpoG99uHWu
1JYxw8KfDJXlbm3tV/22RVk6ugte2OiQR0bX6NMeK7aBj3keknEgkhBLSJGQfGJYLeejAYup86nl
wWcaocDZrHcWJ2P/1Menc0t8GNRGpQhnJH6jjLUHXxzYMcvS+EimLemRa3S/Y4vmsrjVxy3DEqHO
VVdJ1CtUH4d1BHRt09oO4eBq+qNQnIbny+xO5exLk8vVuuuaKIcun8Zly1kYFOcilYfIcJxtBreg
5lxoCZWrIeTkZJ6hLayrkeFyISHaL9PZSy3yQOZewtasGy3BngM+pJAVJVenATNmnKoU08IxXXZ1
MoUwEFvPeQs14KLw74Lbal2UEX2OdDxjpCFWa6vORxPVbBFD6pi0gQ91tDmaTAk8A8tsibLNn2i2
//zll3XfH9g14EVUe/OyZs6Twe0CBD2gbCUuRFkRabEWyW5TNkB2Yy4Q5B5nCXcD+VYooJ6tG2Om
RlUu+nL4/HL0B9nHA7Bn74nzg3wHH+cFm/XNUtcULmiPtnTKqRPD+IU1SOKq8t58E1UahH8k10IK
K/QnSzlZCEBiaRBps64gXBJUNKOic4Vu2xOeDKJbqRZGQlhy9IGLqWzphx25QBShOgd43h+aig/p
CaTXcZ6PzYFMnwo1d6qOALsJaZPAnjGkhomjcREIl69WnZLkBxn/Flj/fyJOV0+z4nQ0XhZrYotY
xjiR4PzwYtOjVi6nn3zThNBks69HCSSxS5gF76V904+GCmxjz31vF8cbtklOOpTUodEIUmO3b3qH
7hLkvPibbiSKYmJTwBM8IxQ2JlyPPUHQjcAqHxgnLsahN+2sorMzrTYgxB0Z4ugXMOXQUj9qNzm2
ElcjqnEuWgs8CcADo53ysFcBOjlg6NwB3o1IRat3xWFlnnQRuajjaplKC2QlL2JTH62Sy/gLOPrk
lDNyVvmj/s9oXnDC9q6/K9iPyizBvAFCYXJecuA273Kn8gy6KVsBetYrck2h7737a2I3m4tWJcRu
jWeOp1wMqksrilfDTK+Y8UEff3HZ+lO19OK1Lb81VG9zqw986URiJ1NKhUteQSYQcsu9dmloNEfr
drMknvkwQv0Ok+fM6ARNSeGnKwDbIgqCMajuy6vj+iAPCOgXmftQ4oMH0hI6QDZTEck7CLDHazIz
bSh5fdnIK4rX4N4OSsjXtAzZPnO1aKbTXOJQNqsnxOyvbLdkO+GUzXOABI1UXpz/TKtKyyhkKVWY
ins5LANcqzSthAyl5ElZ7r3lG8l5ccw4djn3zoVnUIbd1/eN5tjbhsasmrtgNuRKHGxwUDo+PMyb
VIB+md1k1ERnqUFVaq/2NkoTKd6Po3lesxmAsIOrqyylGFqwFFY5zXw0BdnRHspxtFAf82UkzIYJ
+oh0BL0a0U1MwkdbshkNQArwMUm03CuwkiTPhIfIywOegKLxlylhbpDar/7gmPLBLQpi1iWeU3D8
FnTTA311WmEH59qhGE1O6jAIYJZBTRh5AjOh3xGr46vsW3pSBJ/DxTajV2DiDvVxPPVqsG0lZ+vj
yj3DXxU+7KvzNpGkfDk/ZACk0Dc2NS/KtgMsyeQiFvU+Y1lUAlDuOIS56WRn9xogKV4K5r0O08u/
NtzbaexMSutALE497gO8diLnMvClirLbVU4i2AHyl9cs43Z3KGZNz2AdSYgJ8El3CWiKnLYv9JYO
rlep5d5qrkR2aE718pI+k/cf+DAwwkCoOG4/d4y8hVBlE/9VkhaBTnHyzKhq2JkGVuZvwimi54Mo
QSQG/OFned9Dz1RUCpEGsUxLI+ZZiArMGHnIA3C5z+eWyXeGszl83NG1dd7JBse6crvkVhffjmR8
erXUugRkCwryiaSQA+/w/JkMshxHHLEYMKPKoVgeBrBSSry1pMteY7qUNTMJbG3M509G1ovHTAv2
4M/2cKrzHcLCrVPwPHge22Gfj1VI+q8Kt0nnS/6tRFxR/vb9Iynqf4D5qthXOg14A2k3a4RzcMIK
PPSAY1Aa3CFE4mdgf5T/4rQdNV3qHnOLfINeC7lS7beqFoNNuEeJkDaa2uXUFHGhb4F0TdylFXQH
QFE8OHge6xus8Ol0iWQfnftIX6XrF4EKEhd+RU7/4+mreYgndTFDS3Bb2ni9f7yr52F2Eslu6NYe
OSsxHSJOtoODyps71o1FxePuxy2E4KHPR05DW+3MDkyKGE1I5dBBGEuHNdJctNjL5x3lBMRhlD4u
vCHQ5QOycZYFukg+3eym+cpw2EQBic+LhFpjeQo2TO4yP8azj1ToDMu9p6xzDPecylobHdzMC4kA
j2XemjRzVxw8K/PyzdLeL5+JG5QNQcCqeOEJIeFRPV658dMZs99nwHFBSK98Etk1XUTIvOEkdgJo
IrX3efyk31eZSppVntVOokK8Jz+ZQi8ggHjXxyc8NU2OdbRLjS0JUuudSSn+0UetlV1U7DURV4n7
AWGBjFbOgBUajtrnPgj7vscv2kObL7cCFtm0npvv8rArX3w8JiRbRXkgmzHHDkcmVML9seyirmb2
YqbsuMHfvcqpY3+h3O+mLN3I30ujNtaZr4qdO7dd7ula6K3eP/GnJ8SsCQFzNxaPlyNNmWXxs408
1FS1KeqHnGsQj8DfyoBo6h77HdiOvrx5REkzL1nEkpjKwcof4jKkdWHMBybmrcGe/Fx6iG2DJ/3A
Z0H5frU5f5GR5mW9TRB92aBAzx5fMbLciumF5TYzeQDz3LZy+Y/iTXEVSjFyvxAxMBF3J1i6Nqxp
zWwNjPO6vqE2Lj2yJSTM/V1KQef3mZVM6Gbf3f7Vy0iUvFW9eeqd1aF2iMxzEt9W+1jPQCghdE8Z
bT24SUaM66VmDpsJtUSEgIRQ0g/mq3YRKsUwyDvCsBkGT52KCn05hA3KXfuA/pTO8aQvpSAsktMD
X0sYM05q4jybKjjVsKQ54ZMsreFPYpd5oNF0rzQW2EvEvpo0ngXZSPz6ct4+uiuoJs/Q19YYF9nZ
MqyHw5e1hls44eiDy8Kur70/zR3PW7AOE9CGQ4tzDW+RsMcRqT4xfcBnZ1WjLcULBjGJFhB7Gc14
SsycbIzcE9+ObD1K4pbRhyetZ6fiPv4uVPw1xjYwWUVdWN1ZGEdy3K2ezdLYs+DJMKLkJGGe537s
eMnZCE/A3WE+be5O1izi+99y8PkFB5utuicVklDZshGAvYBrckdWrhh091pVFMh7APXiVm3VMdfL
Rby2doeLZsl9/Hgb7UqQU32mlEflEC01aPm8kI5L2DT1UeRK5vw8m2XiyYXj2MsFz7K4aAMwTzUx
J/6/8nTqTgxDV6X3zNSQDUyhTQZHp9QwZV4jzXcnznpgzi+oPwQopNMg05Qj7xXxnQAZtBSi1y3S
6s8dU7PN5t0w+VaDGC+RXD/2B/4Gr1yphVDNtnsvxSchTD8oB2EaN3+/DBbgHEvMGgyURSGcm3rU
qKAon7Yz++W2beBMq3Jebaqbnz866++vSFgi/Fib5tczf8qwmGOAccgWvIhEfzd8cLJcRqwXoZNs
jQdG2ukcoArAm2nJ2T7L+K0Ctal4XXdH4fVPHkmaX06o3ofG7YAxb+/zQSk0cn/wJOejUJNFhhlY
a+Peo1HDpfUXhHrsfrnDm1w6kKJ9TvD6uE+/PX2WZKcf3D+XF6VgCZFrA8aku8b/6kcnSeoTRnu/
lm4wfNb+pZGamSWvE3q5LDDkUs9EH1HmH4vLowXzo8wfR36xG9/HGjT9hxC0xHNpQLIO/r+SQxFl
6K01EFhV/peLXAJ46/5U4pBUWxmHu8Lq/ZLbXQ9teV9BYg5hQ5TRzfuixGraLXPWqvDjI62PeAkj
bTm1JmbfsLMuZD41SliHmADYRDAX6C8WhV25iOw0M+ABakmDQdmXUr3f6ufleZdSJfn8Urp2ZIxL
TyAKlE4vJpGyqZjutap52or+6Bvm4aUFgA2eRvaEXsWQnkiJpaFW+nh5/W8DhArOjUAiiiBdRBwb
H9/n0sGUPnTH3ZeRpaa1glGecEw20NXxTA9VPJApHorGJPcwmaeXp4QGkw5sYfU0vMyQGxoaHF1A
c0Q7aXeHce9EgQ1k6CVe8Q/ybkccul695q7j9YJ0YBrEEVFB8lCXZWa3prhTyHI2FxmTHaVgMKQt
zVbB9QSeaNuvsGg3Nqbu2w0Ex+IyYQnbp42By8WOUfmdNQXhhz+NAti53l/7w6FjncrBQdCDLrCf
b+Evsjcpu7fO1cDRX9gPuB38AT3UmpeSw00yNIW62oShnc0fPMaKtdGW4fRebwqqry2VEhWFBzzH
mcC42maRFRFzcrwzs+2jNQnfFZCorr/VdQGj1nvYrqkT66xzDceQaOHzAlvyilmXVQB0JyVq6xvA
K0EKRruNd1O20kpUNU2wvPKyd22fqOe93VoMIt8K50U8SbUNH9OL2Y4D0zwy1QIN5BTYd9I6xHMa
ffETvhyMAM09XByoPI2tNSELfaIUvK/TCgIKC+8CbiA0Le7ewTwSJQPycGCkmB3JwSJnsTF1fleM
5+OuQyJHhRjKUJHGBwQ+T3caUwlmbdFLe4xhp9e0rab/q5iYp8sVH7eOPT0BC9Hc1Iootz7wBbn1
f3/HLcHCYZu+7mq916JWR3F4FDrSPyUQ1kZTbAG46HXbVJW98Y6d7sSfJ7GXEP8WHbqT0draccIp
UalpAy7vrHyo8Faz6RdV5m2ZHv4lOiuRqURAN/Zitb4JPuOFTYHuA5EYNEMN4dqlWdS0zKnuGDEg
20TA0jY14WOnRzpn+10xql+OpMH6WIdWBGlL7XMOkuvxtw+1FxgiavgMnH4J8+ENZAoLPnQnaSyu
Co9+7gzz7lNVpmqblqy2sGKWmlcWLhXEFbDMgnw/A5KxfaOSiJlDWdCHk5wIW1B9YaVTAqMnsjcU
y92SBUlcr6hlDslDIT3A4ns7+T4jKTPJCwYbOzOkqdAFLTPSn6IcXysIwEWjk0nq3mdpXjk3/6Gz
ru27kgeqgvVb/ZS8UKrJzKwOClA292Kd56uCa3muIIeJ/nxC47TEnARjAPd4rvITISWFpP8JsyRP
JDJxSK2T4GkXC9KBQL3rGSjhJ9aHi9hFEM9o6Frhei8VuidTo2D992huRB4QbXmRV5S/EqL0np9c
QKPpCm6TQmvkzBEaiZnojRMqNz+Nnixl9Bfa4daK7Ux4M/1QOqNWq7HDIwsX8sSdxglicXhHYJ4E
prJi+FaU2Q24RKSLaw9VhenLjS1hhOWh4JChMLaveRD9I7lYRor8Y+UORm1YfxVGcWmAB21OlycR
/D8AXTcG8AmwX/aaMGU9ahgzwAz3F9mgbi1f8GO6Qig+JUSme7Q3YvRjmNmdLpdY/jc8NGix5jrU
H/lBbUcTFIUDwd/HKYYD7jQEWFqo6WMYaTFAQz4kxdJDhRb1pHWd1opAeqWqPo+GFt9Bs/Ns1Qga
JLvk2PbASpmH0HrwZV1M1ku+f+Xq0lGBHrYBCA4Cv+BpujWMHx41h0QqB95GzKnye40rgBBjlT8T
f/DRbpeVEw1p+WrV8V/45+oggpLNYRuSiTDELZqTmeBm/mBG1WngtP6BLeJX8R2NiDhx/1n9ZJog
lLzR94yl1xxJv3kjZQmOa7jyg2Ko888deEf0U9qHi1pulpguYG9PqpwQ3o85BgQLobjIc6sdwELR
28NuWFGVMSrs/vx5ZLqC0DqTjJr5Wu4fcJ/BMXfUX7w8ulyz1Df9apJk0q6HGji7kUIXNGnzY850
aoHLQgjy9t7liiAjXtRHpc62r5WxJP2urpDGRZfShV0Vym4Swct6fU/DGsEpRgp78meHEjT5nkqW
8rflyvlPZr7Foje9fOaM6xy0RzXaT6Bzlnp0ky/QakPpr07c0Bs7Di+XBCQz96G1Mz+lkill7H3G
w+8TcZ15YXjZQ5i2ofyJp4qu4mqM/aZlBupGcAVLMEVen7WbfWsQe3LhS3oiapXi2isi14ma23MM
pRzTPS/RU5KvLV3JKBXOfSekSXPLaH1OznxhHKtTfky2cS9YEodHvtBT6goo1zBoaQyX5AdGgiXx
C5k3QGdU8soOgJkXDEX3JmfloreSSWo+k/z8L4VGlH64WnhobH5TbNU10QSPJBK9mza7xWo6olmr
paE2voWiYArnBqmOMv5BicVEefyuwd1oooUzXkpDuIA6UKT0wSKh5KogUKyXXCMd8M0TjjTxGLXL
uBVDPmFyN0FV85NeJtAj+IQDfvqMi+zyapTO/Z4yUISlbdjGDh/GkIywgKKg4NIpwJWpRJovRfex
AiIMHEqWmZZ3sERde494F4KyyYf23+1/wCJHtszN6f0ilUzZKAMxlU3sYGPkR1IJrXerRhKO1WR2
zCPT7PghZTduQTkrhaBHyspb5vW8wriX+95R87BCDJMG58JkAijeUhBxpCF8F9DHvBNmA9p6UBYU
vX/XgO+TGEJZTB7ZzJU0x5OzDzsLveghOAdQKK9TEQGZZW17LxBy4zyLQ8jYR28fiogHbiWfAmOX
5EeM7cPnnhk7og/jmfjyDjCOkcPr7h13JwjjwSMygP7fM8GRQqmj90rONq6IVCM6EZdyBY+DHnjI
AUwI6XhdrNWY89t6EE7Gk6z6BbWeY/1kuCCpHElgINi9RTQnVw0CKJFX/P2Ur0imxXCO6d+d4nPc
pP8o+EdNoZmrP7FREAFfHF1BuWDXVLSSNaUDpzACrKeI7x7DVlyqe80DGmO4p2FETeUSyRtFrotw
7QomY4/TD4tJBc7LeXjJfwWPQudg0F5Aix11lbkcjELSaNHOt6dTtMDtxM42D2EQXC1IAqr+v5mL
GcSRQK31VOyj5AXOMa2DXrlG+LK7rjzRfZF5c4Pds5LWH/hkAOIe7WcF0erX9VaYJETzJ1C0qvv8
h0HLpU+ceA7Ztap/nRvJIPG1M/5dU2oGWsaqU30pHuK0ryUxjaZDJkZq2SgnNUSF7WdrxyUvZRz6
tqzRHW5bWH242hAkK76xGiBtvRS0mJ1G3Fx1P2DiiVBqCpUMu/sHOpWUw5J2w1oPqGNksczJ2bIb
H+GbmG4F/ctJha42XgpQwEvbU99GrNNhsp4Md3VZPGM/7xGUhuFyWvrRKm/vwf0IjNC6pHPI7t3o
OTkidgSY3OS4OB+EpeLjdbHdBMFQA32bJ2LwAoa1P93cW5+q+0d5Dc3+hsLRrTRUw9yh59i2VXzk
NFJTdfeROM51jHtQRiqLq2MqRgKdCqrtPJ7NDkwOiAefxBIsKqxNWChq1NN+rGYm8vZNFfXathf5
ooqeWYdhl130XBjhgv/cRE3VhnORk0RISGZo/jyLwnykGvqSv0/M5rEB2bPHe/PqKI5IB2R9RO8u
s6USAo+UbI3bVjblF1RHMW6VjIrXD1Up+mdC45c5fpiVIhUQk7iIoGFsZEyYuI7XG+1BMuLVOAxC
pKApMG4qnVyNjEB5MDjSnUMZhRCcghNZ6cOxAuKTFWFCicU8vBnjuX28ckwidDbV7f08yfhGMu0o
PKVFQ+6X8nn4nKmJ9Dl0BKeuH+q0CNjiLCcwkC+JZGixD+KvolkRlv75NkLdHnkPYb9qn70xSS9W
n3xtJTui92BEl7hb59WV297OlJP+zKOJEVJkMtZ7MjqBaNfGWwXNV4KUGsImr9nGcrGOMHjJOXNT
l75dxVaSTX76CnCwhsacfxHLGyWZd0Xvp/fbEiE0cfh9TVJEnLj3llBUXDN74Xaf94Y44Z+gfyso
uCDlEECNOR9Gs9qiN8AwPYYaphlrIBDUqF5Z9y4cWXybg1rVPsfMDuA/tV6GzcN2Z1A0pjG7deLR
ZuIyVK6tE16yUjHnirFoosTCvZ0//9l+LPL8Xs/sCejI8rTnxFGoMp8hoLCvmkjm//0DP9fHj07B
gHNIDE3ptwNvlweS9zZbLoi49P1HyaixVN2b3oDK9474rV5jd+uLULktsyOtFJZ94zY4Pjy2gCbN
iN10aiAfuP2gLfSqBaQ1703d9LlMG8rSCBYC0gyKWAVhZRN1tBu63bWJ2hWdNFXXSWuY7Bhj4a3O
DYoieRfTR3wXtPdzRtt7qwkv6w4X4ZJcqxgH3GsOArlucomlwqYOpTE/sBdvPj7NcWBqNyDjDtkm
fcl8HGV6bHTmbgnr2a1avPo79pmb2pYcpf9ptAw+Z7CuglW7b0K6DrVZQSNv39f3kKKCoPSbmRpw
2aDB7UJ7r+jnvmvvMm4InoGpXeqN0mCPkxxh+guyQPFBYjYwbPNGVz7HrOblFBa9KECvEU7e7n0E
6FnNybSgPzeGN+L7FlfV4BDhcOnidEo/4adWZCZ3OR4QxCFcZ9aAEZfmVFmE0N2vuyD4sVQM5R6a
nULD5Przmg8+rJ1jNqOa5cf2vGUpk8k+7I1yGoVUxxX2PVfigwLf7poWVqyF83ImXwiq6rLx4wOs
bkiJvX4v98ZAkCd8WLi5sZnWNORP0WqDWaoESPcSf4TAnVyfQr3kwHYfjVovZvkqOIp42hvYFu9l
1rRGmdUTT5rESTkVhN21yBExMP1ae+h5be9QH8pHV+Bboxit3pcMKAQ7zhGPfZHxXP+qWSWqqUt5
JCuULFCukjfh9MJ7TgRo3rIvWVVjQH4p7PM+AoDh+AURPsL9HONwdiuGpsnj4AuMPlzrKz76VINS
Mx4FOkhUS5MO3+A2rAt/xRSzvmxjACyQg1Ew0AQG1YbWW+pddp4AuPTl4N8XX6iIj3dOSoBIOA5S
Zg25fGdhPzfPJULE/Hk8G4ftQ4aYt442jE94yn0u28bWB1WfpnQRJRcu8R92UqmFbv4JAyJGkIaz
3XizVwtIS2D70lVDMB1GWqTY07J6tex16sQbat18N1f2BFRhb1l7GQY4y1Z4BHLt3QVCVRbE8JJ/
wyz67yHoJG7SQKaWG01dJI/JcYTCt5U6mqWDTBjDW5AUWqZbzWg8JsMSSB1Sv0ESKry+EwaSl6x5
yMJ073zW/R2zuhEfalE7vBQHXDM9bPd6uvhGljH+aerFcM8Mdjpmg2wes5dOl1mFNF07vQJMJ4Jk
fVogv6iYXyGJNis/OP4sW55709QX8EUMngTc03twgE5PqUPd5TQJnek5r5ueRCZrB1fEq4HJZvzU
qah+y+9zd14wbzT8hHaUkbOS6FhLC4kvJK67vRSpwCRdR7E5mVbcBbgyL8VcS+0IgveU093cW5L7
kblNFoaGSBXRbf/T6rxVAhwLuafkvPgwswUA3pJ/JvJiQ9sS8KK5C87fSdWtHGyHeBfdimn+x+b/
Iy4g23SdIIqzQXOkPdBzB7fonvFgg7t2tMle+lrjAnB+Gk06pfUf7U9jdo2Gwe/ixZgDtR5qePk0
coKIoDKBEy3z2SBm1PFCu/FlFVjUrhGTC9s38HnGR6o7WnXUoTKzC3DGEQeKmyqToPoJtVHba8E4
7tRQMIbYKR9zPCh3BM1lhUVNF7B1EoV6AB/xS+BxfesXyBvE1WYR3InLEyNc3q8O23J/v1RNT9wt
oI2TfjucB5nIVkIYlQCPekS/OAY0MIag9CusL3AhJFtFhh3NUP6HUELCRr/2PfqiWtxbifC37e6I
g6EpGwQyOIhq6JFlBlErNKTRdzAIDoGIKwSK3X4KYOxZ+1la3+4IYUjJzW3P1dEnhAHU5iIKmRqh
wPLyApRGfgtCGkFUq2v9DeeGU1lcVshFbF+ScV8N1S/QHPzfc/LikarvksNu/Fm3mQPTzNHAHD3/
Pjvlg+5Xr/kKikf8/rX9UUU9HLiS+9RMDwjevOkTroAnWl0Rqwp35P2pAlfXc9/LQzuTLhOfOszl
8K55a9aqZAw13Rk0BmavqgDgMLhnIXe6EcpjXekKPxj0HqHNnwP0IQBQfxoDCjsI6cRqhXY5gpji
MDO97q3SLbyvdPmK1+rZ1FkV65u3ESYD+2UTFPzq3raWy2Brym8Bvd+3xoHCtij/J+rx+DzNJdVa
zDE3PAsj/hbKSECjHBbbOTk6J718BA5jKRniEK7ReslQmv3OGmqofWm5SgY6CJxoScPXrQ0Q/OKb
Ul9hq4SBdoXsxEtO1e4CJkVz/5Hh1aCqVz6j9vEsU8H9Pp1dFQ4eDJ/32o69BkZ5uZIrov9Sb1vr
nHbFROdeoM0DODoSdy+xnlCD2QfyBEes1rH6t9P36DfTI/+l+B8xtjqgmdLJ1+7CwcjIfpn7TSZu
XxqUcqVMe5H9imyhkorM5meAkaFYRUgedKwkYnF+alCzXsXq37aexIwKvDDtTRWFIxBwsI4LfffH
y6eyMXEK8TPevjmoMnVDSrNbFao4qZwVFr0l7EcK+h/jw2XHF57RttO4zWiAWz5WIe0ZrV9F/rK1
0LCV+J1T761IE3BRR5iPO8fMaucmJJYpI7IS0ymlTBSJMSbKqnSmalu5OTfiOb+TqmF912OOcXzE
TQ61F28AiMgArn08HBHGCmBRI7qBdjrYyoP6JRf5Ie5dgrEsFJUJmpdZu8BNTlqiCvFhseUVxo5V
jD9UEPNBCtUvkoXho5iK118HFnIjM1iDSoKWSBDJPrWBkPO+bR48X7vvo9BqQrsECar3sfVodolw
iGutdRqLJEwcfcd+HL7MbGR3goNBTnSKnnyrldPlPQrE/ltIgeB02zhr65L8NafPkIgFPDDn58K7
TS7F3LKv5n0xhS/rFIj1p38VhwKB323a3ctCtPhhcpyCluTIXMCzXCBg8slWC447CP7+XIKV/4hb
yukBoQA9mlCvYFY+cf9c3TsCfEgSCh5hbFA34uDvHL26GQnXEsOnwyrMTerF3lhluQ+tk6GxzfbQ
pAnkiVdK8jD6d96LrJIb2xjdYmsdSeDc5rs3PFF5AoM9QhBszo1DBm3KsNujq76b3pQ87KcnwjS0
fxjOsgr53JU128bZuGo+xuE5plaKTQt/n5STrsK7uOvCmzoneFBQRpa2h/A/WwwGoZo3ZONcRUsd
7nRcCVQo+UWww7NZg/RAuPSskwMo6abY/i2lKyQ3keaQpDkgdDZZcKxjrfpiF1q4khAWV+wkqBb5
BOXiITosnCFiaZl4TNTyhJUD9GUsQwzvxeSKMkJZqYUkenIhHdboo1K35XzNQLElMobpTc87xpPF
PnFUMMdnpyDChjP7IzoDMrvy525xK9yVZYctXmWo2IEP9LHjUxRvKx3zAtmyz4Mo7hzZuc1+mYtT
urAt8zq1P4w0Lpr0lIKCPCRd9IRc7ddO+N/PNFJNcWJONN9JuaEwgJ10n6OmRZpLiuoQTrgUeA1o
bSzV3bjw9SQad6UJWwilFwggcXuK5qVwzimz5+RTfsfFemLREa8wnX9yrmpzHZIex4qmH+J0BH8w
d8DhGPDcPlhKQH4mbPpcb82J9RWnTMvpJJ334bljPcKy7n/1Uy2/MPRXfcr/Juz57Z+o4F788PU3
bCDfcoOXP6Q/JuamVTZ7xKf5BMMCzJGXlddxrlbbIAFnDPAgzrUYAywxSO0w8ydxY6759hT0w+QR
31CHqR/13/I82H4TbY0ez/6u1MOqPWpmntGewb72ULEu/lE0wulvReOiqCSogVm5DPf7GaiDIaXM
hCZs2eQCdL8x6L0xiBi0dB+OLCabcswRGvCD3GOkrsXwicsAKphp0CJI4nAl7wEPS2sug360JVdh
sHRy5NMYL116hTFmoBzD8/wfEVImrdmAnlfuz5q7w9fyvrj3oVeGSGnslghW1BA5Pf0q/zyj3Vo5
tHa+7tbifnHwCGMPNopxPzPiFpn56b2Gr/Wd+nNYeq9dN4jbJ/v8keTsWclwRtieMQrIMbAEgBVb
Y2aMWLrTcE8WU+bFCUK88SxbCyjnRG2A/+HAGuwGzP1uxw/Eh5/Xu7Es0Vq4W97f+cvFan6Ufxzp
Ijy/t1JCfSeEPkGE8R3hyuRD71cnZ3Q38O4IGiZIR3ORUDsiEN0eNCzuflYvI0KH/ZNKbUS3N7jT
/zQQTm4nAy3LMtPVkOcVZM79ERZPqk/N33Pk8vNUB3MSCZ//wwGeZ+yzwXJCb/3oFpARFjr3KWzp
n0cAVJ/p9CXEtOBuC3Bfr0Mys00ZtEag7+X9hCgYgRpv5T5BW8j1TCS8C93s8XNOdP8L9ENvwHIx
LpcBmLc8Qn9sYHorc5KD3rOqfEGu06X+gZRWTSEaWKk4PaEEuJDkH2c3CvPNpl9KLrIQlAtCKK9r
AEFplgp+WvPfS/QPWA5UbcwlFCE1KJDoAHjeBZXbfCEcoYNWwJVDXEQdbF0dVJzErKI4jiYI7cGL
FCzfnGXjtWghcDdVENvU417wewG+9EeSVMXnUVs0ACVlKLx6DIMkVWmzMEL07WcGI4581gxqlkzr
NLcCKYJoISoTnAhRTbtwTKdzNRe2El0XejoxDzoT62jSEIFGE6qpKaS3BCIVYmIK4THoX778rVhD
Gf3sUCzgbPWA26cjuI7oebnF5lFjb/s8zHV/ePUmZsXFC19f29wtytMevUncEVh4ZmlSwliRJfbX
oD5D0a0KgBnQIc4PSJRaeDAPoTP7bgVCV9EB07L2Z2/5PLNVTqntJ3iVkh3/37ItsOTXXOEFjr3n
bnl6npLd68JleEBNbk9tj8H7knSP4uNxWteqRzm9ebAg2jeFkA92Kh2mIeHrbwP9FouHCDRrTue8
MjGq/bmcV1ZB+F+NsNLqaXFa734bBSoSrQ8gkOHqG045+KLImWfx/vN6PLUOV0+d251pYxaf1ypl
aDO87mNNSLZ9uV+EhVK19ljtFi2fv9ma419kJKuBdKVgVwcRmrv8j0trfUdSv4XuZUPyxHTo4qk4
UrGf1oDqGsUZ5XNTmZFpIgH38DZHEH1mqC1wv5EH6nwvbSOUZVoh/VeuqIALR+RUggFA6fzasBUU
LcR/P4+vn3dyaDEkl0p8OeYDjjhOggLzBqdKzXWSZqYPtEba4AUF7oesQgEXoWtaoDJJrJXdFSHj
L2r82hlZ5ViROS8wefmmy2G9aXz0ny6bAO9GychwmG33uKLitB+lRRCf5EsKI/qKvl2+W88aiChk
B2qow4IgBpkHhOOOPtuOG27p0+q+uIggPb6361beOigu748Z7lQqt4wGgzes+P4lq4Lk5IX8laZV
n17PVa8S2zZSzjhq0ml9Q9azQMBF+ef7i5BztR16bBrW36gSamLvSQLibNdbl+XWYI5RsXQTMUOg
WJbGCnEPB9vXpxeZuT6uNGRJLlzNfXvM4h6Nz7woNEjrpgK8Z9NqGf+R0rwckrVDkfgbfo8bH1y+
DdGMcKd+lOfP8wwc57e7GQRoCMIY3PWmEDBHB2B7JljbuT/pSUTqA7M8q+HlDRpO3GR+Nz0CiVmc
gVAelHAMDEN9IcxT9Vut4/CCGcTug1J+GXtQGNJ5JVZQbBcQs4n1iroUTjZZtQeuK1aTNIu9hlYQ
cHh6X9GnWTRDzePuCqOqzk1RbtWVoYyRuzDUtvu3kcRxtEWeWthTGxJunlSnDMANH0Wotpfyuj3N
A+0smyDQaFhlcPZHEofW1nU210A9L9/nzFnuUqSt3mzvhtmJ00vZYVars1MPChnB8Ls2EczSG93S
tREc8iufE+yMSYhjfND56s1ii4bFGUveqnxyDEkT/vwuZ862otCmcx1mQ2S57OLqMHNB4AS/7T1B
AEUkGz4Wb0bRottV2kbN0mfl35jxIY6E2j4XzsDfKiNikv+zswEIvt9f0/MwplZQIifbSjhBy/Po
rAcsj+0QLhQHc/UtE9ni51NAK6oGb0AVwIUG02/5kfU4HE0v/6Hk3eZGvoMwbpRr1Pg4n0Gu3ane
0VDQWxQSgXv6McYes4Q7aI0VNPYhAfaRRHYhG5I+3f2qg7LGKncw64BIW3VxOTGazlqdHW4VB/qx
GZQZS0E8C1LT/V4grPjiaD6Crm2791L8vEXS+GrJSXQWWQ4O0WCy6LMrJpf3qP+rxXEQpimyh6SY
C+V3ucy+Zus7O1BnV0h1qlsgbKZV3AThsTFX5VB/xL2mWBJ6DPyQ1DWvnJsusKJAAIpu68bpU0kW
0//1wf3xt1DUBSF9Bo8xn4OR26PKnPw7SZzw42jwYbI7SOU+m6UhScLMqm4gj85rphC86IS8A1cC
/9dOVJXhxWpyAR03skRB+/VEMNnmqqgiAksfPfpgxFV06vNk1VLAuSJ9suGw5DiyDnM6GWGTRMEN
IM3zXg6zOBgwX3v/Y5gZOZJQZPfqNHTsJhN04SQDYSdQpyk+gp/WZecA3m77ouOEO9lSjKl6yQmd
2zYRteo+rbYUpahYadKp4hON8OM9j5+IaIjAfWi4v94FMbg1pR0QpOq//HiPd1/ReMbMXiaFxLZR
07OVL48IWXK6oF2ngcQv4Cazcu75KwxP8/VZYEMmPwDr1LwVl/ZL534vNLIVM6RJVh5GhKk+lidw
Pw31Y8CohGFeLq1q3geIScHyHNL4asBQeWbhT0cJC+yuYRVoL3tphYhSCIG7c/AGcB1q5H9wTQ4K
XtoS4GhiCxJg9XtXXlKmlO0KE6EWgo6nBfP+ZX4nLPjUNvQJfLgpkJjMgh+WH65qh4uJ+mOuDXw4
FzfA+9HiVhsWOSEeYQ6suHZUbkP3A6+QLM2NOoqrYUS/TDcbbLDpQhIiu0mYX68VgTtEieSUoJ/b
j9Ag2aIOO2GxvDsJ+OeAtfiksmr1o+rqCPqbyL9jRfVG3S28zAFzc23PsCDqmS0Ere1aDpvu6wGN
fE7fZNlXEq8uws449rbtNeQNON97KHQkPhOGc5yMpGIVvOeZrCs2pCGnQ9NqSsOEsSnw6sb/2Rwx
khiBfKrNzj0BbahmgGmuU/GyGF/K1ncuKRkuayGHXVMFfa/msvAJ6dFkX865cj3YNofd0LSOkWg9
15wFKfq8yQme0JT3tdYzRzB3mQRvcajyjcMpY5k9CK46CGrCIGE3I7zS9//6StY0fteYkKLnaKl8
4ZLJL2/EUZANi88mT0L6uqwmoNPWNM/2XkV8NPBu/0w+QmHIFu37z2o8lLdeeQgVCT3fcb9kIGia
U0YGSOIMjlIG1N903K50sE7PromEvHxq47UuFctXC9mkcZR3X9gIppugY2Kw6n0qdZ+U4CMfo8BX
Z0O6sfGYP7xHngGrDA1urnzYUDI1RqJ8nAwJx/gCb7jVP3BmfkO4ZJ3Lb9rX23fqOAp0xTyJdDeN
F/myAVXKngeUJhqaPyFtUPpYyjgkPnBvzAvJx0gCweR/iG3rEI/9cszOHakjdaTDdbzTo+V5sBVK
9rms4MJVmJq503F8XZaHiCLAw82OqlXGD9vwCVWRkSyX4x7i7s/Kp4cHgSvZ/T77mFlugv4RdTGN
CvSfgIcdMqdMZ+we6YTxlE624b65iM/lRQFA3lcUIDNErgY4qbLJFT8ArYWqF9PyZOPG0fUDZ/xp
9tbgA+HslhYeM7m4uRlFE9NEGsOknQibCvrnFylVx8JgVhcf0cISWRiJ86zHXh+y2SdKMJpzEXA/
mWiN3QXgcqGNx6Hxz4Crt9w09GkuoY6lo0bdecHL08HZQPrxrKuLSxrjq/G6q1ftC+5NHkTzB5q5
5v5AVAotZl67b8SRL4G34I9UBl0qFx+O0ud0IF/etpsckdpagZhw/EBiSE/LljsPwO9MlVoqUP4t
nZqk+A0s8PoUlAuQH/YvPQ6XFTWjhzP6DMxXb2LuQen57son5MOGYX2iSgmBlSDEshvXvSRlVND9
bzAtQ0iWi6GUop/W6ZOxHn8G0EwW3Xz2Pcq4ndX7lL2bNX6EyQVbxygPC7jh7Ggc59zt+swEoflX
RVf1D+s2AC5cIpT/402wtEolCbTDXUnCQIAgkt90Pwxz4erZq7lq+No4DY/Wx/3+HawVTEEWUUn6
NETVBde/GxbZuZk2YSt0pwWSY6XkvohLCOqciioFoiibrgWGdWGTH9t9RbolXLnigIBU9C8SmX1H
yfFQ/eeXcl/ET7moUeVOt1p7N1+46XuszrMVd/2RhndsCm1GlYakfmSUgYfYCdz/kDVeWxx2Xevc
sFXAQtswQRfKDPLaN14hFiw0/SnBAwvl63AZIzILp70oVibjE8YWG0TsY3yOsleKsJU8c3NCQwn3
1R61I65od42mF2qU4Lbla3zkP5cLfe9XtA7W0ahF+PoKt+3xvd87uwx8ZUtbQf2VsRQ2S59Ylcug
braRZkLsQVW83CcbGbt3hZhpkKRwK2vQ6/fXlx8CgxUAJpE+d3ZNqgdCtE9HUP0VkTvbYesDOLZy
GyBxcnpzD3TrGQUTiMo0pKDU7dMYJKOOiZ1rMYQAvERgmgZUBEs0WDT/CqL1g7+IOixZVEOSvymS
x09+Gu2AXxbjuVa8atVE2IjOQwPXyzo/2+aZtKdAqfGAF3hYED4A+zxoBwq2r3cFvNG4G/+i/E71
BaeJlAJjl9g9bENAA7zHFt6WdsDFfUt9nNY4gqJeg08ksu9UIPNbyrKKt7NiFQ7raW5WRX2qs/BY
ku/pkN7AYzR9369BKBT+13rptl+iA3mZhjOchnyBLAtJz6mY7MDRkhpkAyw9sHIYQAkggPLTNAaG
1ant+9GvYr1yJc/Q5XXdUfg2UPglJPasDH0tlH4pkuFOnc8Ke8UFUJIbN66Sxg0MHwkqMrByW4TW
G8mHm5nRRrdzsw92uDQ48PViXYhGkBK/mcRpIKtgnDxkJ/ISSvS7RfHrflBKNEFt01vb/vT8U24Y
34TYchTBdi+esjElj8J2AnBZsgaVGH7E8Aq0PI3UFxpCCSak9NGy5Iajly9VqL7YsvQyMRRKtsA7
676xDgQKHqGUq4mn24SF9K/TnJuLEoCUwKrIl0i83v10ofpgOT+DIEUIhIjCtZRCSzCg6MnNtaR8
q4chyTbNKbXlnzcmrkQYbQ69Ne51XEl3tVH1p0wEv0mCbmqpSteVXAqvoXdOsx2QtOGlRjQ5xO99
mANhfIIOXwPG3crqTvmLZjDEOC5sBc+lErH4v973wCiiRU0zC78dsU0pXuB9tfmdONvZksvB984C
7p8aaBFWPcRlQ/CdAp+t//2ngJgNuDgf7rKGv6DlNqS2n3FScDM2MCA6ne8WVNKDBGcdFDWddCCK
KA1kfh8F1hKCzBKgKex8XTZbdQ+54H80YGMGXtk1NoqcDtRux4FtFOXUJ6flWHyKMTqjpcjMOcxP
NgoKStQ1qmpeZA532eFD+4y6AgVGFrbi99KbR8iTt45liORvZSXRB0/mw0Df3akyS8Z4iBUtksBR
XiV5LZZdEmdTGnKDyf8wuZ8IyvcCE5hJLWkxEzmZ9zv6+7MZJKrmLN/VTYJg01ANYiJqw2+Qx88r
CjHAZq+T7JargoO/JTrdP6qEzNTW9uDCFwq1dRJpnSMl+bgNqz7IKFPeciN3RsWed1zDQxBTQ/ua
7ySp/HulW/RYUyJ27IoMcEiNgCO0Iey4FOGHVf/3nclt5S/Tj+zV5TrAvzxNdaMJAu3Z2cTDvh7n
KtcfHMpgA9Qwxqp6KIyEOv83txV8Nr3m+EDYaFxdNqRYWIR6WkVOKAYWTMt45OUT6Z7YKFjy+Mrc
ZcSjDi38XLMmmmoBZeyJuAE8TR45vzEJunNmxUItNMU9/YAJxMmO7WVCk3VQDKdVu3BtkMdjV9FB
bmtwGfU1bcjElzAQ6c83ETV+HpN1+kgbTX+sFB1GPyCSUV5qr7oPgURvm0t0C1R9ApPBswpuSgis
gKboNu7drQRHJZMifXcz9K0omBDbzzEwuZDOIE9N1uzl3mDj0KrXL84wAiD0sJcH/LcTAS03nzze
OzcUFRxFsXql6JrZntXL0RnSazWZ5BzGCvqLRjxL2J0tsXZLemvGJb5TVZObd4BOAyY3y0cWnxqL
WqeY63f+eLy35bqGK41wDDvFVeBGE6UmQYL5ZFc/fYPrayNefWvujgra5dl6k/hGlTW1uirBWVWc
/OQ5dLNgjl2d1yFSwAZJvEbP8OLEZeCIhZ8zIpZ9Dtvz6N7GNQB1rzwvuwwliJoTqzoiS/+wT0f2
EavQWU57AfsM0wzshuzJDoGkNRyDnIxmFYC+Odu1nhCpY74PrPjJ3vOfm5/i3uYsKRvGOklNFSR5
ULwfcS03HKGhdVxSKs/eQCIIPntZeWr5m+KuNc5s6QbQfevSr+PeZO83PEKzCz4pRzv1BW8a0JMA
Di4E0k+oMiq7dImld7k+I+Jhs8/86L0eJHReUdSXyt+lba79c7z797MzlhQL4WUTm5qwAXEbme0Z
xxhfSs27nckHc4qAvKyLjJRvR5AiQY5wPnTV2A3adppoxaWsj93JveAAuPPBs4mGCGGO8iNpPVsA
QxsZZTqdd9HQLnuDuN+ji0DTZ1bsf4k0jBAbUE6mScxggz8UgPmGc8FxpX98PJbTuSrtvJMgJm7O
bigTQotO2guIW6gxXbgQrR/ZYGZ+KkumnBitzLZzzLY0zCm0F0G3ahEg43XBIh5MgAOOSrMb8Yr9
q8dn9nL3uQn5BjjL6IhnY1K1ZMSgiktbQ0Ql++aU0hAMBFkR+r4r0e13Bqvd3NQWAkqEv3elA7Qz
k9ntLRR2JTd6d0K1WGpLPObK5MnURmoI0CaXFpVIGKl9Dc07LGaiKOFiqe3m3IvTN7MiKU6XcuFg
AqRlYMopmD4FtTvQRAs+i8ZCRjlHlotV+Uj1NgCFNXk1drC96qdYGy2Jv+uogebKjXe/momseEdH
ypOPcWrJbXJdfMUHvrByVozK2ucYsm2EDIwZbtN0gSEy9+35E9jg/nCWF9QkPZssKYnSbsLx+3RM
kwHBGCSsbqfGhRzYlFG9vYFWLEgqxnt20okPiOP6ZrwMst/FaF3qosk+hqguwqw/SfQiV86eHtuz
R/tvhnuLb7N5XK9IvSJsjgbFR21ccgZ3InBPKXPlMO8yPR7PFQH3R/Pq+AAGv+Ya6WowYZkt/Kdb
68OefHIpbUlIOGb3POkEHapV6eBSHWvrazF0efHLEfuerktBBWPWgJebHFj217mOsoYFpCDUL4wE
SNjni3DV9o0++pvaN7K9lFRB7HFr6xPuz35vDv80yBuxOD07BiE9m1qJhgFcDcR+MYZMMVNWxkEl
iaIgr8Uf4mcT5lZPPbrZ/roKfPDmLNAxS2OWZAuiR1RqkmdkJ4DGNm6G8PJj5i5bGWvcCCmMljLM
6l4qiKDpt5sLtVz5k/UKjlJ1CoZWavJIDji46E1oKycShMq7XdVK0OHbKzHbXtJBx/VoyMZfzNAC
eLhxtS6m/umR5cUVRDVmfMdcAyi2Ug8okvQ7w5P69cSgnkRviFF7arZJZHn86cPlq1Hp+RYGlOm+
29uk4yvteKRUBrmW9Qo/HkhIyGupVgr0/wDjd1lWjXx0a2i3wKzKyDWcFD2IRSN2/qY2ilojeNP4
ndU7sHSZiF3/Td+u+nTmSEVno3sFmKDqxIbwXPvz1kCKbkFlB5VSisp9OB1iF1Rfz0vhUpNvD8j3
hYbjLVqfAtAA5nuZdp2vZaspzjh8RHOpcuvP46TA0ssLZlny2g8kXQVZUPJoxV1FzIkvlMsEoASH
QnHPVI+IF9SIvELWoSJbtZ+nrofYXJd0kd6nO41UdXurb1shKpgOOiq0RSYrrbqlQmAFJrE4EqP+
f9uaeL6VwUjmlf41cgLYJgYZ3x61jWIHCWEfcxRs18JS1Wbw/TCt6kQBvoVDCcUgEInQqH1HFC9n
wkvuq6pkPhL8i3bWPakumHR1Ed8is2jKqmEioBIwk+BcFHq2JOwKn7pOvnyLXkS5N4B8UhVxKiJQ
fl2sd66VkF8255Whtzrdh9DJNol0Ks+aHlad6GKaUZGN5HRY9FKpCT0tuPAePD7T43O7ps1jHUOv
oz4hniJ5H2mYbnAfHNGVi3LfUtThQM/s0IEq7/HorSLD8fEJbrfSPjy+5foJc+Io3mVSMcOpI9E6
8kFjuBuQJeU9vfXdHozuz46hNQmUJYof4zKBzVfcBzBxoOdQb6FwsqypsmKUqTI28CheJTWL9Cye
ZB741EID6rUiKP6DF1NYst3kaqnjMt7x/mDvEpAel0zTBfnel2x07NJJph6TM1Tzmr8jh2/v+IBy
cwmnWYTExPxvEWZ5w+ngzbeyXaLHTTKbKSlt4gVXoh6I/oQHoHH16T93NsJJSo78yznCjQP3G7md
8TTeJNmJ61SOFtRB/p8qNwf/CNMBHLCVEg0a5xKInvuTZKDUP+8S0J6IYHbQrwqnWxWDM3E2SiSH
YgG6c86teujuPkt59h5XNDvNHBJWB2CIgEcuOzD5EibNp30TQSvRgm2GNlLOZBZteFNYqx5mhHA1
h6rhDYf9iJqYiaSWP1+l9fkJuhHagHax3+J3J4J5dPDIsRlT+JC0PztBCt9YzYKzL0VI1ELAhHs8
ihh75No5kXvJQa1Gbbz2MSp0zR+UiXzotv5fLEJT5ee2t74s9pwOYUyJObN/uRrQlaWs0NKNE80R
pA8YPWSMWoGqZEyoPhqU+4KToWuCBdAXkohw0KqkiO2q+EcZ662vI0OGk0tOhz8sUVZdvxVZAe2e
xhcWHoAX9Jyp9fcJgGtv8ZIlzwjVmzYzIKxDuTKptmIQXMWL8d2L2uO4+N8s+Df7xQx98Zkqu2uw
UG6VNiT7wuI8aSdKpLdbc72qwnTcnI99EF4oELX5MDZaGFh5KSoPd+5Ni0L9wuUzpyoTijQl0e/m
C14TQ1D7ZJFCHUTMlo41djK6fD3Mlia/g7ifUrtE/eKfcg1eBdBBU1tprU3GtTL9d/9YuSggK66o
x9znb8KGS5k8jxRyDwWFg4oWbr2q00PRkBNmWsq2uFjtHA/6og8pF5XPnIIbbYOQeV6HPe4YTev/
856JGe46nZQTo2ToLkSKOBKJQR8VveJOJ5vTgvEACatc1e5w2ti8A7o8VrR7Kp3EvbFlplKYDBts
bw+NR/DaCs8iAWvH32odgVNCJEdZM/lTSTZ1BmVmdnewgqwe0m87hjqZ/xn2zgAbAcdwwEw6mHvD
ejW70DyZMHY2IoKypv0Kpn9Yht03t7Scx5R3JGmLG3Gw4M84IYyj3hL8ZzdN8XrAGVMyIOJ/Q1Ck
coQjH/xqvWhOJvZnEE/506DJPeYdjoL0Y2QCILSpRFoBF0CahqT0zH922A/Jxy3aW2QaTtR4l/r3
t+uHjHsNl39j8wLlhMIsF+7Nb0Vn+tWtq6kEf3cZsfhi7KTaojOHJgWSH50QUYdFYmvKcBswyTXc
NxlMdJQP7GC7PQRdy3Vif+ie+5JVd0y06fC9Sa94Vm9tw1Y6hD78NZCx7CgVNjWwageg6vsS2dhd
061KNHMs7SNR7QomuPl9rotUh5pYrznIMABHHhmlTbZXYvHLx43Aa2AK/B++oGapU6IGl8xmDvjl
Xv330dLHyy8tJwp6zAq4Qmvu3vm+8V+RpaDLoLIJ3vyxcBZJWLtpocOKhqK4qpsf5P0FQCTQFeTN
wsLdosTF8+BRU/f/yoeJESMTA+t4YnH5KLLb49I6SoHgEp7We9sqTz5po67vBZMSNeunzTiCAme6
URHKYJcJDUPZOS1c1i7NlSs1ejwsNtk8JoFPy7w5rOWxl7qU2St4RXM6FEMQCcfGCwOb23mEBcpZ
rLimabeapW3oboJNFl3HkZ+/Si8tSRr9XrLzqI5Eg3Sm1W7uoDedxMxfI13m3YWZra66WWwHtDdb
5qNj99d9d8lwSznJniO1gKEuU2PGe8rFJwRzUkl1MT6XPL4ID1SnD3bE08cizNkCNAs3dCIiKcXo
/nSUMva/eeEsXoVF2tKUs5eYHF54ftwM9kBzNUBnfy/V8dknQOVx9jsoE36xAL+AkU7iBtHw8TjN
acqxf8f1Kh7bvjO4oqRgZP6zOTu2YSqR1BC/etKWFZD070w1/xvrfvAugIdGhtLVaz28FOJ26Z4Q
yaSOuJIooIr0h7R9+jAUMcqviDnNgSSvBbvJ9CVm8yKVnKfaMwoVTPoQ5ephOQyrztbpnE//2UDq
s6u2hWHAbKp26nHqwaUnICAJ25MuVG2HIsZJIie79BG2ApUEFeWA4qJTzRq+Z4dloGV/lQIxyJKf
MjUg2xrymDr+A2dNS0F64cO8zLBSgcW3lHUESEVgifO9kaNK+LngvJoAvB/yNPvMnZQsQrKMO3Tk
ykFRpHfy8Nn0Z1R4yTS8aqq/Ynzr2dSv3KrCM4kdAdhxdQfovfRUypjrcmE2OGWhrsx+l1fUsMsE
HVNv0RIicD4DDVvLbe/5sKMWeJT21TE8du+KJdxra1P8DbANMscxCNLsyovZcDQhPlsoloM9XdQh
DX0PVo3poUmeVkaJGjnCnbq/EqluRV7hxIoT9RgezlzsGzLUjw9cBq+CSMsAjPHAp/hasOHNoO3f
qYyLZL+XHuaSnDVNr6KamMlw2JogqiNnIFmRkvo00q7OA1LcL5zYABqbeN4IPfFs2KJQj+i09NL0
tBk87i80dCLujci3z0UYDmqCfMp4FWW9amcRPomIUOhqUlP/+W7XbeAe0rf7KA/XbJ4BgWnqNaA+
JTohfLZHhhpYyWfEP+aNpxK090rgIc8JPC8FSTOJvEbeusXCzpF1bw6j4nQ6f53PvOnBTC2yjr77
RF0Q+9RCCU0DSZQ8MZUsCz8JsZwixAziDvdSZE7/VZ7LQSpveWb4F76WhBtkgiXog8eJl4HRJGMj
2ZfoKoCg9YmweZKFm4jtiiSyLXOZ9CLhe4HZvDtoJCGjlmrSnhA5lSYGDL3zsNcd+4g6jefbY1Qf
oqVjgQ/jyV+qNTpO0pkJLweM6Na7Plv42xI4aq3rhkF7QwHGqUBcVQxbH7j3It59JwTWHhLCKhJQ
7SdB3mv4meJSuH9AyU5rU76ka12TRUiD7UkZJ90GdApRJPF2HfVfs+Y4LlV7mIbTOV55mJPuK/Tj
wCfBtmT2iIBsPacznsjx/UNF8RzSXJDAwLVWWpeiXmSg9tKt73xjeEKvQJ3h5G2c9aNUG7agXBkb
SDvoCFwg9090OQBqZpwqWDFdJxBz/OBjR+ygRibcR2sCxDuLHoLco5xyfqs3tOqT9bdEGsO9X9bA
fsqxQ9qQeOcU0SSzQTZebGScS3EZ6CWIx8op1iFYsZ6PkXCmNjuHvI8G96339hk9hEDxC1XWdZ5X
1cOHQ4zuRSPhEWFUWitEFBd5rr7UdlGXrTRLU7W7CNzAupxoqbcK8WPcizK/Qs/Dr+LNBd+sCVVu
+rnVx12TPKQFCr1BXO2JYjv8n3MKSa1skZNg9gEpo7SVXqQOBHdxil6uePNTeLc5Q1+Mj//ffzpW
QyaIgDteWVXqnBdADcYtm2gk87uAz9JD/9JOf1CLySU0EcyWt1eK9rCjj30QaitCvtkZVUAXrZjP
xdjTSOwKlTmU+LDwrThFqwebQG/jTixri7UAiorCxEeLlnBzr8UgFhoW2jpfAOYJjdiGQ6kCgjTE
PRyn/8KYl0iUDGzyc9uThb7l+jrwcfWM0pX5UMiPoWnGxKz5nbB1cuqLu4npIiR7xXFf/CDNPPlm
K8jvLabhGfQtSFjzeT895l75xIksTWqLE6QHI7DY2VfqHY4hS4PT4A8eOyrk4rtJUR2Yb5t2RonE
/JDUgivc5ZBlOt3IiKH5x0dRD2Aem+OvimXFJqTrquEXJHr1+44XF6wzcWb1zRd2WLCEyTDgNkyA
Xnkc/XJ1i1zIDVt4wRVYnff7wb7nbTNkc4qj/GceeLpG+d0f3KH85IVRMMnnm5JwVdRIaPlFO6qm
ZJLa/4wp+j0RquoSyhf6iadzdSMBWwgSy3UUggQyBLatmh7FHEI2BajqQboPkYdm7lHx9iLMoaCq
wNS3Um8R6DX+eebse5qvLkQTySQHbG8AppbUHsFpa4bUW1puKiEUZKlWch42AzN99EsSVTEEYf4j
v9/G/4uUn0thpqFlkzyxFublq4MmHfay7EywamYg3vwUWF3SJRmxoH7MpMWYqy0lnrdefkGChE+E
1gWyGmissDxBpNL8BofaPlnKHqxzwHWev6mzqS/Lezg+BmGB0o+0Ueiie5j3dY9vd4Vw8Qslf2Es
2qpgHCU0yYO/1mTN0ox4iGPMQ61pFwmwKGvwuiVyT4IJBowRrihhJ27otVp40rdeBXOEJ4eX8e6i
nXFNNfBy/q1rBW4T7eoRXDc29Xr+kY8V4UfAMYV6VahVdLZU3M8rjbqNFAppF5Q3OvEaMTgYHlCS
O8KlZ3O8lFDgm9xabGoxjsFUwB4JRaGYuZqYmhwyd4sb0WWtlSmxcIKKB9RmrxMLinRowaK1X3ew
gc648OpK1+W1WOZVCEAjv4Wgh+fjTTOO3lfvCHy6LV6IFcuClXAnsmJ6+Qq+stOGmAsu8JrKzhhx
w3UWY5/Tu2y5az9SnWjWOO3/Kv1/2Xfk2mJ7q+Uy5GD90iAT4eeOd54P4lKpw04WspMYHTIfo/7N
PSTylmbeNciwHqXadVKYc0BaMkTyTwhS99pOQ2029OB8vYP37R3JRvVyouP8IxgbXk+LelrQw+hu
L/AvQ4QD4IDvLn2zFqQfT2ocUlBJb9JCTmKA4xvgBUWY8PPa+vZhsF4m+2COSkgU/aVQmV3mhQtN
gjFiIo3vq6dNen1SifraiZWyed7dn4OA3sHhwEYnmqZ/jXznho0+LFNaoxT/g47ykqAu+PiAoDHn
ZxMHgHvUAKJxyN7qdGNdqpX5meHnmRQBNHQ9rfYuW1JUzSpTPRV9CMS77dNSoZtag0EK/SSMvBmJ
rzF2myQRw7PEwyLWK1h5YoUvWQuh50XYp0xKW+9iAMxhIkKVGysYKIU86smX42rxQV4Nepzfbyk9
QHGtdz3PsrT9Ngmtxy7p8tFTADstI44h2TJFyxMjr3Oy/8yuqSMmVo+SNRZu9dBJSHSQ3RVI8Y7j
VWKWOiKsdOZ0vLYkVTpdIY+mrF9Aw2Yaa78tpI3F3abeLiIOwKFxtCY5NXWaGWnjUK8Kyl/v5FdB
IM+bBntm+/VAN3Pc+cV81W9d6EcWS72OirffLuknesENV4nVYk5pbwv+f93HECbX25qOkLxqjP44
EWLOA6DvmRtO2Zptn4pQPgvjE/5X8OdEkUw1h+flL3VZLBreV3V/abQnNTzqmpu8xNOEYI5x72jF
LaRgTQXAdlogl1Rch98ZfAPvGbMdiivJXlhVJU/jYHU/wFGa381Ebb+kKVPOvdMzeXqlae5LqT9/
2m5cLQxfMt9XTNYT/HiAnpOtd6tQVDaez5DiI6lsFOTJKsQQXCZmn6qdDFAatdSpgoOWwJ0Cf6Rz
IIAGamXaLHUGxBz56Imakcqup8G1IxVV2bwvXVkCy2WKzMDGBkL+rGrQCmP2o1Zn9CEJl+/jULyl
wFvO55NijBEGItaqv1GCAm7ocrYJEZPGm0SZUFI6EegQ+ZcjOWNIOdc5Z4S4a1IIHLhVDk0ABJH2
ZpYab/K2G55WPknY/XECVky5H6cH2MDcIZCiBPCuNZ0MHxYwZ9H+Yx1gdT/FK25x32isuWwa7WZS
rUuqLMReBEc+KZL7NM1Npc5527AMcDgVFDdIG3v0rq9Pqq1dZ1TjXcgt0hOc+eRFuSX/GMLs8wWe
+KCpIFMsTO08aDNmZ84TYEaoIBy472CQx/9BM/prQFR/9hyHXJRt8Rye0fqbim5Kt99EpqD3YZ4e
v7912ApOJBPKZyhCfeUSLnhwyStEZaZ/yeHFLiUiYke4ylOjF+q5AzoHzze3UaNhQrAXaUHUMEEi
zYON1UL8Lir1jUKQpQCE+SallrjCNJG/jYdYLuzbhpGlKhuReCCNdPJpsPmv6q2eQ9XDAOYvvu9h
lxb3ZZ7ew2Gm6mYQQECldi3dJ1zqlmsQ/Tbcm71eoWPJJjcvnbkTNonYB9efDnMhP955uMUkWeRu
1YpwBs4QTTWsc/mjSojg8aRVXFX3ZlwAZKGqLtGHrapcRCWUyC+lrAKAUrzDfvJmqJx9f0ExMYv7
l+qDFOPsyi9eBeLxgcKXGnq6F5fbi3T60ajeFMhkw14ElHzuEaSHBAUWXHncO/MFDh7FpDRvgsp/
WMycHzAra0E+cBy/XpyHUl3ER9yRiGIt/k+TI3w3iuA12P6J48rglhrR+1ui1QHDoO3yIr1ROV2c
VM3uYkR8MlXYgFj2TwBjfFlhaKLtqrZC3qo+UnImfasRW98IQD9QheZ17yckL3DfYdkw4UPiZvB2
WkOfCSRxxJ7envp6wyFN02WZFt+0xFIdwt3cRwz+QnOgJmQdwR/+b0gwnenhVMHw/cOiTHgaqXl9
CorVAy2jZ/dStTwlEgr9YgI5/Nk4UwC8LkatFws3yH29eyV1holyoNggpI3grHqFLdsVutl1Kx5n
+b3wLuo4CKCg033p9Qsqrjx9MPMyqnNV1cpvzvAFVN+lob3IRo3X/Mg1VRzuu1AVdwOu9T1l40XW
v+hMNumAYdrbdtiwGqgvxzxx3/lESLHmd+jalGj3hXO/h9aBHhmWr4QYM2hoYJHfAEByPCqqRRSp
EtX+xFc2L99RtVOnWGaAnnuSZlqFTdBAyH5+AWtCFOGtvk0vknjM5KNGGkFybE0ohV9l9szuiYsP
81fjo9MC9Um1Qb108TxqNEnvKOGkqHiqeEmHvBPcIqk2lG9KPYGjnQVYE9oF9w8r/r1sD3ULQ2u6
IhBsP0JGJe+JbNC+V6XdqT+R2FntKMwl+FmvC29EubpdZ9X5EoRDs/HMUBBf5eFZEzG7If390hPm
Q3qDMW02qZV4P9gm0f8A2B39r0uc8XGbzbm2lY4ase+IxDGHB/IixJGxOZk3H+36qO7YB8bdshjo
aeIhDhtB2L2/xHn4YyDXOLtTlWGmqPG6vymlEHvxDVSBsIZT1qcn+cfJK+1k9bu6imSQ0PkzwIwV
wo7XEc5Kp3eS1brFoEXP5QR4LsmkHSJGJESS2M6/h8KoVht6WGLPUZocyMQnk0eN1zN6tXAHwoIx
zNF8cqxzSxnPlCq1nUm79j5VfmKZk/0Peiya1xGSFT6/bhYZbpsiNqbfd3XO2LZ2DPVcKSwayQE8
sU53Q+7OSjCCPkg/P9U+l7kEwcg4x/ymn6OJMRKgTK/UExVt0EjPR/eo+9m+azHNXOURrZVBqzxq
pI0iXYcmjJp4hwtxSwsVmA9RUsGaU65yiyw8bnLwKWIH8gaGLTRE9ZS5QiW0xqqUp/IxC72eCydU
PAqLnwVsKqyI/jhaaslU1G8iKWyLWflvJ2hdqz7oqxwu93pesk2MOMgbeGjchK5S7g1KvxhfJQgU
cN0I7Bl4LcSDCxG+8BJuv+39CP94fWTxm5gukMoEPXCiqkKWkFS2EDEOK8LyDx2WoJcjwb4AGBM+
ySL1uX3VZE8oP17wQI5SIIDvU0HeFEDYrikqInaaSyMB7tLGkPv/YIfTc1/tUR0zwIJ7YRMYbVae
1YL0xPUXyv8emK8d99n6sbiWe+ACaCUp8k5dHpMFdVq55/trhajPid2oqSSCcTKMgJKSTRvuQ6nb
wW4sRky1kbunq4TqO0wDXzUaacP9q7c3KilqHeO93E5j5A+oxW8d+22sNBCmGl8VrMLAfbDCzSg9
0UX1we0H0K9+m0WXVmgeYWDhazUX1jCCWHaoQrDR/RFG5rHZVbZQMrR1Tfoc4G9bNL/n4K4BRZ91
OOUBlVtrea7FrgJaYKSZjVUiOcFEu23EU88r2yMFSz8v36vd0S+PWNW2hHnZs8oFb6F8NnVXu5CI
WGJUNpoPT9MVy512AMlt9iWEjShxYAhW6FwAxI6aU3gFhYMYuMO3DNt1YfJ87q0aFCXD5aMRvVt+
XeFpzSZmOtK7oPwLhmTFAc7xScGo+bHRD3qBb5eMYAKxGJtF9OVbMJpjsJMXXlH1A8aTW15+dVY6
y2bxf5iPvBkPrCSBj7+camlhQK3ANN5yYO5EvEFTgRgasy9sxRR1DqEOnioSwuve/eCyL3dm+2wv
W959shTiabqDNlgMbz+NMQd0m7CT+ZQU66In8LPOXQLRB3cyDPvme+GuUKzrtDyycL5QRRaxdbvW
jo1NHWzEXXxh47SOOEV8kx0/GyNlTdsCMO1cmIZ56SXI3+4al5d1uiFCwEMjhavUruWi/4UxbM2i
UwrXkVFShuDDuRwdflGxX75TKwiuAIa87vyv2oESkPtSzQxeQi577n8DqKrxvU8R5I163c3/xhiM
k/0Abr92HMIVCFGoGGW3ocMdQzhPN5htG4nmqYVl8xcDGD/2bIqCBnQldh76ofq+HJ4rHOzUgunb
ZsTYk6KUNwKOU2tT6LSw0rqjm9+cDhWVKjLP1Ur9JfEj88x+xFXAuUjOU/MzLUeh2QwPZhiuUxvG
Rg2Y7+F6WYwt8FN3pbVVt8eHq/o2aBU1dBIzHtH7KLXDa4gxs/bayzgcJoGXygbJE59xILnt1Sg8
Ng4KzE40bwVoQO6m3pAfwia31TTfRIWVWeF7P4gDSbFryTC+uJiBw6mpIopmONP3NsE9fhmjVZln
hNK40Nyms3drbyGqKA09NZz0GuRg4jo1WsBxCZ1HIn/0M5Bj20WCSQDOaF4e0EH03M87i9b7Afj1
uVaD7Ut/IMMIZRkuXjr3D/Pa8aKGYOda1O4jJLD0llBVmH3OKZLXrQL24p3oDrTleFv7dC5XJRPV
UEdrkQTaRdK/wDPW++LObh/YEfmG8R8ECn7xfRYA7mXAUuT+kyTqNJ22TuxLTVAeMYKP8vMQydCm
qkkbxpCE/lKMgevfq4+VJUIJP+poBXbAdXhRVTOd2vvd9MxMHiRTKwLKQKebyvbXmNl32xwgoEOp
p+XbzDwOQFfBfRNYgZL7uLXU0e7B3zflTP2+J8PCYPgsFRHYldhXGXuGDlLbl1PZWISEqDihOZG4
Y2j/fmhuFPBxhMWo8p080GaKMxJnK4D3eUlCV2/9sVNFRW9h8bhP6LVNm9XuwL+ync6F2NCA8nKX
BZn/d+3uZwd2+q6qwi4wFB1/auOEbzqD9GlckQ1ibS4NWtVPuqg2WTCJbpAFLOpHRaWvMLfvgxGr
fIVK5RJdZemeLcLRglAyl3WYFHmESEbcImCaQCh4Z7ooBOXINhz2mgnFl428LMnJVgRsXbNEXRrJ
hry/z+OAcK5DRQCtdIKHW1+aZ1xrvwOjULZ0mHZJ8l+zY60y+rcyVV1mCioZXaE4/SZuqNCaisad
tKlj6Ehf+GTZLbbVkk7qHk+4jtv0oxL+K9vJPLFP164E8yvePiwr4aXqlMMbd+tDc0+VvZt7GxKD
Sd791+NPzyAAZ+02p2QJ/s7/YEZBB1tisz+aznibUrJDTVL4WTloEkTIcUaHzRq4IGalTJOirnGC
lRbIEYWu1EDTAlJY59Hj2UmVfMxXuH99NAkitD0829almXa8kkAJxCkm1GT37Gid4VHNs+1wYYEZ
NmFaeY24S8kLNrJ4SuXh5Iy0pcXqKJFF/wDp5eNuSxq9HnpOUL1bfqvqRNSx8GAhASMXG39d+THy
RIka3TJFK3JEMyTB3+yh5F7WGU85CW24BwER+HNO06vLklqWXs7M30x/XrGRzy/hjEsJiEJH3Xyp
ixF7+gIuDe2CTVwtke0D9Y8gde4WWPxR2D26BRGUDyRWRTyrPKeDiEL8wyoUipCgiGkG3uobNsOy
aUwz7fk1ekHOQzmLznxq+ZlgJeZClHJWj1B2ICShxaFdfcTJz8AbLI4FgqBB5wqV5b+p2a8l6k2V
bXVPKjmv0ejB/8jctkcJ9Jn3DKhhFYhVyQaoUcGEHmPL7dTDJSttUvzILP637HbnclATPNPP1zgc
g+Z9uWPb3mdyPB7RKAgAFexPHAgdDrbX8pe+ckEVFviE9l4sWOAXWPPol6jikJdesMzaXoRPSmJS
ZI5rXnUA9vxRjihdjfPvRHw2rdK1HF2xaUbvGFedTv3ZnBNt1f8RwyzV/5qSWfQti0DNmt8ZPvZ9
CjzQ74ee9cTaLe6U5e8liRJg1qHKfMdYCnmmRTWDs+xMYiaMy5h4JW8QXXf3HwLDim7AZnOTIVx4
N6nwpRmMgxaEVnuIm116jhhFPAR9ezqoKfadGcP9UmBvbhiOyjzVH/bzto+mG9r3IiGJy5emSYO4
Q4ehM1vxksU9MptcJizUo5Iixq0VLrL/iwxmQIFJa0hAqxW0oCZeammR+kEk+vLfpBs43QSXSgLm
GksXtQqT35+dZ16HcI0ASI0vgNAnEpqFvF4bkEvcZxPqOJFDgBRD9lnzUM+33FON8pNBvPdPDKWb
LAm3wxbzI6VXCVkDA4ApGisMTbsWzFShSUGW64oDl+/uGceZuDUkFeeHcniMN+y906Qd1LrZXuiq
xSvnP0JWWBa7DxQgq1GXAToYD/+xJ+oPdm5mmYTb5/nfjSe5maOFlVS3YsdIxVLffrkO+7qyzw0T
oDb0WYFw+FpNXKzTRQen/jZPEcxiwSOx0FA/ZjHZpAiX/ypehcNy5CKEkpJLLSggjp04XqJzSa/O
j+yrGKjYXseQCkIvuaMwgDJF0qPDo2wmmMfi5ulP1V6hIw0Pn1sXS4iuJqJCWNRCdH9AHemC8hbs
ruIgbwETDmPNotg4+l8v8PRcNRVWRwI1ITNtAj3brT0CcW+moRfk6totLTpaXYrlsS47Yl7TtQ/G
MQQiHKLVnGq/xdx9wVBLBkHZIS4uZP2Ny+tAn62taUoh0DQpiODp90E122pKzzWna9QndI8m8X5x
fDG27iZRchNSzWu6Y3Y6ZYqbglrLbS29HQplKfHzbZncI2ialz+fTxBXcArXG6jEeiUKgW9LwLJV
WGC/+D1LgKdklfFEw3kD9nG8e1UmGNoZxGGJXMM7dU/WnnYCPsbOAgobiiDBG0+4nQ+eQCWgZ4mM
v2d8wXAQwhfw5VJ/Wgv0fbuFlsGdmPD1uhVmBeiG0kqDlO8wcHOsbn+YQtyCm0fPAfRnmXMn0NdZ
dkfLrczx7MI1izQ92n7l9DmUtZuVlIzHx9lMgt2nhat3XYnjRI9z/bUFWarUmUDYdIg8xKRgfpKP
BeMhyFOxlnC2qWdTWyqIK0VP+Ps9xebvoZ1Ef05zaQ6xmApd7RRoKBE4XiT3bCr7DUPJ/2GZ9XWp
aztx+NSn95xCyEv4NmvFaM6oeKFuKotEQd+fL22Oj0fjeJliOnpW05QBpddR7hcrzqUlanhJFnoD
sRNvl398t+jdyF8b3hscJGRpxQ3AxoQ3UABAiySCrC4NGspsXGvfnS+RxxafPxkTj8sQbTScFlZ2
UijNTAWRoSlmwSOVxnA+ZSGj/0unmFJ4JOw7Izer1/4cDfBoJjqEP98cAY/PuAti0fdy8+wWtoZi
mojrHVoIZ+0k7dO/iw52jYYoXQO2ofoPL983hqCmKZnwUbDCbqbZgoX2eaf4QDAu4SD164CgYBX2
dqmGqHJ48iFu9QDYZ38kSQUdpIP8RT7UiG/GvlQEgDg/qxdUWeckoKCXPI3wDyp4kr0/5WF4eehp
LB8UC/iTQhSpahNFxZfN2BjFrtzuz53jqXt93/hCgQimdosYTuBnH/i55gVm0Dsl5GIp6T45d/rj
SUS04hc6MopT6OAWjDbGD5FGza6zmt903/4h65lISfWVv3iTRlKI72jjT5la35nBWxb56uGqc/1n
fA1RkAtv277FiqtbiRymIQv5KMu10CNE1rnktmZ2CgP7u8whhEMstGC46mEP/SRdkqLS/dT8WXBz
jZCOJEGcopCDhdMxQoE0yB7oG7t3a3O6LOvZa8HkllvpohAzikA37+xt7CXrBNThA6NNUGZOUF3z
NkikQfL01HrkBvUVSELhUZ9slO20npS1Sy9tAUH2h37nlkqj0c9nMNnHufqA+ziQFugot+WwfDzo
euxc6w5NwC7RXWT4X05TPrSmj51mvA14HCKPJB7IkaFcf8cX3FoSYqbwIho1Hfg/Z1iBleY+qpyD
gWHRw+uH25+Xy34DeBcaeRjhhB7Y2rYq6BBzTghhSHOmBNCfJwBnVf23saqK/Vcbk5RvOBCXfS1H
ZeZ7Hzmxt86NbAJrNRLy31eQ9Ya/Dqggx4mwXiXSVa6H0nqIgTxk41C1RKJVh/YBh7kQfbvAjqIs
rz8HX2AoXptXRgUm8OHnHt5zzrpOhgZmPiloZfpP87pKHuC+6NTKjl7/0xm07e9l0nsOBX8yfBcl
l7ZNSWJeYMJkwETM898Z47+42x0RdHdGAiO5c7ta24wI+Agy6Fmxpi5rxr6w/OWXXu/6C2x9eFJ7
W/g1qZd7rcr/UIy0h3LTKT4BYMYluM9ynbz6q4ZNRBdLiVQlytzZlLGkn6MWJcJ1zug0Aj1ohWj7
al6MxVj5CJPZsplBlXfPzSXQP/+R1sJyiRExYDamMsoir9JNCPQEcssvfczWxLSTNytKkt1zh4+D
ShxktwRD+jFMOhV+qviVUs0kouwJcqRhxOpRzk7LXRJOzfKK282fgA8BCJNmKbd7zwEakdXkmtaP
3hxXIO69oFFw+mpgdQ+VQSF4F2HXqGSwO+DMPznMXmA97ChJAv6BYBxzX1/o+cdFWSaA0/hkmDTy
Q+hnvbJmUKetzZSLCyLKjSwCQmYC5Ot922ThBqmoFJ0ChnUdNrtDkvDbMlqNNm8GZ7eRDigKWpED
eC++BH7MHAuunagVQkGME9XtzV5HfbgUBWBXL923h6oBGl16tlz22ExGmZlffd5M+PfF6ACwl1/x
vnKLY+KAVdQs0yyC3WcpunAEW9xM5G8sANCS1SIAsXD9r/EuXJughilbNMq9F8TyrVTH1wl7dGG8
tUGUOJ0HGUtWZUK7a77+3rp6wM0gbjpNhXKSkor+dMpJb735Q6jSwHAwOZrg62672Gq72LINeGxU
7INIIHGZ3301teNnn7fXSY2205LbHZYawrRrP6aKYNzLp+8ykHB6QONu4p0hdptv7qGkgv0R9e2W
R3H4jeytin+BBw4LuF/76s0bDe0zr7I33RNS38jyh1FDGygDta4oAaJKHw+7Tq94dH8l4nB6sDBx
DI3DzDPTt9tMz6ebqZP7iFlWZRQZ9XxVQ6att0UJCxMdObN+vVKviDNH8p0pznLxYlOLmoVmMTyU
SnoAs/Z4l6zbBin/kB+uePgFh0yBdc8HWsmFg6Bgla6gJnq9s+4efa2lidE3znE/FDSCv0Bhe/oF
tCvePnem8ZRftm3g0VuFXFTp0Ng4+IYaNwoZn+bNvtmqMLqF429r93HDPtIatpSVPTnvg759j3BS
0vd1PqvnkRK3RNQVU+g4An+2LTetTuiI1KxHp/mKfGydJ9bQuKFtgH2aEQZ0rj9Tyff4gWAVqDl9
OlLbK+KdJyemcQbog2jI33YpLibwyPcasxods6zUBYKbBR/gf0R2wOxEy/filN81o9FCQsHgMt4B
GXordkMlE/fm915e4kH5Nd+QdsGhR10PdSKUZmPDHhDRaJhvE2/1cV330JzUjf8spMtUnxfJmtd9
lrSU6UG7vBcTTW/EpO0OaGJJzCF6gIs5gQSqQRYiAaj/mm000NJkJj/0AMP4+DbZgBy9Znihp1vu
KOSF44jN1WZTPBDUtrQc8fpnBF8PexocsrRCTPGhd0xJtP4qYn4WalSX4q9KUGZqDzA4YRIL3+TA
xekqZ+kFbaUTEMhMZeJI/v466D5jb2S6JcRD7zVG5K8aYq4knlggGuYNf8PPkG01vemH3VrwsPfM
dufUIXkmYZEDo6ZiMNZgh3j7WaLSl/8To8eCT1xgUhrg1rpEj6dfW0tlxtKHlmGjIefIl2xIAuZ8
HYXQkNv9ROyWLwGv3TP7YaA+qYe8r7o8zMTTyI+7GaeVkb8+L3Cxawc/xMPiDe04WsuzB0eH5+1h
1AD+qvgBbWARW43zWpTA9huvM0I0GAebVmgWReWucUC7eqY2rlyme7oupXdYcTazfeFynwrdD0Qj
uIdGKlYmtdZ7U3XK+KhBRX0KyBaBFQGoCEhXeo+ZOzPR/OK2UMxkaDRRlUzKXMNjrBP36iXJyoyA
tIR/8dNsIVqEkcIP0fv7f5G2Z0avNSI7ZqWu2RyTq1alfKeEjcY70Y9BqoWOal54ETZlMQCKkKFC
wXHkil8qJr26Y0c4IcHJBsApxQilh3N6fia03lf5mXAuKlUaQrXC4bMZan9H/XJkft2QyvQ/1zR9
kPkNgrhgYehjLuzHa7UCZFCsrU1qRQk4d0My/LobD5drstdxv95HsbnWlNhUtoRQmcb0fekflTP+
otDP8Som25QO3Eyei6BMH+L4DtHrgAgTiQiCwkH6I0xbKyMWF1GFMi9FQdBCk6UE+oFAFDnVGchV
P/AgKoMGEsUiAT0YAWx/T1tESCUAEykgMRTsWDhnvczowLjArvogF/OMU/SO5le2nJT4CRt87zID
rbYvjyF3fDYMT5JPea3xW3JtfWSt1zd0AWKuHdQTYjdrjQYUQEioObSRhC8shMcHrIpOUeaOONCj
sRRd23CT/AEYizoJLgqVEXDmkm3/f0knNEkVpbUNeOZzpf6PJkWR0k8xtZ1S6jIBctaKXURvSOPH
9lg0fg0x8Ma8J9olj5ooewwyunaYU9Vg54UWOzbjZWL9vjmQQecUgZrh04MehyvLuY5RH9Mw2BRb
bbWmyGCTHTiCffm6Z2tYvgMO2fz8+ql+cwM2KnabcUnfJ6JHeLABNNg2YBaW/0i5kQ46CZracp6H
MtiyMq6TnSDCO3Z5gCbWOZ0CBb8Ifr5LNnv1Hs/3Vh5rf1xED87iD4I9KJpedz2WNPjkj7jOFOz3
PxgJmGXuNzWm2JPRuGf0iaWwfq3QPFKvFvdUQfh/LnfOnEGVYB9AwNiZSkdcjcyr8RI4h7mEG4oS
+wky614Xr3uD0p7pajUg+UpgV31Q9WUyzMVgwp1Kgw+HcpPgdguB7WSLV/BI6SUEg/GrRn6nPfn/
kSusz/nrvmSkdzjdqOeEG368jY1yuwExAamWk+sLw3UtNsAyb2p+JJkPqbc/jq0cSgWHyV2DyOGY
RjxxkPFL1nzZ3+Q5XaxocEaogE1rlStj6IE8KB0WJx7LJUtD2d5kzw9Kf6R90WxRQ5v37iefbofx
dPopzYbl2rbQqfaPTMKtT8uGxZ60vZ2X4zpPrv/W2pI8DdOJit5R7TV4rQ0Iopg9WHdGbdAIMNOi
jMaypeGvKcQO21wHNOF4405LJRWndA6Yb786VJV4qcdc5c3+J/e9XHA/Sj0PUjm6tSnmkDgb9ovj
AjBRfthDlf7zMgK24edSoDKhRifRuKJvk65F3LI+sc0cN1UCZSRtYLljzKnSSEouxX8bpBtZVtzy
uS4eUy0FoK9oFW6nxIeR22lUKBK2/ESNVSaYcrOa4vj1b1ld+ebj+fWnVqlWVOHycvr5AqnOyi4N
k8YILQLGYHdeKHYW3NDMa/gqH1m/PDiIAsFp3BQLBsWNaMLvL5Y0uc4aDs39/zGsplaUSoo07hrL
9amnl/UGvnmRGGuBHoZXff9mt68K0mb2G8t1zy73qgvvlrb3FR9r3TJd9EYqaQq/1qh/G6s+tPzu
jojETczG+Xroepk7TQV9Ia/ShvmUpTMhK6d0cOnX1okFKks6+IU0S5Er+laDkSxJ1Y3xa9R4MfZY
a+N7cDjip5nQrQ9RqhHV31hYUU/wRbVqku4UwTHmzftCyHblZYCMPzv8/IBR0lLv+DIIoldZYs8C
anwCY9X3pICVpi9dWHF8/oET06JfhlhxXPXSmDaak6NWUM1rQXM9FIS+OVWT+T5hUheUCx1X2mW+
BJLtsLSyMRRul42AiljlRV14lRkcn6FPJmrgx5BDoL/USn0oulyXt4XiESeu+/m0S64oJTgF+HQd
19HKdkh+8c+O87I1ESmdVKj22iR+J0WolbzAjkKyl9XvkPDmKuoI66Dhyarx/B1ruULDMang8FBx
pNJ0Ra8LnNR4KjngVlVKpj3Ngo03WK0yq2Xhlgd8C1fOu7JfBoIJ312ZopL3IfPuCYxSwKFV+eAL
oSTav0ws4a6SdXHKmDYK6VMUI3S19ooxFvv6s6esSYii9ss91IHt0uCJ3Y7qrpTbnKClQmzIUUXe
F5NRarp85y4Stj5cs7rYhkt+mfFPJtWgaek0D6ZjJ1hgKEj/pqLxYzuhoKGg8WXBoTzKVo3rHdDH
iKaPRsGAK06FMICPoc5QxggzOQAjPZfAun2j7XObrMlXM3fRq0k61y84xNds9MT9IVLi9PtevDCp
mrM6eXFTPVUvK3XyQF/oWQXXJ20/wxBettu5p2FuMX+fsE+3X6sePu05tkiN0/rIxZixGG0HvlpN
028bpoBa6ho5/RaIGE8Mh+UJYnySQ1e3jJVPY/ambDlrchRgdZe54x28EvusrRp0sEMUfPdTzEPW
nFVtHYQdtdtZB6AQ6hTgPIH8xmiBhHcB27ONA5oFmymRmXhIzBiqxjHJ4gzMukhEYkR8utKAff4K
20zTRWu4LLes7PGKue12iCaFatNHhsFi9qpTxd5JgqVSbT+mWGaAWw6jR0JQm4fb8LTtAsK8Lyu9
6NbeSaWcypoJFigYT0+ZAdFXfPBbZws4wKc8McbhyjO6IawSVVSnim0DLAEInCyMV90RS434BZAU
bE8xyxeqYfHa8+m2nXfQDh84Dmg5yi9tc6E7DXtNqaA3ohu7/rN+XN5BxeDfNwVn5QG/Qzi46cSI
QVVuinJYqbZeyWAulcBds1dbGi8DWcL99wEqsxNQRfMfveZ72klbTQ3LXJR/ikMj75qFgBHuAxib
4oHl0Z+rU4lxOD93OBeGZLAJzmpomtLdIQwapV2Bx+NjCt/XM+lCnA0WuQLcW7sXB9hEPLfR01T2
MEXAF3Bo1TV2+iu4qhQdZAdW6bxwWWXnn+rxnS2fVlVZM3oNw8PEpdmPMiFehqU07Ux2HFXGVCvu
iozOO50B4nwdiWXcUzAC5qbPGHhc43m1s1rJO8gFki4iPakyMIcdzAdkrYY1ToRw4zAMvYPsM/Tw
7H9zJRdhf8rLnq2Asl5e9eC346yfq7ggGGPLKehmi+YchFViX0F0/zTIPbymQS6QDQXluse8Tn05
WXvMGtvpSfXL+lGMajFjYS/mgxim7taooTgUg22Js0aMEF9lMGO/GxWrHxfC+d/ukxeiPsLeWquT
KhmENrjZJSzKhVDQUZZeCHvoN/iarMHN7ClsYBRwsyaTIH+F/Ud6/RN1imDR+nxIOnyWc67aHD9b
uzey8rgIvNOt1we2Ewaq+yULsJ0b8JMvA8+Sw6LvI3t61iMGUo+yZ8rkR7YUSMDU68C8lGhIRaj2
kcZ6gq9thuE78E7lF65ohvcDRHtUJqdSu0nvnsh5IjETL7itkoBdOIsuplA94elDbP9GIAFQb+jo
FqM2Dkhdf6IF7Kn6BTxw8NXCi1qLPhV2GQP63n7kU4rqoaDBsM8CTidYnvtYAf2pAKod5YgdJika
ZjDcchYcL/d5xcDYR0g5OIkBICRC4RvumUYkieUR+IaLEt8ULh0VG7gFIsYWcvoNxpK3yCHQ0c9v
EoXgnTZ0Zb4PqMiN28ZL4Ow6YlaAjmk59J7Ny99EFvLBoROujpdSmnZ7GdbapPAvXbmM6H/ihjBj
CZqr6+wi1pelE5L6Dx1VH1+pmM2nat53613pVbc/6xY/g6ttSMF3BAEgznuzq72NtZ6/VoVrPdv7
x+NeUICxHpO+G+8UcMq8vrkRNBHrt4f0ljz9+7XWnJjq6BNYTPH5m7i3N7OSawWzhIDvmOwQlRLz
5L6lBFgFsARBREEN5YyD0hNZJu1+G5F5CME4JkFcwuQOjr9zCq+H3QMnmcUPtsqm2ptAyiCkGUzc
zuqrI9u7/hGjoBid1h39qwsi2KwjByZHTXIcL4v5NMU67v7FnThFEvV5METSHKvpiTw3enVsGokt
27++J5VsU+jNOv+e4SfCgSHM3qrPpbwkrIUTeROAz6p+qEH0ksoaesBgCpJbrhuX0HNzX184NnNg
KVdbHzdjoEns6idj+7ZgEmdXYhA8PtJ1STXAybcVUxSkAYwukqy7c8dYPH7jVZvMRdDvfNVTCGFm
wBsTkZGbvvuF+DmlhPeUS5G/16MYDjk6M+QYgLx3d+8swGxms51GOYRcJKCvyyhVqHRCbCYkkCN3
vTQYzNMp1umsHrPvekgug+rGnSGWkTcYKOpbFYJiKzxEJZWLrogda2kCC3Ja0DdXDZuMz2NiAbF6
shDJor4g/Dvr6iTQj5J1t6apsfzNTpqW2CET8B1rC8mKKuyRdAin09vIlg29uDZyQJJAyE4pVInR
0/jsCrap3v+rRPk1tYV8kMThSePL8uuxr0OR64UW++eEyPve9bW6ov9aPQEXgI13KDZ8BeYz3tW9
I0H5mdRniw1TVOYVQ1E277yTAGQoY7Am4d5da3qiskdC5UcvRECitzV+F1cvIowmHpbcQFat7MVC
25YQY8e9mB4ukfVNJVeowYP0rfAyu2FGULuszQSmShNRP9VPwwO/6A4rBAYG7gFWzgFQEIhW1ObY
OXhP7Lkjv7M1X7PLKi+lp1UN7VM3dGiJdOZ6I4EDG1CMpMe0XGlQNAvPDsJtdMKUsBW5i1JbO2MQ
6scPOK6uQBXypUOOTyqWizZNVuu6z6dE7MP1YcoDPvG6ZUPM2ungYvHZ7d0AeI0cYTJMmMC1ZO0Z
wX01CIwuJPOq8Uzug5VX4Mjw9nKHR5Y3gVI1IT7e/jtCv+Ku4HoGoRobJ5IUKTqbrwGtuqk1W8+O
8OqFda5qtPSWG8Iw0DP/W7J9mTo5/f4GpT1QV/MnOu0xPQ6S0ExgzljowxoTJ70HykoyDGHlUBoA
zA9TdAe05JB/qDa9+aNf3NQC+C+oRi4n578VkIXC7dWPKFUvVGyfMiXCUUFtYwXLRerquNoCYQ8d
CR7yQHd90z8j1g/So2GAFoBUxMQoG8yd3JjWn1LW1PuDR562rpT7NQ0Ii69daaobUp44tSrxaZL/
Y7DO2uqjt3E+jCtrPGwucav2HRwuKOkU4Qu9uhIe5XJ9L2fUO0Lowp2X2eS5UhEHol/6fDQpZrOH
Aj6VCdYq4ntM4vo4qEk8jN7CLFlhfz/Sr+Pfy8NzV4oTsmH0qxaQRXgdZchYml9TAwqu0AAA4f00
wWgKUvyTypbWXLy7oS8MwymJ1xLHQ0OQAAZt/PKaxFdiQiO6NZC3GVQFBVWfEDUjJbQKsgSActgj
pnjjB1xJPCSckK2Tyc6/xZsJKLDFDmO8ysV2rxwSxGQCcaJaBJ8xa9ubNLeDS4q5qfo0Q9SwRQUy
lewG0AtddhlqbcRg4wY8IgbOhLKW3/nOu9hH+cDHI86KTBCuUYLenklCC9M8W30KUZe/PCwM+s5Y
WBDQUHgqULtUveVQ6CzGEAfIwGKb4WUPNs0wNj48BOLqFD3y6ucRL8wsIE0/2YKIcC/OvZST7Mmw
eJHW/P0q85EeQ89k/SGQd5C+cPsHK/1ApKlUZovqmEOhJUJfuqIwFI690o16ZdXq8OZmCzXImBsB
xPksma3ON5JO9UL2svsO6E5JcRI7UK95dlOft4JI6o3zFSDYRXEV+rdMJPA1gjyWes8QmwRZUc12
ws6YSsl/KrUOm2Snf1TAdCX8FRjvVVAcuYKbRzq0Z6oLx5ugEQMwGK9sMOBLEjKt5BC//OBSeVKf
XvLUJfOHpq/EeBZhAwCuMmdEgIyJoGQuZIb4kyANgqcb25+armHqPTw8Oya4MtuW1trX7aeX3hrf
k3Jy0pbPqjDISEJXV98GRmifIZ9tQTHbBymBsa9PlyCPEf2tqRx7XUEqVgdIOn8jOnrVELGWbuXv
nuJmwhGQMma34bLayppuALD9XbLrq2aWh+8oEeaTkztM0Ws6k/tlNytB/QdC+XuYkM583GWYmORW
XSmU/qLOPWZnJUkC4UADFEn4lu4MBQc70ZTWyv3cl+wuDgjNCh6rIxO+QSkbnmN/ZHEGiQljG+Hm
+3tXEdV9gqZPXKxXC/i2RA4fmuGLhbXIxNaoNOJlJEyKBggpsXzrM7UbFvx6Af7gkNBnSV3WNyVn
r6+wZIibjS4x2GuAcbP+9wCeUxitazVe0d0Hogr0iPZEuo7P6JhJ7whAOJ1kW+GIvrvP922zMTRT
tn1TTRdCCvmbmOyjPiWwLRw//naBUC8AqXSTJfPObtp/kx8Qgw7r39J0JwZemWM34fNOPtbaJh7Z
Vst5xHK4GUrW6HpiWWScipEUYkdUCfnuLfnRXPhV0XZ7bkB5WFR6MTpj2vFXkTpRjpxpWFOwq3yp
Ed67QN1D/WIWvpeQslZ6AIIxXwGPaz97AueVU3pfit+9KsoHDcJw2qUP4pzWiBDRg2fgPLJh9I6w
JaEHLk2G3ufxn4m8Ae+UfCf6II/yTA1bIQbxF3uV260IJ3z4o9AnV+IjOZ96gCgcPnrjbpOI/CBa
O3orYYHD/fd1ZGA76sG/LumhCGmKRk+LuLFyfe2MgEXQIacmIKIpIZFnwVsAuy06NOTG0lFWIZWv
1Wo3rmuFO3V31trIw55/mZTvUiQpHF3cKaZdQNUdF53DR4E36pULuMn3kXikrkaNUi0HZOLJnswe
h34rPBrLt3zeUwoNPuheriUGQxxGnokYaqERV/e//4XwO0wB2lHJj0+TEfcYEGvOgSs8VvsQdsNG
dC+WFszUCR+zk1dCqkibKqpS9oWiwItTeG71TKImlVz2wPu94w021nTQVt/btobh3ai6OSrfEhwV
rKB/xO97JqcFpCQCoOxF1/sWGz46P0Q4RaoPAiIj12KYQFzNOfveHN/4xOtob90ZGV7sg1l4qli/
mNKAJzOSgo2ZbaLFMkGofJS6iqY/XRTGEplGMXagT4glhHE2MAtnZ5y6ZveOU7/wWAVegbrEbid2
QyO8runR1LgQopBlYmepb/pRnNKnMHkdH84Q47p4ll6mup3rNxlsGmiv4GoNesUuv0gtnGM7G4Vi
LeE7ZHVnJ0k5AFxJZensi2jjpeakSRbiCfrm4T7sA3nui4IHHby3dGN5Fmaj1ZXNDDn0QTnLByyN
GQfWuBIeMPttfMJHGUy+9BJZmTSP1/JQ0F2cG+RXPFNBWPz1JOvKiCi1AYphYM3Zs+9s1D1NfiWR
lM/ghjEDuqC2utHP9jcUxdAEmKbNpPUdVWPhV6fbWTZ3+OWOhx21SRJs6pYectNFLoNeyrCIpmM4
25mLVBu+nVFfEs+QrdI9WaZFo5ewPKJWiA313nwSLerov9wIciBfa5Zx5ROBEXRChBPlD/lUABCT
lwwWXNQ4lhpYQgLKHU881+e6d8hehJxHznNIVSMQ1st+0+RlGR4fd8mmeByCwGyMj/BPjofrKlHs
1AX1X8LvueUYxbVhhuJg5abTY0+2XMT2EOR4NH6H184Fv7YZSgNolGPqaBT4Trrb0nS5K41PkLur
Q2N8TZFLKXrEb777LcsA3k6KJR+dk1sKgkzyozCyR4I/oJnCsM+uO7K6418yyZFoCiGzmZfxdgp8
3vS4hc/xAPe05zRWUGu6AXFa3L7E6KO/aoZI0yI91RN+mdHmE/zqmfU6vya61PrNg1ewds0omj34
iQmb1Um/zpnPJps9Aad5pCFaI4M4IY5pE20UHK6MtuYuaexN0/AGfrW/zWCP4NdmU3UzipB6zIqS
U05uVWTzpR9NuSm6vjlJH6xrolxC3z6kJlUzekyuMXk45jDz+zCjxjkLbSdYwmLcS/uHVuj6GI6w
HBC7CuZS20Ivdo4NhvxTxopuKnKM4/+klhQShIhO3NvAMrD5bkD9JuljYZg5aZffI4j4DK3G5jq/
Pter725FI4RkacX4gngLDOPHNamGdREDDCCRCltKf+aeSLva4s/uob/0N6vWLGa/VQlsiF524egp
Bra19GQbfjBdBeodsx29oefpS4yKzV16Pt8XUggZzSTLdzesDyY+K87kI2HBVmzwER5RPGLy36tx
GyhZo2PioTy0HgCd/Fj8q1fH48WkVMG6NI90o9WqilCAFJqfpIGOVgn9F3XfhTrORLNFSi2VXY2/
Rq2lttxIB/xTq/bLgzauYnQTYCq51K/8KHOdjk9i3rdwNX2CH9k/47maPgMPEGDAEUBU+4DzGTmk
mIb8EgZndVcSHB4A/Br+Do/Z52Ng31FKdqn2X5M1tGBpzq3UhAV7l/6vjsw7tYISId3f2tViHJc3
bt07q1KpNYzB39LCDeO/m9HafLCTHYbg75bx9Bq87FxRHSvGNHXzZAXBtzy0aUOXwl0luuD61piq
gSeQPwqmDJ82Si4hYFAnbuYTJKD0Ariqt70b4ETbw6BCsiMvWumPxHF8azuk9mGHHSMUKKAdyahb
VMAECSztUT9w4WXgPCIinTHxav2b2XhhO+1QeUHSTD/nIvIMrMQfslOubiP2CgZeHWrO3eirb+2n
QKSfMoGgAA1u/ZrqKhlq8NYCUpLS5mSP4kcSAI860vV3iMD+525QRkiZswQp0G4JlYjcz8yV+K81
GVw/zmiqUdc3rBL32e58EGRCmySt77xogNJu/DQuLUFFK57Fsbyu6+bP1OZ5NZvfKGV3KA/hJKLL
kTLdL6+wdo0MV2IFe1o5NkFgjMJwW9lvlrQ2mDYaYRB1FvTf1a0ZG8X1AlRUD0m7fg82vgMRuauV
TCpSVwF8fXaIrPTAbm0Z/NWlXTs+mLx2mD2GrNNw0Qh1hh/73QqgqKlOPeSGJD5OFubiHDIkVhC4
dSKhX0L1IlR0TwhWvpj8kYicyLRmSTYfvji/dKiD6zu4UdlJZ6OqPMTw2boyabY8kOZTr0ZHv6Dz
x9gIVXnD5PBZcbeLV4lHc+3vBILkvGFQzQPXicfxV63RSyrPc0hQjt0NsM7TQXFAzg3oOa75lFiL
BGe9+L4y+Y1g+Ks+HTI8wK9uJURdIyAZj+E0Bxor4Le6APWXB4FxQsbX0jUr9FAuE/KNLfNyvvwZ
+Rzu/eAjXpdzxwpMulRLVRsAMTVKim/8g6VBsCOFuAaPFy7EiK9KRG2fBsOPSv5cfZmM5CP9tqAB
kEfxiu2Kokj86iAc+v3y8dZzUw6BIK8CwAvaaF6UcvifVQEdO+6X8pXI8D26UFnpDp8k1o17gton
s03WyLbLyyPyMVo6IKYecnBxXvLcmqr+CVDEhlVxvDFWKpsjo49A8+7Q+hYs35K8JOg9UCcN1s8L
5tI7YU7X/sWC36n6Aj76egdHw7zWUm0WvJ5dGTbb3MCtj8jwBRYr8gq2r4Dh/5NJVwQic0LECO/8
zhkxV30n9vNUwanbaxe5o4h9RqzTi/Jl+fYc7DdFlDFToYQCitXjk4/IMcIgVtUohQSpggrN9bcB
I7O0pAEeHBuYGAtrWw1k+Ext+D6vs6bwcrsFfdAPC0jvfGlB4KyDw8tTOcWt2hAeJ980GPdGefkU
OU9Y7JXWwm49xCP1Fs2KB6eJwPHtpZrpUo+J3+PldL65EzPz3o2SwPRy+MypQtREJ0A9Ex5A/IhV
yEr+SuAdWBpQtlm9GFcdjRScHzGzj2BdmaNrOLI4j0/Q67FU0RrnjqDXelmH0gZlXAoLn/t0pbs1
fC1E48xz1bJl8O1RMA1m3krVpu1v6CXHQ3XEi34g9XiGysT+RAv6wcstgmxxhg3cvLgFYNzNyOm9
UbnKd4uEnJRnonEjFypcu4cAoDibxJlCKhujOqMO8Paq83a6XCebEcb6EYEJEDwZkzeqjsxmwfVh
4s1CnAtioiUxZIridUucHHKX92P0czYG2iVrGtVnF9d6av5N4VDTyYRzcT/VVwad9GA0e4afsg+c
nmFGiZ0qWVTpoCgZYmONMOQ/aIhV0Mzj+51Xpk7oz1xI74s8jTgWbaJ+UGgJwcbZcEI3h33VeVTB
X12BK4z/7vyujoLWXgUvYUzvbma1AAIGyjR/qgv0P8HChs7v38N/lXue/sH3xSABztTU20ss9N/r
Nd1+tmd5yvmg6dTjbYwFniO0PME8J+YsxN6GKe8/SBtpqhALcvNqOpbhF+En96aEpcjpuWW/iGM4
ASYtEqxkYf2HyXxZ2q5rNA/dUUjki6sTWpxm7XuxJCGDtbpCUiiLRG6RNaTrlZ+1CfgMOQ6ikS9X
mZIgfIsvGdM++zMp4wOyPMOXTsFdYAaGH8e8amUxTZsJGQWv4fXBnLw8i/p5ipN/pTuYTx8itPUa
zy4tPC1SG+xOo7Y5wTdD8kMEj+SyLvmpH+m9zpTapOtv8ee//bPfIb1jikFZdoSPuvGxWSyRqFL0
cXUV7gWqYZFIV2Fl2eOUjnKdi+kREvPl9d38ecSCzpyDaBLYWrJeU+MUdo6O/sqUSE+nDDeTJqZA
6hiLxcxjc3AbZNOE4s6qmEBxlO2q5T5FYt5/8JcWy9iRq4MtX9vHF/ijxC0TpRZVS6ryxnKwFIuF
cny+kfMwjtlDsdmgx7yPhy9hp2kr3/zMVXVISbILAC9wVccMq52VrFoEWiO6PZU8rkyToEykFfwq
kAHPk/ynFlVAp5uUUAFnjafUmfA1J5apMin630Zq+ZG/2gZUwCusrkGi6rlFbiid/hxplVZih6RZ
wdPuTQcVgMWBpQOaCx/aSb92dz2rZYwZYCcTxdaGQIMBSz+vaLvtm+mReyUUlWWNmF3z9owzAJvX
EJrMUPupdKglzTnZS5riwfT5JRMLHd+2XfM/MJTRBgM8GcslAEQWEGpAPqfs3iR+blbgp0ncMTYz
7N0YtJhC0y8g8sf4rcPCQSS1e/HAUvCznTqgQWch6pJ9+2EQa7p+aXcrF9yppiSDDrCS6vVMWB+B
TxK61Yd6hWr4XNt4ZPyFPflZgiO4tFjvSWmi/vvrxjiO3t/OO7+krdeqPEvpRniXYHjxtV/Vddif
M1mJIYuBJjp4M+O6VFx4EZhm2mAb3sgz8vWrXLC+sMXoVDwFE+8YgOYZHbU1RqrvvlOyBr4hJneU
haybVfYHOtHFoAL0BdSyJ1yDMZ1+/5/oCJjeatMg+Hg3D++fcXZTZqMCvktrv3/cF0BWFagIj2Y7
bcuDfQKiQ3A7zFnEcbADC2+1usfGioA9D5Y8CU2tpVGOWMY0nvBvN/fRLzYK4SmNcaxovTD/8Cg+
PQlEd+c6EQvJhKklqv2tP4ItsCMdtAOU0BrH7rtS9PMpvWfe8Vp56yJ96woyKMIcWfnGS7fyYHKn
hHj4lJ0BUef9Dz1K7VWx/MSWBnvv5Es59HREgkcKnlRFphMIvGvT1BklNobJ6m4iQ6aBoyUqzRIr
bDQ+SuCdkBjulnWd/forZzyC8YDlz6nzxaHVBthDntNZ7e6UhmNM/5cN+dMaHaPHxbOCXm45HJ+/
Afs2Vs+4qW4tZ8O+sDRdxIChXxy5IoBul+RBew5jOuEsnvm3J968f+4gwV1PTI6cTNNEgV6dTwvP
i3DzJ/QeyX8wkHp8cu3dT9LG/MqeDlvy72wuGLLna00NG12g/27jUOOFpaBgJY5Kxaun7hy3gQTY
gbnE3z/DUlvfyy6GXRa3EFYrRy5vc3IdIl3lAoeHglk9oWhEwNIMjrmzsRx6pA1SQq+ntU0DBB0m
K6Kt340JqtBVvZRTzTjK6Uo6B4uny1+aB0/l/Y5tcVEgsOfOWvG09KPNFQWktXyKXvMxJNJqBQwf
tbEqk1UluDSlddqIMsW8npCKbNM1Uj7XV3e+DISa+lGnVdaVdTmTLvHoOitnpiHAjvAsrNEkNC4V
LkJb8KDU8BcW+fhqGtvb6e2zQ52/AgClGHRuCLg6AgXDiWx+lkUpF2+U6Gh1tken7NIZE6CRS+Xx
r65RSiIR75arzEcBunnPC23L/HMnzZ14pxNPY6GkNFYGAxWY1mcEJA5XO+vEXCxfIxCrj7pmYvtk
Pj6rLE93ixx8tjsyr0CPvHDkz7Q5TBiQ3spdlAmx2j2O5Ch4fc6Q+y/ajFgf5h+0GTFyUASg7QF6
EX3PZEdJQwevdo4FENvdObOk0K0hqwxGyuVi6Mh9M9+1ch0rH459rTLtRwADRUnInMWvRWhHyRcV
UTw/OePAR+Fsc/8pXqnyHtQO7HmGybWlBMMXD6X4Lr3LViyMpY8kmLcaALECB0ItA+Mf0plvX6SS
4Vm3GxAz1eRtdryhuddcVL2WlKWoPjI+9Px/76EES/0zJTkwIhyb0I4/3J8D99kKFxINEXcw5mpn
m9dqLkLVwhHA4007SIoURP8SlABUXcd3cxPX3HJ2txr15asWSjRsA7naph24us3rCJLfXbYOQSTz
E/TY2qqk2CMPz43HbSN5IaIGsBxjwnJIDNXDliTeJtjI/YtyBj2rQKtS8/RQEKx6aA5hEL6m5VxJ
K05RaK/sGwd44Wefs2EkfH2/ishjAhVlp7Ql7WMEQ6F4N5bmEm1oR9Hqp5Szz4ZikqYocL908Ou5
mSl0nPtwmr6peJ4hKjQXplQIINgfAD2c1RNbi9X3PxfINEbgTdIMpEMyGCV5RSxgzeRHEd5fW+Us
ZyXotmI1HMFryIwYxZyM0rTCpmI1J4vxoV3m+mzXwsu9fZVmBbjvvTnGPrkfaYDbT9GwisCzilC9
S82cBPwyGxnDXzjbNrLMgtqeGq2QiUpk/tDPrE6eLgoM2VHYiqmqJUw+/4RELZ/AKhj8Ue6MlOZT
yHb5rDht+mVfOwSU2l6OvTB68ZKQZS61kqdEJ3EUhhISoweuXLizow7F/lHY3YSWqmDx+1gT95fT
c0oUqgfFCPY9TN+xCYGLlvK4JoQ3Qv6a4VcO+dJ1JhgjIso38faf3OBVtH3Pf/V+Zppb4BpYZgVu
fsd63xTRzPdLcr5vg/jlJl0mwxfKXS/D/dn1RXd1K5SlWVpgRY8yFoojxow33bbXMkzRi2kH9wbC
TbB41sbxjsPCgfveKYI+O//cs/XitPlJOnj3wJvy9RexA/ZHmcFJupjNSAXnGvsKQtu+BCRsQAM8
wuN+S/fo9WzzKdfFoxF5KVehcxkvWlriQOH8PCIsI8L7T4Dhx3OHk41fD6VSHQ8pKu05+stRpsc5
zRXNuvRdb3VxGg8YLDH5Z21/DnMsV47XydCJx08JgTK4v6O2NPHenSPIiodeO49IFenwJ/Kpdlv2
fwCcF3uUa2Mt/OftGrUDlqP/FTnsNSfz1ESHaakLHgTQAsYOscptRonnZXk1IXU5a3bzEhZQao8R
NVdiC9GBx7D4VS9iLTIeEvf+IZ+vypAVQSs+vabb2RbitrlkrZcuy2KAj8idDheD5YGp/SxXqMB3
TFzSHb4fx7/gkSHM9QBUN5HgBxV/IRxGVzhMbgH6S4sV3TgO28l1V6uFQPDHjortxpNYZoq2Apff
FoUIusqE9pEiBQYZb/KNudUhxuBZI70GMiJwV4Q8dVAzM/UDSABQzYdfzsRBzoowWhQootH52dTX
wEFQe2YQAVrQ48aq9Hw8u+Sa+m/q0xY7toMHBoSE2CryTP/PWdvWD8KTVw3R5xX6loQtiDZaTn5S
A8m3SeHfp4Dx4tRXS4HwybDHXT4UkyRgR4b0lCCtLGY2lJLrsqISoouhVKb+MpmdLs4f3CoCtxrM
+tTUDiGKo3cD6c5gruUenI7WWOpt3JAycFviStK4Tew5KKwk/Wc4SmaKeGO2Y9/2iWOhcqnsdBJ1
9yuS4Ja5id9T6+oLRWoaWLzxFQ6KRP6JcFN4j1Z6ncX3JNdChR537E8Ttgv8r6QfBYzRyWmY9SEU
C9Oztt11B5A/fEtbmqP93I1giOkWEnmHIQM2MO6OixUjdNwjxNLNZSImIY79lbwj575pi+ZcYSrW
NKN5/vQTC70Ab40nVRoBCEvcIicPjWyF5Ch642esQEG74FPvBv2AFxqiRPccC/sj9xEQdw5YoWrZ
oUB7tciXfOnJy5b/QYVudEtGXF5/Gni/7ivVpRuXBY0UnYtR+GFIUowTXkxOhnxt+R0D9trQcUmf
MCTRsE0qYg7bd6VJamgAtPCMVQHPLQmlmr48d8BCxbB2VZ22QwhpQkkfexXi/PuREquZR5vYDV7z
r2s872oTO/hcdADoJ97amSOfTyt3YIT3chD6cJzawBga8qxyCcVleHOe1t/eXOhP/G/1T/vB/gEW
8Pn6adV0jldbdUz47TAREYAu4kIbeg3QaL25ZPzJiefOkI2EFr+RFBmDLf1o2NjVMsqrVYa8lacK
GetjLgpfq6eHbQXHI5RdT6UobhhG7OgVPOqwYT6vSwyXVRQpbfN0nsbJ+i71hF4voyEz3Dn19hmN
mHPXbqoObhC1x4UKw6IoKtJ0vGCU867oWumFaL5PhTuwkXanYsBqNxkpiJ/hDeyIm3oRx2+luDN8
BYm24c8aGGFQmfT+6s4zRF0ys4S6mUiofX3B9u3/Dc48oE6pUzJsll/Zoyq/Dx0C3K6y7awV1lU7
0gI7pi5lFlFeEkbsIyHJRImSaUqUpze7C0YWjcb0ZdfyWsGHP41isoeFrGHusmP5gPSXQMoSiEdW
b5t4AygUNu0coI6ew0PtCrxlxOq+elJZcemsMbW9SlbCUftf7gPJ05K+Vit5Ot4DhXg+E0bOwT86
rup1Ep15XK8c6tGFBzWc3Moc26neaIp9LquYC5Djiq7h2L75Ev0SbimZf7wgAimtVoO0Wkiw5XgX
Qu1DfZ8jEUvnhpxazRRISRlxlbchVZnxUYYtBV7nH3azgc1IgOfINH7plcuPFGXK0SfFX0Ul+hkc
v6HFnPGuOG16J1QmV1TmWFQ8FNY715KGQD6ulyVtrmGGPfTUTGKAmMKkpWKFnTw0/zIpGMBv3XwG
GhbmZjjleSMaJ11kJv+dUkQaPYTRTLoFz7V0y+57utfL66IkbZZCpO3tJDeRtBFPqyBeb4D+quxp
GM21N1tq9A4qDJiP+QY5Gtjlsle41ugkBvJh5nEAHWxeT3KhQbG1Kie8YncBrIcfQu71vkuuk068
Gg3WvIP2H9GEw80zsn+0a7qM27ofiG9t9mFJo26ZmJgQLe4Zi/ducMSgqO4mB3KmyHo2xdh9NrJ0
kRFo/Ngf5izFzKDSG9kyiXzIKBpsCOkw8e+t/q+qVvXvZ1M67eoeAMCaOPmUblcKDhItxH4a/P/w
l3ctnlgt26Oac0t1ywR9QoxfY6uZ7L6phURWEokTd+EzmBb/0k6jRh+AakQd2gv2WArG/VKC2Iuv
R3cbcdxHxjo+r+/cnlcQb/bXlKJ/5r/BJd28upTi3UekzPBHU5YdUe/57vEhjhxAszgMBixMdqs7
nwRrGSas36WaCvm4UKSPBfdPc7U8T4R66aMhupHI9OXSS81zBxasBgy4Vt0i2ITAMrRIZZRa0BDH
eTh5r+4sHLCgm9LZrZWdsjiPd0yOexs6s775MbTGpc5HAzMtny06P34HuhXndx4QVto1YhmDKRsu
aVr3afCShGxYpifslrBPLlD6Rk9pDZpKG1ppn9wKM1fSO9INZ43SVEOUg9e6ZqZcNjrWMBxJBe1x
KC1bbf45f5LHBVwpz8aNxZ4WP9H4188qlXEJZLiyBNBRFCkCxj6IuBcfcgmj2HisYJUn/ULRCqpG
k9PkMRM5EtayAr4dlvHkb5yeFBByCulz34Rp9mq2qswDP3viqk+jXgrvYGnk7JmYdy37SygxVmpi
44Obt5yEnP1dAl7phBYvwv//ElhFV50UiesUQXo3kBNVOJWmdYtmU/xslgelgZM6vKkYnmHlKX4T
W6bsLKzcvghbPKPGSJQ/WbcUEydorus6JoOR+YWvEiPTL1XKxJFT3OP0QZWUNH0/5LiX1050WUju
LRYd7PgWJXoZBTEAAvvCgtGUu+gO/A/0YWCGPeojSrgbhUev/kSjPkuxEQTaggihvEkw1JvX16NK
5+I97QK64YPvF4clCF3iXbdEHFKSV92ljSnduVZ9oxmnUWPCqmtPSkX5Y0SEscMqtyyRy/NVrX+0
VuFFDGO7erps8JJ+k8FiUfiRrLmziJgs2T3rfikIeJpmU2Vppity/Yvt4Exrny/5dzs8x2iv+BRo
bMaiML186xYl6N2bSEtXuhhPI+L4eXO/Nji9CtrVZcVCut4kTVmW1OT7ZEBxbIwMXGNHJ/Yvd8vK
ozwdSaMUHDXLK+mFf/2D5sQSHtBLkae5Ug5RZTMJ8OZ3QOzEd4g6bwyHGvAVV0DoVjfhAiFwr3GM
bd1aA9bnjSDKPX5e/JC6wZ1J586P8AQURELME6JHTR/e2a66eQ/Jk19rN8Bk6mcGG9d/dRfGA5Iv
AvwYp00X9F4ZkP3Y5R0nv0ca8Vz8lznsDFJU4yWfaDXAtXVKgMec0RcPSDees+ek+bFuvAT4whrv
q19uxiDsujjDedoLpxYGvmYeTAOPd6fkL0+8tGtsVcWNAnSWl78AeNtv801kO9VfrNtyj5/qC7WL
e9k7QTuTvRhSUqFUOcBznyQk9x/DrXW8gGrheBs09rvYbSCdE+GSJjZrUcoJvUjtb0YuawDjxQ2t
lpVn+2CqDSwpqFdfKPt+vkxvIzWvwJoJuGy2Qn+5H1dxIPMqtoVC3JXKyIVk+ZRGdJJ4gP0rZ3d3
esB2gDUUndBgDyBP8wcSy3208RWunHHs35f9InW8BCpg0LybQqikw/1QPp/Um38+UM0hKFc6xP5z
71L2jmIFcXUy9+5pldvkeDoJslTBKyiIb+j2gm/hCIyHaqeWS3Vecmreon358rPKDI17cylDZ9p3
l8cfRGLI37H5Yo3HV0bJHJlbslXtczU4HliwOGuxqySRzOiThihZ9fkp3pdRCp/ipB8gnrUMn8Mt
m09Q/ereA/Uy1sIqJGD9yLJtvVOjRz1ELJPX+aEwKC+MNr9EdtKxqwBqeSrhuSqPR5ampgV1wH6z
8J22pM1mD7O86X2f+9WjScjHuCqnlfPSqgPXQfky6IqrOWwr+YYKLu3qapSI2nI4fJwQDXKQzQkT
mxFt/RNNtWTrdrwJwfoNK9uEq+ClxsD9oX38qbYIJnPQnQuC9kscs7TjEwcvb3jJ0SMMfx1Sgkan
85Q8v5vCe3LFM++SBoTn+Sst+AhXClZ5kx7t9ZgNjqypPs0GmtlT3+E9Ujzu3+lg6wbBV911UQuQ
7zehOfkHIFjYowizb4nGNtU4z3m4+cfuyEEY3bp+hQqNJpnS32pL9WPgZpgjvPUw8LPsVhao6N9U
zPlpxI1MI0vAWo8NvhjA+y+Du9L7mMmcreJNO5JvVwGNchb0xlh7ZVQttn25o16v4gbU7bQTBa5I
OGNxgkW9pmt1KCoAY52NlZB7yLw9oyWvoqfM0/cyAr21Od9AsRMRVOK9sbaQQ85wTV94EJ/QBRTo
zEs6PAGNBseA52FjMaGDssgYGKOzB9PuxZ5JNgfxYSiLeT6h/CG+6exKfA4dYW1W/f136uVI1JIw
7kpZsZ9ySyu5voJQYdOT0/25oEr1MdK0AnCbnvqtvGpN8OXsmLpPOJSGIo7YAa6cg23X1iSQ5eup
Tja/XANjOhnxag0+ujHGM/Rl279coc/K51w4Br/jKPTkFr71VcX6jLMDDOSbYp/OE9VX2x5xeOw2
eb05WBJmz+NoufSgUi00E4QOns9aB/GEglXiYLifp/czcNgpBYxkQTjv3/o1kl3r/09bho5kwbuz
4ghSyEDzx+QAd1GlyM2uGlP4FfzAt9JhLKnlIwg2PC+dV+CvxGyVArsZKd9yenJHADUPaX4+Vb9R
rZyf8D5cpmaLRrYFcyjCI4ZHd9pynSYeEkwrbtonSOAuA3LjEz5Jz/8jBoqaE5RHWnddCoYSTA21
1ZIJkSlEG1kPlGRXYt+l2wlKe0ziS6esRDY/EIotTPxpJQdjWK3w5V/sUH1WbG/sneJF7BaxKfqt
RGu1Lij17GBU6oTzNw2e+ypMKZztoI+slGZaRq0i4pa3l447bfUxoW6R5EZb/L297429/37JsZar
HmsVY8LazLx7yzv/vBQ/ZsIVwZVluigP+LOl5zAlWmgwhpxl3VcKiOmHohfAWMWygncpuie/R3Cr
e1PVfKz6XXOMohKY0Ra7szkGFa5WYTX037Uervwyn9uJM9hSMb+G702X4IcIoNU0C51zW/aVW0Jw
xwhfhegLTz0H3w5pRi4/Oo6e7N7P8LokyYBYc4mumfZHvgJ+89sX2SF/M2Z4/BQMWxtOStAszOzF
A517F5tvKj7of/QAUvudjJF7zYj2HWbWX3K3zX8UUbIKrtE8DyP3SgykxxzjeFWn9OCXB5+e64nM
1+CDlan3ARPQJmZ1eYVmZZ/OtAfjZY3rHQYOZcg6KahgzpsIfrBISQ+3AkvTT+1P51695xZVJl67
kpbAtYaHJy9kJHBo16cXHbLNdwyoQkjZ4zj6viTBUZzjerA+99CW4YXczYyDkNBPaCF7rQCBTIKk
4qeSCylW3lp2B88+4esTsZZNweIOMuIYvnCi4I/hFF0/5WY0F/stUy89panWbADco08GUbOhG71C
X4y9/ulvm7R9zy66Lf9vUOefXm8uYpG/tECqBkWJUrYuin0/7mw+ijoquXj4xEN2ir7gZcyw/4ou
bx3bDekvodL72JEfvGKQLB839rJRpffusQ9RUlOns9yWOgE0PfSy8suhLBTxkECERmxoZyV1uPfV
+8IVjof4NwnURJUb1pzFxCiPmr10pOsXEaZ7IqI7oR9REMV2RQ8sppc+VInYidFsLJVXJqJ3Lm1U
FGYLaXaxnRR5GDSERWVfJxiEmUeKfK6CFJ3/tJhd56oyHksutrcIlao2eIuHWyWUkI+jGy2dm0m8
0FrcX1osSjPzuTNVXq0pjo6BPRimDS9UO5qEXg/T2UQL7LXrg754OhO9Xv68yKHE7uoRheOhwGBy
b87yWKdLWHsbSnYrC9i1950dkNHzBILjU8q2nRk7PwJUtSrNSl/hjsVR7jrD6fr2kq6fR2jJWgHT
8eHRKw0zff8K1pkCZcnrzU8fOprxGx5xsHyUxSJAwdn0f6YZImpfiE8KpnNfxa4k+mpBTv1hzi64
hH5jiD1IaoJhtH/+z0fl6p1vzMWKzQH1mF+Et811gMeihGFNscYo0S6JJ4/t8Qng5nNzpxW22IkJ
gW8gpq8lK1YeZQ36fAh7Hy2qKBhuLFM9qSEAYpmkKRlDheJQCDGkm8245/yIEwqzQxq1xJOXVceV
wN46QKJPGg6p11FxpMwgAH7VydSJv0n0QCHoxoCzpCb4DOsTNTvlUjyzeXwVynwXCrVQxiPgYvCG
XkCFVqJkSBQL3wTgAP/2A335zrZWDu6kPrHWLHPugSg=
`protect end_protected
