`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25696)
`protect data_block
49V/aakodeEqdERqUxbC6CT3aRueHDMypnG/ltsMd8nVCMnvVzt/WLhpIRm4X6rpYBCkEelRUv9Y
Y/KCSrCmBoy8YI7hc9OXXVZEMcPaX4uXtTQ7oLAsYENsNkwLkK2QRK6K8Apl+EoXhujlL8swi4Nf
aROzikHFBAMfPtPyHtJOhvXu/H1Ez0cnTpQ36BSfnVPjWmEOlqz2WMl9NJ02NgMeE5pN3aqKKSOP
BDkIZEIYnI4y3j88BZ6HOVlt3ySWqUXj9Pm3aNKqbEi0CTm0kdkQCy1bMlsKXaeMg4NrrEZpSNgC
L5uvK2qwjmSHtCWv+O/J8nhkDqo9hJIXm7tnqGL62ibEKvJCPxLiNCvqe7Eipzpb+1B7EPm10RJB
M0IhuVvSe6o7p1l32nt4Y7cUkCU2l7W54yBx4x7mngMfQ9qpqPG67MVqk45mIoWn38p7JrF+hRfs
PRf6RUcZEWaEvOzpqnESJGvBlq5hJbQquvho+2WQQw1eJM2GEcRttIaIGHQYI2Y1unfmqgYwvW6j
tX/hMKAozNvvN0jqnYOt7tS+f4A0dsA1Z1QQfHqOf56fw+icZtbzEGZXHIddArzHc/dEJmmEXcBh
0XHu97w3moZzXc1psiA72Y7ZSxwmB38L9AbxmBUW3PRQEBSqZ3tGSgV3lOWwBvfRQs9c+zwYRfJl
ip1YydH+RC8JJU/fXNJ6oOT93sLxxxoTZrIjfIqpXZuUCCjQnag+GtxhSvfKtwJ2jfLR8Ip+oEDv
IZG+Gw+omoyQ1y5Yi4QNb+uTHW1aOZyeKekQxLkqS5COF/QrKSTUTTiDANF3qByR7c5gp7W4PJBP
wh5VmzpD1mKIPiDFzXIWBFzLimfWA08QulUs9Z9+M2ZdwiiDx0zdma0Tzr/pvGWgmWwFFibG0oEJ
lxz6vVFecHxDyNfK8itzKHLFBHFqxlinOUBpc7LuHbkCetZFIdJT4VfYQhZ3t1WdYM7Pa8WDL197
bOlQFUp1z0hXIUfx/oNBS9PESyhgQ8gZx/CPmlU+k0axNxFWsg0iQhcsR7mh27+6K16I8gsiTfYx
Zf60YpzIwhje7vFyWRha9/vVttjNW1W4lS0EqKk2KK6mMmAX9ZlH72IleWkxMML0ijEZ9MbGH9j2
UZ8ZlCcBF9ySLcsoNldynUlivgAbsWZ6UAxgYIjRGIFtxLT8hWpdczwd26DvF8RszurIYaCBI5Wz
5AojtPrGuvXmUxwwV0ChMDLTsYc3ktFtoL1XsrFfRIHySaLnuSUI5tg3DriL1oOzX+LIwSTswhU8
i4wpsl5OSORL/HR7KBFepRMsr/xgvSWPMb473ww0VLFG9l+53EfvSx5UHUxHTIu9Yjl2Fwkw0Q5l
sIkRW+k1O9xgiDBzRpkEYJm8qIjqzT8tXaFtxER/8ETt8YfdJsdiDKk/krs17dFdR3UUQ8+q2Eu5
zkmhuv9JKjDV/ejXZUQZY+Y3bdhwh4qHZOWeuuk1kYVjSRrJzmJ+sfk8q/qUTDzBvl6BM5gNg8dk
/z7pgkKJa7uY9e8JSwxilLZcyWOsFs7jMx9CwP/DbvsCvvezIfbB5Fx37Nda8UFjfG5cmv+akUDC
pGHVSnHOHDNdm8G26Y8QbXif0wlf+FxrChGyw2YF43XAg/X+E2biaPfAaDpD4NreC+C8xUoHrbRQ
1obx6a84Ov+BRz4LnTRxWUTAhbnlR9P8ude1X9N49l8ULH9IJ/DN0H2BpbeYGcCjZw1zugZMKkQi
cXkX9ssAXyAbJr9ZK1Q4YrYePDKXghNY4g/5cU/ZTxU26tl6OR5rA6pRZD6xEcYHCBaY89PAKf+v
Gu1539BjD1YhZ3kmzU9AlZF/eh7EFqx9fqAbc7c3/8oi34qclj9Q0JxeNVLbMaCc/fkVmCHrtzUQ
iVI0sYg4LdkyLHNmTMTqPQpjAmAl9+w9555L+6wMDOKJMI3kC8/DKYiIqbZ+nUToR9FUx/SdRYRQ
Fkyu66xNTS9jHOROfRvTRf8Ri4Eu1ntVMI0BQGDoK4p3knEGaCTVoO14Znt4reRYjPoyRgmpRpA+
zBjwstxQeYZvByzIMniO50dvblGQMYYWKZNN9EMat6zEBDr0jN8fbipflHQJtMWLIj2fSn4MKRqB
e791Ux3f7fCl24KdKe3Ah3QKPi2dxNQfBUbjx/TzsYnX2+HAsdtvNYBEBv8qfOsWiHmzPWGqIaIX
m1ZV1p2m5D1Kp5H/HAFMJBRcb13x8rmaUgSlsSCScBl+7PAAMp9siGCWbao83EBHvMIXlj6OAzSf
D2NijneecFeRGHVszuAIyUSn2A1nJt4FnZBbVKkW0TfYuQvhnsdx7tcT7qeutGDTsCKYyp0JypFc
28ASTs4z+UeXHPOVd6G1591/MhKjHl9U+CepLRqBtSrfBH1sOe576TniBiL5vpu2N6jr8As/THf4
/HdDNR73W/zwvVx9jRYjdfcoBv9AEdAeM59yjpZz6Y1VTLmppUkB+oOGRlX6ioP/kudqSf3y6JIk
sk5T78nZvBVlLXtp8/H9xv1xSvVGN856OtqYkXwdoUI+cnQ6Ng0gM1oiWSf8il2dvHNN4XQU1g5z
S/xmZraWJi0GTr+eFZ0QlBfOlEbLSBMePbCsDQ7MAwVGde+iMDvUR6pSDXMTD/t1yAEhLZeOFYBs
LOn61IEJRN3+iQbqXpsvMgPuhYdolyPpv9yjOptPYSczNm4+KGYtYfV6VmnL3TEb+zfOVWM89He5
Y9tD5ClXdCUJogw2f8odM0uT3kmRsVPI54haqpOTTWiUQyT4mVOuiVMDp36yRvS3aByJaYmR9NsL
jgOWkADGveyEUXeziQVdOyVYEoU8OHKIAQvr2u7HIrdM0P4cUJYJPYWbxD2xnAHIUy/g7QLWw1Jn
Drp5330R0tgYvLMvZn5GhyuhUVmpVenVS7k8OrPw+fPRszaPDKkoPtfT912QULfh6I7CIHF3DdCB
82TwqI/M250m+T4vYNLzjYpvYvWgvFJoq/DOVr1B5wetTVZAuN89IZ4jNVcY0bAQsOVBNSVIgQts
+tqlMVdibF5vISeDOTpujU4c19QkSnyA1K0JO19mk4R1lmZN4n38rdq6WzFh/Ovm8GuEia4Eu7o/
auk9Jb4iWhXvaM9HggbUO4JCRxWB834rKdiD8gX4HrJfRMW+FS2K9+hiN6nM/8q9nXbaBdocWJTh
Te4ewx/HkdNVRM/3iTobYD/NPRRBvAFYKLSe2/P7vhX2hbbepDB+Hl/TrH754TMRelumRxoCkCmj
K4qZBPWZf4ZhnmjQg+NGWHTewK2cO3Rn18iB6XxqrY/JCXuOVqsdZtM3626Tk8o5jC1PlTenfFHM
ww7zteE+VL8z5bxf5I+Ec+Y13a80F0CeSlC/oB2MU8lTDULSk6PbmZBQx9bSKOWLYrqhPGUJjo+q
nddLa0Z63mq+coXs+8kC9J1+dzGj7stjH/CBmjKcw5siQqy/sA8ezfWIVxwLl6Tokfor3W3dB74Y
ZeiA4aOt7wSf2uerB8jiWzwCkwAkXU1YcB7g7OulFwQLPcbmMfrmkV3dz60lPTl+TXA08L6CYPba
eJIogiW2jddkMj8JMaHOQ4J7bjksCo1l1XeKeMLs1IN6KVUQksEUDoLgSaugC4+xB0+Iwld0r/l/
1sUbsANTz37qEWI7HxrnezYuuht4Y45ji+PiY2VKPGSBGrs9gIlIF33JQxKhcrhgFK7tBSG85CxH
Wf32N5he+ojLKOp8VD687rHkYFbTdCopKIYDwj7zWiEUOtWKpZ3j2hMOhkkXA9I8417MG4JdBage
cNq0Ui9GcxpCEnu4u+ZUisLVkapUl+MUfRy3m00R6ujPJc1l67Z+rR4LrPoeJnF6H7D1LMNdZ4Fr
eBPmptvSwjqh5joFlAkLZUUqHmPX6zQW3vCe3wypJWJetIEf6sUzCLyiJDn6CdFHFCGdMh5G7dvG
wOZtx6ZMb0Gqw0qjoeYLLLN3s/HR/aqzjHxZiM75QT3miMG5cRVBRPztFTtwND2nPPTyBkyrKAuB
vr4M6FVw911/lOEjsEEt5iBMEB5ij0onW84/7bC+pnrFK7bDSihRki7CTxyzezuUwgCcb0XBL0L3
GgGGP6zgKUcJCD3z6Ajs9taDtT42zSWMPKH/JBWwMd+MSj/ekgDS0ZOa/6oOku/MeoRQ6AX+vuP6
R9kyGEeOU38nsjUnEDTFWHtOdSvs8V+smm02E9qGd/lrHAyiGzchI0X9mGu0kU5VJtVbSk2VBe7l
nqf/4lv5i+48TIWFxBzr+cT+rYoWJ3yJMJLxkvV3HYBmvasisnTSkbtwHwjeHRv4PMfB1fGJ1l/A
c/BRuTxWHYi73yF+/HgKJhm0Rjvb1uEzuLL9t37zTcjEbzBdrzLWIhmVEWuAaFUWg4zEFevl63Bo
4nCeZl5mwP4aMfkMRJIjZLsSEBINvXyjFrQGY78x38dcUb97hh/O2LZt898mNi8iqO0tNn6N79hx
PmzKxU9EpSd6ubCVK0foWoyE7cumiSfB8yGMfjgLOA/zLuvHa0Tqn1JfdmgPHuorP/guJ3IlISf1
Nn3WDrfFHdaLo8nKmJdeydqSbQSYvqZMYJUaB+zVPUn1vfgbnewHPk5ogJTpLS0iBm/mnSzoTBJY
4CdcS+3ST6d6wJ+V4lskCfkFmLHZN6eLkMwwJmpaOfu4uNYeSh72x2f1ChBt2ov1k07jGlxw8/oL
qBBdGvOdHp+a9Z4iQioUGyS6w2rCp2x2GcUAr8s+lPU8KOFmrSNup4I/F/dFbfhQNO0J6Dk0xhj+
KMuayBiV1gBYYUX3uFmE5NxVk8vGPlPEdSqybaqrr9drsUTIbaIV8f7fQD7NPbmim0PNeUwjzUOv
7bhghueXB77iVgIP866d2GYx7aCn2rZWor1hDaLqhoS7mleMH3FfRo7UpV1MxJLrnHiw/VTXF40J
doimhNYU4b6etZTRCd1EP9/qkk6bpbppuaqw9PW25oDA/n3BCEf8uZ4WJpZCRo7iLERa4BM7YhDC
jrg0Usnr7Cuos3z98E8lnS4fiNDEUmAX9aOs/JeD5m2yTROv79ZjjYUo0qLqCwB1qVA4gCBd4BpV
ihFygbXMHuyAkvXbyRlPAvJl43luvBR8xl0YB10AdSAxzvde+vemE/gzGRsYnrhXE5d9CR+AR8VO
UPBNoQbPFxkBMO8PCEMUopLapWMsg249yJTuA/DQzTEtg95XhdebpRaHTPjC7wIBptb6H+0/M3zK
nvgzdTrMUKlIdvTgIDeVRtJ6gfBS8oDW87t9dsSKlFzSINfH+SfEIVu3HtyXhyQEGhEKQMuH/7f7
c8Qlz61G0C2NwpyjZ2MdclEFVFQnZBDYsFcABWxSVyNlUJvSymAgcDE1zTp0ZPKDM9Uuhi9zOwvp
dTJpQ5r4mbDOhSvWkzLlyOvWVHHzY4aDE5CW91Qi73rQ0I3LIZWq8GRrviJBHC7FDU0uw0kacxpc
Dm+Qf/bzTfu0qLB08yGfzegUylcHA20l/ShvwGgWRKG96LHEAdfL2D8UjE53aZpf4rmO6ZVLQtdD
J//hIJEls6BTqSLgr1GQmDVNFXIc7PN1rgBbwfriLy5/s0iZTcydtJJerrmBVqepqtcdShtT5PL4
5dlKv2JRtfEt/r/Gbri7XgeR3dtmyMH3BKj2VlYLWXdKocXBWk2ij1Ey9pcMPA14sNAWgC8E4ubI
g7mXGg+OTOEy+Tp8yDKQbOsRUvpnQRPC6IeUqJlJ+SsgWFNhkQL1/2kkcOCE4cx8GRlBg56pclYy
IGxN9gqp/5cDnlMEg27TPZmPBbOEdiaydm4xgZ9nvMSzYLqILsAnAmEVvmCE2TxhnRluvfNbi8Mq
OvdltGQrScQ5Ml37pFP3+XmQSY1WppJ4t6JhBc2/8dwcNGjeYj0LInUOj8zJ/zgzX/7vB9gwRoaa
6znQN5/JRnEBTKeakou7oZgB/JrTj6r04RqJjp596wM8Gx8md7uRsxKnLD0eedw2PiLcZAp2lnVU
oUVBT+wwr8X8dWdufXFAl0942nAKhMuy3q9tA4tNtnWuhmrkmvRjwFYBqsVnJyxFVa1jkI9bPZcy
svlTJvo7Utkpcj4SGCmeAzsWQk5RIbqEAfcVKs/2MEiJ1K08d151DMq82CBWFvY+XEq7jJ1tFlBc
gR74fSW78KsnhyjMyKFy78/Lnogh512F9Xv+DOWdZzxrkB9zjczfUKRtL+BdL3YjP0vbhpjlVl/a
aqjhYuvN43N5ou/SicHRuQAJK1+6ymtXRzTlNV1ycpiPPWaigq1Xm9fklhd2NdhF3GpsUNyXLALw
C+k88nCwGvG9abEezUncc6GpvPuzVXuqsDv/kWMS6g9h+4wZ5WLmPiQoJo5qUCQ7U9W7dpd1QkRl
kGKTn5lUirRplVNgxo5GLZA1f3Vi92gUJNee+AB3vu2wvr/friE2lHI8XeNg2oft2RPNzFC2Fjs/
zVOK3y7g/6kYim4MLPg+4a9fZ6eqt1CATo/8gwwxn8GokTn6YXOTublrLGnFdTMNSuAUfIT2yCH7
NPI5/aYGh5PChNkx1lDTIokfISesEaW1exjwg0jaZYCdEr3SFJXWeI6ZEFCHJIm1vmRWBQp9G7O6
7DAzAo1lfBb8+jNAbcZPk5dFTMthYWfofb2z+DI6tSbDjUaoxZ/d5CpufJFuUBSx7dB0zqcWg5HD
Z2u3RoyjLAwPFfK7OzoYdEvzfFXZGHRFm387ap5bga2YunubIDEgcnHUo7iVn+9hMdd5fWGnn/dg
RI3ei6qsc8fm10ZdU2zIulnOiFLZT9MS4nnG7yE4AysZE+dyJzJyku3J63kABzcGPCj7tnhc2sSt
YRbMbYG6QGsuD8pjGnUguqbYHLCVeUP15TL5kw472LFGjrdi8y7fL0kcSc6Uza1YMOLCbpW/7N6u
s453j4V77QE/+UsFkY9hh0iBxsF9ZAPN2QV2e6jyr4omHyC5MsXiR03FD38tgJjqPvM7pqmqMrEJ
2frExWN9WB8pheP0uBzFxM6Y4mUPm+RTsRsoDvfaJWGty295qEmfg7SMO21cDHcF+8OvE/fBF1S5
TCAnVXY63FBIunDz4Khh5BxFwKt5uBFVmDvmRe9a4xCJAci8aY0ceV7BCoC06Kl6gY0hYhs62BLL
Kok+72IXzaMP1Po/qMX529riW7Qk9OMrqI+iZaFVuzcoW9fEiaGyEvhlu55C2KN+wwPs5xq4AY3E
sjCx27kARP2WjgRilBrYgjdxT4iXvicDdvRw9osVZiTBKg8Z8sicVvV6k9R3FRNktIDu62reMHdh
ESimu5xrD+DnMucYzveebz1rwGsaYCGXvF3pdJbpK8bltG+FDtUcEGgl5D5AolWPQcDV7QLL+E/f
BJfJFdSvPxbgKhChFfxZ7Gc7hdP2YCrfUgPxhonA7+DW/PzbYce7ah753E7yYx3gzn+khRZh2nEl
47MlDNOcuMjNn+nYdY9teyy1/c2Zjz22wkYOjWyfg4LmNpI6YIM7gUKhRpsDhJfqHsvmlkHdPasX
X8UlvuoOajycdLMpyHDY/phrbv4YZhNGkUSHq5NPyPv77Ek453PT8o3t3jkP/zQPPoyHJFQRAV7E
xLSpEhfhqXaNQWd9sQQYLQpj4NsQr1FugEfvBo5x9kfIfGCRfush/CX5mO15vpysho10SWyeBty4
G1HKpSkKCvs/B9LjjjCDhJ4Sy64WCm+BXqvTa6bBwbbh2QVayV6Pfw8Dbz9IO+NpNGxE7y6xSu71
gcPBul1JdYhK5LTa6CILWdW4N4FycU/WCWFJmXvMtpGpTpa9Fa05xb22J0QRhyhMGzB3HQaD9t9d
RHT6hQCum9A3IlVwkg3QeD2K6Pmzbwo9fck895ID5gwNZBRz9xbIrIeZmgdGNl/9CgAdfbAobCTT
jTmNvWMf9szwatjiekSIJfIGhZy5iyG8mm9E8Fc9rnXQaH1FJ2jZjkHquBbD5/y1bnSYwPrNRIRZ
yuSPVL47dhGEaHbLRB2cR6ztqxGuFspb+ol6LwRp9zbP5kGaK2dcp9DSuVyEHEMCQZ9hVv/LIYSs
nlSaOS8oNkJJ6MBsCSyhe1bw3FWWyWe7YIzqXNvaq3g/ahvx27HlEcdGaVJbQXMUnd0Ahe54iUsr
iGRsgImxOUme99YqaR0BLf1nsgjV7aKV6O1xIHMwe4ot7bthfrNOw7wyvT9FATHPWqw331tb4VPt
YDmRax6at/aaOc9CMM0QefVhWVEbZzVrVTwse/Rqt/EqN3crWLGnD+sjA5GSDZN3mKDGhVcVxZDm
vQF7Yppl6Z1/fqJHXWyIEE3PGPtfFZcRMF0hy/JG/Rqi4pOFJzaGdks2W4v5u7ZIhV6a0yI27V8Q
yc063Zh5N8Pd1CmLEwze/YNd1RFHNgKsDk6OAH7YDu5SIBcGKDGa0rj5OAgZ2toiN5SuTH196Gnc
JSpMWyII6VyRJUluy80z8pqoUZ75Cbq69N4YL3H7M3U26FNr4/uC+l1/Sz7j+s5JhVC9AUxmNljb
TFot4qSco3fG6F4ReQCNXXRfCrixc3MWhm/OyEcFQqfMUfWDxpwKQUR261vnJ8lt4wfN4obf4F7x
RLD3hHAzgvd/hm3vx/Rk5q9D0k2HrYLXV0CYkvHbXka1SKptxfLS2Hl0EBG6Qr+tbVgMmDPRxA+7
EZIo4jQIi3AMJeg02spmgvV+Ja8Y0Rsz9JArBHADiniQBQGKzbLN7CvuzSYpRsY0Nq+9bO3NCWvV
mqhIpWZffwIX3+6fUC0lJyeQ7p7PuUkVANClAS9pFDfdSKY0Y6VSc8aEwRXeg7Jie7619UidWI56
Cu3w1SnFklwUhxE1lKXJLGgb/EA/QfQE2YCrfnVT7nasSc09TngukMMYVRgaKZZcv7fjeK5ioWyS
vKccX3ofZmghDwtm9I1zeR+QG1GBChw69841g52OAQs38VPqzI/LtKkYT/5sUbTOLh46qbKEzd1G
tQXQ9+iUGeiNVqWbZm1aDxUMA2gLz900f+u33EjH8KARmwz4kbEFW3h1nXbp9fIQKfeAVfiM7E4i
EVoLejGt6lUr54b1awAZIY1Bi3t0Y1Jn+N9IUBT+e/0uzg46N4VlI3ARPnfyXLHN70juhS0KQ1X5
gX9jOcMUVZR4tPWvugW6QHUrmh9MhUcT4xmeFlOhM5eef6wY28gVnLlXB7mAJyKDJCRuOXfOEGMe
zlGMuZO+e6cKAUDO9XJvlw4RkxifIDcIMSFHZOnS1bUkozX6LrXDG+9lkUwvY+SCdXUhklmkmNOv
rH4lzUZty03tTwhVftOswGE4wrB6DVU+l9bKM0IrGofAe3xhcJ2vu2r/S7LhkPJM+r5MejIetH0b
Yv6TqorJ5+5Jv0y/6qFoefJ/ZEmsFBh4FXpOrkecSnn8eEhGili9Sa7TqtFVJs330ZVMLZwP3yAw
2mw33Ql3leRnzNSXNMTSNB6IxuR6hL5xDjExusVdxv2ufuyEA7sH3DfTHacNDoAfd/PffvRExccr
umKwANZKmNqLgbuspASMR9Me34SuxP3uPL3UaDUxA9hS/fC4WGQElkLddFkwicKk9H0s9F+4Qbyr
1yFwv4//XalqpC2i90YcUt6giKwqkIdxvg+ufWUKY9p1AzIeqU9BhdmEQJPmdxXV9M3QDlv8VXXV
T+a8D1aump6ilK8E31rZwCo2nU7QsYqa1zGLz93W1k12lQMsPADYdYhumuZz7JnZiU5iPVWUsuhy
zHngI1nocKNHo+4j19trKKFbpbimiXVyHKmrL4sJ/XKS2og1NDOGxnur0dooXsDYhHib2sYMgxqe
kXDH3NY9z+1wGb4oNLXsUfrae4mY22QbgOG+h+AmFOklCq85/9AwVJs6N7/lmnfO68Hfz4BDMiMQ
mBdghEaR2z0QkZBAUdVBlIm1+fA7XF2PJwCVrDPvgxgqAnhKXHfS5e4hTX2TSwKMjKOq5L+mL67N
cKkW8nPMvDz5TR8mvhqlrZPHqgJf54p2TadveUWfdW797dNM/73/mYgyjRT2/O6Ii6iH9XYzVkyr
I/fNpxm8ZRpRxK98jf9B2Y/fIwhPmnsNDV65uBig1O8WHGexJOz3SQJBzHIoxUxQTANmMdu1cL2W
wyJdGNvHqjAv63CbRhwYkpMFjAIhix+N32M08zeVi4m1ZYu1N1E+EVQl5KW0cm06sKHkMsu+QxkB
EIdoJB2dPMbYsG0OOIjoBB5WLkjUOpAIEFtVszUeLiowy/hvUUw179pyQxSfy0a/2DP8ML5NK8KY
GFRdz99xq7/SaPJRLSCF92m45qI9gg2X2DxnCvw5E3TwZX79952uxMvy50cWOc+pBrAhR8KDpza+
PboUr20qM1NI/E/J7odOaAIXXnQZ+Gz+lUU6rYQTb3QHLQC+Luni/Z/fzHmvUsFe5oJ6jPwgjgiu
OFp7LTTthiULUeOTn96ocWh7ECLjupQlgdVBbk0RnUsMjN512QkZD9Mauk2Ybqa0Y20vnWI7osVA
lgm31DvDxhHP8b7Qz6DN3QbkrtzJ+jo4ICnuvfAFCGd4RXyVVrq1Vh4NNLJU94dg/HKzviEmFXFb
pS3Ntyb/BWYeIz8ajuGhjlOJxKAyyhSVvXJawp4sRp0McYtZcLmzX8rVRhCjZw3OnL5sWCc92E3e
0lr4Y+I/HF8s/FBO+9IlZWTaEY782lOPANr9NFsjLA0JuP64IpXGZt0ziJIQcwLtXW6a13GlSBr3
IF/OZzygz0ChjyWxp7tB3rAoVm28C7oDxdqZmI+wTnV/0MO7sgmpHtUfdZK7QPBqFNBb8kqZz37g
F4LWrK8GrfX7wGzahk1TxvoeEK+Y5PLVRmX31ZG1CvqG1bWC2cOIl3AHL3CKVtnF7gXr+/CSdROb
zbISdwX++h3WI5aQpE3JnpPBJPUKquMqIUSh8snJ69h2Oo/q1yNQlNQL9HDEfMKAc5sRtpEVSXBG
D/a5+U9HxYwpWFZre5VC2Qiefeq6anikETIxX2IaR1lQv+7d5gBprk12FJKLdnew782wLZa3ILxy
5QfMF6G36E1jyFYVdsf3ehKB+TMdENRqC18aY0Jvo+AGOh0VtyUvEI3juP3bSvTJIM5G6s0DSoJ2
BUShIn0UBkYkW27JjksVgP9PzD6nvUxMrUgbcpva/YzI/duhQ1MI1HM0wboQn/ZB168EF/6o/XFz
/V6+07ti96j0NMR/1JGmTS/g4brpMmTWP67GVmx3xcwPdhcGvNVnKko5orHzkDk+qUsHOwy2jGjf
jw878qHAbmdMO7napIxnHWJsQrT6qX8n4TaFFl3xiLp9foT/C5w8aUA5HHYTsvS+ueqKv2jM7ClD
OyJJJDB0FtI007pZ2BJNWB0Pj7/Ws5t/K4Gq4zYVa5gh9pyxFYKYSYkB+8RnFbssY5emfKaR0zVd
tc/kRavuMrCPLHLRgct129fovzN5wNGcpj9rZj6CuT0/iNSoQZi5xHjsDp7mDnJuVzN8ASGQblNZ
rhOx9UdudfjoYbzFSArSny2T96us86PoyfxiWq05VPzm0EhR2yrWwGnuUWfitRYJ/yjRIvpTSa80
wl06t0manEKHo1qmbBt+NYdigupdvGA2ZjuYpJAnjF7A1RT5LgcTpdP1oXU1L4Dluio0aEMU7DMH
8J+Cqxl9CufAFIIULHsSxrWbtgvKnTaeNIJreBvztWJpR4OtLUnw4SGCZCUG1v2YrhherszGz4F9
wMR93QJhY5H53ToRoUM8vliP8UyV7Ss9HlpuMlYp7picHIo2tDS8uR40hk9zaPQpuoamn4V5e6wf
cimuzOpZWa5ok17bHYJ7zZk1IPXG/w5BK36gg0n0mvWxH8hfvYsmiF68tzAU1Tt3m2vpn2FFyN6p
qNfJZFRxv+ifPuYvyTmgjh27WeA6O6cxSqz5H/PuT6oF4bh4M5ZhxaqyUrG2ZNyRYbhUFvUkBBvE
xpAaOQHOCCIkpZT8RdQTeqtE53mUvHAcplF+xs853Qey6X5O/krd+lIsEap9YnypzSPVg9eCDdQk
MKwIKLiivpfyxV/CKAIgYoaIxok85bRAFIBHOIgI/ZrlRil0LNfRc9mMiCRNqJO5gR3nmGOou6Vd
vC4DfE3K3hoV0ezwmwxzKFKHYifowUTYhhkzDRyzwDGoqrEogmfykRsIqtecvVS6J6BwoK0Fjzeh
7dDL0DVtRs4BRcFzXfWj16KaZSs6+XtoP1Dsgw5CchPKbPN/H3GuIVLOJ9S4gizUJA2hNOveB06V
Z7Eon1sp+/u4L+W8vPJqlAEeep5XKyWPCQwjXQzo6Do7Uo8E5RpicH9G0XjRT3hI/gmHb6z6vGP6
2Xh/eiWfKTtFHfbsfMTKVgjD2fXjtTVAHDX6l6HJj3M/IgGBGmtFdi3Se7mLbwb6WcSmwXD93XIJ
y43NivxXnHDLRCRntNe2lEFI64pSmwkDUUYU2RIDPzhsNHdkh8Fdypo+5yBX6NM1G5e4fiVDcBir
Q1YMy0U4w31BiDThBnat66EndrOHvpXgVkvivDhp8DlUUhtH+a85qZt0mcmuWA7YUUsHm+TQARYc
JjvY3SFzNnbXbZBmsTu5AXvt5dNeZAn5eYMjDPXofGnHm6RPuIzJ4sBhuL9rwtQcG+0lz11tyZe8
jOM/ugCTCm3mZSI529JFzck3DkMXjrXL43hSmXIb5x2iB8jqk5fOOUfF6dJlORbdsWIgopbbxEXI
OHIJ4Aus4pzN4V5wttXI6q0YjCDuCMw5ewyV6T3ufxU5hQrdJFCYCxRL8SeY3pXA9ZyhMg0uZbby
XgAIlmdR1+pTANTN7jAwSE8+cw02xL15/xxM8D0BY1sPRAyj1W4Ie+bvSY2KQgmJxEgFldmPE7UR
qIb51hOGbYrs24DGh1tkZyfduI3K6yqk7ve4CoJZd3YdKZYGbutepd7lMpXl1MWMM3FyJzdljOmb
Ruvfzh7sv+KE/b8HslE8T99PmP3B7qIHkhqK1mGapUzmSDEa7aDYI+K18X15AisElEYheCwwt0un
tnVqysa4V+mRTeeAQFiJUW57bhZxNX/BHDf+iP7V//wTpmE/TiH9lASxf/CQY8h78A045NjTScok
zDEWUBIyULODL1aq9y8Qv1WdvxrgYeCML4E6uTHHvBONWhP3SRT/inkkMkKtL8w2SsPRjbCnFFJZ
9LSZxD/nly9gfbjwR0U4gAfo2EAUoDWhZoc33AdI07ToLTxxMxo8GJaYamz6TphIMbN8PGAH5JXY
WzZzOEB8qUoKJq0HzIF2Fqxb2JoyrIye9Xijy9xEXRIvy8UdKQtRr8LMUgsIKO9uKX+mbpgxi+/b
AhIYudaVi8EPZ8uNRlvvS7uENh/LZunFqe4PnKnd+ZnUCXNl6D4MJptm4BPCHQhEVkprH1H8uQBv
CL73na4AaT4i3Q27cxZdcgjImYs0Hd24X2kbpYvEx7kt3j9w3wXDTB8OR0MWvkYHfqfVE5rlFL3x
elCUB7un8fbvwLV3x1DGoSVLwt1gA46TWzi3N4So6EYEvICd5igg11ovve/lcyKmnwZcuSXIsPKe
F60qi5+OGSmfTUcRJrmitbvdxaDEovCfWuBZt5X4Go1B/oL+s9my2NqjcNOiocarcqYk3DYQdhpG
1guXpjh05e6NcfRJmWLq7dENou8CGpv0qG9mBbPrqxI2Gi/ao/rGpdFMSNoiCpi7mcrfLLUqZ6Wm
xVWT+/ZUdBDy59giYwpsgLSo2YcC4azwx4HtBQYBXwAz5qJZsDmbn/pnE+Q74z0F/AXc29gJziOV
k5v17IhCWuGy+G0m0YDrhkTmFH0K0z4amo4ccMMm3GUhhaoPBtPgblp2SMToMhkGzOi/8lnCRPmq
A0c9q0M/f7u/6Ky/OybV3LTWzRwy7ojrZM/ONsrZ1wecdC07Fc9UA/eJDDOng88GHlPC7CCn6WEV
1DWGbTV6lwMY4SACqvw5AlwWbd6o7J9zFiwqBVZ/9q9IXudFIK1vK7P97YjnXkD9ANdS2YTvMAGW
tHDQvBZg3Xva1VVMp0hcIXW/KEloPsX8DSj4z03H9I3axSptWYFqlKjfof8AAv7F2jPZyp6afhSQ
IRChFErXNY7YjAlAveigrrHOZYt5jnakc9dxHT3ZyitE6zgdGhcWVLS4uSdiFCQdK0FLmOiYv3oC
q8APFV65mA/yec7aYomp1nGsR7WZDv4+yBkxYuTNS+ErwKW70KcGk+8FXosF/lv84BGpy7o0PpC8
nSZVOpe+X6CVfIMHRj1U1iYW1odhIxKmIkR4rJs8GcayxHbE/m+p4Ucdx/r3uYjjipsAWY5CFU18
zGE9zGwOsz8ds0Vvm2dwDmNJrHFyLTneg8eazsXnTt61fw0z1mJ77sAJq/eskRajoQGQiZLDSkFH
kDswSNlb2k5gtOy/3trR4VoD8MTRwQj5BiFDHZZW4+7aVEOH+TpKd8CeEEBuOcBwAeD2FawkciOQ
Enhp6FkFaiRNom88ivn6/Hn7a3U5Y4Rl2HAA223qjS5Ts2+sXnM/225Slijtjwo96IuunZ/Q7xAI
kB7+yedSQ21oOzzwG5nMo8iDXvdjyHiwZ2RGNZ65fqGgFx9xDN4xFoZ4lTJRvJcQLpl+NWAyFbp1
obefMOiQAYwFd2YtXoIFzfkkSPkNfZi0/HmY/OHS4OpaYDhEWUqWGGmhTcmkHHrlMvFnglqhIK0f
UoE2wx3TTCe8Bx+OAQGHg3wTzOVz80zzHV0P7khpu8PHwCb3+oRQ29na2E+pB9FOysyMHPhR4ola
8cmoD9xUB0/eq7dAtht9ABiTaMNq7xITF6isJgHDDVyQgDTMPJQ0KUYjjXasI2Vh5B9gGUyuBPmo
DzxS4Of1+xiMc3Wfb8U5zYTqD4ylu6Woh2/6zRZMf3PkKAFISviTZW6yEIXUYwq1zc9A1FxvAF87
AUDC0hti70ScmoLb1eWr+II2eHFH7u3ARNsqbnjDFq7XovyFQfo90lXR7eJt8RROpNvSnIa+6+mH
SGnIZdhZGLIwFBsAKKibJrapkpnRxwG33sxdxEjwVfvNRxYLs0JIUtKMkqDbzv8TzI4Qi7DAveZt
t+PV6Wa3gBIFDfWMFfpj3J2/D8uxfnxTr5bkxyb2a91XFe24Vpio/pHl92JXUdJ5XzXhMmZz0Jgd
4t8HhaXK6Lb0LvmzhPTpOhbrfhcR0LDaoNsNHTu324FMEuGH4GZd65bSw5mc9uDhznsRgY0i1ZT7
875TeAAHIqpWA/6PxOqmHOuEtA4Gq6UM1NjEsFnvdBdhlhvHwlaGsMEGHfoRHoVrzAvwMGwEi0So
zrApmgo73ei4+JITw3TeaUXO6KWH4no+qbuIkWKw0/9CqKgUztX/zAsag/JvZoFkcj0Wmmu7TVHk
jivJK899uWBv7HcOYBrtW+p0KYk2eRzx9uMLfJHXGV8cO2ManJuJFJHiaaVhPFyRIMw7Dvyhz65z
umID30ATCj6EB2p21oMDe3CQEKmdOy/ALy6G0B+eml36FUffspdBKN/V94pS1rZTgOfScpRiSdY8
lnFGfjHHLFHfcrPEys0gnggWi0CPI463TiXWxUP9XB/hWrYMJ6CHUTGX9CanONWMvKZzNstr5tLe
MeArf2XfK3YNKcs3Hd2bZ3XaMx1D3NxN3wCSDg4rgYd6NFhgmCvrurIn4FHR/6PPW8ENFDx7iR4T
kc0YLpyKoUE3wtdegedT3dIqE5Z+8sXTKfIXCwKox/WHTeLmuDNgfD5QCh02qW0AdqSPtrAz7Azd
1IvQtti2wbZNBa6ub9QH7HEp0zBlEIkMomF6xmT9DlVAu78pycLrVRYnVw09JZouFgJpMO7+58FT
ki+6pLCevW75QvRwTAfvpxhbI9SJNBnak7xI1NKfpw3THq7b7A7Ew2YFg17uxeWxbU9/kvtStdwq
RHpSY6x+lvZKwzyJOjbK4dYdUKjg6YimezvwZavmWIueyN41G5246/zy5I151JSc3grEZ0bPjaCV
6JoW2R/Xn2zdDFVQr2nF7HE4jmS97fTu8eOyLOE7UUJ5cwqPGaCLIvAI3reESfEJjztnFj0wSVgI
4s6MSyeYUW8/HHdDS9MzLa06wfgItBE9SP6HgOPrtO+jPAAH+pEjy4XJi8EhK9uvXtadBmvcEV1n
7r9XzJfhulkz1aF7OcJa6XXm/5OR1RxsuggeJE9zEy0QsNuqoQ3ce4UIjMvmF+XPDpHI11iF6hN/
xnsT9fHNXH2xhE/ELulx6hoe5PJH7Tt7LhCyGqdcaFuzars1DuZYjl7Nb1O/TcuoDRxwdfuuAgoP
8CYA2H8eYtwhzq5N+bQdUvqxvxqh7s34vGV0BmaKcIt/5pBpCkw4fjz2QzvbmWycZO/qi+v5wk8b
HXGsIiM7f726FuNGuEzrMlCvPdxNtnkUrk91L1yW7+wYnN2N17Xr63B20J2jOEK11L8RVuA4UYL/
r8wXd2iR/bkp0RfxLZs+bmSptBKfhoAaOL2JZr8tYYTybhpdfE5slxd/mM9Z5Duaf2ZhPuZxeTfZ
pSpAWD3DYQVkmutn8imbJ6NH0TDcV2czu5pe6UeVCZ3AEj+gOScvAZqNYIQl9cwLMVkhkBeSDr1p
nmPnxBJq0mjNf1nTAayc6fam4xaAQ+6/3Cy+4ySFO0nj5+tW7FNpaCZSsjElwlKX0wSDBEqWI5BW
8+rXprcZKSlyhIFkgnHb60EfeXm1GcQYiKbn1OGM/4w0Sg4oyvMSoSE+fB35XjHcRf0yvxVF1ouN
E14jWbopimQXVcr+dDjf0MajL2wy44L6U9C7aRlWyYXAOAEfgU6vHDU11IW9awONawZqIBSUljH3
W9TsIR3Q71zBuZGdXILls9Ced0+xXpu2Pw6N26z38yFRPoQGBV53tFV2m0I4ObpUXzu7u+XTr0UM
GlyzwTlpG8LuCnMMSY/JwKLqZxf1DDF7V3zFlrGGCgPvrHRNOVA9UDMAOt19Lm40eM3HtE3NxUtv
ZRSXRxFxot/VQsyDOsAIOSFU5s5oOLxG8w2zlOEZOZ2skoQHOnJEEL6F+1DCQ1xb389DOzcTkc2b
ooknt/pOzGe0w/dOSvcbyTA/eMa3Rtk6j4GnEUSEzw7bh3jU9dLpBpt4Wxziplf6oG6TqPuu+0Co
1gIHNJAaWABMjv3crAh/7NxQrrFg6VSqM5N8lAD6jWLJFdDn76af5s/RC6cBRQn+jdGmmadtJerk
IJ7xbiGRcu30CNU6kc5k3tIENNvpeiDjrD/5RRUaQgKvN0itDctS6CS4HIXirU1+G7DC2C43bQc8
QMkmw6e7jCiXNwcgL1i07/UaPOWzcQ0XRe3AGkjY8ELWY3iulQhtUANbmZbyDrh8x2o1ecx3Q1PO
tnG9lPFJFpHApT1XCDFZSUhpc2HzHTArCSGAwc315nd8OB2WUgvC4uLTbBLBt7DkaXHmw9daigJJ
AziiY0PHOHOVocbsP27XhCJkpQ2aVhhKsg7E13lWHYYP5LPxC2mD7T5809Vk0rlJFV6vH+IScd+b
dK6nq1HVAfS98HGg3KZVNOMxT5Q2z5AmKH2oQ4ZW6EovAzFIiD3byfhx0SO+XeDwSkSyREYxhhRC
dhrUlhdByWAoEwc7ZBrK1z0R6wMbFQuWOiugGFmsvf+EGqdgtydR32ffblawH9bm/rv+B56Pp66A
sG0afM89OC8MusL4gVYpb+blfAhWDkp/8cYxnxqeugV4zIMzdG4n/MA2pg6YqXa2lgCWrT1g86Gh
y93mJ1jIsWCdkVLJE/mDtiURQZ7xCo5CZx75MFM+8wy0v+iuY4neiZdhx4jfLfWRJ+WnGa3X7EYc
0Mp1R1tKKQu6XOitK8G0vUrUxa3Iy3G9OlMGtgdRY0tLCUdIdXLnr17UZ0mnGzWG01O3kQMKIu7o
K+VGuNfOFDjW76Fv4cqNBU9LEX6E9qGYKDSjywEyUbNIl3D7ffUcEHjRgDg8M4PYN3xh5JjH5yyL
j5iAA5fGKJVZ/F7eH3OVR3rau6Fs4VwQa3UPKr8RAGckUeJ/XLG+tuSc721ryjmNw1gYUc5/pfEw
+DRQIpA5dThCkCzyvSrvKo8HPtGIOgawfCJHn+LcQBKVSCVpiOXHoH+vlDe/nbzFri+aF5jVrJCE
EBT3AihZx6tcO7rDH9vNFK696NpuI7GCv+EpIq6bFmoC7mlIFXCEEV6FXCpX65hVXPvnUfBaPavh
sJOIJ7tBC3ts7gAExTZgrxprtXKrFirXixFvi+dwtDHiSGz3pure2Ht5/5dlFUScTj5xIfimUUuj
I0622Ne9VAAW9leJVFKiwwxDMSNOO+D6VeCrI7ttKqefDRb5q4/fPmleE3GxsGfVcgISzmD+vzGH
OoWi5VdnS5euvo84CsqpiLNEWC2vLFnuVSt8D3Y1G/gyn2F7XkknNRaX5kN/UntNSU+eGSK63sA3
UaQ4nycWYZAMiouicq+251ZFRWLzMdn42fVJlTjfph0m0o8O37mM/G8hfBCoom9GCaE3nqoKQlfD
A9DwoLQDr8XTqJaSaDlQMyJbTewUexvCBS+cmo30fjlKMQQQaqmSViWey4ztAqHU2W2SKBuFNGzU
EGeswrDK8hEtk+SWtHAIGA7uZu5hagjc+SF1+Jn1uyXBVq403RquEJNkbtIn+uqslDtOYci05ug8
dVhmKqnM4UL0tDtoE5Jp+3Br5TLuJAhQleGZ/ZWb+9DboT937I1EpKHZFYMnu361O+kb/oh9g7oz
/jHGiqpGods6LPYvgcKCY9QVQNx7qZV90nayKMpHk8zBqNlgoKGpTNzVEt1LjnuB5hsbosIN3Xyu
EGtoMv44oCrdTY8sdnF341vbDWuXmFxcF/0ue6TGq8bKhUh/LBrJqpUSYTbcbuN12XYOpf1T42/Q
JWvYnZLrrYThCcASdKrYh9FQGRApffRDbsCMA0k7iIzUhWtwB4GXFhc74QDk+5cnCheYN1D+dVr5
tijQLv6Z8m9Wetp1ekw6Rci8u1bbmdxJq1ujQMvG0uvWAGonxVYH7sunx/pLoFeVP/ShLqMzjE6O
eUGQ7/+djFlR7Z0IDwkZXqkFyVvcN5VEUD+Ib3ZWmhUII+nGtayCoDGGAdvRrp70rMSr6xzZrH9X
LnVRAYO6z1QrzFeURNS8WEm4VbHtCKiU1wzcPbA7+PE0lxqlp+73FW5RBO5ZMhuxSxZyRCeXPeyc
7GgBRe0J7mD6CxbH+ZQIhmkRsdV/BvtUX7nr4/+sVpOm9VTNcjq/hkuobngkk/iscCYJfx9ZUGL0
OrX4Bdkq2FG1rUhDZm9gH5pJXAvVpcFptoxgK7fRiLEbfR2s8BwrubShgdAf1QpnFUOuFSSaP8LF
aUVuNsM4DN9U9KQnykEkD6cawOfOFd/D7o/awoOtV1GO2G0LwBw8WXhRzs8nxdt7z97xVtwhIwBI
hR+hfUTF7qhTe0fU+HC32Tt270GNy/rJ+BUJA++qzRINpQjq7pYOkUbpiCwHsn22WiEbYMjRksUG
a057RDWQFyxCuf28TRUuyG86k39+L6PHnmocm8QVQ+rFHXtoZAu9+W2b9cOEU69Las8Xlc4dYwpl
JhELOA4S+EmaEupnBQ0jU9fnAOkS5+EcrkYKUw2nWhc1/jTvushljdYJ2NqAXqROrfwuYpZvhJ3Z
ju7OjAcTMCLLbGl42UQ6UdDbneAmAba+zdqUlyDiAMqO/7cMlSXfM7VHdTZ7OD8yVkhJWawV2hFs
Tl/Ef8+GIQg7syYvSLFujCvx6DYmJcGTXPeIc3/R78F5oqOIjpbhTDe+Sn3wJbNzOqGVQhu9jeak
J1yZZZD4I3CFc2ip2WjI3rKsD4otld7gI3gFYYn8GHn1Yk5yQU/8JYYoVO7kZJVvb99BnBUYYbjT
IG31GRwH8hjnrudYtlsyFkRWpRG71GWFykggblSoeSZhtIiN9GaRKREEypgu5ecOHQcNvLmK487e
uxlpuDNHORXIBRAYBpvprcQvEP7TkGvL4O/pIj3wRymd63m+2WZbxUXABEseHQ+jTiUiRWJrQto1
rQOEC3+vUJ++HHngY9IBOMh+9WRWjOMJljCjPM75ENevn4p7B0KP9NS1E4RarvTDc1vjb5pI6kwK
Jq0yb8QKKCpxaBUj39V25iWLFaOnfbEpxOZoQqbe9FUTbhcs++VuNZzakWzIvheQQFPh9NxqoYiZ
03czulhEtEfbH/+SDyuLPKZzL4DhOGjYyMZpQma2FZaynYm+EKgWwCCfb2szGrXIPJ01kmwWec8p
aTtK3SFZYwRxBb6gRUaHQhlJFiJnfP3wwtkQYTjvZ7+jAC36FvoNOagkicwQCqxG4FHOwJP0q3Dd
lcx7vic41PRIqPNzY2K9JiLIhCvx8tOvGQBVcoysMWpPyopd0jV0hj7I8EwW0TccqH1GOthbdbjD
Rdag8KJfO2vU/6HoFf5W3oBJ8/7AGIxJQZHxZpVcsiEpC++9yob+wziDpQClZAlZD22cnQFHiE/n
nyV9Jqjbonxjv/zTw31vhHZPksePQDnfMwH1YIIYjyiMsMx/DFKXTc9i0GsoCHUfT64PlYEAdmpJ
rBel0Ge98PYrzYRjaovfXzludkQZ1DqcszbWoreW+Xkj2fsExjgvtBAqtHTaD/PyzHTt+eyC/j9o
81PH6khdNXHnSJwbdWvQNubAqvVDA65+TbSmFHYeQ7fqJIVi4Soc6pNLrW2kpUFd3YU7mJk+in/Y
LXBI97+tehfN7bKRnsA8OxFZ7SBsfWkdFCUimBZWZ02aIUg+OZoREe+JSkDlz0gHiA43Qnr1R4Aq
CVkjp0FQOdf/IvB78bLigQV1bGlvfrO41CmLj6YCLHFgiEnS2opGhs2WQNRIFwLRm3OYeMfcOzvE
6krPPhz2wVxGuSfouCeOjV7b1TEbweSdhZjn/HouB/qAP4ctq27s/qtpa061yE7pSwa0CudT/vKr
vGP6pzZu3bYuh73eYLg1i7+fCX0z038Qep0XjWpEqleWagyL8Ccv0Kvxu5m65ta5Oxhr3SqdMbNW
54EQM/c/f7bjFAMTS3CatGhOAg6bd18w/uYg0Ac6ggtu7GjmvJ/9ODbAatgfZreIn3aMTR83cq/G
We3GUWvoLnrskznGRTRUCMYmpJ0O3opc89IjVFoSyrTeQ/vAfthKMWMXOcLQPLgidwNTIuqYYVDd
cna0p8NmPgJNk8gHa8ukfMeTd7lUixSps0SpdbjF9QYopc4l4Pv8SQUU766+gZK1uqrfmDnTW159
bbG8znepJ/EJsFpKuzksE72X1wGteUGPT9zTxLzsKBsbl+72G54ZWbbSgpWiX0oB3MHwNiLR/UR4
Xx+5/0g5htDsqmsbpRfsnOAkARaE95KfjTNE1IhEwN4mT9znFGtq+VqC+MG4n8Tff1HqijqJa1oH
87whjZ/3Ay8UNFgpmOtmOohhXae82QrLJ2ZONtdwvCRJWzoXArdFUfX2brW8eQo0AzUpBjHfs/rd
NviQji29OBQaKU/eCGq8rerKxPIA/zt7LFwcg7y0RU8/s9twzhh5djwMljMGw18ehk6fxQr/6sDr
Ls8aa+d60bWbBQ90AJvMNZkOo7gjLlXLBDn+v8P8OAhWIPpoMvKWNn1togIH7W3Er3iuzvAC9VM+
R3GwP4kvofOXwV+inKcrR4Jq/FC0SnkOJG2TbwogmA8LdDl9kaPp/4pb/HPJwnD3bOklL/6c7p/6
JdGkF4/4iyc9lM6TzFM7GkBmFmOE3kSvmC0Pj7sAJGnmcl2L3Q/4fNlPot/vLB3vjXnBsSr0fJk/
qx3w9j72S10ej6i1dW+9jm4iCiTqZFVL6usHoW5J6UvxdViZdfLaK+iFAYzEE3WmXwcEp+py8o68
02frjLFDcGDh56O3NiFtF2f1K3ke1B4Tm6tOmRMu8AhfsxZKSLsRP1AH/4UASzZpjoYfGeWT7rwG
aFPZnTQ62BNR9/Ev7uW73f2DBRMKjssAqW7blxrgrXhb7MBiNrX7ttPpK1ibJUKmbDvrsMWD48iH
krG68LLKnaRSyOlFM8WXZh2CdO+X0a9ojEhtdrv9kdzADDnaJXEnpY8xRTrMc3E4sLY68Y06/iXs
USyJUjp/jpT9rxLb+anPBPSQMiDFHwAsiAXO8VEMYWEe6KBObz18aXqNLndgskQY93/q3Orptvrh
d9vPDU8KMo9M71qFTipf4fz1Fr7TBLSLBEoBaHqQ4RXK0bHZSEJyfQouVREF1SPyLChXtykF++bE
D7hEp7f/ZCMBymDudehER6TSlPOeDK6R434W9Mo4khB1efin63IP1ro+aHW+8TpqAPhKADUIF0Hc
rNa8Btvg/HTutHIGb8oC2F3/G1pQ0mYiCfMGNxlaguB6yHfeiT6fAseubo/IauTVytzO4p8hUgJs
4BWD6qmioJu160GYNz6qBd9u1djKOofKjjSwiF9eeg4BzmM8vJA6+Takz/SzrS/HPNY4uBzvMU9a
j9lpr+jCuMUpCjpzFtu6cJewWQXLx0nFIWM7TyLS5wISHokBpK6xF8wmMzSwjWk0D2XFjSc+d7py
8HTi/xdJGw0KBQspCG2Hh/p2CyGlY3kdVu6fE1+64LCdguTxWAXiFd+uvoMmA5PU7Eg6hlXcGURm
xt5wI188OQMSy6PmzHGIlmB3MfUYIcp8q6Pz7xMMxW+7OXxaxxio4CTJ4rESlF0JbpmiXWue5dkZ
jSz8lQcY/aBSjbSt32kCCCOZEb/3PAw84xF7OEs7MlUEA/JX5580AlhuUc36sG066F8KicX9HT8F
Cj3y2wu9lYI4u/1jL7owXpev2DGGQKwFDdeAlc2vckVZHRhDgo82CNqQh6vlWAgDBudLVXkATOBn
AUHtS0GZercTT3CyBVcqn6DNT2BzIX7kqeyp5eKLUjJxKBhP6AYi2mNbNUtC4xg9FzJU1q8btoTw
zaGjZZqyHflY30JTNE3WwemIaF70NmQiF04YI8H+f+4sO3I1Qg46BcvdIa/UlwedZttcp/fo+HwW
0C9cK35eavqia7cavMy2Ch6BY294udi49VdV7rmf6w7p2ULAbOnEXDPJsMoU8tJttUCsYEeDHpeg
ah9zb1FdznI7nh3rcYDxX7d5sJmIwcQxOzkvH6e9Dg2qMPjv8Oc8T/rAid7XDqEaTXzuhvfwSkfS
2yn64YAod++yF+mkgsNvuoFqSNSjVVF00aB+5LKlgzBvHS+SpBrC1xtlrxETCgrKRB/g23NbgkDb
S24MZRIyGOfnUlqS/NMI1kEt/k8pfqwFUehva/cpqQrEOefIkFW6U1dJh9TP0yfCgAa80gQMycBq
L39KD0No77r2GHV7k9o3su6mrqXpkkHGSEQ7MHumPv8f/tBvvvLnEqtI4vrw1OJ1MwmEi8Mu2oS/
QaX8/DdPrTsOldrwv8G7DB3FHBKxMJe8PD2/VvLQQpkGo1STiGQZvvF/0BHsqr4DBabA6WR2/FyI
sqKNDr/K/Uplj55wy/2eLO87guRA7JNngk8MYGjeMSe9AT1n154p/mxeIZEdnamnlYJ2rD7xAofP
h7F2QQH8t5DHj0y4RJALyeIWVLtuAkNESsFvPLX3Oe+pTS2QllbFPJ6ubapEeovNE+oE521IMwsF
w20euQiNRw+wXxaw2MOfhB19gral1CV1iBn9Oe9fEw7xNJ5gFoj28ENICm2gBTX6jRgETnZdTL1T
b02OAotZQniAxLp7SXp8VlttH4LZ2zMgFyGEYHzAkrx199BNPU0KEWYEZDVqkOUuypKfACOTJAYM
9Ll2PxyZ/8ITOiKO24fERRwROnVuWQ1MM0qN+5rC89WQDrs4akagewrrob4QjG7zPDNujiHFS9i0
jcz8UFrnHgZz7doemnN7+Ro9ONBM1cqWidI755SQqjxkmeer2rLKr0rGSDEKnN5ZbMPOA7IQY1uF
nGCxw82Ox7QpXJFzdAPrxT0/ruv4yjX0+dAB24/eccfTgZVszK8PU0E8WvekLbb/61hMCWIf8TDv
gRJcUrGj6IXRjIt4BysFS/gi5ORXV6z8jn86CZllSnql43HsUK3+tnVusxL00AaLDF52l8DBbNYM
pUmUeVFd9Sgop63WLuGzcUAp4oR2835BI8aonRsa4snAttdqEsI37S9g2/XJnYJ4BG8sNrOjp82D
6fRncXkZEOTHEQtnqg7uq/2GEEWKlcjFWKkdlKYSmycJkgJ87ziPiIsYPJ4IXsXltgkxqfIQ8yRW
lYAUl0fChIPrssNnu3IJ6ZHHzcPdAPktUSgM9bp8yDTocJNGfOG5FbffzCIz25OM0DW1yxglWmXg
B1rmVXXFzWgslynRn5cFZsXLSV9HZK4ISKjCyC8KBKFXXW7cAZWSB9cWXLbNGUaJ+p9z/JgSIplo
L98xeS1pDBZ0zdObXH9AuNN/oxd3xau7oH2OHd6QQhdRtu9XwELK8bgOD1W8ohvPx0SJ9IJNdCGi
Uc4a6HPrkXntkr5bA2H2CslYJH+TFklsldyJ6m3s1O+ZjjRh3BTBONS3EimMO1wA0hFuQ4/02ZWw
PyVhLs1/junuG5ljv8asyHzDTsJpI/SGGjzzq8XusQhNwF9L80vhR8W12bY7rYUJ3a/e+6EZ/Znp
/HeqcRjbITEK2Uo8dTJy/dJIikJbREtn4AvLBkbfnCtA8cwELpBAlkZzNf5wR8ha9/ksGGMzphzw
mDKbmCcmpK2iiePBUMHhcXAm8Hkb1Ry9VJIgPXmXFwxPvIdPN84cwtQxSu/MAkrGHnxCWupSyEy0
H0e8VXQFTfQ8ZVg6WGcVtZVHDjcE+qmjZGpoCSFC/TB2YutwGR8Dbi2IErdHTLhOQVvWBYFB6f4a
uK6cZqppqTcmFMaTRwpNACqLL3dsKANkAIrsysWi+WefJzHNe/QW4DNX8fq+FDkTYA4aLPl0jDLF
LmYpxCsmrZ5eZQ3lx6tI9nOJ4XCIpS9tbJ/iGxRVcT2yXeHpTQmNbafEW8OEKUKz77H59vI9WBxX
PZmOwvZaXcqoCL4RNEj0xHRhPmBmdNpEmArhi6Vh/HPyVxGarGJUkcck4N4idpIVXkUY9xdcjvpi
UcA+14WDBU5OVafM7wXHTgv9RHrmbWQkM4IDRppTaS7kkJDRVnDS5yxh/xQwoFzUbZRRtwrYhzP9
4YVW5b2i923AWkjaOzk8rjLYKvrMmwL0gFyC7Q7zhzczfn0SzNyk6IbHtxlTnaWaYRo7FbkqWDhO
KcmMCS4aS2Y7wW3SK+o02DJMgspb2AMkbTYea7r8Ui9jyfqaWEr5TG1BOpe/kq1HuEh5yRTtD1ye
s6YELp5r3xIRbKHtG+GyQ2gUNpYtrig8zWzu8BRHWdgwoq/bf+mgN5raVIP7yHHP+/ptgEPlooMK
9pfURVXYRTOk5bJlIJZz8NtWcywHksJ95CtwkbBlUObCUe3ionFsTadP780Z8vJzGnPiF9lgC5Uy
zo1EEi1Si2acbrLKEzJx7hvOew0oau5mhF7ydySmZSrotBKfQIGnvjXtMetfWftPl84FF8i30EFX
qZ+PMeTBtdE2703ix3z3ffu9g2m+qZ99TmOzCpRrxQg4Q8csC+FcINvF6jhUzcd/uQROoJJFAh1K
IteK39reC0wqOSmvtDdOR2Ht7xYh9iKIn8jAxQQSue+qS3l6dDcIW8aJKGh0A8+1M8VitaK1Sb1G
MGb8liZgSZKrvKcOeUa4obmPlzX1dQZa8ksfeidlXGCbKgbxaMi+anqbs0KzgXVUuOjcW9WZbj0M
NYcIb5ul4jVS6drs89rU4+gOVSjDVNpT126KbM33HbcLowMfujkFbcFVNR0dqFh2qtfp4V9ngvrz
aWcQ3rRZJmkug0w8F3GGBv1MbqnpldNXct8+0gBrLGpQ+0So6c5QGy4ebYx5NSxZTDKtMq8Muk9e
bmVYeynReJnzHQr4Wx9w/v2C8nzoFzKVv/JD5Wbr9IvAHz9L2KhbpYdHGJ93qqaisNI2mWEVpBxR
1x0LgOfJkEi6/FHyjKDfK1JqGoFR7TYSAKMmaKKyWT0LA1Tn37S+SKS1jKwjZB2bdoYJu2kpO1fR
vfaUwesS2A1be9yz7tA31zV8C9Cw05xtCmMSFAAqd+9KkI4CsQVgRSNujuj5s/3rV9NX/iSnZSmp
WSn3TTbd78GwVfA+lCD1wTCqSfadK5W1Mtxhh4grQpGsa6osLRUjPNr46jQuM0nV1NMDLbOpkvdf
zpuRBLGJ2BSs8XaxtIK7kuoBp5h2rxV1ZwR8gWiSZ9nqSzES9DQ9N45EvLHVqd6ynQp6GpqmfyUl
4UNq7E6H+etAW5lqPwcx0qVzgzrv85lE66Wz/Uf8W0pRXchzciDxqaAYC+hvOe8y1kzt41m46w9/
NscvO1nwJJonEokdLgD9MW8P47l7+j/SJOEnA6dmMPVgIi9T8kKOdFAxuoF0HjD97jgwNmg6tjDg
KAbPPm49QrQ14c1THj4m7KTFGo7xzgrgeRmr6NaCzHtpb+C7KiWb7YOk9HKL7/aBkqElEafykxbb
7ScBhmfe09Wg8YZst6WMs4bPYyuHCXqBt1pbWfyPRupOBW0wyaH0buxgmUUpQVZ/1MUeG8wZa9cq
RmiqGbgtq2Cg1KH7AU+8Ub+qSb+2L5kQ9VM5ETAADiXZtJ6nE9DBArh8cszDWcrQpTN4e8CoVVkI
tFJI2ioLKUBfDfc7WV/NhWs2r5W4uANeIVt82cbS6tkGGiQhnGpQcQ/NsMOzBgZ7OfzOoKAYRTaS
wfXBwyy00IzzpYOcfXuUc+xzbO/BF7dy2Yiz3/DFtfyBNRZ/eH9FBITzFMtwe7abw/ZIcUk+GP9/
iL74nF6r6oBtZx7TjPf9fQgxmivG91PQ3jlDJyqXjxvxAAAuYWmEKa5ifw5OMInj6A+NUnNO8ft0
J4boVQ5gYKBvarwkYkIAIuDnSJyQ3ImPRXY6fHR6MKnKksNg9pTOAqKxcwrtlTg/z+IYa9QllPOH
K2Glc1mSvXXe1t/K1c1YaYLEuARO2aO6cYcXqSAcLsFU2QEEMDUshjcQ7ltR7FnGC5/X6nkJDg6Z
6JDZTTLOfl1rfAZ6u4bu/Ifk6ieuR8nCdOYngT13zIsm+lr/oGwhRsWfYRIqOJDzi6eWgEo2630O
g1CgOYqkBcRgnm7VAr2JywYQxk7llRGH32/NWxsacgW0wbWDNE0N6KQZt8e7omF/21XHbVFLBb7+
3oqSIIt6WCrNq9nrGF5nZjgMFspusBJELCHAB44x9ynn8Up9tcGISVdUQ9vokx8Pn4iiZQ2WwQOI
v9YPEaCbbDIeqmaE+WPxiOh1VzleeITEN334sF16X5YKlSWii/hElqDeVX8Yt45dhAt4KaQdXsXj
L2BsLwNewUNHU2GyPA4+7P3Q4Lg4Y8YWYSFQQ9U4ZbBPJO6xQoxawF0XKZR7anEXLlZuPERly80m
p7R/JL9/38uv9EKY+tiJcMsEPIxtJxZjEKGwfrpIzmimhcALMK2JaS8a01T2Z2+hn3o+b2KFVbjh
MHu0wzSuHea6FRb3Qg8RWkscPTBfw7OppKlrggSRvrd39vFhwcOA9x7FHtoNzL5bNro/C5d2Vgc1
Ml2Wl1Ygrwq9wGypPVvn+KJKk+3iG82b4Dh3egun9N/56a58HyFMLCVdZApQbscW11spx0uONVfd
PhBT2/JutJ+cJ4vofKw+h3BD8oAiL4ZgdfiR8dxsms13EM7qgMFmevvAXqtqb6rMf8WlNwrOnl6+
Eb36SuaiHcodSSqtN1qqgEERDsItT6oNttObCP3b6AsZjjr6ovZ2p3qK17PrKGXCHhTsnOLIzOwo
BMzTdUqlSRjfl8ymuEzqxNBOBUsB2qIRpfDL+WglgswyHyW97tMhW5p+jbxoNmiaEl2G1+ufHKTq
F/a0Ih+EHVPvOslGAkUeom5Lt/HXqW2RPr2s4H83FRiHLcIW9I/WfJLcuyNmowpb+s9bsux+T58r
4s7CAc8SQfTF/Xl/9VoKKy1uO8PnOOOI13NyNFyn5ewO2WMy0yrYGrK5JBE8fivWZIieJcYk7Cjb
5yTU/WVowHwh9fseqwfav990G4ezTuQSkkFwZftYDLgY17U51htVWeIkvq8319cSteqkApZtNYi2
P5WLN/VC1RdWSRs3Wli0Lw9HNbqpo6o3Iw9v2j7+3O0PucUie+OqvFkRRaAQm3UHcJi0W/WClacF
P0YmKQk6A/0B1fwJ2F+IaEXmTR2X2GArvhE5FI0V3CEtY0ViZZurHxKGEzYXzl2LcX8ZBkdzPbJC
VYx9mHq/X8ydxY+tNTPzFXhP89OumU6flTlHG+UNm2AG6D++Z8xm+3ZfBZFZMPDvql9vatjRFv7o
P+C73X5de+DriTJ1P8+EDpgzW+u1kc2aIdPsdvwY2W71H5X8XSxd9ETTSr92IwP0PDhjT4U8N6/U
jW2ty7tc1KkZSnMnNkrg4rnzqH0L8iGR0WVvWDliewxMO5BH+QkIpKvqGzXvkSDy3Dy3PMNhcTds
o6lvaeldyNJd9D9+dHfPx1h804cqaudNsftCf6ZS3eYxh4C9bnh0bbZNFjAZfdwiDmnFtWKCdXr1
KSS0HriWtfgyK8ee05T+UFK3yL3CgOdhnPFkMh9aWxk9xiALiQUWFV7quB5srQaEYDVjYOU9ktiw
9TeWLpKnCZIi4VlWGW9BkT006ctnR5zjaDVHWymQD5k1e2yDW4gxjgscubwAoFN4oSWhZ+9KlkKJ
YfTmrq+U4F/qR6PcPEAnYvEc5qZ+ndlZjo5+9cmKlITbTXAtzVJunXpa+LMWw944yDuzdvZR7UJV
Tx3pcXsnzIaGGpTXuKQY7+yIXrzE7q1ZewaD/60G7tyd2Rlxvlz7A/0vTIc1971co+lX0c/dqcLQ
GACB46Iv8/SCRIoQEFP4BgelNQDkgV7mRudHW1ExT3wdfWTAcIVfguyRxFG2W2Y0L1H95o4VWn/l
kPtjQwE3CFNxYqhN+spk0NouJoYQqBYu6uGzXDmRd3+y+Gj0upojAjtEsh303EL3sgJpmvWiM2u1
dGI+8pFqky3X2SYH06Jt0MsjPwTp2m4JHx5hGAdNDm5+Sct48Jzaw2ydcVhcVlOH8Tn2DsT1GDR0
Jw0OcCa8+7xj+wU4+CHUiD28rWsF8I/o7R0vox57rfN0IwVUW5U1wGDQMpji9pLNYBrPT/0baP3W
tyT4DAQQ+472YwnHgJKL9L0ke63yqkxnVVDnyXhrdCqIzVw0yglVw3B/OhnF3Ruicj9JCTj5dJsv
oCy+OqiWrwTLtvI+zorN1WMBZrDqBh53COJgcrzc0AutqGj7N2G2Em1WaLUrpa6i/UBwcjM5BNnE
LbGzrlxgULkgHHbOfyJmdji5o9+CPYxAElrv6y+kk5kzXQBrcGIdWIBUpsVZFyEOqYlXSLyqFola
6GEY1RE0dTE3MzR29XBsDbKFmm903HhHMVavJf385WyWhwtSUb2zPW0P36vRNROizt/vAA0kGe9b
893WOlO7T59j2wMQsk5NEw5NtlGJFtuys2ZbX+9mXvfBk7ip7fNVYj59VzNTagEXCbwPtYTit1WN
vjzfYoD57ilQtxbR72m2dqNHISm30qAM6HKdfSpqYC0EZu4yFG+To6Owbi0tkztxUxuy/ymChI1E
Xq68LA2LapDE1GId5s6hDcLyI/RutnKMYyd9EIQwGHCuksPFlYy9I34CQFG9Ra7T6+NjAGDR9f2x
KgVyCNbILvnhFMLQe/FPIIDDVtxMM7Ntn1rI60p5fvf739WV1caTvau2WQ3eTrGtF4MO2JCYudjh
91HoWAE6cNRMUw627m0UOBufFR/ZBUAwY2IHcCd3qS36eJ782oOFgHbZRpZRrGnygu+MbU74fwHk
aBD4wjzvS3nS3dh2a3rR0yVKz5Tnc+W29IbtXTzfhKCEsm5xQ0MqMmr0BUzBymkY+n/mgPLqBS+j
ekipEwOlqYDYgDHPyzxdpOiUdLWLAmgCTSEhMLds5tugJ083kAswg17Wc7GYNjoExfZY7DmDijHh
Q380tf8p+jJ5vjyty7zCcYpgi31owL5gED8ZUDPRAlTTqTYGFSMiT1+4Zq8zrnowkVGXtpgbQVcv
2bri7O6zVuKoMzSOfgpn4Y2+FXnn97JZtAAwLahwSfbKdhZb3Pc03UW+MIskijbXQDSXB9+1QA2b
j6RsCn8qwub+0XukPJMP/0ectv/7bLxkP+/hoABHhmw+fiD8EO4/OJEx4TDiGlISJuMJiGUVWdKs
LkBesos9uTqoyotVwsIQQF+toCJw3fCzI+hCoOafyhh6K0rQphDib3x6eiHQ210vI4IzKl67Xilm
M5buaFieKWZEC8mddKvHWQ2dx2hLVu+RhgoWJprLxko2d2dEvucYXJ/JinB0GxYM1CU8loSvQrEM
Anv+DTToemF5g0oF7vft5pCZxyjT/nDr0K0Bc1osZekZ9Es0c5pcneI9BjkrU2OeXtyrRB6qcQyt
3U/h/fVnbRQzjHbFHeDyG3uCad5Wn/DKl+l5rJs+gfooqnyyL1UlbRw13dPNsHSPNeFXAjWaOnbq
VUrLEVb1rGtmJTbHVKU5YcovSRYsuyaMNLsYLAQE+cf0J4onYDOyZ4dM4GgzXbo4Vb3hJC5s9BVw
FfNhw2ivvm7sApLa3WxeMcC/lJEK3WnpNWmaRAh7k9NG7Ig+T53vb9eVIY3Jm/zWWYgy/OM7ul7b
zoZyya9ybV2jpXywgy3fSdCXdudzevYnuzB7xtUKw+yB/xVMSTbw/ou8pJfJ66jg5clMGOQSCjl5
cAgQoS+5xQAutp/APlIplE4Z9q57TqICLDBcQweA2houLieKRVmASrJj+sVbnDbO6YcIn+j4KDW2
e7PAbJD4WjStknKu4l+0QGXFOq/xTR4o0xvm6k7OtzP16netRlsjAl3nLoZSw+f/HoS4HAsMssKz
O5kDQS/ifRLt51rW6GwMHZxdintA0TJtbMgzJcYxQeYdyoPz/e2OCIL7+trJsGDWUpTittLXW75p
2qeO7m0Lf/wMj0mHWTjA5hXKdU/DuhloSmtPiPKXL9Ym2Exe594ttVAWzBf+UP1LEIZakw6iVfAA
ZcFxoZty4CHLN54Ir6VvrBrBCRpDox5MrlP1fnNbep4JmTfc4Sq9Pqwf/hugda/kZeNb+27n8ikd
siY/sSErs9D1wdVxoT0ThOuzLDjwaRvTMUfgasF/F0cD3FzhYLH6cmed87v9UJEyx+jBXji/S8f3
c3l0O8z35RBC95NMAJXsxbklYn4frb9dGPSnLrZ80fhT/763qrU/Q4S/2rRBnvwegsiXBB29NRwX
4oXWmaykyLuWTi023WJGxE7ysNEW9BQGgepmSWEbgXSMzUyU45wQpq01FzwbjoBoPQf+uYXUc8DL
Gxmu/+fY4gf5RdcoLn5yv6ixjn8dB1x9qzCkEXktX9Kq0/sHL+s9S1M05YM7Sw6ptKJbgHzJgFaS
y2Q7rie8m2mvndLjj0Kk0k7TYFzhtD5q9FaBW72rd8TZnuLfhiLBshp49pJvKqWhOVrvzWBBgBv1
PeG5t6VqO9sNblEbZBNLvxyppxLROJeOwstP023Pch4R9UXg0IW+yZIaXc0YABx8BimvED6jHEIR
LxGujg48+yVMQ0p2nFMXn2aONmw6XrsJ/eHfiht08HtBTKkgbR2YEv1sheadPmAbzjnOUyfsdFxM
twx8hKSp8aLTKIIWOKTOZeYPEN9n2agNbfmbp8CdDo7lnOtLBsQeEeVx+j5InWtPeJs7XLWQCsug
eFp4amECMt5prUyv9RAMdAAb/bTn6iZWXsgLGvV4URknAW8kHh++aLVc+9BipUyimU4ssE4whrHh
wisALR/luUsjoMGOQ6hHkWt3HAFhD8ipQ0INlDTtjBcfDgdUeKqAKiR2aAej1Gh0Mu1q/oBPxQkg
gimlLi0gfElKOECvVFai4PZobzGuXTVrIWpcIzlnlcKEmR6EMCcYPDhpxGvMosjewUwAHqzi/jdo
9ZiWe2D+7r9nbj1wzOJDJdx0frffXyT3Wq4YYrSrgjBXS6Avzj9n22jvDaSg+WnNJdWxdNTThrGn
Vz2DHhF2dqrF8qK/9LleeO6i9ePbryaNpPdtzfuqjhgB2U523nRHJU9he4WAPC/347rPj5q4ZQ2v
xj4rNxDhh/1bEgdrYVUYuglKGdrmzUxdkxpiaxuSv7kTKyB5axzJIFfnMaa6mJVrJkLrN+QsUymS
Vuz7TsbCy+NT24BoFI203jko58XP7QCULApdqRejgNfiqMl8Cq5GlYT0LuC+P2x3tdbyz4lPIBr9
OknfXdZNCSep/XopBnqsNWNzY3DSlEpgao/CmtjPK8AYQmfiGMd9w90L7U9K+Z6NpJ+cWm+tw73f
+jYG0vS0kD8gMeTlh9twfztzYLIGpI7nZzd5U2udYCqapMWy587q0hzbZdA9gRcf8YcMUOFu29t6
kMRE4LySCTldRWB91I69czJvt1PIyj6Ju68jzOoM1Q5ir6wFw1ErwP9HH17fMv2LGYqq5z9lM8JV
dY85AUNbIYvPuKN5wlVQd7HLQq3b5oZhccfh3EJL50+i51SPL5Zaf48ruaqgx9ZPHHHLmKwRT5Jy
p6qd3V8s/rhqns8Jw7ps6meOc/oNQU8fg8YxZQrP7eLsFsO7CVA6w8EJ8sGMpkQxaVt4v/MuMmYh
680Ng0y+Kex1jnqULVQwgJXJETBT4SKvAxSy3K2Sk5+eNiqdtf43JPJYy9HiB6bz9zaI1a+3twxW
Hi/snAZrBxkLxlApecVE3cgBP6/BEESYc8UJUaSeiuOJPVvaeNfYJ81wD3MhTkS8AZVL65VoSjAH
F9Dpn7A0iBH3UxTcZcJf6lAzd2tfAo6DMhSienW19eCbLvZ65y6hgbLbaULl4Ct6Bm24JtwaZG43
6DHKtdJdFTqjUFT8Py4dNo2tZzY7O7oZe43FMSl+HVqvFEJBXvqxelpi5Ix/css6Y9qA7NAYLQ68
2Gu/BAc4gEL8+iayuyWXtrmSQrSRWLwv3Nqd428LzrAhMHvTOZFfbeMNwYwuR3r138oYpNHUMlaO
I/cIkrwfgd6t0agdQegTuSQ4lF31nyjmg48u+96mP3RKpTt45tl3cJxUO6W5vh01SdeBtHnCUl80
GceOui1ZS+WsvIXBr1MV77w5Y+/JVzBv/UJuact1J1lbOAbJBoFAeHli3RViDwHgdcBTX6DmniRg
888rmIuVDFVCjfwTO6Mv5Sjo7uYYJhSzhGEwAj5LXRHM28VI9Q7lkVB+SUwrZw5IMQJ7W47Ox194
oJHYHbF4DLQ4q+bMWOM5eFcoiTv6j+F6PkhtzZLXlQut8sZ7pz/m0zY96t1FLL4p3AB8SFPQIfBq
CwT2pRlhPm7hB1S/zGD+y9dXUN3Bj+CqNkmuNkrUBaiLjR9SZZDL6mZ6WiMxj6LMRQRwIKMBSMuY
0wXVEk3wBt2t0At+eC4wq0h28+r37MQZlRj2PjXNSZgnN1qY2/e+yfGuhf/GI4x3rlyAf8G3nybu
VYA9UkYYg0kLEQh29xeOzfy+OFS3mlVknEyMjk7Ble/TW7GOV3m0QtooXNGb3YPGf0ahmraZ8Lf2
F2DhSY933OoSJVKCntlG0lx7boq5fclsc3BaV/05U3eBHVWetIynbRXzrtD2j5MxKNoo44JdgBoR
ER0iRmjyBiqDQELuTo2dOv3/dppHxNDsbrOQqfhTB2FwcfX6TS1wYoaQbI6cRM/37nq6TKLdTvAf
LirzY6vhAz8ArsVceCuV5OftjybOKef+IFxUIN8CQzBxT7IDT8DD/dDUqqUDpTH1lA8GrET+8Aa2
3Xqzhj0QmC9J4BZy8rs8KHWoBlVn+AVA+xO1C9/Bv9nM+qdEkmy2xQFeJ2u2fNvMHQeeaFs9S1G4
JlLwV87lQ73Zi+Uhyf59qJdI2uD/EQr4iupEA6s7GOwHAfLJ+/AKOgND5aGFDwhC+lgHNHdFYOPI
JKBZa7YLvfP1vlcvUKRPfQpcq/Kys3Ivv3T8cSM2ECSYZH9R3vp4trdZLTJ9NHoGl2jc86MPOWUL
UmpS9xxE/Bj8REm912QAzdimLUZpWYvo/x/cyZzWMz9cpIvOmuWCxDfQ8MRLiH7p1QDZ+fp2JsJo
P0TgTPNzWPiBJCeF3pC33+pBvZLUOqAFlrfcxRS8/a3fRyERncrBD0Oytn4teLywv6rFFVCZOIrC
9LuD38qe8bAr5LPTRAm14nv/OweVfhsJq0l3YLIBGKxJ6hoITrvyjfngUMlFGUbdeRew/LPDyyns
/h2/c33GKtD6y1oqOrKTE2GXpNkjhz789f9PFaNu5eFWCSJedwH2JgIyDgftrw==
`protect end_protected
