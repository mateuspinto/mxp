��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���Z]�� �+��+6�8�)�2�<��?:���#�obxt$]A�_��2L�i�)�L�a�/� -V��i�
_k]"�odB�64�<� ��70ɋ� �Œь��gW�x@B�߳��X�-(��;��!'u��/�����<�D�c\>�-"��~�B���A1�|++]{iN�W�kI쥴��z���s7&��,�������iP.�wF@�9���]iM&Tꋽ���1^���Is�@h8�:HI�Ax105�� ���Œ�]K���=��:(��Α������5bӯ%:xN@X�G`�=7B~WA��K6�� �Vr~r�c�[�W���9h�BSR��x,\ /���\��r��X��������t���Dw��aؐ*�L�i�C��(
7Ċ�AE,&{/�q选"��q��2�wr���e%��全v��	m��)�x�x=�/E�$,fqˋ�k������ɠ�&Q��XJy���P_=8���a�6J��B��w�y�P	�L�F�^x���_�@���f�2{9���U)�(�7���V#>�����I�����ξE���?[�Գ�^~�͵g�O\	'�AL����	�s{:��Ѻ���C��о��@GƤ�nP�jd>�~��'\ E�u�ڎ�8�ֹ��μ���\c��dO�4���}�Ƨ�.�`�Й �Qn�1%1�恆jA�]J(��H��ؖ��H���?�A{��;�@B����p��(RK��ک�S����CV����Kt��U������N���=|\��:=tμh�M�8��|d�ZbP*���=�F��(M��-c4B#Z9�}�����ɷs�C(P�;0�֌uOݵ��޻A0���I��泋aFGβ��.a_F�Y%l���.>1`��J�t8n%�;���v���O��](���l �=�-1���௘�0qG���.�aL�/�������s��&?L�Ѝꯨ���?��8�Z��0	���h��*c�V��l�|�T2F>�0��Z���p�/7=��9��9�Q�B����c.[	�fR�Fb���!.B�\��� ���'���^�"��PBlz���4�,\?D���#1�XNl�@�L"m<���cG!�i��{qZ�B$|�	��9��j���ʨ�X�@gr�E���ȕk��eC����׶��|	.gX\����wZr^Y_S��UPz�%M��w��k_������8�m�(�"��y�Ϯ�d�$[q3�8iJ���V7�\ {#��jr����҉e�#�wX���yB��g���_���>W%���)��������#39?�A�/��7�o������FnA��H�"����vM��.�/�%5K ׁno�$�n������oG/�,�On�BW������~�c��3&�~��D��\�!�_�i\0կ��򱾶��G�t���"���˔���O��}�S�l��z%)5�C�xa�١T��.��n �h��ڍ;hn���C���"k�\��[3c�L�-U��ϵ���!9WƱFb�m,p� *���G�t��[�<�	���1�_JN��$"�{���?A�M�:���:Q��@O9�pA/Pad&a�jW��pH�`fǁ�BmfŪ��$����=,]$�ǒ:�|��!tYH*�EG*�zN�^��.�����޶D^�'T���i��W�tbZs�o���)Cf�6k��x`����V�l��[��ϧ�ߎ�@0aH�b��h����,!�������LR&}�59�+ʣ�Pb���5s4�9���%G%��o��Eh�j�D_�|8���{����泸�~<&��������O�gZs�������ey�Ì:���
!��V��e�%� �e=�!�1b>�5�L�.��<e4���-ps��YQ�$|Iڬ��e��`�%:Gf�cC*� ���hi;������A�G\��9��֙�L|=��prZ`��͡��9����A�Y/��x� ���f*��'�~�f����a��� ��ٔ"ֈ��}3�gS��5�|!q�~>FF��F�ለ�J�6B+�!�,��3&E�k�s��53(��y�a&Z�ʫ(�t�>ݑ�.g��='������:?�)�=�ǈ�4���G#�XS�&���ޅ�/5!�V\t�W�R:jt�(�5ė�����	F��ϛ��U��-���@�A�����䯺��,��f���6�Â��Z�R�5ٱ�W�#��A����B���~l�P9a��cP���>�s^Q0�E��f!�m��+�lcnm7%R���_���em�A&۪�k=n+�����m.�����N��r̦��4��0�0��� 9�P'-�m�m9�w��|6H���[J�㎹A�O��vOG�'�r��ߩ$�Մ'�����^�:�����~���ֶ�.�Z��Կ8D���	ROq�\B�Q�s�V��u�l�P~�;���}���(��-"��"��Ydy&��S60�����P���X'g��3��v��m�����PWn������,�p�4gU3f�����WF��/CD;�;�ͭ��Y�����x*z%�VΕ�q�d�6�3��8{�J�p:X��_�yC�D����-5fl�GE�60,���%���$zT�����I�|D�.�<�1��P�ua����Q�Z���T���D����+�)�\�}:�nW9P����i��Zg����Y�L~?U쇈�(��ˢ�/?�؄߄Yi����ޱQ������(5�Q�����yG�6����z,�I^��Ԫ���Κ��J|�-a��/GO�{ѭ?�k;h�_��Yy��o{"��7J�k�<�z�k���DRjW��.a�WɧH��`�9��9.�5)���K0�V]�[��b� K<8��"L-����zIഛwz}B���ަLޮG0�Y�M��n���'S9�����#/j�B���I��Qt��b�>ת�~`v���*��/��v���cB�a�mƩ}/ܷW���'�%?�Mv�C��!N��Z�O���ak*�aTc�� ���+B�.�*�h�<℆����i����,p�<UD���~�n�-m����A��Z��MO��=�H	��Ѳ���ƫ�Ҭ��n!CIAȑ��ǯ�4�c�R���g�%d�H�0b��T%��sAh�i0�
�$���}~_2N�#�a@K�9���=�	�:�!��O�L0Zt�9򐨼Ǭ{B�曉Jq����ks�m�h�!���ӽLf�l���>z��n*��_	!NO�75J?���o�r��|�)8"�2LR�]P!}B���`�����%��Ų�~�2�y�J�p2{���$�0&��?��A!�����Ԍ��6mB�RAˤ��O��	J���T�x�,ڑ5�ҍ��.�%	�-�7�6�ne�l]O���ݗ��� ��s�����aػ�֫LQs������s��W�[Z�+�~���c�=�L.��y��]��,(;,&Hi5D�6<a9�RX�\�NZnL^��i�Me3�۱�C�DG-���죫9�xǋ��|� @�0Ƀ+�ʱ�����A��Z��
gm�]�e0��&�L���n�qP&�vΞ{�X����iGm�,'�b�� ��i�]N����Ԗ�L뗝�YҴ����A�i�y���9[�^}��c��k�4��r >�����_}LE�gt;'�H����q�|�>�������B�>�3�Fz��S�>?��JO�t�솞{��B�'��+^ʻI��N�q\���
Oe�M�C[�g�4"5�%_!�4����1м:� �����2)��P.�8 x������/�G�?�c�0��15$�{��)T̅$��3�_��?4=1("�G%���	3����x&R��$}z?��聚%4I���h��2#5���F���#y��w���an�r�-rLFj�"��i����i��H���A��dxD�����ffv�jj�����������;�,�"�7N[�ͪw^_c�|l���F���AHʚq�}%;s�q0�1�S��F!���'�����������[,m���-ٟq�����->���a��h2츜l��&�l".X�b
Y^���j��}	MHS�̑����0��5����1߿L�9范.V�~��k.ۂ��Kd �V[���N�%t�J�2m���z�ѐU�d�gv 6�縴�7�Fqg�sl�x�� �),��4��RF��\E`�x;�	W��@��r�H	jąkY����wy���1fk#׳�`j�y���t�pQ�ܻ{�P"�2B�z���t�ΩLh<l ��:��^�8ͬy|����g��h|�0��@H>,�밊�8��J��~�@�G����r#���O�phO�S�_�T��j[~5'_�t���\���m�[qo���e��&Vg?�+������+ҘM&�b&���b~"��{}�w�]�ҟ�SF�E��mğ�d3 �N5�kN�k:�0h�Z�z��2X�{ġ�+�L�+�-����h�ʏ�Ц�a�g�B���?eb+��K���g]����c��
Z�{Z�����;����Ot7�]����!ڶ, +-��p���{j�v�mW#:<}3�
/�"�B��}�!��B��BZ��}7�O��\�n�Q�O2��|>$��x?�b���?��@=�i�!�""?i@E��'A~�:�h�
-29{:�O㼼ߜ�E~m���!�O�p��YDv*���&[E\���B�UG�B&x�]u�����ل^\�7e�\� ���w�C�3��7�("ٟ��+z�Z�ZW������_�X%���b��u2zW�g��nq]��6�%�����긑�gBΰ��o��7+�O�@����Q�Z!���x.�3$�a��t�\��[�ɵ3់)��p�b�2��{k�JbL_#��I���hO�SMh;�G�/���6ij�S)ŕI92
-	W�PS���;�d��{n�;
f��?��)�o6I=������W���(�z����׋��Jǟ��v=<��G��^��H��K۩I�Q���	���6B��J���'������A��.��xx9@��9�u|�P�}�V5���嘐�Ϊ��F,`95H0�>�I�XZ��>
�ߦ��Q���"�3�;�^�Iz
����}�H)�{g��b����x�&�݆W������sZ�f'�]��8�6���ʬ�qt���ֈIQ�&ZѺ�ɇkM�]H�y��<�X[#&ϊ�t�峴���ū)�\������ךrk���_:X�QC&ߠ��ˉbІi_v{]y`e�!��L8�?�`��I�(�y�����X�	HZ� m���d	5*g[	F�����}����2Z#�=�]!G"��Җ���Dg�sa�Lgdm4��4�9LPT���0�!�"�oܝ����������ob]����D�2����ʕ�c�f� ����:!�M�Yr�y���{@�Q�//L:��߃���rB9
d�i��ݖ�&i7��ﱳ�Y3�7a^O��3M�����;A���s�w�滛��|��-�U���9Y@5��].W���Ʋ(����oo8��aby���(,��T"�{a�\==�L#aQ��v��(�J�&��Č��k&E�n��UM�~;Eb�\r�'=ena���K��X��WK4 ��N��|Y�u"�&�7�9gE��8lQf�1oW����m��u>�J�-4N ��wJ��x��u��MV	�=��dU$��<+�J����+�N���_���%ֻp�>�I��Ǭ�7�{���t9�y��ՂN75���rΎ(�,1�j������Y�ApP`�/c��X}�v��.�Rr������K��ΞK�����TzN�R�1��Z�t����ӕ������7���/�y���^�"��*8H
�x�"�����py����:�Z���4)Eo�K.�	#V2T-���h��"�E��X�(��䆅�~���i���>8�F�f7�ɨ��I�n��� ,���� XH��Y������8H9�K����S��yk���W�U������I�� u,��I����k�6��1�SC���e@�q�|&m��d=��)�[�O�w�n�����������9��	��Vc6L�����Rq�*�ɗ�P+}%������ B����|
���m������f q�k�X�a��:�As���@;��1�'=��X��g$E{���HN��� g�`��-zV>�&��2��Z�`�b�X>��d��n9J�5��]�d�ùI
�Z�')I�y��Ѷ���1�+\2�>i�4�ç)ۦ���1$�Fws�ލ�#��Q���ŕ��O%CW�?�y���pU-J7l���@�J�l�p�E2�a.Q.����6j��	��R����؛�J���_��Q�2C
�D\�};
�����7_�D:/E]Ey�J+��r��\������y[��3o�[�y�Xu������m8�����@6�z�j.bZB��&.����������z/�f$l�#�������C�~4\m��@�Օ�F2�&����' ϗ�������F.��