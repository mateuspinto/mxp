`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
DsT343niLHjvFObRVbCpXbmOTwmvZMDKhriczqQ5lG4TxiDhdCy/ivb0zyUfoliGJqajDKvfUUQi
LAM+xMT0OKzLMu+Ms+I/zS9ocEc6kR8GyBtxD/mEyEYmXB8WSS8KlWVImTWEWP4mwTXd8zeIcrSO
GNIhWQBibc5uaGV9IQG3nuw/V7zTqbKpAJCrOxcS3LKsIcbuuECO45muwpYNEWkABh4JoVpEVa6x
16DUar9ok1e/gW8+Pz0maYc2MmCYTpdHOBCRotzS4GOPQeDjSTr/stcseBHNasGxCtSEratCh8Tf
3Jy6xPOZ74juPEyX3DaFFJ1Gm/dcMsWNMVeRXA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="gq3UQL1UbY5uWO/OTlbkn9jsVcskkFRWqVmO3PIYELQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 48352)
`protect data_block
8fLYsQfX5jY9aAFUSzfp0TcVAU+ryvMx3Plg22A1chnupaKI4ckQkqrFgdCB50SvSOd0YHGZ0rFu
C59bSL4uAmkp3SgzhgIJNElpMjLXNoEvA3/x8unU2Ft+SiXECYio16o8LNNk5hCghxKL7SHDdeff
NvplLtYIz5bfTJjmkpea/ay/ca4YrHh4BplXgiIEanWG5LInavLTasSYqqBIleP8d9L/JAuWOawe
SQDG+wV4bVFivg484WnSPZ3Y7SwH71Y+F/HqSEwDaL9oEWaNIR+DGJqE9/LYESd0Zok8L7n7Yk0S
taMvaOk9ZRX7SviWgfjAyDuW0YL43k9JS3PyijsX/MeDczCCIm1z12hNOO+CW4WNUo6tai2aVUw1
q7KI15R96g2qJOOcQxqxNtXxPkVxTjIH2WPQClrTAaOmmqAYS+DagK/ytWK9uwOp4E7Zx+M/S+Yb
MTgAtDDIAAlv7ovT7Xy+NXl+b3j6kWbolONRVnGJNLNZ8V/Esj03n9ueizPYfory4Pmh2CYFLaqE
urxkzcU+sml4OXRyT6P/++gJr6yBLMLLw21rryMPaVGZNq1zMmGVG2b6Wn8sczm4xkjyzOMCYMlj
jVafnPtFKhBEqwY0RHjc2eDaOg31HvtYF1uXiWowmhTSZKW6mCJ+XJuhnkck27mRKlRSGaxf0mUz
ysGNhGXd+fALwGlgA3kxsx8Go4gOhkn2tZDqTQwuCRt/ahQxAi7fVqIva02VIDCZlrRm5EFSgjB9
4KsiPRcMLC5Ci1WCPaJ1KVkakfHLwiw76vDmqgSnbp0s/dZ+ZqW0jGYZiyZXb0BTV7Nfz4PD+M6Y
SXelGrpw48ehphn/Y2BetcBTFAR3HOGGj1NmJIVRMxgql1f6l39ry8Fye+sBhJgaLcKC9NcDScA8
3K5i9CFVlpR73y7XcZocv+bJ/G1FtLnzwJSsiQ+UJtZI5IenV6kW69Z3QxYnAHu9+/mAailDtGTP
f74PfCAy5OKAGp9CXzUKz0tdFcvAH3MATZNmxqe8F0BByGG2ApCmcLA74UMEW5C5XbRdaIPnNdAF
NQWA033vEI5C1A9UdA+gAz9td2WM+unFJVinS4YUP2GsplnghXlXIJmOPSPnhE21pDMt7BuQQX/d
6DIA0etYWoIsqKbDfE6NgccHypXuSjrOrHv3iv2GEvh5ISAFUS4K40CHZRr9OZaxD+zOr9ae9tLE
2ZHBOQOKgk7NrHyNqBzXOxsdoKwwAafldaAtsJVQ0duslZliAPJjQqDZBNd5v80pB1uMn44XcyHK
IITV6hviY66jZvDMEsnSjh5xxn/yGSkfn7Ku4CIbpGn4kjwQTipMrSkRzfQrgFTgjkg3uFbJUWEk
G/MaxUl8fj/OIFJCiQ/HkhaEZrv/pry77gI5f/ZbiduW9jt0QXY78xsbTfisNZl8L/iFW7jnvzu7
0uUpTJJS4SFfmhvVxpNHHdqgnmJY1ZodIM04zC7SV1B7R6NQBj9t/66HrmMLrwX1hm1NNBZi1peT
gsQfbXpXSRRo1qBMi+CVLjFCaq+AbGwm1VN1I3xUlAZnspwnRnI8gSFFyofav/89Hmt6MUI+wy4a
DBvuDVTTYO/G/Yn+XcpuB+VP4sWeQmHirAv3rpyE3vB13hEinkEvcbgQM7pepdK67U4WEgHnAxtQ
nq9CJkpByX19m40LQ1tdKRa5TWwBgnX+xOad3IXx7PW3VDLSgc+k0WQyZWz2xkWjEAZ6Qcz34Uzz
8seuPUGgi/S4WNWD5rei5KOefmU+SEUHV+9KBakacg4CiYwUprTT7Eom/S+QrZ2KmEL+XovFqODp
wHo/L43CbyegOkXtrU1HyXFj0YxDGL4fxjrFs10pW9TWjnPbqJzKLL8H6Pi6i8nJ6S6/fbRTAEPt
cshcfmOwTYyuuN1yNGW2DtJwkIYSe0t6BsktMxhzsM1BttgK6ld10i75GNW7ek+VXTMhasUZhpT3
0vdPHPVS/NkmOcUdNSA2eDc4w3NdgFuxiURBhqF9SYzLVnIDYGIuP3cxdqk9tm6UwUoVheea/Onp
QcDKANX7ZXlIu1jhIGcnELcvEN9u95EwPjTabZYtZrGyVjXdd3dfXfWL2KOy1th3p76JLgju5kkx
HTmGc8LhYN6aqTgV2K2ue2h3gl9cI4To0Mfek25o/OYuOc5TZK81eyJggUaG0i3GZffM9LN2wGJs
28N5zlxagx21CzCfrwbih7hiCFWkXtCE+L2xXX/rrCE2U4gjUFYrOVcWXRN2OCiwLrB4pGy4Sln+
JdimmJYOpty4jsP2erC0O7LvXUD5P4wEi7MoaDcljBqUyteGmaGh7hMiAgn4ZJSiFShcnPQnZS+7
ZLgUsMjVz5tAEcrSYFl8U/sbrJS/asGYKp9dt3X9D7dC1OfAKpod3r+uHUJQmdMUh0lQYztse7PD
YinCj39c4rLMefpr0dokuI6N20N65VE9eMfeZfGi8KdEITxwsQoB4xb1uCoD/Fi/v0hnvlM8t3LH
aPofB5xj4PVxF23GqgaxAFt7a/THQJBN5AApJnJki/MfnzvPMAOUpEiBQDB8aHfC3wLpLUZRyLtk
RVXkgMTWgfJA0+ZdbamTHHgD2F616xcBzQIn9aSyNT3LUpPv+ogxyh8xjCAD89tXAEzx23E7mLmy
xHSc5qT4afvAyQazx9Ntodo1X4ZHee9pprBoTr/tYBd3ZeuDskOyO0S8Mv73NNZd4Rr0GLEkjvVt
zZKsqW8WP3bRX+2VpAxXWacO/RjXBE/F0BnpDKAhmiiLXn+fluy1GIdVZyUzINo5KOA13GSzPlZB
64uYoUG7V0o3SeO1NhCfeFOv8yAilfvJyOrXoIHxqpjxSnjttssKATMy4Iau4nFSZj4FkIqvY1s6
DXaCPQo7OxAA9cFAesxn912G1zo8ZqhtK5BB69EBlhVfsPszJ0mRSQ1Tn+CaCwPxpF4kBzCKP5w5
Wef5gQzdjvfBD3t96RYNZ512ifhUTsmaQK2EGlEPGSiTrSxEjK37qsTxcRgnpjXcuCsE04SNtlGb
laaiwquPwh8Y1rH8OdoKF/e1Lg+We8p3NnqAGouAnKtFlD4lz6X2sP4HMMEDBd+wR6TmjM/PZMfv
2hFNBjJSBPO7lN9VBLwm3yKbrfbUzNkgsUTtJPdyjnAEvL+oBDmFPw6hGZu1RSvO+bCvu8pseLDj
7VU4O/TG/PhoJbEhXbRHtdD9CH9bPXCzyp+3BxlEFajn/tJgSh2J9EHiHUqzHx8Bf8hAQqRDK+Ra
JK/y/nKptss6qC0KvZv91nS3GHvY6S2SK1Z4Mn1CuYU0ThlldOk2PsgtDW1+qxc25MsecLTaTJRt
QqaQSH4BUy6WJ/7TOjNwsk997fprPXx3xn4YAaaF3koP7lMeK2Ho0BPZfYEMZqCWUa95qxULXOUx
gH3cjp2oqanRgsPblH61Y71iaZvK8JvyiGhBwmTND+tyee+ziZ+ka+td6g+ncLNnMhMoU4VtZ4fu
1Kkl1+bBhQSpPUIdj7pOxaUVIj/KpNqKCakfSkH0ncahuz+g8Vx+Of8N7Y3UoNz0NxIZagMaw3WO
+xKv4y6wLose1jiTbpFMlRsV4W1/MoDZJuglbg2pLVV0MQWbI4Ao7uTMgnpzdMhAIrmr3HrKhjhw
5Kf/wvPJSG6VFXIQD2HTGa4ZFGU6V8Vbeh0fu+Qeifys90axyEjx8NNO/WM7KdY5Bm3oPArNm+wG
XkyPp2lYZVYSePuST9mr9gkIVG1dEzbjsEl2yAz7LZmi1Rm1+miC1FX0OLgELZph7j4Yr3cXc31c
o8g0Keoe4ixUbLOV961TyeM23TA9MtFXRQJqJkIHUH3IOEefrS9KEQzgaOjtzsyVyjOHfjUsmdAn
K6PLECOAtezFvCLUF6j0Gttu/gj6ssHAx9pwAnxy8rfQ/wAoV9fTLyJbaqYzh8GYr4cRrOzwlDLZ
o7FoAEFDDqMV9YQhIuIGrilZYuDXkY/m+9dPlbRMrFnHJOVBVvU36R4M0ECBbcg0l1XNrkuX7jf6
pd1Kq8orZDrU0b6YTyww3i9okyYz6DHOY/sDihcJXJprW81gXMjKobvHlsoyXuJw2EThc9yGImwA
Av6T6G+DFrLNHmZAPD8GQ5SyCHXwKmYXDa15k8Fo6VtbBtgmVACZFSY9w82boHcqfLbH+URw++5o
45B0ievGarMsbPTtGb/TMzr9pnn1Yt6b2hj/5CrDnexW/mv5CpA4sh8aKKYgZmReP3pvdTEogOv4
nGzpgfU4UdP87XLNWitzpc00yeTAq9sMtzf4tvlOH4GpVTLAfL2k9AqDkqDZTvXg8thORuYPdPzC
ebrUSYLVRhyp3EuKx2gGPmpmnORhmutNXG22bT69vK36EY+n/XStQdb1DY1RuyZ02TLKWRCCRLaN
5YBKQhEwKcL3hUz093copY4yhnkmJYQUV77HLi1ow4HQxz1ueOhUPMhA6OChVuYYY8rItyHcyXVt
G16jfpgt5VMabX1GfIueSwZsG2Sysm/lbvkhhic6B7B1Ld6cqg+khWq5pB2Z0hfyWB3BSMqKQX58
ENDW6DVXb8mQAQiysYHbXNeGlu/BLiw4P7NqVnXSf566xtRaYmEZ+fVe5ivrhJWwd3Bqo/tDjrkV
TSC7U0Pc9h271x+JTQlw9xFquuQS51oyHfqpx5r0No8FFfpcmaSDVM67QplrN8Q+SmMdhGjHiCY7
lBJEzPw29KclO0jd0nzlvCUO0S/9MXLkRHXiNInmIMqKKnAL6swlgcm95wb9kHCWCrz+VLz6XScW
ps3ns+zC94GN8KuBZQRvmS58ALFzejrGWaIP/neXWHkyePJm6YnzakJcDkl7yJLnSE20PuGl0k0Z
LQcG3brrUU/pj3kOG+gP6amvlMOrEnMXnn4oMLy0pyS5vIG+RO8jEPqIKinh2P5DR4XcQaF1NMgV
DVWWyyB+No3z7/VkZZ2dZFg9BS/WiRo9akXUdwohTWlgBfTvqayybC4mJKFLHo9S4y9A88eS7Nph
kumB46lt8TfnqWPXgCljcDbvG96CWWj/TJJrqOnFe3wQjH2FGJzXHDIROhQVjgvYFJ+6Z+n9lp2s
8ZlMInGV6lUDatZS4rGFd8q9M5tvWJ848AsF5ur0ahO1Xo+xipsJYV15x7UZNH+cYMlqpen9rtaU
+ltcLCftLvVEDljTaXOr/98uzvz3/dP/Sn+DoB06i/mYuPLzpQWm7AdJRTsK7Pc7tYf2TmbmqxfK
u/krbzCTK+ddMu58IYzeZqASPU4Qk5wTd5Mod14LxDRNFzq8dILu2oSmswDlIcYKLVGqsOJJIkug
fY8+6Wf4TjZOvg3u8F9Ga9b1pcBKIyE/dkra+qFg7rzzbg8J8PJkaorHZ/G5hKZeDqhlLCTIxhcJ
F/qpht1z3aN9ai+u2k7RUruYwlWL1uRP3fhYAniYbz0AqJDcoFC7K3oaW2qBkrXXiwN5ZJKT0s8W
o0Vni717m5Tffw/9+guhYg8Q1aA7minRcjr+DbdLHVWv9fU2s91lk3WpcZszmgYHG/OW2gMQl3iE
hG/mgi1+MmEgX1515cppWAT89VoqbubG0Y5HgI60ODZb7ARM2jk1wYz5EEcrUUQI0AqOHtlqBorx
QGQZPBTRtTlMKun1XaTXTlHIgxJkJKeWRgf/nmes0UC57iECJRQax8tTb4hLU89ri+T1XNKI5cuj
VEKqvbjutZHK5/uw6X9GgJtQMvnX2e9HfyloTVChUFgy2ExDyaYVlYUxZmsI0H2q6q698Uv4YMvf
Ktusr5ozB0QNLCDqdrEjbwta8EhYlP/0aDwD6e/kZ99kX0i8yiHrNQijDLcX6Fbj0X7tfaPyH6hL
ALt8Da1cEHGmLMy+AuvOIqVoXQfBydsiiZxvKkgUSxShTw3IvDfm/XtcGumye9bijdTovUpX5UCR
mtxdcWEgUx+tromZObsGeLfD1dTsi8N5BmXbYlee+VobCNeEpaK30cHX7RAkDDMNT2oar2uF0PlE
qxNriURANQ0E033KaOQIqvkNqGFeq7UQkGH2OYlp4cFGtMrFhAzHlnQrIhseiCinmiXdYTj0ioAE
vSvhbiRMARiUw5up5U5ljWBRXPVLQXZnxhgesA3UGEDYYD72f/04oPp7p6342RkvrU6umMSsEeaF
5YQpEskkMD7RPtlQzBtK6jqaCenNWxn8qCggYRE+5aqCITMNf2ulX0QmzWA7/9yRFU2pkL98nPyv
i16nUHNmDX8+o588kXrfvIKvdp0ISE5p8ODn/UqbvwFCEAcFQGBAXCy7FM9Wi+Y9f9SkE7Rn0tNn
jGvcAQ98jPx7VvWTHyBWqLkZglGoCIIo4E/tk6TaF+2DGFpOMg/h4El2Q6ZIwJ56xNmfKkPYCZLO
eTXx2Y2WxFuk+ZlpRJX73ipJgmqsi2WrSu6RNAavdZ8tHMpSVif0FQZSCOqEV1dchO3VkzSPgJKz
AStxD8GoHA3n+bn1ucsE4rB7QROo8qsxNvcPx2ogQqaQcQ1L/TANWUOvmYWgjxyQIXjUgDf4V0NT
7cHhA/jgrNCYBkVwg9nvKp4GglQ2YxaLrrtUjwvhh+u+h236G05x+B1jUH7iEv29Bjg5gKNBLaWu
Ut0YMMu3DcDx3g4uNojPrdr15Mv/HvWh/nj7TyzmrmE1tZ1q2fGIMwyk/HqohOBkzHCvEKJfqUBl
PJBWxOmmd9pttKTHwqeTBoXoO7RBqYKtQEcjR38zMgnryrzEPwrE9yVnjTkfFUpYFnSphyds1J3e
WsOhrRA0WrOnR7knoG8o/PqRy5bHm60Ni7oH7p/e1LcebtYgco3twyVy95T1WqEP89Zfpy2XtmDj
yHAPrOtyMspbcgNZ+oDUFN6LuoTBKrHN758mPhPZ0arcY4BShmKbN1ubuk2/gHM7jgmClslrGBMx
77v2UZFYfbOZOmbpQoiHebzJLdwHbdOAlErGV4mcQF6zoqI5udJ5TbRb3iwZ7K0MxLobN2w6NqGk
gmz5VNdPGpF1vh2xa+cNgXJ2zk9ivIEldD6YUu7mGFxNADVNr4X4bEL7EXwp6xUSmtC76i735loL
1pLQd2iXJG+9MYTn6TcGvwyA3dXa7ckuOMHFnS7HB4DfC7osC4qwrSSlxxuJzaI61rNJSVRm1gLm
Yu7sVNWufsqZuYBbCpX3/suMgYHB2qZRTD7fTpsDlBoSdVI5zs8DUQorQ5Qe/eS1JvQMWxLLvesg
2bZJxr/YGrxL2U7t7rdWR47ZsMbxgqHMe9OUHqWvyZjy2GDRcIFqLXx+hbbQEIyfBCugiVpALbIk
sp+h0KAer4TlkTxq2DpWjkqofCYkX+qRZmvqfuRX5UECK3EV1DwDv7ukcJDOdHePe7PQgR6wAAMH
UfOyooDC6mcdPfS41v+xAWTf5KMT0rGjQ8xkaCqlKxbQqnHe9Qb8TmOrwgmA2MFNPOheZq6E06oo
Z1FD2VL0NN9Mr1bhU9uaRu6gaoYrRIEMzsZVRHhZQpkvlb1nJVwQxG9R9lVPexvhdEiU2Gj4lj/b
MrdhPFIYAHWm20XgLtKB/oV2SYEROR5dIpAk6nusqbGNW7nw7h8rie4SHv/39o+EC3Hzde6l57Ki
b6GmlWxpUxBAjf0pWkRrTIAm2dzG8780+K2GKieU/u1CTQtXHRlOTEvByGJ1BOq05BqrHRi1v9g8
f2hFZOVFeJsw/OWKv+DgDd0ZPhs64hPZYPNzGKxQELcPTrZzu2e7Pal+fgBumB/k8fhFACpT4KIT
F6AB/xwJOKz79zEm2ag3zyOYa2u139RWVNvan009UtRFOeAfv/ktVih/cASRjFgV8zs3TZuZJgtv
Ul9x3TANPR6YZ+gjCzekUhNHbHhPL5wbiq/Pq6GwRrAiXPFQTyToDShiGSJdcX0vqbT6+ONDyfG8
JGA1ytUV/TvKhjFdgsrTSxB5n3n5TDRkdw+M2LvU6/S1LF6/M5IlEDPtWaip3FhUB3Ea6wNMf3RO
w2TqDn0DVxLUIIQ3ZMqzWigckZ2FlAScQn8VXpvS4xHD30Eo0km0TFezBgjqwqDMW4ZdCgh/5ysl
xbMABEpL8nYVtB8wPawnlAAl1ZBZFXBfT8zh/DWzUHJppy2aINbaUGKQNf7I1ar/vBnLsWHytpKM
afzTOww9hS/6lFNRSn33oMUvpCBck6++1RdB7I7wv/oRRUlgd5BHSf+qeXJ9XC+WMRzcS4TABsmi
Gigp4A5988gnDUaFt988SIsCim9h1sILEzUIFGWrxx4UeekvzcX2i4vyAxRo5QdqzKKEvybIryce
y1GEqvb1U4xP3n+11pP6jKS340OA35TGbeg4UjVpPCRRstPhE0bb1bYWFdPNf5ZQ/OW7JnQHMxdg
dqAaavvWXVztQNLp/F+Zs7b6ofOWlM+V1W4lKROy6Ntv0qupuJ+ffcB4qnlJ7qJkLgLhCHgtkTL6
FG60DXHiPcTH2dPYJBC9paPuUhWfSHdgPZpENQy2f7oKkTlc79OyboHW6MjmkUBEemqmJmfr47JI
3CttBSinEXcjkUvhQuXHzVw1lFUnSQpMkRZ2YyKP1oC1Fv2N+x8muNNDiX7QkkTkRgZ6XbVxEnWx
v+Faj5ylQAdmkxZixtlWJcXnQoKdM/FAUjWNm6CMf83jzG45zihIZABgonfQ+A+8T2tzNGAnmQ08
AkoQq5XMRbgVWRGK5hH2m2NWQ5vTmOq5gfJLHcXWXF8O8NDB/A3AU1WJVaYUDS/Qg04p896zbOgo
pl2t0pHYNQisxpRSJzKvKGzXJ11lHuv4G+xF++Ti8/Xb7uZ5DSCkJdAitpNWSfblqmDelMQBu9SX
kE+aOytZBMsaVS89OOlIT3l9CMgiZ+YJICXYYDHBvUL47P3iT9kEzY5xECNp+x+VlFVIB4LgCDlK
39rHASLKIc5r/Itlid6/PN2NwYm64eDzABlgYkpybtqOQTUUB/bLzejzpBwT4JPHCsL2YA3/vkrg
9HUPPr2bqcklQCqFooYogCXadHZ8dd1XuGS9rI83V/bqLGDOIsGd4amZD44KxNizdQ7FRyWGfMdT
ITg23Xe/Ouzd2vDGV7Sx2xaxpkB0JSrkLGFY3pVuCUw02GIm9htBkH404d8ZwlBaU9hZfpZNTGGp
SEgi3hm7fPTcq38LJroJXa94zU+CbVRFHUQMlUt6yg99KplLIkD7PPEfjBH/f0NsIc65VyvkDynB
pUVXxarN2DtCFtiUAO1cd7Wy167AABCxHjUd/4NAilm2uTderrb+VQz8rinz4EwnVp6Y3w1vfiM5
89FgrO6FCGw2Ez/SUBWVTrgnwx0oQdrYfoSc3lnuM/IDgpk0eRnc1/c8179DK6H56wKC5KzDlbN4
abB9f43clZQnQOTTH5LTYJyy9L49sQTroAlmb1I89bOSDkyyXytKdTcqU75+dZ3PSUqLYC+XI0nj
0ZEPwKn42ohGq5z3d2sGjhbOOovP+5IGWg5k862Yju5ojc+wiydpVTcgPjMe3Azr2okEmtBoA2+z
+0xpB3q7DrS3uGaztI+v6RIaVkp1znam0Spjv7jsEUhDimTcyUsXGJTobBI87U7bmWIGth/1KtTU
78I1L+9Pzmm7gVJlKTHwuTeIJ8SXnCzrbBTTeRfXsQ2wg3pQqkwtJL6zf1JeZDDhmdsvseqxebbD
Y/ktoc5uzhuxTT/suPRJPXJun/sSwu0V4i9FEMq9faVWWCqBrKr4Bdg2/XhS3V+ulC2gY/f9k95C
ukLMaLl7pIt7r0VBFsHxxhNwA6/jcwzEWSy53oBth6+7xwRGEcsQRExYjINFKFBh77vIgvg2yQjI
/AQTFuL5ykUhG89vLfvBgpLs9Q9T0NEpIoS1hElqZ126G8zfGilC67Tv+CvaGzF1dBuclrTTmPXc
SaAseTl9TrdmWfdWZWBZ15eY4xX9ej/W9xsZ9QOEWFZTuyq4Fpe2frwArXBGOKJPhGlwnkQzFmFK
EccLpAMCz8d4fwIWaImPNpIYUV7cJXCKwgKKo20FUA0vQX3cdJEkLuFhDNDh2LivzdruX0p6/Nxp
i8TKV3geym+3inOvZCKX7QI4X6Hfb/BirjzTykZQnOe/OveFeEYvB8Vv4HcJjolNFyEHDJsEO7CC
DIlEXekLzC5WrRXztktnjM6q+niLGzoAhTQsaTXv57IGqtX286sBimizs9lxQeY9D39e2H8JrXZH
/tEaeOjCzaz604Es4IfigirrejR69Phobb7HeRLFux8AYBJ5himQzXCYOrctkzEW1xmHHRVRx8sa
0yoPCauJLRNrpdwvCkX7AHSs7N+GzACIK3wDRjwkX300FDOyq6vah/qVgPzs4EAto7Lst0zh3GB7
OrdlQvS4cslyrDtlBzb8M1KzB+L9BwsRinEBqgaFWqcFbVz0WJhhDCG9iUvkWQKC/iOs4DOott60
FFPdVS2751d1hCCPeq3BX6tVJDGII31Pso/83Q0Tbh7QfHxhaNLfjkqZSOjAGQrxyGgia908w2+b
Dxt+WT1MBOzUzVmzhxQDGZXcrjQF5xoyB/1acJdmD2ayKsbLvlBuDPmWJpWi4oH3cAJnd/XmgOh9
SoAJ0CN9bMQzhIZF2uTKo/9xfQ6QfCwSOFoPsYRf+EvNO6YUz9TKwExNoL3Lgm3Ar1CKKlV2Fpd0
BG/Q3caFYKOO7tn6eWHDCGyuSQD2Lu0mdlgW4jbQ/TU2DCgzE6FWmeewuKXjWsUTlC5wFKtYGZOJ
pEkqwvPZBaI0NjThYKIzYWF0MtLANkYLM0SjBnjL3LX3XMEQM6o9Uaclq+0idYSDBfZ3NvF11sSq
Iiv2QCZ4oXfGzlG1H3aCcARcLX7pmRgYI0ImwqnoJkCK5GXMdFwoOfcxuZ+ynk2PGhb6/BYNywJ7
k9Z+2rVQdPgWpORgKhW1OOKzUMBl3tQ7QJnXAEPQuqouXUP4CApZRjAN3Fn4nx5mTxCQTlUNQLcU
gTlES2FnlAzgv+uelR99mIWU4E7DPJQnP5rSta5roK/pVDsN3q8Ctt4db+9Ymq4RnSQtqPw9hZGS
+X6UobA+ZIAUBAy01Xt16ut7J21C9Qm9OSfcwf0ItGV7oEMK2LypYC4IRKq1pf9iebppgwNbO1nf
Xo5qWhXJ+GC3rfGfoBeyHAnAyuUV/4dc6aGaFLnN3FsUzbIVu4e1wNPH1QJ5SnoFV29SmSWm0w3k
4bUEC2MCKJg7InyRKCUGvqmdfxh35dgcVd/wGDHTib28m51RFimlvfNbn6fkFcW8RhEFdO8RCvDS
HShsjhB6rhBqEFNqJH41t7Wl6J7HyL+o5ntmnLXyZsPuLwDS2LjqtUsAq6Pm2kQt5uUoIJT7eKzv
vTqh0Nn8ccruHnszaYZgOhkWqRgYVXpbvNPr1f0R0qxqjopFGW9oavw10J0lzjc/hDg/o0weA9X9
i6EGPuVVbye3QnE6gZXzPbUgncc8wEyTzgOdiSf+XOVa/lV6Kp553whnUstq2a4ilnlGUxAdoSmy
cOHhn8iOfdm+zukRmdjAX8SZqEqmdwzqlZrWhXPbHc4kDoI1IAaFSJ7+FzPEmhzPjMrGX1aGlSjk
8YWAHjU0LcaPxBD/byYWu6IpGCUCIb369m2VyFFGI6n2Ie2NUEpmZebPwG4aVlBKh/ktYuubVVJB
9cO79Kl1C+u3DN2iJTNmpT5GaaBNkr7vxS4AlobIcgirL/3zklcJZkNpgPUqjlZPNPhllIqaoNXg
+gSl63u5OEU/OnHfv/j2wamXX/30FmZhORlq2Dy/AIKv4ZyALYx9u5W9Tfl+Irp64kiPyetJ0xvo
M1buVi/2S/CCn/CHgnW+AusZm4xXwfnvd4LznKzdvBT0dZFaiesVlTv3lc+kn9mgohCxboM/F/5g
AomlNj9Pd0+rJ7gbCPsPXCVOks7c31k6HG6kolGqRAdLIz1Wnpl7r+uGnec8A9lEPuxWs84TwNc3
Xeeg9npQV8RbRWI2gKWrkvUYCYaytlsLfsyNCLfGji7t4iaxfWHMiBuU6kIeCbcjooU5Vm6SW5aa
uNboxDk8z/7T6413FnPR8zfYsf/yL+0mt31LuUmm2DFyghhxy5I2ZNBGFCq2pVcAzKqANLbyNi+V
luWB3E5LBTVLn3lwK98WhPQG4PtiusEd1apmhI/OWXVDHKj+n9kqH3tWywLOUtnQWH2nt1YTWHGr
5DqQQZj+VuZYUH6ep0EXAhDIL/Heatc/zQY48v8rSS75FbgDwxLfeaXXLgSk6CyWw801boM5ZADv
MolAAvI23RUnnjdrggEeTRTjhOqDhSZ/GiHIW3yfH70kcAVon7g+d4GNb2xgVIQEMawZCmT5cRD7
vKIUS3oN7YKNYBBzs46GiQ5daxNlU32ynGadd6zzWBy9rNT2t4CL5pWSojBBuerg5DyzPBBIurx5
nTKenBU8963BCw10CenZqA8msGWgwZNVhF9ZEilYCTtDu5CmZyqApFtFuNIzOhcJaFyA7bK2tOTC
lWF15mMhIegTQ0521xfQ+mT/BKVGC2yPInIhYg/+Ux2ffHVBYIrs5dMc+g352Gf14N5VLoCfA4gz
l/TMc32O9yHlfCE54Ah2GFkcjNB1IIALf/C8cGQEN+ePpgkbtMML583XBNO8+9kZOZvNJcFuQCw9
ZEyiLpOqNgG13i6PeWQT426djuwcpflzBSUdJxsFcYPmq7wk5DxRmysAuYj3ayjpZg35V7/xgVyh
Ror5bsNF6Y4aL8u6LVYOAe2Z4k9nssaVyxm+0zcthY3+dKdFF4x6E4cALwX5IsXQBRjLD75UOE9D
FxMKk4/1UrmZ/5dICoNps0JuqujswEdnpndjaUG9VD3lXvyKt3VHPJuI6uN6frThdNZ1JYEjf0r2
9dlNIbBRT4+ji+78tkUPeoRIWE/a6VgHAdrdmFTxbvjqUQZMw/wG0FZq7MafhObhtb51aNdnHqFU
a/EMkTb7WHOWpnMuvDttosToFZb6E1cg6Hr+/fL+rAiqs69zOkiJjDFKhJIBzvWwuVKPrd+JyOc8
HookqRDMyHFKkytNgL1+W300VuRAiFcN0eBDgkHp2RN02V7UfUrY3QQmMet+LF+iYRfYauVFgGTd
DcNZ28qTERqz3gSpfXBs6ZGW+528K/wgP4YmZe3B9/h0r0ZgL62nfMsmsGMX1Tc3rLtRe+fg+pgb
gUSGjQAIY3eyBDkWZuZ5TqvDagWh4bhKgzT6TGSki5peeuY6P4S7qJMvWsliapEFwoXIkwTMHFqh
MzFCzfLqTosihWnje/O/7CihssOhgHTkzp5kgR98VdTSEByY/c+qCnn6IJjwTuN5+k/mRNw0jrEz
JyyBLkeL1aPUhhkoXTpaANHuM3UFnQVy3LoZGZ1X4aKmNoPAyFpM7t/JGB9mmRbisq+okHfaprwQ
0FGnnmslSPHdmmC/v2xNZtksWg7eXDJ4zpC+6VawcMN0ipBUhMVwzPBdBX1DHBAin9JQtkrmhdYV
FS8GiPI2+OKhIBxLYvC6f5BQJ8/wexHUXu4HSo9jXE9o3qWOr7surY7esYY9Tz7jsCY5rsfiz0Ww
Mzw/RffkbxXPdSxSJSd6S5KRtXrRD/JycSnwVcTvdsihlBH59H0JPS59/cdofSrJabkrZVKvUxaB
Pp2CGaas3SLFk4nlIzqh7Jgy6EgnfBJaEFINj/MM1rnv7grCrVXZFJrFV50Mlx2YBUv41dHsLi6b
vah5QaIXx+1vumXqZVdFM2yxcxzQascpdIivyzckth2fy1WI2MdtM6zGn0LiuYOfwg+UINuUcGQn
qLk1l2oXcazfkPMeJgbfaiXyVVP2iu0aakFLfTtXVNbOGhA+cDWLr/LySVEZcCVQ36TD29uwBMEz
QQnhbnZoYA+uf5im4Ial8qWvRwK0qDZGugPXQjE51NUVrxoVxclVxFD7DIms/RypCf06NneElHaw
ZAw+9vlBry0gjICxOf0iq0diF0KQVMDaaw5oaCavwLRamovb4QmCFZRuSe9gD3Dj447gKJsurvAr
gnW4IYS/l2t1xfpQcbBcFR+SZCc2nsnp/fpt0wYBofOyE0GXwMKKfxbCVNYhhg9V6Csnv8ksNfcY
6rRgjxqv0HEgm11d8iyWt7GsQFOxizb440n/0XDI1eJAXrDm10uNO1KGlUVlBr7F6ZihpZ42v40E
gmQfSQzKQKw4UKiU2G9I85+omKyzYfJh5rDj5TGjApyTqZsvi14SK3pM02TnMMIFD5cQ6vRZ93b0
M9vLgDywR5m/ksLjzjdHKolT2K9d1Khnl2b908fzPe6FliT6ydf9D2mkGpkCcDnA9avFTU9A0sMF
82dRMtC4YX1rbyX/ouFAxhvHzGgHKohTMBihGQKgNtoDTfvg8aIc8uqOI0JdCxXBRanP06IXOgSj
iK7A4+xf+meNWH6iUvJHkEtnlmJv3OwAT34H4OVL40ROzc4OXI2YsQJU+EHCRS2jeC/14iWZ79ft
d2zlsd0Ga2ExYkyf7Mn3d6hEiJspOt2TNMeo5cvvucqqmf3pdOKNBw2DEG7B7UkMYx18uZtF89lG
4SJvDKIR9DmwOdVpyM+ROd0CT0WAmEVOzWVonNlWEiaLatJcIWQdRZx/bh4Ibdr1UTg9Q//8xq1L
dYHGfKQM0VmENOzEaaQVKCEmSz2ehSN+7pFiZO0fNv/q0pxpLnh/JfEREjj/gEviL3Jf8jV3zaxY
eiwH8oW0xg7FWB/qTRQsMikjx7MoKTI3R4VxxT37wcuiAbZAw/3TlvP3N4NC4FvrNyW/3e27oktX
8JEA0xwhjg1+7u9wi8IJ15jHlMTrBRUC8eBaIy3pUtx9fuET3wTHGDJzRKlkszp4PsTI9xTw9TNc
5RpRAT8438YWLT+xzORFE/uuiO4C8a/+WQTqBJ18THOlhMuiELkrVnsNejHDhzZWBmZtMjng51gt
yMd8gbL4eROZZtdu15OOW1DoYT9HXyV79gQvRH3H8Rk9lgr6s6q5kZ0p2IsDF/isBtjQ3hLivZGW
spomJR9mDItq6Pf2YQDVsC0KbG9alg0G6cRcMuT4QjAueJvQQKTdoXOV8cR2ANtJ9/Jbph7f4e0k
X26HbONWTphVFRfstTzLBjqPfm6vygJ3owplSaqbqMYTxLQQUfuYcuKN2bC1edUhEEsP5D6sFpxc
w2mDcUtsDPpLLJEgYujPe/uoK4KEIi1KGSKfhNbYN3krfQOCXwFQvf/7DRohy8w2vww9baYFOcUr
oUfMTzIjOm7KLSIZktcqNwixWHfaz6cnTJzwfkCNoN6STTgjueQF0NR8JXs8KxuI/2auZnIk0kNE
5iYurxoXI3XTvSsOSBJn91+Kv41eE9/KDggVVjzG1YTyNLObOw4Xc8OvTUgP3gZzt3itAKQykjnU
g38rM5ngaOdaZ4tJX/yfSXtcW1WGzKrSEOflS+ya75IvfUe142eYLt2UZ4wyxQwAyj5JnPkkrtqC
uL8cY2llzmvATNPocZsE6x8X+H5O8odOdr17+ckDS86GijR/xc76y+sm8aAbgeAsWsoO1zvv7gmK
84iXyGb55NjvAkT+xJiJENemUec+zljPyX2eJsbPFhWDWuGW131zVCj+hLBrvq9pYkXaF/4YJra1
Y1JOnpzaYL6MmuMdGeW/BPU/ARo0pOdFFSgekoEdnP8wwrrUTZ+Xnfvc2oyJswr4/xxZXnUGsKb/
/h7cSWSu2Rl9iEOvP+A/0SPcdLDwnZx5AEJnAcRMSTDKF6E8Yvu/aHzcgNZLj1sT78XhJ5RPe2mS
Uu0LDPLXk1ww3T6Kw1Si8uPgAYypbUBn/MksejWj+uj2Q56MI+N1dDKrW56cwtWv93tFVcpx2m4D
zOcrNu5fYO8uckj2uOCeN7f6wpxmU98xnQnQ0FH+K5mz64h/yI0KLoLvXzf4vlHa4FB3yHrvWdeF
UA+fXTc+cRUp09oqj3w6rEKlqcx7iu6WRNOAiR1Og3Un2aY5Mh5pSxC0n9xq4thQcFgOXyhLUxEa
UOgxmoYboN6zC/dgll9j6WfWLGUGJX0DyZB3CrGR3wipXGT4quqtn41i+unSycmjqFB9EPDX1S1Z
6w7SfR8fT+QOGeIvSSdNZElExJClJ569p4m6VbxfbDLs0Q8hDvwA+Ljv1q+b9+OD5LP8mYgpZhHj
KYq4duF6aqYfnFpi+D5891t56R+PjyZ8FUw7oF0ZhqPWjBXCAS4+UetpV08Txkgm2MBjgQl71h+s
IBvvF93VVNEBE1zgaHOaRKPw1h2YxxLUZJVGT0TG27LElDn/e94DRdbXY0Sb5oGVI9PF+7O9SiqO
qZUm0b9hizIPVrtxuWEe7B2kpB6Kpm4/Y7SmXFR/55Td9YVGx+/OelXQjX1PfwzUKBlxj5zECkhO
rcohrunwABdx2wZFwA5NKh+SHssOtybwkTQ+jncAURxcGhPxhIyMCrCQM7Y9BqraypeRnifENWsb
WnnyZzappxq25uVbR9OnVmuEVCK299lGdJ29xRz7kepjOBZbZ9kWoky8r9HXcMhfOfSgPGOd4Bu8
Zl+tKJaMgfSU7Xe6wQeKFAvCb6VgZgFyWeA6yC7zaxGpNuREvLJGRL5QON7FFpbnnhyeQaC/Kx+N
IixxXyqS/MJ/AotaibCHN009Cy+IQEarYDheS89NQiYgk38tSjYFG+EwApXWljgnG2eLX72dG/60
DY6DIC+wavNmE8rDJPaogFhYE0icXSrobUL9Tb+rH0RizNFVTRL14uAHRX47tq9y6oRIKzoprUWr
VzalcTJ8oJNz6McQ8tcwheECs/fiGs00XLPWehvsyp+mM1N8eiONh/VOSGdP5DeGd32HCXv0BnMR
RkBUvX5JL/erpk0aafO9Iq8fxQ7t5r0IYTSzqACIK+8zgAJFt8RoYzVG5XTFumA7EV2qemA6fLWD
giXMcnTbOvk+PbLqUFc4IYTbuC9k9R4XKFmw0Nf8e3BJd14HuX1gTqPpLXS9V8s7iKdfNw/Pj8wY
TPVrBWAPyreg+ECeGFzc1cx3fJ0uuMhcaofw5SR7pcB0TaTpJvtrPysPsL9T6C9JyBZAKq250PGw
MCxjaHzMjL+jEejyhJQlPTfgZOFaWRxhFeBJjy1wwGuQsGA+TGViBjXKu392PKxtKMI2x25on5XE
mKNbpadHyCbQw71w0UbGNvXmF6B4os35y+nJwc6l6dMXCiHZ/y5/mTGm+etgPSe2Wgz4dHHYU98m
7LJz40GHpb6C9T0UAqpYuPYo+bLkpgAM4QcbS0t3J4GRUw1VQVjryURXuJL20eZ+vQ9dxDWgYDic
gfOdilA9A+Xs2wnnESaYRKA4JqXcX6y8eQxY+onEn9DP75wELpzdlcT6HVb9MsoptPklU+DvaqmD
7pq9ZFXujpu90za9+bpmq1ENblNgnMPDtEhyxaZxvIEZogpJ8EpYxntwaMnceGjafuS7mvSR/5S1
RIkoNCPVemQJ0M4yanWdneDXdsN8iOFX3/U/i1lVs/otQO0hF/WP3kyG+fLEZ5lFjAvw7iyWcdEU
kysMfq2Ub19idVxOXse7F/79U3tU0uXY5TRVmU5TIx2fllWLsf69cmRT+OCQkyshE7/7JLUSm+sW
tnq5/h9LZhkTnrw9y1I060EZ5RXl28o1cib0N72o0uQ8IWPrSfHko1tlHZWNet4PneRU6TQZ7RYI
BTtcZugIuOI2rDyKoZYg0zDSD2gz0DbJSNlcOWQfy5812m6qXemm9Sj6kRx9IlnJmakMByWGQtZB
Qjt+pUppccYfVFdJMYLfsulJH0Bp6zQWmY6opZNWSIx4ppYYDmybD8fyuUpcEJzYPiZG+QlmQfPf
+s9s+4lY7j5ZX8YU86KJVo5mLUDFzCMtcB/mXKCrRpCs01R7xUgPPQWLDxXDmhNEFmfggcWWQSup
DPAa2FQbXHxsn6XjJQXS125CjOttSYpUmsErlrLhAumAkwpL7qMU4YXpffFJTwKKNRSTgmjCa2bl
VXDgpbTK/8hyNXPt+zi6SU1yWlg33uF0nlkY8muv2AHbvRCy7Y5QY4ZL8LXRckGcd+vCGunLlYzS
9HORax/5+Cf2WbIATSXJMPEnlAPbIjnbTNZYxD5gh4rlwVEiMUOEt8vRXyS3yJ6v470Onqwr4juK
/HkCidqmnqJ9tOLURzcUtNWIG0S7zCrD5DpTr/fVv778oTD20/2OMHnDfhIjLNVkWFMTMSUUJJcI
c2QhUT/sUTGnsydZQg1qAjNOkeLcxLZZ3FfJrnuZycgiS5X2f6Czo9Szfgfgj6dFhWxEyZrtPOZF
JmbMdQi32UP3bzUpe1+gke8P/UV5dxJBU9dGJ6JsRANYRFVCb6bow1/42pliHdMZZNKVzVxfjJVr
4wrt/oBCiCrDLyR1SQNan7t4bv/DuQ3czr5AL4z939RWc+TsHjq2J4Q23KcRBHw11wa/QT/oplGF
S5FEj/V1bW3nboXgTxX2Foznj15iA+KXeDSVYaJWhFJzkJRzUETT9N38zDHE4aGVDKQMUm3cuUOU
waUzfGX8u0KFPWmz3MQieIQy9fzK79Ns72jtkSz3NVkyAQxbDj+lIRAQ5NKhzusL9cAydzOh43kQ
qNqoxKq+MIZYauXwVaPOKeZn/ZWqGk5oT8kr2FIO9VRTl9kjR+adaEOFHV9xrjF+CMAYxf8w9TLi
OUD7roC18VsT/KQ5fkkEu5o2NaVe2LhavRHd+oLVcQ/20gXhI2Xm2Tpcq6bTkAEh6igcGUkYIPjE
mmSFtWJHaEfQxWEN/w1TvUfY9PZNnwIgZVog3RNV4vllpFYOWO+UtxcpJclONoEcD+z3OvQhdR6v
gjs650wfSDOi556luFddbj7pDzT3gw8SXtGSYi/hNlBtyKrWEbgSu5SY/wZnPxkuX0VomjEjC2qv
bTlzeB9d5Bp6oMdxhWVght5sqJ33M1JTdk6ONz54o7XWvsrKBHjoWmqsYYnZ7FjCEBzuztpK//3i
rBU9PgFJisuh5XBqhR1fqZjrttRvRCGZilRZpkgItd/u8IQKBRKb10OFCcXfWz812HD6ovyNzdrQ
316KzXClHt6QH6YiWgAMLL2w5f7boPfvUNC6iX8s8T4AkfdJBFWawV7W5/XRa5uNzGffo1NHOPwk
T6ph/BIOufrnqKF5f1HjmxibBiaQe0maUg0D0uVrGwQSM6E7R1iOr9i1gVfdq+pn59forphyCnjf
payIzNdtu46c0L7Pil6s52r12m0AdertxXu9s9n4GPfqnN80jkzu0zI7U2JYmvrr4xHTB+bE9IEZ
koI7lcLC70FS8UKpsMpBLqENS1QZBnBzU/jWUoY4UEVJLFFX5xR9XUtckgXOFuiN41w4cSQyc9CX
D5iJ0jDDz5M1HHUjEpdyzHZbb1AXIwyNbDC2K8A8B610FF+KpxvssRrsuIUuRZGSV9PHW1/n6U7N
IpvkcWvH7DeYpY/2I2UsuOkyTEjnZYjUnbZ6lpB/2L3T5ISP36jyH5j5/fwt1ULVGxDTLu0UcU42
kYyBNeAJ4TkKJqMTRlmm+BiWYA8jpdUPK4538ygwdJ93iBqTgmyq0JvPtfHLjhTF2xjx7cCTWDeS
ESfksDUi1B1xkn34voyu7VTfA3Bej0ZVKVvlVq7MAJILVfKf1aYqc9qd0mKptfrLIHLdj/mGykGh
59BiTVTUyRexmFqfFhhfTHxdA9pp9xd0HLYfWL6JRbtC786r5CuvcbfMdZbe5dMNzubQDWk7abxe
TvCc3j+sDnlEopXsdoInmXqErXfu4TLhvF0f3AlOXqgbKucrP42CBy4K36yCnWGm+X4Gv2Iq4Izc
0bOoGpNiijVet6R/fAOcTd34PV1+ggHPyOCynuNgbMknumg8vi6XwammOGxG2HpnlhON8IUoG0Ms
GAZsFlsumDahB2t9Wu9b+igx/BCBJhIF8+l4Lc2iLYOL8tB2zExM39a1hxnfUJC62olsogb11uQB
YVOQUp6ihf0MdKP96t1dnYUypj7t2s4+TJwOirEGxp/96S6Pc5vbseLP0mgiQ2+cuzji6D/VzfGK
DzKdzi7QwpNfqhCuDGqETPGDZ2kMMqvFJBE5eEuRDnAsPz3IBwLYlTm+i31rUH6A3RLetElpElxr
IcusRyKR0OzUwNqXY0cqrdqdg6zmB5pGqpaPod8iiZauBeVo3jp8XKiebW0Pm2/GWzhCUxKikCy5
ssnNbDrDEpsy0tSbZgJvTDZVTkmv8lpr8CkoKKyZ0ybmb1ijNJTtVg+x/mSfVmCzAncMZQ/WMQ12
HV9uITWgFjbaLDPoHBGuZNNW/AQTk/ZmkjEfcDngOhHslAMKTPiB8QIdjRl9axwWIOt1rjP6LOjr
ZPKlHu0EAhX/bO+f7x3sQ+WcLKCJPiQd/bHrNiRXNnNEV7n93HL1sgun9U24WtnYSAHH3eYFGYh6
Snz2bT/vJYH92vXIgOrJahzgGznlXvUArtyITVk4Fh+IoaUtAD4DRRQILYGE0A9kShdfndlyoiPO
Yb/dgDeae+LhW87k2y2Qsv98Wjf8Bh/8/7zZ6AGQrwA5O+0lI3RKzQ9v4xY1/5YCrHjRep8cZlTn
uQei+H9iaO281SB/4w9ZMc7lHeWYWsGT/gGU/yqePKZ5bXHANUDBbdw6wZ7RNYtRKKpqcUxvaPSc
NG5cFX8C/CzccaDYwFFeu7qcR8IJ3uvSdSi1WbJYdusP4GZKpk6c4TtyYIJ39e+1pHJWJnPdGGJn
ha6nS91TKVPhjRKlSpokBerXwCannpPdkyx8x24fj/jv0xcHz6dIFQkwNJX+ob9jwbaZSjb43MPf
vF5qxHFsb7jJMtVJNV8XkaSXdKDonsPx4DKLVqE/0y9P+H0KRKJH4gXRp4ZCFNhB1+KGC0EuWvWj
Ed1CugyRrI3UKSxGeO64iKUGmBQRvH+AAA/Tb2mIK9b4NM0eET2nMHtc+UkaV3XhNOXXchSs4fCD
Dwayel8THjexn67Zq8ZSSRgkEp0o8LvhzqGIy2xyk63IbYr80g6XKEce2KMnsj5MgM2h27SJDgLI
3TPdJtin25oVHsd7NPE3+MwuIAX5HoLqLzL63hwRlUblJW68uQGQmn1UUCwDpd8DZphB/B2PpF+v
PLHZ1sm0fM4Dqmzviv2YkLeqjFt5ZnabWEJowSsU3d1NcxxPWZDkJ67zbHSYOYRZYX2KFxTbn9qV
POcf+CYMzaBqBkanmAnFzOqby/ERUiBF4rmmAoMhyG6VSplhnAk/JHmIPh53jpuic5XuitglUJnP
KxnstLds0wQTqLLaY4vPJdo97KDqGFdTIbifsTwGCauv7fShNqxehSZmQxPIp2EjJ49t/qiMaQPF
pv7brRqJbaHf4aQrHe/M0bvPWFYnSjInhauZo8m7i2zBJdb85L2L4+H68lXLiShMJhTWQ6750DLT
Vs2t+VT4XvP2p6TxvYD6NrzhcGD2GuNeVaIUQAB1Ro3ji7nElAa5/0B2dV/sL4rOPH37xjF/+8/2
133z/9lXq04FDD5Oq++69YFWf6ZS2DeUv/3QBKMaFQ+VsPqKaKFnPjSFQDKTdXbCM3jIV62Lefne
BvQq1iMIli784BulXewpOiIkRZ9RxcZYehTn8j7kFDBcOZFYIXGChhFE3/CxsZUxd7HwFPmMkG5i
51GP9MCDP9QT8j7v7uIfSAk6low73YJrkv/mAjQLh/XTCHA7D7uKk/XR/xspgsRCvS0Y0TczjMNw
/0Wlj8AF1r4L1hF6YU4duF8FXh0ANBKernBxb/gABj19Ow2Od6zwu4Ufl5goBqmvUdYYUmp+epKG
3JxSWbWcDp9t6B34UDYE3AzDTGzw4Sd1xirVuaFofdZbVopvD0U4jJR9bnvm+pHOJI9g/EPsylns
lDGyLgYSU5WMLaGXrZk37BAI7Lin65Yfpm3RzLxa1h30xYaRKXTeLP1dKSQWDSa/SpA1ETzndooJ
Lb6x+cLeLZA2tvOz6WAGfjtJQ2qTy0I6ZNlZK9HkgZ2SdZJhRR7KTkDe/70Q6eq8tu682VVurdBx
0BSpV98HPFqTm4HllW21giSq6qWjffSir56RNbetDUx1z0ITr98XLKEL+hn02EPeaAPlhkom/iEr
129NoWyK/eswzfFkInBcUGK1u+WyBFyVAeb7FkZTI89ZYuTpPcLMOJXZHtjizSrI4JDTd68yogqr
3fwOuL51Hr9MHg/yI/tNTjdicpDMLZvH++fhrKRU5Lv4RleUaVUU/vmHSbcNSYJEA0PCxxxAho3D
fHCoyLPq0emOi0JKWvKdXQYhgnC1e6fAB4Hv3BeIc7wX/I35fg18NJhZorHyXqJSMwJuy7wJ3V4+
4iuQ7hr4sM1daD4KXPH6VqWuvZuXcMgUqnLdfN1xisFvLNTrXbfLfKK2RxH5KbO9qHKs/mPIgRWB
+9zdj9Ygle45uqxyKgiJ7GsYGUeBCOy2B29IBdb7WV+zme5sP54RevEjlhr7FnSxZKI8bKe/ilpd
C2nHKk0R7uj2yHDCmu70Y5cU65HG1gB7v8sR4Eqg9wxWqzl5aDIWN5J2rj63DJE0TlD/tvvsZyCq
8lfdVgLpwP7FoGH2UjY8/VTCZsEIgPnCssCuN9DgdctA81u2YCBysz42K4O6yacJffgYUZXKQT7l
mR2OGl5oLJ86nMZBpDwBaZQTJjrm4328MHMu1o/qecVweuQG3JhxDJY+IdZ3ESx+21zQCWqkwGfL
vPekga66DytEFKhunfNsRRROyA60WOhBQM9Z45j0+n1NAt/Yk9+1sBpysvSrHwau4sH/NQY/L6jC
WnTT8pkRaS7XUyKsLNppuJIdCELZ6Vbz00MdR7isDff4DT3Z2nrPWF5+033+3jtotiFySqhzJ6h8
zkK3Mz0cZfSIXh0AoZBeaLJ60y7bDHcAIW/cKCJVXVkQKytxBtO+xcK6cBRuRoFXyhl3KfekJWq+
IIIzCLvyUp0Wmx5DK8tBDr5S60YpzX5gKleJ8rnKXcdBgOsDWXzYasiRymo6JXuLEPmTOvJKBSHE
mNL+vMaIAARgtVNcsvX9Vqh+iLavk2NoOOKOUQ5osHytNnIP0jAYvFejnWAc6FE/OLuiq1W0Re8B
uz5N05Fakeb4Z4znQIbiKPe3AIm6ocm4tFXmqQ1F79w9fPkZnaEBkmo6gh+nN2MY+CRp0170OXgx
u1UHUwLWESal78xcOn0JH/cDsghCFsPpjtUj/Adh/re5kuR0sCeE+9QICIItkqx/Ra9PwpQWoaiC
58THE3qP1J5WM8biW127ezzpQiKf509K0qvnQ6Wcr3Tu37sHPk3eC4sxdwGFEcAP1QQUrG4AenDz
nhXQjXdZSUwRfO1tJLBR0JVkhYRZNmsLWZwJfKsgDfO51fKkqqr5EVQaCXlgKQHmG1j5h0C/GZYi
K9PHwjLfYYRBXaSDo6jHMPGQBGXkAnDZyEPpPozOAgrmh/RBV+13dWnqHtO7oD1/MBhr2evOAZXs
9IVjm3s/uv9orfvFtKQIla+XQ46aBoigV8JXuPUGZfo5XKb2sHgWKlgBQw6itMR5Lm2T2Cp4g7fb
eAFgj8p20k4bzucAtij1YHR9LlrYV4vwxMv3taHA/E6RHXp+FtL+0CDwpENxl28RbzuEJRWgB5i7
6d24rz1rzZQzFeWj2rXswf0MKdjZdl+vCfXvEaYR/fk70QZBg17V99BE35aXHsaUJcoyr9ig1ign
gZZIGvdEdVI1k879V7gUkpq7rboNmtXI9nnAChhhj/zflds3UY5cOcDN+t+z+WyVADRIAlHc0z9+
54xlrryNOOwUCFbcFGpTYJoCP+5AzoQQisqRyO3dW2xLYYUIJ0zUo5XcAF3jgjJxs0no2R4EIDoq
yNfx9ufHQvA1+UcAnT95MJYENRRUJlMJp0nsH7Y0aqfKHa6osOaY00FdPDXrCCFQyUIANqKWXQ3S
wSYedqI+4qvJJzo7YKpQZbIVv7UaRf/RfNV5EvoLnC46cS4/UCypcyAtBiwNIzA9RhVHuDFcUxZd
1+4xrsyci8cYCCl/X+rSfSV14MdPfEHXGTlq3L8JkutjaNnrMDx5Z/JeK1NBUPaSD9Lvxol35k5+
QR2pXLrvu8/YDo5KX1nH8mFzjjF43x4E3eWdCtES4WISr8RaE9EROvsgZbWW9PqCbQhxu5eQaZx6
i2szMpdICoR6IsiLH6/faaatkGrseA3gkTkmIDSTmYoRPGI79WhLE7r36V3UQM7NpogP0nEG3a+7
5X+U5DlPP9Qzcx3/MdJpTgFkAVYuCY0C0dZJoOa7vmXIVR+vtj9NwrnOLF75+Gb6hvJCq+AxdKTs
efaW7EioVe2HESVYaI5N4BIrcLAAsmkz2HmPOvgfIupnu5obNsuSEN8IrSsLnrgEDJj3l5Nohy5q
ZP2H8uK9uKTrvqZR61h+LvdVGiPHOHUSK5PsHiDg0vEUcQTGqCCymptCedGX6CDtR/OrwTNgpuiE
W5QB9OS9FGg3JSe4TR8fA2aVYuMBwtEzMqs4S6moIew0vTKeSEuElMt/IGqs/GqJk56qZOkI4XlN
Ac3HFHJ3kreJWer1gEHvxhRnlaDMX0SzVb+pxa9HE5d881jkgnuP3/WW9Z5+NmcMCYGiPsTM9KyP
DixbZJB1L2U8l+CKhO1bCJKg4S/lMcAUi5Y3Avgcqie8UEQF5pYj+WTgv90l9ajuHz/68grY4aZk
OzUVJrR1ZG3ebw4wrlZc0w38OSawxns9mrGC+h/mjZO06jvIZQ5S+sas0Q9/nCCMF8CwvbNIFGl+
2o9rpN7QCRFwQERiAsKOp+kTwl6Gfe48FMVO5lU3xVzzKLNpUvPkRRC6vGIIHIlustwmuE4rsSkm
1eMBgwreJavlYzyYhoP0yXxvBAdNNu0NlyULhlifBSboMJvzXqpttOitKFByiWExeDn0/3Aa/LGv
GyBPYCDqHFtN6bDWVexBt7pPt/JLNey5LbcWLDd9KRwe9zZo9vkcjUZptICSnUqL406tncM30dXl
Bu/AQ3s3aw4WS88kDLUfXFfAtzaG2513kzkmDkcmzVV9foB5YnOkkB5X65YB5jYpgX7elm+p3fTx
ydykzoIwcZ19zNCz1t0sDXZRD59COKsdRue4znj8392Rqhb4kc6yCC2dNJmzFMHXlq+YXBPPMWRN
vpejuIr+HWJ+P/5E1ZSsS0LMgO7ja176j4r63+UgVCT/xJu+RCPGeB8z80rRjE/tsIF8wqxwUJ60
6TpU1ZC9MbSq+lp4tCDFfK2qjlwhUxbZSNEDYghAZKY3U+dYR7KGmd7NPSjZxumKF+yTSM8Tdvwl
Yc12BGHNx7uKWpnVtc99paRffbpKq7OmiwCMjmysG/pW7oAYvsF6PnD+03yncb5JzEVwYtqXqVzA
Up7xRv89pBkh2krJrHDMJ9UkB6ftRDoHberYTbt1NYCYZt/QpVwqPirdOeL2zT0bdF46OGmIagIF
C8sfA6lLcMSrB7KO6bkSK+XItVGuKhy2pyhk1vLWOX5BWF4bRFkPByncXIoK7sanJRVyZl8fIPjN
7kTz9sehopbaO3+uFmsGObeQ1dQIFHfS4sdFx6J/rcI2xqydTRMkKhNs451lfz5a0p/GvPoiZW9x
Bo2zRVVbi9nLelyFQyQvn7o+hut9udiQEhr0VZAX7zDXgErTg5VKCsVmhXRgt8fxx6iu/gzp8dfC
WDrQxiPw98GSnIojOHHHlF8YKGHO6FJKm1HIPLVrH+JlcXRv3wPRNMKUxC4CL80OVX9D9x44cXJ5
I2kLxNR68vqHA56AmUBR7zPvv/4VbnmcbSJyeL9dg9jGQz5YtLlNPtV3BOnbmzxjoY1RLbB2TgL+
+mvgkeNCHK/LixlvwM5wXC6euEQlGuxf3vP8yY5lXDihuu6wJksuq6kSMXZW0yuTzGP3k+ml+FUj
MpHOV6B79YrAOgpbTRksKfn8qYqdBpI+AS2BFd9RcxzExOZPJ3I3Ceb+Y/4VxW2n5WKgzJVGzlxA
x1oLjI7PAsSL2SfZFM92OIpx4HTutJtEbKtg0X3mcJA/ZnzNA/PeSeACOPj99WPCHLpLKn30EHyU
JQ3oEGsel9R4J1H5eAfJ/0X8dleaGAfm2XKWuvpCNTkbr8y9JvhzBYfzDUM+C/BkVnAIc9kQRr5N
Sh/Tkl8yVTnYJTHsOKT/VQG/hpdhZzfwuNVVOewF13iYBL0JveiIUrBkrHQCr59pbqFjKXPZZtxP
cgNjruLkiwjWsbV7aQfmcsh26IOhW5iAHpCzsiT8jC3G0w1jp7bAKf7XplpkDM02/R+I1Hozp1p9
jqsLibXKtxzHm1LkKyAQIsr175MdoRBrPpfrhaZe0ipGeV6PeH5DousXT4EzUbvwVP6DrC4tm/Ey
oA1qwePrMFlkw7TkYbyPO7Goq0Bs3Os39hBW9Vj2aWqtb0VkysEnwwQI+bY0SUAZ2FBZLf5HlTrC
Gd6QqPK+KsMkGm6VEQ5EmMpUDJBOYeqQKub2YowamHXKcSevvdJDtfv/oV3XwFRLxuh6yIdKtaYd
uJTBq4jhiPTAYpn9/ltEPwMz9ayn4X+OdwvZNlC9ae+IW66SAaMW290GseI2yZUKMJsl9He1Z2Dq
sHq6kTy+EhqKDN1+rYvujvcSdSxO68Q0yQJ5EnAr4T4EJZq1jYTX52IhsysfmkeqSWq+xgsv6bW7
+GEw6/4OcYV/A9YBrKWdDQ3gLlPwtqm7kByQsjz/XHlD+PEe7e8hcIwF2zGEOiRCldJ2r/U+dQNA
Uc6D4m/2ZiF0qgcXIWKJ2LhFsa5PN3ZAJq5fFqUflH4W1uWFp70leIrrNYWiIG2+ARwvsKlcETta
/6jHczNPGhHwI5iOrbEHb9S8bLWxSQIX/rHihf/g0uJw/S4I4fzG8ikljqME8dR4mdRJ50SOKPm6
q3Amy3Iv1/Lmr1IsZxiD5xUGIaNkUReKjPLNV+yYK9LT4REWbQwu4Su3hY5ov1Rl0oQ+fHmUagKY
srEn7/LebYbeo4pO2/GDyGFROTOGd8ZhcmjRNrK+yf6FfYAJqj88unxtVteLPq4JFc387f2V3nOy
B2Pxz8VGYIBs/g3nDIV8UoAdTGSXJrByPadHrysGS9+Ycd2BSD8FpC+SBbYSf6jxsNBRJWCPGoNB
skxcpSFKN5EemKAj/WQYcXwmeVTTFxbkhOLmWl09zVMk0hym6p5pu5pcqjEOoGBdHfViu4sGYa23
r7atluN/kps3+G+iqj9qtQFBc1ZAI7b6T5cQS1VgT9KMMh9AmZEPvJ9ooTg6sLWZddG2zb6K9HJP
8xpCCkNLZGdtZRi8hTndn951aAX8FHbtZdxDns9Qt+69X6QxLsrxFlp+pdo30kTjXWLqNSQzughq
3MuhuGPTaVrPiXy+GY5hlGE+p7lv9Ihwxf7jl/ZlnO6vYd+tYufnahinyXQVw7MZn9IXGGRv/L/m
g3EyP/maGJyO2+ivcQN77pOx4kc3GQvxB7lxabyi6gwolRE5BmcW57+3XCaGPLkcM1iOzdHTfHFu
+iEgfUGHQ1gKqqssv3YrJ6j4oW+v6CLZ6jcqFSDJjJI+8VYVtfdnTtYP4w/31nOppYHOZ0k4nQkd
h7L39UcE7PO4zKZOCTtQa+Ot7g4fQWsqiCyqcuyAc+5bBT4U/2+tTbQLALUL8Wqo298w+VyExrU4
ZhRWAgdXUSmnzqpTOg/f/MZobCRVV/G7/oZ1qSHbf7PhpjZwOJYrY7Mtt/C7PAfh2t3gD5FMsXwa
BOcYVnKiXycCW78rxERHN0mQp/HPEQx75NKUm4PcPMM+56RQY1EdyB6KMPT/xWc7mG2Dnz/LEqto
m/49osBQWXdWf8AFSGk821QdI8RkrNS/+umMyHjWe/FhL6JYmKS5SBj0CgJWvNGquXuL7YGYlCL+
i8Z6d6gZG4sekxvu2+i45BvWezdXSmeEjGEFSXA13oA62q885XOp6untJDXSW5Mpdcu7YaXu8elE
N8oDr4GFgO7AxjjSQgFxEsknHCsx5NprE9UJNgsFucGj0QsS2AgqXnnwR7XGmaW+lJMWIlIw8GW9
A6zl8ukEPeeqvHn+uPnmzl5ZBVbcpc4Ewf1hqARFOSkr7EejDt7DOFQL5ki+SpokQuz219sYN2pU
vf8dG4vArwOwoeHpe2PS+Z65Ty9O0IUA36sv+dn/mndD+DfTVHXQaw89XF5meRq///339s0tYB6H
cb6WbPR++Lqkej0V9DWa90KYIZbx2Gpgq+2LvJnTKQ06neQBxurLFTq3GoKnQD6k0wF9eTzwAhbD
zR9utA3F5/j2m0Gp7I/9v9O9PWD31XPgC36REgYj77LSxFVO0PZjalQoKdzxCpqWNhWRRMMEMpWv
+AofZi4C1tu0r6Zh6XDFkP7tgm7Gs0KOck664K8mOLlUGJuZRbJfKYmGlLMgsZaBeMr/9zRWfrUT
B40ihbXSDytH7CNNaUXMPaPiOFcUZ7/OErCWIPrjcy+AM0HawwgGTmf4OvcSw08asfeJ9ABB2SjD
Oqbgez2Plh6ewLOd7SqKw9nKWCBYBe2a9IqAr7qNU96u1Vd2L6Nq6oInNfX6v5/z3X0Q0jT3RkS1
5gIwHHObiBGVTZDgTvGD4XemLtKL8r5xvcLX2GS/HtIcQXZ3vT/kvTmwhYgodfZPJBlvEHK6JN38
J06/SNK0BmI6Zik46U5PzXiqB/18l9ctWj1U7O8Ow+9gs4MnAeJ/PEhs5ZI++jEfV/bB1XfPDLp5
d/hCDvVuhPFOzFjY/4G1voIgBUpnoy2Wm1331t/XFRxgzwAxatrQ3/kl5i0qW+0AzrnKKYNRbGFI
A5wa8Wt8PXzI3QDfmNYoFKvGJ9Y9kSkvCMfVh/XZHzZf6McNHuUJDqoO8yI64vElpY0bzFRDS5OE
uKq/yYDXeAJptnEw6zKRW1a3AHX+TqAwKZt5a2wHOu9y+gwEsN4Om3q+d2lsYJ2tEPvNFNVyJjkB
k2hcRob0aea+pReG4Btb4v6d86EAobgKzSpFKSNQ+7xDjS4hCus1ofMWE1NfmnuzC7qCNDQ17CN5
ewc5QseBTQUtLmWwLa8vevKrvfrWGC2IPFCkogq/joPBiaRXiCqohsshc26adlvfqQYJCE2qoKuZ
NoYOr/dySUKdVuOqBlvzDl1/X1ek4n4dhhBf86lpnwDt2KIE7JirDuqYB5BLO0s/BFEjbvp2T/O4
btU7L8wcoX8V1+wsArIxw1QJgLyd213Cwn3TdUFHkFqLG4MV9SZB4NGgXCckp8SC+a1SFh3mTjRL
loLUT9ICMH0WfRQjwGgje3HdtzrFcsO1eET33R8jufOgXbSjjrGRyzyRMKAZKxyx8q4tVS5x+0/u
lw8CA57Ydbam74q+ahpHATfZ5toGqe4Kfnlf/81D3gT4DlwuVjRoL8GLtwH1FdAQb0Z0JPt1Ban+
Oya1n4acwU9ijBVHmHglxl2agrRLfzWCsBUkLhR5zk+dox+b6DuUUMvTVd6O0LWxc81CgkaepVlB
FEHRvnG9bKbqdDZFP6XZkmCCgMRDpcMFCz/cy+GYipz27+AvPXHYIYSI9Rk7tLDG0czO+dg+wLOX
j/DO2V+3b5cPelBCKyCcXJrccbahwLwPLN+uUuA14l2Tqkj/Q/xcqFDTC6OaK/jNDwjKe1RwA5+n
HncBNjdqi+tHEhkDWRf4MjCt+120aLTyd9OOjqIHoWSf84D48fAK+sW3EIr5iP4e+pUl8kzt4PZY
iRl33cp1+kcw+t5xySvK1bsPoDzMgtSslpSCZtCkzF7e/kVYbFGuNfMyD60oneSnZj2HuKoGUjvs
KW9MIyMiDiq0x4kYxYcHwq400HWSS1ER/t4Zozci775TAfjkdCSkVxygFnh21U/vnp/qXdGEvNaV
O9XpzOS7wi9MM9oaN3YyRztiFD6kukHaTgDAafPaFjROUcFCeQSLesaiPudEYnSoeucioqXz3rGI
9woELFwiyDSxH5Qg69epE3VixFD9+uoQRPS9GyPf8DS9R4lw8q3HVvwRQPLEyLZvai8tjKzZhR65
3GC3GZ9966D6qEK7uDuxEiTq/R4X5hNTbb2/xvEY00KlXEwExGMwo1wkxr/fsu3A8dSwvNfxvFno
F69o7WnocE8saXJ/cX6i+BEEPkzMQ4nwFdM0wwbnKFhk9oujGD5rMn2YDmKXjzSoifTYC5yKt1Zo
gI43WYYhqZJqpThxZTu5qGqo1cUWgBw9TVczd20bCiZd7RjUsSLKm4bo3nVOBbE2BUk8TDKTJqUU
7kLytrRwzROC+MyA8pPWfE6Ngy1EHnnu49qPqkToS/KzAszKZxSU5Bm98WmGLLPQxV4ql/BHWMiU
qe+oOVmv3ivGTKVCqQwjwHSwwTJdqNxBZc0KJhWe+EHfZ3gpPb8FK+d6mj7mAvx10X/1fNSQqUQ2
VfSIEYNZccPSCNwiiBFHnAE74EXsMnEWGuCF11o2qq5V+58UFOuemIIH5O3Fcz/q6tWS0Mcix4iY
R8/+W1eG06jbu4d3TjWEZuaN9h4L6/PjnLKVlIIfTpZPRPj0LBjQe5abIJMBC6jT1kUGFE7GUJe5
rgHE/1jyYSsCTC9G7cIgVcQPss4onwei2nFT6B8oaa7iMD1NOFIgScgenLBb7Q95dNhfhOWBhjij
sFxjV5/GZwZYY4TuSdact36WNlTdjcggaFSzCHya6rBghSLykWv47LmKu3VwncVZunwXw5+/hDsI
SC+5vB/a5ONKLI81eXO8x8U4S1TIkfwr483UCOgOUcLXniIMwvBWcnuwFdh51koK9S+LAJ7S0fjh
XehL1mnzPdqI8Z05UU5O9fmYOKBB7r7k4xgDsLFO7AN9MBtWl6b8m6Wt4H1Z5u/9xmrFqpmGXSdL
k4z3jFlHNiFGFyOaIYJ8q1Hj3KcuUs0t7kG7biJgncvDuA5PF+hKsEOlyetVc4ULRQ0z/j1dyhbo
3IDxjDOtaEKRZvernVFYyQS+X4MzR3tCLamd/KgM4sYZAMlejqsfXmzfpgNd13lY42xL8hFQXZmc
dskKyG/kW/5866T6X5PTEqszvxATxuBzNeqv7XhYHgsjMEzoCrLp6K8WWlgOmBOyrlG46uIfBxgf
9QDkl4ETuRn9ZwDD4YlKzyU0CYrrCjFRmJDzuvdzyXfA4LENaESUMqW1y/57tkj3o82FOU4RAdMn
1m4ZxC1bTGFjeOUYdmjOi+tv2M8N69PJ9EM9SkNnIuOyByviq16g2qOynd6HB1cDpHrg0lkHdOoc
2slITQBVW9ebaGtQ0tnAKbodZ/g05alC4TuxHTZijAGLZP0hWEyclMhKWi19lvLYPeJ8oiR/i1mF
9K4kRLDdHWSohj+BEp4Kq15+zhLQbmlVg+euVNyTirpa0hm/TRLKoqMRnp2LHjPS5uD+scSmO4Qe
psXdI2EXS9OPjHsmAZinSG+hY8M0HKHNldUocUBKYEw0ycQcqjgicCEvXhNq7VFzK2Dj2OOgTdVM
Q1JFfwQAnsh1LlmIAejnmASjnwIrqpAzGc8aOSaXqVwC+mZD7CW0tDg3La2m6T3jqc4jGM9iti8q
NRVa3ji1cMjBw3agEtdVKDP0nb9aC/4VWWvDJGmSb8hHR5ohQg1+43Eb1/3aiPhT+4tHEm+oBYRq
DaO4mgibyRCjfRl715U4cM6M0q7RtQJDl56tupYDh0ga25Bt/Z6RCOgtsfoWPyt4GUrnWLZ4d/D3
oxRKoEu+SAPy63JMBrk8skyFEom4ycU3Kvu26UjqpKeyLmI7nJxPAPSZtv1TqjItpsBQo8ETARE/
229RbQtadAHTceH9uAxK7PH5Bh1z0xy/682qfN9jOhTUGKGDvrKMlUdRE3asHoNCWeq2XN0FDkl1
vMPLyVmFAXSXqjF02eEDZYqms1Ldjfkrs/O0mxN7noAabqcCYHQBhN+zCXz4yiEsp/RBfBGyXzKi
eu/ebgFkg8ZlA6tLQUeXJ236JTaSOOWzDbWOpYllZbAO6gSuSdFYiVFjva2lwatiAEfcOX4rFCSh
NmTebxmdGcoXBubD84KpbLqjHVJXZRJC3pIJaHlZrLor9YXIU8bM9qcRWsABJQv4/dxqGkEXHK6O
WpEehZkGEMHb24EfVYuZAMcIEiv79gWDVam0QuLAX2XB4B7QbCPxPGGTPQJdzLHBLjqz1dMcnTqc
JGQLGgebHQwQdj8NtwzmNm/w6ROaMz4FvRIVf2wkzu51LYIqWZxNkxo9ZhsziCOg1Xy9jo6SPaOj
T4Ro1SlSILCOJcH49VVBTqYes1eBq3/tIGwMvvG048ugxbjCSVO5IKGW/UegFe1iNoEjE+VHptT6
RBn2kB1GJtPq616GBKlBky+EzhFfJG6ASUO05vp65VF9bBcrBl7nnU6fm0WKtF6WOxGdEdSHIbD2
vKyAHi6TpZZ2E6n1pJkJ3zV2wKfxD0/IoIzZb6WnFDVLYxSjdDu+7QFXBZAJNPjKfoPmJUSaazUZ
U9SiYs37MdhEoXdxDSILSY1M+JuEKSJXr+ZWKOjzz2JzX/L2JsDt8hXgkyppP2c2zW3aMwndTByP
FJiRgIlJ6udA5CvOIo3UgILzebPBjQToAmwO1sDJh1FdKUO9phryDxessY+aRpjZIyGk4+H1PGrk
V1ybnqplKRXvH4QVWmNc3/HLWTUgKr1364bBusINEy26BHaLBYFjnHaZ+ZYdJHtvx3yzpkEWU1vm
4I78sxXEq7ZqlFsE5z1YyQF3K5GMWGE5cQ8b7NPctJV4tnhAuYGU4BQ6NbJaBXVylf2LjGNBtBTb
8j1ZyorIEvQhODGWIPsF751nzpILOdBTFiO9GLrBb2nLxCArFj+Aqt/fiYYLlAz6Rdr7M6ZfS9vV
SruVw9JiLLxjFXGoTv5hsMAdb3kVx3ns5+ALxaYvAncQfc3n+qG5w+GaQFNGR2x0x3+KhLExu54O
EpXMS9gMAxP5Q8SSl6mEpx9u54I+l4E1KH4hm7Fe3TuF6+TSIh5ng5Tu+3TPW/7hK/TjQUItMoav
n74LLUJm5e3MYeCJrkHIkhc25QYJNgsNm134PLHFenhHnZrI2aArzGN9Oz2Td6XRIYwaRSrhrnKs
MFHKxMF7sclblQor9PpXzC/5O0udSoEkZR/LKVzpWZnYfO80IvRXtVh0daoqGyj65QikJQ5+lNL9
sXTR6GvXy8tT2LU5pm/hcYcDNmccDHxzo2owspNIv4O30RJHGNbi3nYMpAndFTAGQurxLDmb79Oq
+4R3EW8/rfsBSh6/BOmwpf8/I3I9tYkPfXcjn9ErMQ2oAlrNwbwv5LdEfy1UDl6YkiLWcQXsly1X
YzTnHl8Q7AyIBMyMrnzjbD8PkEXP1yd4GpPFql8+54Io7ByzBQGxEzlJkUxRsJGNiRkMGUwYBc0Q
ts4tRaQzDBuuD+lcO/xZN3xSkTUfSjN9vWtlwp55nj/SzPrXJOhVz7V8zeVAM88siJCcyY8FLVnD
g6QwP/tXXaJ2fU5NKQIt9Z7C+mEwMUhWZEtxXcLSSsmSBt9zpFBVSrjbbvcu5u4vmiilN1+XVyTe
Zgulit2hAQ0c3d9xt1UPp7kx2T+KJW+WcDCCOZLQmszsdG4r/f7r4wdu+NUH7mu9pwTuvzMsKz/u
5Qf2Tlxdx0YR1QmY6BP+V1N7V6EBYvhAZtltzBV5OKEDotthphjEfqNEyTdwwgdJ7LJruSk2Nq4A
JYY5Kye3T/gqiiR63ATyBfisPBh5ua19GBPJUyoYbv381bKk0ZECp3Sinbvu7jmMo2WSrG8p5dCz
ABCNtzQ454LNOsg1p6NoBKfj80Jii6HnnYVVmmCQ4X4ScLUejOaXOm4A4ia7Sl3NXPSLn+lwqkJk
BKYotBPn/Pnk/phprRaTmV4LF06oBbJ/9oZm7+5z8VF+FAO30QbAEb5a7rzdL0SoxwTajqrjSZAm
Jn+tqTSzV3avRDISeXrvK+InWa/oqPk7MYXSzc/4dyiBQYa0qO+SGcVi5WaPYOb73vl80d9f+AL/
5+bFqUjOpdYgYQi7xIIi17K5+5Ga8VkMLrLbmcsOM5R7A7Cqn7unlg6OF+oXs/xMewvjgI4HIu/A
4dWmvRysLigbWsgbRcvBqiXcgIqU694mWa1vVN4Sk0jo7eAu83WIPchzo6mW36KGBUvE38cT/4Qb
hrKpG0WLH4RKDqnArzgnQSub0guOwE2rKkk6eX6LMGGIMG9Rbo6xc9enIElqleP74fz73jpA9SKj
meRHGH1LUGvN9pSC40Kt/xel+vR7LbeRmZfsqzNj4C/8VmW01F6j9RqdseDwVVFEoffLZE1O7WOe
tKdPVL1R/NOGrmOiyghp1YmYTzjauDZuX7+Wzq3HUtwpXBYHPfFmEcz31IzQxX543vxDdrgKbgOo
JygH+RIz6xTVcrztC2XfRhi7NtCTKKZdC48kXmCV79trgaPQUVT1XEbhZi45XPh3iRGCLT1z5hab
MEDSK/1mR9Y0zM0XlW/+N9smLh6qiMxJR7390+OZzWJ93V8NHYL+3hYmWNSwLftleRgm/Of7efY/
+4krwBheP5ktlhN9E9N3dYDt3+umz9NmlKYbWDCp6pEs+TD7IscLVk2yMaqCZqcW5VsQIbLnKlsI
vo37+lmd23yJWzuZmIJ4/UCl7QylrkNA6TqsOXiuLztpGYnNGmVBfy1GSTJkyM6bQ3oRbbssDCGb
owsoOe6pYM0sQ9XzaR2GYUwUIBQZhkxN8Op4+wZFxHpjC+U66w/d4xyrBy5nkDgX9rTLN+4Vm0E0
jbCqVSJANMldU3YctzWg3L9anlBVgmv0SN/5HabNsvyVD8rkNNv/ssaI3gL8cQquWWBo3Q2Zc1EW
XM2d/lt3FOE4sbQbRq7ldiJ/cSsKWiutDlxBFpHwtohWDm5SczdMJvYYAttqIReldb0sr2CsjcqB
KElQFjxrC+nvljbMCzOBOsavShe7UvZugUE/ySDjn6rv32FjG330Iyujga+mhPdC11rdzjH8/swE
6/Z0IzwPmhJJeGuRfCzVoHmLERm2oQumw8lUmcYZchbEFc68z7tsd7JBoI+U3yjeumeR5phCVYnT
QEoMRa9qYyko3/sPuXyyR17AMK0s/b6j80r6zvkX2Ehq1j1o7C8ispcqRGnd6RDvDrDAFf23wdT3
mIsY781keMR87J/PnuJdkYTeLyXqBYy5Y6i9BoVHzuZ+VaEP5dZhYok2F1fE0E/Ri5iWHrl8BC96
FrEqX8/oDd9piMJfiYPtJIlFG43V9cWD2xz3f9MVDNQbqih40wAoKhr7Sz3/YOHX4VxJ2UM58gB1
553tPEKy1I4aygfdDo1j4SRkE/xl9kDJVhuiel2p8Fr30m4XlFtiWZFPrLQvMm9AgAk4xbZE/DRA
RJfjpaxcfsRe+hvvfCVcC+GfVz0BqLsoInIPnYb6FV+JYzyJfku5Tqbryyj8P6tHCkiddG7Xg1uZ
LGDsn8dvJBIngIcrCVi303HRRuRUq0wl8sQSem3T5KcO3Av43Wxlq/MwXkVEs2BF//Q2FdjI3Px9
gkoMIadtAz/VxpYoSVdQb1XbGFn0qkWgUcTYFedS5TPbZNS/zfQ2QiDNaYwXvx9IMbci0TN4918B
xThS6HZHuXOgCIbz3f/fi+O1vyQORyeeBDSAGqC5fcslkC9V3nxhXisQXF2kEJNquV4zhpSXOOPQ
aP/tiMgt6eafuCab300aPBoHFiSfRliYTTg8u8c028eR5rfERXBescJeVR/7Qde+kxm8R/Re47mN
IgUdznIwo+pmbXyyFK6Vi5EhHv3Kla9DZbxZSEhjE2h6QQFZTAYZY8/Pv8MbedkB9uA/w2e2ciCB
ezmPAAFUbHapXXJ5Nj2NXNw0x/p9jkQ0ALVa8fEeRn2GHkT/fbqW+ytl5s7R2vW/kKlmY2rYrTaO
9eC35E1bXwk81XitSK/f+RxbEhG7P6lomg+p1bHcvZ66URMf/tdeszv35+1FrdlJYgnREEbOIV2g
1Jgm/FwKoSBBdS5MVslC+9WDlsyNfuOSwCmeQVLYxdXdm+B7cZ3i4CBOJqT7byAmO3ETIBXdPnHn
mItJuGWfgAAV2eCU7soENwOFns9ygZWmjW0qReXtMzIQ+dvmJ7t81Se4swlRNOZ9a9XR4lWmWCPS
cbaU5ZckuyYDAXv+gr6jim0CtDggHQffl+ukENHIhasRmSb6D1OZNMxHZXDx6H+Vtb+UsMjxDgg8
Izccda2sibieSqwP8FaxvUavJZmpoZE3X1dzgnHgMkYVwxeB00AwNz6nYhoqIdy4fVNwZxaqjPU/
otZOgGTRrt3IrIQuhwpYxms2Xi3gLbsX9MBfyJpiTzfJmXwPtaynptm6r8zfk50oCAHOl2vQXSBj
Wg3iy7ZSe6Py7N6dNrt1LVb6GtvacieDfnllqOiHWn8Lx1WWUqaVhkVTM86Rg7WX0I2FgsfGm2yh
2xU6l+ozBgzuPH3aZV8w0NjmcU+qE6jyjpmO1/FQ9yMaIjj/BB/c5cwWWVV/ua4rwzncJ/aBe/zl
oB69TwhCbW8DBQbPyf+ePkbJ8E0GjBTZSKY4Bs13TYBflb6sRd+kiuUNAO9kZtN0zlXMKygjmPeE
wFH0qsYcWS1uWbOYoYvqUepNzP10R3s/ZCQOTMY55I49owPxd9oa733QZ3Aox/pkpKE9BgC9IFEC
lEur6/v1FtxFJ2ZVpt5QIJY+9a8XVzbDu8pmI9sBbUzYFgUZ8tfzyd8w6ugtr/AWWL0IvDveYN7R
7iy3A0dOckVszMhyH1PZyBSBuD1pA1bcQOYV7TejHmQVcNWH3ds/nPem5jjoBjUa8Aqdt0PRi6yP
NHhe+/JbgTvSpo8uNbJxHV5QWFH9t+druef8z5xqAwrZOpyTot34yX+pidizqMdvJ5TZ+YA6y6e0
sMSYJIBn3OoNFLm2LBTppZvoUl7MNd+rPw5m3lN7E4XCY7MzMZ8TmXYlHVyTMyoMqW3qfGKOsXOj
6OxuD+otur3rQVhJzTNly7hb8PO/9RRCO3QxyFwjZC5NaGRU8Ry0dyN+j39wtlQr7ehBqq0mrFyT
93PvwqzTIR9Mdci1Tc6jBoPH3BMTW9ijXW2wqwEmEpNFTWYzvCkf0+SrYxEkNyS4kDZCZ7B1G+8G
RIYIrr351ZxaGyYcf9wF+cKNK/oe398QI2tmSTVRN6vWyY0Xen4dhVNcp7oDG9Uxco8oC3szuflL
2JF9H7ofSMKX1vxxhNSvotBC71Vqmec2zxLqGZMYqnqi6Fn8rnDR+/bK0KZhaBHxxTxwRhp+SyoY
h0MaXLy3R9FrsFzrGWumXYPOdqFE93jeK3t3EbDPLTdNgE8pnHHCMQy4EnNqbmg6v6h1+CpFd3yV
eQgFEPoZJ4o2PqZVAmy9+5PU0Em7F0CrJLE3s9jfj725i+cdUBl7i8eYZBqL13JSaCAYrqmcexgJ
jbThfG5El6QUL/TCfGbJdguZp084G9pS9BmTQ81i9awJOOGYi8zWZKBUMrz6sED8u5zKQLiZ9PM/
OdHgM716habf+vMKjGa9SeGfDq8zslPwAmd+0o4Rq8JMQjspn7HAdIrSO4qQWffpacFAM7EXZIZe
x53+zqDvPg6cFFK3e/NYzfWcCS6VKGbl5ssjjks/sKdI1HbL8dCt6DBCBQbQm1VsVkih+LZcRZ6S
UoE6F5+SVH++uzXJFiWPNJLkEq2vul3Uv0R0B3Hkq1Z3j9dwyvi2SYX4D9XkaiW4Lkhi9TaoYd/3
l1Te7ES0phWnxyJvPc7iQE/i23Tu55prMwaQyemgYdwOEOrP7h0z6Uzr90oqNsS+ZfV3xpjwY3F1
aRYSs1Cf8FFq2Rb6rmpwlVBq2h8/S+SO29nWhUr/h4q0BRffsHlJ/r5N6Ql0SZAfEW0D1d7PSrDW
+vpr5QwgFVzF68zav26i3xIDjM0yK+Ej9A9CM+Sx8UgPqwYAYu5cBMxs9PwE9oSmLzn0RodeEUBv
MdqEDOsqqd2nIHt8Q+RAuoYGa4x0YHKfNKKBsgjAE7HRlJDIcywzZ+D651c9GNTRp9yPsSB7887Y
Mx8brc04xnNS1yiXFlitfTOFuFawjiU60JGPxjALEeBRZ7xRbbHrYnGOujVkGnDKSRMlnVKFTymZ
8kPSq3vA/28EDWVNW6mouuujVhZLfioicCJwlNsbAAHMjSzjl2UbPeThwFYDu/5bYNcQqzcSvxvA
9nFjOVh18ii+vWe8RRqqIa4NelabynKC+Tpg1a1fKv0kHD9s2+hTn4I7WCDMy7tL1JGyDwFyn0k7
1wj9cQTuf9KnPVlKgQvwxT/x/FhvF9brdaTlLIoYULGZ+UvkMiIDLkaEExHWnSr5QTTI/9NBj+Ac
UpJJi+7YqqX589OrqMEZjnuG7YKK7twwwsg+gfFMyH/yDfQKfOe0zFuOR/O5sGkIXsoi1u1EaNOC
Svaad82IVMBZKou9WnHRkFiBnJyFLLJ6phELGVHvKgujYJ8K4U6ib/24MZEIq8mlUGVYqwA9sMLP
Cifjr0n0G95DEaYm0NAZ1ZYQrr6T5E8xWGBuanOkIkM4K6sy8jP0HcY+VVwX+/IHQjNTM89qsbP5
U3ebe4Sp+LsF8T1RxjhcdYBaXy1xg2VLHsaFLUsRqU54ipazI8ZODE/QblJ6hX//zfOFIf0L97LL
pTdrCDg+rJVKw8b/vUbIl/mevR9rK/ajw8GErXn0lurWbJWOz4X9yU+GAsLoR40DiruUtXrLx2mZ
GM7yUx+cC8ATC01o2HAbR+iYtuFkDSVo9Eo98T1QF5WPm66Oa4c2Any0DyB8tVBdj3MnTvuVnzSq
BcDIcI44bXlsJHQH62ufwdV0UwOe6snojHSO3aTZp5IsnOl0WavTBOcaeKRW5doHpx3an2qilUnE
SvGperyoBlUk1weCdGhc14H4Qasb9eSzrjqw3O45Tt0oWf2lBTV3zAfGw2Y3IlmaAXB9Z4hxTpPF
tn3AA7phAsaY/4VhPa9IXsHdlSHjB70JIZKAS14Xsum0FN+GIFWPZgShhte0kASJnx9XFAl09P50
xawt+Nzg8YpR7PfYFkOk+JLuyE3ewp6+I6m8cchYB9nIh50kXK9SDDuVfRlnsF9SqRobTLfhnCdX
cC6jAneMqKysr0qcI7SO9/6PCFHsNKN5Qc2/Pikjl7mh6Jkbi9TBgPuU5aAd3d4o/4/h+1+C3eJI
E7AHEb+hW23/AIz2hgL3gAqfxqUHGiz2zKPJKpa1R2lHB00saMFWnsEW0dwpECFRFgq7Xp+BTBz7
yZQjbd8Lv/oc02bHcnCqwbO7YuQN396JmP2YJPQJy5vA5/tejE4V9XWOnfpWz47bpoUaXm5jp83D
T30V6Y1ng3T0nK+E80xHpIU4o33GEnSXWlw0ic74yr+vUT3yhV5jR8lUR7LKGYovv/K4T2mSDqP2
LmZpBBT7FdkxlFPFffMKX4z6xGYbdyI0GcXbnzOGIHnMllGmD6+/BJqf0oVShGvGo1GniMHL5Kby
PX697Z8Nr3x/L9c79Xi72kRvWqj8n5G5yyK6vYAB2v0Mi/hqBllZuIWpjuS1zcu+eItfW1ncawZa
MintTZsiidhapN0la6mWa2YPHOC4C1YDlmWvywyVvkyDqQDMZ3vohrHdgN3C+xlGxZG7oD39jLfH
DjcMfSSHzjdUuH+b6sS7TljH4hi5jsxErjpQvNZS96IHlojIW6h7cyEXmK4Byir/rSjuzHmi5lA7
rJE8+Me54tSoYvo86VRKPDlzfQXiofDUU98YQ/9jjFWl20AQtFPN7dx2hDs4svAqqvzTDKcQ4p3T
Fy3kkHFF68poep40lx+53MAF2JryVG0bpN51fAH129Ec3n4BRW4lFs7MgeED80UQRB4KWMfqQG6B
3VKCkFkpRnTk8jEN/lUvIBBlgHa6WY3OWHfV44TkOenghlHV76/ICHfLkFUVvwL+9vef4bWR6zEC
YTvHpMgAsS4qGOYantWfac049iL9FhwcWGKVfUwennzsTsvXeqpppARgOVNFND5svO1qW8GprWl8
sc8Ddkv1kndCKnlmiPMyc9ezWimsmqQxG0KlgALMRO5LdpL/TdiRUzFWLGswNcrjl0ly3zWuQgzH
x5m69F9EAMUParurvUzTB5au8cCRdc+Oj2OSw/fZ0VGhhnmvUEUNmDOuFUhL6go5O9OfF/1i1cII
478B6s7pquPtFuyxnuYvmmYOGRSrC7YP9qlU6N17VyxtCyV03KoNH8hjkWHVWYw60KIiTipDmjHM
ndILr6IpvCFT9GOl8ouM7mvClcVMhIRCs9YBcGDKzu8DB+8CSFj6MojxP10Zv1lPIrA+4XeOhOtt
NGwAS1YPhmR0UVwotfoHUaiOSFCNr4VJbDGepHDQ9D6e0UHz6JCrKfRVHI3URMfIRItNzO2sBcBq
6Z1VOa/JTgbI9vePB6wZ78K9B3bdLlP7b2x4E4vJBRr726ByQp9yFaW27gC7hxoZyv0YGL2hWBqR
E/3of9eJpmMpyZ90xkIxTo0WlKMKgOS4ckY6KFAxVDMagfh2xUQyEv3HfzesmnpI0VnmdLbCw7l9
eRNYiHCV+ALjgxYish6caozl4dc4Sd9qsUphbPTmt2Ed+61j3NRAuZJ6Tz5bhg2UrsmYacsjVn/o
hFxbpFu4jEaSweQaaadReIrMirULOQC9a0yTIRsEK+fb0ltjBmFLwLSZN/swM5eQeh7H47l5XbP+
82yq1EsXFCz3xOdD7jH6t493HSyrfw4MeH2DLRm44qNPzfl9ZVVLipsqf9rDPIqKgd+cFk93UcrC
7/1ucfS/s7fRAtyYWQuWx80sqCmDYzMeQ/vgIzAWa96tCPFoA0hv6IrN80Tcmq3Hdeg4PkfpjGan
M2Mim88YH/+Y2G3XJlx2hCjdwCUTUixBYuFfWlMUVJdvuLqK7gH8RFkbYkqV2vZD0aoNPwe9Leik
y+mck90Z4BrISyTm3CEZjRAwobgSJC54ESpk4G8eutXCwsmf+8Vu8Wf6fEJOQf4pxDSxK7yRrKgX
Uy3ym4iJUeevPet0weyBJe/1yYWHhoQhyFn1AVB8Hn/0ag21O3s1Sxb3htCQyrJCKKouRTQDVxNv
vxOWommzUgQkaEVv0kFVvwF8fD4bEWSb3DUzE+Lx7EDrzIluyDhr+kzgZp9C7OSiWuuFVBieEpd7
XFo0jw/jgbeugoSim69Hp5loxA9Mx/boPtWBIsHFXE37b67dv2ieyCEJnzez5+6hsWvN4jIg6Qs6
3N7B6E0/ZB9nqcxOBmgVWaMN/MC/4CW3WMt/2ZPVsWjGovQW0gTMrYKzbIF6vuvX7CYwkTsJK865
hIkbdhlOBp0rQC2qMno+nFx3foPJdiJWrOA2XcukCXJoKCalM6/BZDWpYXy7PFdbrC7IIVzEZvhG
kQh7SqMJi50XQJhbXVypQKxXYHQeg9X3ruPIFvAmrtVzlR2zxC0zTe1cIvtUY7kQw0Nu2ne4kvfC
6TBvEmbJFKGGDeiAKYA+I9z3xKTrHPj05YTUM9S1Ql0mU/wKRe8rEIuXzn68G81v3VQOmO6vuiMS
hSWV9osZtdTplQ2xpQoYAUXfiVmEBmZshPf59HyRIahX8MhLfcxkc3Uq9xNL/+pFc9yNvyfNGZM+
Sgzjs0HFmW2fc2AzUewdshkk86gr6vwJpSBv4axdB/L+ANQBoDkxDKq181D2iTEOaTOUvNQ9j3A6
1nBoketP+j7tZzP9IIgpibm6NWUzuQBY1aNm20J/aIfCb0HMWEpPI64qVePzuUfG4xLaP/IiKLrY
8kjrFGKpN/uddC7KcK2HnYbhgZ7/Na/EkcURFr5u6Ry2jKdzcwIY8vtDqTJ24xN4vn63meixLTds
NQpUimVuELccAdDLQ3YPBnVcQHODMlx98u/GcYOQewWDdBGIFqwvA+Pv3CkmEc8o4gek8rvkF9TR
PmrL91z2ic+LkDGKJJPg6iqPwXN5u2Bx3npBthRtwOqMRHEOlCt7JYbuDzpK483i9HF2YjvH68mC
lvK8BxFpE92Pn5jW97bG/PP0HAjo7T+1mlA0gu1Pxqi+unAudK9b07I61fiArxowjnVtwX1MtgwP
fEnFw3uYIl6zaCHaaYYld4rlObW49pCqm98zONoZaJunOMfCPHNUhOFNkmg0sTV2iuii6wng52lj
b5UAZUr7nxw3IKitgbl8zdTm2dW4XjfiK3ZwbdtIxrKloHKimSCRFfU+dKzOQzxWt3/ZQJAEE4fV
e94ClVJC+LlQfeGiG/nwVcQTSZEQSCLo0tmTGjuaaV7dsOf8LQatozCMTIg4vA7FN4bc3lGMj2n1
fBDK6/Iw4bQZ89RnEWQzs7qGm4/MuZahPMcRBNAaYUHoEnlQf73dvMrtxjRnKHlvC47KMJlv7fJy
x5asrRLfyU07vc8gFliDri7OZPfa5jxT8QvIOEzs4mQlJMrIsdCSL4/xHW/EDEaljm4KBoNwzSyD
iyeMGlrWJwsiRqrcoPDhJ4XgBKTW8iqiugKKIAGkomP23DWL/c9WQXtdiCE1m5jTIjuOf0lG0aJB
SD0nju8lNOnyH6OX5hItFJpqyC0kbssLwogMb9v2ElVEOfU1w1JXfk/UPKJrQdVotK6ADo3pUT9X
kM/f9OMzAESOxT2ZgWy38OrwmzT4K4ieFnsKBbgHeNnDmoV+g809ro5sh+/2/r+22bOxdEM/6/F7
oPP78qcHGxhyH/GmRvrBHkYbCDMC0osuBCaCkbXrmXpxQzQDdL4Jp4WHluA1Pt97PIFJJqdORFgG
Hinjh6N/wLMYsGeLI8HXIjU5Lp5nc1+1mZBw1uvqdkiyDSzjKvsz0zPuATAojg5hdT/WADxAnIVb
oJU9Swneak9w2nCCA4mawEMsTk8esb/cZ9+pU0JRdm7sBof1ItY5eBOXQyoCCHDovkcT2k0I8kLs
TILgf0MU3c7QLMUN0eve5XtWG8uuZgr19D91sPD/I8wvscijHRy64kANncqqs+hb72kF9s0ZB/W7
pmCMkf/ZYqqSq8Jc2q98KjdYYBuelUIp8KmzeBdAKJ2ey9oZeD8Cej8NPjm9Ok0FUZecQEWpvxde
QCFA5Gx1d7P89Xfnlhq9MK2ED5Rj4uaEygV9VUkNAsmG/e/LJhV/8beuI7MtLulBMGflu49FgnYe
7YPYNmtiHTV/ZRNgRnPQMi1wlvlLtqrokzkkfJ8uq3oyOFCvgWK/BKDwjnm/n7nXjTObwG2sgK39
aDAzx9FXxrGdoPm501KwwypA3UfyPNpl1i8sIpW1aej9i8u+2r9kHYM3MO5x8X0Rh3E4cjDiMgh6
IK8ZdtCiKTRlbZcmSVE/LH+qAc4K7b2pLuKhq/u1TOYNQ/znJ6/ughqZGZ4F5/7fNVSTGtAIn9Do
qVKguzCcKHm2Zw7wD4g2aC/7ZwEGuoiWFuv++uCna/KD/zdCxOjLBUJ/Tuv2CZszdm2gRyBQ0E0h
j6rQl+Wp5oeHM+dVlT2nUrvf/3mGzVxVsGODtzhGDVbVK7fNof9FicKs3JDpmxPdNYYp8RLT7sp9
k02CB0kiBmNvIwYBH7FTYzO7hdETrN65w5wicCDS0o9AfCEnPRI1QHgGhXiVmcyc4wKh0ZndK8F8
Lgzyd+S69L66ygT2LPqgajO//mG4kEJhFFIkqV6XsXLPVKpr3johhSKDHfvk1FAVJuykRIY+9UsG
IxE3vzK5DLs5e/WIQ/7ZC08i6bmGnLRfaO32cXmhODcKVWL9FMcZ+Ib7iJHiz2+UM+92PRmCmmYa
j+Fk5FVJaQeE6X6l/sDHuya8VYvwjkum+pQmD01+xbLNOliR9JFjqvvHBB5npfa9WNBjRgh4pFc6
fcrodBb33H6/GeXac3MrhfsZQ5oB9Xroohj3TKYCP1xph9p67LTieQx1uMMOMN2DEXI6be76A+4L
k6TchmquWni1NCeYzVZSeotuHIwR5JAnWqhTJ1rAV3U/Umc+2SgurwZ4iGA8K06ZJ9Txv/lX1H8z
VMnxk5A90zb7dDVpsh0QQA1B5P8X5ZhZRuoBDiJxZFQFoiNfqFjFAJk6WsqZuPYtISZG62f8zTxw
KDiR4ti0YmxAod/nJhnnhq4rjgG7WUlwxqiYyJ/xb1PQf3kGfuHB5jeQbgWUuUzjjaBC0ufHQ8dm
UBVMkNZIjgiVAc5cd1d8nI8DOqoLc3Of+CVFBvauHVOvscWVUWpwd8TL4u6kEwSd5DeZa22VqzbX
9kCa/mgAa7jJT70N4MuBCRK+AWykJSWd1JlKFXx3cmsW3tCgPg/UoshAno9cktCBWC3kZTXoeK7r
9ORZOe4dfFSOsJvznV8xgrmzHeAFLGLEej5jTEM+AHtxlsbNFfJCgvxC9dqGIM/S3CqiMLMEFMIZ
1LfqHm7KuojqBFIkthFIjCtB7LjLwl0f3TTBHHO/3NobayIfn3+qQevy7M8lgdjoUc6MeR1wBFXy
3ES1yt7g5ISKcM7hsdWenfDXtBWJBrK87ENgjC3IG6BbAG42XP6BugBo4eQQF4xbR3T1hjFOl5d8
DCDSnYe2VsbfkUgxmxjpj7iRwtTlXvGLxj5z+KPQhkiSOLwpwqOjy+tGwhpqlKok6qahV1TjydLw
yJ7gpnLlaxluBIN50l/I2ZbUg9lTF6EFR5hZm0pPwJqCvVYmq+PdTNiOQAOmgTziLHXiSCCq4FrM
QdjwWASCA0TH2YJXWnfP9eTS4vxzaEiocdESBPJpu9DclgA4rWivUC56gbj1EWJ5+IxZEFFUHXHJ
BzJ7O8B3AGC4TEKFkM1I5WGMZLq7/iun7gGE0MsCJi+L2W4WyjUORR2Iwd9Xoc7PNKZH1veA3Azp
c1WlR+FTTT/qW1gxqNFTssdJScwroqbQhfC4AjPG+rs2Oklj4LBqPBLnXUCpQW1YtBzRFKO9nwfA
CvN1ObZtMovko6mANM+/R7D+IVyvrp3qgs9AfHLjiK2dTL64PZ2XnYuQPeXRodDNwrjHd8Rp2/Y1
SY8UOUHsWDq/FgEixqMbR6AwIG/zTXDubOJ2KXeGQUOdxgVijQliYyOHvaFI3JC9ZVWukdIuiQc+
i1T99hqCTjsl+8LgRYOO9OuIlJqUlg8BGym4TK1a2XuO6AU4pMz6TgTXfBWSuD467DPUey4fC/V+
XtUbaXv+o0NvI81skGOF5wOPIvR++sfaMFWOyi9OFljWXrfzMyHguK9YcuxzMojVeObCjB1qTM79
Eyj+Bd7AEbuIUj7aa2h7w5OuHqCCGDqZevRIfIQc++ozORstwJhspREwdgfJc0WrajSuB5O46pj7
CLdrwTj5+B9ih5VT6mRSrucU5hZX0JGzn0V2MDXTetcU7XcmxsLLBHQo02nYuprSzaKVKEWnAJVC
3rgsmFDgyBhK7Dkv8CXfHiUdJuO/OWKcQTRjtaYxezZ0JK08OQP8lD6iOTG00FYNs9AdVniGlG/N
MrxMDvN7VEDag6BwHJn+pUBR++XSNHiFJVHndTaxFlFb+XOe/8h73KgLIQLwFAW7lxjF3x7LbVw2
2XAEYwEqOzmJmhVfTTZjLk2FoQXu8aJSkV76l6Bjd5am1A5xllqG9O1Yl2XUw2gYnUJ4F6PMQbD2
OrxNhXMs//I+qlaW9Fs9pU/G8hopaNeTl0tQsuR4sCgDOt3SS7LC+at0p51Rl3AdeS0xWVFvOn+r
KWkNX6GYLlaOpclw9PEekN1rVcEpdbUvKyHTDHbABuLve6sOfqG29szDAAGX9ypWzauiu+o1vxwO
s28CN/TleTy8P1EnRYYlvHmwvDsth1cukUGZyqYCgefmPeQf911LkJyuA6HTodReGnaUydyddLE3
P3tEglot1gjT/FCD+eKitqX5fpLjskg6nkNafMqDjpeZFsPLmHAAm3IENPqZts36M7ouuioLjPz9
ouKU/d1i6gpUYyI0KH0HZoEJkLK6/GLgiNMG6vUhgOfH8UNHbkD1M/nMK3deeczPWkQedZPalT8S
v+ip8r57SfdyaqJ+KPYcVBSm2ie6xBwd6IwIUbGjFpIXicA4LSOGp3rLAR5RRPItnbqoo0I3K3wx
8XUGXrtkRQ67VXTSa0Jt8BVKMrqMTmk426T2zq0MDWfLuaQiX3RsMEp3qhLNFMxp1fxFa2/zc36B
+APiz0hcduhsbdNIe62/9/32duXjtaZ2vg81J0r7zxgb7LkywOhUZEiSblVRhourQE7IRxAV5YD6
j7qkjxjU3lnwiky0raWnJQr7yAqCoJwutpWhYpSVihJCnTW7ZVHYpIH77crnq5wfig32C3JoC7kX
mf1zO7b4vYIor8r3/x/MJk3pEfZaGGhLWnK0f6WhwswI8qfbHZagZ3TsN7zXOCUGnD50OILaHT3t
HlzU7qFzSzxdhqZZB+ZJyQ1yJ2Y3IA8SKi9m7pXcqjKAnAw2tBvMCT6F9Brgnr7hzF0KNf8BMguD
nyxzNk2WtO2bPfB7Y6LSvL4U1T8MvgBmFd49090Gb3GSu4uNyH2RcSkUdl7WL4hCZeqv669wToDI
qabvRGAjBXXtje5FzSdf4iS7HrMu6aSUq/jEDPej8svLnTiTAzZ+h2UkJsFIHsIjsNiSW0lPH4Qp
mYxPTY+NpDz7u7hacapBuu7szSHCr+jWVGWE2CiWe2X6vNtHbyI+30/ZLJ9NWfiqr8Q8pdNgl/MD
8pXsyZmxx3C+QDJg0OAoqkv6stJU6eI8/FpNzs6BbHN5eauOOTEFz7PMYnC70+lqandbsQ9mSEZN
9r1KTzYTOyDwUj+5IAtei8mZ9/9wrFd4NF2+pypWhFVZa3X6LRm3t6AF4TOhOQeuKK6mdnfQlxCo
XauUKgLBwbOSMj8OcuM9OX3JUH073e1ILAkGnA6zLocK7CblTJY6Pb2Sxyo46UnqAXZlnw7d2xqH
SYSmGciTiUxZJ7BZCdYWm70CW2M7smAp133WiH5Py+dvl3BBsk5FL6yNUetgNthH/6X8Sgi3arnk
kH/NCTuc+x3PkNfpVOpT4H7zJRe6qumBdc/MTumrmTFzJrPhebuTDtpLnWohUTLqfOqPXcBi7HbX
6C9idVKWiCjSKyfkP2gjOoG/SCDmvSELklGHB+L6C9yFA7WJ/crTDjmhWVVGjFOOseDE16Cnn/iI
i+Stk1CFycDiQ4IrDS27ktvk4uUK6kWAESqW7M2ZmM23TrgWYSbiwpLW9MTQVmL7JVIRT/CuBtpx
uFK1f7F1TzAyDMCe58gO86pSWS9nN8wCYWsSPOMtHCiC+oAdDekSrMS3jBXZuVByFXf31AjN0To5
EidGr23RvDLK58Wi60fOSwL/eF1FzSWcZjeD6uAqBWnA+C/Ujrzvq8rmbl0p2hE2neNBhKjS+46q
9PMoLRpmpQMDRBeDCLbU7tlYzrmdPLtG16Wc5xUi6o+sL+fADbnHMSUn95b3rJImUffTQxscCu3H
DWM+PzgH/nh1m71wYN7XKLhDBXeA4srzmN5nuTsbnUAV5pedwSpjkODNm/YAan/POGzSKcCNojI1
D1N/qWYmVpspOyD14XNraOiYM+irKVErSL3R9m7Dv5EfiyQfJbd7CFnFNVt28fEjBLOhVNB2/mpf
bYoyDueFSVJBiEGsofrnLgqkxiI4RAA+z9jPq9cbQ7RNnLwi6vSP1YnhQ37NfvtgA9ZIilcp+Bq7
YcL8w24nmRX+edQgWE0/HS58u7HSaFMBXJRsX5DKorry1WxjQ11zieJDJ7KEqsConelf9RM8UDPI
t/p9esYSbcRSB+rGyv26qEHv1/Mx8o1fEoQCIqTk/eFH7Gg3MAxmY9Lm4MfNXufpVSBj/L7wDDpU
gX+y6Dbcecg0wiiHzudjyOKsyKzctXxGuk3Le5VcXhgIT5lpxkkTGhSRb6IhtQLoUwhn65L/0M+Z
3yR4EVR2w8uR+9U/i3tHHacSgHRZkYJxOwgOUgTgtaC6Wr6ifZ5TwjkZk4+/F3A6NiQKtG1OMHmq
2WtX7FEh+mThJGHpU7KPGXwpuehNa792sSqJ9bB2miriU19cgzgUpO8+fFJmBSwd2X/Cge3HBaOV
H0WcZBZHiYmseIkMC2UGAgCvS8DyYFUrioqVW5m2UcQgL77e09uaw8dKRoyHHuTHImU9O3OXu+lJ
UTMU/twkAcs54SYIiVlfqruR/1oo0f8cD4hPOYmRotwx+BV7O5uQH88ZXno7v7upLDrCxj3mUTk0
HPFpw7A50fk4m+UdRyPfLFrSyvv7XfQ0SWd977iT9AFviTbu3dwta9PR0T6uGr8sTNZyFJhLPVio
vX2zuFwxGS5IyVSFFP9EfubON46m+YvY86whQp8WkpKZN31RVwSyNAcuIn0G8U6VcRNC7dK1Rj8i
bFdNNLDP5g9iX7rixFUPee4qer9nncVMdgPcXux73ZQlWvhL8DRTpuezplvKGbaOiyTR9GRkl7IP
QwjGlK47f1ORc9v+yupjyYOdLnPkSQynAOIwfrrELF8+zujkvycZeMLXnCDkkdD2MdbhIWfFr6/b
/RMfIDT5d0diksRE0Fh4PyRJgBT1qOwsK0zzIgN9hvN5FrXfSQsYzo3bLoR5gcaGR+EZBUwL0VB7
pBVkmyH5zfiDrvrH75/4EbbW/kq9ZaOApqO2k5n4w0gF3dglc6gtvXKusUyb45q7/VTYzm/geN96
lPXjMRqnahiCEtLOiG0Y5uT+pV4hpYVRPJ0hp/VaPFx7TVWUoUrPy5tCrYrunh7J1VAet3D8D5sG
bhMSepAuPGxdd1G58i0lLEgOkVHr0uCGxuWghcvRvLR/Yobd61eNVZdhNbq19T9PzQ6Fj9G/f6MH
Pfesm2YQdc68krVwJGH9VuEhmF0f6KOETK/gHsV7g2zWmJXIZVxsXoCvP1VSJfnA8OwJv6r2Hnox
HaPciAxuL886uF2qSUvImKgZ6K3PZ9BtH1dC5tyKY6p0hawR1IDpSc+t5YiKtTlQH1XbMl+Vss0g
BXRf81q4eMCh+VgGhsnvsRbPiIXUHXTFkaSqoxkuSEcsKVubH8CdxqPJ4b11qUWO/1NGnv7WdZoG
S/TEPrxdFCMvEHKPNCdNi5kp2Hk+G0obNpuPzr3+ANZupJa+P9MyDIqehsGHUCJUWFC+jy9UO2y/
FA/+C7wIv3yNFmGXBaIsHf3eWyXgquJCLU9pyAOpj7wzcBPHJMpA7OTJ35YgJj9QsIugfmwUXWW9
QDLOPGkXmp75jzgCqchTJN2CtASphFJ6GGFEkD1brmJ9fYQx8uWF6DE+cCEEHvlL1z/JYSLhDGA2
ecGJ2RYF9EM8a4DdT0ApgkjTI8/tUsqKGZbtz8c5+XY0ihkyB12JBtVIszx9WKgO7yBAGU2e2qDE
OCXxwUyHa7nQ8LDvtgiIRwRBdFTnFKwK4JQImlynz5LHvEurWaBtVSY27F2rLLkkuwOPG22mPTpJ
KEvTYPPt9nGxPIEVofDCzke1XgiRnMpeuOYyHJegtvWIDxtjomFcx/bRXlkOAPIPFe/Ds/wh8kXt
rt0/7VlUIVrkyKRFTYs8ehbBtDBA+jKjxmKMphk1gck3CZ628EpIJ+o7lnG60KtBlfFrk1m0tdFq
6ck6BT513xy86ZKG8yZ9oMxqOMZ5oaqHIznbKll+53kSFcW7XcDjNrSKb/x/NkH6+uwYFS5qT6LI
o8HCZ2Sn4zm4VV/xlqcbfMMi/6huOi3wcADIC/I85MyoRiEvpMKAKp8VSEId0r8fFvqYnCqLYcUT
9rxMoctjE/j3cfuP8gQ1uXLItryjVpYWQphgaHqLwxvu9ZH+SHStcgmDzqxvh5f0cji6DypqaCFD
+VRrAtCOo6j+kwzZkZ8dyhDR1NDJJF4LXoZUXWh3+4VKOkyIrF/x+D8znSFpSC44QyxoA1D6J67c
hndfiB6y29JRKUtfPl88JdHHLYA5G0HfwI8dTrpPytW3FuuwCCWyw/6pzvG3P3uOYtfLkqw3aw5O
IXoQs7JuPXJw3T90eCcBYx9tXbKes7Voz7EcRt0rxiBOJzE/TiVtfkmah5VFsOGfc8jmPMvs5C3J
SUNPEFXpLGhEBRjXBJ29AX1EIqUXC2uo3Pz2MZ6TByqCZDfP28PHdoCKzprnNofD25Wlptr9Ea7D
a/6Omd1ehiGor+PFva2Jdt/qWSWsAweWNYiP6Eo7JuENUU6LwUv0zYfX0F1q+BoRT6G50SVbq41+
ykL8iG7TjYRSXk5xkPRz+Vyv1rqN5NaTD4wg7TYJhc4FUVkPsdWSNvRCeCtuF+8oHuaUOVbQLQyY
lTRfOmveJNUguK8gxsnhpb194LvNmEuln+fvVywONTmYgcPOTo328ChkkWhpSkRP+bYGIpQJQEzX
5pZaOQq34a1j2mlQvSNeQAovN9b99AzkwCP9PsDx4ut5jP8HyvUwRU9lWyLp5Tr3ybQNyqHFoKX9
DN/OOGXP1ncWalBJEDdAr28w+QV+fmqNu0xolSc16YTfWyDHWSVshHSSaOnQyb85IxT4OqpGn1Jj
T2zomNMJ923ziGMfYGMGYiekm1j085I5ZZAdghxBkS457cmwHowz3e/ha/RaryP91Tbea0fx5D5/
1Qpcl42QHgrZLmgvYyJjNNRccMocHMWCfzbk6fBp+CSSoQsMPCk1jwpFbso+XW0y1fyCOq07Frgo
kD/1sObx92vdyD9vMD8AxoDSVa5Do4495EKhzleu56FhLqX0Zffd2FkuGZx6GNxgr+uHvmimPicF
jZv3ZSZDstgqRnUlvkFu13FNWdmHn8lM0KEwDcmai+ItNZdIjHDgE2lbsGFg+dVVzF2Rarfc/y/r
2xgiWuW/tySQHqVBPDOZlrAMquUqv/mLwehiA6YpHc/hzzUuEQWzPXIHyl/xU7Vbq8SdJn9K+mYl
H/RMXRJKVFQFY6pEnqvH80bSS5IHVjmQsazWjQVK2hRaXbdKp2kfqhq4nmiMQs38tx8ZsFgjpfcB
PdrfDeQtzUv2q5kO4e3gyR012/5PuOPElU9hec2CH0uAhFgnGSaqoOBC2BsdcI/jAzHhM+bRV0d0
cAC/0x56Uwsf6dZoHkFFJlIyBqgQS988qfF8JXxOY8Kg6VSTqYe1kYZ12QTASCYYUtFXuQLI5Tj9
vlCX+1nDMB8JYGKP54SdUKP2Uh/rm0gU1Pp0NZN8ZFj1Wb5emon6kDrJjpqJhY+IgVLd7ivRLtl6
w62GISInz9sYDi8+CaTsFUZqCDI5uSv5gWAk8M6XNxEXlOqVy0BPVwqDafkf9vdbHY7NezP5gOHx
1yXV9Gw42ZqXUKlu0ePHR0lb2MZHB8ZmxTWb5nEMPmhac7u1VF3+Jf4KZmpjIpqB93WsURvmFa+w
kctQtLji2SNOXmaOU2RIhjIoVthIL2JcsDni8GVMHYcXV3RTMC+5r3NsAkNtNsrrZ0wTUZNieRWC
ux0zd9+fSUiYwIywU4+67nVFP5VpizOgstEJH1T5Z/gxflvzKo2No6r+eNjIJWCoheC1DHEEt+IR
0iD+1fMS2pMA34QPHQFsGXVo/5euWzrkITD7E9rTYPglHGzUy0oLEHsWyPxAKKWGlzUKLlZmwMyu
CffWvnBb6Ws0MxOR7HR9NQIhDXxqy2MKbHLMMoUdoMy/nHNyzKZfO+ORnEs5ux4dPXDdtzmoMC3G
eZaE+wehT7sx8r9DMzumV1xnx3OtXoCyGAHpE7YFXPWFZxcs9tyTnsXSFIEobErFQ5yyeVMS2GzQ
1bHnmWc0U3Z/a+/gVLtxEKcfkuAns6zWfo2atqollBVWQCRv/zBf/KZgXaNYbHKHPBgg0CFWxzfr
cl3GbIPFswIRC7KEq3eMFfAqxAEELgfo97w8VkFOumk4e7EVIEKaXwLJdEjpJGfeEOpUcJpSzuqD
NY9ECBsu71cBjO3HhuMOopeaCGE9svPI+Jpr1u4FrZqLK96oYxCy7WFT9IGe4emhgx5Q6avSeOAK
qJcHzEdPhxfX+Hvuu6Z7Dt18yuUb/9NZDudaj3rIJSn6NHvsi2p6WhDrfKtdAppx6LoAqA9XUU3y
15VPfkBCrbAoCTGcMatuj3+boaMRlv99ASES5w/2hHtuxOzBWnoOcqH79FGRwFBcdNeOtzJaB5ad
sjjXXQAxSQAhO329XjLWwZfSTzGwLt4+YO7mJ9xDRTbLjWG/MJIKDMHLsBL/Ec8Ls9IeTSE0EyZ2
LoN2zpvu7KGoZKPcnNI2hMhX6e0lrHdjxfxLjCwzzl5koZ7dak8K+eMdiogtMs0UYa8o5y+FLhb+
Vpc1LKp4S7N6u4mWz4NsBA5jceeJSgooxUrM/gQUtCDeqzjDb5e/sMK36coAD4JF5MmRYQ/x+pQ8
l1fv2qU4PlV1dxGkpQtAjp3vJQYMAlwVxe9Jotd7dtdZJmSqhHQzQCV+0FvgMd60dy87tE7p2b3F
ZJ0KGSGsVPbMQiAkfm8DWUsFrTVU9A3uZHTIJgZChrwkgA6MFOIyEnAg1csekDhtVj+Ec14lJxQA
xiBq+7DMOwDW+nY18Zm1Ve37SyHVpqu+yIshcBnJBdViPshr5MoYqG/M0okLziMqkQaXwzVXapaN
Pm+hF2H7UB/CXi7nICo/MtU6xxNMpAojlpZz3I5G5f+1P+xXi/v3okQYOSBYaq8L1PDzBWiMg/yx
VdPv43qNWVwBq17KmSVp2DJpwsKydI4yzaP6FWQ6qv/W1fr8TAA7YlwU9UrMmEvcytrZEMZt/rex
7QkC6qlDj2od+aIQYMFkVhGNcKTcmsRHPdhiOLpuwCZqtscbqsyQdzVlbkiujRUs9Nge3DTm33ta
tIBDgjuOMaIEx2hRPX1mvE9LiNDOJUuVTvzL4010Fft/4QZT7z16lclL7d0GVomonfhriJ8ioZWC
QiiUjuMcGdcP7NtW8OVMbvkM/L05liXS02CGCJUGLTrJKWN3nUtyqKQ8YX4Pfktl5lRWnVOFAatV
TCjedy4lUSgneJzJuzeKWzC4EoPKXur39l7hchowJYjBFGiixx/TxSZqzkYiZhoovVB7SoT2lz8q
zPAqZRPCBb826n1rnurxmUReyMmTx/+C41Mari0Ky7a6ollr2kDIY8rTNP5v44c/7FB6SLKAjUgq
XiGVUui2t/lqydIHhyMKR/M75FjmUT9T/G5qFK1DaJC1QHStd7RNpq2fATTxzEvASMCyEQ0+DDs1
Jm6wjid155XTv0uVnBQEDJDi259pco4iSDAy8hs3R+ycQ7jmEq170ZNKRS1+BI14mg0qyGB4V8KS
myyhdfej7EFGW5iUmG/FpD96b0+Jf12TiG1LcKCtKRI4uofxTfmONVxChI1rsUBHwEuJqVYomxR7
yUiJMDydD7O224FWHeJhjMNojrPy0CKAABFL7rp/t3dQlPj+9vd/4nCs9fMj9nL6UIsAIzsVb4oR
fF8zRkbkx8maF86DiNyqvlNZBmLh72egk1XOr03I3GMggIPlf8pj1Mxn2aOkAe1EKuoZbormcGEb
ZeCAgDjjXdO9WxKww7ymKpWq+3VeUFhBq4y7ApOln/026P307BowhfEe0349dZDQ/QVj/3JgGpkB
vZWrZGZIcnCgAyqhF54i9vTIzhVHmyDDkpAL5aJXkot5kKfRkZsj2N6HoKQY92jNNyQUfUb7xKPC
bysOK14aqrdNvJw1EFbzFho9Phf6QRLdnakXI6vfZFTxRKRswH89gvaG+jKrulYALtS1qWbVPA1/
n/HBiUOCYcHMRq1B5P8HlB9UPvvGuTcWFRfOAAQGE2iPQysvaCQZ3HkQEetwzkI/w+3zIeuOjhhQ
33FGMFYImBHiWESUiDGYFfUYYFy0rFzNwuDWmyB70LwYV8W+kHO8KxePYV5rlwK9KSa6wH00hkJt
xUjsd7CoXQ9WTrfHU4uHLLEnVnM/AJVlDmJWWGZm+RaLBxEyCegpIQoqpAvlGOXb4R0edrICwG/6
9l+nq2sYb+4oFtODwuhKWRADVl1rxPt03vlRuRF1FmrQXyG3A3ypSJITJ9niM0cYiTBMdBZxTdEQ
980HRa3XKyPK7liLoEJNWK9LnmXe+HWU4+jVbK0lmNkdbQ0dTsm/n7RTI9g9Mv8M9pZuphc2PoGx
4FZPpo4ZwgPYedz+97DPUSGB3QvaI2agYpTFskHmo2MpszOywhfxjwwT/AEH0hBAOM7mfvhNVT2p
ZiZmWrqPYZIND/LuJ3d/lCsHrdb1fXCT4LqC0lXqmyLWmoC6QspwXwSYw4adFvBU5jDkKMCd4gIH
cT6d4anNHJNG+kEpqmfgOb918H/72DmJyXjQ2wENm0b5lUNvCCQIiBHhI+5d7mu1rEI906ZXTfpL
QNTVV4aOUda7pcWB6reb993xAsyb4AcdYGIC6zTE1NUFI2EbHtjE2Px2PHPVhmTsMw+gIDFx3EB1
faYU0RDnAfKQlyDawiwIsCLZQ8QCb928ZReBdYOsQQ4sYugJ55yNw2OyGtmUnLW+Yac/fWbGg2u8
5TVtOnRTZhJ5XvR0xqPoXkmrYhXFFguukSVUJIrcdRucgDsFYlMEMcKowqUwXwZsKW82SxkhW/n+
CKOzHCULIFnpT+jxhZaRyEdTEnaieuDJJDv61QUf0732x2uMd7BxKVJru/Tgt0h1ji9+TDbcNVvh
RAoIbOP7V0CFEc/21HcweEqdrfuNnG62kClLNQjtj1SvIsM9tyAD/vB0NeZx7Nw3pDsliXOqrcCx
OErHTtJWJiXorcAK2A27lWfurwZMODtxhG6bwKQMsm7zQ/SvNGlnXPV1jbW/z8MmVc3fhDJyn9YK
N8w5SBHJkqGzih2a+ON84BYKgFv8RR+FwJ4j0xflHbPRBK/UYONaPkpiHmI9VPppaeEdVe0PsnEh
H0Om6+aCQQT0P5P9Ago04fg+TE8BeS3oKMHH4bU0mMHEUGQJZ092XvEBH7nCQ5w+xYF+oCmCOEBr
Cuy5q16AkYVCvbTNKBk13KJQJ1BHyVGYTuWAr1/91GyO901EkEWVyB3u/Fvs8lJnMHT/8fAZA80p
pGxnnVfYtts/MxHer42KHit9R/CB6FwBEyLNudxPVD3jqUcTpwAiAgHjpAkCX4LISKJYUmPT+p1b
NERtLlkkGNBsCHj5oLv9KNXWdV21r3Ne/CHKJjMA3+d44ivg89XJtZuU/d7LlBl7iCz592uIdGVw
uphy6jmmtiKTtKTtrBydkQle5CP2iNQJA7fTlq/0Ky1jW1E/TfWANAXXMb2V1hwYXwA3SDhz3UTg
gdc2NI7COsrONkAsmIoush4XULnjzZ8J+u7sZyWTdwFU0asUgp0n9dc99lUMpYva3ANI5cupag3J
k2LkCCvsOLchmlC52vWEvMSdYDPb4cX1eLlHzSIK2vpL7i4LzqlWzakPxHmPxuNDg5uTVTrxTdtP
PqmXv+2mW8DRumevheeKX5ZE+4Jwz8d5CHSfDl5xlY41zOP5ZcEICyv+23/Sx3wBoHYMmPd/NMTS
WjMbUDUTE/FLaaIGvqTEOSbSjU5/+9J+7RNucxi41Rq7ZN575jWxyvdhrIGb7kUgvc1VbmFUK7fm
V+J5p6E0pHHw/MIaaTDwETtjRock8a/agmsfLJihJYLUEigDtuyuF0xfTr9g+DZt8HSWw9T8qsfe
T/Syi5rFyRIVgAKA8+YE41+No7Vs3VcDu/ji8Sj9rrjQhLsSCffFz7xqd4KLXLaElWEwL//7Ig14
W8jBzgfzhEE6X4mYChLamX2f4w15YSG5UB0sMwdvdh7KH75NRf+kWLnWKCLZ64BecW2+Yu+KjU5K
1F+kfygo04UYfc1FP5wSwdFpWN58E+bIESw7GSUUvRhgnJ23BXzd0wHj0qnWVemSj//S9aPqfF+J
q6DXiah59qftcG4xE0QZ330hlyAIAxbsO4HnHFXEoT47g8bJGBKvsFSnEVcQ0OuUvI4SGllmDYi6
gEW4Cswn0YvRrwX152oeLDWyiZ8ECh6Ntcu0+HYUf34p9ueCuJhd8ZC6+ZcNR4t1JZE0ugWPCTyO
5KKxtmxVt1l5tOw9feoKCTLiYyzykUFBIRqflwkPkuOtqO7L8Npc+RH81m8K6VfBx8bFm7wfs6QN
97tYm0rVtbEJTPD96DghyA1+pDPboJkGYkdyEFxx4apjPbHtmuG83B8EHKR/EgEvqnNmh9rQFrFh
9JmIbMN3FhqqDFpIyQTCVI9F7rB8IFhEKM6gxRgirJ6YEp6r9bZIqrb7+fj2j5xfpb4iXRusj099
pnoviMltqCcbIUZSq7rvV64z85sHaRaEH77qL1iEtRvykGllPauJ21R2NdcnWgqqLP4zn4sURkhi
NC1DBOmMbsxfZUxDcu9RbOLNl1QvYMBm9EGQR5Oun6JGRx/kByMQSsJdOXdCVoXvLQjJAfuqNtJB
sc7nZFMOghG8TXawdl9qPbsQwvhvFf8lhzbf3JpiPjY/ITEdJz3AxIt6h1LUmQmlJYyW1JpW8svX
jY8pMdYM19OwASp+dLFXLuBruLb3UP7d5ghnCZiQ+GyvFfn2oPhfyMo9dusdD0o9b8vQndJd2J8e
B76ERPtpjrjHnXSTm7xEkdqXKv2PnKOFcFmsGyCHfgn4RIpzIu16vr4fp1VwIZuPZIS1/rdKnQ/6
DJc1lykKj61gvacmRMS9WAlKvEIME+LhWiiDQ1nMVLHV8AFpGRMQ15I2R6dN6KFyRt2gL5nLvTbU
EXrh5u/8pa45chXZq+oOwy8GVVjfK+pN2ivE/LIqD6R9qf9ilxba9T7nPffNAIzk1PYcgU157y4y
JLfneWUy3zlOH3W8ffeDqsEjeUG4R9z4Q+u0SNiWMNhXEfqwo6sXgL8Cj4NcM9Lj+O9Y43NopvY2
0z6d9w2Ms2h5U5E+x8nsw8Y/PeDChphhb1FpAbc/z7ZQ0S26igOXv0aUhoiXkuOvYMbRmKiPIhkZ
efunv/uPo0XSiraQJJZQg7R4lzIKVj8897MRc+ZgY17DaUtbh4ekUbBsqkpiz3LEuwph0Ko4VYNr
mko286nPGSkO3F95KsqVyUyX+CBpOh+CkOKhfpi9OBt68xwAhgqlgttYFAIoF4drcn8MjExOOV7+
KaDlKOU80I4pfb16uKjr/ubc0C6Hg8rsFe0JcgelW8TOODfjSl59TrcEO7EqjskUL/pg2CXEOBs/
adSP6QMGwHhPck0h6sYZRSqZ8w4He3dRQ2JzKujxcXcteoUR77Mxm4fcZ7AP70vKpErm5Z1dpbFf
lv5N5m242W+rxtccbUEPO6qLxi/Wca98vJzceNJzpIVtZ3xKV2RJHopb5O8+HCfU0qsfaQBiacNP
eWhSTZWRFKo1TBz9vegL1pjn7MPTFUm3fXlkjkrExdweqhcQUGzl4wRcniC1AWG8E4U92V/qo8g5
/qDv0XbDkGHpBzGpFHHBwub5vK+k9PLDF9qTszrq5hkrIXy+c5xU+O78qeaYO9+Ryw7fQPiAUrP1
ecDy+LyUjACx2wQVflw9IEcEG7fiSCynUv8qDry1phKA3O0HAp/cMbUmY9x4t4H/vjhTqlahj4cg
VCr67dzkbNDfg3zR7436xSGTqUaWALlkrbAgAftcfN/NTxQfXGZl2y9CzKLLZ6uVEMRYOuDG4MaY
B6fv7RmDCLLaYo3rVqMt43hnJr2oQ5jhQjlkPOYvAAAvhHYD9x5gEPXgwUcF+byXhLIQwPYT8hnH
gBSmm2ikUEb4XG8/R76AJjIdqpCowstxPAA4KCkIG/iSXXKZjUrVxkTC8R+9RN4QLtxLIUnUuao3
6+x/bN/XC2HZdil2/Jn2nbM5wuaKtApIwZA3bzuJjpv6zHwtBwx78ngUhMrWfIbi6UZ3D+HVZvqa
Ec+Tx3AtRYkEYA4aDswOGgqj3U8+I8kF0r+06vYIteqtfjlm6uT94qwQy1SboGqPGUpUBINekIqy
+RW0t17f8eu2qD15GYZQLPWLxeOCUMY80CROmr9do5teaQsZpFLJ+DQHOy+VB7mvTbq3GE3s/S9H
fzKcCjtS18UHs3iuHoS54rXNPfcSRdT/QUzTe2K3fyjpgQDmxkpRMHQtZZ+Qix5v2+tWNbPEK7kT
Zu1dQnKE/eQRdvJ7h7lQhG18EhN9v8UjSN6ILV59lwmAXgnkm4JIaKyJ6udmzlLESZSvogL57Qe5
W36OxNpqqFfc9PYxL4Y7AUVmBG+4QAzAJAvinGJR6d4eVGiSjRWEAXoOgPjGh7O3F7saGQLUiz0I
11wVua9TV/sJvrZ+KsnlN3Yf6RaXPkOta85VI8Bf2clAa71oAdjVQdm1lCAV6iHhr7KWXaQlivYz
9J/rO+QhR4dGj/e6RkfsFuFLP/dbCIERZ11ZS7stB4sl8mZitwE1EIWKrKHqyeZ3aciNAhAYekzM
AgNHqgqoXcVafxj7qVozatgy/ofY05trtM1vXi4OIpwRiKEAWwazxAgfqnWrOv96BrkhVR7XyUJn
tFUbNd3pXCc03bAE84YWgNY7MDkgrrI2hzfVNPaGf24ZshI9DQCNGi7RMyn5S10Su76o8fgT16iN
UDNBlWIPNJOLYpfkbGITsdmP5nSdA0WBasQEI4tt1PSX530kLq4mR2n4/wzi30r+8VlhFx4bFE3t
ILE3buuxOqqW1JexZlJKLkzCiclSULOVKyJ84v9Xrt4ecbM2BIxZvehg+saOneboQ7v8P7Qnxn9+
nIFgybxG5bbfSMWk/vgS72WUzgDKuE2WO8Aa65sZLuVtoKURmAFHqXC01lEGO1QYXFw34O/UhCmp
J3dgyQyhL1tCd4a2lBg51aMKKA1/J3d4moVzyJANWe4idso+yrH8uaXnX0WQTaz11P0So7D6SF02
bdzGC9kCsa4XJOR5ukiiD/fb6AvCHZXRDWQWi8HAs26PKpYg6PmvYuCEOW2y54v76QnuU1FMAoMP
4d9PYNuFqadJ92D+TIDqC8yc5uCZ7hHWXjZLW+E1Gx0ph+OTnLv3aVR5YJs7VwhP09hdzpqiBvO2
63u8yPREk3YMGoGOtI6j7WKTcV6OAfts63i2FLdjoPMlp+8SC7UxLsu236SoG/Pw4whW71iPIkz9
amrZZeWy1DJSD2XWSucxsUzwH1zGja8+wlpNSBbonvI8T1xI0NDi03aJ/EvmV9BG4y0jAm28M8xR
66BrMsHn1K6HdyXeKz9efG7FFs8WllgnbkMSuZRY+u3ZK1VXhjEmpKnbSnImVQHm7iHEh6zb7NLA
MYJngvm+OGoFvZrdyMRvN7/n4Fo+szT06laaEaTApKW4Ds9HXk+eIJZh06Wl+QhnjBZ5vhrDQTuo
fC9/PQY3zfBtBaN7cqHVIIfxIJSUN89Ny33TmYdpRE6X5zyR3PXF/4ZZJnQfhE3LXLK7wwriw/aa
7S5woaSTSXyXAl70lrP88C7V9ag4ip4PtS2kMZo1ZBuk3Oy4yI9C/L2LgOUiZh5+7RXrKA9NkREs
3EreBNjL5lO69TwYuAoJ3WEy/1cv4uVVgzljRNcaFhvWTgyXuJCiBx54Fc193fI7wz8+WJPXh/Te
m0gIKIJggy70mGATs9cHoRcrCyfMKWfKAGfJPNADz4WGiBK/VkrEigOBdIH6p+7EXYa3nHEG5oG8
aL1TA+iDfIsPuXX4EoF60jJ7hcSCx9w6ldW2b+8icqAKCp/lGc+x6oaBEBNuxgaHfzLpKeqy41LC
yRS5OQhITgltnK4kd1UxcKAOHsY0/+0ao3CPjeFTZ/zKT+zffPkBNjtxa2aO4fRwap+SW1YIkQWO
f4pJbLcGepVemXFe8Mi9+QBDoJTYnayR4Cuc5lUv2DWmMn7NXvkW3wL0WY4WXhhAUGrEbnOVe0Qf
/DPeIlKpjSRVKB6pSItVoAnsOYwHU0Mbu58eYEkr96/fhFW9f1HAglD3Vuoa7i2/FH6Faz4vkfM8
iKFlSJndKX/HWYF45e/vBDd9xfQKb24wVZcml6rzMNX830KtNOo98x5dOZUG6InE7PgZAGPy8QMo
5Jg4drA5xWSJ2/shjZMWW2AMmgk4X7eBHUY1kV3Abh0Y7Q9+vWDXDo5Wxn8n74EIEptp92eYbnIb
wDMrVlPUCHjk/Gl29TEv7NizJfFRGOmExojQ4M6auk1bndS8MflAfSAMT5obSSj8x44jMnyXpxb+
seZJAwICzZKqBYk2PEZTLHmebAwaqcFqCXfkyvYEQ1s7G6coel0w+4uYuLX2/6fUXuR/Ewn15k/6
2XZXe0aSJb6kAi4cUoitW1TBzSu/8JNh/esJWwjXf5royTqb+7gq6XRuK29w2K6hPVZ8izXOVUxW
sxoAQZ1Bkeqgp//ZtpWJFuLtuMifzl0+HRG1EksSdJvMJNd3ff6/XQrxJQTkfjBQfmHcn+7gXNBj
nk9CbPhrdg+w93+Svy72MgwqObDN1DZxGH2Rju43vW+JWABrbX2fnGMwLPgpx5Z7akvm7yA+nmI3
k0koXhgBSDMfEGqsOLbWo4XIa8k6gEUC3s1x/JfnsKxSgl4qWP5IvdHrUsw5tvcue1ZE/sTokPog
iG3GIeewSGd+1q+lZnYAqoL+7c3jQ6ciZcClYlog1bsChawrPgaplfpjdTmV1lXVbVvJED8gQ0dI
fyKDtUQXRsg3Lz3ZMlbBArULyEkvbarYR+H6y0RtK1BT0fctmanN7hLFM1AQxyZbjhSTef9xZdfZ
f32E12qDJxam+QkvO4cAUPrBUoorBa/QEqEonXimgxqAlbGeqVyUyqRqPMRqcTXSC2x9PVMaZWsV
GcA2ghxdcF3wche4TBFcHkc+2M0soG+0PD1fZVJPiZiqIhTsuS4Jm8MOwajn1jkYVNqOP0bK+hk0
+2wW6zTBCaUkym4Rc6mc5yHzy7hNI5AxYHIpFWVcj9yQCv/F/zEA6ZGZZ5RRxtok7vZRUQOSJZoU
brPlMU6JI/EyRzAiDhqGgrh+Uj5OZglz1sB8otbs/w9JQb6yh5NvdSWHurI8Rr5r7x9orMrO2BgN
TYYmwX2sULMAe04yNqPRpcRySnSd5Cn3GoRQ5yXHXuhBfCGyLUVhzqj1QtkNwETlKKPyA350lMPD
AeUI9Q7AXmjMzBwkPQfgMXu4KYUQlbw59i95V59zORDWoHIYVXLFADynPWLYJyUy5H17bHgPwa1Z
+snsJf24xu5gnWMrGk4QNxgP/civVybT+gToIJevGtlahLr3oozJbskxxFn5j3AwRHVlomMfO7mb
xvOCPQy3BS0bRqfY3Pae2qiUWOGcsGEpC+8n8CLQEmOhg4FPQl1oD6q/mhRIaVPUQdMKScDxlzF6
YMGDhlGjNW6zFbrjk6iqQf/6wSaG5IMWK6ySC1lJV5k/b7gDJW6DPAg4o/vJFxvLF9OIUEFW4dLN
OV17NUl5RqTwI5aKY6zTdPc63YUUDDLYXS6wMkC8XqYuBHw1p0SmGc5YgJfS9p2cRcAJq6Pp7ur7
RZ6ThJbffTn+mPQ4w+U8GEAxnmM40SGOkHi3eabkiZEYBvVy7tcSzc7TZs8MTIQag3eiB3UGlBB7
jyxapYoCqFYTuuE9d6Kl/YnTsD2uLo5bC3TMulReZ8/P1+acIO6TyideTXPnWrNF+hgH3wFzjqJS
xFNypjIP34KBO00Xdt7daWyJWJzmyjXrVM/VGefvk1m75y5KCNBWP1ycJE3Qpo51qqUv5P+gSSmR
Hha/EKqQiaCxl2Ovl7E1DiWbgwXyDmR7b8y7Fm2AmULpIrUwgDdWMRr1yxLE7OlEX6mWpp6i8axT
DGg6xUEXZbLPqtwWsfzT+QMZKJKaB0dX9i0uIhrHE9t/he4b1SqqihS65k3ELpgKJP8/6ma2iZkw
AbVFnv7tzdho79Xz5LKtDFUwBXzuzphahVKrKFDo65x3NrF+MeaBylDvK+1leiRgpG2IwMnSuafL
bLVZpztsE1eQ7Kizopl2+K7odJHUo0uRbhvBqOCom1qfPCWnLKtINKKbCVkJ+w9i2xJr97XsAcka
mcD+w4UvPxagDaVBNLozFO1MAMzm5CEbOHXkIC93eijlTi2QVMVYkjWoBSOzTAx01J9iKvoKvqcl
9wl5FzPZ+Rhorna40R7m8V2Ae5OoFDv0wfD7SbOiVCRqr9QoDWu0EKCZOiFWJe8GzMeJWoFtDwJ7
5+IKLo1LmwdZnkvdkknrw8EwzTN72J1Uf3926dIejkUTQH9ajhPzrhvnTcrx1Xv/tUIFOm8B6X/0
Z760KCAML1YLZsvtLNTm4K2Eh8dccspygRFuvjgoZVMGtHtvBkKI9RGyiY0wEUleeSmrBg8s8Yho
kUD4MtcGv+qrC/X+UYZiTwJubO8d0g0lu7TxUhkJCX/2HQwjo54Eyhn9+bJVIuQ1jyd4xoH4r7qz
k9aWhJhwFGm9xNZswAi+GS7Z2ogG+zaC1JXGG4KfqYxIyIoVwwK6Ttkrzo5EAdvcM5FIRzV5ZGeM
eZf2yrUY+wHWRp0XgnFnVFkW4haxMla9AJCjOGkGGvoWzH4PCMCS0bC7BarvC9Op/J5TQkUpasBN
DqLvpUcNM13eBr3EwvdRmRtLEaz10a/9bbAP6uZMU7ZoX2OySOATVb1HTAAsPQzfK5wRO/175AjO
bMlUPAMlgH1S+U3cZUI9JuGqO4KWSDi7WPsF1udAeeDYRKdP/OFP8mGqH8fdW7rzMo+s1xeWWsG2
7xxgVDCXBf9D2fHmginUT9d2PfCErxfeya886cAPyO2/+iZ4GRLffog8c0sIAbSKeCMdb/cGUeFt
QQ35UJsWG/9TtOExhL+wpjQq0lb+XDc1pzKcozGfpYN92hRlIobcwaqnG+5bja1SNahAylxJ+ksA
H2iV8JgV6j2lAMNfzFCsUngQPhLSd3RqP2IdV/PtiGPmS0AsItYQA/54lCHIKo8vpDXChCkGkMVJ
sMxnMlOAuCohh88WB7nCD21zhRzZcOiJLpv/nLwmG8ITk/FkYqYYLbLfjz9QGLWdnnn7+BJMezF3
PRkEidTFIKMcn/yHlZ4/V8qL7RPq4SxOdgN3hCubtF33dNgMV688SSZA/HJ4lpRJa/Sjl3Ie4S1x
zTMGqymo8f5mh8g+QvbrMp9gYVjuUma0oeDt7Anvs04c1HmhG31idHQLLbjSJn/YHaeY30jU//Iw
aFOY3G1pLMv2PAORQwI92f+4KRt/HHn1saHw0mYWaqMaNIa6kt3z6UtR40XeefgtABbQBXC+sPT/
3B0x4miI69EZeQvYRRue5tXTfd3Wtxw3V8c1X8TqPX7cXEvjysnOXaqg+xSWiC3qsMXfMdR7H1ay
QbXmhQPFM4F14gWBzEanHKqmrqpR0X9JGpgoSD5qhsOiiytiRn+p0bNv7HttmtqlIe8jEjNunBZG
eATwlt/Dy8INNreZlUV7niQGYdQZmXZhFV/MZJ8HPH/T4pt1wBfq2bsRrFGiSxQNr8zeLjcQ2dnk
hXo69TNPjhV14pP83n2RtHzobRdz/QHUvPTDvZMIqRU3j/prn1tqF+ewnCVGfQYwtTBifKYI8lqv
QvAfAcon1Jbe1eHyKfIdtMT7XqfT8xC2Av1RaHAxtsLQA7VCyS1XURMwYt6hdoQDV+8VbkmVs764
JKFi8NvcKDOC/GJ9Gs/6EohVB0hwx2L6NyCXTow/bKH83lndp62aKDa5XwspuMVkyji5JIpGWjv7
aDT16WRgIr2TYdJqDtFu/BrLjXNdPUEm77QSrrqchjN5YiipTRPZHZ2Eic3F9GO/ZYFcfVtJbnMg
3mHHq4ykK7aGmtu6zPV+ix5Kg3ZwrLB4winktR8h4XDW4men3uvX8inX0/mOxinPnFLPYFgUTggs
CAJXCbT+PcArd9BRZfOo+y37UeG+5wa8EV4tb6Mh8F9LcsUZIsQ1pbd2a+qCBH8ikAcKunyTOvrD
lylr1LYQdJRlGcBvn94GqbA5tDvf1GP9bFWxFcWSoAHxjnOhUXmz8s8b6biJbL/O0UJxO1OQEYH5
I5FikAjm2jcwMnYo7Go609jgvulEptPHguo07TY52DsvqHwfFgoRjqBF+AWzd1enQfULY2Oeq+JC
ZcNmdcPtjriSWnD4tRRTrrXTWdzlBdGbgNF/wcG5CPXxmgbrZJfrJYToen6/nJnUJvwuHTlzC6Wt
1NuHSH8kJmqin1zcGsXW3MJvfv6n+QlSgGJxuSdDg31Ga8rBi5FqMuows87c/Ay23y2n8sh/KM2Q
s4BIwaA/2FYOGVzUHPsgN5jMDazcNk3SlNpeaugTl5qSkb4ohvqxf65D85/p1OBTQT6pFhZRPsal
knqvDNd84i8sH/fxZRyo7iWAm3oGNVpGB0GV8QjHxuJDcstkoUuH/eCW4kVNmBr4MqLIQaEP7qUU
acjjrf2sNWFzlmeQBDQAnVrOt+KZZytsXMf26Anj0SOj3QxROidkwWUAw1M8ze5CLyMwvwg6ec58
34WK2GiMAWOTXPWE+YNgnTqlHq+2RuTweApUiP+2Oyoz5hkzGik0vwmJpYXeI8FshEbr5WZ2IZEq
zx8G6L4FwHXGxhFd7jF34XJibyLKVQpbUYi3TRTzPm8iDChKz7w4eDKkiy/kSfr2pNYMQ+60lA+q
O6ktbET6umgpBELNoQPfc10KzeNWs2NPfOTnxZdDf81bfmenHLrncy2xgE8yQWByB0eUnV93hHW/
9cXr0RD8KJ5oe1IIuvwwRRTvOiS8Xz1WclzrmmccGmCWuW8VRMRZQidyh2+MBzrHfwwolFKOO7+y
i3zS/Ol/t1HtWGDxsvTrBw==
`protect end_protected
