`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
JEhjZ/548BbwmvjhE2/M9SqPO9nkdpAXxJ0vW5YXOpNhTAncy6SjqJtn0Xqv/qW6htKyyc5P0p0e
X0RIqNQVFPXdy5eOYf4wZtNwzuQ+VD+yJCTCBd7ROdla/MKo+blWvieOn1kQnIywvtJdK7GQf3Z7
sNdJSryI522aSpoMYhEiI0n5NoerydF2mZ7tZ/5P0bDcbQ64l9umujdtsWPd5l6KbOFraCQ6FIV3
x23pwIhbqCeRdFtGYvqMVeFAfr/Lj3228MIMokJOi3CkR1TcC0vHJdU7AqL6tnLH6uok/7w71B/6
pxQ4ICqfk/45QJaLj6nR+cTU1ZRXWZujkqW2xA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="SCVhETGgmsdrJPBgQBNLkG813fwu4cMv+DD7G5IDDDY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
l0stoTd87Eg7MxBsAWlarGklONO+P4sGEPgeyVhisgUvoNofBv4edyH/RzxvygjSAZnPm1DDp79y
SDFJI3W0uxPEEK4okT6m+PJTZ+5rBwOfDnuMvjekqQRi05sTjn5L5dtfdE/FAAZR4SKqE0NjT3g1
b/cyXSN2eETEuNFci6cVScna4IWG0NiwrDAii980Ac2yhstNSTbtDEXdyiEClsdcbI1B/K/LHbUq
bNPx+26yvZO4I7vq0rDMFHl9q/jfwdi28N/k7zP6/7f4rCMOiHBS0U8RJm1WByL7Y1aWYJxwtpxU
EMIn/tND201dXmM2fRBByNWNzd6JnIdI5IdtWvuBiIiRAprM20mX+JL/NH/TrCUTbtu077KTex1o
Vq4zTnmFYem3IEfOc3fyrg/fLK5aCOo5ZCcP2R25DwFj86mID/3EEjmnJ+NaT3HhvW5kcucNGLJe
vsp4WmU4kNwIdm6+24BTP6H0if7yeOcvdZipo1kpjQoOd2OeeJvr65w0h4zcPWEW+fhI5lG1MaPg
sDEs8n+nzS5aR3i65acCwSTMq2jUFt16IkHkW0S3G9K3owvCpk4HnbxfDtvoLvk9XeG6Q5x7JFN/
QL6FXUEx67VyXkxacV2DJIEwo9zDggTA3uLnbPPz/qMhdwxLedR34scd2kGPujK4lora6FeoTMnt
DW1HpqxWdtLhdN8Y0SIGbPITNV2Uy50Xd3rv11xX7QkJimz6UM2vucLx/Fa/NZNBvv43+kGPhpfN
+GnNbfFOlkPqKAi0CXYbc3Z68j4CewnTdMTuVH6+DUvlEL93VpU2JknmPn6A4VvBdFCBJ1UC8uVM
aDoSmFuBCpkrKZW2Sv807xoJMvDhq/tepLjKZ/7nHvG46C6Ny0aD6Wy+CpFWtExc+78gErz4AevH
IOYr7U3n049jYqQQtApe5BVCinE/6gRlwb3zoz7ml/SxyTRIG+X/gRQePzaSMFQtqkFB+rxDuLtH
VKUvRrsnfTakDlCli0zDyoHmLhwRPJprGgVpmfItJYeyKJebuof8SpeKJ33DDWssYbvfGdmFGMh2
Z0DBLsdvjqXBaypOb3VgR5e7uoPdaMkzooI725Xbmfbb0NQaxOHu9ty0nMT/ginSrO2tb6hYyV3w
nSi3ZsaKcxR4wcIWL94bobCgDMkmowJYBBE57nrUKchCABWLrgfuJbwcgGt6GkSxyJOWQYqbBKIq
vOy8dwMUT4PN2Q2lOIXP5c3lkXS5vsJrKIlUCz/biDxtD5xJVh+MQ9lQU/9NQhFW7kWDUEH+cSEK
BkE8KNpkvPNsp1zCDCGOioRDrEAtZQTlBjzCqWf2EdIppgQm/rB0vpitut3hudEJlrlYjjmcVhW2
u9uM/aOibLa8CxcpiyesgXfxehUlxdeCU662dveqjzP3orE1s2K8lBMSoLyLUmMAec+31JlqEC/1
SlWUjJtNBQmFLKG0lb7U2hS3k+YW/2ww+HRYGjFh8EbUagET3d1wCQ38e44r//xwcGwR5d72H1fQ
a8n9csFfmQdIx0DGSN4F3kEq2VWkUPISSXYHuTCyIusd0wrBe2YYZZKmDmcs5+uVpve2O5nkOHi5
JKdu0ti+BB8nOI54XTdE0PVwpe4AzuLw079aqO5EqwFnVGAdaDk5M+LU4qu6mYJx9WSUWE+78NAO
w0kR7X5fFw6WwrU2/sYCQ9oLrZLR0NLNBYBwgae4fmB5BS14Mkq5mcukyte4OxV8r/gYEWp0wXjI
Vwr9wCT5r8JibiXSGnGdTvKeTVOqUcGcAjfsHsNZMPC1VlGLbgJ23r0KU2jretWM66lR7y932dUV
mlN9+lOu6aR65TBeqTmT7ybt3ZnnLsON3PuXZUYx+0FMYxcK5WVzM+PjjHnRSwjPLY7bTPoCKs5+
05Yx69Oen0DyTeHQfVHgnsaOVlkmUTCJXA+z2tTa0PXYKSWWDl9wFkhSXCrDVqRyToFTDr6Zj7d5
wO9kvfeNaSdX3QAA+ylzrg4lI3W8FPr6QxwcUz2uFPG7SasMDF08hhMQQHXRTTuk9+L2rpKqQZ43
lem5HDVs/CH4lEf/8Tdr4fJYhHKcEqJJK+J8gU2PFx6/aF040pS8W1fNnx/DCyS62r9dNPhzD32e
YXz3rhLoxbbaxrrSyb5Ygx2Bynf+4izOPd56xrTv2EOj3cKVzhRpvIasEe28GFCOYTZClu+K4KrZ
E+rqzoPys0S4g8KEOVVLFByKYjeu6RVorK3V+9bRXUFe+avg+GRbhAAEw+skT5XppG7B2wMPZ26A
W2x0dSVdcdldR01IVDJZ52c5bV45CRukt4EIODzxMhmW0bgs7I8r1tOH3cBW6JdishOWIsWVaMRl
SWidLDT5v+3dG5j7y+66vcQPS83xOj+wN8yu2HTdG2iPjiW8uF7oUVGVVlyaweWx04VZRuLTY3bK
e74tikTyeq6GNYKsf7JghYxzMIguzINXekAOUCOzoBuc4SuxVT68yS6t6REHpc18Atatw0FlZH0u
fjyVYaLyYAo1PlpLJGAm9Mo29bT5fIU/vqX5rv7NhZ7EoeWViGwOwOQNfZVHP4IRXWbgXAmcebF5
9umhcRRUYnzK91Jr+lGy6EOV+xxpXIq0MjbCDpIZUqd1lUOsjcuiwWcGqs8am1m8sYPMkQCtwY0a
SqyXiD8yvc4WLqGTPZA1pwZZcmaNd4S+ZbhbWTLO21OrNCAKRrPbahEabA6Tsb0BNxWnoksus3ub
DYJpFAo7LI/95n36+h4o/iSenDEIP8kU19UlOZDh6f6MM5asO7hP34mOEiM/9OukAkDyKxB33nvU
H0O8oWrvtOteb+lGbttkhQ7yBydn7exo6faqsiOpsukXc4+gTCLuEXEB+T51Pj/zWxacy1XEmMlB
K4CrQxCBCFW2PrdeE6Z+QryfdoUfy+1cmEhfSoB8qKWs1rv6NN/VMTYPOOlhWyCZgA+AdEpIvlPb
o15TEcAL5sEAcP42TS0mRob2rnrZVHroXlWwq/ky7VRJqqXK3yasVZmKMcSMKjxBAf2+1HBKes+m
t0v0QPSz3VvPgff5ImYAtwwoTtv8ef5AJZIHlIqVwWSwGxpJwnTE4HDUFm+7AePcYpTdcvADpHS1
6Bcs64SeHUmrHpt1w31C9llcJKUiHIS0OnY33wHdIxFd0nibyGvhld5byUAnqn+Q6AaKJwOJUU8p
kmGb5+jw6yxzf1Ju/8Kj1b80ybwCRCrVsM8JTMm+Y9HwrMNYl4PmHqc63EDB/PU0VBD+iFBubhGK
5GDWPrqEIa/cQyV2djmm/uuozB8fJFKyaFLh9t2lfZfYVfWdfyb6yE/4dzlcN34wDIhvjCEtny7a
Feo+ZVgNDi9hbdlKiR+XIUs+3fJuMSVVSif9xzgaQvlGclQH74bjGavgrqPUwU99mc/JmwQIK5Tp
cJhhMZEockv+sRlbti8zGptrvMPw5xNgHxqBbNhWDJSS84OeLxTiQNfmp8Ra6ut0EzFA2TYtvuS6
3e1SrEELfGnP5XlbFPTSZi1jeFUnaaA0GkNMTWXNp/wf9ZTQmteTUmgvHGsSRgYXwOTS7JJzHE9j
o48MX3O2iD5qo3/WGeBCRrVF+SgdNen98v1gh68f/+i06LQ3P5AqGW4LtNrdJHetlPk6SOCrVlhc
EQHmOSohw0/8hz3dNrXZimdTpy1Mzi3+PtExuOv9zD2hf/f90q2wkwqS4l5vorbn8QPka2lmZkyO
ZvsCO3ltVOXg5SDWbjaYtT5TsGdCf23z0kvsajynpIYyrzH2+Q9aRqWP3HH2U0QLmxAzXFUGWsVo
Qm6BZd+qipdiy+QAd/LW+wq13Myz9jAqxpzl4+jfEL87mdVWXGbMSsw1BxJkiUnTZEzSa4h0DJB1
vwOCvTKG7vV2C/E5cWf0JxRou3pQbvzTlnX7rSri9D5qh5SWdOhYNW6qLLytdGBheEt2W/9XpEfb
n9L8x1VT2Oh2VkYaQiTVW+yzClb/qE2Nva73ygOedHWMe6zcmJXLjNSVJU7CL2Ct/TPh8L+YI3XB
NHfVksHWB/AIB/3id/C0seeembBCYrB5i/WjB9VSyUAEcP5SqZDhkysLjsjy4gh+BP6eOmUusM3H
lsR+UU7i1WwFNGaneeqn2eXFzO4VYzDuN2AfCS9P9LdIK3ydo7szcIN5aIE7Y7LkpdNt3K3Yotgy
xUXuONE39IGYWxasvRyt8omB1EZx4gUw89KDZ/bl2K67sit8OazIBNFLr5r/YN3g7a83+hIaF6/O
Xhwuhu/J9QAbylhlss0NkoVPg4rdsvF7QcNF2Ramgh8cvW3WLYDNVbQYq9He8B2uWnX4mcMoCNsu
D8JHvjLizeqJlPWZ+njJ2SkEx75IGoWhjENhBZyEqpS6DEKyzE3gUD3lyoxdDOaqWRwvVBuh0Iwt
LFoZqRWfkuWzpYUoojLT3uUKdZO1CnqbLrn6ce/tegI5qbY+gRgKkRokTg2q2XdCj+ccAbSDQe4R
nJLPFVliPrbAeJgyE97ERDnPhAFVPaoA4qiCwAAT0x9Zy+qURdmK5fQzgYhBR46xR8oltSe3GSgG
GSi9RW9f0fxCmoW/tqe8WloNo6Cgq7w30Ha6DVaF9dJxnAxL2JZ06GmP5xdqobGajMokeiSaUgoN
2HwNsiXIgJ74BTCLPooRkZVLB99QKtxtuozm7Fwf7snJX3lwkvtsfVpLCyq/n61TKTW9KR7JtHaL
4raRjZ3N7z/ydCN//Ly6/rN8rvTQk0FQClqIi7+8rk+Yue9w5TUJjPb39GiY9ee2DjAZjZrJIgFl
f5+oZTLvlfXHi6CgX3h15XHF0Kdgbwm5jwc8+sAdvz14tvga34KVM0k28/98h0XEGlvliArV8qt5
u3aycKcnI01ihHo3CfO5TacFWixyIeNDdOmjbBG5xF/lKzwX2LL525kXAKZU29KIDUzWn4MB+jBg
D2oVLF4EfBIQBqlBfctp5YlEa0N3MiWf6dKr/JTdd6H3zSoyX9or6eeLo/KRutsXCqMCaILiQv+m
7dqX6FW3cSj54Vg228HaKQ+Gu/9e36SCQKdqPwVVSXL7AdJ8cPc54F/3+JS9dFhskfUEs3lQe0ep
9UNwze1r2/ZyolpjZp3qAFDU2D08pIHS0KBLQ6x6JyXFdjwFXFTEoMH+wbyhugVSHxQEAd6egA+8
fLEzsNS/MckWzdJujMEXQ6PN15TXh461CXbdtq/W/d07+H5QpeSg7mAheskWb4V1S66KSlHfyGPc
5Nb23DltM180nx1Fd3kIclkGcQNgO7S0adDfN5IirqVBpy7l+8p1GzbFM1p0yUl+jiNJQvT7b8pV
r4OYY3BGYhHSibh0soy6GhiCLoMle+hLAYlf/gPzju+zoONS+SYounlrxVpfLVW8jHUXEyHN3EJ2
q2AKjHM0RV8QsjkWNJjuoFhgW6rngv5cHV3GX8EgxDOr7t2zIvgITb+IwGEA90Aoo3IDOb2QSRMo
XIkU5KlBSO9bqa9qF+DTlFeXYO8LXTzgEO2OZMdHxyuxFlLDlOHPvuOaSg6lW3NbRhC4J8f5kVYL
Gt9uBIIigAahqa4oWy6zlxxdQMPqUs21105AUGL1AJCfeqgOJzb43zJ+r1ZhaRuUj1uFdHIkfC8x
14uNcflLK+igsIe7T326aH8vZ01zTzVHDftWmu7o+jaN3MYYNeGkj0/WwHcYeeJJwUNN7H0E7Cbr
WFMj+uUBouICpioCpcDN8lqyXEDFemECOaEp5shqShI74iMFGeFUzGtnnHVhVgiuzESg5Mwoh544
PowM4nGybUFDm7ukFhqSrlR8YP/Xp4nL0mIEBIyp7sRJO/o0H04o2KjlWo9yV4B9ca9Q02O/ngHg
T7wNOB0le95mJCGal0m09w/gvEXR/IB2zhBmE+9oODTZlnqE2oAtdJeEJvACHnMFtsPVd3N2EH+u
8k9I3WsBMWKOLrWZ7bElS8N9NtsTR89Tz4fDeEOIbvwWQ7EF+N4TdOMLEmVVoTXEjlQuUqa1KNU7
P7eUbIDIWPO80tHX5fttqyD9yQQc1E23SBZMXXOjs7JFBRjnu0qVGYeXbsf4bntLzgEDScAyC2Ph
zHxy2THJomy+nZYUAANbDDvonTeAOmeiXJCt8k/GbX4QELfa1TE3j9ElWX66jhzyMqIyPwDlDaan
hT9S1CcDUC81R1YCq3qJO0a2ebixZloXB6cKPCsmK9r6WArfXmzaBkTljEpzieQ6buOKjl+4TiVN
KPxqyo9niuNJgCvcFKabTq+d0VPUbwT/m/RpJOBIkoJdrv+dqOM/L6wrJBdCE83SbtFuHrmI/d0d
uyMrwnCfTTx2EI6GYfitMcTiUIsNSfz4MiMg9wXHi9PADch10PdrZ1VDq0DXKBvBwiPpeO2hwo61
0/PmJHHp+gwnCIA6YLQcWr6mwByOcMY/htzFFGhaFbE+In+iadlqR11keXfdvLi+O9BSnIDfliAO
Wr/Spyzw4dYGo0aPERgbypM7crqRzIReM0XFUmetdGJ2RbRaxWJceLiRNYNk/jfoGe+ZWZ1pa0sy
1STCIHi51jz/4QQ72jS/eWTl4auG+mRhTtzfsi088t5tD1ltyFgLe5H4sV25m/0c+f28lsenFe0v
BnwRTPOFM3WioWcE7n2zKnKUro7SNdlqU/vEtgxIlZIFUIlhGM6pzhOgNq+Ou/XGSXbHBSZtMfEH
fJ135Cu9KY+uCl+HIxTBCPKhhOuIHruuadesXDZq3MUqClEeD1eDpR3yr7YbxeCHdekKaK7jclFN
VB6Ow9HdfIRJFf8YcRD/J2Zx1rMc9TjKagRrVG69hIBQKj6YPW9T8+Z98079py6wjrER0ENfS2mr
x8fVyjWidYoPiU+qwBsE21Xq82dtiwS7zv+B5lnFy3YAIFhhaX9UY5+jZjJ7P7pLc2PT55rmnupX
6NIGy7hwx7YRuI6Lwnd6b8r//aCfHP4hDPR+A+otClbXk5JnApzRELBGxKPHJMeHi+AeVbkVuECK
hMpdOeTFWaz0rmNjaTyKUWTGYthpEmcvzgooBnspPDI9AGhFMWjqenCtjdPdyi7qI32hr2CW+Un+
hzhPXOavbHRfRpajq5jNpxfLEo/KRY84UTbF4l3DesjTDlmCUP0wHVWZ2Rdb9xK8fhAicEIlREpx
VsLg9R1g8jIfJ3+/TnQkxDlE22Zc7bn9OrNwkkuh2y2IqSeQahITt5izolFKZFJwVrhoFym7fitL
9gtHcdvRPOuB8AHKOIznqfz1JqPkbMcBRu/YkMEx3lHaTJNdQUqt53M/76xeyIwpwd/k4NTtXR/v
e93odFvMLOd6aEM1fjlyYu7x2of1niKFlfHyFxa68kDvTaxlLtbu4fWZjuocG/zEQbYbT2h6k0HR
lwa55R+E9xRtHhKMezWzHZydAk7xcF6IIL7VKCv0xwouXyP04LEeZWvVpoJwwZQDBr2fw/HXeqGt
EK5I8XfdaC0gI2l1Cm4RBpZMtBqr6G4NqZUuqHBfz2ErMPKsrGNWiPwrT2IvjoJLMGrIGhuBKBLB
XfB54viruLdGmqOjlIf9ave1E++xOSRCYszCe2YMj8VAftMeyWSu952NF/eyxgeyTyST3l8erpuc
nB5PHEzDS2oFR9Sg6zIqNXHjI2CAnV7E6kWYwdyQy5M05ENlPPkCQkdLJ7A/ezmY9zAir5mSZo7C
qC+PSx24uzKxOlYwvxOADIlEVbfyDSVjRv3gpAMyL1SKz01f/zfgbr7rX/208T/TlozKX9YUZM+N
Ni7146FxsjfvUjpiRAvn9EtK3ut/MBA+iYeipOW9Hsk/ihFXB1yCshsHRwbnZRduZR9/glJoBgGJ
gkyKZriR5jVF2isDsFvwLHLswjf09KbdgBImYWrcnCIluUPIqwdWPseTlflZjnzzcghfcGUiaDrg
TUAdhRGSNKQQaCFoq8cxcroQcoUkRO798M7rZm4Rmjx2a/ElYbpmpMJVLQUACPs+N/ksd4+aSFGs
/BZOYhgu4wVB/2DGLyRq2YL3abdxnr9YOow7VZPXvTurpk5xnGnlE781k3IBcXN4Da6TB7u8rm3N
fCXyhIoy+YAKi9yXBImu47HglXztn0WPgLljYYol7D4XTKZZlWrYGFTT5NyButPRHQT1VD7QjQHF
R2mLXbBhIDwc7U+eQ/G98j5SoLG2bMeBp64DkE78jaSEsMU/p4UrYR207KUaxuE2EYkmjFWyli90
LiCflOAu6lhSQTlI4dm7NJ1NDnfvK3pSL9s6ahwru5jcSJBvwhxe9UMKa9A1VNqdkaLYEBJ+o4h9
lV0Wu7Wh+DCMRI+XNjqGPdoLUTTExLC3bfJbScNkjd7M49cjpQ3F9g5e5t5sCJuZka5z9SPJFHna
mWBU2jwijfNmgw7oslh7JsspjXycsg6FamwmQAj5kxvsKut1ByUlvS7A35edQQ4T4u8lmD1+EDTS
Jb6WTGZFw1fq2w5DlY9ttMXfquTaMCjCdsgRLVMV5PVavRkvb6gQkRzMGIBU9ItlcEkuV77SIRF8
QR6MRE5kt0Kxagpz2CFvbQ==
`protect end_protected
