`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11136)
`protect data_block
qEJK3tm8wQKBgHfqGLXmpLTcTKTy5DvjM4UEg5LxUT+4wa5i5oCxdraCo1bGE4CIpJI0Ap9QO37c
6MOGMQyLSHn/eN4OFD2GJc+i1pAjK6BhHRAzz1DeJDA62iZR+BMcwfmWOvEB4t/U4nzAUoADcIrj
5FURxiaX4T8D6kw82tDGyXZG+giq6fgmQXVJuGjHBYSNlv8k1JdChUNsYGxor/Ml3pUWbDKWgqQo
W1heUsR09Fxv6lDYXvhZiQZAhfINUpUxsA90Ct05io7BQvrD6WcmVe3hRrccDjKtqPd0l/DWb2Kb
W+yF6CMGCJOfv4NGatk3/naWGpHfMbGA7AknGtYHkbfOKHIF6ON7FrJJhAVYon7c9bEIQVBMpD5q
gXJFrPFLgos5BK2ByLezz6cjWd1pduBSuqMZmMU+ptqNdtIbzFbD8c9RphZBez/Li3XK23D3IbzP
IJ3P+kifFI6yv+ihq1EJIeYSYsESEo5aOHbtvsleCMdn0ikxPZt6emD4F2D12QPlE0Y6NwW6vkMG
7KFheeqA9vxBcAL8RWdsEC+/b6A54F6rFCZ8VcqBQS0qsgVauYHHqUv9BpT0xAdZTe6mbHcl73EE
3KQaArLtfSzZgCAoAbeDfWeZ+hYP4lSqhIs51tsznb30TEwwfajATVMX8yTJ7CNL+yuHRZY/S1ak
3Ud72b299aTZatM0r5q3NwAUaiz8+eMBnIwH3tnyIPaqde8C2vFH+Z/jXi2KQ8mvXWVovMSP4cv/
sTpw7z92do+8HIS2wpBKU6nVyHmJ//gRbuW34caSkARwx9h9zuEIo+PQqIh/LFMsE/Wa1rdolQ+f
fEaLF+xIiG0VejMwvmQtWzbVHizes2PzotKKZGGQu38WvrP68uI0Soh0DVEivBQtwhNqshTmaLnp
1lyc0989KQveyQpw/cUM6QuumBdmiAX2KQWlAdrTF6RDP6HDwxOnwGCKe9QWSGEyt62v5oMl/Cyj
PxmBmbxXeyJzV/kAvwEtVSbGNSYTE7et6lU5XoLZDJYCktuy3cq5W3fGo7FaBl+37pNZhl1nzDXn
KO3+/gRGtP2SCr3G0UZc6itTEgvzcIo8UoncAqsIPMC8m4eEra88g7aQDPwRGZemWBxNwUK4eG6n
aKYL8NEbJ4EC9kgN1+DAMLfwYqwmF2PaXAqNSK1fAUPio2+myWMORPxzeiGb4NgZM/Dmey2aufii
8D0saU6ptg96uUjxKize4i1hJqt0vCpQIiuR5Xj8V+eqU+JneiatUJ1d+Q2BTr6hpeVoozlAWpSF
uAe+7NeUnaMC4WvPLXlspfGYBUQcLq2hAKiaLPhpyhUcdFhO9wFMB29Pl+4JgAswzJFV+8GOsUPG
aWOMSv5hogO+jE9IOqpAXshutU5hDcX2JTJI9G34QEY1hb8GHGp7VQymKQnAW17oFiK+4Qmv3G4s
hJZqCHujLhyvZ9ct5FXism1j6/1ECG+WVXUlzytkf01cA5RHHB0ITLHV20YDXT8Cvnhx5YcUgT5d
w15tSEqznNrgfWr2tBS2TF9ATxAzbnbohyt1/dDJSCbW2YBTpHht3cFIuMPauqWcoW0B+8n2ggZ3
IMgKY3Cg5U6CdzyxoHhBY5VMeDsFeRn39d2/HlM8MHJq8f9geFgkMH27ouHrGreP0NE7gl7dGGfF
cAHwU/sdM41Vp2IaydI6+519SkLwVyCvQdfljw5ZDBGaPhixU3QSY0dVACOoTUW8hKcyISo8S+1I
xm+0P5KXnrDNfSrvv1vBr6pfbnzLArcjr3iN4dXqq+5NQzemJaW94MuM8vBRpEWjE1zWVPxnmVYy
t6l+FP7Jvacq5Y3n22GQei65XauRa2JNUyPH56rH5Eh+4CQCSSLM1fxrCuu5C/2qX1LlmWasvWDp
ZbjAw2WO7FgscXbDQ1DmQUDpZ2WIeGjhBdiGgCte6QL0Vln5RhaIb5g2QBGwOVdyJ1Yuhk74e0OT
/DvTO2G7AZ9rQMar9Ue7EN92DRLLkJAgC/efqzN2sypLXbreQCjWjG9IJzSA6510PWUoaqioEEU3
p6TMbuMGq2y+gINzXmo6sg7Af8H1D3m3EGMUvZOkKgQrzCjta0y1oLVA+ZlIRXwzpCndyI9QGRh/
RmSYYUn6f0jgvB7Ne5J0eBvN3fU91LxZWzKPQIizlNjGG9tv+hpjk34n5d2AzVAMljNpch9/LTNx
WkIS/AjWUaC+HNcCV9VF00LKih1qu29kA5Q1GDKhFSQZoS2KWu6c9WF3f8zK1GV9GkzwxcBXknqj
c4XqPkhcEsXLFe5YWJ96pT82DL8pD51TnzDEM9K8drFpe9Gu1E2sX6BSNbBd54KyUWOCRpBvrEIr
6H+Xc1tlqW3FHS4m9HpVTvk6wzvcMnM0MXReZiis/hqOeRnfXvmiqlmP9aKCmh95AP1lufm8yl/3
5NARYcLGKciN0BlOrDBelbAzmT/FiFzrWInBrPofUkAw6nfZ6h5nCGae3rowmxUqOwl2t2T8hFu8
RlhRYmWQT3rdDzErm1p0LMfkqUlzuCHLlkspekVsuh2aLh7GFffkdQyDQKS0UG+zrLPin5nNJ7H1
QyS0KHOfiFeIOfcQU+C+jwdOkacSkHCwC8tDSdwNx3VhwpNHyGp5+OV6X+tHxF2navymiFZOy/F+
Dl+C/FnC78uFQr6Y9xiDHGi/+KuK2hsas1Wsq+i8UqdNsA7cW0Onf9Viw8rKwBWK0dzZ6dQTN1IR
ZRBPPgCCGz+fl8ii1rdlc/yX0ImVjsMPqcnLH0f8jqjjW1FBab2PYAzAlyKGQ30ic0fEgi4itCam
eMDWg2i+bairErZP8x6nwOP7EJms5P1l5V1PT8Io5QsSHYENLyP+zc3J2Y0+Y8S0zvRqq9QgBFOO
OCjOgA90ZkappStvPybKNUgIKbFaHRIuDBfQE5RCLbHknXelfw+g5xrdZR9szR3vRmHXdEV3Ol5h
zkKgvn/ZycsVDooEn4D65r/r6xllfbD0eS7Syr2/iqeh8WE1qkudyXN4W8O+exOR4VdGRw5lN/s0
HpYVfvsrC2JAvbrkKjIi0m+J/bEE5BqKuGg3/hGRVzslo3VQUeXdmoEIHpJZVsDPMyWKqyhzpsJr
U856F5t2qMl+EaK8Q/ndKdUM2NvwObnVfkO7IcrkX9zfB2jK1T6TdOESyeNZmlFY3fowUmW0nrGc
5XUHo65WVGzI0ifehbN8nHkQeeis9Q9pAlCVsFzhyo3Pf355QmHGN4qYgddP2Rx7OSOGim0d9LOa
SoUSoQ8bXsZeP6jthL9QyWr0gkg93VT3Bay2s86mKjUyAEkLD0YCUSrmdgrwdjBVIHiBs7YdC9Oy
q+8QP3++s0O0EA+mtDt3YRpiKpYS7UFwVFg8IFTKfNU//1q3LsgvEHv2eJtwl0IsPUtL9Abchaen
b9ikUi/Sg/iuVQQJZ25mEw2O1dMzaAI6CrKesGXywkx4KERfZ0yG7sF60VzpFcFont5ddAHUD+8c
qHVT/0APO5elqqtUKyfOwDbd/igQK99ocXNq9iq+62ybLbn2cg6vDoGJlpuwp5HqXq0YTyx7Rtvb
vcR2xPkW0oIP7Q/+Z2BbAGYxqy5VOqJFkF4CRf5l6cbUzP4BZYlBRXa7qqIcOgSfMAUnQ9gb3G8e
SxN0/T4i3IpyVN2Q1hpHRmTwoaUi6h1ng4D8kFspUQG409kQJn1lUGst5vygAumwikIBnA+MoHTV
xNC5VQ3OklCqvsUHHtU4KwYSerVkLKeH1N85SnOLf3IFZuwdwow1HFIO4fzfKu4YVkZHx3FZBMMB
JPyRbAbCqpfMCGtKzvuI7ZeTLLe18UNxThszXmP8I7m0NSWQH0ONg/PeCZsaAzFR3eM47SqpZH1/
3ps7L8PqydSzRdVD0acUkNoUUaOxj0eM2HfAXZWGcIlAS03J8dZnKYcCNT2PIRhgQbny3a5PHTny
n3KsJvib7nesdXFpNyaNxhi61FiwCcE09xu12qzErenJP0dpv6N5l61p0dwtkjqOCurl3dhRLpJ4
Cd5f5EAVnR2A6WV0V03lxt+YxWwWSKXR3W9NaGE7ZJ7shnTp01vWaaFjQr8+fVtLhc5TRt1T1jXG
kCZHIHpZ7JIkpWLuW0cSoqpxiaZ7P/Fil6m0dQMtL9kvZC/LwvThhZcFOn+9FHFVW0ufTVbXu0hD
LqcxHUBSFoMnCY2A3zPkcgy866cNVwts0dWx4MPY1x2ikB0KcgMV/y3lTC7e8/kcBfN52v/iY8U5
NqM7hPPnO5pYBUeRbITHqsXtwxt/p2oIg3cKlbjjL9J8PZqiM15VhsnnNH4UtmycVU7TrACtkySp
JmT/tiFyVuO2FCsXxoVLbUSnAFccusMgwmi8hh3irEr2xLutOT+NChne5pFomeg4X6MqUfmx+WVO
xLnIoBXc7T8T6yxBHx3hPVAcBDzu2/MhUvWks6OwzdU/XM0HPL36vHELiTzgHp+Z/PDcMZHW6tBw
uvXLz/VNETfltskGaF+TNj0eH1cz5Qv7v9NvJ1nS+HvtwUKsfdCwFlpcVGi4lq72O6y2TDaPh/pR
AHtf619qo0AiHRGBqOkhzfSfygAAoJOYpbE5I55eTncO8mP302QQbyRtL/r87kXBAxuvq6yQDMZu
0zXzGp/RJK9bII+W3M91DMzNYA+WQjYuP5ubWcl3j1ggfb95gfqyaGXO3Z0FlFbD3czbINy/3+IV
ruhEy0FHC6iNiz+3zaW+CQRNe98GCIztqlnOJ4DE9hx8k3G5VO+afH2jTnpGKEfQ1ixHQi5furhy
M0emv7uic4PulTA3rOdlTbU3zss8yQRwecvg8DW/bCVxhg08Crjt6B04ar+QwYMPtZOFapaJwOHc
/Gc8kL5j6hl1VDfqT1oEe7bcjgpRpDcQ9Vtu4ycoHo/nimjXgxmiw1K83NDL86ao6oO1xCPf21wz
OJeChhcLoIgvOByY3L1DlyHflMl6ImpyuxqiVPqHv0GpsP6BWlJtc1MhSD5Z6VI7VxdAqwvwuecC
Y3c5Puawb6Pp2DOUy333aUBIfRxTpQ41iMEdM/9tDA2lf8R5vJtvZLaQ/7jSGFVXlhPdwiy5OI7m
Lx3YvmoPgwj+XmRRbx1i/lJMsVPKUpWFDwN35ytc1MlidMsCcU6YdXGCIYlv6tMoU74Qn7CzXgrJ
34TIAzEGzMx2Yd7GvacMFywYFB3CjhZ58OomO98o3bYqsx6HzvtWsVeZi95WpVhF1KYvgMVxTkTk
Jw37MXGfqvn9O1eoUe3hAp+shGQGh5463RK7NMEICMgvh/Ya6q0vAXq5UUYqho9Hjv4z8+kA/AKx
75Qk+jufg1le1bixzmWtMUFwsMa3pgVvrVwKDNf6VAn2yPEqZrmeDTFF8UT2PgQZ2mfKCfwhuyLy
dqYOFz83rMlZQOH5qxTIOGmW8Ym88eym/S22WNlscz4YIeK825Kb8WFke4cZf3u3lJaIlttidnsE
Yob9Lf9fubWcAz9Br1hzYKJmCYJimVJlvwBjYIo5OUyuqHy/XdTq7lZWe5d5Ec8WIJpDIIMtcEdG
Vvo27AIuCQ1V5NHT/crrIPk4K9mqJYe4rwCTcjgJWfNnFSDZ9rvqMOwk6wkPN33p7oKMxIKrVlwv
rr1VaQMb2IQ643x4Y6h45/z4Dvdz3/b81HkiDApSFdKXNR2REzEEsBLbJyBI3X5Dd9HgHGpe7/7U
d+HuBWzsbCuTFfu9jKgrpZNEwgihPcsgeL2HvOskMdCnOPQXnMrKzQdC6PCYOPnEY+6fsz8FPLO4
EfFJMaIXCwGL82g1/WfNvCbTRbWHuXlVZ0WB4ztmd4W60xidXS90c9dIycHvWxkZHkhTzlwjurMD
vnkLrU6O4SANrhbzbniHYXP2gnJQ7uT4eNsizcuzj0R5nru7BcCnb3yDaJAINEBdoshgS0efyFjn
krmjwZQpXyRkxAA9q/1FOSTlILltfyRY0Gsv8DIO0WPpZsKxLTG2MHJyXv94BRCosVlkkSbwscTZ
h8MyDf+Wao/tFpcfdEhh9WuKRyz8kNE7AnHZGcqV5D3WIf6ISPF0ubwwiXFOXUFeh28WuH0jBng+
ffHJnlOru2+cy0psnvbW/K7RksrWBAQWBEl3PxntBbM4osx1mNcbWIID1qV4eVjvC5ZKOgpfWA6a
JOzz0v64T5h5/RXJ9YrQOOEkViPjMy+I7D3nEnNRpZSlLWr4guqkOtFC7qU9FxeeQrT6L3Nm6USz
mvEWTi0/O0RCFZ92KSEXIpL4pXJWxRu0BSiIRVjYgRlfTxeVY/VWi1iPfvn4w6d2FpbR4v7Lmklg
RaAJl66paITbyq68bSpXAdni7ybEnDvGDSGTGa2+9AvGKB3jXKMqSgSG1bCbt9dNNqvCylBB6h8H
sAE9kZKVnNSJGi7C5o2QiEUJOPszvHEaFqQsc2k4pIcRwwpIV111kp/d+y7R5iL+JtExxXO9rKrm
Ze2DREwRWgpoOfYtSfUYhy0tD0HxgvacYMJnmfpetS8mGOCZ77t7choWSF1tpy0TIamkcddDbP1l
P6UgtE1Nf0ZYWSQxHvhoF4zcyJnqGqqQ3O4eMgLGTgKGTNE+zlT69thfzpBVKnZlqDT7InDf/1vd
iTCx6+yk1BzsAISqnf0F/mnEYOZAK/2a3n3hJJ403nR7FYcevjKNKHU8MOZ22bnviuCalc7LjD9d
SJxj+Sh0htXTzWnsNQZhf9Nz+rVrQ3uMecpyVhedj30AjFOhbbMqC0nhPAAiiurW01yvKr/1m/PH
zFqBMUqwl49cUEAIP0O6vP9cVl2di72rtRo84nc48BZq8zCyGv7Si8lB+Ao993YHJLokmhcruiXP
7UyIPm4/txXC6mF6k1ELtNJ8Tl0XJ0TyQursICqNQlnAlHB812wCJcjPBx0tSnIbZEi+Drc6I5kN
jIoi1+1oJWfrnxCLnkY3cTV3hZIe+daulxytwXB60F4A1g0BoDQeB628lOpIxY60Xx3S5HI8YKVq
k7EU336j3pOCCUiRZojxA7qE6X7SE/mt5kafn4PGov8KGPitLtGMO2pAQ9CjohtFq99NNtDjtJ+7
MmTLTEJwSe7RDpZRUWWfEN7nfaQIaddjNwsPSBv0kHPResYyU0l6jQZu0wZH7XNgBPaWujUniO5p
UZe5a+O4deOLHQUlgQCy7TanT0FA6ttgAe1/C+gxexwxb1DGtYUtCQugxNZU6u5LUpgIkO5tjl0q
VwZcPyabg8pFN9rXVcRsZWzjQLPe98UjwJtXxMndqKgUOb+UQkOW3/gOOhJnJJbnNSzqJdTy9aZM
I0RPFtjRQS+sxNTnGTv90i7RCW5GonN19I2du3KN9rwTGhssdU7+hMiRIPjRq6nKfCf5oP3Fb8Wc
ofBiLJ3Vzt1x3HowHLCE7qUBW6WjSbggy5MIFpw/4FXohJww3l356cgsGp/ceISBlNyrTKHVcvQS
sb1oBygWMKR1bdC9G48erdDMgmjpSmXtd9LScIP/TuMfjj6QiuVc1Pr4qiMXJ73H3IwdagP78AU4
3AGLCcxmNMAO1xPBPSvgmcRg7Ydp2uHKtPUzw0BQogkNr2BWVq0/oDh3Fd9LheV0r7eZ8lqOtxGs
7sEMuatBfxNGKkdGJTD8CEVHUGTIju0TLH6KO+EKo+fZ1dU3bwLZx5VNPPsRMVcAZgnRxe7c1S2l
9OZ7T43HkIjOw2pZGbasJTxj5vBadV6qWQL5BdhmDm2I3ozcCYafG8M2/QryQ21MVyK0DLvn2QlX
EddMhn79MqiUTmtfcnwNGNPaqA6U1lAsPIMZC3ceDqUVms9V3WhqCBLxlHTo6bP/p08QAJmU/N12
3OIe+CsfgXsB9hLE5EUfI4+4FNghBLK6R+qDVeiLVJ62xy8xPtLI8yehKVkPPCYTSNh6ec2Qhh0j
ZKpL0kEEnQTu091n1wakqCWmbWf6RTZmOfhRRZCwuhTPc/SdOaBp6nxN9sIGrj2dN6XCY+81+Wt8
vQM2C2v1zKa/iTgnSYO21IiLONUPwWNJ7BamdgZtVsghBksacD4sz7TiMfCeNh+jGPDKtNLsnYcL
dHlw4IoZgwQzGSoPtIR5ri/o6ZehirsPq4qnPu3w5gDG1f4b9IsnaYg7M6UlTxmF5ghSqq6gJyuK
N/FAzW5DqlFbBIY4r8ubn3CXWc1mvKkisa1kiN3nO3LMCtvnSr6nkzY3w5U5Eop+IEmUSHQTioUI
fw/wzv1OYck1REeBg/LnprZ0WtxCY712Ql/PacfjmL8sbfGRU4zis2X+neBscoacTIqFNVm9T5nr
6OcFcXwVwOOlTSiAyWfo1XHyCy1OwSalJRsJ+1CWiRaj5ubhTBsnH0B2n+KE1yiiWij96SzRuGsa
lfenToU67ahVaXEcqU1C0rtJDzlYZ0KHh+CP3vpzHLTwVgnV6467Hn08P9oD353NfvV4WBTdIl/A
syheCsJ90t9y1hyiin34bXh6LJxM9z3XtMzfeKxhs2RboIUhvlqpkt5hJOC8vyn5xYmW1ebt0248
lnU77XcAMnCTtAU3gU1oGeoIm9FWtGjqAsGAPYT+95bwuWqVF3j55/w5n5ydf7C2cJL83BljrHCt
FaFdZQgzH5szzBtFF7hZTCOZUraLmiQ4SEhN5AhIPQtvVGva94Usq/ap+0ck+e3YdIud6NgBB8DF
dZlikG3cXkAnpTwHdHT00wK7aia8OPgdUcHtVQCs1zbzngmFkrs32tvrRBeMG/NHxyFI+3uu0K6h
o6LY3vcoKDMwvZV0W5vo0DbjqH9ixHsyxdgpkLcwh7H1xd6db1v3H5OWXadUPjVAZddhyT253/Ls
fro/ioxDBuUJy+nP8wNGUK8AXr3HXGecUOKh6l8QbJAxQrwGt7Spd78yWTD32T1TfYEwAotm0NOt
eEXtM8M1dBcYtTCYl1Un6f7zuXKcP2z90OXcRHAg+Ns9l7VrEmETuCGNr0guf2M1ccCSpQNvvBL+
voEGVLReNi9N520HF1OsbyPfikb/xL04wXOUedkWP4IALeiHUmPo4ykx8O8XN6pnS0Y0PCr8FvZs
I+Y1kZSVUdUPszfjK4HVEQhqL7Djrs5fVeozJIogTogCZzp42uwDhzazCPYXG8bwwN1t80Vpni22
/bDEHrX29IZiXj7OSaZTXBd+vf1HEyj3vkA7CkrWHcTpSU+cBH+4t3TgQENjyw1LMUgKTScdojsF
KZON0JQdoFO05AyAevIagoOi+GW4/TJC19JLQ9e1ky3B7LFYDzESGQopWeYhI9Dg8P707gsOE4pJ
Kr0Brb8t7uJhAaPoIRDPgdrZNUfbqdXlHSr9gnzn8nQJ3ux7IoBS4RnFKyVkZ2mzKQWJBTEp1/gO
x8cv9iTqlElUBm2+vN9R3IfgDzwCPFvI+KeVUnrGekRhWvI/ThO5h3wHdBxNh7VtABWciMWRHcrN
YSfn+9iHqkBYSkZFF7ZXEAtwMrMaSZ4IRKRtokApP21plEkmUTlmb9KRQbMf3um7huQ9QIovZkVz
DFomM3vWxTBHk5vXlvczUKy/igY2Hx6+yd/Rv4OjpPuIr49iYC1NfgmMeT53RrGeZJymJki8NfJG
3JYK/GM+YS4aBYCuwbpBBxCLUqWEEC7Zg2kMN6WeQt0oIVgHNQcJNlr6adMXL14K1P2ca4VPSJDe
vAUbdFuw0VoH3f4p8ghxu6yCQfbV+/RPOoa2CVC1qQDZp4VgGwfS5KW0hj9biaRcKH1ylO07Jx4p
77U9MT3YKu3AQwRCGEYmmpVQGPrwoFr++j+y2pnZvrWEQKESaw/0jf93yzLkUH9ZB1CmoWLatmfz
Mnivdbctv7FuTKMbHV3JCui8wNa7zPqAlQVSCKc4mtWH5HnGpZK8aKHye9txlstvtmTH5eJatc8+
fQBC9BBYdNkrrgZoxB1leExxX8H/jlb9sMW/ucDJj3ywHaCjOYHJhSKQ5LOb2t2eiTQlKg+4e2bU
EBmz7tOrhBHKfXGgFpwW+oV8kSeU3iYdrKxeG6IwEfIjgtt5IOYM7ZNvm2ePg2z1aJ1K+15QtmzD
b8e3olalXSi6iYdXxUeNA3UE7YxXwoa5G7SfjlIPaIvM63V65pctANZ7Aiq6puyAIGh6TEqQ/zW+
+PTqymVU8Bq6Gl8mtUqHCg6rBIvx55lcZpl9hpYtz/YcRSRenh2vBVUBofAHLsfp29Jy0QOiCuZR
faB4NqiUcsDHhpm1YaoMtgUwbjGidb0MdxDW4BtKjaNik0RS5ly62TBPDQ88BBmpMjfznMtlFdhL
GDu6V+T4QaR9hMRzphrbq9VAwlX9HsS3vVWvqFrzMNyhkqc0qiGjklY9bQFAlasvP6fJOyFpqWhV
JBI3M6J2cO0yT+dpubgE9R+Nci5fL4pMCFjeRN79uYlyOBs5XpeUxV1KvqkPRUJyoR3gmYhK1Qac
VOvdk/0QHU2lw2yv1lo61asBLgObzVEK45GnpSVC7SicnA+wuxNkstApMZhOv1bnFLqd6424NNpM
uZfhTHr0s+KKtWIoF4QhByyjqCOau/lVXE+FbyRw5enhv3990sgKmwtqmh3fsv1sWbnKE83PTP2Q
3qmClj8xuXo9l0IyYc/jN/br7368xYZnYF7yc9a1wNIBYU4oVvfsrsJ6Di8H1ccca1PHg+0FJu/9
gPQtNzr76gAp6ECJVmIZzpsQHwOe7ChpPIl+PD475euP3zCwJoe+W+jYcSqp+8X8uLr1o6zcQfsn
snfCW6rFzoVyazUbdc7yXOmrg5Zct+aY/yB9M30ffCyvkypfz8GT29aRIQHyfizOYgaPZaM9GrXC
DAUawkfHhVgGY4p0heNf/7kH3FzV0ZxYOHrVUW2jZgK60puq8EMQ7kmDFQUQTdFGAk8bCt3KUn3N
dNeGk3uLRWKdxim65D2rjEGwyrCefluZqJ4bZRSWONG/BeTnKZIn1ODvdQ3AdD4CJzin8afmW+hB
SJOGPHHvI8kewfj89IfE2R4FwdN4K8CpYCo0OnwJPr0p0WuwlPGQyx/o7/r1zm/W61AlPsxPvKRH
dl8WR39YUpcqjGVWvlLHBa2S2emWgmH0y/5HGYx9QwLuTxoVtjRD1YRnUtQL0gqS2X77vYec3giL
rgaRUlVhuvU3L7m760nKVge0zIyU3/DHwBxM5r3u+binr41bj2/TuQyGufOiNm8NdUo1yskmxxFg
wlCyxYeqrPRZcxUO1ykX8kgzvO4dPFA+I/WZf7K10ZJ1tix9A0R19pCx/rRqmCFkV1ycvidIehtw
cjU9d+z6HFhQEeu3tAZiAL3d/AaoaHCqoDonnFuioyc9AKNEwf2ST5kYshHXJbFZvdA7NMRGvod4
oKJ/fyUpnigxFsPobOdC9kCeHnpu1w+5EfZqCPw3cwYn6wuqXuBv9cIOWh1eM/s/c32+gRaieb/7
Zu+NCAL2v5Zuj3N421lwa3EvfSaS37PsYQT4a6Iq7CfjOMqH7Lexb4PFKbnySOhDFBRPQ2L7clpx
C2TJKzDSPndq3Fm1mdQByvZYJGGui8Uu9rHEoWFNUeW/+ckoIzFXH5eXu0TlRaa6LZKJTpfA6N6V
dBkGplWuFWV2IsLjCqEHMCD7+cZy2JpdejfAUWv7NDh6DEr6JA/6Z+lHjF+sRbTcyGGg8QYMbYu0
Eq8WkRe5h0NDC2RkU79vT2eTR3sldUSfoCIupzRBJBlLN+legmAseyHnQ9oUajGwRhghCCf73Du+
E0hk0mLf9rNSbbfdCRa7kC8RnxggucCSq4EZT1lcDdtXuNh1gw9EBx8ZEto+qvblf8Ud5/rQXKDG
r0zz7jA++0W73Mdz3Rqs6KFDjinTiDy70+DWtbz3j+ybNnYJm36oonfSaDst+wKKMOcAwCg3cxaM
rUT2z9Z21SrzrNzxEPAQnmwnb3p6MDpkNHouY8cz7yDCodh0GIHiQXSjPEHSQPp0L2vXyxV0Ps/k
jzXmi5lM5Tbe5i16wPdHf/ORpdCXYw6ONoJ6ZlLE/iFs7btGjOPrNQY1HPd5IKiYE5klxfRzi+hb
bjii1v/Y3JpDtbu8+/8N8L06QrHdf1zHy2z3Y+mSHO03P9M3L3EHxFGpZhS6ctpPnzWDhfO0TJLE
3Ut2KmRf7xXMj6VEQ88svNYypFz3I9FaS4mra2KR2bOhXlscJ6n+B7NZ9ZnY+zzAfMXmbCyvrrsQ
08LJj7WMg/bTjc5NuijpX6RrZF9eiCMq35/joZpW+RujCtncEkAQIm+0VutHAHMxJb6oi3ZYJC0R
ZVqsy1O+L/7vHsrJUp84ggxjZ4CX5OqbTDUvcP3H4iqwwGMdIhf/6rtMY2V26ywLjr4XSkcdbg/a
RWYi4nysUiMuYtgM2qT+aTw6IYExcAkrHP8oZ5X9+g8frLoUUYEU05gSUj/yz7962pGkfIFL7a13
3bmRQlez5sjYrZjfiq4VUiTlt1V3R643ADxFovgNHOm3HIZrCsD/ecSI7vDMtYrAF0yXJuW6kICe
y9FRCX4JGBwMYJM4ciZ3fqmR1Ha+KPkJOHuYLl7G7I0mFke/q/h4/DFvbMNPaaeVw7ZYdFhEQSS9
bJJARd2MaH6HyCIiC/U1jpI8O3ULku8mgTZLZiFqtjDBQClkD5VSNlcpy5rGqAHdvaA4UiCQ6xK9
nkFChfoy26NzV9nZQ1Uk41T4SzRTWueP8HQtIVWnsQjtoe4nkq0/bPXyWD/Bv9k7+AsH7MFlJteE
B0k9WM7sqy0OtV7Prbd4ispuXPuJiehYg6L0JXb3ezQ52xBIsFQvyQC4SA+nRLdIsIsB9OHNP/Rk
baoFDx6VNJwEAW26ChoZs9Pq61WUl2HiLvY9G90J8qyy1IG1m7wYTqszDUrW4mcuMZrWLTd0GAQe
iM80unnnx0LJN044a9KVljRNVu9myXVluJq8Sl7kDoFJchrHtATwCda8r2wRYcPj9oTPDnk4MRJJ
2ZXNoMBFUnxZhJWaZ2tUKhlF7UDMw56t22Me2XAG7PTxYKb5Hc645x592h/TFN6ZT8VXrXZLtl6i
hiIIFwmanngkWgdzNDdSG5JtbvkOdVz2nlIzMr8vO+liqtfSJ55sFPbKuXMlroo8Vfc84s9UdM39
GKge2RrQZqwgXXWK7vI1lmkjGWQ6RWXFsQpai+PE8BM9IFRZfADygbKDTJQAaUrQnf+pWRN/ni9i
XMD36bLO0NpQegGtX0ajfWYX+GggqKaqPcjOvZOxQH37Y+UBm/nQFSddE7HFGRG/sfzT7EyFImTo
6uDBXjzte+4OnzYWHFdg8NTJSE31IWx1g467TUiDMISR2hYN/DBazdgby3XAFs6zmvEmLTRouqKE
W8Pn7qtpTqLzgfxc71QgkaHwYiNgHAKGzWtvJfdaWyzQlm2HxXw4Fz4KdME5hVKZkdAPzdEYh8tQ
J1dV1Tc7wrs4xUCLdqn3iudQHtRIPj1faMB07sJpjLfLPKhXhv2eTtjvMBC+4mmku1+fppcodvnf
g/BnVZXFXmpTnrberVjRuqyOlhBAN/wo/IHWTu8zXAeMSkWQhsfu1y3oIDuO6HYqOL79oF9FR+DE
dVNN7Wcg2X8lhjMs4wGq67tJ7yj9VfWuSn1Ci66J/7LIuownyb8QPw/47GR5oNznRf1bRMnVW+aR
Z48KikhFek2n7+LJUd65C0mKQDsZfbihmX1pz8Ps9dOBKDE7m3K58nzrYUXJnCdF0POnE9E8+zwm
kqJ4D9Mc8yzwMEiyLpAmTEST4VfelEGknRYMi4Gk9HKFk/hDpCduMoziDrGMISUuGVE4JwozYI9r
vkjcSnLCOqzQhDMBkV4nf3SkomnILzwSqJ4pzTAs9906rvL05G0N9ougNPLXh4ackPLJi6N/P8ep
gAPQ8CIk/CzPpn2IELxySNhoAgTadNIU3pJjHJDiUTSpyOD4fUBQ/WfzchvAysMlmVA8sTh0ULSY
00g/LRDbQ8CgyhMAv9xKyKBCb6bpnN/zIwFuLfQvPsCwpoKC+FElra4DxacStFnOu53NhCTbynqs
2xj1+xzWtuC1m0Gy21hyfU2/tK4eJIqSovqo7K5axZNw1TsiCC4bG5tcSK5cgHASKk3jOjoDq+NF
eoRalGlVrv8rejr0IVu+J7eLZRqTJX/1Dm4CGKjEJs5Ep7i5ouOMRkiazsEACnZLt+Z9pc3JPC54
h4prUfB83pe7hsSWbWRq7BnY+sr9qA+N9Pf8slHpzzHoWkyIG5MzAX9xIqMRu1Er7LcUY0DuCv51
/rvP5ja3GUgjUmU31aanq4dj/NudCVG07H9ttFAEpZBB4ftVaEHqZGX3Gn5DcrQE2DjdQbdvxnTd
BzFBOx+4RbzkLwiCwXmqvzaZg+zsunz2tGqzufG5agLl8Taxkn0u36UHWM1LoaN/RKhquumVAC6r
lldODTt9RFyq5gQWE6CGp6MmkcjxBIxJQS+oqm3g9iwWlC4+ixFMeoe5FvWEkTlAY0w2XIH4aJEm
YuhW4NB18BlP+5o/FBUl0TnjgXbYSCNwHNXCCSw93Pyu/lW45/4OSuBud7n4npUwpKILWOzjn5Q6
fdg9pn6FeLltqnv8dEnu4EVnHL0OnmBzaISOrq5kd3Rph2FxwaV8Acf4tmcJrDImfimGet00Nhbk
eSZx727EZQra1w4kK7FpkIt8C2vLvRA+1zobwYZ/PR9XjsAJg3VNmp9gZMZE5IuPJuXzjprX5n1p
Kl9E/sYIFxEWlHbR8lg5ifQMgnKHGBpicv3OQrULPOFcb4j5doKvsVTPnVeDcZ3ky07/FL7TjBJF
mTgC/nyXdPWqveqy3ewzZIbtjQSkgVTaqGr7moCjmOX44iDD6+L1zOTSl+iss+G6JdqSIcrh0d/K
Wss1s7a4SfIX9z+VnicVASUHFSD5
`protect end_protected
