��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���=�^���{3�%���\h�:�0x�஑�Z��
ø�& eW����!��x��c(KAb�( �GK�F{���n*K��f�B�N�bd�f�@��PW80]���{�1i-<�nc?4[�O�����|?W�s��3f��.��K���O��|:�4�f|��̄*	K�攼��9��rj2[)Ի~:��UL~�-Es���R�^/��O��ƫ���D`�k�F4J�n����= #:�^��.���_�Q� �����?P?T�
�*��g1�!_�K yqy�W	��IW�0�L�$FuLg�{fi����t�a�u)��g������{�ksM.�甽J��@Y&)  Ԡ��L}��#��GE56x��&}w�,2e}ʙ<s�x=�r{t(��Ӈ�^�����#���4y]�&��BB��l�wK�U�P�_M`�I�Q�*���^I�������]��)�wz��8ۃ���b
���*'�vz�sRL��L���>鞴b�꒝j_�ؓPC��=������⨥ퟏ��GMٟݸ}�YL��s��%|���`P�{�J�����M����Q��6�gX"wzdU^Y� �kvf�:-ޯհܿ��%�����W��fH�E�	�*6��XHS�N�v�4�	6z~?Z�QP���a�L�z?P��/Q��� f��W�q"E�BZ��딨�t�e�n�kl�ų@}Gѵ����\�}x���^0A��HJ:	c� �¸L	U��w.)�����n*�"�ݢ��3��_����+K�`Z�@m�`	�����M"�zd�5Ο��ri�z&�w��鎛��B�F�J�67O�_⒈�
�`_d�:K6>;��� 2��6	#�n��7a/�$�F�a�~����^'H����x��>�Z�`{��cO+L;����gg|�}6�K�	C��-�(��
<��A����DL��DY�6���s���/�kQO�g�w�d]��z��p�jZ�/%A���FH(�nn��"��@]�v6��������Zd�7��Ƙ�8Y#��0���ޏl�M�|\mQI�e��C�����e<�8pb(�1Zet����j�O3�?9��0�'�0�����y�Tf>���1����Ӷll�����, ��a��D���T)�ۨl��Y!��}7·�������^�8�%�ð��׋�"؄p)]������'��\I�:h��[�#��yz�[u�Z>i��0Eg���C�+:���c�ħ���7<�B�/Y�
�h�Z(��(�9�d�_������w�1={�״�g��h��C䁑�B@��)�ώl�
a/N�_!;�@/�xXy{6o�P>"�g�4�0����O/9[������l�J��G-#��!l�o�ߐT�������pw�G�yęl�-Ri�^t,t\�8��}�j ���t�0l�v*�=�ڋ�&��\�:�Gӳ��8��I�11C���ښ�-�&��������b-o0H��g�Va�����U@�!#\_md��v�$J�Z6r��IY�^�6�"�,h%J'��Tq�m���k�׽�6nrE�W���ϴ�|2z��x}��VX��h����3
>���{�/ ڝ�d���&�;�UH�A�BpCpKA�a_��/�>��ϗn�w�{�_/�VD�~NJ{@0qN�>^0�[��"��ꅦ	4����2�Yv0��å�@��C���ih'3!|W72�I�����T��SM���\S��3���bl� ����\��($�BF�%z\�0����m3�V-k9�I)�9	�Ő�[��'�ؔ�S�@������)���f�����[�vs�܎��/�><q��9���6} q�[ŗ����ܜ%�a"�s���Ӧ�e�_�#QO��SKbݝ���O�X=7j�aP�x^�����Otkq��L�P*N�厐�̜.��h����<�u��[�L��o&o��28z��Un7�:�%�����Ё˨�  ?Xp�ݗ�����c2��F��x���f����P�	ܞ��?ϙ"p��ZJe����æ̣*�hJՒ��f��F��)�U�ySY�q�怜=Eۮ���eQXh6�h�N�j=�e��z0f#Q&�Z36��FoLO�)w�GR�D���՗���O!~����qO�i�K� �����M��x���k�K�n��["7��e���`�����>Ո�S	�A���fY	�>~���,k�$���7��Z��WO��4?��`P���\/�Zߍ5R���{���mh5�!C�j���i��Aw�2;�%�C��0�q�BS�A�f��"���:Sxy��F87��:�ar�7*̋
�:B���(�d������_����k8�×YH`��<8��5��Js�a�Ɗ��� ��'��Z����:wj< ]�V�$q6�b@[�����Ie�a��+j��&~��ʹR59�u�J�ȋ�h5���z2$��#V��`mo���rҖ.!�Fz+�(98�r(�=3��l�ӟ��$�[�ڕ��MK
��"&]!�����Ǎ�h��!^�)3'�$r�7���(L�ܑ����GM�<���<��z������"����|w_.����A�SL��_��p���!1��ޟ�*f_nh�Ye�}���E/��U�L*�밗���2�\�,��@� �ř�k�bYq� ۂ���J�OqXj���D��ZA�>�L-�=Aa�C�\�_��{/@�Y�C8HsS?����I�!d #��>�tP��-��n_�$��EW�0�Ĥ����q1q|�Ҁ�~ϚX7��W���܇^�zs�y����hooq�]8�����$��E�s��o���zrr��Qg�52�4�\�f��ɵNb�����?:�,$�#���-��C��ě㈬��/�dN����[���XYeV�P��נ�B\ C�Z��L:̐Y��4��8���L�-3�?�N��Q �0���l5>�~5�����M��N��G����$$�P��ikU&]� ӁP+�44���hX��K^�L�&ۄ��������R�����RAf-D��ሡat��fO�z��ap��_�)tV��Q�q�"��R꣰�nr�\�Tu����j���I��t=��2�G�����"w���-�t��Ԛ�J��'�v�D$
����/1x�q�Ԕ�)�rM阌�ə���0G�q��$8�����Yn�H:F��J����� Y���-��R����t�U�t�_�������g��K^S��`�nUD�d���qOBu����q�S\�W��j����I3���D$r)�կJF,h��3�CN�2��)0�eG��K��n�|ќ.RF��wސ�:8��DI��g�u��h��a��o�8Tv��vyIӎrŧ}70��|�_:������m�ޔ�A���?�~��>� 7����qk�q8(Cr5���10I��h�QW}��p$��r?��ĭ\'��Cv�z�8��5h!��J紝 �PM�C�n�xZ���$5��[�R+�(����P�,Ԫ�s�J�f�@6�	��a�߅n�K/`u�P+\��'�Y$�ݕ���^��ݝbXV�T���J�� R��f��1�����s��|��o�~�:�5��T��9�A���Ǎ
\����ni�=��w}��M�P[�=]/'�0sFi���3�E����D�� rb� �a��c��[�y�ȕ��r�6i*R,d]�2�n�<��T�	��'1F�!�D��f �#��.)^$/�k$��sv-~�$;*�
�s��&��]7}!��������b��<�sy�����V�ʃ}`X�p�pҕx�uE�s�^������RJ7Sb����>#�(K*Yh�g���F �m���񃼍���
�K�m�� �`�A���;5(��xhAO�blH8���˾�H�������wX�M��/F�4�B�מ�$bk�������̕1��5o��F�<A�VY�Q����f�=�M!��&A������UL�/EԆ9�	�[�j��]3�.�V��	��(˵���n�Y�<A�k}���j##�𝭈BWHA9&S(!x
R��7��%Dl������7�Ʉ��v�<�/�un���_s	+�>C.'�XdX8%�F�)���B
I	��9=+F74j��xq���J���)<�Z�u$�(�;2ߵ�Zt%?���<�F���@��'�9�3�#����vh</t����	9�v0��<U�9��(Z�q�-�6�)^�m3I2��z�n��4������z��<?��fQaL�����k��㉢�N�3�d��@� a
/�)뿀c�
x���t���Z�ȍ��8'���" �r3B����G���i#
�-*=�o�JW�P�nj쟶�)TS�)�s�7袲����K��B�p�ӧ�!��#6���[M\#��o���l�]	�b,�������N]h�=j|����G?Dс� ��Z��8�,���d/�b$ug�X�FqQZ]���I�6apaY���G�ر��M�;���H��Ӄ��� ����>����'��\�)Q��/n�U�"�
J�����Mjyܬ����t8�:2����"�*J��I��@���L�JgmK*��nd]�3�5��At!��H������y�ɇ�$nr��j���P�Dӏ��N�@7�ǟ�͹t>2�;[ۿ�9�����.� �M�i�H�J���֍��*��X�_��*�%Oc�0�	���N+��i1^)�~g�,����7m`��g�������m��N�:�>���J��� P�1�d��G�,;����2i��ADdY��m^Ʋ�S�a���';�F�/#��%d^�0�ʥ�����1!�y��v���vl��ct�!��b�������t�w�ʂ�U5
����U�t6�s��U���᮱Hpk����r=�=4K!9�*4`p�ΎݧJ�40��?�2��2JU�����2�Ϝ�̽�\򫢚�����ԗ��.���3�6󛪐��t���Ԃ��F}%�� #���a�u��}���Bw,��?"�h��-�ȃ�/���c�
�N)���P���2����d����Y�E��fwԎ�U��u�42;�@>w� ����9|T+�?I���V��+|��<乎���RV���-���4o1�ʾkcD[�벘��]����DU3�I��=���
���*5�=���?�p�=4������0>/��WR��g�P!�~�Nl�}�jw_����y�����>�������Ѫ���hH�� j� �[3�=���'�Tt^7@њH�ZA��d`�u��;i|k�v6����uk��ƺVAܤI���1xn)*tg�;"W��P:�`%;{-YQ�����SЊ�3W!{�����f�.�������P�D��)�r�pz���d���U�����ƊЄ��?7d;�e��%�8)��_��B��m�Ck]�k��ύ��H:�d�����n���R�D���`Q: o��i`|/�2~yΠj��iI҆��IK� ��,�36�%)«N8�i>�cp~Y>K���V�����G�u㙧?��r�Gm�����6~M2G?��� 2;��+I�) ����6�C�<IB$`�8e�6g�����Ӄ����?�j��������)� ���4��C���}M�������!��[`�q��Jd��l	��	//�Y/����#Σ4]'�ѱ�45���.@G��9�G�����?UXt�J�Ф(h]�	��wh��7Ns�gQy�V T� ��g8�x�!�o�2���uJ���w%�M���\�W�������U���2_�0�_�{��}j�'x��WCO��f0|򱹙��"X���~�65~S��L�.#J\��sz��[P��K�,-��ZjZ�����q�/�$�+�{
F66�(�W�'�������h���j!��U��M]4<'ӌ�%$vH��f�t�x�L#E�	�:�߅h�F�r�+f:����2�QA�Wr�]i�	��[|$�����Ԫ�I�q(C�%�m���.@�a�`2�8�X���ԩ���Lxp�:���6��,]e��o�`78T!aI��vSE�"�����C�3=�wu�aBN�|0���:]g<�3�E`�c���Ǌ7*��N�A�]����v�6�f>�P��Sp�3����I�^�I�U�v�+�$�vh�&e/�dCc�ޙ�	�3�B@��n[o�	�LV<.���RzC9l��7J�m(�ގ*�ʦbI���l�g���'�]�%-����gH�|y��W�]���u$��)>�W[��3�/%��������,B�
yԑ_�_�����ؠ'Q(,���nS�@��KQ~a�0�B �Ļ߈0D�>a��Q�|$��V��\߸��_.wD��P��La"qk%)qNo ,��L�Y�@��0�J��CV��C���B��PW��u�^̸\�j����$�����̏B���#����E���V��D�����C�O��5��"�����y�Xʄ׿,c���Iq�,����t�m����K��wmN�kG���"X;N��0%��[ľ�~jG��\�W8%ѲBN�5�����7��d/��دN��k m�]7���z�i��p���?=��A���a��d(amD��y�q��kxyՒ[�;�`�1�v�(��� Z�����0گ+�����/����e�(�>�M7��Q�*��d?��w�3��Һ]f~��އ�wa�EqNZ;�oV�TS=g��R�<��%��49w͢DJa�u?�ă.�C��&�M�6�1��^ZFg=��${U6�X^"�0ƽX	�p!Y��>�N����m<���=�{�2���`f��0]L�f�j(W�	���!(;B���.uT���+��¢\�앢�oF���������0{�N)�#�
�����be} rd��b��`n����7��)�BG6.��fU���tk�b��k�V���Q�ṑ�m�vV 	#�Wb��Hb�T�	���l�guyW����Xt��4W�JY�m���ш�C�x�9P�v�Z� � [��t���S>K�&�7�Ԋ%�l����
�Xu�W�Gί\�c������sI�c]����:M�>�ɾw�̉�T. ����;�ڈ���#Fm��4�1�<���*����6�'�A�-�L����_ ���_��*f>'m.�6rr�J�%��{U�;�2*�f[l*�dK��u���^�mPΠׅ�����W��Hg�Y��8�vtjP	7B��#ދt�"o\������W Y%O�"�j��7.a=t����uO�,0#����dु�ő�Ԗ��짥 N�}1 p�/q��\DӾB-?�N�(���B+d�x���� ��� �M���5;a���OTP���	^/�sP��=�����>R�=!.���o����;-�
��#=�y��%�_4ۗ�u��_a�[ت�7�S44�&��w*>����ؔ�f�J!�d��\���
έ�{��
P�����O��'��"��eE�/֕�޻u�^���Y�f���W����i+���E��\&�Fi�2{�'p���3�u?u��q�_�d�����^�lxR� ( �n�9��c�E`��%x�/	TR�"~����撶��EEs�]\"m�e��w�L�?�F��v�a#<�p�P^n�L�����k@	o��/�<2,�n��,�c�[4��4RG���X�(�E&]pd�z����W��ʔ������Bt^N?��,�%S<��/�!ꈔ{"u�֑ZOG�jH�G3h��Wh(C�t��֢�z8d2�����|�i��������=i ��gF���v5�|�g� ���@�,�F�vby m5(���f�!�J������t��,+Tt��B�����Z���<$C�����wZ��߼(��70���md�A)Z���=nj�G�A�Z�}���6���\�mP���M������Ѧ6���|�;E�ǲXv�!�N�T�z�!�:�vNu$FE���AC�]s\�P��x".>�LL�Qr"Dk+�.�ˋHfN���9�B�Дj�w�-� 8o�����W��U�7�Si#����N�$!��89Mq��'�B�p���	�|vQ]i��e���_�Fye2_Wi|\�v:E"�Np?��zE���:UD�w�_z�c���^�].r%v\$_���#�hD�
$�)9,�
������]r��Y��ҫ*����B�i��_ܙO#��4$��PW������ƹq�	�Ȝ�g�$�)Vq�Q��v�_�o�t2��Y�)w$��C�}US5��%âD=b�.}z��],Xl����~X��2�����dcvUv�ٿ�`�"��8�E��E���p3��o�Q�� �W��r�Ѻ l��?�P�u7��k;%��X���qc5]�i�[5�B��ӆ�
� ��E�#�A�/K�6	����wB�����\G�5���0�l3���εZ(�+s�,P�zp����U}*�ЉDW��!�5�+���[�/ >�K�*������Xe���ux������$���.s/>�_M���I��:m�S��hx�k6򼽽�@���^s����¡6L�-��XUD�q;���뼰v޶�@
���r� z}�����5��Z���{Q��|�����ТB���GE���e�vZ�d0��b蝦@7�i�R���r&�~cp�6-�ߛ�9�u�ǆ��W�9�S��IDk�Ȑ��S��>hz��#2:���Ȉ�ǘ��������ܯ�Q��LE#<6~� �������� ���t-!�j�K��r�A�k���؄�ϲ��V<ZUNu�K�"��%,��9��,eW�5Ny+�1�% �j����<�bm϶4&<	Y�o+����^p��Q�pV
H�[𞤣pW(��;Q��yX
B�����J��x�-k^h�[���T�2R�m@1F�Ƀ2��yކ�7��| �M�+j�֚�o�4��1QyD��ad{��H�g�ش�Y���IW�vi|�ۯ㬽���s�~��HC	ޕ���\e�j�2�O���"_NI@����v�'��>f`(��^H������]��-��F� <:A�4YN �gZ����%X4��t��O�>�օ��X9����ZL@�T�T6h���wl���|1�%�VU�T� ��Q�t��������� ��rp�Ե~ ����/���N
��%�=�*x�٘�x�������f�w�RX�+:p��h���U�{%��I�O��|�#S�.\�%8ٖ�_��w��_Ię��)iڈ���񧩧�SX��Z��E.�)Q]v�)���MK�l�2�z�E[��r7��-Z��c8�����䮓�bdכ�1��	�]5M唪��\ޓ�ɾR*�n��y�v�2����5��#׋ˮ�\�&+�ߣ�v�H��.�l����sڌĵS�~<q���]�$�>wu�#\I.��~�<v�jZ{x<h4է��h��ڭ;�B�]8;q�G� r��KSƥ��%9ᒒe'q�jrG ����cE��\u;����{���l�am*���$�eW��8�_�>�C=�i���8މl[�T�W\ğ�(��=���=#]�m�{�\V�����s0� X���f�Br�����y�!,�F�[��(���:��F�_3������w���#uc�/;2�{
1���e)���:�4_���d��=�H,�BƉ�e݉2�a
5Z�5y9�t�'z�@!�m+�ץ� �ǔi�ɢ��<C,4w2W���s�������<���"�����ާ��~N=�Ly�:(JH���I?�Hl���쉂L$n��~�Y�}��,��}�_[p]I�;
�R@�a������T��8����,�"���dV��qF1~LW�3�[�����j���-O��:~��$��#��z^��G�y��p/�F̮)��B�U䐥z�ZL���%��i���`n��h5@���b�=����K"EP%n;ǱSӎWHtQ�K��vz?j�s��N~���!H'4I�`�oo�B{/�:B�N�}��U���ϖ�Ν@���{s��b��U�F�����!�zl��*O�$�wa�#�TL��'N��ˏ0ҁ(�\�u�Mo�\^��uvyU&����F� �V%�s׋ı�A`��Xu֡T�{���ϡ��{.�z���:�"c.�Z�Ĵ5:�l�t�nAŷ�x���S���Mpj׷v!��a�m�F�Ω�`Д�T�I��_�������\<K?���F9 �CɉC���4��r��HF
|��p#��*͊Cn�R�5%��?ۢy_9������ΟK��@�u�|8l����!Kǒ�7{�X Bnh#�#D��:�I�0��-I��ձw��((�G��q�6�S�CR������v�cgo������ԥ_gԥ� �5����*�c�a*؈r��HV���i�q�/lQ��L긮t��C�9v��O/��$ÉV���w�0�^���4`re��Q	-{�d�f!�j ��Ez�ҳ&zU��a�-J/�Q!�^��˚��[�^\��)��'�Ί0c9�r B���/X�Jl9c�sW�)yGi�uw���b�*�����QX�]#��lp�&	� ��Q��"ߗZhl}���_���Y��Č��a�P����ל���$�%G�a%"���J�)�?�Ǹ�x2:Ͻ�v�y:�`���BO� Z|v ���~�n5|�o�v��/a�t�M-.��;�?I��տ/�+�ɷA �7;�|k;b��2�_�ې�R:M3�@��!�I�س����9��\���QA)[�����>o��e����o���%�X����[&Q)O�0��R��m�MT	����q�_���,�0=����2A�W�bй���<� 3�J\I�E���0��.g -�K��� 1{Dd*ª�����U⸲�B��DW\J7)w�ogB�t�$�t��U��;�`�8X�:��!�u;�\��#�J�����W&�xL\	:Wu7V��z��9���a��qo���+�"��F��!��/���T�����5��0�$?�E.�/R򑺿���V��8�N7��qc��H�����6bV�/�b���)OtI|��c���f!1����-T�9��K�-꺛�%���E�zt�{Y�?�+��1�ԣfb\�Ħ�i����͇iQ�=?Z(0}������p�Ys���h!�R? I9����boLe8�i�v2��]���
\�r��/x|�����u���w'���٭̾*�Z�:uګ]ct!FhB�?��	6WF�׹���z���V�sw�}N��R���_��Q���ޚN����j�m�|�o��h?�s�T������Aa7�#������Ǣ@N����Jr���]ܲCz�?���P�����J��3}Hf��u���o����'���X"�@y�؞OX��ͣ��c����'�N�E���le:�ک���`�G�f&qe�YK)�eYx���R��̍�s����#X�|�N�6�ɲ��_N~"E�+y�F��|0'��(��b�`ԩ��*��T1 ���=��A�Re��!�;i|���S9�`��rb��p���4OKς���ИM��ExJ�Q�Ԛ�"��P�Do��|��M�����2 =[����$\Ю�(M.@�O4���xC	��t�{�<�u��.Gو�X�s�x���'�e���aKZ���B�"]�l��IU'�JJN
�c��%����n�dj�Mtg�!�?%�2�/S,N'�����V���9�`��#�u~�]��§_��#bړ K���B��f$�m4`��/n�H�7]�`N��q�!H����i��������A��"�LX�#4��:?F�@0������!Y�bu4k���ݗi���$���ق����C��X����s��x� ���~QA�Gc���Eb�w���1�M�c��A��)H����-dK�V�
�ir4Se�S�n?�� t���erQ��#E�J��{R�񝓐����>��נU��[&W�4&��� Jʸ/8�SS��|N�m�Ը��\�;W#���_��i�3�G�\o���v���޵�u��*��T�v!|�yZQ�*��*�[��Ц�/Q�m���$��W�K�0�����t������C��>�3�<"�[�j,��x�:��]��1�W�4�$Ө>�"9-(�� ���$4�1Q���s��!q�.� �@�tX,Nrl�l���⭝D1HW�-^P�*G�.�=�f��N��8!:���x�eZ��s�����j�2↰��
\�
�{����|�$P)+tVMh����Ǆ��[�ZP�`��0�
��U��Bo�q���.M�w�w�x�,�!�.�i���[H���,�O�å㤇�;�ڟ��s�<|�jnN� [G(�T9�/���$깇���L�*�yF�s����/4Tܛ��&/ݪr�`�vH��n��P�Qz��/�2�'n6dʐy3sa?��:������)���1I�tӌ��-&�i�q$�C��zV�i79?��9�M��5�klQط�m�E�^f��ͻ�EQ!�0�A㦱%KH%��22�G�g���;�K瓓`��v�S;�K��l��l�!{����N
6R;�\}�U�����5�r�e����gС�X�+� ziumU�do�`��5�A�:�~v��1rN�I��߶�A�>����o4��jZ}��e�c!dC!u��b_bhT:X=����� ����Y�J���
��ϧ��̓?$�5-+d j�W�e�0Κ���ժ�Q��96hn��۽ױ���,��TH����t��n�/9:�p��8�����T�A�Z�Hs|�;|�:\�:��ex���M��N�}PM�|�Rs���5B���^B��ÜC��	�:�6ŭ{�ݚ�f�����.^R��u,�t6��UQ�I�>5��D_:t�����6�!q��-űҧ�x��_tQ��Ӓy ��h��T���C���I�<�7��̓�$g�tz�U��x1PP��2Y�JP{����[��)܀�٩(	l�y[�h��έ_���i���e�:iLD# �M�֑n6
��fV�1`�|�)�a��+K,��V�-�s�Kj����\}����Ԥ���`��!�z/V
�����&������?��T���h]�͵MG��ғ!�XA%�f���5��P�I`�2�Z�ِ4�jN`ü��-��aL#�fx�DS��B>`�y���� �3a��Mb�q������d�Aa�ש�fVޟ�uY0����#�d�8�+�.Q�fq�nP�WH^�՞��'��C�Y�c�sE�8���yaӔ��L�fkRmYt���C�f�?���S��5o}��$u�9 ��� �����I��HE�[O��y�֢" ��{�H��:�:�CB�H�S�;�n�w�p'�G�d�iF��Ĥ��׏�|��!�.:�A��b(��!<ҥ��>5�#��p�%���t[4�o��F
�7aàф(�zTb�����t�3@	!�?�-Xk+�v7C1۔?i6�6�vZ~J{y4���:O�	U�B�7���7��V~�Ƭ�Bk�ޗ���~IG$i ��}X��T.~��rߦk� *��lq6�����C�ڗ��|oV@�����z���b	$h��IrXoMr� �����Y4-SB�sRqJ3���;NI�huċWƞ��K��n�.9��Ϣf����0 �_��HcOb�fm�2�2FU�&��0��ZSY��W�(���?��Y/��K67PU�@p����{	�T3۽y��P��j���B�r�U)�:�M�מ��������ܔ�+!%9�
$:�˄͞y!�6��P�4����9k��邋LL*z���k������%h������!;9��,X�3d�0d�;��B�,�����ʒ�{��h:3!Lؑ�̎��������~m�y����	���N?yBڔ*��з<m��;�f��-�W{d��H�$S.��U�Տ�vc<H���U���-+If }���>J%�(C�a��K�<k���7�y<A�]3�k'�~�rk���xg�%M0� ^@w#�)6�����Y���
��&�h�pb�����whs"{��~w~2��Є��{�1�h5 ���Ȓ�}�cb���&z�k�F�Y��x������vV���7̯�,<���QE�Q�s��RI��t X���zD��r�82o��8z�}2W����"%`n��F��r�����y�cJq����ж3(���B*��d[�;ppD�o/e��g�����am�� T�R�㞐�ɭ�)����g�g��Q�U�l�,�,f$n�7Zj� r��,8k��~��L�.�IӅ�
z��v��d��<��b�vq%uܤ��P�?�Β2m{Ah��d\�L�˪���ʧ�����˒���8{ '>Q$/U�t�����O�٪��żgB[W�q=� �ا�[��reb�"��;~�4��ޖ��8����X�u�m��h�V�3s�Ȟ�̨��(�l���2� ��WP#�,L8S{�aK�fVR����e����:}F�[��y3h����rQx�)��R�1�4���{��pҊZU}\'l�d�h�Cח���G�G!�n���sS�VS�;/���%��_�	�1,>��v���h2~���u�L�h�Ziê��oqE?q��H,L�~G�'�[/4�n���o���J��I����v>/�nzep������a����c��-��Oj1��yaNm�%�0 Y%o�7��1���LK[E���3�Z�O���35dM��OQ��ȟ[�z�?�ǬZi^��ڌԫ���߭1�5�NC�t����f�?���7D�N�v�$�|�yUS`�U�f���T׵N� [����ō
���9�ǅ9.�F U[�X�D�A\=�Gw1����]�dc������re&o��J�LM�'�,�!��p��	.�ofጽl^�(��^a�$�5+�c��;.��~�a&D��u��,��Ռ�#W� �|O�R�f��z3�������y�,:�n�ӟ~_Fk�u���Q$@s �(�+�A`������1)X[�س��ݛ������C~��eJ�('�c�����) 3U�Ub������?��lj$�VߐLs���VU�����𠺀��+L@hȸ���</�Ͱ��u�6�9�~Ny��� ����&7��r��]���K��$�b�X}���Ъ�O�2>�W�$[��ÛYw�v���>'��kz
0��o��S�c�+qc�fxi��3�ظ��IZM���0��R/��"��#`�3�(88��@�i�JN4}��B|�b�%���7uB��Z�IR��Xʐ*�\~��~7S�8<���O�ő*����t �^��$˓7�0��?s��8�f�7��XճO!��L�� ���26��v!ˏ���s��1�2�A	g��g�_)6N�LB_�F~�o�5P��T0��9�hx�[�Z�M. }�=(t���ш��h��!�m�j$ԩ#a��$�4����B�6ݰK�FK:���u��ڀ���B�
�m��!��e���4m|T%��&��O9��6����/f9��i�"��c�A���P��5\�n�~�K3dś�Z�	rI���;)t��rPt]�>�:�g9+.;����F�VF���/�)4�|q��	H�]�p��6�����PZw/D4�f��[���WO���A쿲_L�� ��S�3��{O5D��i����>���IH[�4��ɖg�n�k P��߁@5���?26G����wm��d��{>�űhw ��_SD���|Y%%�)�K�䳕!�#Qt��>#��O{"l^�}�X�N,hL�� x6�tm��C��������#��(�l��c���T�O�%�6���ီEsC~�`���k�Fmݺq��j�BI^8V�ҟ������w�F��W?2ʏ�~�ϣ��Z�b"��;�&�8U�B}%v����1���T��!_E��!�R�g�I��[ܡ�YW-���|��;)c��b�͗���\V5.�~�r�ĘTϘ���J�1�
pb�ȇ��
K�����V�a��}��!��.b�k�aV�l��5uq����t�3,��&`��k��{b�%T��z��6��F��c3�.D��$�edI	Ap�'�Ы)ڎ�T){�����K�H'	��ʇh��+J�3�����c�E��P���ҍ�x��Gs������ϑ��S=�F����~8~��.�S�Ѿ��N�>��=������x��˙}-�f"�~�{��F%싊__*>C���y�?G,RslCo�89�~�M+V�s�_��6�&�3�f�0L�P�,H�A��-����O���.���W勩�{�y�CU�^��*�jL�o37-Yu�Y�f��4F�~����~��R��65�T!�JBƏM�QB%+�GK�l^�dt+�-=�{���Ȁ��Z7�(� ��B~����q��ǵ��o�g�P����Wx"�HNRP�֞k>�B��h2�ڪNh�E��D;B�P%91���ڤ<M�P�LHL�0u�;�����v_��P�daȪ��Mq{�5�u�X���;���*0�@4T�|V������g��'G:��D�ҕq}%�`.�� ��7�7F}e���z{�o���# �4c�aMXH?������OZ�ZZeǅ����#���(�I3���kF��f`��(M��A��&�YP���A
�\���;0���Q]��^�[t�^c�V�>7j����K�j�hf��(t�F3�	fX� v�NHք�)�Te��S&��K}��bz�]��N⑳j3Q�N�.�C�>i��୉m?5#pZ{s�K���5�sN�r����B�{�mm�HFd�a��TH�o~�i�}m�_A�!:�^г��{���-�����B* ����|^>aJ_���� �VׄD�7@�fvɛ'��>WZ?�p���+�k�,aaZ)��eU(�Լ�nO�,�b���E�s��I��(yئ\�����x���OKg9���6����Ĕ����V`W�U��ֱp&~�1��n;vT)u���M��7� |�8\��>Ъ��6�{��0M�5�k�>�^a�m�\�>�( JS��2d/����f� Ы]�(��|Y�犌�Ta�;awzNW�.C%˞a��<�a�:�����l����Xa�7�d0�?7�g0C�$J�2X]�u�!d�X ���iꀔ�M�J�Pg�7�Gf��އN��Xd�(�I֑Li4�0dA��!E�J�������Ȑ+�Y+�u`�DQ��]��L�!n�^Q�-�A[)/�k�����c�YLY|�`���o�H�F��QQ�����6.9Kp��}�­�/�v2*�D���&��-����5�z81)�ކ�l19�{7Q�Ct��� Д�#f���`+�k[B�c���uA.a�J����y���-��G	�D	O�����ѽ�ڕ�H'�Un�ɔ(��`͒7ݸ��Ϝ�tg��	�*�_�7ν"�0 ����8�LN$f���'ϱ�PY4'Ǌ�̇|�f��YI�'e���n3��a]�4�xm�����+�7}���D�B;R�����7���`��P�aU���(U�"|U�
$C�U�!j��~U�An4�7:P�Ԙ	�ޚ؁�cs�v�܇12��g��7��y�쿎��U�pm�����t�#����L&�Ut#K.c���\�t���)t:��3�G�����gf0Vܰj�-���x[c���_X��b9������YG>,�?MW�8�<�$=Ʊճ���g��&�ڌ�[�nQ�+��WZ&�ϳ�o�RwM��O�zLL)=���>I��f�o�s,`�$��G.�%Ġ�5�#�R#���娔���	zw����R՘�ٞy�Է
�t-rY�{W"���`�ꇐe]sZnM_A���M��?)� ���q�R<%l�����j^�w֗{�etCY�~D�F�.�̸FrUIxR=sY��-!�#��ϔ������0���<�j-��?��#����	.�7
�[�r����J9����l�u]��Y��������6z����152�G\=P'm�!Oۡϛ��!eMq�r�|�c�(���-]�����+���T��	�:��~Y��;	�L�>�8!]k�yC�c�gJȉ��Iw �`T��
)+γ�W�5G�x���ً��3�y����_"8��;S��B�q?��ᐙ����}���<VAO��;��n�r���_�Q�A�6�-{���-S�`��Q�u����'��tz�~���*᥮����� 7�F�b>J���j�&�~��rIc;�2�*˿Xk�3���c߂)z ���l�����M,�AK�3i��ɛ\곖[���8q�/�J\�/�y���׼����7'R>]��j	i�#���p�@E�)'Wu	Β�����P�=V��u9	t��=�f��`ɖzf�虝��x}~�F��r���G*�ݹqZFp�K�.����7��c��AG�~����b�d�g��1�� ���ʕS0T���@���T�a�~� �̆�������0e�X{a���~uzH> B#f�=~��t�T�63��%�o�~}�2C�b�C�et%�Ǭ�f���*AΆ�������N�'���S�2m~(�V=�X�����TL!�U>8�=�,��H5l5�O\�.��m2�my":�ջ����ϓ��2�z�GЁ�Bݗ��@J�H.U�FP�  p�sY�vFF�e4�	��3�˲�o
#�y!o�
��� ���扦i����@�5��W[g��QEZn��h��q0��I��*�X��}�����v��t�-qN��5���x��L#༜��q�v;��	�k��O��1.v��p^��s��%�4���\�7�?�Ḻ��G�Z�,�� �Ў:Im�µe����}�j� G����s;�c�4jU��Km��j1�؂z��`��p	q�$?��� )6�����G�{F��Ϻ��h��&�;s��#:'^�-V�z.<P�G��qaI�fƭħ����T,�p��5b�+"w�fc�wW�xc�P	l�fr�Cf�[�EE�)g��6�S�-��D��M�7L4lp[�WZ���'z�ze�>����(d0�����2*�����/$ߚ��#/a3j�ތ�q����zx�dH�*��G�;��,�x�� +��[M,A���:ic�!S[D�YF+g¼ p�H��nq��#��'�~�D_̘$�x���5&��Ϯ9��Q��\`�̟�DA�J���[D7ǉR�y��^����X���=Չ�P�K{<��#�>�EC#~Q�[��߇p-_~���,9��1V�.
�N	~d���yҝ~z*��4"T���˖^b�>j�A+����9C&&����-���0\�֏��Bv�fc��d�yׂ��F ����XQi�;#��0s(G�z2�o7
���}����\�j[3�P7ݧ,?&%��W&HC+I�(���M�O)��|�C�1���٦j���#�4�B�F�ԧ�x���P�:��/�9C�� e�}�m�[%8�ފ�mX
xS��Z���I�P���x$����e�� ���h�d%
9������ڋA^#�jN��"QK*A�~�,b�s�N�d�-�%��械2W��x�;���XV0a@F�$�~��gAx��Ğ�;	IJc�'��W���}Z�o�T@;�v]+ۀ�����r��}~y�f+f�7�S��Hq�b�����ȸ����0�o1c�H"{���3��z�p�����ɕ�ٶ�o�i��ƒ�4SC���#}�U���m�S6ժ��{��ۂ-JƄP�1S�Ku���"
�7o��' �@4���
��X�5Y�I�G�c�K��ڔ��~������x�v��O�mJ�j,j���J�Ϊ&�-�ZD :#YX�c�nS�
3!��Ze��E ���h���ҷ������2&�ؘ���;���(��2��0Ʈ=q5�P%v�U+��hfK��ۊ�O��S�D�xxD��!p)m;�ٿ����0�*A�6�B��Q���M�C����J{D~����\0��c��Y"`j��8X�K4�),=�h�%u�,b�a�m�����NvvZ�R\�F߷c�PQ�~?��1��,p�a���G���ae��"/!���%��P��r	 �j�^GvƔԕ��"j�����^'{bd@9�K�l\����(~�N�ͨG��O��%���/˰.��K\FI�g�k~��Y������͙L���>��]�'֛dky�FP����B��}bӔb��3YL��e�%`t4�V��%���аen�h(_��i(Φt <�C��W����g�	� =o6�N��5�et`.ۯ�m�����0��B��6�s��
i�⼪�]��u9�,���Q���غe���J�˱�p9,E<Ҿ�n�4��C��	��O��
�[�yme<�0�b��_8��ϔ0t��5U��#���gz!d-h7<��>�����HEZ}Q��|�IJs��h$�B�� |�M�5`)%y[���۰��}�S��:�����+��\�+�~4�:/@"�F<R{�N���;K�OL�#]-e���x.b���/'0U\�U�v"g���r9�UmT�N6�F��y��qZ�	R;� ���#��1e���tּN]�ZӷpZ��[5�8A��%�}�$gB$u�|yҴf�~��`SH���Y�]V�B)D=��g��K4��O�ޗ�i��4�5�����-�AYsU{���ŋ,�%�fP�2��b�ϴ��@n�Puߘ�F�X���y��>� �L��^��;
B,4��}�R����n�_�GRS�,��ht��)��m�0�$�`�%��]���U+i$�u��������|��u�i���M�Ȼ���B�f,uj|��a�R��0? �Zr�N�x(/'���,w�,>��Ҹ�Z0a�i'��s��I���:��N�l�C���Fr��Qs����VksaY��@=�#f��4�i�qX:�\��ɉ#�#���OG�ќ����z�̄]w����(C\����yֱ�@:>��HA��* wkVU�x��Ū&�Дw��4:�{/X:�X��"���(�K�T�"M=��!��řB͎����4���`(�B��p��	�!✻�&+ٚ!ZM�����X�5�{e-�8�VX����g�OR��U&᣺�y�x̞�Z��i����?��+�~�1K�0�%8Duj�'t���r��*1���⻓�E�Ȥ\��`zw�����,Y���Lʚ$�������hg��ct��zW�ġ�����'V�����&��̮�'=�����-0U�
�(�n��ՋUmD�8���D�-��S�/R@K�D�zC�z�n�5�TY�Z[��2<Q�ڮԳg-�I�
٪j��e[���-as��F|�V�x�q��VI%I���j�w�s5���g"�v\>iih���2�h���`�w�1�"�`��nH�:�P#� etb�1�%�[��'��!�h
0�N;i�(vz�>WqH���l���ϫf�{����Թ��A);]�	n�,��Dm/��Ն��!�0��躉�jm`�c�&g.$Xϒ�e.R<��v��BG	���]�ʮ�+���V]e؞ 3ن�{��i��H5;5��������$uC�v����Np�qC"���g���0�s�|���9�R�Q�o��]d?s���ǜ�i��?���W���8��{v��Q��s���؀w�(��k3��.m���g���?Q]T}�R���ɭW��u�!�A�Lڍ�8�����5�l���"�ȕ��f�G\�D��%c0?�d��:��P��q#��׏`�A{�o�ae9��;����pP��)/@��is+�*nG/�갢�L��C2Z�Q���c�g!�sYC4�=�Z�}�QH�L����������e�i >����!áb�W�T��Ē��>�/	k�?f��@B�"N~xߖϸ3����w�X�.'��S�	���,�7�ơb䕌R�m��$�h�`�_r�A�^0nt6���i w]hI�O�@ xQg��%C9���k�[�M�ͮ;lh�c�6i�0�����R���#��k�9tps��<=Ac-GC�Ke��,�����Xm@��d�z%��P�|i�Mi�x<S���C��(���*~�Jiٝӂ��*��#/��:�
�Jr�a��ZWχR^f�·��";9��J��@1����
e�b5�h���$;�W��=��P�7j��eH�Q�+���A�7"0���p�Z��z���� /.e��(�r��z�~�ۤ�g_�$7RO��Ə��(L�)�9L[ �l4���]p{���-݀�r����p�;��1tim�������WD�JH��E����u���BJy��k:�Ez�mq��}�*dcsOM4�|��n^BFQ��/�� k�����bƖ�b���bb˥eOy��.����PӨr�A	H�	��О�ߎ���_��Z��R��:�!]�;~Z�0�"�K����a���ƌͬDi>��7�7��-�k� � �NFyV�"MԼ���z�#'��M�J�'�.����c-uhWء�8Ƃ�z��v�Γ�A&�c�9����	��d��ҖU�Wz� ��3���"�؉�Ul_�5Q�蠢�Ł���Q�7���JJ3� O�+N�����@;����$X9'U���#����F)�=c
�_	b�<�̨Xv�
OyA ��x��
��,� M{w����i�,�Fl!�'2����u��-�,��ϛ��atw�y�������6D�ͪګ�����l�/�"�x�������^�z�S�|59i�K�%�9lGA��Z6����pw��)��`��{Q���˪w?.���ä�b��'Z�Sv��9S<�?~Y�EX��-jrg�V�A,I����D<*ːOCd����+C���{�Gt�d�g}���c�k�bDQ��0��K�Z�
j�ln���J��h<� ��×Z�#\r� 8�Z�c'Lς���84�_���.]����TY���N���?8�NH�Sw�p�+�3���=��vT*���.	���W�lTWW{ lo� K�[}�'�U Y*
�=$�Z�Wv�Y
�]�u�� �ӄ#u )�I�sn����k�
ZǺۺ�0'�ÿ�s�����ަ�0?y�JsK�M��ୋd����/R��l��P���B�gV�f-�����%��NR�My�����3��{C"�z�%UI:M�i�O&��=i��q���l�F=���%�b���Y3 n�p)��f�t��H�P|zj��\Mݻ�$"RPuf�.;�,KpR�3s����+b6a���3؆.MEHː#�Z!��S�Πy_�V�=��ѣޏ�n��s��I��p�J�a�b��/t�N7Y�^0�[�8k��}��#^c��o1��G�����	�><�p����_J�İȆ `K�+\[�_/,��e-�r�#��/Y#�~xNf"ވ>#i�[]�ZY?Ǐ?�����e#CRh��g)=�P  3h�~�)I�/%1�$��8��7���)��G�	WF�+P�L��U�oџ���e5� �RL`2�B�KjԖ`�A[��\z����uY�rR���]�r�n#�F���7��[r����X�0�E�vĻʥ�|���C�po��%J�n5�����x����\����9��	a��#Fd7�R����z�\�7�Jy�Y�F��Fp���n�p���������*�R!��p��΋��ngz�A�-�R��,���ͬ��Bu�T޽mD��Z�\VP*��ޢ�_2�ƽ`�������TYW��^�Y\�n ��!m���U�P+`ێ���Y����3TP�����i0�,Y�� ��&�������o�|�h-Vl��a^��O\�#9�'�?Xo�3�EM8̾c�]) ��詽=K����؞��u���`|���[����������>�����`d���!�uc>�`x�S��r��<�?#Ӌde���E�x/"G��@�� �h>��C�iq���et��y���{�B��c}زwIŕ)}<����DO�����ֆP� 8���|/�߮��Z6�J�D�|��٫h����F��
�0}��J����K"u��C�X\��CvUl�M�+�6�JF_	<������h:�l�T��T

�We������bU}���L!T�ߋyգ�5���وNƭ[F�zKgW��Z@۽<Zھ�e�*i�೐��,����%��9���w4�C��aZv`yR��q��Vn����4B��L����=*�s;%�NI޷_"_Es�e�Kӎ�)�~L#��2��~2��h�h]���)~�cc�K\m_����k`>�c.2GcZ�	�;7�H<����B_y��E.�yQb��C��FD�^�c��*��X�,��Z�jX�~q���.�#�w*��a�
x�I�/c���C���L<��"��V>RyC3g#�U�z�E)�k�`���EH?ymL!�T�}u���z[k��;�,�B�e�݆�z�����eL�P��=����|S�܂@"-�L=o^� �)�P>���N�����f,��~1��x���"�"���>����<�k^��Q8�9���]��|V_����c>K�߶�峆��v��(��|�����Ji-���Q�r���&�u:2֒������7Z&���a�j�D���4�N)?>)頙�Lw�8}��[N�<��B��v5! ����s�#�tFG7���9�����[�5Yw�A���-͢Q�S��}���/!��i�XpH����Trz�>]������f���]!��v�%K��^�(�/i��,��*>ʧ�'��{��?�����g�瑹@��Zk�d���zĝ{��R�dr�@T9���J�ըL���^pЫ
�E��W�sf�S�;�4Y!��QN��ҫ^̇�nͦm�|嘳��L�*�H�����y9�>��7��T� �z�rSY-�G�U�X����R9��o�Dj`Qw�gŔ�=������=�K:�M����4i�z��L��w���h�s8�y��	H~���N���/��B�W�,��Fs�6�d�����ٚl�,D�r�����'~d�d�9 ���6�7ʬ�4� �PIw����DoQ�H*?�#��S���Tz�{�X���ڝ�.:���n\lyҟ�_M��:e��;�&����p��n�X��qG��	�<�$\b�4ڝ���m
7���{U��Ʒ������Z�+d�4��I�a�<�~�(�q73��;�ں0�8
Gy�"l�3Tg�C��^��ۂ��y��r�u�F4��⌇��:�����O�
J *����\(��m�tH��?�p��9�u����_�n�2N�ue%�`�m4
�Ҷ���Z'`�֔40+D{E��v�J�m�qM����F0E�B��i_�I^��9caOR�V��U�����}��Q�R�{��ZD0�N������)@VYy�E,@��T�݃��C��H ��7_���e����݁�gn�`  �#/`Owz�Ph�Zc��ab����R��o���+���%��Bhu�S/����a�>C2��V�(��ߑ�0v[�y�߅�'�̥��f&�4�qʬ۞R&)���L���f�6���e~W�Uj7��B�ǌe#]��.fY���˔������$��؟����e	�]
wъ@��0g��H����d\���6��|hK��YU��x�Z����dʠf����4��8��[c,jr5T0d|���ح�t���`�b�vA�xl,^�0�zn�"����i�=��=l� �.�2�K���C��$k��q��B���D�9��<����؏�1��1�f2v��R���w�\R�B�"�1�۽?~�`�����>^s@�;�W�{����l�+�Z,԰y�%8.�(������t+�����ڷ.ŭ\Lw<���w ���B�n�1�~���\�<Z��������Ȟ�=��nx�k�"�y6 ��3!���{9�6J�I$ɩ��o2����B�Sk��l�}}�BE�Lc��n���� �t�0�
��.6�]�����9h=�����b�-��t](ܕ����U�ca�������2��b���k�+���I�X�Yۓ��sz� �W��w�8&�`j~#�.� ��6���_��y���T}4m���F��qlX���n�G��H�ѥ���՘�o�ǈ��Q&���O�����,�\�U��"j��v��i ��F�I4rd�G%E���wsWd�9T�3�W�:��~�!������/�_oEŰ�!��:Jho�O|N�Ψ>پө��&�5P��#y�_��W�ӇV��ZKإ^NcI[�ϖ�m�f��@��`�[��֊NĪQ�͵�،z{���Z��Z���y��HgJC�2	x��cl��������9���ͽ�k�Q��$L1[�'-%��y��e�����z��Z��������u��1���8f��?s���!��lɘ�7���*�)(#u�;����{�Oo�7��Q(0'F�&$�����W��N��`����j*���{��� �p@�l�`�7c�M3��>�P��m`�QF�����bdkYGп�n��G��VR�O����>]�'�43ͲR9���#[=w��I������&)&�f�]��{���Β�;21W#�'��%( j���~�[	
2����"��KFC?
�+1�*(�\�Y��/�V(��5�l�O:Z� � �����'R� �y��	�R | l��F�K[^��S8�%�y(|ƮN���ql�¬ZІ��<��qFt@��� @"N�k���y�Ьˈ��q�'T�r֢ t�.}V��|�j�^�x���;�9o$j��^�IN�~���T;�;�����Й��5�[�T8bFz8��4vD��%�;J��,����F��<?x�>�\8s&������Bf� <�-��q<�l��-<30��Z���4�?����tK;��&�֝=��R�8B��=M��~)��T�Q��n}zHY��LhL����G�_�`�s�\:��њ�ޟv	���B�'�n���l8������T�s�1�]���������'�����+���cA�Aߚ���	�;�Qq�����2bA�I��ZJrwF�"D�d��� �.$$8�9(���k���������û����bm����D{@s&�eB�U�~U���qXv����E�&�U�T��A��9>xfa��ӥ���+4�n�x;��� ֤��
=�2�=q�H�`�H�9�ߤ��ԍ+�3.�\��("@E]l)�Z�8��V�oJ{�9E���6 G+qĿe�bH�P����}��N�Ӱ�<I���]��l	֞]�%q�Ϫ�<�@Oy��XiX��gW)�DU+<��?�W>#�nԆ�7`����d����c�iU�R7�%�#+�[w,��&�7�r���2��5`O|c����ގ2�)5x�fn&36G&���I�|���,�Y<�:�@3f���.�=�6�4�l��M�t:����I�t0��s(#�2hL���_��lmsʒIg���*#%��<��n�4"�M�p�m���!��@�ŀ�;ZC�L�8��
5+K�Ln�p��5�TV[���[���1�_�Y)ϝ�V��Y���q�����{����)0h��RG��~��ӓxeԍI�麱QO��i%%9�C��qF��A�4�>����G�⮻�����w?ڳZ[�zgx��?�Ia
���g�V}"/�@8�������U�MT�[@)BHn�
G����%�gp�Ѹ2D�h}�l^��aE�w��~�n��cE�\2�ʋ�$��HDnw������g	V��^C]�7�Ho�`ʩNB���%f(���˖��ٔ%J�S4�Jdϯ���~�v�� ���(q�y��h�y|��F/҈��(��*#�����m(~�&��8	��t�0�\�`\(����K[�m~����������)�����N���+[_�SNj	�.ڱ13g���Zw�����c��yȌ�2*�
�+��ۚ=:���F�Lo� ����5�z+<��C������+Ro����4Z�F��4]���mS/_���`4m{�7�B��C��0�t%�0��$6=6ܗfJ	3�'�rv��'%��Ƴ��eIT:+�%��h`q��N�V�\1� ,\���"���ܝX��������Φ�/���[���K�B�+�
�W��T��L���?sчmx��/����W.R���-�2��yB��-~\�Ak��a�C�qhp��:�;�A�'��!����Y���4�`^�����H�HټO�gǡg@�e��b���!Y��} e�/��g�a�����(2�U�ϼɮ���PD��|�70pmX�<1P��Jil^���}�O��H�r��w��E��#]�;��|�5�8=��zI�Y(8���mo�:.k2qXo)�5��� c_Z��'����^V"gn�*�OYS�[����.G�D����͆M{Ay�l^3�|�0l��zP�1�5���&��
�<,ۖ�'$�����I�����F"{�e0�K'd'� ƵRe��k9�3Ԯ���c_����C��b;
x�b��47��9*'�0�g_C�6�![�VA9�FP��\M�6�n����&c6���NNC>_���[O��m����߈�ug�%#[��e�����$�U@ջr��M��J�o+���`l;o�Wߜ�hļ��?��%&�7x��r��Sz�vN����f�H�R��I��B����L4�w�D�;�^~�7�O��K�{��_���;gNY�s��J��z�)q�( �P��ՒpW�(h�U��ǰ`���{M��� ��1���Xz�&��<T����j�"C$���+
��zC�׫���8ۚ��?�M��o{R��T������8�?2�/�0bIb9\u��K�N*�t�M5�.\�0U˫,?���������e���ٻ����������n�V��y9�G�.Ϯ(���]0Z �\5q�&���l����k�{�2�@Ջ�#�=.�1��cRҲ⊟\�;S�\�ZD�����}�3�%Jb���^���׏�Y#m7vE����_'+. �~D��gh� ot��[�k���! �b���%���H��srk� l*��AҲ��jO�ݰl�\��9�,l��f*�N!���q��-�l�	��Ϣ��w=�H����ye�\�٫؞�������8�BM̦[�nT�[[cN,���:�)��(�C~�{�3�h�/�Br�k��&��(]��U�n�����-fcN��Pp_��4��CkJ,��Wa�� �M�]��h5*���+6X�aI�E
Z�����]%��^q.��]g>c�s�N�+��RS���r:8<�9�%`a���<m��k+*�Ά�45G�s�54�Sw�y�I鯪/ƀ�G��i��K-1�sʱ���-�_PO��a[�(�����2���'L{�ҏ��^kCua�p��Dɳ�{@��`����`��Tz$=���n�z�cp��=
����Q�D����T:�����tK��� �7�Q�?;�w;�H��8�̽���zh�9Ã� 7MG��g�'��LX�j�R��U��t�������'��n�y즙̚Ȁ7F������,��Q�7�ؘ�{μc�8��o�T���?w�N���;*��ƌ��W���U1B�:�͑u�XlBM ��2����#ޤ^��Px��_чƇy-:��4��>��ڛ�"�nc�T�"�tE�haj5Cݔ�̈O��?��e�&%�k���ʠ �y�)�'=�kѳ�m*��.�;��~xi�Fg;C�q�xJm�p#d�{���{2�2�zO����o$��;�n�%.q�(u۵�g���}�V��1Gg-�XB���|Ӥ�iÅK��X�>݊I#�nX�x$}�A�ܞ�j*��A
��D��&�c3#aЋ��%�p���n���i��!揬���EV��S%���,g�!
���q���W�b |8��H��K{�%:ڨ0�i�s3`��Ӥ�W�ķʪ��F4���	<�����⚄���-���޸����q�]:��ކ���#@9}u�
��;#�reF�7lE]`%��.�����SD���<�6�X��"�z��f]E���L��z��1����C0L�(y��r��hx��b��ڸ�>o�y��"�O�ĸ�-��/-�s�$a�d�4�/��;$I��|	�"H-�%Zga
m!\dGԛ����Ӻ<�B���W$��=���@4�&�]F�B � ��My�S�{��^��ɋ�u�)��s�R���2l���A�V*��"u�7,�p����+�ly*� �Uq$jʶG}k���6�<&?a��;E��kA���&uJԈpF���c�
d�w��a����Χᄿ&��	ĢH��� _3Q)����i�B��w�R6	OwF~�y!lޏRO����w�8py3���^rCauE�ܧ�9_�_��Pe���įF�C�%���0�ν	�x��EV:z�*ڒ�󪾌�74��~�7�#�q[��9Y|�5��ģ�1k��ׅ���g���<���R�Y���*@~�������O�o���h�P��E=�y��G�.�͛ZSe�}���2�E�E�s�]+>G!iB�T�G�P^�`rͦƘ���A�	O�i�ǦE�_4)N�{k��SԻ,g����GH�E�&e<a	�#b����-9��}��zm=E��@���0D�/�
���N�>���,_���!���(�۴�p�U,#Ll`�b���rNA���¡*'uG���ڜ(9���DxS���O�F艈3�\9�T����Zu��8��d�io+*b�%f�������N#�.��)oVR! Նe�(C
㑌>����qD�<���R��z�-��h�x�������hm���M�?�tk͑P�҉Үb��x�q.c����يs-~%�
ed��ѳ����V0 f?]4�i	�D��:ow�=̣�8�}��L" �LX��W�w4٬�l%�h�߯K㑄�T��O�y���ii�?�Ҿ�R�j��JE<K[-��o7E���i ����U��)K�+f�~s�'���Ҡf��s�0�����ʪ����E���C�R��k罱	�7sq�&�՘+B3f�u �]��?���@��f�g\�H����]Eg���'la`�B'�^^�P.�mZ�F�$�O�Dk����҇y{��N��ēR~�{�&�갻�4bYb��;̑bA���#*��`��"r���wY���N޻}�7F��r$��o�Xf���T/��ù���w���b3|4_��ң�*���u�
n��ՠ�����{�.#K"������?��V`U��f��wduҿh�U�|�	�O0)�7�Ueێ���N�I�(�}���S���@���c��ف�#��g^NQ{�=���c��e����@�kw�~�����հ��Tv�/���%a'ێ�ح�N���]���y���ъLG֑4��������R$�xL��0*Yh���'2dpp\W�}E�/������җ3��}�l�����/�O�Gg��G�>��Ʀ������������8D�x�w�� B�*؂�Rw��v����1��x#�ռ7�; v�׌�u���WK�p�$����Zq���`����w�@�8<<Ll}�pu��������IPdJ�P�����B2f���MQ)K�7B�/��gw���9xޑY�I$��J�R���nǍg��{��ܬ��/��0�(�e^�Eu�a]���'�n
��P�F�рy�bF`���W ��I��-,�걻=�E���-4Ps��~�ˮ����[T͕��)8� ��Դ�9&u���󓑈��7�<V���A��f#�H���ԹR���K%�V�R�}��o��ʛ��l��$E��%�
ÉϠ��޺w��HV`��St&�s�}/I�4j��E�� GC#���Z�{�kk��8��v�dެ�;9Vf�)Y��C�������#����⯸xs?��ȝt��M�@B4�Ԥk|M���߂�"������2�`��(�;J9�D\�4�*�%�[:��5ő'`$8��r藈X@�&�^�w��Jx<H�i¥tC�9BӍZ��0���ʬ�{ub�#�w��U��o]�q���PCZ�]'P�W�w�^�ӃU:i�D��z�τvΖ�!�<�C/ �첹�"5Og��C.�lÆ��*�,�.�<����PnѰA)ܺ1��[����shQ�ia��\ϸo�hM�k/Ք�zL�wEy�8�G��{w�~�1�p&Z���uK�*Я���ٖ(��((��NR}�}㔷�Xf��i��m��k��/��`��M����@��4������*�6/O��B�ҙ	��d�=�N@t��W����PU^8#�t����+�Y�U8�B�y�P���Z��& Q�����]����u,�K�7n.�$Zۣr�VȢO�N�<Gk��x�G��?Z_��f�zs��Y�5P�Y����q!�!橷i�\:��u�6������#�11&��P7ϫ�w� ���+�W+k�v�ztY�KP�Y	�5s��<�bW�(�s����6v�
%���jޞ�хK>�g�!�#�����e��/aJ�OU=�C�_\^TF��A#��"�vC���OGne�/vB��F���rT���Hd�g��5XvR��XQ>��1M��w���}�֏�1�Vk���+LeE�t�_9>~Z*��L3E0�Yi��}�	��2���e�����HRM)C'JމHN�β[�^P�2u�l�q��"]d��b�ߕ�G�.��c�[LGnA��.(���NYV�:J�8aOR`�*��������`����!��N������`-��B�-�U}���4u���Yun�d?��ܐ����7R�f/�8ۺdm�]�o¸��xo��B�A����aۋ�e)z�����K��_[��Aqt%��ހp�x�$���og.�Fs,�N��t��B)@�/G��6`���FbmG�^����V���fV_?�o�17n�	�7O�IsN�B�v��Y���V�V�� �!����3�t���`$����MGNcovpmy�8*�[�������v~�/K<DS�o@���Rī�Gc6�_�ŅvI6xq˳癭��0=�#�ӓ��`juo� T����Ϊ㔔ykt���;�=����tD�H��� �҉���ıL��׋E� 49!�V�U�� ���qh��?d���%_`j�`�҉�|���GV��~��'�;4�,4 �x��mKÒ������N_A��^%d,�5 -��Z�\����삘l���ʷ��8�j�7�@���u�vS�#-��>��	s�_%	]�mN`�
(���`��� �������$"����s��a�F}VD\�Q蝴��.r`p�~���uf�l�P��I��	8�uN%ӏ&�|�%U�q�5��Rs�e���̘AIB�����%v��!:F��~S?����
������(b�D݈�� �:I���	���i7��9Q�P�y�����.���ͻ��%8Vr�~'�*|��^�i�r�*ZT��0�DH�7��Q}�#	�?&��l�0o��l�bٮZPts:��z�E�.F���	Cf�/�h��I6�������D��������ժ�5�ڲl3��.�*��cc���1�|�t�:`&v���^�����o��4	V4=�D�O���K���:�V�wgE�5��r��3���NN�9'+}M�z����h]ԬP���Af���B\�M�9-xE����,���A�.�_���x��"���#��/���3	#B?I�,�C�_�qi��X�ߞ5�\�@�F(G0���
f����!�+Yg8�)����� v����I*��bbV����)�G�����]��7���_"�`�R�L"��H�Uج�,��'��nD�{����������w-�5�k�N%X�
�f��y��0�>��]����Ή�?%I#������J�mv����5k񣑮�Ը`������}3�.]��eV����qv͑���+�2/ށ��O9�R�qL-Fp�;r3+�ݲf�"�Y�v�VK�#�žb�@&�F�x����+���ٕ8��-wZ�KE���|�?�`?�(�4�|g0�F�[i�h.XqH!��^�j��-t|�t�灗�[Xw�6c��ۥ
&�u�{ a�;�G�0F���}p��/�_q���,%jв���X�8��4��2nf��]������JM��v<,{���LO6������-�Vz����RԾj�W�JS�U���$�������c�L@#<qH��]��,�.O�.p�,z�����L#몉l�[�յ5t��c6�:F���<0Z�{2�G@���:�ߨ+}�^����6[�$s�݉���>WyP�*�� �3�G� � 4��MZWG˙�(�8m�������i�gL�$t-�.r�`�&��|P�����f�^�	�}e�OeG'	�ʴ~��h��$������G��TxJgsw<c�X����� ��>��.���ۭHv<�[4���f�|�dPWո�x9���kE�4�_��]2)�XzP�=\�1��5���ġ	��E��c�����]n����[�.<�C�]���'����a�x)T�R8���g��>H��ACV�h$.�`�b`j�{�Яi-���!u����� �ҟ�u�o�>��^��v�)��1"4t�O��I�v]�����icp6���(��Ի�ja޶����j1�g`q�_����+���,D�l�>����܇��t����d�t����q&/��P17���G�q���z�:���h#�l��`�z�]�s�W���O1�N��ց�y�g�HF}#@Z�s�+���]^v(=#���Qu*įs@|�y�T)1�|�LY���D�O�����E�7x�&�}9}�W
�����	1�c�Gp����E�@x_=.�P69Sڷ��_�5Hv��1z��b���stK�N�$�����[B���?�nd�1��L�IY�����oGX��?��r��5鿃��?3G
�	�0{��\Z�
���3��3�b7,�-�OXPͣ{�Kw����q��YX�����?y&'�Q��0�eeY���w����s+��iB��Ĵ-:?+�`5u��>>��ܑ\�lj���k*�|��;.��k�A����S���Mi[�&U���g�xe]"��F:b�ؙE�!�<7��E���H�_�UԪ�|7�ѳi���m�!�pt|�	#�}�c؋�a�#
Ю~���yy�rD��E���}�3>2�E�l/s�U�Q}�ǫ�dz�mv6yU5LH9�Ln@����Cҝ��������V0T�/��Nʩ��3/����� h�\A��J���7��M��N8\M)84��y6 ��\|@��J�W��{"c��Έ�������ȃl��!Pg]O���6L�� ⽮�M遼'�-��(�o_Ps4Z�Ȉ�+�Lh4ñ�c�����s=,����L$�[E �>�}��6��`o{qm�-k�N��ġ�d��vv�ĝ�ZA닊�Y�D�1�a8�F�\�Ē�1��ꇧ�����a����_m�;u�[IŠb�A�n�˨��;� ��4��T���fX^���,��g�K�	%s���P��KE-��v��A��2��Cp�f�ڋ���84�i1����l8j(��uX���cl�
+ ��o�V]ԒZ��-�ޤd�+�������T�[�P�o�]�?{P�2 Hұ��������y_j���e]!��d6��"�	}�*���c�1�N��}�����B�N5��� {�]	{��нgb�/d�@�$�������%�--�e�J�5����FiI��n)^y�g�R�/z�u���m�Bn��&���X��!K�&)G���|2�AԺ�M� ����8��Q˥t��ėد�o��w�S��d���m�[��@�w�����1I�[fp��.�/��h"�E�s�V�\:^OC ��F�F]��,�n�+Օٰ�a(u;��(�1G���V�b�Lv��й��/�ฟEv>�N��of�R�Ll�bKQb��I���^�S�T��+F$��Fy|f;�Xd����U�W���B=�L]�� ќ��6k(�k������5�$)�j�Un���<����s���6�Z����v?^r�ےu�����F%w�ϙ{��spP=�e8��^s� hKN���dP1��0�\�O�E`���!s3����A�~=���=!��i��k�Rf��X�^��6ũ3>� �|[�gC2��x�$��O����;Sz����q{B8����#jg�jX!��9VP�),���ӭI��@Ty5g�U3+�&K'W(K���74�O&\�r�_�`ʤ`s��o�fo�/��l+�ic��xi�I��x�[R�5��YhJ�OW�p�����ƙ�zʳf�!t(�-���ݑm<c�;���蓼��tj��f��ڵ9�@��'��Ƿ���L��2:���\��7��?u�+�]�u���r���R�t,�!声Ӭ120e�N�Q�1��4_�H;#&9�?Z�r>�����y�n�8�q�q�����.�ݪ�^G�N��U�D7|,o�oE�j����s�Ŝ��+.�w��[sy�nP5�ev�����:G����Q1;ԃ�
�U�!�|u�W�*KnL��o�H�o�e����u5�s�(�%����wB/�J�����g7��낺�4�c0�4!+;�U�����Xn�4 �s lU�E
/�G�ߎ0GD�x��!Yi�k��dk�~4&�~�P����;%"�ߵ�M�����J~s������r��]�j�1ύ21I�燏A�7�N7n\<!�S'=�M�]4��dR��f���M�Zs��tde|�P-,��s�s�$u����O%:>׆��@��^Y�G*wo#�|+%W���Y"pwp?!��s�Ttf��Z'�q��EP9пXqx�Z����F1�솘����0��xX'#�0����z"������v@͚:V�[��A��r�_(�|FM�l��kGC�d����\��g�W'H��@xV�M��k'�b4��୛@�]���/6�t*����fVz��v^�]�;u�i��F&���J������r_�
�Y>L�l\m
��Ng]VQ2��rU՚���3�	��	1�����ϩ�8��z� �]�[SN�vQ���Iw(��<�FLzՖ�C>;ف��9Լ�@��Xё�6�����\2؝AS�Vo�֪TJ+�A�!�+���+Uߎ���J�*�{e����k)�d�{�1�YP��5���t���\�m��V]�ob'랎�Ԡ�X�o�b ѿfԚ��[_�⮐ux��-1�q���.�z�F8n�W��H��'Y)�bc�8�H��u�u[�2)/�(3���*�@t���EE/����s�z�r��}��������4��7�A�^r3F���od���Y2�b��8n X��OݽT�gqG�����9��	�����T�eR[<���m�x�a6.��%o�ަ���9%n;t0M��L`E�)�!Ҩ�1�������w�� �p�f؉��ћ�d�����㈳f��{P�қ���D�P��j50�e��E��+�J��ٟ)�a*���h0Q �Fr�Ǣ�R���K�j6m���7�"�u$ڜ�o�A�f!֯�[Z)`�F��&���PA-e����e5З,O��/F�M�n:���Ҙ�-�������nvz�F��ZhR� ��2?`�:��}j�4�H�?�n�f1Ӎ�3,�� ��z"���ɖ�x�e�P�9����2���Qn�<ѱ�����,�{t��nv9��C}�u�TS!�%��à��B"����3nW��+ˁ�ތ�,�3n��e�;�Q�����ފ1�2���5�:�e����lZ�2_ݪ���"��RN��#Xp8o;���l��i-�5b�x2�Acx�Y��]���E�xɢQ�u���z?Ͱ� ]S��' ���k�����Q��u�p��?�a2h}�]�H�Wrg/�%*3��y�� ��=�[G���X���{�S��2�d�	� j�[�;��t���|܉a��:z�$>ad��Y��HU�U�V���N��ѐ4��G/~��Ay�N���y��HK�(�=H���o���U�@6��fǹV�}9� 	Ǆl隯I�����Ļm>{'/��Ս/8�`:�L ��+"�*����c��k>}�%���k��"3�rG�P"�f�̴u�]�m&���T��8U_��e�9��a����5qP���V��1غo-z,"$��x��ʚ�d�,��d<5>�O9���Ś�`���B\$%=5gzP��~�D��#M.��9|�q*E<6��_5�u�&-o/ZUO(+�B8G�q���n{_���H�2ѝld���[}��Vbpؿ�UJ/��#&���q�����{��:��0����gW��m���&(����Afe�hELx<����ʋ�D�{}�eg���!/� ,޲	�B�V�G4� �+���t����[z%�z?>0��L���W�p��Ha*�>w{;����>gw���3D�8�m/���7y��!��3����S4N(#��U&Gb�E*��`�.���� R�폾j)є��1�-d�ݪQ{3`XVa��T�7ں�n�0�?�Rd%�!N�]��R�*$��E�+�oC��S����s�>A8�j�BĴ�6櫿U$@"�Fu�^�Y����dW�)���[l����݉G��D9��"�j*�ͅ��ј�?�E�;�l@�Z��*
rJ��A-H��`�~�_�Pwq��S�~���#��� ^���K��C��I�S��*55���ju�5�旆ַq�����/˱�~0�$O� ��~:��̈́dm��A����**F9Xx*��U��q��a#:tk�l��| ��8��i\�5��qV:�⶯����H�j'H�&3� �n:M�� ���	�FP=���}ɨ��W��^�R^
e�D��r\I£c��=��i��m�(�5��&*��և�[ޚ;�;�$�{31W����z�٢�iPԫLYd��m�M�\MX������]�b�"��*�I`J3���v�*�գ��J^D�����E�ȓheMN5��Xl,���wJ]���|��	U�pz�?rB��cZ�����ҶY���oʗ�п�Q��<�wB��I�6QZ��h*+E��;���A�����VM�ӡQ�A9R=[�3���H�G�����l#�����яA�P����c�ʘ;ΰ��]vV3OZ!|��t\�g�lIA��6$~�݊���ɪ�/u!k��F=x���;��8� �*� �|��}��X ���i�c�5�A��h[;�h��|#�̵�W�v��R�~F�����H���<�_���z�u:g�mF��D����@�2��C���>c���-�lE��r`��i��] �U������8߉��'��Ɠ_�*^;,*L,�W�g�3$B3�a|UJ��.<���Q�+.O�~��FpA��Q<�ɮ.�bDLn��!22�	y¡�[�칪)�T��O��E�����(�������u����q�텯>�'���_^`G1�8���kn�x&>�Z��!�?4,p��*�i��3��}O�����.� ��t�V[�!9��W�n�"�,�Қ�PQFn��@�q�u�<_��3r@zDTn �[u�3ű;�l*>@����d��/��C������+O��%R@c�G}�1�g���p'ƥwBud6��g?1FaU��M�k
y�~��0@G�V@������3?��y��exR��Dt��\'Oe�8Qw)�a�sb����΃���c�:�F�, ���6sIn4��F{��XG�r��`�������΂�'>�Oý<��Ќ�e�B��u���G0�b�����Ujdm��(���wYX���W������O�p-�}&�]^���^�i|�I��)d��<��w���DY�n�f�y��"9�v!_gdnU�djXƳ����Ս����li�=�t^Z���2/Ģ���'���a�M��a�P�$i�՜:/��J xg����<Y�n8��`}�&������u�.�Ss�:[�?-Â��¯�hq�ʂ�Ơ ��J\�>�sՁ����*x?�<����k�ѧrfZ�ui��ڇ��&.�`Я;���o�8�ɼs?�B��>~�ԉ3�}�����_
0��f�r���D8@;-ln��cU�݇�
�tV��3��<�2
ņ ���}!b�m�����aN�_O
=;�+P��޻��F<�\&�/���z���r���P��tE���t��kG�Z��@4�D����m�]���
�����p+�"ZH�*?���J��qS��������.	��wI@�Q-D���`FwH������f6_�%����ӡ���l%�"ulV��
�/���e��'H�'�VXS��!��hmJ��l��Qm���X��A��|��pz}&�R)�)o���:l	Djʸ"����w����������\�x�)�0_&OԶj�&#�b�us�/}�O�O�A \�'�1�?��Щq7�\o%Ph`,����j������	Z�;mQ���W�+[ހ����e0`c�c��&�i�� r|J���pZL�{O���gp��L�E�z2QH�6[��U	���@���O���2����B�Vn 	񩝈�nwm�Rl�5ŘuO 2'��.qtZ�҅��PI,�ݠT#w#�j�w�����uHו��I��2(���* �$�9 y ����X�Z@��ģD���.�a��x�lK�6	7�B/��T������ZWC���Ku�z*�/m�d;�d����S *�!jg�3�Þ~[������+M~�|�3B���KFA�	��Ǐ� g���������+4��<?��zø1a,��,c��=�5,���X^+~�x[���V�2�Ϛ,v1nD�>J�O>M���hj�#�g�X�	p	`_ȍ{.��lD����5��8x2��x�T3E핊a%�֚i��P8M,�ϲ��1�� �N�L!Z��툱�%֯F��� �MO+��/#(��a�.\�fY�Pc���r�w_r��:�W��Ѭ��I���4����q�^18i�F�����ݽ�kwG:�e��4z��	��$]��A���
�zp����[_�ɢ��b���ru*|��T�'R\�t���ߋ�i����� �W����O��u��X��ȪvN�����v�����R���[)��3��L]_�<'�S��b��x�j(��m�涓z/X	S�кnvP�	�c�J�L����ƿ[����'�
7�n��b��BÈ�D�U
lu'���5���Ok��U_����Sÿ>�I�ne�X�1dς�&��HO �ų��'^<OZ����s����z9��ծ��mxQ(�nli}�lv���j8�g���=��
Z�(iNT��;�Y�;�I�{��[��@��w��M��F\�֟�b˽ys�v \��}�Q�:w�v�Sf	�"��Ej��M�n(����`��ܠQt�Er����3�Q�D�7��躠����0%�E;�zƹ>|�0�t��z��2!>��\t�"4j�bN��)���V�]�ɶi�N8���,*�[yj�MA��R����_�������ϩ��Y��W�?&w��Ċ��G�C�w��$���v
�����b��s�屆Hw\���gB�y�(��"�x��a�A�Ũ�KS�\���UN�4+�*��$�D���'P�g�5P@�N���JL�Zo��$@{R_����?�M*��o���7�^�ʫ�k��<�;�x4��ɩ�c�	���7hBrܚ-�X����� �:Z�mw�-ץ�':B�c��,`�f"�"^2�-�hv�G9Q� Χ3$)�ӏ:�5<J��b֧ �v/�M�M��&�����Y��{:J�.��G�]�k���(����?�"������P%\��E�_1�rF�^q���P��ZT����Z5��ؐm��%�0��D@}<�b�$ܠ��)��'�%:�F>��,Gʞǐ؊i��� A�,y5�	2�p�P�~g�a���A�HmD��a��Y�%"���<Ѡs�\ۜ���Q& v��.���~�����˳�?��(b�M`+P�d��%�4θ$�����s�ZA�2MO��.4? ��X��bR@���\"�9�������3���$�N\�(ۦ� �F>�
��w��bg���"�zpR�����z6~#5�E*-.+��D{$�����]�wl�yUW@��V�(E�'�3"��H$/��C�6�o��d���sĨ+��e3�m��kD����1�,2�7��3��W:�uu��mz7{k5H�괐�\hX�Wߗ	��}�tH�x��'/�!2D���nԈ�s��ڿF[������, �Gؤ�X
��Fc�_��lT�_�5{%��Hb����Ś�ڏ�!q	Cq]�i ��[�5�j�ܷ�d�����|�}�o�R�C �*��I��j`o{o6݈R!Ԅ&>��M.�䡂�#�ut ���g�������)��GQ{�U�:�ͧJ��5��@�^����h�qc�tVe���ݹq�ѱ�[��nv^^�g��<�݀-&Aa*Z���c٧*��B�6k8�| ]Oy-�	R��}�t��?�,��TS�##�T�1nE�k�1-�Y5��zN`I!�4"\�^y�fUR:�ʄ'��N�=W�)<hN���3����S��+��Ćq#�aSQT�|�6{R��`^{6��#O
3�俁���}�JS}X׉@�ʳ۟K�o�W��1�;*�M���.@9	v����!�w��;��Mc���{�XX-ʢ���N&[��5���&��j�u$���_�]�M>��m���6�nכ�8x�)0&nv��<Ï��s�2�r �������I �[	xh����ζ�W���Ƕ��T���1o..�h_9'��%�r�GM�����	�N�o�x�I�0��@�b�-^d�N��3^�Ԅl�;o����3��Щ.X3���]7�0��F@avvGiXӊ�{���"��A�%ږ�Eħ�)��q:%��kc�	u�N |Y�@�Ao�X�%��t<��Ja?�wÞ���x_E%Q�9�8��:`��V|p ��9���⑉�M�ˀR�������A�4I<���v����v��п��A��̯��"��֐�8v��zχ��0��� ZC�r�{����}���9����!7Q���z7�+��|Mn3L'p`
3n��E�j�D�>�����o�^Lb��?�L^g�Ī�?}o��ev��
����f�3�Z�cDJ�Ǵ(�vD�֗b2��^= ѝ|W]#0�y�]�y��	�����/A�ለ�m��[~����8c�z�&K�Sݵܼ�p%c~Q#�d�ʃ��}�Y�7�i�x�[�b����	�
��x����!&C��-��j�0�
�7b�.���4���hsc�u�b��D����Ővj���� �ePP�'�2�T'��m>�D�Evaɕ������-XK�뻷���o��w�	��o���p��I�S��ڎt]|#ED&VT����7w^&An�r�_1��=�mp\���ar'�SI�VÔ��Kekʭ���.�!<���{�(�Ȃ�rm�z���QQ�9bˍ<���2��Y
 �FL�	�-���4k�]�������:��W��sLsM��v`һg:���{{{I_X5�7~���d���(��Wq��t=݃��tq=��ꁸ�$R�u��tG�cb�&:�n�����.���>����HF����}�nO��Ȳ�L�3�U_,{�W��m�S@2y�G����Ԑ���/r�C��!Ū�\��yAhUzU;�${�:Tj���R��<���̓��b�N�a����93��̖ƐM6�+���Mm��3�ֿQ�T9	ϫ��]���E� ��E���tFE}��YM$�-	���<9{_�����qm�"HM�������4�$��7��O=cV�֎��Y�z�
ni�;qj�����p4�B���Bƍ�F���%������퐣<B4'ϏJ'WUl��~�=����4@�y�vɕ�$�˽_:��`x�|��o1���j���$�z?�YQD/���-����=Z�?�b�{֊�2qpO%��Lm)D�uz|"�dK;з�<b����"�w� ���t��p�6	y��.r�Ze���:<N��
��f&Ž\�Sr�nEF�,��P��H��y�ԧ4HOi�(O˗6٤���j�=�z�F�8C�C��s�Z����"T'����f�ѷY��Ծ՘��֮m�KԗKT�l?�B���nq(�e��|
}��@�|~L�/�n�*��͂�5��ʆ/9j����M`�Yo�T��7���}�!b�{��S��V� L2xR�ő��lց��h�R�3�^0��4��o��.��鱎T�,�|6�VQ�N y��ס�gTX���J&�i�O�3��.M��@#\�{�<V��0�ɺ66�W����(�b�@���[����d�MyT�S�|����-�-;T�e�\�=�D@aȘ2�7[Vd�ɉů�	E+��M��2�"��S���;�<�F�l����~WBh����B��`���W;�<���#�س����RzƤT��@�U�t�L-)�0�R�579�YU�ҢY�e��_W8�J��j�#R���T����}v�/\�⍛0JzWĕu,�4ű�׿q߾Ъ�O4ĝ�-�{W�7�s%@���i�j���-7R��D!V�Snѵ��H|f��	�I _eܮs3��=�eiD3]l�xɼ�F�<>�����7>-���:,�����G�f1n�������^�7��4�{/��b���׼x���Fn�<տ�	�3��	#6��KQ���~��BRvno�~x�/��1�C�~gh��5�QBrL{梥7`���>��#y��7�'ߒlr����r�{ �c�0P�����y
�Ĕ_X>�9����]�ו�G���(��N5���%[V��փ-\��*�g�T
}��Hf�'��Zƌ�K$�0��Eٴ�%]�B��$A^�V��6��u�+���]&q��v��9,@�[��Њ0��x�Ŧ({q�ok��e�\7�U_d����6����˛\�jpǜ?���ѯ���\�9p�VF�]q�A�tW*�*��-n�2��W�Yܲ��*�u3�q��u�@2�\�_{��$��h����'(I��a�;���P�v=�z�-�a�q*K>~t���9pe��_��D-���>a���� nr.��W}�vn.��M�����譤z��O7j�L"ċ�.�c*�Z.c�GȄW���Wwtf���Ĥ��_ �����⟆*�JYT"uh]��w�X��1�B����=��K���W�ج\�}s�A ��o�0d֮$T��g���a��U�T�1h�L����x�p�w��s�-t.���\V�3}��z_��r��z�ŷz��T֜Ӯ�^>qM�0C�� |,��ae�����*/��>�c�����$�c@\�mr`���=�M-8Ui�"�Qφ$_]c:�j�$z����Ǥ�ս��iSi`	A��#n�J�@�JD���\��֞o�&�P�_-D����K_o����DT�4m��=��d�� %x�
����F��^{(�+*�j[�;O�����M�����[�^�,�NG��)��'C �E �X��o_�YY���k=��8��`Z7@�+�Ҭ?T@�-���ËP���Q�^��n�ܠ2,�\WIj	%ѹ_zq�"�8�lM`�_ɱP�_)������� ���}�
��1�!m��ٌ���W�n��φY+5�P?91pY
9c��k�Z�����ǤP|���%>��^侢���{:��Ʀd��	�V�6T�v����򁅐޶g3E�W�X���|�r\��ͣx���=�{�!O��oϴ����+\��y,c#��=gQ�4�Զ�ŏ��D��Ŭ��@+�>��n�c���0:˭�\�,�����'���Ѓ�_X��>d�������L���~&l���YM����?�>(����+�*���dj�;\ؒPB<M��|qk�)G�?��j�/^Xp;6j��bqv�/�K�Yb�GC�4��jP��;g�Q(-�7��v�?ҕwz�_�[Lx��&X��D���"B��P�E�9�f7��1�p����5B��6�_k����Gv;a`y���gȄ�>Q�[�����\�LdL+ӽ�&����9�MV�wOJͫ�>!'�20���9��5\f�����d�^=�+<D���f8^�n���8�ơ�گ9�3ܻz��:�U� ���x�W�př��p5��t��'&\��`���4ȵ�{��VִK(,O��awڭ
-�Bi�(�*�P����ډ��[��R�H���ܔ(��^�6�������2x�W@�ìץ篛��]��������Ds*.k�g�onfG.���0L�<����R�k�;#��K�[�s������YU�=���[.�k8G����9�.J7įM0��D+u��wv:��%��X�[�`C|A�8K�9)r�3���rƿ�Ҁ0�ӯ��#���f�6��+����'��Q�l4�� դ��xH*r;C�[�Ftg�(	� ˞;[��[��[o�s���l-���Tf��C�����t�N�6~e��y�`��YU>�@H#	dZ��j)��`uI�8>d���s��4���tR��V�85X��~f�1 FR�/��}�&�+5L�s��L>vږi�d�/p��斓��Y��2 r�.0���x�$�D0���I�p�>(��/V�!?�?GC�r���9 ��"1%�;�=�*<"M#�����,g�TC z��<�d�������l���p6�!_/�c\�~;��m0?Xk\:9'��Ql;�/rMDL���t�b�.��AӔ�{0�S$�"f�Y��+�mRcz!�d-	�����ȟ4�$��?A�6��|}vd���K "#,�akk:N
�h0�P�|�rH�Q2�yNh���\M��r�ȳ<���:��W>�B�4[ΒB7d;c��07�賤H��x�C��Iok. )�|Ȅ�<֧�hx�����8;�3PQ�]��t�-6�b=�3"6s��d������y�Q�n��~�m6(��߬]��z�o��,��yS��?��<�L��e���Ց�1>���޸����Z�S�ʀL������y7{��b���J�?��s�c���t[����<��TϹ���P/1��&A���F�:4��Y�ƪ�4��lTz��\^�s���[�6������6SBnxI��-sz��c<�v�%sx����h��9.�R�H��� ��d�~7���R�*@U��L{+���"��|�t��/K����N�Ȕ����I��,�Eo\���*����M1�׃0u"����2p������{ N�pח�śŦ2_��08��\QJ|a����?B�/���s�6¯k����<�[bu4a�����(GE���������OofS���g](}̿�q��Pb�7�א?:��JCi �#�Fs:�)�P��/�%��ܒ�%�X�����.]�����C���Y���Ԣ
1�-��ހ����)ͦ3�ߴ����f����*�L��[Lz�N���<5�C� As�����&`E�����?��+:���7�L��i^y_�}��e'3�2�eT���79Z;;�>���d����z:ZS�8�'�8B�����-!2w�D{/c=]H<���_ @�������	L�i�Xc�u�Q�=�#��Hlz{�������!p�'��K�7���T�g�I�%�F���FW;y��i"��[�k� 	[)��m#.���oĥV�:?f�͂	�։Q��Q�������R�:��`�BTB2[�[������A/���yu��0�7�����D��lEA.O�b)�>*�A��v`V���/�E��?J��
��k�;�ϪU�#��.h��_�D��[���,.���pr
8��X��w�L�H�%1���;/}[��ޕ`UR�8�42�|�N�m�nӪ
\ ��	��h���)�����HI�gNc�κ�6��1}��yw3d�a?CR��-��`��y�c/��?�#�⟍ �%`m�ܿ�ӠT�'.������˜]�K�QvıD��Ѱ�MT�n|��t���e>^q��
����^Y�ޮ�z�l*b���.i=X�!f{�?�ɟ(1��ZJ��(!k�Ì>\��N��p���67zrs��:��R�_%ԊLj[f�99��UJ��!Ж�W���<�����&����j�R��E�V�9�����)���HC�yk�B�V�S�@���G �(�0G�RCi�/������׹F���M�$����&a��iM���-Rg]GJ��q���g���o+>��{���[�zQ��_��-�	��D�]pZ4�U�촟��	{������L���x5�m�/�㉢�I�&}�r���^wè�����0��pf-��H�	��_�G��̈-��'�j���6��V|��ݿ]��|�i�J��&�M=��n���/(.���u� E�&�/�,�Qr��-��y��6轕�#�}�HA�N���A�0�u�4M�;lA��=Sl���I�7sf��A��*M��R8�	�7d:�W�5�$od������M�x,���O������2ʞN��6[��?���mq7P���˸���u�֢])RX��@A!�c!�!!�/&���+�3W��͌��s�4Ʀ�9\��䬀1gτ\�����N�(�.ߋ{+�l���§Q�R�w�^ݿ$��c�+�6�(6l�46��?z6�{/���!�@xw����hu�J�<I��(�0�I G�"A�O��8
�*��~����3�q�`�i<�d]=M
4m��#��w��+��
Տ{Q1#SJ-S�U�-%K����`���\]�W��pp��G����7����'�*��q�LC�y�Z�"�ٲP>_�I�]���J�}���:o���(LT�X>��rHg6���/���b]�� ,n�:�Q��"-�~?�,�U�&��i=�����A0jQ��r�9�FgԢ�-U\��������x�js��G�w_}*�[���\!̈\_�at\Sr���p� ��rI51�?����I�U��[!�[Emi���T�t�tu��a�2,ƑV"������@<��kH�E�{C0��!�5���ƀ�i�T��K�Ӳ�{\ѡ}%3�i��T��J����9_�qS�| �y)�;G��$��޳,h���s�P�sX�&l�1�h���xLE�(=�!ln��;�0�)z���؀�F%"�.o$d�w�r
�&������yǉϒ]k
��~�>`&`R�״��`l������b�7Z�}���o8���'�Jv��F����]�*#EQ����aAS#��� � v-�8%	�4lQLSB��S_Ή�S��h��dVX�ݷϵ7�2u�b�c?t���|������vї��vO� �>F��Uͽ���l�����j��������j��Tp����iÛ@&Q[2���gʰ5O/_����p��u�jZ��%.�K�.��͚~7S�