`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14912)
`protect data_block
dxqxA8UqaOQ9F1joSxMHUiwvAxPR1Ij5ySKCIymLaABElnYetEZMMrtNvHxNFOUD5OubL8dGBk5G
q1IGNiGdXOd5nko/1oYHZKzS/5PnoHaomZjIt2d8yKykxNxch7oV80k6jr/1c4EIf1NfUUtutFgJ
TFSj1UgxxD1r+yr+0nx1l0VrJklo2P8XNZlKqkzuH46oF2g6v/NUwMtUTTCe2w/GGmUPFOqrGDn3
MgBzQtHZFK96VkTi3OMsVZ010iHfdv9tolsCtWG/PHr0q9kgcNIFv32uUH4kqhRvKtvVbxIba7jY
UkMAYxkwBlZndur1p0kom/Haa9gglAQaoPCmzvXDmT3Po+d4B+8Y2VDljyRNTYfe0Ug4YRqanKMp
2Ez+e0lXuNfs5/dtznd1/+qcJK4bIT2ilbQbI7rn8oxslU9smEeWSabx20NGkdlllMFsQEHrqLqg
suZH3VGkIjCMU9+txc0vsqZ5rI5QiJRQaekV99ikIHK0St3UYh+cx6W16gc5Zakd3VdvCEp9BohW
sv4OUf0YlFu0OCvepHXvua0Mzha67CiKTlkNmB9sYRsIknJM3A/DWlyOWGiFJHfhwLGLA/fNrZoP
jqsfvXyVj8Gbcgo+Y1pGyW5P5gue+Pw8XslkncWCWYyYgoW+VEEjwQA8NzVwEYoWuOvDrNwvbJJ5
2oh7jXAcBqZ+rxLoqK5UQXD2dOzIZ2K64z0iyiu0PAtgKV0LspjhUO22Tsl9noGh6fJr2UGi7T0y
NVm3zYJNmp8ve1h0DJEwlcrgVjCe7RtZc6OWLyEMGhP2YZzFy+2qy2rTQQP1jMHnm/jC/qe1WSwS
4Qy5iumpXz5rvZI5WbN4tGMQYH1gut/e1byKTXU+THCcAT7Ro/tpDC2T8jEHXVP6i0nuyVjgb0XX
rsZvtaMFO1CqykysBFBVJnmTBPPZgP4HdT8qgHLZ+BCQlcGy80Px2wJsobd2ZGCgW4GFQieV2bgz
efFC0QTalLPrHVzo72hFKJamXeMJyL9Xd6PAegdSFyntprIgSn7CMNex8TM3Ey6+e1JLBf3o/SL8
YH8ixF3Bys3B/o0K+aSWVewEbUiFYf9uVwCD9onm01tetvBEoUxU1AtnQ+ePtAz6ZJsV2C9ifGdz
ngYn2sfoKe6Fv/BZyn/tDkRVZDubH0lp22ph2bXcSga/RWGKvrE6J+DUR5rjG3XIGWmTtYNUozPN
jtB1aYwp/VVqX6K6KkEF+2RP0bwzcFN2pi8WdWEPzUSh9iaG6foESbFTXaJyGJk+qAkNTbgROml4
VOEEsnUhDUcSZmWzbKzD4GOco/fFafzuhSOppmMjDKXFam75ZGpQD5ARtZsj5TGwhgWKbLoR9Poy
q27kgHy4DRz+JJRxHTSQsYbdxZz/B5ChALTlC8AIdTtZlhZsM9S9lNlBLHNZZ08sqWzb6LSJqTAS
CF/OL/woiAhfPi7P8DWqHUkcY0Mj3pqwhDZeFCO+CvEAUL8NuVn5My2rPGNc9NY1ePTGJMis21Fu
g8pfbDoStGHAt5bfxzoUkNVf64NHiNrtB6PEWiLDADJg7amGeX3t7bWMV5nXTGzTPoUmvBcHY+i4
xtgp6MJpPMczmNpRe7FZehAaO3KUTvuhNB37nnSowy6ix3i69Gudr+UBiqVxBj+rU4z58pDyY3EH
NOdrofscZMBgCUnp2foXZCdbOFz/oKdIJPJoJ0p0SM0zQjlPhrJuaIutsf5lXLI3pMfr1swDNDwT
A42S2lCcvN+4bYbk1hjeUfgHWpT51e8a+nF8AbEHX8QaW6LOmXsn8OFtx5D57rXgjEGBfzNXN8Ez
5ogZmSaSS4VCOf6qq5n7I668/MofR6rUFm5GGaRqnCVFJPa8ODdE1kXEd+3QvAFPsEVV+BAxCT7w
fpmlhGbu/qT6JDsoe+UibpaNFocYFKNpJRzr/BdY6HSTvRqAbHS6cWK7Vx7XFPD12hW19nNqzSLn
65CjQTz/Rr8mnO2NGVnJEf2ztWKI0VdSBjxO48rqDyq96dLOT1xp3scJnsgbNTWowhBCprficOns
KIQnJCIFWRISFOx8BkHtRs3efWdu1kiP6eZjd1eShZI8oJAlXEIwzGYhbj2gsc8HuGgkvW2pFL2K
mZW3CQPRiOSl4vJ2FBsWowYAPBVswEsnLswwgqHci+7WxzQByH73cQ3ZDMIUukqktSUvBtcV2I4a
vGvTLRWf+H3Z9um0XNT1AQLmJc0X+aIrnIHTl8tAyoWM/I26uIvjM4b10WS9sv6Cl0JAsBCXSY4/
9Ku6IqCAjGIzgz0Zjwm1w6uvbS9+g+z3DCFOFUfVL3t9K046Nfa/6guyM0E4vAScNk1KbVSpeR5r
SZWM9xxoju0xuMZYhwmT6BPSywUNU1CMT05I0+LaYcq/gSDiysGV42eSD0xIHLl4+QTgjocw7hJD
srWS55ZIBHXbsXveVYZkGJEetMzuWlBXgyHeLVvfngyLskN+3kAtoDD5ZhR6cWTcu9UR8+RBAduG
OFCVwBAbL4KqwRMRg/TRCmQKAbTAvgXquxuT+1+nsH53bjOsLIPgULLs3P61gHJSZuceQoeO2vos
JjXchgx+ZIL9SgpZA+MbG0NJEI104uomySzm2Y3hMUFpkALo6vPC1SGUMPBk7NPDm2ELtbD38KU1
utbkR/Q2iD76X33WJf1byx3j+gIrUuNEweC3nctLFLKmIkddRG4y4qBIPZ+dl8qBfycsx67vej6+
WJe0Oc2OJZLUNO5+HEpEc5zga4MTYIuxQ2DREAUWfh4zFNpfYoAfbbZmgkAX3fMpWUSTUPBSY/Z+
6LCxMw0FZn+rfypsCYRlGpisIpC3I/OjZP2VgSLT/JO6ekxH2BfjQlyW0f8GIX/XUHNTnnTO0d9I
2DIAF4CD5mSLZvVLoo6pCxC1VRCfZ8rMykpAYBaIjTk9M1n66GAFPYB7eP+Icw1Mg4quNkCMnpOJ
dOAzHP1DCMabCA/EhYqKQckW0SsfOhrEhd+9S7qW7pDY0+T4XzGiHiXG5EQXEaGwEtZXO1KHzbZI
PcMWt0/TxF2SkcomDDA9OV6HXmo4ysL81JLvrrWwg6tEhSp9Wlfpjz5F0e/G3bOuOAraIwtbvByC
5bOcAbF7SeJrZjzKLU/q1NBFTTFF7rovhFaPH+0VGHmiT8g04w9OgH21zHdwZaVV5B2xfxUKdofd
WOCFQY40UWQGYcxtUMIhPlyHXcG55UzrkaiimpI6hfDStvF6/uUm8wkDVIjObrvMR+zClKLrMCv8
rVNIsRBUR+qRCDGQYJiDUpeEGTbiVmV3XyJBWk+tpdc64lHo9l3OJRa6HeifJt81mTd+O/LbtoeM
1EWFetRNvrx9OfZ9sbl9difIgh3omx9Cj1BMuhCeg2vm6duLHYp2ShysdF7I7sbxQdefaaWMwf7Y
mar7UnSfVD5Y764uKmcvemvBlG9TvJMLLz3wwazpqnHFCEiPjfy5thP6tOg6TkgrMs9CU1W1/J0J
8zaV76drRdWvZ7BISItDN5W5Et7bWwIULTt9XZPbI8l71QnQh1EXllHeBg7RIfURsAcCFLBQYUNj
T0/ZinwqV+NKb5zvvmB3XQ2GQPbwcGkXdluIkHMaGr9xIOFqfng0PYdnxUGWatFrrO8QnSyCUJXV
FvjEVBLhru8FR0KhXfWqZoskNutb8c/IyDi/eM5J/Yto4tlERwt3mmUzkDLiZbBHZZOm2TOkMWpZ
PN30Fz/6PV7/vXiC0rjZOUPYi7QnI+lvPBzML96h/YM7QX1m8dBctDoJhGu5ERfb3GQ9vvPuI+Dr
3TFwMMByUFHiH2fyn5/yiVCm1Bk6fR/unlsf9RR/8zh+XY4hsDozayjPMdfCN+6nygCs14YyUEHs
kIeALxWe15tQc9EKtoHUphlwIV831iupsfajg/iyqTwGkfKm/Ed3j03nQKdERHBY3tzA1Xp9iw/Z
OoJzZYsBbuv9FAf57T1+lYiJHdkcybPjoH9XzuYcgYzNiqHZZcj/wPnp+PYeRyEDU7FbvdZleCJl
BYT2L9krg73JWzVlxeB/FEkEVGg4pHrNuRPlX4tfG6+fSbQEf9ogpeTwD2C0LnQ6gcEI/dDDsAZm
A4aGn3vtJ8Ga6w0z0iWRVVZ/BUH9pH4d91Y1UlAILyzes0scKIypJJEZ0tMzPc1ehsoQLostINT5
GpVaQkpD6S0THJSUoD2NcAnqilkVULbJqZSM2fDyclBu+2DbXwgVd/XYmiB2uKiJvWK1dvS8GkpA
3hpy+2qp//YhYZUVAqpPV2RtKwA5cBuyA6v3+NVZtvviuTgR2cvTCNGEhWQ3LslRaPBKGTDvaTbW
SZX0BIAVBeGCgWnCkgN4JE+lUE/hC6piOEozaUAzporSNrTZSlCUqeTOX1v+p/ytdUPOHKC1pLkb
U+zdwj1Yr93czDuVjzqljBZ6sEgCPimp4U/nUmk957SRZ+hXi1rKq3ipoY+I9hYmuUoeaQ8n3Eq+
MnZZvg7GIr6DInr1dCbgLyuWhEWy4kk2JygD0Cv409k5Av6zcSzymcW0kBXhNZQ6PwjgsCjUxCm1
QJy9gnbK3P/Hwpe/3PqO/1MzsMkN3wfCLdylzynIB2Qw+eVjgB/aZWh9uu1v5pbVlSL85wtdhf8H
Mpkm/+NZ3e757B5z/I0s3e4DInl0vfnl5+N3Ualno7vE6omsFDyg0rA3oTYudyeCF5dC1DuV/yUB
1syhEebWyVhhpjkP49exIebIKNy+d7S10ZrFsepoisGUPR49b1Q8L9YBUL8gZ1dvLOKaOKHcytvu
vr8uGarmks1eof832We5rDTFHbLmF6AtjFgbhQOga3dKJS9Xqu2O9uqHGujLUm56SLSd30SMewwm
nE0MK3lqs5DS6EyQq4x2FK3P0+PUH58GrDrRy6fUOXRhnCgaELxGdkhNW6XG7zMf4bnxmEosBzye
wgDrJIfJKnfYSuwOUmoM+OUzf7aZCyNsFK5LxjFxzB71N2wzAsk9bQqegLFC3W9aEdeU9ScuftxQ
1oAW28ktDlyokAmfprRgqq+6nfbDXIl0Wd5u+2SPtf1tcUtUHEJE/vrj5Yx4BUUiB46A/vpONEHZ
99KG2ix12r7d9czTOzioPF6vSKpRVrKpHnWYsyBUH/q04Lpxw96DNLh1mHG9qk9YdvvVZJ7ookKw
JOgAHf7RPzdI4qVFt4tieTqu+5Cvp91HNpt3NwUgD4qTWsoBDAV7q8E/VRi0Gqm14UaIrBzFUEYp
MC6sbJGBrUjegtPhaVmybHmGXmd3fWeuXkpue3emkFNEYkK372X7fuOXOCW+LFZtu+Ejw60uG4CT
i7bNJlmMpBTypfE86JAFvdU02giqQ97ZSqFUwnza3EnGMzhnApPxvHcnkdl/AT2sZQItsSaa0Zls
5S+/sfiXH+QG4jxB815ULxVrRjAuuyOPtk1BhYIYdIXsOHAjRx1kOkFMqxc3SAweEfw/Pa+2zT/1
jIsT0YeCRrw7H0Da1cE7WRp1ZfZT5YCrvzw9Q5+HcrpRARwV7r5E7ufS4Qb30MiWEnhtzMofdDxf
NTJ+KVU8Oqtdf3bsIWnKde5i280PllxAA23/cv/ZmzYbmVBmwRUf/SpaYGWO4ETuuUmTiYhROFfm
tMV5GnydWsmq+huXfkp91x3ZrgNiRa6O/Nlts3+WMfBuQ8XDU6Mf4eMnGOskcwnJiiTNvwkxbJT/
+o1e3fLK3NKcKlQSUextSIyaWW7o0KCTKRzMo58AEOHgdFhvOhSllfD4agVUwsnZ6riwqESaqFSb
cT9D8+P7x4rvsXa/PSmoHLY2G1OX8y99keIYt2i0j//lXNCpmI3DNCkOrG9gnX2hLS/xKY3qosrh
sADGYHhyuxAuBARgdwy3s+pbHUuCPZsYIsYVbPu6Mmo52RDnDov3NJfSwYJ5Xt1G+zGP5/qTe/7r
ONVnm73rbCg6zRECJsKbrzgle+U1BcKs7CQFjHjmoW3mYMX4YhnEr/Zo2TptAGVZI/SyYufqbkO/
i4jnqQC8N8QowS3LCnJWNI9ycl5zYMhym9b9t4jv5iJ+64iUMi4FBom7rJtd1PuHglfeEuKITk6t
cplxHtx8JZmLgcQ1/0tRfwPDBDs61OOIHtMf+xeTKVthqBBno7LS7+fPxknEUnY6Yu+M6JXuMHWa
M6B08LSB4TYHAkvqoYnBU+mZAQiTXjilTI4hnWnCpS72ubrC3E9OQdsySs0mR8h/mbCVu6ZRQIbC
V1lgGMRh2BxfeBrSaaUZ82sfERcOF98eV7yrRFkV4AFdMkykVCoLkKMSinwN/39OzcxZdQdzKmEY
TApCRgO6GjWZ0Xv9BXtKA/ESYEjVDQ7d57fAu7dfW5nmKbXckbNDY30OGl8TZJ+nvshVe8saqa9E
UGLfdUfdxhtNrCk2lQxn5JRehdXc4f0GJYIwvQ73etn/MBjCrG306tG+v4cNiLStMjZH/0EDcEHh
UxxtMQWAEAF+So35tFh7RXsM/SHN1b/zjWVukSOaajQtDOz6cfgSSSC9FNaEf6hBMawfQAaXaaFm
E8gwyPVuSuyFx7+ULtCX6IIxH2xFv2GMX+vbTJFPIbeDvDRPM0yCvfuBP4YiIS/Ftg0PpSG8d+ie
gURB7KsNi269YfZf/rOdSdNeXKSalVThjD/X3QXFAwmThLxoervi1R4KOo+FYGkyZK25II61eccI
CGCS6PBJ+IfXLc8ljBFRcevkJ4HDbi1XOYptHwsysN7y9XzMQNZPSUazNLerKBr4mTteIKwAp1Yr
UPHLQZxyL4xrsy+P9QJSizVmRO7A6fyYhdRpDnk4ooK0qsh4L6dSgAmjqps6P4kezsMtD/t/Jz66
BL41plma1ZnOBhkE7FfvLxEhpxN7H/voquwxlnQptDJU/YEQ2GbM2bJSJgE2J70+q3H/zN5Tcc4/
vGgmgAHe4MSXv3EdQA2rkNK1SkeDxprb3nAmH+uz7hTMq2PPgp5KV3ZpddLYu0CiFErqmL5YeXrJ
QqbrYsynTLdzjyD2FAEOvmRVrqIvjGfTnWDJaP77ckQuRLdHA6i1Tg5/PoVffMk2Lw/7sNrBPefH
V2gJr0ttJRzV6hcVFa574r/yE5/hI8H6/jWCmwd3qJxtSLyu0ukDnfpkLTBxYOg3sh9N+eIxZJQF
Zk1TDzBceNGFzp2W8nNeLrO7AeXAW2RsA+VsC9AYAG9WyLCBHC4XLVlRRvUW6ONZysI4LnZ2n0i5
avs2GK/q1ZcZtZYugaNkazdCJJ/ukB67kZdsHdjLedcz7ccocHyeYUWiLkbjsUlxJYpQ9hNSgKld
JLn5pIoem7q1pj8tPNU2iN20F368UoXDpwUlb6AWUBF/la8IjdYAmptW+TcgZpHXfaqc+KO+OLzj
3byT3IhJPvJ2oKYtk4K3RLuK19fEmnI2SbDWxQzUtfWxqurGgGQHsLQ0CT2+DraExzNJ7EXkog2e
gtxdDtbR9sUfKUKJ0r7M0Q73y3h+OUJMAuA+xvliSk6S8HO2sc6H/cKpuuMK2ip5c+xSuVSh0brJ
0vYkmxs0jmXAlxx27Ko/yJWbIzK27CGQU2ih6P66DM/KZ7y7FrzjpH+2l8QL840YEd8Q1h143Btc
t31ZovVcQWFJY5zu7JB7+BAGICRDs40nzWmGL8czmNSRnJRqQmb7CnXZtGcDgLIxt88mBwgO78xF
C0PyCqb8qaX4aCPCOxXNKh5RQUlESZPw+qluOvxrCl5xJw3eqkGjwfM8odw06DSTMDubTKCTetlC
eASPxMneBWJ8vwselvLF05m07JkJZZGCnbr7CEn0MH1tkxzYbHpz0F8W5QmI2XGsTYHo6mJaajSC
xQ3wJSwLYPR1Pgac1J40hkIrAhQefbUISBIE7u7Kt4qObhAUWrQ8d+EH505VmAuOkGPKTaDO0Yf3
5GrDt+SpIqZSUTDxMcfju4Hk1CUoFxSsvgWyC1OHwj2tC4QY9eJKVIs0CDXDrovnBUyUDhea1QYd
Kc3ukHuEoc0G9hOiArvW+MLNocmwbfgEJauFamWRePEgmv2aqbQ/igJ1lxEEoD0Ys7C9k0ryizF6
UpNrKY3bs1ZofNMMhrSBFvZTzSguSJqd2RFdkI2qXtQyyY63kv2+ghp+euB5H9XV5KEZLntG0whi
9gKJ5CREz778vSYJuk99VSRfhKP93oJZT/eXApLICVUs1H5lgprIpK+CywIBU0dHdkp55wjvKaoK
/tM7HIJ10EXOjR/Mi9h87bkRaak23b9/4yPMhyfgBv7J1rV8pl/3oS4uCcdNZDLyFw2HIDFsnP42
TP/xT0hRRPeB35WSIn1OpDLlqWeilSYwCKamC08fc9FnZ4NW4QpvKkktX/PkYm9QExebN9xxAyxW
POuoaurgo/aMm0E8+5ZGw3gMSZX0hMFSbrgmT0LpjA08n2BAd2u/lgFKryjW7pTWrru9pTp5F+7E
4BcF3FZ1JKchPvJdT2H7DsZ9dwQMn0yTxtONS+MHPvkAi8Xine38+w6I9n699WoY5QDfr7N1b4fj
4UaRKsg9jkqcw64D09vtoBpUwo+YlWBprBO2q7gTzP/PPPXkkDxii2fnFqwHlylpfPTV1iLGWyaq
LgR7fei4WC62dXou39dGm0FzKx2yaPnGGo3e/AZj44sITLzzSgnWCroMLywjMQ099iskPLVVR+EG
yTKFTNUJMc+sQHVE223CHEPDhKXyWMRKju2FJmOb5qEhS7YOoc6rcKbDUB1xBMgmpZjlj5AbdJ6U
/RqKUov/uR+2kcC1/C7pryWOqWO0m2gEDhbx0H3QKH83bZ0METsc3e2OGP5ulg4M++uPVS57QJkh
PJ4qxEr6Db6AKKgpqjOEfsdW4CtNt9PI+ia2oez3CDijeSPDQNtoQN7MRL8eIP4o6qU254MuJyML
0zm+42PVrlIlvEP6CLFGpLOSD75fztP0rSkCJdcnRlVt33wTZnTwC3LoPurqj9cpW3pclHXMwu4V
dQYJrsnntObzrkdztuzJ1ocbu0o1/DS30JNJNCja1Y+2OznWe1xBJXr4hfGJukjuMFayiv52PVOu
0mVhWM/Uug6sUSyB4N/xxvoJB0pjTqS7Zpb2Qz7EwPKGVenTlf+yneX1qeOfIaHrO7EqbaxHusNr
uT/qCAU163s36jG7mOXbCkVdmOrUk3TS4XZ24QUx3vLfH/mFm634Xls02M8+cyA+fWk0Gtunz5cF
bssZ9AGuWyiW9sQmJa5OALtWhbp6TYSg3WOMv8idhp/3R3RXsIUm/XL3xCfaslcF1LkOXrGKLZz8
BejvGyq2Iztv8w2RrFRW3tCsAQUI2tV9+67sihl7ZsqENEMVF3kxGx/0i5phnJKRnxSf/Tz90o2N
tGZ0DjvG88TRfCUuyuLphCOtFcx9OiUKG3R7ASFB4fApEQp5lqPUYaImh9Uq1LdDQRR5mBgP8dPY
TLz23z3DsSmg8hCqLtxdslmmjq6v3fkFvOehn5M3eVY4wKgDn1QiUemkDD/MAeowy36RI7ceUKVG
7w6FNs78lmrhUpPpgT8moNlco6mh/QIqtCZpEfJkxZZlaax8PirVZ4OVMIbd35ASTHky68LyP/25
XSJm85qqU9FhHsxDqG1+eNR6k/gwqbo31wyqG6thshCgYCWutkzHgp/iPNJ/pD6cDN7g8D2PnuLv
Sre2T3Kv0jEPVjfd6YVFuNfhpYVa6PBWFIO24PJzM7OCKPU2wzJepe/FXBmhhCJeexW+iTy8XQ3p
fD+zYO/k2d/S0pKBHHZ+1B9Jx4UAKz5cOvL9HBXHPtlkMcpALh1+1y4BeAa3GlFmUYHXAkmZIIfm
ZHdQREC8a8T5TF/nLN1SgagQUxlRAdhzDxAOw8kUmou+zlegS2cpc07xE5QblgRUJ5SRLYantZVv
9kw+ZXuwgInnQRXiy236ruS+dNFsGffDzvsVpw9oRvyV+CFnDMQv6+BCp+Hc/JzdF3c96YiBpvIS
5R7vxoWv+roOvtDPuTV+tMVmRkanGuhLvKbW7XKmxdSSimnju9gD7sNc/yzKsrEnuyQ5tXa8Kvzp
Ww9/+s3wrfeWRx7k6YjWdAiIv9HxdmA1d+jlaq/UD9ypy5vvYa/MoIrmzXrriFZ0tA6LBqO/yzQW
/yD4D+obgHslbY3IpIHGtvRtS8HTBsQMRHOMtUqEpWIBV74WvyuI/nH9SpSyijGC3yV5Bd/XgR2K
15fPlxU0BjVK+AA7QUlD+DizTsky17YHifH2/7PmoEZ1fw7syU4KPGD46xfIQ1nF627p3AUIM8Hj
9r4rQq0DPgSsX+Ql4rK7Zt1zL+wwJ8bYbVwYIJNKdXCnJuMRePiij/wmZXDzY+oAlZT6o78gj0vp
RXOVpgbQ2Yh1QigMA0RvVQ5DhXD5yyurgGzpEI3mPbrKTYM7Vpfiw5AojY30wUhivY6z0GbB96rI
/SiZWwwQqznnKbdoa6DT6bBFsCwOSrOaHLGvP4IuI0BFROn5do4P8CUrTXQBak04yB+EhH9BS3h7
vWgSkalDLCv+jmNlJpwxMNt0/oMwMPQRJZjPBmHzAxcM6nvxx9wsaHiImxMS20Dr4w6OKzVBRYuP
r+J3QnVhXrLB3tBviQyN5Nf/gVuF8X/BojUF8Rde4iYFOklqWMtmyMMM4Q6QG88HbAFwC/uSJlQ3
/nRHSJJXdyTE+drX+b/MOk5KEj3J3ZuEkSGMSQKRp28qZDNwbWmvXxjf+Y1yaj65vLQ85XYFZW97
vThMT3fn7wl23ld/oj89b3D+Fd4BV5r4/H4fdNawSoTGd7C7bob+yJm+5xmIFqOHsxPn+OBg+BT1
RMp7cscTvj7QVX64PpZLiGx5viZFrGmsx5zxs96ky7RstonYhFrj/Cb6hdjiYDDQe380E+A++ZLK
lHawwAl7OwTLqSIG/PgNaeTg5aBKxpaqQKKiG6O3LUfBViXKMhG4GbJRvW7ylvwdiAkmSyPLosgk
JS9mDxZjRDsUlXm6A5ijFxyVCkxiSQYWcXUx6xEzdqFjDFHkmC4bb+8p45obGR9Fno0Zl3qy9g6h
I7tJzrLqYcCPCIPlcpQK9AqMSoduMu4TVNrcOUNQ6puHJl2PGBDot7hbyJrIRJpRWa6UdFjA2w8q
g3zm0kJvjxdrqOMB3WTwm0fbTlSZWiKUoivGccsXr9XIVUMMoLz2UPsxedf95AMvGzHcT7xjYO2i
ZEtGYMTrlxi493TX3pPMqL76u5wlGURzaxZrOJc83cBGiqs5na1gYZrY/18J7Gu1hJYLDOKbIlgF
lgOYIcyVbh7m28WUZgyYl2LJZxVO6p8WO9Z9RLfoL+uyJxzbpfoL1yFg5RnxaSaTISnOiEHzKrbe
1ZOw58lLIb1NSVeAOGTsn6NwBJjWW5qE4Cl3rUOnTSpf7Iqeba3g1mDIo6VaXnpLyHwlJyKMqzOz
08NLUoQqdpm0s0CoWG+KIHyrbmov5VGnG+KxMOkzUUwtGoMkNPJJD52DIE6pQBOYrWSYscUXT2Nb
SP9j+ozt2j1ODct6rTxWRHVA92COBaMJ7NSkPg/SwCRwZBy9ywiDDcEpRPhEWu4nyttlAKi0YgaF
UMEvpBtNfhK87IrKcB54jCPXjjRqK83lpiDqF8w+vzWK+2yjt9mcRHFRc9EeJDQgmfKS7ypAxa3T
vs4cmnryH5eum3RPmm2pElPA6lnQdM9MSDDAWuodl6XDcQB+TzYrBp5nUp1OmXoLfVOkL+VTY7OQ
Zu1TaUKIuXOEKwuD528rghYbOM5MVg8giltWpSZhg1qVgTio3k8DH2m21q2gpyrdVt7cEvF/tUpA
wbJsBtIfWnAjQXwoP5jc42eUq1cF6FZsyr4soYABoXI8sTj3HIJgvl23/BNmwUyKBdeuGzM6reru
T39sBcXSj4iy6X+Q9czhWe6Mfs7laxOlA4lrzkSTbxzA9yYQRa8s6CFQrW8aMyBDFelN3H5x/i2Y
wWr2JtMVRF0WmIRTje+Szb2U0G7h+UlLLY36wAhy+6jV6oI9h8aOGZ4fzal/TOddPkXOmFaboUim
3gODBdhCMZI2jIQ/zzJIEyHTTiKafel3JT0UgjuGz4YvndFrSNoqwi4s80AUarJI2LN8JU29fg0v
GxzjwEmct19r/hWlIh3UWy9B6d2y7EWYuaiL/uaEdABK3Whk0dJEzEcBQitoD6vlq/Z1aisX8Dqc
etgJ1TpBraFlOZobqDC5pIrowJikfjKQSCV3E3dDXMs2yS/1xvMVmg0Q0MdIogzGmjZ6UNRnoDmf
JCJ9uetCXdUXquD6IlVJOhSbe4HFP+LqUQTb8AONThxU9cK/1lR3nsRFPYC2Ab8XlMa9GSv78SFV
jQyCbOknlscFvYMAoNU7fxVY2KJHh5YBRayD54ywRHoH5wqWbwXjKatL+zU17o6+SOHGsxQ5Dd3Z
8Lpz1Rtza2zb5qqHkZB29h7WEcwBNBHJav16qf+9reD785QemOQ/i8mA17uy7arQnNUgpBI9OGTn
CZPmzIbt41LRMhKaSXEAGCrbYqtXuzARVkItDjAvc+46N+DoUwqyEslLGM8edUSUfH5KNpGCuaWc
xBP3xMkT+8Hq5XGvZa0c4Trw2x0ycR2+odu2VNqWXdyTBbqkkHQ91vazKi5vqVuSUb4rPUt+oZDF
SbotRvt7BWd7EUYElJNgRQQrSmoAHP6JPmXUm6qtfh1kcWnBefc2fga9a+RdJIO4XVVL8JfUkI4m
+J0afWnbHFwYO2byOZyQmZRzWT/cu+wrHStDa48D6MubX2FkdfOxkta6INhR2bMqPGYiY6MW0r/6
Fz4EVxJTll7mC3AbS5g7lLiBbBGKc0QOzeXATEY+ai2yN0wJ6APD5Fb/YqG77zxVncKnBH8CkgWI
MRwCAOZjjmFAcGR13EChUjiG9tBD/Xvgfkoup/xB3Xllr6M9SG5qgixwXINTKhobnlLjfD7xkLv1
OagtN1B7uQ/2fjRNEpphHMnFqldr6qjGKHtp7uDv4rfOTzO5lxza3rX6eNHiANTrSC3mP6fOqdfe
iz/Kizto5aT0MghoL7YL2UWBkgRfOcbXjsnm1yz8Hac9TybhHnm1XslG2tfwsLqAmqr2EmKJLZgM
bY5Qd0qu75UizGHKPlk9oL1vZINsyeDvNswmDvhVqWCRuFScKQxk1gEn47oVJai5AEWJ0h0/hWGu
9rAK5D/UiXYQY2/3jrnsL64FbNu3Jvrq3sNHUcg7FeYm2p1UTQBaQe9DLGV9lvHC3NAjoyyThKnn
BjopJd/ojtxNNnXcWj2UIG9Xxvuft+Dv6GyeEOtZrlFteBx7qg85WjJ0vbPtjhNJ+g2Ceo7Gvt54
bQAFmJC1xQQfsBQBCKNznXmWC1yZmLlPBm3h3pRWBaCEuXXiBeXsRVbl2ofyQS9/7sfeiivvHpiG
KVovrtdPNs5fCkcUGMu4Vs2yBWGjvzr4jNQS4ipN8OlqcQ28RHeMcffvHWLi9SM6CEycxrn5P+b5
Ow5C4W8WDDH7XU9guBpS1FXwMMh5NARzW8RbM5hypaTDF8EH6lW+g+fYqUMGBP4pb0LZNO39jZhm
xEoQWNrMfUQXfT8fYXTTtR6JLtEFsiKVuES2SsFoY5L7vkMeFLgJKgsj4VNAy2stF01i+RK0dM1T
o3E/0ggq9aev/XdmWqAhWdiTvJXFCu/3xWOTL0t2wBrWacGeJqPTXVBbFGdmbElLMB0O2dmlCwtM
P+N5QBAzihoR7oRsx2I/374xIMAAcIRlg+SxR6Arvd8eaoTsTdxoJ4sp9epE8dEvFgXY3kadOz4q
PiKSNF24rZC8bgJJlNUD8+dz/YVLzD78Mt7Ix4ID97nwmTZBaQqw82iQ9wfLemQ+0/E8OU1uIqxv
7y0dXAWevcMrJx3xJM7zcN2W66HdXzNFcUhcEa+kYNiP6A4Yqk8leiFPei+7P6Oh8UnDsA3fHe6x
a49b6enkoe8QP0Hv6810HbwaW2m2q6UX6yccdstPFYZH+j0V39l3qr1k7WtXIs6As1SGE5KvIvVI
PIvUTz+CpJld/NY4/P45Q6oKoc8tx1HtI33DHieCkPL5STSFd5s86zos81sU6SlZvOmYPudoIm8a
ZA1sru37oNYy2E+sW/Z1EqMO07XgWBo0rH8goDDTMiCZh8Oh8sOyoUW4fWxQx/qiH/9+wPkgIrY+
Stfj7v71x+lHwixWCFY8ccXrM51tonNo0xaTwdJSXjIaznhb4z9BfE477VX1yz8kChxaqpWPlq4Y
7XNT/7tw00ou8OYx1UjDdjrSf7ZktkJ5+mZlcM+fpOsv3Ju9QLofEXBU55i7fxwNMU/lPOADSdET
tqMFl+0yu1UIIjX11Hhc95TlJ2HG5ueFWChmqgDd1S8HUWy4hpAnj+XqUjo124JqKPsWTBRIVJZp
cSAExnYBkVU03o1r1oiGtyslfNRJZqZwybqRGfX2d+ehIDN3QNGlpbpTIF4vnjq4k6VEPo+60EEv
EVpmndL4m3so8LgBWFCzls3KVKSrwCXrCH+3kef6Ymo4u/JwoMGABzDrOGBa3CQ4X4g5Df2j6SYF
s9PoQGlUaHJL3gIankcFF45s8JgKa60T6bBgxaLIJAPBEZgqjlnOV9b63N14TfCXfZuz1vcGC0RJ
niNmxmKWy/XeOpfjftDniJP0SoAb3SyRu4mi2N8/16sE2us+eaTMUkFdMbsm/d8o0Swj2Q1+3WAg
uR5hCQn/n73SE1KpIz0h15O9pARpAuDAtieb7x40R/v5jH2X4PkqOO9kQMlCSjRUwN+vaLrb4ICh
dH9pijZL3hkMuXJcQeiWlBZgCa0OnFZ/RKhq2w5z8HJ238KptmfJWFpMYtYgKd96pQNl7QeugMNS
9W46CzlZl4/EykwCCsx9bpvradZ8DI9ZZHu4fRZnmINCbDgif+lwQ1X4ACFhPn/f/WePUC5VX2zR
fHujg5zjubVJJVt8MnQQF4PBMhqqODqQCrnjEdIOKCiDE4wpeVmvWpwTXgjTksa+t9d4ZXqcBoID
5Bb9P41M0KHHnaIpCzu6YJVhhT/fhZlTXe5JZ1ssrHjxy3iKTYE7Zjv+4oAli43MmmFMHpp+hvAM
r6XUF/SMRElmlgVnx7tkdRvWsxdo7jMgB0TNJcG6xZ27tW4WmeNb3NL1BSSYHlumwAmGlfIfNLFd
K+HF1WqczqvSjH1JiZBwgAp0LhxPyAEykPxLoaMKqhr5QpsxwADoKq2dCZXhQXxpXHxPVWM78QHp
eX6bfg0jHe13tSAX6+Ll+Xvrw1HCoq57djAdsiMPF80Wqt64janPCVsVNDKxjj9O1bf3948vqiNl
rZh5VyDDhF10auZr1jDvx1ZBggW2L45UX2O6uAYXKTFl+GAFUfWLxrsNH3/TVPB1tXuOgLjo4cdS
bBCHdmsaFnIzWNV1d+S6n2gumNcLgpAn2JDuzg89i3IzSIra7GOVC4cu0vm/0Vw8l40TL+lHvn/E
ELsNueWGW/m+Lh1GbiY+FRvTENqaZ8orqhJNdqw+gHl8UG0d1ORbb7DllKeiTaVfbhcHmgUbNrCD
Mzspr24Uq0m4yfdYUJ5+FlQtX661STF5GdrzLPuIELNLSNFLDUeaNIkTiNigrKEkoK3VCDdOiHQo
HCTLwM/2hO1gqsfTHzU3l5zXrPaD69XZag2Mn1399RslevsBZs/pJ17Lev2CVERtPHQMKUnpUBUz
Q7fEPUZ+wZSZWReb2mVaZCP0SQSUYD8BeIXOhQf4f54BCPB3SjyBTisykqh5enamIw4AM3oqg9E8
wPmYtyqDGzhzA+nYvNFdmXfyg4RDS57xV0CCacIp5Kd0QPrySzNMBTGvxJOmv01fKaWf+AsmvX64
2dl00iUmzQ4TUy7f6IRLy4f84qNP/PvE3MCDKeeWYK8aOp68b2/0/KOsl4MsFlZYYFE9Hs0MblXk
wOkDZYtyoiLOPmVKB7Lc+wpwlUcimJpAUOZdTXyuBKsG1hktIiSphszfBtMd/08SMD/ItMxFLPqY
28KI+6Ve6RXe+qfsBhHsMwNdnVsIKXziaHeMgAZTLKbRFwCdiEOMRlxxTQIFWOti72sJsvKke942
xDgPS8iA6yu0gTTSJbe8ufwoQiFusES6CdqQfhGoI2XtO1y/ImWg21rxtnQFtx9wtoYdTehC9gIw
6L5uzYvWWcqxs7xPmerH02Q5Dt4kXHJ5+rkPr3KrZmgXzSntlGwLNAyuyHT0aL8WLAeRZLHL2CBt
LGd2KJP5LOqUbJJDN+8fhx2LNIBWXPuR6qtsLnLTut2SAvsCtCTrGwbE7jnmVVsOtovPkHhvZDWs
tAtpXGdb+qoxesWN+C8C32uzzLw9bBnCMDRFNy9M4jMAB7ewIH5T4IN9UH3N/GZMrl4P1WKohv5z
srYhw3Jfv+z7wJDWgTntu4Cw/XMlzAKFfeYbiFWebDII8ObXeBjus/KSbkb2ofGvD4qKU78WA98a
SM+uVvPSJNC/ptc33BXzQ41DkCDa4gnzor1J9dGUzVadmYXw+KKc0p7+UBqhIH46zeeeFYz4A6Xh
18g/gVEjhgVjTDyD23Ue7UHqQSa9F0xcfKOEgLBEmFfVfphD4eTnicJdo0LqqcGtQtgMUnbT9Uxd
TyPWwEK9Vguf1CQz+CXh+uXLbdXaEpvtA/yy1vc5fAjykCWYQGuUtSA9XH2nq/g/SuoCG5hsrE/7
MRqp/H8UjhjP1LBMnWQEGwZc3zyJ7wp35XQBxNuMaUZ/qbCgJChqf3Q3Rix0w/nbyK0I7veYOHsH
2eMoKlloI3Zb+mZN1iGoSd1LMuNjgX/REDw9xLrO0vv6wuPbExQ/VMS8+1mCGbyG0Mxa7Prhqpmc
6Wj51ABw//3GIn5bSVtcQZDhUkc5AZweyOrFQbjZ5qgqzHF68HVz6/S9z5p1+RV0j88CNZkfmllA
uLuikLnUDL871n83ceyzkCAFxtnpd/8nvdHrDoWtcMe5psBKOXURNZHBwLVmQU+rekhKHSuW5YOr
KRRnClMiJcsojJsvhcTJvySGQYi8xKYhrX+dbLKIgC27jPRZUAORT47lUBHu+EiNRRyd0uIktLoB
6xIbcB+hSWeZNRcIW3gejl1MwoUTjmHflJbBCfXfpPCA2xY0dhsjr4CBOf1bgCELqPP62usjy2Xa
jeq0MxhyJVC7L7TI4Uf8NAIgHcKJF45LwddvQfcxkTrX5voGpQxY+Sg7KJcrCGZJ15DDLsjRc/4C
ldHAXHXp7CuEtuws0ESYtLIBdGSTv1oSV5uWcVzw6vCRfYUtHJnUakZ9gfo2l6QQcsmRy+WL1epw
cpRTlYlmvX+1RujUC/IQPc1Uhvs9vLYrwHuqDQqYgF8pZobBqvKI52cqRs0fGQAVOhWBtUsLKw5M
kpOsbJ371h5DxMG7jFQqI3xYIsmjEG8VtGh3NGJibnH/Xsqy47XFeEH0liD4A2XeQy/t51ySmqyM
vtZTId0abEutCqkzM9Op988K5fhX15ndmMTtdt39xbpg3Syk9TLXfV5/AE6gUh3xSz8ZdnDz/5Ll
3LsHp6XOz1gYdA3sPztO96sMTEpT+rhi32azMkHicrCV3hz8pev6vwvYdcmXn9A4WeVt+IuWUTxt
tt8IEQl75+Nd0u/5T1Bsjis7Wqzuo3FeDQHCbMVRunWbIJGrEb1ZW7Q1hjCeA7ymGUv6/8EFAgjY
4V3MHheC7hQHJm7a79wkf/1R9lsa8VsVgN+o4ELg+jhM3QE+qtEANMrSKGvF/XlllleBfoH4O2mX
aQQk3fX2NP/4crKp3AJpYnvWNkkGlVhDuA1GoXWInMxHU+6CtyYrUj339IWoJrr+LPcg+oFbAUxB
cmHN0eX7xCYu3mBTrY21/SpkMbG8WrSFmeh9TICVo9WQ7wPQw7zjopTot2bb5Np3p4iftYc4Uxtn
2j0JdQVFKb0C9U8+JJqHy0FwU813cQ1VdI/AStYki9PmpnShc0vfYvr9re+YBLU/XSYSPF/aWbpq
yvm0uB+mF7is3veUOYfRmkYf7Yi3VA1dD/0IZVJZcU1rB0iiwnca1fn1ugOzxwXuUCSogbNyPoXC
X+i55bpx2BEQ2KMFYoRyf1S78NvT5nwxlbeiwUyZq8PDXNDcJwv8ulT02fBJrVmwKMOqFEAaRbxa
N9McKMMX/SGCUwolrTjqLMeNqsnV6+eo+S1wIlniMxlhCVH7p5Wkct1RGC4ksUbXGhCDQJwqdUGH
05QRv3r/2Ok6GfON7SnlEM5yQrbeQt54yV8yZaUPWKBPZyyFxBnZemeP8PYEVn/Zra6jiZPavqkg
Aodjm5TS7BtnUeZZTWSbfMD/384U60GQwvFH6ori/KZbWgqUhbZiNQOgfwgtEw8FQ+6AJPC/eM97
JI57GNtf6lp88IUePsZXmSV3fnd6n8dIULhIsF9Nop2v50mtc7trQ7B6oYMvcY4mPdBzyYSgT8VM
0Wgy4qj41g/ZHaV6QGFllweb1X+9EjHk2rV+s2HHwzY9/Gs0x0xWh7WyV5p19oHt+xvCFDJPcjyI
pB/vlX2nHbhxR2EzpF5Cv8LAoes2hH3Uup8k9JD91BMBzuijvaJtrnR8U2uB5tvAlQ4JSn4OF/10
p4tMSIlgQqHIBb9RAXX7EMGWRqtj8hDHqPUnPZPvVnzq45dARGzC6tBCan5AKbg2VZukjPhdeufs
I94H9NDSDLzVqC/tHHCRvVgOZ83m1rdvJG5mlAk0E65Gmx4HxTZGPIl45cMpP+BrvBNZvSmhfzxA
nCLz3wgAgA+fPdcwaUVhE6XvsOWVCieF7P4P7r2wOrd2r6TyZMOIVKIJf4ZTHJ5/CgOAN1eR+56X
Q7KPRrt/nWABg9qfb8VpvCSzVvtE1yKuth1qTg0hf8e6iMf/pY3VBwHVkbMylxskeVJdnmw85Lsn
NCZuresyIqRTEI83WuBXf8ver70c4iCSK0wCQ/wwL/nHphyAPL9gSfRFEc6up3WfAGVEtt5Q0Zt8
xDtBFugFhWdwn23ewuTL0vQkBPy0GYLcso6lh9oD4eB3gPtXW6JJRk92lJLrBQDsBGjljLWjepQr
HyxISHKVkyaqhKrbgo5+7tKQKnaRorRWhUj9BjI0RXS4ySE0Olp6Wx1jU+p8zcrAuvDA26A1Af9D
Te2y4gQDMdpt+hCMJbqzHwev9bw0biiI2+0W/ZSjQR6srVXOzexTwD2Qn1cy6Srl9C98AcEdGbde
JPgdGCWTIiyk676pumoXxc53lt4hLRTSZRB3bhH4jz/x7OaJg858thVFhjnfHe0rpIboM+7BzPIn
sw/3ppioXZigl+1AopbOfYGjoHzjtHBoYVj4h7rEveNPVSYdBVgJUPYaUorURuaiSRRRC/pAVLGy
SxxsJyX6osB3OJJ1WgvE+DBq++Q7TdfwFWMx8Eo81YeT65mgLDG+cl1FpRbPBce35HX6x5E+fxO+
mj9OSdLGa1ruKnks48m8sLUGnO5eRpVlQexvdSFqbTnujI/7TknZKtlx6rjRUa8t9R8sb/zv3gGH
tWvIbVU3wVixO1I+HCeTMIMqY8BTD1bFoxSIeoxFYEEYPGvpadS8G7d4aUJvFRnUz7x3N7epH2wW
pEJV+m2fQuITbIyBQYVz0q8X2/pJcZfcN1m4ce3h9PH+DNHrAzUilwRdM10SBvAKqNw5DBhL0t37
JXG72WrMOqOb0plxnhtW4BMYzOBcE/RWB0qyweHgEliyKJJrCr/K37NiyaQ4CAbTnUWV1jGk3mvR
X8/dnMoyEaE7pXHkLOxqYSl54oTPhjrY8nUOe6zzJmC0gMgn9g//+/JVJQLGzos4hblOoNQ6c6NR
0o5MwFJgqPfmS74wPUKaosuFBh1KOLnTTn6GNdRqOVhw03IJi5UNLjbM238ZTIMc4YLiSYRtVbMC
Cwz6Ec1m5TrphU4hPHesqctsGvKKCIly8Hh12tcRu6mmpE4=
`protect end_protected
