XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��
�������z�(��s}��$L��"z�o.$���hT��qR��<xz�����|�&z~Y/Rfc!�����y���,ݚ�u^\5����c�S���Ƀ�2N��Y�)>��=�<+p�'{�f�؛����k�㷃�M��-��󿡯�ё�3��ZQ�1����f�f�]�-�"=�T��{mh<��5W_&��&펋9
�RŮ{6��,�T_^4EW|�R���pe��"��l|eBF��3y�R�{�D�� �	Su�"�z>�i� �cď�#Y���y�+٬�mH/��hZ�4�"L^��)�$]�ˈ���5Ce8�<db!d���[������aժ)���.;mg��ѝ�Z��x8���7$�+�0��rR��*P~c�f`�&��w6؆Y��RFU��h�ݳFaL[.��L��1��5�����N�H���-�[VM4ѵ���JF��Ćֳ�Fӫ��8���0�\�=T|�|����&�,��cm.U�(tK���:z��#�zŻm���r��ޛt�e���Ӈ���q*�Q�}
	�W!"������`(�N}n{�\������;�a���[�}G�1<L��t �y:��CV� Y��p��ıy�g������o\uRG#;�5�^!���t�ޱ������XS֕��;��q"�5�ޙN�D0�"��IOPz���Ԉn�@%��Ȏ��p�<���H���'S�X4��XlxVHYEB     400     1e0/���o����߃��}E�(�?*�XWx�\ڀ����X�Ւ1�. v[L���:�WJɘ:�Ն~Q���R4~7S�+��?T���W�.�,"�3�����i� �/2��AB��#~L����s�p+�<�9;�6.���Qs��5�o��K�"��8�q'��С��0o�/=b!5`8�*2�9��m\x����B�A�E5,*�J���(�R@A�
�6�B��(gм _�,���2�c���lR\�]�X�Et����)�H��n|�r�]!���M���Hd[���@5I�m�	xr�/_��Z`|XR|y���C�[�bw7�/�*l�wз�N-��z~��6k1��dc�����,VڿJ�fky���cϙ���=�N���#m��&�t��D�(	��a3�P�^a;%=�w5#�L�S���5桡g�p7'��@����(��H1��^5�J�P�[%��{��~�=��c����XlxVHYEB     400     130���6�٨�S��
��tP�o����k���+������i�����vz��8$YUT�^%��(�K2K�B��S��ʡ9�%��[E4"���gCu*�PD�#�����ϻ~�?0`J�1�t�<4�|m^NZ�fx!��A�֘eE����ݨc���m�q�#8�+�]�����W���Ѝt���^⒦�{ {�2Cc�:�x9�30PJǮ�b�u��Ov�T�cb�}�f����r��b8S��|1�hQw�L�0������w���F*h�}g]�6�bWL<YnR$�%Vf��CT����.�L�P����i�XlxVHYEB     400      e0��,���p���)�*��/Y7ֺh[ݴ��-��Le�̝%j�����	�iS��}T�#-p�d��3w�$��>���(�;����J=��������@�D]N	�.~�� A	'���l��I���S�J*	&?���|����99�M��#��q�<�!܈�!cr>}����r��M��$���1���[[H��7/�S������� n(�W*XlxVHYEB     400      e0-��_���-ah��B����>�\�< �u}�Y塙��ٴ9ԻM���O�|�_�#��OR���u��xwP�oZ���:Uy�
oU��@��tw�a6�ס����Πk�#:�4�qJuy��r���Rȵ%����W ]����'��ݮ�
L����s�N.��E��^��*@�}z��`��;�[ =��_<�z��$��CE"����u�����(8K�fpXlxVHYEB     400      e0[:~�xO�Ɍ��_���a0;b���O6�[�O����|�a��Tܤ�"��qT2��.�r.���y���h�F'��f��0�y >-q�u��ؾII9���[�������>5�9o�멛XR�?���cy0�C7�� *2��U�`��+��49K!�.�1_VX�$+�!�����P9�6�B�a�E�P��VDz=Lãg�[XlxVHYEB     400      e0��T�hW?(G���PcQ��f��J�bc�R���W�cՙ�X��"f����	��ҿȰ�x���5J�h�nN��O~E���b�i6\�A�_�"wdM�C�!|�G�3l8+��1�|9-�u`k�����L�&��]N��^t���U��<�|O9 @��fxno��\�@F���pY�Z��%��	��Ȏshj�F�X~3�'��	���q�t�XlxVHYEB     400      e0�!�T�Ub�5���VD�V4<���j�I��p�|^J-�pW�֢�f^�/˃p=`v��߃hw�1�����]��Ώ��̞ �<���2�֢b�V䍻�V��R&UJ�t��N���􌺊�����$� ��+�퇘� �.�ރ�R�"�"&㩧����(2�A����a��|�����G���9w>��
���N���ڊ����ˑ�1qdf� E��J8�RQXlxVHYEB     400      e0�����I6D�����<C��ԥ���ೖN�3Q�H��Ucj6��2B��ݪi��tǔ5��[l��=�Gܾ�!W�L0��nS�",ޑke����$��	�p������Kw_���NLTl%����2u��2[��_&`�����.ʑ�r?Ͼ��"���B�!&Vb����I��>&L�;X��N�сB��FEUj:�e,�d���l�K�����ady��XlxVHYEB     400     1a0��Za�aTB��[�k���[�T�c�-|f���)��${���]�)�>�wK���0�x 	J��^ �J��t<�'�!�,�%�	X�ve��l!�Ɇ�g=л9z����>���éJ�@��i_֝:�H�s��u��&ݸ� �+.��^Z��oO~����{`Ȍ�*�:)af4d��AY�)����ʰ7�y����c c�~@����Y��� I��>�m�Z)Q
b�'�9��~ǟ)���Q�=�:{+��rV����G�i�&�>�c��N������ >9���2P��Gق�p*P��u���#��Λ�e{��E9֑�x�LP&���� ���[��(G9�Cn��*Y-��/���N~a3#�k��eۀ��Yz��r�S�b��)�D�c��� �{?�,�-�?�u��@-�D�J!XlxVHYEB     400     110��ᰆæ��8һ:lPEFR"�np���v�,?�>�gJ��n�B�Wq*7�c�m���?s"�[�T�>���M;_�h4?.O�ZF+��	�4&�J�\�u�c�;﯉�ʛ�

�݌T
D��X5�T"��i�>�����&�"��T��)�	��_aYX@�)��i:�;=D�s_�{Q��2�I(����s��,��[uѧ%݅W�4L���Pħ(������MDR
 w'�������n�EiF��y��$$��7�&�!#�/������XlxVHYEB     400     180;�rݤ3-H9cIG��(.��v��`�pr�x�7��d<b���em�$k�x�;�?%�ePVqC��dT�%����p�Ӥ��;�y��`L�"�򿗠�Q����SS�A�Ƚ��mn�G�x�>��0s-���/�L�_&����˕��tl?���?L��q�-[��5�����t���@gdb�q��m���f�|�����{��x{�i�Q���I��	�V˚b��|rBV�^�V�q�҃c��@�u
3�${�a����%ż]d�pI`8�l'�����]�5)�w͉���eX�(��R2B�$�L�z��֟��y�_���h�i���[R�fҕe�7g����|�nv��@�R^R�!jp%��r�XlxVHYEB     400     120�͇��r��n����}|F�nz}���/�@�{֮���(�ٺ�ib3�>{?՜:�����3�$�kXd��B_ܿ�,-{��,W�aO����qbxۻ�P$��b|w�)���U;���<�x��0�:�HW�x/8�G5x�%

�n��J�0ʧTm�.���l�z���k�S��:�R�`X���Jh�M�����`Gdt ���w���.Ю�%�̞_��yV�/0�;l4s�m6Q/z����D��(�>u˅Z�D���H�V�����E��e�wF��XlxVHYEB     400     130[�S�핷c�7�z����=����m���a��|kઌ�!r��m�'���;��-�
�'�����?>��5��U��/���jE�{�Y��rв& ����ڳv����C�}!�V(����N	j$9�-3&x�B4��p�����y�_M�W�����(��Ci��7��	�v�D%��Wo��rTV(U��!�rIa?u=�uoo�ԥ��S������H�t >�`�ve��|����bWDz�5_g�ef{��JtF(�o����-����n��/�f,���_XlxVHYEB     400     120��.@�*[*�v|��s%K�R�iN�7���p�Qn�e�3g>�1a$�d	^�Sāe�
nx&"c&9���gð(�h����S��m��˕���d`--����q#��"��l�%r*^E������	���O���T4�����>[��^[ɴõjVڦ��YIo��.9|Y��\�t���eթW,�n�߉d� �z=?~��aM�b�r�G�s���rw�Rb��hZ�����Y!��D�T�@����}0!�v��<�S3ò�ćjo�����	�&Eo��e�_:l����X-�XlxVHYEB     400     140^�s���P��-�}%��d��F�=�c𓜬�wCM�3�m�5 (�j����z͒s}2�����&����f���9�k�AAU�Y�4��dzMDzҼ��(�a䡉Q�A� Z
��j�T#N-��)�� 6]�݆?ZF�0AP���A��LF�͐�) �^sJԙnoo�a��+S�*'�I��[�7gN��J�N�a&Nӌ����S�(z�Q�E��(i���J�Qj9�T<'Q���l��:����K���� �I\+�&��5uˡx�M7&��{��΢:��W��a�5�dpa���>�8	cA�wH�iEh�]�XlxVHYEB     400     140���� I�����ǅ�ҧ�t$M�����(���,A{�\\��������}$g�;Ɔ9��V��1��C��xn���
3v6Wa�چML�����>�c:s4���
x�1�ud����L�V�)u	��|���N�S�3�c�Q�Z�����u��N��.Eނ/;���B�Td�A2e�ޞ�v&����nj�O.�'q@�ZrbЖ0��p'�Mq���fkow���i�,4�>�W��7��MP͇�S�x2��� �W�ܚ	����;��v�1�'�]͕g��HR�ԲB0w���Vq��o��![��{XlxVHYEB     400     120�7*�n��u�&l��\�!A��a�b����w��QG��X�2�?�u���1	S0�D�����f������!�i�
_�UZ�l��;�1!Y����ɮ!�?Ѳ�cH'�\��J^���H�9��fv,-W4c���!6m?���{��x) }� ��儞�_;a��̑��r x��IǞ�Nb�՟2A�O�9w�I0�V⬦�=���\X����,��乤�"N6��B�k���6� ��ar�)����k$:������l�ƛo
}�R
�;gB_Yx�DDi�XlxVHYEB     400     140d�v��Te������<,�pS�i���b��h���rt]��V5ɂj1���'�ٚ[6«�Y�sC��Q�zܓ<1Q.�/[L{&����4���QM�ѵ��6s���1%^&�o�����@�Xiv�"�,u0$�,���#���^ó4L�3��{�e��Nu�nd?j�FSu?�K��G�"�P�k|d�<lr�"&��-�=��{�V��]FlT���k�`�M�Q�Kg���@�B�:g�LG�r�Ij��	2���X� ���}ST�4|�"�/EAҨ6qC�=�3���h����W�\�u����&;���Q�tXlxVHYEB     400     120v�,7�JT�Vi`�J���\�{9�t�e��lfh�mnqI��}o9z�����\���Ć��x3�y���%G�r�#_ViPu}Zd0��ӎ>G�B\�gJ��iY��a����r��Fk�Y�Q�Z��+���������w��a��v�kT�HMR[ru
�����JIG�����*��[q}dٶ��{�<���`�)���:�g��dl��\�z����N#E�*��{4^$�orlx)a��8�rw���E�6��r��{���<Ḁׁ�]�/�YXlxVHYEB     400     130�)M�A[��P�7p�RP}i�@�ud?Ҧ|�M�'Ȧs�4�;Bߵ�V���`��Q܇Q���sD�|�?o�E\���©[���݄J�c�kZmz�y�X=�r�P=A�1�X+3��������]��ZL��e��~�o���� 	4~�]�a��P�q��y|�1)joEK(Xڝm-}�5��-tL�y�T&�Г���i�V�-�O����I��Q�F%��2���������OҶ�pi�ׄeW�s�^i`���z��"��,q{M�����oZ]�2(}���NA���X����ӭ����_��=XlxVHYEB     400     120a�����1Ԕ;g���&3+`�|T�</3�	Ʃ맲{��@��O6O���-]��`BH�oi<�����XN�	h��u��ׅ���`S�����#Hٌ�_��BF$�Ǫ��)�Kb|�z���c!k����\�i�(t���n��֡�q�35#,W4V��_��oL�U�vZ�~�Z�*�)3Y/n{�{03OY���R#���(�}0�Ћ��:��(O���Dec�Ԏ���bV�/_p^D�E�irMz��	�`��Í������z����RR ��H�> �XlxVHYEB     400     140�Փ���˳��a��?ؖ5�����>A�A]�I�#�6h�ZA�xn�sԶ
x�.�t-b즂�����`��|L��4u�|���I�B^�!&�}*'���N��=�HV;zu2�:�5��U:�r���Z�L����E����f�d9L�K��և�Q_���'��Ō��!��!n��ݛpGf4���Jw-�z�ŗ�ܱ���B�h�rn
�tq��6�Q������k6s8^)�	��#���o3�O_q�߂6,���PS��CB�a���i� �{�O""��fn�f��8~';��] �� ɗ�gu�XlxVHYEB     400     140���� I�����ǅ�
��9<�!
7�ݱ]<ܨ	�J+!=��M����@lu��Et�-zu�:���ܢ�X��(3qX�8J��٩A�x�Ѥ9��u�[�&!'��|ߞ��?e�S��;87f�?��Ý�|�	 IE���:�Ѓ_*[E�̊������5V�JWF���@��s�Κ_:ENJ��Y'|E+Y�����x�m��1X�_��Fz����i�,���-e�",T�y+��F�d/��ѕ�b�����Vn��`�5�5N�h��D��,�9���k���Ս�h|�4��z9�[�8�g��P���׮���z��uXlxVHYEB     400     120C�@�jB�Kǟ�E�~9����X����N�K��f#Hjd>���Z���Ơ8�����p6�����?�L���� 6�+N'�|"��
��̨�����S�p�W��{_!��Qn�)��\�&�W�r2�t"˂pSh��JǸNQ_��3��'Sn�3]�������?}BC7�lL�� 7�)��f��:twg	��x���
�{Vu� x��vȋp�ɤ::¬
�J�� =���^O�xQD���T.�P{�حG\r}������d�����Æi�eKpXlxVHYEB     400     140Ǌ����U!�c�e9j!<�yZi�����YiFB�T��"���E�X�8���Ck�;?���*+ҷ4]�.]?K�"G�M����&;rr9i8�␬X����Xh����N����Axi�z�t-%��A#mk��)�gI�C�P�p9����� L�3�yƹ�svW-JӞ@E��̼e�v6ŷ�9:yF�ݏ
�-��ؠ"sS��w��j��Gϱ�Yġ%�#�5�����μ{ߋR�F�C�	fA��I7���⢤�muE}_�3g<�/��\~0^!�N��up�XH�-��z��z�I�XlxVHYEB     400     120v�,7�JT�Vi`�J�H�f�&���O[3;
]��V0�3�_x!��j�����-��,�rW^LF�P���ku7���P��.�g���f8��}m�1�uy��,�3J�kL��,������1Plf:��=����.0#|��Vf�ݎq��W�@�=k1_�9CӴ߼b�#��d[Z0L�\/�0q��Kɳ�e0q�KCa�&��y�,��{�g}H��g�y�}D���R�-5^�TQwp�dz���Y��`tIO�B��%z�`r�I�%�l4��,mX�u��<$XlxVHYEB     400     130���g�?�	��C�Q���j�*��ٲ�&���=iʊ5���L/$`��5/�G Tz��� ��6���柗�*��|��¢�)�d	�/D�c��(t��߬�0��R��NXV��Ƀ���3˻������~�YzhtsC���+돸-�	Z�(,=36G�vzU�r����{������VG��~����(�5��+�q��PфK~���l�C ��I�������XK����vF�<(̔�G^
l���xFZ�z=�|�|����mII�_3�p��Ix?����rV.�"��(XlxVHYEB     400     130?7F����X��|ǥ����B�\�q�J��P����-�xSCó��� �	+UކtF�(٢�}�C��ު���A{����T	J ����k�'!�C/{�ӓ�~=�{WK8c��#Зnq�)w�����mt�x��^cݝ��6�J��T�Ϗ��$�QF{)�"��nr��`=.��c��3
W��	�� &
��c��+/��W�L��$�y챗yf�ǤYBn,�A?���S�O**x1E`7L\�X�����{�#�A��$ �b6�h��k��\&���j2��М�� �Gf�XlxVHYEB     400     140-���R�{(��X=�M������Mb��c$7�圖ފ�hω���$3R��{�X�ƽ�����Պ��5�v�濫@����`�<Ǧ�� "x��ٲ>EuS��?�pWwuFz�Dfy15ء�T#�s��.uR��_�11H�Y���C�4����L��̡p�^:�Qܩ}/��P�MU��ݹ�F��Ţ�$2�!͂��p��>J����i���mn�ĽU���7�tCх����a�B9��K�v>H~	3:��ZX�����(��ʹ���y�iN��� �7�j�U�)��_�w�E�\��S��	P�PA1�XlxVHYEB     400     150���� I�����ǅ�O��I�8k�ԊI��ma���s�_�K.$�Un��Ǹ�w$:��F�7;���\�l�a�K"��l�aK�Z��x:�o1�=?��~�4��LUy���p�n4PZ��k��-g�1��qb�����I~���_�Tn8���d�~F�l~�+.a��(V�ݙ�#vO;��9w��b��!0�`��:�eЬ�;(����Φ�m���/K-���:Y�)��
��ЃU�nT�mb�ҎB�ŢH��Y	�ƚ�B��/�^��nl��`��&�`֌���B�*2�d�Ͷ.װAǫ�iᔿ�3>�F�[�9
٬TR{�W=XlxVHYEB     400     120��fkJ���y�H��7f<l+?������[��T�I�l���uc����pAk��U<-�8Q�n��_��c8�"���YyJm	�����$\&�8�?_*�ݝZb�������9�|�	�_�6�N'Yx��yO�Xӕ�'���4\٩/Oo���ו��s��_��E�y�*V����[n���rs��3��G�d|+�-�ɱ@�ge?��j�"��f$**0m�G�7�W�D���s�w"��䔝�٤lHE������℉=�E�ed�?< �˒PB��xz��l��XlxVHYEB     400     140<�֨���ՕqJTa,,�xѸ�N~a��5d�����>�]J�mW�Ře��뻔��,�Z���_�JH*ƹ�r���.��Z�}F�r�Y��|���5�@��X26���� ���rO���\!uG>���#�H'�$ߦ
3g�&U������/4Ili��}�����!�������:�k�J�P�!�_g�-h�Ԡ/g�#��s�5�8a�\�a�T�{�� ^�N�'���Q)��fUR��DA(��V�^�;�>g٠n��B@*f�T��bEy��ݶ��m�u,��8��� ��(0��ݤŽ��(H��XlxVHYEB     400     120F�ءz���:cZ��[<�U�0�t���C��4�3�j
�O@ۗ��)�$�<�^W�b�O��m뛝3��vK�p��!8Eg��R�'#��-����bcT��̖�� �pF�0��!~�����2��^O>�*�Mi��J�aS�Z�|N������0�~O^��ų�=j	9B�A�,����(hI[D
��-R��ʔ#LE�A�x�
���.�='q*����[_�9$��D �ǝ�Q�1|��1��j\��ҁ/��������':������v��� �`���*��XlxVHYEB     400     130�)M�A[��P�7p�RD�i������&�P�ff˚����IJ��<0�&����
���qΡKu�M�鍤l��,;1?��G�{��ft�I���S���ah���4P�P���z��-����X�Tlf/���/�lhhPԺ���1�tF��+R��0nq"�,�Y�r�xL�s��g�~�/����6a��sݲJ�f��`� ]��r�F�r�+:��)��Q~!u���ui4�{mwS#�����[x_����������O��F���S�Yav�6��>�U+�V ��F6X%�qGx���ZXlxVHYEB     400     130?7F����X��|ǥ�C���G5`7yi�-!�M:?���0� O>mm��c�� ,�� ${�A��"=�� �����rI�'���s�k�`f(J����8��B� +�����8_H���]�7�I��`���$��k� 5�֒�%�=��oK�3����Kk�5�kD�Fl��a:�ۿ�K2 �F@8��VH�kÃ��x�dZ��x�7��~�;+`�A96���Uz�(�TO��h��i���{lkq(�?]@���	�<{�Nod�8<�E����J�:݂ʦ�5��M]����`@$��XlxVHYEB     400     140ӯ�1��[�Aq�ת������ˌe�H����WasG�$�������*�Zh)�`�9������1�B��Q���^���⡁
�ڑ)xÈ�� ��,�%�:\5`����+�h�G=f������ ā������2����eX���y��yޥI���TǮ22��Z�zj-ozx���h�O�P�iG��@�,|sà䬭q�)�/��y�k6��׮�Q�~ퟩ��M5��9�a��pA�"U�� ��֩z�T��I��\����=�  �A�.R��s|�l���t-=i��	��)�SDX��XlxVHYEB     400     150���� I�����ǅ�|t2��Z��`N~���|J����H�zn�T�f�>��U ���7;�A���kL��W���bᦒ��mb���P���\q '��m�-�ۿ ���.3���:�6�xZ�����UB~v4j��k*�-"��T��M�>�!m3�e**B-6��l	����u�u���Gr_�辚dM��|�{�?H^�SObE/i�PD5��v�����U�K�� �J��X��&���j�x���s�X^=�e�l��t���/帮ӊi.�6�H>~K�i���~J�D�5Kg�t^_���uO�=O�����7���E"���"C3F{-��$#�`h�XlxVHYEB     400     110�}�:��Y8�����%d��Ã�����5�H�G�r�v& D\�P?THC�C��D���fE��FE�k��d��	2�Ⴅ�$�ZH�y�����( h�,]T�4l�!�Ľ#+��'��̴~�n	�8T�*SR��c�4���Nz&ě%~��e���|k�Q!͎gj	J%��3�-?�޳a �w^�׆ъ����A���z�Yx�F ��������N�^��c�y��X�ڿ��K���JM�*�r"k#pZf�ʙyD���j�C]��8XlxVHYEB     400     140�:�����}���?TMq@�c��-;{6Qdb^���C�P(P!����f�r��S��u�2��{�jO����Vrk�YWhŴ�#pV	��@$l�P��Ϻ����%� QǇ�Τx���f$v��C,e���NefXXc8�qH_��դ>૒@'� ��˚��
��(Ha��Uh�?:��~�ȉ��D�:F���o����N:� �0�<�#�jr�@� ��I�K��HwG<�א�����~�q1�3�h�#�'ZRlr����k3�]���U[��%���O����t�X���7d�}�4��*XlxVHYEB     400     120v�,7�JT�Vi`�J��"����hC��V�}০��l�]\k�mrX)~'���7��g��a��~��2ىr��zY��I����8Bnⳍ�ٌ�PI��빶sǢ"3��=�\��x6�o�%Ӭ5>��(�2������#|�����t<�CdW)����3�W[J�+dF������4���1��+<�t��.���'HTi�nj�E&�� n~��ϵ����3랻�p�0\��t��J(�����bQSj3a��z�@)��ż��s�,�f[;�XlxVHYEB     400     130�;�`6��[7�~�Җ��D�I��V��鬎��|ñ�k��F:�6�a�u��h�����K��By�0M�%��:j��1i$(��`)��W�MI�_���Tz!#�p�ݳ|�i۳�x�͖a{�FLGn���JT�A�t�%5��H��)�����iR��m���Q�Q�Z ���$�{f!^=�a������ضZ����ʚA�!J\KZU��6�@V%��ɝ#<��1�0b+�g�H�(3�Dh��F�ZwZ�~'o
���3�[�=��3mg�x��i�'�ܥX6|�z�bLL{�;�!�S1#��l)s�ȉ�XlxVHYEB     400     130/.VK�&�ZW��� ~�"�j{I�&\����2�l�h�������3����11�-:��9����`�=�$��+=YY>�d�V���#�!��'�dȹAt�-�T���sSҸ/��,-��8<�c�`��j.;�rTGf�Qq��v�C�ɗ�i���ES��T�7XO�l����ק<-��4��8�|�T�}o���7�!�D-�w9���1o�ދigY8�B�j�⣃f�}E��pm������+2���Z���j��A�J��k�<�sPk$-ߢ�!�9�73�j<��L��W]XlxVHYEB     400     140w}�S��g�T�\:�^4��57�f��={��B��5�b���P��;!e�2�,!�yO�g(��NZ�1
B�-)B�%��xTN�+[��5�K�q�0`�0;H��K��A���w�j��}�on)����5�v��Wi�//����LK��4^��6��ژ,=A�W�S��?kY�A�q�-O"�IP���2Z:��U�ɐ�>�Y�0�J�S5RR���;���p�ߞ^�[���ܑ�
��:�T��>>�*�H��s��e��H$�ϗ�ZL}R���i�Weq���e�:��1���=� ���e�{�ѱ���XlxVHYEB     400     160���9`�#h����Ǫ����l!|���><�UPt�;���d�%'8V���~y��R���1��t�ӈ�ma��9�v*�J��6���K�ʲy�8�R��\а5�]toE/�#Xi�̈́����6���U^-)����b��	(��|a���~j`�nVtAO��	�Iv�i|�Q�JS�\9�L�a;��P����K�Kxo�+�z���h�L�P����B��7�sR��d��|�fc0��3x���	���֘!%�{�ހ�ATH�r�n�Q^�ePs.�1����|k�����)G�e����b-���+�j~�!�W�uD^ �%�dp����5�SDU��XlxVHYEB     400     100q�_��ʭp�	�� ��,Sڞ����yNM~4�@�:��X���RX�o ��#A�P��D��▪e��������5�q�N��A�0��=�~��d�p��9��"�{Nm=5���]�//+��d�����
0)j���q��d�1�Jr϶��&Y�7�����J>L�'z�V��/uȦ^d)4&ٍz��L:�L�D8N_kh[��j7q �k�ĩ�8<��h_�7NX�����K���-L��D`�XlxVHYEB     400     150�*`b� �7���SG|��T񃌦���r�c���썐;�"^�1~�I���t�;J}I�|k8�~�M�mp-�z
eΨ��/�˼���rc�6z����afw$.��*3�igE��[��{�M �*��rF�ѡ�d_E����������
�yI��#{Gܸ�K?����̉)ď�"�-cM��j�J���Vd�t�'���5�"��[+\F��/	�|��]�I��;��j[��xĀ�2x"Fvg��V~�A_��L�������b�k:с��uf^���ܘ���L7]$U��)�PG�H����C4C��g	?���DK��XlxVHYEB     400     120���u��o���\%BX����zʈS'R�jU�>�CiӜ�~�,��f;��G��} `#`Yꗋ/U �@Nc��s6�����A�nS���:��cJ~���"�(49����S3l?��XxO��Nze���RaH����������h^��J.8�0���<�*��o��x���tMۺ9����bx	*|_�2x�넕�g�V�*��h�\׺�i��@ǏQ^�ML��� �UڢgaK'�z�jT%]��H�bXٗ�������u��ۡ,�|�Z���πў�kXlxVHYEB     400     130��y�8س�$�O���[�(�6�?
�F9���Ĝ+J�Qn.A���_>o�&��P�$�;�-Y��@��i��a��r�@��EP#��;|?]��	�p�$C{oI{��Uj u�/'&M����ڳǙ��P\$��[���$� l�0DQ*z�z�O�	#��1��Zn�+] IŠ"����Ƿ�|���k��`٬n{�T��H]b^��Iw4AF�t�2�R9�uhO�q"�_&���7`��m��90
%<8�����ɪ���O� V��'�����S�BF=����Br��a�,5�����XlxVHYEB     400     1205�a��)"����e�a�r��c�UetC�08))�V�ǎ�J;X����k�PЏ�\+���j����H�ۦ8q��/U�lB���\<c��2f�$�R�7��
�(x�ǜ����f�2f\��Iĩ��@M.�9^��]N�j��&��"��.������Z_�eW�V����D�uNߥ(�I����q�ǉ���"p�%� 0�u���k�1��ϳz�Pڦ~z ��RA���@aWѓ=�tomͻ������e�ͫ5@�@��zfTf���EF� �Y(�XlxVHYEB     400     140j����(T\����W��xm)�pW��2Sش��n�Ҟ��d�E9W��u�j�f�s�[�!���/>_�
e��pa7ι���7M%t��W�$ +1dl���6m�E8׆B>h�ZӤд�լ��ֈ;R1�j7C��b)��TEz��b���=PU�������>�T$��7!/�������%	:=EXܟ��B|r��nR޼�����mG[l��P&(�ߪ`�J���=2,Z`���N|HiV/��~�x�KT�+pH�.Q
h�?;�/>2��hO��D�/�D;�'L�7Uo���IU�L.���N���XlxVHYEB     400     140Zsl�{��F|�A$}== $�48�2��pjm_����TfL�/�g5��]`���Y!�[��zZ����*߻��x�WH�;Ӊ��T�]�WZ�~1\u2-E�����'����L6?粛�-Q*\�b?ff������[���@��pl�ف̾1->M��rv�	W�<����;�|�w���e��zf�߰�;����y]��VZ�l�����ғ��I�[��Q.lC�4��=O�l.v<A�r�	%r������	+��U���$\7x0
P����'V,��lZʏ�M2W]�:_$��^�Q���?�B��{2XlxVHYEB     400     1200�g������n/`��), Ε7�z��&������v�{h��f�XDC|$�$�:�<l��I���"4�h�ʗ5�;�.�N:�k[�}�[�8s�@6B�;��̥b�()�I�b�i���������ခ�H�"�9g���w㬇����De���r�����9Qr�]���*�(�����q�6O���pry\h�\��O+��Ig��[���A�wMw��c�c��&�x&�3��ϫ���`<��9�L՟j��u��ą:ݏ��3�y��q�+�T:�dہOAR@N�n�XlxVHYEB     400     140�a�"��~�����Ex�le���ձ��������f����le�6D����w��v��X�Y*7]��F�[d��ϧ;���Nq]���iT=��p[-���T���b0�]ң��p|���OS������6�O�o��2���`�,
5�ՠ�r5���>�i�K�qF7�[.��U}��8@O~����g�:k���W:A����~퀌�ceDUI]�����I�Ѯ��rй�{�z.�&[�h�V�G�������p-� k}��V5����a@�5%�Wy�G���.O8I�ņWU硣��r��Rp�,��l�J�u]	��XlxVHYEB     400     130j��9�8��E�yI��`&0�k������t�fX�W�Ѐ��+Ǹ_J׭+��DQ3���:�0��G�e���g8e��_�bf���j��SG9}��N�_��z�r��_������(A�h(��<�8Kd�:OZ�mh�K�tz���,$���/r��;�N�c��_�o�J��v��Q6JS���^���<�ێ���i�G/��	=<�kd6d�fwX��{7��\)�%N�|k!�?���.�� ���S��0��6A��b�1g��WA��7C��C��C����$~�(%��XlxVHYEB     400     160x�)�'�2/�S9�=}
��6�A:����ɮ�����G)@��|T`ē��VQv`@��{"_�ur~0cz��m-��)�מ�ak2V{�"��)����^Sgy��Ѻ��`��U��"�If��b2�[g[ki2��HC�4)z���(t����#���lRH���I��e��'@�uSY|nYG؆��Sں��i�>Կ����t���p��=�H4�C]^����_��m�G�ݦ���`sQ`���>0&:)ŀ�z�ʝ�E�����٫���m۪�0��eh�[�'<�eb���,��]%�`|M4\�Ǡhe��4���xa� 6J*��ź`qt����^^3M#B�XlxVHYEB     400      e0`ǗVM�TЋ����_�k;P(�<9i����x��|U�CRq/�=��5�d�e}WT~�!,	w�>����6�%忆v)Բz?���@d�i{�]�����������w�X�6^F�n��ND�%��"h���流�s�fAQN���)�mT��
 h��N����I��^�J��������rGR}t%ܛ��W5n�,a$rn϶�Kv�×Gz`�f��&_=�XlxVHYEB     400     150�bj��;L&3V�)��	�1}۝H9O�;;�lX'�w4${܆O]�G�	j�x�6�PBl�(��|�]zM.	P)���0L�Z��NC*as^`�6���'G<�|�⣹Y��2r���u�p}~ñ�3��V4���@ M��FwIY6��^p&��s�����e3���oF]�E��4خ(=�~=��˕.Z��v+�kA�g�n��=��O�>
�]���8 K��;*{����_l��.��8O�v��[lJ0��"�є�tFDE���88����7�ݒJTTH�-~`hӰ1ވ	��8�!��w��Vd�Fd�ȿG9km.��XlxVHYEB     400     160���4ʱy����F���
�?p)��@?�N �&y��e��61����*2�I�$��@�y�!c�{��v!LC��ËW�Զ�IX2��m��v�u�=�N�k�`t�w�$Aѡ䲡*��>�)*����2��߮���ƌ�ɱ���bY�-��(��@��I�]���1�;}e>R�@�1�׌)�M-�%��T��Χ?Z�q�^
>�K�HM>��4qW�s��R(FL�E]�Ѯ� 7S��Q!��?6��WK��c��yox;�.�bě�� ���
�ŤQ!�O��>�m�U����>�n��*됷��C���)|�@��ċ܇+i��8�U�_����W;m���D�XlxVHYEB     400     1200�g������n/`��'VS���7"`�Q�Y[f֩-1�t�9�3kJV�{m	\��쇇�!�n݊S����2!��G�kjf����J�?�^k� ?+N��Tرׯ�)����g�����CU÷O��W���y	"8x�M&LxTB�q����nǅ�Iٚy����U��|����l���`/j���x4n��e��u��w��K�q#Wrz�^67.o)6&�,�(��?�7Z�/�\~�V����s��<����?&Ny��0�������j���b�8XlxVHYEB     400     130���!�,Rg��R������WѲ`;?Ш>!��U�/�S�7���)Ɲ������tN߈�4&��n��Y�E+=:�)�?��Ñ<�EHf�DKv@Os�VX�� \�`h$�{� ������([��R�m��
(ٹ��.����I�M&r_R@����n��S[FvMW���x�����J�	�N���8i�A�����Sl���zI�X*�e|m�'��E��1�iFN��l]�eej�D���M�P�7U��Pr���X'�$�h↿�X�*���3]�LR�q��3��<��C�P�)`��Mp�XlxVHYEB     400     140.un��C/gtT6H
�A܌������ �T*e����R��M,*(�#�!,s���(�]l�	O��c�H�$��x�W�� �{(��KF�t�e��R�'v-1 ���L��M��B=c�1�nG�E�B�ơdf��F&Py��D�,����-�o�ʍ^�t�}�\@R
O�cn�G��s�ڮ�+C���a,�<�-2YT��J�L�84n�Br���J^9q-_[S�Qd�9��c���͆����05�rc֜kU0q�I���)�xT^YS˓:���
<��4\3i�Mc
YV+T�m\��c竔�8wXlxVHYEB     400     160鉮y�4��6^��C|յc��ײd~��<-��=>�Z�]��&jm�*��[b�D���1 �>2��V��l�P�|�&�.!�B�	-���g�rca���؂�n�'�R͏��>
"
�H�䔮�h�b5%��\(��lk��J$C�9��y���_+�#��O���Zu
i�.��])��)�)n��A�Y}׌�Ha*8%�5	�6�#��8=�Cg$�b���j{�*��sљG^o��8?�j��\v#Y/��%��U���d���ӂЏ�
�cI��h	��G8/�,[пٸL�b:�gyD.h�&�۔����nu^D���Q�O@��P���#�����X�~f͆����Y�XlxVHYEB     400      e0t�1Ja>��X=I��ÐmX$C�a䖟D��+�E�»@�<yD'-�.4u\���נ��p�C��a�ޚ�
a�;aI����e�!@S�!_`��:�w�H�1�͊7��4��5��X<5�\x���1��gJ��N�l�֏=��f3[jo�Dx�$�Z�$�]��!�=�5�ﴂ��(���,R�a�v&SQ��n�_\�����a�L�����7XlxVHYEB     400     170��{�����c!)qg5��V���.��5�_�!�y�=MH�}��z=�*;J�X��P�,�
[>;j��<��K\�~<�aC��ߔ;v�BN�ͳ��aG�`��l^��Q́agG����iE��I34�BZ���=�<�����a��~2$�>i������gqm*o�ѻ^7�$+�l<�j���[�ك0��u�M;��v�H��� Q��{�v��5$e�\m�Ħ�B�2ٚ��7(���e�c������RO�9��5ڧ]��FH�.ؠ}��{����QH��n��á��K�f-{�P��Y���rz/N�����@�T�3*A�>�R�����[4�A�nba�]u%5a$ë'C׫�v|�o��XlxVHYEB     400     150M�iJk�l�[?��d��0�R����=�9V��k����N���%����T)b��%��U��; Ս��0��,�켫u�Sf��J�8��eˀT6)W��J_�K���L����!�ʃ���;�ʰi�
�sL��(�����k���9����ޱ���#�xQ`��ܬ���jfWA�M���HuU��`�%�C�}b�?z�B���X�#5���Ui"��;8sR��g��;����[{bն太W�8D�dW���޳�(��O�7�C D��.����e�c�,_�����O�0Q8� ~C\�᝼�(EV�Z*{�	�ګV�YZ��XlxVHYEB     400     130ϒw���1�d��L������m�H��0i�E�Z����E{�!�k��.��Z|+����������?b֍�i���]H�W�o��Y�ǟR��	baw��0��"[��V�[�����pg�,���L_��h���UL�#�',I0��h���y<�@{PHu�Q��y�͟,W�Y��wu��ы�5���˼Nd/��L�v��&���R�2�ӽ9�*)ɢ���PBԩ�er�7�hI	@E�__U��14ٙ6��Mʵs�VUKu���s�E��+d��F�]�VB ��u}Ḙ���ص�XlxVHYEB     400     130�w���QT~���Ch��Ղ6�qf�)�a�`C��E�+}�{WJ�����S��3K���f.����[�p��4�D�jc#�83��?���%���$�#|�����ʪMD��h�S��!ܰ,"���m�ʹ��?���j�9��K+���xǜ�����E7�^��e�'�Ƴ�kܞn;W�ԇXӫ�Y�!%w^�*TjoM��%����p#TzK��5EF:Ho��8��E���
R&�8F��,_�V�[���ҎT	;(�ߋ9��77.V��1�����o����:F�[XlxVHYEB     1b3      e0�e�3�KֶRr�0=�G�����.Bv �oXs8�1��eB��yN��P���MiF��6�&TV^}H*:ě�o�&��9���"T�����i�ˌ��������<��a� �e��M^�m��"z~��!qML� ߟ��Fr���'w"��C�_���^�O;��"�>�E���A�B��+��O���0ɀ�`��w�?a{ k��j��