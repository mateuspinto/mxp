`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10640)
`protect data_block
Fi6eyBEp3Gv5yPdE3jl37xZV5Oe0LjmMbOfsABek1wpSzzwt84f23+2gWQ/WDCRRwd4/x3zHtT2R
ibgGPfSSHeexCK5HrQrXhTICsLtjk1yeWiQlWCsgHx1sdlFNU4WQ69rJd36xC01rx33ikzbxiLVI
XXPMNOQC+8wjGiYfcVX8okyFk+Vz/oTvLq5m1rZnaT2j7fqyh+NL5nUKDu9iej8TLSuLUKPpD+mu
pyoGGY/4J23cw8ht0Zik8aVztg1tDfy+MZRS/Ro7ZmpEWmzW+PXVZhOf9MpIkJIusw9XWKtEAl9s
zOM2JBkyyWgcY6LIIl7ZJ29w/a40Ct9wbXoHPGaYV9dB0+VOfnkn4Yr8cKaT9xEH6VzENIxssxoy
jrUjwULWPz0vEWr0UlmlkuO5mrH7I7LZgM3TfV/R+tlEzZ1oxpLReLUT7K9S5PRcPIH8S0gImep2
awWPGSAUFghhOqlGlAnD7iynX8hLRaOuKNL1yYvUKUkkfVkX79AiFVA2yDGixGOZBksslepkitfX
5/Uv+F3LA3SJaWrGfsiYFSifSisPGiyHwIcA1ZIeamQIXNg7wCe88iz3apVBGH4A+2918I/ojoDm
AntJlB1lemhKbrAZhLyNdWL0DxSGFDuCGOBKS3R10TDIVlnyQpA2vf4yPxmUoQsMb2UqE4rWXU2Y
afdMJiEhjVIhhDZkfAm5Ip6MKyx1/zlDckJ8Hjo3X7Vc3PVooIOZomNCNTi6IyW0IzusLOqX9daq
MnpBnJ12FxufCLrK3Dd00rSzfP09B7gzgzfqo4FfleIOfdgNrEKaND2BDHZVm1hz6tM8rc+244Y5
dCXWHivh6uktweZvy6NJral0Py9JOIu1ypbWO5BsAAsuMw8tKmzbhVH4k+kS+nj2GMyGjalZB8x5
xWPoN9AwNaRD8Rb0vE/e+A+A2n34F0NdCFRYu4qpy/1vK7KGTEO7ziuiXdAi/dEA3rdK7Ug/0c/H
16j4YAGV2jv7Ay7nSt9K5FzPHTxABaaFOLJWwDaeb07wslEcBecrjA83zCYkdarjibimB55H6n/v
fXiJAC/vPJVCbBx1MTp8KBgeVQEM3WBKIUKpieLmVha5rXuZ/56wT9nA+t5a6HtG9EjBf8qVsoJ9
4sMNCwcrZ/viL27/B6g3hsOLAsd0Yf8UmAH5iGv0c835z14kVhkbXbsWk7ib20nHSSL5gayzNjGI
TG2eTYdjc+K62Omo42N4XySP/XwIWGeBcbOLCFMb/MPow2MrnRvwgOJyHGGr9/oPa/5czQiuD9lH
TH4UuKvV4LylR4dbxTyVok7QYg6h4NmTrVe7If55ZEJnIDuwpGBVbpozeff7KarR7cbFZign2kaG
9KoQMjeqyz6i/FdHOIYTlHy06U7bAtEOYaNEIrTWiC6x8sa5ytGlbpexC2YWby/p8ChUGOQ6luwA
MGr4EFl8Lx2IlApyiO764L1Q6luhkcN5by5bmXv5SG+r6Vc01wVNNOuUfectI9EuCfcXUZDDDVw4
u9hDsDmgnuO7CUhyA/clFskz2d0YmcFqwYcakIvxLEBnRbrDKcUOiNiG6MDP3KMPIt3LNPkHhN2a
nHPDfTBmbTBXFbd1nIirgmliFm0ZT+8KMhpk6YOLGKNd0tfh/1crHCpBx45yhntbb6F8AJzCJd4a
ZRLURiGc1nAsR8CvVrfRbAizJxHbIBUA0D9YA6iadh3O79Ym90OVHFBztFyc9QV9IYXGs0nAoNQK
4DXDW2MqQllNmDx3jwWv8QcXf/etSIN5gIgbPaMu8RmBWeivnp7jfS+gndbBDGv0Tbtv6sKKWQ5T
OYCAg8JVZldaslQWqNsIgNdb6RPjckIq1L4fYMGNGmN9r63YqH8xtC34dR1I0+7FTf/7RIYJ4PKq
X1YTdIx2Op224yw62/ofXdvfdkNCdJwg9YH/SY71seElr9D4mXFzgkv+6cY04blOmZxkU9mMcQ2x
CkLXKxOUPno190VlxiEOoimGlj8y8RI4EyexCRasvptB5hdspUfZNkWoA7D1DbwwpmSntycCkFQy
rPha6kcdWHyLkjVfEwny80oPXH0y+2CJCUhGdz0+joaliOdNIJ6vaVEXCkr+UvvQtx6aMJ5HYJt5
8MSYr+nlzta9RSeua5YizdUKIZ+r8IY8HZ6Wd1fYzLoRG1BQzss289au6Gy6AmqIBPl/jdhyzbEp
XNyzp7jBWGRx+8qTlXbCrnUI1+KK2gNuCFHXNgRxsSARtXcOoXSu9iOKiWB44tPvOv9AyzUeLXb6
wIrC66jnvGYkVi3A/Kf1r7WHqkNtpbUGdFY7uFdjMIJ5kL9lRE1jZl7MuY6eORCL6dgm0mjlcwGR
yIFED2Z201FK2VsVxHA0wSn39nlUr4QWsUb1V65mAJeQhHpxrfbWxQbYLjVb138hUfmMQid2mH8z
GGjxQxekW2jYXa908NYFAGvJ9Dz18bNRTZJACMF42tFAE0pSG+AoTxPdS8dTHxA4YgSBPLBIXND3
9pYP7PnwCPLNN2NYdVxsB6yBY9n4Hc9a6BzpMMI/KdYBv6ml/iBsO7x+skyiKh5bFCMh+1kni3tT
QO7CrpuKtzO84MNhTyDMJT8z0RHv2cBCQreOg6m/tWXVG4pwt3EyRbpG75G5gfZNO/YMZ0eukmZH
vXlB6ZsG04Pd/16Prs7dtJWHMgPRE3otzCoEfdK/NMr066Fke3k8zibl3UgbYPgrvbHYN7a344bI
DgKNos3L/ACbussKN0XNZhyDmM8aulRb5jjbMyYdpKT0XbQhZbNGsIOxrpnpYud5Ih9laKqfLbjE
dvhr/fjH9pTpSUN7z0lO6F3s+f18JINb44lMhupm3KlZb7WlLFUZdGcXyQOFP6ATjRLo4CC4OeVR
lmPqB+of9m5BZx49kg/HRxcWeDhC8WUMNe9mN9i9Yw6vhmS/TOFVHVQpBF0bIXe7W/LYDdfVNRHF
KxYXFX5bZ9Mwa2jHeKJ+2oq6ma/cF3H5yJvvjEz1DFE+geW1VDexNTzDvSDoaAWnUpa02MldxkTg
hrOB4DC202RzWl2hgxNZactE6yCl5CJ0bQ0qv0k5i/BBfZiGMdHtbsdOCwe4ZsLckr5fnmamzIFX
BI/BqvbqkmyGZqsTfI6Y1K4XTE6CYmjsToAUAbJUMuPqHKX3mzoTV8BiaglMBTtZ8rNmnEp1CXo9
jbg8qiPaXCK4xzmI8sekDL2n1jIhg5UiST6J8a4xyO/ObKTxMSTVUW4yuW7XWXZDYP3llj52bOmz
4sbaPQ/t0tzM1NbjILjeYfcPdlh4uFznQvLBWjxEy5SdQnWUXW6nZsy1km95QldTu1+F6ij4iefg
bLoUmwoh/DjA0qGUNb9+m1ymHETnuyBOreNMXcHvuWcRuj2VX+KgSqE0GsheWli82ZQCzJY1zir2
dr+v/UtqMplpNucwXo3Kpr1jkjtWTVSynsRHi1f+ZLW+icgX+G6rZoEmktcAN8gjgy5eTP8m6Fwe
jrncgPjTPVnazYQXfPfSLtmmRnkHGmltlAIR6tOD/w5Rcd0Hgo0R3Ld9nHMIFiMPKjH07YRU7rG+
f5yHU2pc8D+2Fv9LET2pfdJRLAAE1AeUG5kH8qFLjsh15kCElBh8fh6MP9PDM14Kl1e4Ttx40XuJ
kMVRjEAQxW41q83hXqMlRVD93AE59736zVcVb0z2gK0+BCiQQ+2CKfLPePGrbPr015SYg3iMzHju
VquUgkSteAPTRSTx7S7QA3wg9lUAPAN43ooDuEwcYIZ0nAG0FygV5Z0VmgB/+BoYYUcCcsptb5TA
q3RdcgtaWEPcldYmZdMYl97pP9LPar01m7NyxzVcSSVznfecGV5ghULv3QBe2od2u0CsbW2GPw3S
utbIxW+sEyCEgbchF9b4n5RtizKNdgW2ZNa1qbfYXnGJqFeLyVoZLoMjDetKTo60AB8DZ18JyJAi
hfvSd+raXazMGSutFi1omajdQgrOJv+2RYWFwh6Xuv4z9Qq3Z7g6qMRYSo9ZkH+Ut7o9n3jdYBCZ
k8SuskeI/OnNp1Ut5AEprMvMoFipZkeWFZXKAH43B68iUpQLcndSTZ6XpIDKu8xHf/CLVSZQ5eQn
MtcCc3U4exWxfbps4oyRoFy6GaQ5DnILBr/QkkAyI2WjHiyR4xNGIBAaOyEuOhkCb+0rRdbnP1tv
nHxoszNQYKi41nPvg0UNjphJUdkQWVyUQxrjFNZNU/9OoRbXpVdimkIzoTTgNF931hJlcJiRznQB
dgyTHg6ICRUHgur7z++Nl8xAM/tBSqG12o/xPqcXsi3kN+KZIvC5HiVjIurNJuNQgqZ1cnsR9AEm
85Ez8JAlQ6vFJG0ubjesluyl+QFkXvU2FRRIp+c2qoVQgE1vOiagZqNkoQKA5/3i4e/tyMw/CNWN
d5AbZlzOvZOow2p6N8Rifd+QQgFdN3JZvJ7cDo8Vdzvv5zx5iEpM/55NiotlGv/eN/lQC8PK9GDX
95MqpQoHCxdVqarvEkyc5TWYtuPSE9TFHYJf1pbe0CZuf7KtPoundm/A34y+NNSe96MOMUTCGXJy
44DNSdb/gsQpY6XBjGEWd1w5RFUEO3vy0REjuna51nR2FZxIuYZ5YUQfv3wqTN1Mfzyq0DevJKRo
Q6XmHajWVu3wO9vq6J0e66DcLRJ9a6z8bQNZg6NmfBBRjEeQEiolnr6qhQ2jcMNJfG5V9mtVUwfR
94hdojHi0CYIeA7LPBZjle8tYFuHQZgVh6ZisLCvHTdu4EEHyk6dcHNxPpOkzOAJJ4J1Za80lZsL
jAwA3ko20mTZz4weE38XcSL8IvvZhrm0KXycBc7hkIZjGvHZEDr8p/pLBRhJLEz06Fu26J148Szf
iHeAIZgAJCrtA22ySZtfPs+wHjkUKpYnmCbOIebKH+uiQoI1adja6G9rIDZomtIKxo8P3kUibgla
kpuOuVSzw12LZXixdxUTDwbJxEN0y8IWy0bxzTRDIW0hkBVMp4YnQp/93RhdGJQCvIXO6hWP5exh
WUqrIOTlpDFaGCPEdllQzIK01rPmhBWJGI8cnfouyEmnxHMK1Yae4QQaYZN1JojlNisx4aWH/UGS
sjVOeRj+mxq3+/EbQEPs6bpv9vo/vUhzZa0LVtcdX76dljlepikbKoXLnsjVIWKSyPezpOD3D8/Z
RkO+XyvjW+FYoG1qI7S9t3xwkh5AgNrBPsejsCdtJH2dud9VffMGTy0AN3YhRohcy2ffC1GuhQSg
ISVNTphWp7YUXQu98RFISvmezqfS4ghB6FXzpYhl8hhTK39UDtWM7m0gV3izH7DdvbJyCHf3H9ir
71z9lJyKVML7/EnZA+hrfiX9f3thCVxjxaUlZNhjhKHcJjpBwtImohqfNFDHzk8/PanpObcYrLMK
Hnw4HOPz2Mu19jfdHAmuL5j2OhHMU9rMVEVQ8DN6gypV0U+F2UuBInOBL21WllBeK60e+0k0h019
dLnIEwReXiXEn8jDQCx3nrhLtN4cOpcPwuz2Sf73GXWJYAHZgb9CqZwkTeH1KYSr6gwF+d823w6G
evPukvF0TFEUWwaJseBI1f3mWncvkHjiCFGKBjflS0alhfEDAkavdkpZeify+LlshMOlH9CYyMey
cteofeMz5+y4XfWDnqhISfp13srjTQIN/+G6BlC7hwDxGm0JaD3E1zQ+kRhxcSu5FR4GHLA70g/+
1EcNihyPSV1+ct3ksFZvRnJOeojjgaiPuxIvfrbpQzRBTVoJR39qtQXCJdfwfzqWIq/3E/xW4gzn
c9EvqfirnGLtl4robDOaE/cteqKcsBNPEPxCk4tcZtKRF6IMpIh3oXz3V9ybj9M8gwz7qMVlqP14
b1yUh2F+QkpfbyQMzq4UW0fg/q8VruLY3NX4jjc20ascyX3mILKhNN6WEb+CiLXDpVJ771RnUlCF
Y2psRV17szBvuJ6TYuewRk2VXWuiXF6sx2z/OxJi3eEpPW85TCNT+EHSuvMFPBVKNyo0ppUYWER4
QA5V6BljK5prdtu0ZvwDTYDKQW7zIndDW7UZZ1JOOL5RTlsCPefXiRcdDL8nSprXSDB/sEXzO7hb
60A4zIb4v6y4lWGM7gHGCUD4q38vVSYgWFMSnYofNmJCw6XOF0O0gSpISQs6nEAKxI11sSGVGgby
muGMqbe3BkBA+dM1pWg5zYwbGpZpK/1MtQ7MWg+KsOqHBAPoKdcLuzqi3qt0RyHME0PTzaqOXSVP
bVgn1hZQZECEGSbW+uQKAcLr6rBUwKECN6Hr47xjjrc249ulAqkCvp9JvjfwatDEHnKdbjmLI64X
YwBBmlFZ3yieGA4KScq3UeFeA2gomzFUEz464nmXPm8BwaCtZkFd0RM2xJeL40RpJyqbhaxAdfi2
0ePQ6rUYJ4mM9eC/5vTdoA5Dau4rf4alR6KXOyL9KKRn/0Tvoh8cFbBTAJQatDTQtFOv3pm25ult
jj3rvJap3lwP+nJ4zs08wpqMFSNrLCCsRrJnGRg8xrgwxE57dzdYurdD7VUvb/9ElMZGv0hyNb00
nbqHhSycysKiTrOgXgzBoPx08kWJGDwyhGtWDYXieH15I1DGsY3BIEmf+PX6uR54elv5KX33x6X5
hriRlW6cu/4R89j7ealNZWUy8U6Q/qBnHYM87egiiQ4PxMOjSSAYX2x8shEWU8LcSU7i7ztRImlW
CplDomW62ij8bzfCTihp7q/n1C77Ooj6UWCoZJ3HpYBivW9GSWiSxNE7NvqFKQutC/u9pEBVe00j
yqV7TJ9MvppK6ech30ZgOUR9BmbeiTAc1V3ly4ET1WyEeYE2WRdBaj1YDAE/+tPigGKwWlNQJG+3
13/aGPNNo7freyIIpd5pTv/KSP91fvXLk3LhiPlL+/mNv6Ww05QVS0y8peb7Z1M/7M8Q/xqovfns
RGOuXEWT/wd8tE4gzXMz5JQ7Bs94wVJECq7jq/aqdECzVMURAsDCVZ0GslJgwU81+sT5qauic68V
5gowZm2E0gqh03thcEVCtXRELLnhhLQTXcXkU9Ymck7clapaQm7rhTYM5uvZ5u72Pan3Zl5qUO+Y
4WwAzrU6cItaQ2lLP8viDBH7B2YsXMwQOtWp52IBQtF7E7tqUiur0biGg8ncinsf2EanSW/SQnS5
4i3fn0H5Updw4VSdPcF39/1fK5aSb+hkcBmkNiKprje6YNZWuv73bcFGSUpwhnPaJNfsqKQW4NJf
vn7oJ+DTyzF0zR8U58zZVl1F93ij1Wo6IDzbFH5dzJ53KbWVwR0GeP38OTh4gtX6HWHBNPVAPLgL
r5Ew8avhFSHWRuUe47ao7phr+3nNlrI4PRimwnosJenScDNsqhZzWwLPL0SJwWdVdh/obrLg+YJ5
umAHjXzueXlwcAfNGTVHorpd9zAsUC6neeSWx/WyFHoHFCU5yTj8uAPSYZvkc36cxU9vDjtUzZ+5
oRuL7OkLtYKNfRDkzdsKNSMyn+TsUBZqpWpdNDiSWXwhRlTdMpcNdkfowsLt2VawcWFngslX9pKv
lCaqVQjOo9luERjkScbjVlHs4HKNfd9Vkb4diRbksUP3dX0J1s9ou34fAt9Pq8RszTdgN/pm7F58
2ASCCKWHHCWvb5LSwKxqxsZwk5GBQYH0c7aOK0Kff6XAbOMzQf5+mYaJUM0aqM2DGyDVBdWY/7IR
FElca7n38LX7o08FWfZE4SMcd/vMXEz1CsN0PncSHg20NIS/OqnWeWpTLKfEBtISYw6gyQ04Ek8A
bIG/ICeSteTIn/UgStg8+exWV2V/4g/hxV24RgEz3KbGd7AU3mdYEUtjoWEWU9f23WtUX8vRawyI
tliQ0cyb5fG2zru1aJT+Pk8mvnQFnU2osvxX0zqYEgvtzV74izLaZdj1+u2T5Tdt4p+eiIYwma9h
F4ytniTr4lYtpJesEAecAyQffWZsJr5JsFflZzC2k12c2sG8Aq6NFZaFus0SGjLfCA9eyObgw6cn
PkkvLNHtzzZPbZAqFpFJXF/crC119BGWSUhANDncffF6mswNdDxhjKJYfIOD1Ta5QPksnPbQEV8a
Ac6wtQaPjJi1k63xzSwakMdMmgKMgcbwND5McdbUuMu2cFq1+zLyIxxihX/fKbQNkiBgKivxCgHq
Lq728qceHHZAZLEXsXVXrmlkLon/bjnYIUk7Xq04KjNvTjvEAyaFU3Pt4fjEJFxxujhMnup7lqxz
Cqw/WiVMorInzS+hA2YTv2K5BIiG2kHd6KkXa/MCBXvTNjbEF5gjuAy+N6sQmWfL8hw+y6oRPqqg
t2zTapfUUfInWimfE9FkXtTwJMLkzc/w8WEbW++CAN7SET6i8g/+gGgSbnE5kWGMw5ytqdXTnRLl
Rf8ftKe0j9uHgcLctmzUHxOqSqjdOFb22tqP6928rWb6n9EVV7Th6l831/FLlhadKIrqJpAE6AOD
5BeCRIz5XiIPll1Fbc5n5XZpgePwE08CAhOuy4xlATFe4xVe3x8jeWq6AltffcOr+Y8AC5bjFMxc
HVifwFYDmCxgBazxGeyEjNAIJntPXyRVSusdxl/LAjJBV+ZVO+rB0z99hXNJg4TjrGhD4q9DYRw8
QuKWP+ruFRT6QgO0oCK4nO40u/Qvp0NilfWOhEu9Dpof53sQU4gVvZj8gtoZhVPDg+kcequpeROw
PZeffGeqi6xwmMjmRcxKgwqo2qCyr71X3TasEuOymEWV94r7SFHqhAx+7djFZtRXoOu3EE3GYTEP
Pp7rr9hr18bIjGJ3YNqaAOrc5ASBZ1vpC6yBoTgSR5JWnCl/JdQODrxr9V51KWhqz/gQVTwxj9Y7
sIMf/bkfKJ+ntYWm1ko9agQIovJV9Wn+5pijwOytZvpPyLBx4aXg2uHgAMfLggyPtiMmhH40KDzF
IMNN7Wmq11w3sVN4BgDxT/63U8Y07x/xJpsMnQkuLIowsMdFjSoxvC003oPlyYnPkTBywGh4EEwf
SNDiOWBz43wXsBZ6jS/Klxp3g0sMlkLDTjAPk13gVC4GgLDZjGzKQU1WaW6wh69P/t7zol6MGlh4
AuIvIIpiOfqPn1cnmpYhe8TbLPU28C5cBMnY64/0gBci0fob8dCdsCrecH9PU36t5XC48miXK3Ff
YTcx7kpRdWZVbIu9qW6OnCysDr2SBzabvszRqbVrnzC88zXnGkMZPPw7ilON2pmM+eNsySr1TQ60
UYYC/AdT+Hd1L/KEjC1zLWWWK2XDWbLOjI1ngfD83eSNMh0wr+P8BEz8E7lKMJycTNGty77D/x8w
L5ez72jX46sbPk9oQHRujcbgEb1r+35H6YFdPzXAZafkIo8oy7OpMGuQtgFkWgCeYfwmg8Cadvgy
IckdjbOioOvAwOhE1tSrR6trSsQ2ekyLkYVbzE1UP37JrDPtG3SVHFVOtdvhcf5wBBTBzTBrlxvu
nqPCyvB4CTjESzqCTqUwUgB3vhsPnpEIGJ5y9iQ3wmwHb7DrPQ5q/hpt7pA4w45GOohK86dwTUoQ
YBMKaT8QE83dcsNVuiloQGvxwioZV5J+ten557epDR/24llqVq7I3Z64IWsecPDUYTFC1Lzt5Pqt
bqaTRgHkPDr9lt1xleRa8Z5vyt158KJi53yepuZ0dhzcXVbbiiao6wqE6jj7LiP4K1Q3ff1iAzDe
WqVA+gvmhiW+T0LGDxs4aiHaXmnNaTTO7jzDEwSipzybS4N9o25eEzPoGXfB8nGJEu9vWDWfEhbw
1VLbGkLk/MYEut4H9BAjpdrw97pVO+I+pW9qTJ9MvMnxS5Km0TWN99fOrEOLASrsuDlv0IxpwOMl
9I/sdm7JDfTgDNhokPASM11hNdHYPcglEwsgkry/sRwaspB/FC+90PZ2OU8adB+rntd0aioJysqn
S6jp8tc32th+0A3I+EGYUSrrHPxPAThC++y3sMgQ2axswtGmkl10zsEdDOF9YMPJ31HgSSpl4BJf
AKbOW7IsFo1BKDoFMCv9gCU2k8+AVk02LfuU3cP1umDZpzjeVuD3Re+wVEw7VA8n5ewLrcK46UCL
dGNR08rC8RiBF0Xd+NQ4AxkPpasS7MYMPgCCMJvSlKSJLo+zZn+fvXMPFMdUTqBr7Oorf81XtXzP
JPKpuLKPX2+SsGJpmBJlHeZqwFp5TVj5sEjsSqF1ziXR6yyg/xoCRIkc3Imtz4aJgSgOORExDG8x
5JmgD3LoFCxLZU1LXNMZrah7kAvMQRpgkWlWDxU4Iodyl9wA8pzgYbtyXH5rEk8tsN2EkFcsVrcr
UtBx9zjRz3uLAPYRcT5vLxJIBj9qP1f44CSadVqGyQPeW7W8VnRLcn/ONRMX3KDx21esI1a4iIMv
CbxbJBsKgoPVVo97f7OhJZKhRAWns8whm8NWaa+9q2fVeyUzwwMg8UwHnYfrpWtSLFzehi7Nk37E
A4WfRRnLzVbhnhvCYM1tiBROJu8zXOV+IxBub/yQYpgK003PQ2k0TJYsJkyo0lxiQIzzh3u7TU8C
Ek0CSOYhpASayRj8E0O5Bq51E7Udb/epunpU2mdxeE+iQA/2Kyzm8WnVneiQEDKm2o7fE45wZC5c
YwRotQYgNlcce5kwcKMgtY9cIwWEaGtO+CMncrpd9z5PsHQDUMV7d7S+eD2sEa918LvqedbJasrZ
zebd+9IXGfdCv4dRRKlnX8r0xiVGo/t0T7OgZoX8NqtT+o04wTfDGpDBn8PNa3PbY+S0yKdSfkxA
qnpGe1zR8s/y/k72Z9gnJQ/ndIOcFHqkyyzo6RFJUNr7Kw8ixYY+GqGGRhrYpBA/kXY1lUG6Dk64
42kxuCUdxNquiIEcFzXBPFc/wkU69D/Ylg/rk9F3+qgu3mp9oIUfze/JjUzU/RkDM5Oc3yzpHcuF
bNRULchV/fCo0EnpDx038YvyVP2bEmqSnXPmKqaSZRVhjIZh8MP2A38nXvRI7sHP6GtiQcK7bocr
UXTYf5driHfRg5CLF8uPnm6+FQexzfBet/DS3IMnt4WNHYxQj0RBaJOirgLUkmb1yQ1/73fkzXDR
esAoOtPA8GlQsin91kIaEFbhb125/dBzqV21QtWTJXNzk62ahQOnArUQIM2iOvigpsIZFx/duRbD
XhYoWzg3dLbm1KN1TB70RcCWU+XvJq2mtPgRDIcPsu7HSiHTYgduaExFBoFlmEG2+OEp6E00i6Dp
M+Nri1r/z7Q5+7LO/JtJIWH+/6ZaWYpOz6dIksXuSRm4y15BD44nA5kB1zqWPd/9MJFAdrMCcTZv
D+LZgtFmH0rbx214f29BB8bdqsvPQKKg4j2AhidkcxiyPXb4W9d3QVVoo5jFwOnYt0KogEBQ42I4
cGT31j/DKEjDFZTcAGX/dGEABuGIcT6mPHFcrCkc1pn1ueCSJ998s0aZkI/L9eFfgLQQ6Y0yWaPe
a5XQIS3Z9LnzILXD8kNqUzpx7d6w+qQkhqLa8poX1Nwbpcr5FmDuQM5ESmP5fOr+zOxlqHeu+z4j
bYYBh/g9oRcOBDaTdXdpXnRzVz6XqAVMXn1Wm/x0u8cTQpF0FNsuC4rVgToKwSufn+1Wl7g+liuN
aPI70ymOsdMIagxv/gnJdCQPbKFoekgcsbkN9hMqIVyA4KFPKJwhDLRF3nArRPRZLSPJzDBJA8R5
NbaEYU4nq1Vl8YLXELgXv84lD9qNPYeJK/x7xYH8oIymqkXYpuabyoj7eYbqaakdb8ycyQ5WTmBq
BN/63ejjUkR6I1B6apyE/ToCP2mmAXaYHr6/7lEnbzSU9UE+nG3TT47SC9uFZkclVbNq00WflCay
qy5CGG6zUNvfFvN30LgQ5wkM6LdTidmxOXJusKxGK0TkyfuoN4UJghqjVNXBUH25mMV8CsutjkRl
I3enafJ33PXf7mBXUw1qkZjHDAGtPgdbGYCW0Dkq+lbgvrdgrgHVvT47Jq2OA6ia8+HnZGmBjc2l
0K41f69GSDvEkqP6Ex614yA5BMaRAO6APa1q9k+Aclg/tahzKEQHpgVTjjmQ3WSHsBXAVUUpUKXW
yvRd9iEdGEovXcMLLDv2+w0ytTrqGsVplq1lazfkHMfDPMuOCfs2n90MzItHQCgUpuiAxVHONG6s
E96JER7NZdrkaeHHG09ooRL47iqGq26VswfiiPDlqptSVVeo7TD2TiuytpnP+x4ibjnLw5gJLKtm
HdVuP2u2wcnIAg0IIB5UOrDe66nv1TSLJSgGS4abUWGNUYJDJsL+JqZD39vNK/3G1SCdum8kYAa9
3OWkgC6JEDyqeWwt43DJEsLE8mHNLP5fVVqmeKsPyXAyMBJLLlJh+XniH/mF8nIq+qFX/6sr8FQw
oXhxxs0JdFkjoeX2vmTl7lWAqPtJt4XaKjYTn5yyf9pxZgbOMzZ6Gmrh2CLxy3ctzlEJILF5H7UE
vIj3llv8ntSCeIG2vGq4u5GWGmHNg4iga4QUG21d+ZFuFIfOO745km4DPwxjt3eq11qhlhYZlpo+
7OPwqu8j4bRNCg2wGC4u8hIA/kJK/WTdyptnaYEWFmtIYCbenuBeZWFoYWhi2PXsZ1G2d3P9fjxs
7Xa+QwDx2kaZTFnG23/BzLlosxIR3hltPCeKxZJCajJ3SVMpVNNjGsvzdInOK+6b5zGg3slBnQdg
kCRKgZS3sytZ3QzugVwf2A0Whjduz8Nh90+QiHgff8/uXeGCjR1fYXVICwT4Zh7apuwx4IFj7dGG
/NfUC0NUjp2Iul8+fChvv+7mt2eT861YQlw/B4VxFIsEcH2CqJVcEGLwN/3xQ7Qxmr66IGIzu0fn
25CNkEM4FTBLwXUH10oWixEm2pAPHgnI/hIBMjN/si8S4kDSqKF+qAB0JdO9PSJU/zCxii3XHLFg
d+PyU+DfTx6fnkMFLrc2sqlUEfICrsw7T+DxCWeGmSRz8EgJdqDhwewpnUTK8uPKwvwXTGLRneat
qEYLG2+pM22Hlc0NR8I1fPalbhi67I4LcUnpMOjZggJzZY5dMFzXWibZeO7//j6GMPFHtBK2Qt6o
peKw5ZgjzuWQV+wv3hGgmwzLkOBT2MRi7Z0KWLgm/pdo8D7k2cB7A8HrAMUpb6QI2Wyaab/4oEP/
qWFL2pRgjvVrrBF68uPtX1/V4Iuk30vS87O+un9MfsXSznfNLdNYq82+RhR4DyKmWV6UJsVPTAAZ
AvP1z6xcF6op7eZxfHJrw3mWUYBmDwfyn589pNUG8I+XNK0b5CTJcP4hrpmeGEKT0+jYfLSWyqil
cizzoxAfPJLL2kpXix9gLoy3MkCjcWqgA0FxyXU/T9TdRJJzRxTSJSn62v5khBKq7lfwqXHi0LnQ
atEWub8ScxgCUp6cdnIkTtTWyBKSBNKSyOhbDjNm0KnvrygKE7UbHjgHfovjhnfSzLx+dO1rNzmI
v50P/15xYqEnIyUF1+jSrc5z2PySGeJU/jUbV3HoY8LJ0WjqrLogTwngm+q4jEESAFkAvVNadNHg
g4J+Pgb/+e+g782DHCe/IwE6MGlfXgQZ935NZwomgBEieg9jkvYEZPgTgoPU3ZInai6fyjnmezB1
FwbS6+OC1329/90mzHjMVNjY9zQsMhvMsg2MzaK2BBCzCJW/zMY4r8jBK7KSN/cy0p5COGkBcoqG
b+Iwso11ydzjDnwz45+nZEd4LZ3r2GiPgO2PftiBdBbW7mSMKeaqLJS5YdL8AmZuUTxtD3Rw3Erj
/UHV2fdwGAxX1/U21ow4/xLmosAo7sAuNOVY5bw8L3GBUlA/hO1Nx3MQDaFbKBFkGMJcfyOBGB7x
ZLSOBnNleGPX7O/k/Sz44K1zXzRMO7VqxQd9CYnWIPxrLS3qadOmDckK+kgccVSPFjZuRY+0gpjO
hRzEra2pGbBTuxuq6+JGyO5rnTjMCLLDiV7Q+lh6v8p9FiIOrlSu0jldeuSRv8TPfSrs9Ni6HeB1
HdeZe2ve/cyAMlPTjLmP8f+LdR0x6Tl3tp4iLNTVmSClrXSc2JNwjxA+7qcCuu3dIlPIAIaiWbkr
H63hVdYVDGhY/wk9x+YegiIMFRM8dzkPEg95UWepjhStVNw5ZswaZr8PgMuFR0j1SfYrm7JZ4Jql
ogrlCtmJ/jVRIcH9zS7UO+BXxcz/sZ8BKtIB42UGVFqvSE2+b57VF2pgu0QrEP2rVv3IgxZxGoH6
6pT3DLCSgFYy/sEYk84tXX+gB5OvPZNBH66zyq8cGSFXcYluTpQ=
`protect end_protected
