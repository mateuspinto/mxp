`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8400)
`protect data_block
8RkC0djadlXTXSB4ZKZENWQ/pgYjHF4UgpvHfflRm9l2YOPihrztJYapSz1vtS3DJeI7X+65nydH
KYRJj3zQoum8zvo75IKFsPfFGDduzIfJHwlduGEx4IAD+lkeaRCYnXVCuhcxRrArTDUs0veGq9vN
7D+DDXJJ0JFw+ADdP97feLEt5fibgqsXjs5zHb9kKUAwZFXtHI91T6SsaeGWfSf3yCFH5+OKDB0y
GopD8MJCZv0BAaFNeJGhPnMLKbaWv+GX2gqdhADXfj/BEcMOoD8sFFNquZgVrwin4fbdjMpP7PMC
MuR6ecmHC1+eZytcLmKSRtO8XVL+IADdmQ4Y0KXiYRvb6IoIpFdZOE2XtYdYTrWXWHnDsk7Dou0O
t8ESQUETp56w0+425qgXQmbx4/kRVNtwhI9Egtt3znU/SD5W5yg3RwYBkFZMXDssMikl/i3oH5hH
MaLkSykwW0NqllVPNMqqPotENvSJPvhNuWJopXFNIFNEktX6yGlNj0u0WSvG2inaER3QHkO8mKzn
nJ3eBWXNvkCN2TJQFTeeK+D+F8xcHQCNg8SkgZoMT7qlEn4WLQzh9U5290ycIkhxpJl7zuqKLl8y
tCk1HwC2L91ZUcOWJdz/FCI1yc5L5MHvD0MO6789JsYXNQxhkS/w5KiY7c606XTu86wUmZcdTElh
1UgSu3X1KpZoXwjv45Gw/DYcDBG92m9A6KRZ8OpcQdJr+hwtRSOopaBOFHPe+FGCwxP7rLkh7PAY
bq5j9xbwzOvGOwq+0flupc3WDcyMQyFAnBxgLxnj7Bat0ENje00KYmoi/jBeQXGJ0ylQSKXewlb+
wAd4dYJhfOEatrx53y64D6l1QEPAokREFLjQ+TnWLB1/059CtHyTQlT/wu7N69wZX48EO/tCNw2g
TZmtPaPmU6JMBz/TTZLl1d1AUH+N//WSaxtJ1bDXBO/Y+mkkZR7ifKdLFPttM/Y21Eup0vIUNHsJ
Fo9UJWtUo0SLSgPhN18ZVTLfc6cn9xVOy/p9BPwwt3vMdKInXjNJP/AncmAeGT64SNk/ggXpO83Z
mlP80BG3I825fQaiAI5jrRjoxnhs6Yrx7E4B+sSqDodGkjAEUFepjrGN+Rdu6HikWY6j+Sj4cfj3
Ul2bLbYGVWsf18ErfiVvX0mh2xmqs/TrmepYPPw72XSUWOGeymdeeRhlCwemod45BPpnxORCBASk
Nk4u+yJUtyzKldKQO7Jd4kLKadi9GBKtiNYpi7trxyV94AXPiVSDD515VcQx1+g21hauOipmuFST
P3BwcRQUgvtY8IWVDsfgr9ipriLtJ13+fLai7Pg5CRrvFmYTQ64ppoo8B1CC08ECh++n7PWP/+l3
Ulw5Lf+5p/SrtSADQAzZyt83bD5iC0gV10qNCop5lpHa1vCVEsf6m5lOGWsPnb5Wh+qB7LKFoLHz
viL7M/+H3HhKBw1DTfthv+BpU2YNivVC41a+XlYUJvZBD0paYN+l52RaVtO0YmQzkRrsh0l3f8ob
HPYmv40KEMSsSE2xua/ZrxsUzChkkGD7xBFcY9S7nlKRVU+qSMWItvGN9q/Y6DPDxp2VkYeGQ3Mp
mQp19TDmWjB4F36Q+xNjU17vIrShEtv7U6w27T56moizzbC7Ln4OXAOIVs9qPqgvRr7eaArC0C1C
gcvJtmJsQ2a5pZMsS5RRqNKalMcMK44tQDeROp8D7Exu/A0twsleBryyNGIcx64R5W6xtKr2Hfms
4sifCeCO0pjwQ8AsmGQHjMBwruMbNPYt5DdBNuwFa9jfn6wsyIKEK3xlsnDxK1qfSBMvjiL9U3rD
8/vn5ebdWXMHETN7Lo0rgDqpMk9NigXtLKMUF8UxHjyOBlOZTlA7xgsVHMGYQfLhMraISZT9ABix
s8+D81VHilxd/u2e1e5wRxCsgefWTMJRNrc09sr4alhyFkdQcTSrOWhKwd4kRhWYMlvbkclMhu5d
lF0jtPgfHDHHcVLw1v1DCTemBAKKIu6jjdC9KzuUT2xWazrw3kmqJeEP87GyjBsVAhkZSa3nKwR5
kDjzUHl9I3YQlSImWB9y/2jXKW87e2CFcUm3fsw9qz8ammj8Ws/bH7+9R8DWOl4ArWCJ1BVZQSEX
uubj5daWia+FrpLc1zWK0+Y79IBlZAZpf8C4MigxijhsTU6Qb3XLid68KOd+TD1udl4dy3N0RSGI
HAMRTDyJZs/GqrNKYZTJ+ILine55IgAX6e07dWBkaEYulfRPmXvvTvm8UJT1pVMtK/CCQexjoA/6
gMfvGRSwjibCZ96lEDE2o2+60cbHNkyN7dfXNwfiCcRangTM72NH34aUHPMculLYeYcz9ITQioyK
qShDkopKl33pdlJIhMfeX81xSEOTdwhKxcPM+gsGOc5BTyk2BgqLkHsQVZgu2A9QkATNbvQruBUs
5KuicvnReuVNcSU1FQ11eYZ2noBkLXDqXjjaR1KylvGvSV2L532HDxH3jh7mEeEsMzcD2TCRFdOQ
NUR6K4YKd3telN9FubI5cTBRYo+jAZF5epRBStBqRnoxZcOtFtL05UWXFQ/kKDxwwVXEsHlaytzw
Rjd8YZ7r+5AwKL93EihFXnoqN7fNKQLmRSRKSzKjXIQerYcE+wc2jdFnc2uF6Uu2l9uzdw5D2mBa
ZE68CGnxeA9xEI66h9GvRmz5jJCphbE5LvmstjreyBUVaW6fbRKeyKKGBnoSEL2LJNJf8c3QvI9Q
0BmPdRG3mk6cBqsBsISbxShqSM+l2aOp5uX8H57BcqkGfS26oEWoYX9996Xk8m+wjSfzFuuSzKLY
BVkOHnpoksE13JoZjVukk4/YA1yNlVLsWj/37By5rv92qjlVhLhsQb49LM2r2KFxkdoDWBmkJixx
kpfEQUIti3DB5I9el2OiRZ8pG9X0RlI7OQx+rRohwOCkdybhGPBLsFvcJ77Gp5O4zdCcfx7EtV5U
xxAUtfc4zTRYakQxgDva3PP4peYxHQmrYkXzzyEgxRyAiVfYM3GBk7/4GGd4b4nZuCTgYrCLNaaK
5Cvt6l97jXaCF261bHCTAUR7SbpU8mYwADf/ea5w8LzbC4Pcmj5YzLE+yQxLQxQLVsOb8MVq4iUl
pf+zXF6UzmHHiAKax62YfSRNwKv6r4CKzfKu4r0Ib8IqykpE5dnOt9nEL42yD0Hflaqi0juUaV46
+ANZi8heLJqvefQX6e8Wz8l78VPyV2uK0Kvh10TenRII3sfEqn7rAV/WiuiJbFM24PjyfOZwyW3i
/g5tFwW+5Gyz2doXA/2CXRYyMbDirv2mYCn+tKHOSg8N5XUTutmwh2V3sSUqY0NOTvjIclUSMxjX
May7fEP4gsj2KSc9IfEec8lVtHeRXo6WDX9MTTqhc3XKr7mf+mry8jchLTVwjZGnc6Ff2W7lizVi
xJ9q5R55xnnFP5JW8pkgUYqB8yG0sdw5mUIFVhv0H/CQRpMVozAvaF0sRv+A2+6NU1vWEiT/3pz5
H3EtG0UIPlkHlRjcH6mHQ0W6W5xoPJtwd+hiVsJI8jRE1s5viWxODyvaqwZPuDzBEVZbD0xjmhrd
LRX+LORVfYSKyLnc4T81BBgDTMHjTjM+tI49zg9PLMzdCCtr8HZwx/BfOpkaz0V6v4VdtCpoiEGK
CZYWLfr8eDFyVA+BIVAb8nWXvArnxBhXT99anCyJ1bw3GgGsCTr2tN+8rrw+sRf2LcrX5Mwua+TY
E80+rdPDdsKnXK1BzAqpC120kd6NBrE/SWuf2LPQGZVHS9N+vSl2JrbGY7cHv96mveoRZEZFUnr3
l7MB5VVunXvi44Ke/XI7e2GDu1sL9AJF6d5Gq8j3lOMoqsotvnORWc0bX3pfHy/jdp2gxdTfUuIX
5v7y73P/CIfrO1V7xaN2jXzn5xLYI8OE37kBxvuuRwrgo5j23Ly208e7otk6mkauyPaSgGVg7cyX
2WPUDNNoZGlPLcM86a5tkRGrogZVF7CSsj/phJkebveRPRSgWEr2Fybuq8Djjm7GLCxgVMlbi6kR
uMV1xMeXZVtm1FRGUg4wQNGb09EvAxcCshTnSvwITL8XXTEe9WBLfm2jxhhm/GexiHR48zWZIcJd
8vZaXVU2w/ozpO2Ot+A1IQXy3WLkV0vYoQAexKCD8toZasBnBG2iRjYf0vzZKuFeCsxCSyMQuNkU
05Z8ieQSc2uMV11YarqKJjVt39+dLdqJ521x83GTZQhPR3p22hdEnr7KVYPsaIyKytjXWxTMlWdf
hd4SSoVFl0Sv1x2T64kJMJMY8X9Le6N2ChkNexv+Q8Nnt1DB73dHYyjn6aIcDcBSP8/2QzeZ5Yx1
r1IBEcwLEE4tBczIqCPixSgsV6SA0OSKH4VFgn1ABq6hKYqGaUAaOaCUCMeluPMrCDR9twGrHusZ
VPjyxdEY4W18CTFmQAgN3jP5YfAJ57fukOoMr5ZfQnBTBsKxhq7tiS5ygkIcKv7Lq8ytlfhf2OEk
YmcnR7QN1sTphVerRr6G8vBJTmjE9HsYtFYVzrLH5QRvnmiHbEHUmE2nuRNwHmzoQ4K5qjPCLq9w
uAmSGBXNnDKazeH2IjRb2JC6k8yiKH4PN3f9hKbJn5ZQHfX7kdKWQQqL39XpifCpuj5jhE05IRAz
Az5S3ilK8kyfmoaF/oVyFKz19gisoYuY68jgvFvEquhGi2pcmqwSrvBNi4BuKdYoFOCLPXKpeot5
pzM9LPfJzo1Nh3YlBIbKzRHga7w9KWY3cnK+KbNbjpx57CxfaYmHPni768xpbZN0EUTujor4+Xm4
QmvAaHEXxNC/c+Xe/cTyvqrcNw09Ggz3parKCOXYMPIc87FwSHLujyT6CytZXu2DnQbNUS5tTdXz
xASOBhTZ7Ruv+VWfy/fcWoxpSsQDV+z5hb4OnijQQ+3vDyTkU1fn8xxMdN1p1eUgPfLB2txeiR+r
gJbv1ne5fDEK2jsKUTibMn4EA/CHIcplYAGOB9CZYqNhXZMges8fRXiyY4yZnwo3Tu7EMrlq+Ome
qiOqquhwL1fQbVdSvGn+imj/nYrN+hs8vHJZDKyOQDH1nJz46jOF/nOD7YIuKZuqnp0jKOfOjnys
cOJY3BY2yBHXUYNizO61uBMFl9UI4T0doBBmz1Vc5AQlGYG4xsjXrndUup2EEyAZR7GRm2aHpCHP
7CL8sLtbuqNxaeQdRA2RwzqQU0w3L9PU5U0D0ftmNKkFgr1TtxpIyYGnJyq3VSXA9vTNiJWNpG2Q
yxdIfdhBElfp4OhNUFxJ48OmViq+XZuFX0W2JN46iBLb9svZt1pPY6i37YIaa+O55YLD6hBS0JWh
g4sYQYYWU0E6NgV6npXNhzwxRC+6Xf1ZK5qWF7JnPW8BKtQctlAvozWuwlUBg3uSbHlF3hOFAjTU
6k6YrENetE+Ow4ONl9ExnXJhrORgpdpYPANCPMXY0RT3ONfZxLUmTzaHGZcEaI2B4Ubpe3lfnfCx
aHsgkr4p3uaiBi+hD01wCdUbCYe80Ti28rK1FxVOlGAiwP5Kq8GgxbPPFRbI1GmaG5KGTzTzXSE0
RJZtt0vtvOAgF2PgKq3VFgETr6BiWbD3cGcTHI317Q9qu78mPmVTcZsgLqyj4dePkRNncUaINF9N
VsVmAKwoGF7bOwSzlTBDDD6sbUB9K8l6qYGB89w+ze0OI/Ov6fHUTVLa3FVQX1aFjAYCFB63b9Wn
ebKBx3NwtHS/QFrfb/q2H71rnlwJR47dXgeMza4Eq7EwOsky7mpvuN4Y+7EZjKLQDdWCk6sRuk8/
5CkNYYG7BMI/JGydCM+L5MPBINItzeKpb5ODgQFRv0y160+v2V0Ilcc4bd2laNrpHq6y60e7TuCa
BEZUYbhN7atZsBWhdn+S2FlN4pwxWJpLg/AUvYF/GV5CWEomJBAYMoz+ZQvxF1+PL3M058Ce6rt2
Dba+ux2XA7DbSZUuAOb0Ryqh0MrfCQDxXr+Ex1qSdR9usVYH+WvivyGhbAQWBhANMv0ANZy0TvrQ
PIb+E0STSJnBBcp0pWRXBanY72M1aC8Id60oVU1rHtGXwf9+rk9mwa7jLZjDQ1MQ5UY/fWinxASN
LZm8wCNWhTo48S7d+a1Rodi3zn/koQMww9++ei9kMi+M+6+UUa+EmiyXwKdP4XRGCpnuCDTNoM4G
Y1aqda2DM/cZmGMUKzdtom8KAyrwoyKefBt1qU+ztAjPQYEQB0EGf773RO6GzB1AHLMUtFKbnUD+
C87O9I1IAPsrRXFeZjLxEN1PYMlE5pRiNvQvDUSShIYgW9oBoaXfUT6RLb5+vxG4EPY9/lryDZuO
b7EB+6z2Jq0XEjHNZNo9ZuAXT3jvtRSPF1MBHrjsy7ReucXuhEC4x+L2h4cY3ds4xJeczfW/Pt//
JECjUWLJ2iEoSwOIsk4+ofCtynxKOB5N0rzdd8aRd2v12AbxVK4dzQm+LJBKrCPp+h4g5DWhvv8u
/IP4nY7zlJ/1YPtHpI7FyBF/hIfYBEbTG9csGt1T2AO+KhaKozb4+d6huerGR690aaF5bm0V5rlk
S7j34CvrgPsH3D/7gpr0u0eTLiNHr+W7xjvLNG/s31DeboBZ4LQ/3mAaHKJn7xZy1SRtEM0QoupX
5ks56HUVH1uxHYpixiaZNXHh5f1fso9TYyfZ0A0VZTZiVMIeqdOUBqLrTBmasFHNXPYWNe9/dBAC
y7q4F8UArcAZzce5rnrH2Zussr91Ian9cJl+munqJB3YVJOs2GcwLzOHQ8SqtSLY8tPs8n2QyzPW
9cJbTJ7mbjoS2dzM84Sd3fFxauiNzc/20pgh4wjaA+f8/potR6/ueaKYDMvCoT/CJWLgZz+O6qCQ
bnyUy1T7GwHTTpBqCDrPXdTP1RQwUdAaXkpNMW+NdBmnwrguYXSzb3yV0TgbFu87u7u9VC/A9CYf
DXpZPJ2kVrSSoaxR/qUHOfk3BnZLwnvzAuY/pp01QykkS65Lw/6gWFCMYiwFyeIpYvokLvGal7ct
U5Ku6CtGWpnnbHw9pNEfc/IadmmOVJErqCv7nybLyYI3ggAc2zoGwsdD7gxyOUuDhp6l1r3cC/FR
vbSwloH7l2TA4ORBmDshkposc+b0TEbfY03Mq2wuWMN9PghgA7XfAVj8VJ5tDO2NiyrYo5bE/2rq
jyTfVNDiMLFbL7aMrVoxZk1QqRB/w7d+5mQHP9rHxVEIJpJ7kY+DNWzh630MW1UH8nAQMrjfxfDb
YIsjMYPhqNKPGb397ZKUa9C00OVV5rMOs/BXmvNHOGhmo7WyNrnHrZXh+qvuvDqZnY7PGsA9SEJl
INpSjbEDYbUSBO16zzenzYofuvOXUy/i5zDGcgvaQ4X6fjjEBTmwW7Da+eKOxRzpZH3ZYuqnbmp3
GVcuJM2bp7H7JTwES/nfvVBlfBRfZ+YDPrgJgZkixtjmWueWpusQE4UZ8so162xZV6ysmZAXy+6/
frmyyzslXzwRsvH+qIh6AObDp3D6I219Mp0XW/imXyAk0u7ave/xjLgOy87FNMBUj3DHO/r1DQbk
yngH0ywh1AquXgZr1JXb2Ca5gSoMljRuPd1YRbTfiHb+mCj5ZsQ09wQ98hItEU0lJrf6ZB0YkIpg
HTFveWRH1s1KQBTHB60BKfuYb4rL30dsViJGQCJEGTQxMm0UYbJ/z3n7ai2Ee6PpOHelg5GvDpZM
Mm1w0TWQRXiVQenXl0qydxYr2vHYU4QmT/YR3CeFMP6O1KF9RYC5kzNDBI6+nddwGlxRSdeZ6JDB
wDoU7xklwFYSgjK2hZQ6cIaTdpe4apWWm1NIntnb0ky6WikOtEZGCgnfV9B+4B0pdOUCzjYkpB/m
qFCB9SrN3mI2DjrnOvFPppr4ONxvTsI1baVrwj5tnZvFCE1eT53tnfJV8RKXlZRBL75fqwUVE5Tb
7kgKNMdMWW6Qq4lfOS0hVfynJYjvyw9wQjlWQ8q4IA7Pui/opstQAyLhA4zQOCzDqvAQcA92smSD
BRl2FK3/yiCiNJsV88dQX1wsv3hoX9lW4xHyzxZKfTFbgItQmPQTklrfPF3K9oJFzXsVcIdwxwdp
wK7POVHb2JIGOK65rXZAXjf7tN+ulUH38HBERU7Z+vOh6C1g62rCShV8c1vZSKfJNZMl1nHUfqic
KLPT5RsfwoNQoUGW2pa7WA30YncvBly5YFMTpYBViOU7EWJAjV7exKMPQjPy6seZ77OyKpRCY/mV
J4/XdMdc073y6gcjhmNzWfBRxWS1o/qLIue81SbEaw5DzJSqaUuU33i0tnqx1LuI1Zq+iQAd0Ioa
mkngCR57Ws0CdhEZIuANZrq5Cv3L89MRkPU7MX26aG6kWowDcxR2md+te2QfRdr1X9eJrli2K6/x
J9mlVDwxqAK09NnOwrFkMX893EQdDeyKhy1wyjO+NKMiUDRu7PS0BUV5Btpv6cH+r5S20VqsF5Vx
IJ+aPA/XdzD088bGu9J17tgYJ48zC8iroUE8PEns8y7MiH+uHQrmYmW8QOqe/hn7Z/TR63RXVHTn
9rLNr1X36BQxj11bp+foUpvgERBI0ckKi8EYKaK1O4sQhdIzuK5HJwuZvSYF5hZ4hIHS0ZgXSlMf
ItuNe1OkhMJQ6u7j9HzHsrCUPjthij4TlOKTVtGX4ku6BYJCzZVk3v597f9WdH0vmAz2QE6dHlI7
Pn7tSoXEZEnC3bdzoogBcrdtfdbafHW/hQxyIRfa8xYW6ZOgQ8EfXndwNfei1UiD+rufDYzk+Z/0
LZ3EVWgVu5d9BxQwBSe7F7s+2vwUZt1FRGTb5i9i1678uJmCVX4irNDcfNkyvi5N4wAEazOugSZm
hM+nYMJJ7IzoSZUbpjSAlYan1Nbb9UK+zQVDlUKip5v7vdQFCom/ahXv/9SXiGJAEbDZyp+KN4++
gRZuFq0mJIJlnjncbw2XUW2ngCaQXE6Zuz8qkrWBvoNAIkyTNF8ev4Wq2shjXyps25eOWyO//Vc2
Xl2KVYUlCN/Jaan8gUZVAKJ/9xRnxThVCyWg+naxl0TBdhYc2aOfJTm/qfYjaXIrDYmexjx5mzoQ
T+uO+pxNL8cL7RyTJhEG2LloKo6WTcVRyN0yFjaXMGTGWoSxJBH27mYG6CHay3Ekph/1K+rm8/+2
qoY8Qwo4+d7cd9LkWTUlS/tCuA4WraRwyNTXYvzwc2kJNrm5zsFoh6dLX/LCvE+HxzBqYQD21Fn9
PR6KAS7dPxBsErsgQt0jijXC8qEv91pTMkmaPDtU4k3UJyKtRQh4HObTjKkekuo2jnpGLxPUdAYZ
RfurVil+gwfS7QHGZPOjSafg+uDlgRWadAZmSZdtkEs4FJguALvgmN7Hx9GIf9H10i5mAouE/3JS
vkxD+VafI1l2avFbMw0Rwp3fk16rqUjPW8Vxvz53qaLh53cM6/O2hxeHMXtR4Gt7azxf3yBjkp5C
k47Cbyy57q3mhnnJ3Ac0wBrQxlL/NlUfG4TQitswUt+rb5UzFReGJXYK7VEyymscem918qZsnaOV
xtxgkxGLyj2YAUjE8Wk6GxkuacrMJ2pyE3V1JnT5bKu7c/aAbm39FzQywKhAid/QLAaGZ6lC2suG
IjctnCwtuFoF7viVx9cWrGE/ks+l0W3i++Vf9bQNhRhbjK4mbF7etHC9Lx5aJbxZKACJuPj1vbWE
ZKalaDcOArGtdzMqygBbVC5p9cfFbGXbRYyUiXpIRDpRtV+ONCGebagrCyJmWaMc52HNW2bMoqVy
79edlOygIsk6ehbcCXxHpUFeVf4C6ZTILI+WXbVtWies24yywRW/Kx5zuKNcJPoGNfkxrdPhUVEK
QQf6mm+rJHDfdrJSA3L6dMDuLFf+IMU3udB3OSIz4qN/xsP6xChCuU4bTk3O8asJOAjOIr9GNdLX
cwORIVEXC+DaP3wkezSckiqYed9LyufuITrFuah+d+IVn532blYPAh3R2iaphqQhoYFJGt9NPdWR
Ayhio7/JO9X4UJ8rjpdueFAwnu1P7x3jn2TIJg/evI3F6IJVJ37jap91QawY8YsrC2+3rnru0cxU
Npt73UFt1O4WyztPKTrBssB+c4AEZT88AphXLR/dDt6rWbOhAcLkt7GOULehV3/x63bOQmUDgeV5
f7bAXENRPMdDEkKJHmg9eRZMQdE7HhxphCHTx0vAtZ6Gn540RrMoXjQhc5QSUUBSXuu0cLbAAXyG
8wS+bZULv3POCvG2j4muzA2bOZqb49VER+INlKq/oIXAgI40VmP4Fm9KnKJI7rTIe0O7RgCiVcS4
Bp67XMhBSZ0cMhfqjv64tupo/SaSM4i0w3KdBbU/TShMgng0LJSQRN33KwRMG77ZLHzbRhjS6A7v
xlAr28pxOmbrdAsfqNN/bswQ4MXhaQBWYs0CnOh4+QUR/m6mVbQJ77FJ7vN8jE38b+SJgPW0MBgI
8mgTILBE+Z/+oYIXMyiyd4BFOb8ilX6gCC7RvMciur/s/Ms773exuD7RPwTGzOqsOXiEbYD0dY6x
XeArbgX89fchSTJZ/B2QPd2ldqK8U0iTKxGxEZH3DJGebLE6LoRTE3/OfsqEkUbBk5Y/S3vhVi8i
wwYzYIluSeA63bm9GcaM76y9bz3IXHHJ0fIf5SbcgYwPmbbTzHcSx73n/8uuufpzXAwHA4DZUVz2
Q62HUSTb8kdgNRbpqOl5jfBhKfE6Cgv6ZAKdcL6f9cnjaDs775OKMJkUJFEAKJijs7SiEJpgSFW0
iO09Vn134q9ibq3al7WhOGydxNKATr4Lgz2ycQzDdMFB4HD4Cw2jRmkRitXtzuT4SC7rcYRRvjqy
nEmmkut/SKXuaya2RQjJyXfVD0QyMtntG2tX437nNjaxJ6nUiT8TXEpwOgiJ2v4ihFLoFydyzTSl
SqscHEdwssc4FycXHgxmW0uwS6TMaY/X56A9K9BGjf7tjVwrIP3YXWO/7FHTmsAd3X6GdTZ5PPzP
v7LNGKl92UJxI2ldqAWL6EmdeTX6Wn9WiMKQpxVw+2AHkJtfMN9aJnHgnMs4T9T6LSqFFdMH+fUQ
QvjJFflAD/VhrAH7LVV7t7eEKRIbWXKbA3+PrQpMfqu+Ft0xZ+5qIhM0R7gMt6K68mSkg/xpHifu
8qxPYXF3j8mkv0+9ul+uPMLhpcBxojXlPbmzzxwuLU1oENf/5CyDsoFYx8xhs3e5SIuvUJkWiC8z
HA4Pf9h+yPVcyBLDmVgMIElzTxZL
`protect end_protected
