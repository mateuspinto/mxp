`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3168)
`protect data_block
OxDTa5Nc9pUI++tRvmRndeemX+mAEWp07cSLio89/THQ6mgCJC3gBU3p2mRrRhc0/k1uvibIVuCM
8B5YmOUOu2PpP79pmw0jepZ1UNE099+LzJOEWArfWdSqrcj7ZvgDWqaPMrUQvObeNrJM6JVXhjsU
+37b/rFtlMs1wCgKlVtx1ZzFRDE5BiiWrp9ZQ0ATTNL+lYBPlSprZcPzePV4/iTLMMVrGdXcQALd
vxnWpCJNFcA2uzYPseKXMLNKQ7qWCxk8fGd5N2GPmoWgVIfPzAnQz4+em4lUIV7FjN4sx1DdRQQ1
NhOO3Fhp4vF+56WDIfUuZpaE3WgFkvTp/Lo3Dxc2hqNpcaUyUlSncTqpSL1EIzrpeqwfT/S2xYbc
C+vJ+Mk8oYJJfjCsH4jre5g6X5XPSNBaJimXE8vdUGvOFtHAtLEJjUxbjX3cHgc82WFMrx0jqU98
qAeFMi2sRVym8DIFWJ20Ei2zCwD7IK0Xr5MiQBzEocO9jSPfw/dd9TWGkGDaxl4YsAfA7fV+BCeL
p+ozkDN7H/BDD68ivu5HFZ1xxOjwGJjQOLWCYOFyOsZS4lsyxm8KejVfFyu/cn8Q+uoz4wQd3Qd/
OVrN2I3KugFRShAhwaClxyw4fQAMhlYyOpN++Zp73UZ5jhGsvyNajjWcLe4MptvAGqKtNtD0Gh2B
NNmfv4zLSBGPnU2dd16EFQubAyCOdRkfCydNCF6AomYPq9yY0aqKug0iYLuWJKNlqLasrcc4otU4
mNjJuEmyXhYZVW/Es40swsdxZagoUO/m5nWDqZg8fjeJi5S/dVjXYeXBZpE372/5D73GBG4KMY/F
jAbq06J52e0XF3t58mgRPR3ADbntNxhVe1CXHg7VhLHJ/Jdyrr0Arob0bqzdkAisWWFg788+1CIB
6rKpNkYd9KXJMHKvEA316Egg1Q0sPWWG/b70nkewWFV2HhFGXM/vqjwR9+IJ/kQubAMTPXFdbnVC
ZFFMhNGficTr4KXYI/nFp6fjuI10ud7Bt02gufBhhn4GVaAFeQxh0RotiVwF6U/Bm077OCqv6mzX
kX9671fLdCKF7xDQlETdVIrwkCk1osr4hKQUJyxQP+fyDZ/ltOsZdJokS91oYzRplbDEmrZ3/3ln
tE0rv8GMOHwGaIroc9S4EEFiJwpop/7bJ5y/60OsiOrQ6+0vFjV9/9mLjsIl9ERdTIzAMfhNVjwr
KEtbUl1WV5HFRES5ujomJNI7zsVKrCLNDeirPorZbAC3E47PFMqrjBi4jgNv9sRMCGctC6ryZzv/
PD+fpuSBfISdcvh6WVvOlb4aOwwEtesU6G6/40+3CuxTteJMdMIuLTajZb2GSzojsMyFlZMbObRC
i7xTdVbVtudNfccLkJkku7TS2RXeDySwjrknix26WA3lQxD6OeeYfm1//3v87uMf39eiCsK2tE2g
dyCQ3aWPZhdH0LtgZBKFesVSCaUeNrsggymRfLBHHhV1JOawP0giaGmpvBe6J6uEAqIVDL1s5jnu
p8yYgtNk8SUrhn8bv/CHoK5P4eq/ngd+f8Isd4JwD6O5AwdtemzyXgZiUCyhhvvFT9BmoE/dQFtk
06xXRm0fLs0w8DpYTWPblqjF5bSZ/Lglr1iA2Gz034jEF0mDlwhfeP8jw0IhcbKG2xxrwdXlsJm+
xq80m8zTkcuLPjZsqoYlMuWr2bBlbb99RsqtBoHFkXMewiFkv6CHZx/nRg088fRWLC1W1Fxsfuet
3xXEXFNOBKb0doKHsjBHB1VLzUgOAufjisTMJoNpN5t4jleuj1i1Ey7hA9xhEQ1hreejGYFAuJXD
9cy1cPBV1lWDeglkacvdXKfDuN7/bazMvy0YWQPNMh86gxJBzTFq113uIVf84eQkChkIcn9McmMG
3ETlKgV0NSOYPG0tFNf3/vIOE6pEaLg2KhBY2rmOy3zhqidQmrpEhe67HifqtvNHxzgZSM6GN5fv
OYTzPJZa/iUt/XIt+PEMLbmRZNiU4gczWI9nw2UgsXpdpLxP1ZSXfs/R2c8xb8XK59g0USoqS3ws
Qh2WKCBtYBFKUD/zzhsEoBweZ99RwvoMelhOQEOh6lljIZmn+mjPwkYVto5+2MB34leWY2jRQexY
e9Mx8ART6Jt2xQmG/bgGi3cNBoYnXR3rXMDNo0qIm1uNkxmaH9PPqtqBRJkbOFH/dmbxMHigT5T+
ag7vl3DTb08C4232JHXWvfNvCoXHZ9dRG3J//T28yWSdUq8WieLh2L0emVPOoDe/WXuUk+Ey1X3s
4QoJdjM92WrebXLBcaOWqtIgUR2mjZkCAvyC/TuUzgxCf+NeJKNjQ/NzdsmG85vcH/bT4eVM0KqX
ZmMlMja9YcuHZ6uVWhVPjWjBR/d4Z1PbW2g88u/r6fNacyvQ8J8stM/tLk+1PPx06zDRi2AtZhbQ
jaHHoyNZ1FKRGQrLHilJCMHf5oCpQNm/orOGXoXLoRWQWK58IvHaFrUwuF3VSIAcXf7PQCK9wrsn
JNXrd1EJwui0v5Rr6tJaxbu32av5X9XfSPlzw0ko6JiRpkUGbD5C21lJNHgqhVpHiWgEmFRjhcUK
9tdOO0q0evzkLSDguFKzdX4qelT9n5dOUZ930T7pW9qvH8jPQL9C1hAe6ChxcgztfWiuCDse3llF
GgiyoGOmQ16wp6cpGJ0EkIy13NzobdOJmB9eMWkiplFqckzFpvnHlbychay+hZwU75D5pjgVOBhE
jdyDWJ13dVcnyU23crANmzaNiF0KCREU62BrV+TOSbk4xjKfhE9Mz8GRBCt6o5h+5/Ke9PqNPcRg
2VCJp+ynoMmP4GScIX3ukJCvsff0bMC51w1Wzdqrd9a+Rv33FM8g4+aMDnF5IyQTHRhIrSsuMj1o
mq8w+fHvY+1JtWSp/RuIIUlR5NoQe7MURipSiVUTIG2okaz2Bj2F5ZNHk+W0dVnBbdFCIMY+kCZZ
leUCZc6yDKcqXmOCTEUE1eIZejH6p7TCo2eOKYwFYW/i+JI9W/xd0Ee2Wj8MciDJX8E8ENN4w3g6
q02A0JcxjQwLMbAdsvT5KzeIByyVnJpmqiE/O8weBbpQzsqsuiQAWWQPYteAlHNT+U45AiILuqZR
nTZ4o/9d1pW6L20k4I6zWYoNUMlW2b7qlGWDwuOdf9RVXtNtlFUMnz6687ybQ8qNYM8dnh5ZpsIJ
Ket2oEgmBoH6J5sCErZQ1xThSvcj5yNtPfEfg4qNYByDQ0H2PMAe00394d233wjf5ykFKWhr293K
HOH7IY1QN95KmUgqwF2ouyNozDhtE5RcDs1bqu6OTj9zLZFOKuuBD4mWcVm55hrjaW6Lc/hsV18P
uRfeT157QSY9d4NJ11QyNjJPllapAJyMhg+nnVk3py9zwgeMmZVy3uofUMv4R/VTTGzN89pHlB//
YsDIMzg49663ncH8JBMJJkqAazKICC2yeoCOeYSvnAIdt5DST0a+dyf85C38JOhSq1zIm3cH1XE3
S7NLwi+dgALk8XVT/YDvRfzW3dEXKr3QZzOpQhIFopWASuu/zq5Qv92y+u+UYPd21QzfTtSLoa9s
toyLNdUDt2SHT/NwDSG8sP4Dm3PktEiLiQ1bXI/cRIdNhHDEHCCOCGHJiYrQ2iWyQ8ede3nfFJc6
sn3vlzkX20lOUWCVcflZ7SjZPi6X7/HGZI8xWOV5ad0KBSLK15nzRIww2WDmFwFpn+L+IGVuWTdE
VFaff+EhaprWKOOPSRwI1/pRswPbHQLmkhMs5y9y7VgGEO1Rvr3vmcpybPHfR/PvMmSE/iWwPbyL
WLS3TxzPSrVyRHEVxhfZFwecMHZMNp5cMsnPr8V3X8f3TNr8+wlo4EgMhfl87Yy6DgUlpt/m3I8Q
s/I/j13/9qrm+QlUNcPhULmRTXxB86/qVF1eQv/KHr+EQ+AL2W4DqLAqkUCN3ARDwCeZohFmpoJA
p7GeS7VuDf3VG8zqcCy+ElMm40NU5YRE8owRHzZly98q2Q+G9i7L5gh/XxT5Nsyj3L/5pNhmYrtp
INbEq1KCUYy9Ewmw0YOax9BQ1v8TdpTiudEGCaej8B7n2QFHOre4/MQlHpEUKu7As30iDTB8cxhA
FYJCQVzqC241lLJwA4hT2REOc5e9Sg4y430oBQ5IPt/tT4BRp8qp4rS0yuNQmChj6Gj3k/nN5FTe
AyJdfNELeOAh2JWZoj3xkK2gysiH5YDw9QD+pq6PB3Ju
`protect end_protected
