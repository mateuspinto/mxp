XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����p���I �Z�W����{+8�Ȋ"��r�cd�0&�OK�g۽�3{��;�����5],�jWO����p_���6�hT�ۻ�T�Sqz9��9�L��-���RA3O��5v4��(Q��TN�tp�2_&����š��q�L~M���i���؟>�s�5.���a١!%�]%��w+)�{�=x
λA}��<����Y��pR$S�1*ݒ���hXDi���4Y��������I@#�	Q�%0���~4|�ی��c��"=���<�4�ֽ�ĺ-rZ�ym�K5#��8�1ꝋ�� ���1�(�>g�%��S%0}�P���!�ؿ�i��2*
ꥴJ ���I�N��5�1R��T8޴��	0R��;I�5[�uK�j�q���fJ*8�&�;�1�p 呷/W���4[c��6 �7��m���,�+�4";�Ϗ����
���#�	M4�1ϋ�Cl	!/Q6������/��*��I܋�2�Ց�v�2�2N����W��Mv�d2�D�����A�Y����)�?�5T���d���`������,�~��ut��"� *tȲX�Ed�ߏ*ھ`&2��].&e������b6l���`	�@y}�S�|�2��A|���N'�P��O���n��%̣�G�x�l��3l�	���bJ�e��J�l���6��-3����MWWY��6ȅ�4�[mn�7�e[Q�i��ݯ'q���Q�p�2�#�uܥ��.z���k�lTi�ɵ��XlxVHYEB     400     1f0���c�����`1ꆤ)��Vp���ᚐ�.�7P��>ͼ�\���-��ɸY��M--^)~��뎦'�3G[\º#�!�CH���i�^�E�%2L�gm;�	���j�7��3�y��mb׽�]�'��r.s��ۇ�G�忪�1W�>���V-}O!�A���y���/��ؿ;���:i�-Iv_n��h��sػ�aS������b�ҳuֈ��1���I�=p˗�{R�"YY����*�~}"��G�߭�g�.>J0����	�f���� �/�jh��t6vr�BV��ğ]g��sӴP�k��d���//�Q=s��ʍ1�3��0@��M�Օ����΄��8��	Gq�#e(���x֚��L�;	�s�k�r�-U���VO�h�,�T'�� ^�m��Ƨ�/8�@s]�s��㻖��h�߯I�N�w��kՑ�p�49CK�#��?�ŗ�I`��q'h5A���v9�Ƈ� ���XlxVHYEB     400     130���P���(�w��E��F�~N��øԽp�\�!DA�뮜�;����ˤu�x*��'�$h����ZZn�PW�<ޛ�%�DG��y��s?3W��xDPa�����A�ĕH��񄁩`��-6�9C2�[I��[43$����V�KTF��1wz��t�������ۚ�W��=��|���zj)h�D�Q<����2x�D�#Z���m�1MOc���V��#���F�H�«7�?D��51z��̭����w6�<�����eÍ �����)���U�v*�����Z!lި)XlxVHYEB     400     120���-jA�����Z)TS`{��Ԇ��8����s�?ؠ�x��ga�X�砯��a�R��v��p�G!0�u]����M��:�n�l	)�q��fge���Rf@��#��+�g����/D�]�yE2�t��У��P'��޹:��?�5�*��̴�����0�y9�C���ʵ� ΂��K`rlU<���r�i���{�r�P�K0�)w	�&��&���v9�`Op,_U>�W�H�_��	kaۯKH
���-;�{�w�0͛
��[����>���"Q��XlxVHYEB     400     130-O�(�d�a��#μ��)�g^s��Ht�S�~i�'��gs;����p�{o���F���W�e�0QXA�o\�*�x��E%���\q�$�M=/�٤�DE�Ԫ��M\�T��`0�r1�4W�N�S�-��J�����.��P�������z��?Q�_��hL������DC�p� Cfx{���a������+B6�<��*E�T��	�d�y*K��(�ͬ�ƴ�m�����2ir7�� �(d�s��۸Z�W6�ȡ��Z�$�޴��;�(f�c��+ٱމGnWl�Q,0�fN{fLy�XlxVHYEB     400     140�����|||r����Y$���l3��&	�<,md�%�Z��wq�B��ƚ�
�E#dz@��x0�P�Y#2h���Wh�h�*�t�+YΌ���z�����ċ��QO����jh���;�^�a%�i�B
������0>χ႞�hX6>�`��=��f���̲UY}6I��_�Y�\C�x`S;$�E�ށ�8�@ILN����$�49Յ�#���ҋ�VJ/�9a	_�􀃳	��� � �j���Q'"���J Fΐ3ĵ���:��JXր�N)��TC�~aN��[�(���E���m.`�i�vvN�/����J���-��XlxVHYEB     400     180{�#�.�ry�(��4�-I��%J�:�87!@~�n�o69z��2��j�3^��T	O�#H�R"u�jr�8���\����GK�XbJw��f�Ec�m�LYTR�ۿ��jh+Z-y��P�շ���2��9�+�	��n�E�6m񫱀�(���+����74[,װ�|�#+�AtYmzIX'��ul�4p���ܱ&�6�ֻG5G�?����aդi��bߝK�uΑ$
�BF�Ҝ�<�W-�#�
n�ÁՆ(�{?�-�-�򨷨�)�3QJ�2�4V�$w�܍šgPW�^�ׅ�Q�a��`�5#x??uk��ᰉy$�s�ޙ.t�B�O�׷W؞�y�!��2 ���� PW�ɍx�iIQ�rEm���!��^XlxVHYEB     400      f0�`�t���`	�S�M�m�c��9v��&��R�Xp"+�5�|{��!r�X��m�KO�� a6��֝��`m�+������Z�T9մ�d��E]��-]s���']z?��*��u��`U^C{:d��/�O�nr-���}3�T�'��.����G����wqd�4z~ C�'����2�GBsvx�rA:5Q3Ycj��EG薬�"!����;4��|�p��[/�OnJ<�	J'�XlxVHYEB     400     150����/A#����J�
���gu���I����� H׸,�ɽ�j�O������߲&�Z}�x�AM��� ���H�`�t�3��I}��Y$���|Y%x+�f��%\Z[˴��Uw&��G��9�fCB۝춵2�$�i􂃰B�]�by��;؆6�Q�F��k[f�d�:4�olB
2;������$����K�g$�Q���,����"��=[�,�Y`�O���xN-I��R,���� ް����󧣐��UKɡ��J���	{]�Ҁ��'�{i@�K�A���3��M����!����_��3g���T���j쫗hɐ��Ʌ?��M&%]XlxVHYEB      b5      70�����l�S;^�>=ue�S�)6e6�H������=9zDd�7%}^��T�W����쬃'!l$Yٚr�:խ�w�󊉤�'�M��Q��ߏ��C�jIІ��*G:�tE���#��