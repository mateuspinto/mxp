`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
l5kWVpRKra1SrwV0beKw/APJtGBLqa3UcBFnPFgGF5wr/WM8KRKyYs8QjeSC+PaEf+pwfJL8rBZ2
yzpI2nL6RZLE2lXWl4Or8wmnGk/ai57xnAdSXCI/0E1LXwThqwSkgNebWiiBnuI2CndYOFLQpwB/
kNBE+1BxpcUpd7f1yx9QYhBzX9aKZsL6MTvl2hZ/LQC/3sdU0fVa02l4nhL6FfZZPJyWHqOU1RAt
tdN2W8qzMCfcnLXMK2SgnOsG1E6uSj7zappBcX/fyjJzjjM/U+S2abY89wB8QbNQ4D7AY7eu1tU8
wfKIa8795v+PVb07x3sC/OTfl9Is8tzCwVHJHA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="XDCWRG4CNRbSRKAPjS83z2K7x/l/CrlQjMbTAVGg0xY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2896)
`protect data_block
M0NvRdI0r5eo1YVXY4+Uqo7Cy4m/3x3x4yn5oVTA9RTjZUuIaA/vC//n7FLjWScRuv0pjoHkVrYW
hjk4ikEflkJxuUJZZuqsDfJeoU3LJye0s4TlORcaIuFAiG774LNqd6wa6GpjlCACybDgG212M6/i
28XwE+sMHJy+Mr/xZdLp/b+n7nDmPK0E4UqgVjLP87b3xynBxI0pAm8SxGwStWkR8GiM7te2IFFp
72K0btRLqMfT7rSm9iuzIvR5C7OmR/m9ddxO7NHsi3UklYSNzWUsEx5AD8pm6miuT/cu/RHWOyxn
qGk3RlGC03b+t1yg+T2iWG+kZ5RpTonu7TQ1DwSJCAhM2W2WNkg1wpjc6AmJRFc13Mg05BInEqep
MPnT9i2/OdesYbb6D5ae7CzQp5pZgo9pMYoajH9GM5WuNbyKj3GTHucNo++cysF0g/CLNFhaLtJf
PukF6neyrdKxhGpUtWU0eGvq79OkhmtTogDEvepHuzkD3jaxih18obz2aWJ2ONu0HJlfpJrCfMCl
jQMl0Sohf9CNXIIL3lWPRlLj2lI4NbwbMiZD3moC+NFJFwIX18MBcXta74pOaZ9M30B6qA9y96lz
E2I7YxiLbjBVlXpnugNVKHi8NewP0QZySdXmKZjEj6vUoyq5schyZNqGiUESMH8nmdokwBWGWEk+
aVUEmY0n8l2T2tFQQkAm8sWnE5bUeufUQArwbJk3EK4DHDMpw0RC29EQ9E935VECVmA2MIJbd5pg
TyV1VKKqsGyOVgXawuBDX9NXCY0zKxvvh+pgzohscKZlwOYiWt65zDtTIPULgWLarTHWFWH6vjTG
h/yhXxdydBqdk6hXzjbdG+7JSBE9FUopGh4hpZWIn6it1Au8EsQOcbuHiOjwHMUO4z6dK9dtfJif
gvjygtK7fYoSTtlHU+m4EO91MF4kxwX+3DCFinM0VztwupvtQkX/mZc2TnjgMfBIOK36t31f7S5h
YmlXCFvXrguhmwPtjHWbCNt3fMjUwuy9zILA0ZW7dvyPBZPCpB0jKrAXAzAc6FyENfqGqyloHDgi
vOX8BzT5edh13FpOF1zxG1d3vV426kgw5VGE1RVSRjSHhcBJjou76TFPtSerrG2j3bDyVDGFPxOS
jvx1f7ErkfVwmy3Hf5EGtwLH0mM7l5IoEfNSFX62MEDIQomC3hz5Z1vaVLO3YGlwLG3D4OyY8fch
cAua3nOt+jE9Lu9C12jTyYR4YH0NSrXp3pAHFSyS6fXJ0EmdDuA+miBiyS+4ZrS6Kg/RfO3k36Qh
TIycjzQHdXV24+ZV9roU3Vr2Bvga4l0j+Tkgmv4+3fHYQUqiXgDqh96kr4e02bX4Dr4svWU4TpwD
sJdcZhy0ebWmYpptyaeEFkNb3GZqGkdPLWmCOLo1bMzSDgW5Jaw72MRGPkhbcNXC1YygY/8Rsm0h
1V/SFtv+2MH5SN4TRTGV30sSVfyWnNKk2kY9P22OSPRdA7puZo9RtCveRQu0GMZbIUWCtamGu5LV
yjKvAA/7J+aSaEMt1YPqydsPOogqgwHqQ209G+nYbAWkxDXzb23ru/UT44UzVlfw4JgI43SyMV0m
nu7fHLlS4UKHU1VrKgDQL9v9T94b09aDhf6Gdi1RREkknHJ+oVRiJOlOBDLSMUyFuKhtoRwCGvOi
pOLnFjU6PEspTFa0p9RYU5T5m6WJCxYBKzqgHl4nSIq7hsUzS0F8hEj0CY/tL56fPTcNcUKtyFwM
djc9giENp0+9EnMTAd2nvlwcjc1Ami35FTq4v2L/u6MmGZQxOELHqPRtT4YpvYN+ZUNsgloHCzWx
9VMDp3T3HSPf70sbspyusf2PPR162UTkwk+Xr38E2hD2UH0zN+GclI6UGEsij/pR6Cw9OTsTEZ/b
9fFl0Bjd5EZt7n1wHaBbq+/qMLG1lpdrFxzfKidrfPO6qxv7wfobbd35qPQMzCwLO3hL7DKnzAk8
xbKwRvLDSwbeov0wHkv7LF2l4ime/4DmNFexxs6/lNBQllX958gDCToTtFEbA07EPq+9xMf25qDD
MWAnik0/wMusicoLAlM2XRHTujcsIIJl7V97SkT73/bV4f2CCL2mLtXBNZ19lEg97bEQLbhwZLRz
V2V/BdFcCi+Im8plHrX6RNA3eD6ehBZ/E9mZexqw9cxi1S2TFnISjmjIdDS3lW03UC8s+pKcSP85
iYz/OfObFtIDu61WxR/trnSVrcc6LaykRNxfdFpmX9971I5wlXbYvfWNDpKewDmYwQE/Bh6xQ4Ma
pGPeZmAn4r+VdT6RAebCeON1EiyEWRWKgb4IktLMHwbop0aTFF7Ulr3Q6IlSE00FYBTVUUFgnk5i
Am1CaY43oQ+CdV87CDbcoRlTOJVMRJT1ycvCbtCCufI2xrVxg/8c7zBHEBabI0XN7t88ShlqyABM
v9FHGBV0F6B9j4TLqp4VrQSpBcR7zvkid16u3MdOnH3RScFMyS1V7hpjdoLB+ufTKf+40dnVgY3b
1pYYyXvz5mH8RNV5I55Cf4qA4Qosjrem6hTpy5OEM0MtKSyiqMbsMdLuP8Ru+1s2hKup256i2IXp
qHwBZ2vImAAR6IarpamR6DSOtbSQhL60kTrb9u0JWZ32hTo/UUGKOzHrePLzBu9CYasdDDiRf4Zo
jbGskSVYCzgihY7ctM25bNOT1L0IfUPvj5DtjWndOZkxUd0B8mHFrnFLKC5D9CWhTJgIpgt6wJvZ
wSpRan+pYBkA8l2o/1YKDzzNP9I1MHHedxHUa1FAzc//dKzSuaIZyzQTHCb/gXGJzEg5Rb1C9X31
Ft+f918Nyz3iCFfJNYmRbdlZzTxiMQJHgLHXk+Q3xhzFBiyJ9NMnJ+olTIb/X6HJausgc4ttrT3C
J18hg/YwQVkF8ztqUi90+ECNb5mE46ToqIDGg6aMBcqwfQOtQIYZnD+EnyNll4qufoqwB9HPRKQ4
+8R+uI6rj2CVk1zDOb82DsD3Qie8IXsHqrGyw/FZu4Y+DwoSjeKzWheNr8uJeowQDNr1IylnuGfU
WpXEfAesHKjh3stYBy+1AayTBVWzFLPPfk4qHeA4qqiMtT9iuomLJunLyUPN5Z4i05efg3erVjvI
rceFbMBC6slCPup80GTotJbMNl34DHC5iK9GVLWv5WtR/ANmftnIpdymMYqe8s/tvVZdWZCpdrI5
Y7/CKkTQ9I8aKs6BFEyG+u+6mXzGau0HZehg3ap7A4/j5YtEmLPvGwtAzuwZwUaAeDP6xmckZxTJ
nuYxQXsH+3CI3FL1s7geMXMrg28s4GVbNynuMi5p1uuBDeZbNulaggKKzVc4V/xvYa7z8syWVi8Q
pFfwcEms5ISiH9BP/o/du3dYYudPlUPQebNlGDgyQ4NfhNfMLmqivI9C2WMqf6/V5RdzPqEJ4j86
ZegN7/WylsO9Gwk8lAp7sMxB4xk5VGrH56AwYWtJWucnvqDgF9XYtfWd729wv3b/yo8yXNckmfPo
hRZ7U4+2EKTAJoFFvHd4410Vmn8WbzlBBXVPYVo77se/TT43Ww+ZFotPtZhqr5vacxdG9JLUrhkf
l4qNKEKDPPj62TqYevcuH66tco57YE5FPtoHoE7ZxTpMcFVQHVUCvRsW4typ2DBADuCL9ILV/HG6
NmzyJgTWRIMfLtAzXgOwKBOhPkBIOsdxXTLAnPmB/ssGc7peoRtjK2d11fIE16IvCB92w5LPLg2F
MXz/Yy05b5wYyNqIuKv8+xB38hJ++Oa4CB/k7/22ovgBEXxp4JDtes7J3XXBC1mH94cf33Jy8Qep
ZEr4bLlZmsQ0llW6AfQp4AVJ6Vj15uSSv/jX+YvkB1YpxPWRkd1adjQWSK8aTw==
`protect end_protected
