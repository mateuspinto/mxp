`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
PVklwLKanX1OLU4iqzcIQol0Rdj87PJKN5bJKOoWPo4pN0XrdiybPCBM9D8VKFwipm4U5YcysVz1
ol35qhvT4pU1T7SDCMiobyxCTHOSMm0KyoEimWy26y72dSPrMC8h9px8Ndy+yaIQmWUxG4B0HVp2
u5NClySukq3N1se54gonx3uK5mHNgxYnCXeGrIKYyVqXwlz9iJR9Niv8XAmlICtMfVI/HKDugaCp
1K2HKjg9cUOTyZr65E8F9J/t70/RCGwqYP96W/am0uplE90NmTMjxmyq0vIrTJZULzkBCGVf1OgB
9SA8U7STIBo5ybDk363Q1uYqhsNF+nH/MyGFHg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="l1CH++dH+6fXXN3fHjiGDw/zMZPSpZedbEK5i23NHyU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17728)
`protect data_block
4FX6Ix0H+Rdw/ey1N14ULBVQBNzzrLst388+zCZL6F6ti6U1l+yjaR1zXNE1ikETpYxiRfuq8bQY
/olyU7I5EZJOmKQEg6ei/PGYdZyXIY/vbwq4hE62mPuJ5k8w1Eyi0nI3Q/Xs8sl/rek6o7VqX8bQ
UFAkes2SHVygI0dxhHvwymkZ3V5rZXQSjr4fK5/pASPmSNBaiRgKBt8D6h8g/UAC2RislKmwreTO
h+db6nvDRQkNvEj/a+Bj+WBsrNekfLmZ6dh/hSnhpn915QzqVNrbKzg2ptI7KRWCNtqLuAbABKry
+mjNYi20ysAlz1rrrEfhs1ZcWV1vKUGA/O01xeBPqNMhyRRUifwCIEitsTiFnruGlIzz+pHhp8Bv
KWXmCD1cUF2RKUImQdJSn6rKxtR4g9MF9R2v4fA+zy4Yz7kgtMkmZlqldQpUoCOHJp2+fwDTg3y6
LgA+IiTLDP6e3Tju/t5nTlQ8K6EtSBaMhFr78JrUJbzpLY80nQ2Hu71Fz6HWDZuPbD3xDqdbF4pn
IP6pBMnMdAC7Hekn3G7MlFKcdzmRDa9KmgWj/uCova0trS8+8K0Vu2SdKvHCJ/oXfrHx+g9Zgy8b
hC0/ddqLR4HQwPQgQ4WkXxcK1INOduYAY8NsO08Omc3EkMjVPUIIOJm2ZG99OYwHom/OxnpER9yp
DCadrCuJ7VwwfIg2pTRnywmJnd+Vev5wVQCrnYvk6HVbV8l8WYstC2wSLyFgZw9QQWGy5QEO168A
Do5mivDt9bk2lqLp2aDgtRwwJkaihIWUtcu2RlXQ0UoGc9V1aCebukpy6L0nTSE4k4Qfot8HWAC7
0Dl2Nk3T2UNPo6iUK513EM2DBSKYzuiVh5gVN4nEvgZOrZv37yp4Dxq2w43aIe332iT23FzTyvWh
4eGPFX89HG5aaLmSgjRrSesuF/whiPF6sj+Xho6rV5nqDtsxkge7QY+HV/3AoDsyIBXGdgw3YGF2
WQ81Kn0Y4e7IfX15JOAoIV5MX55QloWKbxwcVHONiohaMzJdj5egolz0DjF9oSh+Ef5AiBymKEPv
zIOaOhZVqck7oOoeL6N1HgMPmz6v97gJaNnH2QE37viTBE7jYmMk38JbPmihfUDQhS1JHTK3PGDy
XCGcxxf3XU/5btg3OiMiUqc0g6V9ewE7dgj61hqVy/gmG0UqPZe+04s0cftILkWNsGB5U/sMEbaa
Qk7XGSoQgI13rLCqEPI+pRwYyjMNPnXH5Asl/dCbg3pelyv8Y9DECMflE23QB+JFe+7VU0GJqJcG
LhwVzmPgYnhmu+hjqP8MdGKwUpc774mEL6E8Mb5K1A+KAK7ErI/Haybp1UNCorMKOb6lwmB0JqQ/
QlkKMUa5QP8sJCAbnn3OOTCwsaJZ8MNaaRlkKVbpeRxlCFgkPJQ2jHMBmgXevCnzTrDgzoOPXaKI
NwkN5VcKIcaa+c8HvmSVNKb9jIGmYKYJqfpzJHwYVnvLnzkz3Fia4BcmTWI2mN603XeyKpd27psj
8NpBSVukKyO9VvPxXcgOHZ9MnxoIvAUhl2KSI2UHUMiVK3YL9vme8J8JBJ4rSeY/RmbT2OU8NPWz
TalYaPqYVXrdyBMd9eCzO9rXNhP6elIJZkS+7FwtwmOwY77HfxJLYwmXj8zydCA99afMUs5FMzUl
zs/kVR7CpdXsTfEEZ68rROGASvu1ffpBsT8a+9i+iDj3wLQ0PDMeZECm3FgkmW3lZYSR9JrZTeq9
yccb81UcUiV+vF9Xn9jYl+UhE17vkJb4SUzm7NkHA96VY2Mx5qEI+NfE2nxy+rhJslQldSj9nbeb
HYOarqWddmVMvM+SQqonpBTMDJZtjHSwyc8BSWGYxZk9HyxC57BZ+lGtENLd9eimsbI/YyE+W35Y
NG5wYCedVrGYnTe578x/q9IzQdfxCVEf/Q7MIApuLI3OPRzL9ySdFsSEQj9jpKlwhFB6woaxUZnt
/etozqOVhANnXQiE9BEcy99oupioxFAegiU4ouUM/GvdupL4Y00+FrVrW1z1iXx/+kqQe/aRLpyp
nk+C6usx9R4wRmx58n02E6enMGaZB+XfQEtVuvSCqwFXMeTRVKuN/yrJ9jlAc/d/Ujyzl110C+eE
H8N23IMrN/jGBqzo9cwn1+UfjLhwRcnS30y1MF49XKUONRulyanat61v/631P4H3eE5wigaR3+Vg
EWLEq8BmN02RyVwHbedFF8J4wnxYvU58KurzLX3qKx+eE35Z6j5orCJEFp64cdlGMKBpP/yW1JPY
6dURaDuFMvK6SZY6PDQfW1HIEd4syJXXi4doASFITJREpQ2xiKKv6gGhCz7DFDzCYwpK5xaQz9yT
BDHo47A+9LVYMjcihN/s48y5mbin5HYAnf+Quru+8ishk6O7aAKjRineQnUpnEFu6N0niAxLPB64
E/ifHvt47PlCmddCKtJ5EwHwdOWWBb1udp061c6ILiL3ll2aTCMCrcVpeRAolfoP0A8UblhudWdL
QIgSzyPL2GBo2xSqeXOYE2pJhDGzyZeSjyGhHUUjwGZD4WywbcLGysu79jbrCANN5cnNxt7Z5LeQ
ycxhFeymBfO84r10KJnzoJMJY0bMEbxS6r0isuEWEcnumBsnGGW1ZtregsuyqQ93ppsqpiDQsIQA
OLTInsJXK30vCbU9OedO/NOIDS0Rq70LcM11Wy5nGtveAd1KHbS2NY9LVcrsAYg2pyMLBJo8v/Im
pPgtxaGwKiveeNkgW1l16bZeZC6lVE1d+709EzIuG/waVhupQtVk5m5TaQXigEeEuLxOzmO2ZjFS
jRBmIEewg7j6ubfRevL9Zyj/VPEhpXYE4eN7fvK+yCbk6m1SKTK/K1sBMBcTHOi46F/6ql1EpuTO
H30bp5L4reIaa0z7TZYQS9MsqpAOHLEkj2omz0gkl2mip6qKRsyJB878QLZdX5rsU/VHQfu1phS3
ujWA1uZ2xMIxNOsiBF8P/JqZYR9MbY8oQ6376LisOec8R2wORypE2Z6Hq1vP0P7BBF7OcZSaa5in
iudnpKfGpfYWYDiJWMXvy/y4uqne1GtJC2uHl443CrlGRqTvc49PUPgyoa29QUSlKvV8bCfVMtg2
F+dsjohlB1upgyG5caH8NMEfmPklrDWQ387wo3/k+umX/wvk737pzeluVJogJ6j8Onb33m4uy01q
Loxg6AA3Dt5vxcrHQK8rw70ONk3hZHZ9Ei5yzkHbjEI2XJaNubIzq/ktgg3QTioEHmOgpgUNJ0H2
p4YbQa6W5ndujlGPhmIyrIeAWRm/w3KnE0MMNM/q3bC3l94Y5l0c+kMosBuDeYaBwCrKQU/hnQYl
HB2+5eZjgAIjDggWhOnTP2S5Y/n4XnbVCeG43ddO4nagDreLyz+Nss2WboeY6ojLH+erD/sh+hDz
iXSGzItf/fCSgS5qQGzBUGjbeErQ1qvOjoI4SK7KAT98m6f5b8n2QzBXmGmZ+owTcyj8qK3GSzgo
oGSbU5GGQSXoqimr4v2qjbsPMeZfZfBhqSi1quvAsR8sqFw5Xl4E9h6QgFiI235cNBh/bQa20MKh
84VzksFLiNVgk/qctwLWjCsQhlTg0IYM1qHPQAfPoF8pb+wjfOk9o5uZnq9SrBBczTcZ79+jrlT9
m2lvfnw/tUoKN3Wgtfwz08DI9gLi9bN6XYHJM8riCT1E+tuiAqxwBcQ1CEVoxnoBfQmrgXiAvvmm
YJPcpMDh/eKk1g+/ZwQLch1NZNo4IhOtNpx2QdhjY+PDTu7ABEczdkZSBZ5YW5EmSDnd6Nkc0Bc7
nuQt9xcf+oK5TuVRzkjKqwwXx21qNlU4Na07CKLWJKDosqKfviv0FfLUc9O27dLBnZnLMvzueivH
U46ch471jTfoiyWPB5k2ZXQhMcp6/cZR/tArKSfV7+UvBcliRzNuXG3HNkMXF1RZmiFEFc4aZ1hE
sUVstD6+YSd5xl4DQ7RBKtDgFEvuMdXRSOs+LFmHTyMpMiNXP9gKij1W/uDYg0XaMQlJB+r6kVow
FHJyaDHRk701NWgX8Ib5YVP/uRVQaU8v4z7URh3aMYXBzQg5SR8nqULHgMYtdOp2CdqBIHAcGucJ
y4C0x5v0weKMjuW77f5QZ13/B7YakWFvIWyOPaII+6yCMQLzClnQ3MJPxvwnH+9J3RcTkGutJCGZ
kv/OJ2oTlI741valvSl/N5sOWVOslZdRiDmPS3sIMQXNd3mYRIqyz0OhZwMUJHmogjHkgetdjr+8
Z+ops4s9aMfx59UBS+5aLFWHrc2CjXonCz7FzigglJh5Pnf+UTVGYEYNy9FrLIf0A9xZfnq6zK8m
hDkpZSzToPT3hyFSuCx2nsgCM5zoPzz76gwJkrD+hQYvMnSGYcKh19VSqF6+gZWcyWclEpFhwQjs
ci/0ehtsiHqIuNihlzxgg7tlNuNbueOrMqZwKwbbRJ7K/hBx/UPw/33nCUPO9Xa7JYVp5LkrVEQ8
2oqgeVx/Tijw3ahIiuuqaqpkdfT2B/jnMw0KvNFhJYenTE1yQ5cTA73L5QHtyv9t55zKLWU8UtH3
6hmBa7fPjV/01cMnPldFc20+RFPqD8XWsk0rPxDirMdHE6K9xi+AgXrrXUCcoYXeR8861bik8EwZ
QlKIESYkSrnQwjTGry8NOfzV4u9TPdPNJbo8UkKJD1xCVOTZkd2422thiinXu6FCbtgYDPUMnQdF
tgLOu7dYoMFQFzsIjljJeG2NnVq9liCdxLQO/gCFTdiLrOVMRsC5CmLcpLlJK83RoNYPzE7vhj7l
ruWVkHL+AtpuJr6yRMT51c4QrQk9hZhjgw2x3Qv0UTHfDpqp+AL7jOo4K1fBI1BZhJWc1FnZWyKk
Ts75Pp7lSZ75uFfDiVO+OIH8LzqojhIWI0AV3Crsq+akdp607tJkvMbp7rW6DQTz/RiL+FGty1ly
GQYxkvqujpqj9q0lN6/xAIUj4akkUMCmgJ4jyDxNP/J7pAVFfj5BvFDffuXmhe0DHe0RxomBlER7
QngIxx2qw5v7Smn07cB2yzgM9cYEFtHtiA48FHP/YXg7sFkhB1+PYSXi3ZplP1+VsIuz8MLetDAx
3CWgHwlHzcBNvq1MYiBjh/8CiAa94V9RAWj8PzvMULHUoMiu772nturvmJekbn6dEo4Rz3SCU95k
fLuhydX7+draCau7Tj4abCLXneAHf1JReIStFKpakwaRcplH7Y5KyDl2Vv48JZvjkM/MeXDDJeFo
IoB22OH5+SOezE+ZtLgA1Bic9CxuuziV1Ixwtsv/nAYDg7hTnfnt02hD9UGCi4Yfoc7zluWj2j2D
3tSq3o1a7UxVs0C6f9gHmxzOPqV6c0SERQKLAEcZiHInKN6coj940ZfummAZO/ttKEYA68IVwELL
FCV6HdjfBpUwJ/iEQWI6HeoVeI6KwJkwFNqtL9kMT9xdlIFnzgNoSl2T6VjVbODxfIeZQx++FEjq
v0jvfaPcZjC5axM1KFgEhKTbVGm9krD23TvJyVblWW4+XoqB7s3/mal02lMWFzNsmpAJsvjm87Oo
RGpBwuivsT40Ri7mJafdlERiVyldD8wxrpC5BesQ2cUa0Qrgll+ZdeKhgTIWyxRKECqvV4Ygk6OX
EzVSnfo3Wdy5I1mLsnaAjZX3kpL7ShtfSO0bAP2V/h72kYsROf8e39KZPh6wpRnYwVKn3N5avyyP
Yx/bUYZIvNd12jtkvyT8K84GqW+kJNtaU9PJiXSHxB84O4pcMKJ1a1yjvF0uUyWfqoyOsk0MRrUU
/+eRoL3/5fAeRI9T/dzfdwLevlR6mHVeXspYz7+pyaqrh0dkNDZTPVV7Uczley6Y95jLAHkLmqwF
8sly7iRcM3m4b4NsZDvj41iiH9LfFqUO5tavhvlJ/xu3ngGMCxEpgxybKP5OQS3IKrYUYzjLEEwL
J5iTjZfptHtH1chORfnP1QD7omSJwLWuFxXgZvps0lE8iH757DdQpbI9Bp/ieriSh/36qIQiXgFq
QHgxfIGn6UfinfZ6llxVFWgjTGYA/uPQ6BdZGNUmp7dt9pilEffL3buJWTc2NvbYcx1Mf0rseRyn
aOG/e3KL0EhMw+ITBu3jGtsKP4vKyGtvoe4RsuEEQy3xhuqCWF8BlaOWGiud+F3DkbOBFtJokjZe
K4Lw9iLm5Dl8GtY+gPoRRqWEfV0eKJeiCBF2msWuRyBqqp8xQVjCIXti2Edz//HMb7pWQCyHJ5Mq
UMTthmHehIWcPRjNM8FP6tX8lDUF/Rv6SKrcCFO2oHE2K+F7MqgQwAQzOo9QUFQqKPPeW9/gearZ
8mBoK3oYN9kkidKKKMtwm0zq8LTTt67kQwyuVwoGGPG5hnSDKaZtC2gnIfJgxxD/il0Kytj71k7r
m5ba9DczDwKKOXsZIL+znXpr9vDVdP2Q42qj6lN7k5IzT7j5J7DS5LIjM/nJSMILoNh9eUKO6pyA
+X5C+TYFP6ZV+N9T3ewhwsyXVCvyw2dSfKhIVx2llMrcVJw4aIEAlRY5Js75+oUCGMAM5qt9KhsU
QYbEVQqmpmAgJJsgaOKGyhPg7X2Sb8x7FaADLXGTkPfGpeRMiPv+q3ueIzLlTn+fDEkgn+RDKl73
n5EfX9HHIujIaJJykWtNFTb+mg7jHvga8XFEYuHB1pCf8KEg79O6YCEbp8MPwWqc4bwxTX3X9jvu
XQ/saJcI8aZ+RSPujpvJZse3GwK81R+vcE4U1aOomCgapbtPScgQwtzqX2JtzVDMTu9FtaaVO6gA
Tcf2kSFekTmbD8WpQ3WMsBVi/EXNkjtrhQyQoR0D9udpnaFCdPayzGOpiuphUZuAsyHkoUbRcErb
UAUNxwK21P6Xqg4hWFk4jLZX9RHzrmKZl2HXF4jjsptIyWAYk8jKj1Ek/2kIumGc/vSNHofThBqU
VScbXaPNKJUFgf/TPyumJ/MRLL4zfa62ts/2uynP73GRZ1wkXoKBw1UHNT7WAKPQq3FoSJCFX3iA
QfRRRWHNUJXXJzChY/MBBAzH37nPlbRcUj+JTLa6pgx9uYWEa27M7O6Ep1uuVcFF4jEi67rMIjZQ
WzW4kNQZxrrTTdaINXCXSm5bz6t2S43BgfxhfOXJm27fdzN8I+MgeICV+edbzKp5u9SvRlvf1I5i
HeKlKWSMEqG3uJgeSF5cCoj9hqRFsxsaZnReYs4avQLr+EjcBcJWrc5sBY+LyVkf0wTriGKsUgsU
gNMAXGbJWqBkbR4cDO0FKpjeHHmpXljqJHKQZlfQPVe+rDO+72tXKVXmWSDvZOwTl+WAIFYX21C7
jOtYSvDSYKz32lW8nHmh8aVPseYHmLK2/rWvV8qcOEhFOnSpoPEnQI6S6wnkpCcMk6HzbLu4udZm
t1tm2ps3zvf6Uz3Tj+ikjo0haCCjNWYJ+b3awnw7VcQaAHTSpdGHm/NOwKXHlb98arb1Zc2tQ5BT
oKtrN6u2hNmAG9MeA/llSBgmxmB7Sqyh9eNscF9eFXAN5mC1ZyjwwBSU308WscHMkW69O6/XZTe4
IyWiS1MJzFoH+HsEUkjqjruLC6hCh6fJn108twWtLhMbEN7Fqju5CMWoWsKd+zG2KZnfRuNSCfuY
QA5NPa9l6wvTqPZndL/d55QkBixuLHggABG0FvJSW3ZOfRwZw6wwFGIPJbtMA5k2HnMKzAErVUJg
GBWBdT5F24t6s5MUDEigM2o5Wd5iRzvMuZ9KEKw5BU90C6CouvxunOE4YP4AVk+24Hodx6t8TPG/
IBdU5r1qGo0Nl/m2UET6zJi8iNgHQ8fVfEg1VoBGqCUISw+FGTTwBo3SD1OQu+R4Zm9QdQFhQy0o
db00kq9QRlxmrAWhzcvrRyOExRM/CKGHSPE3fT+HInY0SuQJm26n8x/msGZW0/qKLLsE6/ikEqnS
GvxWZTLTrWf80qH3RcgWZmrr7G1QS1Cx7EETWW5alv7FZIUEFSZF46g+S2xQiFSDBEgVrlj1/TGH
y6SY3ZSFYCw8gxfYy0mTZnoEiEKVY4Q2bq2f7sPvvUpOkCv/PhH2FgBdM1RNQXVqbRJoirHs2p/U
P+UF6uZnj56xnd0xWxccyV3zpNeyD9rGbXMUho92XGheVVNjsQyZvtzm+nS6sdqJ/jzaqh0VZdC1
4Wz5MllNRGN4ZalA/PnjzrhD0mMhNZgj8nlhWZf88aHhuwD8eWDQ82Utp38KxKhBbcbv/26erep6
H5Whturb9qzHUuYbSyzKGbQZwwjX2Dj+OgwiVCfMi4pgg5IQ1+OieDZI3iXnI5QvVisL2vpz2yoZ
ZfOCjUi1qiylMkK5972YOhx+gpbsqdYTWizRn9mGVaesBHSfcRxxC5MgqULE8C9GPnG+wOOeB9kW
/D8NvZYdo4+dCuPLYKIhs6w0jRd+f1I8wWl3nPXwixF9hIZFSRg9eEX9W9/Irp+xbQEPqj5vYcNH
XPRMJsZYgGrftW8HQck0yvTBJYDVukjJSsduU7iH2etZ5nBsNAH94Nk8grvS6sOP1QsotBRuEk+M
HZyYA4UgGn7q++6ylSvnWC+1jMmCpaUWFiwf7V2fnqvUmno4ue63J8n3yfHf4LnR55YYVmIYFdwb
VsjuOaDib4/CF+o0eNHKvlSpAB3G35lN2mz7+3/P84/vri5ZnGZ5EaVn2QYgx3ZoD32qVfB9lbMe
4798OrJ2844NJSIJF4m3/tT+3SGMtbgfOICq3vijHuMrwx7pdl0ige2PMLw2R+9e0wwvBjpkFLVN
h/JTvRw8kdNdrPLQgZ9kHpg3Ngf2WmXCj3sF0RKwzVc9JzS7hxPZ8wBTif1/dIEdZBqHGzFMg/JW
Vn6haGZEgLpmDQojS4UIEv8dw53dw2smZXbH6nHP6r3nhDgp22i0YV48aihlgLmbMJcaYfZFQuQk
FgsgdxlhU+HjEjszXgMCWxaXGiLsJTgOOT0I/Ii+P/4Bnf3VxD49ruGC1rOO5195WxCoNE4pNg0f
fwAnYEzorot/QAxpmeJVb3iMgjPJ8wajErUGXw1FNWI6jEFb9w0GDdxSfHQDMln0JY7NIzm7taIi
mmgc3Q7yYQ3HkZTGclsWvHP/nqwlMRBWFQtxdQ2p/sfgWYAMmsJ+VDyxTka3yO1mnFa497+UaTAg
IMRHh32aTVUZV8TWgTStz2H7VxSvG9yFta+TpCVUwoGel2XE7ws3287BNtFnPuACPsLV0AkncI+1
/m9XpweesYOcqi1xvVSyKSaQGwxJO8wx0BDSV7OeVLb5uKdZruU698lzvvG30V+J+S8YC6MGh1bg
YOSFGBBJwr96NqRNYP0XUae2AFX0ysdwa2mcjPiLyB7lGfcxuwFnL/zPVD319olsac8zG1uybl+3
oCY13ROO09agUPekb7Lsb5uaprrTT2F3u3ZAlBnPFKFWFeHNrvuKiZFiBUVSxxltuLP8UQfkxPlk
InJwii9zLEXGDKeZI+KqWhSb1rMxLyLUV1LixP3SOtZ/s+pouTc7ZH0r7fzTxTKKlVusG9t8GTbI
5uR6lcqMg1DInnlxhDRnOA/LuPs/61u7mS9WyL5lI9f/sms8T4tTZTayi7jod+WeooF9F4sC/oF3
oNVyNqyHV7jxXx1SMqfIOwCdKUeIGKWXgv0+JkjRNPaNLPFUMmzJxlCEeW2jNIO8i6ikx9sCnREJ
z9eeuTC+rrJPugyxjryxz4gj7h4BCdEhaHMbnkzqjBNcAHOqaf/OyV5HtZXCKw8AsXN/B1t5w6dZ
90b9aFYQTi/ktW5jlWXhz/y9v0hIbBtRJapwQ69UgjNJ0IN6xvFLK/Bf931ubXX6WtIGp79H8jgJ
RDwgQQIU8r3ujYJt5MZfV3pRrRRxNpzQ3RwpHN+bcKy8+E4ZEy7WZvvVuRATsmMY85c6sJpF/Azs
L30SpRdNdW0NUZCHAFABpKqaA4RVcdHTh0bCBv5l/S04mP6pXSZDN4c1v4F5n/QzrqcTtRpcuSqB
HPP/20CCfBAZ9mxBllQaJuYO1uaqIteH2UNxuTTcpJPo3DFe4DHdkKbnarxTNTEaxnyZdiYiZt5s
1HtMhvMvlGrWJMoy/Ypi7zEetfOtShdQPhD64GLYTA7NAk+b4Vz+TKyU6YQu+6hXZQfzr4eEU/JO
7AK4+WVEg8p5NEx56FfsgqRoYq6a65cC7Ykzuxw0J5FMYgs2O5n65lZk5KNoYXSzNKf1IzmuZnUq
t80J1eMq/3tXe2Hf/sSSLq8xllY7kVgmlvK/7Y1mz95+sybsZQ3vgsMgBuSfPvyVHawf6W+GO1a5
OKtes8KFgVXaHkRhNKja+j5KqFvvyuGTShdE35Gpc4LI0gLfMTOk2QMFLbEPzINXMKU5U+WnZwGk
22B9MQ3B/f9gzgR5pV5Hui7UR8OCvOfqeErPtozXg2OIczdQBmmMXXXS3cOMJ6AS6uTOB/Bc3sKl
+efCDhCzD0vdI+cqQUF1yvI2sjLxa1jZZWCBdv2K8kSBl5ydccdCta2E05W/R0MyOieqzPW2YRHA
W6bwCm65zqkgOpOacpJo15MZAIvQif2yPmCzcko+YruSXBOH95CJ54bpq+r2usFWQdae1h6D3TF2
eU7jfaztPfZU/DwsISQOt8MUSuVAWJAgKR0AX4Cca8ny+aMCduEN+1ORrqDokSMrh6Gb0X+mlNRe
cwcpYoO4/HlDxH/lKAwOSu2nnBfQXVXjjDhbOSZi2ZpIc3ZsMBrFVuMMti8OIJyHPfdwQj8QgLRm
DaNP7omrqtDbvIlvsS+TW64jMZZgeEM3WZ2KhnJ1Y9FBQMGv6vddk9qyCH/cHkgL4/8F7y1J7YKv
LQrY7BXfL7D34TGf4fgNmLr52pKHagd1F4XvvsqSaIsYJMfItCzp3iedRRtM1gqD7zCgTYnQjf1O
16uiE6SszRASai+E7G2Qt3bic+zkGS41dUfNQQWejujNZOnSvCPgnxVH76X5JWOa8aIBNEmbQZKy
nnZImYQseDtSaCntSrYQ0Se2JDrP7dkRzQmK+vLQdyecqJ11VeeUxkPaR4jJxzQB3rV389VSHabS
kQKOUjjAYY9yLQp49zwaCSOOPa2bl91sQxz2NnY3eDJi7tNutq3eG3/CbjtDQ6E9KlmxotEvgsPU
cyrJRXJcQo5W+C0OMuTZ4G0BnMvwfokBPmpXHZaJrMFR4wNG0vUy1EfvcZUdXZ9bIHRZPgM81rcV
DWW29H8UhoRNYUVlQSYsv4kOyEMaZRDAS3UROOGH/DweZJ46oLRoJOYBDUBCPwCL1C682MO6UdXq
OMQGomeuyvS1rP+Ti35TBgoa921xMzI+zHFX+SaAcNHLTzC8ipayNbp3X1P3Qgt2k7ExuiwAyGVP
drY5Wqr/2HlnJciECwChNghZaBFCDikrtkDFUEPTBpGXNhMxiyLSPmHY8aQLZSLbiTKme6SlgZ6/
NCFdhrBrU8N+hzG2n3wgbJhy+Pb59O2++sC1GSJ/BgYK8uH0UqFMhF/1RjCYniRKTc9pVmI9A7R5
3Jhk36gaQxUmWUw440IwrCgn7DfTlbr30c555c77/BHxrkqRyK1Z7otRphJR1eV/A4/NVF3TQUg4
6NyvPjj2FqChMuUOw5OAsRRab+7eWnoLbbi3jXp8PLQFhEjGitPNA69aWq/tWKTqdI7+js4cZZHl
xknG8hLD4LeBz9dpHwkXarNxEI51AeScjE+vaBRam8s3dAvWrANHiibGtg/G0hUkI49vmXay6lUY
3fHU7zxOyfi2StL8ZY/GS312GK7m9Nm/f/vxXJhAPCTFYygQ69qVdwHPd4d/6yWiQjy6zZn5FUzs
VYerehpDNPXk0US8zwgEMNycSMivoW1nvvIWEbbe04+c1SA/kqR/dVdDG4uFlwFkRt3ez2lCIEkU
X4bWFF2KMU/XszeEB1AtFw81DSmKwNK+qUBFjh/V1KOlh3cY4S0kMtaVvsb2f6lmG+VRPYD63swi
RempbowHF6o64AoiirMyjwD6fnCZQz7rP+vmF4zt//HtBrdiG3M7BJnfR2ZZ/rpUU6TjoM4ITkVe
OAw1iBeitjHVdS6J1GhdhxDXdfpdthT+Lklrr9q9oHYrJcMjI1fHr2AjDRd9P4Ma+tMWggtHXHJS
2udPskeRU31sFlbeqM29WWg3bgcRm6sRJD9KxF5VoxuCQslAcv+wSKCZdfflhhp+tfrzCZ6YBRY0
Z2q36+VTwBGw7c6VwpyzzEKVVHj47rtD1q1k7UO4FjVnObWoUXaR0XIeCwAneCp5VgGXO4nRQ7EX
CwtXoyCrAk62ITZVwAwHKGxH0ZIdLITKmKimdieA67E7fnGvU+MGWrYpXGbiCvR/CFen16Xy/h+V
TQU31glnjRhM1/AhlfUSMZLNcFQxK7KNey6a6BGbCKboYG9/HJinsq9B+6NI6+9S9e/NHpL5LveM
3BQlxJGgETD29dljA6yt0KwmW1kHTgWXAaGBYB59BWISKNrYt2lMl6s2+giwV2pC2TksMzxgUt8f
fUJprI7x9ziI7+6bNzP3l0j2RNbXj9CfOtZitkbZH7SdTS8afKyeFgd7HLkdtQ4Yy581W7C1DkcI
OVoL+mehTDJ7HsPcV46MGHVh+lMXIc5NFgahH7FdjWPvdzQUo2x04osH27yCTKm8Q1E1fkb1k1qO
Gv9re3VVr2b2NP2Jaow/TABC6DRv6h02yKLVF59Pdrn8aWjQOUolmB15iqAvT55P65U7EC3i2sLW
xA/bBvR7IXr72G3+8McLzSsupVTgJDFnsq6JwQcIvEQd59f8HWXhBWsAiNklJlfTDcTBwS1eSBlS
SXKYXSPwyGOg3qUsCYmmvbqWHf3pYhq2pyrjssFvhij6BaLtqRH111JHbj4h+QQdo5rMVPHEeKMq
NOtdMxFOHq0IJRNBXIBmWQ+UJsYgyEj9z7krgvol72niS3W269ppePjtEalzUJsvOoiTwlx0703r
QIC+6Mm7bKVOKTVyBUkgmeUGNI7VWORk5WNdHq8LVJTJehO4ZRIOHtxyyBp5OnlcaFlsEghgTA+1
j8h68jj1RL2BTQweDehU7LWPli+Qjfvoh4bsP6OQo6Xa+lnYPv7nPioAMgPpD2C+NZOyCR6XiNGR
X6I1+I2iGu6R2oyF1ZkYCYjL13UUuN3TEBfvWMyHwoSbvsCwdepvjanDvR6Zvy4wd0XCh1f08fRy
qYspNpbq+z78q/gfMGLkkn8iMzHStT8LzfrdLSTwZmR+r6iqc8QAUh1AF/CTJ5cjNMZTceOaYVeR
vgx5kp1eK31bdPD3EyQz99CZ4oe5BQRqnRZnhZMQX34e1/6h8eFzFf0S469Bo6RQM96hK3sA9pgv
r2Um2AE2CoD6ca/4NMWeDoHncMc/o+xGXK561pjEWmMJi/PzKcSQcCkdImPnGALXFLwLp6vjcJiR
cA/e+cfRuIyNMlV4+TUEdxMZEPNwFXXvDpvEfv4/dAig5Ie3mvDPUQZrIBBoc8Laa7z0xdzj29Ow
PzKjMR8OctN+NhPlemIHrsrODgRz2oQDvZ1tQpBiUZN6oCg61CcPEno+fGol0IdryH1pQX1Uui5+
6ngtOXDR7WiX/zWku74PgGdXhzH6QQ/fqWtYjTclTze1RafyZ8oF19KDAAzikeQ5gywl0Xh27gHp
eEdX808kdnAGQ4bsPuFaOpnZ/vTLzoK6Dh4vQLg6xQ4sRB9WGwsFhr5z/C+hAuf4pJ1vBF/8cMzH
sjEP2dQzDPiqZpRy3i/zQbagwk4hI6LuW/Na8K5ormYkrVzxLpvcIk+Pt3LB+S8pTvd3jjBboTs/
lUO/YvysqlxjwCGOcJclrXmtDpPeRn93+dCuWQ2C3IB3Sp+cklK7OVKRtRqnKPSB4/HI2t67DmrQ
db3htjSv84sfEyshmzRMY2pq1M1aFuZ+Z9WBklfg4Jk8te3vCFiVn4dQe3TJvBnxQyFngpMAbljq
ARudiDydcvzAVZ8pJfuUXzmhYrW3L/7u9JP3pqfUGtPmWlRzPH+XNpE293XaacKFjjL8O3kS8HD1
of/wDATZhnKzGDTXiwaxfu6J8BC8AZ57fLIAqGwkX4Pnl8qbURZ3JHdTTH6Ht6+U9We7V2lniP4a
XpMEquJSm4iXL8ihT20d+7t3rw+4cNZ0LjJPfD+ro8x4ca0Kn6Re3lTBtwPSi2d1jnf5rnt/CBXk
eI8eESJC1n/LyrTsBRMIfGGsIIlDtfNTUVpGZBFpHUsICgYFRAqsPa8hYf7YSS4yyKG8GDWsL5DM
gyA48tY8/Ln6fphVkQ5mjSm3H0FG+FuHVg/oX/E6t47PuW+ls6Um5+ZAqKIosl6jv48GoBmSH97r
QQFkng9BiBPDSjSS2VsKXpAFkGzrN024r54FMQjN6pBdldqin/LJptNpXgGOkqeJi4xWEFR+TE9q
zq+JJjqUMjTmaapJ/7dyElJekC+je0B2xyvGkSPnQK21j8R1gUoi41L93WSD/e8gT4dcK19Hc54s
1oBNtCOfK/nHERg/vg/d32v0w+A+ROPdcl28pZqjrplCLC3PT2H5f5Pi09Wdck6PB9be31WgOWpo
mGp/zv5ERX1aAXevI4GHVtWQJDHWPGxh05xgXtjHDLJeWD6DJoftFJ+sPMzMqhcDtWsBbUm+F6IB
hF9xGpCjYxF6+qWFLlNYF9t8ruvJ6k5t0ypD/ntgAcMcKmVAH7PNGMKdjn/WNknziMpnTAVMO6LR
Vmd+efq1JUYaa8ZB9WUk45WNA6ShFtQpElfnHzbuvrltTehMIsaevHaG4GKjV1J5qtl40ji4YHlE
nRH3m0JSEcOHY04uuxR2pbQZ4Uc2CMSM4bq9anDmyB2ptj7xQJxK2x26g8ckE9pcbsx9tYCi7Hbw
Vn0RZLfJDhncWLuYgCs3idqZBE5cfaiJg1LOutr9Rd+fCrJ+FrUXnGGyJlZjjNsvhBFmjU2w3V1V
3j2C1poA9QWtG1NUf4lfaW+QbOiiebhXN9Xb5FbCvMTneS5XhuqpWC1nc5gwxCDUOuBzsnMijO13
pHo+9SD6u5IaIX0OImG5s1B1wRHKCZ27DdhI7WcZeGx6nvBrU1uOh0LnS08eQd7oqmXZCi1msQ+1
N+Dl9L9MSsXqA+CXA9ssoIqz7+yTq60IYK/7iaGz4y/ZOiHhgy4Pi/Sp5WdcI9dcOPN9jR4kQbqs
+3hfwwIX+oDbI0i5gYCSnmgLHDFGXvtxTPUYWhQFFEGK/jXNUA+S2DjDgQmf8oPbtmInDDxOu3ro
+6nwZHyerw0wUE40l/jwRt3Sz6OicwPUaIefjdWLxX3vZsIVzbJkgs1UaviRPaxdc7gobNXgkb6u
MhqeRQjkS13nWktvLIhw/S4wDAwUF83N80lcalWo/6WDfh4n2OUbI/XOcV+zAyiM7iqvTO94j1+/
/sJwWHXXHR31JJiSXntvpJ3Qfzp2DWVnLIdG7PQb8FOsmgFVfO1C0CGOQJseQ0ljRSIki4ACme5S
OlvXXp85R2R01nP+jnfnFuIlROauZEC5Vn8UQFf2OgnIoV4OV6HfhR6rN9q/yPwxRUh1KPLd6GJT
8oTryWgMXocvMPTwtUjf1sLozZnFPOThdd05NQBaPmu62OnC/HKMjrRDb0MKH8LZ1YQiSh4KVmsG
HxfdVPn3/lP6ENaBBEWPAPEIytX6vbw1Ts/NwHWVTum1BkkDMBxEDyyRyiH1AIiTtooZUV3rdUHz
u5gcLsVWC0QKHI93Gj/06prqgFGhF/SKIj8xCROG6b3nwoLeX5HWAVpnNPfFRPIYHXNFdMW6PTF1
IPDgowcWXtVjSYajO0X/K3GWwcvJIZppkvIk+D24zINyBJ7bLs2W2FcjAyf0DwY45UXlVSYKAmmw
QJHRujCue0XxrM8XTjZO3hoEimQGSP7oW4tNNv23QurAMSsaAu016xnSyVFZe6utXTECNTQ7Wssb
ufLakObJyDB7eBIU1NvKyMbmbm00umRA7zxJiH1B9li6J10pBoxAj6/BLpf4G89FwKb1a5BkqK0L
T6yrewFLMXGq1QqdhNIeK2E/OFWMHl1ZGL+31KbcqwRitNmltMkxu6x/O/uU0d5QpOn+p6uwzzyN
Q/wLeKmXHqI1JWiYfrDLtKRDEVim8SpY6t4Dk+Eu25/sV9vwXvlaJofbe51a/R5oTbe+THmQejj7
XrWHzrAY/eLT6mzeZuCzEKYxKGCdsTiIRJNF7NGbwLd0YaxOnBcfJDKMw2AuRCQs/3L2AFLGaWFF
D3+An/quNZ2N6D8AIyD0hl8OwHHSJuOrhzhf20TizOIbzig5HXF7MIXRYkDT0cIYISU85YvT/6Zv
8+QX8zPZ//sGZotRq0VKXokBlZo14AE+4S6LVG3kQvVuevT49zmTBuzXos1LnsqFnAswL1U3BFx1
+UY39V22zAqsoLGCWElAJd6Rm13SXlimg7wyzYsfWP42+RXHu130oIc6Hg5L/+mKMovppaSmcCNY
1D2NpLhBxrLS/VHpD42PNSxUTidWlyUWyHfD74ndcPp3nWBthjB1Yyp/ebqHPWqEfbjfQUpV5o/O
JKlWJsoerWjXAvAHUxkvPlHk0A12n8WYmJwQ2DCfvjsOPQQqEAcvxGvx3kuiq8h536IwmkyvqhLY
OY4ghn/8xiGR2mVgy3oAo9CT+hShFlBpUNZE9NogRXdlREvYjcR3UUFIejp3WiMY5jqxp4cg7/fY
td4shPJnXrs54HeZhH+i8lwcSTxeDjEN0HgwvEEbxslF2WYD4TaImEOXME0OkNJw5BKYSkwFMAVL
ACBciQN2XHkxW48KCtjDnhJrTU1eCNQedOkrCJ6U6Qt1QICoAI+sBEDjwi9M5RNZnvaOi29a1W7B
RpDUnADd60sBewoaQASuB9xe4eK++9VMmbq5artA+MVLck90vuunAeF615SsZl4c1jv1DIJANma2
nzRVNQiJCvNO8dHM26c5z9gBkzuD5LmQkpLoaRHKxEbsxalJe5MuIhDQ5kTtHeNwWIKkrGH0vzSO
AObsQGW3YRJ7OA8H+Ih9cZD9J6A6J1R37W342PlUJuK8G5/EEunjomy88HJe2OS/C9hFbntHqEJL
Chzjvft1LpUFerjnnPB0hXlHegosQdWlRobwO3ca8gWdMbK8oonZKZqzAxprYSswZqyEIwGUjlqf
TqV+LjO9Tx7v5/JIJMC6/qNfcxXq7IthZN6TrQ0tnwza48aBhiAobaQPNnYbgwbrUIpEOMXDrazN
MoJ4IsrU/G43AhLU7XxIDWmuLKOUYnx4y1Vqzo1HXGX+R3n9XxLYGtNG/5KN3eX+XgdEIO5giyk9
seVNqQD8RoR4fxRa60qlRkivvhc/l36HVBIw7xiba2DgFmjALTeAY/B2on84IJ0zLr2ohljiyb8p
EPd7qyFam+ggxkdUtX0l5GWEaPS9ARiJHIINdCUGEyES8dsO9xIMe4zOqkxGEky12BdyQifT+xPq
qiQyS4x7JCNL19uTLhE8HRhAAlUwWKhMlqv7u3nDo7g+6ZfTo6XlEfReZpk9fEni98OMaqfZS+VC
E7mocCpa7werTz3Y0NgoUfVfCNzCS7CicxEX4at5/cMba4hxE04rvNdg4tkVdMNs81H9PXQNVWoK
fb1+DjHbqUJ19AGSzgdh64Fwg7ooEdJK4V7RYh4KBBS6idsISRyDnSSahsrxVNe6gN5+MttJfmj6
7L3yXGL4OpKXYfz9mRxtFDElQidkSPN7DHEa5/8X0onNAMlpfN2OfojJ5ewXqiu+EuVVoVdPrXB7
M3wEqGHH47GwvbLSQlWmGBlu0F4RGM/NW2av4L8kVZhvkbMCT4cPjVJWdB7D7KBnh7DbYMyVfcbh
+5M+hBNK/NPdXrTVB4llSqFgm0lBKnM3yJaBV8V7VXh6EDjT6A/ciGnPVHSrxQznkOYKwxtvKvXG
yDdtfWsvk85Flrzad6CAIidReLj0BDd7dDYsLZah6WBzbdv6bkmWLHicYwPcWzsfYAmSZc56vyjA
x14Qs1Rcf2lAZP9c4OaBdeV7+HiSgSKHx0e5umF1Pbywz53HU0xy0lqDq2CajuNjWB5T4hBpxths
VFztM7u/eGEb9NGv1t7Hv41N3j9/WknWWqmrNj6k/sbcOwiFFgCVBhllTuCKuWYjv8Ph5jxGQA+I
MW/cX/j8jqLkx2MJ30/0NNo/SIfYv+TRR8BpsVBqEGTApQ/UHC0YHInY2h9IxSKN7hNfNxwQt/TM
bh0Rs89pjomZJbVbYaVgZqNEI6sRRIi4jUnwmDzKn+hCkFXnMygb0Mq6K6BKsgsh1Cg/ztGg84cb
TPyly0ixxm0eqKugktc4FgVzR6RpfhfgAjmNSsxyGFMBPAxHyTx8f8+Nu1govP/mE73a+osSF5dG
2vIqnzseIUeYR/oLfkk03YOZxawmzgOLg449vVd5yBWMK9EN4ou74XZl7edHAgql2aBd/svJDS3r
Q3Dx3ixNf3h+oD4CyBX9aXOVQkKzWoIYzPsRy5z7WB6omkJzvyH0DhdCi1C0G9CEIgqe1ZrWygUk
6+8E3riyHQHUgM+PQEK+bj2+Vyu6vLKqYyFxf3ZNGOpHJNg/U6yt47p6RevDIfKAArP9y2mpiMZi
jgekngYj/KLiaVKUMJ3ovM1n6IFnsBuSGD5z2hnJbHTBrr2/zVkj/bAexrMBXz7p1R7ju2u9v6uo
WOSBa4eXYELBeNDB5qINFBG6TpgWTnEOWQpy4VsEGdo/5CwdlV+/hEJ7OuH0GQQjDruHuLPA2Y0n
haV9Q01G2ELT16NIESdLCg+plfPj8MZgcezREsK9BnypiJEMw7LEdsndpEQzNuogocvNA8FgVP/u
02m3AXb1MTIKVcmozN2IV6yq3VxdXF/D3rJxtKnncqmxSKDq1YrdAEM9J+WUq4BRtE8o98b8BdPZ
UyO+9wUcLRvEPMKuEnTIjZKMKpn/SuWYJghIoGpIDU48inT7gwtkZH30e3wIUfqz7jhZxQaKgyV9
IV8ctmKsgRMN2FZzB4z198nMHmmxOsVCHlHSnz+9onl5wk+YjJq1d5fUmGQcQQKS0o9/tGAjF0yz
oOc6AWw0XbDJZ5qrIEPiZpDTBuBkeq5pLafitpNgafr8NneE3ExGtbOzSSAEeFxEP/fSxTmHkxtU
/LCDpm8sW0gwn1AVjUTmkwsnvdeTVcdV4byNyKnwOzRJ+BgEBxIak2GYHw2OZ0Lg4adMHQ7rXyRa
lMX85RQlWWtNEQbsm3D5GGuWe7ors8KPIfn8jouDC/JghBZuOfZ3+DBsYohlCw1BEiti1iOcQNM8
x6ab0PS8YOaoHIEOnBlPQzf5Q95KlQZ+f/IUPdd0lznMdkq1stklYuJGtSSJgCUcsOOxJjx6mGy1
d0mm6LMSV15GU1A+vWNmoYcMLi8kHYe4ZOrFzrtfRpJPR2f/1yMR7WBmUUoXGfMmvl8JLWUeSFUU
Y8xHdobxm7AiBx55bJUJ5WEeTAFXpIyEFyp4HJOFzVkxxF93UVw0qx9y0wmEDRjGQf05IJV+ZPxh
59NPmNcHGjxHn3YLV2RJC4VSBZKODyALHkOKZDMB6oOS7x3bS7dFQSjUU8zK2iR8JS3Td/JUHgFd
JWjaffx9NndTC38ta1pH5CtVwyiZkjotpKYZuBU0+nbiYUEVh0HHMcDNBfJCBjLbrnr4X3LviCTc
5iuSj9PPACAb0umw0sjbA4XUgwJAmHz9ulAkM3wBdH1Z7FoVbw2xxy2SRPxom29KYRIykzCCe/XX
y1n1Y0HV3wFNuzci6wV+AY/SIIKPzOhrYDk4mRkyY1k3feqGpVWUnoIELaLiCiPgIJc11DQC4wob
EIzcNGNSfJTHLTyyNOLF4gCFRpH30Tg2pdhE8caUebxy2L6NpMBwUEuo38U2+yN0nBumuXoqXW4c
vptZt2yTAGs03Uq2Y3OwKaBNeu7IcbRr7mvOk8tmZvW2n/k3ZEaW70G5r/R5cm6aHUgFTs/Be4h6
vqyM583yzr69vPGJihY0UbZniVDu2irGlsSa0gnrhxgaCOZ/1xbTW7NQBsa3oO9d7xVQX5brHI7/
BJPbrOJbh0XOPxspHM4H8Ct9sgg5FR9wv+tQ6PgulweOZvNjp/OcF31hEGtER94HiHO3aPBsK9AG
2y25oeh+uNhSnJbpbr4AEYSJbDE8bzJs6u2ZgeJ5C4g7cWZQQ8DoO0y5Q3hKU3RnibZA3XG8hGtl
wDgRoyqniKZCNiSVEiPHigHBedyAmCy4J+Fi7sLt6jCJZNRvoEP/4GP5twhl0iSZlzjMbuSlo4eX
SkAGW/2IaU+6KulSbV0mys/6f8LfHy7yxUOHe02mREA9eOP3ypkg9PdGgKqoWBKWycD7kqmsyW3a
uZEjtsXCz2Rkq4d0PstzJ0EVQZ6ZKwl6h+C4yKDfSBa0wCumBjg7Uc6+S+HK66c+YLS/b/qBYJpN
bEp8c+uR4V6KAyt8OED1bd8H53yrfua66/GpHRKEPa07naSqwmuezchQNhXq+4rjx35PsyFleUGP
7sne5mZYmuVAD5SemOUxtmLtxfADjglAR/CyzPy9Y0xuDIFIyQXNyFsFr0H6IXMvKi+W9G7v6RuG
dlRND3hjlSRVvm/7HykU2L539WfvALP37N8uN1utxa1G7k4bau49/z/TdiqOu8hPxPAG0JQ2cos8
7ypCNW0SH7AfzR/srcqJq5gfzCKUMImC5b8iE0dGZsjpIW5x9nwHI1wDcgyVk3FF//mFjIuxG8V7
uflVcbHcN6BRSuOn8UWbtz5iUVJdTp9AvEiaPzPuksRbOa5ID+FSJzErQT0oHS2otW1LPQ/BtW5A
R4tV7uIXFd/zQYdZiBecu5hV2/y88xrjysJJGQrcZD56z8z9ptd/PxifefaLPgtRpDnj17IcdgOv
Z1nD+vlEv+lmhe6lF7Z6yJyy5YQXWLq16ZU8v77egzZ8/TWuR68zYxcaOwFRLE/z14gYFqHX84sb
z66+nApGP3HyQhE4TxCa3XxlpPXEpFn9Ag4ShgM3ExNMmD+hRDi4cOneEeQkvMiRDKukFtBLoZ3u
Jbi67f7hWJkzDNPhyq1ZBqhGbP0ryohmjOTzHQQ2KzWXTut05AD9yZyxhaLomoSHlYccW8hsa2+L
VEGXoKwp8bDGTvYKvFPS3RpwGGJjY3EPRKXVOFCyx4GgBVx9mDZpI4Af7mOlpNivqX21ofzojOrm
9uI68VjCy2tMMwmk3m20ieE2wHelV/FsdB7B4nULVWl6Zg5AkFQViORZOoUY0xf2LJDdYq35l7A7
8IL6vTxlv4fv8QQ4J8GPZ01MlQZHedX6Aea0nJtOZunIzKauZ/1Z672OUGl9+3NUBYlm7wb5ndK/
lRrpZW788Yv/hHKsq6TLb1yDaSFXB8sNla4KVcIGSIZVU4kIQMF4+vOGVj/esX7jNSbGkBuHDo3w
Uls0gwNSAdeHwAVsbX0ZsdZIQT2TWiiQTgOKMcoy8OcP2ZT/foFhYTXUi2s/cZYGIqd0lioq8Z/b
eY2LEW8Z6RoyCAn4uOHvLQI3twW7CLbFiwnzA54i9wJtq+qdJVHaWQNLPGyMrBQ74hKysUTugLlP
M2J/XASwSmYsrO+tB02Qac++0MKXbSEeN2f/9p9KToM+ULKl+5Rwgu43/i47b3oF+xn8X/NzpbCv
Jh/L266RslxFd9OnxqbAOlLBvB/vohfLaJ2MeV/WsNH7DxEJRF4LjZqIwAxZJRCzIwFWBztwDUo0
cCYTN+Bp+sbB4CBDRxZ8+joMAVd65JwpGprv8Vp5d2szCU7nfZ+oRZnYpgZlEAO1qDdzbTEmN0MG
LWJnJPWyh7vqnomv8WL6tDE+xb7A/p5M29QXJ0u3WJRhcDkXLiENnraFUrDo+z9Lf1MhD9klgKLf
H8GjBAR8fQrVpu7jXS2Cm6dKccpOcB/mcPuV6cy/1OHDoVhmHTmaMBjAxLX1a3HPNTYAuzl8fIjC
H1m6dE81/XZ8vzOVdWIZ1NpqWpclbOj+s3Kf4+SvMe1QOJxwrjOpC2kmQDLyWCkFkk6K+sGgtCla
+Eao3wAJL6UySHnDrK26BS3I6E/7zrdRP9QxxICiOORlOZIR4Tb1ky3zNZws0O8EOEfag6DVyL6t
Hp792uAQpZbODOnYYp+zptKUJk3v7+Gvq62/DzZWK1ukSKwZHFZU0jrCMLwqEA7kZRX1ZuPp4LjR
exJ+fuQESLV7Yn6SoJ66nZBDwypO3poDVXoyKxczzNGDWKA8WPcVxZ6o+B0FFrMrI5sLr+aDm7R/
Ebdwahkl2erC4jI2jy+OvILbbhSw4pKuY5yt3JQt3vjXbb9HDr8/9vCslswQJD/JbaowDZYu1grZ
VwNU+3sXGauDoysk5iIaicLy7JftGHsvQ/ow+vasK77jkTxPGkmBoZZT7haROMHQuu12a8XsoBzH
xAtc+w+Lz1xZ0xd751E/YvXbf9cDJGuBuqI6YWRiXuNdNNh+3j5PuS6TVd8bsgCYhyljdy9uRxk/
rVLS4Ge4Qj0G9FF8iva3CyiBTFFetJVwGQSUA1GEadscPfDrt0Tc6vkEgc7I7t7JDLkafznuM5Sj
NUXyA01O9ieou8yG9c+O1N2kHYAJbvq1WWms7NzYd1BzAvBnPcAkyd5e+6M+9WpUHa2wKOCex+E/
ab/++WaUjRYh8ZAYRzbA5MN0+4SgEP9SrbQ9KtqER4trED8WhXtVHHTFQQNp198KyPxaW9LDpkiI
Me4rZinab4qGkunVxUASTpefIuJ+z0NrcMRbq8/qfdHeB/hvLy0N7TNNzSZVZF4Xt8dRCq30be7h
SYPYZHabNN6XyOiWkmA5B7bVjbOBOaRLVCgSQu4zOheJM5gknNUfFowCm8HdgGVi5Q7gFHzCETyx
1o+TRdSYV1D1laMIEC7nbgtpKI0MMCncIWH1BLgM7o/vi0SfDbZHF0hEhcxvNM4epN7THeiTij0N
A5GUKqSt18tUCwcc/IoNnmJvNfQhq7cEJo91bkAN6tSYwqfgbYBes+lzep9uQKCUm8mqVPPqKq4+
rCPz7TxZSTtn9F6+GJBuhwBT3eros1OOu1C1YFSWLQLXbN081pMlWtBlFrSRHAq46+Pyfo5eyppz
SbrfEDSakocjoA2nIjNTAFxQFiA9BaZa5LiPd1ihOAPI/xr8jznhFU6TWDoITvLestuj41zVEA+p
u5N+C/Xb0PVBJb3tbhCCIiesLu3NCBlkSWufzlFHhkfwXRtKkNsRFq+KrIXNr0FZEP9z0Iqtpkwo
lWfOn50nNXCoB44j/W+ELKrB00ijZifkb7DiZpo3Nf83lwDwcTv3dDg0t1osWnIAlOlb/8FlO8x9
cpvKX/qtDXiWmgsmzWJ2itOeox3gx2Cm+P6J2KIB0ezYsTRY+mpvXUnVISeMgaI2fnlTgoaZKjG7
pB0KZTn9ijr6zI41OhTkaLJfMnLk/xijIoFxtK2HLCrY+Hb1gOZgP67z8HcgjLdKAiiCOA/xd9we
7BeM7R3Vv1WDzo+mMb5lEh73yUPycltfkwV5HQXxE3b9Cchi015o9tIw/LKNzVagEH7hNfzG9tbD
T1Lm/UU527VC8mhYj0zlKkdM6jiPzTPvc5urjWgfgBweYphgFxE6fK2HrGqb7nMePHbh/syog1li
UQts3T1TKtl4ahB3y/zpbnoKuLYT1NgyXjge8UeWu1sYG8AWsc0/nqxlzji2q2t4G2qwccJJujia
bg==
`protect end_protected
