`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17056)
`protect data_block
tL7ZEiOlPGhz+v/WYlxHkujvvgQMeMx8y4hV5LZ9LTNnkF5SMUvP7HusQ3JndZDKUXoUoyFfpGbm
vpl4XMkuo+omA9XN+z11BgEbGCZcPmiff/4UkF+pOsyP0KcldVlGyAv++3TZ6i7u1wabR+jp4EYm
nZQpwkHy2zP4t6Z8LVnrjASzqS5ZKGvqm7Ee1zk/81NsWR1bwhSiNsd7FsK1xFA4S5BYY2ZbQw2f
WyIgt+VuHyvIARW3VKTxfuplX3Sb+FYdMvgZSoAmBdLrnIANiv8NbqTt1j6o2h+VDwFomm0OaXIU
Gi3coR9MmR0KMDfs/88inJs842R/W1StFZGmc2bgzaHiTuHnZHmsEqbwdGZniRQyvFfGdpk7o89A
RaRIeRKM7u5/iLnCpyOw1Tlx0C81gxCkNnMA4zH80GRHXv6J6xy1DPrMZGd+wMm105wywpIX/BC1
RYDIC2UdqY+Ei2WpJWblG5soG1TULNbb+kjE1+WoPpSEngBKWb8v6WLMRaDcW4ZfXCQJRWSNykcs
bPCztGgfq9lFXEN9+EMlwXfh7ilPpfOYV+z7R9Maw1pWWAtgzJmGXaqq1xufV6/LawTkqDLNPZM5
qLnTPmm7E744hErIpfJb03qnN1K3oKdjJgPn+0SatHBW2dLITR1PH47f+i+2rlRmlkCqidCg2xu4
DMIWsGinrDd874oEKZ7l9pvb/7dSa7y5rG/bXfRfabdjrBuNzrkVnUxHH/H+VnAJXXVuL0GP8vch
Yhw+GUJWGGYI1xE7BO+WaWN3l+2YGUd5pphkf0Fy48r8+IauGLaR28xkAUUV5bpG0BT+5Xp6D5eu
b3U487FH+gZhUzuemb9QurKJippNgpcliE4IwqDdNTvQbGJUDQb4bEzx/3d8aPTaxYzfLHdrun9x
1GRN1yxTw7DwLzsnj/mrWM4B80lnQdAuAGRtRXu8KaIanOzOya9TjCBzA+hDOvfBGAJTjx8dlR8x
9D5LZCmAH5zYYJGMcamXNrw1e9v75c3PvjuZ6OCKm23xnR2iOy3k5gOCfV0IPSv9fLL+vz7a/xGk
UN+jDmzsltQ17cihC/90Otzzs2Fi0YD87aColjqYjcviiC6f6orwXVLTfV0nU516NurNdIW99bOT
ySZK2521Ozq0JI31f7UuLF3uBOV/za8RdU/zY7yOyD5V9b7RLZPksrh3afFOmprvvuD5jZ2Q9+oE
gALVXUT0i1+MlfUZ+oIfXgGE8Nznz7ejFC++Iqchm5Py0gu1WqdPaJFx/CHgNgDb1gTxzE/d7kuC
dSxTeVF1Ffi5CVyuoptEON2/AeCHuCPDeKUBcjro3eOMtDh3uvjkurOLGQRLQQ8siFxjfuTxVHKS
3iGG3HsbghKznfqBggYBr63/NdGiIsmtTl2h/APKLTPuuS8GYtvFv3mXz8T78vK2GTae/fBvbKrK
lek/XX/KobcrazYLc90q+HkUmpNvjNK/GY2xagJ61+TJJBrwKE++wE/QiZ7axR6WaTeoi9fcnUVV
YHiVkLI0garX95Xxsp5KN4qFwDko7s+jK6X502zaZFcefVencLKdkv+rKbUHd8TVoaI0rt73zChJ
M1SkASWWdwyt8xbGGoUk+a56VJJ7CQNkcCQl95Kr5fxy4s/wdvxtbj5guoywqfk2bfi1rttcMcll
RlJrcYOznfITLnS0sgsRV+cfbh8DO/kAAyMGNXUlGWPpEAAUHfNxkOHxNysUfXGV6dPPudBrdzUw
I8yJzuv+iNfADR+SkeOKRscvbeywVRWkEK6B5JU3Sk6gNHY4Zujq1WVkWs5z1vTeI/aiRI2qTFND
Znaih/UUPzN6Xsjr8cQisgRzLVsCoX1tk1I/Xyu4y0exJKwBap8M08ANvfPqkiky4wEaJwMhhEbf
HJSGo1S32qRAtAQA86x4U7OMtUwAFFRgy0LMwPdWsq4E7EJusqUY5TaAESEufM5vWgt1FeM3d6tT
H7TUmI5+Yq5jVIMce6haFGTcUOkZcXveiXmMOhZHTaTbceQgsVEFb3I2Vowx6ZY85E3+xkXotI36
YGlkIUxzGuGgKs/zbdl1FRb9uxBNYW/Z8cvdAxXgYKUPMyHuRRP7sAVlRg5zL+d8oFBFLhUHUj+1
tALPm5y4D9EQmuxP76NeTm/wxAP6x8pn6InS9G/pmqxaoHhBwCYxBgOzAoaBCm/r+WWktHp7rImZ
vzVI2e4G5lB0Qu7WDVnLd9F6DvdSaxOiW685LMJ0NSJQ0YstxjQRP/fXWu3/mcCm+FXhjl2nud9b
+xnvwVwJ3CpmHkdnjSv9IWCOkc/DhhPXoKenuEMCMHVBsXpPpVwhOHwkjAp6932F3CQifMPsNuT8
M8GicXmBVKRaDfaej4KJZpigboMIW4H27FTkLI6BdXoB/afXzOrnV0RiaZUwMnSXeOaQSfwZfw+2
kubRsd4E6b2ikFaVeLxwiFV+9xRd5INXDn+SLeghxCnTv8M4Qew1Fjv0ModSdGIW9BfTpGBgR7I0
QTVYq6u4Qozf4J9ioPm5qGFWqBs6YUkfZ8+XhW8JJA6yjFzF5k1Xt2gYSC4DIauLhzvKR8MbrGdX
fdqPgdE1SZLzj5J+pBtQpdB7GfYkoKE7AbZdACEdGD26jbY7DQ8DJjQgaoWp5cf/zw2Q/s5cqs5N
oEb1UDSCMcKIfaI/3CA8Uk33MEZpjRicRRF2h2sRvp0qUmqcCKr0w8JFPaXiDddcCgxKq1Fh7krh
w1gRMO95+ejw+2nGJIUtqkElSBIJR9T2R2pHAGU8aRJq63kw9pUiqeADLDtUq2ibfNwSzFORNsBY
ATX2eETASW9Sq1DxGCeEmK8YduDPTcNAMYNg8jp7e+k1Uixhf8DdtsQzuEugo/UDi069B8hT6T/I
zYFERztgyH/I0ABCWl49CE/kiVE5hoRojvVTmJZx0mSErBirghYrsnLMAkqlvkIbNnNDbjx9Wp24
5SV9jGhsULfXtCcHorzMyNMn7Cu1hSg55gNjgguvPOmo7i4r1TlB4gDIuHwPo2crsc/F+/SH9nyG
A81jcL0hyxct5DENRTXpyArhz3P366wAiUmfvCyvueyuLP4elkIesN7qW8Clx1suqAjHJPYMy4mj
JDmi6/5eu3JDXMFWubLOXOLLuUrjE0ibKfM+/R2gUPm5c5kIID78YXgtb4Itu8ZCXOmEzGeKh9Lo
cIzSvATzmfahc+jJbzkupv43MR5wX5nVteQd/zsTlg5i1a9Tu74QF2ytMDQxuhOGbrezpHr1az70
/DnLMIEV1niYJLdfjKYgHI2JtLagAZ4hIIdj+k5SD6NOCITY91KSblsEaeAJ75JS44LD5pF+4v34
2q9xjWr0xzQm3wtPBT3zXRTFmSvoqYqmcu7rsxOxStt+Ww8u+bmQCZ41sBlIbfXJy5Eyd7ZIognD
4OgzGBohXrG9QYEdhQiMJ4t1twVZpAUrLmPMUJ2x0htxzpzyPYon37l4qoL3l4y5H3JM76yUQHsi
J2ZwuAyNqMyjnktd3IEMLA5ZNJetuP9ETGdaKF/GLcBGYwvBIqfM74hd8/GgKNsLLk7vVVABEDGj
476gRsfsPWqqwVDL8fYg2y15c0y7tXhUZ60dIhwXw5WuIDOJ36yRJSZKqP63QSotrk/ossVioxN5
g51JZERCQ38Zyl+WagvgRcXPBTNhxSXeymiRYJ2DrBnUMvUw+GtunsemnugDJ+crKbS+eu1qlePB
/dvOSeYn/hplsfsuHboENm013pfypW9HCr/LXKECPuh73zmbsEoLtyOos+uhOkUASkaGpL83Z//t
a78i+KsXa3+Q6HJ5oKCsIclBp7ehBko3dPy8RcCe6/ju3ZNsLkL0FIyLtzviszYABgXfFi+Xq82x
z0eps85osJpHiKXws5ctMke2uZqkT80p+iRJlipyHFq/Ay+kN4HFXQivonwdInMMRKpypijNBqYH
onh09+QfYcDGl9WSKvpfPVP2aAKhRnhC2BgVhAy4+3x1JyRXBymSu5yRN817uOfa5tbDYmsfLCRZ
zgtNOBsflHGOVXIE+S6uSV2c7GYx+yKgFwimI3C2HBbh5lklykOk74WQeLIfahOFiZTS+3aRFmS2
stCNlLEjsI+CUuQDhmzeC9u508fo/+fr1IIRzJK76lf7jMEPD0kwWde0kAmTp8FsQNaIAHYwQYCz
BArK7++1XHzXtPOMz+/0Vfxfy58O9iY98jKHwjSLlcZP87pddtWk3iX8vXdc0LoXNzBC5uwOKyQ6
zNqlUqx2yzf77fgtVsKYE/3TKI3xkjZuzYE07zqAl58k8E4VRS+4lw9IgZKcqv40Oau5Z68OLNwH
hQDACPYbv9CKz3+5aiA+MHDbPnG2C+n1N+9l7KU/6s2bDEbJ+SMJ4RexVxC0znLGOc7XIv95rnDG
MJvMBMGmvEuT4HvMLvKoVb9xIGlzmOGr23zNW5VaXiLDM3m67nkQr+COpZLis0FfGMKxnU62F6i3
Qh3VivdIbYYfuivtUVGF7KNkDgdF0tuLAwUQCMIZuLD3X1nsJj/w+UAcDYUE7GuZwOhKg5OQvELL
c3lPD9tFbhdCl0v1V41O4NDfudjBxuj6GvN4HmSkPjvtiO0RA+OVywMGGwxobPpEClhZgUT8ddrP
LDCAC44aoojhfpCY/fdJPJ2AFmLzUsaPpGdPvB0B5W8RNFUHzQCRQ8srlypxZt27imrK80ho2ff2
7FYTPJUGwrIAYW0m5SWUWiaLvvnDWAZH2A983lETKXAE/UehySgdYvV/GUQCx4pU4mhPo9Tp/iJi
/JGwpAqleCrJnlvxxJMWeWIQd7o9iSaSIan8wydR6nLK9eTBhKARQ0U4L2NjYiiqpQMnie75TMjS
tiT9mvnha3NFP7QhuaKJRL9c17rcDErJaIBcn8pmfmtpKK23XjEr0iR7gP0XXBwGF1mbGKAWVPgF
AGHPjsoyM8HhN2ANG7vulxZ8TK+1UGj8qGbNlsOxyddqj/egJScFG3TpCdOUmVRYtqifalWKeYqU
0j07K42RwvoR3KcTC5132d2DyrVP01PwdttHQggq4PlWR0jarrqpDJ5QU1EEUhbbRKlgLZXmslOG
8dMRQXEq8qvd7bHhIAiWpGUqRPdOeG4ZehZqy7897sO6dMDmP6FGCxDmhX9TYa6QrKUIgqkBCw3I
1Y7H7KKlwAk5HGbOfTGqDRWpdN9J20ExMAwC6V4dZ+MY2RwjsdZJIYcedg4nfSb+E0+9BEpQFImq
gf60tBkjoA4tLUpkfJHxvOuRyXCqH3XaU1Pr88KU7EJVoHb0Gj4IVt9Q9x2g15qoWP8GiJHrX7mo
CGdWNa3hKfjlunfXCiX4UflwQu1OWJETu/l8Fu7kyjqr309nrykEr6QsnGtxuDyUXq52nRNMYcqg
rBko+moWBHG7frSb6XRf9mhvnMclDE0XcNjcuTSOeuKrTs5tpcKk1rrW8izwBVjRQlBN2b5eEjXs
/+f9+te7Wo6xRqM/wXSQl/JVA15oTkOoCEMqP1xcjXn+22K2OQJG03pbSJEKiuPnQtzXUWfjfMMn
gVkrtDVzpyueZTNUwvVht1ySdZ3vswTcFSnUuuscvzGiwBgLjZBdADIy5BPPIZ3C0g6c/r86UfPI
kFdxF18E5oyAqKrf0ObrWcE16YJS1jOUoz3/0hOtL5C2KEPa4JupRxjUoilBXfcsgRZgwNJc1Cne
M2h5Jt2ZS5/qI7r4hmm6FFZPgZDNI3eyOg+97ZyVJ9mMrZviaiZZ/8/y3lZ1Idps5LS47dweQ9N/
zmpG+ULAFmuFvMLszZHi97PofWHbYTlzi89uojtraxcv5bufhch1OohzQBwnFU9cWWO2J/YmG+qG
CffA/Di8DT+mpY67qTscoxbgnpWOjD325/nW0XGNeI+f4CAS/jD634fuwxSARHuaPhir1mHlyp+K
l2af/c0Sna9J57u/tvoxM+aTPs1xsobJwrnLFfNfQNKAkF8hqcuqa6tDb3xAcNkOI4os4xqbxvyv
mFVKit7xGMKvR9T+12wSvakrvNu02BTpt9GVHGbSLnGZYhThoRVE5hOhMgmlCEFo/gJ/Om9dpeYg
6RzC2p8V95rzroDYv4/QCniJhVLM+NJ4v3+cvh2nFkUcM3wkuoyQa84l/RbX41SBMgk7SuAe9zs+
W2vPvRUdCjCyeDiJkNl/0VTiLBjpebQDLFuRJpvOXBUZaYJLHSl+4geHi9SXtgovbzbt5V0V7xCK
fe5Bm7BytrZiOXe1fncK3tQcfSJFcPUGzgaKGBfYOwIciuC7uNXttfMSGt0z6/EoB+CT9H/kr2dc
F4EdWFJQFGE20bz3t8AsatL5UDT27kdxqwliE2dGBMPEi/vE9teqJLYjqkmf6mbv2mvvNH78zUE9
IjoK46v3TiLb57gh90gvRRrP0oMdNk1IoeXiwX9nxXhkhC3SHLZHj79ZhP63/3Mr6xNDTCh4tWpf
lcH/ybZQaEg1OoZpo2QlsMG/IrjNAPxeE1wckTyBBgJLNuqkEcU4YidmaZH6lmdKXb7ksZ3StqXa
ZcOm89iF9cy7UeqY2EOe/Svpx3dJJRwuUzxaVmgmwjEwBSLkJ+mx7phNHRVrcXwpVUAGl41JyEyl
P1BX180LPocXzUmzarRbGXQNiAcJj2CVFwbWReMVecesL+fdIjF5RgFMb+bxEmdF+ogsY3GiU9Rk
ah6iHtDNRIg8lOTocj+Dp2VXfUXYX9LhyBTNeRTPAfiWCpd10bHsPuyBlgtNIKDo/rGK98HKFnKE
48vxxbZtpB5O7jx2G0Zjh1PUQ7TtF9FsQty0xaQJ91x+8LZvOMeT2RWI6i71RDvJRM11vXZQUXgy
feayu59aNqlk/QLMVBzJ8I2PwURcc/OhkNRRjR9H4fbrIA2HZWRLlQek4LwCW6iRvhkARmzPc4Em
FeUtr2TAN1/lzvIB3naBB410dBJrCBjva8jj5NHHvrUKvUpyKFlH1g0Wnl3RPPgRUi/exoDngnPk
u8EWPtd9nLhaCv9+TMr4LXKlfjibkuam1TYKpl+jGrWKRD8UTkV7jBfMNNwOkL7WOeYCAvzKdwt4
fSqZFzENqHttE1/Pfdah0HUUNwYnmh6thHchISO37jULLEA3fLjvVywYjFLHSjgspY4GwhIKoMxk
koStbWgo+WcbURmGZAAJIuinLec7zWRMz4JbNoohUWDiai8VA0d7AgyhE2zFw2N0WarBzzYgzdWf
inOLuGJ6axp5pHaspyCEW67rsIcOZ/CmXKElJV1OMZU2SZOOUKJp+EOGMttLy3ebqmAdtABmgFXA
tKgiDmPn0r1XgV1VBYbB1/d7sK+KClp0ZT9LAnPgtXFTsnykgQkY9s1fgo60/BsZJ89F0Qy7s/TG
vmiYFQtbNlbew1w6WqDCEK7fAdLd4W7lpJpn0WS97V9mm93od8yqGgIACxuEyeiBmkvU1DwgpneJ
jngOAE0pqYJgnHy5B5C1f1BUQ6Y6gjDwS2fOgbcfTT2UP7MKP2sO5moHfjogKw9ujdXoZAQ6aPtZ
m41rh5+WaclcwYa9lOfCsB1BBB2OG9GQfbkidNGDwopEc1dF8/JfUOWzHI9PxiXwpQPkgrdjtpGI
i2l+VooVVfCOVG4YSBGLjnDV6ELLLAhomA84wRb76UvrTt/t7O7zCXxxuSMXuIqzyng9DhQcK0lV
C+A+lvCkJw7GNM3smeYMtjnmz8+IPnfLkfJMou78W3paHvhURITWF3wFWX6WISj0JA3fkdAEPH6s
VbztsKzedj7sOrC1kJLwWx0Re1kmq4gCMI3B8T7oaVARybpxhmkpxmacxR2XjAnRl/PzxJHoALiz
0pVTt0eo9KE9q1jA+WX0xZ9LmmscLGMDMo+rfzDhUJU8p4rhdVhosTPXfh3yWnBQlGwhMvFPsChF
DcS5ydCYIKarc8nPLjMCKIF8al8CNODe9d1vfR6ErTrmZDmUzQMWXeDafW6DMlDtwPTGB3jr0DU7
YGyhws7yEivYH/EV0QbzN/R7NyX8RXEECs1kEy2E/K8qd8oPq3jVb43WmEXSzZ9T3Z7cyElcsyGH
UdypHGX9vj/BZcHER8ttA/BXchWTSKNOwXgXK7VjNh6aLN324sAHNeFnyimRoPFQIDmr8h+NGXqp
HiUFn+QLe9VcqJN1FAFTZTxrTIpn6ri0W0af7WKADVdoex+MgGZupJHI/Xpuan6qDLBZN76jXMRh
EwUiEML0uNbvfrsFPKB8pGzRVtpb86P9gqT7d+z4KaU8ZvOOBJyeRlQvZAAC7VZGMmZ041FDh+qr
fP/R5NdNUyOJtPjUQTkLX8gAKNXE/zaYfNY0vlS8uDPt6O8YPgesWkoo9MDCkC20wvKFYi9JjSRV
RnjZ13Fxmt1LfZbgzuZMN2m+wMyPO8eR0DVQ1JIPg7K39FiZhxGNcVVzhnJsXSxdkOCmRZYPpED2
j/hv5P+BwjANU1rOoG63DT8GiEIi8ulsXt5/m1paXi2Luk/v01UrGx7gNUJSqC4RbmukBNa+82SA
LmG/qB20mNvsk47teiWRea4UD5hWacUZPnDZrX7jD24ykkIxR8S3SxOR7E8It2YG3g0jvqyQXivQ
JG99+Hlgu5cTDZ4ZdWdRi0ctumHx3gltkKp+3GUVWzzB32xHAdLXRWl5bvLeo/Rv+exLAHJ7tpv2
dLfNL2Ahl2Dmgq4bvsgzGGtmxqSo1zzso7h2NDfMo59lEloBxvaPbNrwU3UU+q872I8sXNBlzt0t
EQjQGyxMtsR68Y4coPIHlrqd3MDOfmXGRrUj/aV3NZSdNO/vAyQcX0V9Hy4H48GsZNhmBriiy3CC
cKgk19GrUqE2E6Y+y6wWDwAbXkf9YCRpYBF5OnZezoljEtmw593c8Z36cVB99IdUxtJw0BmdfkNS
8DKyiyiqqV3eYWn2wiFD3SAMa23GgZdkKDF6gqSCN6xIvH9DKljg0pinPKNr9/7MOdYHlPA/q0Q5
OyGN6jWa6U3NT4MzhOSM/IrbV60djhib5ItM+E423h+4/64PfzxnItP/XVz3Fa3Si/L9+C3SrhJv
hdfI3wbK/pb5GAVuxUpS7kr/6jgHCWImnIeHcZ3qjDzdH9NerKdUT5TfmHGQxO/uRcCJYN3JxoGh
ZU8oVs2KRUc1/MGn3vVm2mgIBCaxTiHoCswUrA0yVRUp9z816p1GPEWhgE04rC3Z9WnNvtN3jtRA
mVoxY/hlfMfYjOJg1ctaKf+Y31ZET3Rxc7uR2HQkyGu+wOtzu4IHT7yJqZOLXzQVR3K5WVQcsyr0
fFGiwGHazzig1kyegUJcKIuamYCrAj1slUoFbTPRrdRCkk0BbjkWMcKfm+U6Ymh6qIZuOAg7l3Dy
CmWNNBXXluk09838HNZF3ZSup2sD27cgAFLfohppks3XInTKEyIktBjH5w7xaObVzjXCHI4ySwVQ
h2wCdYSIns+YbOw5H9EqkPtyvKYCh/e6/7ICPipLhYACNapc9KJl6wIMpZSghuJ+FTPm06+oHIqA
ixehPs1msWU0BW8SrJ1Zfdh9Ko4NeY811xHs7T936E/UKI59X7DOd68FDVOOm7+B7z8A8gjBTVLy
od6SxITwqcmbhhqWOGdWXh77dIiA1iF5ikTd2Bya3Qv7CAod8/tsycY8cfjkWJN+yueOpdK7C7XS
7kiZQ0b+aqPRQ4bRYTs2jWQaqQz7L12ZPieeIyePlJErX8XJW0B13j/ZBpEKKnVIqLOex/h5C4vj
IVmepeHdJjp7R4SnwEtk+J/8OnXTGbuIYcgJMRy/IazyEwFKWYCD6AOUmDr56A3k0HTHVyZWuwSY
iuEyi7gR8pSzYdFzoaJedjqdxlruhU2M/TOl0XgJ2WmwQb/L2JV7AC+SOvwpcXaFt4hNlvoTyeNl
9rNdz5+214fHAZ2/KRxMEniB61Qpnhhi9SExeWvRevYYG1ev2lmx9mUBCNhq4GiwDp6xSk0//d2v
+UYKP+PMPegAF9xassLOMkZneJG/6KoFMVN42Tpl59E6dfXCZXpHevEQ19COH/pLs64OsPC/Ng27
G0zg4nKY9Tsuy/mpvZEN+GTqs99fomk26tYZsCZZKpLAps+kKmNDaWp6/pju5MTMQsjz9Umga3fC
zjqB1jonqa/LE6XhstacvrI9mzXVpTVWJOaFYc3xDEVGtI2ewtZ4xTBty0COoEWhmHwmjLIPhLPk
cqcmRCTmm+3Ytbd3AWITR01bqKufEQ0gCTtEHI+CTWG9kJUYLxNYpsjRQc9TlcDJYpHqKq0qIgx8
hr2KlLBpxsN8EI+075Trb1RoEdHyTSzxmRxUy70LoRX5Tl3zGKwJdz7OyrEQ/ANy7hdYhTZBnAJL
+ZulbpO4/eb8+IB3Y+uQXTRLpkg8ItUG4Xf5uGlSZtyHc/LfXgfv2cpLouPLCEv29AUztgdW54oW
VMtdP4cYWi/1+cUm1yXZ/B/5z7q2QJ+yeX3TgT0hrCKzdPlQUZEVYA1fz+1kZ0eniSu10sTZy8QF
u/FMdoGCz3l/P1aDWMZxSjERB/b84QLRmshmY8gXR8yW++XIhewM+qWvIXFCoP66YUaSvJEG2vRZ
d38WRg33OwY+4Bp/pkWuASg2sseMsJZ/bw/Ejems5NEtR6lZgsdtVzJEWyzPtlT68Pj8FW3at/p5
JPd1H27FlwFuGWSLT8v7JUOjJZHroi2/Hb3YyYFZhuKkrGLrIuA0ZFX8BzIcdNbUqO+tqJvrV5Eu
bNB8zJY6jYe2WIokbzC1bRrr0+4p8vZ7KNliRMKQLnOyVvhEHuHiFASk0Lo4uCj2AettW1lxGG4w
Hpz3qJOZhfBpWSKZWHyyqFIzV9q6j23neNtkiIu0MnccnIxXkJ4AWr58s3wZk6Fa2COB83H+pGOr
GvG6jKLn0Wwq3TDxpQotNIHhUj6IOGMZkea8jozdvuw5HQBfvLFbdIEpM5QD8Y+mymoiynPD90sL
joAZTx0kv/PhtvMJD0wzHR1gd+CaFcQZUlW7oXtfHxj6qDNpBAZzZypxh8HbWX7KMA6wRdL/lj4G
pbjzmPH0X0nAHpXk1muSlwdtgto+9bF+Jczs/nd8/fOup5diKzwg5AAIC+lCTimRn4kS+aiY8re8
Et7FQ0HnYfxQRwSNLT2bIcqy7RZUxy3M+gL1AqNe0AQs/Hz5giclU9ox6qNNiKG2d0CxgKULS1v/
yQ90ynl1rW9/uY8HKqLydN+kcVpbHjxS0CyFhOuMB9ruNDFKA0zb/QacMrc33Czj0O6BYnogNW5E
Pbur93VKRSlLsLEYnkqhQO6vVKo0SpLv4MA2WTyMJp36Pd5ItSOqBZUyg6iF5y20q4wiTFJNn0Dv
DJ5C0CPmpRXAZ+ylhCmIqQrVCbDkyJCYAopNG1J8MB7vuY8Kid5TEp5l7ZO9nWN+KT7xBdZgBGKK
ue+RhmyBwDeQwtJ9ko4D0URHLf426eP5/QQH34VsurgmKwqGF8u/fppfpUrO1hudBOKrJFjygzGQ
R9VOu9Z2+yE10m1IixdSo3Ub8oUrWcKiA2WFQumQViQEQzZ3J8e9J2FkUho4Rgy0VIw61IPKIpD3
cpCc+n2zUAraszuUg1tyiWStYgaI1ZHzpf6QbcRe+wNxh1LUA38i9DbzyVEcj0zI/DikIevA+gHE
ya1IS+0H9e8J6M0r5Xfvh+fbBGGWhdeFgLht6Xy9+wUwPija/5jTRhBPYXhbwOq5rNCr+GrzL+Dw
FxP/blKWdf1N5S9IVIP+5QhGwI0SZp56y/agWgHexseCcp06bP1y01QVqpIgxsWxp81Oszgw8hKP
Cp49pFOb3jo2piSywbPEBK7NS/DJlwb+PZ7pIUGHrFeDjsvevQox9hknaOsNsDba2V6/djm3ynWZ
j9/etoHJXJP6baybPoI3t60vGVgZ/5/OYCv0eEctXAzIR/OVYmQLB72C3iHfqWiwkdqzoC0+Rbmn
wns56aJfQMsvHQV9rY9d59nk7rnPTRlzjtiUs5OJmqh5Y8QDOxqBrN0q3nhBkj75QnwYUz/wLuCb
gOvjGX5dLjQWDtDjkD/7zGd3nPWdljqK9eknnEnDQp+ObQZERiwVbE+a1MafRV2ehNWIdy2tSJZr
CncklU8L+Z2nWgAUzc0m1K31jLc/ky0Y/HY0DnmMoCZQCLnEcxxnVs9LSPhh1Q50AC+ERLP1XKyD
ckwBeSla0hQMzmiknXLmTdoJolp8BwsmtxzBM522256/AEaW3M2vDDuxTq+rZ4oNfCtD3QGe24L1
YLSkgk3pJXER8qitPW/xKIhvGGcXILI0vYrf9vzZQqORD7W2qbWJe26s/0C318djOux7Lavqo9Lr
zSmAUB8nJ7O/wT0FNCe8iNmfCCJ7u9Rq3KoghgE9PoSfMez8fqRICnGSQ6mndxMerfI4luAjAnta
om4Uv9XrzaytIFHZLOSZ1qlWitL0nOND3YYHwHVDRLsTtbAPAy6lR4nrUvu9vz9YPKwY9+cKK5Lc
/knyAGXxWOlxYMgjMpzmpaZ7DYb2TWwrKtPOO6GVjwFzXZC5WEW7h5LAgihAR3TJgUIDkPcaWsut
hB3kYxx11LM6Ku6TOpYL4bT+g/dkz5tgA6w1vG93fUUZv0CdhPoY/z33DW5m8ZFqh9kfI8cOK5bo
R1Rd2hXWixdBm2NaYfDv0PZyHMiB7LFhxQQ1zDhinq6pw3DWx2N3YT1w7Iae/xOv/2LAGbuWzP+2
f3GdVGQyhgbpFEFXoly/H8JKVvKEKRbdVw5H8RC+ZiHTT+QqQPpxQm0okCEHR6BWX8ulfIC0J2db
mHzoa7qIKBfEoq9BbNrDZOQAMvpSRZ56BzNEVJFOd+lJMM6LB3UtVSVCBIa1tPhB30SCG3Egpukk
vOqxCiZk+vrcCEJpyPYVz3+LXNdKK9AS2GuV3Aiu8FkCY0QKldD4/06XEl6xk1e7x408fBo0GMVe
nK7K8ccHspnS55n5D6guY3Lm4bfjrKsv0n/Y9UuscBT/G31DItmNVzxvsKN340PYX+0aFgPov03p
ODOH6HA4Usb2mawt5z8ZMiOmnijtHehopq8Dx6JXe6WTdHPMfWyhy//jlWfpIR5ftddNsO7ttXRw
daTlj00/4VNrLT7Qep88XNpiWAWicQfAie6EBpEVx0gsxXMbTHjtJqzV2azhTo5Z/BPIkDUSHUwI
QCD/o7dcwTwSmOHP2QvgABLFsyoV9N+6SxI6sBgCdcx3QG4cOzCQeMrUcQY/xG51XfNv/QqotRNn
ZSRigMHuiQ+PUdApS/FjIbMKI22YaV2+o1AbQdDbqRgmZkS0D5xo1H14cSvJ2wOOLpcw1mdYqhTR
GZW8hkgJBSzmQPkTRgA6eAx8HQ0rPKCESqW0KtYFWC3qRua9rh7F5eT0xCsFt/KLEOWVk1qIP2GH
vTw1U+sWDguAQTJsyGhnuKNAXk10nB/Fx6vlXX3nGe5N3IQgYaEM78YyBy2ZsNZV8ixvV7PKLavT
e631UcCv7jtIeQG45+8AE+9MG+piIs7aaxkk9KQgnkVw1jpaU+TAfaT+DUSVZHw2SWOfyXhn30WW
GPGxvPglROJPe0vtZPC6/tyMpFBHqTJGR+6MnfTkE2g0BkQ7GbagIXqtjKoXXBjn/JNZPFmxVgtp
rEj1V0BVlUxbhkTTj6rbhWBuEyi3fWyOV+i5DDBbBOUf2zrrOaYv8HBh2M9rePBH02mNcjqUsJhN
6rCKyLavTdC4BQ6XtUMh2VnD2sCu0ngf9OhrW5rGR4gZx+xqT+0ES65ry05/pUteHcEZFFhnLhG1
B1fOa99S1tmIHRYrMGYaMafyska7tIYu7Yw9aeoLZIDlXQ6iYYJxvV8moCkGrO0B0+2H7geL3WtW
NMSa1I6DwYu7U86J5Sc/N64QvXhvovvOQ4oTgbF+QvJSbRyWWv8gUq2G6rIK6AO4XvYRJIqPPnpX
zrA8aLDAjUJ24+Ztu6tXGwe2G9koHELczb8US/O6CCw4nZB7IjnWSGu5CkjbRcwIzbxa+TsXPXbg
d79IU9kbfeRTyTHEXrFQDGsQoyxlHONcpvjt/7c4woCcOGUX10erX1Efx6ftpOn/yGwR4eRYG/C4
E3+ip0eFcS6Q/MF9E7UwKyXDvYILDGsXSJIzEGhlEbaTtzhXiaGPdpzXe83lATloU5j81YM0u3JT
5vC2rBxdZUeX210kWWyib5M4Z9xN7p4kN0fiyk9ZLmYly0rse5NMTaQuXeCLpe3jQ2CzAAsSMGrm
tCjRowo8S2EiZqfGIMKmqjInB/HEpRADbowYcSTJVL15mpZ69CE9pjXinNnDtKAg6mhwMTKyc46S
Nll1AXsoDD69ib1bPaYEw9fa1OTVOBA2ckCHOWwukDBFZiYK3axf+hy/4Nul4C+PjojeQLFX5D7R
3RTj9SKl1qSAZcmPJ2pFKYw0rNnWiu332OE+LML6jVYEHnAi1DTIrDuVhldLtbMyX/18mlKs/FfA
Ow9DFRnTzHjyMRmcuYF0LrXfBV6xxwbHF9Z1Kn3E704r6kjtdQKSXC/oX4hQkB25AizcVCibsYEZ
ny0vHHBAP7MPBGi6GrXFFs3ipiDo3czrpj9YOIwSoKphMSCYj7kToO+rTEsyVBZq5vYqqH29hhb6
p1ItkLrfQ+vE9nnd9hmYTV8pseBK4XIDw/P3Sw8UrB1jifzSDz25wHd/YxJWHZRx1NueqrzaISQM
bHyKJ2lIu2E8vYbjO1C2VDjYVB/wtWDZ9Vb7CkGDfozeQvwxqwlvSLQ7aFgLpDjhj3HMioPC8n/J
dTgw09NiWjaY8+LeKaJLX4fdthgSjWjP0DqEvCP/Tbehd23o2eS4QP95h9NQbTNiABBXgZMVwlX3
9gNkH7CMHOJsl+DyNycCVx1iYqRJEuMPWiHL0hjVVqdrXoCmTckrlaii2uHeLImxqBxAkVDNZsTP
BCOY0tY1FeZOtRJ/ZgY23tg31vvJiUny/RxgvXWPC5OcVvbOrHGRdHKNP/DtJecb42Q8p7GMVYqW
YLganbpVT3SGvnKM6dyRDHrzxlznuDDWDq7JlLnlhOBRHQzNMtHKKvZb1+WWaG+adwUU5wHmaKzY
unOr+sD120vWcNfJ2Hff7Puk4wClAulQtR0cDJXRqbchyAIcrR58hEwCjAuPnsXj/7ECYuzdHJoO
hMjxjce2OmjMpwj7nBh7k+k/2arQxhDgT4cY9B4Mr3mBDrv7bjyL6ba35x2O2xnnCukOvkBB/7pU
bYKcuLsDSG6WgbnP7QF6+272UVtxOFM+c4zEJ4hEgWSsRvlvJxnXAOiJWhCLZvtvgjh/xLUaV8o2
eyJkkRjk5dXWFOoVXRHJ1V3+ZLcfdYlMajOSRD81NTZa0sQGJRDqXc+o/zHjJX+ipXwKSl9dHYcE
k4hC2YOTvh9ayTqItsEWoa/wGwqPNFnG93/F2Q9rmX/TQZQzFaoV/MxDmlDVD12RZMQZHoPNQAov
YnQl3kkWYU78uiR/N/7rDa0bKqU2yivEvAuDzs7koM1evvy0TQmJYN/sXOrf1yl8ATV8nv5EKJKT
AayYsymQ1uv6fzSbe3S4zp47A8zazfRZRFttfpXqP0eFtHe+gKMIYzRDXV1H+PvVzBaeHgrLJLby
3tD/YaoZLyGJziYYh0zYSDz2bTKEbAskBmIDN+jjbFOggjAiYqcsvvcSEpPHm3O/Ipipje5RwMVc
nEoWhp1dYN4g2yf4lRyOmoY+yTNNjQVZKIiY9B0iMO+EaMA1s/KDRNWWxV/OqKB5t3Uo0nStn4Mw
Mtwr7yCZ9esJv0VGqXFCBmzzUHDpUvIFGle6OK+vuY1z7I3OcuZP91/DYmiB2ZGwJX/dTafngmn5
UatE4IfMwfWRjn8VaYYtBEe0CS69GUY7nSVyBaN5wNtCQS4CiU36t41xAK5QauR9OQKVjpAeNmVA
zsGoo3GZnEfLNjnl1DurNVSdErLhzCX5n6PuMIWjv+O4OKsEY8xcVk7t12xxRhUHxCpNVKpZ7Phh
OpS5Bb+C/k0Rd6yLrh8ZknuVLvkEUg9YOV5WgsSwuKs5bFLu+kLgeUuBKouYTWIGy66NSXefVX4T
lQBBgb5PiWgcd3vZ10hdKaQKewb8MvqqR+RIINWbncB4+oxOFx2k9UncpBBejylLXPaPdTrixhRK
aeNXxkDg6rfi9ePZHYVcTqO6oowL+jS7Cwto7miFo8pjr5fodYq0cgS0fYKSbLN0Rhqgf8iBf4M+
5+j+oGofiUWcdDXcvJQDK/Dku/y2fMYE8Rq8CXSM6x37sbdJrKsFRL6axA9i8EaVmczV4VH9skaD
I0xYoVpAGJ9xyvrJ9xRXrlvqO0vQj5EdVj4M4SDsQhF7k5FLCgLhoy35FVIARplXmS1M9w21nHIp
JJFJk4VJQJUQAMn6rDqVAY/OZS081Jk2zizvvfaxDuhNsXDsF67DYKUvxdh+6TGb4ryW+1L4jGk0
NO/g15bv44+T92KBcFND3wCik43R63pIgx6vpExIU0XfSeU7/RFdjq2rRQU4OK2DPfZiHvH1zVEc
3uBEE/5NSJywidgIOt8qdQ45E4NT60rRRRJWlwoOWqrD6hrn6XDVWobUZ+euGRtw4ClD7xb30iG8
AEKMehBwaHOf+X0igN/gfSIzggbL2gwpMGHgnqUSjZXmn5EDhF1S2Lnt263MOl10+c7QGn7ABtW9
k8BmIKyY1ICOJ0nXDj75P1OAVvqEKuwUl2Rm1Kt5dfoPeEGmJT9TEvZEk4qv8MO1StpZpKeuh4Hk
sqkHGxJpeb+O3jT2Y5NK76Qyh9JGObhbd9gNpHOgFSH7pBCQZ2JHRsAzCOhOayj2FXeMEqZXkQSF
KI9oPzFgY3OYhjpZRAQb0AcAtvrW21a29HsiUTcCIBb8IcZomwdvT561ed2Qd/7+lgSel/WbMVZa
PY7FlVCtrgLJ+Wt8x7zhOT0DC/fuAIFwxA0G+Ent/Y6/ME1iCOxJk3JDiWB+j8bEexvJNdvyF3fU
ZMT4BSkp9mn2xViWLgGAewM410TNtPMef0AfnmsPqMDVM/0ICyzv5paNEXFR61hXEzgrm7uTNk4g
wS4MARF1cZuM5HdeSeEZx4SHxnsu1D8DzBC+GP4uZDBPrUnSvfvp4q8EGCsVowMusgk2Y8CLomq1
5umaY5xEJuAxYo1ta6xjCzvh2JzACaWK2yFJmyvHw68rCNsP1fXOE5uGNuqgGArdIUEmtWruwJ/f
9D3HNxn3lCiAd5vfJ6+q6p9hcsnqDxR1VpTqNOQ9SG9D8fisykBowYrHEh7BBfpIxgW7NR5wWT+R
B5GaqJIz7iXomTIsHGspsTSJ7b1lV8lSugLZUtmZfldBdupHhPsJc1Xevdyw2P5jH4FJko4gr9SX
XAyndH59KtTM2NEqfdz5fpSFzu3yEjJMHHeoAxCzTI+JouUlUpv/SGp7HAJQy9hS6JdVO8HHe7Oe
2NyCeFYQH3PTnTXnZpeQu3LTAwuhb+JlPdiR9GhbLso29r8IEHImV+XQsbAV7Ub8yfLNXtcrbyVw
UXS4hPTg4GQXyeE90BqUlTWSVxL8jOmwMw/3LtnPvP6W9Xq/nRHi9Iw8R4XIcTp12jk7uYKbBv2J
JR1YE5GIApzhlTsrGYTUvR/beizcEMiz80hnFG5rRFOkQuwPgosHzHRdxAZxwzL+ilK4d5RfPnxK
sDeppZE9szOqojSdv6QYeoEQ8yrAFZmL3R+kMSzc1DuNq4MjVh5nRXsJsLf243rr4gre5TEzgn1Y
Ji+pcrEKgtv3dwiLfMF5qp2wijO7oQQzGkOvrZUq85BA00dQLvj3hHwOdNXqaopS6WANAcxeayx2
u29DbB/DpbhOyVUhSr9knwo7pAjjdcsFaI/GXKGLKh0TgXNvrYeez/uhR6uNlOWOGfXXBgCx5eIf
XQM6ifudauWvcdcOrj37Ym4V3hNY/ESBYJpj73bIuLsu8lxY97lyeaiPuN+rDmvjPNrAdFFeb60V
U6bfCQJhPTL7MljZ2jZUQjzf041tpP8Lz+4a+fnHgYmKNCS0IZNWYtfCap21L1a7HxQAt55a602g
9xPBTU0AidW+h7Qcos0wCuzFfGEKcNnPZmMt+oWFyqxAHP76ShYkebWUj64RzXxCRKUcsEZy/1t2
D2R5q3biec43zWRXxqwJdK2R54SgoICsy102YY1OGIVKhqLsby12pHNx9dPBSXYwJICnuvoNEw4I
EvAuHV8chSwMMBhtFyfzR2wtctv30xcl/7lkzQp+16gS/LSQuqCG0BsXEqYTQi/vLmRim38W4boe
xRUycV7gDVsPPSAeFRrWMM0FxJW+AulRI7Qyz0QPjzcapOzfI6FKnS2TZg+oLfIuduq8uhSka4ph
pLaz63NQuvuJ5EzWDupsg8TuqO8/AG1LsBfWLGH3/U1zXq85WwKZ0RR9LAJO+qH/QdxwzBa3Yfor
TUb+EdohaCK0gn/5r7NjSyXZUjKR6PCqPHhITZnxbCMNOxeBJZKJKVUQXVlN0g1lXOkWYfADgs9U
+JW7BYoQjY5c3sJLF0omRR93jKuIsqTLGo9HWD6vQx4xpYKQwZAV1RWozkzr3oD3mINSo67LwLe6
xG6wrl9OzVeRqk6GiQHWBBFMQaUX8i25IkLpWf02JYw7xu+laOj86ge6MaZnL5L94aMco8yTgMeS
DX65cAbIDtKfj2q9CE/AyiHQpyD/9o/vi3BJhlGxS0RA4aheD/Ao6/HfG737goIaO7xQkabrWESV
q1mcMg37K5vfBBz8Ltn5ILkRSw8FM+9xthZ0wBbPCUeRNmVqHQTplzEBD/Yg8F+Wd0OL64ZBSgtj
C0xcbPMsjA9MPyzmZL4TfmJad3OUHmrruU6IMVPLm7P0y3EFsLGtLeARakDLN2k+vi0MTwxIgpXw
HqhNdd/WlidHleLTc1xC3pa3NP9r1sIs8UF56KUBegbro+Q1m1KeO/heao/o+ysROXiw4i/teTQh
UHlWdw4drquLFqMRxbX1lKXyUrxvxF6SzBMaTaohRVeSuzhUvWBQwOIX9XzVCqh/+27LORIA8CEB
coEBnUgu0ymYicSiNj5bIbPle1p+6r2oeLyxcS2ntiLYkM9KPoh44NYQ6Rdm4tOEEK6KrlC6tNJF
NE4ezfxhAAFh0zLL9+ie90k2BTmmqS6h0xTNwtwelzozpFphj8+ONvIms0dHby/cItUNlHnTUCoj
p82nTBuJ/6NDzqLu1O6nnKWiuPU7AfVvsezXJOHtzL1B92Pwll3d2lvlPCHlrCdTDhew5gz+yosc
QGjVgmEqXZlasuJJ15/D8OV4ndsNovcxWUFi+zy6zlFjjwimV7edGiyjXxdHWwoj8aKWOAyyjUtq
rsXJ9V5GQv7++6ieQjU3zkuwr5b3txjQ4fTGF3MWRVRmeJngAkIxgU50zKbPoEJjMUny8bD/YpLz
y6gbHVnOcxIl/Y5ljXKkf2x0jtZ2pE33XfYVHobaiKHs2gDRHor/JGdPbWyRgeV+bvRYjiqtLhzd
cPhzKpL9x2uSMnu6jpl/aQLC6Z37FD5X/rNmn5ZhamBg36fRgA25wK992HCq04omc0L1o7KVhQBZ
XuL/0QHAkxUUp70WuQAHlRDLWDKOcz0wUDvXtLETsy/S7gp81jwRQXnl1s8FMXx4YKWYasg8fZqY
4Feuam/eJ6ylg37HgkucU2/d6hqZXyYm24vcXDNQkFWA9dEIeFNY+j7cyuciLgS4n/cpVymNzykh
RnKwTgIkfXC+tl6gzMTYs63AMlY2tZnQTIgsJXYZmp2rzn/ZPDlF+X04CEIyoKFaGfi7P8ePTlrF
vkeoynn/e+BfbHiRtnkLy34AYoF43FU+z4Tm/igOXh4QRO3JG7IYWukqy8x6/9Hb+g8oXu661o6C
OGIJQajq4ohe7bMrvmyqEKexRquAd3KcdRh4gyYU7YKIY4YMV4odgk44cXr0ccNAO7JnesPaibcB
PcR50HrHXRmKEvt/KvLwDZYM0EmQ6pgWKLU9onAVFYVkeJEImLgOXSVjmrp3c/ANV24foFYgKNIf
HcEw76JX1Cn8edYeOvhNdK+ee04E64EnlioFtESvlejXmpLM/FAmU6PUH5u325U9ZEuUOzgFcQjt
02qJiGB8n4fVz75ASJBZVLW+vlP8lOXnRsBUxhIIdPGEaC9TaNedUGvx1Hfre3is+/C7l/pb9XWy
chXKQsnrPm9frgWNNyeDYlnAEw2REUqSNOAs5kvqzgTQkJPcqTevKSBUXHNk7OspVa2vKG6Nrnb3
FPCz3r4VNxpsV12QHk1GcTf6bZOENEG+xQmxVGakjTZfjSRo49er63gflnQdaq7H49NlPT4nUFFq
1yRGr7U0jxBjR6745F7YO7i79W2FFug82Z0xfmOpNqsIc+KIiyoxiz4PszhWjTIvJyqVpNzChwN2
X+myT9CVZ0C5qjS1f9Iejyo5Ihg/prGK8v40zmbHc8EZ3lGLzdUCONK7PllM3tG8lAYcU+x0SWq0
Mn3aMLjjCqioIdVDJvsIhA53M8NT1WzoN7MYI0+01oXTwbc2/iV15xvHPZK4vZedl7XniFSWbxQ1
5gYCoExJ/YYjmL5NnHHXg8hKJQJGNowhEbW+lIQKrPBJ27GsotRteX2bwmHZzRws+RrvJt1aYgiN
v7QtqCUgtgZ/+lQW8orZF5f6XfJO/u3vkZM/DVoya+RH0T8K5JhRWvpznAlpjJj6sdvZfQnilS2W
p2vi+OsrXvTKUKNxpvdHs/lWqmDyh2UV5PCniwVG6OAibDGlvxFK7422iYigboVey9pQmFb8J2X1
z6nJi7l3Qc4XsTeyk9oEFO9TSHngaHwuMIE9C1u8G/i6Ivgnn6yAUnptBnRW1ZhIk8MusZJFSRDo
CMt8Oppv1F4BnN9e7rvZrqOc0lN23gdH6KpkMUnn1O3j1usycblEk4cvBKPQKRlOdxAfZqYoW4Cm
nDtcddkFVGoBqnsvNw53pIY/Zy5CK5F2n5oL5YlEjCGghqHMhZKVOBlbcfd2up5543+hGplrlNtn
7bixemVnxNMVCCaZyFzVeUEwan/TwfJ8nTpxck+P7gW9V6Yfo0naDaVsWszGS+7joL40dgUs2Ik+
40ukYeh1nfyzOLa9nJhfn94fZymg4LIO6DwLVYzlIs3S6oSj5FZFmAINNtJpJuFZzAGcFCog9Wvs
KNe8hjimrcxwAaLVo59TiPkSj7W7hyN0UnjKQMgETBqOyAxeAVz4gkoyIaTBl5pyPU0/ctfXY/K4
u73LKSYfJ+45uwQzG3TH/0l1VGcHqqJzgfsdC/oYotNvCw0WpJjTry0EfavUNuouE4OiUtmmmRM2
DIG2T0T46utq59wM6hqSWU+LTwXNX9t1m/8+6gvalJrPB2fR1MJVWjcunhWbz9wOU1Dz6wDGl1vd
qX+LF6jdvpn73B/nmm+fsIKORzhUo9snXrt0KjFMSYVjxlXwr7Qc8AlFVhWl1vGSXaHoKr2k97CY
hXXMdtz1xeYFWen1IRb5KFNW0NQ/77aF+nqsS385RTdkIqD3BUJj79Q0tc8ACoo+uw9HFbGjwCjM
9FxrgeD0XlEwdIEeoXhk6HCbLay5zKldSpwu8mrg8+zlXKuLoF3AYWPmaFGifh7g8Wlnt5XA/ntI
E3c2Nwel4Wd4E7n6z0A7EKi+8MY8gZwVxidASN9AjcHeOc1Ir49qvAYpWnPrCgtdkcYwaclkGzIH
sZ3Ex9H/L+v5zqQJgCi4s9FhmACTbn9RZMnkcbvcjygFiI3qlYR4+jxs+8FgUU2VFwmAiNHTo4YS
6ClrAY5Nz5IAElXBe+ictHSkep0VxrKfXrx+9V80iITZI4Y0/8lHsJFdekuF8dxb78Pa6LVeC5xP
PvFk5PVtd9OFHApI/iRvHKVBHmj5cJ6hKcVQ6XS3MBDTGSd8ZWsC2AYAuknd2zmBM4LS2h5V+olv
yO6y0sXo/4z1P474rdB9IYBG1i/mk7gfgD2D/z9vvgyO7gyz534lynbR4+jo1xODj985sh5Bpdfp
yWtCapNIJzZ2TXAr41jwsuNxRJRJTF7mWLpd2Kkc2J2PO8moNTpRkjOy5kQxLfORgOOXyefMEylx
IFxF7a6yyP3/tv896Flnpx2KOl2GMO1sFub+r7fsztdQe2BEShUuLn32st/EsrCZ/bwqDPr8FC9V
9DRM2jkvEKCC/kcW+vfArvqBlSZUlw6gdhatjdrVIM1Cxeopar5Z+s0iUPtZ/yI2i2w8ZV+K+hii
dwZLz0INre4jeTIfNYS6vRIo7+TylAkLXD9/nvNlfFPIktpuQcFnIsoKm+0gyQdx2d7uoMTx3hRE
ZW/v3HiWMagnv2em3TNP16586fqu24VEJJDbKY8v5JAYW54E1ZO4F/R9AECBklRxStQieA+bJiKq
NQycIyC//Y76ShX5L3Ndkb++vWKGZB1Y862hVhNaOYhWlhsw7A5mKFLJPp5pyEqzXiAYZu0d9tBk
F2xUSmzj4E7WfARii/RwVbQycJCz0LgHwtlTsUHoWSZIGj9jVgW3oVttdy1ICfKw/BYT6vkeZQbn
35ax/sovLNNj/n5nfhA5USv6REEcZjQVwhoh8YcjSlJ+g/4RPHISJz1dDMFFtrUzfWT+uBpCGJB3
M5+wZ69LkyHxUm3qcg8rp+ceQWAL9kbUglYD3UT8RzUpYM2Dz2F5wFHxWim59X9DQEndBltNYFwJ
E7EXWDdYK1Y8mVPtmN4B7adJrncVDuXlQ8Mj3vIiZhLabJgRkjLk1L27VopvOTELAOOrOdC6LhEC
pE9enmM/G40f+osrMQ==
`protect end_protected
