XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����?���H��7|�d�}��PY��+V
������C͋�̽�]�X�ut MB�÷䭿�p��t�m]��'j�Y�]���L_pR�c5 ��a(�+�j�QVm�Ў��q���_P�ud�=�XG������7z��y���!��֌�L;��)�b���ܑ�z���+-k��s�VS�^�\�a�����2�i�-�+�����-!�[�5��]ϸ{6�x��yP{D��]�^�ޔ���\,���:/�,�
��mi�B=���M��F��7�2�~��^����3f���ql><q�u����4�s�q<)G�noɅ�Q�O��e�D�9���@����1^��6�a��m�=�K�M��]�G�� � ���a���� ��R���<4r4�w���qӿv�$�Rzᛆ^?�h��hڬ8�	�j���B��t�q��oI Fq\�o$�H<vܸ��� �1ƒ���H�S{x���$Z�+ю�rg�n�9vҋչdU��4��@u\"������>�dI�T�QJ�z}��vC�e���+r0�p�|�_t�Z���F�Lڈ$�
#���C��+=�����'ZH��)H���l���!�s��z>g�(�E(�93ohw3x,���F9�,}B�$4@�O.PM��1�S�&@D�ˡ3���	��=�ӈ�(��M�Z�@��ș���<^��d�KCU�[�.ċ5Y�;��e��.ml��Բ%ȴ����áZ��w_�pYA���$���w�z�*n��XlxVHYEB     400     1e0�F`�<鑃9F��Xo��uz^�Ȭ�:
�$fM���H\@Gٮ 2�T�	�-����-��'�� Ӆ�ֺ��#{3D��B����M��Kwo���=�Ј#��_�@i�z#�׌v�q�6��'0���	���4��@g'�Jm`���q�x�PޔX���b����_�0���y�A��z����T��R.^��`�C=Ӧ��a"{���=����#�[�,/�|�f�h�����9��?�>T�$̅��)�yh¡�Ϋ�X_���etd�yӲ��ڑ�?��ΐǁ���K\�@OO@�@���!�b�B}!���Mq��#�J���ഉo�s�f|��}���qb4>��`���#khǻ���%?�k+���9(��P�R��L̀ߒ��S�kO���բ��vǣ$�`�|�Im�CUVX�t�,��^0y�2,�GӨ61���u�����ļ�m���*��XlxVHYEB     400     1a0i�����g���������`(3%��w���y�%�j�j���+��\�.md�(��} ������Bg�qK�
�ʑ�H�j�Et�M��5��B�:�̠�v�������O�}�z��h��@�G7Uoe~���w��J�;�ٔ��3+�x��mD�R���rz�O-�C~�\�����a���<ʰM~8	��XP*�o��6cv���6��Hm���]9���bX�A���Z�+6� �Ft�����>;h��Q2�xT�[!��'��2
0�=-�]Sp+�1�D����O�>�j8��p�Ćg-xU�=����y �/��������R��yY�Ө hgby���q
�c<~��'�.�7���s ��t��;���mB/��H�ډt����T����e�#(��L��XlxVHYEB     400     130�	p6'�"�fU���?3�~ׯ�^��k��Ñ�B����V�ª�@�]1���&1{G�z��#��eJ�+z���@�g	5;L�mDu�4�ny�#�v���QNE�� ���p����3�7���&:����p��%o�q��+��D�?Cyf/'G6�@����+� �[k�d�4c��O�i�:ݗ�r.!�ׅ1� ��xc��c{��aS1g_�QPQp�������"��8y{��xr*.d�s���T�QCb6�G�Kh�;�7 ��w.�wǩ`_�R1��wD�]�XlxVHYEB     400     150͂g��tFI�N���tm��ft��/"5���*Ѣs�ꂴ�'�@�����>潗���\�� ��]�g��g�yw�:�f� ������A�[�&�!~@�R*/�"��CAT���mbǺ�ōghRD\����h��H@ԥ�Af4����\/�vT�/��K�r�����k�l��~�8׈�ⶋY��=���ڞҸa��
�u�9���ϻ֠哵��tT������5k>�e�
�7}<C~��U3|� a�F�v�t�C�<�Y�H�p��۴P�NsfP�1����-���z�B��|��$Nb��x|=�gC�^Mu��0�8YG�lXlxVHYEB     400     1a0���K��b��Y%b�}�C��#&!�Y@I�� <�3��4���f�Q�.��� E����^��d�?{[��m�sSf�}R�͋�ܮ���EϹ�L�z�q;p�3�ׅ�֜���X �M�g�_+���b >r��Y����VC�I܆��swG�)V���_��o�<�w��F�ݒ�%��$%U{�B��s�7c�Yq�n���q3:\�Z�<���1������?2l�p�Wf'�O�B�Ұ�b%@�_1D	��o\��=��m���ұSa��ţ�=9&�C2�蓊�<���C�9�Xsۮ t�h�. �?d$������ݳ�&`2��ih�M_�(�4t���{�Y��;�|=c����g��ģq��o��z�QZ�Z;��I�`��[z��:�¶Q�XlxVHYEB     400     180����7h(��3:��5/�cv���	��jfc��@�M��[�����߅�<	dwv�r����`:4�o<K0�`�e8h*�g�A�P8쨂����D�����2������H�wݩ웨���.��2U� ���;���nM���'`���G�4�ҷo^7}�S6<�H�����{J}^�b���k�a��g��t������r`#U��n�.��.�z<i��0'�_3��q��Nem=�P�����������ޕ�þ�|}q�+���O�6>0D����H�6�e<�25��J�1�.�E�^����2y��L�	�sh^���Ue��vg �p��זՑI�V3zs�te��e\Bz��U��;�ժ��[�WR��=#�/XlxVHYEB     3a0     170��R(@TμH5�Z"!�+��_�X��(�@��y���%��K�֛1�]� ��D�{1���3�!����"���Yf^��u6F��$�n����!�#]��zrL4Τ�?5�FN��+O�V,�a�8��A��N�Jthٝ�����l�_� .-��V���5f�Bz&�R8�sp�Dì�2A
D��1&�#��N�g�i�!^���.OR�<����FoSL�>��հ����Y��ry�A0ɴ���y�����2K�h�:� R=��~���ٳ΢+�>x�59������'��֩�z��~��J�J��2�1ԧr�c���!!X��Q˽syw��B���t�I�g�^