��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���� vU���O} *�(Ӛd�ڔ*?�x���*�m(�e�Xה~-�F�g��Tdd8���3sl�%�ڽT<|�4h-0���j.���M���⌬(f�튆s@>d{�6ɹߐ��t���5~�|kbPל�;��j�\$��:j����^��(2A��� ��+����KA#C{�+V���t���I�m�'�AZ)w�h��:v��٧���G���O��!sH��$)3/��8f^&&����/�&��b�Pj���\���E�Ҝ>4�Kt�a6�N�'�v��
x�ףAoh����r�.>\>#���gt}�U�Ĝ{e�����4� ��8 f�2:�^�3`��Im�'��(��
9E�D�8HAW�z`��й����I���Dc)~���������{[�DӘ��=&{<���ỆR~���Q�.�#ROcl#6�ތ�懺�k��[D��TF�ߠS�����StA�����1�&�`��l_zw����n�,�g�a�z�K�4�d9�U���v:�Уeސ���Z�,�����?T�}|�M���A~�ա7�C�|D~,R%}�b-<n1Ԙt�!~g�9ߺ�ʊ}uT�H���rP�	��x�a]7�8U�֪��n���h���!�1F�m9���?�|�{�4�02��%;Z�M�31�v���tC�n�i�Awj ;\����I�V7�}��i�r�I��GS0�)9�2��4d��?�sZ��.�h�\��
�s�_$��/m��r�^@�eDg_��<��ƃ	�w�#���{�p����7���E���F�Q��T��������pf���Z�U�|ww��2hkX�1	��_֑W��o�ye�Ή����WLS:���"C"�Ί��T�������;�\�̆@>�������5��(߬�L�ھ,p1���=����+�IDU1�	"���[�}�������\DN�錳S������������ݛ���O����
=���?|�r�q:��ls5m��Ekw.�>0�r��,k[h��թ?�2:��=�#��6��J�#\]䭿��<ՑT�X�-����v�TX��v�T�!�zY�S��̔ cI���n ���[���Y�����>��;��F\��R���M�_��0�� ���v���(>����(�n���{����7q���Ƨ��gA%��1�J�71�TH��� �9[3;q��njg��t�Co�l�b��#ƣ>i�N˝��Wl����L(>��C"�ɟ^�E 8��sO ��<�}7KLY.?@b�m1ȥ{Ahv��S�p(š[�X�5|E�x�^=]MS�V��o�y?�z`����x��\�P�7��^ǡ��F�����E�=7�C����h;
\�b�E^���KhX0�[��EϝhFP��� g\��W�|��,���(�l 4�~+�<�khC�*��W;:ُ��4V��d������waW6-Ξ����X�u��ΊT�F���|�p �	Z�mSދ��$��s���W*�gB�NP"C��OO�<�) �����i���a�2���pgH9�wk����#멀M�,��*r,ģ���(��7� �q���[�<��������g}�@%�	"�Ӭ�RYL�Nlj]�@�b�)f~n���|�=|8��y4�%�#R��/�X�v���)g�՚�fe� �辝�!��da!��-�-�����`��\)E�ùxr��,Q�g�H4^��c��e�0�js}\�J\󩧶;�jbA��i�%_ʅ3;�o˽�y�򈔆�I�1Q�1��(��Z������!��b����؟���-����\u#�\�a�_%�}�.�-L89��wlu���κ6ߗ���_z���>�VSˑ�bˎD}���6�'��n5 c 3��e���im�)1���gu��u��	�H�h� +�8�m�oo��H��e�v;����T�{�T^�Ol�@���r<�LT��̓�H�tf�0}°"���XC_��-�I|���E1z�����X7 rx�%����h�]A,���ctN�7l�;2�(�8F�GٓC�\e����(�V��$�O����.<Nt�(jm|n��
7�s%�m��d'�c�}�~(�-�^m�?u���Se����}����@İ��S��_6�`���b�RQ�$�����������N1R�N����Ȅ�)�#\*�;����]$ݱ%�ѵ��`�<!��"�� �/�q��)�ǉ�C�2��q�\�]7:A�ߜO�Q��l$d��_����кW�ث�u���TѥP����6v���A,߫�A۴��f���wq�h�T֭��{��b5��v�ďUFd%�\7��d�����~�J�� '�h� ��=TS���Uyt_W��;]Nɟh�����k�j��i�C�g��o�����x��T̟d�͗��
��%�'�q1�7EE��$kC�c�
�N���r3��ڀ
�y��({-��h���߆pL���,���l�wS���p���0�4l>C�)�I�r�;4�B�dI��6�R��^�&�oV��f�M���SL +�Dqe�"h�*,+Gf��c����U��T�i��2��2��#%	%t߷)��3�Gvb2e��Ͱ��s��{X�OJVQ��M����[����B���3�R��6'��l�25��]\h{���c�4���+ѻ����Ň	���<*�x��#'�^Nյ����5P@���(��ʸ�)�m=fI�k��l����;�����t8�CH^�תf�T�m�cDk���;;�!�k�J#�8x(?n@�3��?]������KjMiEΤ��qz{>W�K�9��a��9�f�Pt�����@1л�%̈́U��H
G��W����e�8����	ul��J�֖C@EѮA����n5-'�A"k?)HNV��P�h�\��_�`inf��vc�������ϝ9��T�������� ȩ�+��_�V�� ��QW�L�A}A- ]=�Bt�?@f�㏷���a͠����`����