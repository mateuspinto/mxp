`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7104)
`protect data_block
o6DXWRFU4SBV+7oFD4vCA5kAl/vnIy+sQwJSSYmYwfU4zoUti6qeX8jnHsGI62C3ujgmGrZi6vjS
xZz6sfyXABRsepbI09VYItPuHm7DHEPDsld4pnsV6SeEPSudVDDJyjZQbAQ0OMoM1sW0hPq5+09k
ERnRcbqTCCiIz0UuO0V93C1fjSotVFis+ECXXYBoO+yda4DqPxdNbFyfN8inYy5eRAybd5C7wkBC
dnP9RzAzRHgvJmMipZQKyJ0DcR4t4tUusXSTKh7uDqOS+YefciuU0BJVLZEGGTveRRSi3zE377Sj
LbZS0cuDoG+EUp2sq93njFx5xVq29TnqBOfGhMTsl8nFONeDnJAYzX/UFL9LvdN4h0VKLtTBAYGo
tcJlwirqHo26VQZkOmPrLygH02TYU2hrrygrSZdJZhqaeHwlI/aBsQQ7fk0GLDTGxr2/Re0u5XdU
fHGa7Jam/86PDA3T9JntzqLZDR5mGZ6U+7jbwsIrzvMKr7tPWAN0A2o+1okMVyxMlgeIrxFvMdPF
rGYeXkELZi+VZW1mdckbXa/rwOPmDMTfXRXJVwSbiKITyEgzT23wgCGSzymqEUIDpuMEml4CZKmi
q9wehK95EXJMGuZiTnmaOGj1ZWKxUxZSfTkEfM3JWG8vgFGZR6TALIYnfK2DaWbjAJ+8cjsjENEK
7/rhbeOoK3UlyQg9SXTOijaJLTnqqfuAVTxWLIUDYACgmF6AFrsvoEY1FN+WoUCtIpk0aTPUa7h0
rLPEMJnUZeCp+QbUPiwzcakaDimRtK44qpsWUBkdOcPqaFrLyZYhJTjmiF95pCtp8v50w87hYYZT
RzuSh5mU5XXw9oX6R9U/dc9TZBDWLcKRVFBjRBarK/ppZwXQXBMIt7akMaRUvncdE1XupP+jc6RZ
8LNQ1TopokKdslwobWV6szgPTAYwhmAle8YHL2GYRjoQDnW3gy3R8Mr/uY5ySZ7QbiZpQlhHWZVR
Krct1bZxHchsjBBov4qSiznpkdTS24zg+B04ecnYqF03TtK51F2YdaVZ51BYnfptpGUOKOt03zbc
On+OWq8MnXUe46n+S8/U+CR/i9HNfGgpNj7AWBI+fWguJTm+555BzPu/0GOy3liiNQSKsP2bcxcJ
Htg5THULQEMRLjkA3bPeE39+mWTua+7MnoMUTJxycDxo3ovJolJRCZGUS0QOKlNN/RQT0HFvRupj
iLbYdpgrbSBiU49s8MLwGJ7z4ON0lrFhyliZ6T3heX/XRtXQRWvFeqZqH7nAlzDSbX99IdJ3WP6B
V9K17QMWwEsFZ/k1Q9SVfFIQx1aaiGkoWpyMOhJ8Qukt0rOlFcgQftjOLKpn7A5RvcwXazYx6hH/
Y7QcnZfWLjzpO0ySKjTrJtj+oMEGrw+AY2SUwj/rwDTZeE6ZfCKt8yBT6qLgFwKooJNiAmXIGCuw
m9AWFvGaOPL6VrOm73bP5LwlpLePJC/kP29I45KwP/XISetRdxnjfaobADvAokCQ0DyaOAJaxr1f
SP/OJDwy544Z9wQjyR/SnqenSXLeX6AKGt2rmIdyXf6g0F+t7rV1/xLcnWkSwdDRtxUxRL0VDxMA
eTUftWYHmNQAFwiJ0yqXchoP1OxIK6SN1net9fKSVzeo4Nh8TmGJgwUH8eK5ZNplUAPYm4/huodj
9qzMkz0khzVtdJ7eg5nCw/OJxp9a2MWGnQrlZC5KdQh3aahI4XfnEodJWvSlQ8WUkJAXZ27hNPwp
IdT2xSw/zq4hFfnLLzJyFgjO/pIGjv5aY05EHGbzxyJOkUvWim+4aRioH0J0lh8GMQVtclGVMu4u
Cv/w5Eg08hQB9GpCcrzApjQd0sBhfjS6Qj/gYBM5wgosu/Oj1HEZ1JAO5Sh8Yyacq06cWQTiDcoZ
yPJ74HFilgLahHk8b4hZl2wD/SmqrZ8/+PWEPVdM4HT1DYpzTDlOg+37fPjp4mRCYlzLb3Kx+JmM
9DeKV+/AsliC/mhNwOCGL9/CjZax+ltz4aMMCfpWhID0vX1ToI23V623R7Zm9bqRtxhY/+OW1vjt
mYKxwLS6EUgcQuxKf6O35yDV1kklsrQ5t+uGepyODM4ECYxcvF6oiakC/+iUpTXyquGO4daleD/L
40p4oGjiEq4mZzxQUURmvTLaubJMeiOyfRAurWPrCGOTu2MAWPDV+pxhYQafVWW2OCs8ghxal3lR
622ddSk+spg7BNrKKXzl6FXh9tFhpJY6UYvPYU8tqFpFDQXi0uquu08866JyLLdqT+TgOt9cLQ8E
tFMXdrEpjznzI4DnWJpaa4HgcNbR3zsHa8IeLp+L3HI1VN/7eWOkIYzczmKeV/h1t0f9VBo8K4KR
6gGpuLijm5aetEyNlxB+Ww8R91H2tEJF2PWt3S9wUAJRdzdFvCYrbHZaKACi9szYTUIEJ1qnWe4q
vNoGjPTD+ql1H+Rtko+QDjsnjf9IdDECTWGk0x0OGtaOuBkBdNcnkb6yu8YsOHej51q0SCCCxMNh
4dhB6RrSRUgtvMfnDgUkWLXnBlkFqOBcsF8HSNM+FcBkskIc3KK8QsOUL1v6WZxMHkO0k8V1lGxw
AU21PzqPyHl4FNQscUcTPAryfSJsun1U89IhgSzy38xTGhP/zDj3sKres4erRk/rPCDXi+mZ/a/7
q/TwzMDfjUysRgGZsKsRS8QMEXwo6U8xEIoKTvvBtYFQiCvWo9114XvgAGtw97T3pDkP5/yUGAu0
rPt/fOiX1lMPC8gqaen+EM0WM/Ti/dUMXR35cDn0/23snSeQjWzkivKwtc+mBQG1Mzs6Jc97+p7C
MUWZDqgR7qLxfSKhFPBLO89pj8QUIm9O00dqn/Iya8FP4ZSUWqTisO7KQwtDRAA/OnaDoKvRrxgo
KPyXgpt6Weoke+HEMpk3WKxPFWm3lbNP3uY5OMMDzCDgFAXwQE3lonso2Q7IxaZD4KMgm4pVP5w+
Jdtg9aA6letqoj+0u4e1vGe53NGaz8VrxLaubG7mW4LmZTsQGAKApDR0eGm6cVmC/ZgCwBS66WE4
V+RPqOuC33ZqzLAh++3CL8ua5UJBZjZS2MUmNHb0DnGI9a8w5hEwwmI/1YBfK4f16jwyzsFrz6ju
zKwbbtQdoROTWFJEmTi4mKpcKkqQS3XhnwftOnBrhHIm4A/4shDK/1f7/u+Kk9SKXpFBhWsHwxQC
ludWlSp+xhV3qu0jrOzn/1issIq+NaNXOhAnR1gOVJ9F1CO91YmcymmIykIsqvn082EjyzbIB9wS
98VsTq/+9VLAxOTTOyf8zSEK92yLzGD3C2C0cNGX5vHL3WjJ2FebWVU8EN6heAvFIVIfSokJZknB
FmgwBWDyUe4qaqktf5J18gi37ghkGAHrkT4upyL6x6N8+aLaZo84Qks4ohDtSBkvuadV3PQFapaw
8c81QLjycz68lTWWOsEVxha8XPvIxSpI0rfOn2yG/8jpJhC3jEN26kA7pmSEBKnbS4t1/M/BDVe4
1Ln7l73fgNBa/Ixh8qb0RGghga+yZmKXP5ZyPVj21VmmsKtOkHhNn5T5vbHZVrPtwb/48nczKN7W
Kj/3jY3frK9mH+r9gQ/VBth60/NKHfYmmbnN0Cw0I/RxMIb5eU8PUraOrz8EYQTkb5J2wSv7R7jH
8GtUIi/uy48sD37uSi5++ycfWyvt1VlZmwcc+aWK/Jj4eo7uYsMbCBzc5ckagbagJkFzHbNcxZ1E
sgzxRhHeyzXqgI56oJwpdo00hcHuoQGVGC1fA+ufJzIKFCRsYDtwF+RvxXy1gU61tWvLjymXL2C4
8w8bdWEeDFpEbxLhMC5QuPANGw7uM4MiByCHDhNMZofCUKU9uUg4AaEiosYqJzcuUon646KuTNxS
hB82Ttk/kL5Y3GBhnTWnxsKaM7pmaX0z1HB3w9R9RM+47txfiVjtxBPUKEp8UjKS6H9yPeR3GbEr
Sf0s/SndeE8N9F6p41JtwvlOCQJgvihhI62fK65t4uEYX3qNynnG5PgYcOdM/VEMfMwrUfEHg6DC
TH7lJ5B0VqmRTtGk/ArQG4SyA8eMphrVvpvds/jAgvZx8bxSpYOq9+2QQxNcU97RnuMRoluDSZJl
PdPmEJU9jYm1Njcdn6La8Zyfgh+VQgYc6A28irONyfrz18RSQJY1E1KE3GHAMumFY/BcresTrhhI
jWDFfMrE+ZVOH/jfT/8uDrlOdbOo8jzDlqOmdfFu3HttRrvUpI8TKZVCRWbXtts+FCZQz/wMVzxN
uDZbQXSycHnQMYlIf45KHvVL0Cknf+TB1jVakHnYpUL+n0SIHhPjC0pj8laPrVLJrHiQf+DdLDSA
re8tDQCGZghrngfn3jMtss+cpyFx+p+vdSkOelmmGrwj50TtHd3GbQ/9uFCIVdxYDfXO7HcWhR5Y
oyertMIFBRZbentKu/iG9Lu09WjcssMZ60E6U/fuHO32W6rflrB4zGUlVo/8u47R+FjliAR7L4r1
gkF7jUFmYD1MFGjuHs3G98bButCjk/rMbB/7Fklbz9FbI/eW/Gn469Uee9QAcOlknITsXLVZJu3h
IASGz3Swi5YmXLYyKLF1DCXkU60rT1d52EbcfKkxaIYfB7NvA63QAj4MGI8vtAxzAFpMgprvutZe
yXtatffv4W8iRtQZAx0kizdaAYL2JxSrLL8zMonfrGII///wO+aleeDp6XKsHuAHbCQZ+Up8PNwc
3O9Rh269rK9z7oFFkd58H3ZlNSkpIUwpwAhHssaL4sXc7wf/ZXS/oAzD9osTDUWORmumPEGd7JT3
KyfTRQA5FiCEfCOifeMjJkA3Z5lQeeOEDDMbB+QFE2dcdBnSHeF3N73XKbcvaPRKOH1q3v1y0F79
28w2jfumzxOl9wWJ9acl5T6Kb+v4nzF6MKtdrJtPd/1/LxvG4RnXfXz+FPnarxzp9VctXtRcFsJa
T9Z5vKvUV/r4imMApG7wWzWHSscLfRvMfiJ5oJ8n3rm0ByM0kmEorScjuikbEDULLgmREbdZ61be
/v0XEqvCEtt7wj8tpCYlNB4Grxj5HquqNxM9h9arE6qDUCt8j4aCtoLS6i4fwmP9B4gIGvGyVUlx
94jYsArkp6nD4U9dX2raGnlLkrduRLSDDFbpN6L/FbHFsNHrL6NttSQEQmichM6HTM71OG47F4j6
o+m9gCYpXrvM3Z/dTnhkwM4Um1sG8WOY6uFReHl5QGp1Q6PmnB3RK1OeDR1NfL2wiLQ1k+BUwkvr
bsEBHE0Ngu5qIazsZA0Y6mKR9KZCcIpIRdYW2xWHi/V/vU8te5+HaCH6TkG5muYKO53AjEg+Wb4n
26SRq27f9gXwuJ3r9hY58STzZYZWWHh7xQMUHQ2xDok5HGzGUv6pwquo5I4RofTcL8i3Cuz7WJnO
1f6DnJ1mLA0vNshHzT+c+E/wExdxn6Jrj/WSQ+1Ma6Ap8ChNIXBGLlNj8nmJX8rUEXXF71HrvmPe
t0fjsoWHVRY+TcOeoEu//my6Rh8eHKpTJl1oHMTCUp8DbUUKdWYNCP6fLd7sFa6OBCPHzSJaR5WN
IlSr6LMGxfv5yOsQ8rzWGeM+DdiUsYk8GIVh/XmnPQF1ck4YeeCTKbEwt9oAAoZVB5WqG64TmxiG
DdllhBDv/Z2Rer5EQW0MgvZWxwtxUmcO1MJt0VUMDNmFztMolEwxJZPxNgw30mFW+zTqEQYOXdoj
6oZ0BYmm9aYNQUNoFB3LJJZkddkneoiz3gUzL4rGDDLwD70zVSVIQUsJHo/OMMjDNWwr9rEfA3f8
sKiBsTdTxEjx6phPvWMKbcZoWEQxN3Sa6sEbTqc++O1Ru+EeUa1YKTaZQ6I+9HRSel85Cq4fSFjY
cm4sz3dWL9BGqaJTPd30mi8BWjZkcn9PYbbXDAF9lc3uH+OaoDNtvCmh3qG1JLL5htBhlvhl2QIS
4Edfte/Eto+JI9uApIc2ouP/dVAd7ACazLAAzCivhVonIVqvTzJRfL2zqXDiGZ/ViIBkKN+V8TEV
VqGBUa8edAFP0IL4ZwKrLUpleJruvCPmIQHItFMPmFWyoZNlQEAwneOZ85GjR7dwu+f4f5ppAhgL
OugZtfDGnRFBey1OIxQoMPLGoM+D87KyiA6lo0tWJA0gSlusyT6MuOZo6SVzDOPu11Mn7rKOZUS8
zjmr37d8G/i8r9uakCKIDaPk3nQsEGLoBFgspzB1qZXSBS6izKn6dgNFRtTK8Qdj52UGxAazd56H
9RcLfNM+kVps5XBEe30C7HcK8elOo62tcNSkid540iqwV3v5ZxRTLUnPa/z+DZLJH9Ay5mh26csv
8bKM7pcY70ID57155chCr3FVSSPoLqLEI8QQPuEYUGpeZJZ929KeDRzitVOjRDG+zESEyz2TBeSt
WkXosJeZvstMy3hYRytjqJtb+fXANVSCdfK6kUKivpZCvopBasAe3TxMA/iTR3EvTLd6zYzx+0qe
YQnBN7jdnrc1BNV/Mypwc1wC6KIqBtFVITC4JFoArc1DNo2iCfl3z1qqk2epJnzW3L7UvGhQHwWN
frYFSK1ntnYy0cVFmrKWU8l7tqD8rTdFpQbI1EGHb96qOEpoH5NhZwSMlTbhEypUB+XX/Hqj7Lne
40zBYCchLYQdxKKBl9flOVEALleKjtoydsA8r5u2dnCLqpFaDIkmBcFPoLCEL1SH6ask44DIUJ5R
diq/vbBIVGDrlqqdJKxpsvZMcajP07RJVcAuFvrRlu/i7G9CEoSFkfruhUkUinKyPnfHaFip+U29
TxY05BAE/X0s1xKAC++PJFC8+lkuyaFoazN6h4y/mdrMQwE3CgVEGdbIqb+p3mhSxz2pDvsGULAx
UA5ExWdEzTphOfSGjjJVM7GSWyxAIhYcn78kV+PU/+HNEel9ZNUZYhzNGUzBvHb9iTDWOurmo2SF
qUMQEUWKmwJnpVIpY80P2kn41j3aPuUMbT/oYGMkl59wM9xcHEJGrsgI3qOKKNPiMRH0kj5oUK2L
v2v774lq8PZybOPlGGfR+ChFVoxFeHO2mCd7pHx20k1ZGSiw19Qz5DBOKOyBthce8jKVnOUzdeCi
8LnF3aJFiX/WibSE1ue+KHrT6TWOcFLAe7XcwJgyC0PDEAf23wYah3MVSfOSOyw/h6Y93eb1bUDL
/FhTxNSjrwc6BZWR2QVVy67yKXYrwmUt7ByxnBkMt5JA3wAAKxG8cOU2FZSNjtePwqqTJDRRBc/+
SJYn0pYCebVaPT9k0jUBCNz1i6yxPiKGF7oKYf7WMtFnR6WUX6ga+tIFkiOE9nKRGRCIKnmfebBg
6LMqpkmsaGwIVCkzNZjSNZ1s95VQsAJFVRjHbuvakoRr5MyfLGKJnVdi1L3UESeR8kg4jVbe7Arj
zT1gGbt1+sTfbNTGJRFOGbsSz/5W/TJhaqQMjz9DS+FgqQkeKanCG7PIEMEIzCpcMkX3AuSE66Fv
0YtFkQHq5CCrmSI28Cpq3zqyIZca7zJab0pB6p2QzdcbEBZAalpNCUXbvpL+vE237nbIwbLA//Vt
mR7vQQbTUMdLNt4C04c+0EE4hrOJ8GcAW/DyubuGVwZGSKQhHAmudjSJyRm01iKnSS6f5biqGpRF
hGDky5Yrn8wn0mhpGJcHMOtjJhpkbrKPqLR5W0tJnjyeOO9r3cKR3cdq5bOwn4NAZEs8lUVTS8BQ
CJ/gLwrG2yKlsHTDufGh3mFLJvgF5Jjz6mLm3KJHY5bHCnM1HxjLLq75fRhUtxW7ZHmvjQ/l94lL
yb8v7SPQYf4jJ2ka0C5kB+VsDGynG8zpE2X4McLrb7bFq97ruBK8i4O5YS0GX2ao/7qKS9Pab8Tj
lPKVLPIYSgY4hOk/k2UEqRy06JQ4EQc+WATSnSSk/Qh1EHG4e/ZlTNAziqapk+ak2c4ZgcmmHqtA
ShOx8VywJtxHYdQk9XoNrMq8knz7ZMowmTxpboCT3SQ67IEC0v33l5bE1ZcNEz4Rcx4jJT0FkHxa
4CfHLlFNlbDkdwB+sgLMcK4BQrRWmF6x3i2ui/oG4or8TORktwGSTxVtq9/PrbH8oQ9szvQDo+Q+
Z6B0xYJ2kyB0klypuIiVE3R/yZSqxWXfWEMpYN8qXjem0221wVsKvAuqmGclEOtnDJlpRBoZVyWS
z9G/ffxdcuX/lPVKpa+hoxCOasLFOkdZ3Xf7RrYjPUN16Sx2oMqtFC20k+Wg+T+lgFZ6hruRnsnp
rS/WjgAAJclQanG/JBpmi/Y2pNKvvAecT7j+0SqZq0+taIZWDpBACXXGV9tgg0m6gNJ9bFAwyMvL
8DGsvZ3LOivZr23kaZHyN88ktgqOImv0XwQCOvdJOZ8vfyB0lHjFrlDntTCptDhd7h44sD2hFmdd
s4dQFlVKCX0mThiJ0kLNa59UoVLaHKnYvsUKCLrx+DgQ1Awv4gIJeQmdMoNzXTOKudEjoOUnBC/1
16Fo3e5DUhFOiCxBbIzx70Ks/L8q5h7f6gb9WvKvt2/KH2PzCk08MINPsu6uOYBiRg8fj5+8/U0r
V9eXDZaOwTnJYmyCyMPWP0DDHPnkaanYFy15mm8Iw3Y+gIq0xV5WnmI9GwVd+HOI/HgtJ5S9Ny8g
s1Q6HNrnA2khiegCJuc9rlbDwFS7e1gu2QA6A93NlJXmCJy2NGilVJTqk0iBQHC3WhpWQYeKcvVq
y8Y71Ucc83zpIgJqyPh151XY6XfQ1Q6OYXeMasJX3BZOb2Sa7msvrXrOZarivZXSJHMJZ5bpbZfC
fPtVrISZ5POqHSPy0L88z9jPG/ayZtuLuaH2KtvgULXcMiZIXOf0eNv+5DcSVQbaOWjN1pGy3chA
YWHf8qZ0wgrIJptnhL4rqc/sj2HfwiYotp+3TCT6k3rUlvpoZJtbKcaqFuGh8DhP8wErYzlzjOjn
txxNYU0CX1gdDFpHerF5oMQ+dSBMKHQ+LvDqttK+9wcTHQ2sSy0WMrsfGKwY+KdNQqjcH/pn120B
8HWNQw3eVwZcA2l9h+yizdek/qs++uapix70F32d6q+ztTobCudkXsKxCnEeMEwwMe61oHM5C8tf
t4kOyVx19eYhkarWiEADgzeZp62yh0E6YVTE21YjwHr2mj1tCwOe/f4M4f0GpsviTeYdKFQx8nad
AXbXinNo8kE6TZ58lUXXTQmVKFFtcpgKbJ2TsLdz/BZXxX2543fpLXCeLTzuNDtnU1rlUhK+0P7o
f2VHIrYRbVe7F6rsOGf6fmIk8RL+f96EbxMjtuBtLtCsOCMvgiXs7iisZ4eB9lRxho/2Bdz7t8B7
xGCv3WuSwMxumFzEHQBqleiW4x6Zc8JRTcNdJ9/akgY2HS1iaFdjfLxN8Wy6LLL7UZ2Lovtt8G7V
miuWMNcOF4mthHm/4RZ9IVk/BKpWxNHeFmvdxmUuwuORtsVNq7fgMszCNkmSyM6G57rlpJdGlbSO
vbcd6DqRu5DoUrEfVo5KqteQJPmyHO3cjLtCMMdcwOEdVPdE
`protect end_protected
