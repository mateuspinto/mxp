`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 50912)
`protect data_block
ydae9oxdMuO3Gv1vcwLox016L9Pvt+m1oYcG6wDjX0hCA1PU8pxcO2YJGIPFyVXynVuC0N6+FNiA
KIw9L/QBneA369GEwuZjHlDdS8q1tiejSQw3Tss0ChmCj65mvwRD2a1M78gVSTa766vDHrH+5pR0
c1B9zsPi7dmldd/jtBpFUHM4fn6Rqql3L/CZ8WQsLk39/Y+IBB231QjChVewjTDfjfKVtWDtoZQK
UI8rAx9IRJZfb77PYCGnh1PUxsM8V0wh07MI4S1WdwTvsWJF/gWtQR2lTByEH3c+9ABXbGRy/t0R
DhhsgE4bxAKUAFUBxmymuFRp/A9xsxgc5EQi0NOTb88Tprgk3TzLeIV77nDliqbLFdmsiOe3K7YF
G4aQxa4KqUQSln3us+fty+I0CfSCsKzTV2Rjp9fC+GTueaLQHOpzAl1JRlPtW2gxfTTZ09KQI6rt
gRuTZYM6VfPL/gKM7nsvbLBwaXEWwkCCGC5fCnUN0ErYsguugmkxpO1S8uolHho1mh1OJGDCXUAM
rw5KKUqaOS2WQiFbLKB3r9OlJHBUEAbyrE8I63obEGNODirnNF5AKiNtHZ4oOzVvfE3EuMwFIcIf
c137oA9IyzciHfrIWo1wLjETTH4bi2AKCieiVDPECARyExCiJAjnCWyyDx3Rg/Jjoy7miXyznP1h
NdxVIJlv0JoauQ2lpyjeSk+KSp3o9c4TY2YZ0LnAiT8T5xFYWd/UtFacNrSaY/QOPq3wnjvIluzG
Gpqb4i3tN1qBY5Q7mTCKVcvG5M2ignl8fxGjN/elTl0GyHg6dx5tRjkYgbxH/+AhFIoplHaHY9LF
R+C5pd3bYSsTk0BroSMGYBvxFSVs1zhFKilRyNzVkPPs9Vctu4ZMXHGDgk8mXlb2tToCUrwgaBBz
yIDKqvSBwMZf3uqyOBckzgFs19WDWcDsDIM2dtcBVOCXqgbut2wqXsgyOO+7b+6gGF8XukYroGIt
Prds5ua0CjlireEWXFEqtCn6YLIOxP5EgzaHrj2dJAZXSDKFsdagwEt4lFLo7uxOBaVH+8lMZIfG
l1wgt9EjnKegDdBQW0Kw3PN8ABChun8jxt8F6PbSkNKHoyOWF6arRwOBgCzBpaQ08UM4SufXMsmC
cffcx2r2Yu1YL43E+wtINjHuzsqi1zYGfWURAYtuWLK+unHtaGHAyO7TRXA2evjf7ds9etXUGRSV
i027nH3c3Oha+zgzLyX38qD+POPARuk7twRX0CbOoGcGiecC82dkeh4o3fbdytRismpEW6yTA0Px
m7nAPUu+l9ctF6H6hYFm4GgbWPUfqCQXzRXN/b7cV4yhllZnEEt0iAQ/YuC/w3aH1tkWoGSQsH2O
/bh/9f1Pps+wvx80EcMGhZBuXFE+GfmgXCxyJd5pNc6ZSI9+AIHnHSOIhuAVEVA+pZV8nMOxGiIT
1cenu5av9osUh8mtIID30C916N+Zx9wd3TcZXTCckjKdcTjXlHX6/pIM2lLa0VlNXQGItlyttCDF
DRb50cn4ot6tboBP/UVr5bB9cNa+kObcsSYvA29gN/xb/yoKURFPjnzr6/aBrLDMojtVwr7mArDM
Bri4MNHm59gMLxpq1sfxNHwNSDV4OFiJX4HB3OYPHSZ/dhub0XNqDfgz5/yQ5lqsZfUVSK+K8Kiw
7XQ2LQfMlq33wZErHIQGTYLMlJv4SUZtpRR5S2pXdoNnh3SGQZHX/hUHCwXCyd0/n7PDQG8QilVT
dOFtLGNXQiax8OoihSVYeD1Sh8CbvKX6W5xk2sGU0dfp72EOwPLJMmzQZt/v4122WSpR/OCVsWon
TN58x+rbLlIXOn4pikLM/24HYXi99S+yZI6zsAqA3u2HzbxFkPVYE6YfyAX6dsOomT3H+no7SZ4k
+SyoZ9hPOfpROpz2BdgOhuvLIipC/rztfnEMK+niABCEljS7rYYawU5zMZHLYA/fLqloARerK5x+
gDtkJ7zPOnrvSwKtZzO9g7oa2rq+ewI/W9hAQuUO942M/A3Nt0TA9lL3pj08DL9g+/Pd3eDH1bOb
+qOdTJU5w9PAG1kYgSiFyIWGfBBX2GPWvBvbfSU7dti0DOhQCXjpDgxEEQio4oRtzgYgjVZ2xT9V
dgYlej5TPijuM18b+nuTUox9pclSBUafDqzKPH3nWtJK2Bsvu3XDnQdDhcMKEV+Eg8tw6FiHF8sA
2Kxs6gRhwb5u12kvLmB782OywDDMwy+KEwPuv6II7iPw5s7wiOP2Z8WfsPnO1ZSDoGdGTFuUHcZc
1lyhxdMOM6XAchb4oGlJIWVJHU8WW/+TRdp9jJXBMUepIqNR2eforhRFQLZG+6GpT4rRrfNLaHTs
Tpq9gg1SCv1K8zIAFSwPM5rv9EoHUdT5P0oP6efGax/jbg4WxUTKdPvqztHADCkTHwUg8lfN00T1
euJZNQ+KxJIGvU2d1HhhXl5rn6xi+KdCBYTf+P52arRsXRU3nJrvDvBAXc//iiz4CXUD9r5mgJfM
Z//vueXNOUS3NGZjeR/44Sh/rJi3K8GksxvdZkhudIrU9x8U0wJ91G1tIJpIRdqiFoBCK4cqvL2Q
9HqV9U1HKR9B7KLMpuKvVpXCKaUPHEBAzHbiDX7EUa/803/DO5j9Bw8sNJp43PGlcpp5QQvk0MXv
WWFdZ2ugJf7O6GATjyUoMFkGjD4isDi7pCk+poO9FLtYR/mjRyyE4P0jSP95xolTaT5Qs+mD50tF
D1gGbmWkPAe9JsAiROeP3EAKUMIVYH5qFSAh/iqgdBwFYrKS87P4qhbA/ghfh/czrj5XpL5YxZEh
1R5oquZjSgsO5fp1EneJG0MF+t3wOVx084asRp8y4Up0XTr97XGNNSgKbZjc+aig/beTARVwZ6g2
09UvVJIjx9isw9VHLDEeNlwTbTcam34Fo4t8KfijB8wWcf8TT5zJSMbApWxmC1CmAEBLEgw2hB1P
qALC5hpNKSXKL9WJJu7jCLGOCUKaESziztJ/J8uY9vzqExJoPgYXhE89sj99nN0D/JNeYA3VHzTt
k0VKN/gmR8zuPD7dSQwI1p2MzikbDmIW2OIYb7wsQj1bASAvA9vO9KOhnbtpktfCWUx0nMXb57Zz
dN6wZUrYWSq615Dk1JG+Hjj1qoeIy4WdQWGZENznAy/4A+oW+QWdKuwxlE387+rj441VpfVMvhxG
2VjrgxvnWDfXPMaF//vZcJfzJuy5V1POhatZs+U/YEZm5BHdym7XnONYt34TvVVFFex4rB6+tVTw
kM0sumh4Uy4SaJUoG+L4hSbzY+AR/mmDFh4Z49xS4bhv6HNFvwUgW1JwleI5+hv5UXtWLpTs4Try
xM0I1lcVTDdSe2RoeCAnFVb5mpCMaWhwIKgRLm+LYADX4X1G9osVZC7K+FJBOklJHgHWKnG18Cri
Em0PLjT1KHgpKtBKMzRxmx+U22bEaB6gG+Bk0wsdZlycEYIhNCWhcAWtewDcWgEKVrxsd8uEz4Wy
hRE8vvU/RGgp/12GV9UPpKPZcwfN7wkMQmtWxDUCki46FdabVD4JZ1Ax7khXvbLknBop1By2Ib0S
OLt0cgxHebBt4Jtonr6js/mqjqnO5XnfZsBdUgCayPa7fK0eW7XGq6ObBpG4W9aVbZe0uz2pZFqU
5QLXzhsRx3TgyjQUYZVbnt6YBUExHoxRBHk78ooMh9UlxAtsQKy1a0Q87vLyI/pqm+KvxtlVx6xP
BjHXcqJ1Qd1fDpmGj6laIqbFSmiGPZJiRtjcQ1mBI839l1RDR78O2i11LIlEjTMSoOz5QefOm0Ru
EitG5+tMXRV0sjfii6NIQI1zYYfafNGExOI37M/EiEDYlA+3F3RY4b+GJZxGlAKZse7PslnBHlOy
qGOZCACqtgtpx1H2xWy6jg9tMTFebbL/IALxrFmPUhaJuRqi02IdAFVFl4u6ot78ALEMCc11Nm5A
A2w/cG32Op2tvYE11uDTY7OS7yJfMlb0ADlwvBUycPA/drWOfao3mGk9pEufW4qCH4spTIaWnS3r
yR5i3fQis3ikvuxCYavKGxBUEdU9I1dyikiKsrKF1Y2WLF0w7/5CxbORRpXxO60iQaMndiCPZ+m5
2bA2mk7G8ygqS5zy1fYCjheUoryK/mP6OMC35e/w12nLAGaEOSWkMGRXd3X+BQyxj5B7bqEPIUXg
sTTHUmyfWGYhW2podDIuBI+Su/xbEKTWHSvyjiG8G3CBCMuEzWkRF5xDQoIq7xS5BzqWFwPg0G9v
3ycbrXqXAL8XRV4cbGxeSs/6/16OcoQQy1WYpNa18AO9HZvxlWvuQYcpWGs3M6ZZzAEiHaIaAkaQ
ME/X1rLw6+t5LIal5M1Zqm3B9Ttjw5PXGhZkrAxbVaM6e6hP8ynV1GhnkJQrZJkpBsKeWZQ2gl0L
6woWOl3HYhywSlstQ/2I++8GnLK/F9QJTXxdQTOScuMWERCWgKxWVRW0qydCYrBQyyfoicdHp5t8
id+dny9YuWE0xoE4SQb0vwZxPMY5CZx/RvBMKSW1RDDIeHa/eZCYI6WpNjCYmlmDoA2pfSe2cZp2
Qve1ho4SqdMafcn+KlxVOHnz1qDKeNKqfWWqNjGwiUmZXNrJakYZPS7rVO6JEysxw7uPhYc6pR5L
fyYxOlAl3ON0pFNcnWMSG98VJxKYtIGKxkQg48FMBm2Yt+TrsM7/EQH7poDMV1huUO+FuklIkGaE
HC90XcoJoEJFS1VdxxiUXsKOTWxT8qjlOZ71dWb15dlKVCa0n0W1DqZFcQvJBfVzpMC0QDnp9ggp
ZdeW1/K8raHLHCSR4qKS53WJvWZoo8jo7/rcKbLgKBMvxhytm/Gjw83BofDcavMsUoTG96EE4qd/
8okHkf6MPQEyjLFzEf0oNosJoF13+5BICDnACkXDtSPcjo86GhvtmA1uRf9yC9LgflXwJCM+wPqD
VAH64LuyOg7zPxiX7MeWCylcJBlozNCxk9sTZphB3cKgDkn4242pFmdjlagZglA9IGLncyLXzJWa
Mgv5YS3ld+EkBgnqRLmZz7jXFIwRpGAV2o+MvkR6/F6oWSGqS+GhlY4zmhenSEnVD+VmVqBnhPZc
WPKE8RnIQp2TGgolSK2sAUEtJL/IK1BJNV0Ge30KW4s/coUMM+weZeG/i+UZopqczC7SynIZtRGW
MYPyVpE1eCiaIZplptC/3ep8xyYAj3VkbeNJS1eJAJXehDSH86OuDP7AI4ovCoDxssrwFmKeF6Be
jPVhxQgEedxJpHJT+64oYkpY34kLyOlzh6UjGWRAJAoRIGiLRQeuYDy2ZEb08dVksD4+rh6akDF5
MykG4TfVAUqCKnhhHAzbj7vOZsEXw5iPIQp5FxMgIfdJ1IoO5b5g0qHKY3Cvtcu7lyGUS2C2fLL0
6nwAZAyCNfJ3Cx7E9hMJX9hpAmevKBz3BhpNNV60d2wCEwfS/GkTN7Ct99xObF17D3+LTs/seobP
c1hX5K7k9xKF5RB8Jm/HjnpyRHM5R1yuZ4FxDQn8qcLSxfM3p4+OcDAAmJkeRUzn6uZDTQQj4Dn8
4G3xRNhkdtgS+4nG/IaOuSf6n7yacGdYpJ0Qvtuys6MI+ludbwHdSD9hjIpgeXQ2fj2NFbYWVvX1
AHioy3ApOKk3e52Hww0/0PGtkVTakfzRKS4zBrpDIymb/s8EObJbwMo+O1wLdinm1evW+AUKw3RP
eQ8Q4lkvrprk6syUphaeuP//Ni6SvpZpzvg6yk83T1sJSZIFtB5xGiNpn5U4KytrOlL0XAXwpy6x
boEKBHiu5OXX9c+lFKpgIJY/9ubvNZ90YRTQa+4ix4sLZwZUSwdDGNQVCRvdLcDWdFCmxtKJfQYp
F5c0Szg2BQDNCb1E1GBH+AcYKTcEhqEWKmjowDZtOxcZLW26nMJU4T2gTE0A0MMR29FDqiSI4KUo
RqKEsv12STZJHUCxoOMJAaBkpCZj+bEouEgUhRjolsw27vHsgWXnFM3rJr6L//cPUYKdCqA7Ocf4
UlqnSCSDVrI3RdlxCofXH8Eq4REklm7vfpshdXcywjY4+WR2fJtfe0a6P+TjDPWg7OuSbIf6/hhV
KkLyzQoVGAHSyneMoV5CUVPV8dc4sNyX8i/XtFiPAk9t5i/EfLl9w9H4owA2VpQ0bB0Q2MElIxKW
H8rQ70jaEu7AKhe87V6qiNq0n+T+jOThOSOCj1Q9xc7JVnVCJNt5ZCbAA34vsFefrtRbRB3+TMiY
6k5dsYX0zju0gUBdJhVCQRwt6TbEcJzcEx5PI4L4Sb9ww1Jx+cPPeHBgWAq2DKfAvQIXb7bBohe2
01ifQ7v0FYUNdBDJpAM03FRh6zc8jVBkC5JhkpRyGUjZ1ONGfituSqu8HbpSQ8kMd6bmG/uFhJ97
y9v8iQtwQgJiELbKMwnlZurwFJXmrjrHF65b+8jVkzfcItX5kVaATvtTdL1YiLY6jsXR5Z/f/3xT
Uc25R6KtPltK62hyzLIDCQbxNgsAWebJFrsT3aEb/Zf5F+L8tCUgyX6oyHXPPxS7H81m0M22Jwjm
kBfX24waVSprqTBXUp7UcENlvspL5Pbs+JNMaUksbhG3oi9C8Ez93NvOZCw616KnJd4STYZIGU0L
uLYfCURtgD/600hzkq9LCOPLqmiGGWL/bwwB0CHvT2Gl7utw6ZSarhefrCLGp3Fh+n0HkhDvgrjJ
s0+2jqMZ7KiUQwDqAnEfK5XeR5FKZTSGcrJjYJ0LHeONyQwcuc7rPaiAKyEle+mLiT3L/BfUIJkp
h1dFkqZIFZ8AZdfBrbFdVaGDSSPTqAMe1/HgXmEdXFaCx/Xri4Tzv9iXr13qmkV9LAZGIk6VvXEM
hTEcbXJaLUbyZZDUIm+5EPEJjtnlIn/Fbkogx273H4p6PyHxrLYxxPXsq1XH19QZxk+FZ5TPxmFQ
loA+9QN89RbB62Cb2gPunqk0pdLwIW9XqkaGI5LcbtuUU/ulaWnSbjbgVoRblL/kt4Xvkq5v9TsL
SbEO/YYCGOyEvMCjw87F7RIsIxCmA5M6/5mFjQUu1vzKpNU+bp5ftHQwwXXn25tYxJSDZQY28ehs
p9xcySjvivCbV8KuiTpGvsNHn23muZ5HPfOJxqTOaVNEgXnwx3TKLLWarrrHip/O4GPLV6VTGean
NKQ4Vgnz6tf/4da2lAj1019mFQmV2yZ9TwO2PqS0gdAasxF2kdKAGD2i0OWxyq/7bEHF4luS8mMQ
9g8AxQol3t4mOdYo02+/yY9+9ai3WX0EQV9gBy7SJs7tjw8MhD/QANC3YF0W4VZavq3ic6aNBLOS
+4pb/ps15mvQuEnvEYngeZDdoRKRClA1Q/kSwvFZcPGypyPYQRoG0meojUMdtpL85joI22hFYKhF
6yItwrVw1EPlNtOmCUqemtpijU1tzL5dJHsv76mseF9aDpvR8fnxSbIGcCFGT99tFsdK9J9PHvzq
XE9zOUsYfe9zBj/umX6LKZHSFx8LIhyqTA5TTyFq2y7QYhiC3PuNZ9Ioy6rSTI/jXECqswbSo+Uk
7TNwZw+J/OtHxxGVjFu2eMdin3sCnrVKdFTjitWwmlw0DAV0zjpbcZy9+woAbQGcTx2sg37APLXW
w4/Yyf4UdQ59B/TIcqT0/P6h1F0FV/DE7ZOos3i33Bm/AaPpR+0qhhVRqDJj3tf6gkClSUK47JyU
EDeqWlaht6VH5/96z7fy3SgmC4gjkdBQQ1lnO+evBBJX4NZx3Apj8jMW2D5uD6I7Zc1Y/qcDYBKS
aTdGvEJUVRiE69cCRzOkjdLG8udy+CEEHAJqGQctvkzaUKl5T49reHkYLAZ0zg8L3g+JkwPr2uKP
3wklIhP6uUlGAmI+vx2pYH7PlQSPjnZX3UONbvKEMBzuZOuhN5QqPktZqyjtJrZP/FgKrZ3b12F+
lgC2K2J2a7NbN8tPDN6OpNieXWunWKKs697c2lAJwSOeUtkU96WkJkuMkn5GNpeZoXs7GRIj6zrM
2Ss+zmiVCi+UQa+UpjFtp6MSLZs4JJ5dU8G9zxUq75dOzlSqtU4Gyax2vra33ihs64aOcSkqs6eH
dkAFJ0cDtxhZCaAd5MUF+GIbdiCe30KVoAIDjbLGwK6C7ZNd9QzMFYkmFRBzrMobqxmLtbX9bMkc
GofYWEEp5HCA0UNWiCZ3mkOlEfYtgOlsXw8F3Mjj8l7u0tyP8Tggd8VHV/gM5dZi6IOKn6NYi9Ig
amgNRdcRKru1yuIBfn22UXyJg4MaW1g3Pq75Yi2KFDrb/IlkAfMlN5pe56L3470x1fZdt48WMv0x
TlYAANG6sOid/+vo4iPQa5BmAr+A4oiOeDW7Wqtl/VcP2yZGzqdJg/ZmuNmvp1cLJX2tcTqRXfla
fNRb6JzdlmlS/Pf/9K5J1E7UZxYcrQKgiVyhkcqqiyFZizaNo3mtqfdaOwgvcUT/UYImInDUid76
IjOYM+/Dy+F8qyt7iv9U33eRk3o+zet4kunoTUhwKpyCmaD1mnUc3YIZTKjBc0ZIRmONTGywu4zI
UsvHQMaYADmvqmBnHIirk71YrUNuDhXuLs9lX42ChdPwzFp5KOImOfVY1F7ZQrMWu0IxXxlEonxW
W95ZodiMYgmCNjMhsmNfaOdpXMmm/5yu/ygHpDqn/iuhG9HsGSCCOcXulBiI57qPo5j2mJCdQ60G
U1w10787xAe+IqGlp6VAkkLzX0UEuxUtWj34H01ykczxyPuNfMLtgAblSPR2u2ABZg/exkyqqq4N
WenG0JX2utJc836HuOjgAmlEIdLBbVkE0kyCsWGLPd6j9H+1GnWtuDJnGvaO9JRT4tU+XdknHYOM
iu9s6oyiDx4Loojhq/iUmu0nqk54ahmK50JE11TfssYjjs8hMHDxxaL7EpFeAoS3p3K8bR5r0Zw9
k/hF7EhoNrvN6XZ1gQy6eBJDvO9BGFqOiZoKHI2rAxbcvWtXRm457OoUIYG6i9WD9zUpBR0KNRdh
T+Rm9bDPU1bGEjePPCnJZxlDSH1vn4AxZ/nZtPm77O4gfsHjkN06LmnRvCeJOIar270hV/CaMJaH
n+pkH9neeZY0eJJSDTyYIFAC4eeuPmpAizk+yUr40uORYx9ADLnnTJzgNRc9KVs9FKH3nweC0uly
K3BBS72y6R6WsN1rvu3d+9UXaQv6H+T/we2b98NdY4ZIkug1TmAaWUZoOKZkVH4UQFZ4ywqKYx4u
ehENxaBp3ywF4dts3B0IDcoaYm8qT9qrMo/goD8V7jFzCSW7sRl//vtCbFdn1qOwyBQY6oDeDTCg
9jyn/ixN22ZcrpS/XOfkdZ008Lx+EEN0+9moUe/vOu18ScKWO6BWfSwcyiwWGogp3TAv5XKPJ9pJ
AUS2/QwkSX7nnoAl8Gjf70lxCRO5OxMoiVpluATpZwQwqq5hq4LcJUgm6KrGQfm/0nhdfjz3/fSr
fzEHjRPHYRUZ9Coyg4Yb2mtph0bGvnoeSMJ6qGn7Sl4aLIW+johc3lfyuGfA1wXW8L4wSGqGOrS7
dDi1zSBgmjbGAa4yDTzAIb+95jcJfq7RBWJpqj6MGOqkPtkuW5hYnY1vy280WeBymQ65E0gbSIXG
MQvgEFph6oPN5a5+8xlLZV0qWqOi6dPS7GU4zRyGLmtFAaq7x/iVRu2fZngHTUjpxWKnyCNhgqfn
S9zq9A71qN/7Hl3pYK2ihqLZc+pHXtBMtz2YQ20v9BiyfztuRZGDFQyzZwnCCa3vPMALVjd5KkW/
jwrAG6flJgT2ohyVvFNhzMzx/I+XIIeH7x9AiKtvqVe339urBR5A0MypyuBT+bEmFTnnWJKtwqww
kREFR0Kj24l4wOmw3dVt01C1X0O7qKQqaVPzNk9B0+4ff3xUPBIyhEG2u1+kZ2N9CeFVEfBj8sUd
xeMfRBY4MBTck/WPabhJ2FOuoEChLziSmJY+hL0wkZexIUOb9i7Nt8eq+liztSLGQfOCLdsFxszi
wlzsuqgaBoMBsSjsSPXpJKy65ll3WOOVUkvr85zsktJ9sVJ83XDeb+lupyzZBOusvXI3MiWVbZU4
AGLkoQG/T7LtitoDyb08bKU58Lztplz++jsp4W7JaVqslYDiVZ3ZHS0+GFOIVyZeiGbQI0tZgLYU
IQTJ2jWPTyaxKm8OSjnzrdBbtUr8Fzlj1zh3AnZKcWKrYrtwGa1x08209gazilt/ESobS7wHvtQI
RFhms/ZwCBWmibL5mxLL91Eyw27YzAub/BqpROUkuMVcI/kpdJHN5BujetAWV7Hiaw9h9JaIxjPC
277iZmt9+XAr6QGmuX3Z4sMZ7CzCtmPqaY+PV5i1QkXnwVQY5g+4x8bOZ9aqTr/orPnXEwuzugq5
dtbP2nfiPei5RzAkRPQ/gmiGlazcJzTHejIm0kE3N7ZEmAbaTAzQXQXdjBVyeG/Nah5khql/OZWn
nsUgcULgnEbk1kvq3Ez2/Ct+AiIEfdMYJvJxk2Ku8lMEmDEihG2vXLe4Efl0p3Jey6sjkGmsv2Hw
nH2VBkCl0z9OePKDnlGLuHbx1n985MX38DEV2b+lDMUNfnyYpI4+PxLgt4rKXBT8c6CzUNa7kSTn
6At3or/msvix8hpUzVZDbbaufkVKLP1nb+5lyFuHxG1Hjn2UigrEsnF8Qlx5UdyG6fbmMHLXsa1k
SaN/h1zn0nN+wwD32Qnp16rUof0JE3bzwOR8qhYKmYIMI9yRlaFQAafME4ZwO7v8AF6NrPMLA/ba
ud3fVrZjScIpl1lEbO08LpOF57oNGg2Th6meaWPGK4ionIPZ/Iy8SBnqZSUxZT7WE63bk/vV9aTA
7XH7VIPecgS3dq8O5qVPWYmkgm2jCNCyWsK7rSL7zks+XaMSHA7Su/g4zOYKbRruNVVaxrwX261N
1DoPXbF124vGb3JgPLuHL8QKnD5oH+dul/FKCkIOHM2G2xJcYea7QITXggOXTnWtewevnOLKDL1d
DSH1Ictos5DcWswIgM0NUycBUbJ1Z1jBDIFr2GuD06JTh1AhIJykJf9IFPpEsXHOIok8Fyc4BH3l
gNORFnhiMZGuILDVWUB6PQvGA8gcmPDkwDGAfUdJNk9VPVu6osQAbFzfURAsDImDzfTKThgFZv/6
dd7ZcMuLb/cpEf6N/WSYKgZQj+Ot6chxwVHMOSo9elleFvHjsC+9wB+ZPCGVWHBmCE0VDDQYFrLv
5ivLTnfa2j6hoGS8+od8tmekIJp/WI40os/Xq1AzC6Y1CuieXtanucvvvDtoBeypkZSaM1B3vaLD
MFPxqdzDhuT+sNG4MckzJ5vOs0W6qOJ1OMLV6fUz8pEvprHsda9m9l8OCoaX/WotGgXkwhfYqYkD
h6PRkFHzigDAxSojxH8OGB4YuHZglmRXX0geOJHaYBLQzC1jK+QZ16V+GzBxx0zVqUKmgmMbWpbe
iBfu5SF0lE9nBMYR2wTFry8lyoo4js3yH+cuPMM9WCc/O/r43iuwYL6pajLd6DOvmEcuuM9PU9AE
t56YwPqrvTmX3SDHVxwuFqLBHYlL8V6HrfcRIsSwh4bCVu+EW3Bl01Jw1EaMATnDjuVCGZvyOoa5
IckT7dIP1Hou9W9GqsuTZ95K/CVF/JLXhEOw01TzbrxQs4G51d1wW/L4iJPE1RBkdaHtyKr3Fqfb
JC01WJGhTR59TkV0bv17OQg/plJuLshkEWstKdJhd/wAeCPxDVFqNnn6lLie60TIQJpNmPRqS8dY
tYjGZtoz2YabJFwyhI9d9lOhsF8YqQVZUqCQK8yLjz7odCl2grJMbkd5rZKRqvs1hT/dcbeVY/80
D+1aoP3z6RhDoM4GngzYpoTxE3pCdS6lGlcgiWgT3dvi9nDbS703F4IzcoT9nBEULW9X2L/pL0YJ
0vVMsfL3kH1HijQayb5UreXQ+lAE36tmukMMKU4A+o9Xux4X6jTUibzJbmZkteKDPN7L5RpbjIGD
9ij6R8QSoSFjNWbp/1VQhBZOfE9MPovuhTT8QWlB+yzJsKJ1vA4aFNE7RkQY543+t8hoaRrsDz2U
WucdXUzwV+XNr35ssyhCMu5sxu2e4ILmoR47gmuTHNi6/Yt2Ss+78E3dffy8mtw3UI5RI6PC5bDe
dlEUolCdFbADYxUjSgbjxW3Ya0f0uUmebda8bo66S0ZmEdQUsh5jD1X/C769i57UkDzXHzoQXXau
UcyJelRQHiJOxY/CxIWOuLrRDJXYaMX+aCKXeQWlqqEY77/boKWz8McYWgP3yD6l3p20RTs50IuP
NTnEY0T2jvmiH9Rlw/+leCH5KeUinTg8dE5/4BBj1ktVeAQ2ea01cFZI45pW+l1njtHTEnrHYt/U
1/ScV44dw94E18tqE3+7yf6Nz+IX7djeKH3k81zJ4GMlFP26zCDSyXDa2O3SHLpghdqxdA1nqmDw
fesou4boi3aiRh4g/TwBbFEpQMDf+iQ4UOiTa98/5H74rTPrfxGu9W4PxIEpEyX077EoNvwmJeoH
8Rd1t03+48kreGf+GH0bjxo615YtV+Sc2YRQWPNI6a3gVwddKlYLd1YEW5fKyoHqQ98OT8WwxuXG
ssD2HmXpO0VWDrhy1LccMJn5u4bHxLtZFMhUt/Q7aaUJJt8aVavxvnVMh+XWsUiTA7OyZE3eI9ru
hyYHb9+3uKXCJmFVV2GTUMUly55Y5PmaoXawRGA9R+o6ADHgYqnrPp1QAxMEW7znWppBM8q+/4MA
JY/2x9HZldOxi43qaeojRxmrKFiFexiJWjEdlH/iE7KdWff5r02ObPx5tb7QJdXqttIsRO5vCXD1
W2Yc1V5aVMzycotNIAaoAbxpMFkM9jsITOaQTEJfRMcTwx6mrOOphs19PQClDNKoZTJiq6Foh2So
LIlJemmzS7yYVfC0YLZzmk7KAyzhdUqQkl+A9SefN1Xug1EF08P/xBYroyFpa04L6jNUZt5fAhpV
L6Uw30BTK7KzuQb2f95K7r1qc7lpXbAJnQhYO/2iwt6lWjUD3qgtal6TQlPcRSWDxKmByCuTHFfZ
9vgFgOC5WFCz747egDWlJL/xUaoOKGI2KZu5SlxqjyRhyCjX1DiCin7Y1v0sMggCTk75nHwE0sk1
tKOxC8YtgPXeoxrAuzU1EjQMutTsnTlluYskIpziagMENbXQtcP1JXE9AOJAy+BmsN7Lx1Pe+OA0
zJtVJCOrqHC5si7klJoPsSM4nEY65iyBA6IMSZI6YZ9f9zJrLIf8R0fWLypjpb7TYHHEWTBuk6+j
CyMsktSjGMGlPWZqthOuTDJLrAAfxUG+kBji2L4KdXRW17PcC32+g1mmzqA47vYEyyEKop8TdPle
2oR7kNiZ5x0+iNAJg34nljq/2A6IxNPb2yZxr3pRRfU7edyiffAjEJtnepjNKoE8qjdzZ3FTaW5Y
T17HeDEfiCcbfCqN6PPN7jGYkNDPde+/wP7kxFbWH+o9P+wpykd+dvpNZ0zYAtvodEgi+m6xbyy5
MysLzFuLevm3agj9rI960m6CkxnNGanYFNHQNFLKm+/lmHIlKXrnr+Tmhskt9Lv6gTHxfxuXKdII
btj2fSEbSyEE7ua0rxOogAuvDHlxAEtxmMYwCf7mt1EDiH3gSvRXqt92fX80xrj1QgvBpDq65CJ3
atmqicwNx8L39g1qEybuntD6RodJhFzokshpt1aEmUiTnkKj/c2qfPahQdwNrA9djFHCCZ8+2uRj
4A0w5SOAvqziJxY2+VZDPORZ7/n1+3P6XUsYnqWO2LSmGzzslPHsksxpdDycSfH41bTtJGQKBsgt
FY2SvoDz7r/ke3ZAOt5bB5CMbP4O57pwFYsA1WxaWNlMw+NKtvKshdw4KTnhAEhmfhBn4/b0jWD6
N07laVedxKaez1EaPkagFHJ+sqCj95ML0rfwG4kXgueerpLzHpItt7nnE70JkwQXFJtsp0FNwof2
k39ZB4k/v5CEaKZfQIbXZVJIEsEEWAEmxQpSxYvMkCKRRqGl9N3NOsAtrEDzWMYGyecUULVQxzcU
6ZcF2VIWYdR5E+smw2EzwyDdsCLWNyh6HdbEdiJiZ5dmxq5Vq8Uwhw1/GoMmvyuntFG00AlXddRb
i43xl4dbSXfQqZszzoldz56IaqZeb888n0h3AL6tMQNtqRsSPuv2k3Id9oeMeyFXfCiyb32lP7Cg
7GtB8MTHtVRgY7Wq+E/UezybBZMAv/yYaGQ1D0b11xUm5Kw0AiKm4g+lbbF10pM4NxN0deYJ4TU8
8CCkg9XcsdAL/6FCwpUkdX1HpPgBltZcbc3n44TZt8egU+d10aNn1Xlm3FsNcPNKsxWswYDhUk+9
9HQ1OX/CTP6AnoxA4MqPuW0Xoie+zioXpBM7NaCYTzeqt6gCrgu+5GLTCE5OTFYDtnk8B174QNTN
K3Hs1AeF36ANiCTlq1RjVnIIHeEgNgegIpeik1G7qlzHCJjeNn+0gJVSUnfOW0Z/plqQyBjxwDVh
9vtrVXg+zgYedlWdfUf45CMQ72vag7FI+vVkC7CeuknVMYPNI05aez/JEiFPdU0HR5B7JR2s/l6l
LYMbJMAz7PX5VFhDp/AwDs0coOqCCXjng6OPuEFCXiuXO50HF73a+tXk8/bS4A/d1BjsOgANiMzJ
cb7ZlFxXjTlc2jIPWkM11NmE69/tMaj6lmMrnn8WNLNAZn+7hfb4S7jvIwo5xxeKjaAEPF6c66D7
fLLVs0yq2FQCphu9t+qw/Jy7jzxsk71tDNthxhgRznupEn0mtEsXk+R87y3qT6U1NeBk7twUspaw
PL6Tgson4UvESoDWoO5KSdGjAdZznhUCnutKOt+NVGQfJerM4ykOqKPsWUesz/2PcJxjhY/8BZld
7wOumwrIwimIO6W7o6VkZ24aQoHTEBQgntrJtMwoXqgOBEJV6RzOvx+C27SpqyzouErADr/C++Ns
sq8tBDoBSSCkVqgDIUJyyxMhlIHgprj0QCfPPJzR3RKggnZV0Md8F4DgNjSulCo0zh5tnMtsQpFA
sJAhYQdnwfqLQsis1NoneNIgPiFzcPMVJyfSeoq9Lq6CKCw7FVut8o7Ojlg4VwkGeuSDcQ3lOIkS
istILVEE3R/KrxPQwzslXveiM3Wcdc+K7U0yaiAfPHX55WKJW5TtAPjzX3IcL/eDjjWx8N5X2LyU
1qGcFHlL6h7yT+8UX6h1UdSKywjOXhmFa/1blD8MCtuAHOUKwjEb0orj3t9mQtSPAMCpbLBknmhl
x5zjG+lfEZ6+iT/ShNSJ9Yg61TdyrNxS09MOT0EZyyrtj3atdrI3QDc+PXGDRrtMteV2ryISCO7m
gYqRVe8Jk9IupH5XJc/Cm9F62P76f6X5EZfhxdhdHLC0IFa5tKPnjR9gEGd/btnQArG4FotFv1+j
QqkbtRDTyAreSV7cVfivF6n4gjMceSYjdYS2YwsRddHt4JLjCNvA7O4WEuWjgiEBTAjRnG5TFpm9
19bQE16dtYQ8DXUXpHTYxD1MUSrWNNYwgJ5g7BSo7j3CUhmilXXbnzNh2CNG4rSHKM/H2JgWyEx1
NQG8f3YUArTNPwVJ5l53wJ0w5nHX3fyuffyHh8AbwRV5tToe69gMVkshNb3MK3/9jwcJ0B51PjYT
dcETFlNgG+nTgmQL5VfoWp1S3A9yhyjY11EbOi+9FP5/QnrQCnjtbUAjexc6cNachUEHN4EEI7z3
Wcibfm6eE2S4DjOSnFrKJklRY1oQOug40iaymYpC0eFDNn9F+Jl5U5qYMrq+JydSm2EyXNkCf0pH
TYZEwWG70gnynRgyWJ8/pQJWi1AWGyWVJ+4+F3QT6lADMtwO5KKvndhIcb9jqpPRfVU06uIE0wMG
HlzBeSb4BhIJPvCUua8WuEyw8utBGc/+55/28XXNe5KohZoxRsWPNzt/IS4VlKBiyq3spv5mzC8v
E7wuanRSYaNh8DI1+Jit+mAlo56dDeerMAnMXgUb7B5Hq6BaDWlLL25iGbHhnQVBJt2lbsTr/Gki
XGoEu6m+pAcz+gMHlhLGBCxjC4QDbEogXJzrRLgLIp/sRpBrP8Mva52Y+jz+lLBh1kvlXi0E60Oj
ue6txuapRhqemWIwt4GQwVMqjF9jdsHS881qQNILb1XugjinsHrBaqyziZpCtyAz6DvhQNrRP9he
S21IoNvFYISUUmZV7uLabkWpj16Cb0CIm8551PvvEJLpIM3D6qm8f59X2gEyagw6nJlwpsPvPkdU
hxovqMB8CWxwyulZmDh/PIZyJz/SLol/GeqA751mSY7wqMLMIMFLbNyi5TP3PQH2zkl5nmVE98US
41m+0MJ04T4nQ1v7lWoCW7B1CAUbQLcRks6MOdXpKUue9SeTBYGHW8TsIzN7Tt3Qp1LwJF9UM/uW
Bmq1aj5SOAnL+qayy+ewRzkJRKMpv6IMKjKHjBO+8YxsfrQ7TKLrAFGIWzMvnwpkvZ8jWD4mhA9m
ZxK67I24KkVr1NongKSBucMqLN2RYmYFRR8Fnr4EhysTIttJgyv/4avMRU6rQ76+D9UUgHXpPHu/
j129btiYqi4NLhQn2HiPCFA+UdTzixPYUFogbYkj7YeztbXZupzmMag6EyXs5ScH4xU26UChDQwK
UAFl2KmLHUg65Sutda7Uu3tui4lRsSKW2Cm7rxq/eyGk2TJ/VjUqaeuRauTh11hrO+oN3Xoh+XFt
0uaHGYqh+pWmEkMjPj4t01VE+BVlELWNf2/m0VyEe8IWsDU//FfrtFBJYcVpPW+zkd6J7sjRWXHo
7t4A5qmYUpCtLxm1fqL4NjuEHNjbAEOhKxBFkTVeXBa4ObHw97ypdtYMEe+JYQFfgLFcMKz1w94w
49CMSu+qM4bqGWtiDjRHPks3jLB76IUc2mAuFb7qAR8HCkWB+3A7Eihv6ru5QO8aW9J2lx4b/bYo
RXxNn3JzxVCZLehVHDJR9zNrUzvrFqQAJPuU38HOptNdwQ/zQwLqbf+X4SyFuyc/T9yTDRfWDpxq
RfRBUTskWvcoOeuOIcfsLSiI9jiDQW1bTXVe5VihjxF4b3Tj3YoMAwb5PRvhPv1dne+nB3iW2uhw
IXb9CgW1/h5nyhJRZVeN+dglcgx4AUS/efkwOQNm8Wt3jwbLXrViLJ9PScIKHNhksc/SpLLdx66a
1gX+X60IIUfTOFyyQcsJWRz57cwsLo/1JYeH7+Vx1k/Rj2lFgO8ZnslKVMJe11ynGb3N1/PK73CA
+Z/xdxiaCv3omZ0XrHfdgIaskK30jle/s65wIx6Gj2/woDdOUfs3WLHmiJ/h09nGy5bxJTF20bpE
+g3jDsWw8B25S+/e2Cra+d92263zr9jASIi43UBuCPAl/URTBZrX5TrlWtG4eTvj0CzeaDS4CjuA
7wDbR+VbKR0ZSREhI+aT0EoI3QNw3tYJXgs8nIk04vqU+M/u3zE23wXz+dT84ZGU0znR25jBgN70
2HtAdaVAxGqajsdIqRXVI04NkOIekcO9vuNbF4B7K537HP1tV/6BTDqx3HVHT4NX8ZwHVcSg07uj
SqNsNfGZ98+SG3n9vkC/1jhIjHGOrmFecp1A2ZrnPGk5+Sa3Mkm7ICI8KsAYY8nr+LkkJYVupCVZ
W+kgQ6CtlteI204v57ihWMgiawzviTvuE/KhWxiOxKh/lpzjjTQO/0b/VqzJeYPhSpfKqr1r9NZf
iWK7ubM0+QaVeVRNzfr0kJ53jC24Yf610Z0MIxRswYA5ihP5t8tkog5A8EMIZo7JE8PSAM7csng7
MPqm+8ltMDeug+ElJm7gjehtPjUDOUScVrt/zBKB+QssHHv5vR/fQy6HJNDtO9KkChW0RVXUyeKA
RRFM9tqiiRXP2Cw7fra3idHz7wSn6c8e07AmWT5ZdqIzKDMaBt3VGca8T8ZAZTXdECEoyJ7qAcXo
ufroj5wlXrsjXbg3wh0Iu4EjgnQoz5+KL9Sqp7cKHlMPGi2zeby0ibG0h+CNm0J/C2poHMPn0kJy
z/j4Y5BSOMD6XjLrZvnEPHg+1/avxXwkkyo1pBpH71nPcUEi1IXD2JsW9KQjNzFVXfrHhKNHqqh2
Jq5vB6/zrhyMa82jMjLy9MqNdvprbQQDqDx4u83PvIQ3z7E+WKlM58FNtwp9zURcgHRShvNabM9U
OW8YtvdRW1ynWc11879lDgDNgulOSg771McfckWqvw0WMBCDGk4Rqbl8B5cyUrRSRWRw2NGBON2Z
35ScpGQIDKqeJLr0vkO0Gf/HBbmybxS/tKxhtJ9mpk7qy0tNmLUcfgMUFqDaTysV0FHFn1FH6//W
PUSf/MDaO0ijNxf9tb7lln1VSHremoFh1ZylRa4MzphlXUChgfm1ImAobxPNHH57seHWYWt6FZHI
mMWlm2/mjB7OmVJFOTUmwRB5lsTassE6cHpa4jvcXEVo3qoUT5kkYV1gi+as1D7+zwk0IWmr8fS8
NmyyweZobaGPLAsS6Vt2SU2WzRuPeFRQZV1c5LmBovNNt4VVeA8tPnT68LSGXb1Xynd8maSgHydG
4+jgmnVo52VRCtjrTlYwpctW82Vn81+uuNceaVUWd4XiVN5OWiEpbTrsRt+fJb37OrO/leoGrhVP
tTXCXIep6KCYeUDbRa+dMysbMornQ4MQbbqy0HbGJEnlstBjp3bvY+8WJBlv0t2zQ8u0Q5oRoegw
IQQ4a/oWbFqzGtj7IvKBiXso/BPsPAewMOhHeW+YYEOnM3jIdAzVbiffor877A8N0RfJBgbif34m
7wP5hEAs51LNRkC6aRzPlHP38hatG94xUeRsi7j84zgDIN8I1jqncWBn0RWDAL2KcV3fY9LcDatr
9sYBUzPycgdbN/kT2LtNhF7LPgm4+oHbvmjp9t/AT2OyOGzhv62acWlFpyL3YiWhRdabhcQwVqR4
aSZfKSaB9Eom2LygHGgD+8EvnqaOy33ptJ4ejfDuYxjjTu1o0/N6vlC/WI4bBrO2wcvLprlLO2oB
D6xPl2XYsukpzjyKhYJW62uPDecZft86ldLr5xvjjGq+FKkPyb1CUem1ANdK78aTfm5/nGUwn7e3
9yozgSM0wLnmynscTjYzspavYFLvkDepyATVDi4+4qGiDWpIWBzcLLFpRfH2+8szDh0lLlyT+W4F
zCRD4xB/ZhSX9tgpPqga3RFm0+fszrN7W0fOijBMxEsgkRlkzVt3p5f4hmr0JUdmMK2EWyzfUq0x
ADvOzSPhG/h61Zp98o3yINQxBmXf3tr8ah2AUQMSaCJm9vnMA/5JprJ0hU0N2MiAxe8Q7exEuffz
w0pExAYiolP9QRHAKwwzJ/k7gUWJ2wVvdV441VK5dTz0xlwuhQzBjYSRno2ia+0VyclEYA/KrYih
1Emn0WTrMiOcWhHCdvLLXfxD3x3aoJgfP03bQOqfEPAC5emGPkahYskZYQqq6DPB7K1+i1N5E3sO
sxmifv1kCsGz0C7kQbp0fMS6BA5h0PzuW/ayLoVxKJcqV+tqP4SSYCijagHLZZR6IMaNkRUOdtdq
u08n9N2YJ9ftvUELGgdZXFJCmNx2orQ/6KJXiZKDXpVkm9o60dEfhQ+JmoPjGOsFbwXcRQMTQBjx
KGnk3P1Kssg0wUgCsNbHrlV1yN+YY8nzlij72qS0HJoBlU4Nlja1lIehhbfYAnVf9rEblwYM2Rfl
MqfHrhxF19tvEMpBZO4jVqdEEFHozrqWfCPdownGWwyPs/ncLBf47vu7S7n9UsBrK2S+C3H7Rw3r
qEurI9nOswlXT6k++x3m+4Nfu9bVoa/l2rgaoySz1m69Vq3ZJOrjwWXhQuMExSqYccQm2sf+dvHN
TqssXftBnxVn841dWKEuFjyzbywKUd75RE7XV2XBdhv+cxJnKeH5/kf4mT8PBNI4/S/IxIt8kOpL
TQCVoLw26n21lTxu6R/2J00/mDHyD7xBEUIvcvl0mNblj9Ax3l6yrOBWqkV5zmpUZDhqzEc8dIUe
iQ88QsXY83ECZLN68SRXk58gGjx4yoLUD0gseLuOV9ayPfg5LEuKqzc5oquMZ/OAhif92Fq66wIg
nfsJX8dI0BvRyoE4PuVQ9/jtMEguKnVGh3+qWSshxjALxOyLVtvTuyQx0fcHK6U+B6+fz4pXbQfe
XARF3xVSN43RcLEzltOXH5MMgAmtFsSaK8PiYGR1qxn8H9LrSMkMJ5HOCHRis0lWfhF3VpqRVYzZ
EP0A6n2r7TVpzRhJq3MpYk8qUzfu+30d2yfqlQXPTw5PwIqP2f0d8Uz8j963UuDiF1RXrt7ZN7gt
p9ysJbj4lf6/UOj02R4zUpghld8bh95JGh26jaiOzAz2xDyGv/vyszTzeZ04UQ5qd2OlhkPiIyaI
kxSKFx04ots2bNbN4jTaFDspBMqjoX4cEptS8wcuRtr2iZ0uBr0WzJCVpCNstCjChW8S1ytDavvP
VWD7m2ciZOlEkt6hVO7yRenpugZZjf6xOFbnT9vlIysc5dSewckiI5TPZwfXXndS5XVJMDEcksgU
l3o5oJACCNZKbawRzi/MBt8zOqEXZ5MeLb7ZQhCj3M96NcFmecxjejlK/E4oflp+CEBHg0Ai4BKO
htgeqSOaXPhAVcWDlYWiHeYLXSkfIbh9H5nEa/vM1R+jWO5f7cAKYA0g+jgMEgo/gGDGMYC+m3OR
wDFiJWuHpsLdnSaSVbMiWcuXZC/5i6WJopz3OwXGsg9xdZK+RhetaOJ8Ez5t6jrCRbXPi/WfWcnq
6Jqx53pnrrziGwtxdKIrVda28zW+FjFfrHUWC/eGLEpAmKLRervkgrQYRdPUwF/L1Mua0y8sHWiL
4W4wYd0c3Cbl1YcJ+U6e0bsAUsbrGtn28SsEsVqhX8wrkc2GueXmANTNkfL+FUiWUiRDUJDBxpuA
8BWlV1PoLb7H6a2LajiT8MEx8shN1dFyY1ljBgotGbkzAL/Ch6HmrpxliMKvIpFT7/fC/2e9R6xe
TFDQnPv7KDZw0uiTsauZ+r3gr9uD9ilTT4B/vL13O8T7Gk/tNizeTddrBrnl0e0SFu7Yy24E7Kgc
woHgfqqcMdanP4aSF0Gi361OB2VVajiwXbjEx27Z6v1n5PqwLUgkxYmGgNK4LlW5dwqWyGMpxIDP
l9d44rmVMcNH9P5philFCTxks//qpO6i92o+SbUnST2nnQvhmZe1ol7qUeKGE/fM8NyOcNMfRi+o
MSDK57TgvoC1BPRQm32j6glhAJ4uBn1VeVgIC1NuK48GyyEp6addHr/hP9zXnwxUdNBxzcRP4OmF
FZLsfDdiMGHsfY4t8+UIzq1vbjtXap3T2+hzaRhikRuX1Qs6uwzKZPsUdEWBVdTEAD+57m9Ckkyq
TgULN8iV7YKVyNPn8m+P+8zAesr/BKJYQrmyAN/8xXQRXqhlFOmkk2YR41Ix08zNMo6PNsbpNDh8
zdldPxnxfv1naQoeaUWNIQepro02fHcTbRL51q16f2WfFs3Wqiv76aImL/fr13hUGKA14mllHdFj
Z9g8rgcF79DaxWcScf3RkKuWnEk7FPevZA9oeGJqDmttsVAa/+C/753X1kVRkAHsvxc+cGn/qCp8
curPrM4PpNX2UIgNjbMOMfZRE18KoWZTfdgtkJNGjl9+lOwI9fSbPCBL62UMqvljnxXoevZO2BEZ
0jQzIpy3719vO78/aW/NBwBrSFdIsPL+dHcsSUJspX1xPDls1F/EcuHO7DFxBaGYQNylbbOUeldY
ful9gbpG44YLT8OC309u5FAyoyC5ZVPohkREC1RwyilZ8aFaa5xgmcqI6x9pIRq5lMCskh46tmRf
VN8MnrLLA8itnd2/t6tSIXnqtU0BZLA0aTkvnQ/V4r39SrPoY91KqnORtqkrzphdh7Y9JTAG3XCR
09zRhxN24l0aqzn+V8m0pqHd4sO23Uu83jA4RHLJpgfnQlhgCA85cZUuenm/MpaZFLK/aqLkevni
mmEhSMN8yFHZsJ+9AHvmOYc8Ez/Xpw7NLxY8iTHo89G7xYF0mBx1v0sS1nFGPQGPgs619dMaZRUO
jQcicfCFMwp5XQ1GcWb3n4OlaQvHVLOWqTXcT5d1bNTQfTvSXCginGNHPPA2kFUvruCl13U67Agk
uL7nOP03Hz3vOHsgZe3u5L3/INpO8HWaZrvA3UzJYhbtUMrM4JOiSIyAvwgdBjZhjxdW0X798wFh
VTfb4an/Fq/aboYCffTkfD36T6SKEosoCFvOzk9V+JX67jotJeBEQU1lLExKITkjzK/ziVtrcqIG
3+dwceHShpBAmw000DtPj3MrJx7jfBOSmxQ9V2iof0OW1O1qo6ZrBHQbjQBATRekF+M/Q5bft7QE
s7jCr08PGTGEF8nzLDofsN/mJ88Muz419PZL7GpaoEE8wwyUEqFrReXtpX+/w1duYQHtvNSvQHfi
51UE0sJ4qxSN6qoEau9H2+kfI3sACWba7b2wP8ZJfWAH4iJDmqGWQtK6kTpOskxKIB9+N6T0sRsB
9DuHlVbw9se5xc4ZdRkn6Bv4NxymHgNuCwvFhRXJhy4BgwV2lgF1VYSOw9nvo5kLWhNluQvhytmU
J3r1r95MKREXUhcJEWcMsZUh+OlLOg3EtwkG+FD0nF/dTb4TGraGelrxt3TY+RxHs1Dd4sOPadMY
B5lo9G5hXBQ37w7vbQzr3cuEBTCSdrIuCG/kf7YB4mLO78OfU5gkWuVrRaUH2sGyKmK6vCgk5SGu
Bbcj40z2mE7YjJK3uGhfiF1o/Sylg2zJnpkLUU3i0uF+NXt3G8boYKAP1q9vFOUt0x1T9pOLRFyi
O+E0QLY+3KUV6F0pRiZpFkwoplM0RcxjgwNyR5zJnJJRxsLEbEeYtPXH322tcaCxxFRBBeDq2piN
RARhfKfI6p94XTZV//furQFLw5XH0qrqgYwW5ATer9VNqqdn1d+eGPLbR5W0eMqDnfZvfuY674TU
X0R2jeG0HaeN8U6TWGPX+oW0nw31I2WiHahOHQiwrb+2Tfewy7pJi/dhD30c5H/uTtWWk7DAufCd
2xogjs8h83/CWrzI0N7CkQZwpiN/rTlkZbIE6ELu4Li2MirMvyLbBwTU/zOzgVCJy3AZMRjwbCVL
fhZzsCyCtSu7p8Nz/EjuupyHKRGAgM+yqSWT43+Wvar2CuDQyCIWf1WXh2s2GlPC0c9pn20pMUoi
I4W1DQDH8cS9RDXMHYGpzpik88GBhf0pVwzrsBh985PX9hQmmgzAVoBJC/cAZG/MMQWB9zrzqviF
okIkAszHF7vT3Po3HBmOeAl+ugYz6PzOFSWkIwevbeyfFkoEmMs1HfejlU9pppyAFzLS4ct9Vt9z
bt6LvzoV04c5gwchK3sdycZEW+TtNBaSrWtwtRiRQAoTjXunXrnrYLutJpttKaPXSs267RdPfSnD
jwy9A57l/6T8tJkjtVJyeEjVNToY7P3ChlLhWTEIVvNcHYpqFnSOMeJUXlDQMjpnDMmFTVTM+smV
F14jmz4CvghUvfA82rixj7nBJGOP1eseNgctLu7lnVbbkMuw3uaLM1G7+FQKHefM6YtZOwsxY10X
r1XgLPJ/MHJXboehlhqekp5DMj2PJN8rimqUS11RSlEIV9EAjy3k0Wse67QoNNsIFNwPVQKsak35
Cirs2nITyASQea4b0DYIYHalceEXs3Okb2AAiVyrNZlT2qkiaEBWJRxxthJhUnimiHxVyVWyKCIc
Uf12kOQoaaw/VKEzAUsuk2+yxoVppQfy+O7kWrQlMKpDhg5BCUXEddFeW+SG8opIm+cBXKrPps6Z
F7Z3PygQbCQbqL5t9YQdaaklZT19MgFmrM0MSkXhS0/bMVagvjI6jy48EKKUgo97P0h5DPv5VoGz
hNNl6f5iO6u1wsmny4D8aabFA/SAJu3+wcY9jgkyVKgMyakoeMwfQuYMSk3dqe0iMYSrzooVb/af
MHaYm/1qEWs6hj8SWDI0sx3bByPvJfABk5OYB2TYaR9ScfPWpbrhlYkIhPGU1070vuxUmtat/qM9
jbrBCTdXw1F1WLToNMKSmZa1BVCFqbVYNVp+995if+zdHYeksa6cBoh6Q99Z73340xZVVh6hn9GJ
hMtoUyCMRE4k5GenzF1rQa8x+YMOaUnk5hcULJEurR0yzp13V2h4RByoe7jKjgDnBYnTghCTk4tz
rEnHqledgFNE2cMBqiD6gQETs3v229yzw0Epf4slSwof+4TkNlRlBVSLeSymKH8dUTlzTI088Kni
OE/tmZUSkegTzOKNVb9o7e5/9DAYfneUvFdxxGsE9jI3wHYKnKA+1NxUlyZFddTANgdTapyDoZLn
gCtu0KPcoMbrSjDiPNBxxuB3+uMZWqZAlE+NQ7B2v0yG91UNxHMFJEUPpZfU+GV2W5pWtC15D+ID
acSb/2F52I3ucibp1Rb2kwyakLjCJfvKbdMj2IO5dvTSpRcnTOySlhB/d/a9qjTB9j2gs1JV02gg
I+SrwIp3RJEPLlH3WrNFwreIKZJFnwX1SuN4aK5/oJ/mcYYun4KssoXeZvWgKJ92AJrU1ZRMah1n
f1vM43wrslNk1P9oq2756VeIAyhf0ZPWhsu57o2dCm+yAdxTP3BsruwOVqv0fVvNGiT4dy0wBRaz
Z412N1doe6XSLsrjExMKnCsojLB2lsrSMyOpeL0rcsGrzzsrw9dzBgZmTNx7+BMFScyHA6ZwMyn9
naLtYL84uVSzuFCs5qNl7pv3XKn4WhRCimfaQJeVAzfQ/r/NR1hDQw89VDNu9p6dZAX6DzJXvxUy
wfsmasABn5eZzSeewQnT6Jvn8q0+bsefK8mt3J38hUKGdRRj9QOO1UjSJ/adu19l0eStMmVmv+gQ
EAb/YWJJZ32AJH49U4KGf7Ce3t9duI7KMW+JAAY9nNuEUxJyJqAGOP/811gVhub0lqfmEDmRTAih
UVNBX2H+zjHcQKqIe4SkkWZJIWA3La+AS9Ho1kwUeLDvUdkYGGzz7hP3JG6RkewLlF/47SW3LV0m
Sh1ieaZn16HEVNbiIww+hVe7e6APK7dhTsJ7aQIaNI/RawozO7/uzq4hh21+zK3nLPJi8eLLofkZ
HllDxl6fVm4MW+KPQICTawbVeHjSV4sjZHOOwkzE5DrXqxyebPL5q6npPQNrEvENgLfYoxl9TfvP
mGa7yTSmBvxfw/foMxqaz08Rnrq9SDBIitQYE2tnx3+Qh3Wm+XJbdYYHq5TPX0XfFbBAFwoNRYvZ
nQs4xtVizP8QIaWm9V2Nn0g8IPOGKOpRfUfyW7HLw2vddsx1yMkpqUE44eDusjYGAWen1GFRASwh
f5NgMJDOZE0x8r/lqzRaq3v+PX+63tzgkPlgmXAegZgn5XbAFpstPtbeLoy80FeoAKVHFG0kCSvW
FzjsSmEZC761cpa9AjgM4o2LT6YXGuw646PQ5HOucBEjusCzGreSTH4YA554IGURFsWkbNQ/VQcF
6lQNgn7Z/cEdjoqDPq2p87dBrTlBg/jMaajzKGHDR7wTBvJ46fjNmSXiLNrFMXbbhgCIqS84UnC0
65DgMUN5eYU20P9udn6hatpEE6j9DVT/3NQ2Camy4cL4y24+meryh0CcyyUM39x+YhZ372+tRu90
81bc/EMpywYKlQz8wmjqmy/Foz3bqaqgY4omIIt2AHJK9J59NkvGjto5IOPaMbfLLoJ6U77GT/bM
+izsqdgmnNEXmb+obOT279Sw4LpYxpJyBGQzNQWhTo+PwSv5zNRtI5nqN6VvO0lGUad0BNG69jBB
yqX7UGIalE3prHkXS9b9LnW8DONSdgI0eAJ6Ci3F2fcDJF/2CWSLPhAPps0YM+79CeeLtT27xZQP
uHzoZrCb0YJZd1WN1dEc3mQJoGdluvsnqJjD77MX7Zztt4Vthqz/nqjV4U07NCdF/kc5WccMZsxZ
NnyJWxGYfgYmrkNAJTWrPcFCDnGl4AsLdhnoXSj7Rp/FdwXIJNs3he1zeSb4vqV0VdH2rPEjgZrl
nhMWnYi+Uz4Jpgy86hoZ+xgYBsrVbTZQRa9ou4WIyerIcXSbrZuYNa6TPs9q9KdtL4c2giOP2U+d
5COfe+1E+x3mJRWxNZ3aPepSx77q3Ou9OQf3LS6P8QJtS8IKIMsFNB5AI6+YgxQat1T01v5PhvLU
vv3aDaN2P6/focQ8Ogze1zWbYsHmhj0SDytJMgSyejGvvEPbwXUt7ym06q9jfsvjpT+DXlCSN3be
QDqNCWLVzuDDlPb9wXuszWJomSd83N//Pm+nmvCJS0+ERoLHjGy/hhIdbCpw1cBRM7tYoc8sprr2
elXqjYc/HI9XyvCMMqysjAUJs+lf9jVD6x28ZqcXLs/585lxl1GZ6cwuy1ZIN2q0keJFL9I6r4yo
ELSe3q9AG/dG4dvHTVO2VOUvsrSRcRpe2QQaDkHdXMfEyYJjYihwOb4yCzLhzChVKETO955wetqA
bgzXQH/vL7tTfzHuUfzvkFjSywUI3ExLVZED3z1HTl6Fs2sZTzwC58NoWMAnFSITqS0S+CRQY30V
zwhEHAlisiwyV/C2zGWX+geWAl+R3EImLfmDY+TsVZe7mgj7yKQvWWUb432pFCrB34YLJcDsxJwR
eN8DcEG5wfiLbTYz3BuxnzAUR/EyyIiHdUFbBN0ilz47BZ9wJOWXzj+Bfn+cy1xhhQsN7ecWU8ag
b9bcqaVOpVWwEZadmJ11jkxHuYlBtazU+fd8OK/50MR6vps+LsbddUZd1gUDFet7pepqRSVZHslj
x8Bmu6La9mYCXH9glLP7TI2X+VNRM7j1IPPhI5w9pNOAsOkdR9cWRTtS0VGG5MGSSJlktMwL+dBb
mMdyGfEVBd93Pi/6pIgXFCPNakxzFWpGptM/Jotpi0aQKJxfnnj4Gd8qE0ygV1GUAWd3SYuvsw1E
EBWF6CQqobzfA+CHdFerRDwTUyR3NLNMKu0G/4hySAM87S7wWJHMu33ugAmHpH+uYX1APSiUCQ+j
8bQYJRKl9RO+4LO7kMfqenZVAvSaKA/1fK4kQCQmkHwL0rvnlZJXvTJDXSdwnSIS8QsVNZ/3M6p4
DdRKEwQb7WqbMSnpGHjuD77lypdrUVWWcMfzF1LY7/S/vIde+oJ6kBhqZMiwwLKgoojAjDi1ZHkN
OQF0Rn+/5Semv/rODJispQbcimKPVbVWIpAGupgEy9kCaMHl4pjvQS+xcQsUtIMJLX3htxnZ50NS
hlgKZO7EeuSqHMkFDliD5s6ml4HRz5NQ9nT99pv7g3MArJm+wxSIZW5GkMFh88wDZgJ6N/F5gF5O
rbfRixYrIO8RC/wb9QvHyeNg6T+Ktuy1LLi5BX6SyF8QwcFHAAAK++nKpPwgjrp9jQYq9BF0jlsx
XhoeIZt9ly9Pjbiaa2mB3RJ9VeCqhUalj4eWzxQUwiThqvFzWJ/pMHyqARIH/+rlrCtOe/ASdzvH
7KzLD/WKJyElc42ICxfSF8T6lz8EwwKs5sa4AO18XuIXi5HZKVz5rnonXvrWWv4Cyh0fMC4wVsS3
b80ig25E0a7uuSAuwSLAOBcPcStpTBlopIwzWiklUZpGLb7N95bl8VF/mTGGlHIy0C4U1NKT+wuA
Wnsh0QCcpaOTOy632bwzAieTgTu7Jqnm11qwTQ58wHbVygBVFb+PTlYsCdFYH4hyWoDYIWRtRMj5
RIhm2siI1fSc2aIdQAzXtVKu4H9qcDNqiVJjBHrLoKIDwjfPLImWrQRT4imaf4th1vs32+JUaby4
Nj6ePI8s/Zjz6CJsKNzddESdOLG7RJMZINDuO2e+PauYIWhZ/bAd9nDg5XWAaprogtNIhRXAjo/k
TxOLa82RGiQudW1tGm8G5+Z9qWBCn1PDhFFSn7Ac0Um/+4x9WjDtGK/rpC3mtFib3GcKcKDtOgSc
MSTMVy3hPib+IOT/LcUx5D40QxF1XopqOrcYfl5LgTe7sCDIn7NCL9L7uB7N/fYMduan+fnhsPa2
x16PdhP2Yvz8MGGfloi/AxFjZsU0qtreaGpEYQjzNF70IsUVgvUev86WoYraHGe+LyhImLd8ftZa
nB6LL9jcCpFvW9waIz0/juWR7BWPG+3xLtfmA9tVC40sW8G/tBgeJUd059XKeRY3Ecpf8fQBxLBk
Ajo/h7JJIUd84zEwZS+2LpzgCSZIU8cn2n3UEVUVymTe2uhv+o7hgvkxT212rTvEU788oARWg6w1
L7uz7IgDbBnj6pRti0UeR4LAG+gpiL4OjGA76rmw1g9/F/0amN0lu10g4Fj4KFbs6pCPzeFXFLQm
rl3f7DQ+SSHS1rwUC439dDXatCgT5AEDBsNe7LDnZdaws3lZZ+YgtIOTC8uFpllW2zh5cHctkqXn
WBGbEXcW63wQQ1ZgK650Hbizh8HzjHcpwgXYMWeqruXEuTAzRJRGOJA+rU0LocHuSK1rl0E2oyVG
5vbltMN3ff5eKhfFFQFHF0RQWQCAFAEVXq+4rR85Av2JIVXmIV+TbxDbCndj6N67JfvefpDw/gnR
nuZTfSHFkA5isBmO1ILwk14ou6Z9j7SCfFzk7hI3XZDYNsND6SpW9xTmTfT7PJwXVdMeod8Trpwl
PDmZYOZJSxfu+soeHQgc272SCBokhylj6RiFwy7DCZnA1aA6rOeL3KF8IgjZHxRahR/lkY596jvS
rkViH5E/dG1M5PBpX6ahZp7NH6nFR0E836ksZM5sRd0mH8pRdapuguRZUghRXnQ6CGzoLGR0dMKI
OIoz14ltoc5KS24Ok37hNYOQI5b+IgiytcBoaHRELFZ1iNHzKMprD+u0caeNjfWMJ7TxU3654xo1
vhCydAqQQthia34V5NIA31mnFPHkqzU5H3qGUveUIjfroBIZn0RTqrrSCW7pPv9O2n/lbQ2nND/2
ckFVDZ0NyZGRd+vwNxjGi8qbvnw2dhrUZHq/PUoNQPs9XDT5k+M4U4VgSnyfclACuQoo30mKffLj
KGdgVy5YqumTgQnU3ArSzexuqPkXOARfp7BvF+uJ/2w2dF1Nczgg6cR4v8Dv+uHZuCD9OduVlopb
ypd1D4hKwJHnhKkNzbIrs+DqnRy9o/Vg9/UHq5AarGnf/D/+SJf16pO1ONMmNQ5LnZJ2DX/VwG6h
+JkQrtzLcVXj2hcNkKcBfHIxfFKZ3Mzkx3AYMz/8mNPCk/mEmkiPzR5e5ew0IRqZnKfoAKOrFpHG
+JK6t5v5z4dDgT1MzzuUY0o3OoBB91tYeQyMn0tk/8U7rBcZnCuQYijjqkrHQjiH9ZkrGgtlYv8X
QIbMmoXBkvVWYGZqEEtnSKEjEXxCOsqpBrid9ncjI+LKpZcSNbLKT23mFKNIz/oAZabGVqDEROu9
bwvnxLR7COyOp39uwVoZ7YoKrdWWRlg1OwXpiX3lhKzW4zqShkBlLCXKvTI1BNCUblQyfLkQ8iqQ
yje3ga5QByJ8VoLs8Fr6aMZ1kucFzJ3PnmFJO+cRjknTr1JN1U4ok7iaobpIJaOAJtPuo8mTJKYU
Gez9ji/7Qn54pV9OqKhPRycqaUGfKpfUOf1PkDMVYKxwjLD0O3AIdrylMoDkXgpMFb22sOjaQOHn
6DdgXvilZM0XZO9nm/549Pm3DMYpF5F2oWh/VB6FeVSkzRXNkl/hMdFl+TVboBW61Y8OCL9CyYyi
l0xf27wQlW/JXKD6dp+AIH31dbj1xoFBRDLvH0+ssWF4zgbchY12O1g3ufXItbsT4zejBxNz/6Hg
fucOEPvWOCo1zHkeISDaef00hCHcShHstKv+HmiW7xp+g/BvHTgGdjudYo9JNvBQYx7GEwWKt7g3
NlaDyqUW+u49cjG5SSv2k/cblvzS2BwdKQp8PXrVDyrE17uUffhVtQ1fAKVXwdkUl/H/p+oFiWeW
DShFMpfDBaZzqMElyv5IwRUYAFoCeAxUhwEQzQxjrty3zzZSkmGe9ogouRZ6zrY983f9iel3XUeI
GeO6qqjxcZ/3ZMm4VA4crmKNjSsHvFq5V1Lt6PV0QPffSsZJk1Gc41qFBQOUZ8m3k4zNFvkFPprK
TO9EgCP4t+DwcCt6sOFRftFp0rCX0L30g60pyprFwACOvFhi5zEUuPrfsy1af0EvMw86SgDUUgbp
b7FAp85f9rFBU4iPuMZZLF4PiyPVZz+6KpLiOZ1xy8AEPLFmeeZfNkojT2GPbj4Hjrshg2niD4pr
fb8l4GVVH2av7OnEHBm22GCCQSA48Z9qxgfvbamskq1EGmELktf1eC8hQ6tuI0aXmNJL68tnko6u
b0M3uBVf/WMmze/BnBZFYgIPA7yYy/ndnzgF75LzGMlqwB3HXTQpcBwALQZfteR2EE38QbEp0rZe
afspJSqxCMdWyzVr/VUjp5BWQN0zVfuKt/98IX/q4+NFvwvGqoeyNEwbkIyunqTIepl6H1kGIlGW
xtR9W1RYV0TpfA2I8fRDNpgOhtjNUxFpYuu72rOjhpJbzkJYYEM893p/BkXE4ipRQj+FB3tT1nFS
GHFs1hBrpwJmeZcu2bfSwd9+V241eJPRaodnbsthMBKn8Q7TkD8NhQyZEt8xNoWxXzI+AiKGKpXk
oRq6AT8o6CaTGborBAYzDdU2XSry2EgLnV+a1nNGebqHvpasqqjKtenQWatijiu47g3CoNFQ8u35
ocKMPJs4HCgA6ATXMaxoN6uLbbIogyR+IoZjBhT0SRLUzMi3Y9agJXcfu4kXsysAfiquKJgFwcyp
MphFdIenxzeAHLqlZ+RwNxbV9uAwdKavYbVWq09zEOYGXYaavVIOHJUQCq75R9qut4rJLo5viIMP
I+GfWngtAoH9DOKx5ynbpeSzrRdJOSeRy8L56Bl4cM/BFF8ptGUmj7eqQ4yZsEkT9MLNuzm/4oqu
A+cYJzEulXbNtVQBVbYTPM0GgosPK4tkCUzhxow4QHKoLyfmIPzwJXRoODfKdJ17lFamqUtNk0Wb
ho2kpAWuEjwQXe8K2WuZmqXcLpGj0CYCLJgTLm57uNxHbpXchxmNWuASJfWluhNIs/TnopyETmpl
4auKwJ1YtGBWIZo0bQgy5lhvSaKTIZUU7LPxXeHEjSBljXGGJSx14mRNOZpuO1dTD/zgJrnr6T8t
POxbxp1eACtyW7v2tQQ9AiS4Yx31CYjLXCKvQN3LaqkrOBtAcmnH96AnaQI++ebCFh0tgTVLXAtB
6hqkBDirwDGmJjNIR6efjkX2hCeqNPiYJQDOqcsnpo2RcTDpHqVg7FORS6Wux5Nu9pdIYRbyKqiS
+kWAxg2fQh/ldEt5BROd/+zf3DLTLlK+U/315aT+WwOmpSwwg4Ta8l5/JN3Cx1K99ev94PWrHLh2
b1KxXLhE13rdRRp0RJ4fP53N9lh/8K7cF4Sgzq4UrrK8HYG/jCxa9T9DYrGwjar+ty1HzIyHiyJB
xEwJQX8hvw7FewToINhlpbzL6PN4Mn4l6i8b9ZPeslEt8OmcK6eP3XDXUfC9QCR2dbvKKg2b8dEs
AfecBBZQU/QyIhZ7M/lvZRSPZ3YqLntHBesL45IvTsXjKFeV/IOkcfsh/6vtdKs3tYnuUD1kUEsN
yaJ6zMv1jW8LKxwpbMzzry44VX80wyLAAh7TzumHbG4UJ/gnt/hzW3UZvg1dHmq2gWn8YIVvCGKC
xwlZQq/sFFoDvM9dwTQmoEtJ9axByUfMU/0B3AY8PsxOsdt4q2hEUq/LnH/knOmUdbDV8pySGQCh
YZ/OJAMRoo9EmUM1pn1WdbWuqBt6GoDjALkCuJAsO7c6Hg3j9Xop7dTZ++5lACM9DvulGdHyiyFK
AbQuto7uWPyQE/sRulZdOWwZDYs/btcoyAlwiI6n3clwF+5fJLxYkBAklyrHMROxvYj7hNRvneRh
kDHmIW/6BsUVkpmvcS3ssYwKypmy1UD+lRFa8MR+VvCMk8nqoS/pEGXvlbBKohkuK5E+DcadXdwf
xugSjfRc8c0vqW0tFta9dTTorgVRqfJgAct1IxjazFXNspBLd+71xtLztioBkLww/lBlVtkNtnnN
zOKFQCOq15WgGGx+DFQ6ok508i9C1CEkkOfvUnrCdmW+7264ZmqYMReZDLWSOtTuJs8ZNp64SYha
TM/90i6qHRcobcWPCS0jXE1sBVRsupR5WV8eRj63XtJR2yjFeFvN+IMkS9xGLLjFxrdjaSjuKGZv
/NTQL9z9mpJm9dmXEMpJPMfjHjGMjBB/wCCO60nXT1S4SqECwytlaACX9JBAXm5HtI9O91R/uLTA
VUs//6gTkUHBSEjl9+vKyVPObzpysCJzrWeaAvlnxDPfLFPr8ZXSJpYKIla2//1xiPBOUToePAL8
5FsxzRVUp8jefPXEITMdSXJK9vwem2hFDJTCFU8cU9T+WHzQi09D5iQcL3KkGHny4UMNuk37kArQ
hnXMcCbxWzF2e4H61ha8gCYwbAu1aXhAieM2g3FaOOX267OOV97qwrdlbh0flNLf8J1dmkOIwOYK
5+ueuIMpHXiqoV7B/dfKithXjHzWos/H75eApGB2+3bVmsmoZ6zNtXTfxQa94Xs7DDkCo2RmSNgR
HXbEdr8gxx4S9+gv2cGhEXZracho77gDenynGloEBsJI9UF0T7nGgiDuMvkOylO7X0eTysRD7E3r
UNIDw2iLOD/sUuClnXyEV8ou6YRDWlOU0aIIeMiHhe3zgushWNSru34952k7cyKsQlC6lLhbU21/
RmDchWzsuo2wV4xKW91A6Hu/GF8Xq24Krmh3iEAE8YspE1vQAvsQTHdzeGpCOo3QflvGpGquym9A
M89e2uBmMAxyIMgOlftHubsSZmiMwZYKvg+gP7JPY6I+Ly7ucdg/O1B0eMoyaa3t/INJ8FTrib/e
wlR72Um44vg14uQcwx3iVupqcSECE8+yUB9OZPtemwxS2u24R0GGdi/Y2hwbQyWzPcKzMlluIf+1
PjWmFSR5lufWpsOIaZ1pf0YnoGV4qE2jvw5gLY2OOcpDYcqA3aLxsBX//8UWLBh0e4yx+wLjICfr
rL2K6Q+Q5OAofzlzgxHSGOZbD1i63IiUmjAr33O/pBfhH0HlsFIByUAMGO3cxCOL6XRWdvLmNB5P
gr/XezQLy1Ol4C+HmmfYeY/t+9FBhxoY57PGB3coIYwklICtheIMs5Cb/Yzc6U7zPulSaBBs7buy
IyimnwHqYh4Vt0rGVEmpa9g4sVkoY23KXLJHUwrOlSAn+apskXh9PdmJnP2dqA9mNvBTk1oCQG0s
bChu7fMMLgkk6krP7Ym8LLDu/kvO7vSvQHTPrK8MlxFRsBKtl+qBFo564PYUCFBb9HXzYcbboOrx
YYo6v6SnyRcuGA1LxpVmNl6+/5MF0FYcQ1uXqMo9XmKiRXK+7eNOAL5ZPczms5WOaTlnfjYnAZm1
fJ/QoCTBquKAJM8K06Db6xM7RU7c6CJHolC1rCKYXoEpwfw0kc8YGmsbziDzEvDE4KihHhCBWk54
afXryxY70qrZ2p5wywc1LJEyJGRCZeqcH1Oefep95l0DDNI2cORGp/1eeDWOOOrQZFeCxG+Xna2c
L6fY6gL9kg4KRpEFaQWOQ54xX0joOULPRZphioA0vbrh0ictV/ScKkOAITzEwT0b34kgPQCqCVF3
unesd54Lf6ZIwMle47U/BgdJW+yilLhJGwMJoxByHRX29D7Xevj/uNOsfLjKV8yfJwFSktMhMU4m
5Y+zf91NkFcxl875ynjON0BxQHWiI8GaZ6FYBrD/eLFkFQN63+Y6SjSNfJk08e1lP1a+da0c/wdd
Dnt4HnNhMnftkZq4RhOgecIC6cKWOmT+qwymILFGeppcmUSXjj8btB3AllpSxybPkq6utNDS0nkG
3Auq1e7k0jQo0apI1W3G/jAATj0XzEpyYEfKzHgMFzQ511BnwiqYEIr9h6hLTbqbPOatg/M9uHWR
1qlwkEXJYcjGd8X0Dz/NTUH3aG6X/VOczQTFnDZ7HAJx8NCK4GnKnCY3rMbSvTV7o5dGH/381Agf
mp4iyaEM9c3+U46Pke4RrDlsx1Dej9w/8UwlCnmKTnj3tmryaGhI0oiHqahOR+RHEnc/XEMKiSh2
W4y2RLNTZ42rUnkF5jt2/w1/uKKiLE/f6Ckg5Z4/gpNYhv9EmaIW34jwshPQ1hk+Y/k5KBVnMpBa
IT/9AZbzgUuOP8y1q7q/hZ/4wyrzwIuomcfgRWDzAxc42eU001QfYaYumwgYvXFGhPjbTJoa0hXX
sgKXI3oJgLRAVf2j4a64CVxyPJxY2ruqpbdN6Nrh2KrPtpiJymF7kdmXQ8nw7uVXVnHUvgCllmJC
R8bWkS5QLqbW0idoZlh0hlCSRQMJUOj6KqbD34glS54b900dG7bRcGhn6kFPU5vmRE2owgeMWgWv
zLuPUayqEzQBqLkyg1SuTVx/NL8hHdjZNo77Cyo0PkuNLI0xdH5Y4Rzn8fUHYoVJOoIpKZgqqHx3
bpqSv+HYJpag/7WCsE6r2nNJ7wZ6NsHn1UW2tEtZbkvx5o2FpXYeKWgKjcvC1VPtWVXZ44JzgQKA
fea/gIN7l2rZ56O3/ehKCP8eLqdnz/TcTB58E2ACWF9XVpdKxKT3LGUWe7EHZBdPECesSZHUM1/s
ec6TrLB3wHS0vX4ee4S45odcIgm3tmBdwWZFA33PMEIK1fLSJBhcnCxWLoYO6J2MjVDVBd6ukf4V
/j1kqJm1TZNHsmcrO13TFNM0t1ybakFHEMi6io7c5PROFlB0DifF5p+0R7dJAx5fRKvETrJv1s2Q
2PGhxWjrlG4wDTaDIYsPMte/NmTSxWuZchXi2rRRLT8X1UzUhdcCH6A4ao+WoNqN7BJksszsThZH
UsgB5m0zSBRWfQX5V63+/+lAnXwYdVzjAC49NZXbageqy2Vz2kRnkp9obNwlXYCoIVOIUmaRdD9n
CoBtJmGtuJ6Ym+D0lJOHbQAqdygn2uVhM2QmDYft9HHlxeQQxk2WBtE9g6HRncV4I1A1iwK1DtWf
bkf2uOLsExOP6w/4r0EyDlJHhroch4ZSYzsbrqWFt0mQVXv6uL7xdlhI0pVydl387himXay6S3On
tU8o5np1g8wINhEauXqTQoMgMEobK7Pw9L8UW0GiF8RmHl9DqaQ5yunDfsFk0rDPSq4b/XOElwTC
FEGIvwxMaoVKmsUSsRCK+H9iA1IcvPPhjibW0DaxFRZGvIfW1aTm/cEQwpwoQBLynwwyqP6BUXKi
9gHTpwfXMnAqYw+6plQ6h9J0jhO6gUmEYVIlwGoMVTGOOc7W4JerrhQI5ub1t3lAHbXEyebmZwnr
OTUv3HrtyNBqgRE1lnjV2jDWCdolugZvrt7HqKuzy4gE0Nnfedk2z3Jqnz6R4A3u/ROX2yzaCHLi
ZCz3W0Bj8tlBoCiqeyudQBD63gROaLmEB5U4uYnlAD4oP0YEJgthAuD3tvaq5VJKpqWO7urBijYG
WITkZ38mQGxMCon9eQ6EwKHXrxDc+/Cxb3PxqGHqaHT8g8fDMKEx3NxEr3zsQr24EHfWdhpasPSZ
ILxmXeDau35+Rt1XBIaNXqDWaROZa5UTDjjQD2LArlFezmUi90vovhnXsl3c2lrrPTCvdv5OKIKa
gcUAskpRnYoCv3LZL4PKZHdnNTorNxSyFQhuqRveGDKb4YeU6bV4QqLGxRju9RgDr12aHRWDbuBn
hegKIx9K167k7jJ2pNTtcitVqCjzPZt7WdPioTPiJJjmriyVPqDpZmUAR2bGHlswa2pq/Az7M8rb
Am+VTkbLphKSJlFe37uLqNBR22EbLbtpXB2giST8sBMgXXteZw/C73dunIahuZ4M0Z3BjTEhxEYF
K45bqFX+60kDHdrNTl7t5FmOX31/zkRhVLQ5M9hugR48sQeiZUR7FC1ndS+6KZyDSPQzGUwh2Ftk
h0Gw4wgW6O+2txc5rFrh8h67cJXTxjxpy9CysCHtmNsl3/Y6xvEpz4qzeiyml5XLY+wRdHdQ+Y6L
YphCvnQrw35O4SGMPL2Flvk8TEmJqyWcXUyb175BxYc/80dbfbFCjv9JJACp5yePEPxIRg8J5xN+
b6CYV0LjoB/tX+zgSDLa76oD59itaW0UdfpC9Kanu23nwCuZktrgEenonJqNQPzYde78lnDLAFST
EKc9hSHeTMBvYp/6LbimrAIKJHyXIr3cVSpjd9PjGOFFeJM8oYd2x4UzulBbp3F+btJk9fxLukDv
yz1yzACmsnY8H0kB+FDz/a6NKep+eCEWhAM4D3WXlA+9KFK4UK8/9Uaer1vx1OfTFIm2FHZeK/ES
ie4v+vYOZel5orirpkSE1dKoxd2I9gUFUXvO0XL/Ub73ze9d1JhsmJt5jOUQoyeF+nJbwhlJyPCN
0yKtoZMJAwcZfzO96KRqRlY7/I/6Z4umzSIMRt5KUrRCM1CrvFp+7EvW6Khw9gkGuNSZwneh3DlY
uNen4k7IPzJ6rRLplxhlcfcZSZwmu3YbZnAouWlmakIiHX2xiok9s3iC8U4tJEkIBcMgekge1W3i
m+TpXfy80hwJPy6WMaX6IwPPinWl69eBBjirDROATz4oETWcHH1WOCsPuRB7t1g3KTuRyVtwnZ6O
Pa6yxaThfdIKJSu2rgxIknuukkrQ3+lufGeJYQB20+yEOpApj1EXoCKbopDp/I/txNKdyJaEXT8R
SJSNHbHFobEFs7c5b4eoUQAaFQ2IVhYfid351BKQORPdrQHNdzf9btl6fRxyzDgm7nATM2CQxw1U
HdclhdMV5+HorFqcKJT+6Elz7M8iW0O0CG203Whfv71Q1tXUd0SJ2O86pwK0Qj76zqmr5VhbsHNf
prLDj7a1hc6XUHUcUeoB+TKHLMqmeY+vEYPTE4MBUDz5qXeY/NCLzgYhAFRa9DFEoPlQWUbwnWce
rCHHqZS86bh0sC+SFJkuVIDMvnt0jDlUkx5I4bGJ6us7OLwB8SEePzmtxFYK7vejHh3uhg2Vn65u
S3+CsZ14a4Aoc5A/uKtCoIGirEbJvT+CdeO+A+49+DqHd1w3ZkIqgQqivE3QsVYVRrlaGunehOMQ
Y9H1DzYB/ZNzE7EV8kudY9rl02zDN9Wncf5cun+cinG2by6xdC86Ilq9O//cqKBRAe/FndYAe4hV
xpEcsFHkBftEJgGeF2GSILvYKHIIKhj1wSlbkdBfnd/hvwnGX23l3Blko4JNzSbkkgbSF/d2pkVj
+1/UNphG1Ism8cInE0T3hMpGXzTcRSUbAkCF1Y95XlnPxVZUEiIOfefkEhS0VCG56FNUPirZ3LsR
gAS4StgO9+c2tJY3AlFf8kqDfd1nYZ7Ih35aZeLHcMmfulYxQ6kECmL+mAL8Vj/fNspN1d6mAYuY
Qn1UZCMCrZljM/uFqxZPbMhPwth9UL3Ytvitjff4n7UuHvQSaXDAlBThrNvgQKucWi42hUmaRN3q
NEVa62yCF954Sxipr9iuX9mAwx9fnOXzX4k5Dh2D/vhxuoNaNFIhqTsU2esW/FvQPii3jYNU/rbq
qLaHmGyeMX81XqHdMO4ppPyURLSqi3TBMi4CQc9pJsVcrJbZR+a8KmcInHIJg3myTMBNDHdaFZjx
nIofTrG4/675SJQbxxI8+q8teeJJ3jcvjvWKPCDhYl+iAJsFf2NdPOL1gXsYShfNjp3ONDBtbuws
e49XhZR8IpDxZAyYKMH86Yz6kyt6S9B/MrbQEkrEyk11BR3t80NUZtBlYWt27Z4zAEy8woX6NL1O
DDPE9xxljaCkCxJOvley02krk0IAs3ua0cc5pkrrUCo4Vv529kzlhOuRghjSfV8MpwjJRzS1hO0N
9P/c/DYvFI1epdVt9XOD9+h3S2QyYakwHCr/IwaIM+ATm+4x8dtdUguZiwoql6HWJNiJY45Wu8P9
o13cztNkm59FXiRF9QlaQNDDmPCEKxasngxkbF3MRtHWX9wOafmkXR3L0dl+tOaMci/5hmCPOYej
my/eL1C7+El/jy68cpJL0HNu9sQDyRVIIThy1WCPjVFYd1XCR2KGfYjjbVGXQYVLkXcS9CnzQT5L
5WsUuNW/f/0wlX3OHkHhYRClBOSGmpIM9tIEdisaDTI48Q86+iBzHdrV9zvPdBZ+hoKdu5K6zg9U
gdZKkeaY3LqPiJxny1N114n6HhNHfQa/cmIJT1CWpWtTjH4kZS00li4Ej0qM8THWbpRjrxwP08hR
dlNRz9yvO5pp4OWwR62gOiC2kwqQNjVd9OmeNfKND2zXiAwqKHkAGrOT04CUB/cQr7eTF4s0EM3u
ajHvcGt3r8YAiGKlt67OOUAL1fxC9PYDF4yyC1ES/H7IxhuHchev9KnR4NQYs4wImgQUAXhprZ8V
nJI5bXDWoOZupvTVEakME8Y3LGA6yRRITy8EpSYdMRKxqnya1145l1egPTXT1zzGWaL97BgOvwtR
oVNd+6I+6cnRklKQ0qgpB6C/rJzSC3Ir7Qs9sT+VTx8Jol3hysXKvDiMOU1Cz7Rl5tst0Fs9IJeQ
WF1cohNP0iRbj/MI/R4k+O8usMIhq5GqilktbVhgG8wDaHz+xN2nkgADXjJQXSnsD+/g2n3WLIop
eeVZAFHGmN8MAH6mqGvUrgPoNa6frrezUAgSxiLljx1VvoJUt5m32INQqISV3Iy5bqEBLGZPZU1T
TH7xhOVjO+1ipNVx/41/ZvhLW9H6zL9iLLlm4oWePBTe2cYJNEy4OuIArfDqCbRPY/T8A8/MqKzm
k/A/3g2dUfgkNg1iYM/sgE0N+ta3Ck0FxxUVCTshKzAK1vF4SFtx0ixoUJk1cP5LIwZt9oVnjRak
iqRVDPd3nDjfKRdOBDQkeaBEbNxny9GAx8bEPg2SJyZkCJSksosbQLyFEhsE5AC9kXt6YHyxR8y4
n3vrh4SVb28UsW0EOEPkR4vaB+FimaR4dSjWuUj7qGH1wEtUKKCWK2+zDCQTVAXcQPFy8QMuuTcv
ghqMxtnyFOerjqGiiSalA+n+00ZepriGnJdZypsS/tt8OIFs7Wm8yG5D0bec3D6UC8iQ6U+4gGPq
+v6lACGY0L4S8wqLesInhBzCuwxZlj1HXJbBuy4D3A35pScrlZohSgvukt52MyGqX7VUDt5QRWBN
HEsg7H5LK9B/dX2fOJ/SlZ/7eBUkELth2nOjy1t4Q+/P/zMg2vI/UknLsNIGlMa6CjIHZ/S+VCA6
T6qozEVoj8tsLAyOH4H1h+fe4d1KahI5a9x4RDE3U94kzMDu4uTpij0Pro9yifBVinDnDsfadvM0
eXy0uKfDcMi4dSUdud+5nSAeeujCfgYdT3GMg2gMoOKVGAqYn8QId0e/leifgXICompGEw4cZjhI
0xAgM5CUOz5MZCvrL3mQWmlZ592fChI9mVGdS4z2NCVLpKmiVoDCYnR4sTSlOURx7mGdlXZCRhqk
BTqdVDQnH2Ak9bpJTVjOQ1EbicOkLII56Y51iriCbOVcqBb4Cb4P+SPWN0gweqK90JtytUXvQGLl
TJfiCyMyVIz1rFn2JRLmW4aVBhc4ddNw0+XcOWkNs0eGIU2urPSi2pe6vnw6WuNRHSxw5r1aZ+VA
wit76KbsrGi5H0NLQ8StLdVQXFDm45IDVKh7idIR+1ZtGIa+UPRtvHcKQ0Y+xEtnviutpeWA/qAM
a/W+TKz95K8ji4W0P0b6yswASvZeCTRcgxXix5FmwWpIjo/nrJ41Jn+hchsn1AISmpHdzY6ostUa
+8aNYeYS9p9zdFJnZ7kg+IXhei+n/1s3vHqk2CTpoP1j7HS2kgH2DLJPdxGOYKJ1zTTCCfqGSd0P
CUukMm+AaDhg0DsL7irN5Y9iVhqn4sGx26e8F2+8M2NCH1AyWUWZtLiTmQgzU4G4PqtAgIpAt644
zL2u+IAYCsjH/QOBteV5QydMVlFAl8YvokYJY9OqiOaIzvPVWuxmQsBKBoY+G18bsrbAGKQc/XMo
JaNeDlNAG90bkYSXuHJKQclwgtjqcUdcPKvqjZ9FFwgFuFgoneSb01joguZ/n6bSGIhz9HCnI4dw
yDlSzuLo9+8XivawXEByt5vuCiyiFSeTqIZF3GzJYp3r91M5con/UHD+cVHN5qYKX64PLTroUyrV
Lkg16t33FGpxCXDyqbm8+RgFXz1/VRj4ajvX/uAUYJqxvmSopakJ+ORN2IXcXLhE+0LJD81BEIIK
o4SegUBtr6XC5rsvVET5mHmgfFKU5t8k4tPo8t/iDO4UaeK2pqQ0eIQI+2AU5Nj4rLZ7lOHYzAOa
GpzJfYWrAAl5n2bk0lVrBBYjAVKRFL7r++KIWdfBTqv3257CXiQ7f3yWsH+GWgOuAtIPKOO19zVR
4Tdy2qX/4E0f/bxTM4deBAgmRpPF/AnW7ssHUuuTJDPAxRMtD27H6jMMDIj8imrEe7GvwjYUa58n
wx2pgXBbi4zyihwIouG/vMxHVB6+P6y9AFsp5Od99VhqY5NO6jDLUuBt67Nlq16UVjWtlX4TZmXQ
T0KxT8s9csiDKbdcSGO7xI2M0MCLbWunN1PouStsUr8d/uzhAArurJTC88EF7+V1i5xRCTqWl5dJ
8EBc5NdYtd+hQsLiWF+6X2kadjZHYFs23hy6hwxw77dJzKIPJLmnTt2TLcYEDtPJunPqpsR+8zLQ
JU+maDsmh5ZzqcSnpS4l3eBxbXUEwoGEOgmjkITstNJqEkEYGRJRTMGW3Zw3RcAvWBwxy6wE2Wzy
DmLDNOa0TYFsW0AIDhT0iZrBFRXF7fhQnm9wfWMGraAFmUZrGnmy6txtgwsS1nk+iyoq9frATTSE
2utkaGFXQa0oBje9lk/mYbIcbfZH8+7JXa1yQQ6VFEB3bjZPhWSLLewzvOnqOXk8qp77xzoyCJtL
pi4Rhe2KQfxfeNHS9Rc1Z1JWCel0pIp4I4jWIVP6SPNhxyDJWaaSh55Zm0XZtTSnqF+QYkJ0Uu8L
vOPwB5B7C/AuAaqMHOfLIwNNUBQesQSWAQHsNq/ai8hDwOPyo1w7esOc288BSf2EirUdzaE4GKYj
Sa3T6JEpLHYRuZEasWmQhL1rAmUfLNPXptt1GA6ckliqIW0PjEZ0RVYkKF5m64YceSttD1fIY2Gm
lUEOqi7kxVRKUN/Qix1IT8xmf0MtlGiEF4YLEI7ajR3YssluqxAoAune54poTum+cfxh04jXq8/z
04dnrM4UTsJawKvbXhprjxmEfd3/CPw2QDLS0cywABWyqe9+0gdq3jcvaG9IJTLnao8kB1JOgCMU
PAnuXLMvTCRW2pYKH4ZH6vBzrM+7Zlego8FjUH4RAa7qbig1i+AdrOKclwC1FMrLRqRjetf7mkBQ
5CrcQnUv0kD2Osqbas9A5JqoKmSdu1kAkYXyem8FblKjugUFnfQryvibOYPqadQcqJIMYZSXe91X
z6vDqS4c8vC2KE2nzKf5FycpgORfodVGoIw67CFovHARES0kTlWAP7QaMUtXynjo32v8DlAvM3zX
OxfkFG3wTMvjMIS+1v3hgd1aUzNAdsUiC9hQJgffz/e1p7wIemabCTKM4xJhTv2c74FiZJdilEqn
GY+RkcAIcaSvWJlh0RuutrQ1MQk+IWTRixdYfN3TG9IWGYFLcMDyx1FMIzPP0Smo1/dg5fGZWhyK
xj/eGKZAsE7ddi8NpNO+d1DBwA9wPqXaVd4TQcEawd2QBUK/je0Ihva1koNY0mxPsA9b3ghclORu
oPCxvwekiKR48ZBNJN1VOD5JKSbi8RwB3oHXhcuRuiNuD0EdbhFsrIGSuMvvTh8l1cDkUzgIVNIl
SnrgySVW/p3O8R/eYi7SpkxC4YxpFYkiM3UvliI+ANi1CewV7hjRbSHedWKDzthjgFBfx1V65vXI
6t7d+nwNGCa27baG1tegzBwP0blf74t1zDWcDZJkqHpE3LbJmD1eTC9Reqy/yORs7EBUBRVGEu9i
Tk0w8XZ7lykzHbeiN2YB9cXe9peCAIxYi3imhfSLlcOsDTjzPBZrhnPLN7FqdId/fom0fuOsMr9u
s2Z4pTcqALuKKAatffy0wggpnLrFxk27qNkV2PtZSy0vQPOAYv3GqWZpm3zQQ1iXGPurnOE41yyj
MhrfCtvOKsckkT2HMzmRIw5C4tQPkXPnqUjw3vVkL2okrae8rAEioyTdTgYSZviHk3w9up0wzgwM
vTpYMA5qPVeKtD8WDFWQLMG761gfXxuQIfZ2ON7K4aHr/G7WJZ2Tl49fS3OaCxjblKEX1Vsz2wT0
HMqq7BpAvzruwUCTvd9VDlky3U7h0BwiB9bq5/Hr4wVGdwA5+SdCiUt5y0RdAmQCoTQX87eUQZlB
Vqljvo7PLKXG3BRERZpxu+C1bbnKRREJl/3UpQgDIFlI9i5OGNCsQ9lhAJybhrpaXWvu3bEqO/Xx
sE2VVyYnXWYETWpDYLWoKyS6WJCJyGSITvNngcI4/vs0G6VGz4x94k4CYT/5SWr5Tn8MzBHTLy90
+eXdZrMnBtz6jBm+dsUWm+EMPMv/jTeOV9ehsjLuncESJtQbs2enULONEqiH+XAkXRh4e83v02oo
kpjEyQx+YOCP/eTUT9Kk7hAxs7+bWiq4mTATaB3Epw/rnm3+vBQvpejx52oICoAj/bhp8ggqFrik
KDlH6b+1IoQ475hC4Ky9nOtdwCn3mpfztpbDgZSk9GEJCgJrLK5tYUhLA+ZmQj/n9GzFjR7Y1yEP
3oT32NcP/T+LcIbE6aOSXavqC2edbS0FupzT5oJHzZEKdq2S4+r4mrpIG3q+URVOorU6CKrRrniL
IEXzuINAAppyW2nZxr/cRnYnC/KWRbEDaTN0F9xQPp5juF8EHnSRReCxKUF0yzNBzlnU3LdJykpR
m9k7/N7wz2mLQb7+Z601BnNG9d8bECEKbclg0f2N+dTYUiXzey166NrJnhR/GRkBOeRL4KCdwnTG
EYwW9fC2HTV17CXYA4gpCKW9D8E2rx55WjjFNLilqUu+NLz20Lq6VEp3oA2kPArm8JmxKdge85eg
cI2QZ/1pxW3NNBf8azAq9Brfw58Wbxgymbo/HBXvonG+nYHAYkUjbmSZyF8BasaqySDOKAMvYL3i
RVkOYTtGqxHIPHiZT6CKYLdgou0cS4dFR0e3IXuzUgosDANt5sOeI3ZLjDknpF6HBilPDPUDQlML
gXDA6AquLOhBBjzU+kVuB7sFtbVknYgSSsJuJyNPAa1CK+xPgv/c10NPqnxMBVZnCs+JM0f0YB8N
w71twMaCltZj5MjTAcEU3097tAQEGfQR1tUCKF+xzr1iDOtPGbaaEZjfbR2Qht7jkQlhrCB3ZJ7Z
yI6ysu/yDOMmHkG6hIn/F583FqAf+H7iyQEsTtPVnxtumyarvz22q7RdSCFwATIPR/YXL7XeGk7t
sIpQcUCxlO7P+BSkfV8G2b/dqwrHZe1n8AFDlwG5JymSwuKZ0dNprDec0RycUqo/lfd6XTkSPRd7
nDkXiDuzhtVEDlT4/MnNR3NLbuXoQRLzEOM3TGmYAzwm4OGoWpNdw2hbakNynQ6So6yRIUZ5WHGQ
br585hoh8fVW3KA4BN1SXSFkGm72NNJMNuqmEgKgewsdIY8l75r8Q/RHwubyimyRv3zS3sJ5sDRP
mF750lqJ2qu/XHNzyeqTXTr1vmuPrNEUNMKF4FLpRTYwrhAvYVJxZj3OIX9Mk9pklZn2yaAIfHHa
UNkLD1a7ikRkhWPxPfNwo1mcLG5Ya1tSISb9OXGL6X9HzVKrTZPGipkDr26Iq4Bka40fahfARENn
zoNnnQ7vbo0jSnSgLVOlbh1oweyfw+fC37T4dJrBlyFulkcV4+V3aAuJKOFQhw8FSnclIL1A5EDU
Zu4uWQ76miVRtgsnHyNZSa1bbqTdNceRXXSBWiUmJQB6zPHdpafgYF0IoDq0JUDu9wj95h9KMAEP
m9fmz7W8YANakdH+7aFGgO+n/AQH543HZfnb1WBDqf2FB4g2kRBvKjDGLGlqtuywQWLfroJUh+1k
qxxsQa6H8OUm2fSkD+VxcLJ6cCzuft3NlEUxgbOhc3AOt+Z2RAXKDiUjq1eyKnsmb6vYcCBBkh7e
syHM6G55ycNU/DRozApGbupUJ2m+RuBFPMC1NVfZLi4zFduF47QwtR5+XiPzxNsrUX82oLRozXGO
RpLh1LDjwArYma5sXzj7/PsE/3mltpm/mapQ5prTovoqMV+XedTSsb3nzwx3gIuyV1ZpPWDmkO81
IE+AArvWPchBTIOSjB2/WYD5NIii8ZQR9cuz6PkmNxmmJYUAVidoL/hkZkM4yoyzgFja25bBsPRl
vmm22WEtC5sQl0wy0vpBv8BbMXVwfIPMvc8Xgk42Ke34cZfbMrr4eLpj3OqgJEvxurKR/Tf+NYAf
uRw+9ijf4bWb3V1S9NPaGrcxmceYCRoG7xPL64v9fgt31gQHyWKoAPpbE7UKFkSINhiG7vtmStSj
ctBiYEPYYYGrAdAncknabbXC0xe6XvDncp0DP/cce5ErtKWOxWjCzU9BoZXsl46ao9kNi/m/WAmA
foWwy92E2CFxs3+v6C67X0miYzPMML50W6zu2smf+2qh3fESEwpY0WK+UNGCChxU+LicscbRfw4c
IT7EB+071ALPPso6ZKVokBMUk7JvoW1RYHor/vidwiwuAlOvFI/fZ6a7nzCU2UwpEYfXVL9OP/UW
NVWv0gZOj++5fAjJeKZHojZtjO1puteldo+850NVxTgwqt5KNhYHE47Cu/hCQF4nvwf0D2vj5POJ
ioCBQrflHB/LbGiEKgixdkHmVQdy26fj91oE5nU6DC+E9BLlFI0lbx9Eecpfq9PCeluy0c6yxXvR
2RJFQovHGeA6Br6WFsBJbItlUcu4ZFtSAR7/Y4u/2aLxxYayuYBz2HVY6xOzbVJAzeVz62wX/RUj
YWnh7j6FiS4cUYboWORmKTgZKeyBZcKjmjlxvx4ZfH1FwRheZ71/9bSj7+ZZQHzSWajXWe+loUpY
WNOtpjYPJaOrtRBArLk4F5X59u8VVBMe6FBDxUy1iU6fOjLde3Shn8FVoFL9y70aW9OJ9UAqNu+o
P7M1rK64ZPY7Lm9iM8yNPdtYKL3ks2x8YBsHHD24Q+siacKhl+835vN65lTj+d4tJKsC2Q+gBxV5
L2bByNTJt/wTsliQ/IVTWQRLms0/wtlpINZLnLaM3NqsCXRJJI54Q8kf9n4YddBJlF+pkoNLdiET
qKg5BnvJZuEy1jE4dgW0irEAuqeZxIAK+v9ScHmgbObytzZZS5TS3lzquCKVZR667ROrxx9vmHnZ
rCP//1yIAlZXgSBGbNTfyoyqT4+lkAfUWttXGOZ52QgaG0sSx4KEKX0athsI4Uu3a2N3rhlUDJHp
4Z4ORdirKMPXSon22z/3/RWk6NR2+zzHhsYv9jd9kle9TGzMYSMn/3mEz7i32NL0OsUR1KF7oGve
+rlmIdGcqOd+z93uEX5tEzuLahrAHz07q9ixvgDCLLFYsWijLaHaNJ83OpwJHNfN/iC7VHfpAJtY
SZkMKvEeQsVXen2BoGci4uZ/uRlF63rVwHLX+VzbhNpM8aclc/p45DiyKo3vpeBKKGZY19pwZUJp
piFhSz4UL3Rj3/kdZ+cvi6uzBIroJDas/tz/rGgc0ht/Ahlnw02XfnBlNFpgswHl4ipMOJa0gUMY
Y9jV7xEUxPCsZMax9OfgMy6DPCdjz3etahK4n+0SNaZnYTj8BfjTWjd55Yyz5NJw5rdpKaJtMJFw
KtUtInDALkdqLbU4HqGVwwNkY7CtqeZM3Q1GF4NbxUeQesNVSQbkCIJMdQdXIiLyE4Qd6hBTj+gR
q0Sbm2oXXx6f3nf7C82knIXk84Wy+cejtgwZDyD6cJ1EtQB3+gS15AWITFyRgA2X3Uclio5yDaZl
j2CS8z0PKRd/RkvHDGyXvxJmvGpogj0ZhadDokyXMNYxdOAtXrbJTZ8ATZxiIBE+VZKvzyUZWt77
R+6HlQXLPYKS0TBK/uJsyStu/blAZqqRPg59Nv9OxWbYfNLOILwv1NOn4r7E9sP80MX7Gb82dfEq
FQoz976yzTvorn05o6vb3XQLWgfCzbYQ8eEWNu+Xhs1Z5UOJSTpk09kSPY/8KAOQIiT6bd9U9aFi
1N+Cf/AnrXwtVCgzF79XyZw722a4YgtReb0Uz/xNfsSfstP9uBbYTXeQTivT72+0Ll9Jkmyp8MZS
KT1vJXxELq21++cnNqL8E2uBsTx76VKgmUqGp18eD0eTyg7G9FQZ1yXF7zS+UzhpvT1l4q5fWudL
OD31C3nmHpGfXIRHLWvqNwsdBuYeq99l6O0701XW6gqC3cX37aHkrGs3GkdEMUtnLqkgUKk7H7m0
+/gq/x2ceL5xU+0mxUxIczT5hffIo+rpSac2L9aumP7gSEOa7N9NQcZKltKS3uAHJqEnUsETb3z6
y3H1ww2fhM75jwDsFn/3b+4+QARDtBM/RUXu4LpJRmel3CA8fJzT0k1sCw2gqo4Q3gqE1nP4rybt
e1Kxxyxx3rUQhCUw75qJ3KYvfSVQod5TDdyHw7FJhZi6Xp3t2YHfz8XSf6wcyukh3LtRuOc4FdpI
NSJdOYW4M++V/WpBV5t7pxBW3PiaOKKnbspwwN78VZ2PwKrGKuztdge+w5TQ773/5yN9n/py2dFD
jRQi5sn06KKGEm+yjAgS7j/orLY0ROPESdGrN9w1+IltH31jiq8omDP4i3BV/72wWT0SBTzks8dl
4/l4qEA7cIuibwCKtwZ/atkYnJOWcGOBwHBFh7TfbtmWCPVHNxcXYUs8wRZ0N91i5ePRrYPQKZZi
I50n+i+WHhSov+7PmSrmeQTOhn+L5XGA6DdYdyZfL8/nnQAlfQZ8fsCAkq/wlcbNllqvNn99Eo3t
iLyXY6jWrrH9FdOl6KusrLrJ9BffGGqLr/ShpvdSAOeaNbmU3LN8DVH+dfIi3wfOW4naCp+txXTZ
8AG1a7AyMoFiszj+jdJDlH7jBdp/R/JLs8aWl5T0J9UCCiMaxE1c5TK3tzuTjm74AfKZ8dOSTyIg
JtF2TUseh0zuYpR/AbmSDg4cJqzyAzvlq2Czu7jBwhMUA4xunvfGPQqvmr8AuJzijD2R38izVi0r
ywg83YyxMKdnUAkTUqNmPgksNnuzxBXjwhJ8QLDiqhvHQZ7wevREVO0LDRhht7QLg7Qik1f3x3ke
Cp56n/m95+FGAeUBVeo5z4bFZsdTxZQfXxV/urPg0OOqu2A27bvmLg4uVWUAAdsT9EQmnMQ5X8+b
U/Q+1VY2QR2uX5XW6xfmdNeZRTepwez7qezWIIvdCNYsVhRrV5hFeXigmdxlCZfycvA4XrnYrDA7
qJEQw17guqJGo9zkMGaAymVNdMAH2MXjkT8b96ijPfUvMKGoiT3kIexpB6QUeLExg6MgGa0uygF/
7UiJlxDQeQZWMXmopjS4U2q+rQiwd6qWmpFhXLx1AJk2zLpChcfEGn6vGzozKHihkg1sP566ckk5
fAAyPSIcfY4e+NHpPdoyN1WQMnUvsfDKvSLsZul+oEufuZvUFiDCDZ3j85xyNeMwtBrL1/OI8FFe
0mXfKweeBcigNHEW3VF5bKw0wu8pREjCMdGfQ1O3LN8AILKyMyWu/aGtM+qAy7reLlMr4Gw5XSj2
S6zLxUujJK+ANZhhktAY6Y9XL/TdZ91UFCNegJnYh6EHncOqOl3faKYIeYTKegoBrMp5HTGNTOzM
a347A8jv86CUS8eVEimGJ+lyhrTq8/npOQaahht93RdCtunMCP1fAI7/8p58QIDFGKNn51nS02mj
LCuM6N4N+rSGPusq/K5/pFkCJSxYCbGprlBvxIS3WfBq/0pUVSufVJ2iysYu94hkUIqLURc9dmm3
aTmJicGL7uASbZgF07V8ZqYbxe2EWfXSKs5lGwb97Ij/MVl9xrOVs86a+OeNgi03gqQWnGq19vB+
ocJFElVWUXe0B+eDYeBQTWa5tQGPyhne9sY7gvuba9Dqo+flEspcxyUlyuk70AVsaEKdtoIHdGZl
TnSL69eU73mjsWFAXfONaebIZSnxg0wjLpL83HMs6H4awagYn0fi/mtHtuALInOgRsA+7DTGDP+c
8jBXWbmnTa0A8n+ulNQmXiezQBYPrn4h/hSZu7nXgeToMDNrROLWtsw2g2gjhNS26ZVfR2tn7bOq
MWNjFyJAtfJToD27cCswtolWwp2eJJM1vWXbGPN8hvKeuTrKyzDwcemXw+9J4tp0DUX53w69vyiW
Fnpj6q2/zOvWZFi5dDYyQhcfH6GA63h9YMA91LepbDqKIFZJ3thpR+967HAgpHq6FKNe+OWN8TnJ
qMxX+OP2t+U4R8NmeePMjn2YybDcABUmWOnB/oWGrjiHMKoyFRNtTqxNNaqtbQjiWvG6AhGovUAR
ebS33xgjcAlf6HXifX/FQkiAWUaAw+69JA1cY+oeluxHa+mhxfe7hruu5/yLCNX7W6R0F0aA5u6Z
ERRLF+nEkWMU0Qet/JOVG+64DcIKFa/LetFtNFZFh+kE3VAKrulV0nH7MO+nOV1Z9cjSm+uFNTx8
cTKby+Lc7q8/bxUw7DGQsb3HMxPyJalgjUJpxNbF9cbsXpSOz786qDKriUoKgMoJLLkeVOhx7Jho
2NNzvB5L+cvJHlY7MmMBAAbEJiS1Cr1bJslTQAuCGzU7QzF0L2ppfzXbk6W191FcrLu1ASCj0VdE
2DW0oS9OmSMVBWWzKUTBqIt9sIEByQcFkS1xYAcans9LGni+V8Q9sAAm2UHZSryFL0bGGOAxL6pH
jx4gfeCXPDCDJbPM8l5wgbvHyd08JWA86AmEAmboTTf7vWkGTx5sccXNss2OpUbe3Sz5rRjLYCDF
YGOj4skGq76pZ5YB4k5y2EKIZkBq6utqoTrqekD/S3Q1PTdNjz7Mlbn/9WM1c+Kb95MEcYNZEkZX
nwjr1t8nBorUoWgZek49HwLTiubuozHxIGDZqfR0MnilKHTkJ9lnO4dVhaasqTVsWbSbryJFLAFa
CDuyvA30Dq0/B2hgiI0ywKVVe9o+50yWU4ohdLINkD91oBI+AAgPlp1QsacrMnHSq2PmxjFXCIeg
Zh6YjBqCwcp4iNZezDVbpvFbOGPV8B3RwEacAqKCyWuaI9H9tD3roIm7Wuer6e03hF0Rb349id5X
/daj+KeIHfLhTN3AjQaCZyytRig7rv5MmAZrl2dCipKWWQVPi/w+uSAiX78fO2fOox6BZCe4oVmA
fVNM1RAzhgnuLscNvYrlmRC3Mrw9BkMyMO4nBWp2BIRYCvMS4Qjj9nPCiKVmgQjNX7WMdoL6kOFu
HRw7oYviMBD6kWAkU/wB6eyxRr8arYeY0tomwLuhxRZg5ckP4h3UjlmsZq8wUYoPQZSLc2+/rYUP
A4SG5zT7PX8MNwHO7vozw/Ysy1XfKwWafRGzmTM85LDfI0A+r0vB/Zg7IPqPrWl6cv3jPG0YX/47
dvIrqmXIiGMx0zfR9CYCXQFMIjZ7R+D/vAr/ge10jbsuJk07tme4fSC2nbdORC3DbPmEwCKPQLox
8zYWWFHHQeAymc3CfVInZ9dEJrLjfcb/PFnjGEj6jai0CDzXXEQOhIY/YVecbyBUydSfrKGcsgPL
di/1umedmTqvRTKOjVbsULENfyep4caSpVEMuLKqcB7ZBmTMc50TQshDUYjjAnbkh5/2fwD2U9oA
A4v7HAXHVlhbhxxmwdHUrh9DpMB2Y91qPtUk9BobcMdvdgv2phjU+GbjjmvPfkHn/HtxBRN67XB6
zZFkjPAR8OWTQteLY8xBIHAS6AKh50MQDgmUVCAvSv7+mI1nKhLFYoHtv4nGaxTaL4RErMSMd11N
F6YhDmf2OX2cZJ+0JmE4SodYCASUA8w9HPVdq0DPXW5ByNM/X56BvYBgr5s77kcx9H3wn+5wi2YN
vkFhKh8YilXJAfatM93Tf39hMtgBfTxhhcuPHgdJcbmaZlVm4kUgf+i2KvEcbWlOWN2bTjVwiHYs
UxIy+63UbYHWsIb0zPY7j388APrmmBl47lxadI9M905TewuN5UqRhsD7pm4eotl3/M8Ua/In09Du
iguVQ/ca8+O40L2tmMWpIKk4uspVzKy8UXJJWeIafpWAk9KImC+yPG00p/C54O6SkCE7HhcsJmLe
ssxGCBzMw1EPhggxETGdr+hN/+Qs9ObjxNdU8OMHnKtl7YDYUIk6UiA6ORCy9o8w/y/GIXavP+t0
SyFgHhb+vQ4wG3VosU5JV21osIz+dMsi51PnBdmAhc086E+Y5a+tXoPXKTsNPsRZwJB0vmTbSTsn
TdtTGS/vT9PoLIuxP8Vjdbe1pAdXgUTR7rSVEcL3GcMVJmlNB0+WEZqntDE8FuFtE65MbwzBOEmE
Z9/2MKHVMpBa8kOtOveUUDZTwieS0QROy9tt0fCWO2GYCWx/ZJw9iX8fIN7sGzN6lPasd5eay4Ce
JM50h1Ps5cPVtpzoy7OkkJTvmBFB+l60iE9XhIvX35e9hvxAICj44AIrWS7bEKFYgsYzrPJ2LjCr
+mMhvYyh4XHhu74v92jyWuBGXLs++gGfEi96U5c8vfGAGt1R1hScVt8tdzF6hHD//t7/0wQqwsjO
40eAu3CAWP7+cLSFjH4A0YqawrTTUc5Yk+jNV5EbvlDqJro/6l61fkUd/8SPLitqwsWRApybQ7fr
qTR7qtBYp1abv0uWC9cvpViW1mQyUmPmY2hxyqteAvzY5FQfX5khNZ0msf+M/giGCFKfWhIbI7Gg
7ZGHHAsAjp/i61pDM8WU10Yd7C8fNFXcF7sIaUb6vpUZ8oEEAU8dg+v06KCmEf6W/mkSUa5sbPG3
aXB4ZKX/XMLBtkX3XRQJIS5tVzYpJCdgKXw6jieXgvkjWkAwD0thaUD5pE0btLiGjXcf0bvAfN0l
DIAOGtUnKpai9/CLVoXg52wvwP2gcqzbnH/TXlOMYN701vUlTxP+RKKGisSSEz3z81KL0VBw2dmn
Y2UnaLFl3kgeBUtP/EL6lSRJv6ElCGB5SFPuiLiraXYCXQNDmHVEKv2WzdJKxvRqsC23gUwvAdbA
VbB3WpH69qGAyt1IFIVnQdWnqbQEf8+pxbNQQa6zRwVr87v74f4NXpSYqvYIFDrg3E8XtgYY0Vd4
UDtACRtQQxFq0Txuu7xB+45tPPkHVrvptV6NPFZjS3gDE95tLc9WlLJHNIqNgIBl/6/ZbgLl3Cqi
3bwlQ5/XH07zOZGFGNLJ6QLmh5Rqg0kbFGx8DVHEDQItoNC9ICQ9SPGl17KnZEStD0mEDC1t6hdQ
7e8LWgd86T3pzCTlbm0JtKyDl550MrijmbmEw9DeX8ebOciJMTXsEIS/6SVIQOnjjAZFBZWtJ3Df
fgTmSMUm4mHRzM3j7XL1+FN6j7KI65o4UQRYnnXfrcOoZgKwZ4PJRBCdjKsMy5/sCsY1cTXSiYvc
iFigu+BI2WXJyAL2O3wjx6lizbaP7l9OF0IFz69em82+puceXKYoNK5bxuWmzWKWfMLUdZ10qcOg
CGwYvtlWYRZgTC4BU688y1NdTx7oCyWtVToyoN0aIeR51y98npY/geiEd6RO7JCmZ4XlZVaWCyR6
unaQ2uVGJ1Vys2s/A5MbLF0k0ygcUy4wA//mnxYkM0P5aDHF38HurMcB/RtAiFtVprH/CMaqAjLx
fbdXTzdJx16EFz/4Ku6/Peu09uYzsJ+s1y4DyBgKbGzHzeXjc/1ohDkpOdO+WCixrfWDElmWOSiP
Kzs3AgGoKCpBW2/fiOOEfhiufw3jeF5BkkptiRJPcVF/7eGcip/HHG8dtCPJ6UN1qwxRwXDU6kCc
cj5vedGV6v/6RMXSSWVaavDip2TyzoT3tdYFVQCnAUMs72aLfM8tYF2zT8Z77TnisfnPGONHyOYX
cxLmM/Xh6vrc2reGJjCf7XxP8MmcQLCkxQhaOuvNdv6EWzOHeWukQg+XjV7eVYEKW+zzdnWzHRNk
zLRZ0EAb3ag2w/Jsxyn3UzOjH2F0FX0oa9p8I3ZObAJ5gnBYPPirvb+jGX0yj6MxtxXKIpYEpkos
48sA+dObsLdfPvDLVNxUE0TMll1/41jMBqt8b4OJz5u324olS8uJK5j6x+sbKrogixsfjZ6UQJVj
6itT2UBUD9OAe6YDt4esitKX2k/QbKg5YXEZKie3sfD5MB0xezuRNj5Gj7z6EEV9Hi4MTZGjg3gx
t9kYOG0x02F6hF1322F3Q6wSdksRdk/UZKuqdC+Zu5YSXskT/S8wdMizW90j/y0m45WWn5CRH+ns
t/iFTXw4eduWWlog5Qq2ONcQUPCqQHvMwix65wXLPHVSU3FG1ofMlHaBhR+NWiChZMCQf5qpfU1l
uUskR0sSIjAabgd9XUK0snU76Obztu7WReaK68uxM3tuS0wiTpRwAmJwXIwjVh52JXW/TYGyxT+W
+oKvQmyLYe6thmFzR8KSKix+IcYnPeiUMo2N6v9YAWlvK7L4N2d6GLCG+WpMP67MV76Mh1MYubw3
jb1ww09BAUIV7CzWXWg9QZP/PXx8si928m4mnaMvN/Ng6fUZgAVJkN+IcEMybAKk97NGAQIcCoWk
N+XO+rMXOiO44P8QKLeGqQBRTtsKsL4HrMmynAvdyzwJr/dkG42wTHtxTR1B5yNH6RMU4oEh35VF
Fymh+hqkYovQ8K3eYPhGu0HMWn4M/LkJAsHl4w8tpn3ImOtYcsMhG0+Ly/mnm0sbsa8+w+I1E660
Ure8pV2OiyDJWmNX5NxB35ctwugy/Vmetgl1kT8Ccc8NVkTQLJToiAW9dz8o1SSA1qwQG2Vy+JPd
lTf+cUV7Z5Susc53A9Hs0945D7Ttp6CWFLWYeWDA3cwmZURf9D0M1sLZbjyiONgD47xvxGKCNnvb
tfxgwPiZvofSNJUXpx5+2dWOJzmCpCQ+2qhLyvR3XO4Uj/5IuPwhE/dtc2/nQC9LS3NiaGpTYqBx
QyXKQL4KDLxdJPZ7C58+ADbBKDbRDq41rvBjrhN7tKbaZGwNzAoXcteAJf66UYHi4M9CmbcE8nnt
eKJ0PzWwRB2itxTPyckrZPx6VVzeiMpktx5Ay4fFB4PdXT9dyeTO3kzSMGrUXm8ugW42bbJRmv7z
UxBCrh3zHQc9AaeH47y3H9Oh3fW5ZHhaWtGB+bveP45QyxVL1aTS2n8aYnHnMzTkUO8lzCtRAmL6
M+U0vYrQ2/0sDw4hRbLxwa0a4XQwrEel0DxFi0DhGbXMNAhX1qYTLv2DOSdYYZtSurZlIax/hw74
jeLdXft/6sBdrADnRwGYhsA1h7ZpFyKBoXNVREFNDS0YFEYr97f6ggbCWasuRtldLQhQ4R22U5DV
+HGC14ueo9b8O6n1xAvz2d9OWpSeDcjPQwgQKTN4TCX2kkGkgHOkK5LofXKvClAW/cqciYTgBvMr
cLAXri/x2cNgwk6LEkUsvZYPws1zn9pIziSbbD/letYS1fCB9pjTuM1nGWpSSDlGef1UTEkHxp4U
Xa8Dm4LhtdbdjcrdeDTV59BspsQgYay4VqILR3Ezx7lKeOC0gsBp/DT1c0Hv/aRmU5t8F0ogZwT9
Z+zn8KfDaCaVxmjZAOH7RctlZ8s2c+fuoDKEAjfxMtwnwFByfXjVILJxIkqd93BB153yC/cbJQQ2
SCsrTlU24svE+3i30JEoqOYXcbhoxmkdyZwoiqgBeYaPchRK7eagUVFH+IFaxjLqmaA/cyxv90Y3
2bjASDVntj9Yn/OjJL3wEJS9cAiwagaK7K3eSyfqTUwfCZuu+JuWDNwOu3nfboR37AdFnevkYPOb
kXeZxu2otNcrNuLZBFvS9bDVBluZTtQ7JHsn2SxrzY+tKoQqyipvVMxF1TCGCy8eJ/DM52ykoqQ7
8p9/M7Sc7FeRNnzUYCd5RLwmTmqPGYFqFR7enN05VjwnJDSB3EseOWVe1eMypd/wKQh+OfNoTppK
/HYTdzFvmDQKNMI6t+zWpojU7ksrCK9zBKI9LRwW7/SCD+j4+06WyLGhgiZeRXgBZI0TfOQZsPAE
Q0acAPhYw5UAgBkeQMHitEl9qc7VSLOAoiU2wgN3EgSQBSjvrB9h6kiJEdbSZzvFeGvBKzOo8kKc
/LjeQm8t60IHNuiCg7Rm2avb89/4EjPvNPr2ouSNcQF2NtL1KBCyaMqOWNsLzycvRG6budJuJm0G
ipKWA7fk1Xx9pvWzBtY0QeCrcMB7rwqZmIIRmRYG1CvOdVJPbp1kEh7+W8Oqmq9IK75F91UQKKbB
dTtLHcesvDyDks1rlsmIuTsinrl20nz0/pveJWWkreRYInmseMgnjoHsYH/C+4D+L7i8y+FQ+Wu1
fpfZZ50LgClTCN/FkLNK16N9uUP6Q1Lna24VrdhbvZix4pBlTeO++D5V3T6EImbQGbsPsgnSn7qy
3lJTYUZwoBVeSIOAbgcbea9BB6yn4ObyxXj1DZEb9pHNFLaGLSrBOZzvbD6QUnSpLrtRGOrUCVTm
ycV/BTM+6lsugZdCGgft88qRCRPG69OVDC6ynDhXirlR9xaukWsdSecmkwCuHdVVl1o8YtFS3j3Y
6JWH8moH2kDugGKdggkwlfdVb3wkAjXzfHpvZfOju7NPuzdItB6ttj3HxgHT7GfyGPwG/NlrPSbe
CZrdpF7RjxigJzZoSAAa2KceDAvLW+EIhO9BYUY5u0hb4+D+vRLYOx4rrl9DIos4HxO7w3+eWmGl
Sj8cG2UAdhfbSgGN9INJG0B6dw0tMoAPUwCU0q9dDqIA9wAY5pPDafH+/IdCUfq5jEjYRn9tXtFw
su1HP4hKpXuB+ngcfsC+t6QXOpGGKm/0gM9nvJFLZOD64v82zecwB2EH4SnqbV/m99WfmVikYA8+
94GxcI04HX63dDErRZSOVsUOBgZPXu8KESS07KOWtdetNkmL6yn43yRlorcIWgdOnsslTJp6VweW
sW49YvJ5W2beFGDrDBLQ6jqVL2Evy6UnM0XaQ00If0Es5xkSMP/fSfzWCefNPX5FstcLiYUtgH+A
sl06YEQ9jgNpa9w0UsyGOu2pE8S8o4us/bsZDUN20nYthwQB6PVozf1FErIy4Rqw4A0PxDGkndZB
yICzcqp4h2LhPiq3CkvmhwMgmiXm5kQk0darXA+iRrJKlnA107wQc40LF4aBUOlFOtMQ2PNWqtVF
+qoCFjNZTBcTWxYOssctW7/JCx8VSf6MV/bHmpU6F9+3N0xaQbdeYlneRgOyG9rRJ0xAD3bGQtLw
tRje8hAie+hdf8MQ2SPvYE6VyvjkVLz2y/J2z4nWpqWNCe8rwdyVPXD099nsx+ryyc75k/tsTy94
4ZIWVrcn44t/SlPf35zjYpkhcN0/UCmeeqw41Aq5MKBPjJComjvBfYoJKqjidOlrNDQkVKy2SJHd
M1OlI+oaRXuanmNdQJM0CDwhHsC+un4kExYsU0SVCFPKGQYQ59s3pS0JIoGZOB/+UPXhCy79JT4C
QMOzXrYp9eC83FfDYwWkF8sSDxIch9gEzfkLwLAFCyrVFjdDZH/HqCHpuifzhiYhFTz0Otu6tQ03
f3CxO0bo1fTzLjAScAvS1cB/g4bZtYaJOVaixNbu1IJd2yJLCkCC3GkKIoI6tPxpDic2+B9NwDMN
B7aFBP85h24tnrF+LRIUBpRdHRmoKQq1hUnP7qd/VhdmZbFmzKX68HsgjzBnKUBNfpe8KI8pwtUU
6x3RlCO5obSW6QUm6Fc/Be8MOBZFhSRu8pdBR9jTfco6DG8fDXj8S29iVspqCT15JNetpNA2/HQN
LvRIp+7TFvNrcBumzf3Tah8YMhrL4AjAtCPp6WZ9DRzrwPQsA0sRzotWzNg0BXZ4KEKzm273vE58
ezNetCNPYxw/5oRvCIEHq6ximSfO106Erxdm0X6aWCsXVTHQsRSnYP4b7+VoYQEhPW0cYK4KOKu/
SFJghka1pQyeoFpEYiyLEKwod5JFGidCtcXwaZoEEPFk5QYFlIpVS4105hS/pXHhSMhpDkHmiYiZ
PJf0qnqgbSqO+pj4u5oOL1hm6WIrRnoa4dzehdWfHPgn1ifjJA8sugLLXCBiHNw+vM+eHD6hwzkg
j6BnNCLPBHAbfgc/Ao1JaaQ2AV+iKZ5QZVbNTULCbsemRF/oPytpMrXKefrryqTkHftEmrm8uQ9u
IDTYLhXJVHcLA4O2scv4EO76YCo00FEbMO17Euu8PsdnmMaixXQU7Wx08ahuMH4gmT4NpS1zLT3J
+wegYYA6kS8fdIkohulUMqbbV+eMivtbArLSwLNqqY8bJF+6C5Pbn31ZSyoWaOtKQd64hywnnIq2
JoaZrenVRnkcJcK/WjpMlAt66BsHXh+hAcUpnwrQ3HDDJMXkpCuubu3n4JkZy9x5yfC7aQk4KdX8
e82aGpqspy0+q7w7Wu+bpHMRa8SDOR0ucgRxUeqGlhM0vDlpPGXMDvjvrwoIZEUz7BXlhFd/9B/n
w9XOYk3R8EgkeX2IZEagOFtJRxCXe6NLcGtL5y8k/6+iDfBlWTn6n2twi7hKkynfUe1RswcQmwOP
Sb2vSXGwYeEktvmGXDGBc7Q4UI3GsQYtEhH32ovV1wKSl7NVdrhKH/F9qMmFjWAOG/5TmY/GTR9Z
9ZYFXwXT1F+UwN1vlBHZdCz6oEJGDJypDpcNEP+kKVUcslfjM8SqrH17vEc2MnBQwmUFC/zyDoF2
HlURvSmI+Yg1C+kwTTVhbZ//bz9CjJlafTI5fhvDeiajAv7/DZLCGfX6xrLkgeme4ApONK/8TT5S
pOeku7x05/HaTHb9QXf7KW3UuNzF+gOscS0GKvKhldFkfOm6xGxUoieopgQcXO18uH8oQEYz7+pI
///iunQo5mUEohK14zpPYwFKO0QRXEysbqrY4sY5FkEMC5Ou1rs50tkK5EbpBU0zqOBQQmBkRWK9
4uwfl/QLF//GFaP+vyDk2lyn5K2CmkKMHtjTVwrZre3m/C8i+3cbN66MSyK2swT+0sDMFtmznh41
310r5DCSJvzuuLvm076leeg+WMLmMClZmY6RzYgOEFF3EJsGmjusBpn3TYJZKGlGgToF84m9DRGX
AQJcTec3UUSPBsvL3u9Guuyhsp9J6JQU6tPjWIBua1dcaZ0NCmC63Mpcz9r82la39A1rpJYv1UAC
BOWoW2nCrqk3SU/jE1RglF4dCrbxOe3WC/JJBxWsW/DMeA98gB+waOABWaePZjyZB7DI5sw1ldcv
ta98SuGP8ooY7jV4idWzsDe+akwla7VpUPWqFFG8Eq0JynMl9OwhVOli3jlQ6f1wDlhBy3dOKTuX
MoYr1FPd8vhuMBY40JvV6YKhBFCZwKU4b5CD3fhi/iWpThv9T/z+dS+cy5XS2qXjce+KluDrbsPK
fOgOtD+Ox/B8xlckXss/rggM9dJvClEi7Q5zQg/+H8Ss9XASBkIqZ2DoqoPXtvb98OOLm4Jxm1gH
Q49LmIEV6YdXeu5DGCbB/fYxUSVNmJdqzUkdz/dEGinInUV+Bhr+PFK0zFLfMN1WY6V++wP1wCre
4W70vWJaLuUEY0fCB5jJ2dPhU/95XC489jbFUOnnrt6i1tJPfdw8EtfsT2k97RnCi5+ZiwtA6w88
6CtOdOi/0FLnwDXmATxCuijsohWtdM8/Q8Yb04yQXGhmdW6tEYUyZI4pRO3yGGuifSVVCkeCLDOT
8zHs3lZog/UMWayufIwNray9qG/65bExJ7bg2xyNU4o1daftiEyErAFOF7sAtD1YyDwnuao3c3aw
33xhWnSZD7BsgyzCniYK0E8Exp2olPYbTMGFn+jc9LcBVIR8aQHyDPpY2dz2yM5YQ9SHW4dgXRZx
QqHGMUrBTL+VEi3pw5fO5c5P4MsKNoilUnWGYdjqMIzFCleR0XhNPI2AQzS0he3iIuSmp7qN5fAd
3zHNvnKVTzkMTi6NcZeTXs04PYnFlbTDuFj/ikJiSxrxoXUcr5PaBGENnaUPlqpSByHXKeR41MVS
ZFxLM4hSiEX3rs6hzzhOBWXTo+aPXsajKxCYy3rMEFGiT1sak9e0VypV2lTg8YmO1FK3hyHJYvlY
nuDBhhP0pW3h0dlflIRgOGeq/vP5N9NdiN9vvhtQefJhB46jOnDUnMvLCX/Y9tdQG7yV1yyEBmhe
9pfahTFlTRi6fyTzPT+oUr6JUWZHCrkWW8oB/6rhp16mKi6Z7kuWZXaU04wLew7iNQICzk6yobmh
PwTRoS3jreBIfbo+YER/CS3tOj9otySxAAmYAz3eigbraKityXp1BvdW2Sq/gidlkLJ7bvpboeKE
WsZLoH6mP7cw9Al3FOhX0p0Ir6LtucKdRqQiz1ZDpww9J8yHfYEvMpTfyFbHRNXSPJlsoHNsIUDf
ySfnVGuzO0LhPeLoiWf+qgkxvkXPzMP/LGB+Pk93fzpTCmwCdkHooxLrWiraVhAyQguRCoqe914L
ufO4D8nP523QHsy5q5yFs0yDoJ2csH/tG3/AnkYfNJYXagVbkIOFWIB+iuDa61J4Rm/w2M90XkWk
YCYnqpEoQwJKh5G79YfcUH/Zmkg7ZzmXOYbhdxgl2HbSYDo9GZnPXkd7f+D/RBm27dqfaYXXWQJY
u9SrKd7VMzAGUWDJxhnsEOG1z3fvJa7LIVtvUZnePpKpr5QRvrn0J7luXIw12PmfttPjrQah6PTy
leA+jAlaRkXaCCDVMwUtrz9oTRvogzwJFCDCVscwWgcTEFTn9/DrKad4iWRvkZ+t736fnC7VUoVD
Y3kXp3A1WP/O2co0gI8EeNHsiDXfNu+k4jyCbC4pBVDi95/d2hXh0TgS3hhoij1T/AdEWyV1fxFv
d84S5SvQ7MhRHSQ/PEN3AHO1BGzf2S8fCGk/AFsdt0osJesL4lsmNsIUrR0KsU5fB8d45vBS1pi7
yzBeaqBsXzROqLfHcuZRTsH+R0NBICykYhPk2CAO78vLWVr93WJOuzA8Izmm7DMPmBjcROe446bX
yxWQKVUobafC54q2D/sg64r22SaBEj8C7axrBpR0RoUO5IdTmjZFIizHg4+g/U44ajGUBvhJlQL3
HHrQPd4Zc4mRIeRPjSjwqurtKSJHyPcEDDm7Ap+haOkkyYHlTkDAYSGFks5dGl3ge4hPMTbwQuxM
afnqgy1akNau9y+Z3pgwC8/W4WRjwBJlTNvMuncnGXFsxv2iVGW3wBGVeMlpx4ai3ATIjvkT90gY
JZDIhhg3rUu/SKWSLUFELq2465O09U8p3Nc/hItxQYlxToVjfF/Tv8Z9Vdkhm1fIdwjQgBr86/PH
1xPEfXBaJphwhqP/Ccso2+NGoEinY/McROmo5cY8CRk5SpS7dGa450KZ5HgAMEn7+GrgMhWp7EvS
QX750zg7DaFuht8Hspd3Ue6qiYl8xcGIhepNgZLBRpGvTq2KHWBU3jiEnxYgKtY9wCbznTXmvtrY
rNhWKfBW0oIbdVkGS5Vmz533jzejnkNLwhSQzmjImx+rRFG4tdI39U12zPRXoCluixI+sn832KbV
kRPIz/MOx/rvffp1OxYDxQ+byJTRdAf0EPQqQEoZm4U1kB0W09T0CRly23UUN40XFcmegqBL/PtB
UNxjCNYTRrbvGTMQN3rZATyDosFa9jKDpQPLZdFvHUOm4laZGDbKHRDUs4tBygMYvUDk1j61fpHe
22VVYHR7G+E7399jLPX95Z91Z3bipjQA/XzA41rQfREPkM6+WQQQYR7giYbXoLTQuKR9MSLgOsD1
W2GS8/3dSbFWB0udTN0OAQnD3IVMYG6VuCpjjgq802PhsoOEnQ7xyQNVjqJcQKfqU5XbXmXC/E0p
hzjssBTd++/7uvqCpKXUOvbfkrFusln7+rJNScQTBSidWzLgppwAEibWvPmQKhs+EdTtCHAsQKs0
k3LjOHBtcNKaiIcXTtXwiI+BLaXFJ+lATybd98kUO813hr/TMIMyDqUmz9ZvDCnalG04bOuULVyA
IwDdH4FHgKykPYVlcQAwAXtiPlxFLt2kkD2/zjDclYKJPo+mJ8+83AjtpZiF8xhwdGfx4hMoeMOI
+iku3kG3OoMo2KhIYg//HBAn35Lj+sH9xEkbGC1ASN6OL4iU5OEGRKwga5PV1v7DkSxYnef5dfug
vE1gjZHgwROJocdUS2RIxcsk9VWsxnGsFeUX5DPjJG2o2xLXe8jJUzQTPibfZdPyyStDoBKicHu0
h/mAtJmDpvQscHMxpZGaizilaBQlDTgQ3fT0nFSP3Rb1VnAMPtg2DdoM72JZTxAk7YvOXglzDBUm
3rpi4MhEXr/H+eTGS6llFeaZT8lZawEo+c3q81uOu1FnT5Zwkj5PZHL11HlUWxHi99mEaC/44yUV
o9DLjbKNFrtpssmYntQA7LPdzclbv7nb0lA6ZbFOIGVhOStbBotILeqyi1Tkh+BwfcW/cmqxVXEW
6Pfnh1Jn/Un+zTPiw2l0r6hgMV22Ipxmx4DyBBG5MEt3F7ltCGXfs2fMt7RoRADR1ScuHEXtN7kw
q2w9V/aXMOg0yNx+AgYE+Z4qCPimcdzOknxXbXe4lxxIYNqq449F7eqJxChPGpHTsaaMI6Tr+9jJ
6RHfufDgttVJHVuj0m07+QsG8LsFM62TISXSL88uNCbEz/OBYrXJ8ycedbN+gwN/RJ5R9IDqQqeG
2RKnq1txoe9mXWkeQ+vItXuZhMchIrX+HcrOn0S98x4zEQLLmFzk0gs3Cl2jXkdxzzIug7xEiIFx
W9joa3AnzCLtoaI2cJGghIxiH7zuAban1ETF5prsFhWJznfKIx9Vi+6atgE7NFq7d3eLQEC1A27/
Hg8o8YlD6hmSzUrxBENAcQH+qj11n5bs7KM2Mu+xCkUz2g24XW1uDNbWg2P/NzBeqvA8Kd0GMlL1
0jsCvsBFGfHlw4J64VTJuooxABRqRlRbXjTqo/iyyhs0aFUgdEePCvzsauk9s4/Yn7TouHuF4M9j
ZxsGtBEJHHzdqCLYMb2PgMBTT/LsKjkhQUJFymTT7nx2K60K0mI4z0WuAoiz/3VVNTaD0TVaONpx
bx2iOde4/7xHz5HTd49Ap8scALlcZSNPVPCJKN5ugC0DWvKQ7Ks7gHGwhf4llVKuDM0fTiVQDVyB
g8gSNc+03uGJy/po3S1z3X+YIb9voOKDpVrnNcavxdPaDUORFx6HnvzizBVawj1+BuqxWpm/Fvy1
DDroKh1kUsV+CXiseJijIbC/kp7DelaLLSgBDDZiw/ZpBiM3Vi74L6zJVkTf0mAjdoKlOl1o1SGr
EgId2yK/a7LqQnJ89wR0MNuyun9Hv8mpXYRrvZYdapfZDmxeCtEByszjNLLHVWoUP5zJaZ2TWoKH
IDrmhG+C1WztqGAHq5h6GHpghEGZWaPuQC12R9jT6A5FfneYZhQ1h54i0M9FN7eSKbNlIur6aO0D
CajSdtkNHTZcbONWgubK/As8JQGldqQ94XFAfHCV1sVqQfOYOABGaD/5GdujVjn7UTT2VIGEadkd
T6Le+Jkzu7YBGrCgEazXOhys6eB5wq+Qi+i4FzD2x9363mLohpXU9fE0g0TPA1crxQahbTSQ04wp
2T2pcVD5jYwhlYXHdijxOX6TITFnu2PZJdK5vdfL9XCV4CRwKzI+D8CVi7ykNaVhqoYi5mFqbQoT
OH+M0beIpDLDIa6GAzWlZNy76fji+E0Qco9tk5yOBSomwk2hITomySFXcLObSG5AgcZ27djSjmQf
LNNAmUqkO+EZWoU8mQSqINFPA5bSLGqtwQ23xsG5fwQeyuj3FYRaYfaOd9RfaCGLBP+aCr2LO3Nf
+hQ2Y54PLokCvD+YuGa3D1e1pXPIN07XX4p8RmsgN9IggkHznXKcMFSYiEroUwpBI/xfRkrgWKRY
OxB7nmpukRvq2BnJivvY/fqy1XM3AviLViME85xv2GwYYlheAmiAf6gZL/vuo9/kJiSpkuF/hoNz
RpaqrpfH7brGbpibUOG8qdAZgAOiZjxemlH9NSGUJP+n8wshWI+xOWsPDacC9tUPNZYk5jWn6+t2
06zb7eNO533SWpN24jTnY0byTwKyq/ekCjLmaUyy2sJu9Y0iiHV1cunFr96JqdKuG0OH1AWU+35a
9ebNb/cUD4aKYMkugWRF9FcrHJnN5+b0AZwh+gUe+ZAAN18EU3MFVq64dkzP38ph45u+SDoLcdNx
TvH3+4DYUS3Fq4jcMWnlpF/GE9hWg0K/01ZaQdHnK2vPFSRUJV58mz6y0ynT7TOi7xUO5UnQ4Cu2
0SbwoqP3wdVwPOHe1XayNCLh/zUniRoL/CDwHkcEQGZ0r9sgydrhjQFMU6wbrKUsZQ9IU/ZO96ug
PA35iHGGvJa5kcQmFX1lQJ23wMjVKY4a50NdoEGRtlDXEIWE3Gd4JxCYbGVuj8fJaaufMqvE6AEE
cwbsqnjIQlUhDh3T/2zNK0TJBMgUvb52TEFel1wsJcfi1mk6ihiZJy3pLBR3ZYn3DK3KN72crCwI
njUQYHU02SQFT7oowicRwsoCRl9J3d1ViBWkJMY9J9T8RHTk4KbwZTyhavLERgz+r3wXBcxyqKFY
cF3kORNy1dQMncjxbrLD0ZjWz7LArHh6hRoE765cupF8NeiU0iU10aJ7dNyTghb/Ovg4dhSrsG70
rKP2S/Yg5dJNW+AyaeXlB+S8XT026qRmfPznneEtJ3vbQ3TRYb0UIXwXfVTqUOIVVcWqfks0q1AC
9hOShy8S38kHIK4mekp/737gLCjzs1K7TIkdLN9E0ibYnepkf9L6cBnhhWlD9k6HxlEgJiUi++89
PwD0febdxhQNkAGgX33HbCGjUTH4c7xcrngsfDVV8z4hv81WXp1Q4z6xAJxXxTq76S8U89HAv7Lz
l4eP85wJ1YIOlrxWLDbp8727hd5D2Hr1K28Y20CS36+6IEt5uTzGgEUkjrZM1NJ7EuebA11B90jF
nbs3GwCHwuxucb5Atp0LR+mQMZn9+5Yhc7Uii8Sc0m2bQc4ymgpTsuVDcyQS6XWUGndueO1znQik
DQefImmSMP682GUKYUp3wm2Xw1m+JhGSUq4+y6eugYOCnIXT4MrgWbuzwavzq32rw7946PxwrQbs
t/KaEXLIdWQiMMfmoRJRXAMT/MsW6oW/200ETlSJPaCuABT9fVtEvT4x+TiuGRFGAPQjiWKM08rN
7feAfRW+QSV1FLT2P7nnbmAfYBM34byGdmFMJ2lTNATyRJVPasp3UD9OWaSM+P1ezhO1wvyDFOa7
ueoOQNHtN7Go6KDCcYEyojcO+BA60eRvVxdzqVa206Y7ZcHJvRIGyhWK2sMfH28kSaltF94IEpiS
beyMN3TIIX7fa62QR+8KY8VKk2Ok3vOiXFsWMssSnXY68gUaUKDHbIJltSIuaOzVNdWK4+UwmhrS
jqwSzdYILmYSQpsT/Ifrohhtvv9MwPEXucCBrkgpCuKVINQz7HzllbT+1nQT6BDQZKLwkOxiYWES
5yDKqdbo92UdNEO30u2GcBGX/2XhjHE5/Bd8bjLV5Ngc7O5rJiNU4Jjs5zxAZsKKpWjiKmyQpuDU
eM4erOnWPQ+2QUIneYOFOWnCpeYr+TChL3ZYTCffq1EKLO2P/hrRmKKxsC+IJ3lUtn9wS6ufo6zW
rCMWC8dHNjLyvfuEkI4/x4PIJAJugwus6v8PidcAuDhDNArDUjOosXztOAlvi7DMYxC4CStnkUAC
ZSQfQqtLiP6Rh9fnnS74upyniRFqhk2zj+BGDm2rCgjM54UCaQOW7eAA+7HWsIkduUiAuWqIENF7
7XPZBMFHMdb6/HR0Gg24f2lL/9Mniu9kIelOdwfpPkgQ1z4yhoqovCFn69AjVZBdtvdJ2xCF829Y
Cz6iYO592dIUTvrpxRH1PmakG6w9l2Vq6Ga9jCgFzPMoNoL84YJqQKwXQz8ghBUbD5tzKCRkxmwp
60tgSN4PkmARcpqZ7ahbQIhyR4CkpTqbNHMmmsUVorZr1WJrYi01/flQJhXRYw3fR0ijc1vd3ohA
6aWHZaWf0XCkooPjFRSAMUDHexnk4x9f+5nZPjk2rFNttEt0+aaDjn5qn33zQBs8VxXFBYRoURh6
srWhuACSoXqx7YHI0Gi0ofog0UDhbxetiPD14jk27YnVgMxQIkhoQd82Oppa9qFGCEUGdWvmMg3C
JMfsvzzT0juBxpXUfCLWHURD1mjEFPrMv/t96L0qYaz319JzP5bu7me8mHb5xr1TT8ycUVwCMwab
wscRlCdgwpmwNx5aNbx9kne61z3q/o/NczJjyYyeXOICo1+HOgzE27futngz0zUOxroBCQEPD4xK
U/irU0mGuTCPvphoFW/wWvJCK30pdjYidMXaAMurLlguwiNoYFIecJEgucl43D55zQSjrH72nzZM
rVVnpYxLmvrFVri0pAa7JHZ2mK7syhjgljZYte7FUHUOiqPvvCNz/K1vZhoPxvGBxZeyf1FPlBOu
5hq73teTKQTNWjpkXCW0siERs66q5T+qDJMCgrSqaFPqhDaH7Pc/a6MrYCPSWknYHpZMWPXATlkn
Ye75756C22nYMjfXma5HC6YYwOdtln1aZBSguLXbZLQuHVH/ZojrtUu753We93QSD31OWwKe1qel
3wAzF6Uy3N/sQh8Zya7kNUlAkanA4pZufKCufqR4JTkYMBm1xkAg2qIbAtlMjkKrGkUreA0uJ8kQ
fR20x2CRHVAogo44Xa9ljVlQ+iemiIK/deWstAoE5eArSuPJEsx+DV74DRTF/UHaMmsV2FFqTB0d
5Seu1veFZ+lnPE/aU1g0RYKb7Lh6MdEFbOs394MdcL22csLCXIaCcrS/ywKTtTzZdaWEp3n8XYBi
EJrquVHZKQ5qDq8FdCCbCHqthWZDXr3Ssg1F+npmmiEfmi9ZJY0LKz4wdF4IVQiuyf+hkaUlTgnY
DsGUhLuJ33/1ejmCIUiAc9WLJysN+df/AeNb2m7wtZoEY+ypfK56p/KGNPvsH0/ScglfHbRtXDWS
ZzVIuT9ZnY1xs6He4Hp9Lk2xuyyGUH5vt6OwIlq5RPccfKh8erOCK2klWkZgBXqrGDNsmS7R+gRp
sv47+X5XEdTGIrUqV0VHzW0aaE5zEDEHPkfI87yYK3wwr+m21+hbRfG4Jci9gRao3B86ltqkEszq
ZccYEzrX9+82h93PRI2LWCopuzQkcVWfh+nDleu01YTmSU8+PfRatCdyB+0AlgdtngMlen+jDiQJ
UklKNJtfm9/dmRlK01iISXBF1uW9PgrfXicB63ztdFo3KO/ycSs7dBbDD5D4HsFhoHhzEtNNWM/7
LRXt7wTiUHztCwsMtgo9qTRnY1637HiDCjmkL5z6fWB2Id9E/IoqbXLR+Hzf2e0W8ZCYNP+gyPe+
BgItz0KJy6M6TP7Q4Vfsj7MiGxXWb90Iu6QbNbMoqqvqSfZyCeEZtEUmqbS362q6wfvjs+EAh9Gv
9mNOeBqVqvaVKr6VAD27XMFJNgGO8EUtMbLI6LZUbR4QHJ5VHJFgshgCp/Y8YjlHUjUweruMrhv/
oEuCXBbWJ3fYH0PhI/IXGzmbPGQDD8rrZmBoyAZhdMrMPU1DmI8GaRX4SRkok2kYbqNFwnu5m1ou
nWYj4025hztV+OIW+Iw1trAQMfwE+gft2FFsWGxP4V+c6GIgaxyOXi0smdgErdWC3/IbQZPa6I12
MieuOMiTC6Pb0zAUn0lkdQzT04jxCEMCQqid6pXjK6bGFrY2On+p6d/+ZOtxZfwkGACuO7hunL53
3ELpkYBKJTFGsl4G5wTZ6z3QMoG0bShhBtvTskEU4Ge3gJNeVl/bENS3hGScPik6yDpkkkCr+YKf
uRrEJRcjaMP+BYfZjVTZCmWMrZSlBKJyd2dQQxkqZzU+VmmBcA2Lxq5oYP4JVhslTo/Vhtf9yKBS
G3WUF0kFjDKNbGWRDn5H0Sb+DRcFewzHeFzYOQwxEcN8c33O9+y6GTa8vkKQBMcLSB+fKuh88agt
P1IATZKeTO/ljXihj4//tlcIV4L4YYULjxqgSfMAjXMQuoD2kSbCxUVqC3iuM064WinRABem80zx
bJoU8eULTHToVz/cuf58VRtndIxAH+cZ+FNW1RDmpTxHYoi6rBG+cCQu0yuWf9xMDraKQH7f52uR
tBwNTVQVwuVOd+mwVdYmmgiVwJ+SivSCMzIOBq6Od0c3xrr8KtEmk0MNeUfuI0ikiNAbn8nzTeOh
hOfKQ/W8O5isEKhzIUYmIvq0fwASeUMxILyS7hvooIIVZ1xmG0Dqq0uUYksJGulIuuPm75eBDLGI
XtZpFoAfpD4hvKaYqaXTbAdZYcfJXCH6rOqsNz4sy/P0fjQ9Qae2YOMjlQ2Auel1ot6LjwCjot+q
CNrcVmhLTl7Royle8Z94ytVH11SVhAWRdu/7NXVwp5pgAPcRXwMqUqtjXRxWxC85q4YugvCg/qOM
zgp+bHo9QiUR4TQ07xt6j84uq7btmEbd9o93CrwNNng6IWNpGf9H5fV6e4fW80QdXDAsKp4IX8Qh
fgW6myqC/XGDwM2nxbB/ipxhWEIa92DWbUgTvDTrs60WyDL44mTuqoZxmt/xB3BRBKeRG07Sn8oB
ZkvMi7NX8O2qetzdyGQP4LMt+maTQ0xWTm/athMiqjpw4I+TBqbdZeetQQImlExlm1rWl1gjP4nL
GJinlOaNvJgqzwi8hV8xPTd2OIqC7EuYUG0uLQd85QrlJTKRcfcFPS5obJHtw5oT3JI08qhffMPa
k425MqDEUL85EaoYGoR+hjU7h5twaWvXD29Lj/MOd0ixUkXG0o3/NoWhf69ksr+knQbQwGMBeB+z
qUBsUGMywUh4+PtC60QPMFdNx3rkmVWc+JPRliyPQ2GNyV+CAf+4u729Iv5CC9EOdMwKl/iAvTgK
u7Upbnwdt/hcg2wa9n8yjYfbRA4IHqaysLmhOaYUg81d5gMOO3TV6t1qN5KMZvB6bDWeS4yboQXS
uZ7AhIF/Spz/ayMIzZnP82nNgW/zsKqsGegQ3kP6NHMsPDXTyZXPBM9O5+HLZiXNss246+G9dAb9
2UXxEaF10f87Zil4edFgz7WCg1ZtsTUmRPGaD13neo/jStXfmCzzqAdFRV/6+sP2gx24c8Birz4g
wxV0j5QtUHmVCZH3l4etr7UXZ2Ra5zJ6Z+3/xtZEb75xvNIPWkgxpHLKuXUp+Cbhu4SE4jU5Yxx9
vmvr/SBJn3iJnbgDonS3tgveIu0BQ5nFFd62XDs0rbELSz4b/SRXrvFJuVo16ikQSAmpLk7EhL68
3LywujN14ImBXu1fcxQDaKMwxBt3HoXxs26WrlDLFoNoWxooyeZvUE4h8g9M5HhFTP9OcyMrj0Nr
KArWjCHpaI5ruX4IuUeH1NmTnDvaTV9O+AIf7G5KeW7cGaMCCP0PrzrUdmXl4rWMB/GruIOLF+1t
3rNNHQHFIxZI4+iVcC2SN/Kc4Qo1yaS8tSoCB1LzGdZpJ3NciqFYI/CL11tvvRy7Glhk2mlyjfAK
enghWaroMV+j5XVbh7gfOd3AFBSVMe9/FuK7rShwHe/l0SLvfikb3hxoBEi4qhglRTofM+9dQddL
8ydk4vYMcg1OhC9VEAyO8jVQKvF99XJ21CaHG5s5yHmpLSJil8JFzmthOFp9OlTyO145dLokjhV6
OxCTLX5WJc2ASfX80tRqJIaJgOGRKS87esjd24NyleCRFwS4rwP5DBQackCOzgyqdd/TqGToqKv9
+AWoUYDO45NqW/1IHdFzNqWXSf/KtKSiy5lZN42EEz3JUgJBSMPC0WiVhGHN07RX1+xZUr0slRnR
IE5QdwFaRSK30j0ES1H+aqv/H3vbFjtV+ppdcQj5r+Hi0qI/xmKtZzpBpVVnKZovnxtqpmX5ZEY4
pLbt7kBTNhsnDBnl60pBHjLRopzQj8QwdcLQlf3gKG4uaNLRQaXL+h7CxUrngkF7ab6YmwBGwCKR
pEYi6FPqc6VMVoN/ndqyeiUuXqW9B7/G2MWMADQRHxlAC2Vhc2CPoXUMmd7kPUTNlsRxrhVBbo88
skOu2UXpBUsPrBE=
`protect end_protected
