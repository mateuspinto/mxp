`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
SFqLNAWB8R1v4JnwmlIuptRVU4YHC+57+y3iX2BmrpuYkRsvoTbduHqsoK83s/Q402gsVMi6QqKg
/zaqnoLbca+bPiVvsnYldg8w+9iC/f5pVNFiIrKR45rMwLIipiZUTq/zD8qVn1WvCJrj9PEz4pU+
BtjP+tqrxTvW4u7XsToP37L8waehsBimdm0pTOc0reQF6AZjDTAW75IeVF7bRIfj8aZrbUT3ytgi
6QGTipQGT3d4pRWbFmOQ3ctnm7rxJHjhVa6MsRlzOLgtcJs2mp8qPW/ezzlGHlfVz4u2hLbYoIya
zilFqCiYFlRMAn6jRKDfrrvjgevscV9jbMi2hg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="6xmoXwSuRRDbMRiBeY+Br3Mrr3js6AlCDpy1Ey9fuYI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26112)
`protect data_block
pvPXvJ9QuQhl2ruMk83KYss0NUQPviObQLsvn+YQ7j+JGdPV0jZ9tzU0hVkwzgxIp8oRc5sCrRYO
mwCIkOMMSZeYbsFlSod9rWo0FeScAKZzz+YaD17Cu4ABEzAXVBZRQijivraG8cO2PZhxEYmm/YKt
nfhbf7w4ZtEKVzu7h6muO+8/t+qdsmlbcuH5pIHHoWoHKNoR+IAoy7gv6D/v+ofT2+Xq6NvFShbM
vRwbOzhM7jbLEOliWB0rUhCJ3l8ULUTlSVBluy67DEwyBqn1n8PsvvuTu/5E76Yp1HjJ8vQJ60vI
hH6+YKzVSM0m1AczolZFetDEetYjiKEk0gcmJHrjI/YrPRtD8QTFfmS82yv0WhM+sS92m+o8cnAk
pwIcxLmHH3yuWvFFD1CXdUQMidY2EFOMIRp2bd4O9M8+BUkiCrYNIyfaYkmhliVnnM28Gk9AB5Fd
/SGjzjEqDxu2hnpNLZqjYo2+EI7P2RxrsjW3M8eRhHrRELvYcvJ7xTSwKeoBEAQq1iYiXt+4T4ec
FKKin5g8hUR6kvzYPypzEhbQz+R+wDyfNKahr/y8Au/WLAr/JW/G66qNor00cqf1x4NEi6s1Uobd
RTSlKwdqHowHsQn2j+pFn5WPQGGHqjvMzp05PsoOJDQpV0H6Daa9ZuWgcPjJud0bqMBUcXwEmG0c
7MHG+imuARwbqSi0hrMzRL4eHmhpRbS6bH4V3lMJRxjSne36dvzXBGyBbOqjzVy184kwoqY2mpHf
+WAHc8n5xhSna7DYEjvIM4Aa/7bEh8W6bPbS7+alp4m+oXs60JxEV7QiRWjM+coasQ/c/JJAPUwv
7rL9wlMHJbvGpnIrDsKsUhBt1E5pmc0tT2Bc4yIz9lXLBiIQ9M5hP+toqMX2L5M265keQ6Zs097/
fY0Gv3L2NVK+YeQreLc+e4m50PkeVv5gKUUeemfpbRDya/8FjpvpvaFl4I/6n284Xx0qMJlRmXdB
DkG9y7VKUds7CJhUOt7YCqwSrIJQZDqg2ae9NhWXN6M6s/10PjSsDbUmxzK+Sc29JSFxtkGN5Tq3
+2VxANhhstmSB40mvBTSXwPC680cwdT9ySGI3sQZGm60+gCF9KVOZ6TS3YFGHcB16dFnC6OqBYit
CLYwDPFHs28uFOLkwJWg5xIm8oNyfvjdH9KdOzxazo9fapE+nGyKr5pOrjiyCrVXH92G2n8+Q9MR
CjV1ZBmMU/XxTgMm50a77fXhTIelM9F0N9sJRGJy4hoHlIp0krBQXXWeOlQZXdaXKM8T9mMOzYLS
ayfgj7NZCjwSREAbEjoUeI132ly92AU5axRn7dSIOqFwIzpDvRBc2i05vhz2j8RPqOYCtgEEr7bW
PnKW42ffO4TPmSAep8T8Yv+6QfMPig5hkkoqjCb4XluTj/HWdbu5BHoWud8kdLe/40W3O5+6EnPV
L52SL1aXdedk2YzCRUU91bPI8dQS0PWjuJgQGc39F7X25bDYjmYWMVgf7eaNB2OSQNM3kjVxPyUl
wbG/FEQftRWONquSgSIBOrERxxQLWdIM4+VuzQu7w5fbTLu95wpFAzeo8czRjC1BtfF83BXmn4U+
CCOkBfKML2PyNYSIR9ebzHBkPNq2SghSBwGtSeqCCNIrzsmLSk8xHtTGdyWX/E+Y/q/uvxwPd6jI
GejM21IF7H7uas+YKeCzV9nHLReGn6FdpZXHk29t9obctgvgMPlauj+ReTGlnJ8bYmT3K9tJFKgw
vPCbyTqsJgPJhdZCdSESrG7Kx0aPMG04EurQq9Ifg5DqUqafvPtA7R2scioYYq1kPdmvFOhzB3SQ
W8GHDxWBrBYxmndaGtcRob3viKmxN4tGAC+6WmYMQgnWB3HAI+FO6tVhCSW4VLmhCZKgqOHSACTF
0qw8iLqRlOHxemA8CPir+qSCh4tOjeLr7wmMW9tDU/78ToPpbBwRjAT13OyYYqslLs0/zkxXjYfe
5CebGnSgEgr+XzPyiqemMmyW8sRmLFk/SM643iIwYzjmI44EUJ2ToioXdj9BcXIJ1FLnutCsAu31
t8S522VJyPFYOpam25vgUTmzeWGbluC/7Gwi0xd0bgKP2rutS2eakl9fBa9PoglPQsqny0ksRIL+
wRfbf2XbpWMznO+SPi5/Ke/K9kC0mqUzwRds54mGUb2wDtpyq6bEqWF7WfjINHFAkkSNAkvVutnl
szUC/fk2wTYaFiMWzXVckKoabtu4jAUvh+CqSCcwB2f52P6KJszpY1cpmk9eZfI7MLNda9BauQmI
r+Sy8j8YLow/CQzEu3CrtyhdwHmdArz/iI/b0WftjE+MajdL7WQCg5wulBlVQ8n+YhuuWWTr7pMt
kTe2WrQ3XZUOuGw669qdNj8nkcm+SZe+hRIsR0DXj1yDDEL1g23mQwARu5jwwUZt8jSTlR2ydkDC
F18V9hNQrO+79FMikhHknx7m5R4setDOJI0X8iGgAEvzj8FQMTQTtQAEftHMax3ImxgitZnp7zG/
8ULVxIdC78FTpm8rFRigqTrIm/Vk23SLkwQMuecYqtq+PUEI3uJde/eKfXuLSyz1n9Klj9uIEpo2
Wa/1m7WzUqZr0TVjHkDVTtgmhe63ht4MF1zP12n1IxAerI6Vd6dIYIaAkiexsfhd3/J3InyR3z1W
D5RSikVirzk37iwUXHXAm6p4W9aei92cNFZz7kRc4s0mb4t1AY8HBlyAkb6UHi4HCPfcidR7LJDt
sJj5T3NO0z+2x2C4VTqZZtH2l3OddOD4YT3rWYR6FTi5AG9oQq2lJ3CiD76eZZWsnXIQ6traiySa
MNHqn40OPF3QuSrNIKcQlqBKO8TG60l4PbYWbiLzApzH8ky+MKB6qjrOgoMm30HGoc2dbId/nWJx
j1YUxgh7l1Sm7405vX+LIee9eV6Bj2lSKA+8b1hHgEVzXAJTILIwiTRGPeF7LEdcJeHyo9ZhKLgy
8Qxe2Q12jLqHH8OYpRKEjwLyYwUPyetQ40QrYLPzIAAMQxtamRFkMXSQ43BVMNvSfyTF3GkjOYMU
eDxzz4mhyJRpqI5yqEvJt4aqK3ffhzNKQMED1K8KmbuOxpsURMecBqm818zmolfLUiyXEtPW6WUp
TFS60G7EpFlHwIkfgDCP1BZ+DRe9tNRa2OpFygCvVplb94mI6vgMIQ5KFIMmSPmH6iSF8MeIC/s1
+IIVqnSu/iwMCRNlryDqFURWdafPAGx5kg1h4FplWG3SNflAYbL9ivb5kM5WrnhtayPT5A+ixiq9
awdZEMqEGhORgH2snFRXjpqNf8epMqhNrZAUcBWqmCW5GUE7U1YPTSfIQDjiTBu22iwJaOSenfbB
DSGKcRztLtJxJHg/i2k0zU95qve8MI+So/cRKnxjKJ+t1aTlPRYb2LwpqB+MIvOIauERITsVPkmC
kZKbFiOBOA5fnKYkaLKQXpuN1cTPZz6d7DrRs/zjohkUPomwBZNLdtcuCq9yc/whxBumIpoKRIYj
XRQHhKJ5KuNcg1FQY5zumF+tOKu7MSLaB3tBKVs6A0KSDap4v3N9FevKhsu+YV6vx/O2gWCVPRkH
tx2BBodOlsRQDK4tIqCV/iiCtWkUJUHEGM8FdHrZX3nUhMybgiP1P5fT0H5jRi1sUWc8/syl/KK/
JY/7sSeRbw928ViuD6l3s+mx7+jJCJSadkW1+TF8KA1/BfZa9kTThfs9HMYoMMokkpgzaBM73BAe
TnVylKt7Xw41e0RIkds59LIsTe4RfRDmIrurFQ+3RP4Y37UJAYJgql1f4gtOvfZlAXE6hQS4MSHu
Z/v2J8BGA26wmR2rv2J9+Ahu70ntAcZLM90MFf8VHEKEWJTd4eHZxyHVF6r3a9d+VSWrQGpBv/IF
8mpvXDWxZiZwvXOkCgqEFNby8KqLXjS+wCDNqDCqGMWWJo4TPj+V+9ZheqsSJse9tpV5eU1a2jAe
Qu3B/JfXAC5kdeqDSKJce3skbX9bNz6aLOoBgSxcSKz9Xc9FrUCFOTQVnwhJUq/nAd5BE+c3jouX
J/iGimP5aHpXa7JrJAtroZNBE81+j2P5IRnDRswuFr+dWyhpSiEbNM5KXF3jXLJNLR9hmeHybCds
9BMdJOTBYOr07wpVWdd1XZfXAwUvALH6CMKJJBWCMkkUZd3VQEmJuu447D5GJvZnaGqe267M3zp9
myEqiHZO/DD7HDQlM7FTvzzAkdmrUuBrLOARcUVtza35T1KDOE+LIb2fqv9d13YDBsUqPscC89Tz
9cDYuAuSDS7/qF7EvRKMV9SE9bQRiYVMR60MKcS2IVECUwmHK0VRGyDl//qHGksw3GtOZHUijaHw
sUjVLbN94fXwDYoDs/3tJTzv/eqLTjwqOYxUDTPWPRUS2w7ZeCLRGLLX0ikEBggu7FEsnsWtCgL3
Un5ELHhKwr2ZdWYgotWpP0trYukbZiVZx/SxkPzv/ZU/U61AHCuStZZbY9LxIsFy7bheWzKOEbzU
x7Dndm+6nGsawpUTCerqTnDqE+NqJziPKZ1MJFo1CqF7WUmtlQOfdzSzo/Pzfss8ftNbRxSefwdo
QCmVtVJzHXQZFPOCdJXw1i0/OnbHY+WGxzHZa3uRX7wClkxiNBu7Jxe6juUvMHiodUFF1Bgl7Bs2
fVPXlSXcinRDjR8FrFNugqZNwBZWCF/WIZauTAZI9kvNzjdKKwi4LNTWkIXjCouORHPx2ysZ3h1k
mx5kvDt2dc4w4uurplszWHk+kkbNBNGCw82g8AuniN6KAoAvP91DgD7YXt3ItEH57vtX0aNHsQ0N
9twN/Cvv0osCEFrWzhCEKzQZQ5Pxk43vO3MYXiWeDa0BXBeiYfHP44JXZHz8vNw96BwMsKU9RzeG
v+7ZBr48F9NQ1aupFLkcpT8obd5rcOFDw9uopKdOsWuIcbGmXCmE21d6HMHdwocTU6GAYHC7193Y
EJspi20zDLGsOWmpbZMEcH/aayema+yggWWy6ExyZbdyOFfuE9iwWZmXzg5R/k3JWtjceFOMFkIY
ATGZtFhclNDENVYcIhW7o91tl9r+JJw7jsHOzm1SVPk/XSjBGF/jyGVqpzFz/wBDlfnyIksDmemY
UB64Fl502l916SmYoouU+eeroHLkkHX4xTFYBjnl6CmDs+KvquuJy+r4u9Ch9JsLJJ2D4o602iDm
OfBaoug7zTbav5rxNjGXoAzY2PLyy7F4atP0kmlAfbXYsSCLkjcBKvvuwlcrzdD+9vQRtG0w8nEO
Xu9puIfvXEp4YSj/yIu9Or4KeE/2S4g4qhmZ/IG7cD1qDcIoRmwPlI8p010Z0iaRHasDn6sk1M1d
nejTVXUXmyj1Ry6IHcd3JVcJDUJCFtIiS2q53/LBiAayVSIenCwALPnlwVYCVHBM7B0E/9y9+8BS
YE+lPPxasApEXkxtKPjQD3pB8chL4EQYlrnOSuu9lCPWZUG54YihxPSYoGFAUoAlIfwLTw34ntOU
EwuqCTDLeKS3e5TVkex1P5TBIpf4ApbUh8ac+b+44jj5NBBfG9D8qoBLAN1tAKBIVRgPlDMfQb6E
mOco0h8kB3+d3GpCFswT3kpkvdjNsPhx4UYRx7P5U4ZKkUA9K16LzlyTkzwY5WByzC7DFRmXPmgQ
6jkOROz9noKLFv24LcMLnegVBFxYRG1TRwk8vi117r8MKhoEe7KKo5HPmbuLp1riY5AQKtwDcy7v
Fi0w1DB1opmWIUwFPVG02T/uCI9Z0VYr8OitI8auo6BqYcPBF7nFjyT+jSXQ0hEMfMeSskIGvKtp
VDNqhVCY8zm8zh+5jrYsqqUiBbmk3NTrKfxja2ou/CPnScmCnJ4H0HPgKhNZjdWSCfuJ31ZUUHQv
AE+ZIzog8pxDk/KSXkuB+FCSYdduuQ+zcLVYMZjERhEg/wvJX4Jv4BqDYd1L0U5BpXQPIdJt37qO
E1ZObhijv8LzKVFhEGRIZJ9ZI+AP+L38YIQdtarkbUpcCdMxITahaJK8EumrWAlkg2IKQvTkUoj7
ugnVWMQfButme40rGQ43pa/uGmIcBejaa0FCUDAYe7wGMYTygABpCSBtr3o1pwCKlQSmMVODZ8mf
V2dvtu2gv4foPgx2DirdJGJRqlbYGbmFTB3aLuemubt6HfByy8gv1+5q61H5Y4O+yTqQ4T6MM/vW
PRhRAV02cqy//Yf5l4Vajr/mHJ4+mtzF8rwJYfJv9suPQjqOHXEANRkylLgKPuxsxTdGvrI5vYhS
DBWc6qx6NtfwEjX08r9PllxyKPXRQWrtuXaJGWXNROez6Dv4XqbfvuwYOw6Yq0mVFl5AfANIuN7t
LJ/Wr1/LjjMtdxATZiDbVw6oxqON0HhBfvTA+XeeOrqw+26PGefnG31fUq4xEzPf9aD2QIGelymY
fRm1iF99CTs4n+CKsXlek+oKYwXbg8adHc9hrSp+qdZZ8nSHYybAaIvub3/79P9bxIilNHt4O4yE
NRAcBvhS8wVjSKZjW8nn3TB2Ec6baUHu1XgO/Kxud1LmKNlCVZh443AqHjtnaf6snoUSJ6gXnD7x
PL/Ews4W0TnQhGDXWK8kJCO/JHTmUAbHjJnA7KibTAgeJqSsL4M5iVfWH775jK77k/2Qj0cBuOFN
u9pAWZSXpp47OZAbHfyYo7gLa4AXSRU+aZREwUbWuTcg5uMxkVRfp92uMYe1Bn0GAsNjdFZ9tVMN
j9Pw3mUov1O4dwhVbpzR+8pd/t/JLoeobL6OyAZAahWZ41NhkKjuC6zao3Tv1Be+61hRGts1shpg
5q5r0ZRflL3P+64UfIOmkArM26cYwolToUQK/9UwepcNt6iaD8LKFBvcSScDH8j+/LqZ5bJGdJq5
mFDriCIBALTxZVO9Np2KLKSMT/zMEZmnV5is/FN3bs2IL8dGrJXl+lEtB1QSuwcpAPkpOn6zjE31
dg+hA5qKRZBTnGMg6QmflZUxT44yUBfzF+Vj3eVF3HgRyjx6dP7tSi9/YHAiz1MjT68POrzCMFMy
N7N8jM+e6L8I3GrzPOYG9vS1JbQYTZaz16O+6sTJfsDDW/UZNbff2iQDL5qTHyYCiPn3QvGNUa4S
AP20EFMK4R7syID1hspU9+8GXMltVfZ9RbenfRw1QL3GePsFW/tkXizLT0hAPt26RGMDGym2oCDp
mPFcCsQ31+epDUUujfCcB1ok0/loPyachlEngD7zO/pqxTPBRzJ0mOOePzYrlPqOP4dH/2Q7n0M2
d2UekiQ404brbUZQedNA69ENSQY7pez+OH3T87pPMQtt1wpApSzarvb2TuPzd09ejeEdYQ8CfBrv
8ZYctUUfHCaUXCb+aDWdP3Wvq3JvrvbuSFdWhiLlLz0sZWQGrIVoSSQVVKi1o8br0ClC8MjYHu3W
I6EvJf6UCKQZTCWfWsExS3r8GieTlgA3pSmcvQZEWd/kpM2eVVlxd6dCElL7If2vIt8+JSJqBrq2
2byhBHwiB01noiro520od1xYFIdE25jpgumyD0tYjlNz1gwFIyEkS2zF2xWdDD3EgmGUIdxmndwI
GGgRmJh1TXGdorL6JVYxxJ/FBF3wzbpb89Y8CB5vJYey60Hh8D4pLOLn/Kf1i6hBmzPbzdLbtk4/
AuEuzJOcC4eVxBxDOTChCed+AufCKN07wFfOn9338vApTA5/8dN4LeKpFPi2Mb26lltiD3BCyQSm
XjGAIBJFzzQpVf1JDMukv06vZEfSdzwCmMKUI+VTqcc5xUjCMzVjtNivo6CelpA12DmR7mLKlmi0
0VY2i4DJeCuclhIgX4q7EIgUDc3WkMjWNkypnMF2gZYzHVLkyNfZXGAt6bpK3nXLx7Uz9vDwjJih
Tpnjml68vKkrabH0BAhAaQyUIGEPl4+Z57ryTQu8XwA1OQWH7RoavB5B4XYitBrIFP38UDUfwamR
cUXPcltuvM8qYQLOXFmFZpoxBxWUykwuoR14+hnQDWoFInm2HWGUnkePlOcvSjaqrLDufwtOOq5w
2umQdvfV3hJPU3PWGXWzjMOFl1Do3Vf/pUndd60I3GIrEJb/lcIo6wMgffoIvN/msaThuRwo/6DQ
A7zE+jMuikiWjGEyTXhTU+xs42pkdZaf4p7kwK7bFdHW/4/QLJa3NhnuTDyUrk8fV1L8JrZVtN4T
bVR5vEpcMk5IFcEeSUfbSITiRWqfLLzPUX+zeYvrdhtggQXWT79ZkYni+vttM8Y6DCJYg02lWO0+
Rqu6m7p6usbptm1JWhYWAePdvze6CvQc7RFS47zkkB+0yJxizpIVZu4JqONHqNNCWzMUa50vsY3M
3H118bbnfJlr6xAXuEevYNHSWLOEwy0SQB6JUr1vj3OzdQYi+g9bPrKeXN+Esz1464e5sFD7K1Q8
w3+jhGE684dnxg+KEDJL1hLEvzsVycFdQBcV5dkNdA62ZvWwka2nor5xDYk/dk876+uxR9g7CjNC
AfvMYjU4jbO6hIr8OzYH1ljcL83N59+dKCQtCfSfeZyt1uo9N/OvCulVDmtBL8Ywzq2R9fH2Yv7x
9hkvfB2oYOAC1myHBsC8rBU8fqnV5oCMQdZroLnAXsmc6j/blBL0AniEuVa0nl3O7o0bwqVE4E5T
68tCkJV4eNEUwmQlohSnaG9IDz5wBSR596fVuIcUdJX2oy8wJyIc9v7iMh/a7VNOhSTK1t2Hn/w4
OKc6hhCzLWlCmAuKgplRCHulm2JXUfiU95ZnnwP6wCQTqEvqkA0X+8nvb32lLgw39e5JeZ1eB0+z
eGQb8ElLUjmIX99AIdWm2Qct7aF4Q7dFWIAVzQ5AQ75JGQYY52QJ/LKyrLle2WLDQiTATAzU8I+a
ggoIWqlsN8SNX/BW2r2UTXAT/fmUWD1YZoyYWadu59GRLO8BDwd4fI2QNK7zgFJB5wbHV6dN++YL
h94yCy37hnjRLg2G1B1gGF4kflOd7tJfzdls/p0RZHIX7ZJukX71xnV8lVReCemyumyvvh37c/DO
WJsjXfzsWdrKUnL9JScnE4GwhSPxUwiIxGALY/2a+7Jthb47WeehOHHQ5vKuS2F4b0wxTQz7gC8E
9KRyojJyEt22e7jOZHoXyxzwQ0ZSGJX2XYS5LfOFPJiiC+9jANTV/Azpmxvo9270rjLKQnu67/u+
YDuq2y0tM2TiIULkCm0lSBZadThor5XM5CLs0gX4jxLVLPWE/xh94WOsy1Fym01eYUK9CmSXMjn+
uES+Y4Q3Dcpcdng63BlX0bf1IZGZcIRT6gVqbBYeLEBsGA9qMy2KjrQB4OgWRdDTlqA2/tdLW6NI
K3+EjilOFiNc50pJMPq+j/B8/gVA3zhVkC3KLRHd9f0x7eXOSsUj/XLiWXAdLev4mrzIaGboLmif
huyybn1823/IS+ZNNf80jyg6lErdqIgYmo63dBsnR2qfUtD/yROQhDSOdazbSw+CKlU6gs9LQo1I
rxPuDZZ3CfkPLMrCOPK5U751kUglCfaSu2s1lQNyi7ArRWt2okq5aa+2T5M6PDzthOeHqI/RZRi6
gWcQnOCoRdvQYDpHIVT8RyHixjElEhHm7Civ5FMWgXZIgK359S5HwCqzK7E5qhmOtfCDzd2Y9Fx2
5+Mcz0iFKa7Z+ewVqUOn6YLHBOMHJION2kUG0Wl6ozSFW2u7H3MlWPHObcZAfuPXTSjNkm5hZOdU
ilbiUYV/jks7DbltqYFSb0Czt3a8jN5aVnkq2cTauvnuQyHWd7i9QKvVL4edg0sWhOhxx64ksUgI
Rf18XgWlBBnQvPkQXTqdWduOUTI70lD3A75DTT2tFalunIy/elCKmqqTOEVwXD1nrQou2aZk4K/M
BLaW0cDWnnWXQcifBHe5Un7lq3AG6vn0zvNlZN86D44afdPMImLxTvt0DOZogBAGuaL40u0HcflL
N+kzu7uGcN7EXczsIgesgxYLxdBU6hJrt+3MLocGKifSLgVrSAmC0+pvYIjMNVVMzWvlfBPKqkFe
quc6npZMg2TZcu/PWrcm3T4mwjdrvKlpOuFiIJ+FKGzGNvhYSJqeHRS0n78T+TWxGK2WXMhS1E7k
qK+FnKYn2FSB7RodHd+QEkSV4o1ktTYWDfVLtwQR9wxz60HZe7jtS87I/0Q+cxxyc6ZSrlMC2kx3
3pUggt8RyRlpYaFLEXwnd1rr4OvMd2bJlM0Q8kcffxStGuEuOfsbzVNdeOhxlrXNQyD7+xgEIEdC
OdZXjg3PjWZTUMVlKgcMy8sveUvslncuIfDmthHOuPJBuo1pNM7ORPO2dqKSqupK8APQpugosLze
mZObbRJjcXx/p8p5/idS1la+yJ0I7cmwR2J/LxAeRsT2wSuC5uOugSeFUHGVDVUTBLTZ1nAY+82s
kr0JNdMv/h2V7RiYXMSmAKNSFKOdD5n11eAPuweYe0awnHjo+HYgqZ9ncdU2QgJACeNpqibYr8n8
st2Fw808tzkui5JzrKaUh5XJj30mOhI6go+g9TYpzrnX6sZWOc+QzLGcJu9viAYRMCXRYbuCo+Ek
eolY/eRBf4mhbRv30smqHkYUJk4LMn8P3DNcnXZDJkf5qnwar00QJ6J2UPrKUKTO8F7aqOcW4Zgb
u7kI9+BvnJqzOIZjG/1X+s4ZY/ir7D7qGpNbFBR1YpzqaeMZwJyHuXsB871hKgqMUMY805E+bXie
qm/fHo4BhtgqfihOga58bOGU9u1KIPW6kHmwcmkKoPUX13lL1EPok/nbNDedFV0CzFP6Gs9u+ymF
TlO+PyKkzh2Mx1giF2YX+kxQdSvae4IsWuK4JX4XNbQm0w+dOqEVmI1AS22NYM/70JV6ICZvWhL0
UKQvHNO0MJQcvm7tNXeXgsQJ/Hy9+NBJVyATstgbHGY2OXYo0hS+2VY6qb84agN1QuyO86WfVxfG
s3GQXQQI/Ko8BchpRRA9MXs4p/T9CNI3dZuR8MAIsJWqqVe6t/MKBgrz6B13tzCLZnDROrM5uUvS
058X4cifYvQOOCvUM0dq4IxrbxCac8cn9Jt/7PcB5wh76POqajPYI8P4ttFB4a4YFn3AlJzSzmxn
dUoqjXiNAoa2d6zcyHV78xrt4xnHAgVmNnBR6+xaIcKTrkwTq78Yj2P/2evkT+PpOkRECztSwZyI
e4Wsq2vB6KURdJGJFa2pQqBaBWPnVBqE2gHetaOAec5H1jfBWZMoogJZfb8+oPe3gr5G0OxTK88H
MQodkKErz0jHTd4+p7bTU/ynXTW1LxC6IauwA6hkxiuV0x9JN526jG4SF3+r6k74W0JNtCA+Lw+b
Ywvjds5NS4y+gAz5gmvp7V+5wBSFhl8wXuJzEhD/9OzOKoaM7ZHONReMnX3APLcNFCtCiCIdozBW
SgVBY8i/A3PeD2oYBuX6K4+ADf3bXqTgCFDyo/4mZk2ChxzfTlMhY2WkIWWqPOghE0A22t5IonMB
6ENgiUbMyAtDU+TcU0WtqadqIkUfUb6VXidHyLTjyuYBfE0AgAT+jeLguVBlkrTLY5HhRoHT8igv
Z2Gad10GvoWLXmT7mPzi/BS0U9Glj1gQXfy905CZlMi78tlzASAQCafyownihuhe0yRHOwEBxwyX
WEkIqO2Z9dxfno2nV9BwnyivYB7Pf13vaPKqN1yctruMg9LAxk9EEPqtLmp9DNuu9fgDrwJap8sh
AjOtohOx8m6moceX/jSWhwF+tuvN0BhVbPyIpMyEPpulb4a2ekGiqHrni4m6k7qMRIEMnDFA05Wu
/kln/1aLNC4AZj8GFSqfIwACOihO3QjlkMXMYF0T3ESOuuPyg5wYCQuklhWrThhm/NL0ATzWqgue
UnwCC9GBlDKdZERY3w47NOOBXe5chAfEFeK7HMs1wbmDyK6TaCBKLpshALqwuEBzQU8SxvvKI4xu
DX7DxhmoHvwxFevZk74rSM/ANQEnJO0ukcOcFg9kWVuJ63WDJgYiFTq+Y8dyFmUjKXi9JqQvs8jl
nOeGW7BiUdie0LfK/a01/StYCgCD/SRGdNpxKSHLBKLP+hsq+319NWNLrpHrVCjzOcqTPkt+Y0Ub
uIlQoDInadhvy1AQ+HCQr11QcoV+5WfjpPFlmBaf34xidh4YylRRH25O46c2LkW6Gd7i6xBS2OqS
Z4sYIv1YML/0JKdkrqsyoBxWIEKXlCYUVJB76uaXCYI+Z0d37iuc7dptl2MBZA5PVfODTQbPG95s
q6QHyKeuokDng1FYn+P09fjzhwsdHtXqPkx/y5xL2vUdaeh7+6tp+nXvSHcfdf6ra1Dpi3KYeoBe
Epmd98eN0FDaLiWhxmuMSuZ7dSeD351ugorXZdo20d8ml0OqRZPHXd5qVQRJDXMHRYuLVQX1tvPI
XdJuvT9RfVEnCVX84PMg6+OrOnaFlUk8J4wimyT67seLd/Uvn7NSfKEP8CDbIq6pevo6Usw9pfPR
Ittt/vKZ4TGu1wOil3VkFHh8Sn8k3Kx6EjeP6fD8T5u4BwPhC9qNKHwTyXq0hivRDMDddtAUB/ik
qY3/9bJ+EAwIsFRItV9h2Pbt94C+KaMvYuQAENmNfQNOcdmiXBUpQdPByCgiQ11axxrFtumlUT+8
Ph7Z4K+GohAW5+AsMF0Tb6FWtOdi3RjXEwzn5frzCjZ64jr6NbxxKUQutu8awdfJvN+E59qo7YIn
k1IZbGEBmsPGDN+IH51c+UMcfuHZVM/ni01irU6hyNPlqU3Thu4ma9mR0g3Df5xBPhtKhs3n6hG2
Fce5W7PcBmeskL/p6fmRYHmWxsxDCRMEs3YY4G/pL4m2oBe85ntRwgWzmBZBvOHhw8OiUvOdrPse
ykoRy3BbuDviOw6usthnoQ/hUOgUJSP3MUSxONR611Lf/1nCZO1ZhznBqCH32Gpqfy7guhKg7I0W
h0QHUQpp12RPGI4kNKJFpPeQuIw/7it17pVC9fKGlpiqqXm97SV7lrKSJ1TnUvhnswstPeXxc0CS
F3VRD7hAYfgSFfK63Z+qmY6owAKNlF6M+CvN0iepmUNGC27DWJnPtIieFMuorz21o5MlUS2qjks2
/86G3NumtBKa7Fg1P6UBucwxnvexWrj08nCN5O3rLgjgh5gPFZ7sTmWuWpvxAPWULxiORNirBdjc
pzd+vGDvAn51xckZstefREXXf0HwhafesyHUEsq8jnz177Nvx+Q/h4+E82XSe5Nm25Dia3EcBIbt
40aNH1yZou5FMQnZI2glCtymySgbrPB9yiurlRAgrnk89nsThFrLGd1EbZq46x5slW7JWIMNbyPA
xGVkjg9PyMKYVYo0wkwOBEIWiHPVN3rbYgHUvvHm+ZnVX/Ndu08c6Nke5Gt6/Jlsftonij9CtbP6
4zQ4Jdds5eJgItSgiTS1NcIxcXcYdWNUHSuNrl1bnyKmjEEy1/DDGFLQ/OqXMhkBNB2Uvqtk/HMp
gdiLM2VA4gceyPVGLkwZ8+KZuTYjofeVnClZF4Uk3Pm3ixDsMwPz6+w+7R1vU3ukYKQ2kLckbi/Y
iip+UtLsaFdZMrpZ2IlDQV8AtUc2EQvSGUoSwI7IOJewcwNwV5HapKeb3wai9PKUuEAKSCTcQCdq
DBne2GC3lKMViCXzs4Bv0gIEMZTkUUJoQdl8pEoiQJDHNauDFhxUOinbKkWA9eEivsIVFGKBJiA4
x1oP7gjOLkkxWcOsNAS0uTDaii++NS76RkcFWS8MNrczJzXPjb8n96y3f8Z2gJ3xKa3dLHIzVKdI
FrJ1XwKhgShW11KpVba9GTmB7ez0Pn6KAsAxmAkoezsPzcFKp3ZYHfKq7D066e3z5LCFFi0/zVC5
ERdxAhV5MfQ8e05eTloEBl7cPf0MxQwW+0EuxBYxeBgCA/aEcwXf9vBJX+b6RRjbi2/WtO9jaw5r
znMs4eWGfndUT7ZHn/t8TJlQwM68JJqiFA8U5HGFcm/Y1Cho1k02imEGl63pLDNhA4/5Xa5Nrr9r
gd19U1qwhrnp4YOjsyrRKTA2jpz5FSF31cLoVPn5gSHqzIqjA1osp4rNZAs6gTJBCR0DD6721v4r
0u2g5JqqiIRClMHbvkxjCWZK7Ac0B8ZepxxPvBGFijLSj4shDmoTiyOn9wxJVE3rQ0Ckym6On2NI
ol6p0mmEd2I01/j3wXt1B5MQGXFxiHSB19g2Ap3yZ1RPyzoDRqsjlJqcdZYxia7dmLSvGoc0DLtu
soiUCn3CMpAUeZs0hUhBlOj/7OlBRGqF4vv/QRkjqJwEQVc6A9TebyvuxAoLZw7PO/kGPwthkND0
prkbNf0xybu+lzHyBm4+l3T8tDDxNvNAp1lFxVl51kpzypa162ZwQHzsVbWK1EdmpAGuOWpzlIpp
GQ08sJBxqAzfHJsyuSEQjhz2MQy+e9t9ruNZCo4T9FFqRQ6NQS/WZkR0N9Uzqe1wjl4jivUAtmZH
hLe/dIkayIdxCJoUO89602dkTf4NoNO54hHIGEju9F+Qt57BiV6vBPV8tQPk7rPVbpaIP4cwLGcX
2jO7LF5zd60S82/zQYv8w/tENPx+rW7EYuPmklUSVfcEHGCjKiDWMRjzh/Z50xUewmUSDmY/7eQu
cGiiKeJSv6WuQVjF5MCQYJhCqVAF9oeuLNflbKuVgmRBkz23340TjhWE6kXsqcgk7xjKYe1Aahm0
RzgebH6PHRE6/yiBWTk66C9PY8SJd7RRz0UlyrdSoUK5hCNUvt7B27lrSfwXcv4SmM6J0o79YodO
lag2Mir9qGnxXSi0rCbeHtCED5QiJZjWyCPZj/xgqBzC7v6Q+hpbRMbiZWtFRTB67OfitNtdXx5N
hxilHhrilwGV2/mnyi7r7CYVqVtlPlNJeTN8K6HZxoiA6SKRY7hRx1RPIGmnIzxvWIgb6kW9ZktS
FiXPSmTl4HQKbx19Da767hJIMXhJpxCwMMBpGdp16/QF9KUBWcElMNmhNgUh/8YsBGHM7M9Gu1vq
LoWQXWu85N5/Yv5Ztp/3f14pv/Fqyj0vRVBdS3ukb1uqY1ShDEHdifyIcm0Nrb1jEtUwMhRtC0EY
KmEuJfj3xzYoY9ASEl2ejkWQo331xmbk9wF6pY4eAZT7PHxV7KiIx60ZxcspqtW02aWuEmIDLBl/
eDjoFivQW6OG0g+1jHEL3sbH94x1dJU7gLlwEJgDBL9n79bB2nJQmw5t6qHJluS9WrQBMPrpvydv
ys7fSrS7SRgh8BfpFyO5Mxr741rziXuBQB3lXPHemZbtplseeuBR+bTEMA8DgcBPU0uVfr1mCIDP
FayEuKkuwrd5soaIhj4J69cAk0RF2sA6SnZiNVIOAm6MMrb1qf4x0xDB12DVDAfa8TnHBG/JLm8c
DXvGCw+kiHx1SGf53IYdNxcjoTkTVggZU25+vWeSrCc65Rcj64FuUmy7NTu83WoJOI3rNXjiNGsU
cRQnSTomEg1khBLn9LCnRuyEXqI1xA/Ywkz0m5YGSaSgNSBVEm8NmYllJg8Ml71WLsWb44XwnXbz
6BVY6TUwCNO79/9KIhiP8NicWLmGU/Ju7rox0ii3Wpd5vpUR74GMuSGNrn1zqv7SFMC/MjwWJwIK
H7tTMW5yVnG4XK/JPFJImRbHdnkcC9PsbN1BqcQCShxKHHrSQRjl68EmogpX46pxn3Qw5ZpASBNE
fRozNJXLjddsEbRnFCXF27Os2M7O5RihHfJRGxQ2qfmizFvC2f7rPZgrQZuJhV1hIgheEHKCzDJk
BxbUuq9IZfDeHlRBkAjYQ6qXzP6yiyKVGQh1XI425hELn3yMNnC3v0aNUpebrpWsf85ahYC7c/k3
nKCVdORl/3twhzwWpZi/ZEq6KhZQ4VheafVYtVpKW1aA6Syj/4Upxih6gM+A1rzwtjtTLUcAbN1R
k/fVJ0izWbYHzcgg78rNKOQEtSFXG/RWl4vxgPdIiBGAmThdO/Gt5NIquS6PQyQf4JMFug8PUn1j
+qkMjd1YsE9Qvfb2iGCr7J/yEQ5oRFSB0qmHquN5dJEzf6RuUZtcv7l/Xq72+gFET2HDK9e348d2
h4vTIUDylyd4C8fPWaugBIJps/KpPlnDKeg0MjwEh3DYrd4iGD7rajJjU4lcHpVEbWBRYH2F1EKP
FK4ovSzs3rPiWHuB8bInR350pmOgK90anc8k19x9XBN4VFls+DMztNwSHHGH7sOGiI5LSq6+WC8F
T4fbrBryzmaRafmiIyErmIP2Cn9TkX4gvpT3SVHehTt8QUhrtsQlH5rkSooIFMoKQmg3HvjSRgLh
WNf/Fz65/0g0diL/UkQ/+VarXsBzEJoTdFsdB+4ChmE2XuITkDyw9bdZ/Y6q16XAQEFo7htulgki
Ijwrse4SEkWfg/KvfgH88t0eD4kJjiitXnSvWVgTm9UosLuCapvourAl86vviKnsrg8L+gmTA/er
8mBVsK15Ig58J86KNTBTx/PlGpjjNgcLU3cnSFTPZp+7ulYnDWLulaX2zc+VAC1UqCcLtOopj4zh
yOA9taH+FeD8oz1aGgR1kxNi/TVWw+GdI8nJjMGwWAqjB7bT+gqAVeIx32IAbPsyyoA4ffLl80sM
B9R7ZUoCHNk9/KNHtPRfXhL7H8sAIk7PEFaKmJeUckTfM1vTp9AZS4Fq0oGcEwErQ1g8XhZauCFG
jHT3GU3xzuRUpXTDrLXxvcG5P+GZsVGz0oFIeNtlRWgteP0gEH4ipnX6sYEwd5aI4h3AiJTquqW1
b3/UpjBzqOmLR4/hqjxg9sM4yJYAc9YIu+aOt8ubgcxRfwCcXVqs/2HOnX9I8p74AY6C6CUnGGKi
fSkmJiFO7HVYgHvqwL0NEqRVF5HxLIigP2xoTVqH0i6L2I6XpSJXvgqkmhp6aRnV3M5b9fWurMyr
SBf3OMUjUyN+Nu9eBL71s9doLf4gmYPx55qy1tw7UAIZ+nucz+awCydpnTk3LPPkHtoy0wbvRNLo
FD6T669euxSxhxnOi+wJXmGGDOAOoCFVjdJ0VA6ZcjPgHHMzBHpAQBE4+oJGxOFkpk3UkkY2oBbl
nTzB09rU9JirVPYTy11lH3a8UTaxvSjmKOjq8O+0Ssz/DpEv5HFyoWqOA+DWYAWHPx2OYO+zuMxF
rPGg4uUK69U0AR+WVNLFSYo1ueMmK9lXy4LU6hZYjE0XRdgVdLif/8nkqHjeAy2iQTQdPaAUIyD8
5RK0Rzrz2tWdIem8/51Vs0d+xpCTkpTyhl7QIJ2F9s+2hpoL5UBuNio4oh4oKUdxoPEeREyp0ubH
jr45cWCc/HK7FnbFsxpb2fA04g8VdzbEFCcE63ayua6WVAK1+2ODjXiIeG8n/aSvbLLFVluTV5Zf
HmpJkN92B2X3SBwHySGaGWUaf07BG/to1uGFVAMupD0VQeZWGgwNvtkoOkY8d7DKQEAwZWdfJjiP
N4l31va2eM1tdTJDEELxazCRBxktvkTju92Wi6biKGqOI9usfmmvzbPtMJIVGtj63isoiMpO/LZw
OyjFrYguImByOh2rIjm/JvFlT1qt71jnn2ZxjYL78+CqbIbZBfUvUztwL+vv51RMLW90XQqNi68C
7ysgxQvG9wJZC6toPWgYnmYk8ae0cPLRDOzaRNaA+t53TPcyvSgTBmdP40eaoePDy+2CmNcWhUWx
GcwDp6uTbSTK8GaKK2a2i5sdmLjGCDEu4a0Q5NRhteVshM6CkxlO+Kx6E8K/6QdDuqCpulrv08gV
F0EkAdy3o3IXamubglK7E4w/XNgutopzhaU2enSOiNd0buAiNKordUcdkSajD8GEB7TbHw0MUFo+
owRpySeeLtcMor6A5SWg0qicNHFmBMz2RAaFSC7nc0W90FokaLG9yVPUXpALPsfqiTa1vegJ2bJu
XZQiL4VXPEJ8F+2fFC3+S2vNkoQeRpNvdtk9MAb+ty4Ip1M01dxTJzicUZEdiovjt1zJeAXrGC5n
4/0OszQ/lKrRsnAPxQUSdANGikJnjrDoQfMmM55ko0JYopa9fbOJbyHSbfIIdlIxeWDYRtFaWQ7e
lE0FaGQSIETDXR2tutGJD1E+8Wfyj2rQvVEFVhuF4ALJZhxJXA+9EEkRbUusMrsbGfP3qHnh1NV0
u38V9q308N1gpSvV3XrhscJGhSfB5Ry5yoL6cbaaDQVT+NXJWMlWya7NHOrdi+QOOFTQf7TrDWHF
9VaBomLv0vHxshmYRQOYquKE8/meHTXKnPYsrWPmuB01Juduc/SQNzio1Fo9MD10GI4IvtHefQEY
ZeoKY/JFh+qRv3R++MfKDKuZCeo8/bDP4y1Y+PNlJyw24hRI7KywDRMVT+s7WGnrMZrwM+4+QyVD
BimnPIsAVgU/vEL4adzkfC1MD630ah9oYfROMQOeQI7L/mIrReNTmJXWmG7SvHQED6D/mxari5Qv
tCLytg1GNmXEYZUnsfmxbV9idipbXpwVUTh5ExTfjw/C96/gBSOvzHIn7CzHBqanl9ylagpd0KNK
tBCW54kH4p2Taj65OAR3FsSU3aCmQThLXU7ESVW+jONn3MxO5RbB/Z7CLQBmY+ZebWfT9FG/uB7+
8kSrtsaSmYg3TkD/U3TkaxDf58ef63fRjn4mO+km9kuQXa41KG5Kpc2CWI0mqJI0oHDK5y//rOrm
g927KXR8Sg5wcSWaXugyIof3Dk/qiitmbo57/bl0hhc0F8c2eF0UXa5wOlL4mNeyQE2ImPICPFix
707d7dabPT4UHV1vagoPLfXwXxCQ164gMIhQyz3foaHrusrcg+8BuPMyk0yDDaaLylmKUN5382u4
l0WWLeLLBqmWRSLOFnkhljAzZYXJ+wggCKLCvTf62J1pQl336/hE7dQ4d6Y/NQ5gjyJeEQfb7Qr9
8EwlZCcqJp1b5iJlLMOyi4fMZhUrQstzWVywHdKRkj+SPO1CW+pnhPJiFhM7M30CtWrYpHaN0PIz
odAlhJBLZzIVBhMehuU2DB0MuNo90Va2qWbR8VZpYyMo9XIdpTYKzL/QuS2OmWuYk+cA209AE81O
M/Wsn/BmeV/ykQkcXjoQUbjPlj13rujgEW+QzhzEp492a54SdY3ZuVUNnfXZqtHTVDLmeBXveD4o
nIbPHdwUL2EtiE4sWrEGnfhXUagblhDVXZWdmx7Tmp4nQCPXjj9yb25XiYycvC3ZobMAN8sxziUC
ihxhR85Da5aHcLAP1nLOYMjz4qI9jaMVWZctg1B4DALeyqWwuBFCQzG4Am+16YgqLhUCfjtqhAV2
0zurJ9i/atpYQoDvRE84b4kBNFrpKKhUqTmUMeoXo5jRwe+X0ltb8HbTFfvDXrN7OiqOVJCC3bp3
TU8OOENFhTD1QL8ds2DtgETUk/F5KDGhmUUvFXGa9L4nUrBT7cMcN3myW1F2Ca8Ll49BxAz2806L
2WqfCL0+g7By2AMqHBjGnnOHNzcaTMONDBLsRYDJU7YRtef5nw+tyAWlPKcmudZiQOyWuYvZXCBv
esJKtxzWzrYE9NvEhWxT71nzHQKopx33hXCz6tR2P31GcK8NcA9D+GURw3ZHJHj6F+OIBMOZPzAU
1pNH4UMXLARZDHIdUXalySX9l9RFrGMpDFLR7iXWeiefQOUiXNYMrXchxvn4wTR+dMKU/J0x6Ea9
GhTnfCwA66JnYrw+soMU2+lrPXmpGBbcV8r8mfNlc9JIWquWn0SftoCn+cMGAc0BbjC8WDsSAquc
fEK9eD95kc7tA/PDY27yOJBIU0oG/sxZiz7Od1Z6IRzEHwtV2iPQlWFqszFHuPkPBTwWVrSN/XUS
jAv+QGGu9Z6sXCy/JJMzPCsPe21HdjWYMn+XzHCtyMlgyOWGi8nmY9Kdla/Cz6Qnb3dxnFzqoO0t
FTb19574qg2SBU7NJ9xFqwXi98jVwqikFzdkMHaSHGsuJ/tlCaXm/xJ8+fVODinswHnb4w+MrVes
mVoA9dLnJT3U72RgnBsX0Ac4fWr8sJXWGEttoAwsRuymbZnmtpH20DiRPUGqP7fe7f97FrErVlKx
Z31cU0X2NB1GaggyNLd92Ka2J7SMlpVdFbtZ7KwYAx0AIvuF6rOce0Ej784ukF3oA7e91rUhWVsY
zZcDL2LrKLSw97jKFcMJ70Rx/uGfW8LUk3N62ScIpE0FuFz2afuGFMAPZOuOtMoh8a6SCrstB5s5
+8AjLDSFtkKCeHSOQw5Qu2voxK1GPWK023feveVebChBEuvDfbuk89dQ6tsn/ZTDkIR5iqtWNDSp
+75e7NF6FBxctzYXB5W9zpIylGjrkuiGhp69LsJKFXhwxC45aBT8HB59YMw04r6Lq5suygFDkdY9
U5W/y5Jw9yDCa+O/xWN2IZqKrlaETdggXxs45R8jYlHdLxrc+zurSy5OSuMi4Da2H3HgTvs4c3Tj
P+tIdfcYuJ/yz/1ax15F1iu+0p6Fyo3v9yVEcTNaZL1QXqO1Xz+0xHcyN5ulOk0hvoG6/JU+pAzw
N06Z12McaK3Z0mSIqw3kEWRNqNO4lRfH6eU3U4JN9RSNgdfTjH6JjgBC6vDm4MZbyafK+bq0i0ci
nKKI5c+YWrP43YjPc1WySgwdi90sPrtGFSX029qNTecuc1HffPYjkRgw+zvjOtJtzi3X4ABk8SPz
YIUr/XTTvJb3P/f0rjOcTxRj+MgHrVdACEIUUcKs2SsDAk341NfPNGWM8Y+EYHiqGINvJqNkpxO5
EHS5zWzUiyiYNqJWx1P4SUNluQ3gTLIzH3IVkgj/5DHm/d7fxPVbnlEkSqWcaCFQ1FK24/uBkq6k
pbM3K8rduyUn9Y1+zym49gmTL4H1CAuXofsxTJtFfK/1tWlhrjRh280X2V3IDGXWL2na4IH+LZt5
7PERCrWpyof4jPI4ZlV69Vcb2FmX1wH4lMiJUD1kUFLfvrSlTfOHiEmS4DrBBkztbC9eenYTL/ka
kBy3eUIUPbZIlxCStAg0YieOqMApYHYNVKUIJ+sfw7hfolCYwPVHv3EvHpaZ0SevUQPkM8esAnN6
bDUeCUYpwrxAyXNbSaiVc74sXsm0xW8sKWnW9xCOAYDypa0b/SbiOob00evOccosxvN8wiP9X7f0
cdmKjC2JBMUNKx+pLKP/nFmTQb6PHvGhbT20dU9eFdZezRtfa2Ko83FcndniwGBwSeK5RH8F0K/7
BhfSIEN2EBOPkLrMXr5jVr/GhjXJBJRQsE7RMsnxiSwjywZ4r+vbk7ope8T50Xhnl3eXUJJPu0NO
keHGVIkRtDicBTT0b1YMAXp7Pnl+AY0Occ79cDwzRRAdD7W/Oto6HwMZgEqW1N309DzVLqS3DPAe
NAgI63+iO8sagcR4KHJXow0FZ8Am6S6qG7w8W6RqcTSpGgHvF5E7u1OU3aLkIsS1x9/5y7wzS4OQ
jnT6alHQbIg/I4zl3Mgzcv1YhRLq2wR3cVVzxLmzr8YyUfMI8xU2zXOJnpM0qGrVYxh0ywXmXJkN
Y8bK9oAZWx9v6rDXB5qLPrNAnGPup3wGmtBwEm8YIWEs5H/9xXrf4qNRGnENasqLcSTiGxs/cQq5
XnVa53fPreGiWPPFdYxTdoELeYJZamGVp/O9/A5bvEiBxN7NnMR49Bs3e2RfAUbr8wMGywSOeia5
EdmMDDLRPLDxTsx5X+s5pqvSkxJBFZiwVWu+NMKrzRalRMjvo6m3fzo/qeMGbhEQeDdn3UBe6I00
g3S1jnofdIYi/fp0zQiTH5s5wa9LfK7q1WM7wZjTDRqKrjgl+9uDBXHLmt3k36FOD7S/v7wWpQCl
F9UjSqOj01+9LOc61jLPH6rTIzyfMVYdRA72WCnSMEkFI0zoT4qOaRCNo0CC6CD64oVm2Dc/5bcC
oHM0S4pyLytsZ14cSWn8J8SDcDV+5nlJyvpXGu6up3A4b2/z8YjlxAFj937e2VpIgUM44uoc1jpf
Q7HfMem8zRejESOa8QmUjIUGcx65cs6WXMjTdxgSzSNCHMdIEAATvPrDLFWIDqYy3tQ/NKVxBFRk
UxprpCBMKPEOeJiLIRbXxRrDKwo+qYkATrqhJ9+b+cGSQCwRRwan/DM14T/H8yDxab6QACr6QO13
P4D3zgTyIsmPjpEcEH5nv3BBjEOjyfS5UkdvbgvUE7hqpUxuvp+9TL+mPIwfxmsyvtDEbN0+Wy8B
NMFhxFfUGwQfm8ycJ3MXWLjYtgnSEO/dB3ZbU4ItQCwtJ6YSKzz/4PyHKbo73JuubQ/cAw4Rj2Wc
8nzE5L/GduBBTsxPzkBy/PL5MyQXPsf81IikcMgmrTVbNf1BeZDLyLsPtTTBoLpb7aiTJa4tWIGH
sieMViY5iLP3B2eKFAdGm52vqQ3ImBcSnFCq9KJcLYYpfbH/6etyOhIqtr4XP9+pj3fopxprlz3S
XMccJTcaI21GSOLSw8Mju6sHeULvvqywEbGgjzQQIleDj0jCDZzh12B1SLwwJ42onX1G9DzxGo5y
ADEx0ElEGBPtoBBMyg+IxKpJyVcF7TqtHOnuFy5+7IkIW3j5y1oCGG9DbzWUvhId1zS/5e0pY9lS
E7V8DUoBOKzmaqSDFH0E8fw9BeMM8vRcGjFYnDvcv6ZBnT0e7jOVOiqhgd13R+1E5ECRVb267hF8
jroSO8YvtSn6ZIN47htFH59ok17LQI2cc+F3SUggz/8Awp9zA8j20DVHgxOF2u043l+g//tWkEBI
uB9TBUxCE2+WxGjOh3J8uub9KjR71aNXv/X79lVOzYGCr7NJGvCmByPFIfNWdTabXknuS7p0PwOz
EYBPl5kecKvBeTzMwgf4WUQLxW/zdqOsRUKDd4zWC0WQ8Lg210VmtcN5GdXDEvH0dLYaQmxa7Aa6
bK8rF4EqFw3r1GOYpetfcqeSh3Pu8kPzjztHAXL895P7UDHAu5Qoz5g6EOfXGdtV03w4zWRkitmp
MYZB7ciWfWZugk98o7uf3RB3cCcZ21cxTVWpj+hdPo6wLWDXO+IJS4y+P9YIB/61uoYJMzZTA26Z
UtS8Lrl9Mr9AgIjK9w21+nr4/NFgnH2r7NpT/OP5NRLiU36d/vivwBoOF5a/CwZqmhzBq0gAE9eR
TxyCAsvnut1mrXI7ghayBH15eziDK+NmGOliLLkFXrAiPjk+9r5cMuimX1mba4j1FtD/VI6elBR6
mNkkf/wfg9btvgurMJ5SJDLtobjaR7Cqna5+Y84QfwHmgZAXfOTKakkcBEMBYbQx7M8Tzt0lI2lJ
fab+oZKUIVPdwaDXC0V1iUq+QDejrJ9bcWzNASlOemTC7gvSrt9v6jdM5L0Sn04wvyH8//qeVji7
CE6r4ioL/rs61N4YTRrgQkqI6DoxIB4WKmUzypW8Frq0mrT1YljhWQmp3rt7Z+Fv7NKguwpG91dz
GIBz5KZcR15xQf1Gdb64dRybaUNgkw4mMQqj4infSrCaDiSWfHZM6SgDZusBLYLtWrdv6SwhaKOk
Tn0GNZi+evnhKrF/+pzYrwNjQmdSHAOHTN85ve+ITPSlQ/nQJaQBD6Ahg4nMC6Jb/eRMXFz5Iho7
oUGVVx86ybzkbRo10Hev0Ztm9rYfstygafLaMSZTTAh+M8ans18mu/xmpt1Ua3o99dgrW46ih2+L
NPoEuymSwD2AzQbh4rcMqm4iNNTUwPs0KfRCVuPhIHoy+JZCkZLXvc+D6gNBsIYCbaCqYZrx31Bu
aXRtrFkOIo0LmAnxe2bbmShW16V8e/sAvhrtXBk/JhLztUMH4nhg5/z4Q/gjKsyxT2576CAoUkYB
d53KWh4lw1fMuODb91RRFfuhQDiP02MCsqjNLjPkqMh9y7Sbr8iDnRsXqbsRZWfKv2sA8YsPS7/X
YaXctX433iisDBEHhgF5loYHRObxWivIyADoY3Nwaq+Xt1e+TgiIBN1Lbq2YpF3wrzQPQJ0orMDC
EZGiGVPd2ETBNfTt6tGjs2jiSn9mlC2CbBkWbVrHCp7BJ9s/+YZmUfwXqsEUnPmstWHTghumbrFh
6oJstKq095Oy6ilcgkZnGBi0+8qqHSd0Zk6v/Et6QJbY7nM5RI4OytzjdYZvD+ENX3zxY1FmQZa4
+c2DDXGYOrf3G3e4lVf9mYPvxjD4OTNrta4j0CSX1zpl5o4N5exqthTpyyaBEcHz7GrMryx604H8
UVJnLmMWmOjACWLjXfuM9klfj0c2rA5YFLhs16MmLnsu/I/THTE0NGarba0dm0my0ds8hJ1bd1aj
BMXly/o5CtQBQpB8BW4DysbDFJiGsdk4e4CWe/OLel1cBIMiSeH5pR9ra5yKRwOJI0snR7cswCJd
9skcw+v++Cm8bvHlkrlbzYIp4ME5M/0T4tjYBtF8h6sIXFeTNCOIcYIAz7R4O37UXfwxItlzBeUP
cnNb/6Wx36y9Yho4hR9bag0/XcknzKX21jg0JklScN8tzWEw2iEy26Bne4iEtKVTudzB9UpeGv3D
nOXNwp1HaJtIzOS/APpSaWn9Mq0dwaQgs6JaJDOK0+3+ojz+3ay98gHpVd7yl9hMne7/57tCYnYN
/8Es3l3bn3fciS9vzBE3yZ6Ob2khc+XGOxL1o7K5Zfsx8L/mS0Hn+Sk7Ne8Gqa41GSHVOBg34xtZ
AYzHeYz/VvBJ3cp/OMVFA6IHXJyJq/EYI3tu9yfoRadPO520Nl3nSZop5eH2U0DrfQOwXV5yYv6e
lAwHMxXxq1WB5LMn+Bha7HQZMEOnKlmvv8c+aag9SRyQYT7WBf7+HEm7G2vjllTyc6XQZkPyFh0G
frz5aKvo7akir6qWjHvQmGFJbYwNvrUTwDe8Z4W7I9wqizUoQ8zQJ2bGxhBzyoBRb34Pe8N6qgby
J90WBunIc2qP8w1dFIs3jVRlyVPEIT/zryOXlmQa2xeDcBJq4d6aFJbcippBwUDiZOtXo1EO9vsJ
e9fMERD5e1rukVY8WuW3PTpTRzo+rj1BUQR8wvwLXqbQrAiWuTm9LY3lsZvSa5frn6Dcwb5TOQFi
qlyKZEqdCiL0tP8Fy0zcgSgamyOxXgd/WmI3RPDsVbuVLMaMq9Y45DlKeXNFxez6bXeuYtpozcDG
vE93Mts4bCnkunMW3J9lQSng9DUGZAb/0a33OVkKdjZpk2FpMeYNY2Kvctyvw/rCMIABzTcilmU4
ZSKw9UvY3UG7wLatvdb4t1xxXmSYs8KZgZm0Ml8ji0F3jmSFpyYFTcYc0gxfV8lgBCxafsPcbYt6
+M7OwALVRreqNuVdC7sRPUqhbT1R5uxSW7EH5bE1kAQ4Co2ec4rZSDEJp+a3IJCBz2c+Cwy8JFk9
CG7gnI3P0R7GQmXq+oLnC/mRySD94RRR4kjUsrZY0eWKA1OdlyRSvhgw7PNmsgndcBQ90O+rAnKI
fTMSJb5vUGPAKt+uR6T9R1BKa5uXkBQbTmnb+nzdAKuuvN59GvDIGj6H8V/ZXvxSH4LVehDES9E0
qur4gejPOwBfXRLmK0qlwTn7+7IhACODwTIcEMRSy91ayqq1CR+6Tt3o8fIhVZiVyvHGbKGOvqO1
kC9ym2+rXXaktxbXSgbPR1HwclZ9jyr7T/D2pn3foFSaY1ntWwwYxpOsQCNQkKY3tlfILOIQXYZz
Sia+Rkds0lBS0jdaxdl7kG0r9gav01TvfGPc5YuTqM3bwBhzVlqiH3bGOIB/4xRdFTs37Hrp3wm2
zPGiWwBGMJQGqn6JNtLB58JEAw5lnQTbwVgLbF/AN+ts3/jCa1fhPSmQtozgiCeuWvLZ+//d0WfN
fzSVIOCBcsTfKBRQuJXILiXY4ZsKGq25HMZA21At8oCU7DACcsyMNKDGBDUFcl0eJC27EvCsiwCs
u5rj1QLHIccIwt1USbYb4H4GHnKMl5N/klIo7MNLOOgjxoaARELCCcPkH1Y/mTH34hShJjbUCP2P
cUOnoYr8vET72Uusxy8H7sRUy3ci3w/V0tjKgwE3W+SVkS/VlrUqbnYCmRvESfsuEF2F7/JjyhLq
STfn+OjdB552LrzLTEFiqGx+LlGAmobP0Cx4wvvQ7HMLFfqNRy7L6+vOmZHqILkj68AZFkMbl4jw
QTH8/tESy/cUTwAwodvaRmlmcZEZbE9XcIAkOkV/soDGZnQHcAxEX6azReje0LIXJ1IvKtBpNWG6
tJajREIiQfK6+yH9uCVd1oGAwXagczV6nYHRcGbQESjodyN2zqBZ/QVVMsmuVY9zBlFWOoXuzxq3
RR3pwbGDpqP1HUixF506YXjWp9QOSnpexhkOqwF2b+fLvBZjhrfOeobXBOFLOY88QFCT+ZwYq2/u
TYnwVNnR3lzrbE1NWgYB0vivCU9pEa0I2ip3pj09tfdkkmJssz8/ne0SOmNv3MXZHSozl2KDlpTs
k563Api5uD33U172ugZGli7yKyhTXhtJtwOdUL9IYHd5E168tM7ju3d9xHfA36Ui6c55+6utMc4i
Ca1qALYXnB0qATb1xmm4IdMxIySKdUbzAhm7SaCcWan5GWi2m2EKFsg7LUeOYjp+U4YTeRaKVPs8
mTZ5oeY0kofrU2ivb6gnKz+c4cDueJjJI5+HRHQkhCwA/CU8jQJ5nJmHhCPD9nxu+Z1IxZyGEaIF
YEnRxq0nmsrrx65agYpMGI+DHCx0vpZBGY/XK4fTeE4FMUnGxgYCLkeGKHd7uDrmoMaI/eNunhyA
DY7J9VMx7+70JgRm8YqewGaSbFpShLYbTIGYOy9irIw0VQBoaQGdbrOIVdpx71MnokyrRbw2bLL3
X2rjXdFjYm+L5/xaXm0u/mq5tIuw1NPAtIL3zUN7YFMaff8ZFE6EnL0ZUS1xavGKETFe4lwV4osx
P9Zgd2lZ5f+op03DPthdQbznyQVJb8rGMJnCZl5jv+SIySIhiLUUiCY4xnA3w3j/HUFrunwh5W0f
EAWK3C+/OFwzX/gTM+iMopaZCP7Z4szKZRrGtR6NlXU3qvaFu1jc/Yx/xzHQ+INHF9btc8L3uznV
Wv0Z3edjS+29bsHcm+ktUOvx2XNS2d1Ex9ofvQb3KLmErshP7mnWmAIuC9TT0t9kExDHZbiyImIM
Uuf+DThrPfSBIv4VcyaFPGpJXsmORnsLQcDN7o/AWfW1447/Lornz776ck565ri4b0VBV/G6tCzZ
HHyDaM8E4UF4Q3BVvcpAW1Ey5YGn/UqEwlu/hLg21U+ShVFCOM7PZlEmfNIVHDraRgymvbztUdEP
CoRDGxR7o4WsXFRycNLgXM10JjhCMAaRAYw3KDDaf3zYKbVWSsmqrqKLZm//UEmF2l27woBMxKNQ
vO8D3I5c7xWltWzsdbmP/wCHrf7yHYwr0UqeWsNa9cetonxx/va1fFR8W8qtkStqa5l3FvmOzvP4
3Hd66UypMgvUlvPUN905Q7spR3ktWshyDrmad9DYkqnZJr63qp4zfA7QljFDsB5/lWYGv37G2Aun
D3kOTq0NCUgi6n9ckqqppRiu9EYNEhu6orapdhbjPBsI647yphTEI8L6ejFEDgcIljuEpBP8kzd4
FcVzP5+ldbvR9tr6BehJ3c2uzpZAcVXbLMHouNdDHHBH8Bc7rw4klDLv7utFjtxY2TgyLXFo9WtU
eGsJeo82ZDxlHmN/sOcsAWjXyLIusedkAKlHYYF2fmmIm5xaovOq0UKpNTZr3dvU2TG3MiM6x1ld
lZWqxt0zJ0+roDKFH7vzDyEVtB/FL1/DiTTffn8MaSnG07tFbf1dMwU6SxyiB5y8kL/B06wDiHMb
LfvGCd+q84S7T+SlGOS5pVApYFE7Y6fC0iTAa9Ky8ryT4CsMAIYyOwvi+9xiTBoNL6tYl85ubtWz
2volY4bSqe6RFds5fmhaITnBj4Qd/SYd8EZM2K2NI0/bl+Zf2+eCT8WBNQNpn3kaoqSbdObwi0oM
VtR7UXpZSdsdgUSkhkPOK1gu6VvgB9ZtEqMDTQgC4T6bOUSRB9la77ByCwmP5i5do1rZT+TYYZcD
hlhsjLd4eocDalRdTPCpX1U8Sw4USFTEfNAeoqT5cqVxH+t+EzbPr896ZJQ3upnSXEOfgljg0ZWT
caHzoWWQNv/H0yzTwtFPO46nekgUh6lHF89Df8ozIA1olyhMYVlLVbrD9qlYlNDuc5oV8MTI5yvS
UO/p/GWzhM9IN5+vcPaBe+MZYCi3B9M2XFykM/zg2FnLerjy8jgazE5PVuWaFvyCZ3D7gf0iM2YL
YqMYVmbgzht3CCP+5oRZlTRSJKzCQ3S57PYVliV5AYX2/aMdANiYfE7kU/cvWerMO49TNJKOHh1h
eIad4YiWvqFxpf9xoUPfOOY5e3LGN80I7Fz/E73ZkbXCBqyz+BUvfH0yWZbQRwTl2hI3NnozJ7h5
ol00XMzVsCNEKg1BVXymLr6ds4HO5MjvqsafV5f6Qj0nmwJvSi+ylQFMcFtykQywA+ckM0uBUoCC
ETDZCGQi09awmcmxnvYKTvlhs1QdmJtIro9QkafYNOYaAbooeSZbwVWFPN8uDoCtXaDCEp/ggJuD
jk3ReQIWbl8NhJHGfQUkkLUAkukrTceQc1tXj3r3pYQpo3OY8i8xmeGmpK3HtlUBd/nh67E/74vR
82uYLl1LfzvSxoB0EilGlA8cK7UBJOTZ54OyhImLbxS6rRF6Y56GEGkkhr3mXUczQ9gU3jzRDOad
znuwEGsxOXPoYKgWPtEG/oBvag3GZfQZs/1y6yvFiqKG1bGPeJGhbsacXNjggvONyly4KkaGl0sN
GNN3QVOIuG+QMR8+z8W+o943TMu1nJzu++NcErvQ/Z7wVhl8OmcbrheUvSSo8Ca2VxrdoCuXY6Qj
rqFV3H3H1vZJxgM1pratOPMGMS9IzI3H5wgdtjgBzLVKBDOzvpvzaOulzGxkKmQEmUJ8ftdpIZzj
M31EtcXLzn7NsyHreH5VIhXff2FRDAKSKxhgZNIonuBH7ttv25eoei2Fkfxgq6/GjuK3l4PikaGe
iU3WBuFh8G0jp5NOF1cQ1El4OKB8eOA3Yn0Wlbe6vP/zmviBB1+xOrAPsmdGLDndzBdnbecYQBV5
CfbqkqmbiTZCYP7bjgTy7cKXvwWHODJ+FYL73yeszeo85po+nu+RHh6WI4K4xlYgqBqqKqxvQrG4
OsC8B5JCNb5ObqhtfS6FOPhSWsuKv07WP292zEGl3+NgUGmD6Pgafof+OL2nN6aDOWCpFHtjFtKL
V3DAABYzKWVv9rXhO7rSgg1yS3tZYZVsyWCnjvrN/OmExaMy605mgx3jn6qtSTlGfUgcEom9sZDG
pluEtfWZweC6QFO6/eMenq58O99zMpkZzO6DQiktbLz+EZzkA/3XIghS1qK7hfmuh5chDW7ZnEll
frbE9G+nykflBEGX8V2NEc/QWfzlFUaLknFXecvzDp+o9Lk7SOWgo45M5xsEq15EnkaexxQak8pU
3LfCZC4nojpGqOK2n1/9pTRMctg67CCiMoz68h9hzxXluhAtHk8nql71Ckmt/pTePMHkvH8+J7Nj
SMvNu/weudJIikA9xb+jQISq5fLCReGtfuGvnZ/oTDxXUT0qW7MIgY3kCzycPb3ZYh6HWyzI51cF
KKIDHz/0OWyDrEgtpkym9KZx/b/bC3hmeM2DN5WwyihT45njIXR1WwOIOXCi8uyRRlmOEg1Fl/nx
uHIMzPmtup58RNc+gk53KEBTyGFT68tfXRy7m1AZjzDo7THP2RGiP6kLy9guvLcSztjdQEUBrAML
frsj4fmZHojAfCIdv4dvyD4eAt8Xc4QjuxbKwZtyMuw5BuD+2mnZRFiD7HXIXnyLVapL39gcTVMZ
RWdOjCCS8JBjA0gN88XUzfJzBbwOOPfkYhhBm9CfdKgq31GbAJwoBx3F6PSCEJYrkNjk3qs23m5e
rlfZEfk8dcAbC4bhlQ6QR/7JvzWyFVNCFuwqt/rGkg3Yxv8FowOYwqHErqciA39xxvWpPat8f644
q543mfX6CkLJ18tRzaWQM6DUV+es5tJsl1ycd+PtTWrW39fZn2fWZd/nyHdJ7yVaWUfnHfoh6w4j
zYUQW9WbwPk/UWTmzBncKHvj6CR1EJ3U03CSeK32GDXzgsVuq7QI2olQO2SPol858+0TT4ZsIK/k
QhiD+d+r2zJumXze74wt4sbgUikhyXgid1xL0Iu6SlLfd6yo1AYv5xkrmg4K3O3WGlJl2OQJqbW7
R6JWNDdE3yJD0H0USzQZ8xLdqhaxBp6kijLCsmmsg+wubWUWlmEEzrJ0BEPjnO75AqkJ6x6P28zl
wX6CxvMPt7duEhZePJc7C19uQ64jJl+4yX8/xmDPtvMPpozlFedI8KeQxnfxf/nPsohf3Fu21pzu
H6+3/6aFGfK5vc1CZwssZlULCrx+uMK+k7IuNZ3DibeZ1CFfQSDNjiIxwVtg6/OStM6041LQMrCK
ylYirRp2Ow+2I4dmVwQxsRVhQpsw6VUVhnkiB6kxX2BFKPyNaprEnmFr6wZhAEmI27Lrdv5aYpAq
KHgkqBXEqCgavx30HVeq5zRmCH/zn3lgT1oRT+aFihYTb0y7RjknAlnQLNYlq10Rlio23Aad0EBX
H9eRcyCq7DNsKymuGrk25UXQLPU5ZB7z7q4KdQacMQNEuvvVymH5xGA7cEAMriHyCmQqy+MWBvnm
DQYfh1nNTA6TPFS0ZKIV2bDMp0fz+j37L1AWr5k37Sa4PXA7yPUjKWtXDt0045+cnUqVPuo0RLmY
JcP9uWyXsg4IrQfx7soTLSVhGVwIEYfW5fQSAV+FjAToIecxhoS0KGybGG96GlPRf77y5I6oUKP1
qzxXWPhoQaCIVXmOrv+HAhkxvBMAdjaCabfJxsctKGlrbTYY1e4DVcMpYJ7Jn5vDgaH315hGBBXw
QYcPXvyJjHgKJLJ4vJFu3O0ffToqNh5RjLfaNWHB5ZwbsLXwKdirs3HlCaY+q5ke9CSLg/p2OjcP
RNsx6ydSQ0J1LuRZnuucbn3YDvMpx216eYgXw1GsiNSVbp8g0xApO0CIqgfm+51ywGN6VHGQ7F1p
zzhbgkhixyfR6+AGJalI/9Jt8CS1jgCFxXDSuDlRVmu1RutorEOUWE8DBT0YZ1863g+q/FdIhg5b
zBMaHOUfyI2+a3BX7HTYZCyp5SUOIKS8Sb+PMcVbZTI5Mn4FL1fQ0l4iXJzJuwCJ4B+dVMej6rmK
iUeGy8hJlEpcrEPhPiAbNIZXTeXzg3jU/ifjKDo5D6TVDbuqIL2WrUl/F87y0EvGAByba9Er7h+V
yHdyRLoiA8eEIKBFOKrGKSM3lsV1o9FeDZc+sGfQ5F4cGS7HrLJWuL8nPvHglsgHs5v0+by3zpbQ
GP9Ud81VTLwQxYqHVJIIWdPi7eTsivG/2bQPGSClY/CPzii5xT9NWpmojm8SRLLz+ulJEc7KvQvu
nxBITTotODd4aV4JgKjeIoWyBmna1QFDTDbHgGkA1UgnYWrAQm5hcCe5yF1BPQpPFef3477jtfHA
8C96Dmjcv9KHqSJ2nVxqV+BOirf46z6MCOaHaCA+Vf7lzYsEQZdrxcr4fsU0ISuZ8pSd11qpTjxc
atf2Lrg2PWzvmLcj2ALD5l5sloyra9He+2rf9dedTW082k+6V3/uP6qXqm7fuhtcEZl+LLBh5piR
+r9JrxTCcOeMboc27VbnLHRXz/ZB4+BeBH3qful0qf6y8Jm9cRJzMpaHSMI8CBiz9baxwcI6H3n0
K3R+Umo87wXBjIIX6Qyea3M5QgF7r32XsTiiRuz5yuHzS6TcfRqUt83vKhN/ugG47Y+UPnVzeesN
w9r29GoZgRqMON5qVYtBOVk+0XWNeuKGvTT3x2GOYPLs7iPoMqchBMzBIiLfYyxx11joW6FJIIqz
LVdy2MuihxNQw1jg+lSnjoUm6ItdB7sgQJNN3B92fyy26nDhyzLR3laWqKbvOH8V0Mgg9Pss03n/
hNg8PAu/8VRUt1HhK+Kqog43dJeKemo92SF/N8OXBBXRbTPjxxF/VMge8gse/NvUUPOWM2EjBG3C
3c7lkhubPIKaLCVEeAsjuC5EWSsw5UqSePlRjQfPGvVOy38Wclg/GF++IMLkhd/AI0wmG2XvwsbX
w5acuDwNB55sZ3jVtsojrGY0/z52NCO4YYzZIkczxhTc0m2TR9t8I7gv+78MnMD6wHXXyCc7UXPp
4hTgVl9JsgHl/ekrkKwR4n5sXIe9kq7OgAaBbSCqSRSA95P7Y2ijJ9tJyvkKe+JqLN2RJsloASoi
kdXO4uyU1G8o9iUpFoAE3yTxLAZ91ORHMLpbvGCH4kTmqHiZ2/+zsvcdj9gNEaehM40rNoYNznU8
Baz8GqwEUOotIkQQMrewq01JOv0+z/gz2rMy0d/n4ayT3FSNgbucaYq/2NJ6UC3e83n1KFWkSFqK
Llqa8qFss20Yg9D5sGj+kAEojzmuN5qoMYO9dcvjGNODnBZafw1tf9cOKLG7DKtdxD5Z20b1WXUo
nknka4G5NbG8ZskmE7bdlqcXYtUzukxTRvs8b+kDp9p5Fifn/8TpftbaseQV+me6j+AgkHaqS131
hCBWBIxJMgDHXkbCvbYMqH/uFdq5fktV4ges/uKx7MCbNkHnL7JxeRQAxVhFS8tC+Uizv8PZm89s
Gqwyt0RXh3UKiWzO1Q36gxMfgVpSXVXjhbQ5EUV30pHOLZ/8fKXtF2Mb2wiHI/WZrsAHPN83HTRO
2wNfzkxOaB0FzuPsp90Rd230WwgSwMNDojLZEhsSQX7QHzLqvGWR9IFcdYFVSVD2q5eJJGKVzzWW
OYTjkiKRW+izLoHBvkLsXUrdlbYzkhMDLWJk3dnl2lIiexfXur1pnShuzSSniHbAxxwAGG+fU337
urtkwUwfdas0aGrQbRkJoXtyMvCskSOIjMYGaYMIFyZ5qyMF8Ua6cb77GbHJzLp2Sia0Oj+3dMO6
fQxPdk+PmPtE/Sgw2LXHCndR2Hw+JvUey88CFL1gUzY+ys/eUtP0wthCCGxjCbLEgNFhBpSbRlB7
wMYWk+7rD4ixec2sT9Nq2u46thx4wmdhwTYcqOlLtn4D9CSkg6GHqJaRCrpLmM6e3JxRcQWRwO8r
rdn7chb6YZCrK0yHAKow20ne3vbLWllZDv4RhCkH4y4uyUQAxut/I30++lcUv7xUY3WluX423zvY
zJsMMD4camOMsuA2wfRTHlXBwE1z7jQoUfQ0S5hsJQP4fIQupiHi16qyzN6c3+s1Srieb9QG6Ypn
V30/H2ZgmBEFuSAdjPutg+M6wawK6p2ETV3d5wcwMwrlE22Wgn+8Qsf7FRgK6eLeURGxAcTBET3a
bm1kvSe50i4c2JRg4RHsXiVae7+HjEvMBWhuP21vokLI2ralvuQRMx5rcvWEY6N+PIsTkCzURBsW
jId/lME7ZySvp4CTy+Pt8o2vHJqpND8ulEcIxUh3totmwgbTWzb0iuYS8/Bfz3V8A5/E94UXuflm
3hLnQ5WLhMbp4I6vAoMPiVJWHVx1T1SFOPi9HIz9xiIALDn4Se5MBGohlYK7Jz1n2T4qUtzqodMC
H5Lt0cs7dcUPYWJgel/mNWD7M/f9jfcRnGXT5e41OsHvo6RGEIsR5l93otsOXx+sidUBWhw7cGoF
iYcSj3wFA+zObpGjzmg2i1qLeyDDti22iq3Du/l3Hng+8cniBSOfNqAK9ERfu2tPGpwEaR7DZW86
ZYImD5Kb99gjx0rub5f5VS8XCLfPnbfgJhIpxO6gmsqWYkXSCJ2XspJat/i5ITBLZRcvJZdUXyQ0
/C6tF+cWw+p/Q+N6bCzQaq/+DUON4dyBTsIBYuhOcHr1phTUCJ9K48beIyS4mRKA9MlP+g9sqHgb
Z0Y7ZUwc5iG9qkRF70ltkiviH89RjzfvLC8/YHXhlp1n7Cfqq+iq/AZSwscHVDphp4Zi+za5bCqd
QLllvzmaMLYgtQDBHBg3vsQwKKMFfSTEBL6pwbNCroV1TxE59Fh2ajReU32xybPEjc2f9qoefvD+
FaXmvmGJyzv9TJh6WvpRTd/fwXfTj4Wdns/2hLjEkXLGL43EpQXeNXa9EwWwHvOqjFVd5+080/yj
LM24ebVlfiP7TvNV9oyENEaoEqwdNcH8yBldfsDOAF9mOMqXXbcmOD3sZDf0a8QtC3BK/DEU3LKU
JFVcCoegf27Du+9dS9Jr4XCFJxt8GwR9tiupKXwqUVW8IscCyCyIUDmHI1eiBvPMeDcqeW2Q8Kjw
W+xFAk2RH/ERo/eImgF2ZGdycsbywrwGYKH47yfGIAyLn9/QKATUoly2qy8FlbwGSaW3W/wZTwv4
zhEAx4ozk4ggvqGK1NSppyW+s+afeztK+4b221hmt9VUgxNnu2Y9UnynpY3l+e0qlLqKFpmmkRpg
iBsyyrrhRYrkDtCFecYIvzCAOR5cUdgUjFdvA+RBlPN47Zs+7mRaE2FLXRI+ZJo8y3QRXIhDfu+K
xHtECfpuYKgQpz3GKY+glpnP5/ARtiTGabFytoS5+hMYjftu1XDLVudpF/LP58lO1wkWdilGZxvK
kZtnC6xYKa4rLPIAAwI/lJ1QQ3GHyJyOAgm303RxYQDaRbw3yuWgjGnFwXUYg6pP1PKGQMppo3N/
o+4/Qb3YvBpxYZdY0/HUt+1xYs36/hPp0Kz6/12Mh8HNRWUInaopSMVE21DEdq9kYYKQnN80rgsI
dvVzGkdkC78YPVvGGXBz1N48PC+lR3EhA0zBBNyPa7jihQFdOFKCLiJy34JrIjdqYxIDlWnexUK3
8umaYyy+TVvEquB8NLBuDiuAuLRiM2LaFr2pjfAVJsa298e0esQ07K8AKyW9sDsOllCme1tiDjm/
dWDL8keLd1WRtnBzPOGwD5O4fD8B4Ojg0zxGssOHkbIYC/78afqirPr2SL6C0yZ/EqFV7qziXt4o
64b0eOC11COUsrqflyqYMuKbojnGwDoYFex/9WpXM/vQjXP5bDPo0KxmahhimOOpZbHDOWTG88ll
D7fAdWf8
`protect end_protected
