`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7472)
`protect data_block
UkQzrzzOC+6nAVErMbqXXQ4LsmetlyZyo063++wXcvZOdNvGTDUoTURrLYEb9XjpwvMCrjujxCJm
40wQryGdsJd6vJcu/qxjLRa/cDIgMzUnmi3xfacxd28QBIcnI8Wfw2pswKAqvQmLla0cfyhgWvgw
u5LaEKPX6B0TkQH2OIxdFS2f9XJ7wzzfBN48xdJf3bJX59kfEgo+KxQRCRFmzp6SH3W8+1WS9xKG
PQm80PkUKSoEd6zKDvfWfFQQSUAW9ag9Pfr4bHo5oH1xmUl6RaGq5y2pSsXgaee6gDtq1gpEwPEI
prO6mK3GTJx2OgYxjDb8qZSJsFrWr14mDbtDnnDMbJ5tq8J+49I4cKfpskLadjdDPTe7cwDNA2Ls
DQKthKVd6kU7jQqk6yw5Zu5q/onTSv1oxFDLcl0t5pxy7sm59tOyTJkGapzfjMdRskyDW4AWHyLb
C6ljJHHBa815EAvJYpDwD++3Iso+z/Gk8p2LkPLXONWzh4HHU5QyVe1ImqjURyauarh5u7Psn/N2
wSonKMMItuQZbZlrD14vdiaPspnfHyuO7RbVdkgxuGA9LDQslWLXGKekK5Q7Dv20/BaHldXujIX1
h01PJGhH99z6MITuzLjxCnmwwRFC7I8Em6TwMSA7DgIjk1vftEiqhkZ0YKKneMVbjiymNWpyQeG5
kEKnk1hCv4bNCuAy0ygDFEhebivBlrY8ObhJdOkNtsCitnLhuQXQUbq7qc63bRrO58Rc/DbKVyIh
3VW+h9NLdoigWOBvrmUMrp6pj0ExiQSj1nP0jaDv7IJPq5LmQqszqJWU7hewb/bfKG2mXAtjRfop
j05ggCfLoXqapIsczSLTt5V35Im7Seu0Gv0hVg3aTIDxZP6MvaZs4dpuN46MxAj4ztGGRUHwRTuX
s+YwDOVzKEk4X68j83okeBmHvniVjAPuNZzpWq3xoxI1v33s5NkBObxm12MEIFeGBie7XO49AJ56
Rdr1VO+igwqpNfNKBmQSvYOqOSJD7aOla9pOwfFggpZwJCgJt2EI8EJrFKHqDhN1PFv45h1P4hmu
uwvSSoGxKUWCmpExbHTb63xoyslDQKUBdQNvshUvrH9OL8lKbGWVaScxFsM3DA+o7/TZNblONhHC
sGjEYjhcxomedL8c9j5VNc/QmwTMypZUcj+bFz3BBVc0YP6FUliBtjCTMXP9o9A6QYMnRUtX182L
Og9f2nLWTcWyA9gkpfDhMlImBO06JFmY0mJQ+tatNGzojaxJMSXhqwWHfo74yeFuEcIJUR+3kmKS
56AYsRWV9bFOGYqJpo18V7h36o64XEPNYp/ByIVMKb6UZ5vFHGTyuKeSvhr41Uc+rCMsG8Xx8Q7R
woswt/pac7ykkZJjQzQGUpcWU64ykv7JU9ndotKXnlfxiiF50i8jx6SaaRyhYtv4o2w31XdDC8W7
rO1681YIkVUJcsP9gH7qwBMWwBrgIsbczamUHL5bW8xfRJYrDCwxjEspLofeHYh3GTgQFh8gUNLa
7/eAk2RokJQcNM85BUPCbnOiCK2+WeZ538lyK0RT8ZBmAWtURTCVVvD6Q1cCdPkY7ikc6y2Na31Z
UhV6NNfIu0UbiISLIeW4nnGlEv9Xrx0ygpXsmhaJuZrH+4GHO+Mgt76FuQL0llikJ5bxzAk00xUc
Sn8TAW220KQyYlriEMe1yxJSsXJJzPQVqBW6lfEBJmlv2Jv/o2r0cnx1F04AgzaSndCSBdt7Wzn3
bEAhObvLp6Zg+/5X9o3n2geDc1KVL7VIKdVUSTLJIDytT3/Ys/mBNjTb+To6Ebh10rbvnU1Brj6E
xdAkazNX1cyoHwqw+f4tkSYbsfb9HRKRKrEVgCHi12LfFl9C+qRTXQbkdHb1oWSiSYzIX6Pzy6SN
JJUdFmvRYAoZfSl3sUYvqU3aFwTMn6W2e/5QrlgWJw0JuZPAgbcxLWwv8wQ1CS4exTwsp/Mz9D89
UZUxkspU+K6GiG5BCFWQe4+0FwPjBBaDRCETit8mkRYWHJSKhQUMUqTeIZBqw/eGfYm40l+BymHH
+6/ARLYK16aTnmHIeYijl2na3eUL9A06HfctcNFs++aMAMQvWCoybZ0h4Gxqy5zinosMAcim1tWt
r8o0ASXUAQG5NaCIpeaUnnXfCtBdZ2+1/qXQRJp3ttyne+AkWscgtvK/0K5ROtvQb/wOI22YswKu
Ut0zMriBYH2Vqrr/Qau/aMvDyM8o/unDcccrxAwGXcjQ99PeUXXPEpflAIkVQsPTdv9mJSkfX96R
cn+gcWQkdQph6wfyDvLDn5PChxS+dXd5Z1Xn6u277z00NB31Wb4jem/xXLRVHRUOWIy+yK3nrPOK
zxaWtuCT5mw48ry+A1VBvl8riFbVV3VeoTgCBKK8XAXoAHWXq1888y2PgYO5lQ3zUwO29QaxHJHz
kg8+w+u0gIoWsTHQ+7IHaQY1wT7EanXe7C1M0SGibQkwRw+Fwh5E1GLvbSVxe4XSABu41tJB8CTu
/f/c8V12BEkC/6CvmLRFeGWnOrBTYL2XjBrDrc+EdnT5FkoOAmNReIrQxoO3sNW+rGuWFXj2Dr/t
qUEail8chhYyim8cYVi8p+zvx1FlNL5VlKneexWuaD+/AM6HqcwZ6G2mkBffrO0w0pqqsajocoBD
MoXcxvOFdjbq65/eyeY4z4Kibvg/5GYfQ7xvKlsWJgOYT+DhdUilR6nord9WGjoKGJR/eZMf9gFY
GmONteZbSXS3G727fhVtlIGe5Wz/JLThJvZQdWDfNLkctC1msmPyw5iyDvOgSUHJtfrKVdowpd1h
LLCseamSUPICbTd1OTsQR/0JVuSS/ZuUDVMHn0/JCNYATtQlhNV/YFR/odo0LbXaHvXYf7iVVhNh
iZmTHmACYZ0b+CgXCI8VwurbcKKH4o3SvsLipTZ9tFKnRpqdQrvdG22p9UMv2PVBU5Ajv+/N9YKp
5nNG2mLFxS5MHwrA25NXZTLOXuTixjg92o6BqUkD+iVHTB8AAFiL5s68iAlDm01W1fm524lJ6orq
RpuBom9pEb3zddlZfsS+ksB/5FgfIfLsO5kewT/eF74BVK2OL10F9/6IszxT5IERacXMRU9iGIdZ
hNrjaHFXvg1/+baBZq0BYqD1dPL9P51XKdsSl4QK+vF/KUxeiNTUHNv/rzEjceL9cw7BZvw1SA8G
upyU52aSpI8r/+drv/CNJtX0yNxKLcaPxrt+RwuObVhlOxgzW8h9r5AtIw2pMqzNkBXkGudLlnKH
qC21Cn2bIN8tffA0gRvVBkvHUpK6xmKEgOZA3ZFBvZdxyY1Yg4rQy26deGj+TvzeQdfW/p5oL6sN
ZJ/LW454aEsx5dtYzdkAmTVR8OrLNx/Qjsaykvghl1hRZiGqp6ISqtUR5JBVC9Pqa5DOez6oP48T
sEOzAYt25HoIH25/z3+CCj+DqHy0JxsmzGMowL1wfvESZEiG0lEIsBMubGL3vEiiqxYlz7Mj1BIO
W88KdR2xZFP6kT/7S1c/z5IGDmuoNe2ccLo9Qjj8s4S91rNUtgCJvUksx8cXjGchClpkz0xTSSXG
Xb+dlPia5Lei6Lg3fRHLsMHTUKFkL7vH37vmNUo8xzJOPDbzzLXfFyS1//FHYHNkKr335fneFx/p
TD/LH1+WYgTH5usPV67JhP6K9A4lsC0c2w3GQIcuuuT45vQBO2BqilUFskszsfcpppKsL8FYoDdU
7lMJxTQA7YrThmEI1GiKC1roeZC7ERDSHckqXiP0AtoBtv3hO5KZ/0LalfQRXgkHjlE1v6IZpv7S
FLYgmM9rDK+pQo7pXVSjdhy88Mny5+8Ifu3++FX7YGzb9ySlulTBjOd92E48E+5CneSz8yxO7j8P
EQK7UPiOD63qQVbZUuvesmrQKv/eMIei+IWeKArZ1Zq0DX2x3uFk5sr4CnNMFej4f6N9qLFpZFcd
u3zOXZlI44vV86G0BV8nxskDYfvLxRQszav5zbl3dFMfK4mc3CNsDWZgypn3A/QCl7KO5cAHLsUl
i6dRkHJueEcFrlJPkpjL9iA0nkjxxLlwaTJbGNWNDHxHNk/2ePhF0MCzTMGqmfShFZYAVEiT0DjR
ezGVNhUbT0LL9ECG/TC6wlQtnXy9kCvm1yHTlxBjcQe4M2JDMDTyHvyoW5dc/QrED5nPLJXToZHB
3oWKD+OYxLWwJf2fNdp94W5VVkmuUkg8xxYmzldBq+B5sbZ1jUyppUx78iGZtp285QZjXpyxeR//
DVc5KxyINyd5BtS5zrcVROK/3CndkVyqYVK0MuaSi9tcU4XO6PEliAXxu5+Dx5/8k+tOhN0SZ1dW
RmlNK0r+BOrsdpWGQ17hQdfB7QDv7H9kB1VLrrl/F++YbJ17FUH2hXSblVRQ63ltEKQ7onFnwrqW
Sx2vwaOlxhcyPwKnGRIWjpM59/0Evj3rN+lFluyOjWZlk2CNVjTvYGd5+uGop59lKKCEPTBOUC1C
PdOTFSddBCubs9HlV5WOwhQ9+goL9rfk7VFxMXmjNINGCz2tq+ug/VJGz3QJPjFE7VyzhxiYNtd2
ymNBGThdlifTw1W0eRgGEvLfMaJ8cRdDcwZBYDQi0fRS2k67P7of8TwqhAKVi5ejFMULtOXzeEvw
QrGlfZXJNGtpyhUaG5y5cDBJfBGZjCv3u5yFwshtLoUT3Dn9ABH4ZVtFD/hdqudzGasvS8Tv5Auh
V+kCcz0Gbz3n/L2cJYfNuuxlPDMtEZmsyl+5vnT+TRQJxIjfz0GR5z3nsTbJHUaw0zvUOQlq/HCz
vZvkI+pifJZP1TbGEkc9O7F0UPZBoYEPQ0TQlc6JEikwWp15lBtFJMmYUaSEcGvonEqopqBg5sh0
E1S/SiXs6Jhh+66QEHrE4jQ8ELPJry7D5C2BjVx47matS5wKG+VINeqr096FwyvsAOJOIs+a19be
u1phT/7ijZvO+ALwOBML0XEYftR7s1/UcIldHz70xWR+GOblt6btRagiKS0XUhc6AI8Q65zkC+vF
dl2B4NarGbYsAVTz+RLQmsOlZ5ojv5e7HeT12PM5C7rlItkcKEUy7woz9S7qHJsfrx0/+TIRTvPu
0NFHCvWWR2vVPnQI4XjKJuGS7n2084wZZLZNIIPNHUFfmTk3AZx9Kl6wKnGimxMBpSOTwQUPLTxn
X80gLuciSSifyIj040EsH/EaXgHfhNk5VxvftqKdgjT6O/dN5O0A7CH7ez8ZfsCjx9Oc3FkrfOgI
GVejwEudtfSNduA8QvT1v2934IUYf+55x1rtlo373hDV3rrPWWy9LAtEyZPrdBxBFLtrX00AAXnk
RhpaVpc7GFOd4YTQfCnMMb7P7koJKrAJBQfWQl7wb/rSh7i9jxyidZOiTTSWEWd3JOF+PXXVRLgV
qiSN6xScXNFutlBePneSRw9VWZytSTkGzskjwbhh2ztLePhXkPOH8E2A9X8yR/+iqwSS8CLplxos
CfIivD0+jtU7HQiCdTcgnjFpqBLP2D/0Lsf3pC7wT1zI6yZOPbNZRvF1LSXuYUN9sQ2BH2GPaBg0
gnUTFUjmEow/y2KyUUPO1Jm70ZMz1yj0qxiif3SO0jaFQKi08ms/Qc7BW4DXRbxnYghwBv/nZHBf
sL7Hsv5ApEc+heNXKr+61qkJompdaNnuC1AX+sarQAffzupXBOTTaeWiHHRGoA0otKkkvosPMRvf
AIU1q+u850ONDTBMYFgcTOWzzlFJt9ocJkCfXGlEbGdXd+IkZjULeyfQJkGM6k51+N+bMDA3ro3Z
/cxMhFhQuEERcmn3apESHqjreXoY7Z8e2jg7k8/ksKjJsU/D0p/aSq95GP7vQBla8TljWaXpRuE3
ViO9o0BfcWcOlWPjOeRuplYPaXxpZRZY6xIxByz+LTA9NycSF2KPJqqre/1T2dQBUyZyWOz3pDyj
aiVjgWBRIJYGfC/WaJwOSy3Azps59HwzmM8jmz2hYBmzKeMo9j7kamuskj8fxvgKTNxDtWcoboNA
FdBKuOsZh7QmvnsroGf/pSdQKP4KBLhB08icW4P2TvACpJGD/pPS2iw5y5vaxSANOXduHcQEwlUT
DuWjfonLJhmkFhHlAdYdfZBr2knV9pdTRYwoGQQRQ0QdBmi7lItOuSkc+9xJ8e5IEx/2nwaVtJt4
AhjsIfA8fbLsnc4MscC77oUCIs09Hik6kPrVNtN9STYgTFzEaUD8TRBIrzjWEZlFikndD9Qj7qir
PMXROpNiYkhpzPEd+U0kR8k7msKTO8rXIEMmADzaQeo1+wCfUWr6+pGxDNMfPz7ifPzqPRbaCwpU
iMJ19jjYRodjeWcJD+RwDtPn5mg9fNHk9LF13sJNYeKNnA7cEWvgdfKYc4wUAZ+A3711yoHlfami
XSPY2MXPRe8g6HF1ShzdEQj6xn/ddYpl3yCpB6o4ApTTXs1L27+sq2pR+8jzsrLyQP8MefBWyqnS
VrMmjPVVetVBHIjynPOwETzyDYyWmZO5Tyhy4KDulG9vnrjpoY3pY12Q9hFro9aEKcRhTDPQtU4f
afj8Etuqqg5PQrSBnWQX/XoBWvHDOQqwDcT1LGgqCJX+9XlrCP6hnV01q0H+a0rt8aiWUx9P0yAV
7TUMxd+yFmU3cSxUBB4EtiVL1VSCDrPAgRc2NXjcDBiox0D215XYu0jC8o93Rf+LgVMKc9OycdsJ
a/LAMI+LP9zrBS5XzOGjsdh29gr/kFrZZcLihJSL8yFmrCwg9ml+S7FeRCiwh5irdqkr/jtpWnWY
PkWciL43jgNUM32w8E8mv5Xl3zhRjOL9OZ8Kd+74laIvkZ1hLztNoCxgMWYOkie+L8uFAogCpzff
H/Lg1aMoXWi70BBLzBInf5PZ97YbawxmHvI8WToc0WOTsV73KZTelIMWPQn6/ef04voTOvtHsRgh
CGASUzzpj86wn5YDBs9Lp8mzKv0CGMz06y+b5tMO+W/I2wj+WZy4OTJmvM+yQxiob1dOZLVFfsZS
CJNhWZONYTmGYTDUmMZMbFFbu8W5fVSbXqbdiq4F5jeEoWxJb0cZNE2uDJABDPE1D+ygX/utA2lr
9OX8TNvWuCmMY+TSjiQQfQRismpZ6e0pz8tkVBex8KNWVeSP3TMVYeOa+i8Diq49iGSkS3jNO+qf
8TRdlquxDSdg5tpBcJzxEuhvXWmyJEk4Bj8CcygoVPESFH+56KGEGWYH5P9rWCIMAu5jvBK/Eid+
nuA4ukFMLZq+JAKdqLmcgQ92bpyrg9rW+95ibiQcRIspDS7/M4KywSrIhzLtetQ5rFdvqbudduj2
qeXGwWQIQ8VCJOdZa+S0VY6so0K7TyU+9UJKT78sM031pzroGy9SacwggHMery5R96T9bzMzFdvK
XObhUJgtMSdEdxFJoCcxbw2bAtZqc5Ac/+DUNs2851bxypSTGz6CJwY0O74rch8oOrJkgRg0nu71
TrbCndflyEySaY4f1Y3GUqFqyo0qvEknNZ4GorqsaJHaqYP7zv8STx9Gg38gvxQwRhdqadCvexjm
rVCW6pUuTQhO1ecF2bcW3XC6MjfRLEq+aa6/jopO1JGaS52ANmuGxr3eRQSqEg2pe+F6zrx+bpP+
8/vcxa87C63KtKwv7hKOon6qiT/Ec7znVG99vjrBGNCkHN1+o4twj904IIZp5s3USoyUz87M+J05
ObNKO4tA4yNZ/AHD8HrONw92qiNP7q1s3Vwbe92OzgxQd/zRYGQpaHw/LCYLJmQl5JBZVcPadKQD
Ln2pwOFhv7VIlZbhdObPG8crFa7lpkYKdkrD9byhHjxIq5KRQfWAZsPYVSb9w3mP3bXu++RPy712
GuFN1C8rbFNV9LhChpqvEkYxIHh7B4814uI+/rS/ZmRmLJx156l58vvXccb1UVxiXcLRRaHa9kOx
7EGdfb7328VDsrCQeGdNoMRNrCvDiye/Z9pkMbFaAC55V4of/MkySe4cS+/bQz4J7bBb1pQnu+1R
CqPDL4eOm5uVg74YUQwr+q0XWPirT04Kd6cEf+uvixetv64fT+2QXLJlPjNmbMeESRN9N4OWBAyD
MVLwqQZMLpWH+r67n32+pTux1XyrRTlpO5h3HWFG9s6/AAOAiZXjdGEX3zP3e0mSzAPo8zN5Bd+y
WPHU0CKWESuTnld5f4O0i8++I7DzVZWrmDDgMQENUbKkRiOzA64Fazqr4IfV7P1Sx5mSqSgwGgQG
wk8RVMot4zIIuIZdNtsUkp/+yP4tmGkhvM8Z/lqyQJ0l/djP7JLMoIzylw70FuprOJSc5/O03DwH
Bs2RH5PH0Mbp9jJkpHbddw/hVnol5XvQNlxyRZBxYYwd4vR/8WcHcttMhKkyP3KU3KwcFrMy/UQy
+DcT4KppL6pX+dZMr+UFm4Elk4521kZPQ8S7blap+SwjIYrUV6Jt4yHCYVf12ABOcHdYYv6ZzVVX
wdaZabFYNPgXtb5Pt08FTUCCDJV/uNcocr/197IObyoGc0aak2ablVH42lDYGpCIDS5YK0Xopumw
Hs2fHRyhBA5hq8Ce+JsnuyA8jfM7Uz6QHxZfuKwo1OKwNNRbo/MwF3OgX4oWwNzqDZtsPWnj4Aj3
iOUjP5tiTdm1vXJWSqlCGTYg+a5f8Cz9A99fd7RrhpmEIO0FxET0xDmtwzATU2NP0ahOQMPwk2RO
iod8yjXEIwUSo6ZmlIWgdmGsRp7fSOO4xLGdK4ZmPqIP5JLSKe/rLfhGcVERBcRpwNn1O1P2FKz1
ApdfEiQwPGBwPkoWSbaZh4oVfy9+nG89dcMrYIRz3eyU3ViHwX1Jyk9yl39PilqHoQY/G4X0TuQx
2rApWOXqZqGE64jBNWj6K014ryMHD6qjx08SFa6ENJanSz3N4wQuRBF/AljkmJG8OvJecLWv03lr
BwOM8Xgk8AmQG7IHTMiIWuTNgKsR5D0CuxJFWVpRR+5McD6Hr3KWLwIn9DdVr+ZxjXZKrDU8gW7e
+vY65ph5NkDZ871p475NlZR7b5vGnR1gvI39t9hBf4AKBIxptlI0U03We+dNNerDU8ZT4EUKawVa
M3px+oKx1EokT2XCWQEbGkC7PF28aAPIS72eejRBQv7pmTmJ4HznfKvhK65RxP/ex+/58n36xE/5
xYNdiFfaG26eAaaEsdVFXoF1JYUUgug4Od83i8Nabw+7ACbCsNSt1sHLt2VwakV4eqCQKs/oPCa2
a7GnURTIvzEJw+1ocFgIqc+zYo2FOyLCqD6ttwpZnUZcST29ZaRcZqdfLwmb2gqZLPjETOc00JLv
aNv8jM6wH9Lgxbn4dydtwdoRgUOBnprX7pH4Qs+Rx3nB6dlIEGYs+UGDlD+7ep2xc9LMvqowbRZz
SDpg67ZBpiuu+nSZETdCZsB7N9eS+CEmY6dMG1W6RUBt1d8/YPzpE3PlOzN0ZBQwWwSfBQfXi3xm
WNjAgRU2JEEH2CX6a3Wib9+HQiwXpjbiC+8Y+vPpd8EHQCLu8YsEsvXq7kyL/O2fnaSTZTufGsXK
k1d9mHZCot9ZyWXpqJIifnhOAF4yTBuhmKfl7AY4cbEcWaoSJkF8dlVS7r7yQnd7de2ghPUdbS7+
cXfc9eqyxd2VlBQ2HtJSukVi4r1kDfXnaqtOM0AogEcXMf+x8x5HAvnZnTf52wobQlHMA95Dhnak
ywSwbxRndwNQGPZTt2rG4ovdyPYuk3fgEM/vJEXZ34oBxKHahkGxgJHkeOIivRUt/G66pbJZQQKP
E2IbXYylM6yp3LRvXrY2vah3pqRpjru0xaBkAof6dEzhglm0MFpZWdprrYHkA+FZXubEzDm7Cn8m
86cVHoDyEWdAZVVpGLDMFvizFFCtNuKRagNcj3/im5gLIDjlh6fTEg6cFI9+T95pQP0iimqmL3L7
v/GoHv+TSaWYkPJ797pCldc7jGM5s2GNRwPisi0QtO2dqZdIPOtt/CD8P79OQf9wgYts1ftuqqzX
QCLiQpk=
`protect end_protected
