`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17312)
`protect data_block
0USWSUGxovGsyBJteYpEoZoMYTkNXR/GTn+lRlGRKekANJTwz2MgNnst9CoiV2BBl0enoK5kqInF
eGzV+syfqqc5CTKNx97KhnmBlKgYT0dhGgloj9GluUw+zfb+k/umttwFcC2gO4QkGSrbfb2b/2Rx
5nc7gCOB0voxEBUpdlfEbPllQDZl5UviBpR231IQuK/eNRuNu0tza1gdIZH2edQplEyTzJzQg9KA
kYxSGwyz+64SuFRuSCcZC4jKPyN+muuHN8Wxvnf7TDLZyzHWwKmPpjp8a6tucFAOrFVZ3YW/xlei
gyFekjMYEUkykx96pDMAOdBnR8Lm9dljZre7rstoPnUY0wn+pbYgTAVQNiVka/nnPCHcN2lFMQEd
2rleNp/MKLyLpbbNFPcxKTMyaqkbUFXAkHggsUlKQoqM0BgQKqcp1fb8HppivFsMwEmJVZ3VDwtI
7nA2id8LhWdituklHubJeh8J+pGTMMCNDyhubaoWS8abMkkfJtXCgSt0jFv+Hu0yKwN5KjqKs0KD
7W1cRaq3j1pb/1ljxNhRedH5kpX6i8MG047QhgssIzoyC/kb3ZDwrxL6YACEhILyRKRjgAApAEFa
1uuYduqYUbCW2uQozDU+a2vJOk3EIKUFGi7We4/lOYeQKno8+JOCQ0kuBGrqMpTXEJmCcYMtHO+2
eFZNvt6DgazaNLkSRzrK5brLlK9Xftvay/JFAglC1AG93H5Tr5e6d12cvdNgXmxwZyheDL+G4jzg
AQ0IMPJsNx9eaQKKH/dq3+gjLUCvisZUAg7cSAOZN0CfCyGC2DaSfjuT2GAiLyRHinOoCJEMS1SW
bUSWch/6uyx0PjXJ87WjBnzQwZpvJnbIATvqMDc169baucdM9B8oxD2FapPFKQ3iFMs4Gq0c5oqF
l0MTmFvkOhPLGdZg1em01COt6kyeU6cMgJkjiXZQD/EXnDUvBwWlWnn5aO7XmHKN5+NXhL+wwHhI
pSeskT7pHRGsx7HBDUbpw/rtsqSGaaaIONGU+dm9VSYmO3eNaL5/aQNSmH9iUVUNUZP7+hzA7OJk
RCOp3DYAifkBozh4KPuuqZBnOcsJbwJ7W0of5Ts0QdmD/5B1N0sqyVvXVX4ypVBwaq5IVmo+VNRV
GqyjtrEFiEL07Fo8sKfeS0PRpFWByHSj47OEJ/6nOPfRQMVn1Ck+taPqde06F1qXR+3dNGovNhku
hPvxjZxps8GILPoDIwGbig4Y5q780Ge7r6H9qx52n/WTQ7cM806yIBcX4909yiZL9wmlGsu4yYnN
ikONXCkQ31k1POqk3vtsmLAjR5cyAX5FgV+0rzfB7xB1LO9iNDIT0ubti34iWWm7iltkM3IKA1/4
LqED9OIGi+qQHIcSRsvsRkSe2kSqtEXFBtl4anEg1d9qkxOhBaUrQzFz60FFkcFYZD0j1ERsozge
W5mbJlQoMneNjdhO3HWfLP/kpKFslF8ZJ4R1zYavGlKQBm3JUBnNcTvzDGgwJg6tuzuJfTVrLRoZ
RoAQvRhylOQRnn9XGp8kyiMnN/RhwWHClo+RbS0F/xpBfx60Sg2/C2WzmePnYpA1nDV8mpEx+wKF
s7EyiPI0GHNTrO/mIhH3iGigC8g2ay6FEsDWft0PCjcVUsGv1hrXoIQ35IaRa3O1OllnO8eR1C2a
3y96bNGL7IgcRNQPODmcbARzbxktr+4ks2j87M7U6A7Ha8Tfd7IrRxMkjJEZAucnplQ7V1LOIpJH
pW+Jq8TOSy/UFKvsxZx/OnnvWRnFYAxh8lqhN9hAkIsJcq8QHZ/YhHUiEpcDwnkoWac9zEcJBOY1
jOS4Kmh3Cynxnpgpk0DNoLJtq0iL4KvZgH9s3h6E79cZCMjeQDe07MI9gw1njSeqDxngmCOWzkd0
l8uQx057v6H/8VKIPrMX1iRMOSg1Bb+D4GH/pdRyiNVNOzFB7nABFSKds0oR3YAyZmMUp6nbf9Kv
1QyUzn6qPYysM9GDWPMoaL0m1AhoJVubo74/x3nAr6MwR/euc+ZRysFjvlAHItyJnSGGM/R3X9dR
mCF64ss9uRZItjiPMq8KGJi01G+gb53+k7AgQVAYkWvOs7aGBbm6/4EFfWAmUe9z0YVSwNRPjkgu
DZQ6nQWjXVsYpihpZbLw96RAeazWHHVmLdfOGe7ptnUjFZyo0U+H9iYplwHhGoXeE4nuVmLL0aTs
K8cJenDBxV8qEGTbZXfv9FZe5e2rK4HJUIHSnDGEDGltN0Ap7ohgQoo135ANVM1ZUX/2WItFdup5
Mkupq4HaKHSa6eZnHXJiz9hCafoitwv6QMbebtdDKRGiW2KKcAvlk6R7mbgF3dTyNcN+SZvR9TG0
WtMVRe9F/InKqt/wR8q67hNiJtv6VMtazBluXmGjWas693RqcRZJPo2NdW6bMR1OLkbtdMDhX6/c
YFbOkFEjSAWz1VaSEMZ1ortsB83u7IkcaGAXKGFBQ+o30kxKW5SxPmNP30xL6Hh06jo6QeSjxeej
d9ZAZeP5hmh6ux+7AMY0CzyE4V2x+SOW0iNu4RnVG/JRFrPcol0YEO1vJ4Cz3aM+1XX5TZd/dMj7
o3VBspR2La/jd9s83SofmIxVD4bzykyW4hEwreyOab3Hygbi4y4ES/tLeleleNKJQiubwvs0/9sE
KuOKCAYCsioIp1WS1qgMEcAdcAwVKWqFua00y+Ioa8tkbO+6yJ0m00Y6yvJ6cUBlyC9XO4QN8w/8
rWCFwmJttQrDb/CChHkCBF0PiaBIv2VT7+cf4s0udySo6bAT0oxBQvGyDlJzVUv/0q5jn2rRRi4K
/LynZp0BBj8cmbAbhT0G2+3nTK8BpQNLnTVaBT3i5ZYSishtVVbhHwak3w9TUWL5pOb1ZS0TUczg
Bfczie1xwEZWO3tgQu+VTRKX/NyTxHJJpO8hT3aVxDU/rZnHSd6XmvR+MH/ys3gJaJppoNwVLuS/
DXqDE6o1FRvKHo7MeoMkLNNOysi9W+qTCcUtDLbSqVxp8mluXBQTwQRL6kjOh+E+wtBGUwG7CNHH
5px2m6HpOg61XudiCjLup2M6M6Ct1zui9RNcW6A5HbqfrzevoFrDCL+i9WOgPFKRGNbKn7+t+7xg
+HpImASP3XR+gVsXD8VHQj1ywJ/lOdqFLPhOuVyBBd2XADadUjXAqNrvJUBl0x0vNpMlR1tgt4e6
pw3DgBxP4Bx07b2af3wuJe1+BeHT0q3OlKcoayylsrGVR5Pj9er+XZ41p16He3ax3ri+077MjMcv
nnGVO+SiWdDEIvjHxR8oGd2FzGjcZYo997igwGOqEfOCAzIm4ufh6RtBEI2mm8aqB0TXm/0Lpk41
TYRp8iOGf4JQ3MdxpKkXoFqsP43xf0Hba0HepNoINXD4LdQV6BoWFexm9D/uHqfhGiHEP4yc/XZP
SLaUn2uc/pBla/ryxGbA/yibTLG7KZsbZZcWi3v+k0tqt3Tmn43eyIlfhJz2Vx9GCHAYD73HfN3y
pmpbvg1/z8vkywpM1A59LW1TGaXp5UvoYxPmbiRh+KKH6EpBfyBzWSfTMYGbMxGsMXNj/3pI6/HI
PI1OK+S0tPdVdcXc9hVL4INJqws+siuoocqeS+dOrtcn4ADFR7xg4OBX4BuZHdU2QbIOctQAdpuM
eXU/4mHn0M9UHUF85grI2lWNq5eyZ7Mfx+HU1We5t1J1x9awz86X5MOlGvk103hVk2irWJZq0wu8
NPl2MAse5urEZbhgJyDbYUul2DJ3zOC/XI64yf43xbQcAJWlUFaAFAw1Sw0rxcj43JfEKu88+dF5
U6VDZEaNj8rzKnhg4cOc5gZO/ig8OTk9fKBSC4Y7UfAjB1mpKjB22c6B0TH8P8lMuFT4UNen+xYP
RBnUpbrtucBPBeg7g3QtK+Qvzmxu0z1Qi5nIB+YDAaM9/Uxux87hjBOEC5OxWFD13iR83YZdIm7w
288ULBfYVluAezlLYa1h8LCztaX9svaZeGLoRFO0kbyhWPuzN6FhdILxrEyz3KNUb2MoUZNpkypI
7iRYsgn9aw9b+dEDySM8CJoxnpDk1EUL0Ge2/i42JpeezY7yVHzpPCAGvD7KRSLVrYpUXtMBrrKx
A952NPukbDU8WjkIbbQVdX7M4DGZ8yi+ECb5rRkNLbTmncY9GgTDB1JAKOUxDNEIFyapbvqUilC5
rasTkFNesYnLdd85FzK6++Ly23KpaOW2KqKtKo84yimKIRUWCT4Cvx/RFFCkakIS7S73bU9XaSKu
xHFaDKNuA8zihzc+zfn7F4s5ghYUtZGgEZTQZQ1y5+S+4oB6nSDpBnH73zAI24XfhllBVIAsQugb
L5z25OLiaK9Uc986BarTUQpKk7IDVwBtqij/Iqy6cJyF/U0DjSKJX3O+u4+hDQhPABgoKdhdxmaH
Dd25mh5QpkWRoZjgx2qsYUBA2ojHmejp90VQjtV/ZRQngqgS0DoiIsKAI4O1sS6Aj0n5WLANx+Mp
5iwJQWrD0kpAlnE6ZSet1err2XZaI8PxXRv0rgculzsQOxXxNO04+ciMhJc3Ke2YR/vlEFlg2e5s
vTmSZLbbMoQNhkWRG9euX13P2r4/0BagoP/J6EC1LpL9Vx5kAwMDmQM18az6lwtQD6T2h/xhmTNM
4RkQ7DksTC3ODK28XU2n0JpyWYfVbj5cwzAK/iy+ZtsaqCB5R6/XWqlhpBCI5v5vufklBDyhbXvJ
DMjHVMcNfH6EywgzFynAugnQIe8qI2gD2GCdwhqnD/JmG0Kvt+2p8FVSqt2AqkR9889QC4UJRxj3
c7qQUBhw6TQGldVTB8s8yNmqEYfNh+r1ZABmdJXMnvq1GSaR5LhRxRbX9Ma/J1NqOzeFxwZEz72m
pW8m/fxSgWBXqtcL2DtK9+g0LS1vIwSg7JhSgikJ+rIDGGPzrH1e+KYEmANbGGECxL+LIWmLqhCy
YB58K3OsRZacWQYLstt8i2yMz3uZmIMndQw+34ayYVV6EmwUzrhlWLao7PWGkjTACK8LLwIJpARz
8U+jKOhFpEKAr8CWiJllpv/yBnUEK7KCCCAfMtpeYdhKXCSBUyUi2zkBHkPOzauu6rI2pYLACvJQ
g7YEtwU4XoOa2B5CWtJLnggHDFtMxuQJtzso/2Ab6XEyKx1aDNzG05czFeGir0cBqP3UXtDkDWaz
N+bFjoOhGH1J929T4pGZc54zfWpEpAzaI2jf2AEkLfwM5aZuj1AGo6zQsLH5m1y0RFbntWFEyzOV
8fBbSmu+lYV14QmHp2qoI4iaoZZMGPaRHKrq8C5cTtMxZSzD+SWtWlE8+rhfJHtJPOSk5C74t89/
US55DA7FkLsUgkeNU6cIdghor1iMzA0Vugym/raOvjFVf0x4pZiANzxyC1MEMlHlJ0FrmW+TZsUn
Pf4AMP5fv3+fqZJyE06iK3CWXjP1ScWtB96i0kSGNp66Zy8sdaJc9JXxi3IahhvcikWtxKyviRJd
rZ2wGgffdpgN9Fbs+DOZiBH5kqz9j5j5PuSYf1tYueA3L+N2+d5QgD+kh2gtFzksL1lkym7g8iOc
iXp42HVATm8jJTWr33NX6QHP1M7LumQqampAn2Yyf2xOWe9uy6YV/8JSAaqg5kerZABAjDaIjEpF
EAf2CPbcqCcSQDyr4SSWfL/ol5vR/THUWNeRavkYqpfdd10vbeIIsRwGLQARy3TeWZMOkmOG5gyo
XiaGc7vrsFjUX1febrLFSNlRrRlIo0LBXdUUAHaWycYLNsK3X0CkNJVSqaLGB4BxxTZNXK/uZwsn
PLzE8P4nHzgtDdKrOJJ9RcmdjrVMwSfwZDhZlB08FjO7tJ53g4KtjnI0bRTXaO+x7x1JsC4XYHzP
CLHSkoVkxFQMGshpxRPqG2qwzIx1k685xwCajXvhq6xAXVPDGYgfq7jiE7ynw6VEvES49suucSfN
8U/438u2sEssvGjjeSe3OSqNgyPeZ7EQuLCQ2MQYtjj8j7uhOZ5IUbHBgMaOvucX4AbcYQ34R1Pm
aL8hbEQWM+Q5BfZxE2TMY4SbKGuiLDwgv219ahDIOLwpiRu/3e8fOUvn6B4phkXLpadwZQj2WPYe
ukqzyBQZpNIEknnXF5wzbnslxhzA1h+5mNqvObhxaMDKmap8uIJfCKEezsrEZd3Mlq6ovPlDOzXV
dSqhDr8WYN/8AtSby9I2tCEhUMQ8DdU7CmO4OZrpbJ8GJSZomu5zZmusRy11tA7GAj/cYMijpmWh
t9KUvm2J6Q8ggfjQvUqYSKwPBvOxzavQn6/2o5Gm6CKrZazaWM4QK3ax5opmCi+lL77uQ9TzxOfo
wb7H+zDwQY5ah8cejpWrwsHTyzhajVS1eEZ0L81K8EkOPWBGnC/kO7makLjROuOr4keriC8n/VZL
Oilj+TIkv1kMGID4raTLjAHXeDOqLxoPnd0hDOo+EkTtETNxxFc8jjhlrdIqvPBX15kj1n3sYTri
qZAvlWsdm9VALku5z/V9ZUhKqTg9WJrkPLasE1+PZ3yp5DR7ODeyKwYQi2M+j7q5bfXSwzoPjKGS
yPkLdu9rWPzD0OX1GxfN5KrVeqclmvN8aT2Co8DDTIhCArtKxeAjRkuvn0Gldai6yBsHcQs33JI4
Rx3ojBcMWwnVmKKjBfUAqlSe7iIYe2BAX2xccrG5wmEA9i8X3fxmEeMtp3JMgHOpQD3IX0xEdLez
pYv3gj0BUNeJ75O/XPXogm/SlDG47nlDPaQjZTeZMWZm26un7gV4tdeDHM0U4VMjUvXqCoVSz7QM
GkHGh41t1lRjubUNV3coosqVOgVpj+EY1zj4QzguLta+5kjqUEPP7cLnkc2QHJsIn+PIrpxdislp
y/c147NJG1HCS2UNwt2lHj3JSG/VVy958Az16+sZEkmzTkwp2iraNm4+3QMlcs2LpAyydXRwg2fj
6puPCF77XtqGMhBYlMi/yyYuqqA9AHKttr6y2U1BjNWCOt0rW2QiQqt55VimCMcJlXYNbjC1rcvd
X129f9YPhPi0Gun85GgLtyix5iCU7GA5m4v0CwHIAn/teiZxHMXsDB8NUs4pKK2CR1Zo2etE6f/b
9DgZ5nG3O9Ji9iin6vn/xbi/Yp5J97TIhGMjRvYrMvbo1gASGeKPnvhH7Fw1Vtjc8jDAX9aFx/2n
Nzi4d+qdy8GegwGNiLpRwMwhmdJBJ3mIgZ22R7k31ODsM+LF4+XLV2Y7Uv3Dw/olTw+UdMMAXrEp
3Icxrws9XLyphMulGQ2cfd5ksKDLoKlbYR0gB2KFLDUhCldbv0h6v5Ey4qKgskQC5/TuSCbQ9ABD
5/NcUoc0tJjqaruueuZgLRqyA2L9ELa3AFyfnvzXR1Laox8Q2ppHlBNXU+pDVkDx7SbyKg5usBs1
mhY1Bv+WOv/G59o7TQI2EjudM2s+NuW43Lra4pQc9KnG2mlZAxmrf2yoJ3jWgHUp5x3CDjMbz7NT
Vg4JRTgpa/7ujAoszaycHdQht0B0G0/hAmLGRoSNo2b19tBPmZtAKRXl5cSAXS6DrxRQps/natLs
ASmGlkkNT8pjPS5lKswDVLeXHtAlonVcNSV+xnYn/xkTm784Rw1ldfJ47+ViBj3kFFTWbnR55aQm
5ZO5HGX2TLIC/nvI0XewbzcMH6K+SA+gzCc6L4hcuxWnxw1LSoLQ9xttjqaMchEX6PrbV0H7ZHNk
MRyR8VC3u2m9tfuTND+JMbGVVDjJEwE8FixJK8+6NzkQHS2l54fKbdcrsAu6TFXN0rh3Z2Azjglo
fjzl9AvxqDqyS62mqJRLLOOG3xrRXC0a423unBd06iHHtd31m034kKQJW37tnZAsT97xmnZ8KSB9
4JtENGJOFcRLS5SoZFPPoPyngT6kNzEMdrKyf7bYSSIW5PXFaG6uytiPz7lGRaUKofb5grZl+cOF
Xb3j5Q3aBea9ja1jjYlj2Q9ZtOSsgOxHLHy7HuKkegqPzglPkvzDR3BPTeGAykbwftoTAwOKzTdq
BNu8Cpc9IhYb7ZMriYIeSoLiRmENfdCYxxT3AnvBUa1u3UUdiKt0IrrfXqU7CzTyKwupWoS9lhcw
OUJzCfrw+b+2Oui1BJej8dypd+ebvy80U9m46IdNPvNyfigShHEmeOEiVtTDbEEZH1ElIO1Z2qPt
BpiYhFclGBp95qHfgRmncRxd8zWontXqGXbB8tagMy/NETV+AglSyEZd5L4onc4Jl83GVvJ0TOAO
52j2jQg2E7jULLfganvaL+rPXQJVG8ugrSWH+aaLPeMhaTFowa+3elf86TepaqxrHC7qa2/7L+Nm
cQJ0s9ul3NYLW5scfibnDAm9rmTzl0jQw0vKIXs4UDe3KkjgdSfIftovsm8Yen0X1ewSljkI8yaQ
4aVNuX0myzo4/Cm94TXomdJLyakk7SXX/ioakgMHldx8f1rjtbivP8Yw+ew96xta4cVWMa2vKBr7
av6Q5R7v0znTsEpxWkUl0DORqDRwI//V2qN0m4Y7KFPKSwfuA4siIoTcsEchVAKvfNAPKBdjld3I
6NuL5B1/t6UerMca3lAOckef3HGQ0FHMHlh9/KJB783ykMoPH0uydln3jEq3kQjAuTZcXluKpM6n
TAVBpfDC43m5lnSd5TUbOtq82CGzCw8pJICznsBqrnEFK3i02gfCkDShfJDGxaXW2se1nhPzkVBj
Z41XS9zGi89qG9Jrjiiu6HZnvkMoLxSMwQTEpKJ0MfClXMzTasgQWMorWpG4y35f9weG8YScyKwS
fv1mfcr08IQmm5xKDZoEmfpNfOv9CGBfixjUqbcbOGkZ9PemfdVqxyClmsQLDzrKmDBPomdQxabx
dHNnVKIIj1ma1sC4iZTlNMwSfqs0GiNaDHWneHxnsehThLO54h7G+wi3y4WfNY0w8aFYsOdgA4PF
hB72xVSPU4VEZBBk1yhtH1XTe0UnKdALWERxeAtTsI0FKwRvJp7kN6rFCJn/vYKch6Rylw/W3nG0
KUXYuN9UXqoIdZdFxDzPIvTR+43LPhAydPHyLL7oJhxbMypkK7QspMQ1hN4E66Iw1JHb3DhXsSJ0
658mxgu9LwAZU5rhBNqHyaU3GwcrzNfqmSIX7boNpxo3FQ0li9HRYfT40F1b090mTu0x6r0t/Cqw
nwpO8guX+q39/ND4cOesGr6VHhzmtSBSFAkHejwyAbSaQU1VhZ0V1kzrt22Q9rT2lUGj6Vb3rvsd
8YzzR+KIYNpGh+HDWV64YWCDvgErGFb23spRvULG3akQwZp4pvAV43R133Y8/mVL5jiriFOHpAwe
mwHdxchZ5OFbycGW5MZSyCX419VH1Np8B1lOY4SZkaECPmEemFSsPsW/fmMDyXdRfFT8pPMUnCVA
Woe9wUpS75Lf20onKCT2uZalDkZuee6vE0tDwPx8j3mdq1oCYIetGLMFhxkdCzebvCbc62Mfi0gh
d5o3EUR61dQhJCJ3FzvxXGR4r5FBXE7IvHQ3rJFBwEpJAXER7iRdpWa373ZJxTXFbC/eWXhjpO/Z
DY/H50TBYKPhFjwwQ1fCEkYqGomQrbdPXRnBu98DkR67ZH1u1I4PTZLZCNBSkreRCSTqGaSPiByI
rlfgXCqPTY1+h8pwcah9vTRc8Qe1AKUoBifTDp8UpYFyC53lmfKh6h6IzmLCkNRa8T02yMdVyoSV
ahrGAoyGbbq+TjU63lwn5Qy5byb0MiAqL9CSnuaB45aKRWF9JBYi1LQ3gr6OxUcdKAuHaTtSook/
ud0Rd7s5mbwaBwzY1wKY6SvMguzIK/flfJzHrZZjKMC765EAtTRYUItCj57M+dzYc0nq4m/JuWrz
wr9zy5/mmh0P5uwdRLK23I6fxLUXWEr9ZwPh77AL3b71+OqYrRVFyaNXQmsSLqCHtGxE/cfaa8GO
/l6UbzHgIH4qC+yFLV5pnbIXUfWk0RCWYJVBtn0grs04mU63krKvjCMBRiWYKN12rncZsM7WgOy5
y9gdotew+NIteyFTyc/vg+rF/B9cIyaVbnfYg+kGOb8Im3+qN7pV2NFcgpUCxwfkrbcaSV/5gs5d
LesY7SAGVUiZdoFMwQAGIpj5b86CRKV9JhkuUY7ktz+4ShIh3hxGmRgseU/swtUGxY3h7O/f5W88
kLNLU1/Ygk7jsgBGUFfrP/Tf5kYpdQ27771AgHoFogjinuKp8W8AOd5+rxeTRhBnJ93LcFW/Rz3y
OG24NjW4IlaxPrF+yFWulYeyqJk0tx3QK3Eo/L10OO3G+02eFuP3X+c4pGgUlZ1y7eXXqV3eA5Ip
kZMMOsGQedHfRnNGIqF/gVVFiSlZp6Z3wBsL6H1Eake08MDgf1i+1tYnrTpGWLzrYYsMIx/p3Lnq
fFaBe/Zl+dxtP5BXC0dMxnIfVskVtc/Nf2TyOgWfZCK8Nf2BWIQIjCm1SXklso5sXdccWRjiNroX
CL2ku25naVmfzDIRqcyoQLXNJi3seq7VyIEgTXNDBo2BYDxam/tzMeShy34wv2n4WPz48thnsANO
OWSJP9snGWmm69wAg1ijG/DTsohCIqg8e50BDXkKUo1COA4NkIkmkJviVyGwgBuhno4SZ3PYc6Kh
3DYDBfdL4adU5Q7rBfkFmwlM/kjGIz8E8Rjs5Yld9G8P6e859FEwHJw1CG94jSkSfnR2TBaYCKrq
i0lEnHH+90581RO5vUNXcC2yrlS6ztnlvLmaHpki64IGTDYzxSsiMTAsDOasb1vO0nJSM5Z3/oGF
LMxzAJKYbLmq/gEIXQ25l0+f7lfAmmiDMiWugRTeOOtELGFtojfq0Yt9MqIgtXHBcAoJFe/jepBz
UC8AX2zeWdJMYkPEvGqE8bUuYXog2CFSRaGFahC/5llHVN/B/sPPoSO1z2U8ooAhCEOayTbI+QZ/
BsmWbqZAHLVwQiYS0fgOlkj90i2AZh/7yHA2C81BGhhjho++ZZu1vf0WAFqCrwkf0UR6dWzHX2um
GjSM57/bcX4FnBUhVIHNjhUCV7EWBWsoDqxhjxDkqveDXI9zdPR6lf/BhcnPGCeK52kdCLzJTsWv
3dT1sInI5oPYjPr1r4v145VfuKLRaFbvtLuC0aCl9gBn1l2fffmPsXOV4ycYIg40C1n49WirM0cG
Q1xZIWNG5XfV3IdvLSRUAAhFAH1DHVbTra58TzgPLcC+VfijCNI7fIfIxALDTPpnhpH959yP1y43
cVeQo0pk8opQO9cYsfArjhVH0P9WfnKYuEGpzY6PzGTwy2Ko4lMXEQhUMSa+6QQM1RRQ9hKefFEa
aNZJSS++KoNKCzwxCYLCd1xyMteFAT9vzkjQuVW6K75nYxF79g3oS4C3v1MBwB3Pq7S8jpRaWRvN
FjkLr4jOkKQ9taMfE44V1IeQzBNwExmrfnM/ysfgLHVnLY32ua273JI72cxVchfRYib5/ylMkmnj
7lEfXQfztym189rF7uKtSf8WOWuJ8Zyku7c831YejiIW3YcRYVXcbEsTNVdOOelxkz9ONFg3UfUH
i6RzZgI0UXcpe7RNaxSFl3HWDD31rimjlYOf27iI0ShpKMyf7SgJWxz0feXWBTjHKHiKV4OwOnp9
JJHu4WtCoZNkl2qQcyEnDavSnbjRM2m9UL975bF9eU7F5kqIUC5vjsODfYoQ+vQEDOuFu+KUmTRB
q1xLgyAQ8nTXTtHeFFqdY7X5i/6HeO2XWvzCFxvWlPr9Zq3DFcIZQWdgV/oPUjsw3XbSdIGhGQR+
KiGBRVB6wEnsAqTyNh4sVYy0m016VxjngAIc6ZYBe0e12dMYHFmQCqo/P1KsAUnvk6RYV/4gFZQ9
cn9Ivd+Gb3+eQe4ivv06W7YH2JiosGYDQi7i1Kn+xy59O2/Q1iCXQjy8XCiOAHwsWM8wsXDkT47j
cGzxqy3UD5ebf3RrFrUa0vE30uOPh1AqWXupuYReJxEm5X8hEZP2UVh1hmoPLsqSrpetYnGgTTCT
grBn2xhMJfQ5uKwB1NS4mAIz7Mc7sEMNPokuQ0WV+lB7p1s7lR8MeXkSYTZu0/BU4TUD0KxdUO9j
MMegExFXfPTR6gdRc+ScBfIfid0zyElmbIRYVSQWJYGzzWfiPI+21+ygo8wR9f0MOgBdKHAkEL02
KsgmvWbbK3qR2wPQ7QvgZKjmg0iygkPNCtDMZee93ClWdsgnoboK00NZqcU60UhzUT9mLxZqVU99
7+hFbFAkVQS0++ggo9YHDj+LdzdnxQ9mAZCGSfMfY0u7smZ+LB7CybYxPVvHUQwaS1EJDAkjOOu6
flQ/gjhnnRZKsHwkMYRr0MnBUxA3r/Ee6Ipx9d4ABZsSJz73YexSTdmrZW8347ajWBKtaKYcpjjG
THngBEz2tHWq2WLuMnfIVoPfHStLFXcp+5iwN35rNh0W43+5AKooc3vcjZbnvapN40amPyFHq6uD
BbKN4hE0I8MFqWECON+1DxClNMF/fH90k7XmjgeFt9Nr1Cx+labwKcMFM8WbiImBn/b5vA8aXy3p
BawxVMUeeJRtUMpe2dbDDt8jEHnPodDa1zEnbu7BeLkv8dsuYMC7EywyRMLgGBFSDvnyh2sR9lCf
UiTM5o5pS9HHTD5a15dcWvN/6Wl2TXQdiivL8ipBTRjWZMJTZTsb5nwIZNPb5nyAvnXnidzYkxk9
V5KPkLyxhaoZXSF9C/VrCv3mQ4IINT+4rz2lPFFYRk9fmU6v8pVmZwRbSkpIQMoOvq7AjgUmN+L4
vVSGFXPiY3lXnRxsM41CncmEfKvOPUJRnkPQVST8IWlsYECc4N5xemhdNA1tOY+b/Qx3bAKRCT1G
2/igQwW5+FWMlk8oTA0unfpr8PvEY1y31Tjt/88f9Mq3x8nWNykXQZb1zpQBGxqm6oEDU7Gzjs3B
y0xzLZMX0S+9NLwTEiyI3wiNKROKgr9PRxBYw6HtV8ntS4/paK30ccwWKdguSYY1NwibBRmY/TQ/
SJ6XNJ3hyMkPIx3yROqNov49kZoeLyF5hcYRmXJTCQSsujuLdlJzQ6fSOBf0rMyDtXTeR9lC559e
de3r6Q0+NublF6sAfnBrWZY7FIuzEytepbrCYActFNwirrzkPUPbuTG27YB/ZAMCBK8xmsa5utdh
/xYjIxzIlDzs/qvnnfb1yNhPTpDhVzJb96nKJw8rhna2XQzzWi+mItpuu5/DFtqkm2Zb1Jb6b+BN
1JRMkOw+IBWlwm3OH2/0tkHHQJq1XsrEpZmFQuHnKkrJmVbefkTQVS/S1Q3/p2zinqgihsvGMp+v
WNiWtXDcgNYuof/ve7KvSpFDyW3i+dXcUipJ8/G1BuUJl/4XSa07Gh+1yUqgiF38u6RlUBCRi8qS
ZJNzNEu9oOOvDNWzjsMDW/ewVsir/cplTe5lzhZBnRn7tgMr/xYGeobUh1StkeckOrl796pS044W
/r17f8PXWTxy5lhDxvTaAozvNOq+mY3G7zk+JOlXFHr6UENTiqEPbD+L9Avcf/DciyPzmCNg15fe
EFOlznK4Lc2MF2NOJthwfY+TGCN0CymPjYZ+vC/sk+WldsibWugsm6iLWkM68W14+8sN6lpS+fkG
FVngkQK7fAyMegSeqeL7Agsoib5/xDmt+c/Im6Qh2Br9LThCpdRS1Ie52TwezMYvdv3ycAcSupV7
iJgPwx+t3bTWl8O2pNSeDznWdJDKOzmks1bhN5831L+SmCQVagUKlOpLumlJAp3pyXLG8GHN0fco
RY84vx6tKOZvt88arf5ItC1wwfyxT5Jqr3vwtstwJGy5hc7n8mIm/5fTzjgJZ17/l0RpblBBpb0P
Omm1DAvWP/qrwDkNLqHejJ3Y1kfUu+HqEZDLLCXPUKBhTkgatQmc1n71SR8bHBtt4BO4tOarfBPM
+uMWeuGIoKFEJu7W2J/N2aPEoamGvoWqgRkMmSdDcCQZXK3FbshGEzBWGOnaYHaOh8My2F9uoWve
6E55KvfMycx6xxi2GALmfrhNr+P1D2ftkgO22Rpio9DtkGpCcOTNsiyW/dtKLNnohnRLsJzRaqe+
hMsi54V97sRPSoPZTTtiLADDcxsqhm+wgusPAVtVixZC1k92G6M1CDqbgeRprYSkX9bYGoUkhyF9
O6gN6u3SyZa4WPIYrImDYQHhU1LFWEsgRZnXEiCBixgzWG5zknvEAIkrmlra0IyUs6M9Gw8Ikja2
/0XfrwJVebBVPx1SMA3SexM9KklxT8df++zF5al4ABE5Cv4zipbkpBhBQEkauemlBcLUwj+oaWY5
x20ius3kTa1ydFnTFId1c+FS1gSFcNrjyCTRYJGVnLtaUQNneHaEYIjM8cnOXBVrNwHiHrwqGr+M
OQDLemf6p3KMVvO0kbjt8Pi6ajSY5899RKsjPCxkk4ufRRA4gfloepK+fVx5mceRkIxyMLFDY4DD
ZnK1xj/SawT//1/Otn4s5yKMtoVPRWjxK7vLGFxIB0KBWJuuSQ6ih4nYy5psDeN/+m+xx+SvGv0Y
Ze0jdx8Xtldh/PXwhhNMqsl33QWSPDH/FKs3xoyKFm/h/Y+cAjRVia5q2UhFBeV7jA1jxUlIGCni
9qLRgzQNfpZzHpbZbKOqDYzk6tWNaNrxBsXuHfb2UBGaVYolNUB6662UnK/45L77dc0o/RO34Kf6
NHrH5LBSKCyA3bk+4AJuKkZ4Kucc2y/jdP5QNZt0q4dGPCSyMAamsyuh7EZ4PeslmZfXtuj72llV
3mmVVxQ5EIEGOc9unNA+iEXnqimk+s50/cCykMATDORyNALVGH1tdlz9NuLAWVi5cC2b8aRScHjl
0TOkhJhQ0mWiUW5tO8qQ3oBNFUOtaVyNSTPmCfqDOI1HjhhKMGlpBkEcjmJRZhne3mpzNAq/UZuW
Vsk+wUKV+WqgvUg1QS8WzW6KApGuPwMzZMryzxxgJaFG6d/0Y4F9wh6lDpUBArdNbQ+n6+n3A3su
ExGcDyy6Qu/Ug1kmbBJRzzyXqtrbAAcA0y7M4jua/dDgbv8cA4LnH3rVfM9FOWt8sJ8AAFnq3dHq
srFajbfX7qB2nl6HljoWXTcvxkzvtoHegZwxr6o9tHt+6qcSP5L8xBWxH2U+H0NePHdUQ6V6d1Sq
S4x1dAlotUQwiRQIKUPkRu2WlZLzP1ii1jYYcqAbrHdHctxgQTJhQqUrsJc9GZCkjqvp14O4BnrD
QsKd5hxkpYmVlPW5uIV0+oGLJxi+mV0ZSpD5npMH48Wc2Bz/8C5hRGSMxbJcWyJ9bmxLglE2N/aV
E5clt2P1aMB+7ur2WoxUMdeoDXPZ0e2TlpGSIb8oUiW5/89QJDW79kR5lxWqmiFSUXYFTM4++3UG
ZB6XCFlIDuCE7ch57yAqxrY8ZPvRXq3QDWoTsIXmXNJuJISwn9uzFs2PJZbgXOvGGWB6HimUZy6V
XymezNPuOhS6geAgRDc3Bj61WCz4ZC8mhNai8bRxjkjDhvEPrLByoBuSyD9ny9ekvytS01S0Rx5K
mMpK1y5JRCyBCB7Egm46VFkzk6YGkmvHYSWo4IRGuJCQNYBW48GsENDPcb2HM/wZOqGkN6lnT8Tm
5VyFbf9s31qjMvxwiPESuT6I228z41n5V/7Dm3Iz99NzT/7AdlVhvRyLxuJJMO8aT2mWUXWwBJ27
pxe8gFjGLM1U25KAf4Z3cNE1/Kf3r4navvAfFlT7KkYLHpqPnKrNeYrBzgGRpB7r6E4YBwrO4K9k
PXJS9u2fc9yVrKj0+Ev6To1MTo+tcAd/MRX0ydPu9NZvHvjl/Gpe2k7dqvnoP/BZU/i2YDH9YPDQ
X4iin2sOODHU7H6Ug+6madaiOdSYle+D6PIJzec89gOKs0Y/l30ImXWpKr+qtVJsMb+p/r48gP1n
xSZcrdVNcWb8fwZJAY1OI2afp9vgQ6ngr8kHFyLu6DL7AbFLRZ5g0DBvH5EKVmHIAp3/5IWRbdDE
yVATVdoDzDu/LpF3DWmQM/2b1VJu5t/y/x07pKzS9RxpFMTt9Hzc+30v6bv185bDSovKaF6vsjsA
BLL4kMVK//ZRTaOeC9JvPI3SvLcyvTXooIxaXLMN6Iysbqky8afkPSjemm9tEgRhpgB6BM9aZ9hU
lZO0oWs3w+e8JoKA5AUM82HN9oKUZjkuk4FnuExgGII4dCapgSpZobBSwmv/ak4jPTzy54Eb5wH3
gYDkfaaMqHyWWpghKGVIUdGmVa3Px6rm7BMeudpzc3w+7kApJpjBgTCTHviUvVVRtIPFJQxvS53h
noOqJ/9yoZLt1XhUsF4gG2L8JhrCMwuSgfJJpg9FogeXAMO7kTpylwsRIUoszL1HL6yHapIfY2v8
tIxjoqw2R5D+LPH6DOfV/dg/iCoNwGBQiQ9AvxD1qswMjsGigwmw8Ak6c6JrMheD9BppXW/G+Sgg
RfG5qgFSvIyIpDLY+zoKv/O9UgPudt4ogTd7bApWRwoFSIQueyHYzMhyDX3nt7utqno8B4iet0EE
vyVlWKRxIYqeaeFVFUzoSlttfMyPQqbmF6DNJMMWNHH56cMljH+Bdt9NP5m3Q4VTeu4RSdBtYde0
FqY97zLWxWfsQEDKksO7ex/ARyQgIsrKVXI4zcoP0Km/HMN3cyKAItWXLtcMQHMyzj6TDVgF9vAX
aojFSg28pmmSDGJ2B5CS9eaD7cDqV2WnG8JnQC60pGusPUIwf3/tJ3wDrJP1FjZCBc9qKvXsqzBp
3+CTW/G7spjeLLVAAz0OhuInVgT3as4pBJY4VVkWgXzV8vhlNGoWnX5FteO8uU0Kmj/964hv9r0G
0/8QC5cIr/Z9WgFRhwjjtSr87WLETLWLefeQgSQDj72sB2dv3kK8FZqAfIDHlnL+1e4r/C+F7cbJ
GcA0FyeYNMpIEEBJj6SlNPDlf1DOepcnHVh6ZvXj+Yb7Q0b7E3x1JqkbI1pXGUgUGw+OwoZ5Ctiw
DxjxqtKX4FKU3ktM9z2riUVMkYFJuqaxwu5nx/FGaV6O10xGaRMq07tMpdOBl2tJ0WhrPubtCuuA
hAEQ8gCqGt0iZ0/853FS1p50jaGcxHDDW8Yhp6ae5snaLKgJgfv9T+5ANt7amJNqx95MV3g6GxWe
9z/UlMIvkmkW1RNQZ2kfE0OEey5bwCuxcsODIhBy1RNjfQW8G+LG1wfmu1/eTfoFuVnp4pUDGI0s
nvJHlHkbM3qppzVY26PgeY50I/nnCHQL3Fb77JOZrXrPiFcIzcT+UhU+B/cS5CTDqBN/dpAbeVQk
EiBnwYiYhoQE/sGIsU5LaIis9qiN/hFSgXxLTOZZASZIiOj3iipAgpX9f964YsOo4ZAg+bmt5d3K
rGEncrihfTOagmgJnjtjEKWlwIVqudwKTe0Uxbzmh6MF8A94ylXvDQG3oROnFnWOpVVr+VtJIJ0G
11XUhQnNdMc4ukfWknHEJxtPn9IzJEfrY+hOfpnhVZtrF7RQld98Mnj7x0Bf1c04JCT/vorgpG3j
WRVowheEScANEzXcvhvSppz84aitue6RmOkDHK4LhSqjHysqQY90G0fTFfyS/Vk0NBxkIPwSfb9o
2Ew8WzrybJsIM4s+VleVCLH8t8+KGHC7P7MgCXIUYrIbFu+pV4xhQv6+H92M2DbzcO3U2rAZ4uOu
g8xeh1DFqpHkHK18/PxSkKZd6GoXw/4oy2TfAgQvc/ctvbsw9mfw/jOXUMCdAaWSW+ZSvClxcXwG
c2xsEKZG8W9jASjugPJoycGyRpPeFd20It4HrtwCaUnW2EgKItBeppBfHXubv4Nag+icLUnUUV7M
5qv+0uyLdIQ6bIb8j1SvkqTUC94nk3HShKV6KkIjwwGaVEYt3DO7mFmZoJ9k+0dj80DB7Q3FOBKY
KmQhFLIUFw97Uu6Rt4G+2DuxmQ1K8vyd8QN4s1wmKpreQ8mm+qbPy/5ZsFKm/CGmthHX75jv7rv7
/DGJ5qQdg0KWbSNJrRFXJ6eTbn4ak/QDej/leFa+uJL76zDmcAVSfaeTlD/ye4JsdjyyBWNgjSQM
z7d3AsSrspELmVNCB/MwChOXxBQH7t9pFv593VUWZHrsDYTbmjml/r3blGhqOYBgHQDCZaiH4EWl
4KdbdBWZtnjLhX4t7WrO6+54q8oPsXKNhNJx2W66xHEb043nno6vjYmnkYzdUgA5MijzwBCTuCUS
eUnZ9j6h9tdeo69EawIOPQGCYs+R1NoSmB84NAlHPRQ2KYagLj5kXImI6207dfquyuAHnmOgf2mG
lky2DYzwc/GEsSKzulbWf8ArXXpahmXAsvY+Zmrn6UO19SXqdipP9YTobyiK1vSF4OZCO0f1o0pN
X4isHTPBHQZhRbsWp2fflw7FkiSZBjMqc1lwbYveEf72AWmxM0FcNpd+wMbGpbTLA49psagMfPnX
YCQrusoPAxS675KotKk+/FmWT4gaWULaDPT7JR+phQ0F0YM3I4TIMneyGIL/XkG3TWL/eELQ6S8D
ZGZXgj8dYrMdOrdzWExEgejIi0pEqQUT/UxCNv8VuErOJkZ3YCuzCvFoobWPfc9QKlOTmvcb5Pf5
jK3BLYC9cqWsq/w9A4tjl/IlAzfv6B5WsU9R8iMRbwVin/6eIT8Srq37gFQ3tcjOpN6VXGFwKH1M
u0VfbDp7DPQYpmm8qSOTAB2lyz6ggshHqyRCM88+5Ey+wOUKD3g230UEf/KGGZD210tjLzj9dfLK
IGIy8lsKu5V9qEsvOJO7oiX6LwQvxjnbuB61Yas3GiWAAH7Hcdv/F4liu8dY2YPXIlqN1fSQB3cW
e2kqunClBCRo0GbSDjybqEtQhI1//67MQTQoLZYR8ZElWHVwDHuew+n4qQgAHWcaAZ7IivYeewfX
9g174kTxx9I38THwpLe1qEa5EONfCqmzRh0zqH8ekG2/9++IT3Li9QpwgB50CoSCMaM0J6G9XA8p
n9I6/8DWa2VHei1hf3igyiacXDp03+JJVJhdKK5YCsbVkbNgXR3ezgSClhKkzaBj+EBBOVyrhsyN
g05zDj+RpKWUuCpYReKSn8iGRRF22P5gHC4sNFvSmS58YD3ONpeMM+EMEQpeZ6B9vgRpnrj5cp3o
Tjqi6bKfeg4wZ+OP7CR0TmwSjQfSMBljhC4qKUywuoeH5CmvcOCNVCdYu/mcnPNDgTwlhTh7l6oq
Qg5S2rRIH6TvCuwpzcRPTtBVML8zKgYDmZEEZigpnOdVoZu17G/34RVLPMde/drgA3w6wOypvo8s
SWiNTBLL/0VNoU9R8aaJZzBk9t+Q9yaOKrwZtxeWlGzO791Q6eWOjxt031jOgPIpV3+tMDHVKObQ
b94DZegeIY6ye4B93iC4qgmklpoQZ+Kze2RefBbBxx43jKthcxCdCC7tQzR1oLpSjFadVOq+pBuQ
2sphxCr4oZA5YC0aaYS4z4gactT9u6bgP0W4VftAQ8Cq/RqMsD1aLAzp/B/xTuhGPHRVKTO5InOf
YzZGLeqXPZ1jZipRNQzcpZiflJApGsJpDzKB8Y1WYOQ8GGoJz/PeyrJv+LlQankVH9z6YM1Wi0O4
/vVxtHXPH6yd8DD+bmDLfvF/GrCLhuQlKNAPobrWxXIJTQ20jBpYyj5kdnHEC3i4JrMzQKebArs9
dhYZKhGZjaaL94y0EIx7tg+vlJ8vyWjHpwBXrLoF9spyXLCQNaPx5/KOIY1eOQDCXJgJCGsW4YkP
biuQ/oPJ+M/REVLTmCWD0LmXnqxzFR36RitUyP9wZqtwbZYWM27BgqHDDV23ZLsmAxM+XpC+G8M0
HdMLieN0fBewZWOzcTvwb5O0SA1D241ijf56KAY6ubDWZ8DnMx5JeB6L7V6cZEoPkTJ/rn/mmaHL
boiL93UlPy7G1nfkPH13UtDUUAmu5ttuvLjUwmvZ4f8s+302vW1WCBP6kMJhcSkTLlq/NJl1dTkA
1t4HknrSBhoNwO0JUIyVox4Fg5Xg5n3QkyPiNFoK+stDfkSHMtddSoCC5hWhKTcffgiFa3n32p+t
iMKWLfFf0+xevRrOBNgZKuXIU7g854uzWQL6ayZq3RDIYQ3GdAWHrkQvTPKucXBXpjVwUIZLCMfd
XDmzgPdbZ6O2EpJz6khtcHwdRcFtoCcrPbcZmlcXwBEpr4ny/1UZjogQmSQCDwkrjQ7Jnb/MPR/a
GzkdXIJvh8hds0vc34R5K5SfCXpqGjI/SzFThBZ8BfOClnj48uFHsrhOoi/YukEv3cPJa9Uyg6bh
Gaj4G7WKkENCgFRAodoLwAe4gkeuzGwn5oMcijMVZZI/L14Do1khN/a5uJXyZWeNHPKBffoJy14B
hUYrVgRngcIgiKdWbmepoORrCgmWSmvXDgdecWlcUaGNRJ/GmZw8Z6UP6dSlFrBNKkIj41+x44A9
PPoueWWCHS/kpAMAQgtc/ezRRwY5wRG3epD1Mc/UzPyq+TdrjGEAhaiuT5ItxgL5BqovP3VxDqKs
lT39Bp1JngVkHgXZRJy2kZ9MjKQTuLdblGZuL59zOK7e4ESkRzjjS8CgdhNIhbYyt2pegyTOgkTH
WSQnxEGkns8gjgV9HP0pdvV+NehgQXin/H1alb4OitcCfuP1UxpaVv3yiu0K54ofqYWWd1CYSzQq
RVEzGEYQ5/CWe+y1s+nrS8xEXYASqPk5elbjwS24o5JomI5Dda3yRjbu/b1c8XBISI7g8P6XV366
SU50oIrEDXeC1tYGAekHfZiQaGHLoeipUX63/4FtrDAuQwalkWvrxVFk3n8wO6BolcKu9tBbBTfJ
2w6+Bg+Q3lIRkao1yae+Qsf1aRvkMlY20UivAylVRAAR769rN4h7d+sN5FfOLMxmXDqHJ7RSTstR
diVvls1Uro6PkZTLdRMH2WBszGIeoVuYEGiHnlQ+Az+uFBCh6MvSYEC7aZaUCJDG071796rio9dQ
vXYhOvCjTIDIkHTfTHUK/5H65oYWTLzSLSAL4SUP+Bw2NqqUZ6VtLuGEiqJhLIr+e32HEyasv9I/
NejRrmR1yjgk66iTcCxH0wM5qLpvnV0gOjMmeyNrzKHjEBPHhvidMdJK8Ef9tbrWlmpRycz1XRgt
947ML0xoBVAGtZXzu9C5VrgecitCkmaYVsKqklMs5qGwgazs+yXysxe8jb+jZ+ieBnUGd8wTro6B
hbzssFBnu6QYnrG35EGzDGypSBxZazqB2wLiPHkoSIgIx1sfeJNZzvCB0Khv5gEyv0/OD/xGVcQ/
lvA8wTLUCPPND0giCHEwTZC7+dHsb+qdH+NsaksrmvcQnIBtOkk9WH3Kqp9r50wCl6SjcFXpZOFm
s8H4ETm172mW4bp1otnRKN7gp2sPUc2sRvxCvaNdD0a4tRtdqMFGdz69K57kheaHQ+QrDqMlFRfT
J1jyLNyt9uTU2uVRPKhKhIpcXFvhK+NpGII8w2uY9Lx7oqS6ZCoNJCSd4Z9ZO7lZ94lR1N2WwDcy
8OeUnRPParf3S0/REv2CX3vXuaIykvYXI2DuMDe8mSBOeRJ1bSDz1r7BfbgFppvFESuJ2Z+JeX1o
jjs+WDusJCxkZbdX3KU9EDxoZWN3cyH1awVFR8Ze4u2gd8dsnn8ZcJb4RSHjHGE+3aOvtqLDVYkE
cykJOfi6MXIYk7/IipYKzIJdQijIsHpCxsvwFDiUk3DNH6kzyY1fFMPpwvdx8h+s0B/irh3SbwgG
TOGLFeCV/LZn0aJISIlBERIr4VZu/fpEbrfBSK5ZUUPL5igNHKAUtgDjH0c+Iy04wPpUabpIjqSv
ahFqkSjm0KNRcvEtQr0W8mYmkpD4DjL9g96fQfM6f788QA3Hc2LE6a7HQ8dmwtSIW8tji08OicVn
jxdmSpWcXoRkyP2J3LLuPUdUfe0fNF6JiS6D3HgES6VddJKYiHat43WSRfmFaG7gVYrGkcjivncW
zXmzwOTa+kBuYw+CzSl6SLSoO6GPw3+lQU7bv/Bfx38GSVNvWIHRsKgnLXSiEsg0P1TiQ31p1bcY
VdLanC0Ke/sOSH/4KTWpjnx1D+h8DXVD8qdkj6WAhyxt2mpvJ0+xvYnNVEkDi8OJ2zZ8IXMFHRQq
2H5HI9Rv3+6YzTa5UWHeLkT5pcM1+fUtKM55A7O9qRZlmxNwHl+UYfZiKIMH2R8AbiuXcwGviKG7
8PK2bOMj+DP6lPa5cQen4SCsr/VWeqm+BMsO4kehRBXHyLu/NF6SzZKoZ5Uwp6Sa86gym+R+D0SF
5qL7VakLbFIEPUnF+sXRnHrFORu+0pYk260P2nfKRDcwPkLggQyjRdkLdgAe8SMbIPuWFqMgNmBj
xXxoM8IHPTBwIFdp4jGNdNhFyFRKu3BWH53FNDu7e3pHcR8c9KiNgOkG4Ze1kIGSvGGQGAJ5CwwP
ICNfrslA62UdUV8pl8At3fcTAB3m7glxakHFnaX3UPxSDv3nxxuY0HyLtYXMEFQ2+MAOfmfGFeNc
Jns6U05zX3gtxNb7Ifn87Ms3/icEkq7F+TU6NjmQYr+uYoRyGPv/GQTONBpSH+T8A84XpXG5oOxW
eAHjLKOfGNMc8d6dy2cZ1RMCTYW8NNQupI5WDFiGvIv62MONlKuIN3F5jCJzKS/FAjp4UpCfdR2G
zpQgJ+KDum9TL8nqCq4oRmADBhBBJlIijt5VzFwGXw9KIWhempnkfezJ4f/BXSPe3Zn8IVGwlI4X
vKB0sFhp4eBMxS8YWqagdFJiCk7jdzt7KGOqVmfquQDULwj+TdWEyWYIltsSJCHD50F5jVP4DuNj
k15qluYHA5DAC32t87Bhb5lvhO1AvXUPvWQP4RU2QtknftLKcTAF7nj3MDpy8NzUnQR8LehTfzBI
adwM03MuFqRMV1nZ+HcDdqyWxc/CmysbrmwOr4FUnuM/ys7PXNrJTXB7LsTAwXZ682jB9IFCJM1S
lfvzgsk2CnuXssN2XvpVf89YeFXuT7gptUWuugCIqaU2diOv27BIbCsD+Hv/hDjrR0ZmFZbUDijS
MvU6zudyGmcaDK1FfG2OJ27TDboDBKgP5uDKLlXa+2k/hmIYtd7AKlgtMatlD30Rv97gfKTcV3bY
JZyLm1nugoQFlnOVN/qy9fg4Hh0TcBLoPMp2Ag+9MAvj0VNjywNFEOkSDOhKeWGj6lNfyaDChyeU
oWn8RhY5gOEB2UDLjB5LcK45xgORii8/cOGydOyshBXWu2/6h/7ZEaA=
`protect end_protected
