��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���{C�%�P��%֚��	��3;�Fr_i�<a��R��\�}��B�eO��`�t�ZN�ˇ/��m��Dq;��C���E�㊷9n�k�N Q��E�X#��3�^�H'�=H�6�)I�F\	��a�p�0ޱ�i75���#���C[x-��u4��L���aI��7dJ����?�7i��.�a1�@��wii��d��_S4t��" ���C�%�8I/�cnM�;oǴ+��\_�C�̸�P�!t]00�`y��)��S�|�P"2��X��I7i�@Q�]��:D�I�s�s5S�f��]�@�&)�چ��(��gT��<>�`@�dg�c�H����;Y��k�Q�L���̶됥���L+��r;�V��%�D�Ľ�PDx@ʪv��$+"S����d�R$��(l��\�@ߣ��������'TkI0kd�<�m/�0	��8N�?ڍ IMµ��f�F����w����!��m:�<����H���B!����:z]��푯�H�Qږw��t�RZ�%�x�"��'���?R>�R�b!�~��� ����1:�^}�Qx��擊j��Z8+TjGp�jp�8�g&���S�!AF��1�d\:��/����B��A�O��ҥ��˭f&M�gܮ�����z�Ir?? ��n���w�x���IH�Vp��cXB��Mk��(��g�^���dG<�A�ձ�Ec�<zv��}��u�
+w����7�sb�X�N��֩�W	T��E��E��*�b|w�RC�Me������p��bZ����� /]�2%t�R�7��|F�Qm$B�\7�º���r� �J�X��dE�Ž��C��8=�I��7P�q��OO��[�c
��j�`�;��5qܙ~=�z
��������v:�N��ZD0'�=�W�DX0�q�S�.��kJ�F�����E*;���d�ǋ�2Gn�GH@��N���S�S��ִ���Z�k�9��:b����Cc�a�/I?�ء���M�����_�ܘQ�j������>����k9�j����I�����oVy7�O-��̾۝{,�M���ȗ)�������s*?wi�G�7�+�Н$��TP�=��Pꀝ"D��L�'�k��'�f�e(~�)�D1�FyCKA��}�>h�?�"�7~+9�*l�	pg+�a}���5�B%ooٸ,|��Y[�C%���:��8�1}S���F�c�)��R 
?iv���.�3I��m�\O	��|ܺP����o���JyyV�R��Yn�k�?�6YTi�~�r������n��u���.��ij�tM=OE���}��C-�I.��6W��(���f����8���5㬯,�W_��1�c��!�１	��FA-_pQ�+;o��j�K�6G�M`��r�B��^�*,1�>��r��$�E�ջ8� 7��C�X�'ٯ �K���k���a��0n�.�^����W]vR3��L:8M�S{���R�n���Il&������WQ�V(q��TN�#��M{�=����G�>������4;iˡ���$����J����u�X��"F�+�c�w�kc�T~ ��y���$=E��Q���B�oQj �5$�2���������E�{���iY�C���{�՘'��Y->x�9(��ۆ���Єޕ#.�f����1�9a��6�m`����<T�qK"����q%��K�R�yx
�0����A޾��a7q�/}G(	X�S�'���u<���4�N�fb�އS6�v|�rf.aԮ�D
����sRE؊(�Yy4�t��C��F?j����3�sHj��� iH��y %Ý+{o�U�����G!����zMw�ܣ�{��������l�4y5jw��UO�m:�փ��:33o�9�7-D��5�:;UU�d�a@�q�R<H9ʡFz�+�=MhS�/*�����n�ofއ���/����=c]�{����U��AZˌ�Ŧ�?�Q�Z<M�j|��ޔWy����������E�
!!�w;az�`O�ǣ��FY����g"��l}y�=��ԣ��p+=~�j�vf���s��`�W�J&�u�����[���Ե���F���@N�-����s��c���:1z���S����2�}_5��;-��uBjx/j{l"����S��S�$a~u8����DG�*�8#<�ht.�H���)�
�Z`%
)�R�F�E��
�l�GC���i)�f��Jk8_L�ն�ݤ�~�J�s�AB�6������#�]�(8T_�9-�w��̘}>3��%�����~o��3�	a޺Ք�X�X�P�s�p��\,���$�F�$��j����K:I�;g������ʥ���6t $ �������/DIc�������\�ЭcP{�0����a�^�U�O&I�\w;�L�k"R���0�I��':����BWy�KA�t����g7�fZQ���%�4�CJ;^��Av#����A�.�;����z��-=i�bI&�[�bu��v?b<<Aȕdek�q��r�X>'�h.��y���C����)��N�#K�$P�I��c�h��A_�\#�Ij�������q�u���9g��q
�S:�����R�E�O4%,�GX*�|������i�GH�4DF�?�'�K}���"��FU8g0ǆ�$Ņ&��9���T<�+���)�M�>�~$��B@�r�U�	��_��;�LB:�T�Rh��>+�Z��"aLúQ��Ư���߸��L���B�Wk���e���.Ҟ(l2�%�JN� y�2GE��zg���3h��&�(yC���!��y�T 