`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
O5/5YuiQ0E2Ez+PAINtQ4Xm2NwBGe195ou7lOLpx0YlDVtT/gUKtRGBhkZDrLD6JF5eMfxlOIRbq
OvhtpYKqHl4qWFEk6u1VAks2MTXxVTExjqwwcG0OjlWJFE+eEciqYFoPzcR1Jo79OGfMCQsTfHMP
4KfTJ52sqMfIWTbV7qCuFDk12+dKXmrEhkivQnUrh1iOESnpTlT4lcfOV+CLGU3slhAA2vTd5B1J
minuM3lbE77v8ZVPZ7X5ZVULe+UW3NcN2IFPgH+72YB4WxV6kRWjJG3df+TCS51aKHaelOKC24/I
97Xs+FWoNPfPgkx8JUrOqS7eaT3jbGTPARqyyA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="1sl9HY6tFNUyKhUO91zG3Z4FQmWyyyb5EI1l1rhL/AQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2160)
`protect data_block
q6ghe13uz9q3/mg3MR8tyVLCuLSkvpNkDMhZ2m9+GGPwERsKib+tP0Oh4CXuwR5Ol6EpN/WyndtO
Fn0LIhYqlDJrLOCBMLBtGt9N0BYfnrhSJ9rbDEfuQhEyh7oxlYoyTQJEh4oTK93JiUruBRF05ic0
S9jYkNfSKG7syV8Nh7/6DJDk+8GiZa+nFBvY4IE50BP7ctrLC81dR6iMcnLoH0TN2bYh5z2gATtQ
xPT1SzbhDG1+zKMAUIkvAxHGePE0o7nJgdhrO9i3TtpChHjpyklpmrNfPjIjay5xRZ9Mig6snonu
6lQij8ydbpKO96LAQIEW+jVjd/qwpgzEfAiYNhkbSaNbm/XN7Q9RngtFue9czh6kAR4M4uWCkqCs
ralQaH/qCw06eALYzCCl3b8WM9tM+vPOJjsI6xlLN8xGAXtMg9lNpvHqUyzVu8m2D7kdXaGN6x1j
CT7LvF76kvmUlOOExiq0DJYICg1vTXGqR9je1Ph9SgoicEDsVU1yjInF4iOVDb2euS2WiPldwZlb
6hXyzZ2/UjpylQlgCRVr5g2pi693ztw3j3QPGLKyM5Aoo8yWzT6ymSnWcDJDap5LGMXq3Vd2cal3
7GUF4wyK9r7ZWNIL/ioj0qsptkE2wRKAmQHJgyIIhlDyHPl1kVxqOsg2THv68vENjHfxxlG9kk/8
xE6qEJfUHwwOBL1N0RifQ6413OwoH7zFzrAKjeptg2E15y+v9Affm1eBj1rq9OIbPwNdv20EptFB
sxoG88a26Mn7qst5eSKBckQwvWPoWeBJKgQlynTo0X8bofMQ+ggTQL7BSjjHPwxxTAKFUioh3hKN
Kj03vOaWr4MvQWuxVGuxYa6cn88N/df/BiC/QkunmD5GyyM6xGVyFEYEnO4T9cUU2H5nBlhrp1ec
znvEYH5/yF/eFEIYoiBk0Eyq84bp81cryhNY9HMTPwZrwy1vvQAkCod2Vi9Vx3Yhi3AtxIQyiYgW
KiiGTtHjI/oWKcpAIpx3eSL1BrANiRhytnIhxTncYbJA+DbwK7jZVarbGoPida7JqKQcs6bMi3Tt
WcLHqOZUvVrgA6Dwk+aD5gnJOh3KCMhBE4YhufKYgROdHoJh3u0uAGBA1pX7E0TTLoSolQ8sBNuE
xpk2Zu9+9CNZDUV9Iaa0untbeHiUXKIGpyBtFY5l0tp8U6WK0kTYeKbXwQyP1bDZqxgVAsrWBzI6
Zb2F+3dgGW4P44ZuHwiwIUnw0hBafSElp4U1zCDMt2jrLLSHE1YbGRlQ3Blb9S8vwG+LTnnFVE4A
MCKjZCi2LXYP9jFCDe76cr4CiRePAjtkbGcyIQPk2xSNI8HPbLeQPC1AJZikf2wkDpFn5Ywam+mr
71H1caa6BHwdud3W0yQJr6e1PXY7wuaVFPl1x40xP2HxpepWrLCe9cImL0m6fuTT21DoLuHvwrQz
Y/douB40C7qs2Bgr6Xvn4v5Z4KhfJlIV0ojbVMVQQgAR5+6ut7xKDKeaWkQ//5YNFaZERovJLvZ4
0HsvgGJ5weQ6NqpWc5FtGmENuz0u9V5HpTHBTBNgkiIo46TDk69sSMWLIV5c4wemYTSuPnqLZPtE
oP+IYBdGAUJpQ8C6uc4hZctBWoJVU6w0j2t5Sgl4tMBPyflBtXxBbQDfUNeGDJru2rvTZLZrcIhz
MtcIfAFeggSkFCR1HvK44nW0hV2bw2RcXzOGnE34cV1zR11hD6GAmnaAYUGYnZfxbAJ8ValkOnGq
WObTbfpauEKPPbX9KI7JLvp1DsWrruVYg7Q/5okNZIOflDRNfi6TpYXD+ZxTIYDIkL4EKUSa35gQ
qcgRPPlJrZiAazTkmV58ZAOKy+jNuGknAQLGSxFMt2ou8FVXBmv5mbYrhmqs12GhdUoMvSSn7lK2
vV4wwjZ8O8SqFQWzkja24J+QuKByyByPYZoC3xZFhn6g3RXIIjat6NOEVCRNy1W24TSG53aZPnYR
+D6Qd3zFCPs0fZCIKi8WQrxxQtcsDLpAtYMpy8SWS/XG1CZNcuVhtsjV9Zqfp7/ql4Bqkl05rORo
O7j3PYPbryCgerEyBtI2BLchnX4vXAN7hRztI7BoyQkv4vTtjbBrPDXZo8cYiBKGOR7z8DRMOS59
psHD5KcFkxAdHweIQHGXiVOaXp5m3U+KZBpELPdErQSRncM/occCurcZIjwdx5osiex6JFPnvdby
E2vg0bPYi6xJ0UiUBovliZiVmLtxvS7cWJ4yHtXs4+r8FpoBgaZnsiS7wchpD84SPsZqD2Yy5DNl
iDmsq3AY/FV8Nccy6ksVygcj55+zT9ffDDjmgb7LDB3WckxRTqbYkWN+KRXKnMQNo5cNVJgajYQr
PS7wWUDwmMkOQ3Zs0PhLxDIWb/pWCJTJ5/6DSGosgDcLhAZEKIFr07Dlbh0nGNLDoVKIESTVl+aT
MyCTDfdvPUMtNV/MvehaujkMW68wOYX4jYEgT1BWnRSD7+pNpFm2jhlVcsM6QlOi4FAzNhNIBlFV
ve6oRAi9CtDJrlEagJA2VTNzFAtr7RWO4wRAHe+ypdFa0vQEFQIWdw27LFQy78vfPu/ZHLPmHq9p
4HduJWFk4CikWaP4ht2rKNrfhcRkoXX/aUK3xHUE5yGJuvca3J3Iuzi3uMg1KlgzU5SFGQlHLtzU
RdXIcGxdXIQX8e6vn6nUmSCoOxFbaaBp6SOCN0NRj+c3EQkc4aWC6Ny/yywCgrQDk2/pu5UBOKrK
I0P149uPPsnirEqUY2+V+oaMdu2WXVUvo1yRU/YxnRNmE7xPPXXIrMtCNtuyI1msRr5ybucKEa8c
XpNXEAjL+H3Aos7GHdbEyqCDMe6tAQxnh2m/0gLBFut0whe6PgNyNAUteCTW/1gaRVz3
`protect end_protected
