`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
6T6UHGVlgilVNvAbegfguONoDS/Fvxs5WEEtF3QvzEKEj8k0JqyCXJk9IrhB+CQkNCJ580YKXIzo
H5JRrnnPJcXu4ME+UxKv+yv2tj9+/91LiXXvA4tanJCqOCZR+DqNu+JZlgYdyTRGm1lrFSR2bVAn
k1jBIoKEX1ZLSkuck0HdfZH73r3z19sfdUDMTgRNIsGMTkdIkEauGt4MXVhto/SmWZFoU4CdZ1cW
UbOLtPeiem6mtkjtAI0AaHgNSMIHUBCvFazLXr2DiQdUOctkZl5PcNOIF1lh339CFRMkv5tOyKzr
7G/gNptEeGFuEnP+Z5x6oDvvLfG3dC71wX0e+BYjMQgU/4D+TFeFgPmJIZmZM39b6Gm9UR4jMRoz
VAiEYcXCcJPfcBSv5v4HBxSP6z9AWCv/kwvo7GDRvpLY6wUTG8BAzTrm/vaQVkDJJXjXoiFCH2dn
NffyOmleRPIxJNowHdtQuR3YFH7Vgru+LiSeTBFMNRr2vgu1tVzXkvD3embi6nVww7Xzlvh0s25W
/4TaRME3Ym95W8SAtEP7+/AjDNCxfdKW8sqxVCwWw/SSbUsCKKnImgeEirrW3lbZf3gmXq0wwXQ1
lw5j086rsrSZn3R7V+Cbu2VDsw3s6DJPyaktdP91AY0bJ8J5pyap97fN6630hZU+feWSl/ySPw7l
MHh6RJS4SjHyCGCOfR1C5jyUZwPpxXG0kUNF00e24rlBvmoa0i94xQh6byYQGa0Vf/Y4O0hHB7UO
Bu5JBLhxJpccVjskUN6TAsmO7nG0stwY4xligEaRjnRc+9PMYmqXKPl5geTV3fjaP4ithyKNYnxe
x9ipKnTQLkhfJJL/7m/B0H2g2ioJehAaBAdyoIGM4d4YetQZnL4LeJK0ElFCZl3qwrQW0x/8tOQj
E17Ovdo/ZA8fqjys5slqJCvQXDDmikfrDcKIC2egU4/DEFPm/I3JUYUBRUedZR7DPJm14kyiBEcu
R4vN71LQovsmWV6Jb+7Xn2O6NrtYnfuWOg8P0gnDhMe5fp1zVFYfJZmsr4i8e4Qvriu4+/RQYW7u
j2qt/oLLhQkQr+KV9HTbGcb1a/LQf0NlTR1RfUxN7xpU9rb7GxuSObz/xkZiGUVJz+DGJHYAsHb3
Np6ir1yaxhsj85v782NUsslrgZjKe24G78BqAQQrQoTkOWkoi6jwvmjZ9p7OV/kUrMWyzmh7netA
puTMghbDejhozTv1jkVVauF58cFWyJgabF+SIVr6uCVsk3AKW5aeJdniDR49URQ1c/41umVOXKWM
/lVxnY7zObT7RFZTVpujC6jaSvrbw7+7dthk/+1ynGMBQqutPFHa5lfxmZqZHox1gQmA8NCpvLCv
W2XMKTJcao0PqSKRC8pipOGfHNT8peED4BFJn7dFSaHAUL261o10gpnfHaT6AL0e+byvfBEGXgqa
oZeKns2njiaXqItgJw6/1jjTs+8nfaR8BH/9amSy4C0C9218k5E+oGGdvBI287RlQmwtWTvgeXcd
4+5DLHtE1e+mgW726yqdnPXn0btbcv6V9qygHg2MXITcOC34av/1TZ0Ua07mbAZ5/UKcIWxS0Buw
bzCJ702HJiaP95CJKM1SXjwmfUjqmKwxnRPz0Q9uV9Q78+he2TTxpkkeqR1QalfZo6vmxkJAzODu
d5vcWuOMQS4qKDo/N0mYU0prW+aoRTAS2vbcVm4lhqK1VDcRJ6O9CMFERokMRLsaxX9RlIO9Xqwe
fkJlqgeZwFti5E03X9okwvc83rj321kdETYCmnCE8eQZ+WFfg6+WzMLNBWa/C91vgOv8gQod7VsI
CLj0zxids1l6lDh5Res69xz+B96dxZ6wclWO7mX+a/ZIyqaDF8gpBFYmCHoJDrGk+I6ixykRIJUt
aftwP0rW5vxvYwp2oXAa8ll0p9nK/Ad1oWbNPNY1e5T85uJus2m9seil2/qTuD37DoA0Kpm/gvZH
UIIbidq4WVBV1YVz/ztEXDCxqH1i/fDaB6sNyJeuDJHN+NHD9dJ9PWR+ieFfqLu3pbKQoeQ1ePqn
XklrXIJmRIfPXTIU0NrZYLGjJ1mAx+oTb6JQzIZ3LfFM3EQLSr+QFc5VW/jI
`protect end_protected
