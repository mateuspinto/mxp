`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
lGj95Z9ffAXMjL5rmj/kzxISUysxbXFvDljkTxMzhg82zeGVq07q+DeYwFryn+FWWl8hftRpUdQq
GaV9GxO0NB07Q3Cv4EmltxtD9vwWum4eahdTgiCk103pBqjICSBZk/nssT9WFlBrxabEYt/poFdD
AdjEei2Bm6otbURR0646nvLlB/3J4HHNM2ksfW096sDSQAdZOQuYV+H73fohwKhVM1NRAUK3dFBP
aTL1D49j5OE6uiu77aMWtlJm1RbT8n6YBxk6vxVUcwK95GqTXVlqllpRCsE3RPZdipcYUY9wfx+j
RylkY3RifyWDcXc/umT9SF4ymj42hnD9qb9nEA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="cpaZpUTg4KpZ/jR8MpzMT8E9UYEh8D09j+o+J3/yYIQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18384)
`protect data_block
LOIPCA1cZO+ugYwudD0TDPWUvdssB2PnIbuTLgi5UGf4YrIJ8GUGMYpqGFBFwtkyQ77U19mTff7z
jKPdJ3UfXT95cb9QkkfD88cv73MEXZIHRjJ0P4x9t5jt5KS/Fv0OeOOH5COUZgrFCu4YHrDSYNbO
EKGgWAj7ft1vE4Gdppz8lknvJoMq4absd3i4VSIcPeMh8Aanb6ZqXnT4Xo7shJ4orkeTsMqMTt5b
RB/3fYJfwfhwnxdr110TGIdDXRz+DDwM7Eb6T0Q6Ew0wgafpCkw1iSCqdeKFAmy6kYNoQzL5Pqdv
b6pHn1gm4YaB1SO+kymi8Aiz8uUK0fAB0ck6/NzoxosjxgKq2WLD/ZvWAXOdldGEoLCJkPI+bRBb
G0LJKhooHUTAQqjDMQWoltez8Lq/kd5zV2ZNNWv45VQg06b9Ci+kwGFq+M2Sts8QrmYIIYx6HeRG
x7FAVbd7zo1nXGIYbUGvKmapI1CTZuDFdE/mDxztYIuLHgiW7ECbh4KeqqLFp4us1M2b/dnnlahg
jaOQ7FEZkdF/2r2UojIlxih1+aKF/mUn0VNWSMM6aoMDUP+j5o2mRzKlyaYCJYHkazsQzXdIDuGV
IFEZqxUbwThwkGUCEbYc/Yuo0ELo+VkmZxjaIrsFNga5SypkGQEMFy7FQmamevGNnurmHEokFXut
HATqIbvtz8MMVIo+EaAB5Lo2mDCzItw+WoYvzcbGbjDYVQJOLdEMrPrF1DM7y2KKAubCMh3I4S2v
ymf/sR8Ek8UxFpoVrUmFwf32b5M8FPWpthESfpxpL/mQiwnyzOWA48w3qFiekGzLIHwxJS5+31s5
c7oNKVPP78BtEdM5v3rlburnwWTzaLou2bDYGGrW+kaz6Npm+D1RWBB07BJBO6Uh9H80ebDSbk/o
b9HcugJ2R7J+GNABryG2H3JfzddkuimKaCRsJcF2UfbsB6/7H8B9VtfiNd0yZO5t1Hgjn3jQm9Zr
vKE+VZk0yQciLTFBgvFqin9CpevY1vCePUGWBPwOpXB/SPexJcQxJtscIP4VW3mZs6KZhyERmKRS
xh+PLy0K4RDt95LPIkZ8hzfrOpPB5s74HELDm/2llRJcC7CvowDxIzY017Egrn2ScMxbcIZQiheM
Zm4GjBZcoznCKXT/weo10Z2ej7DkqXw/lNwRLzgarzN/g2tnm8OyMHMAP77f0Bri1WmiOyRzJouR
ihUABdS/xrAS5gnSZHxsUjw1kef1I4kcwiTKZxC4XipjysXIevgDt84tsLTj7Cf4u35ZOaKtEdKI
rC/li+ZWSnLcVucR9X84slYih0qfFtV7YcPCUkH18CDTgzZhmDKyJdCsd7TGz/v1RWXILt5PSmln
yaE8fK1hlwtRsnXzMGoNHwWlo9i2GazKDKVOENckeP11Zrul0xVD9rKMSOych0xmoDFfGDAdGBCU
uqoaO8JsH35pIItNHqMkEfdmxVFioARAAcwfZHExUgdce8g8q5NUkncZmlBNTbEJ+2OCLLJxFQL7
sBeIafaxyLU0zpCzELQwO1ajSwXVDX4/fCC26moE/b+qFPX7/siRwa957rjMnyqlZCTVHEZVIqkW
o2DXS20Dskg0WrcSoC6ZqZpcg11pVnD/FO47pxpU1/OUS1JoiO8MFHVDtaxpxp/tvk/qEMGxcCwn
1Hf8maGgin97E6+swTtzehiZGTSdFNivVRMpwts9bcLQLOKfzYz2MPueGx9+WguVNAId9BbhaYyr
LJWrgTXqZhGNVIiUFuFfU9VLEfnp873hHfVqHvhocWCDD8CA9VojBIucpHZLAuT1drZPjaPgLTVO
s07Tta5v59ykdpGZ9N3FGmprxmtfv9lpyZqBW/r5GDlHbMxw512HGqGgzW/dTtqsItsZlsH+4oXS
PTJkcFhElbIeKo23zsjBjiX7LZLema1GSPQrW5SdEN9qrD8WI0TJPigXpZ5+WkAIzWhe7Q3j58rH
EuCM5JJKBTRuDZTmqBIg8aE87Gvrl6qp0lUFjoFFhfTrtKyMVr7g26IVFz70e9VG3RPnEI7Nse7p
23pVHgWRESSeO9BKeeZC2BcWs3u/ngL5fk3VfBC8WQJnZLkGznGFcXlb1LhMC3lXQCnmpO7ciHrP
nb0uNIMhi9MVqaYI/kIMOM6xFBAw3Mm6JUhf6VU4spMS7VMaeKsVueQXJsw3ETChZYBaApzgrfqO
yJBg3fvYV1EUuAqwRQpndSSfzggxDeUOhpID3aJKXTXre7OKQKNd7DOOqe9W1UOo0z2DukM26b3l
ED0Y8IOgLhFnnTFDk0eUO/VLMYTU0sgK/DF6I9+gjoqW6RcRykOQ5TgM5Gx+5bPceHCjHeJU6Hu6
aSxcr0pHk8xqN5o1Dc2gthRJZPP8+r6TJB5mstwIhopk8EeIHjjKyXGys/BD4u/EwzU8UvxYM0TY
AKj6lpBTSVO8nmQ/UWSQyadRoJkyQtGIzXgzLvaqCeN2SZ+Xfd8OooZX22NRQVZtyayFs19UN+HU
FICl3dJkJFcLXFyAJFekAGvzDdroV1eLgoMHK2RFq4pWtU8z3j9gNlfrAhjGDjMCMeEjLuoWs32+
EjYbkdlxGa+JPa6Yv5VceJsupDQneAuZRg5KkLEPKX9LBRhfVTrrB5dX/aDPr3SwK4ZsUE09fm5X
HdmcaPRTrLPtp9iPQ/3i6yhpFnZdRw+q4yO8wynP2fisYnwrbmkoisxDFIGPPG0PyTi+fnbzxu51
+xE8ugivKSwtebGUkMT4NiwLV2lc9Yz2zOIeiA2DUZ9hDoL7CBX/ZPKe64RhMpGLTACUTelTryoE
/waFSYDag8HbrMFxdc9HBWIMET1UH6t2NQL5Fig190k4NLF2gYhQt/yKo98MAJQfkfkXkedox8uP
veHVjhKZqrqf0HqGaE3k8AvUgRkkxQy2kIezV3cnmFjYmqsor2mknwSGEnttFGdXkhJj52TmbEuE
sWHQFNm9tQz6yEDRZ4DZdzWQlMrVWJYxBjEyrONpV4sMkDt4Ko+kRjHXMPQKK3AKv61Vl6M2kBTj
9evoXw04Ka3At574L4xSJozMHMRvEjBf1wcrgU0wOVIilMbC8icysMVWsdcBH4ymw3NrSHs7/X4u
xkTmq/M83rEkvNuTLcQA0Yy+j+5QFmyVcuXj2iN5S5TvAMt+SH3/FPV1OwH8CiHqfSSB0XwBylza
6jDyqGYxkl5HJVuKhJy3Jvn9Dz/RFX52E0yXEPsPt0usra97HWgOKQNVqMTOaKUapcvDHEWMAsL6
ldFBk3BgrH7E19zKCy4l8ZQuKkNSgSQQBXE0T2xiuWdzBTE8ZImDHk8FlMC0kcISP1HEyV9L4MVJ
OxywScP+GHJmzXHtx4xV5MWW58mBD6zWiS5+M4F2fUF2YDsx+0DsY8bF/n+sHDYClwU5ukQVuGnQ
XCQBEJv1wYaKZRNGWiB00YoKy3JPWRaro9YotkO0ailQZY4r+YvU2Z4vV8cqfPBSgNE8nsKUTbFp
vH7VCkmPYPxDs+i2A2hYfu8I2r0MV2577xU8iZwBc2vtM/IzKEV9n21mHgBm2/S42h4BkcpJBXh4
SUbzTh95BALdZL/lHQn7sFXF2Q4k4VCncjIxxvWGAPvtIojnZ2Hy7vK3E+rD+s3BIsvy8vxGtA8T
5ySnvFHtlDfFjP4nioGIjtz4QpP4oS1z3kHiVXbpzyQJ/Uzh+2JRnqErQXHjAZml5ZLVdjRH8Wym
XHtEK+P5CPbtbrHjKPGlIUDo+2gHp/yysMvJr5kFSyVyUGErk9SQHKRfdrX3X5Sk9PjD5lHspjwH
/WYhk20+41GUhsIUXYsm85iAw987amxBCaZm8U/rKx0DkscNBuMbjYsUUfXTSQrYxJnOuvPpwvQI
vn8b+R2n9JhxLNV8/7CwCbWi1Pn7ML9DJoxV/402MldqD0R+bPapv7GflD6YKwD7D5158/Ruyo/6
FKF5ddBuF3B5of1UW3NzmSUKGZrd8rCTm9Dx4iv7K5v1k2K5nEBKX9pmYdL0x7sh6xmTcj4CEH7V
rmHRtW/vXz8gvoeO3oF2Wma2dTn6KNzpgrrRJdoQa7raNK5SKpdYuSQDNGp7AITBteQP9LNBrpGW
pjAAZqMWKq+jcAc7i3dhYYf7x9mUXXVS09VN694jd4zn1vahlTDrgKcLsrAThCDcBCmpTgavL7sb
YE9IkVVYhDzJnjB42Fn7lARS0vcoFhwYeHx22cPAJfdjzrQB3iIVPYooiMmjq/gaCgN6TZHomYaz
0B3uRtZp+YjoQ8PElKRLrT3GZDLE218deVnXdCv94TnNzdeq/gXSUr0BJG5VRqjrmGXXxqrYQvxF
HLKTaS1gjTaMLnz7da/fj9QHoFulw3cpwnIALfbpT08ESeCu+pcWj7aWblU//+5g3gD37Id9v0LT
rAzP/qwTRUl3oZSu7vuHUQ+UW4OkZ58Olh9auq2/GL4B6Bpwz+8tcfRe98IGVOEKSvqEWDT9h1uP
vhLaf/B/vGMMQIdkHhNZcmxF11bekWim+YB3GRkRTk15XFjJIRelL2rLuGC/I1DLptolbgWC3A/G
ydokzRFXTKx1fgGehjEeTB5pDtbQ/XFlaCuelbERUvo4pEn8G5nDD0I4o5o9P0fIT2vcw0FTGpFZ
q0FqxkdVAed53cvM2TdTyneP8EBCJIF/qPwhQrfkW3y/ZLf9TTKFyPQ4J3QNQvIM/8PZrUUK4dje
NopLrsrc8PnIA3okOocSucgkg+2/IOUqw4Ce3tXgNk+ILx48keuM52HZLKTIvZOGg9tgnDA3n0P5
d9trXkw/XEnKYp8FGT9cMT8hlYLlfPIXMSOBBuL9W+9Us5i6QOih/TyZkoWm7q8TMIb1YlgBLHm3
6iB0eWCd6j52jiE0KDPPrQZD41RfwSkrmxK1sh3CKFq9uTSY7mQj1aViLx7oVvRxvId62PjTElrN
KKVMTszOW1+fJjwwZNYDwKWSYlTQoBT3OZO99hkCt9d3iQ/6zJvykPOj1Zf/WmUENSx6//edOJmm
G4A/uVZruRXjKO0HsEUPHttNlyuYGuvY1rXKpRqYmgoCKxdm+UuRGqSdAJ7Cw73t3mEjR46bOetg
lDZxW3U0sUfbVy7/bKQ3mQDqBBh3bdvxVXhFymiHGHoqtSBxnGCjrRQdkjWvlbdz+9ZUSALos/Ig
Q8J7qNIPpQjbgDrhIs5VlTwZYyT8UKDxY6g9CxDCge/SA49bPJSGTmCatlEErwK1vUToMnCZlZnA
1n8RJmtg2HmizkoYTQQ5ZdeNdlLWNLZaKJb3bLdzHijWAFyeMv/TcjXr0c3QVGbTtpjhrpocxDdM
fwkn9hRWBRlcllKDCU5ZfUDHfv13Pb92nXkAgMiDqr1B1UoKv49kXFk09wQvO1meQ2IqKVH/fIcg
UY/Ae/fe2Tb5+TzK3u+AvYvFaxU+s3vvuk8kqGmmz6ZSeYWqAu4l8OjT4pbsI5Q1eBJOXvdCRYkF
TOAUSJ8ozC8i8hFabtIZhKlbTH6T1ZmHXJg29geWdmDSkPzjvosdvBWypUNKf1oVCSr13Ri1Yiio
GLPH8w4Iv3drySpCjtLLvkf6b0gb7fJRkm2LWQIRSQypjFyPxxhw26SUSjc5OsAp70GWW+9JrBya
cOs9wPIEvNLALJua5TUzjIITpLmBSJ6gCnEgCQf+mVToQmii6EeILn/+6NFDSO2WKto2NlHXpuSD
88pvhzf/B2PrK5q4mX8vClMz16pzhHdOir7DyT+HvvK67+D5450DHzXhUwObNrN+mMe2vxsQ4X0/
sDshf/PT35RsgwSTvsTGB4/Glp+mEOiQovyKvlgtj99ZRrJvmbpw1hfZO52f5NKT2cKjkut8WIaK
lSjAABIXqzkO+hkmvZLO+KMnJOdJBHZ/HXL3NIhLm/mTvXrvNu2S22tYiLKwyJ/9nv6iXrzR2/P8
sNboRq8RW9yhFbdveAwbibwDdRVZ9y1qFDVGY2EdQgx5bzNdVxHqBg5rcePn3wACyPiBXdJScp3A
fYZdxEPv2MK+WZSchGy0V2eBXDIWqd75QGYuGe5u5ZlQBcRM3VylQaAi5pBavYqeOInf3y9HoNd1
E+XhcZxxyDXBXjsacR3zuPpkHmx1+t4vJWFZWofATuBzAlWLAjSkTUIq2ACHE3ZrlNEgYR4VEt0k
ssCV16/L6XWxhuKPezboSaCFf4nnpmoUPC8wLuzdCZ0x/BH0oSk8YaT53Cz7QJTVwPfgRgUj63mb
K0/4tkEUOtrlT/h2PCjNsjO6IUSB3jv7DKle2tRn9gsOnmbDNCqXGqZs1qC6dH7NiSahgEXI8WrM
EThgXWqw64QCEVC8AyK0yflXFodDinVPG4ZYU1iEjPz8IuWqsZ3RhIubY7NUiwK3NwC4nqAkiANe
tCCJR9+DwwtjIlhv1G1ucs/LTCcqi6QAzQALXYqNsoFMmvN75nrlhapUZGVe/ytn0SQn1z8KpKkK
+VyK37bspcClgRL+1KQ9/QFWcFrIQuupEek0IM4QWWu1u3YLeStMrv8onWoGzpEyfK85Aa3amdAt
eq+Yq/q6cv7AuI/P7GWXtgiZyKkv73pNc/lTcbSlUQ99ttSSOzC+V4Jy5dLsSdqkqqC714cSR54Z
o+6e1ryPnlg49Or1RECor1TfNBcQRu7Ice58cJa9Uz7hpdAAWGuyvmOFSCl6+fUwuTeaZVbMnVyb
UBA8lGWjLiK7oTX+OCCKmh2YR/KLAmemliYGywIaX7sqJTIjr26zOjAINF65DicSLm+7lq6I9tXo
THtEezSKbNzrIip6Kb7tm5dCTi111cCNK5bmHKhue4yr/Pi5Jd4Zevpsc8umolur82NpDP0LItI+
eeI5c//V/phfb0Z+8QaWx23AW+883owzYuuI22ciMq84/OSKbNRLyyebG4lNrNw3xNUMaJF7dSKB
527MQt3XT6GkAPuJDjnpRttdqmJjTRD79YlkxwJHo1qYFM5kh/UG9Zn/1YGjMisAY0AD5vVWLU/C
cGFVA4VBaa6USMbamnGLwUr4SKanW7mGKi5oWVshUY5UOgk2HR3tPMAgTlIE/oykJI4zHWtOa+KV
rr+IrZxMy891H9BSyibwT6VJyGw7Nxb/rdBZM8DJNpMUhebtZsfCZTsOy0wEkOmFe/TZQhjJLTwO
ng5W3NEDoLVCIaB+eWV0QT3kJ9n1SXukIUOq2AlL34x7IDg/3Yvrtr/1eRaYHirkzPlR3PgfoCcC
Tmsh3Nw/E0fgvEPoW+3AccOiCvJtEc4Rt1N1BcS0Uryj2CBE5u0zadmVC8Qdo3tFLlz5OqTwch+V
5dWQeVYIegNBqNo9CaU8PQUP+bcPAjVkWE5nBRruXd1wcBMq+8ORIIUVG4h5CNQ7OgKGKv1r4Kg3
QljXH+O5ZKh5n5g5pfLP3I5+4+yB6dqJcwViB7PlFZHRYOAqBM86Sb3ZxNLWIntjX8pkbtTxiNOi
Y2eZpCPRy8w5fVH83dk/IcIZ0Hkeiqc6qcK9WVBvdN7bq2dDZcfvAB5KFUTy5RrrONsgFNVxjBg6
HXDnttC3wWyiAKZzQUd+Qm9ccAHeVTTfjC01LmWWwvY2zM7sU1QYY6ybO9R7ySlbaYlKzlGjI6PT
m1OA02hY+2EWH1OXnUCAugRPZX3NqE7sJftexXg412R+6a6pkl2HpwIaY0VkYv0oVEqBAGF5EJEK
LH3NMsOUwxBLyRoI2cNbWW9yhWXwV/9EN7g2wdxZqjCcHRGMqixuIPK+cdDKm3ofmERvUG/gscyQ
uPtUR30hG+N1YU3NdJZbPD/fVzNmS1LrL/yrYgiO80iMF5MmzAGlo9KUyN9i15OcttvVbNMzj+re
vy2B/CGHAhoLBcQuKYhsD8zMOla04FTweN1aJuECPw8HsXAL2EmC0Ibt6crdRTYpCghur04C1FA0
oA+1hzDFKF2PWb9CPLFfHRQt9Df2gL678wOUZVxOzl7NKvrOWA6shXnr453I23S3zSbg/XkDLPKm
LjRVra09f6GSUkdCdoBraF2X4iTCvAjRiJYLOoZjvouvBadOuSo1/7GTZHsAy6c4V2a32A+tcbCN
E5i/dXXbBsIp1T1nXEegnPdmSvUukYQqFvLlI0Yr6T0FwlzM7snsB+jvGrLtr1gQGaMpG34A319n
hLxw2zOu2ifYHZSSvWBh6WOhLoTTIq99BXNH0jrzV9cAmpokf3WpSCMZ7t7WbLu6K8GBbKCyzGyA
/2bkYjah7MMaOgNI+2bvS2fEhQcJoxqxIscb+6UAeJsw6CzqYT7TUwBd/Ls+usrLjYkpCBUFe1LN
gbdMflewn/yv+8tcRXsmL6XY18IflqBj8FpKH0cwL/RmmdNLkH1takUKpt6D590Px5X00HjH/25N
1fnrbsCDcKHwVK73PxG16cd3v3Ao00+neVSv68y+0Mk+o6qb2M66p9hvjwwRZiBJsju5IERUz8vM
ij7oJIBmwNPZzXSEU8v7+fXTAz4EM/EtPB5VfTodWk9vhD9Ix58FAYmZzHC8oXNsaPLWVMeHyNn0
RLgg+zehmBAYzDvO1K10lD4bAUF3G8G03KzmLe9SxEicSGJjPnBNK5HOe9eqVlgVyWLU2lyVojqD
UF1qbAhpTZev78xxRwyfIkXxiscfPy9pItaSFwSIUuZtTjvRnju+gh4HEffsEILrQj+5DGgA763g
Xxm2nF7GLEsy61smOxXP0z83lQrIkkxlXpz4FAJeQtqEt1sF3hDKzqOgqqGXM806rS3m87kxbweq
ARTIK/tqU4hlPqspPOi1LkUzcU7wkXpU63LEfHcT99xx2zGaYlK97EnLRZFioziWDPdYq/hn+duq
TC9eJmTJgXVxhCK4ohc0ONLat+8nCGt4V4mRru60VcgisQyyPpHMORNCfknE04ImAcWUF+z4rZ9L
AmkQtYGdRW8sDXA+PedWdbE+DDem3jwseDqVMyTyCMSPGJInacBhPJd4S32hOPDm9wuvUB19/6fq
mq2uwDaqnyyYR4NFQSGcSlAF0aCnF2moXplU16qjkyMoKTQqwjQIFVO5sjcaCMF/w+fpZ+p4IigF
UXmCPnyjjclOPFRM4u0T+V7+aCPvz+OSBa2/r4+VuRtnetTFbUrr4VY8DqXf9nk3eagcdoms+FaY
NundMiIYeH9rSoqs0IjJkSVCnsePa0RB66V+kyAaUXibO843iCZM6eOLGrkzA3lOZYwB2+bXWfmB
ErHrWrb6Mg/TOardRX30mEYQEquAj+Scz/ER4v3s78Y2QQJ9ZF1Lk1iEFOl5+9VgyoO7frjGzAJ1
J6IIIOm9ST2qAnDTVqjGCfGoMeo6qpIC6fPgYMbMNDYcJ08h7EsqamexXzSwi1FayfR9yiUubRZt
EWbgkYplwfD0BWdsnwn8QVBvUPWoUn4QaL5sm1aa3Bu6JOYfkCThwF4hyIWYCruhCsrfnXBtiuyf
5X06PKTndfqnn20gM7lAO2zAs5o3H3MeRJ/V4QDtI84Cuau73yO94nKf5aJuje7xmKudoNbbNT0/
kZIklLtIzQtwH33HIyoDQlrgNMpa952rP7lkF28UBnkjwsc5pZIeeWOmqVbX2Zujab8bC0KQTFrO
DiWRs5uSqEUIce0gv2tng+0GfKWdqErShbKsDu6HeszBQt1iI8t3BLiP8/QgEe5UtGvWOaNrmwsW
KpovRXYkpKuYH1h6nN8vcKsi6GMsRdVi2geRib5JADpMLb7MMATQpb0BUFGF7DHlWEdmwpdNrLeM
9Vi3/6yc7L9L2D36XfxXStzuYYBBg8J3q4z0MaB9UkyPFN5o3jqKeKBclUHgjdiSCM/59519Lfzv
nLC6j5R7fEkowQ0lxfOTpSxr29SDbK6peqyDWXi04TZ3XAs+b0HqCp+nLXbPfbbrSZ1zGOPT5k9G
8SP4DtSsdfT5at5XHUnwuxxWiv249vYJJgbmX9rCFZ0kTI4X34Zlod99uu41ZB1NWw8BmHtAIjfQ
O01gu3MprcpgcBgGL0AM+l20uOcekhxRsnyWnEa6MXzFiQHmuvqczkoRWar8+TBd+I1zfin3D477
9MY9auGreFVxLfsZR0ri30WFbI8VFWWUDEfBuk9Bz3lHVbX9+G/1eyr5Q7sXsIcKa02TAljJVrOd
fD/4efwCnbFsNdhFfkDJTIVI/YL8GC+9eDt4AKUevPJ3hCnZLLizE/oA27UV3fCDl1h5508JpyKl
b7y/dGFGDlKUtBbMyv77EMnhrMED+aPyHqd+p1QwIsRnAHH1Ng+a+tAaccDHZAAoQ41Orc0Uzect
NrVdSBBZR187RVeoPiJNJQqcYElY4C/EjpBKPiT+CHMO2zFLATHGvFiTfuCk9MiFS2pFKvMHvALK
eyYxeCxrWwM+eJHtBPYccjUu9z7xStU65jSXO/O9eKdUMnAxJEa87Xj91yNM98I4iYpUQl9j6xHX
V6k7c4UyhLzV/7USiIwMhSD6GL4If0ZgTgk3jvbzqSwOwg8U00HKqKLiRYxvb1XnWbR6M7cBTXUl
BUikBPxdkuV20wDARMOrJ2WeZq+O7B+PlWETDzPVAJIMR9BcxZVLNCftJ8Ox+H6fdGDltBYHdv2h
AwPRWn0bNipdeXA1BI//+MA9wdmPqdOeW45r9AugEhie/OeuKH04scA+mKESYnH+TgP94F/Y3Bb+
sG2HFmMMeFvXJomuIqKN2ppl2j+RBzF6k9b757V+h3rLZS6K4I93TsnYkWQlJOmQnVJpjgN550uj
8G8qNbGqGOs+XHUXhJYlxdAqpwSyXyFgkfi0ylquIW8Gwy6dgVytyfGAfHE0/9wExAL1V9xLYthc
bUQ+s6HZK1+QD3IXh0hJUFyB8G7iIljAqhjcRhbNFyUtqP8aOAQpyy/e+/u7LXwa5x04Xx33x6j+
nNHNmvkeMYFmE9dNJoi/W95c3k2BkV7FiR6dLa/+KK6HFVuGWIUzZquEQp9f/dFffhqQ2YFhtNK6
zgDvfyp4B2BkUBRecMCipMzChYFLYRDGC/Oi2YR5H+hvMbE9S4myFeMLUeJm5g45vfT/f3tNmfP7
oq5j5w3TzE6lgqceE84q6LIh3Fc0Il2r0bfowPhMjtYl6YHQzbsJyWev10Do6GB46t8Qx/XFvxRz
TT1EHww7653+BcaDoDwnfSMmKS9CKdqFSoSvpp/8kN6ZnI2pUfnFqNFTgXdYoDcvIeCN9tHKyBa2
4Dwwz1/6lX9tjLINP17ObDtrXQH7cD9/ZrOJ7VKpYI7LpDiIehVSyZaQzrRzCRppSi0S/xR+MpRp
yZwz5rhYvAy+zmj43I6MeStuulCD4EMDhX4DTzApOkHCxlszGxCtnifo9NlcsABfwlwjENita+Vl
qe6SHC1uaviP+kPa93dN4nVNM+R70VQyBHNHKJ7kLF8C7lgTJaZ/zd4eFTp51FTi4nBeaGy2QrZR
C4JMgPTHN2ZHbHogM1xbHF0mEVTejkhrlCr5vXgbVA5+zFLuOj/Z6UWPtca7CbSdJPsdBprdurkO
9iX+5nrUTWfptEo1yVyzzPWarN+Cdafx2675PLTpmmF7OX3rLbNLiY9C/IJPXKX4s7GfrRLKKOGH
eqlRO5bvS0zCtkLuYlFnLRb4gM5uMpDRe1t2UI+r0fstzdOVdDipEjHtk86PZx+MYFf31SAn4ZNZ
xORBH9sDg0DVNG3TAI8K+RCCT3bjBhdwawI57oQqKBYB884FkYr7LebqkDP/nZU89neA1IbDRZYn
NWEsEoKqHGLx6C2sV/KlNjCMe7J5xGrJPjhc9VZjZPKGKRxtJcS0Ixwd2VS43/CDD6/lUTKY2qKA
c/33FS23ZcCnxGjRGyUFAAE7UhqUIPz1BlyzQUhlLM8RTLt3bqj7FJYbmilzin1cRbcDdll9pJVK
UMzYno1PlywKdsYb62ZchJnoG+gloqLtezKOyWipuZY6y+nM38mCDNCnZtl/Y9KS2VtRHZ+hB5sg
HkenpyrWBqtgZa+mXy9poe2ATYuhzivVndl9bow7jwhzrQA3iZLaL3wWjZMsma35wgWbgO6X46Hw
SZaybCTLYCuBeKvYg/pATmwviBx+QZzE/o3c6oYcp7FHgR03dqhKfJBNoa+0TA/7wX5/SLeJ9jbV
ukcH+D134MMRiND4SRzuhhR71j/2c5zo7YIvY9mdRLG4Y51LwppLG7ajl480MpmU6sSTch+hFts6
UBIPhzLAPOIOYHV90owNvnvGV7snbCwsSoAgzaRkwEXFVLHtQtqWi8V7JawhDZVRyl9BU+qTF2Yz
9foRWkTPzZJeLh8G9v930T62U1qMGqyPSGsnCvtbdexmT+Wz2wxtfUTyk/AHYJqT+HuyCCGn5NET
bWiJy2ATQCSr/z0Pg7BQrEPQxz7AzWgoTh5moBEvvQWuC5KMY6oFMtNlwn+iAhspsvtbGVFIYE3V
P6Qs3mZCW4eizIShyF0J68pGU+Lwbhc/SRhOdg4TquB9Nilx+/1uKXlBPuBuMLHSnzRxdMCrSTZy
bNB+WkzELF7TU/ouYguil9+lHiiVscdcE5UOR2CPZ3+zVK3t1vbsUAVevxWwxyU+EqIFeOOoH+am
6DVTBldaUKCE7ToOXWWoXvDAY/90iy9Cs56HEu2SI+rWEeBaezqcOdazgfwFIjZ+qENiO39Bcs5M
K9ye8NGF5I1YU1x8HyvMQi8KZlGZVl2SIdBiAC6ugAqRgfhuwh1G+Ltaly5maXsQt9Awxff7m62K
ZEynMjJorYnM8n53QkkWYYhgKS4QV7i36TKJlttu4XP+5FK6TubVVoZhqfnHQbx2ar8WfG5H5meX
qF3RYfnj3kCyajf8FDtOlteT9l36/YhQYTjRLM4i+aqaZDRVQ5139BSoK+g773tSqC3/fTRFb5xO
kPph1L6c1EjBe9lIM/00sNtZrKk2xfntgiAAg/u7d0yPXouWzsHJ0IRwABPXIbmVJc19rACAhYk+
gJoJuIAjQNNTdYfEkJDpbe2cimYsIUhlxoRrFu2K2Cs8pck0Fv70wrrTZAEPeVSOL++Tg3ChY0yZ
Z4sRhoRcR7gXABzK5r/3FSjqp539qnWuNccENzBium0ERyD4V8WWIxHDCrlKJx6KTjjS/i9J5mGh
97K8p8AAQLulD4/qfPWMjBIq2yYuLXi7lDhyR6kEZhF1NCo3ruI/gy/Z8BdCq8UcngxPEtVjCMKH
CHw/dJiCRh8OxsBZ1UUl58q+aGDkY/EsBRoBMCFNAcSI8B/jhWDllW4XVz3ceIrxwJsJL8f3ytXu
AHX9P3KNhnib4ImBPkCmW/4PXpbQ2rAp8NtGAlH7bea+2Cv+KhxMxGXTFMVZlgkOQT2anOAgiBtq
8MFO23PuQRuttyYVWZ7pHiB752cabnVtih74vROgPSV8TSOO5KRIZqqtJwzhi6BIG/bxqZooyQ9b
Mb2Na8uqusdsVNdcBPh5/ak2lhAN5I6yO938K4NoL8QCt95kNu0hIvZ3n0tka+UmtcwkA+IC3m4K
xR5DlwgQpnXLC+V3/EgomAkFD0bnLM6fEvHAzmR/ZP/A/AN+FLVHykfpMFvbx6DnN3sMvoTB4c5D
mvD/jgQE9FZIXc1TbSMntTNuj16s5cNWCl0b94OVf6qn/Qy2hnC3YhB0Bztv6N5DeF4/Kv3taRs1
UPJp20MG3cXR9QFKGI3U5VhvrpKSn2Xksy+L4Y+8zW4Vz5R+DAWb4jnDcsG++6hPr8GnJjH2+CxB
xdGKSWW4QN3Ad0m/cdJ08hEQZaLq+RI86XPqf/pVEnG5pSqeQ+Lq/JaKUaXgcun1v7jWFLIlhIe5
USbUvF3E44bS445Uynri/ZdHLMkanLoHweIDIxKfQ7SAtlmDbB2+8gx8SEMbgnt3yYO/Jbx9CN9B
UnPvg6o7n1DqBouXDumh1S1riA181B36w/D6YVMOg37c1ic51Ek7zqujRoUZk/PpeIUyMKeSOA7H
8bW7lln+VUZ3y2nr2oPp4A3mhbg4PqFO/1nL+76/CF/Sxw+9G2EVGgz++VWltA90LT02mYc1Qgmo
dF+I1qWo2N+4i30SWHSrc+3dJJMhnq0UYJEX61kPwdiQs3Y8Vn9WnNqihiH8itTgQ+MuJ+o1dybF
wJEYurFUSbRTLkcCmxK4PWInYw0+KEYKpaqvAjV5m5wf3yq0AVoDZLb9AHzRMexVAeMPyPomaNRS
mgHkdVSSU3+Iex4p+c9y5zMbRxddFT0qR+SdqQjXj6v1mcQMMAhoWNGuCYE0auSd44Si21osLm8b
lS3Fp6KhqyR2a2pO7otKtRNMfyCiUhYzkOcY08mBoyXzNo/haFWs3JYtnVWxlD48rOEQRnXhw7WT
7YQwJMV15EYiBUmV/ulQkHprv+SNYwhgHNvVGmy6mwsZd8KU2DtzMYeWVExbJWWXh3d1AxHYAB7L
Ar7RzNFuLyQmVxXiRmJj5GbsStCMuEtn22iIq3G6iPZ7SGieYoIMKnMB+FI5q1f2qs63qMqRUIZV
PhahmMU32A8x0ew/Hdvd1EYuMGJBy6O5fV+ewDIf/hvMwziyqsu6vCdL/vzNneFHabx8XvCfmhBQ
pxjpkTtxZtlhV7G9NWwSwTlTtSyWkLxGA224I85jL7G8HepVrB14hJ55ovUePJnyFop5nFs2wZyx
Ly+xePgokh1DSCDKIc/G2FS//svLst6D0Xd9F02psaNZyeYM1I8NNNlbvEZAM91X5Vp/svoGYlid
O2oPAMDeIX7tYhZY25SM+9YhQw3ycmm9MVcbZzyaVCnsPpjf+4KPhiw5kjBGyZAD0dzPhC2LskwU
YvF+IV9gNwe4SjRalO0vIRp2blPQ0ql/AO8l7P5QzqRMlLSvMIwf8+R/D5qr6/wJ1YOWsA5Xl4xo
xHMk+D3yR9ZxXYRZwg1IiVtxkh1UYeaQGOZpTeUmSt0YuZI1Kp4Yf4KQmnLxuCrWsorxpzNA7zhx
x+WqLhyzW2q1yHZnGhw1WR8P1oTZXAeXyvU5jXTTLlnUgDfIbuUXia8AFNKkvog8M1bZ9sxZhRKm
jW8KGCBAliv58LRReoD3tLd6LAZs0QFsUMioRv8mFWhD7nCVes9C2g+hSordJiznuiJJWYAoim3I
o9wsLhQExTEaho4JyvEtv8BoU/eIcs1ls9Z/oGxNqnl6Rkt1Q9IeX2QUMV9pInN4+zjuZpcMGSle
8sLhMHskfIFUSjJzzD0Xxz4SwEmodks7aC52DiQHL9NQjpe9Mb0vPWsMOjQ2Jtz6ZPBbMVEuFCyX
odx5dpbbjB7Lrj0nkuTEJvKYfFBnkUF8vQwlr1i7x5AhTO9FSyOCoyyk+A6Tnj1uZBl1AunBpkHr
6GOZjNG6wgQKBNGV4TOgr8mTplJ9PWAgHOtn5NxPpMrJpxV7ElCFP//AubDSaIUlApiUctMM1s83
QTXvMVuTfaE7uY1BNpvAvF3guu+pRqA4Jt6xiZxfiynwBOE13w1wwr92nT9fDPycGJeKxLtFVpDW
+S0WY/v6FAEs6eYKJ6+vbiHXgnc7din2+LrbFb823tqO3Z3IF5DxacmScy8KlWuPtmUl90ZnAkXp
5uDtv+foPSuLlVYLCd04FaX4Krl4k7M043iIaYHw7p1i1snPyqYzUFzyfdw5BqmsPTQb2Ke7gA2U
MZZHMPt0GbvMfXenFnY2sKqhOm//ftP83Aubm8FaF9QG78+OJiDEnXUMXhRPygBtcK3hKYZuoa59
uqEQ9pG79wAlouMAfT3SlJwGHcOEqkgbL5HphJzIDe5wGdV2/AJQ9YtAN7g8oP2wequulJSNtqpp
+nbJWLfEzFBtOlRgD/R8opVQA1skASAk1YH54AVdO0TLLO+YnKXxovGZvSrm+vUJQh4sAY+sxRIy
R9LFy0XVyySlZnzKKA9+gPhrscUTHQ5Y8uks2zEXXetX4a6Q1/lOThUTfeM2ZRRWKoGbsDYfCMoI
U783dxkZqyDTT6HkdtLYCDjCM54dnafs9wbl64/kpIYQYQtb6VpehUV8UAcBgJ0Eb8KrfDhd+jnv
iIjBiLtQJLg840tKagvtTrhz4O8LW/H+b1qyt/GAxMV0bKmAV+pHZeIkRLhjAHzR//zP+wGdFrk2
Mw0GwmQoD8h5BPRvJS8pUgDwzuCiOWKwRQmoW6AtVKmx1lWwvLboYlASxq1dQBNL0uNNhtXTU+eX
V/x86jaPmy2CEVJfqCNcGo4TSrdeV+gCY1KnlbKVEBKnk3Dgxbp0JVTdyaTwi8VsbuYjoKjpa6LG
4A7hkEE8nhCwjrVDoE4gw27EV+tSNM9RC1kbzh5MIxjhy/So5s9G61jb83cGW1OVkl3/Dmp1znc6
ncupjY742kRK20n1M7v3ogo2pnTLBlkPxBrXULjw+IdlwOYd1bNSvrNUXglDI3BDvz0ygkeVKnjV
0zAiUVxqiKLYZRyGkvnAYecnN6pzy1pCLfycJn8zs8Xyvqq/en7+zg3VZNGM/q24viIifCVfWAgn
3H+FHmJCulnVw7qx0yxrJBR0PSjN7MXiJNUJBrkE29wNTeBxFq7sKH5VS8zXgNjR5OMI13enV8oG
HIuCM2HOOJE0kq280Td96iqGYTAxPqF+bOINsfxX8XcBs5Mv1tMDtfOT+QaKKOWD96gXWM+p3QRE
4hmTP+VEJw79g/w7vG0yEEyuP3v3ShBti+FVZJp7qkA5Af3KfXVHB4a5QN9/JnspgfTCCm0sv/mi
D93dvCsTIbyQH0Q+BBAZ5Zch6lbOwHS1XkfVO+0sm5MSOrrXq/VCaOObVmgKJjZ2E1Xl4Sx/ztaT
7M7V2LzP2oxYpyKasvlyBu0dtEUaEA6ejMcrESgMn88qeQKqO+HLr4yZ22Bz6sDVMCeMKj7PrWwW
a2JGdx9q6O0aZNyEaEAiRX8euv/A0mrdqBFyH8tvhPHJ+rC7/UzDRmVBe3cNn+QTCJnmRv4AJGWM
3ijAkri4CRrn2ke7zcUSXscBkN8IO2sY5f/BE2nRJVYpyCpUa/b1g4IDl/GLNEWEWBtLCRIqCzer
La5l6k3hBGeDJ0CXHHM1QMbN4S7YSezub3h25II5bxJ4V3gSnGeitgH/lxTxsuB81OocKONUKlVk
wR2spcwfsunTDJTUTO8OF9v2ElQjAUi3pArWZeLWbw3a3mlF+IXXDvwUfShj0ZixrP5hApIk1ndT
9Lgt7jRlxJ/EBf1h5Ju9E+f4YBtmMHcxLcobmU1Z2k5nvnoc7h6SaNIa6ySZ9hCD1qhQRvEUSkOP
iG9mRBvyKhMGp/H1VkDhmdDqxZSQLXKHiua2RomtZmGcmWhdX6j59lK900yccg6xKgTNwVGe7DGd
FFuxoXHcy0xm5JPrD/4J6ThwRbqlrqjF9u61uCovNW/kZBBwxh04vy6m9I5ZUigWE6h4mTNWI+yP
P0v1oiQn9QcoZLkRyyVeMWWT4fVy/GdSepSQOiY4m/Jh+HgC7YpKlBdmHBgGP9dqHkTfvmx4y0nZ
SVGFwtqV7+k/0wisWEcCEwhIHvcU0q/1KNQYwkkLae3ox7+hw11A7lsyW1JQEdJQExB5f/B9+nWO
9RTYjeN2Ht/5AokC68ewjtXmhM/lUZkf4BZQJeynjdgXhoCdUPXbQTBtBY9JMN6TIGkK9h8FY3PT
zAjp4jGzsvk/IWUDA6WsqMeY4B/rbMlb2BszzXumfz5yGbmTM8Lf0/qMUmLhw18WFgM3njByGDDq
rPIlARlO9dbSUPCBAuLBAHgXaRg7CppPgMGadr1cERCdU0pSxgOwKJBzyDh4AGAlxpARuHcyBpXS
k0F3rj9Nv41BN592x17/vvWexVZgdCMYIqI6cj2mnvUyPUvwAotwOh7yH1F58b5f2AjC8mBJv/Z0
Li3OBCv6pxyBv3mRO7zymIBkvHu/mk7IswH/sQaXN/p3XQFnZz/jnQ6bS8DRaMjQbsGlHSKriPkA
9AUSEzty7pa/WW+qoiLBbCBo0z0pBzPlEHnhuLJtWky4Xh+bHYZiy/G9ojEV4LgjI1bv/BfhYLSM
Te4Jlz0WjtRG0Gtd4oorXpuP8XC00GMvAAkJFzQ2dtWQqlbZJlaGcIQCMUYSBWGt2MMCl4hJ9+UU
RGSJhpU10xwtVV4A3XH9Dbm+pXuCU3cqVQ0Jg662ftkrMsXhgrPNByuzTQQS6BeqdfwchfkaFlmr
YbTgTwAg2QqbUrIe+WjD3zQqiwCCiz4VBWbAaLPojtgWFmHPFY8eVFCVW+XD8wIL3glZQzpOyd5d
b6tLGTnLnYbmpejnf+pGZDBTol9KNQHghHXklSnWHBTrYRMDZoU0O2WBj/31HbX3pwoT+IsbEmuI
+F9pSOtk2JPksh9vwe8XUmokjcXDW9k+iCr5yb25of2VzsCFeCC/bdtWFMDndIaBuyPLDmhePTvb
mDm7Vv/4o3UGFUsWqEV+FRY1jNhPS3DOVFaKFUmR8vtPCgNG9u3StZu+94CaTe9MfRK/AnQLBlwS
q/5IJWVz7lCb5SL6dKhMzPbp78dx22bOxNvNtpvx4ZajQB9GcA9mi5rInGkFMurg8X0UyDVNr8GT
hCOR3WOh+bSMuXOYGaHYh0uyGgtEirXzK/IiGWwUlT6qj3xu9P8e/UZLM8SRHwFDe5H6LC/6GANy
kMq4UNrgANcAcp/cap74HDmtl2T5HIKCbFqWdeOh61k6d7ARHaHseaiOrxdC1i/U8EG+NfaeYMXO
VD0J5BEDvdR/0P7BWKPBn0IwpKeXWRy88entjbqshMOtFXr/Jo/X96ge0j24xacWg/Q9PmUOgC6o
hrlosfI59/QmvjdruwoAyQVUiiVPbjT/Ww7hl9CQJc9W7MebH/7oXJ8yY+hPZG9ONKfyt/NDU0rQ
4xbL6OGduIpzVvTfp4POY43OUnvUL7ihWmVVuuG0LFIXbdbivD3cxbYtsmtlxMDwbPkVYl72x++y
8khhWn31NW2eay3lXsmao0boyx7kzWcM3LvBQvMsMGR0JZ2VkQUL7cQPzq9vP45AnSm6Fvr6+IBC
oizVuPgKBRQdGjmtaIcqvN/1B1DNglGbRuYuH1MDuMaKBLA1gTEKBg8Q2yFTVMYSCZ8a7aRtP5Fp
Uy5Jv3zUmSJ2Y2fyFYqf5kJVWXr/npIeV4IO44xmvEpYINJpH3R+pQdbSLFhZL+GIBzALBSN/Vl2
PR2eFaVAzhmH0G3wS745ohszCq91GzGGhqCH93hzDlXkwJgNJVvQpvdZmA7V/rv6Mv5ggjGld7If
7jU9XXp2D2AO7FKUWSrGnVHiDCrdF7Chn5MVeNaKEX/SlDTQD1zaYF8UlEy9cwIGDm5gFWE8m8ew
eJ6ZxkaN3rPd/9+/XJWXzfmVq/a5Baay8ftJUfwiNU/6s+6sSZk+mvKGx74z5qgGNGAfs2UfBrpC
PuvN4JVvJsySSZkVXqAl9vgrS+QBlNF8EswmHeO5DSTSdUFlc90zb8Covs3SBH5fvSXAeiDLl6KR
aiDQKcFiiToqCSg9MGt5mGLtcE+bHPtG5L9KIHm4hTbtm3dGZ6zTl7FKdt04xEuLzeyi/hxhdj0J
HJ6mBSxdG88LueKR9F0f6xz6VypsITsVfSU6VAyQ+HIBH4k9d4Lon+o6kePFyTCw/0/KVfxGuRVu
HictgVziHpnvDOtloK8z282zAreCI/exU2kxP1wf5exxw33jd2/PqAQuZXjibpglmV98Gi10uaBH
GOjiiM0Q32TG8O/kgk3lHqkXczv5U/w72cKte8DO7OVZzmdcEGe419ywiyexO5KnZTCtfLR3rv8r
duoXdy1vbK/sFfMQEU3IWxoKBHW3kJzVJbR3ZtH2IBeXe0mT99gnwbaltx4iReT276sntC5kwPFy
uVFVQucyyA6xA/34O6eSFgEvuHB9Izo0FrFcQLjCHPPGc1CQHuKaW7B7ErhSqxUI9IgNuKBo4cpP
IRSVooVOHk9r+oukGRRHnllEk0jyWsM8tCv6QoDxVuYBuZFA28BaO7ZM+jbZsdvJhF2wFnBynoet
BJfytP4ZnRD5QbJjdV04J/viVtZFdZT9ow3El1pR30NzZyGM+3rm7SYd3UOVaXACzxNi9v5l1kVr
qznjjBh0pWlPDhLC8KKf6S+DfW4yzJEW3istKvUTWdEPdBv2e4NoL7nfXxoj8UbNKdE+CWkH1Dx+
KtBot3DWOwmsxPtxwHh5+6BPIguq8rkmG19T5hEGglhh7a6RSRuWQ1S0M5BbHo6PYEfm4Ea2Zvdv
w5o4vU6N9aRQUmOw96SyeMflqcG2eWnU7/A0G57HuuSGqY2uunt/hU/8OH0hH9Q7u3Way9zH/3BS
WKQ1VY8eInF58GMzW1umbvdLVrEdK/9Up2HB8UWZIfNa2blwB/Qe2iXn8RGKR78um9S565ra7BAs
GEr1A0f/GgJJ5XhJTxbnZgJ6v7gxhNo9dfQbOEpQ1TjYyeR86TCpnpa0zsz1YbuZXLEfxrP9HAYo
RCvlGn1EbM4izfqvNPKFTT4jQD5QgfFwftqRJNfok2LPdjweboQ6TVt9VJH96SAFahDlksb86KMd
D/+edf7/VBY86RY+P6Oxfx82tHjz+5w0NwSMgTT7bgD0DxheFiAYplCVpMNpuq5OKX+p5RT1osjj
tdxsefUPJEqYd8YAyh3Rvgs3rlvStsmMv8IoUkyrLPrTGuJF5Bu9J4bpz1fMMHLebzSyXX6iAA9L
+f+bPrTKIra73tmC078x7SumHyHGubwrAJ9pNfeGJwOkiDWLSp60qF6kEM6xBfGxyGQObY83LaOm
Bf3k+0bsp08mo8VUsM4Ajhv2PANLUh7vNqy0Qe0Awje0e1R13pqfs31bNn2OJjqS7gqVF7HRrqRS
JY5Qb68mQBHELMIJhNKsJvwfx/vKefcyBfHM71lcoOUUpLY36HtC72/gibpwn2EiPYkz8TIZ7RBT
w/n0nsMA6/LbFgWJqTSW68oIFZmuf5se/uucpl8SGnQAZbxsObD22oiXtaNCemOVJ+Hs+fiLEUj8
7xbU6x1k0l3+rYXfVDXQwN9ZjGT4N0m9c1WrhGjY2cYO66nfIT09WhAnQX33NJtJt5Bnrcs25LjB
K0Aq7ftSZj5MtCzCiaa6JKkLD+85Ve4smjeHJ4lioSPdkIsso2vAkw/D4gZQEdbUR5SO3mtlisg+
L1KshmDFCnQ8qYFLvzuMcsa3mQQ7IKkZvFis3a1PyJGhhUQ1xz9OLHIkGnuwr2MopvluULgCxQo1
KQj+N9+w3xNhOkvdWPIPI3VKbm7f1Q+djYh0ypHTFw5zGaPForZ5RaXLT0a5n0sO9gPvEjsqatoc
syZEhPP5HCMZqc/NNwDfMEnRyvNFzUuj/+r3C/P9isc6d0mvH68GeLH5wG3Ci3xV064qdlgsAl2e
zhYAe5FtLcKBffeR7EJ/4btRQGaN/El1O8dQebbThTT2gxbpTGD2PtvMQjYPxwETP7LhCXut24kW
iU1Is9oVcw7ZI8p6VakmV0Gn+RQXpVog1A/A5kUL9ayjzyZWKqPZjybveAZdKGMTxjF5n/fshrlm
3YQMyt2lSrnJXhne2KThm6pusVXs8dhGlLy3KSL/qcb/Bx9syS/7dFHkWR6QYuw6ze//FFuw6MSl
SzE/HulYc+Ii4PR3exj7Lt8RuQH7fK/SWkqIvXWIdGqyfnGtK2w8veeJyoAwuBYaa38AGZkudEAb
q3w3z+TK5yUuhCbxC+141Y0BIdlYlVFXPtxpuWzCJraJbWZkF/n5Kmux2KlqrFa25Uk6xBNgUNRg
yGTnLaZZ6SZwpAAbRzhduWBBh44uzzvNZX/sOKqI27LQsORi3Gai6dBkIzmp7H2IL4yOBuJ80qCb
FcKnoB+RuUK0+u/9KCHVAmJpB+1WAI+d7ejqgU/VWD4BoGI/ilIubs3m4xsSIm5NgeVdalJ46j0N
yDMh9qoV3MsJKn3jvbaMBp4Lg2lyCpUzIG7A9xklydLGdTUy+srCtTc5SL7Pze6k9l0vwK1rmmu5
UaYqmThvcFP0tIERbWQ6cNzsLTxAY7a93t+R0wIB0190DzrmDuh6oBE5Rk0b2+kth1VLhihIFF0F
wUEHAdloZ4Q0acAArdCfpHIuiUgL5bX5n/xCo1lY9SAkn1ChqGGy2oqa/3bEstKxwhGmfzWkJiRZ
UT01ib51LAsbTHfDdqORZOHd82XQx4bGD06wZ2okyMz1uLg6KN4v0nlvZ8Ip81loDYHhohcEf8vG
1QftYYrtQpScy6UcWH9miSJ/c//+sRnFH6J2mPU25awDTOZKhmJlvubYrV3x9BWDjnm7vcgXLe1p
eGdH5XncTHh0zd9yc422pryX/hS8TO9J6aFfigecmeAjezsWefYN6D1cMifSxmxayPf+E1lvn46T
c91i+QgjwPtefzTn6nZYhifOAICAS/Ep61+OvmkUjv6GbZIgiLdoKjKRiqCTO3ZQg1WV8bsHVFYo
cZAjSCDCMuM01wA7firdGQ2ZvF0mbrnyEVjP+6WB4GNxgA5+FSV6hCq0WYI6h67SgXlvyvuJOu2u
jnJMf+va46pGg2Lt8pw7cnImiy8xJSyE42+Os+QMnEoMly5z0DGdBQZssDuOxOq/R1a9CTqKqLCK
JGNB6VSjWAVBfZs7TQxedtCOkRe67jB6r9XWQTgxBKVomrPwUtsvSfZAjpbwBGwqcV358rUbFlw5
Mjvgw3zNMR9wyDSgzfO6ix93tL7oe3888i/fDH8raeaL1xJJmJjM5RYRYsCwQtw7GoIaLl1qk2cC
iFz0wd13rpRosr9tFDZi4bsfA4nnKL1s66wWLaX0LLvKpclRW7GbsmPYgHA3PCcVobJbjLjYoxRg
A27xaKbO6s3uuOXJ+m9LTo/MN5sM/3wDZoFWna4N6xPd21qWeHq4TlqHspUhyiCH4CjJME5oxRDl
LEAFRkNa+aPW/8sTmwDI2EB3WrQQabMg2BWkG7rA3pqVrDUOG3UoI5RpBRZWJ9pjNbzB/wRxlICO
BS23YXkDi8HAeniucextwPjKChokD3iQbgM3X65bfKvrVnpEoxpotp2/CAvLYgtCcU4JcF+DULiq
KQCKTotQP+khmJuZeEguTLe5tLjmkUkjkip+lbP0d6GCw+bUtIy++5lJH94uRIhWNi1uOiIO+8uJ
8EGAN+icxQjG3mv6jn285CbJq2km2LiZy6Id7mpBbfV9APUDYQ4atfRFYcZLjOcmoqs/0tcb26X1
hfajtKsMAfT9ejfZHYyZwbPazwMZl2twKQboB/ZBMqlQkGdFP0i5dqigIwAkQVHF94M7n/MjxipJ
fDVx7oy6FTaaf23w8g+/GEr8rQGxepLkCzw+EdRlwHNU1kwDi+OGC3WY0zRB8VDMX2U6I/aMn21M
dZznJA1apLU+qjCBFUeLH7pOB+SycMrhfqQRqf2Kr62HLl51PNEunvaVFWwEkLOPA3ZVxH6EviOV
ErFQbJ8wA3BAJmG8BXR0prbI5evL+fT515LPQPozGsUd6zhakOisMwX5unw3Zjolq01f3PbTunDI
N9DggUpSAafKfs1qltV4LabUkrjDwEnQYQZr0WPSx/mKWkFFuC0nyZ5ZQW1+rMqvD36i1GBJGvL0
flF42PNP+RtR2ol11bF/Nnn0AvyKtWIM3dU+bSPjACI+YwyoV4bk56eVTqy2lB3TzA84ZHwE+0yS
zyhx3f4Ta51ugUQp9l/9SMk7xneA8EiX4eYIcV2Go977REKE8zf+lcz7NFOadfDakYxHSRxYtMEF
lP/kEVDF/1uuLZpR7zvKUXpYzc8wkg9cMsOdQdx7IX9LUucVh7SDVPwb37IhMmdXMnthV/Z0LThg
RiAGpH8abxYIIZHZf8EWbbd/1tuY34J45BKknB5+ipkQ9si3qNQZfX+sx2hcQAVzp3KjnNHG4q/V
qEgCZp39sHHW41mwEj2o3a6b/K/GXNKZp8PIyDv7Af/1UAEMQqYswtPPdG2fn9HDzsPXQ1n7a96f
FjbI2W1Zb0pQktAJF5w4n9bb1FpsH7Nyb9l6eg4WfP9yE9L7O+dcobFEGip6AUtv5KHCRzSpABCI
Ervnza2e0T/iAlSJTde6hs4wvzmX1d64D8vTH1WhrTnFBw7waaB+0L0csmHLo+2uA+0vANpoXYKY
US0WV4gnb5KRmO0V3UTGYg86yUdhvKC15dm1n2CHXlUmn3lfLiDghDaaEMjgEeHC8wEuCkDiH3VN
bCgtl5Kwj/exKsGJXF771LI15AOHSdzoUJPeelNF8tWrJqoIhTkldM/3XEQVRjKzkFbsDWG6WWbH
CHJ23BefACDAdr32XiD4lwrDxqV0yvMB6qov0OPqwJTkuEv9Hh3DiX/jk9q9FkDOv8Gua9qYzpah
clxlFpr6Vg8zHEdbiRDZJCV4TqRz98WN6K86PvbjJ3HBTLgP7Fmki4E6vg6OBfdrYpWF99G5BhWp
lAF9DmrvTwQW8bOS+xxiPi4mNZ1RcPV8I4ig6juZuT0Ms69YR850jayTGvNIKbp29gEUar+QYiQF
kWa2vhmHQ+7nkfoF4HEe8VfEjkS3ActHN3vsbms1hAtmGvuHKF0Wt7nNN1pD/6Sj038O7a/B3bHv
gISdh+1Vmrgx/r40CQPIM7w2p6jrkv5KMi9VgXIX
`protect end_protected
