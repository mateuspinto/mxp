`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 69072)
`protect data_block
R1ZHmoqJq6YudtYgyh4drZY3yiOQshUl8MeqKxRLvRAwmi9uKb14bdwsjWx7nz/HkJm8FGMjgs2n
V3Ct34tovJcbz+N185IjStCRW9np1OpoGWj62bEu3lRWId4E2Fb4T6mxqnKOCt/z94MXrHjaK+kE
maV8hpwu3Ob6PX70g+rOoRPVUwnHHaNRff/N/sa6soVc2eeNp9Xui2fCub+76Xj0Uavpk/c2bxJ+
H6jCjeE3cyswa76r18tp8Skp1wy3tI7bUVscoACTwgSZ/6PlBOW9mzKqYsSRf2gM6CmvZtfuAvYY
S5Uk+l98uBWKlRmNfmp5af8VZVeEKS+JJVWEcBVgdjwcbj2H6A440zSXGN7EpWSE7MLY27RbSFFS
62w3wo6ogMeFoFezSVoRIAeYFiRdDDVW8+kFqLr1eBnPR4bl4zq9OCEmm/QsxI1pxcvWDZJlz+Tr
UtBYojFmB9qqx+PrVWkb2k1r8RXCQKoBXO+3O6ZRPAXP7k/eQu+r/LqQgPu2d1HQpIGTma70liRY
lCjDR9uvb6mUxqFvzBuz+Q9SlsWHILES3Sb/QiFJKAtYTCGc4yGHudFfhmChv0nBTp4QMgRzwa9J
+3mV633zH9ZwzFxPNlbWcjG+ByuapMC5CkrlUvRX1Sff+Hi41wUFQe6jpxlbNxvH3Q74e1P9vxhE
rfTZlVxntIop+bqnUfwJjgM/GhP0ZVf73LY3VQiRRAHkoTn6JAuN6azPpXJc/xG0SPb7ykHfZ24t
Z2D1Lfjd+Q2uctrIn3O+IUhEz0dSXh+dnw6Nri8hWVCRg6QcEES8+p/bpXDGVe3T2PHfC1d+v8cn
QkBqq9ZMLdBtR6xQaUUQgwfYRyTmniV8U+ZCqvQMSMmEUIHY+C+uimB3vdA3/9c+n/y0baHEaDIt
fcwdQoPK0SOS8WC+5umklrhKkOO8oLiCgW43VFGjJPbKk7EcBO5aOuuLdmt1z+qL6EHNr/p++Eme
o2KGojTrJ3aUC/XvNPgTcKz/nJkEv2PItPCdf/OQ3emK+17RgS4QwTV7G6Vq813uG0v+ovSHdE+8
/bOvaVOW+ibU7iY9FFEb+ffd+Vb85ytejvrNfJDv5ZN7lM5lS2mZZNt6/XDHfiOmGcETPZR2K4QE
7pXQoSnrm75pW94mOMyuDNVMsuqjl5GjBqdhzAES3Umeja2GZRIUsYQuCKjds4B3FS9sIwO8gnBk
jg51YoveKNioqvMFF310kT7CqBvijyLG4fW1mZ03eTxErbxx2yz7/cJk/cwqqNQaOLtcf2fyyR+s
8KtbEwIa7c2e95ehPO7km6CjUJHIeSBb2OVgvC5D3E78tW2qdM4qsAbw024hthes+frJdGsnXq5U
HQum92gdhRSTD1ATJMMJRsL8ALv0RMEIxgvXyzPAcNgbPI19K3ckPZtP2wJLzg4m6ennt+mDXUdy
Zl37OOmJAmeXPHVe57O0+zXTL7f1FW5EhwScxQTWcn0I8z+87n8fvvTd6Xt6UxVJOj6dnN8J3jx5
iYmb+H7rimPKSOMcMZEz+76PU6vYO/xc29w4wQYtwsW6vW0KaSZilSif6Nb+YwPqSD4HemriTlH0
MUcVVPQ5In4sVd4gA+Ac+X1INlgxVdt//q06tb9mOrgf6BTkr4aLK3iIovwRevdcuRQzlf5my258
RPNO09h1ETm5EZQTYB3uzTRrYqRvig6vDo6iyKAMkub+Qt74bQIh2p6kW9wlOuVvhNGFxNbvYHS4
+Y2Hb8e9Hh+rwQ1G3lhnUsvaBhAAFnPesSYlv/F+gwFOJfHq6sCIR9ZQH3pB4llmLqBTSCgnOLSS
EDtwpgSZvIwbJjxCuI5vNc9d6qzGMWsxLDHd+boe+ZTcMxcmbIKOi+hBsq3OkuEUz7KULW1b2T+/
wKK+1S4bvDwrIJ7H1v6vY/ICfVYd7Gqot0+UQc15FWioBupCLU9f2pPNE4VR8fqKkvlDTBkxw72E
MXAqzvTUJCgE3pK7EaaNv0+EvL5eBy2DVsEK4Tgq/MxgQRH3dwkOFLllGXQD+qPTL0WnLJmJM033
9jJzs5AczKkYClnUsHBCIh/ZRJ/FmKGocOLDHtSZcVXhhIvqa4vIf3jKWwklSyuTxC5yGAaLJLfa
zCEjUaoST395VnzLwvi2cIUKQ8zCF2Dy/Njlk7rJyr0aIs1Gn24qkrt7GBdQDLIt1ZwSwWbcL5eU
8ZYSz+GKZio+N9Xvz5tYkbTKPg1Sh22Qpt0lQgbk1NRHrLttj6a0BnpinxZ6ew1YXitWOVTA0+sl
Z9pGD79vgsHjYrIL4gsGEOFP3lz+TyhBgGKYfzvLQyeJYqfTQF3WLG0bQWUo8xAAL2NL0yZsYWCo
Cbo9xuktE6M9+KT1K9LrMqYZfLNWWyt3ya4aLJvrOcO+JMFPRk8hrKhn5HRMERJh1Zv4ys3V5xF1
mB4DLvau4lLVWTNje04hJKsIl7Vb3QomDZCyZXSLymRTQezPb1nC3skxqmcVt82ZSzrsMLiJmeCu
0L/O5P0cws5Bswja6+zPq6YhFHRYmF0fkNFcP2pvC7mMhVTMnLuLTOtEz8cRnsPeLTcoCGYfqfn2
B994kbovQXX1RuZ8Neq8eU1yTW7HPxlRqRJHxCdAlp3pjBo82tIHMKkYwpsTFRnl9tCp0HCEUSt2
T7JoGMNClyPyl3a1tf8n0NPvzeLzqgYmTM0lA1jlJPhCLfaeLwuOI2Nr0GJ9teHjz5BWrD0n7Upd
hhqd7lC1B05lcYU6H2+tRG5q6ySb6AxsMrVsa7Q14v0ALcKB0fAci7QJunZEMIE7tI4waut826tV
XGsqNSz+WdhahnIUc3zw9q+PT4FNBNX4f+uuisUuhWLOrIPnsbqbwkwz2FCefCNcLKNdvRljVvZx
Byc8oHNjBjn7C152xG6DiDs/bwogM18eFQHNgiEpG0jL69dzYZ+1wP6279ej5W7U1QqPXIHGPbwx
lLfeXQ2bii3CpdfwZlMGezvxeskzThMQ4IzOWf2hGkxZJ43bvUe5rw6YLJ25u5nH63zXxK6gDw1R
JVQDk54VkUy7fXsnwZ3yQTpWz4WtScYLT1rvHBpHV2P7jGaoAST1KIq/mEOUz+ITkWe+yh1emCGI
8C4JEfH14Sev2svWhTPk8Av3UtZfzFvMUUbtbCCKAg9tEJpzo2DoPwRPzRr2TB7ct4QSQxkSchKa
DsDNgDQOJ2CrkfMEJ2Q/NH41+zMDoC378Bn+5SbCobGvs1RiOZHIN3CwjO+gt03IDSBHvq1ce7Yu
Cqpl2dYtrCaue5ZJY8NY4bwrBJFiOkf+lB+S1YRy3D6pr2rTvOqg9DVs9vxrwtZ3l06TqvFhJ4jb
HE+c2GeUvB2JWaNyIeIcc8p+ZtoOLoTpG28EvVinD1YCHXly2gJL3mUeOK+WFrjRKPUU1goo72dG
nqOGE2g1C+lMC1rox7lzdJ65dUkdzspGM6YIKQwdS18Ayq+9ch6W54kF7VVxi4pYUDSYi2rYeKIu
hDPbY8SFEcQ5imDOLaJg9ETBvB/+ucWk7S0Bykier8pMnjMWbRGmjP2do89j7iB86TEHrJNMoQmy
vNu9bONoPWr2Zr8dBMsYU2eh26j3CqTTZLWhpADQZfkB/m/2sXagYW5W6/V8eJNBexWYoHQ2i36D
tdDJQSzqPh0t0w7oYquKYdBl7x8lR7FNg2yuwTqMocA8sX8sMs20mD3efp5+G1PkuxOfpweujrZf
tSuPvmC5lBUCu798xfJ8gCmenJNmXw4i3gVxFJ8sKMAFveCNcdvXKbSYhTx5RjyyiwoYyxvszcQY
m2Nkm/4APrKTsjVdLAueu7z5OILN5Xg9rp3v9mhY6OGUWIrR4oIkc4TocvNNZPpLXhUwTtaLk+q2
KoJKAf4gPbxgY9xW0Eu59MRhDIFqP/ZdhY6bTRjdm8/TESvX8VWn6Y6CeKgvJ4pRliG9jX6C5KBv
Co2hYkL9j0fxM9ucPC6bhSLW/yd9THCGKdFPXibVeM0+TWXXgJ06R08yYxzW+LeCZxdaXlP5QPlW
hqqtgxuJ0Av+7a3YIVY1vRmINgJu/Ros+I2cDT19mHjDwAOWRZb7qnkiR+qqOWROj7C8BlSqP5ys
P1lfGdV7JLeQRxjbHHUAGtj35WHf9T8dE5TbewVu6oJs54aFSlVipa/Lx3hwi8RcxuxB6qIF0BzK
wQSBFgU8XSzviZ1ggZsYSLO+bOfqRKPsR3HsKCn7ucHB6vpc3PrfZNQ+xxXc/insQeMyHE99ovoy
41FiGDXNOFUTCr8Mz+GL2wvjISjwZhvO4Pyk4s9QsTCizRPrTpu8o/bgeUdyA4ZKdPKbE4Ksjqzu
2hNeRzvRS1BQ7vgZXjG4I6h4eNuyQzhU7j0zUWquFjow/nCf7hP7xpCTiy3kj8JZOkzkIt032CLp
R4ZmKNwPLGRQhigpG2GVI1z3ABCOzlCllflLULu6PQ72qj2WeqVNNS0M/+P+1pVMDxYPWVdCiVTe
pu+Wi4HD7cO0xip5xAxKbugeGrB2n9StyVKWR3uX0idWBiUjP7PFL7mVt/3gLQaNqdpv5FZg+bxh
jhoqmudiyHlBo/zsqHVkvDsO49jf5C7CudEeCi9OwksVIugMQRXChGFaNrqvkQOZNF+tLC204ywJ
MGTiXw3/ofeZYefXnHqUlrz/rEbgAukhJepwUYXSW1ckD1r4pfyTQZhwK2de2z/7ZKrPw/dmKHAY
Ipgrj01FiKe5jW1PPukfhIgZRGmWERJ9kuTeCNbE1vaHgHhPvmiibQE2WGhh4JZXh9lmFh3pr9CJ
0cuznA17Zuy7iamljmYZyxAs6w0BCVt5Kzzi6DvyXPI+70xkDYrWg1vektp7DuL8+XRbw09I5Wn1
ZXHmYZkO4vTSLpBXT21ozOTZ/RpJIMcmJS3oOWXaZ5muB7SK/p7OcgiF3FEmxN6eNjt2gZta9Awy
xFPN5eAxvwQilDJyoqem4/tJeo6n9I31AVlVI5Wgm8c0MsXUAF0UtnpBptFZp01qkwQN41a3ZU6k
uzYyB7SPQAVvg7YQ3hJBTozDokZ7cR+gNmHw0tPBbRosZAUTAnzJy/Slt8pzl2shVd4N7qTidkyC
i8CE/8kJsYC82Ow7MJwTHYE3bYrRLelsE6J8q9JY7NLo4imSYT04SvlZJz0j2h7ew8HD4ez8tmmW
mzCFeJTt6ormas7LqVqrYQRvt9KoSHuJy3yAoft1ztTNgD9v2vgGy56Iz5oPLN0ryOJQ0mHK/c1j
4T+YWL76bOiXyvrzyei08bPvUh9GQIRznk7qJlIO53qxleCC8SUe3KRQoGbYW5XjZpkX2gIig3TI
9E4qhuaSvj5X/XCBOeVO7ZeMu26k4NJKBpS1fAuPh94e1Rqt9IqNXb6wxSn7AfnS30HXzr1gf6P+
i3h/ysh/MPInQfEv0mXPkGJzuyslbEJP99Pa91LDKRySgb2m3IerTWaBSXZk8wugi4fEPYe6F4oO
NZH6D1wE5NLFRtLV3k5X7Zg2QvphP+1PIWWUmaLf1jYO5yIUuEQQL++Q0S1VRPpHHA2ZsecGJMCF
OjSiw/zj0fEKjKfvYJa7NXCIkdWUyQv6heCAHlufunUNNCFc037q3AgBrCpg9VxxKnKf3RB2ittH
gi4VhYBZWV5//h9JEce5UhhCa4DjP0y7EqBhrmYcUIj2nAtpUHMrJr2mnhOq+E/OfLq4xwhK0XK6
U4hH7p1l9IuVzLUREq5V5Xpw7t1eJNtx8o9Y/Hx2Flwrub2X6mM3JcaUntmV8o9FHmbffbSDm8wc
kzBAMobZEsP0pjNMAa2+JMB9BZ0SuiQ4BOkWt2Z0YV8us6Cp3d5NI7SPxNKHIyA+iIDD49Hc0jvL
nTGnw7kQ5eGAP9jAbZ9NEM6R7+UOi9ugX0usECLenAnq3NmwUAaP3/Qm1g87P0qTcDR6PnjXv0ex
BFMwsBLnOs06fKSv33TZTlARoiJGGBbcDU08MPpr+q/oBAxAITu6mWcRyyuUM5nX3kNL2wOebbDf
Mfmo61B9QxIZGEpn6Bt/0ni4msbghoayfLReUnihDj6VO+kjQKrOR2jA+5t+fhIKXgNjQ9vW9eAr
Ul4X6xUnQf7ZCmUQbznNWXj9bRb3CU+R5FbOMXzfODdboP3QTLXvkX7Uk677yJTtzI1Lsh2j7YCv
AnncRnoKyfwaw+Md/LjUL8ZbuexLrpzbYmdPxzA03MIkGtwpSVHbKb+R2VUXH3xqBWCV9Mz5phv/
X/Dw7VkvO2RYkw8XrMFIxrhAusOM9LMiD6tthVDbIaFJKnj+WIbp27cROumZTif3oI1GZx5KNKwF
fiu0E0WxXH9SKi/hex86BUwoD+toZykVhnUUzLsmv97/5h+al3UyI+5QZ3lU6b7uf3vmRbCPcE4Z
YkfBfoIgWGElwMFb2GogoOv/NFANY4wkURx230xMrDySuvAVqXTzvcHd/nTnPo6EKWaQ/9JPDEK2
Ia5n/azOimJh75cFBDevx/CKVOEtQ6Al7oIjxvfnITuqx41cP8SVuIkGATbha76xRh9KgnuM5HRd
ObtgqPd+m8uWbbSZuHg54s8QWnr1lER5lTOc3idaGvwituoT4l2YN/axSNNqNTmgS95Wsvo+6SC0
diz+vY3lAtyAT9TcxnOl4rbwPJSShhyvqdLkUqn8ypXQXvauQDDERuXGilaWLfpcmemQY9vnVJOP
YwiCmet5p924bL1AEbHzieokkpCKLUhuJeoKr+hYQZaTPyhTE/3b1cbf2NE29XP0b84tgxNC5j2y
uNsL5/5PLsw4uh5p/TXMaYtTRPi58BoaJU5NuK/UThMf6pwyC6xwQfSVydR0gKDo9n/JZeMXnnxc
6/2zD56dsYbCaD1SFOcD1/p4UVEnIItDmf1Ax9VAzJ3BG2BAqi6v10x9qY77J5wHE0LOpzvR58fx
23cmdCmM8tgFKqWr2w7/yshxSEX7tSZDQaUpBwhMK0+Ell2NZreTmfwwdL3WRDePI0sfHf9RzQm0
w6qBPXosJziwXdG7XAcHDdQ5gwJZJ/BHyOlbtKPXNqXRrTM0cCNP7V5108zWLVzzM1Sdkwz7JRo8
Z2nm/56kH2n/QH/7bXeRv5VLb0tGJo4ojMCFK2Te384s1e28GMz8KbkG76PcFw9l+qD/dPMuceEF
CViC5qb4+01TKRUXCQAoVf9RTVBE0jRrugav2qQf0WjzuQNasi2kvPsB0MD7hP/tWpnsVzjfrl6Z
D8OKLEA6SuTtBlfX6uygBy+icfzTv861OPD0Dj7fMKfdkGc0k4hgSYiQBg8GxdLd9iqlcMxFbxva
AcQZL2qll5kXL7NMQ7Sk6UGeoeYExIoA6sqeJ7b0fBy0nrgeMuVQKdz/DYxw38UjgO2vxbG86tPy
j61RoRs1a8P8+rYJlQLgef6RfmHpMObJB3hIK2VUpQhCRhJL7ftMU2b1h+DUvMmRbF/BSIhSFX5I
d3nrzbR5eDSQWXGwFU8dqbIhR6b+3yuwhWuLjsKEqATAMcBb5eqP5gyvAzt0q0WCXAhsIouK23tt
lkEcp3rmmEMM/dp6GUTFubrCvTJoFWpDhtpfW4aKfgeaIuQF7MJrAafohnvl2/Hqg1rtXw5WonOF
Nsz0aOk6+KNeOcgvsZ8ZQtDhACSYvwqG+VnOhHG0+YCO5V80fJEXuaCqSTFAZiGba3uLbdE9l2zN
rbmDiHIj4+yEuh5Dp7wpq/R+q9K6I3S4EqxE/+Q0kV5TqORdwazXB4Q9qGQDQKwMt2VUSbOfOtuF
AdYGihtnfXQcPwzWE6ToJ4f7jR7bDkIOw4rP6BKfKh7An20jrUuFMOTZvt4mrkXje7i996HHW4vy
94LA7ISjsoObThJGrJb3ed3SCkNzSHwb51v4YUEcwCJsesQXoxzEQPOcaO2BKgmvK6izyySfj25/
eDMyix8cLF1Cyl62ebeVz7iwvVjkWpDvyFIm0grYB3rvjTgIl+F2I+qVPNBu7n7C948e4/sAs++E
zDEHeKOJdLwiEYniHr4wwXj+p0TlumPn5vRORKJAloAD0AZC7FY7qxHGL0vvWjYXJCVQVltKWvqm
bw3+d2l5YyQ9QaCteFmo+pieLC4PWy1/CcQh5fHrokZ/aNKXaQtISQJnii+oSaObMQzTcY9tAjiQ
knU3Z4kRRZ3a7APbe0wc/RbsN7pRBKwJVINCuv0dAkPXmG6YVcjw2P26XQB5F0PGGbaM5v0SqB+X
mOKmczMqqNCG95vyhnauCvYX/EoRWrpwivm6VZsZuoSLp9YAL3KDNSSYnWoQYEhU/cZQR/+sLaqd
di0CBMIKevOCWAiicfEtjh6OogbnD93f87ac/8IjEfJD8ngdKMNvbQiYjKHp6oLyU2d4GXOawO/R
gw0/nQHQyoisy+Vo/yx2RfLEWf1F5/oKolvCziAJRt/kboCCAj7qw47ewUHfYY46IE0oAIkwfQ3T
BmlOhaF5HU6gOHu3kdgkLSY8c7askV1TV4M1cr3KbjdQhtW6Imo2ULyoEiceqdI5vc5ZW94CzKk2
hDFyiJYkb8+R9Enq036SsIKEdRegP67j6ChtvzwGgRJIFEjP5t3WTCphGrGdDRxEC/zTrW4oterL
Y4RqQqXy+4nfekieNgqUZWy/zZSBXrCQh42CvtYzktIZkFBlAsFgH8LTVjTfzf8vourdw25//7cT
ne83ye2uJQvDk6kBtmfGHzqcD+IORXnaK/UNaWFs0QJ3Cg8f0vV9fT6QHgqTnf2ExdM4JNgpVaKV
bG/UBG4pGoMeIHb+GXhqpj0/HEeieWs/w3BQguYx9ONBsUzSMQwNjdOwp8o7/CVfr91eEleXUWCy
aOoaxNu9AZ5zeK8+7lXv9wk+vdn/aJ3eCb7yIaqWTcedydZCR05N+KyZs6aoDH/34Ouh7RrQ2i/+
B3GYn0ExlqHq8Vy1z8YTYnbcJ7vuv/7/iAocW7I1SD+cptGkspJMC2SF+YN6wqM7zC0YB/Zc422y
goXZ1NDkNfMw/2+ZDrdAOFD3H0FpxCQ9bPoPvcchJGdSmDd+sXi4FdoJIvo8R4fxjKXYMFRbfVfN
mLQPsDr9xE1mxMGdtp6wvtUbVHHEHWVsLH0pzR44A2CN6X1zIOpJSwfFTKBz8HCENh9sxwnrZcH1
jxwCefv5T/4AnDy1eJlcCo2aeUp/gSKTtN7OttU7ctuKhyOzsBwbFAgIgg3GXQtKbN3muJl5bkvL
SV7QB1a6DO9aCSiL84Axkwxvadhq4z4/Zzz7651DdoP308w36Ll9n1IL5kiu3psBfQ/ZZA6QHKcR
RV6fkP6kpFCfwjCB/PTrWR4m2ZlhAlK4Q8QbIQidr0MKARmdGrT2drSd1xua3GZ1UZMmRYJPaHHS
8sHUVmZIODsYo3fQPCi6KdGIdGNVM5gMtkkZYQmhU+uSLp5HLae00dWak8/343Ioab0bZjVhPCiU
XF/ZW/b55Sc4EyA9hSivwsuGX/sYA3EYJKiPBMAFnr7HruY9oqhXveuu1IAH3yyXwxtJXmywkm/H
aqs3Ycjcp4zjYHZ9NCBjXutLKvzhOPRX4+zCcdftx/ohCwURyhOrbQcDfo/ptg9V8lXuVgVEIOdW
9ZYOGw3LRc3ODgLA+DFhxiiprbTk9FgS9TJL4IMkc7R7TVYMG+pONjzG4TW0cyIrq66WGmRewpTB
/AqeSrHCfgDeRs0xIVmKsPldEuGheAXqvLzgnRvk1qWgyFDk5J/QtJFSBZhCuOPanPO5QwYCCB8Q
gOHkduc1FJ6eZLmoO+F/j8n22xn8fKXbfC809Rrus19oeXeB5vugvTjHBI6Ou8f/5RPtZSFl+TAi
LAu4qgC1/oxjKfqItmW7Cx7uRAzrdexPvkwkFkxhsGl/Q02kVWv9ql8MhRKL/nrZRnvU9Rb5V/QG
OVkr/nITeZxCxL0OmFAzdoNbZTIz3nGF9Dao2+yxoYOdBP+rX5UZUF8wD3k8T9pqMxOB5wM4OZat
dJO98bSGnHZl464rYlNCGh0FY1L7aEqphCgg9h5gQ6ieEzsZXv6aWUiaaQC59ce6Ha5gbgtWXZlL
liGDCTg/TBxRL/m7Nzj+IsiOW/KmeZqOQJ29DMYq+ZgT2/mWqO3akK7OKV6tv3t7G7viqJANdIes
hpzZkZ2SIwIZ6wha04MGCGGIrjLFoh5IkVNZWHo2VXQPho7YfHxu4DGei6yST4ht7VI10ZoM6cEy
ppwUatsBBOIUEZcIxkD+UwSEvxwYnJDQ9oRslHxy258rhq/1ISxFrO8K5OaG/RJo8HAhHTKNU2j3
/CYkcF7TnXDyFvsx87Su5MEFgMoKNQzBDd0aCEnkQTYawHWGksFFO8qd2RXsZSbEDvv/Wwz1uRBp
UuvatW5Jz0Cu8OPRj0Aq8hCpcvTk8oZECDOpPWY+y25SA34ivCLyP7gt7xggsoUPifp+emi4Ahnl
UrIqCm+K0Y6QilLy7meXmxoK3yhtac6z6Xcu9vkchZDWOD1grqn7gc/27KQDyOyxZwBGFJtOeHDl
lHtWL8D854auFHrd9C6JXJ0OVPzQrVJTmMVNO5uDbV80TAzsNtyZCLk1/QpOiRDjgioE8sePTPg1
bfmQDx8nAp4SvXoPyJbBp6vM1t8i6p004h2JglKbffvlcX3jafIVrb25DLYSddt8JhHCC39KMyUD
vJu8znvb3Fm35eFYDWbbwRb4B22CAd6D6EC42s5va5lQav4YYbB1bWQbRCKajr2wOLz3NaGyhg9o
LDiY1trgL13lCc9suiuY+DR43u0RlXy+qVWztNIV4JqgSQtbiPv1sd5ab6QvBODPruRni9Lf1CvN
TN8GxMi9m3sredC58e/d23PGtM0pqFnNK62Nzow8suIC92r+f+o3hTX36LKg9UaHp+tIcKRUlz3H
6rTkhrCxwkSKi0UxwaIQd1vHHt3kbMihjIDtzbkfkTIrRQFM4KpEY3FNJvN0p5YFSHgkrOUFujlb
dAM0OLfQsJa8lVqyG7zRrSR8mNMcJDf77RhKOfRiT2VMvbRjQlxjTOTTsuhzViNcgZBev5nhBkOK
RNqhE9OD/Popre582f4ghUMHeBfMHjTbOIiHBRLe2JqfxDP6hRziC5PwZPsLTCsoQCjDVjf0IvYw
B0L+rrE2uLTaAkLf+33N/66ThGxMWheyr6s7c+oFJbbpEKXyHadmsoJMwxc/+82odtRqBs/ZZkhD
FCGMZCYhLSYHoU+2WbypPoOzVeENeA/QntAKcHYMxAKi6Ncx3CZ4My8PkIFqUYiJNCjhVQqWZDL5
iXz8jNZ32Nko0Gnknd17Fk/b/McGIb8CMYxN/N4Njay+iWk2BL02J1QPpzEa+5zjIx69dw+jC4+Q
BwHY+mk6hkw5wGYZGnrkFjPt+J/sb3kODXpOsKjFIQYMmTLIL0AodQ86DXULlDotd6UAjitBJ8Bn
AkYX+CqZhFCQD5EfsD5VU3V1cqCakAlozZhSzx8dx8xb5tvrBp5pxCzG/CBiMhFSwdfWBGfKetuN
Eu3Xz+jfXLzI60auNWfEvv4hSUm3I+/igYBkZ7SC+8G1LIos1gk51DD+vaGb4y0HfH2uN2K6OC5I
tPa3G93QeqXKEmFDZEuauPF96CRPUigmjWqqAgl/gTyM74LOBWAfVCkOH3HN68MXjxE/v6e6XGC7
cI/IfHrRXK18tOGIwLeVXcFw0VUMA8DuwEY05IX4DOuxc4cOG960d0FejHribmnPa37kI5kKnQP4
6vRirANys2nMtjXRaZz6Bj28TkSYztFuI8y4kNNfPwmpSYYRCGFgI7prrqI4LFJvpmIu2B/5CzLp
ZzG3cB8PYzVKsU1mOVmpTBP8MJoKRG1dYS6xBG7Eo3BgBJ0FpUDVwOWjOE6xDzXttI4xU4rq6g2E
khuzKYEknXuHJCbhUSpaZfah6/NlEoalvOYPynzyJcG2pQ7hH1wCZVcjQwR6N9RZPInrONSZ8geP
4aCAP+/sQAnUJCJwJr0ymRNNa/02D84VgZrT2KwXy1KmeO8hE3fziV38/9czZK/vY+B1MzgyHWR9
GRTofsVnPqvv5PTiZ1w3pJQjw5nkFZVQlBG5fDnOTQxlsvTKTjO9zfSHtIXMYITT3EABfwfvA7xk
8lP6UFBwaEJa30ZYcIPmAVTpcLtCKzF9GeUrOwI0FnCsAHZTuZ1UNdl1+VdOiRENjOzq3EEeFj2Z
NqvU2IApccBu1sofUx/pnz3QSVQ0JbtSHvKUjKmK6+picQffyrQHNoItRA8Em7Jot/GUG3YN6l+g
2eEmwLIepnxMva/NAcveLqcatk/6E8sqDPfpfxbS/c9upGvyqhwpMFW89BuPd8es06q7gWeGblFc
GJHORUrXiNRv6Yq9ZfbqRcbCpEwr+BiqYpqNUUFcZ9zsF1gWZzeOiZnLfOb0r8egXcu8Ou9W2lWj
NHtJaMGZ2Q5/qIxvOFJe2X4kJ3pC+l/cxQUzhueAsMBNcD9rMgyR3CsJXo0pQ/1TS52OftmXxLzx
bgFN9WC2ius35zQmPwHAevwCQXF+tIUQnOo7GR0ClHHmBT9wb8mpcQEguqbevqSEqotp50uF4MIF
pmCrryFh4TpBqQt2s4EOeS1o8gEAfQAi2YrrPmzsw2jq0F/uYJzq7SDn82pEAmOaMrFgrPFhUOpF
yy4QHwV+FcxaARRNmvJfAJuyDLcHNnbkiv46P+aITi68HeWyCQaR5xXiMmoxq8W87w9T/06OjAvf
sSuWpflYjKsJNZRf33/htlH1VEOuzB+TDs+HrSw8kfXERNGmNAZQUMj9H2miLVFvCoPCAFnX8sdM
C0hhHcYHF4JqzavGMUOBkRl9CTkCmtrl+vEcRo/BAVgn2wDKl4EL+v5NG6dX/gIPmIXdqc87J6my
7ZmWogQ2JWPJevh8UEYJVbVodU+zhF24HABy98LbBBYQ704d7bIiursTVd3DJhT4hPaMeGNuCNLk
MXRfivkf+a6qOyoBLroTJWYdYthqrd5y3Mk507oppJp/sjLdK08cjc+hWQjZONhqxr6x2YaoVZ9b
K2kN7xAbzJ7HHrcL7GagIiko/jJKPK3QpRnc3ZAmgxlxxIt7JM8Yx68XUCyTMajU5A2yjBU/2bo/
BeupisgjPhFpD59wFStJ3FPsknx8C+GJ3FbGQge2FthGgPo9cOyhQd4SJQd+wL0KBdi+F1DOOf9V
pUiVqL+5nwhWr2855xLWPMB4wyLjHudj24UB4mOS4W3iOEiTmrYiIZrulTOFdYbk7VyATCuG3ZSs
Pz3CR5K58eGrsXOk7d+EmEL9JTGuW6NBPlunK0rBcYbHX3TAeMa52yUEzVKQwY3GWczP/tepiga0
ki0NRtOkLjfuEKTITw+P3mZuodXipfN4tqXm0Knliz2bqv4NJfze1s8jVRn9FfXRIfxJeqmjv/s4
4LK6B900zz3t4sCWxsG5lSfzANYB9NnM2ut1F+pvugEFw0XLiYlkHuutFc9xJky/7ycTFRdmZwzl
ER9OuWRTHB0D4tU++ZAN+60/kAqtLslLUHIjuYss+bp7TyiSqhPCETEdfyAJV0RgE+XfpYueT0at
Mwt7iyR7GBt6dFxVNak/gYHkyrI6MN89Ix842uNUIRc2akFvR62Ah4DBF3nxVzRxGnf7ejN+h0BX
kmhNcKHmFFz0ykYFQgB1UrmmbLmpYlllhLbh4l65lQlEFi7IYB2MuivBnXZzqnH9HNeCH0/xbzKk
GDVIsCvcL0VHcspLe9gyhbHd66RYrnDfFkT0Ho+GePLEcO73zoFiwVbavcM+siEOaJznRvJB5dfk
qCW1opZQ3T6/O+m2R2oUU6Tgl3BGrZzMQHQSqINuqOf6MqTrVy/PmZ0WZ84NRPIHpVnhXJ+yYOif
vfw9uwhOmFRf4vx4YEMh3lUKNk16AkFlKx6d2F2wDlQGmAaYM5luRiE8YbWSFPw5jH5k63eZfNPb
eNPtc7T1KaMzZ5VtZ+JJHdIK2RFd/lSS2LX3Y98/czo5u5T5FuZRiasR83v+6Y5lPi9cq/4SXQb/
3BYlurvBBEaSfNZ7Mraff+yzdUnVJiu1rbghCwWAo+5bUEGRJ6N1vxCS+TPaWh2OgUQk4IcER0Xz
oCaoqWRAQxKtZRksNrJZmngSDE10rBI2RnpHdrEvcRWeMvdgCxqfuPWYyy/pmEJG1NAJASCgMav/
RrM+sjR5qHpuPuH6SL61pHVMywMFDH43ewVvZOLWKXFu15bpvTZG/LJvdwPnebEHY53b81KZT1Cl
QiItR1YxqtklDmHssRnD97DJDYm3oR0iZs4V47KpyCb8M9K/o7JCj8d0V8jjCTcphyBkq3sr013T
9+B2h1JN2LXbBsUqQtKsTm13JY/OkWFecFoJwEe3rvALHEksKWpW+cruWqnoeLeas0foxhStHH65
yfCiREuzsHZntZv2CkTJW8tBAr3I4VxMrhUNZm6d3PDtgGOV/LHKUUHfpZe1W/DAXmMyOGEV7WuD
y53FtyBBlaq6BGLECy1/69uafM2JsFQGdpA1kvWNX1tI9/r5TIb9JQ54E5jJjEl8/bDod71hGAqV
dU/RAFBs+lSeQIQ+3FDBWCL9bhUrfoaBk40X0V9+V31C1DuaLTEWYliFSX5poI8wknANPcYxWAof
HQ6ltYD8mjBS4rkOmBkDwoSwU20C4gksUquveYhyd/iyj/7TVHE4Ubg4DTcp98Kj1wfL2KTdLLhP
bH3cf6RRHcrz59qVT3yvWQ3zD35VrdW06vNdVjfU7Jo8rXy8lhSJauId33k4t+dkhsgdnPM4GRhJ
qz1u8ezXzrL1cUkeyiDTaCyfjrMMgNWtOtv6FOAYiaomACbZoQpra7BW8VCvtZ/owqbVGzL3g92O
qJNjrI8GjvjgV03pt2fIJAR8Bb/JVRGaK4T8JHglABmrThCUWajMbWGA1vFeLLX6tdzIThlsK53S
8EoR4BItVKinzXTu8BcLZnPX87eafDMdGGYbyfUcUffkcmo8/H+6S5cGy/Hgv3cwyP2w5JiyAKC6
dDfYrdXNYKBiuRaexnF51KzEsHTr1SgukWEwpjg4kSWskYHWMdA8zJ+EVT6q2b63YtblIh2+aoKT
C6tm29/n7YJTZCUDDIRmI2N3wmuQNxg3dcrhiKedqRc3wuHis2SqqMgEDSpSI3P/1Q/4xQ0Hz2X3
fzKG6uCuUWuuVK0TPsVrdVA08KaWCkw/TQKiuUZh3Jb2zH3A61lHfI4faswI+X0selBYROxCRa3B
u+YbraQ2+SMRZa55iYu1BXm7lQDlZxhB1nxBaYQSD2gVYrnYyOQWocn4+u+DwZ3sJnvAX4MgvrZY
1trVqz/HfajQ5jgjCW4CmL/f4/D5/6qJ4UxP+4oQf+OeDDwvK/h2A8H/nOvQifVBzLaiZu2mjnKU
Pp2dZoXQljiaHpyq401K0mgrLHp6TdGLDqZpP0Ep7X3iyBSq2yK5IYXPZsO7/LDQi6xEljdSgb0n
L0Uk91mJ2vdFYtW5H2jaf065fSaMKnG503Jup/xT60e+2PN7Y89/bJTpIZ8tLv2HDriwacENeJ3p
dCEidTbM2c4pXZHfTfRQZ9z1S2ZXNDLcCxFVw1i5oIOSD6XAZExpsmhETHV31Q0rlQYBjnVzSbh0
dZ7nPqOXeitaGWe8vCDUsi7ZAjstJLS2BcOiwpirLCxsoSEZM+CLy7iIJluUdMIFhqBMAGPo3wQU
GKv7Tz/flpkrpFi7CR+N5GIinzTVjzOk6zatqpKOEF7+yCiupZU+eKwin+xEsFkwJ0uoAl/BOyE+
g3xSoCN2wwzq9Ll/cQEYUT6/05ocD+0wcidY9tWLJkuzKaiOfJY9vsfUq89cOQOE2LXxWUVy7QnO
YAp6mDUyV6THVTtteAKt0k/kN7pERmy85JFisHXsBtfgu1c39Tde3mgT8agberuAjCs1+JfwXVsG
m4oIxsf9ZnBB3x4moHP299cEZw4r8vBhyroZggIVNNP2a/wqO07BZlKu7tyL2rKYNhTDtb/hdi8G
eqKsmbwyibxxijqfn/v4yFq1h/DXvQky3YbPV2AIpqJkFHpLsZBdNVIm8BtxhnoLmiUjLSWMrn4T
DDb5m9oPZA+bwWmMCU92BS9VF77uk3ZOQvWUX7XVE+WEM3V2qXL8WgMPVhw1iPUFVaozCaRfsIUL
+hQPIvrE38z0lni4lC7y1Tj76Qstt2nOZWd5BCLNHXPSAPESB7KFI/3SMzC2vt3uZr7X+FzGx/b9
zWB0noNdXeBzypO5WzhqhN/3Qa2Z1upJw2Q8KoORZSoSCzmW9kQuMq3MJgg5W4BBE+vzbv1ImHm4
TYlthyNcReO1fkJfAjTa/aRPnPzYssh5lg1RxX+IQZRGQ6aO8XZriR6/Ll+bONwW8Ba5YXcgkMgp
2pbmHKkSP4UMAqwLXYubJ1ibG2Lr3aLjL9YaDDycWGl+Nr2a1j9G9Jb646u5nhqB3TlrmnuE6JAI
maponHtY1bS1FZ40o7rbiEf9UPrMD/YOIE+xFNtU4GbHAIjfEOPQZa30sFaTyVxxFq7oYgSGk4/7
OzpD39vFsgE1RSeLqvwlBSLNwjK0jfMggOGRTII6DdvUL9IZSSVuFGGXsRq2PvpZExToZxLi5D0L
yPaeJj1D3UAuqAS2kkzZmU78Po9vziabl6FWwK6SOS43gJQw3uuhC/DDwLXQW8XHOBdFHsZTwCUK
5OFyFaJ3yJZpKwfngD3urz3Mrnto2c7RXrg32veeUs6DF+L0foGhPwS9JjsrZkg6ByYUrZF0EYDL
Bs9Zou/ifKGNj5peUw+9yHsVJSoIV/uhCMW6tdyFISKAzuaF6b0JFEaX7/ON4Fbu/8Y1Ad9I8+T4
vCSl8wheF9huO5YCEiuKWTdN5+xhGQvhbsvJAd2iIU7LLbU/wqNInOPr33hfvYQGX73ymqQekE23
XKd/lYoqny8WrqnFJTWj0G7rF68JFvFTawJBtFlUG/WSUwof44MLj6KjPu4I6+rbsQLXPDjw1nKk
zUUGt4GFR7oU94RYeBRB8bW3i/Cx9vlsonNEZOk3gPI294cRSWLFFisRM/1qZynMKYRAX3zM3n8X
2LtoPa/vHwxazTE31WWdTAn1tgP1DFA5nYNO7XiNLK9ZjKbCAUyqdF8GStSd8kjufZzE8WxPk3TU
V3tFkQzgUD8cliGw/B0HJHGtiyugM2lFTFv5VN8ulkf8eZ3igyzMOfVlgFSl+WGD3RZMudvbAx2F
56avey44H/BCJ/5fxP5r5yNOxVXWLSeRYVqFopOroog+u4PDiVRS1R7vCtB7Ac526CrJUUT8C8YJ
qkv+wa2LVP5a/ITa53daxaKEIwLIJj/9RowWWEwRYV4kH7lrm5yEUJ/3YPIBNYs+yDHgDPIBogrI
db1Yq8d2rcBWimjtAjFDulQiAGAmhwV9/pppS5IWQU1UGrvuxDYn3s5WCSHv4F2FQZYcmJdTpDu9
2OBAvqoj+fmeaFJKLA2w9KH8DWXwriFF1G1xLcxqBL8mtcORNr6n3W58BN1FN8CMhtI23UC2sbzx
vEDegXrYl+hgLdBdZWrYpJbGuIwWI2xlhK8Jw7RMNkL60vIdC4Je/BzPvynIGJ8WBanADp1MhfVG
UUNS579fxOXLuIsVQ5fh07ynXAHdd2RQsoRTPKZgvY8xGopiEE1Hg57SleMKgTWLcdLlFpCOf1KP
DPKsIPnIT93xQ8hyOOILVYTFHrD2t3y61AosVkmclxXxeBtqVS92EOFXodAt5YdQzfwY30vxPrMz
C2sbEChXJazktKVLpu+Uu77bgGJOIapjTN6VXj+XWaKav8oUTTU3Yyi8fN2RN+hRWxARvUtfBnnE
yB/fZnu5R3uZxw8LxUwMKKl5WsCbkCTSdV4VEp93imETybU3GVCCB+bSW2br7LQX2hjsHV6ZLDn1
nInRkQontVecaKNonIucgPwW4LPk8jYnh8cvUjqF/v8iZYvQ/MXOkJ7njw/0fDWC6j12HOUqWiRd
HC5KRkovA1GM1YTGnGAMiEQPBB4+R8g2RVUuqE16T2sXQW8MnimKMzU5Cjpx/tzt2HjRCFZO5oBZ
kawLCPtQtKQyXfbGnpIiaC5o8K6/d7LKX47Wf+LDIb8wOylnnTGCsPnfFAKIsN+u8pdKjJdvAZZw
U+sP8hdocjSQ4DSpNg4aFbe2D2FpUDwgB1UNxIlVq860a7iTiFO9i7Y/eFT5qSLRUkr9QW4Upvdj
RAtxjbRJ0dWbZSb5K1xi+9VabKoXZAdlC34EwMJt287+C+YIQrJqu5K/MfnavfIxKogIo+RVY09d
piDZrNAvu3d8Zosn3Dm9rCS225fumxP+AhsQvWimjDd1jG9GiDYY0cuxfq6nOgjFaBn59trrl0NT
HW8fm1aCU7boUHOBsdZ4MsIE4DWiVb3fa1otj+e50p2NYYoA/vBudeEQtvQR4OneyaDtL9+PFDlt
m/Pe/+VMztVtfgHAPNblpU4fAmIl3plQkK39Xc5CPXeXsPa4H9zhw6ZHW5mEmORjNYfCH4KE4EkG
vMPgwjhgWENxfV0lDpWokuWQBEA3lQR08uDcpMcVxIGx3tRyuCI8ZsDyCOyxwoScCOG3tXpjysYr
vmxAGi99a+NWuBRkAI/bH3z/q+tTTK7tZE0L5fuJif7gffEg5hbFfQYAPh72J+pbZhCOgChaeEo7
yoF9udQYzcsnvUgEVPFP3ALKOztXupO2d3hzmkrMvHqlAwBl1bHhyYc1I9z0IYpTSdnrC8mXgHPW
uiBwhpQiuvTvWZGrFkPfsnAIcEzT2o1yMKLBsBxBy07yl5cT3ZKhiyLlHdeQZV5H1y7PYnw/KgVc
sH71S0J/Qj+cNSRuoczdUe5T2xlEOYz+2EHivY4y148MDoknd6TfmB4hGmm+zMggtQceLIn08r/R
wUtN1H6NYFgycuDW7Zi06Joyb83r8tQ+/pC28fWSu+siJG68GUopqVg4vxOnbK+zvNFWS97wjWRo
ubFbS1OgwpNGZsxEjgwF1W/Lg9p+J2zyMXdPFe1xiQC1qB0xJpZRo59bqw2zNdPUMy5Bx+4Y3i8M
M9NFtOlHxtEExKselpi/M06fkens9ZtzOSCBCbqwC1PMNLrNEB6dgATeMA6kbVaEX+NGyEot10zQ
G8mLg3YXWS3m6CpBJkOypL+ic6InQIM/md/pfMkvmshg1lwr38gJ3o1pT4JfXEiX/leF8lyASgSm
OaO2YaxwYSUPmOlGMjcCAPoBIM4qFVYDjrO91x9khtzH7SMVUvT6gfXTGbD1LnN/eC43HvErC7AT
SUsA0kxshiN/rJj0AE3jnaU1r7VPHIxfZUZlhdt9rG2k/4rmtBnpY1oNCp7pwI3Ml6ywMiPnVgpf
5VL5c6BIk7aits/4yLqJ15bTGtGt5CZ3L+rsKHZ0nXxnUo/kXUqfjMob/qmLr922BSOeoMt88F/T
Of/jv27mYu2lb/q8JBfGo1P9ls8Ts+ZB9z2fmITdinxtEuD77sRunDU2TIZVJY+wbuv6t3+uz+Jx
GcMHKFBaSE6aJBqEojsN2TnRBwUyoFNxeu7H/riL4Qn3fy4gvK6UjcnqwE+XtRm8UylFSvOq43Kh
iRFXUP2SyCWCQ+Ot2Hi1UH5QuQXOJINdLtr210IndXAdcQr8YQIbAe2gENPGo07ogwHSL+YzkqfJ
e9cYk/R/wL3piAp/b/UYfNWhSXXWwE/jxK+Ndwl4CyZ3xsvD9iUDcUVMOMj6XyiEWsF/u7Sg98Ja
cAioLgb9Xki1AB74WtJXq/dRznSBlSvAaT+Korn1e0ay/l2IJbS1xb50oIFXRXtZMLTCl9wHKdt3
7FkvgRb2/8KkOwM4PO6db7wIWJP3dqrZS9NMros90Ox96mqU14T+vdup1IofwYTECaU5tlPPrNzZ
FD8KiXJm/VAePsGr1rMi6wNSL2Plc3fx9Vs2yzosUMHXpEP653iLqryEfiyIFjl3YvvxnLyS9u/s
/UzogTnK/E7VPLtAiaum+gCtSyoOoVZdaaois//Sz/M8H3Qw9jE6Op4TS+f11A/lRRXJGCZkB/pq
zN0a67xss0QrUze6CTn5Qs7Ht+e5QTlenH97xV5K/kqPnVYhL10M2LtJvHrMSOKuBDjP6RTN01dK
+xi2bvjpvw5wTwBgD4/Pd294nlWM020epnrP7fvLoup4e8C5myuEb7jKmYiCWcu8m3A6zIpA2Kzf
1VFUE3tMD2zA5HR5nCtLJLngQBWfnO4tckY8KYiG9wNt1o9fCKloppK/stpAsJWbVWdwuNYuoTm4
VTI8sC6SacSi7mWu6YCm8FnkRjl8LNw2CYdqw+ddTeiZrjVpTynO+xAiXrkTic5xmtX8xKmEH1X4
6GfsbzmB/x46MrE9P67sjXuSrB7QoKCxC0aN0htXrKbDwSOPRdbrQwoT6SaMmwyWb746Qitr/BiZ
aAst91w41lkMJXWgvro5SmxUZ1K6Rb8GCDS4hc76J2gmlazqonM4JFzawK9VbuEcWJdwF1Vrfu/V
WPLvdVjND53RbI2g0V0FhzgZ6fHU/5oRrBOwjTctzmURfTTfxdkpMkRM/9+OvGJJIOviSiI+CRDC
j0WUOtZBk2vlBDuHpep6NSEF7If7CONuBt67T20hgexUlIxVvlY97uGREHm4z5+xlH4WVM+jnhMY
vZMg1XoYq+6bOSRllBnIxA7cb2inuI2ctGwIB+FoI5BP0afFTE9ZP10Os3XuguTCTXx3xpe5f+Vs
jXs+K5GjQaJVSpHeAEnxVtBJxCJFXLTEzw0zJsIcqqraQaq6YyfzzW6HwzsFz8RUicU4SxUsr8Di
PROs3GxQYvEFspRCC7NZrnjCDl7G3t51EeUVjqNxGQp3ykdxW+MWpgt6n7xP83Agqe0f0KPhab6U
NMlnQsI+55lACWtxg0Ja0xBmhWYP24QaVU2MtmEa2pnU1V3R8DbSOgiKj34m8nsKNiu0DsNLBKub
fLEo2p0AdHraagUukH8F8ug73LsqJ5vro3bA/cYT4HpChQybm9PesOKGF5rvC2vMsAiTCI0uNHzH
Q77h9keBlK1OvuiadkXNRIHwhGrBOmNyHUrhHzZcD7g448mCmwdEXYBH5KZjrDF1dluyq/BGM7Ni
cNfrf3FZFFUAu3IwIABv+QmMGEJrELr99CvsX6yfoRJ7T6KoCyI/B/Vo/cP3G+QO2XyDMlKf7TLa
c8fZRTpHDgBTfprEZHeSbOClPKbvb6i/QlUUBGFoqzfiWracwpgYF4emODspsoT6s3Fd9joQ2i9T
UWpLhdZjXr26dCPxdlGp7eGiubpaQMPCr+mFOBnQCnMGZ6mMNsyKQxQQEU9P2GGO2+membrlPRTg
KQbaV64XgbDTm5IxQXVzmX9Z3wpTLmAPjpbcduZ1XG9vla2DBR2U7ih+yyOMzBauXdj8OohWclll
EJp9Ds+OUaH5uqXItvWs9V4lieMrcCoIy96JIkiBY0gAYXGQof8nH+cFBKc8brWV3Tc0Kr5V53T/
Hjcdc0faFIp3tXlF5BF6ybD0PxPPfkE4a1nXncEanf3NGe3m8LvdxrnwMgHsVOREdygiMsvAye/a
JEfH6I4hOHKmMqReZ18+9Gouq06KDVCz2ZMvqXBLAZVZCIQ7sB9yz6xOL4jrh9GyRmFV98nRQ6A2
0cfyC+cy4Qr0xjDzhiesRpTiGB20X3COuFeIqMfgd7J50dym1E+ehhCy1kRHF4l2WAxrwF7tpSCh
FeCxbdhYwBMrSAkOAoC8zDcjp6tLIJTdUOYyZ0M9D456FTfh/vcDT9BuHBVcGSHWaKzcG4PHLkw+
oYCRFjAeWLMbjEhpukKM7NnBpXqTpdrEW+2E+mTeV1afFhVp7iS2geeKlksjE3rSJzGzvTrykaEB
Lf1GxO6A/iZdlq4CdeyATX+TUjXoKMp+kbifOUFAJKa00U53cCecGU4wvu/DrP13oF2wP2QPTsy8
+DHfv0MgbRMS4wHfJ/OrwzeEOh272NLbgq4pha6IvlHt0EqxTgphotTnuKlNsQg4z4fJfrJWnZdg
0vt39Gi3Zlggxukr47f2S7XynGKfqUToCjhlmigjOr6wbJCPiamsVAeWGqi60ELBvTvkPXfdjixh
jRgAR0wCPslnHJ/mj6Gq4CyPtLkAzA6rIzf0/hGX95nqYpi0VvYsm1Lp/Zzeh3W8lzTZByN6SB0j
oYVRaYtl2yx3bJ5JsFbWwTT0vSYFttG9xFBXR+/Ibcy9tix/Gb5Qv/P8UZBTEzA2B7aksZ2Bv3Gl
PgUaVKWD2TXGu1fSJa7kF48Dqsx7qZ256qx+hoBt+dceO/LSSD3Tm2JHuU6hUJtE3uAXU0TAPLeJ
B1A7j5VN22n+vU1sPUoJnLFXuzev9NznDqm/iQN1p5xw96aQ7ahpCYo537Cy3P9Ev42BSqwty75U
JmDjwLY2b7YJIPjGst2F0q1VozlpSzbcVk4QuBTS7vryC1aPkkscf5QGRfIPlBWP5aNvnu2X6c2W
/LK+VsdDZhzz8ND++amf+GKWDIB8+YCnbu6yMGE5Lprs4357qo6MaJAMdsT2r9CM7pgv5QvEnUQo
oNm2QM3vPbnMJdEAFqs9/Gq+f0s3M/JurbLGCpoerKG4p6tZKVF89fXhcGU/2+PIQ08pJhpJZb/K
xhvryk7A075lv7ItfsU8n5E8meVKrV+/rHbl1+WpVUU7KNUYMOHxg+6dDPdmq0u8+Nq72P1roBiZ
D1CajRsV1wgBvfj+nZgt1YkRIHjDfQNQ6SYbfrwQR4eUgOEeW7f5IJjFGOn3OA4crLs2PTep/spQ
MBpnfQqfdBCMpH+LbiKRcwDUuRDhfo2Ye2xMgbkAXjzRXfIsGck23vDCMmepJnAEUMqnnFYNaWdC
Av7+4gqEuRsj7Nz4xX7iNIaTmpcugz6NnWOwgller0/JhFBfF0xiQo95QzqIAXCUXqySLLZUn665
4sjTxZvUUE5RgI9A+wpbJbadReF7p5iHxI60N/ImFP/froFP7+XydyPHy16sgH/jAENwfNS79ZcT
HoUZZZ2XaOql0jWXKYo1FbfNaPwYsmHHEcK/SlNhPxLZmAWt24hcOKN5oH7RBySf14uxy0Gvrocu
aLkMq5tqXKaV/2yXVht8BNFNrltVy1vRy1zeAGuXdXhmTo5eq8eDOjZhwOengobpBijQvavoFw2s
zW+bW9s+wZCQklbodMsjETlunknwfuD9N556e2oBQt6fffzSVa/dh6t8sMp6r1GlA+qzmzgMCxnV
wZ4ZkQxuwO9IGT2CsmBE6mJpcxCFr/n4XQs+0NxN3ROLV150HlviCayPrpcGFIK4+FYtnmfN2b+M
MWZbkNU48VvV1DaNOyNU87eqqLACeFshMTTTHRXD468nll0VphOWfGt5P8/GZcJgPwW1k95rZj8e
vNXnPcVUkbX6tC08UoN50ZOQ+PJWs1pqVLlMtlTBTjAr5nXwJZTDGGqZQjcvAfOISOkONXbH/5TF
3uLNvRkraJUonbSRNfKHUzYv9pQ6gjFeGNk9EH5nSwmEPVQ9NB0iiR/5ViZ1v1m0br+ldcIxUkJZ
UKrETo597Q297+yV5MwMbg1XlXjP7MfMpcUdW/jj+b+NCwfG0IdT2YXMW2ga1FREPX8tMCiEIsKG
Bmcwd74PeNVeaguQJ8aIV/M7MhvOTmqehNge5F4A011F1ByUsoydCxCjomlnBOF0L3Zd/WA+t6gM
ibL6OzOqpOTcQjoNGWvuETe82KClUqxNibNyNuiAzkDoCfz9mT5C4zI7rYzIQu0tqygynJZdXTra
fWgjLPw1UB6I1LbvMLKaVzLSQMjTj+UadPoXp74Olxi0AW+ni7RJO9/WksR+7lFAu460RbbkVIo+
qwRTE89XUHnxJAowGWP8vlLNM87wZcb5FJb7yylSP3Vu/fTuauT4c9klGsH7AMxtH9VFP92dvYTG
lPbYTC3yX6ytbIUCPSt2s3zz1tteRvP5Q5vYGTg/uuZrUL65qzPpfmE3BaXbq2QP2ZzNlGdA81fA
TLs4sXmOSDQ5Fc8XZu9aKSV1rpU9mnEnXIzta9DzxOLdqMQYKCSrhr5fzvkLbAX0A4vulQMO9r/y
L3PC8lJqUv5YbOIGQCPNXI/x/Bkc8YClRWL3fhnsC3LIuM54xUOtZ/KcO5/VRp0IB2DwxgPP11OQ
H+b7kw1CGu7/+EDhGNRCu/vCQDHOe50XL22+JlC4uAIRcndoiCGU+hHkdVekhgpKssuvWUL7SIqL
XuhBpsgXXHDzNp96cOJ7v7mkzRsL5X146eHgB2CjJ4fFB7jpoIEHaob0jDkJHhpD6ioFGnGhnU2p
rngCIFYy0e2U+wEeV+4x3/3pZEcMhvNZJ05dzwrWLFuYRnOFVktAI+Qy+8uanK9cEC8kzwNsgvyn
LtUAUKbZYjdyFHikRHM30bYDZqp8DBsy3J+08pofii0/FiR1CXFff6+AgqzkJB7sZy/iKAovzMYA
xhGZdIWp2EM5uYON1UHj47jkqsYZ+o2t222ueqrnC8SnwvLBrKrktPfib4JiRDlNR5vZ31pJVcEA
dyFt3w0GP9LdVYzTwFsoU9uIVnj2vw6YMrAgESWuAoQLHL6Tq/5bdTsxwvTAl1PHy/Yc8IdbyoqU
xmsU7M4WPi5OtazemGlkZDGSHexSjXPLVO0P7vdc97BsRQsnH9I20Wa2b3CzcE7YNBueMI1GGubV
08x2702UIiX8w2rKG3Vh3wfcOqurPswa2PqOUEEKdLyMeDRJ5ZTtrw7rgMrcE3s/6XGYvTMWTs2U
m2nY0S6pUWM34hcfdV5UP0yHVt0sds/6lMznWPbzYpO2rmcvGlS6+ofAr+Z5JyD+UXeYSlFX7Wjy
xGG+SkKQSaRw2d0E6/9lOTX9SbDlqh9gOT87U6tg8jlln7AD9FTp3F4x9X/i8L0PGpNIv9QcJDUt
0I+ZatTSR+dZFbZ0IlmsYXS+z6LzW+rwIvJkpLkkEc85Db97RpARoaURuCajvUnjVKRskQkgKXnx
DXKFWcw6cMBTpHu7/VqTBhiEKwdDNzAVawTkUqmMgv4pFzxpF7qGE1T9V0spJU9DZVoF8S5WVO23
fJaDzoZUObP0brYJ63ON5fVBTxcNMP1wOOZgcz7togdIt9Ud6D0jbwE9mDMaH0ONmxnnLaBri7TZ
n/R2KgRvRCKK+i/hZ90aXg3NSeegFmdwrvn7KYW6yOJQ5VLx07xyLoq4CL+vo/8RjbG4peQDC+FM
C0KIUlN54xeG4J11wjs8GWVGGmVKKNnLDCiC2fEoINOgq0ethGp1hsmAr4gcg/HFN16N95kR02/5
zUvfuKmuCvGtL2mUuBKwgLT2t95tEWlEO8CY6KLgYhA/3GCCIz2ua0mioq0zALXVGBvALifjDPyW
9/I1yvNPqjAw5ygciL0qc984OCAzLb2Bv1UgQ2pHNQODU4w2GfIT1yFF07E8R0hRfu5a2h7XA3mz
I0TBWHY8iUkK9zjZ5DiDoHD2u9+Y8C86fztCCsFIkBkHQkqk82QoyDaOWBKboSN72TsGA7IoheJu
HEOGmtPLPPqJJeSLd0xSahc30ckMDGxvctc3Aq14S7qhA/WrtlRZx/ji02ZMCULczCKPM3e3H5ta
auNuEUmhbiNxaQX9jZ9erdBOaIVUqeGNdaEGUB9rIH0kszenuYBrHeJS2ZgkpMlaxPxQStPqPaNV
iJCiIm6ZEZ9MRbRA9KgNrHT4H1cZugnvi5GWyztE2sGYFUrxy5N8Iv5pwr9Rl3ES91d0eP1ZYcvC
91qtz3Or2ZhvxF2ihuMmomHAYk9wsPiLlz4JoXB8YczMm923ugNt9JIu0e5zzjLODVfpPX0SOr7k
dQoS3g/t4RJVUHQOpsWC7z56KHLFMdRLbBWoMr5LDSRUfWnMCcLueV4RZWVRLfk1m6Ow0pDBI1Rg
/SKzE3tCIklmsXV+ECGV5aeSPP5hFpxG3rNu8HFQHBEah13O7Q71HDwieulvmDrAhGhISmq1SJ5A
8evZ5MvvbG+pnE9m1sE7sD2SJaq/WW15sq9w8GEygOHKaRtOTTp3885eQ5v7gEtMibtMVtCkA7sk
oBqzEfdpmE/VUrTbw1DPQeNkJQfpWQ/UmYJPdfhBexK3VqE/oN/Aw2yLGWjTZQIkfVwPGwJWR9u1
2tzQtZMI9gE/LZdIeC0Up01+uyV1AgiqoIu8XIDZqG6sXk2YJh1W/GQ/zf4v6Pe0cPpRk8jp5Fia
uo6Tmh1qsxkAUm4ogKSAqvKx/Ml0AClRgP606oCXck3+QIHVk569CtCZrf1MmNqCJXDOwe41Dbwq
junq4s0vCrTFrcOI8gNRjFFiyY1tCgNus8I4Ftj1Jth2zmxhEJQdQ52m/sR78fMHwvL8HRPCX/qL
N4aIQMxY4CDlX/mzuJQRcDh13S70dhuRp1m+07KBf3VKACtGi+3n6KiPAykBHtKMvWoo3HmF9DcC
NkDbd1FeUiW2dwTbHvo5mQNHsHu56BuvEiRAujpebIsYXIx5tca3SYgAXCrb5TuKSZhO0HbatBLX
oaEYF7Knp2HKyLKJ4+qHsEm1jS7QDFgbReJc8DeKbZdEgIn0TBQ0CyoZCmN4jeRZN3AJWmFMnCsv
nW09O3QzUdjs6PaHP3VM5YrWAdgsXyMUt03rHBDzGZHoLYn/dE99HpPeyVlaM7atfj+g+4skShYI
r44fUulNAmCB61UFA+YsDRDBolUjKGyge1eWq9zbHHodtDK6RimETpWjjDUx2H+AHSmKtSHuziDh
wKo4SIi4xMNHBSd/U8n4xZ5vwW+53pnGoTGc1xW/A1R8GkBPf9MdYO+yDujsJqJNRy8YbQ3JHLlD
j1H70dogA3jbdhdwf70AaxuNB0qjQZmenhKkpZxHU7rMk4AGqbprLnwBHfKv6EJbv34nYtEFqgHq
zlFtHxcHzd9AT8aaz2z4vWC/kY21/qQy2gI1X89/0My4JXtyknoPsVKQwkESA2f7RcK6Nf5QCztd
nWROJVXCm8tlIWHa1ihA0+IXpKU0IlwF6m+rftH56+BsTo5rPpMA4D5L+Lg0+CaEu6IjH0U1PERk
sYrkpMw0vX/cLOpwzgBTp7ce+i7JyLHmfAsz9EBAve+2z5LN3+is12yOt2QKIuyNiY5A6xwKyoAq
7wYm5lP33m/8qa+DAVez9GKx7dxSuZcwobJPB2Yk+UOaL7YHUlpjekr0f4AbBgf0xX9VOJJnsmYS
RGksSZoL7o3XWW+4lnoUFyOOug9QaH784oYtjntRw3criojzeWtxdvL2PDEbR8h+9EwiSQuBYnN+
95MFiGhUECVEvNcOt/ehMD0Obz3XU8FNmceDRDXapjQTWUboZM73sK/PFvKgAcagZjLuQ2WI4X12
zIcedMPkvI31BkaFNXL2YqjrOPOIDAdflzJoNxYJeQHb1PsjZQ4m4w+wj8/ahaWoKgUj02mF1FMJ
526NlD4R/uKEkfXswN406Jcxc8Tz1T15BKohQAuGPGDp15diZiozSs1/Vzx3fyd9DHpMzGRaVh/9
hzFDWv+RPzUXfBQFmCAfaVjQNL2KVf24E9q+y5pQpL6sDYHeiyx1b5njK/Ya2HHbYvcwhfua9ubT
K1wAIatk/biZNSVuQwAm2+PyV7wz/uY0kfulqpJ4Qk0jvDeb+tAPQSYX8BlRL8F2sUO17xgoDY5l
NYi5xhmaGx9rAcdu3MhXMsfrsWiRzyWbovXxnPb8igIy685Pyz6dmpghe4QQRnVN56VmS+qsgrCg
cQ9yEjSXyH98cYeYUsHpADsHce3KiX7luPjZbcYJd4swIXPqZeIMR6tYEOCEJ7qYlpfhTZMU9B1g
N0+MuVb6eyhDnVGjLCuqScqaW6WF3zqrPfi2th0JkfsIUV8AoiVbqGFztWKNzhkinVTIl0jnKOtu
DqkkHCuYwYdDuccbUjsZO6S8Je70i8B5zj2bICxjf7zDWrjGvms7cC0y1ODAMCNAL+oFDFX8a2Ei
5nuEE7yk8eeA9sYA0jchBk8R0ogHD0paCgwB6wlPxEEPR43shpT4splcNuM9dxFwhM4wUJeuj8M0
5+OCor+Um/O8eGnkPSpps+PFUTv7rOZDP+oHuLo9w532Q2Irh4roNq3VC7xtlzLDIippytyWx313
Zlz/qJBNfhEMvPoKm9MEKkIYZo7uBzXm0CeB5uAsomYlbbCKuZ+PqJ5AxV9Npb6y5+fS6kzT3iQs
Y51NmCHBZyDygdza/IuEermP42cnMZghlBPMx1vYqrP827MrBDWxaslUioTGytSHDd0nO6FkZOgZ
VdPUwS05OcZZOs/f345KxTXxup3DsHsWGhAlQtrW8+fRJ3LjYpA18Xwk2IlGbK2OdI88l2cHE8Gp
WpZb03dN700mrr89+LHNkBRlHHASw/cQa7JZCqzRTR/KRM8LXqKmznYS+zT7+8ySHehMAeyOAOt2
uEPL6ZiywACA361J2I2sfmw3guO/8jFsdQ1gGCsogBCvreIm7gYX1tVwfyUAE978wRMac3t8mETm
QGzQqo/iVIPGwA/dOAV1u1bcjoZPuwh+QtytZRrgdc05EryhXK8J+iUros+c6v7Iok84vxewsYas
Amt4hV2319VhE/ciWRmDpA6Q0oZBAyZ4dBuarWdcFy7ZTb1be/s5oY9LU3VUsu/qAc3If4NZS/V1
idZ83MdkWwUrkh7IoaF4+VfPMX4QkPyEECJZ+aVdDXVzZy2lPMEXomsCSubrYy1SU1vrXgImLthq
KSZPaH/LJts2nG0QPQu9lXbhWiKP/GulLlkVxNIRk/3J6aUSpzn2jJE7jIAikMg3aJmkfyd+vj/t
97i+tLK7KwkTQbYl6fOpjXOqMAhKYw1pmagWENgfdGlILgQ88Hh6XvbOQScXYClnr7naRc+rJFkv
dcDx7gXFLLZYvW8PNKF+4K+k5+LEPQDMVpA8KgERmitJhv/7nBnqiGAJuSjEyAlqiT+F5qvTUKtd
9KNkFj8RF3+pQgDQewrCEY59dxVAiTTcFi6z2B2/vUePn8doT94K4glQOCb9d+1FeCJ/5hdeOB5f
aFRAtwO2FOfRmtCBOEiXEEJTkY3r+dw6TU2WVxPRRERLTz04UxStFpnmpMH4/3GuMaD+K5CNZz7K
Ja8G76ctXKNfogIDVrg9HX0VLBaRgM01eJsdQCa0Szioz8IrEQRUwX84F2WHtNCzqfTBwcMRXQUp
wBjq7F8Tg8vSA2BvL+0i0XwS5aTCQVjZYfs00QJYqCkJxIQ/5hgy/e9cFW2ksBy8W1nTlu2Ye4TW
dW2StX148+6vYh7OxWBtW6q4ggWyFYiBBB6P/5rXFAK8x7Gasp9N60C7d6BLex1xitYKrC70z5f+
LOU4Jyg5w/SlcuIeSitTTT17fOqskfJQYnBTdMCQE54I0Jqei/po/7MyErXqd1OWWn+qnkYjm/H/
FupNJMaMtLf4/cZL3YJqZMRFDR1eHFq2YtpP/Eq6lKDG+ksoTdkgIVWTWTZrL/SCeXzm6ElJw9rM
m5C3z1EgiPRSxMOu36F8+f//FC/P8GUpbVLJt3/VWxQP8f4e908b3b7IgQbaFTHS2puRG6NMbl9f
qjunyBsrNOQkTnux6255PlwRFxTlk2rrVqogLGyukBPWwadnf7PG2LJTdlO1tpzGKM4uOklqB+jE
jlXpfpKUJtksmQBmR3jix9jGmymEpwnjbm4zb076G8TAFCCJYgggPSHpRU6OzZF2eYujdzzfdj/m
js7X3NWvaHWtoxT+ib3EfHRoCUloZOKY/44oa1JDjWpMjx8B0pIil/Ftp0XUs2YGPTyfnm3x3Wft
Lwk0/GFmrpIgeHnMbrmgmTuze0b4DeARKl3qKBktIOg/XFGwCRLORR56x2IygvHRmrpMUvGbuz4w
cF3MBJsdbWIkPCYh+GC3XqobVkzfbbOmys3mC4wZcWLW9aqNGnue8SXyke5ODijlhus2F8d4H13/
tGndLxVjcMgETdODxvJ+kAeEvPilAry6elawj/th2XcUSYHhWIXKHEXYCJa7TGJvooHPzpC8KDRP
cYA/B1Z6G+huvFuE02y3IHdXWqbDvf5T4QLgWw/CuoySbFMKYYInwvDnbWM1hyROVew/6xMmiFJt
OY3rxSCIvxmjibbrwjbsFCnJzxVTpMX2EBnYQa/6aEsBgLIxZ2UVHQiKnVv6ijVD1vfGbzbRI3CJ
DGEmy0qdDo0yJZrf9JnNhfmeHpm/zgXhqnnzyL7LEdzOLIpBRtlMtZpaNjHI4bqyjhqzQ0zSIa66
zjxnliGrpYY9ZDZEeYdOpoj43w99JqDXqNwHdt7inoz5SXEmiWLD92GEZ1VKZW7JOYXvvGtO68mN
QzPe1VrMW5ZkT6QxadqhNRiYbDqfqf89hT5XYVXjRkRkR1LINiWaUELgG1z4TmGR3YiP2fgRjOus
bhbqvjq00VE1TZXnU6Vnm3XRP+sdop3urtqJ4zh/1SHQkTSRBdJtT9yO8AwBtvPVLD8v658zTUUJ
kUppkLx0vBR4I8qaym+FkK0HFtqmM43jMnBA1Bh2B6vkthbncf3URvclY93nEkBNdMUQKybxd7x8
0ty8tzYIkOPcLnwkGutfDdfE2QcIkQsMf4mGJvC7R5kMHCdLsjvNkYZvst32JUl7w4pzShrimnEI
3MiDH9rkjwmX1q51I8GBF2BswiK8YtMHUCSapnKFZlc/owH2AT3nyhjum9ZUDTIUOBMyCinXq5QF
1L2ShU8ec6Ck643bAljMpkPH5+zLEvfc07LJepIMeyuyONgaHS2ROSAPfMizNxxtDrvZwPgn25qa
1qXFKlcOfAnofajR05+53EMrlaB0mMlGRLjNH/QPL3JL5yMWjhx567POivpIVkaGbzeXVW8DBjHy
laT0jgtllb/FlKMvPtwdeEPsNCzSw7f9XaFqw9ymRMtOifd/Kna+x7HMn0394R/+wrqZnBjrcgSq
ctmUS4s9FB2SSn5bbJQQ9xg6noK2nOoohi4A5si40r+c0A7e/vdGY7ohmRzKnWeztnxMx+L+PKbJ
nbatGHs3DLL8e/nUwzDiNQmdt/rNdxDv/6Z4uRNycZMpvARqx98+va480WaamBhsWAlqIuoBstoy
wCMzRchL4ZH7y0WAr8q9F/5jRuG9jKn4uBH+hR6cgSF+O2/GFQrAyoNPjIJX4leKW868o5vIAhWz
8dCJy3GRNJL18sdjbv9MHwA6irZR7/Ey0n+MfFJ2kCyenKJWK4oIhkxCW4t1tWDz1A5bJc/sIzst
gYIk4JJJs1AM5hNxrJMKQNs9AWSErzoxt9pd1Fu6sk0WAa9zpb1vpLirsN9enEjh0PSoB0zE5AnN
NgL+kpOPa3++bWiq6HPhO9W2fb4phzvuO1pRawAHqB+Ssbca2oMDNam5gj/WueZZCJWIEqKrfc91
JfT0heMmXMvPjiDFYfn7d7HpYGwUQLP6zUaeHC5lb2TlmDiCjOFJDoLl5xpIboG0cpWQrH+mRa0N
q59+N0bwHuT+dO8PZAqxJ8LwXlcjGL0eirgwV9gbp+P7Z0vx5AGjqHQ8otMWJWmhYuor5Igqupik
hughsshNsDGiz61OhJxKJRyF4iCLeXivfqozUAhtuori7xrMUq2C2dZDlNsiteYujY8XH+7ARUcL
lnFAlh4S5vJuZwPn5Lixm3gbDTyOZIHQMhib8IByTSKqeAN99zZmsnzdeKjbxPvDNKWQiNQe/XYz
/pGhCN/MtJxkOLiUBwWr5w3uBzjdfTzBoSqNhaB7Yn8Cp0jJ1YIkQVLXk78RpXXW9egugAtYFi8/
kHErn05hp82+Q2z4jsVmlz6GWT5EvegULZHmFsMW6oblbQTlBqEAzSpbTY0TRQUuGe3VhuVJCmnT
6stU9kB416wvECpCyJHqZRPWLCW+t5J4r0ia46gsbc9FDyArqKoXLEg+ZFPvC36JyGExYWR7OIjy
3AQgJ65rrG2BfAKWskO2G24svNinPZDX4TzFiqfAE4gurxiJb46kFeknochJFbGei6wwUsyQvG0S
+PL5zE4euta39y5SIrXJSeldFtMKRJPECKe9J0OW34/Yml7UR0QIm5wGS3i74Mq5EMYwryFVZnCA
uCWcC05iDQRRaZ6Te/7njyAuLiJSUm15bmgcj4nfrFHAdkO63WfOU0NqH698e+tnDAX6PG//gnfH
CjckM/IYYmUiAeSv77zXR+U17aUoHi5JEuV9cjcqxCOgDr/E9b1KMjue6LpYWc0YEqslmMp8WDWD
sjjDrKRqFbKOJYOnVBg3fy6FWCg/M5rnVrghbRXkjxpJrbFruG6l38QhVNmmY58OobW3EZwyrAnQ
wkZv4kbR7vbanmQkL0Y3BCkd9TsAOmAIbtPZ6oMRMOIHY+Cqrut00+fO43DmLD7MhkjIWOxgRbSD
S0dB/srzaYBZlLQdcNAktnhr5+YjEmreD+Y/hq3MRZ2xc+5Demf0AjQrquGY5IhULoTyLtS+XuPG
stmS4n4goQiYHwcxbZYR3zGy2+UICFTmdDYM6Wz8LAhCq2vdHq8m7qQa3DNQV+fDfZNnb2hv6EiB
Ai2A/XPTLXz2HFhau05RZq/xge2k3039Sg8BrF761rt/Hi7bVk2nHPDcVfTc4w1TbIxQ6BwPGAr1
2QToGCD5/biz4UcbFdHj0RKtLDPZ+qTtqx2t+9zzudGU33OfeePiMGlOQEKm5q7ED2Cvb6Qq1E/e
ldwNkIS21/HqZfVUf/0Cq/S4KB/Oa4FStWGYiRrK3S/ZaiqVsSMGR3OfvtgGdbfghTpw/1xjQlVL
41N2Xt8SMYSYYoD4dH7WZlh5xeG2J5mAz29agAtNHgWMk0bd7R9VpzfWEnOtcf5TrZbvwz7dux7D
wKK35WDLJnxoGAuww6tDcuVMEHvKxgCVfPipIV1Ia5OEpl6omZVuYfdL7LI1G6K7/gmIwWJlZIs6
6cSAaUP31TkEqHNloxWaDnRXFVnS7kKKMgLrGB4lwVZgRtn3sBZKNOSzGnOG/6++lTh58QsLve0o
PG6XZG15FGRb8tvC3G7bKtPCzV7/iueF6mch1OjQ6lONYbJ4RW8cbM2S73GBy/b778dvhGfqCBZJ
2ThxLI+f0vmu9nB7FSu1trULlND0VyXVAasF/k3djIE2XNsbvvaQUbOpexch8Vx6i6miVncZaxtY
KP3OvEPACDaP+2v+v/LHWsgBpsK9AIHgikquyUJTG73qmhaXKipn5C4lYm1/QXhSxRBBgMiNzaV3
iEtfJJvLsz+7mojBnJcr0DWGm7rbrGtz8L2vefXXXI0BcWporE39mW6qIq0v5e3UupBqIV+PWZZa
cWRxUpQaeVT1biFifmmMz5KV3M8abctoBJoy6frnQL5GCXpArJbReeTHXFsebMQNosdYzwLqyw5M
58lcFmE80CXr04vqIc4Hz85J+sG/HlLrrCfVcTj778PNSYtylB7Bue9pRaHJaPS4zrsgmHaNHfC3
VSKFTEtzM3B8CIIEnxXPcZOdS14SmJjL8FLaeoXsTDdPkCFka/sR0YX3i3N6Y7JxY/MWF6MnyT2y
AVe43yrxovVefL9zKxFYSxEmSuk+sXsO7Fmh3H+KDEaMn3oQjh6GuQsHjklNJehDJuofcaAPa0UB
5VIM7ewwcX6Ghj/rSJtpwRnwmyGwKPHeqtqZ1VBx+KLQNdhaiQHfawNfYffiSoduvNZUAmcK75CR
nI5Lc08l9j8iQABgoGas9rmS6BGLtENA947lEhQlymPFIl4EAiqx8u5FFF7mbMe3HDk0St7ZknP8
CkZs71v1s5N9zWLRKZkYD9Kg5hk70svgyNoXw5JOSIZUEJ5b5LHtm4egaj1AYVh/gNgDHZUG5zO9
d7HvSDzbKlf2YyE38wuTu+HvToCCvXbDd9gT5WkPZclINtAPCl+oA0IHpH1RovWkhKpSDbnCip4F
QPO3ttTr05rCAijYqkwjOcjMS48ypkpLt61MqHp1rSYJmfr3V8KvFclFjq4ox84VaL7bnchyevIg
AEH80hUPjnT1TIBopxjEdobZOIBHPizKMQ+PNz/zUVYlIvA85oG2LV1gF/eKBU31HnHhXM2ziadd
Uj2RVz5IlwsEbnQI9ZUrQgOvPxAh5TXVOd2mKqX507/IeHzcCuRabMZj34Z59ppAui5sxVLU6vyU
1WVGgB2vaKBjgOzkepl9QoHO/ct/+R92QcgObi5yxImFRIxoM4TehBlnt2f/hWslOO+pZRw4B+Is
PsHjLeNtF4sSM98dV7yDJeE6aCgVaIF5U9si3YeanIf8SR8oTkeGqvhL3VRPb+qtfwmQHM5m7P/Y
A2nRtN9P0OYSrJhAooWqx28lvSBqM+4+Xlr+iNmFLclyQTIvlkuD1Duo/gcZTQKUR4Ik6zBkpFXR
ukNZwkF48i9piT/H1WSMOjD2eYyFkbDkz6Hfgf5LwgqPMhLI4hgvPaNzCc0JXJmM4smtuKxO/z9C
TiZf13OxlxQ+uoEDpPbf+S5A3EDk906xNuV0fg+YADfVyTnVb47b5CuEiqNyDbcljrX+Ybpj3M/g
y+WIRy5wwbcg1KegmChYZzQgivXCPq6xGsJ76j+FXlPfGpGWu1ZBbggM/awqp/puj5qWL3h41hEH
vTgrwbb9Rdx02vUN0/3tRecL2k03BS7yX1ACSBgmTdLSeTXAK/0Wj3mtAM7fnYqAxbFkxricXd+0
lEgWk77KfOhHa79hY2gvnZ4lKeEPmE3urio0wcHaJ132eXQUiOTMhHjLdr3L5SihR3Lr7NEFFzgv
4vZKTfsA2Aw9ogHDzN+MKvALIAT3GgPSXoliUetdeCKFpu6mfcjmXESHyMMaV0BIZ1WFq19GujiL
y5NpvUCyNne1TX8mW34rJpRvVGkGGeVnWxbzoTop1VICWkeFr4bSxOytpMhmlyJX2YkdYh+UsgVn
ZuIYaGe+jfrZosS/iEtjPPwPjIEok+2QRXK6DgZ+tk7B3ejNajwMqZbP/RwfkCDCz4SghTQ03BYU
6ZG2HPxneZ61eKy2ToXlrVaJXu01Rwe1BlupUJrAN+VYoDq/uIbOFeaS2l5ZN6Kfm6Z8p1W329dj
3iwyTAxrmsHmO2/lPI/5z/5yrB95mOlArcGruTJKo38RSCUKTRY1tEKlcph5YFGuUpd+YidraiUK
MrDX2ryvVqiMxJeyxr4IcDQvcK9f+KhB6RbRC/bkzpW0ymAvghpkem2A/p8/P1QJ+o5vWs6h9q6f
gLIEPU25plTURt8unUnJ5///znJbikSy5SvJMFTJ8bQCFdux+Bz12KpJ0RMLbVKj3fGje5H5xACK
9T95SKVeZ2aSoh87qGX9GsFBMk2l7bK80FxYMYi5VDet3z4us9S5ojOg/I8437oFJ5i18xZtq3b9
pT78Yr5Ll1flRi4Zyy0htwwcERbmhKWfUvKQJyotz3FFgXCe6612DgYbPr5MKJ3f8EoHq/+az//z
sC80nol+QHuYT9DmgiSod6OInkvuv7p5mEpGio7ZPQeqSTlu0Qk7VIRzre/62Sng1rfbU3Tr4OZo
p/P73fP0dKJ9X81hpasiXsV5qfgXI3DIn0dwtVoc5NRhnTU32Xbu74L/Ng3u3KuJKZk3htlbCzAG
VXiXxQpx9ZLd8nwrIE6yGoQ4ah4SSuU8OhecjXFW1jd8WeiUNZ6MPoXiAtUdUWnMS3DXtJASiEIi
7olPUWbrtJ+UufD59XOfCgBLJn/ZR0wfR8tvptTgq40necSoqeLVpWGx0X5QZzt4LKN8Yv7rq59Z
rgacx4cPZNFDphw2n9TZQDwd5PlGRecjSoF418ojMuJppEllSXAT6ZMt979zOFqSG/FD646LKoHg
KG01EoSIRUJJ29r9nulFwKpCS/0mANgATDrr/JF61XZpsEToZqogh56YG00kAbmDxItQU/+Lk+R+
mlMOOjpaNU1m3r0hiQOYhKGTR6j/CNF6O5b8hxJmR3q2A4GWgR2l5SZP0dQ7D/58pG+At/C515u8
nUXV7m5rccnZUYejtgelduTJX2+kWV9uKRZeobuy2A6rByB+81F381xggrNAche8vhExhnt0v+Iy
aEw/6i6L8YJoKTuTsI/BRYKeVXmHIle4RC0GEuERzKEuaAU8LStAXRPRqL9dGmLvk2MnoMFefo/O
5LVSBVHEV25uwQbxDqQ5n/s+DX5zBYasJnS+geh0quoHQXRMrTnkhyXI1Gdu6uJefZGe5VeEgg55
fOAqsS3eyJdezZVafDQloeihy7HnaVykb2fqxB/KCuaPA2thmSgO5z6MEPcBaTPP3ARGtnPIibJH
ypdx60HHObKV3F7KUADElv+7TT/0yVfscSvVqCLNcwNkk5WDfwTufLCEWR2uPy6hMOUmxcxjT3l7
eIUgZp7TI0vupOdZ6z0bpbV/UX+PDRg3HfuKXdSExnwPSZ1aTNy4jmPecpDiVFLoqNRbmDKAtEUW
fj4P3UQJULNtWMEIjgEnsXnlMZ+kWRir9jyu3rAi6R1bALGavAzWoAGvWEMAmdRaNyfDp0qC+U7m
QtHZWSu5lq9TpA+ubaQUyfYMoS04TiTqCrk4xuxx/+6eFov1Q9ozXPyEHxntfNapCmmh54Caugl5
h4/NDaYLlmcAWK9gZDDxvmBTenBZYNSMhVs9NmylwY3yS5NOWywspOkZLXLSiraTSxbbaMvfu682
F42wi1o9E9U3K3DFL1jiqUiu987tfjRw2Acw7cxowiGA/Jth8H/wLpsYq2Hs7WuPkKeakB6CkQzD
qW3Fhf2ij+HFgkqhFEzdh1T9/2FYp+efx9Ct0WhvrGXbj7/3bbyKs/Dv7TwIrwDRdgSjbsqpzA/T
RYgVYRROL1H/dApSAZ2vj7Dr+8rs8Ty+I7n6gRwv1tlFuUH8b3DsJUwwF51pghPmmoh+rsX6FZQ3
5O8Wr/1zz/NNJLrjXI2qnRMN4UBorwn3Nz860xHF2giwpdvITstZFGWHHsM9PPkE3qcTLWnVrojA
UDUHhtT4rS5dN+6nlVMzu90vwyrYFCao8VqX3ft0BbOwJ9DEf4KRAMiRyg1uFJSWjJHgKZ4ibExU
rmLL0hXBsUN3SFZ3slpWoaMw38RiQmx3DW+jzNTtVVDHvrifECVxY6ReAeZqFkykdE1PRGDmjEn/
F2CikVgQWZHS4X15oSLMTFib9ifjX/bVZX4tCziAy2+Z+uV80L3zaegSKzerVodJ3f4q7NCow0vK
8sd9eQa7FynAT5WgqGCIRHyrKlInO/6FArSEDM3bWYI09ad2Fn6UrV5JfQNPHCrRxfDTKFTGQO4D
FKmAvCLiyszXXGZfZuoKd6nNz4yXd3LVZHYFJ+CllRUbIgEwnvcmRaKvlIISvCUHC8gY/bY08WXw
1gtqzzbFiK5Yezx71kfJ2pSEGUSl/zUoWUZm025wUW7eVSGTAx93ViABdcTQ7+waFUJxGSYT1G7R
YA0rBKz3u77rBrdlXEE5mD+t0ZQl3lf1M2AOqBTn0X6VUq462S7iWKx+w3G7G63WKl+7hBfBsgwJ
unhFbUxCtGLdXfTgOIGftsA6nhI2Zizyqt17woL3EyHAMP/L/So+ZuCGRyUxd4Gt0w2hYq9Elua7
gXgRJjQ8nN3X0VQVbJrwcexVg14LInV2PHAG05w2haF6KDbHZc0VAz3Cuc9D2p/5824RwJTMToPN
AgBvwYUxoHG4UWtbuqNnSioAyS1qvMViN9R8PkzTfNVpPyU7ENX9Gnn1BQ6lf7U19sBltTOySaNN
1Q/Bd2xUfxNNgQmc4+uxtxlRkwWQKBqRx2awla4reya9L5XUiQ/SuNDPp9cA2uu1b8w81BaNYEEU
p2Gcxh7nmbCnZKH9ysd5stxHbGYS1FREE1QdYqW047uTpu34qVPGaF8Grv7kwdyvnmJtfjubuGJD
YnFaydNhMxG0+P/cf7QAOZrgxnfLCfcqaQ1zOfPGowaGyXxaYyTJDvfxfvLd9Ma2MU+smKbZQCGn
RFIXTKGhQMuh88gI2sIg9SFokiZV8flnC7RApxMC90MtiGhGE4U7g+b5PDAr/hxppYqGpReEQQ3H
J2wCsJYD1fbJMALdUlbvaGZ3wKq/zw+3VCbkrCR2G25xENMNXgBArUDAEnI/EwZkd9Mwx8yajMuv
wrd2DIDloj/iaufc9qk7MWt3/NnufXM+dsFGjf5EUt1lNVAk2yAF0qHH40KXNq09DjYItGs/K8G1
6/MjUMXRJk2qEZZNMGzbkErPui6ZiNJd+W4DV6691/Di442anJEQFVJ2nK9fNwftuyg8ZQuRNyDP
+O2VHgHJVnFNFSOn36C93YuVfW2vM2ByIYawAe2+qyj2nZMrwj38VBCY9+u5rnoW7meshAYhlMmJ
Vo9FVsZSWEcRMyjBVrqtqfEHB2F/mwT/B2ajOHbJ9WzWUPanZDmydVkUoHGYSJgJH5YDjgneNwhy
ZmV1zMdYIfVeVgpGKft9JVEHmv71q+DPw3TQYZKZ7u7205IBBTeiDslsj7reaEBjhEnpGm13pG6Q
2eYIbDtGaKe84+FxzeZMuXLkp2MsO3BMzYZcWHPgXr5d0PErWPxe8g08P4kUkgH1cD7eawa7/07d
9BMuym3WN4HGr/yl2OM7H/HbBDK66P70TKssq1nrj7Z7irIu16jJzCmt0jZn2Z5akzX+ADVtCr5M
NgLqMm8lmsCX+O2M3zaDMNEU+qkBwm5n5YGH3yU39tE2/l0XZ5wmEQ/QEB3jT+qLolqGBWuEARgg
MDfbbPU3QPvY9ZQnsLzfcqwXbNRTlgqJUK/WLjmW6JUQDktdl6riHyhBFIiW9tcwyjv4zCLy5eK1
jj323Hf8XuJtVqpjIovl2tKpAJn+OncwnB9zU5JP7wv4YHQMVeOljGoVg94+1MKrxs/n7rA8/A8s
O6tJ8I8RwRDRcLCuSn/PprVSBx5sIgPfnaXpzVaagtfvBJurIKXRUHHlT9Uwjvz//7an0UqgLGeG
mMiQLjZeNKHFT6tuulnHIy7rZisxoFYNMGg677Ax29Yapq/YJlLVHl+KQ/2D3yNKq7mFCSvGb6hL
em8Hmwh7Fe9c2AViFbkIZcXTm/K5CQvyTes1u6N93FCQ0GBq5Xtwc1dgXY8oKn0c3GuLfULr0kW5
+0JMiYjAihxx4UW3xz6sN6uzbtOzi7I3BvDbiKFKo80I+VsQhbJLcyPkoi9A3Sd3DKhZuCQiFREo
yAha8WO4uMFhCcmFGJmmqZcmlirfqRUnH5b7Fe1rzPRchfh0kEIzOY6cDP3M4V0VaRwdKlvraSzb
OLV6sJszXr4dFx+9jGK2uPU52Mbbrq3TEgcShcbAI2ia4mzk8Dq+yGZNsUcPqh4WUXhBNJq6rIlg
CM0KoYX6QyLtHmdwEs7ttvsFBXwEK5lPjKmsJrU8ayBceXQ1TnYd/RF7EA4eajF86dtbGbqJUv+T
qjxBidFYvKMottD9nd9g7vcRu+smXHuqAk3dpjb7Q65kRaoafRbuEaTiWJ9nidQTu2hNPIyLoHcB
v4j84/omYRjiYjQ4cEskRJ4IlRl0+xbyk6o5CsGbu05fIEtZn+dz526o6YLAk/d08Ora7ut+QGhg
pIk105t/P2r1/dpRp1ODXnUcxNDJdsvTfKj7+97PKH0+IyJ9BX1v7qoaGAgDEVR0mSf90AQ8lP2e
5XipbjsXUMqjJwb0KT4jmEk+YUEWR1aNmhbPl3Wle8o4Ye9JKvSAQQaIzm0J5K2SeZP+p2VbI0Bu
+RB0EzplFL49wylUaPrk/eFh5gy7LTDsfaHg3v9CgHz2uy78etsMMt8VSr4t59IZBytOL0Cepj4k
8FeOAHJvPaB2zn6GvwxjrD7jjDRcSdQwcvxJp4wirpupmJb0wUojrydrA2xG9T3KjcPoWMSdn4uU
kOU6xk2r9j6/KDfsGDi3ERFsri7yM6uamT0kchtDduMAE7dY/XvzjXo0cMa6KXXV3bOzN9sut4z6
1cCLwhGwJzB1qYs6sSHV8JA8OzuKZFoYRTL6JabaDsPvwvBfyy2i8SxoGcm4+0LStpM7pk8GGIWj
+mKYPrZowEAWe8XWzaj8Q6Vi+yM/zzGl0HWJCkUqL09buQBvZPx8MaqdIVGDT+0TAskOJZU2hkXa
hoWaUhehLlX4SDyfmzwWOuNwjtWZ+uMnDP54gWLtuxoHVa93ZUU3k6hsQuTwc7U3rA2Jy6tzfidz
6NZzxz9E0I/fz7NP/eL6z72LeukHc+sDSVSb6M5pE9grxE11kDg9a4omAcpqZQyj7rWmsYPIekGM
HlWv2H7YkZTbxVDiN7rysUOn+z5QUq4Mz9ciej0e9ghhAYOI+UhSmtgrAnCyUi7Z8r7aNqSdOXMU
pTC+cMzOreCfYK7ySBStuleEgXVfD8w7P+ulfsunDLBxSdexHFbdDgBsxS7q5Qpg9kqroDbQ+Wlb
MX6pRNfPxSyS4hXCGu1dHp0PAW6LVHg7uYNzzvTHfzATZa77mmcqhgi3oW4JSLxbI1QQsR19q/3Z
OaIKLSFoT6SOzxYbPh8fLkHS2zxUNd1lRMG5zAG458Bn9+aMfgkGKPq7qyqpy8V9q4jGADDRVWDP
U6et33W3uJpMfrLFRWYoE9BkdDi+r+2xLuNFowLYB+pfacm30esvsgxDEJVt83DCNWrrx4QwP3Te
CsZ+Aaq0Y6Jacbl0gVegsfAKRjIWaYNFgm4QSdzG1urxBb6yAVEUkaM9QP+U6ZpkCdTSP3u2dAqG
E3jV74GDvFzQ53nPVMmullRUh5gdT0rqDtkG/n67Uo215ZLfnxlTTiyeRTNcg66nRtvPBa6WyNkF
5qrhyH0tidnqIEKyQGjZjaIFY4Y+Z7uQ8w7JYC1lp1d+yzAk9N5oX2n7qCctVznu4F7ETrfeYtqj
VpsXoJivrw+P6rxUUTHjB371aDZ+Wa9UsgXUCVQ8NY17lRGepLfhawza2yxcfSJae83scnJXr2Ab
RMGF8/tP6FprIxbAMyGG4kQMHBoHR6YGbFaYQSuqN9l3ywg7eJibWFJ4AvgfADkSFsmkDbj4opuN
HZaDFT6gcpTrTmKzsvbBLTVq3hscRNwZP9xuxeCrzmRUlEi3l6o11ANNPJPuXr2GoFV7NVaoQEmf
fnU+FH6pa/ntABDUYwguAMl5tyXGxok/DhUmSyBBVeqPWMNgJ7X6EjDzqKGee6Ma1mq/AqM64LeP
/aDt/xgduX2vnKRjvckUMomdtW1mYhOm0S3RUfz/ki103g65PVRpMmE1VW8ua1MTQ5ibo+OgES2Y
U/II5NFRl53abI6qauW9tXuk1PrEkZqJ9i71GpGeoSC894TAM3rchVhRq2EFtJZuu1Rs2F+s1M5N
IVnM/xvAYjrU76jGn/SNip73+tM/Wh+X/d2/coiajUCcQoVKKa1EUtB1/WLdIYw/ITDUReU4p7XC
53sEzdrnn5Ox7ST2pI3cqCuEjjRHSKFYNyLnR/lyGszTF55hafkbpn2MInZC+GPCqidPMCD/TFPt
wNRfPRA3x/xAszgycOptYIS+H0XgqETLFNnfA2rhgRVFTRA+0eVNYTRc0HT2dhbzmEYedJ03Hyl9
quyRIqSgaect1mfGolvJr8c+0DBmbbyA6YIFf7ximhcjXlzR8KPL7eS6h9gQJJLPZX656wD6YV59
2QEaj1dR3DQkquecBxR+rrPG+omVZw37x8xz+RzmzC8wXnyx51a/xWjFfq5U6WH1/Q4La+Q4olcy
lN4+iiOGvDi60n6kBvvfrsx70jJOzQ2pFDoWhpChLWk1oLr4fX5YjrnYTvKm6Mr83DW9Km7ROD0U
NC1WXbbvRFOjcz/BT5a1D7mOtXoYRjvlh7pfYU3j8MdflgY0Kda5LWj432nD1+d+YMncgWeFz/I0
lFb8OdyPhZ2nswlyrck6SOvkdsry2fPQuE1SNM4lWMOsUjMyHff6l0hdc1XgLgqPCquY12fQkUq9
+NsAyoRMxKVJhbBkj6qrGV2hS34GC8YbbDcOBu/rOMoSbtDVmDR40vVsjv+zG/OYANLGPf17n7FG
5bPNlatmRV2KJ9H9dDtHYokVrsDEJrKjC68hRMDoeOdVVIhVGyvRpkD8cZJdeUxCvtoqm3Gipyc+
kOD3LAx+WIV2otfe4xfjHtpFaJnt6AncPjGQ8JlmjVNGlhM2/idbHZCezBmS+Mx9fT776RCO6zvE
ac43Yu0gKB4ZB1l+EHhosq1yAPrVwDqZgK394em2eMZ0JVvVx8+h6YL921IRvgwM//h14hqV8EMm
MP7DqXis/f0hTQkm0NVB4gIHJCHv2WAiT+07WWDofqtxsFyZ5jqN1CZ/EdhgBYNV0j7ntqHinwKG
Z+j/1N9vvf6fdtg/B16AgGh8Hc4hKdNMbtNkvUjmAv/t4QV43cYpQYDX/r+XYIEXR5LEWI5EnaRc
xZVw1ldo0VpkQYxUa9FVGgd5m5EiSRRgsDgTyoidPuIRt/qI0YD/xU0z9HA+rnx6vGVFm6YeJBRz
QLT5BoJO9dS+uK3KCigVrSO0EY1GTcv5rRTrkbAOSlcjGEfoX9s12aqNCVKdbc/s/hkwr5uEOXuA
G3SSSEt0ZDTBhQpjvucNORXcHD0u24PsWJbKgbJfuPtKzu0D81coIiO97VgDsmcmHcu387nXWzLX
0RSS8lM8fOXZfe/oy4jESCVf6CmlLrigcNennaUhGU9k9fqLFX5tOgWouAwb4arUAaWAv/pIl5JV
gxMx0EhLeUYk/DO1FDgGb5jlghj89h0kwt6k7BtXspqU9i836mDmqGYzZL8TcrTk5KN1G263ZkLM
RoOReRCLNfOh0nn/G/Huj09r61NugW9Z+ZgiCP41YlBrAOzGhsTFXx7HhVhWTYIenpTVxwf2lVLL
EJMQgZTb5sbj7Hyt5ORQia1q69eY+bglCaoAD4i8F3tzHciqzvm283qj3HtHSQhQFn9sfABevali
llMPfxkSqWXFRJEFKrfTCCN9r+wo0EGX7PyWfNRQuenhR1Dht2VEtFZLF8z4N3Y6NXyaXZ89BNBB
bzWjBjlZQ867PViKCn4gW1g1Xir+D7EbazZ3qNetlU1oz75knj0JlLCg17wU+GsbroJv4cGTvx4R
uJVkLE29T2U75VEF+u8g6EiGX5VFJVk7ASHCuIIHtC9BHBrgpFDp4aNTS1ekysKMKA9NFeMhBX9y
epTXtnwVoLdSlD9sVYtK/je/Bn6pqOh9UZh5InElm5Z8yfje8DoN9Se9M4AZxOW8jlkWwWViHJHT
426+YS11dLpbYs0+tuiQCjoum+WRdNHavJ9cHFWLh70X4F3VZsB+uy3geWZiHHNpCeg1Es9oT0lC
MwVnT9Qwv2kUhRuaqZwHRR2SrJD1HSB6R6sZE5pfq2ifby6Eih8ID2rT4rCbfMHSyG4fAVt2IBvb
AluZ9QzuDzbQdekFVReCBn6Yoa3BqIeAoM0kIlgUx1z4bs2lR0sP3I2JM9QLbsMujxWLAy6T1+Dn
ZPq4DJOZFBnmJ04HaC74OD17hm86i4LWzxteFkUxrp6td8BI1YjQQeeHPN/lu2jhIzPssU3dQhmO
pTyxNcMIf7ihOk6zlzvgMJM0vsX5WtcYwJVIt8K+M3LzAcZaSOdedK/pJz1cYCLkYzvxi2k/Ht1m
HOsRS2Xtn4+ZmfM03CXmj3gywBZR14c3rBjOlBYxGwjP7HQPTwx5OorsIF+shUly0C7q8kmKNxUJ
VqKCKt2B+AjhrRO9qjO3UCVF+Q9UZdxVSOqaSaE84fZxta5tGpNJ/6GytEJ6/4mK/5pfCtsiCyeP
9HxyxcjlLlxAFdLkZfgR2aQlINsbgQ5L45bfXa2+7HU+4biVa8c1haT7PGVyVA02qhIBS0ElqSAP
MLOTukdiqcb2qqq4Zx+3G0kHu+EYsWKdRMLnI/t2iu3gCFBknZ2jwiCR38ENbDiaT+dffHgRSjsF
A3ogbAY5kTGlgwzBn4mxMKd99cg0ljab+OSb05R9SAhvM50e5vsc1Cb7XbfhBM/SvSHmmDtLVmn2
/4v/Ka9eivSzmvg7PcYg/Ag8PaVTRaZaisbHv6lxBTdoaansgJDHozWUGyJxHZgJz6WXPWTuejPP
pR9+8A+xnLJ0z2kT0Dk9OBuduR0Ftzx98sYj0ZYW1CnI4Ah9eUAeCqR38EBw4iOCwQHzD67g1jT1
tba71ICPeCp15Z/YN6L/wCazjtCoGJwNiWi66QY61sWmZUy43s0vSYRi3Anyx2FeDK/ldXUA/nU+
7zP6Y+a7TzIuxPOYWWqw9dLa2LAe1ocObMxlARqsCXUiwM10nPEBhWlXKgroLMPrdYqi+7ocOaMy
G0LI8baKyvhNb+THCTtErjBNtQdqCm/OYKkqPnCoKQw/YnZeUVCPnpP8qcQlYcKT7VyJpTKXTx0w
lNpnPVlmm6ojI6ez7Vx/K1X/ok7CnvD0zV807Ctjj5LnDIReK08lTjIlS/9x2x1YUZ64TM6ojypc
3zd6BcAPVDfFHawNFRN4Y6K++AyL8mjlRFG863fe25Xl5wL8JUalYDHaoLr3TF5znmKCyE9X32al
zefu5JTh/29eIQr9jaqtCqwc+oxJsSU5Uf36iJ7Pa/uuHFXgdkWMZZl7CovGFWrLVrjl5JTUaj+p
aAgQ7fD09tbATMauLxLIFxKUb0PmXJGtgMxjisD/3JfaEkxGbOE6eT63/gVn9PWdcrbeRRA/LCO1
t6EUiCeUatxt8Nze+CGUQx49MMi7xueZDCiMTK0h1+wuti9oxrZZxliquVLQh8zTwlfg3BM52NVN
42Hw42AH4/KgHSIgZU26YDqpn2XoUiq+EQ9gSMgsGMeqCcx35rwzVfVKWAANls1mqM2W2Y74YDPL
E4JRr9t8xkGhxQPjGpOSHHePuvEffH6i4VdO7rr3sq8nY1aFGkIewmRClbeuMUS8UHj9TOzfjqGi
OB3dPEcOjN3BgRDZfhSRLXUFGiSdePWhztVD7XN6KewakpzGX5+Q77QgnOks3McuuN6GPbB/aH3w
1oz5aZfgN41tYXSn4F8WG+f1o1fVXJDEsFG8BFHdOfQTxSKNNGgWN925SHA+U/RXHelQzxuCzeBM
WTPz+5a/gr0BERQEG8tKbWFg2jZe/gxaSqGmclfZct5oWhObZATLEkQ4K+p5l7+H+3cbhyvM9q6q
tc0r5yXOxQU5fg2xDkJSp21J5ynvJn8vSdpIjHNVGOzTC81yuGTBgOQcNzEJtca+IoXCWkLdkRK5
5kesFCjjfLOM1LFji/4N8xK8ru81HRlDFC/ti7M0AHMCy+wQwfE3Low9lRBZe+qTqEcaKmMEydWM
pFs3vsDjCAQZRFDuflYiSRbM3k0hRH2BBkoVKjccmseub05uo5uv3g//XpPulK+Pxw5f+ZnVcnQf
NuAZ1HF9MUVwgNYc/plwVJmCmw6PVAbGAysDJeHnCj855mXHqonWkoLegd/nhLcOzrppzeYWb/hN
NQUjYKt/f2SK87CC7OJ0iR4e/eGyiN/fsA9nvU3zXa8Zk2GLs2yXRrUxcgDW4/YHiVY8/ukgW9kc
Inx16g2tCXZFtx5urgNXLwzh8F7noN0Pvdslrwo/R7+5aqGsER50xAKyDoRAGKpd4svcl0n/e3kp
wWVYaSFWaSXcMj4g2rOGHAxpls/Cg38wyp5WWkWCFRqMC6dZg9r/i0AjIZ6lCeJ7pQk1qi5xFvfA
tQ58hNg8EHGUwcERaWAXKHhkS26WNaeKP1icz0CJQUsGmfTpvsbwWtFVX62QtZzpRpo/61WZDCwY
/0KlhCqdbm59laP9EM4F3nuo6gxaXmagW/lK6I1z+FWJSVM/+sgu2OvQU+leQrQEOsPorOsifov9
rx37B9gllRuvy829uJpo8ixbnEGbEd8Fx90ldwL328Nq6mVISaKjXnO+kzL1YhFTNPdUF1uH7RO/
jISfZ0cZWfDTVKOMqKSkWHRJRHrzW0u/Mpr1aHAj7Xs7j2DH2LIK49WnSYQST4+of+lbhJ1SNF9+
NxjijDbHLD3XhfwPDIevcODdm1SALvLw/UXWvthrnI9SN1qXk6XgqUbLPYpmDjmq6S8aKaC3YYpd
pc46uUbxSYlD/hYeHZ3vyFvrHu/rhcO9lGF9/9BGI6dxT3fFHCpibhIi5Hhpr1i0T9qGTU5Ih63E
rp4xOVqxHZVIIMrF7dTxDVBTPAAFk8srQVXSd5JPTZ62Weoj0Xqjv6moSnDljClVtgM0R/LhnfT0
4txWpvmvbiGCaWK1L8/aWt5toGuVJwXj1bqBia2zJVkXxBRAeyGYj28FRHQRsjTFP2iTMs61Ncby
PNxy+0SrjGSbf6WbQFeYa0w5F19LdKcqI3S509nF8zKnDcyPASVdkIBmSjuAQhaJKJK7JFWVunNE
QhtBrOaSQR5xdIdoS+NkzOfWryi8MvZjIEmJ93ZWV2Hpp6H8UYg+sTkyLOJ9OgbV4EaaTgyOX6ok
mQE6YOBsMHJbN2U+G45w5ipKmPVAsxs+Gloa89b8WVBau3x9Tj0c+wHswNFZ8fuRia4CEtPHFz/h
gadYG1Te4d8wMlV88EZBU6kMYNM909PdJi6AZkv3boxFN83G1U5IK8LTBpcsoaO3Dv8x9KJAp5F+
zmwVW+GTzzmQ+fgXrMpYO0LXGzo3lH1dM9vYDxcdbl/zHVSSjxWEiveD464gzJ7xmDglQfQJPQ7J
Yr/MwwyAdIvaMI/TZjUzoDUPso7ibFQiHdEwYCQhcTBMcNGmE5BKsV83Q+TzQxSSedgHNpP4ZGvX
Zautg1+VVcDpVGwnbMUnwLqpHthvVOlSdWaK2ihCGRtvx3A+951jt7jo9wJUeoMEHNH9ewgPtmxG
Ly+MDTeyQAkRAFQYDQiiwl2yXB/sZhb00kOqbJEUxntuLrpV6nV/JOR4lFNU+zk7ilEPNQpxFUYu
9ZkMHvZR1Mzbu1KtI7Xqp17aLsaR1wpdnd0fvOkdrn/U7PYgJR264xfRBnCjr+Lpw2noegG79CVW
L+nDTDJFD+sOGHNb61A81eJOCbLy/07C3UIeq4Q58p8bUZCeunX+K5PPMtPmmyC8qWGpHyx3u+9l
zOPOcCE4fdDtRedRt0slf5UAFQSPCBI0IBrxFOD/0hVmwr8BEZVZao2b44MfXwOP4zNYOW7TpWze
egfaofjBRWNvKn/Is8Yd8jpVYGOGN5vei+47HVqKhNHA/W1b0gtc0dTxEB/Wqt+H+KNzh8oRC19c
whBHqbPXIqZY/pW5FuQ763WNDmkOE6r37O4StJAWiLtlzpXsIk/Afz5XPB5U2djVxFYi3RuLLDTx
fS0W9cD0tV36In+nvg9AwuV+v2+Fu2GIsrZWNa1+UY6bRZ2IaLwsGru+DUD+SZueBfQ9x8vYTL55
0RaCH5v1HvkiC3u57nsYOmwmM/wK2SiBZ/WbmmB+jktNJfHkaGsCxXqZiOdgQQ8+a7n2o2aTFLBX
nkRAKAmMaGD1qRABkZH621kAY/5oVqWWAGkutDfaP4ejvxyKxegFsTJhxyFCi+S0IzsIwAx+Aeu4
s1vgAHmY3PeJf7Y6px+Rh+0ZiBWFv85se3+i4p8d+qWhABEpDisvGEtJhK+CjSf05+RD/z25ZrSb
Thp26Itw+ms5Wut3ze4Y3eCsmU3pC5CH9g2igpFt7IZM0TOPbwFDxdrJllZCx+685dB1rf0NcfSj
aVEpyp9cg+jRqM3Hvu/MzZI+9LdvLOurwztAooS8ia5fUR1x7SVEdrjL2E7l4Poipk48K/9SKyfl
3P13oKSQLoU5YyfTNs4HURJnjoD7fJ0hSVtVMraSvLj+Q6pNPec4qxnA10soEfjRipr9hHpLG+JX
bRJQs0Cy7ZfSVFEi+TKpd0PEw9V5a6kpHp1AI26qfHyKB1Bby+g34F/7lSJrPX85bFZce5Ozb/2D
TLEqtOmh8qg8Ms6eH6gK2hqNhN5RYO9N1WbgGSzbYBv9kW4suvg239o3DSBW9JmqAIkMs6QTqgpS
m9vLzbcSP0whZf1B5p8DI7gQERHaMK6lBrHdp8fSSzaie5hS2E3dSM44Z+x5AAK2Ixamcykg3O2a
G9M1Hb55O0HTHWmVZ2R59ViBF8iakIg/8nu2kH9+wJydSaPhxl1s4oodR0FkvODVioJN2fJROEOe
PYORe7gu3DSuRWXvAxFGAFWf/+L90HYWfCUTuN018qV66i57LotIl6wQ3FTmihDUw6npEW8rfhd4
hY7VHBL4hOYe2NAoeeCfrcxDNwZIkf7sCSR7ed+d81djOY85gWrKFy3zPVEkkzOf0uZ6Q78TN7rT
yxrWgceccKUaE9T1YklYLOCFHwEfN0XUMGcOMAuaUq145rbG8izsc+is4sgBdh8cYmKntJdNFGBg
O+lSB/dzQubCmLIob2kU3zVNDG5Zc1foRORJlI0/1BRjYfcVkpTAfK3uiiNeswu/o0Va4Qf5sMkx
WRuKrIvAs4OLzh1B8IEA+JBQnBo5n+4eL65yl7nHy/0kfdPRJzaqqB9gwcAyM6Wd6/TulWaQvK1R
pF5gGbmBmjpQlmkOX0m+yePydzRGZJm2nP3ca8zYbzsiuCrNz1iEgmDAmEm7XEir33EywRf8l2xR
vSzMHnSCRa9euNj9c+STgWkDu60iBrrgjNVIGpHOe9b7UVy1Wddan6uUIaopHmbx1nGUCX1qMGjo
xSif9RSnN4zethhH9f3qzkJnKckYsA2fggwizn3WP666O7TK1xJlPhMBiU01n8wBn4JyG2XCD7w1
qQW0hsiMwaaSRtd8OZubz20sGwEmazSNUeapCYZhWJJ/qKI2Wj93b6tks4BPQMfUEhqbHKCEgyZi
7aGchxhbmMs/nStysINAGNO+XayQYks9wreE15PVPgiWysde+4rOtXtuSgOoWgU9FLJfW+0nLA6K
EhkWvQgFKyPiyLEbB5BA/xNFYkjqwkVPZYTIjZpSxnApSkjmWkO6wwwWbWubyrlv3JcIQipiwWik
GDm+kTxQoA7fjmRSS/4k9OcTKszDk5A6bsfac/8eFsH3ALPvXAFFzkisEKhf5FzpBQAt8ciiXG22
FEOVL0kIGGl6phL2aLUjPDSq8lq5bDwgF5XDerNbpd1A3yyHZnkags+TSmlOieZaa0+1VnpMyoE4
/z1Qf06T0AFDcZI8Tp9G1OdbQdZ87KEnlZAvjwZDbSJQTI81DCLGRieDuUmZF/pduIBaFu8wa7Re
w6dLUILLzN+iTX+r1V6Rok7P67J/vVTq5KYNyzoaOHpDUCCVPzcXbNJHdCLq+PiD6mLWvzzO64rI
iAYspsbJO8aPQ0wetiW8rKbgMF9fSe/nk38jWDJjP91dE00uVV5FVDRG4b7n1PG1ZUR/PK+tcVFv
B+ZaxuiGglJ84Zndpc/zbXMnYbWf+UrnUKx7Cu92incEzkxvhFWrBdjUdHw36lyYYUBzK9w736/L
inbQkIvOsDPWtrytc8c8vjC06CUYJD7zYauIel1eLE5gOZoUzwC/wbeGd8QF0q//PRMuY8v4IAss
ZFScxNyp74VrKN/lN0jCipWwCKucNxWwYe5GRJnpi6sHIwJWZjAQzs16Df55YmwdWzlTT82jP5mc
lglBHHvXHZf0FuSZ0mDnahgvecl4KXx4Z+3iMbsNbQlivGp9yl5ZA07yEueWpCTBG6I6ya1hMBF9
Tz9wY2rLk6WVTI8RbTq+F66l6FGcud5t+RaPRUej5j7zYMJwulI2rXeoVf5Lq1kyyS8teh1pE06V
Tf9UIk5iVdr1DcK8p5+m96sFbXc5n4FKTgi6jVXrzCF/eQyK5eXMuwZYlfif1jbptg6u3t+VGPG+
FisrrnOT5uHtJjFyTevMFTHt3e43iwj1ZOPOODEsu7TjM6saBW7tJfM1UYxyFfj/RBEj6JcuXnu2
t2ICJj7JGbcCF4n/aOaqoeC5festxWj8/vYs8HQj7CkHHbk/7U9fVxQIUMtRfpeW7UfSYqjpWpOp
Ix6hPCYxyrbs53iHBikD+9apeZ0nshEn04KE2aCJTXEl909tjkHSltXimIP4gGZiC1F3xYBqxKUh
hxdxRDFZdh6g4b35pMXU/ArBSdKlOnwMHhgI2/SOwGTzg/dhlYcmRc/5nicpoZLcBbWZJqSEog0r
dBm/IcsVT/aHEAvpf+2dwkxrLwle361pcQ2adyQhPwez1tSdRgh6O9595308Y2AQzZ6lpTHt5+DK
fQZfv4M8zcBs41a7cScpN02KW0g0mjIT/WZv3/oEStlYSUA6MwpJ4o+WsClff977t86YqoW6F98b
8NqrJrFFDWXrCaSMe/rrZjr2Mj7DH4E7C7+IXvTiJ8QbICkG0cNsOIpqaAv/XTOoxeT3/SUV40wX
6OO4Xp1fe8w07wJva3dTvvSN8uy8aj1XynCFZUM1/tzjAjYGLAqqaqBj0abZCFhMXZUB2KgDkhBa
uljR6dlW1mu36V09ShozzvoBe2P+wSsCBVX0+ulTG8xvqsegybR28YeSf3L1GLKcb6uj8K1H0beL
OZ2MzNwcS2ZAFQdUC0A7CrazcschlM1xdRoWQPutnEWIcclYzLLUrdQW2dtV1zHr6C+g+9Myrh/X
12rPb1yPconHEC0iG9QLnTr2Rtp5XKK6s+76XB13/pju1GlA0VBsG1m3aR4CtDpsyU6ekYslq1CW
rzqvHp8BNbJifqxgeW/x1AphBkXerfirI6d9d6p+UCfXTIewAXl5otTlCrbgprCTbPHI4figbCSy
LVrYbViQjOKUgUWxsc/+QKVXD5rrK1JgHUfCoXHWKD/hx4jJODBUvRpOI4ZAnB4DYP2ggVTBth6n
dmr/BgRDGt5bUeoSXniNa84kf/t/nPUxWjZ2b9pxmsVHECnEPU8v3TlHzTPV+qBc3bZ2Cmd4vpAU
jw1TnBTzN3/QVz+Fy79X0CFaH1VJBLwpeL3S1moY5QI59HPburE/Fow13wZHO4ET4wSUDvzhG1xg
jSNnT39sSxvjAxOAb2QbZQ2vgsnWZww6J2Tdz1BkjUrRYJs6aikmdCFYIglnu8OaZUnL0fMXE3Ns
frqHtce/TFzCICyO9XmtUoZDxPO16Y1w1TRin9Zz4XtFIJxDU2a88PvUVQTWAtPOEOg0JoXx7+TW
RbhnBZ7I/KxentX8Np1vJBbhL/anI09jtuPBMwG7V7Tmtf3tAOalyWuSM/YNX2VKpNA8ny542prF
NiV9CSNVjokzvk+lHJejxgAoTueUWOKCv0ocf38VtEk2FkqQWFhGBVM0/M8O5A8ot+85ZrMTaAz6
ZafTgEHR1TJ3gKwldBHWTMGDVVIHY0Af+HMIgEw4A9g5uRpRLM8N6pir/6YnEIKT3tyCqI3TUf7Z
T6IcZ2XjTOL4j4WFqoIek+HX0A8nDJAr2PPUuCNsuhUkEp2IX+VsM1yD9HfFVWcqBHh4jw3Ub68a
5gGq/n8vpeOXPvILhnf6/wwfI/dC8Ww4AzKCIFuc24zyvs6k++LsNy5O9EaANWkE00aPfngCP6Wc
tsA4+xrmaZzQXtF4IyXUQ6P4+h6pJl4/cZ6c7wApJvVlF7YcPPrbgt9YaNKwJBlHng9mUDn7iwO/
oUX062y1TRjgXtTHD29MFPI6lWoFiZNWVIMsuAXB/S52voepf/L1EAuB980bvHMLBpxmcB3wlCKD
FhVpqhHlWbtJIrPHcVx1P1i3hVDEl/Jo1Vm+kvziJmH0LPsUcIK+txJmbkl3wEwAi2Hw0uL3hXSF
ZXAXJQN7uBkNwYuemDoPjaaR7CnSyKYrK9etCh4q0ryaHMWhIHWurtlJVhJ6HQqzicUHmJi4dOfj
MmbC5SWmWctk/qh7BLgYqxsa0LiNH0eKiie2Eznz0+g+g+OMyXrWA/2gGaPnGywVXWIeMX+abaZf
iNUWg/4pa8jgRfE054YgXg17zvEAAWA+r4O1ohrK7/CQdotp5fKtgnBJVhcTn1/PDER/Jr3KS11M
rLQtDhSBsoCwi6OO/mgsbe6dql8qjZptkqBoAtXw3GERDGiOkG7DBFJKu0wTDqNdWZSYNRyS5V8c
7rflpxjcv05S9Lx+HZs1PTpl/etiXSKFnLMNzTaUeuf+fdAx37ok535FSITwYgarIioHFQGwqq/b
ESvgc91c6WZYB5wK9Y7OT1vvCBjt93PtMrJqmtuAhWaaeA0YuwgpxZ5+RU+PWYN/R3JHGKrKs4gv
T3LSfFidHkJZMksfuTVPR4lha0u3tYTtCmsJXKCJNbQan7IU4C7MTASsFPHadrK6v4Aq556aLXXW
l9zmIRwuv7U9JO5g6FQg8SxN516sPntcyYJk011fRMwpj+8dhr9GF1P5wIjGoxxOoW1Pz0O5JNkr
tKOG2oicOUzfTr/xRe2KYHmHsqvUKsM21vW6YKi2/jD5a6K8OTHt8WtB7gtVs+jsvijRl2WGCL7P
o5xMDIDHLRS5sdP0c8MaxCxGlwL9q5EFRgTS83Wfbu4shbS96SL/fVP/7Rb36kn4MAewtBgXUJfy
DS903Xz+5XSUIhlqYqX6t7y93+pWDu1GKNSf6qtnFuBRsOctOCrXEoX3lCGIS70dfIuSwBX2PEQM
MJHakYiKVrqMTxNaLHMROfljH7t93r0xd6tUoDDRjVndAaKoy2OeN98MUmHn9uNHOjfLQH29nGrj
5d7bT6kjQ/Umzrm5gGd7dTr/3++1rwTaUmtBK9O3rQcVq2duu3wKKtXDhRDx26PD7a8pSydh8UH+
lgyi/Mjs3c54souGIWYxSNaCFuDEF6XthfP1v7073WHV1X9yR42/X3D8Cr1chpkdn//vWFzBepgU
RU2WYXeuphY/3YILw+t0EGpc+WKkqNJpZTbZ8GWgzLh3kR9FZ5MecTlgpCBEwF6WHFHuJlE3nx3L
3QqgxvC1AONcD41Npvw8UNPwNpACGWN7JsiAJXa414fh4NsiwfuSFXFLPSd1ljo6INoFCRrkXUSz
K6wCTFgoH3CXqMXmtjg9D86fKFDppWxZwiGqbrZoRfvUqxHNX4dyTxJFqPaxjc3qb/nEJzZMyJKq
NaNVwnfk9FUiDeHG9AFHw6EcbelxQCZWCBnnm9+uz9rywFZ1TtA63cjhMOgvA86azP60Wllkrhc0
qhe6IqFo/wBBSI73Li6yHimDW3u7g/MBg+dRd+0kOcRtmJ5eyuajnq33ooOwRQDCB6QHJ0EANcMt
MWULvV0kzhI1tZZV9XDqTTmEaqJ0WT/NIo+QOj+7Mo0GqeVdW0pb3GdLYN9jegJDl05BWFQEZxhQ
PPvquhLefmXyyBpgTs98s+DV923gEjyUNpz5gAunftM4PKSgenGTtKiWit1bOEhyyXZsD2+5Lcba
cvrv0E2fD8OtgZR9QcgXUeuE8ztDdN1QXNQLsoJlPF7nv3dTL9h5NuBPRUjW+5vjdBN4G1mme9pm
asg7/U3KDWvWNF20fy3FBiJ3cYtsf+hRui8ipPli3cU/wIz07yooEdHiv4p/f1thP7Exl/9SRwvZ
/tqVSbmFF6iRy11dqrf6X06Dmrxaxxv/mRUDz/572nfUgHqghqsrjSda4bgS47uFNUG2apMS8QDI
RuevgsG0tXj3r2ZAnUBJ6ZTLsI7g42JYDnGy6jKi871UrkgaCDJ1GfXPhYjdWvOYecG4Jipu3H8y
OxTJTZbrmiKKa4j3tCpyaN+8NdG56OdcKxjfeZaPG6/XnOtjtM5tpckMty3/RdA9uwCM9iP2h3py
F4Jzu36sCeRwF6Q+m6pZ4r88b/cM2/NkiZLDpbeSjUcC7QnMXz1Gu6pESf9itl7O69pNPJ3L1LfO
G7aNsViWZFDFd60UY+WlviHPAW3ctWEViXoscpZKuHzr01zhs5K3amA15xdPN2jSiP1ANpXhrMjj
/hD6+L+qu6wgBShfq/FBd3/Z4gGfbKjhsVfkSjs6+javMER4/t3xDtWs13PSLOPKREVhIOgdq0c5
gkI1mlatvqsH7p7svDD9f8gU3V2znrpU4z7nl9zs/PWF7Vdn/GIfIy3T2rL0wTGNAJNpDmwCx4PY
0NRzhk0baCtJ3nFovz9QyJtyMQFF02hBGJJqOuSeX1mscNI9KITi9iqio+A+brKZhHlDjES3C9dK
0c4Wy4WWVcUmzFFfVBDbRxh1uE/aPLpAbc/cLazNSKtoggb35nBDb780XbL+M1kjcRKKT8pk4Vg5
RYKA6QAUB7PX7j3yrTSUIc3PpybRmbcaXsHV2AyRolkGdz3wesQAr2Zcg2QJyL9hD6Mquevem5B9
Qp/2xiFEJtYVW3jNYaLB3qb2meC8zqgEcfs9GSNAngnB4pEesDNv6Q8en5hDRyiwkgHrN9BVWo19
A+Jxsh4gmSTizMdYQneRyQ2vEiXUBhgNOO0ygg/QzPaijxjlfE4iiRym/Jx3ZeXMfdbLwN3hEGre
EMNsiXhqxyY36yX53zEYfukxsSD4no+TskgIdkQTOxefpkXoi+JsTO7V9Gll0RZJwHDAzCX0QAHd
tf93hFcgomKZ0f4/5T9DQQXtmkePeHHon1zMtOBagheCMjTox30GWMB04SlgodkqENKmqaOn+Xjq
1SQcBAHpXvByOy3Ae/Uzhwm9/4r9iU+wgQlRZEMSvrEjCTyCBWkKqLDLwsPAqjGQy8GITbfMTvkJ
FQ7l5rvZQE6K4jSlrLG2OCaZSQdJdx92xt07t65yr4d0C/Rr++p9hlOCxvXfG2fmSPqFSQ6n/kwb
H9e3IPOW9nGsdhhQ+IlI/WrCUWDcGVHRbP5GyTAw7b4GZh2HWAj+IVM94ulYefn0J7htTtxUwQt7
q2q9ymvKNx0vcYhb53/fxDVwEKaWsII0V/2JobgLKO4eYv/lx2mS9CdbA8KhrKnSoklomSX8e2H8
nH2mi9Gzbblsxdsa3YZRADuqoFrNPWFOxv93TVbhzS9a+3lu1dAZHgvoUDPlx7XRocXoXHd4YArX
kCbrXUKAkBr42+NYGsByzuLtRccxjhZ81wpefWJ42Ya6JGGoZ4mb1fpMNksO/TQgPx+Hg+PbJWBv
nvAX3YxnvYoeUxMK0urGmkrri5hgXNpWcB5CSsioTYB01iR/ljK7lcEMx4tFmOMvZ/2eCAYighzh
JZwY1JQ/IUXXWik8BYRJbM9TR5O0GeDYyT8akZgijFuWH/x8AS502/AL40mhHgGlXk1dICJ6ygVc
tnMNIJvESxntoEiNjcgfJVeku+KCX6Fbk/3I7NQRszYRPDaT9jHDK7PnaRLchPIjJVw2m50q9lXD
0QVi7MHXVSHDZjU1xvl/8nAHijx3jSAXj8clkjO7ThvOAQ/FcmN0P3xLRQ5/0bzehexjZ0VhyD3h
npALaOO1M7+oOfc7qwoDnEmYITVInM2EdKHI5G8srkZwGxRCHJ3LCdQ66zL5qGeB0t47qjH/3Q7+
pCKfvoIoS1rcGN8OlqZu2pRpPF+0Qvg1qTNS9XyJUCHomc6AVoLy5ahgkRvL7mmIVLSiDrSgpgSB
jQvJ10sBJQYkp14bk5IdN9pd/KV8262L7phqclzK6kBxtTNDq6q4LwLobKZQtdUTVUPnN+PvBnm6
zj6lwANGqd9nh7RWG9WbO4LIsYWmj0x1Mt+7YfSU+qZ84m+TqzLp9sAB3sKorhfmZjwtWBCPLVLp
7B5YtWqVHeLSu3Ufq46xtYYN34N96UOR4jECQUSZZKDqHpax7dw2Gm4yFgLz8pyc6DiN/VCQJuBj
RXKZhDodJcu6cr1IDOyKdmJGJgDMcGRe8tdN3m5Px2+jX2eaDYoeF3pKOB14SIYiWlckxPiPjqEZ
hLllHsTU7yFqMbnbTB/CvkjyqiO/P4C3MBdE/QfklIpny6QjkACeBzpIH8SXaPVyL68WnpmRejk3
gSlgf+3Fv9QGYV4v9HkEADsVRW+BUwXM5j4OkErBA2hHw1uAT2yim3MHZ2IKOOLaBoCDscEH8PdD
GBf+ZKDt7rKCmKw1f5Ffev9v1NdPcPzKkoIg8taiRC/8E4Syugu56hofxKCoDK3ezHQqMrqIovsK
on1DVrmwL1tSRdQZGaIU6C83vQEoRgID1XJcOR7Hua2noE+NB0HEBijnKuof0Q4sC7ixslZn/T6e
eWtOJ/feHGiac+DzCXm8Qfa+oDmTaEuoxmThlvAk1ZtrmG+/PyKgbHgPArSPOHLkepMOITrPcukp
EGpVj4lStezHazCpGFzPZ1Z30+uO3tX/efefoXfcqJ0O112fCEnupe/pMC7zm0JtoltvJjWoiYmz
kKEcWjIWdeFJj8yO9F7X189kx8n0YVBRUdXLKeX5hNIyuFM2xTqVDnc4JLrfmmKEunnQQ26YhLJW
i1ZMS7WBfPKmP82OwrLMFa8t/ZTMxW9t9FNYX4RbgeIXmqofqk+HzQpQJ7D9r7u8vxuqkV/ExGxj
3A44aTw7lv2RcAYLM+o8VqwGLoEcsgzHFnBWHhSaiNcAvnsrd+3/30DhXIyFYvCrbCy25v2/Pyti
8vrdFYEJYgVhleeD0zzpa4MjvmEuxG4/dTduOuIB6AyfxZdCEzktg3Ts1Qwu4JV7wxuFJIomX/2Q
IQ5NpEUkGz2RI48IhLXKfQ3padOMeWm2ZAqE2VtphOf4TlkwpWU18scX58aHV1ZDKwjsukxOUMZo
Z/5BKgMkKkaXPufAfZiEqxz1vTjDq6TDdIzoBYhEJFKCyqzZPotbE/S+G12KCtXx+YqARIcafiMA
wzktkClBkNrACoU/eMe2guE0fVSEV03Un2gIQ7lLf40he58WdShKEnxevorMh/Lu/TlH5XBDQK6d
Lae5fsOi98PfapWLXNCp1bIjYfzMZsXBU8ZP0F/A5mruCoMG/8r8yJjBAHCMR/p3ejDEBey4Z9wr
dx9vRikDJmOdfeKFYRfvj3tsdgDq8qyvsVTCrnHe8OSbedH1GFgQtn1n4DJFPPWzp7qDo91FBEpU
5sD8E7XWb5TCM2nzgQO6L61iiqN7M12dlfxEHhHy5KK1xAoh7E/gI70I6+My+5wInmUsafU3u8ph
uVvRO5buoPJmGKBzGhx2GEMMEjRuavLGIj9CuM/e9z5lJcIdcqZSr1H7QXLJ1IJNaobfN2PllMqq
9BPkFxVDVfxVp2JrR7aYIu8UjIQM8HpLX0eSdz569u1KOUO2f1b41hk3b7Wy8Gk4mcZ76TCj20ip
XdyEyRomFTrASwyB9cS20/BFxzyZfARG0r10VJmFLtS2JzZco2kBEWsYU772rqoAA8C541ISseES
4KBRF7sJ/i53+iPsh4N8Fxjbcu2kHervbbRuNUNLJb6aGgFENvrleMry8MF/8VKPTgIgm51/eJnV
JKErsL65GlVI5Oflh0rm3oddgl5296SkTm0r9bKpq6hP66KMMdmYEIip9xGUr0tns37zD3MpAQqw
QG/9Zx65IG0TZrMJNZ5dNyAAV/7EXRwDJM+4e66BacxT+0bfg4c+uIpsgyucdLlLyzOml4NGDS8d
xPGABvAWCmlTIGTc4RHqi+tuH4EEXTE3uXU1a94BsmiYbrcvyiF9dkeH66XWkrvbg+k6R6KewPZe
yS+1AvxvjSAejKRvg8owAYOuUZPalnJlTG1T6oPKcas78QipoQkzJ7VZDIitOv88bBuUsSv/AwoT
mkrZ2EejLvOIS9P5yAtcCsioIgvQykXpd/cICLtWBV+S0TGVQEQqMe+Zaoz9NlBnluWtTePVJ/7g
ZUBNdEYGQ5WlXJqT0u600U8fCKojunUZjlzrRdCot4Nn8P2B66evfQvuw8pHk+8+ALLIyUNtZITH
TQwPYPeYt483knEo4GXWIzzFE7VG1XPqbUC6SDnjSeqoeFhvsFFLUGkZh1G82urywp+OPj8z+s+D
DV0pC4MjsKLRZ3jd2kQ5yTaXApUM0FHQ1MLKXssqxpsEgtXWb1f3W/U9VP3xhuMhtXB+JxaT19+6
iIx5d+Spe8AiPA03YJX9Z7vZ6+YXaKVMef394qLDRQQ2nomr4U2VzqVNRIqLQUDgr1Pm82cSQMuG
6JPOiaTMHY9JIUJvZIJnroPwzIZ5/8E2NNAMT1F7pdjR2jUlSUnp9HrpkMEAUpZ6gNFIgX5kqMAG
AbZfjwAOPEk6va8KLrp1dbv+3km7DptY+8tDGJ1I7iaup9BVc+0LBZKJNJICQdADdMyBVANjAGzM
3kcY1zichKP3/S4Y8kNNe2+aRq8Axe/GjYD1ecArCtM50PdhJ/OeDPbpedkHO0h5tv2xXCO04mbD
bMcg2rMOOjJIyjM5FT3b5vbTp4u+mfkHAiWvRUNrZGZZtoW527qfrFh5n/QDy3EvvkyhEfwOLE/y
pxMCyADCVJooVoXAHUtinaG2X4Y0cIIx7iyiqgwdu/BbjIkDCL/uqfy6gISQvH9x74c2OBHz6JuC
CzZ7WD6zRQrmPCZtzKAZzpKr5idaDJQKvzEqLj+1k+iXeCMl/+nrLFVCsBgK9d5FW779d2JKA6f3
nS8/uWpdW3fBhQM0+vly00cude0v8juoJ7UUd9tnDO12hiPKvhQlHLtuLy1HGfFRaelIeH5iWR2x
rXe+L+WIUJPYuSFj4dSfKm4L7dfqF9JfLCiHhWpZY6IxEvUtzI3iExDsWh4PFKgPaqYXDCflnUsu
jyLax82Z0rRZ2PiMq7jMVuhRafeVtBDG8UIK7xk9R6hEQ93ydQJZFelyP09mCE25mj8XxW1Oepd/
6CGKumy8kEao1mOttwweL1/iZ1i2WrxiZzHhHUokq3QkyguR09ITOi6ZoYljyKi0cxFs24WrCrp0
ZsTIoJ8xhYoj/lByfp0Ev0t/tDy1QCFUcRzdYmstEWHBMfqKdmwth8Az3xb565fhrx/ETJyOAH6Q
m/r9K3UJxloSgOv/MXeMrKq4+tEz8JX+bxJI4RHbRqkyaHHl6HVTxoUMUnsN74It9h5FdxDBEN17
pDR96g62yFbcPCmCmajyLvqq3jWzkNRPzDoOGxh3yBQrUdQypJStuR3yFSkiAyMTV5i0q7E3/sSM
oKkmZ/5usFR2QKqGoEsZbf8CrU2mm/zhUyZ0mmLyNz1ekaZZPl4fsDVuSYpiAE/oTYezVwwgLXq0
5H0tI+vtoKZz1CdLHhRQDvqCMOnlDMz53oHPtWrT1k4KblnE4fg4uCbTPTbA007JPI65X3PXyxpU
AHT2Hbvp84uODzH62VDQJeNLf8JediICFDGu9f3kbYNYnDLS7kwiOBEXgQzFLFkMAwaLWIat+pxj
Z6+VqKOEwWGqNZg7OnRjNhnf+gflBG6dPst7Hu8BvdYlis+wMyr1bbxTp8ODLXppagY5W8jRQ6Kn
5iBFzbRtTzA9blJBjANNdx/kxz4x9BNIJ1rK8QeIbesTLRN7bwy/G9c8rBA01XMOdJAKhR1UW6So
YtQTXkwMDlg9TzjthFhSlOD6yL8ljeVYVr4MA7zViVSI9B0gZ7rxzk9LThZlSSSzHyyp4XbxJbqI
Hcl4eEKK22DhFEBPPvga/iDjwHNuBx2KbypZyGzshVNGyaelkTT3RnTq7o+FuBaajZGD2XwW9+7X
wQK0sS3R7GVpqWk8ul2mQZ3X5K6HXSD5wqQWN57r2oowQth6oicGAu3FqFtBXz0TC0zsTKOdNY4c
Q54G87q1BC0UDgvU0e/TeudeTtcIHn6sSMjq4KmAIFbdRWoIrfTerO2Pp3M8VmTgZSFQ50XvfZPL
AkuaUMbRcPj/P05lbxCAYQ91ipCatCxnHrBcA79n/+igaexn5wlXcGVj1PRfpjuP+MbVald8k6PV
ieQxfOghLdALWjVK6PcJmdRw3Ln5F2y0hlKn/keuA9T7IQe2fryIMcZm1/KKMJAwJb6cfkoqY/Ov
WArNHmTlIgL6GBliyhAD7SdyRTRP7bkSBCfI/Z1kfL6y8/CXkgvmVJ1NOHS0J3mSTeMDMMQFzn2B
X8EaGEaSkzriUWiQlEx1crVtmMIjmVmAjdGTMsXDRckLToQJFWC3W9vKbPk4VaU/nj0gNVSVkRqv
HOF3gOZ89tTZLWWa2lihKVprSp/STht6fzrpeiTqSb2vaXHtfRCrT8wPX0tdHteP1Yz4eXU2BU07
oX0y80cM3NxzC5wibXo3fOPd/60DPnPux1Xpnw+blh+7kqETlRGDOf9hDlpOV9gpVa6xbE6+1ZOZ
ChfO4/xPe+kx+hWK3j+8gGvORfRukoh+4qfgLIqznEHO1aMFdYtVGEiwUEpLs4YbJyu360icGm3l
Y9WxPy6o86rLkIdJe/sLDSp9rKmERd158+VHp+coYESss2PFLFSBfTP/XrmLxfSYlxAzLJrrRcKH
YDSd49SweFBxSJv2nEEdm3deEuq9mVy3P8toUl2NgUHP006mRd4ppV1yUlhXXIKVh9lIBr9lnwYG
vHMy+pzlMUDau71fnmv+MUPTBttkQpnvZtO+r36sNPixM8529n89GQcVOsarFSuBhJwdaboIMyDA
F8Dt8VwnvChjJgPt3la7MnMYtiOeKQXy+MI4FMKnxS1Y6q7LkbysYkI1Vb9RTOABBdTGoKNqQ3s4
GYY/ZtoXNzGj6h70Ej5ApO5Mw6R9PwWWRHJJmWtCCpToM+Lq8DYaYQAlSSgmzY406WxEpGtjdtT2
8fGMPZuLF409/d0CEf39tcY1tZ2/GSwZOgki3oPE0OchLtmr5gSt+GewYsZBjRISxrXU7RrMUT5V
2UDhObzS9Amg23Z4d9cwusoF4OrRD28VKyPFCy+p+TPPufAoc6N/chozRLgQi4lDqJvojsC4C9xr
xkGLV+6S7B4iTHalcGwGqxW85tgKgxvXW4icj9eS3M9VpOIBp6ji3rm5T938+2zH+0rbPhYu8zti
DtoJibLYXH1vfkPkrRFSFvj5ay6OCeQi3nyANqNSf7llV4xWwz2k1QiRocSPC58zdqX3jP6FqK7T
RYtk8sKboaYSpUJ1CY3HDaMRiMEdJRB0oBIQ6aNsLPbOx4hooPyWffPeNt+THaNLHO52CLjszxEJ
FJVIpeIp/uat01TS8+O3F+PLpdZQ555ZQSpyvcNDL1BFtFLyWW/xX9Mu011SZjcHHYaPK4JyIbOa
yAHGHNavc4MkLlaM7MDaauhGaz/huIJT/J/wu9EaZi/ZLh4mL9HBG2r6CK6B94g7LpEnUEuLXLfw
GCSa1je7M1b8ZFGZBZpi3ynaJx0ItyvS8VwefxYKzBqiFIPr6jvtBeaHAs6Z+8EUM04Z3IW8HlI/
Cv8T1jNx0QsKam3w44BxuQczWZtairEn0R//zDiiORiUAsI0GxmHn1a3/eSZcYJH+HwsKMereZKF
YKRVidae3vbfkQCMfyyOgCeuUogAzixmmmj9dVNu1brGBp8/u2UHlvQNF5Q572JaU/oVHHeHGRn9
D5iwO7av4PtXYEHujZJ2mc/EHFo/s7FxW8FF9LMQZhqFnqIMlHGL4yxiXeeKOTIWhtnm+cZwdYcu
PifeiYKdM05p95YchKxUjUNftg1T7bZm6frJHafXEfW2153WDmqDfLX8T85cVOlwvo0jNOWdpt8j
rNxtE7O/HSIr892Ebjx3b7DSACcBmzvzWvw8diRMbuE5CYqiDk9FVhJrmpBwsXAAnEi1kKi3eN5a
cMKGif0LxxqP4vauAM4KNa1oJ7SyqiGsHcb2bj+g3BYtfnoU1j3+Exu+vb2If3Eww3SOXc6NUjT4
Q7xGMugi9sDRpLH/rYx5WvgX2IkzA/pyi2kw+bVQEfEVtz2foa/BOU88dkPmAHhnLralkvoDuBny
oHDHrQ6W5AM6zYngBOn60sSIEc68KactEvG4nXK7luGYhd/766sNBzm+r5zefsmEwcXg2EHMbTWW
X2NOG+eeqZVFBZkuPCgtrx0//tcHpmMQQNU5XW5i26dmKUdEVA1itsnZtb8U7f4hd7A94aZCCp8k
4nhFKPHCURHNCZ7IaApV0FY3yU9XHGoywybjzG98Oz78oqJx8B0PLpsUjYdQxkeNYHO9jyVdQJzk
+vwAR8/IoP2m2U3ONojXP5KBXioF+HxIbrmKDZonLo9CY4uq6Y1ArSfwh3eIlFUw62AkLsog0XFu
WoZWbFHM5BQVVHsS5JowqkcEBUpNraaDYCI0znaSYcSKonTFMQHUSIhrm/mWjKlHfIHC7ty0jMZw
/6Vr5VqRo+UoE1WPD9acQb+mFuM40NblkJ0w69nDlWtAiIP0fSuXDGxBkBA+qmhN4zkGgdRTcBZe
EgCdYzZVPGmNfclsCQfWTeXF60I7w6FlUY+nz2RTwzG4r1yr8Ymuez1sjLxLeU7j9xBHx4UBOdfS
mh7hJHOhI4gwdWgffAlJlYIVhM6uPByboDXBps8YdBNkydL25RkH55KHEhRTo3zbowngATp27oC6
QaDW5Bqvrn4Q/ctW8iu8VDLIO/LCJ0bJTiZWHFIBtDZaywMXsPIANGjzEdYOOb1yS605Y941kC6j
KReunymYd+VanGe8b+QH309TEdVde5vwn9xllzf+vbtPfEdIRKE/bEJxJRrlwrP72cfH2c8H0fRn
m4HMvX+EiAMHu3KIWEJnblXvEK8/7EsvPc7rxhWNfIVAKLtAhOEntEm8vwh7xGvLfHAtvRZfGhSj
r3vSFJO3AEIcjQG/Y8d+uzL+D1YmDrYAdgYf7W4vaMr4dOQRL2hMi90LS5MCcOogpvvtPwYAxTDR
zIsYwzgswfEaAO3CUUfyBpuVmGn2+bW5/P2m5SC7UOGsoVbvePk9lmI1xw9CQA+EhysOBuvSfPiV
cxXtAXNSLCVfK7J0EzRPMMTzb6tsbRNzJ71JaQ9zTedQhn0Hfdq81WFtYetAnt8UbpVGG6WmJeBU
L/RHkFe0Q4HupwYSLwBNlBSb66b/9ER53tolbKMAwAQ8mjjHxtXa38FacDMJS04R/9/Yv/zzHbFl
wmhDeTRGI7V7MxLQycR+U/qnoL87c7o9CGzbmqjMcOS+5otIT90lTSaopXR/N9UyN+T9X7TLmIvi
YDfxJUt6rZzck0slOJ713gNnXA7eKfDeypX9SoOu4U40U02MtZlEhD6RJudQ9BeqJKIYpRVGu1+4
szy3U9T19wSSsFRjJczt8ygE053NHqD0DpzE9SZDfN79IUXPXsXAUP7nVHDKvEmUjoX4Q/LCHZ3e
jtQ4jXvfEBiipZQ2+aem3kYv70nkrlJV2x1U4JTrmwWmR1mRz5rbjjNNnX1jEeFCVFfKsVeTBlQX
A2p0jgNvwHbh84K71Z2hB40jZbbwWXLJyPuczB/Uo28HKQ8i4Coal4foPHGNic+yibQlTTPLq83N
jIacAZltb1/eW6Dpn1wjkELoV5oqzWWiTyQz+hRtkyGY8UGCaiMIOghjlQ8KiYTcjJKjkt2VnOSN
GM2Vtm5SedHYfNBi6BTBYFz7jExUj+T/zsO3P00iwA7N2jbz4os/xHg7aO9YtleFx+yW+09XG7+w
uCHuT1tFvGeZpMoDizKak3Ml0ogJxMhAMUdJbjI8eDR0oY8Q8R8Wc24kZ0s6LskH26xlmG1BmX4W
LsolNdsIF0Xx6oy0pCwi8X5bo9+DSbf4bwOuKCmLXcnlcPgKsiaNz5yS/v0ZqhYf2QgtWrFeMmnc
zo3gEm1AGRCPffdtEJqv/ipr95rNulbDnH0QxEnhtwf1iJYfKzxT9128hwl4sTbI7AeWIC9BhPL9
Oi0fr2u8vC0CYiC7BNo1KcMqXXtKNZMtyFxFiYv/5MACJh2OoKm5PzY1f10c2f2dvftTReRAZJlm
Wz9igNaEJVA99DNX92YiA1s0lll9cGrl6MymYNFiMUJwZQkYr4VBfzEjwuqfzq0Tx21klKMWdgzl
ur07FeDLiz8V4OnxYl40vfRTeEZHAdUi6AfjVxgyG/OYXd9LMOdKRZJtOM+kzjom9YCd3vTbFI0v
a/4sgN8Ke46o7HxcrwMqukXlEtbQF36flo7qhLnKTbqC5LDVkMMDE9DHZ7DpCWqV8EqW8pg48rQA
SG29erJ7rpjsDaXLg/MoNz+D8YrCybtw4ut0XyrvxgR/ZzNpHDK1dVKqjBVCunV+LlBiKra5CfXp
RRl9crRrl/ilSXRW4KhezcuyMX9DoBzYtG+E9IO7CpqJnvPciqbuYwatVA1ASeSkdpinHFaZoOr1
oBFd+05xeCL5GRJ3qWTFqz4CCEK2PbIz8a8tS3zmMNEzeetpEFyrfLCD7Q+OHV9bSeiYBURU3GUX
x/1FCr29ayYUqyeu32kF8jnQp+0XUfRf6yQeukPhkL7eU8CX1sWbznUVPsOmIiQv8l6xKh4W8vvC
N9Laa2W4dduUNdMivMco/CkGU6qMWCVaupveC05GU7jIfC2jx3iNVydJ9hCHrDmQ1L1obOuL7YAv
f2r1mRmggktEfRxRwXvUnoqczVpSMl/6ALQOQTLVuicwBTwV+9sHHAbZeXolz8fKvX0P97cvLw1m
gCFFewFFV14j5zWft1fRKb2digpej1k7+6VUSyVstdbwYmQRZNRGHk5C8D0IkBC6i1jg4GM93Dz1
8A/sNuBC9ltEz9hq+rRDfk1SUY6wIYPWe+hgYoSRLCRySF4YKO5CVCIU1rLt27TFLvyhSQqP3jc5
pAIf/zLfzBDrKb+fjQWDVVV7VbGEmKM8AWYw/GXkS/VxExyGTz/QdKmJ3YhHxWLa6CYgnYpRcjbJ
VV2N13cDBVQQHi71yUtwxPQ48dirZyZt9qM8VvT8hw7Ty4W1u3b8D/WnSSRZllXeLimBkkQledTn
AmcMwwseS/KgEWPWDA/nkmYb+7sZtupf6fqmSekvMaHalSM2l6bvfMVDhHtElBJhsgkdnGQW5bU3
3GEM9KCkqV3dYRXeWyZaAzUC83QKHp6pvZokJbrhOz+BHCXAKd0NakOdxeS1oWMealjnk3bie07u
85YdM277MNqa+luyxIdsIkT/SHj1hPWjGLWZgetbwkAMVmQJ9ocSgAzHEwC6Gg3IUO6LfLkbWyD9
TZGEIZNo8QZC9ekkOaZiXxpILyytmQPggFE5+a7T5NV3oqByLO7lcVxWA88Bligia3OUw1+GzIj9
QLjqMjj9NfHxWnQVBm3XF1mU0f4IPnGKtIsMdDo+j7xvnV9EE67lMBsBX3ayxfBsml6dXF2ICU4D
yveU7THIlVTzra+UpU3SZ804v8Ip5U07PJnmD3jGuuhcC5eLweGq2hXQ2e8zwzYqetJhx4p62Wr5
uIq74cqXgvWkk77tj9dwKd7b1tSB9bRzlS8hGezNWKbGzmNRiP5upBESiBHqyvBMBmE2GOKnUql+
f+zMcniL4BjiiNt4T4KDjIAtni2cQsaRX02Pg16IafEy331tqweY7xipJLZ+UP5dz0us6IlyWkkQ
dH4O9Ulrapcq+TQsulVlprqVxjJVzIGZvHTiEzHk5BgCAlswPMy9tVCEsDUFZXOyB1RwvHS/6g1j
kctaha/ia8W1MO9SinY5mG5OV6dWwJGEty0NT/lrfnkUGShZxIsuyTZJMelxYV5q7aQi2rMEvXzv
oHY+x0yj0knG0TzRK1ywW/jVWE+9xR9UDJCe2gmub3MDEbYG4pBu10fq23PIb/kpUt4wRxSdnH2N
hyzrfwbswSZ7Vr6oTk5mEjvQQBqvLoidy/jOBd5Fn3Hc0UNPoi88krOyJi/Elz/IQHEvEMVGMO+E
48I0TfOazlw8FhWqedw4pKLrKon6/axrkPc+1+1so91TwIGxeYacN16I++wtu5S+BHDZT7W472KJ
lYajxAxYzkZjXGqXbLKGzz9Ucyn8C+8wRz3T9BmUPEvuyJeZyeksucxYhzwaso6+UDFqNk4lpHgO
p7cMHr+aRJEH7EX4CZgVKT5WwtEvV8QZei8WVJBXcdpslym/pcTktfDoet+igvOFeNLFXxX9Rvsj
KGsLT8PK0T1WCqmVzi30y78FdVYQoKXDQJBgQo8pWiB5NHgD630TXSXPjo8uHxRmVW6F+pVbV1pZ
2Jcc+bhiBpL9gaf4KlaE64gDBrWRaD9GHud21Bk8OlEJToJJ7zN6pt1XtSGv4TNjPodmj57YoLl/
qmlHraH381MDEi8+8JuWrwF/P+kSG9Dof7hcz0P+Bas3Wx0im4gSwYwhcyqQ7d7mPwTyTS/6q7BH
Gg4gmlrZXrUIpFn4yLH+AP29TpTKrfhUBd4IzKmf/ZincHKfO1su8SuY23yrOmvNliMsQE9XkPRZ
6essZArlZUhflp01l6s+C1TqHH9VwCmIEvVaOIVrdPuGVaKKv8RjwkoqfyCy8V0cBD/y8DtwMADu
fLE+w9T25LT40uqfkMqfcQqosG0qN/iA3QnY9TOaoUzuiz9HJraGKBR9PjTOQtaZoikos+bFOkLF
AmZaE/DRwFGpOUPeZLM1qDIkrYSCc49YccUAXYBdZCI7ktZgMQzq3dBNTzGIDLCpziUfOy7jxYXB
3H6Bu8NiJv471Tb59IxxOt87nqzFctpcxGS2zLxBmi7WhCzgWsvcoKbbGNyoJIas59OzhCRAsgGX
YSTFRIzuU3/qCzHYbBDJwh3nwRVs1p0uwXm0ofMtTtTXrDllVjjxqP5QpfkPC0BqAO6m1fqBMbf9
4jWbAxcMTZUuTbTpgLqPf7n/rN8HM1yMZaKVWGFVkIAClq9/M3Zcwv6yd1uPgTj1FS9A9wMwHrxb
P7DvnIwNp0+Sy6K87aHP/v8DjVFtwTnK6LVt9/fOTw5Uvj0MO4VDwzIqbhau3QS9B0uQ9NZWo2a9
8y8WSkFGvDDTnR33Vkc/QB4cKpSeVid/xlSKPscAB2ACot3J9oDWtEQPXNI9f+nbK4g/rcxmGIm2
76xAepUZ1MygbTFonJRH4DYdykUWNSSIQ5IJsQBOrWMbETrsT73v7twXovPhcxLaUyaJGzReYO4W
6D8zSaj+dWmM2lJHNckiSCp7aRL8HDl+0z4vyoJsMghqbdrlZFUkMAolQ7whe4+FgpHL0anMLj9H
iNBq9YdX5JS2JPOUPIgnPEVxhUiNFhF6ojE28AoRs1P0t1FucgEhuDa7p6lq1jaVvE+DykLs/iC+
EhD/h5O3Zp5afcQBLxHAyU1VHSWZ67om3wDV+I3yyC17Ec8jcH2cg0OiXHM1Z71bGnWT2TRXPxYx
saAfpssfsVX7KGGpRzvPXTtKSYyrCK3JBPFCixYfwbfHTx4mFbWdS3/OBKOKiCYr/0aN50Zy7QNG
zb+iSlBmCaBooJqSmjFlKdiTJII5RnvfWCL+CKDxyjBEOyUp5Ix3KWCm5gh6sujATfMNHdkcJy26
qHcq27CJM8BqWbJXiAdy9+2st4T3FPt5DIzXxoXmO0hehVocpO0SdOyXEPmZD/z3tuZHkyEdyHvu
4N7BHkyanog4dEztCAgJKMhVWGDTz2vXHLYBnqoZN67fVy0jBAv1+XAJzcXd/8ZNvh+cbAk6Uf0s
EJtgRWHuk/BX4PzMCTcI2wPUg4a7e25ZEsQKTGGyBl2smMjrAIqfJiv5OzUqC0OlzW4FhYDkioLr
rPypZiHhmLIaUzROGp/aUu1op6TrKXdp/01/a6IYitI44wrEtl/OFxXDgzlASWx9MYPQA4YVj+z9
T9MuOt55PSx6ODuGBz3xWXCrlt6afL3vPAr/y0WL2wilDPXsZymoKnqeo8PvtvDH74X2tTuEdTUO
jlVCHBi8MulanuKxRgYiCyWw/K/27FYZSnL8lXEhVZrVv2qGQhBbhs4VGIet3h6OvZqgSlMBPfxn
MSKrV3hbfviht5KYpBO7q4ZOeUen0qBMDsO1SVsfY/1RxVqGiHjVqH4T0tGRc3UR5C2cuqV8rEZ2
jaE/VsnAS3xkZ0tLupSlLpJlf4AE4XSDvLg4jJR1dQxyuO/O6nZW82jMnBjdA5Px9/GxSsiW82m1
OOLKLqFLlBaGbGlpXU4mIbhqis0YW8oT0zEyo8rRXrM7t47h80tN3M4HPFe0/8ZY5YR2VYcKPwLy
rjX32RDymJPXi17M8Q0OgTvTo0JnGlh4qeTT0Zc4BD4Ypk/+7XZFGv5Oiuo4LEg1kR5ZZKnbtU8D
fGAAyGX5bCYnCBAn6yXKXG8ltYHnaJ65kzUuwFCKfvFZHctH8tUMvDUiUgLhNPymCYAKiaI1Je3A
cmKNsWSvm5T67LdJ3KgysJOg1gZaHRtwO2X/4wW1UlKXgInmtE8Wzmdij8ZkKF8HNNjyC9cTUYKb
qiS51zv3HQE82ER8QEXVZnheLuIIEmKZrwYhZ51kZkkyy9HbkTQeBktTB9Hd+1c8r5n3E3BawsnY
cpKgEiURN4QKn7LBO56ZLUUQ0CFTubf9gxKiLev5sH9kLZsH5FaS+3cde5g2mc+6wTg2WDOTM61J
2Et1X54EWTEsXAdIOamrrOjv1MaNm6Pjgl64v1bg5P/+uL+XT3baAxjxBwrFJFCWi0rZFue0tsLD
tQVW0ryLsUQHQUv4yqyGTHr3pH2Gmhl3U5XKfvGEAhdj16r4qdJZKbzTJgqQa44e9HhOSWtTa16g
aNj6tZnGwP3HONQ2qRVk2jOIPCsHd+6RJ9oHp9NxF1n5b+iysqKCfwIUs1eieZQBtjHQvj0rSSZW
JMEETp7fWavvGglg+0WyPlQj70COxRkSs97/y3VpAfWATfPa/B+2JWTEzoTVU3JZ33+RSVmfi4XJ
BXM3l8ljDowftuy4uGRKQKURSNSMpD+ZP1Bo4Hg6Hkphe7FUYJVhD01vOi41KePAnoECzCBK2t3Z
KMjA5FlJzuaVITM6tpnngC3fD+pdLZV1CMfSKbdNCQfRhmjkSP77LsvAhpwttBqCLkQbBh0tIft6
ghZTebS3zQJ2Jpdw+PWoRC+KZBaCGjj2V6+JOhDBO11g6kVSDnlEv1k5ygu+kV2ASutS5+xSP1j3
+bdbdPpv2HXk7pnPDm1yiEVXUrEggH3nO5NouXgdnLA7d2Dpwk1CcGqPaY9m6g3EbONTA0ET8X6P
nqiw51CWW2FY6dOsJ4IFDd/LUGVTy64hXbvAyeOX6/CCdFt2F5hhDnj5cXVvUqNhPO89YAuZ0h0a
8S9+HSAInlhkXcNXea2ixkxA1awmWeENOxGLhxYizrdZCiKjUT4vTzq/tntEv63FdJcjruqmX8SE
kAkroZ1gdW3K3Xnu8ivb/l5mv1xWy0l/zplQupiaHpfEI3U/B2ZeO51NUgtdjbqdJPGrt7l31Mpc
Z6ztUekgoBNSskbMcW2/eQA1ZGWHIDl+cxw9Y3NEAEUpwxSslaOM95CmdS5Bi+JB/8RBedDcncCN
l98njHopF6lnkIk5GvSF+Ts91Cfz7+owNnp+ALMTxrf1fhZPZaUzsCyagRsnsdynUpi0DtoZdFEX
KyjC1WGBoD99wt4UBtPWy7sDlRXJC4YqHvUZHpi8luEFW3kpizRFG3HUZ5mwT7QBUiln3GRtkIJc
rTU+RVp8sSJd7RhD+LJbzOiyzalICR0kNIVZNF2DsGVLr7E9PynWwP4AOs4ZJmqP0t+HgDD17tFy
S+HEByM3wZ1VFYVMbwc6nk+VnPjSp9guWTXnPX4PtQahqtlIYiEjVz+uJ0x/zAibtUdBp/I4H1M0
DbdzN16vCUIWo3C4M6tYAKA9P2jpdZuIbQvYaabRu0BGoOk86ZcJWn2T72j8hBJJl/S74XyqoFTA
n+EKYwMpWUTDVetSjtiDp+bjxbjIzIusivTTdDvMCyrBGubu+NvpEXPxoNLcDILUcP5rQfqz3Nky
oVwTjDBAZOMqYyj6k4EPaCyRXb90nqoJnzU2Dfiil9ZVRr06Nu+I5lf3TtmGsxjbfw9Li/altOZF
523EWMB4Y9vybRfxS8+TiuImxZcinjbcjL87JhQu2/BSooGZOVEHw7kroEfEzJlRyiQ2su/03iNM
DLHZuBejipRC1JM0QTgMOTYuru28sYE7HpDuY0Y6p3xdEGRA4TOd6CGUXFIHJk306qgmhEO72z27
0mDzt3W9ulYyZl0Mjv96j88iKY3xghlJUQn79aIX/LbZG77URwkHZe0G702RaMV7FknIn1XOBnx7
zpHa+Vj4lbjkSJID/+0uhv6yvB9PIeyaBu+qROmRD0yKOTbYwMIo7zBJLedIZ5vPN5L9vTghYffF
vIAXMdqcTPOb/wKSuQDTqTrOqxGGUfg7L9DKNIUHJcpmS/O/iexiWEyMg6NaYb7u382UmXBu/1X6
zN4zd3Ljc3Hw9ab46GqwCJWyQ6oB5xfaQjD/0Qgpa6T2KdCOtk0ZFzZQgizXsOC3gLeHE6e198Q/
WpYKg56pCbS2/ix2m/y3mRTOgPRAMCteLxlu+Viycgx/y7msRUZ8XDuVl8njoFvWzU5pp94YG39E
I/3vbfVtdn4u/oJFJSCfYuzzZPXDVi2MldacL0sqmoYDTCclebxfl1CtJBkt9+ijxKQsYIICzyqZ
ZUVH8FC829cEqM6yYNJWhIUWO+zLUb7tRz3mmNlknxAIjjXlHK2uuAvARC4dSACyeViNX/SGm0x1
av0SF5rUYaIkjJDtRdn6OsED7r513h1eHt4MUe8idBkBixqf/26UF6ORNehUuYGOmd77eCloAT5L
jyXGxEInG4808P10EhXYV4GH2PqF29CqYuDJe86WPaJN7Xwzh95EjrOfGnNAsjrKzPXlenluib41
1Wr4x9nUGVgmxChLMbbLUiwFEcG7wTPeZM80m37D1UMhgyG3ue7xSDao6780nmE+gYJLTuZCm8ru
l3s7dMb5d7HttId0ZcMcD4pJs1wVZdvJLkz9xtY8tcukuGl7r9X1V95G/u98oesRjdQ/sajubJqk
Z7zkYrZPZXDvS3F93LgtnptOIeX1qguH/6s3yXBBD4yDMFBKjYn0WSB/iP0apZWW/5Z68cHnSwLS
rCIRQ0rA/grePZNANL3eCJX7Z40yHgAf16HeTKqyg2d4aPFhUBWMI4TjOlPNJ3xgkof0zDAiB4Ev
8BM9gVE+OIh8MwCvtAJCJwidpzP4hQ1pPufhVUAIEYn1lfbqS2u15r7t+rz4QzIIumhRGf8d1uus
aW+5OMHdvdKDiGn+x4U7TVSIv+Hu3Q1IFh/GjJCVG/euArj37+V5ylNZrgdQ4sZw5kLA087rVaC0
U4w4J7trnsB60sZq3HAh0HyXzurUM+xsChaPboCpfgX9UvbxzK+vufHDf25lDvaszsrr1Vv81a3r
PA0wVhNwupVCOtEfjJZX1TZc9p8xynS14kLsRluPIwUccr9Bt5e+e+96+4Cz4js8Bs5q6fNZvL1Z
ZpsoO/16KHN4uf/KoEuJqSBXYGFif/FjeIPVmqt27rYCj/yNhja4GtYsPnR6kbdUGrnEH/Q45IFP
l4VYGs5GIJn1wzC5nehWkhQazCUAQ2VuQWg5JVjjdZ7vl419fJZ+0xedYzF2M9wvRlEuj8BYfGrJ
B3fVPlqdkI+UkmVrqZ4UCbpLA0HazUolyYhCdtwSB0q1fiKO/XCw0BNXo77lY7qgBSxk74rM//OP
Fz5OwVLBfP3E8+gtLlW0+Ogo/T5SKcWAwnUB9MBdMG6gAIxWBDNQuSo14qElB0tdh/6AQMAtjNJ3
1nE+Au1UQeelGf6d63lGWf5cWsCC3m2D4PrsVxTtXAEMkFZ3o2+fUdKY9Bw66vR0pB4Hhfk7yNMA
cGK9uSENezayC6K6SJZdj/1qHAFBw9TH5IAXn4CEAbIoK4kZOH63pZntM7KEW+Uvfg9C/d41ynzv
Ma0wbzgyniIPc3tKti1+GS21VlQYChVnZ2GghsxcPCa8ycgD+YMtne4CMRPDG/kZKizvjbj0QTcB
BgoIcG0JVf4D9oddeuWn20IJaBqlGmXi81zg6ys27nyuUYTGhU0ONMOHfDmG0Xs1bGuZ4ywfGfH7
JC94ixgZw7pFTKdS3J7lSKxTXc2QugveGWWgPjtiAOXqA7MptAXMY9QRAPaRYQE37IK7oIbaSvZm
unIaewPrCTJJhH/oHfUvVijnhJL8xXMwjJg29Vjch+PSNpQ6jEyCbtv4LKI6OSeVm/J3kiGXIKfc
76EZ+dQZA1Uq9nSMh6uRYywDwJl9TISZfj2bXwWt68OA5xUvnEm87t9nByHVlyMTqUmEDLHioeBU
isi5FBP3ibT8xLOL8ml6dg86YWmEM8/95yhiWhYjU3+SQulHLhKFqcB1/zqlvZg44TapDUmW1cNK
VOFUDeoFgF8fCYsAOVVLbYmwHw9ouRUhFJkipFZ1h27n3J05Ts3vGZHmeZjsMhYbcGiOvm9Brumk
XGDnGg864YAenpO+/5OiZ4bxbhDuIqfdWOnVqWop5feO3PO+r7CvtSawCXdcmJbGHRw5ShrFdk5I
Kqf2gnVGgZMwnEoNLzg8zan9Y7MceAd+FXccYWJQiEpY4sb1ww48tFv+gbjgOlZ4qhR0gAA6bUKY
hdIDCuUQd7KIIsBIUzAJlPAjv56QYYXooPfCTD/YluKbjw4f3FdZ8Ibx8hD5EjMohZotsA7YZnB5
Ou67OmeOuBBFlevcZeYNuvUHIhe10iTvYPgzt9Eyt88q45jC38rKQRzvZuAaX6n8J6wVzg/uX2mo
1KBKcBLfncLSK9dj9CyCG7BUIQHKdbHfUxQA2WeI2HJcp9Us7v9uHB4Y4AsPrajP6ZQwXpZxegWZ
kgu1rShYItKZfveldum7Cj9PbY8dyGIoctO/3rstJ4DaCpI282TdsSw01mukN65XrfHcNTAr9lG0
zS12g7NO+AlTM/pge3LRNppPFeKLKBb1hveqkYYG68qLTRVcAhrfQd2sCCtVXJywNNJHFC4V7Rv1
jDcrxOYImyUI992D+B+O7OKAZB3aOi1wig3toicZ3VSEjzrzLGo0RrHaEHmrb52l8H/HrS+w/r+E
6UCLvAPFeSXBJ/ZDeXv2gUiwIui42/oVs7Wmqd4B20rRihbS8htBMUutMfyAUauDLsaoGbEhGVU4
zNouNlcQXzRns3Uw3rNjMuFNsA4jVxZ/bVfNcE2E0Crrx1wGilWRzdGEE2nzcdOR92bgwb/DZoUR
g9JSZ1KQp3Hn5DQvFxH5+Lopv/f8rBvE6Ic8l+NQEQVmqwmZr2OHnM46M1TcT49sWr1702mb6TBS
aMrvbGt2/2BKkDVicDEc+LVR9andr98MLiwiOERtsZ2BQtRfeGWhMJ8zY9qAfAfS17WAPMf3bcsn
1W9RWOT0wV3wiPDHEAH9ABTOkAMUd86PhoEqDGGU5rUmeK4zcRL2/aNCCMc56YF71PUtB1cpaNAZ
FQKLjfoAPz3QZnCDMwu71WsbGJWQKHAqccXaJNM0qV0qgsieWMtu8yqx7YsL9RsHYG7qewaoojFB
/851vWnqovrIEdd9LsdcCDeGysye0sBhf9Uu3YT66BVpOdBHVldaANFczYTmXqIEQOGbts6ZKmax
3/inReamcqZ4k+8iYII3YxPgYEHp0H7NZjRU7LooKs8nPwCk+549qi0CkK9AYhtPetWOyhJloygk
I2aPvC8Z6IozWyl0zNz3O0wkSL1rNL1YDud2POBKWEOTX/L0t4NeUFD1McHQ6pW2pOnTMoR9K/Q/
qNt8jpQ8l/XhdZ/W8EnBDU2FxWOceg334lViFyQkWJcTfCWM+Wb8zya8nMCk2OQwBw54BVnsjkv7
udyz7ulE9KR+an6wzwAJbaqfn4xBIplQsSYnCeas9XOqU8UUgLJl6iN2BJEA75jtoCj5eUlZS5fR
1H6+P2LZkf7IkvoZ12zot9wjLt45M4otEenOxsW2/VlVex19idImyu2goszFwgMHo2PkNLLdDLx1
chJE7sLXgDE75YFFgOx3hINXWsaVBONyk9bb9sM0FgqswU/dmIdFLav0mgOgA458K1J2sZYHB+/Y
4QMD5bEz2Oo6nKnLPnvOi8lku/zzziIAxTIZuC8cJF2FcvEKXK53n9hxJAHStTxObg7fsgXeVbqp
RvQF2sUiJ/XyxxIt8zxvyX+/3+T2BrcB8MIjNGAi47woDxF73wUj4tYjMGRT9su/5l24RMjZkaB6
NymZroVxr+G+R/cs+209Igc5AnocM5f/DWpuuN/5WOLP9tA+uBlVJleDwfHbV3ZpAjji4Yg/6Zus
gmVaD69OuOUAI0GfyuKPzDV4vIAbMXTixahnoz8t/0wRQaOjC3SF0yDyWcYoKRuS8A3XI6wKmJGY
RFiynt6guAEZwq2bHWBhUY7VgMZMv/JpxlkADQfd/JtL6a8tzcuUDqU8TsAxE/XhxyzakMUP1Llu
NF8YbjTIXwXa+RlbUSFzhUpgL4SbzIZUzQYHoHq6iDCy5H3CQ3bzEQKASuxVk/4QcP29mA/QUm7L
pybpaIYv0CDBFsIn0NUVC8AyaTh5lXJbgfYDjvFBwk1S0ZLWTnNq/PJslgrfloGjVysW0z4Nmu8q
DN2jrW2lS6HeZ9cAzElDPLmh3TI1zu5FBYKoI8w93WxniERlcGjHhTq0MQlUIyRXXTRxY67rhCwh
i4gAJZl7x+WNrDSCo0nOGZVQ7W5P/v5f9VC8S6xaUrvqEvyUYvOBNyF9MNamVV+2ibJ4ALLUuLj/
khOx4ZphwEGS63r4a6SlK2GUdYOXguoMuf7eDGiyBg5LMQM2VGJS9vd9CRCR+KF4eu6+3k+pidwU
jlIrl79C0jgfXfdj6AcPHjeppmVrshsmcmmyNjMlS022ACv8nAMgH5FTve9F055I8dJmDhTzEY2Q
IwxPAzApPMj2YHWBUT21yw0ksmiiBU456TULRtLY0onqbPl6Coin8xL555JnQKyd2SGomLGsClFo
2uQxSdE/IroCffy3fJcsJiK15nSoqSruHBJ5qXxk5VBAdOBszEtmgQIXmCd7Qx09BZm4slU/4KHz
N+7h/BjWjQBpKpW49/SYeTr4Y2Bqm99+tDeF77wf0WGKUAd3MbjjtHrgsGIc58Zlf6Rh4+lX0d1x
YvDUUXbIw4cx2pmaIcrHOjZ0Pvw8YStLmFNDNP3IGwNti02cYAmTyJHA9DZcV4kC8JFYPZJTBo0b
qi6Jqy1QNX0AR8wjSdl7tMA2vsp6E81ikOssqFYVdTidqqMLPrnoTHjLSl8MZR/THvNI13Ku5Dqg
a0wiF5WNiqAGSgJxfVN+KFssPN6xOwZwQrKTXHXMMyl5Wu2+DZYVZ/Q4/VgissvgMJj6yYmSIw/G
cFKXn+sw5Fg4BZmGOZVG6Drri2UW0zJHzukKGPh4Ueg4imq4uPj2FDi8Me0C/ODl9Qwfjr0fZd6Z
ghd51HUu3FL5YJj3MOJTPrIXv8f9dPFSjzUh3gR2yeY/7A974W/XIoqGvydFcLswv1LUh/0nfDaT
mKnCJP7VzfnsCIY8L/koPbNbpGobNKPZcd7bmwCqOzktnaf+JM/26qOmHmKYT6QVWcOLB5OIowN5
F9nZiochlMnHTa5HY7TkUr9TE7qxcc3c/fREveORAkpikQzKtZG66UOmYTi1zZUFUoVSl9lWWoem
0IiSqBTmjmmsbk2ocmqBJaunTRyDi9hfEwq5fkQgoN+Nnr9EHMiGLsMlP5VgHDZWtNuOTkyz5swi
PhEhwrsBBobrPullZgwbJ5e2xd5cSzLHH5jvUC+AgQd5VAqUE8DQRLvxJ9G7ZtOH180vDkqb7maF
h1P/aAqKLMpoUBiLj5+LG/sLyfIloBLW9H3jlBfgQrIvWEhbdUXObT/AYq8JBd+Djc3QdXged5fU
jJdHJU0+lTGzWs94V+l4/FgmQE5B93UEjSbIoV2np2mBqwdeFT53KA/8nUXzBeiz8pT62k32/fCb
9HXcNJfBNM6wuK6j64wMp3OpDXdqPBg2+18EvXN4m7GcY34oWGupDTaMYTLUP0kupAnNrkvWwMcc
GVHDeMSa0MMSMNeIMj9t4/3xSDAOSFzjhxkRkWgdGB2ZW3TIg8MLDug2WgDaDiMyi0N4ULIVt5XV
cyamISOK5UiQpl0Zw51rmX9r0h8s4RvSSQl11KGvLoTnhEz21LVT3wSBY0eEX4s7xAsvaaK1ChxP
MtmklTje8gTmx7DHzd0lDkGbqZXkpN3W+kI63V10HaRVNGBfgn3NLqEgktTo1p0Mp32QaSoyuGmM
Z1xwfpk9VXrDi3mG7W9IylyhzpPuY0g0Lpk2+b9PV+ZwcRBpjNN+OR5R4+hwk16IV8jhnQFag43F
XkV+Y3xroNj8YylpWq+28gO6aXNHpuhk1yX3pgUGWlsneOSo878DC7QPt+fpFMNoyIEDN6FFMcwc
22eY2w7psiuMhAEB1s8DbvQK+/Pe3VI8a4kx8jD/LJ0NvVfArIHD/FzzWagbsIeONodrEW5Vnc0W
WC4WxVlm8RooyCHXHoI/MdHKxkAeIMXkg2G+tt02FFM0O4/TvaQEKBlw05KERH1rIEG/WuxrqAII
1W1AuAdJ/ivDUyhqaAMD3BOKi/Abh/6uxZhjSK2zNTjenfbycdz++CWPkoJF+KPAHG4wB/CAtqvi
sTDwZ7XURPlYrD2KsrODrt3gvZM04X165RpNYAwWCczcfl0KM7Dh/KvgluRmocljBZ8V1TUjtjdq
4miFohw37XRLrJLhN+vUYdplzF7c+IWp5ICtnwAl3yd+wikHqeOceR0kbU7PuCtJj774Li0+FAku
TNO6fQGwc5f6w1A68K4XN/w8oZHF5ptE/a7lvwWOqvhgWZD3Dl8YmISYzYY1L015/kia7r4oXqpv
Bh6Hq036d1kPSZR9Bt60HA5mET1WoMm5DURHxMZ1pEj/7kiFRqyA1PjHyAbjEfmIr5N39jr/Z5vz
RGm6RqPR0n1LoRpIpIk1u7V03eTaKPHz0slX7EUpQIGY3RbgGZ6Erm2IqJ8Szg/18oPAkR8Aiu92
Yra/luIgpwjKF1DxVKfPmwt18Qn9KnQC4GKC27loh8BgSv/QvFmn90J3k8U/pNXLis1pruYwCAPK
J7+eHwk8VV3FS+mZF6XNuMNtCQDeTmj7NHuIoL5eVM7iVSmwizi4PrJ9Rhvf3AJSc8CuGyRxy9aE
BhMqFXIA27oZhmnNZVxchAVGCpnKtymNrv2z7mM+1n3l2DPzoYM1vj488L7VtGNlRAgF7SRjFIdk
drboi0aVFecr9HsiLLR6iYQs9boZDr7lG8UkfSiVAFPZUl1tViBeeLZK/NSHA1Thdwtlv65YhrDh
xmHQsYyV5ryk0GqfV1RQwnIoE0PkhyKVBjkKJj70qb33mGQ/gMOSfNvZ7Q8me067y+GjRAJBLJWJ
+KNHOFNP9SY+NE/l8LSKbQjxZ+aMGxMEbPxtbun+MGNfwqVM5RlfQOER/UEVpyIOjBBrg3j7wJt9
NmuibZ3v9TFlYOY5/XLnk3D8q4lf3LyhrC0J5b0rE9bP8Gg90CjpUAKqeJfVdPyTH4iMBLm4+pVQ
3BXMDN0Z4vLlgaZ+ux5kt6L+QWMSXvezT0hT/yc320t/efm8M+HCwumrB5IAFst4Oh05p7QuzuEX
R60AQHno6a94WYcQL44MoaiTnYNy3gh1udxh2FcAVUfZBJD1i2ZH+Mjg15zKQSuzcJPFI0rUXXAX
eJ/UvEKwiteg/x9/DUu6AmCTnDf2dSZ+bST29/lemU/kjfDnuidBTRtwIy43WqX2oATUX2yL3jmd
41FUJAK535DQI99SIwlAIUbFMjX4IRe9M97T5TVN4Gq/WLQfsXAUMhGAbLQiVGQqahHRi+FmeOTs
4cZbOerF9gDMHyEthNf8o7MsK1RRRIQj0pv5FGrCyYUHtHyVcv1gsM4yIpsuEyS624bb9pBdaEDt
jELqy/OVNNdq3sEU1AtWDqnxn/OfqzpouOFYmU4jx7humvM5Rb5zO+tdSguRt3B8GWyG4PFK3ejp
kTRxKimU35pZ0ooB7wXGelpbRWoJyX7S85VbE8kMTcVJj6B55myDvqY/KqxzvVQBCigSNCArO/6M
NsFHQ++7K403M27YkowQdJwpIc30c3EeJNzDZAqIdRWEiamc1G2/jg/TkpLCDvM4QSN6SayhoYfV
m1PjmFECxXZkme6vy0J2gSt982EzmB2oSksLbrne47/GIZPo6TzLP/LAg+AvErh9chEp7JIk9Pap
OswwI+PGU0jrd4u+ouBuGP1e+/iLyn5L4yC0IhRJTSjdLY/Y5FwKc1qIww1/yQoeQB60tDcPPY1G
ItfxD7goqGdDB7itUiu/PUHzVIZzAPBTprlJmrfdUdD7kvaDlSb55rrT4VZAlHjdYW/VSPKdq3VG
MWTTZBZcqEz7nI1wS1p3o59rGPvrAsZ7rziY3EeNGfTHqU8lAN6HMVvYIzV2SIgnp4iyp5gYHn76
QP0lDn/rnFzvMNmHCKL1t/JGRQViAvOcxVt4EWn09oXM74nbdiaTNybpGQCudI9wA8ZSwCHkzWbV
mu40ey+7eRfL7xz6tvolKHiXCvLQ4ooKHNC2LV5kjFSwZVt5xn+UxuG4kZGAcepSd06AGfmbC6JZ
2Br+RCcSrHWNR437FrqaIa2VibDyjF6Is2KC4gYMQonSPPQ7u9wEqLJhMmE0qBcggC1/3fdqu52A
llhOEnYaFP05wKy7zjBgqIgx6QjIciQQsvNlZVOJWG1ike/ryf3TwrcKW5Hz48Tqsu/sCQXqLwgZ
1xR52hG6swBaT+VVTOOqXIZQgukc7GIeDIfhFkw3HgGSB3N6jqmHYHJGhDrqgEEiFK4aT3wKetQ8
OA2kuAtB4jfVPU2h15Nd5NCWGkwFFiLwNSZlxItd6EGw0g4pNs/yzjh1kossywDJOsmOOsib4ZtF
e230R2EALSNlXULTghDnyqzFtLpe4kGWKFLn6nCU8wLmN+jPLa+Z0Tv3OKkwpOew+6EI7KRA1cFW
l2kWs5a/jzCXbv9zVAXxUmEtSvjF9CINM4dItRG6OzEdyBYOX6JZBtKXbIDaItIlNMSfU9gw5yM/
iQjW/6k+3WvEFjVF25ltUygJUgctDxLjYjftDuMPoEMkkLCQklKsXI6tQ4G7O2mqW5agkfG24cA9
5917T3QelHhmsHkJSFnVFQlHfe3fKd59z9Fibg0x7YkWTWDajytujCGyvJYDERn+QyTxXoICfBCf
EEvtWO6wmhgggA/hl9MnbOrzJY+5PURZVl4rApJT9YMwtHjsccP6wagycGTobi+1R/O5wzQ6z8CR
VM1s0CCY3v99MyiEExdIqE0D33KPSUsyETDdtr7aPeAuPpjATE+/4ByCtwdXtQ59xCZWG5zKTk/F
X/u/m2HUUUGR46wCcr/92ToHJLmyOLdr3XwSAMSN8WsxTElOjyZZlX67luhwQm6RI92eC2KeSzMT
XHpph39xilGeDLNxm0FvbDlaqPKT7HfSzKTqyLxU6ZQKvnI9lO7uu/McghuDykqfxtD7nPlLeVcb
ZqoM2UEzJJIkVcnrkzrPeybFL5VYmLImJkGCFYBRRpaPsKzFuh8DPUOAL63imrqD8dV5YLiLfn5b
NCgxo4nOYZd4UYe1X/hRp22Og9igDB9yu77ScUiivlQAfyqZWBMTWymu+AK+yJbJoj9smymzrDkD
25yVYPf7C6Tc43yCoDN7dH0s+G8jbztF1MpkkweLMgjVvHL1O8H/vWFbxsaKfqmtlxgGI+Cto/EI
K73Z9VBEU3i6Cyzpvue9YMQcNO8Y0UrzpyOBJgSclchmBX88ZtL1TuWURIee2Ac3v83fBNpU3jmp
Vt1SjCGBK0W7y6WsbkSKOQfJIxtP33cClSBzovINjKhMH8KN8INXeP4GTUunrcdJOWHz6SgFZtyD
it1eRXMxmCVSgGDjgy3cPbmOxFfC1MFdb74AfolDv76+d8zhnlcxWvWC+/LzA7PGodpEnxExpkD6
fJkQynNKiJFjvXDZ7EM9vZa0mHvr27JKwZ7xR96HmEj1Hft8vW0reRYDnEfsz1xQl1oErYrRJTHN
YkeFhuzCUL8nG8BYWGPx+W6nr/2hw/oxegPBSt3ZjQv6GfAVV5HD3OWi1d5svLid2+X98jpfE9dw
1gMlMBWvLLRi811ijZ/YZ+LlNsTZaEoWcD85a+z8/w8rE0IjIilvpMatViXfOJ/Jo1pIQDLKznAU
XOI6LdkPt/E40ZV+nWmHGAwYGQ9THWSmot36DXVPY6B40Y+5opoDNdnUhcguHuxLx3mKMe7Qjhb2
vOw5w0dEWWhtxVVBgcxF0RYqc1RX98/EVCJHZDL22uV3rJ04j7pFARUQMcpnuHjKHlJl7zDCi673
KAtZ3QvMeKMilgAPh/+pjr/gx3dqoMgLkpcVO/0fSP1gOWz4sLksiLdHgQCRyLvO9w1i6TYNvKvg
a5J+U22VJNZQuPWxE++A4Mks8Kfi49xjtASJloeFL+TPEjFB8Xci/MZlD6MCJt7svwuVcILSAjRE
B1AoP+XfFU65tIVP0LC6KaUwuaKTIPY4yIqmi4rbIXOkQmWRl8I7qstWSGquTxK+HxlC0YFfYQLm
yAUAggpG5S9x22J5pXe/cx5Mh8ACyTyIQNVJerseWXJNRyEYPKFsmqj8wz/mtLhE6m51AzqvrF3Q
wMbbxezOZLUBYJ5fz7PmxRgP55/9YOl+qntsOrw0h1oTrl+S7vgE8eHbPzHi3A1GW1nFhCt9XU3f
OvLbr1eejyo0Ocaj3XuwRgOOeC6ICziFA3+mNcHWY96qmYbmyeyGe1B1izBZbh+c4SPLLh+ck9kF
zznGbskdJanuYilFpmiqriT4O4WFYOXW3/LxtefQZmtT7uqJLHJfYQJZriMDqrMwKWSx9Y5PckAy
0Dqr+f/kcn38u+5phqN6UiuvpvpryPtt9uW7YVUreXjxfBdwD4Sa/dfXbtHpLvYXRL6fhJZhXRDg
jtw4V+aTPYV0iHNK3TLBCWCta0YZvWXX6nHGmgMJFO1+6ON0/H4nv6bNEk+e416AFSkKWye73yCw
Fcx3NnBQCzdNDFh8lNwW6zpVSw935jrcZPdp7psDyuEj8swPbPIMnk46+OQXAl75Px/z53YkPq2o
ecEjzXoft5cWATWnGa48MpmSUFzvVO3Sdn2JnbXZdN6RSfSZqH+oWFDgSzszV6qdH2K/2bIiGREN
QebT2kHlDAOVFMCm7FlKdrSbMNbGM6eMhciQAALQ41ERH0XynuSuxY1UTdTDbePlbQwdF2+vC0U4
Da6QQXXyF0WTOFL2Zzv5gnTBY5TMH6JwW/SkkMHVMSuABk9E8Xp5V2lGX1BK333Eg8PinxibRz93
JMrSOUL+5t1QWV8os1DP6KLij/t4gKjO0Xj+aleCgn+dshEttg+QC37hNzTlsVYUkVoYPq5tAvwH
dGHpFsyq55CofQaK8JNADLa/5ZqvJY5xjxn7TWo8eibUgPnVnTBxNOMYx6pTnPq6rBDi2wUO99ls
S8wJR8JluLZyKv+5m73Sxjkf+e4Oza3+7O/lc9hgGsrCfOf1Uh4KfeoiumEGoWnBXpFZT6e4WuJi
DnV5mcuu7GK8xB7Jt/WmFfkwhWzjeTmoEmAAy1JPd9E7gm7c15jYcKZLTjI2xDVKC/ftkx9/CxMS
RcuAw5gedxuSOCGnCyygu5DkqaR2szrO4UAlluC2vfO0NgEGqOrCfoFc2RN6weg5l3iD8CT1NnCx
enWUPtca0A8h+DvQiq3AyNzXVNTa9yXwomjVyIcD5fmvJDdVBmRkYWSBphhZ0W/Fag8mdf3NOztt
HE/Mc1psiHb2EmGPEFU/JHnocetNH/SHWoJF4sJKgdpkQBQtsXJVTc0G92mlTc1QWy2po8tbSZZp
uEUng3ZA2bMYnDtZsqnJd/uzBel8+ag280pYkEIqpeo5LAg1BNp5gSj/KHxH/pzkEBWte6UH3bLT
oCIGlc7H242EsriE+pfPai0ZaKAJKii/B9fyZwJDSaDbCXJZ3g8jpCNOAjXumgD7ag89Y9uX7sy6
+iKw2SlKteLF5eFUjD+Xphby5hmrAQUHRBqTCPJ28HQgYZC5QgdN925t7UMWhmo3d5nerC0VUXj9
YBmLGvX7x2i9lZshI2KnXAhHxRQXyxUp+wRnAZB1fOwgAu0/pAe73vjJ9awuExLp/WJvmqTQqQmS
NNXaQD31VBAUvZS9rtWSyvFVB9pDq4nw7iwhO2ZhBD++GFbxxf8Vvn0wbykU9P4Wusr7HNRIJW5h
cpbw9LswzaizshyhCSje9CZzEh/zTfzIfyel6Pk9oJdtHS6DHqCkiL+PwSHG/TkgXxuUTfwYxIGt
wuBN5apRFAdGth3tXyFO+RA4JmhY3g9tEvy3BddTcIpn9EKx+SY4tiPK3JbcXaAtE92kVZDLF3Pt
nDCcqgcYQGS/u49icBBn+lWZCdqqRyFvKRodAahoaJcdqsf4QJdUTU7u3T5WRvipSaZ/hQrujBg7
7PoK4eKeuJIQ72FDZ77XKCmEOeQjy44W1LHamv+zJWnysxbfWt0gV5/7in3RbRlbo6dswLZuS4+1
yaI0wMBv4VqjtxrrZ2meRHivdnfKq7cjm/C38kBFTi6aso3qb8kil3uMEnMaF+t90x3cV8E/p15i
+e2osJWf9Vd+HRajAZmzl0PgEoYCZQq2XenAMSFwJL9LmPS8jU2wwS7Mcj9R+j04OFTZr6MQ/CtP
l+Rphf1Romif2WqbKmyeNFZOihtIwPb5eY6jtXPpPFxvHV1kxk3fDNhnu/gR3GyvWwvEgfjLxwdI
HYydk7k71ZGUZbRHasijlG55XEm3Uu3Z4OPVrqrzrE2I16UF5Jpr2EhQRD98TPAVOp1cegbbZwCn
wz3445A5Iy+8xftgaSXS5otjRDM3WPeYMznu3AlK4xPvDrMtSUNS+UIm3Tm6OaMPSWswm72CWscI
AnL+/27y+6Mq3v8Gpa9J4nhlzAuqILsGTGFOrCt0eUd+8PcEV3wZAz/+04OD3vSKYBqF76Hk+xBS
HZFO/oAD2mNQVVdKBirSUFFXtzIt5ZDkwzpAl0aJ0O1WBo4cdsk6Iag3e/5vWaitJ5MIpdyQWomx
zzD657I+wXxsnfkDaQtk+xuuxKGUuA+v2KtYbuIh3FPEJPBO/+BIOFbkAFkTmy7pHbPUo/PpfitM
/Tqgq3Zwm6tlf4sOk+QjwDt+lZPpH+H/gm9XfiVUpZLd6N/XjrW0pEQI0XwsboXnHR/n0C1HZeSb
1nfifdlvdHtNpIcw4wTSUw1MzQn8X+n631LOxaZpPIunOcPKWo6a7ounY4HvuPzjtf8mi7iruqyF
CpdIqw7tnvQPhLo9+vdPkCJsjIuH6y9+X4PiaPQdG5tpFowcCcjUQ3azlvwtjvjxXsVbMhS+Smu+
ThBgQpbxamUuieG6cVvXIL7vse+SEwyY1djNy+J7JHi75YCkvf/szOIIwIpmeR5kufZd90fK2KDe
Egn5FsQ/+Cwa3GvvTlRCa5nMO1otTAj9l9CzfrLGL9Tg7LD7APQD1gvy6/5uMmm5zOYCGejso7KV
KXBUDcTPn98hrmYjyvt4PKzJnfIw3/qPQaw/DUk3/5ch8Sx0QmlsX0ixsS9YJJkp5I8erPEBnigu
wX8JYqk2lyHGylaQ0etrCVCBaTcTq9htYZwY6lQCG2IpnUvtIAzCji8rc1DyG0heTSkN03wsNO+g
/Vg49OBdjt29ie29cbaIDX1gXyiSM302StsZpVfinJGg1F1wwolf2fIrlsc/aaA5gZBvqBUeyoR9
zovfFZUg7kSndm0Nm1NQJ+AioRx0mKzmmy7awgbIEwCnofsDF7YIO8FWTXBJryhAxR/+MHBwUbgv
yZjQT6VAA051saGyGoyJHmOPLvyxf6HE9gxAzBcxuTkNH+mG53csoOIt4XcJFqILsaRN/kONJpMl
kE+Ozk1w6ZPfSL6o+y/IYBgX6dDbU/6ukbFrt43ZtKBACzrOkcl1TGjsy/31DegG0O9iFsJsC6Io
elOfYPxgAksKS02GSe+fw9hAMIyIsCxGqQIjqgIBfORFLNH/SMwW0Fh+a+XHta4BskddUqbN0wmi
HgDtGuq7qK4NycsF8tdY18V1RpuV3o0gPxM3lmpP+7cGXK4kFq489qmDszqqumXpR4PydLcYDtBa
k9Ua47HOJgTKjdExfKIrbNtGn9EbCM60zoEeIGsxO3zG38ngtfOO3+sX12wWrKCaTS08sr8dwwVg
TzgBmFA+zvmWjkyz60o6bfQ5DEMRPVOcVRYsjq6udnxXhUHb+Jrj8sMusZNBCtmyU9m1ZwubaKfg
YPwEmBUASYbuSArB7UsclVY0QQPsZnReectlf/CzTMrr5XcbdDkSatiJ67/rOX63TteJchndwAIh
0rh4YdpkZaqi3QqGGNqk2Zfb2LVg8wZAnli75F8dPm2rbPLu3pPm95PG3VCozJqMWUg1W3issrSn
CbMuHrLNkhVzIUN9T1xCTLWafHGx0snlCIINzDyunvzruSa3J4hWJ++B409Kz0OYbDmIvYmWzMNZ
9RASxyMnxjBMbPQlOuwCTaXOYHhGy7J6BhsiGMYDzRyChrIB/UTjEUuWUkAHMd0lw/oCvI+mwScH
aIpJfN+Hc+GsgJVv/wCgbrj7Bfx3q2QZdpfrgi3pub/F0JqUIcjekZplQDlPUQpM5sbGyn22JDOs
j/vY5bddJc9CXMA5pHD7/gClggISZFIgOScgEwyUm+xGH9i6Pp/0lECBsv+7VCYrlQSxO9aEInk+
FHlWqJqk22+52jp5R0M6cjskdd+FYZKEyytk96sRDh0uzNKIqX/ZIfVwGrPCf2NtI/02GRDjYFHq
vWb8HLTNiOqSraDy9d8QBGJHFoXAvaR/WWB1fyugH2Is7BlT4/n9SuY4Zl1YZyMOLrpYBCKYCEUs
iG5wGdXhCV+3JyUxxzI+w5V9ehYWlntd7H0B3PLaDntgeqOD+6ppOF6Wn4fWCRNH665we9+S7ogg
7AQWYiVkTH+dj0o/PdJqABz/w+2cmQIt6MAjPDYXeJcqIeuqsxAbRA5q1DHv069/EGsYv11kL7op
YP3790xVCYy5Y4iXWieWexw19teYwoO1kZctF1UvXGOWFcZJhKu88hYI6htJy1rlDye1jK8ZFYJE
2MDzAGHtyXgDxAz4aETcEvlu04PvwQ3Sti7TYgLD6UoIwlIEMjtiZn4QgJvqBNB99dIQIvaIHcPc
iA+xBmS1kmU+5K9WXDQmU3WajdwZis6KlkRda7UUJ7WS+sduaKe/k1fu9QzGTwmtuK3XA4Njb7NX
3m8jJ7ZTaigOG/allQNDRR8WnYE6Qapudvw616OQsNyeyfXlef68+Ecfg3KdI14JLWA6f4t+Rbgc
QwOohPPhrAzR/bSFWjNa1DHJ8HQXBhnU8oHjmL0FZg4TqWF+tW/QDWRoljdZNa5K3JJ6AQwkHCY8
k75ecc1MOP4Sj6CNPl3kAJ/0+HwhvtcW2fkNs8MNjFpXmguMW/4QBrPb7aLPtFrRJKWtEjQhqggB
HctrMtEkKF2wYYaB+BGwh5UOXe5fcuKo6TV5j8bEmOYrRBq9S4ma41wJTCZ8CvPLOSjcTswNCG8H
hfE6Ue/8KItT58wJnFn9wgr+49OjnddWYZpuy/DV2aQ4PgFDKBu/ZRdDRynccmf3rfo5UKnmYm4c
hBtYL2TeaMLyVaP47VA98BZSV6WeKv/KDJiMpU8CmtUutCZViZHyUt7sxUF/gFjSVzVeYX4Y/WMC
Je1JvB+GKAdNmAWoGQZApNCt+1E5VHR97/qZTj4+RzYJD0dD3RIvYq2Ti8BsqIq0Qxg2YYmk6oNd
KFupgwtI1JmebE4jCaUNuuKUZwgul2s76faTT/FHkWfZo5CVNU8paeiFwM/MM1L0+dtAss2BWAnM
5H5MSgWM/f9DOp6hTKDGBxaZxDMwSqatg3BhALJBYN3qDOsZQ2pOj3/dAoKozpT+P1oClRpxiMz9
FzC4V1s6rrfSrRZ+GW8535ItRNKNSOdoXUMeNS5LR5A/g7gItd8V57osyxnlpP8uqVwBKAalXS3M
YY4vVJaYbrXrDb0wjqFQnTSYBIE2C0hzigmGTyHpankPxyppv8RHHNxTBkbgHI8/1XOQ922hGduk
hMpNI4XBtMoyD9lb5u9mucvrlYRandseTD57466SmerhjV2wnj/n3rrj7lgoL6Sjgf3cHdexBaQl
rpNvRY6n/5nAd6uXsIqVPQ9fgJxuPs6kiaE3PolgTk97WrLS9lGR08zopWcIcCMzBNwFybPoRS6r
RYsYEMnMyQ3UDZAaF8pAMkA4jUtdsSmuJGOpvbHiWmMIMK+MJgxRocV+KUW9jXY6xXT0zhohWLmv
iFH6KJkjceGvmvKkDKH0Gn39BTHctYdbQieA7ykn34c/dNQstVEm8UEBUjGDWCE+alsrCVPMKwCI
A6yvZkMlmJA7qnGgspp4/fCy/zAlDGvS5ibmFB2lyhMdY3CU8yu2DsVuxH1q+XsN3GbOA3gATsCQ
eDJrn9f4a56wOCMrAOtPumSFQbRDE8XwM1QQf28m+5scwsHORIQpYjvePxnJpUM7KUII60huMmpf
4BzXVPhC0gF+kQAXIaQwaLjb61rkZfSwuvdGNoMSIiEFs7H16hXpI3ueKUjSkZ6aTD8yEHkoNh5V
XhaiWXZTLoTuX3n68dnF7RMdsoaLpiEa/nAT2vhYzs1nSRrNFI/YW5GZSmuzXYCVezy0CS9V26Ag
Q77G3OJJIGLXlaNkMpJAhwrYUyzfhxpx+o834rGy5gEHOYQNt0+ktYocjtTT4NRmS9dFT+2f3S3n
/uxspwdOb2vVF0nyEr10RmIkNHm/gPnFrQz64Lm6V/3E8CE2RmrHBUXzzyf8Qufpawk21RycX1zt
TFbTfnkPBibBkjaOo53fLEIGPX+G5dsFCKwQfLFb8dFWaMPNZs9Kkr1e30VAQ3AcvhfGXh5wtHWf
5Z5prgCr2OTiskC1CbltkX1dqRNUGgHRUxVmWt7TkKgZu8atPk7T9iNmrgvzXHmD8fbJDgQB7nV6
ZDx/FUQZ6AnPx+P1Vk8r+q8Q8jBNlk+Cev+YwlINEKUJ3gNW4y+48DutryPVHJdq0CF9fbK9679Z
9tqZPuTzRB78J8kFF7aX2Ks39cDt8txfc+x1iNjXEsR5AW/45MsWg0NCQx7GJTI0zpCyUqhtpHYP
CM3d2KMuxOZDaL/yW6Ku+XfBsmVz2Pj1T2St8KbMiSVXlMH+1P/AIGndvnO4YV9UHNObahmsdY2H
xEy5RWhqePA30HTHmhZxfI321Uytv7gYl2G3HE9TZv0ierHHvGMUflI/5yJv7wzkfaXgiFpywblu
G+VjEyb4n8SnIETcJFUKuGP6Bz4bUlLpDwSMNlmrd5oR2wFG5fXL9nYfYuqnRZRGgoukkGjKDxa0
IGcsRDng6O+DC34Ofq5gY9/TcFWq6p0V2lwa8CxHT/yRvhoIBPehi94gEBVMPrQ/ZR6NqbSTuk1A
s2fKOqwEJayKFVUzGLrTjtt0f2csa0hEkDbvO08kOnRe3Zh3xTsNWCZjWJY8PXV+WnIGieLyRXFz
ll5j5klKGzI2MmTcH0C6qvIcHVvbofUPUNT/CMlXAjLC+d4/PXEmYNB3S4m0PvR331cHQX+YzTc/
FENRIZshOB3gq1wRGtxAlaALyPZRXFE2cvRoLfjzE3UouH+cB44go5IWnireJSiGrU8rtzFSzWKl
GiaNXcuNvPIjP4LxADiV9XryKY58/2vstmmoRON0FvaciwXt5KNQWJr7vzaH2fEDcOl3O63+eNV0
T2zhM8wMJR1amI+piWIxkuJDDz44OGYV8AKs2vXdnX2cQ6HQnGlRP3UXIMRcKtcHlweUK364dIXh
WK2tPdqcW4NrrmuRRtNvvgD9Bh1Clt8loRLOoF2uAgOGbrwClludchc/RSNaqnw9jCZIfVZ8YVNU
0cAtOQGMZpwUYVVwzvS2VfOeGMm5dO5UN2r7Z89xeYPnkEx1m1c86f5EHUalK1hKQi9DLXgG0SnU
pz9VgSjmvNMrrbpLuJuCvhLwzNIC4UIhTq6DEyDQMH9XYwVo8aoN+py3Qtj4an6r0VL6t0n+Zseo
zI0tQu04ha7efR6+paMKMZBNyWBN9TrasJah+C7eFZ0dQhdg9H/VNsDn9Ud05stPcwA3bf/MocM5
yrgrjmKmd1pnnlDaCtkZLAsz3AeZzp8MiNafiK7waX8gGBHaWJS7S93WLwNOLDggXCHFwVAntJdq
a7J7GqbMMXm9r8vOJkKMoKONVu8VLkaEu2J0h5bPu7ZFSqZyBA8FJ/+S1pnH9YrDEMjcJCGK7PD2
m3Q+FtYEmEOrQ6sWR3tEWXGUNh4fj0H80ZWP/8MWHJjVbpZ/z4Y9HP41DoobKqfa8q49n+XHKvfS
vdalVQTeiHFQrHwg3KaeUgYdyTY+ghLQo2T8J4qH3ziJq+C5qClHBIMR5c4mO0QgfNiHoUp4UESe
9akx7SZT6i9MYXGIhPuGt4n41FwNVW7Mt4a1mMKSqN8eaPy+M3Q1tZENwXY24u/ys3JgA/JQkWkk
Lmu1J1cgmnkbnI1Hc078YB9kKCSqGC/DP0LcExc4jp4FSZs0+POrkcaikKAnrGZ7aCp3KYJVGs+z
ZoF61hDMORC54mem56m55ABu2UEBjFcXD/nHAEIZDahS74dne92ICoxCPxgTNBgtypvaV54KkHXq
8EZZhYeJ4JjToZXBLuXJOqyN560ADxzRkl1yTE6nN+eeMcBlWTsD44sisMYXSxaWUnnsUQ6IZavU
MGDrjmFyeL3/Sq8ud4ktpqyNijAboe45YwF4LG9ba4Vt48o9/j9O04W98a+rfAjr2VMNvYCl8SV3
zQMIBi1RzxWuZX7MWWr8DRIMozNaq/yFFSQAM18Jk/W0U2Flr2zOhwi3jpVOTUFc99j+m+hboHrI
03OttscAKKq3YKqB/M8SoLyrlrNQNzRZZXCGrEsTfccXDfSCp1CDS/hxbib/2Je+LF0tS11CT+pn
zd3xIbRwbZRJIK8ytaL6POpbWboQxKDqw3MKFSvlgExF3v7zKKtrb6EshSz8Icc4qXfCuXP9/qXZ
N2Kok+scZlAC5+4UyCmfhuaZlwlwL1iOdrVku6zIeEuSdI3h3RWZUaDt7tfBdmXC5FKscmbkHDCo
6lhLD1U1M5SLfzP7xLyLoBDuuLUN93DP+QSHCTupdaI3CUY0Fd1oo/jDbuSlL7hYltE4iqzAbiQ6
6mZV2ZWlP+Xxgc1jo89wnP71gxofeoROzJyOhttzVsLED+CeVmZkoQ0StOpiHkeikfGCOdTBfAoA
AOjVKyktjiygFHHdZbWgZwNMUnTjlf8cgPehfbBHBUu7kW7rFrjIAjD2AAjJOO5sx3sS6YzCqkDh
EoB4Wy42C6VfJdU8kXr2Fn0L+IjZ0w9h7IFokIa0yZ2KkFOZRAp3CIPhuaQEr2WeruQMzirtA922
DF1T3gMu2JAnKkwX1R1+5+WwVN7ciWnepbDsgKLbztlG+1MGb7WuoF8dj8eCjM6o9Sg/Tp0Emq3H
VgnbDdsNizAKOedHq8mfLndo3faIwX/7FJVYax2WFJoICKRzEEdEb7O7HrRjTyDZte2rTqKeBPxU
2QIvJZn1alZrxPA/Ni7p9unSUfdfaUpcmKBVqSpLgA4KzapVMKa3qK2xXhIxwhgwqpeX2nAGs8Pe
DMm5zqI0mxosbNTarLBh+xE4vZCnk18NAsOfx5Sz2YMZ5Ot0kHxRnrFqkJ/sBuDBhRP50DI1vZY6
iaOUAyBOvAJWn7Et9jHRAR7CPR4rSqeVDZFHpcI/L8BlON4x0m4PfG1asdE2qA0AZlLRSu/HQcrT
FjOsEppouDZSsIwuJyBU6EDswL40DmYSqAMhk3lhgjIMQkxklt3Ho4beZkRiSpwDmABIBCLOrh9n
fLGxTxmozslintQWJkidzqKn0Dxf3I5AKWkOsUOykvorm+oMS9iOqSCdyj62iewKFEa0GKdxft8G
9G7QDxh7Z+W1cDlxC5usC23k2if8W6jmVhzPKBKYfCAINB3Zw3F5mZpIkZdQsbRfDiq/1YePEOQJ
FaR0crGBq0YeYA9HeWH4optHhd6Me3EGiVjRwqpsExumB6hMrHq6NH3r+Subn2zC0f1EAPNWG79p
cX6ORiwhmcnvi4uu2U4OQmD5DYkCAm6E+smhXdSZjrLTbKuLyDR6NwA9E0yQkgzktO2qg8JblnH+
y2ZhOqM+fkSBnL14iNAzSQtwm/tXz/jfnZj0aKid8lBCHSFz/t5HpuC3V6zAxMadX8UWAUFAL3Nf
8fSp7bcflc2Gpzz6wgFddi41OIqrY7HlB7BAiH44CGGlSCsvP4L2+LkvnvWWxvshv6Txf2IaF6RM
p3NBxhVdcZCIOR/sEuhb5lfOAA05whuUovyXMErSglnlp3ULqG2anisNt5vIzyv9+CVKVLIYtVMk
L9XAR/PWMR57Vl5Eo7c0rBAHH71maWEHdu3Q/YN6aVGco+MWY+byYs/qQ2+UFSPgIakejMEPx616
pR0qw7roE2AoSthyZmUydxMDG/12DLHodOX+M7PN0yN05qEuxhG6CpR06VN/iLPGgyiWnd3Cdrj0
j1cRl6xLsIEyJfK6Q1G8OPiqYjn61uNcOIuJ7zPDpxTezGK7vcbVzwiut0ZFtql4i0qIcSxKB+3K
F91wcbeNR11Uz95uA/H16YOAyBw5X4PK+ZWAGemmnr1nTChmXcYnCi07K/wvMNrhYpbPnxMkHUYN
Uw6ao0Xsokzn1nJUD9SznxsrNw655eCacyt8Q3vBWwucyhTR8dFCRI75e+pjzYw+eoTmx+ePU6MV
vDrG0TaQ9hxKpJzK7XQb/NlvwLUuxTD9rXhqWbbx7BqzK3MbfBZ5gxnDskbILwO3z2yi6BJi+cSW
4/DpEwMBYy4HmDkHTeZNUcsNPRtogjdV+mFW8MA5GXiChQzsdC8Tt2gRtqxjgfZ8zXwFptNiE6Xw
Rr5sI63MEzSBvgdZ9kCalOROEWvkvcSE/WGi91rCTVcKv99hYTXdkxxaX6pOuVXcAMTMuTLkpKq+
xkYSMU2HxD2PZr0TBWQqArrl6zMtPNyqq7thCQbg8EnyKyra48yDBqEZJefnPq9Nr81FuGy6DYMX
9vFLJEApeVCyYKBCtYQ6aYbchsu1HtVLP0f6GmXiG5EGgIdOVLeOu4NP6z4OlmUBAoxv//3Sq1g6
YqQSPxJ508pTPm+HMiZgtIhMH7+jqsKaSf2rZ2hYO5md0340ue7GM83Z9DlYvPgQFgPT9PONaSZ9
sWUrrTev43RVU5iGXPT/xttJVTuaDaUYq06d4I7ASCe3kfenyzZ9dw1z5D2GE5LUdIDdj4jDl7BU
kkgwzRT8mEs4Re8ioZstt1XwwOpUI7oQyKsudKKneYd0YfrzTqEesia9gIh8dvLUEPgRU4M9gpwX
waez1Ao+MMvEq1ahvrOea2/5KuEVI27hz1ExHhbYcyc25dChQMw3jlHCsZGCZDKu0EEkmDe13NnA
X6RH8NaEIoHE5J5dPTeOrtKaRjolrY0M7qr+UeuDoetNZO4/Iva42YdxmPp+KJtXYJovyEYipGKV
XLvzRmDVUSNCV70SIzV2JQtD9iKY05Lyx1sL4YkgUWDDmG4W9QfovDngo8BzNneoJ80nvzHV3lkm
WmoxSrJ0pYF0uXm30eRXGZw3wfde4wiYgK/N9WCFG28O1He3ZNKImSAdttkD43ibU/fTVSnRPdsV
pabIsRxjbBf7mD+5rQ6GUe9mfDD5MA1b43FYQXvBlo9tt65Bcvjut1c/isAfcInS4JAbIvxq/9sW
W7AUe7dGymbOgPOY6sKMbJh7HtZyFuacRyD9j9KdSrtwYvWJjYiDvPkM+nCMbVWWcpEsYrp3TSOn
AeMUasLJdsn1TIm3UxZ+UWzZHPoZuJI2GqEjqrQK1GzJ1lMD36oHWR+4T/FZaAoaq+u3QPDUmRlx
GOYGP1US+DI92e9jcXzYSV9q239IzGYlLk3Ub56ngFjayM346hzlHds3jITUuuu6L85DSmrcMFgy
C+cuc/VJqUGF29Vw6POHM3Rpt/rWjXnBdi9NSbg9A+VqJZ3ow/EW9M7RfaTUP4zaaE1aUPBbwVeZ
7E0ZcwLpz+csPviw3wKJjFG9MdVbmn06eSWVnRyr6QFKEqNbWrdscERHgHBwXw3mAdXVl74i2RdV
CmzfwSepz/Fn+/H7JEecCdciHbTFrVwuEpFUOpPECGgYva24WPkASyCnEeeiqW3f7XU47T02kHgO
Z3JhW9kq85MADYiphJ6Ql/B4oINyANFHMhrCoga9ERUqpXpsiifpSPBvZYysaK8pi9y7s5xSPDpg
jUuQlq4qTcgdbic/V0vxdrXxaOa4QkG83G2xBgZZo89iiQbhBWiqTpVZv27n/1M8477DaqJXCOe4
hXqyQWCPhrmQflNuo7ma7LlhfxDTj+gNF3eGThrO8r2G0kZjDaazdbkv1DP75GKkJKcS9x9OuruL
pkl/Rcaq8bZBos1OqbRwiuibkTLppjy9y/6z7sk0xXBH8O7/QhJqrWKcxZCkD5vC2QewfF8pc4qY
cafAu+Qz2KwWI7oow+tK8o+rxwzwVGe57gpAuE032rFRKIBWQSnT1Ub/ZPjw
`protect end_protected
