XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���cJ|�-���8���u�'��Q�b��6hX��{�J����R�|��&� ��%ء�N�B���*"��؟"�42l
�t�<}�;n�!�u��)B����MTԘ*�tm�4�N�Zx?����vА'�|���Ri}����z�d��2�G��G�R����e������c�̲~���<= d	��l~�s�9AF��ƆW�c9?\��f����|b0�ׅ�"}��~��ya�6$Y2��iZ� �s�7��|(�T�����������Djٸ���۴�ZBT4�a;B�87?�hO�q�b����t]49n��q�H*aٺ]�M5���a��	vݕ�_lW}��L���vWz7��&�i6b-��
���3g�i����Xq-����+�h�}������<H�b��
�\Y����G)�n#���R��%�`�-��yР�> Ÿ�\ڹ���70���3�N�khn�
�[���0;"R����_,U`14go��_v|�������5O�/�+{��gb���t+����kA n���i� �cT�H6��x�*����� 5N���Ћ�p��~^}�d0�^y�����e~��ܕ���>��dAIk��x����V�^��U]���G�h��)��I�lӕ#�ߓrY���8Wg>��iWdl��>ͣ���f��]��Y�|��+F�J�d�f�R���&^���o�M+kl�z�e�ߣ ���(�C�y�D|�c��ˬο ��*x���_���XlxVHYEB     400     190�F�S2Z��������K���q��ȺaD��m�����&������xo�/ZBH`�l�زsB��W�\�q��^&���<T�ɟ5�~L�v��ws��K����i�uη�T��j�M�������2#��ʦ���1!	�CR{��༻-h��9wH����t��^����'�'B������B ���a��������c�~7[El1�E�1"+���a���Qu����~x+�i"��&�9���ZPԱ%�����b��e�7D>7�+;S���u���'������WJ2*�턯CEX��VA�z�SQ"VF����ɂm�;Fc�:Y83?m�Cn���aF���-j^R��E3g�0���������\�c�g�c�:DP��qXlxVHYEB     400     140T�:�|��Z�8�%���پa+�����x�tb��x�$�ST�2G�14�M���G�������'3�6XCW�h�w�.�$f'���O�|松QhF�#��v䯡�F��q h��x�yy�9f����tHf7Sn<��G	�)$�٘b���E�)�t��<;���0�p1`�i�VF�t+dCM�?�[��3)b�e��}�iы�K-٧��~���lL3����{8vj}�G^Ӹìe���%$lK���/�� �.Gf����˛��W�6Hypz|�$�:x���#�)����R^����f��) �X��`ӝ2��XlxVHYEB     400     170}#�ӄI� }�`~�H�g��-���oժ4:��l��H��k�il��$\��l(��3qs'�xMn'��}���E]��P/a<L�ۛ��\>.Aj���~�^�����YT����'iK[/��M6�u.u�zz�����R�'{ӱEE�_GM�D���-�:{-A����#���� ?�U�~YmTG!S�i��A͎k:�5�l()J�T�kiz��p�p`���:�.�Ɵ�#�}��f�us}�a�}��K�$�j�K��<�`H��4�4��Y�sO/�U�d���$%Nn��[Y諤�2&�-�A���;ٔp"�ʊ���Ƥ$�����
�t���@h��d��%Ƣ.��o���Sv^�ƪXlxVHYEB     400     130gf�� h�~8ę�6Gߋ��p��e�W��h+d�iѣDU��2Q�9 3�������,1n�Kؕ�j��E����U5��,<zy����q��]�vT�=�/���g[��W;_7�
 �$1�{��)<��1��˕Y&�m��weH��h#����g|L��������[��sg�q|�����~�x^��D~i/����9
9����,�˜� A�� =��$����X��K���к�����Q�{���d���Utlb�E�9���wY?����u3����oWXlxVHYEB     400      d0L���U�h�ҧ�m���6x㠽	|�<�5;cL�k/�U�0x���n����:�-�L7K�Q�>8�(�����N�p�m���Bn���,�=$��C�Ց���]��\_f�^����k�IcZ�[q�q1����1,�Ԝ	]A<N����h��z�`:,֊V� ��4����'�+���ŏ"����;yJ��S��?�~���^=PH<�"��XlxVHYEB     400     130 ��fY#Y�\��:���AC�����p��(G��Gpݐ�(�ǩO�Y~(��e�BS�v���*{�U(u� �P�*�b��uM>x�a��IU7�U�N�C�6�?�a���H��A�� f��EN���ƪ��1�2m��c�M`f����^+fY�^
�>.&e���<�Y��`(n9�;A��'m����Љ	���&�=�
�cIhwwH�;@Z��[]XN�a1�#g֫�\`��#W�e��*����ع .�Q(���n�d��P�F� ���,CPDaX�tI�wI����>��z^��,�ԜXlxVHYEB     400      e0-q�LY
��9qзn����,Az��ONt��K*�E�c�7v�7@�5�Jj&$��`�иÈ�E�щz�Q��y�W:X�r����\?�������$z�ױ fT �yS?a��0̍+�/&�M���������:xSMǾM��Y=�z�S��9�ͪhς�)�9�D>(;��R�ڮ��>'}��%��sWqCW�N,6����UngF!o�(��:�߀GO~́XlxVHYEB     400     140�c��o	羲�ۮ�F�9@��1�w|��,���l��
�7�Hk�7t[�=�?�I- HIDV\-���	j�
?��d�b:d���`����8����i��(V=���\�޻�*� ��h@rǥ�Rf�ڰ�4�"G��H6]�ө��tݶ�$�H͔!���^Yl����F$[�% �$Hj�G�O�)V-K�/e�[� �ċ������O1i�üҨ���B�xj�c�H=���д��d�4�r�J/��yq�~�u�?r�.�'O�x��{�:����X��JK�2]2;r!�z�Y������W�XlxVHYEB     400     180�����u�-K� Z��(��h�҆N������Y�`�~"ھ��m��;XR���]@2��474xs۰�>nq+ޫl��*�(���y04�C���dv|��G@�5_Cz6��U�DU҇CA�v�![m����ߎ2鷤j�[R�����{��Cp�R�q# KZ����V�L��c�و�V��SW�w��K��F�TI���b��7�����!1�Χ�5�CS� mvc�1�Z���B�ō�.zw�281��.H�M6F<[b�j�����c�����'S��K�y2����(�G�.�MȺh�&�p�c���U�]���Y�di�@jE���KM�uf��3<�\w�>�wT���F��N������,�8��谱b7��XlxVHYEB     400     150����ؑ�l=���K�NB"Iu�T��
�0���!�*#we�y�m2*�`���������ۻ���(ō�D�nB�OE�:2
��:P�wY����$ƚV"�Uj/f����3��ߺ��[�z����u=��9"�ӊ����(��`L`��-e}N�7"�έ2� ��\9�ǁ��i�5��}�(�f��1��ij6*���kR�.�IL&l��2���JW� ���d�*����zNi���c����&ʕ��I�6��\����k(͟kO�~'߸q��H�1-e~�_
Hx�D� �7�&�׹�q%|�V}L�Őំ�ژ�J{����3!�XlxVHYEB     400     160��G��b�6�XR�g�L�}5��H��J��\��e	�!�0v��E�����]jp��U"w��!m�.��Vu7�x�{��π�	(3O�m�M#� �z5}���Ѡ��M&�QFMG�s�%]�ra^� ���:6��rw��^�w�m\N4��[�������L
~t�w������x�ه�t,��^��{�W2蛑�>��g�k���_%|ܤb�߬�\	T?�!6_V�	W7)c풢C�p��@�V,-d��+�1�����"O����s;�&Y�|�����������qЋ�7����)�?w�فSH��u�<����K�*�Oy���^*��g`���Ap�j��rH	XlxVHYEB     400     130Z�g1r>.����^�T U��`�:���Wc-S�ʚ*s8 XI~T�[��P�Zj� M��wk�w�u�c{>�X��z�4B,p -��r�ZF������;P���z4� �RH?�i�,!zZ ��%� e4bpU�w�p��m@_��R@H6&����K��'�>��oK/��v�؄4�S�D-c���,�4m/SS�Xs���3�ݸ�����h���wfמFY�i�B��`����k
S6����c������M_J��\��|�ydD+��z�(���a���_�`d�rluhGAj�����3�XlxVHYEB     400     140�,}�C�����d���+�ww�>YxeX��!Ï���^�0����`�~�ԏ<T���Y������h\�Z)V�P4١��M�B�'��W�K�h��S�rV�}�n�Z��u\��P;L:�H-�~g�<h�ʵ�h؀�Q.���Yb�r*c�x��M�?3,xV�X��v�[f�g�G����U\�d�:��=�j���؞��G靕�I���2�l�^�+tfEOH��vnp���׿�b��+��۩��>�r0}l����!b�U���K����hV@bkK�ӗ�YφS�49tkYS�*`�"<+����aLmXlxVHYEB     400     1a0=���4�n��D�)�FA����K��#�����Ի9?��Im�ⵓ�#7:`F��ӫh+��;m�
S\�C����e�S��~C�4�n�[�@�r��<�� �sJ����"���%�����c�5�����j#�U�l;�z�Fq��������i�ׁ��+�흳�3FM��>�iHJ 8���˧ā�����z!�U�s��c̼$���P�ٺE�>n�^�^�>�Xd�|���a͞����t[�|��Q�i8ҶѾ圶抹�"�N��𱱽�{3'E#D�4`��ꃑ��}�����=�]A&�����y���m�z�F����}��H4:4��2P�&\����
U���,����
�ٕ�a���?]�j��E�NL��C�Q�~ȩ����U]�6��Y~٣lXlxVHYEB     400     120:���N'�>.��3��(�h���f�v9�>�S�,;��$7�j%�n8\0lp�D���ٯ�{C6����c��V|��qZXύOI}g���_�b�]7�����g⏈')K5�"�E�B��4iq�83���?�Ԫ8qls;�e�k/�a�c?pټ�J?���]�c�v��VI�ɮz����t�ʦ���(���ԉ���j���U��l���|�fZK�B��{{j��O%ք��ZCUW�ߦ�ҵ�{�>9a�G���_Rج���(�4�8��+�XlxVHYEB     400     180��l�IB���ӟ��ٚsg-Ɲ�"�'f{{�qaU$�ż�9�
�>2/1 .�C�����g��y�"�$��V�_�(
�p�;�fv*�����jP� }R��P xUk�6��Q�TC&�|�����!���.��?Fؽ�e�\�f�##I��3:%�͒Y�s�|�\��`
�^Ě�p��(:j�L�su"�A��Y�ߢ CV>�P�pAn-�$������P;�/�!Gb���c$=��ΗU�49�H2.��W�v�Q �JF��4>��#�U��q|�����H�)����W�r<V�k��E�fJt-�3�����c�~����><F�d�(�D*�糌��C�*j@���2k����3ʌ�oa��yX�XlxVHYEB     400     160�_$B��Y���,1jw�����-d��}s�6�)�r���0�Lº�W��r^eԟX��mQ�O$��U���P��^ǻ
=rT�8ޙBK��t�ѯ�9�.+��#=}�v{�#рy&�&D[��O�9��DT�2����#��D�a�\��!"����4P��g����F�I0Z�&'�1&�xk��N0��x���z}!��J:��U����-�{��[�A沤 ���v� ��𱉦
���0����7c�<t��G���لgC��r܃Eɹ��H?<��ǤX~'ʤ��1�'.Ic��~�V��<�T0k�y-��VY[t3�3�U�'�3�>Uh-x�2����-Iqر��tXlxVHYEB     400     1b0'Y�"ԛ���M���[R�j.O[�2��o|ɨ�(㴡R�,&0��³%�xN���$2��0h� և�J�Op��IZ���n�Ȓ�VB}�*؀����e9���ĺkyM!�26��A���N1A����eNn+Y����A��I�5��i�\�Ȗ���O(N�-�>5]K�v����w���]ܴ~������'�	����N'Դ�^��Ψ�����g&,�Mj�d�ay8O܃�0�D*��Q|m�,��ۺFļ��=v�i��lù��n�!�E�2u��׻2�<Q������=�;)D���P�猻�e����Xd0`u�I�c��r2}y��f��f5��::jE���'Fw-��`�׍WI�#.��0�^$��BՀr��Zs{���@�XaG�����K0ŏca"*�v�\�ݸql�ڏ5pXlxVHYEB     400     160z쵞�%�<��WXIs%�5�O�gt��.�h��[���5Q8��mQh�������&�Z�֊e����잰��O�7�iZK�hՈe��3��e�T�#Y��T��C�'���~�]w^�|���S=���sw�y��\gyi�'un0�l\7���ݢwC^ j�S*�nQA�,���B�5���|�]�\i��b�G��D~Ե{~�j�" W�&E��Zs�����7$u�_�Hyī��@�T�%�ɏ>�Ū5j\�SA��c��F@�bձj}e�np����[F:�H���@A1�c��
$�� V{�Bxr���R��L/z����Z����Mb�>��
r=\,�z9[��PXlxVHYEB     400     130�d���+����UV�+p�I ��91Uc�8Z���x�{��r{�wy�#�ED�2f�O_����Ah�����V���e(�>aZ���i�s�d���rK��w�g	�V��֘~�#Q,/�����i\�d���ۆw�*�	L�4_�&2tچ�޵����{ ,E1��a��s4������1'QNX��U'"����
~ɓ\���N�6�]���IR�s7�f�����0��DN�JƏ�p����woK����}��f�G�y�J�����ފ�����t(���c��YW[*�<�Vh��{[l���XlxVHYEB     400     140��r�
�Ih���=f]��};�� $��=��#R륿$�'1�\����`��'Gz[��`L�ᚕ��Kv���oW$$H���� XS�;ٚ��QE
���(��h�9�Ub�&f4���I6���J$bH��58����:�'.[���m�jA� \�M�Y���Α���3���}_WT�
G�0����$h��-�%"��{C�܆�{p��PQ ���j�HȀ1|J��@�ʥB�L��{�2�CT���i��� ����a쥗��C�1C��S���6�&_�\��$���Vb�˳�^p@MZ��c�W���+{�/�XlxVHYEB     400     130����tK�*�����]�_G>��h�{E�z,*���&��	Nb��&`\�6�׫Xѻ�=�)�K�+� ��c��(F|ս@"#�A�G��y�sD�*�0����Q��!�wy�J�X"<�['lh���?͉�|��
��	���ҹ"��c?�w;�I������_)�<X�G7�����6i��Q�>��ٹ�A����k�~f��׍�5���.���?R|~o|ɹ��)kC���U�����D�lV��:����A����`�yͫ_�B��}�X�R�[������rH�;XlxVHYEB     400     140�$֒3�f���DG(�IA������6Ϋ8b5q*(�_0z�l	��[��m7���b���ѓU�5�֠FAE���2���>��Y�ly�հ ip�ĥ���v���+�[��Շ9*J�2�Ǌr�CfOVf���,^�����v`	`}}nk)<.f�Sr�9[�4�ET@�U]]��/���q}�M�퉫���ؤTz�$�Lm�;�j2<PN��w�V��t�O/��,OѨA,�����௥�+U濥��R�dkv���y�{�K�#�}�2Ey���N���"^㛠�&��T�E/]�QP�Hm�*60��ȝ2XlxVHYEB     400      d0"���Jq	�uBT�����U76��ިߜ�1�2����I��X����?�A�v����3fX�IPΣ�� �6����1	�FS��]�lY�D�q��k�Q���� (` ��$B��鏻�
�����p s�_`��9���Q��+䐶�u������Ex���{��&{}�ӫ�ū�E;/�Y}�D��I�mo$�z6�+R�pXlxVHYEB     247      b0��x����؅y�@�~3�*l��n\ġ;������O�]�ƀy�rѾ3+t��࠼y��p���3&nϨhX�>�/vjeM`�*S�Z'�~��;��4���/zj��;�U��(�Ww�ᦓ@:(\�e6o��v�����m٢�Ihi��W���6�PJ��:n���FҊfΎb�