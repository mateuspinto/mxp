`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
IzVqqBWrsju3r7uN9ilKFbYOx2Xi9v7jI+ncMwZM8MhO5HE51aBeKKdhoHu5H4OjvihdMulARkh2
d2FsGLKpGatUGSuRG9dMCiaV6B+NOiNSeRr6zKUxmXQwJ5nmX6pAHq46zJ56Y8hKAcEEYo7QGtoF
xaEFU/Btem4ngfJm1hmrM791o9ZOGmA+Z8GKRgAr6HX1fIII0FCucRYm3jwAdaPCyjhruMDVmsqX
ANhMZrk8b/3I0Fk1xplqPHlR9sDWsoY96ZGmEROnOutCAkuNpP2bBzDy/L2S1hLepkd+/11P4AAc
VcU0SJJK14yg5d3EBjQL2hvxhJyofC1u0hH2T/y6bT466MIwbGcqjnS/sU2WFhwF5bxF2sY/CXLb
08ADzZ6cKR/db273ceVN8pLzkb1ZM+UjfZaJqNfy3B4FSut6GVqvvqdJdbKmmWIw0+WY/WbI/oec
nXcqqYbmfmK0vYRRty1/GQWbwkvtgSNT1DNlICzFM+2jPlHnhHXUIWQSUvoVySaucZh40YiFKJOR
igRSzkcsFGaSTxJAuo/3je2LmC5kLj60anvkm+9L2JgfR8eRIDjYMCA6/fQtNbP8Bxm7amy48J2c
/3Wlnbe05bl6nBDX8O3WXfOtyMo2veI7VoaPKxPhFTyG3mPGqsjFvdfSMkPFJBrHVav0IMsyO8Ao
FGFjJ/lzTkvxZVI7i1uTAsbx/No0B2wTBp7ONWy3sh5rYfKXNbkU/JVBOV+C1UtTsX6ufGqys7KG
bCpKr/kI2ljfBBawwGHZETDeNSmqE4GBsy+KjRKrhU0/JGMm2HRFm9p14bqWjPo9Ir+kP/UDL1bc
HihLs7Flqag0+kmF/8zgxD4wxFN9MAyWkeSuyaS8DFJDsxLCRU3DL8BBuWK7l2D61PNM1c90e6a8
hCA+SKbD5qWMJGJoi2UcAxvKJJXFiXN/ff5pfaczjSexLOx3I5gs5BnFRl6hJrZk4BpZnom50+f5
QASp6kpaHYBK4VI5C2Pj7binUcYGypYXIBhRpWjw7XjN7yQExTN9zETSOgiCMr1XKwxAOp4STiFn
MPYOoc/ZnEIVyFIgHtJXy4nnYXoIBcT8IeP7fLRM6Trt6apRrcyM3aiucWnKc2JSlAFbdbxObbpD
XtkntgBatnnFpGA6iN3JLNyH8nNAWcgiZzDgEMjfdF4o7NnJHB4q2Awvc4QmG+PaYJSAuVmI1/ZM
Gy7axn0SmPXn7yk8sHeLoWcTTeZc41c0TMnoMs+5yPolj2FaImxFdKGYFQsCRHAlfwvw+q2r7+6q
VVKS+D7/uYgtuUIYHguZS+2bodWNgWB3N3otLFY19rxiH0vxo0vQdOhxZrAa+pUIGN5/5kYoNvqw
MnNon8GFHn3R+9blCL8yvD6sHtw+5bMlnwZqLS5eIuyOThKhUJmcL0eK/BCoTz1souN6ivSVt8jO
5jfzw9BrUhlJVSB4HEqdiZ1PqZ6okpcZodoLd/Qzf3EOS4GxsWBvVFgYNw1UCZzkgD3nPK/0CYci
Xu+tZ6Q7BUcTPIAZYNTrdagi9WRsmd8GBQtxEEYimg+7gRGZ9xHS39QhkbWLzG1p0tulDeSbygRJ
HDtSYQ6e6l6fU62DzqxkTW4UW1UgaaEYyCHmKXmN+V+/qrSLglLjmK+R2XWmBOfIvFYWUr7fr4Zv
Ap+ZsfMEcRzzAo47tlcbNZ5JYDSxERvoKSvX6403QJOk2YfeaParWv0SMgyn7zOJQHkSPAr7qJyB
40JTUrla0JxloduG76IOT0ykfvI14yQhruqumijgPtJTK/NaEvTBdQ1IuhQBDIGjSESTL4la56Mz
MPPJZwT0dICVGQ1ywLxvfjephH275/GDf+8B9/g3DljmTcbYygbxDbuUmond7mQBeEp9okGycgPL
YPN9bCJLy6Wq/xEZvC6v/Ks9R5xZ3tgyLJ2FBIBJS8ItJ63tiCNS9ZlvB01OpenXnLOJ5YKhLjC/
B8g73npsHfxlYefytGOPfbsIu0Nm2/kRzt83L0F95s1bXb9Eq3B0Vom7gZ2NXoW50BL6E3fstfbK
iXudZKq5xx710AYe+RSXrDbVIMOVp+if4fsoVNVw5SJzvgI834dDePhW+2mP
`protect end_protected
