��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���6<������LA�H��8�ڬg�+7�z��ϮO?w���b��1b^�b�
����+x�=/��.o7�D�DsCT��EN�@�MPp\�ٺL��S��~.O������qN��������$W�,�)M������Ef�-��e��Mp^��.�_-�C<�/�ڶ�b�b��Z|)0����;����V.7���
�m�ήzum!�"��*0�Ƕ�������i�M�,ƙ� A�̇ D�����1'?�nEL��;�N��t|����i�XOU:����P�]�*����n
�eK��%��)͇���5	��b���m�׀K�Rt�(3k���s��n���88�↮�ug�i2ԛl�C-�z���d��J�Rѝ�'��|����⚩]GQ�M]-��A�A��[�5���y�ל�s�X*�zzE�k�K�8A1ݪ���}�,q�I,���J6r����%P�>�u|�iU�����O���x���-9Y�y�ГKI�(gߣ>Q%��f�&��5��R��93)Ȣ�IV(n�҃q���Ni�|̭e�����l��  ��i��ݞ��<{�m.W1[��7YC�[�ݲ���d����'����;��C�j�r>Kb�<�=�n�(����Tnc��¦v�Bb��-��������əmZ�d�-a��`�0�g{lJ��X������qJ�j|伆ruN*2���}q��9�zӧ3&���l'o�u��:m��=V��e&�����_vL�7&t��2�'A�h¨��`X���\Vi�V���y@�n�	��H��<��ݠ��]9' }3���j;��,E5M�� =ρ��b�������
���O�bg�ZVe/�Sԙ;�8))�@�GR�|�5t�J�}.b�f�>�4ܿƸ������ˎ�"S�[�j�,�i���S4N������*��������c O���1%��gƑ,>�v�ZW�,������,��w�	�@�a�����\t�$pn���>"PsFY�D�e��Λ2Z��G�А{@��,��Ǫ�Z�DM&l�������o��.�h�\g9��3� ���&���{�7���ZEto	H�E�N66�b�Uذ?�$��}��s�څxΝA����o�1 \��)���`�8N*�01�o��6^��D���3�.�1Eu`�n�+yE��zn��X[�[b���`�8Eo�ݍ�a	�|7~R�X`!\�<�H����S�0sBof�DU���: "^����2��Î͹'0l@��aCr�_2{���u"RK��Y��9��rH��/}W�2���|��4Z��Ur�]��;�jG$q�b��L��
#���D���#p�-/��ㅛE`����!�KBe�`(�����~�7�#���=�*��f<��E8fMs���*P�jԤ �P�
"t���s�'�]�U-��>�W��@����Jx!�w���%�I�؀��./jL�S,./�#����2�����X��*��_�%6�I��bo7\[�(��?ğ����๱t�e�C�c��C�_.���M#i���sm3�]�<&z'���x�̛څ�ю��Q�nz�&�]qN`�g#�]ؽ�����|�O.G�)�C�V�L2%N0w� �q�b�r�g�j�l`ZX�L*[F-��ϻ��K�S-o�,�C��.v6'�=R��:bX�:�=$uD8��ǃ�!2N�K�B�������p��7�����8e�^�]�<��p8v랬)Kj�1�-h�j\`�"�)��H~��p%)w�[}y�V�WA����C�HF��gݟH9x0̌\)�)��C]K�_V`wM*)Щm��k�7tpͻ���4�9��*�oc��ՠçp	c̝�3�O�&�pf5���{U�h���$��3�H��Lo�}W�;a˂�j,��@�H�U�@����Wtӻ;��V�8'�	gp2Y\���%��t�r��/�q�O{o�6��U�͍ P�譺�����^�1L�x�������Y%9�p�8����E���P�a�Z�yП��+�W X�W�͍K�#Ƃ*���rg������RO��3ڙ~�އ���s7��'��c������	\dG�8T�W�+�/�VRß"_o�KBXD$��8���Y�����k�X�Ӛp,�a��kѵ�xZݑ�r�׊��4������34��jJ�
�"N�ұ��ŧI�r�a�+7Y�;ۏ~��[!��Q<�>��&CegVG��)��ST�����P������'�(�ZH�zsЩ��fD�6Q@~E�w����)ob��,��u���IݩH2M�~z���̾�4e�8�Z�L��Q��f{�U�G�u3t^�����[q�#��X}H�	�����
�"}�±��'���~�9����������� ���-�`%�~�yz� �֒�έ�*�����%G������UU��ɶQ����ܵA�GD!p�CI�J�瀩�^v`��`�Ur�XI�T����ڡb�}�h�Uy�|����w��?<ͥJ�������Dq��]���>�^0���ڣ��x��TS�@;dJ%��Z�M�2U�]"�M��h_O>�!&�Aq�!�7���NK)�bw�fGw7�����E26��|\͞�r���-� P��G8�?h�s.���ĵ�ct7���q����5C��&ˍ�R��	h�R�;'�j,l��Q�
��Z�\n�l�=O�'�d�n��������0��-=��K�]�����	���Q�#l�8XSSfH�,�����ɸ�
��P��]�[���3gLY7�aҭ��.Q����F3�U.��8�+x�R�F0�S��$��h.��g|�B�20������_R�0"T���^��PeGw��}]q����<$�!8��X
'{5��֑�y����V��1�����J�'�;!(�S-v/N!iPS�tĭ���m�3��� �#���3<4��<i^�qFI�F&$���?̵|�Tur��?xG��5b8��"��k�����`-u�|�\%�.D���P~��������T��W��"ΆT�A�C������LD�(�YD��k
&|�[4���l}n��D$:�
[K��cu��W�'��_:�㱍�ɞ����vYŠİ�}Mt��i��\hfd�Cc����A@�u�#k�n�g�j���>�}Jǟ�I,|��칇��I�R�BHH~�5�Ѱ���d�+J�
7}��D��J~��Ⱦ�0�;�<��8U�aJ��^��#-Ī���ɢ�N���8CA�G��_ru<'�\�xy���xӀ����s"��;EC��|:�y;�����ĉM��#]D��<����'sF��[��Y��3��%P6>ϳ�Z��B#�-���C	� �[75u�)3�r�_��r���J���?q.���q_5p���� fn�=�v`F�C��J�J_G�6��:��zj?��au���'���ǘhA+F�?��K)����:�HV�/����Õ|����.�8e�f�\a8��Y[���g�x|�E��@%8Ň�������Cӧ�0��B'�ѭ�^��W~��?!0�}��-g1����H�4�vĨ���H�|3+�$�S��t�,�i<�6P'}�`u`H���?!��*�����ЌS$唉 �
�c�&���;�']@,>_TޅĽ6��)Z���D����Q��>L)�W�Dעi^Ҡ_�x�򼕈6B��[�yc�(�T�kz� R�^L����K?q8 �Ȣ�"�?�ͦ^{ �e!��BkMB��;>Z��8���'�:yS�[l:���$۩<���E,q�8("�+W(v����/K���ƈ��߸H̃���t���N���i�p� �^�9Bs��;!-Y"�3�dM����J������v��?�2H�R�%s8�A����Ҽ���j�\�]�ɧ�8��O-3 :�y���I��+A����
�d45� lINn���UC��\���Q�����Eߢ�@�n�C���3&���D�� ��}�W�����D#�+0��?<aV����5K&��`������]�d�!F}3���L]^�&��Z�W`��C�J�w����6A���9n6��_4�?V��Gjo:��s��69��xc$=���ʺi�������>_T�����ج��b=�� �A�u!���/\�y7��m?��^�ǯ��=z ���̝lՙ���䔥�ak��J���^&��Kf:�������CG�v��D��E�!O+�����n�g�E����褽���:Zl9Vk��u��{rK�&�)�D�]�zM߮%7�E��^���G�}[��Ds�����o� d֭�$��d�2>�'�A�RA�n)��5KYVu��6���%�G,rQ���*�,-�ɮv�Ɯ�H�Lo�9m�,b^:>/Z�.����/%�)Ϫ���۪�l��yE)���i��1g?W1���} ���g��]�F�xV@l�ל��weV����p�R�����ҙ���`3�XǊF�F�c��^���T�(��)U�Dە|Ie�1iL۵Qe+�)�#�Y��%���7��C�X���S�`թ���:Apv��0�qDf�/�3 pl{/P�
e5�ޘ炻+����N��(`���ܭ�N�W�[�a������=�na)���#�c���$@�3���7�$�����I��W~u�|&i��9&����]Q8���NyUX�����~1�Mg���n]k�)��O�����[pD��&�԰������ئ�����㳅�,� 4&X^���.���CN,d�=%%�o�� �������t�[U��8�*��f�+T!���
 dW��	������)v��C浇�㩯;v|\hI*w�z	8��FpN�{�j!�lt�Pq��ѓл�Z����5�\Ͳ
#Sq�L!'���Wk��QW���$[����O��� ����i��?x�dAq1����*��k���ON���f/���<���=G.K����6�Q&.�?��\�o�IԡZ�z�_���.�L�=Y��i��I�^��Y�#�����5��B��Gj�|?��i�O��Uφ�-�r�0|Z�#b#y8�U�F����לZ#��,�j6�W��נs�� ��p��KB�=F1b��Υ�����s�9d5ɵ��s��2����W�v �^�/��Fk+���g}N���y�"UQn�@MJ��gP�� _�� 7�^,z��}�Y7z]#^�\6�ȷ@%QJ$�w#Dx~v� 8�!������Qc}��R
F���^�N-�܎�dm�sV���[�T�^3���g����/�[���!����{���V<߾�f��k�N���fM�O�<���b�� `uP!��¯BX=K�e!XӾ���@�\����7�&�w7��Ҹ0տ<��������̑���ޞl�D�֛3��y����	dx���⑏�n���Bx�wD\G k(	iB	�i~�yR3��ꕷCA�ކ5���c/�;�����/I�g�o���T��S ���x�~�����sO6A^�H��"ۭɀw��z��[��=��&�dF��ϵ����L�줬5�D
|%���h�MSu�n�����:��u���)�U$U�(I�����~ܫ�<Z1&�H �{��Ks�����̥�hYS�n����Z򩲿.5��[�.%�M�=,rҾw}���h%�b������ǟ���%<�4(�����`3�Nz�RUW��մ6;a����)��ȷO���'�#P�h��:>r�O&a�9F��$����È�����I�� ���4:h�-��i#�N�6\B}��d7�Gڬ�a�}�����Q#��(�r=É$�M q�� �;e�D����D��P�7�`t颞3עx<��@��.��w�D��!|f԰� ԅ�w�(�P��1ۡ�����J�yq@xX�S]t�1!)���.�'B�.��Z�ĢΙ��_߸�9;|���+K��d�U�dǷ,��H_��h:u�ZuGL��;�zRO�7%C��Z&�8�*��9���Jx%ZL�2.��w��<TB�5}o4$g�ih��ϡ��S(���L���[���q���5�,gG��q����HRUY=�����⺙���.e��!aplXQȢ�Y���%ò2�*�&[��r�u��PT�q]��g�Ķ�v*��3]����f?8�	�T�9�3�,ɮ����|�{KB��Є�D�dj��!q;t���=�$ NAsbg�WAi�V�c�U���5�*�����K]���_R����7�ҏAafR��"?}O����o��{�� 횆��L�Q �m����ʖ�HV�evN9��Q;z݁���D���*�@r�R�=H�H �<3�)U�v��/C�T���K���c7������8��A�g��Oi���4^�!�-�l2�I�\vSd�v�Q+uk�ǖ���������*J�,t�y������\��R���E���U(�T�v�n�:@fM�EJtU&lM=�e�=�t^ �FQ�
�S��^=G����4>��� }8os4�vp︦���̼ׂ�oE�9���Mo.X��bv��zh��ֿ`\���b6�yXL��"�F�\�}v��-�2|��c��OB�x���Y�$���?��y� M�	����Ӫ�|b�������d����Fr/�R���zԺ$�<v�[t������_��k�w�d�� �� ե�}d�x��~�l��9P1���,J�+t$��6�a9��{JL~� �aU�E[ݗ���>��d?GRkd�b���jҶ���d��H�2]Ƃ]�3�5�y�*3.����+܄v���z��}��L�H-ȘiWm):7s�1T���mJm],X��ے=B�6�h��*�IL���H9$�~c��O������b�������m���4͂8�s�BGq.�ƌ�T�����^��}J �GLL�-n]on�Gè���4�M�56���b>�g�a�`�����[3�}a!O�ov���!GSSm��W��4ez8U�3��n�A��0�H��uaxU}\�oN��� �8%w l��O��۴|܋@7R�8}���e|�h��x�j�E6��7�l�B]�\��ʤ�V
}�k����&�I
����fg*��8�@��	t���4�O6n5ʜO}D���_��|�X�Ǡ^
��^���~��(�mV�[}�)i��=�U5F��(�2q���*�\���%��Kv�����Fл��{t
5N�F�f�_o=�Ȍ�ve�`�}vrH�<޴J�V6i���Z2ih&n�o��2�$���'�	��)6��n�l�[(_-�6��[Ϫ}�%�dI��*"���5��� �%�)fx0��l*����_�&5�s� ��&��&3�����g�R?���0a3M��R�}����p���������;��'�%ߟ�*��q���4�?��?�X8J�!�{���O*\���~�J�W�)OOr����O�yL��G�^�*��7G��kmF`�r��o��� ��>�����k>A����K�n0X����3ɳ�fX��ZЇ����I�^xݝZ�t�ۉ��T�S��v�ċ#��դ7�޴�O4`�����4�	n	��9�s廍�\�EȦZ�x��
�ϕ��(o�ܐ�Gr��!~���J�V�7Jt3#p��H҇r}g��[�$Ryr��m��Z����k�L�ҤÎk~%��ae��R�>94��r�Owc���7	&]�I��n?�zc^"�I���U�v\��?b8�����d&g� �s�ъ�tmr|F뮾S3a%~$�{s��^1�i��Y��x�UO�'�;�G�=�a��D���g�6iN��׼P���Laed��;��;��
�I��p�5�c���R��|�)L�vf��_J2��f���hۛ.lt؞��)�m^v������v��Z���#f�����-o��R�V�͍2:?Ig��b:�o��u���+�=��D{L�>J�ijF�g�z�R��j�h[aedU����"c�|?}�,8��H�w]{��
�$nN�SP�L.�EP��M�E0n�Ci��v�U^Ϩć�F�w�l�nV�8	Ⱥ(���sd�n�|c�FB�1Z��q�x����yPVJ$�S��FnaQp:C�B�oF��Η`�sC����^������G��__��M1��:��k�C1��	�0��m���� ��b}�P%$��8(wc�B#����uPj��J����k�&��Oa��)t����������k[z?��E�7��Jo'mW����=k[�oD��j�u��j9�����d�	���q���'O��lj�n�o0��d/\b�h�@LC��9� S���s�FY3j��0�c�k��R�;��դ����	`�zCa�A�)�(Rp��k�6#����g�F��)��]EAtX~*����qVX�$Ւ������s��l[�\�VA�����*��9�|͛�,�-��j��3C�U��"�$�-[�%�*r�v_��*��m|w���ϡ�s��iF�����+�u%b�Z��c[�ip��g�դQ)(T�cl�������:�)ĪQ��*0���MY�ϊ9!���K�a�nx9|jk8Ib�:�8� �]}�[Ց�ܞA��%�
�??��^�t0�l����,���Ar�������k�7�c�OR�F�!wy���5f����my��H��W+D�eH�L�c�ʳ>(�ԩ��18��Ql��:q�ٱ5gr�TZ��j|4Wi�o��d-娭���|O��EK���~��a�;r52����e8xRp>X7ol�"��wy��(���m��-�Ѷ�����(6���Ъ<��g�) �7�e"ZM���>n�JY�Wύˉ�2���΁���`����9_�=x�e�*�&��ꀿ>��L�i}K���8����n���t�gL�q{)�m���Hx�Ã?���7����aF"}�pc׋�=�46J�3-��^���:�Z�T�hΡj%hI,\����C2�|dgem_��g/�U�Ұ�+n�1%I_�*MO�w��~��F}��|�7�~���(�g!�#1��[����R�#�֚\6>U��e� �ˉOjP1n��+vZ��D��@
_�0,�;�8.NeU���N����6`�\�2Q�ԁ4p�c|�2�bX�lҭ!F��	����>*ô�1-R;W��	|��?U��:oc����NZ���C|q�R	W�\�#%� -�����u	��Ÿ���{�����?G{sq�V�N��8�EF;oω�V�<6R�Z�7���ܹ]���c�	�+���SiC�vf�3��K@/H�����o�,.W�e��8!a�UV�.E����X[ң��G�Mw4�*<�(���0�|:t�������$��|QWj0ƕ�u6MD��b���f%JN��3YVI�Ed^�^�-^0��3�s���yY�O3�}a�?�؈�D�J�*�F���=�h�t ���nY����N�$~[;ܐ�0��1�����p���8�qE'n{n��Z~ F�h��;]��;��o�F��ת��o�A���R�)T���]
a�+f9W�B��H��K\�K�!��'�i)lw�Ux�*_��J�{s��0��H
�Lkn}��`t�]�t\I�d�:H�>!�B��ȼ��i,62�t	2��2S���-x֗��=?4����ڻf:�/�i�t�}Qio�Y�ᯙ���vlު~��ߌt��b���CX�e���qd���L���a�~�J�r�'Wſ�ǖS��WX����OFjQ?��4a�.�µT��Awp����\(�V���Դ�E'�1;A��
��z؆��T��dy^H��,�" ���T��Ǒ+�D������s;Itl	.�	�z ��.x�A<;��wsaz �s�R��?��b�o��������H,~3R���������hd�<7��}g��K��{�@�=\���o���f�zÕ��W�/�ϺU�a9��w[������ J_2��E�?��J�$^���?�d�ټU���K1
��1���P�b1br?8�γ(��3r.KJ����Z
 hS�MM������$=�5�I�A����E��!�
I�^��ŭO��8I�`͈���)s/��t��
C,!���"�e}���[���:Py?�}��[�V0�#EbZ�F$;h�A�S6� rUq��C�����7k�+�n������>���%�e㇭�"�282�.%b�����+�l��+��8;��t���e8��N���6(��E�c�[���Į��٩���Wq�8?�K*2��3̝��k�z���8�KA��^[�mIz:������͉ڢQ�"}P�|�<Su�v\�N]����yp��N[f�S��|1� ��"6�cL�ځ����#�-Xqؐnt}���s_���XS,�`X�<V����|�E8墉��?�#X��1�"�Hd�3"�e���E; �I��g�<jӎ���ʀ\"�
�9)"��#���F���d�K��,���K�p��2���"�1�V��ԒG�oԏۉ."OY���j���K}�9�Yش�!c{�q�i���¿�S�R�Z��/���s8��^iނ�J�.Nry��8
�g�������dP`=�HZ*�s��)bף+z�(��wA-�����v��c�J�ST7мe����o���B�Fy��E�D�o'�|O�T���,)Rk�4�NS����!�S��������4J�O��@p2g�pk�ݸ&Թ+�K}�	���遙��r�ai���{ڠ��װ|;��yu��L��g�!Y����py�������X�$����m�T(�(���������s�+�c�y��G�����y9r��+!4�r�*|b��.�̧3�����с!z��d*���TM_+c���(Vɂ�٥��Ĕۥ�ŀJ��l�6��'<:���!���aq,O��N˫��e&_rcH��O�(t����tdv�6�Eñ�-��ݐx�B�����=$ބ�|�_��]���[����Q=`�ۊ�̎� �Pg4�-9�HU���zG��ދ��4>T�?�� ��0����ڪ#�2^E�p����5�OPYhB/�/N3^�0�yU��y��"�g.�:��)��C�ϒ˰�lP�(1��t���o8?�]�w:Z@0�6���-ܸ�8��ntۓ��Z�q@��&�f/q��0ރ�B�7/3`��]�"��8�w��a��Jod�J���)z�V�]M��+gl9�L��]��wj��Qg��2�uQ�ɐ}ȧ�4v^(�!���*ڡC�}]0�Ax�&�)�Hh7zh����@p��9���Y��7��'%DV��Rsox����B�U�Lg4{�4vD��1Qۤթ�4��H�/�T���`�,r�'�;����|J	�2�#�֍՜��W	?�����4� �ħ���4��9^| QG��O�����qG`���=K�y!�gD��V��ƾ���ÒĐG�$z�����P�Z�:�T���+w�P�]�Iz���BD#��8�2<} U��+�/r@�/N	�Lo�V�T�$�Ty�P?%�=K��щ�B��6!u��$�N��۞�!��K�XsFp�C�"R�@�s��9><�V���t�c�u�5�cEc�w��#��dx�X@j`
�)�m+�"A����
��꼧������Q3f?�5��v�� �0 :	,+H�m��:�`���4�C�cJV���$2��Op\(�{��8�5�ۦU�?��pU\������ɸ&�6����H^���@��~��S�=;TKSkL�6ʼ?5E��+^�@8H��+�s�C=��4I˼\Pr��Y*c��>�D���Qa^��^v~Q7@~1�����VS���[��\p�;K��?�J�8TD�E�P���v���\V��s?9��d�������k~D�fôE�Cn��'s�k.��"P��aDk�PJsQ@h鵩��2<6�Zм!&*|�ۏ��;�}>�↴D=����H���u�C�lM�I���W�C~\\4jQ@������m`%3	��[��c�R�n��� �z����#+��yOe��ߦ�+_�Y~S�b��Eh�����*N��l�$�LI��l��^8��=�K��..��Uy<��8�玓,�F|�`��ELؓ��%�"�X�i΄�Ze���G�9�\*�C^�i�P����p^�;���q��M��e���`�kaS��1=r���('P���$�����b9���=�9��WIΜ857�tx��1ҋO�ջ��B�6�tw�g�G���%HT
A-��M:��չ�0G����d�z���+�Tq���.�$��(q"���7�{y:�1�g@�� �F���素���^���ED-��ƣ�+���v)� N/%�-6�oh9�ySY�)���$9"�g���՚3:�k�M/��1���j?�q��ν�7�{���Iq,��K�&,D�%q&!��F��e;r4�\�绗��gמ���H���	�'�}���6�������-6�&�������D*���O���I����X�#uj=��c�-e�Ǻ�CDщt�d��p)���ė;T�h�h�5#�M �����<.����v1p�+�l�
��������>u�D�(!�zR�3�-͹�ٴ���p�m7:����
0��O%�g2E>NC�����P��T,����ڢ�)�@Oo��]�~]���P���D㓎�����_5!���F���@�K����9.�f��7?�q�G��h��ҨFw����ٌLA�#p�o���ۖ8d$B}� ��$�M=� �2�:R"�b��ȚC���J���6"�V/b����ؕ�8����|*�)�.��O3XQ�~�E�K���hu[���bP*K+Q����M����9ؘ�(�26�M��XÑ6�DZ.��XxV����O��57z\A�BC�yQ�dx9�x�i����K�F��ټ��P�,L�\�A�b�C�X�s��Z^ADн�zP�z�����U�`yd���J������F����_���+�es��;r���Ҟ�x���h�E��(�~PO��:��n^Y2�\����;�^�,�E7�!���:���~���|�����v�ɇ��.���������W�k��.h�	
]hr�&	��C�����_t��������y����Z��ʞ&&3�M�|¥�O�NM��+�.�s6y�}Kz���)���߭u'�a�̩�y�PUej���X�H���$�%��)ܷ�C4�rd�v�%d���C��Uշ�,�o0Dc��ir�8%JZH��u?޳}<F�䂣�+�������7�lKk饣8=/����k/P,n�%�o��n���}�0�U�y�W��z�����_����?��ICTE?��$H�%���l�Eu�SF(c�������:Yh_�,��⟍Y�]f,��+v_�B�e�a�n����<�(��+�1:DtnI��ৌ�:��2��FT��R}������v��j����c$�u�P��d���L�ɘ�W�ϡDĀ�9��w��*�*>���������T�I��}�'|��m�	y|��Z�%ml�ѧ�