`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
r62cbS+9jhzz01UhsAASpDYyBYMvCy50K6RrcHfufoMBO3eSP31+FqAVtPCneonCYou0Mgu1wGgW
Lr/P9jaXu4jUYMQ5mo1h+X3+RBsg22+4TtwqNYq4u69FmD5Vf8O+X1Xdytlr/LYhMK54CaFbgoGB
kvWVj8F0WxUgBtFa8k9/CKxy4v2juHsYFMJM6Fuopte6qGOiE8ysrr45hgD/Z+qLF5/yoDBIsyrt
ZScGgXgRoRRXjcGA3d2S646A6/zOimzUs8QR6n9VtJ1JCvQcnqiltvwhf4Y6NySnIkJHU1xcf/Us
m7XVhhToHnJVXzv+hPxrZtzNi8nQl5mQSINTiA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="e1aZsPcYLFJkAO6L5uAAMBR+XuacM2up66BTm+709JU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3056)
`protect data_block
YzWwUa0z7RiqBjatQExye5qHEELJ1685pYDMGwR75QjGiAQaV46DhInEvBJHQY6PCkA5jX6WmDAP
OwEUms0LaBgMk52PNJNa0t0PNIJwVq1FIirFsVY6EE8LPkiubp2gOQp+t+ViPfPD/RGgE3NF4OhD
FbB76/7wzAmDmtYsPGp1q/sKkiStPqRe5oZsAgw3o+yyBXURBJVX4iRImi7LFPz2QLOiRY7rAORB
jLkfSi5PcOHkzymQ0e7MA4DtebOF9VhE2/ZR+rIOj8yWbYkwhy2asDfvabMAqDljN4N5aHgWBKYW
j2S+mnZuPqd5CZCamcOoO09ZhVhPjmr9YksX2mxZibbV5XJzh5qpacBPKscIrBoSql2FTOX5bFYF
SRjAwxF9/ikJTkKXGAIPiTV5eZ3OEWanI2abzhKY85Wtk1irLpCp/yTBPx8F41xqJ9AmkKigP+K8
ZI033sMs910Nfrw2QilwryIPkpM77EoYpzl4mhZBa4b88QD05RWa7z2ApvzZRwqj7Xyg063r9D+s
6nJK6UuZIZX/ypALzQkjMvRsfmmppPTJ2QqcYxsMq3yKxeQP2tTTR1+Mtvu1GfsWHC3D+GG1xLni
IWFGn9gnVVv86VBFGN74Uxi8C5OR/G3U6gCeSl+Q+hCPOVA/y3o9rX6mRi+9Lh9oFIaxyton24OB
4HO4K1Zc3Hx5LqQGXwsCSjb7rv0dliWZiubqa569mWGrjPMDHevVXF5iWd3TBN8TjJoyWMQiWJNX
R+elQWMkufTb9sgvFiY/yjsVh0paeX0vV386qqIeuKivXnTC4R5RBTsqW2YZTo5qBL/4nhQCDrFz
16ZHE9pLWNF/WbTrALeKo32GlTtAr5FXBXfHxZps+4LdUGn2Ryc3vP7kR58QZM90u7J1dlULtvSa
zylAX2N/eSz3QQs1/n1xjEdeoJThCRQ6+Gj4ogBEVppm1vPq4e2ggI0lrLPj/fG0S+pXxeASxBPm
i0xG2awWjLM/xcLuYZTr3+1LqRQINgMbdwp2taq29IvSkbbBLIxc4felMuG51W3EHAnr2m+9u9uT
Brs/qpBVGiZf3+ZGPEUDl7CU5bGGsUyntiy/ICuQGB2dETeAPMO+z5dS4FUWSSb5s0rbOrmIYrlV
uJIw3sThYToJDfW569fcxNLTn2UsPUciVBu3g3MnadCeLwKqW4NSzNhu8g7V+XiY3zqU4bYhCftA
HLNqZ1aOiNyd08RbPTt+yHak56UEsaaLwgowNqgZ2hu0oK4vvnv+VK4abx0TAVL8HOd4oczpggTv
9h9thQv99dC+LyGA8kuOFcYuP4Ud+ULNb/Rl0XH2Fb4/ya67GXDWTbbVNWQz68jfZIrK0Y5OVfIM
IDrbOYAb3oam/+ckh7z6jPC5SekRJIWxfw2o1vv5N9669X6w+6raWrRoXJN/355MD82DRxSu6Xyh
Fw7zkOUTxLxpCZuclhsg3NodmnesG7Tac2Lml8CxKGT69arxdFwFDCGZA/R4nyDi4nderXuH1I85
xKEUYnx/iUGiyrOoXW4kuKUML/TtH9i7AKXrK+Wn+427itJQqa16PyzfoCKeHErO33F+D4YNhGcw
2lWbBNus7WqTX0+f2GmDv9Sb1dBNS9WfOhYko/o8uDP1ug+foRl8PQYyA6geILfch6ifFd3wtZ49
MPL7KHEBtHEJiIVn7bw4UFbXkVnPAs5RekLjur7dclza7QHSJOOdjxcdnyl+fxs3VFYd3FQ66131
4Q4OXD+UToEQErZh+33bme9rYI2sN+YrXDYQOskolVsqvl7I2aYi++KYIkuB4Wh44u2lRc8zP2uP
wTXPYw7x50IIYEtzT+oPLiOyX+UN1qCIMwusdL3FqHYQgcJqyzSrUdGGAhrqYd3Y/ZsbzROTMEWx
26o3/qTgcQ7BJbu9XrRJEvG75MoTccfscDQvd/C8nBvVsEwjbSY/JQAstC6EScOF9qG0k8BQqsAP
99UHfSWMK0nM7O7wbWl8jOvUPHvxMynTWbRfSLya/rLgjH25TXjR8SZdAbjdGOqBY/QCwwb3bkGy
lo9cf4C5vd7aOc8eEvUdltlKdZ9+xQYVtoUD0Wte+oKwBI65jmMpru1abarywa1IQMsU5+lwKLQm
lH7kiblZvKJgHNn5rMUJ1A1VmnS9wXhOUEqMN4t+D7T+J64PCP4yuasUSLvUEEy9xaBytddmdy8c
SV8WzSvPG8CerALtZ2dT2ZIjnriaIO9ULTdlcdWv+hJ68cgtA2DZK2f/Lk3xadrbU0uXgTBXL5FL
u9M5vXv9ypOW9R47kH1moyrnp+CNeMm03zXq9FGP8CktOw+qpsAfVZAkNuKPxAePP4ev2yvHq9yc
qaB4uIzko/ORvGP0H+yUc8hWEf30+1vKi8ofNB2RLmbMvsNeKXczNOn3lExgbHsbBHn1wvB7Px7+
QvN+w1fGFLxJ3ZA/vI57dhEWmSo6aWzjGZT/XGt3CgRQgWl27wEMVKmry2iw2cE7Oizehh7Ze2Oc
TKvagt9/LcCoiXbaZLj9v4Od3JwMDPxsg29qla9TGUVUzdX3yVWM1Q7Ex17e9YCYFxtK2CksAXgV
1ab/haHVvQh5+b28QzCC11MOI3OCpWti9YgYDV56jfeiST8rvezmhU2w6MQ0oWWZwf54K3U/dbwp
gJd9rvLtM2u/zlW0lUTvG75DfPVH5WH+qXYAGjE15ge0ZfpsUF3ANhRWRwpqswC+WDRYZ1G5jNtr
13WRAMVtDm7nmHSLTd4ra1DEhjY9ZlZyfA3rregb/EufcAP16mPjQuxgBDzNqYHTb8iDshEWMjb6
gfPe68nvbQ7TTnLisdVvmGlNOcbiDpo2tglE5pXxiJEUkCAmwmK/yV47/S/C8G/lC0UOw1wTndqm
HASzqlnwmjQ3PHm21gjbX1xdm2RvSA0cR62ckWDaimWIQn5u0ZuUiEWPBgncMe5sXOhMKPOGIzwA
CEnlxmIiTq26cT2rutSFxSibd+jw9ZIz73G9Q7Q643nySrl9q6o3igPYY8qSvz4VBitwCPzEGvrn
jPrsBg2Ypg3+CGAVQEHMy168XdQ0hD0YasAPqGchHu1Q/xGJnao8N3JFUIFfP/W+eQljfTwGtSyz
zBpZpIFMi0eS2OKtt9KRFn32CnRsiFSlRB1FJ0nt/ZQAUo8dAl56iLzPdYBYFaKy7I05QyDtok+P
3Xr+TevA++9SgRJNWTjddn0FnNxWpjWTB8qc8LHr/NoP3MYWbveHjOia2D4jepE6CqNc844Zzc3a
uZd9SPPQ+xl2Ulb7EpfekJnApWmaULPvNUybP6TIfzSvcq+VcVNMa7Ol4mOlveHEQAB7CtpwvAy5
A9SWjKOHbC5oVVXDlOL6E/1mBVix82M38O06Z0m+16q+4IRLxSkJVqLaSBg0bpTdPeKKoA3iySdU
0qp8pvvQSc2EIZL+WH+8Q16r8cAqBBiI5pWZhFZUlKascSf1ra5gENdd2+yDhadMz0WEf8iaGbk2
OrSXfqr3Lo4YeWDKZY2tYKmPWVzRIMWPdS7PF/FmyUES3U0PtGFaVeI/nVI/ZQFMLjN7dBUrJ8ie
g6Z/1LI/cd2nxuHs84ybs3ymAKCc5HmBQ51pK/91Xr3ivZUmlB+BZmPPHZeTNXOsvllXQGwLrqkT
kGPKa4jVPmzfi90n6gtXLRt2UdzfejDrvulMziuB4rKpIXlfF3KetvYgyCHDOk/HwBpwcwjDC1Y3
Uvudukkxmnv2QJ1e2aK7W8NBw2qrCfp8+pWOx6mnJ+7U/qoJrNL7zhDYYmAjl1oenf8wJBTmk+mL
xYg6L1Agc8xuc/IjoQE20tWCMB6aulaJ+/YuwToXfc6ptR4/syVTMr6UfKjrZxhvM11Liwk7fvOA
zZuxMprPQBmKHeigfzLc6sy7oI//WQkd381I3WYsqtmT68LDU33Nar503yYWt/hxRLF06M14/acN
Y2KgQefmObZB5uUdStXXYwLlgSBomkdWeER/Y24sxBfwaSHertXEsHqs//EClsG8+cvhVNCjnJqY
7olHeeQuEmk0+CXIog7Ju/QbiP11DBiKfpg/5F2cr2SJuH8=
`protect end_protected
