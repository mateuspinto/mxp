��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���� vU���%�]����d�S�}�� ����#*����tC!�?�}�L!���RB N��(���M�}6�Q��� �Bڨ�V���B+����r�����6��D��?Uf�3���R=����&�*�y� t����xw���|�kk{��ԭ׷�,Z�1�����D,*��%�cϋ!�r�N��TG梉��̿�ڬ�>g�@�]㴜�:M���}��,Ag��R7���w l0�*�\Ot��|md{?�m>i��7
�:T��¬�z���Aj?�`o�	P�F��'!h� �QGB&�w+L�y�R*�3��޶	�mg|�;�,᳆���b��Tq�j,�_�1�`��6�c�o�u&\�AUur�]מIg1�Ϳ�w6
�XM�Tw����j�7�a�j;���>(���4Z�]�񤠧:�t��G�^v�}O3= t�sVC� �b<w�b��W�\E�k7;��7���@	m>;���_3��P`)S�٤�P>R�Rn�qd$ؽ�]�*)�#t9���ğ�,�A��^�TA�lg�{�GtZ����������ɖY��>�o��3��$)��Y�A�f��2�_���:L�[���I��iD�f�~�8zΫ�O\L���G]�b��u
	y�'Զ�A��!�J�]���H�����R���ëѧ97zg܎�K�\����VE*7~�}�����)s[��Ա��X��1.n�[A��=��7�w7n�[FηOۖ�pFJD	�rr����Et����JRS�SG[Yz��d�Jo�}��C�&2"%�V�=k1��>[��^~2���k�ulo��\�X��š��~xr���@��F�l�6����RA���t*���n��a�Sk����W嶷����XKe�K�Qv7�箽'�f܌�.� S=����&�꒼v�D��a��ܛ`�Zowq#kD)�7����:_����ΎW�.;U �d�S��sk%�cR��\�:oA�Ɂ�Ĉ�J.&����*b� ��s��p�3�p�y@X1}	��g��2>�	},�'%�7WɈ�OI�9$��Z)��b��jc,�#{�Ȝ��t~�����=#��z}���V�yP�Z5�#AHɓ�-�$�#료Q���~ԭ{���RY��U�ڼ�q�|�~2��ȳ3<�.��=~�n*�3�0v�?�������]ʇ�G���:̈́J2t�P��	�VE�r:}��_�N�O�
�d�� �o��R��=��1��� ;
�x(�<Z���S����U�&�ꕜ�/v,vӳ9��\v� =к����֋@ڴ�8bdW`䝢�>8�[y�D� �X|UBe��zG�p}��9̅65\.h)1R �u*�� �g��y��IԕW}�q�
t�*L�c¡ߘSd���܍�N�!⟏�<��	��Z�2����྅�3{�X0NO�Mv�V���5�1Ћx�"�;��}I����A�F�RT�Q�4Xs�ek��u�}��޳�û��N
��e�?��@�D����ר�;6��p��2ظ��	�|�I.�Q0���c����<��YB��>a�	�w��+ts������g��d"J�R��$�jH7�f�>.��Mo���7e�ej��6�W
Ƒ� xL$>$
,�u�6�3%ub%�����-�k�P���,xɨ�3�b�J�~���+�E_C����&�^yW�=ȸ��m�d�H^��e��n���|�#��J��m�Ml�A���U�(�Q{9�?b�'�h���H(���	���t�ϲfZW[��deK���Q��=kz&�@�C�$���%*-��L���`�ם�}�i]h��oi���@�?�L��"l��*��	1T?W���a@-i�[[���Xo�2+�-��AHb��|�YKB��x�[q����(xz�̦rR#��@�f�p��I�5�Z�X5b�P���Κ�$��qt���u�!��{��ͣ�ij"ʌ���J?�e5{�Zz�+���2�Аc�Q�nz��f{wI)��f�k��N�R�}L�6�1I���{��e �{㡘e[Լ�|���s��}G٩�,������<�@pq����_����a�!x=XuɆ#2C8a�&���>S�#�~�˾��/������9���7��F2��E�L��;(-+{��@	t���+f��:���K�$m�f����i N1S�|�r^nF�P=�K2������c+�W	K�ᖊ�e>�u�?����N��߂�;G�hx����hMɺ�����;wK�'���n�. �{ɯd7ŏO�u���r�W�9���I�3� 3i.�8��nrJ�x��AQ���������0Mpa{�kȌ��^׫r�8�b��u���+�-j{����-C ���Id}�.���~c�EjD�n�h��W9%�[��Gɍ�F=X�t�����?��aS�����a�:���י���������F��T~�%�p�da�b�����;�x��;���cxu�О�=䱉��7�T�$s�UfD��4cl�|�7���/�k�4�� f�в�ƕD�{5D��z
U���n�	h"�<%�̅�֕������6_��2�\_S5��1DF���3"}Ok�G���@�m�����
��(�+Ķ`Tl?Pa+b?JI����HH�%�R|��#����:�7��N��<�)F{8U��b_��<�H�u�M�\��!dl��ߕ���]��-|IQׯ����Tt#&�:lAP!��j딚�����YFZ6`a�؂�U)>-ˊ�5v^�F%�7�Q��2�ڌ���E��s2���=|,{r��]�� b�$��� D�\F�x� \���6ԫ,-$�[�}W�?ȶ%a|Q!�$ �_Z%�F�D�,��z����}0�5�c_�� ʒ�RH�
��5�0q���v?�al�Ź:T�z�#:�$�|Y)G����xڒ9�o���������y��t"A#.�ys��ԇ�;9\8��@���~up�#f�ÿm���C�@9�d�kG͞nQ��w���b�|X�a��.W��?<P��װt�>q��OQq�E7�|�5�����γ���(�>�W�t�.�j��U���_����J��u.шƱ�4�tgñ����R���'l�J��a`���gt��f�d�������l����pB�-5{���?D2�Ĕ���w�&ܗ���AYG������!	�I���\o�q�fµ�G�-4�9-�<].L@�ɢ+RղCM���y��4��l�k!�e���Ɩ���BǷ�e;��ǖ8@���M�P/��xedW�oO� /��_r�}Y0���8��:�á�����]�Y��*`�+ӟ��'�غ��S�� �Y����j5���V��?aG%)*1�
~ԗ?Q'�[�+����1WJ�Ҳ����K���O��x�^36�\~�̛����s�������.�!or�� ��nW�u��`(/�,��Zi���� ظT�NB�ǁ�����^�����@�F6�;�5�z�(�����.7�[��O~�c�R�(t�5;ݻ��U1:��(�Zy��ѰI��s���^��؃覕�)p|�Mw��ˉ��ħ����
�{Gr3��~��!I��o�qk�Ez�r�V��i8�ݸ���DWߺ!�*� ��P�d�G���b�� 6^:��F��!+0�qt�����_�>2�?�����\Aj�*�S��;}���;W�0��B ��cV�;����Y������c��w5:pa�f��<M�Ν̎e�˹��j��;S䧄��LD���E0)D?��-VuY��>Ɔ����SF�nhA�r�4��`ȳ�0)�cz�^�To�=A��&���KT	��~�uR4@LJ�����#����k���'<	��7������^Q(`�ܭl�1m��=��v�c ���i3iP�faxh�_o_��y]hն��:4)����׳d�&>?��$]����[s:� f��SSo�x�N���S.Z̾���^�nQ��o��(\�))׍&GM����P��M�q�%m�DT^V�P��=8D��rk]yצ1��wƤ�5la1��?�3te���'���r,U8pu����H��H���1MЭ�"�;,Y��c��f�o3�٬2
K��:���Qѹ{��&X���rmQ������`���@1�f��?xu��po~�Ybz��7c�,�a�_þKdD�[]�:`g�jqE��Щ�!�tz��QP-��#�j��4 ��������T�΀�9��ovDS0���B��>�B 1�b�Ua�]wo�CeD_d�m=����*��������ujH�����|=�_�S�Ӧ�x^������b���s����.���N��X���qB��K�H�9�L�J�p]��\��&���gAW��袄�%���oL���^�BB�pl=Z6S����*y�X�[2����}��N�I�E՜�y���b`q�W�П��&��_0�I��i�ʳJ�W���X��q��� &{�B�L���A˅$���'�i�dB&��[]x9��b@�����Ԕ�
�j������pQÚ�(��ف���?����t18|�8���s�νЏ�x&6�"���)�Y�	SM��a	a�]�9����ߜ[��WQcU�� �B���vO����bN��ّ����o���s���D�O�zk�6�|&V���'C�ŉ�nP�� ���qGi�3�;6��0>\"��庛d�
.^�S�m,����=Q�`%4�'�qtɺ�?G�!�= ����P=bƫ�`�"LHEGw�4��:pdK��m	K<N_Ù|�H�+��:]3aU��%�W�n{!c��Se4�~i	_�r��	�p��e�;s��ɷ���h��R�L��m��+Ep9hn�C<&ɛ��OT��P[�Z/�+�B��@ʈu�#|�M�<rv"���� �u~�\Z�B�d��g~:�e����w�� �[j�����-���O��y�>Z2�g��
�r�n=���Zc]���d��Ř�����)��N�-{U�v7��ƉE"�d����lHW��Z��a;�c7�����6t1�<��Z��od>g�'-o'9�0���8b�l\���>�_I#;�Xބ�X�<8�"{����-��a���i�R�Y�7�`Ҙ��]��S24�yX�|n7��=�WR/��eE1z5}[%��QN@��@(7^N�*A����˳C��;�����*��������Aܑ�♅���K��>����d�� �[�[��z_�3{lt�Z��Z���[]��Z�դ X��Ӫ�\�E;k���ܨ�en��q!x�,/��4)wyH4<V(^C\��s��#�&g���pw%kZ�c�d��2p��	z�4*Zn�o�E�	Z�@WA9T��o���rк�Z�C=9D�Ê�#������������3_� �т����� �kYR(�<�]٬+���MB>@�
˰����/�>q��*B5Ab����_d7_�n�.��r@JE�ϲ�T,��/)�����%���:��W\�7g��E��*F�>>�_�.4b0�y �s΅�od-^%�o�ФQf��<�V ��z��5�u
�%�ј*��2μ�<w}р��m�\����9W0Ŵ�Ko��y��v�q��h��}��	�FC����/�b�9�|�6�x���Bt�]�V����J`��h���}�c�y�c,�=�.�G~�$��m�M+��P�y��8�������b&�)p�GL���I1����y�G�Y����H�v���P�`\DBw��o��%�H�"1B�
�ߝ[k2v)��ۅ�_$��$a���)��[Ћҕ��9�҆�p�q���O����g�?+;�,�;��IG��'���0	�أ.��# R��$r�e}w�\0��p�������?U��H�:��o��nT�7�Ȗ1����u,<�������.�܊	FR��t��.�����8 �̀��8�۴��_�(�����@sͼ��_�jB�#E����BS�y�ЄL*0f��k$���;,���6qd �(*��m=B�oN�B�B�!���|Z"A�J���w���ƨbʍ��J�t$	�{������.�����d��[K	��V���1_�K�𖤽�(�]���-�] ,;�Ӧ�@��p'��ވ� Ш�5��-�ˑP�>\�< x���<�܁U�J��8=����ǸW[<���t�X�zsoٝ�YG�A"�atxS�D�}��@�����
�i��g$/{?D�`��E��n�8(���Z��S��(�@��͟T�ϋr�|z�[P�Z�FQ7��x���T���.t%��G��RŹ$�y3+_���d��{�x`h�	�V*�������\�:���J�:I}�p"�:����ڝ�����"h��+���	$>$
��������$�D��u呾�?3.�l���'&�v�l=o0�3�B��`��ʯS3v�N��
y�n9��a]X����\�g��ݳ��#�:���)!EOPV�\%}6ݯ 3���ri�W;S%��l�	�}k/�{Z��gx��s֌c�d��H^kr�B�`{#�����DԎ%8a��;�ܑ�TbQy�[�b7��iU���g~$qu�@/��Ĵ�t��Z�����Z�H;��]	�=S{����B�����k�"
�ԥ�e�]c�hbm{ktm�K@ɝy,�	�-lz���݋t	.�e<"�� d{��R�dR
t)����r�j3ҏ�ޠ�� 1[=�(F�p�;y�C�_dч����'�L�#Z_�]TS�����)
FK�葯��3�B
����UV�R��9��Hc�8��SQ���N9�A}�S�!똩����{�l�tL��-����ۙ�g
�	7�91@5�t@Ř�ת�����H�@M��2I]"uG�O�����{T&�E�#�f'��Qq̥ $��.1���w��o�^a���#Lԭ�/�V�A�[Iᴪ�u����W!7N5K�k�}KVD����Omo�� ����љ�<�6S+sܻ��%3�ߑ��M���Iu�6�������T�j�2
����M�� ���l^*��GB�e���\�X��� <��[�3^���_'b��vh:��n�+�%<�I.h��5��I�-c�x<��B��Ӑ����zȸ&��M��Y��J�̮�$��L ͎:��خ������F�X���Pa��1}�����tz�����U��:�?9� 6��E�NԨ�� x��:��ҏg`6Ty��
ӭNn���p;��	�k�ω>c�3�F~��8�60I{��S�8�cw�վ���(�.��!l��E�'g:>;�LZL�K�`�JO��c/8���/ʊè�����	��HZ;���+*^���|�������y�)��}���_kC�ɊRv�5'H�K�34=�zY���8@�3ɫ�K��*Cӏe�?>�ቪ$�e�ڴ]��S��Q���

�P�cm�`���r	���x��TlW�Z�[��bT|V�?�B�>><hU m�"��%�L�ǤeW���� ������!���"ܓ. E2z"��]���z���#���G./�����_��9��;�T��W��o�Л~Hŗ,�A�ɹ"���$%��Q7��
�*I��ņ��<��Ͻ
Ƴ�FP�=kpx��g,W�{p�d�� k_%���
�Ȁ���ڈ���-Uç���g_�����o%6	\���Qo}L���U�!A�w��x�����ad(�Mm��D���h�g#�ob��V!�l�by"&��L��{#�{�A� 	�OБ/p�-F퐂�Sr��� ����TL�J��V��\I�p0:d��t��&C`ۍJ�D�PE�!��#�ðu�Z���9�ʌ+fN˛!��4�?]�G<Z��@�|��	�n{�Ar_�<���Q'�J��{��6���E�4���p��۰��n��We����=���b�45�%X��	��^
w^��KlƂ[$,wf3�&y�H�wF�����b�H�7w�%�Y?�F��E=;}�zN�3�gv���\��8��n��J�B�D�s,�H�y���vqŅ��U������u�[�g�����H����M��5=i7�^(2����aqȌk���D�9-nsMQ�p��~�m�e�>���lІ����I�׼��rခt����r_�`�Z1��P�[Ҟ#�2J�8+�:%v��h�ɀ��NA�E��e�Ԩ��Zʍ��o��K��@�ŏ�J��yVώd@�?y����M�t��A����~�
��jl�|����g�Ϙ7���(Ku����T*<Mx#��>���6�:�;G�$�9���҉����C9%��$�>��)-��8PrV��/v�udA������#dX)q��<�q|P+���+���
c���tY=�G]���62h��B��Ǩo��6T��a��/��"v�\���tR����J��`h�g�~��5܇�w&X,?��!p9a�X�Hg�O�M�����E /���N���lņT:V� 0s#͆��R	h7.��t"Q *��s$r>n�BN�,��`���Tz� ,;r��u+�����=�)u$������9��BJ�i�J�N|U푶��I` �oo�E��jZ�<����H�T�wF�_�@Ԃ\�J?�3��H����'ڃ�O��X�R�DJ�nGs�i]pd���Y�/�٬]P��L �HL��7�v�|u �΂�U�T�ď�p��T��+[G�m�C�>��Ѳ�cN��ry�_ǰ�e3Z����6�ƈ�;~ �^�I|�T)C��%��W�W"� �<���E�2�:��D��@���Yl3���r�̲��^���Ƌ��R+.0�
f�C'T�$LC
��6�oyp�w�Bj��A�-�?L9A���P����-yOS�óf!`�\����$@=V�V�G鷞s������--��F��%o7�n�d��e(E!Xɖ������VLQ�Ne�$|m�C�}�%��_��bA����8�Ӂ8��:���c��Q����C%���iyb���i�̵����Ͱ��m���.︠WD`.
�%i��e�o��V$�1��4|��}`�gP�s� �����(q|V�ׄ�h�Oup�AQ��Xln�9����@���ý�/Ÿ5ަZpwMkTJ�x�S!8mk�r.�s}�кd�O�^��D�[5�L��N�I�k�0}�'F��0/�] �����z�PW �2(�R���-�G4i�ZJf��&�+��:�,�0���kBdv���
�PN�9\�Q��V+���n�@{�nn����oc|�}���T��Ǘ��rnz��w�3P�OR��	��W9H�V�s�>���~k�ukk����M�pX�h:ۦ�kf�a�i꓀P���ף�ɋ���Z�>����:#y�7�=t�捏K�]z	D*|�RF��]��ZW�s]�ݝn��oДw\�O⯥g�X��`}S���n����f��jQ�@��N��	"p*�&��&n��] Ϙ��^��£���@
-9v�_G�*J�n��jV�%�W�b�[1�>�cB?���u2���)R3�7��"t��~g�����zD�hM]@���صĤsK� ���3�\��ʀ\��-�G> ���7->oš�ohs�Ƞ�;��]h�j�$��KQ��JC|��[J��WI�ΐ
����n�S�kR��8��GX��?�g���!�;[3�*��QC��{Xl�4���'z_Ģ���*�R�t��%��4�=Dx����<RQ	E���2��f8,]�m�e+u��
��C]��-]I:��鬽lK+2#�N������p�@j 7YW-mD�j�Q8w�y�fR�ya�j�:�b���E�$��/�68�v�,�L:"6\yp�<�ԶNa>��L��!?@�bpS4o��OLl�`fZh@|�g��m�u�/D�6�S�Gj| ca甅������E��x��i�wU!ъ@� w�����6����-�o
��]Ҁ�P�+��1���,�	�莥@�/��a/:��)-wS�.�Z^}�|-�m�_B�3,�Z7�����31Uv�|5+-a87�8����(��,���4��QB��i�<�=���������(����Po\϶��-���D±e?�$�j���9���i� !*�-\pm���Zڭ�^�|�
ڟ���|\�%�J�W��m�XϿ��w����y㑳���z
Ft���4���Y�H����U3ȸ�]�������~��p����>k�^Ez��<�#���K�ts���UD�l�ӕ�R�昹�){�$kx���h\Q��(�������ӏʠb�Mj\��(��i<�W����ۦvӑ��c��Ԍ�"�a-���ZP5Y�޳�+[�p��K{Q����������At:��âO���KB>�i"�����FG��_�A=s�vN�%:w�2��")�����ݑB�����ryùdw��^2�_���`�����|��3�\p��D��U��r}��h̟��WG���x�G�_�9h�����v���n�9�-d� �(E�h�¦M�T�_QX[�]xyA�ȸK����"����e$�?�UpB�l聹"��tmk �.��\�A���]q)0y���KpP�H�Աq�(t,�fމ߽�v�j���8NEm�^� 
j�yX���
��kb�YN(�ڲ/�#UR���PY�4���5qVt_��'����q�I�Y����ߴ��j<�e i�aю�CQ@�����f�^����9�K�Vg�AH��f�˩8bh"f���󩏌/�2��{�^��0?A*ʣ��t����3�B{�=�����2lx�,	�o�ʂo�>�`�f�NƓ�6�3D�30��ۜ3�g�\��II�+<����n11��e�l����H`�!ӗ�%�)�4A�~�H��Wx�CƳ��[��[\��Mjꇤ؛�2īP�4�T�x���V�^U��Q�e�E�ͪ�-O\���0����+\���_&K��m�e����!žA�= �8��7�-
��j�D��o�{�'��R�t������R]p�/Y���;�GH�{|Y�퉸%z��y�X^����7ߌu{��'!�䥻��z=W�R�|zY( ���_��0��p��nG�pS\vץ���� ��y:<p�9���ƒ���6����!����`"�;x�wV�㼅�;l5���z��wp?��Y��di�S��/$t[7���ӯ�����:-+qꁲ�u�^V-V���ݴJD�G���י\��u������a(��mlبInJ�kp�_ʸ�F
��;��nh�,������LF�^�~����e��X\��7jB�X�-�����4's�a�I��{D,Y緀_�\�.�O�y�4�*	>�߰�����6�;��B>k��G�3<R���⌑�����P�Dڱ���
|�5�k�8!^�!�M�3����2ö:V3:ջ����s%PR3����-��v'�ȇ�m�oNc�Q��]Jњn���Pb����*_f�;%�2�(ܜ��66%4J�uI*2x�O���I~�b�n��yt��MO��M�5Us0�Q��bU�]ER}���<L0�dV_Փ����Ǖ�2!N
�X�|nhpVC�r���~�k� _���ׇ�e1&5��@����F�O�eiƃ�c����W_U��a/6�\/�8>0[%L�p٨D���J�U�`�ֿD���}�ȶ[i���H=C��W94΍�
��� �f�?��{�O�R5�몄��Y|D�
��+�{d̈'^^���w�q��R2u��1������r����]5p���%o�����%!tI$�����~��n�_c�1��̔���!�d�,؇�n{N䌿��0�3Px�mӘ�C���K�ʼ|�$-=��K���A�J�^�����|[?a�⒊����*�ָ���id��K��1��~��M'y��!ɠ@��S#I��Μ����I$^Hg� �qO]�7����K�7L��&��� �<1�Op����'��՗��şr�ŭ��F�� ��e���{��`̤ŹpT^{�9!��	�p/�1���N�+��{?+P!��%r2вS"���
]G��?R�7%�u�3 �%�Rp���=��\:����e �U�Xt`���"��I@ҥ"coȃ>���g�6g�[�G�z���&��1��.�mg�gQ<_:�ƯX�dx�SK������e�B� z��Է�ˉe��ӹ2y�wJ�nM[+��s��&�or����W��L�F��A"�J�C*&���0d��EO7�B�m��;�	F�qK��_��-Mܜ|l�!�վ��!���d!rl^[�I�:%u	L�'�F*���U��φ�}C�tv�b6`��gȢc�RtϗG�<���51$�}��k*_����H��u��j���:����}:+��b�\򑊷_���R5�� �FҎ�C^zam|ҵ��K�ה�ѵ{�	*����4x����S+p�� �b��O�u����F�B�a��y��J�' ��-	�`C�Aۗ��%�r ���H]O��Qj��q�-,2�J(��HB.�;N5.�fS9hC��~۠t�]��?΍���Z�C:#jb�ΰ���������x��"t���	MS�<�m9�����K��nH���P��/�PV�@�脊��\�z������5��Bd��?�U-�~}��itF0�r=?2HȺ����ىm�fQ��d�T6�j�U�K�n	_4Z�H���݆�.��Cs�-�>���,�aL��z+n{����^!~���_\��V��d�~a�q����E·��se�!�J��p�	����;��o�����K#�>�J�&*�|E�>v4W$�����Pp�1P[p�_ֵ]�� (E����#Y�Yv�GO�6�l���Dz���U�F�K��6����ȅ���J�\�����ea9����;����<�;���2�*ß�7�W-ٹ�R���R��g�ч?��ΩrE��+<P]��,V�h�*���O��/3UL����<F�Սh40Z���^`���8q��?I��Tt*�e�E�k)�"8g)%�7��cD\��-Mͳ�F2�/�MO7�#��C9IB��l�����G�C�o�A��Ȁ)��H$�#����7<�*���l/\ih���w@#��n���E�uU4��S/�i�?��0���~�ib̀=�#Ʌ�ɸ�?���g`�֐c�MuD�?l~�� ���o�s�6}T���tiJ����md�M�ߡs
k��7�OJm�ɗ6�Rػte*>��.:��V��U��TC%���+n�t@���:$�9F7����v�����������VOQ������{�� JL�|�'��3X"�Ŧϛ�������Vi4l�q����������FR�RQ��pj~�l}�>=_?��j�|����q�Z6´!�^��Bߨ�{�HS��0QVB��C���+�a���I'�Ѷ�-��X��o��\}�X���)W5V����n��K��MeK.͑�K�IN���1U��IQw�b|�ƞa��29�.�����ᓷ�Ot���< �5a�U ���RU�(����5O��IE���t�N�z�:aI���'~+��q�AQ�]�!$��p��|�:��Z-�
���f.ͱ������]�����o�@F�o��# T�G�1v+��\,Y���M��H� @*��?��D���x)��R^L�u��ǋ�g���5��d+��C��bZ�˿��:�*�heO����d@�8ñ��ڱ��cFJ<	�G�ݔ�?�AV� �stG(�۝�Tu�#9u*��AU����1jG�0��Z�Kq���%LYB%���7�=�aj	�����l���	�:� �+nh�Y%��~|�d�*����	��
�01� �}�8���t[��ɲ2�ݻs���r���Y��&��/�V�c7�������-5:v ��&�j�]|w��
2u�79���=�5;fi&�U�JڼE�wl���*��ٜ~Qp6���~
|���z����I���<s;0�OP��L~�M��t�@�xP�H#�������S��o�@�\=sY��ִQ��]r1sx"$����6�3G�]W����L6�6��E�!�Ii5h�%��s�q������W�t�9�4jnde��	�
��#�A��B-e-N�����]2J�����/�U���J3��5��E���.[V���Տ��1oX ���#]"�!�<�!�~��-��ze
˗�3d�j�Hb�\�q�p�����r}t���H��.L>���D��^���ۂ���/Orb�tY"%�g�d�X菘�5��ܸ���ʶ�e�ȑ;`���H������q�������AU����u���&�V�	L m�8��nW���y���$:��L8�~'09k5�����OZ�Y;���ͯل	O�J��MΊ��w9Ǟ01G�V8��c-����='!~!��B=/�$p�e��I�W�8ی�7�����W����9$UGԍ�$���啭h��f���"	�v���N����8�ﶊנ3G���T1;*���,NR���\K�m��=ǣ�5�$o�Q��zzv��?��吜��$����P���~�?��\�_�Cgر�G;ܵ��֒V��+G�����F	o�����x}QP��䅢}�	�\��n֤t�������EI�Ba�GP���Q���|a&P^�6FK5�|��lp�!�3��<�xi�3=��J@9g�vnk��C��(6�L�~?��J�j���2��	��z��8V��Ϸ�EN��a1�l�;�bx��Nk�N��$�s	�.|�6�MWO��"�b�y�rR�{Y&CO��&^�45Q�{�ԓ�w����\��4'2�$��!�(B5��(bQ�=�a���+����N���q�Z�]\��$����}�u�p$MA���#!�](���"�^�ɾ0��.n����M@�B�I���Þ�}��y���.�Oל���t-mQ�i]�9���"ba�O��F�ЦNV��zy�+��^�fEl�h`M�JvH�3�7�o��E%�j���w�����VmԜ�}P�?N W��aA��t�²j�M�$Y�S�Hu!���G��g��Ľo\i�k����=ew����=�EzY�c<����7Q�m�a��"o���p��_��B�~��o�u�����%�r��*�������-�𮑫,lm��@4G�l*�0��j��U����{JZ��[\`z���4�=�뽸�>���&��` e�j���8�׊xk*2G�G�u�q��h�h.2���z�h:��Ly�_��z�V�J5��G�B��a��t�U]M+�4�Tؗ�ט%��o���w(�Q��H8�bo6��6R9X�<HRLi�g�u
��++w��K�r�bEl�=x�h��Z��F���U���bl�򟇄$ęvr���ݣ�Z6�P�i1�J��X�=�����[X^w#>�
�T�d���N�:x =OI�E?;5�䯬)zw4`Gz��^f��d�H�r��((�Ě9��}V-<�1��㟢�$z�a���e�oҀ��G��Q7�q���y�C�P�te�Yl�3!q�G0~���]�7:L����2����f�����B���m�5Y^���i6[���f��Jl�� ��y���� �$t]Z�r�!b�e��"{�z�ںD�!�E���9
�3���*���Q�Ft�stW�远9Y�S�I�Z��+���@_�_��R/O��
�:��#'��3��2��0�%�c P�#�넎���`����}���8U���h�a�YC��s��Z���\zh��[P� ')�d��c��}aZ��@��#7�&a;�%R���	��^�Y�db=�@�1<��5��`h�յiY��4a�9j�m#������1�1�@��b��siZ�1�R�_���T��N��/��f�XV���%�3�3���Ca��*�@�$u[z��( DE-�\~Lzgw���P;���٧��mq���D��e	�1��3��Nvj��N/yt�LE�E7S�p�jY���/B��K��<i��8�$�#��$��:Ν�2�3h�0����&;,���%
G~>����0Ζq}���L����>��(ۯ��T��/�>[�F�����<E����i�w>U )q�س�| <㜓���M���6�z,M�I�Ph��Yg����#�+���ͽ�z�>Jջ8	k�1�J�o7��G�J�	��:�h���hGʵy�=��	���
}G�*�K����@�W���"�˞��%	�U,��kv�&�'��U��c�p�����^d���⨌��;W�W��
��pk��{�� ���&�6
��*��?�%�M`v�@�"��@!�Q�	|� �/T�>FA�!���`��&���^��|�-s)�^}o��\v�#��x-���OXv`����M,��|��)��،��f+�R�tVX0|�
.1���Z��>FU�b�	�c8���y�4��V(�Uc�����e��،t��ӽk�h��&���lm���py#F��T��1�[���+��(!g�����"��g�̋��ZM�G~��.����#˒/��$�����¦K� L�A�.)�:���toLv��j��;Z%�����e��s��0׊�y'��|���Է����@O��]�������.���4U7�m���F( #��0�zY2}�Y�8������ ӆ���yu3�b��y�y�}�#�_�X�K���y_
��^p�,�&c%�a�み���f���a� �ٞ7F'S>FZ>� �{�ʗ�I���Um��c�Kh��W�������~\�����]~k�뢨�����G>5L�8�:����PM��Ird�@	%��kS0�+�9��_�OIv�jD�E��."J����9�٦�1R�ba�i��AȾ�TʩM�.�>�d�4F�m��oz��a�b��_�����)�2��՗�$@@�u���3�_�FRx{o��`娳�efp\�Qo1-��p{i ñH�)qkM_��]huEhj}��r�����V���f��z�2ҁ�&1teU���eݞ�Ԧ�O�E&'����c���~��ʦFܛ���2��&n��F6�z�����|��!����u�G̛������������㤆_꧲N�·.,�{g���r=v��mT$ٺ�K��p3�������f?�'}aNl���������g�����`����~�_���>�ƨ�������ȼ�S�)J%��(�u���i�4N��;�[m��yX5{iK�]v|�˸��ƬΘ��>�D�������IO-�P�E�?�0(�����3�3�(J��l`���E �[ǌ�7�7�צ���j��6o*��~Ϝ�B�j�n���=�tEaҁ�����زa�sus&�Is����M�C��Lk�Bm�a|@���(��ŰIך&�)�Q��f���Ht2 ��ޡ� �W�p�4^�+�M�5Y5�ݹh��������OV�z-����m ��9��V���i�h��2�Z��?Cǩ��
�?�5c�EQ��3ݰ�p^F�\4����&�8��`;���0������x�r2]���x%"�p@����B\.��es�C�00�R�oJ?;І���H.�e��m٣"�z�T+���b�[ǒ�J�{RxY��%[mŚ�	U�cm_��4��h_�>�G�&:@հu(�<���b�q�����ң�Y�u c�l��n��j7f�d��+�y�.,���mwB9d�5z-��B����;�hAl��ʦ��
��+��o;�<������M^��
SQW��-���t��ө<��F�j�lړ�*"v��~�ǭ(��D2ul�ب>
�pYD?�9,	�@���^u�C��	2ʊ�e�n?�� �G��~kA=����~��!��gS��_�v�fM������Q���^����|q}#��_�*�H�D,8!c����m����m��j����,Dɮ>2U��ӎR�M��.���{l��~Sخ � �֛Ȍ6O&���P�~Sn�^�����?&{�;4o�`��TVg�*#��ɤyT������gQK,��1�O����;UǬ�r���z�2E�}?AVĭJ]Ɂm
�f�N�Q^��P\`k[ia��$�>_ ]���ip^
�G�p{���s�n1���4��yi�4�AS���'fb�^=�:yYb?/L��`Zq�I��584�^�L��]b�>��	u�:��W5�u�!˥��h��l��9J��Z�D�57�&8���#�,d�������G�(�O� �f���f\ˮ|�}�ȶ��A�\e���ݒ6����<|ur^Q}Nok�}��ߙ7����� b�����q�=?ѽ_�".S#����7��f��JY�@��6_����yg��:���`�OJ�1.����dV���=
}������X;;�Hkb���܊�<%ҝZ&�#���0��!����N�\�wt'4�Fc��Z�e�j�2���xob�\��0v�?{�I7|���sT㠽FX��6�e�؍o$���7��?�j{D/��	9��W�}���Z*���,��l���i<N`W��y��p���砿���MD��+=!��.X��Q��X����P�'Z�������'��s�	9��� ��gN�d�$(eI��ү���ο��O�?���Zc�Y���gj�R��X0�a9�8���<K�^-����g�GP۱�/����W�5�F�B�Z8|�˝0)��6^�3l\�Ӊ�Mi���uSV�@.�d��?�̊��T$�M����ͨE�� m�xhZ�3��k .�x��{�9�A�zgq�)���f�;Zb�J��nڐO����?x�>&�y��zo� �4�΋�˛���+s[6��fQ��;y�MD���U�k�`�h�e�A��G]V|
���;]���K(��+��#RI��x����4�|�]�K���S�E�@o�!~y�:�*&�K�_�-����g�X��e��b1���j�y,�=�p;���4-� Ї֛)X��%k8��1}#�p4M�+��b����E�,��K�|w�@>�aqz��$���y \����n��7ot�DB�OX�������AY��W����k����zurz�&�7�=��[J��	��cr�hr2d������u�-aOXQ�i�s�ы�c�C�|M7ʡn��v��� ����@}v�In8so�װ��\zg�H�<[ظ(�{�_/#�r�=?|��p����%N"�Z?{���I���)�p�pa��)���I�B�s�E�N7h�����;t�yT*���.�W�mB���AV���'��دCK �!5|t������'I���V���GM	YL�q���&�fg����D@��f�/a�E�k������a}�s�DT��2{ј�IϏ6�ܮi�6z��t�̳=Yp8[&~����	��պH�ˋ�ȟ���?�:?�(~�q�����,��7��a�C�]A��%4�Rt�#�aDv��#	�۔��:&��T���a�O�^)1�պ���#�8����R������$�w���)G$��Q��b����MX���̡on���	?���2n�or|�c+<��2��fhW�f��.�XJKQ�`?�o��b]��ً��1��m�Ŏ%D��#�-���4{����D	���=��%��^���i���E����u?=�9��Pa㴘J���C!`u�ӧ:n��D�YI�u���{�j������Cv�u���	n�)Lmk��5}p�6K���AY@<!K0����>��j�+�	-�G;]I8�ȣ����y�xWx;�lV`���rR��ŒG��T�eͿٯ��U#�����VT�b��݋6؊��w��Q��czX��m�2h�r倹IP#��R++�j��c�RO�!�W����AY4W4��4����7��Řf���V�({����\���3�N�<�G�0�p�zƻm�x�_���y�D]T�|.0��|�|3����J���̥0�.�X�~1���*bT_�'�m�E=k�^�̋�C@I��Gg�Kq�?E�V�KE�Ƌ#�H�i@���g�KV/��${�����L�r�����_�k�$ S-���M#6Zoi����:���Mñȑ{lQ̄�f�A�8+��+ɎX����Y��鶴.@	7�F��ɒH����#�(mEc�c�6������.�Hr�ܙ���['ƛ�bP�*�Z�>�9�L%=�K\qǛO���Hc�q�:���8���U�ٴ�����.��V)5�5:��^$_�{��b V�9���㟏��6T&�f�mLhԩ��K�N�TK�_Bĸ$�ݩ�[帹�V)[�[���j�����AO�7��wdZ�W�5Bxk�J�9��ʮM���u��&x��J��H�j��j�u���#l��n0,�����d	�ܹ؛�R����=�b����~C�?��U��O["��-6���F�!���
oOI�Ww�y��`OVۿ1LfZ<>u���덣�P��u)�bM�t�OB)������J��$�Z��n}T[���J�����g�62��zK���>�?)B50z��ａK���Q�c�ɓ9���I��̬�Ũ���kuV:�NS����`c1�Ew��;��1�s��jo�}r�""ۣ�8h�;/�h��M���Q�.Ԍ)9�#��J�d��c}�vO�be8z���Gx�A��./�K~0��A
)���J��0����rZ>��q���r�^"�Ʒ֮��cg�[P����'���9.����z�/��Qb�
}|�U�.�XÒ���+�˳�2���Fd���NP�b��3P��XJ��Q�0���W�¦��3>���(w���ki���0��f��W�y�y.q� ��Az���(QwL�X�W��,��tF���G���⹗�����4�_SN�(�L$4�{�X�Ji����;��GeXh��	-	�ćkp����ۊJ��0>>jtERv�zg��7�L�D�G]�_����f�\3��'+�kTk���=����{��uA��^1mL�|�+��չ��?�G���� L��L��G,�޼3��!+�mefr@�!���a��A*F�>^��g%)�)�K#9+Kx�A&5��V��5�4A�,p�9?�lN0	�z��;ST5~HFHgE��E�d:4��TDtޅGwRL%�����f�Ag�:��� PPgn��u��W��R#�_!�#�֨M�y��ipF����ދ���ĸn���	�h�GR%�#�׬Lv��Ud#�v@hS�X%,gԐ�h$�\"�Τ�?�{{HI9���#�d���{&L���a<��	`kiM�Uw)�\Q�w{�oC�1"�>�#kb��$�?�/J���rC(�I-b
����E��L�ɍ���eP2��_�r;��.���|�è��b�d*]���	��*5#=G�n4*�
q�ACaj6��U�&G�K��ב�1+(l�`�p{)��B���7H�3̪�)�a�@f�N��l`7(���ơ�1��p�ٴMhK�Q�.sx�B�a���.����۝�����`���p�J�n�d���"����uf֢�ɭ������G���Y1�+��w������M���ۖ�N��I\:�{�Q�Hg�,[[yZ���R��Dz�NO;�b�g����*n�Y�q�D�B�Z��~��{��"ǭV�lv���p5,��]6�ݮ(�=�f�*�J�Tj(W{��!X4���ItX�� ��Gv�x?y�77'���vR��9&<�<���H����p{��x)B�z��F`:�N���r���v�&5�,��kƵ��Z�TY���%e���'����0�~�N��f�-'��a�֘����ɍ��ǟ�_�'��*:��z�o�0�Ħ�G��|��bK1EOv�/6�I��Cx_�O�_��$[���,%� BsJ90�ZOKO/|������&�/?T�B�͖��vyi4'�R+��/(.
����_<�e�Br�2<�ϙ$[��^F'��
��H9���9Ԉ�p~.$T�@��#��.,n��8���6��)�ʟm��Q�6x�Me�	����p���'�jZH5��^���'
���b��F�c�s0����l^3��CUo�k��-n��@	n�:G���\cn�X���_�m� ^Y�~W�iY��n-a����TT	���V_�lK�x��.L�9��vmD��g�𵄴�H*�,^�j�"�"�$��Y#�x9)䈲g@F"d�� �IGI٫��yrK��1(+�����X�	�`�Ue�n���/ܗ]���EK�\��3�c�N)�3� �u���N�����`�|!7�߄�b����~����6��/������T���C��/=�B�������'�'�5S*�s/V�����:������#�.Z(��`g��N�{~c��Ц2����A*�KpNcR�+]�@l�/��������;7I���h�VM� �X����ӥ4,�&kV�s4�S���T�0z|[�h����
�ِɼ�����-TF�{\�P���
�^�韧����q�dKi� �+��n�H�kj-wM�ɉKM*0���@��v�A�ӡ��r�Aeur��W%P`��4`@�	�k����&p#�#y �W9��B�Ag�Y�Хm�,4�x՜.�,=����'�,|(癿��l��:� �	��EF�J��;:��h�hIF|���DE���� Ϋ%�5;�B�Xo��%s�L-�C09A&~�:>��"Z����A�Eju�5�~w���J��"�d�{�xAkBa7���Q]��~���sr��������!:g�N�]�[��������ռ�8D/�.����~d��C�+��`�>�[τ@��/��X(v}�{��Jt�=�&�2S���.-�I��|M�F}���@�D��2|%���A�V���(������LM�2��7�01o��Do_�e�j���H5
��B��+�n�*2��$�Uۈz�N��K�qT���9��h�=G��nb�3v�xSz���qkm2�����O"��&<��h��e��e��������A�����p^~���5�f@���u	��'��R���O_��ɱߟ��v�cܭv�ـ*�,O��Go���%<��m%�\��QN�M�q��t��y��G�v��0��wpGO�l����v" y��*��D��_U����t�8����}��@6^+���$�=�
#4+�8��on�DI���p�pK����9����Y�o�*@���LW�yc�E��˓Kc����p1�1�azk���pn�,�t�=�K.Eʀ�%��y�H��
^��)�
��H#;�����4�~�w��4N�z[��}x=����5�b�X��$@��.�iZGp�ڪi���f����,��3��#`跭���t���7��:E��BaH�m��@��Xy.�oqJv:��8��,�v�u'�Z"�w���b;)� l��=?;.�~/�xp�ub�BPs����n9ja�EPnH#�&��IhQ�/�''��>�m]��3,(�4O^��#2 ՏR��/E������E��h��cy�C�]@v��P�0����6m�2��]kqi5�q⃩fn6<��X	���˥6�#�@Ó#*9ld�#��9�r�]b*�������aT�/ �F�����V*�����)�HC���Ҷ�6y�0��t�w�;��ϩ��y�Ⱦ�v��ǧ�V��t�S+��1F&6'�z�>ģ���Dj�"f�p�lL���>y���~��P��L/�3��AKl���U(�DI�s��Ȉ�-Ԣ����o�7B�}ϝ	πĖ�G�0�/T��Z�\e)S��+��� }������adү'n
���WI�a�{.��	0H���	_��`�KO�0�·e79"1�N�5C-S{榤.�M��Qm�~�����3H ��0Zq<o���s��Z�I�{-f/�T�@�@�����Oèju-*�\!�)��:�A#��q*��	6o����ē`�p&�;����1��Aй��`x�뾠h�#'��Q�$�,�gm+�0t��:Y3N�O�l������+!�R��p)��Cr��pZ9����u2���d(]]��"���)O��1ƛ�P��Ɂ�HF�E˙/��;k��g��.� ��08�á���}��m��mm��(�����w&�=,�g�R$����s}�	PZ�%+�	���G�o�g��ð��Y����!v��T$m��)tN�%M�j����M��g�*Y��
��<��NO �^1��ql(����^Q��lƀ�0�r����)�<!ܧA������M�K�|�_��_2;����_ƺ�w���:�A��,ʐgj����W��t��hG'��!��)st:t����B�ɺ�\���(�X�~�['p�O+S_2��}{�,�.��{����R� ���̉�=�Kt�~��[��M�m�Tp�I�󞫷�Ʈ������B3R A��^ւ\��d^ B�]xz��	b2�7��������s4�2�Ȗa����l\��	�*y,u���P�� ^�N����qF��0#���H�r��
���)l!~?����|��I�R��� v���;�I.�ʖ��?�-�},A,��pFBC�e6�o���3ao����$� )��� �zs&`�⠸��1o�I��l+d��.�f��˃�V~�jz�/�F��"�)�S��u�S�����g`��N9�iz��(�v8��'CRq�*a�tg��~o��!�rhMz+�zǣ�Ag'P��/Fb/+�>}ܐl��}�n�8�E��B􋿀 +���>��ab���VI �����2��d�j�Bg���-,П�.,��x��G9+�wϬ�����ɑ�#2��=�Nw����l�w���ʎ��#�O�|X��(�bI"ر�Lx��%�z����Zv�~�͵��hýB�$�]u$R���V��N�\���Ɗd�����R��h����"����r'��Z'�p��?�D�N��^ԷU$�XHNU1�T�CKSd7�	�.{���gJ=�����ă�ߍy���ϩڴGی"�Ȱ"֑�����ҚyRB����L6@BEçw; �o���r'�"2��BEr+����A������-��i�R�x������yݻ7��V�J%�?a�)� >e?��U����^i���[V�zd���gJ�}��9X�|�D���ts\C����.ܫ���� �(����+ �N���jiF�fi	T�лh�lCp�L4��m