`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25184)
`protect data_block
6oukF2EH5fBbYg4CbZAVsIagQjuC/3hsYb+qKA7L1whtVxiWrAr0FBWfRGbI3O3WbwOvcA4+XJm/
lwC/z7Gxta4QEdKFhOWypDgpsIR22nVNpe8pWRHpSfwydx40Z1fGXRL+KAYwn59PZEVCNc7IwQyX
CkZIoziLn2Rwtp8SBbSQjMlxYdUodekaeIzAbu8ysSLDmV/5mWZ1OEPJBkHp+/Eg0KPqF+ElFOoy
r5YfBptGnnpAT+339mfcOqsYFRYVrv/UYYFBNgML5ZssXFGzzJjxrBeXjEnDlf5gDFd1xB3CHmuB
rE5GJ/H7TuFBwTjoF8I7uZLlfAaac3Ubj4T9GrRday+RqtBn8RHQIJ0zszLGTI3RG8xdNn/fo37t
rH712FVmua2mDGvZo3JeRfHNzbkZd5FMbudb2XhP9WYdk6kBOHKKZ8aE2BCrhtabOUoadozoKV/i
pEBgkPrylm8DGhvDlEx5qJlwP16DRYJJ8fthDCgsaZQN9CCoB/cjcYtgjqIlalus74Mu/uQDc9KR
A5qyQwDFTjAmDkHMDIASb3uSaUikPgEe0rWE4pQhN7iSswgw2HO3LRFp4C9y40TzzIbXgloHXBrW
Uy/RaR/kKqNGHAydb0Df/ftS7+vRoDd3XTCqyJSSjRuE70lUV7uiIfxYZ2MV7ktBYiGD4Zxv5CGH
IcFxbI6+mVgz0TApTqIeZXn9PEguXd7A0eGZa4zX9mTPEO4OICY5+t1euRl5ESo03/zhST8U6kiO
CP23L3/945ZVrE+HkNm9/k7hKXAqCROwYikHTDigWuYWJvmDxGE8pzWVk1E6brVf9GLIpWb2J3JG
URulba5SzbES8rKUHXLKXtwUoa0cqeTK2TBeC1QeXXJOyyYSpKUwByjAfIzwdhlaU2B22EqAyBDo
W9wuX6GVNDc0/Weqcc5m6XDG+Na4GdL6PDWzy9ApBWEC5/I6OMWYAiO9fXBiz/9GUAndXhNjkdhe
C7wn0xFakhr8tP+eAaEmvIkxfx5W1pYa9WbqhWI/cVYZ9i7xuYYWP6WVeRCbX3hiOJa/45dP+1D2
JfR0cKaNoFzATjkQsEI0UtJBxoyNZodwFKqUKq/sE7sP2n63B7Q1JD1s8xthDcCE+bMR2nfPSNPR
r4ZPiaIj2tzwh5UkK/J8p9VJG2JeH2P6IBrBhLHXS2qNNHU2YKXeAmjpA6aV+JqOv4VPDia2K5VE
9e9BUSjmWw1eh21YJVOlYHkXQ7ZlE1Di9Wz8g8LL9CutFUZj+Ce2gIi98fSxIu3dusXTC/CulI7O
oCfhjD77cI4txwImDh2CPveNcub8CNpvi3lhy7tn3z6llyPoM2tOWPoxQTyae0IoS0WnKHOv5SPH
TVX0nJYGQx1YztbTv4m922LGRdNOrtlydPZmZCihdFku0xX6Xe/qrXj6HK2AC3WLd8L6J0j/kdCe
GFBRuEfQ9+GWvkHl2dH78WGk3Ss+00kpD+Pzpi48TlOVPCX0I4OLXdP7PGpoOJOb9Mk0knGgs2rR
1aSyj0utDxwK7+GfWIImCwU4QRUNiL+1P2c3WbEY2hGgItFUCAW4beQXgkTgJ5tjOuAbIjtXQuo0
1s94NU/itSP+AHrmv1SZP8U/Ep1MNLWRrNn6xuNNg2ECJbAYFgy/q/3GMNb2SUB6MlRJvVWM6nwm
40scdDzZdadCEehKYrhi4VzfcfLt9HL8tS0p/n4oaAXsFAnlXu5lWUhbiY5Em/CXI1Bsqj4ho3p7
tMl7BCmIlTyPtWNoD56spngh6xHTkTqLycR8JQpBJduvZg6LPMyuVkxn7ZW8SXMtI7XxNut5xdiT
qHkUcNSe03ivAm2no//l3xBHZ/q7Z3XjFkeOehrndvzonk6UHMevEINHUQ53oeYSfXETdNIGz42d
M1Ktwiamgss3+fgeZp4LVE7xcwbX4LTKNOcVJ0N7NfasyTT8p6gYvyEx3AZDUh8rnUeqJFAjyX3i
E3Qw0C+yJUoKEY+q4RomxzvWofSU0OQrIUv+296nb1lr0QoKGI33509eXQ8jUaavFse6YeSAmNHL
bwzm+C1x3M0VGa74/zzyO6wLl0Ku85LJw86Sp6s77Ilx5kcEi1BJnOd7e7iLtZ2ZiGD5kBP8p5PM
OovOXHM5oqfDVv7g8vtCRpFZ9FqHFgnkOvWJk01w62vnmuG/rb4IraWKLhVsMVWMnhtD82+75xWa
+s7jXxsReXceEvxzXapaasE7+ysUT+stXa6nHPN5JGYecOmPXq9CIiU6DInxvrSsbWxbqg+unsxU
UqoXuX6nJbzqCmcmcR8JruagFqgclcmvOiNCjLNzH0DpfD2XrAp2t+VQz6KqUU46RGkE0DIW7xyT
asTR/o2l1jcXkUCaymF1yEthtul2DBllF2YL+XJL9NTWUfSo4tg9VOw5VN/Bafy4li1quAtzcto5
eltopn67XhW9Kdmk9FEFUcoTRUra5vqTkvRh2Y8gjCxI+GZ8vZCHFczIzUU7nbXhGBZHMMkl/G8f
vObB6+dRR8AuiV6Zdz/NEJnmN3AG7SiWw42Oi1IayVoclULc6uXXSzmn1PWblieXqN/x3qESc3yM
VwXJyjyEdZX/GtV8h17qxQK97Af6pxjr+eQLTLnG+rjBJmuxmN8kDsuJZNjUPc/gLvPtL2dvCtHA
iuEcljogoRzNGgVyH60dRsXH+S1kwGhoWSoCy06BJWY/YX3TLAvg6omj8NT7VXml+sh4qK3inb01
vR7G+9jFe0D1vWyGSQW/Cmo07aQtoJlxqQgvR8Bel9DB4mru677rnpMd3H4jNEzG6fw1+xji5EE6
7kricn6s/1wk66JLt5m/Lvl7eirNf/2kBew5E28Dt+UYveGCrc6PzvUA+wgHyh1zzfC8H8ohnMs3
TO9m74bQDFoQsgcQBK3QrY121d1eZYcF/zZH8NvDZee25p4Uk48yWuPR/Nh9gDX/rkdeHZ5O/68A
ruNJZc1LJGLEkMg9SeQkurylpWaOdpRpS6q3eq+Lv3bly/qsXvytW+Wwygh9Z2Idn4VCV2ac5r38
i0q7OarhoRCDZp9vHAQmADPDS6lcK7JGgRAjldX4q7tDr0i8rsUBJGatte2ajsQcsxEZlHJSKkW8
longWt5i7XSj2/VLorWQIT36C8NTSlLNpn0X4FRztvjJ+hFdTDWC2Wx9n80LvstxmSicc7RutGqs
Vo7JIFCgvXodjStOi6YRRqWTeqcLn6ymGAojGeqHcnOe/FcIBqgBD7StB4DBPJfx7UpbM+MzL+gx
cwejM1CIbZtwwfjYaRUlWCq0nk3pP1dT351Jlml7V2Bbzjz9ObVbTG3kkyhLDIgqOpnCS2g4CxHK
A+uZi/cBwj7/XvT55jKxnq3+oEZKFMb+WZkRoPtHQaHLFFMe0RxKstX7IpDTjbfBYj4jjXDEg3y8
ctnEwgb8uQltjp/jr89LcKUn8bW/o+d99mDIalO2SSiLhO7QW7FqR6shEd9y+W6tSgvBIZjxHsGj
VFnAyPlj9lqVuBV+dSSnEbjUzlnQNsPLCOlPbgqZ/zjIdJsEvvH/gLj6t67CvaPa2sIrZO5gb40z
d9mNLBLPGc54OdI4q/t+Ok9uX8Nx4202LmzQ9FWeKmgzK1EzJqF/hxn3BQ+0qto/TQupH/DhOXoq
QKTaggPzpFB24fjVBewgL74DoqM2QkbccfG7zXageeW40WnRX5Y2etS8iGTCFdITtR8ocBlCPU84
3Qcr3wUs0imJxzceDSNUC1GiwWbPk6xrgC27z77FoEbZtglXOJVTjr6mDVLTE9gbfb9WXDxSYl/p
/LQeqxQvEUYEZuWDWRpKLivEXe6lZ/lvX4rAdxd9gRvwqOTVnSZV3Tk11HAoz02AVm0wxj8vf16e
lP8EJQrod+ieeB7Hb+92KegypLVXPeiCXlVvlrCvI6ctmByUkvlYRzdcdXvnYl2j3lm6ef1uUa8s
2ke43udgrNoYcaTyTxec0SLkcNdllWrv9MvXbAxyL/xJ9v5Kg1BRT8Oz4qVyYFQ/iDGTqMz85vuS
nqaUDRf2Abr4sjiH0URBhZzh9ZbbB+t6fnCWCn124fQKvkMgvVgnHnJgfQAAh8YQAc1HIX2gyjJL
puoKhSnEP89Jfi27pTIlmXYaVUCDmf2TpIHnrR4eflilpwn+u7yNg08pQvsuhb2YMEvxorhsaG7w
ZaKI0HfCoPNN5tDWHLAfje1IMd7LCK8l1nwXhEALNatfvE+df2zIR0Zbs7W1Lvg7ZtzopI9nAgEz
gtiFpZqEw0vMg0ak4ncXoKhdq7Om4qFNGoWHjaeU3MJ731T7y99YGeiWMVqXVxqM2wvaiJQnuFy/
Gi4fB0r6aheCa4PHc6EUbjs9k/zhkeXPTFOG/uT4PE1CCcgQtfabeGgC3x9XNqUvjiS/7gP+RYzi
n5tyTTJDGGxvI3awfPfD1z9wNYX3SU1GHORZa0inE14YAHCrB/LQ3IgAQArTPZAy0PPWHwowkFYf
FG1kh2WhbcVpw/eFlcvTtuFg9e6iWgtBvRNVl57oEKYIDxrJ2frRQ2Uj3aw8OeNaz+Hq+lkMZxYR
o9n2NPtdq2Q70az709Kkp8lQIiCpFr+uvajbxMuP715xYOrtccYhoEkLuO1QFbPXJXdySaWitc8e
zxiKXEwQC5DqB6VjR4YiuWfs9cCl1x2WrrdgolJLpdhwwOqDd4UtxG24ma7Y3l0wexRScyWgiSkk
tPdBT8tN1lG3YrgGb/Tt8Rnpjjz3UX8C53xeD7smocfjY2zIYGutMCR22Qi7i0B0WnVLVNRuG5fO
/hugahJDAQpm1JvWeoodLynwbyyrA9O4Bl0oCOGkscPXRnXIWjzK+Sk5PzY0W3cjK8BHFYG2BPVr
Rgb3gwtte5aFWNz7/DTqowklfWUcnrdZntq4bXckp4+h6gB4+XyIQNKB4VKNEECYrDuYwUi9JhNY
1Vw2b0G58ZrmYrmT9rFGRrnTzglzLZUr8wzZPzkPyViNF9DEiAl8TPr2lA1argnVRzgmSx2y364n
muQXj3Izp8tA8DKxplZc7pn8nml/8FP23VLzu3laGRwfRKCN23BMBbzgiFenthwcYVsSMNONljzZ
LsS0NzzCf2KmqIWITVVFwSP3BEB7cjTXKUXBahLOYRTMji7F+ItpYoie6ZZnuoTIx3/v0pBUDF9v
DLpSHpDiVa6A1FtpXrT2jYUsdq19pGmUqxBdDNqZchQF76fxIG/cPXUdfpCjLnItwWUiDVkXVvzw
T60Br56LKLQ79+hjRovKdQGHRsn/NkvpgOWs6P5BUCnz0qgre7FTI/cbFRpxX8VnvK/0/JJEturi
AiTezzR+5SxjubqDPO+CvBeNhmUN3CxwNZe1hUQLIvM0VlnUfKkRBV0t/4Umrena6bCpJR/l9n9U
A+KF7zMLT5tYasfALF97vIn9M84wq94zs/ZPf1EdJZxxfTiBTaCLPTND4MjxPM9O53jV6BtzwmAr
7gLCHLSPxTzToiYj++LBUViYbBv/x96y6k48GbeBkqmLWGfVdQqnZGJ+rsF0q26pC2v+zt5B2JV0
+6RVIQETnL3vJSJehEteBjeWKv9rnkbU8HsgN8E3ScSJMNlKUExDDOA6ppQ47w1fyJgTzpxbclZ4
9DymQKUawWR8dOs97SsU6X72ZW0uGwTUn2nnTRDxvBCNpveXfXXz7sdMDeUy+T5mzoZKIslBFl1y
I8CDtrmvLPcZaeD9xRJJ1LJRXS7tOIVeFqKuNmONNL1y0+FSwZaJSQTlNlrj4ZXsziOQ0/DmvkwP
/eg2eIu5aFMfBr+NLnGTa028u4r0K+CBWcpRDkseD/mCneCEAFoWQWVvKSNgqxc2sKdA+gVRlcFt
AnqBNRGqUc+48IT3DHofhRXVtrHzjA3824kodpESSXx2+KNU+dIMGRZZm9G02UZ+1DwdFYhHCQdw
KFqQexJnYT+vNIa31oekaptzLuzFJ0YUIL2UgYh7+tg04BTcJ+gbrOGHT9/AjI416uqCbrTeHkc0
9vV9SICfj0T+gOR4LCarw3IpaVz4mAmNaIkLkRSZadnGHsi44w8PM/BHG0nm4Pky9SHDFjPz1pdb
wo2ySmkwFqnHzVoDGSk1thOuUFUMCYTW8rZRxNxEcbJ6ufYn0Emx1QF1wrAUaAyNjirsl+9P+255
RYS+0HJSUb1L/PwKC5Mjxsq0JAstO3DG3z6IFeK137ahUwGac3leEu8rKIIxFDMk+GJRoA5TUUPA
i2LCLkR2Wal5csAJZYDkA+KiuJ3hmka57HzCJwMHA+PBlETHAMzttIyPLdaBKETEhdmKFWtqjrcW
2mDCb2rB8+BNQCmT8Uz5QZgC4bSnw+jzLLSITOjag0VOl3rF7Fm+5xLyd449bCJr307KioEjt9kJ
GNovlOIN8ZXoeSU2CriToHJrcCrx6txMiW2gD1RCy0saKLh/4nQCqCR2vjfDCVIVOomvW3zwuUAl
bzLHqIfK7pwelsaa70xzTvBV6OiRykjRuYjQldmtYlB367SGdbaBJ53JJlihXi0qMMezxduztyEe
fiXXyJU2C/8A9hTZ7HfC8wcOPdMNWb0Q+wSQFXgHrljc+i6IIcswyjYzhuss+93r2G6m++8uK736
L3XzM/VpvMEsjb96lku84ZlzEH/jGSc12dGA+T0+yL7mGMbA+2i6uLnCPmZsoTrjNWIH5KIWq6I7
kqSrhdmewLwDu7m5QHE2ia4c5d/nWY/R0fzEGkVfEqguVdAyH2QaVyGHBWnuwepUJw0q5SBTeFm8
BhVJgv6KVUgXwijl+01epN1mKSL5bNrjwkhfUiIwi9GP/S3hE4l7EiOQtdS2Jt984bRRPhaQSXoP
wmdez+POhiah3eT916hSkDC86uKc/piasJCSQJaj0xD7BaKx0rwbXx+3GhC+q2lFVijJG58DjirI
gGMumQ6aNSAZLGMY8gLO0qkAvyy/VUoo/lr1dSaXZULfXdGX1ftfZNgJKseYrUjXy/zEvJlub4oH
CWofyK2acpRt/flaCuk7fL3O1dYXc/FbLmq+Qktb4S/yS1oSDvs9G0LsIqagmGHxFpSUDcStQyf7
hP7f3PeEcaLL60u9gjZCUGSmGmSdgOZzKjTCPm7bbRHJldeWnP1CneQFK0P8WLr1XY8U3z9Fi398
n7dESVQSJT8bGVJDHZUsqJTtUuyrz4nE3/8L+udMAWpD04GhJTSbz2t2UoI+773CMluVujiiMEAD
F9Wn6dpn9HytvAPkqCMMp0NE8ii5uRwXG6+WBVxC9yrksq8RIZXRSvJJXm6K8M5OixOAxxYR3VpW
QFxZdIYTqFGVehSaytee1HOKxU3ghf9snhZoxdlGJzUpkvoP0hpvQ0GNtyOWky9HPF9k94+bm1/j
7JCcMrgm0wdaeWkuXzKxnBA8jRFzjZcCrWn0j8KMEznzUPAPd/xNE0b67cnCezRlEPa/ZOqyrV9g
rwmo1OChxZzQ6HdDGinIrIYKd7r3IaVX170dbYbOrkqIkuVAYfx4FYIh3EApkFhlaA7XdqTkqm25
B4swHCDACNLnSxKZHkbQHrOeNlDWoUi/EloQweifpxL6JQpyVOVYlH9V7owzl5gUnycbvdMaE4gr
qWdH+GBOyvAUSwWVTFsfVHoVD4DqzOLbJ3MAeduCfR/837PYvYUAvvk+OKcnIIbQFANtES9DYBU/
lpK+cwvO2Edl3sx8PEHsyiWljdVnWhsO9SsFYZbAUrYbvDgSXGxHlD1x5/ED4t2R9R4Ogx5FagFd
p8kcvTsRE4QFtWffFUNmPGEy3BT1M1MA4ei9oAo2z9+AJaZ1GfwqZN4payM90BPXZ6iPa50psH0f
8ejRV9iofm6ReOy2l+UfoFjFqFXoueYks6iTiaY1G723WB6LTwnNh1Kj4wftQsy74HmyOP5ZDP1k
OPH8m3tsXyafDWPdm8WCGoz2XJgSLcPXn9VEXcNs1b2++jf0NPJozIjQfGlzoJmouR0kMY3UptUJ
hV4zuCIKtaBAT4a8TBjKInI16v1wRrPOxDY3WQXBS8lfhy+tvmnO39k8H6uvKjf2zvEKb5qV5nyt
XqbWDz+buypdT109IkWnCov+2gVdpE68y+m0PxYCneW4y3bMQkXp/bNw+n34T2ACT4c2sZ8TaOjD
HGSnPPiEmO/qxZcm8C2ZMJ89d4aXQPWjnyWlWhm8psgmdqfq/P4fdKJE0+zN9r6gqgCT1Qhw80NA
rC4wLI7ZYyfe1m50PpQbvD8zcgRPcuf0HQx5eaEwuzJBMNzjig+r5pHVTbWfdFBEbXAijGcc+LkO
O1lzbB3+Kaa2CKwxP3iKhqwCJon5GZpnQZAcJpsWO+su6loIsL6/CbifR5x+Fc982VDj6/HKsEfy
J53wa5hmNhmv2wgVmz/AhS1uh7+MRb9Vw8ED14Y0oEhDHhTFBqn4R8K8nA1VBzic795WakYBMaw/
pQaVFxbBGIzbBCN2MrRI8xIYbeHeTKLJG924D1xDY3158fOLzWGXJQfL+RD02vRveqdjgYV9NtKf
4gC/oEU5f4NhnrK+xAfQV0P2n4KX3Vd2utiEwgZr8w66Bf+XDBqYIhhfQLPbP/matrmCDW3Zj98W
ZJ7+U6ruvUjBJkEKa6qtbkWGglx7y3+w4TqioeQHm8yWyWkx0/zfRCGuaUyMSiYsbZPp15yuOgjS
eEuTdmh+nxypQp9n2BOKdOe+JA9EvNOKM9sx7SZeQhS8qqcROYD0Z285/EPSqtoPohtKfxMnVK9v
0mPDL1H7ewHr+BAWbMt45RXdxQD8y3GXspjFYH0nCznCCsHYb/T54+YR5S0iCzv+Jt1OKR0ApRON
8pJZxTQF95MRFOfxa6g1A0KXHxfiTibMEQc8ONH23yjDQr+XGIiAiezY2RzzHRXxOnB/1z/NiaPw
ygrMahHZHQWhLbDanq09Xo+rqPfh+xeaxuQwvVEAmR9ApzC/NUqjwqPV2j+ngnbB5aU+kM4SOxaZ
1TlXTW4ndF1f2k3BB0SbqHPzedwibwV1PlcPoGvsVT/C5HmAGuTk2vYhg4VvzP5aS7+K9B14DsNc
CXudcsdmn8+BEFPCToINh7VMPWGRT5j3wxh2mFAu7vEmlsDckur/TJJ00Bz6wxLEKdn0qeRoplkJ
cpb993RyW6s94rBgUNsfUBNp3bcc56TpEmw2bPB2Mcnw0zI0mFYaU9sqBxFhZSkzxORU/lM83evI
+DI6P2gkwh9+w9Kd945l1RoU5EXQgS/ed/BjEN63IpXmLbLHuwbPVd/dWYPfsGGfrfDgZeQWuD6b
3Etmz0L2iL3LouXmmLxpHtiQlbHGZcn46+k45FAlnDdF6xHcdoOJnURXWHV5KvwaFw16/JLGsPne
p3lDcqHR0VcT+fg12KuPxHBdMES2Pon/wkB+hsAw2jOFrV9yxMc9jFWkIcEBRHVmVLwYo0waML6m
8sHKbmM9uB7zI3bFGSpZz5zCJmEGwkLB6J0GgRoqLEmwLoTQiDS2qGi5MhY5UNPNTY7znYZaCtqL
ovLfuOECwmX3uTbPFVtkgLzOm3gzHJmL/2wAm0mwa0j/2yFVBa7xNoYXwbNyRr7CLCqKRBBVhE4o
G7FjJwcWlAYRxbk1Eqi27PsnWRXCpeEHDPhJJ0K/cYQJwvOnVZP6LwyldLxpKmCvf/TXsNo/W9Na
gimk+RlYie0tLTC7pR/rRfWmlstdgk+Ct35Vm65YkNSMnosXZPKJRa8Iro91IYxXqHc7Us7q6JsV
7GnxPfTZ2kg1klIAky4WdhUM67OjLhnMYi2Rn7ooA4RFDUBRg/hFXq7krwX30GR11pRizN2t22L7
CTxdhsGXEqDNLUCE25McIY7M6lbuDb+4f6ze6DDBf8RDBcyeCuv4xvxVfpYvpAUZxJdS7DbL2aJJ
KyJ5FBGi7x8qPUZuKgPEJXl9o7EEje8XgO2A1pkFhpmBJml5N/IvRozmS1mKClwvZ/OpLUPiImVl
HH/e5mEzfov1OQY3+GCpADZwceRsAWyVyOE+8+C7YNBggZURYvpEww5sHIrua/1oZ3f3xT38OmUl
JHYzGCIVK+bMPzacvxUe5KdVbNClfL7OF27dDoLaaogekwH7zE5ZjK6JexjYyEkwQw2xjs1bvuce
sGhmyy+jTb1PoWTjD3BKIhctzTJIpwQar+Teq16XeUyLEeYl58ZDbAVr+SEbPwSCcVe27SYt2JPg
ssPWyPtGNZXNAS5ZJLyutBF8Ji1dO0aBhJkpCsvlclvH1TJCJjivx+DAcKndqleEYNQQa4MjUzT+
+w9k44XyMKDCSQKTsUdyCFBnKD5Dnj0d7yDObPa/76Oit46uGZeriIVCfUh6IEPER/6SsX5Wnv3s
tu8erVIhRjsy2UBt/K/MEPdJsNthUVjngFiWj8UPU9K1XSJR4RRoDhXShr8wCsh3wEx0Jqmvy0tJ
tYPenz8RdiaqhxjSbIwUCVrRIyM4uUMjoF5eNh7/gtd/WD4a6aefYcHJ+UtYN0FrsmheimqCzwqB
5iwH9LFhFeaJ9nxLHygD6+te7nq+i9U2bPWDWfm1mKI1+Mhq1eRSaLb3qZ7qJKb44M+StW5pHhN3
vlBYrbDKlPlesoCiwNTWs2BnkrPYse4VhlS8JfTRcn/Tp+SG8l9PRVDdXzvSEtA8bR2ne1WREvOB
zI1vvJgwFcXvYhxtL58C13E2vmXkKwukWfEGZRZ3xZgv71tIsguTgs5wcSCTmdIfXw8v2ttrRk07
pdNMGczMdhQFEMMAm7rIQSKyZZ6pNPpQWosArwMYN4+oeYQyORpoMqUapvlBa2InX0Guwo4bFNli
nZJDe0OhDNOxn5eTAMeereh2+W6v0o02kh8H6E4yqlO2ASmeI0dnJu8sFTZs/OuBKLvBRtLuXmq2
kye7r1hxZH9B2sdhPYiyekTtJXVuUada+3c7+Z10ucgpRZKNxyRapfJxnMBx80sm+QFzZdf3/UDb
iWQQBuBK7LHhO0WhUuXPpJIXjZKbtdDIEDGTEpm+eCY2eT++2PxmV2E4ayw5jbE55TXa30ckwoyj
fuyWmMsCpXPP8ut8yRmSeSznFcD1spF0ErWZfApT5FMNrolqfetNtFYf7TxjYomnxrqjDWnW8/Oh
HQGb5OsneVTUMmX+ZAZ0NBDD6CN2G4DdIWP9/NrekUaw73FzkRkbCAzQYVmkjzesU4I8aGXCoDkG
oi/0zGatTG/AoQPY/t0ZYBpmm+FBCrq7EaVhUCcdiOw1hyg+uRsiMv7n59wfIia0L2alwkErGlzT
51VO6dD9bE8t8/pR5G8IfBnNgdK7n0f8suH1CyvJ0F8CGjsR2IQGVCfvKqQX0rpw8zvZSqIo4w6b
2kIsTwxm4wDmbaGe4zhJxpUMVoYRMVkUNnPEprmHt1JA9sY1ULSP7Plb/U98MBZRHuUbZQ3RJVni
iLehRV3Qw94bDkPWBMWCPIKW0YQFk0mYr85sfyVHKS490rCuQqvSr8V4QZ/F6QUFIo6s815xmnCj
KPIvmK1j217wNZlDhCBZQPShLG0Trq1m9arrBkHHg8R5jx5oWSlc7IQtbSasraIIQFPweSPKhLmF
pSKm0BUXHuTu4ekKgMgA5g17J9aL8vGKe0ibrq49D9cZlaw9hgJP0mU+uoV1x04ud/oDgky9xbfm
L4tln7NR745d+OgmSfZFVc5JEtFyk3a/osoclexZwYlalzxZqJnjVp5Kg/blcIW7kL8QomzZNpuZ
CcoWqTXJQuXGaC2EL5Kclv48dXRKqK1xmcal315O3ZhVPqF7fg31mIto2kceqxNjGtXAtXaOe6pT
lsoo3bqi9Lz7kpsW0ci89mPLyE/rejHnfJf4xbPyGqtvF3BKGz4pxtw7q8ZeQzeZc5rNG/Ua63Ih
owdPVSWROdAADPrpAU2EbxIGhhFyFebUEQZ+i5oGUyLp1Yf2HgS22PvAPw3HCuQr97URKJ+oJ9R/
gaEGmHSPTeb9yYjp/rsaogsHp6AQbrLYeS7JqYhtwCol2zOxuZOT2kXdbM7vPFZuqFcuK7ZzPE5Y
3EjhDiPfRoNRCUXJ6VChXImli/bGmypkQhpwakrWfjTZlJg65/v9uI5M3IvVf93SDv7fWIfBatde
K8e4ytGJJmu7pvuFCPwH2sq45UD3zCPe4ku2uzcIxwU9aIVqXlBKSDLOci6pRy2OPFLjfQvVI0zZ
6WjanzIosot4LuZ3xBeTzb0c5K7l0QmYQ869veMuxEK2SmyFQ0v+3t4V/pRiw1OLZ1oVZaOuxvPy
8cJZ+YM49XTFVpJV46wfGiUGpDDQxXlsLhHuAPdaLa5jBIOjmL0Q8bj+vJEsR2reF36bM1vneibH
xscvc2rZFTs9YdokrhmIY3OfhzYaPL5zQ6fJ8tUfiincNqxX9hWWnIoNa7yNW+FciYNfj1fZnZpx
FuMJt6EUl9CgqeBLhbUtu059O5akulcdXsDW2wO8Q12wgxKOHOk/bA1AoI0UjfrCLAoB3I1XQhyy
StW9YLt1DSl95P47lfzVhC0c/XXSCHeng+i09DB9qWfXc1qb2Bl/ColQN0c+PgIiZKuxUAotLF/s
72VD7cusoX/ddOJJ6ZxSsxsZf8yQNQ6NNSEj3mMFV9/72Yw6tK2cLreE+HHkqZ/ycWlwjrtnvObt
2ltuNqgjXxR1VzBXI2DfG9w6nzLHvWJLJdyxAVS+IdC+fgXwjAXtvP6+NZksabeZQiN7yMvjov11
e34m7DaVPwYkqojLHZeyvOkeqc+SnRvSKjT459lOokkOrMNRpBRydgyVFWiGPceTbTeKzerh1+xk
nMrVmusn6m3r6yKA6EpdlffF8hXk7rV98w5y/bS+WtfH2oZjVC77OUEgT9ZWYmbDgMlrJ5ROpUTe
IihFRp8jAtE24zBSUbY7FJClAk1XBy+CJ7S6ig9pAddAiBAPRn2MFENC6t6HPEcbF5Izuc0xCNcp
U9D059Oi4xYjscnzX+Z4aS6skQ2W494ypiID4+7oQcbXaX+vxLHlrThqhj8ybOHtu04jkIh53FsL
e8oE/Z4uZb12SLZxcTGjT1m3HvTXx4gq2FKirU4vIL+t93xxxcLTA9WmcStn3yUJy2bvu0qmFGCO
zNCzYXxqe/h7h0icbH7Flzi6VrvFoEjOyaaDJZPCTOSAlfLWC8Blk4HFZiunNupZTaUkIAWbPqM0
+BczMHdTxVh1sa0oCD7xIsXb2UUWmqRZ9saerj46gc96s/CGOfUTJKKU3Kzg21kMCIiFLi35OrKZ
WPFCSyPmVn+JpHRvh4zMqokilUcQOFNxVX9/oKdMQ0vGRzhM6nm6H/DPz4J6NVdrPZqW8/vWz57R
+5teuCaayEPchVF/nPZ3V/iR6lr5CNZZ0nMos7Bx2zh+8+SrCqesKHuN2Yaec6/zVB7YXUnznWog
C6rscdssOQxj42a0KRklMQnPDvGxwHcRW5R1HkaohdsJ7MCprti+5INK6oQvrmFZIfqJp0IZd616
osAhMIahec0hhezyRCawmYiWtq8uAk6XYyXj5fwkBKiAWPmxrWNgdSLMrz+scNEws1OoVvg9xCKs
hytyA3mxr1so6JbTlOEQDW8G66Y/EnDp2Aq0MDckR7I6Hmv941EpyBbfaG/sAFyNNpqYJGlqxZS5
fa19b14HQUthSxD7ne4IjAlSWaLxAwwx+Cemvsgir+gp9s4l/9NBAlVuZxSHzAW0oZBijZN4R7Pw
wvhAeHq6oG6NwKNqlwVo+m22VSA2vdTGJm6SXu2oiZbRMyZG+GgHraw2tGCPu2tD2rnTj2SUK4lO
toLtZby8YgxIa3UlSqVE5fBB1FeB+2ZN/c19TsSjoOX7tX+y1YJJEpqgfo3OLo2CM30DbRRpLiAg
fOTzhzh2kiBRD/HXe+ZaDaLsaqFSKM3vGX/ok3faCxhAI1yDzhGdpzzAn5wYzA02sYw4mJ61GYVv
RaM3WqAr9rHb8E/BUoaCboo1qrC1mEVJAU4PdR6s7MhyDgXLe7N3AWvlbomlWFa+RJZcx46QOQz3
VSSkj4VpEdwXU/Nn9eRdveczMjIG+rtl9N9lJpRSku8iJ3W48h8q/2DingL5cj5hAYHWDD9SIwHp
JH0naXY/wwx/ypTUDvMdgVXJ9JQEDu2XdsSa7Lr8UnFc4Zhl6sOpK9lv6C4QQOCx7wk0D91tLIRi
Avun8LqzlpQdVKNQyfUlUWpwHJeqHZ+gwgquqZgzFQy07mgwlhrmPFOEXt+DZVWctpOnIqdW1cDX
D5Rlkkkd7m5C6w2GqTfggho0QNQh58tmGhw5NNWXiU/2mp0Lz6KwlaFqe7Leb+J/vu72Z8X6EOlC
vgU+EbWi5xIBewA0fiIdIYK9b0eti5M/uvVWiJpOHJ6scGVMic4p4FZWbMSVLFAVKiJnd0mxH/WJ
47+/N2+ZS5qIhGrRbKegRUP8HqUD3BhRPRTUSxpVxrABrfAP88Kr4WOZsK3UnQYvpOVU1if9dvLc
pYFKg7XDOMOd4ly5+/otDLyubgdV8ji1Y+adWWG7hF0rbfRPz6xJo3vm2nP0C/ifjNzpBPpCSjs+
pcRFeSH41OhDf++3lEiQWCwbxs4QJTlDjo/UYw+HKCi4orH8mog5vx6e+lWnfyKNdZ8NXTR8B6I3
jcckGkznHQofUkuMhCCHoYo9TYC9S+UeGADxIou2uzKOUTs0rifSF7gE1WBHvOej9F3N0zNhErn/
w/nvNbj0eFhBOgT+Li83DRtVxKogpM67DIjkhw8dmFv/4ujV5gGzPDMXqn8IhrkN7AZ7tBBKMBTR
2XC7I4yw4j8y6/NGdR0nKSGLmwVDnirQCZYK4ygjTo/WfsA7CWul/71wQkWV+hhksPWkixEDcIvi
24P1sgd7LoIpiujNFpI2+YSl+GHCQve2fX8Dj7WPS4yUuPvxTXVrsOAj2fUORxf+hPCzXxby7AlV
yBdwSvYxzvA3I5qt9NnIZNbb0Y+rDUZyc1AmPT3Ok2m8C++r6YSad8Y2V9z7c1xgQ5XydqaoD6RU
bTWFqAGGAajWn6z8jtfYNxcEFJ103+TlhRwz9Lg2iXZZMDIY2C+8pbcWL/P0OMq0y9uITONr9g/a
HvW9Flr5sTljBDR4RJtCT1MuQZ/xvXIKi9k9wXat9yID6WI9UsdbR5UU/Bx0LG1vAINZlxfdgqqs
UDN2sJSHV4KM7tFPvEylJ0J5EGs2bdjl6yjiNm/azMOtwYHu4RA51vmJc4gGOQBaig3144Frodr5
LBFMkU4e33KIUwRt5Vtdm6rKSWBa3tisbui7CtRaFmAZJXo1ipujjRep/6quoZS8k7iovqi5HNJy
VFStRxWaEGLwlS/IYaRVJRdUx9G9hL121CDnTF28b1gOGdg0QLZduvMYVAj6dYlU8PCwe5zWYc1Q
gpc5aGpyRye5GX2J9t8VqchiEhOL/l/mhhjCCcynITG7VK8P2ZbosTRDBQZxjJjKWsT+nVIZ5Wnk
fgLxjXliZ42SukTOw8SM2sxcOs8HCwYbwbuCgiYKqEkT8/LHk5UoRitBIWt0IrY6vWYbA/mlU/uh
s5Gv5+gThIDW+1AeOsvInRhXHNqy2CuFCDhsCUSdLD4+vvODElpvUEkH3riNI95CGMYFeK5Lf2A8
T6206ML8dJWXszqzPXLcWdT5xT18kjYpaPHvosdBSYZaZ+31Kec3p4bOCpJdNrD2xRDdL7gylvxn
CpIVZ6Bog42AxhG4PU9IbkX2yUCSFm0KKez0TUytUGTg5bdSddedAh15LePdK+xOWY6GUNtTi7bj
K2vxDr38cO5Oc21VacUAgMF+jJu0LhHE3o7TP9SOxxAqBT72m+62HDM86DIsU3luimF4zPESA5Ve
j1WMSCTFK7aZoa33N0KdQfI/9Fz6/BnWZ4h/AnDxT05N5H4M8pbvo45NYWU1pUFVHUa3EIfKIn2x
7aDmnB8vLiJYdOwHMvrE/+N2XBLPMmnZuI/d9v1R+PI1a5cRV550F887zyLqlDgd6pduBD+1Ognc
xrHLof9b9ehpZLpeZozSyrb14lEEsoxPTPMJ3RnpZRV9WQ3pJ3yhAIpUyzbOfQTPEKouXFwfw0xK
cZx9OaLT6HtBQrpOwhkMlpfOlji1I2mtYXGpPYYmfBu2Q7EYURGpUK5wrjLd5Am5O3vA2mH1Y8jJ
BRAoIy8Z04bohdSxEB4gprUQMCUGNVaSH8kWoxYlvoLm+w89Zj4IFT463KjKuEu9yjpMU3/erLo3
Pre4iC4nJpM05QRtqDcKZBKHTdpyYMhLyDzcviiUg8E2o5t2WvtRzGoSOrX7R7XaoLvSBdiFUwSj
zVwlu/BmAIs8g80zYFMsaTrZT9XXuAm11IWAmg9hVgdjiD9l3pJyXVWAVq7LfKWfj8duflMCqGpM
J9ZNFqUfZELpWDDBk2wF7MdA7j7S7CN+9MSPBgmXYZRpXQ2shhXrBixV0u+7+8iglmfNd6eVHSrZ
9o1tLDgfis3NAP8NnKn8XZjuLpO+oL8W+CD4Orw+W3HhhcP9lmlOEpFeKugMKkvDjxDsWGwgWfWk
kZtlO0A9EC0wsyuwK683m2LCkW5GNDJl88MlxIRRbtkxlukVbkYfm78mSmKtnGHv15kqXi/7qkqY
oFiziO/z8XR1FWD4g6HAJv/D+sAbH8ppOuamqeXqaxT7HRIOcAYWwEevGY2qaZCgKV8zB6Mu8GQ/
pvtuzrZEXwSStis261vURPbQnBLFH8r3dGiJhhDZukOkvFNa0t89uGB1HTZ0I02H3iNOYJ6qGf3G
8fTzpB0JDsVCdOs2j7t4rVNkiJGJHaSFdlVeeUNYrkQLvrzJTbnpqI7V1gAGGWJAmV8uEtjONUrY
D1AL0j7DydEoF16ZoB2+sod6vDfTi+cDV1N7tbnFVl/SNdO4BWyMJdhsbv6WgnOtODS9f+9m1rSJ
wRi84IuRfza+MnYdab0+Rj9gK+IGhndqC2L+coH4uoZ8Qkgw5nIfC00tlXg+FKaNksjxZrCd/fyX
Vb6WRKBFlaOaw7YZVuoy6sQeHXMLBUWPgq9C4yXs+AOObOLGomrYXFXMVY9mMLOu7UY5lbRrN1z3
95Ligyb0JOgk1gnFQYcaXqeuV9CTiKczrTEJA7ms8uF8K3yL7LJnCY9SPc7NUnfLtIVbUGuVi/Eh
YkePNzKLdmUv4yw1DYBGolT1wzrnPryXsvG93Bjw16lszsnP5PmzUBwaRm9C7CCkXEwpyWqqqvXb
pc0gEZKF00zIiYbHXddir7n8yooxL/BawZxqRrYWsAa8NixEsHqw/umhMFkAE1BquMO3p5Vm+Yy9
naxIZU+3q7GXwRZGZiGkGYUmiNzgDKPUArfr4KJGsWZluKeoDkzvX9ZNWhyaBf/IvYIIJovCA5iD
W9rJxgV6/IOuQIkR+FqW1eH4rbXj6F1bsjiu7qPynV0m+w+3SuzoYvC2zNMcCG33xK/kpVgm7X0I
LccGykAxTsGFZq4h2HJHYpLZJ8bV5+vWOpMUnsHOkWWcgqB3uNGdbzWmv8rzf66H/WtlPPJje7J5
C/Bs/7mXABfWQumuFnfkZik5QIoQaF+S/n0ymW+vMkvPymORVQ8DPGy8QlOtcFP62lBvJH8MXpqj
WQbb0e1sY03nBFXEXb9dBVCI9pD3aswTiX68R1LSc9ceS8RCq0Y5GEdQwO29guUJHKHKFXQNcBH4
Hvm7xhUJVxq2Y851vxrA8loUpR/+8fXL1gVgm0uad57sDm6SpIfSXVUH9lZwbipW7rM2jcgh6jhX
pRcw8hPnlgCk2XmT+tqo6HxPxBvYqCYYVWtmNfsOmz4O1cPqM0klRqDgbgGeecWQXrxbEwCj6MfZ
K1yjNVW0xOlm4bwkqFB7D9xZMlxbqaZusJTppP5DXwInQdaU7TCY4VQxd01f7CLcbRm0NJ6XDo9d
GcqcyUS2e7GQ5o7wEzLUzXu72OvEmmaP+avLXi1dWu5Mwr6pUgYa91r7JhhYTOBROrLJ9RIdIKoB
NkIRAF8BY7ecYJZ7SyGKDO3e+H28Vrk8Mw64ei8328/FYK+DSoQFFmzgZRc0pmTrk0VScM4oAuL7
ntkNLNZhF00pr0Nrdp7DhW9MwiuP3I5be5m5AEjk8syFHeYBaJCH7LIKp3SQzPf3C8zjT+pQOHq0
I7QJXE2HS/CM71VGclaUubttHSvhEXO3gH2dSNMtXBNU4VEEiwxNZRANTdbMYD2PDwcGlT4GjQUk
8Sdlt/wyxPWNgrTki1YcQ2TTbMBrL0JfM/J+okBSt9xQEGj+EwnaC/naWO+GkMvsvmcfcu0ofU4i
NxsA4fA0xc6D3B08TY3n3kG5bH+4+/ovtLrXMm6ucReUFxk2RpJ+vfcKekEhIGLxvEbWLve2m1T9
rXlTwJ15M8HsQKzD+WGAoue258M0+P+9tM1wFYjRYDdi6MF7WlsYPXedpRALpdq2yLKhWYAy6t9c
p7PfHhv3oEDfXmrS9rFhNedcj1Rn8kAYfz/kG2whJyp6+Wb/bwiraRw4goxTXi5BpN3iONH3SKea
qCtLisUINIDTeJgeFr7ecSsgjtdNP2P/4XlR+/BgSBTS1ch32DNN1D+jfY80XNyWDvHc8SMKIYO+
hqTFVywdnbt3CFVON2pM3uFtWWhrp+ZVVvEwBN7GbKKsMoKM4OQK8BzCW4toNd2RYNKarG/Pxc/t
1Ou4+mCCQ1WrzHS0S2t6mEuRtmZqT95RwX43veW2kdUvQgK1KuaAWnAJ5u8gn3Wv7w5MQ6BN9Vqh
W8h0QA4pZ+mF59Q2fbhghncHoJilDE0aKS9P+fyvF6P4SZpWYmYOZPBLFd7mLcJ3Ms0EESechcNU
KPvAyHEOUJBwQFYOnhi5A84VFiDVoEAdzNkDVfdWHT2cbGxnyYV3sAmSEnn2FOiNzlbyyc3+2dgZ
kcUw7CiN4CS2wOa9fCPHiWlSptfSmNJGHc0dFU8azhDURKw5buB39VOvhPdFoyuIZ6TBbU8cKoRK
bIYrJcfsJGnsfl7sPLty4StWl7mpo5KZeiTO/eDfMNtfO+3J+TmzY4en/R+vX2XdxJJrJa0exXN+
8XhH0Bn/Yitb06Y29rfMGvIGEXLd7NlJEVyz9kVJAAf/2M7a/wY68b7fXBCyokcMvzdzl3ISbcbA
CaFRxeXK9b75E9CvvyWEbRywiXzLULYV00pP0ZAQLbABo0vAHDD/4FUiNXjAbHqgrXN+V7ApHYHR
Oe9Y/TeXVcPzV2AuWRJS3gP7PfuZ42/PfwOtNY/c3CMxGUWIKDBOlVFeTT0sEf+W4uYmr8fjZZBW
z1YTL7ULsyXqVAwX5i5vOL8p54ehK/jP3IpP2yCS8XcjRO7bx2YCVTJ04XrF83ZNXyqrqqp45j0D
luc9+TcmQk2i4vUihnMoyTXO+bsKulxruekNvYgsJzwtWXRSpjtIni34qaQhGnOqHuDLUKoaQ0x5
MfxGZIcFHzCFvR31Yn8D5BjeQOp8yJ64TybC9YrCeMX7N8QB0463rvVqifduMXD2X2dj1RO5fafr
zT+RXH1Sr9RZR9mpFlCw2d6GbdVloAjFuZiXw/f2y3e6JSIpfjqiQwU3wKYsOnVE+LOpzkvvZOvq
WrMduLG8j7eRpeUk1NrwB8yhcOMmeFySG/wRg/61QbmrAPj4JZ0jRGeIr/8MRByVB91Df9M4BHdj
eGBIc0AIEIUzD8wGIgGpCGMcH63yLk6YtzY4sPWpXJ8rdDM++iG/DPRUEcAK6nxq9W4PecgrIdK0
UawVQVt60vTzaugr6Jb2Q60MtGiIlk5B7dwsfyCD6TnaUr/TX482Jm8GAOFgShLeJmEIKtx/3wEh
rU2wnNl3FPhfs+gE2w9dslyP6tCawmihaoLO9llLrihjrsxegI65yNZzDl+jF561LQNovLSIgSg8
bUDKdq/kt6D5VdJf2YITN0s8bsU2nwj56vK3HrmTxn+D/jT/bc3AbGuMoZSRXtDZr9DUXGZjxBTb
7VahzeH3OxmZLK6igGx7fd4doPi3RmXGxIARTS5InR59R2Cnap2m5qN+xyl5BOHsknwY4SOvcS0x
Jca1o8ZgE85h2EzmKoRP3uiLi+UFFPf1M1KwadCd20y/+BE0kTfnttdiuh3LWO17tuMUUO8douIe
PCN3K1UmOZnaj4U62LZjEX3P/YOFrUlmN/Alm8ja/pfVicued32IZso7uu0WkHoejPSnUk3Uw/jI
C2JNc3mRnMcCadLbUKezpWIbZ56iAubEtwxDPEMpkF2Qf7rJi8gu33PXbeZmo8C0PWsFpwdDS9tc
nubFmnCU7CQLQn/3143yvBbtJFcuhvU33LvZK9bAXWrt09FthOgS/IbodqvtY+ZG0rGoV9fgTnX6
Djz5Wj+ctig8PiJz3irU4UR2Lvq1UVMwlO/P71SBa3QK0eeMtNS1syRYvYzb81NN8AMjPSYidmWK
6nOkkYB7p6+qsWZe7CU5xYlRGFrNVH3nOFAmayDqepdK6hCpK0qbCZVo5DJd2Ojet6YIL5hNkCCL
95WEPTG1/qfcTgyP5JXoFOMu3h72oIrv9mA0XsaQjBVHtMDmvWQo2nyQWHVObAyWhGtNNAtDfAYc
QgHxFGzqpmDMnmxEkbhxPdFArsP3GW8w4FrAovmn5kuPVaroA/6TlVDR57mBGkL3UD8OXH+D9bpq
FMPLM0rZs8fIM/SUWUQswUHoYkQp3/uKF+S4uV8eD9cc6FM3ixAbbUgmZP5dNto4JeWS4kak8Yn3
uXo5iCZ/muKBoiKyZguM959EOmaJzjBECoNn+e+By7lrmd/PyuQ63FYE5FPlPfGqxYtS6TgZ0ikg
2GKPVE20sLIlufSGjGtQNvMwTPF1p60Dh3mz+iodR34YFzGNcryd6/0tOjGl70vUDJebC3r0zIHg
V1JGadzmAI4jtjWI1KeQggRl99gblzf27+pbBw0fgEMlSXK8Bx3MC9eADHd5xFIFhpGYUXBeCnPh
PUMuzDELyDzecLI6md0AU1d2neEXlnZvHP++H3myla/pNd8KmaA7PqkEZmJeCjDfoGrC4Rmvsa4c
+cXo/AJ2yhjARHKr2N4863CD2QBVgqCYgAJyfFHSfPmTDM7AUMzzIOTW5w+4u+IARyrDWfki35NJ
KQrlh723NmgNivBOMJogD8mZ04XRpld4EPwfaaHSOvI/nCmqSULbGcIjSjf8Z2SRxFsMW43lqm3W
/+VA3FvFForIDZriyxmWuxccIOZW1Naqa0Wp3XDXdUQAMh1w74jOb/W7fEv6KykoQds1spuhTNLm
cH54MG7YSfacVnYHCrxwPL2ZByvly1ezGNb+0PT4H1DMlzh9C2XudrLxJEnVtzzdwqFsKoKqFaua
h4eGtWHEgK+qQVlUO8a0En7JDnKfOSXEZIEAYFC9Y3Gaqyl+HzpYluMM55gjb8AMWw67XuDwwDbX
S2yw88WCZiVOxH6v26ZFHZx71VV27J3N1v006h3Tqp7Wq8HgyZt3H6zmx4vv+FNBODbAN5zJiNwA
J1TbiQI0hSyVsLvrWFafGwpv3+e+rld884lFmLoMU7YfV6GEvQI6y80J8aQUr1G/F3n8w1Dlv7tQ
v1MOybdWz9AF08pO8v6eLJsdd425lzVLDyH1BtqI+nRZEq22c0XllmU7IXFA8ja/OcbAtvsSnZlz
AZRa5tQHDsPIrIlfDouNMW60c42gpnDDCO754w6RdMmB6uJlpTDpW5TD/wn/yKfMdr0XBgpfq/76
2TbG7pmHeukOpT8gM4JKxXTQ6rln8CK445zgOyoAsxWa82hVF3KYyie4vm7oxx0LySaqDI5enp92
D/zRksrVsOrDG5pxF5IRHafaDma4dfHs1awpM4A/MCgMOrNelqIwkBaX9Xj9CAw+dnR4OzDdeV7F
IAU0+B0MYoTDpXjTEFBMSsvVo2C/7vUXj9zg43iLQeNaNqHdddYk+3jnLrnDLQb5HTfnDIPa/W1P
MVGfourNx1L0UFedTSjlIG/VQ8vfnqSma+v19nnbI1NLRvx1k5Hc8l9qi6NoGExvwAT4MQxQLdq1
dqpACR9u73e9vuhsElAvdw8aZOb0zscQiDowKGecQN1eDEixebVI+ZjlxDpIfHaIH6Kfy0JCOPhX
GAtMJ71HRQ9ThH7gWoT+vd/Wxwl8nMCd0iZN0KBBiALOEH6abAAJQQUH1IW/CfoW6gdygU7N6uTB
VjnLMK7cbXva4DPtZ50sVHLyotRZnSL+sXAkYdMvCDJ7yUTBLbhzWtA3LrsofSmUxvO5FkQoDn22
vCvUFZ2FHcBBj9oNR0RU+GTVzNcGv11wToB1EsGjoY37sjyBh/bp8we0DfgV+AzHcCn+acxqMNCV
6JK+Us8COr17k4dq0orGOhRmppmIRvDFHkJ0ahL3Sk2eP8wuJ0pI3Qvfl40AaDBEeBeh/0Q/l3Ff
6IYE6iv8tBr+YUVPPS19zFJBxZIFks3vuVPCAqUXTcZrqql9mNZYcwGw7xFT798MMeJ+WezZDlc8
m2mkR869xY9kqK4KbHLMKSwUptLUxop4ZiNcA9ebBwurS+H3ZmjdDmcPWSbkofTxnSlLmClFhaCU
8QJWJ+Bv7SdB/17S/X+BGuR/crLF/eHNhWe41pHPjk4KfREMS2Icxuxyz9cE9gAJ2Z+xu9uD8mMo
pCHrZ9xeuNDifXMFDmhWQZ+YBApXab6QUAz629VtRCKX0WVR92OMsjOHx31NQoHJtJEPOY+5saUT
uOy3xF0xlaFkeJKr9EYSvwxvm+hEeC3XphkPSiQmVTDCKS36YvWi4P9D18IOWGl+5P8C8Cde+gMs
H6cnQ3FrmCAdq4TbzFTgpP29i+u79jI/9Ll8SskyWxmuLiWOEIjrWn+Z0aCK+mZeoO1/Og1BWgTg
ahOIYWNHTLf7Hg3398gY2GEhlfeemVnSZ9GnPAyHrh0QGfY5IIL78ULtBgBfH3d2hoajTHeRp7Ct
osRV+7vi5lg5UF7LUtK6Hhmgew+Sw9Veq/Mbe9i10VgZkrPjvlwsg4S/c0jifogwJ9TSVoDrYF36
oAL1CpRed7TnERdMl35DB8UVLZQfu4l9xtytAYs7NK9LKtYy8tdR+g9Rr2sltKPVEb0YGvuG6RFn
5I2nen43TGyiIV6XQsi79dL1kVPD/4li/i3JEkhgXnc1A7GrVNg2YyuSN6m+nqDE0cqycpg0zBQe
DPjXMoogZ7Z+XcXjN1GaZDB2d/Pk5J/KI7o0t7zhbZI4woT+AcMDaEkixI/Qelq73jOGx2JH86QC
KQBU0ovLss2XXuiBzhsZB5Z2NAMESgQDJI5aSD0FZfL5ORCXITVGVjP3Cm1n6HPmO3RERD64UDpv
MK6ozWgGqzTD9UjSXUGAZydcICaaMcJXlrWtlud/Y/e3cCL8tNDMNwfDyH48iYOvBO/xsPf2E+YD
g2AarhUzoceRQtnfTGRpNHYL+DNQa+Kb8QZeAXwIa718+F5MxoEo2lIHDyL79wPr+V0rQZOABFEq
HBZNaAcULeUtomT1c8rC5uShbM3i4PXX38Yww6yam9S8pnUp2b1UcpWd5OEcs48GMoTAD2Pxtk6s
CufET0p2Av8MdM6Hy0ZSq8ay7KNeNHzujPE0RknY/d0T0KpV/51J+cv+pGyCBO8IKZHUKM5Mcv9x
9q7Ebi4UhZBddGgtHsL8mjvZPbQ/bZjEp9k3Zqmd/1gyHBeBxWkWEn/bPKZ52diu6vIdGH5vlwb6
aWoVlMfCXfah+6W1JYdtA65uQpsr0/od8U++8BhnOuovINbaVaY9D9zYLoePZ0L5eOKPkv8Dap0z
pWFij4sAbh4TTZgnNGF2JEP2/T39mSwqyJnXZAQqVZzYq8+Tpv86YBlTHgQ5Zr5x2CSIETV1rUEV
k5tJxxV0X6iX5prIuYslCTRAfbF2X0s5tOKCbUHQ04eENuyK5V546wXqprqCTFkx9phgXcP4k3N+
VOuNUGoUCwsUwzZYTG9oZ0+p6v7PTtmIRUJj6epLYDekpfDqmg3q2mFuNoyAum9f75aww45DlGHO
Fm/grO6vjlFOF9jh56QARNNzZgrGT0ygTetzdDO924b07J6rA0sjAhen6/Qq7QN9kdL3k/73HRiP
CQKRk2CNTLkvjnM/xmxm5HFwAWuc92thjO6aChQMU4i1lhsXqoW9Ity0CiyPjGxcRWgS3Vf+fTiD
ZGNNqJxL0Gwg7wuEolNYB1RIwYmADsMBBSUFl6sK870DIL+qnZ2gqW7ZeHKxM+rbbPQQxtNyIB9G
gMGpydkkZ2UAnvza7+/yrAZ4Eq/eTPAn9u+fPNQMHZIHbVZy14sdjAK7jBnPryzbqwQgcyujnOww
8IK11RLmF0HVk207u4nnd0A+Qxnrd7XHV59Iv8mo4xHg7AwE+3g2QKmALgOsDtPyz8hCdBxHkXkf
FrCUnTMou5r5zPU2vdGnNYssH2WNXJXFN71S6B4hLBBEPHb405If9xelD3ufXpqa7OtGzh3p8sm1
XfVVAqjrO22X1sBFHTRSGLUtQFF/qYVIhi3t7TD+yIfHPNv3wIBqx9rhrCFGIB2mF1Upu8CfY3fN
Hwvn6JgZ7s2cLBvPZdfpfqG8F9S1jiq6A0TGAk4bBCQXVO7W3rv9NTh0d3kGzP/qV6mI5ds9/ej2
uUvuGOhNXZRjjAe6URArBWRnpktr+L3q9PJy6lAV2sohHWj3dQmQzYKl1WOEnSD/ht0PNIueP198
QvWTqvx11NRkLOiB+NzDga3LQ2+kglCCDLXOpoPOkWshU3VZneSANPzc5dA64n2oAnyj15IA+x9F
knu2jeiIggSfy1xST77WBafEdXhwpRe2SwIPeu2S8tHHbDdwbKZUQ7j4DAqfg4E1cxOkZLkcY2bl
VuomMdTam7DYZJ3XsAaNsPa9tpsT8r9BxuGhO4cNc2Eq0zhrzK8xtguAznEfi0aDBAsQh49PVL+j
eS5+r51rldHlCNH1wxgyrJ6+38uJyhG/Jhx1lJbV0WYpDmWw5+R7J9CU3pGbe0cUCQnM6eLSJFd0
bRLPtg/J5G0f2YP7uNGdHUR7+p1DAR4ZKG6zKira6h8HdM34AiWjlNNYzQuuv0/TSu7415OsHZzG
kV7yDgUZv4ZtWHsC/lwlK9IZI3c213/VxUkvSXNzi3g0ndX1X0DeW9PnNpahqZZu0DQaGPwBFVSq
k1mHIgVR63VpBN2/rgJ81n6jDTNs3Ldwl+zellPmDa/ZkT/asnnFK5Ns8Bl1uM2aXmelB7n/dx2C
VXCsQK7+ty0bUIBBaWrHnLv6PdqaUNrhdWmE3juntGsFpH4pJ1XgDGwi9mxSEEPrH9wb7EL7aG4H
m0jOn73GlrgPJVjCj4WfO121DlQUuVghciWXk/KKB8HUtYgPu2hBASXWgzCLdyQJbedervUCddfx
1dO6NykqELuh3ef3j4mv9vxAeCjIUUJfB3DsPRreL+B1Ah/amHbrzVBoRTEPKhdEGcXKWu/9gy+X
Mb2Gfvw0/D7PdKa68YzBuj6H8h39B6fHm8lI+xCn8+5Vgy5DXw3H/5tuPEX1mAb3q/RDT8WQT3OM
5jNMyK0vT2l44Iqj9RGCq5bGd1yMp1Q8PxfiQ+p6yU3uILpWfmMlgapsqVFKW806SlTEPlXOiNTd
Gdz0p++ML/a77rirS1cSIpndZQsmxyamZTsHpj1blA8RpGmefN6B6DmoAwxbIgD1WXK+hwh9UOqE
mzPYwSRATfaUHyJaVz80ET9wZy9Y7lyEVIuRmzlv4EH3nDpS/Cqgk78KDwVsMs0SlkWF5h0sTh+2
k6w2wuhHq/WYgfm2GBLbXOhtkCbFxEuWGBrXVdKueeQCn6Vb09qgY7/llZcFuuwyHtC/civ7VjjA
LwAJWTtzq1Ui2DVWadDAjiMWXV8NNLFpbcXwGLoaf+tDN9G8FPSGHnFoI7y4+sgV/vbvBfwdNqc/
VoSehwdlXhB/RdNjMvZYNsm5EGtm2DannyYPMt8LUKBjUEIrlD5ClTX4sJxXiwRUs/Y+VZgl5r/p
1eylOfr8CRjlxq+QFi3bWh6iTOlE1lQ8Nzb8lGp605Bc1fMGzj6VJTVn/rRLiXHwD/1AxN1+/rHo
0vNqw1L5G/jQPrWDi7i2jUdH1bIvEQ7rwpgbtXCYWNuoIj3yHAxioGPQPlMtnn0oIm+D6IV2BOPP
709vHZz5V2FEV0wa3zAZ6QpYNgXGn4f6ArNtekkjGRfTtrQ0FRL1nVo6ibnY1AcIOiWd2kgMsFrz
rlLsx/ehWJxGrVblBA+A8blY+aTg2/vPyHz/BCrfqWzl/2YdIRrNtmxK7ZqT0puzqoIqQMTbwQzS
7woCPkUNEdQmLiSuaFsACGYdQt2u6XKUuvE3tKDVsByECPIBUXDAntFhofNRraDbV70aLHTdxcuW
rTiw2HQ6hGZvA7Z5rMf6WyKcHJH0Tv75Vnsp7O6T6ix4IHlidjr8La3I8IuOl9NgcKUV3uClCn9G
2mea39rVDV+V0fq0ei//BAKWh0D6tpXvo60nJmI1y1rpVoUREwTOARkuvg+O7ZQvFXV4iS/QeXZP
2fddzTa0j8cEqUipd9qgr4rTMjZQ4aD33dP+f4wOtUJxMLqrpNa7UE0jECGG4yAsNgCfDD4MQpUW
g3Z5BsHgz6Bxs5N7yjRLOQANbFj5utrmhSdTcPKpoJPHBFX75wmplJNTGvBKUw3WMqze3jOfdYNi
IBa4SraZtJIC52sQD/S3bGP+A3GONex3ZURsiIYJD8gDG4AZpCdJXz4e9gwUaGBem7tyGCHySnZJ
NWzzc+ptJAesPBp1piGs9QwMqCQv3Wm/PQjxTrjBcMyPZjP1EheDo2UtbYFWkXHgElGCP6oVgb7N
mELqJ643MWT7sBLUgiAY0ufoqLOVbOoML1og7z78Q69xKMS4plM1WnbSMiDWSOFTQOXZr1aXnROv
fxDdULTt3sHKrXTen9Y0bZhgiw+5zrcxTPGyubHVkq/GjEWElcpDk+M2gKhDTX2tAs/kzPPdL4I9
yJY1rDd9otyv9+HLVWFhxt+Qex+a63uutKznzUl9DtNvEWFAGqMbqu60F7W08WaaocKh9Zt4pi/M
LwsDhir+XqfH0LWnyDdIITquAAUp/5oUO8FrhVYY2VbDcAXPR7CUGcX+4Yl6CmpgccjsQHaG+9qL
U2ED5sysIGH5GmRg8cTgE/vI4xAzw994sQDkmlMPH/GfimMyUgo51R47z3JvLOmkBQsWC03SGkMo
YFfdv9/Fjz7/J37LfUwkih6Vsugdlt0f3Ov88IrIQyRhXjHfFGLIXrrM4S/pBk0yBEK5UUlS9O/E
5UZkDzGR70/qoV43YtgkgNdOnijzNUe7QKdaUvTIi7/zlwSx1iwDuryQNs+nBi1T5cvQAUhuK1WK
oeFZc/1jVndHFJZqfIuJyOgWJRJIGbOyWRGhtkfymjgfrNJIENq/+uhjujX4R67zyQfP19Ijh+4U
Ye3OjsuTkt8+rQd2+NTzTF0XYJVwtW/6U+QPK1bzE6XmSeb8KWKWqVwf6RHJjsysFacqCDIBeCQ1
MSakLZRt7GdNWrv30bzxu+5EtaKlwSbnpWfnLDEPfL5fOib2+yYR0SPoug8DexfEGziS6jaXh48E
lmOEnkoBg985lGWRqJElWjbiGFr04I8/s7fOjRLlmqURiglLP9OCk8ki6VgieQVs+88T9XE01h/r
HluoOfUIvvJGuP/eAu54x9WuhkvavHXnXdsMiv0Das2cR8N1dP+fNutygncuuCWHcCA2YpxfLBzT
V1httQZVoalEkr+HnKsrTvlKSl0diWR+1sRM0gHqhxCSQmsoTjcw+AT5dAo3gzaVnv+OGksqyCqR
OwO7C6EMtYerAfYqTzH8z4m5NIz5EaP82ukJacI5nVG+n8aboiIwAppWOf9uAvzHiWdI3lUj0tID
N46hzsvVazstvMdCZ1A/72RDvzM9XQJti9rLGjL054SZRiz5G313ZMwNdGJNEWtjNB5/S3vuRIyt
HFUpujyAQpZOycLdw94Uz/Hle1ASWFOfBJQmNFDU7IcmCZluYuQJ44L4FeqhdczhsHT5YVAXHQX6
Rvk85o9J/5AVTc++fenpRrd3aMjRmUECLG6A84Kd/A9LxV1Dmb0E0mrusF8X2sucQJdcLRaLbkaW
zyMOJlxVzS74aXhO8rYlMl6RKqfV2ZFMLzFQQ3grYynIKR+skBiRyfsUa8DGko29LWRNNlgf+PR6
Pxto/6qc6t23J9e+IYKKHT4RbsWvpNSA7WALAJOdTjWvs53AzNF6kGSry+7M1DJvNIxq+67RfWrM
IjEmAnaHh1PMGTpPpODZ90IMS9kLEsNhzGoSi+TaLaLe13w0eo7bdjn2HV/qfYSCj5ASc9H2xbnY
DtJBXn8/4ZgzIH++vgSr7DZSlZ8Z7olMIOdzFlecFr3obx6ZtCClFIcq28bctMMQTMYASzHm+ouy
bQ7ELZ5xU9XMd1SbTwaKSD/ukcjdnLbTrOwomjKjxgXdbmmWTPxi2cRJEoYPrnvy+4qlYkUoptZH
RpJDzP62Mq3IJSO43aevDIIGwBOOlWZ8Zx/GmZE88T/DHf+TpL8Y2mCyBsZeA986hwVYc5+ddN/X
K5sdrSaNn9+yzPlshdoXUBvjtSJlkFJBDSVc2KKM2lMgJkgYt4RGrJg1+AzCBmK4f1D5kBRoVsEW
3T8SmGskv14FIyznOhGHvQPI3pRxcsR4OaonIxaYdYlDZbVc/s2RawiB+wd8Tl9Uzyb9W/3qjgr1
wBfK/ARsdoGKlvQMt6WZPwfe74Jhm7VlrPTX6bPMFh9S1AMrvHHU2rBAj0DLE0DEqX2bmI0jkj8N
ML7ecK17SjRFo+J5qeOSfCqhyPYtZXXUmDBINGsWW13rXz2ckbCeh2sVLOQSCDVd2Qhj7+p9C2Iz
Dod/chf9lyFCPmPYdAgr5dBwo4JMmgyxbUBRauhRKzrhywk3WjvicpGsRW41Bh6ZgWC1PoGhFzBF
z+AkPcnTcPCLewnlx5n97lgdHVCnV+5tXMWnQb5jVztxkCTbq7gbpcgQzm5VEOGC2ZunhhLIGbRQ
r07XDR/vMd9H1Vv6sirfsYqVt9e0UuuCzcjYdAioTxgTcwiLm/rkfUfNFyLoWQUV8+sVRt4CZuOA
nC6SxZr0wmLcuibGbvslwh4CA9jEVvlh8iy0bR+XWVSFDBBBMT9pcIRXmKSevPac7pnP9tdPi9aD
O6OZKyy6SQAQTGfVhkTbWQ/gCJIaFzA3kn7rpLUfvfTTyCzBPZ+FL9t29EAy29nGQzJttgdheDVy
wGjGZ9GMzJKLgmx7sC6TNC1YCcPBIat5RiGwUaB45BQDE0HGFQEJVe/zcr+W2jRMapVwogjCRcgb
Rw2MYmNlz8HuqFB24CBoNbj/kawHNioFNkPef5ZeamJmVZqKNqAotLxfuuONMpVAIW+HQogMhIDO
VITrGggQR55EDXaxbvEc/NiHIi6YDoOErlV3J8OWLgiq6OzBqPzTGIcd1PAv/baNdRmaAo4s45Re
m1iUVy2iWJflvSZdkztOcmZB1gXv1MdG2QR3qOrjum03ia5WDr29bpV8XRQ8kB7BZucbO0dsskCi
OIJRMM7PKLAiRxLX6+ZYfnB1MJemHs1CoKs+N5dIzCHaiMMwd+sXL46Xavy3tB1xn2ZSd3iwXgLU
q/F1u9LQ8uuqSyw/JUj/PZHHZd6RcR70eFdBdHGkvP+3nz7jQcV8oGg5XQAPnamchT9B1m7JXiMU
MS6RFL7qVtJ9GIKoYlc/G3Km2fO/9hY2tOY+6tV+0TVbL/ooaC4aKY7DqcaUVfTP6w8+7HC92Ww4
j0x7wZr8a3pvkDZr0dudPQKO+Im/di73nAX0AkKOhN705sZKof6N7RNXerO/9tdfR8nzEoKMMdAW
4vEO/JZQJ4eLmrrqzl5Ls7P797kYZMGv9GIiu83hvE6S9yOnCRVqSK+wrhRINnwYU/j1UTOI+y3O
eACbnHzg2swQ8hD4zLMORTYX7MMniiW2Y+9CapSe8r873w6EaJT0BSJFiSecvi62dQKX0V1OD9io
vCBzpD2cW8RIbhnLuwRy1zsSZ2weYDlecBwCvEvQC8FolS083QWA/zW5nh0BlDKSpxC6LxK0z0qP
JpgmcjAfzByt2xw5+pYpxDQDD11VTEGZHXJEBZpanEA3h4qeHxLyV/Nm+mVOCTk6HxTvnspDXENi
KrgoKVIjcH3caF5zB/GB7saWa2qwuxoNzCRMGNdQkHW+wBCs0lCaf1zv3j/1tJ5MIYuU3VhlMPEs
KqhRfIg+7RHfiP1UQMhiHqykg4RQfgnlY6mhVaW1um72YhrBzdQbusq/FpDn07APU8idWVkKWQc3
WI9kVZKW1pQcKTyv/KN5lssa7EEwjfaUDCsM6crcQz6JBYp3W2RU6u3PyjEbmiGX/Ei15BjUugG+
Y6f511H9UZyyiMwye8UXkhpD2oXVC4GnRV34z7tuNEHguKPCQxSjBBYfu5HoZZud1KtWw5TEPMT/
ze0++UF95SgGfnSHJ2BUEHiUQqv4AUmGTr40Bkwxj8f5YigS5Glz5ihmy/zTEE0fy9NTA9KoNKVy
j0g+Roq0qFjCqq2Y7yB8peEnqg+deZ4pYmJK9urF2W1M/VWjnixlUFkwsHxDYtDV2fLwXtjXz/Xk
5TtWFKLBFtcDpo/EA6CuALCDuCffX8tpLBOdS8lWZ7ITHuN1mO7J5P5IOZegHo8zWOL5We2XOp2P
mof7HdaFIvyUwAsfSoU/3P1qz8CpBuz4A8jvHIMqBNWP01Ny27gppAyLQsawp0LIHxtC+uWGIvYy
C3V8ecSEGd6uAje8K3liHPf5EngEDHh2wX9H9VOB5uRULFlZ6P9Q2SpWYHVAq+fWzbQPIglPZou4
H1HyEEPGy3IdExzkN3BOESZYuTPWg0Ybqdq3yo7zeR9SO3oO1eUoFJtfXLxAsqFjQOCkbW3vberh
6BKzkjPMShsAdUF9ij0AoXQat4+c4hUEqMJmCb9OBdmhvrPodFlvA2zHgFjDeQmC4Xo5mUV/1Cal
WHUXzdv11Iak0hNJYvTKf3UqqLxOds+d9GW0qw+yp3d9b5zia7UVEbRGhDegDANyWxCtHE82R+Jr
tbKEnPkd4qL5TzVEDEzTYeh5MAPTlU5Y1KLBT87bFujZQnZsfC3vI4UekmGR8iGrpyIIYfcgYtZP
x7dEqJlRQAj0ShGhK25Y7Ix5Ar6/+JYx0aibUR5awDliIiXbK20Pj4uP23SXa+f6HlUlDd1cOoKj
5MwjOZf2EZUwO7NFexdorTD8We3B0DtWP4K32eyeXGTOW6W5GvIXHPJSPpLo/GgNt6J4ZuzPMw7n
HNjCDA932HNohpKyntBfttGke92IPVt38o5z/Jv0heHkH9WdhbY9DK2Lyk/hAVwZx2vVxKVSE+Ct
jfWSgCCI141xkx6xPyOY4fC40DlWy68WYFydDIp4/45L90DL6s2v1F6Jo47Hq9Op+zSBBVgHdpQ+
DBrgo1dapBHjon9TlrSJRo+d0x/Mjj92a5tufaY3obulLNT4tzPkfhzbf3GBan9W4XwEnUQh4Ag0
BEDA8bS439Jo3mRdHGrUh/RbS4PQaRX2+GeyOR66AdzOC9hrrlcy5w/PpEBHyo40YOpWWWLQefhV
nc+thda/FGazSDwDDlVd4mb+IdFjtEAsDQfvcO4Kl6pIVnvDUWc5OmVk6n6/4LGQD7E8nxKSYDjQ
rxuROFOEvUCFUj8q1Bbg7Jt5W4QFBne0Y/2akqM0AmYPkdVF86UPKUDM2PtJevRkAkfSRGiuZcnt
LFFI6SkBFdfqessDtu6MIYs2uJB79+4MjKjLqYk/NKG3dbvKcMn9VAcMrAnYd2BK2kAuvFMwU5En
Kaja4/6XQ+aX+sRWkzT098AhBI5eslvJ16ImekJUmH46esfmCFYS21QC8mEKFdypkonrtMnamYic
6Xmisj0klGWTkrCyVipJIZbha55g86a9m+RyynYcnfN9RfIVxnPyM4ms4/jXDKw2QJpSbDsQq7Cb
b7J7vZFxu6qyKazxFrG/T3zewvkBOdGj/kAhduiKYW9IAWR6M9Cj0klLZVQ+D7FY7SfAGClrc4bI
mQmxkt5KJ0rID+OBAzf1e5v8Swhi7WBUsSepBR8TZFaA7G3Dfs6nCJNjnMKClO0NsXJBnyILspoo
xUiDdxwaHIqWT/VptV7IIN7JeuWwxY0of8Z4P2p+NvHF4pNeYrh++uO7ZXIaELIcUKLCjC6kNtQI
ygLeA5Aga+L0zeGlwUiiNq64mNP+S0QPUrjE3MCKpihFoSX7PCrVQxMsrHJrlLBwBsX6Fn7UCfEj
bGwKA7fh0QzZCJEVz1dBvhO4Hd+gk+oZulaj4VhOrB5HRW6bT8CgxWoR1bjKzPloCG/n0610f1/v
fCiBZv/TfKv4JhovtIaM97K/sd73Sh9Zr/+deAjYoTR/5WHMjvLH+OxJsvdQnawsd1W+IzS91GDr
gyopQ+J10LUL+iUQSg4m+0zMOgrGWZSpr3ZktJz43gk9Kn6h/LQz6S5Eg8rzHqfzFEyQbfPIsvrH
363xMLTpXUIZ/jrkr+iDdbD6rCS9ppe0v6bZ3JNL8gphXdaWNDaeQMt5ksitzbP5J3TwYBwnrJ2P
4GF7ORkR+fK2k/X7rckmmbBwhIiY7U5lZESiiUCXt3ASkHYh/3NZLzJcXcwvOdeZz+ybCBFBBKbd
6Pb24n4SJCXIjr8kmVwgYISRIZlW19YEaAGsaxGSJisx3uWlh016TkSM/8gwc8wZV0QvBC3jgsjI
zB9svY5+RgigyyXun0T5jPeUF9o00gpghuE8/10lqJp+8fP77+Pv++OhCcykNGkE0yreVZfExHfX
FHvuYjD94dbRr6kD0JcGM5Az6ZJ4CBFasZSqfWeFYp8gRNMn7MVNQM2XnkrVyZvFcGSNBXGKYpgM
eFul7dZKNzcLgq8lj241TcGbQ8oHC5AkD8Kl7FiVA0YpG286xXMxwdSXCGwwETmeUtggqBQRK8tW
bH0w4rrnf6yosCanicsX/HMHFuF8TDFnQqt4Hhg5op05rQlZH6zohoO/aTsdwc/wr7sqrYZ73TwH
VJSV0maA3jEKQMRGFl9nznO9zEAmO9PLNO2yi0+CEgCBhllShx0yvEj73rKqWV69HGdgI6ZTJjP2
dZRtd2e58oxbBOoRD5YyQ5YIqQWDOBgg8f8FzxLOxRrdvcieJTSyUMDdSbYifZrmOP/HrQQZuSZs
7bcJzkq8Y+Wz/Iks4qOg+XcZYZbiPyavQMdx7rBeLBJze+YNdjSkdLO0D7dplBF8u1Y9ZKLudpYR
ey04LG8nhx5N8Uac7WweCGX5cbVoYQnwIg58rOVzqLDA0mgs4XGj5l01HrM4ZiYI95jE1nt7rmvV
KQJs0VA4gqGTGNvRQw/d79hyV2AodKkenLFMbHiNPv/eHLZOjXHxpjCdtuXf5Z+NVhiuusbamMH2
biy9Afpl5HQdHceqpzjCnPYOp2SppjD/wZ9ZbDpFW/b2PSU/dxVNn64KBk3ZbEzQuP3Ci5br/7wb
xfENl4ddNqeuIspQLo3o3PJwVDoNSZXm9LMOD7+T4byL+g+ZqyS5xnUdrDZRSGoEqUxyMHoUIKSG
1LMhBPmTP30vfdUl66umQEVT0GkZqqm+Fq0ANOx0Mmm0eLoQHanwsp0D52F6wyg=
`protect end_protected
