`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
JKH/Y8PMm78dTPKgICJLm6WdnV6dYW6cyfdQ8x2rEf7AkCCiuFikjSiV6asLlN8ATK4hKKyy0XQe
A9g3Rlnm446X8Ng/erhNRIUX2pfdlU4DO7S1nh18yV8KyYwxiI4a9QljxpjKcBEyLVmyj9sVe/uL
J3VLCeOOQj5FN30cJjuUW2JjkD0kog7QgpUgBGjHe81/1CWYd7v2+EuxaGxMTTGmRBidSr7WFKR9
hSfDMpEezj5wINfycTYF4+ton4WyIjgBUXV2A2TP+VAhz3NoqXK76w6uoEeWzZqUZVX5WuhBoCFC
53/BIqzxm7Fghr9Fdyybs8MHG/Sf+4KMSQZOYw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="2MMHbqPSz8lfY9BFYyDiTIdgn3TpDiXwcOp/wewLMwk="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26208)
`protect data_block
+5+6LNvVdqu4UZWx0CtwBEOqBJVIHWi6X9YPLBZF9peM0+ZtZxEj+lj/me15dJHw3Z0Inkr4UTqM
9TgoAFa5v49NiffcLVwXQWdo7RDE+UbqkTumLl1fUCJx7QdQyRmasXAkUUnqygk995bF35ahHmkY
88DBf1vXckUoin16Sl29lGu0pms4eN7NnoTG1XfzqqLMNNitATmMHyj/HZy8iUjfKICmq8s3UnU0
tB7LeV6zkUzth8myBoypxDFfwJdnsOGyYHk1blgEEBbeP12V7W96VnR2MMqATQfaKa8uLz+2uAaU
Sgr8Pu5zeBaCcFRAgBOy1AI3m4VW0CoPSORYSwJcWnYuAqY+1v/KLL4Gb3b3jseA8PGqmt+mGhFB
K0WI7GaPJsfWglMlzuY0uGoeo3HUmDz8fkonOx42tMgetx9qDkt6iSh+vpq/XbcawB7PoEeLVDef
7mDnJ7I48hVV7qXMPTgT5OiCx1xW73Ea01cdXxEnKx9zeB35OnSH+tS9qhNStx3eW7jctw3rJzQc
2ciXg28EIc2wfw827kqM+48HI8jecOxVL0j521QCMiTj/NWD0DlzecP9sEoAcW+D3HVq/DQggSpX
W5rvSMoRgFyFWGHx7tLpSop5anGkOBnSnK/2OFOTdilFRz47prlMSoc1ibSPbT6Nca8s1rraA6uq
8hi9t7LQUzsV4USUZvP4xteqIP2g25q5ULzYuJVQlNVvQME7o3jk+Vt/jVbfERn+lQSEjOcx7Qxw
vnBY5uJyKRC/tjL7hOoMIGQe8f83YKebaO41NWOkBhrh5nFHOmVf/cqqRKMvPWd7GCbJ/r/HsYKE
G1M82RvYVcYMC6D4X55HpffIzaT5kJp3UQZJNhUU9iyn5eftIbNhl7LqPUlf5ZoR0CQ2MABauX54
qUOpPqw1KIONNLAkXzHeC/r3Vhff5BIvVpOlviRRCNyJ8rMUkVspYOl4Pq+u8odZlmdViCLr5Epp
iLkb6uKOT5+TpgbFXFLi0gNDTyKZa/GXsrreq+H10M2v1T+RzGU5TnOdoD7r6lnpp1UgrPinrPvN
u1bvni0Yw+1FzzlBvmc5HEAMc4OsoVz6tY+IOrmC8HGwyiEiMxZ8awizwLqodWpPHhcBmFsaSrVX
hEEpVQoR6MFNM/5Umct8o79C6PS9DPo/iX5Zqe9XGKZaYQrUjRs0lT31ML9qxhr6my6kZXAymCVA
IVmqm26oq8X94W3AgBa8cl9LXtcMNBUWhVRijVeIqkfOwQbsyc4GkPd5GufmXwn7Z7GONVEgPPkx
4k4iRePHyKIdRMte4IHfSbTwCxBf8jCHUFftTwDOLIR1j7Y5kVHvnQTdTnIvZBBX0d/WmC7cOcsK
45QFa00nsinKgOu1ODGU/FKIKT1j0gpU7Td/mIx+9WDSbUk7dZgF+Po61x6BEcWKNA8cfWx9IPvm
j8tTGAuPDZKRQkAfoWq9CQY5XkSu3GKTT04qPsb7AmsFMIWxgQRpfAYkPnUSYUA6GPIbUoJh6d6y
Xbmpt+g0AoVKIz0XkumERRHxzewiZdhAEdKHxoo7VaKuAZJ3oL5xq3kwt2iKop9Zn+sx+c5Qm8Tm
m6F0VqGqaYWnZ42nB1GjcfbyV1ELx9suOllZWyEvl58y+b0IGTjwPvyvqib8haFzKCZY2U++0OQB
AbxjxQQ4j8EA1yWAZMBTIaRuZNfkHXmSSD2GFHPGAsF/oGVMuVxVc+Ghexz2Ms7eCDP3kmkEPkm9
nu+33uYvoSVI0f1eRfIyoPMhOVG4EsUGPlJZAhX/VKsh2H8dKQGeJQjU6QmYnwMYBdkebnB1K3e1
wD72adkVZgPjSCDGzzvSLrXSx8qRMWyDzG4YxYxj07n5NlVDVjmsPopiZ0cNmeLDGVzW8w+xaWCF
wytNIJ7uwEGvVOii73GZVNjiqdAKNtv930/6vDqjxbD0Fn6a3AbkcGpja/qL02a/c2D98qlD2v07
L1IcEViq+nMZfsqoX6KyhW1i48YQGuE9RpVx7uYy2mjMxcAQor6/qSLs0nbkzO3xfHHahLnu0WEL
xKnmMXde8YzHcatJd2gwCPHelz/5seXQrzxFXpVmQWxUYRn0KyrbOo9Bm3xO0pXruL87kfgcklVf
znzpmm06DywrObt3SaSuctvlAmAWNPFlLb6ffeHmTFAcEv0eL9e66mT619DWhvv+Sbk/+xSXoJOG
c2j55e5c676BVYosBax8cZ7luW8DEWw0bhDZu0U303MLLVgPjfa025dF5Lsj5Y7UeTSug5cDjXq5
hnnYw/Hky/XD3Cw0EPC3enk28wWevQQPgk/JnxR4n26phMd9BSBmiQ5+D+FvrvBk+GgIuKhRGmA1
MxHBUs6R/eDjfS9oQwVIl8gRmH5VWevYnlnuOA7F1pqf6hDDpuYA1k/hWJP70haeZEacr/8OU0ZB
JLoQiKNxPS+pM2mS+FgAiDkQrs6sVKBU2jpo1ldExIMTa68tcJZ5Z4uCTwpJ4dhDijBd/8/AMRBn
QgzfWe22yQP/WOht12OGu5jO3qnJmEq4t1dpfHzpncghZkQ4hPlCnGIvboVG1myZbOXsxH8FuvM/
jUSp/1ZqjqosWOwXlCAvZIqTu+z72KUetca8q86fNNaolsjzNRLjtsO9lRNlIZp1BF6M/vH/P+re
2sAXmKDxgr5LKd0txYyphQJsvUaxFOPBmbP8PrExRIR/HEnUsc0Sv/Lsl8Gx9cbC1am7xu2OQ7ms
XmnDGrFMSJwVLeNm9FwvQ+5745cDsmgoCglXy80WhDHI7hAK/13tg5vJjz3FHYGos+XZDFgd3dGv
zbhEZu8xNWi+Ib53oy3dIVflhvR+RDTqwOivXRdFg0hSNej6QCWKMuOBM4ZPw7WQOSsSiQuKojLb
anPAJv5Bwn2qGSHyfeNSrci3rWvJwp61OGP0hIrckRBnLAbvMafNH+SipISl5dgFgsj4di2NwXVl
/b74bkRku1e9TeAPXjC4LPYjt1lBrg6VfzkkFr5twJDVq18osyLL4tZi8XS5oh2s+H6lwT/VjqNg
sf0gH+oWIj8qmdiJo6k4gz/XoRa5bd4XiuuJQCaTYtBAMvt2lAB7F5B3LLL3+PgdgLhnYZZCzyf4
WbL6mhbsNCi6OuFMg9tFGXdeSwOmw/iX/GC86t4txwuSNvRjOmBT7cf9sG+Jf/pPLAr9geGftw1z
mXcPfq/1kz30GH2e2Xlg3A34RBe6PDtYOiMHqra3r4BWN+nj6jYy1JNUFkVxT3lXXKlFPCYdAspA
3lYjdF/PljfUNpBYb/4fNbYhis4p8A/zi4ctbMMqtdHYAH+ukqhGvQ2B+lWvnE2d0XrOJY/WKJju
O3LKFQ3OrNf7194s0EPrFcZ8vfPvR6hVnXFbi0hNGXfISGLi94ZPDJpc5HFiK7KtHHCNJ0tixccI
xUqnbWxOTuU2ZQUjucPav8a6rIM5/69piBvCuRdE+3Fns+NQXvt4iSdL6VJXY2vdnEiIw+3AYXkP
QBJzCBt8HTdGN1EKkfwyAkO72ntlT6rukEU/8EktGCNGmw3oH4LqBssa2MMIFOn5M7H34T/MMk0s
tHqE8ucDcCUElaSZu9VsYktzEY2rWUz02kC6tA3rYV0GtEECsf4YOM/P6ZDdUYYQU4vuA26N20Fa
LT4tihypLv7K3+UbgyvPypXAjnqzvfQGmiMxt0Nubaq9F8vMCHzLGMvv+j6l7z4oq1H4HAaU2isv
Awu982kJUwz5FMpQwzesBeiydJv0D/bHjzhuVIAPBsEpWB+13/0rmTkWXzfCe30GogJRYNgJVJ4V
RZ3xZI5De3WjBv26pU7IPJAD8YcKI07X4MU+XpT2ZLA0DHHi/kFN6X0q314uMduc3Cwat0L2YGxu
cA7o0vMN1ODx0/UEa/MEwxd1AgQSCgOMv4VUu+9+w6cIUFbBa1L1LEksbbp8yf3ePdD2Fc+N26C/
InetejoS+SsM6VGdpKy6Xua7+CVjJ1h7WRsi9TxwYv9vFFLoxkfboJ+76MC4ttR1u4rqiersyiSY
ItXiS7hI0XnVNpbDt05BIlbhrE9oOvQuknDIlU0psN3cqigJpHutlMx9oovDhFE9o3uttOXh6LYf
/1Quedt0lXyRsHqKdfkpb5lLoWiMHXvi6plm6nZlYaqM2dAcpHSiVWx38NrjmSAjh31H4OOeSCwy
eYHwbxko6KFSWYfOzJQloo2A8vXayH7G/tvxbRXBPDc/dfWMlZ9v8dJgjo0+O2lNRytP0IOl14gc
aabVAnCHGgA43u9pVYvaynaJqhSHSSyOsVyzu1hnYU5qDjrXzn7j3p0atmAV1rWmJFEyLPUyQCVT
r4UQ9hMrRN9i9dYzUBLyNAK7HcjBvF8nmQNtFKd7XOvZCH1vX7+0vcl7SxeiH87cWxReaHveL1jz
4G3FcxOcCL/6sqH0OlramU8pQXf9wT+9lIJO4k2b15L1YESXustP4TK8Lo9/1Wru0jXT+RmLvW7C
430nBd1jkL8uZk0j2dayjQEYErDkAaV8T9DvjkucHWSJGTvE410UkgxwxVArDpVH1soe+HC+GX8O
ShWzJjh+wC2ZrtX0NisY1zcH+6QzDK9UHnEpcGBkg/rua/sDxZHs5HbZJrhdcF4gX3+HkmbLYz74
Jqg3lH5oV0tngnV2x3fwdkk/W1vyOUQEC/a1A19e1sIGCrUfK3cuYDXrr8Hmb1TCz6ATp1MqLDJQ
pnPM0wslNES9u3DA4ZPjRa9oGvrBiaoy0LEOvC42Epd0V8A7HfWkqpf6yJbjl4RrGDKDIRazJJDz
v7V81f0h8p/snSz2lz19ikAcM63QVgTNksSBl0J8gyaukx4oUIaoyXqdGckMF4USDaFMwuRuiqTY
Dbx0dp3lXKT3Ubdc4Y3Kc/ca9I/odRrn8a5XUUG3no6Zogs0U06tqwHYe4gKNvDPyG4xCxs8xXQv
NmX5pVzdgLBacWmkZGvVs47ME5Re0WOCU2U0VCnE8vtYuNnknBelxL1yVXFBCeGh99Ed/01VPKv/
hA8i9uGPSOh2LvN42pgY2rZGKvmJpeeVSYqqyaB7f7r4JPHb2Wu7cqMKnAvuiUuY20XtgZSkty2Z
qov1V+qhZbMqIs6keurnsPXgpQ+ztY/rHc+nT2WsGCUgC8skqXonYBHUDnsGnQl8+tgoOwHEgl42
FMbFQjLBaSB2/6KNKujJ6mLBBTDR6KOZuILBtQQiA8EEXz1py087HGMsuqYPbny79jCoyMJOYM3a
zaXi36Zuqdz+yqswzd+En6XjwzD1DPsG01p2nk0DIaa3sCOrkUS/GPaH/FcjHGK93HedCJcpzmBQ
CfHU72dBYXlm99Ow4AIZ9ED9ZO/X5FhYsiVE2k9fIpbBQFsE/04WlHwOEOdSFTrwGprdDeCExsnL
HC86fQk12fkIpH96R8vbgdfb158w0pkGEL5Znk4Nhif52gGCDjsgFfNDZkkskSAX+A0s/bB787eU
Y9EEo6vOLmCTSRhenxDU5uA70cJwDjd/NLymEAEkKFsNeqfWP6ZHyrHWJ6BUjvENkcj2iyOzXvvH
6z3OfHKd6O8iiVu8WinZrhjxxZvUp3fvAtwEOm1cctVSk3uoZazX1/0W4Qum8nABXZt5tFwzHnSw
WxLODsKttlqybyCroDqlFkdxwOVKQThnRFd7uNePLsTOxaAdKYbKfnfHStnBuGR0QznPWGAe80KP
88FPe7HNShw9JsvfFyvOQ9jQD2IPboXz5MvN8+Ky61LJ3W4sTR9aJ50hzkskMv2CgBzKnDrmojog
hkokgV0H52gGxf7yJMquJPil/HQP0TsvPiaRFl9jVNiCgH0ZqSeR7hMFZg6bGjZMYDnY9rAps8Ll
R1sPxPgigTTGuvdgVMwFjftYttluLFUMtkj3ZpHloG/PcilFv0Agc9iy5vXTVpGrE9+mED5QM84B
DVrP52fKU4in/PGFjok3Yk30/F4ixqHe2fu3lsvHNDwOr6BTbHroiF4QTMxnNBgzp0KLxvV5WIlD
gjkc4AhOaBBBgUMs+48K2C869eMraBz8niSO+bbuSaNvzAmJDGqch2HFGHE5x7IIEUHszQEAKI3P
ApR3z1DCoYzTnCVwVJthZGLUPfLDHQ+V7hch9tFXCUIBlySZASQ2nki9nGwWUttnIRNJKJApO25d
Svi5s9CGaOuGkzqTm0XtJhq7d8NWQd8EkfimQYmTtNvTcaXgtGgtEyo91Fyr1vF5klaayQQounFA
apCx6I39Sa3NJJXZQV7VewnnZ5Z8kQCafEi3ADVmwY8AGXZVsFlrYB1XHlY3CV5Gdw8xHh6osw/m
1wxGMU5KezvecDsPxVa/0q2psQnvQ2pmdZVjnALJQMJ01JEyX3Wq6NwFtIzRHP1ITDIoPDe0Nj+m
Is3CC9CLPggbQuja0eN8qgY0boSL28ow5t+rerLN+w7cgOBKtZVN8lmTCCoHLNFo/CCZIcryCiYe
mQZOD8loqqpnQOi/1UQGTD9Rqcwm6btlfaN+Vag9SbKzQZ3eCkK1ScqyJASiWB9BdylaCblCmeUL
fH7hK079LNyIAZ0JnmuoN8uvmT2o2AnlEmszpGtQMHX8F7+UZ99OdjxHTty2VhOwKVxvSQDbyb5n
LPQC0rcOU5A4MdCLBEXkLiWBsiS3GeCUDdGVAMlz+b6TqCO8k8OJr+mK4ByyMTWluRctfxIED4HF
YlEPYjWHlfJguCJSF4hVuR9GxVFD5Ig/BjO0CAa4S/hqKWkdMG8bfEmZCni8z7Z79p+ygsqM7IKJ
++guLrXEBEwGA9rnkpz6unCcKp8ImSBALltiPjOM75XSw4l3gKddg8Jl2aWuIvF47k9DY+5/hlmX
6LzXA5f7OZTkCP/AdbrZ6mJDsHO/qnEBBSklwcHtWwArGBPy66n6vAGlKK+pJmrXA+FP6YQiT/e3
7X2FIcPsPFQSYCHHrgyOWa5eaCcAgIJXRbDW+fILImW9JP/Cu0fUfMhLvdbCaEwxHgDD6iyu/eAk
FZJLKDbHEqu3ugfRspoziw29oGKIyY2PX3wEEITHs57Wi3aA0kbl+1wZfGi/THhY4QDI9Uvy1opP
fDRqp3d8Q+eYLBGlRp2HDx9XawBx0+RJsVU+OmTJ9SJFVpiQlDDwJnvlLOwRKMjP+oAn+wu7n2JQ
axaETpDM5LHwtwAmZ6Q95zn2csWoUVQehkwFMOv5KKeoqxtQDbk/soIT5E+F8d3b5TJB3tfMqCBm
eQsL6Bl5kQZ/YVUWjO2VINUbIe+FtzU/+h1Ha8Qf+0UJ26hNwGj7OK/xeX8Oz5Ksmuzoess8P68y
/CN6wMPaRYhYDRZNW/TZRmK+3AOTCGeqoPj9nfS3QpzDJYLOAaLlGnC60hYXaHiFvpoW7wYL5wcj
LFWJqjc8gqTq/cIhEaaNFb+mTRkr73QzuJ/9Beydeo1dBrCiQf6xskuqcruSxi0hv3ZY3OWftRqj
ks4gWbPd1L7SZFKGaGfZSrXXnaLEuz5rcTZmSgd2f1tyi/Sax/UvgYwiabytazsWfxMkxyZkygBb
qA1XWeEbs2Ow4nF9J+me9A94k/o138K07imj0i7QBuC8paHl/es/svdFHAN4xO0h19zJs6brSSq7
qD+1cUMYiaGYXm/Y/OdMcJ7Vy+dBqOaTdyqViaQvaRcVjGyFveCfT09N680NlMMZLXpsopy7P6Qt
8ck3dfq4zzKqVAhxP8NmM3lzjDE/DSmu1jIrpa07yVICoBubgYpb2YdVKvYDE/7gUOlaAV9JJSnz
EBHD4EwDN8HebpIU2qAZCwKHBgOAllhTBaSF4Lj7Qcnwpv8dI4vOXCC0zINX2McV2K9YJbNoU1Lv
snxl1H55O8DpRBr2xlFMc0grBc8s5UMklBERPgQUqU9kt228Ej8KjteSpK+7CQhDnBbYGqOsmjbn
cP3yFUa3okl9znWU8Gn9ny+lz9pXoqzITRloK4asD9TBKab6yIr+LZgpe+AUqpX7x/V/vXT0uvZZ
Xu63pOrtWLeFtLwekkgxUIw4qxkJgxdNpVftFR1fB2pwKTU3quldVX2M4jAEW0zEkx5OaRreqwfB
A/V/BfQnimYCkAJDjEIBXsVao9bomn44Vmw0dkMm5VLX8O6+DCLB0waL1XNz9XtgVDVHOrQ0ijBd
9a0Ym8cHERFRhwf+pPsHJN3vP2fEAGuuO0gm2Q+aN/RSFRdsmd4DUVINr7fiWqcCD3OB1ShuHSck
dZvkP5xPq3Ugot2xRWT0+Un6gE1m9iSQsTBAHs1NeTVp9AN0dkygTjuwmqKDVgIZ4x1EyTOZQ4z9
sTCwu0YMNqOcieUDLJRYnCxYhQ296Ei6Emr2WgrGesWvf1im7XDvKR02cQW42HbYCEt3me9CHNeC
/eZnqfi82jdlvzrK4U3L+41mG4r7kLbcNNy9wscAXfvw7UvLEyyCnC8d7LKn7Pyms2WFhB597liA
N2T+2a3GP1qRTy5Y3svELo/v7OGQneoNa1xnUvW9INhQZhJGHo3jYu2iYm62rkRFHMaE9DBQrVWH
TtotSFODDYB5olJ3VSiESOcI5+rG8eiTYpzM9gJaoD+YXshggtLQRssScZ5KtWaQr03Zx3A4bOVs
KsFgimO/tgJrL/X96WgMdQbAeWLvmhgLqob8WGmghusCD1Gc+orvFiFto5NsVZyD7iKobQeDcEep
Qr/PXDZtkTa7Bkni9f5hpjFGCLAfW+vWaptoWpwVI63xsMqcMDU+TmgGTg1nyW/SQKMwaAlMVVFU
ET7r15CGmFaMom9m6zKYJZJX3jEV9C0CK22f8cPw2OnwUDIiROLyqU+9nbJQ1KXzZubC7CbPIHTV
8S50NZAggReurUxAFtlp3b5NPQHso5zHxZQTHp1Rue/xCAxfzvF5/gcglRz/6LYu3N5W/MEaxYfY
+V+6Gi7awGQ0xTiuOfGGnAQ/LZKs29yMor+/slEHTNODcXhXqAIsIiA+UKyIaV2TyDCpi6fQZZIH
Mrvow1gmZpptRJWQPyExR0o6uJyr/0VzgMguG9nDLt74BKb6U2vhtcpipO6Mg7pqm2ivjQWTYiuo
weV0E1byDPffzN/0/7RsGdOcbmSEriQbMQJMWm1fytAqdPs6fULLQdfxBtuLnBnKUjgbep2zdMS3
Lbm+k9Ezjf7Gg0uS5glUTFkGvPUuV0Q/M5osc+8cuJ+kpk7OIzC0KdAW7/kATpqFoDexRDLLOxTM
cj6Whj+gCbh6gvZhtrzRsDA755etVphJ6rZylNP/2czeNOUyFK/sL6xf6MQyl+g9PAQTmIRBPwvN
zJSP7f4SbGR+ghvPAk2sPpZM5UwihbwTXtzLV+WRt+6EM6p5DuTJO+WOLnkUzOsVodFnV53UwO2m
bfVnV674hMcbHCGEi6Bz+eyQogl52VNQmnli3lhDV7Jw9OapsYuaIe0dspWdNClQh27AtjEiiLqq
W+KE+3PvlXu33x1MABLpS2PqER0+vLrJPc8COnH49OaDQ0Nl1NDpzZppaz++kp4+mjOh91PvazbY
tKKmzCohmiqXDEZOar/Ilr2ESNQc40x3I/SL7n7uQvg9utRbutl7dEk+4+M8JnxTpmxeloRh5y5e
5wRYqUd6F05CKYPe0fKUj0N1phWudjDOM65SQU2J5d5rW0QUCBV6+V1zTic58C9SnrDGE4T84Ifa
07T8yjORmLULHO3qboZ9/0PSUNR4sIawyOURNEKxK5KhbOm2qBHYoMLBBWdmLoiqsHf7oWXugABv
jppGPkkPcK/vB5dOC3un8Ft4lzsOZPs2sw4wPqnouQOOwLBM1JzY/C5M4dfzVXRGuAf3lIiXknuU
Itk+BqhWmjOWADyrTb6xYND8p3NDhftrY/ikw/nJUlWlbUy3YP/yW9cDT1yfnNMAe3sionC0Gfrl
0/iQIgaY4a4q9LABiI7V7TmSgLWFx6Nll63gd+BR/KDqYQpvt+v8/+95WlyX8oblQSMkFNd2J8Qw
vL/ES+M+0sayGFYc17lpkKM4iIYTz8V9oSb9fX+ozpgZbI6p6dh3e+Td91mB97jtxLv6S7g0DlQ4
CMTvnaiONy67YexUV4AMx1mzTd1X3Ut1l36ZYEci1hCxRHGMFaPGc1COLXr3iR51yH9uLUEPrWgo
MZlL1ALb0uKDr1XrQq6pu2sTs0IwsxAipg1WyVjEvJjoypgjZZyWyylIfn3xipgigYc2TIplq5VN
POsFt3PMQijJPNgBGtOIOGbHSHl33Bn9U7hqorX3BYncBrrFhygxfRg4ZamvZlA6qE1rNqBehtQs
scmgkfDwzjvXekPbuQ6+Sy8GTFRJtyau3LFrq4nbuocOoi9K6lmTdcM3YJud2z5IxTCd6vhZhuQu
BdEuo6wnAwVqJ+1N0fl8uHaM7+a78mN5jp23GoZzVlww+1hqi4wLEUhCbuHxTENheLtdfGn8TYNl
VbRmb1MHB0BRKEJWsX4qTDwlCgNQ/niX1zEY4zuULx4iiDQW5zUEakvYSbpAbcIP9SFgHfmS5c4D
3Kw5ZoZ9LqOaNllGSXKjBg+++fgQ2CDqIBq4SNdn8yRNijns2j2B/Flye03xyjqowfrEKmk91kvx
Aeoxkm1ny8K7vbTWCdyH1M4qKTtCXCuoUi1vPBUec7yioPVHRRmaK67m5pDAQRUa/tyMHOBz9nps
2bilpplHZWTOwDqL3+Ty5xuMBn2AHSNYxadiEhYNNt20YJFoq4F5/arlCVA81JRD5dp/SIE8ptiG
RAIGu/XY8j7WxhpHQQS75TemD3/UhuPLBxtAi+hmc6LPvpPW0h+q2zYek+Xo9ZJOJlmEwNX2F33F
LNwSmFytV+yRrkCNXWlckabXbH8whS5qR5r++P5dS13DVTtP75gRJrdZ3Ht5Z3D523b4MS59T31b
orRTF/JgLBFLAWOAjAHIYF8XTPhYf+lfCWxjENPoS0T/PzhMtKxkNknlbsF1+XJYAu7gYQHHyHdV
Aw6sy/wEGxxBogknN48Z45iV02WFUgZXHVMwrrExY+pF57z0nbFhRdn2wKkaQPc3QVQy0Uxe7x4Q
zaOI8ghYT53n0iNVhkKvDpNjpb1roeBTEJ6DyYA6mMljazH3mG62wU2EgDcF9hcqDXsDw3Kdk8VU
k28goTmwJYihORJ6J2koqblvFj3W+X3kRggQW22LzRPIrMDegekFJeoy0CgavSrYwdaCSBMYpIS8
xqBZ3u3mJdRFmXkyOLsKvcK3tkvua8TWPMOhPdf4nGaOglPb88gK2IfhLscmNuv3n9xdGELe5hJ5
AfVUPa9aH8NDaRFYpH/h3HkKzZDkNkYqFK/b8f7W7h9GGUsQIuA6d79HGzE5s3+ntgrAfEeNf1lD
Mo/FN/dbeEbM1xptWRXGfZtgIstfMGucVfNT7HKZZYC1Ym+cNlKNTl99eTMA9kqRihhw/n/ufvwj
VnOBF8SMzMTydEuTNDDY3SzYbIPkdDUIPYLiujicyBy+2l5Fhxysp7++cK0pevOGBCmKkm6kfnbl
obToj8pYXN2vdj3qlbnrUitQ/d5sGF4spY2vTvzQe560xii/mP7/bGy1Dcp6EAyKu0gk/f3T1OZX
y+TPi8+c79hADCpOCOFVHNj4mmV4MCExGUYvurTJQGbEBoJC4PoHtvD9ZwRJzduk5FiMIDrk6Y4S
DcrVTJqcqA7XsWQAjUMcVkHUS1axnyCEZbiGuPGa3vCpj5vaNo6i+Lc7vUgVIVuBegQTTs/jp2Du
/OEr+wUNR+G6zZKHw3kWU0UTYvnmuqIcKuTGx1rwQvGkeKmRNPErC9ATEjB9kC+K6G/A6q4yMEyV
9IrVUdPtce59VwdtxeRgLPzOa1E27HARwSBmT630maicHP9psbqm1h/q5EEe3ggVT4OiyGHgvTBa
BDXXe5+Mn2xBzt9QTepKNSo+oArR9WbhyN7zP5tgFTVH0gHL7gS2VngvuXXm9U7iAsexf7Qx94YB
Mcc1kJRYCEVx4/d3UhzlM0NgAc01ZIW3gUdetyEeZNDERiaOyebFeBc18o+ilyrABR/8WJh5qVx8
rG6KDnDk06Bd3KRyiQRT06j9SeCGCxRkUInbuTbaCc2xkUSbr+xsvXok13UneMxZJ6N8f8LhJJxm
N4s1NEmtIRfkpwOzA8TdSs4p0O8c8AVlxnD45vfBJZ6dN2OZeuQy60kuBy5OMV621XyiDba35aHE
DMsKEtmrnwmXYqwpDXavgFDOjWNeIzcxJYimAglausDKbG0qj60vYlnmPrAMMjqjnNU4UFe8HG24
074hPepJ2GOyNSoILbv3ZFDHl6lV0GUuJq2Q/N0Duea+3TjpWe2DA5wVPWv7GpV/DSr04alGXaAn
hm2eCa7mL03OtaWB8kTXwp8TKz6TSeJMRaefB/Yay+yEsOiZHQC2BaAzBbzWGlyjr/yJM+mxp+MH
raBhMXe07sOc8x0bb4Go2ueDspLLFp56Gk0+5OG7CK+jKZhFH4x2XgmwgoXypACX/djWWlsL73wY
hckLo98AOM7F4284kfnUCba87F/Z7qPKqrqxUKnf3/yvMcN5VT3z+fchxEKyZNinS3MwQ6PGDkjZ
dmBvDaAbMsUs/BdAH18q7q20KtMBVM1P4+TRM05kzgf/3pk1pbrg3pQRhw5XFw6MhwwYOMmkvXeC
K3hAZhfolduIvfjg1cscjGQxkw2+gJYtK9Oojy2xrOD41GMStA73Qdkfbr6pMzLsNt1BTpFudMdc
bvynU8TkFRe6N+46Q3LVy0cz85wrLFnK2l0KGr45OL+zJi6eBt3qjLPtgtFkXxAajGAdtiHGXo12
eWqEXibIfSL8EP8P3MGZSsva6OOJ/NW4W8AMxvKit23fyHS3l2KMrMh0moYVqad90ZGHkHC6zVhx
7gETvBig8+AR2ruibzJDiDshSinXZf/h70NyHs2pJuzKd49RyvKVLKRnm8NFJzvsw7WkEBwe194T
YAFyjVJGqKqD9C3JzXsnNE7bYy6XzRwlTN3VnKNyrupRB6b77oHsCpsl9PWhIUL/VF2CYLOSFEjF
GvYHlFpB//BMbPV67jmRYWBKojFtZCpPdWv6WttcJYBKRd7nmLpLNuPqNlMynrv5e6Xppi721aak
80d9sMDM5vaiRybHBcPhIoHxTyi2QUOVncZlYdcNI/4ZSGpaGFeqJR6iGYYlgz9ERki8C7FMnfzf
0CCBIYqi/y2SCrY8bXQaqxcA04twlbG9JcMQerJBQPdGJ25ahlku90lLSkTZp1XPClzgkxrhMNfR
/TVp2EIbihlqknaXPfSC6CVP5xFqTxRgFpISpV8pisRoieCxxloVuhUyzJg63janErFlY2q7Hqxj
K7phle6OUiRAngoLhYo2LCQfCjaNmi3LjULJXpmNLVBSKo2GTT2djsDZ8M/lMU/3x2xYWNEo3pih
8OHos1irlOtgv3tU5AbDM7tLcyw+sAvz5US/S2ECeacirL30v/h5ipa/gH1e0Ywg3530VG5a/tZk
+qUMjFBmR9CWe/N7uN/liatQYMPj1gSHDyN6B9ry64HWK7gyXrAE2fv1WDewTRmWhrcTqFGC/QDE
PYj61XKclp7OnCkdBduCB95KRSVT0zm4AfthR/xTxf2NH4KMOCgfSCfgDtCdsOsqJ+l4WbA+cYy2
y0zKosCuauZdh9jil25983XkGNAEdS9I3Uy+yJVAnJv76oPx5a5ozup7AXV4emBrY4osrkPGXK+i
yr/dIT1i4GUkL9uw7PWCUNNT163ICjVOZx+DMj8KOR+vHFav/Z6TONXjDvN+ik3xtUn14PdbG7bw
ndkKJHBKhuP//EeYYHp7ylkabNPbo23DMhEyT6O009jDbI62ihR9eDiF9Lb3T2IXPKR2wvwbDjAi
sxqSI8+a4ZSOh0kSf8pNeQVRigrBgXd7Cc0Y+KMC4lHKUD2PJeWIOCsJ1CXfWa8SrIIo0JImvmw8
Pl/8RlYjRSkF1fFW7lAi0rbCdWonck9HdgBcURLwpaVEaseslZdwUCQLItHcv1/H8HMroO2a/pog
ajugnMP4w0rT/wnUpDOvuqng8mD6Ih+6ae4lOXgR+iT4km9EmTmwFMDsfdce+16DNazlI44gTOuY
Fq7RfeKYEQpQLyhh9eJAa/i4HLLWO+Oo/35YSfr92mRkelBNGAfv+iuThzm/CEyhxa4ZAa6yuFs2
jJrK31Ka6X787OLV4dVJvbsg6l++0Ha8ktlKFA9FxlOO0ZSe1Qo29fLegRfjJtKP8N2jp4wdZQaJ
kG6E44BKT91sdknbB5bjHj0ZkS2pkh1tlc3uNqkTrZDVh+WpV2HqIfOqaFK2CxB7BdWEo5Uysv06
1KcyvAYSuXFFmblwCxCZJ94o5XeV7BAkndK9MvmhukM1iHVCvHTaOFK7pT7GM6nHc+ewbfeppzcg
+NHovWCjSQX4XDlNVgFnOinWQ73Y9ij4aDkzJB8IIC82G8mNXatdZolc4V9cuWeWDzukvkrN6d3o
4gSWfjU0v8pT1JnANnf5T1+lVJakwFpTqBRVDc3czW/k3GvmXM241lH+STKFTOaG6dP1HbMIA4T0
dhIjE6be0bHHsmm/YWgK8h3mI9wyPOIZ/Vv904Z/v5pIYuQpslzXtZ74LeFtbTfxiCIAQk6y84Z8
rkPGde8HBOsEe+VrSf3XPi3RQx1f2iqVq/pvlNBUiNwE9Nw+oRuMz9/xlFHP/4Gjwxb8KSuQU4oZ
cvJqqBESPQZB8Zb/WnQg/LXOBAygjc3k6MXaH0aggMp0NN82uAdjfmoBjqEm+Ir3mVPs6/BwvBCW
NDJImqaqux0iyj63q6Qq1Lsdsto4/WhgmYlInOAa+JVaj70IOJd+NToYfv4ViUq/ui8DRBC23aBy
JX8LD7OByNdAPhHzyvRwyUFc2wPgR6CGpGUpy083LaKDrS5x5gip1ugYVJGAuHpqCEFL6JCueYZY
/rRiddCnYsfOpMaNrmJ3Vjrj0v5tCoSEl77lTYLnJfMgqvs+4dH8/ooGATA/dxHcnuG1gmDGYAFe
Pmh/0iZyvdljr22xSW0NWoSyeK8dT34oOk24jn5+QxylsUfZBzYjxLOzUv3nl2LAxhVdoOPvsv8O
NxyapTj11rbyf2O9SQMf1wKME05iatGmAP0CMkTQiuL+fqJIwYu+mlPq4OccRcqpTuhvRd036+N6
Y94hlRKKxyNz6D7rvCzvehDdH/jz63WbpYkTulxtsFDw7i1z7c4ihdwefXzGC/HOsyBJSKLpZIGk
kVsEJqHMmDhUiwpUdZjAnCLiasjzSweloXUNwLOjTK+iD51co/JGhJj3hLbSk3MLFPeVQn0w2q/M
Q12TJbdr51FZEegt5qChVP5I+IFX8hhEap+U7UhE+uBE9sjJVHY+xw8vVc6Py03HynneqM5SwlQG
GqIPnX3WOXw+su16/kEnnQhlOY6KXu5kiTE4OknN5IdtBAzdm3vSXo1fKBHj8osCCmE7GoLoQSXC
dlHU4ikPyBLhdsuKIVFNaPEU8PiO1g15RrEKWZcoMfsW9MpiFRViVb7jY2nLUutHXI0ujRCAoQPT
AhaKTi22XBL04jBshLd7Oo1jnTtB/+JWCJ08rASVvI6mbnkGiXi31UTa9+IVXAjgSqJE59kpkpRb
ZfYDWlTUqNLNWTNcEJgOEZ/nDedLkOnbVBFiPODDjYfxgSS//Vz3kbrnfZNGPBO4YfrMPBR77iBB
Oa/nx2xCCJZi2GyDvA3wwvZx2/sKGPSCRCBVDqpwPAKTnTtynHj+4zPFbBNdoqyLexkQQUfAQ50y
0r4qyVh1egDBNztVsmj6yl7DichTFr37M6KmQTn2Lt2CLDmiDPYn4Xhkj0KwhHxUMqGtXgXzZyRE
MJrxSfe9nAClo1iY4bwE9PlEV0XQshX4xxcDGU9/IOf2GXx5lQPfqHuk9riJsKQ798aYJjlx/uKB
6VfVaQINEtYwngKc5YdN3lGk90du24UKTPer9I98DwqkBczrDM8B/Nc9weDne/ohekhnv42Tl6ng
HHQ2HBbNrJMx5I+OuOTcZ8Udr3thGomIuZvwjCUgrH4Y6MP22HCVR43NkMHPHIzst3tntbbOb2di
5IFZ4qI9CD4wGwnLLi56gO1qO6/gyvhFeSwkc6xri4dRwijhGRkgC+BCfATYuDD2UVIVoyGlijC5
UYuk0qEB//2FKMozXcKctzjJdw9o7+alaKehkFtDspaEYYYf8KHCKp9p/GvG0ifV/GXP0BP/JCZX
EVmOlhPz724E7og9jEjlLsgwaszsNOd317F80ajRZCF4Tnr/S7XXfZxmuM3cE3n+WZ2roaMBg5Xm
EdXZ3nqlpeh1fvAWy0fQjLSECue4R5qXYJ72LweyNCKv6/eC2hkypzeE9kikDxwteIYP14koC7sp
yIh0Yv7CcHGBMa6QsUAfS5fZ7bk+wmK8JZO3ZUuTCGADK1e4Wa6vcC+ks7a6aogiiVxu0bpMIi/n
9+Juv8SWTJjufocJX6TrQwT72n6v2tSmcm/tYHyMZcnX5V+0+SJvfS2JQfG5k2UEUKgSyTgkOjbp
iAPVZsyrmLUMP64bpoqi3stBnfv+atGtewFNv9DKrIw5C+T6mODFwRGUi/An004qjKALPLRxlFZK
VW0ejd4q+rUvQBx2mGbr7J9FdO9kT0RgiQlPoU9nbC0NxtEGG/ha/SXKT6npoHIZYiLyhPKCqQhG
iH9V9cgR69saqcD5nPTm4Mx0a43lLxsn6uAlI77gy40y6v0Fpr/9kV10JYx/fE6mA5UBp+WGz1ml
rdyec7/V3ThiUAac/NJXcdd0cn0EKcKHr3fZTtZ0p9LKGBEn8NJ46xJ8Mnj9T3KpmK2J7sm2UWy7
QoacQMMuF8aLoJrqH8gP5mCxxbCahp395RlmVl4xFBWjLQIB9nnHNpjCx4IY9mSCNHwOXylO+oJ3
4ABbQKMZk9cgBseIHuPKSJoGhGAMD1QUfKz6viUXdZtY+DNKfBMfvp8FEh1Cs8BFUd3natujFAxE
ODhqDO+h7kALo0xZzIpUScl+QJcqtwllu3Ms+I6xsraDG61DtjsuFl42jUlkaZWxobIoESC1HRhS
hzwmcqjObS9gSD+tU/Oqjbn0VzqL8syIVZYzT9kIlwusvbsRU08EAb5P4tcSGMqAmCgMkh8b7QsR
i3Dgf5ja8zG1Dzw/rg3jx2/23P+QuVTS12v1it8jOR4caajaEnn/3Jg4+4QQzwJ4TLs+tVmHcszX
4GwGIuAaKU6aGtIf26CtZDucxj0WF3U0Nci10uZPWNtSAFMwZbK6jhBGEls9EnYNPwLRam6JfStZ
eIGF06jrkhdwM01V/qtnI2I6gY2rqgPs4rfKVtk3iYkHXfhKUjV6XwbmpPCpEhkSf7oFZuDjibrp
IyxRpQ/8+l1jg3OSuLsgpV0D6DDvZXAa7ECzeieZu3BlwoYw6L4JmeyAhYInlgShUGAS+jJGUlPm
8NH2KTuXIVquk/Iz1hZjfrYOTPWH7lq7yLdbo7HjqFxXPhfO8qT7F9w6e85OBH+lsKNq1q3hUgQS
f3Rw2/pLqfX5RFwHPaQGjAUBDPaao0zQy74YNdVae3are6FXGZgwC7AvzyVMobuO0KtIm4IHNBn2
C8K4b8pRCAMev1JpOcOrX46rvxgD1lORwOZDfeX0BrKtbdfVI8VnGy9/BgLXAvgb//gRqzZYhrD+
aWEv3tMwQ84urWSOUSlG+xDwDzuZERlnG6sVYU+OjzhWp/O4Xc86wDPr1UyGJi15kbP6VdJ2JVmM
iuCtq0/EwbGIwtOZITdJ6Dot3e75GJtCIKGvxyI6IsMnlui8jMyjg4yNoOYa7YDW1w0FUbk070P/
1MytP5gYg5z5Lf7mK6I53k0TZjzOmJR18urDW7rNmRXpv1HMQWRQpe7RBOiQebexxwmO9g7P9pCn
otmqZ5gLzoWxj8ubmu0bk2HBRFfLaFZFS/XZV1rVpdHeUIWb517DED3H/bRvsFMUQdORdoW+RQGt
9IbO/2gTXo5pFrwQuRwUeFLNjkFRtD5JaFiJLNJT9MfNbLXn5o18qzs9070RP6CRjPCWYXXyt2cS
8doGDIn0VZaLqJgsf/0/fKIotDNVvF6fAwOT1DSys9jV1u/d+ttc92OevyPzER0SZqCq0Kif2DRM
uaGNEw8MPI+UkOcXD1qQeiflD0/gISAXBGs4dfsa6P6rF1p0waMheJbo+cYV/49oDAMeRTYP26xc
vE6gb4QsGwf9nbvb2StnN5+kMI0k9zChu8yoQHobAnJP3NI1wLkhChZZ6LAA4Q9yZ8DaiyQY87Gw
1f003YHd2sgf3y/t3UWlU6NaPb7ibctnUq0Z/TL93P+lqku1kwqmAqsEOpiY9Y+IDTrZDbhyb0cR
a1qNeHnClnFaWvSLwBFeI2Z7ZHqlvxUn0RrRI9CB6jsRZWEmpSMg1DGDTc7QorAlqeUkFbqFuWha
Mp9MGI0DK+mkLCz/cUuKYf0KolkP50CVGUf7CvFhWoX4X1b29Li8pHd12UhOlsJHZsbVSK3GLeau
+zy7f3E4ZFrnkBFlpVxTlUYdCNs4oUcOaJCxOdlp8yTRCh7gSmGL0i5pXH/g68SReo80wQu0VhAC
nBvWdUC0tgoyelH/xJKpq8Y8Y7TGfeVLvP2JjMDEVbChVnsL7Bcsxjim/X6gLYUyU6Hjhzm5U5gm
C0zTPKDruA4/NZjUxXTEkxxOUGek1spEz22/ugVf4ucHf8w/QJYeKwp6CRzuhXtvIAJF8ZEf0FR+
Wxa5UAgvdX1yaIdra3KVY4GAxBhEjnunnlrZJrWseyo1ouBELkV1tcBj5JpVg6WQ1W+Ue34V3khO
bYOByM2Xby6EY/89n2Uya3MSUGoJa4nsBlQITqpOjl/kBfPP4vnrbWqJrdlp3LKvZZwsfmLQuolN
1iG3+qDgsUBJbsWfog2PpLudJsRju6bVjMmGpZwyPrjMn82WqS7zjdNtL21nSzfOs0Sv5RFaMrSN
CjkvG9d4MihLrEjQ+UnXjI7aNjlJpxHAjpkZxixQE0P/eDVMWb2nUlRayg5ChX8JqqoWZRcdxl5X
scA4TbbDFqZ8ETm2cJ68iOraaJafu1zOKtSCozbq47VW9ajYEKCYU1vMskhixPLGQW7BZTnFUUJv
6ePBk5zYp+DVSmNIYlj5EiULJHzDZxwKy3xEBi7Ny7KNRg5HI5QBuLxsLLqwYwFQbPXQtnJsAGed
C3p//NQ62YGkko2APlRhELEtJ0W2MnchSWkO7rRL4lXEW5SfuH7tinX7ux2WcGbT2OLMGyUltD6Q
J/Dj3FJIkHmZVkxsiOfrWMufPJ8V//ImdOjZJ+zDTqHhgIy+fb/8PO8ZrxvA4E4BrI2rOWKc0bvN
JLAn6qONux3nQDUt41uFyQyO9MZpE8y1mPmvEx7VzBQDSGbzqMiwMZBI5GGSDfMpMuUorWhMVZ1N
lLcsQNE1vCDnNG+bKLE+q16i4sbk2SS3v43VsgDEiuHlHqrSKrj2F8AIoZp0CiPNt0jkiJusf0/v
NIFQ0ry4UbYpzbX8/2Qfd36B90E6a4I9UO1fY79hfw7tyLA7XnjakRdoj2CrWTnyofzJMi1h1JWH
T+8pNjPC7hREN47YYFbYJQA8x7WNqgR8kpvvHEmz7FkSOMhQBVDRh3Cjeuw7xbrXkVuFdBJt44n0
vvulR8Cd0mtrHT5Is6IJUIvGZYT51XKhvB1VxoOZ06MDU1XV7DvR3yLOg1UQ2N6UQgIrAoJYmhGJ
u1NH5zRHZVW7fDI7fN/cTBXtdoiC74hqGIU4zlmnoBnPIDI46GjRC3lyEWGVmiep0EbUQ+4ezQKN
wJcYnAshZRwqQ37gTFPPzHucRJsvL/hsg1NffTr/01OW6MYAKsXXKLc3wAoLWr9DKzX7jjAfGfUO
/+dodyQZGGFJMTwPKXpt6g1yuQIk+5mUnKiGlaNJ/MB0FwWapa2Yj963BjT2cFw2rmz++FzQv3aV
58bwDpQVtUeu+exzvhjRC/AcCcV3etEht1qop61varqYXvn+OeNBfvwf47Kst9uXSbMxBJSCloXS
L1NsJU9BIQmIlBy/aPxp+V8leSOdsq4cOt0AXS7KZkSfY/xb2Ss/s1hqPxxrgRoaUF4CZpwvHiTb
1m01/jXuOBfaCQZwSEoVc3xcjroKV2C0PnoJHQyxkuGF04hIeZGGgFNcssAEpsPDnDGrYqYkDCHu
qGtZ18Tqb09BipfITyeNDvOQU0ZYxpAZPM6ny8GXws3fSWWf2lTHNA7ctiHoBhSI4zlHjn5o41R3
AREpo5bK7VprSQoHmdhxN2V2+XgaN76rP97GX8K3Em2nAsu6bCkBnEcSN1C8v56N2xH7iEgUhSD/
TrAxpac3wMUaZmpj1+fhrWKDp44QtysGnqnZ4ehOTYCogE9jj9L68g9X+jqP46PLEKWG2MDQMXVs
mas08jOEVODeyXayYyEOGBnNkS0ZElMzecX+FC/NP+Ov9dF75NrTT5WRoTkrjkWw2XgAT0CeL9SX
IOzJ6iVlAwoBZ0xGdERUCwLNl7L2iXoZGizkI3Kur5bIE01RPgpTs9v7WpVJPh/PO31JAEHOrNC5
pVVTm94Jw7b/+jq+AwU2TDBHRalRWOP4SdrHSpLKdo3woQgQlzmME0NjFLh6VWuZFZZddoD6srjt
5XeaKM4V8g0Uhin7+9ozim+9QKIV4zxs9bpPoyzwkoztYnJiEcrQU2MNN4puow9eZGSaA/kVDNMU
Hex8uIFNXoHPAdq6jBEi91dCuv1RefLxyGGYiPmw8v9ihZHQy42U629sepZBsdWV12oHdt3XfWI5
ynLXMhZFLbc8cE8k9wkn029ITNVfs8ZA7iT7jZqK0uqF4+isPU7zDMUF3Tl261leTKkZUEwwQPxI
XoweYfU2o7N6wXQ/zzHL55FQotHLxTwEvm/7LwAnyc68ev9hOcVkNQNba9uFVLfsQ4KI9A6e14Y3
OxWJi6W3z+ccJpzYDZj9WdA9GihMQC3k3Pot1K2RYtN3X4y0WRoFOyrl6Kjp+gPuAXSXgjpwcYr2
fp6uFXiZZd5X5a+sHGQXnTy7nQAXtCS9F6j3+awzGk+vIY0nhWxl6JFSKvIMYVZU7uC2V+Y+BCrR
woDyhlUsLVym16T6JfyY4KBPa9LiZoTd2EDjAgL0ATf0lvFzStmpFvRI4p6eM/aAPatsU56zKxHS
ZZ01M91kdn5hoFxImJzHIkZQFtXfPerafdDAAutrV3qFoTCNIdxiRtfsO+DL5mwGx0N3qB4JY3af
fBgbkl531kPeMo8wfWdbCuHw8L/jBYyQH19+HbTS8tJCwtluGD+ReVqCmEpRrE2cBE006kem8YsN
UqEb+kSHbtOiymzR6NlPintOuTIGMqdXA+oWB1JZ2/n4oDbLSGFaDQn8tx8kumdm3C7agZw+d6h6
4pustI0ZFcxjayxrmU4dCH5VtEyBKwwlYsxYeUZTBsDA1HcNs1KICvr8CC+ZDEkOixy2IO4KyLq8
h5sMS8z9BXvP8TSCAPEqN9gsTfXw7b00wEsrR3jzEadetcpsSN4aWWp9YPUbGpVd9wEzxlTo3o+u
otIXekUYbYCjInaFQHXTeDk0UZ8Y9JbA+Ra/h5Q1j/3Mllqq8ZEFuHFVKQGlss7h4As8kpRl64WJ
x7rdGsLekoncQ1curlEUEIkRjwf1D3lBNESrqiZyI+2e3CI6p9JJxWZGjijbI+p2ICSHPD+v5uAw
cKE81YYE4wOv06Sfm5NUK+n3E+dsbog30B43VqQtdrTzpE5p/uHOsIwP9jx49zn5+hpkc/jGIdB6
7o1ep1Kld/CSQCJZ7wyS3WmZs2mKlBmsPjM2a7PpwXORAX59/ecZBr8OiUn5TIki0aXSYg5fpbvH
xHSlM87YDRDyBOg/Ra9vFVboNFl6UHftvKGQ2rv9/cooceLXwI+SarSoiO664NEqEdsgJr7YPLUY
+O6wqFnvWZpVV/xI8UJkJNqItAlHTv4oS2d+gKAGTFMPLobOz09wML+zhMflpuq4XoS1aXlP6ouu
ptPqZl4hnQJhcFhfYYLU/91S3WEqjZl2NcB+gKyPsz9H9/tIf180Ovrdl2RQzhppDGaO9rYXaOiE
cnZMPhCOYgJ+j7XeTCyK/CQOoFjEtaXCpKQb8ib7jkyMxc6ykw9hivCX118C+lT4RRCabqg3kBcT
FhHjCWEyVFQrDvw+dk9WhTPLHzdxdqaK5oLEcx0AQ7HW0dbHcUVsigey6gKKBulcTAwzSvWIntz0
NhzCRPx5HsP9uCkxibndBH5HkxZVoUA275BaqkN/W/ZbOU4I3sbX2sqXzYuDuOlOIsmgsZ7aU+F2
vrvT+4MWweqcw47wVHM8nYJNWyTBIEHHdcwS+DPUExcsp9qD3TQsfwgu/+F5BSMcbaHV8L4U4d2a
HqhS1MEpdEGp+7pyZqRRMc9U7UbRjKwInymGcSGjuMJIffpE1nZh9VxHTmSmavtpS1YlBWmm4L36
mucsg7L2ZkwhFMpLyRElF84Kkpsa4NabIdiwGzJu8MsQU2sP2OqXw/baZxzNQDCMcyRPaPU18ffz
ogVZ98S3BxxTWkhrFD+z7gxKEzxybl+eoAFO0cmcN2QYWDwRqBDOuVZlPh72zctelP5nQG51yoGp
o0fVu679rFyDjCeSCW3JK8M/pPvBvRIIAMdQKZUX5Z2QQgu26Jp4Vh/20FnupMAS50z2GVhPBe7A
NA9mts39UWwG/TeDyhjvJRBkm6qOHUhm3j+OXaOj0QEqk+f4ULgRMBWhm4Fz6Q+h5b7eebmfspRK
9hHzCaY8u2ImwndB333ApYNHenrhaNIOijxbyS5xqpAyqCAAKt92nqV2v0oXCYGO2W8AA9V30quZ
S9cXpUQpem37QTqV2UMK5U+JlpeKk4x68RdgWW4CExvVHl5oUa8nNOZLeh1bBGf0p1Wkvq0ht/cR
Fe3i6E1WFiIesf9TBDtWkmoBdgbLxSDu1ulx4FpLTq/FAHmBfTvx5S/tD/qVHA9S95QOpVzCcPAF
SWwu89flyO0J7IvPUHYtNgZYmZgeXZzXbs6c94ziEU/kORp9dfco1w1vjcFE6IqQdIEpBARkaGay
TjZ68MeCzdattZM19RWTykMlRWYrtAv6jSHxQ6+jHKZm6MdmWYj7b9Un2qxgW+/hV0NqQh9+5QWN
5q2eVdYI+1ccDdU/6ImFinTuC5tAUrZV7mrxgNZ+IlWhv/p52lO/mqAfBacfGfInaHfyJqQjosgC
Ld+f9bbBtKOFcQ5bL+maS2bKOPLgQ5wG9fGPzStb/fvtMm2yvKSZkxi+2xRqd8NA4IbrqzhN+WkH
QnmeRo7v1rcpl4fuWv7PYjV4OiK3eGdwbcwmObFWP1LpHKdnJr0QTiiD43guoeI5LXnxV0ARQUkR
R3MgQFQnDPS/up4W+QP5iPaiAjJqT6tNn1hZhUtOTf97hu6r3v31J2wkVWr/Zb6brYQTQInPTG8E
epVXucqPidvLU6P/bU6wN+pgKjvfG+2mpaKaeWIlyPtnBIS9Sc+y2dn0Sar9hU9W88oPja8aGWpz
hAA2SbEWeutdDSXa0B+GiaOkHINSIgN8xaMMcJ/0Ci89THnby3nWuI9ivngkXp0zAK2aR0wZDa5t
pgXcOFHirBDVB8fWm+7jNjCq8nDxEfNMY7oonTQbsT/E5yV/dBzcB52k10v/hUjxIArAFqarGtmy
QE3c9eSc9/YM2ESW/b6DiE41zfYqGDw6xlQZplfDXn6EPFvli5srr155Vi7f2dXwMXqNhZ4odmzp
mdBDO/YXTneQAMKw5HRMNiUAzUJOg2oP3dw0vrNnaemphBKMOQCkH+MwvrZdW7gc7ztmEBRBcWxw
U2ZjEaEnhdBiiZGLiA4tx1VRC0d/OPAKWWBeqSeYLhsaVOYIKoXkrZlhz/8ya3BW4c9rEcod+zhy
MgaxyKi+ls5ceYvedT57jeKc7abMiH6U7AqKdC5bsIBnTO1JukCuyJNGsjV7fjatU7kOAAa5LiZA
SQ+fxwAvPbJY/tvh+DyGYq/Z/cN0EJjbHkHlSUys45P2sduK0xEU4joHHbvxO2FhUjf0fmcHC2kE
OgVXkemxmS7WUnePytMPGfDBhLT16Oo3L6oOxAHAPWDg7TeO8GTU/vwNUcI+2WbVr8IArNP51fjL
LLYJVFSOdstj7x+/nxxSGKfYsZM82ftTDjZ+mBsGwqLmpZOVp0ixTC4K/ftCaZOCo4kNDLLqC3Bk
izz/x7jKSC6RbEG5/IapycWNBl77CK8yKPtr/J6wqrJF7cXoQEdKbchtF8ok4biyy5fwtvRsmSUa
CcrK+KlgOlMO+WtTG7GdXKHqS2iSqt305GTTUhldkbb2L0qBP2qPwjZ8KWkp8M4ap9gLSJ29Me7O
RMQL+6zG/9ZbCJZvUrch+UkkqCK54q+nLd82pAOxhlo1nOQCPu4Wlrs4TX7bI/6K81UwBcnELalb
S/T6ViRLKQZagAdJTGF9PkfNiFBlf5HJSWy7uF8k+wppercGHqAbSRhKhL89CrllZWiz+bcbu4Pc
d+iDOkb4W0iXuBcrA1sq7QKhHgcnWMWTv9VSaerNntfR0izeWVgC7fG36bfr+opETDf43x0Doebx
J6KaeGFJN/vGdgDZjnxyMdWRUyCP6o38yVi4+jnSm8JJLIzd4VJ3YyIPXalRCzXi3DJXv/vLkfub
aW0lE30FI6YjUdpkNDYnEqni8GYj+EMho0sVgFLgb0er57b3ktvXjUfjiSMVQNa/5Lk5M3LGTZpG
3FyRX2xXEhgEDthOoHvRP8qZLgR6e07MYQIdVYCI67HdLVC+9R5Y1WNP090ry2sy8y/RtjQHA0Ny
NtVh91ri2vd3KQpFe/P604MyTRv4o3ESdQPWf95uqNYDEL5pToXGM1YEds1PRl8MZ9lARyT/Lu/W
i5kjuZJHFaXBlchO9DztHAw3RxQmov0jvbsQl46frWwrKwA2wsOI7zBl26oZFOtfb4NkQ/taFX4A
mpCB9I6hrZQlYMIeytrzK6ZECHcf2fa12fPOeNrorqMYmj2/wFncp9pwBVoyKVTjuGiwozk+EP6G
IO2XULIRF9VRho6eSAY7WdIBRrO9cwaPGxv2yl/C8H8c0DZoez9OXEzll5B66HiykSuET++apER7
lm/WOoySc/r3d/1oNqQpSXQqfPuM1cEkSA7b+LuhDnCkba1kndvYfqTLQ1KT8SRE/xHq7KRQmoL0
Ix2jNkIoz24mTWwuIt2R6PDegUWlctE2ESVGbfs5eYVJnhH4kMamwok8w7TYYg0e7+/Gx64r0uls
BC0rU3Mc2Jdk+0g6NXOoPBSFGFgqn8CEGwxWKGMlgPEmECz92irbGrfDFQlp+lWG32y/Pdi7W9OQ
UPwI1O0fwJ5O2Cxe9MU8lEyktEDGkCJB9+K6Hw+36xvoCs+cytEsB1KsIeo5kYZ9HcfqygtFsxga
IOOWBAH6cm2Amy+w+2Kj7S8c5k8YUz69oAZheCyvjg5n7kpScJpyrq7xbmK0z1I/LQ/FCxvSMwds
nOBindT+OaS9RjAP4XC3dEcLv+sMToQ/KCC1xeW8CiG6XLrs687n62lTzTsExHOfjLkShL22GXnA
q71QQJVpJRbU2HOvcCwdhZG2c41GJmsysvizLoc7dlSHClGTfoyYHe702tZ6HZKVYX4iMa04SBoG
nmI/ChRycEfyihpXKsVK4anAXRAy4UcWcan/o9DWVWLa0SHcIumR072GfSdlIzBe/Me9B84avXud
/9liUpxNrE9FqRDmFVS9fnfjA1DXxqEpkhMHRx8eQModLZk9cWpwwj0CZZ96nSlVupwSWVd/y6pi
4KnyDKWGMKvldpr7sclt1JhiPQ0jOlbggEOBDlv9GbwlHf5GhKVZxiZKTMFBSac20+0kkHp/wbWZ
Mga6MDT0oAE6QPVURIzxbuXa8xyslUUWNxoSb+Z+VkefMnBJ427bFPsTNfKs7EJCZasss+Khqw6h
xP6/p0j9RDQYgRYc3tLIJknc8bX0utltWrJj5Cpe+VQA/W033X7K7bWl6AgWTWxpCVLWlPwZEzaS
twRJzxWJ2HlG2kaZnxAan2T3DGbZ1/hAtOj9XdOs/rcSeoa28M9Hoc1BlduEEnj03ZrP07gICTqj
XTv5FmVIF9qaDHAgfbpWlg+hdSjaBwnJpKJuCa4+mXnESz3sQAUbU49Ga9bM1qUX8L9aYBrS/l+Z
TJixDtOVlb73z5RCDXqevNNSqQbF7kqvYbd1qH7yWEokbqM3b8nPs0vbQHxenqoKUsxadK7E0ixV
wBv6hrGphUYqwhUgKRP0O+eEeo/sN2GpPrPibp+tVbuBoySVFaqWmOoqiSa7n+CMmeoaW4KwwPzE
E56xER/jsKqak1t2aj8+hb4HzrxWSo4ncHL8VQEOVmx8tZz4zWfJ6i3hZIsvGFEvgk1oZlFI5pn7
X4+mRwAiMddZw00yO7CjC3RhdMX8hAGSW4XBCYrn8zPagpSDPTbzISzFDk3Z9153te5MlJta25hh
qUklbsEilOPwiAsVjr3Ku8hzhzmqrSN/L+2pXljfXImPWGx2C6lupnReXg68WPgQ2zu8HS6nnill
RE/nP5U6MqXciYjsCiQo59yCx4V7AyfxNT65BCivAnleddaGvvZ6Qrd6J5Qt5W35CM4hGMCDJ4hX
yyBNuiEsuFg+qwdVf06lC1Fsw+4YDnV6X+L/3gpDDgu7dZ6zKl/+FSBWJaIVEi7kypUgJFMFdOqJ
XVWsJJ0YTvhWujdNlp2b7qdNoyV1M5mjRp0d+DpIWvWN8aZoSlvRgSWBaEYPN03pEHg93eNp3/Rk
BM+lm+6ThpwbO8o2aF/uzrZnePxAcmrn+HaX8+LbSfLUX3Bb+1+wfk/EVkfqPXr55ZNfpbZt8SB2
lXL/KuIwlDLRwu2S+Bro9+REweL4q/IHjhtPyqOOTcLIYFrckB3e4DYf2VdBfAMNNF7xmCenXRY8
Lb6qbnANKe+1tO3rq9xnxle5TiG2M3AYSPcXO7z380BXOf6AbtsC//JfcF16RzpWCmUcUxLw7Uix
rx1vwGU0iOckyoBoyGq7+B7Ch+m0xqAzXMTAYiSvQ5HvNfei3OdA/BHANLqPURgtEaBcyjMrRmTT
XX0E9951aesq04igRla2cnV6RsB0Ya+KuLUE+jvfDym4O37OfTzD16M2xzUd1MFlh6unwYL4akIe
mQrXoa855xa1+6FCG/17Fjxd01GX88kRmSsA1va7Qhf5TnZTpXIw2AJls8zJHCqSpx1C66SXeKqV
gfaSzMVboTgX4rUBKZ98gZuob4+MTm1KaWUH0VLmfznCABQtkHjO0fmNbbQ92929Wqd4g7WSmkKO
yUizHxlgMzx4BROZj3v0f7L2QiVdUCY8UE2uOPe85JCmWUPTGpt8XFyt431j6Maasm9tEPOmYRf4
J1xW5wIaXsHt+jgGPWXOllH+opmo+NiwOGcMO2Ias9Qj3MBRxcuNQYrLNsSDVscjufdRIDttpoX3
eV+cYjEZCkaicPduu/3mBwQIEM68Dvie02M2mRhak5h1OUCElzxt63rvU+KvL/VR6z1OA1QtoA5+
V2y1FRz7eTLYzy2YXq3ePINzdHPj+MScI1KvXXKkDtRUN6WO/HsMONInKns8NXUPKrAkUQkFDLek
+vu8xngFCkIo0dmQQ4WmB33IdEdpJ5glAD6x+bP3bIubLdvFJiDvLW8lg0pc/+tnHnw2ssY0Yj5M
mMHFH2wxaaJcDY2fpl1kHaBppyfkhkj+HPrB9LYt7vOa4JOaJNMVoqZYg3rhz4irx0pe6fN7uf66
IW3kU/G6ARjcicS0Y95A//hgWxQrpQiH39HKLZKzXW4g8XPNq1JCUawNVT2R0qgXHWOjFkkwrr09
hR5GATuKnDw/2JmiV2QvavfQVswiyFG99hZAfznGSMOIejCkcTD2wOtB5mWBtubRjaoHPghrkBVJ
BiCojZSZ5bBtjqgR4scWLL/c/saB5iw+f4I1orq0bbwIqpwxxfBzZxw9iQ/r6jCFBaG+HghS+ajd
Jd5sMJ+EIaCvJrFP29qBVKFSgvq63Wnxpe7Q6shzc4PbjBZs08wmtmuiw4MqPQZ6IHm5VP5PKhMa
fi1xWqltLHJ9EdsWLurOwbfp293N7l69A9sI72kg7eKvSNNLwOQmiSAJrX8rdKn2zmCn1H3WMLXD
PdG+6fpVytSILq6zaEauSWIlU2RDKSbGzikFp9NbJQITjnL6ejVMmAODs5C/uyvID0Hu7tXvoRix
JbLjG836xKwGveF7YOzNQpSnG3eMZphfLEEM4kW5nLCwgy4q68B9NtwA7e113YO5m8kOAx/nik4J
ObqDiedTVVINBF+q0xIu515LYQRWOj5FLBWhX3+u7WgR2LOh4QOyvpEKyA1MhGIj/fbt9CzUpkr+
qqC7FULb/CMXdAvp491OavsDngy+wIrtaUtXA2ECQbMGd3yxQmfw6uLh6xXJeev+sWlRwCzsWAaV
XuPAAL570+F0l2crXa0J6+bDXKXwiswt+TIBZeyTIMy16TKcIEyemNo9MgaY82GV64lcI3g+zBLV
QVcFTWy/AU8WBPykxv4AO70jaOR41Qqe9S1dGp6OFqGRYlo+XTgv92F2u1zEux+vR28s+a5AMT4d
GaUnEpNYkt7YYqMlgsqjtjc0zb2kxciwtESV7P6CJFeakOEtVqsQ3IA5NQUbx3tv2mZ1qjIbSAaU
PM7T7ZS88iPy5mJpyvhny2weKPVu0IJFjpK7Hy4TUm23LrGXeCyWr4u00xraQsP/k5oRM+X6QDRs
pYYzmVhFruMCBegvOfvFBfJU2NBI7kRyjFz5OLq6y1M8YyLwGxRi1kcImiCmmld3BNXJMZz3w7AI
y8qryQ4brXfQjvgmmLEFcKJiH7+DRnYRuF0AG8EauCsJ1jpyd/X7gsr/U/rE4V4NqOjzHhtRsElH
7iOntoQOZEpS9keKQfuRcn50z+H0rrWutfIHkVZ3jYRvhcIwDJlI6hDh6nDCjsyk1I0wH6WTX9W3
TatBnfB5N2l1jWRbaAzR3g+MP8VeTpre6wY/jb97Pwf+NlBELnCa/+GNpk4JJ9D1cIB0CCm3oBGM
EDfGW5BJeyJuEf7lxgb/1EM+++83oUk7unYhwa7Pw2FSVVFpA4DYXzkwRQoXz6z7f64NOqyRTVjn
uBudCH1QDCzGoWolQivJ8pVk5k6PicsjF7CWIQMWcB4hV7ZHSzgI0AASbYyZAZ8Z/fk0bmXmMBwo
JO6nC9jb8TXtfveU6fcJQ9gJgMi453M06bLDc5ANFZ3V1TjNge7avirAazdbkVJT3un6MflVYIK0
bexGv58Kvm1yO/9LygDWCxgfvindAKrtxkY9DSwNNBvS0hx6Ai2dWBWIxFkPHEJplZ6Ub6JLQnbT
mssMSqjvfb5QIggZS8Oxbf3Ob8+aHuCM4du8i+ASl9IQw2xZM5UQNPhzC5KSMNXRz0hUl2mt0c3B
J2NLe16+V6VGjTHGo7e3kqpyFc8FfKY/VI89xsIgm1HMQtbgb5gbN+5RHNvRY2MScKBxIRMgwp8X
IdD3lVp4qgsJYL4Ke/OkKJe7K06J1SVpaZFC3+0MycsylFFglKEq5nn/01Am/nCVKhtyPyuW8D6U
cuB3PrUDkdVnB+6XjCKbouUOyjp4pKRJCkvPioHiE57CqmY2vka469FwTwRtK6dQ7aO5y5ODeHaz
rmxh1NqxnmMMPKMA9MeOSlBa1Y4ICd35ptQ/wgUSbiECOjN115jVzKykqzfG/UCysaaDgTqZoc9C
+oX+MD1Pbx5rMhit2U6AHh7Vpb8L36g5XC2s7q+IUL5C5Ki9I73DuGogAEBp2BCZANrsSGTuzJJR
zboC6NgxH8zcRAQFF25Frxg8/FzTqgAmPR52IL1mDbZV16lNCm+YovJLjj7D4MGSa41c4gWpAtRo
TvZmgPM5PL4EhA037vn2uUjD1ijUhBdYfUxYchPBIAEkvpe9NsxjyzWbdmp0Oslli0YmL3CeNR4F
k+dfsWGM2XbljIZ8qL7f6pSUpv3RUhJrbQ58b2YXVGBUGUwqTRG9r+H/PjaUUS0VJOMx7Ek/dGxn
D0xaZwlW5/PoQY1GMPCAFTNxSV+y1GrAn/097Z6+5zJcGchnydt9pT3zCZiYnZQunOpCqsTviR1b
ifzJDUuqA04wzHOWRnP3E1zYPYNR+Ih7soymiULdZh0JkS7NryLuh92AfLQxEiLE8qSZR8jpLH/S
Iu1tSE/20vdh3zVxDxjslczbEYxIsCEaYmjcNLtNXVQ2gnDIlKe8VpioNbXjcR5PTjLNMHU55hSV
Qbf60TeMQ/lXzMl7BCA7o3jyKOLir8ziQ/KywApT7qY3I9mmUGUwVSIRRojCjIAPbl2N3pC6JTGa
q1JvwT6opTErOR/Y8dEXuZ3Zaiq7ejp5VXYg5VDIeDWdGXgtZs2bTAOHLoGPq8BdUxfni5DDxRO5
VeSrwHd7vYJH9gF3Xk4fVEnBJM7TRpyrB+DCwsrK2SX7p1x1rAYkLSjzEhkHXDd+aqNcKWs7Lr2Q
lJa4u3HUhkNU/rAWX7+6c51Qbx4u3MWjmHms7E0C4mlTqRpgmUV7/8dTyMgLGOF4oLeppAylrGlA
btViIyHtXPmLyGXvU7a1xJbzy3pp2qCwxGzlFOW9kdQOntoanBP/HxSSfHnx3vIbv2qpTMvZy5vM
VGr4Jgf+GbnDR79WZy8liYodJ4xOletSjYB/e4GCNKutEf1hl6zt6KwQgZa5nE8dNiXVdu5BF2uh
VHJylE8BuavxdjUEuxzKwaKDUh3JPT/anXh15wpvsxNN6jAAjumelVIYJRlQv027X5H/4kmD5a+C
48peHsTTVQhjCEj+rGXdBIVFJrX54+vNlDN47akDON2xdB0rjzgA7WxmdzqKS9lxeNDzKiCYTYWu
ULpgsGRDlOr9mM/VvfVwKs9vPrjFLhEzwBgHUsccpXq6uoNgcQQ2J+2SSOwNQePFLkGLLz13rT4Y
Xh2jMj9c9VIWba0jC1LbTSLgLJd3vHbcQYJvYixEV+03zO7CPSom7qGDv444j8eJcaJGxma4EmGO
cE7uw6sg82LgQaTx/SFNbWgcHLWPFDwNf/a6DpD+QU26kDf2MjYlOzHrutJe+vJWXu/Z5Xxy29Gf
T2tOcVUmgiIBkZu4zLpZh5IJx3IpcjQPYAbgG088nvZ3d2BxV7aRNr2pvNGfcBQJHHlSpRvojXD9
7Dt53/uIDmBb2yMHXZbNwCsbCCrxgVEmp6bcm0jzbjSU3RIFy5j0fqMRD9zD+TjMsK1hF7krPiRt
VDxYqaaM/kEcVOE79kmmDcCUtdurTFalQ1hn7Gkjh8+CFk6JIEJv89BHSzmwBCfcX1C0sJx2BSuK
91dkB3gNPcYRH3Fd1vuqsJEmnWMm3mVRikOjSG8M8Aw0lbThWQchFVcPDaap8isTcx4Sgoi5mpKf
oeSjVEFkLxqQR3Qnzw+dgt+/GcSCNq2mTvGG45HlO10QTIU9WCPEajirM5sM1QEqFG68nUk1bUOS
SDWOhEH9VHpcE9oHyhZu89JfthdVgkwFKLR0l1oqp1i3zXpgcd7u16bINLoyBvun+uFz1cyJKLQn
HpUGQ5dMRFhHNt4J0n7SEZAu2aO+UMoktVWMgn5PrDPKr3T0O58Occ/5JqBtWh4QxeLZRbUP7bIi
IdysrNT3rF4bjvDaJyGacAbSBBI3w2Ovqj8mNvRAxruwrx87n4Zd+7TiR8BOBmxQr+gkX6q8+u2R
YKkK0Q1pMOp307Lp/VloRj+Fymk9EtOdkgpM1erFKxh/4Q/AUGZKw3RLjxwnsbNFy3IEI5DK/4Oq
jkYXiq9JUb8Qpc7aAeMQUy+UvH1U2JTaRdYHwqyrQqBaCrTUUzWcFnzo0QvKQCeJ4Jvg1WC+s/Sp
dBin/rgxO+OLkV8wzon1GENcn7BsQVB5Zq0OOYBS7W4N6IxvFEZwesaVsH1N28gHSVVvrVspDfGl
WgIvIzpkcDYvk3rC152Vdh1uX2zZTWGFoBBYL//zEHG7sVwNSutL0zRzHunq+WVwlXrMR4W7CAWZ
KKHyOZnymFS5BRg7dMzx7Jxcho0kkOeqU1OSrdxfOWp/8sbTIbZ5NwGIx1XHpHl180Vt9T3POxBq
Ocoa27hh8b1dtX9wj9XOiFOR6XjBJhKlMnGVNqQ5XL8Gm4f87av1ZLarjs0nf6pGJFATh/LOV30R
NPj7ohulIWiN8hjcFl8b5pRc8noJjyQM2S91xKZMt32PPawAUDLf7QZj6RaVduE5GHhWZm7enS2Q
wHyyKuM5VFvp5f57/z1JjDgG9i/8Eo/6uB3fxxdqafLF6r09K7sf/1F1tINStKXBL/P1OtFAokB1
NPUJetL3mh8mojYZvvGqhxfHnMNmxMfPmoNzsfR5dSlFVNu8ZtH98hwbbkHqE8LgTKz7q432wlg7
53d0pOPaddbQLkpPa5OVOqfgFDjcB5oEo1EE/Die9c4S/39htAOnupMc4y9eIvmW4IKNCloo3JDN
mAt8Nuxbsad+WIXwuu7DUyjN7NgTnuAhWNe3bI/3P0OFNiFv32IrrQ5Vr+6qB2OpAzQM8x/9K5oK
nA6dqh516vU94F+wR9o/IDG9u6Vko3UYQ7ydiKzEbeOIeN6Uygs+afQRoIDTIoaSe7R1yp5ji7Oa
0CocmlUeyeO4bKkp1oHE169RsB98cTW4A9iAeAYHNPtFdrOvP/ay3HTW+NqxA12E7AOhY5FC5Hga
DnaL2dzL5nijXEi2JZiMzv9zt6UVk5uvDeKM7coc1Puk5wiKbfOr4GGZd+J4fcn/nkcjfyuyz2cl
DMULq/LRaw/4/5dpS1nj86Qqs6l/OxR0SH2LAgZRiJaqNhEa0rxZkJK3c2Lf0KADXQeOf3tt2Y/i
re5Wrfr6KPSsJFU2BAi9hPwJxg3iQhmYMhoML4j5SZCDHb6HEZHwJ+2BXCiWmE5RedTWYlhSmTyR
Q8UfuAc2Yoebt/g0LfhW0EKISXc3pUMcYliRnzHRU8vDRyXt1GBUZlTLBP1odxxMV+GoueoT1EwE
Dy8THmsQ9W5yCJfyI6VpK/O9SRaZ67oz4YWfz6GWtOqvu7hK32qnUziAtD2tSAIaH12q/btsdICV
wnmjMSFqlcc6a2WhyJKBTfXOiu4Je+3TmwJb1QLGjN7VjnSfbElIfhkpXA15hj/kJXGYaX7NzDKj
AoUbScApab8G13QsGG9mtcJFPG49JXB6SfqeFJC+6byjQW3hLh/MekxY58jXCMXOO/u4OOUYHTol
zLvw6aTIfOqHdh7rShhQ13QB6rob0Iuba0iN2bFPt7fwoLcQNp2N371n/13EphOmlJe+3I3XB2HU
+12H7CVXMEDNbvK7TMCDhbhf8i+kErzdZ08PZl0OlEdOwlmCMSuVdwf6wC5OhUYWvGD7nn9vGr/e
Rjt7o2SOmh7QRhVLaSFJsrhO23oe/D1NaYqlpJlI7jzJoiJQwUE5Uy1qS9E2IH7Q2StBrcZ2mmp7
aKMqzKxmw6yQKvok0w1yan6klMrhpBEOyEodFa8ZTbSMEjKDiaH8pn+pegdsqryCwhiU+GzDADNM
erwMrTNR5XBFwbmRRJNoWp89API5rxcmLC2LNjs3IpXu7G+rdl1jQwLeLFGVvng7FGelOZjLm3O0
X/Z9507LGGGjDVbxQ1yzOfd5miKsizaL9v5JMzMzQsHE/cUTb3P53W5z69Rq+B6iNlGjxz/WnTwI
jv1vyGrLgqW+ZXjwaZmJUU5Fi8u3AvmA+7A6tl9zzb5fEbrWvt8wsIRnigSUzk/3xFoMQFg/yZgF
4NlQh9Brs8Vt6DHcVHCdDn8IUihUPd9aybVQVfS9+W8ZjFspQdR1fuuTcE4rpNq/Ngdfiygec2lD
xLFeD8qrVNReHKzPoMhnNo/ZiCsgHEHXW1p3EAO5EgV9/xgJgaVLky8d20FkuwcymaydO67abIon
sQEM0MtWRFjqh8IfTi8e/ee9xkpvihjJdvzwJz2OMoRFb4UCY2EfkuEYskLPm0psiQeggoCnk3YI
0l16sSx7HKRx5L6UWkIupNMSJKIUF/4AJTvzwQv9nhBH9aCOQ02dw66iPZBVzoOlV+9fs423Jbnv
g3NTDdx60/C9ltgWo8E9t1rNwniqbhV/S+Pz2vRQbDoWZdjRMkrk7ymo4Be7dW3IuviFlC1WRxVQ
mctmmW0EydM/0Bg5CAHxtstptRI2Th5otFL/VH8DTR/ikREAfd7/X/WqIiHKe1oDEQTeAVfg5LNO
CyFl5kc0hmqxCfXtLbU6hFgO+d9bNGwrjL5k3cKn62K+47DcAF0nuFaI9cajsgf0oByoLgP8geJ5
jJfGw6Noqn/e4z/zHSE/7TCbFsxSSf1PicnLo7B3jK4KIM2qYv+usuMVjxWutWYAc3gK2YpwtW2H
XOUii1kYDmNPqH1FFaNi4gP6pvT6GczP9Pyaa8p4tllwpZYyDzFMaKBo+aFUJs1qkr57DFLDsnG+
zwjZEeX98Kuey+KblVDRzFN1xozH0VFDUmMblgDHVOyOZOfYPoDdtSysp8BbgR7u+u/LTa7eI1R1
j3nsaVUOOwohZnhK05eW5F+5fH4e55verMkwjc+13lP/bGixFsfG7HO0AK0c6NCQFsqgCB4Xtgn5
10EIs3G40JmN6VIWjKbjGeKRq5inCHCt5vokW4RzLvlZpmaXL3S+OpuoKNPj0dnnfzk4by0RqCEM
1GlxyvO/kaArOgB6DtOvWRXmBQ3UqA2FQdzy3IimxeeLgXrWbELFzvjFXyPrl+DhXFiLFbS9iimz
vVh9nOJX+NpfRC3Uw5u5NBsuTrH+mjuGpR4/aTy+DCa8pWChfBRFycmxs8mH4jzNL97dJd+MSTaa
jbmpkgLCus9b3VVJJ9GkzwA5XhQaSTnKWalGAoKnYs9JcVpgKmkJ5XHto3yZJt/X8lmQlmDc6+xi
odPcIYHIftTuN2+e5Y0GLphBeaZasKBhvd8CB2O1+X6CenbK3p73dA3GtgvP
`protect end_protected
