`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6256)
`protect data_block
R0MVZjhA4mJbCLIhMdymey0f6Eathtqn3xwC+YnxFZNj6KSXzxR8NnuWxgReV4ajzqGd2wLV4HPM
/XN+evwJw9gV2BZ7ufXmHjA7N0/qjhU3YlvHwOSU58uK/O+1alxi4vQ+eK/A42moOLtnCGmmvqGr
g3OsZG2GFDx1CXv4knCVn5WI98gC9pZbN+gMLD8KguONfgs/3Sb0epR9cAN8YOuXZVHYRbBEukMD
uErD+2EYsGHcvQhZcL2cJI5LipPw37nyBaGkpinxyAFFGNEBaH69K8NUumY6Pbshg136O60bqbL1
hugb75RajtSUuB0YiIwYQOrs5zRGiVSLrq5c3kUaQ1X4dKB264fdGHeInvVdI4PNhCSz4DOpJ6dc
Q98lzvJ8KjrIMjKSRWw+DXJEaLWKy5XP++O9tyh40ogqG9cb+i/AbfGAtW8Qz5xJ1cVSnvCKPb/c
bPxs+tKMS5panLKUoDyhvaNNyQzyoIAaxbdxuXyU8O0w2opxo0/2qf36xdrcZWfVyDQ368DkYB8t
na4yKE/w0/CIG+haSmk8c63djrC+z9HpwtlqtvLFZ9pOsFdSn0DWrXJjQSWYrp0ZpGiapPyq3CwR
aNlvNdcw983TLcYsjgA+d26So/wRx7tbUq1xX5d9Uoq5N7Qu/1EIasNZsuE3xF9y6m67bqRvDOWn
gyuKPp7SJCEwErmhE93iySW0+1RbKW2ivmzNQ65MrtrTjNk1Gh13QIsoXKAGFEcULD3PcQxP5NXM
WU0Ivm3UEyimZAmvVicRTK/8FRofuNxjpraR5bd9BMdbXCUpayK9BQv/ImNZUJVTZWQPGBXQ2Kvx
NWOJ+iCHqiONGhRgakCAcrHIWuCl08ZrMk6jOlJ1I9D5OKozZsCGEvww1E8fgxGYcfg+dDkFpwfc
ZTFjTtOCkvTUPmgKW59zm9f4Yc4sBFEUfnJsT+SYZWPX3narWF+Y4+ZIAjyni6VWgfEIMGmTppD8
X3G5WWa/Q+ubhR+KpmNvo9A9WVhZ5cyjtrwfW7XjQHr9AM9Bp93UJk3kcXk2N6Yfae8gFVCuAsKY
5F6tZWt6sIxhabQgAY76ol5jiY8Do+Mux2V2w5v7m8irfv8henkxqldmoNbBEwoJCxzysNWL4VJ4
qh20CU/HA6oU6Le2HTy8i+Nav9q+HjtgcKYsOD0o1DhZ/iBV1x8IATtPDAhms2ESndM7aN74Kvc0
TMPRuRR5XubGhTToySjUpZY+Nnzo2Pe9C9FGTsqgseSzBWdwXR2CGeUCRfqVkNShTh3caTiX/92H
sGJCqXUrhAuv18lfYqcDNIG0OTDNtLGbZyeUk2uEYwj2zmLEn2NL8D3UaSLGmsxaMOmyCpDhANS8
XiGC/LvBHNKgA35p6SnHXvQxLD+vtwaCEPGed1KEyNhuiBYTTYRmeZ+b4N8N7KVjstdpBG5o/qa6
YREn6Q6XcKSgxnOXXv63WvTvAOJGnOaXM0oD87ej3ChpfQCjvs5R9AzBSrWaa/ShIv4cFe6x1p8+
CqHuAIBTxn9fqDBtsoY0ISzy12dKEvwwjx7RYSEDOiPhZVEMAyxxNi5EbHTo7THm4Y9IYTtrOUo9
8Q0A6+jb6oJTo94M8EEdpGI2H+1YGA9IyuFq+VfaOHvcGZ8aR/DKI3mUiiZJEqandVoQX+uvHdA1
uURCXBPxnh87lEzM29QHD4Lpb7xH1rcm3Hmd4tt1cdP4l6pq2hEkXN6OYK9MKR8luNk/l2cciXLV
xSnsyMzzKZE3NGQ4135I7odBefizRNoCxpFZ0dfRrQ6dP+djp8TwNJ7Lb4eEFAt7wOWxX3xQKEiR
vV/Fv88vfm6/lsPdTHQGn1R7bXQ/R0O+Vh9fz8OocO7encWkT6AON9NxDZV8zWYXxgisIXNJ9cx8
z4Lfq4j6e/nAaUIQktL/zRqZz2r+gmYY81DyVbtiawmeIR36cXiIdOmKSNm8g/9ehOIxr82lyQWc
NXMth7iaHwbotTGJE0WZ7L5NGfQ85qAZBavYrgR4oTUrUGFnE2MsgKnxA4eW419S4XxlB02ZmGRz
R9iDLMWRHVs+OTABwhfYX+KCw+9aUL1F7OHTjwcrWgG3u5QfyIoz6vm/Pk079W1vmxsPHHB+HE/U
Yyjwh4YB0Jw77kgV9XvmpCv2sNCptyZPxtfN6Hbbh1yaTXGO0nM2GBHihuf50NrU5PxfJoVaL0YM
HcEFl4mihVtPG3qTT2p+xIrE97bLD/Pkx6z0p6XBZM/CxL9crCM/uoKQ40q1NAuHD/Jvs8ObVibH
MjjgWdyPpZ1S29L1Rtk2FksjCIhzSfv4pOjB7qVZpL0S76KcGVqw6OqYUIKS9I626/OV8YX8OwvD
fLCh3jbpdmK1boyAH4I1FLlCoWYT4FPgSUuGPvBjlqWJFgfI6AhVXeJHk0sbVD868b+Gn0GV3WvX
YvCswymF+rAN4a0+aYvyRAA9MSdU8Kudj7hT6XK7bqW468wCp8uPVwiIBzCP6InBvP2BoViOYtuI
AM9j+gLtG0aKLsi5DGfPucbUyGDErWgrczhxoD05idqu1EiiGea/vy8WUuhBx80IFlhXZ9GO0bYu
Selr/uqJkwKHjDWUrkDDudq+1xqoONRUzXWXK3ffRNWA4JOCYeGbK6EU7uQN+j6koAdqjkji82bK
iUWWNhEtx3i3Q/bXmy6aTAkfR7B8+K6tjXRyLHbE/wQGKhFuWrPtvoF/v8XsBzLaGc+2A6wIKhkB
Ds4UILmnHKEeLMKRYvGbmiB9ReWa5SLsKU2f90gIuJ2Am0m6TlvmjKZg1BUfx4UfGK1TZFituLzv
/WNqkbvLhfQ8D23vRmgkCg5vrg2YFJjV75xXz7wH6MNNfUShNfFGH1fEWGZsEEAVUaOcgFxKUbq3
d2ptuHjXRmvY+DOFVlwNPLDHh6l6RUib1aXyqnfwrCfWidNweJ3RDmlll4Kv4tu/fQnSVwO2sELu
GfLKQ8Nj8Dj4iaI0svzTkF+3s3AaT/vEWDxcPZpUtMv7OTUusTE1SLeoSDh6st5Wk0bW39L1n/z4
L7iN96co0DNvajK1SU/05a3GCyWYtcwgye5itQ2ZUNKktTg3omv+V0AzKkX9tpcJ4s2Nsk48UZho
ToAWo47QTXDK8A5jySgWszkwpsb+c3mEUQQ9UXb9I2wzr5MuVWboYlZ7AiNDOXXp7X9Se/or671l
HT3Kw0NvLLwHn+QouZJ60cecH5Rgn3AIp6unKtMcRStFHJuc4OTEpVkEmySrZfykK0rVHKLdAdFS
K6scqVz8JjI0eMC7l9t+FO/LmJCRBZAoB6D3uCpSs5mEqMmxfbZi6sSBn5R8LOXO1M+EuKc69csY
OJSe0GdWt4S7SQtxa/ITKUM8SPhjz9GFL7Otq/B/Dqln5qAVgnTLzqld0K+rzHpfUWWpdHGPKm6w
SzzQQmICMf4JD30w1idFL0/n/mULx/ITs/S6cuZHE62QDqjEBQawAbde3G/mb0iwFFLEFbulwiVa
N/qfJXIHOTedzJEn0kdGNl7tMNFm3Z9lUyXJVQ6CoSDJ9O97Y4y8uff3sLXiO67ewjMTwMqAD03m
LijM1awfeIJKLTHg3ByPP+2QiB35jU8CwGxXsOxeSPoMl0ERezgu6zFPadtxAbCeZBh4/MN6+UQA
cd6ntCVln3PShcZi4HkATHoLCvN3emv+S2nHLfwxAhoOlAo6UvuTib4NdUJNbhw4lg5wdZgq4AdN
MpaKuGhaMZejBNq/7YGCy7c2xI1RvxIyk3gmR2VhJnJyIFXZbUg/O150zeTuuj0YTVe4rfvCp4bU
H90W4kHp2FefLXX5PWLg+vA4dZrxsa0AAWt/+mB87QrQjEkLsSoyOtoIWpHyFt5lS6widHr2y6+q
5B4QgmOttTApz2fhyTxYJyQkFWpF6f935v89KbdMThZk8JgbOUW3JpWXB9FRK65/MgdyWxmqo2vv
/y5rCV1yf+1EuK/aJ7qtGDkfmNAEHBIya8B2fDpG4V2wJTbvYW8JmnnqCkgZ8It9Fr6fAQ3qoNty
J5dAPSCg4q3GolJj5aM40KJUeyJQTkSI2lSmJhSYxGZ1OtvpBqKN1e4ygeVW0X4l72gw3pe0QnlE
XlMTT6P0UeProxx2uYI48neO+zR0kcPC4xQkKMSbyIIYFd41jEV0FFxStpexDaChRd/3DL/Sk5HU
huhHZD1B9++YE3qCM+o5fixcYxkojxJRQSNU8ZGILu3qPpaJSHGk2TCTPW0+bSEZfDb/DsKLqJH1
/CjxK2ohoxtttonuhrk/zc71AX8Wpf8Z0oObUlWl/QEHnK1vajCVcAXKQdCOHaXpHOmTbMBpHl8A
X49fEbIU+60JS1JqBDthApA/1i7bCGZTd9wAzGeNk0djYYZRnwN4uEfHMMO3D7HCn9wUBxBZw5ga
omsV0+yur6j0llefBfBe5ED6Bv6vDbPLXV0v93eefCjfWZ1bbCUzFn3teM4diiJnkIIBo2BbsYg9
0gvrLRY2OFTzwk7YGdJH4hWYiHg98ve4OtmjwF+ra3F+e64hvRFh4Tzlh3edLNd8X3ptfq4DRqc3
rhgJGUsvpbBq3cmEmBMWS4sTGgVR9TjDdUCe3KXR/ihek/GWqtK0BgFgBSXx3Gw0fKayI3b+i3R4
DbbGIs3BEBbeHGO/7CYDrIsvNeR9RvtRuCGK+fLls2KL9opWVKRgwvodsnAxGtVcfS+pIw5YhWrj
rAZ6hW5IhAs20v0GOhCkG8yJWpN6Vxm5NqC2qfS/L4YUEiqK8X6Dzg5OGRb8NhWFU9xoaIiYib5B
oaE86OcWBbhLpHBnjci6Evca/slJ9OdhhzPyK1h/vNtR42W3J8d/+dtVsGt8o/J24Ht49QHdgBul
6F8+bpod2mpfDcuWCv13upE7GZ6j4RWSGq5+G2KcODD4bkK8e7yzIlpI/N+RcxY4cunaR6UIp2p6
DDxbZ5YWthDcp51LS93F7KPTAlQYXwgmNcDXhStTuAEYspfefgceL6r14Dp2Za6udpRimGwnL9bD
ot3dAq/FQVrtCtRwMTpLvMfQaeQBwxzio5gLkzONbeSjM4+QUiwjuE2ek+23B516hwpy9brJrVxS
L/Ez/GRPw1k/N0JiyyD5pEscaLBvwYnhNwORbmNcQ7Uv5e3NgE9axcj3iaE3ibLTULNnQTxu92vW
gXAaxFZV6RIU/sfTPlRbTIlaCKTTqcO8gGBfaMXFq/U0m2V93/NRWulGbt7hjB+ydY1moe89OpCz
ycaqehCQSwRs+bJZv4iPmGQSvmnwG4emwNfMsoKyOofegkGbsm1KRKqnW54dhL8zJdlG7GygmrXN
+pRrwO/lrhP62Yi4WH2wXKaajAd3mjiCXnfafLnYUzbm+2VuaGYz070WdnYs08YuwfVIoz3P/tvg
UP0mIKq4xkZK5rt3FoqaBekDMssNFhcpYsm1J1vi0CWABpSmTVs6JXzneTvTjehJFn7OCroNWboV
sxVsKxG6VYGAkoaBdnzzrPn+ufLPgf/sbAfNYC98YM0W0MAaflLzGcsIRknv3VxN5mB+eh33/rCo
RQSIKOFJS0kNwV1KxUsp2ZNfUrZMAXYvgMSwTjxYUTqOWUco30IA++ODrDQ6cDyTlUV7xf+/qMW7
b0OctPYicv1fE/P4BQxlk4eAQLaEAGgLlMGryrNIa46Qsn0L5+8Hd9Nx61Q0L4J8SLA3rcgNs5BW
gCLM8c3rx6VClkSVFno/tiYnGVKc0q6foBay1DkNd96gtkRo9hDog3B2qTP6Cf4zh2Z3EJklnOXI
9qr0+dRr3kMsamLf1ItTetZPjZf3gvW/5YEzG5gdFEXZrCfo5JcloaihwQTWenWuot61588cfLTn
O1s0sImWP6wU0KZ7/cy1u4VxUbumRDBCfvHKc04q/FvTydd+qPOXgHVOKMyINA5dVR5pNPo1Fhki
tEh/e8fAmtUi4R7H4nY+Lq0TqrONzg4d8O2O9s13LpOYBiuxS3/UOKv9a0F6KHZ4xEo6Hx89DS89
5NMYVtgX0RAcii7NicD4IFwglWl2CJwolJdE451ECctenTEYroqHHz5DPcheRISEloN1HohYMi0i
Z4/Z+icKPTVxcIKLiRDGhAVPu6ix7Ycd+X4dCAyefhkU+BJYcZkwdUjDcfwCmsJef8TeYfuf94XN
qOYY6KPTW03oQak4ipLWPPoBOuMc7tiMO3j6vJCmI2k3NoIMm2V7kCMDE0gg2fXurO1kX/BuroxA
JUNgPaxIzac4QOSBpO2rV5pevecmE2z2vNAeuSSDtEHfwRpwnMJRoEEPOyVY3N0z93TK8qQP6Tyv
JOvz21BIL2l4Hd9AdvCV6PvNhuafWvWLJCfpa1JRk6GknE8ORkcceS6eItFxxW1Hbs09hONmxWAk
xA132or5c5Wlbc7A2yk+/qZXr6pOLZQ7BaMjfHbSnCNEWopvBiZ0HsGayVc9aE/0MBZ0Al6t94pr
nl5CpsxJmZVO6DyDvFLLpQnQo2TUAh5+KCkUPPHcSuqgy2rmS7/wCJJEvO4Lbn3wsJv+pVPGvvrZ
p6GPhAyeUNoUZA7Vk3nBTDxGRySiTD635H0V8hlYFULi0XOTvcbiTcUCHbU297t1Ga63hws4sERG
PKTFV0okFIZoGF3539Nyb2REAHK0Xk/B1shJTxmimYbqgNT/jGcmHo15zs31TPnrXh01CYqF3AUC
rgfMVfxFy9blVzOCJqLrwecQX7uzYp10gxf93QCQ9/nmOrTR3fqqg7y673W+ewlJA4Hm9462TJ0f
7m3fBoVVJ5Yv6oGvVVlpb6hI2D4tk+SlK8MrOalln5SEJcIwCwxBMbMhNFJw5XfSyBH/qv6y4DM9
c/Pis6i2b2YZTm7f2HSL6NBHNomJQ339WY1NYk72F6ArOroH6jMI1GPVON0i6DhWYuw+4PtqPH5v
UzHI71c4B4kUAZZF745nOQHOCaxkTj+5v1FYTLHwawCW7bcCJ7Sf/h9Bxl7AA+M1RNZ2idw3dMOh
72ZHpyvAu8VFI5aDgxBqALMw+8BopnHivrOG1dFuqSk2YbTXL+NIiajjCaiwkrFAgk7ZBxofxdYm
eoyPoDmYu4bIfOHFSe4zsmez7UubRzjSRCqFbTE6eT/GOZnxYA0RJ3sZS2XYEPRKUtyc/2cmCPkV
4sr7T06FhTQLSRO53fI9N/2l26itssDRLZKsrj42BOq3/RNOGgP0gVu2mivbb8eAoxMw0SZYe0JB
n86Mv3oc74UBbgHXVY8UdWtL8vHNg5khxX2MitOua2UDsMGV/q/31/NYV+yLroCF6Om+XBiflE4p
Lbh4KaC28tnpy26d+cRXQJJvW0WW9+TRbhr7vwyWEFn9SkfPBsjo9PSnCXr+Np7hW2P7tAur7fGl
Pnol3/zFFTpVj6dVEepBoxzUC9BSK0lIDG0aiLtShtmf2J1iNvuJNYMKl9v0NXVaWmC9KO16PR0r
Zv2xuqSgJklrurW7Gq8335ks2/59oicFj5LOi+K2UdD2isHRRpIM3mzrNXuk6JLyRurpKtY7gjtM
31sZh0doXVYoVhs8WCIkSjfqtbNQILVQuckuep5L3eo2sKe4cVdR4Dc2dcaXhoLDY4lFNhhzNJMP
d/Z2e/rfk4k2ZrbrI58qpct8b8zkCqlfRHGQKas7iaWLFFc9XZsK224h0XSPQrdL+crKrUOpgJJx
9CsFkUQk/b0GtNrd2q/fT+5/pIdr3+7skdkPPSOO2OBvxjBs7GRa5McVQgQafy/t47X3HEZ18uZS
HvUOcLMi9jHRWrGIpMs/TLIU//rTFGT8VcGecPcgeblACRngOquliDuTNaKe+bRk4i8gnA9rSmVB
93fVKNsQ466mVvcULBpMK5yDMv/WuT5ca6seM00+OTauiia6BsQo8JJRNjVBteSndYt+wj+EfJT1
bVntMkA60Cmoyk97f8yG1xvfmRE2CcQfUv+D19LSCekINuKtfjJFcE13qXDM5b4KJXEAECm5/Oir
/O+roNd+mATy9p7beCdnVDvdaQs2bpwQ4I0gpUI0fKfwRcKdmePkgX07QRND99plsC2rqEx2/1XH
9mnqCVm9kte6HW7u8dao+QY0DlIMv4eMETn1SkRhhTgKfRDS68EOwLvAkUT+I2KxPPkesrAUVaSe
4SkZlR1/XkHRM9TiqfOzdeqdPWqLzcpzlExN3vW4FGNeANHURM7renqBo+ztu0M9oN2hk89RGq4t
bIXAQKSJMkpyVH2eQJdROJ6koqdjVlIcSuG6jGjhF9NzBuU+YHrsIi2bmV/Iw5co5TfRBC1lvR9R
iMKwbAaUbVs7s/A/S5pD5uaf0YC1gL2g3OkdwYPu7YeNa4CbOts3MovLpA==
`protect end_protected
