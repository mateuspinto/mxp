`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11152)
`protect data_block
0USWSUGxovGsyBJteYpEoToHr/CT2JwYb3pHYbg+Umt4b4ifnt/Cn/EoNBEIcVXX6Zr/gD640HLf
ezCKYqkuWLluNKSlidQDajt9p69M78Ll2BZaOrB+PZMg3a2kkuezl8eam1mkbtlI+cvQ9q5uN5Mo
TXUoW9xCLXnz7gE+xmrTvpwj5D2UJMmB0zzuuP1T/B1gNLiPWJPglS8PWKy+5Yb2+rl0EE/z5zvO
6NS8rSNs2VH30sJkxpbDIqBGTB+arpRhNUcQTtzOLpyogl3RwLos9l2CiWwdWu6qTFsOj9VVg1zq
dP0h7xxAcfQiMo4Rx0/rFMb+eaioooimFtaJndKhZxx1NZQlxLLvVcH9X4Vky4bqHwCnFW5HRTsz
JQ6jglt4mCDP1VH7ZpGcIpFFwTEWIxJ6zQT7udaE0OriO7zHqbdfK+M2pFv0DGrcnoPles5bP6oB
YIFloseCrQtASfXJrFCrcIVmIYrBEV7WU1oc19RqpfMyl2GDvFY1E+Ot/SRFKRDNYUTtSpj/bYCc
QO/WWfVGxm/nO5Ofyl/lVTM4LU7vjuin4YPjBn9qo97MyvPmiHhRjl1fY5AV/u1o085PItyffU3m
BZxf1p7md7tR87H53KGm4NRpIOqhQSchCU+FStSBmRFl5qgurlHqZIHmeiVp/ZNi/b2ZgVy6U/Pa
ZUKMSWrcAkybdr2kVzprw93os8yd0RX6ZjnPBQwngulrt4iumkQ+ZpxEEeieSlPpUh+ePVv0pbof
LQB/5189OZ/lt+4CBXYmCHgmrIfC2DExOPY4CE1yvSAYfS/571B2d65lh07/+rvd8dmYPVEH4eKP
oqaxQzXyL6TEsBiqbKEd6HiOneQ98LZUgL53DCI86ar4oVjSk8kipQ/RIoIKcvW6c/EIz/rCOYB4
qYS6/ImtViQ8/9m9B19QjHF1Iptx9WqJ2Rt+jj9DD0w5vMUtEOdYp5P034dzeQ/eYelGzgh+lhTA
ElJ3hNiM5i7d5HAo0ekbw6JrjwsLi5b6kMm2Av1b3E7hhUfTSd8ekIZXeHh+Q1FXfOntbgszzatd
IKhK71uiBiAXmvS/scRe8+ZktfTOzFa4w5lbHmuOCxyHgXWkTEfhMGoCsLZPxk7/BHEwXWLTJDRH
ynP9fHpguBWqfpQdoLl6Gj1e4fVqEwYD9b86DQ9r/2jXmO9PhjrePvb4S22Lu1xofsNudd6bdxnZ
r3PjuHapL/DHu0hS8fT0xamn6Y72MJ6Bw6bPLltFeKPkcQmwOwKDylFB8fHnPxKXZ4hrr7jhvQiO
Sca2wTXRIzJnQ3JX/+8aa7VxjGrHSs2pj/RfwksZpmewBieT2VFcPuDlfV1dVrtYxP2g+fgiizlc
lDgdBWC7sgmbGWyiEEoOKgRwMDXX1+I1WAPL/kwHRVn0ejaz7L5PKcbcDzPR8h3ko6yJByKbI19d
T1BMQinYCwqa+t+6ch/o8Ar7R7ymN1CW5/r3e7let41uDWkzRgGasqmNla4S3xMT2i5dpPpn/BDu
UyvxwmGz6qrXAkc3UIqHtqDvQ2A1WlXOY9OiMCcwEX+D0wOrsnjGxrkH4aJ+srDGLO6Rg1OYDStx
VlJX9wQhwzE7htaC4rQ55YSW6Glv755v5UjZnNsA2vt3r2J83PaDVtU/TeZ7B0SG+1L3Zla43iuA
Q5xU6IDEJkbHvDTQCLKdjNr5eBxyY7oMw684/DGstBSEt3fjgcHkf/3f7KMFesJuDThNfk6WnzP3
I6e90fDbgfmaFgzltTo3UGvH0aoAAPEG67uXwNc/czLo6M6tJdE1Z9H+3GR9XQTFfaHeBqy/Lzer
3JiZv3lFuDgXCo8cwC1sNAEckOO9J4Gl1IDmU91HDglobLLIeL7E7fsZTLejz8v1RUjCnANNN+Ub
weo3beTCsSZY5kl55QXhrIhQmfyutcBYzL+lCeNTzS5k46dE30UTR5970oj0F20TQSNE9FXizfSB
B0+FoMhA5WVecwewT4Z3m4umxp0l5r7Q6rpwnoNr5R0BffDR4eQpMDz406Z1GnaTnH21wdAsZJWg
rxg1v//pIAf85dJ6SCMH4Fs5C2bEBPi4QcHxDX6OsvlofSreRAX7SYLmwXDZezzxvRtLnZGtbA3a
0EszSy24wHh98Fv5wX9m3W8VAg+7MPDW3fAbWMwz4420KTGxGO244guZrv/bqZw6EbYM4wg5AOBL
pLr4YnoxHC6hTmOJb81aSmTnvt77Jg/ZrBepXLv4SaQ16+fyJaZNU21Spdp1WLCNWSWNKnJBzGQW
8wBPH6uO9id+EY1X9DgYpoBPTwPjgoxFgFzHwRsjoHL3muBhVyVHJQmWjRENjh7hBok8ZuyBX1gi
a42RADHSx/rUN3HGNdixg4SfwPwcUO1oT3cAOPkhfCTx43xRsqZIPwrTSntzGFtSn1g+/K4LQ0Mp
2aNzsqEYIWosxjWZi8OGZ3EPVW0NUHpL2ZJMrlCqmyNOLDzZl+gxS/lRVK8jRhmjr9C6NZvgHuAA
fU5YFMM0UEFYq2rRs/4STZZyUX3B2MyLjD8bKpMiNuoqRxC12kbRnjw4maLpw79+x+XiMYPRnXUH
TyG6PX0GuKT9oHvfEm5SUxHHdFaFlxu4//xj+8hVFdLDig5QvqDnpEfQxL2xUeSPtl+ZE7vZyC2h
VVNDRTG7lVBT3kpxZ7p36ytjqnZjmAlk21Psw2tBV66m25uLMEAulDZ8CIAaWl6BbaFgScInPjWi
7q0Yp+Po0gsL9DwfQAZYuaOZPMAgfrpbILUBY0riS87DLs2eVzs6Frztpz6VdG/mwB+uwCvWl7uU
a0YJzTD4YJOTdkWQ212oydu0q3jCGjZ04LQnRzUPqGeqTDqxqcY8yjBUsme5izur6GWk87JnMvu8
4Xl880aFnxJ/SyiV5N4fiJoGbGpZ2fiC5D1dhNSQVaHN+ef5U6vcMvrM6ZWlzvmhXq9SOMatNN/T
aOXMil0k1Kl5fmuHSB6DF5JJqcv4mHSGaPZ8sgcZ8iwBKQGVpf3PfHZ54hICmUmvsTW9ZcnEftmV
FOBEtm3rKQ7FtCWiHZh/hd9f3J6IHtzAlVERcgOuKRKqJ6Ru0lC5NUQV7yXyuCo53UJJltFz/RbC
Ti2p8DJ/Ewn2bGWmqDQ5x3ITInRQmlrQ7jUYuv4t6xBtXkDMg+3rKdyxDGBC5mQw6dYjgkiXMP7L
rMHrKEg8vKdDtgfrczes2ueJPi+f67wWqjarnrusQbY3mTyUOo20hrppOGGvKQCK3nqQbdDZmT3N
oNiZJbYEums0bpmFXCHZnBFMQDqJ4qIphXoUsNzAA0eTNZufDJrIb3sTOMXkHjBQWd832UpU6CGh
S7BgXdGk2z0BFHUdgTNSeaX+HlYS6NCUatZ/iOBpQr1ViqnCsaQNuIZUlQQ+6JHCsfoFVaTuXWLq
ZDO7co4ekICd0vq5mza8M9e7iODBXJdeLfPmz/GsuD16UmGK6jnXPixPB6rSI0+2wu/KvnhHoziU
7hF1Ew5itOQ9HqLo++zoC4UEXKHMBiUkiFI8PJb8t4WmHzeWhoh4By7fw/3SoSiWvyc0CFHGNAgX
vc5Nh6sr+3Cmw4K+5skO2ciTggQbjFpoZNdjezGC4r6iVWLalwxWvj9FdimrKH9k1QTBU8L02ED2
NIQewTY/xzUKAE0VBcyGyyxBwSu6x6NCL/4Et8Sp9l66FEtRYivYuxRGg+7eawJLzy5+dWiD1NGE
hH1j9PCA1vWyHD3UyuPr8yuH5vqJ0uviPJnWBFNo4fJ4CvLw90RPoONN59LE/YL1naqY/GnbkUVE
9MRGdlZRTh22IzdeA625cDcmzf+PwL5+3NefDb+kJ48dMNlgWehLl5hU5KniLhxHrWFJxJXsKgB4
0zZAWB7avIdOu0uIkq5zYuQS1C788LD7EikH66/y4olw79TjDZ98fyDRqm7+dSdfSy1PVPlMoRfo
i7K1xOivqQdCAsvtw3CaNj9wgequA/IKpkwjMp98BWdgJDIqB5NJOIJf1b+A4iOVWrIf/vxM+ySn
BHl4k197Dt/Hd17U3NPsVhsoHz2s61vo2bhO2ds0KWIy5VE/DVjLtwC03OO4/EOqBgjRtyL3axF9
uPRAAdCYtUzD+Lem1tKkfLonIaDWig2hwflawFjQcYcalrP1vLY5rDmCGvPEGhPJIA6rgeKKFpbr
f1GD+idC+fkWzQFW5d/z+aErIgQPA4G6CYPbtu0fmy5gg5vEV4glbPaZ0GKeT7wGSbVxZmId53xf
r2dbcqVu7+XmPl+joTYbWeQRMuudG1wJ/js4hSSoBBBk54OuPBABONcccmt2RoaISbzk53Bcy+rA
S7+zVzAKEzc0jVuUdQLOFgv0QeCkMx98/6n2GA+MgXFN4eAkfbIG/N4QCK7tXh+MctKiaDeqwmtt
WDrfT1x63sHldsVdKOiatBnpb5Jll+9/mYsomYDNFDBSk4I14cGlTET3VSTwqSQGogSfxHeMWnlm
JdikkD+pRAFhbQlnWbuk6ukIZg9VK0sw7cVVKFo9hsRFxWUrKAKcqRsHNnuuHiybTq/jcwt1cp1O
CSgeiJNc0LtP5/8wc1GXD10rLDo/CogxpjxdB/NiXKqDU/RpYXAPoIBv/Qsus+agClK5MVDqEs/0
0wsAvrH8fuTrluhph9hWAWbox1oVwYxwYpQaH0ZzzC+KFrsj1UIIaWyotQgQnrQ+BLhMg21EPCQM
cx2ybAVHoNNkJ5/ARMr0Y9eWFFHh1yOlE46KzG7U1HKDW3D0vDehnK38RC8LoI1khQ+ghYmzKcdK
qo/xKanmXNBQHLnZuSWAgxy/GuYHRNGeX23wQYqOUKJjjCextbCDMyHe5axTTdOkOz0PLXg57PBw
pd8YC28vL7u+hZpSxPJJH0xvt4EpdRCnTo1+2Xs1FKFtjTqgO5qUDndt4rS5IFgy/onRey4t4sPU
pkJDchlCbfvWFV7Ss/JmoXRCLgGQ+v0waXsMQ+gmjqbg5GjYUzuIZzqseyDjmGlqkhj0moJHn80R
mS8nPPtczIb/vUjubwgT8c1UQgBa1h6MAT7k9+cDPCdwU+/RLUy6ELe+G323U9pW0nga45ZYqT8e
UUv13r8m9ZnHLEezjtMCsWVnErEMly9jswqUgwafVe6b/NCQj/4vcH2iCXUQqvSKcvchE+0whlNy
rzfxXh/Y1Mi3i/MbNRoxAVjiunHlp9iM7iBw1SBXFAqcW4awxczO21L2tQKIf58nNnHvQ1vyw1bf
e/7P56DhvI3L2Xo3OvJ/IaQCgrX2mnavjDSJJdanNDACK94fZSr0wA9SHEPhSJhSckX5rjb4Z7bJ
nYB+bli2RbK6rdmBj0/nyIunyjJNJ5sIxuZb1bSO8kI9uYOpiRiVo3EswW1+HNLzAhtTbZL4zbXf
8XExh3ONtVMPj7cvZdM2LHIqPqrOuH0qKRQ85+3cif4PPeom5hLEraOQm2Tk8unvpHRRcxOHB6Ti
itnMFsCChCxrCZJnMvMVX79/PEUbIG/8lVkEphGRVaQVItE0L++J26M+97v1N7Jl0x9KwS5ZBTcs
YqX9oafzWpUOlGcHKef97o8IFtlQFgc40A5FQ8IBYOAEfwPfe6LBcM2tTv1Y4gMGBk+nHtjrl4Dk
7BbOa/d19cT2b6Dl8DNdF1gCOQGdJJYQrO1ouf72gxTwA9KqF0fJItmMPyLj+7LRn+/obMkirpbf
Rg56ztKE/JulEZ17vTzMovpFcCPoA6IMpMO0gQ/etZKK6iWlOO22w0WxW797hDq7jS46gB/yykXF
t5YWLS+PZ33g7kZ7O0VE/2P+OUBBvkMQiT7VwM2ennvg/HoaW1LARFPkrU6/GQDdbulA2l1KcN/t
gOoWu2rwBDcdjjPB55/0Vszd+eW5dtx2aefLdJpdJHmtriYz+jLqDekfyrZ1BuU6TktVXD6EP8hK
yv/DQtKACVC97B0JfmBRRS6D1B8CmEayzt6AHxRnOwrjILNVdFqgwI3KOB3nZkc0HEc1mFkBO6rP
I30+cWr4L6NnTeFU8QIUQI0cnY24h+QAKvc15E5gsoiInnTP1HSeyC3rgoITvUkVzQWBY46XttOt
0ZOLvM3efzSTxqimwtoLOTwiXXYIHsRPvariEpm9Lt3HATsk6xrZb+Dl/QE+d2WJspZnys++sSJG
RzLWJAxjVQmZem11adowo73+7D9QNTYwAu5R8ETW4HzKDwaY2Kt5jck3d3EXDB+uRt5glXUtyMEV
PvUSVSjw9gS0g1R0ltogTVWO9EOH1gGujKdb+QOEGj6M73QVY5bYdZl+4Qd4rUlCijBjuVOytF3e
FBAr0EvXxqDWSs+gkPfaTjgSfKLe/C7HPozQCYZBFctTCcnodnl2SFMuhghKs6gNTtIEeIg7B2D5
JFYUMfIvfJ6hP6FuG3hK8X120ocdLBdR44AcBKUhdXGJ7lseZ/kBGvtw7+Mhwq0kjNj8isQTn83W
KriVDklrZAFPMJi2OL8qadGnYTQ5GXgWHLgQ46nEw9aSpuA+BM3gjVLFDm0szXbJfFyntrkAmNu+
iYWamVQgowqwtUoQuVBB6guNynJ5u1+N39n8FHnY95sOKanDaOqdjIxRiu5iTo90Gp2dYD6AsQB5
ekFdKaEqHkx3BDTwBRwSVtL/Z5rLuxJ9hUfS4BT/eFmdKV8rS71QqSmkXexRvMM4ygzNNLOaFydg
+mNoGPsYY4ieHr/TrLdOK49fZoiSMdHsHwcsFkveS4gDnsaFiba2tq+X56hJYAbuUYFqiO+MPHjY
8q29qOqlGAhqz3oBApm+T0zE5s1APK0yRrIUNuOogj907lqPm2ahMnA+Ahq2wteL8CQu/45y7W1T
1PAVcBwQ2JnDUYPwWD82224jGAk8F9fkTFLsRsMBiEnMBxrBf+PArVv/CPoeF90nySWRt34wLvy2
A4iBZDDJg/K7uMhaLWghmwNx096zY2dI97oc0eEWUP6sZ1BJhgi6lLfhPmRKuTMjq8q1tIRmqlMV
y4ppylZlZAYTo5ysQgqc8krvdpLwrm3GW/ZgQ06CG1iiuIQ756iAJAFNVaIQS/ApE22VP63AiWEt
vhV4EpcD0NxfrszB4EPvXt4lk7eQfs1Kz25YsTwFSiyFMCksmWKBFhVVvuCkPhnKQqCtsK/wyTm1
V6+hJ8ep+eZxM5kn0nPHLjfaJhKIsKca/LYVMbFcu33u+TLW1tTk8FK0oskt1Dm/rl3R4enAr5c1
qp6UMM5T+HKcMcpuS8SUO7u1guWQEC6FIiTPRM7enLMsCFGbmKyiDhyGahDTjHc0O4BAGm/nkYGx
1TnvrpYRXDPWATGgPaIy2HxKRUg5bZkrFacAgdqA6jocCEWGwigudXigJ7AlEX+hiIZWvJ6uoz6Q
RVL9ho2lKmmHoNjgLlBltiNrtJxWKiCz5YdZRND6QszDJd0WuNRHfBgStACcVHRIDfgJ8pyyzqJD
ohOLHETjfzgTKK919pjMzyeCZTJaO4HepXqFd0lwbqMC8QTG6vy4VbRp506nQxyAKeUILJJOKoUm
EDmiy8AZfeSGeYUEztBcr1rzeGo25Qpfh0bOvzVyjLN2gpSGtZkQfzEyKpERk6OlBYwrEpVqBXU/
lMIkRaIp5R4W8rG+3si+atWLZfOWvGXOvMxMm7jNw37LIOKXYAc1zvuE6fKmLGi9MmwA2Ci5xPvJ
sbUUmm6yhz8EQYaAhWm6KrVt2uX31sr2IlzLUyJ7jfhKqbt65j9rwGzLTQ0RSvp+PKpNbHD7iiio
lZh5RDe2uFiqpnCUIGzZTK43bHzreVXoPOnZJCaQB1xUOgkygNjfM/gsjPVva6cdIbWUu3mMHFJ2
4iB59usAao9iF7RZi7mwWCDRIubz8yYXcdK0e75tyMqE43yHu2MP63A8J9HqJgiRQvh2jSAe9Hv0
b/10Vq788xze+mqAs7xyFFQLF4lMbQbyMS+ss85DWu3o7HNVCZcpqODzqZXxChfeoMJdlb9b1j2/
aTjVjHel8gnKDk/OumikZfNNzxjA3lvkGqfrAf8UK7xozK6KjsCnixnrLOkLn3hzwFLCspAE3HQb
F4Md12Yj9wKJ5Cd4W5ArT2jbUP3nkUgVaSxSvm85HwHENojrZbZY2kTygZUU4Olj5mG79cSxYnyh
ZpcsQDMhrF8FAMX8sP/wbd1nRZ+iKmgS6okU7NFX9eLDS+DQPdrfg6yFkAgnyYw9j/WGzK9uYhKe
1h3j1keLC1VGfoxq5wq1an+wOBx94S60H9GEpHQN6ikNgIKlBb9+I++nn18nfSeMNYv31eykf7Bt
4a+zMbTA4PKteUzpGH8gJLvsg3B/cQeF63A3bZbyydi/HWg7ZJKSobOsAlGRE029qZIfKfyl/AHB
PykaJ/Ka1E37uTzBOYGuyvnbpL4H7LnhIQ8k1Fml1TfaqQW+LUX3gGIq1q9vTP+Kqb+Jki3Pns5y
fblr4UeZVJxD4wLRvxXLfAL/VujPdvVxCXFBL3uVNqCofjXcmUICPajC9F+RRI+z3ZBkihKuWkKZ
C3V4VUIfG4Jj4sJmcxeyWmsg5NgznobqyIz/AjorjsSiuLEzRrWD7ZdU4d40gr/Bg0MJpvu+KRz4
xggHRoyiVJqSHdUkkxfNR90G9RTUDgVMEv41DkKFo2Mpei+rKEf4ExW/JaktYu9j54PWTf0oA0lu
CCxoUgNTY+IfoHpIYNacb9r5lnmOziXzEZoFUE0srU7SrRkW4o/90s9aDmwcNzetOp4Ai9kUSsao
pj4Mk24wLL+6X2UZHeaYNHjg1lCfTkBeO7S7kn5nGdAyXTODYIpndR+CaYMnb0VJVT5QYLFybQT4
FNC2G2VbN8bTcxG870xBsXmoVS43f9Z45YbaXv/zMUwWMGVxzh2+PQt+OmOK66Ofk0kIpuE6WacB
q5qysdNn81w9gT2Ym9qKoUCj34GJQJkpoqLJDSu8iQlKMkJByfs1fIcWHgopVd9pArp9J2Cep4gV
9QWuaDpInZpVJGZ2Hd/e8FdHVfRqXchZeJ7M9IDjOgiWsfPliv5sodi8VRxaYAO5lvKJOqEf2wqC
U4eIPsTYHImMA2nt5VFWDSiv/fNoa+QLwqXxfJcBsohWlHumnXhmlPiLdCyszxzTZhXOmPwDO6yL
GNh7kEqbIY9yxnhz/itUE5n36ci9SF6SDGhGJ19Ip8QRfS9go0Pyz6GJUbQuvoL8X1omgNmYKaSY
YTWlrPek+8ad1v/ywt0iaR1R4vTuEC7sqfMWCM9gEALhPVZplazwTUaJ63AyfNjyuQAbe+25dQgt
OYKWOcCRKnZh4LPVCETvIBLFruAc5YYaIejaMYD6ZOoalj6nskyld4jEDWtiiTkpaRpz5pIB9lnZ
dpUmgkf93W4xBnRKYYEJ9tkLTUHdPrZHY8MDDOhNefJ1/FSaqxpswPb/Q7z03vVlqqs36HwSOwh9
KS5AKVWEYd5TVGzP4rBU2IR+qWN5XDrBXGAISKKnwrG+WKaa3RM7RZsqPLUeOG4k0e69+W/TDIDC
AiGeMrIDNxeHy+/PS3DscMQwLfU3wZDFcnXVmYZgM9lG1e8UKnVLvOngMSKSXnJ4BElaq+A1r2I2
zQjMDisY9143f0codQW4S+xQN0lvUePlfiXNIhicL+oSO2/zZ7JYKx6ojiWQYjEPnQhxxGO0OZBg
ZQ6o7AtD0YDl34woWdwyYFCddJdBiaghjD+gIqSMvM43ELUfgitW264rG6LvM+z9s0OFbVWrAmRv
HqWQI6dPkhiy7Az2GMGx/WJ983ExhwsMI7e+6ingC55smH++uxqstUjXeFEfzFrPA+tGIOIxhgGh
Isqse2//x3fRgFH8FnajSGQ9ZEAtzdxbrqyrepoDM8aH2JGTK7yro5IHoAxMv2z8qY7FAqOJo/FA
ArPZFjx0/Fdvi+p1/VYA6297ac05ZaBE/CUl/iLvB7e9TgqV6BOPF8cQdQ5eyPuEqNMkw3zWxtin
nH4UEzTLu66oLRC3FbPDovmYPflSshI1CdMQ8KdlnhPUxa5JIsdCeDzRjv0/upFdM8YH5n8uN6eH
rdmABX2zTkB45tQO7WtiUI55prEnc0xLLEdHvin4mmLr9J/llFl6qsOFEtxxgYNkTiVkVsF1weAX
r0iNUqLmnTaXbLsSYhYvaOJoCez/kw++xMiuYxdMLKC2eNfy5lvpWgKN7r+NIfTEQ+NyF/hljsZn
Ig+x1POzZz9NNYINbiGMZ1bPCBII4T4S5PRsRDwhg2I01anx77n1Nl+P99hMxBiioR3meqwV2Y/J
SdlXZyuqcO/qyYe1o4/xgrsPxTt4AHJjvYh+VPa521Fj3y2w1L4XhARm0/OmiZSc/x0ULkKj17+g
vEfFT9PpbWEMrl45P3QRnYjZwC3RntmKTF8FYBgyatSZ0O8mq6OgAqjJ6XBs8NnWgIhZANfJMC8j
mXCheyZOUTjXX5lkYu4rrSh6CVj+VInJMT7t9Bpu1jYXbY0fTJQ9YGnJCsfmj0vDPvaFq3x7zOYC
cFX6+/YMoU66BgtFgMiVGTjVWVRu1VOkwDZaiAeo3d+T2VKEPmu4CPYOe3csMbyV/E3fs+OFvrVl
Ybig3fJHMP3Do3HxDntxXFjHfMD7tbOezq+OfcKVbbJlAdi3IF/FPKyKqI8NmL8RO1cJIfosvujY
zwpANxxDkkMhs5D+2qsgcMlj7i4bwYe4VEZNU8DXGfJb1RrAeEQyeIaaeZJz2JPe00I9F6H62ZUO
c8pq4t8iMUSPXbN63n0s4vbDhyqxFIqyNVrqcNDQOr6sb903Eadc3nl1sHkkFdNh1VCrI5XilklK
4F2e6wFzjrdSWzmtj7xvkLnn22KnqiWZMdXkhhrm0/qI9tUFyEOXf+0F0sK3PGCiNNgGh4dbmeMb
DZGphp8Matp9KizCQXrIVML41VE/CLG7+/gq4llqB0d5ClrXsMpSSmzSKtBTPmdC+OieSAuKkB4x
17pqOldKY21GPgqAzl4K/2Z5iNg7okrToAdVasdw6SIWLKt8hiE5du6oxzz88/jUgJZd+FMKBSvS
bSYRgZV0NOeKovO/nMrGeJVTaq9fdJhTOVwBCYOnA4Tty8Vt8breWjsnI8CbWK1szLpnZgp9aI9+
RmP6u/iWEIslEXZfr+tel5apz9hshczeH0ng6V4PCpLzrwOUpC7PATTvjCHfWf/5OTjVhyW9aJ5z
c77IlHOpu1C11oNbSTbqnvsdLldtX96de/CGglBb6vkF89k/PufdgZ4BbmMeAVOHbsg4b42t4sYA
mYbxay4Qcxdbk15GNXgG1XP6mO+NHBnaF1QviiyUGHy6LaOhJgYOuQqwtv54GN1/23xemkR9J1Ur
Conn8wsj0W4uZF8oCiHh0s/toHz0q8czpM+xQegIIUnytoaEiBmt7YDdzZ/H09F9vnw/TqyVzHM+
tSZ5XConxkYwe56ePK5Vh6rnUY2bYO31LI843HhEq40lSlF8P41XlbHdL6T5b9bZax++QTp1HVsW
BSQfhU7m6B+7Wf12ttGII0PYswUYds2/lFbdQhm6t3iQi36wiji4a3U2rkgan8RZyam9KaQJJKLf
QaeL3iAGyyXbku16C6KG7H3qj5lx2ErRWYSnNOjMH9bGi4vevPcFOB/YJvcrq/ova2Unid5Pz4L/
ORMYeB+NU6zpseuEWYnTj9Vyxs9XkAfzSv9acykCoI6rLwcp1km/Pbk+SWTf9Pe8szmN8eJ3VW5n
ZLpejtI5uR1kKqfI/klLqSEIg9aG/fuZ/bcO+fViZNWsEsVh7Q2WFYPEFNYZoAhx5f0FlxQuLSZ4
1mjS/P2au1mJYOuFUTFXAvonkDsXUIS+bSOV4p+Zy60H6Z3CQn2rLQNwSsmdYSNp+FptsleSsTPa
DG+xATt849rsaxFu4UXirqc6uzk4ER6Vbn0QaEE3V054xIgfQP2epDGr7icBCIwOJ5aX5sdu/wzr
xVNLJ1Jlk61/ZyhMoBAdgR6/OtRopyN7rJaMlsYDCsip8FmUD0IYoqpStgtArkZ07XJkIPSAEFHN
aOdJnNF9Hga0S1t3nl7Hpl0ZlnmqKgCEDeKxFrRbxIodawxkR2hpyXy/PLHRXwuom2n+5Cz/4wph
VQznQu872mDgZwTjzYw6Qb1T9g4GeXSt+hBjTWykbXcBdjs1sAvHd8DnxgYwEqDnKd1vfGU8TUoJ
hkKnm+8VbJMru9GBPEGdM3Cq8avLfaXPnWod5Qbyqjv/va78RYpZep1r5chLshe2m6FK3bdhI36v
UbDSNEhGu7uRjHW/gwqxWFjRetiui8jQASBGm/hergMHLHDPCl8OD9QITdoKZPz8w93L7PcJMbX6
NgORV4MctXNo80Xo/qajuojqVvFbzlDkKcRd4ywMHiiCK+gBGEOTeVsB/SxrkmwF/s0bQ/K8VRWm
aXFMsqirRmVsxf3CecwIDC6smN+DvkjuDNU6S27lC1UZTeGOFGWzcZAzwO0DkLVJ0g2Q5p9ETviQ
MWpsiWTmbXDr38U7/p9WMZxQB7n2S3283Wl7ZHPrKV1AepNnNdKq031j0xlYgWhgesR8Opzk6F8A
DmhAWu2L9ghurU63dNGD2lyF6ZvRDdyBoCSBUdmXSto5pLoq35UM8x6OhTi30I05DIu/QguuM015
jteFno+5gwIKeI6yq+A+iI+7eN8VmExsvrtAhrRe3Tv7Xnl8ohqXJgPn4CpXepgbUkMnTsRO5dZN
Wv4sYzIjTgk2ePHEQ/3Iz6xSVOvu/uvzcygKzdxVjZ6tuofA4sij99BNWzqcsoejH8TUZWcrM+1Z
LdKz/kD1mxO0yxtO3fezYYbRLLQkATQmbP3RjBpY6tumscu/sHSf6vVq3Xm0gqoDawopzcm2VC1k
9ZQRL/gMz2v34ZlS/9odMsT0qu//1Wgl061BuwiZyjwZl+C0p63eRvai4bzjzqEJok9ALumnU3oH
yYvb3xpuAngiVOAwFsIteHAyPeeGVcEXUGB9o4s5CCh7a6PdbP6sszPYNWBbOSRq26o2YlQOrLQC
dlO9GOtX2Bhivu+Y+NEIXCde7bUrnO31BnR5OPhNkh4HVdBu09uQcrCUd84hg1Fxcpif+Xl1/abP
9Kg7MLqUqrFMUjCYUgiAJ2WaNFxqCoM2dLAsbflsl5EwgdMxKgvPh+qzeyf6ekRGDs5ZlbolA8m0
mJr0JqGUSPKWIiiRBs9EKzi4z5KnTXGQFKoLXgp9KsiWT17AsXVhbg9m4B0IuYANMjlZaMS49nqe
1LMV7NaHoALUNLgS0SXVzawONqQvua6+f7soeVx5U26FsnUtnVxAAsh0ew8mMqbW4KoiBjTreVux
FPgkYOkrGmjN2RzjIi80bnVMRNqtQj1JwMHD5OzQRolF9cCDrptyxojr8wyVTufIEaYW6e7gbzG2
e8Yd4meYTvrs3xsnHkWXwady4FV7H+WWy9lcLPh0jYhPXDbqJp+qLYQDKO3oPmD1GGfe3DJw6gPk
p1sfF6+xwx9AEzmxQaQRcIIeiivtp/lgSbUPj4pCKRX2F6qEOLSiVbcZAa8s/yf0YDVOZbap6ONE
VO4sqs3guC1uRnEcqPbm8XrxWsOgeHS/Ki6Nkw7CuTblepr8C9Nq4k0CRwKpKHFtyfCqSayhZBob
eFPhCkzk/9WRs4Y0Ar3K986hL6TjRlFGrAZJlBEQqMEtFRiB5GyM23FWMyDAA3FBex/TtI/n3yZF
IOJ1CKmTrm+wsFBfhg9NI/xbFv6nbmf+RV1VCm76IWMkZ6hdvZ4lJzF10qfJlP4EsAazT0ag7rSA
DI15+OfAizyNy4C1+DM0QvnJDGCce5cVmzwFlW18TKV0hb9SQwYrBD50e6ZnBb5euzQbhnJRtNvY
or6J9+3QZo2kQJW22UVhK0xN+zMiQBOKtJJTVRLRdMM0FZZw/+rWlrt8xUpKlc5iel2id+ZXFYsA
Qr1PFxZr8RfVZrgId8DOvlin2SG5HSjkaR30R7ZlMl1XJsR86HlmhfrPrukGn7wn939XmJNNo+0Z
oDS3qk8qAUu+N0bc4Q7MqHM6LM4ZYM6fkchKBM7DEcQwvapX5ztSy+0/JPG5+CytpYzsQSg4Svmf
mm+cqw8PpsJBiYeSBAUYfKCYTnYTuJ9XQbTEziyg/WtneiNom/2LJFB/8E06rX3jGE31SRHhm+ZA
fnkXN6Ui4Gy+P/YoKsZtXCVJOSWTvmcX6pkcqYL35TzbKqONYWvcNT88/n4T/pUM5qC2gDDhVG+u
sBm7EjWcSwpzA8Npecw/6CwJEG6UPfgHE+kcNums1Q+T+Aw1bvOIirAfNd1K7deqKvV0/gzABMgd
25505zNdCraRzON7aqX4PhSqhoCDwsrJ/deIHbEQmTOUD+KhXhRmmif34rOgyzLOtKtv96dq5E23
WuiCLg7AiMIc1AYCiHHoJuLf32u2KKgB8su1VmfdoC51JFZ3XVHpJV9XSiP7P9E6B7VQhKHSmtT+
e0DIbWll5maDt+8w5ilimRnLgRwU2xn+Z6CMKfApdUp+CSENkteb2xMUTiIwxOMKkg9TuugYBbtv
512Bdcgc7kr5/pDacMlW0B4LhPuvxixiFY+LauMKPTI+L+je92YEVBg6OWdP8/ZJtkrRnoL4x5k4
6kt9G28uql76LCPgr+BLdEFX5U8/an4G7fbkgv2m/xcftdjpOh1bq+QHD1uqG3IM2oTGrIsQKP2X
QqW4HG4v0Li+oJ+AGkLfGZ6NQ0oZfQa/bjqa7tN5HN4Zs6q0PFpcX7yoG3vdZgrqSubvhXVf5Nl5
ycaK6o6Rymk+tFu7CaapyTk3IIQWQe4Y6+2NdHEahQLaegw8UojCOR/LziYDIf809cLwiIMU7kky
tNT0UMU3zEG3rAjbQHjxApnhkE1+uTCm2pXscJFWuo06STGmXA==
`protect end_protected
